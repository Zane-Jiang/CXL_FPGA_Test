// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jCIVsIRCfaRXY7Gwwl0vKxFEW/AUaz4Q6ukguEqsKYh0Hz+ucUEvBO4sBlp2
q+hLDts/LXhiT8eEb2GUL8vVGO6GqjRm5aOg8L4ZK9zZ3Zb63KGb+k2JhfPr
gSqNiZpbLCFCrJpNShceZ/0797BKCuKxY/wrGdp9QJS5wEiP871nLTiIZ6D7
NfurzF1mS7IcYfCCnx7GDPDo5TBu9X2g2JiC44M24CrtwUMvm4mfqe9Fh+Bq
4vfAVPHhiwC+UU2Xb9Vm9E1PPkbHGwdxW6OU/+MD52EClyJZgGrLkwd4eov4
xtQJ1HsdW+qK2uASMIVvhi1HOUW4eDv8Cz+4Yxl10g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ld7CeaFqw2Z8zBYjpxwTRYTX/jhEwxQZ58bOTP1+ONPWhegxqisAW9e/f1Ty
Aqihe3A3/OTm+o1hNlPGsX11iq9yRI2OUQ4hLegaGt8/QsSJ20FKUrSHzYKC
nPu2iX988SPh1/FNnDXWr38HR+LmHZMAnf0tT/EmTGccXITXg62sYKueyIt+
l9Yp40uR3fvpglGDxVSR7UBkYNBmbM4MvTQxXg/QOYuKyQbaqBp7EwCaBWR5
TyOWWGdHIeB8D2Gjm7DD6ONeUCEIV3miz3HEtg/sxZrV1sZpDaoMoL04kB9Q
CFS5I/J6ydbWBSC1Lyfxz1WxdTwL+Gt1XSXKc8vdbg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XjZq40ozZzRApXnmfdlY7Fg2YrRNNENX+7Wiv3aj26TIDetxv5W1zMq+MTuJ
DMYZqL04RRO1tcWrIPp0CudOFLR96VDg4Dfs1Zq+DvNcagJFZIY1iQt+yR2T
d41UOKt6C18z8gUXqCXpRErEUEG9jPrgKF9JTOY/ccw79QVhspdhxTN25Aeq
bOUSS6dCyY4kYH60mVtHiRFUwyuz6VfUIgPoFSbhlB5hFfOfGw0Hu7/hnCpD
VPTYcp+aF9B7mIA7X17jqL630VPPR0Hht4w3a+wtAGeFWvoO2UaelOBOeVHd
npFTvXMJfPrHd+LHLUmGuCM7f8j4WOLuowwmjH0CfA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ex8PChQUgwyzJDw5nlvd9S1bm6f8w8B5ztikFaft5QaqXTgFxjCAG15wNt4J
ySRdANUywEhktZVOaZElTldLS7XoTc/IEUsNNQjkdw2xbaE+bOZqntzPdK/x
16LGC7qTILi/PptVj9cNkrkeikS5152zSeSTssk3jWhatbpx9zM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Hbr0HkSNbwhbcbPtfxCJfvBcKgUc6T+XKDdLlFiQwrm4Lc8aF8Uc9i8k06iP
W5lv6srRa2dmqA7RGV6riD0LKtZ1/ggO2kt9GdHncdR6yAESNMmge6Qi7hvw
bKVqevF7FvhJnoHGVjsNcA/29IuRbWWblBiWdqHC3lekJvOYXezzEhgI4fIc
ZuvqCM7S+LczRulPtgevbpWWd3G14nfhZjrwXhCH2Xs4G6kTgvni9uKAP+ap
DQxkbTtpk5X+PizgT4SWgjB34KwBqMdacsUJcQMjdjEpQHMr920kBtz5rmAm
ajYoafeFEOOlCx53hQUw3+IKCNvHopEwPOTIYbXk9z/HIZ2nUZURyabSoR+X
CugR7t4fUCyvbKMINEW6Wmdle86wFHt3S1zQqag04se2JFxd9Wbqv/wzCZGI
2bzVk6Jl53YIy1tQRNIYGXFGUwjasXpuo3cYE6YYkdPuFfr45Hyi+pfddY3Y
SEfNpt1hvmVVqEpfPY3VA+3oI/GE8L6e


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e1iZ2FWxfiQsTCH/5ATZKkqwR3EqlhoUcv7at4s6h4AoooKLwBh1B83MFzas
Q98vZH1Ra3diNbRQWg835l/wZCWv2IykDKlldh8xyrrHQmzuHv1rVqdITJJ+
LUEhcocLi+MmX2PydOT5g4VKEZPsNL7WWTaVuxU7Vpd0Vzr8YbI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lU9yQDIeyY5ihwzN1Q+V1MBP1YSXAZg0mbIVAgOdYEswomdpAItX1HarpRb/
4P9dn3OCbrIjAVe5Y5uY5MLF4b1/9hO3vXSYunoZC4MBCqcoKHw5lG07SqTD
KpFzxLJ7U1sdu115WNtiF4HARgIOujgrj0TLj1dnAGC6izpSYW4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15344)
`pragma protect data_block
DtZg8Rw/yXWU+WlQCHSdPuURd7GxRA4tezRdQTiroXKar/UXuhu8TeflHeJs
kMxrkv6yDppBnXsJs291ER7gZ7CJf8joDcHzh33k9kYOB9VbD+FBjIH6Rku8
tgWCeyy633ZMysBBbFFWyoZFMeGX2jazwW5PCynLyH+c8Wz7aK9WrOlx9ygJ
nxMhF2I44SubzyeCQXe1fsH/EZSThWV4cUo+4pLNLtals6DNhB8UoWhO4lkZ
cOmDbxvyRaVn5igbXfviFoOe2SAf3dr5DO2twpHycW+QxAHUISkSN2bwd3n8
wD1bDLboj8n6GAyDcVF05bO5/RgWy6Bv+6h2WnUvGIX0LjR6vk0dUFmy1ZIz
p2juxa8ZsfnLXxK8hLmgy1myoNoNPT+6rAuHOILbmHmQActXMqql2BUQDwF7
PQD3/MrfBW/q1dup6Z3jLcrTy/1NByFC7Q3bPfrMrpX8zknZnFGDh10jYUe8
/lzBqmwGC3ounKalqjiVNzYP9+KQX5ErKvLz95P73EU7PoHUaDKrYdf/ZwWm
hr6bcBJqZRIM0F08PNovOVib+C1mYNATC32I7tbcO+vOXEs0IsaDvQXlmwHA
j2jZpw8kJDVUqWJRVoLPcF+cj6fX9GpuC+0SEjLYDb06q+XpgwOJk4DnDdDB
oS3/EjAeggtxj6C09x/kDTGeI6pEC7im+wOSb/s0kX+mePDI0I72Nzu3anVX
s+hRVXClQ35SDRDvHxpvj5S/3T2UvKBId+/H12zvSaB6GrtnQ20iidpaVM5k
VozbCUznt9pZLNC2jBH1lLuN70Hb5wfsT8istVyFmSRckfYEN9XxpP5lXc97
ZYQH4AftSmnORo+xBbcZZECLtHngEu6HfxYtwa/kNvQyZZ3010yRkb4yY39K
e7S+XavapZe3O2YDUn1SUnHxmCw0KXHBNp/tm0D69nYMg7RpZ6EgEIhwpV+j
+SNLmzr8wJxCPQD4bWNEBAFSlZT1K3YScZKI9pFKVMx3/3D6xTSYc4Uaa1dV
h3OjuFV41qD+vSgXX/pp+WnlqOvCzKx7+wuNOUnc3d5wx8DA/dsCx8EMM8jQ
Z+BzQ5X2Cy96qTlsZJbiugNzIKcNwNfiAGyE7SrdwDDS2IdXkIHoCrJn4Kio
WBnMtr8ip6IW6GsVBS1nLBwbPeTYXA4bJYhmRDCp0xzneuXX5BD8gtnP4gd3
m8fQR+T+lcERSQ1CyamgsIGVBhFfhIkUZ+jInjdrXFMnLV2RGGIsHuQqaULo
R9Ep7EYO1lO5C+AxFDZ19otaocHkPoej3K2LRY5K5WRyBx172hm8j5i77SRV
BBhpF2BAs9QK/8I+4jAcemi68PZqogBmHjOl183FjXu22+k58Me6sbr0m1dA
CW5iHTEH5iLy/1WqmZhUv29ojTBGBZHwSPnfNxrYsfaOJTvZ2acyHqQ5dssT
2Rl5L6NoimBBZucjlsU8XJHur2mjo4yjdRU5qQwe2vVoB0EIPfKZtfWlAsQM
JsTlFqhXDGxQnU57bVi9MBEEt3xKghmRusbhk27wP+G0FTPge+WsUnm2xf0c
1nXkJe8rdYsRNN1Q96jYwugFfjyqdmdXOZpoIkjh/1AvL4QF1uT30rwcBw70
5A5LhsTd95YXl2BMav++fo/aGS+36cwuYKhZ31KUz5mbM4PPcdEOdz6cDIiZ
aokh9OGGTnhY/KjjeBuiqo6ccVKCf1Vp5wDNZJKkOcd3UVU9TAPPd70ckkjB
mYe6WYpmUToDHPIAblJhMC+HH6IT7zoXZ+qnVeaxvMJElqk8hNUes4qr7+zx
8T9VJyu/45OzHwb1tip2m1lM4rEmDiruzVd01VXI5R1bwHFcQT4zRmmsh07M
9ABkY06SYjiUBqUSBCGxWbx7uIcMA2/zZqoMc8dllNe4i3FwOqvD1jOe12lW
s4D2fFhFZ9L2quPRybIVivZwmTpQtsi0hIc3ZooUhZnm//hqBvNUiSlt9R8H
ciofJ6lSIv0WVTMhIU0CaxYCPmnUlJe0Zp2hoO7pyhDJ5JJLcmc3zhNzoGQQ
2JdYsYmSbbobH6qBsHhthbnCcmcE/o936qR4vPDieTr6eFNGAoo7GJSXY14J
9QSO+KKhXXQgsWS1CYN0zOMgYA4g/3jg3vDaYdjJRkHh/W/FLS/UzrBy1YKB
NQBORkybSINb4goCW0DigPvd+3MeKgQ5osqyfWGI8vEYSmjbiRxSFw5TwAd5
IjPzUu5uvovZQOpudyMNYDsJXjkva7gvK41gmnR/pEWeAgKGd4Io9aoYmJrT
U/Ar3uEFLr+B2SL+qsbjYTX9n/5P4z0JpORCkJ6ef9ZWt8v8VjudDWMFq0E6
fQTNxk8zW66a+g5UUM05tIIw3hUFMNSOw/HGcBzCUf9f7VIIdN1yasuX7uCD
VoAZk2BOvhDdpBHSxa/6u+abFV8I7CQc9iMRaXIWFVMBrvHkXixWy0Drg1Kn
pCDW7OkoYawN77ulbpJecbdnqZmCIalRo6LvxX+ditEP3PqaoQJsYZ8jfpb5
7nOyt4NPXQ/7z+qckoZ1ImmJMSVviop0H37eVY9EyvOXQ66qPRN0129jyC3h
KPNg+a8WHLOGFI5J+fe0sb4LSPyWR5Zg/x0Hv9LC3TA31+85dv4hzsggs/XI
aemQNm0k6ysOUOJCH5RTrHUixubsqOugm0F4lGxxhe0G2jLBC1shQ5tS7qyt
v/bfphjpS/pjoINda+BJepW4pJ8B0bamcsWE3J0hi5fF0fx1pFwnuHFl/8/V
tezC+V6vCNnnw5MbGXwva0CzTzmJI2b6dVNF0d7p+NJSP5Lna3zasMK6+Urc
wPQLgaede+mZfn1x1/8Viri6joGfmN9S9p/xLsN1CnxfSq6EIE0/0uyiR6pM
d0GqRS4dO0GOwrXx/YU5Fw05QxWmN4hVK4ZOZLqaek74b2huIEQK/9gv8FRl
sMmk2wghEvYl2R1eDzwmk383FMSGarN1+iF4Qpy7CNdriTOgSD48zOEkyeN+
JapH/OiQDpsu2dlbxOD+G/SW5cISdjZPFt3d/52L0m8LSM/91h4olxF1974o
RydVo9KN0eNqDLJJ060ucEukpG589ubHg9zJkvujbbrzOa38oZSS+K6GaE8y
7Be6fEkgDS4PFpvMCWRZA6niyayVQ1enUKJQkOAakxCqqxT54bEZSi64N+rs
kfsGQnFJ5sLO1B2Bjj5b0TX8LccRBJHo1b0IhG2mFt1B3rjyjc8viprYyL8b
yqhaZq1WwGQPZfz/ccwrdFzE8+uJ6/cU+TEMJPuLEL42QExSDKRbLj0ihzIU
RD3UXEbcxK25UZUAj2taza7Agx2YaZ+Hm4j/a+KPFYTrSzAQ3Gp218lfFwT7
0qNpjbBU9vLG8jV0pl8CTay3Vbqh4k/8BbnbvcFAzgoZsAl6tbqpVT4Dhe2G
831Jj7Yk53uvbb/oS9FnKo645cmg7x0LKJ+OtU34mTdwdbbOP+XKQRuCI30k
8C74UzeBziaW3VZJ/2JW96IXvR6KINtrlLh7IKorAN5jH+q09v6XsYBfWLwu
AX23yVBLTviDooc1ffToy/YMq5lFBOMOfeAb3VmKwhUSgBOTunZlRnzRa/kC
IkGINaJyDMMmPukca1w3d1r7Kz8xH4pYDdevLOOPiM6M8ahd79XRG1JHxQ5I
DOPh4ZQr27XBRlQgz70Qp9f0E5TMebvDaVYkT0w70nULNrjXj/04zyTLpeAX
jX55O/g83tR8jyxBWxLvf1/f0AMAWL7sxWIXgX3Amci1c9jnAA6vrURSVmb1
guqHtn0Rct5emR5im6iWWjKZRmmhLVEXNpiGQO8JDWZzK53xNK4bvEljDfKG
fOlHPuzbh0rAPjpO297GoLkGoNoqL8VHfu9WwE2gqCRAdQymIB1Uh4wiLVS0
q7tSOFk9acx+tcyNIz3nmM7snX/Gugd6+3T+D8eo6JqzI4FhpQX39/GzQL8Z
0+cuFigq57JiD8Wcl04Pix2JOrOGG9Dv+MuPaY49pxDKMFp3po+XMjuYsXRZ
quqJ/+aTE0fPMqM2oj5eLqFTAVobGlE5vZeKGqcNn9PStJvMQUKdv4WU0/u7
9y0rYtyBm+i+w+lMPqptmw3OGdjXi7vmP19WbfuI8+CRKCGTsK/vF+KmWX3U
kx5UDGE41C7zsnIYkOlBkIVzvIRpclGgXzIb3ymTLyG+pINDxfjbSfFZcjmo
YfEZeDXNnMYiMAV/nccRhRqsjkMvg3qh7JiNvGRgXfbByiTQkR7dssW5mQ4T
4kmwBo87ORfo1Z6fTxbOU2ciNhSiA610P4m7tptQ5XaUqe3x+ukGeKDWvAnI
FLRGBst3EYZahBYIPoR6SQ6Vzis0PnO73m+eJ4k6/d/tYUEvYFxN9IgZBsJi
TiciDjXhg5AwoUwa4jsvaOlHUSwWHargcPNS9qhH1RfroitZnQs3DN4FU+W2
AAKbA7O++ybiMdH0N/31RhYDZvRYGmiSMNXsP2S4Bi7TWgNYxE0zBZTi8D4t
4L05ZOk+4inyxx7prlN/q4wGoJ8mpuZpd9JTpizavaloocCrcew1Edt79iVq
s34gyU+t1w1i2gxmZ8nEaWSyoz/a4NTaktVg1wdW/pS0VdOirIj++IRs1/GL
ItsDxk1X6f+73UlHq4lmY9IAR9mMn7QxhBhG06Cq+BPNC7+i/TFgFBPtfe0G
UJDyr1DVbqwwC5txCCeY+KXxFBBkxKUlLv53ZiWDMLOMXMirz7pjy6Hbvf2m
8W5aW489TDrzgo61o53MMxu5Sv++R0GjWYPNn+m2GWa/LEL7XmqbGtUHEQnt
WncWLwB61GaubHug00FLR9KZmkJPpOxm323LFviqUTvQbup2wNSHGuRc54Ki
IO1UE81gk9UU9VYtmVNmkwsxEYIxxLHvrh7VChJ/xMRnK++r4ZzHV9qsnt0M
8ylDnuZI1MfZmqezuPd5926YrgQwBxUumU3+xWs/Zw5T+Aui37tK1IqMAsgs
VQpSURdRw+D4o0HXhhmt9/d1tENjuemJM628VmX3hy1d6KrOgTvOlVqBHEbt
7nUSmOtog1C0MY+ERMv/a11osjnl6AITveX3s8gAr4YXxDJG8hkPaQd9JxFv
ztNYccYFWBrWwxPSLKZ6fSXYwFI2Jjyt0yovHPqpEFNCOanfkE8FQFiZX/uA
qeLZw1AQ67KLyjZdvMAaZ0y8bZ1sOHhvIDBA4gMzdDejpfIiiBfcQKFXw4PL
PgUP9A6hqF5t6v2jujbgEyS/62O4U/u48MtVxtrZ6D3ukB0i+zHQ7Oisc4on
M1/G9vK9/rwi+Emiv+slq+olywojZsvNjKNS5gHN0CRXr69bsO8cknaFolHT
S/0gC43Bxssp8deuPt7xg1XlAkISdncwwiSqVpRdTMyFHYuzYt3XaZF8rQxj
UPRmZGAz/oSf+xEwFVaC3O5YZjY7YjwUIwf6FCe6GssVhiIWvhwsx20iTfKI
KsCbhHUWOr9/g0gLdbsJI4VZqsqKgNuF9M4UWeJe0htUyKjcMowrRC5oZRkH
1NEj1IG2YxztcjUI5XCZqoOzbC4LCmyHZG0RJZ8SvoUTRiI1m4JwyWYz8x1w
cHNfoWVYvdb6R9TqvVI4t7QrZkPj0YAaFLPZ7Nqtcuqo17dORDLh3ayz0AVC
GIyHYuSqv1p8SmtPR4nbiwmm9ESjAPCqPSUS3VPgMyKm9UhjKXk7NVbmQ0w4
AgGu7XGljkBt4YB83DXisbF5uNMILu4gkLZ8PPuDYtGdmk7orXkgzZPWwhVj
etKs1aZLh9iuyQ5kknajk44XVwsmuyvhl0x2oTApqPIuQQlSE4NwKvXBNW9O
W+LjhxdsDNhjEFyXVD2Ha9a28HBEpnKYy7oqHeUx9f8fGQ4WaHDyiWwY8qXT
ULyC6eWKIrbCp/XjcZQDh56KXdbIHjZVwkBPxgPWnrMVNrQ9p1UYpXGcNg5N
TJkO9SS4IKv/UU25/DzdbvxBVLyVcgqJcHgWnOTybty8V+0ycIC2qJb4e34Y
acFUxr3u8TmNSsjvXVrSfPtXrqEI5/vuB60YKqi/LgX0funENPqCTMMrfREB
aQWrBLG/FSJg+hAOKF2TBo8AQAf3l7u7tKa40vSliOA4Tsena8UQMbfic38C
GlIWGGqBh5T7Xl0pN0HrzNK5PiWKPKvLrIgY28NWJoPKb9cCT2fiHYJLFwLI
MqGpmCVD9edg7YjLyXP7qKn/XAT8JYp+D5e4nXaZIHjxuaocAY5EuH8c/Zcs
YEMhx7/gYw+FB0PZx+Yk7Q08wFxxEBGM8F4XOMDKZdGjd33Y1c2JQ1EUDRWy
Bu4Vlm3QdGF4RyUjFMs9lBIaWjoGYyJdlzGDtL1O1/zG9+NPXhqSPY/RN+nK
Veo7DIdcs29Omjc9HCbJ6l6j70g3xkZQ8dv6GixmGzu/ggOo0zuIkudv8chQ
IHoHPnNrs8NoruqauX8RzHhHX5wOQRRj7ckrUhnNafX4Q72vIjbZDC0x31vP
qoJr57P4AFUvXgAYh4zxbshom0y9iJ4YZn9WluuDEXkcmHjRRa/Gc7mIR8cb
luK6El8jrbhP2cBPMr0RFX7Dz/alTXz1ED72MnkqqybQp2HLFEzD33d1NWkY
eVM9SYLf9k/xAxc4MSmqBk0p7CuC4KIcV21vNhhBnQ5TsPG3fdT4n70eipDp
Dtjd3pVb0dTfuAf5G4wX382edC6m+9Xh4aRMsvmk7vRJkpbm2PTbRgdfGuQI
D+Y3zHJIigZKJWs63AiIWMQOTlFBWT2v19sL1dXhc8o/LQe3dmTrinMWQEnh
nKKkr6JdLAAqKzsLpc32t50Rllefy5jCE8YIviG5ssC3GPXD0wtN9KpXx41T
qDTQZcRrsd2x8Av6NVPJcLOK6ucfrt8FzVPTaPECXWxytNsAtPhqTcI5j/qU
NHWjtnYeb6GF9asdKl0ob8y0BAWgVCYx5qSn2qBlAtmFJT4BTiKl+uj4Oo3J
XoUxj7Sqsnk9d52nXHmwc0WiTZFd1eXtnjwmND8D8pxf3F92oTvDmRG0Qmff
0GpxOeIYMTg+z/34CNybkVzTRf2kDOcXJDxXb1OkMroIlo+YGBYpu0Q2M47Z
fmjBsBSODNH7YEJhFNHAChTIV3ntDT65O6GMNQPY/5HK2EuqvC50j8q3RIK5
4DCT3f0fTcOKg2zqc7jDl2s93atim3DAqbY58QYGd9sgi+HDEerM9yskrbox
3tKc/r9y9rlfDCR9Dfu3a8QU3x+tVEW/6yfFgD0zaU2IuidP0uS5kLUBlS+T
A72Ekug7SX5npyqH9qmX7PEwgRtZfwbBUSW2UqNVyvifQh65uG70XQ6m3cWv
xJm19MFsSnSYWg0qFWZB5QWXh4FUjejmK2IzPLHSO+xNj04feYS2EyhOdPdF
yClD4ZsldI+wbnwbIWDohG3Zcop62g67UIirYlMp9v0Z1Nxhy2+JuiJQ9nn1
tSEzs3/3e2gSFyUshMAH2EZweTpRf0gJ5QfzyXGBnzNlOhjHEO9J/xpAdIEk
ivNuIk7CEo9K4i7LJJ+e8H0HcbDAYm7cCsJ2tnQakXqDwAiYubPnKJWFGUq6
TdcS6kQsmowz3ji2hUOE70b6aiqYs+N7v7WyrW6SIZG6PYNQBRECxRriCegI
AtSqlewTSYD9Zs5+L9XGCPFWkH05LQHdS9tURVukGgoLJ/Llr1Zj7qHiwAfP
VzLb42CZA7bmaNJXAtwxRoTFbV9sE8CaIfEb5V4ctTRptwfD/ekZ3FY5ywn6
JYJN5CUs0i6oOfMTQFzMpsBXe/wWcZe2JJgeEJdDRrZAtiImUDbQfTf0NhCC
mi4c2HGdxL9vSRDD0f3NLVyLfOjrpAqb9TzXc2+tEoyDE7QQxTLQ32Z3EE6J
5QJ0G6R4CdWVzouYQiGX8Ts0Xhj+OOQrkUPBWM49BMecwHYVb0Ef5OKq/x86
dOw+0JZsw0iHhdY5QL1HfB8tyKfzep/1BeRInM0RmXaZQMhAGrjAd5w9WIas
w8y6cPKbumnA+Xw+PCQxIfYlodRHLfzjbzVgKxIYNA0qf9ZU6+/AwWuW+YNx
BUZMsXeAFFyFX3pNSfEbbZQZ+GE2oupsUL3T3FBQB2Ce53ULI4ilaq4zDG4b
Oxa54GV1Ltn7yq4WBYx3rAmpx3bCUcXTzxXri9U1Xtkoqfboz6VhobxS0eJF
u8Rp7GdHc4D8Z8P7TGi820vGPJs3ojFAwGM38tn8RDP/xNgyoRmKDcgcDfLw
xns4j3ACo1kbXLle2hdfAMK60dzq9B3JiLRAqhXa6R/7sKqjJxyJRbdrrby1
kgtjupcJ8OAjuO1LU1Ztt2VQudV5l7yf9qppelQepo/C/CJ3Q5QdHNcZhXVp
6VC0Ivhyk7s1/fUlXfac2aTg7JbtVIMZruK37RsV5csSQ9C/bG0qQL/LuliT
jXkAqIJohJjsQpn82FVGbU3xi/X/328a6igSIW/Wdzy0z8esiVei937jCmIF
ZQXsnmobSVyU8vNoi8gclpS0Sj1h54vviIGox/sS+23a2pVhWNaTdOrsWY/Z
A4Ld99iQA23+QZUF45rQpL1ZmhggETLwkxnRLgrR2vC1ewfgVVMWbr9S3EfG
IxbdzurRE0C2UGsAuLv9PaUIjDjArhjl9xD8jwVVK7dAOk6iUsOVmo47qeqT
KvrrGC8btWxVhODzkGxwzo4NiLDB5NK/O0Kpw4pvBFAvCUwRRe2qcW6Twdel
RHccV7IKlsJLNsg3euICEsJ8myN29MH+SZKRgEWNOdju7EhbvwRxEMHK3adl
UxoyNsKk7/NlO+c9XqLKppmPY3yUyV4jwnC0ZtKEswg/Pk3nBhu6dR9OpVnr
9tEcO+VX8MGg/RvatZWy6ZQ2TZ3+rLWfn4pz8ChdlQhlmT9RRu2oP1mr1OnJ
J5JkLi8otDzdKK4I6nWNnr0TG/7U2wQ+JBU53+xHf3aZ5hT/9DWwuaXRvmRY
vZNGj6P2olQ7dk5wD9iM892kDJH1EuZZcbmBQfOC0RlQecl87Ymu/bKOPo+S
4Ce4l5FVorHT4D/6xY2YGTrqzSHf0JLu87F+Z968rjDfqN+8ArBc1m7BgBic
ri5U7/yUK5rcyjdOim8Og4ACcTK6CaJ56BKvCXLnW4gvSk8UL3qLYqyug1dx
XV05Iw7yuwq2wssplJc/2H9JFeUqp3N8eAsnpnp8Kk42RQyGXwg0HW8rL+Qj
BOF31m6QYR/PuKEU57wdvNf+U1HXVmSvQpktH3l+U2UY5WhbUq6TDb0sbbx1
ybhK5UWguXAQ8kCAuK4cfF09feTWyO9weKfdI/kYr4lIjqP5pxlIlc0f80IY
9H+Qu83UZQg5NlFB5tPtS+8zFQC40EH5EyVDR+HI94fKzPWA92EvDn6wzc6O
ADCMx/Cc2Of8HmZNirXzxTnjMq7QQa+TreHVQxEHhHNzWb5L64e3lUURj83H
ZQNoVAHDgaYG3v/rKgkZ7tHafSdKBzJUaaHSKRyHVVtrsCv9HaO/ekQceypa
Rb9HlLK0n4Q0nRKkwABcRK6QjBfLoq7s1ERzrNoBGkmeVqeh0lSEqidGuY92
x6gWUe4BnRBVzGD27Ql/wUZ0AtecmTCHJ1zS1J89aSlI6bvfT+oZSKkWgubv
KsXEs+7oZJEAVnW6Xx/xDZKdxzQBmthK8xc3kcqiQ1RiPYFjwCDiQM3tsDWf
t2Zu1XZqiT9JQRjX+0XgyRkm5UheFCxbuiufzQ7avgHMB4dvqg1Oymq7DbxX
BzLm1/BfLDV2xsndGEOHMYR+AZc/StIlxLatebXYHgcc7c9q7MBI6ShAWjqw
L504hzu5BEHl2iWIAEzprPgb7SAwaOjEfiHu8gi8pNCq9MMpf9zAIux4lXbb
QKB0R35Pj7ptLOdVmohTiJvZkHTA7BsVayVfFB1TlvIaudTF518FYr0JO7W1
/QL8lJyOt7IGP/6FRt9nmN6hohIwzS++fYzbRUiUizVMFf2cOf8Wst1thjx5
I/W2xerDVzTUSDP3g0JCcXF9UWtX7JwrOt9fLMIYJo23cIGXD3rP6b8eZ3R7
a05fqyCRbqFQ50SJRJm9wcHx7WKfg+SEWWA9vpshtyaZr5c9Df6RVvlk4VtR
YhN2BubulK4SXG89Mss6WrvMP9yX4UVF3XWZTG3f/WUzYg3mFeFrlo/RN84r
Q1b6+us0jN8CBr9AffCQw53H2m4BghHsAC74H1kw0N5WvyUfskTx+AXkT3X2
nNTsYv1oAVgqpB9Ygqrr3NrtOaLawkr9EGpJrTAYFXFUZvX8DkxyfPKrl0b/
bpCb8DNdwRM0TDlj8qo2FQmEaTkBr+fp5v1XUL1Ub5K+szFEP0MB/RJ09pPe
Apfu1CI0NvD6NHIeEqk62DYKAHNgn+j/MUOLHf3R8efMWJWuK2QpzbkejMb5
k4XajAa7GuDIs8DZNhVZU2yWIC6U9VmMDnczfcoc8rBkIZHDBU329c/s+YYr
A1pI7qrh3zfjAdLYc5D2A++gO/g7NVVpIDhUMXNrzZnxfYZTtdTKiwg/wpRG
xe1jzWHK0yRgf+5RSBlYQ+smslMFFiZ95BTO9F5ec8B1bcT7J2b0L6/RI8gB
qa8vsE6giBR9dkj2yd4YDFv2rKM23wk2+Iv+Y/alRUDvd6aBvMKyFjbpQWjF
F3qUGa0zF5awSBoHVeS+MFUBnksyi4vaUaPfV/ayeumXdVJxRZZ4gWy4H6aD
zyZmFA8j2iFV9/PvkqTn3qLdnNd9u0oRwECafZiLa2eRr6PHsS5yKs1vxUqO
kvfAPVBsEdZn0GROAmzLFr2ooFlmaTDj6LYyjX0KfIaDSRHb2ygfd43iGc6V
dMzq3vIQJuMfm3ZS8vELhUtKr9JoYbuy6gT3zFYjoUkg/gTOLRUizUMT3DgU
rNNaXtfWWOutO6fSlnRLfTu1FAgmger/pXK9JaVMze3vP3ay5jhxrMZ4x9qj
EzesWA8ufg9AWjSPfMAJDmYgGb8YMaviL5DF+MuxNe7yD7OOf1JQzyFR5NV/
4K3Qyg7WnV/jelGridC+ruKtzoc4EIO98xjBCRZU8aZOgyT/Lu2+Ibvv5Zr4
m1jQKlsnC+n8Ve3Ae06sfowdLBVZFELShexSCI+L9YQ87I6SV1wsfshYdjVn
e0CUJg5W3oTwFHxheEjdqO1S8/4nw9xf86wxqVO7Mq0BPWxsoDz8cW4ONnQC
1E6NZXMwOz3LcFQT5hik3K/2c7+b6e5KlcakTPIS8JcDuoK+HJ3y/8Ez2G2V
hwBw44ZKk1kWNnvsw8/XrPgoDMth4XopJr2tKOXa/TPchTgpLnZLG9nlmboH
Cb1Ca5hYNw217nvePCdmQPuIMw/b/i5FqnL00bXWpFhZxeW7dfcEfwefyeSw
qnNcg5cUdBblI6kgI61dQt+pi04yAW/XnmpTZddUz898+CGktLmz3nEuam3V
rpuLHh+kMHGUncZ+9rSm9N7U8ZdUCway/YRV/8wOZuQN3l0fqRVkeMA3rwv+
sYPChJMKnzevJgWPC8Yn2nQZi+zNge+ohviy3K47NOVdgqvel3KrTmxUEnWv
vyZ0bexF/WrOhJcl2aWR1Jnl17lkn6By6QUo9cW/AozMix7K+aSEshyU2cJV
6nOvI6DGDLrDP8Vj55kYio5Gev4aUG6h4cI/MfOIYWYpP3+n7znIJ4/8mhG6
5hWvKSeKPrUOj5f+lxrCLEWTthPahiY1W0/quKoOxtPFOCQERGI8OB6MfJoP
1MkjPdkZCGsVbO6lFj3586au3tloVSgj3z73QtzutDSd0D32lDwjbAnipz8G
VPol9St/VXpY1dbtnAFV+t7B05oUr517Sar7yzTSsDeDlVAHTN97BRghB0z/
/vc8duLJTd4Xzz7jrV5/KG2fheHPr4Y3N8OQ2DJIUbrus+r/8nra+lj7GQdg
OX4AL5ApRcyju+CD0VcNKKh18vmjsOaq77Ut8GPPSwJFfAVd3ic/4BMs6MqH
CMHdnigquqOJtD0qKnDMP7DEixmAjSzisu4+xhSS9qR8hcYYsTgy2dlJQWio
oXfhFgnhJ4exhZDOlgUjhVmkXUTU+lsVMIznMY0meldb6+gzMQmHcobfrSyt
WvDkk3FIEF1JiOLWU7JRags0AP/dKUbKp1nn+5h0l4smUy7CZ/+UXx3c7K4M
2sH9tw2d6j/0ZWwoRFOkg3rEetoX5P6Noxb/ny3O+Rk0vv5/AoTQc57rIH3m
JjsjFy/TFANDj+K7cNKQxHYFDMEMvbom/P3m4Uxl9VRPM9cAyfluNCenwHTe
hBlJa5UfJDdmA6S4/f1CYlNNUuJ4mkc6hYe9XiahHEE4QgScN+06EuG4+OQ4
GZJjnQBl7fyM3ZGO6HnBoBA5DL+jvg9PklQorEFbJA3P/Hn6oh2aMNBRECh0
7Bh7JuWnTxP0G6GSPEpm36GxApYelroiPq9+wW9jOVga+/rSUAyO52p5WPiA
Xtwt2udeqH/Px3t9etsY+SD6ta3M53ZjVTS+B/9UXUxsj07a8LbMJRJhLP2r
1O2DcsQRCfPVoZmI06BRwD65mY0KHsPvaoGP1Zc7SW0MZL8Wd/eIdgqyRTUN
qm61ba6B8P5sssb7MsZASkp9XQjaTyobsRlPBijfyI7uxGpfc+iY5G7jYUSc
J1SSeYP2l2w0uCYhKHw9pf9PIEwUJNP3EOygfMoIdeCTUlGrVUCHgl/OHg7b
oGzrjea09YITA9Pg16EiiykaXtLWgaAWVKKrTFdMVPYyeNp0rTdsCUd/Of/7
ugmUXeCtZ9xjHeIn4pUW0A9ruLF4WZtzdFPolSHMhgOsWt/6dwZbT9FR2RYA
orbKW4Dir2eGwgAVK9/DDdIHuXVbmYjm7OziXm3VU6rT8CZXc5Du+s586A7h
wwrNLq92eCTWRVYDRsJ5pcCzvLH6UflFd3aSF/kt/lQHgj5IETrdiaFi5kdX
y3fZWbPFozi0N8sWz6Htgl7C7reOgYnR457/2WLz48QhX/JlEscIZb1jHMxv
VI5gtJMyQ0YqG8wekRdvSuWqokPCzdltSK4JyeBM0HmEE2/4c76n0nCP9xHL
8TsW2nwf+hsznj5KPUzuOqxR+qqNwi69OJsgx03N8qtFIRnr3wzxAy2Puy6x
k2FpdTwMmDcz74so3FGU1S7dtsFH9tBJP77HnDrsYip+64gNm+78lvJlFmWA
NXbKDOj/yeI+Av417BJByFqO3lTbXOhraf2juY60ZoV9qWunQyZ2Wj6WGTsi
rxGRsPPRzXIicI+qs8njmOgVp8d4ij5Vrj/VrmVxBN41GLH8eVWO4Nh4zE/j
vKbUpCOu3NJN2wJ/9DjMjkIpUxjSiSc0asE611Qx+mjMW+hVsOXk1+SJjoaN
9CQIKhEJRXieIjAw60xIIb7ZSjzXvMf94seqf3/Ld8DWR7S5+Ikoznz5wwlp
GRUuUTGgPoyUk+y5bQ4vPOuilCeSH9pDuFB3AQ+AP0dTJm8sR89AFdp6k3lx
otNGBxP2s//hZD5QArcotqSp0t+4iDdZR11NvjxPDxbaF4qhza37CzsDdoLx
riQoXSWZDI2Wn/B/ShlzPpbX8LrI042fCPfUKFy01KayqffT3v9mTNAeKFq8
/QOGknkzMHO7+Kdy4tcvA6u8BPowtQWgReg6v/P5XfTFEPkhMPEaz6jMRD0Y
K16fYrr9UMLiaWbnfQLAKN6yacGAfEGydfVnCMe0nLAsbgU4S0GHwD+J+go+
a0FBRsWH+5/pwTRLiNK3oEBzp7WVw5lo9Xu5uq55HbK2xRvj4RVBY3WK7Ihz
nniLzi3zz/3vQBv+DPKZlV6x/xFxchWTxPa0Mw1QTfa0ZaaiUtFcqWwb/jxu
vm5AukBPVAXusHZpjUTunf2S5QX9FUJuWSRK0SeDjYHrIQwMKZdUEKdbmQNq
LzwAvwRXSfW9rQDjKTpz7U9iWb298WIyDT4C81LmT+pZM9VRTN3bCeAbd5Gd
wc3HQ3PHXCvmymcoOqi6BFhSnWq2apyP5EM8bzoLXTCcC3cLL3Gti7+P1sNL
GlMI0xpqqbJ0cJyvo+7PgZpPe3wdUV13WIKcml+ld02eoFbf9UypGYfE1/8y
7Pht3AzWn39K9HkoV6i6lbrVP2pgClTYaKXETwfbrvjwRpwwlq15jUgWs1pO
TuyasSAQ2R7wZo+oxE1lwwjXZFFb5FVrdm1ayzt+qiPY5CBFoZTNOIUx1r+W
+AHoaDva7zhCEighRRcG8VnBdalVaUw+VJi0y59Gl+kCMaa69BXRTaW8NvXZ
PRPgVAI0XFTWpWNhGRSn6aI4lMso7NNhLiQjvYg98qwaz01hozASjeb+7iR0
4kTUHryyNOQtipuVvKpH9BepzLXQMDcy35UzoSZKhRWYvnvqv1L8qapb9CaW
P8GLt9mu0Cf2ZID6gvqhzgSG1s1IXsqbTQDjgfKZLmoRFNsw+vCwTijuj/gc
sEm/JHzf1NCI15m2lsXvuX0Q9om3yYzI5Xf7RN6S7Tn/Ldz1ANV+81oqYdMm
ajFqr01LaN6RtZ+a0/gaX7eJgpXzwCmbK9QFi0j/sVKF0urJwMi0j0G0k3I6
U5Rf7bnnzuwzwGW7HLRoKCL6VBoX40nCuleYkTnGDZCLSuYGhJ8KxG2Xz8E2
ZIIw6dhHzBVeo0OyAHYttlwZm/LHtB59bLE6K8SD7kVm7x0/+06RmErJ3M0a
6uM/9lD/9PEDEp0ac2T7Qwkr8zIPq1lUUjpnjrAoAAZNiv1Dd4RqrUdxbV28
P9yxjfquZxDqrw95UC4IFjTxlIj24Wa7W1CkxSRsnIp08ahcdXnAmeO4ssrY
gVdFkEq0CIBGkXT7ORsigib7dGMEcoyKiZo50tT1Cervg8jdKHunA3rP7JDW
sQRNvH8QUPGUp5qcQSriRnPXaCKk73HfYG/3PwBCNF7IJWHO5fxyeHhC17ma
1mKa2ogT55cDHMC9bjojFT/8RGISHIczqkbkF53dQLmRJbYj7+KRvLMA0aJL
BLri9o1YktSdqwf9DNeotHd0jhdLn1FS9rWaYbYXw+XwQjTaoPVX6P/0bUXd
9w1p3yFUr1VMPzAFXcBSBDV+n6lMC2GGxMS9PsPs/mk+puyhgWCt2/ABJJPr
phtOHG16cgc+4m05BgCJH91YlC4SYadQrnlHxuKWzik9a+02ASICNWoJxFdF
v254CYx2tEz26lfXnYtWUUOFMpmN4Joho5qFKZU/IPU6csnxkXPQdYww+T8r
ORb2AvT54tFfSWNmeOmZaXgfsJ30AgL/4GfVxJSGdEH7Ulq85zPJMtiABsij
cSySkAHxdHoo0qC4IzY+JVMVfnFcTZx7t0oAWMhZEnSfdxbK4iFffE0U6jnN
+jTrbt3/RmIalY24djnwSHSIxV2SFVKepg3BSjlutJLeD8fWb/3uChbIENf7
6zFr6Qfy7SDtK0i/vXtXbzLfW0txAXrFGEoevotnmpaf81OR+tAH+bTTWDln
NQU8Sq1IMhXb1fFXL3KvRfq90ow4ZLt/nAcZOVP2I+QcDttFXfOikVMMtsYB
HTJ4YSgVYFWDAXKy/DuLXuTKY9p36pQeIQQXOBUIv7YT5zSGprftwhdvo1sW
4/EoD8pVaWpjxBCX2KwvrMVab2ZgV3LcaXE9/+23GCmdReysSWaAoNm0BlvR
FyxOmt/9wZEm3p+fVFd3WcxMTt0fYvFFt93MCjnw18Gf34ezvexZ/zQ/kYgi
J0HN1Q8r1K1IFuRuNF3J2u3SKbpQVAMcjMrAdSBwcrnneOByxu6R70oex0Cu
A94z/+fr0CW0024GQ2TPHaea4yJLWsphf5GRJ2FUemd+rOwKoR60s36yMWmw
aKyg9W+0nKYGyfm1KTQ8CddTzjYX4SLJdoZIDbVJ2bj8flFr/hu1fWrRPJRt
QCT0Q/w7I3yvirKY27/6pm4kxotyAcn7Uor4O+OEmqi0USjPuFs2mN1r06yc
27rtbqzxZEIAhsRt+AmFrlt2ZP+GMaaHWkaKnzv6TY7bxAWIf0Pb9X3w9VJR
S9IM3ij5ws8VydotQF+BatVE+9a9ZawsdQXQjlJZnU9zGriflkXfx+ZYORXO
oQ0PyOfcFWXFFma2tojsuukzB+JoYe6MUvSUd2YgfX8g1ntH6E1cOGA8S+UJ
AUMgvMupS4mnakkL9E9K2cfMiDLNFT3rgQ+Tx7r9pMxBuKo8nYhsvCHXFOsp
dmnY1eCJzwGmDNalGnXmJ2nKbCqi09Uw9OtcXsDpnAruY5LYrw49+pnB4Vli
ArLgQ7U9AwI/HYRLYd9CUCDjXdN5EZdDfExJAC5CRNn4c2L+gfl91bzgNbAX
C5uCf+7JrzZQmWFkQgXd0kBB4EEF1SELM4Mb4TX+kxm3zRZn7JYowJhbR0wA
qv672T+OXigRszGJXZ1kVsk31a8f2AZAYDygfxLtagSRj0QnsJSYPiX5+bHx
1aZAO5yiawStLAOS8cohuRduj8PIP/Dw5C/2HnwB3YOL6deheTylqfgoXjk3
tOfMs61EU4/q/LXzl7qabJrV+qLcNw+VsStJAMcHUOM4F5pY+3iM9qeLGtkp
SQMqFjnzhsA25S51qbCPfseVSkG7DCA7htVNZeTtrgydMgjRv+AC7ehWdwmN
aamiPsNdkfBE4tpIvepIVLUdHLkdPMusXe8LCmPIGl29sBQ6Bky4PMrP4CSj
92GWexvQdYBOQ/rBsnths7lZF1VhCo3JMomGC0VR1fO1HvwtpGEFI+bjGbYC
DwgWhxCJT81wupPzRaZwV9xkjyDDxockcE4l7UtYmvHGesPS2mRqR4RODPWW
ER7wIFoMX7N8kd2bZv1gmR647rNQUI0+kdNs16lcozbDfeaBfQyHzf1XhnPe
9eurXUS6eTBpaB+7NOKn1Qkw+yh7LxczpioTs3LrdSEW/vDWjrp5TQYPfEuL
Gyp9hEF52NEvj9piVp496WANaIj7RdTV3hnvIEq9Wz5ePndz4dKIVYg7tbdB
kzYVNu5Yk40IygYBNOakzbAFI1sTW9fLGUBz0fZwh5GyplvJ5hT4IpNUBB0r
W5EqFoCJt/k7DkkLJ35io/DOnpzGQ508koJXILdvA3vSA/QsUpktOXNs7pLS
8vYKDengEeTL1Hs6hyksNvMK26fQH1P3Gb9PCMz9mFBvcnkvHWiNQkTgU1k8
6gM6qJ2x8Exa5vIfZes5s6hZ2qq32wEI9DSj4qSfZYIZCl+xdzSxzWd4YBo2
tEZ98Mv7dBXdOeOhjxrkdP08d0fMj7EkDJxnqjsin/lu9c1KqyouzmGAdhea
VbN6hEsQgJQ68H8b74hSqtSG2f6BATRpJSZUz5gXj66G11qjI6tUsUPnlzms
rdI/b7viIMda3mtp5RQOlIbSz8NDwM5R5Kn+CKYLJyYfvmf8Do7WaaRMegBa
oQRnvrb7YZbZeedXwNGX5qC0KNAydgCTLaFtRMTJGNOM3WMQ4pTUr7kGO2gZ
APs6i7tnrhT8l6HSh55e7bJ4OEdLczVbuxtmV35gRdQS9kPkBzhf4FVnDmLR
PlGH62Q7i8cs5xS4BQphAitJz2QEDJXXDXIkhJn+7J/jsXmiOmIHItMlLIGz
NiLMXPMkwPJX5A/SiMZEdR9j8JHzOc99EJpg/iHcGMl850X3b1AaDRR2r7RT
GkXw7vmHSOTeBhreuNclXgaMDqnNzsmhQdW30Zh6rGShmGVCQlvDPypSurpK
nLAIBi07igBrtZtidJyibSzdti0kGmt0CYFCQRhAtfUC9CNDPASsjVfdV6/X
ci6BizNeKM1hF2IOEBG+ZTAsEjcEoAsabnNky1oqJvXnY9XloWWwBwzTqHDy
53mpwRMvpaL9Dtj3qrzv0Ucz7jW5YKEAdiMmuUHH5RqECbgSg2AHTS+ZjfnK
hxsgz+OVTcOwvjNhmlQcDCtaHGQHSCgZiBrdDARDc/E+vk0doCUecUyL2KIC
Fll4zA+NzJtfrcShA8+orQQE8RC3m20L1kvIzC9VJitvTa5Kr8zVWsGRx0zV
riPU09H+kHdykqBs3rwIiPv1wb4QLnOrPDEueiWe96PU/y/S/izH3mnjWDZm
hMeT+l2oMweDKknWrzf5S5Q0mMT9hgVvMe2tEbReNEHvAlBf1v56vfeEZg+W
8cVrO4x3+4loLtJYH6nlXcGo7DKGGVI+m8TOfvsD5RnibiYK9ShFWusUmv6B
+KuAAyAL6HUUldfpnsEXk0tK753yWZEWh2FkmdDkYNFse5Dv2KJmDb6FJyRe
8HuebQN0YGwv4j3RYekLOnMufmbDHSiO29SR6fsSKUXXAPV1M+ShjjtgiBgc
14KRCVYgaDbYE2UQbN/hnVjKWbbZ+rp6WghSjjG8fqDlWWfKndKNce8Wou0O
EdH7L5rHCOGl8bNn/8reZe4PDBYLtw+UQ3lOpls4VbpAsjCtafG+QWhTUN+j
V1fVY8bVQw2LKEJ5oOOV83j/fPpEnyVGa9wR9lS49c/S6R0sV17/Aw8LmmGv
CzT6iU41/gozJdo2DtWXt3naJDuGQZ0Ar8fY2d0R4z9HA56pyHYDA0YZrrFS
7CDRGHxMhiVCoC0sHdcBwuSELFMGXOREeauULTS0n3NCUKGZKGyxRLSosarX
dlFMOK9cpHdhp30IkTtE5uyYLs2ICZrCkCmUz0B1LRN3OkcLl4VhFERDvR9E
zoPbA1Q3bJ7EMAkqy6HtanjRqLxA/vXJ0pCtME2DfTCKs6qw16cPyQu6AAB2
T6ANDugEydQs7VOpwk8Gic4ZOXRNJKrlEdU7dug8bBAmvNcfxP7DUKdy5zNL
zzXHylQ0VcG8hfjh/iw+P2m/uXxKtn9N3Xu86rHah0qARaxXfliayD+0tTe2
JU1V/xv1ncrbkM7TPsUjsFvGYtczZFXrNxmMVWqbCBP2KqyMfugtqR9yGSyb
NKGaMrCuM+1iAGntYcm4CN1wOW9NQjWQawn5onBybHBQklaI63lWyFniqs8o
WyoVZEfhLGKVhdm3pyrMKuhlBrkrnyG0SwFsbNLatPpMQQFLUhH2rTQL0ALZ
06JZDpaTWYUTV6kI5dn/OqgaWqho7bmYFD6Irx459xOs6UEpFtapKpFBzsTe
eA47qpBvJ0a0/E4vJ58JXsMjI0b19BRxm1qvabzx6aLC+Oy3OxvPXbEMIPCU
XL1CxBEWyODZugwjESQ13TgHOuSPjT2HkOymD1JF0tCarMUlROVMNkZj/yoe
iYZ7P0h+NV0EX4Os12junITSN/5/oHOPmv448pNbpF7jaaBEYuVT0NJ8i7ik
7VkU1/VNp8JrjyEbffqTbot6SZepMbtphis0WBoV43zaHv5r7t+PhUmwWv+G
G9BFNeiBeM+rcC+NDV+qp6jjKD/g/zQAnM7D39/AUZSrZ/zxepwtFNvdeQl5
W4vqTVeD9qEu+diI9EHAOyJOWHxnuQoDZvlONAEezRde/BNABFPd90sXKKhY
t9zrmYbSTUe+wu6n8Fcv/PrRRGU5raRYnxOs/cdj9DIhgxO7QwgZ6i92gBr1
Vmrc+1C2XSc/Ta/4iEzvg6+kjoyAYv9Acmbze7yC8CT9JL9qwYEjmSBIKuGw
0FPoX2cTA3SSgkVtC3Sfxmj87/QWLUCPpCdgzd1evFolQBmT8+hX3fP6LwbN
6sfBX5nlk6UoNbF8Z892hOPWsB6VSFElhznl0HyUMSmgbjYpeGCbD9sd3Ir1
JYFYHJC8ZuIJfue9A8nEwC5kE0YrQso60FlhBedrcQ8P6Ur+FdykbXxPPxDI
/vnRjKBTpTyEj9U5BhRhQLDJMxDkdHikInc5R2ybrnDhMJ9mVbLcVtY8e8lI
Ib14szwzNIWLQLihlYjl+IS2iZFGv39CQWDvKs/JnXk7FXpikda43D+8ViYa
UCEl4yWqWKtUkK+nO33A4ONjqDfOSvFeCrceRnELRf6h6iyuYUaYmlnWskBm
YbYydncR5FdD7tLc0e30wJ2LkpoJQCAdrocgF8vNly79fA/52MjBAqAcujsp
IbnlbPyTFVjBFWnVquSoQIEr+6nIss0tmZVORt892owZpaA4vlokAUks9+Cx
8uJjEFllB8C3rPwn00OB22hrEY9e9U0toAuFTw8k7hFZ6GCUAK115hOR1J18
mz8GLYP0bClTz2aOGruFJ+MbfXMCM/GrRptq8jXrqRX1oKXVf/ExpciHPp5x
Kh92MsmZ4KiHYA8zprIpqbo5VTX/jiGr4SVgvJfoL95ymqTMnmYXy4ph8JS9
ZxKbPSQiP1gVcMgHwm9Ffnu4aFI7Cp0ES//if6ziEoqn67/SktzsWmMbyV4D
IP8yyz/jL0rRb9bBiScRk64CxoeY17wb4lrfgCIs4D05f1gbsBYDlJkaPYor
tZZgrridIXofCVqOIpef/vke9Fx3Zh6XBSmud6fImV20YPr9zi4SUJKNCQPe
d/xPbMDsCO0NHV8AWv+s5DrPituwvmk1u21QQ+ktMDxsCGAHxJj73yN4SzLs
0DjbQDChoSNm3CvF+YoFnc5CkCcszW7yAu9qwpbHy3MKCDHsOKnUDDplNUs=

`pragma protect end_protected
