// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
lGS72Wii52iEIGQpPX9bL2+qTaUGd6Fhpf8s9cnptrfYPr0wC5j9BccR7H7usdxj69dJMWEfV2qN
r6A25b5w7ZTNdYSNKgLmsdfRBtvPHVUzkrfjw81Ces99bot9OxcHS2cnQuZVZ2/cFD1AJx8qAGvl
QqtAxPIwtO/hwW+LNMesKgynD1frrBXzzOKlIpRgwI9gSTpBHRu4RHYrWlONVFynv0Z/6MVpdWWR
RGtrZxrjDLGuug2pbDLwDqzWte53xdcmXx6vnxBD7lYtghrzOHqZYgAehpjLu9HjDma//oCVBE+u
XttjLqm2tc4MCmytBFZxDkuZNsi3/BUJFRmwCw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
kmSVQblLNWnV5zyixct8cZ1/cahpSBMrdYFw9km9z9lHRjPGlhYtx+HYGhDPXz8N1u73udWrZjg8
3vPm9L00UMI4gs01fz/T6lTZaes7D4NpZIZT/Vw3FcR7o68n+oJyVKShp4ib7XuXcpyu7dQN2nsd
ypGexvst4iBu8nhhSjIbUDtFpYbNBZCwm+z00zv8GjZUvGLlysEY2lK47kMIK8570mIbOtRpPcXV
0lmVuofVAQooOgny5I+JqJ/IWR4r00VOzhBxNJK0wb1WvX7q+gLrliyp2U0nJvlUBmwAH1gxJ5nV
1+t+PSXA2BETYXILvX7K3Dw0uMDqkQTgz47nddiVj1eGCfbw4vChHTiEOXzO63CNZ1N14+2glE1a
lNb+nXtK+cNzX1Rs+37R5a4TGcibRnWtJWRlM3nn33GM6L8r/3x71aEI3f89jiTA0k00dpZbs3Ek
AZpJCcgDDse5k8MnBwOJP+7rPN/ex4ArEgOYxKTd3JKq2ekZA+UEBTlbs7LSQAl4Bk3HkZsCdBu/
TWWVZ3UR8gbkLcQJZjJnT3XBizjm/Hlkt7lgxThDf4PewmnFWzWvAjV4fwJ+twb0PvRsaPJNh8E8
1QW5s9rJIkGf0J92WfKqr4fUG6siGoFpJOfsi40tEx9xT1669UpmexzaQGnhdthlFTlmg2rR5fKv
7VZhmaW4Iy60nLzs4KwXh8XznBaCHr5oUAE7HDn98c3Dw+80v65LJFQJCV/p3oe+Toz1pnKh2hf1
n3iKu7zzarwFbG+WrzZAXPQ0YvxSQ7JMFQSnoJF56qj97oDbKMwabEHa3XC8A0WWtpdLsSIcNqKW
x3WBZfmx8aZtieWx9Xiunxw6e5Ll4WbBgKRbqudowsF2q0dfZJ1IigmGPGvl23dQl//HypW4tpjj
MncHI1EOu68e9cVg8uBR9o2YdAziJP1gBRUgPTk896X0kW7PMweJh/fKzfSc83EM6zV7PTFymyYd
6p4Vto+J1o1LuocC79YHWEr8yYwFZKngrkOB67eNaMfgian+rCiSiQl33RV66oU4xwswcBTC+az5
fZHN6Up72RMw9/ZPDP8+f9HazH2NvKUVLFwNMXr1gPfiR/0LFwZUxx6kEbOilUWr//Q4ZrZ65a34
NSvoLA+NmXgVx9UsEYX9Ljmq6oH6pWnwpZB8eqnS0/LdUniVLS8QlmajzR271xNb2JMo9vnc6y8W
oNqe0OZlJXo5vYt355er0HftEHxVk/8BHz/KFh1cP75bePkWiwItpt+tiT7FRYji84YctgZxklzp
gugWN60RggFK/bdqU+cZtIiGUzpTMAXQsZ/JTgJGI8da02Gx27OITklyKE6KiInbiC8rlGEPrL6i
E3MtBRDWa534wib0gRBarx6F8mTNHa0LwEDiHeaOC2JZYRE5w6gTPJVXYPPc+RvkGpRyaIQ3I947
rXC+n7cmrDPEyTawQ4zDnX5QpPvInszy8gW8t4mIP+dYh5C/ok986T9cBXGU0TaUG0Zf3HwI50Ex
EsW1ajolMtTGhg+JX+GUl/DlTs/g/FIya4FXqenjUL1O1osaszBDSwp8uGmKAyNtlog5ZPbxOL3X
3RYexO0WpPX71WVPIHGdNV8rP9/UeqQTqMtWQvQdRBTimxyfq3f1Fs6jWTd0qmhOnCyxsxwn+go6
YhWKHm2mD4+9hWlPARcpGV02G3+BPN1s4ZxO98ECzfoEpfrgoI3TSwHdj1TKFoE2GD8ZUf41evvV
mmZdvTuZ8MzCOTlZPotUFrPMOpALHBA3fAZbmaXiDRIO43qkxPbm/QHsUR0r2KrnTc3LeVA06WrV
eU2l/VNCO25vpoCcBsM+WZvF12EKwEes6wX2r06uFmg9X/U4vYbC3eGES41E5lLHFwJ99tkR6hwE
NQ2O9SXW3fXJnOXhXdcvdGd7A8XDmbFwJGSxMPDx/z5G2RHHTni5l/NLzvU2zQrcGKtD/Z6ceXT+
yoMciHeF1EpH4aLnhRWkjDF9d3g7Nd5kaF57mQmEEXov3EkqNP+/bt8lzUQO9ZB31tKmr8M0m23Z
WxHnfAin7fcTSCe2Q653yORlrNc0cIh4n3ZuH1KU4mc3iK3FY98WnVVOUlP6uMtmymxdW0LNTBgc
fykmxMLl6xUyJI7eRJuZBS9GnASbs/IaE0h/9BRvjFiuWFVxwh1cASLBtSvq4KRiQqEUb9tcUsac
qnwFX0cukzTQszU/8LE3y/762lM3aDAAkx+GUuQGSteYTPhmWNo4Oza2iNuirLl3bAnWUq1FM13L
TiRvU8+h21no1KvjFw6EL4vF610RJV8yR5BXWZhPdAHp3SoNnNAv1obBT0a+kfjHONEXzkqNK29i
arw+vhNaVfmho7ENvMetcoBmOSgO0asmqrYD9TpuHxPNwRefVIwYZz6hyOyhjYRLZ3rqHWgkFyOe
09jldDVrynvyDAfISaT3ObhnYGylC+feD3MC/XGojmPAxrhxjbFX7R5FsracHhPyCmSYXMNnG7vh
51RHWRh0w6KfgVtncyqbKcj3A+vh31p9poE8mPfuLL6f9Qdg0tQN0ir2G+7lwqclDxIO4wM/mzgP
JY/Zbyp1wzhC0dg0r0i7cKa2aWvI92hE3P4dl1Rk6E/o8NdasUQYk2zsAjPxZUCfgSQNYqnZSddj
lpE5i7Gj/fX0B3kX1XTmY5bhbqNkyal6vbrUYUOxbqLv8X8WeGkO1eiy1WnT+/uN7xhzp/iJWAzL
+TuSeXXEieUlY8dLrtG9mG58cSmaREVMVjgQbIiRG9Ii93MF93GohoCMnFDbkYMXekOtM5mjXAOo
BalXAwIsEGm3H8/wcPdQMjgiRM9d/IWvod1cXE41+g/KcE4k4qQVpbGQTl82rO6CDUHkU36rpXM8
QTIW+umPbFfaxJLMuub9yKJyC6WXXsy12Kab6fr/afqiGPBJiK4DmKsN3OmyVd1vPlNnyW6hj47z
Ndblm96y8BZS5npfWLZTznz6Sk0XhZh6fOpK53dVKdPv2SkBYFJgGEFwaI2KeSCSjm2DBRTCFwvb
/ebfvmn2HpQFXHYyBiq8THzluJm5mHxsPY5VdNfIUfkxmdctBHGYxB5dqejoA4uLVEdLq6ETgdKW
3De6Kx2Mten1ujiHIMU0LBTqL4U55N2egmI9dJCmg5FpMfQHsILhnnYIRITF0tc3uIs06A2AndhP
ubEwUFUy8rCyMtroMwMMwRuAOkoF6V2bUpV+W9omIy/WnWH67/MeSRfJ34Mwxo1IZ+bvkzxDkNpF
qWiuBWMaiALdQCzA7hJ/lg9RVgGpvJPnCXiKXfYmnv9B/El/P5w2bBlVSwFXYK7XiOdxU0/3j/NW
BLao9/xqa0cZNB/gQJWqaNzTfe1muzvEYicRn3MjaVunnYecHJA+AOx/2ipx8VzFxz4UEDhhI6WU
b41NZ69RRbp2RyUNm7ptTKfd0cVxqQ+eA7Cr7pGIItAU4zNyl3L1OeI0vRWa2/87N4nbcAwm9rVS
yKI2AD3P4isyMa+1CEeldtPgXPD7Vb1jTi5Z7rtx2yfne5zC21wsv1o5sf7w5EerU7eDt5OgVfKe
XZmbpGMCCi4Fn6i00U6OQpPbP5B+neIWz3GLEtqi+PeQYl/FJzI1Da3wNHcwHodM3GI11E4rmiau
R4tZ+xAg8buuVOc76uqOZLOJleGGqMp1ClITq/Rd3Eda4y2nizKJYuRd3G1lWqP0PjY+nZh6dTK3
NF9AX9JwyKw7GeUnHm3FQBxUcvI6vSPTC1ZKz25Jh6H/XEXr91DyPI49zd2PqM6oT7cQUypiLx4R
PLhDPIGqZAM29N9cqtCxmwLwx4tAy80YUBGc6zwEButZlkoAR3Xt7ULGAyz5A+ng/sBn9rFxRSMd
WQBiEI5VuEuOf+UwXgRHkYF2Gk86oTiPMWyG9SJDfzihcT2+GyOaTATjF7eKp+VSWleXdd8D2Pu/
XUKnPHjnx8h5C1AkFjcnQnhNpxP3flwdiI+oMVqXUicfuGyvh7uCb+a9/qglEyqPNUeef6tslg1R
LouAikuTOcOhu4idU8s5LCqtBpawmBO2r0NLmcaAmegU2s/5HpxugxesJ8mrvTI4tVVofBcA8AO/
0zOBxNCnqp7CJNVz7uG8DD0ZA/0YWfY2DO/tpeaWly3gFqghPSvwGrheuHmOr5Ta14bv2qKO9Zfw
kL1GU0FrzicNPRSD7MQEp6rGsIbFiCSUAyn+gv/WXSl9N1EEuomMy+GqHjPgDuC9pQ2aGaNq5Yfq
db5gQdbQ14lMGTEvma9qStYdykcid9dHYxV4bOPeZHBZhRKYgJALZMvG0muPEovWrP2Uwm1xbefC
TjWF4M8MX/kjmODKGBBhvKOdycFY6xmEqoB+X5msHig8qm9KsjLK3hDfC2CF3k9Vge+kRzf067yS
cuKi6wl2iWGGqAuqfz/W77uVXndyAE6VwW45CpNLyqUrVBG5GCDKflPR+NGIZyohxRpBmJvI1gvv
R5x0AK1rQWYg3C3JgXXm8K8QxwoajiLOZZhbjqHUmf1t3Ig+xQHAdsiKVdcXrVV+1EP0uXeP11BZ
JyWDbi3uLDO6cN8OBp5/veujHEYRRQbFk3Ku6pSIFsNUhqAoNiOirT4kT291alog5SE6y8NA2BMO
tSDCOw4xHfK2Jejsme7q8Ek0lNoVdnwKE8fn4EK+TsjmW/1GpH26xSUsUm0CyZe+jr75k4fKy0td
F2Fhual36B2rLeY3mwytMLKPFbs3FnP0rfk6vNeBQpIb3vLurHM2blugJk/WEpyg7dh1jQ99VZe6
APKFuOWBfKJ7yaUj2kSZIHu3WhLmegbM0zMqjRVG3lcAfWJrlmsaxA9o8uPj+3d5dsu/oXJN3e8n
maeoef22DI2lLovCydoFLnHhKF0s6U/UJD0Df6RTeSEasg1USVkLMKeIooNQJP9km9y9ScmuYFVa
4aBBkRHCB6QkeX9Fuey/d5//sCD4C1X5EaUlSrZ1JPuj0kmRL9v5qWjPGONuJLkyCDzQeHLTGgwy
dmqaBmwO0/y8pd3jv1vETz9S1U77KGdcy6UPZMQXXYGC2hJLd6K8O1yBIgbqZU3IDOQ0aq+m6u6b
hpV9s/5quYH0vC7dzA7pTWpIzXuebh+ykqJUnj82QmjskmPN9g28w5ePYA8/pJj7JOz8tDdffhox
vx4SI6GU91llcv6qSBRxUMtKWv9rszQN3uFCEQhfMYU9/WUHzbVIZNpldrv4KVkUWYyGpfOejiG4
52cWJiT7DLZwDMuM2LOmAqle0VsU3XxBgYsqX9S+ufjUZPaZc+12avnfGFHryknqBkyTqtg9C7k/
dg2qK+Mc+WfLOZNXEoH9xj/qgPVgPdfHBfEB0vw8VXQetx9KaD+aMaSgT58crR5HEA8zinlJuB3H
6uKjF640UIkbFvl0g6LlI8ptrs7sxn/VV1/sm/AIUooRG6k3OBgmUzwq4s1lgBeumJwUkjSM2/kk
5HloGjkuzwYYZFiRkz0f+I/z9drY/IoF0xszQmz1sUKSf3ZUFW42eAVYPgX/akwWNlw4o19daIvv
qv1qWacgXY1Gzk9g+ibI/+V5d23Kvnnay9dLGinFh3eD+NrbVnKtkNT/vPTN26sGjnwSDIT+YH76
t1VFT6cdAhUf/9fFlKyBu6oi3Y6Nfd+WPexkIj4k5VCDO7b9TwYDbSyUys39S6PqvVjcx2jJzb06
zWdl1xoyBflAkqeEJjNGUVI7Xd/sDXjDHoSapH60V73FE0UGKeBEw9yOu23uC8WQbdMIsqWTmgqO
hH6T1rAhejHK2F7rJkKuPNV/ooduyGW67JbQRrkNaOrCS5HMEnJ7UCYGvvZ/N0wX01lygAp+EwJv
GeK4WOKhST99FvTQ0ObpOo1j7/ZIwE17MpoLkZ22ihm3XCiHEuxMm/b43cl7F1rQfMBV0HPbjSWf
CbuN5HCsfugWf575OOC3OAIFIRJCTTjZCeTeINJIAsPMcz3N71ZuovFp5TPkMFaUaQzMNPgTCc+1
h9MzJNpASY+nkpSz8p3ED9ouWvDwPx9wFYRSAoDXw5ysrt/+0VyH/rU9TeG+xxE81WmedAKEGB24
0/w6LgbuFYS402T6fyJves55m03o0EZ8HipDYJl7/6vMIeqVWRLNNEYTHYjjisG+sPa13PNIiIkz
zEHtJ++wmZ2XOmmGSlUtoM4P5MWZ8lg7Y9fN05b//JiKu3ERGTXQzF9BnMc2HU/4UK39BpvWT2de
/OilYA+hAIGxu/YNnrKllwF6geL8q2f2CB+uw2hPIm+pIjPNYDcplR5N1psjV+QJzhsMPp1uGXuh
7E7/d1hzhWDBuGzkBI/F6sqCDosfsUCr/pYjx3/BeEMdPMbEocvlIUyVbxKy7jlgNc2oDI7NyT7l
SeMGEmQ/S8OmNG9rvFtZNp5gXuiPWb7K7eLfcIGq6FAvAeI6t5BXQLjDDWEUGGpSckm4NW1OtE2m
OU8J3zLPGFyP5iLKior0L+Jv0i2QRpxwqXZZPqrgCmiV9ktYkwxAeZzt0CmGh4A24GnAFA6/x4rb
8kHWUaUhsyzK6fcP00ayKnAQUv5w7U0InjnWbjqmj+o4bzJT4WK3+Kq7k5RP0xpeH3VQ7Wkvf17P
i4FO1MP2gYazku0Eqkn2V6hINIqvkRbZ83e7i6BjJnlOf6LjoH14q4fhfnHbn0qBqxZfwBMCi5v+
ippF1+ddOhf9OGRo67vGgri9/izNdHdLDtUOEMIXI2NQn/RyxQQDIIp7G52eh2ZrWgnXD5DOsBBQ
V3VIa5GsUY8/Bgq7yXVlJoBvIoKtDDtZfHUT9M/lj+YmtOJWhsxyuv5khRW6rWNv7MWsDdGmh4G6
szFi21+Uon8l8hnD6a2atzUxqxzCxUGuJHddLR73NLUQixhZyCIb673Ik0XJcPoRi/rIsJhpm+Ab
jDLTalO3IQeDmaUAKWM28cp7n0nTwnlXUIDiB+Q+mW5n4tKHJnd0a7r8TvOYlrIH83IYHwi2DoMR
88GJaEu8bstM/7jBw9+mRfKTTGG5ATAOhOE9Q6sKtIs/s0otvlRZAwgF3tq1zrBrXy9R4aldptBH
AioTqIs8qlf8Kbt+fIwHJqbOXx1DNRDPYE2K0KHM9ACyBFuPGR9BsULFNCI4gWts4e1UKztj+J5C
hb2mXmIXv9ayk/K/KjmT19vJN9Sji+ysud0cOmwQEZyMp2KtS/QWIZABsf3m+knv5tzPsjqFq1AU
GC+lLZi8LLU4XNP07YOY8B8pWGDrgqdCSFWEfhunEDnGMRZhIx9BE91cNu3qVcJIdwGfhubUljRI
fhAU0ykM2ec6udvzBInrvJfp2zE8Eu3/QJhQBlXdaMzC4dI2UXSl1J8BYJZAnc8Fh8k1FWNjWKGI
3t89TlvBrm1ZeoxXiW6NFtx3Wa3RI+ZoVaiIqgi3ECkkiEgSExaIsrt0nyzLxViyS19QwkTOX9lv
FQuiE6awA+JfUn3L0+f5zEcXTVal+A2OUcCqaOQ/BRxkm5D5JQuVxjuRoqcPZQuzDlQgvLdyIjgr
i3XebM7Oo+c38+R8g1H9SD7SzgvPaY4sQmvxLxpxwWAbtS4Un3WefgYAoRu6fJy8/x7JOhS17Y8R
xPu2IOKON0hqK1M4XEk3ZkJqkhSrPeSlFYSdqoolfXLrvQjpP1O+EM/0p6R/d91eFY6jhciPBbI4
zOvxQgdaMqcvamN8j21D2t2ImUPQJY7FA5UedvkojxYKof0JhRfp+eP+2DbgPFINVAGAPsQJv1BJ
DSpFu3hnXPj92uejYKMuin9UcnS6tVyIeWGTM2if49otSpp+XiwdD3iUA8GiffL/ZaLDqn1Gly2/
MT05iJwW1AiNDy/4pRzdt+aqCDGVm7iaeNLvIEvo10FnvmfUorGQHaCwucu2pMlEfLrNeanSBTte
JtBpZ/LUhm7R4DFYzZhJKRFPLXnesAkEFgukxOwCIYJ3YEe81mp2vHzoYNoJLAii4KbiBSKi18Kb
myGLZWgOEbW6ADbrZqnf3fi2nK5zTHdqJts4hw7nVxXUH3Jcu8eHYWcx84kmNuAzToCb5agt3p3E
ysB9OifGLlZLWH8XNDyL5Og9gTLN73mabTs6sfdSZ1CFA2ZPTmeGRMoDcTv16Nc4SoDP70wzV6zd
MWbZCLj8n1iHqrqDHKCqarz+M6sLh9jAvISj5uKI8m81t6pky6PWQZKSTSguU+WVP76LjyV6mCjU
DZRMbEePk1GW44TWfXuieq1F/SqBCGJPNPkmfGjxwhRGV2j1xDG0nvpb/Roz6Jtt3EW0yHWNJOiD
+m2RgjQthcDxrOR1/4vE9oIz3LAQwvWSenIUHJN2lOrNmebf3VvsI+VCpsn9nQGa9onZgCm7bloC
s+zipLgCJxTHBSYMOQG09KcQL+ofrt0elNo1o8f8zwuvuji8VksCvTgsWoX6Kw6+FsZtsaBHcQ8k
b7iajM4RuNfhGHLUpG5woePikK45b1mlfXJYeMc3+LXDPbPp7Lgp2XsDLYP2Jg+/4YTcW2Eumb13
rHGOM/qOzgBRdzq6sfDLI3ZHIqmFpkExIiMpwh3TUEegQmd0adTyeSMILhpwhNnlaFzQEyQGQGFP
oA3FVhPFMfEIKAGxxL9RYQz5Bcxq5Hf+LzKfrL3fayLepc4OaRK96gYo2MRcIjxQmSEAXL7psAWL
erLlxj1axpTg3kH/bk0rKTP1GRtSpLZz20wXLnz7sLUhjxkqPh1QzwywOMUXGa5w98B5l8uikkM/
gkyxLMDdghwRsoOyilLdUc54RVKO02k2ttCywocDFTmiVcQqTasGJuJyn3XtZC0ogMGIXj5ng/dJ
HnOClunjsizWyQtJYQE+VtsqIx1YjptnT5r/25DTgM66y3UGabF8ZMBYjIoVwzVoM+yGDE/ovFvp
1IVG9xeVbHdQznw5GZkoc3m2sqOIA0WclkIVoy3bDg3lejhDft2AcyW6PZrRfom7xLMe5Fr2IGdY
stu9dOVvqRqrXq1NrqswmbYTkLRhrAIDVqlKLewdNj4DSFVoMCCQr2ev/U8GDzHm8CkS+Fe9yykO
BP0/iIg3u+nqhM0pQyI/WEm8n8c1bEfQCIodZueV0m/BV8e0OH8nKL3fuvGtEADcfTy4p7/3laqS
KIgMLCeHmqCgyVybsO/gtrQxlc2dE3lYBRef4hcnv369pXhR1L9pGmiE/OuEVUwutIEIOSIth5xA
dwLktGcVy/I19oUM7HVniAO/OLPkFnf4ygHNyqI5ALHFn5zoh0keeVM2llN2d6x176o5HDBKJVrr
5WvWbP0p8kgSUQIi//E5gAIX2t4Tec5B3NNWCcKB/g6wZIYO+tv9VdfGZ75iTiCPom8FurPmIATJ
WnWxR7H+EV4yb6zwIoDyqPe6jdbrKqgJUnGhvJBnTD1KPwk0Fsy7kJ3nAm8RnM3qoJlAXf/BniHx
j38IQBhQsBGHe76SGxdS3jnFZM9Z2cag55qnUYaL7+f5S9kVGaR9uABdZgJCZp0fuCz1402gcGU6
wqUl8iS4e/uFu3HPyPy9s1/TloTIunRMLijfF54BDJlbsxV8LcKRCeeBF0JQuRcE4c6Lck8WkErr
hyxG0DHTeZDlbgPrBCX2bWQ/MuOpt6oHFCacrJHi3LO5H+uycH9UssSoQRNs+0fRhslPX/8TJ3vE
EEAeAMgGCZ/aYsgFUG8enX1hvmc7D2I6gCatu65oZGFFMqLY+QjnMqxyGjD7GGuHsJqO3vNYnfDj
SWXIXNp/vF5NwSlcWBdEYiAkja1tx5ATfOE+BbQ3A+VOgQhbAF12Eu/74/NJKa3rCkqd5f2g5/k2
SEYPn9HIO91an8985C2oa8MJu4VPPxPu/BOMTrIUzhxfNTv+dM/30mwbwFyKYyzuynH+yEsRJG2z
9SQhypERZTXEH2gCid+PZ+1z6845uoxQVFMBTPralU6dkKotdHnVrWmxp2FELCQ+2yQx08P6dy86
5h5iNQR71dshsiPxeGHDUsfS0pQbETiNepvGYbriT0tETpkMECK4QVXiTZs69PdvXGnSWrT/P8D1
n0S+VNIRq9+5pIWqeMME+57RJ/viOWkubVDF8T4mCrRUb2B3AZomnOuNHMVcJjeFnHLLxB5onkp5
sy8Q6DOofy7vCFMGl5QVUmNlvUU18QEQN9eYHZrUq+arLT/UEr1JAEBMvGmD2ho0YYjPukiEIxHI
krYJmPwizt7Q4Ny/J2a8ttC2W75vR+DgNPdbBPlUF+YGJkhMAFsYoBManEqIPa/suZO5yqec1Vhs
7pwVAMCIeesdQmGiXRYPM7ZYqB3wOSdd7QAOMHCze5+N/T9CSJCF+/1ppmk3iz0aMHMizCGuJfQ/
M8KOxKslc/YnHDa3RagJ9lPeVeEqfw01KcnvSjtAYceAoQNckRWuhlrir4ij7WqHgscYKuHYJyLg
03Jp/WS+sx9FcLxtyVuJfJLWC1CdbO5pll3z4/LGYm6RHllo6ZxqEhsJIBD4j3CwdgBLr8tlFrG/
d5XNxxGi4MJPQ3thjt1RgPA99N9edGpUQ5oj/BuUQKt+PbmIzQ35SDqUqvTlrPJK9hdwLXA2ayIM
CT+qU3uFhNRUpIi1xDe9N5FG0df60Se8jl1VDvUEYrlqpaBiUiIUdO4pP7hcdF+XuKLMKK1Pk2XL
PhYNm20hGAI7FfhLlJeyWDfKeqyHvqopp37Cn+Yqi5LxdtTPMHbTwlpiaHbr5tYwnKRQ7eNu95Zx
gjG3TMFepolAPrHtiZ+sqwxz8i5SsjP3hTdgMkhgNhRXwPFm8zJMg8X/H0sh4KVUTc/dZkNToUCU
OYiEwNM3Rc/Ew1t//H+CQYD/dY6alY4fqgk8m+ZPMI2XXnvOYcz+4wvwO9fDPL1Rf5Nqbo4GU6mt
6knuVFI54iNe8lMdHWZA6QKS1Z1bDY3zz4C8ZLpmQvJFrENvjxyIb95lrbWqRxx7nPdTcDi28QzV
OxSwpyRveBBucN3GXhb9nWR4fDT4o4ooMkCUy9dkeE+LLqkS3Rdd6MEUIGi1jW0jlB2aYrdOBb/P
qc38gIW8vRXzZ4v8Pas1nd6urkD7TYDKtZrsFdSs3RYlqvt99WQYQ7WHuBASk+Vt+EYxFN0lceN7
bQ0BfzcFDh/EMfclUOm/V9S3axNM7ea6UZCiE5+k/FIWp+eHTGVOjAvQWownuWWo3k6bkhmJJgQB
oYnmuXCAGIAjn2TkfEPbuyUBvA4tn+kNkcUbglVe6/G2JMfv7T/yHllBAfvvpMvjrS+X5deHzHNN
tLIM9FHXPGmJI+2C5ukSUm7QXKE7Pejq8mp0WwVElbgIe7WyT5XUS9/9anM7REE70leHMcwbPuHi
O0kS
`pragma protect end_protected
