// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rJT6D2ZLM+wmcVCTDoVZ+sXr2cP+/JFSExbh5MjTTcRBKikqb7E9qUO5UYsxAPI2X8D6D+7AtyJo
MIQ//kBaRWaRkvZnRTEE03hInBsrgcIVyIjTcShNkrMLvUFnxxpeRjagh+/F9r0uPVTkRbJGPBuV
s7rgIbQlIVqZs0TInp6GYFBxCFM9x6BnqhJ0LhMNSq+SLbJsJ90z0FmDWr8lZCLgF4f00TiK2ven
tjdYQes1aiTfO5Ui1cCjNdQYuDTT4MQjNRR6d3uv4oJvtnC2SfW7MI9ZFBmwYuvRMbpIr+V/uMp5
V1kWhmQHHYZ7UFaaAVw2dHxJQsDGotZqnHAxDQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
7+rc1ORp111R5sjMQSFhQac3W4VQ30dumAziy1S/dcrYfM34P7vVKfYjaovF+ggaeJhMoBF62Y0j
UqZfAV8QwB8eO/3ZFjCtFmMW/MwOP9yzCO/Z3gs8pZQWciBH7sWcV3wxEObTx9THomjzPhaFHb54
T3lkQuE3hQBlOt5BQDWBLmGJfrKB8QuPfRFTHNrkNYgW5JKhf22a46vITWgT6tOdy49S0X9Skt6d
MGIpOAkm0FKRI3w5VH82I11e8v4K4+x5zcAS2IxKRqgBiaywavERBkWu9AenFjvncXD/gt+i/gaj
Nlgm+Zz5/98EMhVMvZ5M7z4CNUB5yTC9l9VWWZwD2iS38HIQHRirLx6iSqMGcswPKLpakW2/Z5bD
8EkZm2okVPibOvl09Ke2yOT2+4B2nVrdRKYKTPM5kJfujh7xReB68D6XJY/B+IpEl540rTT8Wljd
4rguYMg0wQ4MGpWuDBZcgSDFsXKnF4l8D+Gz2xyB1fI6fsbmU2yagSd86A470rHitGakjcPqQIkS
dB2Z2msNUhl2CNpbNZwAFdaQWhd4m9qd9OPAc3GTVMFvb1mnfQTiL0SDALm/qlto7/GK7AJMyet3
BX7uoPAfs1Y9rGdbKap25tNUQk3bLDsvAmDKvY+UD9jp9vSRS2IcRn566mHSvyr6JCfBNiScOE3S
bZdO5hXgs1kmzaN68enn12a73Zprlq6NTdwgDumbAPp8iBf4Pgy5fM58fO3vlwKzfK0/nldzTN0h
WZXCdsZ4RGL4zU0KADibR6H/aBaafox1ydibFoO58L7xQVoOtKz6Zt0wYWdbSOaoFTWVwYkZAIm8
/r3Z92ORC517PY5dATsQYLcmVQcagzHHEe2qaJUL1DsN/yaeIVS7YbEPXyltMzwQ3xRlmm8nq271
hKcK2ie3j/ems+e7E/FFCuz8DApRhQVDRp2qZ8MLEwJpeOuyl7a/h7Fw1y4d/XPqbCy05EYOeyp1
fEI2Plbr9ZUMJtR0XgYi2QdbDHZJl80h1k0nkJ+l9LC58QdIHfhrrptY94FPQT9U/szEQRwydF3i
hRhXrtx6lDMM7DVanWOrSxMHfx/hxAM7bYk1p+ErcA21xuT1ehRVjkLDXIsRcY/LuLpw5m4gX6Vp
omNuy+5yj/pptLg7E4w8MctqYkQ3A0cCtPdyjxsGOXTPjVRrFBvWswQuQeLUm08a1QjCfVSkVHxC
OBXJbejPAYdkF70GNOua0D8M9c8EbHoKxMNQW3BVpHM1ORc+ZQmt+CRZwOJgXOcCLyDLCS3OE5fr
T82/bqcH0aPp2hkT/yxPmRhSeG3PBiq/B+nIFIGP+HDn8frZ/Twy0Op8cyvjcc46K5QjaUdZAK9t
AxCiMivLGVorrvGEd3xwCQ0GmElrIy0KcPUSKoEU28/fQU7h5KjeF8d8XFkw+rzttCKfiyzSIm1W
PMB3c9YxHpRSL1/2vingwEJocG6CLJ+dOH1Qn+YDj2jw3KQEVbKlCn18Nl93QV7M8fSPZABuQ9OP
hiVvE2uOJ8HpOvqjUmRIJhlitRfHKDf8wIYufj2hL1s0z5Ijvgy4g5SBbSr0k5iGIsxCsmvu7FWp
4V0tJekGnhrww+QCOXMaB0qXimXtJivONTWIybt7gpLFRxJ05I/xd+SZQEq4AzVBvQ2d1rVOtkT/
t4VYJhZSrzoQQr4wXls1uwEqeiQT9a9afgVmWu2O4ex0RiB2BRohwZNOdY9Gp8Vvb8u4eU+h/1dP
syw1UNlfa86oVSri/Wvw2nGytzAmVA5w+9ED4Gp6kPZZSSRy1zjEOeMEdqbhuZRb1IblktDsVBDp
ER76XBtxWF5s28s79U9nfSj6FKUa73ETxOjwkasD+jCMlneCENMyCVRaBofsEXQ4UiPB+zCUwxD1
vUECqk8GhHJ448+ZzDTLw6yPAyS59uaKibuuA1V1nnT++7OfjkzYepsVTRPbfN5wO/OWgGZvh366
042QGGP9tGDDmixbeJN7/kPncOwaIneAksJZ+NudbRp/y1tsBWiv9ZrSgC9psOmXy428PPK2tJFG
XB7BJakbSgvmlc+lsCyp9BsdOOI5TXBPwMAqpU9JBvZvwYJVqTEceuulMY02nFKOZbYyQsvgLHOb
bgZgJyD9f7UQZa43Aaprb2wQQ4YMRuMnlQPzj1HD5TbM27YVSEOUDm9/rq6w6l+ohNno6l+dAmDt
kCrxb5swVyLcYZhbw1bWxC9kKA/IEKI761OTIf/0nXTawkfHPMaK0hr34AqyFQ2kMFZH/aNeZP9Y
q2dy66edpP8QTLPia8dIzV+pqtxyKM6gkq0vJ6+rUjsNMAbVYl7SzSxoJfJHTE+Av13TUUqubSuq
oSAhoH5NnpGTwh0rd6weUQAtu17NzsS5ofU6un4m6cotQo0pepoGxsFzAnO8JGZhXyhLIVyG6IYg
zy9icKbVyxKxzOnqJdxwZpU6z4u/2X00XphbvtWtRKgHUTNEdftPnysN+YOxMUNwfj+U2DIBrcWV
3x1VXmPNUq8LT9rgFhBlmF/jmLE7+AbA8Y5PefZyXtWUoJf7tZk5bKyuDA6Vx8qVCT9HLjmq9FoZ
+mpr5TLE8pHuQiB6RgV9TbIM4opIFA3h7qJqG+CUhqmuxBvaiIzFLwBbVNcxRzsI45NVKMOOC4lS
MpCxs7plrFnLgbgfh4+rtomeVWHeiFs1x/qnl6zj5mB6Ph77EkE1/IekE+f4eOMT1yaqaf+va2an
1s05aeXacAM62mhjL17MyC80N3xnSUp/vnXn6scM6baHmsslH5z19bUEfEe2OJkrIHg6WnNP7+o2
9hmIjhION8aCWcvOVRbkJpVi8bkVzIQ1qYSbFq5ns+82N4Ht8n6sNn3LFioLi6oHZNZ7/f0NrqZD
A75Crvws3BdCvb+X0W615jLTxbEGolesXTufbf1WWLBPmizI6TOcoj5aqXyOEpmq+xn9MZvnFn9+
UCr0gaUnN6smAryCkwjgTk+5yCQyND2MF7rnwITdXlV8FxqA8L6p0ZCymfjDChWOg3J/TzrsMKO/
CEHNY0WcLTnToXDPz+WweYTTz4/W8cnVhitOK2JC3kJqiw6/rvmJHKEuf26yw4RW4aTMeGX1+QyF
sdS+VH+77keNz4AGoyyWXPu/mZf7l7Hi6zjbfSL6PFLBMHUwJ+IXlEHwOBau0N9a4aOOJDmYaYb/
oTHUGnZiRebWHv47SQUCCHA6f6DuKFB0Df9dWb9/G5GI2jdaZreQ8kodXsyRWWL90Ot1xtO2Z9bS
J7U5LR3QKFtIwUhjYnwUsnFxFGCGguqHdxzeNe9cKQygSRzlUOceepcKpkaue3rQ8ONag0j64oOl
QLFs8z3zMiHnoeixYbDqhvb7SgClkaz0uzzAr9FGOkB4kV6RN4XsTrzW00Z0Ykys2nVu94MZKySi
tIXE6JbXQ0yxMZWdBSXBc2LT4ViZc6PLwWY5BeXBDVFO9Vv1PdMDrxmpH2BrRsUbtqlev/DK8QGH
Fbypj1XyxTiEVrqdPo9iPDpRt9SmQySmjFxQRhHoYpQov58nueqK5eV8FiO1mM4MlSQsmVPiLbzP
6iWqdBSKpcwWujTo6WsyuKJj3sah9/ILUPoOYHN3wwakDT3hggzE9FSLW2oEfawmyVm289rAxDv5
C9WvrneU1LnaFOqhN/tSaI/+lj5Jr8ZNd6TgAcBL0T0O+EkKqdNebqxEFcYIFkQSjtBda5szMLQs
lWMDcI++CtkUo6DgxUryj98Dn2XCeIpTUF0XHGQ/9lYadzbWO8EAkPyOUtHnQlYqbUCjJDAlguk9
tV9zPZHjStmPt17kPfeYDYoZFsZ5DrjGrqBITFADf/X+VIeyDI/neJRiF+u2h0jwFTSbRSEP06YH
k/vb9oQVguXOocK1bTScPtRqu6nL8Axj9xy3pnwhlEHsWEh+SYohwfC0zsjrntZo/bIRtYAlrTgE
+uaH1xYHR3LWn2JH12faN/8assy8pLtv1i1AjVhHCQYSElZFWaszVrwlkF4i9KeqguAhyufuZsHl
4s1b6/rIVp6RYvcCQbMat7YA6kCEHkD9iLmyyvPjCVew+zwFyijcO4BK7nH2dy2rCbnsVl4Ts1nl
zKx325mM+8PzGvdB4aPVmLeXctIB5Yt1SN1z5kPJfkH+06tRbINBJYycULBJJf4QFqp2whbaPs+M
744z7bsTL+wsxp2HymoFv9KiwdxvabmIpyramreaXGZUnNrMKC3qxHT/XcNSt1062TsjxRQ6Axx8
47JWNUUW/yCJ9kQ8gRwDvX6XqjeUIm8i3nIEYnU8BThbIyYl6KnWEwi/vK2GPXvz+Ogk0bc/MGwM
dIA8GC7ky+gzzR0Qsnv0frIOsoMC0EYFXVmhJo9Wp7Po0cLx3JTl3E7wT/9mAahiRtCrjAvcwVQ9
zOn0TwaHADFgRowopQJe10E05g6r5uWg3ijR7qFWgwtfjxwOm7ht9oZKT9NRQrx/IcRE4QY+R1N/
NzbgKL8rFilqwekEfzcpIFFwkmeUXiVSYbGWz+bqyBTvtBMJVRhSjPN4u+w27Ze6UtHMq6PgGrwt
UNWLucVMfBAGbL6ywEzPnYOY/BHeRNiSQk1tdHenXxGqhZOVg30xwlvvQ8SakOmLadzpT/k4bO2p
Z8ZlRmIr+dOyV/Q1GqQPt8MU1W6vXM5qhL/z0cr4WlYG/+ZgzjXYo1ThK7AIwTQJjfsXld5AwN2Y
c/qa5zwOupDSz/QTQ5BFl3uYVlGZkV5GUqSWE4Sc761zkOsqhSUIxEojC0YwMOhO1AipLw/R6fSK
A6XDZekIfzEivUOgWugQDpW7/lzrdR2WFdOHDseKQnm9eSWqbScUuPcEW3lCyZaGGuHYOy68AAwl
oKMpWG90eC3T9omqrUS0e5uDzrK3tFGrej/4bAmDNFt3gwsdItuWcb0z3iiasa/arRxVd4wz3iSM
wqWNVpK+T/XgLZoDfP4n0+oAWD3hSr5K3mdfFnWwH/S+R2RnwTOE5X16gb6mwMB9662sf1mzV29B
TP+1gX327LiOEfyjA2fyQC2ArZA+XNTH9iecLX16gl2RRqjysZT7elirYL5PuLUS2y0RPZhFCjnu
KzGzFJnz50rHkr2j+0thEW2DNgPJacr2yz3mOEgX1Va6iEelMIqZ7NsBX0kBrYfHuwYz83ivbYS+
KDofGL6rcyedl0ei3n7olGdVh3vd1WkFQedlogg4z7FHTrp5Ud3YdJhXaMmRvStn4LkvPFw9TARH
jB254rczQ+bURdAdq84otNY9nzDhHU4bnFiliW6WLqUontnSYpJFq7z0AOs+KuDlZ/fIIxfKD3K4
XzVsFyBbEqwaX6GDfUKwWgK4pA6ukPqbFB9YctPuMUKZ3NFNY5kFQV5usdrSbL7k0hoAI5TbGJuE
pZFhKUHpwtQekRBgFvbJFhnQq3e96l2GUf42teg1V0xYnqMaEGvxoESxzE6f4FeKVbOmdSyJWOLW
ok68/HodOMGidd0CPOSKeG7P58+pvUykUdkp3rDPAwpVhrR54LRy5wmlooZDbXYlI3T19pcO1fo9
79cxB+jx6pL6RORGLNt4cB4lpNqc+oan+h9y6cThvmSimcEXFsm2+seMO5DlyGwc3fo6+OOXDtq6
1ZOBB5IQreX7OKuTzYOIOvRZDgA1oadlSL5D3RneRXcHGLzyxes+Hkum76yE52c+ZFfSRYGc12qZ
+CoEjH/Y3jLmptLKgDEwxNXdoBKQE6X6CTo5pLkADUgux+hlEhFtU6TyRwwV3cfJtyCZhsdu0Grl
kVfbsEVV/nArLpHWqag/vtICQmvYbTj6AXA2NFmuaKzZUnuzcEh59zG/KbcREe5mYed53Qo8T+KG
kuuYPP6z9HcXEHAHqQG0xhxWj4kDkrPrk3HQIq0u/aYklgQwgCBOl33M3K1g849475O9EhPLTYfB
PFlMjt1WEF4dIPwRoTJn1NcmeWNoArp/fGE5xqAInaU8xMzSeWvENHz86df8dIJ8zeLjEOKGrjp5
wredHpHIWAwfRVYT7Izx84AQca/5tHb7hVhZsZfXFAzfKy3BJJgpmdqe86dmGNCn6U16sjdrHhHL
WEQoYTWUFIgTW/wLdjmSr4k5NLG6gMBk+u7S5Bw46w38T9jlUItHzAhnLDCFksRuhFJIJh/k8ZoV
lZtZ/0psOXzUjDO9TzElyJESThvN+3b7L4BwWSpw2el14u/q+nIpPlQBTkW0ybLOpQe1q0XrcRx8
V8iZ6HVkr07m/JFsz8yC5BIjKTkKI4BC+kNHi2Kndsa9pkYLAoqfZzltgoZ9kYGNZucfg6iOlivM
HwpoHE6ojoikj7X3T19YCDwf/sEdBSqN+XkOF+pYaLVnlkuaPQr1AiDwVJSMVcAct+2sgxtK0ZhJ
QjN72c2OrTIRMyGwg5xARSZ4AAm7z/eYTNMWycosZ/P3c/OjVaYC+TN7wk2oc7k73ASJ1tF2xR7e
UC01BDnXX5dbY7RoTiJuQDFqCIstdfBDnY/57KJwiQ/KK2WYdpaSSXq/2fiB9QGRiq38+7K/3uEM
8yIGIC+ixC8tAo0mD504GZEuAMB/sbFwBAQIeeqpRMgIu210d5AebeYW5G3f2pxbjRxIGT/pmYOD
/0ut4msln2xKviXjpHpV7wJKkIFnGrigjdQ0wa8YMMWK5ApM+rlLXPFquay5VEMFbdp+ty1r6vkJ
hMtYdb11YtY/SNCydZo0RFVAsd/+zRfkhdXTdf9eUCvZWjKzkPbRFGbbo9Q1yb5q3QFAM29YbsKv
WOzHaap7XX7Rl+QNdl0S0TkFusTs9mDTfloju0sxT673WSRdLHhpAEOQPCGdDwTd8EoynEb5ihXD
us9u3DdGF8+6xorDuEeuSorwBsZ94gEqSBPPovKOI+9nlwnU/MPJIg8qFCge20e8zqu9+56hiRrK
k/QTZ7UQ1pHOEdqZaF1+kGdaj4sqfFXwwzHjJM6iD0GuhTYWu6R8RBWpvDjx10cuKp7F8QWztoUU
IP1XDbDoWXod0HBUKu/LTo/w5IbzwoPDftcmLlyOEcz17i6PgXHH/gb+gm4oecQ0zMyOVO2dU84m
2FY6ikyxthJA+sMFuchxFlkoSY8KR7u1Eoh6MK66Stv1t4/cKQgCLhaT+WlddR1esMmTsxK2ZqYW
o4BtgUNo8vSprUaxmWCOI9vZquUKCS/e0E4smzRNE/eHQYVyeXaSyCqewyQxu3AHO8U5E3UpD+Ou
DeffSmCYibX54ohallNOcs6+msZjfdJQoijjlfTe3UcgKVvfakO05xSXlqL6EkSsoGFee7zrI77P
QCcblgtQhdvC4jlgMI5zhRCf/+Dsa+OkviKkE/WQjCuZ8tU5C6tAMrJ8Fmp4hcgYhUxOdQauEyzu
Qi7Y8fNqrl6RefZdl9cxCPjqQUzHTKSa9stjZd7ZiT/z5O4hIf/vvLOIJIEr4jLdOAYSd2R2w3Ku
Ihh4TuEzCrmndGIhjRwj6bpa4X+i71x76YwLvjrSi4tYKtdOAVpFoxqoDsSYLr1oJ8vE4jHPRhvR
HEXXMkEAsbgWYO7Kx5ZsZo9M2HhyZLS4ti9KlW8xPVaYnJ1YS/4tmYbJirWV9AgKfxpypY2EDXVu
++Fi71m+NZrYe11H8RCx3cwQ3sT146HbwxIPdZs5rK7U/xLSQf2zDFMYU6gPhChfHPzlFANwaWLT
9ocdsNMPiZXffXBlC+TbIxATVONuEVgrUNUlkAIqnWNJSQ0UQ4xMx2OuvOMGVrT/Et3alrD3YWIM
O8gUQOduobagSn0IDYbRq+pI+cBHEVITm5X8P3aKdHtvI2nIKnJDYlmmM7gZMUSnQbhJBaiDES1b
xPOZw4L6yUnwZEqk5o1ZEfAW3QhTbg4zPVBibTjQ8wrPXQUg2/QVxPsakhUIh34hUQWC3QwSKubR
THOYDHvrTfFA/XtmCY66mDXf/4A41WggA42D6Lc4PGQCghwNR2ddUSjMOCk1MuGTKNf3q8N2pN+O
z+5KQ6/5t5fy2irvffOGvvjjTR/SPRmflmq6xglsIMq8hqndwSMtbtg8wTL4JX9cLsMrYZ/xkgee
kCmAr/rdgsvB2OrFnZaZYc9zrJZIFFjaOv2/HUMzIuRHqZyr0D2iSOTSbmJH9yLuVh46jO5GYCzN
uRGD8Re9Wragbt/F31i/J3JZy8wMoliCGI7f+gOz+Utwkqbfcyk/shToRvNWhm5wl8ieGwarmvjp
CqLYYH2fuV7vp/zEn1tgDW2YGXlbMklurk2CTQb1OzKQY3RjQLB4LvCxNH5BXZuOFp9MvP7wBeVf
5c3C+QgnTkQ9zz9upfzQ9c4sMVP2a9S5VQckNEwj4BMqNZjTUYgaFXwp81tjUkLOt+gahz4DUUrW
5z8/liLJ3LSklG2EbwjvWDnwxrSX8ySZgW5Nf2z8hCWqLt92DkvYbyVuX3YIDSu+ejEQEZ1MIPOs
phjSBaZ5TvTME8bFZg4PNRs1OTEx7VGcbc3XBN42WSfZlFBza/Z28x9QAC7G/5wArDbFPUSFnHvI
VRwFd8N5SSdxH/59KGx7LymZeRsuP8p4BffoDmEtkrqo7sIRS+aJ1tf0kIfm1nvvHpOunMIXUubP
EsRjFDvGR/JWtzZLVfnz6j2RAV1ywrzI9x7ZGeVl3K4C2Np/M7717q9HXp6RbkQaVD9OmDoxmzRM
yHGi6L0AuIcBGbEvuSENh4AFpF39Vv8Jo+74RyDO8Eu4T2GUqc5MaYa+0QLPocbKB06EJQ/DAUFX
Iod14fK2jLVPGEoWC15smNedwTmSYDiBtTKK5wfS6uQMqMJDacFwTWhvpvERJlBk0qzZSoG65qwC
a0RlFSik9tMmtUZc6S+ZKD//Fa72AScXSPVLk0V20M1txraFwrwT38KmHvMsztjkHmyC/LLkntfL
5KtO5bXJeBOy9VY40ifY5ZjVlmyPZ09BlgtTllaDkuKsCeLsa9UzPZw2HqjYuGjW0iaup8RP9Jon
zsrZkMsFdsHbsV1iqxC567htdJsrQE96euY5RRAg/S5fHJ/ollFbLeqt2gKde27RjCViHdwVH/5N
FKb0ocfnx8MJlLSHzhoDXtTUoi0OvyjSiprCfW0LYEcDgvIO9CPSIq6/NOd0hKlunXvLLOqw6myU
QSt+WJuEZb5tyjpgl1fFzbF9cA1AkTDHco60ln7cC7I/07FB9R4Ntp08Mi6DMsNubcfSK/3FOett
gk81Cdobpu4CYheHbH1v4388RTCvgrjG3yeG+cOUjjqXJt98lV6o4isSCddwJe0g8EpPGz7zteiq
DHblZiXoOQDibPAFqBp+QnmzDiHPXclxktdrdq3X/mYMArZB87mM8qiNGHRxzJTxlW4NOZryXBtp
c9Dxdbf/rLYSb2wFCEdFwHDGRxGUKjyowGbrGA7846L847IIqBXzAIkPCCSzT37PjpgOPu4t5LWJ
D354k/4EA+bcm3UHsUEkkVmJ4jY8wOf5PISK3P4UfmeSDWlsTw3xe3sMlaIps4iIHCCjpc9ZmlfA
4Bd+uU0f6tB/5EFynxViVrJSWNfUdiSr9PcqTKjVDwsYyoCrd6VhzKR/4EYcVARsDY8w+k7ng/lA
ooCAm5WZqDsV2Id3Mv2bjybd6GRBntchJquSoXgoGp65oBlPt3s7UpwZfzv4CzVRM5m3IlLIyhKK
9WpqF4mnZRydc35Lf8Tmy5hshqvQN3p6cPl5eJ5UT1ABWTlhFCwpOuA/O9wFlx14DJgwctT2eGIG
k0KIZgRQ840d6hAKrjgKBqTkqefjgRfyscEsGiUnoUIldmDMUtpLstSe0GBV/Q2o7hUP4x9zJsdO
J9hHJ5oqQaNEHYL2WbUYUmBechcR4ZOX949oGQOkYM5z8KFLmX1XhC8atYS1T+7yFgwWv6vIF1ie
eTMGfhUkBgQfzjOUB83Sdrnwlg8b6Z5QaHHH7YxvzOAbtS6O4EBOpynI3QRdXHQOCpkRF7ck49gR
5d1PYCDPl5PB9c7xgos7zB+Bgpw2R1HKzmn/i0Bojq/afR5Ey9GUWuF/0ruHi+jt4cK/xBsawiaN
djnCOLuhnAZklstcMM79YboewZ+vOS7JwDW08Z3zauwsVe31rYHfgqf11xswbYw5hkciMjLTRnAF
7ic/kgGI26M4uWsG8jl6vkuLyZtsyag1DMX7lLguBEr09JkW1rehRLDvNfHm16aopV28Mzvo5SlK
KEv+Z48ZjA03tYDuJPbP5Rm394Bge/hQUj5OiojWIsLgZ3T7SLCJWPARa5B9N3MGwvfYadRaiCb1
QECl/Gvg7SImRjAsFJPFrQXlG2vyV9bwArpY/+VJoDXd67bKitPZXpwlYVUk/UqvO4bnQtWmd8NW
2LjhlYK1eRcMd+BlR4PS8oFSyD6ds1RcTi3+JT/O3jtITxb3xhjJwdtgC4AcEvwJj2UKMsutd7fs
IV7IAcW2ISfOpMgYLwy5Wcs362yga2OMDcjZ8EwqY7PKYZa3xZB4d+Ptx/5WG3viPaczVD5/9DjZ
0MmFXgEX9tHO7u2wsIP9zRiWBTQyB1M3ZcAdWA/ltZgWGEEz+oZQqlBpaRIF1Z5iynoMj85IXx4o
re8GFSd4aInXChUlEB4rLRV+CaCeW1eoi0168UNFAcRx7dcjexlI3TSY0pE/2yZA0TZkImU5FHHj
vAIxM84YS41bSgJe0oS0Kl8ND8WnJBJQ3eyYQozJxlrrnZZDhDz3Jg1xMpPs/DIBX0NneRocB9iH
6aobz0tzRcMUGKB7127wAdodVBKxBpru4d8Gt6p4nwctYxqXJBPE0ZOW3tf2exCWecmJYqtfqrKj
w+80DQQ9nYko0AYlo8w6rV5H9Ugpo6fBg5VDaK2yy40LM/jwFVswhHR79rakOwYYJSSMQ0f/feQQ
BW51EJSOYKmdnVRM4xN9uq5GkvF5MxHCMsyKwIwF6rqEFWTPmNICYd4oSUK2gqqHhpliLbZMz+yA
ApGWqoPelURRwa9a/3/q2+KdRaxLIpBT4JcnWsuPeeH2cC7flXznpWQ2Mu0s15owTCzOqtnA5tFO
2pxgZm4lc6PzmjJVYsIKF9anuwS0Drw0Yf8o90+yzb/M7F2nFv30asLWf/sOo9yhKUCyHZWWBpBF
4obKmdHL+0z2ro5olSt4LCdJLpWSTakHwSM+xU4J/05izhFwaKGFF8cQoCOVBpQxhARK368zy9Vr
ODsnGw2rMVeHaDuYLd3tGhpFLfNdVOpbG+M6DGIJFjbZcuJF0i0Qi04IiLXIYJ9Nc3k0S3BUR3wu
zZrUvF/ipfhr6NVhjY00ey2RNXD9dr+TL6BhLFrxqde9Q1IoHfT/LWsHHqsSoVWXjrD/pBoNbAwi
QCp4
`pragma protect end_protected
