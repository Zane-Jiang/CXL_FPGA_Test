// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eR1rKPytU+0XUaAOM2YgLMjSusbBlwF66ibQ86g2KELFnfXJ98b5k2JH/SE2
ZAPAH7hSxF+mOnGv/xmml9rTqBvFZKWSQ1MLwV0BqRjxjLCTJXhIDGyCIfEJ
8NRYcWkqNDekzqn2qW0E+NKKFRPi16L8/DCvGpt4GEFz3zXdDL9rIRXq310E
7MkSt97Id1dWnmddKON0MqH1wFZre38I82sDb5g7nwrPF4x5DW43kY9PhA6y
6QfswPcmoqPRCBoWoof+vQE4dxyX5W73/6CQOGN4053q0AefPiHSkfJ+X4rm
KUCwrL9iZzkh95no20ZkhQNmw6Ra4CXbA4YC6XjuaA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BuQQqiTqB6bpC05tA0wu5hSjUHlywPmvjkU4gPxMDioQ96bnEZE3M38gAVES
qAtlF5krUi7gx0FT5dFqKGy7P4UuwbWqmhypnYFaNtbBH3Spy0Q7HpqsQ/21
RQYZoKDIagf5XGUsfJrj4GWfXsEA7yYdk7zsOYf15k2ZjYlAk0fxWdfgsHvf
N+wYymxor+baB56U1d0qNxcBjoGT4ducAavMqSsLqmfV5+PPnAkuaKbSQUaE
YH5BWl94bLqcqv8bjaFIK8MJd25WTi+9Jm3GkeiQDm9nIh/uXeNGEp+FKQst
T/d2l0vZTmyZ4ti4ZAl8PNUlUAwl35MwIDDiHDdM8w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KidfwXfIWCHVaeboLi/FLgpEW4marXoCVu6INDgaduXYQHO4cSzQlryll0dY
58+Uf88KwDjZDbzhislzhWSrVG92KbhV4AGk13GbccFpZLAecL8BktEkw92u
74KFR7t2OdpZokqzcFoA2TiZX42QuVFPMxerdHoFOOIn1u6JfgWwRUXICLlr
sX9dSfyeu88xS1iJ9MxyTUvPc77cmqOoXylx4kbN7dV4hx1mRF1dZIYbVL6h
M5Z1jPxuJ0aXssSe9B/joPPU2F/518KJBxjc4vOwYxPhufVuws9srSAoNGRY
xyBJuu1RiLKoo7ZW8EZ9ohnMUkkgPdEIrZWxEKLpVw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sY33kQd4OkWziPa8aANU9uYlp3N8QIgMRG3OlhXHhCj7NlZ6JTHS58IqDO1h
qoi5oGtnrQv2r7BWctrp+1YyTylPsR/IjRVNkik47/cVanM7e0Qe7+qBwC9x
yHFt6ILEUs/icsBxHyK3gxmPLQGKeyBEJ3SzjpeqBE8c57hyJOE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ioa98xW9LDBdLnXAcyLYWR7s16cdkvKs+8HRyFuaJ0If/QUlqzbNhCrtd9p4
Kh/8PNfHSeq0eeO0x9qxXbLxwChW65P9DnNTeBQK+RSvoyIaLMfODYtSdkLE
11IWS34fnJgENUNJKxfr+c02e51U5PoYsmA4J4nXpWOCGQopz8Ylkr3iuAur
ga2+D8TgGmABjZzBuERGmE5p+cy+MdQChSxO1loxVt9i8yCHS3yjym4yPZBE
KFceNjq280/QSr1p8/DZRH9ixZyLqQDZl/cIwBKfm6jrXVHka41Wd+QVLy3x
tMj9Qwl7/V5N9dh9weml7oAJLbHB5KXX3IsETaTJ6Hyw6Cp6KYYeg6f3f/OG
AMCZwkGcO121dVklSgduEc6wP9548t3KaHKG/DJJclAbWwOI5WnuSe6ymsGd
4esyUHiCLAC1hA/QV5/3p0ofpgAkgEezVgn1AcEa7en9EIt2X/ky5kheJ7Jc
P/ZNaaGHq3h/ZtUIyXA38bLBaSdXgMMX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cWKdijaKB+4H0HOAMs4zlLPy4vWrQXOHXDFviVw3yZh3m8aXtldxV5Usxlfu
geLt0be+44K7Jr5fJ8jJVDs2xB9Gb4n5i6s4Esok1+27fvnOELv8YoIjZHFe
jjRrPOBeDiUn2Sd26AsHNM8BtEAGbla51DUVTmz8KSXi/6uywCE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ds6T5pnZrN2mB8yvSBRJKl0rn4MjEmnNdrRhV9Qu1EJ3qTUEdApliUKutB4y
F3heQGmaZ96zcqHBh8/emKz098Kbylo/wITsWDphy2pq+68xWFxogkyCewMG
znLIXTcWhp/QnXxlx0LjC81GJFVdWJOyj9INtfwQUaPnAKz0Hc4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 73920)
`pragma protect data_block
7WeVcYuukeF7t1yM3jwcpsX9Ga62EtuqWXC5CCOfl2eNf6awE1SK+/Z5BFhR
oG0L7pNDvFq2CrnRSy3SojtY/S46rF6CbS/xK/ZlqonWjhJWgS7HqFYCpfC7
2a6FB0E0YQKmQIIomfZOiyMCitggVxegQGBgf5TYkCTzVx3PHVeqsoIxu09O
NQPQTwDnBV/xuPk2CfkFvpeLLu0cRlQOaWFjsJwPbYANL4NBrWtShsYTJU+k
HZh7YLux7owfgjUA15g+c+3sUw3a4A7eZC6sbf1wXI+/3N/3LsTR/JYW4aRl
uy8Sf6aHTCyjYP605py7slgD1ZzdHrRVQvW6im5QABz1SaR4RbKQvxFodilm
VyDbsJoOrHQ7M9NszX1iAuRo5kXgGDhxGz6XNneDrYCJEAUf7Z8MEMeVdaVw
boMHxER2GGa/6oGSgPpJ/7y0fBx5PK4pv67Ysp2y1EuO1tNOovQHYWv+OMYn
EAsHtqmByQTxYwVtrm4ut34i0u1pLbGVOSgCn4wlOTdxBxz4pphnuvD5j2jc
4y/cbxEhgo8IWAlqGZNYK1oesRGHD7/KYWkAqLBu7rEYMbacT8y7M5WqzoMO
efQOdWa1hF1kN1tit+v0EXr2S6QShrdLdqysgQRu/78t01lLcsufv+YvJjyP
z3S4Yldoy8E2Ut/dehCzz5atbgoherIB+mlTTuCejw4VM4+btAL/0vpQR9It
gv5U+yiNmWd/qNYjpe8iv2MCpe2MIU7dyT9qtRawKA5lI9saIRR1RH8y+GHN
6osqn7fh/n+/FP/1iNktLxFGq1fpajaXB1E7jBe95/IdNn+/pnjx+1tYpprr
NazM+Thy9PryShCfF87vz2ktIDlZuF90MpmJw4ynKNduLOzTtbWz0LNdisPc
/sErXFUIfUztwq7jsHgOtCIeM5PsUMj+QwBApAkqjj9kW/RAWqZzgcTUdc+n
55NOtjgFWdsmWig3pumElu92AOoElJXMR5gQxvQl/+JbVqQ/ZrYVu5If2ZwU
CCOlTVvhTLBWIr/hQ+99Z70xVRUY1Ew5t3U9Cl7/uV+DOLonVvNpSidK4rnw
ZNRkWcWKEOf5H5qQ/lBmCXUBxuwarrI2jcfGMaBRB1rz2GkOQETkBaO0zPwr
zv/qCFCgyx0iv/zQQpgZLLZDr1xYxzrcmEsF/iz7cumLO3V6emX726cgNWfc
RA9pYTdov9YgWARM8rF0mrYcGqzZLodCLT5/vMEZRbUZe3kj1UGS7bi2MV1V
WDkzeGyFqbEK90zZygesqDiSCNayehkHqbdLpgg6RbJOpA2e+5tXRxHj4HlL
WuYxf7/9eGitLfGtNvyFdGJfsh9THNRvNwHN6xy5edjuwJKGMLl65cwoDQMv
iAcEY6dS9iXajGtT1x8NKSUaAr62zwkJlQOGdjX6DGfgxFXmL/uzinEpn/7X
je2igCHTpdc3piuhhzDiE1tMJi5SlnsDJBTtjDvCJuCtpBO5GSIPmX3jTwZV
ituxZoHKeZNRoziUXOrNMaPUmufLAux4/+SqwzTg34M9YVhovRJpqX4ZhkOV
fTlA1wx92gxNg+VU3NkxI4E8bxB/pNyddEuHMazMSbtl5tA2FqW8SEzQrr5M
YvAOQ8yZVge9C7mA0ZUmWuI0VsrbU6Z7wImvUfbKDNjfFkGGTLPK/+8nn3UA
nn0IAh7n8HtM1XZ3YnoLbwhjrNdYblIH5zS/j67fHQYbscfTLUlijXIr2BRY
H4X6gzBed9xoEYIVM0bIk5nKE/RPQkAuaB7+DKc96BJdlyOKYg7x23IVh1tC
8hE24HrNvdTmou3bNZJUI9zokyKdHCWzXv8QbSavNyYDkrgLT7qeGQR47sct
nsuRzb/roDEGH+ndpk6o2hfIPr6ZK651D4kznqlta+59RHAgOnW/dIebzem2
aH8Okoowede+5XWQcWaprx2c9iGS1Vchc3SZBDYXY9alMtLWE9Rn4MStYzla
ijWyZ3llfRYdtLitU33yJRhONMsetNS9tHgQB3a0qmr9tQZWwQpoO+xfrP7S
YnKvljeKdcKZ75T716puo9P1xWZSJHBDok/Md7EC6VL2Ct2xxGK7XT8z0cuU
1+gwcdnAMgBsyMYIPvJd3nA3x8fSYqruKjLmvgXbjpwmdbFWsXweHHF1n6Sh
2wXTm2tVBEVLHoDMaAvbeZygyYHGGD9/I/8pkDUH2+5epQmdam9PJBy4t/OY
o8PaoB87sKD737VSFrdy4gM6vXBmLOkSh8JWrPqIDWAfI6m+tZKkb5LQztPT
dGO0SYwWXuCaGXH2XkRd4bWiPFGqzfq//fawlfWLZe6IDQbgY4CqcBcEjKCh
4W4s3eCJVxjZzZ7lXjXbGzyroJKLl8lJE+wOp6UTxSaIoHGAuunqF6Yc+Wqo
sPSo61+/VFYIQ2lb5Z90N0clDzJVlJzY5nbvO8359ergaWYLRrmaTbPZk36f
pFQkggozwgPuWe4259aiyYaC/Q/6TXSMdM5xhdMOQ50uvBDyxqP4yzJ73VKx
egYguIWsPKvnpC0vWOnHgBMb8C2SGkJMxGRr7SnEFizK64e9Nwf6ECQL3XYX
c4Ltm7e6GjcYj0BOsVq+EwzhRsoWQ0hN+wmmKNo+nNtSxdYb4o5dnhHpdo7q
CstVP0noTX1ZVQXaTnBsHH2AqRWOoH8kIVlCLIBkbbflED2k8OPZg+qCRZ6I
VMHlmXn+ylqpGN/jNAa8VuEAwf/Mf4c0FvlYDWdZ93wf0iKbfFyxYtGvFVG3
xSt5dzsr95UpNFlcClMlpIykX6F9YHmzimCd961u9DTBlu1tMtSSwGYhH//H
OuQaS/CQzHMtv7hFujWPkfiWo+jHHoQHaCk7hUGY6JfANxRM8vn7k2hHD3IG
l/ZLgAg1mblNHIArMF+raww59B6jB8nn+wpG2z4GSEWT8yVMdjIV/dJlS2ju
rUqDmhlDfc5n72Iv7RvpDYB0r6jp3BasNq2fvHYs2l9BE0MYWDyrK1z/w8fR
fLS2g+MCmCXcUkvzimtJS74bcX9JZ1/zNHHKVPj2iETnZ3rgAlu9C/2wXtzA
ALXTErNg2qVzVgucbB4TWvaBSRYjP/niYjiRtUEEC+CzZW/rLH40g0LpAlDd
RnkapqTqtNaU1R6R1c3tIxykgF36BweMt8Uxd3z+MpEyNkLNQmLBX5zQxn0b
OeC2IHwr5hsP/adtilQmKHT+l7h6OewJdSzc8nMhpgZHRNlkG2iA7ZbJf+MR
8otkhrMzvagjMRNZxJQbiU6pK73sV5vCYUp2snlFaF+25Vxsq9IWQZkAboyO
XVFMTuaa/d6dtixQ8EgYCjsM3ASdeFcGC+udnt+KQAm4Icdw90ll7JatZvLD
F7Vxz0fA4//nKLCK3LTfJ6QBQI//hCPFwFZIWHrbqc3I0o60BB18oYg2w5O3
XcpUiwPcuhkkF53PgbBzmRVC1BZWBNTTDMOvtx8PuLGGh+S08xs/xSxQemCG
kDqlzoLgOz5yGYZMaI06o/84eRnyZiKlbPthw8DQmkmEGCp2GgTq3/EVLDnJ
dyKBkU4vXzlg+bAzF7SidhwSbVuAv/YnOlyM5d6EebTLh+SbyPxX/TlHweLs
tkp8blVdeXvNpdPW3njh26ku2lwYX1XNy0CwsTBz7iCqcSOJtncROobIiwZV
OqqHRxBUD+f9WqXZirNXPBWQKo85xACgQKt5QalXAP0F5YI6BFts4EYqqm7w
/uRaIvIEV8hXm8hvkh4nqHyDuSRqvoPSTEO4pzn9bhXGt5ZVmy6/RFsYb2bk
6nIRZ31ZtwIQWz5aAUDPRQ/PEuqJYSvk3s72jln5fn4w6EqrswfUCMqU65hQ
FModpu2e7BwBtvVrC4MMFjtl34x8np6IHf9h8DhIqRF3cKHFf368NlDiB9P2
v6RWywcihkneRG4jM0Q0ypZmsLvmjtRKIN9Pzk1Y/lTSY3WKckyoDKajei7t
jrpf0EwQAmr/X916yyoo72XxaQ7jJMnaVWOO7bYbGJDTczKwB2o5QKG4bCTX
n4+4K13fZQWS5hjtRxgIoaEVpkjH74OPbcdGYM3FUMr5MVOfz1l8gCvAZ1m+
9SjXQS08svaQFzX1JA2jEJyTZBWmSOqGdE+f3vcCdKW9Ser+65uK9kOPsIL6
B3M71sJRdmWn6WwAaoydZ55DvozEyNK/EK+Swtrt4R0tPT4j7OFxZChbIBfA
1WrJm7EiBGdaPIS98PsAoduRNT/13Q/u7wq17mTpCb1VfHaHkS8jpnwsNknk
GVjASS4IpBAnSy4mIxdoldOAaFxK1hhH/WnMaM+gKYKazO8Ebq6CsylXs8CT
JF6pXPJ19j3OPLVZdzEjVmDo8QyayfTmZAH4JwaKWSqFLt+EVurTSgujQCEL
DR/8aED3WxupuIhiU2f+CN0SduS1z61sYgPxPgImCx51xN+NFfR1ohjuNj0R
asUKRPbrHJeaN6aKCMniAhTAnodLXhj4jOfuKsTFIWpVaSDe4BmikrmYHDrP
TllgVT5iW96CQAjLtvD81lomXftOrakN8xk8TXOffF0IcT8Thwj25evMZ2XZ
6/ILbUUSx2UlHvFARQACvdd8PuEGi3h3Nu/Z6Q31QSJAslYoggAIVX0fLSq0
11ngc1g0FeyEBleg+sUU2G+QShNzweOsb30/M14haBxUqgGksfSLrffqxvaL
IzUNqOnzgyENbK4CX1QCk6TQgYPnhULaXalddBgRrXT0p/h6eiwDJOk0+w2Q
OmJzT/DpfP6Q+AgzreaRLh4HWRuKoRSWP+0jMhmR6a9Qwg46m49SHoAqGeCN
z0jR7h5SfUu6zrv+7cT5eU0Fd2u72w3pAg0aCPxsVTkmtspwiESm0xKpSRLr
+KrdTRaHKOg1jGO7tluQoUaWpFKMS/lFeQmsD1tmt95Sym0Hs7IKy/NAzPS5
dmjCUMLaQnD4K43F5s+QPdZJ3Wc22jxYduCT18XCoeSO6r5h6giXHMdHaBHH
oP6fLNLq5aL6bMh92pYTOpGo+ZRrr0mQM6AtGm/2cXCcBG0ZHms1FM5JX5c/
YnfetC4mhjBHs7EWyUu9xHhipX6jSicxoedv1Hf3lsblyJHFuR0NktKv4Mn9
RHzQYulDHwSxAd+D7zv2Ji02LbqZDLoSROAsUoPpwU3gy91TwCj9FJiN6Zgi
dGnzMOQFYLbaH/2Hg85uBNnkOOMVe5a+FuCYMD8qanVn5BhrNK2krxf+0tyr
HQoGw174gKxzp8PO8HdjQATWTp1w+PUhTue2kgNFmunypmVm0V0iBKNxD9/6
5EWEV3VtR7G327ZPHOqnB7Em7my4AU9tzDjReQGif09CtrSK73UFqiDV6SGf
TCvr5wBV9EfXH8eUYwi0QvieO1QGp/6yvbrSbDUEst7roXYj4i27NcS2j3tg
/g+x1TPhjLZorJsqObDqBfam4Sg5yB1X9IVmDgsdzCSMidu4m9qNzUF2ON5l
W03PVhI6sM+dkcurmloMSPMin+okYeBld2uvw0NAlCpqhRQMpejyQmCaftC5
ZZ9NhHm972km7cxuiO/pSbLYGJo1rlJr/Z2h8R0kFByVm5CGWruk2d2F9QJR
ZLm8OMBBnhEMkRAnPwFQB+oH/sRqILWuwPamLgD3ZGDkURn8nVoZHY6V1ZOW
OKMX1/kH8CxYcgAXSICBrrNCkwA6Tx9MMr0BtF6qpiEIcZFD8kY1QK/VHSES
ZtcfdTOapYTxjwosFKo8yM4SM3PQ1nPTgS5m57jjCZ7DcX5wxjMTJdk95r4p
znGej9goVdGfTI8faYYmJtjbkIaMyGMvtg/QHf49Ne7+UrS62xrfZ5WOO4i9
la4E/0N4Y4iXq6+UGN+CBEgOp7/z9Q9KppnLbvh42XXz8ZhnKNgO9Vz33j/n
z1VFwoP0upq5yxf7aZy3PkS5IzCC/vkRngB0YWfA3OqCswhS+UnCeLIMAGMp
kfvrvrCHcfqG7abhDQg3fl+aSwD4xL8o9xngIHrO4orGpUJxkVKo+FoaYZIB
6oD0CH2bmrMoJgIW70+LAh4ZoLJt6rKKyvcDv5dgP/OTL0/fKSs1gZ7mwfhL
Lsg2fNJ7le12qaBcAlYKV5fkxPiZTz+Xcfg25xFPwaau4lGC5A6oumt3HRYv
swBoQ/HRrxIDEr8PNr7VYxonADhx7Bgya8N04wBpiBBTKzrwTKfCgRoLLjC4
vNR1yhk7KfHBhsXx86+NbO+rlxIDYYlw+dE9HAJe1QEkcEtoF1iliuD/Mlxb
Yas1dtmTmkhqY2I0pRG7OmCF0B9TX6gYJ6UonI7D8xcS5R5RpgydzDTAN4td
PRVxmvU40s37GleXVs/xYvqpIRst+A0bG+c8kdkxx+T2Vh0uJJ3W9LlA25Bm
s+U0SY/JQgOo2F4B1OGWdjuzTyz80eWSRAxHgBfFSE5IzcfqUK+E+uYy9xzQ
M/d6raXoAZCCEWF/wNvvz4UNlT4x7hYdN+P2YlBh1m3gm9ozWnW0ySRB+JM/
jN818nrRhejIZqqrGJk0Mb0Jmi4jeq65BcsT6mq/K0T1Szgno9JUggglbhZE
AQw/eWPs4iqS6D0J59f+tyyFxLTqowYFJShXIkcTO34EHHCWM6ldT5te7kXj
UPsc+6Fu8wEi/C9U58QmOn+aLqcVR53XtrdYmnRlCQNhhvqAUpsDOUH0Texu
/vDlLRwb74vC41zKuqH0lc9KxkxD6lWRcie1r+XFSHnLuV5OUzz1CbxCFGvm
JIeFLn3aVEJb1QcMVDCPhqZX4uxZGEdS0OTbs/gjhL8DJpKDtMU5xuQzZnnv
DDmBYccQoSkigmZDpzDl0vXqVqPil4KCBC4DSrlGUbg1f+Jupdlu9WoWZe/t
mcDDB2bePiUGEZmdte4Iskcw5G7eEwS+mpNYK8DwSIsYO9suEDjqJSS3mipG
cQbEzfZqDzoab2Oi0GePAZfYK4g8b35mkY1mwKniBFZAjw+dPU1SapQFlqV0
lzK6TBstKjjYz/Vc4mq7vk29Ma0q8ncszNA4jKDN9CCfGJLE6Qwc0aMc1OI+
D81XeVSmMDPfGxzi5glbsHTphKy43pDw3zWYTfRJ2TBuoqo1RN2Ogtor5LhQ
Cf/rDf4rfAhAL+HV1v7/rvqM/dZnK+CYqySqtl8+ueBzwdgAAYf7wAhhiyma
bpOZayGEnOkpEtsMEkeNgPK9AoUKRtDNUZMg8wOISAbYnHTZ+5VPakmcNsme
nzvyNSbmcFBATd3M7ic57DMG7rw6mydDgqf9WgOkKczAnGF9vNULNTuKQctM
mBm4xkjoKu9pICNMIoVqRhjZku83UApBodeM3/oH2v2kMqj4s9t5RNphIZmA
vhdR94FN0+q1nxg9tCIFK3LPDlriOvCu4KorcfARTOJml4Ag2WQbPKgewSiD
s1Fu+OGq3eBgZiNd2BEC/8GMVeu4gcUJTqaCpC4qi238h+UEIujwpG7D+5OC
LqFdDOqGDWYinXDeznpCoJz97qku3FrLzJfKIEckSSe+4zdtbIv6qleC9BYQ
fMg3E8dmt19o1AlTaTbBZeRuMjgeDCF44yFru3dlTV4++OPxlAntek4mJmaV
pLS9DE410f6b4jn2ve4gykNRZ/aPv0R5Qi3ICZfVEE26v/MNDNmCuNCyo3RP
SAJ3U2PU+2KQ1WlnfrKIMXbJldb5PRXAGfyaSw+jAx6K/Xf9VxFSVjPOcx8F
MMTNQ5DoUfupti5qri03dlir7gOyp1x5RVhNxJRMyTeFJ2u9u3/aez2+hmPL
L82tVQkVjm4L1zH6GQEOYWyTpqMzBLkSFC7pxzEDWZhd8N1XEPp3Cg+hDbtq
s/ZjEGobj//PexonD/F6U1PhzP5OrLSGZwtm/TsC0D2HWkJptiLc1rnxf2mT
usvovqnWkR4aMjEcT2RuctmopUvSB9roO7zeDe2PE8UqZlq6j1tbrRo6fUSu
7PeRKi5c6ppWRjFqYAN1mW0mODqAwb1oOdNb6UeRqGAnE+jpIu6Vwk1MVH3X
jt6RadUKKuxrhTox+SwsRqeRP/Oz7d+JoSk6Mx2Iex16UgZB4pqgDvL++ji7
r/3LhX4+4UCofzTbUyZ8BltxUDKPBXOUwVb012SF3MwOC67cIwqEy/FfPyIx
s0VfPSkMQSBGHHn/JtwDUEkWtrtSWKQhBZLBb4uXsHQX0rvk7A6i60gM2DWk
VrbDPLVeByNi3B0ZO8HmTjJlnxMttJDLIfJ0w18BvpX0Ytyty6IxnnIjTqVC
B3EIkDVu/42hFlcbquk/ydkGtbtPxD5Yh4zhmBBHSEe0JVp1QNMN67jRG6hY
bHB1zPCSJZeurnazVvOzyMpNAL/tY2fgWEvUBujzS+prZ7QxmphrM/XlNuTD
63dxHCFi+86vKG91aYecwVmJTsXJgo9wBXYXV4vgzmhz9mdcpIns85lDuGTt
dO4oDQzhVhEUjukYCRK7RUQa9199Q0/GDte7KeUSA8uV2tgbGDXrlwuRPNbv
OWdVO8TG4gdbrjilN30zuO3i9Ye7yNb5cjbpZbNuJeGLI31zZ34M4MwCHLAo
z6DbBRQrEJbg8gIxcbHIJawAS0WpxySvGHLF1EtMzfOKpo0GFvEiCrJ4i4lX
r+KEOPxfxNBuebG5MZzyhvBA9Gxe1S6XhBElfCpsIpfFcdrQ5SSn/ceWP7i+
qStOz9k6lmlnbiNqu4sGg66B10XgKc/FaJ1NOa//HCmX35RdUbj3Nsvb7GXH
tkG4RvEHJeujAjwM/59alE/oq2RW61PPUK1yda1ZPxJ1ej0SwujVphkdXm8c
dcVrjzobKU/HgDd50KZbpzODWyt9O/FUf8tQrewAW/GYJOiKaNf3tfOkrt5A
whlomR4gSacUsS5iTalvcmOeEKhs4dVaKWAviBJiVQB2wR8b5q+NK0WW+e3n
ygj5Z0/CWZYPtju2bLEruSGswDcE6BwFr3ErK+oSNakh5pUc2zbavqTvrlgu
Y4p6e4W4SjEIu0/jEpDp71Tf+Dhong3tGCnV2yoi5Y6Ms2LrAIVE0n0+AS3+
6oMwNhlUOoqOKIpc8KW0Nm29VQgXYU4+NJ9tA+vKeGG5Tnymg250wElRkMXP
TaizNWKRFMqQW+1UIVXH5gIJ0a3BWYGGE6Ekjl5Hig+ww5f1yCEeBaV8pMTM
DClNPjpyScpgTotyxv7Suuong2V8irjyn4JsmylfMToS5zXe3hxBMm+1oV/5
iGOYHOF3e5sXzzS1lIrnSsjOJT319MPeb/5pvT2twxZe2VWhmQ4+GZzr0BOe
xEv/QtWQe1EERN5Up4Z0xTC5/MjHdTEi+zQzkhPWXI+yhlKGGLuIceefCREx
gKjMj0mrY2fqRPs5AyZ/SpxKHTIHNOfAT5vXuOhOvocQG4+HLyFuNoVr/56R
5G0lRHcMjh/0ep5hGqkJXB7UV98VfhA3/WcAyD9RdM1lxkruvwwl6PP19MEm
VH0vyRwBmEvRblRpV4N0Tcy0gwdl61FhnROkarVbOcnUXaR7VMpLKTGdDfj0
8AjONQrZeoX5LIHG7gImJ/K2z6jR9Ie05XSCqZyc84A0NVBWucE9vlQDnjuE
sOivk3o6O2GlHd3260p+wLFDVy0CzH2UofOPONVxGmNPSaVx/Kgc4alt5kLI
wEeZs91KV5G/Z/jKhxvlLICFGMV0Mban7DBbiPdQLEVf+jsHIslxP1rcWdha
Gc+RlNnB1r0UaY1luXNPgUuAq445XUtyV/6YTVx2zLJxM+NaXU21tUuLfK/d
4uvtenkI0yF5uVrTdpds9/N1Eh/vFKIqKi97pI1ordkRDjbRezFBLNqGs9UF
ha9LSyZf7b7Q67TT1gy3DLLuZsc3nmCCcYMvh7FAgzuehVwLXa4KNdxGydFu
bpTH+xLjoT4rc/0kkoH6hDDcea80eEVJRMbPhl43ql9c/yiqb2uTiZiwrRWj
aWJ1BHqIVnSvg8NqjUDiaSEbb2ei5tS1yFmOM3yB+7o9urRFYpXuwHaFmZE8
hslDzTnjAn+DkOCaAoqYiIF+X/EReEK1k5rkjN7B88tJ1HW82IY6zbQntW0x
Ln+6fzfVkazNnNAbv3wibf11mSlyqfEQ2K7leAgr0YRkrgwFQb+4G6PtLIgB
22ha2ITvIt6npSUHKYEk5S/yYK6a45xBDvtexuWT+Ejsfaf0txzcbf2E4ktB
9PQqqHBSVx9WXAuU2upekUP1uRTnWtIRRWCQbC76iNCgXQMAsPiriseCyTev
mzrYyEiEQZepEfY/NPRdqp1uMtQmeDFvMBCHxg/r6lrkS4G6wGZaxEgzkB4U
MykZoZX1bpB6ReYWRoaGhuKFzPSWqxg7XYErH5ooIVGfrrL9aMcXhFTuk885
gnoLjn7fpMSUeKnLHH04dIolJOfyIOK6/yGlYzEQZaE/mTime5fQgouNXEEi
7/6I5F1dG0NewBlVTrLvXs/mEFm0zTGzqd+SC6ukuJBRzcz523G4AB9uH+IT
l3OMmScwLz8UBNSqJctQ5ZR+57XSmB9PvCCez3CO4S0IxbNuaUD/3yfukPFD
qzbe000AZM679DDMpK1FoERSd4p+LR6wEgBMZwdTiaFOgqOWhhvazLYrexOG
TbveRo+HUBad+AkWIdHkOzw+XQ9tBNi5Ub67plyy6LLdacRqxl0ZYGxSzqTi
l0waSFKIHY3ei92YMpOJoKvFKhF28wsMMjmXF1MVFHIPIzk2Ce7TZQGwMzFg
YJ9ZKCmlWFDK6oAnnjnsGKIcmKFD4vKw4f+XuRpoefkR3uCYQg8yG9w6InKw
+aQq20GrhEpqxHj8MXXYL7hl4xItdaqEaRXzK03MsodotrbkkiZG/uIScbeA
lvs9ivz9htCUpyGWVcuynpOrslCAUisCjNy13v0CohdsjRNLwaMmtMA1vFU+
TQYXRaVjsDIRrJWi3tUDvLSxTnQjhwyTtxGq3MkGwOVactSpTO/gdSS/vlOE
d+twQTv4UmQ9kioFMfWBm6uu+jhLNvIhWRDBUhQrzbtF/hlREEPwCqySLC+q
Tu9VdoSk0kOctnI88vCyimjVnYD6f1aW6sTJl4ydLVxLSTVryt5CCUv9uV3+
YnUB9yAhryjV4gxpAMbHzR+FVGp8A/fXxLDDUy1LfK/lJItrUEMZUHpGDNTU
C3Cpex0PQak2DAwgOqzVHlxtK1i/56ilsNiueS9UVhxXyuAEVlr6EMYdMm3J
NqFrUHclG1NEe6tymmm8NnF4PgeClEhP8J7PfRY5roOLwadGOdbqgI22Zsj4
NcRevlmncGwOSnphoPv+gR91UXURLVL9h5LXo1w5MaKjjqj7hRCC+5qFZv9y
dl4at8inV9Y1cq/CA3Jibtn9HpCz+GJt7zGxOXB9zU6sCQCg1/3/xv1xwgoE
GQc2KcK4QlRLCG0UrVxHZlxPVzDiKROsBzzs+fUspkdmcupUVE0QjAII8ahG
DQY/Ilj61ZyzJzq6c/loSa763x6u2oQSsUCD2V+6cAypjijiRyQRco65mhwt
0vzO8Ir9nDxsVZfhQqpfcxkddatj7PZVPdsu8QI1srdl8TT+tFrXMy/zSh0E
lMfXmFNtp5w42HGOddgvetQYBAWTJh12wPgCrp+8ixigNRSP/EHBvDGGZO0H
zI8yXvCtl0Ow0xnkC973J0jqjB1gBTRMy12SvwbwuEOAT2bDctfrLaiwGTUz
H1P9XisBxnqiG+7kb4RO59YTwykrBt5M64N7aNBeaGbb/4xgwNx2BBpji+4u
BOqI6Hf30mbSjwkEU1GLUUtWq9f5CTXG4kZBQcYx6AkBNvNPhYXzQRkRZmgp
npaELMAMGHblGHVFE90j/4/zKVAFBPH+De/GIpHmmuEpGT26eIVMoueToYSP
N/i0N8EOwIpGmWfvq1FKuk6C8zjglvsVbrO4FzWQbIxyEkAm4+/O8Ymi2klU
pBFABdG13+cZLpDCh4RD84oPnk1FdhUUWPYYG6dhiGGaVqGDITM0cAeskIi6
Uof3sUtmFYdsvBo/pNLWAwbCrXJLh5+DXI5vCah0URIPHdvoXmZng+a++ilH
3wYw0+BxRDJhanN1qf5/sCtY1U0/bzo13Lb9uKvvlmvSDPU8jfm3X+u3U2+t
5UhPvB/UZ6M6N3RlyeIrLSHuV0+teBuETR6MWK2etBlmwnVQEDrEAv3qzDfp
klfvzcn53eNKodoHyTHX9fyR1c522uQkqvyaYMr2nbL0dOEcgz/cvqYGSxVS
ZxUe9n3i0hCAiHWG9JO9NV8zJiP1ZVs6zgVys+RkoEnnQrhBvJezlGREKqts
asf2jYWJLwIywn2CJJxivRvKretjZ6C8DqlMvR1T9+GtNkkmAtWQoOEh2foF
/1BAvn9j8WYNkWuMdUi/ZiJeL0981NMbyPqLxQ/S7N6TKWsQYHikZk4q+3DA
8dCjkj3NaoaQk8Si4DBa9ow3i7RR2ie2d8n8ceRJVXlcN3yF2e6+TH7Yq1f1
nDkb+kxgqkrpvb62pfyBExXrPPeT8d1JJc98hHdcKBFdzCcU6jWIwohYzwml
OR8AagHUJItQNOtnEpgl4uq7XtnV0EcLlWv75ntT2qe6A5FOAi1qigczuL7k
A+BwlEccg34GSq7X6yQXB7jS/s4qBgJPy+ys1moX+Laqds+3z4m0q8XP4xJj
pCdNFH0FuyVKKuaD8UX75g+sbiyN+/glcIliNMvPGd6hIU6FFi0vn6rVbKEt
3WjJ9ntvPpIZlRyp+smYv7hsrrHrdT83I6ClOoqdEAKeWF/d2uPiGK9uCRwJ
ZeOTXg+hZ+gfPbq091eaw/KHsvVbexoDdXDejAbF01YR6QJkiIA3UXPaLC/y
CUWFntwXjeOhI1CCBL0EQIV+HUfZ9pE/R2K1gmi7JHa3PPwLSga6ME37bYDy
5YqxFQPqBMs4sN0R/NIJceBI4I8IXXFDf4V0Po2yGPqGsyDERil+hM3gLHyQ
xq3DGcygSugeB4FPUiZLNAMLLC1JxIPGKqcFjpNGxbRYE+OwV14GBRZIbMDr
Fu1NKNMpJcQYAHux2S1gee5CrOVPqRA/jJxMSRAKAe8c/LLZ54DB8Ot3V9Oq
9uP2WNK71Cyeh16NliN5h4IIaJt2bmdEQnF3wDu2UjhcLyL/hgrLvonUKRck
nKJe7Og6lVbTe45OMtNdvYXvUwx3uJx+wT3M48brKKK5ERzjqI4AfSMUF9OI
AF9XhIyv1RBxD8/KP2+NEB7WKQ6MgG7ZHNpcnEjrlbsBTKISqhf+TB+Fy2Eg
FZDseO5emtAjZVBP0t4Bksh/TUn+r0CTEeM81Ap5gsMdOBqJJbfk7iSIQ/i2
lMKcRYcu1EdmvDyJUeGOomsNamU/n+T9SMEteTcE9V5DGu34lthWYTBZTb+E
cK+djAgrU+D7g53rNZi40SLojt5AG7W98gl44IfaoBL6Tr06w9yz4s6xkNTL
1A3ZY0r2BoQZ35qA0FjKYtJeMWktzsfsWpDAkEwHjr4+r4PU9SWNhz/hYyi0
BvfnLbx4wUdUBTbeo12URSXd5Gve3G3eiFAWWQbXBjvGg6m8C6JeSUYz2tjC
dwLsPWbJ4hE11PWo01oeIgda5buj8XMRio/RHhk382RFE11kiePLnCFTiy22
j/bhSY6Ob7N6rnb4WTKx0D9fLfRttBXymSsWzbtu5cM3eG05Zijbq9suA7Vv
+IMJ0v2fgRJyTYG+s4Tth3VJoPVtIu+7YtX7zvlBVmlnaztmXz+pD/HNNZgP
1we7w29ZkMMHL48MTVmehoRYeCuyqQ6fVxkLU5zCRFyDEF/gKtc/jzUn785X
aLd6mAW0OF9QEZMNmWetb0QkSzbt/vCcvVlSVA3Lle1jLp9REclqJBCKzE9m
oqNBjyNxHcNcpkMJx9qhUK8ZGY36UdbRv4uL3tUVdolMOc5T27Lfo9dQDcH9
VU7ZzfESKfwiYifDxbX1rp63WEu+xBm6PjgOjaZn0VfxWSeeqMJOSI8ouFQg
kfWKe3Eg82/2PgLHp+yy6sgJ781XCO9nvgEfvBg69xJckHI60swcpG91HkFg
TwW7BBJDJrlqF8aqtALOmuDygBq+Q2eexNpR+wHj7aAwSxtSbijTvG1Yfnai
HdwfSOBxcfSvwBWTdqNTVc/2rq93/DH0USlCwlhfQIRh/JErmKCu+oHJH+d+
AHUzmoV/hD0JrWgYjGRerJPyQVvGw/gewuM1n2RIC4wwtZ2TrHriMiZPY1XG
S5bXx/oiafMdBdilQsG2zN92sUMx9s8icui0BJg3p+haiJLnNJ5Meu4jlXh7
8RIPfxioOVxS7cfKV4GwMiaJv860GrjlYOPiX8UBh3z+sIgzyVpWVtGaJC6L
brFBISdgekVWCF/uKIJeVgfpS+LRaXGebEjXveXFuj4wk9SLHEyOxsNQUYXy
KqPS007dxztC3kVbNolFo84STQcnOo4YGme7krrn8wr6E55g0FHoC9RYzAPJ
acLYfO8eWwK+n/40BF8bcd1ahEJLUZLc7i/u9PehDrRXkz4guz+KAr/6Cw01
zWwvHg6ePl8LFOKYvpf8kNI/sVgWv21HSH2Xn2uRdoSHkcXhkd3JWAMNiZEx
DYK0THMYjnISxOmagIS7BT1KN21iNTk+tRFde4ugrcdN3vtJwaQnMS38pEXI
Kq81ElDQFduxHOMk3K92L0LZ0/Zy6Y8I8hg6kB2ZAdeop9psxjAy6Sku3byg
RO3dw8fx5wX97Dza3PZ2tb+v0rFFyEYFeL+U3DGXuUAVe0NrDmMLjMhlM4iL
wak+mDsr46w1q3G+2pKyHEYVjcmAidMbrdDl8hJCpXncHYMdYbvc50wpEXQl
iZQr/4GynYuG1ZBjXaQSJNwH4KA4iNbJIv3x4rcvjQXak68MfSL44QTOP/x0
N/UayjZYo2jE8M3Om7oBQP7WBRqVjMKrAAZjVE65KQQK52L/nD/dyOIVxUhd
ugZDm1a4GYx7eLXPzPbP/T/IRF2vawwwAjbRxrUESWlQeNlK1Khz1HHDQQKo
MxkOr+KJy3J3PpxSgJ4x1Wfdhs384Dg64ftVLjIEl2F4k/M4Dcd7dGW/bz6B
2y9M7z1TB7K2WjHP5S91FnCYC/4t8iZFkJbqcjD8JMZRVWOUEczPng5E1cub
uHGsgpgD0dWvNeB+aIXF3vE//ilvy71IHTZQ/U7qZMqfmQK6p69D1EDDNsrR
DxmnJARnweTsVBTNLqposCLpXIZq0GGlrXki1ToZvcr57z7i3fG9GgyE6K2G
ThkYBoZO4HusZfirVXI1LXmqcI4b4FIgerKgcibdhnLGnIlW9Jc/1Kgs1O/t
ci/sWG7zJgqjhDJkheLDAgCB4tfHwtOE9pDk4Y6KjIdUMa/mZlArsy5eJ10I
4ud38VFCc+PMtQ8jMsceVbrACV59uopGti1YzkqaPoHGvehpPB622lTil/wl
R0WZERrex/buNDNz0BerpM3Q1+HTQhcUieF4b2zJ5iaWx55KQsWg6WBKQf4E
c5tod3Sv8YYeBgSDpL/xI1+jgFXUM8Uhy6vt4q3ug0w/3UOGH2h/ZKd7/R4d
CTblF9Q+FkkEneKlp1V21Ybg+V1jZz/SkFpMcD7awCZh9xFxMF4M+EyT3Iw4
5ncPQzdgC/GopiMg43qf69ckPR+yl7OR+ZQf0q639bO9SLkXVPSHVsEAkKvA
rjmxzMdBs3GtzlvsC6i0nwxfM9tnYd397u6zwXPNc17uYSUHeT5ftqlwegLK
khiDAiTbOeRDJvff+CaFmBaQ9LFJHWTEgHqWXaR/l9/Jqf5Uyq661krDl2X3
bMdeRu64F+Adr++dH/wlw7r2LX8DdG4jg9fsDlPZ7XRqAgafFVG4qk3R92bR
X9DeTWnlvqnqeGRtv2od5zUDktg7ZKgzUjadiH25QsSzYkkiYlMQSz9hpqcB
slTgioSnb0CLDv1kf0ivYlt7fTCLun1/154V/VBWltxwaX8nVQEOSOuMoS9h
RQsygCojtVEQa9rZWwFezKgxZ5Wu6NfM7vqiabEayYoqgysh4HHfjbUVKR1R
wtnMrzEjpRPVs6WkLfQ2LVV6trqGUtii44oWAFmvNZV2F0Kg/C9grif9+172
pBxc8iWvdhYja7H8+DJYkoAQ/Kl4/ysSJ3I+ckV8VdY7u7aOeoZxZVFmYk+N
BqX6hu3rsi+sZoEPc8owAhgH4der1GHUlQfnW+3PyxauXyemXZNit0FXMdBs
npqYopEso662b0pBgDZXrrWKBHmjAL9IhwX/7jC100PeDJndVgWC6bIc3VDZ
9dcQ3ourMynG9ySE0mVQq254OlRxMsaXnPat6LTyy5u/zQcmmwWcxauBzOVb
EtwMHsVYf/XmjDB0rjNHhvRR9iA2skJhSGtUaz5leS7jS4C5pvnXu9zJxYZu
uBDHPml2U3Tk2m2Z4NNW7ENZalFUlB1HFPVryfEoW4Q6SXskKBWtoMRflt/e
eD5qxuEtjVmyAub1SaidIp7LiV96INZJwIgKSGr66dCnV8O2zDkG1Lzy30LJ
Zn5ZUOGsQPxfmIHzhbj+MUVk3q6zq7bv0PSsia024p7DfTVJ3QzNmW5zOuL1
Y+SkNqY181/cpX7ycD+UPyYNUDfFeLxbyHDiLBL8wk0U7jMWvPTI8T0TwpBx
qS0ivlFPi7fobjdWd+cbs2k7csyi9gm46OKtJlDWWNc6vg0jiLI5ljDD1pqi
UxvxsQ2N2Yt9zcCweE+K1Zg2Xqi3Wtsztu+foIHHY/ilfbjrh3DPEhOGfiTC
MRxV7mrMaUupu0M7yRgFDVvmh6twsHqAMTJCSOiUTSNuUn7pn0GMWFjMPkDN
7xvTv5HxAsVm/bUP1vzG8rrfefG5WoLd63mUYtx7InWpJYIUXH7FQMrjAFZR
nBSnqJ/cZmMmRASeM38Xd8BlMNBmOvPyw4MjOVE3k3T4gg+1UB8EnxR37kN7
jTPbJGmLWUE9jSXagV+73eAj68qCKpLvKNWG3Y778guEapFpWrwUdmVwPNcN
nYTg4+bNfwUB7uQ0YjIAJuu6yfm5rSUwWrCy1GoB6L3RRquAebmJKXW5M5F4
1Irj+f55yi1BOY2wALm9MbSK1pvSnoNBUIDl8kRhB+9nvDpN/NfbqKCfvyUo
cMnNjevwCsPwESQX6mCViLVDEKcqU1Fau6UZ4cwm2LXAuqaLUbCr549GJhQU
jFHFpP22yJopmOT/5THQlDJupG9rfBLoRndKLaWnJS3dNxNKD6E5aTHbBqko
JHNri1uCX76vsKG73sWh+IxdTxllF7i5mw6Vgp+tzdJRfnhVXE74U57XzI98
dYXfosqSoW4AdGJjR08JxsohqmaKb+k/BIlKRJGvrTJ4H6sqanarO7BgzZfA
HCyVcQ4evepXIKHEWl4AGkAWDCRR5pZ1o0sEvdy4Me6ppCyswf+gUzQDfQJe
RBzuF1Q8DE0NQi7ig7YfbeGp4uplY9vw8dA7nFmPQ4XxZdfp0o3I3UkgwZp9
FO6803N7wRxPaS10W6oZncBsJV7B/K6vYL0KLAkp9983U+wCGlVPu7gUdyRv
f83mlPGpT8qrL81tB2ALomqvB9l0oohC+z3QGoqJ7qzhMJOR6mcS2PNneYZz
FKn2HwJ/c7s0sAWQDo1V/lRopFH1e1cktlZ+oiCLxihu5Yunnav0w5SgcEut
Of1t4eqAlK0WOCqTdXlaS+xtFJxSdKpRSeSgFYdLQpdtNPg1NPpU5Qn8gJQA
uXJMuXB82ePSBIo475wR+vSt9EgbdB7J/goXo6BqPUgOh0SGix1zVfXZUE0N
e5Ea62DlXgcL4ci9a+333tCCcgOlpK7myrCnmJftaXJp/YYd9HyweDexoeOM
IZhmMzgiBZr92dyE51rC0X79RMalqRMBzS93P/Z6H3/TH1JR6+PG8ZVvL7Yr
Fw8oK+NzPLk3W8OVOJRW5afRkzosJErhBmwMmYEjPp+aVrquCt6yrwLMPHOP
BCrjXa+UZ1FkBFS8Vug+Tt47JIJYpH4Txw1UqU79nFrpRuH7hMaLpr4yRp5j
2SYrbdfb84VRTDLISlWnGGVuV9heL+WF6fuHHoSgHs7goVb9fNguH8uROMbt
BL75Lk0LM4SLsGlz/EZl3k1s3nQn7lwMuVIbNlOqNgfUSQWS7IVNpI5ulLM9
zMKtGiqkkYoT/7Nbq/QpusMydgEdPy23s4sBJsL1JpVFjvbLo1diN1WSnKA+
po+fq4RVQOye+V5cCHFbLUO7tE2yiafwrhQi5/NE73qzrKcoqLUCLfTX5hBZ
DCZkMKWFh8ec2/7YTqLOCbz7M4zDkMtMrBeAqM9WQeKhAPOX2ZGsGEQCaA5+
I7xC6nbB8G4/k66u8tA6KpnpD4PIJWUGgOUKFs79oAKtU5K1b1qR74vUEwTw
nqRt5BwTDEl8wDrZxo0vIm3lmGNFWKCocDIK799CIVZdxbulxAqnVeHvpIiK
GDeML3y533KekHKrV3mEiFvU1rb2FqfcP4bGZPSsGX4LCpvE9qrmeYB97aVc
mCqxBVK3PyFwSoMRXU21Zh1saXngyIrv3qWSlFJS163z7nhAW1YAOu7z5z6v
gyr/WszZqT0x82QSusu89AjAeKlbO5IQms5vNrt8kQDgzcU6/y4X3pbCWSYD
gAgjzNwK3z0Oyw3kSIZ+n3d/TiCcwziPbKgtxLRI8Zag/jmxY5egdVQhWHrj
WPmYR+ya04EI8rW+MAEUNDA8EQglURjEtCTIo4Yxzg0OzbBGHTVui8ckx/eW
R1dxvB93T+YczsKBkHG0lU+KUSyfJ+RbpOGaA6XUlc5izjH7YDIKS4TJQGrL
bU6AaXj0Jk4yB6sNdSiKHrSCSqAJINoR3pHS5U7kp6TpNQ1IiIAmvDoRW0Ed
FXB9c5qQrw8mPH/00k93S91eVasXBaDBNnD3FkUrSwccAFAhnIfpepcet8z2
tw/Ktch7IBM4MP9c9XXi0/lQ/aE7Ayguv4WaoJGNgaHjCVGBQhmVbLEMulm6
W/bjNq5z9yEy6o+s/zkJliNirnOO4ayEUk54On2E70857nmSBK+1k7OsFIdk
D73Wy+A7kIaCHUL6Np/LD75GWKVeDg0aiK4ayW2fotJLradC4bgRyDndm3OW
PunjB0Y9fo8AS7dwQBDLEp1gPd/dy/CIq+zJ6QUvFdlvF1KKmGWEk2UUTn9w
Jyex4ra1woPb1iYg1OJ35Cdrl0R/lDJDKEk4LHgQaDfc76ZFzwJvlt/soel+
RFM5jJBqT0TKz7TLkxKm64SUaFb5H+PEG4yL/bC5/6g4NW5ODnrT5kI0gSw0
LoMUbAtNnQgjjKW7bOeLciiONlTppRsSDPlxG3riVN8D/wRcws1+ML+ZwDiO
X4am4qsQO00V/qAY3gHIUscpEz5u9n58TVwcJfamb8XWCBawHV7dvwC/SvWu
xolahsLp/jU/3oxvYEWQPUkL1wFy/kLD1QhMZoBRF9sP5U+0JfGxUzy7pCOg
K0VMBg88eI/OEbMjJ9KXB0O58noKzmOjyW0lzu3LCBkXTFASvb9IvHf/WtQo
ufrzNIPq6EPsctbQH45KMxlu3M4Xdch8tOX4K62B7o2kseKa37ih+W7Ulj86
IYNvsnNyJ1BkLUri02+qO+sDLDaVYd3nSmmgEiqGe87OqeoVUaeDwkYTYqRD
YANrw2w+TxonrlmiwAYBLxCJ6+itvTY1Drm0kGhMfVcL0ZFD63Xh5jFIjpoa
dENe5GdpLNiZ5gC3f3yozND83U3OxtiIjm7RCPJSUe9hAYsQJBlih1+7A4eT
GmvQyBza07BjQ3i+ynHDL2jYq8MRJA/6zrDPUDEoijtZwfmpObuOXyVrU1gZ
r1ZyDzjdMptarIZP+rf1HDzVQ1+mq5Z4W3ZCgLdLb+7k3EDTy9jI/adio6ss
pJre5k2Pb+WL7/rJGUQIgOeYjqOPYDFc++SVUB1EzWulAFhwT8dVkfQJ1Cx6
gVZrw1FzAfH3qLtESCP7d/EzS3XIHYWPTYMay3XqnjOFC2oYBI7AlPaulPqf
VeELkfqCuPXnyhPipMbUtJ0+6+YXHLYzHBY7zMDqLiGmxWrS2N/b+pQzdsdC
E+iNDT/Sr8rFl0/KyjzYmDcvs/mIlXumfWhFmoL3iLpk9FN/C9PmINldLNo2
wkF2g6yb1V0mMuZXKN8tikxwvdywRBVwAIy0LexYxy/bANiCmh/SCRg6r0TH
fKBLNoj/VBiP1wk3hgNwyGix4vmBZsKYRc/DL1kkm7Dr6dkk3gXqwf63UEXH
xVZxjRU5m+W4XWrLKMG/oGFmjFeRUQ8WQbcjuBWoGaAZgaogoZUeIFRSQVRf
MJtIT3SXkQ6w6fJlMGCIJsPaS24YFMx+kJROMNDEmuG0HwIfX0JfxUzsJcI3
Sgl1dqVQd7IJXZkF72I+r1it4plOV1zZUu5C1f3SU4mMSYweApd1w2sxZJCl
/2PXxeF3676ch90fdfYRA18UP90dY0W0nvfWMuQ3uf42uKxR3d/+vJK7pVUD
c5BQ3ooTFDQWhwX1uP8EcfYVLHvDiJhWzBXh6/LAf4Q84YXHzSw3v0FwL0Wx
xn0Z7eI2remcZJBuauEDMsjJvBcJ73QoUZS8Os+mC60JpA3mDYJTVXT947U8
3NoG19DiWxw6GOWfvjXmNZspr3OVAuNNHV8ojD2/KcgJv2zlTiGkjrj0uDYO
RBEl8J/eDfTkMv9DRBtg1PCASvZJHdqZlhK/Y084+9gedt/tAmLfpIjrzIk2
Wld80AdORLC3IGc06srexyv/dPPGnOhrvU3q6rhQWhQu5jGQpJa4nq04dpnn
i8YPtsWUOpyo8wvFH7KIQJdBWEc60HC/LsIPo+tDbQbTFknifYgms3sGbCKV
bkTUg2K9MD+FryOpxafwBWee6kx7NND2VDoXOTWeTTQk1Jwdhu1NvQY9zXLJ
HvHzB9WWzlVjYleTQ8ZKDFb0GSOjxHEk+nPgRAU0fgxT6G4H2VB/s5zn41JY
MWGPiTNyW6ZYMVbykwzHYN45vyw2bclpogVoSDNuIHBMBgCHU8RJ+KYUf1Xt
YAvZU0226RD6/Kt6L/iNZUUke656YJiHaxbPrVAjkmG8dTmbHl7SHfgIQw3L
TuFHr9a0E8sS3YIE0l1mlGxNc+jzu9nSt6sY/FZGoniLhGHFHO4qe+LvKhPW
eGC+TXEwBLCIHvxdcEEtNm/l3Ml3OqrstBtQku3qCZMvArT/k6Jfy0Fo6411
RApel39jqKMTzqzLbxSaPAMahU6+9R40m0/nHJncQjlNys8rVBwsStDKQaA0
lUtDcOLz7w4MQ+lvP9zQvXneoKI4XyHVX1pPmZ4CmjgZYWWqG6LToSkKle3v
N+rDcSgPbfTACu/8nW9QnIgpYD098CLHBotlxWCHCZRz0xDv+eH/65cxcuNp
ks8UO4JWpW9zXlX2a2KHtaO7TxgZ//N0xDi4NKcCcJZ+m/y26Bo/sJ2aA6Wu
s2rpROkKjvIHCG9CRLKT9PUOXgQ/ryyxojc77Fyg0IBp7iP/LzBZk7j8cY53
ck/WwXiJdnWuj3SOXkKK702NyG0GTVi0USBzKG4DFlrORmGGJCVGa1V3bfjY
rzGtegRTjYdaoVXJtH3L8WHR7L3mXKl2caO6wkBZ3kcKt35H/p045eiz/Gca
P6a2dMMF3Hh8hhN9Q+DthZjfnhsN8A5VAz8V1HDgCftzW2fD0mOG2JGisZg9
eZCEW81C11JftRK8IrYuR/wPs03tv+Peh1nN2KrrRxvGLDV1Kg0S64l/PG22
nnLaaaS1JEc3n89Jgq+kbgrSySk+i4uGUFx6PP6exMBMBaxvCBshmcXMpFKK
/t4jOGcFEBAEC86sa/ltEpCKNVL79WgpAN9PT1iYkcNfLno2T/3VxjJtGLAR
oYYeYNII4DLtsz8dNiirjp6caaplKCUp+U0+f+ptSBVvIM0UvHwdP8UycYbw
myr7jbUtqR01DQcTHo/2YXOkWGWoE1nKIOSsJMO/dpCmiZZvrN1uA575RlcI
jXuQeG8Pwcg7nODWCuylGunykyxlEdfucv/Us0b9Pil1Oel8w3CjxPByDh0z
AZJP7ca8pwzyNO9b635Ss9fJF3hdBzPbRb2qPkVR8aH/W5V7/hJ/Xs9cE0te
vMfnzpHnPT8VAa/KSJdhyGmeIVtCAZIBjAUa7dbF1nvroSG0a/XuX3+K24+d
GOULRpRbHu9XXrTw81xTbFbo9l8f7EpUSMp+r+1vtQsLo8/Y2PebFVCkLfac
boeSZHpJaRrZC22yCf7zdGkIRXgcXm7mnxR6tTONjy6gLHDEN8N93Foa43Pf
Gpz+fs/9LRs28Pp7iqSEGZ6DViF7KIfQzHI12JSwT4d1n7qYw6Op/zrzi40j
tfTzE0XjXpwbMWPUEZoS6UGsCqP/Cw5VEZFSWcoZOimn3z6tQ3WWRW4svTC8
jkWB5c0Hob7U+sryD9GZspK8Eo8Z9QHVxpiwILO8OLunwrjSTUeqcvWNV8UM
hdnt2r9XxKT61mzU8uMG3vR6HrHAxeitgu33WgBLFHu/UUgk94qzm7PMmfT6
PJXg67+Er7KiDKuEZ5f5kG5tNCbr7uc6ChwStXdz/ZN/lekH/2hIeGrO57TG
4OoaDBQng9ezAgG7grd6g1WblKdEHpxNcUZdelQvh5R7FdxdKE0PBNEfGMFg
eD2XP/hCN7pEKGTmFV2UXPrYBdQUpsQiC9R26qSfa2RKsUZF4Hq0Ond3cpeW
TS45jJjqlGaAjmxdESTnqx8IHDpGOqx0uN13xelox3eRgGXiuy6Gd1MUn98p
4uOnuOki9CfsvfzO7jEPFjSB0McNOndPPnzFfEB5lJEV+7gLTI5LOkEfEGtX
J+w0uCqgLvUTis3gkYydWqZ9VdeBdc5TNhToXkPKp5GEzZpwYzHpcJw5rKko
+KVdnpLw79MMSQtrWfl74lUyTWyVxSQDw2RO/5cfOKJ5n/3/287LBzN5fmGf
hw5gowqt0/3OeAa38uDWtOaFQ+S1rDhEg7nq71YiMxJYHUnmgKhAkVd/75la
9BwAHfaUI6JBx95tfsUmCgd8RDnQq+orJZrVvtkXAcI7Z2n3FImAj98SfW/p
vUP6nEZPFjGIZyqgkT4bqeLIdEAk6wqqqDIu121iYpOQzLgJKHumDESve+LC
ZgWkIhr9+CQiMarKtmvGDLgZqEiDzlys59laGzIfTT2LO6s/Aw4dDkImOa9q
LlH90WhhanZNCvA8xURizjxjAkb6gi9Nzmlsd1keD5Z9ALpdbW14cwCZjpEh
akN/6U1UFzpSjHOc9Iz2hbLpqq/x2LqU6MAVJ26G/jjvsHTySL4IhYTDhMqC
MR2zQXucewJvMeLkTVSvdCBrFIlbbViTsGL/qApZFgSAU8kzscxyq5Qp9q1K
TWwpN7xSFwMsBGBJ2GGFWXiQtQt8ZCD65JlYqk22EuAAZPZeHmt+0XqL2MIg
SO91CzQ0WBuT8SM325bIdXcTjTaRE173+baGbpN8Cg1BwtoA0KubcE2z4DOz
zZaXVUaxiY5RdkNZ7bGQF8hgWClSHwCONh4Feg983z9axuUZtU6xtLIhyiww
w/vf2zJLE77PdU5I61jL0JRYDfCnt7KLOCqUbQb97xjWJSA0CoRp4GV7xGlu
x70iw8r4/ngIBFmMrEROVxhwNySTaBoQ9EazIbY55mlsdqEO0vXbHjJh4lPi
1KmBB6xObR8f4VqROVow+jiTP6m+PYShTohyfUZBlFKWonr0qVo/GbC+vrQU
wVwt0ABFf36LOLVT6lTsr7mIx+WAkdc+8JoPL84er/gu1ZpDtNiGGB0K4kTI
nMFHzXiVshov1LvKQvypl6ifrq3IsJ5KjY7TbFuS3HCVipcADj8dTvcwb7Ww
9ncN7Z/dkXe1uZBv0GK7+zKyzNc9BODbCRKcfNVIBtbdgTKuIckRvK8Hg6q9
vW9pD2X50EMlag2MV+ASPsCl88ioF46MboY4WmoLjH/P2kU304hWUbQA1ia9
9F9Lh8Fd6erJDfyRGzrOpXOeTH66CRprsPExgiktwmHkMLXyXfrrBnAE8KDx
kUX1bnOU99EpdWzIRibmByVGg7b7r8RRbJIkiX8f9DnPybIA5/5h2NET8zE4
mI0YmrGu7goVfpRixw+gqOcHnPIvQA1os00hC2yOa7u9BlyI/EDNMBlZ+x/v
rYrSR96kcfN9NljGapEnSzT3MELA88i0INK74iBCweec9HS6HLCm9RZZoi6c
J4O8q7Ka7/Xwg33843yNA9zU0+EADS+dcRZx186rfWoqDoh6uH5zOcBaVZnE
MICqTe6gY/zsUYtp/AbB4/VzxE5Rb7IiMUdVo5Y7gk2plKM3ANjccgX4sIO6
rhe7Gk5WZg1Zt5SGTiG3UCi7I9uU0urCn+JQRC2pfDnb4Rbt9a75UHQPBktR
qCuGSo/SKLuJcOoYZZ6onwDWJfEPCtTwHZcsEuefXjq3SXPKlvRMYJvjhI3g
U5DaoRtzAq+P6oV61UFSDBPcjMAqjHn+dyFMKTPHkqEpc090zgRSOkNCJDrk
ZNFGrw2K6iCpKtc5LnHyGnnX3mrcffYB46qLzh+cj8MaeZpFGd80BBEjZbR/
7oorRvNYrmwRJ8pOwSrFGYIF32pmLD2IPtiVq9lcSz9gEELfRtuPUoV430jn
eUEhpWfsvERWpX/18ix/crl7B9JfeT8zLr1/whRXQppH+yF3+dlZDtd67nIn
5r99s/hCc0NWxu9apCvToAjdGXTPdOllf9x+TVgYbvGG81SlXA0aGxHdeCSp
7Bt/Wr7OJYytbfy5fu3zjXc6D3sMyBzqO5L7TmHoWuG06BKuos4AGtg6n9RA
iCQrvfE3VNoxHUjWS6wsq+33wGJVo8jcR3fMhl0yxBW1lgiLO6P6+9YDhmnc
pUBzenKtKlGRW3oJ/fa2g6/AstRu+QtOMazVSRZSZ08Hnq1TS6198h+S1tnv
X6uHAI/yKkPLhlTu66uWMbeFAkpP8gVsV3D5K4TxuOh9jVpNxQSBuLYbcAd3
NQU+J5+4DMnI1VeLl4414Z4Irfyrlsj7QuYAHKs0RHIs4dtLe7jn+Vg7DgFI
lC1lPe45B5/MCWJA5BD9aZYbuQd3x+coRM798Pmj86FFGcLhUzB5leFafRUA
QkiE16fK99NIzmwnH4XFCm3JXvfnp73ECZdhsEqpFveO6BAxc9p0pRmOy8Cb
wMe4FT6wMrnH1Fr++BRXYARQGbAZMe/rdkVdeuQRuFjXnkdFyx1vRFHv+kre
fonF2yx5CH9ZwS7xGzIPox793HZ0f8t9h00RSNXHHxAbHBrjF93MXN2DfA8s
ln7NJp+IoYbyTuO2gXAlzdq0ITS10BNxTGD2MAvRQ5lHlQgV14naKEVZ5A9n
vN+uZxMDwBbFfG5Wwa5gokgpJ/VBxirVIvXDwagKsSiMpcabOEnEkD7+kJW8
ZiCgp9R98OUF/bg2AM2S0RL73KdwG+Ax/8n1rNEgh0uteLpkH2L+0N0XLLD1
PCQitMetvdqLiSw7/c+joKTplWLvZ6fwTce6ALjPXHhoA+g7k/oHLcMw6iI1
17M3RBF7gpFPas8h1jxsSqvcmkFXq7wLgBPAMoP1cAWscWh6JwrNZByOOOsC
zPTrdmvbDdWz/6bPORxtG1pCKrfCiMng3BFhEycJNR8cI7TQfffv3NlW8S/c
S6H7yi+EN3xyZByVnVTaOg+JP67Seb8zbHEMAv/LaCbqvf2vbLsl8OFVKqFq
pBr/MMUlFk1U2LBmlcXGiaB979bsfBRWoQCStVCQM2T+kaUTmmWe1Lbk5Miv
0dVG2jsS8y9NNqMADbc0SCFtVo6hkPI0jRDq9PiFUEWtKnD6lN7UzU6ms1z/
7j+YKQYYXRIrawgJLIB6k1GxVXRmGZQsX+uuvRzpi0XPHurYcMQ+52UanX81
fqrbQ3wMpCuCyzuH+OLyIIGnIpYXx0O12tsZ4Lk7ecMtvpSGVF/SP6QyvliZ
cEF5Wknd3IuXk16CK7hBvcAACkYyX/5xPkQQJbHY3DBNU9VmbeYFYteDe5Vt
F7Q1mS0glaAoRLumx5gpcRinv3iFaZGYpZs+h5EW6ysEGf++llUlnQbgGOiw
tcVgIkAX+ZkL0ocM6gF2CHrA6IKTPiCkbkoagaaNgIdIThiFaG7Sqx6zkXr2
o3dXU4/WI2+huxWQvoZBoHsE3HXYqMf5ymgtG5kg+mwNlL8Gb3h2bLP0BbmG
dOTaSjorUREVD+Vz1802rPPphgiL5PtNqkrM56UcFJYNHiwQ7hDaFPV/X8vs
YLZbafICn+sD5xC9ci1JGZ8NqyuaOQfsYlS7xAAq8BU81jNh+ZZK6wzVkYQk
dIjyJBzccbMHxv8/2W0aN20HtLBbGDzENDzQj/OWarNW4pVTGwpysn/Cy6vB
LDTV4qFeqg6vvFKGqCv4BFPAiZ+3qGPnl9nvLDpwvr3KnTDOe0VDxkp5wiQW
bUn2o/fqAYTizbUOJ9/eV8ZTu8Uel2u9nIItnJ6hGKXcSUwQfOTivO4UKa1J
L7gRz4BU6sQpFb0FjPEaIFhBpgwXIc8cUeZD28VBjiTwTgmG4TuX6covyJQw
DrJCzarOQSmOUhkpwcO3YOx0iPW1BmUC3gGogLk7XlF8n7jqEFskCzzoHXGw
aHtQ0flb5E8QHSkgQacupnRjIIMN98OPTPWXDpHOrPMQp+5kCb+BjnN6o9tz
VMhvZSvMNWzwWl7lrhjkWb6jdU7XrOfh4sTS1xx+hj1s0RdYvDzf/G2xkQue
SC1RUx7a6ntm+80GpkyBJ1YSTNRQaZ0CRwX+D9fXC8RoLT1SccqGYZbfOgmH
PFP0Ip25758x/PSXRxZ1rKNgyomSiAIG5LYajoOUeRc7tUDJlrV32FSaNRPU
mMVjOTvVxuek8dEHN2Iu+Q9H0pLPps8ZwziDwqa5rUUCx8zHFyt92vTtDKY7
3Q6/PRsDa7TNJXBhB94FiIgWlf5OfY9T/EKbxcFNsjWQOjtwEin7GqIfmhNx
D+58XWmJcQImDwCIvfrb+Y+yEBcscW3HRQU310neHQ5juuv5vFV4CYyii2eV
KJ8sKdqMR5KYFaXbIQkxG11fEWQ8VLVPtWkQtahW9GOtOAwJGR4jlGCx52BO
M3g8ydPOVxTfjrcVNuc522wZvTThAzXaHIt1/itRExbUcpiErtSp8+eo2uVU
BFZnCtVxwY4o/hRcN0/rG8sn1DTaEJyfwJJL5kzkD+vk23Lm6cpZ4+rew/nI
3xGlSJOthJlJVMtLStUM8U/5MTh9+lBToFvOwwn/kJTVFkx/+n9pbvMuwa6i
VnuvcCVA+3mr37iX6jEVpQvN7qHA+HTXVlZk/LER4yDff0ZmeXJ2T5c6gg0N
/+ElyNBJMMtxIaGoI6xvC8QpOo2ikHXH+rtLuGpR35fKEEhju7pKQ5B7uVhN
o2gWtn7mS3su/9ursx4JJmuTfs5Nw//dIcxe0Pj9gCQC9ZE/S/xmFunx8Aw1
Y42WhiiSCIy0PHPQLJ7TZ9fyiYdrwMuto6fz8d3CSc4JJcdcbqbJFeMDki/9
vXLDycq5ERKf2jN/6cR9znOaSPA4mH+k1WMGxwgN5OfVLlL/QD89vZTVBW32
cREvDetRhXyvfkKzgEnujTcX7Wam9Nq/Tv0uAe7yyof32elwnD5ZPaLZxK07
1m+IBKkg4GklAQSx2pDI7AJ3vW9xlxd5VddQJ6WGIO5HJrq7XxPBl7cagBmS
M6GDx3Qh1vPDM3rC29gOyPFfEwNxs8cTlWVdjuTcrx3uiylgxc+EDLCT65v4
4Ibs3HMxz8EuOw1pH3tc/R/sdW3k5TSsoUxq8CgaukVoSf7TD+Mu7cPhWSOE
330LO5iTvTlL4LmPE8RqxidQzRp+bs+dR/QcklaRL2SgEsj9SaRymQTIS+HT
/R7/dWlET2NRfOyDJlNcEBp2q7dVipUOcr5e0eET8Ko2gHkLWG8T5w6O2Koe
mr+dhPsxXxq8S1/aVbrFoBywllrSC9HWfeR8m3KZqjSn4d+9dMtwzRERcqhu
5y0Yp7BDsTTBlZkYXbEUTwowV2Fvif103eViYLR5jplcG3XdOiil3Jj+FmL1
PPsVVYvHIrRWi9KM+ujGQth7UmL0zGJQPZwgDDbrZxDZ0D+MqC5ROYmdRCTO
ciHfYum/kZ3OJg1xP4JGrek9DvemTZZT8LAwBmXr3Qa4Ln+AJcpBE8k1O8HJ
leLA5tmLjGkpdFYHQrWJR5Xnt+SWJyhQVtZcR9BIy1JBcpI/xz4Z2L2PKsXn
uzIpjfA3p5i2ahaTDO4JBSpWCnj9hx6gvceTLnK9cK3fE+jVGvdyQOswmb26
rXz6lY6mlctaeVXUk276S8RQI7cNCKbzhop2UAamyuZfabiu1ZoHIK50GheZ
kXWolipg2HVWZ84hiIbkT7QF5DmFRWkZuTZgF1R/wPISOK+G00lFM3e9BGJN
V4g/5sd6eN0DWCH2tDRFfrbYk+/leIRrbOsdbR9xs6SMKb+CPzArEDmBaFfx
8ZHeGIRudKfYmCU1W0aXkO990c8/d307rEeeZfxyPfo7nW5J+CzR2RzH9Ym0
YYkJCSD6PMC209Kq4PJ4yhaNKu+6yn6jpNAp+sizPG5grcqR4gCgfGHya6bD
ALTojIHWZr4aT7i+pgREvVs6VLGFWav/StE6xCDKagqQmh9TYO1pCenpBUia
s32bQcwhwT4iwTq1FrtUfj30dDCVBi3mpfnRdaDDWp6dV5+uIt/6bk+aKJ04
0J9ywR+qMB4dlRD+obfnEFlpFFOmgMzrvXR3ewh7Tz2uzoMJBOmwHgc2l6Ko
6kEbXit52ZtmQ3eYgd7i1nkfY2vu48xy8Sl5A/20ae1724gltkZDL5jt39XB
lcixHrHJXTvzoooUKGmkJESTFub2Xnsz+IojtvLZnnzjDe/KX3SsVGmeLZek
IuRly4344NHBWc4afGIi9hqoWFWsfMv62EBR1wRkJrztGrdBameftlKbW9m0
ISakvlEjjQxBQqXsdZNRqwYR8qmLcUC0hQzdDiYOWBLc3L0ivPkK52QF6TDk
sHweqQuXkhW4Ww4LpbyWBL6MVyMBLV9Knh5HBiYnav/VwC3y2cuC288+mNua
JQPSC7qYilR5EDpAJ2ADN9UBuOFElMwi9fk83gWMmIHFnkwibrX5O2pOLxKc
V/pSw+/bpXGyhrAIoi93dkKwesp19ScxXTKGqq0KcbF8xIHPjYJMyIfjLOX6
yZWpNWuQ3mNdlb2KiQ118JlSnVye4zncDpqapMTOKXIxEPq3Bp1gv7MAfKb4
tCoGWwEEROYFgmTn/ZdUSmtFqd7SqOgILyRvr2YapWOD8ogvSRyQjKO1GC/a
NyxGyt2PNqHy1TfJkezdYKsp4K8f5D/B8zu1MurnrDpC4gkJI7eN+eWzTt8T
7uVHtaeuaNiF45edhSAQ0iw8h2AIVSMzft+oWsyvbr9x26nl4K7jvLpzmPIx
PDBzOWB+N/P71UWkYIbDhROXcTTPA3FyVNgZvqJr7zMqt6dm+ECiuMHwltvt
sxORs+7dWiA60ft7ENT7HromJLeQJEUIVwR2ucIpi23Y+xz/0xVlJDRTqH2M
8Qo8qyuY8sreZFahgENLiz97QoYyfLKmNAo8e7LIjuAvROVlrbPS4yA+dbP2
1hJ9dyNiM43gxqX3e8Z0HQDHq6v3UA/XOzyt6OnFLFV1ZDRR16+m/iLS4l7r
1syPj9/uSngPP06kNp49QGT6mFpAqWuhFxeVkLLW7tNfcFqa6KYBIryrIurK
n7jApqSA0Pew1eCSD0dtpAXp2QMivHustG+5CABDvWOaBCvhC3tQSnxP0ONA
WiAhsUoAU41ql44QGxcIgV1pZyMYulI+0hd6EBVSw8/YMlbguKlfMIgDFVRC
Und17zo1xCyPDNuOflgFv2XMt6SLcgvsvDNVpGHFfPmHsS7tp9OB/ezEkwnY
lQeegmrVz9XGxqzOCEh7kSEOmlWu+BOhAT3BUNzVQmaD0p0JKRMmRn0eTlAL
+jrWGKzQx4tAOIs2efkyn+Nx61xKT1Y4k5dcJWWqIQpnR5KWFBDbDKJ3M5C+
cvMtyVNOxUGicayagUQ7pik7orPx9nGOYd1lEx1BmItQ/fOMuLcjF7zsK4KP
K7ttmLax5LdoPnVBpb9CMUMM1ehAQVX0juOXXvBzA9dBRaW08PVUM0ZKcVLE
NGFfZEpVfSQ3GlEN+MrJgKHiKBZnUjsHo04s9SbB76527gkHY3QMTi4g5qtX
xtgvLTN+Ul09PpRaUqGdXcAdiwzQgRqWkL8sRYZJrnFctBVwaqRFogKqKTFs
eu7cDGsykoq0+idDozcYnZYcbiIQlwszfvyEOLiDhEO0P/RgKOOw9xE5CGLk
GRgkXBOtv7tpOL8JUOVF+gHeqFKDk7OPABxCYCmE8S8sL+L+35bEVleHzPKe
WUVAOGZF6uIXQrLSruCAcjfPBBwBuLwxLKBCJb87l6NV9AEEdCpDGlERXeNp
I1tE8bCetaBYAW2qx3kRR50JGF3iSjLGn+lmHAYxeGvPZrIfBiSdDDElFFMf
b27NmL+Z9TNEXqNtIlkZrtSvABEyl+5tOd4jPe40PqDYgNOXsF/xr6djO+/e
u1xRqX3ec2Hmd2tmvojsNl4Nz/2rt/Zl4O5NqvHI3C9StCSbqKBrnWtddNTP
oi1WF2EE+GqWw6S0X6DvhiDsXwHI15HkkwlunON3lkt3rr5voV8qc390XnO9
VPg/8yaGskB9ZmQQX9kukiXZtnxeuYW9dKg2k316MoEcYbTXiS//aQT9nH78
1qOSuvTgJ6PtvjFe1M09sigTwAa7T7jsgyhAlt+yf7Ze+G8sncpsu6gI6HT+
IZnFAVNIfUyne6UBWgBaAXi0ly6AJA7RocD0TVZmZOmirnh7KXbSHXkZj7J4
EdN3nKVG56QtGNATFsQ3ArvuJ7bWJSSboQQLweesddACxY/iUmU+nT6Cw8jK
u+8bR680HDC/SxoSEFB3RGHAhoMROz1uCA5hG9jTb1i5LOe0bvYMlY0wCzhS
HdOHeucoiLpzgw0Vun1eT+5MZLFCvkfl6FcrbwYe3hSeuk/HuTqKOtcklakv
TbVPaJeJhjoocHVhaoZwiVYHSbgycQxS9yiEPOFZaudB7ZWcPhG9mqD8YmpK
WtdAd6tM+XkuIyE8gajDSgaC6VYHpgBn9QcgOZUkjOazrAwez/+LXMzp2j43
yQNH3cqyExrXYGFwlqjiJMnqSbmjFB6MGX5My8Nti9WB2A/iKzVtblAx7ufZ
uPerDMIjQjqHsUh/FsRi0dx9g3YVgDNl9bh4MMYdjC992cu9+b43+ujyuuKk
OYkvSTOwo6ZhtwAUNhw9+00QVjzhVyVJufGKEtZbNO9g1fHdBxJSHmKR8oG8
M+4Fc9ffYDCh/UozZPDySe/I5fj09mP6eYRO34dSAJ9T9kpYySEoSCUmmjKm
TE5MN62Xl8kISkMfyimnHGlftMJ1bJ2Q5bHU7RB9IDMTTYJVVA6SpMjPE2L8
3mB6U2HU4mGN7WUVAwqhsqWfaZOdxK8RXdTSDWxe7lRd0PHitdrt6dUHGenw
uM3eIz78O4nz1uO8YrgRkdPHEQ06Ril1sq6uSBYjM5Tq7u17BPnFJi2igSMF
UmbCLATcP64i2yQ/CUYzKWWLUq0InhTy9tfrR4X4iZJ7Hv53VfhTdG4ZfOQH
UwUBkIjcMjsfEGSTvdWiAMPcCNDoEW84zG4MbZ1fdNb5iTwaaDPkeM6Gq4UR
cYCqNqlcAaWzXh/T85vQAgPKy+P9+GMP6WHuhRfHKHstPt+3L5EmHcH7WlK8
jllH9Xb/sffRFOithGznMx3AXvhxV3EHeWB0bVk1owcU/RzNrUjsC/pHJW9q
Q87T4wjpWD9EtoaZSKPWHwVWnCwMYBczcdXWjK2LO10PSuqg70QW4gulaaT7
0+XgUm7EuQFkRRd45QobFrXP9LDWTGzdlNTz0oFgYhwywYvonecnsNMd9A++
XE63vQIophn+p1SeY6ePHLBzp0ir3BU0+e7Rskc/IFBbFtikB9oO45o16mKG
cIrsZFMbfTrWfSvFrm8uy3wksmnkkSfFlAbqXkvrjKdi1t6gyRdedZ3YvqKt
SvDKvM/XO92bDnoyCC4ssiPEkLlFNK2RKS658jC7HQFTHa3IQLNB/Ko97aVH
oSGNGz8zlp5ActvARvjqk6rKrSqXOhvNtwlsZUMc9Ybj6e2hkz+bPoDZQAwn
OZxaqm39Ob2hGcr4fXMqUNp2xhBroJcs2NUjD6PK0bYo4VLofAzdYNvUCqxV
WoFGe5WQz3NDTGZnknvl4br/krc9MP7pRPloBMLxD6Uonc0a8V/p700q/TIn
Xx7ZtLPyinImRY42VL2M1RQ4grrclCLjyGQDfkwSHXAIlL3N9nzWko2X9DdQ
xOk01qZrPHDFiDjlxrZjEf3Pw+fuaTY+nCT2d92DUv5HW28OSX97gALU8Dma
gb6D4F9HHFCgwdUD1lG6hA80URu13A6FrYdE0xMxAFxcPa69OqpBXvXjNHnc
Ak8W3xggRNULOrGLcZDFokyUknU3fma4j0WMsZvhs93qSwt7PW2R/UHF0NG/
OaxPHTO0Y/Ps9oK6gSgCN+UB4UIDf7GxFdleqrFpU9Cb0vlQo455XYa8hOJ/
Auv46Ts1HeNTA4hYrdb3YelvnW9OqmJobSTND3fMeHoTzJnBMyF6g6UqiEJT
rG3ErzeStiW+lsepiQJhqeZNWYvRK+h31CJD2Xd3m/FsCK4k22Go8O9j9f/j
sElXbTXOcIUDe3FwV/T2Q1QmZYGTev1XFGq1MRE3LvLBf7L82vSZsl6/Ry/D
vD1P4kufRilpGTdrP7oEKORI2rFOzHK80nLmmY/982O4XBP9Dtf65lhfvnMP
+s2rxfHXOPlcOz6IOfelEq42kwXbU7gTf+yI2GKjVh+qrUQADJpiAyx5DAfp
LGbJ0yF4pq/0DEzEnulkR9XSLZwuWySPUN7rjJPdkG0eqwj5LJjJQ+IIQqr9
yvdL2KZYmopBsCtxWaWtFWVNqllIPkx9nA0+ohOpfMCn9xpW7qthgUYoJIzP
XWjHkUNPuk8eKKhagY77OQPzQDnF+Oq0TVQqBHjAGeyIcJmzSYODeUQ2zcqg
dAjGATaL0FQIb7PAlyB+0v9w+S21ldtETqukc8PNstlV+OAdUaQw8gxRjwYq
LJMWdjct/BYda92wi1QLLKoYcJiVZVZAUJMh45As5+VncWckXzZR9eFBOz8R
eVlyake/9h/RWq425B/TeYn1pdww6XiNqHMUcFRwUijKysBMn0y7foZZAdSa
7BPTnqP3TzH5TygpqFes9AcsDjkTtrakJg1zTV+uZ1+/DIuxkhxLnTZ2xyE3
JTvEDR4OipE8tAkVTQ2WLM5a9jwq6BPQTMXcG611ya424Owioys/NRLrMGLL
BHAVwsj6oY1wnjFdTD1s9/GpxH2VMatHzGrJ2r8V4dzS4ykLHFYwcrMABfRF
F5g9UVUvgboZhzsykXq2YKZvjtz/gh+MiYW6nsx5CgLi5o7R/e16r2vqG6kS
78CIAQf4vOMp02m4QaCZ+X4OqhxdCYiRwoXXeIN04fLi3dO8oM+snKCwvAUJ
fR/5sHB7MDRnjOphnS3hDVQe1zGOW8wJGS/aCnUKSPSAHsGVKtM88W7LQgmV
MmtdJ16i4gBcMJ0G9bk4ql8Ia/ENdWWv2mNa2zFGUDhk8s5MOn9w0jlhCukx
YjcPvUbYh/AI5N5iSTMWDrSXVyspEpxHRxaWocIK43T6Qy9SvJH1pE67O/4N
uxa7anqzp6dULaf718gYTzI7Lasl/cCUa/WDnb+VIjazW3N9FCUGlXWQoaHu
cjz9dC9FQiinTAP/kAHOgTcBS3pIBEM7UnPkG1FuwXeZvuAMFPuL8te7V65L
CUoXeiigZXSVmBS9CYkKpp5SYECcOWFfHx0VUYCCZBT3SANHWxlXG6YJnQh/
orFAH5NbCVOg5xgCar4JQb+x1Wy5B/pWIYyLK8zZuzZMOJrmctYxDfl7R6zp
n81Xmdt/wPIIHEHXXdbWVGfRrKqN/wtULYFiPZCUS2+SByP0i26gt3crdjLE
nmhHXKkjwvl7tx8cMaGKUSn9U7fOdIb6nHmniMzInT6gxpccfRz7pdUX0ZTO
ptrGQBAmWEjgcwup9jYhvD4dYAIZiyQcTOzGjdpypSe2CArFRkdQuUlRZG/0
nO51gFw7JtZHPqTzVzfMqo2SRGi1IZqBx+R3bhxc+m2mz8DUmeBgexZdAxPw
oW/wGXIKQzp4/VPMlTuEhSveCP/EWHwqU/fsiU5xK7ERkUBp3f0jm7njCcAf
ppljTD789D7WmNAsZosgd87S+hCU25zCk06LH5yYAY1YFRlMUnrWeDGRd2tn
2PE6zCp67v0VXvRrBkLb4lNhF3P3xKPCR3Q7gbAHjEsQG5CilBUdsajlWMZE
FAGdmqsggVDZm0FmuMCxA17gVmX6WfQs9ZGMyQ4qFEFBZFRMFxwZ5lKOdBd2
0Yy1VVojsPlS/HMEswsUQwi3sNqJl0G3x9Zlezz89m9WfXjv6LRc4vfWFs37
kAymXrq9o6oP36c2e0Rh1EaqRYhfLSE8XhBUblDQNwjxdOc3paUGKgF5s8ug
bfMp05JKWz+cPHVQjVgjKQXRfsiMscO6ZnP0EivMJKpCWkGeCLFaceYKfrym
Qn1KZSvY09WFYxm2gT37MtZ7Vn/fWmgv6DkVYUih4whOoadYhVdare2a8gji
hAfrUsR2CgXXvnOggDbdybakc2QJy+yEmsJxNL3/Cl2e2Gum7IjXzeIzX0hi
fXLyf0SnUAdxnxIr9HSUQJRqK9W9D7yuzkEqTWibmn1BbGCwDGkfCb2NHDjy
4cIQP/p4j6eQXWzrMBN7/ZcQCyvXRcAAMEwwkWrcet8RcP3GKVGOoQl+ho0d
0VY7ffaHqSVw5qZo039A3YkfSBzVL7QhtwG7ykZUl/5LQjsU5G1Hb+BKIcnm
9819naeq7illBaaSRT6Ii3U4bPQZ7xCPOUyPu877O2RMWYm/uH7Zarxs4azF
we/YM0ONHV1eP06tZopIYzurpUyqXYXWOKo1ssDhB3EXd/fkfNTwYPvIayE0
+BqUdfqkNmkCr7vUz8XLuNLKHxlpTuMa+w5H/W6KMZsmH17aZQbQoJvIV4EA
2LZUcTybwQ1QUdym3MzeFIua+GiE86fPeoYlE6B2HUDkvep7oR3H13egYlft
9Fn1Ano93OXzx2BYtMR3HTm9xvQPwfWcjUjRitZeARV/pcRNklYPxD+KsDIa
BOduKsUjh72Uz4tzHhl6sRTNm+ZO5wZDr1axd3Ew+/gp4xa0vTq1WRxZrVEk
GxYJWOmCPY2llMIAWD36oKu0BRhbwiVbwovXzHUNPf6c1Kn85zg0XrgahuSR
wqCTW6oZ2fsbySGM7rtkyxfYGaSvIWyfo2xv7aEhlCezKGo0xqnkEbHud2Nn
CmEYkV1v/rcozz8yHrcD9w950z0SMBuVs3cOGespTf8QNWYn9uVKsWNTG+rt
fC2gSS/CBWmqfHzijGcuGahCdXwiiHxd38Fpd1864Tt8V59/HcBUn30/YaYI
6tRKkxXmOJvONaBazstXRAHUGUQ9u6H2WDLo8Ah4u00U7gHzeXuXqHifripn
NjejQCJk53qyCdVyRg959NxnFCn6IZfNrYiD078Lss7PD8ZeAm0ObUjhjTMS
KPdTDcQbpCknj1Gi3oCcaJ4EZXcQgjYN6/QGuPJONMF37tDbcy1EAKPSUvMx
rsKdEhE8J4e1dFfZuLmv5TcULTEJP4hzIGISLckwBQRDcSmESFUUr9JTyLPE
DJaMwOYf+6gwpfpEd19HllRZlyb4omCeze0D0MMwEppb/UseIw5+4Q8h0Aek
HQwt27bKC8te8Gf/jY7KsfHLVtyxntoVUzc+glax4W1Vw0uaUIo8M81+nvPN
i1XgnkZRCt0TSa0JMULJXJjQ8hXdFN9qTsi7ZV1YTAXdjYlHlDvxCSrAk8Lc
tDP+MYC8ey1SFHJr/77xYrVZmRPOS82pR6Y48qPwnfiZFaSJe2zyFfoekcN0
BMbqm5MuhrEUdwunK1xG5h+bJBe0tfz4RjfXjiJGWeOpUz09kG8UkS9ifp6l
LJN9ym84NRvKFl0YcMa5x8PdcO+Uscen09f0ZoI+QMFXRtxVIHcK9+oMU9op
HfrsIMEZD9xLESsu8hBpqJP8CQ8mAnibGB4YNM/cggF0TWKK8ehSxh8kzQUG
c91zcV8mTImJFI+QGZl06P0NpU0rTqYMdh1hVNFzPKqy4drRiciJDrHFG4UZ
VtsieeUwllykJrRkSIAPqqMFreMZ93LtKQCxG7OF0jWoMtY3FkGJ9snNmybc
1XgVZ74xt/Om45kppp90KbyIhQrDba0+IZwxJWlxg6evt3b+VrhNm6sYYx4F
rOBdkRgIIRLh/O2GXC8LHE7MysBqY8gkyJMsjhfdSOiYAT7KsmcQcq9DaUub
Y4pHjXhEbYkU0mLCrSSUxvDr+FV5PB8sDq2C/cIvx5rTkksfoLhhs5gzVIYH
fXWn+mxkhAh02+EDocix561HE/wyx8yku0j+WYBaIPAe2PQ5kaVXnxslHpP4
/5ihKSjz8Z1q729SwMHjbNPGMi3vpn86cuvnpfgQvqh9mwwGwXxu+pkQsRh9
HluaASM5aFnRT/rFgzum3HJtg/OMWLHVX3h+fcEL/A4ex4Jm0v6DOR9w3sO7
98I7aofhK3xRjLxi3bwpL0cVZS7lPlywPt9gy5x8Nv4YLPl4CjL7caBD0QIs
nfZ0bECIl0gryc7DlScKAE91EFlDf+/HFbMz3ITfv5DOAhYTmjhfOLi+Flfz
wY3SnAxZV3yaD6GUemoBjsGZjtcgRU0l+WrlzVdaPjMEx2cII/LGHHzvWbj/
ybzkz7NRt3+lV4P/8ktM2CudaTMrWnWxjELCZly1kMguZ9bVSQ88K9mxZR1U
hf7NQ0rtExX+iC8y05dN0wUxWXS/G1luA9ELvL3jYLYCKTjDYblmk1yjZEwz
fQiCexJmHr6SJfNjAfn/mG0IpLXb89PE82euEJNhjz071VlF5bnPohi2u+NP
kmVW4ihQ7/pOB9DgKP+MMDfkc5H8ypGDOREXeVdgTMT+3WCU635pdBCn8TCb
YHhqMP78eBcht5XncVfouzT0x0aatQ+BTlQ7fCZ6bKoBrpuIuQ0/1w2slePn
rP6YLKM9/HnT2UiozS7xcPpJLfXlx7P2JBD+0/VrueHEprfbk4sHcKY0QjVl
2hPLW9ycAmI97GzyPoCaYNama0Ycm/9wSoRzQE7EBC7XrwefGJP26QTO/0N2
XiHZR6eQJA+0KNKv5TB90AU7M7FyY2olIpTfeH2LDVdnBGaWH8uxq/Wuq/iI
y7AM+wa73vYWoscw3RTA7bNbIEM4lGaAgasTtjBqADEYt8FncIIspHsr80ZF
5W1jMmz1OqFzpyOGr5vZQkzWOaipWldncd8/rPiaDVe9mxGHusOHMHtoNOnh
xOPwUpeb0Ky69W6PwdBYO2T1Cu/K5JyMx5tsYwW4qzWm2ahUW5fpA30wIh92
oZ1apyRyQm7Yn7cypiz/vRzwBFtPIBk71Ypn6tHWYiwXCtNvoYShnhzr4hb7
sLM22Wglpru0RZVudHQmRRw93+JQK8w+bv5lrzi7wKZEXUUH/+I6+oVpJ4T+
3X/qYSfDYZueDcLgv8YZNEiHOkd96bxERKPp3IBGZ/K0UlzcemufyTx4+7Yk
eXmfwR12Va9xygj7bb8a/9D/nkojCqTq68ZVmg6Xr2gjV/lmhcIR7RInfYqz
W2xO6lIheLwwIrg7rA+xSuKOMPF4SsL8zuDBLUQp/F/pp1BAXy22bx+4ahYJ
gYihogziF3vEC4FgQ8HH0sgLyNCaVFXT5QgXAIZe6Xqv03qpCpOlb+eSeuS3
ZWZToowr8n87pjrMwad28Ysti2Md+GdZ3kJSfoSTaA9AeM+wNDhOHE+wvVsz
zLPGiLtbqbItSinreDDCkKg6UYDMCcgEt+8N9sTGDq7S7n7yRcm5mGBsSte0
7T0MYYw5QrL6rVc6eQIL+1O/oQUehE+NDO2xXZxNPHSI7ZUM6WjCgXD/h3xo
MgdZOSvcAUfvhWv3MkQF7Nrg1KKjqEgTvyNQVtjNZlyxLcvwqWWAlZpkgwNT
iyc+I6jycuy1mjGuj62MELGkpCGSEXWrbeMchNUsKdwDMWB18Uq+lj3Y8Klr
U2Ts+hRUbvjW1obKvfxdniemn65BN7DPwECFG6ZHCp308hYoOgetpcU3DsVo
j5BG6grWclVmiWn7FXlQ2dl6yGngfSV7oPs73GsRcjXyXUMv+2lsdT060E5p
B4odYMZ9dofPmgOAJw1TvjMB78QN55H7rgmPtaFjlb+zJsqjLTBK1Xurdv+w
SS+Ac8q30giugwVyRJjnNKQUBebLNs6XZCghwJX7BkS+fv367sjL+PaSVZe0
l3S3rGN5G8QjLdyriLCnIgNtBHqFAJwSu6TIAh86XP4c7rWE8hL/wwlfjDP/
bE0+plT3LyDmcdHYAMJ6uFIyQl8+KV7EN44hiDKiw814GZJgNw9yiUF26lUF
DwYE8GqSKjM/cbnslG+QwdVqet2NRnSQ4b9Ri43SqIO0wag/IYm++3Gg202R
IeEXw3kwB6+rED9i3KIJDi4FX4Wn+r177Z/QrxVxfDytwgZRATIRvVp2mnQj
FY3R28yYAYuFjUzNh6EOFbuHKOBJzOGnioBW7FwSk+IbbRplDBuk3K7xY0hv
Y2eCvWecHPKifv49YP0zMoeKEcXGH541T1mb0l7HIPwfTGKoXdDh/l/a0ht+
1ovgT2v58KPll0lNTIgGgQdzbXJ2WlHabtbHy13VGD7CmZDcHjEZKTVthOjb
XQ6jgDXGnGBzVYzyyXbusf+Qp/rJbtlxYRihjwZ9TpfnI1RLNFUbqJl8Em4c
VMo9aw9go2gCqBt918g3pUMbFvnSIcJqOFyT/y1X1RTVjZfYyntuIjcVkXkw
ioD6RMy47S+zc+PypfskUtVdCcPT4pjogjH2E7RiNo1nTB9C3OhDckRq4pu7
gsUoQ8I+UgC625U2KBT8PBPnDk6soYvDwOfefv8qB+17dXu0zHTtSYR/xCrm
ewGWP9qoKRQ5JVnn1Jof6P6Sf4lQn/LIbsZnOI+FNfNDya2OOka3GkiyeNN4
jziOyGnxctYKFA3dBM6KgpwWgXLMhER6p6clDybIAE+EGSrZhzv6Vyaiffoj
7iDNijJVootn0AdxUp3Xxi+FkmT8/L4hr4kmKYwrwFh0MnoAR5RaosLMqn/d
qOR9H+TfFN4ep8574iipGk6Q0lSK2mH8CSBP25ZePmjPy4pNhayki70czRmH
9V455jwXk7FNNYYnrALkpOYgD+08udPlpGhZk9JfuYG9fdaGdSAxSvJDmoUi
1k8WciiQnCkvf/CQgkHJV5lN6U1XJLLWgmJL2S+DvpshDyR+X8+lvBWNG6df
W+kECsSi4+XSXRfWzAkPoyVj3TAkq0KG6if/fm6SOfuJVFxc59bviaFCAjPa
Za7TPWafU43m0UV3Lo32yVY273W1a8sW+Mji3UVSoWlq1JyBO+KQ8hY+odaB
6j7AmMNUdLoB33NQ0AfPW+qM/kKCXBPM4LVIwantmBjBec39v5IZPWl2g9jX
l52oLU1oaBgawlTlbNGiWN7V/rI14QD7nuYlasqBDFcI3Yn51T9DtoSm80Hw
iaXAlbQGgF3ItSdPcekIBTeZ3wY1WV5FyBk+ugalg1GPN201QHnO8AoCyov9
V5Csd7RRZKpnXnFurXdbNUfvr9EEer7GzFGHD/oPSLwHLyV55VSLqgM99Y8p
n0mb0ax+sCO4CzNcLSJsPpHiKjMKksJ/pM9vfmFzGQp4NBcQa2koEFGEYKjw
VdrvjHYUtuC26zZPfiRRib3+T2zXAiGnH3KOixWNrNTrx82R8lo4mdbMRPE9
AprsBOGfL+snqwuqanK24ostlBkCvr0nHgiExndtl8AV/NvDUqd0x+zoSVid
Gvk8JHuU1ozyX/ejJ4n/APSU+OBLud28GlcExJz0oSoxv+juQh7dwghtCsPh
SghnAzfGa0gaTxjtaKVbnl/SIf+in+VqtIWbrzFlBhyV5CHXAhLzTiuKDbKy
FS8/GPM1w3Hu8FBJkYj5UoahqE9mw1At+fTbGFajdTgV7y/YPgS3bvpWSL67
aPngx8uv7G794bNHfUoywq35VyVScZRNQVKNCljpY5/BmhRhU6vYREoaqxS9
He7z536lTHOxyI2kQHEqoxigHxVDpi7U0D1do6ljdu1Ig9D/HINConUCuA7s
vNOZizGwffYYDhTbNTUTFsTMJc/zWbGDsIK8/QtEDlTtRC598A6CyXaSVwaP
sGkYdeuQ7iFhdshb56CEqvuA2s+RbOc0zYtLK9lNxOsNSolFIp88EcpJnfDy
VDdayxFvky3JPv6Bqk+PJ62YOu23TVu5TA5+bwSo77MOrUCRBDF0MRMInCNM
fhGBPW3x5O444vI8KLyoJnHVyLXOIuoeBJh2630ybJEwEWfoVXCGBwSYQR9K
+ljbWushp845W0fos2HCJhPcRQdZkQlua/2IRQjrNckRHasFB8nZkl594zkq
4npv/ADbnJOm4woXgj9edXm0UDPfH7UUz/FfETXHzsrUU2SyR8Rk30Dx2xON
6nxXHSRGokmwM7i1SfN1n4HIQ2VV8tRigPCWAoIC5VuvaSsn3LwXot8QXhqV
bmGJZx5NIAbJNjkgXCrmwZCTqXETWC610gEyGUW24K6NwBIMgo0o8LjDzZ9h
SrrViribwE/K8bt7IB5ywSvftk33YGkf1TJJZlCnFuL9OsrTW84cNNfTKqdj
ngJ7GgkBVHEELy8W9q8AK8AQfEPmx493YQy8ZK1Qkla7OHEogFTcUVfazIjX
aa2rIgwbyOBQjmufako43fobYBu0OgmeoCC/nOx3Vi/htaYhIbQYq8VAZUap
zz4Zdcl0cCA0bLvDhdczsD54Lys7DQuxWZxONIjeq2UDYNlJqA5G54lGpWEG
Z4oEVd5YmslvUeZE0m0qYgGLnLDxYAMolK1sgL9mRde0QSzdofD7eYZRgtpn
Zjx+8byUdgISVqYlM1q3anKZIC6dBvRq7v2P8pRYvHOUtKBrJ4TP4+Axfrmv
93Pn9DMpQ+z+ZtDdpQ6MskXQzLqrOO0e/vRPRz4B1v+DVndQPzC4+zSjLpqT
349vW9QpGzzHNvCvqfU1EL+KfFd0u67gBIo6UYhILkwVng2jUxU43YKrp8BA
Ke0Phq7cF1PAB9mok54/IVxoMITEX7XVKtC6SOrKhKprnKlzgs+YMQVe1CAY
FxQW196ncKwf4GMzZ6LIBYviJUbTcYWgYsBVQf7XzJcobGb9Qthn0OgWjbkj
F0kbtAOfv1BgTQ8wevWB1oKNFrSRKBXgRycPb+JhAvlIqf7VBAmhs0l9c39D
7NxtaE3QG8cCRxK+3RiQHN8BmkQBLwnDGH8ZXkE2tqLp8dx/KeQd48lAC9es
AJUgnT8bJDOAurQxLlWvZ02pDlYjXHQ1YFPw38FjNMV5FIDwlNOOQAH+EQIw
AwzPkbUdicOYIpMVqzi47xmaXCPWwnxwz6eDvpHvY9nuFjbF/+OoiNWsIESJ
Sk2vTDDutYTHDIY035vYDOk+XLp5M0N8g/6wJfNZbSxkFWGv/4EV3ljoUoiY
vUTdagLwjMFg3oVMY4cCAzrA4taFC7wgB5Pv3u0cwbQfFII7c2UXwX+ylzDC
3b8g+CtD67SLkHO30xnoQbQJ7Fk2v1Iy4cwPe5NCONwooOigOAJfxPsTixF3
uI+iqOv2/aw9TPPBUU3DVc0llCWP7JAxW0vIpfrIbppw6qr566tnEP+Xb21y
aL5U4zby2WL+hBGzxRFKgmVJFnJAYgFP33kHm4zHyOuFhbEeHF1rnSK7Slwq
03SwbJzWoXLX0tTLJstyt7H+SOKesoXgWT2AuxBdjBlPbDvXQBJMhwVXgU53
vEW/q/iE8woAGFHVx9aUQKboPXds3dhnCgsmMdWrKAZPNqiLe3dg7f6iDJXX
/sBrrWJvC13kesryXWWhHZMuisI9k+4vXciqNV5cAQC/i2jiYkMfeldlpxSO
loUJCKvT9q5pbO71GHvZwqtPfBnJ9siZ8rezwe/jRyQQeFZKQp00gKnr/tDR
eWoXn3IfGLZqyPGr8DyYFhk9xjrTmWl+MqTEfNBnA1xbSZg0nMQJa7TVIwV7
pKBfT0FaxWwlXO4ffoNgn3TSCi+HsC1FD162AcVYLbQxe5SfCiJjUL73ngrn
Er0HSvqatphxNUlwndf4qslogKw3MrNS+DVYQkFKfFKxKRnPx1LTsEL48/w3
+yHMdOetsueJTKphJe+xxNTW/MI+h6nYgPxXPsiGi/HE+HGkapxanY06OYLP
h08MEOm8THSz0hZQyYtyVjV1FcAoNW1QsJmZkUF5WnbyiDYQ72NBrMS/4mft
qpmL70Rf6gMS/32urQvO49BV6s0oJb3tasKPWy7gkCsnhxEPZvjFMAKHAJIj
c+ZVGmbqoddtklKWxovNrDD6jszGM7ZbSutHTDzsvMw/lpsRfBIhGdRbTt0m
N+kfFQGivSqjvK4OEyXlb0/ngMRzoJ5kd+9CQulrojnc9P0RyUEktIXSg7SZ
6ivd+CJmNfkCaqIZGLFsCGDQLTTIRWGa/j9HJZ77wnVEkV59ciqvbjlwtqOq
GiUUlapGUsXZLlC6++i8oe5u3bJsoo0GhQNnnUsPuEhHuG4QbdxHxd1BF6X6
9V6f1+3yEAoBJa9E3vcllfTqz6N8SzfLO0038id64B8GQb7X74GY7j4wXOad
CoGwTHI+dNd6prXfCzaUzKOfg6zyrenq2DHuT6sGT977awuUqcjlsA2rr20g
UCAk7KIMrTxTee21e7VPwZbBUIaz3j+AaQteU2UZ9wzzIgCzPxb2ovQmuLrM
6dp/Knu7iNWmduuTRyaHSNMX8PJh7cONiePq+13Vpl9xUK542OuJDUMpyYBi
rlBHbSJ32Ljx23uodPXvXb8fkqVbEZ040j92nXcl/FpBy6gSmS61iJSJD6tR
uBip8vLOXRw8y5skE1OZotg/ls4qmrbDnD3HvjOlZwpUYfcB/BO3gpBjrKMo
ftyQOtX0pYagTurLaCVINYbkvETuyUSOIAj47079H7b3dOnHk7PqmsV/vdq7
HQ0zmbkF8Y3Z2MFGa4Dq3JHfJa/nR9IAWvgO/GNEZSqsexTyUIiX1KSuZC9D
maWkDRIAUC/ogX2VSsYBp8nN9fKdJ4ITEkrGLrQwUSUCInjoIxe6HzLICyv0
V2sdL7JFsWPadSBEbl28h77OyTJRU9EtumJALtwMVO15pN+dEphgyCMT3ykB
+NlFbJ5whcBbZljkgfNuqSqYBW3SUXeRfuJRT9lfDAlwnF6Vmfr+/XGvq05l
dBCCk8aNAmnowuMB2BmzYYo3fwh1xkTS1n1qXhWZ/8HcMqs2uacAi8PgU9Cv
/hQk/9jJIKxDWaK//G1fLgE3I0UXbTZBTPvOBEgAc3aKEs2R3Cs1aLhXbw+X
QcNkZuvg3PeYy3SM+mnIjbYtDl4ZKdHeQ6OOhwL3iZTWbWmSYLBHjQlITJ9s
aGWKU207gBD0Z1bap9+4FLxRZwQAN0JHSWf24OeMiGBxaocP8qS3VfnzHX0g
15IlVuZymHNFgwNUOAF1p6lHrlHQzXQ6zPTWI6SKBmDzdMIlDSurcX5nkKAH
gjRhtQ8I7X9+Nhg7lhHhFKTR3uTt95RQy1jyzVy5Il6GS5IjqA6pYIQAWfFh
bL9VhStt9gtCQWl2gqfIUInk+PiOt/uDhRKqe9U8w8Dh9XTdQMiVLYv1TBME
CA7z0q0DVk/jwp1Fbq+f1fZKkALPy06CcH/YSY9InmgTLJX/Xm8F/3z2tdN0
1DPN5XKqlShEFFOf1gD/U2QfkZsmuN4thxI4A06PtWVXQ60SgfHpLF1O4ka0
0HS9xJDeZqH/pielUPc4mF54XpFAOHRgW/Fs4VUiE/qsamMccx4t+m4YjYV3
sKQ4PEx/5ECz6HTtHK9JAwrf9fTucKTKrKsP4TIY4Q97cNxVVXhZUq93HATO
te3WWm4rjsY3sy6SQefZbYKb6Il6D3zjW+f/CTmgJseJ54wKJaJdRuDbdCwn
zKGnOborlAU1CIUt421dUipDjdtQuVkYTBuBFBzq9KV1sYC7kyt2d+9T1zZI
/N2reAIPRk8ItXXgJgGXLG7XiQhnbII4vMI5bO1JZ0m9DPCnoIYqmoB/1VZI
zCNBR8X9GaG8VonI+Rh7HTGhYSGemZw0AW2CeNUyrKuiOXO5b1q8b0E3xoyW
Z8E9E4eU/ZIyPcqAFmHgyv5PSY0YVOyFNesEXu82RSME4lGDhjCMo0wMHCxq
ShUM4f2sb1c3AnOaFLr0XilIlHbKnSOqy52aDiNWnA6dItS9XHzKEknfY+2G
513ILIbT96iLpvD4zpkKzBvdTgnNQ8eG1aCp7xxa2/Y97qBFh9xMSrX2/Wdt
FPbNixd5OHVZKRlgpq67XMqRGsQxy9HoSqRS86U9zdFO3Oju68RZbcTN++LB
3vyQtUCyCC7+LQjzkib7bT6SMeGyrGf9bS5+VY9BVj2VDKtc2TIBSSE614pk
pwhcckW2RRm2cirESsChvmWxbePR1ZQqiR6GjFYUop+cWGZWeeNkLssgnwL/
zvzfoVYTKlG+ReftpXE4cx8EXUi5RTI8CYNB17bN6sHWgBlKErBNhB7gCN68
nQJGvBnihCFyT0hfzlZ4GngLAljQFx1uNjUZIhw0hJveeOl5e4K3KDG+1yeQ
RnUxzAFHPIx5WvHKb2CCTFWax14nO0vxARRPJJLAnDcgY0+f4EuuK/VTro9J
iy/1a0CLSCPx3qDFYq96HLFk9GGmjMldqF78Xs78yvFjH4aw2db639n9zMiH
w3ovqSq+8KeSVRc7Tkyl+yEZip5Jtc+NAHcXtul2owgaAdB+Gnr73gnYc2Qj
EeYTr67DbEUAL7NjrP6BOlkmbxvj+4vEcEx/WkpVpE5HKfEnf/vU3sqtsF6l
vLI/WbW/HYzpQJI5u8Xxb1l66b7fQwiTU+imXzzPtLoI6dnOvSwkxRuCUzfs
YcpXsnGCQ7NKJTR2IUG9LbEvTvs5dzIG2eyNZtj292wnWzAjYmNM8TOTwTIa
cqro2MQBVhqs+elmp5neqL+Y8iUmDvUucZKB/IG66tqJCSjUbtak2V5peqA3
CsO3qiS8T+wwtSdz1XP5jI43MZ/eOjev35q7ZnXBhTIrWqSqRCIi1n+ptKwi
f8WQVZ0XSJKj5EYeXGBmOF4EnoJE4/zemazBqOcQ2qocAxFZo/U9HwAlp2kB
fvxowNpBcZ7xlNTyCuvJXS2GpqgjLmatq/ALbM06N3HEsclN1jYjCUwkm05P
yMXQwcgYpDLkBoK1DweVXn033x4+aBz4UHutcXBR8I8aqMcWuoPbEd4Rd5RF
klVFNPnpXnIKTZNWD0FUKD++JvKclP+drp+r9goQw95EOhoJzXYM8uNGG5B8
yrE9Qi5Yb+QrDboroG0l9NQcEfZWM48sQ4ZNpP6Dpm/wELRHkWOazc5zdpmX
DFPaqe8h4tfH4XEaHGmAxTsAH9loSX5BfA8kjEsiyDynb07GMG0KpHsB0hbM
q0DESLGo+J0x4cHQUVBp/mO1bSnOZVFngDUg8wNxoMtIctFqN/2BOCAudlnq
NazuHJ2+LB2VHV6elxkxbn2iIGZ6hrZgTdvKDdI5pvEeOu2mfp+wvfwEkLow
3Kfq6UPXq0IslbfyVZcpm+P2fpr2TFwt9k7/R3xzmtuif47Rrd1WLMM1yyQ0
6uNc0zAP7OV93XoRLlW2SxW99ODkJVbUMbyYT3ob7/71TUL0zu82FL/HXlO5
bjTggJ5YAXKo7PClwxZwUZ04jRvxrOKHwRHal6wQhRaamPlO52bSmugMmpr/
/uP4fJ+b5zfFHO+L6Fzzyq0ymiTfybvGDP6FnLhw4mAQ1r4xMGPpT3+a/oHs
Y8dw7fYnGllMcC3p98E9aWkAaPrDuFYUxm0dGvRVTl/GZydIs3prFweNvtqi
8DvHNPNQ9MpiwsvOywqzBbpdcCHGXRXkCdH8qGSt0lMRP55zjgZW+sOluJvU
nFLBUN1/S6D3K30U74RuJjGBpnjcS1BUdOADyC1XgwJlLLoKEaBKCYjvgvnA
ZfU1vgdsRuqbD6ht5KY9Yx/wLnZkul5/tTWs0e5k5Gl1YAcrCPywsLFkDJVU
nsKKaweIbVvYvd4gtI7e0AODxqRv4Z0zqvdSzZCVivEqsiInpw486IzqMp1t
b2FsWR39cu2uO1t53cbxZTKO5TW9v4plbCnZ1guUasJYutgynm2qdVPnTqzb
qe6TYzVJmJ444zyWAK1IX7ZNA8eFvq4Et4k4WQ/xK3f+uO1hr9xgYufQr52e
GiZGwziw6JwrnVKfQUqhh/u/esIxKMk8WDurXJEQ565pMfgQ55QOvIbzwB1j
Axn8I5NnLEHY1s6X2ZGGw+6WcjwdSDLiDtN3xphITvP6afR27HNdazq6NVBb
ONeLco9u4lRP/k2h+r8x/b6ea8iic7Zed/YmJ1wd4i6ii4V6bGyHwgq74M9U
5MYjYBRsNY66+erh5AYbjX/gxLMD5TO3T6h7niYay0v8PS5WMcctH8xSCO9L
9DtT/eeP450vd6eEAwwqUryXz/l6z4k0a3UJXnb5HSb6io/wljbL9NWB/fCL
7Nw7mPjgJDE6abVqYvMpBrNFvflaixm70W70vO9L+uTGYnbPM27Ce6K/2Pl1
rpkVYo0V+snr9DMN4LxPq30o8gr8leugh+cNjtIO95OjVe/rKIUnLrR+dqWJ
Y/GFwt5vHibblZ9Jh3de/Xu/Clq1guMTz7f6n2232XNmsOvOZeRw4aQIGOz8
P+YC94q3goBGBGHb196PskF46Odw03/G4yI3yaLAaThB/Ct2fih8jQ1D4H6w
lEVMgFVOldFbGI/D8x51H3CT7rbnC3JdqDceoWQLq/t1lnkxz3K8qAkhe5ZC
wSgDk4l7h4qi6QDo8XPGqs3mI/6zKlf9RaBDOrTwCzGc3hLV3plxtwmz6O0g
jt3LJ2UsZgE4yTAkkKmmHi6ODRXsLy2gqU5Zn9//l1B9ywSHuYZbXDGByzre
LQg6+JoTR2z29Ga5yr0dqShhPjF2u19+pS1kuDTdTRcQ2+brqrxYeytvexHG
f7MtWaKa3CzxAGhU7hx/0sJn2/MFUwPDgQNlUV0qUZtNyBcuyU+PZVZYVqa+
XlH/WO8P4BosyedTT5HagUp3iN7JYAuOHXddDhnlpAnvSk7t3p/ujKndp7Ua
5dBcNclTxmFQsrpTXzFmapnPKe0+K0pmYBT6y1mbbqC0dHEK4thOvHMOI4Tj
RLYsLMbScNO7APZ1RjP0q5xQXGcAwTb4LX6ycuBoBg4Tk4CUxs4/rKQ3nIcy
dwe4O3jfaJmF6jhYTZGdwHB1hoQtbWjQA19bn+i7ahko7UHbBpaP9SeCTGxI
pQFChUiXm+U1a4vbCEoDlteoGQr0AFUjoucqsuX7qj4F3K+BxB6BUWIYyM7r
PAKFj1KOmj41/zNKGzEnB5H/iyJ4OmlJvcadxfte5c4x3kDPDhuVHHzFf+bi
Duf1AgWJtyq40lBnNCW5+MUbcvSVCDzRGFrvzjHOtCv9PXnxzKq0f6syH6DC
32E9CQm28DMFhzXbgCbyGz3ckO4QxuYPMSeKsqw+0kZrSA+/SrwY0PaC7lxA
JhPNsZZGQ7kQQcS8PRcPuBL4buf2KJ0U93IEpRf7tIRKHEljm2S8tmYGS9Jf
kwWFf1hMSXT97kvQWOw0cDYvdY2vwzmXtG3PrNzapozITYopHTJ6ggDXwWI/
ZC7vIh3HfSYTp0HfRisIXjCFBe3uWI1+OJOJtMtfdRfkImZIobjHbExLzgrW
o8YdbMbSwNZShnSqZ5wNx06ioY4+kilCx3DDJY3qNHRkFqcYWM8mBXwQamRu
TetkEF6xYW7ej9OKVEN3Xmrh3zwexoxhQ7Sx+u+pm9qJp44hoHra9cJOZtgd
SzgFtz1QRUg7KUVCgoMB/pEjJlZ9JsiQsQT3Ix7ULpNGTk1E90SFUS2X4gLv
BwXU4CDSZE5gTe9k6HKQx61g6oCHilAwoPVOob1tji/w+e5n1h9OY8mueI1/
98EdQ6bLVeWb/tW9skr7Qx7auDdRTngZHPquDRumnqSgzazMZ3OrlTX78vl4
23MO2nAHAZhza8WsgtiyWfcXbuGRW8AVPd5+3mmM1QM47qKekRCduN8/ZuwW
yQ2Av4yU7M2iRVZ7UC1TTx+Ig5luUO5tPKYBqJ0QnfP9cPsdZtoJeUo0F7Kt
m4Waq19OQ25Clkv5DtamNDk5XiaqbaOTMVEULZX8/aeSxThoWaZ6vaE7Ddcn
IPgRNhSrIX1jtrKjkGJhdCKfQLUxvM7cpapBnuTN1lyxBKfaZn502CrqvMg4
k6xQjnGLZOptpJWTbhQMFmcHTAYvk+8xqJ9t0koxrxJtqWIUeeL8sxKPXb8y
Wa5vSPdkGz1R3ZW6Mf6bZiV8av7kFi3RC9pZ5UWDU4NbkxZvDQEIaYDC9S27
yNR6HM/1rkI0uilDiLKilvU6kiIgOqbxj+5u+FysG1pwxb77c0m/CBp5hEKF
pA8TY1kFPYOlFUX2f/FK5KHq0RA+6CmBx8hOY4POb4H6Io6s1GoxuexCrHGm
0G6y2CE5PwLmVVQenCdHKHlVn3qyeVSE8FvSgdPzazRl3Kg1mCcSA+v7LRx6
KxEOokZhauej4YsSHXZy25HCQ18TosXaVQGf89eSPkpaia7Qz419PvV+6CJG
+jeyF67WXbruL8Oi0gW+HyNZFs2srkrAZGKUzpeCCFMSthqyiuRbO1NCSxGu
aXbdGYpvugJ1ZExVx6lyEQbVpwP1XD1wii5ohQS5AQ0RtYBneRClQpimyLcX
+jrozKAIfk4U8xdNQ89VhPje4bo9Hoo0TAR3O+KiRRliKElUWgQcJ6YeLCtQ
z0hoSzjZWO7EzPYZR+MRRJ10VCj45NvqfUQg6ncyBSY+kKckXfw14V223OEf
jzk/KNF92nT27WcSVSAR7na02Lt7df+yGYR3jp6Sp+v8vhFCtNe571C65vU6
mRdVdFJIWYw+ZdPE2FYo3Bm2MLwa7Smls0v1m1Mr7uu0PehUTSMm/TtEsEz4
7OlPGiYANqp7bhu66Y7PB4yuYlNwUoCorCaIqY6FkOUZumb+NWtrFAXrS1P3
w2JpKWv1bzSEsfjVs45+wqX70shQnjqfGEQjRai0XHe98Af6E/zw5lerlgbT
GbYTVaYaXuUukYHC7F6RhANnkB6uLM/5rikq3PqMY9BpRW1/TK4ldXnnw3ai
39yg9gNI3H665H5QbkN3AKhbEIG8B5CpZ1fBYPDu4ZDQBOn0hXlzqjS6/93W
ulYOanBzDOe8/1gSwG+vjJNU1Ko38eyTa3DK1FrTBPf8uzG6ePmtUh4eOiGR
U5MUTOJ991peYI6b7uzWham4YW92R/qib0zLOH60g04eY02qPWH+bFnLt7+6
3pJlBfi3Isu8LijrJs+r1dRygDbiqvAUsUlvN87b5A5cLWmdOPJsJVP+47g6
kuwfcFBovtwqG8ezPFXs0tn0aNIBrAM5z9EJGC0i/k4lH5LRX3+OyY9z11Hm
NxKTEjkr/w2iZu1qeT8RN7Zpq4OcHkz3pSL2DDhDuGdkL44WExRu86F6Ydbi
r0Ir+9gQX0XUug1I7gbvv2M6Kuf8MTrjfZ2fBTEuSH5OBu3Qknl+ZMqzQ1iQ
kDyUBf7lBsxY8HUoGL8fakKLqxvJNwaceK7inY6URxIXTZHQnpy0/O+OL97j
miZ7opDtgx9X1F109eLuTiHJwC8gnGTVyCqz3MelFR5L71OnnNgberS6w6bx
IMXMAW7HiS8lyoswE2aXeSrV6xTUbnkBEfuI2vFsaQLG9iG6cC3SXpYIgyeq
M9JXtqtA2/e8lNFDGahAgo4PocsOwXvSk3/NDgE9wwj2TR9TDEj9w7QL3BIO
jVRI0FBrieuv4r4PnPs4AQ/bbQ0m3IkcIZ+Ci/zfZ2W6zbjAIqy+VgcDaN4o
TuihYIPNDY9ixcJcFAKlWZtsWcv70oFbXfeiK9ZlwQ2xmzYNheafXxsrGXwR
Js0v1vbNh+Z9EJSqN8TdBwD+ZqVOx/tjAJUZZ0bkR2j/patIWFN+Te6lL9wZ
Cg0nA16ffRmlNezzIgkmBqyJoX0vIFKdBlTFazVvo9aIUOjOyjSEq4sjfjQc
I0tNJOSYrjgK6EijOtXmnuGCFQiOLPURDD1sOMN23oL7kUR37fpTm3lm84+C
R6kuYTkO2GS/3cQURFSS1pb9cvUBv/9D+yheAILgBVcLdiG7jR7Sf3H39iic
5mjtzZQZBhAT7mSafNnct4JawtVzzb090PJ+EH1I1+OoPlnCs3it2mjTgQ6v
mq7g5Xv325yEFA0CGndrwLsm+3VhjMmQRD96HJWiidIrMgNNypwBGZJae73N
cWoatBdEMttwBihs3nhlqiYFU6awxO/L828DFSPnZqDLxy4MbqnolGNh2fNZ
T9LoF/3ehPVo+NFvtCKmXoVWmqRgxS7wqViUQSoNXjUgRduZ5FYoVJ591vkf
oS1dRW4umpVC+gs1S1BhI4RTPjBFiRyIppBxAFrHPoQ2NqAAYYUBmviUM3WW
zhgsI6Bntw3ps9FFNJisUYOuWner9tiMjc+3HQpL4ffgdLx5D53Kt84zwEsl
Sius1pD1nZvgLbDHGralv40/9xbf54P/dlbAySXOOITfgbXL7k6ZuDVU2FGQ
Rq80yN+iXJJUqlDi8KstId6M042NfrcLcTpnqdFvh9ZczAbqYBoOLUUQLB95
LsLzS3hQXROcqo9665Pol3Tv5zcp2zLHGxMu+KCKIt8eGxVEyEnStnd/cFRT
iucViKe9NLHIOrtoSPgND83J/M4IFj7jxqLNIn6FiO/2/mTRRwjKhATpJLBf
JJCVp8huPPVaoX2hqLcOZzVMkpoZgQaAXjA/GSq54leZD2rTcs0UNxYUdIKx
AvBtIwOcBTeUj+2HTUFh4W+wBnCSLnFDhxhEYEmkBH9Ar8eT8PrJHNZp61xv
93FyYmBc+6L942/AuCIp9p0C5xLyhDWrMN6g3AFonsjMOSV3Vds36S+JzAwK
MbnX+lg1jD9Nvm5aAY81gcrFYtWMSza3lBGnm8wavNWZj5YeBphqrXO/XaF1
wKfUqPNQJgiPKwXgFDPhe7pzA6C78Mj8oExo4kq1+aJmBgYmTJ9T2+c55Dsr
R1wH6D9njTD2ZP37Hpg/jDHqmNntuMw5UVeoNTKoWR1sfDgYNZOQ477xeyTB
QHxiwmFwEua5piTgml3jwU6bbtBluxWVbYT9qKqxd98y8+yuWAs8a+PCr5P+
6O1AaPtV3yNEh9zurHjggBuMd9ChIRMDFSyPrN52q9gvRjbBaZTk7QjXK1Gw
XlCRc4qphwU7quhecS/QsNtr26wZFLuFSrw5N+tnM8OMNg7IfmPp4j60s1Bl
6M8F8B6M3lqNUcpAbSEqVNxxHKtxZ83mwOvdAnrqxj91HjrM6f9WK4B+6jLf
oDEFZkzM7ipPh4Fl3MDK6sHI89H0qO0Gu+m81OtxBAFtIpZL0kbQ22t7wWlt
2lfKHcCYDCw+CtuyzbaA7XWNuaRd7z7AZQ2GS5nphsAasy2XocikfveySzrR
0RizlrGKBwHVzlpWgOhEHiQiisfP85vKCJ4r/52hFqtfT0loA4g3Dp7GuL/h
vul9AElkzl7ZXNWZ0g8aE6drO4uB5shSG/3ql8zZBc06YzadKlFz2ipsk3BW
va0OZpYWx47oC7HjfZPvg3l6QkDcApW9vgCQabsP4VSwx1aAjtPqRxxtjQMd
/fanrVBRZsRR8Uk3rG6xWvji+1orVJbFCIRRxEs37hNN49bfWheXH5II77R8
E9kj9G2mVzwv1eJCsx5W2REw7rHEcJnkvLlSiDM2yFfyq1gonGgdfSZikNss
D7rP1yKCEEKORl2suKzUd1XVNvqxN71eEVqPhJcBpxPXIrhTCpgJ8R/d2fSz
2FkFkoHfEJ54NXuXpYlbbty8Ph4lIcavJDotu7C973FNa5M0lGg69mkxaO3y
ubKxVErG8dmq5J385/VjLC03QKvIGaz9L0vfVCNUhVYl7uQKv8Ow90eAOcYx
ZcS1j+ylHYQ5+nRjy2swPEi2nP+oAsbW19k+iVB9oTGXgy+ctrCowz6F/gdQ
hvM9ArF98OVNaXWqtiQin2kP7SjljADLmDykP8bjQ3I2JzgrT59F4ixqUFm8
srMJCg8zwfR68PuABYLm7bZNS8zoSS4ZRZo5b2ohS4LHb3M+Ey7tSXml8Uw4
rTpizsuzruSNpbZg+xct3Cv5gMu/EVMysNC1lsZAN2fSUmhBduMEkyrHukFi
oVRGtP4RVKbqjFEOSGoVE2cpEtWpnXrklPArMG/BdBvZLHjqQG5pTb/mLRxM
TFbmstGeJB/8zLeMe9U/0ltKa6w0/aOYHu7BkDlVU4uBQ4my0OxDULNokXjq
an/rf0u1tANvXPsWyzVYjaDqP/h2ENzawAXNAbcSTSnwiQDUfu6TpcaARUIu
wwMebCSovIJz04DowIByLSN0+4mTG6q09Cv7wI3qWnljCy3BxjE5LZtF1aVq
l9ZvRUYB1zdJuFP0bhmc+O1COu64p5wM7g3DhyJe6OxXR3H3DgFIsRAWxgtl
aIHyciH1+v4hNaExHA7NlHRc+HzeiPeq6uWnwctsoQ2GxQHckdX0WbCjQkYz
a9IRZYzK9dYq0sx0l9Nnj2WgBi3U2sz4FiZG4fkvBED5UgIOwB33Xnn794mb
falZlY0vKjCQ6hrmayRZ3NqQLnOheJLut3k5WyV6K+S5Yqcc2KcXzrzujPri
1AEzmUXuIv3TmBNIWjzAw6klD+De+z7PC9Quype9bmU/dhRwubZ3NRN/xyWz
TVpW4kK0mhnpgCDPAhzSGdwmRsjMEJrz6/Mv9uCmPcSdCDsVMHxXBeOWrxgy
HWnDDvn3i/xn/0VkAP30bnKnbsUMnDeH76HFUYPTrDhMaq6Mz+R8TYdTsYGP
8RsOlN6Xo6CUWN7vwfpJ+d4jh15V/6otvUhpyTIsyhWdCVGa2WlL5coUfzse
LHvPIdrkcZgPJP0xucO/WxnsveAN6hV1LEP2BhptCd0sHX+wDsdO8zIWb/qU
T2HjdgNQXRSGG1DLznzkYZS4h5EXQklTkHpjKFcscC+Hak6iGC4OJ/3Er7F9
GH130nR2QGlrZ/z4XViNUXsouRKHbJTMFso03PPyYG7tbrk5HT/Ccmol/UJ0
y9+A1Bhvf04cTPFTQhgT+OEh16xqUt+6Vtxukron1t6mFwMrLJVgz/Cj/93o
r+4UY26EjDiYBJo9GT0PlM46b0w/Yq2XaH+aVPTmTcKLhaOwOz9wP1bVrH7V
Bz5SSvBt4hv3zb83tOn+z6J7X8SjSF5tDMejoPzhSjRgfmC+b2wDgrluZsoR
5oJQxWp6TMkwUzpTTmFzPvPkQiCK6GeSUlPDo7L/fdAEUtO+fWtikXXYpzxI
RQeJDO1E8IaU4/ezRVg0kt4dLMim8WIxZCDWQQ/tvNjOlPDdurOhM2x7fuS4
eYQY9U/adfGDm508PJcsiq4Z6zUYOIAU1ELBSJnYV/R6hn7r0EM1sAP70x6g
5T20ABbRK6z2Gq8ShoP8G7LuBA0+5pN2gOIbxZwMi0etPCuNkCD3QwThQ5vI
hmmbkq+HntyOzf/a3RurvvV3iZqbBzknelSe6LHf1T+QEHgMbxyinq7xkQLG
VUeG6AFIm661taFCr2B6J+V7CyWRATwQMwWaml19tfZ/SYF4oYE7X0skvIG7
YgkY4qV93T37nI6QtswT7RKAo6NoGTaQhewE3RJsfTVtrqhuJxl5cQGVBtRs
26jBsg6kYhMLjfVeIVPUSIUvO5yioeSZkqABgush2KXEO5gicMzaOyOGbNtT
XbB6sbGs/4qAg3GvDMYTqye+/w04ENsr4ERW/tfoKHyGF+Y2a/zEx6/PZbO6
YT3hE6qFPPZq9dnoiY7GE8EfKj07tw2RcXzeIVvZJsP6FRyM4pARRP2afLyc
QT3tPbnoVUmXLnBvNVxPVMBWUx2Zm6rADKgccHpuGXFQlTWe8iq64kYCNgmZ
4L685rkmy2mkGChPmtDx2GSZ2iYH3smmpEi9kHJ/1ee9hwq7vbLdz75b90fb
Q2YsbEmdw5FynQg6nmZ94AsTK7N6ghLgVHwUD4qBIwgPpA7yEpOIoTnqH4VE
ceNSZmQ+crLhtEHBdT3UWZhkaD7LzDK5ORrW1f/OIWDKgGynh822x7I7Jl8u
KdslhtwMxKCbkxA6KsRsuvED5p1o2lYkCp5c3Z57c6QlK0xUTQigLk7xkmwZ
/d/SXolIsqf5NNwRoUDUNSx8C+sXVEIVfp8o77RUhVTg6cUswbXSrYRHqD1R
EP32FZUQNUkNy0gK8C/ceRLuvwfR5nwPV/PAuJYm/VT2sYhDidQmPH1zXFdm
72qKp/H71CUfFOnqZxXdMqS8PwdWIpqB38Xf3/lNbs5eNtHX3Kkxjt4lWVFN
SyZluaBU16H251mRQbLaMOp9qfZdtvmCW5VnMCDNLVS25o7SRCvfeBJ3kLbJ
eDNxCeNuD6sW/dndrskF1ftMnl/V5owo05OYdNYwOt+qYa8EuFSETJUmgvJl
dzE9bQUgPxTKv5y1QCkvFgDzy8PoOynKhcHHJkZYOUUUKR8/UH6e23/AzBvV
Ah5VT+q+7FdBBPciyrciHDw3oyI9ddWfHI4XiU+RhyURjwk9MIe7c9yATmeh
u5kjOh/YJHqtbyx5gch1+yRLXAFWJYi25iJlGlOkuMT66nsMISccvZ6PULRi
4+X96a9iFucNZik5/HKtCdpbi1X0wbQLgD/iB2aUFwTO25hXG96ZE++EAuQf
Cm21AJlntjCso5CEGCBxqNYDdika3PioShOeU6jzRBUtetTH6zAX1B66AE7O
yp031mUd3prYQIyKf07Ex8LmrLTqOe/oHMKQYHZbbOJ1BEWJFSXhvO0vicC8
WUivmg5jxPvSo32a9LIBzHsujkq1oKyDOoGzcbWD+xsc0vBW5rrCo1MUqi2w
rT8ecqTNOZ6DoxH1SRqvcaFY/ExG5GrHS4/u3XCpXYOLK6R5n8+fQ2hN3JjD
27dgLQA3T960Ezw7ipK6+g4Xn8JFjkDxH6HDoFjiwk0rH6oWwFT+AfpUu2dB
glnNy1fYrYSmNm4S031xe3Es4DdspaPWxU0IievqRayNEczpCZxDUt4QO38M
ovzRkhquYnqN/CbnDWX+mQZw506Qbpm6mQ65xHttNbcUkvO5Y8FqjtK7fCr+
wlr5td0djaDucZojL+fL8VGRqQBxyuXlzE1FVRWhtroUZmi8i5p1KOSVVrDU
JJnfgdhHzUgoIS5bQgOAlUSGFVd91FxaB6A+X8Vm2d6c+c5+OQaoA8r1Ubbh
6pr7LZsIqB9KPGr397rYvZaHVxFyNrivQ8Uu8+qrz951jiDfmJaDYDSJVuit
iosoVD7zinx3NV0cy/SYk+DA+h6SVoamx9v8EOAtRXt5VrJbNK+fsz94FMlg
4F5C0dMo/zGbOR5yN/gm5q3opGoheuyebWdVzThlOpdUm6ZtIEQannmQ5L8o
6kM1biBV/fZf9HYKG9fhR0O7smJMu+f57oB+5sjazu8l8dyilsl7TPc8OISC
FM7wMC9haJazV9sK/fuQs0UZH0C7Ab/1D4EPYUu3nKcClA0BY20+oD0qzvbW
d4xdoFdPAAL+/e1xR47KP35F3+QZkNrQRICT+f1C1STpYMwIyicIwu9JpSNj
iOFPEDDDj4zF8SgCbZMDvmTnxu8wpFrjI82o9/K6EMUItyuXBG+WDyhH24TH
wyjKFhBgRQ7yDOFj/RE9tk8oclae+KrYqYwGvlqYWhsiiludVuwsTIlY9q/I
424FtC64UuAb/hP8jN46PncidOB98R22RTehG99wRij1ooIPm5LAZPNvn1sY
34buyMRs+Jvbzz6ABiHJQUTPkJeSga/JcLGDm93BVslVRHltNYRqc2I0R6MQ
T1nbugsxQ2idAugyeWbFQ1chFyblZlGwTgUOb+vDdDkjp5ah+VfBi7Sycrb5
MxibnAYi+RSFhaWanrX88bJPv5rEUMsN8RbTTxSbRHegRmWkznsotGtg/UUy
IdmukBEORdtopgzQzJItJJ8IV85+x0Ri8c/nfcC2nFHwMGQt77O3SWVDHch3
hMDHxa5R2SomhkZPl+UXvCjPvhbGjbwTqirCcOJUvDt/OCR0PeK8nEByvEZk
A3gqh+Tmf7osCwApcYb8U4xQbgbEg2Exye5dwYvEZKY6Jn6S/FOpp3T1isi6
vmmRa45zK+D2H7ce3qPG4dr7BfKPn3vesBPmWDlxg4tLy1QhFMUHaDtoVwQW
QCU0Wp/gu1v9ZsCMHZv+ThjfBpJZmuBSW7uzlglD5IhoWVyQznfLAiYzfTW8
Ds3MrjMRQHqB9y7UmdXFCqHsOwWotGhqjcrjmSf7aG2HCrLpUwEudrmn2Suj
Q1abg3MHiNagv0HT2QwoUaoA9PWOydWNrTQYatctSR4BhLBUZyK06SQGSwMd
hzVHiaItcMN8GF05l+pJV5ZcLm/xth9/J2FPpKjn0ur2UY3WRd/Ny8FtLqMn
Dz2CQ1vNRylNOJAf7FI2GBb4G5G50wwDe3IA5cUfRS25/86M/ZzK8oAT6I4w
sgzae0RCimfuM6fQWF4Vg/fWhK8yz2caK2+h/BAoDgA/SGdtG9y4alGXNjVM
SVsdJdwJSeYP2uremqy/f+f1HoRAK+GRH6yZQYgLlnwUlOh8rRefXb9nFUXY
cimh6DJmw/kBc0zrv1t6kGWzmjchUv5HtK+7K37t7mnWf5sMeEzpoQeiHw7p
eVIS1RPcy8oowPqGeVeQX2KcQdy1QpwMdUAIxStZzceey4LpNGV6pKNknaG3
ihEwT7hGqp/LYRm5CouOD5eW75lnKcRh2k5gMd4Zc+hCMe93BB46O3fQ37Xz
0e85/nV6gVRwy0T58H2XuxebZUis6M2v6o4vJT15nKPb2OKRSILsjR9uYZU1
crtTiaTmFQxf6wXGn4aRzYpm/myj8VEqPSoQZArhbNOjW40pvKVHUMe8LcPI
bH2ud8zZ3aYthraM8lnLw5KUFIzcYVz1gXGQuVXeXIImrvCiAEjwnIgMY9cc
uDdi6GuGkVTEq5SNKWXrV1ZispTNlBWM1mDSop4D9TJJdo/yHhO63z53e27o
ynpeZGbyf76ETkWqpwSoo+2aXH1wVRhjkePaFrJZ4UDOESbvrAMDX4at/6Jb
5qP6BcR1zeXjehhNyyEdoJOYJlGWA71VtHSeyzvJ7mLtSmWIwe4ufXdaJXbp
7IqaxTE0vpvZqrfRmmOUsCRTP1hPFTT6opnUzD5uKlKOPr25i6XKAgp4PjG9
VGIGEKZ4/lAfU0BftGXQVj+RphlIdbSpz9FFtnR2LPi6vS7nMZOJdjJcuJnh
GSQ4gpKkrINKAyLLtnMOv0mWS1Augx2XDBgHtYbDLKVdwbg3mH5y9Ys2++PF
8Eh0ByZdzyrosQUHxDs7K/FEDxgc9PRays76jfvdftux8HPuAfHpB3POqoPt
lzKbnUnUtL2sSlFSpMGT9PNIlDm4v5rsnuAb17X2YXRI1veHQvkjukXlKF29
TUv1Xx1kfKsayvKLq8xDmpSop5H4RdofEP6OFoiDxMpKcRuMYjhkWzEKbRBT
5g2lxrhM/8N5ukwl2ORZPaNIrOIb8nDDk26xnkdfMiL/T0rXEMCsRxGFP+BJ
F9scPrmvo9dUbDlYI+ZxCqzLy2V7Nwln2RKJGgIdOemuAkWWi6PkcmGL1uGZ
6vdD8YwfpEwrVqAgBzhmSKSX+5DZu3IVfl94UewsXmb6tR105U2PnFqtPjuE
mOr8jVdEFEVqSDUS1t1pkv5LztTIMVdjJ3daQdHbyMjYL3wPAeiOnr0v0N1V
OK3MkIoQD8vqlLJM8HYXsWqYnRFbqFL2Nu1qTpu7eRueHlO2voEkXuylpcdE
/whUFGguxOg3OMwwdDj4T/DUaVQJHi0zDt8LoH22rZLqLrX7k6sEexh87Xrs
lzCw+bJadhpGGaErgvgH7uhcpHQ9pj5bYx2qa9NYlrya+Kpi2vOtBfqr1S43
7+c2xzSQh98MiWNz1KJF7h7D0/EKU1crfwVH7QvlbsUnvrn1uTzQF4RyeoZm
5wYFou2sTejZhWkMiY67H8ZbxP4D7tG7OhJie6AsnC5f7u/h6zl8Jid4a6Vg
88QOOsX90uPVRsko3xMtCL4NtOGSN21YuKTLyH8MrMKTmGlmA7SVPhx5lVcU
DjxbPTCe8qREKktU/A2FxcM5rkwQtSMPV9zgXyDEmUOQch0j5Os/SKXO7UqS
xfPOII+8vOopGs4Z73wxmto2dhbt1NmTlxAug6PsO4GfV0y8qKXeSYqw2J7+
KC+tKBOtrN0qpq9+8Krol+atJQPO9h0M4+SMmtgEJBybYaIzyW1TwA3G4oD3
aIB3oo0CsQOYuarG4sfScLfqF7Izvfz5nMfjY9+fK1rBi2uTaqbLKcgjTOHS
snGzfR2LzuWSq34WpUoJJEVyirmL38wBtINRQCi4zBysbKJ3J1gB6GJ2room
Y5CtsjsE7fOQACoR1eQ7TYPOdDErg9pHdA0NYFs4OtjUu4aidya/lWJ1jAdL
reMOJ8xqVP2XVNmSgU2SO2lG5A1OYmq/40UdZMmRGq+rMDRxNsajLPQWt/dN
j1bTK5jT4pioz49wcyLYCk8JxUBfihR226s/dnIFoyrlMHdD3F0++HiOSK7V
7ijywZGqMJVNSJ5t1kCCCuQX1hRPXR9Tb51y7UHfC93+xdGgn6bVuGmCaZxU
cXCgKaPNto6AZFBMo0vT49renK/dFi6bphzqfDrFJXiXtSrqpQngVSxnDCKm
F11TNMBit7YyElrEge124tHjss/RE66LocEnq9zKKharKgN7HAVOApEKvPPy
JWmaCZ4T9FVsjV5yoNyk0l5t4l4C0IrMs8HOrDIWCkxGIir4nc+1hMHaPaUR
fw5th4slIYnM7Tt1SUO4FyxSmBYnkf2d5EmmA92bKB5V0ImBfGj4wUDF16ck
l7331RfZPnstHeirguT1nOMfeLa2J+4GjRz9nxzmEa2BdRtK8RUj7TlU2gEf
JUBreSQqmtDkakOfU72dLXGStdiSHSdUwJkwvL6/a28mLv7Bqomi33NcGsSA
VWb4o5/TVyFcnBcW10/x42yhJTggLg6RjoWvdPmnCt078x9l+Ue+OSV53uBR
sBhSXB+lSTUSUXKWGifDVkGPTiOFsoOGIi6mFa/zuvg7dcg2v+oD/VdL57w6
pgfRE4u6j8R6ahDSkMckK3uUL9bRdWo68AfhE0H53IBJ3kvYVeUjtlp+g+Pj
BaHWryFBA0YKq938+0cCq6y2Ksq2oN3BdonorKRHtL9wVRsWZi04RWDY+hJ8
pVDDZs/w4FBRMqwjzeU977I1YEx03Ai/98mn/Jd/LCCVgDy21Ch0/mukKw6q
tCYoxPx9Ijvq2Mj9M5HsbYFctNXCEvXVqVT6WnDWef5y2TGr3f/wr8o4XohO
/7rsPB87OGw1DaR52Go4pK3obNr4f5Oxpv/LaJTxnZcRPkNz8VGi18GtntE2
YljHSNMgtztoTEQbFzt0WJpKmtUOfwfa2JEvGgSaiFe4k92Z2Z+RGh76QL0r
Hvr/J4/3YJfyAxolRQLQTUq08Imu5RAfdf5obo5C/4e1Ur3jQoIxdxN1WVw5
s8DKh1vwvw7fzG3jF247qU5SNVAwTnI3RuUtDqsLLRvvu8xtxqRWvR2TCw3R
HHjBS1Hzp6yY/sPmKeReDFs23bJ57hkXG7TRBtYOl6J1VWFQQEKwq5LFt67D
0LO4RNHf5zdpLdU7c0mh0eBghPI3taFpWW6eCH9b4UIl5oxwYE2xj9zqQGUS
cvYOO1BtEGWmHW54nAbCE5iCm4DJYw30XJEaiPhvHE5iqNXuySf1V915CNGf
p32SqD2ovPpSeKQvsI+kJcFc06VGxUYQxhTi0b+nmMPjFLApfrNw66uy+t2f
pMj8mZrfaJpcoNxpvS8wckCGmPnRyYMe3aGu3utraT6menTHgGQOMfU2JbL9
QcAMj3AEQNdMPBlk5fzVO25KiJMrMx9NIthDwbbCKlWchTgTmH6mbCQ6esko
F/ueraJWJd/H5E+HgE5YZt2bXeN9YyMHlJGpV5iHB1dOMMLL57h81G6A25rg
+q/egfCH4FJIz69IrhKEwYAnOW6WuzXZMPqZ89G16eawSr7m/Vzx2ZM8wN96
5tXcYHYHa8V4MzV+Gf+/KSBTlijqCgKPd8iZZLAL8NCRfX3IxLTYgZJp8jPN
O7KJRN+JEBhXXSMu+P6+zUXjTWZe761OchQLKiYN7bo5AWSgS4t0zRnteydQ
NbVC3VuU5U128YXvHWzNRi05XVY2i4NfiutsgPn+8ZXK+ogXAtZ9Ee3S/Zii
JdRNsv5KM+InGJKQDwPGFPvzSb7yZVPk9AniS53aE0uHox/CFCZwZaI2vPCY
LuHtnDo9QO0WqlyZgp4HaP7rMwgM49oHn1iWaf2JH69awaLTO+0vmP2r08X+
cPdGE2tTHi1uKWvnziN8OLj7yiH6gc4ihJB3/wt10f1xYT1mdKive7/n9b1F
UAZnivngzzmhyRn8DC6gppNQa/au6c0fAYPknkSuMKmcUOHZYm4RDXrUz4Bc
cmAkstV84xo/Xx9ABi+9TQ1zwbcisxssp4N/r43GC5VJ9J6vN2SVVUjI1Mya
bmDNn5W5uPJRcxm6kb/lKcRGSGMu+KaeKJRLfhRaQfyC+jWJaOu+X6aE9LKd
Bw1yQ+Wi0/+wLwfTIlm1Pl0C3/qrjaeVS7YpvESE3ypkIZuzXzT+56CCuIz/
/+r4Sq0YQuq+x0TxH0a9DqPxweTSngDmjBoXxl1dHs1HISiVgICAwQsBUa4I
3Z/HGG14yPI8dovJ4W7MDxLGSbjF7wlL3HZH0Q84qEFR+J1aYGxGnTKuRS0t
d7hOjicBtUFqY/D9fOzEzMYRgp4T6B0Kd3Tf4uYIhqjRV3uYImK0RfqYNDEF
+iad5Saz/KhwQF3VpLEdajyNO9CLGHFHhpBoyhxjCNURVuX4LW/IfDtRflCg
lerHg9jbd2TEfWT/Odrd7kzXj5UK/LITuJzL+N2eXxKS9k/phM6nFvTcjxot
xkqWNzPY98UwdnEkF0ib3/pbs5HDN3OK8T8lE4fTfPAJFj0m3QjFFI2RiUbB
sq7IxF4eRxmBY2ZweelN6pEhpeccTP0wZuAxWfPvh613yj8VzYcAaw6og1Vs
Ii0UmG/8zYFRRomd7/ePqJfxXVbq4LgfBdTyR96hR5UJEXyKI64Qhtm28Qje
6ekkqeJzRKkg0ygr4+Nnt5sS+2oZj44Bv3to23iywlkV73qqcE6zDJu8TtHU
swCjVTkOYdkHOPYBeAraKnwzChcEiARJkZrYxykcQq5RAoIM5CGVCv7Sd0mg
9Cbhujxte27dpFBTtZfqx9YUAr/BzjA1JdE/yTKTuMsL/0X63lc+pv6whCVH
PFaOSDoA2GuAcw3UKuEW2dVO/rkm3if7B5c/Dwtw4mDzNSUz2HdOVFahbOmw
JpmXxRiFDne8PLWrlIalnrJrXCcEnVVjUpspmmnt1FvOJUMOEy/EoEWFf2or
ZtUuFMVwBUV+nBf+KByvBw3YW5OcVQA4FfsElgnhmI2mTfq1m5WBopjJ5T6U
Rp64SSfxKVqRYczhzqDxrQnogcYDvyr+pr+O0Jv/8ISXytdgGYIZCdWjZ1Ja
nK2ed1fMpuXe0QKEEdVgKIVOs9JliECAu3beqWxNTg7p4XrnPuV5WLhGIO/k
O3f2ANr++vhjKGTmMCiisK358I4fQ5yGhF54cCVK4ZtX7lVVPgkz5jG7zt7d
bfyHjt5WLWGcAW2rF8xne5+p76ml+4T1jQp0FpdL2qJ9+7ioUNdpdK3lk2DZ
nTf8rxvP8+Vs06/Iz6xveigEM2gQHWOix1HuTLl0f+bNifqynOvO1xhpeGU5
Qe8/2HUZ2+plaxGEovXxBIGdFXdOEIfUfow7eAd5gNr9EI9YeoG81EuilkGM
nfdl0ehCVuL3nSCYz72tRZePEEU3gCe04NiqUZtcXJ+XRPd+13ebS0+ZQjIB
EuIhA3aR+yvDsfj9hTBC4X9zZ3RbgTJbj8jRYNAiTo0juF61sbeHZ9IsqFOL
xLEHE2En17hJoMbSqFTng07iiWeqQw3oFOLFaGIhCfhKsf7EM+T1KBOhkyiE
8KQWy4PQlB0eh43F7znmmHwu378FqxmQgm2Xpm9eHU2UzbRbSzNGa3uyexCO
xbQn9UQmu8fO8HO/Qe3zaEwdPeGJum0aeTk5dslekfXQ+v54K0mI2ziLs17B
0QQdHOYQclHrulosjQyaG/cDcutGuUwedPmig3Ll6t7XwEAqIT4lpwx1dtxs
ybzqtKH59POuXt6IYu79YG80BLQK5jK3u6N2boP1Jw1fjTgi+hTgI1d1GBrn
p8giDPTSPGI6OSbL+rS7snvUbYDGGpOzqxWOxIOdLLzY24uQhIa0a+JGARi/
ODP2/gsQggykOaHs4GfZZnMwOADGAUKcnnHcsvYMCkTpS8tCvXOYvciiy37X
6VDB763K7xSL5uwy3foZqhjC9KHnI9c5Bfkd9ZYNIR69iTvSjif1AruJfDEn
hShNRIp20yBSekxmPJT6q9D2dM9JZmwf+/zcHKABhY/0t6JlxeX2FlDDNtxW
EnKSXNEvm4mXlbhJmsF48xT74552gdEP1bL0h7GUnIl0II47//XSfsO45MoD
XPEZdTnrsqdLJd4FNUtBnWvYgV65OvQLRjJoCIpozqG02MdevhgtQcLsLz73
sohJqoVXkRJy5pYYz5tWkwno+hE6+0pTe9yLt1YfcoEMmGbAxwTMAbJlnKRP
E5WcZUWAmBMy6UXubeEFqvnLmwZ+dMEx7y7Uu392t39Tkecm50n0zjlWvjdi
38PuToiVx/AS7rXEmB8YgmxOIbMX/6JBYLTEC5uxVE4yC0YppK43gFukbpsM
8NuoEuAbl2VoG/dkjIst5R9rotPf5wfp4CTpP9uqIOzQ+2k4Ywh9gILSraN/
ycr7u6rjt+zWkTB1vtkJy38c+34Rk8kf9neYOI2h/tx7eZZBLoRc7B6OYkj1
wV+k7vPJ7yHTxrjil+5R+JrGqL264150edMjK+VygYKnnlr7/sPe8REMGdxT
GIbc5miM6YlY1Ja5nHgvvzIHpmAWdicGWnfNtwjj2oQTTlJievH/7z5gXnzq
4CEYp4Z1xw6Khj68eJ1NVVlK0lgspK9xnUixXOQ5ZBqtc0+ZfTNrOewPmW05
FDIjVuT1CPtKtZt3m9RRhTP7Lj3yZrJOviv75H3ihj6HDYe3bKgJniFIhSB3
bIB6y24ua9M/PYUnq26awtuMuhU7Ybbgym4rSI3CqsNTeZGOmv+QgxkdwUBg
RXP2K5icjEZ5VlIMLt/2fcOIHH5ES+jfp43cOnmkKAsNwvS0FlppNKxprhfm
HkHt7HHZRiZ/4C4Ok65ls+dc2hjc5F6cl6gyrZngxzaMZd77/kD5mTP+Bk/C
BKVY8FNAo4/cpQKwOWnJw63M9Al0KYExQpBt1EWHJxW6pIlz0RpoisBK/qFp
afKwK03Aw7q3jrem/JSgJXT90HdrwjmjggqllctMK81CQCQBKKPhW+LHwRXp
H6M8m1xWQ1KrTe0tH6aogMuqr7//FXZ3Qz11p+nJQBUL8eUsAV9o+h/YuFVw
6LuQEXBv2DTkQne+tUrU9CvyAqmUp6p3r7B5F7T8ZlEXUBaA+jwf3L4VPw+3
8+4rwmCNJGutdBdqW3nAhswe11wFH7/Ec/S4DVgidXchseySQd1q6a7SawRd
SvccXagV4A3i11mvdUmmQgdK0GKa7jgWtxgMn+7vvRMJXKD1RdSl9BRq6/5J
Gmns1dN+b8V4l4aVFcadyuMDHXtIqaYMiUpZm+xzU3n+5QHQXKkjLMmFAd/z
BuXjA4WBoA3nBys3xlW6mkZQRbOQ9RKYe5mXInDrEb6LcKulbriiGFVHnToj
mtt0WRN8s33YH++x08vwm5mzuc4ZlzaDjNdwkjGdK7iiwZjtwmXWzSQ83ljo
OWpVVKOYdAnIIf0w2QOkzvfBP0bc5Bb9Dj7oG/qZ7nQfjySw2HS+h9LP9rZf
yI1DXqOr1ZtGkW0VFLO0KN6L+PHOeyFvyoNlz/6rG1XiaIf0JxObUhtkg6ZO
+lrD4DHx3OgPYrQxW5V52Ikc/7Y5bSp203cHWPFSz+p2tek29UIX5xSwqfpz
RUUU+JEmHwRii7oAnjRSRb0StNVGD+bo0oHaNRm9ytyqtOvkxhq424Ulm39q
qJVvWIdQjjFmVBF4vAQ4WPePTxwHxzdYJKx6MbR9Spj8n92wpjpuXqLo0lp9
qmj1TqQQ5VZxd7R1Nxm0w8N9R20orFoize/cX6SWYVRj/Z54DB/Vl3DPkVnf
9kEHO3h9otXiCgfacV/is9yIaxKp1S3fPYQzJr/FQcilyRRONHlsqJcDRVsL
9vOmuyVmlZaaiBeiI8NvF6Er3ThrSQzHjDUZA3V4rdpgWSQulOc1OFD+URq7
HQoYgbDeVJRVOQv+4q+avz+2uXm+5Wch8BqGdvm4al3l6kuP62XmssSz2k8f
8h1Gbz1lWz8EhcbC8jDlnm46LzPsaoDWEbnl0H9AlesEBcMpnMhRCuEwA2r2
2L3EKCmBD3gMSsyOO1VwOxt0OSq19RjywAJVnBGFx+5zgSwyoigHg+FTdmMA
cb+uC293pigO+fANfXIiPE4WY+cRoXJiz9J6RyRXryFEq+mCtIXhosjtheC3
84xdqe9comwlpwvaL4Nwc4pGhGSFf93VdZWhL8Ewo0goLRPGmWO3x/bm2jgn
rigSLWAfXv4T+wcbeDg9hR50utKZveWNTVJ2aLQOWV3vi6jZxc1Hf0VvL+Ts
A+mVPm77CzEpOifjQgpkX/X9Jg+SpdiSD1qViGYyVT399qm30Fh+n/7Wh2Gn
6xxLRt67H59/FAiPdH+lLsist1wL20bLvTIBklbrSXxxdqLh9cYgFxFk9UYd
cqm8Z175KmgDpJehif3VOFfJzgrxJXrOsNonDrEwqGFBpkOaDq5sVn2BonNa
cU/eneOaMKJed9hfI93H+OewcNcWcHsNnJ8/ljIxRbAZZjaUd+2d4vTbRpyR
u0+SPm7ZyrJXJ3SXUwFyZTheS7dkR+fC1ku3A7WeSoYtLheBb70/q0w6rK5m
YllqDkv9VWMbCerergUluwpYazy1w4tjqXP1BJw1kopqzNw4VIUo6qPLWdtL
8qojvi3f4/gdFmz7CymVnC/31omzQGDDGOZu4+Gq/Jln3ZG/W2OO9cuRxey7
XgrQkY21riYsbPEZ4dcMu9U5SHQRiPtSUcpfO98z8NC3MaHxihg+hc5PULbp
tRLXedhoqXUrY90aRNIcVpVfYWV94/t+hLgSz1nileCxfLBiyRHD/uFsWAkL
7An2JLG68Nt6bsIRdIoELhVPQ5hmAVfmKskvq2/rUyxCvqh6fO3vwaTEOqJy
nOT6XIgCf1Gu/2I47ngJ0gTq95l/l+p+HiV28ItMIhnt726EaPmJW0CB1637
ybP/DY2bEIMy8/LI5o7hfQ6ouzE93SDHsGpFDE4WFyi7LHKZJzeTbWH+CKlX
MGjjlLghRWBZBh8dYSbnN2GVWOv5zfCS+B8NdMNMsweiAGHGrWxCloYp13k3
+JBlIdUIlKDKPn9vG7dOAvrJwaIjQ8djyDCetq6dt0RgChovK/6GwYI5u/eb
UA/MEfWet56Y1mj3VLeC++pEz/nlIgzZ/W2xaBpEunMY2ooFJVKvvyz5XxkN
QDfOOffXzCZdICF2XB8QApadg+QuvefMT4vFZy53sodZBL0EOob8Q4nvg2DH
1NtXaf2tqXQn3zsOwtHWflB71eOc4Lf6MXZNXwf2WTupOgtAzI0az37CIHjG
PJtmvUXuB1TI+GlPfjVKcm+jeRmm94/6BeJlbi/5vGyAOT0NEdbZGIkvb6qg
BBfQzOtcqhBUJXLWy3fT0tciJuaxXKqfx6JBeeA2V12IxD6DbQ3ElRYcJyzN
sibJwBAlzJKzjyst6/fGmf5NxZ22mTpCb9GfhZ2ZgIgSBu4VAqQ0fkd2a8rE
Japwirz2XCgjNNOm6UwjbIdTdjQ/Rg1kmxTXXBglqvT8hgUdMNOUr5+Jwm1F
Beoim04PtKJFRMTE0fqXH05qhcFLKEFiMHY4+eit7o4HDrvSBGFaSTFTYKEC
VblZ+26J17J+jcK5R8n85FxIol+UZ1ToTkbBPxrptfI/ipwxISui1XP9k09l
OGq/2t5ECq2ysZOyZ9a3ILUScN8XU1wbCebdg9rLlS9aBEeE6/dypnWlw5PS
JkoJBQeinpBRhyMJ5QGG8HtLTbMLFbdMtC5cOuNeos2yQFrpNvK/3afoc2kB
30X5BMyxEgQakU274QNSyDgsvQumajmurzywt631SNvTmikxQjMdFsHgYS/B
S4PIyHDNLQcTi/pf+73tuj0IvFd0u3xWCoDCmJ/YRtqlTdgnrOk7siWT10mw
kWCNZDkNFQpUcMbXup/be0rhXNFuxgwqpufhOyWAYQnDxC6MBoIv8ugfa6TK
ddd002024eue7juTB6eTF6xH22EyOhYclgSE/w3DDx4WP67T6TRlSdD5VwpQ
9+huWIm7YK2GwfDkYUePwEcjcofjOvsOWkvSdvigR7O6tjYTEf204VT+/sFk
j6gGrBwuqwQ7SCpPppA1ei671oB8cpcucN4P3vyzbp2QqEOhQZ90GMTL3QW9
v0E+4Cq1aFlKKoCwSO+DItUxUXePKqvexpKT2tzegD2O7cn9Y/AkMXJpMCnC
LmGFOdL/RZAWf0ya2JAUv/l7KtP+XLeayifbDwjmYN0EtBQU5fER6AqjzXGp
hxnzTfxyJdSaYL/YyQw0I19WSQzr1ormOu+0X83BlvYjfzCTIkpQjkk0FnoF
qgKsUEgUFv4g0TV1H8xLNa0mSQbdfEv9dKrHOD3J8Vc9cI9fcIcrTNBjaX5J
VhLj84IE5iPxQUnsNpWUxOyBhia/vT4MSrvWXOWjoL9dxLSZJQbZiNL+ze7U
VRgeAe75T2seYSYFJb+bQZhP6It2wnazkQkasV4cqTPX82ClWusw9riJszlW
aqPihCOXRmB+L4XExurmREnCpOsTxCMB6c+w6RPcm7ZEjXqXtl30l9vObQf1
EFoOIVmjhdR/8xxD3YF4grVy1AtkwsdPVZo6BCCAOJMWjTCjgZOxWt2nLAPp
ZVUV6uS1PtRHPOfcBv1SnYMLLE9tsiV0MZ/PrU4MXO8KFelxocxQN5RdheZK
b7cEEsYBjF7KE/7na/UmIH/2Oago3racF484xYnBsikkJ8Iqi+WiZkLgpm/e
cubua6m5DSMdZoqFOCsbtLzGV+iXCm8OAQ5EdAFekred0IPQMd2ldkb9IXjT
hR+Bua+Gqz3nHN4w2KMWbf6msq4X/T/ltet8MHUdgd8hm/PyzM4RPDX0w7YP
PH5TdbSdTVV20m3EFls/6M8eqwaIvpHjCHThpwejYFYBPkKwJhfXsIrhThH5
C07Hv/AOe+1nxQEztayH3MNJK8u8mSV1A7sLpDMemX5qBN9EXa3OmVIN4tWC
SL0RWsV+hXdxacK5yQqu8dnw3p9o698GlCi4mPjQnkF0jyxnlGZHfmWBExyK
Alat9VEpkZ34cw75ro4pW0JqLVfqXPWiKVIh4qcBPKKl8nB4Hc+WxobddWQT
kyym/ui61wKlVFglBp17YV4XqQZACVxfhL/qWilbSXfUuN3Odd2aY80Lu447
+xZqbqLJHPH0zZXwBFyYCIzipXf3xV9zSsKZQCRydMiDWEO97Z+dGWZsOnIJ
ziubtbFOQThGyOKvihuldcY8qEA4LTspe7qdiOabwjiJLn+8X8USW2O4MFj9
FUjQ9VrvMCEkpFwukJOuR39W8id/0l/iPtsetIFIwCQ5lMPwMY3eBn+SPrgT
UO3wYNvTzEJZeVHNdp1jS+7A5+hwLE+R5JnteDg3dv6eeQn8xdZFj5lmCTlM
Qjr8paCdsOxmi8QYKg0F3G/ajIOmHRSF9+U3SpSLnw8VAi/GDTSIQnie+CfG
40ooXF8C6834lbl/0bsbAmlK4bhWOzO8o8WiKlJ10Q/JdNpuroKIDchY2Z+b
ZprHgLVXVV5QH4V1qwtx+DC4SICEARz4Dc5r3gsDenpteKEInIaNz7ANZXKd
QzQWWCkWFNVGmurl6Mv73ca5Ib3ZGvUozjiuUcQE6jdq+0lS2URNWGJE2Dbp
Dxx7C0xGZJLoU4VI7zhkJs/YhF4mPtcprt9KoJ12U5RkLVm2kWIu6Q44hZay
vkbFqtpw01ubJBaubVHewBtmEYvG+moBmva3nhIDVxM0Yz25DRqpeONGEz2P
UasQgM05sLQYzCme/1XMiPQhSJcOgns4OioidpMNAD5HJZcHerS9baYnSMfF
RV7OGIY9h4tpfYA8sZWn4mvKP5x87sijdnHbpRO1iqvw2d16qKgcpWkhVtrv
gA7Pz4/NubYZWMXq25GKzLecR3NnpjLroXrEVxELwJT5O2CSrftuIfdp57vd
fKpN/3HwGWJ7hUTrJxQlbRs3Y2ipwKVTwmEvIUod/MjBMQl/lNvJFmCtTwuG
q5Y0hV08rD4oRRkN6GIngu6NtSH0XSAb4yGWhQd+x89EpQgrd+P8U9Hoxij+
47OlIaRi4YJQcx1+z3iLGgHMUcjIg0d+DLCltUweXYlHFLT5xWvmRK7R3+20
ukSuulSvEBhnaCh7yWmY4jSviwwxsrYzN747uoklpyYUYRpyy5njjPHiP7iO
HiFFompDqKyv/1PZcA4GIygTcFOEUU9hyon5NgavbajSX4bIaWAvJrxSXsR1
qxeg1yElpZsTerh8g7ISRqQC/Yt+1MviAag25XiUzSkmpFHACsu3HhOBaDOw
iQXbRk4e/+J/5BqMpZWpFBMMivENn1vJG6eqwGHk3mc7/OLobO6GbZwGo3H4
gB1KjuFvKbgD7fsDTqVeMYEFSjXof+VwiA7uVWwz3RjSPfNkqrYRzpjaE7zb
6dER6kXbp/FhBWDwudN2hVP2cYsRRgNVBDm+b4pxWDuBS66vmS9Kfb/VB6jo
O4LmJhcyaRW0XzhG5RaZlUZYDL+l3bilV+85G+csk4OzspFw26TUqDPP7f/y
agP5/RlGZDQP6PlXUpUsEx7/RwojwPwSj+TB5xOL32N/wBct9D1CLlbXmT0f
KvwrUpjcKuwoRYfOC8LHxa5xrwmOgT77aJAFReXQJyIE9YzBdW0GwKWzlIu+
NweKEr9YrA/THDTix1GEyj21TG5VdvD49v0/wq2o7jdKR30gDSMVJygGov+e
86sqZ2aioLvqVSBqzrGb0dDs8HtrEpEtBi7FfSNtZvN5qW5LKw7kOBNkFcaT
K/PW80umMw0xUYXkQ3e5Pqe5Dp+Q2a7qVL6IDLtKILF/HCV0lgi+9wDgMGHn
xbEbRyTnXlWn8HB6hPsBqsuUbCpl5f/fx5JxKglpnB4ENbnfrBreQT+tkCLd
W1XH26ZfeZgxnkd93h6sNIgypTwuc2REKqT3kQ+IpvC80sTQY5xFWQqhDxgj
GT4+Q0D9pdfZsOn8M6Wy8BQmmXJqNOsXAUyFdtdPo1d2OiHPcXsSCjfxmPKP
DwuBxZ9VjiNIOWf3bYMdzdtLW8LgJWP7bEAZcg8tlrdiLerMkVJOhwfdGu0M
osqfZCEAYfIVSLTXye9VqQ6I3UFpb/cGdciuzapXilwKocZgBs+VJsEd1HWN
W1CNbVz1YEDxqE3KyvK51LAYPIdocFeFu+Cx8r3S7pf9uiqBCpA3xUxxmnye
r7w+G//MyerM8mpbzlVFYud0O9slNpuk7jIYzSBbzdJiwTKBOTF5S/ZgMb5I
iMKXtkmNiMaB9L+Mu3zTZgvANBV9s/VGawnAllLTuk4D9UZtLiWrHH9xlw5o
+vbFvoje642kmEnytJIit+d4LJbjTaOaIks6XhZxr0cxTOk455NDAGLWJljh
x5g2MUOAR7qZQdxOAr1OYV91D1JLXvQEJWIK1X7jRFaZ3BG1XwSSO23ZEojc
dfQmx8X/fGl4ESYb+6DtS/iXP1dR7uld9OMvtbNYgxG6e58xzShs5W/09ftC
8gcPbXO+JnCZ1BQs5o4Qi5VppailfGw+FNsHVLM/RNnXRiQo4PP2J/3hI4+O
LfORFSuSRJVprjKSIDZ9iOHyFGLMbOd6RSgMkYCll8OEkbpdiuYcHujifQxy
LLwXIkcaX72sfS0mGGyIqsBfnXAHRAoAdyrjb8+FaZdE2z3BcO35UoGkxWmA
9O+Z2cGGP3yVvcV5m3BShi13S629jSvuC+36JPBCKvk8e/tGxcu4JOkirjkc
CEcL766YvvUX9ddqLl9m/QR7pYzDn2unW1lh4/X8fMJeMUfXmxjKGukKkcSi
GVWNx1t1wovQkezcUUjCB8yBkcmTs0rxj9qFKDNCoievTXBN101cDu53yYIQ
8p3Z09aj9FV85cPhp4l9BzbWcUmkWwxeE313DSALOjgne91JRaOjiLFAbdqQ
ehi2X3Rs5UUSzcUrApYNmpinpLqpKPnbHKXhnUnQxsgHVPXSCbaTTZRY14QY
2TZd6p/Q6PGDcFNOfyPA5DrgyTn1ClF9K8nYnivgjhFGcOWlBQPbyQSXMAu4
o1+dPco28URCosocM3uulzNux/wVMJANg1+6mrJVTOs4XkQpBLtiDJNCBDB7
UmWFfHZ9rQ4wAxFn+6Hm1ur3+UMeInB3ucz/svucHSLc/WraEHhybhvattTQ
h96XHOfc019TLxz0ugTNZYxObkGDgzrmTqu4QxyPgYBU82WGzvywFD/lZiei
SEGlZJX9s40EGyD68OfpbkAs1Y2w2ANMdvd29DEkCId9bewQyCPB/lMz5uqD
ocF1S+wD9x87JMc4VRmiO8XJNzdwjkQrT/x4D6KSne9QyhLSOkCewETz9bCj
yHJDeXOkEKv0e9G9WD3l/JwfCsdEYamYCEC0Rwd8RVH2jafqL2AI0kubwQb6
ICY59dY5ldxzocg1xLG1rsV4eAp746zNkzDst6oCmfiHpkjv828OUkr1VMve
FdEYXawbZhSnoxQxCN8ggGEY683xEuPB1WCQSEelxn6hXQKZtdzUhntcwvwC
RWvsfkkR9e2YShIFyPwmfJfmVsZGKKvih2SfAEp5p/tKCG2xU7f7HH8qXbs6
ZcIfeXGwc9RmVpzWCCScHvNTa7qkly+Tm0W64kwpSCf/eU0PXLgOYqgja91A
8UsJUK17rggRfBwEI3g6JkwQy0tXgO5WZ49Hm2+Ldk7s9aCaNSclzoGS0de3
1DtEU5qx7GOJrpNRPqOFWVb9Taqip8DsYZp/Uy6GAXeoet4D4UmPSzU6YopT
zWyWnv7qu+GIFqGYX1CeNEP3hDImde/xlV1fLvnzwZ9IdxG2pbrf+leN+5lM
icHA3Ochh71uypn9xjaePhH2Ah45IxFf2jowMrKN4UIQCSrFdoIkPLp3Rkk9
XiZfX2haFkGpswHRVKp7+YovlJyW0Z+vDN7dgl0MalGbTA41V4kAxrRiCZj7
Fm2PAsLDexa5rYUP+cxi2vqwHsip+v+VrQllpsK/20HdGzvWt/u1jbccV22Q
8D/pYxaL6qmmX7FF4O2t7DXZK3kTpMKrT1HyzKgSjtTX/E2yzT1lNzAZMijs
g2sXlkvdRLb4PvJxsiZXm3fP8772t0MJVMSxH/Aoa1HDEDvXG9rGiw/nOa95
vq5PsB+2C0VbfniyeTZz1aHJUY7XJSjPXS9hyzN+hxQCWpewllFyXLL//QAB
cndmZ7xoOf2q0KUOyuliY1X6eCU8/kkrAm4q7RLPbL/FfrNa0pPuvcAEHNrm
eC5CMDGbF097Q0aEDqZWHN1RX44eW6kZBWgchXP7bGRGsE6soNAUO9F0O46l
sR/59Sxu1+fkk+Kc8KXT4Of1WtHXcqwZGj/ZbHQ0mQiOE+/vg1r3upjkJldn
rTIdYGHMAVp4EUprV7XLuWQOmSwpaPMQ86MapgtBNhlAVBMKozRizKdN7rFc
aSKOgJUAwamT6FyxCq5WTL/4jrX/sOBc1pKMC07g1lJQ9mtdG8CBJ23v93C0
bB1HAPMxaLFDFFiFpzmmS181ZKMDYdUziF6XN3xpz9PNkCJ/T43DRw9L/C2g
k54H9z1NEimnqooNupX6MAEdBxUgtQ3SBjlVcnwPgEKcWugSIQKqoVmLn4ll
L/GSYFXmLrPGimrnSvWTDQ/e3gIQqyeffX8/zdqQB5Fn8W8ARscE+FE2Obx1
Mf2Gk0xEUz6u7EXciD4KTch3lujlvgBTHs5wJX/7ucKZ1JkDoWDQilyj4xSH
tm3pdgUOV+bstYG4l3U6Mu4+dzcxAshFqFnK6396lhLFLBijnjQnYjRc0ioy
HvGqDAI+DE8uFQ8ob6OO+bZdH4qPUPEpoEUj5hgnU7F834waDK1WmGGbuLGh
5tRsyGvhHVyoYamFXI9lFENgLv54C9+oyLFDwoCwIao8WLFb1RxzujB8Y+Ko
eq9gaRRU+B6uGYu/SVNfuPh6FGZdf34o0GpAkdQj0ruL4AnPtuax9a4r10gn
GLJiWaPmZX2hQrIGVSqYU4zLTPpc94RmfnP4DEbuMybvVrmQKzwfQ81R1y8o
sf+FCZgFjs3ioED2isDyXsyCXilcDF929yiQr0jT48JiVzSYUps3Au/LpJ8P
V0aVWR9H6Z+djJ7OB+Yv7YQT1nfuWbcUvZBYSlwHRDOOsiK1vuK7RO0B68bR
gRAmmOPwcNnTCp6W0g4udIcCjmTR/9+OM6rWrX+BdnuJOYa3q5c3tyepTgN6
obKZKavBaAfeoBBRoA+kkXq6Mif/jcSxvPjnpqpg67w8Zo9Z4rV2R6nZ97W+
T4cZC2DcoERgHWDnWA1YjHuBNTs64f6iWUzHsS6XwADNbdObV9vZu6ePpwKF
Pz7tsmXAJ45uDVjBm6gazIe67dU3i1sTRfGLq4syyjxstFQ0wfcjzLlhKH2t
XDpHi8wD/ok5KRVmQe+9U1SrZ4uu7Den7dlX7rVejcYkpO4cdIXM0swpbmqj
ONlYtNU2bwx7xYCKdgb9uvFylzs50OXTIhZuy/I2mXiLK/tZe8feoly8xTcr
aLbHmYZBSHYus6xj49BZTTApTgoD8Oai/Z6xFvgqHMpcfWkF5N44JshBCqlj
T6OgYASkmHySV3BQgXAQQNBa7Pi/wHIV3fQ7HcLv4yOa7W56Q8rJveIngSvX
rrh0b1W4d8GkDvyyTTyYNysdZVqoq280b2DI2doJ2sGwHU5ig2Oc+L+EkXEl
fwN/ehOnQ26eU7bKEXGQq5ZlL3nI3rOfO563veT/sp0M942xesO6UgrO2V2z
4Yl2TmXKf1piuDpPiwYXFwZbnmVuinXc25PQZIRnibGwv9bRgP9kYxcKAhGf
ugmYQmAKlbjJiPYHs080EYKrwEapIklfdMVoKf7mY5QIaSXKcZ/FUjj/fBh2
iLuj5+pDfbN/vv8vlsn2hXeSJ5BNTAfOhka8hlBNnTup8Nq6rallkEPH2PAG
fCYTVCZXfgs/6X3tN0zMhZtH88HWyuOSwqNo//crdWcYVuJ7ChUoXgBiUqPE
tnSksxeBwkjV1lgD+A3APvSjaXOVVEM+XHHi8jLKvVzsKKe+dGbqUjIqOqBh
fLo/HSWju/2xsVxzTXX+zRhnvY1Nj7eEgy5U4Ob7lDdUOL6McFW3jexncjG7
QHoDqhe3p7EhLlZzEKku3zhZ0TgGdh/GyFeSg47TgOHN6qqQId6HHYT7QjC0
gebThkixwXidmO2Jv3n9TLeGm8E9pPb+hbHy0GwhUxoznLodi/FmWFQD+9Fm
qiaJcYRsDAmRVr2sem1ncPULsjSorfPiLZ3cbjKG6BG3QCwcN+89o70YUGQZ
8fWecw1E4gagk5xOdX65JjKGP5q7wDe4UlOonRjj+/+mW+T6EhfhyWJd4BIn
FHjEfWyVAqYavI4o9JqR7Yoa0+l98IU7NV3okusq+9N/E6dD/KNwDVPfVpWp
p0OS7LwGcCcOp6d0a9av+K/bE9SjAI9uXdwppTBxNIBe9JrUI6g0M24vaUX3
0A9P506UPklTSmbwyzaZzFp+0MTSJJI3UenO5D+Yw7Q1Ul9itzs/lqEW2/48
1Pr+5tcIxgNJlddjt1DcP7EdP5rolj4xU644QFUdPS9aZfOwtxnfa8/6A5Y0
E2ETk/JQSMWuOiujqgEYTcDRgUiIy2xWdz4E2FmsHWziO5YXnkN+w5xV4Igj
9S5ZiNKmw3/kR5nyI9wxIqPdp+Jk5JnbpqfWttJR9KVk1QDHr1+qrknsIw7p
2MW4q8E5rvdACOEZsqur+/h4IgWFLgaA4AHW8dtYux/mjYze+KxXR6AaxwoX
dU9lFZMjmIrJUeVPor6MFDrDFzcxbq8j4TvNyS10xP4BKdVGuRbzDHV69e8b
wISWnaC0uWjwK6Z9f9XYSOr6yBZ6U6NR2bIB30JOrh9g9Nurt9vQi7ayxhSm
GvsGfuudqMJlIuzEc+5x/OvIrfI8IadW7Pm6ql4x68zlR7OzOOH6rCGCThaC
TFTff4fPK8uH2cq/OmofTT+4sbSyNy2EfDEuE9+X/PHSXCxLCtDE1sHBfYJT
Wtwp42iOl46qGLF7MJk1FSZVV/zHoI0a6ATqpEY5OuOy3JlckBOQPPrDhgxR
8t7bCdEdqQhvKad/4xhPXSiOaCi7g54rzQCNIvGPiRwlx708LbGSzfbR6JLT
p1C1/mx9dFd7lQS3zllQDvF+KfmixBfQCRG8f49e3OOPWGBbF9luEp/aZk+f
wUmnRhBvKw95wARJmUuzywOm7fbm8cfwZiqJccgMmLWu7NUZou2wVkJ3cB/P
xGvDy0X7HKnzu6Ud0aggOpt10F6NETntoG+WwPeIYCJCLac+JLxEkTQLwVsC
hskUV+/3jPlHBKdeCnzjJFfZ6GbL4pYn/rrx2v1o7nkedXcDtXfH1aY81x4C
UCeDU/K7wbEZNBSjRoakqaS3e1HSKCw6U3t8WmJdQI04qiBTx4X0cLbI/WJ7
z3xLOm46D/FjqEmeXDWPG6e/TOHfUoC7mtyBsMaEAzYsGvI+INA6veK/z7n2
uKVoR6QqISf/p3Lb5sIwyw8THKoRABjZpei0uUWUPdD6Z3D7c8G+rh+pRJ6c
l1IhudgbjGIX8lCh1597bHHyy0w9VrmeMxKZ5+Gb9WLxZWc1RgDz9ajd4xHJ
FCa73Z8efgIdCjubtEE05fhTdzqRUWesJ39ROuKryNqB0dPqiA+nmFk/c8PK
fngz/5vZdFN7JxyuLCkH+locWXQ0e9i79yw+jAV6ctf2feFE7RkPC435o8p6
Nu3tz/pbpoegpj9OQOgGWmz/rc9B3UOV5Y69/UsEC88345JulYqoxkOstoIe
i9qyB1xvluWP9RZBo8g+0170DK8tAZkeXr2/8Q2rf9jsjfGVDKOxbc6m3MMb
XycMf/+P8cMqjZhVnxKqepLQzxZNcbvHWCsqCG8kixrl1hQv6rvpVp2AiXSG
d/VWNp8Wsk7XN7kOvLJ993V3+9SlM4sW1H5Ckv11W+0U7cZU0OQefMLqaGJ/
wKyssQ/HQY4Xl4cUV/iznTIxKev25kfclniEoX3vOCbIzX3dSixOaOspTt47
ABCNHaH5X+kKDDtEyFImLdjlrEKXFXv4PxAFIQ4wrfTtmqrE0pK/kDUP7Ls2
3NL/yJF9yrkaA4+2uvctcgX6Zlqwfj1lKUCxsxpDkF+d3KBw+n95h0lNXHcI
Ow4gKpjEZ0s0oCtzqUycSLHkTwoR00RDthmUTtFxacY1SjbJzEavLmYhXpyr
R6HbpNZhDl3RAREkC09KO90L7+LtyECzG5yhuoMaVlgFUNEB/l/hWTyCcz9K
it6i5dUBXRHAImQmM+5lE1uJdqQFU28Qb87thex3Ksd2v5h4TE5pmU5wZiR2
85i9R8oxjtV2B+GIlvsYCznAL0KU0gwBMZmEIBfiErmZ7lVt8CsZV9WefdjG
3s1qAzw679AxNst/bZJ3+U8nAXCBQKeSmx1aLyD812iRgxP0IEpjJvYqPVOe
8c4umJfMkURe0L+LieOmjI6hEpgLR6fIQsCvD4mv9EkHsLLyu0TlZsjl8WfB
FL8emp8Alu8quxLqJqAbb+3IRVFW63GE2CJD8SrX5s63jt6leED2Os3qMP/9
epuK1ZLvVck2yap08vPf5IrVxoKZfuxgLL0VtPRaQCjr1OMcresVfMsczZ8M
58dgment6fqES6sYQx9uuJZ12TqGTy85D11QylWCNObeG+Uz+D48f7TF8W3z
jKQA1IFllxg8yHzxIM7+4P/i/+im8KEGDZkXauFT+Xvr1IycFDfdJQypAcak
JmTi3lFZ4VgjF3jyUEQ4XBWwEx1GMWq10Vb4BB8LIBFFier8waSKDexbd+T9
6kG3dTjIzEGf/1SyKOalrxxKCPjRjLK3I1ML8odTQtbyufmTM72R5JH/RIT2
RBt1m+TZz0YSeuTMUUPScRgL3Fh+V3JOZw3ltMZn/znblr8MlEZTMw2gxQyn
KJYVUmu50bc0575FOGb/FXrv2cUBTD3QFWbiCNah+OdK6Qm6rODrqeI6MLnp
SbRROg78WiIE8bWYn4Cdyl0lXwfgrzqH+rnJULaM5nfkCgfDlT8ymOBHyPIM
d6vVVWWhgLb143yg//w3vt4RvfevwPvIDIVnizFG2M0O7ZAmy+8lVlBVZVDV
BeaFFr99Mq8u8X5L+vw5wmFKPr9SKlMhmtKUgf/md+SZE04KW8jxRmdEu3Tk
miV/EeXp82InscQNG/u6a3RAiGQ+pCjuzXBrGyQS69lbQK0uIobwvkTQl7pu
+jvi+ScBnPxyT1VOhCj6fbYE1u19/3dimEBr6G+w25xhkHQ440WquDKDo+WZ
46axNUBrTXTnwyFMy3E//RcfeIl4Tx7EUiGE4hZdzh6qWwy+Srvmnn/a11Wg
kjrM7RjS20Q7r4+VMmWns14Tzu9rk7ASGN3745Kg6Q30kKk7TSOdRvrLZIdZ
aDYtzzeSCpIII6bKYzL7dEZWnR/WWYHnnL6+50T1+1o3WRMTUL/RMZqf64O5
bIfvDkv/Do2YM1btCp8iSZIVQYv7cR0saaQ+Ye255ytajCS+ZPs/e0YUZE/u
2uNGVbEnLlyIgAHdx0LQE6j5uChGDBSQu4AUMBm9xLQn59REvFoX3QVG/ReM
zMhmmxxdK1bU75Nlxiq9DwMrtbPp4dY3noIPKZ2/EjUlqhykTBHdl7nXzWTn
/pupb6v33nloOtxiFgsOOCfyqkApFibTju5mmxYoiChnKzhO4CvN2gyNw1Yv
XXzWa1+epUxoXbeCaBv/MftH+uHsat3v1vcCkoh3okdx80OSlAWtzM3Rwe9h
IKbW1pVeRbw4XZZw5nb3vqU/YGkr+waTH5v+k5NRtb6VvZlyz0fp/jLOHhhQ
pw0Rr/7M6pWzjOxgexTK6eVaVmFiLejOnF4qyqZ9SkQlJEM59Krt4Ghlbr8l
Z1nBSSsukNk+NxmkpAUPDp7KkObNaYjyB3UiCxmclVRc42GkJB/eqy4gzZuL
lcFj2zKZBQ7XKJdQMQ2zOMOLwyV9tMGYbJG7kV6CBV2aFVfzXOf2ccQE073o
bTynA8wjOkZt1zhZ9TASf+boQKQjb78q56EQCuGJeKPNPL7xt0yPNMIhLUpu
Jls7rjNjecYXZNb3HExJVYp4o7aW/6clYuTreyZrRns/P15VKdq4aQpbn1Lm
jcuyOkVX0/d8hJrpg+m12bYu/ScEtoJvNz7FRML3xJvNUUzThmyiaQjHE6Qg
e/5OepoUHywFVaB0CdF2EeCle43XlpH8PkO+2zBXsSDxK/L94Y5xmkMY6OAa
aO9CTXYSA1Ob/wUQL4x7kmtrElvGuFj/mmU2EeIkJAgB2uT5vRpUbholA1Kx
HItbOH+JEevnt1KbXu1PjZ+8ivmgtIlPRlchQi127mLr73bv72ws//NvIvcd
MMzRQSd83BcV2m5vvsAsCt50y64WY+OlTp0HrtK2/YyyfS8nEVKThmQNBGFc
AWHk+M1FX5YPZvf8Y2gJ0XJSBEupF+awu4OFAOvY1oHNTlMSLGEhQtSbRbhn
p0WsDKsFhlYG4sfR5ec8r2zzf0ZmKEvQ43Osg12vTHQ1F6G8LoefjHMhTM2e
SlngZMeQB9mPvzbcCajDmV9sRLPCEtQkFMJmyEDYA/5iVeC8hp8EauAh7rIo
ZszKNzSDhtbzyUG+kCvT/EUNi7LTfLO1b7uqM1TE1umDUmnytRI9ZXYgG7kS
pjWp0AbjbGPFqFhsBaFdpfCSCcaLCIb7Rmv/eHJJoU484zLS0jgBLW/doUTl
U7+m7/lm8tBHddNLNu2eDoj3SarphrZo37VD6Qy4bCifCGIpYihQGU29m0tA
TiiAeuilHaF8o6F/MOFQrkOcWkHD/FXY6kQnIY94MnrjKonFnQa5eShcGhYQ
A+TCao9FMjXIg6LnOEMx2r+EwWgBLdaWoDb50FV6eX3juPiaiMumNquhYC2C
DcinR/4e1S9WsbKyX1MuMCzY9pWG1OtejCOcVHxgptzGdGa8hfhLfWDLigCp
w3HtclO8UoYeGDwbygX3laj/byryXnMH6EXHeB4+rzV5tL8FBvBCbR8wRO/X
h64RFOfCU5dbWRNucFHAORSwDSCc4EXrKaQ8uymTZ8choGkoN4e6z+QDzCnZ
jp6rWElFBFd6ATIFJcU602cq5M7cz0/DEPu7gKr6JUvdY5N7/vE+7PAH1E8U
btQkQd4irPSgYC0g7oNZOLeMoxlhAnm3WL1yg38oua0MVWY9Zu8IiX6EAzAp
Tfm7s7wAtBSWG1tzvu9RLw/nx7z1Ox0pNSRzBwKKDeQaPixF+Rtbch21jGfg
y74E/FK6fWPe0NATdShU/NDVMFIBvTMJfzthCHmkFcYLXH6qAIvQ1gcAa1Ab
JJj5a2OHaXBczYgCANVt5AZFIsTYzgl0hQKfnvln7qnQ5L8Tr+lNpXaHU6on
PnIJz73r7bP2SnH3Eyw0QwjzSGVlbXB3LyMaqi0JSPebAUhXNpoOU8DXnByA
B2/0EdrDmIW8SKmOwClc41MR1hG78sBQhU5v7TUMSJ7xUakGDgqAEunRqSdD
9+3krwUUkmetSSweg2bpYa2PKsZSDuuWLMPQmE/gIBIE50o51KiMAf8P1E28
3rsvg6tMLSPR3JSeN/xuNUyVACEp38cHpWR+5qUv6ecaysLyaduZuDfWq/un
ovYHOUIuhfoJteeOUShoHeYhhHUDz7fRP/qp6tmGK7qu3wia+m50+LtZkBQ+
8YiWIiNw75WEpCczDCVonKFBixSgNZ/2wPeJ1NY4QK6BF2UWaY73yANuRfqe
zD5X/E6iG5qoEh4Xl5MVxcsxm9unV0cJ0wRZj0B7/ZDck1sbotR36sfOT3AL
EDRE+rCmV3xSC7L7zV8DFPxk0aRAcuvLeHGIQqkSCubVZfleyPsb3PRgVo8O
YRSivgoAhGsF31bdszvvDpm7W9a7cMTiSbbI87YYvusKATaYwt38J0jaqJxe
RzDpgRqnvb0mGA3eIhZEayKpMYm4Qb4lLhmatsH/mGiV6Zr9eSkz4xW5QtAV
koVNqbFw1eOCHrC+8eJg4FKkmqh4RhpsWO+V7jJt+ekWmtzsehd0h00ogHwT
838TAQA8aPFEv+Po52dJt9/nQ4YvTbHaW4VQsN9QDrMrCCVWL2w2geRwAOZb
HDYxaoY8zeMRVTkUfHrtOrg+GgvPJgx9ts30j+BI9gLoAPiXVrd2Cpe/LvHD
bTg48CR2zBu2iWYQ8rj6uBugAyAvRqSTXYXXI1+lwyNX6uidh7c6S3eJKNKu
z5BuIpvC/ZVKVdEeUjWiEMvcsfpOEokX5VPuO3KNytuNubNEbelh8+AvK1r9
hmOBWtX4sLrrTNMydpQ8ac5KUEUYYuWtJ5A6OUF245jZmnPtGPdrXtP5L/9m
7Z6y6ae7pQX9ntxvI1qdkmg9WsdFBUrmJCs4SJCT9qWL1zBVCfGOwZiyF69a
qFkGKrZpWVARjc5sPkCVesztWQdafXPOEof78G59wP2ik86aYqsjWXQ/az+S
l+ox8FWu9aGfoKbb9XYq0ztDCW5qivqnSS9Jd55quxs05ox+M467SrHkFab+
TScBP7A4jqN8OWei10QUCFL2tRVdO2Lc6dOSVU+a7KS6oSQhzwDPw1TehmfS
dhyhrDL8G6VT7TAiobry6ybDFe5puGlTyXNhwDolLJqgjRilhX5wy9EsZ7Fh
PFPY2mTTdxLkWH222HCcKlWx2PNXsH7B1GHg7bqJkN3tozIymGsAPDaZhb+h
xMD6rfwaL8ozEY+rZWgWaWFBJUpXasqOHoDgeTZT/xMxC6bIoE7DzHOaNqRJ
EnAbkNWTZ8OJvSYI14b5BPrmuo6vhG7s/chV/hj3TMKNWxoDApuKcAMmIK7a
3HAqkUyj7mm4uZudU4NKZh+DZRlndghRnOu3SPmA2iP1y7C1/NaDmPmqHIWa
VXLQief8xygzb2cr3kgzeZ6fPUcZCSug5bac7eJ9g1We/z6dfJx5m8yqeT0q
zM51azIOQvx9hAyFkqdZpfPQPwM8vrdDlDqGualt195AnMie2McUMafEOkyW
tGdJlQbTpur9MofrVi7YeXYY1tfy0RYZGnOSt/lzM/vuWKJeDghTx2E93JVq
S2vKLtrXeAeoLhUBsGv5Vw0BTi2MZzfGS5aodWBX13cIDbtPo4S3Z4aBP/oU
detK6J5mdp6XO3L1t6hXGKs4MVR3n90JBM1EVjF+T/ZQ758iHilkCQBbNWZ4
TX9hd3yEN9NqtB9Xb0oUOTsYKTyMByiUg1JQKiwW44fcjcLSgUPpoHt121Wr
fNpE7sprq/e0AIKSezQKjuboV8bT41CBrCk9tNSuaww3UrGx5IXjCqbvBNQB
n7x6EBC/z8NoLGgdcLRaOyyYK+UXdx9E06JEgXfpSHCgvGlXSfC0MY5s8Brp
NaxtA7jhVF8O7dd6S7cNCmSqN/+GRpcjh9WTp75z04gfktpZj3ULJZOPOQPb
Sg+JGm8KD6mpY6Y9clVQSMLN07T4imMYC9UmYLC5KryUrb5yXa51JOWicsD9
yA5LFOdpg+15WrgfNJDISeUVK/1lK5huaTcAJqO9/41H/OnqF+teCe0uiOKx
QjVmrm9UfqFqVBXh4TZ787lD0rHey2GyvI9TVoi1+d4OhJtuZOOlBZUbfvD2
IHgnGjoP/4FFiTOJJpbYYPtHPB9D/iOdCJ5n1UZ86xwXeOF3yT3JHQsAyq/7
WaxB1msrqKqqmDn1H/CJdYT8aEASFaI0s03pt338ZDkMgcFQ77ICK2KMhwLi
QpOPS3qBw7WfmWIcpADfyLNW62WSJbxttcXpvncRuNQ/saifO+jZh1Q7qtuF
lu/AvVKqPEljkSCLQuvAj54LE2QOXhlAIPdl7ax4xH88VVn+AmvtbE4dXJN2
VL2E6trMiCIHcD68vskTW4XZRW1y3Jwpfuod5FmXMGpwZAL6SO9fRGUS9ycy
DarRIlHa3Z4KXL7SjV/GNJpXLo/MD0XeGWp/uHKG/iq6JpQGDdxJIcWMa650
g50zChkoQ74Ia/yB4QWoWcXm38hXxPxZ3fttNZJZX4D0Ty8w6jBw0L518vVm
ozhytj3Y3SvTbzdcq7OvRO5oP2q9hsCrCEUoqh//gAATm1O7Zyk0GOIyW2FD
hMVoqQC99J0ljxE1Lc3eejFj2K1Wkj80XEEBpkbITnszgsOWs2SRMomYuVmY
dEiL3zdoUouiYs6P1qTvf1AH00aXUXQmTQNjtm3ZJFV1eOh/4kJ0lz64xihv
ardTL+hc3DF0/1/vQaHVYervWuxpzF6FY78pzBGk4PQN3KcahfeGYEa/HIqo
DJXitpDBqYCnMrHBTeVEhCBF1rajxQCCbmEji2NGO+izAQv28GsJhQmD/e2U
RniTb0ad/aak/gImR7F2GLR4JvbCLguMZYUV5tfEr76I64XZvTt3RFk0YcfV
4LYKkeMkQ9LoJo0zr5vw6oGVQVxorFFaK7uS+DV38bxCjVX9byKUwC8j4d39
nEWMpNxJRuDoUSdzHyQ4npiAjvX44sloZi7j5hlqJWPgZFMDc2yebAdaz/Zn
ejDDJlg5QSqNn0jLi156M9bXKHxT7K9J2z7JtrnPWEqg5i9NRD+m740rdGjt
L1IBK11wSGuLnC7mZZBR91RL2V3VybgwSjrBVRJl5lgOft8K1DVDfL3n9TBD
Fz1PjgENC9d1JPI48E//zpEUUhbrJ87fQ9Jl+yVy6QHWzU+pafuKn4nwIOID
48ZDSZDp2pR85LwT/ShVmNUzFSHwDD58uuHqOyE/mgCmcopzUqmkpnbYJ3LT
UV67uNTOUm7LXN0JJ4pqIIhL92nGjiM7WhSTJkKG3ALQll9IGAPXRHlz0eQl
1X6czOtnPpPfA2J9JEIyJx0DmM3Y+8ua72HDe+XBGXqGM1ZbScPWfU4NvkWw
lzEA0US27J4AQyNRE/ccY2fd1w9gvOKAfRJhqKA4KbWiZNtvvTOR+WPFDEWG
vXeeZF3HV8dRlAWt4zijR8/3F6vSQ+1QSejAvptQTmxhUqH+sorex3a9tJo4
GlUihJQ3WTxpG7ECpyqAXOHUjijje4tRrsyUT+rt2res0wPLY2N8p+6Uptm1
NNtfraEvII0x8FKVBcLuZSvatzu6o4P5p1Ie5o42/pvDKqLUJKeQim13Xw7o
zQirIQJb5zGkGSpSzoGKH5IMQdG+MFpPctvjRANE+kugZOa9huZbjl/dtK+Y
mFNFWu9CU9q0H0EOlexF2Y9T/naRK2xtaFn/aGHN3ARjylVXWp8oMaPK9DQO
7FXv1waqcBbgi8BEp0zttb6Qe80pY+5TKqlArWqyd1roCP04331rL3I9NQHM
15rn6TkEpXItFpqSuGGwYEuhJbva3DRyNfQT3lBA1l+mX9w08OgCHqbkd3dm
iMD8wf4LllsLtoSTmk2FdvW9nLSt5xNYVaQllRovzHswQLlFuMcqtbUhwlNy
b1JmPInjyboRmuF/aslj8Yvjy5jEBcDvSfg7RqTtiVeevdHh1zC6198aWgjZ
S0boMdw19j417sm2HzMAyhYQpyW7kIVk3sUYul1g0HAjUIMoyvDixmHNw6ut
PN0dNDjd+UfDZWxOApsSv5R4OqYLPj98i61Hfxmb4u6rwerr/aKKsVwgsF/l
u/zQ+Ug1eUwUID6opGBwqMgRIAa8I2T9SsO4vP4filILSRUHoQz3Z+OiGOhL
UGePBXy5g4pfN/UFyEcF4mAghVaH3E2kFbU7OVKHgmDCFqqEr6V3q52aWuMk
x5ctdLqMfYb4e0Z1jONQsHmpKdbyhVCrx9AgOltQEmLGhr2xjTWc2XRED4hP
aMZkfFO4+eXtkZpmtGG2WYRodejNbi6Gy6ZF5lthF3948LL7V7d2/UNZtfhi
2B6Siwh5ACAiAb2YuOVild3JtdWb/6lG8d5dNqZzDeJ4DBduY3OK6Wlh9AB2
nTJ/8kUIIx5rmuYtXuaVFHmKcP4LQBSHn5c+wK1RQiMDhdO8+WCWTblkOW6k
O+K1hCb1HRbppB3euD7nkZKv04wxZcBXfEEOHjh0qchHku4HkRbWVLuyWY4i
iErkpBfaWnv5sPY1772MLvrdIkkSRWOW1oMJ720sW7BmNii/wGozQ/GwsDg7
LKR9m3MCNIPpxzLvbpwuAZCTK9J/2znJ5kCZfzvTLAQLDebT/79fqh74vVKy
sZZVuFQX83gIokeiKFnRH6e9di2cQMxYhkJbRZ+Q9pAM1FE5b1kXgsU4GddA
LVpV6GXSIUGrkWYqOvQ6XXc3yzpBTm7FoTJgVmisEgnfkwHH2TsDjkoH2/Kl
mroVJdAuOFwLe82yj6dVFWjTs3SGbBgdYe9Blsf3WoAuzxtE5hTOtVFmHqo/
QYwdPI6wgBJbgM1btnyOS40X7C64BfFaJDLpo3T2b0nsGQg+gKE5bBgJnceA
E8klZGrKLVekbeZq9aTWK1/fYJKMPVMAbYxqTcoquF3ubXPgYMfJ6IwBs56x
0fD1vZnplNRhfpC7/XImu95hqBMuMaTK0rDoIvyiY1/xXYffdVURbb7/AJa3
S635KHgqKIy1Phai4J32FP0JGHXr2ETXoPDomAX38qdoxuN2On6cCi2O+6fh
GHO9FegYW6RKy+zaxHvuIqHDs3gWhSmfMefpIQ5Nnx7u5GrqOpiguvaay04j
WmygJEXKHRjzXOWPiO2yIhiQazsG21rDZiXaqOGRftQk5gXBZf3y++mFMpTg
s2okL3vkyIgg9Oll8Ga47I7DmHpDz7pfSJoa9s0kKv3L7QA3Ddc5R5DVQ/Wd
j+l2cqt8FM3nQl+D3qX97ogWHuSMh8UE9WAdI62KLoMzpWCX6zAgvqs60Ev6
GxWOOZvaQoYhvgvwWSvPQ0YWVY8tjezPTkUpnQQjZ4TW5d+BGMmdYEf/qk3L
rBEAbvhfDPP4IK1tkthfnzI8qg984FyzGR77Oph5fzVjwl9uq7/ny9eysiPD
JAt/9dkE4lWuSgzaH1iTolNOiyABcWsNSHLgWIL2rPBbltvhHb8E3DinuL7+
ocGNS/InkZLAmJ+shFJjben92dUWest1mbZ7Oh0+aqZLCLIvAAi7VpotlBZP
SG0y5rmDafEPH4Mb5YRg0iT9P6BM5HP3J2Kxd6jKHSaEyXL+FlPS7Cr78Cn9
wgusA6tYjH4OoiQhnYBo3/Z1wJMzuTNIvkKvKHTnauALNcmYkjUgTqs45qQi
GyCZ1WrdNE7kbfMjdkFU2yu9KGJYu+nSnb86Aezm38LBkhe3rRjlOtTtnHzv
tjrMBCqXxK9+4o+tFnuDa25ORygozXWG4v7EKs6I0yFGLTi7VdFeJhcL7VIq
zt0E4vtfbnOdXuGnAhRsk8Ad7cmuplR8mGfdV2zCmeIk0T+KewNKg6JZc7r3
Lut5xvpSMWwCh0gZ71Uedcl1cVp1ldPefB8PiI0W/CcjPwzsh+4m7ERJJzZ1
z0qzjOvDYuhjWU3dUSDE+pKUzuAyOkwrAOTjS4ttkc+aZicKksl7ZcKKD4vZ
GcOXpaXatj5Flz1Xg1lroXj+V8MjJZxdm8f9YnGBCYl8nE1glPTlvkN6ws2W
VGyUvvCz3tvR5x76zBbC068w/fJxJP1RtH6k9seOiveUcrI0Vg/MPsWGB+uk
r3hyDt01ee4Yu6h1U3HFA5LkyQovUyUhaVJjTnSgiruvB7Snmfc4fnYPzpSY
70YUZoEHsnTD3sn76LedAhqMppGfWkaiFmeeNSBJIC5MwVXw4K/zABvVbGdh
EmTFEQXD6hnT0qd1cfHFMx6u//yY/kNI2i2Sb+LKnxt5Jy0/M7/aXOWCUULB
fkubgk6XQFNeiJvw4f6lVPUDnxA0XECaLUh+QdynWfWPd18JvACIdiyfP474
YvUps74DR2ym9+utsQqy9EuC9vhEqOI0sW4DzrOJye3vtOHvDFPB40aNykJc
buOxeCOMAJZMBrxmurIejdn335iRhHLDHhhyIl1xl14dOqUUR/RyhwrmPzTi
IDx+vv9SleJ7SXK3mi97oZaNScpD5tDfPVdmGfF3asg0CW/s4qVuvKvBjpWu
wbqc3bUtTGg3Eq1bNNK4PW5XJa8ist2G5eGqsbTyURYLzoUHf998hNZQtqrf
iy77TOdgakVMIZx2yTITkjbBbKbScgxq8QuoOGprKQO5Rm1pqG1xlrdNf1RQ
9tNQm0xDTbAzP606EAEy6XdNZUDREdjCVeEEgViKq1Ltzc9bw2fdKTqd/jtX
0jsljUsTHsmfn5ff0ok4LcAvBwkbF2PohCCRtorqdACPJA6Sirg/n5tQny7U
BNgExRmmDUTW23QwL6c72YKApE/yZHGcLSpzaWK7iTYoW/ti+WRA6fEEOg7Q
9rFCNocv+5eCF+eYh4CFz7yMvlvKmH2XfF8YJx7tZIgf9SXphvNOqlT85tVq
IXJR4jE89+k7t/Zr+VG+Y+HBAi89bDk+rwLs7epxpyp3xmri5rc7ww3Zx+W0
YtkDSUldHcfwcU349xnI9uJr9c/l83bJx61rD0tIntjj8NhZKAQbK4aM3FVD
qaaBiqSruXGhAqNwK9gpt8HMy4DvKUSeLcHPmHGaXGK2nrUhudKavsKgeaVP
eHWwNY1K3x4VgqkKUR+tnMWzvHVgZIb3PjXlGXjtLe0CJ3rW6OP05VrAfPGj
bNMVFU6PitMChjtirxEY2keZOW8ZoqZ9W+wuSGrKDtp8kago2L34NcobASPc
2i0Sz8hvfwca7rDdDAB2rynqPgZWTXDXqgI5jo18RwliTX4Q67fgIcowH1/U
iqWQcQ7+fkB01x8mtW0BzdGKBCsVfGwcUI02yIdrpoOBZP880jjkzdtR877f
7VjwuaxlJ1BW20fnrU0f1bXab6axvdXBRWAF3QudbNK3urdyebtiduGhPjaX
32W1V7CNBdi6QwavDHfHSJM2I+D73IDqnDyroU2Yq9Xk6Mjy8Xgv1jT6rKYD
C6EA5Xqg92a3Ab/248vAVedjXqfgryjJ9H+a858ZMcJhQ6PhLtU9ViwkUglP
Le2DiDZXsG03HhJlOp1vOWRlMXMkKP/iR+Ha0xuKHI8BaE/4vvuHgKfnUteP
omY719rG/7aE4DQ1N4oT8ZJDWomWq9E6gkKPgv8cQNVI5uDsnPGzngUfNNO7
bkQR7czrdHkbe0VTpfjhVMXh7oP1Ws2H51ZHs8EZcO1bPvZfSmn8QIKUDbYL
UmbJ6wZNiK9sUVSTMyysH3XpIUiYrfcqbc5rRxgPc+kr/rCUjX/Hol1+qGX0
kdOc8L9PU+WVUG5APIZzR7MURu3mJcd8PjNYUMAyKeo0I1xhrIivcGYlLEQ7
dyMpqQAFMMthKJY8cUnOx8xkSPAvot2aiGt3m2fRe+xsK9jyP9uA5l71JtPk
vqtRJVsIzDNtJuH9Nc9lG4dElL2b180wAlHNuRUOl3ng9YvFVcUfyFYciIbe
fStpA1BBycG0hg99d10pin1PB9pvGSbFfBaSEbklMzUvmaVBan38J6dGzNMs
0O50CU7GaKAUWyjc5fvwg0hJ2cK9HCr9QcBoqryqtAKYqhdzbDLV1WxIYRYf
VJJVS+JPh4FSsgnmlVzK54cPqJs/hF7Ijs7d2Yxqzo0mG9eHj+g7lhcJfvWs
H033/0KNJ5T3nQ5BrYBxBBqAqWjYZTrvaEaRXU53HvIbazT/cOtsUbrdqcmh
MhGxh1Z+MO9UqOFNxLmdXqETqB9cljh8fIIoQ7bp6z+tZRNfY5fxG6dZbr3w
3hPlwK2ACnYV287neJkSV7inlZaZrFVUi5edoRqYG6KV0sIrdnQVq1d7A+jQ
5oZH/F45Q9l2ZuZciVNgwjFoFCzpTjna6bKYf9SmJzm5mozDk6rjpYrhEWWq
tLpo0mdtWYWt0IVJNyAtWCxuSKv5fepBAGOtstVTcm+n6HRjisTAGe/mTaI4
+PGak+hHGnTgsKgG+qspc4ZIaYhgb1PpNc48iolqDk6BzDXA0m3iCXME3eFj
jjKzA3cYTaE7d5WXw4pzheA+k9oOZ3Y0mD3WAPUHJBYhwQHCPxJIKzhixoTV
fodJ9Y1hARELGj065o7QBR8dRwpXzjeFhF6tzA04zGqTuPC8/+0nkUScK5/u
/VF0dEV0UFhyqASKUANkb0N+FVjCU2jMlD81fV4Mepo1+erDYrAbywmb2sXL
BbCoBKrM1u6458On4BpLrZqHNrHTJk5nip+8CknfxWpeWKclacDpcACpuPT/
wmI16AiBojPPuqMlqsSrf9fSKkNFcX/9F46QuHpJaXTtP+vXjIvB9BsmKJNM
qJYxmaFGB9GdLuY7Prrfub1cOKuQu9wvGzaGXlwoU5M2Eyo8y6hjyS4cI6vN
3VgOxwLqLaog2H4VOVVfKzKyTljawug7my27c8eX0JPxhsCmSxd1QxPmCoCe
yrgsPz+mKrl0nlHhzuZKsd/y9Gn6jpq2NNqPsCdBmaRDbuLnZKWPCrExbc50
KtErZZF//kaUsap6sYb7f7LChUTjKZMITJN9Th2yVou6/JsO8cKulr5XSftj
PC1ky5EDXjtdqQqMnpqCYiOkm5m1OPMGpsHBixM9Q3ph6UPMaGv5wQBtoTfp
2TGY2IZ2pTOi5toeO82LkKvhuZGYK7VbNghMkLZ7qrS1insV94D/O6gS5yKC
iO7ruXrZxHawzx9OHdPWimkp1hitVtq7168m5sO8BkFTyhtB8yWpwx791WVk
FEFdIChbG/RNF2KyUg1D7ij5IxeHrVZZ1GoSPbg3XRMKJL3JeKI/cyPTJwHw
R6zNg4sOVNmw7T7BfgqkVAvhRxlr848EOJvr2JMBIiigf9JeTSgHYjL/RZMm
TGoRwz1wqK8LRsTq1HeY7vND3uknNHABc4IBrVc+/9gCfPSXrULEjGT0NooN
L/TZ2XPRthxUaJYXcjnaV+Pp6ZsOqz+g8uedL8zjhALBEQNBHQSo5SLWgaV1
2Wz76Mkp+/BYLR9mPAWd/PW/MODGzDkrBmAO5UN4TiSkqXn51e4gvR+/17xi
KeGcQ/SAP7UpfcGzcdxKsBQ+sHTxUmVgqI6MaZwm1VwAr4TqNLQ51Cwf8+qd
Fkn0svMhwDgFA5QqDpTF2cHMQ0dsYB5z1YImHayJP+h12V/ZgJYckwjjE1FQ
BHjuB5mtfUqaI5fzM6lbf7Ea7sGWPjIdF4d5g02h656xtFYAqiab8pK+2J+B
t2B4M8DGa5wKZLNXLpnAlHb6TMN4AydwIaMfnM4vZb5bzhzBEZr/TpxJwD+N
Rhs5jktTDPzvPuyDmpMAFanzcmThLG57WZwHGZPcXdmXqH9Igc4/jnSpMUE+
4YaxlIeH1HwZk/HqFWO3r1HwDZyaZx36l5UGmzIBDVFISUIobQlWfB0HCKdV
/r7qzoGkSvZcnUYy9NcgHhxUCgyeOjN6xnKUjARvKvvREpzIQlggGQAHy+aB
8XUxMDpNR/cFGgJxihX81YeHpISmEWDI7RjfnVLJz/IzSRTumsgaSM/LBYtq
+FPVoEunac04v018AtcX6gG+dcgHpfzog1A85LGhKhtwkRWIOMtv+HD+ugBr
Lg++I0890Qaa2Saoabh1giE3Q4NGxsuFCOadbm2BqBvJUgjnD/15edxdNHhM
GhzuhgfaFI0A55mfC5OY9uSjXzzEyUSLozQq+qbDH2etzJZlebseCcRyHTw7
zyRejLx0DQ9x/KgqoUFhZ3BSX2vms/WQSnTaaoItSYb+zsd8rp4mzvN/d69J
AibGHrRQMgqOxECyPqfmIWjlwsQzhXgOU6iW+o4WY2TKI1rYtg/K8lPtotVs
MajfYl8BCRQMXmaiQn2P+VYQpsTODYq958vZHqpoCR1tASQzz311VVAftLVh
26SiNulgyA8IJhEHM6MksQnIHizCzQwpTUCTKR+NWNvRi+t9BO9Qy1+LOec0
9JSJdkqISbv8nhLPZDKA/jchKW83y6s4xo2jGi1SG/WKGoTC+B1glmwvC/Uk
DMqECvxNaBZJuu10IY2jpsRQnNrGNst+sBjEX+27yaFERB3nTdBM3Wgz5EFo
vcfvlFisyvXFzJe58AgLKNodmo4pBAT/g9grcb+CmfLWCb3bmYi+bkWxeuTC
eQALstbt+4sAdaYVAgUdcl0oQ2t+vc83YrruJap8X7dOLnFqC5SWo0vid5Tw
o2fLhfydT3goebWe1KLjHpIsE4egbcboYYu5b+suLN7KvGOQY3CDRZ0vnTQl
kPF9cXKQZuNXFq9MEpyBhgHcc16uCIWWNKSfCpuKkAXo0Q9gKMY6GnRtAUkH
JSP1IgPNe2QGmsr4/csX0SiZ6ny2b6e56Qsm9D1h+sqUPPxnwulCMCB2FC8D
lAkNpkjmGXxMxPlxeLNGVTSLsHLlh6NQs+DCV6fGkuutWZd2+p0lgmq2arlo
DgzPPpD6PyiYWMOSSu6VkK4t+RY5FAhv1jm2uADz3upCgwOsGkBR63vFJxGu
73aJuN/D3oCPNiCyaCSTt2Y1OshQj9Sin8x1pBC5VVLK6YTpzSJLBYPgSk7+
IoDAEk1PVQHmULSbTQ/PKwKWTC1S9ECVz6qeyG3p/7+2cNtJp85rp/mi1TvL
mbX8i3HVY+k3m0fmL+mATv3D7l2JQqmBGvI+2emppuF9xBRc/Hs9ApdzUnbQ
eHa8lDxT2szLMcUtvuPfj4ybNzR0euYfjPdf/umn4TYzKAHoM5oV8T/0A5Rx
8MnAv8W2gg7+fOFNDQwWtqFxxpPGXlhXIXW8d13bY5jad7wksbttyu0f+5g0
mG6Kt0CcMZ+2FgA9q+kdRfccKbn47WmuhFKdpOTdPgvDHKI4P3xxpfdg3xzr
qt+iCSNW5TbNYq7l6IQe+Q2L5YKTk5EbD+cFgLEsZCSacYHMAgbDF18iMGhm
k/t16W404gYHbXuU/Z7ZlLOlUsRSsnc3nhtMPMzYZ4A/P4rsRi+yaHnbU5s4
zVvEWCCCH327l+zwb8KsvsqSkW4PGa1u4L+WN4kZcglQEXvIVq5FfeNYXYsa
LcIMZpHldsInZuCcxKa4TudDeE1ESEcny6Zz+myWD0P5Zzs/sv3mMxTFM332
QGTJSBy275KwmDsJhmm53QCKR6K+fqOTRScn/gIHQqtJNB6Tf+JHN4/+136r
MoImxFXkpXlYZ7Dm9kf9mgTMQWvx1rfL4wIn6kaycpVCdj012fz81cBjXMF4
OnnAD3PejGvf3Hb0zSzY4+Owcnvrsm/7Q3xDC4mlgh1pMH8saKp3IxiEJXoi
IyzUlX8i4o8McuKpmQ0zljGvttZF2MG5NZFDs9fPwAeLOsJ7iNEve3INtaxU
x9B16eiRJJGO2pDK8gsJ4gHyg/pBGIhyPvVlBLzocdz0eJpHOayuq9JXEhMw
pF78HMVJ12YUwVlTtf7AuQMyNoxtpsw2GorlWlFXWRdu6wy4AX+2rwpQf6LO
KmVoUbwtBlkXspVSvhiEwf8HeYx3120GDtzmku2UQ0whLyMGTaHFzxrsxfcp
T8rUmaTC8kuA4ba1BDHzUscnoHnwx6XoF0qzB+6syvt6UTBTv64IxlSajc7+
m/XMRT8WMSw7y6mQFHn+xFrCiN+UQ9Oxa/apqiFjgujnDGdGC4Org5n7ZXdS
n35X5inOAmNdG3stn3ERJvSOn/Y9mdXa6Hod/V/vgvlTLbO37+vPvuVCvcyV
IjZ1ZPotiK+kFR303f++u4eEpL6+gBE0vrFmk6KnIgjjUd5viRA5sQZO1fS3
tedJSPLHFrgQSDFh8bkLQ4LGAG7vo+11cMDnAVwgDG9NZfLseSGErurezKkl
PEXSmfSX0IASl8g1CTMN3TlWpSX0+TwVaPxe0qfUvfhR8x1Dx9JZgQZqkV3Z
OPaZ5PFnLDyO0CtEWWZxXAYzylT297qyGf8XUBO/ftiJ5xf4UPOnpsPQHxTk
DVT9ZqkXyC+RCYAAqhM/sxArb7iswgIYt2SzRR736CAvEyF1HHSJ/lMfb043
qiKQiMPg33pcOfaMX32aNdzWvxeIoclNeFlpk40mTKxOe8MKz+jdGPeMDg6I
HLfKX1t291hbUbjxEQLlRNW9cDqY6LaLbPfHkN3qsmU22UfSPI9PT9gXJrLA
xFAfhuZvAu/GjAMICZFAX7Ep1mUsuBtCpqLD02C6c3ZgOx5v0tW9kk6WT3ne
ot7IY2Mrt7n67Jo1am2GmDT2BfVpRPASEHNg3eO/An3rZWJOcc8SsaRp9Rf+
MmJEAgwXVO6iteOzzsbRtxJxyz4Tnc/mKtvQxfr43EbqLSlQg5rnStId4TDH
2tnDto2YrExdt3teabdKJ3mT9FBlPqqJMnOHW523zhVLxvkhThMVQy2PNT/x
YRaQNxDVTKnuaSZwkLQAJSwdRNiwlRS+uM5MyREDeW/sI2Z6cPtLJpMQBKys
+bNAGiZOlzbj7PELNC8SLeqwGP0tZc5906SC6eWXl+o97RGkvGzfwh4b4c6H
sOu0wqQiPsnpZD1g63xGWAHjbGK+c3HdIXYISrMn9rC4GltkeJ1X6rBLX9VH
tAbzHA/J+eqGBgoxYKPEAcssC5QPc5NbX7AddHa7zPWIyclol4mmp+gsAT8/
PypnmHflEb/D1Pci0Fo5tKe6qcTPmV3feBg6ukeuPNdda7YA7Uq5phXdNjan
kW6nCb8ZvYFLRzhDH9viorVHORJL5k681sz+xAArvjcqOWEI99ABA3EE9FRG
MpPdTZ2UVRQlh4DsdeyyhH/GejRablJDv0Aj/o2lHHr5+A7yIciwv6QrfLy2
8C1Dsl5vUQipSiJ5nt9ySgkx7P/Ow8UPCAw+8QJ13J/oGvELGWw/9pnz73m1
2doSq4OMjKBCEO18k2PUCX5Wu25dQrVMT0wkonv1YhtZcyWDwhlK6Bfvn2Oi
kXx3ny93k20BU8p/2rFQHXzR6f1uwqOUjCzjmuIi8OvlEslLc/IdoyxMRhPr
sMJOUjgv7DHiAF6sScNB+Q8rkUqoFOjHHCGxT6IcD7Xl2MfKDMm+TxQ1Rz66
VifXJrpSQRsaYW54JuqIIDbMTBjBJyU59jBoQDwAywIziz9ascYsUhjiAOBo
rWG5WHcoxO184IMlfEQDBXuXSnveEZ+fFZ/iYElc+n7/5JEybAdogUxtuYBI
65PMgsD8PNBHMMbPEDlF5AUOHwdxWwzcaE7gYgPZZaIU16CpeWs5/aO7DdUw
jyMmL6q/t7MumbCjaLgSeRGgmFj4T2jZSm7IoPShTn8z2o2qnR6/IfO0jkd9
DSh1JuJq7husd7/tTHBChSoDT6xAZm6wHdJTb8ufxSl33b0LZvoBGLNU6Kk+
/XsaVu/A7zMPJRRdVC32m6DmkGiAb9XUT2uoKTMuYTN9/54J0XUX4hxFFmHg
8JzpWBVvg1MyvwEuzOdYv7yA11ax39wOKv3bO1MFiR3/2NFa1P5Al+aAjQE9
UkDJ8w2HSfiNUoT5R/3GYYYREacdLcskc9yYt83chC7eGCKpp7h3EASLmdb7
i9cflS1Punhs167AAkIjcuqy/DZCKy2V9Ira1I5aF3YlJNf4lsTUlswDeTFE
j/pRmmTITlwv1taHGoeimoHMrNpE1GyQVnVfjkEF/Z9MPPPqu+jFUq6f/V2R
Ow3F9bD/EC0t6v6eiSJ2YFeCTNtE5nij3nxhU4faIvSn+fFtXmjWVhsVvIzf
HROJyWsQ3AR1axMYERh0nGGAiGwjle4QL89vZShm15iISzTRV1AwNQSYDyxj
7IYWZHo049ut4Vganeeo9bmLRmQXFklTMIScktYhAFC+/NNAWWLJpUFMWIkO
kccFIu3BokLClZoz0f046N7ZmCQTrTSy3OnQkGNS89qgqMT8fCit/OFb1xay
LvMtStBijmfXuaVb6OeSmCGsYm/XwD1b4ZWBJJgftLtZrYpg6Z3Cy9FFtfj8
NpnY5OsGJcoU1RTlcaUgaSdtt6BwjBcc9Dsy4+AsYIBTsQRmuCjMXMmoBVRI
3sMklS/NmxQ9B1Sy3pyv9drapemrVrolo7/Us5yD5AvI2ATD1j2uWKRqkU5o
RevTXC9O/s1J8jWrkkuH3mWazcn+z1AD/IYlKl7o3jeBw+A0bBq+psoRmHRG
nddswCl/oq2h4DHC7M5Oob0z8grsFrVLaUNU/HxEpVqKlF0JbRewBfNG566/
p5OxETnulZstx5asVRmT/32GuMlpCFs7XnntkOa9TKI3hozSfNu/hOQ5uYth
g+SQSKmP0C+OILmXhlCFf37gp9p9jk73tM5m2WnOFPf7Xu/Rxhg9TtKG4EGq
ai1t+SvBiaYS1BbqVNQb71JHC9FhHHInmvLrw6y/A8TIzTCuq3WBnRDAvpPj
ZnNw2qTBQJay89z8HRX2tIGrzQULVCTpMLnkMW6v6hy1qDyJ6ytxRvSUe/h0
yWsWiaRCYpkdE5V7m5G8hHuR3+aT18GhqYXJ4HVUda0vswC9m34sOEPW/P/X
beBj8E6J2T5podh4xKcJmen75SvInMPdfWdL3sneQBcdeWlQZdOiJIAUVHWw
AKUi8Jmqe+qJHJNoOYE6WMlIznN0j7hXRlH+sNhV+XHLEA/hMq/2bGTtqfas
nTd70U9WrqYL/VLyisK+l7ur9CLIfvIWzR82twRaGlfG472DdGHG1oHKszks
WpLnT9m7Tbxh7xKJ94sbScKXHeMF6gbkyij5YghxhwEVA7fh1CMqW+YN4vQ/
99BdQjs0xtFAVfNgZTPFi35PQbiR50IBSFRdQarkrNbQDBo+MAKMqv5LVcXf
CV8z0a0+2HBdv/nNr8zXTwWkfjEysUuSGE0AMPTNPHX+oUcEvLDfnE68cEJL
8AVmpoVWll328ChQqiFggUzmVsjnniGN6u12KXfceMEY4QUsQO5MPvz7Ws5t
MkqTDBsm2f6hyF9RlpbAG1P/KGs6YqWh/hvVybbkyy/8Nz9+YMjwE4tJdxWL
KEzf9dSr1jHRLpin+WJ6cgZiwG4/7YEKq0nMB8yDaCdsv6O3kZJpFSOsbCLS
wZ5//ASCxwsH8PiviV+rKcDijjxX6QPhoKByGAR5472LElY8sAewjWxZF7LD
fftHSIoNfq7wZ52ZyeGYQDTJ7jP/8v26c9BVWdH2VWoABe4Pz6DbRapCaWHE
sJ4s2dYGre2BJY/AILnVjO/z+zQjbdB0fBAKJtfefhtppS/+cLc9dhdAJ4OA
ZZAtUzcAfV4W/k5TKK9RCJcC8PDnpodoxtvw8WyhaE2seZvQfPrZiAsDczJQ
uwvq70ewLlCEtWxt7rmMZmb5RySyUZPBFY26B0WnGUphAjTj3l9+X06ZYE+D
E1RLIyC0qQyupW+X/HiCTsvsudHfvs4P3C9SXG6c0O60uFL/kt3HW3HB4Asr
y1wjb2Ju/yUTYakHI07+wvqPbSTjg02N0uMIsicMpI4pyxu/x53qGV4yIe2u
ofUYI/B9DrCQ9sN9IMcoqGQC8wT6HxVnBXxCHLJQZBJurauRrVhRfP5ClnsJ
e6HEcd2c/2+A3kzyRcckpYO/Vo98S0Cr9T+nNz5xnzKQa0Sguf7z6WRtepk0
qfaHfJC8a/+n0lexDn/YBUJixq7Iu/058kFBOUaqEpJQYe75Snu/i/qcJQYJ
AYzslQ7BYovPBOlznmE6z+y5SFkWQ9v6/CGAa9QQmBLf6V0P7YesA93rCD46
aBkBaE0LAsi/WSU/xu5nop/3k2bzyKGJOkDokJ24Cpu7Z7rEw97YSU6mgRCM
pmYTwODVOkThXMTj3tNklyHu5drxoqwEt+UdTtyi0TQH3ftWP5yL2+F2W/8E
8BkaIQyWor9XLiXNP5jrgTd4K+dW+W78TkhMHDysr9lLzsV9QzSycm7e09Vc
kn4uRw3XIefzD/3dNrxafbLQic+AlLfS5tKF3mUONr+SxB2qfzb9CkuzqcPe
lvrDvs5JOlCS7UBK1BTdNmY1t4FMjR4Naio2glB58Q+bAUlw3KB0QMp2BB0n
1urNb5OPXz2Ulkum0yCTb+d6/OMS0dSAr871FTelUhL0ZcP+yeX/d09ci002
0CyB6OpDB5/uiLmxdFAv1Cah7AABz1W23N5xDA4O7xiSRvlr0B9EbFAKf458
5nnCkxZ3xY/0gAIAphDEvIxeScQIR4gbR/ogdokgIOmo0V0HUde0QQdKFWRC
PHTO9QZzTJFSh5XOY0HXtoLUGVGD1IUvefexOkqqo7xIywe6Lc5CbJD9JChK
5mdcVn6ImePFvdoGfbpAupHFYDlMVwhEkZ6qOR1KnSyCmpyKYnptJuutGamL
nNZWisHHP4/V6DZqmxvawr9KbVm0XtAwI+R59XQ0uajdnLMU1EjrWfUl6cKD
zR6/iNgor03MDGjvYeRbjy2mcMmHpjTYujhXuZ9TbbHKTcPrf2+EhqeFBAjO
yqLLT0g002drSMpqg/xkh/PdedpxJxwL+ShMWLp5IHlLNoQT3+7PuuWfuIxp
QMJMK1l5luFAMnlyssJnSUn7YRcL3/nxfEK/Z664i+8FZLDARsHOc+hPcPjV
ekj4DwJ7uHYrEHLAH7ZJ1z6ozKA26zIMyCTkO2xiJJx1ZQDq6rDZl3fa84bs
bWjtB58oB9/BHURuUYBb+0iOSO184h8AzUaSllFVKILXbYkW8jwSzXMWgJe1
buq/++w3oNY1/Oy7GTrQtaqbMAwtq77jeQZJla0Kft6WMFwN7svgXcytu9lA
+5NMaEBstVCzmXb4xVXrNbAJ0aOWwyp+h1I2bvzVaJQVVULlR+B9NRRR+HNA
LjwQzseynVt+Mk9wtAoEz8YWPOrwVpugN6NuR7y4ZDC3f43zBkeKwKCsrXsZ
f0LWk1arzIidhNeGDkDxoJ0VL3cUJaDzMPAThsxOYn4PJSRwuYQcqW8Dj9kc
cYW9xk3yeDxa1IQwsCXJkSkxXaKUNb3Kq3d8ToNwcTQveQ1+M3NRn/Q3HBX7
iB78JaJOoIJUXnmiWJyzN5X6CbRg0amyci0RbVyDJ7JOrMTJIoaRfrJVPRmY
Wvbpa9gYdgihHQBD5Sl9H2VkSMDIRoay1aEdEEgOmBR0R1VbamV0MEyBwmrE
kfj8xNArtBUlI0dcKpuaboVl+q/WWVE2V18RNRtaRHu8gDD5t7uaYwt/ERlx
jHV9Bu4pVQexbZ9xlw9hivZojbIG3aJnPeOaL/zvmXUTgRrFU8anXzcNP4fB
g+RVpgFWhR7jfekmEMsxVvT8Cn6VF2WuuRoy+75w6f4/XBDrWKuInTA8JJxx
tv6p4QOPRHhwLKoov3NFkgFwhpiYvuF3pLc8qwd6Jcls2WDeFeiE4nPZ/KmT
HLEsCOXKwWHS0Bkk2df789Br54byKmrygSkS/YgJVEdBNUtWRgBnvRGODhJ8
XY5la2IMS6mGLDy8/85vZaNn3rr4VXG0j3lYA0thPdJGb6oR4EdsC5HJ9YWK
FI/GlMWr/xMcYf7YPfB7YKsGqDlB5ggFLYJHsSAlBUmhhD86a/o4lzqPHa1p
Ctl+Od4diitXzYaR+cYBzBf53v/uE4KnuQk6FhMuyO0F7wZqo0/qxxeTaoDP
HvtaIDmXdYX7u9MooRWsb8zY9/j3WuF0Xfw0xp1BEdmI6OOMqYqXZlb/7qyd
JgoVZWXwBbIA+bsOjDkZfVVnQE2+EfczRK1BtcLzM80LEL/UB6EP+vawS+3D
BWxM/K0aIVseeYZWr6uveFNYeO5oubGXHlw05q2TZ/84MJjos1NCmW3roSu1
8Yrg82xpQhYBji6MO5+5CebuhWLiNn/TFPPkrYeO/849B7+FR+g8yEpPoE1q
2zJwHQHwMRH+VZb2G+/TRB9Bu/jVK4YA8I0WpSDLrp8N9tUk/VyDOoP7wcyf
TtW3B/qPgk29KRYR/M9tvQ74jcUhBOR+wFLWJhLx94XC6DwxGI6PRZAat6cM
DcG0T7tc1fpMPTaUK8gLKVoBiUG53tD4qt9bHgBK9oZ6urDiKF1sz8rZvz6e
rGQpwdHAFwvOQZrWD8JceIa3CGdkVolsnn66AYNndsfY+YIkUiX3A7Mrao67
lp//LdOJzupSSJLDnWKBHwhFlRy6yal1XG102hZ+/jug/6JuiEV+XimQt4Zg
8d2mFpaUnA5WaSUpJgHO1pJf3aWao4Xjj6nMQLK48EMNWHPGcLSNTf53OBK0
EaZ+eFetc9ggDAq1ObK24Nl3yk0upmRHpjmoj2lKcgrmGbjaHlQOpf7mxd8A
tVsIjcXzKjXVl/mZY+h5PbMazv6KXJ15pgSvaOMLxaO4rfkHWt3rwfdXuUF5
3pETPpEakaLeNDiUg2qHgVrqByRDfj9Y43xSyfX6okqImzVKR4mkl6u3Q/aT
xxvGb2QTkIP1Kbj3/GQzABrIGNux9f26LvdBOB4OyeiGJ4h6zooQVijOvO9j
hv8xehKrSOVUR0IENFCz6z4zw1d4JBsLDrF3FBP7DeNEZjdVhRD48VnSUfkB
RoiZTHeQId/dETRZ13ffgEqRtEhw3z9aKqI2Z+4sUGICU/OhPv7X1zqg/2o3
bwoSfhbiD0bSQb8B8bqo+/och3UKW43VkXPcUKMnEutAPXgy7CY8yOWot5DC
Hk69IgCTu2aJbYg776GkyQBTE3D0TNjAkpPnUr/o4P6k/fSKwj1+xm8Wkm41
8Wj1vLaewGHfIUfQeFJwEUfzmYcCa/w5qHuxpTCC3v+4vjd17j2tVzF5+/is
KlW2LhMt8j3G6DgNlQH4POHbd2CYOH+pBmaBO3NS1BxFtVg0n1K/r+LeuLZ/
/Wty1tFXfb7S3O8YzqKfUPIM1n8w+8EbskSUUGcph3cg2Xb0jnFkQnHOKpax
XU2vjnWMvM49rgj10Z2TVoXgkCwNMa53PNvs/0OCNlhzbytUJhJr4Qn0JcKJ
VzyN6vv1N/pOpt19nhdNEE3a4rjKBVOXPYsRBoIjvMM8kUan3NY1aQ/wFx7z
zIj7L5ZCG9qyEM27jJDfmyRxQ8FUs34EjG4zwSRTNbAgZopDnzMbkNTJcUE0
V/mkzvNAv3K3B3QL1yKqc+HCs/W3rnXiJBoq+zo8tFN0YqYFXodnG+yl04w6
gNuRAPlINfEknFTsY5O+adphWt9xRwXG+kGyv35G

`pragma protect end_protected
