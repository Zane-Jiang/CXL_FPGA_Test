// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qOGPk74bRHdM+oSlEUvlvGG4oZA0Y3DWKlVc3qk4lWj7ceV2HTh9uE4Ae8Uh
S1hWb0m6tvu42ebxuWSGSnfbuxuZO3xAU3IiDLzxncmDwPBsI/nM35qPgx3b
gz+6LjqlkeDiixmDeGPhHq/2HyC4/pVWETos5BXXWX0RESqcrROmQJUY6BLL
kKw9GSRcpky1kcMS0BJybml81RhphlcfXl6qR0jo3z8sZeettp1n7nqD5cfX
f2JmNBIwKKyrFoOmmVZsoBWlLz5PrMWDpCgFWc6Z8y3VzgJxvI+xVGz+74RG
aYRCaduARpBfmAYQWJ7QIfBO01OULKz6NCnun2Pr7Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nieboSjr+m40PR7/McOPSqOX1393qAHGU+0j9XIJ5wWq91/7Ft+p7ElKhP6H
0HLhKq5DM82I7LDmAuQQwUlVnUfZaaTCJcYBdT58VjsCU35xMPhmsGGP7hOc
eaTg2HOvknnuzh1RKzWcZk+K4bgiUUXOwtG7Ndx3dK4UZ6pwkey6jA9RIlOV
O4W5Bk7ktusvXXif+86A1uf3qBFofOFx6WVoWoBuTUw7vezzKna2Ry3lQ81P
zQj/7iWdGB6aa3Cn5gYSFy55tZ3Oit/n285bKP7xF58DXgLdw5XojBPZ3lDo
qYOMQ1t5QHjNa0IaZLD7bwxNcrKHxhRbXE9eL72Ltw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fTRyfh7xKs/VFKRFIeMThKC70M6p2pNTNOP58JUuMGswsKi/hlj2FMPQt3in
c3HLOHfOFCiDh2UTYtjC5kQkRxmULHfgqPTclOaMfwc5HurunxNSNp4X/NL8
5SrSfRPuR/AycsO4hHiVw7+y8YHreWaJhScwfN5znn7FX+cGfdrtqu8n3cly
O4cKWveqahVRfadVb61pMY3KYpXgvmyk4uJAUMjs6b4m/Ts6xgJ8PA+sXqyh
5ph4pxol8OSxTNisNaFPsOESfgLItfQlT3+jkujJLYisVG4OMsse4R880rTl
XfBj7BwuwW5Irb3lxC4D0J5q7gvaGyLK361fzeDu7w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WPT+PKEGHF1lhLGWvHcPocIKnqNJyLWnL8NrFndyE+ItMOi8ZRRb14yKAQr5
fGYvz0Zt/f61nxPvocL6dGhc4giS9SFxFhxuAdUibl2aLRx5MRNVU6ofuA5S
Lh+NGlVZJcGPRbhfzwOGkkuyoQkstuwZ9tYXaXRcKnJfvmfXqaY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XgS8zYMJSR7BSfVEZWWFkSg2M+E1S3rUrihQyMgGpOhCfBM32pK74UMlyhA/
TJb8bEHeAxbSsPCzwXjKVHpIUqHlqjFuACSFmmpODjeg92uk8Qp9JoND797e
1rc7AnJDuqvgpt9/mt4hgj4ppaldLerkz9JayIA52xx2W9DRcXJuckMrxTco
FdKa1sCRm2/CN2NuOqH6/xIt9FcNvLkLliSYPIO6Jo+EbxvaLtbD4pEDfyC0
2wRLBvs6aN8dQrNF7JFiESs+vJqffqlElchlzy35jiUUlldWkhIQ4q82/KSo
TbFz98WTekakBAkRh64zhv6cNTrblJA3G8ORbo+UIv8KAeH6kB8378nB1eab
uod6QlzPyB5AJcIMT2Vq6tF7kFleEjP7hwVHRy60oeXoqYdRhz9rezhT248O
SjZvnDK1mPLb+/OKFTD8GcINWzbiPQVl1wOcajRQrndfK3LxNkRfxnW8JYYg
RiGk1FnUNpJH0ITIsIcXxa+XZu3b5Vuw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i3cXBzpxhWZTACuArfRA99REcYWLqN4RL/qq+f7Lv2yKypaIe71kKvt2yKA3
phkFGZCecWwkV8UInjaAmdBPHo4dBGkdB/aCSr+aNbWQcIyLF9y/hp6UTxXV
4AB6O0ZygxQHB7tCC7u8SgjtXcjlmQXm9/1nTQjSws7n74bLrSY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zhm0QTre45nr0xkC+jMh9OrsJ/Su7VdhC2Fa2WnW8hoJYTGpSr4ZUlenDURG
p7HUQB98wgAS/+CiJ1DE0dXcRKzkwaxJFL8L4/8dwRDzKH8TuwE3prayE5eJ
YQjgovNstGzacpxrjczLql160SU2S+v7U+CcBNOys8+QZ4V0atY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
FCt1x11WiafdqOxNgQh+MawcW3V/xaI/xrr63w026WlzYc5Gxu9Va6edeJPG
85qj5SK2SBTUzIWCLn2aA8XiGQ9M8+3MzJOORaLtNeaXBMVAkOjpT873ZJwK
BIAN1zq4JkzEhJlU1PGG1UvUiZcMSpGoR6l/jzzamqWMb32mGjDLA5vTpCU8
eaWyeZPF0Mijpl37Ici7Kw78vTsdO+H6hT4BztpsB2tTLSSlS96ud2Ck4SLB
Lol1RxGL9Cycc5MJJT4BN2BYO+D6IbXlnP5WkS8PnEhqbvYBIhImqVD9N0MK
ZqkYMRMYvAo85ijxLmhRUIFJ15LG71l6gKP+q5ocsmxnJVYeI+m9je6eBhSt
Gf/wXXlNNvzay1OXXTKskfL0eLKkAxJOPJHTNTUw6ys1uEzWlje0IZiGe0nh
IvhWGX/+p+kZUM+1Rm4LFo+c1T13RY9np8vbTmW67arahb+Q82tAXzR6tM0G
xJtc7fo9XmyDzAsor6aRw/ij7AsbZhOUevPPkrTSq+f4eFGriEwBiGjIcso3
Gls++Ml7HPlAAFFqe1xEE7OlYrbCD3/Uk0gDxAz5DXbOtpqZSNiZtJFSsQbk
lOIRByoilnIINJGLsqBmHx7dc10LxmMNHz7D/NDwmaAoleLBtaUKXv9cMq8l
ycI7/1GA0pPNMAZrdFLtNDZMUyiacAhaM1TlZt0IeBqwIBMpXPxdFnY2hfwH
XNKecDnwJWULkL6K+RuCFlHPnvOFiYTXRWLI+oua4DL4HUUaa2078/wyrzrU
qoO/7geO6cybPvqvlycYU3Gdu0zVByeRw6ywg0UW/n8VIYn/ZqJfSKCj91Bh
RmitHMuPRmFaQ7nZI0uhukLunNtp2xM4Nsd67w0bgd2deumvhkCjIZjNWVdn
ZktHJsCbPEVdxJf8MQMsnZ89iMJWMtKKm3BDGQMK3B2cdVRxg1hajKpwwMrb
R2LfPZhExGsn+87nROUoAFQqhak7JlSB1bJPl7+NhnAHNg4p0Ic88dC1ylAZ
o/peQruq0CPkeCw8jSVbQzBTHmZaeDgQHTCJJ5mkYj3EwB58TTUqRqZRKm6n
Iah7Iw/0SMk8CsFF6zjtvRWcO42ckdlFcF/4rVnEd+qOP9wakNZbt5GywZtv
M2ZvFxfcdJGEtgtRW0wL2AeSbT75tYBxKVsph49uXmDbJMd1O9R2eXd/R119
e+2dJ0n0akZI12IrLwG4uPpOm9Q3hcXqDp3LYSQD77bKqNg9CEwjjW64eXoH
CclvnCc0jQejvRSO5ysRtlckPnhRdrfTbPelfVn5oqs9Xz/KVELjP6bqwBWH
+m9bX6XHiam1IlAzgxeY3z3WGY5UjZ0BMfrJCDpHhpExw+SUEHsYAIwquPEc
qclOPoa92OinywLZ1YGTD32ixZDtWI4NDwtXnCRwxNKehBdPb6hT9fJbu8pP
kss6VuldmpucSYBx26HJQTc0GZW1q7Un9pvPFxMVwwMdZvyxpqvTT99Zd9Tp
i9MmyVtu8Fzr1zvi2D34fZDQqPmRUuncF5K7y6HhBMYBvSP/IMEupxjqRp4M
pVmh8g6q0z+lzYV/UqA6MtwSBGzdV6mICWdcQDHr3WDCtTA/6IP9dAjFJuvc
M14GWwplj1kMRy/q/dKlqXubh35j+aYpaH0LgFqUr4j55RM3i/hchd0YNFbM
kImxFgED4tkAv3AKOtIwaVSKjxT8nnbpeSubtmTOlqEnS+Y5srNLN6UzLFgU
DCap/uk8Wg==

`pragma protect end_protected
