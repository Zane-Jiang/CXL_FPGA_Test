// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dD08djt40ANS6z0XqatMYqdrU3gMWRQNZM9mrNK9isJTGt/hm4vkG6xyFTM2
XZYfK1/KFQS6Jm0TGRczU7co91QW6e72PK1+ebUUqwLHhxKlAKyJ/vTym6aU
ooFq4eaEufJE3J3+F3BzHCUM8RkKBpjf8LPOkDsqlvWsUNeP8qyRPcyx2mqT
A/5tgscp2kdYvywyf0ygZ3UmBo39GBgE/9oWDCmKe/GKWghhQKubcwZx72OM
UKMsp+kOpc2sTOqRt6NftYvsfntxNgBqaFj7Lv3QqqxRi8ryBhPor9jrDC5D
UFy3+gmIZ33Ss5qd2FIq9dinMzkJDtoou6GaguMxnQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G/fXiU52ILPYywvmj3Vw0SVzShiqUU6E+M7Unwjiew7z/eRVTcCGwiIaYI/p
OJSyIb5yFVNHg0vZSrBx1ElvuDcxm4F8bqKFEgk0IJc4CVnp9Ntt6awR+jat
/4klWj+L/pj2bldlFhX4/w992HO3HgKlKiqvC3FUIzXdzjK978kf+NGK+jGg
29CVhVxVmEJyTgk5M2JjlwkdKGfhW1OU+mKTnqLrv5gjccl3yXHAXhdRb9st
m1RQQuAD59mAAAe3LRYNEfed6ATd8rhJwTgTX2B3LiVUYeAsL+oWsdibvfc1
dLszGWRJ552N16Pd9ubzBIWHzEYw6eXNF3mqy29vgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DH8eKpgKcmRPhkQo9vRvYudKBBYndsC1D3K6ZVftBdZ8920nKoDYQC4xXLpv
DlSY1F20W/AEoB8ZhAkxqaVJnqxv6SqQSrsFAdLKbScK3M7XPlmogukWHaGE
VrrFrEEpdIuJfqeQsVXhvmTEc92XOnwxmVLzouV5RdY6dtf0glJNeJgRXIBl
HaL9axfXnk09so1R1WCoeWEZHBhcGSDHKZ8t8YfZzmmOG1xM7nwI/EoE6bC6
diDaaPnLL0cNieNAlF1wB7gwPGH0dr5sbaEttJMtlDG0XBY7hT726nUViI+O
9nCQ9IMNGB+o9SRmEjUMFJxqYC296h3P4iR73bi/kw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iA2khcoHT6FQBc6ClF+L+hMBnaD/yWc6+hi43BlCboZZQkSff+9eEQCd34l3
mHbvKtSmt80v+5H5ls3qtYjuMnPB6PAZ9y8rI7Vl60OeC3QeLQ7agT/VjmNl
ApmxdK+Gi340nqj/pxBS08K2c//QvqjM5U5dQFFQoUTjYs/QHaY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
q0jbhqU6I4F90CE00xkl4V8g6oS4Yxl0ZC3XHAXugFmJEntugZWXWsbcDsTf
87s+BMKxSyTcTNVi51HZ1yJTIcK2yAP1yzMr2hIJ+zRbSd3OWo1QRO0TpxUy
0TJHHF1Smh6e6C3p89bi+FJhz/4rpfO+XaWBop+xuug0BL9HgUXDIOXFndSC
XEa/awKVtyxfGtNdnRIqoocBmkbkXdPIZe5xEIDdPVWZyU68JUk1tGWxH+2b
iKJP+Fyao3Rs3+fzb2StiGXXIkJZDkiJ+KRDCLTfO0D02p4Zdv2HiY+y4WVx
KUGHBZ1FelrWXqinqcgBEeuoDL6wvxwLA2fX0S3vp1068+oqFryoMZLdm/TS
hxDmpbZBNAHes7/ct7a9xXk9vU9qRR8UgCOiwK4QEEUE7VPQExeE4eHxImB4
8KH1qLZH/BN8I0ivrKit2axdF/d1Iu7X2lMb1tW4vKK+U2db401iTxRFc42Q
6qnEMm6pCkjXie6z6d11McqTp0ak7r7y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L1vuEGv4vPpqbLTQTIT/KedD9TKHEBJ6ARnoMGr6UgsQu+f64tTzyvBU5MjS
PofFppqzqzAdfvfG5F6zlW3OQQ/LADx2c47qPbq0W1Q1cuPb8KNKiMsyHEAN
yhPGOxy1k0xqRAF/MEES/BcLHhpJwD9PM4L+Ulv8Di+iY7Rbd3Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Mz24CXLDwcpyLDyD6Ody+MBQy0vspu1U+l713bUcFpvPDJOi+84UMDWq4WH7
8NGa+49OuzSEL7F61mS5TCBqtmOHCkxM/4Fu9cAvQQzm33pAr7NlED3MQIhH
U+JH4JMrsipxUMxssAbO2mNzMkJE0Pr+GmajIMi5XB/uxn6fPog=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
0NNkouUP1fW6ZhP+sarb3oFGXI5Sg1wdnTElhn5wd/idKRNX+FTq0v8+ygp0
W5LNnNbeXmmfryK1+f3JnO4XzrfJSpLFpNbo4V6e1oNLFkLK2y+qXvxscZNa
MPTOXmZU7buYnY+yyN5OJHMFnRyh467EC6pPZCjAm0jDRVDE01tT7+K/ttN3
S30FkO9naPUjUhHrhUkiTw/kL9MvoLXUZOnqDpA3AyDMafSsg4A3bxEOVzZ8
rUN/Q/rtCyKoIaIswWhaiuJ1zLKsHGyXkHjuJbHPhETaJ1kCNTspg2cHfv+s
T/F1dVEy1ZwqDZKakehu29+1h2tbJcL6eZPkXHBIbIY+Et4scvtlGLsQvlps
eYa9TGt65cbE8CXneqsTiqrb2H0llhj9K8drtHUyB95Zimhwe75waLVvo6mR
nU/Ifepy8UA3x07T2HvCeNRQBtGJxIU8P/fVUTQabsIC2ySKmTHDsd0uuTuz
Mr9NE3M0Txab0w4MVyd8b9XwKS4RdA3A9zh+YAWDkQGiXGk7Dk0lvcrYCS2b
UtBRtJkhG6CX2oNFlKr9SQ3u5wCwlItquhELvo6r9pSfPovFtc0buu7map/X
HpPwKR1iU2zLDK7VnMmAnzr7jZuPI3OQC2erLdDljwp2dGZVwfNvtM1FTR7I
WB/i2Y+qxn4oHokHRrVrcSpTiKGv1t6VWKGnOZYtTy0LTZgCR8aKR7HQQLBf
d0ihyZfUupKafxxjtj7vg7H2edcvioAwBZa5hMesYA5mcckcYkjKQITQX6b1
euPHi8G9Tl7LGL5ffW4E9ZDjbCfFpXFtjun0zQvfV5hvGzknVnoKhBuXWDOg
+HqqzOUPtDwVOk5CwidxvX0AvRnZBKCt+OCfB//ANlKBioDi07C5lth/h3FX
eH1VgcVkFzk5GWL0KZuG018spfM3WSQABKfexzx7+BcZtpITBawJfhkLnxcy
OrmOehr74BWJij1uOsrL7e0Q4hkwn+hbHJ5I12qNXjHde1eunUrgUJpvwSuH
m11l+z0xTdwk4EYOAiJu3H5WK5K5JcKpfaazn3JLzkCQ/3/AZF9e7/FR3hgk
mydcQsDUhMLnxSmDmcZC+RlyziJLb9IlqYku9J6STzFdBUyJyEOWV3VO9uRl
mpzVqYRYoOMFcI/k6Ma22uy6nMeOCGQlhYL9a4MdYBlNvio8TzTE9e5n6m07
cVn+3yqWaUIc5EOz8txpk0LSp6jkE75cIzw0C1wRQZaBocXqovZ3d1MNQzNG
sbLEoXzlAq0km8qUS5wz+POpc0oh7F13fESaaO3lLl3KlKyOaek6qwjvnHMd
1M0OMrrGoVP4nnpreg6JME8kJCTS2KBip5pjuRldm9Nk9w==

`pragma protect end_protected
