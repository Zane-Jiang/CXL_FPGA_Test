// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qe9umj97gI7xa3QRGrzVtHlXYaigJixIJx99LVOzDvubrKrBlZ5Ltqy2KnROw8Rb+V1MD5BtMxP8
jDiRGxWQMVyHN6RqF7ke8r3R1iVonM55wFCiigWE53+kHx7ZpEDYhBeiyW/BTVS5YeWen/t4ne8S
V18QuOyea24UUfr+1DT468xam7zFpjw/F4q1ZnkZy65EdhIV8NN4SUe6g/on/JWdA4rzMHH9KMhy
50Leg84RyDO3uMgrJFOWtIPuEDlhcS9bzEO38Q79rnxYTtNs35AQmNZYUvDub5n7vjLLJx7bu0HZ
f7kJPTOZS4Gu52vQXpG2fUjTuVW3GWNfc96jbw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 57664)
Tn2d36IgQ9zERrGhq2fmlnfeMfU2q1Qb7xAZYpXXtpc4EaqpnXhlJnOE9ON1G4WmU9nDG5icyjg+
3wHOmezuznENoTc9xkLISkwmUl4KuK3/PvM6OkaBpzVvIQz5Z4xG8O3He3VQk0mQfCrlO0JuDjgT
T5RtCxsxAGakp83EimYnqJLQBavVvevBIYIKbR2xZgwHAtUwTvGIIxC4w0OP0Bcv/8bwuA3mFbaH
6nqkOFjGOOpm5kVVCoJbsW51MM3NKs211AYMDU4x+M/hqV1BxZQSeUiYA5ooUnT/56Xt9fkIjdPb
8JNdBB3hjdKUjRz4W03Z0hrgCFUGg7xeDqGBIWOkTffY8vBV9tKzhfsJ6FDI0Qt3VY8cieDoKRCc
+xAvECsQMGJkwft4y0LAWNnU1X7FU+lg+nWydWajSCWUIrjJiJx+O7ZnPWVbmsLZAzapJa1izIRf
h08IljUlLjjVH+QPQZkd1tJzsxCg6U/kTy1R0h11x5R8VHRvV26Oy26QjrRbSkt1SkSTV1hB6yct
ck385zniFjfsfXHfKgzcxLe8fKRcfMyx2qC/3G7BuP+mn7HycCNB+Fl+n9F//mPexuWffDG6ZXDi
oLbYHLfES60AhUbbFNRL4AUmXskAxQc3xtt2uhQPAeeLFZMSDYMACrCW0Mj4NMRkXYq2zivTiza6
F2Wbroqeh4O76OwHryEeGnt792mr0Nle3Njzh9zwtRwkxICUYRoUFDH40WiZ2Nxg07ZtBesR2ah9
Jweyy/qE/O67jN+qSohxpf5MAvZ1tv9VZuOAQWMH+Nj3BzN0uAjLvgMxV9ylmFsWm/az95bRmkUA
8SSJ6E+C4QwYszNU6W6v6FZh/EENaZuyk1HFTkqtR1mfv55O2ScUPn7jo49qTU2eSuE9fYPn4LfD
eNmvrNpf3gNYY2eF9vXtcqTJKu6ksBWjydRE9XW1uL+mBqgdLF/EZ4nsV65F37TQdZOkFVlZOwMI
0SOfLjuIb2SS8iq2hftKOfgjiEVwqijkgTcA0kyHhx69os5LVNNQ0sZ5XJ/f0IPWEMdjjNVIYb9p
tnOHo4wmUCqfOFcCKU5af87kXJrYHfCEec61GcG3cj27JQKx3ANmpKFaNjNQZLxBcuwo9UzwDiEY
ZJY5C+7E/biPiI/hpVFgmb9+7c9njWWN5CW7RmR/mBuHxgV8fNjnRLUG+2bpwP9E/ILsluDQMlXv
rv+IIS+aRZBpzsMkDo6WNxxCr0GpQwUiY+jybm/KfJH4/JE9yCbpUr2r8vnZpQfNZbpXHFWJAPHq
Tcjr1CKRO6yZaZP1zIAI/CEEhC6GzqWA87wgFyN8CnFu5mLVvfTIlwkKql6ctezHtQRDd3Yt8VWw
fOJ3k1xIjOLE1YFpmYNSf/pWZKLmN+ur2pTYOzbgy+x6Mjlv7xW347u1a20qSF4Z9hn5eyqYjdmX
X6tvfSNLv2AGXwVwxJJwgV1K2u+nDHrKDDEeeddFnvT7gFhjUtJz7Ic/LkWgIm7RE60CxTX+dQt1
LzbTLP/jmgw/8egqZG6FDBXXTBJfG0Bv00uCrS04e6nuQP77nVxTbd2KaEMjwg//ywoCXgxmfNm1
pgO/fUkKXEIz5Z5NRoI4vc7J5Ny9beuJnwOl6k7tHX52cMWAV7sWvLh2go9KShDLtbPDE3/srX8f
I916N0NOVJU9Q3QdMhTNUbk7lXkPR/zRTfgx3SOsgX/cesXWCRm0iyg6py4ZFyMuk7+aDziCYw7U
LvkXUMuEpJGoAquPj0UneVrHlBC1Jsuvm6vn/dPs9px/vsWpbkpzVEo8hLog+c+/lIM20bI076jZ
9H54KsdtzXwyyeXcYLop8chQ51PaOCO5nmI0DZVBHwkrXLUjNg/AQgpWEAg6AAXNYNzQZbQXrtML
kdVZi6KAL/xLnSk7q1NxaIceWdXHNMcRHYM2tFNFCRoTzfGIHbKEmts/EDgGXp5doF4oIMls35W1
wwlRLSQ/3kwESdCG6+zszdG1E6j24F0eCrKtlZMJ0L3ZCCimWAWPHnlZLLhY/fPe4KeXSUsMCa0a
pdYPk4RID0wVLYPxEUXrDY5TSkU9jlRl9AFhAkNC2SnS5duQOJw9HgjXEhaoyq5OOCzRVddwZpxa
isq8ehGsNRwads1RSpeo/JRxQG2AFIZT95FY+7TcGuxRiKWNFeoHmUed1YLRqRAM0zGuBVbpMp02
IaB1jgu8ftf7nZ0PRLpoygs83vAMeHO9vcav1FtmAbwl4vFlXGzTQN7ZBF1Dl6505G8fUtYXcgoG
GUiPFszon0XFKRLY1sf4dKfBDAmedXK+1gExPz3G2HZS2NVc9QMkKWG/sN/ejAi0aoQKLTbdT2xJ
4/QGEbGDyXeVRo3dYLy64ftSl8Ib2kEBGmMuGb+sQl1nBq1atNbSy6kqjAceWKT6gFBL/DMNRDiQ
begRs+yk3Wa2OxHNpI4NSaRw5g5600jcIHjcg10okMITMwHF6Ek9bh8FWGgFDypjcBTChvW/Nae8
CZqRtFtqYSN6KV0ZvTWU9tSgJmpQGeaDiKi7uRdWd14l3qaxnGp2Z9X/ryTYlZqe42asnKRG84+U
2W0x/X23L0w4a8v+48wOUNyaQrdsSzrVbs3hjd+naM2pd2vdV4WJbV76QBCCqtbt49w9QKwe9Khx
5G8mzQaPpGC3KtOeoOmTRcj4BV+nys6rNgXVLXVej+u9EDXJ2oUdQP2TvCgwmeeGsquSAPHTJqpu
rmX1JIz8kv8QcOWbVZ/2FEbVm0tA8H9POHiogjgiAjLyFa2puiBzQ+ROJCoWF1SnZmFtvHHubCL8
PLzdQS2ouoHoHcBAqNKlN5h1ytZN1qkqzs9e3q+UGSjNuBOLMyz4f+q9SdF8CnwFqRs5n4XayCRs
m43ATKplQxCJn7DK/zctKsjlPXVx96Ppu3kE18Tn0LKN5V4mqJvuT8FTxJJmyZKIQksBSIzKzZg4
82Lo1h5Aek007zSds9aoXnC+M8Bu5kIbtwP76yiLtKFex8i3UgJ/OjtD6BqXm85yyAJ5DUFDMP9/
+5A8Ii5dU5KfLvvBclY9C8WAN/3ORFqcW+rS0PWUgZZV0i5meXXvUYWzeyC8rnyHZ1dt3+3Ly5hV
vqv2zgPHwB72HL2qL+bVaJ+hZlQMwEalqP/gSS+H1yELXt1tLt/gi83gdk0HMoXBENEzTbxLF7c6
y99pB/j1vovaxA7f0aZQ8QCFrzPAM08Z1GggWCZbVGcnezL2CWPkS23iitzcPb6qnSI1xmZiAa96
IhIAQJJiusL57t4bY/gHHJZuS6tR4r/DfR9L8wUjXcf6TzHa3W8kDDY7H2YiIcwp13ZHUJe16MRA
i5i2K/0Mix0VksSmFxiQd8xNvnfivnPI0O3QzSrYJhrk8lV6e2xAi22JyF1C9zIozm3/dsPmLXsL
ySjMSvah7HE+rqljlv8KC6NC1eYqIQbrfwMV7pmJaalEE15WtJLhQPbXwQyS0Ect2sRNhx516rO/
/vY7ksx2QLtNdtVoAhnB57BcmlUp1Disxv6pHDXkbDfAgv1p41UvL3mOARz+0uH8nWFgVSJOZOZ4
0ZC/cc7GjnzfuinrpezF7ns+qKilBBuna3uUJGNPyzD4iqg+hoDwyneHrM7cPPFzuviCKcE8aAF5
41Ho2ka9sO18OGeynY6PqMwQJZJsTyyAP8g7HLpys1PfqPp6F31bLe6yhCSSpoJYDjPvIcnUt5Zk
bx3KKEjXg0LEZKrLJDigd6npQ5XoroUUuqL75kVgPkU2Pu+nut+DllBzLvhyN2XeIlyhaAVJOeAZ
/icMEm3z80ZQpZ+HL3VuhWWWtsAOERygiVcX4N5GaKmFXpkY8UInrG7aWhfDsh7lsoe9JAB/7E90
a8RGY2UQgMkM3aAsbzwgBT21cxJP5Qmu3K0Wa9rhfVGzVXKHh+I/m8lF/u4mgFytwyTFpY9yMLic
6QM1fK87TtHOoIQw+C039mvZ/uwXVxzSmb+nBbgLwzAdG6bZVfqRbhQAIvldH6hW5wHBPJ92hJFv
07j9TqKNme3Wu2Q9HJCChBiyR09GnIJuEhW1gHwY4tnxa+IZBRuVaspP33V9o3eL0KBo0grMqBAA
G/84ddNY3XlNPJsfcXoIPV16tvdFgh4hWzAMMQ9AQYZybok6ErphEBWXfAM0PuTbPEtgziLnbCNT
HHRxm12FqSy47X7L//c10H5qTFQorHchx9xpeX8r0vrtqwXEi5lZMA/0yVxOD8FRi4pBFZm94TOd
+CwnQKf35sxIZwvx9GwaUjqAJyEKe75GEqWfwgED4rg+0jivo7Ozbw1zA9Mi6dx/osqZ5fAfs1j5
xlsRCA0WEEjTcBAoi+BLn9C1ofmoSeRt5F5RGd0Xm3ze4rytk7DPYzhzsmZcvtRmp1cQgQQ1500T
WMMNwH8o39iu7Z1JHovIIl2vQzo6wxDAlz3C5mR8Wblg/kKk+vDpf986bMVcQn9wbZ263DUJ5Js9
BsEZvWNqYY4T5jYDdpCd5E3v1olkUOrD+C9ANJHi4VzkCLD1OqePsEtX17jA138XrrUOfgHfq85e
hC5z2gGOIxqG4rXQzK9okaeBebgGkHhoYLEcjbDTf/9cOAzSNbSTWHznnOs3CCTuPtfNkBlDmatb
9CYQ2hyhi2LXNMmXNDlFiKtF+8yP1BISgZ5USx7GJjamKSPHWEE5BZqwGCk0nZ3t4fyu4MaocHOH
hp8W3LSzAzeRM9F3gDuJZRdLweQ/03UUS2UI5o7zZtCAUqgZttnT2R2fLrrIlouybLrFYh5oJgB7
PoX7xWhwj0q/wlrjI49t+zQXctD2p3VL+clSjgu0rvj1qDhCO3OiGWfBtJzprU4jvbbP1eXmOSRW
SzUZ+NWBwAKp6kYOXVKdKUn+Zv7fVErOxxYBCdjTwOGrOpczl/fyCK4czeKmbrJlPAbYvE+I3IHo
wKMpUkXhKCaoUGeliyBqQQuk8O8SchoYexqZWRWClYC1tP3t8lhG85sneuKM5CTnts6D6eB5FwrM
EG4aAp3p/LpGhMgFDIDZFjfcB1QDHEd9447Lb2GPnG56DaLLv677yh6qmD5bmXy9Fm1OprTsrKnD
squr8G5anu+l4zfOJ/QzkLbzgstcK564+ZBxr9lS/o/0skRCnK+8pLbUkShyFaaRmKeV76U4K7LI
ToJ0LL1uD1IkqoMg21Ucy4pSn9JVO8vk8muO8HkbBsyqKrnkmciBogkPClJgY+7HYCkW/hSHzQ+S
T+n9TljC0II4Lr1yIkhigkTeznNktWSa5lW6wY6f2PPEjdCGC/k45H+sxrbgE2f0ICzQCsWq6sDg
xoO5KsQExi9gh02c9gxsoqPiGHUVub/M21CWm2Ap5rGhQZew1Gs/KV314VQgoxQlSeuvkPD3q4xv
Cae8fm/aEnWZtkJXBtiUCan6iDdH9V9KhkX+NPzJU5ZAxckg8BKkmfWzBxj7P7TA5u4DISgFxGB5
fNZrNkA4+DWNcNaf3jIySpM1wOQYKH1sLfSjQbwoe3eafVgeWmuoK8sLz3lnz08aJPL4syzpspA4
IkYslQ+fmiFkqbz0wSxmi10zl6PQyii75JaxqOQwHDKpmY5jCyLjeQ3s+XnYglbxBMEbdFBlo/0K
51fFKObDUY6WnKz/1JJlnJzheFPTRrSdjKtnqXpKWK9zmsSgc/j7DQbvoGPLqNOmKnpEgeOPYV/Y
4EldpJu/2BsjHWqgCVuh5EDeCtNvdX/WEBxQJxe1InHG+A8zkZi2Hvpp3gMz0uclwuAdAYhNw1Za
PlCCn9iFNaFp2c1gorZ2AfmBVGoFYJDU6kw9x+hQb3Df8ChHKeV67igwpkFA+QGi2a+YwHyzljVg
4Ww7tqvUnSpY3OYblkt+pDuQifEUwMp/4TIvmjtVGwpoIBdkI5fIwo9ftuDwe7FlvFFGZA+9ZllF
BfQrkHpVHcWxWmEWrnALwVlg0nYDRdJZRzTZrtlo2toSM5FVowm7mHTdHe9V9/yyoKHJ9W4Lb5Ob
e/8yl1FMCWyr9Kb4CQxAnXrI+STYTAAQh2Gat9fUhIbX1dV3FWYBlFswHMW6WreNy0KWiR5JU5T2
m6PWPfytqbrhw2cBxjtQYiZUqyPpCu4kUZYw+A/VE+XqnY/UXJHwbWPd90fcipfjcORRdVAIfzZY
6dMKE25V4KAMo3x6GirgI6qXIAKafiKMxFs86LnSI9X3TEojNJktTMAJlKsqBVfAHVhI02g9NlXP
eOuL77EmFZ5An/DJYGrw9mw5Qk0djmfHRM4GUlHaYc/RGuof+UeGv601Rv/VK+KRbhQUAyQK7q4y
2jXEOMk8vwkkIPvqNS5XZ1jOM6wSkOTV4I2zk/2RFH5zyOSBkNyWXm4xqpg2WsL3ZtZIQDthU109
tfkqJMc8DYie4u2s2s+0MWwrFmq5Z8+vrlLgzdycS+ko+w1LCPSG/+FHzHwquPTVfWXE76BvZk6w
kf5GFILGnCP5HuRakB49xbeajl3V6tF0RwNpj+G5bN4hR6YUYwNL4Qf0WyhL/2lH//HRdHK2FSGv
EY5MTXc/wMhXCBOfhG3TR1kLLU3kHar9yYM6LOQl6zR+0YzPOLG7ib9SrL/9myQp8it+188Xu2ZQ
mb/iY8vL4WmmW9nAgodiQH680M5gRGm/PNeeY+qE++/dgYe91+9qylLEiX9IsH/FNTSv+f8hhgoH
bbQrOm8K4yof18z79jOpF00zsiCBsXlBARr24PF2aawHp3u3PYDrwbxuwXl67TPcokJHZQEuGbvg
5sw0h4uyQA0FI9y1Z8411F9+LE0iwngBVsJkQ+I0znOsfT/oZ4z+egYgjwacpV3Wd6ptathGD9/5
+jmceaA2w6z/A/LO1yGrbpv0Jsn4mwlvaRVV0g4+ZZOYh8pd90SECOON3HE3i7K59zkEOIYYzX5A
sF/vLNgQ6cXwc0pzo13vlzX/e8qz1oB9mgWtJfGyBe/owOp/Pk49Yi0mvMY2dXWznFYYOi99uXof
7iO8iZDaGIOuEEi0F2dV4b8Lr1e1d8hsFUH+5o3oRH8k8HDB7kIRz2Sp8GREXdvC1x+QqUWUx3VE
seQiZbZj8e9O/gjc/nZmKTEebL/yK1CFz6NfU5vAnePoe2COTLgE+8wiN6tbPAquii0o4Q2O+CuW
nS0sPqbC+/+R4MtGQL/FJ7h3U/YrrmzfCqrOa9vMaBeFr1NuZN540jSGm5x4/I8bJLfosdLbzpkM
nn6nTd4+qoNOGsCJTAgPoz/rINl9TCIILlKvpyPbYpd14NnZfeyE+wLU+XHDHI2Xe61opMK29Vzx
JYDhjTGuFLuOLe3KTPQjw5cIH3UZhFocLxCX5QfqvaPE+PcIr7EJISkrip8k/f+OSlqKCXo9V/G7
qME+5PAixJdOxosNsAQVFxpWGexnv/vtIa9yvKnhtl8SXcVHwvFWLjd4/+l303NYVff3ayFa7Az3
3tmIVvmJ9TADg7wazBv/9smmOO06RxTjJBRM8LF9f2jFIUtUdf3zl94k2qgc8oWnn6e30g0dNC3G
86ilXvlSuXM8p5X+yKkbdCQc1IxQAR3TrxcHBF1pGZhVDHhmJwRBgWZ/hXsNYrNr1RmmmZ2dKIIF
i28vKZ3aODrvk8Xom9/u+Pmnjw2ciyY8RyThM3oJfE90pD1Vm1Z+TrTiY4OV3i05iaS1mD/BWM/p
2C9NWWJvIvwyCV+Ea6aGwY26VIfrhR8r7HVvoB+76E9+FcWhgd4t+XMHJGtgAOGDdzI1Z3C3cDHx
m3Gmk9QljXd0sG2OIKkiQAwGJaN4VJfHrnrVncDQ/gXj81QKy/Rm2vExM4Clq7Lw83QWWmKH6h+W
38bhpPjyOAMS/DVCPJ/6WE1JAJEsmcIeaEC4RG0f2V18xZ5ipL6DC4C24YO3mtf4ivalLgGnPDdS
RXSjJ+EUleU0aUwUVo3RuftfUzvUebH6joiiXtIt/SGYuQH96L/k6x3z3nv8S1A0mqGrNyhl62SD
UsvZA1hj+/upz7VyMSuk6NG8tIQSze04GcLWzy2lKAKwP0AeEwM2LikgLU7ey+c9ZbJhrVLXmpWz
aLKcz2fd61dxW5xL2m29sthBFuhaKFSU8xD6rA3dth9br3rIlCnHsCcRukGT7DJJzfSqjfWcZ/C3
ItmYcuJSB3elwl2OTxOYDTJ3UwgDVX4zhlfiJ7LVKybwqZnEIoOBsnrdjgqKmxwDXjJBW1U2th9k
MX9aKkGCzcjQr0XRC8v3RdLsweIpUqTWK8aMR5bZGY2TlR+Q0UpG7BjfiKSLID9+XwwLyLVgf/TG
ZAkiEYYMDd0PzGA+UT3H7QYNI8dpDqGtxZ964Vfv6ovnjgCSTv9a5CMUdCpE3c1zzkM6dRGAbbln
mG/+wracEs/C2X0Vv9AVKI8f3kZ6S/wn1xqyW87CEhKDZkyAtzmCNnDX7KBAwhMKxIJO7/XWUquw
HyBmRJwbW/IxccbRbqsjqY5CWwePgFN0fHV4yJdQG+bJmBv5BBxLePP0xCk93r8il33oYFHtxnLH
pU6wVFGOpkiujDlhN0oXgmg7jYZA8CfpcSmOpZ8DR6IKgdhbYhRZYYNbLV0YGX3JvL47qlA/artn
nUmAHSAYSGk5boOF5qeWVM8QkfZyLb0rCoglH3nwxdlLEi+ePA+8+NeZoz3B3qqbRTOyHM/FDqU2
JaeO06gMI35i9S4a3LLHIqJdO/YN8G4svztNqd8jGLxPqiInV/8rq0QZ4YlciyDTzQc/dJIlSlQQ
5ACjagimHyip4IELX17Kvpyb0I8yoCRjf3/mCgri7izuq96+hsYfHKk9JOsH3487fKUm67Af1GW3
cmhQ5NIgdzSkGzjk1FArU1a3P4GoxpnTOv7K5Sjm6ko3JAPJIJCF51/1XUfAcTgs1Kqez7ShTviZ
7vxxkgXmwNiMEYGqvYk57t+G/d88FpiBUPG/dT1NuvehNi29Y5sle5cLU3yT71dkaNgFQd5N3b1G
x23ho3uhlMgaYkoscTy25bSnL0wAysWX9uCR0y5HhKTyj3eQMt97vANbYxCFYPoa4Tu2BLzZLFXS
0jLj2mTROsy226SPkKTSa5dKPuLX03X4sxswVzpuRo00obPor9gyzUy+vBAzykgptNS81q0FlE+o
XJLpU2kuHnQIKqVVxYuBAPbaKyiZ4E47qXFJHGCzbUhXof7AwcaRhR6mm4Wx02rNUpxR3b+XyjTg
dVauNxRz7Hrjc5n6fLxt/mG9bT/0vExif6EFhesc/C4ia0M17owVRqnbO2ZHHj65OHQNVwX5zszK
I8a/TEOPNn96bgYnob1smHTaw1ifz29QMnkfwSm1sxtUqyu2ogBrjVWQVOvoNuUTD7Glh65a4LtP
UO9dGxrj/aL4YL4jf+S3zqYdlV3SFTNjHv7YuxzdrItNNHPqwI/JeesRn6rxlV9sHQLyehvk1Td+
vr1s3c+xBYxcTYfvA5flo6Ouyr0fDYpfM/2b9YJ9Xq5UmUNg8hcSfbiUziMwfs6QKgUmrC9xThRU
zr9/F/dLoF7/GnNsXuKpVdnPpadQaO+nhUAp5bXcWXUiPqE823fu4IshCivoLdrLHvlqhQhsrP42
nN3rXT247HF1mUKOa6eKZ/q3EMU5LFMejtbX7YTBafabcfW39YC+CSXs4VGBF1STt8DT/fdixhIk
2ESS6TkNwMSnA15O6z5tRoXOyow4aTS74FvE47DzLav8lKscRmTM64Pw7TGfkrtG4e0l4d/Gip/H
npBZKdwlMA7oaJZKPh2bGaPtsZ2DGhJ8ZIU1DC+iM4vKCth3ATnDkHa0beYWDKzo3lN85ZCuKLS6
ZHVP9alLw5uIpjPoBEbxrWqml2UsAaoT+KMh7CAtRJw/TAV4sR1EeSKOWByCRCyRxY3AprIPUW/i
pgRcTL2dGQJb/zCc78y4NRVox3QjuK/8wv6STXnJwjkixKXwUDtGdqH0Qbe+KkWPJatYMhopg6ia
C9+OqVLJ/iBXOfG1ouH5u/70PKwHXE7uhFtfl41GDvQ0gBklIE6i0uUp4HD3JLyrzBMpjQAP4d16
K74Djrj+MYM30FoPYL+FD20MoW0bWMR+aVbN4mxkPJdNpucetvMeR4JSNHOZcRjK4evpQKWttlty
Ki3L4SMis7ZNipsTtwIqkpsbYFMrijckEnnY6rf1NaxA0E6st8DA6IaoU31GxWfX8zkNGVl6dK6n
cZxhdc6LppHcMTYp4K0F9QLL9sHQ5FprZRS2bZ+xpmd04MEHTH8bwswY5s/4TD4kiSe/Fa3HlLNj
vQB3xkQT/ejlpvpv77VGdym5f+ppPti1KLUZIhnoTPZ0FI8DKgdilUO96zmDEjCdz0PfHe/4eOaT
iezlrY5oY+LgClyilvIIDSrOIJe2qwX0h95Ls8d6gUGmobg9CT9bc5wPRHx9QTDq7XDsMqvAKM0I
raHzDwfB7EgplOI6wNsykUo+sy6ICSOs74ss2oG8vpYCbqkNHmAbrqcNPc+t3wMXk8jQHJPr0Gk3
dk60XCI/CIuzL46I3ZspJJB1T3xYQJ9Vj+dnwtZmjOiIHc/PntGZLriPmXrVKEj4DNBNnO8lcfhL
mENFBhIgxAIldmRCAi1ZsPRgKgu95iaf0TJ/37DboGUPDVAkvmNOJO5P7Vv2SWdkeqXAmHPia/BS
18zEYZuqJCPIPBtPURFI2dk94GJbg5UI0lhi1loHjklo601zWgwHYZbLOvb0RmTjy5EnYpnMkAaJ
sSQzdo25k8/34rjuq0n1eJqWN+qGxd/bAE523uScMRhZyDUVxfTaMC8SXk8WBysdBu0OMpVMhdPb
5nvu3jJ99+3edqH++HSOs/HdRzSH+lSfkLM56V4ACBthfGdzem5ENUbZcKiVnjsUAGTIVuJjIeT/
Upjib0IGVStMDUwNKrmCilE+xrKkPUnl5sLE1tfxNhNcRWGCcB7pvUOCQNy561D7YjVSo/v8kFTF
Gt7bbY8wBHmduR5vTvFuao8zLpTef4we5+Pqz73dcQ6LJFIMGpRn/nbnmbnKZ2fZA1qnApu3KRpK
QFg1LPAA0aInetpQHaIXUG6D2qH00MdU8yXNuhyfxVsQAUFpsiRtNRHpUsClkYJMpZw92LmZWR/x
C8/wD2aHLm2mFlUrhXYQIKV1/xBMM1ovzmeTfVMepFpOpIKU/wL+b7qJF7zkL1sYbqC+AvG3Jph+
20/vnzkCjLd0Qkm5IuWNG/1oR7KIkK626c8UkNw+7WtZHdOc5pNFNADJTDopXI8AVfTV80HntJcD
xUfEIybcsssYr2CyZu7G6y0AS9Y2CMw4h72cmehHpu/eiWa/yYtbOr4dHfNuAuAOpqFDyuA08dJx
1R8dgaCK367SvZje52CXqXvAcnWP+UdXVpk2gPwlzvewirPRSoEq3ECZS/oPX1wcKfZxT6XaWfoW
N7SsXJJ998MTMYIIlIU3MBMg0oUiDbGxSot99zr364QVl/+saum892C0gWbIzOnePyUa6pg8z100
hkfidpP7xEEc+5ZXzeet4IKq90Cca3QEWqflzcz5YUZuho9TXVDe1123OhlSeRbhArG58a9AyMvp
KYM9j6up0iEfnXUpOu8hkMhmKpoUS+kwM8pPFta9HRpw2OAMDD+JGkO50mq2Y2hFSXzEQkUosTHN
gx9ljtnV/gZqkrBCS/aBokwiqcLwu3/IJ48Dt/95A5C2017QT6aG4SrGnlt9JCDIeqWOAxPVGA87
uhvkJkdKh2b0CDrEwMJldvUf65Orwqf08+r26AsDlBl5Olzd8qR7rbB52mXDB+RLRQRkeHpZOc+L
21aeKnx/ma4DkPtTjolbjqZ78jbnUqX4sjPytGRLD8315OfOJKkuqjQhhA3i83jlqBIt195g7ebK
zPGHYx60dgKChv22/4eNgBEWk2JYIGp3L4x4Y15dKFIS+Be846VuABvPQhPUqWRttxkvJnxzi3xM
h9xt8ik4tUyZK6KQ5p7WHmT7R1DfHyMcMqYa0o8NljuCurjNSpzbYloHfPs1OoSe3fQIm8VX3cSw
S+gpPQwoSgBHnKDTxUh5PXf3YN5yiRFfpPYQID8Bh8WmAAEegl1fPq4PkDPYn7Ntlu90eW3jRY2W
TI5+aR0x5GJj5u+Crjpb334d4x0MNvIDNui7AtJk/Tb6q2SCkdFKY/MB13DiSaegyS1yyectLGhE
oKtvoKWdWlg4y/GotRHpBcKDcwNJYZiLuNg3cQnuQLnlRGZhFnHxCwIQZPy+4WDXlHkPEV0Mu+py
HFJ59oM8Yxi7MlNH2AIE00O1T6nvJRCmrQRZffkBQ5oWKpnTgRpmEn14H7/a5l0dRMQ/HFfEFTf2
paufME4lQt3LOPZCC3H/j2te2+7kffEdJGq+rLD/sG6ohjTx1C6bXMOeaGK4kkVRTBH/h/vYv2Sr
Pt66YHKRZ7aydThVFlAU8Wc3ivtKzr8aDwk8ncHViwQ39Q1/ltU1U9pYkfEDLO5w4l0pVlqXPWaK
zXphP0aZ1FYXB5IvyCM+YamkeAlgFf1Y0wGTB03NbYFl/J1QhthaJThxtJBSTxeVEYM1U2F6emYM
vnLkToW/5GxZwEYvhfDUU9FsJcWV4opUqF/k6pw0Ll9WbQcM9i2rnzWvtaTMWlJDCxOchYY2Qlkd
DBaPPFghWWD3lxpR/tnx8kUcEETWMkkAg4QDE+hdOp1u/L4jAnCEbKOJBQZxNGK++SUzAJUJY5IO
+TWR6uyEEe3F2ZDfNSU4+xUxR2FvVWxpDTb/kAgJE9yXoaZsRL97EYP6U9Md7sQMQbjnUaIQOxPb
sC07SlOhFQ3rOGqRZXfEgYNi1xBJMFHN+3eZHgXezIGZ2v6EBgR+vPQS/xzvwEmFwe0nuPlyiFZ8
clKbryq9fcPdCyh0yAnHC7Y2vKL8gRrlk8oOuY+ts8bZOD1GeGHyF0Vnw2gIBEMbjDbS68GDkYd4
ddwsooHP6ESQLC+uKnfn+0yCfUWA9V8fZTFIYrXLon2kQfu/mX2EpQMZ8v2cgAOhvARQXpvWOBBs
xvmxPuq1YYR0VHlnbIbTfNWxD6dNrYZm/uu0TvVzaj9+C9Wv9HMqTX3DTP3qoPRpGhxAaaqQmS0L
J+/JgG5US51Qh/mOw08yoCqk3cQuFqRZen/oR86pZ5rmagVaSQL2EKnQYFbGocaU3APGN8U70Ayr
mdMNeu3wXUN9cJOaaa+vdPWmHhCrESt+GwaYKwLAz48COnJQlLxUGYLHvZKw1pxb3yxQm3icjOOs
MADSMY85xRUcen6nNNf+PLhLIqRWPXgozL5UhfSbmGqCNUb3mnTf6zu26G+kCYyUwJWfa2DmR1hM
+WCVw4yRuxt5X3fTLrtZIay8LHT2NBBRJ+rn6HPpAb/TjVqWR2iXAWJ80zUq3vdmnuOxAXiwV2AI
lsh4rN744G+CoHblHYCh285VcTfUaGkDQID+Kr6TySghHWAHYEWxWogHszHkDcoGtCP88tWrIxrD
A2vHyE2888WgizgKd2aO68HOWWre47kOQKOP/5lF8h2Kolwya3u2pUDnZoUq7b3IBor1eBJMbZXk
WM4+slyHsvh4ac7/sQ37sdZ13ooNQAyE2KHNUd2wsGYfqveK1f/qEG2B8NqBeg4rxFXVcnGGXqJ2
bw2DjnW2F2PU4DzA9nv39B1jbpleuXufgqBRPg7pc6U2CJd2UQYrs3dNAdKlblBS3e7Vg6FPfWy8
yffFC/qo2vqQBqjg9OsaaWODOwelr+x/juJEktGHj8hQk7BkY4cZ1WECRU/jtUNwYAnZvFX5LjpI
44MI5jRVI6nhMMa7Ks0JRwH2bnH0mjEOv70TK8gG5bbNGVfP2zBuwoXJVA8xfAD34ofg7Hc/AUCq
XExqhVF0ciVu5mK+tIrBzknL5vw9g9Okc8mzYaF25kyG4vg8B+TFVYDDAZTe7kb4SgvqfIxW944a
8FQJLFS1O5GN5VEbDtWuTTcRImx+1X9/AyTtrlb7DqwCTap8p+tS1sq1kMKve77XzXJCvpbs4xdP
V3QuS0ou+9eOUrgcgMvUI1+Jg35TMrKmv3G4I0TlIDstJCn7W8hy6cSJvUw2B+C1frds25+iWOgO
EbhZtQxHnf+zjH62bK/s/BcQDLEwg994x67Qm00/Em4/gkKQT/2Eu1Q4LIvQJwkFXxhR0NpcE66w
p9q50QErT3N9g23sbYcL8o9oBF39KpQTOCHHINlTOA7MXPN/yBSNqbvu7bQXazfDUzG0Ucqa7sJg
TXDni599hGGKfk4xKlBmpzwkmexoCD/HhmNzUCGAxTXXne9FcVN3PrU0rMU9cweyf/w2fkX+W/uq
Z4/GLZVEB+/H4UCwjuGzG13ZT03tM4uHtwyoYwLFa/zHTU6xMi8dHx52DzBgEuhK5IMWT49N24fK
ho6gK5oP/zGBxMVb0vrmKJLQnQDc/Om7GMaWrBSlMsEGs0IW5pQlfhdaHyRO+djkD8GYCVDve6zk
GITdkcSyYFT8PLSmlzBlNmDcBFOoZLgoHksG6IwB6ctQhT0ONZwjYmOy/XuOzPnOt8avlHcjJyC7
aYgKUXqkqsniCr7jg42fgB/yCHOQpegNJZUVRbVujCP9+0dhetJs5vLpFIOTsknVS6tTFlKXtPrT
JjKi9CFtrjg3nSe9Z1swNzw158o48SUhac+nlSTsgfb4VWNhTuz4XMGzNwugbO3wDDuQUAnJXuma
gZGe/l6hJ2vJlDfSmxrZKFEI1qpH2HazDzkr2VwGF1OP4QYQiVUzC2URnI6lZuBukIxzjgckyJYm
HXkBPo28H0KmcnB7ZE0wteyUEdm9xvlHhnQfsvgEXganEbfnNHtYa+ZFxb2vGqRmWdkVio3kCnZZ
deWDtf0k4zv8Uhvk+BtGLZ+5DEefbqm438o1yubuDC+VccmBo8AJKYrnGE+Nn/g6S5f5nL8Lc8mW
8Pfa9c3WeK9OfzyNeA3rA+Dl1DxC/sfuXozCPbWoDWZLv+ezxfkdmkVTYOwGm5fOzRl/SbkeisPq
bhNNCuvhiqABh6sM1nFewo41ijlrJytYumv9m3D/VkYa69XvXIeod1PnUmvacVJkm7sReEkwZyVe
PQoXBYzdanzWITTEp7qyPOqZSVRxYf5rwG5ketFNoE/Ur3HnXIw10Bt7QbGGflsd/f8KnR5Rb2SI
7a/jRX36ZAcOXo24aspzEzGY/fgyDfHBa3wsJRZ+3BgBxcQUpSgQC4r1oySTterNeENnZSXIpmKW
mMCyrGDXPCU+haa6QRmzcHSjUeZXyUyNh9rdkhzdw64doQTQ2T/or/73KuxlHacJuYXynco0iHtf
H4CQShAsaImU03KZlaps+GMICum1HX406/Js381JtvDAvInh76MdBTwgMUQYL2gBYS+27zdkobCf
6XFgT04ANKrLkbtjOX3wbaiJBIrQocQWTy8OYcT/F1dMPzlToUrrIai9S/SHI8Mz33zEjeiXF8VB
iGpfqdGJ4IOAE6Ch7CSVQ3f/f50hSvsdmrCwYLkXV2g01p1MeaaBQ49PHJtx9k5fiFEW8LNw2lT0
wongY1a0TVUvqi+EwjYOuzaG5urpewpOzDmhKSLDTC1pxYGJfs1/E4HxIYZOxeXVw5NS2uLZCYnC
Q4lSGKotTzwhY/yJcQnjHiYCpfLQtxSi61NyuLnE2skpYfzKFdMCoqf0Cuy4yjLmX41bN4Y3y4Hc
rH2iVJUewuGRwRkQ6NjKK504vFzbb2cWTlXb31/ClZO2BIKPczaoAokRYxFnSfopDru30SLJF7uu
DLG2jIufxYK6MGBNK5Z5SbkPDTgFuL5Y6myPvmzdTLw9hHpo5sF1/oUn0RYsp5xirWFeeP1g2nit
P1wWj9kwvBltif4jb/+0ugKmpgrhRKyVyPhkP0EPJ5rAmBZ0KsRrSf+Mp+uEb8ArQp5zjOvVlp7U
IkjFqt0YKGt/wO+Dw5o/PzyyjxAkXpnkkjXrukaVcKPhfy+tzayAH2W1o0b5OizV3VPmV249jf60
IOxCibicgH4S0LYWzV8nvoVVgyR9N0jt0FWKXBDA9EBK6uqeYlQflCTBrT7GucJYp4YRWzz03JIE
KweQocwTeuWJLB5Oppdm73XPr752+y2LyevK+4qWIHrgah+bv+g+iaK0W0WRBoU7j65Q/cInqrlo
U6YbowXXllbtmBdRAcKxZp0hMTD42DM+cI9ySyE8qyBC59RRdZRS+whE3jyQ3++YnTmflAiZ9YOQ
J4SMKRDt9ETbuoSMUINDezN93Tstrjyqy1ZeOU5YhE5Ngq4IyggBOJfgEnOaAANqmHL6++3A2X3T
d6VqMBjXqG/2KgQOfF80gpSgzTb2yBBSH/QhPK/FGy807blJPvG5kwAztQeVhmakzjCwIFGR2RXr
iRL5fer2oqC4DC8YvFrGHzmH1PwaU4A84/SkuNeB5nQnxSHHj3hRh3kPhTWz8h0eUzAgfC8W9dEq
qKh9DOpnzlWdpysTyn5GEZKQU5y4758sbAG1dseBTIx/fSOH1m4OB5tl8Vsob8+wXpCEfPyM4xA7
7yhBCxcFT8WzqT3/f1N4T0n5Plaet29eNbpdblGEKPH2vUFTA87boCyFNnO5zhqoqDNq/XBiDMRh
ZV+1ZCNaNJOF/IL+w+UFUL3DTet/mrrEhCy1a0TV3+btyLme3rzriOnj4RDfc3Ijb9yGK6H8owKI
62fVnBWGzCAGtlwBcWj/579XEcpSBK8FVbIE1BhSdzAQrbI76dN3Vorxy7IpfiIkJWkNsNTywJtd
fegoKeeB1yFsJR6IPxCuZhPOMF/HqjXDtXblPmBu+jdNH5ijbo14ezpNuoPo2A20E629HGvWn/xU
sBfiAcZ6jSA7o4bzF7YG5uoK+BG8axrzR7EMf6GDrNhXhjyCLb22rkYSWhKoQZVhATnzNaqLpnCe
HNVXhc4kVWEjbL0qOnkZ1hQUKDYAtK9q+I9oWuflZPJ4uAIFiDLZ3hs8guFo3CG8WKVUjEZQhEy0
GoM8IatHVpBHmmBsty5W/+flD5zuABlbKFntV5JbCpuk29ejB/IiB0FbldiAOVAalLGJ5E+W+kjX
Mku5QxqPs1KXmnvqFK9rx/7SYyq/ONeamdTXsaGePkhE+lKfUZYSYYP+ekKJZo9lU2wOH62D9RhU
BCeRVju17FgsxAxJwAzBS4nij8ROWgcZ2J56OyPVhnNDZYlaH6k64S4wcLwS9o39dvFevz8JeZ2w
aDYqOM1wwP2eL6hPKgJPug1rslcwvxWEZHgbW3S4GcxLyZjjoVJyEszadYocUpeSsFCyIGRCbZL3
BWpa6ICIhWnn5UtSTSozaOoukhYJQipO9eDWh3jgLx7U5KGAOYEVXVt7ZZZCkmgaOTqJVZet2att
ktg5DTpgokwpwW3/I1gcAChKsq4TbqxVSA8GXWQUnzrA94xhaNsbMVxK9VQSZ0fkUHdE3hfgHtj1
WLlsa0pzBCn4vmY79F+QFtJIb0RzP7hCz5v2zlMDSE0bzvNNmvGKTM+lMmvudyWjfmOhaPPLGmhB
kqcFSJQZYf+F5KhQkqoddyLAfXVIhhLtV5yCXIkP1XX8QazKWbl0ND3If6eDrwnjnzfhYTKDeKKF
88sfQAxWF11YcJYDZSlsJv6/P7is4bQ07tdzzXkUcsKwBeMd8bYB0UKVSYggDMZQ0DezbNXwcsbb
4I3VC5Ox2DyIQinv1McNehE698EarHkIahMGT4rYXRM9+bjPo45wPJjgE34El8Tc1N/ToUDEd1pn
AzuGftvPwe5d97Jm/wYvO4vwMStd5UfFscMKBlhByp2GuGfwRuxZzUqHR3s2+JBQIct9w4SFIv47
dcWzRX6xeAZenrBYWIpHuboDJ1Dnd0/J9jBtLSyrDfypKiXnIqTk6pItBB43+9R9kcYyT47/clW5
9pLisyxt8ztHSjykZyZHRMSF1V/k7/4GC3Be7VJZhbP8IosCQkFcQyJO6IAIzC/IKBbvLGlfdxNv
Dqn0OuiDOKhMOme4ve7Rh96RBmZobNfwdVKylW+0lr2KBu5L/3xYyXoFSrx+Uih4aE5M2CGue+tT
lce9X3hnwdz+BvQP3pYF2odXCiBEUlhvYeDKOetfXerEQ3vJXvRdUPKg1zES5B6LrxDsBnC9AK+C
rDiXSK2qMZh3QFD0j4dzOGaEtY84lGTEbwGsFrYq7KREoIoM9LmV+ru3rd8WLzfU6okYCUvvklZ2
Wh8HEpLPC7kujqAECXse9ky74FxqEllv4BQQmzwec67DWgW93o0jurE7k+SEr7q0d6Dt1xZPVM4e
Bc/flPsTAUYZfiUZMy7rN4EQECPgm1JrMtDvt/HAMgNyqfwtvIFoHvq+LdOWxrKndmpmSgPemvCE
IediF9krysUPMa8uoMPhZZI5tW56lfvJ5HQebb11bkxAM118rJrg+Ktxs56ssIQFCadgc2fL7GKW
Fe3X+ZOlW6bbpCoG01O8/MrSMSCM+mYtpLz7SloqyEosmiZtZLfYo8N6tSylMsqWuo1jRzObkfXz
HF0dm2hOqZWXVR3xMgiMltPwXDi7taDdKD2fU5mGkviexFtfYgPerJEGL/XMXKLz9zyDfllHqb4Y
QmLzd9RpJJ11IV8NWjgG0ru3SA8WtIhjDNIro92m5xD/La/jWB6dtPRN2bgZ65cH4CB3myEgxzxp
GzrgNke1fYCZJLtFhLot5Y6xbRqbHEFVsDy1WjPZQRGCJUT+eg2gifBQXQ0mokzCWg+Nxamcv3LT
IvurpHvbBfpFZN7B6SAbYvDkFBFNFfYhtleMxtl8Y3/ilObVkK8EE4yFI+XiJxKnaU1XB9vcIwYe
X2bvBN/kSCB/1vK9PBH+Bmz2A0F282LLEYQfKkI9NC6or6jbK/xgNyLYDZA5bdqH/E3BdKO1M9d/
mV05BbTFxVAMRiuNeB1Pjn7eCXpyflB7h9+MuRsoUaJe/Ct7ZPIegu6DTCh7ePZump4qQfRn3SYG
/LVIE/pzf/0qUVFT1wtN7mh7zx2cmCzxkF/rNprG6D6GpHVn9OEVvG+/Ez35KJ2min4lGKPPJ/xT
F92KBP5qMkxoYIayhjXDN+QvrXXkqYhO+XjkcBxiu+tW9X7M22Ow7Px8LEpBx+7sR3XdgG9U35L1
OzLeXstvOXPmNV/9Kjsg+AE3biDiSkNb8jhmEqxFSEp4z2fXZhGmskQLmIbTyw8Kmg+65lSmGi52
vWFx4RgiKEwRI1b97xq6tl9X5jo5iLzc9CQSt7hiaqmjUrBFtrXEcetNmxGIwz5+uSN9jxZbdQ6s
Ns1yjME/jWci6Zn/qOs7/V9TMlkjD/PhmZF0WgO6RlumJNeYTt3esBNsJ5/cXPYOQmoNxHzs+TBU
3YgyRLnGZ8qaYvG0xPebAGNuWFJ/B5X9WEzwp5KPOMwqcy5BWT6y3x71Mt6NetXBI1zS+b1gJc5V
b4CJZdumWqiXBr/7qd30eAr38Kj4aLtBqoj7LhxgtevtA1DXQoOWkNtZTOAw7LuQzCWMTt/lrOoq
v4m0MuabWTcxSBox4DBWHF91IF1vIEOY3DZG/58xhdIzQpdgiwWJDUWdMXYRIveKSt2d398hfUCf
NGv5R8FYV0QM+m+oB+UADNk1LBfR24LyakLmlK+oFeaCW2fuBc21M5Wpb5EHLjWTAW0wjd6x7ool
O0Xvh7awRLBkPjjvZWPnOrUPOQLvUdlWi0hC291QSnTYwpI1aF570hTxB0fA3dAo9M2/0yBNASU9
DfmdKPA6MiCUSSYYqzeKZhzZXbD2hCYTY/n5SjW3Hbt4FEE+IToWCTpl/Uzgnw0FDWCP68g/u7Gg
ZGbbgFzAA4EutvonAkFd+IDKMaVZz9pfAiyeXko8jW6V+XQxw98VyCT9bKmKTnBts112z1xh9gg3
iChELZj8lFlWajw67bgaR0ujCbwXEEmlxi4VbTPl7mMHNkdZiMi+qILR6OfmrDKFSmfCrNVmNx3N
xNp9JVnlypVucaPsquuotxgw7wbeSbW/mXDr0VptDxNC4p2OQDKqv2TYfg1Wokkj2QK+suBB0vt5
0LjVnRLPPXFdPFdG6CQAcJ9C1FGBtkG3cXzxjiHgc5UGnMHEJm5gQt2mi5fY8wpPTdXALvs8XbXW
goV+EJChY8MOyE19K+40uIv/owU2s96H2jDQaYsBrG80SMzZ0NQsHz+ixZ+j+r+vYakWlOMAnNDz
ggvIS5k3T0/KNElvCjYOsuKZ+YHaX0LzvJsDnpmJ2FWi6v4+D66JynoQrniv4I7/pViHy3Iobr6O
NP24ufVJYFwPmV5YLaE2VhSXWJFlRwMB0aUR6qGjLbbdz47AIeQ2xIjfp2Z6he9rRoo77P2Lv7WD
TdfqnKZb/mTe1E4Pn3VbF0TkqhMrL3IaC686ANKekuP8NEqNMCiTI09Zcv+8zUm1DGioKtRDwb6V
9j3V6Jhx9qXNXPjNmAQw0hTQalg8LzM/qX6M8WbKip+rfyqBnBJiFAFDLmilPVgtgb+N6HdmQTNM
15HZPlRMvwKk+6gIlNQxbUCw8lsPKIIIoL7a6ilMBELSHkMxdzX2MGRHB+PM08bObcmasgMAgydH
AyjNXVXg6o6mnLhAlw7EcZeeqcKMzTackeNfONLqeXmPhu7Rr0ugbj45pHO7G+xF8eigjT3aHn5U
4Lv5n8NKEE+Xhlf2HYs39/ZpUDrgydcQws7KHwQsyHhQGY4kAGV26AxontvFoDLG7MNF7my4TsgY
QCzI2iLtrqRlrQoR0ZevP0xN8rXzWFzwP8UgrTqjYVGl9A+OKZnLQLiszu+Gjd/C05U2KN/T4hRX
7iAuU6In3Oq2kRCdUpM7lLfOpkjrGF2znANSt7qY8HJdSdJBiY5YJ9hYB8NqdkDrJdbh7bcSm9u9
CPqQKYvxJTxTdB4ZQsqMGWqGyt4+cV5EBq2RrA9qsVj262a+KUKR3+u6Trr5uvuqB/hHVyjIipPa
zI37ufoka7MUWVVIfp17VLVrhovZ9aKmnfCZZvGiw1+pOoC8J5Egr3eb0LQ9KL7xE7PLBEbYOpwK
lJqlVEP34TFcrScviB2el7eqFBKuof47ReNEugdSIwCi2gaToKGeSFppqogp0QqTQcyPj+1MijDh
bOmQ6EFw0p1DWBy/JYsqUEhiJFPv53CWWlUqj2L3qfej9wiUpaBfOqM3FAChzV7NLB0PAyGT4js7
6csFOa9gl9uWuaTXpjVYF6YaZwD4t4ku9VooNzQiT4KLBE6Rv9mD7fsrAxSgQ7xbkH8oy+63bNAc
91AlklY/3xQryfTENDEu5iV2PyhasmpIVLqXYa1EmDNeX6OlttHeqwbLzkWIkx/zRoYB/l+PYJZM
Kb66fJzoM8jyZTYYy+QEs6j+ooPMtB8KGccAYknmchDcs9rFSeHMZ1wXkfqA+FCrc2kOEPpHNeky
HvuwHln2AzCZR/35Cg5iTUo/ihY7RGeUmC1J+dfXL6WD1P4eWrQa1PVV6/BhGSd40nZiOGV8Iq6Y
LqICrEhAt3OAfwTPMmWxd0sjemnymSTWU9ElAixyAeQRvpSmHcCJA4s1ouTgd+IN/2MuNOV+weIR
nbGCGozfhlLQxHq4D+Fb5TX3xHUZ5p560R1OH5DGfXbb2QAWzAW2+70Q+bTJZAgiY8Wrnz2HjW6O
3iIpcd0Rovv9gsxGxxTTCJpdeVEhsjaeXcGN3TGJZTKSHy5Kvv/qjcVwe+58DrSCvQO4PIVCeXxH
NnS04Pp/uyw7lVrUc+GTeTHskFrGIVg7/io3eVf8fvJ7hhgxiDyJorORdKkY0lfv8w5rNg3mgtsY
NC3ux+Y+lrzW+iZBL9e6YnhrEiCeeiWLuRYHOJGa79cWvF9DJDDoNbMvg4fie2ODrI74iEYwQF/g
A4atHmrUltP3T8aUplX3jkFGP2YC0Jc0RUyGuPlaXzQ97EsC9psPnz2xvB1wMdm4YunxT187vEtT
EggrVkLgJC1KoUX6gip2lOxzOqVbJ1/oEjyQNRtFHuiy/bOE30VR6tZESdnJ5S9IdetYxziKcNKI
q3GZt5ZOQsGHNlI8zMJgDDPNrctGQkMHHWwthWJ3CItH9+0BOU2HfA2VSGUsS+RGjP7QNWAmU1Ak
CSOUcA7E5B5ApXy3iJdR0JdZeuNeSFugw+2i/GAeHnM6YW5b41lbQ0BAFGcm7tbBHa2EKIea54SY
BUm2wfOQcy8lD1BqKDK1zkVZm+ILU1ZdfemO/4ISambd9vKFsVR9dgArFWo+85kfYohH5uz10oJR
HVH5FaOJ20SDz3xiyYLBjceGd6+JqVh2h92v/fTw7jzarDJ0swpnvIY41X1ssNiLsbaXnJK3QIkY
y4vQ70nQxLbouN8oYa4CDc3IajlzLFnQU8tHfToiM44aehpK8dWZY/uA6KT2bsrL09KDqt/KeXNV
XKgHau2N1tknFEiAZHIlrzYh+baYlx9MnU9/HNLvXyx7IevpYon+Xe3VzQS4aJ1xwxxmH4qf6g9E
MfuZW7GyPj0Z/lmUqkfdEb4XYgeqgrcaIrrHGqSCFk4GkooZiT71aYFEl+xXZXY0pXGEAqDjlzbi
yaeooRq2MCCYDxsq144Rx4xEZ1apEK4QwtolBSHb/vff6oXh7M2bK1VVNc6XXdGlzMWQAUv5PxQj
w6vfE1KFA46BSxs9b3oNVmrxN1Pu8pb+9KqAA8nt+8VScYP4YmO2+NRRAsaZiuWtnnWUfuO7X2KX
MbCHEZ2hnWCiRhU3H7zRIWqi/SDuhm/a/uXQbYuYFyoXtFW1t2fV9G7o0+OYfOmWHunNBEq4JEPq
eqGXbKfMinDhxDJJusKx9uKJquka+eHq2k1/WgWAjnZTDrQRwzcUo85I5PjRCIBvoQS8NQ4AgwNF
+zyE11nji14XzlOPwaoRPvZy074wxnMnoVlhPvUw7mU/9H3ZwIB06df2jICWYjm/tZOgw2G4Hf08
zqWkffDgq84G8OfzoKI7D6s04ofq8R8svFEyYKnm3sAjpvtZTEfY1y46YJjy1T4fRrE+roGYVRPw
OQSJWTdtXkXoj8edg4AmotP3mB0aPOBRkxgKFIHKP17m4ta88Pz+9dxBKaY1+GO4Yb97/v7nr6eB
akVdLOzO/HdRHM2OH/j60KRscEvpn+jyxKrQrJ9otg3CHwgjoayEWu7CQ9FXK22Aox0OTRExqHTS
JDILeSytbtlm29M2YngILFBzyCuVEDJuTqOOVQMxa4m9jFA+RsQMbvwM5o8Rx/UfJQP1pX0LtC+G
VnjpKmmIbzjJl/XFLZXMUxkZMEW2LOEcm7o7xRr29rFn9ioBQtqnFMwwgxa5CirWm6ja92XMXqho
hvPKeuiKDeZRblldzHxb0Xfng2z03TwPgrLVwjrcQxXx7759tQkCLOpJrldtm2YSM8Fv5N6P4WFL
u/U8j7xry2zGJGBuHeMl+gDkzK55W7Z2jtTY5t3U4EtwNV+jC9DAPdkG2yz5m+6RKw4TVv4ei4io
P4004YdQs8xJG753DdiXpr8HEjGFgyZsCzRwBH2nYhrhkhngrrrNn1eZzI+0f1gANAfHylWB7XVI
e8yjMwvCGuoyUQJoVEKMjMkTTna0e1P+BhvyT3ClNQImOXTzxucw/5SboTNEknVwWKD1a27CoQ3a
z/g6L4F8T6zf9+tNxXZ7OaQ6oMaHWjHUqOObQ6gGDRhDb8UbTy4sP8vZC6xyNaskp7m89HyGzNhI
59AfmbmvZ90s7jYk6BM06VW5G+9bzuQVfx9cMRncPiAt9+f/x1zYswK8nWkd6dEvyqVKPumAfeAe
evYFl+9LWKIi293xTIGG48tPFpS8sofcG0iKG4qPIkBwRh8wMocifW4ABVAKiCC4qj94M/hoZFOD
mUY8ery/ezFUFUfY978CVaJNwEUoeV7+2ZgzVAjBixx+c9LVXDggoAk/6v1bpWPml2J2JuBK3nb9
UTfdFQ9YEyZQu00/xJ0fGN4iRp0Na8NZqPjYzXA4yAwaSvsalTQ4vp16xsM0jF+INdHZRBKLhrzi
wyG5drpERbuf58Q0+l3s63RNys7AoVfAgnsDoql2vyvWfjePTjsZOhaV84O/xyanyH5M4eqF/a+u
MhPC1dG5TWewLgSMu0jK43LDvBy29eHa5Tb2f1PL1QIvH65+udexhBW1ZtIbercXK1mbqaYbj1T/
4lx/Zznrxw9s3seDFVUwMls3LcJUx5xexI8HtzpMAuUZT/b+M9oi+fpP2+0oLSpKF3V26DHKiXNh
3F3q+2JcjM5cOU72kZ33dpc+nxF3CC2XRoOyHDqB/gctO6qegNU4tT2ut0LrC1A8skF+gqY2H2TX
XJ7f7xb53ofA/DclVkJ0thh51EoaqxbzG/vxLMNMy1Euc8BNGeDg+O9/WnErttdhPHokJh/8bw7J
m/EuOhbbnvjAmXJBfCd5z7MwqxV9172yxLfE+6SHxwpijW2hKBWB73FgTLZr5LQ5DmoXg+j8v7W7
WGnpyyGUkAa1ZVlHCrDAfxtfHMcYUy5ShHKwD29VU6biMWeBOLyUGtxKR3apVXQDZ5SjzSCQEQgx
y5tjeEy/Y31mtsCMVEw5lp5j3VGTU3OR20vTWE82BfWIOhcwU59SLr0AVnpHxJS9mCin1wCD4Y1X
EQ7sNdenvHq2vCFGsEMGHDiKBR62q9nhQl9oOxLye7TuITz48LZugy8FrsV9fXvj++nHmlJo4Xtk
X9bUDeiruR1UgMOx9FIZC7wSD8MxFFOBAe0FW1Qk4OM7yV+sE/XdVOMQGaBASqahCQaDgCzB392F
fCRPIbonff8IzEle2mILSQIUO7DvuZcVO4+aO1hUVYM1897nNd9SEeH/qCHR1pB/EIQO15tvYGjC
o9QgOMshBpUgiq9vLwhom0/VLWdpckIxjhE2mZgmxCiftzrFrmr5BjmaBgdjAphKrMHYGJkZJsIw
FCi27xk5XVrl6iCRQN3/hgt2KXltuEeolLUozTxpM8vvwFRN6IA3hx9awqWUnieG0+TJ/g58jQLZ
tdR/ZMnEMR2c4D9WJ3WuRD1LOc6Iza2/8ckKSUOIZy84JAsOW8Q5KlhzkyUoIB6Sg1ossSQA4wsN
B/gm95jRhYPzPWnNeSEWEYWdkIqlgOPA0T3MP2ofIjAx/1LPvMM+LmO1tGwk1jjk0GM53pLDcYdD
nD2OLDKx5Ye0A8kWIzoj51OMHFbx5hxcEiwqFPEj+ylsPb98qXD+L9triW1o8IjWNspFLgqrd8Rd
96ied7G2m0ubHIBZhdO9H6qPOfMyFeOpLEfupDlvACZLAyOwFYtht7d5WaXkVU4IRYGaIeUtzWwz
2+NndwwlCx5C9fkcOxM5QGRWdSyVvaDlogUkM2Cqf7nqsh56KBeteKYJUb9yYavZHwONpZ3jgh2A
x8cijCExFDswSD7z1e1GtQPt3kuOMwPNoHYu4fLjCbD3ac8PegSacM1vZdJVpay1bIPkSugPPACq
dUB7zp5M+1jC/kclWG0xVk8atfEgwQuHAqh8+fnrcsk8mmkSJ9+6Zyw6OpA+LBJ7hlEAvX4zc/tZ
xfKfMsGmXsGVHn1h3aAAGbVYsBCiJKcVQVbhuXomWGuoKJL/NiphX9ua3sYZC7pA0bXCTammT2pu
kwJIA4fqxpIeZTxBVqzS3JscG/3EqqIgR2XbMQO936taSk6itxoacDB9lk1BPzyVNg33CtotG6SN
JwPmyvRU9iWeTUoBM9AqJ4oBZ6EPtjOD7/STdGy7EcsyRmhtEF857TVYoZctZpNZ+DrW+hw6s50Y
Wtttll9bK9iO0YxMFQe2dMUA+SmjBNRG8j87ejK33ClJTpp3jZVo0hjN7vB44rSgoEIkFbn3lGaP
Btbg1lMw19HvamrmRocyfZyl/jXRlKmPtpGyyHpRVcIybYQ0ZJGN1B9C9rDoxBCTE+eOL7QE99T3
fDe8i79sEh4eo7h4huzRQDXloBwUQ/xO+iM4rX1lgAlx9ieivS8kBGeXPpoI/2AM5iZbnpVZMkV/
yA1B4LMb2/OYI/Gk4QQqKZU1vckp5Rr9sUHgXC+QO3U/PiUBaSaIASlkn496Y7CRrh8hKkrzJa8w
6dtP2bqOsktD3KsiJMgZwZUATq+tbhB8dWp9Kmd6Gfs6f+D2aRyv+lunjvEL5jK5JsGJtl8TruML
U7RokieEKllDFX+xs0ztEdsrsqXjywKkPIDYawkV7TBgVuU8ftUzbcrhGqX+xBOfxlpxNb7FN8LD
ovBglGbRIGiF90KCGiSt7CdGYTUauDdZVTkTWjx9v5fy+pqobjj0pCyTPAFd+7e6O7MdTQFY/4/0
ZeHk+Cw66dkqsGpHOyYCPIb+P9ik0RrQxs/3HGoRi26SvAmIf36nBNj28uo2JfO9rapV0/F8h4Zn
C1uktqUZzeBI7YhEmhDOvzqIYJoGgwpv/U4ukh8uCIDbD5QGRsum2oEqRRmtqZiVKVMb8oQqzY5L
pjz6EQxXs5r7IzktNRnkdpnwotH5i/gRRKAfrFacw33RGOEex+WCkoWwuu24zYVlBlrOE4qI5XRi
s7otJdF5Cz/LLX8U5rk4q7eGVObYBkw0Kf+tuZQ61gmEKt4r/Ty0kqnDI3Fdpb9Z+UrOF9o1MMNN
f0mgl9ODgZKJ4e+VHLkqO5g2NGesIqE/X7I49MT98WJ6K3/D1ykaBi1GHqSESWV9JlgtXOXdzQtA
kymeTkLUN4xfWRSKgp8unoMXuRudHgI4S1Wl62uSL+tyNEUseQJZ9ZVA8D0tKXTyObaJfsdE1njB
Rjekgo/LVFx3oWuwtGa2KGCqZFqyWh52Q3C4qoJ2cItFa9tXoHyWkOJCyMFP8oq8KqtJhwAjqQ8w
Yl4MuH5eFd7OrIxirMyDpO6zzjn2tG8fXEm55NoPqSZpRao1zptRt2Opqrw3UNJciG7WgS8mazZH
1d9hE8bgUK+yxcvwnsnC9fyF/mtyDLRB5ixdhQyMPSLQGldZ/+RBRjADEbRr6Sz7OdGtVB8joFIk
6h9Sc3zuZdDw4pDm3eL1Nq5dsMDFJL2wGCoiq4CoeUoZEm4/4605mk7Nx/mNWREJF4+2SIRikvLv
Z8SYOxHf5dnzHcchNmpYqDOxox+/NDDhfAdNj5N8b49l92xJ5QcVtTv0QTPZaQlPXyksCp5qAgLo
dU2d/R4AWyeyqcP7lFSQBDm0x/lcyGrW2C5Y0BemyB+JxqMuvkqPpPowyMQvHI7ais37fSfHxcTa
eu4ihWJSB4EjtLkn9ez4gcbcLJdJZA2b94wAX7x3YvB/M+N9+4BXrkZO2n8f0vzj2p/aAWsyqV0Y
oHGZguDDs7RLY7RjiTmqpZoiDSQ+QNX3sbu5LHuh/INvoZcLZFWQiKwbSdL1Xh+8JniMY7craPvn
Xr8ndw3v22UuLNDkymzE+Rb4Ib1VegZJ1aho4/8Z9wOOiHi1tNcQ4xrnVu8n3IeDIewrZKTSjhsT
3J0ttf+9ICLESi/HruLZhdCfMg0X9tDI13VJDEqTjR14RIBpkZfWKZaVE9pZvlD8bI72Mdfrtale
skk4MqjlRncup8kFwjIohd4CvYeTmHxmdDkuhm8CZRxqYvSfskZcxUZP820HKfKexOASVcfFxVog
i/Mho/WQXDkw1sdtXdWkq7m048BDc4r9sIgCTIG9XtevWBJLZWe277lK1KfO910hA1MfbNCSZVLK
Lk+OjwuFzqeSAYDfQtVlGpDv83xEI+mZ+f5tAZzYKc4/c7eXtJaCxUBzfrQA9B94Dxo5msl4mA7N
C3lPElc3Q8PZDFDvu1rRqysvaqlEtZRtjXU93eO5j2VG9PBiFrGT/MAwlSngQ7kHO5aTHi/3gXNE
qx4QRP8Iozkbmf5qeg+j3XvJh92OHarOTBcAYWLSpuhmy2FaSgI5gL9vnRJwYLZ7nlO4x43oZSwO
InsSwhw2X5KIpaIKdvTTnxABmh5Kyxie/7gh5/ac+DDTVGvqAhDNaGd8ihZxqLlTh82/Uc9dU9p9
VpvtKRDuKJ+vo9YWPRr1hp4KD+qyWmUSwXwwCKDUfg+MI8/sd1lJVYX1RU5j87E5rV+eJ1AaQrdk
Go3kQ6bjOI3X0uKv7RnzspAH0RANIBpboV8VKcUsww3JOxhZbdWUVJ86Gk7/W5pi6LXdJ3sItIlv
GgUaVZ1TdnSpNMwSu+duwy6OLz9jaSkY9uiFkQ3L1xjGxX12L31S2dDyH3LtxrzLpgCtxs7CJu4t
W+BVUiEY0dqgUJZEVYCixRseTmjXj3s7z9V3zqUJ8G9Gz2BNiA2QG/RD3gXyFgb3AxFUTB7dyqZk
rw6ZnUMwxAZV+oP5UIsoUw3ssWl7UjOtbh1NIvtknFcS7Egz0JvGnQyVKwPlGr6c0ElLoLOETBhz
Oxr4pK0WFvQyQr31V4n7xVlWFLqBJkaNibmLii2Gil0EaKJy7k/OX/uaN2wlnQjpjkTuQoC+3tR3
C1rfTKHlw2y5s6qH+w3YoOfbGSxVih4KgrG13WfCfvxWh128FT2YOfGmbwbaGcbYTCiBdo2GlFtC
8clrDDUKDIJAuX13WlD4w8mUgBS5kmLuoWx1wd7mXHCX/zpDiVZR6g5thFLPq7XvZGZeG2p0kZ7H
m0X+Iq3GZzpNOp5CFU7M4WzhEzyef4olqfqqtz6bJ0/BjvIZzuPU0PBTUEPQUhO1p/JxjiLh/8VB
QH9eZ0d+QXuC44Oh5UM7E+kQ2GWmdZHhZdzxI31d1pkzkVTIvKACY20y9sUIR5g17RI6gakXBSmI
qEUy4XzbqwI7bxqdORozHg5I5xvL4NphW0N9HzjskgyU8UlH2CXqDsr0k9QQw25IcHsxkcYNHtYh
DES0/erbIQkCq/yuVN9mC+X4jnpMQhmCtq4rmlMOpRHe/JK6jrgm3qD4OBexkn62fQEGB88IUzTd
iHRvbMYllGuA2Lak19llYnGLVN9bkSaE5wGvjmRTEED2CHYDq0xjeMJmXkDFA/XNeSNq+zayUPey
tDq1YUFNZjoR/HvAiYiNcdEVczQNLEd5iX/RjS+yWShBCdb1hbMyqHay/ys/PVd+ndqZy6Bqek+/
8FI0Ox/hcjcKiePPKWrcnWnoxBL8kEv02Yf4DnK8QRJWtIDaSgjQvRqVzkvxEZWPZobXIaOAhIVk
IQ7nCIp1iFiuNTsrlXNG9YF3chY3vHMNq/nrsfhLE8648ejPPUgXe2m3hKGEkiku6g7K1tn4okRI
yVJxuVth6ZvDtcvvmKV5K8kMHvUoiHNcQOgdfKc8XfYbS/W+Z+ee/Mn/Jiaou+O2OVglMYLT8Vn6
p98XnTpAKUj66u7VXwaiQB04IEGkIptUdJo/xO4k6bzJZPvPQAaZGzTTwETxkUFDWfRswZ2H/u16
gXCgucS8LNWitc04IuTlkxwOVJU+c9L8au0xyUipNgHk5Typ3lDcynw5hA9Mm3ZcNej1DMmW+QVI
Qka6op2rvm4qkHCEfyZRXGlh7NbFuj5aZtjs/s6G7qFSGaxp40dW3zqxrj3vDGMMITHTqFoHt3PH
mmwlickhN2lbPez3AnCAg7f1qMJRTRdT2alP5ZDi9JqFj8724XjrxIJSeGXaLXjBTzC4Aq9KMuJy
RYjKFxOmZ/rZ7BNo99o8nNszEhZgGABi24JAJfAtf0U2kMdYmxO8iiXKtKGOFeL+v+62/Xw2040W
+Xs6lMRC/NSjTbgv0A8X36FdKa/3V5lqr52KwIeUOsE94h7R6fRQgZpkfOcgr3m108B0SReqz4ii
HQHjz/+BuEUpFMCljDFWSt2fOpFmIkEABTVMrio2dJB2iP+oVTHJZ+OJsBbJOzkzcpwD1DS6crV0
9wUpQN14o8JboHt3i/vNLg3GSDrt0s9meENECHHfhUmsgv4A+beLvhLR56R7bV9UaWizh/Cxg5hK
V9yjIoXncRnePtPuepQFJfvciR7Pz+tYt/AKPl1GiVKr4UJbbLGhGenBKr/27zfaS9NPOMxbq4ij
EZ+8jYDykNXlb0zd/kwdNDprG0NcAFkoBxwjshUMXntnN/9Uxhc1VkTpari7tH9nTLYCS6Adb8LU
ieAjtjqwxi7EwBgPiUjalyUB8Z6cGFthiymKpmGjTJIyd/i2bMAB60G43efFF1SciMLfFTuCoXoi
zpiTf4fGzN+rMlgVxhxdaxbopsHe2zLzN7Ndqlex004s0x0VSgJxxN4N9B0CP40/Ofvtag4IbUhw
bNG5HaXt5OT7FaBFS8lSHH+BOLCZFazPjZFphVINpORPgGQKpu/fKd5qZDNlC7w0Lwyc1tdgc7eU
9H1ebNnpfs9eR2uGUxXoMjSZcaT0U7wJSZe0Vk362R7EjnjgLx1SgJQw91MxX0z1lwSZo3o9RcZa
9jRVCQXl1Vfj29azjm5BK8T5Am9hWUt31hjl9cIaHZrsOII0mZeC+3gjV9kHzt1cOJOUSUjJBLwj
EXf6IobjKrLvMgOYrENv8RAg06rSDpXCxuJG+fQpgDuR+6C05yEawH7T7VdzwvQEdeyqeeRojw/b
AcHv7fGe3lR7FhhEBte5MCLN53rONIWAekHwqsKSDyuxWjs65Zg4jIFSDkLt+/ny5NMv1Wc+M+nJ
admLsmgQwOLQvwAdP0h0vxXCrzWcVRlKczWe/jMpHNNxl7ZELgSkHo9V8ESGzQTY48Gz2gx80Jlq
LCoIhCpbrKwJFPy7XHzn76qFq/xyZu5O5F7RgbWYUqCxyIvzY+HIXO1B9tmZXSUUFupsG+Yt7p7V
ApXJ17XO3+hWAmLOiMs8Rnxakb3DcU/6dWttVXijenZJtKSDRl3lk4sGuFdo7IopVeeeeIZqMFfE
vjfReTI3HKOJMHRUpuJPcMU4QQfpe+/Xwi2hcZiHQUQlAukU1KUsk9hGrjpEIPJ6IDpaD2FJkyIq
or83BFdZY0mlaBQz7JlYWNgchWKPhzIzA8LYE59j/Fp6N889cR/D4cuSNUU1EKXV4ABHvLtzhoY2
QVmEEz0N0v7DNFQoS+h+plJ/ghGRBFwBCnh+OnFsDD4TFaqOfJ17fW1H7cYrnAGE/MfRSS3rcWq0
0ucsTF5Mjq8IB5ES4H57Z1pgswyp0glkX7DIrfeQ5P7D0Wybj9MhsqE/AlursgDhy9zYuLiIWecJ
q7wWUdpDpRsWpBPfvt4AmsUIQnWy+8IEM4fDPxag8nHzQv1plNJyK+/ph1xbjv9mHGgPeCscIFGV
fgDvPkHkC8Qopj5qezudYpAUGLQ5CRdvAbd0ruKCWYdeG2PnsLHyfI3ErtKVJpIa8tYz48RuOGY/
+4Oa2Wv52AIoLO4TUM3YnStC2p0Ub2UGbd5hjASBnjZcDZoirnFTzuD/Yc10SlsLTEUHYhDpXCxU
6R7j2uhhdMBlRQWH/vzYc8vsiC4ctuiNjp7/9b/A4IgbqUcQOiyJUkEK2hqikHFp2oMVMGFNihLS
HWuQrKlq8P+0F3+9ygUbxgX3djMSrQNqR+UQJbkDaTi+oUm24qLYb+IAsEBCPuVtVAEYqcJA86Bc
szS8tLDbZMj+BVGx2HO7wlBMMPZsmIqdTWuM4fmPuZjgowO6NWtrAcjJX65MIum1eKY+GbPltaXs
86sw3ACTIioEarg4qSSG/82vL8TDGmQxKpg2Z0iv7P0egc3Y8XHVGVXkoMIr2O6700L7I3h0djpd
/+6uXc3inDHLxT6PMgCNNVwyOxJiP7LetyqNBv59P68mXcNeAyoKETmgk331RWVT4F9iXtboWmBj
dUmVzycGGaJNbXXbnUfoRIQf/TklC5jAUvb/NL1YKpaGzVwc671DrYtxnuQkNWwcYd47Ne1nF0Mr
cwX9NDSjrA+K1B4QvFge8FjzR1pcx1kOJ7ts4hdYcJJTUNA6zQAUL4DV5DRW0SsfEb4TuUt5NLOT
ieVbTVRkGU3mmupf6Ha/xwT27Znht4W2Y0sfG3XNDzG5phOs0uwZuK0sUvRgLDDOlM7mWG91aUDh
kbkW7ClIVMdrWRUCTsxJ+3COhBtJQJYtmQQpCBceXsLbB4k9xefCRGkU2tR4tpRt18uGBV2gh+nW
hgPrQBlpnH+2w8+oln0aSA3wqru47IZrNE89DLDeFj4pUiLFEaTuyc/Xx5kNFLwhZhwWFg/JR+hP
l8+N7+53uP5neWlf/IN7FNp1aU2eeN1u5/O184PkSSETDRgc3r3dTQA+9z5I9/dFjYFB1F470aSa
ppVL+WQMWtZOpzYXfnquFcTE8+uBwdQp5g6ItQA5MBFNM4npGWvt5MNGuatgm8sU5N8g8qjSirvK
9j632pymTwSfsxCTBpgiv2XJCn6G+TdpIrE0c3EeaT0Q8B8lDVohlUh6b++FiAKDNyNGAhXHkHz2
rozDqxWQ3aqrkguzk06fhwZPllsVwQ0OztwBVhOsFhJQ6nAbxhYOcaKidsHVB7XcGmxPMuo0zgRx
dTIdZin9+6n+CXA/ZDkOdS4sK8vMg9kss06fd2hk6bWx7mZTLjWDgqRVzIbVCN1+Sbhj8CkTxPRP
JGOTKkMiZljjVG64dfAG3HKltz6WhptdjbcLShI/KsNdVvfLf/WWv4SpLWmqJcK4lPos3gt4gDXF
n+lw5SAEqXake04L8waurqg5zInNUSoYYo8VBapj+dEwnemkptttl+YH8rx8gqllP0Zx4MMLYFOS
JRSRghPAS3tU56Da2lmwnXL39jall6AvV/4p/tOryGh96dKY4T3inlab9wXMneu6BYvo4hIC9IXR
Z3jnmmJK2Bydpt2BcL1QomP9yfxOIjYHRHf9YwoR8mGxYG8SYlCNwljMcznZHl1lnsiD7CwDbS9q
jsoO/X56epUUFS+WmVA+3aC5VYcRARswrTjynUuVCW4Gtcf+3irLfBpBjSjfe5mJv9m1y7Ek/Mf4
lJrLaNevMS0tdUjmzxvJZXzY9gTsmi3CDa07/tyg5+7drC27YCol0shswFUGRVl9KBgAqEys9VcC
jCT4wUXf55uxDa5U6dOuIauUVjZTEhAiUWsEMCPXSXywNEGnubIo2/7tfTla5f56Xg6BSBHNCHq4
mbrZ354tGBnSg+ly2Xi93PunE0Utv6+5aZXiV6OaiUewn32pU0oJumOHX1fiYeIwEb/V2E6vmkKY
Kyc2tIEgUkXLV6jYq2VoHlGCmNHvjL5DUQ2w0elttf7OocDDRbNAkHsJ2DS8xVIcx2Qt+idJXJUe
5yWQ4ryluOmec08TOj25Aaj56ySXtflHEOgz1bwMvKy9drQZcvDVnc1dKVeNoyIWJSU/wZAqB2mu
meke7LgQXQLSL6at8lQITmPQKAhMWrfS8E/68/0gDl23FdqQvYOR6WLUNczxa58vM0R+QLaVXhJA
hseigaX6cosVI5TIZk7P1LDNLOF/dmysdc2w249gqETCWFFJ5GZaYTtf1O6hiUCqEE3PGRw0FHHw
Qa/1pdsx1Hj1rkaV3xLsDMTOI0t3eS6gdNwawSIc+vPVMPb4LfO5ZnHifPsQl+5qFi/mWjRVD4AU
KZpiDeR/SkWLmMELXtQ9EgOBzIWoBN+l7Slbufc/rKaafqYYq8Sj9YqREkHTmFByEd0SnGdyfL4q
BiV+dZyTJZ+YDA/TrodUqOQKUcf5186uWJqwL0OqjqmM/CXo4EXIYOVtziJtv9ip1WYZO/rTO0yN
zZDZ01JXIyfjTJk7/ejPnTu/+YJwEHzORPl8ix/9Htbe/PlOil+pecBWv30DH1j4a16h04SgHUeK
g8wfcF/4DKQhEo0Xr14iQm6ybhOAavU+Vhf2btjPNiQH51iTcY3z/p7ThMiBBWixUUOxGblHUoEq
sn3biF/F9gX91J9qub84PLz0MhZZaqiKMsJi6s916bjJq+WNRe7ijGFC0Lx066TrwnEw4oOoydXn
RtB4dZJaOt1btm12m613XN5Bly8/Wr1iVH62W3LoVutnIqsgt5I8TlfTBMtnI2g2I5NHxEwAP9r+
0dCwSMsintrqPLInxYCJzLjcYJdLkRPKJ+0ssP3hs5JKukzzlHO6kEROWNua+w49YQcY1+cLI9O8
faGPfLDZVdGuCN046p6Qj2y9TSUMGrSxJWXTsLqqLr4BuPPiWVxaO59B0ssWafE8twONGQ7JSD1I
3lVa1jp1GZe+yAw47U4IxDNLmhUGmDQyca7ZjKyi7X9nQeELvfa16N9ZEZGQkdpCW1leHAtNAugu
ywugAELXmbWzTzoDLJezPhS3kQ/NP9W27bJ75wahz0BbZL7Qml3wlw3VkJ9rEjLJUHK/DX53ngSO
VnXAe7UB2wl074hzLJj5Tsijf5XKGb5eNKvOStSfx8OJBCt3SvVpe3G00JKC+cIMOzCBNV1luGQ9
x1U931oFxv99PXgPptbJ1cP2iXup/qhvlNj3UM7m0OeuFZqeg7nuj39xpt/Ub4dWR2tJndVXjhoj
X2tKoTOr4tl+0A2ZNGxeAfUNJvM6okBlT6PWMJoanrlgLyva2nYaeDCfLVK5n7j1uYHeejnkaPN1
5GCw/R4olLGNUzb/cd5SLrS4n1w5c1xNYIV0xg2SbcsHMXVGGXPgJ7iNkMLTD4tXqPrZwbv8TDQ0
aGDXMr5XTG4dXwV9Xi8d3L5c+z31xtlkPzFPXPWmJf8L3HrET1+FHtxmDOl/iepczJf0fp9WOnGU
NtYrUaB6mNjPieg527mmFYcPQzA0+qR2V/+xbiqMoFAgYuKE9tz5KXQOvQnwUPOms2J0RuFL8Iv5
Us6fwufNzqnhIYGysleLxzbnVFpGLnyWumBmcJ/cMnL1WGkNR6nVqVsOF981FDKJdJmYCwzpfFfG
CFGKzkk1aXMy9i380KQYNzKcbk4m7URV/JXjvJWcHHfzRaWPEAow2+/5IzuW/eQuYttOqeaRNsdx
sAudqGJ+wXS6A6oBKr33nUqhJWh4sbbJBMl+J0r/nM+lrYjjM/nazQAaAk7fjuA/8KCWIGg4fkp/
XjjlKQ2lG/PdPWpfA+GeVJ4cMN9nAj2BkkJqixkBRgf2Oh+WRZ5xooBOgYb1W3dIs2+vmzqxEWg9
Jrofm91RiY69iLrIVnjjTjAoUqPZbvi90d23hdWKQNy7cYBfnIKAXQyYq+8e5w5rYiwRAAv9rj1P
rZHC9AQr3N/6JolF/xJmn6KRDbQoR+5dKJRitKDk9N2bvJILily/UqrPt7QSeASj/3dVwajow6Qd
mokFe/JKQ0RtWiUB8B3/4mufTcbwGMRwnrQ4fRsqlkO71wCwkdjGZeEkiacVVH5JvL9bvkFADFjG
rVCR+r4NdmY3ASi5OZ7+XMY2ZNZGhGon0eJ5ASFxNT8jvE2P0qA7IX+mzjsOsTwC++fpjWy/RWGN
JhfcIzwagMDtMsyu9dBxIc+WBGCeVz1D4kpBYtOa3vE8DcEYCDljUqXvzHM24Z2D//3Xb+WjPvSF
kldD7bieMMegfU/YoRj7nc59WGvtp7yFFHqXlUkF7mRoNaPfqM+l+lTtLYOIjrkiD3BdW+NYSnKI
H+U48VLCwrThzGi5cxf2ZRU6Vn6wu1F0lrJ1FTWtsgWopr4hGzbOfgTbaajidpm3PeyLxGp2+D7J
s5dE82KzndwGbTF2PX7dUKLHgLpH6ueq70vWAKn79N2Qz8qE5QSN0TR9ZDt92+kYNtlr6tFVdEHh
sVCamnHgGMy1nvcMN15G9gSHpMF65f9gKBtyYvSJPHT2S/FdF8yjLilPBs5kLDyxgM1pWjtr4SYl
m4OXQA9u6URT2FZp0V4Q1R5LL5b4p0P6E9I2EdjeIWBqEQZegXf5IiNWLFvAlafeqX4bIwscT7QS
a6pDA2a1Fn8gZKG2xcUpXnKI1T/iFS+oPdBJFgBx3Mud2C+XGmy2aQpCt1ngA6eK2z+XUpPxGCFf
6bswCUy0M4DoFheNtBpwpTKo04Ca7mlW3ZIfvdhkk+26qB/bEG8ttsCA/UcQ+jZTIIdIUdKK859e
f5GmUmcZsvSwwQr1txpYjeogrHyLN58XtWqOz5AIGHJ0VF7PKuQ4QInnhl1l1jLC7jaxYw3+3UK5
JanVDmwZLXYJ5DIkoUR0wd0X+l6Mmz0CN6by/oczTbkIFnnWixSpHLDUJmRQ0pPEYZ5dC6zNgcWT
RYq3UF7pgyjtVeYsMapDz9zZ5cv/2tzIF9Lpz+knx3R9OJOXlYFSjdcE0HDY4dgewhKmmvlxSS0Z
h3ZxKJJw6V7Aj5RkyEs44J7FMJVsumcV1zKilOWdMXT3B/BueqxyxhzGMmrlVeeM5eX95+kkR2hQ
xiiG+aJIl21eN/wC+I/t4gwv1dvD3fVrp/RgLc6r7zLkdQjRhXEwsRBiS+LDpjQE3fdJSVDl0GCf
rB/xL87ySTHZSKNh1I6NUz/+nV/QQ0CgFkowV5+AsscDeaiDZpvuJW2FpYnfTf2l4wIQuj+qVlj5
EgGMTGRNQ08tROcI07UhSARx3Zwgoif6nwwP+w+PEW43HohgpUdSxooANzEh9Z3ChSoK0TVh3wmz
Rw0G0aY/X+wTHbFCB9eHSp2OLZ73wv7XtfPt0AtsS9Ho3Ao+MlZm7sM+hCYaDFsl8VmscRxqllbX
ibrTf7dWlvN9+k+h2UazAPRbfMoG4KDBN1e5IlB5JNg19PVQwIsEWeblttui/v8R5geT3y+IG/ml
eclFOTA+aU8E1ALnuZE7cLi2cjj9V24RbRiU22qOMNUa+6lCVURrf4Z4qdPdgRV4TwU0Vpy9J5fl
xbAhJi2Y+K1KdbxPYLSr6pED6ykNd6oMdOuV+ognTJ6jg+8w5p6DehnK7Jk5+xG9XnJbSWdO8rGz
DuVw54KPh4ODH6j/k8vHdCsgImZuR2uyKpsRnxs3Z0oSiX36xOwQK+VXDWi+iz8TI0zh8Vw1unzY
rdTZo/sRL7MaG2MtHAazJevjFS7QNCIA7m9Uq4ig60k91LdWXpopcTWuqMkx34H+tdi828PgcLee
5dqf5TNp/Pk3cRDEkMeRN2hbYSrIAlnW7VgMO2yl9n5M/r9KrtFXTzo7yU7vLQlM2Jubx7PtlfzQ
jWpaGvVdlJk+GtShsP6VyVt5HgB/34ThQ6fvf1sDmcammtNR0tqdBSH5E2JHC10e0e/v2renLa+t
9dJ5QIEQuEk8JdkKZnQMevob8VmpJaTb2bmUX/IzbJSEUqu4dVmz9HR2oR1EP4l5dLjbqNXm9ijG
KHqeYtCbfFmcMAJE0Z9i8GRpLl3r/ixBDJF9LPykZeCMbZ4dkBJugkjeEfjBm/Qs7UOEQeKYZGn9
PCxltivdSkKNQtRPNZpLFS1E+bIeEHGXflbP4MyuVpmcwss3KKJMtjoTnijFd+je2fHJI91TE54A
sMWjiQtLFhyZrkjiqgz1Y0uF89vUMKUckk5XTlPXMfk61FBOu3iA02AnKsCrgU+6ZbqU/TEkqiHv
8e5YmnGu3GOkQrW5Pw2IEQTl6oY+875h0cWzAgyneXKlVso9fFpdAu1qbwthnOGvzSuZ+cn07sZG
tcIdLFqXpLj7QJ0WrKUVjBeZP4o7U4aTDnQ0s+C82XhxbjLdXz8If3JbjUrhtUAGONJxtfCWx9my
JuiuRNEsYa/9EkDii4sXjUkVaYAYV0Xo4ZpMof6FB5IGM0yg2sbDvb+R79Pd1e8p20x3q6XJfLUu
mZpIQHpvMKqvxHNsDzLV2/hMbdzni4rq9Mg2wyDaNWDwP6gIJ9+lkNK6DeYc9uV1Y3Oeb1qVQyJ8
5DyhjQB/8mutUTv0vjyy2qrEmkXrHihIwvZEmm3uDKqoK60l4vhicMry+ETysbhoIAIQ90A1D4eV
3wk7j9xBAjeMa+GN2QzxNYWs1adArlCtpPMtoeCA54niA928d3YcXQczUGe1XOaTsh1a35HeUNej
Ly4qlL8bdcvp1SXhMF+ovLHXM6JKHec+yORlSHkdZXIvLTGaim6R8tesdA5I3YGDGs52UgfJiAQt
GtJQ5dXLZl2mjKivCg2WaAocscQmBqtYISod+dNEinaVFvt9WbHYmp26OHYSAd0mKmnaPj+aNG02
r/h8BnZqk8eb9E0Gdl5+hR4XX4uZH9DT37+E9IaVRUeWT6UVGuPwYQyOXPFwCrLJYjepG/TgaUa4
bi2QHMOx7p0+m45G8BYP5vxGohOxXgFETisJxo8seWnYeRrvpWo/k1Q/mn3stunoF6h230eRg5nq
22WoM0/aWcUIAYinhZ3sj6hXILvCfYo4dbom0WFetNDFBuoOYrC751Ow81nwc9cxhDljiwCgl/Zh
aUW6gVj1D5CHnSs/e4IDa23aPxPM+PBJ0P2s/LWKmCuaMMPbHCSaDSyQatGii6+WkzQFzrgHZGvn
jA7QR35tgPQyrpDTS4BZ76EigsDu2ZBw7mGZX3QWAZyZnnfdHveFVSVFoTVi6l3FDdUeQ9kQA28X
QzszZgOneEZUkWmRpMd3NWkK+7Cm1AhGZybRHNrZQK5sRUXvPw8L+0mySpgLC65YOUkeoak0HQOD
wI8vJWTbZyca/dRfTWNj70DOEzZZ/DuLYbMwz+2wgEhLsKdMeT7Y0Y+NZhPAXA4CFbrTdcnFe2QQ
+9THWUi+eaYs4CsevGNN9NdFNAFZE5QKg0HzfAWHXkd5jkkBtdRESNMt/DUUTVaknLedfOaqH224
YjMhqFFnoEIyw2S3xSzHgbDjfh/INRm9gP6XX5YzxC7woOcSlTM6Bj34ekVrepu1kjaTMzAWxM5H
4L4PzdqL02GgwRtQAaJjoXIn/XjgtbQF0Tozy7lv6DcB01i1cgdE07MHsboVRocLSUCSGjAjUyuw
qcMLC0MLoFBpL4tCgBcGfpbgGVRg2/wdeivGKyZZ0M0ycNcXKOi9irW7DYZhZIB3JZduShbt6Ym8
lztbhIAoA3QmpRUuZKhpc2JikVC++A4yd4v4tXCI1LbTPVLaFCgw+e1koKX/dfy7OfHhfV2uD45h
w6M0sTvUujGLwhbIlosPNkmpLppB7Ajbfn9SLjt/fz+zhY1AXh1N0gS2zozm8VMOZV8S/zzdkb82
ipDdqHKdI2VJuxX2TlfScgdI8NSg576TG42GcVvoXfOKBeuQcRUYb6xiIOe0+bipyv52+at78i2Y
7SyAFwPAqk9mesaf1ttWc+uz4fhHMfNvPmrcfhnZjeAfqAzZ1fPfPzkEmNlDkmaHwjMRO+UgdCxR
1NIl6GPWS06NXPVLVbyX5eldsySZ5GyRZfiokWJZwysg6dNOnk9wyMin7qUL6T4sYPYasQkRwXpr
/47Py1NC03EVfOvL5PtbVAh3QVGm/6QstGU2qSpFqERmGzNM8kt05j9oMvUeN3lmIJzSegM/sxCJ
KnkBoVUcpI3QwxSdrnx/uglJERsAO7cpsDZBve5+fLor+yTIjN5MuFGgDrCCud9WqP1j9k3MJOIF
OwyT/ZvKoWn/8q+uGd6YqTgu04DGJGW4YzuvgHHG9b6ovDQetnbmtqcS+T+PezyKPG2eNe916GwO
GGQDCGa8PqRtipTAw3u1KnvrjgeLh3XsTuOOhjs80fxnTK6a9hrurNyRQFmJ5Jj0aBtyWyklqsq1
d/srqaeuHCsP4I6qOjceDTkKAsKkzW2WdJVuATwTcufayd1kpr8zqyEcpEL7qiWUBAS5dYZ9TlKD
m7PP4B40BSJ3c5JN05P50Pi71kLCSaMlk4oOU556mq96qB6WSJamYBIJMhkW45Z6Gid2icCdDLrs
Xd8WrCVy05fByQpXVOqEuS2W49qBklMGBDtjz2s3VU7uH4FipUOTjyaLlaSGfP3W5FIjlUpmo7vR
+WwhyRju5ImXStp42K+5i7tP172JAUacRIbWLWduE0Mo10W7zSklCdSppkNSwM654qmup5tEagl/
tbLdh0/CyXFhZLHEWk/dhqUrVQjSXxbNnoUZFMUiNDD0McfZYENuAZ5nuZDmunmuNkM/bGZ6K6dY
XZa6bjW867alUv0mVRHe7vobwDjUjWM0El6THtv8BgHCIijJrJ+lF+aValivamtN0gebYi08fifx
Wmnt8zhK9hbnTmxWH/z1GxtTVJNteDKQj/nWlorjptdBFETTa8ziVXlJcP1HzGdya0RMIJxTHDMo
a3r90ACUXRfqMxBmEQPZB4SUutPM0SjRGYcXhFe/X9ImpqnBTwAGcnyBoDa6cet86/03lBmhvQ/L
dfVh8nzXlt9KHSu5zMfJCtyzwfeaFuFfY3XbKWa2LgycRjNcoqo6sbT7FiCETt+suhw8HjaXkO56
lyZ27NSvCj+U77qB6PMY5Fs9w+jAKTZkT6J7rcX30ADwaTn/SaOZUZJAsTcKRlWBBX5EmBJzrcsb
FzHOxgw/VNJ0XVsJseuM9y6d6IR0RWEXAfNnhnsb+DN15ZteRAhpqfzpjQ5US3GFh4eo7k1rUJUD
X+E/OuCKTpeT4CJdPQ7HoOUcYnBdpmJ+8GLB3pAzM57k78cBI03CeDQ5IDLfpEo6MngxgXwmgiQu
AQaXKVmfblqVX2d8HqiUMsmwPBnv1avXlPGsOW25JsHDvnuMLIc7ALILWqPbmAQJE1OHGaH/SyXi
fw73Uluz4b1m90n+llS7Q4LEGLTiWhOeo+5XgUgpytHBosYl1HGrXdavAAdQL8l6PLCQmGhtpDqI
kDipV+uRzkmv5zBVrm5kqZM+jiZvMQ5swvRgUHn4MVjum53u5KaE+32pacpnmFuN7zF7HwXVQERr
cf/caADX6cz2NHTBGFRp0J3I+MHtTWCenysyru/14AyUn3FcHgYpkkrptqTX0Eh6FD66rOcK7IgU
G8j10yTMFjSIT65dBm8xzATbRFpiXgMJj0Z82BcuMs7DCeGjWGVViLKrf3xNyPTooO2VWscMFhGS
Wtm9c6dk8RU/2fFB+CfT8SOQNlSFu4Di03+dTa9A488eSwzdPgrqv2sZI6/Mq2HZjAJcBch1cJgg
BSkkZvcGiClDaOk56yxAhN45XwFHSShzruxfeKOnEj92xV5goFBg3A5w1OKN+jTGYadlLl5JesGp
s+O+H6a5aUE1vT2UmPAVY5W4+2oo6JLL9Szrt/CJ8AhVrb66e/VsD+RfZmV+ebnZrTdxo9p4L17+
vVsuLUGXWDWbrhtHvYrcHh+WlzXtmcqFbpSm3ROv5tDEh91Ch/zW3zWuJM8MIGhz/p9kuxhOV/zR
6Q1Ahv54LKTQqMFTO6AHPXpYT5P76Ydg9aQN2XJcZXWV75bymmwjz++/bC8lb/H1NHCLbpaH2ctZ
ZRFfBd5vhGKoUU1nxmJuEUNpPqtwth5JT3XzLgi7rHOh05oX9oOZqP5vFEH9rf495j0MaFd3LHgQ
/Gq/dyTA3Ti1FACduIwzV7wxoW8+pilX3PGQ26C7soZwpY8cx5XcUJaeDjyjgUj2JmGTrSKEv9km
n8z+t/o89nnyXxR9eX/iqFXV4nLPLmFJvQbI4XRSRBEDUSX/LUpigL1RDifAHuyxvsQf0OXl5Z86
k8YZh6pOlQddEWu+H8dgQB93RRy9X9SiOzTvZ8iyQVOPHreXv6cdF4liXVUvAQO4RHZb/mQBg0Yg
SpOo7l7qGy1NDAYZSGB/qFKV81xb5oqoT1pKSkMM9epaqlZ+s4th9g+xD9+EoANJ+4RO/kstIzZY
k7X02Yh5s/hX33hAqNKgFHtD8p3JAe6vzCFh40+jjcFFs4ngCFKZe2ILr1BvHgQIzn0mre5Bt5Rc
nWL6QwsZ2iNnh1Yyv4Up+xIiUr7mP487BAAtcHKVT/1MqxQazdYQw6bA1XWNojQnNMbXojhaU+ou
AyVqj2QetCczu7Bl3P4Q8z6O9iD53ut7bObsVlMDQQ/vXGddGNei8GaDx6qkB+bhhcWLVAYw2m1a
yL8SnXymYqasYIv1VMR68o/+ZGfms0lw9Utf4R3znUnsk6nFH/QuqXhZFU50VCmq761Z9b/nU8q5
xD+5emdx7NjSQYCOpOvnUheu4dH5vhu3vuXiAZGzMsYHqjd7b8Bl2qei26LrwFpTp0Pqm+svr5sy
ZUaAGXgZLIiWz3GpN/jNMoTxPB49PvT5Qa49csW/81gD+xlkY5gE+FA1RrHi+mfcRjduwyHu7kyC
hg4waibbUZ7W1OALBN1S7ubmeryDmfxT14ScfCLufDornDYZodSIM5dFCvNwIPGRNbAn9XdfDgTq
66frwCSLrDqd2PXxUZ3ukag1PF5zBCawhjW5a+Kq5Dn0Hr2PhYljgxHwgXCMLUxPYOdkU1tKL6kq
LpuU4UAgFFoUKSCKHaA/F+4hOpLpocHKTzP5rJvjPuc0g7PJ9neWZk4uuiLGsdQjajd5IxA9QXv+
HxoEeE3foKGC/kJtZzez9Xy+WUvEECxlt3onQUsI52vSjinYgshY43b5v0hGlzmzs4uY9ubXGM96
4wllJ5Wvn++wG89Qjogx3Ylsmkz1CNHFWWRFLJ2umSU9TZeJEn1+JYyZM8SYMGhQJVlJILEKx1TA
L9AgfqquE8jmY59BQVm4BKSB3JVx45wHd27xCiUgQ41AColNHpn238SmZ+eUk9FI2n4+f5yWjIlT
l/xxRGvB6DFjLXC2eTPyqkW+R79BAf2uI8rILRwR1xqe69aYVJiJYlhLRp3PdSRPzB5YqyuctdXP
hgEUbLcnNtrA6ddibP5Hyd0gjvz9sH8sM+Bdy1uLJj0bSxdF7VrjGcRkboC7eMeS9N8vUrfviJai
coUyM508d5yk/kf37+WzwQySar5UmyG/yx+znSzJVLpmRHjw2ht2KAObGvKZHejch1YcJgIKIPbs
MxDQYkTmO2iXnza9T8q9JcPuPRT7y0J35K9PGW2zBfveGuaLRtC7cMMhwrxQm0B8A4CeMTua8lRn
mwVd7Su7YRTh1On/IjSZcBearB5WGtJ6dJ3GQF3hlyow76MqjqerlURLjKmcCuGd/dECuTL9lBd1
nNCAo0GRjZRpRCznHWcwobvMmly88Akks9rgOD+Px/TdHIuYd77hMuFHFFse6ATG266db9URgF6M
/BxWVd9LVzhlG3HCVlYoFJhGQPHTJZG46BAEqBMqrLO4AA5qCRTDwOHRccLPIXCwAeN5p+fcYgNJ
mI4v7VDrUfu0cFkxaSJMbX5SE7O+MBFI7kO/4P8VcZFa8TFe+mFd4VPSFqpzHUjan4dvQuH0RBzL
+2qT4iXUmD55Mt2aVOFFDj1RV7uIDmi1G8Dzjg2t0d60zwzDAoGjT4GLd19NlkZ4Ej/o22UzMqWq
SgH/JHwjDty3dWZ5C6guhgs1iiv+XsV81AR3KxqGelglR/N96KwA/b3P+r4dysa1xNEGjKtOPw1o
zdsa1PzNHu3x+aIyntOY/6KjMlfoMAzZAk2Ko2/j+RIZRUHXRoC9SbXBqMClcBDrYMDE5n4wFp+O
wz10Mqcyx0Fr559Z8Jy2Z78iPUG6qjjTlMm+boxiwx7UVPVv5wJYEf7Gv7UjmjwgOWdY0Zdna/hp
vOZNqQLQWSXpelG0nZKruX+SeASl7ItoPlsZARiy69JYa7lGOuNA9dfMIk80SNCDIKyPYrFpsVag
ZgzrC03bH/3OFs0I4tvD4leIkxV2N+WwOTKZy6TiiDwqZ5xNAJkmKM7vkOEb++ZDzfCmUnaBUY6k
AJHzOtqD5ehJi25nvVnjcGtYtOT7/nMqFyj8YKdN8lCZ6dfsLOMoX5adgoDg59RgRIGUNZSdZhHq
9Ae32jpULaNT0LJwo0uDrbBaJP/DMJnwhEVlcW2QVpUhSU0lBmhluQqXSRuVbSUYp6+FYLAgWj/G
e1WJlGKtysNVoFHRBQ2Rfh80px99AhbCSk5iRNXoVopL9GuiFRCdDEb/gihXsweSW8jWDwcE48yg
cLOHsae9EY7NqclT6ylIXeEmNAivsC4y/E5U15X0P7+fXLgkSE9RiA423ItI0QovTlfZDjiYp1JI
UhjLVE90e1OeDEljNFPxrL80NC/2gpIN1sR/HAh1EUyAGHUVbVUAX7GC6cCwHxh8tJVZ06MTMJ6E
eMIA31gzFrChpzVeSdVQPM6ffCZzpkwB0ZIuF3YzSBSFNstEnVSfYP2tL1a8HbPfvvooIHj5pDQH
2xa8QlrLbtQuDoiF7e++rasKacONm2EPIdLpsy6USfCGyTwbsevPW/AEdVy266i4W5CoOwzAxOxb
Sq7KrxRAS6ndmtzCfZTPM0qIrFEAdvdwhieWMYDpo2vw2QJV8QbxKYCyReXqHLbCBCKUew6jkjss
IAwKRrSJjl8LGFdPjWx8fm3IAMKo1skP62gcSUz5auh7m1NkCe46IitHhs+TcKTixOB0T5Q+dE2G
78hFvmz9qfyYtG+E4vCgj8/aw5FVsKjGeTXMVpkozuBNk6/o4SL1ExQBzHo1bRyUh06ZUTa7uPss
4Hb4ujXKBn6JKCj/EUjTkvPnBGaxD9C2KgdJumymNZGvJbm6ZqFfTULzejUQlV7v8hBj/h89HZJ1
2+u7zuz6VVLnXSXaNvtPtAfOcVYbSYf3yeJVNJiy1d6lKCWX5Oy/zjmRYyOlADpHEmy0FjR7xaAV
wdzm4sqfXp6T5obZXgcLXNvFDFg9GYpiDvW82oOl2YWkLLLkFQ1DJMS1mxlHVspNZMlu/1ABydH7
GeYDTYKmGTekHg1g6GTydwTQo3/oTZW1WRNHFXRKZx1yP0kMinVgFej0eD7O/hrVfpo4FvLpNZjW
+pZRe0EM7dHlaBKTfIfxYjlRPlB2r3BUxDr0L7vLE9SF5SMlgIJ3pAwqwZI50d40hRUIUqMzndpl
w+Lg0L/X27hmLWpaTmV9nTjfQVfmMreNrPC2KwUZsxzZMRmSqOfLsBmzSoyzz2fdpREacp0Co2sD
YJbkieVwGZ4Q4tyJDi9x/VVshGPkh18plIuHXOPZLG2zTrvA7q/Nc2gaM/3RLOJOcagNCIxqPl6l
6Bl2DJkY+XecO49WkmZVC7sd3mpLodYNCW/tScfoji8L+tQwyHblu0tQFuKaRcxHOOqR/zxU7506
98JM+YEO7Xfwm+ssCuyfXfl4uwHlO3jsOO7qWReD5JXywQTKj0h3xCxbJokugnW/dOg2s8yl2HyB
zsTr7YZJQ0PcxRVZEcswmzPxotTXptv5hyJ1+8HDKtF3gfTbZIdo2NECgotmNhe3qoFYsgxpWBhW
8EdSpnkBCZ/vC2gZLtOhJT7CRFJNMsUvcFu4bEqYTuIYkQhEvUtu83BZRUVjizsjgwR+wn3L/7JM
vifRq/7JeU9SlAg5/EvnFzDnJ6vsKLSwuzHVHc7UYwy9d2eI/M3KdHRrZVLhEFnWL+XUyea1xQBd
Qe4FsB5jo8dgjUksTlzdFfTd/dQAbPK/fClqhhrqhQZHCiK1diWzKPlt8SnmTm0NkVcSrKSPS3Vt
liMCm0M+F+ysRabAe02kftz6axETH24ixyV9Hc8MOuDufOw/GKNyob33X7ISQoP+EUeNqq9dQSqe
ho7LRwVITauGpb7czroN6CSZDysjZ2MDPs1pDbRPGtKcVJm4yUErnhnDSuR4FzDOCMpyXO5Eh64X
oHZHU0hKMjc3XpdH9E2jL6fyTTYqtnAM50Szb2JZFmF416MaJ2KY3mB+J1eM0vGiv+6/3QkL988a
Ze9D9zepuRCXkKpOZNYXrkvVURUnx7ivODgh83DzIEbF0DLPWeudiFB/nFR3fHtF4VBiEip8lrZL
M55yFJ+K3r6p6idcm6ypvngG1RYx3GpEFkc4EfBT1EdsNBoMYXdV8YHWZD565dP+4tSmSiKJqQg7
VeY40e/cbzIWRqwuWqygiVV+UlbrzoQrDElFODJb5wanX0PTSagrXXznLiLvZeIaUxcHPzu6hdpW
HTEVj4fOzzySzp/E/94JAAS+TR+iDDYMtWA2DIQY+NT3JZtY5J0R/wyqnP7AMncHsxu+B15WM5G/
uttadhPYtCwWnxrM5rqEOl5gklPjP9jUnvj6hz6+qV0VwazcXx+kP/4+jq3+ka/1m48yg14ABXMx
D6WX2tQZ/YYx3lP9sWPtvDemgqAY3ZU4r8ksfxd3yWwmV76bJ5FuLm2ZUp43OV7VAEqU3nAqZ1x1
wuyzSj1cgkXS8b2VCo6QG/CGYDZJC5f3kp5/4eRkl7kanREgHtqPt0dwPPK1ehtSe5aSMrvzBHKV
1ZJSwQDZoG0mVuymdp9U0uso+9K7omBYRpk1flDtq/NvtUeV0b0IgEFqWgpftMChmSJBrsq7jXFS
zLMfAs4SgoDNnwpnjv7dDCdkkVQzOp2ygYnWygZkBpPqDLXqTgqK8/QfuJ27L/0CDFSQKX/eCpsv
L45+lkPxNbcoBS2kV56ZrFcC5NXRoJg0U10uT+HpptAMEIpd5XNksGFkssXEFHvEVLmNUbMxn70w
rCJWzUVFl8X4FZdLfFbxbpUs8ILdKhcgnt2Cc7LQ7LEI1aXZ5I2WzLLsFgC13wEP53i3GckoMgk6
h5qEg+hRqfiuJsvBOcPv8R4C6A4YdDbRjbjxRboLHgH+KjrZ3ubyNo92us3mNRWUEm5ZW1umkmLv
RDeOEgH0duyKDFI8/yMEuOjR9N0pfCAiMI/XB27yjoiU87yWjVxdTbYAGO/zNjKUpI2YWEgIwZG5
Guccb5orLKrQoskluXn/fHe+ozj7PIecwXXbByTZ6E2v8RkbuBVJeIKbnVMRerJQD0GYBA/V2be4
f6X+6TDatfz3wA/k0ykh0gUQFcQsjAWptcvoDqoJMeC0cqxp5t4DujsYwjyBrTw6+E8GwAfrYQ+M
3pSqRtzoYynMY4nPBuphCFwPYNx4tOmDIvYAVeHOsTMetWsOojdnkoyleL34P+bnPVuWddJA9LxX
WQrQzNPCzpX86qyrVKaO/lfiIt2qpEXkXwBCN+4xnpHuakZSg0Kfn6RnaS1C0qY+qQSY5P0oJXHi
CYY5NwcrJ1AqvvnvOmrmpvEkB8g7qiAVTCP0f3ZnVg3GZ3tj2zexZX/oNmHZnD2QNtLIPavmxDwY
jR7n8lcArD82AyGtV5qGeqT+ai4emWiPOTsbgnfeYzNRXOFTxxSZt/JtDyvMI5EAk9mXpHwU/vDr
coAQmKFZqXtsj0VvtmDGCiThVKFd4AfEZaTUGvt9dqHtPTqt2hY+kNLMGorVACuqCRZK2hkyUV/H
aUHySZzcLx2SzMLAIinDgjRNuMCI8yDXvp4UrRLFRk75k0rDBDITXs8v7XDkWHrV1+3MgTvx6tnI
Eh6FlJS5SJCw8NAi7udGgGCRnfaWcDeJSfrKi8ykFb9sPtKu+NpLTg7CdWGmxtGAL6gBxUEBRATk
7VI0mSvGUkiX+cOxIRBk1ELM5BHvqxOMuEreklYb1ReKh95x2kyylxPQ076+zmaKAtLAmWyz0taq
RSGRBYKiki45ZdX42wWQQjHfnORGHhP6sUESsDWwl8pZH7VhzV4CInipzycvpw+VoQgdeIEOUiIJ
eFXS5Uf9EJuGRgK+TxEz1Qqn0C4GUilP4bfgTvVSXwwd1zUHuTEMYqeFuHkEgGRrG5ddUYy2VbYd
aNGishRK3l5NSU613xQhRWiFKS+FYjUJ0Jth0LF3O/sX5YbjUR+El1qgvjsQmI75dRlBo0VvqfMp
VdTbAnWHXdX4unK3GMaBcUwSmLJ8faJfQgSeb3/ZmubANz3RNV0If1s9yiVrbHLBowUAyKkyhEu+
HqgmFVl4NLGBdgmLtAZ1dqY29tWNIv5mHrVF2RGc29RRjfFPu2D9CRYpCcooor8v7k/upP++MJjv
Su0tYbSxd/SQNt6zoc6pyNEugcsE/EtPqWP+o5L8Fa7RIjjAPgOXvEqyDs228IZbNCEdwKVS5jxz
T6CuTzB2jxIJKns/h/JMPoZnLQM3K4hC5PWs0vY++4c+7CFlKep0ILFAW2www+G8CKGjyQQo35Pv
DWTa6rA30IxHLWVYangQRFs+DzJuQTSYyyNqJsUl++CjjRpmrIGYPSa8HuTZ4+eELY29xaDFyu9W
e80I+42q047uG5fAli0ZUk6ycnTDTkVGlDobdw5pTz5cFczf36FZAx6ZIMDi1RK1dQWvbE4YoEen
GETY4b5uoaXiV1d+yjQu6h2FIHeOJK5qLEhs037MDGPVMyUHHWyauG5jNH+uN3QGvQDo0N7SpNWk
jZ556UYkUH7uKb+VCamDML6GmrQvvojUfURbBy8qTDe52ZOC+JvCLsMIXiTu+LpehYoAXicaCsE0
oc59TfruyUqj19Fg3KG0gl21n18Kl4SUy+vafSqzykzWxF3dj4SZcWiCE5TX2WO6h6+MMp+sH35a
NWKNmmIKpGApNddk5b30Rv0CZ8LIb1Ckat73s+iOWWnBUaHRHz0T8JzrzJoFHhGGTOEtTw70O7km
LpsSWEyjK+uQmKwXwfo2P8j9G3qHWcIPD+BJf4t1Ky7pzNspjmzfblkhoeC7u8ilvQrOqDE6tp91
O9jMFQWVO83w6LN3YWlVmOAQEXxP1Sutz76R6v82A4bJRdSMaaNOj+nNJjEPdmEsPqOPwxkMq45f
0f2wq9+QEEQPoUs8Zvxw5YWooSChJkNBMVsDmJjMK+s45NYi/ApLWPPSH6KSvrlyY7aP2XgTlhCm
NHC/6DlsNAGO7VIg5TkPqGIFJ8cpIAUUwx4ULbTjLwznoDflfA/XIXl+ueLIjcp8mxVxmYEmG0d8
DeEJqefFMDYgiIKHzmNXcAZ2iQMMuohd8qy04xm7UkuaCPse4fJF3s6G6aCTiEOFUGX9dKAsXMAL
svkNVvdRs0qsfkn0SC9XeP9pl1un4dvLmkPNmUMyUUfC+DK8QLe99UxLdMpeTHuRWhlnrUTSiQBy
/KFyJfR9zRc9I+wW27NnufKXfqUPKqBj06ZEJKhsjDtgAicBg7AfY6XT4v06+THpjv/nGoJETcv7
2yoxjI39a7j23DBH9/Y1HayaKNWYcb4vu1wVZZwTd5wcVwud8IRuXIE8eFHiPL3mugzYmbMgnBoK
nIzvbHY6evXjjXpaCl0+ZLlseKNaIX5E9p0u0XzwL+A2CuKrgl8eDewDv28+dgRKcB9Mi0SdIWym
v7SXOv6S450NIIRcusGBgevq0zh5TzmU2J64JLmrjEuzHNbpmvvZepT8MX9GpHqhV+A/f8vwjc3U
5t3A/ZejR7wDoqWxTKbhHt7d81W7OTsRfJdX1N+Ga4sV81yq5uNnXWX+NbIfNqhTTQ0F9zc1Eu00
XS2iV+lC8N9Jc3xh22VuVlhYNGefzefzPXaT2tPnM6b7NCZCgcZ9nUrOkRn1VwD9MODpAq5SHeg8
UcCvHIKZPGig9KZxQlHhrqL2HuU3RBq5VvA9iji7E0UQdNKjzUsHPIwlgyXNsuUMgdr+Ij6migr2
uX0fIqOd0/6wmNkfJJfKJnxMxFTSHymVLD6raiEQjjDp0tGwZ688V4FIAC+9JY+4N1QdusK3WsoO
iEzcYYiUjdjNJocfTwhV2fPtca+WMnEgnhWojACo0hAqCnVmkMy8ItA3X3tW0hjI2CruLxxWBfNU
h/8MAiEqQc1SpqcXqbXettDOfKorc5DV/FeDagh5TFwjAd1gxhqGwRmpxwqcDCvcSQ6iePXL+rgl
DNYrbDl3mpr3LXqsmLzYzyAIERBUsChID5Srzxzl8nwJdEDvmvDKxeG4C2Q4L7fzf7cZ18qDQ9GY
9lg63pQPsUR4o9fWnfok8WKRfBprEoWO5MA9brMnBNeudEZuiRolahx5+XmtuhMknJOvwui37ETD
eM/YO6G/AIZUnoFiVkfnWQdNNuD6sopSNlE6HrgC0TeLIPy1Spufvttc9E4rtgtwP8w3ER0v05r7
soXtjg8owcs2qyacT1CCLLL983ScpblyGKxynDknYMyGWH3L6uveiWI8sVYwK9mEqiGrz0hVkddn
Clr99RS9T7HRdavahpGWwl9FnEzZ6WLDQn0H1YMXF4hdqurVQn2QVlIJuRkXMciRJPCFQzTfi1sf
IL3EON3rzEl52/B+Mey4HFleJAHGW2D02hTS3bE2uW4PbnJMxTawO0B4mJP4+f/ROAD/ImmXI5Hk
9WpWjX+EgVpRrDcGGMYGJdRoLb3+FpotuWTX7Ghgy1OA0LJmBE7hdeJUaSmt3QkYSiAambDuJ7hP
ZEZhvcimUc4F2P4+6gky4kAxULAcLElyhz56m2pu3Ey0dfXTQ0RZ96rfbqLOtX2alytisHk05dqC
a9XBLXhAPc5Y+iF5zjAk84xla7xz+S4kdCB7AK4d/F8exWjOfLYAt0GOChjTskCbDmbQvNawmQyk
h+68mvdFt51U58J8ZSNAI8i0avvA7lKtMj8MAOR9Mkpnt0nz7IEizBrLbeqTidS6gLBnACe7SVn3
XnhxK2FvZJNNCOpetatVxvKZF8T5TrvwokWm/80pnh61X53enkB7DMS4xWdG9T8fnq10c9qHyYHu
ysaTnZBWUN/JB/dLsavVjpM/YmeBcT8njRGU1a3+gekL2iTXAwC2vdZ6iH+p8t7iyM4iSkz/2gbj
3bi7ixa6HyYiF9b/xRz/6SVijvveW8H7cfG2qNXEsiVoEPsHMkdeh7G8rKbWH+Uer13ejUcUkmfM
da+ih1HMtDK8bj+HnsHkSzMOaPf3AyooBGiJygcmnTkHYQtS+mRGWvywHvKLHbL6xvnETh+K1LiP
ICAVdZHIq2jQ3ji3sNhUKBEoKa9hkJUZKSCFppjMbssIQK/VD+kcX/8rwB1KF9PfHl3nJ2ocX4fk
McYy88j5yGSEW/n43yqTds6RH+N+/EfvAlXA4+yKpsxjYVnglpz5g+NvOgIDFvdKs2vdCQG3KXBM
yJfm5F4t7GYTnpu8Ggl/JZmYW50wD9hKDu+eraZWZw2WjPk82cB9QDsjEsryeSrHMV9H1wUzpJrN
fNT7cyGJNqT0GdGnu1ZfZB1KzCS7/clTAuzhmmqVcCF6XC0RGm4Gz+zK366FQAxgP0qEQtGBbo9C
hkI1naDxAZy9i1GqunOyqfhJy9XMC0+VBZ8KVdvlsxrU8rG/q4nuT5tP9wrIIMvyXjCr9vXzw4ux
LKhue6QWKBLHm0xlOmSDpsVYGstdoeTe7BGpvOKC1MXMqIQ0QIq018v1TtZYcpnBqaCsyrSbYnYh
eAGaJ9jYRbJJ4EommvuczUeijGlF20ohWIHnh8NxT3d++sIB9YN8TtKLdRb2tBs+loP2BofvOBR7
sGV/mK4F2TlSxYO73h52Eq+ddzscM/yN7Sd3LxHLjoPNLy79p5LHRiulOJtSJjYL/s3O4zs6j0Fg
Z9kuPOXwl0FP610cxw47KN7FwxqFduxNvUXjUc9TsC/IpX8NQhdWfrq7hgzdpdXgTfe3luIN52MD
YzuMDP9y2bhFUOv0EQ1XX9qyRKLS6zTHM9lsC7Ghu0yubVt/B/cvpFhVCJLORfuOitPJdoAbPyJa
MAvMRSKYdDmkzktn0y0cUuiNkANfDkZXyh9HyTkNziSH/YWPqPGiMlpzSjdvc0xzcbS4KoMDjzXB
Zmlrl9M/+K4Uvpc2FS9sYAtwt9785lK0na4aFwi4tkXReuC6XXgrAqITW7L2rsOke3JYNWe8WwYq
nh0F78RH8CwlBohI0xsLcR3RFZRnz1AjRVvSQPg7C0zAl+8DsckJBoX4mP/b5Q4GAq+jxF13WZ5l
0egtRZHSxutbgEXEuZ7GdnO/bV013riSl7/A3wMTO0o+5gZ5TxhqJkV1KXeYyBqU0C69C+9csOyN
rR/LyaQJWZiWH4W4CD6YOsrvjfDGPfsSzpjWweJLvET+I+0VJCWDMpo0Z7OT8dZavZmdujY1fPEt
UoOVQysB7NkbUiww9scTJsEK5IyT+ehIuf6Gi+sAHX0+QggaFYmYGGORqf2FRl3MXhLjHtb4jfMU
+/9yTVpiFwkMv4i0gRxb+dVsVgDZWYMTiEaMJhA7sCrDZ/+nvtmNoV0Za/SDTcPPVQbevdKRDpFn
iJIA0iz8R9tcbRziLEUjNzF8lWgVKD+iF486d9R4gSqsYGDCVCCdfEF8ZvSy+0UB6fqQgIi/8/LD
aZ3vgHyqhuD3I5qEYurd0vp6O4plIUF57gcaencvdWcqabZo97TFx+/Pase7flLHmIFIZBjFwx/4
L8se6QRHmheQVCnE4EbIH9nYXLQ95zNQ9vAIdgZx2goWVJwe76zXtIbMPZfQHXM0jNWLReh/+HyQ
I5FpMB4H4nuTPLCspG2TFvUZJBNjkY/VlhKpleBjAIgTF/60Ev+qf5DVuYWywn8lOJce6vLtFaV4
WSJLaz0YCuhiyDFzOU3LLnRnJNYNTZtRm6l7WMVy0wX2TDliiuMP3boEE19A+g7lkwhlMm0m3kJR
mqgdFGok4jl7AlRDjGlwZB4nIvBsrfQ8RwynnVJ2qS5gaoyMMGfsEB9HpJe9CoLwoSyXmNCQM/HB
/LFLifyLNO+HQ/3s2cWRzKLrXAEO2S7raWZP4ZsKknoGBXOe85ilWchinwAzmBaMlDtEfTXDFriS
2kpw38nMmHQG3vIQSxCaXyCWTwZRFHIGRSOtwP1tKTK1ZMJhNygDqmUyviyMy2kbpSM6gDCZ2tN+
IWDHye4yB8vgfPh1TbpDgQO6aOu/BU0sQUnbMtatg70OcT/8E0VJPtmssaeGTTsFDsjXVFyq742m
yGzYDYlqTHETh3fHrQKP5soF/k40hWBhEW/iOW7ZhMQxdDnmKPVw7kvPHBMUhtFsSRFjN7U0oqQy
Ryb++a9HDUByWSN2glMfF9S6ZwyoUoysPdPcMyts8OxXU5GDoUpb6H2FZzoTMoQf3ea0/C5kVU0N
rz0qqibeDkdwYDB8nO+LLvFVyghlgvC7RSIw2QKEVTrUvTKWosVXOCv+Uk7OSp03NQTRwxJI6LLq
XwZSYdEVFKsyphiBuG6eCTKpft58kd/NO0cSRoHILKnAw5keUKF2JAC7BmHonOA/19OPeaMeVhNB
Lfi7KmyhnYoPQdjWSpOJx9QonF6XoHjFs70U3v0P3xm6sF21lGJAmjiXeUbp+8ts5IHBpzAA9l6O
w1F8wLLwcYZINumyvd5XEuUY2uLho/YeBD3vNfFqsW64F1ePkNeS4rmbHxfDDzuwwyqaVkbImcbA
G3rKsArRag2/69sz9k5koD2AQmlyW/jAuRbQDsqhv7Iu91KWEeW+arY5sItFvARsG0fOXyXgI4uX
0bC7ax8a2LfnFDtjeumst0T2dBB/kLxztW0u2g70m82xQLUVeXdCbJpKKROhIExeZx6kpChNBU2J
dpozMBFBN3ywfjlpKk6wtRQIDwz0Z2Rr+h88CucHDY0c3p17/2PTbYqEroMHABz7n7saG29Fff08
NRslUolrpmfyMSxo/7VxDi7+YfRpm0foo0fiJN/5LdlmwA7O9Nd4y35dFvD5P0YhFg2xemf8T7S7
9RVKWNcU1SuphFTR0nTz5lU6kWpzIsbJ4WDVIPa70NUTIbSv4xJ2Muel12ktTSSa31brStGhF9LA
oMpDs9Ppzx86A7rYz5Cxisb4iAV9jQHvVKdbcAbIZfcqv6Re1SaUjcYsa9mF7hJeX6BoHJMsx1Y8
0vh7BaweadkF5c2S5YnBrm+l9676AlLAstSZF3IkXm34esQCVAZkUYKng9I4hjpOCiRB9mX6c1Kh
Mtq+5kcMs0qLLMRgr6O8Rtbw75Zj+FN8mk7MvlmNnvOa8mBSW5kD+RWMLaKGZKF0suMyfuxjLuMV
DvFkF/1+nA/zHG2k+3p2AsbwJGi+b0rtvgkv8FTdpsNLxK7/HcxNWhJBmGi7PLyHfEluQ6kO86I3
yYGaea3T6P4y3ohpizr0a4qr2kRk2c34RRWPeFpNxZxC0LzWJshqpzPyu85RskleWG5NuKnouE3s
TZjeRYAShK2S87ipmN38IaphpOnYyTpPV4wl0CqTgRZ1+VMhIj3Z7iHfUxn0WuvyzrJkUN9c5X/0
sYHqapBFIftL01OFxL31Qy3mJQniMWf5g1cmvPA+nHo9xgqewmSvckAwaT6g6z3iGqvmaK74jODF
JpK+tUwwF2L5wHU+uXa0ho57II8EVv8XOLr8DlOQdX3HGb47WvhCEHTkB2KjriAJFT7SHrWaIKg6
f45l/jtT+vGoFqBwrg2RTFFHsTZ0KPSxfQz2Jhwtx/YtPMNGpxI20NbrF9JlS+AWAATgDFsFNpUl
Xue1Ec7Hf6uNzykdOzQ6G6O+dcED9hX2x3Lu7RvTHEehMR5/D1uCAe/tyCBrH16wkWjfm3q3u4Qb
ZEggcP5Vgt+ZJE9Zp3lg3ulXwYexXovNWR5UxBFyjkWn3AWw7czik8PNTANF16XvDwa2cC6OhxYW
NQAwW9CsGk9YEYzvp0Jt7gatlPGjL1IVC2fqwWZsjtHVj3ZzV8Axy5fs+lOPtWFFYzLDjpBMcIzt
QCUT6q5iBYoGyZ2xYCvKeGW0/8PHYiJWf3qfGyUFLIOin/D5CrkHEMLGtZj0srpB79dRYoPNLaOY
sQdjaZrQlwIby4BYnSRLjvfBUwF3cB037K+NL9z1zX6j00gFwnKBxLHC9UBdfv+b8hd3GF8oZ+q/
t3I4C9O2ui9oMAF1b44DgDY3gQz3M0tmGQQ50q9uqzZWhaTyWrZuMhYv4ghXW/+RsM1rp2hXJLfc
YUZvvolCoQvh1wk9CM/phXTbwgpnAjoO2RbyuuvTaC1lCmaTlKtFdL2al3oN/+j14/FN6QXs92cL
dvcCUxpCA272DNhxf6mw6tlXAegeKZduD5+m0MC3YCKuVYFhym1geoEGv4XeDFlLWRXYQFfwrpU7
jj41h/+uFJ/GQpgXFm9+PyVcUF3hIQFdh5ssVD+646lndZdx3AePtPoblbZQwA1UUUVk+G4mX1D1
61wShb1CaX31M4rOqh2y8fZLJlBCu40jfhYEXHf7ieElN3QhzDhfNJ8M8UZ7gNRNuR+07DZjIL+6
03ItQI7FZzd6jaSdJMM9WV5L9eysvv0YDpiRdWI5X7tEUFJunJPhKsnEzUC9+LmmpMNldm0tAagK
0wj8SZAch0rSRjIhq8m47tzz/vXVj7FGVSr79y1K0CajwshZVTDmULGXfgeXQef9QbD1YVFln6UJ
NC3JRaYmt2y+Zi6da+QzF/MrEiLH5aA7+XHSiqrZBVumwj1bPI3wbGdmq3iZbLlBXiRN/QV3xSDe
kOUwofDTnx3lWk2yhOH0kAzoUq9QUNqk6FR57lkEf2v5Vb6ITG1mUEAOA9XfybvL3KfTDAuaHA71
czdwDX0XCvN05it/cDQSwEJns8Zrv+rbB77JrgBj8vFTGdoCx1Hujdppykb+TcKGxJmQNo9NtB4Y
2sXjFbwG2BYzuhT1vTI5o0mOnMfCMt1HcAB7Lje2PZSKDa6oDlaqjDnUwoeAnotbelANiQSlXCKb
jQ7YGEZ8DrbC2OSCozJFq1j5803BKjsJ1BwBOPXxdHHq1R7Kf+ccPGt5FlghorSpEPcZy2TqV5rn
AKu/a+x+mo8FWFUaEPJgZhr5ANrgtpNTusr9OO5YDFzPF7VbzuMroLYw1XBs8e9geUdoH8okeodH
gsv7o7cj/G/XpwMhgL6HqDgC793hZw1qWMqBn1rp2o/eDqy//IDBxFFYFf9AbB3UQMqMDI+oEa1K
a1zVIK0FNztGbR3Mpp4eQ1OGNyhva62pOGuoZiX/VS7nUHeas3R9+FhN/cNCgcAygbN+5HmObo65
UEvkH0MCebYLrmGVxKMltdZ9FfbPlb7Gcmrs3oMjejozYqF7aHu1Yy5SEgKC9BSVxH7RCG7t/toO
idCWENbZvJuUT+ZGSPp5w9bGXNpR7zr2peQCwyPiS3lVhvva1H6CXmV6mRs5scvvAR6bDOPYjBQq
ZoW88VFKnN9uLGaNbNiFCWSbpoNB1HgAnTELNVHCfwBgbPQgP2A6fa4cQ8g3NjzubRhJfCnBhPem
S5yaECIJnP1uqKBJ2uh531BILpXGtK6TAodrMlMULqrXN2Ls4VI8YwhMYig8YwTfkdWT6VoTdrE0
o5c7eavhg1QePha29QLarofn9hqiWEyxP0lpzvms83+i1Y4f3HTnmMew7F1IEr6a3bwm32D4U+w0
fxAtrbmKwNrb52rtidFRSoelGkMj1V4DfQ0RZj0jMf7svzDMF8lIEyisTpWHbcJrPebY4/QervEF
S7vNUbb5KMClV4V0nxYK5IqI1wUgZmAru3NSWmBdoqLh2he6GFhHXZF+Vd0N23wpWb3FusD2mswd
H3eVKVyiTLzSBB45jETr0ifDPUrOkXO2ONvLukMusdXRLcUy1CHtyJMY5C/Xf8cfcFjzg7queGsi
DnsPGuTTBspHqs0z3q8U7scYqqhw1aNLkAPdJ/CO/jGes7n56/b425oIkeLGvgxTQQIWvjyaNqS2
XPegn0+e2uz7niBYF1AIDGGR+Wg/yFPmW9WKOsvqs0wH4EM6hoij9BD26gr/40WALCjt0mhT/wvs
rzxfLj2JSHRONUVzo3mrzsLxO0YUvkcvDWUH/OUdvY/mXsjYEFTfZhHh/hI3T8lHFqUJ+RCz/t8M
Tot1lAWjJex6sx0g8/4hMnlo6zb7zIC9buoCPiRhBMeczs6WGRwZfpUCXi53H6TlD0qgmgWrgEeE
EDOPs89QGDoXO9ISV3RVwVgS/ow32uOVp4t70WM7xIJ9jLaoZ9Pce2OB2r5kV8A+fvhw3oZAFvU5
aAIE311bNiYzexwrXP827cuS99S3hQKCmkHKzhQomyTxsPucADv41XYx/azuNjE5ZsMJbgBd2TZs
NSfC7h8O+vdQoXsvE7OO/MkCWYTS67PLT69hP3cnG2wMWy2EJQYwSbPnTXLK39DRR3VUmoPqPIch
rh7artNYptnPZoOnanPP7uNfXyC7cm6yw9P63Eo5BYSm+/7eFz9L3T8b+chr/QZLndkug6PVB8mi
3v9ThM/PjsJEjlvwgwrkxkZhMzq+092eQFA1q0eQFyEJtT86KMzUzFqa4Wpzes+66xruPU41aa2p
PTxJlrRQgHhvbUJGUBTJ54wxAZVUoNzLAcNamjRjDcXyGfe0xlaGbHPALjt0sdjUMeBz6idlej6W
cTG5k1DUoU5Y/ByCT/wkLConEnA6B0NNBf4p4SSwoZbgsFT/UgQ6s0yQpSpmfM5068B8y7e8eoUZ
S6pTAJiCd6v2jT3z/Z7w1E7Jz6OXfiALHyT19G3HzcSVN8Gk0dJzqpVsxMJV+eYtDrGtaMrSpsdn
fD/aNafnyko9AmSVvO1jKWftNduL65BrJf1vg6NXfxO9zOcUhhzDqmVy0i3qraP45cK9r0Cdfpv1
zzYxCg4v5W8zytxcHEkJP0GDVYHtaBKt/Od0bPOPee8HziU44CGhBBh5m3na53JQy75OBjYIVGsQ
6hOXKDDgBb1eD5t1iOq2uFjahCZsqPWXW81cDv4oAJZUORJpqIXEHTbdYIZYtLeXfcTUIgbShox1
aLzFliqM+qvOCIiLhUsQ3QJWob89uhssuerkQoH+BgkkLpuWhhK50gh7cIxXfIk6Xtiq6/UNkPuC
XMOMTq7UZclsnk4L7LgoSahFe/rzxEACEMfcJ8uvhQt+2pIJ7dXoTiPjgPv5KUUOKdU2Jze6+u/a
kET4QSa7vYesWOK5GA3P5isxWbdIna9TxI4QLFaM4If30vclZVvZTklZJMbAN7aMveK21/R2HnoU
pRMtr1+CKcHaABXY1NkZFxLk9MUloyoao8M01t9QWfRcN8Zti9ZXw/Thr+NtDGIUlFUtOIhCLxF4
ZGCtgLTWyQBx8GmEVidvVf4gQxnX8kLfXQQX8CEk3zGiIWYKoWuZFFWLJGTrDgAa2kSsC4MEqiNY
qpB6l4wxMcUGSqrRVk1Y0c05b7nCr2QYEZzL5sN4xU2r1Iq7lr5Ew0AAAKwluPCrrC0jsqJKwIdU
Oj+z1Y46xYU+aykS9qloEM/aLYlXJxEB9JqmAf5bEAItpD91BaESYDzYB3CKiVa+eRhf58lAvCL8
4flHV90k/6Z9lC7/0itsMEsjPvr/mSL/Bfl8qT7ZiDIHqAXr9oepZKAtLE/WbeR6bXj/ukeQvzcD
xrBBp0o0D+iYOPhN/Z3Z4X0/8i+Cw4+YPDOYCYHSIOBzo97YSuKIZ7E1Dj6MsHXMKWyoOkRM7jpJ
Ll8WEFgFJxJr2yMstlRrYuJ8fearc3sXheq7Esoy8ioZOWcdtfbn4cqSWKC6vdYRVeMLn9UPhEiP
oldAn33PYuXOzjApkUoklRfUTCr6/6hpmCCkMqXcQBiKcRq3Giy58pFfv3GnzMxSJ7Nha+RThy+P
18BSiVt9rREVgoepNQ7EqibpgCie0oAdb/T0frg8rvcMTXl+YezUF/qAmIiLU6sQ9Uo2wXzM9LZH
WoPw6bMDRxVcRhLN1bwig77rfuzoGMDiUTw45Z2LRDsFA3kKxJF1qe5OIdqqZSxe/xwkcZbCE4pj
6GdXAnz3CAggXOtUfnCuMj70uwIFFn2ZwumXM+pM2F/UEJmrUeUIpEFd1oL5Nse6incUcKvdnogC
44b0J5Uu/+jjThSZllhLqajiney0jeIkJQUZ9j+kH4xlhp286q+4mfQy50fwJhG2V/wPZUPaAUUv
KPhpV06yD9n9ViVCn9Wachwfd6EbjBxB4apzpzfOyhRmybjEFs/2RpElvdOt3handiESlLO+BR96
34uoG5nLeh3SShTdYyejwY9vzzj11z1mXcyN5NJAOvtzsHK/+SIZDVxsQA1dzdRC+RGFtfng+YoJ
QVgpuWg/mOTDDHZc581NroyaYQVuugIoUMcmNtr38D6oCGarrchz07jd8zt0EFCi4/ao55uSrSQB
KgUheCdT+bFh74H8TQyPRJqtsShXQ0cP0HF4VmnLDlVjF/vH4eG6JKGco4Y3JwoPKmJBiC3JJEht
etJSU87aQt7X2bE+aCCEcbnuRbCk78t4UdEUwGotnm2QFKrnjmZrDrE6kjWDKoXAAR3Ohi70XoON
jpAjaB+dfnNISlRTH5iQi66YFa1pQftaumPV2jmEsye3ywTLG6aT896sEk+SoRASFUeyMPvRcdcp
bxSAtSO1HGELDfwjTnkXI5o2FwEqEV5vQwj8YE1+u7qHIJfP02wgJLE1aqKE12TCPVLaKzs0CQEj
nRIrfXmK9J+yVC8OfaCg4SF1RBCV8GPrSRQBWakojlFAZJY/p7AYxwqNM3t9qIdcFK726xMfOJWw
5rofQa6V3Qgpqp8fBxqpjtUHJM4zj3FM9uAxtt3wT9HOifKDBaNdVzx7FvGIoqnWMaU3tFCU+NYG
J4ng28vhoBtmVTuWgJCCgABq+y2Pgtf6K48Ts5hA4NyDRD3Dsg2px0+GPjMyaSohNGygBHAoDBjW
IRaZ93rgJ0XAcwkOD8Izj+ssFBOaqqvp6oxvaES1RVIqIeibnx2tPz3AdYpHLqJEA2aYUTafJwIa
LPHE6Kki2K5gn+1F451P+3chdnFQK/lKwuFCz77nbNxhCw5WW0wCAFh7FQ7TVqQwoLEabPHOOO9W
whgr9PxDG8Izlc48BA7Gse1kJz87/YcgIkvh0NO4wvJroSAXkstoLv/DdAn/UdHGVy/sa1WhLk4I
94CMsELEEeqYOWjwSfjVsvE2sHWz8UqpBjK0ZJVvhU9AQdDv7CUOy8ksuh6/iXJr3AxBZxuV3/jn
oLsEyqdQcRm7EH2dLpnwBf+TBiUfzNhvbmpY7epT0rAJmkpZeJvh24w8onkVBOXfHbS4IRcjkxcj
Karz6mfRGMTfmjXntL7KWIHzkWz+6ddyOs8WU40iw83AIM89qWGeYuPU+4VJPuqdLMeWHgkRef6A
VzP1jY4114+kcTwaulMG27E3gc6e6Tqb79TBNRzn8I5FchPC3zM6SMJh0HemfwN8xklNagEOFDYm
6UDtw8izT0qRMSXQkOJ4ZkW+fa8vhEhvTJ/bW4TUTKX5rVCK4kmJck+Ec4wwnw7+S7vjKxM/5Mx6
A/PuHkDBlGda3UP5Wh8eSWthreIRhTDdn7onaG2dCY00qWOBu013cKbh52Fwopo0M6dVrnMW1/gh
HXpnsO1LdFslh2/P9ZtKoZxFTJo5Xy8glJKckv9PWTZfaNjzk10JeeDGfIkwYgThHDNjDo/aE4o0
zJ6bht06vuFsYbFM9IvEeg4lqCnapLyeclcyTNyOh6BavKygV8xAEok66t2kgu1prsottR/Bqgwg
uWWAx9kwx9d78f8XreKyavXXuAKu2bw9dfYTXBEEBR0j7eRMRbOKiKZv6PDwp8QL1alwGY8JUf2F
B+Wc92Lx4VO9QmU1+i7hs8eziqlycEYscT3e/Kewa2iZ7GqT8Im9lapWH3efEwTUWSJ2sM8KWr8r
4J8xFvnclG33gVbP0iR0Z7eBQnBFfn3AYx6/p8eCXxSibc+SUArlFjZZJGZyE4GmGQJFJYZ+ykAv
6f6uDxock544VcvzYC/+wkKxxm7PAW5YAEHz/XhSjkIq9VxdJhtiF8Z0LUpxQ1167zxPkoNlBg/m
hCy3egotXR8aoDJgbZIsPqlxN3+tYQPBPo8ytD4idxQ6ye1dWISZpq13ZuutEGhuTUKHmierbTe8
HvX1D6I/pPgMgXSi1BJBtxSPD3aLfLBfTor0tCYuMjGQ0hnWLZA30ZP/YqoYLL2VVXZJ9YAFvKFy
2fTJSWggx0laP69FUp03RFgrTHeSbDaZipUu1UNKp32jodPls4Di8l7NyfrU+cGPor3iYVBE+/hL
1qbPJsqRpJ9ysp3yuWKMFhoAP8pZ4olT5xcjluG7YijPhwPmOnQOrgZ+DtlhmPWb/O9NKQgLpiLn
8e9t9kLAMym8EeJ4DKQDrSo6ReeQ/ed6d7Ln/jascyEegNI8XEODkGMV8nAereEiTVT/aMYiGiX0
yXy6L7P+rVIP6HBnNX7E/Er60MVeW2N3IxTS3Zq9vyNVtBir8pq4PigWCtJxlwfbj2A1je/NlTLA
cMV1xVtSJh+943ykuvEJkbCVi8h0xbqOoUWG2jgWAVhk45qf+NdS0l2gZ/a22+VwCiItjW6BOD90
PqV5/6pDOwcxAWGWzmZHTZHvUDnvQEqbXbFDmhs/stojYpJhnzY5EvlsyUlOxpSnw4G9ucxMvOHl
8XqbpCftIUbNHsOF+wYokF0YATviOQU53tE6jwugpC4BHOE2x0nj92itx7IGAFdUv/qwft0f3oQt
z8qWxMyCKEnPavSvYfcI9rbYGiUcgMvdjViZ7lTskqrtPkTnB7qIQMefm3yws5IWruyq6vG0Mnpi
qtaxGVvb612zgtoa4P59DTH3oPJkJz/5fQ1oBLMmmcuZxkjntchxMOvYa88lAEkM30+QxO69T3g3
G1tm2HX1ysOL0uD8JfYQGBLx7pRU5LeAake3KyqmNLhZNDMuEvCqfqbORCI8i0+BlxPkZjGjpJbM
bJewcXpcGzHjaAUTHYfGNAvdfSPt9fjmBW/RaBM3GP75l7xoqAYYK9J3fFBWFNhOE/2vErHsCx51
GyVgK2chcHKUY6IL804qoIswZueNov9gdhYnbZNAhrgey6Sm7YRE0zh+1w45dEH5ZqXmUOm4C3fn
Dj22GAJeuC8SidNmSV6quMtkb4VrIAHNLW1wkvXAE1WEqR6K2D8Q23azF4WXpo6QC2hhBEgh1uGs
ffFSMpWDejWNKU9021bMV98ewceRpcYy62iwrjKs7I2JWT43Md+CeVx7jWVDGqYveR5/mUCzyxm1
E6tKvHu4cr0qInAleaaoKeBeOj1ut45wwmGYtHJtfAF8bfpCeWu+fkJeWPLri7ihZNBxaKFI9Mfl
0/u2+PCFRANhDS9lxwYrNUmOVZnLIR6+Kj7UYlnWaA9pDQd+FFUpNrs26kiIofGctiLrBaP+8Mdd
fh/TnRvHFaRmYh9HS/eh3l8Mv6QHlNY5J9GQFkgCNPbKJMsBMv1vIv1wiKzikXTf1SvXXvhAUxl3
v5t1KvH0YPDvWCAoxlHqA+M3To0sWbrntWp6gdi9TH5e+8b/BXNxSuiUuIbEC28un4AtyqhE/jIW
0z44+tsqPjpmIfbZd+2EPqcQsD9Zg5KboVnJA+AWIG83ukKKeSbJ9rQjyC3mO7JmO2rFq6L7ek4w
mHOVMNu+GSY87UaPJH3n4OydCXqr5lZzKAMXiH9+mUXeunDtW/xrMhxfQXDDm6+ff9RuqO1Fh10f
jHX3J2xUzuRCFAFTjpt0vx9dhqiR1xcgj0HDfmM21RMpOxT5Y55xGuSAG8FzZGHGWzWh78fSmqdB
GQIqZQP/Qth70wtNBDgO42bGgA5JKjoMkrPhWUYm3DSIwpCUxoeFVZfeoGDsC1BIB3FlajY3mE/b
hqdQBdWR5+NbE9i1m0U55Ppz5S/l6EYUvuw3uSig/5o+CCUIcdAnQ8tFhOANWftpeRaBOdev2U/f
2tC688F2vpM4X+wEHDJogRqzfBXfOh4IBPOqQ6eph4E3Iwa6S+5lHlqRkcVBSQjgVmwBM2UbvVSr
igCKGlVnsoPabQTRIESUR1qL+TFB4riRyNqOsZ0vqY5x2qhIclBwldbx1/4njXlhxcINxZ4v19v9
xigp1nB3zwqAAqOcET7akRXwXfJkqxJScHZL+CQ+T6PPf1TAnmICbrc0AtV4jAqfEi1UsFPiu9yO
W3txfhtlDWmMNM2j6m4C/UthEtLa32uokoou0kOhXnjK6VAxK4Sf2MrB5NsPvlsiFxKOxVE1Ihg5
+jFVrHsORF4Tnan2bENYv3SoMyOMkITG7mqWxQGoB+FwlN7tvcCw3CVW7WGsawBGtHqA2uzBAQIZ
PAoZbW9kj91bxVOL+ZQR+ORjp2ccr7Fpek14ghCft3YBTcIx3NqL81mzCKRaYbjbqjvOdN9ENz7v
gLLWbTYYVqU6KVeACHsr3ByNtg5aPLSuh3c/WNyQb5JT+UVMGWGF2+nAuhGIeezX5eAIGB4YEnw0
/mzk5zziers4bh/q5Q9bcjVzG7eN8Xp/P+RiAGXmYanh4VL7iMJhMGRZqzvGRigtiJqdQSid65CR
NPv+sexGfuJ6PY+sHBDVrbt5S2no7/kUvSAcahNiRBK7BQ8Ql4LG+MDiHf+dYFQDJPcRyuBdAN8o
JLyCLV7QxgHOH76bj2BlvIXiCI/+rLzdqdqHPucjZ7asuCv45mF/OxCnU1grYWX4zG/3qp6oq+nr
YxDRBoQJbnpC3dfOjHY9UkhC8faLbeqaeksxWzxHHgSFxzxgG1QK/v42tA70rPLKA2IfCHVzGwFY
IyHkcXJ31wDxDJMiyjf+xVFTv96L/0obYAy+csEfIz+qb3grg+AyY+w5iJCqXrAhUUi74/Pgt09a
5Dz/LMzonBe+UF/1AfMpUFr0XPszxURnOeBgjqPUteRCgswbrF0qLM/QuNkRHZZGfLcdiEt0xOV3
prH+SlN6iVnEKTRM6xnZRGErca9ur3WtIqFKAv9vCEtvD6hwsygTfWt48YqQ8rG8waqxNiR/seHJ
YI1fy/tb+Gfj5g+RSGftquqMO6Q36Qg9JIWiWHus1OgsW/ELyOFl7GsMzWJ2TJoSOJ+a5zBAS34R
JlDgskErZtYyjDaO61e/4pLmsrR8+RqjjYRi931gKfUJ8P9L0l3oEMEeOn3GM5Dg9pxhMCBF59uT
b/yAmq9TpDZAULuHRHmhmTxT3VQ8ulfWyRNhO6GCgquZqb+tfuLvKiTcsdAGIxBmBvKfc9HA7oHk
+GA8GqmN0zX44iCJrs7BdskVxrf8fJHfFXCgXEETn48+RGmFtkf/0ZLYrRziQb8f/bdXECDDoiuN
q/w+Hjfjy5GFqAzbySVo0J02InPtnPu8+NGQoQaESDiWXM68ehUVt5bn8tDIa2OxUqMPG35TK4qR
/CknRII9KLMEFqZb+o+MFVuriiWRzj3BMul3z/GePYEh9fPiaEGvGsRT37lW3408KdjWJewSDHTF
4x+PBQyUUdbgrgBu0/C4Air/4dG4OVbIlXmKkXvY3SihPPfB2OzoVE42lnxEJhGEuCDu8vJMALKW
t+COxCqwT9CGPrO8ev2LDT1uTpgwDVs1SZbK5dB1ync34YHW7qrFKkAD/53OnpYSy10R1wei5N79
kt0DUDJnpgUz5A/IyZaH0GOvAXcClhg+8AI3alp5elLQDzhPAJ98mJrxbDgivIM4nk0rHcl1lab9
EqkTIs4SkQJuFZDLFv/2pJCH2Vtke+Z1fZ6z/7zkU09AIrZHKuzbXRlYX5Q4UiMs//0T146HDtbK
+o1ecHxikM9WhCDgaQJyqKbu9X+KDtL5vv86cxTlovRERIBvMoKG1NMQqd13MmEnc+ASt2Y5NgJz
gW/m1GcwU+FxnkHziZfaFxhZbdZl3oBs76x1EA+EjLzGQ9CqI1BIWvhzR0k18D3NAzDiEG1+0BMP
IYvVdqk+IN0LwfyUQVlVf5LVKHwTsHSd9ODgoX/PP7quqgbTsJSbqXidulIy7VNTFJxGFa0fU4c0
g3l960cQMtvLlmV7OoX3owh+WZJwp20t7fCCuICvtgp1O4a2ikEYMlfCWxYXkKr9GpXx5DYGk9de
wrDqwNCE6v7pYxthHusClxUoS3Wqoi95hKn4boGSW85O55jSkygkgmSjZvnhGkENkOJanV0bmSTc
19PuEKeVmP35s7KVMnq+VbEzaB85jNGcGphU8nUUGUbI/t9CdPyv/vfx+ZUj2aEqyTIGTl7Cwjzv
dK9YtWzS4myhH3iTBdLmVaforFbWSeLsMCaIJDpwqgnlu6MHvu8FiZjBQavvTrXEjYAkgSQoE01e
WPbEHuSWH3t9+1zm46RTzQF1xD81Autn5Nf2xlqTaYxlchzUZa3DR6eZ54DyWmxxJX7tlSsbUPZu
gceI6WWrQPzUfaGLylld5Ej1P5/D7EnLb2Lr+aTCPHzYl7fXNugrQ70Q0hs/7VwglTRLtMPk+JbT
oXev8oRLKzEk3vnq+WnX+Xy3vM+kTvRNFd56S9Z11kv0fv6djaJ0xAEZmIjgRI9qVy0F+BSzSHuR
WSEIgw3UByUACqO89qrb8IRwfHdOnj5zs8ifU+RLF/F6p75RiDkvBlCUKXtmDzwBquoGFzbyGYJ+
p0bmsze/GUpQN6GYTzhkZqHWmSHTblxo/a36SUpxUmhI2O7FhfK19RCVpI3zCUS7K1bIq207jctg
p6I0vK/1jCYKD2sbQVk4aakc7K0vMnERCdq1ic6JHOAyXp5hOZYlDyIw5IoMdWW6A8v77CtFTmZb
7nSwwDjESS6qeHOdhDH1Cyc8XKCi3FUubqXwC7jPR3JjA3MEliK0xpDrLQ6mL2f7b2vBIJE14Ox/
mJyHemkX8dQKFGOafgOPLRDKOknH05OZcD3wuQJlXw/BWSe8LuvSVdXz6QmafRnQMkfZx9zMhykf
+LFaF9szLFQpZCLLr4XZBrYUZoFQK++6227FtXZGEe3mm4MbP9VniKn8N9dLNDW/Y7wCgogDo3pp
cxBI8skeM7t1vxRg2/ctVDEFynSfOHjpMo/2TWpT+iFbJsXtoxzICZqUqJWZQJ0MYdYrv1Rkrk/6
xqIqIP7ImOSQ9L3AN3NusYLkTbdPHQqykiPWViQiMUVed48Vfd56qkyaReDMsKubHPkSUKa/echP
PGncm2OqWM8Bzr8IXCLyx1zXmnK6ymEpaE4FEd5Bjh7JYi5XojSh+2vLxJrnnlRb4U1ED7EVRMT6
UmU1qILgTMVtc78kkj5muX16OxnDET5KJzgx7RhZc0W9ckizTrvop/mhIvabkfq6HMSwNLg+Ls8R
5jE54rIVPByK2cQfzKWzC5kixLo9T5JoC7qrX3YURTrUMfSDhmPzOk0QXoYgeyKGPAf5gCABaCLo
4+hdbhbX1zeto/2sMqy6nNEB19LkTZTs07ebxBmG1/4wJjG8kykcVLC+J+4VnAn3Ndimocx3x300
sSmHWN7Hgc67iXldWYuXraR18joNauMqgS7089UBcULXB6X3bBdwwJ7rfcSbICFf+xovYhNBc3o2
7bt7UF4UELSbiq/Nos1zSAXOVcfzht2LD65Euu9pV6fNbshfreGc+BLINaXq8PnVkNCepMGh2g3b
z0gHoeDEIliPvbFRZTds0bGWia7SaIn+8sS15lkfkQDCmhT5VbSbMuGI5pCX1av6I7PmLZ5ucttL
ySNWvP5zFvgmv4qDN6/kKxv1VPxhZr/PR1BtxSPKChnmS2BpXFsV7hfpDrTjGPylpt7Y3A/ylOFQ
21gVUhN2VtCBPB3apsGXp4c8xixCjM4PNSpA8TNJIPEzRDZThqW78H+GtKDAPm6FOo1s1y760Vmp
8YyxZHNPtf7/7m9iSLrZUq5qPN2U4oIyJjlVLs0dLYRSaxwQ+T171rpk1KYICWoh33j5tDEge8xc
N4LQ9jW5lP+A6bO4L+QYqKHZ6qob4lfjcq7rq5JeOUzhgr2azxjneaOrc+zFuPbqerjP3EoshcgA
Yu/BYYEdaJtOuWxcU24oCKdIlI0WU74iW7RJ3xzaKlWYOJ2AA3i4SF9Hy+VWyfiSs26/g6t8OZkK
4Dj7k+62EhFv7Mn6FAGB1BoBgeG3us7zgbkQftH3RYoBCMeBgDQ5xU215JdVFoTXkf3QGl8SdaMa
VIzzcNHSsHM9D2WQ82Hxp+kivnc37ghztA25RDTiFwi7hbOfPodu1gydmes63b1gJ/ets+tGlwEd
LsAqtPXjnI4kPPFZf5RiXNEkE1pjauE0x8DDCrhHe6k3UAILf+DD+NqfSw3cKD6xV0y+l3K0Glqv
hQ6gVkdCX5UJ8FidzutTF1GeuE/KBeLTkH3YnNxtz+ucIty3a8sHz4KHy3L6jDL0qtcs5nIs1Lr8
JygKR8XpZHuvUyHyhOHIf4IgpeuTqSLXxLCHXo/bBas4OikNbO0/vhp7qXuJl2OOSPiG8KeggYNv
QXEeI19rYYhZKLuUTyQNh29xcHRdquNt3PTDfvbhfaA2IDpS9sBp5WHemu5Qq8GudwEfAWajeTFh
gdz8Sxj9Uj/lJaKwpmK1pu0FjQ6qC0j7gcGkzyiZIX1dXqYtAeKxyisINmzrFEtwLI7V8b/040L1
YTwW7l0U2Yv/c42ZkmuzjJACDT784oFFhEy6R6PyBIDQVBuzqT4cJQ7gbelecpF/ZqywTF1IYDFD
dLv9U/mRsqTrYmLQZAWSXEB/hGN7dq49OM9u9C8wq6BfhhcilPjgQwWr5yaivLUKx2fKnQMQUcmD
GelXmHpYbYUMM1P9nYqhvycy4S2OjCZ7T+OE7Tq7UA39Kf3vLqHBe3cv7smA2uFlYy0N82nuII7S
1D8nhcm3MkBja+MoCgpPzap0y3leWtsiskUNazIaSCBmOh08qiLVKKq2tToYVrLU0OlTxaIA24ye
R64vWKPJIbCRvgd81fZEvaO0eEBeDCnuavMZxOOdCpPv2UBfsWTB3ztO+QASr4tUc0e+mamq8Xgm
RDmDW61D3A5cxqTfVTkkaQ715nLAuaiN4DqwUEe6dF78uZ1m8xMaIHyeYD/yRuWsUQINIOaXQjRD
aDLGXKq5t0XYWg9WrJeXcDTZrcwQAZMVEXBvQtpdMsDaemgxC2Esq83N3ZCI8A3bxSnkqV2w2pSX
1eMiPtf5LU43m/VagSOylEUj+qn0eLqQsUgSfAVRmnpcIo+HDIB5vKWsgBmWTnZWe0q+J5uc4Eyf
XutxLWUyFIYeswq2jpH7610OgnigljfKcaFIEChpngQ2EZ+h1ZpkksbHldZ2gn4WrgKN23SI8f3V
/uLBNXl9ss5Gs8V9oT8S320BamN2nBkkUUxfAwWhkrd0bY1gAXx170JlDpyzXJ6ITzXiIRs0daz5
hHFBYBkV2nfN/xA+YzJbMKun4jAfsW59Mx5xssFK7JYlO8+fmM2yXQD6wk2eNGaHQUF0JunmY1gs
1GPNHiynumjeJ4zu1T6EZgnmpgb1o6fmPwufLFjotrsHLmrQ3k+a4ALeFQYlpFOOjtRkbJMdCPVz
t4/bikCdc54+LjiceP6HCWArRNnuRyyZRwa51U92fXRmrTIPghCy/dTVwLKiv9nQ1MGYKntjw9sP
yoMLc9uVctcdM4rrSylg6n8bZXiWUq+TRXORYzY1XtYAa5b9NXmh/f7zOTjeySkme5hEOAy+klFH
EabXpV/BGh1pDP6ABjtSs+iplcJabygEp1TWZReflB+3lp7k/feNUE+uFXdCRPlXVRf4wZbfLUp0
+O+VuHRe8saKYj+xDbjDOXwwxwQN0OChDhlOlWDZ23waKnxORy/ajzWJFEZoqelXHSv/QtNoWb9d
GuooBLGNO33Db1fuzlUOahpzRVhnLgQLpiaF2weCK07pkf4pt2rTho12fS/mUW6RO3cbeu8sUeTF
k/YoMARNZ7WDWO2Khpp14ClmMbcdx3dUINGEz4x1SgjMdZDvXvNJXik6COQq75faiNZUjdyQKWEX
xYKat2c+/B7ZJfBRHODg/lx8L/GLpbLlGAY4NFqVS1ucNztvL2EC7amCj1GQCu945yPLQr0H2AJn
slwWX8a0AhrjuHhiw5S4vQaoUgoZ+PCx+d1pAr1hBejyR88vdufihMipSjb2ChM2K3tkfvOrQlcA
DARqaLa42GfcmcCXOWkKXQS0Se1rReRrhPzzH5ygyCb8AbV3JbDAjTIQDuDCICE7pJLqtf5ZEwGx
rIqz0D46dt0JKJ3ZNc3vw67gFEM81ugndMv2gjatiI1Jrbol0SZGFE2/Sbt8yXzJWgwDVe4JnxUc
iJ9MpnhJtjoy+wlAYzotKd6KU45qpeBFM4++ZiWKJI93Fjgl/Q3jADJRzBdwfxq5QsF6t1tD3Rwu
8GoTgMZuZJG1ymZWjSLWiJruhbMnyQrKCRvbqiIDKkA4P3hM5dVzrCOJRJXTDPPfZjilDuqAREVl
aOaslkZgftG1AnlbEF/d9qg2U9i19F/OGJ/+SBAzsQO691KstXvbgRJ+9mXT+6a4wK8OGPm2VYSf
glyxydsBr7A3qj6hKK79K77ANqK8mm8gRh4N7MPImQ1+8ERWRvTE8FJhfC4LRbzRFojiQOvo+flB
1Vt9BlCFyQ5z9ErWu5o9bBpyy92lXeZ5FhvQn5wUe6g4fStrSDeUh27whdx0yNEweAxtDqbsKcp0
Fc6rHhqx8XCsoxDft1UbqxVlarYNM+FmzD/kp9ldiyLsxi71XCD6Yk52MEg69HpfTyD7OM0pXydS
OHUzq7N1qs1glL/XJPquycGqnRxGGkKYSEDRr64mDSCY+2JryBG4bExOSJ5iFyAlmNklRp9jaRu0
q9buzK0VwDP3SIcTubpk9GXNUXkLSstCRn7+eu7Uh8K8XzgsSfQmjq9BpbaN2GBIbVNArX3BdQ0+
GXL98Qn7ibsS0a+67IJut0cGucV/J0737PMpX66iMykxAwG2tST9mjJuEZMG3ifHNhgnpM9FGvc+
KHF4ovKZlwyO5oHm7ErS7Q3F2kfHKR1JVS2gKw1c4523vQfDRPvMwoJGbkvjDvEnwRj17xSv0EBl
AhKKSS2RnVX30szF+11BvOfP3lZCZaRfJBTstBfTkVZdWD9LZ40kg3wz3pDNDxUES7Po38LEIOnX
EwVl6q4146avKvZ5VA3TXnewdzwRjSL22h6F5KioG46lCa8dQ0ghDr90BlVa3nFROB3x3DPiBKPa
E1VgeS9gGKJZCgg67Kz7O4rjUS6gxlBbPzWuSI5rTpdp9H/boTXztp0+TN5OfK8nCDA0v2odwfYp
mB0PXOF3uHkX/bfT9NQoT3YumxdZ4qRTBJ4wvD50yRoGFQrOc8zFz1TkCEpmAGkoW0vMkVLG63la
Zz5pXoaJA6Pv1MIZinekn+hQbGcENBYg8ZS/5CBS26pbTqKotveBdzLzFeY8FhA6IkyRiev8CydV
xLMFeKgXftXp7bqfwazqDkpWW/cRiYKtObnP4eTatnHlMxzhdWGkkkrkfrhWB+R+xWbSBpflkzUN
82LrSollLt1NrNA2rV+U4mPrsipzK0mhxumx8T4Lozl8Tg6Hl+s0jfA9XtLOZqOpyGAGyw219Xdv
L8+QNMq6iWDQS8Q24/uB/Aa24gfKmmRnAfvm9423XN5Jmgl9M+DwDopZQmyrRXPS8aYoizgd/B6/
/OTY5kaYsPO39Pc6jKKS31SeBeho4M08LtIQCK5hONBN1UMYrm8mN0fZWNVGDfNKoR2BLD9WQ0uH
erSDiZme2mMnVFuqfkN8+fe5oH7N/VgalwYdZ1sQzrHDGcFEj692+3QlaYndk8N6575BHFbtUj8w
EyRqYzw9GyI8jbMPQOae0U3t725obbviztGxsJxJ/zIqG+ApCSefPbRdK9Zi0V37PlbGY027UPb8
pcowXouOnTaJT/s6nhrSdEE0Q0tvIfsDI5yyFGZyTGTSKSmZusuY3AFXzUvReJfMSrFzLYGfpeLr
u4+ZJqifCZ9vDZbRtwvF7Ck2H96JdHy6I0OOt5g2vAWYsXFXNmQi+5EBaV/l1Eu+c0JnSd6lK/VI
z7jE62VjLYDFBid3l8Hr9p0f2+poiWCDq/dINrBKJjwRVbVj8Q85AsfrHVLG6JwmEYBDRreehh/C
FbfemPpIO+2RRoKAYkSGtxVxqTaxRzwwESHllYervIgecq5S5BvyGquXJsoAuANgkCjgXNFbHvSX
N3B8cmPqcxuQDASENbUhP2NMrKWz+k4ahyHyJ8hEraduVpgpAX0IkwiK2d4qNB49HNEDVwT8+geO
6RXufL/adM9/NfDpS8+78UAaSdebEJl3t/WG4W0B8BcJFFBwP9lDoLtRZQ+JzqR1LaJk4PMKPBYk
d023qb7B73HiqCg9XM6Tr8dH7nAdIp1gDp6K+zpp8kOfZaP4c3g+TlKzugijttxtv0nhGYAnO0zn
3JST3kN/K4vskvcYXDvvaSGWzaTkdEy8lORxvplF6kfyvpWnPSOo13z1cm0SMdEmifuRQA88WgOv
wQfuXHRUcEYAMHSXQz5+2Yk0UsxTNWUIPgqQsYMDVROopEdDxK850WaqVPaPwtNqyDHa8GI2Koho
/Rc8hVUk23U0amR496l1c8kM5X5JPfrnuo9+ZxMXjYo5eauXmB4cNnor/x1kCTFO5x0Irx4jkv4o
P/WX/5mzcDT0QvAdwBs7bZ+PFm+hdnam/PC9HL/wTSXyrE9qlba0POXEoKZjiTEjTjqawX3b18hd
oPb+hxVozizivIpzGy555WTDSCgn0TyS5Pb4qklw+ZJkHJ3z572AuX0+r5upK18YqXLBE2Lmwqz0
wBZ/HbyUAXyHShw8uxborTg+WX6ytA6baiQvDFLHLQlqTZfzqAJ2VT8xFwTUlZGwSq7FJ9FtgMm4
AHZyLSOrqVtgKsDEhptU2yK/QD5BM6ps3oiHUAVCO9zVB0UloMLKzgAUL2PLvmWrPJn3wbUPX+qp
jOUH4i/LQtz9UivgJkjTq1DZ0JIBWFl6wqdg8VkwFUmjl952gEcs7EIYImZvXs6kHTe/EwXSDsJM
pJZudc2eZOQ91KThfhuKn10HDDh3dP6Wraa6Lg1Jo3d76zQSsoybeKRxlUwwpvq59Q3juJ78eDyU
1NDUZyXrGMngt3s3O24bMhh2B4epCgJG+bTRgmpGT4J9fVWTIUYwKe8bgEA/c3M7PORnat90XSj1
97ckcj+bRo4+5HWWAd3rg3cv+fa62lnyjJq68cnzgBjpY5nkBsCqTGx3EmIpTHt6IWqyvw9Ez17X
rW3ie+HAskWF6PmOeQMLwX2ZnDMbaTYNKmI6DhKIvIAYKkf4f64+n8886+l0Afu0+ZdNHlDTottn
GE+Ysh0fhL2gmHRFAWshZ9V6hKRnoC2Sx8jZLu9me6klxGJM2Vjn/YUdorpFwHD79NXARSacsFX8
YZzSPoKRTFBGeRWj7y+Dc9QvOWVfNLEfxUegmQjUf5SKbeADy4Y9EbkfmiMF3enc61OVVCK+Qi5K
maIlwn5ak7VgEFeamk6ph1UvPL8QpppTB40H50PkbM+wjkXFC0+Y0Yw+k2M9uBdkbAbTsiab7uTV
GLlGJ/3ukkfherWHgFWQLc2vZHyl5P54zhQW6GCAMblf5FlFuB82cSq37OCJ4CUS/CTidwlv2Y9j
TlmV3/Nz6JDbaagU1RLyLPwq9cRm+46orB60oaBXbkx/jvnqbRKTUBAxPJ8h+9DrGFK06w+b197/
tIpH3IlCVsNyJuGdliHUTrOM5l0u1Kfc6ldeAOWj3/3C2NAMiXPmtwZM5+9+kVpoh1gdz8j4H4/h
z41BAfCHaF1l7Mi37FxCE7sUTGsqqxFchB8cIgBfhvAS3XjBtbWzpTt4JP5gucQRQebMbSrvAW4d
eGOTuTldm0wfD4nPDfObT8+qOWQN/lUVZjNiwATB+XK++63bYDCLV5nnhsj1tA1CMfrdGc74LUc6
VEau6ojXyIiSpHKuvnZy/WejZ9lpBS3tWRvU57AUyqgVhBNiNZIGzMMVhbXvy6OQNhdpVRadfH0N
n2hw6ogzaC1pqdBs/mPX8OjGkOTKEHiq+4B7zBgaJmkMAJIuLqYSL4EzB/4bVlxCdjvA33en28wN
ODoVgi3QstYxU1HgUowRtul4dtmgAnLYltlyewypILl/5YG3pix1+Ggzw16nUs5GbWBEgtfdWjLO
czsSarmDlCZESvef8s9uCkKpisnjMf7p8hKC0aC6JCNxWkyICxLoCeoGvDdHHEKBHst/ulwD4WE5
do7b+cCn0Hc8RsX927YR5DGbffdPw2w/hhb83cgWaikjZDkX74lwRgqWKZ4pyq0HjrLEkJQ4/1T3
vQzmYKj6S2F1Sb77IEIFRSfoeF7zONFFjKp1w0PZIsCSV0+hl3F1gsOwUYk+ayKap+YmG6awK2wO
CLrvyE9TGrSV7hMbPSXPo9nWN3pnBmIooGgmFVVqC/c3qwYF3wkymtfGZg7+0ngAHRzejowk97nN
llQkDITtiBt1JGuVfKckM5pbbu0Tpns/KMN3xQi2iQRLii544MebKA08/IbkFNh6o1fZbE4KJxYn
s7iJqBJuVsP+2BVu4zIdI8gfygmnU2J7NhIdpTY2svcizW6UwrIL4Hpxo/N2uJ4TwxSmpUGyaGmc
FbgthyCUaE4CsVO7zATEfc8BjRY/xRJM9tJuYfH0Aj74a1t36LaDr7ET1RemNJZWnk3hDHP6mZOh
N38Tnvv4ahTawTIoaHok0FZbnv5Q1u441X5EmAkPyrg+ge/mYWHOYu3MhkOvHmYDFje9z6WdQysA
40HaxrDLONf1VIUcNNMQO/oL1TYlZ9xpVzc8Tj2RLY6TesEJt4WOIeD8iGMCTM0tGIN9rkNn36T+
uXKBsFgyCZXdOuV5JIEDJBg5Ku8azJsvS3Ow8I8b7JvMu77OkvyRqo1f7aZjj4wxVhuGzZTb4q2X
ywSuJTqfUcY7RSlRdnNgzEAb1Ypsig8l5dYcYScBzbTyStWk0pHOehgI+tkrXVH0cmriQoTUz3sE
MyFBs2YrncOj4A22g4BYTcXQXBo22/6sSaNjMqa8LYWnOQqHGZPtgF2T5V/s0+fbW2FMgFuOiIxB
EP8wv2YEwGMmBGAavxtSnhPy0BKOw+w86mViAwDCmk5GLZrNKa9xiBrtRo6n2SVsXewS3EzTEipt
zlx9vnjbniTtl6BUae3IqvOnlhNHkzQDIVE5YQx0/NAgU+CMc7uoOabaitpUwqyI7Toc1rDwqTpg
Qur3N1p3q6geAdLYTTBdiuPoBy12ltGD3aXWL2UzfRry4NTTW0jYVuiDZsfA6UECWVIZBOw5g8I1
vIW6Qf96DbHeDRAiNdulUPSNEbqcEVYH5k3nfE4tEMGK0gGEt5W8caNyp4hXLqf7W18znEeunNiJ
re2ym15JJA8T63LomfKm5UCPZw6KXHqDkUvw1wB8ZoH/64yVOBnrgD7MDjuHOAPZm5dNKDTKvQhC
/DCXRCJd/5BK4cwephza2DDArQbHgjI4/xRSMrQwCcmCkEbKklGeb/uIHe2F6SGD2T/Mll8MPn9Q
kgzfu1IZe10AGmCZmwl38QBEA/qkpT6t67NVj6RH0xzIxz2N2iFZFbCsaqUcs/cuZKL3jB/jDDB3
Bc/ArO2R99BejHdIry1UoEq83gCwV/A+4AkkhxBVMUTGHuqiFnp3G4tLTUW7xnJl8q03R0dafkr+
WNdPSBA81sNwhWmMk9JN78ADo4vAw7b1B3jFaAQ9zepoozTtVDiSxjfYtQqPwMtd3SJN/V0D5RlM
einvd+VLRUO17Ge7ANwgCUhZN0rMLEBYTO0mjbz+KY4VFNwlIAueVnokmatQf02Ghfhb1DzKMR3o
v5vfWn8J9VPKa9ZD6f0GSaQesU1uDM0BaB33CGLQKC4RTZwZQeKwfm/5q6I/zDow9ix9xdQryvg+
m0VdmEmYeVqlkuv5qMNWaFFQ4wUxnLCOXzdYxiK6aoSFbr6XxeZGnQEk8h8YsK9UWLxsSIHvxzjf
Aq4BijLj9GCW2W3hDROAVcRzJE2fvUlFnD2AFmtZeoJlVL0nBI7BJ7iFxGthTUJCcBgzNLo4D6/Z
npeRxwNtKEOxwbZxzipYK0Xuek1nJdRBDOgTwoiGYbhV9ZmPpDZeEmIUEitEL99vIV/aqCWKQB37
p04K87f5LBWzBLHfW+km/u1MItT1ECJlwi82Y5A5zMZDdoeQJ3zQcjujR277nQX1YUkR89cSN3qp
fuUR+a12UhO1FY0jqdjpBri9NcoMXJa2U9yZZiSgD3bChqXWX5uZrYNQgF2TrMLMOZ4lHLSf6uCK
/bZnlTUFLM9HHRPnY32KJZAbWd1UZT6jOgH4e5pQCSrd3CXcXI5UaBo7i0MB7PYbrYbm41W9DeuV
j9AqgBJ8VdXq/d6NJ92FY9kIxjdQERTiXmpqLM7BGxIDbasc7A3JWYcFYpdE+oLrb8oMkfhnofc8
ap9c+sjD23VuqBw3hrpHjFTtYKxB3iHxcVgb+fGP21P9E6pAO7XVOomV71PTTUlOkliuF/tIJ5VP
mFFsxZH5Df8LlVXIx3ZP2SDUplwogFzxz+OdjGc3CLJrGXXZAUexXZyIzI5M+WppJJaACG70eOpF
c2V81i5PWzNQCSEo6CTfiqoIiRykKPz90czt3Zg5DWCCHyoUvXtWMyHyvjViPYbeT4bOnsEnmbHD
XJwQvv4OTGzjMitZscPiXKeDd1NuAgELz8t+FFFR+uWxbaXTKrGJ2QkKC4mzh2LnYrY36mYjTzNv
V5SubWa13YAkdhVh0XudL+EotB3pAzAmcX6HlzQvvJfYapjnL3k4MAVPzDB+mm4lNWircjAd+FYY
F4HvymYzt/akJoQGoos//l0Vj9o1NujypFMF5xHAYgqs2nAh74Se3PzexN6sQUh3CNHHpg4IrWY/
KfFi4VfkOYXa0zuj2tz2pR+ciy62UoCmSwd+HuOnB8giYmvAk4oJDU0pOBZ4/ipJQWSFgF7FB4qo
INjGjl8Hsk6Fas8ryOW43GDEiRkXWKXHaH3ADbxVMjtOndwpMEhCny4Gx11rZS1AGeIMMqd5eJPK
ke3n5LNJ3YNvE9tJm9efMN0VTMo5+5vtgKEsWT/SvGl+alUX7TYhqwkm39kiJNApxYoZvGCm3GpT
H8z0Rfwv4Vot4rwVHpXNJe+QvPI8jHk7Y/2LaxV6Yq0HZNfMF6SVskSuWmz2MwgVAhwVtde8mnvs
NnVu7Y+qfIrcONsZCyqD69e+T8MLhCGdKqlIJD1ukUpG3gILpqE5zz0vDL5wpzi32r4gBquRfrQJ
QxlA1LLsYeyF/sKdFzviVz9Rg6bkbcXLMdfYxPdvojoQjtOjCuAzlybDBgtdGw015HpFvNcdEWnR
bLQk4PUJ307rNJ7zVsnE2F5wTgu0CilOCGw3GivIy/C6iX4SDHIGpNJR9yBhLGcTSiJKIIQj6xrX
iNXoRpmxNtgQ+hSVS0N7DQMK7qaF46JHMaFx9W5NVfB7LXu2ZZhL8sxOdOn4xV9GXE+fSOYCucxW
u/WIoguzd+wtUE9aCVkdmwLwtaLVz30ar8C8ySXG8wRbqQdRKx+vEWAS/jonmFgJ1VB1uqLGYgOO
/geUJXvS4pJZ/ydeN92NNQlJMqx3KT9HwEYqZ+nmP1deGiS758LdQ5HwSio5UiIglwKmV1z2+lAu
IDFxN6HV4pMxUmUCcrPhhKbNLI8Dusz7L5/lWvVTss7mp3atE2rNsWCtMsPazhsTaoKVwxtkApDf
Ujik8OGUpOvE8GWfUJJkHzx6eeSJXj4qe+RglGOp3lJH+LMBZI8ZZyXfLhXNL+YQMiLugroA3zrk
CRgRKVGvoa9nSLekakfM5dR4egeaiduJhoXfu3pJWkMuL3/nB9n38p3UyxLGNwOAFC2RxS6obWYp
a/G9uko1FLAfh2vJwD1kgUdURREyMaefNaaoawJWSY/7I4ZyZokuXCuGwI7WkEXG0oRbn9UNn11j
xxIwO/pdef90Rl3W8eNgXgFoL2EHY7VhK3JUALARIxOb4etAXlcj14+aBTuarlPah0NXdzLfefi3
LO0Q5A5qzBMhXIaH4d/5ta6B55VWvsAg2hmIF+UKKsZyyjhAyMmuTT0DbGh+fxLyr23PfCJSag7/
/IKEewIG+aS0HcTlz+U5//VFpKHbD0ZDBYoqXNv1dEJl2aOXCRV2SiqmQKtcNzZu76TvBTPyLVfC
EUJxmLoUXBRhoZSPH/h183DEEn4Z24WFVBZAnOjloCAAqRP0OSTGEmTzwE8bOKZEkN+SCLp7lqor
bAGOk5262nfBgVHpbBDQuNdQ9Iv/Qpx4OKvcXAvTQbhKqhYfPbTlmGadDkGnfRbzfCOYUE2Fsd29
RrvkRh0QA3+AhS4qNjNOCkF/PEisHBaO1azuqmSO3z0qy3XJNIT/r26eyZe1AcHrz/qS+L2bbyhk
WGtanMkAQ4kPVAu/bNgSTa7OjiNAVPf29nHsdZ6WB+sgpEnbtIRPakgVQnalMBVmi4df5z3yDn/k
bjdgEWT0lDjvQAC2qr8hmvreOL3ASZMxvjJWeTzwQpu8NTiEtrO5K4/NOX5BH7E+nNvzXDEbT+rc
pGHQd/qlluXRZOi1owJHKhE4vkpLMTEdbAJHRDIYw4WigbXX/BozSUB/z9uatO8g5XjcrTv/x6/E
ik4d07vOnyLNm4vxl+7g7jfoC9YPcVCgz4xXxnCt106qXBw09VIPpdDNFAph/ZQ+woPD6/p7WqyA
3SuOLgD1cE01K9tpI3TXsavoyu7QQEhCfbesKiJKXR19fghESw==
`pragma protect end_protected
