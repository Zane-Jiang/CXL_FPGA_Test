// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WaYkoZUS5C8d3sRToGypXUMdL29RPPvS4yRhuwk+j/YQP8VqrbpXr5Xv8RP6v4Iz
SqTAm1crio3Ha89hsG59Zu2qbQM9G51UBlwPj43tkUF5iT8p5MOYQMMUXJbBq1AO
oehuq36Cu5XxItyix4xsvvvzMZnGxtwMggLvJ+pp8z4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31632 )
`pragma protect data_block
MAA+/fMsdJKUrEpgMMhhxQrWs9VXyqa0FRqS/JpSjBrrdkyRYhrKDCgN68aQwkbT
gU3PR+/8Mzl2i2jkpgvMv3Z6iPVRRR5ofqVKZvfRvOZJ66URMdMU7nxj97SQ5I0u
8f/HqbPBnaB/LVufMLIKX2u8wIitXJ5bp/k03Zwe/TpCCFcxYLHZDxp8scMz1LtU
gJSmoYd1lAQyEaq/pO4EhyawchJ8QuCSLmcdewexl5IqZf8b+5ReexkDHaeNzQVQ
jldXWZ02cxXelVOW20gFitnJ19ngAVvAgUDNPBT2UbIuMIzLzD3hFQjQ6/nT9hYm
eoxTBv6c/dVHQH5qfp7K/3G26G5uI4fmssEfakBk5amyjw9wiWMhVbZJOB1ciwzo
knQPOF2NPzd76645nwONCcVH63jyXs/BH8+qdxGf6lNjBkin/Oz+keSrO2sdGQGX
ujpNai/ouNiI1KB052nQoROWjSJdLKTPpYCr2TxhY/yge4F3VyDVjDr8fh4PQ3mH
/U6yUcHS6rHOa+7MICw5Kdpx/USPP1Ay1j05Fy6IPKhmvxp72akYlrTIeJ6nYsBf
MCTHesg4UpLFnD66aF3cRRAS0yQsI6VHvmUPN7+UX/OcUbZ9M2hTruTFBA1uwC4s
RT6WGkZpoilKXaqwbxXAjwhPpzN4TetrnesEA4VlPFjugHwhp/yiNn0FFoArXasw
wWUt9ikaRwqBr3z5vkeq1BqFKdeTftOOEFGQ4PcWzzcP39ZcvfG7em4kHeNFjd+k
qlCW1DTTYwmvRT3hZW+2z8gyCt/uVIPBcqU8mBd6mTMA5NkuMWmQoxC98Od67QRy
kd0KiUCQRf46vsZgjTwFhZb+APklkdvtfSpRcDAypY62mUHumvlL5aNOxeLk6YcQ
pC7jg7Pi1iHnRUPjR3PUcv+FmsC5iVUD4vekxcdWKVoXDfUTQs6wVVannq9puhKN
MYLOrw3hkCXxifM/+PTjVrhNiB0hFO2BB65USfFsAxGKagHSIOv87iZph2od5KIw
mIhank1f/UKk8pUB4x88/ZyvHaW7Df5CmxHpQslpxiJUbqm74QjsEzDjx57J8NQW
5HdanDXh3h6PlXZwC/LI7UpFjNImMtbKptPT8B/yQxVsjmRPlPdO9kIqkX/H7oI2
hoNjBQ/l/yUbjHgmlYEbpg+ZLHqKIN/LsT93w06p7r/PD95NDT1eH0ASr6qj2e46
vxXQsgW+AI0AzrktTs8NJu8FtIAtZVe5R1YufO80WhykAzPdQu5H7ugLrkatsym8
RRGyEEsHqRUjEiouGocoAYblDsylebPh2fmtHPBMq+MhpZ92F12cjN32qsq5GP5e
/Cob3BZTQM/OtuC0DyWhQYHYWCvIuLRrnPSMa883QVqgnH1ZRbm3SBBFXxRPhFXE
8eyazvxCmXFD5h/+FM6H/uEHBHAf3NjGV2odT7ASX8xerjaYDyB4HOOqJreRkmtN
feJAaYkLAuMuq07NP04j/eGARr1vfIw3kY4Njm/z/wOl7ya/bkU7sNTKHK7xrPYm
qbZeD/cqjDanFOc64m8H8j6BinlN5XQTtTCNxMKcXsDoPI+owMnN7wCW17hh/dOG
2uVdHpM/KS4YRsZj5yltXAGPPk4jCRErBijRXD2bnAR0MWT8MUw5/rJBUH3oYbn6
2m7jEyOEC8xtutQTfctWvSBvcPK/FDnq1I4BXeayHIMuMoACSl/zSymEsT1Frem4
NI0WQvftK3Hr3qlVsyDcfZQXq16mW2/cAK/jFd8mSyVvQNuaM/3+5peYyIwbaLZ0
p4y6V3YJxOMgYt/JZM9VgHicVcRyydF7AjnGiL4h13ZG/gCajLF+wuOIpbE3XWd7
5MyJxRigBeopGosAVC+cPhPPc/pBrnd7kKtMnkaJXMp5vqpOJCZsZy94j8YcteJI
4mOGxoyw/ZR1G6v+tMi8Ob8yboqX270xx2h6NJ/qdQUfRKG8+KGAxdaFdCJ9ufHi
rzDOC4FUnPseuyd/7amTzj/+UObCOq5/hogbHVovcGBLzW0bwvRTMlOraBYuZatb
vJo0QT5mNff5/PT5bVKdA7JtiqvjP4LVca3nbCvZQcUza+vaqX4Fu+sZzva3k53Q
p4RtGtARxo5hNxfv/U4QmUlKcIV5FTPNOiJW0OdEajzj91X2Ttzx0afFRB2L6imL
t4iGWQv/DwpWBsEfBuaaE5dAMFLEOmq54rXyv/gEYRKLCSPAq1hOVa2Ij9u3ZyBv
ZO3QZJ0/zPaDUBl1d8sZVyV7jfhNpEIM7XSu/Y4iQvzX4LtxaTh4yWqKl8EDd//Y
83NklAZonpZvWVJlIralIRXzquPFrNF2ycbBnk6ymgm2DoFD38jN7a2QQlsomn6h
t7Wo5FcL1bVjDJKdt9wrpJPR0qYrI80W2QhR98FUwkfr65niKg2+ZCeDr3/FiQZe
hgmYimlwxEajzFB4FYY/kGWg+emyw7lu1SgNn2Jl+pkyHWXgglgTVwIrrxJCH3vM
ACg3my7ca1tmYxUP/wkzj2kTSUCD8ZY0YEbDTXVnOrepl2Wk2+5LYB8OdUutpAvq
R7n6BucPvbL0qzw6iINObEHi7FZQGDv1UEGrXk4VNRcY+0JYPt0D1ZKzqKPvO4ey
34lj3chdkwA7UY2jO1recWE0Rx9/eC/vxXLjHHhLpRkZBX4T2MiTm8YrVubrKpR8
wO4K9hbAsiGYzpwkWd/fdMVdPy+GBYMz1pL4oS8zA/8v5gpvMKUbV/OvC3AZWMZw
D64U/URoeEZ7sIu0jar5wZ86CPsffCLGfYDNo4TrbQeW2gAjjt6Tc7FGKT8wGQtS
FNLshUa6tdgZlm4rE+WzQruJW8FHLBpsCUGUvhl3DAPbKr6xfKUccrZjgc9uzapk
Q1+t5AsJGeMOl9f9Gmft5qxQtcW1JOjG5gJ6LAm1Afg3ZDEshuJ4TfLdIIwBHC0Y
+8l+K2CNBBuGJWCxtrKvmoYBVE4MZwFeJhtaaNKDlmsG8ttOJewsVqGdWzbDmSdv
m/a9DYUjPlLVBCAkn4MCqb5Ws3i/JUnRDBlrzQ0j93io1YnQOJ8EyYQIDlQFlYD+
CxtyEQY/vzjtVLg+MvQ8dqusetJuNFE756Hp+SoEiRGhvfP8PJKs7J2Djb0Z1yjh
6+y3hSslsFdzT/sxZVMFWzN5SaIfjboD16jiEdc8/xMTVxiuZS37k1XbCIS5obtW
3iaI0CEhyIalv/Y3ayoZ5UEMVK6PZH1R/g3sHOm0PkpAiYq7lrye2+9TdQiwJ4c+
V60ySlZQzYX3A0PwtwcuJiO99RGNcWN1y/MIS6ooGcY9vll8wkCX8mSoahX7yzPN
ENhBQkGvDF2xnpNdqI9OW/gBRKFzVyRker+GVPk1gXiWDnaKoFD7i1iftiUa8awp
1G+W1uOfbGohZ9UN3xQ8aAQeacXDsZYaOLi0zz1LsOImR3LMIDoQiQ4XCYHhD5iU
kTlR0FmnIzt1V5roWtjtdCpSuez0hLWScgPmLST14vRAwkhjllAoWFA+8Wq0BQ3K
F1Whjlmw9yCJImEl+nvchL087OtSrGrgfB580lASuDvANHUOP+ZK1eYZFFWE5RYx
DFV6ZYxvw6gtzKwAG5kUgk6x1SbuQ9H4St6dCpn7Obzo4qcZCa7hsW7+6grSVUPG
Ur05CU+vK3VPjB7WxS+J3B5q0xNcmyArZPugtKp3bqjNMdBXSn2hARwMuzN/aqgw
Z63yvzCboiXcEw10sFSB7OXSejPyNuLsa4EZhTmjQfg6ILQ5IpwOso674o6BUtM8
B2xw8w4PQI58YmdJyNT01miR6pw1347p9OZ5XhbNNW3Lk5GaB2n6fJRGr5f86InZ
E+6VGUOhzN0YjAgdXaQ/0+HRbQ9NCb563Z1GUUtQjVVGUTnn1F/88UNLC9Uos0YW
PR1XKQVgxjq8NagXoodQuzqGKL2RtoLnUMQusyRAt94q26VrAWAXZB6P9ldn3JT/
vGirtfYRDLk3i2vZ7KIujJCcjQk9htzR68NiJ4ObHYULiacS1GwS9D4iRTMRYcIN
kn/JAi3q+2462uViH+ifgjprVvaY1g+J9eCOc1Wcr4FAxh/BxkStWUF4iNkvRHq3
oVI0A75J/V66ZynEsCooUBBGQBnSd8d4ncl16rXrp9vOxxRIQCB0UASO2lT51Vgd
2bTbRSdtWcutjh1SosoA5XWh7Ss7u4yI+FtS/3AhcguU9ws3F6E7uczwtPHj4Ql/
jRYhoBIUkrm77Q0VoSU59qvqzaJ2qN8qQGiKbk6B7R0kuc9stbIqNixM1gz1C3Ro
B30T6x2TqYFpuTZ7wNuoHIGWWWifVSGe/IAaHlodFfJyI8J4oT8wIM0ZAjJeaOXH
LgUOCnqHd8zK9kz+7NKsBYItjMNne9PYZUFPR9h7NSshhz22QRi8iUsdBBXnnFrd
B08S32nOp4vN9wi3BA+bpk/ilVMpzQag9upYxWy7uPEDr2ArrOcFnbc2c9fWGxvq
tQBJgYd3FyKxwO80Wuxbf2OzeffLIle83XORlpCNX5QG51M9kVEBmTy6ujNFmnw6
CbR+U/+fjNeaxRmPmryEYuU4zmpp5vTWRXzGJ48LmNvJRQk8Bj6pUrtR4nuQpuW7
SiDnJp/HxAno2QhHKAjWW5cEa2wVPJtBfMZgVOsT1+45eCYW88o1DamdsMLMBpNA
yjeX/CmMuU07FHnbVNeqrnZWIW0FlormcTg+WKZ/M91fjsKlKqg8UOOXX7D160Wj
SgMxSbx/W+Ohybor63nz4IHSkCbEmoJmss0GN+yJQuN6wyMGc/11jj3q/qTl088S
GDuY5apZyKtDKfbrR4n/x40EljD08kiKnICyio7HlYMj9DsVylUE/xEZ0pbTv9WY
aWBBlBcKAl+fXMIj0e1SU0tROf5GpjkE3y2LXA094IN5kZCPKpFtpZIv8h/DSDVi
QpmaKnCn1gayn9m2nYUiCY8gmDmjWlWtEK91ofKNl76/fU9pui0toQcKo9xiJ3cD
Cv/2oWe3UCF78622XcaTH2V0RMd3uc1Ug2bdaRZJ9FbzBnqiw5wp2c9I2lrkXau8
3CV2N7mtlf09as59Dl2OX3c/+EGTOmrEzLH8C1getNC6gTYixw4H3wTU1AHmihrj
DKe3v+8mqsclcFtuEz8ojNjt2Wu1YU/2ulh9A+xXNKAiXc/G2dIh33m1TN04cTq2
IkJUr5/B1ysa4Qju4hKwfcZTAuo1+RszPPNeIMcoVp2FqhWn1E3lXg4PGaIINwdr
qjj6rkMdycBGYW7Nf9vAb8g0j47kyLee29VtoB9oY5I7IB/VEd6CSjg2wA8goaH+
v2kEAQI+Ip5g7j5TEyGoI7ZtFpVRMYDySc7kXo6QQtOfWbZ8LIWQoBj+o/BFBcSc
urSKTnWV0X9ikcYnJYZbdGGnmK8kBaPS/6eFIMYPLECKmJABk/B/gTMVxQa8BPNp
houbKTJ0SUCL7Xb2/3jSlItHcr3ISx+JchkVHdqte/wBK3o55MH7mkMhZrqiJlzV
BLCPeNEkwxAfDoH6joDxgo57wMyLICoaVSWZo59hltznO+/EHF+kopxB/5M2e4tk
neiR5vBpx3NlKZY7Vr8vhYNPAtThCkbaAyhkXlcjOuCsUOIn9hmHunn5avv7UWac
qLund0dN1WK/V6X0J60lFdVUSFsIhFqqJns58GZ6BaRQkmCkuSF0Z4hvK7yBs+RR
LQjXI4wacn+C0RPDR6eOYGOQqt/lfuO9J+vg6AR1ZjMvzWYgAuPc5VSQF+czyn0/
Z0Zfx5eV2UQ+jW2/snZrICNwKYn/3YBqtNQtcmcyaTHFhEgmcHzs4sBj1c8lMXJO
s5bfIFc01gWY+8zR2O0zjzxBNg74mbsBQ1Rv8WZaZVSm9N3P3nedNVMqoj896dYX
E5NqDVvteMm5HriEPnQDOx73b/c1VihI2unpQ08Bm52LYoEHWnNMhXj62jyd0sBZ
RMqkKnSfSm5QLaK6MWn3sUHUatdj24LlqN5AhKS8xkT3He3enaI+CxlfQQ9ozRNn
AFH//vZJpyp5modsxrKupPrV0ydPvuzDj8m6xBUsK/HJc0fMiZnNXwa99vGCPQCq
8rXKIJi70EFrMw8MhsTGB1vGblcLLRx8enxHG1V7Kzq4g65ln+k63k1bomO0tGvo
8MkI4KY1t+wkvWivnPf4URCC+dOeOBGG8ksiLnH7rAAaW5R4pv4s2UmkPZqq3TpS
Ae5t/Zigie2wxwVtXgJOjcYpDkvzfur9x/zI4A/6j6jvEwFvCQkgKYUpCYBMqHIy
CUtz7ZP1sT2mFbhm97hPoFjP+BNAVTIj0lHeGbAFPl8rIByvpPPrBiPhaZep1I3t
+OTHXuofJ0eOtTeoJ4mKfU5NddoWMVYkuu9Bf5aPC0MnxYFJvN2jp35tC7Pt9K0B
MuLOnoGVeltBT0N76OGhh8MGJxrI5ingSZ22oDHFzkzK1l7THs0CFn4xQcCgEija
ZEhD9Uinvs6mxs7TlRZ9AoMEDeGjr+FPWX6wO/b+WmCBThqz4ygNhz0Lt8mJLL1F
/Fi0rrOsrvtm34olR788CRZIHPw5Suoq1GRrhFGSoBbBbfxR1Q/l5sisXKO1MVcE
5YrlrBEHI6O4PMPOwnkSBGDF4+La3LVxpHN3w8EGqZyrR7pKnr9uFOwfJ6kCX/Hr
LhZbAhQhTJESFg2S6djcgaMDKCMuqhcJ8qr+wZO259yIXSmn/AI6Sk/u1vMBtzKo
aAyXOcygIlWBLdmnwOCIs3GmQGr7W92Bj8bnskItuBRNf+c0srVhNLo/dansANwT
ZQHaZSv/BDmviL+2IZZx3PUSIYAboCSjRunUwzkSj6bYq39PMaagQbid1a1gLam7
jtruNrgnn4Uu9iKrnYyLopTqDrZtfTcRxt2Ahb62XRjym4S/AO9wHJlhK9XKfuV7
785kF+73kyHhOAOG5q+r7AnClqvW/ts7PGGuPnTIKFSmdfXHfnjPabc2vyKlttoD
6uqWbMk4T8GCKfNxyW8sY5xw13wAtFDtjhWfdKaDOB4Hi9Wlbl+3vseE6SUKvPOY
jy2xZepAYm5qkSLOGNniRwlc5qmr5g12QXJx+GgYS0bK3l/AwDeeXScx9vVWsiFP
AcoaOmCu+kMDpXZ7lQ4qL3ZdtuA61zU1zxJirbYY75BD9cO0swUO5/W9JG0aXbf7
1dFHZjCa+P73MMaANv8HekxdN3dTWt0lrqR2iP820NMYyGjBd+qXp4SOXN4gK3vV
QPlsEFKOE1SiiLRPtjx27i2ZhCBjjIeeNQVnc6bDiNBCGg+W/HhKl8w/IRJyXhkY
J8BFZ0uWSuf6xMmf9gp0in4DHkYIq6AbrPgq4/w+NLVZp85kjy63knUXxsuyBcMP
bQPqMkGPfF4ZR+RSK8W+z35byRBZrad4q6r1FOyBCR0IA1iftdLIVeMnuo8hlr14
a+oinPvyJbY0iPPeD436O/qIhx3T6KJc3+ozUPeA3ZYn6MJR1U36+DtSNTTo/Pwl
ZesNIBOww2gFxu1CCPsqR/Je/U6l0kfQDycWvp7UaOu7prWiVPe+MebQvfHLp2d7
HuWxgRvpeLVSukwp1ucHK96c8dyAF+UkkoLFJSkJaNUHHWdpBZC5yoS9Oh+pbE3j
CwuGmSAaF6AtsRE3ON8dZWTwXLaoATIMUWfLZKWMu/IbJtEmGMPf5rXPRvsSjQXL
+dASbv71pb1YcWmrIPtxsNHUWyvsRpLBCnnuWa1aqtzG7xUnfGQ3sBom8SJObwkh
p3DQSYVQuuB094hCuVoxUeavCb83rYEHcAQ+3IgHd6ouxpZPfkuVbNuoMDmO98B7
pfqazW3FuR5GUB1nUSKSYFbZ3cNE6zSqs7jmpJQO8pi3bCONQ7AHxGH93wpbf02J
uZxoHLyppwDQFn3XbFQcCPoVPmWovfQnc2twss9ntbLQdnjIGPyhVQIR5UzRyAcv
Wpi/AoqmzQdNBwtPnlIo7N9gzZjSltkbX3gnveycvy2+33g0d+dBuT2QKo3rq6lJ
s5t89YLrB2yfFO5zl9ACog6QWEncfuuG7at0U3Dl2dOK9AfMdpW4hKYOe/mi6I7o
Hs6kJmUhmfdRBBGc4h+OxyNFcJe2H5tzjpKVcv/XkVmtfNuzn9nvLpxgRUIUxPEr
8HAOwyhwXur0e0gQhJuGfb6LGWuxQFJYitYFTEpnXuDW3lbz1TRL4uFbn7HoCjA7
fSpvJD8QCGbbzQWcY742nCu/lElQd/9vjKVUK1i9UG1Y//1ylkct93PPAChrvof1
HEBr2/ZIKd+nXbMaOlZxUpbcJkR3FNq7icIx1f1bQbYuZTyVvPqCUzdn4qylIQut
WQ9ELCNiLdSytOA88YHaZavkcw0xbYcRVAi2vk7X3plaFmtQPaEroTJqPJMR0GPw
cJeGb2zoKjf3OnpDTWOVHEY6XTI1MImYlCjkJ5kx1xr16wPm2gdavvt2ac5KpTVE
ecxqpMHbAKKzGNxY8YHdDEOgwo44Uf5QtjGwDwY/8NH4bVray3g0xV9oSxW3gIa3
H/WW+qOVQa5y6Agnww++5wK6GKi1o0TropanHqcQnvoQz8SsLwjhPNVreXIZvxta
dh1JmklRQHfFSvwFat8ab7h2hh7raOAE6NmStzoYbjF20SsS/DIgSTUqaWd1Y1kf
2S7bSYw6M+pI8VGBHDjcPgqA06m2heGfOkx2ob05uGLqOOaOcaInxrIleTRYWpqA
/QeiCCaSN+1ck8Cqw1O5qOyLQW35YCdALdlY0IM1JdnZZbDRNNoW5JT1Ot0+n+nT
PWbNW8aQ5Z0WIoJkUMRo21bkg/MX51oD2sYU/g5kAeYwRjISOSNL7arC70LEuA4P
9M654GBopJqfM/HcDuRnWXQ9VIaC7WymkI1PVia/0EEgRg2mo5IZ4x5YDVyBHMwi
RZopcGuUnLyB9GTFLUWImf33lyhAHkGl2GfhScuWYYLzFf0THowsoLyC/j8kVjA7
g2rz4rbAhXfAS5i1l0wDLTaanYvx0cCmSPr8Z6W5uqycqBFZutdW4TZcXOpo47ss
79UGpP04hIvmAmBg5PLw8StlMfop6iu0Jezp9SkXkXBCYX6qJiWqfeloz6FsWR8j
O6LY+19dIfdqJvzvF8ZrOYOtUBkgtLsnvBg1PlaM+hLahyOujypOBlVe0Wf0DVn5
LJ/wz3v7HIymleQfXle+XMh1VDWYMU89UgBfdehLH99lnLX40c6S7OhPiNYaU9zo
Ugj3dZq7QjRtHkyMnFaLx4mRbwwepveLpK/0vEwqxV049qS1T0igHCJMaHqcOUpZ
mQqP1M3mWNQWFkeNVCaw8Xa0AJHrv2A4/f4+NGYGShRMayrcT0RyJ5f0Qigc7BHw
E3y88zurAEnXplKVTqR9OT0Xb1TdFwjcS92oOG0qsnKgH5g3YCiR+Vatc5CI4eFS
XcWTZsvoqwofMJK/lYEN+T3rKbmGVDpsL08L8+IfzLFUDQ98z7Up2oGmZ1C0XU/z
wxfZOzaDzSwN7gvx6vcxLxRzJsxBChe7a9FswmzC0nhujh50Cxzz3Bdz4yZa3sN2
e2LMDQy/2miDm2EiAuaGQ4Xi4otpd/AJoTOr1ATjkpkMCl3wGeBj3Z1f0SpgJ+y1
+d8gYT/LIUkR8bpLXQgvJEYHgipeuDZ1ZzKtIsrCmILhJDjKU95/JO1R1IW8S2BM
vWmTrNt0iJFnQRQsr5IwgzAHR32K97U85gYdtmVPxapxGtfBoF8B23e14Ktpo8NS
PDO6nVoyc5xPv2Kr2vZFqyGqJbsC4BdaX9WVYFfIkehncyAJKwkh6VDWk4XMcYVa
4dCmgZQBipPumVF2DHLxEF2Yd5vN015opvWE2CqCNavsDHmbCEyEUrZ+/WgfgJLO
lx24ZIlkxXGEUMzoecQ7HAYsVdkiehGohUS57bLZAg0JZGtNR7QLUk+4ZaK3aTaE
17Vow8Uo7zcPFNXLhhBSfFgDv3a4oIeExjyZsB7elVY1G345G59tmOE2D1ryn+lW
K6/QwU/6B5YbnNFWxOPx4xZevy214csfXNJERyRfFIC0G4EIeJz+8lLKME0xERDw
l5Y4L6+F1GST2TMbYKVsViEu1MnIEGbZrMOk4cNphD2as+lujA53hqQtrtEAq5UU
HppKcjUybajspumYtqdq2remLdokdCEQwyQ2ircQx93T4gY/jmHOsiNgR3YtSIhg
EV60sQSPDDbZ1eaKos8KINZvfWk9GwDqUoSrrmzarn2efAKSGKZMj2UHsLrpVeHM
SEFrquJ6g0qQZw9eePO7kK1PPR8sePcJDobDg5uDY/SHr4f+1raF5Xq1FIjJWaaB
h34rpWDGIj4GEc++kD0E2Hy/PHfzFV1bZV05zjxB5nLeTJmFPeC/ZtIXZaMkk3yT
MK/bxlmVkS8v2H9dVKD+k9UtCofBKCd4MQ0bavXvnsvwFui/xzNYgKNombG1kOLO
srNCjmFisBj7/iyojlJw0IBA8gHps65pfJk9v7lHwMBeIsEWRUgMtRqN0FJZ2nFx
aBRQHEPhpNlj2+vpzRFSwz8eP4O+ByMpZye1mjzfELX/Ax0vm1/gpWkN5aRiSPYP
fXkJpALylWD/s+G7CCEZ9lHj1YqPdymzoBQYgVTXybSocrkQvSdq4nbWsLvl5PUU
6pIdgxt1xVr1ePaeNmqTKjJInSAsn6eEJRDyzydDGFdno6TdjmvxhSqGm6p21KS8
KboY729mu8dliQQiOK1wgiaIM/6dAL1wbxnreTGMWt8PZ/rYG9+d5txJh46GQT2k
O1GAU0JhtB+QcG6d9bDCYvCEz7jOCZ9d5xEA6sZsABQY5YEbajWy8dZb4SswJV3F
vhCPLBpzjq6anteb0VAHeVK9DBtFtvynXR9RoMtkVFCfaxI24slbeWz6ZLlpNJtC
IkOqeKhuaSiZT/BZQJ7L6hPoXMzW54TgJ0m70TJ0P0odPk8xukDQkbmccAPb8iEA
XwmFMQDavi4muYc1vJyKTYwyW6Maqj4skVJvtShnds4Pqr0vVnpeALEdLDisVGPo
vargjEqUQ/fSDPcYMJeOsPbcN0/IuqI3jdYK9PyGqWrojTCnExLOXQJKzDTqs7ut
9nZyiHCcW2yxbP2D0yQvV+7lt1kvqA5OqvLCUIRZwe8BEiVcqlP6RLVRIy0cKzpt
/OafDV/8+liJg8y2PTkIpZQQBerej8faSg3reL2RMgKg2e45RUT929R7AH3igtrp
6OcmAGY3ybS1YV20d2v+p/fqsNlqHfUqFOqYrWEufdbKJRKLcNzBlaBFvmVrXkga
Z0l7DWcUoMRFJUxritn6VC6jm478rWIBa5r3MQBmosNy7I7HAhh9fbrL+DVtrCSN
O3+bl3fF+MBWWuUNhhJLXj91qs028KGh+87kY74rY6eRINhXjst8+6UpE3/UNzNY
MCTAXffmz4Rye2nDvSwvETfr2zTQrYzaoVHVRXcowW4hz4VV5/0cavVo1I+wSOJH
b5OIog1KXuAWI+MqaVBLniCHrNXz4f8zhTdokuLw1gWIOfFfmCB2JuPUBegt55Ga
M/PLQW8AOzLPV0j/OatVpWPW7jDg4Pxl2hK/LCtod8Cdj0EfrrL22JGGk7iYHf9W
2dzbZuJEnbDcM6P1eJq3xb6Pl/WW80Xwkp9qMhdEoTJMMwszp+3BFGhKhK6ij++V
RhfvNhI5V5YrhXb1GsTgq5WMOTwm/lwYCXXlnMcgfYx4+JsiTA9IRu4Lx+DwcyDh
Q+CnnXIbO7MCK5MrZojr7QxPf2UDkov7O1R8Or0TQyn8VlGJq6qFjy97eiT+7NSb
6cJQOsTqcnYyolk8XWZhaLXWVFhyv05/AZXOvu4346ruJOIc6KeGu9fMx7ZnzQuu
IOEwrJ3IXbZricxdTodXfUgxEKR5oAM1GCyVtHw5ASOPQ55iCeIBgBA4bseAD3Xt
MQjcE7j2KOuM0ZuvKqf/V6GNTxEGUGPGOPKJS84sKJwLRI2NI/nSQyTVVLmN6npn
dFtXz2HHFCF9J8aKvxpF0XJ08xUaFXQ9h5oktvOoUGfZJmsS4W2/Io60vh0RxGPQ
jlfbhcHe3NeHZcvUdkOH6tDkdkMVZ3CMGagS+8KuBIWsEvJcnrNv4kfJwG6wfeB7
VvwZ57Ox/H24CX7n4rsDoW3pOPydhAReNKC1RQS+zEqJFcyZHZqHXMKm584XGiSb
GIIgtRoeJ2YZ86v8r1Ncw1VYmw44ujaO68/f+PiwiJqm12o/I6Y3noWHMwMb2xLV
Xo20jXklpat0mYzoy5tyRqI3LvaHGBm3dbwNwM1fVOKVNpiI+PliIlgj57X4pVd5
hqoLaUDB4CP71awym2cgSM/w0j5ke5JjdikspbdjRa6KjTj5dqjNJmhzibrcretv
m2XW7yk40wZaxNgeKqNp/9miLCVa7D+KPnMssbpim2VjoAvFxCVv5IDw6OcHBdZW
MGkFsfHxgpje2EDaLPncmTFbI/q0U3UCSsDgRdqjOrgtEConjX1LoO6VCjpHZb/S
xam4cMyaVAVXxik0kQHBc6x2IgcIVZqGHWTD6+wHeYRQ8igbTdH2bT3B52NBSvLB
1Jedh23F74xpZ/+Oh/EX+Wg45OPkuQ0q7sMkRKLS2ql6T8VgGdwA/AhaVUdrgeZQ
monVtuEnp91oavEXrwPfTRrAx2zDCOok7QHao2zRpdu9sBlwP4syC0T1rNoiqRcO
z2Td3x4XaJFHLG8xv76f14qLa/0ZG4oh/0nKWkHRL+pvW9+Xj5hWmbwjMIDSrspz
CsCglpFlM5x+vyASM0DzmPpPACC64u4iBb0JkHoFvhhOGsQdRbaNnAx5IME81g6z
C+6EU41yZVgl7H51sUNxwwrqTo+S5OjkWlGcuaB5bkOBI+133+Y5g0RUuefCp7uF
h7phFF3Vn3oBA4vWBXsLNraLznSAbDU2cDHNGzU+a3dZxz9O3DYCSydV/wqF6DUd
CgyIOWqAVv9HEdpa8Z4JpiKDZKiHeNdMWIu783/yITseEUCTLwT2noozlQcvKomZ
NRsKgib8xrFwH1oCWqjBC6G0QxPzQU+tOilLQIATIcGSCK+Ehj13cugDrs1oqrlP
8ssHwHtfZOjmVtVRZk6MVHsv3M/pgBPzZ9rsAXqtqNmBk8L4qIxempuG0Md3usQG
NqseTvYb/7mWhLUBnMtHZJOwP7tO+lpsJG7qADY10jBo9252W5rfknTDoGST5hlp
MeRXvRPiiK9LymBkJnKWhx1XNDKc5BURQUfiKK4VwAhPk1UpWAg6aj+pDK4BYVyU
SuS5QCjttm1cITRfDYb1s0Ka+4MyyOpIaR2zBfGm5pseDFWwUYLCfekQ+hdCw28L
+yy22LWi2rdR7vnDsqNJxJBy5QfFhhFCHwN1eTczI8no01ctYdPzC5KHdu5xRxCW
JsgPipoU+U6hrMDrboKv4J9wZigE4IHwFAwd9kjWGPNjKNRIABjU0E7x3EM1MWBb
Sk2ps74lGnxbFvJ87w7/fSEBrF8Ne7xknleMMJyQOUQJj7eACbQWBPNcPLiJxH8V
Mc9hyK88dkHowrKRf+yY5OyPrcP+93EQ7If4QD+yi1/sbC7DoRHVNV5RTFlktx9p
2rEsbeGnUIYBmQC/fA8kuuLgImbdhkmtV9J6ZYv94Q0sV3uEIuduZXUD1Z7SEg7G
Xph/bQ3pRsZGSPVMPQzlVqJ0zKjHwwpLZF5oOXCu6S1j6Z16CmDcUezV9Lk6M6DP
AHLFfTcQIQgQdfPBXvCeXMC7BqS5E6fSQ9dfWkuoT+dfCGPmWpsRATgkdaDvpPxJ
f6VjXb67M5c1ZwEJ2Xg6cCGlcyokRKNTduLtb7Sxqz3bAHvnH1HQKiBVrAk9ftho
hohzCuEII2Dr2okO7Xpk757jCs24T+/fd0vrESO7RFykRw3S3tcD5RBgrEb1KmO2
4gVWaLFms+Qt2tOog3aFL4WEEJMr/au63s2VlLdf5WNMu7P/Pc+un29Etd1q/uHm
4XFyWoV7AXdPmr025a5O6m9TdNgjD13Ul1375o9EYkYcKSL6RVISgbHfnhFZj9PZ
/c46Qq1aUfe8Y360kwisVEBqG22Bjs4I19b8s+eEj2KFcnlYdeHAogq0zKhEdIM/
KE7YGef9YKVo98xA2FvhOez6nVWubi+9/313mDDRAQwJhNtfQtrdDm+gwA5lt3KS
WuGJvA1gFO/3crhNyNdhKfwttMiAi8sgZYUHHeaXkU8jilvs+spn7dCt1xwTBfly
mR/14ZLlXYjJ4lgYMn370ZNOuj4vZc0n6FbKqEt+EpDi7hXyXaYHtJPd8iR4eINx
Ir4m3pdSBlv/k51lMS302V187lPds1Qclg5IdmwyDYUhPxPbShik7yIjWYPbPqQr
OCvR6gspCvOfy72lQ5LOlF7n8UPpNOnGMZ5RXhTWU7u25tp/XtCYjT1phojo+fTT
IGOmS3f6ycfdDkY8tsKAt0WiWhjbCxIXFs666Jr5Ri4xwdnQQbqC9wCFgnewB2PY
LbjT45pxVbVvj61wZMVexcniU04c5bljx6izqQ5pUKacRQRjn2ZSpWHnwxKJKe6L
s+SHEbPM8LYCLbKW4QSHgw73080qeJU3nahANUEBvZOlPAZlh7s4jx4K5FFXE0E5
UI90ih7UaBRHp1sncAbfQ/V7BMrTWTkB0tV/Kvx6pJMD69JZxl/nJnxpvu0ixijX
kngN2m6Nh7To0XLTWGAlOdrzrFnZ6AjxB7R7ilNuSzPM7EK1Be3B7OWHv/mDQEfm
p3Zm15drSqke+d9Iogz4PbnWOtJNZ+PvTnNRK3cYfPxz4wnSPYpA9WoHdCR3hM1w
nEJ367Nu8nxrtA2ZW9gpcxRauM6vWCT3heVfwB6UL5+bsAUfBt6Gswj5GdEXnW6H
A+/Gdu6zx/g/MMllEriV1S/5DvgSUcPpXDmQlvvxuk3kk/XtS38EN9IBQ9Z4RJGm
ghgIWiawdCIP5y+7BrovtJz+hNgrJasE0YEhoGe5nI7GM3YEsf7d23yaZ79cLkct
7X48gTHPiE1zvzaQiOzI0rvVfXh/hMAOshO0zbJH2Mt+F3EYe37IFT2azQvH7sPJ
h8x9aXnEoUsV+8BRtciGVGTKd16H1RMWIMgOHoEHNZxQAAkB3egyeENe4It0qEHE
8WcCvxb6lanBSpIC6EspLdRpwDkB1XL79hJDEotcKK0U5OIiUQZ+HWYOr2LQB3eL
vrDjejhQJb2fBd0qhVGypiZb8eja/nQcYXTRONgWFzVmYO82ueYsoYhAp9v8t7Kt
/jz1mkte2SsEiekubCFLX3PuxIN9PRbBZ2ObKfxbxc/l2Jfu9R6qiyEYrBGmXk28
ltKmznf+lti50PhDK1yKHFiGaJ1BTFDMhRhB9OHgvHM96kBkgr8JwAjYgOUjRoNB
aZ52vxYhrQ7R4yce56fCCQaAPFtLKROUwecGlpQurGhZm1eHkgHI1sxiskZWi2tF
TihRtxYXT6kutnyynygZcbzdGDF52wocyZxXY+Ng7K7faEQuzK1XU2b64vU4jUvw
+ETdK52qMntKsldW3OycbqYJI+P8Ez2e/8oKn9sZ+NZpVIXR4q8ifmyIbsu5uptk
dvmXDokhgOslHfCTG1xFHEZseiR/zok3qlBREEw8oda5Og8Z+zcyt+TSQc7qzrRJ
3Ek86HUTvrxzDggmZfiMbEnCYMMrWJn9EShXnryPtfDcIWYNJSfSlh4u1jeous3V
BRGyK1kvV3SZ+gDOG+u+kuc58j9cSzhun/732JnzvM2MBmWqdwbkcapQnGvgGjYc
AghXG9LAhKSrF4/XBBVK84WfK8+vRQd+zvyqKBeg63i1IogtuHB3hu4uTCqlA9hX
hMpOz/xiRGjolReNxERfTLudLy1rv7XOtvYqcnAT5S6AR18pqPD+2pF7rovm4CfX
uzUDgkK/AEuIbEA4fD95xQqEiXFoVZFNDbk+ROkytWLtdbHzx39JucBxHq1/0K0N
1olAwegmAmFRnK1NynxoRZCqduY+zQtypk4imn4QHqG4SVd9JRZdaQFNr1ua3OJ1
nAr6BKeXoWfSOi797wiviQJtyBnDJVckEmDiWorZJ0FBwoyLEPrmgY2zHDk72bcl
pPREUjK1mD0t85kmeYJBuvMhCsKb6WMBVmMeVdjJuOvjC8g4yghLmp4PhxiQbi2h
7M/ds4JidZ/avKU8G9+9TRfxM0nq5oSc2eWprlwMND8di4GtshPpC9zxBnRnLmyi
qmV2SSYGg76QqA1oUrSjWSBzMs6TJ56pru/E+1MgPdRi6uy49f/b1VnpNdvN0NLy
aLK9HuXmhoqLeFjwBM/UlQ3dMgqA5qCzRJRBmm9QR2/g4yxzSsGa6+jNiNALF1Dc
EK5XE9r0ZGjYUVYf8giNT8oeq80eE0rSut2Gh+DK0B07s1hTiwaHsW2si4+uFldR
j/zSPTg7HmCKaLrur7LN6V0JdM3S4rzvDXZSbZQ8AL4MMOE85CqSQZRgBFeRVEZ2
wHhXdDEV9Fo8KQFl3q8LRUNtRPccQDu4s9dl0JHVb4tNpp8lHHUBewtxY4cLGf9o
ZaL3Ht3URUmJ96c1EI0eh5Njcmc2aaZwGS8k4a19A0AGkciuwaQW0HQ+OHQ6UtAE
K24S4Mm6NbYbDhSUhvfjKyPks6u1ji0dgqdxbmRhC6by433TOD2wcNIYb8ZgyLyy
WzPQO9LaQ13BXZT/a2JbigciG2alCueAd4T11sAK+/WMFKjitxRkYp3AxWac6G8Y
N/0pr+kFdYj1FjuMuqHGllzVheejPPZep5SvyYHxwrzVfuAx8GD3Y7r7ZvSv4eno
TY4EkWJuX8BMJFd92mZ3z1SnsIReCU4QeVpaEl5n3MxUO/qcx6cUBLFQUfDz6Pgw
hIkASLBh2nHN9ISdIS6TDbsde2pEA2MAA67iEY+vYzUQf2JAD0+4Eq+L3w36lllm
edb6+AxD0epUHxjbSx45JT5JW6ojLEB/vlukNV9CjyCbC8i1VqE5FpyjXUPkYaNS
+hjtx60HOzdZqGdeYBajtMkHPWG0xwZ4Ymo3UyAsz0NO9w0qTb8EmHFY7PCZX4WP
IhHwMlV8FjnfAD9y5G9nURmmQ7ZW3K2ohQhZU6Ze64wZsU7BZjfTpb6kxJETevTw
jIZQJIM8c6OXuTOQeDXPhiwuHPqQOzHgTjpLVBgrNz9ChIDotJmZLeIzkZGfAMyX
tJ/NDVmvu3y4ZikDNvfyqnj76RZyqsD1begNPjVRZptHa0BSVXRKA+MKzYh2aP3/
ZdDsU9iDhLhZws6Nq3afzIgBNIHadT0giwpAhuPUTg+tN8hGKXR4PNXJO6Na/1IR
L3snL+80n/sSiB6a6wH0baXv2OUNz+KIQxpUZA8JGx7WXrP+n6RQBSyW5LO7K5Ez
kcodR9OGh9wBl8B2H3BEU8vH4yk3xDZ94x23P4bdwyrylwGMRvlwtMz+lGTS8k5q
M9iNnd+rDgwHhmvx5XVtPMVQ+mx/IkX4A6Guwhzwq0QGj14UKUXxGb9TnPhKjA5e
jvc6Wc++u92JWZNmA7nVaQuK46OhDIO0PJRQUt6JwG/RFDEIZ2UbkWi69RDnygS/
FxeEqR8yPRdE0qFmcbnGLlx/iRmP9ErSmEOmHfrgfAU1X3NtnNp2u8eQ06Y3ezWG
vDGVkt8Rn8s9c7r0Htpv51oOo6KXALUianp8cnl7dB3Ot1gsFVv3qTKlYEH4taSg
VATOB2v0wWd+/6ZEbpNSZwEeSgWVfWiAlkhLyIZ0gm11qMfrr5oeBElTD8gaYf0j
nVtMsjOeS6YIao8NY1MumCidIN5WS7rdRgH2QPO805Gso5kZY8pJI93rb/QLk7nT
RMldEY/En8ywmQRv+wl4IUGSRjwkhc1dNUxJiCjgrB4upc39AVVkIjxd9vXdSfIU
NKFAsRWqgB78/y0L5yeC6N/6uhwQ9FbYVP5AnOe+NtpXrYtiv+MvLerHs8a2LVBl
IFyjDuLKCWsDqsoVUk2VS4A37Yvl4iSSndMxWpNKjhm4fzryQ+xYPaEwTWTkPNdH
tO9Na/wECzHub1uhYPqWO8BKk/AruVEMLZppLAG5WEqvadc0SY/1ckppuN+lQ/3C
VXig0FqF9OcbXhCkgcuBRPjUFNpb0hhC4yHJdBDu/nn40jW9kfIrcaGW2mWSjQlA
lStE/7g7ZWUsYtm9iv+IVRBh7pT7CRZ/4qCf65H4C5Q0zycnscofb9UvTwDBx+wW
psi66V97i6aQ+0Wrx6rKBbhjGwOM7HRdpchoT8EZ2cpjnuz1SpIvG5iHLP3sUFZh
FrjelVKsDnJ2SFqB333683r17L6vOEUrQxPG5DjEj3QSnjPrUwvL3hBuFws0NHK1
CqNrShZlfdoMb0SgH3O2sF1ZiXFFr99Xntb+qVwHxleWXEyS0DgXJSrJB4jt+iiJ
77Q4NbQBgNZwprFHGRo6grddfd9DzA3NAZqTBbR8pa1KywLd4rAvOkfaHdgHXrEZ
nEpF3C8QjoauL3wceOdkjgU4QGiluNPUShob1YDPQC4BKErleZR865j2VdjB0nTI
aM12Cdmn5PQpGzt3Zh+96ZvjDrOd7L4sNwnwFqeFZjiSi+pSuitSwRud+7bAMbFc
e/W0k04t42KlOGaIZeep4LdptnytSML/ypgYWFaDRhIqy7rmzFcb7+fKRkSzdctw
QFh8kKXkNed7CRBRyVMw5B7VNM1DdqVdDalXVTXM68w6OKn9/2t3IHiEpZRJKIuc
vhVfaAnoBsppHh4LA0Gr5FgGzvTrWFHnoti2yxi7YiHAxYAiD4bpI1b+4Oy2Wm1k
PkqE7DsmDZxrOm7In58P8P/9B0hXmOx3cs9yoKfvfVUlpXs4+AXpXlUF636C625T
EZK9vZ4WDUqmjMXu2g3Gid0qDunuFy8FHFgK2UKBQE+MIrDbP+UnYMt7y8liIBWJ
/iphYUpiKwO+F9TRXZ0bONokZ3otPVl2Gd23SXOn3tc/22oC7eUZkfyInHz3H2S1
bysPVfKdukthFQoWJLKf7D8KwhJ5mdf+ABsg1KUO3FqNqE3yW6O+dK+iyjFsuHXy
N/n0ds6CHs94ahYarJsHTSvSvb4KBvXn3q+SgJxFoFJzroAlIxTyimZieOhl/Vpr
nbwmWTTGhwCDdCb+qUDyLbop3ia3skywQd/8XQ014Zq5tOkWHlsVcoRqJDay8Lam
Rv/yWvsjPKcZqOytCYODySOCwkvog/pq4Wb8QQKyaxWT5Yb5/lVqu9dletLSgMfj
TxsQq8/UQxbx3ocYAP5ugKpE64uEVOx5N+NEKLCg5Tb1IwNNXFyZdwS85XeRDRPo
+hFDTJ0T3H0RVBt3VQYoynVnNkgnkGSOO4aZIAuPUo4Phqwr/SnodFkjhVNM1NIg
AMyqGusdOgHjUmfvSND+il2rf+AdiR19vD5Og2s45S9q66fSJWPvgkQtNCmYt0sP
kogHmlZ3Z/Ko+McSyqeozui7T3GlgTSn0RsYq5M+jzsjgORONUzOyV9sKXq6kNjF
65+XcNg65Qzela2V/Y72yxZgXIlkUViVNjQaOg76vnTG1md339tbj2JYB2EUXwyT
7MSHR/YPVHhzjiBUUMeDGOz7bS5oPupcfMjmSPyJ4r5cbW0X9bX3eeUjtvdvYoZ6
DU0cTwTZ7SbhdIJ+0BZIFx0jelweJvSjDMrBH2mGFwjFa0nhcmwUuGFsnewjCX4J
GbQlWdpcBvr/5nlrnoQMHxLTkEbOFQ9/JFh6c3kMWYuW//5kN3WoD4WYo7VZZy3A
JyDmpYwxFazStU/Cgchyracl9M8m8I+rcji5YK9di1VJv0YUTjRneRUWCliYj+TD
M0i1NXCv2xjOI9f4/7MTEbKtahD2uQuEt2MBfgXSacApfLnG4tFUK70y+Ef9j3yC
DfJQ9qop0FVPJfge79D0JSwj9Cl0YBxo/cDnuwcDpbENMK8b5mD+NcOcNCS5AYCF
nxyL041E0Dz3OptM8qPLqtCkI3+p07eAevh/coJ6DQH+tR4soT1tcFnAWa7Qh47y
VrEAFMtS6Iw5+s+vTrJrYW9C+DcBZedCLYnra1ZW5WLdfSKfUG65yzQSY+g9Dbww
Y3VuXYblWKlt1ADcL2w8Q43lqTulwwxrqVxohlfGTSPqqoFoAgqq8hmToMiLG0EF
1Xlje9HFtoUCofgSWwCgP2nk29riZy+irPMrDQ6s4yU/kyOAmxK8j1m4KDHhmbkC
eONSZ5x6r5DfWVmFJvoGpB40u2AIVOlE9VtysYcPMtv8nks8vwKXoffyRQV2tgAP
o+lScaJqIzbLEDGvSHmvFukF8nQ27K1FAPVA8eEFbI0r2Yjzx04j6o2Hp8h/U5v2
Ltg1Gvs+E0XzFQ5hkOHl5i2RpLFXQGF9/BmHfroccgPXU2B+E8q9rWdv2+MAXKs+
kA/Km+19lzyjlMVlTEloIevJjZ7F20TexqAue8Fy6gDWUByvx0/IBZizONz8MNHH
050DVi2RuFphEbMmvq7A4oY8DW4EKkuS3BvXrwr8aYBCQOn/FPOaJQnCgWncKjmU
dHS8cNmxX3OOsmuY7fOpdnmr4MxRprkchamzijAJM3TufRtfslYi1eCc4RdA0sB/
ph8YdNdDG/S3q2hy2hi35FiVQJ3I8/y1o3IUnbfhd5PfH15YYDQhdEuxTCNufCoY
6YTntKqOYOOGVb+kA4aTA1Lw4IHTQmMH7wYvCr3Y2MmsRsu19TCji8v2P5ccAdbN
42etwn8BwvPxxut/QQE2iLFAysKoqI9zfQ2QoUKupYVY6Cjvt29PtRbKH6b30MKx
mulWY1hpE1Mvb6xFnop+txd8YfqusVzQ8/FBcfhSibnAWGnWA5nRE6NY6nb3DFnC
vOBhozzLrEbt/C/7gOPx7vn/TrUIdHGq0vqw59Hq3xt89m3wTEjRy+mTFerPiga4
eL8SnyDpPrvbViv3oNUVnL8vbTWSLTMNWsZwqnibb2EkGSeRa5CaQcMIjeKfaPCp
A8VwhZ7haepV5II7t/yw5nNCVAtq7H0lIinEL9eiiFEf65EvNdr0oocQXQT2AcE1
A5Vm0LEuekCde0IksNIEPGWqeJX2HTFg01nBukRqs5/MBq0U7vOP1BiHiCtiiuLl
JzGuG957oVZZiAgBTvsJ9MDJGUu2Hh9OolDaZz55xzf1nzfLcqD7o0P2p1jG7uv+
bvsQM3hmKKukL3COIEY5amvuVRmKkEmWkibSi2OqU2R7eULlI1y06W19sdiaGWcO
smKrDumb2Dw3jGbLRqn5kPagCzvvwvCZuaaNc9DotYN50et0MBryNRH8AJNykVm2
QYnOAbsWJxGc9P7YBEF/hDzMu4JfcLrPoJEE7h3WpP0SP9152S4PRVsr9x9vRfGJ
5tD3CGjNFzgxys3ilLN0UDEOiW+CwZLx2BTBDimHL5Dh2pw1Hugtl/bYYJt4jAa7
juMHCdM9UQbhyGNzu2axKh+Jwuk5rVbARhYpXgaAwC8SgPDGdIeNrs0PPQYbXXkR
+BDSD26WZQNTKhOlltS1O/+YJfjks/qIWXdhGe7k95fh1FClv6ZWSP0PaRx+ffRZ
FMCCBsnzZVkAPeS4lYQWvdxK/fz/sjlP0Yc/d6uZhMXy7xvKMPI+4LR2f1pN1GhY
Kw6gTxF7e4PhowOG2hbwVd/K0k0Aytwhtq8Wo7g+5mJoXcYqB/0YHL2SQ8bxsNNV
Wh6h9x8/2gn8XLA6arCqBh60iIoaoPT33jGmYsrJpDuDJCmEq4J/5z8xxL+13hCD
kF3oUMYDcs6z9ekzRXggmmjrOedfR0GBgAwlG4yx6c0q5ZIqpnRiEdicVgvpTXFN
f0AcrMfA9Q/Td7C4w76JAw/SI3zWeWuDgO13BVamxRiYST67Olcg6UwxRNJMxCBR
EINpylQZ0uyLxq1fsZOvJ8iEBr/O90vixLCgNXpESxOB+KTtSg+5Luk1ETEHXo4h
Mbh0skXZ5jA+ipvcGbaIRG+4F9yO+qhxQHmC/e9s/T9IXxXLUgX+YK2IHP6N/p1Y
OoxggBR5hg6CFpFeqKXNRHxTcimXSbtQ1b+K1ETZk/ch5OPG+7nhPwwmv1fWAgnX
C6v6gquFYl5G24YplbhODF6SpfAwxHAqfk/DhGxkVQ8t1lRaKL7FYpCxBgwLfJTh
f/YYMi2nWQjQYFViTccdpuRekjObDo8qx5F6HYDkBVB8qy9TreyxJSkizJ+h0nxg
6+wxVOngYGRBO0wSjE15GLL5pUqtqS/gMdwPYMar/DF6mdoZsIEQneBSjlUF3pcE
sDD0zjYoMYRQThR/h7jTQSKlq9QUGR8wT1rURDq/j7QBzFNzig9KIZPTNJreMJ6e
26O/nYKGkdGTtgz4RDYPFfai/BbwRMo3K4ryPcLqX3y5NOXYb7oQYTlBUxXMYzch
trzeFAIzY/kDUJdb5smktWnFAAxcxSWmIropnwkDQI7TKY/TM/ZWQzmX9xFK6Ow+
dM1hRVpdzLzNS0aPqdCQCTRmFQy/tIKcDN+wwCPPKwdUzrhE0whEhZ4r+wygz9ms
VvRymM+RPd/QsNoIqLlZJ3utHpgCMy+pgzAtEKp9qdAVs+D0XhOJY5lT3aLixSxj
Y4rjJpjolMR3ICrIbUTj7w+yaQGbF6IN9h7WY8Ixs2rWJ4+bl5oxcOC9hGuy/Vwa
bgtAETERbvBlZ7zjKadgKYbZ7V6U2Z0O+Ln/lkMHpZzY+EYAzCcypck2JtwD4YLc
dRP1de/Y4st/1gDdvqClYyPXUTbGkFfWNuo3vmouv5Tt2mk4+4qBIkZUIIybNDKh
mGTQZPHrbEheTN4fJFVVKyKY8/BcDWa+MNOyd3bq6x8A/+FDSKp/e/iHU4MkfyqB
QR7fZIAakRkyHC9kX03yFf3DjtiPNUR8/e+jfZahRgj1yFGaC8loUg3VX4eADqsS
BltvpLVCbnbk9++kUwydWSwjKCId3D4nj4SFMJmrRt++J1BcCIk6tWsvriCdLgGq
a4Zgah/vvgDUEOem+Q5oOJ2WKeLZ4MrWTVL8y+4M4BGu18i9igeYW5THaCwgpmYa
U6Pv+wXB6JVER4VW5IFN5r7P8PnnIeTIycEsvT7znbK/u6EFHQdAJcftehqNXF6X
DunHIryZs+uok+aPrlalC0BzFfp+et4eABZjbHck+tdHy6yQ+Doy2C93Xnj4svgH
606wVlU4xGF6z5gc80tbELxwTn/fsFHjOKN681ZUudmphYLwD9tAlWWpGp08Efa/
nYtr2J3afkMzyxqAs1R5lrso9bHlugYkHmhBx4xvbIn53dj+Iy818KJtzQ10jKdZ
HPwFITeqMhYKh06oAohnclRVIKy9DtOhFVTotgOGF1HnxmQzgMRs/G6iW4yLp2U9
Ik9a537vtOC8l81JjQU7BYP7WmwLkOnWOPSsinN44nKHBUDPGfJAGUYa0ILNAiX5
eCzVV20RMpDZROleXrujegUiqSEwPXRgqvzI1TRQtgCOiqEXXnf2PsIf9orfR/7f
+ZL9FU0/WE3Ih6MPzfLr/J+fwAhLg3EaZseQ37pAFcThJ7NXXzViCWaXdMZEWJUB
vfGQUIkvKcNNJlTteROXvoHvTSrHeIpnWmlYHniYuyRxVRUA6HPY0adbd8NrSRCD
I2mpo5x93ZnUgEhOYfM6GnJGhlslNDmuWfah43dbqkNqIk/0x1sMDAyGY9Yw1ET2
bVXw45JXCaVLb6IqxSNSjcBzeoI0s8Ek/fMuMkDVmFIzHeLSateZzxjjxTSZXOcz
1cTwIdpLQY0N3lJx6f98B/jmdVg65unTlh3nb4Kaji0SeHhg5W+z2fQOWIsyDiYv
pGGRMo7QkHm4g/QIUf/Tn6jrw9IguHi150AYHBVpzNBHP4mMpTEHcEuZ+hpLiIX2
lc9Mpv4Sp39W96UsdgoLQzh0a6/3dlYKaLFu6q/9qd+R6dULifJyOKokY+LAnVvG
0W9mMjZJYtkceyLGjRvpyCoz4w3L97VxNgYJfwfd80pfRhMnXKoWLxWm8XtuJJ5n
r0ozxZQyjFUiVAHKXsTvFrrNJenRCpdDCseGLtqu5tAC++GepvAGkImPQ93Sf4qe
jHpHj+17DDldt+Ryxv9hOfX/RZx6w0Iap7eBuQWWO+uMDO1Eqd3JrSSudzPjNnvx
ysNTR42NuRARmjwpX47FNurjuM56Z0/9kIkmHlOgez9N4MQ1kWWRz26biYo8KTPd
Hzri9rgfvjTijNG09RpomHT8rII3A7gjfgFoEgOgbuxo+K9ON5B8qkVn8XaZ8hYB
sFvTNvP9VbjRx9tMx8MuIhFMkslrTG8/d2bZfSTOEQfEfzYF5+SjVSjMTcT8KBsI
UZWrRojuepWVtPCJoAU+ftvkICFlJtkpjEVEh8fxHpnRu7MIyC/7DTFgoSWKGIxK
LFq8VEXOkU06JddWCa3akSruLk/gTsLiTN1s3hgNsqwxBW1zy1fxRVABaZLbK84u
tYx/1vYQzsvSIF8utjOIPpA3Sj7/Xdyj7swPiyX6KMvVYO4oWRJYfMYgeJ+JQW3x
JL9CznVIWpha2urzW0mBPLXZXLJyuBkfy7JvdFWtmkAaVv5hGXpamSiwYQkcqcyQ
YBV9wyvp9gYJC64alkPJGtw/xMXWK3L0IeiN5zWJuu4dW0wDVTTkbG2LX1urHp/n
C0mRVtkM2Yk1OLU6BitCAFwZBeXoUokKEpwHu8QxC3yHoPLUPoRLDCk5A/eaDHv+
LciX9OHuQzHvW5WoscaGaIN/8ffllt5tckTRxPJEdF+F/iYD7AYfsjxNBWnH1KRU
zeW4HUEThs+dkK7IVgvuskUyybmFtWqxffJ4c7YGBUqkgLzqAl5p1y3PSZHcFkjp
wKZe2x5jT11QWZqJB/1eAr6SOCmV7lvoEJFiXCeypwxIekQ0qErwDD+WmXkzQyQv
GOC7d+yjVgkoDcsSTdCvFEhF0BHnZjNjHvnXo4dEpfnHaXttu1FDPO32oG05XDD4
q5AWBORHne7RrUOf+SXyvMGIC1LCcrRNnfczpoTVvDu82bAT+ZiHWV1ibJCuGxBK
hB0zyjK17mL34M2nU1gdfgYeS90xdj/jUhdIJSPUAzs/lUhuG7hcXAOLcIgcvYv7
NUdDL7cqnT+vQx3ULqkT+7H9ZmM3Vej7Gmih5S9wbYdjh7a7v9KaPhGUrKZyH8Rp
aGDlSHzZZpYbTCJgrEVjTkOUr87QNyagkWHL5jhRRPL0/K4sfK/QCAZvd2dX7+Td
+g4oAH9emMfxa2p+XSpPWcCSMS76evClMC7Q1P8Hd1Ap6eqjbBN20obHR+4KD78K
YLlhkrKQFsiRJA/5pUtobTSQloiVbxzO7EsAaN4ZnGZrCnbT4BwHBV+Sha0dXXQ6
4aeMgM5BaSLIfF1CFRCJX+YqpYBgOXaZ7HVK/9SYGbJyJu9qGcuD40Ttv8WMLnEC
gRRppHxgyAqS/89NSR9W6Q05W+2mlmjHBuhYn7sC8Ukm+BeUwQ1FUXaS3iG1KiXy
Bo3y0y4XXBG6NUBQ1a1GDignOc4tbmmQDrMwNtDF/LYjrLf1ILk45ixp34qNQ3Ma
v61RD3vp4MnZvAs/2CT1YRFBkj0I7c7aZ7CiVDcDveCgUmEqqrZ9/1FmnMkQWd6Z
17YwpTKByk1FYQGhT1yaVzVOS5/hhEb7NcVSAkkBJD184PO+vldU0sIKrgr0N52a
Qoa9VzQI+Uf9S0FNswYZppJAtZIjusR8ZKOglZCU2X48Uxpk0UbpglBRNRD5rRwT
vvWDeeNgi/OZqF++lQSSvJct5Y3W20dXbfwOBo4UJ+tbVZXPtGgMFXqERe/OD04x
DzUs9TZ6qpZP9U+GhjjAZkjLxOvmOmrVO0h3ujZFy5vNK/tducw+TOH4PB5EZBqV
5Du1ARYFEK0mbmtNP8qZGkdIGh0mqhc0pa+7/1c6ZRofwbs/zj3jzEeWYEwVVduB
i1RvsPJByQGJux/cv+1mCZ8TQ7sHvqEmQ2JHKNTF2IdvuuVSu404kK5ZKDMsakAI
Iyw/j54isdVpMf8I1UZHpG+OnoF+a1LBfTUevsnuCTrPvmUV6QZavNVnPmSc6ixe
CScNZQC/qhcf3Vku9WvkdAW4x/boeuSbwGEGXtCQ5yX7U6xm/SjxKZl8cWqlAK38
zJtZCZthKobdaanCFNQ1uA7y4vpqXFImlpkgIzEUqAp7Eolr65zX7aQKXXPbWczw
omImNTsY+uk+ZyV7GVnk2KA96a9LIFo4Q4fIS/juTs2hIEkrxVYVpocHlYMHxY1t
FoppbZYxpXhn5lDLcmOS57wUquNZjtTPo+YxPFxeRLuqhhLR4emkwP1O0kkk3B2S
rWluHy+R41Ho60iEg+iCBmdczpPnO/c/zM1owBeak7ARli8jJ1uCIgDq8lTaSdri
AfiLPL8hTN59KVTPviY+UFz7uYqPyOVI4UbRM03hYLtgKZe8zWa+om/90y+YNkSR
JpP0M8omNHAxz61YtYJVriw6M5rZAmZxlxXzAp+RIPvu6SyxxrOWY4yQJk10PQeH
yPeevyEXC3gnstFOjqDSC2rPrfcSBkER6X8CZC7npU14CBibEbqZ9DMla+fXAu5a
njO78DSW9p2H0gTRpKoVarJtOCTQ3OlV7JvIeoYFECbifpac6vWMkbsVQYbeK9aD
sj6GK5VVfJd6XKdIJROP1Rq1ZqBEqPQ9pdlDj3KgXEM27ElvgKa6whYXLXp6ihjC
63NptsXZz3UW+ebIvsSyeSMzaAXA5VrSer2ddF4xD1IgVuE5EEyL4FmIjF0TJO6/
wgNWzRfTQeQc1/j6Zrx+hL/fqT+vnUx0EOZYtwpMcrgXoJ/Jz+ECfIdj8gZeO3E+
NEQ4I7aP37+sRtITrP5MUPisiatQn4003Yrm0OfxcdOenLA6Yxy6cfEaEwmwuzT9
lQw2vzAnGkKS0MJUIZMMP9COjc8c8CYeMiMAYdoNU4V6UxQGNzVqynHLSLzh5Nfu
IFPxjxyeE9/F3IKGOv0zuuuOB0ZYrOAonaV6zfa48bjf/GipaZZG4xYbRTO4xZXz
n4zpxdJ/o2swF85WQW47lA5gUVGEqYjLvTgxN1AkTYqaif8Xc53/QWtRCk9zH8aQ
mKnt2nT6IyZukWQ3HWfjYsxDUDRfPoxl+FSMmpowwWhWfVb9VLPQkJie55IjYiVH
ZfgfEnV9GSWRQ2Bu157sxbKeFjumO4yHr/eHO0Wbetl2BY+gecQT3NMcbNG+y49x
Wlyqg2T6rp5GQwhQm2Xrr/GC9axikaWvZfUKaX3nqcTQJZ7/r0a+pBDNhqf/Gy0X
6TK84YczFnRtghpicDzhi5PDpNDqJqZNZB43PiQduCMJ5DtIf16W7hs45aTHRCiO
K0QEqsy/ztBNt1zxXz5ues8wLcV762TwfqHbXJAj+SCBT9Ddf7KQicWED8DDa29w
ho6xo9BIom695xXUC72jYGBr2Vsvs4X9ptzAF5AbUi239bWNh8KrJvMasXyxazpK
LCharjJN8NHQm4kF3z1ZFAKnOMKQgo9iFXAON+5ca1yA2Tn2DRn8nFc6HzMYynMy
reQlgYkk23OysjlqT6tJM2s67cNqMB8A/GTGpTVdrgryuNrQaqM3U075spL6RRyK
0kWV23rf1PdMem7R4X+bsyav8hU8aUaRM9yngbSNSYrpNmaxWyxLguRj0xVPyLsa
IwCRY+q9YVeKK8IqlfgacVNUhYLMkHAKBBBXcTl4t3CmpLRTPNZwtLHVqWU2FZSr
LkjOmc1ZjEHYmDDMgsqtiUYez6uqJ4LXQr+wMFdMX6Dc6qMREX6jXsz6JOgYJM7D
5OPUp2aNXSYhjyOSMFYzA3Iig9qN2lTKJx+RFsYzYFzhyUOAGQl3nadrC209JRQQ
rOHn48ql8kTogyu8/rvQdBOjRD8cuRZrNh/+i6I1yZnnw8oo3iUbHQZjDQcFEArx
ay8k2vBkRB0ubRIlGhm7D3jcdyOJHKGgcLQ+hap+y+AgCcBy6MumIIWEaJAgWraz
W/18771PU1gnTl0aS245TG/0cHdDk1b+0SfWClSc4i40tLXJB1DRElJgdcDAZziJ
gNplv8ZXxYj6iMjvUNV8Q+4tyB1wfb+Pxuk+fVkoG7vY28aPqbKBFkB4+61I8y+I
SW6JJSxhT5TPmokA6KLf0PrytfyWUUtI04Wq+Su8wPxqPeoefAgZfjsvWFBaks/d
7bOQwn1UPUSu+npCfQeuLCJvXDRm5UzzbEmO+4QeWaMdrZ6rdQoutDPQmyIL+bUy
by28O3k6fwyx2eELOE89MGbjwW+ySAjaTbzOXQ2hUAxH42Iiy1NrzB8EK1ykLHCG
G7eEkCiVoQWJQPaUP0P1OKRbtpl/pHTKu2//uGC5/46KSd83+eXwClmUEXIebdzE
6tyMMOW4zFOY7pLp1Z4G02nsQbohVmmsRKf4vgUsiGs9TPi7m9F9KuOvXlwyiCFh
Wag/rSyMxNcrXe67Mr5FCUjj/Emu5Z7h2CSl/TZ8itH58wAfMP1CkmQZuQA6DrQW
wxsTbbGyK6n4q/qL+RbexzmSBGHZkE1rWWNdmLxRMW9sJc6WedbQ4PuTYoIlgtDl
ACoxujxBYmQR0bW69CT1Atx9iYJMyfh/MaHONmctVzXzKK5OPBkayecOGKT2qDsq
flmz2RbEaC8xyJ2Ngxn57Dnx5tHEhEwXimnzjtLarIbEiMOkXEb+HTDj9VFoRAeT
FdNpLxftJ/DEVMM1grwu10/2+u9JMn1SdbOy46xM2OEPJi5VFhY/9vD6qcvW1/Vm
e71xtY/0shUGyPE5c0Pic3CK5ZhGlUIwouauFYxFVw0PmuMl+qRg0X1VeJyaUDaI
sN+23cx+MxgiuL8XiGV2DDFuXgLNu+8xkzfGVQSiDvC6A5smxOM+DNajhKKIX+Um
xSYcm4txLr5UIAdjDa9C3ELNETJ5t19GqUd0VI/TnnKohaVyFYndBQN92khPUfxe
roQlyDRnRPhlVM+S6ovXPmdl4caUuWNBCu7d5slSC166HcancqhdUJgxb6sXIZk+
cSBYa2iDjeCS6URfCXEz+vubNDfISIEeHs0MkzIK7jymrgR/nzRQddzyiv5NM2F1
ySX5ZK5ENYUIhWGb/JIPaMoepvB8P7y531AQSteC9t23HFY3ShHrxevzLdcr2Rsh
ftA4ORWzq4yugYXfB1T0lDAxAU7GuqSDT1AuOOjrR5pJH7CRDg+qc/bV4toeVdpZ
TTrXQI70pt170FAl902VwVdBfGijFN/AJ5PmDftIHqDHWzxvQwZIytOeovv0iAUQ
DDEhayuEg389EMv4XaGupz8tFbB6LTavdZJkSISigypyw6zS7qSmT1+RhHQ8Pruz
s4rrFDDCOHRi9ok5gv7KnJFdjmUDz6GiPI8kFObcq/0UkIq848Zhm7Yp1w+1XCxd
H3Ou4gMIN8LF355wyyEJbbpzIwWQrHy8TaF20XIt2Ig+0qyEBTfP9uCxpFf+b1Pw
5acWTKUl/ea1ds8wQh2P+EFZElz4xZ7nfx3zmu3qysW3rXvJvjDy7+vbJ+45Buke
UIhCR3ucPCD+DRadttTxia7468NdATfjmAoa8HR4GuVy0cu1etAEswpSDEEKsErc
00Hjpeph8+jlUlWeY7usk0IjNbXdi7cI15+ypbu9951TbjOXY4OoIrQhtbdAKLKQ
jxXEwwj5PWSPSfGGRuLEJhmXQRdp2wN+WkhBQBdVCfenpO3q1SIqo05Nk+Hx2QKb
sOpihc6Xb7PfTNOxrLfPsrngc65k+jWfIQSbbYd6n3O/dvbfsdLQ8jN5abLTHjWu
IDuDHFC+E1aYMJhae6zWwtMEqEv/dQQwd3ZWVHqhjEHz9cVOkfB6y1VsxbKcBpBT
MIFwUJV4tpW6EEeRg3NmDdCNvnIxDZT6cv/f7qO1n5s/2y9XT6b71F6qCgJ+qNwE
KNoEnWlZHazWOxkG/g5DD36fsc/xjYZee7FnnOw0lzGXLuvMWpTvGFWaZePgWedX
sbR7x/GyZVEN8SDBeUNH3kFaYMNnemNP/7/kH07H7jACqpm7JqhKZkF31zHeaU0Z
INc5DN0Oh4kR4aasGb/aaAvOYGxjQ6lZDFLNycWYDbAKdJW+3UtyaDKdCoxc3tHd
niKMogroo1xhQFjlgjX0FCvSryLH2lGwilcLhId5vE5omDlD/w05EsKdTNciqTrP
sCzt8OZ1OJywx6vXpQk1mYGggQNNRo3/BYeCPi5U6ZWhz1V40lHVN0PnkBjzBg8K
On3HrjLyG1hlZpjnliUVwBJUxnWS+fTLnMoIi3lIBg1jEn4hEWxXCHLzU47GeNSi
iqx65Z9Q71FXwCOHdzmqdkk0+xjg2CdZgMsgF4zu0GQESPE7YURLq0+mqOMuKfEy
SUjF3QWMovZUyFlzo23ajMzJ+WGDJPr4KuEWqUARcIf7w7cjzR6KvsMz1vUfYtQU
BemCb9SjrdOZi9VZO6sfm3R8NGReD+xY+ly6ah4jU58gDIkTmeiS+NDxllpxskGw
xP9vYg/XHJErJQzfw2P0J7XE3vHQGpD/85Tb6axGiW2X8Kbcn1JxqkLZr8ueTgvN
hZi9OOGpFo9qhyvngeekdOlv3LDkNUt9DFfVo1UHaMIiV7Og/ZQ7rwYFqu69XXOc
rAOqTvM61nlMVISlKhH0S+gZCVKEIa/NA9P57gtYK+AGa8SNXbOsWJ4qbHmZSIHa
wkfoJuQI7NP5XouLPIoVPRR0ncmwJUoaoga6CZcyC3deHsyN9LztMUPRCSPAhF7b
j41hvyoM0dVFht/hB5XCbeOAMoGre/Jn+swf6BdkEQnbva+YzIzYCTwnvKx461Ug
GEjO+Ezqd5rRT2pwQITZkyYH5alNblMp7YV8jUvbGRqUJJ7jOCVxrS3/0WUKHM0T
Dq6RyCeKK7GkELHud1PtpmcigS9Bn1nPZYo0cApZDgFxN6b/b/3HhZu9EWhjqW32
KyVfTh+o0hz4TpPQBpCJNs2xQZX6DKkTtQOitkiKMzBDp9USvuzJNquvG0sggVw+
96Pj3beAE685eAGC4BmOMEbWm6wTc8ILJ57fJUFbBsJcF/h7AooJMbjLHsuMKnXM
vyzFngeGUA8FUd4X4p5fGnClgu9xb1uZ518nY65XEUt8TZZcKgxb+g8GjRrj9Sj6
SBpO/Gz32AvOQmDIieQx2PMLHgCQWBGNTA2cqp/4p3n1PoorR0nu0u9wL6LmZt0V
rU7hX+ws6th/Vdgzvc/v7lDJUtcVIx2iCR+t/dJanLB7yZLXbbXDGJpjEafh4U2c
Wr/0D0ZHimArMxusPax6visYOcE8D48WgzWxRmaIEUT46yvCjoNN/Ubuq4IytVR+
ySS2SvV3eUh+OBbkYxHH+uoTw/tDe2egGp0Ka9f/ee4NgOAUV+CS8ONSmAk7XIAZ
19zWFmpzIscZAWcRyOYvhw47fplfBQ/CD98wjNWYRFcJ7hIEEGbpAAeqOSkBuvJm
5WTFW7wgWoBb9AAPHxFc+z3GCJZHbxDOyvWgXHC1B0eT/sCOOxchFuzADcrkOx2O
SrQAiN+egkUV6gB2XvZH9ACKfo9820NDk411op2Q+ZVZdm2R++/LRe8/5ztISmrK
OMt8gzi3SX299u86+s/6dJ8AqXPhT2iM9PiSJRTjN4+gWWLASWFgvXUmFniXArcw
e8yiSUHyocJmNX4CWPrPxrkG2uOTqcMEifB960N9sxJAmG9jN2QrTT2BeEDvDVre
HFvGxjMwGD58axbVMlK0ZT8scIcFbcVxMLlrthPs2Pdmkz5CrmDPkC1PUuwzP+vf
r3zlO+WUvhyF5bin+8CQkjzfyduV4hxbu119KB1Iv9+9qXFQDbey773XiE59u2Iy
IYUvIQmsV8IzsPKyYuLb6HF6TdwuhFGwoCwxqBe/lg1dk2+doOiN/bZW1oAPff7A
lPeH/X7groGzxZdsDdwLNXNGwMF0ge0Z66qkE7MFaBR5VXQ7v1L9FFn6vUeySlRn
ZvPnw40Ggf42BnOsP2vqxylFZYIrvf1aDvRU/r1esoUDLtv/9lc0mJduY0cU8Ako
QhqK+w/FQid0KeiJb91oKJ/Y52DCUQNzwA9FCum/7660Kh38bSLdUJjJ0/cK0BrN
6KJUcQzmALYCx9w12WRksJ9w0uiu2zw7uJG1qf7Xu95aIe/39VZp4C2GGNBLyxp2
OHQaBgcpHkJcfJblkSmwhL5zmjtr4/+NDhpCVVpGyzbTbnmeAW5Zm4AMrW3+eT8Y
4k1DKl0QWzy1T3pSmPuhZjs/VIadAMgXHAX2RmPHP798j66OrcK6v1CSMIJ+AG8H
tZ1OYiw5LZpACQdDco69kN/oXzfgp7E0uXLwoD51T+0KGTZwo4qzZiCHrkDRZHdJ
tjZ1Dzcjly8nRJdc7hBBh7zM6dRpSTrK8FHAsLvnjRavGitY33Noi8wEPzBzNaNj
ntC6/RY92ccT1jYwi00aHyeimuHhM5OXw+Ucs7HaLp4URbCfmwvYhw7smBZNPNnK
BcItENlgpl+JFmsNpftxdxrmJF2jfJG0kmqf8Xn0GGIKDFULev7uTZU/O0Jw8OqQ
CqTTXxRHC6KOk46JwLTqPAFu8y+BxL4u00CLYx2sdYKTSNTYRyqVq+1wOmBI3aio
R1sHvH00NHCH7xW86ratdgBHIpiSHjbeYRkaF2JGGd/OKa5dgfFccehU91t6AEfz
fNc2pAOTGBNpRW0Bp9D84M9EymRjWo4b7rgO5RI5vnJuMtjKzDp3u4YqU4T2IvnL
VLzmSKBhAS7v0d0WIZ9k2xGN24uyl95cQ51UFaA19ugijdGDfxJIfWAtRSLOBVHR
V9t5buccxzvl9R5k5Ha9pFA6anDv5f0UNcGVzN30HBTH5n5FLKQi+TDH5UWSrdxs
QZMWDbEgTiCZvcnidylRCq4Rx4OvuJ+5zC4gaTIoYcj5vtecv7n9ZNoc5lmrBYPr
5ajDWxyZZ/ys6JdflYjRtDcLknANoezeEQZZwfFd7sIXlIbxcIo6PZR578PagD8y
jOZS8n83edMeXlb/VN7ylapfe7RvdwRYuPDD9l/8Tm0MXoCepyMzWnd3ftcrL5V+
8NAKKSVaP+pdnSb5MHqAYk6GNslp/B7+WRn2H+/W1EnkZrN4/AhOS+Ic5Fd83yG9
Crqs4bm8mIZJDqPm3q4dc+hOyaJVnvRt7iPivlDalLArtnww/t14l7YYnBkC5jFP
Acie1qI+742HEm5OP0w2MtFXuK6Q8czCGv5V/PlWPrTR5ikgLdteiU1NiI8WaQhz
eUCXvXE8taZfGOVUuF07R+HAAO8B1wvk2OW8ivT66Dr14ZlBJP42YPIYasjIXN++
LEE0zwUlPqZJLNGNHAACYjpnjfvml43F1weHYkHGfZeq6xPPo2Lva19W/JFaDsxb
g7Fm1/yosI85TLVDNX1oG1uBH029Urs97EYN56sKcoMEj5rghY2lgbM+cVTr9URn
xtuqcVg56G3E4fuiffTr1xLeWGNBh/fWf4OEfGP6soaMQ4mpNFw9GTeo+SR4b73B
BiTCpBxfdB1SOlxhxG56fBI5aHd9QeQZqfAZU/oRll8s8IpU9GrxzXkRL+2Ty4dT
AsYXdxqJG+XoiDw18myb3COZ8XVDvW5IEcxBZbe55DxobqlpgJL8hK89v6CXWFOB
V5MugyAG1YMB8SXFskgPPvoVub2H8Scg8O6hiYPX7YdqnGVhkPjNzjI2OD0r0Z8C
hKWirU0XdMqARVFENCewhTQ6WrSk6b8IKH0sRLcpdlfCi1LGfL9N2zY3j8qSsgwG
D7LDhPMkLRDYNa6RDTEiYxk+/P4Rej1U5iEw101QFlu4JTMGcJIodn7U+KPdPteX
PIBc5uGuiZBnlQTvbCrQ1eN5iUcP9jNz0xZs3bewePfhTjJ6Pg/bed4iOeellng6
zs6dD2pEkFdzUZ4Ojgo+CymbgQtswoq+r6haMpKeD5W16vrAuneihJ4UoJ7hcW8k
fV54zx7KTnFB2jW1o0OB3DUu/cRgZoNcGPvqZaqnjuC2n++uTMjTb40yshXyCSEz
WUJc79AKeZByEex05cU7rLiXUW0n7UI2CulacdZ5AnE8OHhMuuoAPrir02sILAa4
yOVqfO5EOmIjPFhC3v6cmZCkBDtfvnU9nTqeeB/brNMoK9r2HxjYns4ZU7C3EbTe
nffujR6YXg+zKVwkkZqTXiZZq94SoaH8vmvHRxCiJLOkYbnxqIyDm+T+n3NJADnL
WDO8n9ED86wuElQJq7T8eyaoyX6G+co7GE8xe3H8mVhqlZtREEUJFPpn0o/UCcMg
KffxL4hoSKZIAkxc0+zhjOttowvhmDK/BPUPbgLDm2Fxx1N79EeF3bD6GlfVJ8CR
wywdZUA8mZ1CwMaCivk9GrKkzyEjlmHOWuxMTMe6Mkg1WkHO5szFn0oNaUmxJ31U
PM1HGdB4WJyAwehzZXyQgzdldg0JWC6nMcrQ8wpabnIYKv+6O9h4YwbDtJVjKerS
CNgxxy2WDZXDyYy+ky4q7S0KnrNfomNDdYFHBvMh3eUY3jJObpauewBglM69bJAK
Y8muCbzMyhfUpqRyopsJrqiOJcTPuV7rjufv9MIBlkw/IHAySMAtD6DCg1gkKFT4
PZOsaxKFWLd3F0pfgqzom2vUMd70+XKCxQTjkBGY4DNsbyipt1vsfo9Y31hTlF6l
VczAPUuRylX6GK/g5kg1XlHbjcH3i5ASajGibiVJ689Dho5ROG6PBQmeQ+P0NcLu
CYSeeJJ0257yC5jx/PCp1WsUAvG/aXQSKNwl5+qX3RPQcTkySUsW3xTWcrEq6IDW
Wt01Wqu4CnCH/rqn7LsYpoVUnvsSkOyF0Vw5gE40ST2kogkHfgVsJhbEmvBSFae/
VJ76hsX9NzVz3fi0OYjuhdvHufpOMc/Qne8j0Cv+tehMaX0hgaEr07fUF7rRX3oZ
VLeQ5U+a12K/NDZLPvFTThbBoHWEuTYrBiuUqoi04zATcsBMDW/KpvKTMPCpwN6W
0cHmXSUdg0zXziUEG14/kvJqwnLTG3PdaZvGHqJAp4QB35JeHJJ2p2cMiyP+Yq7T
LPnutwA9OvofHglRJtmzXVX9MRk17lTRnbbjC+ffE75XM945I7NRV3E6obeIcGrx
M5KXbIeL2sCqK3xPWaS7OtBg7Gs8ba16QzvFOSjnrXjNAaTjDo+7UDPHlNbKczC9
KrAFyCs/M6o2T6+tLcof5kbjzivYBxq9jmjJz7hqgSZi9JwlxqAILGODEs1ILOOk
SzxPKT4gdvt88hBK8NtEzKfHYxJwannHQY7rbOAd2BeKKHJ0sbOQQ8Ufhx9pZkY1
pkhRdMqlgSsHSt4y9lurNbE4/UKhegr9fJJ6wTENRjwj8EvjIp7sKC2+Ce7Y/ScA
89ZXXymLuuz5AS3SDGjfp9U4Ux9/XWz/kwHVOxrD2i7wwQEOZ+NTOHQ227QbhIW/
w1gF5LvER1EEsgUZHoIThpHZ98AjqY4y+L5yIxWgOHUQ4NV1aubR8MKrcmEkNTpp
QSWuKdEH+0B2Ju015ggjSxTaSuy9sQlQqQIBw0PrKYUJqEPLsRrW8EVo4kOokLlA
I5zPJk8xzBSzP/CUiJ6/q0Z92NhsPDFBEYxbZJW7LEo1rVN3DlacRGL5kWxjJtor
M46D1fcre616QL8Sfbo9D9hxHYHFEDAaZ/QeUbjNNGNC9Fzqiw1KYE4alPePO54l
YcMYxvwPkEv/mh9z1jIxicyS1TPxjgcQ5vtOYRJa58p6TbT2v6eQJtGcb32YhgLD
K+aiSx7o/u/Uu9CbPT5nRBW/0MI7MCt9S8PGajuMESz1U/hZdKYwybeJbkREsXNJ
t0UzbwAylcGysxes5AmJVer4RTnQb6Iuv97C7UK+oM+JcEpQDl/caNMmnoDRxndJ
2hbqC+mGLJw1d33IXsWGVZgJju27nqRGnDwAjNV6XiLZM7YO0L409yR6PtZtoz/Q
wOxOGMzczZtzPjDeDJ8l1/jwKvVyH7KNGhQGWg/KbAGohWseJTOKPKdp4I1I4wiX
bpZho41KoRmSvMFLMaDsMpOXy7g/Tb3RA95M21aK9aZ1HOpkZVMqzEUg4XV/8OR2
U2mZygD6Yh5WMJ0Ux6mmmHiXQafFV7XRGmAABXSFp5L4LkNNPkBgFGJgxXpBaJcO
6z4neBiDvP1VCWWE9LWn7M827ZwRCnOFUobgc89V7/gHttTRG0ovy3CGA1CLaJiF
OAimgV8Ptm11Mjea+Xi0LXZveMF2jZyT1TvY3MT2THn6AxxY63xE6Gz2FD4f5Vdv
7DLIxPdWYj7HjGXB7j7kAD0pKzRiM2K1/lHInwMYfNZfShn7K8MT0YzOR9Ez0xAq
nAWKq06OMD19UTvpkNJMSIdOrkr55IthgcY8cgZCv5jz22MjMu2lDReFQjm8W0MU
rtY+WCj6c8uF/PauWvi4sEkRAq9dPzkcB/ID5aXoSew0r0E/tv4tF8Ye0JQv7HL8
9I0z8hQN7rasfvBd814O1JyALvrGJuvAXVPUgRX+dYwMF+LipUWonTBbMnIzg+xs
zc1WuZMo9xA/KyHQXma2UhpHVlReUfUwUESXiqNomh2mNOfwlsAofbHRMPT2MUq3
8RNOAF1pwk6kCuj87bfQcS7h8UdJvMHuMlC1eR+TmYAEMbGz5Es9ZtxmwwmSGi32
/d8W1xwQQeiowlIq6HDQhaib3e/xRN8MY9aztQ2qtW+eMPgWZLXNzyDiub1g4LKS
yojJrdlWEVPCV9Xfo5FgKoJeWjeqQToGvypF7c09PycQznir0rCcoOmeYpQocyki
jyPZ8UzlhTsAUE+BZvCo9cVIyqMqaxaYG5Ywk/YOiaK5jp5X4XakHluIg7ckpELo
3LB+ShUMjdociWxoPBiqGH80D9wrozzqtl99fyorHEb4fj6Duj1/tHKlmDKwrAX8
3yq5JWK7gc9R63jmSas4wtDuwRrRhnwsvYV1ZqGValt36Ki7I0+NfyaNPTGB9PUx
mvVMBX2it0n3HfdEZY89ok0wAjvQCUzBpuDdA6g5wnaBzdjVObEUbKN3L/5fdgI9
zBnEHUB+FX+/oO+tRQdYOW1DxMRrqDrk06bkXlKws6gu4MBI2LbQ8Yr+ZQeAQjJH
mKh9kMLYXm/3rZipDYde7hQ6y6O3YRKnzEvtVLdjkyM1U32MOSm/qKPEKgEU3Wl5
EVpqUx9KPnC1Z+U60ZnZZXdz4f72/FBKG5ghn2H+hUdnRGflaMnI/vfS0uQ8z0qe
ZGwbq5ncL50qdu3KpJDA8wnS4/+QxxTLtMowS9P6NahiDbJlqPQIVZHNN4so+tjE
PMIc8mqVLGMA9XMomO1FxZPD/rGjylZ2OL66JUemOkAc8N+zfGihq/XOGP03v3Ef
I6LD5gvP9NBuWllo6ubZ2heW75h0oWDIuJ0s4Mk8F+WqxULFFmS1/Pm7GPToSHwU
d6ynSdS0AWB4cJQojgEO0DJIkNyyg1QAjzYjDOOe5u0DHMhkvKeX463pFPu8HtG2
zJdzwH7VMs2xCNBU3LY+sXZ4EHzXld9E+4ROKlOjy/+yS8c8G80P7BQuC6SJ5aVP
+zOSQAFqnm0lQbhy8kutgTfb0vfURaHE5oRfZzZYzoU//tiEdpp409SkiWHQaJX5
wrLKRX5TfvCAPtJQ0ZTM+WIROxvQQG3hK8fJVcgtuT9qYv3U36EjJQYhBr+WmQoX
jM+PtaSkRNeTZpoSPBkSISfs24h03eq7BfJUPZ1wvS7k1yecZjVSwdMyqF8l0LMt
Ld21I6TbEWm9v9l14iZpXVGYvfbKxtzJH9wQo3HMUFU1Mc092Zgc3sSP3ELhEvuP
YOqv3fkoNxdLAoWe44KveRpjiEwdjisLZOJlQe9VAX4APdp0a6Z+ic4CPi/o5PWG
tR8lsoA3hCj6VjHK7fXpXN8S6/WVBWJh01RnT8y0svGDwRv2kQ6FH64Txgw5JmYE
O5/lJPdspQzs3YBYPt9mBO2aMLGuV0O0z6pxlpY5o1/pCbpfl8OwKWAZQ5xVqjtS
YGutqFhKMNucKMmANqGt+LV/OdEBWeX91sfn5QGeQELgd+PJjZNlHS4x7iW1nYmC
SCP0/tWnx2OhNTAhHAJzu8h3jlTFvBgZS1aLNWRgbhlNrzQnr/dRELM+ss3juEEd
33R2OVh0jjCp06SoaOBbPIPXYpLhEwjHHXX2TWBBpX3b3ih/mmHAJfcnyWUQfG4c
P/BlMW1JRRQkCSRWfkaIC1p2f2hqqQs3CTDJCyYMPNLoVrwTaz/x39rWBiHUJw7a
Is3g02EvoOoBgm/OTVokga4CJpgCpd5J6LUZ7t52PkCkqrQVDqtdXCctYPK6+6ux
R7r5c0jzdVhbG1gKw0rhrWlsWPs8TOrexcCETKNdWws1wq7mX8MSJcV+EDZaVc4W
MXXrFWdOjlS1rsZlMs4DZTJnbGaF/iTB2nC4k/+m0ySIePyAyPh0sZ/30kJ0HI8x
iUriLq3yQ8IU+Ev3O9ANcxylqV0P6CbbBz3lWsjGUDO4h6Mqy7sgfWjD1BLwhZWF
JM5RZWtwI1m1Q/gHQpu9EmxTAFcEdJQl65Ul5Pa/w/gonWmOtLiFh+Z5K1KymeWx
LyIbHgOKRaVABy45BrGhqUq6SlCZ1O4FlhqT6Dtd6gSGwrm3oYFSAq0AA0CdhAWa
A6vKVmG7MqUKw1n57ERjY4suOSiV7cLLxU4c7vHs2eYuIyAeQRzGc+y+ah3JnaD9
E8SMFePlhD75fjHK5Yrgd84wDSF7AfKMZR5FMxQHDImukQx5bwbIOYHPDmG7kiGx
vhSOOWMlRSP8eLYRI9jQ2VqxcbCKmcvzqC1aEbI+YV1MNn4SsEYOX0hUvI9NtTvV
6dawnmUt8PAEN4tO/6A+r9vlf3DpwoQFn1NeEeA5zHYpzIaRkOhn02JKg8tvotON
KVzXtDjl6yBAPoXmgWQGTQ8rUcFGRTg6brpUQt2lwHSETjmMf6etyH8PtrEhdPpK
BNhtbyPLmX+lbA6G94JnBcWgt/kt7OzpCB6VcEhbRzB58sTmjyP4CpzDuerkPdTK
EtaEjyFRn/MKT72SKPRAVjg0wwnGCg2dihz+58UInzfpUZTzf4dzPQbGiqRc8tpW
yqECbVz9c+2gPWajLA+5o8U2Ut06DZfDLHT9OROVHO5vkcjtKCLOPWgNyKCoExdN
cDB5Px+0LcVdIR6If4D6D0hbeUDABUJ0ybHdkbnSiGtfpChCRlU2M6vsP+onh0pS
BbYdfAbsKztUHqrYFyj0uWUEEZBoe4QA20/8uXyRF/5osxx9mluE09P8FWl2G2Up
c19GuC9ty2eAh5cokgQh38yUGkkRFAPTdCTj5Kd0RiW9r9i5Nj1tm9SD1YBUZsQ0
lTM3/AUxqbmZapyB/xc4aB/4ugaPxt9jqrRer6aM9Q1nfHXGCuhiuwGNTBCJGC4X
aHGxcE8hJiAILH81ViWxDP5h0/IyjM5g+u7iStI7/7ccL8kViF7eu+Y3EjwWXA4x
ddE5yw0DrH0GX4jGQapTffdmNAQR21voOlEAYXhODUk1tHJK15JeKCbB2dsfdSKP
j0BhZkt5vnw9bf2jC+lqXXWkr4N5jwKSiIsUCxO8KOr6Cv8QN3tdeq5COkgzzJB8
tlM23w8wcyeRy3XUJg2Gu1KFKWU5K6N9XRv4y0xDIekIcyo1KGaq25+eK2jcAJmh
Bek/UaPxZdt/mnHW3PbAYPKv63FSP2BPCU0WzySGvAWGxJz24NadrrG8Rf7VBCNP
O3lJpJnk+0R+Qhzh/N8wsVthzkIw+dlQSVdG9NPhVXCDPOo+pcP1yGBj3SVecsC7
MGHFHH5eHZT7yw6SMqstV/EXN1JJ+HEjcKxWBcxiIf8AKga5OHhYrDD5fMO+EOGw
UJpyX7JbQ7TDIREM6sSNQnGrQpwzPmZ6lHr0I6KSzusbp7XmMIsLZVOHdBOzTQWW
MIfx3KLbhUGnh0pNfsvzcr4EwgGluyQGvKacPBTNwBeZQ2ZeTtYdfBxxjpVJKP/4
g5D+/6zAG62jIzgD+RJSBJi9XOQucPnOcpUpMyun042Mwi39s8Gk8BtQA028gK3r
C/8tE906NUYjaERrm7rOKMwu1aEGnXrLYQg2B8UBe5xipNzF1nTI2iDLgMiJ0rkT
eer/+OsuhUj1Dr3MdQkzpAeZacocoiulqJtZblrq5OBGsZfuVAS3lY/9DFyVtBgp
U2Oo6uBMew+cXXx5UbVlGPJFQkLnqFOdGx9WelJQSfnxm041HJq2Qwomc0WxGCYH
/KJ8BVbztPAFDcOLAhIBBaaeRtCXg7oSEk01u4wuWMZ9QZX+ucPcGJb4v2yz4BHA
rDbY82P1HZrLy514NgZrU1dV6LEj4UfpA/4XSSIlfhPMciwrYceOL9qDkZU80oj6
7yn/hj4D/fDj6Nc1O60AGyV1ZZebILodmf4Kbhvmv+hVaROZLtVNoAoK0kmAHbks
azjZOOqNk8qmw9sJbvaWv7Wqjsf3XCIKh3BXKqs2W39++fubv54YhFWNeON9YdTl
ZZdYWR1Qbs16x0S3+i98dvZvTz91KDNx03dQOnbK/RjSke/XXk7CNKN1uLTyThsp
IY+Y0TnhqHZYvaEuJsBTbgVYUSkxIyN/N+E0QeyvFlCoLfpwWfnGId/t518WBAnm
yCgIbWUjVQhd0jQVwPhljje5cBPgAV9tQJw1tJ1u6dgyTjk5LkUkxWuIYI2QOFZb
rzQ48YAD/aCuLllCRpqdUyLKAxOCNYB+yAQiQe2exKqmTYR8ix4oRsvVcvLwdIXn
qRsrZ494ls/gSVkf/Q/nkRbDGXQJyRbZrGx58Yp4ZeJFJai/xksXEsdfQPQneGTD
4r6wSr03a0CHYlQ4GYSae0zEmkN4SF6NfKiBIlzvOc1etysVySFdfNEcAv7iqh9A
gYh4J3pc5j+6fPpba8u9qn4dp4tku7Ky/GMRdbWkblc+ctaafK+yduGfWAmz1mbi
4CN9SdzbjV74+qWskQH0T2WOgmWT0mQmA5GhUB/R6uLYfNcWe/7+UBA8JWMLBaVv
ic9Dv6kZZtCXRT9RFbtg6f12YhYp1oVQrB4ksABb+ma3YXAz3eR6W6PexuSg0W/q
VMavVyIKOLuK9uSmrluolduJn64KMA4TsiW5FhgVtzXzOpLWFm+1uFxhvOOl84/D
DGdo6h/upFYiNK+iSBch/jZiMhBdAEtLKGlctIXppLZoyBlOfSh2EMXoOSE9Nzte
cAan04QnPtQMxehKvW5MCItJuHwzYtrRqbxa63MRoyKnrevGIIMpSTxL9tdglPDl
ve9AIwlYOggCIRbNq/Gbdko7LoFaXF3nzbLxet433AuS7K/luhRTRDrEtW14yph2
k+1W6fRUM9wfJgi4Rb5RKOEUA0w7FN5HVhjHpR+9VjJPObkg+R4p0pt8cBEgA/ob
YyPwvcJ/KBaaZBt4wsSHFWn7x2Ng4Chjsw388RX5UbM+i/sPfckP2nPT2w96WyeL
0rcGE6vc1u/qwkMMGWUgdamfTsE83SBLL3om1vlqg+x0C6UUTGHLsTN10ORyvG72
Cz14MdMppibfGFlHUds9C1wPBNx13yTMzxbzyqG9fRy3sXGEUPbHSNhiODDbTvPp
oT9IlM2F3LGUV6/mUfPsQEi8gmSYzD4JOadewjekPnacao0ghOS4XKLzAqgCPY+g
KupGRQp+/JczCbW+wqLJgFGytxtpLlxe+b8vbLZ9DlTU/v/uO9x6KP2fvFdoDPBq
fRkpKU1zEbDAgPhqYfi3XIsAAXFD5S48C6/F9RsIosUzBvrJzQ8266E/sT6ZDQ2x
VTBS44jKuKS9wh52DKe+LVi+mN8WTuwPCwVxuN7U5OqSmNAthtFpAVXwkYM0X7Wi
gxQ+gZr7ERz0X0r9NuTVPiboI4l795oGAoZJ4gs/V+h3dDSz3I4W7uVYLv4Ql5mt
v+vvc9YcO9OA4qmIAkKRLpujWz50lNwEs73Ka7M7zQ/LZub+g2Q7KHWHImBpnFaE
ZnWDOkVgyG0dbPx/+1D0R5WHrFlaZahHG9cZn7dhDf6XyXKAswAO6QlB02dka+9w
X4Yx8DW+2Ap7nmCRcfKWZu4JOV7aLYpPy/xL2Hpcr0T9AKmdc5THCTVo/qFs078w
g7W05ynRaAPAXkodN1CJhsb5JQpb8MdHEk2187Kwtb9VK9PngjdLxd3vbEsj+Fdg
0Kt5ndcmjVPuaPz6cYxVvO/PeV3uEFvMMWQyXb3u3sKE6rkvD/fkgK6mUmKww+ow
hgpyEpBff6/xnTsPOE2ZBhbiR1EtdeNHvnpnyM0ae9eOBgSfXNv/9I9gzI19fUQ2

`pragma protect end_protected
