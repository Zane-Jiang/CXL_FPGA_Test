// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
PplCTfj7k2/cljSicqwWw2WbD6Ae0vXv6esyTDZJB54yUemYLTquxVhKSGSdIO0i
zW7Z102WIne0MX858jRhI+fkZvJ+SoY9X9RSnOktCnqwaBY6u/QBVwTi93hvVT2c
obiWTDk8tlsZnIy35y+53dyRjYRfal1XHr/fFi3e2ww=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11280 )
`pragma protect data_block
K3Dg+n3npAXjeJwggQIUPykXHYQNPdEB5jPzm1XYnqUXy0Hn55CnvHdg/XG0aIC+
kPm0IdgbBkcE3mgVbXjW28neYgiy/4yhRBbSBH1aGKvHhbywISbcMM1RyO+ClWzT
0aGIqiBKo+SHzKcm/lnR3GeRa3PtZrPfTG//JVRcmYxzeDAwvJXzBAu4PI1XhIf8
P5s2YsUUqDkK3qzCN5a+3oLfrgSar/UbnWu9uvkttRr4PiMRI3IELkll16DwEjJS
VHaoilxhUoQTXKGfeE0jNNarP2qE/oHUT2N8ejwiIzc6JlPKsVVMnvw2oOl7S+Sv
tzvxt186xz6/lWebETzYGvSbicagpSnJg9DJK0j+aYUKuGJy84/nVsxdDnbN7gEt
7dvU16gwUpLbdThJonpLnabJ/B4griGIYhqSlnIY+lWRvSrmoeV8Bo2EESUFekch
cZfnVb9dB7+x7Psqwi6f+MZ5AmXJNDfaIxwGJBkpFLLpHtK6I0Yt6LL61u6ikFjU
NGZ+/+oO29bwjZIjdWXByvNHI8PiiHpjNGW8W+00tHTjsGS3Xv83Ql4u2Pan2+rR
hYRpgRZ4yvN0L+gYsgIdIOsEvon2dkujbl/7VW+AsRv6dIYRZztb3iPlQY06xEDi
x04CUJW4GXn5/G33vIWOjGIXuSIubAKrH1i7BRZ/Q3SUlQUxGFQ56Euw9aDg0rtM
NuQf1z0l3la2DhGofFqjOv+vb6qiNVjI2bONlzRQBy/QIOIorR1G8tUx70IJ1ZjF
dEQgLySsHISGRAMRDz7bMac0Xoi1YSD49JfW1cBGv2mznRIG+uYt/8IVEinTeda0
n4MiDjkfgRmFU4sn1sT9JlBH1oA16+0//o/f/YYZNm4HGb2Ffs0bU28INqmHtVks
6r/lL09rH8bz8E1bUF1gjXHJix8OcGbjtTGqiTKSHhVMrZWJUpdM1MptjM0cHCoF
myN3kQlc0ogqhKQSHVYmlN4o9S9GB/vdyYldtk7rrHj491YHkQXYd4i4aeTNqP3r
jB/ZMnzMpJcAWZ9FrI2G3MHN0J56Tp+u7ADLPobrhm99u5pz4xXdwLjhAEA09Goy
VSR5q4g27zerndoBnAieebmiZleadU8ynLD1oh/blJ3x0yDHQ/xL7hWNq8ZX2im5
oAzd+0ui6KlKpG+lzWVOJPfODRxdGvW5dSQLYMxKnJ+/5W1AgDy4KIGt67mRZr2V
V4Cz7h4PpdMd3GLx5OuqzOeg5P7jSVKp4CiuVQiuaZaMPoIRWCMditaYoxwKZHYZ
3SNkwrQuGLzTqkm7uPEaGRGUgtjJLTsO+obmhybnfiO8E9vbvqbVVX30YT9cPqjN
rK0Z6HMi1wwoQTc+xqoOyx3AOPQB6Fi6HKbeC11Hc6L5cX7fv921yP1NdBrbpuiI
ZWzpFV8z3GcFTlz2q1Qovz9jHNTktdJoA8Wsjpm+CtunIJnrBoibctVvSN6AHxDq
6dOA5/n25VlvAx5me/TGohKsFDEjC9YlwSFWlrZkiCczhCOHkCrwYkN1L5UBUQLX
tmtW5OxKWpjrQouAxFO7qRC5GHuPbqJCqDCICuBPvoVxT1vWiQVuHmGKcpmMA6fo
lFjt8GXRvid4rpqh4P2F/Mh35xj+/h6WoZyyI5KUMLlsJIW5IGZupUe4xP+TdY8y
cSAvD1fpYcFP8TSnG5E2iV/IYPoNurAJaumMnvtO3JS8T8NpBrVz+pjMIcgzwl9B
SRWxBvpY2u10OaRD1Xf7Xao8GZEJ2VPwyOwgq4uDa2Fty6IYRKGVr4uo4eEHrmrt
X8ZibkGdi/AtS/WEw4z/aaqEaJS4zEsWi9Vo1eG2Ugeep/paUwdl1R0pIYCxydka
F9YueWiDo0NEcCfYCJiH+xYobOLqRetJG9R+JyYUTf2xJs6SZpTvjSt5tjWjsM+M
cbrSAmulKZModVhw1xloS/OLfSIVe3JWJRaVrJDArlIh8l5TJbI/mSg0Gw/3fgXz
kJY+FLHFa29L+Qr2XxgwvmTUlaPm72lEq476zw3FlJBwIAeH686ndA4i45MsFJ01
A9lrIETsp8vS2mlHSzjlEPDW3tUOTBAOHkFq6G95u3WKA3esNZTGD6oAJe8YEdwv
x9hrjE+YDuB61QmtjaI3sS1iWXSBBTLuNmMtCO/W+0AX+JFqyVvajsa8zcqG0yCK
tF/o7fk0JRLXSU2+4aGO1c5fh0ymH9iXXDEYs/hQJ/7el3S56BBmUJSzKROV8tUL
1E+9qBr2ysJ5KsPwDPLsGZGQvzWAnVgh0izjP1prMrnAJq7prhGyWbExDF8eL+fy
OCjDjowMuvBSj/U1c2IOsnB65ziLpu/C9M1AzlhwNNRZqIe5w7q29FREA3QuZtSH
3EzlF7KNzBcY1alqOuhqyD3U6yhED1gq5xSw+8fI8scjc95JTqRwvKPBASTIJHln
N05/d92otp1LDs0MST1xSiJZI6pkyxGQpGhuz++9jEbYldjnXnUSR0ID6ujB+Zba
EUMSS+ILxT7pDz30m2FtQ4nlG6mxOsmVgDO5XpeQbHarLQD/j5zow0vclBqH6PN8
+GA+rhTW/4Xrg00JW+RyAPthxBc8tANrIeYgSAbIeAu56VHN26kGvlnMJhMzi8yP
XjIVtf2L4m5+0L8j5rlcctIMRd9vWJszrx3+2fv30wWLlhpLRRYfFVBTakFbg4UY
ybG3VE2xUtiqLDnghWtX6Olg+m4bHGulUB5UP5B/y0Hzd0vBIn2VG3HljG0shWqk
58YMoXw7ylNivwfbNlV1LltaSQPE71bB8ak8zkJu19QuAScQuZV8nM9E4Mqyyety
XpTb0zBcTL58VS6kTNKn53NeV6vDCBDQkTYmhlBiqno/zkQio2uxs2jPc40DqOtb
A/PrRrkf0BQvDaOajhsijUJVK095I/u3lY4PZfHtLJ+9k4X0wxAQpSNxphyrX21O
aby10hAU+8hlly6Dq8D+F4INaIc18CANMLfMFuIaarh1QhlBdSTwP52dyMvnoPn9
/zaG3h8g1C0zko7OD9r32mwfCcgbqIMsW1YG5xJ0ujrB4YRnFlx1NScEU2Cac6NC
GXiVwLFG9kJgTD9vAEaZnQFOrEEIPEuLBU9GaR8GXej2zsDDl6PUH5iYigsPHWmD
5lSc/YAuFdMlulV2X+gqUrWNU8XHcjW0lPIp0a9gOf31ujTO7/1IwIoLGzOdCKx2
3kTbC3teKvlBV1KKN/M+jYLTjp6VSmKrV763sFjgXOlCF7tXunr9X7v63EslRa3t
fJQcnh8n05uP7igP3DKMzTGK3ptq1QNOwx/qOv8FbSblmWcomwjCYcggZ16WewU1
WwBnAnP2w2BHuI6nhTdN9guZpML9B7H/CaZHnTni/KpEY0V+z4IszcIBX4T+DOIG
4E3+tERiS25ggnPv52wlvrSLgcL3SjrC4uULxbFJ50avvNKfxgneL2e3kRyzvR1U
JC0BFy0AoFH46Ch8tA/nDIKQyjFkTTg/KJXl2aDGBv1e7Q3udW8EFt/WZrq6yLTX
s4UaNvPv2mtrKjb0mnK8xHGIy8WfE4oXJP4btIOLKtHKxCSCAqknbU6x46E9f0mP
cdPy0Xd8kuGWqdF2zRyyzdFpwnq3JqaxPSO0ZozpS/aFyVqpyuiTcaI30NIqnp+n
qiWrqZRNyM0xqIbDt/PkNmvPPzVhVcEnLCO9afXiGvyX28D9SvE7m/2Iu1Dnqi4q
PjUyK/v7+GhVvy7GNtQj1mb8++8h7tBOeSoMYOa0RV0nSIwfoFjuTZ2cAXCtTLZ9
YK6GzqdpQO31Bao4+rZdZSoCn4VXRHeSaTsi69ZAOaiI2SFqfzux3JQiTyLkPL+o
Fcu76+dYwPaQAiMnTK2wbtBE+iCAaqX8Q0OgyI13VVtDzlpIjxkpsW+OpqRaXI7Z
Leqg0U9FHpGP+qVMXlx2Y6Lf2D+vzxhcYl+DuqXSi/uayVd3fkmjf8IaQ3V9sInZ
QLyi2a4CX4ScRKmaqpzd1PTrtiXbUBpW9ttzIwS7z1NWxEkNsSSnwCiuI6LLHorX
53ihf/d3FpEYSqI4i+OOyX0XcdovS8hFjLeh8zBfYgrfYvmA1qe/4NG4dVFVagYr
OQ/FddKMOQBdr0RlInmo4oeo7Co+IgfdXJ4Xa3qivZHZDrgIDVFvH0UzIm4L+8At
ztqXNuXSuvB0Hv0YVnlZH6UXGt1a239LW/Kf8jTpLDpwYXvh+tdqZFrRbXsgp3JK
GNSSqq9BHk/VVnXVGe2Dij99Sve8XjGpHANW18GUX8qJdORR1gLv+SJl2kxMh/h0
5vvxxHwCkLQQHIaPiOkZXxeeQzswZ0sD81IEZ5gdjPXvi6q5e/co5UY+WUcB67gg
1vgYJtYcU8HUktlWXxPFvjEIJRqoLoOJTFc18A9B8XlLHA65D5Yb6GGmRtpklueX
PK0QS2t0eclSqfKB6ubQBKygiK8rUX9fgMmQWTjjTvI4lmpiHquGKlkS+RrPaq0U
eDW+Bxvcv3p7SFXyYSYq6I5icbSbUcO5677U60xBnTJt5S0zYB4ZXJ7o117Q4aeX
LqPc3NlaZVXJArjzb9nMGA+W/+4PZxPle/dcWwm21Q6qN7mHwX2mJ2frzLmi3tQb
mI7JLXTLI+KDqxB1dBpUwW6Tj8Qz+r6CrXUwNrWLj98jwPhKPuzDJb5/9ogV5AXE
+CI4kc/HZtn0+bvTG7chpM0u11StkkD5rOlbBg7iQKExLslvL28Tvo21muzxKLQf
hZTnqodkigw1zYMqvRwFSRn7FY869TMdu6dsRyTId2gqT/q3uiMCTutrA2vRO0WE
AZTsdxNjaCM2omkCQPRd7b6q7iloax5/0ECgc/28yd7rt3Cxs2raUWAhJr0hfv59
e7DkIGiW9cfRVaoX8SZJMKFKqGjgVjqHkg9liiZYr8KxzR1p15nvAChQ1Mm2/o1P
RK9wwW/Pf8CBHa1/mDbC1JDxuVAZTcXxg67ZBGcy17ZHj+bmPEVsxG2BnwYf49EK
ho8fQwy0le4ZeUFjIYAeWChO+e4/VEg3UZXvcD+KQdVxd2BTKH6J+LbHRkiVfkCx
HMwFC+O8WkIHkBtIyD6JWCTN6w1KR8chuRoMqBqWnECTuuy/2ZiiQHtavHQMjGq+
sLuwLN4iNDKpgufTKdkWpvHdrlhIaYpO67TwxAKKDTY+dRUHg4Rgbsini86uq8Fx
PThGoMLnVYNgo4OnMpIItRlgeXFhKmI49OMiYHXGIi+MyH3iuM/uQU7PixhgnlXV
SMwHAGBdkCfeZcLflX1TWH6xIx5gxFwy0/unBJcOfRJSj5OSbDaV3TCGVK+wgQCd
Sns3EYQvRPJ57AAsa5tXOuOamasWyNdp/saeHr6nCcOckAi8f67tSnFJlmdmS8q+
44mPWdSm9DoOvOekfe7yuDzzdv9s1TODU1Kmu3fStsURTbRsUYQFgGhodxbscMrR
mhfl/cvkxR82IMYXAis9fXlaKX5LjvPp1fGnOQ87oQK6LhWXhuEOs5WgVCWbDU5k
6lArH2TJ711aUX1y8c7zf4xzmux0ty7qMuM8dd8L95b70ffZ8kjw7Y9pTSR0d+YY
IlGjYPEv24XpwzsCNz33Fa57xpnsV6FERI8DFTOZNp2LyJENGStyjKeH+7JLo1vd
CqQBtpHba1nTSHAx+YK6O3ZMSmsKhQ66tlcwxO0d/5kNfI6eO85RNcRacNDezKh4
9OVflSMChznqyL9FCIupUrn+eca3K25FvfEVqY6DoQO+mgHOnP1ECzLetDnNGFR7
QsnH5txGuodZnuWadnZYNMynYHgCmoGp6n+Ka52Q0yEcxbqf/QDUuLpwOxJZMaEP
J9+BIV7fwTNJFUu03v3NvVB15WVCa3x6px5EEbvWj3U4mqN+uTroI++a0RXBd5tD
puD5WLNTuvPXc/BlXr7l0T8lck0Kg37W251EiyX8AKB/iBsCqeDx+J/gt3MjkAHH
nqo18BoXC8izk60jtEZaUpILVdCo7O+X5bGv6GPmwOZ5gCF+KRFrxrCbPn34eeug
ymrLSlDxtGZ3ap5iFlRtUjJ9IhPbWJtatPaQOU8FcLQfKa+ESf5xYfuAlUOhC+bA
xQ+SSnVCD2Yafm4aJ8360Aa7PCS9MXl79MNiP4n5/aXLNj2r747cVI2vBpafcZ0/
7W0L0q3eTBfe7hMwI8dm8AyPltk62vX/SRynTdPeXPZ2oAxLfW4378pzSOE+qr3u
Ab0au8PPEPbNOFwaTx/GSu8sTBl9VCgnIKVL7AqoRIHL+YFtaIW/5KJncgMOHOKT
8T/++G158dhap3uRMdR1bdBpeejfB+o90QaETBYTJUbZjlD5JDKAamlj5Boq7Cop
fYPSrh1/JE7aBObV1Auc2kFY7V5xxXMRDatvbowb90FW7+eJDsE7MuSVQq+GMpib
GjguwNjkM479sN0L5HvsEjwNgi6SzI3IkQfGeExT2FY/2FhDFxNmUlufq+BdwmHc
gkAZxwlxXNPlfj20NgLuyitYNlZB9oQzcS8yk0zzAp4JZtR2DPmePfov4iAHZscs
5w31Wh/6+GqBh9CVuHJQaSg12B3xuBxCL5rUaiRNKi/MRxMusr7AYGzhImGGwhlm
MXjU7VzXXAcVbUJY9pLt6V+akwMp19flzRue7oba6TB4qrJbxLvUP2u0gsYlD97i
/AR6MpodoMVYOYKElwyZLQNVIKjls+G4xxuH1C4VeHgz5wZGX3dtj9xVim2/dpTA
kNEiU5qYQemIgP/WbfbO1Oi6MLaibpOC8+cpIthiddY26vXCtqHJKbcvhXb3A99G
vFIx/E/q9pNWjgzRA/LdHD4qvVnBzNfagijk05nezYOhoabHF0tGbIqosuuebCNc
xTbZPtV6WGbFuPAhz4c8AUpwAv0bmPYNPuUrGspZuN7BXr1I2Uvrm8tlzuL/3Rfe
19cnK4W9+4G7en+oqX1675YZ9A1yrkUdPruBlUqwcUuUmiLHuTpGbSjNPdzpbkEi
O+ToAVL1LIMsJ0LR0GwZGwzLPbu5TxsnSfD9IJrhyJWvXfcqxjBwSuxDJ6hCXVRF
4IG9O5OyImtx+AObgSQT0ypo3TDkrYtqy6VueUklQ09YoH0lvDxwqcl3s3i9qhsn
kz3syoUhFxG9mvGvORBmpCLHzFzt537Kyg6sMQbiRGRbYMjv1wIxY1hIKifXttHq
+UQk1r1NpivgAbqNA2hbxTExFRqYJmN3rzh2Kksq+UZKsFqmDeObf6vSn+FiDv1R
UP7q+MhpE34V2Jm7pbaMOW0FXh3zmbnxTLwZ/q7ikx6Yk1+z30PmgooVqP7t7URF
XLFj3L4c3B2e3NmCJC/D20CcynGWu8W0q18gK1/nKYGMQh22CZS2u/tYz5Q7CdwW
h9yrpkOqPQJ9ioFaQ2g5e8oIIMsOj930wP8WX6SL5GnQ82wyPYPW0zK9V9H5fC53
yLKdjMMUNRaHX7RO2tmQkqQg0UP4aDtYYqQLrtgLMTlDXAKou8Fwy0AsgdRUsOkO
AWKzqhpyNPEP+2JZD4dEheyQhKKVwm3jDuUJI1Y2j1KlnddCuCMaGrKK51jxhIa+
sM67cn7/pe/MbN8glOf6DUpJhGrlVNe2yPAv66jZhIweiIL6ikE3czicsZoyZl6J
TTA7ziF5gL77mumRFi9TGWakWFKkg+f0QbHmmPNB7M+qeLE6jtwNCzFm8c4fp4Sm
S1axp7F7B2g/MA2B/uo8L7vCJTHxI2N3cqAtFEb3RhT3f4crqQTSsPVffJ5TLX3a
PInb4c75Ap+Rr9oEnta2n855XhsQxWrNgxcMkMRjJKGWL7HgNpIxcJkYSk2m3cQd
kjNbJmm4UVklL7wE0NiNI0OyI3kyPR8bD6ovu1Jlffj324XUIvwnUfGXGLPmdU3o
EbMhp/aEPbAV7SIrHXTVDdfFVg31GTovEsllrjHZV7kfngT5WknMIOSQmCrgagzp
9e7282m83y62zo5/WjgiyQ3K27q71KjQ/BlWTrQBM1SeHAITiKMVmbNkkRs2QrP2
AQnWFC26Pyp5XleiZsqqZ7F4nCrQNFMZ0ezA9oNlnF4oOxeV1hSEARuQw6uxfszk
tysJ2OiinYCptW/j1VlA3qiV8JeJIGcxgZ+tODopMgZwCEPvtHyp3ygrB2LlAga1
ndCrGFtA4JfEdgZvFOvM5JvdvCV6IAc1TYzWo2pTGqeoBzNPLaOMiw4o6eaT9CMi
scHAucJNn40IuP6cmLxU6cDTcPPpkJTaUGcLvWxHjzpVlxVA2vp2wEQ/e2/DTgSR
9Jz8uGLWYoZEtuHhrVoy5zFxcM03dj0nkEEdqqSE8oKJvdHsJOfY1N/vv69jdxjx
lvFYYAfEDt9PKVdJExdAPZ81m7m07+BYOEo6wDIlEdUpHyYCwcp3ZSWwG+I+YM5U
9B4dlVONeulukaAc/2ORFSxXVaRAAYP+kzhHTX/gC+tAIFYX9DJmztp/Ck8SexJ8
pjIQrx6CoFYh3GJO6usyXVxQlJC8vllzgpsNPvh4TWU2l4o9vmmR71HJGtB//xUC
tn5vH9kMrEUbE6GhguWlMGH3fFkQYI8FfVSdY9H+FmmJHsls9IVHKfECDiebD0CD
q7t3UJaoMeMHEsuPtHJD30T9dpzSZy0S83tSCoPBmPqHa/FzXUA0+Cze3q62BQV7
Hw9f+1KuwTgt6DNQY8JmeXY7wwrDN99FieVaUoju5Q65DF3hSAJdRwKwGY4Yk7jB
ZkQ9oEpQVkEur3TUfWGRXbkMxJcYVKL3e/mWZ3f9scljzKpkYTaUa4pybQh+H9fL
8bJB0Ewx+V1zBj94aaM49jRGjLwFymad5v0TjFLEs7wrjNCuf6AQMCOUVK1yJzbr
rmD9OelwifaU5gNzubsl580dZ6XB2zZCSM7wGb4EdVazve/z1+X5TQy3IDDf9sGp
O+MrMo2xm/ULk8WtgXhsV34us3mbs1YRBi51njaRvrkbd3gN8kIi+Fmx8YQtb++i
svJypoFyPBPqKfxRzy2ZeJmgzAIAPUFVwEpRngGzDwya2tHox+CGGdHy1zs9SS43
D6Y/i2BWEmTKTqaTjbg8vL47EoND9/4drcGK2Q/MW9zbh7Da8pS8Ji3zWEFH4Fju
LbTpHacPUsYWTjWIUJdyfXa9zWn64E+XGe5VJU/bo8FGqgOECIaFbbnq81S3HHGF
jRFvG6sN7koeHLCoB6dChd0+I05O1cdLOkzGqUC+V1rvdf5nTY9L4KylNOcdyS8y
qmtvdJiiOXwDD4mUxA/UlkL6UxatxBo4B4450Gn3WMw5+odPUOOFDvYnOurrYp5o
uFeEJRtv0zALLdUnDobbE/3rfoe0ztn7ZVMHz20iwtbIaOu+K5txnYBl42T1jPtX
5nlMI4NOy49tmVDc4Yz6Ot7I/ct+q/A+Rep7KI6aFUgtc3NfhBf5niVs0uYMQuxV
neIgWV9pJxAczx/bvgnfUj3lz9wCfixDZVVPmcDLHFjLjE8+q6JR7vIMMI6c4iBd
DEaKCbRAYKpFWF+3HZSwYggwDSkjw6yhUbMvaI6Nv0Tzlrq74Hr+YzEwhdixW97v
L1wzYYTwa9ai1ehDlcRn9LxAGPWkc/8eJvC98PtfhH5JfyNXy8TCQz9seuLkhNBa
GbaARB5rwCGZ9Odu1sHEC3e66WDwRDTwKwKiFBLkPQzEz/HcxJxCKzEnaXub9/+u
+/1w8Xu8R9HBhc4jkgkGCFYTALzU+fqBoRQAAt3u4O6NTQXBc/4d+UjQ6/J/kv3+
0eZDBh5WRbOf/d/ptoPzabeJ7EyurW+72iuUwwfFX5/fY2440TDjE632PMJiR4na
efcZ3Urwfx+Kbw3MlQH5JEBL351+qKTNKKKDrOsx1nyuCcXr3fuV0no3xtJW7pyH
JZBeMxqRVJfbaQcJ5PDFTklh5oqcJ0LDI4lqfKXIT5FsF/t+fqoreQcqS7yly0Ps
bqWFJGFiu3mFK0NgKWvzn25a4l3JMWCPamtlfqZgPLCPR97iL558hp6YursklQ4g
kJFTcdezAOdD2Kz30+J3rCGyMmE9hc+nSRF0szbPR51+ufz3F0ydflhmQJADFK2c
8n9GQWqx+G1DycIriN2ckUNtAiXLRzHwujN0BgL/iG7g50jMsRDtJhrjmGjcgIZ2
yqqINiCycZjrCgqT0Ua7o1023Acb4cgnryk0FGn1fstQjJyBLRhkcWR4NAAA1w1E
XVG1/6DEa71yx76B2A06wcX6C5Wgtp+AQ4T75RVJU6nN5IbOjnDFfFDkrQHZeFCq
4Q1ZlY9NJ1w3AzVlYFBiaEhn+xM/v7RPdIh9Aya5h0AqbkEM/czaEl6Ei4Fttxio
/YerZ6dr3mNf3FNaXiPuxiRsonEo4R2nE79GACUNrM2yuP2IHmlenMM+OZvYYH+T
5SqkDbQJvGh+KTzPCbB9aVH9I09iQPNYiCz/HXBmtWoxulildZlEaO2buu4o0hjD
6ihGzka9C618OzJk1EgIU5xJRgK2RUkfG73BeQUuX9/v1iBpCYMUMuYZBoy+2Ntj
L5xa0EIOH0HyI5UAacrEOtPkT7WJDcRjB7g9I3tpRjYOXvzr/4WbE1n06MS9lMKQ
D6Jm0iIqeSFNL1XqBseyiOQn+U1YgZmnltvjk7OCmLPkUr6m+CWBJ+19nXklsasA
zB1EVi/Nt+5cBDOtUyPt761nw16rwDihh5URvRh5EfqPRe2zljCd5wJiuwiIzblF
LOLykUHVL3A2IdCMbeYeT8zoqPRblwr0djph8saC1eApFSOnFakqowLIfeU1vkN6
SjQGqoZSY6wwTSc+eri5Fzz5LF9Mfm4CbC3ExjhcnCKo1Okj/N/l+RsS8T1cjOzt
LQqLcr9YgZaTlSrbSSOp5CNCPSwVHbjpndQ7Rl5efZK74y98YfpF83ixF823Aq1l
4SYOVwImb5CqTpLfB8TzRo6AQpraTU9n1ari4xTtpRijJ5EJIxDy1pGL/LNcJ3tK
an2avG5kt/0FNLh/xnAcDqPw36nKvMtaVZ+FqB4KEEZO6FE5n3b1wR/M7iFXqIG+
zoCI5ecSL8US0MpvPfTC76J5pYXyutQu4eVET+zcXhEqho7gxP+//D2LJwOm94k+
SHXkPQnDn4fAaqo+aTrGcHJiZrV2nvoYwOgXQ65XIYIu/Le2ZynM5n7zu8wOeeHd
YNYg3NU0BB/IVvYTnuUNlXQmdTETFEuT8hRB5f4AH+CIbNGXH/f7k5nP6t58+m9/
puLmp5iVhMdVbAG3gfukKJNkjE/0AIGSwdaWL7jLv1pg5X+pdpQhtQgud9qiPBG6
LzDjsvvGz/n0xXrok2Yyu7RvCHZVW44jsCHZqul7sd6w4IZxhAgSd9Y+rlhovRP4
XOzoJulsIONjFDxtn9EdgX9jFeqWO13ACviazUxKwmk3Fh03HxjNQVhDh4D+N1Ax
S2dJw1r+A+C+f76sYlextOMv+8aalAUhyO4EB9+HJMwJSPRnAZvEwjgKntD+5sup
mHKSV9wt8ztydPHGDyuAbtcTVMQ3KpyN8mGXSmk2EbCDXCbWcf88ZsI/153S/dqO
v6mAbF45VCoIdjuzA4h2FVTE7I0CZsnHhGcOjSsfyeyJFxWvMgmXO7x6Vb3kLGIP
A9/4PbYVQ6nmEswiX9gqOgbA/pT2VVjrIOIgfEZeNXTiwUuXEKw+TvYBThGh7yEG
iMttzFH/b9t+XolwTG2jqi50JOmldJ5QmIFA9nunuVSXbkHR28dcZnjkpe32WXh7
RGYEaf977SP4s/+WAH/q0eS3gT6/sdhC4cVRcJcgEdR97d9gehRmb5xgv33XrWHn
377mtFVwddyoE48S6eX9xO4QqtJVSgWTAXJTNaxCfbvnCjDdXMfhp43G6FKhxQl1
AHlFLDu8emT7b3aqPDpdKDo601Py9qi5YCk9+udziQNdANmSGBOhrzBDbBZyFPoQ
hDTn/1MSgbfTHly59HiYo3bQX7J4vw8EQ731YBbj0cs7XPvow6PCeHv38EfFftZk
h+6hamZaRsAp7yNYUq5JJkkVTYDH8XXtiOS8XsPAMDX+rkGRwqpq30vXYbgFzc67
oxdEzEUEm9BeZLQ4OPaM7PFitTYGpYetqeyab2KHx3IGrIS2Va2KhPSHI+KG0Svf
sYt2QrLUqOkLjCbirM1RrJXXGJTmfwCmPhn7WOxp6K8cfNbc3U5f4pYjbyGkKxWn
kfltgPTN3PPoeDyFkyVi0rmhCoADAFf/XGhmc5R8ET1YPKg92FRT96NqPauGltIl
zNbnGRX7gk/y3BKBdLrjZayZge/rzvalW0bmM/+7GOU0bT8C88dxrh1ETRcq6WP8
izjOdMqVni6p2LazFgkbJYkb3MvogBaUfI+BHNuxmBfqWPXfvYV2OImtUsxZnsCW
C7ikIlsJEr6270ZzEgyWJxV4PJca91ye0dI6iR5wR5cXBjyr1npwuf8xNuUQ8hDV
abvd4WKJMpk27irGQ8zfuR9oUYZIZFBxijLX1E1kgW5glTDuDZIzx88urX+ULtLI
xGJKMelebsfDkoHtHZenVjALGyaaXSUpYQ+CLwQiN60ZSk/EY4m92e7ZUCIn/Z2U
yKK/iHAOWSvc2uxoz0m0BiAYGPAP2EZREnqvVKwxZ1D1JHbtQgQDZ1nms2p0NkbZ
aBy/8XyteEGv3OXlyIZyyHr+IUUPtZk8xsKk37+fh6btQIwXRB8EprxswkswwF9X
ap5j573VT9bG9t5h1VrQZGt/MIgl5Bcz5dhnXOOTCZTojJT1sVaj16WyJbpGBV8Y
d8IKoeI1G9vymNw32Qz+kLIAabVx3JBzH3XCYqQo+QMLnwvskt8m3X7bSPXsJFwA
UF0BBXx1BZL06dAtA2qKOBVTZCB7RevxHXo9Mgs+f715DTHDRAkzWKh6js7zrGou
2rba5RRIfcbcMny267n9Qk4ta9jgfGQdtG7W8mKyOgRr0UhUnr80/BYi0g/40CvY
JYJxOdggqNKuUC+FJ1FPiICt9tkMSvI4npWqIAf/4aQ8qrxFSc16EpJtXH0elHUX
9wQWJ+ry2DRl1/251cJwJvtNxVNUAtGjTWUJ/o0nXSHPt8YkPz6xMQQALWRlqHLC
pbcfa1fuejeoC7VkAp9yquWhqr+X8aHjXhYZ535U+VemFGD7kny5ibdOTGQmPgpT
6JSCp0zYwytNwcLqPCtBixKRYe3XZ70mUbzUoLGepIIKcqqxvWINkjsrHnUfZDU9
7KTh9oySfetoXb7Vu38lcvdX97emYjr9iGTxDlbPUYM3mU3VaCe9ZqXNnSdrPMTO
NEdIXVqGGp1GEGtOJgKlYUJgEGzvVJ7mkm9vG33HnoNUDCvl4LQ3Aqnr+CtyPRoR
Op5kqNwSWWR7wdPIJN/4NOfjcDgLQ2TH16JNkCyBjsT7EPurknTVCuUh3xbrMO8r
yS0rs2iS+N0p14w7REPhUYZnjZyMT6yPfom3XMlT8hKD4yzd3HI8X7IcG3LGB87T
PbLIkFmL6W7uRFONuem1cGRfbNfn0f6edMS8WiTQCXW+68aj7JuhnUybD2u69xHt
LKnDwYvv56X5jQ30SuDUtaA9C9PfSC27Ihime/Mz/I4t2F3PvizwOVltzBWD7Wf2
ot0mbyCFW4ELAFutBxK2FT492Q8NbB2RYeXbzNjq2Xzhz59UiM/SHxVY0+2e07XX
Ed3zSKov7bDVCxhOxIW7FTuem9DRUm9iXSB07XTvKKLMv09o68S8mcoZwv7Jhs2G
RqfLNcnOxKghehUatseW+xm0xj9aVGpd0zbmj6x6FES7VkIS84vFKWgq77Ee8547
t3nvJfF569j+bD1Fnis3gZ21H/UKvhgUhXBPvYkkZWQQGAwB5nsDeGWANirMLc/b
3CQ0Ksqvf7cKFIeVicWVF87pO/djlcuNq9gt3CQ6PBqvhj1JWaeFmCFZhEQ7h1bw
B4j4bf8iOOlpsQBeM1uhWzgXN1aeBMJHiL1LEy8zJceCaIzX2ceadIlrKdfY+mCw
ksuH46bgz2BNPKs/UsI43mRnzOfqS8E9QW08eD+HHsIQARjtx/yG7ltoP4nPuG3v
RAOlSQU1DU/CdBcLjumHBbJvT9e8sRKaNufTCxoS3LOlaJmVtiyj2IGd8tp+l9MT
HJqZuC4CCoUBIrsg7NrsMCYeLPTXgviCC6CFv2pbEZKwtovtS8PbDvba7YMbf03p
GLklPDdBPl2Y12Jk2MPR5MJ1FNKckSIaEd+hCY2Wi7AVmjjB9n5MCtkfCVheLpV4
Ega7ciwCUmd3pIZk9Yst2puhMzT6Gi15l2t+B686kz54xBD0jRNVnQIv0tjFnKm6
p2wVzAAHX0tYIc6M0YPDzf3wpuCZqjVsVcpnJgcyF7N7A55kNxabJtdtypzDePbu
sTTH9boVhDJ/bwjFIYNq7UjYRyvobzI/VOFgZtxyK5D32mMD0chLVa0FFrqK9TI/
qVJHjlwzWSVGWEILz3rV/d/B/QSccgz30Cjjk63SHbZ3punbFCXvptzvE0w5lp5B
zwikuE5MsRH/hS5zJ2BwPzGDLE03NfAw4WDs6JZvE9YE23MEFCv/IEyfwWgLBzGZ
jdCFhTTi6g/BXlgxX7fneHKm78N20fQYMqbqcryaCouiFtSeNrzI7DdxulEC6RX8
drhCM2itvyumuGZ5KWNuU/foDUBXm4qaTIGyCnO5BN5DTtToXEkG59GCRhE5AvXc
mKGmOkz7mr7o8iErhhf0idiOHdaZ8Dg1EsXJYXYice3CGG7Ywt5mTmd6WxvkoSJm
atDPkGaSLbmobit57JqeG4oe5sUmmtMlY0TsZSsOug5YhA0SIA5RMCHf56S/NZSl
63EfWW59PYB/Up9KoWeOJWwuRuNtltZ2+p+2ZOfaUjr9u0w7zUbCVvXD6Oy2Ejvb
3X/7KFu6SDRnBHiiPB17plhS1B0XGs2XCpJFQcKwHuJLFur7ZhRwm5qoTz4NiYYv
yYdQD/AqsxJ0Zj38Xz2tbMDpffj5vVqJ60oMivZ5Ds8mUKm3jD8Vz9scknlQh9VA
IrKpX8MX+SvpNeQHbkq+5LWnHn/29ijRGZmR/NXpLXjFahPvr2Mw07iKXTPOIzFq

`pragma protect end_protected
