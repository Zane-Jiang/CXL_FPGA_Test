// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GebxzslXwJL4fg41Rs5KExjgQ2WIokJdBh+1pOAhZsRtLa0tfxl/AiScbDP8gIRmjlQUQ1bTHNmg
mLNcxQS+k/CrbKl5RKagMqVc/+Kt9/TLh4piwzg2dN9pWu+epL89dhVTPOs0iicAc6Ovga2v7gGs
MlE/hMAsRLz/RiAwZ3drVLGdc5HpS7KTH3zcRlsQNn73SBkIn0Iq0M2KbEEqftR42zW7NtpCPLnw
fIPAylKeDpl2yPfidQLnAAzkPIjHFFtmgDAOsicKVbdIfMU9uCghzsRZGr8jJRaaK72dIOgctcOU
P1pFpNqbDNfi89J1r/DgBqwEeVNYG3kXetzPUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15472)
ifU98FZoZEOmfJ9cClwqioIcdoe+3ytDrXsb5JTRuCC1Ep7porCx5Vi4Pv2TX1h/f1k4z9fZQqLT
OJJM3PtxL4DR73LFppN17yyN8/ioPzXBNO5qZnBL6z3Qif1qSoPjQMVU7t/fN0HbUErP10pVTrZC
KhUDhU8tHYiAUoVGLUPq6tAtMtrS0qcdk+0scn0ENQl9d1cronVo697TjXTKd3t/X9//2wdxg+e6
j406gDW7y0UeZ1SZooeJMCSVdtUhsecOeLuT7MdKkiUGExSFNoNOYL5XJ16mfskhze1ENf6nrySQ
FliAZAhdf95cIuwTCG2aGLloW4+2dB4z8GRCjFYIh05dDnZMkKywBiV4MmjKgklSRzUNHAoqtyi4
thKC+0wv/ptWKtgo6+I3bQnZnNbaUP7iQvm0h7KHuG7Z/h7KMNRaGDNKbIXakxWIfyUeIM7qqc+i
Xh/vO2cxQBeNmMS7mvzgVmMr861y45jdHkzqiDLdAA7a4xai0twuJayTuHAV8igvbh/7Anp1DEFN
F/E/HFozwH1pPUU32NimzuFRDgeBOCvQFgsr+PzFNOAgnO+pSAcEUuxJN//A9lixsmdQLQ7wXfqY
BouEIBab2QNwt5RkzDdnWh+0llP3orTOnOI3gGij403f9wNhtInplzq9oon0/GuQDkqS1yxtP73Y
phFsRaEd/CQ0c2SSDEll7lgmm1eGqHHjEb6XSMrKS3FgFzILy4olMbsH52Jv+c6VskKwQhG8lELa
POd5hLgaqAXaVo2mtq0UNAXo4UYzMAHsHqEaj1pgHnyRUDINb1BsvM2RZH436I1lMRaqoezTg8zt
ae+TlywQkW4zKmY/ojKeTJOgAi9Ju5v/3iCPw8v3mFm2CDJwlO+lotL2/aWpSyAH70S97+FAhxLZ
KLZlKa0SJJXZXeOLs/inGjbjTbgRxLEcRL/a9lnuP8/QzdRrVSwEvKZ/mzveEvyrbXNdcrpRztr7
FICNfu7Hw1IPIUCmP0FD11aCx7mJC5fuPSkW93MKZIR2WKnUgqsVF+LL9BaMQUK9xFugQTaoOPG6
LNbOvWhCTGOWGOrCNYiYw5SbHE+yzp/gSOI+u0ocXoc45kb2MDtNnXSnyqRun+ht5Sezut9vofrQ
ktTXfMn5aW3satELO6vJXpGKMG1toUvW/0ElBYzOWeQ2KwX2vP1Qltq1kPXgjH8mSI0GuKRQuOBz
M9nh1IHCOwOi39pQsmLK/FjcMd0JH6lvxaHZydAjyeiMmPsvkQdrTw2HTBNFYjHqEqNQC26BSVQX
Wogw8d8fyh5egr8N9D5k3w071syjCK9oeawTedCbdcJSiyOuKf/8AftnaLk3ETcmpGB0Rubb/gMh
fYmyoLcBc2U8Lc5TIO11NiG22UiuVgMl2XhnCscc1uy6e4hOSDx3Wq97n1KPgZAwN7Au2Df8WgVV
qEKR3nRNmevAFjT2SWwY2bIkZrsrkK+FTUq0mf5xMrUS61o7ROu27rAD5itE7WtzhO097SooW4GS
FK2082rizCo0VjXUfrfd4usuewNOsl2Tw2p4C2qXI/Z/e6znl/l9eszx1B9cc5kIJa01uLy0MxXn
z8l7FtsDuwzXcMaDnxsuy+RxAwYWQ3IwPK8Tj0LlPw3i2QlOg4/iR8CtAedRCe8+TmSz0eG+BmfR
fRqMZzcIcC/imjmJFLk/+HKdXM4gsuNI/M9vDflfO/9Zjcc+YOygQJ+txSiVegj4iayvMOI4f5zj
tfT6waelvhSDE37IcNBoPCq6GE1bWdTGhdCc1VylwRiYhsR04egxF35YrkjVvt4Bnp15Y7TjJnvz
cfgGhPpnInGVuo/hjpciKmdg+fHLPLN/kORKV7rnNlnWLspHCk2OE8oRa1j1ltSubc73RSRiYOLh
utdRU+jDzgbgmyN0G0uzfK0MWST0Zt8GQp5EEpfZPJzZMW5xBrB44IQrxPQEbKSnRuaWvS9uvQIm
ixBNtLlfrElvQoJB/l+o/ct6im7D/wP7wGZy0e/zJSZMGsVvfTIxX62bzk0+52cGN/1P2i6BEdXD
OvPsqrosy4xFxLhvuGxpcb5/e802pV+OHnngZaHBnSqjtZ/4uzw0vPZv/fIpxQFjzhlMVE0XMnYN
YKn/NcRUPiRZcsTufHT7EkPM6ytLiK12CtZwPBKhFK+wTAMEtRO8nHX5qmJ8H0+N25BvG8nGGu8d
nyBl7PBkCD3VaLTu70PYiiEEp2ELhu/0QIMDRwQQiJnD4X4Wuk4w4IuMx/dGqnY7l8edBnXx4M6k
ZoBNgHgl6kfT0l+86POdVNh9IMegSzWIHiHhdDJ5Vrsh0jFjOdFM3Bx6lVR5KodY04PPXQ8lFJrX
bc9hsjmEVQ1ZlPnOKQJNJ1yv83nBtS8HUBm2kIiUvvwK6qm3Xqg0tKsTPZpCTBWczhwvFpGw7B3+
j+APuaSX8ZMGgxF3plNAv5FFay4x4cqiX6Xw8w+p1U2EH270poyJaoL/o7cp0/sL+2/T6dPjpDxu
xpkvpemVj2zfsnAfCStkB/3jIzvrJCdUSzqByGMH9weqc6Av8tyCefuaJcvyt2H9goK/FwmiRTDy
VkYPjMztIP6nVtm7O0bupTwUEY/CzZ1GJwtPyugGacBq/pQcqyi5TctklOQ+z0YjFK6k5PO+9R1b
zyz6Yhmh9xd78q0yJSN00zdrGu5fE9i8y806c1kwnVe66i7SoGPY70dytxgRJyQYOlxm4usvdSGN
orGDdeSPwT0ifC2y4rKH7I3K4Z4NqojOONNHjLKckZnRNgcJ5qSHzalWHmhkLBSVsDvIpUIaYXo6
PJmMVJvGf8Ta9JuA27JImIzsVu+Ui8Oz8VCWiI8fQY47CFodSS/o+XPM6N42Zbk3BYGZg67AzLtV
V3e4Pfa1c5sz5LfJR3U0Yy25FqifrT4BicVzxPCS1Nnh2YR3hbV+Sya0SqWvZTJNmztIPKNUN8ba
EjyS5N5wJGLUpZcXZimuTqqSNfXRaJEn7c3dlX3M3/8/KMrIOg73an4VCKZtKwEjytxXrzP+qT5b
ih6M5YPLrJ659DqiTtZoNale+1Z0oet77dvgWKWo11WyFYDpA+m/7qxxrnc7O4QhMrvjiicVjIcK
c2zfIPQJ9crp2IqXwS8sHwwEvp5RA8MoU+4yW/4sarvSC9ANYF9oSq7Q0gQ/0lOTbMyLz+6ZerNx
+UA2mOtgpZwUm+db5p2Z723JjJuP1RuBMt+OcczjVvDC5qbIL0W7M1o78Gc47+Y/409Yj2WeSD3H
Ze4JFr3VGfl4T5zc+kj0M4mvGEU1XBTZwkKJ1Ehpq1rqZC75hWvAziJg8E7Lv6vokMY1Crpf4aQo
mpAD+IjqGSSWChMPKGox7TxVfjoOH1upkb+dPivw1ZsG00DHxLuTpDEYLyEYOEgVACZryxZgpic4
dXH0OEvaWc0ojOOJInsgAMJrNNde6iRQbzcs4LaQvGO+fhlJSmSxYkSUDkBlEGpkSPrvZsCdkCNc
u/u+zcrhI+r3C80BkTUMCriIoTvbi4Bo2sorWymJ3tfgyUzuzhcrpwzw8eZyo4HWN3vcZwHlhA3I
CPDnenDLnPUYHyPTyECA3LN6XFwXXkhpR1lyiY7oa9gGXmKOtsbAlmWBhusFs5hX+52Azpikj5kt
70RrJ0AzYDvBx+qu2x42IDXXWWIvVjzYmUoHducbS5CDbu+qxcI+akVEvBH9O6eNSd0XiK44QV/8
rFZcYP4kmnQYITMTFACRYmhmcwOo8pVAPsJgpA8wkdWdH8A/0YU9RjaghULlOoPVXPOmDBHnOVHr
mwHsJgeUN1ifmmkcd2JpTmnoq9Ik8oZ36/KNx43KkwXhQYZuMZM66dyqoXzUAZfkQ1Mr1bJWy1wV
P+j0FulgqZBQYDdrjByYQyFG8GuE6NyaNpMLeS6yIoihS3YDprdG0M2FCJOfmt4Ot37ee/dofGuQ
EOjENM7zo3Bvg6LVrRQ1YsQUkibX0QRmMWcKYAtq+kGRceH2oKllkIcaAFViLuteeK/ajNrKhWIU
+mzBAWaC20kWe3xJXcZV1HnRzvexZAPhMNrKct0mnvjOXT0zkL0hvVaAMI3W9BlZqcKAAGlHHQVL
Mwjy4VbKbpxlhJIws8rfPmqd56cziQ2HuU1IAU8uLmksZ3g2GB4APMXVUEPv1JAZcsrOdHyEQdCN
ImnugOsVWeEzw/9ovGBP/qqlecA/Lr75P69TtmubFlAmbi6Rloduzw5XJSnNlgfldS80K2Nq1Vpe
4pNy/KCi+ln8vt/VrPcCQyTLKz1QbHb1P5WVbcwOOJxN3XMT/E6u5+iYjHFcFiqDVgPKAO7IuMoP
9az8bhNkxZ84U9slGLcqIEnO+9CH7tFcld5V55ypfZCalq6gWkEdMekJEFLNbGevIa5/JazZJ4FR
jBIea6X/rvy6CWKT6jXe6xolrmkuGbsGxNp9ZppN+w3eLtMIzRTsdmR8MWKbZd26OAM6CUaIieJv
j5BRRpR9NKzKqVfnNMX7G8BrTojxMusWWY6Wvtq0cXCtmMwOwBX1pAh2v0kjRppTTqKTWsXrKxz6
+gdYsdCgDM59eChEXdsc81AX9wpiQ3ldguTC3kyealuX4p3UIp7ZGyY8/jFg9ia5U1ZA5MzpEpxL
NLXdFQKqptu+Dymt/uznE5794Z4qKYCTPB/DefB8rk6j906JCI5z5ytJEsAP8lhuMp+wkAc4prpX
bU3EU2iITKrMCF6n5lCYXcnYJQqnqmZDFkbcAlF7SNJL3/RQc9CQZWPREMYs2Ta3HdIufrIROvSe
ajbqSLUkJ1FVoC2zierySQ8X3KWdOl3hYrjv7WNH7QbkkY6RdFBsYQq+mYI0z5+snhKF2xSS+iE1
7j44JEUiHgqFFDE7/fJj+quWx3uwKLf23ISrUabgVgmAYSMJh7ZGGMAeeI6IPq0MZF2VyhpHmlQI
R3wkYS8c03TnPPlW+UsXIJyr144Gh/v7VN5eSrKr/46QmwSi5/nRzboLxMExZNSMZKeasudyYG7+
/Oa+NIGVxrlQtIcYNSbRqNWPFILnKFYHvAWwzbBXBgnNMb6iSk/EoKELjD2MPgtEb9VU0pUWYNWd
MRT61jirQmoWZijhBVSHlFOcMsS5q8xbLPQTMGa4E6B6Ua8b17NGKSy+mv3m16020f3fi7NX/MQP
uLztwxs2+xo5Ki9qkXGrqTIP+qKwRWGnXAIilrELIj7+oZapYB7+VSSCrqEjedWVZuRw4R93nHtG
MnzeuBzedYi7Ym+1uSDmf+Y9Jq6CAVH4DviX90R1QwQT/pXHwjMLYngLp75mRoAaiexDap8zg//s
c7B5OOiSmJIXKnB5YR/eBGsIuDkSDEZGbjeOrGhgRfvkQNP4C788ab86fHTBhZlm6xO0DtWjzQ7r
VePHCjwLcV9yX61sOnVOwIpx8ipR9Rce5LdmE+6R0DKzJt53GND+D63k0boQR/7utm4seRsHFZK7
lgNCZWJFQoqpFSDsfHJnBF0LZE88OUjUwRm26nAfsGeHyS9YitgF91JKYqsshmZ7qaWa8DY1KY6a
1v+m1wiegqmQll/HDG3cqbBPx+1abLIf0RRUw8vIx81gRwRjdUU/iqnHay812XGCIMtdt1v667Td
Ag+Y+c5QWpoxBqUo412oDiAq+oYbRzLSKbOXjoBO+kxEqDRmu4pF14n97MdYA8dTGEbIWc7xC00l
v7C0hOerdxeVfCZUC6h38lK5n0vXUxAe+P7jRK6g/TbqDQ/UFJ2JuiT/aq0kKZv6gzJUVrOFiPEu
3HnGtEsW0TLo4PrkJU6NY35vc2nHJXr4d8d9aKKmdir5fvj1rBh9CDotLZtTw8zicNb857+SN4Jr
NQoedxPEPtKWBJvdGhIQCsvY1wejCdKIcCAVJ674Cp76PxR2LmrLlgaiLlZ7EbLQNC0xm556dUyZ
zbmihSjcAd3RYkmxD7N4oBlOc8MuoouOaYPEpNlhN9lE+e8eb/RDALJhE8VgzfxlllZb46Yq6E1Z
qwU8dM3TlG2MXpiKedY0Xg2Lmj6O4nv+kDCGb6dsugozDQ1+G11siydl+0pnYwyTGSQSCE3lMuxJ
MtKW4zEfjGC5Psa69Mar803ZSUBUoVhEGTI61z2g/c03S47i5i6QUmRN1nqMSIyHQbtTTZMoLCV5
WayW2T1wKMzN5RojuYkMygfmGewGNGwZPTBcUEm1NvqjpjRS9yXktbfXvSCZDPC1Xx6jxGVs2/AH
PJdLg6WCYqlnLip1byN8yKFY4GGN/IL46AN7Tn7tRWtb+NrJ+rDVC/O5vihhHeYUy1DW3R2eFsl8
gg443HeTRN57XL3PCYjPlBPWfUYuxneKcpQq4IT2Dw9Vo1HVKqHNWAbvNn8FzGUi/CkBOmtc11qn
yqzNSazd7G373GI2IwvYQEyXAzuQcoQ+QeLFu/O5N5juCYiM0DZ3tDz0OvxYha52mElAgY/ybL9L
JkKvAPnYaW6wE8VsghY5HgDwqjqy93KAxmVAeXF6vp/k7Pr5HvD2z7hZyoASBUCE9Ccw3mfYyWEv
vLFdj/63t1jwp0HWNmPhwUZjZtTYTwTmXCvY0pQFXry3xnzyRjwLNdqFvEIdenI6tmBXvoEmyKMX
/8H+GB0L197TR8Np5Nwi8B9nSgqjJ0wfhBlCfvqp0sL5UhKpw6WFjCEvRtDpKsEGPVOKkoQWqvci
VHu+mlg/pvR6WwlJJHI3VF+QNK+7wT//QzlIcMxwMnMtqWKsdlKt1Vz1MGdcW1HZV+GegwDW11hg
b7rT4G6u/cqFaEdBMohaAqYJZ383NDPIO0WoeAmfXmHkPExuTOyufnupjB8NN0SD43+f1S7ys6CV
xYFMLQ88f9x3DUD4+eSW+E2UYcmCELzTNp0hUSOf8Cxsthn+hUpkQu5ujmTyDFvFg7m9gv1Z7bO+
puGeMSlQCEVn43rqHpUqEMPPUnxYawC06oBhNKL29qFZvXZSEiTHlvWfruTdJ7GU1Vohd1ZbblX5
JVPfoEqqup1En8lH8zIvMbMa/lSFk2ECD/2Tw6M7c4Zue4zm8QpmllIh+B71ylNqMIM0KAF7Yv3A
QoRjFk6D7RaL61BtjdQ6UeVrvKctjPUCBsBp/AUY0CDlaiThp/sP48vQGeZUAfYnnzECQIZZJcvJ
sDqT9JU9oUvmuUNblyybZLQT80pXG+x8o/rTfC2/38yXAYGJiU8FvYW7WRQ+m5vOoHew/bQofyR7
Ey8gtNhlAq38JVSvqS2eOFRtRW+E3+ReoNjLG58HmCGDv052cCfDf2Gwvywib6+CL8yODxWi5Szj
DBP3H3ttrkWzWPP9k9i1pHxgBBDRrZ3/glkLIiccH2W3o54/Ksef2UNGSQhFj7cvxKcpb/FkGq5v
nsPoLjNukciNz42pj7xwiyBDsS73RgyC3aJBUoRdEIJ8Vw2sKBQJ91UCOinhs8KGKjIFS4vymuN+
EEhMqG4PSpBGamWIrfPgRcTr22N36M6YGLcllfBErptsNLLFrYRyMSzZXA+0lc/JkvsFowPYgVFv
66chAlNP3S1CUfDpLUmmEhaXILbfN84VuFqfCt4QNRcfUC+DEXZlHQIm08k4Zwfr1vtad1GrNb92
wE0Vje0JtJOcIcPWiPmvuOyX9NV2EvK8QwfIfxBtbJSe7lq31Z1cmF7Hwg964zX7dP6DtIYOC2H5
p9iytEQ21IFLtZ7dBlg9i6X1GRIlPvs6rnWIelJjAdWYdXF8HiN5MQC/QnBpz1ComI05yQLaOtyd
IFYmpDoBxkEjmYKt0hfgiFHmV8CtmFi+mNDDMA79moAUtTQ4/VnP/oon1UbdhQJtb9LTuZ0dkWQQ
HNb2CbqGPxji2zy5h8bbC3/emsaxYZwW6m5+Q20Fqk5bkVakD4uRyH9LFjiZgHOI2iSY83KToJ4S
X7ONA+G81iGuUt6vpLjjcSP8P+joWdUA45j/6EAnCn1+nzHLnnL7PC+xIRpmqk3VxfLhlXrBrJDR
wOth3aks4qEgpAIXK2mQTyIzlmo9bu7C9A4SNb0q9bQxW8lMN5X/Kooq1LcUEgyyzQ5rud5KIXi4
b23V+II8Ps3zIDGP7rcSsgsLXDiMzzHDR2W5O7iCQRf9VAAeUzQcucVjuV5pazPHtuwswqW8QUDq
JndmhH9277+bTraZAYPQKmPmtBqTvdLI09qBoKpRKTR6uoNTdr31U4NCo7GczTpazgdVBo5GsOra
Z2/6cl+BVb1Lz0cBibUGYqnf6ihh8jfEUXEsH4TXMV3p/U/ZUBVemkgmtdCnpXTHOvBCyTHsXHtx
XR+4j4pur5C4hapjhuxh1ffkMgSASczmKXQ84rT3BJU+ZKNi7bCN5rqVs99qDSU/iD7ZzThyE9U1
Xlw4C6NR6h5IVfJsLahTzG/+d61jXAJY7KfAyX+5WjTBsVCma0cPlPcn43ti0btz70xiqxpExCAD
YEYwz2eJUroQkfzYjeLJ38UQAW147uGBn+w9IGAD0DQXY2a06go31nartZal/izOsS85uuen7oJI
tmamzbRue/7jEZphfuby6UzblXlOq/WPqG8kjW4KNbizx7Y8+p9eWeMkh7l/i+R3ucz8JzkkFBoo
BlL1SKLQlsYjYO2sjlh05SF/jLczPBn8VpXli4hWfaj3J1djrciNDJCQ6dhTkmngRlQDbp8B1fi+
66e3hfLeFmrs43D4vDxN50x37q2ydQQkCHpCPRsWjkXNPbIrboBsxbRVZhbo7W0CxPzfF8xF09Yu
C7RnmG7YKJwmOx9DjbZh45shG3K7QzZTrxo2oc7FFL35UtEv5Q8+2OPXgJ3sDk95Ej7CFyYd4QND
vTVK+irqd25MEgAAhoo9IcUYeQIfAJx3T7VDTeaF3lLpg0ST0UMBVkzxviY4BC+bNqEKH03iAtxk
+cMkdAwoF7ukvQlmugLzehbM1cPJF9xk6wYOHfTTO9Y/BCbt1IjidR9wdacUPBIe3ethim9hvPgW
ltI53hq3n0NgeByhwAiBVnn148KPZ0hxothz32ilTuTJaKRfcE2ynUYKjrWDO/x+9SFz/K8SHy/G
FJgoNxWgxkAC4bIwjvuuVGAYCqILrqjKdJk7zS1jkJsbmqxcEMxDV/VVjj5YXnBj38do+rPvrxwV
JZeKO6eNS5JE790M+24KCbe+A5PpjDIRgOvKbzhKT0DQ9synngHuP9ExKT+76hyt3HcK2oZOQlUA
j+4pR+dMwSGAQq51Kl2HHG6JTaOVrHQDACAr0xGHyjV8GYJ83iO5jA8MLuiO1rNKiHCg7fgt46Pe
xSBb4kzOuSsS93lh+iRDTO1qeryRGpzhB1BFETewzfxGHQZe2q2oG03Etl3c6gCxhmrzIt8byzVk
UhjsXf9EOiJMoK40ZgV8bbAEHaUvCb9h5dxQu+4xuFYfwp3DFukn5HczKLnP/F2Ph6XSQYViqTlU
vxHwanU/+32veP9gPn2jpY6PFk9M/0gmj0oZLc0ZoePDdE2vvYgcXBCwb3RwsOBYjuWM6D8EO7cE
9FAYrxDNlzG5Opf2iVOdA/rwRoNQXM8s1teY3axCTJaAjuYW/SgtSU/SCLa4ig8+EfJO5hIow56e
8JJwSukuHAF40IDJcGRPhBhWLnCcNeaUQAECmVtNajHdrEaiusp6TH47LjM/7atT7r+PQPuYvFBl
fqnt4QlC/wzmeWaDXp87shfZYGXsZtL9yji37NxyyFEugq71oXmck5MtM8eLTb55fNxCi0A/WykA
zamWrVW2d+dwuu1AFcArFsKP0Fjg/yzaCoVx4mOEOI21wITkDcTD/Dw5wxP8z8XhV5avZ8Skxxzo
bVL2lZxppWbU69lzgT+a2t82DXaY24sjCky8xaLjaevwaDj3pxAMQBgD8zJVU8SEwW+zVRjbWOLQ
pKjtUhbeZ41C8oE7gMyh9REbosBsyMFpjgP7g2NPaHLkBmqHF8Jo5lzLNa9CNCrVsNn3RW3cZKFv
c7HShksEAvttHkBYr2WXwy7AvpVCTsf0wOtpfZNfX2b0VqYTo+hSYXMt4ghnbYSvAhMpaZsvdEKY
NIx0Ai59h6r6MS45WRaLnmHd7P+xUdX+hKW7WAB+NF0jIDu50+/VxX5i6yiyZqBqPYYANjbXTfIy
OChdOdeHgXMc9/evf6qvUfmCuj+dfElWr2zmP2tRkozA/nHUahU5t5ReKPTy6nEJCQC6Lc6wJwjb
3MZXlf3FGSTcx1J+qppGkSsQTdSiuTDLMARuI20VDdq0DwvL8giF2h7ddJiuZiZQp1KZ8H4LSw39
24Uhhp/ok591/Jsrm9vCU+IuPsYuqhtFFcC3tYR12lFf2rlVTccWWd4s6pil4uQtPxn6sHau3UZK
ZwOEqJrHEDeLhrqQbJVMBoU+6NEDJvPZVz3Zsq9tycVPg7M+LpDdVtrMXlPXdptFdjCLL8U2EbNh
95T2Lcu9RfLp9th6UOUDKJ1TFF3Fs/E2nxhiJahULd4l4h9iBgu+seMlrXCZ70pbOlEp/izwWB0k
Rl+cpy6pP2afABJ25k2cz4I/pBOjOheIQqwLL5GconiDgB9a1MS6m1MrDgEP8v25AECN3UkCOOd8
kZOIFzDnCY3hw5Tfg0DZASu7IL7cZYI5ujjO7y19TSXFc2gB3J8Tn9Q0T5l8BOWJeLF9dBQ+jHJF
zTvW3n/MCYPvjDkDKpkmcdZ0EH4wXlgDfDkhg4Kfdkbt8MJwVHTYOdYPe5cpRGnZS+E0ECspgNut
Fi+U8qM9EjJzEz5inmETy9jH1inRx21MBZrefLIVX778qqZoWQXWVqC3EAckhsFn7ZT41Jf13WHL
z9EA40/qPVrqrcl2iNuueRpIUjtNuu2DXRZ/P00Si53V/nFJ7I7LiDw8COphmSV403nP0O2H+taK
faEVUDZnaYkhEk63L+aPSj1d3rfY2S5IIwy7IxFC17icm8tbcSXRnCN+reeEhVPkYDJILvV0uZDt
UNhsWw7FRJuWDWy6KROfVKhwz9Jci/i++N4ebUa4UCuB4Mwcsnsa25bkt5kdyG5iE2czfVZdBZrn
Sa2Z8I+Yor8ncwVONOsCqx4m75SQtnKe/OpeGKWjjlOgBMHqXosjch9pnjNQ448Em8xaw1S4gUWz
n5BnYpR8a7YblKy4n1JVBNBfbTUmCGUhXJsT8Jar5fWuHmKaz3Fj6EjoP/LgSE8oCEWNrqoET6OL
pPlt7zN3WfhtYpurxCzWvzqSy2s2EW6UVE18lLb9f9ePeVm5IBaCI6OZW/d2AmaSIHow9oU4INPw
78ZAAO2uNKCj/qb4dQ//hbvedmS4gf3Gdu6iTQR/OrhyKPkyRDVrCpg/hT7+NkrW8R9nB3Cu9QOt
WXnJimFb3cQASM7/e0te/ipWFlCWIcef1tBrs4dW7rNhAMLGKVTYsxH6ArisLTTqMaIpOn2pZyZM
DVAaOuU68+GORWZQcK4MNKL8fNkudBTZKJesyfE9q5prk7Mge6ZWluRipTmyrBoF2Bi06vSD2MhT
36AbFV9Dr3cEVZDauHRRu8eyiXf9tb0izK0myAwbPIjvwlOoAhLvYBAP2S5lJ7hqci+kpLqaPavm
Ty1TcBycWvQrr0GX4Z3auWLzLPADBWwEeQzBlPDcdhClc2VYGySIbLQwKS8CBn2FXPnjLWQpOPlg
Acl5XfGMZEjnJgB909Gebv7fCz7Mhh6Yk7YktnCsTomJ4+NynAaAPLe0WNzkzW7NB0w2+0Q2JRWv
KzJnJQtDKIY9wwOAlZct8f0UVeQKaozcBXs2fmvox3gZ09laf8r+fJP+97DXcTi3+rGimlEBPohG
RsiBmKjn7LUP4TZl6c41nRPHigTCuek4GgT87YaZD5AzKo2LHqaaPeJ3xVs2UxcqVbbwNyCFMdK5
ZpoYbmyorOUrYOCrerO9sVH2w2OOrmSBGlFhJtzb1JFvs1NzNi5N3EkhF/c/1VxEteY3zWt6D1Ua
TkiOLNaW4jL4wPVt5QW2eMb6p4BoqkwR9L70dX07zdQF3sikVBwgXpzhWXjQ/NJvQJACBF+Q+T0D
4WtRdR28OeXsSS0n2fjpQB2vgF8B6O1bnCk1z1Iaj5yqObXSe25rJlIYw9u4ML8i3NxELSbXcmm+
0JNWzaxypdtwHwCJJya0sYJ7mti3pfWxSmiOtQN6LUu9z/zAGDmxP0CLOGq9Sd8tAq6JOqcwq8sb
feGyr+Z5Gp/B/9z99BdrigA3WiyXKoytmhPveuo2xNaaQUcTbBeFxk5fmZ7mmQzoJAFrNZOg/W9T
qpCu5exPWfOPt9QGbgTWMZCQtka0koa0GgbfWBQWo9U13hpQC0GY5X79BA88JgQUI6+BxI14hGzO
cCNU+/MB/ZJde/+r8ugQ+aufRhOvd4A2xgJTT3+SkTQLO5TjOmcJoox4eXBRNhUqPL6C4Ir7WmXo
bgcG0IgcXOHilD12uuasG86B/4Z7xfs54a2pJtjFCgqwyuPYZHGO+d+z3ICYz9VWfRZTKW/wYs79
r7nsmcM+Ntj7AKNbpi1/RmdxxPxfNnW273Q3J1xcSN+57Bpie5iV4pRXi9slkex73NWNuOos9Zwg
K1mVpbfraTno6DudsgkYBZxMlS4pGjGZPVlD0IIzm8qzc+DYy0vVoZ0Udeaa4VNijg1dVbIyyNLj
NKZCr+EF1R0U5AXtub/L2WkWZIIeEljy6fvDoaGOBgGpAPO6yszZeNtRvy8121FS6TQ0YUPDPFIv
8FEi+4dDw7gdCIRnsJ7L+XBN0tYwnWkZePS4hVDVAa4MAxog3vh5KBjJ1VDIk+hX6v2ZVPwAeaS7
uPOUFcq4H88hz3cPEXPZXaWNYcXnbdIkry4ezlSvij7quurCOCEL5CWU/AssCb3L4I0m3ALuLQQI
aBA3GObcnfBWgWTqn/FK3SqwBZM2CoEVBK0OD+lD3XqXm/1/BD8uVThzWUnETBSqX6QgxTQlpLqP
Ch47D5W3F4Q9wDgWyyd3xLOCF5jXZWH0dgKCjzgc23o9g2g6GT/Vm/vOMXcrVBQItGdEBtWq3Zt5
sVjA2zm8quLIzpb7X4j8W3w73AdWyLqyssxchX2q8oxvycEP3a92vKcF4dQ+qnQnnsA29mdRZMhV
a/rilIByZatIfcb26DPCZUVriiQOnFJQ1BmI6ZvH2Cgwih0TgUDDK01YLcL9UQlPMYe/kTdsAeeJ
JC8gVhuh19ycPJLoP6DEPTHXLjQBrd92eP1qObf+uDJvZi2XeHvjruRycfrRsn0/bfM/I7gphvp2
9YcYwC4h8fmRhPKjyofYTCjeHMldWj0J28457N848AI13RpRgqR9TxnwkChSp7Zo6m7B9VQqt5yK
I7vLc4ABYevAmE4XiBl7SDON4m7XNz7wwyZAJATl2O6O8OR7NKQflY7IegARKgMDTyMx2uwdxgAd
YFmSTs9dgiDw4vOKMPy7/6TH7RKse0Hdv3VEXS7uji9qZkotOB8fZzTl582eCnot+HBnN7kScWKZ
UTspdMdS6X1GmDvcQL/kSGStIcpLxq98fc8lb9HPS3+A2gaJlqV2or+ViIoQxro2oQau2uImKFaf
POyMJezEPlXxtsokf/lWv93W7YReu75lWYxRoXj76c4dGHCb3xQQDCq5UYt477QdAvm/enmhBCfx
339L58dKXsavdYRah/sNOIOc04aCtT1HVxI13Few6m6gi0tgr8LJvmpoM1BL4UJcS780Q+tGpoul
05txBliXJIl5XdI3Rgc21ZucEy9AjcGZUmInfffaRhDsF2uacT6klMKJ8zuUoIkli5PbNWkeZNUH
edOtoD1EOsaVOygfR3ynZv4yAZIPmdrUGXiavYlSmEzVGB0IwGk15fyhoX7uV8vXPoRt5dosneER
TRLBD3t/nMVnZ5lPPHAlJVLvIV+io19V27nLzfbC1rMcexYVqGPPEBInFSd9pmrPPV3hcYc2/qKN
zl4MtvImszYVZNSDaiUSv1bUbFQRzOGI36yvnIqeK7S/Kwc6vuWn23wctL4+t4y6mBTXl6Lr/3Ii
Hh7BnAYsaXy4QaC9c/x1JSteztEOkfwgGQfekk7Qpm/LfawukWnVGhpeAlRPE0sm9Q0uFmtXQRTT
nTAd3SmIqce1JE/WlDuawWLUMLAcFO520T9Ge60XgaLMd0Ft+FWsvYFl2dXpA+chHZUf3rFEUvYg
lnte2FIX57odskQ9bNVVhxcKOnTqGeo8f0fw8VXm8pDaJaFrk0jk5ujyq5p/ezAjxoTm5JtOxZ5Z
qoJDPdzmnN7BNmz1T/fmbWZTJ1KLxdB39kujV0/QvjD3J8Fro6RdsRL+o12XL7fY4Uqc3aMwuoJ/
A8tW9/BeqvJNesdlndFHimwlLboVtRk25en5tW4/bELCJfd3a8iJIDvdESOxj7cGJeYlwk9E4YyD
n2WRqMwnSzk+tmVC+IZm4ASY0CSly2mzY64FFUmoojlFO/wVVXBHoru4dg5YGkK/cf5UcCwwdGvx
q/2TXtVVVswWRtMMAKBFsf/fVETLevbb0jCNLAvEdBWfYyOeViRbtGj12v4AtpX9TOo2IhwT0DwK
xYIPe8eU3c/n16MhEMsSzmDWBv+tyGzWRZVpTODh0k37EQvHu4bVkwVbNppT9hBuLXw1iPh98aCr
rCOOwbND4mc4N2vm0F0Jd5bS1r11QBEa8M6/waMG7VaFPSTXxyvABJhZ5+Fkhq97rOh/dJ9ncmW5
2arIAfl0/c/6g1JyHobA3Ssn8T9lyk+a/CStcIi1LEXDDfXOrSG8qkgCrp3Kr/9hOFvs9cHwOisH
vxsJc3bfDCB1ragmHMKFKNOWJA6HEvTJRp/KsOegnStPXpefl1WjagY41ktr5KjmpgAGvCniOwVU
TUYREi0XAn8Hd3VElc5mEkqkaQJRbKwUIoTZ5Ztl+NkMBS1CTEP1CfzAhX1PRLjmAvB40PEdzWT7
nlsZyDvDgSmuwJRhZlsBRds8SkOIRDjLL0XLfrhxH/FT50I6R6S070d/ZEyu7rdII7qtbBs83s9P
MN/KwHqtdaNuWeyWehPF6Xsv4fr8bqKsLwjC6XTQKWcjXHcd2IKYf03ePHGtDO2h/cGfWHouuJHY
onN0f3yxTfEC5i9UhoqmGU3ExaTmULBBkeZ0c72xoYTUZJM/SUJ+kJVnKJZKp+WXHLfT8Mx6XQfZ
oBQWFUnwNiQwXZRi3eGMjkGTML0dFHuisGcll/X5des67AhyTj6AgkdLGNkwBdVUxYsjye01TiYv
x9RomswirTCbrPszmYFM3USL39lwkr/ZQtSGtVYssfY+/yNS0sqpvn2Xgl5NmOBooHDMuOx0e8Ol
3ZIIfq53RmemL+iVv9L+ik/pS0l+UXWKWCj6Sz6ArYaM8cw70FEc2ligIjx1eIHNzRrIXESDvzQT
5hhGgOzjJhiFVtv4OVnRKlsnW9f+cGLy3QNnQZO02V51pfSOW4tMHxTMvv+OtUVQ8sEqPbDMoxod
jcq3pQYbzvxcWeYr/lG5YXUKjusXcBsoaiUrdMsq+mNZwRidA+ajGvlXLLgjZzsgGL7sthRjaCIc
JNgyux0v+zVolfLXGsXNgyJdTHFeBHfpxLO1Xwb2smoTd++z7EAoLCYNLx1x9RmwD9lvFD2azUEr
jih+CjQC2lU1ivKvnYa4z9DFlDhbjUKsktN32/5qkWA4EBXLPhS0LXBK6JsOFtEzZii2rL86J+l4
sxamPLG4gqgh4ckesoVu3lljPskmITcZK1stO86b6KSN8Fsg5X9dvl1EammOnf6F1iCIHtL/3tPH
0JWbMJ8WjBxcwreJoXC3zxK3tw9xWYnvkn1Ergf+zo7sBUSFVnW6AhHlRwrG7nCvFdcvZ17fFP8O
3uc3XACgxJ0nUz9WSEUr0YX9Kt7JkXpdOWy8UzAKC6KLM7/Zb0yGEBQf8Gr+q+rH7rkuEUwVekJd
KqTiE55cd+W3KvPArz8y9MtsCs/tx5VdIgJv32sg8kEHIXxHg4mFqNRecb225qxEFS1w/bkq8gQF
0oiG5FiA3cJpn6nMux6kldSpjiKGHwsSqPbCb8d18X1OqWknulee7j3DW4uGncQBQ5QrJ0nxCxAl
vldlAg7cIS7AQRwqd1kv2FTnLy9EVeYZz1Eq9X/dLcSsLxOxoIyHmuXMg6544SO1jd0DDU7gjLA1
GpACBDf3ClLovLBuZcpxsB71UNUxo3q83xE/WWJPAGkXDv9jq1TTkLp/Sb9/IqTUa6PPEl5hmwZl
IUSnFLaa+3/eN0SWcKWEgG09Hd5m/AlxfU6N31qzEmoqk/RjcICrYzwdr4NHYEj1ladI0HuWXocL
ysExhsJOGy7+5Zy+8/qdwJQ4+rnKT1NwyJo4LLrWg4jt1MN6I9NXy+iXkTNk838m9bzhNL3wajnC
Bgj80MJe4ynQeSq/Sk/0j4lFHWlt1ygeM5y1GXN9I3A6xxasBxoPAmujThgQkigkKqq2JadjXAql
+2jkmAFf6lGCCtH1if3syyRLwlbzW5M1qqVSJpbiGH5KDrCCQs7/Vv4XT0VV7R7f+phHqk07JoGz
AZ0Wc6vtQe896xUGVCVYgAj2Nd5EglN7erOrXK0m0N0tHkIx/jn2Fgd4f++bR2c9kOURLe7LjGab
TWjTWHJnabT6iRGXOnPC6SMj/MWqoOPPrWd7OP6lORROSF0iL01iSCl9HTEL+Xqfnio82LJREnRQ
WTXdNJOP92oQHCuGzmwI6D8/Rm++/iv8nvnjGQ4NoqluBeU9OJDjaawafmZOnXSouzdBt++tqh67
uadS78K4B7brEWQhLfTp6snpPwMTeh57TS0cFLfM1i+12V79M+cx2X2a49ezrpzdf3KcdEDiWmXS
KKVtzs2egNsVmC0w4DDWAMrhCX+5ZCSrodU5Rd4cAqvUI0Px+jmTnQbyl7K8oiS7box+2r5V07iT
8TYLSHuwRiWesZmkOoZa8rxr1GVFDuaYiEW+eOPZS8YPx273PeEc/A5uRDt5jONfaFBSH+s2CJGm
ZvNGtogXF/EnLsmTomkPHDklCCS0mBTQEcNHuNFFTRsfb1wDr06LNUnOYaNycPRdll70tiNAP0b4
0IccOGS4HRLwl5Jr4GXdSq8wEEOf3oPSnbu/7fTwhvPF51JoeZCkHShWBYS7Jm10pjmT9P3VIYPF
1FUheUaLhkz9Y/rxP5e1brlR/pgNpDmm0n+kutTzkUnyUuhOH68uKZ0Y3G1SwIvTwjoHOnmLZoyo
d1Cr+s5yIf3I8C8KZV2GGQ4Z00ObTE+VmcuGpM7dAcpBeocteWJWG5BcAtyP9+nfP5z5Hk/+UxTM
T4YQFHRE0G1CuIk172mEbIFpp/LhjjFuTmM9QgZ3Rjw8U8/P0sPbcyesFXPy+olQq/WIphxoBW+G
Fdj/u1CJQ0x9ftRazud4qmKfj7jxJyPpLtw2JTQdHTcAtyu0npq8Fd3DbKEL2dI4e2TXVDtSPZay
fYPrZvjsWKufVBypj4MmRIZKJXz+veFfWyqXIUVORSI2IPZi6hKRajht63+otN9lXD+dx3kTQCC9
nFhhwtvaM4e4ueju+xGv1wXeBxk9B16FVu/gbLvKAcShWhPJk+IqQ37CJtLku52t+ZKoki/TQa3q
d261ZRAEb2ikJa4E44q9BRK6oE0HXamWHeqSwMMifTVmlP+tS7fjjJNE22yYY45P+h+dMP916PTN
TyC/HY+hTxXSnZlQ51Uv8c19M0EZGEOKiii7ACBzy4eTEYLYlqrGddeSZTG+8Onj9QliJ6TaM4ff
HOfC8mMvQoH+Dze7hLeSbhio2AnuSY2tr9Wf/kXchZlwjAXziTlgTq893ojtrwxzNs9RMqz0gL13
wqkxg/mkSfbOra5Ff1dlBAOrArQ91dOIkYfSC/dYCazyXFkXw5R4rT/o/y5Zvu5DKMF9YFXrnGY1
mxBSGDCqgKVO+GXGSrfevzguKgBAfUvxOoaNkwyjFf4QWf0X1/zh2r7GbTtsY19ukC+rylGdrGNV
7KoIxapXHqoX//ygLDAeb9LVYr3Y2L4BSqw0AZ5RwtBTb1VzaK9VFJs9euhSSETFeP5dmqodmkT2
VB1rdrziHSp3EiqFRMHAyVTxKCrlH8dLLLUeLEC+f4Gzf+BIzP0BtUKkal+oMDAPUWrUr5zO/WIi
NE2toLHhDpWp9cpomQfzpQhaz/sHOcIjywzFHhQp15JxiJ4DrxEpC6mJNySyJcLvTT/2GMuuKgA6
cSuWudYM/BPnDUzmrqRZMgtxRwFNlMSA/d4Qo4F5tcRJ90lSYAOXwdeYbg3XOBFkxZAvF2Me5hY5
4gb9nmGuhG6WqM52yDOsdNE+pYiu/KWMZePwRV0XM5Givl0y3xJDkPb5fhk1P8oMCr06wg1bfzf4
+PQC19gx44LVANQMtj4NLnvs+dnYRk8AzqErrlbGk47AP2/Pm23xD2Zfcdzje+JAsbt8p1kOXaaK
WcIkQYJQv4uqNOSWU4edMj60qTDKrld7+oNt+wZIsiu+zlN1WhqOQlKgRwgeV/ahPOVpfvZYlX/S
dhUzv5R4bC0Br1I6GPPegF4vupVHkjIPEgePmmYBqtY9Pi7+/wigbXfO2svxe/Y56Ow/FMBNKurI
8aqcmhoKbWpvHdx/iTtCOp2A22quGfs7qZAtRxhC7TSYY013+gqnzGZVwWWCZn2NlinkX+7Fi/72
jcTm7fIwb4qNkQCcn98i6NGq/wH5Po7qdYe0KJ0jG/clVmy2FxutuEDbIuJEYzYMxm94cSkg/ISR
EZeSLDUwwW/Wx0onTZXtP5RNztyvWHY7nKJ+7Wak8zVC3lG+GpwpIrNKNUbW1q3/h7AOoDz3qmqX
3wJ2cOeYpDlMyN1/tqxLstw8j0/zBzEC0fVL83/zBDURBwb5YBgI4K8DQur/YvryNn0lrfDTwS9V
ky7U5g2OofeLmASOQrEEk+K8KVgxXTjaV+liZT+p4NrpxjjGVk6qVRQubb6fxp51x/Igvb967Nnv
H5YBMaE1QFNEeVAIhRXsTokS2FoZmBQkdCzHq9gvRUmVzEoJ9N+qf/pUiB32P2Gf6XJpt4GPP6w7
Bahx0H+83kMksLzQlX0Tw4HMZ4WDUY6X5tJG9dFsWM07Seeihn4Ue8BJ3f1L5UrF9k6lAsNwP4y5
cZTqSOt5PB8PlzT+pSRXkc6Q7+YdkWHASyOax/XO0uJvAWL7ISQhZ9B3JqObwZA6eINdi7DNQgSC
lt/AF3qTKe3xgXzZl1XtQKucaVcx0L7Cs3dy/HadlaxykR/Xs1Z/e7ehvhvFbBfPRVmLAvavRQ6h
fguNyCDfMMc27nlLq7rMIINK39nHqkVEVfh9pjyhg8D6y0gkalLdq9DZftoXFtpVMWfjWiRneWOQ
dzXeAClqysIpYSfgg6OaW6tXiNDcNsg9SDBxhYfQEL2lirJPgZ8/doobfZVmu0zYIoIqXmxkjshL
twijz6JHAmMmorhSLm+yK0uJh+m7mwVeTT4LrWVWm4CDogcUwsjQoae13xkCeXTLPU7Hu2k0Zjpf
BBygqtdJz/yc8fhzgNmkstrjVfQ1hjlLqIEy+gUSSKCWXxKKSnoDHU67NK6tnQMiekYDKNA7mtsf
Wz4ypVlnP0T8JjmPHGrMbRo9XLUVbovYMFJ8pZDLh1A4wV2WjBpXs0aNmrtl59z78aF0az0G+SYu
7g3D5c9sdK6rThW7/DjU6RNwn5sJ+aInHWtmXvlg8bP667/7uaRWFr4uAlC5Bh+2Rh4GvrAzGPqh
stlhkSaaTXNczjVsanu2yHL1Q4glJwW7+uE5VyGr+J42MHIq9CoZJQUyhcEmHSGcfr7Sml1XZzs4
Co74J0bkg/awXz2tq42dmXPhDennTtUsnxJm2ar9ell3gzIl37Y2iVdIvvFOqtdyB4d3GE9CEMTg
MmCjA6FJ6Eq3UiZfFZUamr5bJXptj93nwyh+HBqJhPQBu9u2oYmqwMxYy8l4sagJkm4sLMdvyako
4b5G17QAOY/RdIIOcz2MwrLs/ItAH4RfuYTjEJ7xdrae3Je7doGPJRCbyNp4s/DXqjuiFv83gc6F
tEhKhZA6SG9FWVDeb7vabCvKluXma1BBysGn4M4vKpDFLwij0SUDSBP9okgzpUSDOTPFcRm9N4q9
p/YlnaTqmPQ7wJubyfnwbAS59AtVHskk+m/IfwlxgCZT8Fs3e6bbowlqekDvkpXtCN7XLi5JPjU6
rQ8M09fWywsVbhvmWiulyZyXyv4o6yDOuGbpiZuiKo+awz3P+B03xNSLxQ89toKuZDBuzhyKQvOh
gSMEFkzREZsDDr0qUBCT2JkpQyhkKu/RHdqOcMRruXk94HUdYtuQChokRor9Q9vOrW38niLywj8K
6DqEXQALKk3btNZ+4kqekbVc1DdTG96Q+EgO2q4mwgul1vH6fd31pQ5TXfPGWG/xINVa+Bh9wNFc
cbUIhvLRFCy3qDt5QIViSSd5X4Mm8iL2Q9I7EQVO392wcYQ0bIntBq3/6IRdTap9VtHQ5RFEkPRp
zHpMJ73cQ3wZrxcvO8fqzn3SlctuNgAhG9bI7xJZZ+Rd3F7zpS+ixgIBTGO9WwBGbljrlQDlQOeg
HoWz1GJFjJ5ueSZjD8yoEGP19bV4jNZsktw+ze4WMzkbB2hgasu1Ztxtz0RYv4h8WXdPS0B0PMYt
NaS4fWXQZuS7gvSGAr1bpex8HukAlwyoXg==
`pragma protect end_protected
