// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
tY3/n7Ph1Ym06b3M9qFfG8AU9xvJ1J/jWV8TtH6qQa27ITFC1BVSoM9QFs2m9UTj
jkToxrABC5hTL8yBFucHs7wA5bwbSgPlD/7TVYCOWvApWAvqyn/QtGD5LOkXG4UH
gyv4WJoP8wqV15HCA82HUIRhk9JhYiR2gDvHoDCbvkc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 59792 )
`pragma protect data_block
BhRH6iC6G8lrmpV37SO3QiBZQWhOttCwXKcSE81V8qd0tr24HZZIm3GlIQR6n6RV
K1rfy7Mp4GQJ35e8woFj1WXyOyS62DcbLlhLJU4QSX5XsE9NCGY55DCcR+Gbi17G
VkPFU2EAps1ERg8dw/rG4Q2A2Rtt8uAo/X/+LMxOyzjxHrTZ8ZyZa9pdbKSiPjYI
mmoaGQtPGVXSlAX4SUWZlD+iI8J60kcLQSIQo5Gd0M0A85ooEwnuuACllMVNi6zT
pds6AGAksOumyWuBAGfrQV82vrk/hNv+ZcVl5dBApglvTTEz7bQozwm1ns9sO5Yx
Kryd1E+Dv1nGO2Kmi3hpWwwiZ/YDfDWaPcKv8hpTXqkUYDGJXzmjYtJDgaT+vfef
GRPkEADSSdUI/yLK1ioHdDt9fCeIqkqRQS4vDWQj99zyyZBratdABN+PuOV6rZv5
Sw674EjvAb3PslgH4DiP6xkHFAf7tElgTEQqeCq/m1cIrrxdIOLbR+J+Xl4TYQQi
U2c/TR+WlMnk8M6pVWmlH4EX3ISUQG+3GuUYiZ8aFmLSJOGxlhVt+SqcIxnS0ooM
dZHmAGfV+/NvfsgyokiedS4HtKn1rHSgMjacs2cePJw7xfCBuqsf6+1JmoTPO99Y
4JEJoqTlwrucQpAob7YkyZq+4E0q3n3ahH0El/M/OgVHSCLKAnjYyizKf0Lqv4vG
MlZOvIqmpoorAboHQNPaRXP01CDAT3h0VFasrwqx2CybhhK6SnSrdcPKKv3k/avE
unHkbmHbDRXxBSuQuOf6xMGCWg6Y9RLEAtfUO6eABP3htgxqYuJwhTACIyj3pQ0/
aFWsGiiEW9/5oOstQq1iR3tRDYzaAtZfZjL2KkikQCjvJqFxyBL0J0CJbTgswXL3
Y8jfiTBy6PAX18M7aMLhfNb55ENTU6xOnszxB5f/ppdfzhl+ZsU8bOB27nmBUQEs
FozIrFgQzrhH2xXAfCI9SPmL8HA1qh50eq3T+SJd99FL32a5jWrpPInS5ti6W1mL
dwkeDRBXercb9r9NyGQzc2/6TAfSPx97KEPkr1MbmkkUuclIEH+j+HGe4ilHGH7W
BDsCQqXTtXVx/k2YBvPPO4m67okGqYAh4PEs+1Ed45HMusRMThY+u+dQdMLPC7Zh
tce5cmRVaM6rB7iSDm7mtfk578gIt9+vmPYoiaDxDi9YN3aWs5TLxy1TMa6Wak8m
aPIDXrWcTwho8TbjbyYP+vpOxgEaQK8gJNSWluv2SXHJb0zdwHtOyh7FeqTkE2Wp
cqrzEyAfSIgCLoDz/Kfp+0XUAoVCZcWXypT5SDxqeoPpJx6HXfzMiSUf2GE+csN1
Vajts6M99Cq+J2HZ5CIeCFvAgmg0doRKisXLkl9WXXHMNaLN5c+g6i+PqUaROUaz
eDMaU9k3Qd4vyOuYwTgxA2dFRgvktpz/r2FLZFY7ntja3aTBJPuGcdH3deoRcP7b
Nb2nuybW1dfMydKkyyUbsbciZa3r+AQtfNCosbc9j6R8vEff6tqhBdSeLT5kWm7Y
QRdjpiCYopGlWY0/IQRIiPb9LEwbXkEWppDWzGAjY2acm/y0yPusb0EMK3ZVOc55
KLe2KwoV6ohwiAlXNzUKsWRlhHeKR8y68nNCJJOOiMZC9BN3ktK9QoZmEMYmbtC2
E9eXO+HfaI/GyuhwIfcwIFauDwbH2/oHrK1zBa/eRTD7uMx26EcffWXo5Xn0Nfb+
3drFZCYcbDFjVkxcdPDV7BnFMKDJcPyUOCuoWAysRRwdUl0x1WrJAChTSUIevult
EBTELkEFMz0HF4jZ5bphyVRPbXXWsOqQ2/MA83gWTPMj3iStz9VSLgWG4auAe3gD
V/mDAHYz4zIdz8BkUNShLLHn78fCwJnTGPONoTwT9w/BbFj7IRX+oCPL/VZBQEju
WSlx3iV2IyelTJqotwoEQvKMg3Dxk+qM9b1/Y8+9AhpjGSaXnKrE+CQ/4a3fMcvj
HwAleLOV/RTlYmpoxUL6jT63Pz7fmO7KEhKyeTw2O2BEjLAKqG8ki7x46pAb8Vlv
F/EAkXakqfsQdaYfk03fJbXQqRQ0Uifw6wc2yQYqPAJ1ctbc1f4jWgfrFoZ6TL4/
7UTyGG3MK7jhhu4m8uWXEt+2SL4UiAChXl4uqaxJn5LxQFx3pv1+x+Mkzu2L+k7K
nQcGR21jwbpRfeHaXn4NFmdRStYTFuWyAX2T/ax3sTie+OZiR2CJ1h12Yezxe0ND
85/V3CehHpCB//mDXy2x+/Uuiu/mOri7h7H8pcV5N0AtIfwHNjmtjKkPmuIi4TCl
nyBi6lcrjipVeSXJVwVU5zgucVe7tj6ACvsgLjI2jZFsb3TEgZxpx+UUUsHhsIi1
nx3cDif4ISI4ZaOpD5H45OMOL3BSlleTD6HbGe6CAcCPgSm5mjmLVgnfAZOcnUGF
8KokNA/Xk5SIT7Arla0wrI/AJw4k2NjRaV/XeAFqGqMpcIHDnqmYywgua1bkCrFa
LglIIqomP8N/BNg03sRe8v5j155LFr9bgTXgyh8k4dZ8tS9cCzz9D6Jn76QWwqgF
wJysQwjIS7PzDSCBLBI/JgueWo5Q1UAY/z3iWtp/mycas5UGTom0PagQKF3kFhOm
6eUtZtbw5T+jHdb0Bn+e7j800Ev2WAjhhiFTNx3KBRitr5BeVCaQWtjDNeaEr0FB
SC0pFrg/WQKHs+vfPOKm2NvZLdiI/K1PpYlzjJ6aEoWM3IhER0kk1z6MPJjYJpaB
eVT7CBm4DGAqIwX2b5P3pf1UriWEVOB0IXszhxgAZV5ZoqMCJEewvno3csSySeEZ
NXa0Q8CBX6OV2AsY4GYnhCSFxUB5vhvX4rfEzHJjRNCEQJHyFJ306zmATvSzANdj
5sLhHNT3pNCCq6s9skogXMbIoQKNt7U38V24+ISlKjua1NumEme8Pr3xqi/0BOFl
lL40HhPLMGI8/Ht+vdBxVkVc4O+TVD0Y75foAsyAcudYrRkN+Q3e0LZO1U+pQTKf
FoqiXtVRoQSYpxeKe+ZijKEMjJWoSEXZ4sm+q/CE0kZUC2Tx4RhY1VeIaNbEsqGf
1gwWoc4w0XbhqotNTOqVEAgXOrUhPw2DipZoEq5emBhgskrKXeJjSO+85XMUtdio
zFsJe+ZJ2Ex0KIRU4KrQq6EHYnr5KmFFLttmV2ceiKjhGVQFDOeot0JuUVCV7gRt
WrcwYG+DHgMa2p2E16KdU+Elr66MVs631yTweA9dxIPZfIPc9QbhlA4FwxtG1eUr
K4U5ArQgB1VD54eRgCQopnrWLOrkAGe1lm6wjjjZYOCLd2pwM4k/adwHMjMrh6Yw
ldK3mgnIFQWrshrPzrYG6fNLVSfdVGdhO6mJzUURW3tZ30l5BHqlxeTBlJYfxzZY
SHPU59TBvvfH4pbXM0Mi8Evkz5x0xKsDcfl+7NCWCwW86VvxaL5e6fNLR21FBTvb
UaTQpJAChbVmyd4+IWCJaOeL5CdjR5REMcXxzRPuOLPimAJBrd5hYUQ1ZKiTzdhv
68YS1BLDemxDb+BUzBKQNgYghOySdXY/LKJ9TZlixa0i6hsssmag2BmT9Orpxbsy
ObKFEK3hL0IaDoK2pEB8kZT1mYd3DmywYK/oiVciHo/Xq724VKNJdORHuCjVirSk
AfVyLFTwYI2CmSXp7RXdSP8RjMibDzSX8sh4IkYGnzMQdKU3YO9xt6Rf8OsCvMPy
mMc3ZPpGQKUzm2rCDzioY1KuGxQbqqatRuklbn1BQRSZWB4MgumcdVVHd1bYOZPr
Us/s46sX/m3cSaoQ0JTMr7qC5vIw1CVjpbP5AfXyOpl9baJGXV7YUbF0Fm2l+7AO
JbrSwvhGbHWMsPpQCeXOUyuPQG9HeelNRUKSZb9GXDUHmZ2vrAYzG1lLsBhFVNDo
U67PKhTbB739rKkvNC325ocuceevx46nr6fczT8yq4nzxCBuRQyyNYjaKiK4mJVG
iUHQ7jEgQlVWm+t8kYYjX4Pu0pcLABO2XadNsrOqcmmD9ups2Xpr43W1kmp6hrRA
1pWBSGxKyv2guVKpTg13WFdi42CgQiTnQrkmTHR6d1S9Z1AhSHz0uScUpA6XcvVc
LMHXlwUWKLCufpMSS3gfyTgj44cTh1HAEX+a9Ys3XG2Ulnb89/dsOxryZLevXan6
4KUER66CQvLZFaVDcKnN1wYToLfdmI7NE+GpEUYe7dw59g+wiiiwmi/9MeISjJR6
9Y6t4L8p0AjT7jcbsfaMQ8J41GLJ39sRjoqBhMnhNDRFP4VsYvYkkCpWzamlKlsw
Jtc351K7eo//ooIaVo1x4i+YL2JVYnZRN7GIEsl3pxPFtmFT2VdOStNfIDeDAJHl
fO221szUDN0u+ZZ5DQ7VLjAiFCNQc131uiG2iS7QtQ31n1RtUE1jTGCAzkASk8/a
p1XmvclkqET98QlfI7OESiYng6pjqYZmXzjf91B9A6IAuGvRFMbKA2s6FgL8kI+I
oGpICPBMdn3wqAvDwJqNanVsDCxM7M2nPuBph+7Hyed6jsKT4HX1mYrrMFncdeWs
KFeouw+UC6VVBBRKngL8PtG3ZNmYYihQbfsjccPOfnu/3t+Vwv0hSgRSn6vT32j8
3Ty5PAqqWcJvgHkiZfDW7pt+lGnXNCM7kbuXEUfzqTYxt+N8HPZ2r2Md5P141Mue
lsTVFSnH13Xwf7g1Any0jUR2j9APbORYgZQTUD4vaNd6x5XztpLU+XG5Wt+Awwdj
sh2x2mJ/DxhTIRm83zhnxcAmQ2QQdvcdf0fpVwBYQ71cg7F4hnfDvwQPPxmRSt5I
MdiA0Y1AxtfxKr4rx2dxeJyW2w3gceyl+1DvJOAyfDE8Qf23wA0wNrAT7sFhv7yK
zEGGRlCQn1ymZ9+wHPYtPWQ5vP/WqBHi+tgEQ/APHG4XEKTby/iYaQ3WH5BFHSxs
18eA/erldD/aR1ggrOXVVLVmHphFssinm0KUOE75iO8PFdwkirWZKOrCPi359Cc7
SBpPnch0E1Pa/szfb3y7w3khR+17ZCEpP1IV6tTLdpLZdin5HLn+JyiNRV1VEDj9
7bx507t5uUpjvtBulmRbRaVA0wmsoMkRAbTZORnjp+Jy635MgGmWUfvI5q8NfQKp
DYjOrBIt+b5fIR8Xe60VXEpvduRKYrJZHrJ/CUIu8XZoYYhCrDQj3Y428N7T91yz
NFlqfccIV7p/3McQ7QZz6cUWp/yIc+W5gOqkWJNO7pM/M8J0GwSIigMOLBCpqx5C
b/0U9L3ROgacVopFUIGDMTLC7fwdr7UYeeP8udzvg4axQ0FiEnXWzA+sxdaxMx8U
pONIakxygC4sJ96Vav5pL+YZ+nZtG3anTyziVjd7xVdi92N2n7ozq4sgxSjo5hbD
JCmH5llg5TMrvZOO1sQQTQPvUEAsH4vt4hxMH9Pvy2Y4939OveolZsL4FXhuuw+t
9Hzl/NoIrnXFF7Hxy/w2YXovwoc3XmMGXtdCUHQ06Wq/4RBP4/7mEILo1YRws147
qKwjuAZFACiwNk+gOMmfz81J9sKuQaF8Kj+GrwSU0gE5UCiW236p0gBpQXQW0pYb
Zxbjsm3D0NYz/3sKIGQo1yzPkjPXc/Xq+Q5vaFlAp+ySvw6kZ6fDzTYgCQ9dzN24
RyDfK3d9rrGJ7oWA3LADKePweEf2COb3nLYccTaOcSA6FgI4Ilw94QlH2CgFhOjb
aR5HlTd6FU/qEROE2ZV1FKkFUyaOMYds3KEMNFSCfYExMrm1FrWPir8AEuIogzNN
MmS5nQe3+YWoeIKw2//9XeClfpKEttL0gl2XQm4niVZ9K4SAwFg6SYnxqfvz8hmT
/HKym9BVLZTcppw7nOP3B7Rz1ifv2zdvgX/FHv+EIyNIskl/6g5VafVtdr2+2m5n
OcmN4Kf6u9BR+9lU96GCSyuOcXXdG/sEpLo5kD6PfrOhB/WKEuBQkAPhmPgcW1CB
iNHsG9ItJBvonmwyT+IemREmhxT9y4h+L3y8TBy5mtKN/ndajeI+jgZsE5QjNX1C
kni8RKqKRqh3Re/6dNBBNzY0tE9wx7YEZPdCC7viv1+90E9xePV+9vmXHVehz2n+
g4rGiJx4AiHcOjtgefyxMvS90PHBnRFMZiesz4YkCNTYENI4c/xXTglMGtMn3A5H
RjxEQl05iH6qLM3LkwRDn/NuJKkOkqEraAy7OtWmH0/Ok8Kc7VSBv3oJQ+vLpVM+
zbMvuPJAk2OC2Jqeq+uczFYGeCSdxgIfLsFvbnLWboyijSWtpPoDwS0ji4xuTU/3
nU2UVB3ee0lLDOAdLyrjVIh1nDgBrV7vVkrRMOhrst7aXfETDbTkRl1c2pS8oUvV
sv79POKlI/EzjZF7Zk+rlvrup9lm91tvB4Z6ZZ3c4E1HwZlOfP1a3n0LyRws5HEg
lYSthI7vWnH97M3q/VXmuyhLN1xTPI1IIEJS9OgljIKm5yfcfSt1FJiETfO8gXr1
snK/z0NdDX3R+CV/UrwDzkXlbGchc+niQKUdEE7ZP3JeHIbQkI9Llll+5OlFXw+z
YqyY40kppz4wrImRjC16CZYoCP21DqOeItoJepAa36mDo265ytFEc37Aa+R5wesP
56S8Kl88/meoCbZ4kc3iWGKgt67CuO5KT6dG45a6RuD2TlRc158OZasIdklvc3Th
dhlJkUGFidczpxEKHx9JIFDtWmQk5+3B8FnH08bgl+Y4GWfRFDaQrOOG4Dr7BRu9
6K9a/JNEC2Z5f4cdm1DzWiN4OyatnIlXHipMiJEs04e8gpeNAPjUPph/JSaQLo/U
SbistIvnNqW8V7FeF9aJexPrQ6emczKbM7rd2ZtDndKxiZu9iNdrmCXECGGAa3+4
cIMfC+1tJ+UBbYMk/3DMSytLnxjnrcbMMNuAeKBp/s5IBnET/pzgjXAdDU8lg9aQ
oGOx94HyyDQ//w5UUK+yxjmXdEhDKX+WeaHOc8S9GI6kBJXPRnWbWxhLLIbF1/xF
uKIjMoSTNE6UZ6QI2yfjEMahUgm+b/2Z5nvM3VyVj/isVH2x6GMaZe/V0lGPLcZD
TjlvFhOGQERkSTn/r6W5ogoJH+GU4wV6lE4nVxLJWowYvSEFoDe/a3kpLKcBHz8S
ivx0JbQ6esj+memGWf8pWNDHtad2KcZPpfdnac6JmmArGbJIEdKoa3Oa8/fqNqxu
kDedE24YFpQ+iHoNtEEE08KPNTn7/xn1aQZA1fj0d4AvIs48khd51DCCUGkhj+vT
Ng1VzRquH1SYGlUoDVsdPzchb8DE+NlF57w2+XHx/bNcRbwqN1RFfo3Hb33BcVxy
uQC58uuUs7Gpipo2enALWYzDbXMn2fR8Mmx94Rug3i2/XKwKP4d42CfxwwNmOo//
SPQ9UQCMf77HVdI+AMg6Dh6GBCaUl8/FqR1bQrFPx52OCFmLkvhdjFoElUnY6f1b
OQoz2sEf8BBHcbA3qd1u7JedJdUZIutlUm4s2UJaGKzlze8yvBxTRV7K2CPLMY+U
N5wFaxnUlccHRYXeOnSueOF01EIbg3RGabiZ2h9DEVbn73YRVZA8N7MeIHnKJnuO
/bN7xobVHCdfRPtPBFaoMsVIZFCmZ5vvyDMHV1QHRR97QqHg8Yr0tuRVsihoPRRc
QVj5qhgs5/ZU+eod+95chTe6AQEft81YrD2RQ9rXQUghnf+2+BGCyybP38bk8Zcz
/mNLly1aCwPDi66n1CzsikFkYeniXPrEjtpDWX4dlf23Xy3VCUEq7OxZhrFh7ENE
Dme7V45Kpc4DG1h224HRhLA2iOJS2GxPGP0gWswdiBAoVqRvjVb/9M3aVCeVtWF9
wWONI41rS5pW7c3hOPS/XZTEk3KmISnhEqYh97dLpty8SzdrGv2RP2LwlbMBiT41
zM0ZOwLiuddM2K6yHgAt9HNlXE/zMcxsHkLsk31ofKF+AaBCDLt3d+Iq6DRfFsbC
DqFUvQzikKGmX8kKQ47sLNL9Gg5YNPugIphZsGeMSU/bmvK5u4S1OL/7MfSI8RgI
Jc28DpIyf3RP0IDK7rnMtLpFNEvDsFfxMzFGK853UsBveAQEdXn40EAC/3jrdXZ6
ICYJ8ZtKLI52iijc1n9pADkSf7gCWU8Q/ckAiHFFDgEHc3GZLyuZn+CCgsunP2Qa
MIqO2rYpcmMqxPyu0DHRKq5E5gTn6agfml0L3lqNFiGyFOKcnLn63cUsCdwyfB/W
fIpP6RQRmDLu9qfLjGu3rBOca2T9hTnOsDCSgWLU6MKNamV7iFesPKhFNoSUzYu0
JmqRArZMBOCtEi7j75ELpBbW4MBlFtB+80cRLsUylWGgAhg3mBTSbyltbTxUDY25
N7gojomhHeDpxBZuniLTON+6Prni2NTs4MRFrwS+l6M4ztACQWq2NGMoZA9Ngx5O
OUDijmRM0Lc5V83lhL/GeeGQnJZy/qayxHLippqYh57fPwXwkED1KHWdkxeTptRv
59HOgmyg+mOZx3tGefIKFthYZwbdJ0+hFS64ztmHBsPK7huuj6s1cQwBtVxoGXrE
+9+ZrJCkpTsw2Kg7+zlCpwMkFiKEZ94Pqu4aItvU/Oc+2zdbtHhbrkW9UYSgme+j
VvLzyNiz2VtW8vyvd2lHl5napIPaCtB3N4Tx2zlYHXOdA/xgJ3xDiLgdH8ONMg9x
uV/vQ3PYh/jEDmAKIlp6fNGh03rJ/7VKsb+ogo1tXZa/VR0bdbyLdnenSV9c4aa8
0ze0ab9/L+eur/DZG3EyKq2mMPXjSPNYNJx28zcwMTBU29Velvn4S3sW0lPkhtFu
xjMwANlg4E4lTOCdPo53E3VvYPN5mVyrolffVwJPvYStl9A/nfUPeE9RB8taNTld
wiRcmLZtKP0geFPzqDhneaXxCe8tKv+JRL6mB0MUf6DYxMuilW53Ucmnvq6vUApb
j3xb+xJrZENrvK4vkvK4biY99iHIl+VWbT/3g46I9m813ZMzcVf9x+IQoEztCGNk
fzAelpDGzWCNiCG3ObFw0HHQyApJevAsB649HgC58kPbDK+7mkUEy9lMIS4luxbD
ncMxX94diEoSAd9myAZmOHyUNol+q3dWG9fPXORc4qlE95/sN27rVkpV1Fj3v6ss
Gjvzw4AXfUOXikTBLw2ol46eNa+HY3X/tktYweGfSNYivbBzzA+LpGrkKbuKJ64Q
U7jPxvw+URHcIi8dvLb2imW+E0r0lFlnFDnwqypQCcGM/2bOVOp1yyS/AlkwAHGv
J6L2hK9v2vmuMWAjogC5B8tEZQnZoK+KPinerN39IhX2wFSf0cf9J8l5CYdcwEJF
klfz3gJ5JCBPtoHTszsgFtuhIIoK1JWDt721tFhtvAv/vVBdiC/hSurJvwxhAE7K
lePWNO2eZekit+whyNdEnLCVJRV+fOJ77y+iV3JN2I7Th9fOpwG6Gj68+wMFNb+q
19Ta2LHtEjOsfNl7aRfTNhUgJ6sM/j6gjRmB9O5dENDcgdJgSq3tWVAcQJ5SP22V
EoO7kNWzWLn7N3hQmPWCaPLsAVejq8WPoKVou5F2MzAC3CJwHJim/P/XMj+KHDAS
7XaLYon23hPaFidoaid5zVpfEspxb5gT9vMMHyO8qErksPtbjguk0PqRHp5fTbmC
h9HA6W9AEOo9w1DL43vghse8f2IAwT0B/HA5RDCPCkHTwHQTL9PJm639tic9kz3k
eHEHjmUgKTT9QlGYK2yc75Udxuf/NPNGPCYdt7NWBsQdtszJo6dnpdyo5mwkWi4N
ARdnTeePvnfP2gIy3G/xYuFCzW1NwVrydLKltH84MJcot8kbCGjh1yKfp2x27Y0I
dRBH984HHyDrdJcSjHqvZIZqTk0MyqXMMG4C9E7viLKft85OXkdOMtYC4eFwu84F
UiRtSp2bJ5M3h9W62DtcJwCC2d/S5iL7A4iEmjBKMw1OSqGS1DCNSclCfjZ5lIZ9
f9vf+IXd//8j9z33ec7FhQ6ezh20ER7a/jXNPsf0B4E6PMIIDMka+c1Y59GTyjK4
lMSjigm3ohgDOCP6AWGgaTcgD6jCS+ddafQyRqrMsY2Vw/f66K6dMgynPCEApGS/
gZfJAt+zlottQUhdUDtoPmw5SUovohSOqbruEBSPSbqP5SxYyEWrjzHYHkEDiZP3
6p/YmoJnG44b5b4cMuOYS0N8BszLPQb/dFa20HtG5CHhzBZoSwrRE2Kft6F6lqWm
0NQWs3c10MX3EexE7fggEDbIL0sw4EtpaD+q/cYINWTuSHZkxzBsqzTJLXojoplR
x3xvOlRZFlkFnHTYUH5TSxRbbplH8mRmvpsVLKQ40sKK/i8aIO/c+vLobPrqnA0S
rhU6N9OH/wIg123GGhnlDqPwqZWrvp160FCH9w4wYRExSeQNM983SIPklcf5hqyb
5DGKglPZ8U0dEe1QK2ektCW80aRYQPWkMcOYC5O2UuGcxpc7LDETlI4cPZUMIAnZ
tMuE4Nks1qSLTrPy0rF/PTQtJto//1ySw9imDXFQIxTRHjN5ZA85rqvzwnmQlW3m
auLO6ubTtxlEoc65XKsS9iV2Lt1bxL3vHkx6dSL7epDk7vd/CZfBSQz5QQ+Yxy17
JaRmfZefx0CGoVCxJ0qZL2oEtYr/D241bRfFHACugIaohKbmyQ2bNEY1re7k09c9
EAP60DuJ3VgF1G2MBrbMljBm9xAGtX5BJTiMcApWFiCZgDl8yo8p2mvUCZGIAfg3
RDFeyJHsf9TbshGNtmQnyBwHXnWY2ytuzMrQ0GLqtsf8Uwv6+GA26H/8OF3EZAmM
HfQAadjmyeP/odDtLW2xXNdVVUj0HAEs8d57KWLi4a0yggvqvKJnBSqGIjJ+ypHk
mUrayiW3w4wnwczkVLq8i5H0B9sQLrCIBDNbuzf4Q1LwIZq8cOqSi8YkeLF58WTp
lL3sDMOwmy0m8ER6nQGkxXbAdFFyNqDEjiqRJbeal5fKTz4gU6Jss8zQRqSQwJzg
Bh/Wxr1tmwS9V0emtUCENIZHuqd3kzbnLVNMpDav/klypTZQCkMoQoAZ1s6/aLSI
3kXAJZhei9cuzx6iVaXlVlBjzzdIBGJEv/zKvhosZt60EDXPgNcKJEKH70FgNv+I
udizv6OHNQDFZLbAaBgDe7c4phnyX/dDIpPCRXJf9WjoEVnW5Gecj7wRxAz5wWOx
9mm5v2NS37vijjiSIH+dDeig4bOBG0ecYHdgyR+HXVC0fpacpZ2mJ1FjUb6iJLVZ
wUimssUm2AB3uRjawV/CHBnmAn9rj5+8sAE4ockdvn74dbkKQ+/smrnPFjgzZxKj
6AVSTsPqfN/LqHdscoZ5SrIN0Cu9tyrf9eAFNX1nvO2rzVabcy5TGKOIZIaMBLVc
TqM14WXudV73+iQtPaX4SvvCJGV48LI0iDF/lW5hul0VMZ4StZ7lwzrvn4nxMYDe
J6Uyd/HOBsfmlSEipOo0k/2OiRtNUpZxow9eEtNgytvta3MKR08qu8ajqJ6PwsWT
9sXyEMbuA7M0YBzJdODslcVJnKKxaJ/4wbN7wGmPalrICVFbgYgkY1APER8oI4uh
D5KaNTg2maFwibmGRbSbwXF8uIrt/xU+Dg4/RNRwnW6KIAThR3iEqXBMRe1xtB3E
MQBxV/sAS+F5gQworsNjUthdbrR7tP8kMMGIt98NgW4zyMVuF/9FFUo8Ftd6P3et
Dxrn2GKrIASK4424wjkzS/dAFT5zU8VMRWJqFFfwmPEy9PJeGRvsuTgeI9FmzU69
Vrk7zCrWkj4mWC+vxoPo7OCDDJT7MVFIVe5MmUiRLaOJxS+6R4Csm+68xTilYokT
vuyfWBxKjguLbsv0AlkYP31ug2OwCOCmMnHBIPB8VC2wI28aB0QGnSSZ0JNYXIBj
TxBpitAu7v+2lqKc+XqSHNDa+jLxkv6zexvSazCA0gysZ1+pD2KSVndn8tcJM6E2
APDOceq1vr8LYWmJCzT3DmA0SBJKODvUgGt5BeqsaRSFL7j2bSPs+EPNyLN1cbvL
WdJHPMsAgK4s/K8YwvMDGiwZ3nRod03Fkyh0OWcCJhIL/+iocLojiRxbh9+oaX1+
08HVhMe08K2lfEByOmxcTYeH/vQYnp9btsK8ALO5aDsZjNq7Df+9/8a1AyjQdqx1
foy8bYyggf/l67zyTOGWcdoVZpRAH7jbxLeTSTjl4B+1xvnaqFRwWlEFL/C4a8eh
cN3FdfGMQ4nDFjckXlHNPsJK3UzqhzO2uWstmzu5QCYwESbamEesfAgMNdve1vOh
V5ScT45p9Vlwfb7XXjtT996uFp3KCUEAUaTPcL4mcBupkFcOZ1LnNnYk0+c0rjuL
FzLqSrcsvDkXKKY2ScDoPjRaKoFrSrVd0xLutDZ6vxrLC+hHTGiDPKDGDwfa0Rk9
wPMbAStI/vmbw+soCT9r1Zr3Ze/QCUb8aY9w/bczS+EC9ALvgvc55sOeVi+rFfJO
HckxUbRqxnzXrqz/XPK+ri1imgsfDNSJZLVWB/h0Kx3qv/JYLCYvW2XDzRZyEDfw
RcAxfdzqeT9H6D857yrGkmM1LWOylW80vdl6rjLzLQmrQGDHmg4Ji4JCBSsUd7tA
6JIQHJGrcKVcuObXtLcUQA6lZdSthx5Qg7N2FXnqvoxdIUPoUzcKCFZeLzzzHvqa
H06zrtItvJ1y2ST8eQShGacDAzOTjdwes02MOQ9j9DnLIPtQDapqmKWvwmFgLJbV
0T7KL+2yEtBg6Tl4bEIRpR5btTpgiaugECDXgj1oSyujUAlO6XddKpKzpb+nqctd
+w82esO9Epd1mY0wnKjR2hZFRuTpK1KWvvutzhDXK1UERuDZZQ2m7Yi5HniAPzDt
Oktk6+cV0VKSfdkcvaMSUV2Y/Pe2fVHoYdCeTcXcYynOR3QJFEY204tgQC3TGWf0
Tni0KoOu8tkvOSlNInNYyRoyqauXK9AEqcvlsk+1W7hZpcAGjqdRmwzz9gjeYmUw
GqvxcpYwSyJft4T1kfhZsYGNes6Ykr1zEy/H0jbV+6ilQGu4b77q0LT+RfeWQzpK
fjOIJscesRpPokFJ+zGMcVc7gp79qOxMC+TQf0iEwbGwSm9Rjy19KlLDdJSRiJw8
PxMNI6qkt/n47u1YNaMha4HpT3wYTEJOZxtxdy3Y5Ry/vlTsLUTk9H+L61ZRX9Y4
v6iNmQy1GGgsQnE/hau58yHcxZfSewRjEm4BjfAmQmelwc6cSnViuSb+0F7mGWG2
4cgXM+gGYTFJSWfSO3RDkcIpexfbbcmxgDH2xwCHGuqCcSk9iek1jLZeJm+ir1p9
rj9JpTKDoWhYjPHWOJyvaDGyqfMDWcm+ZjFLtMvOVgVm59cgjn/4oBsaETd3nyid
fkmb68yG+ipTfe3q4HLd2LXxkmTEA6WBRHq6fwl/tEtHqsVy2HpnvW14DY1X1Av3
9Ae8HfSjhY1ppXom6qU9OZS5qN3uclvd8VcWYg2Pvt65UyAFo3lstjB+tCdwFsSi
gJ4wgUSP1V9AkTFTA7S4dSN+/2UOKM16NygoH5ehMsIBRiSrNSXTR8I+JdGQ3Cya
Jbo9YtPxzK453pawcI0dCSCLKDDZwtzq5kLsGb2hpfikt+S8zW4G6KjwbMGzHRBe
VXejiPwd7Exe/GdbIAGYzsPElJFvj5Rybi2hZHWxdPzPAUZ5oHpZFtvtnVIU8Mbd
kNCji8FH3bQ0Po43GcLM6sj8ATChWqMopwSaoq9m9Xu7IFAUw6T9YW5GjCrQ370J
5FLhI1XuclK1R9D5aE0mkjk6Tkxw8c6olSHv47MjV7bgnKc5aGKUGWr8SHM09sOl
9mWUwJSZTkBwyAXE3VuphXBt0zQz3tqWw0clU5LAuHZbgDZcG+eyyl+gBElO0Ccp
1q8vQoRuAdL+pIPSbF7Fw3KRib+UmOGS+Swe+7iXtNIfoMjhZllSe+6cBYg6h2jH
fASHNZ3634irOR6ZvyKkX8gI6PimKkc3zWKJNU/DiTntBq7xbTed/Od3ujnM+M8K
P6XxySb8sZ1BJzhaRmYDRk7dHforhpdkZmcZUrCl78/Lk+kZkzIBW1xWDIQT3PyG
k+8AV91DBLBjGw7dATe1hewsu4S1ajpCSf3RibCHtByZ7VQeg4ROYvSeLo7HwAZ6
8KOpINP7yf/qvcLbr8/jxQGc9d+T6jiAqSwcKlY/v3I+PeMRyrJcGfcdGtASgfWb
J75GMb3fXnegRFiXxbMZUov/o2qMf9bGaqOJCb2Xg0WEFURHz5w2/lTzVT7wqSoD
NRNkWLJm9kA4laulf12LzeNN3faxQbw4EQpPGH3E0N92vQ6cVJxmsXiW2NvF7YwW
lV3V3bp5rM3av3XtnIK8ejf4xHCwE437i0t3ISEoCjVVA+jGFEa10MGk3BTGLxtN
HOhDd6tuNn76uEF+jaEF/AjRB6ZeZ2geiWx69h1Ihd6pQIPwKfSWckcS2fRK6DPX
hKRf0G7sjB5y886/jWijLhFg30x8+j/3GyDjiMrwSXMPwT9in0tNIq+pTIFK1On7
dk09z6l3wDqWT5bahpkUW9fo5+QRKemUBwYCh1LThHk8Ngyzv5/+VOlsJZ7NRjOE
ZpDMRTKtEnJIB/QZrDuATIbjZ1JWx7Fhj1ou2cHEdS681CHI9HQJuELoZ8ZVH2C9
ID1wXzQFFIueGED5sWGbTyT2ayRUi01Wcw+3HJt2rKgbPsZqnfXpWTlTT4+0OejK
4bGDNMXNfgQYwmFlELfDXLtkH2gQzDSIy+BSxyWxEsqShvHIY7/BgtKwNIhZknwL
ZYZ4kVL/goTSyTniNrAT95weePdMhIQykCUjcy+qK2fA/nkCli2y4twyfSJPBeGS
F1vAkbKlXf81mLQDQQcYkv6RNXt6zsuDV72AUS8qyxcfRTneMp8iQ7g4d83y/jLa
JDDIAvG6jj69ptKDME95dLc/VQ1Zp+Ok5lWCrga629CAWHUKX4R2EJlosnZk7FCe
20bbAGpn/3/WzBKpxSXKQQnLdh+vlAc+tDK29lBWeQ/lmvJX/D1sjHhwcl2uN/oS
CBriIDeb8IstzTkHqzMr9nPTqABFXeMUDuc6hZMy3kbEDoaK/UCyMt4wrIljBSmw
j2UkpeaGOFyehkRU2h8fG0ZSdig5A3vpr3aD/jzTN4kC3Jtf04fadbVx5iUN6INs
W7ExMfKeW+WGR5Bd+/TNbbrPl44tJf9V0dFLmzTBXPtiJnR+eRZoSZ/krh1tebfR
iXIda17jStz9Aohyzx09eMd3NMs622GjHQXpv0b531+3ywnL1uZRn92kAU0R7G7Q
i4oThVuYB1/qsiNVlCyRO8vI5YAfNugOpRTyJdEg8ndiFDvOIYwHiuDdSzFGZ+gW
E1uDO5Ej5FAeszT5Ckd+RqahOvOqwQ8bDGpzZ/9EkyRMQwYZcKpPuqeXwxouxMOA
rF5KQd9psn5kTuLOgytifxK0GziECBDSXYEtMl/4ICt2j+1qW89WexX1hiSKCBLp
NQhSVgvymG27IiJ4oxYM8g22GnOrunp7IrcTLcZsqcNNmsQcl6vcnzDfJtqNC7nB
r106lm3k3SfruX9+0DoFd/tvs40I4v6TXihY08p2Git/wecqIwFsbKLbCgdnDvqe
qD5aN34ThG0vdkb3xASIfcwq3rkhu3CzuP9x9cmvMuayqj9hkprxqJgQYKjqXQQw
l5XqW3gmt6VAfAKmky6JTWvNmRNrEaOUMSufYCB+d5lpBID8KgaCzxArQQWXdwgb
NW9ynRrMBEz4PsUw9l4RZWLHSI9PO2J7xizrQjY4j5EZAdhPl0kkzb0Bfk4P9JwK
I2HJKE7Ean/zD4nCysG/K1gJVFgXeftsSqoreUe7WT4B7C+vVq/0uiHe5jjLctpt
uWn1CVYVb/F48b/wpPUTyv2aYc4g/VouwRlbAPdp2/CdRT9eEywEZLocVuZu2WvQ
9hIxPvrv2ZLn4E/HEommicBFydx+m6L3nSHauH6P6jUao1mGYeCZTY8UJfsb19Rj
4QZ+10NY3a+Tm6zSfnZrMI+ZBHrjgJEzmxyc3Zxs4+CNRXiaP6xMS9Jlnk3MawXw
GRnRp1pBkbUtxUx/bR3MZUzxJpSwvZ6UdUmBfbwqTAFpIoP3aNkaonEqpYnvmy2s
pew+5qyOnHdM+gR0t8tdBluSzsEhtSqHuCW94R+XV0hw3yp/oKvSH3ju9u+r77O1
m3Y7oAWc3JHPEJeaU/y7pO4dlIwXWau5WzyGQjlPa+DszdrkvyIbRLbJZernNy8Y
zkT2MyACT+/PbUqeDeJd0LK/NMXyT0jt5Ea8BiTviqKT2kKZHgDWc1vyTSZClLB0
ZPakW349YjOKd9t/0odc9sXGUn6ogkulf3pLCenynGjwa62pMIR1+3z1Pb93XHyp
BeXGd50sRPqn7VKXIXt17fWQDt9xZLUxxUesxN5uE+lLvYxhWcqsLr8C5oYG6fGT
gm0eWlBGWlrdYkKlSF7RcTEZctEmzsssNgjovvU6SFXQ8hvrHJSbI8CRRLjW+CsV
8NthFspREBuNDJYc+m+9M+MFcOA5KQUkmBzlLIFxVLlnpavaj7GcYhXh/+/GPqNB
oWu8+ijesmd6X38DvfuOKY9ktqBP3Xgub3JwEXqQZlRPp3gL6/ZswvNP3PZI4Ulm
7sAXEFDexiJE7NPa7Yo9/qleDiXu1yzmnvOWaEeZmtHkwTurJ9ucSE1msBYeavLV
likV9wlhoOjeHJ259JIcOKUfhZIe3sk02H6J9Vl5dvliLElCnPOkyiSshYHQbuQD
BMt4uuZ42KMZEUFLwkV4rNIou5bAhFz4UXI+2m2HXW6PaBXMR4dmzgZSbr+TjlAr
t2VpoZVVMeYjx7Y0W8bgy9svbMosHQKUELPhXZc/pTKV2sF4AYXSds2q7LxO8pyP
IrcqQDuGExClLBXMj5OLVEaEm+oDKDLJekAlpAiDnrjp5jAvoBOpPB8RRex1goG+
uuLPMU2zHxhnaJryhyBYSYYmxg895KDDprvsbdCe8csZKdvXUyjaEhY8S8sGoU/I
UOUvEdXhf4mpBa1CdC4PXhXd1k3dBrAJuJ5MXu7ErrkIUTV55tfHKqsn4yWx9IQP
zoSRYK1txdM10WMa0vKPK2AMPVbKaaGUQ2i9wwqVGt8hntIq6iLgYhSoGWB4Y2cL
4cZBCuek9rcYE0gCi9FWdMwHVgx8z4RWj6wy8CFm+53XZ75nBPIpmsiww4/fM4+o
OgBJh7ZYAVAwwo9AbeZ2x2aZMTkz4MPCmw3lSbV7hTBOPZ/qLpTi86m7bJ2Ul40f
6plh6PKFeFgl2Joxwfbk79Y06IPgo5T1YvyznteqsED+YN9q4Ujp2AMlSKSLN7UH
/4YaG4UFI3QzlqeK3gZYNiITbqQxFAyTe/JfDpOhs6qbWV7F0zcVFNWIJ+VRuBlq
SU5WhHhIGdObzBJx7MdFAmY9Gewq2Mpfc1rz6qAY7C45klhZjrC4qf8HEghCO8cK
rMfiV7nb6TlADV6eUaHMzf6tKYWHqVauvszxq4GsM57J3VzgxcVGyNs3R16s4dCQ
Bj2F6F9wRs3pJFepJp+vI7OBKdIGcd5ca/bAxP8kWRTTFVCQhirjV89vcj7lXooS
xndOI3GN1ack2vzq4jFHpmzHSJj0ec2rF4NhCnDbagPzrH2v7dpu9y2mFcdK3WMS
xOnwgqXqv+onFDe3UjV1Ch8o4Cn5+ihti06XK5LD0KGuHSplkdYSQK7ezwbGbWzy
WKEyhnLQY1+9eRmxr+VpOCnG4ZxKaaMi7GyhX7W62lRFJ4ICcS0LX5iPadRBpbtN
wJt8oxDrj1K4JfklpzN+49pRlj15sjEElsuQtOjtXDtsGElVQP//cekXfwA6kGsw
GBXUmaeTsoKtKbjYoXtAKVg/XmuuGpUgH8Euo0nClfs21QZ6XV9e9RuyKjsjqbnf
EBcmmBh9VGFfzCyH4SLkkzw3O5IlWQxuc6TU03VwfZ/qIX2q8MJi7mhYXMzlgOlK
jrau8lImxTuYqZD6DplyuxRLUvIr7W/i7SUjDsafAUOcBmCGbw55bSV7z1tZt7Vr
EAhO2XQ64FptgqwBD3rwRyTxmjIuwOkESzt7ku0K/68vYv1krc4ldnSNgcYQyl/K
uLLhnLcpbL2z2tKNTGsfA4Rav1ESH/n6pttuxzZJGrIQYXBOgL4NJHilbgOOthUO
F35Cu12W1dZ48CbkTDXr1nbFQD0ulwZSsdUiRda8WlJ0JxQRfGjNR322qrCJynGP
J+hg816sL5QIH8ciHJ6HZT4vDcKNc5ViqQCgqhQUV5ZnhdpMnGQtho6uFCU5d71d
wBWQw1ZuHkerG12uxq1a2tgWkSCOfITcUR6F+VKIVL/ngH+QUpT1deTY0XVZh8qp
osopYwdfKrq13Q8BKYQD7Tt8uMfCkdKoNy1mWy4bkMc+ZSEZy1oSTpRGDaDAMIxd
RPIVPWpkORKUh2rThHLJJKnAab/56ttEiuG98pkUInjxA3/qgCXYQS1WjB2RjSYj
itNFMpFGTkz5cLIXqRHkzFcUYZabRXiimXz8rtQTwhjWR6kSj89ixbeECbASHk2S
7hubNBELrQThkBvtRErPCOUIlne50nNSJ59Ort0GatRSQ+axhMP77pMyPs9CMvaq
n5EOz84UKCZeG+A3s2fU6H5aqMhg3/bbhdw9Swik+hoTosCNj8yJJb9aG1FMNFL4
cM7iQEyCmlH9l0G/f+ruHHAPbT14divVTFA+up1qn3gbbSEz6D8Z4pA11JTtPnCD
wh4vT7G7Pus5Y8Sj8eVEPRM0gCAlUv3pw8pfFcr3jMtQSQcMYckEoMVZZtOP0k/g
NzIRgFAPjyOXyDFaL4FxOZt7Fa36FjCPiMZ7vRx+OKaVZhn/9k5Uugc/4ZrnWCzH
s9AgOvQk7jNIl/dmUBiV3SReArZmbxaVPf1CMZTsYO+BEFDhlYCxbh8bcpyuQgql
DWdNoqtan7Vr7OtgF0kpbctxr28CuaAkQQS1qO46rGMfZeIbslU9A27kkBfdidEL
4HlpGB7PpiiF3kjubqHG3ABLFmUYNAhr+ze6SR6CucGBUd4LK7uEJ9e2XBgZubop
x1xhIZxnXxoG6hg/ZF9XPLT2WfLmHYlGxDCCVqyfDMwuv/AMX0OMN/YwXejBtXNt
QfshG72lff0QDH0g7aIZ7saYFiyFr88RPbG28EbQfJyfqQk9syXlDETtprdCwOjP
cXeJFQm0b184MH7bC1GfaO5gz30iJoQ5CaTd4GO9UNN+MlgqXjMe4Xdju2F24fTw
Gjq/2pRxpvigAfOfAoMcDHe/8XP/+U8YPfmG2yJdJysc5C16Pys3k+R71RFjKSrV
I2Yv3jdHRDh90+UBsNrvPchUUnPlChsHrENcsfo52ZqKZ2cpLH1jiLRZfD1Mmpvj
cljKRpyZVbUaasOPL2UnbjXyBnRj6J6NLHgiIVLhZHPpVhelUBX7EJCYB82Gwjdm
S0ceu5QZv7y3IVc+DNX9LFj3qDexCdvTbn8MhcPwOFntDj7VoOmzeijUvUml4Q5d
NaGFx4o5oUofzDsl+pfoZ3dD9RkzdYe7iKSEWK6FheAArtJ00FhBaAwW19YTVoRQ
6sGyLPST4ifxRv/3+cj3cLwiNpwZDULozVIhGn3QI51o/jNrMtEB4r7mAhZ8zvwR
epcsG9TmN0QTLX2J7dPMkPjduIoHVhpvUVvX3uIMveYPPq0kRsE7Ae2leVzTJdZ+
Ce0BF6M4N+ZpVAB1mFx+swsWXkxW9gvNlIIBl3BMH5urUBT9HITCKcEE185c4a8I
fKmz18fmSQDGOK3jEHU0w8wCFQHjvKAsNw+vYV2SMfyDV3tZ9JflG+Qa3nq1I/06
e8Ipug+jBTNChSLhiCJPQmWT8eNdg5y9i9ChVawRwwRHYodnS3jxYN2fNzGCN2Jn
HPVoEzSqvFc7dSuho1s3QoZwlk0lBJmwiEgwv1L0s5vZfBJlyjlKyLC4OOx+x6dk
4FGeKrUpvO8RgZ6cPjYJjRjc3aAJDIa9jS118LKMq56GlGr3TpAarf8k1PgOfInp
OfE2B0s/A0mDYkueqfhF1tGkeZ6TIz0VV2HMW6DJPoz1/M/XIQpwvI0zMmhZE61G
UIdsAfo89g0cAtEeQjg+GEfw0KPJIu2KlzGzTKFNufRiAMbjmjNyfthl6qpZUITB
7HAioZWJ5eklQ5Iqr5KRUldHlRF3WAf3wYy7CN6hVfYtApxJrZ3IrKDpDz97ZryK
QORrqF7LSpnsbrfffmJNMsnQqaLkzXo26N55CJdP97Xq4lcILGFgtAkyHuo4gAm/
ILtCXlpnj0tR+zrtSufd4BBuSzZugo5cgrrb7YYHcVZ0DcYMa8tlTNZyN1OUp4tR
LypmCTL23IaE+uml6sjiJTwhHF5hmS9y94ffAAG48E5dhy94oHv+urEuHt9Lv9Na
2pqToSBrSZTUEPZOqrOerQRxpGR1Ldwl5p/ALQHzVzLuTJ9NYUEKDOCvgY36Vk+z
eaQtkjn6g5KUME/x/cLHqKRde4z2GAqCg4GPn/YzsCWFaGqn9awA2uc9efMd997t
UE5r1myEtQ+Z2BFr+6CeMDSlLfMY2LL5u8u6GpRlq1/aJoVwVSu605f73ugQ319p
0MV1fJhaJJQLSlnvkiDVjwCCDxQsqax+2H5o0eT0W78u9qqKPJlbJYClAi2W0x8y
iBEiqLmVGsGq4T+Sx4/jjIwGPl/Y1Q5rS7lI76IMBzDrLnv95wuKSVUX9051Ah3a
hNENIMVtE1lKT2myWIOppigIfhAhi9zx5GGpoq3GTo3H6aS62rTkmV9YWhgK3QT/
v0or717pFxVotZZ0aGGR/Fqqd+b04jXYuzD13Vaprygs+ESupvfVpE7YINr/dcxf
F1Oz5wslk+tgOlyGuKud0MnNl1Ni5TL49rbfpq4ihjDE8bFBjNgmU/iNojOr4NVs
nD60sRBro926e5SNZ4rIclJuqMsXCGJe8/8c03UK3QXDKrxgjIzXESQwoHtzXyVJ
GABGCjGrCHP/wqip2GZvMheCFS3pQ37Aad9LfuwPrUTReg3nUFo39IfOI8oDhuFm
ky5m0iSmi0UojQ7srrD2f2x4G/eqCxEXBT7Z7khGV8kNG/g+GIfGj2VbhGuEIHKz
OEXamIPHPWrYNTjEnunYYlD2iN4iVMw9bSN8HDGbp8vK/HV5gjJNjXgf4GJFdP2G
aXDj7MPPP6v47L4oug42+BtWgRV2BuPOAUV+Tn/DkcJ6OYvynqMU/Kxc3U/UK7fN
kdx9+ZzjhPqIqzZfLmB4g4VO4eEDwElv6gQI9xFCwTlkjF8mGbzeO7yBCi2jrnMd
yvs6SPLawOC0HCYEXO05mzkK7tAs8sFs1yRmHAxMaJ7LDcvXNpfj3kS1mQvdZLcV
xK1UojBATvvQMKHwhkAsY3MY6FRQrzDePNZm+jiYQbSw68PJE+7X+0Mf0rQ9qS1X
rGz6NOVheEaqQdIOO2RsyA88kRcwxsG/16OiJJ+9iszaXfYoOqDrvvSFby0ANOsX
kdNBC40MVlBAf9naguDGDjdHZgpZzgVP0uX36aWiFyEhyTN4en+mgVfmL1ets3td
1t40k1bFM3XL7PJUm1LrrxbtBlc8/qI88mr0+ZWeYmPtFKwpPhEIkybzpJfKm8so
JF1tJkzQNGmXt2r8ziNKUTeLsQkJO/jU9Tq3ZdaTzVSDYZXKn4TUcjn9coPpngLG
BvWeVmTNHr7fQnHTeNrp4pbzZrRjcdKv9YPf0pYjMkp/bFsKu1rPFr0pYnfbpYng
1RIbRKD5asHQ+YNUyOqhHELOHNtyF4QQ32oXii8qdLOj0mVHUQWi0gQaGsEYuLm9
zSAtX6lGtfOrDmmRH7s6gBTxDJCT6yzxCmoMbv/YxFJ/Pc8wqbF12JhxY4faDY+X
tnF6swrCiryCkYd3voqEP8HeFJWSibBu1K6kQoe2ZeO82fbLyFUVnwNndnq6S0No
SD94FwAh/nLHT0a3eFE9D1RUCUKF67WdfKiphgtapuUok4HpTwfIo/pTQE5tnwLe
eeBe787x7zrCNtYnIIqgTmMs4jaI9h2qk3hekg5KJ2eayzfB3XTlvT/tgyobKEfO
RV5HhlxcV7rK9BHIGiqZrcjKoTodLAuVF8/FetFqgHsfsNJDPThLEO1JgpgtQIDe
hCEoIX1fTomufGW4ImEV8vb/5BWchDtdMW/d9zQRrVf6Aaomx94+xsrJldbUVRCT
UOZ/yLkSU0t7vXuKlYDvcT8yfAnLhE/ige6SmLpOK+ALXlT7RoUvMVA+1k3astVp
5kilQ3n3gXeFRpj3N2b5+CqGUU9djO72yic51TtPaaZykjHYNKzJQRrk+jK7c5Pd
DQ9AyrrX0fQ5DgZf0Ck/gggmP68iicqGYtN0r1EjpRt4fGf602ha5O4ZZCu6vlQG
mJIl6qaurhlFgXsZnKTzQ1msEbU156Rjh67AGeA3Ye6SmbFwwWhS7mTBjwIu8Mrb
igzxia99+sIx1kJ/dAPkvLx0suFL2gySBnxd/Aamn51WsBP3MkRoK80nm7iaJH2I
tZ5QdxnxNh6AimkgYZ1FRMGSLcx3TuXNqnIV8CXK338hXBR0hp6zMuY8q5+DW8+o
3+yfS7xj38Msnq2WLdUPP9e5pplXjeqjVBvySv+37pInuBGRIWBdZLwqbRC+RFtr
B353vMjJhLY7h0SLf2DRoBGcF2/q/Lsq2gFzn6FUdwaLdXXZLC6/FHr0+FU5MXOe
UaKt9FrXxyQFgHSNtSRUngf4DP3T6pmj2GR0wCHvrN9VP5sWyZyzbgAOZw5wssEc
45MBO1TzxMtLJPgFSbFg0QfnPHYoSg1Li6cp+LCfAQPN0xAUhSAaKZcq46afo/nG
Edz4KsoI2PXxR8/IMENNGk2iJtlf9XZd1b6cqAzT/9EGJoHF9VHA1kSs/odBcUmL
/8xaf3y1q9xUGUNJ3ulaM/P2Ma1W3FEBKaqcNU8uN1EVE5x/1BZ7tPqrq/6w1Vo1
j5TbvcO9fsfd+aBwJZNAwQCfZ15E3K0UCoE6KHn1cu8imxOjLduXmfh/btVWbm/C
LDBsHoVqBFaXPS/aWGMLKlaQvZSajGfuHqAZl4p7Yb5z2MUCyLC56uFjKmVcpYq0
qRJyScuMTJBicTRSdJv9DmfGcALwmMOMCHY15rZKNMlPA982iv7Lr8t1pxKGAk10
9liKEt59Fv8FtRHUjPrWSBrMswfKTyqIt8+v1S5EfjlcRPMVJVFSdmn9Zc6OMHxO
OUSuopWmElngTX6XX0rchaFnED1ZK8aIXs7TkTXw/CFRDTdroCQqNBwx+ORTHqoy
c6r2JdBjFSfDstfLHp3NYspxbwXxLOqPGw4WRhzMf2ARKnVcLDKnDxCGqyf7TNWe
IkHdOoGH5i/1+i4wCf6t4dkgLLu3sfXMw/eU8e3dKtM0ItWAps4I5YihN3G/53Y+
QwQiG8uKhFTu0jhkcIw37MIWIxvZ1J/6DvG9XqQYj6Dl8hr9on1hhz4eo6Nh6FA5
at4toxM+a4EV1X8X4mu0YEgP8JOMcNhG84C9/9CGgLRSVfI8PwrAMzYij+uZH63m
WnHwpYN/Yscl/r5AvYPvyffKZYwXkVZ6CkB7PseojYIGqpJUaIbvhJcxcFCtjxf1
anOruzfF6SacoUlXv3+wAcZaekUiT9zfK20Asapf2ssr5dQFoR5+M+rnFSon4KN3
0thLP50Vgh89GNAvv4QEPJari0AKeMUZI00QElHPpYwWtxpEhjs4SHt3H7exGurB
zi7lazQoc+NEjlAWaAGTx8vD620RREeL868pwe7rxPTZUyDorVs/XbDMA5Pxhx5J
IGAqIy1vInuzd4yxfVuEl4wJEMh3RzB+OLdEUZkEM0+FRh8MSvT/y4g08iTmKxFm
e65H+NAzrTM3It0PqqCfRZSP/xuTiw0auRkl8bVK2pRRCjBAwG2TrpHjjFpOHkay
/eXVekg2a7Et4xIOP0kL7jGq8R76F7uRUzIKt4suMujKT44iMHZlibhvsNssxS4z
m7VMYkSetW9VJjoKTN49fQxShIj0KugED/U/Ma1J/XpnkmNKGoKHCewsVufafqKm
z4/zHgbZQsl7ue/jXD7fIVapHwE+CeX5akYcC9+1hl0YYyvBXIe3Dr9TXbKgowc1
UH8RNHHNgwXzHafUOBZ9cht14b26r7pt9dlpVelTMWkZ0Ok1AqPEg2Wq6RziYKPf
BelW4ITz/T5okUXnmUL6cC6wpFG8BFq0abTAxJ4GuIKf3/k95s+CYCHak02A+DIS
SJ8awqfDP1viezzmEjhMLMCZKPfCPL218hDIZPk5c1wgRb8lC2+qXUyuL2lUs9/F
u9BBX9YrTG2mLV+aNkgRwpJwfCjNuen9mL0ZavROhYisldJsGVgNHz2syLN5/4aN
AJ/EPQLQ1AR1gyB4mY/iiYQu9+M5y/mM3lVONOQ7A3ZjDLTi1eASAQI81K4So3q7
gTYdAsi9RklgjMN8V3qDqygWZcex4hQWuhQu6kdoj7kAQIKBqyBOnex3jM3pOFoe
ji5tMxpUDeXPRaXwaRWmc38VzbVj/uo9Lq+bH+e6S5JD/Bvi1gJ8CqKb/I9YxENa
ScQEBGtkM3yYLvU7U0/TbOTkmFNKtgOtDGuTXwiP9FztYSXKPlnJ+shZzeW3Cu3e
Rci4X4G8wL2Bahbi3ppweVcQD0Det+65EDuvYhtlx5bAmVTSDMKZGjrU15N8Z7Bt
l8jhV4XY8SBVAoK/pZ0X685Mz5LD6C4VaMx6ntEtlGP9iGMGRm7whHEm7wm+L1xR
RTA27hu/9VrhTUFRvq6LLkbyY5xPAlYYdGXcwtmQXBjai0zeoisceoXl4eiRGAbJ
Jis5ct1itEIkC0uuLpmqAf3KBW78GGM8n5cRzNqvy/V0+nrQjaVr9q8OqWgy+7wQ
TTriUU5y9HEbUPtbyBC3VG1rmHnNzWkgJrl2GuVlwzB/bChu/yhEoknFiTCUVp3r
/xDMqyYeRonn8BUnnmC5YI+kqA3vSJuFV/iZVm652UaYw3PVYH2HGYi6GVvNgoSG
07vO/BhVCRW24KWCbfjALxfaD1nyujLxbba4+7nVXW+cr/pITw6EuyCMVFgIWhNF
2VfUo8n5ZbdsXYv8PY85vCCsx9hi5RYuJiqaR2AcyBqi5ng/dhP/ZVubxNlFmGK7
QmERBuwYzgA+Tij0AZkhFsfMCSj4ukT/8UOW0lp8Ab3uX0STRFk24ganBJz4U+hN
AzUdB2Ctw3iODm7ffm8HyxNMMMbWJvElVu5f5KVOpBq2uLgdtdaj2gh8IZXevOe7
WU5YxEBO/8Z3KiDf7l4DzE1eQhZQGz5RUR4RqlZuShGuv//AWVAw4ctXVEMS15YV
ZeRsazgE6sUMh8//INjGVF5Hid95tfP+uJWFsLnMprmOCVjwwNs5iAGWbDEOJU+a
XcAWDX9fYaVtUVxlbDKlzgFNH4nNFHm7w9C1d/EdKyEzJ6L3z10krdjIXEha2Xcm
1FXPQMbHsQED5mCM61trXk7veahsTiKTuDePUSm/k6EdqX1okUeCCdhl3CLeOWiR
ML+9M6U/dS4iteEd/tsFav7oWwNn+nwTb+/dCyw254e8vlt23L0K2YO2sPo0EyH/
UJQA5KtWTC7Bi+DVC5cDhloUvWMJ5jRPR3UCWdaPWwZ5QhcVpD00wLLHAfZ5Td3r
IPjnmarloFwXbvUx0i3Ycu1vdUKe4Cemb/etqD6XkrHz5wdcMOa5yMVMkRekCy4C
48P1Cz35vkx3oMPrsPOJJW9ZYA9dbMth8KS/uKUg2T9Ru9qCFXTmW4BeKN6ws3W7
lFRXH7cn9MSxj5KU9Mpkxj6rLC4C6Nx2FMdyloWGw3q8M57wv00Y45IB6bdrJMpH
WpBlR0E1Lu6cA/70SLWcuo7+YjNnOqFA1kBhqM8+iudMNcq3iKxFCzlMLF8QLL87
TAdNEncEHWC5mhdO76FOCmIJBN4knMlkjD5KKtFT5sxUcNsfTUXPsSAc5lpRCPdD
o5XSmhndiZf620iEpmLIZ2/XAyDx+qcqqB9SlAKqcdL0wRp3MokxE2vOEWKjGnTF
mWGM8L40LZ8QzIKTtefkgoLrHt9TkBmz2H8R+5GCJJcpCGb4KsnHE2ZKWJ3xELr3
453vwsMe8WwkKFScmyD88HEBtLdtEYfN/AmdmoSO24AmKRySxQSRF+OQLvG1bgNZ
QEKGRJTC3ifEIPtBrlWMXdp6+G4i2Du5Be6vzHKRY0a7TacYbmCZjn5QUxmGXcW9
rgZMlDoF0lLOzsszV3lHInJCueO+DbVhqbSDHnpKELnRHGzAE/bg2EyjYoS3HeYf
luC0eWyWO8c69Gn70BzuLScpLTT453jUiPfnj7rKGaKIPCEVesRYZuT2c9DFGI57
KcFaLbBDpcoNzDRDybR16qh2bLqucyh1AT6B6gpMeRqfioGJqWR6kHQTlDlFwEsA
7Gf8pge4fn9W5O2hnYwGX6v//b8Af5bi974OoxRiT9gMm5CAcpt3McCIxs6MUsN0
ZR01fYmrL2C/86D0Ths1/rFol9KUQ+wTpuebU4qnt2WOVU4L/d6PSqwEBEiX+l48
YKH9DR0rZvfY7SLo3z+pgjzrBnzzBQM2Hu/udqM7e/aWCJuw4ABa+s7nx+ak0IJc
6lTuws5h20R1kjZ/Z8HQCI7T0KNuVzqhguUkke9j8Vd/C/ZE2tq7BjqikA3/4N0g
e9fFR8vfVa1EXu5pN/3AF56TECAzOyjMjxc28YjM6N+UsDwJry7s/FlbVho3hJAL
xOxIE/IwBbL8e0Nv+Mv3oU2crYuT8PbhiZoEF1FUDt9GvrmMbxzgHFpfZ6QaFYff
em3Ir3fwwc+psniEEH9y0qihD48ZbGSfsh68sswQDEX3wqv9LEXoe6d+U4XtQga4
CmKp3gxSMA688dpgI/cLcR2mOtSnZWmwBnQ37HxqU+KUwqGMdR92Z2Q8TXNiIis7
ClaV498UcYTmzT1O77hOTj8+8db6pL+jv86QICT3jYB6DSEOxUAMJ0496adsyz+0
o/CO7BNKmFkqpBHMwtspSiHZATkAS/m+FtlcHefR5+kJzbNIcvbhpIBiEw6E1/P8
QbLSoyHeN7FMnW3fATxa4P55SWvd3iuhy8WbvkV6VLC8EDbv648NGXLV/5u0nMwM
i/sDTEsc6GwDOptTPvzfP/pCI7LJAdQ81Q1ruNoE3dH4y41f3FpzWZohtgzG+lia
Fo6xa7fR65PNvY3Q40UrqZ/MBKV9zEIZKzBPFQpE34gfS7WSHwyjszR9D1Mx6zDX
VmP5CJpSykzejWdzMLMq8WV+3TKb2nuwFOsJXnBXxeLRNsixq0w88JwCt7ZsWXwS
hT+tMK1G48FOFcWLGB5X7OwUQ6xj/EashOnUz76JndJ8n5k3M4Na6aW0hVkC80ez
2fUInksZUOegr1FZApiJPsNkd96XWXzXT0K+Gwzj4WGUsyVJjXu2fvwD/lmhHiZ2
iuO46b0lbQ6zrI/14V7ji9zjCoQSlaViBsWoQxH1AaSWmtBKdXyYwKNIaw9krMgo
c7/U4DuJztdGZ5Nfzenokfvwtou5aGF0FU0Zia4iUYGGovExHtWBks1Df6lcUV1c
Lx2xZAPJgxuR5kINvKPlFsAXvrmVivtsYUdriuvonowkmYSsMowY9SIBbT8tlRVr
58OO87vZc12BKujVe5mwcgnERzb64gREx896Dwrmr6bN/GQKa6Zii49zMDLuE1lH
6PvLA6NcaHTU6op7lUfHkGC9QSkUYIPr+NHJ7hl3x7xIzgTgOxCo6+QP6XRKfrpe
z2G/u9dRRVsW0zy3BuTXcu4gKXFgU8LKtlL0fE+OpyExrM8+xoH2C0Ku1Q9CBFit
QxaxWMLravrA7bAZaQYlapq1vUwqQ+57WzJqTwUmTnzXMnebVJvvpAnMbS6btt8b
7iZ8sh+in3L0cKRUG9wmhR8Q/tUT03VjvAuLCNC8z8WZjOLN4VT1AF70WDlCmYx1
uM0o0xk6crtuQbNMGs146qQ6/9Olki7pDgggzHS9FtLZRGIXr3QDhXx84a/iz8aZ
kdhymlq3kVWLPaocrq/5QTJiNUsep1SmdUd55FEhgTJAbDTm2D7zPzCKfpySzPop
TGpxqR3tGJo/EsqZz8xh8nMqU8BXW0HUvCuPM0ZRpgjDUjgg+WGkYb+5nA+AWoT9
rpgpdgAPx8v7tlsWUCE9Bd81DGgFtuZnG1bQNFH5G55WqD0XLjrXkAC5wzNwubrn
2SLlp59RvlwF9nwlVulzzeaoHEqEXUIPC1PbRzaxrq++rVoxYGqFpmFPG34CJIEr
qd6oqMDxIdSsHohhuWQOekHi+jnpqUOeT+XwgzX1qCZ2J5qMs65Q3z1/fyHM54kR
ZxN2p0zKq/GtOdoEN6o+6oiKZ27fh7N0yzULLkHRavbcZPJ3bBav+Wyr7/5xIKBZ
qMruEHLDKphS5jc7ACxKW/DmUqLxhJzTVcm6GumdwG6TgmuZd8iYbJNLl3k113ty
SOrBUZO/YY/ODv7mh7Ecd3GdAidCNrLZDGKN9BmQBWW1dihoSEHvbWpahqtE9TxL
ILTDUarzaVJAGtf3hcvZUy/wiBj2bnaqNaHt2QEx+iyFMGgbpLNF3EKuf8IleVnR
c4lDfBKRXeQY7oK7CkCeDe5ytnYAeC8DKhVZ1pFHUGCXRRGamrYpP22SqELeqAS0
suLp0C4tiB6PV+jC5Tnxsb53INJ0fKz8kx3wjdqEwACv91Ep2Id8K5LyQb/BgB/v
ea5d6yJvnv9DBkQShoV5P/o0YPVfU0rmS4TLAaF+4aTRzK4tx+rrf6zzGSRvQwUY
cCAandJ701GFWcMzrmx4YwirblFYcWDoPg0WBTYcdlJNsaRG7CFnKM5on4k+B9KH
8zFw+mei96xuyR0WXH1Bazb6ycUZJUAL4pZDf9bKOXwGdVxBOnVREwvAZgsQUNI5
5BRCYWtQPzFx/evYT92BOknT7Lq4NW3nyQp0trfpG+uqBLhIQj5AUHxsIkhEH1Pg
Jiw1d43K/Fzv8611Im37rWKvx330qTZ7c56SwEWvf4Qn8qyxJ46rZHmTYSEMdDgS
+6Vbfbfg/39OMWraQwj3ZFRXUZ6A64pg2l6CWv+YEF/R38akg4BHuCWakZmPf8mm
oGMgPu53Mof4wWbcOYH1KwvP6J2DwiCmUUvc3lwjjoAUddt8ITk8q4qm+NbaQ0DV
8IVCrIl4XmqzcLXDyBqVNyUGSklXUtrtSioDbehabMkk4hVuJMmX3ZGyfWdlBsJ4
mjxupNyC4Wb12+yq/zC62ksG5hByvzqIOc+yQ8Wxi8bzuqCXfpUA+1K3J408JtNu
FTsca/s74DIQYD8uQS/ECpqYeJEOfntpcqmWTA+rA1aGAYz/dHBCB0qz5823dLGg
lc11eODPWVB31qgwzBpgcvLBwv7vLP2sAHo6KpCaTMMbIqroA83gtMZb4bNRdH5e
G/xegWM6LuQnBpGWS97WWMMTV8b8LaBkq7lECUTU8yOuLn6TXvz7StHYhx0N7z+A
R22gTAjAxYscpEvUmxiBTuN+/CCgn6pKBOp7XJ4+9gIzzH3IUCu+s1c2iXoldR4K
bREXMSE/Pt6+2lEVqFmWef7hQDiLf/N/lAKhOEfTIdAfzht5+FbYqeBu9BvbZN2V
9VYyW6rwX3sTx/A0ZJxqbgfvVN6muIOuBHCF7g08lAQZ3IrbmBDcfZP4PBtdOBZY
3cDLukEnT726/nhpM6X5vve/F5WBV09OjuWM8LpNZFMzXOeYNOn+JqPyGQVpfufO
TKBZJJD2j+HLVQGb0wsLFEHjblG1JSdrgaVZMlazuDTLjc+ak9yvKviwVoAyFGXF
D4lWs+0BG2Xbhe/aZlYwCjDGXhOO+RdI8i8cYNgMYiaHd7a7018fjiMjhFsPOws3
wsDOuJa/32ht4o80BI461Ob/z4B5bFwJ/osSAQRlPA2FBJ0+QfpJJYVO6ZCHUcOB
ZV/gx1XeEzuU+xHo4rfP9ip1vnC9crpHkEuHtbz/ZtxOmL7lpsucnLufQ6VKn2WL
J5yQ8xuJ9SPHjWXSyx1qXG7F/neqVUatWsmnmDQVXMsF4QhTf2bynIlm0sUL7x61
BO/sl5vCNQaJianGzqp3q14V1SQEziniJ8oB63XT0lCcS9gNbrkaIp/HvQbQ26wI
cfIKJLQeAgEIoqHNG92X5FrBZkDTPWR+UajgX9kyKhTDssJ9W1X+icy1rrMnhn/a
i0WniV5fHl91BBrNuEQlKU0dl+kluSDDZriaYpwGvGga8vIbN+j1DzEynkcQvy/+
gtDj/c8OcHmt/BrFW9u+VqyOUSj+PhV7qXr3c2UlhSa+v5fb3Re3l+IRvWbQyT0L
Yw3r9fMimfUVw8XLtPGrGi0R9qLDIliUJDx0s4YDOcRInwLvZxvY0NxZTSNVef+K
fpGy/TxiS+2uIOA5+ZdPct/wycXLPM41sSKiOPBrWhHR0O9yTGzelAP1jwlbLTWd
7tpCrW00OuNfmVSJsTgF0REHxRYP52Ntd4IR7khzTujwupFX83RiVryFpSlCVVzS
R3moL3F5vFHx9aP97msozLZSkyNU51j+mxuB/ZPb+SNXFwoZwmTvKKS5Fb2vfTHp
c8I0LkAiujaVo0M2gZ+3ViIch3wNgyMqWudyZblTEACcf0oHF8uQKFIDOi3lYhK4
rUrbhs5y8SRW9NFtoNjAUdzq9XC+FHzfAL7kVpolOKKblVuAdzepg44dm93paTjl
1gDEMV49fKHc0gD71ZhKWWIEkO8GESx42UzoW+vi08xngA6MCUxTinZ0R9Vdbd1d
ebP0Y+7MKtuwTXUsrMSBQRteBhINUfqhIbEYjPypAjF2qaef3s/heQagCpIaWYwl
pbDaAJpuW20RJTkyldDvAvWdQq9kpB/dtsQUFzEHx83ZQNp1L+im2aXairqBmrXW
/NzCw69nJFkDHBF3RY8kXk+Bqpf78H7zFTNtGN6JJAuXpVKhAN6m25gAEev2ff+E
n5+WGF+M3qA36QbRlgLM52Q8c8WHaaAVMWfpKGd2MNHX5QMf/bFxCrUuvQHKdfQR
zQTRLOJ0sq4kQxLdGamX9CcK3hSq8bKSba/VI6RZVsMLeWSb41w4JcWTn7R/tc2Z
Fv6phsc4vb5Dggme/2zIH3soQsbjaIUhYjdgmH4tbTCh8etdfvBUcPU2MG9T1wZE
lW4k+ZUc54j1vXfKEnW+J2PNWUTNmi7zghg+8zLwGgmGcuNVHVROblrCd8V64LJS
YnZCrHIXLfI+uPs311NzI5kQl0ee4dFrpD+Grt+6DWTXyTQo9p0uqLSRHYSMoOML
wfLEpfUyhAPTTX3f1zE+liMWKrSS5/u0NzvDtD7erQaoirlmmxYsoc77kJ5L585D
NWm+PQWAgIvEzyp5P1oExYu79W652KxtADwhVz0MT85ojediWkEl5gpQxt2gZLkZ
hC6MrbtzYS6vn8M5ecwd6DnI4Sv0B1SgIex7omO6f49unmAatoVB7806WIZHAu3y
VwajJh28Q4WObG0Tv4HEzxNdnB+Adciw1WWa4AgEmycubF9IS1m+gY+scspx1rD8
Hlw0rBdwYQUTTo79ojx5hUCu2Q3uW6tWCrN0UxIDcWXtWNpjEnuH31xMBPj4A7uI
79BEaBjOIDXwEh1HGhP+BSze9YbwBqTVtH7Xp9vu7w3dTCzKwkSiAURNbjGxWiCU
LPT377MWCzSis8gvIO5gRIUdvCNASMNYcpy01NGK5CY42VuRX7YZMksHt4+c+qgv
8Lb7Trb5iuReGxMqy3nIFDXfGzWYIBxF5dNYUKd6niGv6cGs5nmlrCiyndz0fLtQ
oYWmos+BWBpNx9MDxEzl4Cde7IxUUVPm5VmFKKZxvp43gnf/1nlU7yv2l4TTDytW
WG3eAirjGD1crXXNuf3lqT1L4yx4Eu4M6MKyRlTvZIpct0Zx2S5sKiG0QKzVxKcP
FbQOC9NOnRgNSanF7fcQ0KNKmXd4+AqI/kgcnCicftSVlE4GNZ+IIivwZhnFVIU+
GVutt9TKgkpNGOg8lZ3KXhofZ8TZcG7kR1ZK+21HemOogoBcOB5LF8JdbSjNRPfV
5ZHgGARnM5s9/SkrhAtIH4q+KKhW6XyVrEBNEmYz61mkORhLcjOWTILmExl7EwnS
533DPUE8S+Wp1lwQH05tGFmZ2JvLS5MeT+XqZPFnczUs/niGIvSXq54tilWtyvqT
5zIHYo4hwWuF1c1jMl7nK3kNdi790HK0riFE0EnOXSi132X5uAkxrsf4XJZharYf
WDRXvDcVeHlhQ2u3nTY3jW2gGVJyHUjCRN9zt8eGfOpA5c3E6RTjkyUwAKyD2uYX
+Yipfais2HOeYnNNUy1RBGniGaXeaFfR8kBYvPc+Jk+SCuQjRkPIa5vuN5QwQ34v
uj6kQpwzPrPSktDKq2FxpA7uy0GCubmXOnqSo4uVEG4Ln0OYP2KxNT5xoW90eiXn
fvzkrVMxl0n6Car4rrqwnlBKut91GaJsoJH0TIvVB6TF09JJcTkBAZv14B0Ph39I
5KzOBuMmY3YrOtH+r4s3tz00IJh8L5z5Z7V1354vFealRbI5jabfQo+GHcZi3gyu
b5zBwEJ46BIvs0BHCTJLqq2ixPJBqe8T9FoXf1d/GEL6goI2IuWNdDDcQ0uWbmHE
UC7hDd2gg/0wSocFCJM+2t626cf387ePzdMjQOXDBnPq2cFPwCIEQkJzOxV2OPUA
59Tpu+vxJMssn7Wb6jkyOfbcJKNj3ZG9OOWRwNHqDrTN8zvb4UJh5vwgtMwjXBPm
9HHI1pjsxHsaD3kUwWeQkf5yPmaNvBJmlKp07cNggqsKqMF5LRl19eIhz3+dqdzS
1Aiu0iqrIX06sG37EAbxLZAqoGZ9XLm+K2NOiuBVsGiBafBS8QCVspb3ZTsiymNy
UqvfEmTTeDHoy74XNMpnX4BVye4/acqh+2DqyyIMJL2B13PTF3aI194Ma10Vz3dd
ON8gO2aa8ggYUVVr7jw82RrNgB5/o1nm0cOIpT1lJ0kxMTT//dchlU5Dm3ROfRIO
0aA0mIePHk7E/rrtuxxkM2v9icxlXLOypiytss4eGJN7vSwTH2g9uTNLclhwX2ZF
TR2FH4XTNtjHv/BkYMyeFP4QF12MCHLZFf38/Lx9s+OggQ5tpmQof30iE5WdfUsf
z49B+j1HonC5pinV+ldy4FAzI6FhewIQbL6ISNN219ZTIakARSBnmSRn3TSrRjZh
t8myUCZzci4CWLNyc9Qq0zfMrbcvwgiJ/e/t4R20SPVddes0fbJQ5GzawYEVaNoH
DgtyR5EkKP+NRua3DfDk91uhY6uboGn0IY4oBzKMqyW47l7wX1A9zysiYhewNhs/
3TWj7UJTWGSJhQhfcB2E9kbdyrv5h6CZqfeFXV38ZoyGGR8m/2JCjha55Mc1V6va
GhTzBKsfIe4eT010QHrORTNzPW/4OPkYeO4X+J8URrmtvgZgX2k2gRnsFW7pAyfQ
M7aNgMpJc4M2vv1OJ8jU4RFGxr+KLnzey0QKItqtm/OOdMsgl2NXUJDltj98wtZz
WfyR4FJf27o+pG5Ac44zKGuj6+rx4tsepeDGrtgfrDQpRBJeCWeOCc1XhDXXV6Wv
cbR0xv3aC1VG3DBKHfbToAT7nTYE3mHnkWB7xLPNICMmLNHYnnnZFoGNIzttde/t
JoOyYLgZ9QTNLM0Mp9hCTreoH/X9dGl94xJ5KOoLrxTy9QtF9ZIKqcWZqbInG16T
EcA6tiDmeUTl5Ud1houVDMJUeqgclxhZDh1dpC2/4LiAEL5pScHsUrgLb/6MOhqj
D8M2sJhX2epzxN6McPeCzJTq76H29bimjILPAaf6FhuFjcsY8hzbEuCprXhjqKzU
cHFEXm5IWT1YLLZp2Aw995uPuDAPgNoKUEOcIUTWGzv53PRzu+DGCN8Ic176fA6t
ZLf5DgCKsiwtM52RFa0Kf4w17Iov+MFdfypQ3h2GrK/VXnH9bOKTvTjE5r3sA9Ld
VpAVvPCXaWsXgTBHS3g624etCTyplInjxAqk8UdBC7HKUwilKUKoKLyVahA4RgBz
XvETTyvFByi7b+4dUj6+bZVFEvg6mS/sOpk2uoUoqLbVpuTGWtesVU/JkUNNLjjC
6UORdiKHgaIPaH72byW+lhtYNwse7jqVU1lRUR25d0Ou1Z0hlQ/H2Zamd87M4dEf
m5vy7jZ3sxrJUpviyg9mOxjCZYKZbrOR3n5VR//CdoXJJ4vQmUPe40ghJzbst6Wc
SyUXpU9nFQCeNp+/X5LLXTFzN1blYlKtMe7zTiWfsRlKB0JNy1I8G8qvxLcSwF1r
N35sgxHVoLVOAY/Bd/dvPXSwsWPl4RVj/djQsR2ZEOyxEHVzHb0Ky1/FlWjvf5F9
0JLx0IwetWDJQJ9b57LXbTVxQI+rf8XZLOXFpqgCDrijI6WbcNfHeB+Lq1GdOS+G
3Ol86YdFn4PP+fRGWGIrEzyiyde0y/uvKEn1v6dR1jJls+utbjXRwzHvris7WX48
BupYWOsZUu4lmXwLcYJfLPU6jG/ga+1WfVmOog8FeZAxwFHuDjQgOK//tO1y8J4G
/+9Q6N9oaS3xGnpc2Ydcm+FZsq9d84fElNk5heZ5S0i01qXZTTl/rpM1Pd/Dp9Hp
q7pqRx1jMeiVuLfgg969EeSThBszkbbPnhN4IN2k+gbY2bIU3iZnvlBD6S4xSQe+
FivyUsmJJiGx97KTaAI67xqmvUmtUNLoBZ1YOJomx4RxZ2xkyUzaYJYQd5OXZDdK
jhdSd/Df6Vc+it46br8zF17Uy2WgRMyojei1S9AQ9RTn2ZEjSWvgPENEzZXRgRtU
VKTIfUXtOAmUcjMDMXdtw4zY8OHS3BVwLV12ecH34/V+PqnJ33yXbCNiXsjKTYv2
eDMJLOrzf2Op9pNqhl/gxlDFH05G1q7NlTRThXc21DPBL1FbSCBmLzL4eQR/CeK9
r/a6c6z/kawrgrSbpKz4UqWTEpaVpmai2EayQqoua+UhV0+7B9PEUTnAshGkQPdy
fdHq501tgN688QRUwBUW38VACu6ja6FP1aW+t9PqI0M4WKroBtY2bhomxlqn8jU8
gfVRYpQ68pIbR4PcG+7yjqsQX35dKEMXU4HukqwUZGeXBOzoTYjQ/wFplKF/SRvz
VLyG2udzpB9jaY1VC5NVCs7QhkHb8dZQa0BCJxJ0ziQ/OZYq6O0WEde/mi50ZQQW
ds2iECj0GBDoH9Vo6jcoG/2i+dY8eAI46nakDE9nYOr3ziHe1ItnhwXH5CryNfk3
cEQWDc9GTznWIb2IgNjE+O9Rfj9KwUfRiyovWhAHBEobnn3NRzFTOp37VmvXwaEj
Je34T4/0Z1Ta1c2NtBzlThWxGjyeyA6Lx3u47+cEkUcct2gPnVKFHtKujc+UORZS
22qLwNLRSGxDc5V8CKw+BnfVw7wFbg0gruzBm/eCMgxXZQimqfwDrSRDWVv/i6qY
pne5h9jgbsjrnDP+kmzUvUaguFUkeVefDqzeNem1fa6BADteHURYqb4TL0Kp6o3e
VAqz3JdIQ5ERjiZMbT51QlGaVGENV2Z1WdDvy6VafZw0qgGu5CS/770hjD+WNhyT
odBr0BzQ2S/Q99tDjQBr4Mt0+S3WWbkzJP3AW70VUxopVY3hepWgCzEV12iBtS9Q
cYxVFtjPnhlxit2A2J6NVAmr9E3P6FRRyeuKKjZ8bg3D25KVuN1sk2mHXHvlT0Mq
2PIQb5dARSCXxkCvJNiGpwPGSmT2ao6xHymDgdcr4Qq4J8ZsgHBCGZyiQMvO7G1F
zVn9LRIJwXBEvwvLheJM5/1Dm+YsGwiaPt8qsvLExO0rU+pI8gsOZ8Nr209ZN0Jv
ectirftEn+lT10ZyqltlaCx3kdA5fWesFxPJInkWMS9FPBmnPTzf3cX/YFr6RKcy
96KTa+/HLCH+o4DPuGLUUZDI9sYRUMXnFN7T2ns9NgdXmktCAnb3yp4OzAYZT9Pp
Gps0mhFT9kqS5GKgeLdnikRi8FZ0X5xJSqDjCScZT0uTTksG7zw8RzYjsSuhe9ks
uRWl/zyCe0NWq0ClnGpohy3INYt60dE1bre39tq92fC0bZ7utzAHih9LmTa1ueNQ
70yneDBXA6RQpOVyuwpmzo+mLmOlHh1mBNPnhrjaxJHUcbploxhay1CbS+kTgsTg
8HJvJEs0LsIzlln9Sj8U+Z9Tdhvxt09rF7nQfa5B8yZVZysfamCFAawMUVXgxy3e
983UfdoEkgHSqZUOzdFG75dBB0y2CVKPZTdD8yLsdqugTTIR/ctNIAHvMZlQJKAi
9Cj99o5olAz0E8gtZhrR/OQknYVJZ+bswk8526t5wmT+YjpHeew+pdOhN8i2G8sz
BW1jbak5n8nC2F9D9ICGTONkyhFf858GXy67sVlWiogFMo5FC3R+hmP8ixJcQkWI
FEtyuvnYXWl1jDqYJis3xoewvwpd4XAiCNqtmjlZcvQaTMmB9LP3nq0+RdJsBAGz
g8Shmg7x9FgTk/MjYzXP6E73E/HvIBZNg4CSI6eBCZOSz8lRK1zwnOqzHlh+4gFq
M2TzVImadKYKDmW8uuLmUI3w8GwHgYGLCDIS9OebWzwg4bJerzr+o0K9tbIYdK1c
J5MPZXsGDKqQ35UvmIk/+YF5OcPWtkvrLGm+jkkI9gpxtT6m/7eniGsAE9vNOsMn
oL7SfUCLQhn4mq757TwDUcI1bB7fii35Dnt9QVIsR9dK6d0/jgYcDtY1W3plmCE5
A8o1nGrGOsBYzqunGqlsK+dHQa/B0d6DVIWw4Dn/+P6BeFd6YV5838rEbYrznZ07
PQWEZZYw7VjMjsPDgEHsNDVKo3J0Qbj65wYptj3rw8NszYvxgAs9oSvMhzNjucxk
mH9OpmrPNNc/0cSEes0dG9q9bnRxjYYp/WznrE94nQkzF9k3xeaYpTuh/01WEyC+
dO/frwGkaroj/OovXUj06Ia9v6dvJ0aQiz8PxmMEWvoAX2T8CERzPGTPc9xcmGLW
ykDzQjVPkgL1uhVbaUR3BAw+w3b1HSR95JmVHgUjE6FM6CkATmEV8kX0oWMvScm2
9LYLwiWUGck5qJHxNSxGSUZHD/P6BdkLpAdFMZMSP5O8NhmuIZR/6FxXpqbwcmrG
R9YLPLaILcjFyWgU22H3dwc8GNrKamCFGkbForoaBb6Tx7crRBnEjo/xkQoyyKsm
VviDEMiUtGIQxvqqnsyGHi141vge50XYdIWJTAogzeyAiLLQVJug8fz7mR7lWZhy
jsK8vUgwtDCpItRePShLF1Buohvgc5D/VkIVqVmApA0uHbO/5T7AuFJs509DPj/q
WHz/XO4ufB11UgAKObnSh9J3qtYLPTsyphaG7qsfZ4CNjvsSewOzFJlZrQJ/r+d1
DYzQVJsmA5RXeoD12dsKeIU+3caJLUQKlmJikG+dz9ZvZwLnEqUfiv3vupWhjqw0
yIth/0KqkDHm7mss6IeXbBU82kb9IOC1qIs1GCsSoAIOV+HCzcktt06bofEDgoxK
AnZNlALFCORG+zDvEfBB2ToPdr25TW/YB1fT99dJzmaXse37KZPbAkTDGB3DRt0w
U+g0CdmGukCWox3dj6rGbBqGn/+AW8g8THCpw2FAwE2H9nO4l7TMsBymJ3i2nq96
+Q0AwCYb8eoK6SXW7wDzFl+AK8qOFMtp7E7CGpC1Fpfo2eQbgfBv21TQXJ1j0P6S
awgtUowQC+erWHMoHSJaQmZVYxLOO7AiZTOup9+rORrB5Kr349eQ7e0Se1HYBFEd
Fk8HBAFRyvx45/6WiGoopxxvWr35+0N+3gvhJxN5G8Hp67BKvGVc8Ro5ngt5L1Va
49MBqTo1+q31dSS7HLvuixZyb5KgXh4OF30q3Y+PPxhjwSHLsMLtqEEsO87c93x/
2KnSBWs/vVocs+yKsLXPVIXpTmZfrAkEFfF1F0Kqqjpn3Yr4Mn5a7F3vSzRSMV+i
KE/9nkbnplByZKaGFQNk7HPl+yQzsnzcUMFEoknhLOeUv0r7nILt7tbhXOT8z92u
50Aq5wWXFbEMldBE9P/24im+bJriGkK+PP+wl3RZ0V7dAtG7RySVrGxhG7YIKoBs
4LCUqwK8IyOIDdQnsTQ776uiuXTyShh7LkdcE1Z3lusVQ8Ttc+I/DnM75hCeyWXo
KW6mdVsxWvbYvEG6WIgo33JeREVV6w4T6vYbMo5Y8dRGSkv90OjiL7GOKVl8sUc/
hD7XN3ByAp1vZrSUkwk/Gwet/Imq4o3yXJrtGiaKCApekNlPcNnYMK9o+/IjrK5x
j440q20Py6dXMZv+8vxHbPhZUv+Px79tmVVXyVmA/Oi/B9ITOAr8GyiBcDg4bLmJ
fYM9nfsJvdxGPEqpSY05svkXM9KNTX+Pr4fCbXWchKp/m1UofR5eEAbKrB1oA8zg
U9Vo+fmhDewLruBC/s77fi458G3fj+RaZCAsTp/4zy84Sr5yus/vA0QCwvQcQhSy
UnvqDpkSNyGRZw0vHnEQV3FzycqU6IRDrFtGeFMBita1zBK2TBtdP2s9MNGCAl5h
N8Y4G6tehZPyBVvp9ei4yC/qPaJ9LOSw0sUYa6Nl+I/ibxXKESn6WQTDNS06OC11
uVHzO0EJJuo0Y+Fxr8OviILif7VpcwynFzQKJhEPx52NS2AAoGHHr1ZuHe83lde5
JODODVnaBvgt3cgO782MmP9FqyNn4bzN/lIB7kvoTcLn7bC3xEeQTh4qOjJslwgQ
W25EpVgQzs5VVz3Vl/vp6pY0k3W8T1beq8GupbbtQqf7CO2cAIOhq+mehyyMHRrz
xLOH62EF3lBivjoUOifMyYUN8Qpx5xkRTLaqYOkW+Q4f5OSgYYvxYlIEMMIRqRDb
6vzQnN6kevWEwwJiWYnQXuueI6bHRWV3TpfXzNkM6uqvvoiVzK93i6kJN3JpwQcM
VEomK6OEULMivF+2+Z6DLigQXd6+L5Uqni80YG+YZoTWBLsWbHWrwmOaHLynX9HL
kG+U+1oE52KPWGVFSVq2nTDYajkbxDq9/Lf/D1DrqFX4yLdzx8/5wO9b1CBWdf/Z
xUIXCKuy+UvDZ6UnQVFT8Vbw5GcMseqH2bLvpfMPrI0OgLUkRghqFleuHp9WHIV4
zzA4USUeufjxft1e5/bX6FgWbgBr7zEWSIXxmoy+8SLJJ51p2EHZJQspSXq6sZXl
469DNnwH1iX+Jflu+mzVuRCieQQYZ9HrJQvctroBuQqq14V8uOV/foO6HTOMsmfl
P98mEzu/a3xyT2TwN9Rhvinv2FCRk7MdWiTMCkiyjmXFRw245eip/+fiA6lERdKM
QGffknaytAprV6bh4e83Zg+gHudodjxTlf2YfYeh4JV9W/bU79ZThUKkNRdIbNNV
YCTbE7LjjKpv/0k0HD2qq/hdjbdeqkueh5XEawHe2OmbKrU36DbBovYoXsDqVHxM
zn/R9Ax45qd7fSQ8uTglYbY2Yad+1/B2Jg3v5IcwMaCaolfQvG1VpWHlsmBmW9L2
+PTb1Rl5zH7PZ75/QGjcmgf58X8TuuWJWr9LO4oLdiVdFLDbMfAmhQ+y851EeCBK
2j+GJ7JBHLAozN1/IRbkEvH0fTz8/7WNLUaEEzeflDe8Vet0NDR0X5EyFKFl4QHX
ivdo6nchO963Do0ksjhSibOdHhtYZd2sBIMrj2Ic/IpTwjXfsj0wmEdtTE/08UxI
xxnIhyrv4uEdK6x4prsu4TXt73NxZkz374YZZ+Nnu82kV3bS1p6IgnUk3C2CMq4y
KlywhjAPMoVrm39+oqNyLNKBmypaesPVCkHuEillUw+uejW7iCbqWw4k7AchflQ7
s1BxLiMWar5WQ5JrVlNqAnMWgYk4qEVpF2N1pC2sl+VSO932PXTVcCMaUwev+RoL
40N9G2ifJ9guub/+bqP4+AxnKFcoXWuf/YZ2FTa3BY3R8mbnyxwOKppEBCtA5Omv
4CWJgxtLOTHeK/oIGCBa4GHqFzHRfjGBwlk1gR3cChdLRTkgqCKoBxge8+uRewOv
sQQwzyn3DFuOaYE2fu3doa33Nh8ZLXCYrSFB9MCNSfe+ILyw3d/iR3O/jAu+LApe
OPHBQTQcY0Ierl+iLHWhxU7yyIQMIQXJLZKq0b7A88vjLC8UApvq2L4miShQm20H
GF6dFp31JhizQKQJ+2Zl/KWNQ0aJG0jzN5agjxgpjkcMeVkvBRqVfWLUvi0Uenpa
9jVlfXglEG/1f/JrrUzURqQgkCEyy+VAYHqcnWjxPsURIn4ECUAGaSiEtgusKQlP
kZyrZpZxSSb/IThTHan1/QZ7Ff3PsGRatTnaaiuV9in/oesLfcnWJpagkXLLdT0B
CRZIT/U4c+71o0Y+gk+MhAyj4MEnMtN9dbVt+z7eGEsHaK3ltBdoc6NAIC8/k0WD
d+OLsOTiltepBum++ffpf2VsM3SVbM0vL/A0yCve9O/jvbI2TV1/OeKpJCGIwhIG
e6QdNwC3gmTd0JfnixRQD2u4xtl1dKMLzR4lshupBdfileRlcg/qd/Pa1dqEX9E5
lWvAI1TMEtmOURSPdcK+uJyTdJ9teGBc3Hg1gmO/L1LjFMyqT1rnZuxdAEf2r7Yv
HtIcWGZpvRd7BIvmXKU56yawgf2gbwwawZ6DOA4el2Esfx4eQFHrGipnbo4mdQdn
/3Aq9+zUFKDpKnyMzafBpszzhMM9921eyEiptkqa0kdDbyiYGyqNnfsD/Ek2TBBM
1j3k0lwtUvjiR8xoOZyTU/dIrbgrLpczTLmdik8l+CIjohMC26blIB9snk7CpkPe
0a0AVSlcKfxOUr4a24sEVysPyYJqyd5EuuhT08xWqwUUTCS7IASkIrll+2u/jSZ0
qXh2Aetj1VhytGQ9wi8P/UVCMP+rFK7+Z4PNlTI4kJnKkULFZYJT9b88R1ziHNZp
OCHr1pkiA1sdhC2NIF5FgEdJAMR6B54ymH3YuLgQ/t7F3/5g5zfXL2NGQMAddc9E
dHAB4CR/upEEUqZYlJX1JLpvNmyYsE/+8G9jjvkq/R3VnDqtrBNxVW5D7YHqxtqL
Oo1/Xehtd2ZixB2kKKQpy+kJYDWGnj8xNFOdft02me4bpCsopUOcA7I6qQmO4+qE
3EIL0cvk/B8mqrCVtQhkHPftPH74dn7jNZJljp60P06SzdxVW9bhjkhP5cNM0ED8
4tE1TqL+go69AcMPM0R1kzsXKW+zz1uqDiilw3QiTdG4iwhNSv24UI2b5Dw3fgei
Jt02/56PMQ+RfGjjVjaRdvho2jGpjTrf2NOdPX/7SUYZA5hKfUqBHHXmVnBLbO0i
vMLYLjLhogsxuk7aK3gYNZ+0L/l3WLfsKmedpZwxKugEDxL7uyc546TTovgDzn9r
e7lltH/YpWfidbK83FaeQ5BLPkgW8RgjkfYquVmwXY078bYXUbP/m/VD4rkiGDK4
R5MpyKDBIb29majT2XvlQIjRigErdPWRFbY6l+ls2M/zvypmDIpOyMlbAc++lCiT
kiUiZ8DTDWEaeTBRtlXTEnTQtJ0m/igcy7LWZNFrOj7K1XVvj8QQxRmo81zMd5Z8
IJS+8uXOdxRGC9Gcyecfr0BLywdW3sjqIWl9T82gVyeE50o/CLg96iZAGz20Urz2
Vl69cz5EdZ9kOkwckcB75Kk3pd2+ajdB8QnRkU7SZHI/ZImFF/YMo3dsyrnrKWPi
G3XxnEgpJU5PBD5r/mP02kr0xbXt0vKWxQMJWtmXpQmITgNxRLMPS0mlFycFsVt6
8aZJduoeaBkc4TsCjMWTFXj/Raph0SZup2XQ98Iwou3NHjzzH6s02J3SMmi2/k+O
+Hj7tk9y8/1VFtDrNumhMZdZbWNjaNJ1Ub57CedWpBiZlTeJzALLdfrfGImyojB9
tI5DRjtyMh8BIOvnqb+hkd0XXhP4J/J44TOeZHhArA7vkOXaY0kjlzDry5OTKk/R
0jeDhn0kgQH2EE7rPIrRVrvtNE38Dy5dYkIDUcEqV9YArC3gksD2v8OJbuZIMtQp
wBQLRlr0AwYvY27jHZkrPvtHigGaac71XXp5JV0a3sPeHfISDgFsXn0wEK0ZlGzA
F0dokRZNT9d7wKpEdpT77yrXXrW31NTS4Wdf8c2wwKnrNXUrcF2h8PDwjecNZTiL
8sUKNcyeaZMBHYYdrNypAO5fu8WWQnfXgDgTKqGKj6lySmxpoXYyPPaa0A/Txr9x
GtKF3Ccfue9tpDSEkCfTEG66PyRgPeDYJW6E6soXf9HwhkUWp2VY0zKjQL0FCHiD
5CJ1scvyPFn+5gSL8JhtarBuJt/j78P0nZdqH6qZkCNdGSgeokpdH50dVezEEi1E
4o8y91o6eHBtuVVqNj2EptFvVQLXEJKCScsGDD6/D8u2cd7Pb0BVI1HrsgfTwsE/
ikyfMcvQHLCdPpYAIwbXcryLmqhcQJmL0WEcWMIz/nSf1tgZJzZSIkhFumT7ppvY
spnycXd2WbR1JCzepa80DpBzX9Lq9J9mYjK6l5IEu9XznfTw9UO5SrPOKEYXpRJh
o5PiDiMKPsC0XjRJR29ePO9MZy9xpBIxjOrG2cupC3Zl4T6ljV9CFF8+/TRg+nPy
jZHtkMOjVRGyaKPwr3Y7PxCKVvRmt2qwQuRhcD1RyYTLI+xFRPe7dURFEaY/n7d0
cfFTt33EY8KiMK9eJNyft4hjb4P7gPfDhRnPKjo287PGh6CQ3R+HbIN+jBr2y6TM
U9K+Tq5QvHlPJTCivHYUyX+vBm6jU3hU3JFAbnSWQ1vQFNZpfaizEH8NNklPitc4
COHmP5NY+TX1eQQoy0NpOZ2+J8SHDfrzrj5Eco+dGl8o0s4q496G/RwACQ9o8sCd
GGxNxNYwmfFd6E3kysCFiBQhlNRS4FVbEY5ejMwZUAj+OEru6wXGb+Y4NRjkmYsE
WGlQ5ugdqhhol4kHAkDUeoMqpTwDIB9GsoA5BO3zT2GofovZorz+idnLM5e2AMEI
206b2wGFh0dzxLrer9dayRBt37TGMS/ZDyHmd54XeOr07hZ/Ryh3TS24vFtNU3Ho
koC9kiIGr7kNRlPC2R6NakOGETHBTNbv7Zw7GW1hAM7vKahKR/Dwe1WLhjPbkeoh
27uO+Ss+KKoH0gLZ8UCrBqaW1sfZzZeo/U2ucBcefiDNKW+66lKAYQ6FeOYCgeYS
H8iQbFUuWMPSa4wK7+QAD9XIKcMvLqqINeWK6oGCZFUHEKM7tS9f8mqtirR9xjOD
3Lz353puaptZTpXpXIsg8e/XqOdpgNH17GJGWM4YOeJCXwCMnbJwM8t6K/u48GeX
gy5Pw+3BPsPQgdYPl4Ute9p/Mo4qWmrAqpX1Ulodthk5ap4a9SbZ6uv7b5oZOTgN
QXp/vL/kQK8RAvKf8z5DZlkoe5uamkJP9v9Iz/kbmUGcmPJ5iQMo8d874sml4FKC
f68J8t5NjPSpyCOvCGxHfLMp03YlpqQeGcfMT9/xUBM1yZdRYDMFu86D4pONr9du
pmsYgZACTZquPKzVigGq8bSGJQkKHfoTc1C+0uiin8kS0awT57o5Cpki3lKDLXFV
7w2wcUiXp7xjNU1j/lTGiumS8tOCO82+OqP0SO4S4Ba64z9Nh9Joy0F8v08N/b6J
nUdvomKH4ebHU7/Zat6YVzjt5PuYF4+lqwCDm+njlUc9i2y42GrB1evqWQ24qAQT
SPN2lhXoEuEMomDgjT3NyKImrkrRyQfzstby6fzJuX1BWTwJMUEezOwYixpIMkbG
VFWnSTPYgeqgxqf0iuXLdHPT1ffGkCboBNZV/EHf8OtirHZRT41u17oSJh1apYGx
3DG4pdLpPHXC/EUg/rE/Fv47eswEvf7+zhT5GQYMql0CgvZezGD3uu1M9h/tawgS
gfZbGNqQg6QhSrCkbPsdApDS4KjxgP8K46W22x9h9gCtV03FmTBkkpLT6VVTNoGa
i7cgM9JhhSPNIfxIMtnYu4TiOP23BcUxhDi91lMgSQHIbuBqRO4oCtOlheNuGwsT
f659wwsvbQJeuk/utmrkAYj0Hvsx83Uu/WRK4v7QNItU5gsmCwR/+BDSqJy4Dapd
3pvxpAmowABCbIonkd6W3RzRInVQgtq+no08EhvjEDeZJ/51InalMnolosEVBDpQ
9MW5JjHaBb7HK3l5iksADSltbVEP93KfIikPDEc281600dFL1uuDycHe+hgh70WF
CT7bjQzyB5HUtlc3pXX5LqQ2nR3D8ArHMZm5wYlD+89Mee+DKRYQOypK6yNbTSoJ
v8n9SYaK35VjAO3IfgMnuSZ8K2VYJmes5zxPPGHGxo7OvrAlTfypWO99VeTbwQoo
rkpLoc5yM3sY6zHUpYA9Rmonoalip5a36MuJLQ2POQBN82IyKZqbjM2UoJD4076t
VG+ngP01JIG1Gpzz60QpzSmRt1MjFptb3HxRCdfgWM6ER2OmQXGdhzrcfbvakgQj
BxB6J8Ic3N66DIQYP2o7kl8dXhir51JQwCifXKPiotv83t2XYXIAzMH7Fgl5IOI6
dW1feGaksy0ydEzL91IhFQlcDHlW1fX1kXzH5MgmrnJ+LQrFWmB4gNwburt0BOqZ
wyd6ev/+cliGBFlmabFD6r+TZ9fULfL7t6NKpWUd5thyMa5Gyg+9zED2LbgB9kP6
K4aNGqqGiqhhX8ZZabgoy5sumQTD1iXIVBAWYcuJofQ5jiU04AA1YeA6eDPlnilU
ybTOfF73hBq+x24alSDnehoBG7yOemLUN02Dfskmtv4Fq1QrbZxlAmGHILCt+Ipn
4yxVaCBKYQ4IIqKeGMG33jLufnrqJWq5TDvkIyJVFCJ+v6H1Jqr/pYqaFVvnVnbG
GnNVy7bXyNEEBkM5t39V8qGHepwtOwkzCyFYPzoO39zTrZCtrgpxn9eCqrpILQmA
FGMrQ0dQnlKmfKUuban+A1r/USNrE7MfLQRNlcX370JS6am84ThmNDeWv2bs13C+
Q8uc9NQ/NUQJKcNQhPs+sKVuzTu1WTQmMhzHdWr0QQUmNdV1sFOBsG5e+NuSyg1a
ChiOMxkzxpRLr2R60U62bqWZEGzX15oYNgsUm5au4e0EF6JTFAycZcqslsnQ9m94
fHdcAoaVJnbm20ULdogj9x7pcF/kHDHlIaeFZYKSbASB0HZ0BvUSlPGdUbKStsoP
mC9TwYUDREo5j/UpvoCPyPWdvj93WxZ2xehlaBdQJO0YtCHQDYYzqNOL3JxLKK/3
tDu4QHtZC5SVT0caX5h+8caYjOi+B5FeYdhxrDW93Q9vDaoWKNfkb2IUzY4J/Foy
4icfl3SbIk6XiNVczo0EDugMIjTOWxgX86Md62nKIsk2OXbbYEtEAWhpdUV7gpYB
SzVFPr6y0dqx/Jex74DElnLvmtvai2O+YR3ywyRnXvUy9QTbcYPtVt0hi5KQafn8
fvfu7/aBFn4ioTQpnaBwd/Qp+nOC/MhwidqFSGo+B83ygzrgeyZXey5EWYkOu47c
Vp4krRFIt3XoduNytD4ttm8VZJ0Gx1LAX5GB6gP/b9oJBQ0X3ce+hs/+yjHn+NoZ
xgEL1OpS2LpCUmcSWtg5Yd30u/xE45ifqjniu0HilSBZME9jVrcbO2MXovKwxCOQ
8v9CvZozZTEcbV7Th6uhyyr7VzbneFAJpl+of5+sklgQ+AYc88WmrrIXjhMjp8At
SUmZnvPaQ1nV03vJ9yXJfJlnkrCf0+yi8hEEYkLy+nZ05D34aPLN4/xdDQqRPbq0
tE3o5TiHQilYiWmdNEdo/4P9mllQht3/pCkHGanmrcs55HPWcjeDKEUTDUZURRnr
WpaCWd0up6iW/0SPYZSD56GQojGp+nwLwkP5iLUauy7BjLsYKfkSGNAHcgYw3ulH
IqJWDgfR2/eTLI/zPQwhXMrToyyUeNHWuiSHSRyi+9WoLjbA09BSx2eyLYvrZSX2
EolNEbLYYjeLeihVDM588TSx0x/iNd42rHJ6LPdiW1N/rYnwpdyXWG/gnkLmrLy+
xSlFT9wuYsKYxO+XOh9JeKOXAn+QlwUHP4vbEv3/MLFOxKCDxhLPeduconhPcBuB
u360/56cmk/JIljWdBibhzxD233K4jO2h+gD/N97KDcjMJG9ORfwhKD3AhSGdSzh
sNvDLbrqgIWoadPcSOcBlDaTQACK0HIuHh6uZ84y847Sge7cLdArX7szp8wljrUh
h0lJsngMvMAUXknHLa4bkqRxJ9qjucmXJsziplwHPuCeqZWGFvWCNhzlCoxwBZfB
Ja90zxgo18Dyuovmsbbl6BhgFRumKDGK9/tAzSIG5lG95VUCWp8I0S2/TX/w/VK8
m2R2AHlwB4QUhBCb7aUW2EJFzCc6+xusm1FdY1epDBkzF791BOD0poGSX42pyoh6
GO4d30EYWivZiKAvcd5O0MeqdUIUsZrhla/jD49+3Oe1VUBrsqMif6gyfMO3KLRM
bNO/hIUuaGbUCLTjU1SII16ZZaoQcPIRdByYdpIF1CtgkCTjdznIQX9g60i7n8Mj
BQGDcDiu0f8xuvWQuhnc6sjdiHfqGfDIyCR0tyycZ4N06ZX0UNsXWP/Q/XswhVoY
AU1C3FZh7BhGrjNnktf5Qln+eldFVp6Cc3omuAetXu83f4uWgjG6T0dRbqo8L722
FOnwsjP9r5nmxPnYvX2izpcrfe0WB9AvmxrRMJmXSohpIF6lpKTq65IWOV88O/gQ
gdvniJXDi11tr5UulxswbN/g6qczgft0AgUkYJOExjj00NehNyuUIjeMuPrMZayC
3GhV4IWtoelACKUUg8zr0rFHX9U23KVrTOviRB8E/dzjrvKZ3U7HQc0QeEJVeS9Z
MlYgawEcDT19Ll4d7xhQRT/QUbO3qg1gi3ZplEw7UcXmVvLHRwV6/jAK25YMG0r7
+mE+nG6G6rzfi4hs0zwTt18F9BL7YsCsvVTUmpozuBap+o4AwVUhERKz2x8LRi7i
Weusv20nk0GiuMwx9GH29rdS9EKO3c5ktvJb7jlcAbNE0tBw+/Br/uxkjk76ht2R
7eQ1Sj88Gv5nQueHHQLQRCq2rvRzU8nqS86Dvy2U+hYjoGGgDdO1zX5iALWwV7b7
nUVN+stgCw1eI2iagvbGwYrQEl9IdttN4MptYauUB6dDsAkjgJyA+jKSq8V7GkZG
qhEyvI0edcFQQVDd4qhOU5357BHaEsMwK9z8Y9VVDvm9a4YSXVfldaESdgTCLta+
GkFu058SEciJFytotTZwjdcdLTupfgD5I8SnXilxOb7KOaefPHeXiTZSQI25Ra2T
Hry4axqGzzahIbo0QzGLn67mkFmFcXvBgmfUQFhGeBvl74Tfunsg4Fx4FA24sSsN
KUguM0iNSzDZV/6pKXJlOpcudCQz6QsZB3OHedNloa1BGV06h/qgqoHrqEG0v3Ok
z/mAVeZsxzx30+++3H5aTokogyBbhe2A1iDaRLChuPoEaDT4bXmrccYz2tkvGqkN
98k+/IsznLyFZO/jjdGWX1f+PkoSNJDAeNXOp0QwaZY6uj5ZOPOIuTbrhC7AWX1J
FKzrLDnJudDENRtZP163I4EyKGVBUgOAU4cqtZBQzP7YjEwLw+E5ZbgzTJwj2HYJ
TrrFxEieOW6rONFhk2CpveW2sMrBlm9aM2V+j13ENwTHy/a4cZ4sNKpK+bLt9/zr
ueV2xkkZKdPsJCDBW9MP8AJprl2MtnUyOIYA5qAaW3thEs5cw1WTOH1VrBhhKG3s
fq2xiD6JzE52ux2wLbCiK6DiMQOKGm7aGCbQAzewPupoHjm5+EPG8ZUJWhaV106s
fD/78XM+5XlzM1M4NqnHkrV5i+r/9Pzy0qDVcYZEciEdfCnzfq9WtD2bosR1loeN
uQLp7V+WxEs7c6jG9vNO4Pwq0JFDp2Ssddlqwp7jD8DEGtbQeD3Q/ZTAfVI7iqnF
AV3SPE6dKQ4YiPUbPKHh1nVtESkFUmbdhH6zuAaTPxQ/VxpRjfA0R/7x/Zug/1np
Vujd+aFlQoiyCDVlFFF9lcwwrwMLFzgBhHx8dBhT9xqUVh25HoC/09Yy0qHnyYHV
1Am0CPICIg8xXKWc2X18mifqLxhVq7TQtkiWFTTBTIVGl7pQdimbhNsLwkyhnrFi
Qga8cx+4Br04uqUcS1XSCAz0Pr9ooBnEytamVXRtUwmrb4/LQciX+zwnkWbhUUGC
pF51Wi9+5yuvQKnvjJiOykO4nkZIoNGcpPdP7QbX4AzjozwjUNX5BvVTdWJ98oMf
b2H51zZ8NVt+wVbLKNH09gCX+hBtMpAu7qsmvI+21PWi9iFER5en5L6NBe5cWyn5
DMWIis8Mp20FwCnpqHVE65nvfEGQnYrLP+38mNbaOpIC01ho4aGVOS4HxCP1PQY1
9Oyu5Fk7zH+LE6Zw/sa06e3oqxFcj8C67yHwvWZ1v+88JQGZG+WvyPI+xVfnlMPY
1G+PBqiELiqP7zokXo+RzYzIvslWyE3JVATZGBp8XyXCtKueoMscXzZUE0MJaf8g
6naNl84OZi5Efq4uH9VsYC0tYJIUg8OXTRcZDhJ5U+ueTDLiVc+rTLFObzQPoW9C
dRJz3AEbTh1ZqXmmaHmeqN7auQzZfxIq3yKsdBB6+lsGYJp6yzhtdLhVzhduGTqz
LAsO1EkDkAsh8diYEcS+57/iTODLy510EQ0HvEIlIgsXE/TzSCI6nzWo0zlCtoRW
tkA2VUq5WtTzrxNOYQuVQ1nBgvcAp9DNr9Qv9nEFoWIyQk0Pazlr5OS8QGJnYiE0
t/kMycGdILg2vh2ccatCk7KHUWOuip00khumRBCYcPW4k/UTjOYGuUaGfinl+9/d
7Ah+4z39D+tLr5DVzvPp3xZyLIFuuUCPPwEM7V1kbHGqSYBp6/4fivTYG7KeDq72
CpfM/INb4+B5SYq7oLWRMdQgGJquq3/c2KVOev2vhRQL+oKGi909AEdaN525PV9y
qidP888SEdRUGkbnuy9AMHVAPhz1Cfm/p+R3iuw4OQcKDC4dqYk9pfGEIYDoXc00
PL02/7Xd6cijLvDY5gFxvCDq4UbONEX7eiDTZve/3c/1L+MTntyQxgRbLt5bQ24i
mU1tSU1CG9x4nlcc3WdDJX1BRKLNe6xVmzH/V7xQwiGFY3/M0SOJa1xwJsEAqucp
9b4DL4LUeLDEms2spvxbAxMvO/PRc+t7FaOYsabZqe11kbyPgyadQqzUhRIh44O+
OoIKp1gup5IT2wc7H0Hkjz/ehzrggMVTrTBZeOBvX+RNcccSwvIseLi3FiFMNrBN
lC/Pgn4SVkb/DqKmTuiLf/nPJH1iWUf5pZ7FB0odxebnkbPr+fMnSXI2GzykdlJ+
r6iGAPWo2jizjwqeQDTQ9s0Cg164Kvw3RX2z7EtqNx5kIc/9zjVk04yulrliKTcP
U/2to+5/+mTnA7Dska2ZNRsgGV4tOmmC/Ek+inVWW62nGZhOvVA0LmcG2JJhtxpR
WalCTpnt/0W4naRdO//+x3rnpSZvCr+H+0pNxP2ntUEauG85KRHxxHdNI5jzsTT+
zRMOPEQRv82WoKwKVncQBg36DIqk0U3A5gkUVFPuPqFG3YAGaG7wgBjbGjYopQmd
lrR0C9TCJD4JPfJW4cbOOHdMjDaT+0JL7R6An2jQo0qTPlqlRAIrmyOyEjXAoOIp
5uNk3tMXnMvv8TfEkRcn8DBXgcZ0MOzKHYIq2YmduMQ+QSOuxt2mJdTAvDeisFk1
caw0CEasTv9pQ2eXzK82I8VjQtezQaZIEJztLMRfb8Fuo5yqz08QuXAjchUr4gTd
0LfEloIuMoHddlLJaSHq8U8NjuR0hIA++sQOB02R0X4PRptdO+1j9K8BajWH3Q8x
6WbVr0KZHAXOHR5GjwCrGsiOnrZxF7BjjKKoHRaTUwPva0JCvQZkfHIND87NMvCn
amGcETb0tNvAqanXlMI91QeLln0x00DkBe9/UM1We3ayqVfqjYHdtb5k767gcUSQ
InBr4Nc8fxAAAOJP1yV46hf4j9MOQIL62GnbbJr3GYshZOF+R2cwUZdK55SeDnBh
ED8kAt94+XU2mleDUcvPVDYFZJwJpjVfNpTwkd65Y6tNNHFWn6f0tVmHqVQPYqc/
jxr036w910sgXMMJw2dyDwzht8heNn4mp4Z4pN6C166+IN710BKjf19dZKUOnAWv
cGNMtnSNCYaUMF3T9xToitY9Wkj855lULUuNeDfAPOdQhnWIFtiDc5pJCdUXYmsm
ap0BZmbpuca6OImf4nhY1E0On/51Yx/FKPTcn2Bz8DxW0sUybn+lvS3EuJJl83zI
MGouNlJ2qyLb6OQkfXyqC3hY4IDQMcdscKuW4AreyHYJ4aeXeJMsTbeX4j63ic7t
EZAR1ii069EYMo8kECewtQHoaFi6xkMjyxcVdlSRpDftuG9rX0q52anRZbJhbUei
a2+bLfid1d9PeLPj08Vg8yjtSroe7+K8s0DZA1t6v1P29PPNcx2SI/5dJWDWMtBf
NY+f/WIOLbkhft9R9WqTBBHMtWmfCvxuwZVvfyUAIYk/dnQYKZxHTQDY0leIND3X
ycqvvc8CYrUcc/0vCLTrbGYi19ir31oH7+gBnv+t5VLi9so3H5PDGvjF7GoE1Z6B
XSUAufRESWamWonwaG6jAFTGDnpPKjKK/GtylWdrCz63IXIiPUT/7vZFrtPJE+VC
U9Y6H8Us5UjwA9rfx5SHDr/2yC5qvD1azlPiP8cQrgENgYv7i0x+51BJZShHXH6B
o8vIp/y/gM2bZ9UR1o51g15bzaDMNsSnwizfZshTz+aiUSJnCHUrYx3H6qhmWpgu
rnmMK8sLPdrnghJc7vARIyVH0b95FspNXgSbz9TSJbT++XFh8Qsi41Hufcf1bHPL
ISnhxbogDS1qqBWA/nvj5PajljivG+OVAugEIb+oKilS0pkGV9480UbqM+jKAtUx
dA6pRIwVny0NtU15rQoyXjo1zgWjo83gvMYPvG5SdJ4cIsHQwBQ6cWMuqK9/pnv2
oomwT2TFS5iIUdBGyUdGAmMf2eF2X5feN+quK65nr18i994DbIB2Lmva2GSNAhQ6
5IUeJFQIzRBjsC57OuzwX8clYTcJyvDJsD1WTA/wrW0mN9E5NoAZ0GX7Bj0G7q4i
r+CuBU0IW7WkN3nQexrV42TRxbYqWrbW9D0b/i8UmYakRDM9uRVW7d5w3Kz8rwU7
I/KrfQDBkwWJxVT+nsziqz/aDFhDnmFivfPIXJsLEk5LOsmMVs+YZJI5G8zU/lCd
BH9TpugxFcqmM5HRctue+v1vMJfUbjUImbY97aOzplhSi4ecBw4mFiJmIrPFLvXr
iKSoSUBwuI8XvRoLQddzlejC8CO7QTABaZwF8PuXn94PYzCk+Lk8zG/k0gxb938+
FKeFBMrbsJKIKw4OshcH2nPT/kZQ6WWILWQ3p2dWO6LUY9a+cEo6Wn2rR47YerG8
lJvX9ulE2UlLJI86qFEe4Yp0WIDRqTGQUpWsC2w8TTyyTtrrU0PKZij6ATrK5yCX
p4QecxotH2U02jOap9YqNHqDCDT71kJB2zXnjVR47XFZme17jIXhGF9m7RRtJ/dM
tpxfoV2NDYO49QUPzKoAwSsUDeRMd9qGf/da6c3o1DfJAiRbhGqvmEoGNpeobxtc
9cdVAnZOQXbiHQQBEp6an4PQfftIYRIV1c4Pxgofn9tB0ERCD/8D0atAumM5kl/Q
w//f10UlYlEotX06+129hsOhscMPjVMLxwRtJn/1IEbAFmFQWhfy6FsrreQrJM6P
dKUXXNCJFqU1211rFlV8dBnFiKm/VFYmGRYI8aXKX/RbB0V3WnsASIP8fbcMgQf3
PCwooPJTotkYM9lyYqFqYQym2NIyNmeBYKsw/AX+CCvRCdcjHeY3MkRX4SGvyhwB
kGD++DGifaKZo5pqyj3I8R2vQR+zrnbsWzmHaN3miwymD+4Sv9nIaHn7MxtSq1/A
Q+SUTYNdEMENRDJLloaKGR5RFhoQTxGNeIrCYyuPm3ubK6/+HaAQyXgV+nUJSo5R
U3Yz5gHXlwe5pVpMngLGHioidOW+2cVXDptm052GL5Mioe+zrx8E2ZJuKyKhpHcN
Thcwhym2mOJ2T24kz/qY7ipDB1HGZTsGUzZEuqteNKll1YFHJd1lQI3WhyKP2fym
pVrwhSjE8GJFTRJaLoj727GnVqXswaF09gbSnkBiK0Uf0sEI0foh51B78aRc3OjZ
0bFUEYkyeE0VuZP7OT0PjAPGyGIVXcj/7HOfSXU0coMbLGU8w2w5pShl1F0l/Vax
mqKbXdo8xUAdX1wio5DJjCZ2OmdGRheA+aQzqybPvBu55thlYmYvP03Gm6BXTtqd
5oRito3VubeCVXHQfi01prMqWjTWwLT+kyPIPJMLII9he0MbidyFomaFhl2r+Aap
SY1Wl+xxb6dGyb7NmSBjtjGIAgOoJnH7NtkdvgPB8T+7FP3n7dzHENkb7As3l1Ts
76+VfW15hQQn4ZmgkInwcHnqM/UuYqs7pwOCbq2lrKaREIylk1xussEdkhfFAT51
shmSZikuV+FIM32xF+81694cOgZFEwmznuj5NiyIHw2q1IHq0wdQcQ8zBElqwfaR
yFsjrRJbAvnWurBLs0JoVuA8G5OOnIU8IgZ3R2oex5z9YkeK3/kXlI2BWPfpORuR
JpZeOMv1+7+Oea4pINraCgCFLzPYHHJoyhUIZxruk934Owl20aGdMNB6AsoSkgZ3
Ij+h7PVwzuCtwhXvY4pfrK8t3EXHCXVzZdF+jsV1zsp9OKWRcwwEpABaKKyr+0Cf
R1sOiIq79BGx8GwPt5+bJWbaWqJlTeRdj448rNbsSmI4XCQ7sDeZgR6Qri8BhWXq
QS90Uy26fUHb7oGLRIWIpj+DXAfvoA53sNrzwz0QsByx1pXQFCMcxcYw42/FokWR
GAQ3dBveVN0TcM+mSRiyxXfRwKutAjllhEiZmnexysuL2Uby4jC7jwOllZ4tCOvQ
fAZS1scwzdZNTDwZ1eDHwfAMmIe9L6KsKqt509FYugBdT4AZm/4WDCpFP0ktxLDT
fNot/BpyfVsgqG5Rcfq1m/o5+beq5/VdAkDABrv0Q+iWrCJ4KM6TKl4+Y3am8N36
WBcwrSdIxbpV8DWequnqFbudsLOoU26PKmRYEeQrzByiER6ZcFx2qhIqaus1ZhHn
mkNkKLtbQaSe26HQ6UuD88W2luKy/BiRLjbZw6LvBYdoevy4+Cucaa07lMBDq7yU
IxB0wuuakZKg5Km3/QUIMAqc43JO6nF/MXy85HHg/zqUZzbkBXTrRzIw1SRyRNL2
7l8JPvN0YPglAfAwpScy6opFfWJN7fX93P3qxSQvvfpkb8C+EgKK1oDVnEIYO5G/
SZf+nabiaZ+RDD9S7gCaRE7UHATxklgw+Sav2YStwYGrV5KkS5UXnypnbGEGq9D0
0euOuxnzTzCRfNj7Es2w98B4jMSjOcuuSGmVLmipyjDHZXvgxApue1tNw6SI7YUR
+lZi5Fic6XA11Qk6yvcsYep6+gXG35De+9J0Q1/ksh4cI/w8WEF34u7PoVma55W1
pYWdS2/QgyGxMz+vzIKvSWaXE8Pp62hJnSWI6Qi8Xwxl2px4GEzGjdXaMjvMw77b
UpFRQSM+jnI84GaXDch0I3wyjgjAyBEKb+GbgYxJYVVJOPZVCn9qUL6YRwG1hjDD
Puw3fraomXwak08YMvPF7PeUHJDfrhEWPKcPEUBJd0ij6h56XfnCgtuqdPbvAKLq
PQI0MrPPOppmodPmjP5Rp+/4jJLHalXjH+gYFcGsuwzXNRKyaE+PDCa6Z9BqKVqi
QbxkLbdwRlPHuu7nfcvF317w7HX0EWR4vC+X2hc8Yatl1Vrem4mrguLJ+Hs8S4QI
AwFdW/esvNO0COaCwb1eTVvPjXpQiGjph9Ae2DsyQ/yS//EzBQ46LZ6g8ASGpwXl
tL9t7f630lYm57Nay4qQVEqsoqsbkD0w0D5RAl5t5KhP5m01ejvPntYSPSUiKrAY
XlrejvTzMSu8/zvnWdUNnBqSI8nqZyzdLr0M4c8KZdfDM5Op7HAs0Sg536RIsL6x
na0OUrHoYi4lHnrSEeokeLoY/QXnhWNPQyS8cl89knmqokYOn2Uv+JfhDtnxtPfs
yHKkhWeA5Sig/QSnDYLbfk5AbZ/u4B5M9PuCo5Lo45E5087ynhWj3SnjHXsHKLqF
Y7WqJFqaXZFavdmntOS3c7D12K7qa9EUwrD5VkF1ng26hI3TXlVTDdkOnXN8JXqS
VQE4qZFH9fj8H85o6caVOSoXrs+7Wrx0tOICSDK9dcXbf4PNA9/O04rWig2wzncW
2IOPjusOxbHXxw5vdNQ7lH5D6v7i3Yq3uqWJGdOLOuqff3mg5CTZgAY9FvSO9mpA
PYGGXu94axKVmNrgB1Y0ac812OHSHF4GoKpBXDSKL+CE78bzWYtymamt/vENB2y0
8CxH6ufNnLMTKd/1dsWhC3+McgEo8EfaMuq16G9Zos8foKsIbx2yhZMfIummT00p
bBzN0ts9dY4eIusTNkqToQYPiT93MBtEmGT71V7ocCdQMs99ZNfXUvi4untsifqZ
qWyM5JhIzZbg2mNiYLQpadczeKCGmfMSiY6n2s0kg871hMqn8g0VWwJWjlDLeXWV
juAxiScpicffwKxz1jfpc95ffEarRMbOY1/jAIQ+vD+HlNyuVCt8sM5DyZZBjkmo
fZx7C3cErESM3jPX027iAc2GwcA0G+1/vwpKLdOqyFIoxq0k5dTG5FhHUUvjHYDk
th8Dnn+Qvru/qTaME9Zx9Yd45NMQeaGzR3PciebERSIow6ji5qVeD277lIb8WZeP
ynZK0daHKhz82wmQf47IejvqlKA3mIGBo7U/rif+cRMuRiQ4wglLp4WkpqNXtSKC
Y62bZh9JqUNrLK6bgCJECM/i278RSZIKwRB28KxPUjPC73wXj96WFGhp6Y5Lnnod
60QruDpgiTqJLCIcH6S8brTgglNiKSWpRn+butwHuTcNb0asITCrEH57VwNUpXTL
GD/lyDCTqdMSvYbm+UP8eNO2OHGdUTVCm87Z+PWFxJlOir/CnhMRu/uqTtgRnC/W
PeSb5h0UHAJ7nFUjd+oV2cR1NL8wn1wNSKTXLCct9diB2gHU2LqRl4Hlvm/6R1nm
V524OdAB2JootkspL/OWZcde+FVLckYmY75rbKs5mVnXk0qnRybkgu9bzKDkwv9m
ZTM8vqsyNOkK9g/nzJRF9H9hng8stkd43hKDGQ2PxP9BhALVLpcvNifW3tEAPRsr
6FCShwbH2iPR5/t21suVVUFAitSlrpyHC2c1pR4sIDhdvmDcRPj1I8ywR8fecxgj
2fBacbe0rVYLV8zj5TQQK4BJOq27YvBiV/tzRsCun2LE8GklAX2xwSj8+H9xtHmJ
4fc5xMpB4BcpjFw4R/ZiOPebTo5RwVr2elrj5ip0lanBbo6hVm/2slO1VHB1Iqa6
2WODB0cs3eekkneTx1IBhLTWExIlaMuDCMvaE0psGDYAxXmljEeLKeucWqRJwJXT
QuPa7tmmqQOBPiyg0ykQmbxsNH9gVLQpKQSLOQb+8/9iEi/vYz5ScAtDoaai67Lc
MUVn/poQy8CZ+mDfrw64j1VZGA1zVkL8j/R0ti1jjGRZYSl0nUHBtvPhbKhs3HGb
+YkO+CgqbV06WWlLTGwyP/Av220Zp/7GBzez/X+cNkV0lPyi4FQ8Aq1G1Pb5aYd4
UTAh3jLfo1VKFYosFWTnKKeqmAu3gaeaW7KXdviKV9B66ugatJ8bEhxQekEPNE0N
KpRVig+9yttFNa8/rOvroN4bSZJjiObxL0WRefcmTCyhzuF3bSPrGlpQyyJV4VsO
Jha6Wl+5KLV/u5duTa9q5OoF3fPEeNx2BnqoLGTVp6rMkibh6bCQFakXg2Vu+/9S
Zxry9fBMbNkjPbuKXfTTTqO8jCytRIKvhu62VE02PDhUSNEzfxjfn7TCJHBW8fA9
zmxm7EJai1UT/Tl4nnIxfsSnDXzuwXnyZxbtMRIWd6XhRwEHCRrpoLrybgzkyFtr
joXDdpehZKwFSSRJyo4VzBajMTFZ1EQGG2V11YvG2TmUqkUyr6K0snmBWLDkZpTZ
erI34u8kScYUzFapq5phEVUMt5F4gPISFgNeeqQApyZBP72DVwWUcAQMTwdBCqtQ
ef5fb2h1SLITD//rWiKY0JT+TuH7h5HFR1XseMdg0ULnoFq8eyTyDNtjV4ObHmVB
IQmV4w6if8duA9cRYlcG7mP0fgLPCq/thHuRhX9H00x047wRn0CkTbQTxq6gjZaR
W5pm1dr005D6FZs0bXwGsxV5eJscL6xY4sMtZ2+j7e/WL2PwQK0H0CsZbQr2uwJt
V0+2V353qzOXLRW7E6t4ogCodJx60xvzSUetYlkexHK68IwqIcpwP2q7xHfxqYXZ
6OT+UYFk+ZrjwfJF45VuClezCu7ZoR0sALXYiOE+4daaGLwSIXBKrawXupmXaV0H
KN+KaNVCGFXwwoAqyE4gGVOudPHqngVyLUHXT7aqfxPrz5eI4gbYSGO0awOJT8Wq
R7vxG6PcuKdwcEGJgP5Sar8fFfcvyvJ15nNYvt0CWRnLn2Yg/K6CLXoaZuKCQwN9
HhQAAcNf4GI2mRjugpFRpnMCnBBc4Be6K2iudIvjqBi+T7sSDe7DYm9eZxIa9mIO
i1KXdfFzivllYAweBuwx8//zMmYHHZ8YfSaaJFYrX9bKYD+u9MX3bL1DZ8s5qsz2
uUVHz7MKi6qjYb6HKWFj2UUql1tuHvF8FWp2VDatfQ3R0w2MWv/ndD8BuvTTgBtc
FZx2hYh5oUTPF/s7HIFCxU0+MkmWyX6HH+FYA9V+rsMVfIxgINdWRXQ0pKbR3D8/
k8tMCmatE8wntsA6Lwz2XPkPExgnsmHe5IR3P7AmaPCGsdzEpT1e+XB7hW1NrnJG
5Rm4yIBq1o0MUNm7ISjo9H59FZnKzqxlLHEOJGXQ+v/yyd+3BS0B3h92BtyZOkh4
ls0zWYKUetvGyDbeIQKole7ZeFQjEy+G4OLdTDKG51KhzT4xVT8ZxHpOby6mv3Ts
MjmqTKdQrS/RijdhgCaCmHWCUhnqDMCl3GTXpb70N1hvXieY4vSjCrKJrIDM27sH
LlUD7EQupRGRQbWP92kswMHFPk4y6Jfft6Wy/JsJvvOoHxPJA6y9dzdfB1r2gm/6
Ia10NhaJKb5Npvvhn0gVdzK5+wlMIKI1JM+bznawPgzmcUEU5ljdEB/n+98XU3dk
2yJ2CM6s6XMIWV65otM3HPvOdm5QScE4sk2x+0XJa8Kv/9jVKF8I+Z29RTkMPefe
3jW/nwExR78RVuvHsff2pke1x10YuL+3NpmRSjMBWgxeNN7PSqi8zS0MkNXNdgf0
gQrex5GYCDgnl2XKDU+5oHy8Xc3qeSXIgPxACTvlVQOGp3V5CJkUw0yHnWbT3go8
kiD+4GoIiQ1TODO+PEnQ5N2LVQEVRxuaH7vYVecL0qFEa2xgM88AK3xDvF+tESQ+
PVzi0F+An9UoZBPMtKE6LsaAf5q1hb7mYeCju9m8s+OMJkdTeBM43bQz8L63OaPm
HRSUzX38DMpi+PdToexJr3kTWixr4kFsvYahM359GqtTgGyeguhhb4kQQOLYipwp
qRovv9sQH/AS7137KjMAezPMUVi1E5I07Y6KT6MQdOONq4L8rRHYfTmBnSa/I+la
4pDVhF6c9gVw7ZzJuOV0vmn5Md+PVGS1frEU+dowahsgJUSYvK+77APoS4jqWrcr
JuhxbeOLsQUeqVS6xIyHvKA/lkJAiCRS3NZxHWVl1JwMWajgzok1ifb4KxHnKAVM
9NMGqTxCd6emXdygxnmUJxSxpWuxU5bt7FTtH/d/ZBi+1WKbEr4WBqC3XuuLw/4J
+vsKMMVAcDRcLyHLW4MVyLMBVWf3JWjuhXhtBh3pBWK4v4GBZHuL26YHBkCIs2ps
A4jA4hNs2FM6RGL3hpBi08mesBCR5eFRBRgDJFZtoE2gLcaXyMX3K1GRC5P20JyB
ZI9vQEvUKmWXvYnBxYQdAVAcgtDUZCMJcrgXcoX1cf8OnWY5HC2FvBiWUCka+vvf
UEfWRStY3grBd1yf1ZjeZ7/3k+g9zAtlrd60gKs0CFbRhfldL3oZA1ckx7VXeT89
gg/cVvuMM35SKZ9BY0oU08Q2ebjNSFUddx+O1N3G0KAtALH6bq5iOcUZTzkjXScq
fGp9vSc6xUdx22+eXkFoRsXo28v6v9STbOFrw91fT2wPzIO1qzFAciOtAV263Jz9
Eb1weQIl3gupJHsWmHlk1ijRivqAhBOv2z///HOGYjCeWVnG0nxU3qy04caUatZx
haZ1mG8pQe4/Bly+PNJzO7fkf8tQkwizLK/ejF9fEuqs6N4ItMqhhf0eNkHlH1DJ
oEuQ0moCaTBVhc4FkMgWMQ9QOGqR1b47Mz43mkPGIZBapMs2kQY1yiSTZgHkBO/k
k0pzMTG5+okFu7TfaeHCSOTRiT4MoNAxAeLkfl3G5HDhxGoBgOrPCTUBpUtEkKmu
lh6aEenB7z357a2IhW+FAoTBSiBKT2F8WT4gzizGQ167dJ6mCMfhQTSGHAPGjC2F
/f6MW0Bph4rpQ/WQetZcwfsCjnzh9AmM8I4MIy9scpSUwvKv6/FUjNIfArO8e06c
a5Jg3eJFJ7sGNqnSP+NPFGDQcHQqJ21NIDrkgjH9NCHL4sAzZ5g0kShpoEQzv4+9
I2fupPsRFbI6dGOf9vKVKSz7zv2QxkZCvz8x0CedJ/bdBVSUprC3xCJO5gE2MgTx
e7QLTCQfG3eYWGAkRrM3p1YXfWX8QwQcO/GWckwdAmrE2pUxLA0WjYRfnluRCJf8
yHGLa1wowrl+cCJCtLj44R/XmOER1KkX3zpH9JRBAkKytDNAzh1DEsH3pFUHuSfF
TI2yRHt1eBuIZdKk3jUfSTnlyGBSIjvfvRLbCAsSlVKuj6w3q0wbiQ1t1FkUG8a/
kJCKL2VyaEZaZ+JDZ4XCftGUba7zoXFtlDlHJm3WIIQg3z+STobJPdnPgD5Yr1Dj
Uv2Ly3afTL2RtUfT42aNvFjgqHQadC1w02qwCXbxj+u2EJO00Zy+8a6ys8Nw9BOn
2lmGCaR73MUyOsHJvRtaf3/klb1tPWA3cjlf1GAOGSWQAqu3hfZK93fjrTLoad76
x10yYasvWm2ghfPhQoApQ0WY5c06eFlTLZu8s3CZayagVnetStf2M3wfDgBZDEf2
dpMTQVj9Qq/oS+BriekPh+fH5DXo+L69VD3yvcmXv1WTaADmfKNwjNog0jMZwKaU
hz/EFux0tLfErs9x/aJNWPSOgHUAmQbEnBl7JE8HPOXTF6CbVxV7gh7U2C9+5RwS
y+NlH3TVWRMQTZawRoMQY9wbbQNg2DlkjACi8BAl1t2hulPb8t+WSqFoGfXy7zoU
3jQAcXnejQUApNMnTtr9Zbu9JrkZ0uoS3bQqdNJyvmE9mJVAHPOzAp+g8R8GkcWl
h2uuz/l8Jg9iMXRAWmHkrR3MnG+zLd54ngvODCObceJgeZgjRPNXnlB2iQ5VVYgf
3Zgay36IXMMzDGsM4pgUmegv6MqSUwg1AERvA0KspW6Wh8i1OyWDa/hebRWA97/p
Jc9EzqZX18iSQ/oeH6J1QHErlAPBQTrCccdETRrAaq6/ar5zIcU3Wi9MFkipFoZ7
tXNu4TbUhUbPLrI/xufeHU5TzJv68raB/UyoOWGOQfPX+26jWxG7ukYH3RKDvnYM
F2xB19rn8nK4VYeh6p0zS/3luoj+aooN38iwbM0MQQSSp/lW8aWm1azL+2J2Dwo6
6V08gRtW4rTVGFFg9Je6txSGb0XjVL0mgb2Tq2YTX4lBXHIW7BGhMlJO2CUQbbgp
h8YRZxvDh1M/TMhAofl1VUf9zNB/QKYN3O33n1b6tlfsQXrjiaIC7vpALVBrToSx
5tF6WZ4HMrM35oq7/rrYq8K9pdlrdSwnRCQHzjOiPeZQYxIDZX8HTPJsRIHsd7S8
peR5xG55Lmgfv0q3vj5X7jN9IO2eaZ5LSoTSv2jsj+BvqgvqCyrZJJo/pdKcqzDK
mCvpSHv3b8Csz+47C5cV+wUwaO8seAdS8meDjez5S+g3vxyrkZPD+2+NmDKG/vO1
pm+ScI/j52+DJW9hZHp3IWhiTPzWf3R/t5yMrbvV29kIn9sH6G8eShjezXC+TuSt
cNdr+ZuOd+m+ZXyXiMrk6TqlBzv7RUrngaG33ad2umn6dCyeSQgjAJxBJaUVPhcP
274/VF6xBtAMhOEoeemUnoVQ2U10w+hB9J8JUWOjTPDiw8T36U5IMA2ER4LmZbzn
94XC1Rac1jPLbSOkPSgSIyVqG3GxqKom+wyhmeBVAUbtKUZYA5zbjXq0VFqkjAL5
Y45MGnsoIiiKdJS8kf2w90TYe/m49FocE+WTEJ8aRen/16DM+XoW8g7S3f1MUUbn
xhR4WaFyNpB7nyxVMNmkFZvXU5gSnrb6rLdhyek7Bpgfiqhgb1thcWKeZO/QiNJX
oulacWRvRhTb46W/vZBXXSARit5l4Uky0umB8FZ7YrOM3yTaV1bF1Ie3Q34XZiuq
G+MUphRZ2E1G9M3e42shNXGvqUDdjKzpQNmme3KNmqu7UR+1EHVB4hq1be424olq
mVS1JZis67D8Zc6V4U9NSSwoQgSIfzviaWBMRi1mz3NzyC1xLnbcI8wBMdtFjBwz
wqmS0MPtD40jqS7f4c01LWsaAc4oVtuaMlgrbKKcUguUC4dbrtneGltTqIlaScMF
cClU7IzxmxYw+ak3ZTGFBssOU1dxGJozRhAnhvTzumPnKHn4qPapmE1kvmeDfJ7Q
fTZzQpqvNo7RLkhqjCpkvxZk0h/sYqT0nwFXl8J044blW6pVBhIgTGSdmh7RSEyE
WjUrp0DyZbliUfHcCg/AUxftq4Y1xfCN3nhshsRKNxM+J8epZqCGVZqWyzLHArrc
Uts250fyQ5XXv6bsYewatwnGwyKudyywBwf5OZb76o+ibOB2pskb+7VNej/G1A2d
L7RLxN/ffO7WDmewNjUZbJBDwY9eHsxW3qTTNcG+ZneOQfI3obtSuYm3OmJVrKp3
Pno4Q5sRxNYyImNnZ8aXqProBm0UfkhZVvvR7d3CIGtOyRk41OKEP6OLHlhIDig7
9U8Y9kbMJCRRmrqnWeKWQMbmAvP8CdXfNufKdP33ylZPISzXhwaSLq+103ev5N8N
QJdakWmGCPSsY1xYi151peiM1zETAlqwVRcA77cUHgz0mBVD+ob2xMQVLyHUGOU/
4kLuzGKuGno3WyHBkTIQWDlIot5C/gh8DCttqzSy4inEfUzmjevOqvuXqefGmp9V
kPvCEl98kFB5M4ErZQxjgbFobE0/qwnjVp116c+L+lYwndnhGG+YFQbAfZ0G2bEA
2qLvh1wzePf0YGM1sODlbrkGvYGViSS4F/rnU5dBzyygfx41gD6JRuPK+J9P0Mtf
dPhnfZQplAt6ykc0R1v1ZD0s7FBFIColNC3nIXnt0EE2F4cC7RIB1KE6RD6/q29M
78ta1XTTvBClXj9moeo9pf7jUtiVlOrWZx4336pLFU1kAUcmp7E+G/8mxzDivt4J
wsZhqxWWyx5WgsuJZVYQ/E6X3bpOhY6me3CubM0MYWyTyDLVXp9QSL0Hn66zQ062
E+KxhY6z7xJLRu/kVxBKd32nf05pynDZ40c3uh9KeDscqA6TWfy3JcvVue51yjCN
3nBg8xrPZ/xGPie1LLVPq09kiGfiMXKNqFfo0VZYgq9WEPZihCzyWOaVw+KGMs/s
s5QMN1uiC+2TNqDEmLIBsoVfyU5YjuBdA9g+o4+LaRmpGGoidFyuDuWgDghvyP/7
+QH+Q6QmpR8WFLwnWdl4+ZVwkIHuYUHCpiOSnOkJB0XWCNW9Dx6sUVcegZQ8J+lv
I93lIU5YapTBHBus91Z/XwlHM5pXGKmnCF5Ea6kbvxzHZATVfYao0TtiWk7Mzq6B
Lo9BUBJSwjtAuyRcUdtDxHAXNZpfNnRMGMxmOBo0DvUxCosAjcxeMDpRECp5q71l
wHGOPDsWoAJhNQfatHziWO5WnngFVBRzg25TePYOmFU0jrlDPbEmSvQoDeRRB1jG
7hGprNMSg+qty9CP0a8G7qd1smS+OtHZukJmwTQQ5LIYrTFiqa6scwRL4D97q6cw
1a6yGQCf4I//S9VIvzWDOY5c/ClDiJvC2C/xYMUG78RuLaNhaTCbLgRYVSnPhQAv
idviqGOU7Hk8fwcox07KzPqbHVnYLokyJz26LTTr55NlSxBGnokoHmmXUJmydHGX
4F7vkPpk7joQBjA4YMmbaH96/NXyGOGSpqV2jaN+TrYzMBOTjN9NyhmbhXOQ+Aem
7ZRJyxBblH2j4DvBa4KJ90n2qyVEIGK5AZZMYrTTnffJ5A5Z0c9xUYFtHJvkF6aB
IOES3u1fAX5G32JqUy2gkyQWGRUNS3A70p8hpezXGbChNGacGIJ5rv7JTWrVvDdW
ZcuKN2TpWVxh/0UfFda/+SKj8ZP5a0P78iB7bnLx3h5PnlbiLueNsOUyCkD2Bgnt
gFjfhIhkcDwWl7YFH8JNfBgRAFqgGYPduYHXSqFiwVwvzaVQ8IHOdMCu9SLOLvlP
/lvvHOa/DfuU/3XSaGEa7T72bVyE3IJ3MLG5hX7K2SQbBF11w3+SfIxBXFANQQIu
AohUHrVMaWrBypa3Qf2tijlgRyTrxVUGdrD7qyZeiMXmVD1wO8+JlG/Zxs4le4k3
kdly5WYM7cOTiq6YiQpItiNGRcxe8R2QTzqYQfu78CYOgCU2tVWIxjvIAym57iHR
w6zdqsQb8T/xDnm7gyWpQhKth+DCtXPAcacZ3CeFh3u30VtbJUeagsoqZBVk9yWN
Pi3/Snn/xVi/fI02AoLjUUTqS96ejvBkWQYikFZC3boa4K5yY9VJu7UUSyIBBB4t
+hZqYvYKtD3/aTaA4diWDKTKpL/xOqDwiuXeOf8BNu1hvN/cvNQfkHMmtj/M7r1Z
rdcr2+tV4VxldEWBY4GH20o1absYf6nFWc+j5QKfiZW7EVeT9owwmnY22mF636Mp
jwtOcFgLyRbjFP5udI9MeJlE3TVrmNUf9KiV3ORYU1omrloD1vGF0axVDIZ6JzLG
LnsVhfgTowKpOUMSITy4f+Y10sQEkExtbBT81vKMnnksSsjZw74CefODHUm2NwMd
G0jFFqTpcytMYd+jt409srEp53CZYs2IJkT7MDBRwHBes7R+STS2z2qWtL9K01qS
pHSeRm4idEj+3XFqaLN5sWdvXnKG7FTgKNe9P/k/2d0dTgUnubXZk9LI4UEaFwXE
JT7h4KJcj8qKazhQhazDcm/W6Ktr3ycbR6Jw+I6+bixjnYm+iIrm7yTNlckAzNNs
ZyUy+yJSo3YDcc3nKWbQEu4livkqQmzFZ++6D1lcRL6AywviLY8jWIQwrTj5k2tb
ktwje7C3/2l+rL3zMltarUhIN3xHw2ql0WyKf3XzBVg1p4ZjgrpA/3M0qb7pVYfl
9ERjSBowvDKbM8kMgv82qhfl6qFrGFhFBCHeA14jpTpZApD3he2IPGYNWWe93HiY
9nYpwZ98ytTmGo3z63MrwSExQNhQ/PMjxCUQJy5W7Jplt0gP6hFl5drBLjyYsIZs
4/hUP5mAeErDZ+rgKGRi+vBFIiQQDoKefgdaMYKk7GaRSeXbHdZxfmadk/X5HpV4
eYKa9GXcr9Q3wjgF/0OCur9dzAlFJjWkwNpL5kffy9tuOeoxwaRHj/IynvDci0QW
jZJIAJ8hjCmX//jRsU1AKe2V/Q3Jgu9K6FHuZddptpX4gT5idq7isQYVWHpNv9BE
fPj5XMC11aCu90kG5zMoQb+xYBlgcEBZn9wrCPs/bxAKEEJDrmaUkKbIby6zrkrE
NtIFezkWI2pCPTtgIH1MLMw0yU5coaNCbudScaUaStL/35Q6mAiRTjTRfEElyjmu
xkWZFuakAQLzp5C/9mGuCQ2ZwOjpdIYXFg+tWqe4R29nMvM/UNCqKuY1F0rxzV4R
9eTQVdi4LGfRpyVMKZGHW5iGCHPn7vrVQXSCYxPEmZE8WibOaqxkwKOZPkoxVhXd
MeORa7C8O6G2b3b0HSLyAeo46mvXNijELZOJaTrrAGKu8uumVUuTC4WFSAtzenSf
OioWirA1m6W82WtYBbwynMPC3VqQPd8wlLkGFqVoUFW1vcf/s4nMqm6gSEG0Wxxa
y87PKB94yZBLMJp0oX4TWtCOYSVxvRt3z06f15cEMOiGCN0QFWNpOC3anJ62s5Ls
baPihbcdfkleiZ1xkZ/YbuLhRswjINEmkMrdtTe5gPjUQc+hQYa48T/iT2DM4s87
ePWTS/xOsD4M4/7XsbNkC3CL+gn2SiTJ3AUTJxoVT6CHtgHec4IVXbEoCJ4VWokb
CgfHLGtrGPL7iIFjagXcI7Bm43DIxt1BJ5mQWu2TW4RRP89xJOo1lbNXQzPzgeW6
4sn8ww3Wcu8VM5EHsZw2qAf5wE3NHYy+EQhgyrpJaLT3njnn19hXiYy4F73Q1Qx9
+BRdsX0KNmTGVDFVknTtm2dZZxPcIzOHEuAf0KaNAbIbyDn1sdcDXI/B5afca2kz
R/ABR63gdGtJlkEu32S+6JlguV28PuvOJouxWukarpI2C5uyv/3oXqDN3tuNWXZ3
hyXeU3sWsUPwvw9gWXLoDbwLKfKx48C6VI3mLlLeSYvE81kAiHke/3f5xZLDObRN
WP9EMd2KmJ1FotYOVeozNDkAd3Z5LUY5imzfF5jUyamRDpKwO7y/dfjsE9q4+iLg
uWwy4wIYTEjobpMkVZGG/xe+4FAtXKqoHoFjC1Pz6TJCtyFBIwW81B2eIcoy8rl6
XnBYFFsk/lKDuXN8iAmpvvQlvyHGrEk/H5qxMyYAeaYMvoSqImwkC1UvIuflm8Fc
U3EtikuRDsYezviEx5p5dvkW7ra7Y6uBePXgJsjO6iPc1CAe7oVipu9cBgWOCpqT
PR0PzxHWEbCXqtN71HKamC/FKuiuNocUmEumRwHtnSuPpmra8WkDcey3p9G+BD2O
bO4uYnh/JaxzbnFnISoxP6sJ6oTYHL8uG+wdHgbOSaShGmYobJrcaPSshPBHk0lu
4OhJ47t3RODOtyNY6ETwKsk3D5/iJ/0FZzXAmFbw8NonUFQn4FNefHicinlJay99
9ZWJqRj6+z+U0GaqSwb5sssoThITPqH4Y+hdTs5IdUDDC9DLiDXv9ZEyElIc47cO
3dm+YZ8G8hCfS27nN4fkWjZ4CqFyfaa/jYP7Z4z1suQeKZtRwqSMUlTA1jlFNMfe
heCIKWWpt/HLX/HgZ8Au2VBne5poabq+9w1zGiDiAcgyrGFJxmvfG90vLNyLzu6w
neMZ3DL1yDNdkllwNVUnc8Bzwki8GX6olncn2aGVj5L/oOwUffbbyJjhAes99DmW
11u0AncrIzcichVxQ0KJdTVE4OuNVGLT41OEhKSajaXu7hz/UmoIXKNH0u+iTJ8h
6OtXgYDLQVjDiFIWi5vcbZY4WWL4/pdjVduRt6gCO7uIjX3K0YXcbarkl4x8KpPn
/F8XMYBfugKMLAyB0IAaP/t0WyzhleyNoOcZBEK45vKjqJeUw0fDaJtzxbkjlzLn
RDqK968alnsGWxOEGE9TTB6qoyf83URpNMSVjWIxkaoiEFlG9x4HtTASQSj1EJ7E
+AljavC46uHtmxs54gMJM2svaOeIeVJuOCKlpARi2vp6pdRBdMNDx+cbpM5Qoaqq
HacscMwra+OMEHijSl6qVbak9GmeEg4/FkpPl4/5S+/ytYIp+fV6hu+MGY1ju6Cl
LIdmHker8jxCbhZBU/fPxbmFZJhm4WGkEy5LuKzml7lheT0lo3r2XA5oCIVryIk/
ixbVPf8E3+VmulOfG9xOpqi6jL3CxxQ6iBceiCecj9V7Go2UgwZFoSspGDfZWfVc
vhGVBSl+CPpnNwQUCOb4lLPLGxqwSZqu3K5aoFJMTMfOiuWmtLbiPayy76leyKbc
53OWEk3rYaB+Dhe0wVOuQ1g+VewC9Eq9UovRjSILW3ZFstZ3d9nHX745ZPhXcLMN
K8GhzpgXARGDGI2ep5/Z0Aj1WBDfnDTiM6x9PtSnqMpBxes89lyeajmVqOUjCokr
7diho+Ykd9UzrH/MwYzk+dAITA73XxWHXudKfePonf+86ox415ODkpFB+Svb/8fp
LH3RpasfXrIkHA8Am2+8B8ApitPFAOq3ANkAMK/A/GaRgWDVCE93ZzY9yg9b6vsl
IUlwGKsaQzV6IdKdkUmtkXrRf9S2lF/W6HwELfykeTJrecVzjQHmICK1AuhDAH9C
puj4g9ciHp+KUC+Bl0MQy9fTzMJaSX5QXUESqtW0UqmPwAqK5z71yQVLjppL39Oy
BXC4BkmM1Lj+2EyyPp3Av+I2hxLgJWfQVidzljdFqW+XigKrFOh6V2/FPLQK71Rq
gRa6UBXcdSeJPHXx8L/s4J6C0YJ/S2XFArF10tzyUOWU4a7T93kpdiBg0ZIvNff0
8SvZ4U0EJp3V+Dewze1pieFeOrn2mWfG8WdVgkd38QeXmhlQIX7S6jGx+8GZmr0+
qVxuISSNHMjloDGYES++JYos1BxUDQkGpITCkhMU0WV5oE03So1ep7UVE4W/Syfa
KuZyMEuDkTRct6sZ/PebMvvv4WMS7kT7ecJ4DUp7cDdfvJfZlkE2cJtSNGTt3rNT
kBYfnX0OHLC6YYz62Uwg2jK1xZf3SUxkYrVaK4+T8dkUEUzI83CJFxMjvhtqgFCr
bkvUJAxTl3vD8nk0KeVuH9eVh7lUqvA0dj5/tSbSJk6fyuBK3uIi0Fggb+4wjVHv
B76sEV8OK2ePFgeEYS7HupaMKNv3vtwBELC43LU1RxokmGrnj+j53+9AKpx2FOuY
dh91lnXH3NBl4u5QNFarx1WmcvLOeLHBFZiWCYYV6WSO+194ENvHnm0Snl6SIiKR
2s/Baa/tbu33fW0exWQcKG6A7354q6MVXyvl6hA6v3KXWyl4XXA1j2zdy6pvIi9N
Twzl3hmdLPIgWDvbaAWxz1/RYQVdC5AV7nMkW6vaHPhViA0P3PNoZirc5gGEARzl
UDFIfnyoyQik6mf3gc/XuuS69ZNS42ArsRYUoKR4aXg/L0ZDYDi3hbSWXbvRx5Rc
IGMJstMMQtgYhGQgUOPlxIRLgRvOiS9PO1IptEwJdkY4BIBMlvKwLVwl7fNNtUxv
vhlsL1LPsgiBheSFEQuD9ZX9r2Eo0oWY5tuI8dmyEfTcjKa2ChYreY0S6oRfdNkO
W9mauU8H7mZ2NbH1fjWVquNT/U7RR860eoZtAzHKqP6Uv06gH+WbzqHW/sh1zWJN
zsskiRYxYNuvca3ejCgQxr1GyELV/33j2xwTqR2YtBNfOQAQlTz/8Bm8LfGoazAF
I6lce9+cLJQ4O0OgMWYugu9sU+RTmVydqdcK2P3QGLS+c+n5qoFBtF7G933gBqKB
Vkw1QbN8+4RnDmr1XZQNgpKR9tP5S3S4m7lloghVmfjyJPn+1EmIxXpNS2SdcN23
EEtDHg6G5rLkB+KYxfRH4M/5dTuljU79aLQb0NNR6V3JXFsq3vNTy2lkn65AqZOU
8CNm9MetBxmjx3xbGad3dkZqw7dJ8nLiS66nGbTY4+HHQZRMcDwqJhjTbud+MwiQ
c4zyQnGwsT0ukCgBa7SPAZFRGLOHnwyrp+IVoIaKeqWSPGmO6Kq5tBimR1cY8XvZ
Biu2az10PPAAVVAYyW+Ks+8j7tLJAy0O+WrW7nyOgN251M28k6yBpYMYDLkvAlH3
fFls70FFGw9PjVTSHdZRTOJ9OEPktjla58jemDLdzux7to+MeT3dLf7od1Wf/iIB
T2OPiFi9lLh46/xOcCUXyvu74MOAVk3nk9dfydo3QOLFCghUsObp5G/HMCJt8adP
0JIlhJzwYuh/F2fDWz6B72ofHd7AFrjx/ndkc9wKub8Ny8bThvxwNesSQM40bA7I
ZiLu9BE0sY3X2+1IhWoF8GwxXNBMriiXbKKmebYsDWCesja5gB03hKkY6W2vhhRA
gpmtgYk0PXgybj8uf5K7i06uN1iQofpvLrkXSFJpDFqFygZ2n5QjZLOf7D7r/emI
8TaGVLddrHDN6DUhkxtXHGc4T5CrL698ByMJQvJXIe2miKxOokBtzcE8ny0206oj
Si2Js3rJfW1R778x4L1E9TeZbq+FBGpYwGLuw4Bt+4XLQjqqR8LYTQNJKuU1ebGY
kXgB4ruVcoiAwOK7NXpLIQSbcBlS2Nw1+zjf2FPgqLMgxN97G8HbAikTTnJrfE9p
P8Nptr+oPwDL9mczjOaVzgJrjVwTGEcidB7gn/saJVTHB9fMQx5Q7HXoNG8Gqlvz
r7k3Pvibkrzip237Xy/JyD66LRLM41O4bZ222SB/BLWX3XPGewqORvsHT4+FRd4b
VWl6CgbtCDiYfEjEigbwAhbjFcOrdv5hlUaWfNVppYMw8JE/kbKy1ufMgCLSRBHj
XLE/8SaRtzs/Ln/TEYVjwz8hXhuS7SokD5yYOGjy5t+3wAx0NJUhLDuthRebLZx1
DdI+GY6OdfHcP8TmcUbxvqK0tob8exmsRVYGhGVk6jwUnA2U1HRAefKkCFDu9Li6
C2ynL9u4KvDRfvTkRBcNk+VOFDYxMoluLf2VR3Rpd/KuIYLDzLQaxrTqoS3ysSta
ELBVVh4myO1KZrkBgnKOZwyL6KpdcEuxRfvNe9C1zGb/poyWE+sufKimytVzHuDQ
Hnaz36OyGdos8DagljAkPOfpNlfjaP22JtJdFMRhe4JKHLLeF54aIq9CuPCt7u16
7XLrF/OUlMkHz/j7n5MKTDAJhbBEYdyrK+3eBoDpkxTPCFzdBrsQguHXUgSQITkS
l+8mPgrP0VhHGMlKkpKk+3claWb9A3sdbnl7KmvfXyw0Gbs5eOOA6H058wCT0aeW
/u1tX3Ifl4PlG+s5bQEaAK4HGM/2tdYbfZxLtVhZPkASmmQauUrvxnHPuO4O1DLh
YXlNAKHG8YnJ0RLjQ53kizl3EEPgVWwoY5Q0swOtbeCpskp4sId5qFfMvU2ZUg5s
jvfhKu1upkKkko1y57Nc37LrZSdqJbIW0AdHaNMHsNVtHhqEq048WsNt9dYWSJu9
DiB2cQOEYsYNyZb5ikfy+XNHdUlYBIrIGvAHLAv6fTFF1qL+It9EOjZFM5qATHQs
WhMUN3xkfiN8x1d/YfH45EFoNig1SpULIViW/LPrf5TbtcjF41lxRWThNOiD2E00
3BK1oUES0SmJ73PRRvAYkMwdrE95lNkDDUYcjwpJrWawQMtiFaQmi/Fm0yGgE5CL
eUvS1wDkB3nV/PWg6GUlE6jLEeM3QZI9qXB5zJ5KtdFOyK+CPexYY/Qf20dwAL32
p+LeL1YVoqZL0By8qUUq1FeL2onR8Z9spsndfzt21ckIfK7isnemubl5vHL910F4
hP54AEhAyZYY/ob75cFmL/sI2XU8g6gLj8o6zFCWz72Qw4RYy6ONfpS2EJto/35f
3FVDQsB615gfPNW9C4ZB8Ee9SPr+Jd668+N6Q+oWdGz/6Y5w5ggsx3KNU6rwZVgY
O3yExEHtUDaX/47HYSQEeX7SLndGcHA+YXZL0NmOF42e1MkS8Fo6eXQAVcQrsm1e
K+wcSfmHg8wK7way5gXwQJgh37cNN17h5jFkuCArObMLjRf0E3BAikOeLBpVXuWT
DWyLP4Zza/4I007iJxm2+lFx+OUWyCVYPop3hjYAu+IJ1qliAFMr3c5rIphxJt8v
LyKIh6btWZe7tY1MZP5kpXOxWyEvwCtQvfypmDqj6CZMEysW58H4xUSz+5MlJ5kM
fqicLfOqWub6MDM67Hy9QvbL41onwHKb6v6F1JW0J7E0AC5wtJWW5IdWREWK1CF5
j30+G4PRE3+0FzN9luS5qHZ8y6a6JqXk4nL4JK25uO2Cvp4VTZK9sFcCIKwykj7T
XXCIDeq0gEhFpWDvdRB/R655w2v3PGRItsKbp43XnY6xGS5WdKYDcPBA5rZLTWl0
TsF70gl3o3CsESUZgqtiZ3AaC05nLF8fq+NbEJB3MJcSzMJSklaMSw8AmGdWA8YI
kocObE8cTd5eCSjhM96rfNtTtk39DA3pQE8CZ+GtaxogSwRj/ByKm1XrU1jnttT7
uVBFXsm5gp5KZx0XdNbN3w4dc6ydNz5ni5slDcK+XTPaVNiWOHMzBkuDa6hbfHu2
3cfDWhcfZMUHmhUgTNFwAsM5CpaIOJr04zfQy1SnJrYFWg3J5fMEwbLKc3TQaL/v
aSzJOBYJjT/XUMD6ZpzYy86dOa0S+9RzFyngdiAAOwTG4PwWzN18fMhj2CB6AoKj
Es3AOf+VDyN5uhx1V9uDWHNeNQzSiMjyJk7Di8SQHnEQmqsJavlACAH4zl3kGz9t
aSmkucd23I8Tdp1fSuQB3EPp+6DnshBG0V5WxlIYJcxH4C2fkcvYX86E6yv0kXib
BWVwXDKL3UqPPkfhIecOfdz6Rg8p2cO6Cfj8zvKNp2UeERivwvg84PXWO5U46hMW
K+HDA9G9G4PJ6UHVyetnhMwBPBZh9nlzRRN+SATSM6T1jHyCrlqlu2VNfQ+luWxI
PU3QWMR0QFOHDIVaTTsIWgVhOfUBENf28dATOQB4hVzBSzmN2hdC9vJSo2V+Vsc2
d71QQ9j9eaR2yVKhUMZXDG3StcBPO9tVAFUhrUd1fbMSvgcKUIKGSFGisaoffdfr
x2YoW0e3PJesAoUnEeildgEmBPH/UOTUmUs3eiONHFlwl55Wo83XvoED+G4N/v0L
p+UEyJU2LH39Mp0JSZs42PjrIyhEu4miCCNt2iNiW+FbLLOCn5GhiZAIlHyLZse5
d/ptaJlLhv302OYgVkpLIYyKjjuGq8wlHi6hcsNxDRjDLQBxgAQZcChwA2XrPVxX
p5dhti8LISMI5HZKXzm95CwyiNCXF9odfMpQy9KAQYG1Qj7XwG8YXj5MgzcuJndJ
+FKWQIe26r9UrLiA7/yHKTxuySCRUAT3rXAXzJbquGQuOhgyGks3yWW9NO+ekmCk
f9ZarvYmjAlfm8H0vFT8bZgNaq/k6/DiFN+LlAWY5NnH9+EIvEenY3rzDr+9BHfC
rtshWGucucNywrDtK0suzpQaPiPd3g5zlgfv8NPIBvSnncBMJapk1BvvdKvUMTPK
VPDNimwEOEEssXZlyYuUEdvSN6tvfEpR/C8qkOwyGTHJRquq4vujaDqvq6vlkpvC
sVz1TJkHMznqRtlnfISEjZbYj0WKjugMzR+I40pfSiHXB2TzLVUUeBxCchVIuCIM
IxyaIi2FzkjQXUV1Wt9bl9PdtA1ONgJPGgIT+qnu/2Sjs/wxOE9NL4E2Zi5OpBeH
nmuJp77k0WIzExteR7APXrAvP70Ch+IntUi6NHmfGc3bkXEAe/Qty7LSVc4TfdJN
YysqxEC5k1mncNNF9/OJwcnUtILcOn73y50GhN5xx8W+VDV9GZIXWAfWD9l5gHaq
DnSqSEFD9rRhRsn9/9kLnk5dtLRwkn9zE0OupLsbzCLXPGmmMbJt5eUcd2lB6DD0
GOmCo609t3cT3nYcnUCLOVTOomSt7dU+tTMAmuirwTPokRJlOeM4s9BhHvwWOSbR
LzzwuNNfMu9eHSt9MuzMEWsmmdclFkSu6JRnS0JM0KEZNE7vKoUCiyqUhFbnCHHz
1LCjqj5+rRc8j8N+6tIoRCopKa+/D/TY6Ea5R7dH6vL0wVgSCxll0Zc8dfwiLodt
Zs3gd8YnxFhjckNfbpp+2NnJlmqME2lU5DeOt/EG1ZBuwWu/3zKDEIYeENHUcMjt
CfL548v+0E4a3lc2i0n1JmjxhLpodkUvYOsG+aF2iGd7EQ+1Mky7c9Ssrznyx0eu
MKa6tnXCPwKNKvd+KUS5KKl0iDuRT1z1HmlWxlpZp/f8J9d5cGWQnaSfPyvrrvbZ
MSF3xz70sIHljkSkI2e66SwG1Z2VJMnrqK67n0rhFZ4Ld7HCKb9p81J/pkRnZVj8
XpQ6R6Z2FeCReAgWYDfuwPBgoboGrFoDBYde8yShJCZEdADbFzzJamF5VRFbxK32
xS3ONB7uUPOgkhPF07HDDAkP31Pe+RkW1Z8FD3WV5SuEanvVNvw7BDNKgWLUViOc
ICf4BZWN2zQ+nLEayNbbGT4SLcl7MShc7KT/+e1j8Gx2TFSGEdd4AfTt7yYNl1SL
r/YFgGEQx6p3ox0oL7/wHz9LEzSjBu3aaoyYuGLhUhKdqu5z8qQ7rXKM4pAfaUJW
+LONiuEa5FmA/HlHVqPZ7zThvYRE0Y+4KWbGa4Xund+k8a1B5qc1U1S+pyr6SnlC
Hd8u9xDySs1m6E5niDzQvZLe0ldPsRzzmq/YG24giQY9krG+JaIDkNIGOWwBoe/x
SaKVnCLfPEAmrvS/sMIn60sfQ++3Viv4qNLwHgldWx3g8nIdTJJDirUOHiICzvtX
c7N6NMAoajxRz236ZndUYlvH2VhPDCAFdOoYTKuYHYPIS6oDOfqD+VLq4bDWi4cT
SwkHQLN0vjWYgLpc7SwlqQnzpqvSD2/jDUfF08kHDHLy4wzsSZp3yiPH9L747Dij
6h/b4J2QL4P93IbBBCXZDxrVVc/Zn+HhwNTRdX1GrPYW8Bq6Dx6TfDE3t0L4DGNS
JE7wmZonMYP6nXUP+ydLID+Oju3OY5d9ImBLuF5hNWUi0EW52bH0a6XlhMfkxC6z
UElg/gBmcv0WXjZ4fLFIB38/LCxtK17sVxachnVb47X0t2/VS8/+pGtzFNU0HPN5
h3quLDM3j1I4s7cJLq6hBdLcK7hk2g2dki9V4vCr9Eei4YW3MfpmOvPOf7US1gtp
lVl8ambgOhOpzKbdykpS7pBlgcYElpqBZhpX2ern7SKbMiqboOjPwXbDklIOiMzN
gGhsGGzAjm8FbcNZq6CquryIc3Eqpkx/+F3/L7tT4vPno2p5gW4+w2TGvtQZKO9v
w6UkYqkCcOpOY7yzINVDwFjBNa8v96IbJrXg7J2IyO61OjD5SkHfWEGLkng1H7x8
nc77PCaxxew3JhCBbKb0QXv/otV5J+cshBSzNIsNLP7FrPdgPewIrEAbs2gjQCrZ
QhWb4RSJgIA5vfWUloCi/kBAdZzGTtjZKZSfwZXie5nNE/FppwQ5p3kNA3y9YRkm
gcnhHWik5Cm/esDffgp7GYxWWl1Ry/pxPQOXGylWdZlRJbPLncFDC0DH8xf6puAh
oLUAV2yFxXIlCjpzKHdQi0JqJNaZUcz01rlo8g6el/jNIvkY9IgvwY5727zLxKtx
+bn0snFhTAUVGtFMZsXM6thRn/05PE90iiwABIsmMlmFyTTMI/X18clU8BPM90SU
WH4VoyOwt/mVVnU7ksCuYz0n4i7a/zLAa34T2kOMzJ4XA50k0PTO6fqTrfihgbVi
YjQiueJ3OpP6isGg107rpglKaPatG1BhspK8tPPfOGh9zeKn8UK5SIm4uPxfWg1b
n19hd8RT+GraxnpHzoZujhIRmt4StBn40d5tqUWTfYUQzG+LNWOdMJJKlSrSs3kN
odYsO5ZLNGhsfG4v3Oe87jaBjXBhn9pDNYzJ2lbZm8BeQ7OuiN5NfIfniklpbw+M
5ziPzj4beglidW5BUdi2X4IgvLZMfUyzGPoBklifrm6P1tQsEbqa3xrHKEl91HRv
aIVw+NXEJJpkof3Aul6dz+rDZOD0UOpIY1AbcpiM3XXu67omrNtaNcu6ghQv8V5A
R/XaHBmV1u8c7IzkfXo2kP+w+AI6M1M3/eZMWPEVzGRB4QiWsuWgk9xRDhxDXMVU
hOQtEHQJsOtAmYWVTO+5h5bs8dk6SuUyFdDPbdSm5Wj/O4oAxeu8m+gU6In1FYoC
LB58/Jjt9tuuerPv5voPRO2mAN7wKshjisKosKaCAsEKH1iX9HImCWDPr2Qr7EXJ
+VY8kDvf25Hre1vIxt1769Kb76gMszxKpgGIFTQmQp3DJp+l62C5rc+vB2fm30Ne
QwWPX9p6cl78WD/LgeThXGz7jfCm++uN5CV4MTCcVbNw8T22S8OJR65G+eRIcVHt
x44U6128il+x/ND3xGyk4efnzwtURVMpfncp/aE3EwIaCSBC2GmHE6iKNvWo85dd
5nxQA2XXJXQCIOSaK0gwzZb5hf1flhFsQBN7dQw6KjWAxysAXMdULZfbO9YmBVzu
rU/QEs6ZHLG0EYbHoxGn1DVs5MfL7mquiCVBRyLifYbck0mu1hoD+pRP4XTo6zbo
0csOz0WKA3PYM6Q+J/thS5F+xFYcx9u8Ui7XwpVL1/+wP+PCretIPI4X80fcsnBo
z/H5NeUhYhASVW6WPkD2wES0Hjld7VA1PMRMcFNNrkv8d+1nGwl+Xjf6KAnXDEC6
vvd0eT6VkQp8kog1s/d4zIhExphTPmNk2+rzightewfxchcgSX/8hl64tUh+GPi4
cJ9Hp8RWD6EDKHIdDTnKn5bTw+y6ZsHDH5KCdv7bY+52DzSgZcCEZG35AaYVcnSM
pBZGZ7P4X5WPRd++8C2av5PTCQ47yVJJXHJbZuY7h7uvNfppFfuSJcQ1VmlDfReJ
mkyyjsf0AhPPHjFVULXJ6NtRxcx8wIJ59M+45hpj8WgdNN4YI7kz3OUr1WdYAUZ+
74hSk22h6ZfdLzJHSm1JdnasQm8TbPPeDRmiwsoecGo4ossLdkf77scfV8CU91JK
269sYpk+WHjaffmnuc0qy0DzaODNdqfUwSl8FSevF3lgCeDlgYuGLtG208UwiCdX
YIBhXpvzhkBZniD/ysvhXy+T8jX0NJBiZMnYxJXp4GTV8aGom9nUQ3S3Q549430+
KCV4C3GQrQzML9bun1l4IOiQ74VrOUBiRv63otj2HB/VlvKHtwBNbNT+ZXK4m5hJ
LGwx3jMOrX4f3oAbGQ2QhtXpg6Er97GgNxrW5xJ6X5qL3iTkOXnKcqjp0I7TIMDC
YD0jmf+dbgSePO8YjROpEgoWQFYNpI8QKt7nMZIJ8RajY/qS01+mVGFkl5TySxF9
7thFWnUxfNbXlhDVtQvjtEwiPkYrSx32K4zygUQYU7yfOCBP4ewWE6GUEof4YsPR
xJMWyQCRq/8mhmwQgOSVYDAOGCzJf19y52E8iLi1db6b6kF+Z9FHpTr7RptYHt8E
iiLIXRgmvd5cRs3z4oPIBe8GPctlM79wdfHGVs6n4cMpB6VU4hkPAHJYv+WYi0Xk
OPi/gJroeu5/mnLLmoc1zt9/r1t6fRD3gPzstCYGO3CUUl0c7Ay3NdMZePgbMY1T
i8eGm8ltPCazgAPUOAoIDG6UiMl0hg5LC6C8a8WBnHYFGxldrIsrvGTIt6WLNaWI
901fI/2xGOWAZ9ScFk0tdswKyQ6XRahu6knyo4DyUtXn9mm9f6wkJ/tNNGTnQq6G
TAqqszWcmQ0rzC+d0Z4L9OpQA2pGsVtqphfE6O/ko0m7uYZfWuGGxyGj3/vSRNSh
tydB6D17gegHJQ+JBsnI5qZzba+n+cC5GcYBpOIiu5LvBPnctImktZPbJUAQn5ZT
nVBKZB2UgM8QlcQ+5PkXbhqo5Ye/75ottThR/miNJ7uPgVqtU29P9MLa5rRDa6DW
kH2KyACJDLbaEun+kH3D15bYetKzR3Dh7g1T83tNJVSP/7TNvQvS4eaJfdVK3huc
GdN6bBed6aCX1Cxwo9A2yJ6PMiVWSbXAgwFGZP1up8NDbTUfG9UCjoK189mgktad
OqpbH2FdhZi7Q5OZvAZB+QwnamKdDqQb8iFiZw6apgO/4ympecpP3FaqMsAIc07Y
QCa1hPOHeVv40QW/tICNceOwINlNR/JQPQg8I/GRs2Q6pFS1uG3YB4MjuCv/nb9l
wyrSGaMw9u9KJxRUezh6bIGQDa4HvLqnWuZtN4BiviQ7iQmmEz0Af4cYoshlDVeB
UZTz4TB2pBB4gTjr3UkRumxd66B7zcKGcdw4KqxbendBgpArcTJxi+c4vCWDVhIO
bsbnZlJxWhbs+c/ZEJnyUnM8YEY6NIhs1cgLk9EHbJ5VLV1jNFzsaVYW+kEbkjcq
+TG2Coie5RKAVTcJzsgrRvWzZG76yYYKzuIkvSCJlaTTTVhZSeN2vxn3TMMpI0tH
o2rKpZwLLqcYhdf1o7NSdTzVe5mXKqo5emwXYcx7bp/a1qawPzQEAjHXoiuNfo6c
v7iY3odRsf81ZZce9BOgv1de0wr/cXGEma9MwfpHFOPLuGEFjoFv2XtDlKgdg6od
ND70Zqxm/Rt3aNsIZKL8ghVQMoO2ZsGJMUPfMZah42UnRT5i84BUyUJKsauBjBHu
uoLMpwExjeKrrWcr0LUR+oL2YWss/gK3YbxGAj8yKm84mprQnLgopPYy2uL3Zt3l
9+hbqqoyGZLxH6NwuGaKAw3O6/5GiBATOtUQKwk9oL0CEJQVzrRgozUPjDPXW5k3
5dBpaOx5gWHVIUqx7kqNq74FJD9iUGMu9HybbAfwKToJdYpLZCrMwwQZBlYEBrzw
M7TbnuJkv3iRdIbIgSLZ4kj2uaN2Why3hdoDa/xE2FN95viXr893x2F2HnzLaJ/C
uYMA99wjX1OWPVXgj7fjRX/L4US8TaOmdOWi4t/97sBWYYJYBlnKMK0QVIhJgLMg
Pusxaj0iZx1wxXsVMIf5Fufx6p3tTcysVeD6b5VR3e3j+HOJWghRyUNiXn34Heix
mH9Gv3OSZG+TASDS+w/9fgCovTg4Gc5yFOm4r3ALAnU6sd77KQqAZ+bMUK0XnRgM
BjdTGOxJNcPTYuzwN5m1Ody2ViPLRwNBuMJNgXYTu28kzN2lRPHPKaXCNtrE5vHU
PbfGQFwx0fi1KvwjQdIeFU23ItfnCXwWWNfF/OI+QtoSFOzc78lsMG8jsUUH+ikb
KRAV+yRYtdQHEQZAIOPGXE2DKfnxuYXxJ0kyKksmDojmtya0/L6Xb52TlHdNVo59
jQdnf0gvjMA74h0uojNZUdeYJfBRXtmeb4RYhE6vPptZUeAARTLxZ/63uU01ijbA
maDIAhyVwWH3u+YkfD0X6RsmJjZOjvCwbuvii2/+aAGqypeLoDORffG7xN+9hNwK
LqMDXBKRcD6c7BQrZhcoSgZbB9mnlzp+n9RBlKKnlj75dFpLYLTtviLc4mj0wrp8
hq6SWM5NSPbTI/nqx3lIW1I4RYpH0RPR3o3xJYh2i2/MPEy9OXu3LnhrJBmOa1yU
NdxjpmndlPEuQB9P+zC3Ycy5dJGjldgGlOOZIxKpCLuPrLOb+0Sgl/dn3LUvH6hE
QIMi2EDOqZzJ+yEEq6Ta6wBr4H/4NgoHC+tZQUjLBi6k5upvjfM04enjRGbxIODj
/qxnzL7McYRspOEB5GsBfZ0dc4ewv/nAHbSi18KoGEciLxWFnH0ClycehY3tQnqk
YDM3CJTSMCDxeZ7sgo4Jvljw7cjPJuXUWf17cjaTfGLTXorjYiBZ4/6iLP005UoM
V+hyptDDrSMuderrdcfdvBWd6IkUywtCvuPVKLhqBXmY9e0+ICLIXyZjspXt6fR+
n72vWy4vBD0GoaubfB0uh3BpVP0lggf8bK6NKiUJif+5s0uxoePLWQ4Hoh9pYZ14
u1w6eizXQFSluU/D4En4DnhlAcbzOtBuI+veexbh6/psyz/KFger+hw5zwvS7ObO
jwMc9CtfIbGR//wsqdJBzk9aNzvaN4TFrDQ0dB6H4X/3g5DOPi75Vc/5FhLwBpGU
tgFvbAtkFZc+CEjibGgV5ZyQMZZqj3nkfhM9ZmOl6k7mImJr1J6EHg8ocIjjbp/4
jKbpyYht6RUVQAf4SW0SUmWzIFlx16PzsduCR5RPQIpwghX9POax3wkL2U4sy2Ie
giW+V6Z/ZFTNnpSJauqJlz9vb1rb5MEhELZ2jyLxiEzPczrncfVR2zMMshR4l8mY
7gwJdmjQdARmplpP2L05KCDeMRvrpghtYIt5kSHdnDNaNpf+bh5T8IXcn+DCzn0W
jnt3pXILaJ/uMYoD6tsKjELHgYG9gJLuWrhjxgh0WjM2WFWmJyutAVz7d1CZqqOD
tUC5tUVvwBD1w95dRS6Zd6pQ2HF+E4oZ+UWxpODxS5QjfxZPEhnFWhFnBSFFZkhb
cM1pj9ENUf2GvWi2xnBILnsfWRmV0Nmo15hRLuGDO/8eG6r/sU0798xgg3jltEZ/
6dIZDYHbrX7SOx3SXvQEx/q8tnKa3UKCfMb2gYEoeu14xmvQpZ22HvIGn3a8Zn0A
9ROAGBjFGtI9Tyl5wms1gh3rAwbmg7xqANbB7mnHU6liYrd4MmSBeFKLNyW7yjmY
qKwbLGdu+xG8szuhspwhGjzWEK9+pbULqjs/DuR9X34cwpwGqQYxxHgoMzq1DICC
Sxk6Qo/5M9Y0Vy8xn7CqVMdYrTnBI/QSOcmqrtORVTM6BGzCyEY/wnpptUV/F8ln
o5cGzAikL6tWbw3WEY56EUsSOz/sRFURG6RqEoUAejmaGYL9i5mp4gR/tRETESMa
joKrZiD4BwSTin1qNtvEau6D1qsmvVcrCw6NzaUyGBalmvW3HiqPt1GlMklTNVVw
cu4OhwJ1CfWqiKLNG7QK3jCi5JjAwbNJCeHIKl1cYYY+fYF3JUSFnuiykgVxhApm
jXwCtHYfaswJEKURdY10O1bVjeBX4HTnnwbKHr8kFN/Xp55e/z4Du3SxXjlT9kSW
sVqyA1mc+vPLPrRYn+anaXFqVG7BE4PgDl2GX6hAOPs6z9e49PuXlSiFFxuvQZ+4
B7V2j++4Dht5VtcUkTy79cqgoXz8Ku/bfoh8TyrbEwqg6FINoBJdOZwErlnV2FMs
76Jm9KgWvzYpazZcdH7Aka6sOnM4Wgc12kB7idy7GDLO3utjf3YDPEuk6O9Ya2YP
jEvJyHulvqyog8q6gOWSQ5JEOihzRsv63uKyHfLPnOCLw4xywSws+HVIIcNfxuyE
nc3WYCJkDH4tV5vOE8CwiOQ/zp7s31PcWqHiTIUuf5qYHktUWMf1Uku3R2tPQSPT
6YrM6JzfJG9+CKRCbPWVpXBBig1+IMbKA9l3gfw3lyIpverlKgnxL1qb5DF/CiIc
DCoM02/PBHPpM8DSwqeNk5S0ZGqTMNjDn18Mw0pD9hTQq6vgWatPklDmFQCtfB0F
qqfp3mU/kzYuTyorI9CFVMbtjISYyRx+8CNK7033uwLb+RMWRnAr1+sjMKLbzASN
dni9smNj4w2Pnslz5Y4+P7dZC07JQbwsKaADbnH7YObEx0jo0ue+nHDuouHMZheS
eP3Aa6zzEm/hbzIcCV4i0uChspMw7RbjYWSA9lyY8jGje3sudM72WuKWT6EPvXt0
91pv7ZCbEyorpHVHfVXpEfPrpo1ofkrKTTHLDfDcmDi2Idf6jbOClqSeoaWrvOQA
9avI9+aAH/YahGciYXUILyQSOl5eVGWRdhyPNC/PDn/XEIG+poiIHu8GRFw83ej8
nnWBcAhGGiLLg3QN3ppFG40UW83mqCTTV1kUwx8LkBU0bOfZ1k7iCsKFfXxl12fp
kmt2fcjrANfVyCDj8LxclHZa6TlmDkAX0cin91opSiiqfoJEBTTWqo4MtrZWKXlr
/E4FMCMKEIEJn4mCxyXL7Z1+mMh44BVJB5LyffJHJGzT063166scEQWz3cAwGJJ9
gtt2t3shrijvOAB0MkZKWgXJ8XUHWNTv5gXpdLv6y6g0JBrVobDl77y7Luu7f2aA
qb0ls4zJbVI24rIO4PfBAV0QSwsF238FD0ZZ29JlOI1d0uoTXqcb/u4fIph0qshc
KLFOb+gfPriFWvN2SY2R1IKKuigdU2M9sTwsDc8BDS4=

`pragma protect end_protected
