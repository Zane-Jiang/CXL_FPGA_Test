// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KQuv84lZulvnS9C9EM4cLHEWuwPQjtJ2C6pUUZ28I7ahIUUvrZoS0LKVgMrt6TMj
qRvsrRoG4doZbB5QSvMJ9mhuLHZ6Vk0qT4mUrJDb0fWhM5uksITUUVRy35mhBhZu
JDAGzmvp2ExOaZ5FUIG0rRxrtZK0AQBaHzamTm3QR9M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1520 )
`pragma protect data_block
eZ0rd0VZrKiZhdiQfsflXtbwBmBpc7ofBjJqS1da0b6kcaycAdm6uL5h5bT5apkN
arxlf1jz0JRfdMNavPezkMbBLEjzJMaiUegFw+AcTrc64i3rsjG3vymvKZGsOYhQ
BVoO5p/JqVWLOMj6wmkpGpI3C2yyR3SSep4+xSf3WFpbtIUmJJn5j0OM897j16ry
Q7l4u/vSb+DKHQXvf446AhkdRmg1c8amFV0v+L4TzKzAH2hPMcOYxZgqHXZjoftM
+QnU2VFaiudizMl8rzObgkzxCCwH1zQbiPp9ixxM/p4fpOGfQyZ7kinucDES6pAO
H52354T6pdFgK8dxxYBa2Qo4XyGggZZ4HcA+T1VR9LpWWnbIB/+8QtV0YQHTZmj2
nUL/8zU984PlaBcaljMXgL6U6cGWkDi+amGJeaccA1NYsOyURWpyX9dax9D4qmKv
/SSKu0k4Hf01DhUdX+RKVbtENhoCNgZafp8X8yGj58pI5Pa0Rd8OZpPI+WsLc3SO
obzjKmBT3ye/MUfHGhre8qUC6xT3yOPujWmRcVvryyiTfQFUpXsQZW1J2Iq9HC7V
uK3WGRJt4KH3nBu6z8+RIaGIQxSsa0m/nHA/BX3D2ZWuRWpdKyfbmw6KpiKaoBK3
oYwCWcwd3Gf0uuWOmkNFStMa66NdqB/TxOTHuEvIp2YaZFcSemDtwIjRxbzieTjO
JvC9wmZSLfx6+nZTGoPj+dBrn9/hYuxbzMiKSUzi2wKNn14Jkghl1i8qfjHcTwJJ
6ovPln0l6Y2mg+Y0k/PEg9ngXR5AuRz+SZ9IHrsu2kbON7JYwmyqoPgJTcSdAthm
dE4uZwB1g9mc+sQ2M/SPtu38c9UzsidC7BJ7X67CElYs6uCzhMWUEv9hTwRgeUKv
zDtKUd9dn/waGegzsTqhxopwRb8V9oX8tbPaTpLkzCkTpTp0FLCmNvITBVWU2rvS
DE3v25gXp32NTOY5qNXy4TAiIwg4I7P+PcnB9Q3Q6Qk3dHYQmtuA+V8iJGAYNGhh
Oydl8qHXGT9MQJjUw9ERmnNd9PjXrdbezXKIXRzWwQ/sTEpZrQAw2KIR6FX26OEB
TgKTsZ7VU6VY1QRbjQ0GZgrYxqTlxLagnETlUHcmJGg9OoHXbjh4wx/zpu9Y/jFf
jhLa5ZQyUEIIU2gUDt4u9Umi1pHRp/5Sjl6jP4Wpz6YKymm3IbR7gl0DXHPDWOB0
Ol1xNSEeiwKb783TrFr0bWXXWx2UhAfJJEQOigHKZT795jFnQDbWYQHvp7NRM8K7
N/TYY/rY7IbZiNLOln2J6VSTFOvJLjle4K1Syo+zuJXWF05/hBDp/LXM7eZFq1h6
KVgDeCRPY14x2uBJmi6Qg9yyZP85uOk4Ysoox+D5IPQZaBR+13lsvjCM6wtZ3GwM
ZCCaimUHeTH3NJWdzqiB0KzPc6AvgNFlT/jHcO0ZD2hKqp2B73nHVGk5bAccI7+V
lx2CwxYtI0FQ0rejxGK0KBspt3H9dJSbuklatPZP+VEsyiEh9XNcvohU4yiSptDP
MF8cxaWDMfuAVpBprzqrJj/rIBC9aHAHpHrB+iAl12bHNG+YTLXol+eIOBSW5bg6
c4YJsVURmlIxB8hQttMXZcyx6rFd5ckv70+T5CIm2L0ON2KDu5egzgtDn13gqtng
b7a2d2iKMxCuYkYIcEoMNgYyITgPvqbRic7hpJOGn97AHLlxLJZ0+WS/DXmt/1uS
pyHWyze00WwV6RHsw57RsGBTPa8us7E4cintpCxnDoPrPqPul/SSrttUBwFt/2XA
IkFjYKKNY24jKuoI73aSqAZ0Dkx5iFir5q9xWt97N5uFw58PoaNHzkJ32SzuLv+s
nC42cTbO9g5vo62MkQTccwFnI3QgtFKSziC4w1yvdn6iS8OmtnFQqw10BAY1U1a0
C6yhvtsosKJHkcqkjnA+ZV711xuX0P+o3929M2Nt7H2mmFArmTWWzKhJutrlVm/M
H3+59BqCgep3rb4g0cAXpcyKuG76zNdtWeGXq1srKT8=

`pragma protect end_protected
