// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kKjfT7TRH6DlAC/Fwdb6ox0jqNz0zjTEZZjew+VL0o5ROnEE59M5HGhD/GI5
h15psVJZ6m1CItzJQ9VPKontNdI1thtLetu992iF4Y8ZdPoareQZOD//ar6w
QKTjlhgWRmGk2Z+4K/St7hcioozFSYhNZ0vy/6koIUESatfxXxC3PxOEu/gZ
IJ72iNCLuXIFa/uQc/Q/QKlpInneuDNln3JqcwhMi+RHScpVP21cLVuS4fz2
bLOhaKYkQ+kv5Rh4nH1pfLrrt25SGSySjERhoUIIbk0NVe64KbQmZMfUGCho
a7UEn4RpA2Pw2oX+ctVrbs406GlK1pwZNlxUkDnDMg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EyBVx1pFsu+biDNroLE+Rl9VhiESinaEo+gwB5SkwL1Y/6qJYtWAyAUtZx8p
mZpk6gJdTJuu7jw7Z5Zf0w1qpNsXZmr2cOermL25+xmrAvCYj9CPrpwZ1rtq
5gydKX7bVcaJGUMIXAVlRQvAwd0nlcSFXnf2j3pcBnutltrqyciIKBC23gwd
dPkaRcV5qw708jV+KSXdY0T1Im+EeIb7+408yFwQG7EzGRifwzI39fCyz57T
7EIAJresYcWVghkjQM2npgwxNAl4XhMDGMIJrBgA/Ic4qcjYXXOdlnlKius4
AqJGXOulvewsBf2ZqoXe9ZYsYnd+MCxboZvIQfvKgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eCFuYQ65aA7azEQllUz6Kd0AU+VLB6e8lwWOAxfKas8dAQ4u2Y+cXDO85FZg
+08djKzhXu/yaRalz3Et4DVHCKWjTuJkMC7hNWQLVSNHkY/QpqHiB10nyyuU
bWB3aZMagrtR/4mL0Xm3u6G9t21Mv8rWX8nUhKeOHWdJWV/7MHdFvrUnbmO9
l7M2PvaZNM3WUpe0GAgYLwechj1faoOFCB3hsqhAQ5CkaMahGsy9B4CaIGYg
i63GkD5delvlNI8gllMQgQw/Cfn9K4hOn35lA3eSJkQ8MxS4i4CyzgW9SDbU
01zGTFO2fSyvQxhhLcwfQhDGMu/vn4WV/W1A6zUQ/w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Mkw1kVRTizStJGsiyPNMCuCmAxGlEIrzPTpa/dyVHYUf98c+e6ofh6DSI+My
x4cv3qjd9nEOyL9tFxmE4PP2wD3W7rI/eaUkJwSbqsq0V9oz/j5NXl3IphLf
NRzzHmfpIBl2mAVMplLH7aZJZ+1FvdeZ6gQhzD5g2x31mFUmuiU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
j8zhLzz/WKYLkO6Nav8ZGw/VnWBrbwqPanzRBpL8H47LEvpPztIUHUC2sw1L
bZ793G5A59otM3S/AB6XyrQGy0aaEUEGGLzqUx2WWT7TcIWtWyXxbaqXTjW1
K1KlzUiYmQqJ6akwFB1YGfOf4sEMbAMbOiMz22J9yTJuBFQ6LLLdAlsDQUaQ
pox72sVD4UYUH2h9/IGWkYbSy5430dPjJAZypEqYOo77NX20oxDgWB1QCoS6
sfhYTX/ohJSqqSu/imyU7sM+nt4vzbLWp72BIPS/ovoaU9jnxNqc0ZEMY2Ra
1kt/SeiLzrBPWyUS0BgtcoYRzZLtOx4Q7CaIUIo7ehVPpv5xwF56xwzP9A/Y
d3g5UEH9PjsGByglLB43ljRAYhPiGBWK0s473MyRKgIYH7PfseZLSnmCv0ja
PV/FUFuOQOki6hcfLaxfDQH5gQvK6LOFdoNLaoxnDC+7OVlC5b3FsukFjXMT
0Rbe2HpuXw/OsyHwEqALF8/ek7u/bL4U


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hIs+VtqN0MG5FLdDyT/Cl/CGBtJXJm43NdyK87lBsq2OdshSiysuJo7MhilT
qlX+zNlaKoBsej/A8f3sThzwWdovniXbMlLBC1NFmdKsGQrfBRegDpBdl7IZ
qaWjUcSgkEQ60RBle0vlNkfWy3gnEY5DpGFtcw0z3YPclvFPiwM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BVoU5dS5RefyNGQ84EhS6wCLshBUESC4JcBaaV0lKaHWT2s7ANPXTruGeNg+
SPKV4E3FzxjjRzZET+cIQ++oidzZ+Tbbb5L7/B2466yYFXlYDQdY8/DIGq44
chKtH5+KFklzXkJ12rafeyjOYgAycHkA3SingaxDdlbU91KmJ6A=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 321680)
`pragma protect data_block
HmIc+EI0VI83XycE90TdZtgyGKP6sEJcz1uQm7AB5FoZvfbJ4z0qgSIHWsYp
SVAEI8fm5HyjkHdD4rEq2EycJxYvs5LRZq0nVBXjGn7nF8JB2CykzNix68bf
HNp0e7Fg1HXvuFY+V959PIapr/nDXsZdDzbq2z8i7neKn4vHq4L9nRaC/Wq8
xjrZWQeStLdqdTXGL2GoC3RNU1Oz/kYMRZkR3oM4rQ10UKIH4MhgHFtMN7Ld
DsYGEAB0v6xd5GgKcvoG+Lt8N0XajXJDa8oC/nTxw825NrZWH4RqvRlByBhE
jaZElANS7CDzwFZoyo2EFsufl0HzeNWjBp7UhRr1OFoG2PGU/3z7KZdo4w+8
Op5egzj90w5GsN05Pl/ag5Y7n7I40h1TBe2mI3xC5IxlPCbzHPp3U9MkORVH
eVB/fa2WfJOjkxcNpPkwBe8/JW34vS+tKyVhJYKxrZMujc/uDP8e5thcCXTH
orUtFmo0ZJED21sSDxI5W2C78KAiXiOmxiotbyOMGOACQENjXDTQ/4JGWdrS
o+rtojj+8aq484BipD8Qw5fNzTtqwnhWjJQbzn8nUORArzGIvWXM1sKCMcI6
fuT40Unt95e/bg7fEqulGUVgUQGpPwTgaMCVrg7y31xS4SKLjEbyF8Qimjle
6smiAt95WskqV42lu+/kSZZnEuU86U+FJoLXSZj9JKUj/z7TsQ+58cXLFwWo
l5lHNLvg+9A+Whu3xeaOO2xyn20pwqDFT5oyhgtjLor/Es5QjU/Tmt4tB3AR
F8b2WF3l2HAdqDiVno87sXgiqmy53V4AiEglYkt5KJs8mCbuDbHF6lokCA60
F9kDFWu3H7P/90OaExyDnHt0cmbncsLPKeuvGsWaKPIEUawMy0VMCz/9SqwG
w/L9EdQUpDi+Jpy7ex62JO39W/L0TKaJUx4JPbgwS5uEp93LbgGRxJ1Yx/S6
1msCT4IiszewmjaQ6muKifeE71g3k7U3RR/32Lxv4ZZ3WvolsVBJmKw93bVQ
c8FDG5sdG+4bG0SbGfwe89fjdgod2UeltjvHPXyNffcFVLUufs4GkF6AIrqA
mSJnI7gapNFp2DVhIQaeaqycItTen6XDjGV7wOxel6dD0swNfQeVyTWuz/WE
stsoa43UILm86CwtumyAlH6/VEIzaw4I88tNE6TgAVQCiO8WVvCjDy9r34OR
/bbk8kxCrJXkzQRLxb/4cT8xWs4ab3NBPjHtkqYhrLDzCZIfrPOqku11kH06
a8+KatOtQuBwu7p7SDCzDTezeWTWqNeeGXIYRS85rAR/8yWsKGOAbrzA+cpZ
KlhnNfwDME6ftxlhJgfndk7LHIE3xDL1HhRTkNmA0eN1i7/5TtLC0VizjErl
mWNsDwd85E9TstT+7QwRRtQXC+IX1XrIsyDQAFakybSU9PZ7lAENo31Yc/1T
nzO7KkeLdrci6ppCn3v5ItzT0PK3bhl8ohK7fQQv7qvnLLW/CIaOpj0vnVYg
CgDJQZimyK3mBLvpyj1nxp9VACNVr7nD3BPwYpwHak5+fkTApehxfQ56uLtP
uQG0yjLlvBm84p2jZWczorZ0SA4pPqczPKbNn+8CZxSSDDDUebk4pobSeW2I
5Dg7WXdsvtx8dUTqHbtfl/yhhWHldaOzzmQSNoUNQTHE+JhhtQ1zRmcJEA4w
RIEE5t80/8k6ooSj4wqKu9WHO/i1OY+2yWQCamHMO8KJA0tS/dvxWZKfX/x5
GJlZsdADa0qVhaT7FNDY3xnJ+ELt1VGYiU0Rhx8G8XVLVeXomO8Tk9JCnRli
I34W7okqVHVcmG3GBX9UDZFFwRFq2VVWOX+Pmfl8VYKkkB5VMmIXfD6voQ9s
pc3I4btqrj8fINNMecfs8BO4Wh0OOvXIy1q9w76Vt/z8a81RLnjhx4uQW1JF
WEKnz8z1fimK4aE+jnILZNxG83h0YMCBZjRVMihnWnrjre0MDqOCiB1pHZXA
ZRrlwC0NZkcY586x+r3Xofo8HT55B/+nAOkAMtjhnACeqaSp1evNujIbSGyf
h/Pjf0U/iv42rW3cVE1hSNKrUCI/CxXzh6nVgkctvUgX3cDFosHs+6ofrCFY
yfJ6VBMEJ8VOkbHfph0AArKKbRedEVJfMBEQ0wLep4XjWFbw0BKgYVsduq8x
iXBNLvg39Ubfvz1LQ+thz47eDFNZ8B7VsJKkyF3wDcC676nZu6ktgJHcZ9GR
ivyv5gey0RUvhNU3o05axc7oJlaI/Hmob23gXcrBRMPOsJ47SUujkJUEn8HS
3zESurvVHqE8rXZ+aStWKfT4hs2vDeghCCIt2ecbShbgH5q/tEgRsAJm+4Lx
mUGZmMW9zAZPVtKrzF3xFqhkXXgSpVQu31BMVGbEFU2wqSRMJpqmHus6CjZm
NimPkuVnaSRWekOzoH9z34GQkCASdaBcnhA9dL4adTizDrBQHw3y/h3F+qk5
HekRDfeARVWviEsSruTbOs26b2TsmEGSxnUr7UVCuMCfjLPFlA74YyWSVh3B
NX872+IeKKEzezqyJ8EhgKiSnUxzhytAAIVl9BK+9YyDrzxkS7ZOwYD0hfP7
4PqLL9l2NgbrlWL/bcAPthLeygk27MxjABQNcbsTGsrvtYL+vg6NxyCW0eQa
zNHAHI3PWfUpRkynqDCFraL0TwuGJDVaSdfnKJUVKZxSrFEqmUTH7SsaWhOG
3z14KH15A+Fq6OG2lUOHq7h3KrIcbR3pcYIGbnBrufQCzp6DCneJXEXpg3W4
L3VR7qJ9w1Co9fIqt8KrnmCqvy/jG5ytE41EktuLQ6tDE+/fwkC+bjvR+ao3
rJKcnnjmnUmEch7GXc+UEShpcbFJVtkL1QvPF7e7f0Q/GCcS0yt9a6C+vCPq
bCOdLUOnLvpcjcHwqaJaoZU4qskp+lNc7yz1918s/TUptfEBrSBJviY2y6AP
+sfb8X8B+t8skIB3OLkkbE8jAkfnBsfWKw6snBR9G1VJUo+Wmww/h27bxOjP
HeK4J5FRqYp/c9FgSjxq5+9DDgjLUQb+aRc4NyCQvJ3PzWUtrIgl/3tqpK9n
eGvqYA3NN7kc/1IQ7i00c6hizdD/4jgYMfoJW7zSOZ2kC8se2ictxL203ClL
QOTPR5d2YmP2uUdnPUmKsEzxjF9szDgGTIuwgZaKHV9GKR0Tzd4X0Otephvn
ch2yodhoAe+0p1mlRJdr06sppDyzLXWlSMYkYQddkFUFg7gFmEPV0wg8g3eL
WTAxa2MJ9/vn+H8oEbhGBuRua4PlYDUJRpy6Wu5uEmG1gTrwMDpkoxaacRNG
E/lMOcOufJHOSlumtE7nBf1JqybMr0G4njm7jEhDWj0GWxDaf97W2KbEY6B6
uyfYA04QSmxU+tegWQcDLmbtGQDSgcX2FAkmb/wY9iiTTjWTpSg/WVI5oXMJ
ZgenZNuFptYJ9Tr0k4vAj17SHdqgxw2IHQ4izJ4dpcpKZUGEoXKTAE4G/xCQ
eR/uwR7mAbzxj1toqZ3rXNHYC9PtTBmMvHGXFQXUD/ZTSst/Kwd8bge7JJLq
deJ1HpYB4cvcYv/c5BmGzkxVlbfJtyicZ9s7ubdbeodFfmHcCyg6UqwTPzfE
zvdCHXpswDhhpFXWt3g5J5TCdjxccL2BJkRBeaJL95yBYWbF//JRGt5EGsGN
7UrNxqpJiAkFkdb6LNTC2fx01RSJ/cbQB/R1pNiAx59EeGqGx5rkG/8gTuU6
WZAA2N1sHhNeSl3q9bHAtcljZI1yUp45WkA9ybEc1rqQ7EjxooWQ++0pTsvL
D5ZgEbrs0jjdV/MjjS+ZmbYV5KIRTbAVmO0gwuCsGjGkWQ9mFRgg9tUx7LpG
gGpzm9IO1iSc9ayQColh1ok11pGmyo59gAuokWv5DKtX3/aZKSiHfnvwIL+F
9MUZUtxbFXSCLC8bysQXGAxaYFcCVD26l+ZwKD17pPenuHR6QDv2d8bHhz4+
vy+cXw/1RWZyTMEQJ+pPove4Xd7Ou3LH1yTXAx+U8jwT7Mr7O2qTp4Daxkkf
d7/l7nXOkJRsR6TnHnnwPuFRgDpI+e1ziPN9RnAaD9C1zs7Qlq/CgaIVd5N5
BqPKLYHeHzFyC8lO5yXwQNMeroucr4ybyrfXtDGpTza2btb2LeLZQ/JTZyI1
C5YL6eAY4y5T0kirC9Js8bR5AyTssEAa12aijEt1g32BekBOMdOe1PIiIRIF
bFEyl+YBzKqPkcchd8qsNABnFMLGKWeFMdt/sI2RcIwp1QaWRcscYDPitne2
iwtiF0kN2CJp5TYDbtbhl9HGt7buRAR8vltBwbL2EQd5VLkNY0sGGziJGYpc
o4fu5JtEPJ8m17/4fhfgjWzDaZLM/iduvSBQwIABhNUvdILV6OfQj/eSLW11
CgAJOEguUfcRImK/l2u2mJrjKg2Co3GeJM3Qhh2pvx1RAgKzkaSKup07Gz57
qSX6studVcYuNPUEx0D5RrGcJTvY+oEQulKE4XdoJ9gq1ptRA1iHQnD5xnEq
Ucc9gv+R00xXWKourw1wurRf2mux556YvIaqPZqElKHLcAMREbV9Hd8iAAO4
2DPcnWQeGdZMviG+wtWe1yUFzWIyt1n8PfDmIVXMnSEqbu+RvVaBHBo9+Tf3
+wyba+g+7mCYbKfChrmz8VdSxanUS44UdjIQJxsH/+EmGOA08NgAIKIS5Ky5
+nbJ4K3oGSB23fpuH/KLXO8mEUqO08ui2Dmx9gCd8VUEmAelED30fVcMZMde
V4+9APkPCPMOIpEuGVfLwlsWASuuMMX1euwEnIpNAqOUr2DtRibCDkN4+VgO
fqFpQXW6HVQNFcCGiYAgyWvVCEl/nq/1ch6e8d6LasYnwZNfHunjy65lr2nR
kmSSTFw1eeqq7kW8yM+S+41WwdxRIgqsiQbgKSfmSKqfL08srB/HeL3Rw058
4+NfNUwLwYunN+jXFAeVPNmfjeh39lHiBOd0C1J03EOGDaJ8d0OfuqLTp/PY
BJrcrYrz9mIb5icnD6QJFHFM5arNPRWnkd+K+rMuN+4mi1SBvJUTogLj3RNY
Lw4JGEeBmegZFhMhxviokBtuExi1Le29DrxxUteu7W4km2agTAMRk51A7atI
zKIa2dl39ciwraOIYDkMSLTrgqDwI+iSoD3H6f7Y7wy4udcgPF5yEjrkU04z
wSZJaclBsrpNBr3fVFCztKyUICh8Zg+x/pxtWTpWMdz2qNdBX7oPM9QcqSNY
604cjxgTqQBSopkFOvc4xCS9TaE+BlHjwGfzt1Ejs66RCRGgBBWv+cjTTDgZ
Yo1JUU2DGwSK6TVnSZyBiwiuFteczP/B3rhBn0Aj/JiNypYOfgFHuPSyphFV
KqySMMOvv2fVHot5MgQUVmTBSDHEx03YFqcIGw0P9XKtXQsmKjqbjS/kg9lm
jSbt5roR8BDRO832U7xUA91cxt7qQJ0tmnQ/z5UGohvmzBTInuGDINbkO96B
LgzsBzhwKhWM9qYEaZzs8QWvICOsZELh6UofjMuL7hfV8z3gmQgvWG4NzS9P
mYAXJy7hngYmpO88GnbVM0/oZ5loUMg1oZ2tv7vHE8rnrSSLFtWGHwZBrnR7
8eJ8YKBGPCJ/sA0k5qv2k2IKKLNOYQPTlTJ6Zhc4ZtlwQkxMW9Txbs4/++tS
Nx54os3HT+so1aUScLfoHfnSBDl4bUjhCwiigeFoNFA9nLlprS2qS/DScMn5
6mp2S6vZi8STGfca9Tbq8F+6qwMUEr51HDRH5sCeDCzD6VzU3CYAaebpDR3x
0be20DH8xBxc6TYoYmmCAyxNmMjGEnPTYNKjlkrKqUTq7wvK/XzJbwxnoqmC
QX0ueX71OZWzsEeD2WpcnplDYITk09K+wSYBOWPQ1917dmiFF+UReEjt7vBj
0YHa60LMltwtkZEgdJMym/StSO1QKFbx/zZtzT/tiqeb/f/vMmx257v4PyBY
qmcOlAsVpOMpwY85eCKDUNrSIE1W8+gWZ86r7umiRpxWCdlSoHl0u57iHSdH
15DKk+TTCmtAnTDH6JyUAWcTVSMROP6E9c6CsFX+5AA3Qq4QI2gpzYf8hkmu
IJDa1RyB4TOxk1UeEfJBhIl4+Z8EXGx7cShkqx+ULivbWdEWbT0JO6u4MeD7
IgE/4thdVhl3p5inFy535Ules92fbz6JcxYSkH3RodeBN5Rzg9uD84/EYgQE
6OcZvQT21a/bUI7KMS54lJ8ZTsEOBe/EZNv3ujtvi5D7bAZITwvaMqrpqv8y
z+kHc1wSgYvw/cAcvrWP4VNHYtddP0aOWwjoauA8G+a/Hm1OnG9JID3vAngn
HRFk894VPzU7IU90zsXXpfzRLyRMyz64zUxcUpGwMxx+6Gddu1EhzyOi8CZU
CQbLuixf2FMIPdzdHWVDKrcERN7QRIr1Vw4Z4cAOtdr9Zz+2yfBYZm1EhLFk
5/UjNBwLLmZrcv4/8pmvYdxuhsnyVYgG/oBZkAUY4Po+TqMkpJha0pCO+Qlj
JQSJQRWniEEDGkNXxqI0s8AH3kXp92FCN+NtnqSPb+HwuOrgo2YEUoMlUyAj
n6JSVJuZ4pW1ujso5s0B7ClwtLNJEvbNAQW/fwMxl0gDMUlCikI8DwulUcIP
JDiz7IrNvowcSOKS/aZ0x/t6QPmYB2+g2dq8VegQQ5j9MAa71q+5EwZeilw6
PMm/KL4CNujpl5wIv7h7fqiThsUQlk+BZd1l1Rbi5r79AyGJnL8FRjg8lXDt
9wdzyEgC+b3S+LMi+1jpMH6ymlBkLtHZK9xn/o541c8arm/WFomU84Wti+G4
5m4rYMZcIOkFDBZiDSyAaugA+r3S2tM1U/Y/uQzabkgquGczbJq33Q3mLz/q
6gcy8bK6TZy5RoRffK8rRqIpm7WLtrMbUYnkMnZRzvFwzCNCzP6kIRTHw/bQ
qHKjyLTkjXGke/wNQpxE47aK7YPdGso/sPzzCl1nslaY/hu2uoinvfZCV1wk
tlqZF7ywzgorCZQaMWSCoyuiacjw/PJzHDFeffdhZeXVDRcJNwmOnpl00ZbV
WmUQIWGNWENvhwjEbWmfeLsLeaU33oSg4DWal4UxEuBfmtNWAot5fqPprpZr
wwT/NxIIzgKSU8lPFrjm4No/eCjdCZaO+s6jK6kRjEw3YY0/YUdYP2fZIYfa
GJat/NHV5j3KXT+yMVLfbulZLaiQjgcs1r5G6Sr3QD3h/gO3ES3QxPcKstKj
Iolwt/7O/f403ELese1IEXCpKVYZkF77JFNdxH2R6t/xf5dt20O6IaKIDxHT
4s9gPegB5mFEEAHHhngkgAhkErUF/858h4t1gJcm4/9IcM8LpN+9OqBTqHFL
2U5Xi8lTs91WYE8h2TX6OT5EgQbcTtgnh1OMmRZgrUT+Qbeewy75bATRtpom
PbuPGfeJ3XgYokzvEqoSVEYsnz3cLhZmH0D19IeVzHZLUqNKJXfCPjcGBqgn
Eo3XzN3akCpD6MlpvYmnDyIiyTwLusL+mShtJdcqbGCCttaBYOAQ5Xs6kA/p
9u4VBLNhgcIzRwNoX/2YUAVL/ZvKfqcjIv23/fg6spSl+ektStRV0M7RTQ6Q
bVvZKHp87ap1nGR2/8XPbyIg90T5KZz+xf1WiLGzfSre3nLomZrrrWlbt2Zs
bwXuthXuyeE9aLigUqJiiOFUO9ruxMjGbtLC9/HGQ94fEigBo5DcnvJWUGQc
+5bhz4FragNFF9MoJ5FWGVPjfCwnSuDgZuOuOuTcp2mKbFve4tRF1oS0O74n
GjJ42eS+Ax7xD2ohPKETH8xQg+eYZUsXbEfpdM0wY1IFTaT2z089kqSzl4+e
ToNyuStyZhEcgkgEvUchjnSW+lJM6HIwIki9wPVj0zMrClUnrU5aMtH35KGA
mJ1QSTk5uQPXm5nGIyIPDJil9tEldgwR5VNzTzDYnKYT45wOjsgDXZ0U/HXP
TlfAvYiVrSY+HFdkuQGZjIei0Nnj7G8Hq8WvsFE0YrYN5XOg4zND5lqbinZj
GeBqvUyy5m2//r3ViI+ZjSBeX8Hzbl3CK+BAJwT/wio7MJ2JlmFxwnLlySjv
oeIaXCS3ThQ76FlC+RuhvKkoGzw7gvCOzL2zR11oPecEVX0ZevEJFwIAze1M
3iC1nf9mSmajcmySmxGyh3q1Jh2aY452pt4j+iVMKE4uS0TsWZA8sVtDNsNf
o4zY/nKoI69Ne/flU+71Chuvgk/zoo8xLQ7gXkxrmQMVtItVnT+rOEw+dPQN
olRzA7NcriptMH5uE/hTQeQNml6RLLz0pQnmwIdGrALDh39WsRgHmQV11BZ/
CKHm8cJE4Kl1G/V2WrxwxR8fZNGXWvMxVPTYyWM0vAiFgpQDy1KDu4iLmnYO
QFuqstPFvOAUiTmK24Gp/RraAEBy0+k9ACLal/FR2x8LlLCGQC/BMpGTTLqh
UmhbP8nancyKWbOmERCePpuabaktngI/A86RfBwju6eQunY0d17bvOqsHYk8
edsadLDhsVUZxo4snq4CT8lZd1DItY6KTAtrCXJTXq02FU7S5vy0kmRW86Q7
84NEGOXdG0QAcUrfAYeGLedc9LDYpzhD1fn/oNtoNZeZqy6PAznmPk14zyR6
bpomIkqRBdE10QalQkrrEPcZTnqkkCs6uI2Es1rTubhL73d07fH4b//U7K/1
XykP7MTOikTItFA8vnnTkFhPhrZj8wpyjyNP/sRd/TnqHQEnQziCbUvh5mrz
DFV4XjUZUurNo66bgWkwxWfXHYQVAACy+0DGgtW0o0/qBeLjn824KLES6MJ1
7Dr3hXw47FJwyGMq/HIQpPxuV600hyQLmldDg4h3fmoqDJdvSPMXGYakP/7X
BKwViMOHSgsH8JxatjiR//r/u8+h8ybsBsw1Fzo+ohdT1KcTse27H6VuZC0S
Q2raa0XZSWqxY0OL9Ni6daOnvR9u7GP5QtBVoAWRG/fyo7xmnZk7hzh47lhx
DckZ6zwfk8FKWSTz6fcmlW/pYSzQ4cCh/fLw1zFW0aFNey28MfVl2bsS30E6
Qe+twQkVvdEeBeQsdp5LlMky7pS4yTyztpRQC2BEv51g5Rrjq5PKFi45lqXU
rkGRKBIqiQf9igH+VFE49VZbm+uuVrue6a3OiNbKJAGCGbIB3StJijgoT/H/
TPghPv/UIFBtN86XzsiIFVwZfW92++BnuO1dzQlTlmHqeO0eWPu58PdPHQuF
oLepbmIcbBrF08S5RlNpTzxzSesxCcw7ucJwjsIjH+ogFA/rCVJDxcHfmNLX
mSHmkZYYg3bhe32YH4RfWQE1ziP/octVpmYkPi70O+Q7J3ee2UdFIlkerZ7o
SHK3kOCxLjHm0B6oCRrqotbc972MJby4TzoueB/hOm38/2kXqIPXIQh8QN1H
irhM6+xchfF48vuMgka+40UaHCRFm0cRglhl7U1wSU4bhxzFJG1RGLUpWx4H
uTp1nfvzOqdWZaG8Nslicw+FRDIYieY1YR1WJgYVo/V8Ngm24tDUn9Bzxbng
RLF2J7g2wqa09eRhkvZHd03erCLN5NS9pS2MDzyGbehDX9D01zngiciSCmwo
BvBjkniB50dohhyqP710QJrt9R/5iNi8Ii1dIsr3QzcZfvA6+WxJnn6xdcJK
7iJ+5kUYjrhWbdL/T5jxl2B6ewL9L/h/420f21AK4s0WxgxG00OZ7UI47UOJ
pJ6y4I4ch7621VHeKTHRNnrJ7fFr6JCTonaIG75shbP65fW9xFh3CQu5WkVX
va6kbF8heBWHmOwV3XqzSELANU6Uq+m55l45cPWin/i0n7Ol8+1+yzyGqoSG
AlS9Q6y+ZH4w64dS0/6mkNDmYdC2xRVXqfdYWcudh++bU6VqWuOA7n46sSRS
phg1mSf833ZMVuUsqyh/jmoFy+zvfFj+Oz7j1vHIFyMw0Pt3aPsyFMGcQewR
bGEdmnRr5aDOMEjG5wIl3Jz89JRX4SO/QZ7xIAMH1DhhwI8iLkTczOtJPZKF
xge8JEd/xDghysZz7QZLyjAkY+hXkTF7UOY1OQT3dFUAADx9yAMWvM5gnEf4
2D5xE5n4ERxOTg+OSbJNazdElNBLMtqvPHG20QBv7ijBjTbDaekF+V4lV6st
U+5i4zQTdkcMfmvJ9kWOZxfMPWhl/gEWH1x4Y3q3TqbsPG0JQKLF79YTBE3s
93oWQIsDcUr+nq4cxwjOSefXd9q/AEmd2NChO5rOJDfPXuPOYt9Ui4xX+cxS
vB00ZgdRSTuTMefL4KlP38lfdlCNWJB53kDAZ0ozTSysgR2Mkl7pz86Tz4XR
E+/+Rl4KWWnDQcW7NOlZ4HtXEAU8SZuSW322/YbfD9Bq5oDLNA0cYhrwqRIj
hYhcy/b/2VP8Jtmq/o9kXfOJvC4z8MkQZrsqHRNDsuIzyKrmURtvj03BcQp5
7UQbCeKzdANoxQ893BAnECVMcnCMBZ8iLko0tmXitFBT/ft9sOCU4Wyy1bBh
RP/gc9lynYGeaQK5XV6x+g1Oir1d5Bd+keTFr2a5nQRDwp1uW1uA8sNGsAYw
movueR1InTFJXSOurj/N6CjvqD9PsirHJudLWMdv0izyWI8fQb4xiSdrbq50
1vZ9UjOJQYyJ5OrheiB5Nf7LXEa8aNbX7oNA5JsWyImv6Qax7NvDmfVzuYdY
QEA1CHKurYSRGhuM5C5OeIN63i2/CzR/OOy1w+815CCZL/OzRLcnMrCVuUp7
abVXTMr35NcOd54AfRDQnlos8LnWZPI+vJrKIKIpQ9Qd9HdJIyq34f7jUgUu
dhqEBOwvpeImkWi5vNzJkJPzX9FYaFIxp8ej05W3/VD2gJqd38YVW/yzUbby
YkYOfIyzXfHUWoEBv2gOKLs/iuwol7lrg8W2aVjz522puq9MxEIYuQvmHEjp
FXJ8dKUR4dYrHL0fRzuSPbaA1BabQyihIP1SdzrdDYd6GtO0ohLzktf0h/iE
5r44aKeR8LXYOKOR7UQlxkIO63jw2IDgr/PXovQgDa+otoUDic4nJfLeV4Ck
Xg2hQPYXx/qnu8WJYL9FGBymCOJTj/vws4YXzrpsg/3/RbsiPaKB4EcjxM2R
57RCqunn0iqInXMWbMayaK7Pw44Y9cR+gXmGMvgNn1Qd401vIDb/46caBO/F
UtdpGcuj8S1auvBGwZrbHrKL0NWZw+vPE6QN7HDqf4zFk9RTqkubijyUAmSI
Mn/wMQamghaccniIdrVO6fv//aAYASmJoOuQIB78eNgMuo1VHtRrrFreu9cr
G3qTZ0yvaH4By6nzmRfMiIrTzGM7FdZWZ9hLE1TJ4pTOe1/6AyJwt9j8biBG
yXDBEP+SUjyPv1fxFWaloh7XFwOhRo8Ts+d4qBHOF/76NaXDDV+BSxncsSZx
eyZ1ObYD31FX0rkldi5YVF0v4zczBLV4o+Un1QQz4uXRpTyzngjhwbvzet8C
tHxMeds1qYr98AR3b5VUztfRJWeG/gzcRnHDTgfwbQig0k65cmPpfIc/Xxp/
jxrQv6GV1wzg5c+mMqGFC9owLtPX5stykxxUKf8frm/8w1jLz4bofdzEBE/y
MgTxFJX3PoI4oMVpfJ41W/doJMECKDl6uES+FpX0ccYap47ECi9Pyb/V8jwH
piUd9XFngE8gEz9JiT/7E7zE2Zyzzs53dZn1siDZe3KTnl7q6R4PO7MXUmwu
ORNP+xxjABNqVSGP/Gb5alZcKfxNwwzb3S6Z4NOeb1biVZW0kXlKdHXf+xA+
+O9bwiGse1VvZ+QdhICIQ9FW19F6YJgh3To4FbJnv8CtX7nSf4jDPCDx92EN
d1IMA32stmRYPBlSFRQjfZvotiqQOHp9U/anTp31I1t/fNZ6EJm1rSDU6hrT
0B22awUB5v9W6t84kxl9IL+by/An3FvH3BwGmj5pTuBqTywwaI5CtI0vo90a
DNcu14xu6zbWIRbHufYmAUeLNimyVyIZtTArU4kmDojcAef5sPY4JUZVf5Jc
sk2yQMKyX8/jdBiZTNgk78/ZB3f+zGmJ8v1iP+rGXfLyMJmZap9bqLBuVs5u
KA3Xp7M0EX+Myw7QFbLGsu0uqhKCw8h928wN5dW/sqk4OOebyIKoED/b/mE1
LZcCWLDxqjKjBusN4IVEkmPYlXx0ieyMZtHo/W7fpbzXEMDYZci2+H5WSmhY
9eRGkCfHVVOrovyrzxzwRPiHi6Lmu7ZvoFAadQTUnwOPwSrCMTrLATt+vm++
TpYK5R2S0Sn+8fuC1rHs+UIRwkho81KhEMWd1X/89S6c/2/ZtuYnH76ujE3X
VyaA/J/VMS4XC8lv4DpwPbKPs5ozc8Ft3OmZ/oEzVqcwiXS0dQ3z3hWhFMN9
6/xboUpvZIX3+47R9wzASK6a6wj07fBGTLdZtb8J5BSlYPBqgIzXr/0dlIGi
7tsl2YhO9qRUjzYTq4yEQMmYO0dYic+TC+QAdORreaLHjAQ2Z/oWHUdBfDiz
l7jdOpAHeCtuMOPF84Xm+2TJBsxcTH9NKYIxNQB4EvKivI6Y5n1NtY0o2IYA
TpQQZa/FOuRyxK2c0VR6OdIU87diFGsjTxR1VbODuiee9s7cwry2b/EZJLHn
EuAdn7GJ8k92zhLF2sgIELtT8UV6pRVkfDiNMMCO/woqrifG4gi5HmuQOgdj
uda8jWYZsdSep2+xUIMd+1tCWFlMeHAh3rTTIEhkL/7q8Q96lyWVjfQBb1NM
QZyl8YW1mSvbfepyJd2pOUeHqM0cUH2IED5GaDgLvsQtBMQsjNM+cbTmOnLx
gUhQw84d4DZXohrAUWIVf7MiSWhXFPsuEkJSUcZPcpSqoEX55hu8CkRGjyoo
FUm9jTw5sbobbQcfdCVYg4MICI4tS4KWAQKlMdGEgg8loDMzIf9OusCdgUxQ
FKvTS9gJEio28GnavCk6w7tRQc9iDq0C5OKircevfWEpjweukFUCLJc8q+W8
gFNia83KGoBWclDCGTuyDgC7cmZwHhfIGqnP9lnAR2S5k1//6makyE0aUTjz
RkNpjdbAJ8HWKEHWgFkB9D8igFUB0Q0Mf1og1lS3CZNouUvntxYp8xbLetHO
jxkFlkCkf2UzBnO0QX0vcjPCgKy1uRyMVLRyqzr5KqvgL6wogcDRsjUTy/8e
PAZgBR1V12Qwa1UUPKb4hObVzPuyzZhPIlsBFhrHuG/rn3J7B0z3IUwWMuIO
cRcwJ7DiV72MwVaGIDVaFVxjANpZrZs2KlaeigKhYrpUrfYkygy7ti2gRxbV
KfZ8Xt7M8OT4kVWZonhTg7ktEcMtCUbtFg8OuE/VWN0kPYejnwp8gpofWVSj
GiYp85emaVFnTmeG+g8sLshoHFP/jx/BVnX0g/e+bQcWJwNTl2SuwBNVZI5b
VAVxuwx+0xzMQPq0IUjHwFc/4GjwDMfAHA2YVGN5Zk6D8xetpT2VSkPEblPT
1EEjndGJfpPiWCcDANybZF2bQqly34pJYeop94QhIwjv7uHlW0j5xgw+q3wL
pCxMAxkLpm0gAb2ifQ7S8xVgUTFzJHyR9Gfx2bgF4dQb+zqdl+pYGIc+rV4W
Iis0NPSUPlB7VpBKwWKqbRv7EYRf6FtG29PeBhPQbeswr4KrqmT6etwXDUGo
Qyp0eA0e8Xvy+FT3Zt3hxVN9Ed0m7QGLEBSCT+AhW9hol2vfe9kITMAe+T9j
eTNeeD7B7jS8lHCQreWsQH+zRdcu3NGb8sSVkj9AYt+meTZhOq6q0xN1WVUG
2gW5QHAZW40UyonAHAtz5RJfTQWufDLeV9RHG1rTZnAy5zyAL41OlpgFDcU1
tjP+9Jr3oFrghADw1QYCe5MeY8vLZVbP7b+pzN8kF1VpjjCvLP4BBj3rA2uB
tij6P9yVkTgYNuj9MR75cIRna38FwOcZCjAftXVqekHFh0GiDjX5JvrOT8U6
3wcaBfUtFSUfDflj17hl0Ujxpvo0iXiXfpUZS0kGWa/b6Af530vUnsDil91h
FjM1GXiwB52Gf+gEbHVGx/3JMhpDXFOtz6WRr7cy0/cBotIVImRfkFPEPd2d
4G66cLsz/OrArHtgpVJFy1X4e87sTaypCMrMDiTPZWiDe4xwKKRbCddMhpQe
T3mKAk7VmG4asa3/SPwLzlhh9jD0gy9PFgr5UjUWQzbE0QkCFI/vvg5joyxL
qe1YaBvwM7D3VWE/A+7S0K5WmGMQl0tRn9EmO5TOgDQB8hksLfvMnWs7Uvzd
y/1LLeXA0wIJ62ilBYq6DYVsj8SwnSMKoVxTEQpCzhneFWWhrZ3Kz6dKWQtb
DaCps7rqhEhM1TVFHsTXTv3X9Lx7vM16thdNd8h5WNHsXlkrmO3sAYN5+ISA
0OozD9mi2XLTpQ6qV1xJJ/apBzIjja6CyQU1SYxznk0XlIO4M/+dhv5/sodm
/dIUQdz1rkNZ0t0GxxcK+y51fI9mfh2CsNdR2CKn95Dw2mwvh7dSs8LTRJAC
abaMzAsMZXSoqIF33ugHyxPkDaYWrXzoFkq41I14nMhZhqHMUe8sF3VKAK0J
fE0g2pY7GKr3ols1SS0EDpkTSidglFMMWV3zHLQypf99dHceHrPnNGCGQidv
vwZEbUfxTbAJtB7D2lnCv7yU0qdhyozPI6OI7c0mZ46S8Cfqcp6SjPWnEdgC
iWSDTi5kuSg0JW6M2+fFrgAH+DxzPQ3BglEtpTdBz1jnDq2yQB7NXDWNJbL7
2SPnOgfn47erhvXkUJxh79o6IqBtqClXTmNkpi4T+z8MSW1pWQvge1RFeI2C
vDHHjds9Mhbz3+Cd+1e8VN1owxArxvGF5c2eYxbwOAFqCuU01XacPVGX8YYH
C/kcpZvZY8F9L/Bh6f7j2vGemZp/CNZfOYxttL/qFyFq5dgulzbDkDYxflbr
l1E94SWop6wEcgfGDUqz6WeV5nf5CzIKKbmckJG1Y+EH8MeCI8itLsWed6ZW
LMOt5iIe4wU5nmkBJWPj84UnDI8oE/lM/xaNwYJ6EyMq8wdKoDWwlfjgMqdJ
UJhjY0H/hFYnLm4e6QK1TXbm70HgpFeYVje7i9B+C/xKmLvIQo9QBxIRbN3I
A6V/WEAh1qwTbYczoD/LLvhMMxtc6DdwbhOQlENGtft4UxJeTXarAaIMJ3yt
uXgX1FdbyqKdf9XcyRgOLtb/LOYrI3sG9fZzv5f5NuOcAbTvAkz4wIaZQvKb
xSQk7hQmcnO71wnJjexdXMcDVU1jxlgCh7pnW+axDRiHYE2+NmstA1EOJtPT
M1uDUOfCFi10DHRD6YnoYgUIbQMcyN0IfIqAbSP4U6MNivsjUJCapFJStkkW
nS/g44MtJ+EOf2BlpGDOdSCjI2mWOr2Gy1FUI01q7OzOEx1w7/OD/2C4Mnuh
fUYSP9d8di/nJK9VKfGz6F8QtD3DYGeXzXSJEsbxl7mPO5hrVOZzbn/KNMyH
+sBjg5tBr4s8NcBB53wmlZuO2CKl8tW29Vi/yWzhD3jlk1mtmuAHGwSSkwoP
IYnKYEFF8lRCMPQ8Bmcki2NdiQ9r5zYD9kR2PreT3G8IrFMEzyu3WuUrtXo3
LD2+w6LnqA1JHxRa3N/cs3W3p76vek2LL4aVyK/gCn+tYlWsOYgPvm7S9tCR
4B264a9Ptm3oU+3BuNanuhQ7tTKAWbVABe3os8wzlJoSEDjv49t/yJb4r/Sa
pyRZ87vQtTKLjV+BC6LhdGXrXSEzkXmhUvw376gep0zQUzsf8zZdKE3f4Fbk
9sDqcYsjhtpeYcsKIjcjImmO1ISnI/sEIrhPYhd0ZzmP06mz3CnuzBR+MTru
4OvMoPpBG9hwqObZEVm/i1MST5tle6TQvS3N8Gb2cqXLduPsjjj3xSz247lo
x9xnWvTGWnktMf9H84sCuRLoyIQBTnp7rs9KTpCCGTdkg+4WKpT1bXoPglEt
vzkvPsBgMq9JQRrKpumIsRWxCKP6vrj5v74p81mOjAeh7cUdV7KInsVgG2CW
EPxiunXoKUTtOR1JOVVp3FvIQ9XVcRvOJZ7I4UrPRlgQBaG6Jvm6b08nd0A2
p0+XSLip53IxGozefEduUlmtCAwrkkV1ZopoTArwMuSsvsVxH4BwjzEtA47o
UftANcyMn+XyeA0WUIes3k29uj9luSrX8ZZVB8Qz2xC2yL9EbGusG+5dXxQd
aHKy1Rpkh/UqSHPeHyaMd3uixqmnmtg667nt/FxNwnrwOPFNScq4vQvwP/Ig
lGzKw064VpkoMAXuOUUDBaRABxz5+SSpKF2eRec5q46bedvAYeZ0/v1McysP
2uoFmlzHjdRONvSBUVKFc0Zyf8Kq/pN/0SUrFJAbiWD/vqzdfWCt+oZ3Fh+O
BJSAQXrlotqwExAooTwpVwLLxBPgVruRpiZkNDHemmrcEpTgBh/cP4Tp6X+Y
hzoGtYGRnnloIpQYJCPt+MfBVcbB7se2PJJSYpZHGUjhr6Hfnjvq7DqhM/jw
JWMfzC0uhpeQI+ZwV0k+e61fEQBsRxQz42btDO83G6OY28ujgZurR98PuQLf
0hqY9sFeId+qz2DDm3q0ONAefEEUJ0Uum92g2UFgT76ONrNStbUB/uSnth9z
g5kK5x9gy74FVzeLDtXwmtYStOurbZwWCb7RBQOAu7+JXnZ4Qc73JwnPi44/
owWt4kjK6OYHYwaCvKWEiHftgGmLR2Diph1JeA+xxZhW0+U58JBA9pX8dB8f
p3+rLe5Z5G3ksgl2SUhCLfNTpKXN9NlaXrq7cSr4jaZPanVUwTGj1bDIFA5s
rl7aD5ilazu8gJ8+ZYAV1HwZMRFtq027yoWgpKLjoBz0DBSOe1yDX0uhCxML
dBcaiHXLr1/TE4pDrAnGYMQMwctdCF77m3uiVf/0UJZHzlgIoEN8MqGTsEnU
UYexUkv2qWW0zBJB04+iPFf0z+kNPAOqx9XAmWv/TItwndgjN0T4dILH6rgZ
rRJKtohTptpIAzma6wcYmZ+Bca7utRg1AiMOBsDEQckc4yjMm1BzSVR0wsCL
9gcmXcsYDM04Budy3obfIsynEQa3MQ3K48pOvAcO9NIdc5Y+aKpRnhN/ACbO
L7DDZxkF1k2TtxDKExt43GqhhQmAOl7X0lKPnAfGcGf1y1wTnTZn7Erxlgmg
TAVHMpU3BmGZzFFajuxPytlUHi1mOglo/FV5kbbfQhzoHbZGbI8m1EXxgtTv
vCuXy8wyGFq7UvZ444ZAMaD743XV8WzFgWdGTywyS2JKtXLZaEgLTIPHdb77
H6ADH0btL0VovuxkMmETArJIoChWZWt135PV5E6/rI1xbJrUZe75F1LFNpwO
5TYFc/AxQbOr/OGWTDjU7jMsVNLYWgP111ZeyVlFC9OABSThc6ofc1zD1Vgs
/7Lh0/K3dwPnQIQt3UATxvr24F+5OZnmY179jtaCizhXgIAh2l7X8AUN473u
xIAPB2r2zeWZCqgbQDJWrpye+97srWtZyryTv7y8DcAfr6PDK4yk7Otnn2u9
Dc10iVLMQFdqVERQVDvbq+HTu0hv0nsa0JtbUB3wWaIAm0yFlWN2/ZgiJwbj
u037rPrLiaEwNQgrSj48pqYv7IGzv6XEq5L2mZ6kl1BBCYsrAymg0X2nVK0S
nPIqLUl6x6t05nNosvig5IJOIYstXNzmUly2oJKiuwgcKFB7QaGCpVTdMcOV
aKfPIqTfZT3wF2UG2U10slcQXf6+njWHhwXmaXCKWoaoyM3iubPBXMcLWiAC
3jri9kJTRUp8w8XQ10AL7E7eLjjC690PqVCSxDSUasVeDTaRTmIQc3rD1w3J
YUWy1aZ3M3XCz6co6HdaaocG11U29Xhhp63tNTQz19AL1qkWUdAnOzM9QVbu
sgP6/BuoBJGxDjmfiUvTYDOVP/aK/6B/blVy0yXGetUXZQDtso8EP0CMaHdp
cJG0OwUP7Hb3c1vGID+YrhWbWH0F6GcTfrYcxvD4s6iw56CuiExd8LQeKkGO
IPGhuwaZOhfwhQ4JXYiO6zIKqGLuJ62sz6pzUzdd0my9gHzFfoPDUwzrwZ66
1SDyDIJBY21vFyKpqdjtj/UFAafh4TdPABt9ZC5XgdeXior9axeN0FabIMPq
LaMsQaW7RDuTKyu/QAZAyJg3/7ovu6lOmqJAyCquRJNvHRRTt1F57cIGjEWO
2DIAsxA4j7mlPYptfKnzVArB3tfXdnKWqrhdSG3U1CJccUvBvTmMj/mxw76x
dNHxf71k6WSoJ08E8xEDmZuPYcaZdBvm4jDZCe+jAhZIGcBH8DFOAgn+ruF/
8KuG6Qt0mzGlPzLDLhPPtXDLY1bDRRxyBgQkI6sdeMcFETXqeAJvwrRLHVJ7
CC8IK3aiZ/TUKHjDF+mhzQkJLq728sERSESjf1tSEjy+y2l9loHreiRIjQeF
XYkc+e1zTV9sqZjgrwMVD+dYH5NTpRqGwL4cPxfjsTwkVTkHaEYlHqOl75lk
awTIDp4oHaXwMwpf427JepegjLE2gH16b4q2ed+mpIcfm3yMQJ1wqFmbGGUS
SIfP8N1Mlwe97jLJKv/qi/+7qCVL2tTNLa215zBdV3VtKYL1gWA4gAWUgAct
kypN/D0MXE2p9Wdi9ZMPB3xELGm6qlsZhLKjK3dhM2rB9yTfZNdjvg8aZ9UT
ezH6Ract0YlcYx/vw0xNLCm7FWFu2wNaHuYYsIcVqJmvNEvkt5O1+EvGtKj1
dDdDEI1/TAr5OI9a9bjx6PWosGXQ9qhnRHYhXQBPEk2XvyJM/dNP8hQlWuNT
3tyPPayb9cwK1ZQQfMK7bNuvCJckbREW3auCv7DQiNBM8MWUalpgMw2twBFB
qP/kbR/oivqBR11AXujpVKNJtmrDjijIjyzKn9hdwqzEGH1lLiaj1ReimDQ0
Vw4VLnKp1UH+nwwPFGESRumwV13mX+nvR+tCfXkGqk4O4jmyC6d2FcyKzorg
qeaAy3QN8lUAnru515tVpY/Efc6CDIYmtWol6uVO904kjX19nuQq/NGZOGzM
JbAxp8brLBBNESxteIeOLaXPCi1C+/zycaGbxgOtfThWzsKCyuD0LqOhV6u9
ujyhijjPfbXMU1WGIGDaXAapeLVcH1iiXv2XT2CJ+8inQzf2M/ZMQRHjCUac
eaWRbKfcDZyTLciEfzKpSe8bmdxVyi5zcDj8szrFaaVm1q9G6VZ+E2+079qA
L3R5ZRxjjy1X/3U3WEypcUl+H7nluFFbDDbqT9VxgkyZDbMZxsCVAWdT2OaO
7U15jTjdIeysX089JzPqSCFofZP+rd2EVVH5MWBfrA4/IZI5dIHRPAcRA8zw
cVCZQ7tCzo9qHU4slX2sK2zvV4sf4aZFoH1iOEebDRqBLngWyXbOYOeu4Iew
A8jwZ2ypwD96t4bhQdWxrfMHP5xLxPpX6n1o5Ht6Ws03FRuzRp7VaYkvZDmX
kennDhAF+XTBaO4zO532p2Ec+Ofu2IuWxge4wokLMVRA+04r2G/NZD1jkf7D
k2p3kNOGfgxWE7gsBjtYFdm+IPsMZbpE3ntpi2PDWD+xhJLAm2o644gls4Gs
y7HIlyfUcSSusUPa3fhOQ4cY7VuOZzFxmP12n5kR9YzBFDPCZ4TF94igtGGZ
mHhAxlO3ceH/Z2LRo2Ls0W6hd7OVezb+atAORF4K2s2rpgrLRrfbgs5oMRgw
X9SH0YzqTBBOAoyiif6QeEKzl+WoqSg55WlitewVCh+X7cD/Hb0xAr3g9Y1A
0ciZMMnBhbf4OW/sNBruDFzzRjyAuXfX1tG6Y9pESJzk18bsaRj/YmoaPnj5
sWwHz4+Mthu5BJxYpc5ihCN72nnoZmuIvmgS2rwncz6o9DWHy+2BpoabP7EK
FG8fH/asMBmNlHF/Jx6SknT8+I89pu1TVGw7BPHerB6vNCU4RqUVj+TSQ74J
mHt5/yaU/LUq9lgTWg0/bTm84Qke9zl+otK7KWhDbcn8YYyib3RFYSuonfbB
Y/Dd5kIva1qKKb2VdZ4N1HPS60q5xBAoHdtnW6sVZdhBjrFmAKivIO4/zfDZ
NoWo+Je57liHIHA68I3M5LoiSPESK2qsXzvb7JhyygDHnpZJKI0xIDYUVH2d
L8G/0A5iYLwGIi2TGrg6zMxX3YRK47sGAm5XK7n/DUp3YmJ4LsbASe9NsX91
ya9SH0WbFgDngg8HRg8DFZdhC/y2aeschXRF4EZJT0Dx0NAilCotqJYE6yVW
jZPnf2QzzI3G3aTkYihj+W/HKGeB8vw3nzmmEzTlkphG/KdEeHqy9jbNDAJT
Vb/6/Wo3fUBRgZSeNZK9fAlJ4EQe47mnvsyUY/m1KhFICqXstZSjcD93uP75
4PJhBBzlReB10X8gfRii9kml1FUamBzFIt+01YJ/eFtZVZ7bD0++Fbj0Ps0T
aQThtQPGruddEOwSmkcz2cBOKVkN+grBwY38uH+33yXVCPtb0aV/cU0u0apv
3TrHRhEp8PsQucvLpfuGM6Fj86TT00hR/I6nu4fnLNT8F9Tj9QKsOb03sLtD
ITWqnYmvi8TcJlz3yciQBWfxF9wO+XBj3wv06vb+baU87R8tI7HipQp20xfH
R3xnTgUCe58kIxXRRWA2r53yIXCL+eOim+7p4xIg4biPX/kVZvM+K1zrI9ys
7cAI6Ww3gKuXUc8SWe5PQnsih402Wtyp3k227Oxi3szbOfz6RXZIJnNMl7b6
JYlDDqueHL55naHGh/+hhn6sv5N35/YX55RJef1nN6Jy9amU8vD4WWxUQefF
Fgmq1q9jbGiHJkJeA7t4BYiB3rKfk4PuvKJXIVL17bxXm2OY9ZWXiqRL1ipl
TbsmIKUc7O4HVYVXmIarBYDOYd02HHKGKCOHMEMJc/99oKkktSi1GSock/W4
xmRHyBpcdPz5olYF1CsWmexlK0c3bul3MdgPauq8RJbZI6ArcZuGaFthh5PG
bZHWXSZ0tdr4Jpt1qlrdh8aPE52t3G2MDIcsVOmj1R8UwKqp+DyTPxn3m8yB
1WxVKc6czbKysowxsQPatoW6mupTgmqjgCFZSg6Vq8m8RJG/Sc+rSja9xE8Y
r/atwwshDonpLMW9nviT8iqIVPwHWwpReyPrUr8k3qttnXXNDK3JIrMb3rvK
u6dI1XobCLUma2GUCmo7o/0kTF6AsYeclx8hVlCUF4KLLPEfSikBET/TPT3R
Tyj9V2Ht2OBebedOet3rFgp+eKijsLwilkY2NnDZzBe8Q0qE7VXxMg30JIED
sqoa0kHM6rwmTxEq8ucUJOHRJJmRBF+tZrLBsMfEfrTxTaRZArhQmhB2C4L5
PrHhSAgxemgowvxSaJ1T4aDdAI2t/kDoKNjTTjmps8WqdUAEG/ZWwmHsz1fp
kG4DyqQIRLhhOcQndqzQwRHKxZbcSqSCGRi2CL/RKd6cBcbpuQnwcCAmZ/N9
ScVxO3jHGwbpN+EGaGkwMc3mVXvVbbz+y2hpvFRduMzu0DU9U1yCmJlofEHr
vxr/nw9ZvnF6q9cAXG7AKRPsB5T9w3d9pF3saz4nwCjJR3ogvatBot1MXvDn
0fH6uvb+sSK9oxfK4udInR5RZ81ZPirKGv854y5uAEaVRbyLw4uq5KZim5WH
PIRovT6GCtPWPB+s7hycJ7C4Qnm2cUhYQRcHpAcHTkt9eQ/xRWOFSgUCA15D
75HdYSL02rAOAmer5wn+fr0xoP0ndeiiF/IXI+FBw9nfp33kRHkxMKZtHlFa
k/ZhmiKZGi6PqRbTrHrRwX1GmEqronFfRZGf+4ZUtzy2Y4hU7ZSWyEftinCT
zIeuh21NLZlmrCq581hPt5bv5FU5e1EFd0sNtpZKUZYdmog96cwOCgAy7ufA
O/S4+aKbE5dhC1+3BC+DR8xKmR5BOPirrRz5YvLWadgiGj52wOD0LOjnVE95
+ktPg2tpteevGIP7x/quSkQd5XHR8fi47HcigggQPKjgBxnv5yJ3xUSSjLfd
qpm8MmlXeGnLXogeLrLKb3GyC1L5Ri1aFVSC6ZJfekfD0IaO5f4zpL5lA+CP
kcTbsKEpdjqikGB/nntx1lRLzWbyHdt3zUZjIJFE2q/I2EhGvf2MIvL8a3RV
Bpp4Y4TXN7LNxKhvrseMvlB1MqtW96QXzrxSBqB2a7cLkEx9a9l0oyY9lw+B
KHolg1X3OfpaFj5y0jDue4kVTC58j30/JdvISIjaps1jpRvrMuNhBGSkzrpm
S0G+sZaoDPzxsIrNr9Gq4WnWMoOdJX6BpAXONHuZ+v8hvI4Ke53y7jkKmstq
bHpV7FdabsOEdFjQsw5bJJAvKg9sFg2ri14ypYbKyD8zEavKOgg0tl23E+9p
K1t6E+uU2AUkKLvsTcwYrFITGmYIuJKviJqu3ARmHCj7DyssD7eF7ZVeEcQ0
MnDAwQHGJAZGibQIH6XhFICBhe3cEjfzYRslEXuElGQaTQkHUnV0+y4tymNs
t6YfqDZgWstiOTa+LCdAHXTi1OhUn8XdA+oMg23PSU+TToAWUM7dl+CHGS1/
iC/9VYnpYckqLYaGYHNd9FN6lZi7LHfesBhCJ/fchss5/7Vrja16648F5BQH
d58DZ3Xn75RuI1DgebuD0A72uroJe1x6zYTUCrjzPcfDKxVXKNJqc/CE6jpn
B9aUrOJBoT9ZOSuVmYIX2KqaLG6dqFW8SXmzVNDec5YoRfWvtUyIpiGAThmL
zThbJLw1NQr7hEKFlDCdVzbhJ/JJkydRqR3OyTgAX8uN9HUscP3xJM2sE/SF
1XjcMhjnllTzKJAOE/PIgUuU297tbQ+Q0bB4pVcrrHNEMYK76KZf+R2LP/XY
FGELyYb2vfMR2I7YCEhbGEaZZe6LS33MoAZT0jlE/42/n1NrXFo5FXwE8Vyc
py7LJUcS9umN4fuuyXcrUlH1n3CztgFGN4p1OsjdTMgHn6o++5w1OmIOqmQZ
Fs+OlGZzTCj/1sMrxyRgl8beeevBvPWkyVCryKSHJsW0kh2D2Zhz4CLsAnmS
dpapdn1to85NQ6rotJkMdaYSPQcnfgq9ZrVcqeBiuJYBxaxztCBSAJIZmJh2
P1cCcau9vZSMeqgLzk8fe6hZMTwiamjqyuYSJZAsPVL99ICztIULztuwgCNd
wCwUN/9UD3o3Al5UZuFVd+Bcr9bOaIn7WOPpWh81+6u9k8n9AKd/+PNQ+eM4
YzKWKbSGD0UAv/h87qQCNPqRq1GBj7ODAjBl9EjoDviBgFTlhu1n4/Zf5UpN
0QWahYwx2bf5FIqHDmL/KL2MjzBxtTyq8sYPH5+n/Rksl1ZgpyDmrkmP8DXS
LmMqwUlSnOFelnkpsEqeWKthn/wbm3y2mQ9WMBq6T1RW4c855chubCTpYF5W
mOEztSyPBGSP5yo7GBRl5ASqif9thNh++qi6kh7YmxwBsBghyXqb4efg/r35
fkACVv3x19xXAbM/m/QIUk3f+yA46TP9MHe5zs6hjNqeKO6P0FwDUysVHbiv
/yQeJzEIn/orzQpqXGp4u7aGfEdRDr0lPpvNfsz6AY/5/H+HaCb17Z7gYLyn
Mnp4F5vj5oAt5LonKKwqmLNJ62AQB4LtIbOpZi1A7MmTa4pGYlF9z4nbva1L
lkVpWqxN0Sx7apHHrAEIc2DwxUnsvBmzPg/xX76eCYgUZJH4y7rsZGKPNZB8
jCagSrzYgzlIQBVj9lyGZPv3THdy5AoW2PAGNFSRovdwCqSb69CvSSRLPFIA
JRQ05fpvsFEzdEobXZRCXHsTcJsAIpT1IZndCF737iUob1X0tv1c2ZTlwfXA
ORZLaXy5XUUZM49v+jDII18aBpwB9+nXa9LmfkGrKWbsgujm6/UEvM7fP3td
Xi3LwFQREzYPux0J3ILFfiNvhoYeLX3VFDuhb5sp+ebr+XyO7oaQ/6zMQGqx
/jv4Z83H+XvhKzhMWlcrZDqcr+Dn9/5FXcbi/tCq79dj5aL2Q9Nom98eJjdz
Y6VH8A0oL5o/pVl6Eb7cM1yhZV+0rnjo6JhgJZ/2Xnw+OG8lZjF7KLK8v4+y
yXewFnXJPIcVE5EV8C7/NwMMblWnlGZw5DXVmhqAXY95RxTxLChldTKUxeTE
u8BWkmXd91l03SWOrRvF3iojVghhbB19jQGz3TklZ3p1/ffqonxx7+dKvhpH
tKnhB1v90l+4xw5tb87NAD/oyLxJp5oA6mHrlsWO5EIvdcDk+t4jcddjLflK
BJTu1jss5V2mvRik8BWoJZnxiIEPuvLLb2x0tz80if7swHtk2x464SE7G2XI
xJMIfciiutv41NuNwGy0s48evTaivzDdP46GqA8KbkoHcrG46YSMvCIyYbjI
tGE7oHd32rDDv0edOpvFhXUlq2EhDHCubRriAgXisAVs8Og1054uKOPUrLeT
dFttqx6HayWkJ/doBM2kuUllh5CpjfH8O3ConvgxnkrTpsLUoBmqYrPxjHbp
ILe5dflw26e8NX7l276TTTL4I+YK8gP/kNrjMqJVggB7xUyJW66G8RhsRNvx
Xo2Lecy4KplyRLdlzBArtWc6XRTW1F8eibjditPyMeYy6F3V6iLRGjIaswPi
ndhUlCcIlWCTQVK9al2Yuqu7wzCKMUeu+nZDzOJxOxF02s6tZMerwYpIxy6k
r1FlsBMe8r6AffsQw2J0iHCGwkJ7dquFvwVgo5ZrWaMxw9nPiGDTzcWZIDo9
d7RHobH5WvdCqDZV+KnJHDOpuKVjXImXgCwSjDCqfEMjZsX8MQErxbigPer0
+LDhBg6D1vJpKCxh0/zrwT27IStyhDVL3WFPk4xN4jNNF1DH/cSbPE5fwkx8
vsoCDu2tsGLPsVKlnJ5zsRnG8flA3U5eYCuZFufsnQFu6krHxxAId3v1oFWh
aDipfii5GORQIOLRvNC2k+1amrjgtK8w3n1o3/onbXcj9qMYxbCI//piBgrW
ccxo4+eL67vLor3krDcWJsWIVA3sQs9XYcN+Pj22hb5XFdoyc9W06lRtJ8Ng
93bnOAeLnXCq5DTHHfvcpOiHNxkaCNXDm9k0pehXVtHyVKfQX0CgoOkR05/Y
u7060kq0VQyPT3wnKoyto9Y1f2WIWIjexcT3w+XY5n68M1bbvVlxtiCrCdjR
TtDM1lLhpFCoLvp3Z9Ixgn6vln1hTHRBUMV1QRx3G7dTirBxAPCc674/1Ge6
wSj+mzQ5zyZD1WtqDJIuc06KQqfC2P6xi37YlHzRH8KYj2hdOz0kx4GjEuxR
JffKdCft/FdI+SJjFCxsBfE9YbYRLq2T7bC9SUoPeCyTTPOefuayliInGcrY
0ZL9cf3RHZnqQK1wQb5JJiVgDig/wP+CJ9Pzz8VvXniLsA/jT+nj/wADaCLK
OSTFDdBlzG9KlzzYsxM9rJ4b0oUVPCCMORras1vOmoxGnzffxOHm5+qO9o/m
cHWB7YI9/fLkHR2qcgau6fm4A3aJAhalbBdgKbuchYVnSUjSLeTNrFMQXNVx
WbSfEuzNTsO05mgYAtLdQPXg280PhM1eTnxhCbUydedryhECIu+vE6fdw4h5
MTjrYZIfVyveORjnmS+iVgZmGVQCTncYrO3ExOFSlESWF7DnGGTzcRPLS6qM
w0b+ijwbobff8YsYpKtnTFJGYbpWNqeXYgTOhEYwe3gGY1k2vSvLnz2t5pYy
IlTybaARoIiBLnYwxt5gE3adbK5txJvVaPOdEHTgL1le8w9xzvQlmLIGupGK
e5pqbVekNtdEii8cILajex83jBTu75nGjjZ62JPfrQzq9CqsqQwgQUBDygVK
Dkz6kNNnJ5y/EN6D6JY+mUAAz6hMLMGmUzXmwuSeKV7uanqEkDvVO3wRt6cN
5crN32llO0EcjXlMndpwzN6Xhz7iHVZ0Y41QFpNsx/MwdbFcBNgYCc+WkNkJ
G9Pbi6uNvADgt97b1H4jX8OcbbaoSrkNpU2aoQkYqlicPxRsllnP5W88sFYI
IE4vkjVMVh/zAy1b1/5zFPeyQtriE/uJSVhYUQ8RGgog1dOQ9MNt2iHBHV95
WNPh5c76l+a9asQAZfmicMREYnqufU4cutY0DNu+hjvLeOG2SdidNX9CNCjd
oTiP5IIOicaJMCoUWzaA/4WL+/TO2vhKkk9pNOM5JGSXfh0STO4TRXQS1r4I
YopIpdbWK/y7X+I4LC1XB2HXRoaS1Vu6RVnuSyD97kqsk/EIAwNgy6gidB8k
l3iUphh7O/QeKGYDfQCaSBagzI6sLLb15TOOn3W+9T2TX6xtz+Ay8f2yo5r1
z+zBm+eyhqoLbUEd6RCS2kHqs8hFDBAal3eIUYhvO4PkVIEJeuUAcnEFu3P/
trgI3br/HUxlOtnJ4vY7pWux5B4YlILcnzWMdqeXzaOU2hcYVHH0Uw891Pwc
HKr0CYzwwP/NMkMN//b8u549jHTkgrWPxWS0j9euxjdx5DOnaNeebBbLU9mu
1rP7RLFO+gb1SPANXnoss9HXVNZoFPjc7dDnaKoquN0kCzzKlkb5c97znHoW
tZhSW8Dj0nhfANiPfr26zXpyK8VLJpMOzr2venpX+PG3sJ3/07ObLrP02fdi
1qkA57t2F2vqr7NBGsG1mkYXrzTy8t65ITB6zCj5dESXmoPlgqQFkk4Rjdil
/n4yOlU/BNDEN50VP88gJpzLRGqX5aQgbFKJDvd4DxwyegXV1EOCWgOZXzAD
Sxo7YUXMbGev1nnUPeCT5zDBgDGc+kazIk5IFVIzdaS+td73e2jt0DnXscXt
K1CldJQFSIvrgPsCcSvRzw/kF12UPK5htHNSkZhQg86+qiz95ysc3zWqJPTt
/JpvO1fkUP/Owy9aOOM9Cp+EvttUinhceiYnjbf+Jc9LcIkeU2wV9B3ZJskX
A8JHEHW1ufYMQt7C8N5X//P+zesP0b2Vc9K1uBU6p8N2S4OxHYf4uXMCG+Ac
Ex8eAjBJYsBrty1y86u1b0AHJaCwxkJcYzezOwIXw8neG97ydN76Ey9ddRjA
3QZ2Aq3i7ka15Vi1d4fEfTFFVYvmns4rDH2yj2kSOeZkavzMK+s4lMpA0nop
JEH5Q/QGCih1CWbo4zp6AD8GresrDn5Jp4CZxP1ZsfbQSGYR4hQeUUtept3q
jbChJ6HfNG61h7rC/p/36AaOGMVAKNXAGxapo3dfpmbgF9xqyY36o+dOomDV
YWtevmzQX61slVRFIxMKdWBUPbHNSkpdLbAQEyeEisH5yx9s8xxF0uLu0hRF
dBXsImf3pAc+nDqKQ4ZbMDKnZsByKYoT4PNCcP9llGYsQiU80VPHmfkmIEEI
Zbm2AszPNcrMwK2LbayttugE9pj9PooMXAJVOwmz7ay+nwg2fr7I3JskUFZy
rqxkK+bt1fTTnmWbT3ljCKCT42YbkCHDCdZNUH/HlZxWgdqHNyLAac9rajgm
Rzx/MRHTLKzPZB98LdcrsLF42PAEMwt8OcPZKNHtS4gpNHO9YvpSonUT/LiV
m8uieBJTdfomLxcHIVJrD7rLBwNXhX4UjLa4+dDsSyJEKlFewV0MlHNw47oR
K2YzZG5yJbK+M6qomp23FhZKll/+gDfeReTRuKAiPme0eox5uP+BY5ypSMdg
TsWszawQNg9Vpck5Ex0e1Gd8F7YaOxqRWyZPvcoix+dklx3D1ZdQ5QuDk8YZ
5JlnTa2t05024MWnkYiyhRAjWWXYCmRtVltvC4e+RJmLzoGN323FYrlYOheL
8KscO/N4v7I8jRtLRZh0Cg5puREWM3cNeUHzEG9rjpQaPlMUTjweuju4PmzW
OCWeoGxHbhnmLfxqDoB2a8/4OuWjL8AWZbe4ZbH/RVnyXBiYIXP+IwfQGxCw
PvcGinJqpqP5OC62kSUDHzPKfBIVc0A1HhhNfUrDt0V3eQHrNAuIjw/Z1gOU
76Iiat5LaGLdPEil9ziBoxh5wvotlRec4d/N7oHrWvkAvFmUSJwNIbDPz9pi
q3Q4Kuex43J85CHcAfrXoLZLpZLnmeVXd06tdd4ZwCQIycvoewXjxxg5qODc
tH3b51prwejuFANIdGSlzItBW6TUkgh5dYaEng8K2PTk66tebgWqPsl2rRUU
31ORH49m/L1K3y1m2kibwdAOjGn8jUi8jIkB5dyofkIROM203N4oD4yry1Rh
FdA/hpFYYxW79x77gCetYQkgHQkekIW+fr+pXEZuAtT3+K4AxkmFojhSWJf4
o7J+AilUUMdmzD02rxc+eNM2aEcyu/yU7heG5movVWJxySWb3kgVPx0QqMyc
JxZsDrIw+iOuE32MQQ66mDco1hmpff7GmvxThqoHUzF8L/ZB/OuJgOtxgZpf
4LYdnOnP3R1uwu8L1edG06dutSFjfsl9KuyspWWyP2pJowv/PCN1e/4nhEeT
da4p5vPqyCfKdVU42EhyVWtpk0Ei+nUWh09Pq4IucDv7djCghANPKuGd09lY
4V4IldygSiKDhjfuIqFwYoj6KfmhjaIheEYL31Ol8uzfbnJ6D9RQ2jGuPUY4
+PT2Gf96glo0n+mxaHaNXA7QvVI59F45teY2PoavZ1vihn8pYWp3uk6hxRNu
7FvbIdHEuys4/ZwTDZrYwnRNpJYu8b7PpyjY7wu//VEyiXQjJlAXU7uz9ZMI
/fEKvjXGdW/QGtMe1bcsTaJgR3mZ3a6FvQv1ub6Wmtu9qCGHIjuqeap9IKmu
lozjahdKgBVRMjw+LgxIF0HaMNWb2QXh0d9NsF24PLauAyuaDgFtgT2xZJHq
uNt+KDxbmxzc28wR7N0P6Rzeu9wHpwdN7dc+GLm4XGiJ09a6n5YsIaBBkFa7
3wMrKXBTlDFKoJc16PN2L8Mr7PP1yATeTL//AJEQ4Gdkk0LUX7/wj2Antt6l
qPmdGtaf7yDAlpUc4/FzqlplmA2igxRfrlj2XcN1Mip3GAYOS3/+PsbSABjX
Icz7aa0jUU9sd0InBQtLJmO+A7b6dMdbDdT1PKvCC9WeogpnZI7VZfMgvrXH
fYGxTmK61ge558zWsYsmNqzk7E5E6XmG1yX8PB9yVuCmbYCNX5j2ugzOQlo3
ZP7GfQlz3DAUUjnb/PM2l4WlKBZIjc62QC8+KZh5/uDxbVELO8LeMAQXtO0A
sOXG02ZesFhJUvoZ1Oxzj0WGJLkvMMFqJw7b/W1n6dH2XrauOc0vqwB2d5+8
UGk3YNESPZDTQr1aQnN1hVzjAxWxY7Ea7ZClL5DuAXJi43UMBCGcZQQXUGsZ
UlOAGYOiPbeBqoGXfFASOsSTV1iqcFyn3MTMRVwcapmIKD6+1x/D5MrxVNGs
kN4e4qb9t60eTbbFT9hNvFqZjfGal10x3YEsvIw0GwGHXLH5cTWzvw+UIulv
LhfUgf8ExUcmhk0HlRQ/TnY4p3DZxePnm6ImEeWe+5ANPhgQ9ntitWdtGzmh
ckHnL/8miLroNCXbQLzahgVe/HYPwnlIoPIcWu0l48UdQP1DbhHHWu9SZ2yN
/oSZhYfMZUDMkRqFTMbGk3TCzwSKPisZKkCSeE6NgW2hdjU0If+oFH89bNEj
jcEb1DooZboDP4Oqtknb89nB5H4wUqVMtYVUCf95y9Nh/zrtfLh0B4cloASW
cyuIt25zZd/L9VPks4JWoGK80jo2pogT2LBf8+Y/2PUam/oS17KEUTBE/IoT
oNdHz5g7qDOuGGwtPoytP8ZLxUkldZMdjILx5/Yvq2j55aoiazFzQJbCjjnK
SjOZFJ5SK+uI7JfeYbLntpxvSfY5eEUgSRSgoobfe3/e6NXAUuuCpGz2lG1/
EivP4g6dpzqmGEaeaV3VNJKXbekLzovlwoBPLy0QYlqEVe5BhIzsNj4Ztgr2
HHuL38iaN2pE+zhw4XDPKU3SUlbv2HMmVYuXej+/v4OH/gBRAClmpAdJhkbg
qd691nyXNrDmeFtH8g7iNLPmj1ftexMep+OJae6zQIu2TDlaqM73LScfuTLU
0aDg7dN2mvetCH0J61MlQ32U6OUMEmd6DHOO7+4GUlCHRqqCnaEz3nSlpZfW
G1pyIxPx8LPdhEeECGDW8sUGfgGmuJGvF2LwlrA9c1nROuDxoyfoyln7Ou3F
iqqJi5p0zvWJKjUqbvfUMbJma8+Ovaesq6RJyijO09PcOL4CcfgyBkfRd68j
+w5tUx5qpr90r9bd5BIoQ03an/SfRwcubPiqgAZGjDWWVSfDjgR2wWMdoayp
MCg9A5hdCenNJNb0IM2f6jev9pamIWJ2oMF7o/6WsuNlfsGqVb154nrXYBSP
j4a+xibRniplQORhNIbSfRw4cYQvIVL1rWwf/1w/Xbvz6WxFPGWekBun7Ga/
BiJjXlNXdTLWSRD5zezCrLt6T0YUtDIxYUWlgDFciOAufGV6Qd7bv/BLjegg
7ZSI6r0o7o46LkBXK2PDCpgObEGo6zKiHpT4R48von3eveS/+AwNS7/Wqs//
vbRO37ORonw9bcrEUIQCQGYvcfGj6S5benoPm2eztDzVV/Aj7uCXk6XgVTPp
7KrUuB4DNIICU+crysTswce4j1Q6rJhotRebzt8YxVSsSnUNUhe0zp0qRBar
BTDEhTuzo3J7rCD5FRc8GJifQyLw6Jn9Wu3jKpOh3zSUws2ZbHaCSTO8Cy9/
5B3gpn+b5Lfw/zIm1cfNTJzfX9Uh2XBVdGop2yA22aAffnPgreSnXf0fpluk
9luG4PUuFiYX03wdvaPoVWZ2pVot8hZWkXnIaxDL3mzxlnovUGauCLfMJbop
SahHKfHvIY6VJEmH9h7XJQ4DNBEUULNxe/EA9Zlzt3Q0NphaPIL1gB9Da3ER
fJEUC0pm3N2n+HvcNfagau/Htmr9vBZ4zabQOi6Ozy7qGT6Zdx2a4hfIRPwZ
JMH5JgWZSdoWRKOOsoi9ax7JhJhsGd5IxDLQIO1iRjKKwg1CHHEwOJUboTrG
OFxV2iDnzeU5BQlQtAtmGWqU/NGnqGssQf02tjs1wztyVh6pO3rnnOtkLM7E
R9wkHSqjuxBOCmPdip1sb/sQptlayLOW9UBPMwR/8NQANNxrDvvhEEmJRDJH
+2K5++HVzexmpXQ/p5bfYCNrOKIxJZLutGo+4k89OKeM1801Ch9s2ao2vJMI
PtPo/IGkYJcjm31ynH+X1dU2eKI4cKsPd76CIiaHXI5zLbFuvDl/Kgq61sZc
62JIdSDpsgJIGe05s8r9X5jp9BKW0PiH7hjP+AyN1Tp+IYyUArXDzcagQcEj
l2QPPJsGauPO6HI3pBi++9Q6S6rzNnNFO0pWVZFVz/pYpB4FqWIbj+YP/pM3
xnWAOoZE8//lS+OS02nBQZDT94zWX4FxKwUvKzyzrQye+oyLT7d4bWa4TLCv
CsbqX3NrLIJNcQ5OO7clbvU4TgX/rAmbtTOmuyw5GBiIWphAKmCSjKBtfF2C
Hz7NEaR7mqZKlQeHq9P03oEuwQoWp1WWD8owFKDVJB9l0S3qPkliD3C0wTLk
Loj4oIws25qXuiBmvKisF00qq1b/4rjgjZGNpRiuJkFGj1tXEAbazXBRbeJb
aW/TU/OzeBbTTDP12knSn1D2p0KULCzoOU3373LWnixsEi6N4pYcUKxv+KE5
ID3TJOOaOEfOUlB1Er+2Tpdx9DsksjVvrhizWrdHtdaGhNwd+JTr48FKmLrh
xK2CjGVNIZePtjhhD8TxfinQsFWHht2b1NYIpatNDo+MzO+xVfhg4nX5EKY4
2tLnZaJpdDr55c2Xxdzb8O4TGMMHib1MU4VwpVnpLyArF3kDP84axmQXoqUX
GDdvQqLc752/m+DP+IiMoZMYO3aYSfatRlcrOvwBeK9nclNHASlsDCSjqypV
wDQe+bnpmRhQusZFkjJJi/Ky1qEvLIiaPCJNJG5LvZo+aGMXB44z5cdjNHxp
xRe9I/btaKsqPGUNqkTQKvemRRJbF0EpoMSJIjkefcml7ROK4x/yarv8lsst
hSJeFAf9g4Pg/GR9fVXArGj+eqTkRG7vGpcP6AFs/VTS5igaILOH90+kgFdT
1dCy/jBiSVQ5SIogQ/X9XBNN9pCkDw1qGqADjSx3ufRVFix0/sqReqcxr2ph
/bys9LCHWVMxgQEPnZCNc61GK9Rq7sMu4hZbzZ5fAMpRGhR+lyIIaqYjSiYO
TdzaqENlTlU5aV4lZ0g14Ipyimv17zwRSQKUt5RQbc8WXTbH2ttAkzxc2z2L
iQBgtfzwsPkDmVlprj6hg0kd9QuciZmoH0uqvEFW2yl9Pfw5XV2f+xjC1ekg
gYlj5Q3fhc7jz6Bp/9CKXGGCPNI46jULxvjX7IyY+H3a+TTi1q/8UFE+Kgko
AoT9w/8w/+zuvGecYa91151pTqdoXyzdCI8EfXWAAb89QGiFujBVTwGt8Hth
DibqKtst0XqJV1tif5SUstDb2YSjmukKc3F/Th5wenVb9GeVioCIr4Vc1lTB
klJ2bS1FnVldxZo+1MFClDrDrrNTd7zvVZsJKef5IH30ordSLq0SrZJlOdIc
J17x5cNxSyNnRJruF5BiQX7egaV/eCkhXPXBHTSMJ/SgMs80dgG1dwOD9OMs
FZtw0z6IIrm1aBedRhDhAsNnQk0Ga7u/1FvQN3qTR/cKOQ/ICnKMbeXS99MZ
VOmszSPoaFpvjW5eOoUOvokvbh/MOdzsXsjja22mMBMsYVUYzkIh7sLuzU6X
SUzcGiHFnTdknGE0haRLzKMpdunC4oiSqnijO2sdFadbhBNI8WM5Lk68k/zK
5U2pR2m4Gf0+S2mxE7AvSfqWgzABN0SYqGtGc3sCYvlv7SvzudgoIx1N0ZqF
JSOg7oR78t9wkVXUFKwf5khsFUsuKCaJ2kVvxsALaJglzCOc61qqaBen+oBh
nPWAwjcWTdxuq4FSJtLFj+Hl349a4kyoEBfIdJt+9FFXYE2gqjcwN5+pglqU
E6tu0hO2s44lf5kCDMoAmOKHvsB0FpyIYqrkcnOLVnNTCUBoTT4XTTTzHLtG
jnYqZQmON93t8HDDaViP8c/s8q75xxZUsZ9wHOIOvYti69nSrxGdLqxkDMOb
+IEzZfgiZc3QS6oRCGLuolXCRatJmkk7tRyJWsEU3I+URXXpSfrVDbSBLYHc
WEHNpCBzAojHkDqz64mH0Tlj6Z8SSqQ5tS9V+ZaI3FWTaj9RgBNaLpu4m12b
x4DKYQ2n2GZn/tdlNTKimxjhis4PtMQT0ZcF4+Ez8Kl1XXqZMWLr0HFeJiSE
VjEWuI1c5VUaTXK2hxROoEbEJiuDu934NJSM2kYpUCaYsrWlbJBI6EYNZJd/
ZloeKqc1gv/hxZimDcSmzXTakIw0gfJ5nbwusFOfozs+HsRQnOIxDre7TKvZ
0Pg4WagiVu4TXZkPmegFc7e9CTfozTCyFBMV64tDo7e+HfxrhJXhP+W07dEZ
1SCpu04uplsQ8VfzQlhNLnUTRUg5OZ3plcLcfkZIXdFl9tq0H7FKxkekXw4H
PXU+xp51FzPY7AzM2RjpYXCXyEPBGmONGehpGgUS4tcrMW9VrSpkp0bSvRmK
AEQmwc3JwdGSQuYdAH4UyCeq5/d0ZQM7iq6/r44CSxZ4Gy6boyrzqVcjArVb
nYaIRppy7vYfwCvmlS8KkTTcSZQBbbb2ZaIb0GE7/b18zJPU5H6BVI7ELFNB
KB2Pv71M+uHPjJJZCnpHrdtXni397g0GD36QPyUdUeOIwcA1lOjj59msrzW6
3jChBfPmuip+QIIttrYBDFP3OLN7cagIPwefB8Kz5oZazXBTeRFl3XL+k4JP
XdjuXNVBYGwIK8CG1DCWznPmJ5ONdbpxMVIrDDahYfnBu/mggnuOH+jBlMeF
00Rs759MByKSFEE79i3KLi+BXD5bkE58ocVKE4jlsyxflSahI5HhpPECiHlx
BZ4dOEcJT8TuScDnBMQnwobjNQeD9LsZsBduQrZy7Wgt+uphRkCs2c2kBNHq
HJoWFaPTnix8YmqhTHwakuD7ULR3VIuDsEHCpVMdJUrR61GrevQV9MldWvfv
EtuUMcirNUiqBJ5AGmPHmkvRpSWlX6ozBGQ6px5oL37R4QcP5DEwE15JXM22
h6rhXPFDb1W5Z+j3OXPmwJk8kWq3ajK/XYfdUU1HdT2kSx4I319vcpio2GiP
7/fNCnFv9UH37sylVlD46w1Vme8NNlRhe6drr87Tl80jLE+wWZcDGo/aaKDa
d2lvTNh4TYJcN1jE5xyfMmpDMXzVduUemZJ/I4jXiyrfJyaX8ZYFjJaX4Ljz
tjYfMh1tkspRRATgEzWjyU6Y5nAaPYn0B5lYG76n6ngq5pbMDptRNASniDV2
jmYv2yVbnq9NJafNOWVvwA/KBL0iwGm1TM1r1/6Zl8RgKqqp+WntlQDAxewx
F5LszsCnpyUvWQtBq/WwTSxthdlec0fV23Tfrm0zBKXPaF8NmBPa1kXi6DX5
O1t1e+5vDYkvy1Sj0IFN8fksxoTfLr/ptEE31mkq4NG6a+ZnC5UUGRCe/qaA
PpFnVnrrK4BHyeCTrIVRoj3N8uvHJO5Uv294b9wQqQYX4qsGNdLxW92tsgzw
PpZd0kMZDLxRihurkn81UwgjE2i5C9Dz/z+WT7ICDM+LMcw1Ec+mPYRSjtDo
y76J56l2WSgCdimr4UvJEbUQ1p4PHJ/yENa0mDMrfmKx6sQIwhE8gtzqlVaM
BfaR9HKMxtGhGaFc8cSOm/r/9ppaLu+9IblNyo17Eils5wocI8hMuuH37rCD
8iDKVhafY7LuuWQo2U1I6XSnw/H+tKWX8KCYtr7Eu/ZaFwQvRlCe3kkLMIm6
JQ0IdR6yhDC6rJnQ7doC+q3rZAxKYxNtU/BbSlVnExF8HXbeG6aW5bjfmhi/
GOerTSjZW4GkEbCuUpkJaZRSmlVEpspQGNGmeQohN4DHAG1pD/OYtLiGdIUE
gpfUIkj81qxXiTDXBh0kSSiHukXPF7RaDspPKQUQV4uV1KILSpEaH0N2cRtu
7zOZP0rBiQC9cQIy8eh05/9Y447zW8Of/31Xd9evGs+NLbx69700MPL62gDl
zrmQb40NAQymn4uDm3+8mloPI4gThkbuwtT9+0W/eHj7/vQ4jgGLm9fOK24Y
S2L35HicrlJLqwgmkjLcC/onl21HxWiEfrBHmBfvKmt3qbTpS7udTEnKSzAF
v1NvQ3yDGFwJYx2V1gd9QwUaLJceHN9Ty5h7tKr5gzMwX9fmXVt99ayhnivR
UJy9e4I46aDV2VRxod8nuJh5OkSWQd1tBjn6OGCu/JfiqmCpcMeEPAaBW/zn
+7UvrCveliMF0nre5MZCMk53LWAgbwvsgcoa+N8+PxFTmXuhBhaJB3rd4VDk
5bhDKdpttFEkDNDtIPoKS7z/hKTZdNEc/WxvwTn6kT0yoNsSnINzvJqcYtsB
nRT2aors+//iUtSK+QcVv7wRRtNjgnX8jt9Dn4bRFKicIrosWpUXLzHveCBZ
g6OYNW/R2ueRZEp5wscG2UIZoJNblpcsUcniJ9qXZleV6GtVavzx/wCFCPOZ
Y5KjR4SOm/hw2woARzjnli78e/QF40CcvauCvEF/ChKW3TTzr64t0iRFtTpK
rePmPeDY3yrffKY23sIY6cmZ+jomfHLkUPsS+D6FN155Pa6sL9C3CL0KASdA
kvonDmhbCKlgLcF7VucJay7o3OHLLPEJ2/4zlfbtwI89zkbOedEPEhLRLvCE
rByGmVrIucCtqZC0UYw6BbXCTBvQwUbAVGcIFdrqwNVAXIi/d1FirEIk9tY3
kLhPIE8vOdxfMB7uJ1dmIuYmCcYHBOp8Wmg2pGK8F9JHg+nOrAN2AVwqAvhb
h1vzfBhW1eYu4IRxPQX87LzeHlFdYwDV8jH3LVbqUiOfnjMGRgwwt/N9KGsJ
5Y7dimTSPbr4xcC8rwcfyhnu/RjeTdpW5NEHwbDSx883orROVds3MW3UD8Wa
BqYHykjSE1uZBAHIylIt8kCME+H41giBNLHmWTEwfCPWQIs67MTbzyxjPbyj
ze5BiVaiJCoz7GE0UwGn9A+SzwRVYxxCrm5oHwhyZZv6XWCuG1QtTXHjVUiM
agZaFhjXk075rkcDK7p6rP+xW9PKrVyrtAbNQ/83rkPReOYmuwslGEfLAN9I
QszbMgCFZ1u5xU75SeSWBF4imW/7kmCtGd/sXBs1asdBjEaJTRFCbW1PzeLH
8tQHOHTiogEYaeYaytY1seulVK0D+UIGZgAU6Q2iEnrTE1PaYp112bEidWqC
ufuF/DnvwtLcX9oi3hAqORNjNU0KDEe0DxH+kEWn91XKhRV/5dMsdFxg/2+N
D580PFYuu9UpJUe5dGADKOkVExyseHcDw5bl+jQQEdOuJxAFDtoGugZeC1aJ
9O65MHnWVZ1eAtePQFdvUERFY2KCJPme5YILHisq8k+nuqdSw6rVEBBXQBGg
O1PEE3Hzo0sT4NqZ44EXMK6UKwgk9gwxCP/WoMGzu+KLd6+eiCSbHJdPLQZM
k4VC6VEspotw7pHCFp6MbopMs3wr9TIPB3oM/2Ao8FC8jdOSPxAqx1ATSsB0
eNxwrxvVA/6z/9MLzVpdMUTo4bQYR0dL7Fy9A60yQz2FFQjdGg5eJLR1YqlY
9PU09sAZf7/Y+gAFuJAFoDwKsyqGpw9zbDPqM/MOmIEzh7TRZOD8+PBuoF0y
Vk52dB1Y+tsXrArp0+stOkrOurjF4m2AoMPpG02SCMEM37s6ves+4KvIazjk
3gPpiXCayLmn6zbkMEs6Xe3JnaQ5wJMvzy0MCDRk0Rbo/qQc0Nt+noT0aq6t
ZAVRd/knBTkzAl4iGoa6ZICZ6NQr2J7fIM8yCPk4gL0VOxZfcC+fY+2dpOlh
NS5vBnKVfdiUXEFCzui6g/BHd3/Vli+7tD/JAhYwdLJv5iUYm72x3u5XwyAc
c8SuiPNj+uM3YsKPAKunHPAh1/cxYKJYai6FLAgGHpbZSFqR14JkYh99RQPf
oFxBn1NVbmvLdpxWG4RRYXrdOf+rypcS0R7v2PlvI836BSnllqbIbwebt3SH
tcG1Sm8C1i3V0A4V4975e5lSAJCTpONHT6OuIu66kUbqB3WYMRPj2iErpBDn
dt1c2VcTIb09Oa9GCDB4TKevJi04/T5notd1HRq8T2fnc/luAw/LT2ihzIUg
1D965OKlYAS5FxiNZvB17fP9ddx/zR53zuylqaa0krkJR5S78SM3MJPLap3T
OPib+tWlNsEiFJWly6jAtS/EtM6O1PXUU3hCFHtKXyiEYmYrLSWE9/DQjDNh
DLcIEw8TslYfxjV55vUzWn70Z45D8jsIr6ca/5sQ9koZ3Dmiz3G+tzEJfoKl
lLrZ0j8V3vNjTN9JtJtLmzHhHQjJ/EsnDjEQD7YUhhXp/3Emxqz++INBl+St
1V7zU73ddWWI6bGvOqliKhZrfDC5mFeST3Ipz3tCPYOIRLA5dJfMe+1kGdVg
3/Mk2Ka/Gf5EkmVlc7Pk47N6hQ6jvKqUQNNBgQ7HoCLrN1VlFuqKGE7RHlb+
1U/WoaGk9GiOktf6NIyLganVPTxZZSqbR428IA7tfe0CJaFZ7TmQo1MCVCs+
bXB1xjdJ6RlEVPxEG8yrMjRK8sVVGOjXpHdcrhjLMkelGZ6LeGqO9TBiT/E2
7YR7plb7l6hWt/LBbFlZAYYaTkZItToDPVUB20qzkcezi97BMcJpx0WTABrr
diuAicutdMvtfgBQJRaAanr0N7Q6RvRrFRy9VfWixo8uqDhDx+whwhmHLOjq
OfnBqJn+ppWNCHI/7ZYVTXHSC7tLhXKvHOKj0d3F7yh7PqI4Wbo4pVd3HvCV
IZb/OaitrTNKb3ysjMrghzyz/kSDtrUGhg7RF7d52mMfAlpbWqJuvhiSMVpc
vZVS9W9ffCE6f5gvbQhFi34axGyMB08ISTZI9zgCcoQ/zwJg1QwptIvuYY6x
ZtN/b0tKU3ozw9/WIbiIWSdfukQFiD2//ZmnKEIvAo1Py430CeFUF66+le7P
FJN4CkG13RjgkZZVncvJ3ujItfKOBB4mmeZAD09Win05ZhKep8Zi/mr0elWL
XU+TQWpgwZlLxTlAVdzCy9Qn+DA8bhnnkNQt0v3xSR/JXGnClSQx88oqrZay
aFZnFyHYe9Y6E9oey0P/6V+tCFUToZ68JGcyiCOtDldfzuTYUBRkEQkRapA+
1TVjwKv30KJRMhRGt7LbNAWVFdW8C80MjEeQ0di+buVaG7GjzpK6KlfMern1
ehwp0yaPJR8rdch0OxElGEr03S658JREERWlu1TI+gU3OKzsxjNajnQO5odq
OB46YlkkHqaAhskvmsWtSrOu5L76zQWKHm+XkVKpjH+avEl8P/REl1Zde1O2
UH5RaAiDbbZfrcecp85E2nDpyC9NVY0vt00VfIkszBmzH6REEXgpetodOgYT
tNTbC7JVbSYsl0s1njkK5ulzH6e8Sk0rTJEfks5u8Mz6mUTHPg6dwqNUJVsG
99wTl7/Lc83buYp8LkFZ+ZCyTO80oIH3M19qIyaKnYSs7GGfZ3WuZFa0zTOr
XOhaWSmw3OJovKDRMxIWgJD4hXB7ig44B08cSM4k2nfclnKfbkWZ5r5XSI2l
G0lkEiXw0wNDhQi/QP8ycjwLyN3yIvo+o7wZ80gFw7T6BshMcjCdj6COXwi+
L2GQ/qstua1/NzUJUSXBc0z9W6Ygardc7b5mhXOv3wDsfaTbw849WF4zcJhp
pzHug9d3jxvDB2XUDz0uN6TGR4vRRLEWEH/qOnGDN/cSXmP1zg69eXP1Stox
JIi3bKv7UHPHyKm2PyqwWX1qntMQqnc44VA6uuJ5wWfgpqUYKxBGOM3G2Bb7
cCLCrs1x4eiJjY6Whx7f2alTkoZlnG0U5Bi+ueNuCRxPg0DGwigLLDz1odvY
UM3KoQpN6z91TOoIm4TNJefsS9e+P/ltSsVVEZNfSTBx+wjSVX4zGBpiBVuu
ygTAgbo12dGP+iLu2ok1Pd9hkpouYqouVhj+pzwq60ByS97LPS1JO19jI2Vq
SIwnebGYOdISPxpgw/ERNWpvsN8CPCK/pPWGxBfF++TeS+EV4WDaWyf0Vi+V
rACb7N1Lkoq7kvsDR+reKn4urG4mMaaaEjmJTcTca7N3MZ4QqpZ/jvUd7ObX
R1eursdwfqFw6cjFeMVkPUlk1G5iQF87g3QkBPTW21raaPyoiei52ikAAjza
hRa01PGaFWAVwQUvYhu7jsn9wUAxMAiyuaK1/A4MVPEw3iVD3qNpauM9bTRx
vNSTAsBUHExb3CNkSWK7xNVmXPg19vaw6JlsUa9ThLbP7/sf5wE6CZni6HM6
EZTADCsuONtP5Nc6fD/mAOFT9UbXc6ydKYRoFu24hPUn7tMbkkLNwDLs9RqC
gwRqTh8aWWNuNoQ6QMU/yh9qRPcrwnWvCnL0ClUiycGOZNelZ8H7ZQzVdv8B
xXlcaVK5muYD4v1rjQiNtWSf1D2H+pYQNK7hnyxhrunPE8fWiMJLGBhcOPAf
EQhoho3joeJFtBTqEgVW9rkn4TSlhjQbkfmYtEeGU8MNz9XlBMWrpNufMAt9
kUu08R2GEX0vj+S19/52eHFoB8Sg3Cu5wKZ8Zje2xWrNyhbNNHMgt3954Y6k
D5VnbRUn8yUtgMHPqid7FMkwK1u/85XNtJs+ZCUGao4NCajbI7AkqA+ztEkS
LoPLcRnxB/nD2OBIfLzM59Zl0vXLW+G2Xm7EzaUXbdq+TX1wz9pC04ubL6Je
8YH/FTCj8zd7nbiYh+B+vgjkOGA1p0BiMHlrbsIcUfM9++pBT9Pycpw4OCHb
ES8+HacQ6xIuZK0x0LHu9jRJCZA/7xBCz8rJKRifiY7X+OMuUNNHJMeAvCrC
n81DVe0I5w5hLb2xHd/HTd7dEXyaIVBG+ndy+AGKJok3vs6giKCIgubHfiqw
XccUAfUCTLhZE45gTISNRlkfl2lHGlpzTaiZHHNib5MFckDI1LuKGjQmu4Ak
Uo4/4x2bf9vnNNrMzY55o+rJ32yw3HTUJknWH24WmZgp78Lc33f9l5vRMTwn
mXUVYGR/37fUvj0PdbbfsMHxEoBwY5jOBZxptH/bIGFKYOynRFUof14ESAcO
Ki/dgYJ0yIMkSoyhBfVbqMnrg+P28lWLy8vKH2XveVb8B2l7D1oMAehKcKFO
nmKIJ+bpk7P+Xn47eIGDfab6Db1esDrSSroDOCSHXZ4PMm0DotHj+J2S9OZy
mRktlWUGGlxDSxuMXHtrreZ9Rcj2p6NVz0esxFn5Z6iWUu4GPuikXnQIWLEX
ygFW8OecUFCYKfQh0iSSEzURm1u08R/8n5jDd+02mltsjOb3r8SA/RgqAicY
fuvTddMrIWuBdDbOeuWQ+GHb4izL1hvHlz9+va/xXAlO9Wu5rBAXNI4qvD5T
sIEnA4hIrshN1sIgelwff1PVZCTDhI0uUMqVi1xEE9TLDCKcK5DgsO3WRjwJ
WRYY5bGU3Qkzfr/gLW8FfJJ4RZKYU702YeZv6ge9dN1JB2TozAo+r6NEZD/k
oeyKIxHFInlCVmGxbLC/arsOSLLOfMsLuxRyUHtJO5cOZikAFyaOjRB0UFV4
yCw47hdfVrLUFaAwNd2rdYsv0r+vJLiF521tRB3JnRmXxsUZDKyZ/z/O77Q1
em4vFn3Bb7BmJoAb2YPxSAe41oBlMlpFVexBf7VsawEJa780TGFz3tmHBSxf
oBHo0zfgSjdz1Fx8FzFbEgbm1uhAmfQeBQ3xLk7hOQIKCUavd66pcaMX3PTZ
UjjB7luL9/ZIYHTWZQJqTjfmjRAfNLe7c4QnXL692GMUH6Wj6z03Tui3KEKf
23blUixX7oDxDsfBPoCI3JydUFmsGWZPpVoDjuD+fRZgdFqCT5wAloNvovkM
B4uDs+4N15RO4/SH+XH/W8+F+E88/fPspVaBb2Ay5fohvQ8WuwGL5zFYp9ch
t+AHpXV/9YxU3aVwpkLAJx6jE/N2Sx6lOHuJHgDONYbTVb6ujdKD9BRFAKj0
wECllat1WQqDyV8sQkf+k2d9hILkUbB7R85IOPnJTAjw7FinljMvIAisBUv+
QBF1Sljfe+jqQsFQ+gaA00NUqvCA2MOGSkPiHfUsRAg4jjHr0IVxwqXFy3Dy
MtvX6zg6pCLSIlucLgImLS00scoHba3sRjZCBzAdjhOuJu6CPlAMn/EDgM+C
9arPtdmGlgUhkuxN3RHoeBizDgpYa1Pi9LSCZH7iBkGEmuKQO/5wgpymUFXy
DNxqdvX1aWNNoqv/9X3xV2OMZz4QEFB63UIGyC7hOUTRfwDmgeJfU8Xl877H
SNe2PrmZTrKBrvfQAphZOXbztuGuprvNOowmRzeLebB1ETE1O6qOqTqpcSXy
y6TScPxIbcsCjr/RucKj5tOvolqeufqCBGmcPaYv6OG/SNTvG61t8eYu9kAS
Nu34phEuiYQxi8O9aDcpoDRr+Rh8VV3eQlmwQLoArvE7+7fRWbqI7iidVOhm
SDIZbadNh37cEZ7QY4H5R45HkgKF59LhNoTB/ucjFBWfFjTchqpw7o19hXUq
ioVKnA1L9QpFFam++i/y/QIztRdTkjSvl88DAPTLlhEZdoJ0iRbKwmeiEdsu
pEljTo5Yr77WCVKtW2mreTwHiTJCwZQa+Wgfi6X2meVXADNfDTsy7v4TRVaM
A8qv+1du1yOFPp0COSw6J4XeBmohmOM2tcpPvWFhGbUw8D/AiEtOr/3NXqzq
rBNCoic4CRa5wtj1+/YthE5TSkniZv5VIjCRqKc7XQgiO6VCzAbnoq9SfXSc
o28vzoSUMsl5IdUGm9AKdtI8+C1vqS8nmtQCZbDAJJK1P/SqTQsNtEarlyS2
B7KHhWNqdgNzqRuCESWC4PJQVHdifrrlGXroNjSdAcQy2CUi6hLJPHo6k8en
OoaRcQ/MeMwgGgtgjPalfiYadHGXex5tzelSxBBjW4KNHIeQMNYEG1znGOTB
98YANh5vopK9AMdhYLk1L+ShXQ8oXoxUFMaMV83SgAfniEANLRf7RGAG1g3b
YU04aO6BYuHowUcecQ2fO8Z096nvyMoL61cSLb1ukBWgSNe/JkRJTGMWQIeb
47AqhY9lLnc554Awp+n2TjxXe7br2SL6jlI1aPmVrYRaCcFZqjfe4mHBSWAX
tP52EnOh8b+JHf4VX/wsw/5m0PYCSSk34TfqrpqlKIITkDUZ1T81OCJnDWjE
6FRgsBLR2bKBzBgfEbU6DeCY5fDI11TdrvAU1Q75RB4qlde8tmlcfLpsxm/b
tUUkiayA6uxK5NySOfhkVQ+6Pkd9iN3yFaoKqp3IXTgHW2cwAsbDu07eQAWN
ZbaVxP0ZwOzde0Ig7ypQ3yM/fX3IBos+eBMjmTg5N/2b2gCjbe7adbl2zJug
V23DwOVy3jJYQH3a/XIsrSAHOSixNPX45gO1V7FP6Klu/uTYco5H+5KKXU8J
KHO+W0ygoBEU8rs6W96WmiACKEER3jvs7nYnpVnJvaCNqTrO5O1CSFRiR+Qi
6iJX3Z3sO1OVbWASDvmKWmjMQmZth0tn/YbenricY1VVSUXc4i43To2atgOc
poZfsxlCo9rUf2OyUiPvrLdjHG5HnULsI/j8jT3R3F2elQ+tXAS61WutlTdI
oquw5mM4GFbMCBGAzByJOoZ/y3qEAGJ+LlcR0Gih/LrxXZ9oYeft7xxGucnR
05mp/dqdVT0fnnjyh9eX+IFCKeq3zssrk5zCVVRCSG1HxH9P/UjQIDZmRxbf
6BYHoMvRQLiKnj0Li4a7z9TgqxgygnnnpCCtSG+QiCy/38aEE/lzh6db2n4h
MsM0oZObro/vzHWtelWzvUltBw9EWSBRYmS/a3TQ4c7F6LQq9AeC0uoypNun
9SehvSgwr6jiSFJAiW+0Bpu1E/qRAxjGIP3xzl2+gdo2TTpoU4xOF4XZDq9F
qHTjLTT6j2VbJliT9FFbBWu0qx8E50F6B3E52zw64CN6PYtmF897ZuIHCoak
Nb4fA7sdyTifsyLlrybl6zOqGTkEJq2L/r/rO0kOd9vmnpqPqEexHcB4UvhT
dKZhSAspAyazFIxAybU/0dcs3BCfxzts2+dA4dOZuysiKQD5xC9QY/95yj+6
uvXLxky7gn+fFMkedNvQjfzuvLS3KqaGCF0GRnF9Es1+rAnvkGwTLr8wTGpy
Vf1RWj7j9zyuRSrO3uya0XabueLK9gTWSENZJkg74PKw/YgISoQz8pajCtrE
+JcO4w7KyR9+AOFxUblhPn+Q4ZrWhvP+lMdDcshziWKlNQHeSjLBdXkanrsp
2U86MTNEPtmbUE6PDifWKhJyrrLBxsXyHmeYy75zqHYXmEVacYc99Huc0yCm
Eb5luT/FT6OuyU8DGXFHbwcvRHTcAh1E0HMsZPxvi6DAIgncuCJMUjJsWOkV
aYOGU8/IS1xsDuenvcwUtN/h2K90DDkQgU1ygLrzDvZQdTdrv4bHJ9q9rMFq
O+l8QwfLZQ0HFhTA3RKnIklS99zsNFnv9xdkP4z+ynY4qICqC1tolqyhGxiP
60a5OrYJKggyIN/2spCY0ZMvfyFfwkCnv58fttMQVfeOisqr4GiMGePUCqcS
s9mzgLnGpodGGk+rI4qb2Og4r1NQyNToF/PflcOqP3kIvlE7u7dCnEaED88Y
boR0VTMPxPVSihuyPeW8I1PjwopITyrVClw1m9LUVbSU6OyLQxI7PTPuclrz
QZMw2WBt3XPdehznyWkVYVbYMM+BGVpq7KW6387A9md6OfKlRRre4V6e/ys2
Ys+f5gz2qXaXrWv0bStvEa2CYm2fBLeuvEZXbqlO7l1heY/lO4di2YgQBRiy
NnTDsjLf1v0oPAor0vpjy4sW1LAgew4+nuUXwCsv8jHayDUnrGey0W+wsMsl
exMna4MTljkLveKndhiJO0mvpmeXaZuuRYNVrR0fFKORSUbGQ3NUzNGJRILH
PxyFwBuKAgukLZKXEDgHPnWMqQ3TbluY+20jEQKhaQdb88q1SCPPswU04YRt
C9OVwhIJ6Ip4Lnzh0X35z1v15nSs4gJ6BETM6KGSZPbhzKsuP2Y8LMRJCgS5
7Kou99dIpKf2D9IbFVNmaSaSvneIT+CVfyudg5ZjmLaZVCLPOrvCIg2vfmfl
v+427k6wvfe1TLPsLJ+wKcxK3e8q/nnPfMqaPwNdc7FkB+8mnnufWoFiIWz4
X8DXnDP3AVJNSKFpBKlNfxz+aaeV3cKBIQiyqvv7dXrBjgQyXwiU9xs61S1H
p9p0jVFkFH1AJVaNux913DymYdAx40dwKyKeM/26yuZFFP74iZGPi6ZY1617
HGcX0ZlBCbVad6ONJfPca12KHfUuFRhcM7emqT2nDCbLZec6FCgfm5pv2k+x
KbXXHFUZ01nUI6iGkcLKwdJ2s8qTphmujBmpMnswK42OPdFRgHrW0mbLSZqc
3T2JaCho8qFsz8kpHwulQ0oKbhcQVoI0ujbhs0I+OMs9wFe/AlZ/0oj6JoYY
CIJd942YJhg9VxmdMKBrITXpDysG6OgwIOuy3bcQqDOs6HjJwoFUE8Ig+BJt
ZCT7PRiYoG7wWg1YEjWMNMJEQa/lyUQogqZXuOPCVatS7FAjMrNOg1nMHejh
0xiO61xJTJpWuo0Za9rOdcyO0DzOk2KZaqPyDJtYkfhO+r4qt6U60J5yOvER
oAQrdxINEWgzHuyiM1Z18r0t/yKNMkTqTWuS/OnLjYCpfBF+yD07yioTx4Ve
xtgUGmrtKnue904i6uyN6nDUnO/4j8vv/XqewREFAY8PTtg/PYfJO6fOB0/H
uNsLcifAtEx43UqkS6knZYaEMnJabqEuV+Gd/t9uLmf4LD7lZaMWAuk+OXl6
fvCI7LkY3rKpvoQTZ/+A4DGid9CRaxMoLrE0/iasSjHWzmrCQ6nucUzVRNlj
6MbGBkzC3yd+NlFDj0rEIO0gMN3Bn5ZaCuOYe5IbhqudLbmCRC36mOE9lKui
DDTHXo8j7diJZlKyHVQEX9akZ2LUISVLBc7kRJKM+NpMsaRofFaef4sH4GKH
KNOetGKYz/sdkaGtn33RbKuiJ9ANlWUg5kk6WpPJjBiIpsibOjdnC3nUJmNc
jZHmL8Kl5AGad6zQEQFpVh4FU8W6yFqop0b9yV3yDDCWqok7RWruNcBbtyN7
yFLw1sq3bQ6ouUHK3WP4CTnA0pJR9GzT/4y9woXKAcBlKSQxcSjEkS0sClDH
tW/Oy74xA0cLWNnEdCV9VxSRBicruXGwHbOjaED7kdiJwdI33MHiFCxD5Ctp
c+FgIpyrRlZN9ktfbI3jFl8R6DoOJxu8/XdhoAvp5ZraTf2yujZQ87rEbTHL
j09ZSk51JnOHY9ijAz2YFoltqN+84PzX03stT8NxIG3TNit/MVuaFC+bxvhl
4gnI4W1T4Rp8h9UOr+303OGTHKfjfHTpolgCLhaUGnJSrGwp6bXITmdF9dyV
zmt2qRiGXteMeLebEqibAMo9egS6Bq46HSrwgb7calCOFiYm69OPmYkjelcP
befEhskQQzhUasmjcUBML+vlZ0F04K8oE/n6o/XBXAOtb/IMNpgI63opnftd
1NhSfn1xwxHCQaq2bZQoTZhaC2559e/6rDNwa1nTul1F7zEy4+BEElFkjOEj
mp061veXcgpjYKqLakMiQ6xIe80Qf4rcIvQF+htHyKHrEbyoljN2H/zxQq2f
7g8T+50zz7YalnfL0tMpH224ep10LjTpM6sodZuJfaAlw8u+YR6/otuUHDjV
oPNdX3X/kqS8GGoged8srI5wOfmwpYJzz85xYNUJL1uoC5c4IEe5/wONGqp8
KL5gmeYnGA5f77ivjAfphOfIYrtEIDYNkjJbAOhyttEs3cKTqVSJ+QIEdqRl
UkQ/hznSTY7rw6Y9Hc//BqO8OanTg+FC6Zmb/jmFAn1Jak4cJGi1k19RlVu1
+C1jps5Zhi3wMEzY2S7XvXBilkT4JnYz4uCwfuOuHcmPl62BjKWRRvh681vz
fUiGANSojxs5h9+7mYlXVWpRqypX6/wkxDEPpmvYaW/WY6qzoXrr6akh4NEf
ik2pmfskBx0zT4hfGAYiCLp5YWVaLkWl96DKAF6asOAC0KGLPh8liV2VuQks
NLQIHBYEqI+Yp+j86YTA90rp+YjpGhhYkVJqdtlZTmo6hvfezIEmKLa8ESm4
T8pM953YOUYkSBPnv6gW1MM06J7Mn1gHnd8mgU4odc8ebd3k91V0l8+paDM0
f534nUj8ucAONOfgpqJPZMGh/ml5CCS0Yie2E2LNt65Fs6EOLzpMgLP9MOmv
w74b/zwU4fAXApB6G2U3fGNOzhUDvdSh4H2krYPdTqfruB67Ehb5fx9iZSqP
W532ixisjJnppwSSRf5VIKRhu9JcOsD8mLvo1Ht74hhrbozOBZ4a0O1Xhidb
FPQ0INCc02LkPeSBazt1yrfSS71sRJzhavamwkayXX1hWo11QIaXNbFPRHbl
prbLaD5wF9zk3tv2m6YOHBJ4FQKM6uc0us/3mrWzi/NsfLgJKaBzcqNPnIKV
U6bSvIWhKOaLiuQQWyxNUhlsCWrnY/evXZHABBrRQn09JvhzFakDMtgDQPpU
8AU0yq0kYaw0CbrmJs9KTahhCjqVI1q7gWsX6/iDmrPDbMxpIyHkAyfJgvVZ
LwRx+cr1sLWKLlKeSS6VmqF0U7FUPMU4VY9AbI2QbSOVzLxuCg+iUnCvrfEt
C+n7U5L8KIWw5BVd2m41ggcFGfRAcWYN/t78CovPKVuCgAIkO9oWduL4h1nY
/pf2kwjQsoYqQwM/Lb60MyuZOi0PAD9mah2Grq/ClVPLx9mkiHRgz4VQ4V9h
wIltudgZVkLxkt1IIrmw3odmwIMQ3y0uOGcfeFWnnddBn3eUEpHCp79frhJa
g4fmUO1HobYsL7qD2GWxMo1gKKOV7Fjv758BnLDftQhX03QzGSQnNA0kNn+Q
EZvFtHkJXAa+wh9YnHtX/WckdYChhfvDL1QV8ZmQIZHGfiEKbDHagUM/6wuY
CtZsgclQ8XrNCPdaD70vFzz0fL1dJPy4ZwWvQQHGLkTwrytMF8LkLEYGw7jh
7h4GyhGfFtEwCqq9SfD5cfiOpzc4hrpaPKLZ2dbs5h+MB1WdS5M+1T3VzEvR
oxfwDJSfzRmViWNp5JMTgiwRznibtd+zsTuFtFksvUyvBa6l9okB1M1wGGKx
7rH4OP2sbtJmJiCR1AOToZjLVBEcMWOnzoxKnDQ3/irXJVfx0C7w7TnMHL0X
ysEMgeqBVT0g2u/U0kr81kyPK2CYAcP+pNtYAMf6vLJSJ6+QHI83SRIIGpXA
veTAYqB1g9k4NERjKqWksfPwGEICijlCtgQJe2shxUBVjs4g6SAgKFbU+M3d
iqtOSpFjAnZLzCS1DxkGUEq2d5Nwx+RHwACYH4WgPoKB80+k/HIleqbPaBJw
7EJ9v0dq8o17C7mShvxXePaHsYZ8uJhapUohs4B1aJLSDLDGKsxlcp5J64oh
G3J+nP/4CaZgi8KrX+d4UZOu/ZSVWd8MmMwzc2fKy6v7fM7g+cQhhXV91daZ
YXoOVAx81B0tsKeW+RhN/Mb6iE+qtl1g9PSbCyo3AMseZy5dqx93S0IPFHg6
OTTz+XhpS/ZP4uODfnnfyQNP5NYS4abYeuv44mAc8U2tD61tA22jH4Ca9E/z
eYFLY3s/7RPWvGiITAuaPrQftyKTmeSE6L9n2s2BGzBZEOiee/yx6dSpIAmn
WG0/3PapWTfYVq0SNhgK3VaXhBjAhU5qBMHZGLvwNpY9vQJafvnF96guuVTg
9mUV19r/0SMo7jeIMs2LZKnWK28LvwuCv/7hx67ZAxSIXxZko5+w6lMXkA7B
gtiHpQCj05euVv1WU0y3/tMVP91+ngNZwbJ6ptGTJ3iZZhDsxI2Fe6v+RlrX
08f94VYCFgoXLPYFuDmakIiMP4qHHGW7Zcd8N6M9UadayWRm+Vi1KrHeDKD0
LXlGm7TH/CLFaLPz2Szv1todMQAMKN7Nv9s4T4Hke29JD/hwcR5s6Ezm5dhg
iRYQn3e2zjhUj7Wz2ImNOggvj4nK/f6B/zjHLGJpSS9iw1KlrMlXvpIe5AEv
Wg0OyiVlWphZKGhxfgmiwDnbFc2RIKrEq1TSS+crdZ7fsf00lhnjRygrx4pE
maAQjA47IaR/M/84ruXLN4Ukrhaldf58LxOm1M2sknOKTBKjgW58sOZXaycE
G+IW0XMRd+WAggLpXchqFj9tfEO/f+9FTKUtv0lkejmlzGSnSYEduVMXKomM
kQzclc84+lPHXLg3yHB/sHg1RPQw/4D/7vKLM9c6yQy9QBXm+AlneDRxlFX/
GaEC4QLc1KQTP1Q8c/pCVPFDwEjD/UPOh0wJQvroGj9ql7aZa3vBukRuKOWX
gFvWpAvKSrA3IXq88K/YPMVjAHletqjSiSws7RGvcgssolTjLXsUPGSK36ub
QO3fuPBg5H2avlb8cqaBS/RtR18eul8p2ffmUnnrOSR2xVh/TvfFnZx6+uEv
OPO79BE+xV0bqOs1RFNZy7arDlYJ+TnXSFWvhiJhLEXy3LwSp/9ITHdPORvv
KRS0AKeB19IxkT+vcLC/nyehJbbzbsRtZpLvuXDTZt0hwGsr2sQQR2Npyypw
aDcaXlulQRcWF8G2C5VESk3dUSRwv4oJwHQZJrFNFzVw1rlW/GhuvVo7yuJf
0X9PhrU03YMEaoBNYUhXfdJyEpgV+PKNTt//DyGyOlZ51b6vD+1xlMlQ50ev
+9RxJANnxtpMzFf9Tjn+xQ6S+Nrzw4g5+RimdIRSZXNbA4IGVc+qg9Ccp+L4
9/yBifNEn68D3w1yMxPMqt93seCr1RO4uAXjyqADf9i55i0ypDsXuktgXsAO
dI43vc/GcReY20hhH1P7ue0nfSkFZDCtHTnubjtOCVTq5Jso/2IxdupgCf1Z
bvvaQj6xhJyZeGndtn8WNXLnCA1C+XTmKA9gzzEhdwpO3INefPbR7HkU7pbq
7CLf2LqnsCsfzAWD+Egot2vyApoTC+Sq+kczT7JslgDcDKxIJfHK1/F7ybdS
xdPIXKAbBhqqI5Sx9/O9qsOHuG8h8HZAmV/tcRFGVJE0pYxvXK5v0oDhADV4
mv8lpVGLpXUu+nXrlCVZrNinpMXL0QnNTVaRFStAAObB9bEpLqS88WucZTcl
GAbgg/R5pVgUo+VyJ1s+tCR7DsLXG2quMWxmFKCFjKQTmfWDuoHQ2M/9CkOY
UNE2D8acFdjInTeNH1QdEIONvicuYiEU/SQwaCfD5yplQk/o/z05NVsrnHjW
7nxdVpmLV64VoWRAwx4dNf0TLX3AwHRDh3MpP/x8m1VYmf7/+vyWQA2K/Rry
rkiJQs7U+nOQIOZSyKMbBECH3j/Sk1dsml8u4d10Dq/Yc1HzkuMpSHjjxhkT
AOyYGzxymVl2QJPzmsm+2fokC1HVlMiuP/XMi9ck0ic6PmcSrPnuJco6/u9l
vZnK920sABOPIEPgrSo5xgCd4Ej2RRif3IdgcvBtYee5G9h9fgUVouWPKEUT
Em+Yy/F3oAlAeTeP6ILNDiOPO2/Aw85Vafjlzei951PIc50kTXnSJM+bH6g3
q6VM92dauzWZ4BDDmJB40d74OzVaog/vtwk067bIy8E6mBtziAT/yebhPAND
1hLyFKeJ9lzg0j/0ImTpmQnihGuE0qpb4+Bd7ROX/TwU4P2CT5TkocgB0UbG
W7jFM7Cg4VExtoXpgMEx3R8QORob9uDS53WOE8hRVDuybLjAR8F90EcFkJ0V
wnfs2HAYzSmTPNH3hm7/DHTJZPhXSJZVJCGQYmdfpLH0exWYq+h9LtFg1dZF
Ug3KMCeZaSNaaQvu9wNWfjKOySbK6SZHez2lTLykcrysX2yKBryjncgVslNv
5FgWnH2wHVsuRvU4iTA8Ajkv277jloB+8nBhHeUJ8foGb6q9Vxfb1Uku2XlW
xE6cWT5cL8vdpwBeyi0ItAdgf7CZ0Q/Yz9vf6eaYVzKjCHdQjWEaTPB6XRxx
j2GRHPM+LyPlaEkUzguHrqQ6l0Z/h9OHZaqrJ63ToOzl5LKaY1wA4C04U0gn
bOc65CYjWH1Mc6v6t2JO5aqKsd/Z1ZSEFuS+mn3JpI6mWVPGj+6sktwzKsdA
xKqzEeBTJlJc4EkcGQGp1dJyPOlETWOuxxCj9vdS2ec4dEBylHc2jtwGUc3c
olq8dIYS1rZXiZjlesFgDEeXAY9SZg78FY2fiw+Oc5Q6Oyo/XjdVA2k1kIYL
ClpHSMzeVIQhVMz1YW+Rs861S2vtgiopjEx3uJHlm52C9SQJ2DOyNvb6TF3S
96mdpuRvIVfwvkrYnsMths+2yTKkOeB8IheYFIfTqSZtL0AjyFmKQoA+CJxd
9yLn8I811V9knQiVX2qxF3RCX9DuLePumm+GRL9Ny4VcqGrryJPen7H3AXA7
RBrjRZRKoLa2idJlrAbsPhfBLWJRw4Lpil+67d0FHB+6poVBh/qJrj1ufiyf
fqswJBAcwAwUvdY8KsmH+WSoPS+dpiac+mTM097tFi3TUNIy159pyRXJ0Mtm
EHc0euc/iZbyf8ym4zS64IZPgbJK/BR6sCCjfxWYtWEdQZTDcN71jMnXemU3
ZLev4YQT5i1K/UoXVsTerPV52CtBj7I4epELBRZqTPzpcZ2lRJ5vRSsYwslX
G6OU6LTQnBQrROFCly56woNUVpBXWo6N6OCpp2LYB5amBS0Fx8KBm9NL99YV
xMAx01uwKjo2snqqjKRbEFJU2I4z24rKg1E/SLuBjT5cYUj1d1qoe/nSrIx4
Bl90AfxrNVOtxZ2WvDM2+KQHTNAlYK4ntVeR+d0KnX3WrC0qwIy/pbHKL7HG
4hIS17Tc1d2SBZUjHaZ0/n0dorg6kOiAirp3tAEzIOpLCdEqqZDx3+N/jxLc
GU3q2WM+k6fpza3/7BdvKESZhkqsvZyUqFqNZBm3Ar8sATIoz2Jd2EzGgzf0
94o7MHltaaD0eowZEqQz+R5X9W71DtyLiVeV5cVbjkUnViOUk/KU/mNYqcyl
I2s7YRRTsbTEIXUtKbRHbsQCZix2OkQLWeSz1CKzYwAmIRwWXdouJ8EC6C2x
EI8rpCCXZvEaERG3oNYrjCdrZbXIjSwOxgP6oxG+r+Wzf6AaFrV5y5WYZCt1
+QLatCV7Sj+RAUlOxhtWziNxcCHHYO+kQ+w82D9K+wov7TIRJN7DG44miFzH
wz6kShLDNpu7vScdnIAKbamwWWiPyjiFXIoE9NDjnAyQEJ6PA8CA4LIrsJFs
lqh6m2DgSX382gW4aqjJA4acg2/ZwGKG3o6MhH7mbyUZtIAAgeJWEZnVAeJw
0mHNjhbFnOhFRC1+GN7Y57Y+g7NPnHLOEEkink7DgJ5HO2N8Db5KOxSMWbKf
rqadsNkUCyt8pYYvX9y0zatqZ+WdYNlBewyxLPWZP+FMhlOghJ4QLgMtqowV
W2+Fcz496y0ZxAfN4FPippKRYIuk+I/IJPD72z5PBEPBrAXsneJRebsgzMPn
cnrkYwWETRlKKdIRlkheZLMhwvn5Gr/d8hZQ1qTGbrpmkUxwKwVCqFrIl2du
JmaLtNu+2wk86kuv7lF38+qNz0rEh1tPaHec+QWBpOrIOiAuZAlU8DH8TVvG
jS+gLGGRC5V6BjvbNMKlckuqyuc9XoPEHXhN/fk7wamcQHv6E1Vj2762LudU
sUxValB1yuLVudCqCKFwEgqCLUt2jPSNooAwn1ETTQaeOMmYgH8V0f8CvlQV
JounTF3XWLr01/r8E3kDJBxf9V9s8edxU8KWBU8UOBdyDWxHht5CJGWuOWYU
iRt/6Oe+ZicKKp+OazWtylL+KJbgQOB17XDVTqe0h5LofUb4OMZUwWxj0AFX
j64KI88eTPzTXJwE/568dBwkTw4szn0wqyUpMllEMvrbmH62IAzuBQGvwIhS
4AGacT+nLbuY24E3cdX8TIM00C8xgGcqIMzhHJWiyyVWTyG3ETJWoo9RJFGB
MHjtiYgy46Vi4i0V3hysz1hI0yGQMOkFyyWj+EFTkm5Tem0ls+udhEmClEp7
kPb5Hwn/T3IlQfodqv9k6Joz9qp6mlJnJdIXuem89++imPHFG9rAgevCi6h7
MvNgKirbV5yKgY8Qn6U+x/x4qG7eXmB09QEzsH7ui5d/eXONZL5N3m0SbMPr
1lGKSCyx5XWEwCyjh0llkBIQifndtB3E4ADbPdPTsgeiCGsaLM/g/ugba+p9
vij4szmnV194GuK6/6voT2OtTd+e1ERUhkUMfMYDy5D/eJZFv5lczw8kZHvD
DN99in3I+ygqSX/W6tz8wvxO1UWYVu/DsVzz3vFwsf2ZFCqVsSFrWxXtTddd
fk5CtEgsmFxHgpYP0Jr4ZF/Mx/y2lie99qQK7hnuOe2XF8Xd6XE/NI/jUR6q
yli+mrNgKTMVEBjvsyQkB5i8Ri0V694SP5FWGVCW+Ss4lwPtKjy2ALsZU1aH
IQsnuGBwcAnu+eovVcFsRen4EfbxMpAen+46hp8tUSX4pv8LMd+CE+IzoOaK
OFUYHUksoBOTOyQwEufKsTNb4X/F9lpCRvLW0C3RPNT0cdPN6XcusnZnLS3Z
bkwhCXFd+BQoyFxkaj4SUVRp6cPdkVRSfhjiT8u2c8Ofofn1YB/zj9rQrtGm
kwG9JsXiIztFTLN46et1EitIORDmFaJpzuuv0WCVOZfVQ0hPgyZzEsWdKehD
aU9yqGsFNHVg1t19KZyXc2dnepKcnujiwB+L0W5scLRO3wMsggi78722tRqm
P9L48N95m7/8LX1cbs8MFE8oEl4hF/1KQ17bZHCJxgyv3GSYNVHkGS8h8o8G
m/EwIj3zkaRotDy7wOVO/YY987vjoke0tLYl7hI48B0AVH4j0mDn7CzmrMRI
RgWyD0qG5BoBJiVFi1UC+86PQBVT3M6YBPQRzCidrNePiqIGqmlVt2zX4ejE
PRpJQyda1gn3qyPOa+ZUj20S1hgVUTqVBhcjOv59wKg6nVUyzZO7UF5bsi3I
aq25yYOX+5ovNzcrbtj05LZpOM4G1F5LXbTY9/huRfgiPThCTT7HLwYcc4xP
b6saoaQ9AAhaQKhoQVT/uGE8PGVyu5jOCEHPnMBfzNWlb9vPRJ0wwKm7eo0+
5j5Mrr2i+ub97oRTB1fEkq6h7U9JaOJ5q2ZOVzhbDgbQAk0mKvgr507dTuuC
oFoBLwOzSY8wStaFOHC0OpQLDZ1NWIEA+cGSslah0vPUjxzRTCeJHku5tPQ9
w2Ec0Xxj7qW/ZZ8+lBFqilIaVeh11Vgz/0u75O07wbZUNMPvD7ZOIVqOOKhh
IwXKCBS/UKJnmL9hXGOKBVvfLW8ZE5JITDmaQ1Q8dcJh0WSOzJ4hzmu+D7a+
4UFneZH1+NNHgyIJQ2647w3kx+Tx8a5+2tDBJ9SnT0qkBr2hQyfMi0uk8mj1
5LtJmlaM1SZdYno2YUHmB57oiE4Hs0S/0/VFF7xqOzhsZLwke0AbOFBxs5zt
pRaP952obICcHeVu8DBuDM0uQp77pAv0Kf7ejwra6OeO1bOfnZUfg7HwokL+
sNkS7quUUXPIo/Y6YOxz01kWYGMkBo9sDitaRPseA8GPHLMrmKTO9HbPkuNC
5opGr26Gb1wZLEmUZtXea45PJlYTMMQSCSfCKcunQG/qODZSy3V6u0ZB8VUf
ykVTTS51RYM4fUrsXFtyEMZkTe4I57nJwgrPa+kGhm7a5UxzWCvq1pUJcBgx
X01l2F8hSYPWz+n6J03Y6w7aL3+4FLmOMkKHexuXw8TNUVAJKVzs80taJTHY
8Y7HB/fNvA2GatyzYofe9qaarwz6/Qb1bVAr0XMy5E90xbuUp3BoQBeY1d/a
WE1YFwl4WO3lSyUgt+zlH4kOH51PZkiAwU9DIdDwxq5wVQ92kC2tt4zG2W3U
y5x8T2OetGJhLffPeTqiBj2EbFe2eTwjMLenDsEuQfV/RqrYpFQrZHpyhSZM
iffCiwO/3WX5ax2aOrQf58MQT8OngHFXchPz+AQZraANKWQ4DHv85co3RaLZ
nIfaQdGZd5f/mG2rWL67B3BCtGSUv3HbOKQAFXfQbCu5vpaIM6Xyymw4KSXB
U+AN7sqGU6msV+IQbyfojd8NNC7+WokcZu5KJ6lHIMMjWfoZOhHd7xRabzBX
yp8yumasjVn0FXxl9Qyw7u6vc4Dr6PUbCLpTh7HtOfJh5r7ThSr0NeJJRkmT
cBIXgJ+H2RvGGlR/8b7xQf8f/AH8IMUuranPpo1yiLjFySRQESiaER54QFJV
wQtwuwzic4tgdIiYHNiaTHHK4sgi0Xkcq/qeUMMcy6chyaHq2+2EfqwVwbkN
3cLa9A1s2Jzx40oy4b6X33nlxGk/D+EYCupX6KEnjHIfa14rcV1v1xXsjsH7
cX+VhYxLznjtfivCICLq9KWpT5P1gwFiYqpcAhjv+1O0N13b4d6o4G4OheU6
cpi2c0MqvpNPHe5d/qtI5JLFhomNLZaWmN6VVOkYTcuFGz7571cZyFOVU2HH
5S1HflL08RwYwE/9ZZqLR16cKYvcqoSItXLpGtEGjvzj6N8twtvoWdWqm/qI
+oX8wscohGhWFzZKh7qaX9kU/gXPZt5MUtA8XWBXk85KtikTbXwHVVKQB1Jd
21UZMPdX5jPVd6HB1DcI8wfayboDU1uW8vB+gCH1BQk6fxJeLV8k5CBu+3mx
jFSnTlHgoCqo9x54yiDxdjA6v5od+T5cAGuFulTCGrNsj7uHer2ciu95mQKm
T+nbLOK0jTfPf1aElMdfSznF/m4KJPoZ+dGKtiINESDhg/XayrvcIc2BwaWd
vPBEn0EYH/0vfnf0gHB1u7pwwU9PIIhkoXjwYEhc86xekTFw+Cgl5EaoMkaN
pZf8zyu+QQsUgXXut5ppE1gRw42wKovvCsh0OQRuBo8QHiqr2YNQSqkevppV
07jeGEg5I8SFJEnHIM7mFAV375PEdd1PAo7tW+yNDB2/0ILqNI47Y1ONmBp5
1zI6w7D08FXjkZNw4+gsDVxFgBdpY+dcTiavHjW0mnePUbR5xzv/n8eeDnpI
vrZMnlI3BWqQYQi5AWY3h7sF8HkY4uJV4o10bRVDhFRnRe1GaCeGT8AN4s5E
5C2pdNJif6WkonT0XWGqQhh8nWVdnBJ3J1HUDV7Y1Q8GKnjkufdWX/9PAE9V
0x1E8i7PUc/3I4kXCCXcVC49CngQf7rgk40gOR+3St+9vHANmpnS/CwbHM1p
CkWPwMzd6Nnbr6eqKD4g+53k7FwigiXmUPKzpoAG2clsj+H94GzhzlQVoI5W
0c4253Tmaq1msut6n5WnNkKWI/Py1TxoaSq94IFEoDCcp9SjztsqtuQZ1iFf
4iJq3eySYUNclwQGiLqVDMqP66eBlA6g+Ya8QHTBOlSuX8ZpJFdTIvwLU2uR
Aiijlr4EC4FG6mXcYTIeEOaqoAOG05EdXnhB/8rRvo+o7/0Zsd6Bz6+W7UbC
3AFwH//NMRl+jio2vCJvY8HkNBJsCgEh4iC3v8urYdKfXjaQFJxvWptX8eZu
4wsyrI8f7i2ujvdHN7JdVdIaEmwS+VpeQtSbtRJM75kqcWNYPUXj+xxX/vus
JIIzNBz6TMM0rJ/5D4CxIqYyIMatUq1flZ6Pmc2hMWWJ43/k7KVH0jXNsMZm
oRjvLWFOYtFWcVo3JvIDFQRIeRgiGfKhNZZCnKso2rkqaekkPsZIb8L/HSV4
rGYdJSNCHEoCR+VTlP7N08hruny1v2jMc/y3NjuQ7k49PNgtLNO66zCWDoW0
wlvFdw/X1/IkclTsvJ8C+EyfdUtMSg19b9ibuawagzBH5xbmBg94FuC05WFu
FFM+lhaz8kJG/1UpbihRKrTElqSbfztys6mGu3/uFAvEEPyK+ZcD669DYp/0
yx5fT9NxA0/68hyuDoYN+At2Z/i3wxbofDHNXTMdLU8lBce//tonlXH/Nc5+
GQ4JPVH7gxeQGkf1tJtPtTkAub3JfGIJubT2AWJ4VJ62mYhYXsNaiMjSlxzp
5cVCf5TEd4uDGNFX3ru0FWirEbVvvdJeXuQbeX/gGy79SPFpGHMJxU/iNnkx
XtqSRNEAiqbaw15eFakovuMrgpnVFyI5aua/rF3pb+0ul7GKMHt1u44gEvMj
UFWY1VSZU+BSUKsvk7NedcNhjF8ENKcfqhLUMG06A70uiPRpguDEuUgeNKGj
AxIXfnpH+9X2vqYiEAIKo7vjaRoSHTOepxyuzm37SgjKS6ZWwpsFbHvxw4xj
hbAmlIW0ww62wXfQG0gAl1uLs3G/j/VT9RGCLqAp1Ly72woeD3YRsu6Qb57K
htPjLNPKZjE8IgKauTaLQOBC4/bvkSd9L6tEeH2l4q49WruLh7tngEJfm0ji
T5z3nb1XEyJKktilQlnwwQHjKKF0sk6sqKl/S+B+b1VkIr5nAP54tH9begkn
h+jArHmJN/y/SvPgSbGXemY5yCWNt/wJyENPbfsvENUonENtz3GnO3dv8rly
b4EcnqDFkXYb4cpqXKnhsLlAVhlfSU8z6BAlLfOEiO72pe+aKd2xG2jTtoaE
Z5ius+OOk471FE2ktdVSOCu8iNJTH+rRm2OCdSPWDJHEf3goJndUJw5mS0zt
UpOGAaCGQzRa4+paajGPZc+25dXQmDNafBsK2bJQDH8kSrSA1vybkO7V96YO
j0vV/C/HBsNOx1SFTPsANVRfQJf+777vs9U+OTG1MC4b3Png2aXMgWuwQIcV
sZpukvWkVCuHsZW5Wzct1poiihQFmuW+1gHwLyqP3qHe+c52SucrA1DdqUna
2ntboyJdZT9I18QHk0fwbsB8zTMKah6zZ4E/3ODZcSKgOBmk9YJfonnXgYBB
SGvMh49d3G3UjvAtTf2oqCs04nKmAGi75/j/aNbHcPpZQw3J2SVFC2h25RwV
OhLWzfxSu/gi6snzhrosN2nk00BZvOa4AOmLK/uYCOjuAV6yfEHYVia6o3+L
ozoaEMMtdM/GZ9XKg6BJZK1RNEj2mak/LaTGKNTOV43yUuS5L1h+rRIdyLOR
Ez4pM0ufeg/Qx9VtPE7AnvPehx6Dpq4D/vcdHt8Nin9Fo9pQzCMf9OkEoXaC
LSGzMHyK5nfL4kqPwJPvs1gfxe8wHGr63YVXyGyPefS7bapOxl8JONqbDUxi
j0HkILBBppW7DpvMtZZn58RyunJIcseLtQihvEsUqJ4rFmakTCLA1WfOcJof
Jc2xMYmNhVQRi6jR6HkWOv2f1zR9WcxCZmQPmuBWD9VIqJuXzr+xI1PqLS6m
kfy4WZhhI2dBYHQt/aqrqTFBFuOdidaSf1hZjUovIi7fXYyBIeO3U2dsUdA8
sE+zqfDd2babkzHZA/KGTIcG1GU4bY8FjAWUHX+pNTYG9ZX4P3/lG9vSJyU4
imNeOhIEaSaE9m4toBajYkv3/a0nxOnU/eN8aWCqXzaeNXEN1BMwHXRjHS6i
FBDdrSbj4peaJ1raRUZtMScGgJ7NTYVMNQ12FCEd6I1j74o6DPCQ1zPwEP9f
UhTTaT1U9SYNyWSQfBo5V8aLx0tuzJNIA0Y95vY3whdi3AkH7FBfS5RDv1ZX
spXj74Hnj/ZYEAZT4x75pDtgQ43OQB8RwV6nyb5t2bUjltVCUIacx5prfDz0
8PeXcMUBg4fJ/Pb2kD3o1an7OiqKNbmGmSGMqxzhiwIUSTTqloPe13qLrDwL
++gDTxHhTkfUOqv2Fohtd1TfDf+9rTqw1Gp/MKnUUFLpWek/N5SxVVfVIuNi
STkeHw2tR/c7xnBnVaOKNysl2dA6+EU0e2xs9NzkazU9FSsJglKIq+HN+flQ
so42v54nQ5fM/hoiB7xEgSsWnXbAmqP9FDpSN9T72nMzIx0/k3C68Fu8MyLU
WiUvbg7zawM+oncWPwdSp4CZOpRO7/1XrbGQ+NVUcSJAHj3Hs0FcxHMaIYJa
63ZXqyYfrcgraTidXH8g7QlX4hc9p0R89h2WoKMKcgIo5vMPEz9b7c/0aJam
2fyw0wLgASm5CC8WbBn0dG2tfQnkaPUbmJmaF3mdCajRITvVVGK+ClxdZfIe
N0Gur4mjZuhCw5TvUdId9XbtuU9nAYl9aKURFVBApVUxuxJc/YxlxCtELyNS
OLS53Hnxicl0nIbh9utPMhkA9f2GRGmNAmV8DEd846C2SvgtwMmUbF/pM7vu
qEplNGdOdPXC0D4T8EHjuEVfUD0VT1O3ZtZJA7J/ubbPC1tFg4jfMeAI3K8L
T0eeYuVXESM8Gkb/TdWDtMX4JkcRGBqGlUxL+UKhf1qJXSEmeDLMHuAqWl2K
MkAT2SuAq0gI6ZE9plaPdBbnrpCiAkOjyH1+yID1Kg69u1V9TTiKLzQxfJoD
iS0zCZUfTb3tZ3Eq8MbwMTDOd24u7YQ0mvsd3k+wg6a2dx7POXG5sFy1cyve
mu4mm9OtlR2WhNGhvGzpdkeajsulQvpdDdK2o0nzj9KmZKntlZZdKCDY6IWo
ZDwYfi6vH1CirvXyEgR1gMAMG+aZ5N1BhlS7AL0uDeeUe+yj7i0rIWEZDLDD
L2//4+XIcPCVYcxgI+cs4UcQB8b+9sHfOfruNZnnyKpgU6Jang75AlGl96Sl
BgF6QolNLNxTqkrIiqNp2BMhADYcjhG8UzkfVPEXNLCNTYVyrSPvFHkaSt9E
TWmt4JKkWecG7jhLadEg/lWkmPNxcu1xqkVenyTzSInjQPJXGhtjPWYhLVQF
7Ztgt+XW0C2BK1zPiKwxZWG7NydmQ+qkMt+ff4TcwIbTM5+q4BBqTDBNhJwk
anoW9Cs4FCukIpOr0E+LB7L8zkD3HvtRnb4wODWZUTvJxsLOVzp7lMwc+isZ
D/sKo5yOWL+wolIii5rAZZSEhslFY0L10kz1TZ+s8rwoDJU/tyQtuUz4ALgF
h59/A1l+p1bbiDSVYC05slTFaVG6EFkVqkKFVl2BSMtqwCNW5ifgLXgDcU1J
y+Ux+o0AzOHZBs9ilzvGxK2DYxY3LgK3OfQRq7FXCbwhDRLiYpK9ZFHovMno
44QX2p9tDxfp+rzDv2nhfQnP7UgOf4M6VgYipukY3rxy5KA7dfhk7HGEBY2t
77WkwEuG5ygY0cxEjv9KA4zgrE+lZWj6GQZS571+bFmIdHDcidzOkgnf/svQ
X4isl1BabV7mSydKaESkzTMVSkj1cIwZ+NzH2i1eNVAHF0AEZzypMtKanCyn
oPGQ/AYzeuIUMJTIzYO1K/+o9Hw5SpmlWQS5V72CA9Jxo/THcRQMgn21KJ3M
Wpp7Iox6uv06O9KaBrqNoYCnuVHFhD3QcKm+qiHTxfrlu5KzpjZDRQJYa33A
vRuxsriBBk0sJWO3kNKaG27eGbzLS7za9CTzgjN0INHATg8wwJ4o/30X7KIf
xXvktaOUe9vpOD+aTYDgoYN3/duXzu3mXtukCALX88hWbAyoKAUqghlcAFbJ
Pmzfqe4qzXOWlHCZpBw7H1TOQ/CH8q24Fw4lp02qDxW7jMZ+NWXjHg5I+xFm
dyKxLazEEm5HDnNrAPa27nIDHEX51OYxCUut8aRoQoFgHj3Uh9/YMcRACc49
NavnZDzphuq/10qoNwPVfNwtuGMXRVCMZWNb5xqso+5wY6VizQAAzHeqDGGd
GV/myGJByL+z8ey7BxjWu0vXitvBzxUo5RJXNmfJ/dJLZw7cT8MgKT6MKuie
FQEAdARZyQjp/MREmKcYWZcBB29KkEaNTperKCzwitdQX193aK21YENUWDrx
+1QPxzbkV/ReLWQV836i7ucSkVDRcE2of960hYq/bDEnIXG1Ie17jG7KQvjK
R746qiyA7m1aa3Ae6+DgEOU1DR6iUT1oFfZR9Z/qw0U29kgs9pmlT9+dsbOJ
Xga2JE2bTw6yp92WhVhQxwdUT9bG+RjPKCI5eIX5amPwPLrHyoNnlHonclDk
f5ivDVmCLYaA5AbfJm3IMQXer6CU76kWRhZO5SLjJ/aRERRd19QBgFN74NYV
Mv+YgSsINrPpnV7kT01WSALQawGWBAcVBEHq/lIMxgZd3UFkm09aHA5EMGeK
AJ4Tj2P7evwa0SE+iPaOmRnGTF82HG1+QW6wZkUdHLotx5uKi2eiI8zDWL24
Ei4yr4tvdibEXYTg7Oq0Pc7g6bzvjL/uBkjDfsveCSOpWak5desFgjTfR9Se
Id6vUIUU+1jI6Y+2c0uwkMxVmGpwt1X5ZuWrxtr5mAWOJiRogzHL7Q5MIlfD
RaEt32l6xT++G2Ong6/mVBy4J/rDd7h9m+2DCVAnNWErgF5WbxhQ/jv/jhzz
RhQZjq+XuHlUs9oCloMJaugMr1t7NT6WXFCHumoGngEvvvk1UTrdcn6QJ+5c
6paa9urvfHah3gsjnYxEXwEemHDFOIEEFiIt8NQdpCwcHEoWasyrfM0QZmHF
R4tURI+AnqvET6zuh6yGlnfIdpyyqEkKaGviZ7PF/Kty1K9j4HChvH+juQGP
Vftax9K3NimuZye4GPHMs1+cPrvmDu1YLhKhTSuK3e427zKBbgNf1MGDH/oE
OmRpapnEH9x3+HpSuhRhLkLKIu1vV9RI6FmEbUOS0yNN6BoA6gOyJxm+LyYJ
9gkm8S7lVcCe3hWu7Ag0ELc7ETsNjUOnbbI6+CjIr7704qJCU7XEOCvwW/5r
/OPugDlXBnGfVTjQCBONie3/VThoNzgtVRfHpdwyANPXleDJBDq52QRdYeyx
8btcFNwjoS2RBBqniwmQN1QVxrseCba1uGH/MYHqITbVX7NmopYcz7/AYOkr
GybninrvdC3xiTR7IC0btNUwIwcI/90r6NcvI+ihzm06K0iyiw/4+XzFP7yH
Va1LHnl0Po6H3OMQIYRPbP8dgYAjf9IWmHCCtgIcE/CCgSSfKWNZy5rfc4tp
DANUShALdl+ZMYg6cxuVXG5TeWohnuqTNr08cpHbgk2/CdQH6wcZal4PNDnn
H/whnFj2zvyVjKYe08LHkTh3ckhJYEzuwFcUFRxKvAn41pP9jMQQaccAbvdX
D4Ld7Od23OPyVgEO+W/u/98lQ9GnAgCi+r3XyAUn2K2fzOYBHFSRM0aDbFGK
03tUTUQAkOisKvu9B94fgHQKpqWX2fUhYxMhiLeTvD3FRaxe+fHkZN7m1loV
wyiGRRaemkq1nQ8gd3X/3EzoPiGSShSjtHvdxg5hVeB9ufXPbinTuQCAn2ex
fXuYuRc+Uuc58h7/hW2ZCPfgEYaszpvS1at4Q0BrTYx7ssvVi9dFT2CclzyF
ROfMI2DXwgaxdg28f16ink3gWTnIT6O0WrV1NfxvBvcxJ2H8HSaC33B/AsZO
X4NTLxQM/N5LzqI/uehcKN8WZcqZSu0mvtVhUlQujTS7RhZwEYO3DdKmg14C
HDxh8/3k+qX95Qhkkq4swtABOA1TpmIeIxXnHwRysE5Tf0mhv0D2HDTEQ5zB
15/tuHJFdvSnZrdAc53pszMGup0rALp5t7n+txeDxn+22VYGJsKI3Sn/33a1
tfa9siO9sze9EIO4bLwDARpy/jF05p6aKQCxHEtPRmzwy/Lt4peWCh/2WX+/
NHI52Tq7T2MjkBFvdLzv6lKajqLot8NcZTXVpcxRkbzX4OQPrlZEhDBeXSsO
IIwxxwPHqtCkZTnMuqNdWqJZbLVbxKUnPhNT0HMItjj/6Oa9n16vZf2WEhIe
yXxo7vXjzOZvLj34yW8vWhgcRE797+0C4tBK5BpuhuHJr0dTcr0GG0wgU+mz
rvq89sOSOIk0RL0yvEes3XRdp1Mqm54UU3s85af/aSy8VX2DnuT2XP+fEZgY
m6QD2Sj3zLw2uXpzTFhz6UhFxuNlr1hDstLE+F7IAqZiQ1m1iPVD0Itepq4Y
xTm+slqSYdQS1JQscbJMxNuNYcA8PWc/kEOCTJbXHMfAvMS+/RhGhQQbdgb4
urJ8jdqPoAuTtRk4GtTCaEijRrCJfre4FHCU/G+pDEdL6/OOXQ0OMwFVVSDG
IRi9SupDcNUARCHEIr+uQFaonwogETxfZFXB5aSyoBffLHqkxmAOIKYoiL/p
tkqVOGwvu1264GruxoyCZj600m22F+Gd1kiA8kNglXDoMZC6Q+X/3PGgnzWQ
R9x6IsxXq+tppKZcXbucTA5tRLu7myGNSWjvLDsssauYAnZT5p6zJe54BR7d
evpn8P0Yi21kCNywc4BhOnjsUQltkG5wHhtBQ8cfcNIdmZHiVi0dm8FTTBOT
k2mmsHd+vZC3fAjHXXIL1hDvjFq3AsV6W1HEs9wJ7cWX7dMeSwOfAtiwwR4k
t0xS/EnG/oQ/E6Wm6OxJrhhcIVWmu7T8IKyaDC3eBxwTBO+0421WOYDgT36x
BQCtBvzGTU5YviRuEZ5G3FhZNSVy+QpjnnNI/kmA7tpqVuOi5Wea9xTW344A
IBR9JYwm2k0qJuedLMyc7DpbiJ638hVuh+J3l6PmYqBO9uhrDBl+swx8kW4A
NPYuKQtanTEKdUuPtq62vpn5VRv7e5QPL1Mz03gIGJi/T+kqEnVmYf46VuDm
X6CeXM/loxqeWSf7KcA8ONh6HbZcDSg3EW/IsdShIm1BcXWvErMYoxnmfKfN
VbAWBsw2iuLmEvbbXEhIuWOW/4GQbLPzRBPAA6On7efeSioQ+WrpPfaIqmm8
4uuEdeLnX6rI0Nw7oz0fkdvXFtL7EIrRUJsEmuvvd/qRuMi5CSPVbR4sdBh0
SfCdg+AVMMZ+wyi4MOjRurz6cnQkS6X3Q71Wlm4mCUbA/hIIFGB/Ie1cBDdD
qyqhlaqLZzmJPA3HCcfz9onHkGEA8/6RyjSK3H4VzruJIuqsx1HUtvPv5MQU
EwGuaMW2HjyrBXC6Fxx1dSAhydcRsE6usrXoMp+ddxOb5qyIGEpVcvSe1o1F
FnSdEosnPXw7+fZyp377jQlDwu9Yc1iYhUp77Pf8mD77ziB6SAFg0NbRS1XI
5zB2oXWhjmvaJKFSVHM+8fQNrSeZpob5sweO/QZe29KMqMZbr8SHiNwWwuqv
KBtEuajqMQwIeIUsU8x4HgSsymZDOvLDP4NCGDiIFaMPCY82j0a876EeQ7+0
V3aOXRh6ZKXuavfJbB1MZ42QsFlaHSPcRAPWotjbFRWER5gNJLTvRuocmTtJ
Vi7qM33zucYQJ/TOCz37PhwjNcL4wML48oP5o+qrOy6xulShjMWB6Szl/dGT
9dZ5+qNjbTT01eo/kjsvgYjs+jqOWTGD4+4qNOTaHeujri5eqOWrlct/9Zhp
DTfu6hiQS4yBliIA9IjzjftX3G9bAOu6KXLKr6DJ1oVerRjn3z6TX7N4JhbV
pleAKMgmTmSRY/bqgcTj6Ng8hdaJEu+dutyWvl8tFgEuI4u3BmjwAbaULRE7
CsKENihAlb1HdA/QSyuRb/5Mh/RpBhI4ScQHsV044sJZcIeHi8rU7DwdgYJJ
0prTsr8lUreb0mMh7iguKPCIjiRoOR5Xo+xYxvbBdSjF0l3pY6jQXA/X+L68
pxHqWVWlDaWUpnGsgkcPBnCE8Gh9JwcsoRZ5uiXgr2Ckxwn2x5qptAXkMAAY
rVfJPtA6vs0rttWpFH5apygmTx2npLk3hvxtMUa0C4qo/7tyjHxIAKy+9ro0
PogrUBXPQ471yKwH6Z5BWro/9NgXNfAKnTK0VilCoTv8FYxSb8ASxOoEbGFI
+khDhEhiFlMnC/lzRHHONCb5zNvGZ5uTk8nefruJmH/SuUHIUKyEeBlLfoJF
wMXTfgQFTqjd+lTDIHuYgR1KCUStaPopsbTfHeCAjPjzlRdBFQoIG8GHS8rN
sxf7/0VtvhvBHAc2mpuhDb8to+i8BJVJdf8+S8yD3iMCGWFmmvTWuZk6EeYY
TnlWYF2fLKDxzD3HTBujd1A7LsJE+nFxUi2rAvYDDw/gDvqp2Axicj8nn3Ou
RD5Wgbwe6cG2qTdQMqP1V1JdDRPRM0samkEW4pCz/Gw+KTBalcf3xDlO7sjo
FLalwGkLdFi7juYfD2q58pisiMRzTRJxilQ3UBJH4+oIRWgMDh4avyhiV9ZK
ViSaL6VTK/LsfPhFJLF8PRtsq4PeHCfRtlnShVt3WAs8eQqOj8dmBBCNCZxT
X+3vhg3qTvUlhW/dctnyHR3NS1ZFsrVGcw+QBKo6OQBZ89zr5xjINUM3OJg1
SKIU+0lx2c9oHQ99Lp+gimTGDwNxJog1zh1iZymb24hhDfToJ2FO7KShdE0N
nqg+DmK2BvDiLH92aVxm6qx6idWy83PtGxA4mNf89Kdi0+dzjzI/fIwY9o4I
rkvbE+S+S6AKg1e7i8Jwktm9/3FALDUbO06UMj95LKlKadctQZOL9StQ7cdD
9UlsbmErcXhfIeMUEb/82bzVbTu+vcYTpu/oTGvW/hNar+ZnavgszTnsYUJI
xKpKkHf5N4FFXcpvNITMHgBbcW/8M5U0Su3ew1J5sJvbOARczcHQJc3RJl7G
rf8f7isbc6k6IfBgGeP9+KjlJycHj1BRW2fbffqwDTiEQYJbgBgZAX/G8o99
i/kHJLkch+lxLy55Y90P3XfFmmTeL0B2lzPVI1BBIIuSyazmSLjRe9ZToo+s
TQNtdKZ3KVYPW1QpgNPFpFk0R9gcL9nsjxsn3ZjUVJVtueIxFS+NhRJiBgKt
srsJVm5HGJWHnezKtRE/t8SBNzy4CYS52XxaFTAlMm+fkgY3bvfKHhpkbaVu
TaKDSc55BXWteCH2/2hVAiaYl8BYPEngb/IThtYr5s4Dq/YXyQcGNY4I0ZIs
hla5bPm4Jp6+5YzTbtJHPDHM+uSl+YRvltqDQLcmKV+Cwip7EYbNwyQAljLp
irj3PnfKX3722uEM7CMmtYw2WMi9DSuhuwT47WlEfY0y4Hlvw4+8AOgp6TzO
vVIor0igKN1c9iJnHayxZgVB5Xi9DDD3BMTnrcT67uJsjfeWIf96aMvmznRO
h8Mf7stxHgmIWxK/n58YfQh/aNUPRNsE33JBLZlhJ3o/vF518Rc5YMBn5n0T
pctBBK2TtKENIU0azF+RPhCdlMEZKD3JbikTe/AD+pAoSae6pcRKdrnHE6RT
TDgRGrNO2Zwb/tCL0ywTIHdyxGPCEuV4POv9jVI7+lENR9oaz8x6gqVsRWh5
lV3Xx7/Jolb6De7mRaML5uvJgzENIhQcoE60u4CLjPiah/wm5iTh6fNSxkZW
8L/LBi5AFdxXssKkSo34NajcIV8swh9ks9rD5YS3xmDxx3QZkyTseOQFfC9W
4cibPLrFaAEpCujmSs7xZSy031SnpQQFZoiVisfD8Sr8N2l+EPigCc5fLtaa
v1LIqMaG4LaO/vbUYzzlUAs+QI0JNJPzmeQwh2m5GEvVQTjkKjXH9Tyj5y7f
kAMV9U1alBpLMu3rHKv6F5ZaEWt75HEN+Y6a4Dnjpf7QxscAJizreXhE25Hm
NwWT1UH9BawgggcLAejJJcTFlP4bhhHZFPPIqFe9+Uv13ivBE9uXGkjDGPuq
UnE72tyo/juVLXntdgaIzTQDyeqnhnaVXoYJwQcV6vms3RuSnkLbpvTMw7aU
8MQO/SVwGBYOnbTga4EzF6DtBxMkCOlZJXf3muUVwV8nb0+9Hh2hbG2Pvib6
+SXH22jxYo3/Igdz8UN8MpX2fOD4Ff6NgPi21QMn7Ye6vDM20FtuhacHMJeV
V28wvIADra+/nCMkS0kH4CUB0nP1s+X/jXb5lXNKQaNW+EHbh1yw45HIXgH7
Jb1MdfhdHvTlTNrTVavdSvtrdMJAoDsGt6JL68NBoFXMOZcg0x1YETCM8tTL
rS6/MlwqW+ExdFphhs75ec5f0mAUiWwED6IKv3PiLm1DK5BsonQWOmGM7p3L
Qbk4rnfur/HfltZiTj0NczYtmqcRbhDQ15oirpwE55+AKrIcDeg73HX1sGwj
rZsbzsWK74vvbDy0ob3q1uPqF+yiNIjldzN/Q0K6fuGzgmOWz6zW5B/+gG1L
Cn4B3sTKYlUhm3suRczutNKjiqcrvd6zvbU5FsJae6vnl14r82mkMrFOcz6b
hKZCf9e4ZYpNsNHPg1BgLM+Ne6cgi0wC2IkPFgCp7U1KSQcaUKI/RcqLKQC3
PAxthyjTRpNNmESR6/6voag+G2Zm9WjSJZ0NxG+cpobRpnaHMYklTfe8s26z
OBm0SV74BeRa0LuI0JHNw/iYeu/WrqArJPMS4+y9Bfoe0Uwc5TiHKs3nDEoP
NlOH/dMcXVxN303j18Grj8jFVjVJTZvBnA1eDI9p/JflMOlv2dOP7hV/n/ts
IeuN9GQZuOKc0cNSibd9q2xfK0YbSdhBQ2XryduG8lDgbwPX8kn9fibLDv34
M8gbkSZ5CNwNwKZ1fQI8U4SfYcXrb+ahNGpQtBHfojzSkOaPLs+LLf3uvAue
UyAdgmUhC+VqQq1JiMGisQV6OV58Q84eZNELOJItBCNgBHLpZGWcCTSBI/Yc
+lHoo2QRLPB2aE4BJrUTYVWzXBVBM5+hviGG5+7bObK0WDe7gQBZWlKGcVSs
9pdvnJ+mhZ2v87gwSYVTx4XPzFddp9SkNefNmwOOtHauHmSfL3vaNBl2dXQo
/NSfsEYZk58dqEvZMBNY2dhRgbxxyWQutlTJ2+yTna+9ylFb/phTSYXpzraL
RB/YV3KIVp3tipIanCmrO5k0CDLxt8voSGqJN6imod+cBeADZH00dQzBjua0
rWqBBcXdGtc05pPhwak9NKa38dqOSJYor7srMxtJV/R85fAt5RekoqkOPzUo
aqEW68A+R+PnrsCpI54JEb7gP6jB0K2pOQlvV64C4l6HyOZBVlZWO7GAl1MW
28WvG36qVPOTmoq2bkogL93QADzsFptaFJAdwxGNeqLklTVv3x+ReIl1KU0D
TNzjPmajLkomXFmTTHSXQoCcwB3ZMZrBuLdfR/LVN8mCwQ7Ce9eRrjjPrYhY
RKUwWTkVmZy+k7Y4tyVLQ0wrFut/LCcISI+wMpO8hn0JbaJTjfJKigbEwtjM
H382JdbO23kW0xw4xtjdtWWLCiWx7SSn65/bJg/fSIF1ZtGmmlqaGpPwfbHB
tWSwUQ2kRrgpqCLcfjJHQk1ukCzREQhXoNyVetkfnzZ1AM2sJSPEUMoDbvFL
Bg6PnThKZSbL2LUxeNP9jBGJ0myYrISDw09kie0a9YvpfsqoJDfLSJDl8KcZ
QjgGSaVSZhyEF5kHyoce3H16JURXOK4me4+AqXk+tCQOTl2mstCwPBMv+J1l
6/N2a+RpfruMZ6+R+8c6OLPhDl2M1/MiUMO2Boof0rb75q4AS5Y3GeVc95Nk
ilu1eK59npUFsBurmMciLbuGDIWaUu2sIW2YSYjmWt15XDtdsTPHC3A3k3wO
SJhzpsjFKjVS6u6/bMAQSAsytDR2FDrhlcn1UCjc8n437k0j12BQOjVQiDzz
7Jg8TUzoENGJvEvKlz/zTBvcQ++p2DcsYsp7pVHCmEElvTC3SejA2J0oTd3/
8HjbZj6lNltohze7s6ctE0ehDfXc6JwsDpvzpQB2GuY0NhUKvmMWOeP1Ikq5
5s9QblLs7vYrGbaKXSOa/0Il0JSQGmOqdEw1BXyGdHRgwmiFMfFiaF1gcQON
3ebjGO7XoP+BGdcwVnGJiQWNw3DSA8IP/9N6H7yILK+QSBGdETzNHE4jwKNW
t0NIM77VwDs1b35KaYTT/Hn772z+UN5DBRI6aFcLbPIdYqUN+swzzYPxcYfz
UmUzk79RMfzAyLH9k5J0KgoUWIan4S4xXyTSi8PhqSK2Bl0A81Nf40WqSSJp
nghO1T7Fs8l1292PNrejEIkxD6+COiD8FbXcPrhYxawlGNa4Q3WtdhZP+jMl
YxK8W9tJrv+vgtV1nIjPg/azHxfzkRJw1WlNh9TpqLcbe0bcktXPGaDLqKen
3fKuXjf8jgSFVYuxGqB4tamufYw9+KUPq6ikIOhkv0TFg0Fv64GanFnZMkFK
lKIEFon12rXFhYCIz6J4fcdKLZB/SGUd2iNr/qnoPC3jz/Kv1CQ4vA2fAU6W
/TvSL/fpYte2cSzn057jUChh9u7UZylRxIMJEd1QAVFn0jsMW9ygL9ybQ62B
xusq6CfM3W9VKhZfKb1rlNdYP15S5dCpBhRF5Q+cebB+eQXcLTPHGPiPAp2a
s5uEvMpzpV9zbJeR1tasmb4BtYdJFmWuscB9JsG3V1nlgWcqy0qG6R0er4LR
xDjvZAMzYwNnd8tO/HD6yOTgC+ephV0xyhIJpK67Vg11z10+PRFEVYdiKtXg
Cmo9Ps1jMHy9OupvMYiTZ+P4jlz83/oj7wr9lseBYtuhOyxbiXmAc9NTSPLq
e+AS8fUD6YQ5PQVuhYhqg/xrjuAyGicss3n6N0l1pEuVeSQfZOARyNiKxcwa
lgqK5P6Zac/NDrfreLjRXBoDLA2kjTPOQmkShekxMFGJO3o0Pe+DlF5ftbiX
eWRykydkqU177r+7xnAHVN7ItQ1+e21slqOYqxBAfeoWb+xiDud5cAnk5Oxk
Yo1YHVhxHKWr/e9LcG8b70Mb2bwwtxiEV7kbdxQWi/Z5D8Wlg+eXo6A3tbkM
VaBlsXd6CU9fnS3gbB3FUGOrELmjGp2fRaUlWi6SIPjgjW9eqauHn/PyoOyi
uUvPCcDxI22M5y6WE52MKsZlW2Se9ZG3Havdt8T+P3z6CsydXQTRjonJinXv
/KtLMVcBa6AEx8HG4Xe5eH8DpxK3GewxKvr7kvIPxl1K2qKZkQKEXyLof5PL
VkHEu6JedaGY2FAA7kC73cBy4hEEkaRwpK6j+YQnpXM3Jrppy0rm+vwb/bQz
8vtjdpzoD6UoSwfost85L11GOk0MnQ2TV+yUyHLqheBGZpiMuSuxsLUIrXCD
0/sGqkb6JedXV/H79udqgkH5Fc1HyZda3WzdU/blQKFutuTbndQ1ux6ZbYGk
VY0GPMad2xY1HTQ3NVC2p8XxYiYJ3kQC5sEwG72m/oJhq4gyLnfsZEfoXZ4x
u5AblWplNdNN0tPteiuhNnI+LkBET7M+GpTJb7vVC5FtgBtCspFMrRQmaX14
jQZdz/xlZdFsfrjX84bB8ZjLDiDjouGL7oZVhjv5jA7NLGPLBvNJSt6h3NjS
Qkl5PmgtyuvnItS3MmFC0kHWbH4MwqNpDsHjcaDpsvuw1ZCe2qxBzAT3ZToo
6x7xzeyegfExzgdnIp82gHHp6rG+nD5R43GkR6C+Kp/RrEm12mVgPdwIo/GE
mZl0qEmW8H6XZCUqKNfWkcZg+eD6l75W1U9dmwiUJq5hQMh/XhGL9EEERgLe
mcg1P+UbPOMJeJZobGIUvjHeNak8k3itfskEzJ+KttpgDzpltXM6jdAmGchZ
RtEkb6srlUoQlBoCJx89/fwrYQNzZAsj8odAVmz2Jn5Ukm6mM63AHlg+8Lk7
Vc4VLTZvoluBKSkzXp/trog+9AuKkPzuCvbpdFTPbDY2ymBKuThLsncKJeay
LB1N8bGsI4a1jlKCncHU3WBjP8hqkTyBtD8Z0Sx0uRenlSYWws8VR8pzTsX0
LAw7VKROSRYErpigfuQXFKXtSixdQl6+X3RSyc1/JIginyTz3x3m07E5+3Mt
grNNvN5e15Hd1sN3UBn06Kg/z7lAu1rdjp6CtBxc2bEpQoPRHL+XT/9TXeQM
E9fVWJtHUcBEJA2GDX+SKxzFazO6mVxKtRaIq2FXu/Kf222czxqoOYTPxWjL
XkNl2buoPh+WDHePlEgnv20mkNCUtrLnLypNg6J8QYmvMAkfy5GHRsFqlt0x
+DElDmyyk2uyvElGnWlEd/cgwDDay239QAw2Z1l47y74SwJEVyg93dQkCKkd
79KCfYkRRYs//o2lm0RB6Jvq90tuEm09y9vm8H09qHFbkfsYT2DsNfBZV8bi
hPccuGZHRsqXL6aIcQIIZUqbUVq/IP0Pz/RGcPata1IjEr7OngCENzbQZgo3
PqoatE9rcV7nhykiJjjzeVAIL6L17jH7COZ96/BWUulmb1mZeBv/MlbkmWjt
FLzSkX9j0XY6+wtVeULdJjh9pxTlGnwYZIamS2/IxGsjdjyx97KAf/9J34re
nFjlYek03Dvnc6vJuFhiLkCGcigceSp2eyN4gsuZKYY54Y5it80q7he+E5EI
47ZK/5tSkg7jZOOHZLrRaC7iIkRJTcpMU6vaP/d732MmlNX7rwJ/qbuYVV4F
kpZ40Lz5eezqzmp3Hgdt9dl45d+90EVy7gKamVG8ZktX7Xt1BhoT41LeD7l3
x/6lGXOiZ3Bxfl02Rv88OA71kY6Vxy9vp3rqorQxCts+z6yP6z5+U7zq8sqX
jnFgPCf1gtvTKb6fiXL+Me7rYH4ljrLM0NpHglDuNVyR+KbaSaFa7/ANaoGe
LJ6XF7vCTjYYBzyCsxDJ42SBYubaMHdIZbKFTFZe+BYdfP2GHKs1n0U+8QsQ
fCjoqvyIH5DZ3GfVyBZJ6UjMIDlgCVDLzVNxfuXMUyu3C3o/+HkN4H/ad0BS
77vtpgO67GOysbdrtHjFY4bsUIeB8Cyu4r2g9KnSp3p5ZKVduVJjrx9EnRjP
7WqwKtohfIoFEl4pTZObr6FduaAU7iPGriERDvO27G5rAm3MIUcCp+K/2QHR
94IZOGsltUD0BYBQxHc84Bxt4XlPj2fqstxaqFEOzZccnnBMANEa+l3RwE8m
LPi+GB9Bhu+nJKJUfwH4IFDYPBH8jKrlOIVDlDlAgHq5I8qjmo/vKcZ0BjdD
l7WYtMYfae/6hRXgwrr2M5219mhc+LA71+qPyVYx7lFCthny1WnazEVuhJQW
R7gqeGJJMVk97hRbmXqL+EtHCyHD5aaYpokbuQ/VblrWEr0v8TSONGEA1PRL
RuD51x6t/KXw6wfwaMoS3dpfUqRd9PD+n2BkPST4ZIMyIPLfs6xGyivMxnnh
BODa9wmZiXVFjosmTIGfeieNUXzEPNlcHezNMqEaFzdbQUgoPti4z4MpxdWZ
1UMiLHy/wTOyFoeNcX3OeUicYV7Cg5bXHRk2ve0FuuyHhvSP3yv2iNY/kB0Y
e2PKsgIKNPGGLicr4OAO1SUX7y8hMpv8g7xU42oEllQ9hXgcNxyrTzAa4VSp
r6MooWiihaWh/YP7E+CWhKU/7Gq4Qv4osrZZxCkSQr1wX3bOFMxVM7wO2eZO
pRIbXPZ+C3Bfw+BLtisd/FpcBTXd4yHJyUtoyItflQvU8+95XCTYJR5t5Gbz
vWhzvvBigMNLOznwtrqeb4/WTJ4hy2QMhot/39w9gGw4nwZP2GDnKUTMChql
wUvyEiU5UNJnKcACXZAQck9+U61DvGeNIGxGwPx/UsuSxdfnzMTqvxEVca1i
/7JZmL+Hl+6W0a24XnyS0OuDZr7eFWcybIXUuE4r6cXxJ3zunLceG9j4lxuz
CRc/uGG/9XXmVnIbhmBT7x89SjrWpla6qPO8i1IGdnucmg8m1lHQs/YImT0V
JC0W+dgVBmKgwwQKNKXGOAzXZhpLTfsYjiPjq97lOcmoWAdebYlqallA6aN6
9NXmmjwv2mbNhBH3RsBbJ8hlxvrvgDdvRr5CZVKxl8YGM7vycqoV987vxGBF
DQEoVc/FMbR4qApC/FEkzjmBNHsxsAvMnpqGiH3LRxd1TQOofWyxlLJeE6Al
nddi7rYTzZYNqOnYSy0+AUpPOGy6xWKep+cBxSMnKstAYhrej7ePqys6swlp
bZRz6o7bVm3z6od50iWr2yV4GOa+CpkOm/ZS2TzLaCqxhvX6TX37reNNX2ia
Qfximf22p1SZ7BFUD5ZrQpBbCwRqAkJBny8D43F9IQG4Tx9GD2bIq/xwsHA/
jeGkWszKzyCrCBARBBmQ6xFpOUClID/tBSNOg1obCf5+QZBxbZS7lwm3zR/2
AB/53+eBuqw7Fbe+tqH0Es3tHBXpnAPpfYZiZd/E4C4Tnh5cPcHid6uPP+EP
3fZ+A/lOE8gUG/X1X5zqWA6KD8fHgXYdOmm5njKzBwYBtKEs7YD1/PikjemD
pE0ESL03Rn8k3NcJ+8+EgvB/kPQCNMmu35c6xrZR8lbyYJgJIPQd74bYBdhH
D9f+YoxU9t6ZVseNAsUPDsq7zZTN+SHSk7G7IjmvsYsAmJc9RiQqDTOs7cA2
CX7tguC8XlLSQtEmndJxEaOYq0w/X6nwy2rSsi9oclpeM6wCJmcR6kxdkAZh
9uxTXbdNxRC2Xs8wK03UZlFWHrpQfhQPHEjpghPZ/BjmnnJgX8udNyUYLQ2U
wYVHakJWeiLmBSIauYTDhODePGg1uMG9GFTlBBOVlObWtyMSYx2OMJbv3IPs
yVTjAcAM2Yl7S61DVVT23Tgxgx6O0b03OTQ97aDYlGIhzUyxRQLNSE4mE3al
iSRw5wS/+0tl/fwO1yQNpxhy7mkAdw7sIrlRrjHB3e8nDo174H+yM74+dzNO
FeqLugL4fzcdKuiOpCMq173+iL6KPGepbgJYTSCso89aUsXeXlsQf0BjQi7r
uYHvPBa8pj6EOP7VONT5ZyqtIyqgWTGkz7e5tpJ2uY2id9+PTW77KLqw1jx3
KziArklBMgCew3p8NIIeqDEFt+DV4mMjz+fJBashjpiKX4kVwpNj5h9ql41H
ikubOYD8so15vZqCeD5jDEBXkUsunk0kuVfALbaalyeGDtWIj9/28LWRRvME
H44HGKbQp4J9NkTMi46ifPz/kYyITRaMumx/FoZnZWK2vxBgplWyPvMySlOd
U0SzF05t3zbwSmcvXP6VQbjkNEnENdMg/CEhgLIUC2Jc02NWUldkin/Pf9Y1
HJXpOjexgAdYQ/eW3Lmrw8h9r6qZtNiw+dYtRSI+gX8Vl5JqFsIkoxfMjx+I
5SbZRoq0cRts7GNa2kjk2N4DaLYgbdas9ShhBDZ1anSXQtMhyrVGr4gG1ue4
pJJPkU9Vnh/8tCHzaSC7jhtZLiJD809z6Z1KDpIF2FqwLqHEPYwN1KS4NgZ9
55tdqq1qf5w48NfBl7OKJMb7jZobGNHigIto5ehybgnPKhxecJSazRiO6ttv
oBFdnPr/B+iyucegUo2O3QNu5NuEnK709bCEbmyngNfTVyMkUSBQ7+Lc+Wka
eS1Yk+Zk3jVI0YRkexrbubgGDwdZ0F5AbSGPQeZoCfIowU/qH7z6HHCCHZIK
G1ee+JVQzg5QTiGH6f8aMNSDT+7PUAoVcGAsE0psZXDjRoRf6N/ZxsYth7rO
mxvSSyO7zkuWTkwWVJh3Sbscv30Pyn3oeHbPyvFpUTPOJza4rUC8lOj1m4+l
rvZIN59B1956oJ0V5l40EP77XxCWFzRqYOP6PBJtqgtkssp2W+ViBaueGpuB
hEU9izNlT0uttKZ5zUcqLaVg9Mu7+agQw3n6YQU7hXC/KyR+n34Pl7DQTs4L
9F60oDn5nth2yVH8b92OJVGO2DzkCGOJmE2xhkwRA2aHeVBm87/1Hy5iBHrX
Itr24Fh445IM8s410ld6s0pf5raayVOE25eMNQlJ0CT4awoRM37EQSoKrope
7DtnJeDH44p5/QwwXTmJVjRo2VQ+qshp3ndFAjEZ6tYruiPjC2FHF/q8ynES
BLK7JHGllWQklKXhuULMiTYsbQsAWp02rFN3XFWChQnyC076jOIoHMs8wxmu
S2c+S/O6YR7yH4D8rsjekAI6Q3Dr6z8J+PIJah0NORAXvsAXTzno/RY98xjd
twztjXtHZRWb3XYKMylIak8KH+wYhCH7GXGdbEtrUX1donWKSpjsu7Vf0yqM
6yedBDdfncUDrtxEmKdT6ilkpKB9m8HduOxjq415HfxijjEgJObZrnmYAJ6e
gS19XLeg4iJ0e0u+1l8sMG2RVHxHfiaKk6IILobL8YuTRsBoC1iQBg/gM/kp
MWxjts4I6tuKJVNgWm4TZlCq/56U1/11jMGzcKFcRRQ1hOGy7lSo3aT48sFm
XXYw1dgICzjnMxEDdNRUmsM8UH4Ay7GBm4Q4b0D+zoZajD/I3Q/iGZ6TAT59
fI64rfUzKc2YHfirdpNoaR9UDdn2rfOySkxPd743w5EtVBXURzjp1ifv+sp+
wO2F6IGpb7DEVNA6tf2UnpmiAcWw1dcFqYgJmeI8+U7t4yenGMQ8mNY0EIl+
pakmBc9qA856Rih83UONc/OIo4bpAqK+ySfKCnbuITQ8LIGA5n6iAKHcnfpS
c/Wz0NY5uP/jBQuwHPn2mALgKTK9vfm/AGTEQpUI5s5+39O4BY489QN3+REV
oq3rGA1eHMKXK7mSpIXtITWdNIWZ2o04Dyld4eEAEcKPQB44lggPKVopPJZ5
5OdyDMcRYS3Fn/0bbDfT07pgUYDZQqoVyvehO7P47QFhs0J2tcw4rkfRkGJc
uWSWFRLvc/mSWeBWXPVKnucqdG4s4VEgJ+9Kv67RGYd/jwCIzAmd7bpYzcNF
fMW76WEMlGzaqHsHmEmRPdtXIpjEQKtW0Bg0ouLOrtBmJFBKNIll1RhEycB0
yA0iLoHugqO1yKdwPevy+hy/Axnv7yfjchksPtPIE2sbD2HcNK5bvFzmDvGj
8iVRHe88YcymTDQJaxwMrKYBcAdvuLK7q/CiEVj5p5dAlr2lBD/M9toIa1Ko
ukYGcoQD2loe97ylRMYOH+LlACs5oTUoGZ4kOw38C8yVPXQt2bzZux2c07ER
qBc3eEbRVMEtgYWfFuWObaCamI0M6+w61YSEsz/DS39REqXgEpee6sSb1LfX
jwaIrHc7rkY8/Kl5ku/vQBP7LTO2P+3uUrf/bKNjTDOO8Jmi1rnR+TM0tTNu
8gKqmwVEaaCSqkYheP9b9yihlgUrlHZQ65zdDKy5sJA2RQZDeW8ZTJOQJXtG
BAqvQJL4fyCApcsAjNfD1/ydJP/kph2EKrgaR8ri21JDo/1YEeibQxXoVcNh
xOZCRVcow+5deGTYLVBlPMhbosCODapBUDiHUYK9eH0asiDH/caACRHzJtM+
p2qUolmD53tQxDsyRpGdYkoAjxADyOS9feiawtCmq/XKWJZ+/LX1Xvski4mz
wv4ZWxQHcn5adv2UOjCW5KTczU6QBqm2jMg2bBwmSYWlOKG379bHIdh34w4z
SJYfoxHdaunwKNp9Ma6AA1msmDA/X9mSahIXRff/iQVEdhJAbWaW+2neyr9V
93YBVAAJv8bkXg5W8sOl0To7HOmlEszfTSlSy5RsanDIFhZb4YjXeYNNzI56
veIVqXRF7CWV+ofpZCTWxU0wXz/cyz7kzeS96aM1BKFmO27RQpvzB38WRyJ1
M2YusuZWrRtWZ4zFkngMTOtYUD5XFToXxPrT9eJWE8krPc5drBv12AS1VPL3
EAZKqCNXz6ayMJRotIR67adskghdWSVb47qnYv2tIv7CycG9+wGAyFw34QdR
tVMuG5v63/c4m/DPBIV4D7LYjo9+MdwGNhsY2p3vl/cw4hPFlXjmgeVH7fbi
0RbdiasISSObMKxgWiCde2HXLPKtGeTA6pBTc6kiWVLsLBozcG3EDQK5oh6k
xyX3DgiJR1SAbakq8EbgbbnA1UOAqQQdehhh4z7wpSeduSRJ/XGG/m8diZWb
a4TLtaIouDSxRxNc03oZnlzw4ZY86RhUKCiyR0Rn40PwQaASFRCD4JrH/mgv
nHsjHqBnKC1/Lvq4uQULIw6qCuKLjSQkoM5Y4px9kxRbnQdRu6pGuI3J0pgk
oO8ubw4bIhf9K4AOnk/GeUP0V+bcH+qk+y6g6+hiDPKzZjh6RAwqc0Iwc+Pq
aM132xZm0MVhXKludZKkfWYKmhhn4vlrzrtnbKz9T/K7+bxuIHN4mFFefa3Y
lXVRknTkNcUGztOnnFSfFQgjKukPJpf+9WJZrSuh7JKBYr5/GPl3UIBu/EQh
sOhS7TguO0dd8wU97XXL1JEaeGYkuJiMxPSNNe00hB8IDrqyfqVpnxrWQyp7
Ulro45gxUFuOF/0G8qRCdOsN5V37tSfIi8z1cqHBDk8fFhlbeo9NO1IKJFkv
3T46pX9T9jZ+pJKZKG9BpanW6IcQ7caYybdjV9DwLR+f8gzJdOoOEHDZqgHH
c6gEZwcS3cCq3Ki0AgeKL8eZs4JY4aOTD3+I6NGEnBxMgt3Y6tnlg8a6ctfP
ZVZw/s5b+lPF5BuY1ULIqspkVR2pDHtA5V++Ja5nLfP1hexHvga8G+zl+qJy
vItwC/iFvpAEBkJsJJd9viQZ+5htAzRUD+ZQV5LJRjLYj3PULD4HcMFoDLAb
rLGAZiRGWB/ZbaUha+c0QDdX4lMEPtTPPD+/9FjnRpVneFdW0DcE6L/8yf6J
I5oANM7GnsTrl/lXc4jewcZAaFjbXo9h0EpZiSnChE8Nzr7IB5JTMNcxo/fb
4ZUENAgfXCvb9lazwD6isV1TSD7IMwxjw1BrAaoN39ElMyxN5D0qBTA/tUx8
IZUXMu5mmpTGQNHkeskVbGbL9NWH3DZDLxExcvWl2nkA4NTmyU/HoRF79l1f
O+205lZT+Ttiuqf897n8tPHyIXXfERMhJ4P5ges2Qg2w5jLVCkwu88rrGuI2
BA1V1rxXhZCgvPlU6BvSul+MyrHZtpicGoaKQzsCM8tUBpOHY+FhvxGAI3Qt
sokVEi5Iri2U5HcGceCKF0aPAaFKrOldEr0dlxeZvrLdLkAFBDBbcMm+Y2xx
7+9tcthepe2Mh4oDLDijIfaaPU8SKI1GRUwvkb8wnpkkYu8+d9B4FndxTp73
w5J+41h38/wEXodbD1gNPsFoHoswyxVtOlbt1lAe1XryrrU4qv5o3UHpTxAe
Y6ZaQa/D/ZMuN2xHO8O5SAxMd8iTgOEheLVEKl0RlQg1sgMM5A+w0WtZY9Jd
ylDorKK07QpYG10GOzqvhI/emVqEF7FIGbw2KBAVkxhbDId4ev19ulYgrBd3
6/MV7fTOsp4dk10OVinQVhZHggLi+THkrxFcyy67dA14QvY+z6+kW2fuPm2L
B7QREtCA+bsK85A25GeQavUh2KKHFym6WQk/GVNdA2FBk6SQTg09Cbnszb1/
OCCf3YABVJSJxbpeypKUTFcTSk4FvS+1WN+cC/2WGgCA2vPsTheF+MLH14ig
OB03YSoMdnEKOWFS0ghqc02ds2md/lWTY1RWcN6po0d0dre1k2N1qO2MhOXE
ei0XAOFUVfXDxs/j0G5yqqlvySQdBx8lx5ZdD6QOJPIh4tjad0C5O/GBpLiA
MbzvXfLCF44Yjvwk3VRFP++ePeWMbF5iGx8MC6JM112m8dhBzH4tFe4unBIY
ZN3Jy9SKqKuXtTEwEhtvhSQrnqXHQtZ5GLxjaJFhqOAP6w1LRn/ekYCdzAEY
LzJ9llBucKTH+68vZ+F7Vl03cg0WtwiJk6v+GgOlM2wMlORk05ZTcr7W++7A
1Zpb+ti7vst/oAd2KZ18Z8JhkHb5UV0+dYFO4VyCJIitu6hxd9DhXt3pNxW9
2SR/iEpXs/a4oZd8nKDIT64VrSatXMrvlYXWnFeKuwGyvrQ4FmfX9KL2LRWG
nGAkv43kROO+dv6HshHczoI5TUZf+sZFSgo2S+vel8jI84IRr1Sp7+TKvbnG
FeupocYF0qRMZcQWIsNJ86GqXwRwjJjRw/qcSyA0S8KdIZyrJ6tO9tjiFKo7
qIi/antd0d3Abq+4qDSNcL/KUZWfHAg82ZVzZfHvjyyUKfGXu50OrcTu9ZsQ
2F2WNz7S7Dz56wa+q4RpmZPE0Pjzzq3LY0h47xvehRk0K+iEMI8xJRHOCN5C
UM6FAS2DMZbTsDbOvCyWzngjuHwl+X94ut2R160GV1USQIFfZQ3Bn9h2Twrf
itZFgc12Rco+oPgrefriV8EybJt+8QE7kjIGPlcAnp55XC9BfGB+3RyScdia
NbU9Y4QBbI9E5aXAtwDbtaL2RxcL4gKBzgRaBrwWh13ABm9S4huVL9X+TcW1
dDujIX6UcNZdb1EjEpjT6colUFwISDpza8ijAqLOCkAy/jWElW/gTw+rp4Ew
UbXlt8E8do34lLKs2f3rDHc+1AUj82+JNT7f/zBPfzzPlBKQYKVUzl9aaeeB
MO/ogaGF9UXRJvVq4rHF77HiDYSkZJZ8BW+U5oPGOTUhS4ItP67K1F3lYN4e
BadhoGP15QXjcd3GXA2CQKfONJk5oEAoE0/3t7TJQNYXeoNBIIJt4DLAb67f
3uAjS3kyu/MZo+jTOOc28WqOQ2/r6EvHJoPbN6li6ukOr5vRlxO0B2dMjBml
3Y2A3fWQnANX1sfMon4aXDmKp1Ti72V+ImyGid2qeJJTE6/Dbo62seez0rEl
cmjp3qinv0k5xRwq5euiLtF3fBdnkeGFJaongluhGz7P9rqVMyR12rBSSh21
rJgU0zyXh2Hgc9bdfq6yuWNGDJo4EDoicwtz9Ern+zSp8JWqZciaY6qg2BJf
POsT0IcRh49dIh3kaKS6PXQ8WmtM1l2najqWdPeGwGZdDuWccmUqZT/01Csl
bDzYokpwXODHbCD8hHF10Pns7lsko9l7K6RdFm2jKHMES1mc+h+YO3brZRwx
V8oo2TyMAQQZqjZzHrsFFWaLIQRJ8P9JhYgMQxmCHP1GMS0a8/f6TuUWj0by
KlsYBYSSQ1/8jvgWQ2EsTN2krm6EE+jt/9uDeBToUR7HTPQ3pTne1MdMPT6W
Tc+6lxvUex3kOt2czSWeTJcojDB6oC6uKkdO5qItohI495kvDXts3rOxtD8H
TvOwPaBMPPRDbha+9fNUHIUeygogHfeAIkyt8b65JIeQzAhl/IuVPyecyH1P
OA5ZOjHWTpO743NhrlOujPkAVqVfqMG5CRTOyek1dD5HxEiKB3f4lU4Zp841
HLUVGT/VOkuLjDzOi0ZD7+r391PkmU5RFuxDcrGasDko8lKZIRHo0608537V
W0FsgTOsOH5Gb4QwJcBBvI2gYDNJAhSPT02+nedZpt214K9f6bTnI1etWKw7
jl1ja5VBeHg4et0tWwwqqquVSC6I8f0csADS80e8geaVcby83ELoseK8Nsbl
dCafeT2lakHiTho80bG57X2sO1y94nGE8u1GiJ1Sp5CY8fFBMnKoCoLzGK9y
oTcDdedXTpTfcYOMS9ymSoKIs7EslUSdIKf5CyxaCMJaKV4NMJwNWQ0DSmUm
/GnRxeyZhoMz947iqXIJMLW73KkuClMh10CB5p5HAT7t7fHg2lFVDyXMl/e8
nIva5qoxwJLBoYnCpIlLarUGNSzLcEAVqlInfAvngN+KJwHhHRrBSsyfWXTs
2eB8JrHB9T78lKIip3HOEXBK8pCEUMMVnJYCJ8Z4T4QUKtZ2lRWvvwcoV/TX
IkF+bdoMEnhF+W8x3QZsz0M5xgsvT+m+C9oaQe7kN/hC2NtNjILV8h5UOP71
zNW6bHCkGkp9IJOHpD5M+kLprC8Mhl4WjItnXU32110LrlnOwEbh3+/HJsr3
VK/zkeKeAZ2Kxu5nl4ObnJNo1yoxVooOyGCyrNEFwK2FvXuuAOQsPoEidJgi
7hnH/OEQtD8KUJTknvCOl1sIAd8mha4WsX1B2kzNw3zc9BrpdzD0IZ2A4zgF
7fpPiGHIPDl1TJa6YiFp7BifqLA25OL8/EoleeRpvGkUqEq1bS/JxEriMVGe
FxVzYptDO04HJ0+IzYV0KgKgaTtBEmay8EJTo65Xvcj+4a0jEeUdF4mcZfCO
OrRJw18vXV8itjlC9mG30MBKlrp4HRRlQLuyEyJRZ0gxE3RgVB8ftU/4yplC
vIeIXP3T5JFheI91iFpX0M+224PX4FhvDiWMvMMHVqONw7O8B05/xEmOASh8
Rd+6M64YBPMfVcO9j+wjF2e8JNMyCY4hby0HrHcVAMIF6u2GRHej10gQqbgC
PAyIIWcylxoV5boN4gE/1RfwaBlGZ2DGR65YAxJkbOz3cHX6e88YFD9K+/5U
3mPfEVk//bef/+PLY0V3+3pM4Zu7u9YIke2UJ815UFcRrGjIrXS8lUqOC2Hq
pOjYMT2OoiINi9o8W29HWm4Dr3cSUvPUDwylEY3uH50mcAFP/m/iw9BSvIOv
G3G/QSrFKKwN8w9FajP8tHJ1GZSYRw2+CJcS0ukZUnowghT+uDvdIssnA45/
fslQHSpCbHssWZ7QM4eZC1qIzXp+szBa7hENVxnkbf8nWtajQeCkobSGp7nz
1RT3RLYrD9r667jmekQ38sXe1elD2ldazCDxxqgf2767AFo7srtNKaWxmK50
W1tos+FlffK3fCXe5Ow3dVLHqE1gqLmxMonhA3qOdCudCLmiQeFyhE13AN69
8b+AAZiu1NxS7ked1CTJfOVegQ4efvF6MGRjzMJa5wHy4PHwcSwp/7hkwCnN
sdA9p0WlxEMK3KWCbmx4oKgAarJCatepe5jGfQ55tKsI+ON2+Nff0i8wtBvO
tR5qQi0weIXkzZ/baU8otu8p4do9DBXDtBC0fyIFNYGLU2zPV6VripH4/ZfQ
I4/bBSl1D1yUgEDvs3hFN4oiPvvC2hb3OmNEmstcMEr48Z6jgI92D0JPwugb
5t70RhcU4W/Q8wIC4MW+z6+xVU91/83c11+FV1KU9ZAtY4Tq3hbj4M8G9Fha
uGiSNgZ00pBtl5r8M+gRbfGGct/5H72TW2PnYoiJUua6i62OA1W0HWm9A9SX
cXL9NJmnEsVTf0/9QbFuXwvoJ/xsfkHZAyV57Ud8+KQ9TN824KmCtSBYSJxa
Y0OUz3rurhdoOuwFTxKMLhKpwGtdjlPVqERdFvKBSFILtOAu9mRtK5k28Qdn
h94aZe2UWAINhAzty3jyuXm9IP/d8F2dA5vzvsRn+jgHAe+cZ8H/aJTuUO7M
O81T7k9ihozsp1gE+GW4EfRyXD4qJx7FBRE79neZcwP0OIrYNGYt9TtVveIw
3GpU02TA8RNU9fB5gSzpJsnoGCQq4ARbBuazZK9KOlyqOsoVAXqbze0qBsr5
g65OR+6o89iWuCIt/S1sFgXhP8CzKx9VmeUOpQH8Ab42B1B61usWi0HW/kfr
ZrnNyEQMxs1+RI53mlm7wlTjGHJkE7zBliyIkNS519JIIeJ6BNrlk0Sg/HBa
/XcR7NmnInstmKM8hUdAn4alAbNJVvOv3cLiQn3Z+dQTEXWiuRrKAPpSiZrV
5Vfbxu2l+elA/zy0NQVj7WvJ6g0t286707QTeb0s6Msl1D3T4ajpX5JwAc0h
GN0FA1KJQRReDaZK8+EkJeUcJZjVSr5sVOvx+rv/r6U0eO46QM5ZbKYjIOM9
FXvfqIMpNsVSvz3XE7t8LWQql+NBYEmRSC/7JwGSYvI165SFGiguQYlgPTbd
GTQRsOSGOoVoEI1b9WaqmF4UTxa+0ipBj6SjcPcmImzq8skQpzkYe8pspb4r
mRGBmPMWVUgsJTlbIjO6lBpOia8XAKoYlpQvDec6ry5bWEdopjNdYL438Q6Q
Nw4nW/dito103Bt4jcrYdcAYynpjeTeKFlDE1JEWqBQlYhsvyxk8DHqTxRLs
jAIl+CDRD33oOR9dwVmT+7JpFelS8vc/OMp5w3FCe7YUpNZJwrvFBDQpWEOv
+YV0aq/lRiD0yzV9CxuY4kAt1xb9/mTdLmpguAdO4/jzHsQ7/3fMpYxBR4GD
WgiT1m6mwL+UMF+FRTjCL0hg87ukJkIyrlvOB5/MNqDb/paG+sMh8UQpg4FH
k+oCMqkgCJ1IdmyW0ijyXwRMIs8b3XPKigshLVkptHrzSpwT9UChy2cLGQsR
yWCpeANm0bs5cp4ERhMGqt18JhIRFeocZZA/i++e5rFy2vAz4u1Kr/CLvXZL
yBrg5BFR/nsMUO9LxfHvtUkdeOqHaj6f5qHh99aAh5iNy+ez8NmPRQoh0tCp
LPQt6vScDW1Q1AF/ebqDkK6hh1ySO9RoJHHGIknBL4VIjDBVuEKsMzWG6see
DNwx6VwxKucyzu0uOVSdUnxnt2vUjykLK1dlSWYdjGCS499synhrUl1mR9av
21U87KEFgSqi9lyzRAbdsJZNFbmp/OFAPuL7prr60XlyG20YDNrDiMALgj/Z
+Hwl/a5mkdm/zOQ9FScNQobh3o/YLm7e8oreg8VbsAylAlDK3tXKX1rgay6z
nFPd2bKkc/O1c9xSY8VWJ2Ab2sxqI0OYMMsjaFekkIQXpa9Wt71nAmeDnGe5
2VHRRcfElS9oscBW0+JE9jWfwxzrnK2qy53tTcXPs5SOwKp1bE5u80enowai
s6HR4unp91BcOj7dMDUtj2SyBt/XIKU46nCBx/zmmdCs/PsOdu49fnnwrd4+
F/nDPFZHgehRo+/qKi7YSHXLmbI6DoH+Z3AI0lgcsCkCJnW4i4k5a5qYyWRX
veYnuNLnvLVanBN5Gd7m7DVCHTtT0Wp/fl3MBQg4RE/dETt+FZ43bwQ8VPE8
bPbnXUooFokM3N28tgZeeCPD9fJhF71/96CCDSF2zFb2UNRYyVtTQlulNfuv
rTprd9W/SVWZTjRwl5P0KPntRYUh6k0K8TXK2Nvvq0oWNRsWMMVvUjGpYlDF
IIm2v07lGmqlNTzWjSwyefUJLEL9yw4fgxzY/xYu/cRkOA/TYmewvYEZRgUX
ROQuBW16oRcYG6/KH/hHbSN5XM+I5xYJDUMpwmE21GHeC0tYbY1+AL1pKTJ6
Z48mPtHyCn0z1oYip2AxwZmbmLkWPXtUuHobI0X0FojrfYHYsc3MT0f7nYS0
r3iNAFbT5MwHbXGyEx6BCXx+B3GY+TB2GmC7jjqLXSIr1hVDYHjIcvP2PVsn
FVpyi8mcWjSZSjtViHt49bUHeHer53ann1txDbhRHwedV/m0j/WRRla55866
FAB7oT3y3APQPQEXNBOqsa9eT8AA8uwhJtyP7+itMLs0or68+ZJRhvkuJZ1X
kwMsuawneqrDRuRghHdp+cWgWGbpUqSaxmRgyT8gkU0lNkGnD3BtmfBiFXd1
AFhc2nK4YI8XYDKd8A6FkXGEXvAiHtpf9Lo9waJZ4C9Fs+WJxJNgMBCPwmLi
YTbuTS0SkWvJI/WngBs6SdPErAF1sPeIgA0QLyy7A8EIoD1gHP/boeMKGoJN
BqbF6TrxzbD1vgwNaM7+MLYLf21VfyOeE787RFqXPiUiLfCN4ZL5Y5vJS8pw
q0iKrJm5yPXVtHVPXGAv5PCxorf4Bnkfv9huFoynhgYZTSkGo1PxyBk80e5m
UZ8AgcyP3fhB2wLvpdquJHF8l60q8eAdIPFxDpQ9sgrxWqM8SXIoCtjliZs6
MbPFr/To9O3kqaifPepjWUg5dw9qml/rqAL/3Cgeox+bQHWbKK+Sdc7PoHe/
YyAsxcwYg248xsQ1IMZtKdHHTcLfR8O2O6SyJd37oxFDXizlcQ4k/Tsa3hOA
JDwRs8kPJKELMQX1rnT2CTeTyaCZ5DIgnZ5ut99inEmzfla+/I0zcVkUw354
yMROknLcKBAVKxaGfihANOIGozpVhXng3LzcwzTNCj4X7MmRbwiGKGopqnbf
LoyTeknBcY7U6j8qGDuzHkuvqsNbFqpJBJAP7Ki3gGmDLZGj67ElZEa3rTUm
nh/nKBUIgJ/0wxqJSx83p3aoYoxqUz62lv4cCHJa10ZA2kTWTD9sdhXyWSZm
0sxowgkDKi9UIrDEWfb3bKuwu3S9b1e4twCsfkbn4lcGquXD2SGH/OpMseFB
q/+79YvDTS9ZZyFtKSWs1fBVTA61KDps3dIDEzNQcGDanm9xk242yb842VFj
hJf0fnaXx+Ltn9XVcN5hy+MszIzNIBcyp/jPAYGkoDzCwOZp04yWonXfeJqf
hr9jE/PpzX96+x2D179vbgCUrvRDJXoDPPEdSs7f7jIsZkM/1NnJZ4HvO+M6
WdNBm7sWmFe6/45hZ7YJxN1J2PJcPWv3R5OH+9A71U4zcY9v4fNhVcHMEVFs
TsQDi2VYW/A9SZZBNiE9NBQnCOic/UdpA0453GfRCEYgCMBzMw9SCmGLOm4d
NnVVRwNX8l4R3rlrwej6IW1dPQQBDxH4G/qlCFjQ8GAzP1+AMkGnqzl6AtP8
kZJt+E+nBv1DGBiC/ZHpbX+0NKVCLaoOEdI0pLait5cv8+sAUSkEg2YPwaFa
a++t2ZOgFamjass93n6sYX2FFkGzocsXE8Wa4siflRoImgWF06n672nFGu2H
yjZKWd4n7gPKcnPCLXopGD+Fbzp9Lz/Ac8XcNB4P1mPursUcRwVMsq5lyfzq
4xk2c8scHUOy4UU64a9XH0JlFsu+xdpLTppdOWN5d9d8j1O82jyPMw6jfQgE
L+F/GMyXMlFT9y/Q7X5LE/RqtSZBqPqNXCosDD3MkQ1tr5EjQIoj5ipZySod
2fDPCKTnruNokS9nYj1M9KfPa9FQNP2W5qXgsy/kZR2tf7sIYZGQWvkp/1+u
XNNNDvClePBcgjaK7EB07nSs4dXxNiWtwaBTDOsq78+JA5es9vWqzIDgwIff
zBeSm2d5oqSeoSSI/IPSLEiZAtI6Ui76BCtakXnaQLeBGAjbF+WNkky8FugF
MyBsjDzFP/fwjz9FuJ9QhrgMnafNJTkxcVY/s67S1HbdRE81aoJZPQDP61VT
iusqGJvqCOrCHPnOGPzQGybfEHrvV+DxJDRVvGgFbW8CefD10st3+5DmjKSM
o+2eiq5OgTgy0KexTS5LB6H2vDC/iJRclG5VSwGIh0HIglOs7L7zuIKwM+qU
L/XIY10gHNAiKK2N54kDTEZ75rEnrQlL5r1WeDfbsQsUT+WwPZF9mBtCbXvf
gRM94omLserf9oDPnC9PNejGyZFawbIZ1K7MZafX95ciO3TA+EpkAYxnWNgr
CQL9Oov50Ryy5Iudxpz4kVQlKCFML2qoUffTuioCeAok6F/Pp9w1KhVaQmd6
eHiTkW0m326/Op2qKM6mW3219MJ3DXG4bFtcmwloyOSgQPdQ4uY/ddPSegYV
P9XHurhzGwF6nW18ROq18yCcJfSUjxSDhqPiZmJFUY//gbojFtnXzqJUL9bP
DGDPnpc0fsHlrPsfx+ZDkAS2f402wMql8yuKHaDLozbB8kINtTC+SyrNojJ2
5cNMLglHuJ4++hwqVvpb4E2N4COkoc6Z/PKLEdXXCNew5wuL+Cj6ziSzljRX
+z52fysLnfWTsy7WJkUKJ/x5F3HeTV0PPwS9ztwyyr8HF57G5MbGLv5ZyJZp
QRiT3tY48oJTjwDb10ZA4UOlyJ2spnhYC7DG20LeAdM9TTm3F9zyOiOv2es2
9szD1S3hBD8Rpxfj0aQ9WGp7W4HkoKdTtNxerw5NNI+27aiywvSVP8AogKGd
0EIlU4xlkTQ5vkfKPy+iCdtq0xADUShQcyMmT4n7/gPnSuSbFHO5rpVZ027Q
ZOb9Y+ZnurPS0pdP6339dbff0Ae5Dw5T4sziqp0f2dSFYj9L9DGrJ5JB58Zu
DTHe3E4MlgDM0fdbuhFU5kCRiaci4tEKoAGTIDzg8VavGSKcU8eCzcniwq6/
+gErMPLIilUAqozygCcbAp7CzMX6WqBZ2rfEYoiUID/oGuT1Kidrujn5vnM5
I40YyWZRr083Omz2Rh9E/hOMI8iHvixnBz3XjXRpW5PMMHbgfnkonzV4xeyZ
LN6FgKriPwE+t5U7UWebkikTLZDvjhWoH6s7Cwe2uClLK2LtcFe41LA6d/kp
nIeLBo2Y5cgEj70RW1jbKBHF7SAp6uRWSe4QjQ6XN/jnrWGaTK40eck6Do86
FWMo5s9ldvAV488pQo9jvXm5IgQTeto5FHUPzIjrvuUEKsqQg5WEJXwbSvL0
HDo0u76CDkNCWTEBUR7iewle+uHXu+SSgKYsw3H2LIW2Y7Y9tk4wueLejDqf
eMP/ea63xJXrCDGpqyl6GucQV3Ittl0FYN3uP/Ij5Kypri9EEI6zjdXMK1Ao
qKRISSivBEDmp95oNBjb4dhyUtzD7kK0AOOhk9tSD0GatzDyf4CGeS86fOb1
LLfH7Y35m0aPIe9nj9qIZuFyp0VxUXMgbvmXE6NYBLFgavvSHiRBCXZoAenr
Fos2Uer64hjyPeLmA5RYUr3ZQdBgCL44kdnVCxVR6KLSc1XVMtMOE2CiHWSN
YCDFDsjt/QDCc9+HwbaMQUvRrLp7n5OLdODY1VZVKhhDg/vxSFzkiwJaIXb2
36/fOcgPNuurw8XuI0ldrccImC09yD+fnr1Sedy2ToPNBErVbmlzHqbhIzBR
zIcTVM/bLolse74axC4CCZSyGebiSjnK2pCJC1tUtlAr+wPtM3haeDrzxLBz
je+eeH7vCrFVQ4sTO2NXz5zF7m8b2v0qiPRsTHk4OAHbNB9lpGQzwQPvTwds
5CJSGfrjNpismH2ATIgosRP4J+gL3JPm7DdR3fYNHDV+m5q78lIZ53iF+YJQ
7IoJ+prZR9g8RKjuQnfqdBWl0V33p0Y6xbHGG1QMX2KjrbrQS/EE5KN8n1MA
aee+mnrMFgwFEgk5+KGaSpgO94rKR5mSL+LaNg9bo5twYs1WwBDsm7zTMZNE
WnaQN6ejwsTau+fwE6C2iFKViphLMuzlOy2+ZaWfZIitL+fmMLs0iTy90OWn
3+u+0OYgwAI+mzqjEEsmM5VfbufxS+KUAQHVNqQSH4Pumx/KSzZllO04qwtp
VG3KqiOALJSU9Meyd4lh3Fmb1yhG6SH3Ri4mVGbb4zlHkPY3yimCuCWpm+DL
u3nzAdqgeKndHl1kXf80R6rFS4ZLsizX9CnMttbjg5gZKxfSXRI1hB3eu5Lr
qu4F/M1Q7x+NDU2rCqDIcgZar4sJZS6CQCjYtSOFynsb1J8u18kdUtjSY50/
kQizDbaL96ZSAxTdcsJ94hbHbJbY5RaZindVl//SrgtaW0FwD2T1PkxsW+vk
vz8fcNrnrfHy1QHKoG2rnw0+baCSANCqVK4cz3KuF8HeKBMgwgCBlgDtcwgb
1cNPZQOz0b24tfUgt1Hey+vxKpBphRGPgIxU2yUw3qDp69D7jeGOxz9qGsKj
o+UvWgc+jrQXm4tknySGp7j8ono+JCuuZpOm9l9neZaisL9vZuBZ82k+cqy4
altbghM9BQaawOajIzFy5ruRG3/z2GZxIlYihghef/LDh2KMm+C48jZLorZR
kFExhLrDN2sVGM8+Si8Q8cf/lG4fWkQUQbFeRS/oddDDvQJgu2lGrUlZx7Bx
Vwbl07ScxIeZnVQFezcLdG8yuhtH1BGDZETsZ3z1MRWnHgk5QiF4yvW+MBGB
/yf/RvwRtjSJCatLkMiV0UUlvL9EQPoAHUIB+6XY5sFmjJmN0oe0JPSO3pl0
iMdcuMOfcU3ZvpcCyWj1yxlv0XvcQcBXnzDjMp5jDNtPxpFOpoK5tZmJ2iEJ
eyIL2JKuYyWimx8kVCRPOk7/iSyQV5dgM8dYQ4QGcfkeANStDR10eRCddByS
kzpccO0PZHsUEvLRoOW+1c55uRmLw8n4KkTXeS0/P/mxADjwDbFcOjHzhZCK
LtYbgZeoApwZZECLE06maGUBEgd+KDw7t96CLAenw7No1Zxr0rlETgXVlcH6
EjrTUFcu0nffauYndmowevz3vfTjVxx6gtTZPe/XRA7ZiLZz2NZMlaNDjhHI
mpcf1dM1fcIZ705tF7d9zneo/ya6XuKFC39ExgEWqSPnIR0WrD7Qaazf7PYd
r/uxGFoc4yJ/YpNkvgHHYEujoLTCfPBpFF+Li8B6KtaIUdNdleftLgiarH9w
Cdvw8500iEkWqoJkfvwOzLNGWoXyW0WgjrEqM2O5WKSMBo0TOgrfZ+AVe35D
bk60oF2oG6XHTfnXYXCKXIZQMXebK+lUH7c2UehL1Tcy3glc738VcXb4Ce5u
ZcT27PFM3NPqKw4c/x0aW5AYWse082WIJBOFPC9js7exHwmdRy0a0evoMy1f
Qfrck+4L3bKXglRBtkZ7JIrNTNfdvsq0Yb2rQCDgDRCwpWNhYvBNqOAcIiwJ
8KhlTTynA9pqgb/SOIo6MzGWwMpySwGr5wKX3TFvJH66um/9MYIRFxd5rp2j
1q/t6GYmaMbrvxvRTfN9OKWNLU3sqVIZPL/GgTTvB7mvFjje6qT9HEuCkNUa
YlWaE46a/Ul+gGdoAHN/jR2wLcg3oVFGKJAr20yQdn+i8jd4v2o9V5wZqJel
rNc/gyquKpT+3UNSQEVG9cbgxS+1aEA8+S7qMgFsnO/1TmTEsSRctYzU0jf7
SOhVQyZrp5rzUIb7mFyRoAJ3aa2svfNPooR4OBZObl+fGZ2rZqXneg+UnY2c
8pRIgQBfa7f3s38L26ysOeCN9mH4QPMbQvhXf8HLQvoPGQ3876Jof+FFAQgu
cO4pRBOupmOqWY9ipeZ7NHkwIvmhz7LQ3/hQxpJH6eRwNVof+qC5HOL+pqoo
LNftCPSaL2hJSlvXJD7KQRX6hDPsWa4S43ZuoY3BtRYFq9lW8PrrG2L3jz2I
7cRAIQUyhOr6Mlp4992uJPIlUPZfCj4AAxp3+td++gn8kFR57l9HZYFb6oiL
AJZiYIR5XF6qzKqNHmigSGf21XoZjkwpdjkLoUhOcTHlNz/BRzqYRS5G3975
xKRKlYmb9paaw+FPtd2MUyvKrm5PRaM73cZKdWaUDwgptHERIEO3baeJr7h6
DUEnoxtMggulFjW7MTeSebBxC0yAaERu0jX6mlooEV4r8K7XRgfvSrMyNCrm
p+RME8hWF55vFD/juskJnYHvjBI1gFzvuoR7pa/FHGqDIyIe/2AMYx8lTG4/
DqJrJVv7lemrBSmfEvPYAcFQ0gKlnjJqJH+4EKu8bBNFt1TfUJASuEUMPPhD
e2pOuPxwlh3i+yaSSSwVCbfYXFHhgoicKx3Gj81p7UUa5LEQENwjb5GLmgoU
nZ+K5PxNkWHFVaRrioeHccPbOIZYN7l4KXJS+1AKv1LdUItXCrqezTVAviwy
fKwrmiyS9yqBYJgPz6tXBcPQQ5G1NqKyNIedBq/0zgv+KscJj9xH5v6KyO/m
afHHGc1Ujj/g7DO/z8ll3V+7EMuNEIV3XFStj69ZT/lE7yQjA4XUe8R8y0cS
FPUvbEV9vwKN9zUBh1m9DFRUKp8WLTbtXv6ggQ5LSx4NGQot/Hagcu07VT/q
PeyXnTuonGIobBbMbQj2lbha1DcITd9xsJMQMVmVgLh43K8T19hDW7FKzZvn
dcb6KBey2vFkAXN7/lO5cUhwth9DqDyz2l/NEgILtHQeGadZw0csYUKMzBRO
u7Fx+BTJQ5Mhv2y+zLTU0PQc2Eyy5qQaFApuKssoZ/ieJCvzMXNqBdIhS0z7
cMPhnK/EJiD9ySklyDeGDlPYOHo/hDVB+luu052B+wYDMaQO1nHqjHg/MWAO
vkrjomRLH/9F/cnSuAezCP1vG26pK/0gPKlBBord/cizLD0EJ9IB19i9fsb/
3LQwf0vepoI7s1W8FT13DbcTixerCUPWBLYlA4UUR7PR/bKjQQhj+M5I94eb
euD2+DhI5FakqXZ/uqC3Fe7yg03YdNG9QmCiNmlJOa7f4xYlLoeUgiPqAJfA
r9Uj+krS0RAvY0Yz2As/HDMQeOWMdrHMlH/QbiX4vt/5hDj6w+Ni5nKvPBQP
bPlZb0bAjSu3DE/HO5yljqGSLU+YL0b5JWZ9np75IaCQFbvjvJ0hmlZaaZt5
NPsuOrjA9WH0kXr71OhoJ+3izpX5+6UScXpeB0XHExyEra0oeK1CYAu0iZ92
jsfDAK8rzaZR3wTTXHgdggpRao3DdUPkOQ8uRuQbAkhda9iDZtDFwFaw3YEN
7yJS3IWWH+lEn8Mii5bNcX8DFEfiC7eAGjVUfVtTDop8TeFNRnyroce9STTQ
SpIISH1Ydfa/eR4vVUyL0IXudh3TwYD+ZsFB/lefO0uhMtNsULYQBeces7bR
Pwlr92lxnbe7oJHGxt7LdtCMccq1E1TiJJpwDoahcxoQM5syCfCzAb/SdpVG
XnG2KKcDMDSCOUXNQ4R9rPYGQR4PKzOLo7UNzrNNdPAZzI6xGzy+mB/7Im0i
+O7vKz5FgdJwzvyY1YM0YUBDTzWCiyWNccDwZPvvgar/KFFoiNquOM5Q3Ms7
/mExoPB6gSwsjtSuwa+sW0hD6Yr500kfly1NZyA5Ohj9HdEC35iVSPszOGVc
l/6To3hJM2vrJj8pfFtUKyXTY8szuaAUKIsZ/hZsRKjRgVWIWdrLpzliVnQZ
S1GrTniYXGdXIK8JNuTO8FOjbISFZWI0Nh4HUxlIzQgxUYsAhBGUCV3OVr3d
CN1WkElxBkWkU+3Bn0nD60YRJOEH1Ewcp1Ovrd29PY1YGHO1OET3np8vVZjF
XziZrBSLVHjRfL1OOkZE9UD7vejRQpPtcLpuEPZ9F2CGFN2KDcGoRyMXZ7IS
NBqz+jszxhMQqs02/baaG6msBxi1dhGEYwFsEh5e5cOr98NE8t571+a7zovI
Dnvzg5MOMyvR+Jpitq/IRJz7bU06VweAqMFn6aWQS5CbgKC55haXGIIALRJ2
QegRelPlzHHIII/Z3UN95CE4PqKi5Vb0dJH0p1RQzhhFPmQbWOVmX2dYHiXH
tv1jRCIDMh8hw2DWHTDZ0nnCPdeWpBPce2PNXkKFfTnJm9nskulpKwCMtYqu
K7TZqfjHMcSSMBpm4bZV44jRIbIVNhXDc35vLT34h6IOJUCQXJeEvWEWK+RU
H9N0Lmu6IQdxm0JkPdQEFuTpVQMP94nBx/+ApQKyvj40i7Sv5kdW9Mh6fn77
YOYqMmoBqjg64WIQIDdM1cYvyNfIEKrgcuH0F6KngA7Ei+kgLlR5X1VCtzsV
gdtz1VFc3io1ltafVa3CSHHF/ojGRfSkviLQUvSDTK+5D3j0+wW1OOiG7laq
bHVYVpmPC9e7/N8ZdoZxswPuCLbWlEv6Uz+kJ6C2yywntV/5PmOidnD38fho
nQbXFIHyWPpkNku5TNLJ2Ge8xADS+3p1+z7i3yZGO6ckkOQVko/olBtoftru
qLYdzadQxIyexnQH0oY5Sf/vltG0KgIPEywhugI3i5CqqJcd+ZPfOpWUHtDS
3jsr+dmO/A0giU0cq6x+c5Dp67xbLaMlXzAc5kfo2+BoAKg7bfMi/PrSYRPs
K71fCV6DJAk5lQP0tGiZx6PylOcqs1ZSlGSjIAJ8cUj7IZtvHGQCT8yAwBIM
u/L+HVgusNPXI/BCAIKu4oakV4s6f0Io7aQct/dslxJocJPZ+hJRc/J0FLc8
/RXgNHjJ1px9XwmPQQOZknVPYehJaisJjMGMT8/gVsr8ltl7l+6DJ1D8nJyL
r0LEr4ZURsMzBlzsmRoawtOoiihU6Ymnd94Mq9ILaemXT9/FbJCcJJSa8694
WecqwVtL8UXpdThBc/r7Nc+qq7Kc/si7ymXP/xoJwNCeFSzTfuN9MmyJ+Vi/
OvHPeg+pYk7k/qj5mbcW/chQOfv0ii8yK1h51sXvcBcB9Ej6TrALoKMJhFtE
G5K2ntRwQ6nTVj70k4hahxGDZoNpR2vDonjzEAJq18PPT9KzpQY7HlJr+Ypx
x3z2fYW2NSe5hyBwKyWHDZ5cyKHXV5birfyf237D/X9ijld8qj7JybwkWWWw
pBqbfKHtZowMxlh0WS+YirfMDGmTLrB4FRZXFu90sP2H/+WBlh6HKW0vsvmF
HLQ5fNgNRY26yYkZNn1fs2TPrPIqIIDEjM80UPMblfd1GinyQn4PqycbZR4s
GlhEquuEdyNAOzwwEAno9iMe4UdsY4Es/Ffg+YURW63vY/IGRHVMmVMlbe+U
RggninmAYDsUUeA6aMXBcw6HyiZTn34vbmK26CYwM7QZ2+fxzIkwhLiV3kJw
nc/9Ckl6rfrVnDuHKZmOLBZlIeVIaE+Tgm20asuUJagcpSsPcDCAGWzX4Xad
S4qFuft58z1z8c2pQnBNUbhaIiRDSzEmAu8gK+sP+0RIOHbRta5vGHAkV4B5
ntM+DX8Y8S+pfZAYcDbNM2taHP0FSuydixgbkwWWSONJ/JsWETkLRQbzljPe
tsTJaVDhEkHcWgBnMqfbZspazhYzvKfk2ewmZYKSXhEQZYeZq2Axlz6m0y34
ySkRUtKBe1Bhm1amSvTXqE3BZXHVoPMucityFJqNWefLobcPX0umZcQ/Ti0E
fsQotQwzHrtWS2nCMoTPotQ06zkhWUmobz9TI3cNIyTWcD9zEqXI8zYE81G1
FqsKZ5kRy7SAHy10VOPu1haPqFZvIjbHICZ+YyJETEVRHuKr3oIzfsQWayXR
5QveJHqHs0V7w84PMM3lHQ9YtPVY61Z/bpxG0x3WEMgICj84xfWYR+/Nu9VB
sZrGjiliy1HqZjbjrcMFhljRGY/fZxd+0QrU1RM4eCqfUBSkCa0RJm2if2vN
U2dqqSLGGamoUY/IDZZeOfzxslvh6vwkgaaiT4WEp7v8uWJScgdzg3g5rg61
OLu4Z/L10NrICzN/TfMbo97j1s6k0NaWXdqdi8jHuKVnxnlpN7X0thvZ+H+L
pwphkoSkBIdkQhRjwdST9qf0DFYIwdPkpRrCB0c5/3xv5iEuou8K9JpesloH
0oTxLm8iB+KI/8HQDZNFjx93Qvi/q26v6XT+MjAWZwrGk/9GCVex/zO0O4Ki
wx83SpM5qehQ22pWcI0h0+p6E1Zq/YLfv+6D2A22G9aa3cLinz2Ht0JLrZuA
Ysi+i+uLLdqFq5cXaFXVtYWaDDLLuP+Ps/pGEcecB6OqkBZu+eSWSeXvDCTp
1idHCBKMSWhSU2WFNPUNwKa6phIetNfWxzJxtXqqRxgNcO+acGOePDL7zSSo
lZaqPxm19SAXY11ESkA+dAP062k5WsG64Ocnh1fbcgyeMBCSbBUJ876FucwF
2iHBT8aXTZUiMvYGosinxMQ1AoRJ6ye4RMxEQ38QAV3wT5MlGixXZ7b8pII0
jbzI38bi8tPGD3dsTxqmjl9EqbbvOt9Dns1GqLMGhhOCwC72N7oduOciULB2
j4GXeXcW1QQ90WMUZmDMvrLv1FDYmzvMTsPJfrCfm9/xEsUkb9nfHQCgozZo
2Irt+ylic1dHPpDL/EnpUw8Db3XnC0I0u+N/eFGChaaR3jbrV083vR7AThDH
anLRLf8mCxH0TYSn1Ivd/qmNR/b3FjTXoTmcl6TG013jOmsaoD4Q6jno77NG
81l/bebJ4Q1E2QLcvzpOszLJb4H4dGBmqQNAIGVlpdpQDXk2kALuQF9rENIP
VSxbtKAs4iVE4gqxenCQcUG4BXR+/JGkyXHPX2xkUIsQGvS+YwS732NsSGGn
00S8dVCjBupC9pHuewml0zpWfZ2yx0O7EligPwUGHHBHcypzXnsEBjzABc7/
WEqS/vlnXmnpCXFyfjvN/NoNjFtTmy3A1Fr/1ZnENyx/FOr33kn2uTbIneDo
Osd0z7CIYESqrAWKIjqrB9FvjlTyCI4y8CTfL6DnQSv1NZhEaZvcdNKBHDsc
1xcxPZnoBV0ddiM/BmjEp4ezkxYfYXsozKdnMPP5FFdRWkgKAHHmCowCs/bU
OGPbCMQ941Va8cn/kJ3llb7Jk99I5EiXHWBJaED4oyM6sByfcwvjFolO3T+Q
1CquhNDBvikXHua0o5lmhVf7uyzTJ6Tr/VatpMwMDzMVcLhllqfEg1dAVy45
VTkkfvH1P7AzA63zap/jQokr3gLYa1fEu3EMuqjC0+vl5W3893CstnV67HJs
Oe3/qA33JCiCsezwcAo0OtbyCOB6KdSh7BRwdpdpIPme1ypWJ/v3qVQcrWZz
piP7rf1aoCVRsDTzkxSOpaF171/DbgymJ8to9jdQYw2WAVku9EmnsVRZhYSx
jHdPOBfD0hlvLQX7mksGJr1CR1NyK/P2xUKMTcOI3QeXyTdxL9nXhK4PMv7p
PpIaLL/yuQ2qX8mBra5vtInHoShoN6I412uQY00P7i5dnwN3xphPRCKT619I
5WTzHZN+QYuF7cwOj6W6JzxH6yOwhSN1xmcJzDe2NEuYLSDZjAl+T43V1HLq
ikMj64OcdLLR6jTHjjvP+pK2Q9pDfw0AXnIL+nEBNONUXb9OwH7x2Kp6lG03
rAMjSpBTSrrGEVcTVmpXvJuwHdcpMbo26n+FYK8KSGegCD20YT8mBRmOJAgF
P9vO8Mw6sKKdu1U1k2ZSxhb1edUz+kJOaVYLphzq7nD1vYUP3XUTaiwCzXC2
xEYSHrvIrWojNTYvLeku4agBECLC7njFnx56nFQbHgGP9+fdBNe5hpvic5AP
3Y03QyrTVgr1FFchtb6LxoVp7TKTqLvw4fV+lItKnR7L9sVNBPOjopU4NBU3
Auh8vtRL/Om0sfoqj1XVX3vRsghx3M6inWnL7jeVmung3X2J5GqJtojOW9E6
xs00ipM47i7zZoysY0kB8U1rMu9d1kixS1CFqKAMqg0yLyBGa60+EnKLWiXE
LLVmmbbt1lPLNwB7kxHjfdDTFYS93uHDob6s9qT1km64OsxBo9KXVuZwBfgY
Z6QZBaxrTd3TE/E3vwsqhM7kFEeXIf1wBTML8ej8vzG0IC4YSwacJi20zAbL
znHFwa/H7Os3gwQWtZXc44dTciLU8U3kNTg3bp0cxI5j0yODuj483x8UhebT
daUXjM3LBHCV/YhBV8/A7kzJAKsoQzIExIOvYvcqoX+akp0EbH49PETe1pSD
IBBaNFTC/1hs9iG5JAHAouEtkUPm8DUxABggU4/dxm3ioLkGcH1lUU6McPPm
/JbRBCMTQHZY7HIUXCN5s212QGYnSi7bl4t0/zBPHHwwDBGkBqFtDnsWoGRZ
jyKRr3DwD/SEZhCz4BsejvGkIQoChFqZAJpo5GnO+S21KNO4a0SJk2njLVK4
VnhhzDFsL4QxHt/up5hDUQmySXiGPVefzes55GC+qpyPkYPCGOR39/7I2bZg
zm7wXD8KYHXe3/oNV6YG5ogjS9xEDEneplI5+ZJGPq8Q5jWGIX0OU9UD9Xp9
PvuGiQc0ZUa6heKZcwpK8dplPO7TEIEOj4VkKN3z5BpAzkC6cwuDbXqI4IZf
QQYafdq3iaQRG362uEPIqpuN5856cc6RlF/4CpgMHy1UWeyZ/JZt1xsriqBE
vsq3ipAeml9RBDBvMOLLQhknGyzcp65/qkZjiYxIez0+tBWtNOw0GBCTp1Y6
ShokxdBGJIOSVYM4AZJl70e/P7ZE6pi2V8mTGTcl9+7YaPnVvKHtI/uZO8ot
vcdkfSTzb4mHEZzus/5XnX0xiQcyzJDOcc6l99gh06y1/UhoLUQTNtQP8A+6
rlzauoTR6KYpjd1W1LY6G9iW2TrexIRpgWGeP+MMBdNtUkoFMafY0vYQpxo3
AeUFCccR01w2FnlRnw7Mxl8DXbOImXw1k0P0CuUwe0UVPqz8scyn/xRuCaQB
VgvQTTAJoWqOyrgsb2wnGI/GJ5c0wWfZqUnsdrkjHbGoawXNu3hAuQTSRdPU
8yennOP3TTV1Dki23UDVz2hpykjmzHKvd9BnFRSToyneYEWZ9VTVjQIqJZBs
S2ufjRopdBTYcfGgD7gbL+xBYfvUYjGPcZQls3EPRfrzgJMvWO1x8kohdj/8
GWMLyyaAPexB81DiwY95lJCqQkHL4tQHoljXf1URinx4PD+rZ+o/BTLWfLn0
Y3LEmDf2w4SkEhz9CN9Xqv1XaUJ8cUiP7HkJOWY0K8ds+uGF1djG2NvzHKRV
zfAVMB0cEXm9Qi2oifq0cOVSrklazmqGptHcPCV8GQ4ZtZ9mYqpDQjsVRpPU
MEv+woTzXYF1Hhje69uzyFgVxAODXA2/v2yPpp9l8SPTP63yib95+cbjkjRJ
6fnho6WNaOhn2++thutXiUliXmXROpo5jlO5e+TXr9XSm/QK23NvZGjhQnKI
9f95fEctn7UfWaojFKjTEZxTbubGwu8/VcpXgyFMjNrsB4GkUlqRPX79hZfJ
eZ68x9a9U78EAWOiXJ16Me8sicYML81rWSO7DvXIsN2UYmbp/aMc7rYnVzIi
1LuqI2Iz1bYcKp4sKkbcBgfo3h421mOY8kcUye9afQ1Y91aopuzi6woNoXw8
awRlCbQ4AxtVJuPxQfubxv04ntBC/XXA/yRPOLwqu6tbCDF7GrY4/m7z/rD9
yD8OYerPuRCK1B9Nfn2MBqrZh3jd8VgALSSlOEJ16a7KYTQk1cCD6m8Nr8BC
On2DARiWOs+MOyMXy/7WEgRtv+2xbCEWD81rP5lJuIVJlNppRwpnyZdyeM68
y9wlZfJioFBxFNgXhXy/aOYlFtA5zsU3dtSBSYXvBQgRzDXCmzHXT4WhjUYo
OCvZWBxhvfVxdP4wBYk3Skk8sZ66BgnEg+h7MQajKso7rXBo1qktm2wDLs9a
ZMK5aV7VqKrtlLwyRJf/odM0S4LnCvbD9y5Z0s90vCEYS++r46JKnMMN850b
Dshqjkj7eSGT30FWpLH8y6B9R1PMNGJbQET8bweOE1/Ymk8L2i246+gUizc9
BwEOShmkLv1XrSlamraGdr+50+MUIZvLPvmw69g8yWvXCR1m3S18e8SqPYU0
mwQ6+llWa04yBy4zUtJEQDomlfOjKlDJH3kBpbXLsFTBlUWgfGE1aWIS6Wy6
/0yRqyfvvlVZsDYBYQvM+aKoc8fecb16w+a1zorUMkarSxfaA9kXaVSUoY5c
CEUvIHgKF+vFXaPlRdlVuIWsjHWlaaGIm/WSJBaeNtiDe8tiyDurIGOkz44/
dlGCaVprODFdq2Z3lgTvuCnZQyaNxtAYII/wVEI5I129n7XbtgsNFPBHMeF6
WDHHwDkvHIlDS99K/zhMtavwFQFQZlDIj5zx854z/Q9V15PWi8hO1jAexLbc
yz3iuntYGJEoIwAaA5hOwMG0AjUAypfvQ4KbNr7H+FqbWoak4Yj7KGpWyqfk
69ExYCP02b857Kt82ey8OxQffGTv/2v/EC44xvRFAa1hu7wuJF48H69qKjH5
T0GeoG4BLCkRnglVzrMo2alBtqgPo1VfkIYmQ3G/KMVDbOdFH+77Hj90Wahj
oW14apAVTsEpfXqQZG6LW3J5f98Svh4XtEAPgDm2695ssLKG0dYpnsVvY7Ol
fa4H2nFBFhPdLe8edEaWkhPfsQAcQU1k6tN2AXmOS4pG88rHkkc+8euPOH3A
Kp2/3WwIXeTHyp6r68TUJw/5R7FVcwLISow/Fg6V1ysUP9wG/QH4DLNb8Uvd
sccp5lLCTFam4Ie+AP5ZyCXfstswiTODhpetFdXNP6UwdMR4vZSPVdrzKvHa
bBmLm/zw353n1z44MnD0b+YaTPPKm1I6R2UzkhqN++sdz5F7X3PSQM/mtbK3
p0OmLVJJNTRpP4xw9HWvnVnzFumnuZPrEEZvkgIfl6lnE/fzlr2tnQOj0k6o
BXegpFA0+gfzse4Tlfs4SUjZGnoYunMSXFUr/+0HdtWcCInO0HUQN5shALWu
zxL7la6GVgRrt+lHsquXp8twkU5IXptCSopMyd67Hbd/rtKoT8Z/nIjBDqtH
lA4n4XFQXm97js0bHUNTHw3P23fCzYVsWsZzbDU1AFs0iZrMFhKkl9yOBVpu
Q2R1HI1l+n6JQ+jgY/M+xmme0dVm0uAuvHZWH6yzIAwPMjMTuOZL1LvjWrul
cGFsZXKG/PwgyUUbV5vIGYGQEm4epAxnnAbmTDj9zVhkzlORELFCjyfcF7c8
wNpksq/MZ30zvpxGV3KdS0tYxqYowpbRnnI6ysV3GL5IOmD3A7WtGwsndydy
t4zt7JqR3X8TVpMZyF7Tzr13jCwuzC27ryoAWYsh5vss1I6NX+PL1hJTrWp8
7qJQkU9vlPqhN1M9MgmkJdLh6S+4RFumAaQt8vXENQ3QiXjwATLkVKYAL5AC
aT2LL2KYSPAfabNJWGHVjjSG0/E+RIRt2BEXwhoxtxE8z4fS02vumks3xnuV
qu5KcvT+huWBkhsjs7l0LWEMTT2Wd8FjQMXCaS/dImAxdFFXmF7ZrDf+Z83y
HODO8qQbWiDk8/rjdIu0jPHbde5Co+m+49BBnEUWL4gS5fN7e5ORI8AnPBXY
NVr+YccWPwDamw0hkDmznPznYJX2SiBQm20LmORh/oOD7Hc0keYkO5BDbC2W
fCNeg30LVCjlZda+Y7kJqmt8X045pXdDZW5zyHvY32e7Zr8kQ9WMHn2FZAld
M7FNxPMnfJzTPTMZAo2925VUgVL4mlu8iOdm3pzqjhM8jbRzPBNxnZNGocee
kjsP/AWRirSTv//5bCkzmSxwcf4yOBwOWjK4TmDU17i1c0AzXhW9pbNYbmVP
BOrQ0jYKVrSeODp2MKmeH/fyExpUamafH4S2wuuMfRmS37HapqpPwkcQy8Qv
7owP8qqikd7tTuuNFUFcio2zFjc1x2f/hTpXciQUBuDMC8zyBQkoC2Y367dI
2R6kGrVE00XIIqw6GexNTA6f+6LNXG2uSGlf4A+M9DBH3bF2rq++kIBAAc2v
g8n/stKRSyx58hW1Uv5MPmijh3DQYpcbUxkPbiuN0UDmAt3Ibd0GqyyvziGQ
0UomdjSZNNuEjU6uS+BJi6pRipa5jMHcLEYBg+QFtWa+Vd9a/FN2tOdo6I2e
hw9q5KyN6vcJC5rCJNdYIHgBlWsOF8V0/W9y9N/x8Q7PfDuKXk7jR62JuMk5
KJurGXw9NlrmiZevHjJzf/NwvniKjMfHZSE960XFIoWkVgDLMfBxPDiNxTqF
tABBtimHfYT+/VYo9501jDy3OBa6UlsngTa6lACCMPIpPnTk965crzmJq4ur
Dq5K2BPP0qRRLnfSE4qZ843k6zo4C+h0fbe6B0FFa2qE8s/nBN6556f2MSkt
Ou9sas0j6Hg7gX58NV2Gv9PADVhb47PD6Hn4iih8fUBN/JiS9T5pI0V/0EGp
5RnwydWPGrX/Ft+4uTa0ntMHVxf3rDsUnb/PnM2z9fjfPkAkqh44B6e72iZe
k+UX6zTTGykzGF69DDFPZtoXwPFQDhBcj5oF1/cLaYoKopvZpAakQf2O5Cl/
7yx5PHQUzIypUdoPTYipmV2yAPMyBXkVKahtO0alR+nRiMKWHlX2On9MyRzM
gwl99KVUHXSmC68jxPBREj6AZaBkSV6Q8Hft9BWlsJRYOV/UIR1Bpoe3AUvs
s9ADaXMXQivJ3qqef1foNB3NcV6Ij3q1s2U8EYQluRp9m/ashp2MRbkXxUYt
H2GKkgFrexrLKYLyu/jRQy8h4Breuk8+Q6mEg0PBJOU53idlWTYpbpfoxCz/
MpmUqo6jWfbuUP1BjC1AQvWz2iA1fMZ150GRL2dVW6AmvxgyXgUNGlKG9xY/
s88KRcaU0tN8lews6kV21A5/0+ATgDF3KGVB9DK7NMM2Hys+1lMt/cEPXdCg
ZfXe2VxXUOgNs4lpxHSJ67TfIkwTnsG8s8BFfO8r0zoyOcScn7xuVy2BUO0Q
V0w/xjWqQnDMk571u5kjp2mEnWwrICZmaJy8hJVOi0tO0Pxiwpd7ocVw+lnn
/KeS1FFZmxn8X4yDmKMibOvZePyMdBgI6yVR3WmnMgzdO57vR+05sEmLz7iu
uVeXjdb9CSLiGOaHtyrUTZoqU7ZTN7njYQEckArtwQ+1wbg6xQ39m+zXoXGp
vicAKocYjxyrer/9LaGkaqH1GdA+PIHigMMdwAZUobHuh+7UM0EjlYa8LFFw
GnQv4rPP9oE8deXiTQAr4zz+/Ep34hr8MVPuO07s2Wj1Fhx7HdjYZC41uYFX
eGqrqj3UBKn0UCRuslBc8Zy1GqfsLBKIFVSOSqyTc6JvbY2n3JyawTOTqEFs
TyEJvsVHFzEXRaT1ZuImDd65RKcnAuLOGAa0bNEiJ8FxuUcXDJkCUCpN7vQM
o4U7Zdo0Wt8xYzuD58tHxR+E2JqDziA21BYcquDxxRO32qXfvz420Nmnb9lM
ocYDmPSMzdNEXef3jXwkteWX5Tb8KY5LYjI6R61QNguBI1F4bj1UXhi79iXj
cwcSLbLQymZH5MjP2YoqjgsY8des61o8wdtStLXBdN5twEmcqOEJgShWCNmM
7yE4zOqCUqPwHJlJ5ONUfgQdlEvrgTMGTG26j5o4t4QshTx0mqXhXcoXGh34
cc3O5Z0UUlPNMu9uW4h+lNsw/CZKEZ1PfD9AqO8hxzymRwp5FUlqwcTejKIU
lRVqkOuX2B/TInG0q4rprY+iomcNobKTy/sOyjfW5bvnVtW5xoY0PlBHwv1Y
arYFyVCiHi/ooT4yJuY8AVY7OW/gkcrBwICLLQtCW72C3B0pIApKZ4v/gt+2
n817T+8Qs5ogtcwMj3k95t34RdloJ6LBDlEnjiXavLAitNSQyWGcwDlXz1SM
CegE8FgE02IuSBJxsTiwEAsLrd4dTAJf3ej0tUfYzEiHTqHkx/tqNhK2YIHz
Lu6/WuMc003VFsNtJ+ROc4LU0PUt2x0pras0PoPSWA4b84lo3CUKEvXorugC
ciFMGtvw5rTjrDWzTDheWBbxVboAMgsYmyS4hfUJKF8efbCyZDxXOUOytbQ9
fobMDHaVTd46rRmjQbIG+6WCta8Fa8bvwQpd6Os58JAgcknj3EMW88lxdpj9
5daDyZWhB7V0AZH+/H63ix8RCBnN3d8TiStltLf0ORnfiw9eCtxB7qF9hiBe
+6bw8xAL87i6UM4yWwNVzZ+TvbFcalDkF17xaqjA20fx/MDpG6NoA41/ZjMD
tPfmEGf7hyw/S/uE91FvQMYa31h6+VMSWAthfTnhB02U6FL5aZ2qPw5iT63Z
1Vy/8CtaOSdxBNBFC5F6PNBDdmuQInD4WrloPmjUPb+/SUEN2fBg9ppidRN3
Xv/UqMUdeDDu+l4hk6YyATXwUmccAgAlg80+LjajM+4pkyC107fJ9qEelRnw
Ia2LfuuzP5r+VRcFOiXRRp8SZEI8TPExYNTyOBigbN6/oEuxxdMERW5NfYF6
Vy/O2pOvHUv7V/Wlw1lfBm/TMoaO3gcxyVQI4MIm2gROy8O9g7S0cWqIonff
3/BFOx4QWGF8ZC97DJmjcQj+bp09NU65RSS5WmsoXJ3IuRKiDeUrR9v8Jz7S
8VssxgdnmmlTQC7+BkMWHBGs8stZplUNacP8SxATjhjOPp9vEUXUF480XzMo
X+rVnSxeNUe5TffNnnYEChr8vdD0+jXbMrL5hm2be/6Ar7256E8sh4YZxtAE
j1kzyUj2IhJ6Ts2BNqToOHMBetKJP6wVFPN95hqcuDbP124vd4qpbe3PQAyn
piSVIik3BPuRDjDsUCahD/H7T6iJruaSjnA/4dheJPvTFSUOisFzDCMuEBST
o+3G8553HCtwNP1vmuK8F+KzDjHRxcDwirYS6LwYpNXS9JzwO43OKznTgxbv
/BMtq4UC1ypPNx+HlACVuZ2HuR8P1N8m9L+hLA+SBNtkjO8Q2T57MgHaFX3I
L/XKUXlJQ0GG+ECsWrE0L5Zn1+R1rdugKGBcCJ4o9jH5+b3B4N+EDsL7f3kj
i0EkEbz8GToCF5ToRDP3V0wyDGtPaD1lyI+E72+iess3lqOxmQaNQAXDq9jE
nLjcdxo6qi2NVwr6Qh9maLpPQrnbeeMURWVnJS5t+ylev+9LX2KRMpta7xSw
dMKjv5xIP1hNLNmBPkFHohax2hbTGSZYKmHswKi4cqUObOCJX2hAUDfHkYUK
mAUzwSqK0oLhk/izoeJkOzcRzbDcSBB/QfO+NWdxnMSxBliG5OsS0Vi5nvoE
rITkoQgfooXGHSfvERe/oNh6gPsDYWYM4lP26qXPSbyAu8Axw1RupoTonK+W
jxzeTwMWrjjjhWoUGnWaJJrf8cpogV7sLQaHyBi1BjTZ5ML05SOLGw6GdiDt
RMEJOtLOwC+00CHBZnXkdqKIqlD3tHrSYu2cjZEkusy5iW0c1J5i/4Qif64C
Xuxxv0RRIkrIUjyRPRAlb4ozGZUU54CnI+OUXB5oG/dVgvGBrhQXys/5QJw2
0vMmZa3FbBpurUA2r49xP8geVBetgCh+/yGmjMaNBnCdBRXpSKAp3Zr2mNpQ
lgxEDsusG5S5VGrVcor3uXCKOvqgf9h/dQXts9U7Ma+6X18AmY+MG6d2FDlU
C/LtzkY1X6t5L6KQD2lp5r8b3nVcbpKceJiMXxcHBbhcrBLLIO8HJa/iLV0C
5wePY9V0yIYODihJ7e4azSDIiTm4NCIcXHRpj6IKl0ICgN8nsEN/xxiBy7sB
xCdVIqlV65nrf00/uiS7b7kmI2R1DxXMU0fLkbR/DLL6fftb65LIt6WpLNvp
6z/Kz9yHoIwUxxlZ2lJETxREXSh/DMqruZWzWltpj7xIy3eAmqrgYgMUDMz2
BKGEC5GM6XLXmFlHGZkZA8GV518N4lSrVRmHahc2478w3k2gcGRflXn6EOZU
VBCu+/tCwfZJw8ERJu4X8SbtO4Y4sanccUqYuyiyL3PV4IGy5JfNuhiG2JTE
qUgpiYptLcQBq8eq7Cu1HRsqVFuazrDBTkqyyLdDuSms+b9vJeSe25UKF5hK
DByFqOyniozaRYAYJNSUaWby+uodyBaWVrbMqonO+lo+6gL58iq/qDVSYkwr
EppuHbA5eXYjryvMnaTHdALaX3BUkANwixFriiRGs2b3lDIBWLkPjmiefU2Q
JfRJjP/O5qKt0Sa0u+MGal14S8GONST417azJvB2JUm775NbBj3Msb2b8Oke
LIX30+omZPOIZAH1dty7rmsqciY765ZanUuzmGth6K//7/X22YxPkTH41pOr
ywiS+h42BBruka8N/LcSv/7FXX1LxWDySZz+g961Sy8BGY2gI14PJVSQs8a7
reOnZkdBnGnY9KM658XER2wt+HCnFFOYafWplpndgog1Gsa19/J53RVqM0Uy
GZaC8npRl6Tm6N9xfP8n29XiJx6W9ML6ib8qk1FoWStjrsbVnN/6xYGnk+3X
M3dzWKKZld7yApQVjijxLYnDjE2koAd5iKh54o29Gu3D8iHmcMT+688H56XK
7dAL4IEkvc5/+DmFfRVIriSl8X7aQXzXxU+h8eczvLuzBwIuH4SJyipRxUfg
xquLLVipR63qvZ33lNsd05MYIMczrRqBkIRJO6ibeY4UrP4bRIm4NxiOYWbn
vCQuiFjODeLK/tduaZBYzgWafsUDdCu2HGRcm1NsCsuXEPif151stWuzGzjN
G9ktK6VIAVGIiGiEbWQIb+Y2u3chAtc7KaklIkHh3HezHz5PwEWVZiTAJszF
W5D+7M5HFk3PwNUQPl0kXHGXwMfneV/hVzkJvFK1OBvBuLPC8IqMg2dm5X2u
jlDZQhXKUds6GvI3CHZo1G8a/MfSC6UjK3hDr61LQ43LByUIIbWr3pRLUSxP
T8D7mednH7rrgzHmJFZKMemxdiPp/YM/5ojhpRUbE6upYETUFC8zl1HVmvPT
EX2ub3NRNZFVQDVsw5PtT/t/cDAQz7r/zoxHz7gsclK7J074KUccv5gEGilW
w3/aC0cnxnWvlqfuWCILNTS+fpTIx3S2HKOPnz6PYdj3/h0/fcPoYcbanEfC
GsEO25CuVqoxYiQZrJItfe/U7k+A0xVqxKJ16dI9wvZC/ZhspwG54UcqNLIQ
49UArdIkIJ12Rvn92U7oO0Xb1rQ2w14TAlK0KLQjih1xQk3x92mAcEUQGqD8
q68BSelOW85zkdxiupVmOfXYfju8hBQWnigwz+tZ0z8ol/Gb7STLrFLvy20i
0jnx+dX7Cu5CP1mq32hQ5Y5jMKBDwhOIu1N5shc2npa8twQKTDLplG9qLN4J
U0Ah+uDpK1fXNoJUZwt+gde9i29jSGiFFVwc97xpbm1WaSB+WBG7HBGG9peS
PxwXRbo2PSKy1R6Z4uWgM7Ck06gXp9Jz3qDhrwDXsEcwx4a+ALvksKDKAZ+Z
ik7i9WyQc+VwV2zDGOnroeObMFoktFt1ryVKOGZ5ApGj75ej8KRL6/fX34vb
RCmHb8hAdOvUyq6iSCbf4mOntLKI7xr5yAH2MdA90Lf+I/A+JCZuqeNeShRl
SGUmOg2Se7wAq3JKzNUlL+GqYk+uMZQ53noNS8Fc0/3GTdrvkVKVt7TX+9iR
3fRqzmbmPBwWq/diyhNnFjkvpDyP4yTAYjR8XfKHJSmvbrX6gF4ktN3ax+hE
RM0eCctUwRpjHO7Uhvu8WXDp6Um6FtvahwcqKb4zxexMcduMYUOC340ECnjo
kcZ3kBxuY8M6JCz2rlJ65wG9a8JuxnlX7KKXP8WMLzNfz2Ue5lUZGPG18M9l
4xJwPCZOSXc0pr8i99KFHOEOXkfBpUKBhjCgZ/eNHNgpjiyZIiJWlFEGF/UZ
+HY8jO0yQwRvP0I7cXANat6YR2hQiYpaau6+h76SdsmHkZUw76K1mRlT+CzH
+QSlnM5LEnSJTIoLD2esnxDsQ9E001R1H+FrZiFqbBZ4JgzMRxip9qBdjNDd
UFnCouToB3L58y9yemWArQSDe0PqRD9CX4/g1oiWhWmMeOm9FDSAcbHUKRAm
FMw5oCdqfh9s4zy128hmTnY0m2jzKbSk4QZIBtUoMjR3nBxUvKBnHI1FBuFa
xJreboEtq9Hb1r7gagVzv5RBlgvwS5ACmfzzZTeFDcY3s7o6+vKGP4nvs5xl
miXNTbt19SgVVmTpTtUFQp5SYpAHPANneOTxsb9gA7lQityVCukgJol2e+Hu
O/8EmzgzZox9/0fJoU4LSij5wh0/KQtIFFmX1Ow9BTL5fJ8W+3Gc4yK9RtbD
JqCAb02KfIe0wWtfwIu4b3SptFxkRYTu3z8YdW9letM4ggWAc8ibwkRu9Y17
Wguf4git2BzCIfto4k1AAt1yuUmr5Zx5fff5vV8zJNlNraYwVKeszjTkfKwE
YN79nU7zkyNRvFqQRD5b3gD8j64XpYie9Dl/p062bGxe2adnjWIEcU1amCzn
3kIk404CZnH7B7z9DjamFJmVO0T5jCDR7bh6En/sQmokEJSwe/gklwntNSGO
qdAu3h9AnffdRskvT6vhdfJd7WkLaRnLWEg03OmVxUE4OcJ1WZ0iPY+uEadU
B9pAGmGdADK9KLfYUkVQSJNkERrp1aeA4YwDVjp6DHkcCvQyB1ejdMISF88J
I0TfXbOpmzeAHQ2gpUSrhEwISptZpxm5WYlqjm88C7L/y5jINZy/onF8mu6u
H8GoEt7al1J/sncpSV9nGBHEaZWZ3YdMiunoigZhL0h9Hbo/Yoc9vQ3BgND9
6ve6Xgx2U0SRGcyDgh7JrB0IMa4UTn0TqBfnXhD2WYx/ii3nZTlrcptq3YdY
DiJubhke/rjbRoX4BHSjZpKEQe6oKqfIBQIa9tLj/sCoSwCTMS75l+kkINfu
Uq2GdNq1q/Sv/dsKShwqrOdu70w9Oz2Y9MJ71Pri9sDjRIVVI3khMn8nZQFR
Imsrw4vf03EDko3QbzikP+GH6wkT0xfPJhgYGoLcPC/UBIOvnJmJboJN2EMt
mzukq4Huupd/8zRNN5pVALwEJLHIt2W9oZhuacWHjPV1VkrzUFST2SWuqq1B
O6tr7v9QFwEWdQdelSdieXkcwY9ufIreEuE7zrK+DbjulPsRyl2CihMv2jYs
8aar3bm31eO8a5U8oO2y3L04ojbModOD/N+7FuDE3U40RNRaj9Ne382tbMf3
SX6Np1msAW8Nm1wBGaXOYL7GmS6ykrb3F+y5FKHVsd9EEvrKVtty+3+czuOU
pwFpP7U/34baSBF+CbVh+bRuOFS6SDyh8MLlVxherBGMncswxrBqI1NVVsQn
FJzHoNSPl5PpAlBVkLQhJUuAxOxcBQ0avsy9SevvUZcbeJiAd5RB8G5Dapgk
R9gDT/NDHytySjnze5HufBvkc8YfeRz2lTg3NaypqJZNOvaHvEZQBVB6Xp/N
8+iDvxF6LNJsYkSQEt5ZNSOr4cZgmHLwL7cMQIXDR62yIz9baGDKaJqp5PXI
FLL1bB3Ilnz12+Y1a7W1gPCDZP8FG5kPTqv4TPusUFCJHRbOyN9O/72ph+x6
auXtBFhDcdUbDFivyebDR5eXXJXibtaAaWChdj0jZj31uEfAhcTcBuCRwrai
DWEt2NnvD0nq5Z0zqSG0PB0SLdCULExTaE1sDvW2SLYW/b2QZl1LIQavzQ9A
Zb5B7sqYWf+PE6o/BgknD1FdegEdtMpYowWTAdFlFiwumRMP8e1DSzELrL4J
M3af619gtPAgZq3bgPQ5CRP4BLkXtx+/FQ4FoA7YdZU2llnVVdpSCYWq6Tno
YUBWtqhl7O2PGx/L5ZLafMKokMMWoOnuUxt7+P5SE0ht9ksS8wUDZz8mJEap
DcAgJjJ6stGGd4508yjhjVk7u9Tp9fMk81+Ur96JRF/yahv45I9aNFYDdr4m
3cbRrBDe7vDRjRdtQeG6fI1k1Ufw3NV9aI3QXudeZ+KAHyb0wDTbVAyJglVC
52cvph1OQKUZH0zHUfdA/8Tb1DAqdg5Q0qfoPYCFfRc72tR8kCOp7E89HuaQ
Mb3uU4Qa8mheJgnsgUg8mEKTq9V+nKwdu3TGDF+CqHM8JVx/oHbuWc6JUjYD
yFxdMJwzoYXxSUGkGDfZ4FzDoYJ41JzLKMN/jH195pYGHn/kCAiT3gU3ITJQ
JxCN0TXx0PHk+Lt0YYewdaYL5HO5CzaOH5B8IUZqX/1eD2piV/R6Uc312hmY
fQdGkwIvDKBGgQ25+PoipFTG82hGYC+aPnaPshvWmgf9jyJzG4XBj7+jlRN3
c9OhaVasCVijOA3TCok0zPGsx5qZTssQQbnLhVLJP0pqkYzFcuD4eEJ57muN
oGkAiaGYHbTnoNW2thkukdQGixHyHe2OsrrDfh2Dc6JWm2Epq2T86mrn3gwl
Ao6LjVPCewZs5MkEdmj3bVsPVF4EIhTJCJM6+JpBMk+1N9uOqArK+M+utJVo
KbzEfoZGIeWR66iCqMaSrxoJbalU7DOhQdTiQIabWK8w6VYHWRHbLL5f2EKC
SdmdZXfiVMwU8FKLzmBpgZq1A4EvY9EoC1cY8lB7nIOQW49naH1u8hKDqXR2
EvQBdFvFBe0qGcecWEVK4C3XEMAOBxY57aKxYMxvkIj8t3estXNEfBTQAxSa
mr1iwCQ9AoCz8iOT4FFcpSkPiceAtUjydLnIgCUKKxLMxtq5of123zRexX+K
5jCHmoRqqQmgdyHh/4FGs2An4LSnNYLLNv8OAF9Vqw6Z+S8PYinlN40Bzxdu
DTMqCULxDMUuPnURXNlNpu82agvTcXSjgIwp7Extdf+v2CdpdJKYfsejTBBu
sPDuqpOivV9abLiD9doVE7XJvXppvN86pioJiKw4AFyPS87dQrr1ExqddEQB
cYIWPHpOoX5vyyjdDnKZOoFt/Igl/DjZ58HF2E+q07PC5gdBJg7K/CLTXQBM
KNYJmsGsVMNPImdf4XHllT4SdT4ERXmfvHQtwijbU4jng7gWfIVGFFMYNcRD
DkWssHZgI3cBXJwkXUjRQGhSpxk3ELywVvEfQwCepJkYXQJzQRwm/LOJXgy2
b89/fD5En0DPK65jQBheOHwIdTO8CBixbSDafeoLIb7JMVLkW36k5MkfeJmR
2Y/G4c9vHuJS/xbaQV1oCHDmvv8p9FxTTcWWdLtPojsD7wPPg5q98Ldte+Oq
/9pjd9GgOuiFWgAw1ObDbDbG9/xyL2nawcgPi+IYTPRJiTRqwkhuRsvWQMMO
aW71aeyYcFww/lo62erWZSA00APXf+2BG8mS3vY1HXiLagy1Zk8hJQ4foowi
cEsKQVrW3RS3iLrZznPwiN7ZXDxJlD0+dL92KnNHNy64zvcPBUPnJjMDQvwT
dAWbWTwH8Mkq28go/B+4qdNp2TrBoNypoB+dZBmghuZLYbNSpsoM4unlKoTs
+evQ5FgAnSsvhUHKhJbbpQal5MsWoM3ofGyb3lsMHphfX8096YKiYpoaoY9g
9j6cqSDfMtSClsLMpK+neGUofsAC5h0St6wj0h3gxZjVlsLCUSPChcVcde85
eP85PtfRL7zHfVXfKciC1yiCM8E8JOBQw4hZaEGhivp8GGkCSs4y76MFOysR
3Q+Sm7pc3zi6CWF5safI4+IuYjdXRewMfrzLcY+BiW1zUbFmRFlZ8wxPIaZ6
+D0ZogmBwAXAePAlIIje1Hj0KgxQh9fgyiFBBpuwWRwrcK5ERI4360mEvQAw
oyFPHuzMlqlEvWE0+M38zlx7yFtzjAoDZW4LLaPBkBQOE9cuf0vJHEv1QRT7
sVH300WE3PLw8rOdlBchmhXPvLsbptqaZBOLUaL4Ulvvda7VOh6Bfn7VtIwP
xkqVQaXu6wCJF5EbYAbWtk15ORClIp8PZA6iKHT83ixAHnm9kdUY0dwPjFy5
n2GHiopR4OklEhz99PnNdVpCDXR26JZ6ghcJHTu9V8VRpIiho+jyWoXGB7Nm
NSag5D0RKf6JvYgD0uZpWZ1I7C4JOsSEJLfYRKeJLZQoSvHWa2/cgiWt3e24
ZxwAmJyme3o7i6/n9O8P4RVzwqx+Cr0LKFIc+uWYvdFq0ecWqPzv9TSJW0Jv
ZgDNZfyjR791SxLiz35rgHWw9oUBVVJ0aTZtLYUrnsl3Knu9w9f5x+zpUedw
jX+ZXk/sWtqOJHJfhTftUoiTwECGn56RmtNl2Q6KMdmO82hOQUiNiUB7NXia
gjfSHRmJSxv6n6wUXeDsJbAHgyo9fNIjhLFrXomk4JG/BjvpEBhPQV9fFmuT
rfekr7EfHxo1x4zMzgAPY/oRl0UIetXEWrBNh+xUlUM5/BD1rNfAa8EHd4kM
VrfHssyoDiHlVDY2OeF+VWeYD4eSmFrnZrcJrDbbTOtrEYMrst4v5Bh/JW5W
dv1tvVt4rtOIuzIyVO7jfPOU0DlUuXov6i536HFVAAHx7/Ao9FzvrASS/b+I
wGSttENJCuSv8WieoYIE3nTJEnfh4y1DImkNQuzvq/naTtU6VRjQsoqMVcxz
lmJ6q56nMWuFRvmd3VWiCrOxrBYHRbiaPJcB3mXeDMeBYko6IA+Y+YyRAkC9
d1FbH5SvxJ7yO0woaS88QfX4xuQmrcSrkvPZYDGj7GoVe40piX9KpRih5fzT
xcyYdZkbmKysAsroSeFNSezpQ94vVLah3GouqRXCEdATYBj4JCaUktHEF+t4
cL4Kt1YxVHjH5NofglICfQhNGmO9mJp65tb+N61evYn7qO0vDNrsWRewSRww
K3RVwN77PVc2Hua0rbzt4/IrtshM+iwWahzOnXJkgAxsrsxh8rPV4dlx4jwn
kvjWNkXC90KXSwLBJrzoAFTZGAuDEI6Dr8me+TpOQ7hKEEi+WuMLeDbI1hPa
jd4mOCEH0UvvaVanry4ZW6hNnp0wnQ3r+EwYWTXKrPzUfijZ2HSZ0k0PJdr4
hMBKGYsGWpMMh5+k3W6GGTNj1A4JnX4vKGK7K47DDfuBo0htChvyXKRef9iY
uE5MTGFNiU5hXfHV0QRoRqmaGGc/rFqycpGC8eZkF6aG3RAvHK8X0yvGPEen
Au8rxsycJ85xuv2r3hMzMjnaDBsZ2MCS6UaC7IXl20zpj7LOnopFO/SP+4MF
pPZDCGXhbLoTsxlkBqmQdZEJwWCqIlHLMm9OVYTAOC6sTq210XbykJ9TJR3U
IRk18OC6WmRRL63rYiImp9JAYl6RME9zNaER5ZjQSssvTviHXzD9I4yVjSos
ULM9xeFzH3xHz9pUT6aNFy0FfVNyZ8R02IJZxD9ZcFVaH0iBQ4VbAM3v7XGx
+WdfQe5o08HPKfxT3PVmCbTdzi4lRzf5R365lZNkD13rb6groe39w09xKPkr
yv3rE9Gr2esO7ulX4N/4vAIkJxK2aGSG9Wx9zFEy6CVRRveIenmMOhEmMq9J
tYYyOTEqIzXoc9zywL7tjwyz3bm4CZ3SVmmJEacGePMrvJdSfo/+1tdIc+AS
6OR4UC9w457Ozwt46sTERREiWNervQL/9pkB966t5JsvADKhX4hBDTKelS5s
fDGgTH/MtbAFnaYJ/BNxIk+v2dYcmDvXMkhVBEa4+a2jXTPyDWNIEB+PpodX
+kXgNlt0Gn4mGduNomf0Mu9/yujfisyz9IpmtYsgllObaYHYAZq8szMaLUx+
oB6PChRCEpi2kRpwXwPv8muxiJNsIGqRoaPjm5auAgfkhHkqOm3lGUum4VeF
UBB8QbPMQSasmSfaI5WwKrEHov+mQ+9zomLZNPXyO+bypuzYrsIfC27gyCyC
3nF9VuxTl8cfGLMsjOmLbn8HuIqrxTY4hebY3JN3orz+iSLBf1YS3amw0mxJ
XGqhP7u0/Ov9V4LKc7IFDZivwkc74cLagZoZZjEMZ5v1/NkJLc0zlgrRLoaA
T/OE0R6NI96f0D36jMF03GrMLmShIIJEpdPp+fdka+/Ct1gslYkcyqIsa/Fq
ppnhSbNIMHNqSEYsSRNpgLTkA4SayHlAfD1cZj+VPYpy7WHjQCk1QpWLUGNQ
LtsAEeOkBQa8z6Okkj/BQaUzDDht0t55rdBuGGibbsdqg5Ccq+lqn2C9CKoX
oE7cpkddbNBOZW1jMfwROvJtHtQ7n79b2e9A595zmjisI69QtvnJFWfM4wdA
FIBn9xNwu58pxOGMXCfk1id508fwi0SfxikmdbIYwtyh2/Y+MtOzkJ8mMzQy
sQ2eKuYn2P5K2I91YqHJ6cvp6b9uYI9QOV3wDhmAnJ2ZKZST9Y7fW2SOTHQp
FbNtkAH6i7vytl97qosCSmz4sZfKkS7k10asuBrvA+IGfdlucGBq2xh0tOb0
3VcZdmTumkKP1qyUSH3+iVfnk9ThjX7HFPVCLZSUf00urENetD23ZS8woTvK
VxHtvTfUOUkjMN57pLaCGFKRcUMAowvVmcKHOrkCM/lGiCIs65kdZfM4Lwkv
gzB/dMSt11rwjTAa6mBjbnB78oIA7Lc9Hbz/jY6IHVHPwKYMuggkNBuFIEjI
T8F7Vw8pBwC/Jc7IQ0lcgxYlV/yWTyumSn8hI1OEAkE4wWFLLL+dmLzj1V/M
PBR4nKzpoSLUUw+lppzJlz/fFgzu5tg/8kzzv/NGN0vfNBDDpwWR9PYDur6a
ncakc0lK1KfhF9ueocryh1/azoXMotDCJj4QdxApCsThERl89O891eS+uECI
iCUuxHQoK5WGWnavXtwlUwwxn1FPEdB9A43qfnX97aHsGz1GMTAGNKoo5LT5
aRYrGv6kpia5kic2K86wXu06sEW32TiZiOWJdZ1rX7k/xx9HYelYbepHq8zs
OpyWKPJI+SOiM9/I2nXS5Z5j/f/kwnBexyznX0NUdk6BYVOwvJVWzbV3yk1D
1yctCc2iAORGPQPeFadKWGZTS20aF6X2sXnxafb7LX5lQXfeuipUdy70Yf3G
dJmzEEoLbfQw8QE3zbe7Zol8Vffu5WHn6oZMFZH9Pj8FQ1Qumh49qagU4xT9
N/FYcrS6telNRD6uOr4CstN59wAU/u5VhRjT83iSaUbrT4FG/PmwKbYq5U8Y
EdURRbxo/FLLzhDBzbIH8KzHM8G/YYLiTCACEG2rYjqaP2N7ijFkFdHZ7hGF
BHNDkC8yaNoGyLZFiWWn0VgMsJB9QgwMIq+l8lopXd00Dwn6EGzSrCxkx8I5
iGPA55IRyeBvgtPBB8E5Mvgul/NQWiVImrM50mCeyFjuXXwOZyO7NfUSHRwt
A89ImDeInGh9z6YEULGxRHnFqBTqv5vPXA0PcQiDPwbajHAUoUERrQUP57bY
eLtclc8wPaEgnXu8VuG+L9qzstkcrsfHbQOzrXC/rAOwKuZGBnu1xF6gD35t
eK3I9ojGP6MI1IQJtnojcJt+EsHIoVX7Y6W160ly+q+B4jLq8JPFl9AYdgP3
s4zkp6vBxY1/O1gpeUhpl8C+EqL7GwlqYr2FIvWwgy1VuwldY0exIMlG/mig
WSY3VGxEUBbFumPhNHw3Eg9SX7J2tChsnbRXKPDtC7EtLPhMIheiQxRCQ2T4
yaOjRQqnVRHYgmU31H6JVgerctJ/1lZz9jd/k/WEDNrnRXHDZgKrBmn1JTJC
xZdx4GuaRuNlNPTsRArkrS0BgvdEmZIqs9AD1vs/8T/aintzOf7Pa6vVusIy
6yslZfyec1L1PvltjUvlVJzZUmRh1UCXQeRFaROf/tRNM1TAu1zjh6NTFszB
oeb3CK0nzg6kKck0LNbg1RgSvi1s3ljCBv0MUteObTyJYjqKt5EHGZs+ry+B
Lvn8CtQG72FKfeLdN9/KiFBy3hC9w5CkLOB+78GdB5iXWJ/aB9rvccbAZ4M4
+jnLGN8/OGx4ZwEmaDHSHPitDiIq9dVI2SYuEV+jkknM0IeIyQWOkDlCdfl+
IdjN0SyDAe57No07FqlLndcE0cAMoOOUUJ27HxnAuFGUiF41pKDCdXp3sxt6
gXtteWxCEKIO9ycRG5zAyUERpYZdZh2/t4psMoUNYWB1nvDycMhTWeH6tm1d
GUtrVHSGg7lo+X6H0tWIvFrxdM0kmBtU2gg1qNmG9k1Ek2oR16SHpWOlu8xC
8Zib69hnd+UrGUdMBdBZs8l4pewNJCd4xG0k3lOdvc/JlxemqGhvAufZeWEO
0zcicLQx2XdbjwIoH8uSd3S05Jrk++FcvGlMw2Ucu+/i83GBth1Mx/QIrMWH
SUlRn7uXIpMNb0biqKY9Vtm6R6MGWLwg69qrkQCSl+3kplRrloFlgjLdr5x4
u5wzCQJfbzPpKMW9ZxkN4GLh9QheM2VULfaq8JUKL4EdWJr7JxJjGjezZoLx
xNNVcUZxXo83o+OjH7o0hnyFIhOGakqkeh4K25+CG2pFvr954pEc1Q4HiQXU
ZsGCvVaMN1eKbzz0cs3tsXfjdzhHQJTW3ZMq8ZJNStMu+931f1TIGSHYyAUv
NMbth5ljlFCl5dRgnphp9cRYiU1nY61KGCPufsUmFNrD8IYBFIQUGpxR2GuX
nCsAuEb/ZTUMFjg9VqvWtETPbZFEV1qnrN/uyiKu2uqflBCOCJHzkbxvR2hN
DSPGEH5VkGY1YhW0E4UhxqXaHJzqMITnMCrNEPQ/VgaQiR+RXTfaVR4aqwNo
cz+abW4JI5MsBy2Ywnj0uUWL7p3tH0vhqNEDNt7gt4LPdxBVlqV58SwYdNFm
qZINFsLVjQJdCl6wbK5dDi7DsmDR+rW+HqcTCiOw46ngdOVg69XkjuLLQBhS
k37MjzfY7Xxlf2PTk5F5oPjG606bvnthMGJKTx4kT5hMEPbOUs/IE/AjCas7
BCF2JPZuis2MhDvnPEkGztxFy9tzlEiGpeT/FqXBS1Gl13NEsAUqw1UoOdoV
bUZ7FK/WU5lDMqSbxKrhrkivOdRkhLtV2w+H51O7Xuuay6Wbcyd3eOUD4i1e
hxLc4N6pLOMTRJmDQd9d0vT62w5etw4ymJ9czAd+rmCIcagq2Qkmo0CVfbjC
oi6NXi6yEs3F6Uksw1HKUv6J7hj6ibrI0EOvO9UJPnt2SXeiwV7YOzst07Jb
ZCPjwFZfXXun31dk/UKxC3YAcny0gtxSPx5v2wU2dss4XWE2XpBdvwCCl123
7hI1QfrSt3s0vMn24ZBBHqlnbUNvcQE4t42Itskn+DsdNLrJJDO5U7b4uzN5
n91D8b7KDifgNQFCiC1NbCYoGxqqrsWu96QZbiDdV8kLcUoNxiBEsf3rtBSg
hgxpw8l5FR5dFsFG2wZvU6rjCHDjARSFe30OSVz0jPBU4uycWZuuPDRU29J6
rtnxXvW0CvBwtTpHWn7qs00tFe/vZxNrd0I4R6zpweX0pXBVGvJa/KV+a44q
9CKO/Q0oKeYoWMxgB2ZWEBzEbsqT0YXOwoA9sFxlAjpSNi9xSDYvN9Waf+WK
lJL/hc3BCkDrbImH6aQI2Q4dub358NyMmPz65OXeRdrKnWn7WaKJNmiov2JX
eVALF2fCr15anluUxTs/BKFN2xx4yI/oJFzsCKCxE9q51FC3HxyrDOOdBnJt
cPSJSxhiJSXFK4CPPAZ64Y+e+Lf0Z2svhg9yTzxBzqcECdpRzPEXBKqH6P6X
Fupvk74v6iCAtID8PlxXEj7h3fYE+8x59ygm6HAxVQ9I27SY5LANue9+BdjY
/VYaQi+qpWVzzRVCJC6MNzwP5v+moI/NcF/3RByBl9d2ap5sxwi96L7hgN1k
Z4h3oIjOoWrxRUS12f7OtoFT31W5oqKoAKefPa5M8+xYEuJoUDcWnRcHQ6Pm
Z4G5crI9hUx2sFDDo7+0iOZ3ERzCXrpGiu9jyhmprAVda+dlO6u6RXrmifQ3
obFZE2ZivcBJ0mtt682ldjWGJYppPBTWqzDrOic+78zk+G2VB0Gsng6j+wMu
3Ougs+UGz7p+WjjuFZ2r9bjhuVBpKooZMO5FfDYhtBxdzpI/ytt0wy/AzSGT
h/wssFsHQfhq08orZmUxmolZGswdEiBrj9QXOqoFhC6PrI+hpl/NdKQce5/Q
c7S4DSD5HWUXPMv4/s059+hcy8vEOGEkJ98meL6Hr4r7R6TE+zHcPWBV6Ezl
xK5bjgJDXFNB51GB083YuKGG7wBiBtvgQFz72/QV829HoZTWMJv2vVfy519C
x0Ufh2Am5PFJiyzO1I13qRKxcDJnUuo4pXwaoM4D8AyCLOoP2MxcpDft7l6/
7wvW2eZfdctsUt9J0e9u4iGPvEXkFsRKhbq66qGOnaOZRCV0sf+rcDGBFGSp
nkgXrdpp1BPELjUTWMUWVerYOra9auetd6BD/XbMQt1FiLiK7Ehw3LeX7Cb4
/SLvfTKkzp8kha9/9CmMom1TzALhPQvJdkjPrAMur3hND6CdfHCFQ9ubAQWv
YZ55eVuVsvToMknczqeInSXEDuSOpekV0Vzq1IkSK1uLncgDvoJkAo+98yiF
QLAfn0id9RaUkbfRSw8JsLCTzckDdl5ibaH54b/0w0GJYOtCuBG4My9th/lt
HtpC79bfzZsDgj+aqdp2CebIeKc5ahIEQbfp/u+9b5vOa0vKPKc9HjX266MM
Qu4OFVk9Lbeg5l6tGFK7WBZzaR/jOZIOoJUZn34JoAdOF+lCIdpn2OV+HIbg
8XpP1mj8LGL44IKb/HWDXUi7ubb5K8WFUkMw1DCMWL7E74AyXaVKUgzLpFXA
angVb20rCFFW/hht2w8c+hnn4xAzF/Wph9jKHnj5i/Xq8C6hidahIqyC9fkk
J3G8Kzx+2XMb8Q+OUVqPdsqbPTO5v7u9PbKpJr5NT+6lwisKs6TTtcDCyX/w
0NynlzqIk22YSBIRT6NwyL15rctVTA0sAj9WdRJ/F1d2r6j9i/hLIYYxWsPt
D5mTyEV9UtqyuIEvZXEJ1HD17VOwqPhuYiHUhw0ZZECIFGak6Mu5sFm/Byit
NKFPfGnQ9Cc2W5EXyizNkqPS+x9Y62oxvxBrLRD+LSqUtt+TG6E/3hXlQ387
0sPu7Pf0i3xfOZzCAw0zgmEXoOmTRk/FmoQ4IN1DcbuNkQAISRqhmjdE+8JA
9/1XAMXoQknUwUwVGBKFETECBVA8uie6M8gMlj7BqK4TcfV4FdIuSrX3VhjY
gWjpqT1EPwzTI0OMwpDfb5T+JCgLlh7fKrWB6tE1xiIneEcdmmywmTEYcx13
fQ1abGiykauXcxUgw+4Zk21IFb91eVHCf6W//BDDZZpVCw8b1/EY1C/SbG/5
oXnwv0MsDzE1bQ3kDm//29YX6Z40pchpGykW1Uq01uVOO/JCCoAkvs/egfXS
cbvLJi79SMdMyQcwJd1lswpcN4FbHlRsl28yrGyrKEfC8xPqBjSTwhFAXmcs
HpwnGou2JjqYVCmFuHAlSozZxU8kd4M32kxgIayMP+vNE2muftF7tOSGnKDU
zJk+G1ttPDXJJaty/tNyFJtTjA1lWf5vNu2evCz7lx2ETJ75RE4NzFYMlCXH
ADpW6F4xmEik2Lc+Ai5ZQX//a5IZB9QQnJLGOLyWDq8AIhfI8eRWtkBdaA1K
gxGahWWk+GsJ5K7iKZIrJiT0bptXc227khubSoMLLYiyRGxbUqalzt2MQsec
atHJaczUW1ytenifBIIpcgqAFM5Xe1NjDjNjmzGaOmhYU5sHEQQM1B59j5nI
OTykAF7ZdZo9RSWOywigEm/40/KY9uNGalFGNPQWe1Vjd65GOp4FAIKj4VOf
m2JKF8aKYenhMfgTX8XOHAP5p6jVXLHrg8+rpNJnCtezsQohdaXyOXJ4do4r
nlo8tkx9Wj08veJb1+DksuYZNRCyr+Q70FHl8b0Dhxg+zg/1+63sf9HyrliX
ylvfDxOqiBQNZidRFHPvfPQ6lE7Ei4pxrAqC6OTJEQv76/y6wpj2i8eUaNzm
PyvntnYTJAr5GOBmxycItX2iG2SKdb+syO93hlRfHH1BekYmAmWRRF0Qj90q
rUgq2kAbJfP0trDQT65SuCpAQ0kuJvRJJKHsi2wQT8MAcdgtzjFdVv6f1a1V
g8qTIFUJGop2O7KZQ6nbqdG6LbheBgL3wTPPJ+JCsSs8UKTjmvbQR/ShVPzF
+Z5BEyUeCeIg59SWAWxSRVRj6qhmS8URMnPx93wyZxv/RmyuBwWSNYFejPb4
HKsZKHkYtaxLUDB8eR5ALkVywizRsOEM0uJQAkMF7bjI9Zj91luYRBgFYFNx
xCqI/7mto1dagx4RLUDqemRCHa+wJ9b6BuXUkUTrQVW/+P7sMrvxg7k8KS5u
wXNQOc6jxZMbuaUcZzYfUM9XGY3ZeCypwiDuaBF1K/Fls9se/RJuMnjGOsMP
ZiH/M2kPR7182Df62FGeD+K318htxCRdj4/kGrfKkgMcAcu5uP7hW/Z2u+JU
qmhXrLH3+cREYkyl+ihxBEWpA70bRE+KRcdT7nvsnTA5DSqjgZxaPWL1iqwI
etlRIaBwy2zVIWloz9xVK47lEpprvGth8DodK+3/qjLOIksqsMXFCk2NVrcJ
AulFKUX9+udr9VeDLxTBiITlNAFl2hQRZnPXgSM30QLBZJGPediEXBpK0I6A
p1+S+x9EmiuSJ2hO3qGVkNm9ZLn6XWPYtUuR7ylOtKglCpomn/SnKbuPTUMG
4kML2vR/GyH+mfw6yAFs6xYuOQliVUv7eq8+AkyLYcCsdMC9/eRe1lDFnc6j
klSnN8rx9LcSiF01NtU8Wsf/si5+y96vZplwY/F/vABD/ReVTGAD6J9rgvg8
rDnZvpoY4EyW9+xufVj3EEbIKs/e4+IHv33XYDEdVGVRQwOo1fGiSTxGTKQe
QfLlgN8KMOATLIe9cC+XXtqLqBth3DV4wSRaeqhalhCyGpRWQmKFb/BJDK8x
6ByiitdDKzYLLpmJweplfSjSsOikzwFlmPNZXzJWiTlO5CrgXOZ4ve8wePsi
1k6NiQuklKDldO89VT2zQm63I6FNq42WPvo5lm27xNq/Ip/vCuSL3En6s1y3
lLUwoC9w3RgL1s/Q4WdHwILjD4qY8hwNKhnSrSnYO6umbljxmyNnB2VdMA5v
TuAW0xogM5dqDd84K+VznElvlN7UDgOn3mpRbucbj6wUilO57RWKRD6QOnrD
JuWxaYx43w68VtqVCEZPM9dJkJ+U/h6xfCreFV+4VTf4+QKx6FFnqM0A+Yft
JlENX9alLpeH5Wi9tca2rsP97+J7wYKmUIghLqGi0vxI56wxdI4pteczOHjB
OWFLlz8pdNO6WUKntBH8TirTPkEZzYXbfRK9I2MSxGpVGmdI0PuPZe7G3Hrc
gtqZyI/Dmymx+M3T4ihsdneDP7YDmP2mFovwX2L1gJ6sMc0R++edG+VrXIYT
em9E21IU4xF42QlmuX+cDhvB1ZYNvU9ZN4hYBCtlYkNm3k9Q1Nw7C+NP6mnO
e9IFXU4RAPHw2ZMRK6B7yTMUWoWIEPnvroXC0USIt2suh038HcKegaNvfJs4
Qgjk+x/hDZ4rJNuC5hd1mOHmMf+djmLqoTw8SysnPs43tvYGkkHqZtOWV9Wo
83oz721mbtRj8Or4HIsAG1V/z8J1SeMHvAgluyUhCTC1egnrbkKcwWTpJb0b
hrruLWLkeSQN1FTeoscHTWxyoQlMfZsKs0PB7/EVo9cT41GFzVbC2bGt01DG
vcmqt88NpsPmCCMKyI9Clg+MisQwnrGURml5VdCxR3F/fiP8r72tXSua/dD6
zvKFmTdHQgLYPx+Omuea5w0bCK8Tz33hLjxmH14blnt2jmOrn3X1zlXwG40n
lLflfqXYVEuNztuvb2fx/9G0wJHKv2P7+SLMuUCnb3emNBiumBPzqUfNhgGM
1164cTd/mf2itjSAajrLIPbf3tHkvZq8mp5JuYymrMUeN/xD3SY2ZrDG+ZV6
s8Ua8jIdelo/Fv7z2ro0e+pdh7bKb44xFcrioilcBgnu19+ZtmmLl9c70VkY
wq8DPNQ8G/3DSQNgzPluTnJ1Oo0AwhvhhRXqdM1WBCEOqvOP6ZnOPBUvieGQ
iZvE2dz1Apd9g9HD1yILoS61uUKEDWrBxfe5PZf4uGNmFUw5pavpQznfzH3f
fjGRs2ZRyyIobBk1Jbou4H0haLkPE0gvC5YPLtjFDX/ZHO9zsuvd/+P+YJDE
ewfnPLE2KMFlm+41yqufZ+LOifDypHkiwWs7q3OIzouF+978qvqHU/kiKm+Y
EWclNRCo63sYxlXnVsSFM322Ie4SoUJdgIRbcuDXxN33+EeSV03+4aAPGElq
q7Rkc32ZqmdoeXbZ7KUCy0PrNtUV3XRgZImErmM0ObTtkAE4W2gErbxg96+B
+jigG/uBjW+KGhvvDYx2zhZKveBP2L/AntfXpp497FNxzRvPoUaM88kw/W/f
yO66XN2UgaDvqBBJOlYfwpqLgrshJqUEKQNPCZdJWqcWon1Wxyc4ez8QzoI2
SNiIDoaz0ATGDBpvq3VST6cd+o+68KmQyhfMdoMEPAMUyTgI/EIAbibXZ4Lx
L3okZF0ByszN9n2d5Q9Am8/rzTx1JFDFsRgJGiMCQ26h5zRswzQYIM0xAWO3
7dxddwiBd4MS5HrqQLo5e1qiCVnW1YUJmbG+xvtDGGBaHDzqivr5eHOB5VpI
APehJjPZH2f/GLPCcoX3BLaw18CJMId+ljI9ayQN3MGELgvRI+mjq0DZ59nF
4d6swSflX1vwBxlQjZXDXB5wP3tw0IbS2LHYo5UOnPFvzlMeMe78y/mr9yt9
P+hzphUdKXaXdp2sMkQTNeLZYxjn5fEEFnhxYMyx/Tp4V0fVqdyWvbbvvKMZ
PrxKh7ZWu42dPcoTpsLuvhmSwcw7ERA/qLxIYzkhJQR1zrvWw5C22sccqw6I
EVAZA+gqSnBmZF3hb8KiyubrsuQyskvFwjTujt0bDXuCx0ySfHrxPXAJXKlw
vd60Q5vzDLryuv1cfFlflYBEc9pihnjk+YZpXtwQZ6VfR0V6RWJSRj91XYs1
4E0Bq9tyuVXnWlatjKTyY8w+FO/z2YfdGVDIZ8MYzXp/x6YrBCW/gB3VtTLC
w1PTW/Xpxe64YbhBIx7S5tMzPVs3mlOmc3OjzvK3yUNTqhsMIsEmgjmHhReV
wHOzx2J9qOM5DXIA83sNl44jkrGNo9wcMocfUJEHwvc0RKeNPwg8dH4yCNdv
QLGzFsj1gqCYqt9fmg4HUsr8fsXvd1krq6CHY+kZTqk1xJDiLE6CMrk5OOOj
1GlK0BfEUKp35/atWqNo0UEchYXc4x/UcV6OxJk7I1bknXWVE8xRnewS2qi7
jQd/pMsi5FBCGQlCNjLPHq52YpNQEeuhDVhrCQm4YVzsqfmt6B+H5ZIi74CF
zOF6VsigzVekazVuOzPga0cJO95rhwP0d6pD04hk9jdKOMqZ2206v90eUCDV
C6UXGc7tpV6HvJST3n2imcQNtiNKkOU1nOVvDTIoYOQJ2cgU4lr5FJP5iq3a
o+IChljED5d/0q0KQYrx47m6K3OAwY7kuPZ6o4EMOqvIO/QaXGEYciYtKIiQ
2GBkPa9OV8EomAp85x43E/0FpbldGG4AhXSzzQ4SPm/KmUfggXAvr15ahbKx
MPtAs7f2VX9yFNR+qwt9fEAJpFtBy1bB1aCzvUl93tjMaYv2/Z3Us1zq8x93
jb/18DkA3mI9iHC9Ka+ZmN0xCRqXre3S7e4rN1MRzIFsosrY1OUNKnCNWAN+
4KqzYL/oB6+D97CsZQual2oQPdcRsORqYfC3Vt4cSYzbk6HdjNBvn3uKpSQC
3qHungfxdtvyYYDv5oty2j67w3I3a5ZFsM95kFjanxAolWANGxdmS9BPhqCB
PrOJ4qY6O4YvKxK/INyHkwsLDRIqfnMJUKuD7Pms9glt6y4NXki5Qmhh0lIe
lcJLLcZHh9FMVj/8LxWVjPAQf18wyq2WiAnjP1sug9LSWlbTHz7jqXgImR3w
5vo+J/cmSL8GLy6Br6Kn7IZ9jyodc8l550ZKAyZEDrxCNQgGtOqwgno+IrsW
S6JqhukC9TLDMHvOGStPmhAyuwFX1/FkczOK0e/fqCS2zbA5r76umX7Gvu18
Exx8Cux8WQ7p9kbyFVjfnmcHMqvoMVQW48OmbR9+VQCAmpGYHjRkm1GADU9b
VXBvnsVgDH3tEyUzVwNrgBeibp49nbcM+MR5wsrZGsqQgFti2k7cN45fC/J8
SXOZhru0i3GamNsO3qBA4qBUcBfzAjnrP8EfYSnWbTb6ZRHkMUa8W/Cwmxk7
9/+2T6z2VeL+Tq3RVkTRdZQk+UR4eW69q7YU1XrhOy3GBLDj+LFyUWFtehyy
klyaSBKTtg4VVmrL7QkX/SQBiYWPSBgI5CcHtbKYAC45qM+nPkQZyCUJWTwF
7FcIyo0z1XKB5qI6BNKLaGjb/v6WjaJJEuzYLee2Gr398AJwAQGNla9cIhi4
04Yv/tFaBTCVVNK6acHt4HC8yoPpGZrICeWkhvjHfh0irzncTNA/LpOlCu3R
k4jvPgKk14NCGtJoAEfYg7n1v+WZEdfikSyY2iOEGGAQS5aqOPfaK3rynyB7
4irPR8g+qDvJ2mDQ0FWXKqDmDUvXevfKU5KLWh8li+HISSSlDERElPHekH9O
Z7frAojUFi+25YEyanHT0bOkDhg2iLG+m8ylz2Less96Zjl/7Gvhjwd8e/dW
CAFdRBywQfbnpqxTevR9nXBO+zeM7cVWRxdtHhKx38hlOT9feQZIhkrecFYo
OxRpZk0FpzPM9cbH5uTP5ylCob0RX6wpnX9lVe1CQ/dW4uQuIPmQzoHzj9lf
h/zQ4YfaKfm9SjSiTimf6tDtQR56NEea2kFH+dOjSfK2xLs6UnT8nkMXSvoY
YHVxyW4JzbF9iRDg6p3JxtaNNCTxUIyrv1KuT9lpRG1GLL9q1FtoUdkTkNR2
8+eqYzf40UNFKN6N8mI4rBvGRfeMmRFgwF1RTe28yYPipUliq912DFdPNsaB
sTJ8+YRto3FvuDEkJEhB8lUGbv8CasptgNzPi0Pph/RnyNxbcCj6MPfIhFwg
TkKhOporquyxeOQZrEUaKpJ0kea9Jde2Ndg9GEoXHYHEZOZeiBVBt8pfoMSo
Ec/VM9JXP0MJHhu4DlCAau35xfH+60eyxlwa+IzCHBx62ajVT+7Hl8UM0cej
bcSiXuaz+ZrK5myp/29nHkw5RW/uCzhbN1bVYBS+XUP59wZzdDojYMphaPbP
vYRvkOnrgeQRzdLbt6ralNSS1jKzrmiSqh17UIra/EHJi2uR8SEoRI4oyDz6
+mvNqKJSiLFEZTWOcQtEmPW7HXM8SC4Uu7qNJUEBDeJPMa6vGmPPulqhOvej
VMGK3/We+yPBEcOfH2zbtOSufhRzI21EA7p/iYXmuEc9NekovU7lLwAZXCMW
YVfdWBNKSEqFJ+P6e0alZbuukwMpJ6zhVHcggHq/nKSneFYzRxf7On4BCZaS
HxX1kRoG1Oyxt4fzXKzRy55h+Thecv0XhnXKgccT9rcaZhjaDrbX6p4j/etm
w3RRGM6MWqINJc5LPgybw5TmXZWCzsatUFjHEOWrocx4/Q5VRobRcUgCV2AD
KbuGYkIc4CytWXfRG1GaTdDWYsz8qNrKF69/nW6cXW17Wbe4g4QUeU0AsEf+
5H78m66pK/CmZZGuMKgp7Mz/YOhn8qPgkJZFRHh05/jjODPd7O2u67UF8Lbu
m9nmI5dNdyAU4F+85QpYldxd/ZNOL3lItv+PhqXLRTm7Otlmc7XOCBbDys6D
gZHjxaUIlAdMja34NgsF74D4nKTlkpNKRLahZc4WukOCDWSi9GvDggJzBiZk
czQZFK4USk3U2p45jNuN3Aj3AEB8uCzGBMhXg5hPBlILuS3C8WRHnXDkXuRI
ICFM5iNoyee/QP2deIQAX7yO/QmHY14hJaQ+wW1ZzQVjWwodq/E8h4aQBFrl
HSeDOF7GiV+Ip4uMz19M+ycDDNzx5uNKJFxZnY6a4Wj+1pPKpoDY9CjrLU4M
Phx/64pLRnMUgJE998TyQMksl9VXYbIF+4F2StLoe9+HmN4ptYaaqq4/zwPX
hcslTVRlAXb2sUV3cOk5XsXx/DrLJxhXGtTr5d8OnRcLgFT3u3ZkA5qBAHzF
eVIGjrkeeNP24wZoE65WtSfzFnsQbqkA38i8MTjQEvSpcS7MYJEFhHvzYGnK
4w34QdW+bgiy1z2zzjbQD+uC1/bgP0dJF9Z8kmAaIdJf1tcz+96eJ+p/ML6J
JNWytyGA0WGkSnyJAwDX/JOaLUfLvEgd2L1t/Z4xjcp599PxsbkEslEUYtw6
L4cDMKORyxod0b/Ak3O2cSwUwZ73jtiJhWtJGY8+mqwZLuaNNAigB89Yce/v
dpCe9iKMQ5WXurlyv21Jsbsqde+SGqSFMI9bHhIX2YM2xYRyEE4OQGkrRVKV
zKkHNh7TeCzlzPIAt6tkKb7oHYF3BRUccAkUlkMUmYCuX+4kMHbhDLXcqW8t
XqQZ1qxEWD5aT0D8lZZQakY0md7P6p3KYJ41G9KUG+07Tyb87NyH8Z0VrYAr
5i0pjov7vTDzoj3wbDreiKan7HuB7Qwafo2XgE5rHQtpRCC9fy8IMrdN0JZq
D1HowqYrMdAjAzLoJmAmpsH6reAx2TB4E/iVpLqwPgT4HTT3skPsIui0hyoq
8YbgTS6XyWVmYkWaj5ptTMcXOL965ZmGjY2jQubDFY//5WyFyyfxusxkZ4NE
8JfhcgPB65Vu04JmValFshukfKc4DYBswrrWQh350OdUCFo2JxJqQFTY12yw
cBe4Qn3ENtUmVWOslL1EQhxgQtVOYfOfkpzQGXmCQrtgcueKpq2DBIc2pIyG
2gVphpWHbO8GSQj6+XMv/Eve2sAmGcG+8/4YqxHzrhnY22OfL5D+gxRIHvKV
msCfP01cYla/PLV1R1GpR2kdVEmffJLnjLW8Mx4XKz/Fb1i4IaiufMoAzC4e
Khxat/iznVO4wxXvuCk5MOwvFVFZe7EBkDVZgPyAlfPHA0MGcqsWDPCfk+uB
HD21EMGMKaH9/uqf0juWfetxf7Q+8fmUolpk+70XSe385HlKTf0wgJYD+K2D
H9b0tZvPfPa5JOrM71kYXqmMrhBBr+ptdS6uY5fW7EVld7xc82LIVMKIJZuy
ljBHLUnVZIgEhOg6RMN2LuABnyj7X7FeMd9ElV8PFLLIimgkV4tAJwosTMBh
XEi4FD5a3MUZ48FwQHPWMr/5169ouaN4UpWLn3FAKY8XzVrIbSb59ro+lgcH
aRW60Ypv5japg1FxjnZ9AqpWem6TB7okeUzpbwU8KatwcmxCq0O6m9jQ2miW
/szK0umaohMSHQsrdSQXabNf6VJCpaNJvUjcIN+Nuu3mpG3D6Ax8SYROm1A5
GxlYrF8cJBEdfVbzg4ON6MM7O+De22zWkNiMekDx/11EP090DIfrxA+1NvYc
J10yslhiheiYc94V5lucBN5JHhsQyW/oMS0RuInL49PKuhHNpRncVYgG7esk
TQtggEd0mdukWXy92C48AF/9h9xvC9kdWSQPNz0lAXnciPmuhV+ZMPX2U/GW
7NadrePTYl5WIjZkMUjJWN0ZjbC3g++QorxO+MCAzKziwGNkaAl01md+7lJQ
2fA9hjIuvfFxUuqjj8JxpL6Oy8a9mA27zahKxdzV0r72IaxLlYgvNrD9yp2v
nLKmLtgRkPQoPkZHhmrcHReiKHNmMXANAP8jCwmJ+He9bo7rFBrgFFNfaVxf
/EoEnqUq0CL0UjTqVFXLUjGLcuAbJAdOIhdvhkqUSzdvX1TrUdHQdJO85kD8
WffXktawxgjG5j64EvYf6slSxigSjjYCattmH3bbLHeImDkEaQeDeHBdUlMN
73cO2S7FNv0sQhAQ3O6UaI6U8sh9QfAbC1PDsZ8U76fBpxxar1jRslqvbeGu
v4f0CbmhyCuDcbW0iJ6bTCgfGpnm6HT7Zh7ihr9mEIEvZxXx91HM/5i6Sobv
6L88ef8J1d3EWp2i64uOAQR4Pj5gZbXOFLD5jW5kPup09cbP3bQDqoP3EVyL
6j7DBgf9VqfyjVXmSf0tau12eow5bfDF77d9EPY9tqxtPlhDsoQlOQCFIVGO
kg87/l/VapyglFdaGQX3xUs8fqii/9lEiHywYJ2fyym1f4fzy7EmGC4Vcqjf
xkoBM9iqLz06IFanKPgZu7yFUjWLOX8xmYJTKA3nY/0fN//rBIGTmnBCVHfX
MzAUfj/quqE2nzI1KABQDwhx7XXh6NESh+9aILlq3a8LM6sbzDZ5oraMgzTe
VjNkzVWlv7URwT2s9uUJAGuHDhvdg4QNas9IZpVL4R37qG3JBiCwfeEBqQCe
oky31Zo2H/cWUnZNxlimAYaoK/R0WgW6p5bD7XtteG5u1PPmDQlxymXYtK0O
pGIYa6KbdYwjMSeqf/fBQ71Spj1h2uRcVvZMcviUxybPiC6fUd9u4Oiub1i8
q9X5XHNZrRFcjjPkFTDtKckH40NKbVYCUszsbpP29U54/9oMrLV1P8b2+82r
/McLYEzitcC+9UqDAmJ5zGAnyt2QV3BRSGLIrLqq2TwJhTEnwVffxnnTbfKK
GJzhqciIdoQKFNXLN0Lq4BAzHNUbnqz+VaOtLoqOFotG5NvN8FzXmK4hOcQK
HXde3+gwMJv72CCA1qO9oVlg9JqQxPMhRl00UwInz5DZBfJh97rcyn8VhY7g
jATMxRXZwCprZRzKgbCLCUOEmmM2Tnvt4tiLvcVbjZ82mw8HvmzQjqP7mq5n
MC5mRwAfVglVrj/Q+U/PLxL+5kq7sYNXfM+zJ7C0wvEETQ+Fo2aZKYOKXCTJ
ZeApQ2V3IkBSE1SKcIjd1BzSOsFHMVx58Ez1UbTGkIA8J1zp+WmgOS6ZREL2
DEylgVLEyxAuLtvbEkvpHlYTq+ejro4mOV6eBXJwEcNyzM02kXRpuI86qaxG
S9ON17mF8Knv+NlOHRSLugpblNdEnvgv08KctI+cfDWwuVuiq00R1JhoxBlm
8y6zdsu2xqwAG+bJsrMawKARhd45jrUM+4zw86pU9jnijNgD7d6SPkeXEPSh
Z2pz4bF9QyjCeZgtsfuYAjxX3JO6AvGVTnZqTkHC1Psw6c/kt+5VY6FFsxSp
ieb8e/co0P9ThwdWmNo6oidVVi+qZSvff4HlUOXa3dNNlb4g9syhlVTFaqaP
rKJm9UNAGUdtAJqLNCLh4sTqg4DOGhkPPjo2AMqjTg0qrwgVDUvjChYm7X6O
kI1fUPDjfphgmLOXK3zqrdVGxxOZ62ykSETpoF+46nHDosrDrjRgk/+lqWyg
nPunfCsiVm2iVgaSgKMuU20XbEs7dpluwqWtqwu+jZXcOJxfatlH2pDOHhex
GokvihamlUCvj5Er14IfjStSTZbwikOqicWp0q+qWGmTJ3nJRKJNitlYUE7n
uq2aP0aUB3ra4YogvfgiVTvtYszwF6SB38k8zqZemzDCwnQd8sH7hPXwfHF0
6fFcfZb50C7bauyR3EFuo53LrIu0Bm/GiWDf7MbnOtjVVzXSXnAfwMZidntm
HI81XJUmZuqH/hZYfqDPDqK2ppXYAveY9+rOza9s6eEDvDQSZxf/o6y1Ix0E
1LRFcOnlZCqE36yrgPPOk9YE/PkqRfmqG4BMHPqjPlGzvjVvCtpq0Glo7q5s
iFCQHL3vvaEkfYKevGDlhr7siLD32FNGVcO4UhlXDwOD2d+48sXlzpmst50D
HPgdT6ZDPl9T3Ch5QxBnyfEAzj5LaKWCJsk6rJRg0UbJAfj5rIOhTK49Nw2O
ZSW0FS4l7zp2d0FDhn0ivPPyLm5P+YD5JA8SmB9nVwVZVVUWXq/+huSKzESb
Decp9zzDNVExbMGlBizE+z+3s7n94tAZDnfzxWxmV2rvv4//g6zIdKocidy3
r43T7+6nvCRj1RrmLymQS7JDvqMKM728OmrtXhVhPR555D+LbPZD+7ZziP+6
6W7s6hpOd7lsYDZ/weKIcxad3VFt+JwNBZWCpgEPaqYodUoH6hUpm/eN/G3V
M8x5UqJiITtzgk6etuG0F0gILSJ2G8O44O0IlhbaTUT7yg6Ua5OwUCYCe5RX
fRxOKf5LMJnEPmAqb0cgxsxVWttXPxPFPY5tWgIXw1KmjMdka+o2OC7gb/kS
Vjwl25SkCUAGuk4ZlUlgD8yrqsBWmcOfnJhqLx1jRxQl/OuZqu2VWsmJfwXo
/zh0oxIiagzL0aDj6FuTHwkfNT0vTIRMX/QQvodQfK5CCkyCD4JTTvj54no0
37glKTKhGzcExQquhYLYWgMnjHZbDlRoV6ze5QFwQjDdbLt8NUwIgNNcnsaL
0LT2s5Ux6A2avCMDjFBJMtcY2Xvvchpt4UWaFkpuTZNW5OWXlm94zdltcMjO
rG6JHkRQ6bpKKUKR53HpRyFxi1PTY7jR7sCL+xuFw0vOtv0SszUlrnJsx9Qx
iYlEoZkyCiXW+zuO0WJJCmLw7pH9g/psCjm+quzPmCqn1DGo3RGc84AMgQUa
Uf7QeUIhaOwjc/ej4VPTHNpu3gWh7o482vwbEkmhfJ1TvVV1cJdMz25qKUve
paJBPTo9XDFeNmyRQ0sH/2BiXKpTP7s+V5irKh5eXL6f0Ewk9997tljq4m5j
fT1yeAJBjF/lvegyTEn5eY1z5nC+JJEkO5fONEY2HnQt2cVhIka8+RAHdMCO
e0dzLqBKGCfZTmyJ78n8FLrHF1CjzWTunMFTGCqt49WSTy19pzun3goz5BKc
XaciRk+ef7uo5D5B3b1GPr3rxLlTTRZdtIqQ5okqEKuv8gfR7xYptM8lginC
6Ylc2VU1hLMblicxKA+U6b3AGe/NCmEuR+mesFWCw6ojUO0CfREV945Vr2oc
digKliAbA1nDQOaRNmttIlHFtYFmJg21P4wjKR3TIbqya3FfX7G3HS1Dil2+
ERLqR04qfukUbhSbV2g8CtSWF7jqEmXcNKUb61gEfi45RE1cBYz9leZ+89el
5xGgx5S8xCDVP+5XNi2Dp4hgmvI4yYS0AImd6Q2FR8bJB3pTrXXihDyHkTk1
TLiSN6ZasDyrUJvRPiw5+RbeHEBm03GqUaCKBx2KdkUdR8NRTXl8TPoAeHOx
okxEM+ut8sISoH9CAcYITQreY5e9xwkYwSp7psHRoHiChoLtzNw8huGlw4j9
nv9tnKMehCl26kF327KXTvwEasPs+xaZCFUU7CL4I5fJUW3fb4zzVSGiR7/9
aNVfhlGgKYdULDeCWoCeOOtN8UhgjLU8e4CB4WnSUYX+YUYQCaukWcqCoL/F
0hosTynF5DJB2O3KOa2tQVofauq1mDaEtyx4DqRnfaX3/mSsPEzSKu7RrEbq
cWmJJf0G3xGxZjrj9uz8ipmOB94Y8cucQY8ZzmoM/f+NORYsIyRfDRi+8AHC
MOcgddc/AKc1aQiMNOJZbhkyEFkH6TiUPuWkLo2PX/HIaw1OuW+GjhpxN/Ct
xNfIIHietyDwdQcly+9JdETxbd6oJptMWh0UDmyZ2F6aKbAf/Fccs8y38s6c
ahjenjNdOla3OtCzBMdD+u+rQE7KGsCarxIDxV/lz8idalDV5FFdXVKXxxhV
ebpOY6UZo02bzamOldvYiEks99dhIwOsXdC/Aojx+9Eitx9E3siTma97PBKp
Z3WD27/u8uWht8CMgxtn0QYa9isL463cpK5nKJA9Yf2wT+Cy0QhULuxI4iSn
Jws0ESd/NAA9mAOogRenUzpFNgzCR1JXFJairVhpJZl1AdFJ3BuG/dg3tRQg
nlmrE8pkxwRiUavuQVUsidNjcs8JckeEiHdKjy6haRrgT02Ry9NvUMbisdRa
/pXLW1/H4CekUBEj1xRxCFmigPFVdAHTfiX9rYVt24MC1ja4DSCjd2GnqrWs
dBSLZd9Nq8fWyz/VnzNcQ+QtAc23+HBrY5prg04Omhs63+THZZSyuuuYESg/
wH2uRlL46+HP7PsvBuiCQw4VY178hpB0Vre//rQ2GUwtWpeWJugGu1kGlVek
RXLAQrnSUNab+sDoUMBVxKlqJ86WdZEm913R3zZpEFzM2YTJiHt6k8YmpPIn
JrxNAeSdsfyGC4veYgOdtc90mtq2Vo+h4IINN+MbrIrBg1YJBQ9UvteghfR8
7/1L0PJ4zDsral+PC0zxDXsKmqM6+ycL9Ji+sny4bdzfP5NlpvMcFJd3NV0h
1RRiDXM4/Hy67h0iDtGLRVo1mGtdapO01qHFlivIRm9KnCfk96GoJ7PoPJi/
P5aRhp/fHm2PwFkXQgY27C59NWcWqJTlI65ftXw4fvBgjpmuZjL4aUp79ByR
F6bQTCDrGBCvo+UYMwOFWt7G/7dUAGnxCK6fNgs/tm7iB1pYU8anfyTlCedI
pnxQQOXy9kk+ea4naYXFFw6aq58+2puN9G7IffkyqMdZs54GuBEu3d2JoHrE
NoyX3meD+VnlbxxQheK5lTEAnxXvq1NYMUcyg2KVruLgsNFmDWIqDGg8NDdy
uvc/vI7e86Es4MSphxjXsdqe5CKpLkHmQqb6jAkSNLYxnJuN1tRR8qrBhiWy
w3i/kgYG9cMCu+Nv9lOjz3XDc9KaGaJykY1YF7VE46lSmrHZv3g0ac0hCxuI
8OdvEcEVFmSBb6ToFIfvMfxgSWB26XEiJ8gjdvxzupDvPiW3jA6hSePFhXqM
KbNtfxgy7McRJ01VvpHdghOft60X+K4s+ZIS22D29qEz0HFdYMxcp7uz5LBO
uqFjO9ggxQ90szj4XHy54/vr3TvglIjVppfxmMD/S0GpNudvWAzyAL8RzO9c
Q2lAKk+bHVMon802bHpDhTcyDX9NxJIzbJopLP1EovQKcM//nMO+uQ3N4iAO
YzInMR6edn3o2OuPcJv2JF6yEFXqKWy9/Qz3uVpOigEpiNRo4/J4oF0RhBpj
eksJ2x8mqvCuUyDWs/KXUTbHqaiY18edfi0NjSL7uFPBrx7bMOacf77WlXMk
3CHkb9ebnj8+F6C45FvgLsfWVJSqqhrsl8zz/BGHErRbmpnFAWVuTcAxHcZ6
83eMjTzPdfMVjvsqiSst+p22l9IiSkOte3UhhbAj9ZiEXQTxS18ljKIMHU/X
wH+AKof1rVbpTVXcU4fUlacj8qIX8lGAwNDPoyXEjVkDRZPAy128gVAbAUDE
BP30TA0AtnmA5xdh43fPcfLAL2K6Ko5i2ytzUvj20vFR18QvRfK3Sakwzcvy
RX6VVWRuQGAelfHs6wqAbN+zMSAFjrvXF5Dls4FMWCm6vGXbgsQMSRwtmntQ
nsA2x1sG+cJ4tFiKLmicB5/XKKOMEDYPZqHb3apJtrPc2R6CYmxjagHyU445
bA4jaSE9BmjDAHSZs6bFJujw46U7DiUhAGzp6VUIzzUFmxaRmF8xpJvRTcLh
TlzB2edOLFlpO6/8DunoXegVZK9baoPZU2Or3l8FDzmyVsTggJxxLlSEdqVq
VCMS+NZ9kxvzJVqOJfYxaku/uER7XNMAvRUhwX4zlPxyeFsllE2prkMuLkp0
35lSLLGuY7bixR/4M9tSW+VAHaZd6ddvTq20Klz2GbixAq8OKSr7ZKIKLnYm
/rjFgPCBMfxT6fOau7hv0+O4ZO0pS/OKBQ/reLXdkew8IRsyKfgmJa6qrl2z
l1VMGa3bHfT1uIJuW4V4UT4Znsa4DfBaDyFnEoj4aEDWvajTS4hq4pXCKjMd
umAz8SPHPPb8lNXxm+Bstpn3wmj7S7J1ovA6p2O3lgOBqct4z4NXKRMuhFA3
xAHBIDae1ndipYhbMCStzKfskcp2szJlPolBzwSGaEvMhG9/GYSOdbZa0MXq
LLJB0g8xDVNTstNMeF14TGI8fR9MfnXq55+DOcjbhX9Ck+ckMMSXMyOuMY6m
ja0sAyWzjgRjY60Rdf5AcR1m2gijBli54pAhcoSTlVsxsMl8ZJfG1beKERYH
pOJ0R1F34HCVA8BPQ4E47H9zQw+xzP/996MXhR4DxL/CLaxgyK/yo2DT3956
30xrSN9Fm0//o4VGy4KijjCAqMZYJOg2pFHrODqnoefBkJR9YlqXMbULenaT
wKAMcc+NZDOaaty+CK1NGvGVNvrgLxOimwsV3yqc4/BsZND4ibxAIpD1VrlQ
pkrlAacSnopadqHucghiwjh+D3m5bhU4UAfyhu5YwLH7iktWOA/eRafVRgak
Fb5IwjfCY85rbV9hv+oCdz3GpT6wQKr0otY54fWsXFuVsmZpLlUvnQxe0rij
jRgaYRytk/sVCasyhvWD+ZJNllycckdTdZsl0i+swRi2Z0J1LDlQFc99+qBp
FTbKplLChF3M3I5LwZJkaOrDPZ4jxuGRwPHOsZjX1INeKir3vEyqoBVXogi3
x/eOLdNPF2IOGQnlHzxzDKR40Fd0xTAK+CK7Id7zEIV8NDlyOPDoYLDnG8tT
hX50U8gXgEZ7kFXxtH8U5l91pse29PSPSe0fVL51Pz0BjmQ62tqdGbOpaaiI
QaSI3V8EfwVKwl1UObp2skQLv1yhlGfcLvm4jKG6s0Ao9m6KrDs+KFiFvgBz
yQ/Ms3LRxqhQkKvospj1Bn8NIsi8ljuwMdaGGkAhlPUk+2b6RUcJOKfMgu2s
bpPucS9qENorzAt4wLaCsR4sV27/ZFoUNN7SdH+D/fVeFLvJpP81nQez265u
gXdVRIgzPHfFasMdDQ0Uwgm91Mw2wLdc2SY4Ive8jsITQzJXtAKIlYupnrDn
hp0WR6cFXlAsp0lgV1eyPtGtwWalMdFnboKg5YKZn46PxGuTTXhwv6rTImjy
v5AkWIJ8gmbZCsX75nRxd9cz9U+1JDenIDahzeH0tmruESSTb9kQAhSw8mg/
0uudRORiGRvK2GgfMxNM+GzA7tlAsuym3AifPbFDKbHNnwtIoJVCUtorr2PB
CnDtj17yQwLqDW/GokzntNZwpjze/8D9ke3CxExOu1A+D0U2AbXp1fACEX3g
5NrSGnph/JIIo2Wt7pVn0Y/AAUfTcey0vR9IX3fBaYaIwcu70gQ2IZMjPqej
6wZlILGeQwz1psN+U1OjCiTXqwmWjMfffRNJB93jxkY0Q9rCojY8sG0zkui4
ZShgO+OjXLlUXXOiHrOdDyKS1/yThQesjaiaQyOvOYx5If8TS/L2E5BF2bN2
XaRVJj+6R8QIljv8wG6sbQRzsKYq/cB1zLor3x802QiCgtCoLDvNM9T/0cqg
OBPpGYk4JAA4jRUFK4zU7b1cTN7dypAg8eByeGKPHbsWFxRLT8nP9gjFK5HX
YZoi5tmggyN42zaXdZsxTypVXjYa5pQqQ1+aXNjqagVWZu5DSC/LXfIcPVya
m35+obwl9853T1zeVBfbGm/wIRlEA+NiuzuD5Iu3WUPW9+eJfI0+btCyPMMG
vFZXBzlzv1gxueRe4hpekxdAwtBgAxAdhRSC/nx7nIjjHxJjt9p6YTi+U3CO
sWaFhrzBrcFbWInfHZhxSYPzqw5XX0e8ZhWjyWT7nrSwoE/3oiZxqQnETCAE
6HlVugNP8TNMLBUmuo60ZL0LPUqpG4JP959O/JM6Zcpi4wt0n33BdQIDTgDl
kV14BRgHLtK7I3UT7pNQ/V8kN5oQmPecfJHvxk3xzDftcMHtLm00uTA9kPLA
9fVIRCEPDkiEdUaSfgIOGi/Kb5fyLImYCqqyx7Dq1+xBGVA76kiQP+FoobBp
Ve1A3TDzWTho9JkzKRUuzwMoVyxeQ/IYj38fzrtwJxO0o4zAHLTqf3a+oZir
9j4/gg2rVaVLUjlpzouPbJCoL4QJ8j3me7+OwQeoCMnpgmg6ZQfSb+7g+RPI
gBuAKvewyJv/EmuSGGIVuM/dFCTT4lynfFkQfRDpOKaz5ETdMG3kLl4ymsOU
R2o5A0Wl3/9Jr+oA5GFONQib3L1FbcFTBbkem99zFrUG7eEgN6QLDMU8mqow
mInRq2dua5LviADV7K/hg/hjl+245RCMyW75u/T9HD4FzLVXmg1j/mWPHWbR
Ct4LmH2iO6V8CQKAvktKdBMiTRX2Czn1QB8pFjzt/iotznNbt1xAp75WwCpW
HKerOHpdpobmfXSbh4Cbo4aD92mq7VQzKzkDBmzWSMBcpC7riUbzzSUg20cj
9rIWs6Gg5TefnkMefmDFldpUZrvV30XoqxmtuG1adf+9RCqzG4AadB0izByF
aQ84xbWL8rEnigPqgB1u78j2jhKvS16/FKE3LYXiFHtYwAvL9dr5hwFi5Aeo
UpIPpKvPG/mRg6wcnJoTn7dEHT+dJeSAZu/XYVd0hXAqdnzceivNmCdz1lNl
ma8RXHZjk3W77oC6pvbV1GrUTYHNExu3wuO31q2Jj/qiZv1PmSFuuJM/gISh
dMNaNNw5MTJRpCacpG+nK7QGvVVBnEtz/X7usr43ozxZMGK4oazHlYeGbnBI
7lDAL0GbXyUb3FAXOcbjEf2v71acruQgnJrcpEPY0uB0oBfdkSVuWvLC+gq/
yS13tMYHcSd3W/3NzC7QNbCWHE6U4LoR0bfOfjYcs6hMfuqx0DLv90BA7VbN
vbuSPZ5Cfeprm6QD2wfNf8WDafW3bxottuue6GgbCP9upK+yIY/f1igloVtJ
U+USwf+yYNzCre9y4zo1clouXiswLkzW7n1M4Atzejxf8qqbk0D4H+rh7WuN
X6KelJ2l5ZjWKEP1uwbbKefLSSQzkb0nRjOxJbDcGt+oIGnfP0oOrhgyxpwE
8HRpkdvJ47pOWIwIk4YDPnSOCHjcqHpSUq2gecTcApW4FkXeh6T83t4GK9QL
jGITZ4bL9J/rAHAy+//pdYyzqGXj382dFYEWcV6z5flqdmMIzQPY6Ip49Nx0
Bw0yk0yWG+GDzQcMgtEpJWS02vHk6jQ0TwtZZE9Y2XFOGHxTaTpABIYD55EZ
/8isz5O+V2vK1duCoq3OYCsgR8JNcB5Ei3oaWTdWCu5/EPBXo2EiNInrvC+i
4HwtEDvM+3XRedS4GaKPdueIrWFBqBx6N/ubkz0dpEceF/sB7ntFT70sja82
hlUSGVGIaiPeFyK1344WhSHuxHDghfQ0sRXYLRlB4xrm7p2igLm2lmONNzgh
eMszDGOv+I/oukKngLeeaKkMCatQfIYxYvTPdA1Y8lTjUk2rdMUE8NIimEzZ
w8YsdbOsO+WqRDYC8nivbVXjyx2vShU5JKo/wXfzkyNfUHtQP4ic1oQWsVjS
6jKfsBB1fkjCi6WZJbeWnpOWDLaAiwKduIl1pVdiufj4FSdbnjLKAnoi3WMb
ZI6MdVMvaC6lCoBuSFJwMLm7h2pbSBsEtx0BHF0bUtIDI/mNSzRvBQT39+an
hg/xXoPGJ3qGp9h1PBhA8gh35hOXreinD4+fybNeD0YKNPghnL2EDWzJe/1z
77L9xRdBzoW5LNqQ3zPqIUE1PHvWZS6EyLD6WS90FtaRM/pc5hhnLqqVFy8Q
jRO3gQyLBqSMFMhmvOdwyi+VvEhJYjoeF2GeOqW7wPDvqpTG5csjeohdhpXE
ZTcKaC0C7I59YXDn2Gz2V9iUp96S3y1ZKhfwRy0o8D2A4iuMah79uxHwnxKK
BWrQm4D9eRT/hJgDLm2majDiP+ltIWcuOMjx4NoTtVV+qGzrtr0zN69bD3V4
xgjSKMUpJRYxq+9vMGC1lkxqXJRtorC+YypvTWsvPkQAqpKPLGfXFLVrgQ3i
vWaOcF3hyWqOIopLbvOcdN+7zqJRt8qOQdlj4dcEBibe2RbWylVIis04Zv8K
AmQW8FJHaMvvjMSCKKJ5nazlSOyVUVdRMh/UxhYERzkU5067rUgKZdA/htRQ
JPulZxdNeah4AUn8wKG7wnkP3Ll5ckx38ZoKDPDJ8C9ns3iCI/Il8MyD5CpC
BB740JoMPhUvzu4+at4/R4waIDi4Egd014AF3WCPVlMQYGu64QH6cJoeHtIm
ISPzzbCt2MCgf2ucydh+1lo5j4QfOVfl2ubOCZZPN9iqgYCIcR6/KGr5GXrg
bwrLNPfAG+033wG1g6yNy6DuH4e+FYNZ5BxqAyOGjpD73Ft67q5GRy4GjZsm
JxI+VstKljLiciDEPEsggQBWoHXfCUCAa9IQKm2iHpMP2QNSpHKDSDxJ1nRL
yppxCbletgxEa6+CZFS2av5KK1SDb9hDhL1b83YyvKuMK0dtyzToe3sI9p1G
LAfO+SnDmG7w75CLBHvw7s2klMV5kf0qv04u0kzG8llc/sOj3A60oupJQ9OK
hoXAasMZW7KOMw+hb6VaGev6DnnxM7KOE7Ah1ZOwI9qnz4OtSZgOrqaXbIC6
ahhQB+bB7n4SJICKN/t2ycgp9YufKos/4Kvbd4wGwH0UJXu54p+0yZoU+hTM
sbPIvAE7hQ3Kv4utN50C+/zgZpPudWBvQb63BujMP0342KILDSjiikKflpxJ
hlmF4xotbUezWzavL+2P8LoBvwDraDH6SvKA4Vxb/M5A5OzGMEfCkprwb+vf
rF0CH2UGe9v6NfQYyujfCnBLr++mn+JTkBkhyQ+nJCti3tBOHUrZgBMs0EZ1
/e7+gtwmeVwy38nbIuw9HImUiUMWYn2C03ve5g9jI5nYWW5HrEa6JsFhi0GH
pxI/kRK5Wn+COc+DekN7HNR1q73pr0h9DSDqW82rwqEQ+hoagHamQUnLBrPI
fpuWOcuvxiJhWBkHC4Z44O10UnPPRSwCIwr/aFtBrZGDPgVP57OY99mwXcFU
iOwK2fKweFIu6jmqARKaaVBBK984eULtiVwKIZuZBbxEL8zzjDmgnRy+lVDr
7Rz2N2XbhLfIE+SBr+DdI+VGfoYhXMr7GDMrGwy7pdnMgpO4UPrQ6FFECute
TzduKsAUNY3E8sMPx7Yt//G1s8Q0CWgYTaHkbsVOekOBBOTUSaVVYVouSIx7
VOLHGE7qMyzm4eo/+yyvWpzwXgX3jlzD/+BBHf3lpRC0JL4RmNoeTYjpE9Aa
GGygtyARnq44JpF0Ld6sDcSwx63q2yO9+uZzkag9q3W0sMACwTmsPhUDTfUG
EPlD7U8lYofc+X/tX7fHh8fbsrmDMghxlnOF8GUpPnfHwkzmzLgILxyB8vll
HLgttiz1R1x7C7v8kaGALY28UCQ+wY9CnhCoSXsetJiepHpSg1PMEtpYaYn+
Nj5ozH45c8FcH1v3unuW7yjMbQhVZvByqYAhI/Ow4xiu/Yq9YoStAUXY+BZ0
zUdjUrO8iOIthKUiYMS8ozpqVasuorxwyWH+y8X4We0JHKr+Ga1Kv3baK+R5
vsQw9WyZ2xyh5fzb8nJWHf9RyFduSwkvvEn812H49sCWSptTXVCsfQec3olw
zV3Kke3PY7LUx1UaXcr7Q6egljHwU8vrgqgySgNATPxztMBYJ0SYMdXivu99
5k0cPKYC7KVuioJE7b6B3QTFwxQkVfQMKxBQmC+QcxG116XqQjIJp+Z6O5BW
R6atd7KTZ5PMjaw1c+aS54uErnPzLecB7nJoqV3ZMfB1wKb7hRl8XNZa7lxA
BuHtUwrFuUBcfbfxE6fxnXkSbGS1O2wuP9Rj0ge6VKQdHuEll8q5CLMoAIwV
SGDyz92RcxxxhhiTLsXakM09e4TYQtdFh5p59GHmkXmyQ7JXylGP3cv/K6k/
lmeoEKWhfRcPlWBSXfbUyOnhTm7qM4wxtPOIPAe/J7KQ69cz/JJuuxEjTvTe
4ODzmJfNDbFL2XEOWrwV5Gkce7hS7dA2KL0BommjAje2fMNlVzyBgHVh/MZU
+Q2oAopgyrecAOHc/guzjn02VpFr6/PK+tdhfrrVANhyF3If8vu2MQKYVA+2
FaQHSQgP0N4zmneYMq74FZgWX4UlsiPta192dJ/Hp3Peab4/bMQnchtwNlPP
3i7/1u2gudT0jdF72LPrFYYcvTOuBVLlo7F68m5kP5YaQwXbQtW+2YCTcFKK
n1WlSvvhHZuWqFHkgcSTic0LjxEHRqUEITq0ZfZXPlt/6uTYhyjllMC00R13
5luHG2reqgMaDWV2+JW2v/O6e1p8EyAy5aCgVyg2ntzY1A64Q+JzJZSCjZv2
QS7Qsc/9iprJO0Lz4I7M27btLVhuA2rquyWef+R83K80/1s+uLHrjuGBzGk+
T0J8XY5MnKi7yko+L2LPlW8fQ92rJgx8Q666hWW3VtM5JZGg3srR13LiC1IN
M/gqcTUAroegZ0EV8hXwyqwutxIlCymvvR8c4tQoiNSX0MeJ3jEcm27M8ILF
490qll0Zq3NdTTiOY6eI1YGXsIF6u2Jh5t+JY60LCdjXPW0chbvpSGm6CUWS
2NDy+agpzczdHFzvKKNpxXuG7If+1FW7hz/HOLjLKVdmSLJ6ciwpxe/k+Hgy
Bxyp2zzCZKzhvR37HvL0mVZW8LlYErMOkmIVFxyIUIkblV/Zd7bbGWPQzpug
Z7xRysDr824O9HBKeNrnHNQSc62HAqe1Apne0GDhcvr59zcEUsQ5wSPIva1Q
jsf6KYRoiUrwcpdH+/ciL6RRZSZE+g0hDSCVNsMrWWXWvi4yoXFoUE2yH5Vc
Cdo8q8UVaCKOxVvATwcAuidgy0gWb+yBb/KzUyPiwWMTYD1kCTFNBSA4AIF6
dcRvW7oq9O6g9lY5/AzvI5NUDMgFJcuuk74YRMOu4gCHqXfgYHa3Vcg0/0KM
QYzFvz80LnMJsIlM+9btnT7laUA5P97tPnOmqi2pn90qI8/asC909ZqC7pmV
zY3sd28j40myn6DaJDtVnwZMGagEcPK1h4fUkZ9wJHWKWyHQHaLKqJbNk6ng
+6BYI0YnNPbTd/kIWF/Te3vtycTahX9b6aLbYKsROXRmGvGNU9JtwhNgplOR
HwraJ52eME4UBL5M2SRWKc19x6xS7DMyM9DEsU9uC5ndzEo4wKUfkuEsduKA
BBrc7iuIgOKJOFejMFRczz9ILNA1JY1AVpoFYeqVKrTz9FVStWgOPh8Xg4L4
ggFXuo7G6nc5twWEUv/YTHl8555jhaM0zf/uycVeMoSNT8nJZ3mCnvpakUXZ
jD6zDc4+Lf5LMXR/dRtdr6wCLGJmydtf3i/I5UfyfwddDjRsq5E6f+dobMt/
KLWQf6zMDCXi3tX95yo2BVEUFXIzk84IENP1HM+XMzXlSqlWPYABZXgSMoim
r53UAIrGmbueSaOt3Vtx2S+IlCPhSmm7a/ffCId0QZNOV38FT3KnMZlcf0HC
wP+0sGE17I5wbQIajxUny6CPMxQLuGvwKJS/xZoDE/F44rd6VS1WYAoHzGiM
ygsuvedVAxTIdlO9isnBSBKO4p8w3M4/FmjDpOSeus1+PW5JdYwzDxlIotZD
llSL27zBCDQGH9/onnUXN+BDLz+HsgSdo9NrjBbbJhmtXpKHgZoxQEtD2a6j
i+CdJ0xJkOUpLzG2+5LAk/uMGVUcd0iMkIbwQPxUWvC1DdM++QiWJYUTLy69
J5xIqSGoIT52qigIMk++7hJ838IgeulNusia8cHmkzPDWcwzKySnUIKIG2ep
5ysBp1R3FOocUXAhYuF3GCPRMWYII/wHepZPAp846YBjfjP1z/mIA05sPzCL
UmxAErZnzHBSiWJkFyDI3e9LDK+lOzVpLY4X8bCcgmv7eA3msn0kibbw3Vf3
b5LfL2k9UaxcwnhcqhkQjH+b5QPifcwURKtiRRH3ik+3SyZ3211Qx2sCGPdI
vs2bOKIgFDrHkw5wIcjjZ0P0z+WscexV2lvjE40RzLu+tKxI4/KtZ2i0C0ou
1z/neETwIzvlDobLYb04KTx4vXdlhk7qunAPblUg8Tbf9KxQdAVlE3tKAIS+
EtEH1brRxFpniIm/34c2rPJ7YMDJAU3nB7sFoNNG8caiKrAM7Ux98jF5224x
uypNXBg9DrwfJyEUs7RcJou9YBZf8AdkfAoPxb1D1nkLRVinXoDPPULCArwQ
zHjE79bbXJ9+ZJOjZgnhKfs8IZGHWz7cnljkTLk61JeWOoxMCD1HAzA5qBT6
vJ2AKb9++HTqO/vYhb4IE3VDmsBjph8RrzMqyiTlpq9OjFmFFXk3yLbC/25z
xGjYwa40/boJM4gJKM8DXBBp3RYCadTkFMyC4ZL4QJolcKK1JaRIZpmYHkBl
a7yJT2GnfmCpWmAyJPsLdvt524Pj57nh76C0+0ug2oldBIAQKzF/fe7cuhI1
qZv4E0MeQSXo1difbumNtULo90ku9jzrMhb+PU/uiYFTHhBtmbfwaklEBvQL
N014IuqekshpRXvT3+w82PLA7DgZDgGZfCXOHbEWMZeRWrUVd24EU7CiSFQj
mXioKF8a3r8T9vYSP+nZxPiBpy7kq4TeqjDmMdbBUkZoUXUanYntzy5KEq7H
fkD9d0w3Uj+Dc08wMHOVFuZN+uUgFD34+8Sq4z3NMxKwxTy7YHTTeCFdnad5
0mcOisZDvWZH6JaGSPE429HIvhf6KNTW9kdvMQW+Nf+nWKxN7s+AYXvx8Gnm
ZhjTrvbA+DoJvbOJ8ckRBXFOW4Sm5ujDh/Mz3FKw4+Cq6aAyucoHXNit0LgA
f5LZ6KGStZsREuiyWjT5yD711BEkkS0wHXXO6u0Benl0WxTWfwQLe5WzAfnb
HzQWhxbLxmtpmzWwFgIQq0y9mMOv0Fg/PGrH1fp6NatB2hYYDRCtu9HwKCk0
/JphwPzLPkSLqmYDj2HjWhjqnA4gSuIFTZr5DPXRUlitAmn/KSWvUCGznn8U
SIpmaIIreQ8iVpqDgTwIC72yP6Py0G58W+tKZe5YqvxZzY3ptbAIO9o2xuTa
8Aaew7wHQoJn10yCrpr0+Ja2O0SJF+zfJDdzlx/nWW7Kc9yUeNET+To3jA+d
iE0Vh25TNuT6D+ssvRkYwNbcwDaD1KdIPvPfDv1u0X72thrBnFPWGkmDpd1y
48ctwJLk96celZtQIV8dV+y74+QP/I3NYfyhgWAM7KCKdrIzwY0uh+AcIJLb
Fb+P3ssDDF2YA9UyL8OLJjf0c2JwLSDSZFEjJJK0qLPRM6wMMWCSZ1rGgh7r
hlZzAWTKfCSm9yLteXHfAPlxXPdPGvZxl2BOMKp5ARP1iGwjxnmIeJPAYkpx
QoT/UuKOQ6bZb5PaCcrj+uVo2wTWlAc/EvafZ3Y9KEI5iw203cJrsUHT8Mx0
K7M8hTH6PA3HCQeUDFps1BrqH49F11nSoGuAu9Xxpn5ZJw5Eq6zY3uv5HWL3
YqzNCyaxQ4QB5Qe62BkdXqGWYiZ5rzpU5t47ApnvWEcl0p8o5DMlQXNS9raz
NzMOLOm8EJ4xC1wMTsNlgEDOyJZLTJrWVI/ltwHsaqbsj2UXATSbWXbxUE66
K58IHeV/Kuwxcr94IYMtqwCxfswGN6q27FGmnrZ1nRfjOhsF/pd8RKP5ERiE
l7hWl+m3QO4o20C/cFazfGlk1eRZmGHW627TxFSvrPISTk30JucOOESKCY8X
6tKsTWQPg4NZ+uk8FX80TheMzISMyPLFWsJg7zNOX9HNnUD06PFI6+tBJ/Qg
+3hyTIAzadzAtkUQjq/BcyANq2wykn6Pfy8WCS9gvAj59W3NsjoS+CHBRiy3
8YZa5h3dutE0EAjw8k0fiSiMI31rn9S7DhAFFano3vkDoJanysj7svhGqvcP
Vm0z/KFJUfvLI7RqOEW5XQ5HMRRdJrFfjR5/gfxo7RYFCPYlR+gUqYHLsvuC
UBYme67o296ZwCY9Himm53jS1ptdggERFp9INyEvkM+IYmrqfE7vQI4Bsc7Y
Q6WW2x+rDjmbFZdCVBrFZCRMIl30xXB9qHl3zfpBjPwkWb4LYCKSDJ9EWg9B
hkWDTGWNRRgpeGWhElweROe+rRr00JM5FG99jc1zIs9mxa1NVuB/fn5iSGu1
l30pvNyo5Fr+vRqO0H/RI/A8T2IamEPfm0FlS+2BowvvNSdh8xArlBNUKFW8
Ki7bHlp/+Dj7PQQBJMc3OYtPzfDpp03cO0/2v/e6QhT3udsZ9dUdUikaK1jV
r3n5/nWwkzz/6NiZGudRN01nNvv/HM/oyalpohPrFZRCmrvU0LkXK2Cs2y/U
t3bOioHjjGMArLo4wRcVaZQZodFAlmu69Uq6R5i/27BJWuLMAVBBuVbgCxeu
4eF9HLg5xJqlK2mYf9id1HdwsUocWR9ViWH4tvj0rKLq47aJwIv8+RnNrTfv
BZY033wPV6QGqUoMFEK2Yw0wiArn3QkY5RnBumyiQcLb8BLkh+jdlzaYbc2H
gDl2x/gF6k792xegF+Mqq1HnsPI7/qKCy15VVAYJR/vZuJi2eNGzNkO1N9+m
iWbJFg/yBlKkJk9CyTXVF1ONcconicldAdnZXkC1KwP/5XQxONOki3hFeOld
MeAZ3aRCSOOaFK+I8eXjnMigngsKpaU2IpI7YE8ZguNlTw6iHjHfq7Sf7piy
/ZhI15SNq7YUQFIKbK+wlaF1K1b4v5I6++m+8N2rmrSKcOQijnx33vX/HIUx
RD/OiNrhLHByzDSKQv2BMed18INl86YVwHLigxvcjp/+Zuht6QnrCQnKI7uP
HWm6yOhyU2mXhKfZt0SfmtfDoup8L4MFijaemA5HxMSu0A8oeacalTPd3CJq
tZxGHftYeBeYnILpY46ag4yVPXUhuxxfLwt7a29gl2uNzqJqw2CJgWH3heCc
r4u2ZJoquOIoB3ZptGRXpJbEaIAjaNXDJDA9GfsJnsGy3Zpls/CKpLTOdQ9F
Yp+VyY93eH4IFxnnZnkmQnokKTBu0yM35JPbwm6n7QwyyvxwP8TItD9C/fXT
nEqBycnEqs0WtbggHKdYMefq7CPCPbq891P+V1hSsm85cxMdjP3mwV5yPdls
QHtseP3xeCOCGaG2ubjcipBioNWiajNYHMkZyhMSMpqgs/nboSakRk2r0Yqx
RMP5qJcq50Bv5dV7fxLJve1GVRK/ITAIGiz8C2ez112Ly9E90UEBjDsGjBJG
oP5xybXLed6zA8POidaKgugKBefZMUBS1IvvbQnMC44QjcTtiVoiwXcaq+RI
s4wJJVNBtXnUPB9jwZTADxBF6EamZII19m5ovn2a8GnLT4aTD97s6eyX3YlV
8bTQlh/6olGns+V6EBOCjqzzNKaiIU5uuMzpgE08UqgFbHTsBdUACqvt32Qz
NlodIpfuC4MBCalOD1GKcHJoAeusf0SylT/pcWeMsxq5W2/82NPaaRwsMJ4R
O5is0cB0Ag1iAjEHqm+NZDw/BvsOMlXJkHIJsX5yM9ohmY0NAzEQ+7d9WAfT
XXMtoACJ6L3Xy5rDUQIyVGI6rdBGJYq6zS0egWBQhjtU/V0JlBADyL2wsMHu
1fwGVNJAtvecK2+dsETCL6kRijeLfzn+3MYUcDj7b+un0hCNyBzjShGzxyex
gzwYBBdtN4P3LWSr/zUEyVUnYMecAeWkvlc3A4m8U8/6pC1XBMo3W82hPJYN
cWV3SfVXtWg2sE+D7uyoOfOA+rqDcuM04aNFaIp2b6HMV+NSHFoaS2iWmSW1
1GO3TuKNHnz8jHY4V6h0th9gt61Fksx31UMnps/iFiz+jhA5zoun790Ku1SK
2vyFwgx4xlSOTxuKzx1W9MRZsag/Fu/Q55HKHDkbDdaNZtSTcm6dxytbfNV2
5xKYDtmwGehorl5VyOvUWu2c8jW0q5oQ1rfwK1rTSXOndsPJNWJDBYWcdFdj
ssCmzXyWmPt1bIsDV/Dgf3g61HxrxTx9+7P1ypq0WQOJ9vAIautzy4m/z1x4
r2kNNSS/2QoV2ybyaMdMnMKbDVoVmuBOmN3iKX3EXoWLBny9RQI283ByOTh0
ilJKSZaW0Nbf09200jqcCf6cnIcuRJ5bqcu/MuUtQnxuTqLHBnvnIrWeabnW
m9O214lZha53ZZdtubz5IjuMgB26ZbcLdDRob4lqMBFZQqMyO+ioYtTK7rnz
Xn8TwYjKbDwAbTHC47QHar9KMDk7ofKkPQsSnW0IQrmST3OuDaC3u1T/Qqo5
0sp2U4vnyxLIDa4/GhK9ffCBVDynpMy+qAA3tAY58XoCMWAeV2765eNvisw3
xr4YTGBJDhOGRtqx5SzF7m4rH8Y5N/YLlBqnkM/W3Ybpv0LrSnZuV0jpr4hy
POcbo/W1/UdGl2wW/c30YYmduZpNq1x74NwVPaBAk2tpKBx9G8qhZK25MCyb
ShnhmDDwsrQDKYBFmSj5raNEUJrKvH8j5l9tWkGNH8LnucJWbTUTkA60rFYb
P4L4/+W4k3whm9ylA4E121T8ieDzn1FQvQUjflWZMmJOAMy4ZHRxjVaOUykP
DZbniqGVcMnhNnjA68ZNEbhQfypSFErt8iK5prlXpgfpAWwyOP3srofOqqo2
waHMjZUQP1ejBynVNTzxRibSttLDhySE9ZG9fHCZTUKC8sx6cZt9+pp9LaLt
gOAMTt4YN06qmbGgB+a0wuVhg0CVYxQv97kCi7MABT0lWiCXp3iOV8Yow778
g7XaPg1XBvZ2muyt0EobWmrHhjXEE6M3OLdPXF6hF8lTXcUiIiVRwpFvKf2I
pnmqIr+DVuqq7eW6gudJYdBUeOfIrNZVKNuLX+v5UYiVi2QLiNhLtKlA8psB
6/ffB1Vz871/76s/VCg/h1o4e5z+AT6duP7Hlh/vfMTAb+7ZLg6+SPnAqWlJ
1hyXliGb7G1Cb4dAzJLbxELFaEoNLgh2KZQwdeHC+NHMwTsDa85deWtRGPEw
zarsVYU536irnIw4looGkiZPXh4tvZbG5ua8gCfo1QlcN7HR3mg+7ghxAyf4
RdDK9X0MMV8dOMq4qfkLlfuq5971VYbwyCxrT6YbzTsmCu8HqkDQ01R7DQSc
0wvFTtlQtzb6yr5bxb9tElpVAzx33H7gZJGEa4Z8yHVN+Zda/Pc0hu/o4sKI
NSBdERTrw3Y1/ovX6qwfXNhflHqSt4lszKw42SRcGxLXKkTsZBw8YUbK0rmu
X43DPTncAL94vePQrECCv+IaSBhPWifAv8E+3BsK6ahTwPjVE3mWaKwIewgd
4OmgydeNQi0vaVz76DsiC4P0uAZWUqVNR6DEL2+qK+fPNzP7sX1mkN9JTPrS
7Jbmz+1t8Hc4+p0p8X6Jf5VIfmj8bV9QzfxQttFigeI3gEwHiyx6iNf8mXsK
nd/sFn23AcIwhhHd3FOvaj3H4Q0N3jE0pkXn5hxGkk2/FdX2Nm1tUMhwHXcY
C3CWb1a2x3bCb7ODs+gWIhY9mLX2SoXOM+fuIl3IOp1s1KXszVUfflHrIF4z
igBURLJ4p5Viv2p9UkJSy4OgA49dvMfz8cAX7nAyitDqkIWjmtVPn+Rp1dDh
8K3z+qz3J7SO3+IcF+QI8z0UDaLDRguXDHfG1ULaUNF7g7/leOGYW5X6/YxC
Qc6c3r/TCzSldV8Mwav0hArLwbDW+QWjn4o3hODWNM6cH/79zTTHal5XFJF7
JTlltAa04eQvWVomvbRqgMQqMHhOufeIXvON875gwjMWSCBjpXXtoUCAm7du
L/9giENWr2BV03A4NabkSYRMBuqcABsZifEPfsZbF4ZpYlkqVej+b4TMITja
ANwf0mQQ+ywMILTWC90VZ2pXo3DRQbN/2qc8Jzw69WdAbdPn/zEVu0qFx7Pp
nq5SWIAGxP3aewOY94ejN8/dlZS8yb8JR4glq1pJAkWTsR5AteCXUOxaM6Wf
NaAgpB2bFB+uhth11r5VPaR3UkMVCfww9m6d3FaZki4RRdj7Rc9pkGzScYkG
57tbAP3Fd/lFg05XrxChw69JquJKjd0XKsvESvLtspYb3QH4yqjvppT/hwgk
R9gtu43P2OuZgYYtJILj21hxOJKVlgxD/ZKoIT0i/g5OiCe8wrfdLfLof/PR
zMgseoV7h2f4NgOLfNKD1Cd2Cf29EnDYAMtefJuYtU7w88Ho/CmsN/kB1SUv
EDq+nFXhf3cxSwA38Dfe3ZZtz/2v3tgIibZYXrabkdtz4fF9Qp9IT7FmNy8h
QtRLHVNiP6RfzLRqj4ZP4u8Uuz4y3r0fkKeoleejvNphuLNk9imslNxMkF20
KhboKkIFyefRiSdvJ4yQaCoiiLBGOTEZCJGibNkuntDzWbwMzC2RbvJA4VcN
sLmLISdPrNmHahBtFnF8DV4HOl0V10gQ5arRiZD76WGt7p6EWrjRC1+k9bUg
0pGlf6bOmwcgrDx4aR1k5Xy4xQz9hxeB8OiIWSORTLFfryR0WhdvBYCkbVAl
r31xpAO6/Jwyk8eE0WYe6Za1oUpl8fk0oYyyepvKVwXJdphTH987JV35FE1h
sQDgrk7AFAmQzfYRWMJrGiSFUy1KjuhFukWdDFTI9QX9m9PFnIcL82KbpVxJ
Lm6wqfmk+O4m7vBbajiFdfVYPn1UuLEbu1Nr7EhkrrkrEtQOh1TChnbmzXAJ
DKqT18jCSjWo/K1Y0qHZrQDpXI2vmpg/OGN7advF+RAgOXkX30uzP4xrA800
pD/6JcULJtoZsdq4IznNW2rSnKvY0aaNQt1MzQPZh3F/xl+C+zSLas7kHnOo
WOAgrnSmd7egCO4gml4v3fBNGeTrJU4B5hySkus1T6ZPc/Hpq2ORC5e86Ruq
3GMBdfzcirVAkw2MFU7eJ78TVjCxu/E+nmi+tM/aWSTxkglUC1deeKIqH9gy
fO2Kj658zegYDXEjhdI1xCc0u2vaDBsWOD9BZdmxdvFAhtMrKcLbV3MjMmS3
ZGgkh9WhANKb2XDnqBaYzN56x3QnZP2BylyvuDYBXBl8y3EiAPu3FPx2WGjR
XwCg+QryEIwSvxQwDsOBT/LcbOrn6Ht90BxNNFsZBiU71CG2B8UHz6u1MEI1
TJuSbbnDpPxG5mEttxGtTSI6ENRSKceRDF7LJpRQ41dsSMLfJitfYapJctfQ
/jcOgfAhVN2Pu3/t7C6GT+rN1/XMdZxD0Kw7/mBcE5FMehDRQ7b1P+O3X6Mt
rfNUl/M+I+Scc/LDGWrxx/K4XTH0leXGQJ1+WQ1EeFqqbY27obOh5aCrTpol
J88iDO2C2lbcBhNN0dHyL935kuOZhyAip5BjbP39nzMT475prIROoJBuKQTZ
EerE59Dh4DZuFVuP3Em1p0PZ1pTPB/AJCka7e0KZREMyELPSSv5KQcxGM6YR
qRnw1+mnzZnodpfq9VjDRlIpSDBD+M3nBnkNt5lX4aPr+21yWUiA2JWV/M3a
0657cu5s2jnBorVKq5yGImSY/CW1pXf2ixEYSd13fuiCpDFdYUOInmAhXDbs
MghHuX0z+yR+1640xUBs+whtTNjU/e/GcCK1FYmLZgW87yY4qjsrP1FY4Y1o
ySrbdzSDve5Ym/66GULv25Qvuby1HoU6mfqsbwHUiR/NdgbfLlIR/mH7KjEO
g2bPhz4eSzp62hbd4+OX4WoqYrAlyIMQbTeHStg85J/zSaFd75aomW7KJtEW
O+UwHO1Af7DilAatc2zlbalBZG/9r9Wy8fnOyMmRyoH3SCom2rkmIQg7KX4U
qvtauYpN1PnLSeMZDWoVBauQzhTi+RNsfIFOO1EKiwJHMGfgKIAlK3sWYWm7
Xgteniyr0V3joCUQOKKQd9d0RBVPXGcN1L2rFHNv2wBcHbbtqCu7NObktdQs
rn1tOJC9Bb1027RDXJxlsjr+R/HX63CyMIxslSgPNWC/kub2zCKFKgSrcZqb
EuZUhjatouVHGLDAqJcj98LqJsg26fzvkkQ0itTCinjOKQTeSs6VLZKZp9cC
FabGj1q8Xxnh4yEdUDr7JSLj7krY2fHMziSjVMkrQmcGCgVkXFghj4tEmMww
5P0AV0igFMe0mVJuAyLu8LlGKvqrjEWKzVlEh4XLoB9WsDt06sd8iK2XRxzn
7VN3soFx/ajjPNwzU4b+vXaEZidh2AJhtB0jMjOzVINm+OSktGpLSpOSkhyb
w+fy7l6YK+k6eAz07cgpUxmnnLOAC9ssV2WV9512NN2svA+yti/m41WEjoKR
cTN0p/Q3OBqpl/47kdJF9U7MXLggPYbLyq1V/R4CcSmG3M+VeCHyWmi9XpDy
mk9UmxvJaknYpqo/w+s3f5+0wXQsNuHS/cTSC/ykbk59s7rSWUazspQTS/RN
drhDhZZ00i+HDfBIMnlggG/HbmkMs8T43mFKD2sQXBgSDcInd+I2Hlq40WT/
GzvEQeunyVkE2AToZm4zm7G5Cxj6ZsrQQ1A7ODzEYK7ng/2Vc6Srp3hvKJYy
M7GcXzWjT4JMyGkb9N3pU6y1iz9+DgxLoLRt/D2+wStgOc5FixA4L1jUTQxZ
tjgWJ0EToOuEw7hNMNrMybKpF/oLXqHesDnJPOU9j8tTSa3mvntDXkgVqV4n
uguEIwboDWMkw+aM07LmQRUO72tCHaJzDNC+z3aBoncG2cU/2qpwU9kJRK2T
j96LsKYmJpoSETJjoRmhxiKLNZubvwYYMTSjdNxXbZW63nXcrdAagZf8uwfw
nMhq9jeZ2zhHR0IBYII54FjkzuqZznF2t9A4G2I6W9dCtV7dfw5lzjjw2RVi
ff6S4LrTjl6u9+rrGrTL3Opp77FXLYolkE2c5Qdk7KuOdhAxM9Vb1dncrEkF
/TWBHWjN8shzWyMtNjqoRqXIC2UdtY6Bh9z4EDQqxgDa6AK/QS/yKPuyUOd+
3413FR1KyQDHsmuzToKJUC4xWQqRbu7JueBpn7sK4Nu8yY5cl/TI8qVDohUZ
jzIiqWv6Skwkn/qbMVvZwN7FX7kngY9+EqroJGyz0wTp5SCnCssbUQWH8eAv
MR5lcm5LpKQoIsCgVVo26oqIV5gisiLbW4dKXhPpoMlmajqVbCy8RHFKC5fT
8asncoVnYFc0EeYXYIVx1ydhAn2orz4YTQsBkSvINaxnXZnw4g2MQo2890Lu
Jp/4wwSuIoEfr23QZcqrQnlbK2S303BpIaQUi4l1qcwMQUU3WxMwZt07XqUg
FStsytWtgcfec7wHsqInpQuTdfDv/MQEDoU6RjbhoEz/KUA1p0PuGF0WPgkF
jFskKCLGYOCkiC88yK8cqwnJ7J7h94ifwTSO2LmAWyvrAGgG5zyN61SKPv3V
NS/Xb7WbHbxJSWYNtAySlGs4+rG2QOEihF2fQV4NLdc/AcHL/JeheTAX+2dh
3Hn5FKCBW1gPlJzzHXXXgU2MaP+ezhTH7E0Lar/EXWp76d2IC/HkVwes/Hqw
t18RwFpXagQ/zPMMousJs2ynhRu7ezy+nNozIcugflrVrDrsYUpSjffSpK1x
K4pc3A8//zECzA+JZVE+fXwkwK0BWCq+Ak+FtAZq4u1ltNkg+0fcwujXhCyu
gb0AsucwUf/8SpEHlgy8gI+Jr5EpJTQyj0/HgJFV/nraFzAiS4Kk+6ocIYmT
1q2M4q1AJsguScdYLScweJKq1ZLWQ9oYBwiccRzkGyXIYJKV5YTg5rvs9+5u
JmL7DSxEHSIyNshoK0Ok+1ZA0/bLHP6TOL4M+Lbe91g/YSXroXFYXKm3vidQ
nSHx+OiyXctE06l5AYGUbPGmiXLplAKimM4NkAaaZGTJ+b7RUvKmEmG8rtRz
vJZHVjV5krYkHKX7j/8D1qIlPJ2v/yVZ9S2Ei+BbBkBePKM2arfXFze4SjqL
Tjx7qovr9bKwYVQttj8KHJdeu0ChlUxIjgFIcyPuxgfrv8YWYYKaMHuBr37Y
KqHzYNDb7rgjzRMCCLrxKi5g9fVMFPapZs/At5rHczddrh3HM0ycTRt4Al8a
xbVPfrvb16R7/b4SIWvioPU/FDCfTXHMe0x1f6E0qUinHygj4VImdrj6kkJx
m8FcWEC2u/jaDmyhdsihiqib9+zfQWC14jN3ZzfchNlSnBQhQEC2f5IMzknI
VebPrxyAiCWXBKkupTZzF2esDCumZOeQCVbPx3tR6MmCBb83sBojeb+PZW4U
UJKA/pLJ1Oq6mFNZNX2EprG5aSXn+dWHSpqHFjR8a/rIg/Z+Q1Wa6EBapOII
wS1FIk5HjIbXb4PMa6r6+6F5EEx/u7j3SjOULM6Rctlv1KqlKrf4qmFbjweI
Js/QYXKcAS9p330B2Y7LPKoeW2xf+jyYlct/CV0eWkfZz472vSwkcRlWTM1Q
mOZa2kEYHEUnLSidVJyYrO9tAgIpsv9W5NagoTN/LJISnumBxabm5quuEn1d
wN4+QWK/CkOC6ouHjNa1LY+rsndqgkecuiYQ1Wd6NJUCz9yvmMDZaEa3c61U
TuHgExs7U6ubBb1v7KBdzrXw+JRWxm0bjrs7ZFpEE8F4SjaT6RAAxNYXOWjI
UL19JQxAB+pzvQcU7cG1rVOw0QQF+s6cjvwfT2WZmXiitTibrl1GnpbAmknK
pueD8vPRvbj3EvDqfhVjD5Mrh5R9aZTekayYEMmkkyBY6CFYmzdCzk9AUe1a
rSt6jcGTnjJrSxbUrktGDRpHvp9jqJ/GYHWdq/wa7mwsBL5a6qSKi6vZDtRu
5hD4+SbLPwwbd02iggpUY9XaGr1MGfVr+kwq07VJW+1mLK8aSIIV1JnKaly5
cOefohv9evgm6C1PJxfr5kEVUh23idZSd5YjTveN8P3C0b1VVCzBfkSBZkf8
9VjJ1p+gx1U2ygkbOXLBnuAjkNYOPJA4+FLmlrjkDvIvOHa8I0VnwhqAgePG
vM/k6hOrluXUdLk72Yk93vk5Zyjs+SQzmOwgmQzTgN8R0kXHQh5+0pQ43Cnu
nHd293NTS6qhfHfu9DEASmZ3EqQwU9Tf1cSgq28BiGiMZDkZmb+kX3NEQC7R
4ZSNFjOXKkpbPFsXQLSYEeyetS3LZelZoGKqX61eNn6XLV7F1fBHCN/Vr5Nu
KoQpGbdD0UO6PGEBl8GxOXx/xSocG3l6FJwpDCyvlNGkDt+WlZ3zyHUGiPe9
i6fJhS8uJYCNkpCwXJnNz5XNtzKljI27N59yZ4bMaija4s65Xql7eeDRZ1Lk
iyXsyf93jgnMHuZ/726U+uDlswsU2h7EF+1GzMtpj11GEc6rLK9qDnDy1+UB
NQM8LX0jkXvPsR3U+Jo0RepBkZe48UdAGIIrCjIb6qnzqR5xXnZeTBAtyEHE
56ANsCUNfEeLXxYx5fMX5oIlLxdBs5Ym/1WULT1GBA0YDB4kkUnw90dq511t
kmY0+HP/YktjKwelHZWM98kls58MpFb5UmmZpY8w5WsJWbsB6pQVyXFvGACa
r+T5hZ6IXnD6S3UcyC4E+goUASL02rx8LJLH6H8LCLeCE/NYs2ZkhbkMAsVA
8tqmw6YEs3za6Hh/2E0aGg5lTfIrbaPjKLd/HV3Jb4fbre9v2iHHA063nXso
t2MFztPLyI1wH2cg7xzhzujmBWJMRDTbKeIoAn/xVSGucBWyUQFWCwUd4rvF
J/dUpHVBkf2AzyojSgNJSwT4FhmnhWBcG/Q/bdqGC5tdpj9UN/xxIJXG+CEo
iILytkDWiF5xdZylUIKdyQDzqRdmFkw/oAJWv7jkx2nbQDBV6EJQ1HoOyDdu
zTR2tVio+8265Y6QXD3nlZmUdsPHKpo8Zj77lnwCQLsBdG9vtyX74ZcbuO03
fT0HpFsO8LGfaFajmwmKEm+zu0oDkHxSZRbYeSYFqeypU5JoZr8H6xQSRklm
3zzYhtr5PBPcxPlt2hN1QtM5jZeqGzs7zLHIMNWZKeU2lsDtXazox51TPAO6
3E4kauG53kgzuBj2oalKxyOLli6p6rPWaO2jhuln7hKCHerC4cjnaYyPlLKt
4r14ggtLrjtb9x2FLO6JeNaTZ4q0FX2qqpCRpk7CCqZCqUAr/2Oe77A6d/b4
ATuWcc2c8KTYmtpblWNde8OFrJVZkiYnAWonAMrMC2UAvMpecqpGckgfJA3P
uNf1jLWHqobBevWcNE4gyXnLEGp6A8vvkrTFW1JvQ2OY9FTb2ZJPK2SW9m5G
vKx05Ym3NRf/+edJfhr7qlb+gAg6bJJaERKcmeefhTsYkwEzQbfsnzihU86k
e1mUMKq7qV6aluqTfTMiCQvukn9CW3HwouilmXS9eCE6j56kAtP1V3x+C1D7
3AumbZCliwcZ7MHHE/bCFfhDnW3xyMSEcURZCDkv5E38VoXSFdqavJtlaDsu
uucn2V0IVddfMGAz8iIp2Wo7CREQ702yZeepfbGXUmLlCEVT4AoLF8KjDF+5
+gnzK3OPTBC2GZP5gb6PKF0SvWTDbcDpmvb93wQneKbSiMYewH9dYsMiHiMU
Rxnvym6pdlraN7oKJam2oJ9QBF5UWpDqylb3isfR0ARU4IMWrikxoUgxrnvL
b3H+LwXYkKcpjurCy89tIbBWMRc37qKmaDrNM4avBk++i5ttINdmSCGek3do
h3zQ8GocENQvi+gS96bGpkSCN6Y8BvOf6VecEw7T9CKuPD2vT/VKwwEKUjNR
54NYOD2CzdbCABOZIVIU9heE5yLJksixYHDr6DtGDwlAsfMaHTD3IFfyWbce
J2kVLMNW3psgKSYxxOf7kfaRAvA6YL/gtLhPCUAwvOvSITAXvv3kxl6SQNwf
HPv1O6yTx9VAFRiljQEQlybJZkYfyPe3trUq/KDQqCOXPNaVpaSzHyo7SwIs
wb7mRfNcrPjX3OrxFrV0g69jeE9oZS4hk4QWoaruM4EIVDozdrqwU0jm4Vph
BWK2+V1MiDX7qKa3w06aBlXrQqF8YKdmLlI6h0fDYIG3VCh229xwtufdnkU5
bPfHlHwBTohQJJNIZ690p0jnbZzdrRxJaEPgXc5WkJnpY7GJJMgy69SKPAP6
uNT9KurgTjdZFZxAkcZUMyCK/MBKXuQt2pz7kg4aB3sa91c1b/uyhtoiDcVs
mn8pOF/egciqUnQLOkT6w437Ls9KVGVYiBBmE3MkYUO3jAACwUyziiieTyQx
7pXjfSTCZ2T0IgJrMY6wjpSPiUuik2MGjIQWfcDeWbBGzDWFbyx2WcnSm+Y5
6qrVZF3p4lXFzfrFz13zcLPstpAFG4FsanME2NKGXlqziYnU452nCYfJyZqN
ylb0FNNc89a6QeRRh9Jacnrrtw4i7xBV5zmCvO17q8xcA9raAiAAcdNfftGx
gaiZIo8/9QqnBvnZqCRKXPwkXFXV8tpkvqnpMPDLP9tgLSv+ByK61rv30D5h
upiiajY1wzjC5b1ccqaRxLZp2wd5G4VXNzjD3h81/K5pbKIxspS0mDomd7GM
2IHxs99478FFyqNQteFmdCV3PLlwde/B376m55sy8AY6JkHPnoLMUZ7ZINQN
xU9EgfRK3Y6fGny09j54ZWjj0EK3qFkWc+D/90vweWmdQMuVgEC/4laCBgdd
C7kC8susRo+q2O1GpV1DXIolZF+6vVl/l97yNlbGYKYTl5beOGR/uiNXjcuo
im85eW2YUhUimPH43DULbBWqvHqe1SyReTrm5hjMndtDaKIq7F4mRE+ghSDY
6qkc5m84xP+vY/ep9p0f0ZiPSA4o07BwDWllDjeBPwNQ0I8re9d48I+qds0D
r9Z9XqZe9jVnkgl3dB09QsTBuG1fp37OkFZym4Jbio0kkXGKKleUwEyo8dAa
AiljhgXrjGusthbJTk8A+OWYr/ovvVuzZt5ayUB+HGwW1CMU6NByg4c/62IU
oB7iRX+BP2H0CJneX6cX3NRl9ppxZrLuSI8kzIk7CAHP+FuXYSDAoHw40YJ6
d4extqGFJWg+chZcGnpvlxamueFY+hNx35sA/kum/xgve11Qwt1lsq/fkIbF
lFlgKwpS97RofQ0Jxr9/gNGjcBt5c+Ojxbb+NJ6ZdI0zNd/NUin5Qzd3yxmd
W5XjlBesfDSX/0jOXKBWMR2VCvU63Nqf6YMdbTY3MsyqTtskfK0tBBTj6e+U
YmyLGaL5cnndFrStBC29jntOj2Csy5VafQs4nta0QefDEJl2SIbxJXxdCpkN
NybgQ/5Mmjz6Z8j3UwTG2Wq8y+24sTaMWSnhS4CT1i5/6zMLo3SX3BbtT/am
/sYxWiWRItcjdu+alnGB9CXzcOEyLgRMNgr905b2zVgRrCNcDzQFEXjhXEsJ
FoWInOgM13NOF12McDP6pFkuIzL8NsdLk8wSzebqidfI53ThRE4qCp8dzhTo
woy8eHP4sG5+g+q9aYJ0ptiwajSpeHqFH0Ueu7BfW8c2svM0n77yVBzakj4x
9NjVAy16KTt54Psf7nm4/zCKIhzvB7RROB842uNmIH/DczM13eXTH0TQZT87
cR6yck/EkQz+vM05VlsFWddc/wYgLyfJsalOlrs81uanPDQ/IJ2Ul4O4TT1r
aoDc4drwbewX/c9bzVi3LxQTYaQIifRWYF22xB13C0EEiJjxmHT3t03zYTpC
+h9qD3NPkQPlQsSYaZdIL02/xHf3Qq6jTsaBCKcanrpIvFQKuZzUWobbAfAf
gvMq9dXE26PHzlKZsLuornRiG2T+KGG7Eep8yYTibP4zuDsiVYOxz6irsuxC
UOKeBdgr+W/dxvKsut97vNrMkzaJZEhcSmTQs4Sni4t/an+26VYkTmEgvnlf
e3i3+825598de8wi2ErQgdN8EdVSK8A3sryuND3dMzSc2YGSAP1dFLqW+Ces
Bh8eqMqxvG5vB7M0K6gAnyiYxhx9vxWp7bdhFc4zHPOoYhd4xHwXSam7ViKH
x3ZMpshAurbdQIBV/yo9ccdoMeuA5vuIqt32V/3+2+AzO4wuEd2YXbkqVdhn
9n8+eEynN+u45dmGMw34eh2+ZC/5LudBTaJVu3ecX79s5u0LqS6FeqshqrG2
Aqua8uzj8NLJKlM/GmzNwAxrPAGDqegPDVCNrSIST/zbV5e7TTz6jmpSkyuD
pXiqXaRmegbZ3ieu0SUmhs498LnMudErXQ5i8UoQk6nz+NRpwn2gFDnw9mGS
Kjo9/y341l7SNPyfP8iIvgb0+AbJlJS2PltYXhga8hnM+LqPKg3+y4Cv/dBb
SpHn9ZlHaxXZesmm0Ivmx+zlLVW/a3KyfInR5FgCBZ6pdVEFDWPf6wLuSqqt
sb2eFry5IlZAxqSlRuzYDXJFBGIYLovXloJNVbYjj6WWM8WL75X2Z4o0Nz9E
JGnu6yXwJwQKwsdoqjamMwkPpYfAsPMCRzCHfih60VL0HbQqDqpQwL0ld8ep
EPV6KzCorMH1wPA/119O5YnA4fbbkQl0ZKwHCvH0ySrLuosYmHpaZIP/o7Gp
OxFJDgFYko3bxcqoyG1JEVGlMPa/0p6oVSsnS380a4Y2IQRcRa4X2ieID4ZX
lPPWo2g2KptftYQx3Lmd/q3P8R/FM0XOGzVf8NvBTrNfdla+aCq1mqT+LeRp
zCoyO4wqQudNO5/BDJ+RqbxBTS2Of+mmnPzB00q7BorFUfENegflG8vBeKHm
cAV3Th9jCK9faQcjXSo8haCLjd2Y+20hDDCJ95idDQhbZ/qE8KIslXQut3Db
KblHvYfuXYcfg5dnJ/GTQa2u5N9GVzh5fpiHgZdLhRbCjQXzAxXOYwfN3Nut
hAZa4ZxCoJmap2Dmw1iwl8Y0xEzQA5Hro1UpguE+0AYs5FfHjpK4TRpnsg4u
F/Cxqg07NuqFDOq68f8cJteTFFpsyIqDx1T6Lsd/0Xa3jHXtvDn0LzbOl/Db
SGrKO7NQcoPmGBwPSeo9xjulBCZHSvKufTQlkySFhwY0AGnB4mgbb6ordPHD
lStqfIDbr6izwae16L5/Zii8Xcb+hWVRDbw3DZN8LFJCZmlEQMM54SiyaKF2
JijK3hWV7XqwLzBAKctnL9Oa85OTYbyCQeDU4ZBqXZ/mlrTaDdSHQ1yUAMqI
deikkrb+rJOfLceSoJgRnhtHF991Jn7Mb1phSXjjlt+15RY2l//te+kNceM/
GkYBLNg6fiSxK2h10meS1c+nNB/GVMfr7h/wZhRsR0Ur/xJb7geObN3CHDni
Ysbrci6h3+Bm/CH0ZgSTQzPLh4NFo7Jqy4+kMZ09tjoJkAu4rKB8BpSXi93t
8Omc2FRyszQokDyt7ydCK6iRhYGnMBZYbG46k1pRE5UwsPQuXanu7eKcHcNW
CjSnMfi5reoj4kaeud5S7/XK93v3bkucQ75GNPGOVGZhuj4em66ZnAgwmSP2
qgVNPytgtgQm7ziWxaSeMqkbuJSV1Ak/3t20yV5Riz+jswCLxjHLYj0Akr2F
JrRGkSHG21ripwn7F+8ColJ1ButacfqZPJoOBZvtnPMpeS2ebm4GUs+eClwF
xwWz6GEvrpH9PYz2jbtHrA7w6GY5fz7JX1NRBGvKEjhbYfHVeyWhGbJJs0jS
lYswqdssI8J5IzioVpAUmRojz6HSUOQvFxw2aYvVePGGiMG2BiJ1tm8iWyew
RUIuI0GmcUsg7FjVmCfLs4+za6vJrXEDmTMGQFgrdmmqwLtXUx38SazGtH00
JT0bGMFxCUA0ZvSUeGoH4dG/WnmAjBS6zwaBSZv8/B0DARTLT8CCaYT9bEVV
Lwe6bsFyuBm4orrICgz3JpYv4GgGahTLikte+8bjhAc4bZ0yekHE1eGOsOxm
GixLllIUx38E1YQNf6Uv0VtvHnU3Soy1pQRmv3Ts7UQt6tG/FuYe0Ki4CdNQ
VtJMgUlrbbvmtCWaGqfPyGyjVzYjg1Exn8XKuZBwOZmwW9O7vGDiOXgecQsR
0mu/57I+g/X4Xvrm+Z1ciNIJFI0nlM4kpusBGKtFnsldZhYZD5+n2QdtnY1R
DlJf3+SqIN3+lUawiDQ/hxXWonUOwgbEXU076RsyVzPZLxvP9qkYvVw27uCL
S/3QjBFCS941j2TLDblz1IyhT7QxYvsptwDOlkUX6flqFk4VhmRU8AKvt5QF
PCU4PUM2/tCmqxrHIE5ffXLVHyou6z5lZzK9tr0ylEMJ8Vn08q+8F9m/NZgG
tJgGcq1S2Zt5Rvu2Y4usT46d7x0NO3MzW1o2GyG08STceGTlP2k9qzKv0V0n
QhjVZ5N1asxwRGh4ia7/rv9r7jilq0Q/20THZQjraRtDx1NyCDG7jfxHCvge
jB34nznoYMAW9GtiR1Uid6FWpe23fRZm8wAvMveuYI5npEbSRymll9CiPgOw
v4N2o3QHN/sdVN6PqJ5x5SFGYDfwzv60dXgJY12BFhQciwQPIRvkaK5YNVWU
/XBNCqchXBFc4AGiFV8+RelBRyyM9KFZoQZliUuGAt7KGhCPdgUZ++PmsJM9
UAo0h0dCey2sjPOyKVt0lj7DQMwoNvdjE+WGQ0M3uswH5+5yWACGkBKD8xN1
h32p7OT5eqSCVCfERyquCobkK+Kk4QCNGpfXBSSUBlEKbAObl8e+coiCacMk
hfW6/d022mon6OyP4odjVVDP5b/g6UcwRcO356pkUQOFgBt6xRsJCdX2CZCu
P71U4UMDd569ftez2cZbBphe+RAaYF0r/zmHYuF17aoz2TTPG/goLiUqOaTt
rOnlhMZZFudLHSAlgJHTF0dwnGczdfsE41458ekveZh9nISuzdBokCBzdryM
10Mv2RPpwmQA8OM9O13wJn0n7pOfNold8GAWUdI9QdwieB2hTFObUvu1WQDb
8iSkMlzuSRUKAvROQ4OMsWqboRRks7lIoNnPrzH6kQABNZ20J1jJ0kdTL1ne
Si99yxFqFIeNL0Ig2ZVZNMg/FG1fm1ggz7YX6ufAzNVakmPlipz9qLxH/LN8
2ZoNA+1DinjMirvluG61gf5wUdnqCybxYQ9nzCqlvIZgqxXECX7fl2y0NsCo
znLRb6ey/plYOcooh9kfg7PymJo4XYPC8K2e1HZLhCVh02tD3b0Q9jjXEAda
xKUXxDzWQFmq1ZmXGAslUGsVhShoJdMWdj3kP2msQXIHQnrEyuVWCqedt2BZ
j3Yv0HoJexDhxiZAf1Ljpagpnplf61GiIhz0SSw1cc+h886Rjx0WPatNrVa2
CJobh7Y9FZxRfFqN9U/1aV7lpEGHHkxe4hx3hYv1svbPI8zA6MupPPw232+v
VCE1s1WXm3AE78tjn75GZpgusdN7tlyaZ/3oPh7whJqk0tspByTzGqzUvC3q
l+p0TERprvO/nSNBNsL0bByuJzmPge71X56vHAk7MAVXpKs9huF9AeZmliok
atYyBDzRzObt4AfqY3Sy78yMxs+tnxjRJ4nJWeALXTJc8IzXBhYfjO0CZm+c
Te2Lj9kXhM2FzsKs1VT954ZpCSbtdjGdcGSa/ErIzLk9R3UYAEpCKUspigQ2
uoCXgldx13Q44sW/2aPbx89sE1CoNCvdAkbWC964Lq/DSLpH+wQ818IQjPzI
lALhgZVjSDmFF08pKViTaSatvKwFMn55xMfQjdGSr1eyCfZKnBTQF8VW0fgt
M1qa8UqCxAPYni72taad8vRJFb87CoykauzJDM9OxYerSxClXCjPCFQpBAoa
V9Uudk5+xzaVuaDJ0/QNPBEwuRV83WPYduExfRgloF5UUmxjBg9sKYuaa97/
hAOMS5fnvqVxbD1uPbTt8sIYagXvXfMfrxwbDuF7RsltjQyzF3Oe67sOXGV0
6A4Rubvgp7/bDsY5csbCFVF3derlVpRxCfW8aPM2SWk+Cibg3KBSOCc1WqN4
tKy0X/Oi1nWDKdPvmn2D2pX2MbKxr+HtjkVwpFEkHPfAM7MzS3teK1qCD3zP
lOGOuEEbkPTzc+mBoiHXz9g/KkyNeFo5r2xFeQj0vj5OysTRoWp6SoNdhtPZ
2ZecVt7UNKxt1AUTMLt9LBk2lTZV6UdMsbL+w/ZueThe/veYJxIxky2OSKFX
mSKzulgXwKx559HOejPhQ/Vb7xkH81C3chJIHDgcG2QxQ+w9f1+fqP0pqWvJ
cxiBr8xdnN2diCm/b4UQY7TRrLT2ym4MnmCAui/hJAkr85Ga1dKpP70T9bO7
qieXeK1H2z41gMADaE6xbxdpXremG7RKjPlT2/1E1jlcSOC0urMyZ9NnxMQt
KMObCA806yymhyWfDSJTl83e0rl8cnzcvB9mZ/GnPV+6h2cDRY6mQKwTXXUu
4ZTCkilVSLrRx/JVvgXcuGjFouPKlfdq5fyA3VItm9YvSty7GvNv2tM8U5I3
aycWCUMTOVuHR+iFZqZdepTKrMBXb0YObwm1n8CqSveDjUPmWxJ6q3DjQzHD
tSi9TEfKK9YVuc2CBWH5udk52euWM2hf9ZwMt4c+h+jRx5Okjef2B/PvSDFt
K6hduagdhWmos3jsHABWWqblX2T5PkBbjowwS7VYAciCLn3U2QICpwK/hQjk
hVgdBy5gE/mq8hBcYxG7OTOluI7d+FG5iQAPtRVeuKWJ25DHCfERYcfHDRNO
7G6CnF3iHA24RwMZe6ATjrFETquzg54mHM+HlDmJqIrTq8LUPgVOtSVAD2Ai
6xzdzhvZr4oqH3q0+kRWOZisQkH0RDBnVRsRTSnJ31jZ+2qY2TIIoJI3sYAM
FaYV89eANhDCsxxUXtrL3q6b13LAn+lswoi0OV83ZtSxxpVWyw0IGRmYJ3AF
fyPb3FwGpuHowUvxSc1hn46YVApOXiKlNul4gQPE8cSjM807LozbKXmGHwdV
WbpHKcKyE+1TQYL7ojJEjA6+PJ53Z2JMGreRp1RO46813kcEW/eI9zZNgl54
nLsXR/huEWjrADQg8Q4+cXJAAJknlIvYUqHgVjZ0LhNKJ1XP4nAb9uF806cV
w3s6fXJZRq/0DxiDQeLAdA0z2OJQtK1unsnEism/Ske5ZxHjCXdzKew+bdU3
PMqNck/62mC88UAhkP+aVQfwh3S+FHtsPCiLPLa8P2mF9ZZVc47Ybvk4Yh8j
gWDVyWbEa+ipLj++8yiGff7AI9D1eGxwZpx3q5GWdUU7DYsiXLtJ1mTKdcLk
oowONXyGr5lUV4Ts4jmOH01oWyeSeR37eQ2GXkUeEBFvgzASl3JsUR35oWq3
UYTRY50g+vh/VQXYkJ6YAcs0B5qS802XWr1vqBaF882vKlTVgHnSKkppY95w
RuA1Spnn+9Ci8dQVkDXMm8RVzn3cSmOqSRaA/TEkJGCoel/hyGmqdxhFWMhr
Y07wC9fxXGwKF38zVCBq8shHaV6cX/f5n4d7idPOa8Nk0z+df/6cj053cT9Z
HKRUtUFoh9AnZb4CGntqfO4eByon7p4dJKXWPxL2RTerUB4Wc8KldgGqAoPn
BFgSPIdp/vYnt+SxxiKqVLFeSnEhsaLPD7WqSI+RZz8eBUwfY4nK3HrEV2PJ
SZ+o4n506DHfUYaSByUH372lfS0RsDMU66x2vNjYXiQv4TJhs5csA+cUPgb7
BJDg+TKilcMBRhLLfPcd8DnSTmySawwcNF4ucpKSLApqzs3gY64k0/8Ro4rD
fE72hv3uPGbQvnWt53IwMj7MphlHMtkCalps6iOIMN+FFwlhfmB69rvVuelQ
1YGHLBiyjwyGtHI065r6RpjIbPXU6WHQyJsFiJ3VMkdTPi4ZZ6y1b/+YOLOU
OVkxPA/PozFQ1qJ8NVWsyiMMl9zZO9oKaLStxzYnpLt7nioUAJeDaSHC4+w6
hIhubuWSTzH3a8f73K+gXvOVi2yBvYjVnPLbRDJkHxOuSbRBn7Cc4zCSOdfI
KCDDsE7Tvj1IxmG/95RgN3DBr4BV7ok4KZYdgB2UewUDqGDb26fK74EW946q
U3tOhJqkBoNGJDmcfPFI66Qtood+R67LxKzjYbHl78povTeRQiPdiv2bozA8
vk4ZxYmkq/Cox87g1CvLygAU6S9XdDA6mjGPvoRwNO0a7Y6E7BD6bIKhDPNT
kG3lPHRp0OFU7ALVMRrZGplalAaVaUicn2iINze/Rb6KEclde7K1Cyh7FdaJ
69JcmeK1H+kNJOdBwfImO0Zpzd26YziSh16zyhE8g+06+0RIQKuUwdgoDY5E
9rDCJVc0et65grSujhPV7m0YBDP8lkMsqP1h+qbr9ASDxJUhr1SYAas1rxIJ
+CsI/jaA56SDudgJJSoWmV1WHdu+L62zrK2FmKZF7591Pssqdod3h2dhNDla
dAGgn6djp2bjQhRF0ETfS0pxHKrjoA8o3AzIF18FZkrZMXEZZh65bjwXGDCj
jdt7u7uIE3ws3JQjtNvvWN5DsQ92c1IESDiiUfl5KsLF0gOoq/MORqR0sPFz
mY7PyFo5o6lqqnXtWlAXKFnB5uBbs2U3U9xKufMEp8kW0vzyGzueS+keZHwE
uAyiwhA1F2Y8zs5ZumkdDNgJh7Snyocxf78FT9tD8qzxZMZMYicTcGz8buBJ
I52803Sg3s9Cwm6FjtCMOigyhtR4H9HmFS/JWlqIqMG/eqbZb6WY2ANcAQ8N
Wq0P/lQ1c+JwjtsYvurBoDijiKXJDdCPWk9AJZg3EH6P2btFokAkT29nKQ3d
/n3QEDxS+Vso9/UJCiKM9FLhLic39AZ71QlYCkDCPYIwYilPIWP3J3/ygxD1
KFm6997Kpfu/pF2lEwLKP+5lKy+4Fgk8bvPwfA10JRBf6QdLYNhWEyE4Hx1G
CvJkhd05aUFyMuglCBhiH1NPLETsFtcVqCkV0II6SoM5YpXFlX54j1nfNpYI
A6alkpTogcos00WakrR8zKwkt4PJYr07K36VTz8S1OwLJLXCd+RZM2bDzViy
h6hXqZgK0gHE2Ey33a9CXpF7HVsjBe2fao+1EiZw6Byn/bpwg7H3ph90QfoC
vaVkoy2TasR6oUAmQujEz4ST1Ppm9sR3paQE6xslDbBALvk90LTF4Gr/rAFc
xgzn3iejBOrNo4mU0F78zEAa4M8zHcSXXROUzTbkXDfhsOkZr+GhXgWhEnCn
kT/j0XIqrgR1JtSkBhgQ/RuaIgpG0L80/N4bUMHV9sUn0EfTuzX5/GpEdarx
fjPK3hLMo+9vcPwVVaRkMkzNiMij+LGv85Zm1JWL5WFtvVMD75Fdjir5t1OE
NIpB1bVCoMnGJOcaKGZOaAiW2s1x8EjttCQKXAjq05kx7tvnjBl9xg+I9gVV
SLlNpDT2U8/kFlFGQ6vljf4XtXYTIkVdX0U2XKu1DCTZKhh6sayMmt2Mc+Uh
kREtH0sw3r//eQU0xdQg5R8jv+LSfxJYNl70jcZj7ieQv565wLB4raeDCoV7
YVug/ZJQoaQsAH2uTMQUNLwk3C60VY4aoesXBLrC3dX9VYekP22JPjumpkuY
7CLKrSGg15b4Z786roxzSAF+8k2l3CCKuKYRr6zCzSLER7e3RHH2LND/cnHx
BuXnFwuCIgoGNbqyR+C5Bprk4Tv9iAjwJQ4Tf+Qu/Wpr9CgPYCZ22qFgI+Hp
/1XD+AdZ7uLj9UnHCv8AyiHuaoGcghl8Kg144LLgssrnJ5SRI2ihZNaW9ADJ
gbuDhF1/GTXYDZ64ZhiDOwBi9eEUSsfnwSp7EINm3Vk4kGpfUUJCNoqFcDrY
Tj3RoxqZSYIrropuhFS5Q84OUxx5XRJanqB9MMwQ38oCT3kBPVJUyHh1ZZqK
xSvj01kgdqvLEo41y1sTDZ7xBEQDgB3DmE9sZrcBMLPPy4s8pvWOy5wDHulI
AW2QuOI5AD9EHm9xkSfLXKbdRR5COe21oBxljgVxeb2WAySfVTilBs2ZjffT
2SrjsiT+TWqg+YWqLatR9Yd5X/ysLP17Oaw9WCAStfH/mTUNpyR4677uK/GL
7mgS7mw2d60vKUf1cwSVu57kXP/t1n1/t5oYtbriioJXAUiJHg71ucRGASXS
iv7yq5Jnx1DnmpmGRrM4Kab/OQezwEU7+GIggeAUvqVQPPsCemalkBDB0Eth
ww5xuj94GVxmEni6xHdEYy+N2CEKBvsc6HUMJ+a5mqxdsMn4CCePdiqAv/Xk
q3Bls2j6xNFRwPAGE/0EL39SfFpap09gkIKQo6UteH9OkIHNZXWWDijfoRb4
H+CfFJBqkISKSE4BklptiL+A2bgCd1/O+pgFazABj4ZIW53/7LifbeWxyUFr
/IsnUKQmJlrWZHN0kfgOwFcLjfNjQ5PRfpcTJaQKo9DlD2kXxOIEbwTLqkSS
CY8zrzyOZa1U/Gm0zv1GYxKhsbXyj3JpfzeKKFPXnsSGFFd8EgHsIoy3sA7L
ydpUSZMR889+Y1rde8dsdjAqYDsAA6z9wvcJ1ExWG9HLcGTpb5hL41tptLgY
p+kCA3vYuko5+T1pKjqJWErVXej26j8oTEAU/UyFpNgT08uM50LA4TxMOrYf
sa13EOQEKe8cKCd88FXDEvDUheHd/voGnwQNs0iZwh6IX73wMfKQQyvJ04wd
DTOl8LiuAOa/04Ra3ZhJx8Nsk8iTJb2wfAaZuQggL3J2W0NQXdrIhSDYfUAl
EAPiJNbMr0V0bdhKcaoR1j1JGugjUTg9jP4nkMJhadOiRKgTT0fp3aPhJ017
3LJp6wGl6bu0cCSHylWDzD+dGTi1tA4sz6CjeNF7OO87rXEE/Tim3Nrr+VV/
kYFkfE8WQh5awOJg6JqeCrMB4D5ghWYIqF5mJrqyulqonTADFTVbiUCD5Spi
AXx5kKKe8YPjx/R8xaizQEv4dsB86pvRIxWofW/Z4seSaKelviNv14NCzd1x
sR9x+/vvJ8IIWxBpvSEGH5tSo3qr6pFGN8X24CR1rvwlWPxME/KgRIVKWqHI
IqO8Wjr2jsIaXzqOr7kzcmapQyns76brFL4FIh+lOeE9kgwaY6Dt6dok7irN
62BaxW4uXciksFEVovUc+Yfch3Z48/mb125qkdQsTYLCa7EF8L+0lnjBoXe2
kOJA/3937ChBwLKv+Mo8K30R9L4JB7lVYJp/vpILQB6jeDEwz1tInkBCsSZ1
hXKjlnXOS8uMeEg898V1Rs9Bf3mjWFaB04/ub9oI96rS0eK9L5PSKiT5z9NM
Qy24eVtb/K0B/MnqFPrZm2eCItWMeiSY0rInzUJ6ToL79aJQb+vZFMIEdj5M
6p2iGtk7EJ5ykZ2tU3FUSBcY3Md94Gq0gfJW0RuxRl6McmqUIxMGrSZNHKS2
5znimRS06imtI5uR55JTV8qOwfCxz8NBJls4XEfESQ62plVqRoRgmxT51PLj
Yau5Me3Pk1Gqjx0qiSwb3CfJ/ZeNYL3PRWF8tie6T+NKvIu2sWs4PzH3seJa
00aliaVX7+UTTjuOmobaFIXFvfec4isbaXNeWq3QI3TMSmc9yEZazmMMLBjZ
0u0Op1i1IZqqj/uMOKpqXox9poww9YIELki8Di6y4xokldsrHm3KnzKWhh3b
sp28TfJDbYY2dKVd1x7g8P8+CZqlOBIke/U3p46vnh4unuCtAwrfNxYqCp1p
qIhFWRB3gYsxThyw0B+XDLVxttO44TuPQj8VpIXfnTpVpaOdB2f2D+XiOAS4
pChUWWpUBwI2HUlfz+JlaBdwqYwrXYQugQvS9DF698p7wODEg3l4xxe538am
5zbrPRAWXNurwnaSXxQyQ/eUCxYu/D7pfNn48t8KqudK6ricEJCJcmLUPzY+
Z06Cf/RyJTxOppAnzL5WrQKK4f7KfFNgVMpQSpzK7w+WGlGorSOBddVK04i8
YEZ907RBQXT1r/uVdSzS87pbyy7isRhpGKLw0D9uxEVHsk4b7aIX58v9Rb/z
Q2DR69hiRYVZ0n9lFDBNcUP4XWXaK8Gwhv1Z2njLTwx20Tzmy1zUMipz/3Ms
1Hq7tznkyN7Z0TETxlhjq5xWN8ep2BmdLdlGj0KbDBnDGEC6hqOcckZPqIQQ
96xIHqPyOWt0Y0pTxkhQkbjtHpT+yluBHVdiNcKyNiAF3lNvyVeDGcrarcpZ
MQ4DONiM3bhvtmhtd0kCxX+2PyLM5rj3j6L0yyJBY4c1Nqyt5nGFMU/bJ7+Q
70mGGOOY07BJvHEitmQ6Y4uZx0oQ8sBx+JWaJ6BdcubdmOeZB/JJeZp3e2hx
0V7t5mCYj/hXOXToizQfMt6YW73FY62/+I2k2hzHWbOnVwcYE+rSk1i4lbyG
JUe42mN2UIDAwlk1NORvzCBEZQ4Y1jNnx/oj4reA/8oN8+xHs8vBOBwldl4f
dQAzJ1I/8RI8jAwhV8J6UuJ1ASSF1dF7l9cpHRvEzgtcjtlOBH2ukGpii0P7
8TfoEncUjaHtihwsI/8nIz1UQwRtBXIE6sWIygbabBsArP1AC+tmr9lYGnLb
N5jTAET6tRWOxBcr6jpCq4Hpmv9gpZjdIl4K/5R3lIoK5LgOK2uASetFVQKC
0TR4nEfVzFZ+D5s1uDctqZPdE5yq3SUmAu2euycbFUc1uNJJAZVrewL03jS2
ShprCfL9fMnTPV5q9OIpkKifq69dJzy1OEsB0O4G+ao0fJ2RNM5gRY6OWxUj
ckvY87V9kXSX8ifa90zsk5l2h/25UlwFEKM1OUsgAMas5qbbem6J3sbPiapq
7qlbS64MxGQt8lQgISf5xmN5/Z663WeIhHF/PJpGR4fHkCV0vjdTgJKfqqbk
CO2O8Hy9n9TihmN7pyuMdBxhbCWWwkaV3ljKUX720f6+m/D6xalXW6L11/8H
zne1vmUz2gtroM85imwPlTdglBB/zJ6Ns2vaWhK3ldsAIIlnaHB+MUsqsSXc
STQRmzmcBVYXClcw6vnRvZNtDqhu+GBLsIkYpOB7uYvf2EX2pbHoqAnisRh/
NUcdeGw+9IUZL8Z0YAxcyiFN8mZkK0ivMcSnudLU3/t0rQd6Nlpi2cl4Teg8
9kBBI++kite9sWlhTsOxx051/Jssxl5bAVCwmyrgUhajUqNBjZmqJ2eLpeNX
YQB4E1r6ScOrLbifb5yWtDpjDS9w4Yg7VCG7GmqpLJ8zb5tLmT3pyV8owRX1
b3yDFZdDv7fJ32DZOxDSSwZxL3VyyWE/pZrZgdFHy5xvwYc3ErkC+B3UBK01
4OC+Gh7bx2oQQrTQMTO5Ks8bTI3+3H9eqckkR2vahut1WPzLHneP/+cf4Tkw
hD1XUyPQCZw7Anwp7vXNQeEB4iflixXDZziuQaMcINDCW8REYgwNsCrIuB+m
4GIrb60Qo+AmBs5EkjH9iJq43DoIDGMSL3beOz7tCa/i0sxx6zEsq4NPP8BH
efbihhlMeOJNU3TtjVhz61qSZmaDpcv8C2EBnojqbL/VWMYZ/ad/GWHkE9ta
j8qf7XAHERst0fYL+gnQuPQ7/ewY42QNR5OYiWjdg7BCOt/kAfN/b+45A5qG
1wLSoiFN9SKaVvqr8j2iNhTUqRRHGvrRukRtupeC86x8pU5oAVmFRZ+w4Mj1
dOsq4KR5Z2dSVQZ/X2sxY+OJvaiRJGQOnm89b4kLBWzh/0Mb0L/BNLCJaUHI
4xj9A9/3KDwrBlWz9zKcEUR9KiQ1crZ/fMxq4Wl+RmhdIJwo4n5nzYaZNqsz
QMdGHxns30g0LAnAxSr4NgZwOjAob6VaCK/eJ4cSaWp1s0933uPjDKgHw2+U
HjSJ8Uv/rReVoTbYM0A6KmjiZeQvscK5jLX6q8uvSgha4uzxvYGLlWbXnNbu
KEn4NGD50/PjQV20ca04laUismoPhc6RUX/SdofvWINgI6U2IeRySJ0Pk+tx
R6GT5y0VJcDb0Q5Tw+9mKTfLGmVBTZeUppoRHRt7ms99dSm7tclp/K8jcGAM
AQIjcccR9wiHDMBgECixJiKbTeZPVj6+2iLqDeKnF7w+xISTrKWs7Vv/3sgR
KDM4J/ZNHdpEjy7NUY9p6y3zvgNb4I9qb0eKe9Op2J+8H98v/p7oRxLVZqr9
6Ru370WNlbQW6JbdtIhrl5+3tijPB0jKzuh3VMLj7+CQgM80MPChSeuD4BVA
V8a9j0F+sXeHOrSjntOry6yDcMe9FBDc0LYxCB52dd8/128AN6zbLlOU5pVO
3kUKOCcevMcp3vSTnjHmPyBVERmdDD2kcavIzW8JBFmF70lXF02229JFPuOV
EoMkTXXSoA9JCBImcM94jmRjulA+c9M27Uat07ocy2nQ+4dP4wImdy3hZ5ir
+pCmGalmSsRsvbKfXo4QuD6y7PIjWug6AOvekipvY9so1YfdxIGJYleIYDmi
FZA7nb7hiWDZgqIKkE5PW4kdxVtFAHT2K9JX9aYlWBFQnckMVYD2RDEMjlkZ
g50Ixaa9nugwPvwaIWfBNIMC7Mpfm7PWAk5hfmUcDVGtQVgpaR7yA5RMUR7U
vrXyZQqgzM5r+LjcuY0anieQ7A1ECE05jpvXAmiUTkAjsJ3Lg1pedKGdyUS1
WG2wdTKEpiH6SBEqPGFO22ZlDWG5HwtCOzOsjfHkMEFZ1ax5PphqEhms9+O5
6eTicW99I0f/uMpcf3m0aVNIV2YTJQaMLgVz5eEW61v/Gzo7Eh6CO779lUR0
pWqHkHNj+BEbYnnnzwHiQn6cGwFnrT3eNbwUMQlf0MhVp3SoqunOEIqPPq4q
/aODN6uPmDpvbtkmcmB6HvpSs6HYOrVOCoANsf5zToIIYtqMRKPCwYGmK76C
IYGqP09ulnpElE+XbdAxt1V/3pCUBUIyppGfKBIPNkEIW7tIyBSmPZeKCblJ
7vowqxvwJv/IGw9VDu6Ecszf4/IMoNjuziB4xkIkffrBuHn0xP/BSZ4tsIQl
JBYefVY+kQ2sXk+t3f5LXgCFR7VHFLQcqMFK4hIj0OLiJnHOGY+2r8Pbd6Il
VxeyeqyIaAmj9yi1XuLmQQNIG94NbFix1/qj02lFIsgfubmAedaNp9L3hcIl
6zyY6cfnZS+SPO6YfEcVZ/5MyeeB38MUQw5VPMvWnVoaYpLK9EMgI/m/TNNH
b0EzTPnmxIURLxnROd+Phro31SyKdWRu3N0k5GnskaTFpnt+KROOXg4A0X26
vimhPLz2cKr/MeWtsxJSKOKyh6jxU5DsoSiOiV77NJWsMQlHBtAcSXM6Hf1t
OzdARhDRW/v+4zHgczTPz3iHeARJLYJc7LzyJkG8d/VJos+0qK2q5VWoOL+7
v+EBsvahSBQQSVTJ7xETA4s662LAsUbZdfH15w+h2rjSKn/m+ysfnbKTptVR
w3gwlZvFXfHp5Tq44gNkyHCt3HgFKUSJfnoLtL5psJTndf7LdOf4LVHVa6h2
Z2G7psD9VQjAtZD3CAI95Q1rg4dlVmrWndj76lWzOeNCasL/5u2iDxO4T+R8
RnFPNZM/5Y6yt3cPCU9mGOvpogcyMxzHanD+DUFGPqqf2v6RYFwwyMswAb5F
34Hq7boDhpSaI5OQUUCCYJXr8N7ClncEswxqut7xg9Kzirw1CPmMvFB1+c+u
sAIm7+g1qvWFNQy3tk+fqgcKBRoO0QfQgORdXWcfL48G22bpTkRXHSX9iPIJ
MvJRu9zXioCno6+V8x4zTUfVPDhsaySVIn4Ee08l5BG8CZpfX2TqonHIL1a3
1h8wbRYvooNktiomojndSsugpiycynVB6p2dBax6TE0dwzJm0x6avUmLmHHR
q3eMYb3FE5Og4d4beVjBbjqZyheIuFSVBsGjy0eWdHurW2HzNxDZRlSq5Qdi
mWmdT2EVmTNhHItQc36BmTFaliuaL/eP7FuhEvCRegtCt2bjnGJ1fR5rCTMk
69LWOL9SQltzN98hhfSharttfSVew8eLcGmVBUxKGukJOGESWNK3RhntSQ3Z
fmmULChDXZGQOLcCky4KvaH5U2/ONiWgCqMDGJRGLSrrqzaj1tVFixNMZtAr
kniiNZN5D5bYbq2V5EEDyzq96D1FDYWASyzLFZqBug25eBo9S5BrRT4PJPJ/
j1b3aALcvoY0m87G5nkitEUZa3lAVnCWrWWm2VXTDUSOttUpQ6s48eUHGLWp
OFAH/qEAaGy5WEqphozSVx2Tf7SyckokGFF9JSwzpo1J1qujEJ6HlDzQKBR5
shROba4s0760jiR8tm2Ul+AdUlI7uHt2YE1ZPn7QhG8PyfaP/hc4fDYfKRQm
a1YxbP8wNsjdpuC/OPFYKW95b0M1HuKJCz3MSHySzRj/2EveGNgb5fQlO9r8
NwkalM9fBAvwsDoN9ehtc1M43oL2e8U7Alqk/SDGifPZm/KVAvA1ynQH7zyA
8I2QBe3rbNh57teaDeAUElgHLHR/hbVamM0IZUHn/eaaZ6G0y6eVeGTJxPpY
/OVX6gFPaYZtpy5+Eq0DJjB9oazfro9jj0F8YIPoy5HJ8pfSflzOr7m1tQRO
6W2P8hj91CFSlBwYA7fRSi8JbNZVOzWDZGtVoLsFP7RfclcPO1CqJRKJ4heo
kBMM8q9GFtjHJ4GO3rOyeYncdCjcYWG/ORQuxNQo3D9AoXtrTkhD/jhqvVB4
KkkX+HjJIwr7tj/8qtwDwUxJLpIUkNxf60y4UMKNFSgif0ReaYOlvl1BSUeq
AhUodXWACSGLaEjEzMWSpk1gUQ8MNahryxcsgkIg5MpkP64aVt4VyjpqvTbj
OQL5uwLenvFIE+tspeneadrY+FMlmji0tFY6FQByD2tRmSGG7Z/vTSU6gjrZ
jCSQwXTS9dbiCp5bKyYkD17mcz+PMIFDAmM4/4ZArSbOn0EKVz+7Ml/PAXam
4WmKIc+D0yWvIJCPx26l4CAjFLSNgOOcOlzMuTDJ4XYQZlFLLUN6XU5GGm84
oLP+dJ2bb3s9rPPaFuBp4CBmNWjXQNXCgQEm6H//mX6Ir57//PrOOkd2JNa9
vFRDTRU1MEBtAQunhoE3UPJcfN37+S61FG2XjpPkbiqnHXFdaVlLvf/Prue6
2JNUOVfkg8ZjyUHr4kfLnIzDRMqe/1wKGR8+t4ewFZbUk78QHVvnsBtYEDiW
9CpTUNVvcgAMX+A7QeRJFkQe08MIkzSTqS2FCx5pw7hpTqTUDZZv0cNZ7Jtt
jGgYaMlvqFf9ItwU5TCzqP0AP9UjMOAqB7CJNZVUnkuBSlVW/wBqulAZ5iSG
ewAjxZz2gKijTw8RL6/pYBBsB5isxS3nD1NFd2BAKILGtbZUle+Df1XG/M6h
eYOXPtFF0YtojD8OO/eXcBZ+NoUbNfI21vs43o+Jx2pVoEQdNJ7IMZJ85jFg
xvGa5kDd5+wyWN+jz+cKh0l6zkc6qm5Ra/JB30NxKLWJKAS70l0y4V4gH3yN
IVZ26O0a6wL+MQR4ZiFzFGU7bZC3kYGUxQPSN2oxC90j7SEQtVh0yA7VS1P3
sVCUJqAPyp0Dpb09GkZwQQyQ8B/fYyXGGgauvfPctfbXpZabr9FIqDd130Dj
ejZmoP/QtIkUgOEDHi3RG7D5N8Br3EI31il1E8crVRNGbIwR3JeFFMrrQ8BF
AIkF4jQSr+6ZbmojWvxlLGGd6ebt3iKmjDKXuHN8or3HzSE4hnkRvf5QqJxW
hR8+GpZBiiBhcx/q9PYlUDEIUjYzS4KanvXZvlHIqJKLTTWE8dCwIQUePJTq
eM+LwRSXSLrZL4BFZBTzzW66MwzCZEfHb0GQhztHKsq5xO4mclXc+p9jsd8s
raDAU4IKFz5Z3e0LdqQK3jVMb0fgliOikLzw6RIdGUj26rxGwGQb+vjncV/R
I6Ui8QdApCAIIuOMoZVNOer1CIB9PP4fwDSZA0HJefZr8d1+JVVqqf1DHdrT
6bbncD2i1sztVXxg8bnWWRCrFCnUR++8I8z2iWU++FVWeGctzmwpyKO1ZkDc
Ce1sY4OjVHypao+1crTpiwbf0w94L+YJlTijA/xZTLmQ/S8Pk9TX3BjxBc7b
I/h89c1HqvczJO9YU6Slf3GywB2vk4OMnuUhGJi8tGhpfPXzBMp/aojioxNB
/Yfw8pqpH7rVzv6X+mfstfwEb0o1KNx1gdx2HkST7MWAwaoc/5+vWrfJ1VDK
G8dGDP34V4/TcdrxDPX9zXqUGDHdTXWHbDj+ivFdvuHu2iLuzM+p/gtY1L2m
oEKXwX1XSq0/Ym0fP40rH8+PQiab7Dhk+XZVWQt1uCx41UjkERUdE1POYHEL
NM9OlStFSY0fe7Bl9JDgVSQBDQk/nI7dak4BBxEKEdqBV9/Kw2vm5E4KL3ft
KNvgi3hjhp4Ru0z9hlJOepAiCIv0KJNiBipK/r1bSUTtPvHVUifbC4wil7Uy
/57Ljfu9v2BzwmqX14AU9DtLPk3KkjJQUVufQ5nlmCdUZdjFok2JXo5Vq02h
vsTInP0DGcz88iOOI5nKaW6xLNPzASWyxmGq2ZXOY/I6/cW+09qoxHYCsTfJ
k/GsSxq3Us+UBZYxVdFSCH39DtTnTv11Zst7KMOaF1gKv63hx0ti6vgKWnq4
q7yxQ/HlctalYDmrBAg9wG4OzqFeW+D+yTKleRmdecqKTnoo0JzgrWiJj5Gr
z1aRRVsFzH3YFsPAGr3g4jyQQDga6lTKUhqrjeD1qoe5MfaGYoqxbzwz3ku+
VhP5RFAWRCPMVx/fXbBVQLKF2UISviivjgAPHu7o6N05jbJ4bFCgPg3tyZE5
Mv+3AcxSZGCJ4WkpWcahFbPz34NhK5uyCyoS0FgfMGLr2YFc/rzXFlFNLjK1
SuURMyqlSbV8nCASZtUms1T4oBG7gqNjSVaddijZbSQkRt4thnb34BQeUTHs
NBoSOb2q2JK4QYRrEbdinkhsrzSXslOjImRNNK5wZs74grSoCDM/30Kz0crG
LwOWd2szJz0WipZCjBcNfB7+QV9o6yL7ycc6YiZYysgsBYVRZGDQSRJ64zqo
A7cpVQrkPba34H7WiXw0dhegzei0CeihcwaXvT8jq0nL1mh2YauZZKXuus86
Cbhyl5Ok/SG6wrZao6Zs6LTcmLaeYJmqcj1Zw3Q+NvpfZWhH/EqBjHED+sav
P3VYkbOK8WwvBGSigke89/xrM+tJfCqmnHW6fBfFcz4CENRKZSlR0Die20PD
4dpffwankOQRUxFU85V5oMvQUdF0wL1DCJpRbgA3uTlrCGRuRlh10Aglgisv
fl2mHAxBAdwy2Zdz/RFpAkNRxD6HSUkoF3D5gEnuS7jKizf2nida0TToJXNO
dosrt7X9Rtlc3NIwJdddddmnTL3c2jpIOiXQy0OqnVrUMqUskO4U1RONBD2V
7I2MxTCi0lUZMS1a9++LrodHD+fKzyHvBQ4DHymJjL64q2cuOm8WwDJGS9vf
prlI7OzOECrBK/vaACxmja3ClZXA67PJmvlAtKCTTdPV1IE2XJjRxUNLSXjN
JA/xEbLs5tcGeAr1un/G0djAOKd1j6xgfuUnJ6zKoB9nutWX4y2ebh8EcfZe
2JtKf+BXqGJivzmz27Cy8zFMzcaV+fJpr9nxdaCf2xiMF15d7jMfEFoT8q8L
dQhbLsAD1J4ZCC3VGX+URlvg2bNF4GW1lDfUdNDUrlN+/XgJBhLIGQZ53jwK
JnWQNbaIfkNX5ujOcR8Tb+NsDEfDCmiPyfJZEdS4Jes0w28UgW1cA0s844vM
nKX2ma36o6CQo4mUa/NVIVb9rCodtivCYbQFiRfA3PWFtneftMeGnz7q92nd
55DTSzMsQXugEntQdTXtyrAP+iRszrW9nxoIXqCoErcngJN1dB6MzgjUrmUl
KiKOtGhKW7R7bd3+PKyg1uhHcU1BoK0G1hsStF8FdzkYShISkWQgK+/+3m07
aoWRjU2Pzts8GGNvzZ0ikavL1UzSOnchZJ47S1ZY78/cWPycr2PUUkY3WF2+
Z8zSP5GHYNhgU4rhcd6eTYdHQo4IgOA9G4gJQ6kU2mUn3YRc8joY+4Nahy1d
gLaDvWaOm8KVWtL6NnXEb85RE/6j7inOMdUOHOvSv3LUPFYSClfnzH01zWa2
OMv36VCnOx7gbz69UN7+QJ2Ze0Dtn+oPdYKWedi/FOF6wnUpxMKvOikYKdxA
cPsqRId6E6Td+OcFt/9OnGFxIz33YCE9ALVepiyHeJ+qW17+Ws+0HFOyUy9e
5QiVVPcH0kkBx17uVo/NWHSMsJt/jArYXjugSuumMw2lwBOy6OjAMop3ETAS
BKso6MEREFr9JYNqtHdJDKXY6Ec5kZOYDdQqUHU3amyKQ+42iAe3Q48bgBPB
Pgkz4zeK0zPMD9m654C9/bUQNVm6GGZnTXX7KUsckROX5RO7+7SgfquUhvo2
AqQY2H5krt3/QCP2EbbxzP4JgzV/ha9my7uDySdvn1OK69PbidFVDqv9p375
dgwdI4kSSIdxh5FwZ8zugWCf6ID7whJk+x+JGbyDfXSM/GXTuj3M3XEGD+cV
YWyFPtzvJWbzIgxN+SLCYWW+ZmpKDQOyhMk32UlYf7qSoBWGsQVmu23GeD1k
+nzinCimh3N+HpM+bCATWbaj3kVaobvzk+qvbSjwRILysSf1cC3QWMb9Dz96
gni40fB+wqGda2RviYK/mEYTnhNfrTh74ixIpz0hE1W/YqYI01kF0Mlnrt0q
U/QzMnXse+Sj2NMficAxNGPe40vMpC4QK7Sv+RBzvSVJTDGS1Sj5NIkk8/Xh
JLXfs+e7b9TcHye1AaMZzAB1UnLBDLLyPph7oPnf09qO7r1+V0PDERB2okHy
U5Ckk3gYiP9kppmdkNwYpaUW9a3JMJJmmx/E6VpMHd2p/Wyp51bDvqCiX7W8
5hmU6jAVuBw5icjvPh0aocmA4zzr2ooFm/448/NqBSQaF2u65+nE6maCze2g
md3ZzHtrGBsPWm+GMmIxIYDjC0oJPlkfV6gWAspqoH6Kd/w+eJhCiVRaETio
ahKIrcAIc4+P4dGDM3Be4ylIQXFsu3vgfsniv+EmOdU6lLi5aiZGRhwoBspG
D0sK1HT5EgYsMvkUTD0EXYNkEBvC+yiAfmE3mSLF53gRFkYtrt27dxodGC19
09cXhWTSZ6kGM5UbOYRODLjvt1X5I1M+E9BQeq7vZH7ZcZYTTiiFu1qNnxCZ
N2hjcA8g9PihuLRayeyLgML5PdrMOPrutyihKBBcZpB0uP7cs8tFKsx+7yRl
lp4KgXRKfgxxqjJkLGWu5J3L9nyBNgMZ7DY6bY89KRETbpkW+KjHNgd0Gf6p
MT5gARUE9mbb/NjaqprQfcwVc02U7iJ/kOlWJziZdy3+qc+FwhpB4IKjPXl3
fHxRl+cUls7Ummjp/Ydvk20o9gW5Yjc8IXBGyWspag8Kxdb7WCpDwlpCdZF6
1KdgE1uwIY8UIYrkFepPR5LIib5eOd7dvWkFsO9Mortb0cyrmj/gAEA66cSp
SxrE+wyfeMVc9dF1S+Y0RpnyXLj8q6SU5+Il0eGFMdfzrLrTLFvTNqTAUH8+
xYj5x9LEQ+ik7lMOD6NNWSEsowRAlQl8MOgoqetlY8p/SpB4NW6v4hVDp3fu
lrlYi23Y7uViBdZjqCb5qR+N59UbPP4hxf3c7U1iHYhDEjJTzPVD5+pbqIxv
Umwmw32JYcHUpf59W0zM651UV7rp+kQkXm5KbIhqnC18fVojYmSUd2goO3Rt
0onNe/+95UynnroV7mCgOMuk5YRJdzXz+LNgIQkK2CqlzGnVMMYS2jXvUsEz
XK1q7nlZVjgQaE7NfRV5VOZLhxHF0FbNGZUuPNCK8BusmrGp+BH7nv8iDxwr
qwvw3snLg4/SWAiBE0+CS0LmTjU3OgZuRg58JcoiPvZZZUx2MhPSt8lFdJ2F
XzTjWunIrepLRn3P/dYh0Ac43FT4j1+sfeOZdGSMf1vGIBprJbsxQbpmesIn
9SB1+u7wmt176C7whFgywHc8XG/PKX0SsAjFNaziabCUJyPCmtDjQMzWWsJs
TkkTiWhDnX2SwLnVJsneXQUgtFqaxs+46CXCnxUI46zQoNCLAoASnRMl8Zwi
U1XzCWav/iThk/ykiqQj0FyKmGLW8iNRffFNJQqC9BIiccLbgVSnjYxQ84iz
DiiGzjrxyH+Nqtjv9e00UJegdpmPUu08vlE0NLhK1uKm2Vb5rMiiabFO8SOs
oYzfQnr51q+bk/noasP7+uqRM45u58Q0V+5GgM0Zyo0Tz8hR/kkFyxdnShMB
LEPq8Y8maymPFHgNOfH4ZTAxEu1wruhiE0m2NbDvR0mi2TVu+XIU+2V/jrKW
LUCZwp8NVGadKnNdsZrOzY3oWxXouD3BYCKmJr67/0EwmdozQRP03nucnjOy
nGRhoJKnEXIL0efu3cQ2dTpbJl8nfH/O/BvpleKVJn7cwxiycpWJU4ty7lht
LkhrmhHTMUxhnz+zaSeCfJ9JTdVRTWgTPL4tiPimPXYi88uUDUAUkL3Ut/MP
vRIwjvXi9G4Rva3/LM3AEVdTKI/CibA3PUQampkOx3bETk8DswNps5iPPfQI
gyVaJbaT/NcS4caCIwI7TqA+Mb7pgKygamVRYQokLwO3ls5FDaNwYaalaJXl
7+OEdkDnwEXNmIiDb5Wh6KNeR8mNYsf5OE2AACjqbQNSC2mwLBMphppRHoCW
Ki0RFNnHGHch0I60k5vv4MTOzHjah6nlCHkUfKaM38AwiZPRE/87M3Y5RlX3
0JCfFPl9USmnBi1t8UTPBQEr7g4M1ibpiBIxTi6/ohCc31NHr9YpZvPfruks
Vw6YmjL0v88TNszWkNbqFTmuglh7b3Q7Fdo6x65wooPYM6pI3Lrx8NCstURp
5nGrH2Q7sfJ9NTMpiRguur64CymIBbXtqmt0GBxHck0Ql/hLLNfYiN2PZeJC
wBaMg4YZ+QmHJb4iGujYpDNa0hebeaFcoU6ydFpAEAlW/RU/e0Yr3ZAHDPRK
j4B8jSK37ngI+vyZrDlA8nRpS9vS0CCJVwMz/QLr+u2ZP9ArFPXfqFOp+c5H
sBlejZo9R1tD/zoEWJuWrtQKhw6atyTEBiW9nKqR7gZwVrWaIBVxpmTXzvUW
0HbkTj4s0vvCpf+kF7+UFC8tGdvsHpwK2/yFYW0Oe8A/km/bC0Wp188TEeqd
SXjr7y+sXETQp3GoDkwil1ljCkSUJErR2lwIJjuuk7YR6yAzv11bgGfduDyH
mR3IoEEZ9c3dE8qSCC9qISTXXsIjY1uSOlxfYaj0pjO5tRzNnsHtsJcN7vwt
A8Oi0aSiP1Kz1ZgBOYxeqxR7WCJKiz5euqif+Sg3+VBRA/VIfKqkU+L+iKlq
I3EFk/MouPcCwFyPy1OtUx1ZgQoC0M0xGKHIyAPTtTJuU4yAYCvUVDRiyDtL
e+tmpv01rLMb0g34UdZkuBxCWKPwk4Efq9FzWmMsYHaGSQmjBQCOl7HgUBG+
nJLHyhCsrw4woBfYmMoay9ioXQeDBpBV4qtQE2FgEIV2zGyIWpsmWoldntpm
FbY23NYmMStp7csL83Fl+QXvZPPc0gfoe0vtZR/ovK/z38NP3neOv4ayVOas
mz6dkz8FPwp/c56B/gI4pnIfvuf3lPsYz7uPDZU9JXWKs3Fb7H4eU0BKjUkw
Yd/lPUUv7uLVrX6XI3OkUwjxveDF8O7g/9EtgV/3eUOALMity/JMGtigg2Im
YdIaa0V0NaL6YfzoSFQbDk8SkQoMZE7pWdNAr0Xf/ljopK38x4sZOF3mvcDQ
3+RsWVgpGnfQfbuaYmNDy9z14AE6A/mOZmzGhRfk1bUfWakY3J8AOh6Gjw5k
BkgB98Gxn+Fwjq/h79Yy+XMlQFsTMm9V1kMBkhXfW+woDNRRrY2AOOyjCUuD
DchE9hg3j9wrSu2jzjhKyz1+4oVjBxj4UiZmJPZqT/fHGdfTwZ1URqrgqsXn
93MRUiF4+XVWacTGTVESJoSuRiARgt+1wDyilGpp2V/o7iszuQTJ0CAJtIsA
lNY966G9A1omG1CqYFPq7PM5FDv1XvWk+UCjkpFhGeaRzklTE/YbW8fPpIWi
t7WDXSNVYeixUWWSSAoP4FPHvZROjMIBVbQB6mpSZkf4/BI0ScGOs2aZNpBS
wsQSpWsWAR0qi81ZKeVPrN2yXae4uEvsbSnIsh0gfQN2g9E9njO9UEB0t46q
1kxrM57wQ2TjJ5mcRyDWDxUIu1sLrohvmI9GC8aYFTC3RR9OsexS7M0UXvF+
kjteOzo61QEII+0zE8uiiURcz6sgw9jNWaex7yryiLnjPKsQe3KtDpfXWaHm
KCZkYx+CoLVUvsQf3TyffWbhuDjlU4pi8Te4g/ImmfGk38NIgQ26stIqVfGg
G2KkhqR3xUhz3AKyGFm2OnVOBoeUqAgWy0/csz/VPEJVSeUld9rMJH7cH7QS
UtAVmfFQGv/mCNJWuy2IydilWwWur3QPOU4sS69pSvDwZFOYXvCb5JDRgZyr
c46PuMKOU/J+hXmAuT/nfIinrMK38E5WYkDbFMi6i86Ct9puSrAPmUTVZW/9
JYanxwwO5hSoQBPBSLH+gDlxLMdL+J7Eja6KCKeFcCcmRNNdy5NRE4+q90gB
Qnp2DDoluXek11p71P/dK22Y9eRBxB2T4JhsFHHgOzLAyljS5aNuPOI+b3X6
BUx6ppei2PoW6clfifMu+EWVML30jFiXzl3o5bmi7jnt16RemXhjf5DQUcob
3QpYCxgj38XKxMb8R3f8tYVHluf9M2rBKgunHqzY1oCIe613//P2PJZVe04R
NpDwekmXYPCED/fqGcNiGdECxPwAz8gdmnCoKD7qFwHf29Rb56ARHjmuhaUx
rHmQyCNZLZHV/W6O2+l8wAS2Z9/NR+maQqnWqawAZW1RQr3BpjxjH2yCcYNU
1b1w4Ss4hvJnp63feF91v9DMvgZ2wn37FZMbWULdeRrlo1qcG6rt5oMB4aAa
2GK5+m4ni9tYP75iAAKp+714dIGbtOm/7Z7B+XZmPsAHEKQIW/QU+nxhCc4p
xblMeDfOj4a2vFJ/TuEXjXoDhXokPHITo9WnYbw5pqxLtYd9hVYnjbvZkgEL
7LPydsb1vfmWl8WNoU82FYS6dN8WbzmWlIh+4rQ6g4XRvZoqPE5vPppaeQPG
jhVtiRXn13kj2OtnH5e9/xUXbUbcI39j9BeiIHBh/ZdzWelsE8Hmemn3Z/QF
bPRKsb6vg1sdnYnEEdiNCSnTpf/i8d6jeMuR9EnAaeU1cgXA7Gb4TtiQi4Np
4zEhHC5WfrhjHgRf3kOrkNj62s7Q/d1zpKwq53tmlG/KO8T5OKY4gvIjCsml
aasKZxfu8QLDbAbOcDlgKjtgzAynvgd2wMT/eF7Tj3JnBWRlVsO3OfnUHjq8
JoqeyA+9V8KyFUrGrgGybnt25P8sZPd0qZ6BG9oSvnfCyYo7iA3TDGq8Y81y
3NHM9wd97DQru4G73defDGh5j9ct5vimg2GTvPdA+MFQUY+1BAco8C2SNaOH
S90dBLzHUAOqOv6dghYpGrwyXC0Zbky/xkMIDALK+bDh72E6ZgbWKlUyCvNP
FOZj02auwziz3sRD+ghB6OR1UfHvBBb3lEYLdlrrYreETwQzYTr51dgrCuXP
T6C56NiSzKmywie429nxloXDXFacZjltRCjMezHFs/ISvLbcQi/dzXf8wyhE
EwgusizRi7kGVeKaDTForzKnYVy3QXgw8wnSKTFhgDdDTEk2uK/cvSeoWpl1
4iYe+3Fr/YhHkB9CnQ2JoSViJMZOAgyp7KuspnItZcR1b3mnAr/HLFch3LS+
59lOVL2+/mgFlEWGslRIpAFavP1+ixpKWB+2MKcvZlxwfnTIK60CFtcavXhy
s4S9m9nIb7dFwfairMV+J54b6kVWkjyaFf1kRTdIgpGdBnfiUnuff+HYzSTB
bO1dXJ0Wa1SrJVhHMB0yQKBTzs/IqsllUmaenXyg8KIXbKQHTbBEbgq+YjyQ
y/CzQUO4DZru9fkL0tbS6uKy6mOx1B2Mb46QyVqpBqLkwOyASUBiK+Y3mu2e
LwgVXBv/oapnJ2ptg53BKOYd89ALj2MTcI3npJvwF13VQ82DJmGUgmfke67M
vu7sUhIBLmxHY4PJ/qPHH/qmXT3FN9hSus1GMTxL0vdZMV/CVK0/CYeGep5N
980JaMt72QFi60dhheBQ1K2fLycwlZknDIi67zA3JbZTlZ/zlmMAdBrPRs7s
QpPuD0+QLkbAS7V9QCecLtMneP0FD8w1c1WJjtSCKhyUaaRmFmDMC9kEBLEA
v5Mx6qiBZvihN34aSRwKSlXOHNU0i03Asm6QOUWZAcP9DuXFIu7UJWXjKNr2
bARiq9TcdHKXKT8QmM/4CB565RyiVdhoYRRnGNBYUb7dvmr+XkVbQ+Sur25J
wlewpWS4OdFQMGqXgl64us6M8rsuUcmW1iatpdmzlH9SBJx2Gn91k5ILACIa
Om/bi4YGtrWGjeeyMb5RtXd4mt0jCP2onMDM8ZuNHJy5esBw+atireVc+D6L
u11pooGCSKYqv0BZcxNPCXm5vNsa1uinOqNXVws1UyDn+RgQXzw2Rqhb7UuA
GWbmaibKmKgwdj66zh90CwUgt0qO6q1k7EADkoPwBB+usk06RbD0SlYHrydb
0hJe4fzJavNsUQWS/DXY7qopsFcisI4JnyM7bC8JJActY47rG+HYDEBfnyKA
EKqktkJznuXoWbm4WcWDNFRMO42nEHXE86CGFilk9/52mXPfRKAH+lSY2IrF
QKyA6kRYUSgomhA8FJphkMAipluiAp8Fv/9r9WeVdiqx+4oHQOtONhm4o02J
G+FhF7CwJXLZ296VCRuL5Jwo2UgMacfwyNWFZIydDTBJ6b+5Sfi3Kt4DUt8f
+plShOS/N6URa386va9xIbw4D5kAvYCHccT7kqLnix2aECtQC506o+vt4hkE
K5qqxC23EEKqBU51bIwQNMdxSW6Py3PL4PBW3QHRcYSVJHD0XG/a+3a4as8f
G09ue3QgSIsraH8XXjC/Frxe2N8qLbN5RvtvReAYyRVc8+PgVqMeGV4UHzVZ
TKEG7Rb7z7nCG2CZMQxeKFPVvsW6lCZ8RZiK+ioKJq5k44ziF2PDr+PK7YLW
nCzfuGp6CmSaIqngbHwR1SPz9RS6GoOHVUP8PL8a84S7NRZqVuYcCB9OXm2r
hp9J9O15NIT94NKfVgccBmiF9AkHjbcOrBay9wiKrHnGx+Ok6aPAU1h+YnNb
3bH8gciAi2fPXGReZ6+m8iAK4PakvDMgAwLrI1XbGia21iJlpmhnT0HKiUOV
lseAg1lc/ZfiiHRWU/JXxx8PWOZBxP6dUR6ceUIaUoOwm6xDIQPG026IwSDW
YuA4KrxAO1em2owtRe69LPLeTKwDvuQUMn3pS1plvu/Hz65ncj8CaA+LBzPw
HCGhD/djDoYU0ryU1n3oSMcxQyJHZywr+ErtaYMpVUSywKjpaPj7G1Wx5cD1
7U1F6Qsi1meEZRoeexciABy2wrG2cNEjoexhtX4Vb2DKPk+ummu1NDGA5p+H
McWnoUeoM/PVmN+Arv5LL/OOtCukzJAW8YSqkaiVd+FwwXjXINWIpe5yRCa9
oI8wNFNL8e6XE0111GZtw5AbiNA+3zGjUAr6bDZHEt3ejfCVSVO/psfXAUju
uaoS7LqJ3sJNWSDjE8jui8LfqRnpQpeC9E6osHDQclDdD23M3c3JIBXezKPQ
cARYDb4VlhqRkOkCIu2nKFm5Er46RwsxhD47nIu+pwDwL8q4zpdYpsEuJXuJ
dVD2Kc1gamlY1qDrzTbfAfrgV1r3LdCx5jDDE6e4YHjD7psakSEQLLLSYko7
dXvUrVel14T363TK+fWkhM84lE04NawAkO1ROrWZxi7sT2IbJYwNdLtvjB64
u3XzuC8PpSyQwsi7YBHCPnNzDspWa+K80amlkjCmMW9F+dpR+Bn6C13xfAa8
Bt8ajpEt+JIcyTGLJxcF5oUIFtmvkNM0y9H1SN9Jdkwsaoh5mgX6om0c3HEQ
rUzEEQ6JU6yn73gDbFa0rGQ3z6oheaqJejyX/jeSTcJidYaXPXDXqJJywUdX
uZXnSq/eLWQIWP8+lhhD27uO+qH36eaMnvSWPnvXd4m257dDQnm6v3GfWVg9
bqHicd7ZBbm9HZuQLQRiyHm5OZQTFMpu+VA3FHVdfQTATH2wEZojXct+HceM
A1YhUpdBbCkXUQ/4h9Rd8cjXqr0cNPtiQrervXRgjNOB8eyL2VRHWry6CsYv
RJq6xrQSCenF82+QcA1kkrxdIg7zZINdWnEy7VNZzI99VGDTPAIxA0SP/S5p
LDV2dJrOhJRdTHezecD/ydiRDST2FJ/sbZjleeVhm4YioQl0DBAzSORmTv/j
nbyN/y1X5+7rZJPe6t12pI4/zGb/tlC4OiDLr7A5gX++HAWWP/VIBSI8I+ty
nTv8geDHa/IVVjqcxFHuzMA0zKd2ZIqxHvxtkUCNHNYeuHj7pO8/ueDleDb5
LmKZf7Kph3dgpx7VyoMG3In6qO0fyJT+QB5SrVXOhZhG7/U5SKejL/pIwz0o
lA/Pzzqd+q2qrYXgLk50NdjQhyb0Wn2f560Bd/iV9I24V2pvYFauHZ+1oL3J
J1uYDKgMYxs5Lx8K8M+EldlRt5GDhsr68kmGNgsGjsD7t20Djqa1XHW+KYvL
ILuw0X5+e6uXXvhLyWJXWIxhZG/A3fEkXoXhZg1nVe99ycRrAfEUvWB+3dNh
5i+kIWloc9+nvm9pVjwSb8aQ1tBCqyLwp0JVk/r6A99VglGDKi3B+IPcM8bQ
ljexmnOB/pPM0zpkT/L4u7H8IaF1Zlw2CqM00hdypW8W6o8WIFAg5ztktrI2
I2IhV0kf9at+3YNhgJ8iYNMC7dJ/SgREBHnvaOFMXvMahkGR2KY3s0sVj8De
1X19y9UqJ27jV0DzSdXF+zX4mae22l7J8Sl+Ih8psjHaZWpXXDc8dD/XbUMF
/no1U+ciSpThslKGvA9neoUblzaFOKvvObWxrwGXVixrsRbBgVVkPWQ/VL+x
qvsjEHZ5KbHygHrAVcY109XSX5i+b+yJTSkfO00TwriuUtkfIdn6tFYhqwz+
eQR8OTCkQeiXVKMPX17T6EkZwSbuWHbzNgL4HiwsT2JhidrW2kFrKjmvDbzr
8E99qRoB3qXup0+e0F5+oMs3ntb8TEio0mW0RRvKlvjn4VUj2ahmzqCKN8Uh
16THXhrIL1mnt777UumLaqrSV/R/Eerxr2pWgcwhATu1Tt+BFURzLy/s3Iwc
ImjQu6E/BhOQ0t1NmI1hCywCTJ/xEvuaUIFMfb+Bkm98ZBwamOb+fJbooAov
T9PNxbAcMg/7shfOSHsTIpHo86NrHIIdxk9i1+B677kY20X5WKAYuuE9kDnz
VWxxuwt/qJLpkVPyen2NpEsHC81eLd+ax2y7MmYVv1ZUaGjCVah7j3p3/ymH
+XhTYV2VafIAzVrciPlOyDZ6GvCQAj5k/qsW0G6qxNkaPyo8gEMZdpIv3W6q
1Up5pKWXsFFjvrw3fdLjZsxWboRZuf6pOlI8KUUHXED4gvsSuiG3WXq4eGcW
LwjxhMu8Q8EmXavOUdUH5KKIXkbmkLgDzDra7CmwKbUCM+diXQaReJNI5sZY
9HHtwOTe7Xq1VYBwmY47VsICSJC2NgZ/EkSIBUg+5muQaA1xa5WtG+KZB+UK
RjcDoATGacB9L0r9G6LIfEXJrwxLvwcv/qy0opQ45F/FL6sW6RUDAT4cG8z/
LFopWpyYTsXCF0UVVlY3ACNMowO6Zqe9zJ58egmO5wdSY2Ckg3UVtVxhZa6G
nqzgnBdzrPPysyf+B/Bg/obZxbw/XTZi1DXtu02dDFUbjiRCfK6j66s27czX
HxVicDyKUqwZGTyU0OKCxdIZ3ebR9q0r+B54sEBcuafvRY3hCjjnHSxDvqYo
g+6D9nJnOptnm9QlECo0eDxLvwEllpYDtjQfGkbV5aRVE7KPlyHbeMAG9WOg
K+h8OPsJfsPu+k3vaE9egnEgEHeF2lCavqBIpw0UE4KNo86eIwvyYZWqAyWK
4tw7GkNL5VvqRjFrgn+XTJWzJ61S2ypKpViwMk/aRtLD2Gh9rbLuEnpDWfFq
oBCBTnZq8qfHPZPhbx/O/9EzHu7HLVrK7SMJxwLiCNKjblZ9Pdu9jJosw2oY
EQuG6lCiZ4TLEzTK53I5lZ+gBYXZGHTCZunLFveJqqyOP3dc74qcWYz0nVr7
0Utv3ABUWPB5nOeaOEl0JtCFm982oYW5S95ngzkh0tVO0gq6Ok/ZqTIFUWIm
tqAeqQgiCDKsF4CX2++bleZ4CmzxNN4UbAixl8aPWKzq9w+RzGnM4Z5/jJ1H
z37VimcvaRxJhPNNqA/JrTrCSw9xRSHHXxVIooJNoSrwK2spGe1RrgkSRdqN
QZyh9PVtVaxqfgPywAzkm3mVjHAJaR+HFkA4yjUMVMUONh9xpeVVaFSMCNKv
YsjUulPjjIauYABIGLS7G51zd6GjBrFaAMZjhBh6iD3HAvxeo7LP830UTxaV
NVPf1r4uoos5nn9UKMBArJbyOF1Xo7MiAfpcOKkciALHy8hcoa0Cpgtlgyo0
5UoapP7kdiV5Xh6HFMoz2FnNHYSrxjTxB0Losj7mRa4o3g61ba7fOvuBOhBW
tU+TRqgsacOyMYEzO7yGN4PrPn8i5kd8t30SJNaAhyzx3xOyLW5ZWh/KtvgW
IwcaTsjXejId4y+9D6pAk6GKyKfaU3d+Wg//p5SuT8wRObZiu9vO0C9X6FHp
5+loYZ/tcIrrij93kAIxrqpfsRLgVdQAaqDMare1VIrd/vnkgKDX0Sfx0Dwz
08BtXfX/UE5ase+hpNNUwYaSpNViv4QQoSjTk5Cg+85HgrjSo00KPFTmT1cW
mW03In0lDgsQ02GHNkFAbBwvDDL3+jF4iGa2ijMORftQ595y2+yVdmjCYJjx
x/zaIHG7QRr9nLCGvlunIDcjk4sJKWVr7VvWQdZx0rEPnk1qBJQ7nN/SdUrk
9FPTYCGYR3OVDlmCuoN3w6IMvlUn766G/lhvzMll2yGYySCOCYTEJpHS8RuN
9kkf3Fvtt+IwzlGRXA+HiJSQnPpbg37HLtfGYIoWN5nmuRy//V7pjAb/X94N
x5DcPCGDOu5DzjtLwCq3IgoSWFJoL/VpLZD2NBPNKCg97lzBMCO54VKp3y8W
k1z91IqLgdADi9+TtoSPRVsqw76ce9inM/GabXe6MfEzb4KnUDERV/IUsaBr
jGyZRobfi+DDFwTsbA+eqFQWxGsdbakcn3tbXkTKHxUiwdMCy2Sha8e3+Txg
ckFn1KEG24W2X+0Q1CyZUIBVnCpIGsunBy5VPWi1SUomFSw8D90L7hrw6FwS
Y2SDwiKfyLXDZOX8dFujn97B13z5gP7PpmF+9SXdgKeA1BtCQvk5TrIbpIn5
ZN9lZ6/mO+VkdAJ08OQIu0atuigf/+ZGHrPXr0QrhNegLiJh3aOkYuePukmO
Hu9YdfYyPweKD/HwYE21KtTTW0Rc+qAbClxk6HyohghQ9Mc50e+luQTZEr5j
cjesKa9I38e+R/e2RrTLKJ1G8JgyEOysZ57Qhzclo6U7QPiLmByofWkNqftS
0iIxShqCuJJ/dVPx1Rs3sV5mam/fJGS1e+Y6cTrSk2rkeHM8wQ15gYroqgeF
vsBkAIfZ24Q/W9n4/Yy24NTSphwFCkPnlxehpBpaVNznY4/SgE9y4W8nEv1C
D+R8MMtFZMY6M1jnZ3Lv0IXuett1GvLpykiCeA0eJedKidZW7/enf7cjJYkN
uFe7LhdSXW3LMc/VjJUb10A6+24EipgKaj4Owh+cLyDyrF73CdfsXZWUk2Wz
Q5hSEGnk4JPdlkkLFZIyTahbWZWKL3rwQjucTOz/ZkKZ+EExlLjSMOoCMhlw
DBiAH2vebnWaTdPdtLfw9YI6RRx4YX4bqRPRhj8NaXAIgm3k5OzSvMkz582j
E9qCEVRGCePOPe581UMaZVF83TXC1oPyRU+9qfGkXbNwyTjabj1NiR8m9hiW
2bwRPZ+wT3fIrzW+frZ5Uhgr5lGFNCMaqzkuVB3E5Wp3YBS7ivlUf0+5OSg/
vNo8ejD5ddeVv3uXA/vbzqNnG4oBiUxwem1NFhgWZ/xN/zT41syvskBqqYE/
+LidhmNFTn7Grh66ndMwiEYmGwcXa2zDmp/CWpTC1wyy9uJmSiQUM0eYWzsR
qiXv5WMSnc7yUFNIsF5TXtgTrXFY0yxAIqD75goB95RSrxvSl5N1BW2X9rwp
RtMuwacyB/QPdB5cAVt9PqKObEE3TVipxclmQl34b9kqemYLOSwVpiQ0x4bj
NxKWeZiNNylKdhI5aYmvOycGFilw2bIvub2HUm686UrGQGH4z8sYd6QKbyu/
5ZyyAzB3ZKQj19CP8GFQHZY5thnlfyiof0HfSwGUQqG/a9yjaq949D9LJAoY
0l5o1nJgp/eY3NBegDf521LrcGgC0GSelfl9NehgHBnNgGz3bkWK/RUZ76cu
iia8Os6PlsvzGfjkZIytGdazk3GF+Ug4pQMUqRPgdiw/EwmlUm3RhiD/BCX2
B10D2o2gIDX5r7BEzhw0LXddEzi2wFIj5sQtqpckvZYNwdZnALVzNDxXF7rR
I/vP0Jyb8LZimouuHGr+0jCFoh7mwfdU9tpmCprr018WdIAUOe9YDZnX5xiX
0n3n8zHViN9+vaeD++qyDnyG5A2H8DM0BNU+54UhSh1dZgD5TT3cGy52d3MR
qSGfEuPvp/0VPA+7vavwE5KjeyI3q6SAZ9mCdy9PWjRv5g3bVvlUqANW80r9
S6buemeT5rv6+LVuXR8flALK9vC3HLwpqpjVdhsymBOKTkhyigZTn3Mv6tPy
oMXNzWxj6WGh5oEYhHl4CUXY4n9oMnLQ7H2Li9I3FonctswFp2yK+FIuZmOK
oH8FR41i33pijKPVq7VXDYkQX1GpZsR9tbkJt1ompSMnkxyoDo4ML4qE4hdz
6WYSFFCeyGhBInTIZDLl9SJRZxEyIDwci9Ze5Nj1y/gkXULkABMhWRhMWGw/
DoDy5IVRuSVGqujfQPbrlVb3gIZ0a/Bme0QtnfKp7FeQW7josQiQcmzBEfdY
Qk+LBMYpunR1Ro3tpKrD/sdyWOKUzTooB7JbMfyRZQtyBET2/H8K/9mJnWUj
7u1FJHnaUFbbgvhd7dppjWrfDdnr8A5Zjjv5xBB6uLacyl3VM7fI40vyhwD6
rVvmSwzJ7ngoOvWWbHYdCezF/UcCX9Mcfgt9UlqVukfQ/5TSWRe14qWmT/z6
CxE7pIJd9fjuAryOAoyanS8C9PvAP8mGP7ewaGWQ03lOtLnl4NALndgWvGsf
yMgGDlj5DyCNHVpoamqiLYD8axLIwjlRQrsbs5rLq4k1Yv1GdNcjnQ+9RcEA
jBIAm2ZsegTQ+fgm/0tkZmbl9KfYmP3oUF8MrwMI7n2Yw9+KA3u5TOyXl9eg
K8GNGuWV0aWzedplwZdjkEtmkDJ8Z1sssdn0IEVehp4loD4/RN25rdPf0Ide
fs4jSNMZj1kEyh0RQ+3VQ7Rdg1irCm97y+4WVSpgAfCP7eBB+HiDG/9AsOPO
jBAhklcI+IzUgJpSonPNNqbUYpq4RuVoX7fqcVWhzuNUr2ycjGzNzy8F9LSm
NON45Ii2L0gvXPiBNYLl3Dd0rhJ8P2CKjgtL5Gx5kd8xN1A5vH1cgwjRylUp
axQnS+m+4cpizI/Y2PHzPLEwhJ4WNNzsjC/YpurtDZz+yqXnUk9LlVnPagbr
S4bc5yjX9J5TOn3YALjEXm5WSCBgOCq8YvfZcWtaJ8E88+e9JOTkFs/LTlIY
Q4eedD31Q4/S3Cf9BqKJCU2iykrD/Bn5Z6yd1WIISgTtv7ovh5iVLR40Ihec
W0x6lqY3wHDbVKroFk5hn4mRDLJcH2z2ZDv1Cbn/FXedvmk6WCk2xMYmee9b
bGi6UKq28JByvQsEqp2j+y7GhrSV50M/f+jvvDz3P7PVwc32zTuoqOytF8X9
6oJ/GSoaIJw+clrPqcpgJNM1qscdpqlb3jJlMfy/UXW4KQ05gJtKmHoSQXFG
o63vtwiNAXmNnf4ijwwhkQ5n9eEk99XRomw/ACRxfffBKay1Ichck08ZVKwf
xc70EyB2lEKMLqttB4jz0RkAsETsRouP2AGIGKkUDDRGCcb22NWeP0i0u/4+
ItaMEFfnvicZPw6CESWHpdYTQADIywcT8iMG4Zy99HtcjE1YmQI0t9pXNYuL
AORrhWAbJc0mfGXVvyqjiHX41+BIop1hN/Qb2H/9JAyPxhPJmdD5xupNDyE6
e/mfxiJb6L9McOtuK4hlX5jIzS1sy4R9maOAz3YhP358nLOTFXL+wW38ZULw
4okqKyE022l98JFDCREGHXYm0aWDuRKKdYFsv7taEH/VNPS2cHuXyF7ZOfRh
sPhTfzO4ryPNc0N4bjUJQw7Shu7AQ1164R/n4kW9nGqbGCLDH8J+vBqYyekM
5EJmCvCq6w3OQnksMtBgUZydSfiV6R3gLNrNTJlH9TMaWu2JQPVSkpoScTeq
xO98qMPa3VDVTrPXvdQg0QBNOE+rGwpJESSZxrIhkzPqLpRFJjFc+VUmRxZ+
0UUjkH/fSYz+YXRkOHY/L5uuJJL/0JhnsTaCv/anUMfQ0PVQO9hC6EbAaNLW
O4tqvFwteJw+67sNIwentSMIOZiQ41O0LiKYKoaaCfasVDNlUTAS1H605ib9
dwVxXQcueKvQx1eUHIJFwJpjJMDfShnqtyGdOPehtTBVeL2f3FQbpk9DZWuX
nvq6V1JbtJuW5GpiR8uut8DUrmbYe/j3LY/Nk8VYLNg9xKnZ+ryjtTVkxBdr
ip+q4jdUN7HHE+bOH3khs1CQQO/kCt5vJ173XZlSHTlhCLStPRUBSvuAkE+X
MJ0IureIjH5CuN3R0rWsptaSgCWiod2l9KBuRAq3koZQLqzKLrKcsoCqMvpA
eo2VzzsfzQ0eBziv/w0Ga1kOZAxaFjzXmzIviXU+zPEzF150TPNsa2TZOwdk
brA42dqNtwXi0L3ZOS9JZUV7SRtOnz4T4zUNufolla4k4uUIlJVXMPMYDDDG
lTCdH5kAYw8BDLwqNdwyOPs8A1Ztw7ibvBndk86eyFEiiqi0CwRBdZEliM35
ab+91jr7MgKOhKuP/wyXuJvmT3xNZUMI03LuYh5t45Om1UegjRsAsPjoSLcU
ztVIjCXm5fUl6/yKRZH/34Fzx0NfCmyHo+qmUbQBIz9+bQyai6f0mc6+2oJ2
6eY/t982dW0tbKHgVxzR6nE3sG6t7be2/ZphyfjpJ/ECwk6arifoupqPpPUy
PrH7FM44O0Dz3zenP6U0fMjIvvv/GOiDTMoNcEjYEvOsBZo/POoz/gp9pa8A
VsNb0twI+Y6ubCGwraCrQCbt1avSC5wLzTdInNuUnYvxfsM6NqFkzgik5UiU
8lY6eXI/cDam3Q/Kbdh9lDhe2a134OUFznNiTTkf0YD0ysy3e9xgZCbipl77
4t64MPJ5hqrxnfl7fko/FAx7LimvG+1Q5gXkH32MR60ea1kn0eOfGU6FZmWu
t9EvJOw3v+jYyT3MeUgqtQ9kkJjkDQdV+H+RZWdPDF1yr1/TBMgPPoDqcOnB
WklC6OUjysG94QHnTOoqN68chcyi25+X5p7hJyA0w9DBAUxoQTeayixF/3HL
9M9f1bcQKSldYyReoPRJ+fjXyB5SfcbCiJXla4TJEp7w7C4sbWVFhwLuzz50
BOHPQNelyqyN0rTL/h8EjOvLFIlVDp8UkarBMsvigbzteuitEsBMEwbsdbuC
zLErxlR6FykONXfyQLLfIuG5fsG6BP7SgGMI4YOAqcccyAx8cSUY4KSE00+p
zSIFpJJefd7sgY+WOpFLRy6DDXFie6ppm7aJSlIebO6wUutqaLP0v1X4xDGS
oPOADlLTW7H4/OR8ooscShiJXY4LzJf9IZ+gsQtKGRw7vhpZCpwaaZ3aJhOd
yvc3r/wnZJ2ksh1yuJkFzbhDedTKAUEqjd8Iknlg1Era8C4jH2JweAeeiYsA
TNkC8nBxS7unCj6cdaUia6v0ekEcnZqH0VbOMwx2KMOI/NIreDukutzKhkTJ
QEE8b6mgQFuuPR07LbGLhzCgxdSr9EE3jiYGci/EQ/iFQJsSJLlweKv7lP+Q
JK71+ePY3b1VHKPX4anKHVRQD1ZTxZJxAuqsnvqX4/07YEnStCXTsaq7d93q
YQ2rrD5nnmIud2qioPT3yPiy0BtKKeD/yDAEAD/KI+h6rhN8KzvLqZRWun9d
TFqs9uw8M09EIzQvWUPki0o7B9VeTJTPe+ZXLpQjyjODT+UEKqvyrAphoEkE
Jt9DRICdQkgWlDuTiYKSoBV4YpAOhFmvgosuq2HFvVo/098I/4rI6HSSzuhC
DdfA3irL1ywlF0aH4jguVfJ/FqnmtRWq8b+Mq1U1yAQ8gEN/kfTYtwnndvkr
rXgha8G7RjXJsFiS5Tf2DxG7DcP65ZVWrRX/nmYfpBWzTZegPqF8D8UI1580
EUAqYhgdYwUa/ZD0iyIxgPc6liNbk9pond7BdohZJ/i7ddhRThYNVSurLhZe
Dav5w6tyTkuKfLnnioaUQkkk9sJJ3WAd3iTHePOaf77ZNewmV255VuzqW7K1
8OW89m6NGnfx5cIVsbsK5eSgTo13md1l6eGRDdqO7Fnk/CDSerjegp7CAh39
LrdQZsUFHXugl7b20arCOyHOthjskIGrTIo1PdX4D7ewx+PkjirQfg9rOWcH
yoDrfUZ0g9PNLW6pOvAugYtWqyMocmdtWKtdHQhqRKQmK3Nq/AcmBP73dSNx
ZtFYPch6qGjQ1SrL79Ni/eH1Iq4J4NVxPILy7sSLzH+L/xNvmmP5N/QVuM/z
EpaPhqeMtKX8i3QGCAexFGhX1H0DZP1VeMKFKsE5evsnwgiMXoRXs2RsxCDd
KPcdrUIkEHbX5hnUnDMj82sxEWzBhpPRPZMI5XV+Fbf2YEMc4UKW+EFe8LOO
qEhkOni7Zt7BzZpbygGfslu0mAHaorSEYHiI9aW9baftPEHLoNTsV8bl6SeA
B1uDbTWtmCrCbLQX5D3iQAcO9DnzReWj0mQ3ArqXekriQieh1lN0Ax4s7j2e
+Fkg7TLQpzz2/lc7b4x283Kkh2SkNra0TveswWzPOxtY00TYj2CczYiwYS8M
mcf1rafpaN9tj5quAggK2fhzLu8aZFffS+i7tgWHgG6NZIH1t9vSkL0E71k8
OHifyJizRL3J6VIqijAbNMEaappEV3JXfSoSZPtHFEJqQikn/I/VlqO9yYLB
/xDHwlY2431QyC90kT8qjD1/kMxqir1wpWUeflkrIzYVivxyEHNXpYuX7ttR
PNgxQ9JDCeDBIXiOufb8hhpMTrc/GpR1EbJNW6uQNyYVcmvA8+9Os8nZu/jG
jgaOtAd7t2SJdJ7B8BjC4FWJNQozhx5kilP/M1Y9a83XXZwyqCZsQO6nq2Hq
0VeQT1f5enLZ3eFHRSgggMAkUG5BH96WX2fiXSm+ssA1pFIiZm/I4iaqizHb
A0zzxERO9ea2fOFSu6wHkO6xssDdnCUg36amAIFcbLvBO20GPQ2AB807nZw3
4O5quc92Fbk1umy0XAtuNiUomt0zIkyYGa4RwgOUKsdspyXMyjqGLsl/MK51
pOPlrrZhnLLsbbV/fDI3xePXGyRlMhydq69/Gl5LS9CgwbIDd6BfiUpAMG6X
0d99a+EvKFSNzfA1zeSRGex7DlQSRE1L/tLSNk1m5ONdbYL8W8gmQ6NslFw2
OZRHTZzdYG1+kdCQ3q5k7sgqrrRofyRVJU0tqKKOUenx5a9BBe/IGX0rviSJ
rWcte8dwpK8JXsh9eDQKVES1veIkDptMH1R0St90O/MEBYJJRCSScq2wceY0
5U/zmQmx/u2Ai9PRV7tJJPtGW5dFv+BK/CPfMK5Xfaoc3fbBWKSj02mqExOR
ZL5NvVRbjuWlTiO6G9x4g5mRvir/sQZDlYz41VAVQbVXlyyvNemruZJeePCE
Zjx6Ne8t0nrjCWilK8eaIOOSOkC2+EGvG+6BhkziQBwxVl8FOfs8S66wj3nv
hUb/hTAjhtR/9z7Q8HbqB7dCrFsFZrwCWHlRVErr5qpVUidxXgJ5r33utByx
wrJPjO1Q/an8hglbTJP8R64U36Luq58e4IQOzgxnnSJOcSsDjZYsEZoXvPy6
otB2afMfojy/5oljx7AMIdTQ34IYUd0IxE5XSVFRKhHou1ER85cjBbZm3soq
faigkdxLBxtIizfToR+aZUAkMNRHhRW7XIXCZM9mNy8kB8pgkYzq/hBAdkbv
EHU81xfOobhO+9rz/Js8TxNu6+pPx/c0rVyNSLc1kzIik3mhTAXnc3m831DN
slbuSJ5wHxlxLbwJ/pl0WQLftPqALolaV/BL9LHJKE7BoL4KfoKgdTg1uEDg
icsjcd9HDjV1a8oJq/eIQdye+/geQf1k3W2GmgZq2uzh2qVUkTmj8YMFhYH8
E6D9JTazWoI6+nlk4d3NprroagviNKLaEjgvDF8Ae3//evP8IbGI3zBEbTqO
+VilTAL4bkH5PT/MJ9ipMqR8GWxdtBR1g0wWakvfg+DHcws0M3mKwC2JwOss
O91quh9Ii53OCX5HjdZsgguZknaMI14dGVNbnhVQUjueS7EyFZCOBKbbVTg8
rQ8KJvgQOv+o2PVKpVOqVDFi69W67U9pNUdlar1hu0LFMtt/q7hJ3zreNQTQ
OlfdSCWLzNQDjhxfXBxDBUb2TQ0cKWouVpKrvDPCmgCJHnR151+N2UQEaul6
Cx8orV/1O9udi0agbauICy+AYf5owJQZCvkEEt8S7ZkcLktCb/KzZfjKnpRx
U1ch6HotF+EdrQtL4xqQxUdCxEj+wvOGpNqY1QknZXYFQc4QLn7MCn5QdEpz
F00pG71dDttClnV5rbGIuZ0m2cWaGxlQNP9nHP9+uOeKwNpLasezMf3RRH0v
TJ9/RL28CJ/s94KDqHk03xMzxZpujmtly54DNqczmLOz4P2m0JEhdzYutgc1
ucrKFnnzDxhGCswsaKT0X1mWe1mFQ0lVNOFBWGI+fo8Br1kImboB/3n96fxy
Q2ml3fPr6PZ0Q4ApG3ZRAFDcdAFgzyCkMscG99hghPiSjHr9zU1chj16mGy1
gGkPM6K6QnI5sAJPD2QHd5DyDfXYrw0WwMWexRzB3j6HTnTpn7yq9+DEI9Jf
n5ShSlICU1+wFnHKpoxVvGim31iQx9NFp6SHjxP//R9Lr8ovNnVfARrtUUhY
y9k3RT8jBafIlXb47nk8rsp/dNWZCmaTWuQQ/oWRFXNu6KGRCpvX0wIIYjqn
+7tA+OgBCQ9FvLcqZDMoFb5v/z2pOGOjRQDf85isbKLd51TQYMomsd3FOm+J
ZRmqQ7Qa0geDXzx/un3hTomRmMsU362nY8fDoXfyu2meEhSFO0ZBnFJ38HUH
0RYTM21sbmonypwfrC8dVfEPm/REz9XBVHqcbEmPj0N/gkJI2I9rDKp9WulJ
DCvDFxvBQ8QCFb1RlC51ywkI39gRwPAyPGHOCwYlrowaCc7qvsOtcaXLa9hc
AHWYAqsUgI0+b5+vvaEq5WhSMOecwo0gWxR+dvZH2AadTNOBYgUquVJi3V14
hM+Jh4TJT1gTVoHpd9qnRRzjQXOFYiCPyuWXnxpOIWF6z9eSQqc/yWvI/Dr1
4Nr7zhoxPPPLrfq+WETY1/TEsCXHEezF4cMiczDL4Ivg3lVcYtALwTY/Qyjx
nWMXEYPOPqP0mpfW3Fwv8klJ2kg6HcKvKQwvetI97DkigVHqcurMRqU9kblg
TbHBhXGRcKjL3ZWcmGh+aeYbZA8Bprm4zGRlnB35e5HsM4BdjZ75kP/x+xXR
crIUALoUCLqtPLK00fYs2QRDISlbcmrpIKsoCXmtlnAniYZQJ21M7QBgITLO
/CsIyOHTbF5e7epX9pKqacFoaVJ1+JElvBMYCKtyHNqGR3lml7CQzzNKiIxv
sDTfmktJRBU6qOFClDob/6qU7qNEZ65IB9VTDWh8SHf2UZWOd0kebjXseHG1
IcqukSmtZhKi6UR3xSbCuDPtMQfB9e3vSuEsqjkT+6qSOPmAUYB/CNmrOqU9
zJ16B8t6XCwAaG0nTqKVVowucFj469fuBOlSQD7moAO7UgcAe2U0FWQQrgS7
UW0wE0uIauSep0JgB0BMBE2muj6bfYZBcu9xECCinLk1+88fuCiR/u+s6OC4
MCL9gRM+pMqI2OCPvEsHh3k0v8LPAUgB5WfV0B+bH7zTxCi6OzCsjrH+rhV4
WV0PC3wn1K7OQLyheAt7PqhohVE+CWH4QTkmBBsNVNcgn0KWJFJPhOb00DyZ
Yv7QqWfMDVCqFeuVTfE9tZ3GjyrsF6oglZKlfUpauQW15xkzD9tsNigY4sfU
hBvK49ol3V4s8dYt/KsgA7wadphLBCfe9RaD9BbV8GgDTKzlj7VG1q/r/Zed
OOTmYW1Kz9juYEI4xQCzHVNuDbDzYGqA3UGNnTOOx6LuAO3F6uQoNK5D/hMR
NGTRd5RMf4MDKUfUHW85NeYELOQ8T3KhVWU/M47o1rexzvAQ0TFDK1oVckbv
0GtIVa35xEyixt7G7O5fQ+k01i9Uj1lDiiHuSh/eYEm9V2A61s5cyzMjHomu
EbV0/k9vINLvns011DUpE6zO3MH36W8eTcj2tSAiw/GnT66TKj2bxCpjxOg7
ozMmzdaeBsFrx1ddUhTxbLD8kAHgs/kJqcF7eoxY3irZWgIrNY8m4hd5ZsuO
J4i8/pUMDG1R4hu5Ft5eMgaSM0KLnNhSXYhEdLNMyQkpFUmXJZzZQ4Z7MJje
XmLcIZMbsJwl+dui3PFPEwcD0azLTJks5O/p3rR/yjSe59VTL8JZFIHqtq7K
U0YFwHSEiF6xlAlzVuRYKeOi/61VhRX/41Tuqd5oAzwFBXOxKdaotzO3v+yn
GjjfAKXnMPz5xfYTOFTaeSadum9gj9liZdYkLOltiOouzTSm5BATFvaVPr9D
XezF7K6e+vJU4635By2mEgTcsdZ12i8ksIx+pWw+Aucd/22lHGUKGyho+aUQ
4lf8DOLb/88Mv/DWHoknNi9KjOzBq6+FURt2IOb8GKiV0QoJ69QhcpBtKINK
MgwP56r3iHRDvlOs40305R1P5lAzBL+Q/FHJPS7jYwNVLg27Ler0IB0Awij9
49E0WwdNIgNtWvjbtHAFTCNabU60z/yCc3qZY/LNeohwcYHdBwqOfRKZWIgz
4lOqkAvDueskugFL66Mz6I6Yf9G0SzFbnQIDVsiojSJkvEpsNisGyLI9Hx7A
hcAO8wK8XZfP1q4nlYM46FRq2jPEI2vXgzL2aqCsYg6VC/C9a1x3NjFPPY4q
zNqKWmDisPw+ujp0G452gia0u9kdqcCMS8U94Ws1lnepzW5Dwjn9K5SNHwHw
bAEOLDBXeScgFzsLdQZsGWMPHYMapP57oyriVghQ45N6Cp2TTJWa1QXY/Bev
A43IuSxqQyiPpbOq+prL+LH1mgFeo08R0fncUUpaLe5chEUO/6ro4YLGkCy2
OhVoIUt59aKzRiKoNvTInGTjL7TqDroTGSQyAbBZi53q4bbJQiVvoy0zP1Z/
abssWGdTgAc9hYMqaXBB77RzRdjcDajjhwhjJi/3MtyPLp50uMMZLTQ4Gbhp
o7k/3k0IDmRYLaVply+G6BijW01jcrL5mLYyS9U11IRe+h+cmCxuE91ryZei
hVw6iw7Tg7v0+uGd19JlKNGvHNWsZXPgKknmCaOrZJSo293tafvPN42K1wWm
Sts/Za4yQadvbeMRjKYswnrYc63NuNleDJUOmP2vt6u0JeeKsnykaHhejsof
eye/TRZMvMRiwIkkaX9V8jWXfExWkD6rkvsZ6KvLWP4Obsa0RWdU5Ip4Kj5R
Kp0+KCfoEEWL+swjAvWfjizaw3Mgao6ztHyLZO0mgwpkEcN2vm8YkcGS29KE
zK8Zo92/4fbbki2McLsZ0yRf64kOGR6054eZzp0Qoqg4SlXspwJ9D5WL27ip
jkqeBq6m3Lq+mOEWXiBW6wOuiEAt4ir8nF9jlcjxanYRmyRORHaOHjm+0UTe
+6IxvintQ1x6dpONVdYmxn8Pc/CWtVuAJrw0glL/eER6WPwfiGvOBdsPVj1B
ADIOwi2xlKWWW2lvMKc+DFBIGqy1qWwI7+SJ907IWmEAlf70MK2rsggomoEv
asBUJzkdUsPRNMKNgoodjvWsOm28S+3CQwgJqdT86qMdL84BLGG7ercDXKD/
1sgyFdRKBKuX5eXO/6vn8X0pO63LthuhPjzSE6KmbqlvyyBr0Hfb4XLtROoS
7tZ0fNdhJG45V1wdfNKMbTruHibde9wzVAHrnnInXXlDlI10jUVZvEhnN785
T65LdkGk1rwuBnW/4SnnS5OilASWppugmAkQXTUWc/Emmd6lS6Kx8iTPXty5
Mh+LOM9ZfC+J2i7BA7LgAHdnN8u2IWVPO5Av12F4Imxui8D7TTg46H6r5cFm
ekPgfq1gtk6pXfeJ+uLDsF12fjQVuobrBNusm1VjPgHiDMzXtsGBaKmSv/eV
RETHTy/DnaezTg59VKE+GzedrwRTEbGXPEbPaZsOPfhgc2SgVYaUVD0Rkumi
T/jtiOgaTcL7Ik8obi5oLoVJ0+CjfXmZtnZFLJ4mZtgMRerNm9LRffl1vTVA
AoLr6yBDEzbBy2KjmjANcZaqpuUPOTeX2Eppq0II1eAMVB1PbEAW14IciLvR
qod3CWMjYCYSAKYyCYenr40kEmywUp5TdBXe1lNLYMZrTrS25onSiey8Fk39
rcUtG62zLXGOhZfNoJXh3AnCCv41XWBnRPRwawYXV/i3l2GSLMyrTPde4juT
LFKck0ejAsrjAVAwtg1hc6OiGuE/DDcGyovdhrrstucCjQt7OaXAhgRgCRFD
4BTwW6OxR9f6+DaAm1PTU/C1DHpBvIx4op8vS33+P1NOGNMn9BPgheRMPbnG
tHiK01UHPwuNTeAKYGX5q+M1KkgdZoemkWGRMKyWzS86AN9J7iiE4XxsxCT9
SKJG0jNKI2aSqSmsT/BkUmGacw2Su2xrHQfdL+nd3xkVboK7OLpV4uTguP6l
78vsH0a4DbhIrbhiDiXEJ1WShgBI4gR/WYgdA0UKDtnp94E8m0XtluBnEGar
8GYbMxeHPclBPuZIqP7n9BB1QT8BPicW3428H/tLhPyyyK+2d57k18qEI7ZP
YIWC7wcB+0ylSv6VwnIVSIwhUi8DadqADM+xP1K9OFuzPs0zk97TWh2409lB
HZ1e/Ul/tBPKFc8TP0HVlE4V5f9V4FkUlPYcCzxh+8frmA5uHEMh4aT9j1eH
hswwSZUYndbA0ddWMpVWTLNBuwbf5+PFI3hmG+oGXsGN5q8n6V6tO9A+CJOD
G1UgvyxvwC2puxPhx9yvEy0qGZcRo0Jm39FbRXGfFSZrDPEOaBsAq4AxsdKF
KWPXVlef+aVTEd8lLTb4mGf22xl3pSg/6hBm0pHg/sSAcft5rB34UWw4j3Jy
cHDBk6/I9Ta+6sSWp3K18dmI+KQlwaaEJw+3UNa9fx3iVS253y25HHTTvvdM
2JlF+SbxQbPjyaPl7rE0l3MCVKCiQbFHiJ6PJDK+5vybvdijp4JGqk3n4zDz
eDQ6v1Dp1iIadjB9yDRK4BMDuTog9paJZ6o5Cc5uWd6+smAFin8uso8gZWmi
NSNIpCZx4fUTrkGU1oD+4R15JrxXyhFUw6809ZBrQSFM8aOryXHufxzTwmJt
njP63EqwPIEx+4jM98vp90IxrGYqRgdat2fk2filvnK5t+9zhIOt3ZzikNeF
jccNR9RRHCBIA0miO0ESyYtmEA6yY4K+QzQX4Mh6XduWL19xH8Ug9TTGL4xo
w1/O/OUfGne3PFxL9ur2ovuzKTxBGqNIsj/ZWg+vkYmFGBDhWv0P2ylDZqbM
PR37QmN8xYf+cJxp6Fs3WAwYnOTjkk09GeHuNXpL8gZKJhsjvrH5wzhIjPo+
iYsfkAAj+6TbahnqPmQ+9Ad1IsL9oN01HR6/ocvoA9PkrZL7xcU4+PberI5E
u5vfkgcyh5xlh+VjPHrN03oCrXGrkkwX/usA+sY/rEv9hOtRzyMroNr+WGGJ
I0HZb2nHmHpI1IcQQvEz34PFxoc/3KIoZuzx1zyVAWa6UWIDLWRtRu5ejkjM
gJ51zXt5z1OYK4GK3TPfoaOXQY5WWOIj8v9my5kTT8CRZ1GRIA3PizsNTPn6
5yhvo2QTseb2wplRK37dKzjlxiAdTcxChX64+sNEsATyeZFVpzOnQt8bbYXK
Mr7qaxCKHQPexHFQMOE2PJPCY5T+OWSTW7gmR7w427lF1o5t2uZIDbU1Yl3b
Wb/F+jI4d5deTBpIo2QX/P0IJXKpAkzJYc+1MY9SSeor5thBGsLiFXaPYhKH
fOhJT/+3Vpomr9LjzGM2FL7TltVR0qmcjov56RHZ20RE9ks//3SvewcHW6M4
SgnQaXOYMCu0YRspmEIjy/roWtJTCg4F516xHuiGMyVV5rAtAz4XdOH3wzl2
UEQu5to9TEqMYICM31xCBYmrGZaBTBTRqHwW8bOmhpaKNhsi00BOv/GVuc5H
jHjAUeAOwJQ7uzC+mtDW+IcIA01Xz4pH78GjNrivTz/yrKaxvxQ6/SK7Tazi
d5odCaW+5mIYON2TJaONaU1YB7BtEx/RfTBUjQwxc85w9r+qRwHdu5wjxd9Q
zvQDas5odVyBG9aoWRhFyd7Ph4MLR90CP0tvtD9VrWveBXKvBjZsxNnEtF7X
C609M5ZjoOxV/CwYsDelc+jnWlFzzaRSIod23u5XslkkKD8FiOlJlEJvXy0M
yzl36do7naxYlUPk0XhJnWdA7APY42YdHDN7a03RHJczZJ1wnXSHgtdduOXo
80YehDum3gb3mBJqE6j3HsqKeeqbsIl8KE+zsj9ujs5Gm87e//U900SjWsKE
DQsu143cq6qgbQVQylDstdXnylyhpznOtd2R2Ucw8p7FK3z1DWKEVL6+buKN
Q1bdhc6e/0gE0Vtw7vTSdVIyrBq7CGZx9rVH6YXUMTw9026uImoa42iGjic3
DcK8qRuS/2RYIwO57TuKyjb8gAwGY4zcdBv48+d0WxSzbAxEjsSH6GUSGp6B
bFs4hGEg9K8ZCnny1oVjsxJyUXkixG/41ObcuCEuCixgPrpSSOQLl3gVJ9P3
zXBFANLm0TWWXLyT0dF20niijNMIXpJnk9w866rAvfwmmHutw8zT2RSh8pA3
85kciOQhI5IyiXZpwd8vGqpcK2O7gbteqcprawoRe8rkwnscBltkFDDNwSdW
WU1OCpPPYBReWBv4b2+1FonRFAADVlgFvSw0oSxgyD1pXYJt/omiAsB++T6f
xKJjwOobIINgLegLKz/lhpmssM/8Fd7HoFfCCpVltZVYAotWviGzLTGqa+9D
vz6mYwiNObgzsCK5FBOfU1SLRIi8tjf+YdHZ8i1UP/u2CUgNPxURB5HvCv/e
WjCcmuTxHjhrwqZAISva5U3kMfMEU/SLhKhArsc0ebZMVqQ65iSD5WN0otrY
GpPC661m+rF8oXaD0amcnor24gZblhaevvp11Z6+bIL5og1GsDc7GyMEK4kz
qKA3EU6VbJ90EygklDCy2TQdsXy4It49leaobbrEZ13kME73xr8ffWkwQEEY
2NCD9/dpQhBu5klLLZgmK6emiPhlPwT5QG2eTaGIZ8NhOKC2VB5G7L/WyKVX
tGnz4Ecd+1IVcBG6/IcFESPUZAHkt5/n6qR2zNL60/g3f8c36ViMY2haN7kX
RiwejVJHc2ubRoGTucIqDBLzuZHx9vHR/ZRNvLbECefTK3INqq1OS7F4XS82
AFtfjk4rT9wetjviXNy8WepmX7MBRycx+kyBq+cds7aVZ7/xUu0gN37DVnzr
CMSvoAhJ6LrlTRJUXWmxrHHSI4ZhMySvPa8+zMtkFr5sT2FmJdkFDUKklW/O
/1Vou0HWn2ekhtFFQqdVnh8zeMu33zjr28F8RRz8OLED2OCBYkDeoiw6fGqL
w36KAU7cqJzkpuT2xNJ03fJBhIhhOB3rgHWeNw3KQVVlZlWhtSwnZ6lKMZ7K
TczP6otAjlDnd51ViIhvgK/E81Hh4u8CpU0zqzj89PEvAd2ftDdZtozZ3Qb4
dkFCS38WPNJQALY/e+wnHJIY7vII/AvMIm4e3js4/r/MCXcgIsgFL9VhZaRN
v/0hBfOER5eo2WDGH+zmA7xmTjz0YvyrnI1icIsil5Qfp3BjJit6D0/sOOr5
FbVBeczHBhvrexFz3U6coZHxU41GUQcs3cDQqxeuW/17pFlMxWUVEhFU0M7r
zosNmfcqk5yj5WPxHfJ18stkQqyxjIolz0BWF+sEx3QlHHA2tokg8RUwkqIe
I2PqoxwzcKPtj79RwoTMBLYeSK1a0Wc2F7liGJN9EFHyWzleUznXOfI2K0fx
TaF6FhMF8Bg8zWg+tl8QVXYIP0fiACo2wCd9+ggCFBY7cjmGCw5fNDBjYIWq
hJkXtTySXjLIgTID7yTHNpzzCYHqCn7K4qZWpkCGWHvt/O1SNwoVCxGX4sno
qZjR9Kbv5ftpTq50vkOBeQZncmlzLN4iNBW0k9uAVxpEhWRZ/945k1eoZZkS
R3GrBdgSwf+F6B0op6i2uO6vtZihOQJ+MNFJhRDak2XxTqud0QN5rlG572/n
wUAU0yfUsWCkYbWd4lvzdPRqcmP3HoAzrgtiyn+6E55OK2t3ve83dZQf/sIt
fFFUwmxJkO5tYhatXD4CjsDFZ2n+EASYMP/KswOWyvhywC55+OQw1e+K2bsm
0wufeiMuSB42nYLmI50o3XREJTtgO2oFM0HsdOJ7SHjReJT49GBFGzZZryCG
KHxKJIj2dlZwHhpD0l+nNb5MXrAjQZqKIL+TKANvFFsqOXsd9ZaZryB81L87
lXW/EPxMl+I9Y/EmMdOG6p6SWKSIL/7xqFHGf9jd3cfYgl+o7ib5sdR6RhjP
4cGFr0FdCg3fHKaUiDmbm+Ekz+hGrs+zkinxwwWrNXVUqQj5FnTvYsiv3V0+
n19TIxK+3cJOKApXSYOVwx7SskO6j38bCPM+lXONm85Hs2qlK4RXNQnKPvR3
GvrbPGhOQgbUPJKzhZpR7SlYy50XQ04Z+PDe16Jsagcm3TCvHp60PS70d8G5
PV8a0fjXKlhF63ifArKsZA4R2oxYANCI6W/oCSOqwnJKSObNs4rV48eCQl1m
YKr2hhSTluMw4PeplnI6mn90D9Ndx8Eid4pqQ61+bQ0qNmGqxJL1wF4X6Wlo
Z6eLk/1yYOtS3YMs9V+pWfkl6vCYrvUtjzyBOd57cQ6pa4NTSWifsNGO0UjN
MAbCSsoXpiy9H6HNeV2cYszRwAHteLEb+0Q9ogYo6pkjzQL1cvLVT1bf7+bV
XaIERS8yYjbC/GFkLnGX92krfa0Hu6oHK3cq328Iw62QdNISlqhMMcCcfHsI
g7cf/4Nm86DlFLdyuDpCfE2qRQZpWN+MMUiurB8VOskODPLgo36YQnOB6xg7
hudV7O1hxIkAk+27908ETUaFrwefOKtfkO9oYAOvRWEJ9PM36M1iq0r5ZKBC
asumgFkJ5eZpJUxVM39fTyV0E+JOcjn7dTldDOW6mZy+1Ka0CiVc69g8ncYE
gFwWu8k2N9UzSbN0fI21LgIeWGUi3mR058cfKN7r9e0m0+TbJeUAa8viD2Ur
fF3XjGZTPUDLEzPA/EyXto6jCNK+twmuGVKCQ7I4VMEubxRM1+GWv8Ai+eFw
vrlfeRL95ofoy5YsO8MAcdpPOw9xeLQbKFL9zdnkuijMfAzm3k7uI51JuS07
bPb/anTxh4SWHlYPgHLRYVCVS1Fo3XjJiArbGzyrJDuon2A139ApvjM116lf
XVmnJQ///DL/Jf/b3BX57p9lSm2zMlaYZV677EqlcFFjgoneur3Ekz4VGgK1
JSl1yCUt8PiPILpVJM+lu4jU4xS4NUW45RL0G7IO44p0TVtAptOE4n14yhcV
E3OIn17BpJHrKkrDe6Fi9mPXIxW/1Sf3qbtWIEHQjT5uoc/hluX38X0XsQez
FDNQznh0Yp0TnpL+kbVNADk+rM+BbMt+qx/pHMc8VazplyZbZQ+u9KI1Rcja
wz3vyY8ZvesMZt7/KK7DPl7dlPFX3Iyuy16k8NMNXUTUGk6ALXiG9k8jSzgS
+sBYm6XPa7+esQD29ueD99/90ihE0AJDTuCY8IIncvPsaJuc7REACDEzgXnn
oevkovL8U3ksO14IN70tQRBQlqrI8Y/bdaKNH5b6FEhDR80huV9vaIUIKR42
2DMl69rG5e5GTSRwcelXkHPLRmPpyknDlyY3d7prYYeuszctej8TaYuXfYcP
1+BqSUgeHrrdMCwMA1V73nb5lBwfQyq8Vup66XkuoaKDJZ7IISHnz0DMhCpY
y2BbJUfKa0i03lcwOL9XDWF3fLcTJH4fhYIvU53H5FZISbPBloT6p4hXUfXC
BWL1k2e6xhuV6jOzEQinxQWqXNLU1qM9WS864D0NJ3JwrwC/PPtUpEPO7dP2
flCpfPafkzwBT3bPd/u6MbnWpax/Xf0A4Jem4pnAzRmOMtsaxyUjm+jD8Dgk
s1MlYDIvyUOUV8IQhR1ehQ1gNbZUfCrFidyt7U21/V/bC1fFz6Y7UQz9bp7f
7V4d03TR9YtxpPx5pKzAZwPPDxzeycUR81Yk0AWmZTuXu0YTpMkEh1dL/Sq3
m5+YyhzU8HOp+z+6L/2TUJTLvd2MpK9TvOJlFMYGNorZsUwTEG0oE+5mpY8o
wzQqtO0a4kdhfcI2gU/h5W6QkKfSsWQpgozyBwM2oKTJXVshoNuXp6Mps/9T
n5071ocDo2kBVW5NXiCnreKjgrInMBwzPwZC1TuZHtjImiiNoojIkwK8EsPj
vqsDpH9yGopowpYJnnByApM3rnvR2OZZGPAlpzsvVYfAdYiyDmWCdvCZkYym
Hi0iT0eBG726qJE8+Loyx4nlT8trj7HXJgSbqmNTKQyzLCmJcymhAqjXfgQf
IS44yknttnYSuJTnVAXr2DT0NkfI3Vv2erQ0mMrc2cGO9+UdLq5Chv8Ya7bB
lFOf0aPKl1CiZkbjTCjR3nkn+iv2vogTUm36sMst1kgiksXcWRtiFh/uPzCP
aPLTqKiDQDnoCF5yeiTe7RtxX5EKy9d9CVkGHRjNuBC/gI6kSpjDxXhv0PIj
0Nm5egeLv5tvRkDP9nmSp6ZXnnzr1TGNn8uIKdZzykTgXBIvyCLVMsDnFhvX
776acCtX6CpPbdThyP+abjRMRXyFl9WCPlet61A0G9WRBMosbkeBaQd+Iym4
V9EVy1y3nOBlHD0nXizYIFNPBG0G4aryjkhBH8DaveoKyzfU6TRTNItUmVSx
GPlK4MZ8UzKR0cE3qZXb8i8T9yq+seZM5wPpTHdZhTUvY0Jnm6qvd+tuogEk
l1sV1O1TYs+hxdk2RX/aFRh8olJTNrrKDIflCWHx4LSZI3sUQhcY926/pOlB
NghTGRaZgH9FqqpG/0pR6owLXCUX7EcSH1mwt/HSGdSzlKLHLlodOZKx1T5V
x/PWjylXw/CU6hOZhDYeYMyd6WVKvBSO//bCyr7qwMEWa0zj6cSefyGjEI5/
7BQqg9sfN6K4KHeHpcJQnpQ3BfRHjNiJ+SbdjNJIU6oNh7ZsMIUKSjlgpV4r
ZDjgmtlepPBjCn4DZpIQ4rk9XN+q+6pViuan8o6FWdQlxQ51dtc6/ZATGV7n
Y/uscvEew1KJPoL4/Zcr3RHbwTsGBI88ebq6MLKSzXUas8RJIpMo2qyD02fC
DIwuQMl5SbrmFJTC8JS3wCUV4F59aPGYOvLsnNFfNt0uXNavb6/+TU8Xhpgb
fFsoFeSEEvC+U5glgkWvQwg9LBDYKdBFy6o+08sEwOhet2JBxkLN2Ktys1vT
kxqONnYfACQY8U1m7XM4fWxYmAPL99Vg6ywCeRXzrDB3FWudzvAxuFzNOUfJ
mVg6uw4T4OTfwzQqnPk+K6X7tMH92X5TZvKyOYmXEjxI61FjYlrsNFgvISv3
HSl0Y5LdtHkvK/1/8/lXIc6CKTA3myWpunDNhE5Dst0OXRypN2VDfqnhBxGf
dMPAackKCKr1Gi8OFsZ6OtAC20CtrDxPd41YK8ZsIlWO3ExGBHR13oGBjig0
fPivil4KJJ+TOuUjN6SjKkaHdRR++K7dyrCYvMJIXvSM+XQ5mHMuVQIldukm
lk37YTI6oXkVzlJJNjyZvv+OzjfS2U/xvF8xlwm3oUK/WlELA66OHQ5QOH0J
Tk2B8k8CxcJPy2lzryk2UmAYA7k+2qytXsBTNJvOcizk1UlaQr3B3T/epZuD
mvOK+L48jadPVlrmkSQfjl6nyTSnj3s+ayNOGbREaExAnCXU45h04HkhK0xE
EMlwHioq1d4TunsBP6PfUCMIlSuZhp+So6V1KsTi6N32wxlKFoDpAtIg3oky
+2J3a3n1BQuc9oCvk2HRo9Cf2lhUGmNDCQKD72MuKbX2ggi4V9RjYPikAM2i
Lz5ANPRf78VMTsVm3l6pYAgAGvukwFknsN7ytxIdS4nJkLSfUdVrIBFWKMyM
UhHFfGIQZgqQmCZucjWaEM9ifqVO2/LyCxNNYg6PVm7CMms4CrOOPH7enm95
BGt1h0ob59mA2xiRXfjkMbvmUhFG8T9mEACV28alhN3pmpMan+4D8WG9+gDJ
KAbxms+VX+Ju7sy2EBUS65BeSOfq6kaRqvwqcUCwcn7yapuPiZSADQcYXQxw
Wq+JuRxtC7/4m9GganEK7H7my7r7dOyB4+z8W6Q1ruonTUXyg9XQvMGj9rnJ
1ngKQ2niLazClYiEm6w8flXYZjhRoJKQxYh2ieygY0SXnZKO+7K+eIUrdnEh
mYWUH8GSdy09lBr5V7KzQjOweio4fhsQZCaD7W/O7wJCSoYzRrs/8y33kffZ
XdTqZrL1zKCsqKGl5ME1VoO8nFxkUqt16bKagEIRljbT2tSBljpvtGRfMriq
G1JJ/90EVTmXLQx1mLNhbz98XcciZytiRWylLLE6cKCokXWiGAEOlhXN/Wc1
pB70VkML9RCDulhoWbIQiOiLWsZIxXOJ7+vywoJZCWiW8frGr6dHDyufCdDY
wxlIzmYCuSGJSLhD65+jrLVFEKOIc9/OCTBd2v0/9YwcRA2ZMW5+XvGINEbO
45rRW5LWkfVNKr+uivDbfhGGMZrI4yeukIdmKIZou1kiWKxEOLnYg1jl2V7P
xH4Z/tDGq258YGrmWF+MURRUUvn6VJ4S7Oe27DAgiQ3u4jfbbFOcROHpFb/B
cP381Wa++HGLHcWEtkh1hRWyFsahMCmKKR5sL+/FlVi4OR6kWtIz4t2FcY2p
ZIUp5Qwl5IU34dEfutZN8w8BihiN7QdhJSV84vEoZOq08e/WqqUL15DSo/ui
7iOmZ5uqXsAd3rOiB6cBIxoZdkWqbe6CmVB1+inca7x20yoqt/mupF0iDnA5
1LERICxXwjSEr7C9Ndink6QIIlWmEfSZ7ocD5/d8TwLEBqEa0zw/cDCHiTC+
/B0FDfq9RMDaxoseH1yhI/A18OLnu+9/E3X0LoxObpetOwksusbwVXxZon1Z
ZaiwyoNculDSZ5Gz2iyzRCSgtulw+PuO3KrY3pUrfLTu2GKSmI8NQAEY2EVu
LzeI0jDqOqVtmy/zJiVjOGNuaBHh0Z3uzZJdnGdGuYXLJfXXpAz5C6AL0jV3
4iRjjuL/PCtPq9Hskyo/EF1OyAinlxzG4JYlqjqBbjfhlY2u1p3xY73dMwUY
Tqw1oAP9EcD/DeOr5oyLSJ4oagSJGwzGvWGwGdbb5AMvwc0MYv/Kskro1d0K
YskePbKFa/0ItkZPz9lqFXlMCeg35YyzZMSa6tqk3XKgtipDSYgFXYcI4Iad
Mt/ZrKnVQqU4ry+NRKRMRexl2+goeoobp2NsKVgoVIrmYLtnBHLHiJhV1a3X
IWNMQTuMC9Ce1NxYPSbKTH/96hLlOnhqbXcvR+to0FcvNq9F1ZtCvER9eS1j
j3JLALsGcaNQnK8jWcZnRVPrX1k1I5klfHTYBovo4mKXi6HCGbQQzCLwtc+E
YG/cozvyMFr1f8scWUIw9zfBY0vzSRc14QdM0QDbqAzou7Fp9qLAeXyo7aSc
z3UkLClZw6PUpZnJCRxE5r83UQrS+nkTx2VKcfURa5t1EWLn+fhrv5RpOuNd
YngHcQwVSrRloPONk+ZW5EMA3zGgWGAC6J/Zf2LpLt86s5OTduiAN4Sabawd
mV7eq1JorD25jKCyjP4Hp6vSpmDtBcIus05y1fzrEzf9OXLud5xY3W7Oppfs
AggnWhsVgxLThLhp+hzOcZ3z8PFoGS+cWqF+ZmbIh/iD7RcsFqxkujXeTgkL
jSynBUgEG8B39cDYoNWSye9t488V9w999t6ChcaqNxAeQ0qj4JSzkZ1qX4GN
cYFXDCDSAUvlYTv+YRgV8D+QE3iY6aLCL+y3DrKvbvUE+n3QcJkpcclXEQsM
Bo2rXfgenAMJPjxtLPaoCLBDSfLqKrcv/h/jIPGIp09qkfPC3unMlGkD3y59
pPLroIZO3hy9IuSE7/1hxtQktrVjWbR+TCBoCkUiAKy4kpyDf5bZpUZ8JI2k
dhvjesen4wUa2tNnWpCNsY9zZnhcsvmLO38tYTWVS2Zv7szkGyI/mujRFUbp
urdoHBGGnE2ut/uTJnZcR63Fr0ozDkCrgALKwsDnzhUL0pe5E/kTjAyV6aUK
OO1fV75KA9QIs9QHyYTZWad0VaV4vooklYqoknCDngG/XW0g189Eox5xARms
fXcIFVUMsj8RVUVOAxXIriitv4Sjjs/jTv1xvDP/JaG8yeGiX9roih6Khe0n
Nu+1Jtrvm1QABASXU/hrL57MSt/Lc4h6nHPnACJ7AIrhBrWGO54R3NzCWU3l
wHgwxJs2XAfsFwhN4LrgFwqakxGIijy/OPBygKV1wu3DeTlDqdgPCCMW4MpW
6YlKt+Pwc8E+7C6aMG5nrX7ZDHxgrRgvE18dmRVMLDgYFoo8O+WyLGpniaSh
ecURWOGvpsnp7mPTj1xT4tYs+MS8GI8bUc4Qur02HUMzngDM0lbFHPUWZTmk
yUiFiedF7ZTKhspPTE5ygZBtZJeI+ZfLajefl3RXOEKHWXtJgm26LA0FF8nm
nJFnUcwEjCtxt4Xe7OlaPnf4vEXhBgk9JbGwcmHcO+ZaMIIinViEYzc2i3r/
Gi8gHsDuqtdfA4r3mpIfBGYI2mk7yUoik3jQw4h5Bq+IFTKgAeUW1dJogdD6
XJD1GJ9y68qnz2JHKVEUHvAwWgUfedoXvEAggA8ophD/lGy9lRl6EIdp0Ka+
RQ1WZj4bx76IfmX5rm3YQtKWYBuczmQaGUdNDob+dbeTKZIrKnKAV9RSV5l/
ziDx4SCZbTz3aXnS+2ffbieSB//KTuGIhfw++GvWFSf5WDNKuRnBzTbOx/F3
FlX410ClnyuQZWNBCYpf0lVhwLBK9+Q1D/safoEgzRAEpNUAdQTVZtgWHJFJ
d7LrtR0ktbAZFzHU18fTfcPH4IRkPedrldp8MgiDPhM56vKBmslo/OrnfAoq
OjnTj0jDwy2B/LUCYUnAyJPOlklXGfJ2ZkZdo9z4key3YXn3hUaQw/GDbxIZ
BfAB2o2bdt8RFdZF60YB/qBuFsf1gsCsR3saZXi3DanvBaMuqNxu192rMWs6
XxFVYnwFq3KPZRD+ysKjSFac0SQ4OI2+Ocght3hYNTZ1M/nuniFOAeB88ehd
IPgaOrBAyjwD9oxbj0uTRnkusoQ60WuY6jqx+dsGTrxF8a2HoUg2OyDphDe/
eQI+9okxisj0XJGgfXYj6kj0smJrJUbrD9z0T+xxs3ndwnM4Ke0tCkrjkQLg
+B0G2ZkpvhdsaDuGpTXySvFAdvvcW/pn+uBlKDF8/GNwY+aM47SiSkAnpuSv
9/e41NhD4vJqOivtbVBPQnAdmRpd6HTuuD01zV2E4mrwDrZBbTdhYx7v/clC
bORwY5C/qzMzALbY+Qdw9GDxXKwFGZ9BI8PcIlRbO7fCmo1WVm17JVVHBz0L
xgmOHIDBrj9cIOaQ9Tw4zosQCuNEVLNymv938Pq6X4laFkO2TA7NZgHpLSoV
BIhZFAkFukJx+OPKrikodtjEBhu1iwNDTaw0bw0wOiii+LiKbRPcYQcyZ2TL
+DtiOKzXSbj6q2lGn82KxbUUYC8FgOoWQqdjZclwyb3fga1KUDgwnuU3Di8h
NZ8Fh1r7Rj9T+eEQ7rYU/EieqkMWkXEXTtnuSZdadCjRP6qJQNm0yMe+VusL
Pg4V2f4j8CvzlvKJ5LulSZOIeA9wh3Z9xeosVLwYm6IqzBhjgBcAO8qa4U16
+RDbZe4tj460XcYFXFE/zLRY/HHCBJya5DilWKIcuY8pvqxIlSnW5iLrx9+1
TbRMSFhklJ84BwfS5mizoamOTXnefXpBDjzz0bNi2YsVODuZHLhywX1VsHgg
ZAgFsavM0xImFfK1Lf0wowPq2ohgpEpWy8PA7JVg2g5NFcW/dVvdzsjawo/4
oEOKSC1miHbdoAGhx5VHPug/qDc2vXBWyl7li9F4eyaHeo89kweO9iT7ra1M
hK2B4cBy9zuf44MBBPWVKRKfP2lP967hUX592EEd3dYABqFq3PvhlFE1HCL4
TJiL1bl3cbuoI9GtaZ9gD8TZSjX2EpfKWn83Kwl9doAcciQCwDkYCK1t6lS8
/aTpCuZtpo+G6LUNSUTBT9BqYKNtTvVnp4iIATTCkvtE86uW2F/t4Zd94p0Z
CpcTTQPGpVQSvdjP8+7WjtKj+c8eUbXizLvtmpFmvJUfcfQ3uJggXTN/tW/w
ppz/WNlEeL8dc5sG+gxtHO7BQEYwMi2M0YbuvrSAtWoKogGZNkEuKLWohLq9
WXjJuD6+U4VrMHDX5ZCUcDGG7hianMIxLNeLg9priuY2+tKPwbELRjR4qXOo
CIOD7+I8PPyyNF5lPrLX6UhVUqZh6D9F/eyWAItrDOJw7S5HAIQTlv84lRdu
ALtUBc8kRzbmVXJH+3OGB0QH9f+z0SeH0aVG8gUD2kJqH/3XF11/sWKcHE2K
gE68ro+5jNee0VqsC3mPV5pG9/gK1Y/L/jioLpfROvOyrWJS37x+S/JTEBQ9
5g3RMCdhpeti9QZ9UdLNyMkaRYW6AVXDelP9Q6436XbW6Yig3cOrYkA5P6uR
oug/L5H69yaqEyiD70nG0RImWm02h3Zy4O67lVm5UbaApW3r3XQ4pDyts5vy
QK1b6jnt523mHSobjH5CL6CyAb0Za8AD5Z9ca3TGcFsAj5eBqZJauUnJPn8F
sVPZPGt7waGfUIcDsmdejnCLupHwhLaOPd2vPCANB4tMc6hnAtGNO6W8fu7x
Llumf/u22VeKkh8PTD8HHi9QPVRKTcOtJHtVKPn95P7xpP+CI4+vYdPjXq+w
7Fv46+lcCuEQCpqXPJ0OnaBXdmFCkPkjjbBr49z5zLFgI0p7Q1o/hm9U7Qlt
ijmiOymqGvkRgpP9PKAukCVEcOB89jGiMMMxDLuHdXs7eCfUGnTHdBRCfFtN
CY5PN35BqmlFKoxX85nV9NKJ98I78vhk+PuBNeIYqFwVlIBISjrgjPW6QqD9
KjIzRjwkgJzcBKmf1xwk4r1m2g9H9cxbdZrE/lniM4yNLV7CPCNjBzCIxcrJ
KLxLpmnJ8pmJuBf4rv+wv3h2s3emSrOLEMWayn3lpaEZ8rjQsXlZXmIYoazO
zIg3Rz2kD+nfsTzq9YaET5ecUuICa4JgAIhohZAZ/NrGMKXU7Y7tWWsfbyQ3
Z/1Y216QcNloD40KZwZyhh2Tho/D69fO9sCHGUehHAPG6UWDD1pWqs3kpeNv
GL7ie2et6Hgja2ZtzGdyr+ZEsvMJQ8nx1RAKu+e1emSmERff9pvM5pBCt+K0
llNMBFEeUGXfFW+j6yHbxIFMlzE6ut3dS249pnE3LOoHtjpKm04QY4z5/K1W
A0DyueR7f2Yc3VNfYXRWEh5cXpkHb0OOKNQybW/Vn838CCZAYpuplwTdQtwE
pWM+oLrwhZQ4pwLz5/qSAnLdhSV6YrgsUIkpwkHz3a6+VD5Jgvuz/T9+qpc1
TXCb5ijhrU/V5mZ3jtkKQ6+SoKAPJgDutvksQMcbA4tuxJoWrm3UUbnkJgwq
kT1+dcpx9qM1uliHorJ+ttAw+VzT/Ck+yOEQpzSXlFNza07Mxpl07Rv/WN/H
ixpWRCj0BtCB6Qa5ehOL0NQT/zY2Pla2lzYCnCgQ7mH8etFXIL8U2YxmhK0R
a/ebSi/kSarmnff6DV6RahJgz+DWTD3MfUR4/BKp3TrfdgyDHtOvgvYnJcvZ
GydKkoCtFo4Rm+8dkAjJ+LvP/+0HdMO8OxJVzozsojyZ2oGLOMRXGvVn1VYi
CMlsZrNm6uSSVAw4Tz32MzzyME2bABbSgGNCNFzXA/upjna7/A4HJQQx1ems
lg6iHCgs9W6+qRntKN9nV/35g+FJuT3mvUuPIaeigWa5c/z1dAyQH2V85/wx
AferkIlTIbHqhzPVomaNOCWv7L1BZmsdOi4x7LgEwXf+vAAFXqA9Te1N7JQn
fUa59khK+lQSRfIGxRlEzKplWtHnp6fmnt5y9C7yT6syfog5Ew2lF3dkrbm7
K14l2imnjDB+QF1NHqJPurQZzqa8Gm0YRK6rH7+k9McfoGqZrbCoIAuGZVuB
7Ny/omeWxvXzSjh7GZXE9Zan4GReRaQA89mIrt1Zq4x+F4pDOTW0J+Y7X0sX
H7z1a3j8BrEKrHKc/JFzpHjVNAwe5nRVQR0S6ppL8dKa5ymeDAG9NUvkk+NC
At5X74NWRtQ1uNG3MD3He0SMntPB+xZbXe+I+4kd3lQfDYfSo5QhCgvLoBoJ
Cx3HR/kOjlXw9ovvN+aPKpifck1sJAxqMNO/TUqH9HnAyybZ/kwrBMQaP/VT
YOqT86UO0ACOMvEvgStHStLJ4GPjzd/qbZnDb3ylKWVDaHnXDT9yDCkTb3m9
iPyDHm3Tk7DUse4pZ21Fc04Y4tXOsPzGkoLVbuvGPO5QbDvj0g+IhuHecP85
2zov3RY9olQlrqbXA+fAyvDh6sBcWCQ14SN2MGCMBmcuNV2ZpPOp9S0eQO+g
BPQsBCl03ZS50kkGGtD4Kz/zzun6k/GqyxF2tD+ROg8jlidWYiWVmfoQ3ief
ZjAZhOgGmoIH7jglx+VwUk2jPqTEI6FNA8HVPKSZ6rW9ZkKQoKthltEpFjpH
8NbL91Q7TyXOXQwTeJzPTbcLLJh6RW9/TcR18geV8SIasEDG58PakeZXMjPl
sMXQyEMb2Zpl5esTM4DEBEvmqCGeBbsphGSHJsnNyBUP0E4I9/sUtF/4XPhU
4UCYRksDihuyV9B2al6o5vRAbPNfwtd0oOj9urEPUCqF5r1wGj4hhnw/Jhl+
Y6sNnVzUbQQ9fifiav3K6estT5FgmOXQ3P6tzNKfJEyXfjCH3n6M9r5SmwKi
AJ1Pdjup7bRQQ0IYRM10HBFUd2zeNb8vazA87fMQ3xzhDmoAcPsc0CBSlaKu
1dbCUsSLw9IPYu1lu0YHOJO1vqs6qbK6/ARNFW4X7GLupoIi+o9GD9UdIqCB
SeehswLWpvaa+Rd5KyQ9wdAP48VHlDJJb7+2U0YKkCpup98UsSO/tbbl/X2H
Xc37ojtt3aYIcLe1WvXaFj2NIpllmk7hnlQB2VTEa2tltpABikB54fyZBGso
iQUIGvQGV1KgYJZFznUc5sy9DrjP9IWxEEvzrxiL2jBiZTsjoZPmhlsknMZe
Db9AHprfACS8yqaLaPjyyN+0e6IsuL72OdB4WH3lO57LszJ1u0ak0LP/GM55
1dqAWvTp7cKd1KlSIYjdG4Z4oNHOQX/ndzSbkBGCPTB3jTWuWOuzY0dFdqkX
BJZxgpJx3t+uH8s5FWBIwyH4fTV+VfPrHPJN1QZT/I2x7wOTf1jrFTD6gHft
6WXLo0BG5LOX2u+YrtuEcuEQ2Yygu6XxWDKw3hpWE4KLmRD/TZ19THkdedRE
X+alDmHqzcUlqsdevEzU5cc3gBDmGBQtbqrb/cKXapmP+vN+0FJyDZF5wyn8
vKXYg5jZp2TcCEEDlaNjWJKuqwITfrYJO9HA8ygmLgXC98aMF2G40LrprXYy
oNd5yRWwR9QOaVDXw6oSlhUMNVoFBF48bt489EFMXebxDzSY2arw0pAMoBQs
RQQSmLREv5snAakVtMeda0Tok89TTZsN73HmJd7B2LVv5sHT3nRPALmSWmfI
pbHuIJ1wzoE/DytsN9oSxr9Gzpm7n3gwnEjtikLvCUSamRiUWvBs0Ib9wu2O
Pi02LgLJQ6p9Mb5Es2+aRXGYjxLclLVy8XX9RCna5qdrS4jbeMo0gqZ/BkEW
gzzoqsplimGjGyiuNXUCjQJEdstH3s57avuE3xRtp/JSumTqbGhOKLo4A2pq
6aoFmlNihFXHQU5v6RsREG3HGkyHYo/tPt8RxZ7ZT/8t1yEc7QBRXJ1WVV5K
d/ttYMij0HQKApOdrYmIRfHGz+9BPQRBsAOX4s+6hJkdi7Ys7I8d8b/DXpgJ
QdAag+Vjc4luDGVAm9rtAlC8xSjI7XNKPJhH7Vwh1CRM3FlVaMWWg3wcvHw1
WVn8KFZ8m4ChDQxnVLh/ymYRBDxWUFfTov/8o+2z/SyuY8+adKLlZAu/ounP
C5mTFGFkZq9/gsDAo+lLNhn/hslTb8tBTGyPwF7y0Nm0cIMTN762dC7Oej7+
ARmcpsZIG6Pd9HHL5xaXsE3xvda+u+/mU91z/ys774y/thwKqi4a4Nk/iDea
erT/kFLsc3HDkZRvrzByISZUK1uT5UlXlGW+fyFDSuaGnUFH0R4GmV7oAfys
KVWg6x3czGrLLpHfIbs0P2mKp7+fKiw8ZKmL/I8zaBHUUC5zmWRd1o2BF/+M
LRNNsPA2yYotOMrH95H+H/MpbjBLoJpZXYvK8IBIsxju56ebPKLCDqgVfQPd
ZQRVRDxEewf84UtWLsOdS2/jdFkJvcAFpcQBisZ9rY9B25obi4nCjMepzZRw
oSgHvHdK5gyE0BopfNymYGbUFtPx1wy8NaC3jrhTI17Q9PrgCbh2idmiwWZf
dQ/nG2z8IdHmI4f2Xgj2x4vAFrIPxOllTJhsoYOVypoMGS0IBhVZWQOtqyvg
BjTYXdwEaqDXEExZgUKlPaGhsgs1Ce1LSdgi0HwdT94Bqg1OUrA/2l3P9+0k
UxPY/Oa2IFP7tkmHEdaeKkMY/2FXiP7Z1U/Xx80dsiY4HOVXIQH5p0VbRM8s
tz3U6HPDA7Yh68FwHCyMNWuw97zFmokA+MpLxK3nAzdYl13V4v4IHQ50IBaT
e0/w6v6ucYwMK4qkjwZgE5kI+ItaHVocM6+1uV5kfiAijVuuZ86ymljJtBjT
6Pl6phlD62CeWKQDuwQTW2XAsPlQqK5U4Vw2s4elQuOzDUxFsOdGR9vr7PFR
4FJ9Dq+stJt7x9iaKK7bPZ4eUMDugL10Rd0gr/DRqTDvh+dMMzcPCruUaksd
8tU0d75jmn+j9f6k5lu4DnuzfHCkD/DcOWX6pnrXlecKU4ttaWZ45WRhJbXH
w7RseQbK2PzI2E6PvXxzw5zUM/U+ZtZ5D5mfHK4i/h6uzNuX28uCjteA7G2P
ioZXLmBRX+Doq6t9YiR3Z7hl8qL3LmT48o0vj0bUkJdDyPhgFSpw/rKkcCs6
3nNNmuo89McxeTaO3j+gQptumSEC5Vm8ZKf3+0RhuqivTO2tw84J6aQrtBxc
TbxAP8ivevDZYA3GJmORJLWB4gEqS+DkkFHqsXLloFdoTWrZX5UoeSJzcxzJ
8f/SvIqVO+JKWOBHZrbBqqSbZSa9fEddax+oPAd95Q88veFOxNEg9zQJlGAH
43+Cu+qw7sPvbG/P/8ktznuJnW4RJRuRRhfCa/7hzEYAmrICs56hp3flSZK6
DR7gUVUzOWKsf2ZtWp2+k96KKZ0HaWV+yHCduMn8inO15pv/Sstm5MsWKcci
6eyHR0PVkJMUepeK2AFXtBlg/KKnWIxLghMCh5WAnYCbFV/Zu8+1tHNscZ3f
GNUsS0zt2LjNU7p/x6MJeKa6n6kHvGFPy8KANfCiEuPiXz+C3pGJYbSifbo6
rEsIk/7npJf0iKNV71IH3n1i1QtzmqdvQy6NhJexatUuiDdHb3+d1E/MrTwS
uj6RkJs9KhAD55Qwpd+f4BizPvExG/F1dA2N0YGkqcpBXGgOSi/mT2gDlA8m
yq+CLTCq5KGBEay4GCy2goTX/uGPpN1tvoTIr+i58tnL3FfBsbDugDtk2YBx
wuTvP3KybB70cIG0tgwtyKTC00Mp83DJGnmZglSn7dVJrsBGbQwYQ2GlQvR+
l99tKWlBUmJMNAB9X7iEcMIfCHyLYE8ctX9Uc2cq9zNtha8knXtG9c69xAVL
qR0qbAxL9quOFQroqSQP6M6M2Dut6SGamKsYmnV6vejvW+/KgljcQSTGTMtG
K4PlMZoVimbJ+RZWBIK8O1pOcVlDS209qCdtjHbyPJy6YSGoth1WQ4YhLkPT
Jwn5S8bknl13L3lhxTzls96cO2iXFY60+tNxbnqiidOBaDQejLTShehhr3zW
SLPURVYVU4SZNgKPcrJbMdqHYl/UDw7eKl2KvpA+xbZ39CS9I7qejcB2LG6b
5S7Ijfg4NGs3CS2tq5royDBh8PDOCEyOcg9wVvh9GQI79qG1NDvzneowbOW0
rd1akVN+ZzycZ2zUmBUbvCD2Qc5ZXHPXR0WDuKWR342UcsM0QPj17uS3Cgoh
p0l36diDg/njnrGI+POQ62q0ZKT82b5lxSNvFgejItpTPmNEMQsk+lMWXA9/
V/Wpk2u8fOBg/DXzG3IDvNHfEyYRjGqAr6jkEMMJ2g3Yec6RFPaiReAyVQH/
NhD97rLi3FPOOc64ANp2v0bftqXqQnlk10iLsFtNiWA1Xq5f7tBZT19X7vpz
C8O8uYjeJRrqiDOm2FnDi5keZGhtpknnJjYE5yHoTmHhr4XnBzUX4eu8fT9R
WRXL4wyTLzoblyLvWlSLK6L/ucAUtuXXUAfw2v4oUVCI0LSEgpzag0L/J/ZD
WTPJybFZ09GtzzDpm4RXlNSXFXQRRulIlyM4Na2GOwM4bX7sYjg820+EVsw3
nwNnKdfw2JXqVLICaFqEGBger3h4P/58W6catEiPCazSRS9obSnSS7URe+M9
4X4QWSNnxIIlWcxJLDFx335OwbIxrrjrXEeG60OvONGb6blAqakvlJx+3K4e
0TUWM8Nbspb5hqJ7DJ6GCBHiWM0yauq9Ap/hhaCoKi0w6qep4I4fNQLW3St7
dZ09N/mZFRkkFwxMdLBI3vmNs6S4axcc5v2pl94nxMcsEcPqBAEKyNhaaOii
8f60h7Jx8zbnFuIPDTNLuAQuMSOhUILRTBLM5Ivwrx0rsqhY4Y2M6BMouG7i
HvNKw+EDLYcPLq6nJwibSLHgBhdNFph44ENk3SRPXFFuTwxRyx8CFOIow/e8
kyp6rejmCaZComDrksHU6KXMHqE5wY+qxSrSX5puTvwZxzsNAG+Pjp4WGlxc
KCP3JEiJTB5Urev4XWjDo+hUmg/Pbm+ZcgQIeA24m+MB6DV4pVfGnhaWo+6O
X3shF3x9uzonKZoPSFRPM5M5AKGtsedeCMPZvL7xIy3c5vy9U417de6E8CwM
6a+3UJUduoJcDyvHtckaInRfSu7pSb2XFdqhgzbnD0tjk4FbYi+IK7JnHqaz
06j5nMByZh6xWOHCh2Xqmt6+8hLaRxi5MJGzPOP27K759Ii7m9AcJL2Jv8Kx
thPZDx5dZF2kv4HjbaJmRKnyO/Qr1AQykOwaPN8b1w5FmiW9yH1fgeUO11yn
OevBCQJLOC/wunkFeuqdxaHLNdzLb/13j3aCVXpWsUcXEwfmcWRDecYwLtKE
CLUSW+n0pJionpjB9Re8+FXHOb+0N+1SPvcAzeCHLlwgaVmSXwba5GG/7FKy
GD1Y48C/8BvHQ3tUuHyHybG+ZpNhEC1dMCKnwL33GnngdmXILY9dfv3TIP+W
81sjzcBu0BX1USMOvP22cuXJfo8QmW0r5Jb+dLyBI945Yn7GR4KIFG6lL91I
ci9Jghe2y1QqbjNoSLTxiPLOz5kqvfqbN308urSdKngzorPjYbw59lPSfs8H
PkYO71DHEmu4Xng0ACVxZY6I3mH+e+te2YULKnHD4FifKcTPxyYpmaO9+HAJ
rZXXKwTs1MflgEo8L7On8irXNHTI/pH7aXD0A6PC/G+DP5/9WZ/mchy9vDwM
RGCcBWK0PDpZFV7zLVNm7hwnx1uI/WPM0lMRTSYGvjE9K626Eknwq9KFlBsg
qi/etXiKwUK4PHkC8+v8JOev6FS4R1E6xsmsG+Yaf/AhBeMT5RQ8K7IE8tCt
eCkT+lueu5bqlZPjjXe+sRaiOkRY6gVi87n0OK2lQaqN0X5tvQWqdn8IUC0P
P+VBJPYwmecA0qhAcxcoltWOcqZPMaJnkEkWCDfalBMGmZjuspfwLGhZQs8h
FybQIQFUckSSE8eAKPe0rsnisiP1iXBQ+zr5dozuBW699FVWHHhdLHnGhFAL
UHoyqX992z9jdz+RXCubdn50Zj1gkuClNB7ZGVJ+68uI+xPlLcb/SyGFk65w
tz7qGelMsJ4Db4fRu/sPlK0awsTc3mvjvXMClHaa03lxEi/s2CfQhAknrFQi
MuvAWkURQXfarsBy1sU+to1DUbIabcafaOhA1XeB/b+ULLZqTHCFBBsk/ND1
oUbo98Vns4ch98EAl1iKoJ5haykEsJbWxQv+HqNfsi+bj2JzBnMxsAR4Z5J5
kYttttAuR2cNG+8GCXgegF6OzgBT8zITIofnm6NAcaLR7U85tK4jUwwYJFoq
ITKNbzy4pfzYiKjYEFxQSHZzM9q1rZsFd806gqceReckBWw8N2puHm2WBMwe
3MYRtXNvEt2puLIFo2EV+7ao80d1DLROGpgtZGT7n5Xda8U0BODtZcYfb+pM
StAS3AIqNWAJcurFVFYsf/wfkl/KwKdkaepxHsBrz82kj+hYWqtu98qwV0Zk
TfVkztB/r1R1VOLWv1pXeHQYdwEl21ScohzLumfHfFiTeJ8dRe2VRf0rSMte
ofpJPL+QNayNojvb4Ko6ncMolJ4pxJRseRSXq4XG5wwq2QLCI/NPuxuN7/BW
7E6D7B8aZYALc3lTeyrAGsTNk/FqQrdo4a5c0XtqpNPLnOEhNCgzFTIdItUb
SCD9pPDJawShh4cL2fMbjgFiz3LXMGmUL/uY+/m1yVt64wB3l+OjzFP8Q3Oo
1erm0FlNFaf7A2ZkmEGAjMJTBzH2K17va2zyyH51tqaJ9TFLNo0q0BH/n+wr
vFJznfZIKMwMfqOw19+EcJN0Tt65yHJxutMoaxPT9T3iixavAtKg9oOo+CQT
CE8oo2gSzfIeOw+3UCVLN9GDT2jXqiv3fI6WF0OT8ymjPr9GsJGrMLlNPURj
TrSRyG/H5XtI5nwrnNDro/GmS2odCORX+laLGAMBrwmOjExoeMyP0rE7Xw8S
AFaUyVWcj1Pr/QQPIY6OAwIDqpgpRIDHjE+fEfIhkTWS3z7p9yvF4wVQjNK9
HPMXCgeTeXBrgDkm6Io0MX9rAiSI+KPuqZDU3CgU/QbM4SP2avaZZ/nSBR4g
2OrdNloRNjGdicWMXaEC9SQS7DA0BDZBsC5UgpZnsWlUizeUXZw9JtUuEYBU
D5g9FGN0Lis2JnEdLmIH9DtiyKa8fYqtjeAiXj2gGdYs8Lq88lhEbi0YCgQh
TPKk8zEvoiJ8B1in5np/rIDdvDlVvn9qBPj2FMsS6gR8Y9UD39crZv1d8eET
7dJHm/44as8otWtswLZM8oM/AjDKhgbrLFdF0upkfLj+gGbLFxlBGJFe2Nya
qg7LZfxoNwjZFvBOxCRBIDPzfwSDHs3tOntXxVJDdU6o3Tzfa/fHPwxnk4N0
1FHvwhQvyjlli48Frv57sTUnZ0ycjbqjWrssm9ZIUvhjeR1qZDl0WUaWbwy+
JzWNGXmigbSl3j0qrJmUE7elXUE9F6EouaqRwtHkbzylOaK0UDkgmtudsz1g
2SBbht4G+dF3yRCFHzdzy60JdUYJ649bc8tzrbOJW0OPh5BmKpstmhR3fwb8
fwyDUKo6BzL3MR+Y8SBJlN7gVRNq4958ounAFDP0K/sMeUK6wAJluwfK2yoc
nH/+iz920IHlGLOSEpgjQBAF851g24wufDDLJyq7rgHrRijDwGzBKuj8+byk
TSdoEYZ1EqzJNXkjfVMhdqBZ961BS+8jka/gMXeT3PdwzyavCHmG3Mp5KjKP
G+6PLJJHHkNU+jMTCX55S2SPOI+Mg6iKjMV6hv6xuW1VrkVloJpt9RhvwoN2
fF5tebGhN00GF2QT+0ntXg6RknDEG0gArZzvesgDd3p1dah6tiLUbVx6WNDC
EB7UQOZvxwfMrM7VGQ8BRYzXeyTpxm9IM2oLFMF7F6NPCH6w4yK3r5c40EnX
H03AQlaUvWCH7OLOWlBSuMzldbn1gXzL7p5qgMx5g1WQT0gC8wTkdZum+0H/
3Enj3ulaFWgsyGagS3o1kUkhK7aWXnEdy5q/P9esmU96sUTEl3JRz26AkUdD
BQaKImbUAFiQ1VMR6UmFYOXvZg64TMM7eYlp7IyJD4ta4GptHu6D0Xz/gYDp
1lbTcPX0qXIce3ZhjUshYtQDBsko8s+mavJHnNL5dc3Ed+XsU7PpIjCiLAmo
DQE8LUyxSR2DnFY8vqojNWG4IN3TNgb2MQIIWiu3k2gITO8X4mvFO1+eZJAy
HL8HfS8ELj1nn4N/HSkgBpMgLn+gt8DEeplmda2zD//8fnx7GllmLiBdXHXq
Gnmtlso2Io15f6LC6rRw154+enCQB+SWEc3yCE5wwP5Jo4yh1qwHXj+0sBOu
G+wgW8IY2RkzOYHMarKk+xrbIgl2SR2sc5kuygrxRd7xsJVaAwpELgD/PhMX
HXKOxvmVevv8bI33zlo8o+p+hrZBz+Rro+7L5udKjbMKKZii5N4YZxLiSubs
MPmuiWvJ1nKaO/zsIuPTjnytNgpdvy9SS7xnr5R7RnMtzjqYVG+qL9bZXb7M
OoRVUjQdqljdqK8FUzTZYjYg6V5vnLpPlAher6rtGfWQ6Gaqd91pWOkZ01rT
nwCZpK8oguC96D+XyvF9aDTksbXzEuXoIW45+CZiSDiQ6MYLf4okYgg/EHEO
T2uUzjPGJqyGozscrtYUk2i163VrFwblzSwhUYNQEh2mtlD7VQGwKlNR31Vs
O/oBq4iRdCjAnYxgLINhEQXrqDT2ZzwHNQQUJ+JZbPYIGNlKiexL42d8a9oa
Eosue69QQvVxbgwZ1AwNBLIXDszT8vCrfycv0M1R7yRyColbz9Oh8a/eg7In
FplhMoZHgZ1FT9lsLkHQIsETUhj8MaABQGT4p0dt6UcMF9Z3607t9ws2nHSH
G3o6o2E8tBUUBasDV18uB5DRfzUBd8HmGEYa7t9WPsARLloTRWkQ/HWQKLGD
ztZKcktW4DpMdxIAsRAFSY3Z+71nQeMNmCyWJJh6VWtKBzk7MAD8e5X6VNK0
d+etqm2gE0owQENtXLPhsMfixXHL0OQ0bsswgFFRBSVCo5+1MF2kBPP7A9KU
JZU08dqaR8TGXXgQmZTdLgEq6ucWJQKNa+9N1g2iP3iUMbxmHWcv1XvU5H4x
1VXHSM+LQ++WNaTMA9Bs/aoYzR+VYlpvDGDW8uzEwDCrqiCQQGZ8IpI/iKso
OLV6D8ZG+XGCVSzbAN2dl6g7GMlfT6h23G45MDFuLLBmsKOMQNW2Nx5oVHF6
SUFHrxI61NqIOqVXo5wDnw/Uxnmt5DPOfX5KQK7WPRZrrAJGKPwENs9eifjo
554I0j9SZJNrPERwst3uAbwJovKXXOUyPVA/sB79PuLvopjJVumUWR5yKbeV
OHrygaGAMAJK1y2d9odIEh6ShtfzInPnCNXwYI2v0CeWj6nbMGK/PA96MiS3
AZcGYFR60RX9kJKxHha/d/3gt8o2nYY/tXNMbKcTYJmCFBBRBOSvjxFOONFV
LqZuUO+frQ2h3r+kM40hRcMLfH+0+4FoCYazjAPT1E4SUnKKjuRRSXBJ/EA9
fKRjU6A+QZtRn4etWe0rcYM4+JjmFwkNLQ8S1oKxZAmJno4J9RtZ3CWFWnrt
UqbjopY/L6eb05fuL/VsojhtN440oKwxBrx9rFaJ2wnIlSHmtz2PQ37C/Gt5
wYSFdcrQ6HBHckcx9O9efBXoxz6Tv95kzGlhzgDB9ciHVt56gH9uEteyG9fM
3FCAZjef0GQvie2iEjp0IPQ5te6P+959qqZ9IW698tNFscAdz9vBUPfOq0TZ
9/0J7QQT0fY2tO8bKkyHahs4CrqnRm4pt0W47sf6wO/iNsnB36QF7TRmjXKN
sJMtEVCESIt/e4Vs+7pfxXbGWGY3T/MDgdNZ8NNaYzp1Cej2kmKxwFc2lEyu
B+rKN3Jscnk6gf/5uYroaJUKkFjEW69svZX3ml6lXMNg2JEXd0uoZfbcV65h
k0aPDAgm9eLLbzOTie/PfjvBv2YU9ZemTqi6/ZEX07Tcdu+7gwFxPImR9e0a
VuPY0k9FaU6lIDMbyqP1mKuKTGKNeiwy/NA6c9opeJa90ucgL7zFuc75IXxL
ZY5tafsBhOur8FTulojLHw/WqWNju6pE1eUiKNHZ3Gp0yWiRNOvj64baZ1Kx
MgaDAxPemw9+OL4pBQKUUq+g2ILVue49Qx7ajO8TkQsuADb0AFyVimfbcFJ+
snNfyhgOUO3RFSvhW6uI0uq6YWRhe0vVi43fFjp5onSXiek/5+8QClagQAIb
poVzuyU8KVBBVoWiMAXIRjEKvHZTH4al6XAkbiLRoLCkiJKK+ttnzUfdzq4S
yKkTEUSoyO01yJBjZupgKi6ucBEtzIEiaW5tEV80Afrf7VYwXbrxwMkEJZSL
7v8EMAPBVP70QqFBuaBG/1UXKvWmBLBBeOgLSmitxNl0WnjYpKJq7q4oFeEj
3omzV0XDA4zDcMDQd09bwLWklHnkjHGBvVt2Ci8nmkYblGC/Hmho1rnyZV1o
lTp3rPE7LNGMTbIH3iO1Tn/XEeP3eItOFEphpdElaaVdWtIbusFwGens4zVj
x1KdgbLy8yEzU1/hmB+qy3HRNTSrPQU7xSuK0xALrN9+Ltk88RjY9eHmPY8e
yZyUOtgpyEHw+SwK00tH0z7PT/VfKDzYt1Qjvqm52lteUxBvL+/ZkcNIAZAz
TrKB82m4XlFm0ty1JTDdIXa45QcDn8uXMZT6RFcA4YvFktlZXMr4As08iSV1
v7HWAxbGtYy8jEgLHLumsSwoPrrWWXKfnC2l0bcuZG9Y7/OC5SKN1JlCIO7Z
t385OQP8/hR5NX0vriuEAIxfTa5S39augfFbCVG0iU6DEPkWhiOTfpZOE5El
i5cblcwU0RVMeJ9O2VgjxzaQcRQypOrYZxZU0Ex7SMRRXZabk8sDCt6fkPQy
1m6xGkmQPVVZDtgMrsIw+2BGaZ+15EtoMddzUDC6LYrhXgRwq78FIg26JVjd
3mC8KRRDH/UqnGFeVXY8ZAT/BfNFw30MGuUAu4FMCYws5UblOptboAINY+1S
riE9ZXWqyTxancNK6jHZxn13MliYVJUanD/YyitypQglo2JeRkvZEfkV8U1D
2A+SkHh2fpMjae8Y2AVEzfizzeNPt1gpRRKOZ3vTNVk4IPpaQhs5VK/DYaXe
Tc97lsX6DHFEm1Io2+3FlGAamIIrqqz60ZPChlRYi2oTiyrLB+8bzAsHv4Bz
qJcMeApyiMPnmMpLy2UGwVRxys/ciF0lS3pIKQBB6HFQRu1K5JEmhOLoqTTK
dv3kAsC98D6ierS1cHUlXGK4cfzrbD3d7aRsBJwiDyz5U5AFD3gOBPwNk22F
N5BWaDP9SWRrO/wcXwxDYBvB8iEjOMzDuAh+5X6LvtULVQP2Zvj3VgPMunNt
XpINYjxkyb99f71DHRbcgPwOcZ0WxXl5MT1teS0+s9pRhCkclscfKRI5I+HG
3c3U6UB67Iu77qFV4QUPejAEQNArupcGuBwY8DVliuthnp+9iTXcTivM5woT
LK0TSHorv9TNpffGKRfYys/DGKqQ2O1NurlAjnfbNDnFDVrbWDjozIPUiDLQ
NKIgByAcSir44NDmXAOT3hVFa/KigtS8rmGE/hNURxBOOENUAVJZqBk2rFi3
OzmjdeUYXHRjrJ9RpMipTbcr2k4xYzVJ07Z2KqpOyBJQ8ZtE7E/1KPmDaI/8
UurRzPDQF3yWjs6vfOiWSWT0pcheJGIDCJHe1edizn/ZA2Myz/iL+fzKpbkg
TNG9qIKarH7dd3zP3KC6m4Gso90eLIsMF+qTbwcKXF9mQzNT+7uzNVmeiHRF
g5pTDGf1pfh3XOFe9kRKzIVeLqhpmjXcT3GBjDmwwwBVs1eCsMoLVxzG9zzv
h2uUYPAkY/Qt2g2f9KRYXszuWQLYRyN7gYnXSw7CbU8gYqcJUCmAC4LWPfs1
Wne5gi5v5onnqSByG6NUmXbyiAwxMDCpGpocMXWqLKNu+KErTHvDEtrX2J2v
+gkraVmizPY+jaFY3dOoW5cyWN3Qizt6jyNm9vr6A0prwy2UlUssY7Rvg0oz
s/vRGbAeraSU4IhUXiIMIAgSQfrIyx/p4dXHDdPzHFBah9Fed/ALrIOuwEKp
L0icCYap7+oOoWd47as7qbebSySVDEsF21QxziADHlL1qxaFlvw/BIcvQK6f
i1hWEVnxRvthwK9aRNocFiBQUFXQH4wBDNJuVH1FqQCaeQZJFfbxkWYwjGUZ
2Po/Cc7IFQlE9YfvZ/Qaghcstbc/NdFudWRLjOd9l1gUJmx8wKUUXEVKn8HF
kDqkJphIP4psdyHeyWyN8BRCa2K6H67k+1TO+XbsiiKWTFUPT005nBEy0Gkg
WeBSz8V4wZFjq/vBAkHzvDAuSLwxHp/qC7ZeJWb3D1Je9UIEeUmlmIrkScaa
Byt+d8QL2LLDX8SPSjL6EIQ/aQ4hhx4xH3WBrF6NsEi2oMaeAjEJhhQeJSl8
L4+JBQgOiE8AWo8VXrzF8y8vsW7/hwdaRkog/ozsJ4SlwLvMRAMjsHDjww+M
Bi/YuaXXGc7F6snijzQfmILgbH/7peikFpiiK3up6/FThaZytw/Uj9iu/943
MFr9G6qPrgff4/brt95eo1idYfiur1CDZsl7fAsNWQUN4RF2ayaCUkxhTcR+
30OWMYrGK755XX1b9vSpfVysdT2w8MqIw9gkWXdY9UZe5F6fxnaentl7bJVy
HL8WDYl7sW16wdw1kcWuFXS0Tu2AYyIYSKKAWrUvge/QLdiN0QrZBUHRDz6k
B2n8DGPkEGIIhTHWykoa7DF8yidNnAIYYYQ973BP+rjFLnDuVVLywk8gwDmq
Sp+BIciWqzwmemWcN1MyzncEx9B8TTEt6OTkrRpE9hFn54bhHpgiNDsonRpE
XpI6Y51BLiTfG5L1jpEHtufRBm0cs7aMvTj8cOvJ0lz9yCcVzcjidCUduPpr
CAqOeDQuEz4zwAAWbvBRHjI348xCxtrYbObcEMTYFhaf0Y6UOvTYDpHzTkLh
iopQjpdUz+/49FBMgtaq3Q2xJL9rUZb2zTdbWwRNjMBrxJ0MK3jupi97RWo0
/TJsmL0TLljU1TfyKwpYoAjluaBTsSmQATH26KMm1s8Ve7n1qH+1XlQzQnGn
utSh8Zkk4Yot/3XCXGv8jMi9LUs4B4APbvZnSfEeh5gnPa09e/gKNvA9/bZN
zCqrYNtwdHWhXch6cGdI78MyFnt4pjfomAdcVqVaK/KHjHjyMaPzMHzcLFLO
EpTkzUQ1Xs8h8k1HIWYlDhzKY7E5v9woHH1Xb/+jYkagMRSEeTgmDTXxMwPH
Sur8qwx2l2z54Xj3/xZUKebLQTgBwZMFPcHG9xylmVR0tRZnNnaQF/ATCXW8
KG9det0jIjmHB1RIsCOP2DPd98xmaq8Xuu37g3jOc+CCee/i7ulWyUDgMGP1
V8T7a3B+XSJR8vampo7Ho86roFrpnBV1PGxXxi8EkqUMgAiUfkhAl6YGhNr4
oL5gHD693Nl8LU7wZUc15zhAbEB5FeVgO2ornWV0ngsgNBTfqkFidRBUI6xp
kIMb5qeedmjlqM0LVmdvaT/+68LSp9WRUrYr/AISew25Cn8aD9E/pz71lznp
AC7fR7ohIOmu5eqLybvJqcjA1WZeKtuILtVfmY+9/zjdvojqkIPn78QO1Ccr
Bm0sC0/+pqRXGEXYjFLwHyxOZ5ol0xtQ/6X5hWFBWtCIy/CAkc/3At+6R4RH
vNDlpChZbzszbChsqaMh/JpvLrKv85ze21EALv9PN8CJKXId4YrdJ4Fkb8wm
Lpkw8GiuBPt/zB8Zw26ksgzZI/iz8hdv4yxv1o2SYkkktRGHJo3PUYTuWEJ2
smrXKkNRHhfGvc4w9z9yRnZ3SNHjDYQFebDOZQEakOArSKSGDmTaMnh+MsQH
9JWsGtunFd8+fjO9We7gYYAmn7LjcdB8bXYr8/mOglA8RYv1mAy57pEGbtlb
p9Y+x7sa1GJ6nNqbHgB9srxqc3EpAFU7s9rTgo6bbf7E41Uwk4L9sN9DWAzb
sD8nP0+jTjZ9qKBCFX4rvtIEDuCzQ2ArfVO+iuZl9IPBhgDCncUXYROVdz6v
rtFSzFEKJtYwq6Lgcekj+/Dh8TUb0SYhoLk9Yxnj3nX+MDkqUfixS5+yUQgy
U40fFqVYxugn5JA+Sz8tPZs9q3XVGMhgZBpgfT8Ir+dD6w1hri38SbkVH/8m
eL8lH9xU39nzY2JwMG/y7NoLlddO7x0nN6Fz2o7GsD0myxVV2heMAUh577Mk
o8uGHs+I0q1JhdN7PZNwWYN+TfwMTHxmOikvIYPM1/w8vBIWZ7T20GxHI6sk
qzy9SyxklZKbUaVZ1jmlU9rNk52pQySZx4QxiRrJNwejZUIuv4zwgP5A4+vZ
MAbCfkdrDzz7YAvhgoXByfX8shXAMez1v7zFrdIupxqFj/PDKAcTEyElo2Wb
ur829TpFEkgJqX8RnqFQV7ItKvkUA1ztXp4NtOT6ZvL8Ob5gnJNcggFS3jba
mcRLUGhpMIK4fA2uhTgrLwXQc/23jw8zUEvF3RC3XyOchQhcxKnNOdb9TGx6
jPWl8iXC+9/AjmbZkji9qKmz3g0A2n1XwXG8yqxjZbgqEKwaQFq0ICSGw9K5
RqrfFUUvNR79rd8q6jeyqdBo164p3EO99XWsiLLoVm2jKOMWp3B0z2KhCIeL
rABdPBM1ObrHP8F2DCRWkXH2nqZzNlXhOQp2wcjhY3ND1X0KtwEKNnvRDcW6
ukHVCZME1xZ4xkfVYP+Kw0kjXSyUfPfy7hJyugQ4uSgL37lGz/I6AwwzUG/U
ARt7hKdWn2j/W63wK/uDqozWDMSYnSxzy3Mg8cxsGWTgnLisVgX32uLsvjot
jlraUndtFMgdDBg/CW4tzJdm04AwGK8iyC44nUKmyRm3Nm2/PNmJ7M6S1byt
dXasjGfwGEsNLae5hJFYm6P+/xBqIfMFzqS1HcfLZRCWKYMiHFCa4R0goBsl
8QDuEXXwivze2YkOEsQENpLvJlOGDZ44MWGpJWna+2MiQDRZfnxXWAd2TfDB
qZ7M0fpzR+FoM6xkDAP++H/KDVBS7E8O10T5tqOos/d7/qa4lIJ18Sh5tsYY
sZAikoaXL/pI0ioqEnhcfJAz2WOGTw03K2a5t3zDzSew+XmlToPgqNBylEpA
ycLN2Q9nxfbsTeOczFAeL2jKYWizcIegQocFB09kS+G2E/n3RNUfc5gIa66G
Pn00oJMVXBS1itOzvaILHWHTRzH9QMMfJnRewnMbgQxTQzLmaxJw5wvab7EV
WVHnPWa9tPH5uR83k3451Q6ImuB9qKCcycyRqbSk3n4DBK2EPE9p2s7O5qc2
2ag8sR9IslA5ZqjuwcIF47/Y+O+0pFeQHBGspX/WuCf/jS8iwR2vyYp7fiIZ
pIAIRZuWweAXHbMU/vJBP90OUt2tX4GF28jIvADUvLZPqo6UnwzROXD97add
CvYqJtqITRm/ACYoYLFVmthXqBBuDVLz/5bT0VTcKDClg1xAeErckOBhesUw
6r49rAvI6i14JB4Ec2WuEzYwYUb4qGl01LpiiMfiPmxWKzpNonT3a+EbyHhb
EhYUtklgfuP9eHkwBVLL2treoFuAMdFPKeMkYAUSZEPd/G5lHTIS7nmBbWsY
rklW7CnojHG4sadfLJwvul3qEbBY6GRWOKGzG8Z6gDjF19gZlHBKodm5jpY9
Hwlw5w2XUS+PxAFwAVd/y6Lm56HAfA7XBxaRDy1LXTzirExk/WYtuhr+sGHB
J7Qh2+sXQeKIhRnENAqvEmZY+DTQOMwKSyZf+7vH4yWOmVa7JYdtTG82aQtK
1IvNO9cu5km5mZI/2LlCbhc2w4hArBC3x8RVdZD0Cf3TsrHXaDzYdGUtZySL
gY1/m1XJAcxgSrkBDhFS0mUuhOwL1OnIlhEu6fiJ9Q5JlfM5pMycDhuNaUCU
EDHZXhHpk6ucrcH5c2kFERVUfgn4gjbvgNfcAvURXC8Jg97BXcHUJJh6PA+d
XLVUXJijmmshjFsvSne5u78KnOtF167946NeIctn6gwW1XaQc6WmsHVB0Qsc
l13dnefNM7R5Z8OvlOxRo9jDXOIGjmnbO1ofTWSTzLahXGW3KFcoHHqCtd6Z
u4aCz8rSDkyfuetuPsDuoJZ3IdVG9q01X+TOHg9pVSgY+68p9MbJOtrbvhK1
0/r3atowBFeMW6JqXNV6UfPLqRPYZJYQgKNb99vI2d+bRQmFUiqtssdn6Gem
CntyKCpJmBWT2Awd2VU+8gdHxSMk2yXMOYnItaRLjj7AUFmY/P7V7V9cF4Hj
6m3lMHpgj+NMh4mmgHkn/8iZlCvhygKsCWJ3SKKKzSRic7U9rlgQQaFGCRWM
Jo42bZb0QhUYlJTfTM6RDJtfE+nVsyj4/9Si9IOWAoRtaeNtq9F+eqUURRQv
SjlC/RnJy2M2xsY4ymboL87dFXlSaH2tCGM1shUDvopGvVpZRDTDiL0SS+75
BRfr+/slhnv53S3XDqdfhicu2ZV3xM8KMCHLm9ZsAo+dh0f+tgM7QDCYb5VI
Ri5kobAhBJaGnriXASr7azgDBDaoLMc1KRQ5L4Cm5vXhCEusxHg6jADRVmKZ
ygZy4TC47EMkWZ8tQcZGZDYKco3aU+HHa9+knGT1Wvdt6BxEYdlkw4DMNriY
kgpSo6B64KYGH2fVbICopjoz5zWzdF96BB5zXV0btrOqweQqhcffWrzM8T5t
5X7GVAbE5sWW0gnkinFZrTeGwT8Jo1n6Y0z++dNPNxREU5O0QPRtms44pIa4
CnoQ4h4P9wShpSMrmSRkwFYkwjRlEZCDHHEISAsv/u25m/m8Kft469W0u+Sn
jim0XO2yfFyWD4SgwAR5H5RoP4PNfENho2rS9poh+6K7/lB7rnJCtEE6i8bK
NnyCZScYExaVd+7+t0YmRN/viRIMeHWGwCk7F6aKlbZsP4I/lgN3ytQ2uyvS
TauwT54jChlan8zvN7JXNZQjgJ8Xq5gzvNAzRAHbrAORmlNlcWJ4KHG6YiBg
gqnfZVvY2+eAY33SBf6bo3UbDY4mRg4ByebhXL4V0rJ1Zadh4wbw2jVKWLlU
3+1GlSpcXoeDTckx+UqWNYYosvvV5UaexLmSmTSaZIkj3PXsOLW3Hnm3KrhR
bBbPU2VejAKHGDxNZvm/ZiB2blH1WHq/eiKC/CqC4jZpfjz+Pu5FNHlot4NO
t23hkdh0Lb16wzlwcpPbbEfG8LtHK6R32s0zYYJq5/dg5J1Z6sD0Q25iTqSG
MyvGPS9rbFwBRaFYhyO1FYKTz0UDedwv72OzuU/iSLUe8nz8w0JqCyH+fnk6
dnT680hh8ehhwX5FmvS6mTjlh6yt9nS2ekWStytFsu4esNjxPpT5LP7jcxhq
GAFOucuMu3czkBmAxm84/NpTX+1c0DoUd2fGgFtlSM240E/vxmRlw9iPKDYM
1Hoo3jGdJIgr8EJ2/FTfmpz6joWWGL/x6cVeZy7BT9dag0nVhyduhFoh9iSB
hiw4fYlc49zqhe+V5Z7CNzXFj1LcYeTB/aqQ6Z0vIzVXgbvoXJ6fg4s9AnQI
OLYV3RoZj57BJ4wudzNGkyLpIAfZ0RMXCIPKYBFldr8BxMWo8j20hOBzuu3d
KrVi9Hgw6Wno+UUwTbp6L3IHaZPfPLiAFdkfrbnCt1XdgmsXZNApTK1VF5/Y
7qcHo28flwMX1HF7T4f8wy6Twtfv30hxWru9q86xR+5N/mQtroAf94/RT6ho
usObippDw81jHjkax279Wjdth3Om6rx0X+YArkDk39Py1l6F9E7d8KJZ//f7
H35CdMMtIDzTW8IWqYLsSmWAmCFqbKu46iDONdZ9EKKiOHoXBmpwnDcT1nvs
X2ur5ZU8z5/+HtVDTbBSKAY0E0JN1czh33xCdJdSEZHuqBAxSuMe6VKYLJNz
yuEuS7j5tOOAlddada/6dnTkOJnB0kFqxpZA+44DyQxozUEjSOoYb2ZALvGu
eTtSxyO0vNgiP3+9XYTqJtf5ojVRMoK/G7EqZVlurFDsh6KPSpE5FulPAqMr
OqLGl9wd3pnKb9ZrtKWMWytUECSkWkhiBwXv639yplcd7djivdCHF8Sgd2sV
iJEmZDJGXY7/NHDmEzkTICidXXo3aszl8n2HAUAoLP8CyMK8VXyTT7myZTPL
dAVlHX4wwijCydVru92yh7XM5RqsN5C0325DnJJhJqfe7hBxbcSu/mZWSsxY
7mdVrdsENK7/LN1XSHbW7b1REc2QEcv6ZupdX8UbWuYxh0E+38+qTanWJC1Q
XJzAzscHDhvAHo4L3omXY78uop7UBkP6wRncbvS6X92GCrOB+bXzCkIYtYRE
LmmSI8tqdvbCfyinZpTePml9rAFaMH8zJh1NgJN9jHQjhpYWTa/FB/RmKzuv
TdjEFrJ5bmuKefefNhK0Md/JwghlrbTvLfB/LX6WhEv58THx6Iq9vfYZ8DdQ
qw8hmISGZzmgTpsqFiSSwFOKa6R/urotcCUCt9e4FBBpQ9fKy+WfpqCqQVtV
0UlnhwRrPAxuyKHrN6FIdMPxujZ7yLVX6Sw92pSgp7qfpUqaDGurooNptMj5
aWh8sgqajbPYidQPnu2pKDg6BOYVIakh5wPdLfmOBW7mlM500wFSvX7pDFyF
G5plPyxtxYpaw3URpuodBGl5f3If5xF8KZK1cJP8A6RLK98Zokbo/HiMyIio
7VsapDtvxpU9RZA3D820IZAbPq0n/HIBcjqdhVqD0weg2lbaoQhKUJUQ+24s
0Pq3n1aMs8lKmmLUUuyFQ+WB7J0KlNBxXKgz92bsDhFnUtgFqzBaPtqVTCN/
fdGuBAg0N3arAOI5yywX4LSHghkO/UCvhSibqjQFbykFinBFJBRqBfZE+wKv
Z/ky6aB8vpIhnybP8rUzoNvTh/JH3V/+0ki92A9iCxhQDdjg2Ui7dyxih4fG
2Fs6o4tufA+25a0w6mhtth3hfDbUBBUYIFQp/MzcchsNksMG1oI/ER01gyL3
Xo87+Z9e+BNaAHjKBUsQ51dCnGGyCnPcQvp8eSeIXvsvZXMLxqxXQnqKDgPi
I+YwG5Di9AcosfCLCihqaWc2m+OJPNLQACY6ygiJa/EmW98Nqxz1rdaHoltK
qmm2SaO7+3dBTc41xenIIbJ+Zmqok9ueN7CWlYTAehyQYqZBBtW3dM7BtuZb
2QQGHyhCg+M5PX0gWIZK91kUFD8KAYG+i79fhKaUD49LcnPMkADQQ+TByGFO
5EPZn04PzMWhNdxA05+StOJhMBCiHw7fFu5toQFiTPyG+KgHJ5wKmZ+v3TuZ
zaWcH19rpclm46Ao4m037jnBE6liiNkFMW/wZSqNkk1PsvEIQop4FnptAhkg
2Cf3SjflCo5NTrxk1+k7v4oh9GN0abSWA40JMKhZX1XPqbVt/K5xXgjbSh7J
jRB025YulTGbQDHUTiunCTd+8+uZqcGm4ie0inYNzhi9/8TeC59BKEjTPwQ2
AHWFOP/Xe24DzTIaPcrBDGgB52SW5FjGprj5YYIYo154LkRNjKNcfQF16oEj
4x739cjEqZwtritegxNWkILOC22+DHtS30n2aPRM7tUGpiYMzVaYprcA9Gqj
Bip5KQiUcLF8IHzoDmcrA0FvNJvsib4gxPB1nJxh7OZ/5O9kBLgn8HlN2hWB
GbxJlbZjxB+nRFvOUlr6zuBXzH2mZ8HEhzjsdVsD2eLmKpzZP1A0KK8+YKYQ
6TUObF25/VpTx5Tw2coDfUx6dyFfbpJUdmMBxa/TgoOHijq9a1jBfNMLBrtA
eRx+rgdLHO+9TERLTLzLp1emLC4EEtDIR1RHgQgeXofUneHy7i+pBnePPf6K
nUVDgCJXk1zrItyITrCSuYkv1NOGAM+SmdlHdEEwwsIijzbzuSZvYfIPfpee
IG+gvDuOxHzHAQfKb0eY0+Rjlwh1XiysFbHtkcgkkdaQZ03+RJ58ar4e3RNB
83d8mJ8QBBN5+y0eGmYlshhdUVUg7eMNauERBs5xy+I0q2EU8fYvXnliWRjX
8BNstMdFFFeinXWMzy4RSnyc34wvfPyuBfTec2/eovm/cwdxpZmZPwPY3/xw
oiGXCvUjVi8rbSkqUGD3RZZYDKzp7yQTwal4PsGTAK5s/Se2ajACBsJ5tAfW
2H/d0n6ZUlmOmini0RHnseq/S8GsiZ/Bas20JGjt6KUIPTowOlzaR6+YKGN/
T91MLXwjIN8VJPQIRsDbA0y4tyg8cF5qWR/nVgubb8i1NAA2fAxC6CcVSll9
887256PMc68fzLRhPJZxzQ0SL/ABnn9Z+qT+yuNfQ7CF3+EuMfFgr9Mc5F90
awhauigPg7pVwXszTzdK7AM0HtNLAB0UURmzMB5/y3bwbIyhyHizAmiwb62h
GDAYA2C1ufKug5dlUrUzHq5S61+k7xo2q5+B/Cn0jOaFRbPWegwcLNLIh1Dr
E2QynIeJ8ZOyQjV+LxBcHLEE03QWDpgzKOr47CihU32RlLOxZ4mU7aBS5gjx
bH2t8Wfro09JZku0q2ofoGkZEQsU16DGPY087Qf74rWyDslNw5pjRL0WDRm5
15pUlY9SFo9ST9fin87UXsyPoxlDLV3PDao7OCumYrvKAM5dGSfv1cLdsn/Y
w1tOC7DzIbhrGfAYIXrhQnuuZmPgsGN3tKgUmB/6DTOlSvLREkXaLFUOkcyS
FEDqQ9SEe8YsN7dYAGouDR+emNcNwqHnpeiOYZOJH4EWycIB5+r2UrBVgcq2
5Ny/FT6uka5f8QuToRVL2sBJQYpQAWsHt0Dt2Bza8YnyW8cwklSGrC4eNT/1
2NPLoY6c+ab0o8O4tj642HfwhiGgWqsqYV9zschemXLpUMrQthdCE+BuxiIV
TDZiwTILwRQIEfv0Iuo5PqhzSQVB8YaYvC/TihMzOFWMqFF7fsoHDCH9ki7o
fvV1sMryK+SMrpfucVhvjRtY8A5SAwkCpBSF2TNXSy7uh/yOsd+TtsuH+eee
Iie73b/Wd5pF5h8KOquR1lgBmovOS2sEQ5CXLs3pqejQb/j/+YL/711RdLL0
q8qqBPBifxBD+IJkC+ze9+rEANKcrq6ptCBOY4nPHCt/5GySvVf8k+WJ5Hvv
c6HSWALXbxkPprV8dXnBXBiiZa849ntrSrsW3EdG67BS5b0Vt1ndHTHnHZ4d
b2dkFbF/mHZZdBTZKvU/i08q7+8nmPHCaz/O17iDj0ohMxheF2UCsxJueG0z
9N5em9crKhSt/gPGv3c9ejRDdkdqqXBh2wu/BUFOLXENcn5B1JbsWmboddhD
6nfG6aRja6Hay1DWXTWGDRWSJ/0osCO3/F5OYdrkSk8Sq4ftQ2z3QwZo/4xj
ojOEgOSmNmYWEIoW2DuYF4xRsh0FKaddVvt8xqzIJnydu8/RyLqT+7ZV7Xfk
0MfBstPO/3ND5yKCbJY3d8mIxT5KLPrK48eaUuVYwd8qd+SAqvEjE9I3ac1r
x+6nZQWwLUVY59IDI5evKDf35aZkt9r0gs4mqvFvxQhLEPekOyJlrAdfD6fu
0755eiwJqSQVvZNADVXjUtU59BQ+hFxcC1xBa9qGlTIUxuYnqWRZXJhk4d21
uOS3lONBON7mpaUhNKSVAcLc+QXkl6B5D8253OP0huKqsateBZtRhVjwf+DY
moBIuftiPwGdKoFb+7mBvi2/NeFRJOYM1/JcjJi9mQhboSqndixMNv7yGBqG
Z6bH+P0BvrIsNSw5UaF5u67IeKDMdgGBE3LXyzbsWkpymSruMOAUTZCo+0zO
Xf6xD/gzYKXOOiK50oPn/2N1GhfSVfKrpOogvC/ZQ2kxekayt/RFT5vLWfVF
1Zn33HxJp3QpTaNM7401ENDUf4Sawvn7l7n5Zo/Tc2mbAWHXD0Kw12yKypoI
aafRy7UwpDDE4Dp1rJxLORwSuazZieM31AY2ucVTJRDN/hVs/mnTS7E0XsgB
EV1WHUgd3mTdaUOg/NZirt+/qWlDCTeOT9KQuo+RkV9zEU+y+Ogxfx2TdtUT
pHwfUrGWMVKddWZNFRiSteckcxHhtNy70+uurwyCy5eeJr/8XuakIgBRaDpP
2k5ASPZkVnEpdUA/uyGwMhhDnaZWLLEUtJc1npn1oge3tict/39tLkox1aai
vmKe2/yHvkXfOSebNWUAMNl4zTcCMSVLnJx+Dd7yFr6iy0xJYD7jQ8I0oUzM
+9m+9OKIjx/erOYRLb0eEN5r13ehoFRJf0NREjFhcLhcH7+9CIi8a1BhrsIX
cFwmPEY/pM0VarPuoMLDzJNB0mRzpg7fW4KvC2cwN9SzykZOEJLn07bc2i7B
fIzv6zhtKW6TkaT7YzoALhSDKNitpdU49bPa0TOjcJWoa8xH9WEZZ/W3OgdC
DHanFOd5M45QwlVBBJ6LHRQqs/29OO9RLBhKHygKGR0wH/21YUEOPIxPA0n8
Mc7rgZnLd/Y+6mf2zOvqlykRUOFiL+92ZnsQ3Xx67j3R2Gw48VDqT2sWkuTr
0Go15wPV5JBzog3Hx8dfozzKEncjKtpQDbrxsFscrqapVYgbB5YHm29HQ9Sf
emXcEQm0KWsGvRqZo6iDewVHx2gNn4BFktloLDcU6QpsVyfL26zuj/lrXlyV
O4rq2nqK8hXYO0RhiZ1s0Pakxmoo3ygDlwJ73VRu1j4aFkMffjbapklgRmJY
qsglvJaZcfyXmGVmzjVcH1B6RZ840Y6riwWcDw1T6yw0wk/xLkMoM/VGCOzM
InJaH41XDzmDmIHNAzXLFvPS4RCNVWIx6sFvrbPYCZJEbpNV5+qoiEOCMfhW
zwwKwCRbQ2wzwZjbkHfi9nbRvxVCuTLo3CUwmhVVJbT/MmetHN8x6s+b00+C
BFEBcFFwNqN0Q8WI+6lRnrm6FqKe4IunFr4vzylrhn0mrli+I23LJg/agv2E
a5ZdTpBdiEh1lTKc5MnbIoBowR8AJkRTmHAtoP1uVV5MXpQ4oa7ssmEV5BUA
eQH/SmFL8bF+V46H4HoocxJrFx2YOWnu7fb79CZ9kw2Sluyn0iKgN68VkUCt
QJq0Ip5R44Dvk3UACr+44K43wpqYWn0dDslIej7enukYZxsQamA5pIeiNV4O
c0FiCpKuMCGEKduEeMA7XUyeD20dEYb0ISllAwLtisKZQmbQWZryXjan/G7B
wgwk7Sk8j9mTfXOBm24c6fnB22u+G/3vWgjS6ssEoF9ZLmJ4YrmxdHobNxtK
XJ1Ki0L8Vcg1KO3H/eXQtX8HDgzWUewayE0sNELArOuRoxog1m3ljXGCvPXi
xuEtzBjaDicICqqt6lyk9tGffCWIaDKf2H9dTfpMcKvGeKZzSXay/oKZqu9e
IRbRKp4tCX52DEFoQamHgw4kH/zSm9ldgAhoVidFcNTLaRfMVEFplhKtATwl
WcO0VZY/IwGfir/pW2zcwTPOJ3KSwpEaOkSoEU+XYKUtvwP84DLgEpIhNQMi
50biNo0/rmIoaJutMKJAPjSYilW8dJ4s1axfjQD+EKEXBcuvpIiGuqkCfsEA
QPwrU2uE4jErsEwy3rwBhMyQcoqSkxFQJFoHqRFRBnvPdy9Cax0kVBdT/cnU
r+7ukHK3V+NwfpZaxYY/XUWYc/JMAYdUHKh0RYwMvyUwJwSrqFOLAGwN8X7x
KkT8vVwIaySZ6oA+wHwrwpF6T39Ajhy2wOXntj1ik7MRcTHd5C9l9wtUcRMU
6Cn5y3lwz2fimc1p4HuT3CNqvA7pGg8UhFu18NsKRgaoMWqRkNGn9+ticoYa
P00EDIzspkb6727vr86iNsAm5wECRM+O2FU74NjfG8aJ4FE3euWfk9DS2VoX
fDRdSc5q9OYcqq7VkCNTdvTEadIBrSVqgQqS3IiY7RGYfcStjoPlJ3L1q0HT
AddXQ3Apc941N6JzJL6eTcJXCLf6hrfM683n7laDA2JeP0ceh6bhQfRzm7Gp
WS6SWoecRRcm516v/Mvu5/vZ9iv0iCEutfmGfG+uWdPQvMbt6bSzG6ofTehu
fEnED6q/oTMaNR1BXrOx9OcZXVRA9/TVKnn8eDjxWy6lhxHFfzX2t6qW86/I
DvVVvJ+Ky7XeflIb5kHll7WFUtuiV3cE4dUorwFvBhaeqP/E7t1206dqyAol
tgoi6NKqR+4DjkkMs758DADjsRldkGvIutkC8Lj6Uk+HQjh6KDEiNXmtn8+z
RiZv50Oa6EzojoDWSl+mN5ZrfgnsJT73xu3Gls/y7tdfS2xPhfO+QL4MHa5x
f54ls9gXi8r8ZoPu4UGJSHhunTISK3+IBK4f2YdYYN0P3393xHWM0b0xDoWx
umu9NA+OxXKgxc9gWKgU3DyvVfGAOkliJ7faL+Axbu/+oy24XdPaTEQjDQ84
eJ27BXc/bE2L1OSU53uGGD94vdnZAZ42fkrt+h/8pfs73pIGjzCK97OMcSXg
ZbPDGU7l5EVfkBbHypLFGATIQxasBCfecSSI/eKAzHG/xO0RSdk0LxjJsrzC
wlvKwga0efoXW2+Bzccl0pBxKIUHpYJRLwFWitI9bKHaTmLwDIcQYUOTUBLM
X6ukbig5GPOO/I6/dO0T3BwkOcggGM/FeuCHO7s9JUNVz5akvt0h/1ix39Ue
yEwAKkIfBKjwETJF3gzrDq0oFFLwsyWbHqW5oIXYN0SVe/JTMP6zkhY4CDUY
qozD+ABOgzG68C4a83W2s4PHqtp0QmZ6WpTUU/SaUqrDL/j2uyNR6nxxYI94
Wi2KoxY8BsiPeOXUX9PvGVCFqGUH8qyQ3mD+neGEDMfUZUE2TT+9VAf2N1N+
6OaxBwg5dg42d85FaENDD7Y9HLBJISCD7KKUyUl0N5pRfWQ97SMtl7HtVzlC
V9OSKT+3IyqH9Mxtn8COl9h0ouq3h+MwvVnZ5PLd0iEynK382wPAfGBrLZs+
YoMXlR41Ub8834GtTJ7TYgMeP1PqpuzJID52HpnBcAW2gRRBrFWgW31YArb4
bwxkzUIq6MhkPT33h+2epTvQ7WIUVuOA2HpM6brekQl3W1MH7tn2c08TYeur
lauTsfWMh8QmioHQykcwAqqd3xT1c7JIsxAN2MrtbOvPX0JE3LHs6NQpmCWw
S7xx9ocAKloOlB8PStnHEYdAsehFj1MeQRWC6RMrv0yd5r6iL/kGSPGkbmyk
b9ffME/5IelqV0MlqVMtNUzQW22ve7pcA1D/uO5+VfUwv58YVGgcFORrFVfd
GeGHE1IpQ1a+FPopKXQb2vn3ceEpbZVnquapkGyPx5iPW3staeLljZ2NlKSh
PsRPk7ObJzU1VRAgak44S8oo9H1ig0nhMHPWAwlm+6CnZi5we+41yjiy5UVe
vZjn6ge3xYrWYUs6r/6jsCZmO5PDrHdoO5oTCGoJqqqLXBfZNoqKbiP0qs+c
UqJQl5WPbLoER10/ZHUWhp3rvU9u+Vbx3TlnP2T2kfjGo8l0gtoqWqr4hVcP
xPpRcRRVdxKq9kIel+e8WiLMApYem+SYk9/2Rr8YtTXqeySW0VpOhM1ugCcW
5NjvO/pqb3MgTMcUnFElZ+134IXEDbQkVzgqCKnZoYo8s+/6/ablEGx0ze3e
vv8Szapx79TtRgqQT2xb/zkl6OBqwxlHCIkSPPe1l+I7WLmvIukOQ5RYMWpv
d/KIgakY5D3eIdcaVaZFWaJg/sXH/3dcTI14AigDd5O9lIFrvO+DnGrHVm9X
mJRlZiuW78tnq1Dk/cR9+oYxSSqVOGPyDn7Ku2Fb5PVViAREwxCX1GrO+H3k
jnQnEg7DHzGEuefyvKlTt8qxxBgcgTzbMvaclTGAZ00837ccjfTRwokmTC5C
Gh2AtWE7q5m/Dg2nWhhhGXb1FkVuUOV4wiVLXwVU0A9KYj8yAbETQerDZv+y
JFZTY0bI59scJAZkQpnRtkHnG5Qew7NXJB50hFoM4jDokMbNoVlYMYOYQMWX
cQddUQCw/Q96+rtsflfxHTVvT/FAtRHxe2OdpnvC7zdH07wvlNYqxICnqQpC
VzbDeJVtgPI+K+tiBYGmvNbWkEDqz0asyXFVbMWZUTcBoq3oA87aPfRICYoA
4lCbSGiKTypiyXU8XNbUoGaxBMmgnN2PlCVCBKyMRpd3Ga8W6Xg0y5XHyFm6
z8T8MQlpRit8NLHVtG97CfRIt5gxCc5yey2MX3zRfn0gygTGkOplHqdD03jp
QwDGPVxwDq7ds8UEG4wamVmP3+j+NPwe2H7hhZcrjeH3cpqsPN77VfYYklzo
dKMMwyT4GtkP95P40WyiAmXZUKFB2bMIeEwJdyow46dqg2bp5w+j1dhAdvh6
hjNvgvdvx+dIIwry0ImKK/lZOeRsnSJIU9zt/xFuNrShfLXdx3/nuxdwYzWc
46nD+UzYnKJmhi/VFNKiS5QjvOYn7BCeCiUQzmIprZwQ6Ep7pwDWVBlet8mx
jzowdzqJR2Z2hqAyN1pFNIkd33CL9mRBowmoUdqZXuUFJhMlYUQKuBGQIH/o
EUCwIrF3CvYPhUQjM77jPk+/gHes96xsABIB6U6wH3DS2L8+k6xdeX4mwF/u
xcIV9xQhb4f9yWoIoZbgIcjAgMb6BXVt6MzxBAJLiZhLdSdHb5Sk/tru+3fa
j4IIGc4RrTYRT0Z7ZXE0mOVpVxxoxoY2ChFvfgfq02pV1SS9/H/Ji3ldgd/i
lfJMZu8MeLZnUY69Xeqg1dHFik9NPqVxZoNZJrrrMQrEVx7fdzpy+oybJM92
boJ80eEXtEjNDYzepmDy9hpS2Za3jJBjMYMVUh56Piv96zt02Vv0h+PrglbZ
zPGPl2JszP5uibFFSdpO4A2OZSA0ock5VMEUtA6VQzw1IK28vQXeVVhVz4Fx
2AFQKi6BioI7JI+3h4uWoxKq5RsKDCYg+qu31CbNOjsVfeICbzb0Ec93tuv/
Gt0rYWRJnd8BdJ/xO3A4BauKzGzfpy3ED7kiUZIZQ8ngXJkblL7mYWSR6HwQ
nmeH0UkTiExggk8Jz9rvWmhEZa61diBgSLk9+Q+rcihNr2OVXUVoR+C8VTgW
OmqeRVt9m5BX7jucRc5GWIpoGTT+y/d86gnQtiD4scUZhW7c9+k4u81+0UId
xVsQD5/shVZxmL3MYOzwK2QyN0gR8fAq9MyRob0mNuVkCkGGmh8/EXS4kc2L
tXpEjBt8kxUNC/JWn70XUfVI9j3Dy2jYRVcf8w8UO09seWkAVnkxW1jUwpeK
DoZf3cXsbZbJLhTytIIzfD48rlpIkqm94y/UucyuqhCLgYnOhdOWqOzO8bLm
z7A6Z5HbwfpNvhMxt9HTDG4q62Xzu+QEO72Sk34L237h1qvrx0aewgs0QCpM
m/rvD7UtpSF/kW+ZXVaz+hQtRjQJxkaa2AKuoS39ppuxbJ5xvpG3BI4KV6Ez
RXUcC/LHtyM5wZLBjXXFF8AfVNEpfNobOtMmWCN4xzGZpd4WVp1qKe+FwqhU
9miWpGX/0xsQ+jeJYk+Z7jljg6MeOUH35hgBt+hyRNNyoZ7vEUETS5HxHjHj
a48+Vs9OMAQGYu0l/FfCQoUHMkNDrcN+kS11X6i99VweWZtz4uiSs208Pen4
g4pDnvnpRmh/FG0FNNiBlA8IFRBUep6d0XW+LhCwZA6BtCrdOM8YiWPI3uEM
URP5a+ye/TNdG5ukBNX2httCqKN5fmVx32rOLtKnbMbsFKrOfYIaIcT/EQZ3
2tARD4O7mHE/iTDlpZKUQLV0/9uVq+6BQlBoPDqoE4v/WHGhxy/A4Q3jo4Y0
DkS87u/hEohL5VwGgehb4KJqwEd4vivH7SnUc4jOA6HBl1x7lxiIx2OQi1gL
H6ff2Adin27WqP0/j3jkpQZkYU8GxBKOJXlELEJuWWLFU/xgcu6qsUiA7/A6
/dy2qREJ7hZTCcOX/onoBvcQA9c/CWPJN3tVVGqWnCMKuhAnqv5Ra2/oTqQM
ZRYaK3armew1RxOvBFcDPNmXaLvcnq8H4DnO71mNPeHBkBGz69i4lzZty05t
aW7wWGhjU+SnbWM4Vngg/zZx88aAv3vnjyn4BNrLQ1wqNebniBZEtaBpZien
ZDd9n3qPFYk59m63FEUMbi+vUJQHIWD/QsesXb8QDVxFQEILr6lsoGnRn+GB
xjJI9o2K5ix7VmDLKvdrEwlvxCqMS1XdSr23dPncuJHsq3fRCuzeSr8hYkF6
KaIl6l0KuwZQMCD6vgIE4X3dEjDYnl2FDLjVxqesLyJVydJgOPId5zXD+y1t
QiwujomtVhjvWxXKSxy1jL2oiWDIlJpK3/vi7WkQW91tIm+ktbqQqUhHCcTu
9YnaMNdxSvvmqxQ0Ajz/Bcp491H9S2h0kuAo9PhonAeiqzzH58ICASZmwohV
bBGEUc4FSExCQiyMS3YMDyU0Y5slRjjqIYpdFh1jk9roKMInmeg04GZ6xs1p
YuJxH9TW6fmy1ngUFaAh1SoZy46flP4sm/+VAlKhFXGQTCfLRujColRbr/Yc
4iXagSfmFhDV8zDmIcwRXnhOPPZ+CYQTGKyoiZB6gpSATRI9hBofvxf2ygvK
OvVfwY7i+G/Dus16wfDoNBP+Oex1CbR92Jo2ImCDn31TRLqteS3oJOoUhslj
0Kn9Nid9BisRr3oQ0WUw02deu9IrppME8YrvkoJkBby/mYudKRMKQWeF8kmE
fKwMUcy0qzC7QDcqS3w/A0Yr/8t/05MctJBnyYLinnpkvkdzxbTozr48CQ3r
MlGNrD1Q7qqaLhPkMYVjQ8XS3mSwIr08lBul+Ss3NxiTR2mcqBscKeIP/2YX
XbqfuE4EcQMSXyj6J8npvhp/ILbc5C9sHvjW/1/iAzncb09ePwrc4FwEAKob
gWMKbuyiJpBPkherCYHmC6L7fOo+q2sJ/qfnG6Thd9wRNjTNrNWcCCDoyyR7
VaoEpBsB7sXq7cpdMRbjyjIsf8XYqoFSC0URpvXbKVBmJv101024pwuhaAn/
7szrNZAzm1mh+oQ7OxGGAClAEvFcvPVfng1mVp8KlKpsKoC3BBZLC7RxZ7Bf
WEdyyo+Why0rWXbNEjGWQx+99dTjTHhTGXrQoy7S1Uel53qtw9TNGbhlRVBA
gmJNiSJX8ww09qkzRUwRCVec+WWtHCKj+jwdya9T0e16LMa657DXhTwRZxVL
vdUWZavPKZPN2xVf2uPK3OkQhev227nTp3dZ9w0azujZmhmrXjdIKYYMFXR/
NOvrJx0xdo8754Ac3qS+mtyiplrdZQU5pUl3ub3+Dfjy1HKD/9QRolamOJEt
XFFWZ3as7SdGvyb7mclztJpX3NdU67cL5IoNVfenMdBfKbTJeVMKHPAR4u8O
/l+paYMf45e7ZpSTGIMQm6HCNnj6cZrtel6hkkHLze5u9/fhHq57enrH2O+6
tYXRR6YBqpMYXSL3ZPHaOLLDJCOZXSqhlWrze86dZxZc1WUeKsc7onTCLe71
tL8rB7bUJj9wCeCjCdooIrR48iH0HlB+LJkVqSYSzyRuNQG5GkAQ6iRGn7Pj
GrhJ8COfOQgsHqvVDmyBMxe/OOh1ZykzB/A/Fv5YXczwHWsCLtpUzS+4NhCC
ywZOr0X0gfbsvU9stnEb31uSgA5AuYfkGzHBff2xR5FCEpPhLCegIZvDVdP7
qwwZG2+yVeN/7nDCREpjvNy+P9o2rgb3G8CfFDyte2lnhHlF2E9DutD95mu5
oMb/y2mMCWFkHVAkr3WndpdOLD/lF98QXi+fFJiWwQNJ1wmPAnhu+ZZEkeYy
iYSLN6q3CaGRIoOoAJEkGB81H/bFSfc0VkPaG1R0pT6n8KCF+pS9TWFhRnNO
5NSRl6RU9tso5sftWC7mK1M8kYnB1eNL9qlFGsXIJ5fUoZkFk599ZFJiNYpP
IL0E7fU6v96Oc//io3GEp0Dpt3x79HQJR1KYH70bFueGbzXfgDeelxrJ952E
ZGrnDgiWVhBde8+h1w44xlc3j3IENl3drKIJ2Zeyd0/wIcxxi1Nwg9pzUV54
ZbapsV+CWw52GRPUWjKT19EXlcbeV7VdG/jSwbXiGvvQbxYheuzBQxTCQZPR
m9tlzcd6by9wIGUg8yM7GsrfG56vkDjRucFofqJYwdBqGpUghRjQ/nvGk8li
FIeCwosRs6ovv7vSToax1S9wYtn3KH1iMqIJ2CgtPyAMrY/Kagp8iSP8Uo0y
vVVNtji2Di6F1+3tMGXjqwCAn7refYyfe9mG01Tlg6udvXE5EM/SPTbKFojM
iJbujcsPKWXKOShhcenAtRoXUm6Hg49PjJ7A0u88cqpCE28NJjtaW7/MnW4b
teZFF94TAdfBTxawGwYlyspJxs04D3VRPw04LPErquy42Dx/4Vp+dJNsfGLK
NYXHDRAgz1kXuo0TgYbfICmMQ2K9a2I8fszTD3l1edlp63C3ifELrr+aMJZm
unIyYx88aPDbYgeTsv3OKo6QP2uooutfXyqM9GAvjpKR3AqOKw5bv+7/vTY6
usTUDt/e2UMwA84BhTNE2cBdhPba2P1IjHmHblwjxngFHYxaNdujBJ7e6Hkn
5/rt//gRHUROiVGFK1Nryg85Toj6L7Uz29F03j85KXpTo9yemRgtJBZXaI7o
mwcurFAXJIQn9GrwsyFpES6I36Poi/bUcORu7rO1rr60YtIUYYWXdy8WTIzn
cdESFQWWsihV4hagmYTsprK9XEYi+WkoS98+PflJA6xEAiPLDQ+swFrPve1O
/OwTtzAm7RBtkmlKwXfrdHL+evABIR8zBEmJPtClvYieOHaK5j147ebzPUbL
C7Q/b62/l9uQgzfyQaRuqJTF175tgY3r9oEvLrPlifYMOJ/r6gieZBQwB58b
tKkO0JfN57BLxEzJZFjFt/QUiS1EkZDPdZXoxVMKNWYg/n4iEkgjDTswTxzR
hd+RhrLdH7Y1pd1TPa4v79EFqB+jbacG8+C20x8kE9LkDGWKzr12MaS9Ypmq
Ff/4osMJQX9VrbPycsSiFY0MFfsmBNVP9mFK9VgUDly26lWWsFAN3x9khZtb
iraFbAgzwf+FDah0QKgBdq/pn7HUR/WyBV7/5DBpgvcu2XQujYSfrPhn1ONB
vQv92Aj8JKcSmBo27IBmXq1lAh1XSrriAiGfxlJ9HNPstJjDOnxrfmNkoVgq
EM/9AqaXjY/My95XH2GsY7aQLtm12KwbTvYFqP1Z8xJrZwAHgRjxpJNPVSLm
VcwcvmlE7ofCiRDOmS5jj2rxCF9jiw7MFEs94vyKHakbpXXeBorLNhrft266
BkmkzCE09FukFZgAJV6U01lsi2Ke6oZfZu0fY9PKQUav8aZ9OOl8BJ19GKrr
Gcf//3mEHcSOJ6Z7SAnXM41p32Jfjy6XRqP+6pNu/bPUA06K04bTDxpfznAW
jmGZ5tN74R7ZdQ6lgeH/CkCRJ5MObnURnFxaAHpRaGZ9CAMTshZObjMjrqnG
WH2ZyOJA9Qv1TQKE/v8jY+NN7Smd0PB9F+VWygbyt/Khgu9yZbkvfGjiXjA8
XH450x6trBs7LpAx+Nlak8qK7hh/qRaSVnLIeMf1N/VEOCT6GJnQkjO0spF2
xt9Y44sQFBR0gyO/H7hwnF/S8fhhqgt6O/SV93711CZPQ/gmK4SlSHpt0qRG
VUTsKCGASOykWNx+PtzAv4g/3OmoEmUkQURaiXyKRFfA9CnePmIrXE/OV5aF
oZlNz51fxyXbddiMTtVM7LPu0EjQZTyc0NfkJVJ7LeLLiHY5vL/7YI72OBMR
tPT3YPUuvH+gdTj1ddmGY/Bqh5xYKzhL5DgemvuTcpW3ep9cqpXA3Nsbk8kB
mU36C0A9I3iut0MhrTnKPiy1Yrc5Sp8M2LU64PKtvrj+mr6fFRrkI9tvHUd5
JdvHzstPV6FMLL9BQuVNz+usb+8ov31wcD4+HvHiqdYbtdK8B/9fw3L2A7Pi
dP5OGuLhaeZJdxhEOrfQ4g0R9OMPAXjwUPQpmUqmDOM9sC/lf/p/1JWB/Exa
4DgWg8fp28XQ/HszdRVbAm7DWRO4oTKwCeCEzVzxwLTDfpL5SwSA5KDSlpqT
QxNkdkmbBvV2ZU5T6r9+2TxudEhWBq4f+VHCCNWCTd+06TV6T5ATSSHMIQgf
OG9MboogFLzMLjLmwMVhKZ0fI4hOfeXf97DF5OEu9OzB6KcXIFFQkGe1P0fk
uPWQWyOTNdU+f/MfLVcU3V3yme7jT5HFJJpBM43n0pLtMWRZO7Hts+KGd0t3
uMDbaEH2tScKEHpZtItqLEyeTN6y5n4E55Gu1wt/V/ABVGu5F1Sg5KgVztuY
oiuI9dUX//33qVli6XnRvoJzap83O4dZdk/kWXzGgGUwnceXmKdZviYhlFxu
7e5pxo15nFje2TjeV0eBu8+oS9URCPfmRo9XDKhH4Ym8h8aVpcbJBSXsFs4L
0zRCuhSaSJ8YxwkZ10hQWIx3gu6DBR0pJg136irDLNy8HrQQZbm+4gzh0/MU
qNjQUJ4QDkwUG/RYfoXRpM9YuqZhHerBRpSALuXpcefhi3ic3eJzeN6updI1
ALxaeZniCPE/ASc1oFiXkZYqRo4uGb86NcLDLTUEQeQYXr/NZWBGl6+3jH7G
eqyEfTPims1Q9gK6j5uNJXknni82CpkguyX3O2mHZLSVXsevi4MvPDLBs4Bs
QVcRaIWlZOHwwTd9S2cFHCFOrOC85TkH40UuOpk55WLJ8m5P1czfk+kKjWy7
8fY0jHz9OIOtDwxyvv0lcRYSZn5OowXmyHEA8i9HiARNxwtI2KxXHWVP/c3r
XN1p55quHL6WhpAnt4XLxVt4GXFdgVV8NqaITZDwwXC/ZdsZcBK8HOhSUPyh
Ebkiqfc0yHHXs93EjqtlXHyg/CGFEiha6oevMeTlxRk/4jueDz+6iLeZoLz1
UkMun2sGNcF3y4ztDdFkwBE3i/A34gOoloDHaCOQ9uL95ks3XtXnYrYs+w3y
8r85i6Cs7i4YJ8JYxqhucwj+Q2EeWPtU3eeaCHk3Ai+R+W7N9a//j/NsRI9i
0KTcmXm0MpkKRUUiblIQge6qg5X4VB4VLyRPYK6oIpoeLJmPrtjZmMCzAscZ
1T8PpdURAy4F+XAMwCVIS8uyRZRjle7+9y0Wjgaq3H1XeiTQxKiBdK2VMSZ9
IFNZrEttvyGrc4HYkttqMszhwRp8xp86OsKo6vlGCi/WLKosmpOxUoaie2i9
DndS4BJeyHMM1bIDV64mcxFKLr1n39eTG1PsywcLF2dgctS+0BdGWsUA52X/
ziZbyb5aT7ChY9SNeSWF6DMqlszio9G3N05Bq2LaM6n68VUsU6dZuYW1IHb8
g2ZWWL3UFyqw8bTwXcpvebvmtCnjW+QWDs4wvSMGmHqRAcUabXGN+OrCqezV
h01aMc8g+NwJ3/lB4W3L8S7DpT4dJxqZh+HJtbSZ1wW3auby3CTdeDmqpg3Y
/PcYXAhrLCSFUkbleH9jLbtvIBe5U3PQqTtiKiZ8TUhcQ5cbyisq0/RkzcSq
ywZzTmZC5CMj0IdRC9+GN1nwZ3Bwi6jgNexrZBm9dumvuGCic7MW6abpQSwL
YwVojXUtgzfniI0Awhu9Qsc1Vd6XZqNlZ+7JBTPCMBZR0E/lK/fqtfwFUPqW
uE6OyfX4Au2gxnYI/cro16QhYoednDRfDBJn3bW/zl5xy4xkGAgp8SJGA6RN
HugXTCLbW+dLhJ/IR/TGJEeihSTnn/EXL22MpopTVIW25fxgN4ugM3BuPcZX
+VgE/0seT5497fRe2h4utQYbE6kvxKP5FgZGDSLmWkerS1RXeHdtn8NIOZuh
9gN+GpERgdiSownETez7wOMGvncN1dnyXZK8Sjm/uaxuRTdRA8MUELOxZGbj
p9Za04aIWf7WZ3VeI16JnhQS0KxUTMEnrYhF54h1BdWbjrM9G1mBFiQWHK+C
8Z6eNSYV2kJK3OfmhpWk321Rp9TDV+q2nYfEevtnbwvh2DFrrWp+2FFccK66
pQbSqgfJ7Hwrr52vLPqjGVQN/oyJ9S4abSoXGiubiu9acB7qQBYhwGkFYJFK
2yocksKf78SLBicwzXaTTSJxw+eEOsOnB/IrZCpV2wshhr+y0D6/8iNnd5hg
S6fB/28ncUB6/WjbZoWecfuJ8FfMqaLed1Fgp0TMHnMJS97p6CdVyWVRCQsQ
a+09ZDzFzgFHn2Yz3DM0Nax2SLodtyF8ZEtdm2WfTVA0SXw8iGU1zG51a3ni
JFJJ6fCbD6hRrEneQ8VozVwYdIwfa8zbxWDQ2i26Z3ohZDyriB6ydkSu8S9c
x2Zp4p/OeS4zXO37CgEwyR1zfEUirtcnei3Jf2Y1O66oTfkoNg70rRWPPDwY
3bgsNu6D/j31YbTPC00HJxgXNBJ52VGcpQdKy3K9By0c4Nxb9iUQaGzj8uPF
MuocY9+mBt/jh4h7EV7PWf9WXJr0RkrXMRGmjVvDTf6yXRozf/Wg6zLsjhnL
xQpR6s51MV6WihX41h1iRSp9ftD4sbORdu0MWQgcV5ao9xU0PYQTb9QEEmTJ
73XGGQMKWFxXKpjAPF5c9dSetHZKUTjsFDHXTuT3ol9A8Jf6+U/vnj7rGg26
DnhfKmorrubdyHzkzVy8OhJrmIkH4zwiKweQp+IvpnIRI3t31haPUhK/wyZ3
FlS2WPnzrUBYC9Fn774FBR0y3Rgc4tpbckCwKbb3jFsxxnvpuMMAx4w1bJQ5
aVbCrTDhYH8gU7bGtUN2XYlBVcJhiCCTqNy5O9XJS2tJcoJnvuH0+9RgAKZt
6izta2+Kd053J+p6W81JAmZceMT5UHfShwow5fJ06YcpBx2mOJjQK3WEqW3P
qxIDRmkGE2+aEVmEEkAKzq61lr+GHfu8UAQ+LT00AwXVgwhClHj9BXCatUYK
adkTWkDe0TiDZC3Aucpc4pmURy9kDb435mMzSG3qm2XIXaa99DB4d7FtmaRd
6ieGU0k7w6ePNIHFK6exhzjyjU2r8GYDrk0VymXJ+y12JVJs35VMedkshdzq
MnAwYlRNIAWEr5MYl64PLBKlr6YUVAZdGycZ4bHeJltVxVylHtcx+HuGWnb4
7mYIyCYGRFpsYdN0i0lviARwU5a+ncD0PEXrPGnGULwFbo9NKTPcrbms9tQj
06IOzYSe/2B50dwmgVKZ3VUfYKRLdiUUIG6OWcoiLkUjAOcby3d4acTcYKTm
5s+DWs3aK+5/skm0pkl+gAH0e3dNp9Y4djKnaBYc6Zbmwth/ygH9KDAqcXDl
9o/Wn7d57LB3o2i9jJMrBvEeAC+1mJxVMajRkZZfYGgMWrz7VbfNXZB+3XRs
sui9PLSMnCt7ZBaeN64HGdJ3vBY+gzpk2A/lxPbsO1oLVb/uT0ieUqS7dV3W
NsoPCkZDsBVPxrmwNWZOV+CxONDm8b+x2Ir9lfcfUWtO97QmuN3iYC+cGzE/
07YlTRYxpAy88siUtr3eCScqj6XQL+GfZHzQkP1t2ucvGSdUvwonwxByvcAg
ThqrxN2FNHuw5jdzHuYwp8OeClB7DgS58Io6xJdI43w9j+b2zP/GgviZjbv/
WvfEf+6FaHcBSECE5WYfmDeInpgO7rCAWtXNJ7AvSScewps3q19Cf9lKptMV
dWE5Z4ePyKthHESgCOum4SzmJJKq9w7wST9pkyIQg5PntOBKvxNwJnlrVMgz
fq90CH5xq6hMoeqR8ifosJZi6/eVubhY+QbLkA2yaWrHzI0rhWItV27v4+X9
Ps6qbtWlt+mrY7Tb4S8Au4fingBSe2XSwhMHyrbOgtQMFnamhCv2j7ioC6va
J5N5PypD0jh19xOBOzIsKJMlRBz/Y9AitbbYoTJjuSCDDkzl/6M+azJEfhtb
ad6r22B8A51Q9pgB+SxJgv4WqxQ3O7VMnZGe/LkPdkQ4dankv8Ul2iytNgp7
ZDOCSPiCo/EynVKrdE97+jbigVFntHMMNiLmTELt7K0ePvP6TmIjpq3W7QkP
ypyOIxfARlC2Faf7EdIOx/Y2V6k36+1xormCoXvhYynvjWzbaer+6teSVG7Y
VkNqXmgErYNEvJ008q4Zdt9w78sPYtQrSv7mEgPZZNZOCwEdiiR4P/PPxmJA
ZXRZrSxB93OEJFsR9L9GLVSf3V8NysYKJxgtMeZIvG07IP73+jfTg2bd77Az
wmP27NayIVJag7feqvZGexa2J7v0vBDsc5fqzJujhMptjRys2uqS6gtfCPoE
osPfmVqWMoGQ9lKlgP53zuLoQ8ZDNoK/YKaRmCS9wtVXES5FZo75tbHALmeC
AZMSExTek+JM1XXJcD0aIiHiKhuzr2TfEo3aPLChxTykBLcl3i9Kgngdr8PS
Xigc72wn2FkbozsM7f2ZLCdVOeRBhJB3U5M9kXaRzAjPAt8GE+4WJ8Fjtqs0
/iR1ULezjdimwmbzykhgaCo+u6q1Ew0vzqaYCwLzI9pmt70Z9EtY8JDuMCTP
KnuWP2+znu7PJGnhE1ud+1dQqMMjRWvO2WEpngkrk5EOSEMxA+dyB0kvMHRN
j/ag1eS7srzBlSJNYWUPZLDIO3gbURk2PptiNzOpncsrRa8Tg2qIPmPXpEjY
H3SKEvRJzcIEB56UU11fM3XRN/Nh49kQfTum3E4T0hTFobct6d5KpzrB/sWN
yEIih69Qyv0uNFNaMlHwLiod5hIUzgI5FJINoRpslIwvrAbbP3uvzAPDeuzu
iGBF1hA7snhy/1+YNIs8gMA6FsCkCmIGvv3gXesMW10VWJd1R8e9Fd5DCZ8R
v43llP802K7TGWJMFmoyZcs4u70GRz0i9gWDTXUtnHr5iVTfBTLLtbjrQ2HK
fOk6Lw4ot8SI+CSkrpI2DchZKbQL0nsxJwyeWJ205j4LfYQwts7o490LXv/x
B4sfJ/tBB/Y0Yj9RCwyg3tRSBhNT14fHUo7BiYqQRktfm0kjAo5qxhn5cRqv
44XwXvyY3wLh8KH+jPAgsmfCuLHcZtHveDWCwta6lgpD9n0eVpPaHgzpjskS
k6MleRVjkN7M1QS2CxL0mm5TKMWiyt+CbwCXDV6Um4PJfzvBwyr+InmsZ6Z5
B6+rksh7xKc48a5XOH3HSvjrC+7o+4grIHmAhe1CtOVCdWrAQPQ4bzflUU95
bKBVqFoLKG1FguFUvJgeh6+H7BkEDVCrcL0Cuio5ED3yqBjZLgTbRBrudyEm
E83gcWzaDi5VVwMGWh/nxyF3jrGtUN7n1pjFxw/E+8BpKpXMMYdN1YzO7y6y
Uta3/bnMS7JFulkCBpDtzK2vkDGLKxRfIQpWtR1mqp9gOp6OvQzXzT9M/ouU
ixpAqWy8W0ImizUxV2y/lIsh5cv+2IcUdaNCW6087VXlXcDYLRWKrHbT/f26
6Lnwh7EdMDH2AVx8ayZYh4gy5v9hZqSs41mxRd3WA/zvFPwrTKXvKA3nE21q
xzj1L1r6kcgQ5RqkAvFQjBHIyQ9ttinAQCzui6ApZowjk0Nw1o3PW7OmEW4q
kGHdVAV+8iXtzGD9gnjSeKnuD2RHOmF9JTNgea6SHnyDEOkYcnrdK1crUDDj
+cbFDJ0/APdCoktOdzPmT7yYRO1SL0i1XTyKjHUgUi3DZJH080F0gmMKRBZG
TZnNW2vwWqvzlSTY5XXNKqKIr0ZAv1xQq34m99caS3soei0f/d6VrCKsvpjV
+eS9qu+nNjWqtq+PwayfO4MyosKG+uJoy86/vMUh4oDOLL1D/SKrfmstiLAP
mZjntMSStbXFqLAYiCY+cKRgSc4rbU3gOW+xhBGw14dmGgTW18wQFe+A/+9+
UDviAqSMOWPgS6RlL8Y2GxSpulNgCu0zuobeG/rjDJ3RerPcooDfbEB2Dcro
ODEL45jopXXjoV93BT/I0j73vNOCtJFsfOTX0KmPAbz798UzRmPyeDf4Zdrz
yMHuLMcEazI1qDbCgzipQCrYyLHr6c2Yvl65bpvm+TgZ4rksUQQMMM0/puaD
Zv9YvHGM3upJUODg4Ow5TGahgoaRpm+gpugydfCI99v9ZorqkMg+Fvr1LTmK
yY6pAcS+Ai4CcaNo+PeL+Y9sqwiZWWJWBrrDk+2XzkSlEHRBktj/7SPIesav
/tfGoqy5oEWfmNe74e37z3/ZniRGqnkjFFWL9czAWBEqiMX5vZvf/JdMtGQz
fTut4F7hD8cQUhBaZB81G9sUfCfj1J82LUX/YHCwHhG4kXSlIj/0GrgAn7/D
VZLj5JvBm/gGzmEuoMFurCp+mbeQ3ogHA/ycJ6QYjQzEdcilxsVIKeXSLphT
99zyndC92sxuBRaJRAQnkY+pvkqqZ57OMBgUyxfOkSLQv/fXiSgyhNM91uUr
k34MmjRPTgMeIwq6rsOQGQ6Pmt/b2+nrsUStI55Qcy/1Olw+2+fxW4SwzLxp
thKjNN/dcif2+Rsz6mLNzW2F5fng32DwFY98ewwoNmSWaxR4Hh6GatawHJxc
wB8nwLchyllwPUY4Ee983AxPHJtznKfVuQS0y2d1kWdGUBodxEeiqU5nVab1
Ybj5/5hNIY43noCxK4fObHDemNnv2dQc6Uj3uThFcuDjpeFw7032eftLq3Ua
CiY8ogs0MxHmUJCkfrPffSBsgTcOFM7ce+9odnnLP8u66dEteAx8F21rEyHQ
dxpnYFzk4q2vbYXKmHUih8UHAsOlyCZzZSFg6qNsf2AjIoxlMf6dh4Fa1EYb
NXwUcEpmNi8w05WQ61bXp5oz57V4KhT206JNFzYMK1n0ODKjKdDg7mdvTbRc
XijwLZ549ymsa/9DZHJgChkn/QPqB3a3YiTSR/1aLRArYFVl0QEBf+QTHhht
w9ArDDumHflrC9qp/ZO0dWqZ2Egt6ubbvoOyrZ7Bu/SXziK7KeBO8cahXexn
qybYh0WtxifbqGYWrf3Qn/h2OkM36AN/lgP1Pox5DHjldJBBQpzKY6YA5d2h
UX9i9A7X2rek4oKSikSA7dYvEhB2SH5YyOz29BZpkcH5Ug51ipbB2tC4UOkG
35jstxhlkXxpyla6ajsCFoP3H7L1Z6XROr7JEv+ab3ELBC36BSasoAsx+1up
P4DjJI2ry6255X/A17mCgpUlcTT3gG9T8V3kh5X1Wmne3ffpr7iaggklWCZf
orJ64dCwkMw6Rx3ipK/1yE1yM9BBQAO+ApbhNeM/henkrLPTHBFv52lqZlZ5
/VVR7Q3F40cRsuZb2ilDkG1UuMDwFBVNrv6huHSiNnPhy3iobncZgn2C0EBJ
k3JdwDOekEo796Tv8JBGoFw3+NvCcgisAiI27smFwm8rTKxojux9EA/a58aa
K20NiQdYtovtrYG4705XVYEqtStZP9LcwE0BtwYGyUwezJK8njxiziCml0Nu
01Mtnym4yL4NX7i3CxPperTxPlpprYSvUu5k920f+o6xU7yRt4PRxggtjnPz
+VFv+4pA/8ZPatm8iMxjHbyqpFxmuACKDgMrhkwTCK/+rBkg5wH5CgrwePh+
vQc+h5kDWyKWnp6N1WBrFdhAgb4of0lhz8bzitmyK/vIiM586qG4Q9vBYNTm
gVEx/kqWbd5oKmyqpY6Fxfe8xvaXssVHhQGju+iDKWuCXweqGo9m+Xbwjh8j
SRaN0PbIA+7Ewjw/MeIo54Q2Osbf9dXx19iqO+qP4tmr+MpqAHC5vMxr8IuP
HlK1fqxxQwlUc3M9qks1xMPT0KNZeoWTLzLSVskmuHcx6GXiErM8tTmKImmd
tHlZ0tOJNbm84jb7//Uo6uG5pYBxTHNydHqrYperdS29IBy+gQj58U3zKzGt
qCKcviKMT1Bo5zImJxdp1PbILdwMj/3tkhMogL7AJramrmQaCXl0oaCvFcHv
zfKgjZOv/vCM2dBGzRWVNIlW/9gXML5jSudvhjaEV+yuWCxXbc3rF19Fwbza
fnnKD3VR7l3ZUx2/hum4A6M8ouLnWdytAVZMGu78cdX0jd9oVUj8y9P/YBLc
NnLH66z1sk4zaG6frWXzmka9Y8VS4771QJd2rFlxi6ilCUd2eDkGX/1V6V+g
y3c+zGfcQxLcuxXXsyWqIngEEnzeqdHuiRdfN2k7SRJeULoPTBI0yleUB5GG
EtCoqmG/BHi4cUrhwOCOIGLDI/xFdPQXjMjLA4sO3wGlw7hr/pONeVwlTyhm
SmKnWboDB3GVO3/SkqmjGdJHwuMvx2UQz9oh4waGGJu+T6lXEhP7vr0yehpZ
ANw8v3fY/XnsEo/4Q+nyaNmOHNwp+mmv4AJoqwnef3/4XM4WZphMACEUU9QY
ujTSpg8nZjr2PoHyxSmKW5QEViF+a7BzcwL+OdL9CtT1j8aBV3NkDiJtshjE
ZxWrtoBMlXaY4ILulm1hZARTgfTNr1t93eTDpAb1vR3NkFLLK6XsyYoQ+D0i
NpldffNb84wF4QM7jFp4NpLSIROksCtODnzJB+HNSF+R8FtiWDXmui2kO9gU
e3Ly90FHbOuC+FsUn6vCKQgeSKiP26I+/2vrGxLktqElew4Ljy4DFUJxrXDJ
WJYAvM+IAAphVualy8/FuaMadPAoLEw8HRMX5lJ4WB+yjPvKpjFqUxVxVNur
3+xOBKoPlN1QWrUjJ+K/JC1FqLs6nhihYAHuro5iPvbgZaPqTRqGBink5kUA
5Mg4mhvDmzjYPQVZk9DFXN14F1sc4njlWQj6VYR3JJ6m7sy3GiJA+nI8Qidt
5lbFoVDF1+/3edHlHxvMpdg/Gv0suWrUpEnsAtoZsL68uTDQhINC7P7qdK/D
cdVin/jSk+RGc1/+msh3S6mPJp46GSapvmLgokgmvDKjoTk+H5Zzdp6r2iUn
1UOSp1DcPfcfOkhgoRrzgu0JMpUky7RtTmwF1TODIUYD5AuU3Ajlh7yk64UU
LKy8AloiUYXMGItuMnfFswVaOEkB2n31jVUvq7aNN3+x311EL9C//VYxjWRG
ygmA1APEVSHFq97HRzjKLNaT+F0eUiee/GLsRvYuIkqdI8Vy7Y1L92nDaIwf
B1/3npLqtOn6CmCmHlSmxLXw2yX7a2mtTf9f1VvYBYK8LXpryn80GXGlfdWF
jtLFbXUnVkJJgAHD6iEOn9+WbNcHb9Ea16n3iM3DqS9AJ/i4TcmGOikE5QJH
NyhESVjUfPjfocyrHz2S6qJLBtB3+U0sVThyQtiYddRzCZH0ZbufgnWkw/zm
dnPhfIByuxE9PEl1BnfovCsVcMJHOQMIesf2i9mjz7TmdXNykPLnNKN/dJxq
Zqs3Z/V/Nq2PUPtnUBbgAFIT1HO10PKeLNuje8SzfcPF7DBNw23CgcVI+rtu
wBfD6uMinMrhhCEKKQSG5PwY9gr5HmONsKkV2rpmQXl9UDcCV39UD4dOZRxh
rj+qEqCTMy0elG26Ko5WSnJ1A9o0JWF/TgvfHGs4vnpWNFyBdkfyKwJQepA4
mNwS5Sq9exuSIYn1ocftjhd/NQhE4k6RCRvTzPQD3jBBuHYpdaoPgoIdCcOm
uydWgVgIUAnRLF/FqBrwKKYmY3nHanXlbpeCPNX+4fewcGW6n7an5T86F0Mt
yJHOoigp8+bqUMKjw1bkL9Q0yGi2c3E7ud+REVjHVK4j1k5i8P5ermYBKZcg
noua+Hdk02TKEjf1o9fQS+MAg69Bvv8nQiTUtz/NmKHp4bHay38lV++3/3AF
jXTRj5JvjC9BMInLISPW5Dk59OQkGQnzno/h5Ea03eWJqHh6q1l17SyT+omi
v043n3UUuCWU7KQUVEeFu3T0jSjtbPg9B4kbCuDOXje0lBMBDv+r9E7ks0xR
JCaXXJP/7/v5KrSI7qN3wjsWMUU74Tu6yX4uYxbmMTd2fde9F2Vjl84WQwcz
JZAvxIu+dZsQxU1ObeC6FD7YdKwZoVnhx6x8/gyLZjImN2Mv0NnAvKfj9TFv
rUT/SbHpyDVhz+OYI/bjtoe2VG/+i/G4pep0LSIyjSYiKEO/Uyji/IbXdUtZ
zYFur4tzKeHQR30azmZ8fTDrKqc81ZJnTQwp6ltyAm13axx0CE3U/Vfelqq3
4Cy2AQOUgvSHnRiOpZBa/N75bsANqa5EUWIa8oXQueDPaGXENw7KWS4ou0t9
MyAl9NTW0mHW1h4vn38qx/hl/j9lXpWE33mIIfAt6yu/8JxTD5kTyBExhkQz
H7g90BBdKhzikBtlekmglbsuH0iGmM82qJIfLurgmlCRAtHB5VDtUhge6qf0
qjCV/xgWfVXpEhBRTEQ8507aQuo/oozG27cm4vsw7tf+hbU8tGJBF3ICOqzJ
3lUtSwjOXj0SncYksjMRKM0iLHxnOvOMX3T3Qa1Pao3pn/U6PAjn+0K8h+44
HLrynOOBihkTLKGqSvcaNOb3qPK8H3I609uDXjwtORYcvhHX0us6yCIJxH9O
vFxj7zieJ2w7TqLybL46Y6txIEVmy93Khalq4y30JvEUdbRcxK4pR/I7OViI
E9CzkGi0sE5YOv4GK170Idr2d2quEwpsAP4col3vKYKnRUrutjDffEjeKr4H
0aH5EOR1pI8c+9X46nBK3Ix2pClLUH4ik0hsqtFFP08uaWbQN/TqzTIuMaJn
NX42VWhSQVvx1vG95u2lbipg+pvc+ZTNf9qb5YUjB1PMm8AIQanNmFhN1DV8
isliqw9HjzUwVeMiHv1oFNRQNnLgqV3CipiHhPPKxZd2+aR+qyeiXwwx2S4N
MllwvGEyqBu1jThsHpYoc5flIoVFw4mqVZgMDOWLhUbpbUj9lwcwKIDKfSde
6/O2cuQWAAbVudOojLiGkCNe+JU5XU7on4BVUEDrp67fZGSDqq05fShDcDPR
coIGeisqz+tioETi7NfcdkbdmqNi6qMBl2YG+mRhNAwjGJSP01nJyQEJKCGv
nVsdZEcuqt3fveD2UiPmNX/mLgS5K5nqmsuTxE5bTyY5o+0A7MNbt6E0Ns6p
KMCsHA9+7GyTSUNaUQz8MHcqk6bIDDWvvmPT7O7jz8vKxgZkW2gm/e7GW7Pk
ZFYLS+0aH7kCgzY8gj2jxblpLh62EGOLlMYXsUEW8rzOxHJfiR2yj76RwwgW
TsIdt1Pjtb0eDFHGkDfPiQhEVfGtPXm8CnteyyLNi54pPDy2zT8eAkAWOxIz
7n27S35kznUOrhg7fcMKx9YGl9mal2N5+NObTvfvp6cg/2lBBKcYybfFCbBZ
LN07+SgHlgL+iHlFTAHEYGC9vopuCMlp61hiKOTyPr+bnyDeGU2/G7IjB0pG
Z+pP0ZBP6tVHNydGKpim6xU7uxqWL+9jID9/2L2zSsV8M1BK5SG+J0YrO/p8
g7EFrYjZ+H11skc1Nux7Fk9Xqlep5/lnk2FWRv5Aus0sfoV2/2mIVcXpWIk8
COzbUwPWpZC1h86qpCE5buirsUMYd9sV8geH7X9xPV32cjDKT8/5ApF2ssME
Jm40CPe0tRrFv5mnoB4dWgJxrGkQngtfDMLhDfSYNaBFnGU7xJw+1XWiwJmd
4Qjc7P0rM9H/15A3cZGiP/bzn96V5qbXXoxIyqjzIwEDw1ovHWAPBcX8frpL
Dh4eMqPO1BrPRKBtkprRyaWpYx8cBftVok/4orXHv6jyo9vZybhxq++j1wVF
A8+trkex1ldpU/cDAgBmlMttXjYGlnKv3SDuXnzRPZkMmB4g/ynSKmJTbtWY
g0/qPuH983hD/ueZ+6hLgcIo6XsLPEkhZ1EaQmDiFl45E+8zERkNlxk82RDE
xEcuFTWCsro5bIxoY2W+9nNOfmYtjzofGjOUvy1M+dn5Opl+hfqgH5HUHXwX
WOXQwOydEeXQ1ixG713QpJ9yJ2nI02IicF1ChFRZ2wjcVr0hyyLIoUsDqqET
WBniTiR+FW1VoxePL/cyNHNKJMSAS6QZn16MWWmKldJmdAFIy8xsrl6WgBNE
Eqgl10cjukfEgsVeDBwLsTpL4ZtWMN3iZY3ILunXPpFtvBCuM6kexy3+dWXz
kRA444YFqOfYeoXgfiC6zsy0qK0+QHVn3JoQzhBqQLEgY3u4YAyRf9lFvOv9
UpYsPV3D1Ot8jBfcZ2kF1mbyhrPrhpaKYqxsKUpTwrCE3rtC+mgm+qy8vH/G
82ZnoUoF/T2h7p8BertA0Y5CfsVnDs5Nz0cwQOJJJjUh3O1lj6jy/Widh3DS
9lT4BZo3lsI87/42K0sRhgVQqD+pF0226fUsXA68KDRPj9TOvIuu1u5uQy5R
sZAufGxSOXZv/HW+FVBvyW4SDAMvQAz4DkQABrNBFCbgzg9Gn2Ign48MrSBn
UqU+N/rDFcBSZrmQfY6OvY5W9KfsoYSw0O6YQZZA9cyUycmSE7aiLQENeM3y
GSe9C/y8o5IOe6CIUYdl7KxAfXRpo4Jo21TXYWB0n8LYqcbVbIBSLKqKTakU
IXvOa/Dx0uI4hUNABhigLMMSPZAxSB7ObjSnuuY8o9TBIvmSqSXF8210AckR
4rjXnUEKWsH993+gEdcKVF8IIypl3+oPP6e9SVuI4th/ND8FR+/8+FdIEsw1
nZ1t/meO9D4w7cA6XzqwmtCOoNmd00TWM124b6i0xF2KaZoMVMUKS7hVJmlf
041vBImzB/14q3DS4Dg55DAB3NugIUZe2nQxrPaw6fmYUZZm4A1GHutN+5Q6
GMISqGCsQBQT1DHNPbpHnsrXJBsclI0HnR4JWw811hZrFe11fiEDEJr/qZtv
wvGix+CVcFXL73MVFryyBU8wKODQIyuSGrJuYAzz44hgPBooR4f/f56DXlUT
jLF6wkw2KofBVXVRyrueqxfXa1PUnInNMlaPbTciZbJRJixmka2FqabP7tBL
mru2xE72TJIequ+E6VVHySg9CGXtG90Yd1txyyQ4PxwyFXwbRwcPWXnCnsWo
cCu2E0qjkT11odO7NkOIIibcZk9lzb2LK26voIMfzWM4IWrmMuiOt2sZcwTs
hyS0jOG11xb4K6D/XRgje9ZI0RPuS5t4BrAHVCfXOlvgi2ry5DA7w73l51xY
i1Qze/ENCmC83p7VoZs5v+toCdZt1pgrOI4zACQnK+ixQmj7ftlAOIBjF4VE
CluHHzLIg07yInopEalSPIEt2gt9cqICGb3TTCd9WDpLuZ9pMcQ6lznbTMKO
3t0egbFQXOSSRxlR3eZPVGxJ5srwT0zLYREIlE5eYs9lu30MF15hah0CgA/W
I/4S1lOJ+WuEklhUJINW9WOBy0FiqxtVKzDZN2avWdwEip1NWRx43TEV6h2i
SoGQiO3qKcvYLBuxHtXknWo/kuQUVNm60K5+KeNOZnaENcrlzlZECCEzBM8i
wGO3WvuVsIwB+LSCcWDzWqtL7R9AeH7JO3kLsqmzlh2+X2cgmTNHqVHNPIlr
T6KOEdqhiCB1ckPVhQBnUeopjGb8jM0e8YJn9XqjzBnD5cr7npWzYduCeLCm
+ey9pKLrr+4dFdRLf5RXJfHVClSPNexKhCpgTcj9XBayZbPYW89Yfzv+QqMS
/jEODPJ9JgloPXWmPeQ7nW0Q4MNx4zuZD5zpG/dFl5lZtoZgweJJEqlCSH9x
//aMBS3PYPb1Ldgl+FjxJgIdZeOWZeppHoADuOLtbYK2DuNC4/AlD4hSyfjJ
eKX0WjGX+VsC9Lvi+gWE5P/quGGFZloGSP/6bH0qh5hWT5NygDQPd3I2xfn7
29VIYnaKViDNRRS1hITQ6hCXb5VsllsTyuxf+eYC8Da9M9SHYWQf3WISWC0z
xPqQWntS5V/XA/HHG/L7NJCmg7QJgDb/JskLpRMVlxICgDrudjmYi7x5hGdD
9ho0cRUQkQLDmI1V4oIgfUNv9E+xujtYoE4Fi/CceDuM9ye/mR/OhQQDw8xE
5iUdszYMkOm+WxhYIoRgyozjBhc46h9iGK01L4isGKgnSPITb2y7E7eSWAO0
XzLoqr5xW5d0DyKrta7Xlaf/S1HpPMGHKfEcHfcDnnE9iuKkXjeaqKk/Sehd
RYMTai3k65nvbwYIiPZHk3H36ETBRE2SdDE55ayfc2QU3kL1OSXCOzrya3HL
G5sebgoq07BhqnKiLIU28XD7CPV2pkCztWTbtIynJi1PJwfBrG85TmGxVHyW
3wEVBE/mKPY0CT3qLnsceNemBYz+my7UwJ6iUqZYR35Dskt6FTnKYoBRl6wJ
o6RJsHbh5T0xCDPfLwltJcEc7NNMsEk7rjL0yS/Hby3W7INXjy5CYBt14Vex
I3RrJPuXWJLPEj5bnWkRDMyWhrVrOtN5GdkFS9tjxIsKGwoaIAmilrLNgNl4
wpLDQd3VhDRN5kZiwIb/wGHphH2QfFX4IcRvc0gpEobREF8QXI/b3wsPbLYM
rkluxVudu6fctlcyOoNOzB2wiWZxYKOC2rq47+8trhdLlxVHoyddWZHS51Ng
xEcVu7gmCt2D7G9w2qsGvn85O3XLu9YhO8E9OsvY7pAoHDF2ufTEloocRAMc
Pe35t6lWPtL07nzF5zc5Glotl69tCRhLTIXOBjp9LJTsCRhIoG8j+DSzyQ6U
nqtQ4hEHAIAQmQnJhdo+OqBD0Be0C4lkmwSltE1C7A9fA/yF1sYCrbktFLhl
2s+GKi/QmExfFOgOZmL8HapiZrhnSzZfmmiqmadalhlcQZtZL66zKMPEn1d8
v/VSK2FkO4/ehZ621Wvzb5ujuNIKL8CnyyOOsgtVlm8kps3tGTqvF2LWkp0o
a4/2A1jyEHACbMy5knYSfDPXK+luH7ZfExgIjuU2NYB4OhMG3jbyMzP0By93
yn2rcCyGNUEX0K87PoPI6dUspvWADHwt6iI168pxf0ox0vH2O4kxmaZvPDMr
zVGKk31OUlFHryHKZrLdzw23GHmyHAKZLR8eIFoHqjkE8fl8Tgr6zabxcOtT
3LHEThNbGkGxH1PF0MEpRk+TDq4fSfUva1qPngo536HQRv8SazrilSGCT1a/
N/YpH1PZZXTbeffqlezAht85bZmpr+24lL+AwfJT4RBgyHGB/XDQr+9S+/yx
TnmliD6GZYM0bRzOD5pcUyilamxA2/rZedeaikedv8zs8WW74yPdiTwGjYc2
URGLcynkfuAzZiiz5Nii0lo6b862gFJ6Z1ggjNh0v5KMIiVTgd7oN1eS6clY
XDYF0uoCAdyVzSkgjkVtRkrNnO9iJSRhL7o86oB5d4dhNe/ihiKNAj62AaUu
ewJWF6aOLrdbAj06NYfLoa4/7ZwCoIM2KAdAPswrcDzanENqyYov2WNxL8BF
+wPhsDpOWK8b15wfNvlopl2VT2ZGMuH9hrdJ3NdxXd9GC+8IvS11J3CEYIKD
leEmqyNygfOZyQIYmt/lsTMYBnUoXet/oT2O23nhRL+yfbtWOWmWEASl/FCb
jvEXpd1K137LgxcGyXTRokPnMtbe9OU7CI8EGyyRmN+BLB4Yrmv9GwkzR9us
EznYZGKVEiB/oIjeigUDxVzzyPgJ1LKjYdZOd9717gtzK3PZtsw5RrLF9VFj
GSplpWpiXmLSfFNAKKMr/lnTefFoVSyZmrIMknLv4+LEnfZP3Hz1MzHx12nP
Mak/DNcv9/dEXqrGnTlsUBu4cnTridWgHASdBoQnX+d+P1GVNNvRa1Q5nCGC
NOxKfvEjrX4xknmMAci2GH7wPBPItoU7NxRK6bimmGVV9HaSbjHpfPF8mAEO
k4tqKVk6WRV58u0z+IMsURdiApm1+ywZtxuVr/SMM/cuZxe7aZiNVQHPeM1I
ke/2PmegjvEF0A6vmnsEbxh07nKpZX/cOXME0YmOUoJY55TqJ7tfDBBcmkFI
YCaP2e3zVUk7IVlcn0xKZV653aDK5ECTOnxeu99V85ausQb7d0whUYwI4DVh
DC4Vh0A/rcRfqKvTQFVldqfyeOUG/H0/O4opKHdfz1do/RQbTHR1OUgWCZUX
wOy+WmEtxj6cjMxlcZyK3DmkS+H7yQFFECrKvDJ8Ef/7Dhl/9uYVcyrId7Yr
78nWy6mg7AhA/nG2HZu0V7V5NKASspnRw6Uwr9lQDJoP2Bys0XwfUBPWvHog
WepC2IY3tDKnT+uhDAldeQE/P3cycgQdsTVG+hKmQXhsTrRxlnLovxwdu/Lb
nHOy0laWpPei1vdQF9ayNuRjJqMgCfCMcE24OkrZ9+iMmTEyMgyugLr5+V/5
+tmOvGyUj3BUutvtYoT+kiPZ+xTc+v74O8Wz7L3VwvuPdlhhD0XaU+XPpthI
KQMMHgLqaZMp/YYBKg8ln8IO876sS8g3QS/Q7jOlKibi82xcLJ6R4/fnACf1
Z3kKSAYnVHg98iMu32teiSzE337nxzy4o5yCv7/7/iWQ2nbx55Hfxdqn43Xr
l0j1DIBmpzdUGsXkUbvhCfCrU9FgzSD3WUN3D50M3I6AZtqE2T+J14gUv6sJ
hV9ad91f1jTQJsY2rEyLjAs9EceriUU7OwSlr//PenlzxDGIVfdbqw6Ri8SM
iMfwmtgWL8/pwxKD2JLbsxRFnvRKdjV8Up53iGmH0sHmKGffBllpBFtx6DFh
QDqjblHawcDPfW38nS3pA8ipPpmpbTEd3kMUh6guK3q5wJsB+1ExIoBvElhz
oSsS9tR355CxZODiD0V0v94MHsQEqLsbOyQjghDW0t3DxWJZcflSzTo0+LRX
IgQweD03ssqV/jnqWv1fdYdHZE5qCnRvxyH/M4DcOFHJCCMCo/SQDV6QoRsB
bQQQbFV5Lygewb3jN3M+/5hLylwgcGr0/zzAuEtYpkZtx/R8bo7AzCqdCbwh
g5nNXlY6E/ziH3x1WObhSwvHUnYvFI3DFVgfmKWa1JD7fHlh4HYaGM4K2vKW
izPykqbipJgSNzyixGqvmR7R5BjSWmh2aHxe60QwPDH02P+5WVrQDS17ZQkw
53mPcMTiacjFz8UYqR2hrmJaDKcdFtxN98wtm+1aV+WTTMpDMv8evrBqmV6u
U38hNggs0h31FvWkjHsq6EzWveYgCrIUTN/xFvNZiRLU4ruOcIVqv4Gv+Yh7
IJRontEgQB1aN/Ukmunuvulk2w6r4jUuY11ds05/WJMzAghpdHLlt/8S6LIO
Ih9wUV4+1vzDFHexMtoaxgoL5BzFHRf6H2YzZrhgyaMeScWOPutHxmyy4yMS
PoBdf7Ik5WpDr902EISM6qQp41+Al0jU4fD5FYkMOcijXZlnTauwQ51WGwhW
bqCA7Mb6/nxcz+rx238fmoMdcM6hLSefdKMp16BT8XEnmI8FVxMCZXo2uktj
4tHzcy/C9z8euQIsKBjA8oDrBraaAjh5/Ejynxaaj8tHS6+K5it/f5Ou3IOI
rdQJFLgAVaOMrw6CHOAC5z125/OPRmfmJ2T9/ot1ypbOSsOys8skiWURFAAK
oj4HgRzEkaQ1g9f6Q4rAzsRs6NjPZBa+QV/ZaV5SifrNCtAsMrH8Q0XOh+y2
icGoZ4NIJARpmAMEDbdlMYN8UBaDf2s2SIKQxaTDfydYQPxlH0PlQNavU/a0
7yCOCMil4V4GdwR8fx9Ul856e1hrtamHBSraTl06kFEVKraypwut4SWUEFRs
r8GjPesC0RDuqwR7Fc2eJqhoSyxR71Q+aFf+BTGuK0kyj7+Er9F4JQU09dKN
tCVI23y2xxJU1bizXswnStqQ3DQMb57y8muA5XZH0I4GSQtLigMkXS6W/7Ft
/K2mTwtTEu5G+moEfDLs7KVAL6gvappOZq1paF4qxm8/NZtyeeii+aqZqeSf
5oqfMkzXI/ZImsafjK4EkfxrN1QEnwlM7YPZcsiRYUn4kFDGX2hZf7M6P55V
pLBqWGlnD98ox78LO9Ud3NRD0irs/X0lCbK1LmSe3twgl0nQJx0pZhHoSSwQ
H8ANTO+DXFa+qwmkUYhDK1o8pv69Wa/eRKpxmI3oI20cz9RGS7TjRz1ii0T2
DbbczbP4fEcumqmEUkVKNqznGiuZru5l/hQT5z5AFMLrEx+f6V0YNazybVwr
X19R812k7Uv0vqBqldwptIQQAddMuOZQBbB6ORvJP0CXm4Wqy9inWplvUrkM
ZoG/PstofqcqhkORBohJ/ld7cA67rvmK4CsZmArwg0RPRjJzIoHqmCZYKO/G
HV7vQFm6n9jmZ5Dty5dRe05mO/72vRYC/Z3CjsPKaFvAfYbMhcASpPNXHT07
7bpWtnge5adst54AVMh9VrV26eRqkKunIwfgo+Rdxrn+IkQUhkVy8uHOcNB4
FVQgl8W1RPobEip1TtTE/sG6s/f3LD73GzGSFSKxbe9iovCIyxRFj1cNJWNa
nfkuRFmFZT5DI3xlkPspcCELzzKKjOyl0/BkPfFFI1C1mdZ+E58pLYSiWukK
4/IfJlRk5vgykSuhTd3FLL6Qk0vXPRq9Px+Edv0ay9TtShtA/3BAHfAkgg7t
th0d6CUqR3qP/4qmtHoUslvCrgz+USWHmMp0eBymrpaEc/aSqeTmbuHo2plU
9bZNWIZfx9BbQjD5Tu1wZ8z2ebs3kTSgEIETx8qOuKESauwQ5Yalon9416wp
8t5/60D8u3bRza4WQrTt53dvO+xvgLs8RDsjDAhI/yhd7rx+y6D5BZTY1J7j
ZNlmEhdHlE9DM09kecTCMf5NNlT+jYZ1+ug0g9auoN/QjbXI/2bnLYXt0PQ0
GpdOcKKOe9roml41Va2lzwRLVuCeOph1d7B9C63i/a+QAd2J1IOJ1EXpRjU1
AMSaQuDpbl5R/uFOPQVx7PVVwl3pn9x8nMOGXER2vQYAhiNeoWXM+3fUyLLW
GFOsYVDLD/kFwUyq8LeCp36LR5CiNdkRurP9NBgSttG0HI6ghzAphC88ukhg
9CWtWdiAqixuCO8I+zI2C511/QiMJFsUn6rrckNhQSZjndcI1xTJ+nEk1agc
UxWOWvL8p9RR7Cttii0c1SSVJ/CWV23i5ubRp//R5nPtRPWseMN9X7q15szb
4+IJfYOVeObTP9d5Jx+vwo5ZrbqrM7WZSUHRI8jleo6cUaiTqdNP5D/Ttfia
xVMWBeF7OZ/fwTbsMqgyG6gznNI2ok7fYh6WLHACrNokYQU7NqrIlvyzqy60
r350q//cBGP/YZvW2TyD3+JHzhQkujp7zK2jh/BCwPFkJaOohhQjrHCmUYIG
cYsPqtJxuJZqvOxNfjQYyHCPSzfnBn7H2iEWTFMb+R6yE8sS7i99RO9bhRhG
C1kPKSvI2BhQ4I78wECN+yQ+/iqzKGf5UjjKv7C8h6RY+SSuCvYiHfdI2T53
dw9rvYHMLFZgTvpBxifVjTqTiTh9KBRXkE0XaqmPjs2PZNZmfhQEriOGxSw1
ft5CJQkO1hJsY+MEuzQlVjqKUIH3DTlVCfIytB//c0XisW0O/8Lb7c5y8paT
OP6NCjygUmOD1c7SpJolsYw+7P9dB1Gw/Z2vOJX01Bcfb5sjTSfUOJ6Y9w76
LM1IikVAY0mEEm0EozzWJQZp7sZzZeuJ3lzcsye3wDDNGUhufSV/z6tESRDv
9SRDA4eq4eItB7ROxnd8TKrR/9fPi3w8S/NWI2OoXOOraybMGsLeWucZAdZD
QRhHbDvZF61KJ/COaQNNctiOVOyEKC+U30ut+fvar+CaFZN8ZU/q3KQS37Vn
voayKXSvoD2ibJpQE3C87hXEI/q+Bugg3o7Yr3bCV9BoEGOBLsAK9jmcJPpg
ebMWx0XHcEve3SPCt6xFHYtQsKOhs0fZ8gGiTzl9VR4P6ZB67JA+LdfHkwc5
8GaVwbCIjYeAcqBBwtcPrR//wOpaTNH6BZwSu2v6lUvCzxPB65o4Jo0vUx+0
P62F5MhOkhctcc+0T5tRB2iWpMJ+zMrMaKyC9gQZ5EyhooYahfA8gsi/2w9E
sU+VqUHbflay4GZPjUJCU7UHv81BCV7nd2cGv2CTQDslEYGexkq5JgCGUsPM
hFFkTFg12KrK0oQ0ia99TFGGt5TLywLb4xgq+eHLVkQiCUjpeFw/FQ/yAZfd
dHAYbM3W/iSwcCSCXK0grzdilaXwoMUTfbuso1rJx8rtjVEsVpXcP4HKQ5oa
T9UrWPEw5lOLUL02MG3wnlYwC7Q2PPIAWVek0EZ3c081KVwjwhyUtI+JR/55
h2JxND/HHuI2Vk5XRi6M/wCvD7ODuZei7Lulg2mscqoU1YZJySGBfxp6KJwI
QZ9mnrb6FPayVnBRC4foJZkrJKJRmclim9xbQ1JBGOeayo9r5fhF/whqUGaP
amBAwKKxCp63QRfRY5CL2gzh2bQlTw2+cPP+ZH7/Cg7yqCN+Xxe5TRxs0WED
U8FExYIJYJ2GfsWyjjHjzz1pcLV4JbB1p4tQDTUSi5bNTNyXD3onlDEuTeeR
a5Jdj7zuBhovOy3L6abZtepB364LP6kk+buU422k8X5a9J17V0cwWQNAbxCL
BR83vQVZKHrHU95zA4W67tKi2lpkHXacfKfdpj0vNrtdJy3SDdKckFj6CFvz
TvTCTWCiIaiK+qwKoD3yfZaE+QT/XMy+tV028fz2I/dOFxGzRa0tcjiXO7Ck
0eBHupMoIRj4qNyRlW6Z6Vgv/nm/8FW4b7vnJ85bIrHXHW0OoJmN4UiuEsBF
RHn1ZuDNrJVX2t/buX+07f9jPODRDgoy3yxCYBLk2bA8hEubRzjbDf4vqVTp
Z75dPHLjpDrGeLWhZ35affj9zA9YJIMpzW+ov1N23rHRZiHy8JggwlyDuU/s
+88EN9Dj6E1rsj2uslzjfY4YFlzdrs4kiPbc8h3+AeVlxgAUHRenxhkEj1ZJ
LCLOqoh02o76ZskM4787arkPqpXye/NeT6sn3lxHh8TQ5JawKZJtvA3r2xfo
jk/3qEP8kHfVlRe/t5A6QXkBYSI81ryLID7wW/v0CRu3naZLyo1JiDP3kFxj
xhgk0TES84dd5Q4lCaa1QKWpuvnSu+7mROofN2egk1gJqvHsa0YBBRMrV+fM
z5sTMGvfuK6LwXrzNalfjqvxGV8iSK1CwylWTzEogVTrY58YfRjqDH+l2lcz
DQllzsqtrM0RiTgt5I6N9E/iijrggMZAqee6wD/Rn/3jgdTJzHuKmdvyQjgh
TmEqvxCr7NNdU7h4n8ZKgbav7zzGkdt2Wm2HfuuYDasUWO6CQWucqa0VL60T
y8ScnvJDFQ13rvjS5ulscKWIDjWUTOTE0uotUBQss6ckqBm0h0RLAFiK/XQo
88qVDVqFLiWM0KBQdU2dBJdyNoYVTg5gnEJWEslONjrcNNpIq10fwhbJtHF8
JTfq5hZCEmqnRilMFqbbFG7vs4ey8bwTBECFAaSvG4eZXx+KXeUcrePTyRrn
fi/JMrvsuKJ9UZ9uzE3gwuqW5NHAuD6jmiT3ZqhHp9AOgshMhmMgP7D2MtBm
Zd2pl49x9YoYediJZBI8J0V2viiI4NTFBXg2akd4VuBHN3LhSL/A46j6im4S
igeKH1aSOTrv2wsTGtUzxNa3AsU0a1bZKLp4v+emjOhTR0ieEIsVXUrmWUWN
Ptq8yMD5lHzmCmdHDqeE8gb/CifHWibsQGjg5O8xCFuZpQEZ0Gyb1ZMAD43n
TU8zzIfQyKDXrn5OaxA8k90BVqk3qmUYhpEfwt1dNKEBG8v2Z3V/7ur1K1dY
89wxhfGxBSGFo4ZNFS1jRNP0pVldGc6WcT+NHnyBPK6gH8u8nDTzpGd+w+Qu
C19cYp5+0vPXW7RMW9XsDLrQoNQvoyAe8GsoZgGwCTIkiphQ/ozA6NQGhg/0
NhX656ELCXN1wtsepex4dyr6uDmy2ben15wkOwp6UlvlpQX5UTPEULaQ8Hcb
rfmoKIOhyNrDGg/VOJsbritHzRcLgmPv9jZ77jWqRi6OFUuHdKIpYwYOcnsR
TGUmPGfLDW/AAFTPePQdVU5Hm/TpvrlRVJR+jtdvfq8Hp1vD0M+7sRBCkXmi
sdqiMtt0ENahu9klxshy2SAoJaygOD+ZHcW5QqPsn4DBpZLfoz0Xqt7nrzD8
oHovMurDo++kmBDujggekmZewYo+Yg0VXqPyqmP8jhqzvjI+q0lZI2nb8haz
P7Sjlob2BfT9HRZee4vwiZY79h89U8VF6vKt5PDqeGJUgK3SvVOLzBhWbLJ2
DGm0HxFgvrTsW93HGBMNBiYOiLjmItbUmSXs0adO5RUGi2MWglRzKZ4LNGLn
UbtUn6LgPdrU1dE260mCqYK6jpVgKrU4dv76Iz0zOuEil5jo5mFYLlMXrn2z
fEjeBYLePj3WcujumDbDT8m2p6M8414B6Nr1tdJW9ylU1+qDyJcA1ieXPrI4
mYJBKffQxQwQ+18ZO6qv0FeQo9TxIzmttXKcFM9x4wDmn0C84PrGfPNq1Drv
N+gxFu52oHXUqKL+riIfHNbICMFbOmnHZ3HsetlsxDl8CIJ0lKfS31SzDqCW
ZDpxmFfU/pcg9kzCAoFRcnXXL1quqdRcVBShR43wxY8x1d/FG/pRpL9txzBV
ljBnVHYDOoxF6P5C/9maz89/VWoJ+0G4Loi3BTO6/QzjFQ+WM1fK8BVjFUGm
zKfAtI2CywPvBa8PzQBcyBGpET1mfUeJ8fKtJWlbZIENYV8jDypjudD6L3ZF
YH4EJxnEyO87vndmSvJyT6zqFjnimCpkY4kPzdm1wEp7ZLXQ/N9i/8OYwLCV
OM2Am7DSTGJU1Yv8vowfTHI35VEi3pqriRUlrgvTfNMPESv5OHwKk90V1LSN
vvfoUOJPF7UlXEXFEr5tyLoC+97lmS0V+6pTmX766x7VrfOYHHG8WcFskrL0
PXMMbrUUKcFx331ZJue4DUXJx6J/oavig1cWmABu8RSDwO3W/7tNhVuwExFX
MVGW6+WCrQcQRqt7h4g4zsuLeGtpl/g2MpDzbvHfk6HnoW7VZZI/yzWPslr1
M0MIYAU5WUyd50LNo4NrTox5iG+0jQZOdtVQaPw7Dd/Bk/U64nDBVVrSd8/2
2w+YAlnNFKfgl0O8BK7hKOPD8FHs8AEO1A3OEJKNJQzmkcYCbQx9cDMfnNRo
WVB9oJsDt5eXvBkaXR1hQHc3AVr28j3A0MAL8ht16N1KZBK9gkl0gJMpgbau
hmW87/Sp0HF+bqHaUZFSbpxuO2GKUE/24IT7m7X9kVvNCrnzt+DMxp2ffMwM
qAHeuoCnevTm7scW7/NqGzufhSxnUbVwokNQh0gYZSQsLHpmzJKhLgfpDhdk
Ti5dj2kp0NcTRgT8gnaERsuEfVgWPKmtB7CARkzsJ/66F2j9AcPo9lGvLWZM
9uyFaT53FaH1aJM2kji78ZWkWF3ZxPZQlmxCb6e4+Kkg4nvp+2rwu1mhUDuq
weqrhOha4OIfiyVTjrL6DVFxl5g5s2/WoxP4PjP3VIs4vqNQh2i+8oI0miMe
d9cSh9SAObOkic+z/5aVJtnwogKYX0duK31lKjEy+DHUwDJjwfc/fAcYGirW
BwF28Ld7AH27RY5Vr5POtbFzugCZrDQH2lbhAChQ+LziTWJk7SXzNEdcetBv
S0OYdNiMJzGkvA3AeSlX1y/CaZkCsTOYa1/CskPy3hAu4MNnRIfJPVJbTKJq
juSdAo1hLdJMpTIUEygf1CAIu7wwBCEcOK4IPMehHX+VX6WdZ1MlnaJSzw3V
s1SVNAd9n64d2m4riN1+uKXGhiLsUtBKjumgZ72b3Df6y9Kx+gEljILPIog5
C4OQzfTl7qt+XddPUCu2RdqYePCRChF/dhwNpW5IZiYz+JHTHQXz1aKt6VvY
SJj2JXwU3Bxqr2LD8nz6nmqCU0Xpol3ueLBoOfGt8PTKYK/O6Ou/dMOPdNur
vb9d0GKevKQ0dmA1HQDSPSFE2LFhLiWbGhaV/VUsRde5SxoXbYAgHAevu4xs
DmYYCy3wdyAB4i2+NHqXcmlN1mWJ8hpQtC2lPJRAUhzdKuPKYvChwLCeD1cH
7jFGy39geqF3uwY1IA+zl1v4y8k8oa/EVFL1AFDEx2nHK7ceumVymm9OR6bH
Sf5ea1/mlaONgCfSrbsNvlM7mNcbnouaeW9XRkI8qcQSh769JhM+FRysMqpq
0JdFOAU3vhHgJEgagQe7Np5IbTfZUS1NtmYcteOvcxpDiq55OTZWKBjP5n+7
l02Wm1e3hxEefSJBfA/55W+k6vWNP/s5H+cO4Oq65OFNFdk4uAvCkXHvnfJC
r8IbpD7kJlscc8SMnNOfmOOMpWusRFeqd10wTusNI2JBmf7UYEoIV2osTKEa
5s7OMIjnoGsTPKAe6lS1mRIAspHdFneGej5CybMPLqVmD9dlPuUVZHXrQ2Ii
Dpt2FuLkwm9yaRRzj8Dr7DTngfvSoU7/7+G9sPdQ7uQy9JI5s4FXQlqTiOv1
amu0//xqRjLWC1JfrKnkxNHcUKxA70M7k/ji7XdUQFt70yuXFd3u5j16LFv1
45j1Dw2ML5k5h32vN10M6fJf1sHsA4O0h19EF62MqFEQlyX7fN+KMHwoXLFl
6+Nk3PJUCH5vzGbGY7RJcmmC31/igZWnpM2GiKqrYoz6omYe2BzdQQd460UB
yh/f6ofct0646FKZ/JTTNpFDwVbuI6tCD7IOybDB08oDcpbA2oFDPNogDtzn
3lx2ovzdVW0T7QgDQ/l9cvyjCL+IVIO792Ifh8wCwMVezYdD0oc6Jqyg5lN7
V7qikCRRBvHrUfMGyALceZePs6TubiMB0lOYfmM/6zZkgXWVv8JuQ9cuCMt1
ZB9f2mjRvqeeJFASWmo8osxVrQzrDJrlFIjj+tuzL4l/Pl07GGfDfhGL7HGx
rR7RIF8whrW+mB4a72lTHXBhSN248QASGru9blheBgyLVESy4lvjn6CyrkUP
jCJjKDJ8BthWRpxtxP/Iexol7hOvIT1MidipEhZwSIKmKJVhKMlnDva1Lska
Y+L5eAAJzkj6zNl8kqqTXBulerFZtMpQst/sFnMZjkfzt5Xb/wpBu2vC4V6F
usy8dSVT+62+u2SOcKvhCg2J2VUJGEaykV5H+uEkSImrteKSgkYV4vXFjxgo
S26Yvx5F38xQgUQvIUOqNb6kqLDj3850Uiy0L1gN7R0SjoCOvjHSIyimj9+O
Hh21OrYeCiFTnkcYX9EfGicL1yhq7Y2n4M1XUOPlSCse0rda55Z1gh3ya3V5
NWQn8d/ssU5kAdk+88ywJcy02vT5GyXzwTZKSTTG7yOnh3btqY7JkYFcv4D7
CJBaQqYXcHP0pkT3h1R+9Zw0jphs+6jZM9IBgAnZWKFFGHOaAqm5pbXIST7n
eDmjv33t3erZvQLM3lPBAZCVwf2P9lcU+7snZQJQDeCYa190QuCQv7HjoH80
pAog2LvK4fsajQGE93OzD0p9jRHMMyB4h2Hnrdv9gZ442Jm5/EPR4U8LRqae
X3p39I9oAr8PZJf4xwfa+Voo1gHwdnBWhSqQHnq0p2LXj1LGo21AOuA/i28T
OCROZ9gCCJ9WfV6khBZLGsSCARUHt4mmm+jv5Jay4HkdVEU0W8INIGA60N2a
6MOo/VGTJ90IdrJ0hAKVuoSwgH6g46m+BYmz5VRGSSpbZl2GAeBT+Folu+lN
+VmS5nF02s2JEUZEItHm5fex6p3l44cYxIuj0mDUnLL5gfmwcVWJdYImk88I
OVBVNSCAkZ4cFXSGhz/v1ioCfMymNSQMdqkQPRDbvPYurLklqWcXmk1XuFtG
/kDwsWGT1PLnUyDtVF6UmR4EgnMSqiJVlm4JOU3HAGqd17Kl8uX0gBwO7yuk
jqSYKltLMDRJsL2E5+wL6aGMDACIp44utdyGkpOPnmZCmAmbe5Z+1NRpcVIh
W0Mr8E5sUWCkahX4mv54By/SQo+sqS7kHMTdvrGodNTG82pqqyL4pk5+G3Na
tIVak0OcqCykU27X6hN8K+lciH4TCOg+yt/98vQWBkFIvabhyDPnohr822s+
4eScxWOUlBs68AaQE271zZCl26qKGlRSBZ71Uk4p3axEq4bgDOG3p1ElgXqk
9+plm+/nD7R9tj2q7stjlfmTc9boqIhUWddNcyCKsPRwW9nzOJBUpmGtyaQC
HfZKVDEfBCeP8BT9hWB7f3rN0atCj67S1azXEjlaKObps6KtvRfebZsS+i8m
QCvgVgji1wiNIkzLUpTvT1zVSC8b1mM6/U7PbLHWCofwg6v2aNJmHaAJ3W0W
UTbXw8EPYG+SzE8TdG+haHV9KwGPKSXm7AUAxgcsIfFd+6WpnIqKW3z9qFRD
bxaEFkvy910aXK62RGn0DhfeB9VH8rmmjXX+pvXVDQAPMcSxauWidyMxHCAW
8FQL4vYFOT6+IiMguAGMJC2/Ju/RNtQVr3ocO1q89wLpcLSUiXrdjuayJ3j1
JrbQumHs6EQUvwQfP6AOMHKbl/RtM+Vt0Ju4roeRn5ssEhYrfMbcSKkGlicd
3BCxPTrrGcCtI4hxO9iGCBlKUHr+mJdi8oiTwknekRF2R23205CJFM6EJrXd
l03uxNdJ5foNq42IyKEPneziTiu5jy1dq6VQBwHMH4xfIi1Wo9PRHGPlUWco
T/BaA1X3TfNlR/n6/qZfKSLAozUb4yLZbQQ2K/XKctP5zqmnWaYdd51whpJ3
XTwPHwh2WFILoH4jw1/YZfSNx188NYN2z19Y8cjXkeAEp1eTmtfwQyjYlHVg
md1K2RghASvSTmw+L1DAgKX2uExGB+0wR8RtB7VnNnbkVGcYE04oaXbv5UZA
XP8bV535419wQLx0Hq2RcxX2zv3ogxFi3FxdnkY+zHjUS+Z+a/zrgdaL3wYN
H2vshCRUfx2eSG5jC7OM5t9RlgJMrCglipd8w4jXJC0LfH93ORlk4n2tM0ro
VstVLIgAxLI9ntDGyB3fCbWGGZDMp6a6aZ4Ux7uSBR2ER8ZmUSwrMM+mSDIe
cvsHyr92Xtho48pekl4Q1B5xeVU5vubPUfY76ukzfROZDo6tQhPM+61lkL9M
2Cg+BO36EbsOIQ/Zky19nZln634IKUnDbnj7G0zcnymPNTbn4p+AQhRUENEw
HNwId+uBcwpYgkwWlaEuhPqYn5rjgDQQ6zZe0jnh6JeaIj5q03rd3iUQToCz
n3ypkszcf/dkKm58z/ea/7LzrEZiviRhfFsGWsBvgIebBM7nxr3pzwVPFhB3
Guw3oHN/zAIbFPfQekjM/KDbRInCsU6O78lnWzSF221fFd+sWowlLgifAE6i
tIrsET98sT7pv7RoWTb3rKD0oKRmmq2O6Z4EYCpVEDGFi4t7vtK3nYIm88Ok
CldY+ULRIfrkyKcQvwrHzjnrz2lVN08wXeoKn0nW2ol1K39tSrPMunwhV28H
p4pUz1Yg0ReEC2B/+XKVwEiSP655a5itxLYOi8k/15LCKK6PN+lAAy+R0i7y
j7pmB5HE/Hnyo7Qw69l0w3gjAwXLN4TPyeiLI5qNupt53nVJqCB22zSvD2w3
Ds9avI1JhFWe09DfOd6rLm6W1h8tr6ucpKgh240/8AzXK6QcTplknyZFaUT5
NICV1yk5AnJh8r1elzboVWbEEwg9jTD4RB7Ag8stNg+P3S8UB1jy0D+7F94H
RbmJQavmWLh8ndNR8Q5xFn/tBIFeX/4mqfgnNUh3IDzCP5rspCnBjY4uBMwT
nxjPOvZ7s5UHzKHi+7cJogKrrFFRQP3QxaTe7bDiQOBFZmNzLHw6fCd75xzG
OkRCReSKRX4iEHRwwwxoQMFv7CjYK25Lm0nGsXpcYQfiTP6gSSjDNg0avTyL
55DXTmYR04RghVk9N3xpaAI636tk8zJokecOlsOtVZ4TWiYMPnhzbxyQQ2rX
iyl7VaChWx2g8M5nNOzrNNodvSvBIpMhP4HnksKbLf2LLz1G306hJT9UtzYz
fkMw8LFvXrdDoxyylM4B5RXrjeo9dxgM5L38sLTKmScmRroDg5Ue56Ranvox
njLcspni+ValLDesgxB1O05rqs8LFV6n+w7ncPVluncDHefbp1FwxZymk87p
KVzg6Y1brf6Ze+SuSHCkLawH0qNtoLllEz9j9GlL9elQp1z3viXZIoC0B06D
xc4+KAVUtlX+a19mnrA8NIhbelQvGJNqwk8Y5/WdK2LDeh0f10camw2MyWEo
p6aOKhTouBxZDpfN2+rZOLw34I9cqbAmDseKgUwEBDWqBiPw/f3Zd1GXx4f5
IrnlCPWOuePeIXJZyG6D7IHpOOsDifGd3GKkldr6WgF62svEOfq++r2DMmEK
OnlmFNtLSmbVvXg7OxjT6iK7sLGh+2bk12T3S8/KpAVvVaR5i+KaxJj/olbc
p3FuKlOTSR+fSjF1NIYXr9yrK1f4JFshQjYpqAnFlG7FpOp6lqUwI1GjkZfJ
zxRlKdVXx0PlAhWBrULT+nji4jun1j6wAQrNs+3cgYwbZQEVQtSXa2g3/A8W
A93OoflZbn6lSlOgPqqSQUH2BiPO/Ng0aU5HhbA62jDP9eQGASJQhSjSvM0v
mze21u2z1AwxjyMyw06yg4kg4zN9OZisRGVWiv1Elf31Bee/OL0GcCAXnNYU
Q7bRAZBK4pVPE7Y7zRUAEnm2qg9/TjJl83BzasdEXJ1uQ0Z0GJwWnUf1+vKG
vc+crK9utFgMoRy1H0+/WqvjH+ARxe9l+Bwqb2XL1fo3RqHfR/vnzbA8yMdX
5B6zfieeC8TdsvbXIrMdlUtodDBJuQkzomiJgQAsZZ2lfmKa5BBOxilsHgGX
H61V9rBVm/TaagVZ8oVS+hrAoGo4F3l655O03+qMMR5Pd2KKxevXHAaG85gt
IJ0CxYAXjpfJoEPouvK9YRv61sEh7iFC0XleVp3a0FdiGOY0JVjuu9JOIZqu
GI29O0dwWk1gWgz6m8Aao65EFENmdIfelEcMPBGRPblF1GOhihEJbsTfx8dR
0JqN5vV1yeeklKIip7jhZvS31I3Iu2BULDPqfK38S8PmLYncKUHGGkciHyTL
ZwlXj22oxiapNxlBAsVPnSxiT0TUyfz1cljpEdK9VhT4rtNct1iFxNmfWzJI
RheIBCUMBFezlW0CMmZewXnvxTQwTKHBocmJsjMV9aIriP0ehPUUi1nmO1lP
IRUNxUS27pvf7a2sBQjf2ErKnO9Fx2XIs3QYvvKlLAJtxWzYDpGrkTSvzCcu
FuvhlUCPSmkMPpc5ivXkIdb2SPPCg/ISC4FYpR05VFLWEwB5HQMJdf9ZqY8o
rNdF9cHTiLTiIB+LPrw/lONIfP0XCoRDb+UwnJyndt5ULxb+jJqXnec+jPOT
kbYH+T3sMbYp9nV0y1s1TRpAVSpHXkn4OqYrRRuALBApGhjqw/PuLCe6Yack
BYHivnVK/R1rQDGIE0s2iLwRdweDmaealQzNhGJnBAfoBWeq0pkMxTfA9Fda
hZ8UTll5DY4oGu0cgPfab+m/ibHTxttAptK+YHEL0hXJty9FSA05iWfwMSr3
frzbAVUNLjW30A07AEc1wz7LLIdH6Uz+igJp/62MoD0u1xWEcw61RcJCkmWv
ZrbBV0zRaDmC52Rnst5o4LhnEE8D2xh7jhwzZgtKBOm1tCnJHJF2Embsis+d
1vvTbfTwBG8uUi+4QVawUSgfdCbDWBIgFPqtkBnhvGzCOdSKYakDW8X7hRrw
ocxIQt59kL3cPPDNJ1d1ncm0eiEVF/84fLkQG11G1YBv0jVLUCeqvrUuuwCY
oYtEr3k92fgQRxxBxbgiGBxFFj7uKSROeqQaagWxXQyt5byxr78jl8p1W3OY
eO6wCauBi8NTbyKAzuPElMuf/v0dz41VKg9t3aO07Eae6Oyj1jpXO0f8qy19
1Da7Pf/OEjvEGKVHGNeMzQiiGxUJYFOFM1z4bL7gvkTaeyudqExXQVQnOnPA
vxrIS7t3ThOEhKWw8FhWc3UC4C8xZDzicCUcJxdJIOtWooKSLVofyl/dAj0g
FR7M48hGv5lYzco4mSHcGXy6XEzCuyXIqTnyQ4q5QRpfAJYlm9c17Z7d8Z8G
aPEgKGSt5+0PZ/tlgRCXOkLiliyW24mEEEJfA6xUn4L1G9M1BbsIXYOi/Y5R
E/RXpcbR7R7A7c8pzCW1RH375pFYyPEgVe+Fs00EWPFJzISOy8GVeu6nunYR
WRnRcVqtcoCQhThq6DcOOZ+osPCNO76Jy8fGesSCq8/mGN77N3DKbvcEHvUh
xx/aH6dj3KO9l469smUbW3mk3bTp1Cm7YZdfGD9RIVIqh85ltpSXQZ7QdWUo
PQ/b+HauZXtGA0A/VNGtRKn3WPPvzX4CPP9wUM3wasWjfo84pLNpsrwLVo3e
BWJOWTnBw3VwXBfaUyjDpA9QZkMvV73z9mFVx1irKwusKKnW37RomMEJKOxy
Xlxt4PmJO0RcRAXkL3cYo35lI6+hR0Iczy6g2f1X+40KfNUoNLCSPuuft1sj
HNA5qoVcyOmGKL9HsAL72mAk/CDPKzAZzEg3+9FJ1gH6KZ2+2wK9ujra8XlH
0qODt6hZPD4IeId0mbO6IoSiOfrHOtOBzaXoKYbf6/uwh9TJLGyKF+YRzdWX
Pq2I+r91+7flJSG20u91QziUZmU7NBqkTxSTbG6wUyADktoA/Hh5Qvo2xYia
uE3e1xEbrlu5Y2ZgB2vEi49umI5Hrp8kEQUCFJ/lmOZiQ3ksKhja5CRc59Fz
trs4ttlfdz6uWzKMskMZy5A9R4PITTJhQt5F49R5Q2h4jDif0XcDj6ZPhgk8
WxJD2w6y1TYnCL1pZLiqywvizPal5WWRGXF1hpO9RdWqHK+cscLMr5cf2ljB
7MOHY6KcU1RCV/kaV519iC/JdZ1yWXxQLx/vWiPKRdXLOYRG+ByNIeS3X+nq
A1rawVArt+Y3viRucJrA9hb06T/W/lOAIBM0YoNirlnfBMCZsmvO/jQ7oMud
UNsyp8x9UUtTxgwtTIMKQ9ybMhHkq1iHZQpcaZwyGiOAy0hsk5C8BPRPNkL3
ZAbtqHsuXSSDc+Tmt/deSWMe7V4iSginBvvdVDkax3BWgHuWEjThOOUpmB8A
ptMmhM2shuV05Dgbrki2gNAT2+04yRrwYSrXVVaJiKfaoQz31gX/2vk9Kpov
T7C+6LiQssVnSB6Ml5xNTmBU3To8ifeeHd0RTxG/E8w0kYtdRIMn+onpUxEo
yIYoZ3OxzzU/Eaz3+QilXNWYbujY5+8vQz4b7n03v1VBVEEZQAQlIHU8FBO0
8KXuDy36/wdML0o0ga7PYwAO0oFWonrCA6/iRBwwgRv7LNsScoyWFH02as8z
jdtn5wL06eREzJajcuERpuZoU9OirsjCy0UvS6812SyfXq1AHQc4GkbfV/Sz
p8BLLGV/TmiWN3rcjjUL1+meaKCWibFKnPGIYdcGUswRZyg7e//b9jhrjiFc
zvlqs2y2J0Njt6YcXf4q/Zf2bTp9g11/60lgV8ck1FpkQKy2kNPxcdRgk/oE
XaCfjblGrihlwxdFVQp7/qxDWSudZgeS4d35SlAFnuCoxAk51Eb7yq+87bew
WmD3JXzZVgmx4B+HZLIhFzOkRYWM2qPIMa0iZXJ2siTg7POD3GxtkQCpiNDt
RmgAazEq0S287g7m46goAZCl8WkEtYIJ/1dDeWdYNwAu7o2OgA+vv6RPU8sP
K2OIz0VdYuZodBzIRcMowq97phDRgf9mGbYCrylrJeNXFQ3JXJlxowRKDX+V
EADc8SZ6lMKAbBWddBXlrOB8i/eGWRBAV3UIUEL7A1fFy7PkIC5I2CrEFCpr
3aj91cmmtmOPs72p3yc7wk4aEPI71LK3YENFGZ699n0iqP0KmmT8Iq016/2i
pF68DQe18sx/V0u98foY+LsR78GRKIhw43ztvHYJKrHKCb+Ud1xOD4he92j3
v9ffIjynnuRPFoM+vG22ISEG1ic4fccV5ju/LavLT6I2JfRkjVRwK8On0yys
V/VCEQT0bbX22ij9I6mnSENgHposW9VVvmkSq6NZTBBKShKn/RWOXW3RglWF
kdJ9DDrXBJosTqJjFyFwEFNuRy1Wl52zuDbDzijS0mDlXwDRvTJIcdQfrtLJ
74koFXF/VsHhQOl4xTLOjamm/h0XIs2Qjs5vYyNDg+JNesp4YpOgqWb9ZifN
gKQ9vQywo2Hu4DOfCxypWeVjV7bqACxknIcR/yUNSzBMZY1lOPOHx85b80c8
Iv3ehYWh/jrXN6LLRaGdv6r/RenCMKq3nTiwlglMypoH51GjpuwhJ7s86b6s
2zlXjqGid4WDz0Xs+FEJ8orx6Rklph3UhbG+vXh+h+Z5ZPYq71y86ZTyPUrH
kfiUWgofr9+Upo7QokaGDCNOuG0VxU720eMVWi9hk8zBUAE6KnZmB8/ILRj2
6+9XUU0cjpTb+iS8jJxGj+c6vvNMblyt61eHAf67zDdjK33gbezLFokrS4hr
qZIJ3MD/yOZNqllEyq/HusyBlY5aYKm10oWewnADxFtWk6qfLEHSC826EyxU
QpyPyM18YkYsxTYVu9sYCbFcFcw0V7L7LF8qOWgutVaeCX0x6xaoqMYNPuKs
o6qVerMukqkJm04GVW7ybI5v2ipBFFYNC+vSqJD2x5OkkRIFENhEt4dTpO8n
nitDngejjbMDurh3u3apngEoBRdc54G534bCCbS+6PG2+FUUjq7RXbP0m6P4
3tprSs5BKhgekNvPaL8IfHW4TEa+4ViS7Zd8SeoM8W1KZjYZXKmTyGTBPac9
5TgqHh5cJAS4aROELASBhY9UU1twJWr1sQ7ROS0PlkQjqjaWRzhn5BDgBfm6
JxhMRljN5KM97OvrMb79Tao7rljH2wE37MzHb1WCuOLp7FKpKqyN8CzCCmFE
8zhoC6ICXn0D14Ubkin6tOVX5YcRU0orW88QJFZVxmmFwAcX4UAdkUef+ay3
MAkPMn2lj1FRtJevy4XAtfBvlo1BLUhdhTCMWob83KU6uIifudLqa6C18eE2
E0wvJpPsuhk4DH6ITNzs82tk+LVAwtITuWesxgU/G+BlaRVxlYwvBtsdMfoq
zxRv2y0w7EDHbK+d6BQZexkrcSfmGAdBY/EziTT0XtkAH+jcGo199FKZODDN
HEdiVuZ/5ZZWyNCI1Kw4UEUCvctO+Ia9DK8mQ/XEHjRKI3YWeusxVLBTnulH
gRrImxFpgb8m7wuXHfYV7+WOE4jPHzZw6x7A1f4lijjXIwQCteWp+BHXiptR
9zdqaaEl7x+6TWn7hqKNVduGp3bIeEkbX4jzZqRlJAu7ZL3CZjXLn8teKCyt
s6zH8Sr6PrsBmciL/PDokU2F7exGhMnqszI9s/j8tB2oF4oJtdcnYSUWqrFZ
efJALY0iDNr4q6FEWFhedsz65Z74YyuCD2cCMt0Ax346zIgtz1WRW2vlLOr9
r643QxrEQiZbysFYdXet6QWZyxjc4B2vba6/ZxnK8jtla5aAuxDJDGZBGRGc
MkHF2LkUUyaYQXrf87qpQZd8uCtJQvdCrsmrr7/WkifmBkbF1ENp3ubaLUG+
CLXP0vl1p2MyHOJGip7IbwrQKDLTFiISXoY0xlqbTV6f/qbsc+9TAVqgEGaY
QkzxEwI/5zhRUSvPq9IHDNDduXbHFzzXJ0mHGSw/7qtjxpcahxJvZFLspHmC
DllEDqC/RP+O+mvHpkiMP0O+Jvg193BeSo2IFWBX1ti7XD9lUrtFq3nk3wlk
yxi1Qju0MVXQleBThnAnLxvnIQ+1jU6S721orKHWuJS8cMGfWC6Wpe+KgdT7
9tsk8sWVOkkHJclG0RcyomXZtgV0PLWYBiDXB9grGfX1WQttuq32x7ftWUeR
mrRNqhZt3ff/I5dS42KsEZvhrQIgQoZHGcqchyCD0uktQyh7OxkYvtGM/Xam
m/FDS2592+MOPK977Mb6dfa45aDwGMbM2GziWPODvat2JJbqUFEk+B6VhJ0A
RLPwRQQXCZnnhaxPvYwyJf8p8GuVSYSZ+iMXfZ1xPz+uTBqqrkBYotMoh75a
lY+5gYuy1XTKK9MYCSttaGOiYZXcDSIKNrP+9rvX/1eZiNqawsdiuVsBpSJm
jXeOadAt9VQAN9/jJbCkksBGcGf/waXFO78USrmU1dQ9jj79NlOJCX9txWD/
ZDKLKfr6NoeitlSfDSrdXjr/UPNQrx2Ewa1yk3jenGGQIMb4c/22nvAspFiZ
uGaOQk8dSW6HS1nmsIjNyrAaSdF6Pz4ZNA+BHQIgKp1W6s661UQ91yt7pqMQ
iuXcaQcp4tkM26TiWvH0K8d+4I/Uz1iptST8L/o3auD7xVIMIB1Vw4jeU8GV
+z2fqqkcsHvUOWd94iXDBKuPBbyV0BQVbfkbUQDamhoZKYw4JWl8xnyJQ5ou
wgGh1tKwMSbGd0ydfOedjFTASAldLx49Z+LMKB+0+ZhIowDcUI/SVLANFiCq
1VK+N9N5xgMUR1t47bwQLotsDp+NhUDCJTGpLu1nrlZvEF6jwiHJkpPMCgo6
q+0C3Ez+L+PIhh/Yrq+fAYIn3zbkiZRQhnaFAhnIyY4dtVvCqhxHgHs3TPx7
tbX2DFvhfA1iMePjujtEgGmmV6zPbBAFWZpGhuEQH1OZoIIiB9qWkvAOJ+6B
rKA96YMLYMQ6FEtraRn3EFgXdjUgzR5bK+qPI/Klwm7Ejd7CJmsb5XZwABi6
062vrJnKmYenacOMZWXwPOAvilRSnc1jYh62vrC4Pla/WjbAdufv40RZiqFd
fBBrQmK6LLj2XCh8po/bIHi6TAv7+OpvLgSNlqpKpPfbIObgrh83t582w+Nj
aZ4kuieJ+SQamTE45JNp+Ukohgx8CT3RzTpQxGij6RxzoS2t+GpVlqSMG0I6
fktS6g8zA6aAGbMm6CyRFia7sy2/yUqP6zrkKI+LKJP7zY8vr/wmzfYJSmSZ
ERPwWEffeQIiVweMZ15J/oq7HmJrWJLO4TB5w3wkOjtVOqc2pXhY3oGIjFmP
+BkLDx60pjv2E/VSaMC9wsA1fJTD7ZlT0UEI50QBW6q5TIrbjo91DUBLeS1k
MeAfCfc55tY1F7dqexHtxWqyefVQz/BE+pngbYCOYVueBiYh/4O93xxGPeEB
oifkX10MS14RDZWrUG4P540yhbZz7sVq6TXBdvmaw5T2JXIYvfRBfcsb8V/V
woVMeDpgfdjImms4dOEmDqk3jtgUW7PVL/VqFLvCVWM5VhveD4Bq7c0+hKPa
PGXh4S4pxZi9bJt17fitF/Dzc5XgBT1pDXX8w+X8SLb+Q1gKnWTqbdW5LU6q
NSKqpG4eKgMk+WNI1DGLUcCQYKGPrW3Wnw5C5mclsSLlS4hgarUjo832Z9OP
Crwb0aLywxft9vdFOa3iMNacylTMJNZAOntppzDwgfhQvoYUGosP9QLPchQQ
Bgx2wNzx+Ph6+7xNPLnGcRcprDn31ZXCe+W1e5ArwBuvffemhcWoIvvKcR3x
OszzGiusNFqHrS3GdC5+cXSI/sn4k7sOp9Nrk3LLkhHjU0U+BXTYrrJTnmC/
2NFVuR4r9G1OEG6h9CQatnD6IqoWCVqPjLS/5w1aSBryckTPkMo3NQpCHsXy
k97kKyIjNAvMhjKxgUCJHVxahZEKKgW2RECEnwj7lgE4iIgHfZ35yeJdKPWK
phsBDyBfTH65zlBHWZElHxcAIubceqWs5gJz7E2Hkl4V5Lewe9nqfFyUkOXC
GAnzXunWbCnyL7TJ4pPUDy6KtBXJ7EDvnOtPKWjwqtCLZ+9W8hvJRAzA+pc3
+5o1YZ29fEu9uXAUhpzaXjd1fXOe7d8iuewkBpzU+UCDSJ46V+pvMN4IVrKf
Na62onczdlmT519ANbvHB4OYA/XwfZJg1Vq/r3K0QCpbYQ/jQMyS1PMZ4rE5
4nF/s5FfMEVpZ8S2Vbs3oJ7MNYeIQWfe9oGmVbQ0IcjktEpqu+/3TOkZ+zE4
BptmkvK3OFxPNIPiENdRV+UG3wo6Zs7P26czDgSPAl53kSXHn0ko7DYuoqsq
Sktb6Sd1hPcBARu+ac+SiqLGv0JB2gQBIOyWH9tKk6KNT254fIgFLnMatBlB
e6hcZfh6DIIp2J9tFDXUf2q+04ry3u+756l/s4ixrWjCd1wnT7epXa1QYrrw
YXZz/pcj3Rya/Mbbh14NfiranF0bxDnmsyTruMfKhfBw3BiM7spefAV+vUv7
4e04p6LkJeH0XKmlDtXwc+jJx0W7FEkRK1RNg1yV2vX7DUEezeUINCQ11tgj
/tnupONDKzr79Al+ZLonqVkJ4H1aZ0wfn/pEbAq1BEtF4hTK6Wv/1lb52vjG
lAN1wIQcufyxxc+tvKu34hNDAts9lvF/zkvDxy5I1XAEDO518nhIHsAgDJvd
os91NLoBhZkQbAYrS8Fk746tabAoYUYogReOraE8m0hOVfuNaQj9WVBO8wr4
xhnVEvS49Nz4iP23NDDGb9eIkSIrV8LbeRaWs9FF3MY6b3aUAc2gd+s/hEfc
YEzh2tF6e4pcGoPkAGKBwUkOtpoyXb07w2hYwyEQB0FntE8AnXbH/9a5Zfyi
a2tLoPy0zwQxTyqWG7/pcggeTBlP1v9bhnAgJx8UXPHbB2abVRKWQONrHSKk
4p0BAj5wivWpGaB1xfPygnNXU6xZJWyL2pE53AVUYT0Sx9oay/NA4rXVbt91
rxVPmNOTZp9Zz0tamaGgZZYFxJZ4q3HFj+T8/Uv3AOEUxBXthjAwl0C7ubTP
mmxahHOJ+IImYcmAQONSg1UWtk3myYL5IVGwcqH/38sgjp+OvQRrFaEI/SUH
OnOFqI7CALPi+Rk2M3m9/nLn6AyITE3dNW2hvSVbUzbMsUfEesRX7f+Vf06w
8xuVj90GGcKTQr475UtVimN97AelkSIAWxyaW3OHoDAEUZQVF9rrVJxqnIWV
MhHzo3RhUlnsCZCsoQXGZNRWGxYyLb0lxiCrMaSr5X/ERbklfRTOtWcHuJpV
39wcSfucqOchW9ZJOEJ3+sEdKnMccMFXkzZukL88LYAlMuokC9W5l55s4uWV
S4qCsZePLg3w7bi9b4nBT3vbkus9XyEJnDXOSCW8NMEVAsyn1+x2nvD8RcZh
24j+cwQNMLWS4N4TdjVf2U03ycD4gVk0fKXg2K0LCvHopzJob/pRfsScR8XU
39MwbAMzssKdXm+qDkw1VA2yeI88zfEgNKOkwJw1t/QkKoaNRyOLuvu7Y4Aa
8ywpVRiyEgG3rpu6H4LQ8Hp7HeAGmpKt5ZSEQC6nOwavGe2vFB275Z8nYy+W
AAV2AkTGal08RtRijymmFE09dyKXj5nmGM0nHQzzm6OSHK6gEFtQq6HQh2yT
vktfQach57M4vdiMxvpc4IG4LQgLnNbYHnlbv+5JKagjdQIkuufCrxEVqPD5
GvCX+Dndx0ahRQzVHdm5dPhHEOmFvoDwTl9v8lSjQU5Sg+6SlTMMDBDUN97t
+PFAgZa9KyPARVMkfcAiMxo90tK6ljiwxWPrj7NLKAqRvW0FDAOMOwKcBXyG
SH8qW/WfMDLVtb8PeSEz4E63Zhq1R5sah/gWcnroZj4nBV0UZmS+7BhupOuq
KsqaCySW8Fy2rXn2hMuZq+tY2zawtSvGj7/abBvs4bSZcYcngbXVMolLbClL
Uy1WiO0GD9lgJgssw5FyIfqIQzxawGL2ER3bG7lA2KmdK+dHiQ/LAWeFpHjZ
6sEavasKd2435/KaUBL4GBPSHbv74mErrkuzdZQ8TJQ/YMw5kY9rMdnJ/a4O
VJIp9rn2m9wvfPwCRGBv9oOUte4gHA3S9nuSmJmLc99HDuyDImHBNRiiuMho
3a6lvgUDgqZQgtPklh4OsG+yEutmItT92eEJ2AdbWRfkhTeHEGQaXfjuYKwz
I6bduzYhb6BstTkHWZMEN+JKLir4Knhw8xbtrypGZSGGJ9vOqpgpgi0g07zl
ZgtIOnOHCsyXOeIPZz7HKGvHEPsI9OGPEvC3PU2IVu0WlVbwNYT108RokCoM
UApPceVMMlC5NP8Vi330xkkl1DCA74MEjaSDr9JKRcqXMm3herw9wfOv5hoz
gnr2wW7SQ5IyM3xR9oKx4yp0/ZxINB/CelpS+nIE3tgSKtRMsWGZx4jeT3Zr
MIfMaZ0bTc4jrmvZkI7bCx+5rSZqywbtwhLtsMtdiOowB+ET/Jot5YLA2mIP
oq6mgy2M/ofqMUJf+7I3E2F/vbztxJ+gRAOVH18hO87jszevSEgXjuDKGiO3
MnG42UhljZohcZe/h61ovq1cwFH43fmJplp5KLDy0CzrcjSnU63PXA1Xyuxq
tWAKDM+yDPyg3yPQsJ6jRz268M9SSa/SYVXgJLiaS9KbMlVdW4N51ybww2zc
PYrAyoZVL9qUC/dBgsMQ0/CToO1VIFUuCJwUiRzOIO/cvpOx62ldLQ6uNcg+
8NHedfx9uvr7qfCWtKh8cgMd/lKQEdZ9itnLQfO865snFTMgpkKxtGpslXZo
j6kRrAyJvccq/NyWT7HPM2BxJf5aBO9U0TWo5UU64cdH36Zh9wtGmLCXsYYV
qbgtEljZIDuuEosEueKu5+9fSmnGs5F+lzjTntlrjKJg/rcpQAvPi4JPzTxs
AKBi72LADR3lQzEuTn/Cfsy25ifQGQ0VutoX6DNWRS/0y37vnfYz6qLrGc0Y
LCXi9CgbLRBP6upD83CET3PE8S9IIrAU7gCcbiRIlxdJQn5JienEjtfjpLa1
Pm35gLlptqTNcGUMAtcWeaBqdIU3oKhDAK9wFWZakeik6jaDwB5i7I0yCLAt
YLm6eRQmg14uE34IMcYgYd/B8HLgTN4KjNZF1N6CrqZ3QOF00ULL5bu/MpOQ
WPqlVMMdJkcfWegrDP/Vy9i/beG7XcD7MAuwc9cggR7OQe/oX3IeiCApKbgy
ombwaKmpM335oSwEspupv06moG3RmjsZBytwU6cju40NYtiP2sS2JmxOgOGC
V/e68A1xZKyuwqdpOTInBBj0BcXuF7iYXRbnf+j5Gc6a5b6+Tcir1YZZVB7w
cNO1RlBdj3BgOgiR8RaCkDZIcH7dhxxMQguOWyGZ9k67kQMTAQYZOjqemtH7
bZ+TbvOOn5s3J0oBnKt062pHbr6w+vDiSc+V8SL3XyDMfJGIRxblKiYbUZOg
lJMN7PxuB9De3yOJc04aHS1msFykE5FpilRohmHYkTr/FUbpUYtsN61V9ZbE
NG3XSvyPd1Tk0xa0xBdYgxAQ7rUJE0HbdFt/KnnydgWs5/pKjHF5AHDZeWvu
I1nCFldEFdqIDp+/uL5TBTJcURjPjF21VuDqaUyHGORDBV124aVq/W2tld7/
DmIGjJJrflrUfUk4FeFaOAkoP6/9W1OT7Ylf6Kh33jerpTnIXq0tDDpplmU7
PCHJd/Nwad58M0AwIxByenCTR8b+0dQOP+Vz3BMQsYFrjBIO4hnhYAoQgRAL
zhhH2AJfGDWLP9qzxrEQEMYddQaO0GgVdCNvqys1c1T4esZDFOarp936kSAN
P8KtMrErnTR50X4fvH4bgchKjh5pA3le3ztFiv4nbpe0acCxGmDCis7Nfp3E
l9sHa/7NC+5cS6hYg0bcLdh5gw2ZcRtp8Lp0ebJDtGeXwXoRqeWQH55hdywZ
3lptf7zJUmPKyNO2CUSv8utSEW74GK59Mk8I6WEvl3cffJdo3utSj1yVGWKG
nAIfAFdgln/kJIViK5f0WWZIswMrDcdem2+zWnNmP3ZLVlQREKatUNKebHZZ
IjgAq6FfBBW73KLb51kC2NxAB3wmkaorRn5zqnVLNTOZ7EODzrTod8aE+rBz
q1fvt+lbJrJ/yicdywCEsQoAwWtWuzJQi68I1q4YzZr0T0VOMTIPVZHTkQOG
Ev39amTSg0Bhf3Wlr7hy+GdUbpFrh3y6Y8USvu+VVTGSrW+Rz2C2JVx6sGxx
Q4q5O2dooY2zcnHZxc3iTROAFx3cZbyau671eV+FzbKgqwWPdOm3qqlJ00o0
AuUvoufqRxCNmio0Hpqf1S9HoOcLWKnnjDMeKm6mJxYrp1UEyyLzJW6uILss
lalE5Yy23lanaYpa9ovX3fgPHwW68QpdGU6ZU0Iti4Huiz0ok5uehVhdBdaw
WC8u3QBhWSUSpo5Rm85irf0K0fv6iZMV72fkuxL8tJJIU6TybBuIuBFB/XMO
xvIT7cGlFeW41sqZuXmp1cI+xG0O/TufKH8vc2na/YE6oiuPhhIr7+HT1E8k
zHWbWxfZa8fFNg9xsp8OJAKS3cSnIOEFfutHlpjgW8Tnt/l8j6HxbMVgi846
VZq8kS5kHRfoUKRPXGPHh9tqq6sta3iDe6OpQP6PVVwLR588+FPSuzyjpuGe
YRqghIIuYu87ILqLKkqnmXwfjiQod0Hsiv+tIR1FNQl9CPIy8vMGyAre5PCV
VCMlYHdhWIS6LaH3+H2ryXAJXVQAzS9mzEVS0Ghu9o1ySbOzjIRcw5crF19J
oE8H4bK3tWCtNLwY8PdDhgePRLm4C+f7TDpb0ffdYJ+NAb2dRjl2IbAUxgcX
xBtBRU+TYAeVyLKXsHer6BB8QkIW6A1aUUvzZyRg3KhdXL+21przcCVUwe9U
M+ugMm1duE3TbStXw89cmUohAJHCafMnMW1uMOJflzuYxCFELfZKmHdfglmT
8GlBT+gVn926ZOxNQbApTpzmvV4ZXPfXfkdz/Oxg0nRu6zQUcoLWhsqMRDA7
eMbvEp6ma5Qi4l8JA0UoJJLgWh/cWrBTnLYiIXtWyD8JEsxmep3Yirq1yoRJ
xEVIT2NywsgDAqxdQ1DJ5T8GrjlDfwlZsTFQGjQhIWnDagWwMuRs8DZIfOts
dVPXDJ3drBkcw1H8w+Az3gTSNG0BO+jbPrlIpdBjd5pnl2WQeekjdKGqe1XY
ytm30Dj4b4Y/RuYrvJejHkSWmlYWdEYY47pMzZytg1okPxTnUOjXGHhWNUkO
pJMEUnmGgQa2Hez1ek1izz5EtSzKN4uUxEoztv8ROJnSYlwh5xA9v1+uLqh6
POcagOZ7jaLmb7AOUsGcGC/OIYaOAJ2hv1PgfWbp/K4vEGUOoYvOtcG7Iom1
PWZ2yviEzmbleY5hJqRv1EeZRhYCKzT0G5K/Sf7xjYnoUfrtHklurAgyYdWE
G5xZ9hB7eCmRs4laLbhkAfyXOFTSDVANRtkbpLHuF5/wHCPeX76kFl1HRGMH
4xIoEEFkiIdMkVhKRJJLZeOBZeUbQ+ejo9I6tGtzZmH50gPMjnrqHq4h1vUT
MdSw5i7kAiKLL2Tmg5nLkKu5q95PxvzCw6YzFkhAiYneW/Cug83SbaARsNem
OPnhvlQa8RZW6UQR2sOfHSq6JSNwlc0PbkLPMcqXO32fUnIG9YeUZpzNamuh
bZSg05BE1qBQFc6oWRC5VIn+DM0cfF+1gWFrZNCoFMpyeE7iOTpkoS2Grojc
oHIkRjGAChFWNFCRTQ7geRqYy+6NAdHk0p/sy7cxBAQcKYqzhGge2JnJ4Lxf
J72d2EUFLZW7yur7IwPDCMC5nQWW+4LEJliwhvpxSMYxs6MfArW3x39McOqa
QS5eGEMFgSW3Z7qD7rmRDeMCaqjW+YAWcKBz1QbtexbksRxqGUjNPGSEaO/n
vA8zVZymNVxChVX7IvhNIveFO3b/njuDJBvY627XMy3+0k92kG7rTqRSGKNm
iEPdausaM1A4CFe2iZTIdP2mOe58bbv8SrI09FUqDzDHaYa7/x0HZE3xSu+7
V/q4xPrjgPIIIKlU4NZlfAFaVZdnlZ/257c/3DRcgFHH3h5moJffHQNzXTDk
DFBVOtaSoR/V740voS7gBr5Lj+cpJi4v9E0sZFnfKeLuUH+y+ZotjT8ebPCJ
Of9RZCVcBT6Nzm+rFSyJcjJmKL+eYGpdSGc4tc0O9KEiuGJdwzCstksUxcT1
OLpCOLsi7kvBkBjgGb7GGqoIpUiRNQumX0Pc0vFMo3LNtzNcm3YeKp0IFCh8
llzec9tdpLsfEGVGLY63FNxLEkYB0c0z/E7XvPjvfOioGGfTimGPUhE5Qh5+
2oGKUUuUCWJY3pK9kwOzgYRBzzjD3UhMup4wdphrhVVeBtG0q6OkoQXFZ0LW
BAX/TC0WpxHnSZasXxqz+tDoDqfBLmRjJvmVLAVXt9V5CQFa64wXd1Hpv92P
we9lNfWlj7SyToEK5ODBBsJX4bJA2q+rk5DD04pDh4XZ7YYGdIC2wuZh2r41
31MJPCHeUwAWOCee9kh3gsP6sWNSOMtdD8bkYJ21SNWFYicRBbhhRU8G6CoG
fvzh0DhBDOajPtGr1lpuE1ryNnBquE2K8exbBQ1y0tSj158jjeW/E/hfCdcx
lsLDI8Vbzc7woOLKj7F/3SPG8B7jZO8GwMNXT1+bASxbuBdJxnP5UO+J4rci
OVcWFjxCXDr7gHMWqjRiWDVPX0Qr2r/LafOJr50twf5/bqxbfoJsj2kJyXtf
YhNlHflI44XDH0P2NzaoIKtV0G9eymsrpTfZT8x5ZSzkQrkAg4Kx8c7ZrBuI
5x5d3Er6yX2npydQsDf/qoLyscUT2zIOvHof2hag/7C8ZEnc8Xg/VKaqQA0t
Xzq4TBzQIPL9w7yRzGyTSn/GgcqMdCaUyWoo4V5aZRQqZ6k/tELIIx1HH1k6
66Rf00O5i8wVAQVuVMz68+FKM/4D30eHamLZtQRnDgJKt5ttd6fUAjwrdsJa
2KHGQc08qeEUHlIFMTKa3eBGxXbYfYpjULoNMh2UwmBFFOBvWIG8AGCGd4Zz
SuLHLdeavYg4dY5f0uunEEKQne12inQtdAVU56gomwjDS2IA8ww1FvpIkjyD
OB72kAIU/uRtBk6bX4AZmuYfj8UD1vRoxOSnWelBPM7ZZgGIOgkYQv7QYCf7
yKoxyCvWjdIDxQpy2TLaxtLBoViYkbhnBHVUXB4tIABTxioxaqYBbUi8XKOn
aFiMH/bhuPS2Fv8jE5skkVlBN9ozWhk6P303S3ewhoP19EzpMgpMoL6QZKzm
0V6KTFwdF+4vJGjujKYIQHPJR0zAI5QQm5m8Sviy44e9i5+K3OD+mqtvyioR
1NqsR0TjXp5276lPY6HWoO7Al3Nm3+pOwKWIjGvD2WiMbzKjkumdfgXRBb7v
KzSkZuks3xMGYjWa8bApJODhOcyZdiJCRrLgB9pOZUUa2Adi1NzDH7K2Qk5j
ii3nDNi2g3+D6iQVAsP4ajKWfTPoz1C7HGl/kkaiQRhstXzemOletTq2M0kl
JaS7iFI2NNyIj+ZWKjxnnO7xarav8fDQan3Zd0hL7Wt2X0e9t+t5nEKrW8vl
slMV0PbUTR4Rn17kXbKQsNZvGyZrftVii1AImxcGDN3vs5hP6F7UFH6hXV/y
0fH1yuIM9IBHy5libPVVz9BS1Ohy4aFaR4mxTNt5xOwgNwD6mbJeo3AMCaG4
a6+wFA2pLla96Ec35OfYXoAuok0gpYcHnjoNuDbvIIkYh00Qh6wPHAqmkrx1
bDRYIYGj/E56JGn15tp19ZEseix3kvGFsQ3JnnZ9Dr+YvxBs1tH9u2OGznRX
3KUkRJCnz4lGv5/JElnpaJB7rv7OHa2JA6OLFs3gns8gvZ5ID2G9zqtgA6Cy
l1BFuyVbyZSIPS6+5VsEVQ9VtKBj39NjyXE/Z/8j6Flcj28WM8Pf70jmGyF+
UStbamqHFi2qzTU31DWOC4BO17eAEm5q4Fr26F/ZunLc1nAS+WH8Xnr4EOK2
OA57mMYo3xwoY9OwTzQzt0+Y9hOPLBHI7bMCd2/mXbt1xcSbzloPimES6wNV
iQq7Z/aVR9ZY2vHH1jAXIxEtMuUyN25xPupbQ1t85IAxoA43I9aL0488UHpO
DaiD2K3re9mI7jtw/YqaJ/jJySi5QWaZrZ8fOMLsoOT954/2JhFbBWg3gX5s
oXgp9XHD0XzIsluwM0SctbuAycVt+oGH2ye+VDxIbjSra1p9e9FRCDDbOJfV
GwbXJmXi09FXV4QOHCQKfqj7NIYI2PKdAorgT1btaePVgALGv8EmmGhXTGBX
dO5FEG6gVifc0ikr+PmiQs3LFzcn84uMSUBrE4uIiQqZXflR3SK4nQzT6ukX
otnXHmP1W7F4SWpLft/2PgZyHCWswDhX0RFcwE691UQ4CLXovLah0NNaP4no
0pWF6WnH8gAzQEKFiKykfsWKn1wAuWCgdE4FUbEul2sgbqZMkeI/+6VZMa+l
iLD44ZLXxHUCAZNIJujc0h76LsIAVpK3YMHd9izYVf5NyaREoJJ+4l47mcfp
mu0H9OUaAVu3Ee9shP0uUoweMqvTKrfMNbSVxQFIaaLtoH1wo0QlzvuCaWjk
hciJWW0G+MrIOh63HBVLIxt7b1zCxXqY5BuaiDpu6It7DlpuCN/qWx1Uviy0
qO73hxMhEkS/iPLkFy5WbZsD3wp228JvoU1JczONpQqajWKzoJGOnKTO7GZe
1eAVqj4boPchvKuTga/CSGh2AnAk64ldnnq2aMn13J7QgZioR6Y2Tgiw/7V5
m4YbQGi5SRM+N43FzmQ33bHo/gu1+XqtubNJki1sMH8ClHZ0HqMfKAYSw0lT
jPjYlUGDvTeg0g71H+VgEyUM7O1Ye11X1znMbpnStV3thjxL9nmTVTbpU+G8
gaJfTLFJrQsQic2Fssrcyhp2DFeuZL1xVhS9FaR3W4SN2qIBcabZ0vRmv8tE
M8q8K5miWy/iMsKSGnLndrSc4em++aIh7LXQgCCrnpCAiCzcJzi4qLEDmO+T
BQ/gL9O6wxq0EWXwtwPtJ6K97Ld846lm9CopN1KL6JHAFx19UpiWewETgfWo
CCUoC9MhEN8dZTXzrXHqTy5csSQgtLO/clbUmAaXeEPkWJW/61cCvwQn313Z
q/sD3W+HBfJb5NsNcdu6fUqHr1d81EC8aXNY7aRlE9ceH7tcDbjru8fJYNNF
v2Rp0wi6NCavBzJWrZJWgaUx9tBIQEXbE4J1rMRBlsywZIn+3iNHSgwaGMY1
4pEGe3ZWh6/809Ft/WmC6E2j5Ba2Y7rFI70V0knrTKwLxg1V9ZYQIqcyhV3t
4fY7JjN3VW30haGvYsOSKxXoJG+sLcmM+9Di1bMP26Mx5LFGp4TNYdNjAhSb
xHIs6bToXbKrmVqudzUhSSDFM8vWogdE4zMJYli6za+Er1NzrM1vFacIMVDy
Jfv+Zxr1zr5fcnHmyTP18ziAgEWbbkEv+4aPyG5WECbO/ZqcCVVyukOP7cy6
AdH9wjsdk9Xp9Utfr0oxpQffWDA+nXUQfpOqKw5tYnJM/Wr5XyfV/VmE7RES
SKSfxzLPYpyxS1LgQbBTTGZ/zIlm3Y698QjKFGnigIQuJVe/z8I0yKdpTa0p
3ykMWtzEi414lNOu3ULcsvy/xGmpdUzbulijLRVtBdgMgM0K1Chwi2edSqPf
Wj7Zm8MHKX4XZha6E9Ec+6HLm9PIegKlUuUaX8tyPtLd1O/Fy09vkO6hzI9F
wrTwwT6MMjIaSn2nXTcDnH8VSv2kTrvfdaVmiQbEsbfiNPVvvhzPjbC0NVRn
REY7m4PZngA0Q9efy/aTE7xHGC8nQAQf9WMHT4enocQ/xRtm36OvHLrOKTKa
znNXt7tUULhVZI0rZs3/iEzWR9o90hH4xcBZGpRk4xPzgA707Fwv1bv9aOvn
+l8BgorO9mqVFX+9BT3ytkfPQoY5xqnDRslJtFcA927rXHiqMv126L9ujB7p
aor+gsUmCvfXZJLefUWPZeQyykPLceZmqNHTAFV8igmPqjE7TZmo4fxZgiOs
rrGKp47CCl+VMIZ/9yrZJE5W2i3AM7OayuR4K3U65BYzg1TtAkbGxbGbUpZj
VIWtvZ1Z0G6y/bRJQFU9btD9mQdTiKxKwwzcnlV3Bd8ejbcUeRcguqUtaol1
UA1ure34/aBRZx3yXMgevuxEzQItytD5GPWsEs7JZBe1kJerm/95dIMVmRof
xnrco/igqgImQwyZOi05QjQDrbNkREcpGCFUs0DrM2dDpmBkpD+OTtg4VHUT
6IqXF62b8v4x4VJhllgViRI7IfoI00XFoe/f3eJXuBERtsTUxSxSQI56q+vt
sOH8a6rPljuoKWTst73sM4mY5Ypr3vmQDLwa7TgNpkACwDb2m0vaLhtPL/L6
ycJFE3lOfGHJY0EBX2MeyvcRcXN7kdAi5jRmIDdoWaN8+oJGTv5nkV/X4deG
Lch7GU7NCCxTT5DRbENfLGZcgirWA0cBFxbdfrpbbRXx2bOH2HaoShMBr2I3
b2jKU8FdUkcjqxTM5xQULmKWoGQgJfwK5pbSgGMf1v409CTTP/dwCV5cWqBW
iKLPlBtCjm+4MvHC8aHIUq/kc4T0zU7YwqdYw2cx3PHJtVIBg5vSGGWbDbQv
ZPim8rMJ79xemtB6mPTXnI/lj0PdMK2bFnAqIbXqeBnVQr3wVnJAmiCcmo/5
8HPjWiNfLkaje1S1NdQq+nzbew9OWQwpZjn2iRl4z++X5XYYqQZnymjwAEbu
/xJ8VlGSwTB1AfWglj+5uKcI5G7rQSOLSCS/9MgGinuqYcF4xtTO058RGOZF
RlCqSBQsDP7P1JyUehOUn/fIhbgzlrSs2eWbWkP8e6xSWCEj+Q15B3RvlweQ
GnTwCmmm8Jpsm0nJLwutsozzgxn2feeMKNRf9fUOLa9uwmK3gfRe+Z6Wk3ph
U7SHKn7N0bRTrA3HbZiDnsj3HcNY1+ctLvKVA294VstB48eRvlIzcDxp5IrZ
GvkydVOPhfl7EH327146xHNWwxiIZAtwqFcRUBb73X8EADuWBjdk6j+vbUFb
Z/6btFJrT/QpN+HjwQM6F1HPKnseaBrG6gPHCEYyMnJunjVb2QxMlN5vJb0f
GikklGe9H2ofd9fAM+UZfkra/5OxE2Vo2h3UuvA9GudhGsWNSJjeNkCRxfBT
eyVlZyUceb/fjoXSIDnjaImbWzUPqtmrE1dSGivCqsfIIplJ7hHtcfVCA1HL
XGpB2tWT1SBjAxunj8Snqvg7I1dOkA/ZUPyFN12B7pA5oQCSt3lvcZltRY9l
YEjwk0fZVnIJgAM0tpY48T0xt6HcjPZvxBD/i1tVQwCO8GK+MNQskkpto0t8
bl2inrRn5ovqMCP45w0ZmKIi2ehu/5WwtTZPWNiSe9n3d78kga1qHyXM/6tr
p2hyyXd8WiupkV6//qErMfUoaWPZgFmQaIVe8/WpbOmN0AkQ3rtw3sri3fT9
buG1BtiUsIlnITpD6mYrUj/WC0fwwq+UkJ+N5DCk9U+OVQkgff4lWAUMoBnO
Kdy3yCZdq/REINDFf4vdy4JqqbzpIAgUlxJhRvWHVulwSmK5/hK2WzfQYxSI
LgHLKZk4V++5bgvTIKSnKQg4O0yrZREy3cAC+E2734zz0FMoWSNb4uskEsjy
OKJkpli0jp6vwjriTRZSXlQO+3CCjJ1ajqMAOuO/O24zfswOgP7v+vHHe4hy
T9s4T9W7uSjLqnjFxo/hpkpBt3CrcqCmjYRW4k7DBsJ2E38qp3xNUAv7NuzM
Zy2mzaX2I2TtjaoiRZ8ixNwX9IvYGv/arZN641+/peAzZ9NnmPyA26FYAPpw
UUcWGXW+RyUA8CeOohrgEM+H4zW4mPgWIrG2W5TmC71PxMWPt4STyZsqIE9e
BtJWOISJAbgVQe1dYmBLPY17AWgyNLH0Hnr/wvIuB/N+eFcpaFgISs0s4RAN
UzD8O83xU8bphw8bZA9E4ZfpsPEYYUZUM6/c6emDwWdjhincUSdNpxviumG6
KWGkNYjdWcUuFQpl744pXQCcMza7jku5wcY68PIbxTlKJwyVXs+TZbvt3Iqf
BT2eEIoHRzN8xDXdQM7v6lbJVVKBsGJ8D8vflJvyTwVSGx3lU7hxINCWk8vY
q8iqqbt9MlCGto3Dyf4Ix41dZc5phYgUcGRGekYiWP8i++zmoS37DKVRzPCg
TaTnOGDhsgMmtHsZXNtCpN+vWQUPuuIwWEYCoaMYHkNnMcHuXsjT8QMdgWql
7B4pZCnmPRDIp3B8HIISUgJr0jM2SZSrZGCm6M+1TbwXwlKynOjAtpjvBPUk
B2AaHlNb5+ablCFaWRmdqWHAUkUpriFo3VMk852S7uhn+v9XpT39cMoFEB1k
QNuoSSO+axpS8QWRC55pPeamYAIviwa5ldkRdLuiY301YLskwEQyUY2cCYMz
hyaKQyIjcl9+r25kcuRdMpGFkWkKoI4DYy2rwTBbGREZ11xm0CFzKJc/KmRv
FyGrxusvGcxcRRhhH9kHBJLZy6wroCaZqRSqhhez3IFnvaAbJIW2Du2BiD4f
/9GUo3h7/xMKtX13+YNIp2Gz+k8p5/LKU6JQvYISBAtm9umRzY5awk9QKxCE
UDwaooA4zKtUzt9872BNRki3LC6zY0BQwU7Isq9nPci+sdRJTWVjgbnvqmUF
PNsCyYKnnQ4AedI+ydj3Ajl+8CBuZf3K///U6cXnGOKRmvrMiTvs4JxsuiJp
S1cOqi0Zv6RkwczljxkEe2vUTg2D1kt5r7UzX9AcXq8vwMFEps88/KEUnnJ2
X10nccN8L8rnMboNK3Fw5HvF4nkS7kq3YChTjEQ6GDs8lotFy4C83Ox8nGCZ
4XytheAv3wq07QavP8GD3dc1fCXd7r5+5CKwhc4pK/7EOnMihURV8DFO6oGt
sdoEl3eFQXfS4F0OCuyD/KAog/zCG5IA/ZmNXp9toCbDJ+PIwADNeWqqoUgo
HXIUdxOQl4LL1Qwjl820hlamFz/kIpzctukjuaBthXtl1cz+tACVYqRBklj3
UoCquVsZxkgOhzbG57hPZaBi458ItE2uzQTC9FqRa6XeGikzZaVkDjZYf9FF
uh7XmROlojocEG0GdO9VnDdElvKAQrruYZnL41tPKFy0uJOP/fr5PqNN2I1p
h7cbeXo3enXWmrMk+ST511pQTxFc41B+5QyhDDdOAMALGZULN2TbBjzrPcaa
W+bH4rWYzquNrafo/RYKKVFSg9Btg/3zb15MTGAC7fTwvqpjN4KPEP5zCm/Q
IOrQDAJ0ybcax340CFkoWKSDDKtDutDNkgr2I0DXXOOP4Ls1srIIm0O4e9U1
pnpTnktXW6iwd4Fm/354ADpfdTfHuQ+J9uB4iYtIhH9/GmvwEfbezYeavPL0
PKqofoxB4hcy2Q2Oim3H7H3U4WBn4yzK6ds/amRNII7tYEai6Vw79pNyd2Q6
fAGnBlZCZ4A/EZxoTl5r2Hii4JD5TzeotDm0tjwo7RPQsoNmgy7oq8mgKBtK
wzwWit9C0XTrzSIKImMp6MgbOqF+UvQ8Z1Ls2jDV7584PUFmp7XoLom0YcNa
33g+WYCsO8haEZlwelVlaQeVXrfu2XMzuTnxi2hkW5PrC3+uB7qIwFlPml9h
yaoBhmHWm//wCLl6PUuj6NZlSKdBZXM605xgrSwT+UF7SY+nkXJnksRcRACE
vISsa5i+0Nsi2SwYad9E8xY85o6pQlk0B4WYjagaYEXXPk2IDeXmqC1lrtIs
WRlAnT90Sf+5Tb0/5iZwe3u+fn79anh+2Q+TKM5AkBUh0Iv9uy7n4nPqwHvr
Fnagm/miccmVER5MtmTN5aIkAT5EOiauB5uWhmNrFTdenLo178l0Y5x3jXj9
Gtxl/o7KHhF0YLXCHHN9/Lyt5Vpkp8K5UlzY1Hgc7u/+L021zI5l5usu52sb
3lqHk/fQGy3iYXAHTyZCVZl1wJ40525Ovho7n611k4NddyFlwoQ94jtiEipn
oAvVaJEACZpOVB2jXDTe7cm8zjnkTrCqQmJVS0vNEqqQu8xBDU8f/41rvk1h
JkgEmfh4PZInEXiFAMoMl7/WHcduwUK0n+Dy/51oKmF30ILhit32fdFI/nS3
CeMpk4NjfnKp+IN6AX9ogeppAxdJAcmFaO3P985VQuOqXWuO14HlujLWK343
+dCKkYiL5TOpy8jvAzaF7nsR8GFR3RIXBBTE+2tB7URiizDM3sJwGXoTY7iQ
fOfCp8T0RYVXs1wjylclN724LPL/H9CFBt61wH9OJh/9HokpwZfHTBEXUwnv
iUOX363C0xcIyb2LHxJy2EDu9rcdx1Gmb3Aqc1p+jkeP7xXvKK5tSd/yuALO
URdU+3hdPMt10EHkzCWRBWfxopp2AoL06aP38/9XNDIXwN7StTkWfiHOrPX/
s+kJqSXvmCPLI0zJeHT+8fDaPWzEx9BghEr6p/Ndl996Aa8XgfUx1onPxm1S
jgW7t1m79RsgdXhsZqFpmcMFoEJTRqt1ZPcyHIbzAtnndXEDp+zmawaC710+
OHbjc75ayuemnLbqTE+BmSLHcqyQOxQSJp74AcE4XTWqsjMyNc74ELa+Zda7
FLn8Cgm4CPlM26RNIckLejoQ18WlQbFzMFMedVN82jd8N593RTH2jImeKj+j
2H/YT1YWeofOMtC6CDz0dHDaCO3bT3kgf+qhocb8yrAVvMVqlDmgkzGaheYF
istts1UNmhpgfDQJONLjr8BS/DXHduG+nm5fWpW45v3iFt5FzMUlzMiyvJql
jGXf3f7Vdx1Y5oMewKuutv7jbI2Y5IK9ksHGHsXMRI3DzNH61UbsveKhx8qe
R+/q4j0Y4xREkfR5n53BMzai/mqoHa8eEUs5fC0lPvKPm0Y+FG2dR5u2IPU0
9LlZtVVgTrzFueyW99rrttdHeGUrlVPdAzRO+/XShlwdt2VsyjXrX3yKfnS9
PT3l9Hftq2cLd/eINrLvM1QOaUo4IaaadOA02wQ29ed5inGFZb+DQC+fPTqn
gIWZPfWwbePT13Yp6PeSHf0sNwlF24OFsgomQ6XH3Qq5WUQ6QX+PQdhwmaAL
XOsBO7sxV/pTvi0YE3Z6m2XeZn3KI4eAEA/X11jjn3R3uiRKd+iyNPOeeJEQ
qbWFCiS9alnUxbwndMt6dhrpBoOAeIuyJLyKoX8fKhJhQYqFb0rzUh2SRBb6
rzhyZIgrTW0nh5pMaAOQ/3GrOo4fqttMbe4gIwyVmaVUzxNYrYMMuSawIOj4
HPeIV0mkoMoWdpFVdMrI0yMROZJUd8EftMiiEct9KVjYBqsXMEzBb2I5Hccj
f2awwm9AvchIfK9wJhVB1+9nxswBxt1g6tmOdSBcX4unZM2o1oZTc53OpNRr
9fUHLe7RysWp5mKHKDVMc5pVZAYyb62nb9Vm4xgHo0CzwjzIcEdEf3OWpPFb
j0MUtJ57+CLbZlErEMGXQVhMKzKfxNHxN4osotU8Tld/zSWhgRV6pqcOz2bX
BDAVIa16j8jaCn+otmpm6rI4WbUx65Cyqd4vtcO06G4GTa2ZHm0xwGdYiR4V
jICMFsaaxm1nh54Tirgx/j7nbkDTdDHxoRGGCO/KikUsRWMpVjQK3zFfley1
2rgkFh3/nGiA0cTR4Vinu/HahBPB+b0QVIVfC6jXM7i76w5zi4ns+f+H/SAw
XduDTQV0/hnPBC0KwQ0adQPpepiYDvcr3yLS+FmsrNGqPoB4OI/ryjDv/Txp
lCoiv+C1WgtcmJYMmFG1TBBQ/rrkJF603osJZltcd4h025IovY9dOIGrTi2S
paMhilUkLZPZln4Tht43poMEQuNGkUIpEWGcHdV9tSK7FTNr7b4NsJSUP+qg
M3o3uFR2XPNB/yBCL4/64dMDJ03jj1YJaOGAZegVkVCwQVUKYkOnoUYuewL1
DAU0DeDcOD8PpW0I/5Ssi9I0vomLbuybfmI1pA88d6kmANZ1ZgLfk+ad09uS
25+YkXvXYr2XkiV5cq5j1Vwj2Nryzr/SS5VGc0oiexSPmduTGK3CiaomAFQb
0sn8g3YbeQjeSl5n32LNyF4w8QcVMpElMJ+/j6lEYfG7MYezgbnAmrO557ll
mcRpQB1HP7eojwfgS8DvvOq+XkkjlllmBQsilIdxVgUVdhg+beJoIcy0W2EZ
jGtsxkUarsX5P74TeCeD/a50EybZjlYwSQnOjmd69c1zs7J0i6sozN6dHw/1
F3WkYsMA+0Xe0zVrIVT2eaPztrY2+JuK3pSyefwkEl3e6eCHg5kcgdoVDq7A
ovp6Ka4FKSdyjYXQ/mr4Gxp8Bw+RbtNmMMR6LqthSMTy3NO4LkzeS/Fo2Og+
jR+32e3MKsJzVZJDn+2iqdUIZ8uvuiCRmo6Dj63lj2GR1rENnbl+8iFTrJ0N
h30EvjANqKkH1v+bo1xjxbat9POtrk3e/1ntp5G7dOnQZ+9wK5VU4GzD2r2a
LqadMPW4VW1UM17eL7ba7xwIVYdpeO9GCGIY1FQhJn0HOoWc1UxPLehCtqhn
kzpIu5wRgR8u8E7uirWsAja/IH/Dyndn+89bgp56a9jA/o9RJHKQLtgK0ld0
1rVH6Pcz/NVpzKAp+/eBQCCiNJRLbYCdpzT2gZ+dXxXllRIkE2p85dL9nh9q
aFssa9s7bUXAk5StxZqJTab39qxBoR5HaSByR7G1faoPKIGlM94N9+j12yOk
QjWk/kEZ5QgJj26TWy96Hqu7KMmNEzOmFMecOyTUX2iRKJwuUV3rLE3dTUl5
fo/uwMNyqytxojHqkhNr9VWds/FQzV0zJvoPIzXlAr28p1TjvfBoPONTFoPB
ZPRbF3pekfu+4/REOQPGhMBoUyKlhI8RTQVWAu8L7LkoGApuEHYpPmCmEpzJ
umg2kk4ytawF2IQ/c493Kj1wCyOQvt/thSwKS6J2HTKbdGjuioafyUOkpln+
iVMqWRziTK2Ro0NX7+Jk/L9+SZqJ9bszokzW4hQeLHD6PYgpf98d6oOfC68n
vNKfagPNIDhR8nPHTgTpwLwRXzYTlDaquP6Qmz0KXxUFwMGNS71dfnARJM8/
g+MsDQfK1homwI4KXE0tmiwtR0tAkmUoLU9AND3h3eNdeZQQAq17LTgXlZWE
ykd2qhgy+rM9s/UZAxcwyyX7roWRpxvsF1kJJ8l/q3KrZVWVf1nDizstcWTn
95/toUMboYxpszFIZEOltkHLn3bVC39UNTkNQw0CMYiyZGyqqQYFNoH2cncb
NxwxDf01FA6iWtRclZ8CqA6Dpwz1qK7q5QnXWksetVTvcOMMJMCv3mX8tmOh
9agvHeiiinvK+KYd8RbTxxc4jySMxAi6n99bfz0Y6B5yf5X673G7tpsiWWC+
bBer+wRwnbVFtU1CrPSesLbwA4XD8dNeZhe66DSQUxlRkUMKbX+WXZ6mX5BA
HghlD+ZTMK2TFz90xqRw0eO6QBa33qHwQHiV7iYyL3j1lFqMPW/oD+PH3QGQ
7Qmb3Ltvm0GPOoqLtmkEpkRDeEYhO+40prRjOEIYoDyv4jA+ZnOPO1e+Az0y
xu/y2omugibo+4LlXv7u9e9panjYkFJyBmeY2DyfW+y7/JHNnP4zsEz84/cj
IVmkSnUd/NgkW5DsEcC1BX1AtyH/g5TBcIW6c3dw+XsmVMGtm/mhJFvParYo
lbDNbRKUDeOi/suRwAULKi5SRHaQIhP1VX1NZwKTFJv1AHHoK9uUMcdn8IGR
A7QZREIyOSrr4ah803yBXivEC+BTQgLyDIqSla7qjlu4qjLQlamEXhvRAPrT
WEyBYwXGNONsZnmOFsbkOVlIrAK/1ImuBM1c8ZplF5UUGbgrx14oGz0kMt0I
2vkk7b+JdAVbMmVizYZCeFEMXzXf2VTgXG+z92WJO4idl1lpZuzTX80qOsle
IeN8yHyFPfIgUvB8teMoXOtY6z8GUXymlmtQglP5Z5I2QNHF85aeEYD51vmB
qtGo9enoIYDK9GvaqfHf2GUguKnyYGr4M8pOz/sSWzk5HZ0OkOUwmQpbEgoA
q/fpZ8vOvT3bVrKnFAHZ6agBir4P48INEpUoNZn0NyMHZGHkREv1AcsDpjv7
zWCxe7uSmfaa95YGeTfefuduLqyq1ElaS2BvW14L/ESwKhzH61XRxuynAcId
Bl/qFANHoz8cOMhnOCA774k8QJC61hvCqmB9lfrH1mqtEC5PrCHq+5yFWz4K
MBy2XilFpitOD/eUlB44LhCqQsNF68vOsvjLedH7j4WicXmwpnxhn5DEo95W
9imt51736uivEDQVaQGU2E8+CsSRsWTe323KPAXJS8OZUSxUoaam2xZZ+wyP
raXJMj7G7aNYnKjeaIlcSyHEetiGQULDlqGLEF9OFH113sbIsvIHUp244cFK
4Kp910soKnIqgLobSauCS3glQF/5nRSfVDjksJ3k0ordyD8ceFZR5LL0LzpJ
BRUA+kjtPZug0QSFrZbWREFEDKRmRRCG2yj57NNMY0zi3XBHNFzQJSlfdq20
0eL+CULCQmubzvJWQZAHjnrGaieoUCeuk5Am3goVaptahnCXi/vZh4WKv5v7
QXn7jzdR8y2bqkQap7DYccpt6bqBONP45SvoXTqHezkqQMNhNZLDMGtV2CSZ
L5J8VBM57DT1yMhws4gLyzGFSPb3RQ1KJku4qYaGh43G57Nx8QnjiDP/1/ij
VqwT4M2LZrNNCEjXgRwgtSlg78EzQudrd8z4ALvCyVAN4Do3S0h7nv6ERNEj
iMMbzSDvxeVGsfL4/d9iPmML2hWWydRNk8IZlTAoCM6tI+DJ6FIKWv/PeSL5
Z0zcW5Fpn/NSsq7wPsWnYFVUb50v7UZBOCAUFQ4frvwr/uV7DP1wlL5Le/zF
m3A2/YneKsx2ejPtBRcSswQMPQLBjOAvkY4YZtvfpi+G1sbtTIQ9X1r4vh86
IX7nNc3qAOPDK1N4cM6G3L/QRrdyKb4wJhBQF/zo1trGXCTqMtKXSb5C7PgV
1BscEXGnqaQSDDrerrpkX3A79NLlQboTh6IAOZzTLNunEGaSb/jmXqV8LF3v
yJAPtLfEVKA3xCYCve86DuJncRTx9DCMwtzOnZZ7Z1OEAdK4zMAa/827im95
ld5URsvdoo2oxhscujxSGOPJizhLZogwt6cofPHlOR7vZWlRRZ2LWSH9Kr0U
VSPnhjg07SAGAeP5w469RIOMIFlmdrOGMRerr+qKRcqjyN1uma5l/akfCU/1
6tU+s3FVf976+nOdguczjmn0dJu0LcoMYZvo5OW9ZxB6RAr1qkMTCL4DKWHO
kCirEBthHGvKl+Zu2ZYMH208TuOZAIE9V6l4bu8CiGFTDRfjlx0t+lvDSeh2
5EYAMWQXqjZK2DmLxGhvVFFctX0jfOIFUqzwBxMNhwjtfTM3rUNA+zLuLxvB
xoLfFZHAhBb7zl1qt0KuLAH8elC423rveaNhjHbLn0lQPXmulgTgxiXIh1iI
Kz9Rewavqmq1qx2xRnNvktCtN6ySoNFP+8I1D649JSxpJ9I2b2gZ1aXJosjZ
sRdfqShOAw1Os99ifi8M+x1ptsVkdXzGxV6fqvk7EPmN/HgEq2JNZaBOkSAk
+g4ITy6yOJgshcc4vsfP46IQsmT/B2KpYbaRL4u3HagpNZ7tsuhca39Wzosq
gLC+PYf7227PQEsITehxc2Inz0OlChxDRrsIHaNUr+mm/nEvoy7FtGpUPJv3
/FwVIho6uT+LiYskhtQlqIQe86Msf3wWnCkSiWHHFlicVSE5T24buiwYdEXC
mR0aulc9nnQ1+lFkYMgmh6kZoWOCong/W2R2nYGX0QnGbAMWyV6OQ7F/Zrtj
r79TkDTrAHPKlzpwp+Y7VvzZhNp1RAX680vojWbAjBjZ1/UAhfqE8zh6y79I
TxFRdVzb88+2JV1Yuip4YltXqeby0bFKlf6Fzk5yuRazdvzs/71I80MtaXvy
0xCG0ZmJ5Qxrarr9Gn5DFO/BPm6IK0QzVYbUEMHk8zbssIh1kQigWYIGkj/T
yy50BDGuU73ctDdzE4f/YvxWqxkzVH8vG3piElyqCTVSMWIYcL0povcAdbdp
bw5vpy5XInuS5fmx5wpRaiIEWu1fQDE0g7pI8tDGpt1tibztWbpBcE/BpW8g
66hrdKNo+ln0BbDXOJvhqId/6pgCrsNeHxJMhtmvYaQyCxaJARnPat6pC9kd
UYaRWvoRqDgWTddf5jEA+tncH4RlMxhY5JpIK/rCn9mC1Ba0+olSXrSxJFoM
Snvrc0O0scr4rPN7fla61Oz9zYQ7tuUfMoLzxqUfxj88JvzHpt7xL8qcnnCt
+ICrqij5BMUbKBPhy2voXLE0lgncPNcLuQxMHOks666KM06qCJN3LmRG+22F
EUQxb1u7aWFzovxRbY5tbt/ZS82Lpix54GQVyfQqJh6hVDVWWe3mPRCIu/jR
l24pxNjXFlc73+PR7VnqYnzFONiEzI/HM3K62xfQlKGZ8vq1KTKikMU2yqMQ
CuPHy4WhuHiRDofR6YspfMqN16PHdT4eJ9j556L1FzOa8UE+CmHJWgc55SxE
AG8rNWbdUdIht9r8ng4UkorcR5Xj89Q9Egm/NflLEqgS895eDOCfIFOBxzDr
07O2HvmmG590AcDqvMSSlDeeBLatmdHEjcVXC9PvF+BDfSA9CoXJVWCidhJi
Xss0f5fXyHkqT7pRJzH7X1FEX0ycYXs1ce0j50jPmGRWwxYygEB9l+m0fOJi
uxpDUinummxn5RJUPk9wlHF7ZlD8y4MN19A0pVH9+tolj+GK1hzxVDirV5l3
QFAf4Uq5z+zpxmCN5rO+/RBAvKDC0j0hIEoNfQUls3SSAlqsqrqWF51cpMlZ
kZOagI+wpjTJ6Y+tlsC32WuKouXMOjq5dq0n5nkvnPlGzekhQqdOfwl+Ec7e
oJy8gDtNNK833pt9XnoyuRZbglDKPyhgrWG6lZDY/xddX01KBVC1Q8nOI+2e
VHk+SfJ+gBsupY4GT44d9K6uzAbrXUK2ILigr1k3OBQjWGw/c3wU3Je/X766
++kyeGLjWREAmOoZ23cc31s3ykrzTvQf1FCo021TczHaYfDZqk4s/cmJWhYG
AX/7dHowQmAl2fEEinqHJ9hlMlraCtbaEJSwB1hZL6lk3ZP+nqwco35e4tHB
ZUD268HGYkA9PZwUp1LbDVsVM0QTK51UemHH8dCtTvDmOlgTDNCiUomXlwVp
T7DYx1OHelVRUSIjKZHnipivecS6VW7hrzZyKyc9sphIipeXqyDblzk9QOQR
mRLh69pjU4W6Q8DVTiIObQuhC/Oqsw+qTdUZor02hYGqGr5ejCaswETlzjo9
Lx0PSURGt8qcT+G3+Ftr5LHWM0sBEjKGhFmTrfgzMoCMzpOQdshrwFpkf1+l
w26vfZww6lwYTX/LMdi4uFa57ZbjkjiBbx0ly49o3YSNqFXtZeefbrH5AJBg
DaigPpowvFEWQ6piaANhbDLRzh01lSzplVe0PU0C58m9epIjcHv1fVJnM6AQ
SUnwr158nbXFOpHyrXGUEcFZKqFHNh3A/DtQ4TUoq/mEBfIYO9E0NAA5yXZk
8+9wjjm/bdC8/8JGgXDdND8hMQ9ytktMieivUHpyfud8Go8yZjO1n5dn+O/b
2BWO5CASJL6eNbBSlAERkm91NcwWHj0MkFNUba0U1FPuph4AzvyWCTTjJ9wT
y/YiiaDMPYMrEq0Tcn5VP4EhyiiximI7LtAP/7MnXTDYuolbUXe7JoBTaDIF
XGrwlPON4kjtCSpuIPnlIkad/2O0+ksTESiXsMFMPHyCdMPKkhj36qwvvvka
o7/GBH+iZ/Z/IQTfwWoaT46fQlaBFWsWaKhkRcfbqyRqqHPP4k5Aya50HsxS
bTViOs1J2JY1m7CJf62x5pJBycAK+PePRQbX7c59UJFlnD+0gDTQcNQM2P1i
kP7pAhhEtnhuADcFQ9frRJGzb2RBy++rlp7J5KJX1qgx/yElpfbUkEgjjN78
o44ie5YCujcS6xsZlO4vWregrvuiTkhhcssnvdbFl72eLqWL38WHZ3aZ7cUm
AVpI9WLJB7tKPBg6CFc3Wt/ootuReEffgatLLOcr0EevBHcj+UwkGg891ws5
sAvrZ/Xf+dPbAEh2R+hHeS4YPyDZUeIcJdhGXP9DBLrgiaQ3O8H1QpexXijn
zJ0/UiuIe+yHRDj95GzT55teSz+eCLvuVcvZBmVRW/TlwT18NIJbmXUERalw
f5kz304VNqE41jx3N3h3UWM7Y96mxEYcSnxnzo+X+XRJu56unXNrf5UEcFNX
qJcW2uaNMKq4z87btrtIUpyLxt6IbwtfBvvc7vDWL4jbXNG4WOyJaRn827qK
B0OFKmho/YTfV41OIurMzyv5QwFOfCvTvejNBU+XHi/bOm9F6QGHaJQFGW9E
wdZauE/9oKCn7imhftMpCpAG19O+9DaYYZ26Jue/6N6udyFv4pKjb+IKh+x6
J7IhiFS1lo9zA71iKc0+2hAS1ZZZKH6GBAssRTteh5LANvilX4hGgC7tSzmq
bMGvREGHyZuO58SykfRnJW01kuEbxeZhaLpTfaS6JUAsfv/9D5YP2YGCIxR5
5QfRRDSck9dhcr8wxvw09ws0cF5ppg/WW3IJdBtsf205RUPlGi6dOhz5SgPK
HWQ8liNGJi+2URe7dgPH+2ZKSQtOV12gI8FRh12nCYvaoehWsoW1BtRprwVL
xyqRlqRsn9ns/NIerGHYZot2dFrx9JKtTTcCKxv6cN3/HpJyNokP7piyMEtb
Vrh1g/g470pmUWRbAtWpBlxzRQ1co50qrpLStFiYRDsmunFEUxFTemPqXXzj
iY76c2L5Y7/fidHZ71KzdxnDNf8R0+hJiSL4zADXPr/N1RYYsNL/XvYGTIAe
ePDj8PK2kGVHW3dOnjVPA4oV60KMhyyNjsEPc0YLVOkg8I4Eo2OLNSSc9c25
/pQnOgN2CVhBFHHqgb2XCwJgc5AN5BEptdwtLg1Y9OKp849f13Y2T4ovn2rw
9xLK2KKJfbuI82d2ihG+xIdQuuUjierR20884RtBoS7yozCh885JOidsftDu
NcG7dwja1C1UqjbQcGCwmIDqHkyc7845Ji8S901jaxVg6NLq38HZcmwjaar7
LYqDKhcu0UJm9cvZ7IB6kjpxIhCPcOROy3wxAJ4belKUpNbfX1cIbXc/n9XW
iH2xyXSceCjIOGgHMRzBaiCa0rhA1ilHTwe52Vqg0pauCfkrwWlDL6BsEX6L
cKp/jx3U35Q+GNn6JwDO4/NkDKh9HgLo4UzG39bz0s02CZC2TnBt40dr4YOE
/xjqWkzV0NtO74ZaD8YzghZcT13SJS/YIMh9lR71+ASnOhAqKW1gKu9+OD/D
cKAQ0HUMcMh4nXqdEG11kYgOhh4T5Q3iRjoui32mC6jXGyYgNurzNHAGjm6+
KlF1pkOwgdDjV0A1SoiZ5aYuvuO8Ogm4U62yFU+POfOoyQXreHzv2bEGPIJb
wfr0c5ZG/JujCJCLWSGAoNfKL17Hhc3yjQBirCtOa4wE+FzJg5yBbdUaf2GQ
+uuHfoqjqqtJ2Vja+z0Sku4zXwe4XxH76ZnDg8uS47T0lpgt3MDyJ/Xl/FUN
6UU9ohJayEf0Mv+ygrLoe/BKFWDR3rrXyuwxGSyZZMNHVP9Roe7CvOs4OZfQ
UVvcULbNPoEeXa7uj7o1toKFuPbvAw3iW/QHabtGYTUySPPE96haJXPhvGLS
aZTNmDeiplOFaTBh16mDVUbD5rLObWEOylwFp08Pd+y+tskmOeW3+jjniZTM
5AeDwTqImSsgFlpgBcYHNBV9kMQbKfGtSxpUbWcIZ/OSpzlS0WnFwE/1wGVR
0WqAkF/shPUsOCry4Cc3U5t3cOBoRkgk3caU9cQlTlkAcRb0PJ2i1UTcmfkI
iScpAfn8+f4MSTIeKhKvWkQ7paHy5EnDxc4AJvWmtnHM/okO9A6HqbO2jKd8
0xw/mdWxa4/shR4wih2EVFVBHY07AAblcbBHIMsmxVwIrLpwfjRN9wWh4G5w
dp++lUhzAR4qtbEA6NUg03BHY6awyPSzOdkNqiPxoftqdJPzCa3C5VCdFIeZ
C+tWft1thqrwDbQzCPpw+AfXWofUSdIMOHiYlwvKPbz/km4UaK/AYIURtiC1
hxD9jqYdeValgCx98Qg03bGL64SNkqcEi34PSmde5IWuAen2RX4QoNcdBwsh
5PCqb/tJ6LpbUDn6Rkazd/NpeZJ8o2sMzfFCIcq4osh8qXvmkya5Gayxy8+9
0qT12rKDnAOZWgEAqVBwONjKT+/oCqrO7bLeNtvoM8707t/exQHCO1iB7TtG
tAGcp2L3IAFN8ce4aNifpitoKVvD0FW508JXrPL+VEe+qcGLTnRYTLphaQiy
VIa97Bzzn8m0ONU8bOjyCjE3C+gZeMpq3kjNThcl4/qcqFPH13aZLaUYjViE
Zjp2b/0U7QYrCo2atG5cOWKXdROA0R646ZM+VkBZhzTZxI9JqVpa+MDZ3ntW
4D25YznKeqn28ICdmhIwS92qo22mWlocsHYsGXVl/lE939KtQ0UdHUyqUirI
hkWBQ6B+WaBhpWseDdhZ5y0esqEOJsP3pI3UUTwAs6I1nNZH8MyTX+Tr1HAO
wE076DWqIjPX0OlFDJLV9zoehTKXrEx6drJG9qqsYVxfsWTg+7M+Q6yAAJLj
O+YcZjWzYD6NM+ocXcaTfQRHJ/9l7pNFZenq+oTLjmfTxckPh5WO4uv/RBvf
jjSDR7KoCG9VA3OQJs5SnaqQ7WbTYf+Nk6ZjtP75dgKxxnWnP7gJDAC4nct2
C18I3osKqmHL2noTsr3EWv3tlzanFXBACk7wWsGeJq3zRQKl7GRzpZmlAyp5
+cklO/kEkOUDAx2FaBsPpm0fOYUB1v5CkkqT8j9pwdDb0UDXRAl97INTaMhO
cjKtAAB6eyXjvMd7CDlvVex/K42tA/PKvLPfGAKL5EqTnwufoOEyQn6BHKjO
nM6dN7XMtJ+iP7B6BIEoyb629Wzxrp+qaiEIow2YW3oeCMSKfsLfElZAtblq
r9+xE5da6svCGa3Wu5+sWxsvlBbABLB/kZ1s1EN4BRaQOD5JERaD/OCrUUcN
DkLysVouytWrAl2EmBItkaxx8wFipRKiXMoT0rJqWYDsYkrfWEWvCzbSxqR0
3yj6dI/3w2s0ajkxrYE/FxPVs1mbWLMZCXZJdoe8ygfq9tWWpIZcmUgCo5wF
ppS/kdI6QDaVCZGZ7Y26y7kiLHcz6WF6FbfmjtdPsYTRL+BRhxv8mnvXStAI
ZvHvCjr6pgNwAUzWx16kbDQDpkmZhaq1vvcATtn68c4DIN2gz5FBiFqSnYrT
H7fU2/p0A9Zk+BmnpUuIxCe/xVs+KKOesk+RMPYi3icbDIQrdIlNpmxTezos
mqtkG9pLCvn3oDw9ylOriLJGCvgzvJz7KDJ8/4v9e7TNbHQW9t+aBi2S8Uy3
GqeigmNJME1bPSwVTvii1wI/7HsFgnaI96p/dYxqWjBgtaH1r8cL2Ac7BOQe
a6yFD/3tfFL9pYK1QB5W61TqQF3wny881xK7vgrPRXKC/CE5tjmSehgx8yUc
7s8aTlboDL6BjvEI2Yp/XpvFrl6JKEg6LpB4gbKl0bCkEpVZC71Xp4NLCyNH
reDB8PBsuAIGNO9tfI6zlyzCuAF/1Og91MOS+KN02gMOxhWqB2mPbXuzr0/Y
Qukq8uhvlqK140ke/9Eom6D7TD6EM/XFnW0lKMbRia1y4QiB7BYQTB64Xrlm
AyJTYYZ0Dkxs7pXsBSe1t8bSj7hEs1rpG4C89SiSyT4RvQmiodwQ++WjsNgY
wAye1VDPYpoLpC55eQDgLzYOAnCKGkAHMpwPJNTh1CvuZ7B59h+2d/5ug+89
C6dd1SXsLZd6/7TT56D0PCbvwjVPhWKtqfvo1ljlhcU2G2XtEQ4yFzbhRJRX
POXs0tCqRNKtGcfSuEdqk3L5sFQ7Yrwg3RgLYDH6DFNQcPwg+u0LFmF96zWz
OlZCb7IuJCvTqEj5XvPpKG0j/xNv4xPVr6tphU0tirN5Shr4MSvBezAUERzh
n2ZZu2vQ3yUod+QQcf+hLBE+zT6mB3niepaedjpIiFCwjCQxKDVMT3an3tY9
hPeDONmisABecenjbjxZWxBLuAVUwYW+ZfenOKXyehDmPpmnFO3JkOk1CbjR
ekl3gnTAg3INWDyhwpfN9UtLR+u+4R3W6tbLWGM7AKYfsW7cTM1YIFdhh5u1
JxYIN2/9WD7x16a16OrEzLZl117iK0Rqshuhc4EEi0hzEeGph5rRbsusW2RE
OyuIKQxwXeevnGDsQFznG2CsE7TjGLPWJcUALfGUcSEbQZApO1rjri65U5hi
9wprIO4ijI24mzN1BcedubPpkXep4GYJjja3N4RB8+dzEpawT6jWcdHjAkv/
n0Cq5pkF408UzKzTh6Ufxgt4aqQGKJwNJu8uBAKu5ZzoGHsgbbJkAfWIq4Rq
aZ7n+CAoND8m6Ae0XpanBn7e45ZSzyvCknARmlNUXKym30XooKyvapipy1Uh
+yJXGuNO4pwP6F8sME3lEcf6n0Fu/yaASCF+7G/zklWGin3RUT9RvkNULoJ3
Vt/D+XyZtCST0Y/5+P6yERLZw/GY4QMOiOlBc0npQ/tIbPEJN96oeAjOZBLa
uO1AwC6rq19rPs9yPVCteKbd8xmh7G1cKdn1drnjWFSQOQzEvz70FAlp5N4Q
k8Msm+eAP7Bnf8tHRXvcowwJ+Py3mHNR9LizRtrqKJHJrodRDDS0dzR+8lOD
IKcby9MIVyfrf8385TSo48sC5v17yo+Z0efW/HbqP8OmpcJMUFwnUJ510Pke
faxzHkci+b2EqDH0Me4IkeHZhNLuKOelMTLQ2P7Vnyj5sUhZQ5EmtzKTWG6t
7yCPIKufJRcLvsveaCr7hDiehvfq6YEzZIG95I9+n3UXMBQs9atM87Hn83Rm
CUpZRX1aZpJKtJWLlSg8xhNvsIbg8vrKqEH4Ku40UaBE9AWA3Y2gYpDjyM+8
vOhfbYw4e8wWh6BH/UnWpi43Hjqv672ZLKIUovqwhfGZXHVWrnijmwyvgkuo
mOoJtVMJ4YbnxwHfNP87BkVDuAtos0w7a4q4W/s75hvGnFeqymF1X6VflwXl
vQS38eoF4ui1/qfq/Vl7yLNmM7AS01RoHWMsnKxlgCe6R1Odn0jme9cfAuZL
d/6O7cdpnLzPhi+7P/fjLitqIg27nQuCxOp+ghEOK5XGrtATIcN3pXVlp+bB
pjaSlSqkFOjs34Mpkx4aigjEy572vh7mZxtyD3OJttHQ/YuJ2TDpaucvO5Py
haOuv/lkAKikQq34EKbvDxgzPWiEUlwkCGO9zuw1Q0pWozsRLl0EW5YPkUwM
JEzCY5YWTdz0896IX4Zs9a0O0Qrg2vBEEdPRtb0FvKJF0DtDybTmXPd2WgBi
g80yYQNH7sjZqy+ahQ0KCZi/dZ0EO/jfaXp8CZlSMcgvixqeNVpGigI8Y/X+
W14y0dVWVHAtlk8g5cTW2Yk8DmMn1lYkJBhyt2HQo0enritf4YfYDMrtgO3W
QKhLAO+1zZxrh21AYi2Sgbdlv7FVLBKlE03O/E1ApixgmzHGiAB/kdeiUXiM
UV6ZQIUHk54FZjY0mmGIRe5mi79Wj10AFzC1L/sh31fD8JQmqd4k71En/moE
vQlfpYsqe3PsvC/DTVZ648Dg0ouWCEJTD6YmNAWSmfnnQXHH9QtQSYlI71vu
T1QVEL43H4OEHRDeSx7Rfeu1U4jQMHUcWD/nhJqN8/cAJ5Y5e0Fzw2uerhmu
+0w+NJvWSjMm2uTwt26a/e8qcKnqFtNUp/51hlUhgAIoBoqVg58uvAC0AzP7
RiVjLaltGHutahdv+8bCrS2dprt2/YqRcQ1ZgyRly+8/v3ntrwgS0FokrCJo
HTdjQ/Lx9xfE9ZV60RKHoZ3PXp5PeCPApOqMv/7e35/dRRX4SCTOzlgH3FMI
c0dhj7sQPdQDnvQZrHLCtzEVZV/hO0zDQLdQxy71ngXEYXl5JuRtquYVsYlG
iKPIWz7SB8tO3+8k6Qa/0WlG3PrPUJOF5bSHaC/5feL07r2aQAYXdJUN5TlN
8NMS1SW8V4NUud5hnPw5UabHFjhMPuMX6YWjMJUV0ft+4hNKGRiAsov2qSMY
7g1R/nAMf0P47Y3Q83P+wOTcAoSSj3FdwK336c6KkKSoFdyl8jgkXjz5rfuE
rPbu3iFE8J4ozkrbcIS2PK0X6/198HlSR0c2MHUaV4RVF9iUrbvbp9iY70d+
udI/qfIRPYqqCBHpzxakSwD8vmAk3bNY50fRUs3LpHFmu9O/5BLKipufg9RG
EshtiDnrEIDmz4QcpcsGqX1mHAJhklAXCgCsEVOIyGuvgZLSrYxpKjJYai0R
x9u6e00yZVensW4VCqW56OJZzB4HASzO1uJ6iaI9HYjBkLayFG4tIiX9l3Pp
O9QJvSkSpfc39ag24yLKXqxVsLUCeXm9xFOfSc0vokJdKU7Ajiaxjd9a+16i
mfnXNu+jMg0Z7c7Ld6ll1VqZWY4tntv3lBw91r1Wcgaz0BnD+qLbfjy46OCX
aIpQIquRk72UfTI/uWrc61YEv7JCO0gyNiXznqNC6T8vRQr/sTAlwlbd0UUg
dKTsjSq7zg1w3JT0TQ6YrsYO6GjACINQnvVKgwKH+6Wmg2XW7HuJSEV0pNHa
q/51ic4XyXGs+xXdAlgSyc5yY0CxUxhkc5a32EFDw3VqW5wQqQqESGwpAcnm
ilKojOO6TLy29hmCm1Kk9oL53lEmoz2kXkVMxwQ3zY3EHqbAr+/NxXTQgMoA
u1g0MnAg4whVh0lHfQQG6fWk2MHvfrw7mzgHbg5Zu91gItyYeZHmVZZm1vZm
QDdC9Ys1+M8aagydsVcxUrNC2byi/zvtBW1QYRbO/oL0rAUG0S6R+Myk2KJ0
8+IpsOZv6LbGBHogzYZZMmNLmYlnjPOIW7qcC3v+K5Vve5VfHRfle5pv1FgY
RVHrseTV2mL0ma9IibanDX0SeH+hQftNuUcSrrNmZeyHj47SasHscS4Gu6PH
NtQuYUfqFepmidFPoKCXaeaCZgPr39ywFRqrDqeQahKOf2m0x683Gpea4dlk
+RtuZRbbOWLCnjW69eLrCHLtv90KvcXZikdr78xSRb3++Xh0SSHi0chobN77
UhOCnqot9oNevf3RkGmup7KYZRicHA8TPo3FC7Y+9SWpuVWPd4ebAcDKD19N
mikbIebZHzcHZuwngQiEdfxnDVzqtieUQVRio9PpUbaggiscJPWiGAdj43eO
x4h9Noe0ketXO8NZR1lAAR8baT4Q8s7PedBgz/I0ds36/+8UBvtAFUwblQqn
DOyJUAwnwYQDKptZ7OMonKWJbFbBjhnK1TgGCYv8BZZ6rgo85gII/aN3PX5h
BYWIPhKfJozzkDFjTmw9kJD4Pvdr0GBga1kpRNM0WZkiP1MWMOElkhr2ld9x
sZhinVpkokbS2tZ7h1v1hft9DmKc6TkQDMPAnZBmIlMyHZHJX5OHudswf4ka
Zo19CJQ+iJG63X2roNXwtaN3FnTaD1KjR00clr5FKsFsYmVHdlE78s5/K9UN
YzR7troSi8A7tMqhoL/tRIf4xmeJJ0UJHeodx6lC/xzm+peMAhsl7gBEO9ZG
HJq0i/yfQ09olOZcNyznElbDaGPg9ANBDmqClZs9COFEjb09KQWCSXUIyYOS
YF6kkmvRLopSBEmmpcqASSWVc+A38zeci3pcvocoZMumtVbiAHvKVkx3MXHw
KgClwFSpZKKXgxS/WvGfna0PlnURQXKhmSH+yQy2UD55qWJ3yu2KjNkSwQ3W
48engb8XtFKXx3uiD2zTQgmge1RrRqOk7dJ90J+cEY52E5wrZme9Wloa1TAn
Jsjo0p8jEdQV3dqbIfcXE/IzCnECkE/Xcy0FRhOMe5RKL2HzwcB3Jebz1SMn
/cSX2eTUzrMsHHpDSip3xNhqdgBw+PeF/ckgf+aw5ZPweVxAsTiXENC/vb2l
RV1qqpGOqtdj4c++fglHUJEUhxEZbsE4TQG+x8j13KrqURcm4n6X6uhRqlLl
vXPUXpUaFXh0nmo4cZ2/EP7fJ/t8Bzj9wZeK9p7c0BI2mehwWI3mJDHUf2Fo
1xKywmI9TL3Qv2vECGZVFJBLzid4wBdy6yx6A6UtEA6umEI/sopKWv3h+Zq+
w7CrVpY6JaPjp5k00AAHTBcUsSoIVvlB3cxL6N90uzJFcKeYfyouf69sEP5g
NbYi3T7HPqSv5AkGlxFGgGQzISJZ9raH9xiGoMvnJLDPYm6hwvk3DcShXo5f
MstAaKmXwbeh6eVIqrSSknAfEeuNVvtljhVnIxik9gsqEBxSEuJ4sQSmbSlT
OkNDxXbuDi53JQ1knnoCse90SFHniuHw9+a6mj9G3Pjq4siSftMxdAZveDK6
hIFI34GwY8UaQ0X38BWbGK2bNNDEZP3qMBEZ5l8buZfpKJ/jZZWeF4mjMq2w
9lQNjrw34l3tSR0VcJt42Y2fX5OkdabHFEZLty8S7z843FCjV+xhSW3GtgYT
Ci1bKPLMi0OIJrBsUFut800YSvl2+GPHX49QrB/Htv2ARvuRQ6ypiMXdCIeM
dnR/rIcONNI11GeFzfe7DpWi+vp16H5e4T7msUjBAz1c+B4u5yHw7cGEKwEp
nITGux9dbun6ZxMwX5yIlHS9HRzRVGZba14DEFECR/BMJ0NxGAQTPrzuJkCY
WCN//yiqmUXDvlXXmFekf5zon1HawlEe74YIg94l5pRynHVUnnMsepzGtBl/
H8jDvs++2bs6/Wo93Ga4WgzznDPgcSezsSkEMYmKdFvi+dUizuTT7UWHOPyq
J5DAxW7MjSwXG8KSlf0aJXaYkfw2XZX58nAykz/Df7zsoZvWRluAKkfbCZaj
VbMZOteBnhG9h3rL2FJeI1RnEgkZVpnf/aPqwNShA9liiKj62SpuD0mZL+TX
wzgjkyDHz0GqY1dEWub07YS6dw84ATrUFHt/mbQMTYiz7gGWcEiD2hbu6Yn8
VRITcHr1JvMDHtM/HKuHi3SCebGQW1adoD4JJhGeMmTB63/Okqj/xfpLHm0/
UdaB4Nw+tzChm3x8B/5Xu5ubDOS2J17jt3m12ntxvk31iKYXvBmY2SZmhWh1
Syj4FV+oPXa25xTVxcEMD/F0ZkMaeSp0RCxuvUnXcRFQgWwmR2POlEfJNhx4
M8MJTS9b/bOwkTLDhCGgGbfYiLkHr0hlksg9o7OcE3sCnxSXaBpJU988PRru
yWrhvx69CwmrCBeqP6CIpljXb5sZSsSbMhgmoyMiWjqImB28HuPmY8NZ1ZDW
8JY5AZkdD4kaRnnKwddOgUD4Xg1ZLzCs6cMjpZKbsxPZVa6uKbcYcTqZsbd4
n3UQjOtWVAw8yTlF/zCJcepHb2zMG7dCq6mU0zbHgvZTKlTfLlFEf2IpgH2D
a9mFA9Tlh+QCkgtYfzI3wvlr7aImPhp2habYEW3d9+FkVmYY4knDQzK+JEiG
Dz/fo/IwU+JOHnFP0aJ9oQzJbrEDtma9tF39FXz3GpKFgqsFuzrVrXLQtwY8
go55JEbKcdOecmjAv9C5RQjEqk1KtpwVSx+BQErP6f+baUIBwySocWUw4jN6
Yya2ZCVoiJhg795Cxqzu2XM/FunICzUA01GcOH4CcJYlhojUOycxDb40sLLC
aIp1NCkuUuYLHnCSD6v72NA+/a773vgTx2GeyvbqCwHWPAD1WXAXnYk0MGxa
qApmvSxFQvkUDIddXlPklujPpWgjcFjgd21eIEzCZIMLQLgvhsZvOjtB9YXN
rNc3ijI+/QboV2Lp0uw6I5sO/cfdeyZlN6tutZOyYjh45cC7J15FvvC2BNVY
E01xKF4wpB+iLltmQFQ8x7vASZqqGjlWD70/qcVpc2lSG4sYMMavK+5A7Clr
rpMVwZAXh+WhnVRrQDdjFR0/VlNodjfQn9u+tuOpjDr9j+d5c8q6bRECLVPn
goElvlKvBZZmTCdyVgwyfGkl3G8TVEkb7BB9jCVyrEzwMF6yAlRjhHMXgHsp
WQyprt8/37XIAyJC9Bci915w4wZzT4mc34dGFg8EZA6iOzgXuQnbeiXXPFYa
Xxh9/7CSHZmy3zfr1FBm6lUCtqhGbBgUeHxoopspo9JmIMtVBLlEa+j4tgDn
gPRocC1gvsOC6LAKg3OVIFat7UBqGOImZpU0epzLDGgGHHzrJ+cELjCdfmAj
AH2KWiGDkERMImxsmeTI+eabyB2tvgr7t3lmAvtgDPBr04Sa8N0KNofzy2U5
Ff6a6r03CsoMgTgovLnS/hKNMtOBGHECN1UpWDp0L1xE7jbb0hutLqpVJtZM
2j1rpYJIS172P0k6gKqJNC0bpvbs3KXSYxFyv92uraeyeTceZ6phsHfd38GI
cOlunDvJ8CagLLctxzUrMywXjVSsMY2SMJvW0wFVVWcIT9/K0C0E8JSfe/Ak
Q3naK9eezUBhUSHt584llO3chedPhZkwpbcQIBiS2MouDu+yx3Pt93rWwD87
E/f8db7C7W9Un0mOeySVimX5mnFLrqaq6fAir0wBqMC5LYU/A+1YnWnEtE/Z
AM7UZYR/AmyrUV5nksSKVkxwtm7lgnJ3P7YP4mCPPeuXbQpoeMJ+vS1u6CWL
4r6RDu5vJFRPheK4i7i6r0oYONkLp+BFzWeJos6GobHjPTOh9JQxvhpfT08Z
lInyFrpQIfY9EB7I7D04f2W3oxMOIM2zaXxV/y0VufU2WlyAUBvft2CV21y0
Dj2kYh18DRNoauiWXtx875JfVDKp/YiCDJAXWMIplSqxYfA2zaem0IvMDMxw
PDuErpDBaBV1nmD6I4eeRkTCY6MCpTS95WDLIXr1zAhRD5e8CsfvCQHzEXPu
zz92pqGOFSdHAENF2ntUbz7bQ9O3YfWYSV6diYyaPeFrnSVme+d1EycCijAB
L0FTcfD9+IhS5sHE5I+xYrO6/Wl07xLcYzW+ZPpAJiDSkk3J4JwU+xYe0l34
ayhRQOF3WvWMYQkXtWGSR7LYOhRBjmy6uyxehyuHDW30X/pORBnjJFjfwEER
CW041eVIBICYGFv1b77oRiem4KITtJ1CzzpAwWgTFTr40asGqdz1O4Uv/NdP
Ez/GHB6O26lnJupKqtlpNMnHOP9WqmMRKvkTE4nSNuX2v1Yxzrhi70DfIg1c
Scz2ZCVwQAJH7c7JhsaF6UdzRYNGbR+sB3qK/hswDSCJNyZzfkgICSsvXLhQ
qAwjugTKykjO4iR502ibZcgtmKTom5y2GDmway5mfIQSto+2GQ0hX03x9MjF
qb3mG3dDnKMRRZTQQj2OLgT4vzx0iAgqUfQk0LqWP5TWl1mVZA+DaB1eTRvB
yIsyvsfBcIeDdPfESpkl/7NLUo6ug49TLHdo3WcloWIha0YRlaNldzH2oflL
k9O/BH26pvF3Zjav1jJcKhvyRPLLnaKGrfLmEyiz74sCwq/TqmrPFR5/jFB2
mk9JhYAFlbVWBW2Nhsm7jFoAazs1Rl23EXmQj6Jo6ikmgtPSI4JoI/lfUvvV
EC51wAyqQ2+ehWfkf0SRo/d+YDFEHTz/4k9cTeyi8VW8jPlGZBhlL8V5CxNg
URw7EuWvpjq7s8iFc/P7ElvzxGpv7+yC8zN9kxhC+uLhJZaXvpkir/qxQSk9
tCfo179nmhMXDJRYkSaIzXdmVkXL4D25OGp54H/ZgRYOWPeCSNR+Pqispdq+
i7EXqCecHkxn0Ce2sHS8zvRlgaAl1+a510k266ksdR+UASP3D5RJw+Z4N25b
k4EfzAQElVhlXUtLmzbGHc1kiBLDqUv5nVIxLBfBE6IF47/N70yCf8MWSBQv
jhxYjnVbCFYIwJyxGbAA4YkPCBDo7n/lAGPgXi35biboS/7Lbthm9lCOaywj
seSnN5AaNuZYRrS2FzNqBO1bxO4yW87lSpCc+mAESPjrdFHW9EnWUWr+OB3l
uiF6bsePQH6otX62WBfz766bRcPAn3LGrXpzAl1CAG4Y1e6Q1LQf7OJSKG2N
MEpshJuc5vYx7j0iHfE+h0CJiBjciDI61DX2p1wgaSYJxuMeA2spDx6xkzA+
HGGpEwDtbrhdY5NW4IX9IsLR5k406FBUnNlMRkx4aKrf859HmT1ZgqLE0uSq
hQCgj2Ji0tVcIRzps9l13BKhuv0lGHlymL8QiXz5EXOD8Go28jI+kC/sPG22
fQyGxK6IB1rQHZQ5dvmthNJYmRBKryOy/NRv/C5/h9WwYztIvy/pavUSYzUT
Mqi8LJAQnABfF3yJ2gjYTR/GkJDt4c6MvZkZs1bflOHb5KWIpeQtvTvZDmYi
+UETqAG/QbqaOZTUmBisABuGt6kNu4UYRIDaW2Hjk20hM0jU7sax8vLPgA1C
zb/uRZMRK3LJGd9GXvHAdfm1NZhCCvfX5BrwY3h87Jrptu41vfG5QwoMdKLU
4deT77tSWJe0/ZHzmdAUe65p/Ch/UOHS1E45zgPeMG2vFvEFKR+kLctfyWiY
wek9I/KkKedmujlZN+EzlfzaTV0qyOI4NdjWdBBiirW5JDCsF8Kp33gJk14O
xvk37LrSVikk7OWogP49XBzaLTKGt/L6j7NqdNcrG2oKLA7y0zL6vynz5XKl
vGYSf6vPdRcg+8PenBnUeWVak+8I4zNW1RL18EE2hhDcRSieQK/zU/mZVDqv
nh0GI/B8RYX01cBYvyUa19pabENiw+XxcTYxY6hCiktTQhWjT2gsCIQ0896k
Z7PcYyNUBDa3sOikYtcG0VC3OnESD4QCC9h5Ac9KD1WRJOcV9uNUJIk+7ZhA
ZN5AnecIeQ5KqOe/tQJnwIcPdka6oRlNMcKq4bfhTVbeIvcsoj6AtoxVs0St
kI7juQ7T3kfNbr6nsXnYBxq3AmUXptdy23+7mQ2iosunQVbBLGo+WYgiEPuB
Y2dPm1P7EcxaHtlSHrf2J+1t/1y6V7ogRiUT+5+pQgUgGp4lZ2mEcwqe5EhA
8hN9KT3As+OdS7eryGQKz0M65Vp0r7QhyG+S/knYfZhCNzWcGZfDUhqaQ9FV
zWbjGNXzAFQGl025lIPgCfR34hp+cZHQv/WRVQZYaF26/aZnqquH/RVyT3Fi
AzTAeGzNxTVGDT6asRQC3y7AivGpb6HaU6DxwgKzpj8neZwDYBJxXixhGV4J
NpD3D38MKoLY5GkrcMB9XeR0QyxngeJBovPVZVc0aNHdOGQ5CYOa/fpoBF9V
sQHMpRHT2n/odXNF8+vxD47f6mO7hwWCitJpyrvdJMWwlWAk3lAPvUX0ce4e
nenZWzTObNxn/fQ28OVqQD5rXGpzHPfo216w7+pzW0Xo70hNBu4zqOenFHgg
ItH74maeIU/MDkEkZ6YUSmeh7qj+gc0tSLVR7EqoSfiwwP1RZfR9tRLswGOr
1bUtiKda60bLnzjoBbGx+k67a6hMaeNlb1GYI2Phgwm1/RYSVWng4jBNJqSq
CfDV8Z0ZA0LAV5p3U2Ihiq0QD72McEWvT0bRNQywN+wVJPGkqVSGcoNTB6kg
SQAJt5/4+0XMZ7FIsFB/w8lALF6cRCGPshCFrNyVGULIc8B4ixEfm++vcHdV
YWh3jvqpKJpP73KHu/zQ8+XDY5FxSLuzyOM9vxjaELw9C8hBo0JfFNUlzFBU
bZZiKP7vyq9mXRsrK6Wllq+xNRm3fDOYwXwqqDPHj74tFwBJroNvBf4MKSNy
P3f7JtT2InrXkCePemWe83CTK95qnBnRjj3s9Rojlsrr0KKMxuP9WuGKGmnW
hKQYaYjL4tEM8EXoMa132awO3Pv6pX3uM4VDkbk2oVVW1A1XyNSElczDC2he
xwiaI4Y2Vq3xN62IGAI02Cy5FTNvVF1558nR3phxhczC8XR+j+4i5V/eTVgC
Jbd0dyOP3Yq3rkmADj7vflx9pyHEX1Nt37RZchRw1YWSoUMJ/PAuro7THRjP
tMCILzx9ruT9sIfEISTuRJK/JPHNexdJIEInCdAZQa8gQGpVB1wBsUZhWn/C
0NtGdKIczS9Zujyjn2Kk4OYDHt6ITj6J6kFhQACgGefdwG/kRcK7HDvlh1Oq
BoS9qi34mgrPLxaJbZZ0pGo7C+cBcen2y98xI+7y2/h7CdvssuUdU3QV/X92
VBe6CyWaJaAsyOCtAli+IAwKuGSL6ItRsBX1IuSx4nqGPd+MdiBjO9t20KjB
lDyCe/3Vq8yp6X3ew4QzCWZ58NR+pTyjKDULPUue9rOm90MbgbOEF7NwD51T
HyG7DIqjzcKyqMpJcWBqii1f/T/fhRHUNifdAk+/d/A21bUrVyO48cpdNt3A
b9x4/qB8xSxOqAY3pH02bF5rHg77odp424Wrc1OxQqaICxnVjcWdsDlHKJGm
hRCTArNxFUbMfeJi10RcWrfWmJuMdnSY5cekYQdT1McfxmYEPZyt4f2VwC+6
FyPb8Rl56O0x0fs00LYUY99gWTKuPGnibfAEGMoIWXeisOrwtYKf3WQZUDdX
DxzymKUIP8uG6pm5N1E3GdEaagf0kM/5dwOrn17ACokqTb5o87rSWC+QBzyC
WLt6WazXkujqRekpQkRHBr6xWYQtjCOuBniQDkmW8USWhabLmdSh3UWt2z7Z
cXKU5Le8JXJ9wzhSoh0qiWglCnKmF/kRu3Xd7d7U0Rwk4fCrBS70rCZ9ArK3
acoTxEg56IC0l8KiMIEPFl1TlGu/prl9hPaP62yAtNlNqX21lKPPLKebNyJ0
wnVRPwupOENZ1niBJcgVjruj3+CTMu4xsGBqdgptOhan7xj/rNmvfhWYwTKU
niEzpiE0LIEhEJTDt0b1ay3gX9zPZp5xu4Q67h/GGQLFAi9yPjH2LLahbr+6
VH9QwnklKfOYzc9HWty0dqX2Jjt5cimE3s6iyQ42DvanbMNueisMszVqMImO
ccBWEi9lvrX+epIEoYAgR6jotPSn5jGbWa4QiMLlHW28mQuIHlDjbLAo3KkV
stcIw9ae3UUGfpBZJUdlVIenswVG8Orapeo508cwRCftHEm1PnqU+eyy8OcE
xVD44jEndNG8lA4MVrc/oE5cuz84j4Eu05X9v3f7dlKTX4Ol+haASVDNEcKH
XVpY4yAuYJq4ISUkz+mNv5J63tzaogNFhq6FsUST7ailPwVcVGQ+PL8lgTYk
yE7KnIbxrtH57hTUZIOHUMo2+DJSelIwfEYH3MKqMWLDuJy7zPvPNkYv95jh
ubYbqtQEvpIKPN3iBl3UfllgUvrRMxkOIJ5RrAfLsyPNtKXztozRtWLhjH3D
2w89dBKY98V1o5HtQtTaSRgt6OJzMc/0KagOrz+v623XN2UiLUYpOs+KV7af
Rt3YIXjpjBjKpk1j1pQTtKWpGjC4JYfq3QoGEYLDYI/IXlDM3OTWTOoy48XC
MBB9OFAyptrud0LnZSEJi3th5EpOI0Dyd6355c8/+UYNgkmKfj4Z/EVv61l/
TudRb52Uo/odsoIxQXCwlPmDe/czjpBkqPtwSMsoSGFDgdwevEWIvqhawuxd
jm6EuuHP905VyaEl8wpE0i2CvYzo7NFUYxt/YrbFg/ZxoecsVpNzRGKJFDfr
55HDn+Lm3QJKwulLWpP70hW1QM3ffDrhgQZIpiZ+DadQgJV2Ylp4VbrT12ff
kxabEevndeMnJ7N52YOhpmTpBfYjL5TMsVGiV5LIb+QdBAgQe9fwadtukTlL
kFFmydsZYGhA0mKqkE7DXhFkCGDedR/eWOdN1+EwzfvEH/hNQyisnKozfIsx
aB7hhqlWTWaTNv3or22h69osRUxFDiKPCYqPr3ajJBDm+YgbiAGFIiNfK0bC
3D+wZJFor0y0W1urPQqoVpEc3Lfi3XookIiy78jpb6TxskOfcjFvQeM1Si1z
85B4/+VI7Yz8xSOeu+/yfpZGQuxRKUwE+BwDOzJUaEsR+uErp+PZ/fwFU98c
T0SnjP8P7SCCdiWg10wx1Wd3KkYcbUlUxE3UfADEgPZxsBX2s+9xXGlR2E1D
v8NWMO4gXEg1wdrpTy3Y8SkxJFp7AjxeHgJzTSeFB3TkmE+aEA5LrR0fCfEX
gIhEfBR5NE6sLgTx/bUDUcVlErvF6SVdtjgZgFKn++m4IGs1VZOZj5mThWxA
65l6o0MxK2JvkL+SNsEo9heAIT7+5Yk43GLoxb3Lsg4Pv0m5vGw2wCBq6Ji0
Nddjw0AeBtuIi7sBtwEFLVF/G8qsaWyoXv5Ol1cy/gAGZXAJ//RydyvV7CHa
zmsmNlF8vhCMgNSuoz/H8gfn3JHlGxgpRNgWXGDZlTYNo01OykBuQmklLEF4
sOxOk0y0ORon1U0VMk1gSm9Jgq0NKuET+E57u5umQjWY6odja5PvxFYjn0zK
xQTk40zVzie20558fpr+G48wVud8X4y49F8/qoVKyacr/6n+VMKFr1KeuKXX
ixkIYa56MTbT3yTbH1cWfaSCDQViM3WTDrypyXvu9m7Ukit3pF+E4qe4UzVJ
byDVMpwWDwhDe4OQZfLlFrmm3zQgym0w6xBjzfPm4/utdr2UT76bh0UdvLZm
9mENqYp3iyE5Zh6C1pKqE7sWkyT6SN7siLkOhQ+3EycSXdEqEnHqJZLH3Bgi
FmMwqmtlXLrecIPIrR3IiuxTMza7nf2OxBcH+pf2syjeOD7GqfQHYNNqxOdU
k2HpLafQMt3X9BkOzuXJONIyozT1YbS20gU6XtCLaExrzhkUAsX18+gAoY2D
BaRgJ2uCgeX283e5kc7PvEDo299XBK/0J3nxbLdfviCXLqKEs3hWePdyH5vP
hOxRRhSq4KSyvBX5fVO2mdcH9yRs0IUpLGLocdDRc+oi0tNkohcQmG3stE8Y
/jPpMSocjdoo3mJtULxpXonh+WGMl8oz8+zw5iLqaG4uQCwQiDwfGZNp0xEN
HqShwn4ufHa+mboJWv+EkC2wH0h+KASO+iD5i2bpKy/MDAt7F2r6ajWRzprL
StxDpzuJlcMnnTLN88MLBHy6+5DscYlIR51W4i4NbmAgdra3uzyj7j2+X1L2
/+N9oJvIsrKLAy7h2oVYCMQEt4vNQ5YQqApgslpILDCwjxLUGtQNf3sLANip
rqkTvMAejTD0d3VlHk2RCZ8kCh/tntlTKX8gaQsVg5e1/+oKG28Q1R/uhBlD
ky6ncHETc0Cf6x1bLSBwxHQnZr7GtPyVfvlPWr3qinirlz8N5BbxSBxOy6gO
dSfCTXDnR3ISGM+YzcB8c85b28gzKMcnFk3pnxu2sSQY2NScxpx0fmzuhjYH
o0H3Oq/ixqTKqsRRAnbYJJgwmBGnKdjtcnKDMwiy++hbtcdB0yf85KcEPAs+
ccn8yZtqzOoOT2k8f6W99i8JXkGnctSGshFG0w4EhNRHkldQvV3BdbwYxvQU
MUcaRowDLk1S8QAXMNQIXflfmxfQHTHMOsJDA+3uYI+uaVIrmBVlMag/zUnx
ccL259uOiU6GokwVZFFs/OzvJiRouMpa7YQqRRFRukswACd9v7/8oKebmda6
bjvBuuYUuLp/tVPRGLoO65xn9Lu0YAtT3vPxODL7ZdUJLWgXqbSG0FcrY/si
BLtiSlLoDVx91LYN6n2nQnC2Lkbdf+mXFOTFVn95ZNOXofekKRZxLqvTHTow
5Qr9hXqca/86nZUDqJDr+KQZGM64fVavkuFMNwPsguKXS+syH7X0ukZFscrD
jJ+nXF5s3ihpgu55HqvF0NeeNkJ6fQs2UwtHEAPwBXXXQnUt10end/F8veq9
d9CC6AViRuigrjm/OFpGo5SjRf4P/etF9YpjyMQ7C0HRBS8Ag/D53S1pd7An
LrvunfHbdD6BM95prjUv43bPyntZr7uIDgvnQ4Spz1LqOqqH+n/W7KIopt8X
G4g8s8Bb727bElm++95vpnWLHnPbsOXxCqf6k/3avBZ4gX7LI86fqjeROZEV
xvvD82K3YQDSAdFL3k9eXeuqAQPgfpBlAOHW2m9l08VSMUrlSRMxCOTAAorC
/lULro4ie+0inYbZDOVRUYX/+8RyafCljY9pV0pGw9znYJlhxRt/J/ycDjUW
POi5FfrgCvO7fieq5YOMfBMh72AwvkSMmFH/BR9pmwuOUj8DW60m/4yBeyW2
4kTIJg/qUa/be/jjzFeE808XSsOoI39VKHPtX6kcT/nA8mNQr1eLFi0b1gh/
Ikmaz+UW9fo031WSGXI9Mei6cS+8fln8yAJtGHe0lz3tSnRGbVrnsLBtUAW+
DK0sWOaX8FG1mbpw5IiAtv3DRXD7PLduwqC8uaHUZVdaZOJx8eV3E+CuR9Mq
4cfBEbrI5tGStjf+G77jOZVF1OQKPGxXg102Un3O5zK9e457dsUW2DUmto0f
iQL6fNnROO2Pih1QC3nBT8c4JFWdRWNYLh4WFBc2TusPujVDEerV8TzX3jn2
FelP4MGqE2JgbBPIyx5iUVhPq3Vv/K6mpRs930+SOlTA5J0jTwUYxRB25SfI
ccKLo31kG2GCMB4t5Ko8qDDu7fXyRu2nc7r13zori/1PoQY5Bmbl9QS7JeQj
B0jR4nERO+exZh9CVSYsnfQbhPjvejQBSBRwepUCkhmqoYIRNxGUJaWmo61H
agaNPQb5D6ekNCl1IKFRqf4joMplrrTcmlOf1zx9CXJdYzvLQQQvbGveBsxb
pjzk0FoU7+JMsKkjEvWrLQuJfgX9o54SFaLRI/Ivzfcb+RBisWpRFaXtpJZu
vl4Kp9Ed80vdiTvTUCt709msXBGP8rfrzPqL5rImaCDilahZmWETPvIDnaT1
RYkjkFsv1KeGXB5midSbUq3LtysZEgEJcR66+aAf4hABZvXi1ibk3VzfQYL9
LSZmQ3K3BN5YDfbdXY6/ojjkcJvGEdxVgyeD6lG/x0c+lqMkIHJTfMdk2yTV
SD6qmkYV98Z764erjX++p1sPk0WQn+1kavsr5GB35lY7Ko3fhuZJfHgMgU5l
391mliuUdcLoZquSS1oT3ITGN8D/kw8Guc/RKM7WnadZzLLIa5fxsvA3NECx
v++yJYsJmpmOuQk4NaCj15USU2f2Rc0cA2H0kkn0pfmOuxPy8ksoEUyx3Jv6
glEGninlR5nXiRZYzQgev1PZXSRpxoYKMDSWGMZMN50a9Z8e14FJ0hRBKsSE
llFgdyxIzb+QR0mqJcvKUlPvaH9wRjKZ85ZlHeIedONvbmgbQc1RrSfbTQ1b
b0NctXOd0HB3+E1cxee2Jk1qU9iyDX+C1CRejS2DRRn8871RBY7Qg54MFVrv
zomRI0S1wf2tgZx5C8A1ri7tcUWMroCB29rEilUtKrVP6oMkO5/CgKFhHLoK
H4T+foe7tQV4DW2hXEr0FxQtalW38x3FOMrDshCtr4NGdlM7l12iaiN68fKe
BUuyknWD/C3/4THEMUcvNIsKZSBXPk7Jj9xpieHwMZtErcljjBOvWieYVHLq
pnYUjyh/xfz0HTpZ72uDwCNb7gcyJujVMWxuJk4zbfvdA05aO4WBJmVErxV5
7QBzIlRTkG8TOTmIK+kice4UdI+zImxc1Aw8opMXUuKoxMfwl9Pc3Vh0xebL
WbGoMgR3xBc1vu3IEqTv71EtYq94466A3+fqOI59BARV3bLeAKFTO02kO5b3
w1DXxTShB1SjkkFe8yiVtmltNvjnIdw7FgyySEwQoubnKsyjFQnub2/CWtJQ
DDmdV+BUbH/IDWrkSWYxLTHaOHFZwAg1ywquZbbfhwywN6FAnMoAuMZC7I3a
B6PsNhkd/1iIRi7K8PCfqmkUxFO1y/k/gnJNGCO6Ao2ID75hYOgrh9pZTofM
aWOKf2G7H0kUM9X1yH/WJOlahUNLpNho3J4AmFW8GTCcOPAdBtit2o3xKIhe
p5bMXTNCj3ctnwKBpGAMIWVnw5RU8XI0J5R4KcnzPJDFKWBy+emiqNoDiPh1
y9OLIMkpIGzkGhJJEDibCHHyWlqL+3Hli2frAYAqWmY/e9Fm9roy+WA+0U6I
YlcrFf+SMwP7Kq6EccuMGDY+ApDLM5Oi2z/+1PxpH/Xnxv99HCUHIhSRRTF9
gJ5VYtNiJsub6ReorgE6KDeKjWK8wl7mDF4nmMFfTCPF6MbkBvfe4Hjg9G72
/ihsc9Z7Ogk5u3JY+kt+LIaTClOgCHk0PQ94cWs2UYO9ZBfqvcjoEX+ZDjdD
CSfG+UfOEIxA5/2yAftcO+vF5SU7Eii6RQOObWagby+8mmOcSfG1aSVC0PXS
2fPOES+4Gxi3OT5UlwRiJV5NQwrt9IwzmhCOdMMX1gRQD9cC6f+HxmgSCUHC
21Sqw3OQHcaU6gMRTxoCLxzla4FYWaPERdR4+lxPXXx4o69McaAqmJx9wMvX
14Jukeaa64dNsmFuzJ5FP1zg1PmMD43eD9S+LKGffpPwckq8uxTJPwAXP/uX
bC6eJTCe+ObO+xpi+LLCPG2BvOv/gj3uh6C+dHPB9NQtMuuW2uN3acFi6fz8
86HNpp1cDzmJCjaFo8EoCkui0eWkz0qWeoSN06sdGjidTsb79qDJV8ac2Evi
IkOUfeYVjrEJcRV/VXWBOqP99z88q0eJMbZVcA079+il684yQ5OTT9XL8klf
T9+gSEMuAoqh3RIqT9dqkqEWUTwcWetXEuooz1lwGyRmsd9z7fYDLCilvtH2
AG7HIt4TDevV++Zlxl1v1cM4GYEc4ekaxcq9QpVhY33GFjK2V76+WxQr4uHR
ua35Nkwdmn5oRDZ+dkytv3TNDr7VMMyZPfYySCj6HOawOVInOMFuAnD1Dz8K
hnM+7MP5sdsDSPsgrArh2G9lUElRtagscOJJGTSzRbFc1XKdzBx0MSjhpWn2
L4GCOc9otBa2RAamFkNIkg8IsavcA4B+L+Ox1tnHk5RWMNsRnCqkje5Gyztw
kMPKVO3OvGyuF2j9n6C9NcpCgn5Cp9K/1Pikr84jLryTQm8FNumMmmjGP3wO
fJ8uBHCKUO6ZJFG1yWmF7Xqxm5OqZ/qG05oCGeozx1g+JXeXp5c4UYAiVOkk
d9uwe3sCy1EvDNrRgYJvREEDxWh3c4QQR2ATx3V6fEIIYXMZitRoAgyjub4G
dd70HnQdJZ8Q6tdGeRml2bRCEM+fYwkf1VNlCo9n7q/iLeVVwAgE3X41vbNj
3xJC0kuq3+b5wRKJi9Ebl5tcgUvGelEwUrg0EzQbynTpOhLZMPo4YJfMjqBM
MBCP+2LigwQHWbRDNU+wgJgKm4iMmkG4Hu/7ozqkUB9niJSjLymkibmZGmhB
IVv/zIJQeHIM2cC1Z/piDyOiv4iGaOu/DI98VMqzyse2ADT1EelpmVRdiknd
KSVydIpWeZ9uZAp3yqWsq1SCGNie6kLHvu8TD1zNyQdNdNK/Hiv6dUfkqez7
QdKamQYH9bWNmhrbj2Rnq7kCWW42a1FVvITAMeiIf7K2j7hbMMg9d7qQSxCm
TJeXVIwv6OvgtFCxwep9C+6QeLrnoAoKmyE9D2ZS/JVwv7RhjjtekNrqnO2a
tYV1RUyQLirgn5lfmNXK4hWjk+axzmUhMXEqAGs0llRB7UH81dpbFwzIRGhA
EMmThoxcQPzv2TFYqu3YqaC0U90+Ry0rXLcJazogtq/MH3UM4QgR+fCJDvy9
JA4p2wEma+LTKCypHIFtABoa4BqqMiy5I+p/PM4d0lMCylwujRwrlO6/EOWU
C23KL49r9W+l2zGvBne/F/9FalK2PfAVCksihTI+iWVlkC1WFE8aqL5Gsh+M
qz9VsZ1b/yykLlPGEoq1wzqKHW7UhBGMWtBQHWkADk1iKHJ6/Gb70PbZwrFg
wfu6gDAkmmMuZ2hwjVtO7EMYjz+rvrmOILzVlFx8ElRgs9aN77/lZh8aFPP4
Hh48H4v3Rw8/5uIHfHOzWt9cuAgh6HM16assJPp2RB7bWvaSqKNVkgxyyjpf
1lqly7hr0zvSh/p0NORcoDsHbyxb4PaanfB8/Jf936nrP5CpIy24dDzB3JF7
kL8YSZtPLFlpjAaybxSfTW+SUnNVDW957mkdoyF8Y96sebHOrwh3Og5aLSMI
a34Qt9MNWT97Mvvq4rkhXlGHvSnz5FrH3a+e8MVLUNS2E5oeilbRaiT4rfGX
fZatffPxcnZf4gEKxj+bNkFFQoC0HYAnJ0YybYV/FYjy4RxlCpzSDaZAmPSQ
ftLUTgV7etRQJHKYQiX6gmUNthZBdOEIcE+GvtI3b8QOjpzfe0M4SgKc0+le
6Si9mABabVAKZmqGJR+5fsFpdzCmy32ZSzN+oP6J1KmTOYQXAOT8JcqfMe0z
McRmkbXJn2orZvHkGYsPR11+3+h04GIoIWsfIOXj6mrrM0X1F+fjH+9W5mnu
KbjDl87zlPDN8lAq52kKnGUzFUvQD3Dzlxtvn7YgbD7d4mTR4auRyxny/Z3f
y+1MvKVCOIfIjTBEpmPrEzBUixtToxc5a9+kILN1SwCXst2vuguwWJpQV8KR
egdcfid7jiwXpvgXL9sEuQFmQ34v5mTnly4oAJqUo41Pxyc/m1QdINlcWM0+
twrs3ilF13wiK7H7GCNOewxvS+SOfpigr/wSDFcRcgdNZfUoOAYnbhhdQDOz
YCXd+dCSpfFGXxy3nPfaE6Gt8wzPjCvPMl6cZ+M5v97UcemXx08UsIsKDsw4
6yiBNtDTrKQ3CNJu0kQUcBXfK1J/csSkGBci4JxJHbsmuOZGShkBRolDvaOx
e5dfRjmIeGTEfuo++q5gtuaBcr1PDlQ5bzxyk6z0edFaHiKpb/KPN61ArwQ3
8Q68QEkO+59zvCsTO5tfI/1+kOKRHMO35IKr+bTPm1PwHYo9iopRZoFJIaIK
IyAfiGh47JcGhX6Nh43+EHaY0KzHKVJXdBrM1pQ+Pm6xkH1w/JhK8rj3PQ+4
bDNcLFuW+N/nEwfQH2oT7V2ao4MC7nm7nKDE0/msJpbHlgbjVtRP1zHRm4Gu
NBGaRzROHCtH64Utv0AJo1P4ICQJc018hykHwVZGGMgDuo/DT4wlVbpehmvM
K7QWaqUx7dZWUFkZcvp3iDBN6OS0IibYS1X6B/TkHkpD2G2MqXohqIWFFvsi
xmQo2lz3mRGqW9RO125ogOwa7h8ieADYAMvQAUfQgkfmeOWytjdKsQ/MIX+L
GeH3LAr2DHdwjVdyNNZc7Hw9bgWGKD2O7mt8zb8QKhqZSFzj9HEGp/M/59Tn
7o5+0Ki6IIRQzLmHDHACgfP3RugjEuCNyJau+G5asoxDCs638/kIenb7WlBh
EwOEXyGwlGpb/Jpk8UgET4YsZoUhYoAqOn+KuJC0dB/L8yk/LhZO33vYfSGW
P4EFDRb3FiMxhoFO76ZTUbCkDbn1YRP7Sb94GzwZGvWtvYTvFEWTtORmUWbb
gh0aM2TxvNyPD6ySLeHlmdc37z9ZJqLkhmlpHPb0suRSwq4HVc0loWU1P+MN
Vwnm5WuokfUo/FKSoQO3NQsBy8Bh1Rn8pQ4Jcvoh68ldlaeAKt3CDgWyYrdn
KOSiyxo/BFbshKX2c0cjuEFc3gR0r+7v0xnyJDXu0poK2t3idD/ioBRH0rQF
UH/OrZMHwffnhjSQ/+Sgwc0/4WQjBlPG7NkuSNgs/+H5d4YQ2fmsWxK2JGPJ
ESr4sTjkFrkfGY3EVHGwCUB3hbcD9hH5vUUVKIK7yCwrxReDM/fpIl82yOcj
/ElWA23OeqNmyHppaHnn0ytcNBt08bBAsrXR0CGZKuIaUX3O/I/mHPpwkeLN
S78egaC7aBWw+F/IwdHroDCHBmmC8+ZVJ1Hs9ls7+jNmNFQTrhSI5qVZF9/A
n2aHNBQIs02APXXHLLSabtRXOHKbZWv98fcgDtYLEVfCFvVzT78ndxmdT6VD
JnCx2mn5X5MPzuayCrfmWcTIpyP9Mb/K/xNVlaXJDTXWMHOdCf7ANruTYZK0
sGkBANN+XEMxHBRGMMU8GI4WFpggqg8jT21H1ij+yyyYsudZECeZ5Ug/pj1j
dnOl7ixjm01U2iLks62aMV9sozh34QE1LkJea+23Erb+8WXX6dzZqm/1O7PL
WPOkVzYRdPvgVQdd6hWongg6iz2eLq7qpa8P1JA3W39PJc5g8B/DccOmUXHh
QkRPbFt80f175tiZH1V3dYt6Be3j71PNYMM+rmUCx5QROSPrAYUlwHyzDlyI
UY5kQbWRDOXqbOGK85Z5FFybnTxP9t2/yAwhDWzzopdr1OYHC/akxmx/c0EM
EHMfid5+neWJ5VG1ioqNzEtfWSrT69j996ns+VhtTUVdCqYeD6FQRIoVbxRa
UhbsiFqsseem3dMixGIe1g9SeLB6doG5yIB9JMT8g0+lE6yrIzUcrHonhRFO
ZQ+83BXv6lxAxXtYIwIxkD/IIOpFoXGTFxIGxU4nUDVlEghUpc5ilzPBumFl
N4ZAYRu5UxV635OWiphoDFHi8TR8OheuSOXx4zLUHs6hXKxFsKgDGox4FI/K
Brwp5ERFwxvLdiK6rbrtkLyLjRR7PARUunot0TrQYK26IOYlOUEQ/MURRxN2
raaQrWxQrldaDnBng49WkIuI0N7UHUfw2yKvIFrQEHa+6WH+HPEVqn/hz9vS
bhcmAD6wbICLgrLlfWlAp+Ql35dxwFCe4sD4nw15o7Ormw/yqqVbLqktAUJ9
1zLK3dnBCXkaNyY2xHC/KajWSdD2MvzEx7BL2GcMLgHZlwXfddCR+mzN9MCB
zUiKwCdv1loK7kt8UIP5oo6yv+DIZy3nfbDSFE1+vc1GC7Fy9L0Eh1bq3QsR
ZVwWQ7Grnq5rWbV7R7gHKHJFRNcwqo4x1WGudUxQk2D9S85ZUQl03vEJQio0
RHK8fgfmXw8OA8SXyNKdngd4rzsUVSgYsDIPzhD57vK1/AxcMTcDh5DDf0Ie
FA7mOPTD94NprHofgukJFFn3zg2gxQFFJjek58Lt0Es3YncIRudQFYktzVR7
rgj85+/ZFFfLAEwgi0Yq6IRHTeAEQ75olqMbcWTuJAd86xw3VLyFwJHYxkz8
UXT4tsBQY1BaZCwesXTaqUEZFE3zO7D5Q0B0H5qLnKjmKvkJAJ1m0v9H9I9/
oDG7BLOP/pAXCvRcBvZgEQKQAb7yc5plZcRi/Jru/Gw1aszY8m6DD60Fg2Kd
+Y1kTqp2RM0C9k3GCmKnJ5floDb2uHYrj97OfqjDILhCCvlinXLaTgvjZhY3
vxZp7gRRvVO0QyzYNveZ3tjnEw0QzQP9hmxusc9dYOSoBICX4XQxt85eHoYv
RusPjVE6hX0YHP2ATsEzWrgDrSaw9KFfy/jjudS4mXhp7aYW1nWlhJJOGtdP
OGm4N7E0NTMSyVY5eUmyvszWv4vetPUP8Kl9x0L7FGu/58Gyveh3IJkXjXyH
rY9oJBtd6rRWASxPVveBwMrEtxXf/nBxEojVJalk9XmQ3ogOzzSYR4S1kq2v
x00cfrxB9iSr/ecUO8BVFpPKFbplqklzR4JXIIwkjb0EANaVi8n12TmWVXkA
yaFzWdFWpmhZ1kb5HfDZlUe+7UPslUjRTPgmiHubjyFaLC7Er6bxmArvEIvi
lYgeDdF2T7bH54zKr94FBvaRPSadcYbM5KKBnTDtWf72eP96etl4vW5yXjty
P/QnUYvwCnD01IzBFz4NCqZOuUcUoYoKFXy/mVggWsQoAXjdRz/YZKHtglix
IEaGxb3o93T3xVFn0ZMXVJ2frKe1laalRcjJ7ODHMGMLsvhon4ZSk4K8kdVA
cKSWj37zaOUtYizJ2iBIrC5eMCOCdjpjpETuOrRuV68yJWhYNZraght7Ii8d
cHSrrwVqUI+SK9Xv/EzGzPzNsWd4Yyslz+24JFIVc08P7QQ/NtraVp7Ru/lK
0drUPhHp9JCUNUXULWNFxuZHxElG7CxO0vBSKjK8mdLIOUMiV49E+6OzhQaM
cmrzlJ5COoaWQVprra0GH0qgBoP171rz3nzR8WnqJN0YJiwQE/55L281Ogvt
0RnQjwKUqCUYZrz4VF8IHblsQDSBre33g5AK7BCtM0pqS1RxLcYLL/M7DL4J
YW/AP7MXfkxLWDO4n5PIP5JQjmfm/+kT+NcOewo7eCmNnRKaNCzUOFFnlE1u
hXzPVjompNNGdRe7zVWoWirUeFFuztQEAHz6R+5r2zt3r+A97X4Z0PPl2c5o
jLkPAl1atcdz47JDm9LHW3aeNLRfgfMrO2YQwJDUJGpIjOgTqjlDaYJa+4tq
X0pc/GmRwX+/smFmspL+jinQZF36xTHV/P9bMNtKgsNr2w0CZoArMBnm6fXT
Cs3HsY52lNuq8rW1iNM3JB08bKVJsKHnFrYNlJbKy2ChcaJ/rRH2nrj8Dz+E
mH2QfpZAlDCrRS53rSk1NBQd1CfkL18/1NN2ERpQWuQ8Ca1B4cG982wnD27n
fL8sYquxXBljsySA4BHcFK0+dNXSoS9hNP4jHEMT+E4E3sTU08Gfro187hpr
EQ+WwJTcQiR04iozgQTDO1Rl6sXuek9XOVYwvLx7RkOcCx14nKtBGNIEddMD
PQ3TsrHVhw28GqNRgAayQR3XnKjBNjOdMn/Fr1S0uLOa1mg5N163YHn/E9xc
iTxlRl0xSjUHYQKlbM01c9tNX03iFTlw4A4PIxHmErkWwshpju4wzwTFEdQR
hxqcf4YMbwo296LokKZ9IshD7ichOSc2b9CXaQ4Bt3sx+7gj0XZqkZojrxTx
QC8DmLUrFR3mFSasDdbsDmUBhC0mDCrf952xobmLZpgVHVOFJ6L66h5goVWF
6tkTbnK6nxoYUeKNn+xozi8ii0nT2q6Cb/+PdGAOW0K5pReYY/utov6sWEgu
NkUPPTuL/TKmhY0zdwtPX10k1jx/gtcgknfN8yIHvqICviJf9DZgHAhFqZVG
ufkMzCcq8EUFeZC3hrU1rmuETnoLhqrBp+KxD9IND5U6p3xfX4VKLMpZ2vdY
obl3lPmmd+eGl63Zph9BLrcAHY+TJoAngRTODv99yRavW+gXNSqCFMpVng4e
A1NCG3nw8JzNhbLfbvitxOpMI/ZLP+1CMicx0iJhn22Mfq5IkYs/c23cCM2X
GlL/Z+fwy2mEMtKA1jIxsktAuZEuSPRwf5lKNiMna3oFU22kldcbjQnYRspg
+o6DfjYX5FvHMgaZLdkCh8jqs+1g03TqmuzDpmQ4ydHwHZi0NpuYzcsxnJ1W
HHFS0nWWT+JD5dm/eL7DIq1OV7VpyZOLxDwCWPeL26gvyaZ65y7f3VmKnFam
UyJvRM+tyS4BmhIiUZtzvVejC8a01SnBSm8+9uwFtcnq74Jo+hV92sPEsZrO
Q8lkqkANaaUjrqybjy9NDTdAyUddkhQuBfpf0nqe0Y3pKUQF1UJ27TUy6jR4
kzyV09xVUDoi16wKA9CifTwCBfpelY8CdNZOjJdeeCTjqSv8zjAx0MxbXhdc
wwd/WFN05/RajmtMeoVPs+MjQXq0flZw50e5YRHaO2aLYblM7TCfo0IvOz0u
j4zllfJBqmIgoM1EAM41sV86wTLd451J6mbbeDsS9Iqb1WLpgGPMstXquluh
p0jt66onWrlzyo/yN5Te5dSl5GDPQ4y0hZ8eL+no2aT93vQ+4CFujosTNqxJ
VaWpABzARX4ETJakuMcpWDesA8Y8tSp3ycJLZqjuTUPxmU6lKF7mwJHBydEb
q40RP+eAnP8KtxETaun7Y6IUKdL1H4/R0YDKMd1AFLparlSx9qnLwVVXQ+HR
KimNXGBRozVXn9IZi9NVtt3NsxrRkKOysLgm38u0UuOSS5Z0bw0e06HN5TU1
X5RMFMQsoLUAlK7dQCkvv1pJaAPVCxyCEnBjP7+9uB//hoe5jgp08luws85H
CamvESLALnc2Im0w6rtEKQShnbWGoq8SaHCAy7XoBjcCJ0aZDQBs2vDaGNQM
wQ1V0wT8IZkUVzy/LyG21g1446gU2F9sCpiJQHr8A54i2jDbFBt0d9bGcX0f
ed2PkmfiRUK4s5LTEotmmWulqd44Joo58XczWbg6xtAybWOj8Ci0A4OE7tR9
YaS2e2EYgsePzzHghuH3KFkF3xKhVvIBZkUGd0IYYDuERrbhRq3B7thi0wCJ
l7cwFpGqivd5NmtF1uDnIOJgIrWHbZ6+YVTgaf6aPE6a1vruMD6Ca9y4YCgq
cuI0mE49cwyz358//RZzfimsaCX2aIdSn38ryhrs5vqX46UcU5FvNOmQ+J+9
OA6h8fIxmAH1zHd6SxBu0MYsICXrwlN3ZX8V3Y1M1thxpPR6TNRcR63JNuj+
QUhqzJA0rCNh9gy5yqRtUhbURYjPJc1fZQUJY3caJXbpuuNhYd1MApZUOeRy
39L9LNjZC2AA+T7X0NDLj/08wFMinrfOI/ndy9WBX0GjhOt+eoj6Dg0yRAGU
Amvs8olYFI2gkDY3/tMDD3U4M6dmFjQAXHxNgAxUoH+IXmjzegPL2y3SmwIi
EB+f5Jq0ttvDt+nMYk6LAbrV/d5K7zi0gDmGolAHsPhTE3/670M2D/RjygC9
/i20gjlFFYBHttKv615OhEAFNSEABMdeFJe2q6ZA/KiS3oDZNC1DwNhI9ISA
j3wYYn9CKxjV2tDxjdOZ9nt3bTrmCrvJL4ZxML+l2TIobhaiRTN4XbA9ym/K
8HwuFTe5h7fcbvof7+Oqe8RMYrUc15FSYTyEcZuesFPiGKM3mF3dYkZwJCd+
yUeAkI3bemxEqN3i61E4UjN0hpRa/QU5fJJCKCXC16ZDEgF52QWv3FDEvmjG
s3yTGjoXJJ/3j2xXv3f/U0G84SidngwI8Kli3EpIiO5NSWbcCEVV9voYdJVW
gPbO7C//9ik4izwYVTG+i6cW2N+0O9/GP+YMjy9bmH3teabl7j/Wi4JlUnGB
4nWAu5y8mTPXvzTIn0VnNBWxNZpQSTfoTaNZBLGrYUpJaDWOduEPp4FOpnUV
Ynhb+jO6tVv/HngkhqBLXXTmQwfHTxUMG1+tt/dCUiYmhOS7pgm7XaaE6MRe
EM66aiCbeCAUx3KLnb2ubxcJN9SkSDKT5Lhlzwdse2ML527ecbmUV5W4GYJ+
f1mWVZdwUfVJmjkqyrZhB/DeuyI/DFmrKnbfYFgzxsni9YG5llmB0/weFo1q
ImmKjT2Wk+W2fs/BZZqfowXsdKnds72wIyxRvS7A9c7obJe3Np2gitp1tAL+
uyUv+PfpUTyuT+IyjLsKEnzJKDP+ZnJrYhUu+8sdFgcpOwyofe9rIbz6+xpO
qwnAFrV0qqdp+Plthp32dS1ydKRlNDUpyBXNl4CszVE9mOJSClr7NVWYTFmI
I8meuqaY5oIgY/EbUL4uUAEGxTyYeF/PcZU8tmUj0IOewcI5OUhl+QKpyuMq
1gtLOxTc1mHjbAV4U8oJzYPDkHhBqwPVfWbNi0uezcL2UsoXGpQkGEJwOIoi
UubcmDiFmaLyXqY+3XdrtKCEL5FD+7988eRQRdNw3MFKxMpLcp0R9yXRHBHv
Fjbth6R03h5aS4RIMGNulwVrkh8PjD0CNaE/LzDNCscfWJdyqBSzq0KxHUnk
UrTc9xq73lEMey+90PzqsmUk6BAsgsS9jqQSj2N1jEhDl2D1r9Qu/e0HK6Y5
hRLcSXr/bc+8UwHKKxjOjqiOJT8iQQHekh124fMFgjbDH1kFLdM3EEOeJA7N
4N/Atip78jUwWxxHzFpYQ5rvsf4QyvcvUpODg0wqgxOCUtBwZHpBXVHSU1U3
SusL5kQ7yT+xK8Fv+p3uPvU3wdWpl24h/EsXI8lJtXwK7aUNGuh4Wr4HZOd8
QxfE7RSkWG9izWIrqrmhiwNPom8rU+zfmOW0NcsNKiMkj36Pm+7E+zr6mvcZ
zqWOsKxGj7/5HHYBgdI7aN94U30NADcqQAeoen+JDel8gPDSL1C9vj+UIg4o
GvDkbVd8JKzeQ1KEVU6XCoqLXpKxEu0oLyp3YNl+0v2Ake1xQF3LeTCwhsee
uPCmpNlzIsIhlgE9ISXO11MD978sfs837eXx7HJPACgUSOWLGHEC5LKVErhe
PPa8g/HNSXf6M9mOCkeOMcodnVjdiSOxBJmcUdVHOylRJJTw49jhVHgEoVGA
lJeeGBAfPNGWBqcfUGINqgyDFOx8d9gGb9sFp5QCEG3mQG2f9vedfErJTeFC
39icXIHz9DvuyhO+U8PafKpttxwgNwIV37S+ghth3NCfm0rqJTUzWt/lw2pg
oQFXd+fEZnbhrpA8xXhzgW2b69+yHFq18ezxVhGol4oufgJ7InnUvnwKtIZJ
HMseS0oketXTAfbQsWwohyNkb7ZGijU833sKQyflfzC+TZyWErjqGafLwa1O
k8L+FuS+HBpqsjX5r+c/pGgJdvijgdICPL2DHJUprpolUCZpMUhWYL3TR7gZ
uPI5hINdUV9C8mLq+3NMo/hbjziRIJoHfdBfQPNgzTJSR/z2/ikT4QmwXM9F
5ypfejQQplqlNr0BlU2DMXYpW5EhRSTJz0/Hjfvm+GlbdyxA45SB9jlFIL9Q
MB4ivNuLKDQBHw7bBojbvFW63tZS80s2wWD3kRasPu8E7dHZ+DjmT6cppJpV
zSgqDaaom8rEOfd446ykO4p7beGbbNZAilUo3Bpb5IVdP3hq1sY9MilB8UHL
Cp1lWdpZFmGzF9yfGGOYhvrJQVWWeDikjVGuX6h3fhRUoZFsb9vq+WZIFLpY
BYqPzpOHY6FNkSU26MSG0ek9W0juzWQ2PUbnmZgaJwwJOQUYM2MTdpvXcxhb
JsKc6DB6Rfd07S8JOsBe5DyseJmOFOwsDymZBnASycPxXaiUGCmPuW01Etgz
0Q+YnZbeH8HGfgmNtlJFdxeTtROEE3heV7D3mRyPZv7qgOVpK5LJKUA9VwS5
MNXvos/v+qR3ng/4njPpipLincjXfUvlGGU8jLfNhx3SHsJoaaXKMr8A2GAs
DDKLCbUc41aljyLFHL7R+R35zkRWzsMc6JqCK7cKw42lR4xbS3SRDAEzmgE7
qmNfEGi9N1fdj6MmRBopxjup6X+XaaoyScAPWlyqVQTQKFDKZeqE0bOWvqsb
CoQBkfmEFWtpvWpv5NEzb9UDXhx+82AQpxIMx4RiWHH/CJweYUAke6yzXM0t
e/qS4t7VLB1k5Znh6xpwZgKtCgodlwPX5fRX6EJFkS/fv3B1YPhNX0aEEC67
+dlLIbm4cc+CCI4QgqSnKWwGvuRnmqi1sdFh0IUmvenuu0rCUn15gPQNrdYQ
h1d3Sl+j/uQ+AYUCOA+oi52bHQj4os+JNW8BMW2pHDnWjcIQ0dZCUSxkpeQ5
zEO5ccv0A/3wg7eBNbRV9O3UzBWu5j8e4ef6dGAgZ6IGzfm7MMks/UTvECAZ
14uwVngt4tHvbj2y+0D8ARtRLDsNH+bSG4BkEJfILeOWJOhKtK+oTsKhFfnI
WjpIiGYS1gBkNOSkZwhOVpkbvt6MZS50TWvSCON/uDszJbWyhWwfvZGvVNXb
jpyELRXUKV5rjpssJUyJomuJ4TDHo2bYNlQUVcGktqpoPz3XXpFZE973PBWO
PPBuzRQq6ybLU2OL360N6R+4LUy86c4w4XmX9Lz/3Ic5O3OpqnSRWWIpr0MZ
oQHW0rMLgvpY+BwA8C4REJK+3uK1e8pSfqvxli5rTGkgX5uQCLOiIsFCkymW
HOxZTuDejIq7gCTUwssR6vJVJfa1FK862iF526kVZZO2S33NADeCsRL26HqK
DbNn8TAyxALb7h5SoKoNgMP/2EN0rNuZ+GDmfNcONxztBp3/1VrlLofAI71S
J840Xv6UZWM5E7QB9/tfsSeM79ve7WFB4D0T9mPS6ovd6OwF6gcCUjLAby+0
Qs6nIE4vOjAkGqdKCeHCT5M79tBNA8LbRcKkbS40aa48HO3NGYnqkz3F4UdI
f/uSv4wJ6oCHfn9ThLf5Ss5SiQjat8PoG9ztM/BFHhbBrfvSRLt77eGii3NS
VDdaIbDMdfVzGhIF0oW6mw8p80+hJqrF/9eoy8zDUif3p6UZ1PsTwF2/+itt
r3vkd3mRx5yOLS8hCC+/G+bq8iruEt+8oZ+2If5WGXC/xP05S352xcM8Myp9
T+f2adoGe7/XgrYBOs7ZreIR/LCg5QKBA4U1JnfYx4F4y1dL+tzz8oMw2mQB
XhJIx/5KGn8I6FffyUT52cgJxhIfUilLFQllhEWskXAGUNKiEEfYLq1oJNNl
LJR37QU7vReXxbhNzXDVDsK3Awf764D7mKrHOG6vaGRUuqVpDB7jLI5FRegG
1RLSQhL4Wb7sLUVsyHlmCeAKaBZ6Qj4uIT3Lnm54SNN9yL/6HYCzDufRxPci
02SAHExgypoq5QWfSwBhEXrjYBWAzjE1jgsBIjaglUF5MGaHWlXxqt4xSg9k
oti1Wr9U3pN+aX8klnnD7j/bczSDCTDvtz4kJLbJNN6kxnjLpkXgL5kGwd8I
kJT74SixAbegQ5seRoNMzkC59iJybordBsG4gPCPw9/dV+/sna1kG3xNrgzY
+8oBHjQJ00RYspuEDlszIJOMSCxUYAKWIeJpVQ8d2vtaHfaNFsdsMFvvWxyB
Yrrb5xqEVLF+8RZLt2RB26hMV9oFeUNuj+yjJ6iSSv1dDTYTw3+cdsqtm14Y
N9GDFMkcXP8bAccjThMr5Y0TTMjiOuxgtoE3bNVLBwjFxgFkOZHGwh2gzAoe
NFRfCGZe+d+A/ckBC9/w7NIQ0/6lHnJcrrQZHKGn0NStRavCsbHACQvjOAtQ
qKvFv2+teu2ZsnnSospQk9tywMmN0WnULWdJoIyf3btwbejSeNByKtLf87HI
i2vomSA3+VZe2Di2p1IATozQDEW8Udz0hEVIs/0rg09aUy2kouXuizr0i2Py
+9e+16tSGGqKigJq14zpc/zI89aqtQpkw79FB/z/geUNTaU61VBquuEcgl8d
tS6Fikjd+JBJlemumK3gC+cT1JV8kFWSqDdjk55dLhmOWu5kh0MUGUhM1W8Z
570mmJXYnr5KFP9vl7wj12pn8fChan0G6rv/BaAQvW2wZGRXd+ErXgpH0dEw
noYm/eJY0mzlMVpJkAu5jBKWH2N0jI1e/7stvTzxi9KlMjz7DN/4JkVaxvYO
KTipuykgDL0k6T4KBzRa9mRVMyRGAgIJn7QO24qruce+AWzp2HOUQzJesYoB
WHtmFE2/kIH0xmBwvCOGRg9EATBHIIU4+T85A7TYSHTVZY1LJEvOoNQyq647
p2jeT+I0fhWMYNBWkHQibOBd2BvfxASy+cVwA2T3atXHtJdZkJb2xTBOaKKz
Z6HVf0DPPPyxKFeww57gyl05SOg+kNJLAhbj0qg+YZLHi5QeYJdDzNkAM34B
vzCEn0nPqJKpUAZzveIBao0S7dehw95osaKGhMTgp81buL/w1bQDu+eeol4r
Xuo1iBEgRrE+LdWE5/n5nOrXhYJvx7K4Ed5Xrfqc8SOZMvduEY41Vv4jdL/W
AcxKXXphV7KYTmqPpQUSm3QqOIQoFl6vjiwWSu72KkMHAo0ih7BYfsUiz/8k
8skAOwRYFBAIV3TGVUAKnc4tqn0AhS0IUSXuITOO39g78fdbir1ucDueFkvF
kAFcWuSmvwoI916WyddzraoGjH5NlWjFj9J63ajWiFnAbU0FA/2tCpglLy83
rIuSoLNNrfmwzL1goxcUBhBJvCsvGeV4o6aZm8PCrxHWm1/EtL/u8Su6JWxh
a+A6yaumXPhXJ1qj6eREVi8kGdh47pzPEdpXQ6YI+rTIuTWJ+3sf8qvCiN4j
sDcvk4rwPSWxPCdnUanbn1fLAVdYWNTGRzyG4t5Vi1DtL25gb0zd9KTWyGfI
ZZy8+nP4HJNk1k4kfI4PchI4/Vx7FuDP2aH4MDQzOhsEFlCUEzDJY8jGx1Y3
1qxfUuVLGiTse3UJa3k5PaZopGc001kL4FkXRCYHJndCvjXF7s6TdpN81Gpx
31FroKJPIMSOcbr7R9MMKz7UvhM7ac8tAKceaEBv++nLdbKefsz0u05fNB7g
1lUkfFPr6ifsGkCXXiBhDo9X3V2rU8jnPq8UqC1+0yOwoDoRhQe/VCPT+YqG
4E1sIHvv/PMo3F+/tdkN/cxDyxRbDlRzjkkRMlzAHSYAx2sjYDBVX5rLJVtS
83pZjTbcV3H+PLgcmSYfTT6SAtZcrbYUJ/cXkUDuADAIj8QMqTt4OrecujO1
OWji/unqsq5T7M5w3fbzAynE+PZA2I275LEz7FXgT76ggvmNZPK6KOBUcpZ4
mEvJBcfeFMhgL2oGEZtqYvahQF/ygBycUjaAR+3vS3zEacgcX1jovP5D7Kia
sSxDHXBNCOL+6dlJXAhns7uJv0cLBOyJHpkseVu3IJ3PRHjh+wf0+jpXJLoS
Yrw8bMqBx2rgmiykzi9f6zKvPbZdggNWLlc9XJ8NtSuC23QisZR6AB1xlqUo
laoO2qBhAGnzrnVG/3GYHxKcEtMdYj/WXj6hKUWqa1yCQukjYifhPuXkfAve
8vqvrtxeCzlgmEvJYiUCDNC8368y920CUDkPRwFpfmAyEcSyoca6W/35m98L
NFpgoHm8NFhajqs4GdecoepLRKXcuEWpa6kmIUnvspJIJMvbrkXiYB0S7WQy
F8VfTzzQG4WFdtEALTxvkxJVgC32tefdeDS8tgyA/o37Yg7P3VMtsgOwcrDZ
A+WhUbhY0maAAIDb810I5cANxQyDsRzKrBKQ3XZpWvAy+HdK76Xd2ZjgSjqK
bJcBieQBVwbU9VwiamCV1IQv0WaeWjI2eRTnLTFEGYIhzzas9aRQSvs1Ao2G
ia0Mz6MQvVw3GE3b2DVzu5bxr6ywChitGMBMLOHiRZPCEiJFYGbaMV0/mO0c
lg9nfw9B40fsYhWh7PkW7Ydelu+gV2Faxow1oVuMl97BXpe7jGcLcQAGHbif
R6Ivr26Da+H8GyxVOlENr007bHtL6OFpSLw6hBICkGmt1g0nDD3YpM5cQkJ9
XnNDcCDnNthK2oXtYpH8tYPHioM4SwuGg9OO0GsYEE7Zz++Fq4OU0kesWHMm
IajIYhfDCz+62IwSm3cBjXOuGB3WB3G3rswYqZR1Rzhfop56iEhQpv6HoVz2
hM1y4S3tIghNYKc8xtT0+EBQhYS56XkrAzAEog7m94OWxBbO6NSuy+Bgxq1L
LoM0ZMSawwx3AldOlhRZxzErODcIHz0vIUpgnlVORp2W4+xZQwZbsGsmselX
6k5SMljGOBsjXkYfsVrS86NX3Tl+MeQlzReZquS94loI/lYeltQ7eF8Rn7tH
chLzI30t+ZM+xSZx+zBUksldG0gXda+TaiiShzsd9EsK/i3u2yjSyrP8I+TR
/5Z9T13kg2TKgrfdt7GSg7LXHdQ0nKf1nzwEjkqMxGyNhzJndQuL/M4p+M7y
EboKEBw77rCK8oo7E/QBj2ierpphLPhVdzcejyq5InShlYjEpC0ioZyI7uJi
3NbVB0CHFdf4U97HZZ88y1RR2RhDZtL4utNUw8OpfAmpx19Enx/sg3nMWwHF
ftfMIQQHkoSTNM/D8Cr1g8dC6M0sXLbV6wKUeTHaubRa0sb7MQr90MdKWjP/
bLHX1rbCqW7b7hs0dVge0Hq8SKSQmL3f04BzT0jSSYjLb9WzIWkcp3wZwpeP
qR6npfASL40Q2uk32xi6xKXwuHGP8D4egBNcGFwS3vV1u1W76Uzzy0/vOEjN
xKC0nUnDcAkUzLH3pV+PiI3JKnT41n1BsSvtXGB13IBH+wUfrzy7hAJbLPzO
eUDl61JksAKZFxjLfNjtx2f/Aumo1GYNYq42ImzWh1y7NaWvGYwz6CVC8/73
n28v7igeVzuCtHQCGu0RQRPW/5c/MC6EmYzxTy/NeDGmF+VuBGw0lQ4uuqks
FQxrSrLAS4HDAnNg4m1eyVfd5Vv/kt1cFPMHsBqN38uFiRgHnkeUOG6k2+Yb
JeaDNCCAc/8ngzqPtQazkzIjqH0TwyAQvk+zNFbs70oapRYNSGcN6a6eJ4Hy
VrOy4dHCoJW0020FgMOquiqYx5ojZh3kyyDILehZRtG/CRtkJ8xDM6bsUbbZ
E7vfQF0m5jPgme/KMgNb/O7FCmilivPZHJss6VOTOulZXaQFgHj3szbQvL58
kDpdUmbt7SdJHMPiosoRgtf5DBHhlqcFACOFOMFjpJoMA+eNhnRp9J97xToA
NA9Xrh7g5LmR+qBxEpvqDWUsdOqiocjP8ZX9lzAYSA3ZfICGnuvAUp3Sq3ob
637wA1oO7fCykmq7lkQFBzhN9wKg7abKqZx0MqH776cp6BeO5GH7Xt8l5Ysc
GzQqwAx2N4zf9og/EId/M4QvXk9V/MeQjiCbIYCCDpLjOPKv1ef1+pn1KzQb
g2nOjSKd5dgLS8B9qIFwcO9VZtimK56l+Jnv5b06C985N1M3s/BzHaE7sSQd
n/6uMoefGrKy41jV9qWAoNDznKxLJbnpf/PdybBlG3co2t3BrDA3ZGUts3qi
FGAfQw00Meh/2+rBLu63no01tF18EAs/8G0372FuzNi1cA885zEP0FQnLpT3
G3GBaeSvitW3IjCniHFBZbyDZkEXDlhEVxdyeOoqk3Pv77kamUZWyriZJZym
MDPuSAfuQgZbfgVhQsQOeXy9Cu+urGpNvexEAyHa9IYgcOG2SW2Xrr6twiW2
+dtjQxMhJV/bUhxj8eN5Fz2Qcjf1/KQL1HEVuwbPJQR0a/OcG5UblMnKldcS
PJ9l+RpbzT+9A/pzbgB8291RFKjpgrLJeNLuLi92WNmTc4CToVOHl6L8/Ko5
E7kwZfeaGrBYSHfOTySAUx0ga49l+YQUcdxhU+LHKIebSUwKoPjFE/sR2z15
6++eB2NEfE5FMlzGPoqR+sQGmhPU7p5YouL0F+x5HKwL9uXmB7dlT+J+DuGh
v0bHL4C8GOy4yiD5pjbXzwYOHixE1CIH8ZEhfNeQK+GHiOKDG8rf84K7mkvg
G4SUI9txpfmCrORepthJLuDqTijvb+Pcv7ACJWWg6Wb5qheCxGMuuov3iGaG
cm/Jolp5vvN5NUqOO9vVrPlDgJbETJnwfu0StPEkcvlcHiOweqdFqmjabt1w
vhL4Dxard0hew8gaWtosPl10U2MTY4aoYlSGRzeRz5JowCbj5q1Sk5aPC2RB
ZDD8/+PZhgi+Neu70pYK9geHtQSsh3uldxa8hsWgi/X3fpxAXxDLBz+YcXwc
0HXQ5U6BIu6qeqIxUICnS6CnMTh6SRzK1EzSPST9kyUd5co1eN7+zyqUYF9i
P7DFZcmC/0SvDOEgRma6va3cTANICN1vn6wIBCGzS/rt4KQdVVplrFsX/j5m
Srws42MzPYYBGwfbngFpLUQzV863xLTlprY+Kgy+pNLRyfq7WNzM6AWDwfj9
0Fdac1tXF2v6AznBelM5tnZotRdOer7h56zk2lOhUjh5pE5XAb4iPApmUQC5
JpFD8+DNzxY/fQWEDYZNwpSgyw/2Brf8kJWa0xgDpTIX8iWQ/DHnGyI7rpvi
XuWoJjz7D0MzdPCBI/EEXCl9BvhcOQcEb+ELfCBBY6jLzcVCz63F4YYm9x+f
QZBc4XusDLjxBUvDSSdj+NmC2P7+1TtZetOcYSxUQOp4WHU1B3a6fm5BUaPD
5vyW7/4GouwDoXUCY5UFmLy+Yyuc/DK8cMsMyphEcMHaSaLwzLHKq4g4QyiN
tdqgUrqob4FiJzWVSXSM8kYCrSLtV5UrqWhjetqLY3HQLQSHo1BP6kEMD2P/
G/U7kt74BpnXZ7p/XCCmMZ23yv+U7m5kzopMilSAXghvWdQzI0Frq9XhwxwD
tq4lyUsoHmvieGSJMtgRnHW7neWecGqnfMEKvN5UUG7LErdpiakFnLrxQFVV
CrY6WNHTrP1O6qvbJhc0VViZiaxPttW+XdVN+xJoeovxryxWUxKehu8dvasT
mpkh53WjaKN0hvPYotzbUgd/QgOcUW7dmmMAtM3MDjJ195WS98xdchgsTshR
Y6QXxO6bVaoa5Y1pRTTwePrxt5qlQmbNkCRB+e68ZKXyj+X0xZGYswizJZPN
7EhR+tF3zdE0zYBc/xuMbXgN84/dg3AnGKmYozInAGwGhH1pWY1ewGDns5bS
2hrZA2WCxnEUC6H5q+HPMiXAMD2qlhxvGDtvtlTq+R7FJwBjzgh1mg5MZO3v
e3eO7kGRDAZwCNPDm6/C2UjsURf0Q2uxvhM7kZT01kzEkj7FT0ERrtaZXAqL
LMS3hdfWMUWwMR3RkL6a3K2gN9K75hNeOJzqxG8SPqNwsrPeXtJq2EJ1WgyE
vWNZLU09DYVbPUy5Vw6uQ83M395fKwQ04Xbp5HjEEGG5hkyk3ZsGvUKPNi4J
e2h/soYoaqasyDY2tqb1qoeJUTXiXme/TFKVRwizTCQLiKXzXh7C1S74ogIh
HQHhPqrjuKLjE4J+7c7sCTDtpcEO4v0LrAJBdyOZqmXKbko/MWuRUjmNg22Z
M94VasuVf8mrtGcHr2S/dPMAMH3xKtb4uW0Dw8FL1BEYVQHlS7qQRLSFQyKG
TW5Us8k5yviCNh2wVrlAMhVTcQCGV8AucmYzQwSIxDENWZl0iMrtwz8+THiF
tiSUoAUA4DC6MnF3cjd+GpGfxpMZxVLJAdDS2ChHO/DIKtSauwjkhARQh3eV
eDdanrdexbfNO1henr7XwJ3hnd3aXHAOykLZO1DIXf8yWFL3lmkrGhfjVR0X
q4qvmJHqPBrqv4W8xaw33YrmhsoctzGQu+I4mXwA88sw3XKLic8/ml4h8TMo
mjYvidYILjdxZE6wS0ajRBGixkO+TOsWBtiazkBtepauDO+r1lqxuR0IUaOs
2fd1ICbWjZdAXtXw/wMNWZWfs/zDdiM8lq0SFR1FT8QYs7pR6gf1irqplmkZ
+Fqql99n/OmXwyp/SXQdQjvPB0M3VrL/EQjS/UTEaQRqhQxHZgjPwir64w0H
Q8h0vxpFFdT2A45ImsLSBbH7n81QA0nVwS6O/iIuRbKMC6EydqamSjf9xC7c
7Wr+PE/eEH/2KqhY+Oj4QBxgfaZ9pDoJy7yholnXvpw6drctzMMdYwaTVO/a
CApiSAVtm+ueiDTCGpNm+RQT4RCxOESU3GWN7Rvbt5B1Ffrs/ZFrukN+/pbv
68fGU/GJlyPGQZ/P9YG9+S6sPvX68sWKyzmU0fClSvxBAJKC+lhnbBXS8SyN
Cx5Ee6UaB4Krwx3qeO4XNzNyyVc/wgD4DtwKvKFjqYEDG+6VMuz81+Hac3Ep
T9xox4K13xxC4nIyoiedyxpIbtHpcFX7HjOlJD6b5WI+TJMhUbPUBf09YAT8
AAPPDhlOqI4SJ42DGdvMTLWiLzFs8pzo1zwbaAr8OymaHHFdS7uh9IKaO4V4
4r4Cmi6f1cUP4dq6i/r2cQIu93/2/zAhf5YOmaEksd0/QmMOH4645T0K5q1p
3YzF3o34BlAfRRPyXcHAPHVSDjHu73SHF49T8+ZwT33dM0duORrTTcbL+2EN
6bW7Os2PseaHEMW142g+dVZdAeAMrSkCVh3vg6pT4ue5Aga0VRfStseuRFuM
17UmpD89R2wv+/KVw43qvDPCfQQ4kWZaKbh7KvQiZDbXsFxwFIPmEll9g9o0
lsV/3cxV/wdSnfEr2Z0DWYljueyl6jRx6TOLqos77LHW4Y5OHl56kcs/KXT1
buEPFJzSX6i6BZhGOJ/kojF4n1n+UD056qvi+5e7rhwUmgsWvsgMnaViYhW2
uBuEB8xQu4KY8xAM4cKGhJgSIJSrctXU4kRubgsk1ZapVBFPgm5pwlCyTIpY
77XuBL1bhPiTrQQvEOa/CJKU3VYXD+2TYbrzjPGP7rZCjVmdJn9T/onsL7xp
SbRJt/K5ZwVuM8Asy8EtioS60LzPdz8TDlq/Ioy6rG+czpaT/bF9HYT6rNTv
jZBd0E8PIdMTxxYsrJKrw4emnWlgmMU8J7Sve26elP8HeGvRHE/L0CFwg2Jr
SktmngEDP6d/6TWbaG489xdnzXopET0iu57zK+5cD4R3j0RV7NswTu9+Ncr9
R7VIGaVJ+gLZwKEdlp9V9yQFOFHOcIkHr2+nXD0470uHJJQlg9PvimRLTrzC
r9kMTiSdjlFJZIdKEVGsvJXzDcHIIxVxGjCgaCLeuwq2bJ0RJpRIcD+Nk0LJ
lXf4Q2gevG3ihirBgYY2b+yBbcilEfcdx1mTRml8Z4CKwmrdYgUY0MLVNCBd
/qEUuUZMLzaVbnGiHijWop2mGnDvQ/jmfQ/4EmqEtOq7s7G95jiPkT6qqsOm
hyZ1SgQXcVpmm/NNY4+dVsueGXLGXxrBPP/b0TUns3re2QHpFPxXKrW5QDU9
J/BpoPXP838R1M3oax21ws11yWlN1h5SWCeZI2pxy8ID19tcTfCnXd7/Xn7c
pepQBZghxoFfPVgb+m70DDTB8Lu/BkneLLs2luiBXiFcbjVKaFZSG7VGFDfk
qUcay1hqh972dlsaDVn7jbMBt/KuYhuc6i/hWBbxOFCpm8kEQvlUjZzRPM6j
m7J7rpxm3H9WuV9BfL82+AftYv37YorjZkiOGLsYxZD2qQRLU7uqjHEHUh9g
SDhoPhAHqplNNbRguMJDeo11DnCPw/bYzQPXtqiWfOUmUZpxtMLR3WsYFc6B
S9QA47vJ075cCpy0zVMPq8z6P/FCy9VqizlhvtwcF8symtrMUWokp0QGtVS6
fuPwVS9+ExD/4Ad+g4C7FhBLl9e2lufhFM1fsFVzGgL9w2CR6KedcIBtK9bz
Pi2TLaZPi8b31/zu8OcYzD5wknKLgpwYCsnW+MGdXHMnLWXidC9146ZgXOWX
DB1bPulb5S5O41ew8w9VfaomOg/g+gTiEr9HIMyU+lo2LtqPZAEGO9rAKmGZ
yiVuRf+N30E+NNLV4HJi30iUVF53Kk6cnbg0Eaj9ZtdWq1S7ZWA6vKyIssx9
IHcb+9WYW6xO2z7+cgY2aesB+uI8dJjM9ot1mm06uMzTX5z0BnQLxrX8xuW3
UDEwlPr1msN0P1WU2ToVuA/O3B7E0GYAHgvT4wAv2T6uWSXKx0oEP/90UO4P
Oj3S/7AGQTurcke1g9o/+OOCXHIM2aZigjpK3qZ6IRAIHv2Mxc3C5SWK3qX4
DYVrpQTgPx+wNo51C2wcsfNfW6UOhCRilPlXqheuK/uSXf1g0xj0POvpGVyf
K6nLHbHaBNDlLr2Tcq+MqYmXnsFVfXrI/PH4RFE5v0TIEgcs9kaQJRwnaAPP
Cr9nuJFxz92VAT1dS9Ayv7Qv3RxmswTPHb0kKis8fxp77W4VHuB7KnjBG+Q7
kNnzeeWCJ8Uin+1BM7ANXWtiWZgUss+STe/hbE5fEekEDgjL3yJibY8HeYhc
XqTX836q/kAj2te34adOtf5IWuXanQQ1LcCxarLyZjiO71UCbcYXg9tzJ5V3
CMRHAHwIqOLUWf/zxd5udHVUdAgl2FUftRjG4u8X4yVmi8fQDiQOIP2FlJvo
KYQqQa/DYSq/UsX0VCDFlSu3idCqz7DXdpowK4+PqcWpL2/B46KN/Zvy5IH/
1qqTNyiGCTuWUE72LeQjz+yqHHDPA60lxX6YXyNL4Frdx6JZwNRLt4b58tDZ
PsQgzPBA+n/Jt38g3nPnDtaj+Gn+j4hF+CzgMEbzKHXBV+XgsUmen79i6QZl
91VpLduPcyjpcm84UH1Z/kT015ByUJakPKbKvYjN4d8+g964xDHoh1bIZk3c
/Zm2A3k1o6sDL9PV56BjRXc7aAxk6WOwrCtxYWMaFYjkGc01gvgSHkfGqPfl
1Mm3t041e+Pilan8wnlJukJYmEo3bkzhzaLwC7+jRVbDcVEQULmFkP9biWEe
trhGtc8iCLnydnOn8RPIIAoyYgMiUE4Sy5R0zEkYK1Z9D9Z9HaTwXtz6xE5o
xBOJjdx/DvS5UBaPLI3lBZbMGNxpSoo74euqmn8TLNjW9YiSP/AY+mOfBV+l
wXxI9krqUP/iGhbCG/h8fY+/pKrpLVxsjO3MOICfFV2UL7euXjEkMUBPBZ8v
cA0+CVOSZqi3fc+Ull6+x6s0mWeSY/A9fV1dApPUDm94QeslfsJNMB7P9iMG
wmBA2u8Io6GlQ5a2An4VZZ+OhAwzr37Ux7kMZV/sEf+3vVDdk2pJkuW5U6JI
z4Iakrr0x2YUhj8Ms68+Rh7EJySmLwDSz2FOJR60g3uafkwuI4vTREtcIwPc
Po9IiEOmXOZ0N69geTjjzd6OWV7tLHoNKVi/42UsHGlgnDIP7FXZebbmNqXB
ex/Js9HYsIizVKs6qihifizDN9TNbKeHEE2Tx8B2eU3EycnmQNOTPZ6OzIS9
lWD9PnHaoULalwfLhyCeHmKg98Z+kIEYmq38H2mJ/9WmHq/6GpS+F+zugbXj
seAPTO+H4oBWOVcmAequvtslMU/Z/Bixl6/r3OkNOb+/k6U19+iL2h5HRbU8
ozdJKq2GO8ZQH8K5cWM6GMttZe6q2YNBhBtniQi2ds8a+4veQU4tlYav6nyP
H1HgYQkET9qolRLnrrCAVQBh1IyFnO3fT/WGG4bQGVYT47SsWm0KhaG9+B1J
kEYYN9qulXHTrZ8rxxlHQeCGhHDnKR6mfC2Z/PJs00oikiWbLx7dG/hfSeTT
QeaAsJ0QLcH1akb3bWJVdxBViagxMF2WkMzw4lrJJ050HrvTXbxqyZKKrgv4
R7q32QoPg47dSraGJpQ1MWFO4XnfwSZu5SSGWeIDE8tq35csfZgkVX2CEPyc
fqTRLrXzgoWCIZz59W9okvsu0LHnyfgWHvUlt7nHBjZAH+TbSFrlDwmojwzs
VhhwlifuOf7Kk3MnQO49DXnzVpF2ws+nIcqYgslC47f+0+UIhFe+RwLO6p/4
RusKCY155ZcOY14fCEUmjNrSoCHxtnj4WQzXf79wv/Of6ZFGHJRd4XfHBg9r
dLYSmych3Pg3UkTwbSr3fM6tBspjpTazNLN5iBQmhB2c1/Py3AE+SzOOJ/s0
I39qBb70Aoib4zARcELxWftO1BE8FtT4PV+3XMnUhGEPyK+2oh/cxFL26vO0
hAM0NlxShdO5gLw60PFXZerQ9ISxfmDPuB9EPA7FVb5O7SbN5B3QOoZ82kCh
RkYsI2hBNAa9cdSBvumVVVSeiqu2jeNVRyc1RTAUg8JGHmq5ACddfMa7Dnd2
wRx8AQAOVr1oOvXamwvTPesBQ40/VwJvjsIG1E8zI9+tDQr5qdxOkGNtfKV1
Q9UMsqQ6KShPqwHItErixCv5Lx2ytB1h4M86NWDlwmGf0LwLllfht643afkM
hYD/vaTzObMCgdnTIy/ZnydeguqP4mmU0/NTyqJv2q0HiD9fGn7/6y1YeGXf
fizC1iPBeSaR3DDIIkhtriqz14MH5zvhVu5+wRqUqZpBZPcsBiLnNQK4GqyD
YbTRoUP9txJIfllp2oLmWwsd7tlMdaqHBj6O9B8UhFvSR6ZmSgdQ/7M+v6ud
vjYgL83mQa9/Iubb+eW3cLqWgCNhGxRB54cf5RgV6Lx7t/yh2BWJbGQdiDPk
/r+wu1IvunGEUdP89DBPSdsk5KlyA64mCJNCJk9mdfFrKl8MirMbgykC9H+T
rbzEujz7pwGBDrVVxXEv199CND5o+s33P1dkNiydPuYTvpwT7KsAxPDljGIM
w0LUmr84m3NT8iS78PQRr2gDIesUO43Jvj8VrlFpVdVfZ9GDxzCjAuGpeY+2
TE/5rJ2WUodHB1P3Zjw3Z0pHpyRXxQMQ80cvMu4VxtuWHTsiaP7hgz6Bh9Ly
PwCgO/9uKbR+0h7YobRd60h8jb6D917hVf8yWDA7eO4EqgNbjPUWLBkgFJBH
alUyVwb5+qDDVRifGVahMt8+1HOj0oIxV7A+Dwm8ZcEBw4cOrJQjHsou6PI7
FCSAGz39e8vVKlod+QOasqLVTyPsY0mQZolhNp8nHfgo8bM9vxowYGzXajx9
YiUcbjk5H2y5mPJ+cpq3AR/2mjl/E8OzY670GjTkyQOuByfnwf4AIwZi+lj+
OZLgwKNtFEIbrSPIM5fD/WLimNn46jPtyWiMkaw+MB2Q3nT7ULHitkZrn8xp
m+seWHqkFb1jD72k/XuDG7+Ulriwwnko92dKhVK2cXoL7wDgaBY+WnEyxyfi
LHIOOLRNBAxk50lfxtb2L8cFkJ+QRHJXJh9BYZ3lu0u2oG5BwffjDPwC2sKb
vLwybMti8yMLshebupIQokABh15l8jNeaBKHQ6m2rEEMuKXaLKb1HG62DOuL
ptA6YifjuqK3Ir42JS2FWVUC4fkRjBLs5dr4eMzIlnjd8We4bWVAtKIJ348w
lE5QpFcPy9yQBxRjDxLGIN1q8YytDyB9SYuE8eoF/Z8YeaTPUubjWwxKkLP8
lciaCvx6+L5f6issREuv/1NUb7KslhL2Z5kWlutPuv7WTsv95qDP46n/TR92
T+7xIG7Zc6Jp0nTwNHGfsQuvpN+9fuKZKt2yEZCqbPKArzFkqLwFDkgQSCVf
AHsGG2VMBQLCR5h7ph5mpCMg06hrcl9qS5CNDpyhh38ctNVMFNO5KKGDqj3K
DazhLoc1z5k1z6V/44inyG/rG0E6pZjjTiBAo3qpJ8M2c4OFPbXBma6OYpvh
ihcE9so7y0EB4+4Xsj+mu1dKIBDiR7NJ4OcuDBTI9/3plk+jWQ+Pkh/IKxt/
NJHazs40IW/zA0GhTTNZxlLgVDufjBAqqm7oQzwuw7F7MVm29GScyUd2RqSU
EDP3XFPHMTbi+ziL0B+9uYHMuorpUFSfgMVP0CLfW98ELT2Kup6NNuQi6Bre
rYHvqVQKge1t+c1bmKnRWC3VXl9htyTKVXrMiypQ4on6hzEmtl8ef42S1RFJ
suA4yfOjQjITxyuLvvc24W84vh3KsOMpTTpmNdxTc9aGwbrcQ0JUsDArw/HI
P3BejDSxnDcEZx7JONBaKNzSErqMX2JmQTY5B+ZWVaoFMROYN9MOSzcmoELh
0hJDAD1/vBVwz8MvAh1gOnqPBA1FrYIi5g4xvEMAjmXxDMGYhnJ/wql+kU4O
mKT3RwlcGBu0KrrMt1bNHeyF/oeER/A5jYY/lcExr/zIOCqY/ZmuI9oIDSTe
yhcqvXD1NYcgjpgwJe8biMvbQAd8q32aTIKwJGNWsjaf5xvcJh3A3MyBhaKE
zAZmq4kF6lHQxfoS7ZFKniGD8BQ4INWR+v9fvunjpXplnFJEiWmW12NsTNDG
8zXxU36ibUmbqJZTut2MhiF8TgLBSQ9fY76BhvkcgbwKCYkdbRF6dyjk04b3
ZyVFI63c4e08VGvUMCtnGC5PYAK6gBUpCljfKVtjdMdhQKzci2VArUyWWAK8
mpabHInHmT5xQhdRLx2yKozViKh5tVX0U4zAZP3mphyNWiDt2EC3dZcemWFv
MqiQ/eBoksiMFNTiLEAj+YzDoOOuy3yynilF4P7q9KR8job/R+h0dhzzKDRB
mGl/LlXkMRTfqTACNhZVsRVgdN2pmbEmaFLQV0lzBeWbB2IO/32BVhzKLCsw
GFV0nsoyE/Anpf3Zkz2McKOd2OJsqlliCoRNjZE+fHb1Atlb9uNttCb8keE6
nckHDDFPHintZ2HpvHI+yDOC2DsSiZs+U3Qlrg4+Vbt+a/sgxXUbRvnRiWhW
JxoIP8X5aavGPVnYfAV3BrmcA+AzEqFXZS9ZxbqhAhDpChnMjA7IbB7tJ77Y
HdC5BAf52I61cpX76CYloS4LTi2AN2/enSj1lh4Bse5BPo6j8goDEgmPeT1I
WZn3VC+G+Vll3s0NFL4+3K5Lia8HTMZ3K2VBFUoxa15PtuPJ8VPlK+aB4KcY
vPFbJpGXygUJg/DDLPoAwS2fmtzq3xRe3dmdwGgCkhYraEkRMCXrxQTjNVi2
NsVmbjnJOKrUrduEVGpD4GQpDjmMQSiC7BG4mCmHpAwUTksBDxFhDcvgnDpy
0NIURje2Ha6gNyHR7kM7AgVmNiMCBvEGx21E9phIGFYQwQEbA+K1xPAQK2zi
ND0C+nJT7T7gpAtVEmsqL5WbVKuUs9huit6FAhGYzIZAMDJy7b3MzaMYbSEa
kRXZtMRnlVRKLmwcOf43RcWPoodT64zHL5Lm5IXVslcp7wjk9XlnFhkpHsAH
ySBSnrw3RhEeyuuYWLS+d7cm6CF3nZpdolS3pmUqZ2sk+Pg80AFfAe5FmgEO
FdyuvMP8R71QapPYDoMLXLX/d6H0s78thW/7SYY06+XF+ajjj4vpZuRJJ2kE
ktR+6qk86LYL8eVpA3WMjyaKewtM3PMEmpm6xN6HJMfSIFMECEO6uXkjSi6U
CfaijaVjjQ7BIih9VYtcYcGoDH9ZqeLK2qF3rB4R4TvkXq0Z5Jgz/bMEBc1d
xG/Oz6yq5ygAqEQ5tPsa0iM5L9BEfXU8552ElABca+t908QJAj6i8iVIahhG
tEUgTbPeHSJ12YGsRO4vtH/RdfP7ychVoS7jdxe2Idyg1kIbxZElyW3EMf8m
bfvMCUIHkMsX5BW+ENqcC/w1oYUeWiBE2sCiKjaaV3YLruN5qS0cHvpyZfYM
3DviQtOd7pET9xM51Hem0jufKnL+wZRX+c/JEkxMwz3dgf5EmaCEKTneN8tq
Kz6a9ERPC6QMOw0VydooTnxzeOHTLR3qgqD8nxRaghDqGUUgfe7gTIdffE81
vtlbBqcVmA4ljE58Fun6IL/NqG5gczRVmKYPxncw701Qfxot+VTMIyE3y/ge
OC7CMJrHRNQB/1Oi/RNgZitSCs8acsn+txry55dN/cKfGA2NQUWCeEJ4Npl4
DjUHgMKTRAwCcHMUZB4kt26PTsytm4tjBqIoJcAUH/5tZDBGq9SGfOBYIrsp
lyWyCrZ6yu8u+ADiL3FU9xuHa98axTjQEsEzKVAYUxVDmwkFX8o0yIQu6u5i
wapLsr5UXhAyO8E7xwb+CAbgZRqRPrbAT1cN1KtR17iwRasLuQtiDIra0Z4n
ZOz8Rrb5x8puxjPtCCaMjy2rSMAyGBI5aAcDtLoKL4D2S2snaCRVFFcK+9N/
vYS72pARaUhknSQq4A/8brNS9ExdewpZcAp7Zon0UhhUHa0SM/bEjwqffERh
+n3JuoxxF4HoiRls3myGH/9cM6iyEXOD2nosxsWC1PWspbdaF+nrpkVPxrwK
nGHowZ6ie2k3KLrgNbmS4fLq2A+pjfG16lqobodP3uCNQuUiMTG0OAYfcorM
dv+4AgRSoe4PdSLuaEMuhuC+grCZZTZTn/WJWb/WejvqoCkkPdpAv3HCsnQK
IprVXeg9x/vK8ResT+3F8vniyJ23kh5cm4/0pL/GAJbCxmlmP8Nk72Bp8yNa
v1VIY6a+UFSUjIBsNwWJ8AN5iutEHDHkadlH/da4QXaGtXQOvpJ6GVg/MjFH
5HqDZf1F0YYEeeHTDwHf+PGnFlSAR4cnga1MJppXj2tkTQaW2rx4w5NZ6clQ
1M+joBbGT0lleBvemybZ1/vPVn8tdDCSkxkWEcU9HranMq5ixdh0qEJwg0Z7
KL8o5qyOMEINsMZv2fn/Fq3X+TifUVbpHgWTwFv1wOCevOmtYudOpZ5Oa2XT
gujfUByqO8aWVz8J9gXJb2Ny9rmRES3cRBziUvw5aQ/4mnZYwS4FN0Mtx3KH
+y7t+LEa6TF0UmHBlDWCPCzxsHvZN0kcXabvgj3FoNsQxJLQwhNmNo+/WeKC
W8xQA2aNUznItqs2e9mIpcixkIGy0hqiryj6FDms29R9gmHkBn0N/qFVwq4b
7MRucvf418YcDVAhAL0IdpgDTs6msrQ7wR5xGNw+z0HRKIrTLYK53sHD+9WY
swnEBfFCFUcXIT/9mPgIz0Thk07HSIypIEi6mC0zelfdvacmdmCylsB0WJch
3AuEWGkJ1moTxYZf5p3UFKPUxpnsU3D+QaW6YRv9BLDNf0XEqqeq2ltTP3mi
RzjTbesCPnmpsLmZMLHdj37m6gdAcrz6DTs/mTuCKAwPU1OtXRxYKpDPAc8X
y5jjjbQpZ9Ox5IQAuRMKRxmnNcyfpMIvETAAGsQZ2BUqNlIpB+j0ZWGzpwOM
nSDhr1DoC7YenUQaRLSQ7Gx0k9nOZIEfOToSs0e4RpromFTADK2UKBhzR8DL
eAT1iPdf5kmzlE2yVxkjWR7wDV74DvysibSYoBen2X/43uo3NnaEZzDuXLCL
wli9gQ0KBDKgyDWwH7V8Flak9LtkKspMR1Obd+pTaY7/uNliUKsbOcu2fzQB
nvejZ4zeRSxVPJmC59tyADXwojz5iVdDBhFFO39v2bt4fEl0aC3QjsFdalUN
iNeC+WFDU0r5f196cUcnyGTMcEl7PoVW9WwZyU31e9mdEFPTHnqky727jScC
geEODSQi6Zwy8+qblNBW7bEJPsrS3dLKt7+bZy1eMVh9ZPRul/VZrAatHH0R
6fPyppd7c6KjoDHvgzd+H8ayNmc7pgPg66oh3UxtW+7nEbpug1PMAhKD90gp
dBzvGuiWIRxb0VNDRxJOjGTLQ7MQffvi1SvDdXMzEDRhlKGSqsEj+Y3KinPu
noRjPk8Je2pB8wT3oWtwqEYql/ZrRuZt0lU+6hrHWke2KNLNaq6vTiCpvma7
mTT15oC9FFhUMU5voJfwsEVbkjhNZJuH/5G1nNlfOJF+8lr6uYn9CPra34br
g4rDaIWhZp6+tvQWusJAx67le0sZSVSxNO8IyNfPvurfOVKWgMKab+DBMlsQ
YYuDd/BQwP48lZYw/jiLOwkcS+b58eN+djq01CxtJSJ6bdMZb7wITcQPOiwX
OdmF8sUlFrNOB9jU8rIjKoDZG3+zuAyxOfQ5ZWQ13xWNkKe6xViBLdL42n2B
CJy9Xp21lYll89HyuGqmMtoxE88gmKw+6y8VADkKjwwohVF18tmWm4tGl3dq
TtulzxslwizpmCJbwmI4ZDY93L44gDSX2fnUecH7sDk1lLLurlBEFn6ixlbm
b3aZX+kapIK+Fte55pNyPXut6sWR+R0ERHvp5AdRmr51PaIO2luaFvvsuY+9
jRBbjeAPDlW4G36Xcke056eei+9FSTH03OW8JxSVQZZPP3VbLudWLW5Cabp0
yn2xIag2vfSucHxG8wt/cSIdvLaxJHH/PrV9i8bAZygAAdXQu7fo8ywmH1oW
gxRvnhPgMoh15YzbHKAPZoB1ksAOd2QRTXQrx265ngC/SNw5tYApfckd8IC5
MwoW96GqtfBA5VyBVIhb5lrmyYVl2VDhakMQoL/AixBZ7QlavSiIMHLxyxgu
tJm4aSJsZONiOPxpULuhUobVoA6DJWaZ327NaBYkYDvS9ThkFTgrgrClH8yx
cJTesC3Vtena/LnDGQqgx0G6UOIq3ximcYCRx/ojBlh2V+x5sYYpzp4fm1J8
+3goqGGg5RlIPEeccb+dypWxRzNLEJkbyUHW92/RMk7mlXa+M6SJiAhcuU74
AmNPl7OGRBCZ1RL+d8SrJG2bYYqbY4dCTGzeJ/0BX3+SSSZJpldJCZ6NFOfa
gYZsyXlnZ3ZUPU/vqjBkkifZptxm8IYSPGPQ1zHLjFpxl8K/4BmWzZDfu7rp
uio5roVmHHohQ3jFX8/vsEa1H4mVLIFZYZhnBXbjLG+bNG+3X/NiNn3iUlNn
1ohReOhcGQcE2Zbl8tXrhmcrRVFnJSKVaAC+/RZltsqVBblTrkLkK7EmNCsy
sRZ7Byq7Y1z8Exktlx3ubWP20PoTZ49con/emPjygTiKMzCpwxND/gRJnsaF
ecGjG6p1fqQpxknXExkxe4QcKZJRwdGeVWcHRxh4fR+F6TFnrEf8Fc7/AG/X
Boe5kXY2iGmCziij6GERwxz9pevnU7mm7+E6Z3SP1rbpiXaphtOGc61bLNON
Qvr54Nga7zfJClFTV8YOpuJdGef9FgcBt85AvFkoVgH17fvlSe7IoewCndBJ
1i43GlDzjbQjoaSff/jc8sRVTtaAv2221zdp+P6teGLZxHC05fQUWW7qJRyF
o0m/uRvUSfzPcDFQaFnYhKNfr93CEitoQeYexGBNpDt53xd+j+F6uPXxRGgB
0M+XFDL2F8LgcHY/54/PyNjo3IG/KdXQMGN818Wq+hVfo+at/INn2BgNNcI9
KWUXQqYYr1BlETyw8TWqXytPIfctdvjALfmbLlG1Nt56Co8kNKJtbTMIMTMv
53S4PGOGtpiDQ+rp7xXG3IkTvdsvLSSPq/oj4QZJomexFH9sWolYEf5NYwnd
qAYn5zpjac3OGiGF9v4oIVUYCFoFDY3qiIf6OPu5g8F9LPOauPqDo/RJVY+D
RFGbhDAvj2DzoxWYaasuq5jFnIEHjJe6VYF5Wfk92YjZ6FEgdjYeVt1f4aft
pe+D3MJ/mojb4xDAuo4MqhbfU+4+U6Y23KnYlT2IjLAGS3K+WDDn82TB4mwF
hGwbmZDhhPlovZKN5b6fjzaKgJpz3HfmsM+WcKdwdALAkipdDLKdSkFTfILO
jzTwGzuwi55TsE5tj4lCQwD1RHQl4xlM3BU8cMfD+BLV2iIp5GGuIQnnKAvH
5lJ9nf99PQnitTwqEt07BgewHVBy4zjP+6mmyUEOg2Sfpvu9X4Y8f28RkJBW
D2KC0sVJwSne32+LgRDHwHH85gyEogGi6ooww3bW6upRjGaa8X329zCGcX6V
PxYOnb5/ybo6Ev3NckBc9e0G053gaRnI9d/zBZ2j9hvKi/ZiBHeKa5hQyKdD
yBzTa2PcU5li/g0coTm9zQS01kyo5chQgmpM7NgYqQKEsBGtMm+yoCUXAD7Y
Tf3lpjZi8UjhGrnRSP9KTLXIqcYUJRgEJfzFi3gtmiw4qMGR55HjvxDbfy4D
Gd4lUqfPHrKyr90zvSZukfn2QFY5t5Q6jGEYIy7oIaCuzAHvoH74o/GCzbg6
IxI/M+MRtNjC+qfD7bhCiOjfbpFzd4Fn9bIEWxlI2vPhqtxb9n92z3hQMCGA
XkwKCiiOKNkZw3FSzlRTzTVmoIgrdpT18iPYm9cIC8LePzvLP5mpGGzCl52Y
/LFJ6SVrX7xaKxEAMm3m9kAO/EH6sElQ4ekLHv2Rmnoi+xDQgfOJRm6Qolfw
jw1x2QhoMBra6I1C7s2OQPQqZ70PUifT4JYKIJA6YI2yOH/EgGZQvjTnZN24
M5lCQQAT6yLGAGuP4g9QKR1U3b1c0I8L5UeP9tItqKSmZjeA/qIkM1GpjyTr
3qN5kZQg99UYbjXBfbc2opSMucW5dSwMCljDxAt9BAGRcBJVTbOIf9+ZanO8
SequNlSCKo7b9/IpKGXQxOiAlAHCDQ1+NCHkJeu092F3zT7QJ1+d4uvxZ50T
+fFmHGRMgi6jGPU4f/AfpN5mFycqB0gQzaSW2GRIi/EM+2wbFascidvY2xbY
JZ1BukwflXJN3x1OU7I155vPloiuK97oeMb6fSGyjjI2j9+bs5bBpkejxYIO
3rxHGJh/9OmoMgIBqCTYYcnv3Qm/hhj+mqq9usF0neO0CQA52f/+16fM+Xin
of6mNIPg5BXzLYYOR6dbdxYReipGLS5h4co5uwdiinfNkbQmB0nyE0CoIwED
5LjRBzEUYztKIBUQfV4RWfQvQLozFb9TZNpJVJrn3p2s2Hn5XQ9J7YfcVrW3
1+CMOrmiLl871ti/wOVNN7RMRf5OZwbWcWDoOe0IyvizvFKg90dM5fFVUxp5
gEQwy5qjwi5auIoahmma7VBqkfjwusqEAj0VlnerZYABs4HvI+H6ih2UEqwv
+XmFHCXaRFALmCDDi06tm9hwvayQF1W8AWMoq2SjaqJY7oq0Y8o8yLfAg5QX
gOlTfWqDQ9CV3krCuZr6DDTosSa8IfyWSzQAxRfE4vmxXfdCQbNGSiY1BeOs
/oXDiAC2BigY7iRpinX0uCFoLRX04IOwofw0JIdg276PwmWBqr2a81aBAngk
L4DAXMksOojEYecbG+n4z3HfDveTwSXMxWKyU+57y8UVbaTwuN1tJ9DFECPX
tbQ+8Ly3YqbyjdKLgoc+aHhwnWkwoqlWLnZU51zWGsOvGDfm8CzyNVAAxaa4
x1nh13r4j/x298O//ZZIpGQHV5JvsqJzW8fS2ndrzf/oa29f+ai9CQTsDaLA
fq1/nRgkC8pWoehh6czFz7UxiOddOVW9eqMGiUdFm9UifTKhuO10k81+M3fF
TkHT1N/rzOBp92/9YESejxYp5Mo1ta0n4QNgp7RFS1XDPpFiV9H5b0piskks
PW4+CzXM3pUt6cjmruNHmr70VfZceNMzWaXbTbr2Ts6oyx0a6RMWU3a1WeaF
cF7UlzcG3mKHOyTEIWXZraoDIWhFwNJTPTJ8TAate/s8/O/SuFz8Rz7V/YIo
HbArTwu2/LZeJ0QJtGnACTNyb1Y75/ApDr7rThJq7e2gnSVhIiwSeACd7N5r
t7s5b39CHc8QbnHUkLcEi/q9fXIkpXB3wsIQx2oMD1RqWp9xzmhm3Y2JtbTa
/BFtlxfJXpBwev6H2wHZ03dNK4cQK0cYxDEw/+MvVqFaufLTX/HfnuVbmXat
0l6vn/TyXFyP8BfYbBkO3Tn/9KBBvQP8dWnwm9xO79uKdYWiHsyVyuICjkXZ
z66xuqYA/STvsHweJq8lfnjMSYOwkaXdWUm2gHcwN1te1oNZa/0Y/wocjgAH
8DXXBlNTllqHUv+f0UzGhdYsHoz01SLpNkNG3ez9Gq72Z0tGEa/jqqoXSEpl
yFOqtPReBj5KrCc3u3lW/5O60BzKwTETR7/oGoOJHXmd2uBUhSKaui4vrgaB
1nZXIZo9koveQfKVfifQTrFQJFKwJPDMdjQpf0Rer7OS1nLrvvq3KbhGmp5E
gwTeM5/B6EmROcaKSO1mTgZWioRRS/th4A+PDZFneYVlRpJ/JPwsFPRxeyde
h5riz9LtO8Ji4fHHYmqHEIDW4G10y+xdoXUVvy16f09cZ+vdtz57MXAGWw0G
+I3jCiBy78XJWHvbAhmuuCeQ3tU6RY1XzugsODGxN8LVXI3XID9slgrEmwK5
OJDO7dHkYxj5RwKYGewHNVhf8f7DLiZjDWlpvsKzRiLqQ3m/n/L1mhaEe9EU
kvTL4OQ1qmrJ4ZQUn/kgllriqJEb5lT4YbxlsITJK/HzzEJThBSimc+dyK1s
ZcL0mXwS1YHUDvnaQFGfNcXsdVfMtKxsZy/VHMEMYxUYcYy+yv/Mo8Knf3YM
hOKSmfXmWrVGfFAnLkikgEyRir8hvso9/G+c0W/v+KWDPqd1O364JKK44Br0
cYIEEvu6IxtFR3qNaCNAaxVRxnqKI0WLJ+VZq5y+tBMxWTH4Y1LlDi9bLy53
RozB0MjB4YAR6/9T3iT3UGR2gN2+9qpn0piVc584hx67t1RrfNhN/kbcj6bv
5nTUToVjC6l9T23kZ4Dum85llGQA2cpKfKloS/CicSO+H3cOlaKapVL/S7Ch
HvLtrnnGd+XavkebcOcjapTCekA08tdsts24xDivetBt4/pZJyr+jWHNlU+l
9vdqcCcRiVopbTopBztLdQON0QuHbbRA/e1xN5YWlnNXe4AlsxsFBt8m1lN+
Y8XKXcg2uWYbDRgoNl8NdgtAeOy3xCxqMhO3UUIVHUrPxawFWl8hV+A0eGPp
PD8YO5DPjGrR6FjcimS4tVRAi/jXNmZJXDrYtlCdsckkcZaxNw62M4E8ABHo
DdUnq2GDJWyF47Df1l/fPJfBXgPhtiMpGMc5Z74RfcIyYXB3pT4x7odvL/6M
q1xY6P1VVpdAZ0Z9fU6fgRhYNyCW22jvm1TqZy8IxLWehknWeC3UYbPiP1QN
YH1nsNCnuGHY/Ju4sNG8CKTeA3x+qHE0V5hmKxI4TqFNw9/sXdOvf8DstbQc
Wk3I1IUgqKabyDzMx7pDmGd13Xd180kJfiH98qKxBDFQmUzJaeGtfaei0rLe
cXhdmjRBn63bDh4vpqlKsmF9n0CW7g1KVYVUw6bB193jwdcUjG75lqnWd4Ta
lBUVFGmn3CBjSe7gfEJq/QtP+TS0FTMXdXaZ6k4OOk+CX8QV86JORSprH4/T
CpI6WHdcvuHA0OGVtUbY2QSFLhLeVCxbIFNKjGgvdv6iE9wuec4RRxt+AiHX
U9AuUlQS1D7xUuXwtVHOs1DIFQAilFwVkG3F4P8XDdalK25mbYfG1rEuKST+
Ff4+ehrsdiNXQkEKx9BUg9OEoTcYnvb2nRG0Up3pyK7Nv7GKlY2whVfc9Avt
ZGKzgzndIynHKGx/kge7E151P953fyP6+wyJ1dFdyX7G8hUfbGd2CQn1t9Wy
YRjvA22Soh/ufqLTLE2jXqii8sYlV5oyfOfV3kMRe3/go5q+hwkdqZg0vxUP
QHpopqEvUF2NfQTM/xFMIUYPo1idzeyRM9P7TWq3EM0/JzfmM80IsesRxtrM
kmRzsdfR4H5urAkqLUcHOfQUbRw7WpzT6NtWDx43UHPY4B54JSCa9VOhbEMP
96O+XK1DJ8N3saGco+zeMigV6cHDM2/Pa8XEhX8AF+SrRxSAsIGxRwaG7Uah
Pr3eeMP6ti5ucbohQih6CHIQdjggevppzrVEwE2CKAWZQB3Q7g++gn0zGcja
JF1Ydtqt8UGPSnMtyuyoC+lWA/2G68gkbvu7rgjzN2ygJ7fliaiTDun0AzCn
zFNx+b+cd7n+c5OtEHgvk6hSiRS6eFQBqyonENO1REZMxukoAwXq5EMWkrv7
TwuPVlkr9apieQW+ugHCfODTPxtC2oIXasj5KkduyVwEto1Is28nWq5wT1GF
xZK92AEUoz/nNpVtztEXbF9yMl/75ifSMC53h2O8acGYsVVLHEQ1ND565NN4
ZqgngicSzZkg8BzMEidpRxbodBafWdyMCelk45dqaBXIVD11DwNP1JQBuNfk
1KTK+c0P9FvroHulqd7apaueEm72wneHEYKmlRkQHsEbA97e6wUyUK7LwxuF
Z3y2MQynRL9bRlkJo85hLs57pnwIhZ3+I0zvVeZ1bQdBtTgeI+LXCmH8vjk1
e5K3Gr1CdXYXDEGRdOMHnurPF7o7Q0HfNEvf8BTmRhk2sA5g2aPS7e/L3lPQ
f7ZSzw4GJ0+/0PdUibtNmeOVncwRHhKx7G1k9VGgZ7saZ2mkmiEBDafQp2uf
gA1I/vinIBETJ8qfy7trSSahv/SotOCotW1YUTfeGzMtSdms6/UyKXIiTRyh
MuKp9Oqgwtk1A3Q0zolbGzS/cAbhF4HAyrcBWbrTg5Jp7LpnS2egXXFZuuO4
kWtVWge9a3lGFwgMnuQ/cRBoCwkuqPvRZAx6EWoH1nC9y1a55pQbf5vtZHKX
gaWBwcHZPVxh6QdVzz/d4jAFgexCY93JlXhLJHBCRWn1nfQKcJCob1xcXiyF
r1HcNGvfk2Co56BxlDb0keF4PH13ZwBK0ShX6O/kk1ARkz/R6Xo56j2qFr7C
9g/MMPvm0DMsXJq0SKvRct4qWB3g6P2os2Gl7Ilqnu5Kkg0LbZfkk4gg0G5G
AEYZayuMWX02NqrkBhlgbbh7iDUKeDvJIBkGSV+XrAPRKE/MMnkbIbjvnk02
z0Rq9Z7UEcrIJgnq5LTu0lxxhxzBZFjUDTLZC5OuDvzdf/w78k8DyZGfgfX5
O+arVWqpH1eA4XRu9No84WMHRzDrvz2QGjPJMr7sxZeczbaJ3tNRkjNGJCW5
ih9SXrcGH2ySI6xB8yOAuSubHIfgq0ENSzKs3yOuUtav+fT7hVa1RHLHYYrV
O0+tA689POz5F2+Gh0/RNFAHio7cyI/JDdO6L/lk5Br+yixOsuSgA+bOY6u9
TnE3aiS+te8D7jEE51STS8rTVcK6SedvV88Pt5QFHQzfwYi2mlQvZDRRnfGu
Fo5dpFQuqyx1PtCW9NVWFqD5ta+9BYj7nqS2Ee0zo8OB7HyKjWGSRXxHy620
v7Xpgrb1SyEbe6ygAy8mjgEzqB7dd9hRvuVsTtLjZN0b1WsXSCdiyTMQr8gi
mcuyzaOtWLYqVXMShco7WldJEcdgui53C7qj+TolYb7BRFgeIfbm2qW6U9he
brH1qWsb1LZp9GtKpQL92YRSaN3NXi3RgBJOhWF7bBboQ7t91ps324bf7Vqe
QIO7z4/Ee/LzVs/fPcY99ZK8aKaO7MsMDqVgIjxcRwdwPTu4x9QSLOVrY5Z3
RKIcUyp4fPPtpK7kTv5pnH8HWm232uYVvgUD7fLiO32VymRs/rP9h7xE+ceT
O1nzSFvqVxN9EoAId0wG8Wf36EPWXfdK3kVnZxQDnS6s0rQjk+9QAZh9giWk
ndGfSu+pDI1trxB8NyQV73rj/X5SdnN6sEv4Y7KfAZ4yhrzznFumADpHEJKM
6ARsxymcAWy6Te7n2z+e7YVS7ec73evh+KorWUWQl+iWNpdw/Weet2E+iEsP
gn/WzYy9ZBtqO4qWFGIak3D+Da0NTiRTSYXgwtRG4gLopifCutAK15rSD0i5
C8HXgSmlP/H21PusgOjx0irRYiwN1Ft0f3PVWlzLaKHkYF3ctCIeK18BFhyU
bYnRZqlnvhNMH2Yxtq/gbhpVYIrzeJlf1iU9NGg6958s+uUbE9uAdN3VlgGc
p6G08TzHR9CK2voJZeonKDQdZZa/k6k0rAlpMAQktbCmYblPX+GeD++/db6p
fgVGr5sWshohD13n81KE+z5rv+npoCeuTQWpK1IX7P99DfrUf+hFadcpQHUO
aAwhQiv4P2UxqsNAj93IBhCU8ew3HBmPnbJyj7bz2zaKGXfnwHYQi+kZYBc/
g2iHzM5RPoAq/+ErgECHkJLaXdVEGTYVsF9EpsEUkFqOjZl6QqEqhmSSmggm
gC1VBuu0WrV/v0GmzVOfaRxXS4hqPkWyMKc1FHVCq8Etve7Vb+vUY4qW/Oyn
1NGwjVHbWdn0n02s3Hp3hW39fuuMjKiCHn9F+NOCs7HgaNRlkZ/ZGe62ouA2
OdR7QVtrgyoub1NqQVUv3end+kfo8m+8V5lbOgHCM9aMhpi2YDnTWjCY8M9u
73MiVgXYUDpTT/KxRtS+3pIIYBHDRpx1D0SO2IXy2Fw727OugdVAERklK4tn
ni7KCQKAM6/TQfgplqt2d7zujRjD0lJzwOiUZuCCXF9/y4JIGJHgw5OHOhHK
CLfIJNM6WBtXTn8NQQIJyCSeLsYm36I3lRH+Hqsbg9zLRFUUzyfZqKlZnjgC
X7B6j3Ey0kyAgxkuaWWYunK4A3337XLwpypYpmkkPWGymqoXRqX0CZbZORoj
aoWE2PwVuLu89ow2QJstuFUeKdFn3Bqdu8rpo3qx2VG3RG/3CCZxD6Q69pe7
zK1/2KBvfGWxyvBqfEp/7yI57CeVY/3/KOUUr8xBhU04SUObPvFAOSdlxidJ
kM0AHAWxefoZMRLlqpePOyFhT+p6NVpo2SoofoQWLpVHbAcIns6PF7PigRY9
RK8KLPuIaF1KZgCIMHrNw4Ht4StQ419uZHRYHC/xcJrrnsFa284VDLJuyXSr
cCMjrymfV10VAVwQBcBFcW0xoAkRcfW+r9BatGVUBkpgliIyDREwTiuP+q76
5lxPsBNBZ5n57ey6TIHBIo5XO/6gmQJ6HPzLYWZbTNttD6HYjH+vkQCgRWR8
IvzilQM399YzIcIyJq8nhc0dEd8dD5NCD1Dh9cgDAWzxdP7qXcphx/yJsLD4
4TGCITnmzvDaEtwwIea4oTlfAYX4u282GcqAo3RqjTKHwsQQ/ipZN0inK5Ww
e8ceASUfGBgjajqSpz/O+B9Pf5ktGjH4jlmZ1jXrIfmxi4S2teaIQcbrirLM
FkrG7cpM39WWdMEKcv+QFyTaE0rxk5mJwef5jr2Vf2j8W1KCtwg2dfgNA6+0
pG0K3UCfFIOheEpYcNvP1AzsPENkETJsQgq+RTx3rNkhR9vA7ZbPZoYs4d7d
y4xBQMZwOju/BGPYpKmGczKz9SIq+SaszsdvObc4w3/lMRZ/52ASe0aNNr9O
/I5rcDySj3pHRe6YVFoNBbz1WSmdeLF7H6euH5413RPdgew7zrbN6PsjD7e1
MfJFjxBAFgmX0O6kKGI2EISRSm1/FtEpuTIsMeYN2/BVs2EOGYic7OJKIpJn
S/5exF2zKueWcD8+9nXwgqzYlzv/5QNaO1YxvsGpabhBsHJEFVsYBgeecFnc
Sf/GUTCFDg95iR1tRIjlOkkgT8tTej4F5XvPD90woGinV9iCLNjhXQSmlr3M
kv/ZtRiQFUvBRn5zp2opoZe07kY+uFOkMajV3Z6nShiuC8nITnCefPJ6fPub
zRU4IJE6yXZEsl9NyvcL2nbIDfSus32Ep3pzXDrMrImOGkxOR8TliCoZWqvM
0OMhhl8wLs0R++UdqlK8pIe+wheOngBIhoNGCbakNsQ7LYa66VJeRfFiwylT
UPcP5sr1F6qIzphbifVkJkS/Jn2+mdc56oV+IRuNHS5UR6TD0oZlSrl6Qkdz
v7V0+NKXxNztFPg96y4XV3TrEaEGX/zDl+2UQBD8uFryWjrGYl5K3gmcXBXh
MVkDFIy5BhJg2kwvp19E/QFX3qt4ELhca0L2k4pVKkQPFOMJVpDFVbgHCtuA
gt0Mw0I04kGPCiYqxjN782iBNDy/PAZlv7pWYso6vDkYy/sk9xqnfoZu1TaS
SVgPb6bTG735/jEeCHs6w7Yb3QjCnccG9ofT8r2yWNLyAFGcaRC0lHLonAFu
ZY6LStRlYYyFFuVfr+kNMEIF0TEZO1HEid02WtbYXd36lK2YKpeUWwGrenvz
vA9c0gmUCVxMvYZ1iWJAyvLB79dOzgQmTSE6LcF8rYHZpdtQ4+TrQ1j7N5ep
DUzhwMBYv9yVQ4H6t2BucLRrdPuJbFzt40VB5cukfJETEdn4G6ASpaSn7TP6
atfZZNHsxdNGTpnusXnqbfEW2SoJ8cZpGG77WYUjAfp+h/6x5ZACCWtLHXaE
5c1e+SJJB9F0fhG3rGd23mu4qX8SBHqr+NXoeLkn162gB6r/IKjwxOq0E6DG
aZfaWLNveK6JqnIoM2pjlgNeiV4PyHfL2ffiqxJ6JDNW6BpAmZ0B6mGKSz3Z
yfJd2bgl4oNc4GovnLAiVi6Pz5tmYTwmSFcttJ1f3vLZ/E90bvUTjuJxY0Yx
zkqLTv6e4CYG5+ilD2O/MIMD/xHLA59GKuwVFuprs+z5f/DveBYBN3petpkd
JDjS40umJzBwQt6Kh8Tb0mh6gcyPpuWwuGBcfzgeI1UHTJaz6ls7soqO4Xgw
3CRjyR3VXHPovA4h3nFaHJ4pFnQuC9pW/eCrHWmdooWQ7Gj6mY15kDc9y/nI
/k+cPHxY3yzTnNckM9YSFw0dtwwGUUB8tvpaP8G72qgfe3RPKHgMPH42mlSQ
1BxLUPieB6bp/UwtGFhKgjV7dbvUX0m1HYZxiKpuyO6HyVjolF1yISBcuvVz
XAEdlYqyhZWdP559yOsLTtRr6GY+DX2arMIg3jtYqgDN9svZ2DjgBsgerYYa
XKJAgR9ePMVt5d5JD0VvmyDy9fhHT8B2n9Nfhn5TJmtc+qy2SSo2wQdlf0uL
zhmY5jMWj01lp6U6ksRHEBxoEyJqAV/96bG/uW5yxuKjVZuJfNaSDCVw8iHf
o1MwHIx/hwpTHadjkZ7TqgyDuXoB0UiNkMynupWxLkQSCAp53tjVk7TVFXEq
PItOs+fYJ3eJsaF95dZtjVWozWaiay9wZDHXYxIuq0Enu8cJliHZrVZsj30R
BUK/KUGgztGaXoewuM9NAx34mCy1qwE+8D7yLEtuTXNJFjIqN7IadwQtYEQy
9Td3YEYPO1TpO3XSq2dF9N2Gctlcwho1gJvyuiyOtczubhPLm4TLJhG0JV19
1K1w+8Y/X/TtA0lwg63vfuOws8tCay8WMu/GDm9uYhcJKEoL+3A7NNGPQaUx
jufJU3POJnYvDC0dqulFWZj7Jcq3rGsSGFsyAuwOnr4TmkAzQg6woxm+nYlm
HxW4My8uASU4taWmnqWpQ07ZNWH9vzbXUNnlRV4jk2ef+uqPG5IXlMaQ1iOM
XwVDTiK7XnCfQauPGjMmgKhn6vKyXds/pHiL4Lx/nVIX1KdNVeZBwXbW1gv9
+ronfjZl2A2fKNVa5eWElKCD2+LONnT9WRgNqUfjeXzf8h3phkPuotWZnXOI
NNUykOhdt0ZwU9ZaWAcxWJO7zlopVO/BWNJYzxjwyOlZCW/4IhgZguJ0j+KD
iV6DQh6hniijaTeXucYuQHDY9rAoGc5h1imDYArmlWGZtXChEC6a0dARQJQA
mxFUv2TRSkTnAXEC9h8DmobAMKKYSQ28QbxCk3Q/f4582WmhfbZG+hSPvttZ
W+Y8PljiAAUNYSALGLnf3Ry+JKayU0ppA0PGPYtLVYeznPYhZXQ638ABOhkf
TU9bNjkYkl4SyLVPtlel3ggS7Q9iVzIMDb1kfZmQlvFwrdNOEthpBmLIB0LU
NOBofHMKXkny3X7o/kyjb3zwG/B1I+jDptcXUBSYAQbAAeLMtLdPzD6TKN0P
MIQ9905uicRF6alh8sGYxpuTLtrCk2PxBV0YFEkKWHYK158M7BriG4lgxHnN
za8J1R1E0h2/mC13pYkMKSX9Www/7hgBGDJ0WlNCeOY1rI00OVR462bPBmMx
G+i8LjlWzhC2RSvReTy7pXoznkLzZPjhx+3hHICgtjWg21NKXFG3pCRWZ0gv
8MY1AgSUaNj7QzWzttA+mx5II+LApie/pAhXH5ibcUG3xmGPYQ2+2WJ7RzQw
JrO6x4kCS+m7OT6SVxKCr1pZ8MuVP57uWJ0b9jc3sBZySZ/qusRfHbmmEAiX
ilJsOIDqbrrb2b1aSaPobJLQazHqMB8oH8mNrl8/3GWamPd6wMXC9lbQQZG0
Qq3Wy5fgOU0WgAVa6xsvm457vkOZCGFD+otv/Yyny5M6S7EIRH4JXizTlT74
lszasH63YyN7J9IqReDgaXLtdQhtTR1aH/lQjWrQnspVsjXrKmi8hvS4BsM2
qTguQS6Dl/5avQW/ltHeb2zd7IZWiLIdWv3DT72KKcvZ3RPm40WjerEKUbxr
YSeDIi+BBGC1ngpIU23IgvHA+7i0uLl+OpKDoabTDQalFyFj6h14QumT5jFI
UwZ1KCIglunjC/msLdbp6WiwJanBiPG0y3jfdhhGp45dwXQapVLNABnA0ebA
AVQEZDGo5ks6b5xCrwdo7YyvT1NU9NkzD1aG0nXsaFJlitZB9lF9wy+ANPKz
MI+eeknfKg6HU2BtdLhsXx77CKlY7KG3w7lXXJmTmTkAvm5LYAoJBDgMU+KC
4KpSac36t+i1YZS3x0UmRZEnRCY2o2KbiayvTfXvC8mzbtSEUhiOIM/UnGls
turyIoh/qGAGRsWhfNjWDkcBMw0PGkpBo101wa8IJSp0Rs54mv35vOxP0bcH
epeM7KSRtvI/WW8bL6MmdQZkD/gAlwAszFnxTtICoAZm29V2L2910clHC7oN
LilHaqcle5p9xnh6GnqKxeyyQ/gyOFjU5voC3tw0sFrmSILdun5Q0gkdXVpw
VnaZUZJIF2gLfCSiSDuFeHvHX0sm8G4L8XkaP3aDUsVjD/zye46Omi88AwPb
qjNPZr8avEv0uPjd7JNSjzPBptxLEIiNLpAUDPY11HuCUdtnEfSUsc0r+eRE
EGupDEG6AME0MGQVf7Vkw/UPKKA1flixo4GgNaKQk56PPX1VjFnu00CLE17r
9n+7rfmybMhDFrvFlaCnUO5+kzbpbvyJALAXeALpR9SRJI8rMQz60NF4Y+ky
ssTBUMoWcu9w/sHdEC3IGpE4B9oqxcTp3KXyrFLPsgL7R0W/JffMDbgz459Y
k1kTAgd5XVi4CevcGBMDGje0eS5ULekjb2E8aS3Gv7+buXcXTCdhQnOjpy1s
vzjPenYpGH6mJfs1BnN8er4nd1l0oztDMtJnZs5cFFESw5wpiCIgFG2XJRab
GodnbLAIoJJJAiW/EJE8Pm7Yi6YS57qfj5C9iCi9DbebZyPx5B3KZaDtAfB8
B6vziwG2njmtCgGHGmNaQirWPCGAXkSpFshse6FPlshXcCe7/gAfWJGS+c7g
cM61/BhLWLDbIEqnTOV0H8WibH9v+Qe7+NyiEm06CRKEptCF7S81Ox34oX+7
/EgfF0e6YLkgsceFAWpDbiZAtoxp6dWaY/gkk5QmEtVMCeJo7BFY7n6VXQWa
osy45spBjAFM1XYdxQkkF20jser4/2F+2aRykdg/e+akCj7BiR2+fsLLGfFS
BbJlF8NIRF9kBMyuuauhYtzRKfA3qJsGUWnuWLFiI4jS10mOcMFxcbtiixrw
ZaZuVW9lawLGT6U1yj/L37wNuKcAC0hjV60G1oYaiZf1BwCaeswJcJClj78h
9QaVFB1rlrA9CfAaBfgL+hFG8VnJCnLNaoA1y1DhJo2jsrGmWmi5FRp/yNlS
XD0CCRP4udlnTzkiV8rZAeoXZGbJkywPZ5PzGym518j1K5Tv3bWBi1hJDPx2
/MhaSOiopQgLVUTTokcbzhFnxct+CReuqi2Jxx8+m9bZpLQlyTdBRO5WyAxq
4YypbUfk/f5FmjhAIqoPR8UYtA64lj5I3QdikemV7eoq7lm8keRO2QNO2T1M
x3xVZ7cd2d7c9fUASkJe30AHlPYcYdvMLggxX00B34aGKbr9CrRklJPSUDDG
e8XboTo5m4lfkRnWQBbV95JzYyn6aDVSh+wSEXJZApJRgQ35n/5vdXjvH/t0
Pbm6lpAsmoNyevtl8ERGK3ERkocM4aB+h/hibgTUTJjBFt91BBvL/c2ROeJZ
F+izhFJESw09LZujPnjFjjYvnf8chpJu523mQj/eIwG9tBuAZ5jWwPAy1Z5k
nto6yhE0DxG2hI2uWpHFd7kLVYklvKNeFItl+lXQl5x3mq+iszXtB8siUZyR
q1nJswzhNVTknHOXgPuN7uhLR6j7eppRHLCzdmlVCusVCE0cjBTBLHqp2RwC
DKDK6hLT1ZJFhqt3Bm4FOhcgWFzJKpML4HK6Ni+E1PlHU0zr+X0Xok3qpZzq
ZeHWCdCXN5t64IuNkWgtg2xIplxR0YLLSpKCrzYJUkbIr69A9VEleqbeYd0d
ypidlau8HgMpZ3H0rHtO176fLOH8UCZ/xDx6kMufZOw4DteA/tbERq7mmtJE
6R55y4ZfPrRljoL4vlIt/LD4vKMaocEphAIwG4ft+9SuAknkkKZoe9+WDMwD
Rdr1tN9zNUxCf4SQrrZFfKjs1J9OnY5biNEJraV+eCCCk0BCzLLxjzgBgktt
wwnMiVjl7HB6ohb1qPo6FW6e0psPt9TnE1S1yL/nCUN//FX0V8IRgFNECRVb
/t8Jjq1jSqThhhvPxHw+u73epqSTDmrzehFhVfjPXbT4o2j4TxXfo/j8LexT
rps4feN980AeCHFe3KO5IyhjvsgZo0fMzE7J1HPOKV0SAbINbwnMuxPae9rj
R1i7nikaH48sstSJAH1QUD0Y2ZEMuLLsp9+pEcJj6+SFk80SQcyNGfWZR/uy
ZwHvPkVeBc/OmrsR9q6xmzTiBYAy5HTvXwawNELHyAjUSQTNezfpWJDUdzDL
smxn5qNUErEzvqPsPZikQAw0a7LQgLXXSmGBpcfm63RHy5uWCf6JLylQL81c
GWFw+4n2pxczYfQyoswO/xL4fScoC5B67s5Ru4Q2FEQp0T7gFnoww5skSZ5b
HFV1DpdpFFtf9BK1x2YCsGbhxfO26fgqjsSPrHGTyhZ4Y6SDWE/MeB3wdS/Z
m/zhJfpu2RJK6FxSLcqRH7Mt4iLiTJZRHla147FYBqrVjcdT79MUb60GCHYi
tYFIAf5IUIXUJxhN/IeUSuk23n+AdPP/stJgheH4G4+LH0OAg/5CiV3qpqui
cjTg0PzbhSyT7WVB7nHvcfmdUYT5VMHGCThm0y4OSn+qMG+FtIctYrW6Xoq6
xCwFhBHPzzpHripp9H2zdtSsHOv03wDPgLnP2OsGEE7Njg+4puu7U1W/KCks
PLLP3I3XXAEAtCr/BZW5zcsCo54iTmwzQAKOABtNw+xWOrRUpZuklRAdxe15
3lWNSqFt2KpZHR3QBeWkKqEVhNASKpy3HeLmgp9cpHaOQS2H8bDjWdDSF9WD
W213ZTZE7GfnSApVw/gnxDBlOztBPu4x3RbQaS/erSw4flQytAFXZO41pHJX
bLCjid3MsfnfQH9y34TmmYFxT0rChH+xbmbPuHLayfkdKuoGxVNxGgL5YtZS
RlyZ+IWbne+4gaG1v94OEvAcItglfeZWAG1SVHLOi/L19pwJaSa0/wVXerGI
WpBEMxEW6Ss0/Vk0jx0zUi4X38TdcPE/Ikx5vEOtSH+hVFK2H7i3fC/4u2q0
LVyAEwevJURkXbrMy6cstt6l5JCKMC1JyD7znZieBgeB3xEqVeoq3OymvR3f
z1Uber8eZiYnn1J5uB4IIWx+JLQtVGAzS/1KnoC26+YiDCRlt1WToZjbf1z7
7UMH60pqXQreZvF3vH2lBIX0Q6RRf1KJGB7r/PJvoN4xY8CVgtFMfHybVtui
zZ3+FRioLSNuR0mWNNiLucFXMK3KNqxB0tndV7jmcAHyyWofVbBsrwhussZk
R+6WppPDJ6uCM+kwpfAMi6iSUeODqTinBybpNdKlybWeRFFVVKvxygdITd3B
VlgBMQL//NUNFvGfPtmhKt6KEN9wt2ybzxK/cD6l29BgzOKEYYa7Ymw1suoB
N1p9NuS5EFrhvu+Hrf22d6rr3Yu+lLk8UV1sXD0jHv/ehLs7dRapfYdeQjXG
ggdAF+AaOD6o4+pbuoO3taVGk0l+W+VjiW1OAjTeuOfAp51oBn2ARtq5IghC
kPR3Y4TRTAUf9q/9fiZmjeSK5Q7f7hjR1cNKh7omttUXlFtNqL5jZTak5qZc
izMibgMN3TXd/z2m/pryknX7feA9vdHGTeGxFI6tfTEpb80Sc1ISoD63JRO/
hsa+Wqe/Y9j1MTYDWxT89myqI/MzZrVbwuP3qrV1XPE8tAUXgx0wBRLzMwIj
nvvKX76McMDRb1hyHkurfCp4duGT5OYHiBvcw6a/NNS+IMJ5CFWXAqANVBY2
xoUYlSQ4TjDtPIAYTQlt+zGkHMSE1TIkvGy8+30okOwfhmUsLRolV0PdVMEF
VBOS6EOSFzu9w5zxSJz4GNpNcyQxjvNi7YGtqFbOu0WSImMoZfXdCV2+TajL
g21NwHWuJ64INRVpfix7l/8qEXwwsNjlaaXeunPtQcqPV3Ys8z14cGFyiDi1
v9bzkPd3vRtqc3/N84yC5xgSkXZMyU23xjADJysK9PGeFyUCn6gbab7qogqC
7t0uWPIsMiUzAREG9SNWbv0gB1wDIg6JJCYNXFnmCZznCFVnLphgtCovBOnt
m/U5amrjVD/k7pL78iD4Dbh1Sygcaf4RbTKaXaMzurSLSjo+ohMQJMkcxdly
wkK9KBhLXPuvOIKYy+sFKI0hXDjOPBwG6Qy1Wh4ERZBnymKCxYaEyDKaumVH
AikgH410szwUvHiF+NQMJqJUzN5y8Lhu+E8ZVW0NHGEZZX1CwvUxolpSqpb9
AB0jlvtOxXRXZ1SLmeliGsEAPuqKZ/JUF22RyqWwEDuOBYaqXBGnPfz5oXYs
GrSppfxvM2erKKbL4dXKrD+FnTtCmYEdgNM6YfunrbPttm7S3ZunsOKnJQvb
Vi0YAYK9k99gw30grkiOYdb3iEVrohtM+fPEXL7V+u/0TmZpu1X+fCE6vnlu
/K3APuS6ne0+kKiMBOjm16AANh228FnAWKyW7UWaNsrrwwgNMZqi2BqO07Iu
YFV7yGIbaviRnYt8ZHaDTObBrmxOakUa/XDeulWYTNjcg2dJW0ITvQZO8Uys
j+e5apRzDZHp7KAp+8TPTz1Bex6k3KFRy9HyT9dXaPEtsg7qaTjph2c/WAF/
dWKwLEDmo2eTDoxWZTObHWXTn2CzLtms7bMdJ+VLeTdH0b0jaMFsz+ij8eRk
e3sotvFB5mkcylOk43uroPXiw18bAk5cdMFxJNdXXwbeGlBmGH0PxmH7hUIf
FbjSqzPEWR3ql0Rkl2chu/PGgt/iqAhDRYhTJL64F5sNycdHU5loFX18aQHZ
GpallKMFV7YZ5UTAEFvEhhpRKH1ll+5nutn7xi0QhB2f8qkzm6FR0mIx9x82
Jv/zHKoCE3SqrYF2mirVQjOCm5Wwy/FKWhPgIs6z/RvbmWG69d+wujoYu4FG
BjEHwYyk2+jvSQxg01fvXbEnha02ThMTsqGMCpHNgtwJCpZwWq42LoqYA5vC
z5mn7V8xU9tRSWGnrcJtMgs3BSg4XJrW/h7cwk4d163IDTgjvWoIFYfJIN5f
oRyURr9WrHKseajVgJb4le+om6ikepsURGaOousPg+V0pxP3Xplxr98Iijuv
V/l2WRLLNkfDvrQQxXglq9Lab+awMp05AHqrXJdsS3eHRci7jqUrMW84TV8h
PqWI4eti89EnPxQME6ilaQX+xdHPUMADkxssaAqjKBraijFhbMjYSUMN/Ljj
bHIaGbX5UvZH9vElFkJbgiTjQydRjbt2UiGUli0lZfsKhppjWNi/wEEfSo1V
bzVZCX9Hb6on0rBlhtxcaJjihsPwl61ycwSAA9fmw/HXLUSv+HN/57CS/Ff6
iqnF9NhcplPOfNfxBzUITeTL1lCc5si3OMgXbhTQMB7qgL4sgzjJF9/h7jji
xGUYVzJxFKCQabWBoTM/iBjeCbbphBCwUDtM84OMTPToWD8YqiEKvYxq5KLZ
i0gufVxOb5hkFt+BKSsqkVE/K8yCxQtLwIDoW7SwIceZTBqI2ysxCHJwR4tw
wUpOC/muv2urdaPVhrUfAmn8pNv4BicXDoh4RLgCysGjircsWzZhXjFWGpFK
VyKsvjJnNlEkTN/H0tOwSq8SrtJjiuGvR+Tdn0sIVg+itQ8lpTuhRslThuGw
ylBRMuxWcBPC0uKdbC6fWkKwuDce3lYQgF1YgoKpARKY5a9mE89fFI/9yWKx
tSopi4ROVkXMS2Ay3HnoDiRU1DJP1mdXzp+QUcmDpXBMWxPK0JEfBGN1cZwS
+xGMvuBQEcRFLOCL8JKy9K0cl1/BzgSemaXfFbGtyafsF0XC2HOhBYfpvYBs
nPqesAHDxjNc1Je+6mPQTilLBUntc8UK7iPd/4anQQmEfJGvt9DBnE4QrMPb
K3JkwGfP799nTsYjX7S2Wq3BUiY3xXOcVfwkNtE6wMSZ2Vqbd+SZSId86zGH
MHszm599oW9knAe6VmrB8qfBy7duv744AxJjo0oKn3VyLSqbN9+8XychMQTV
aCgfJPF2MjPcz5sqybezBi7w6NMyy49heRFN1iKPy6LaRy4ZxICPkTGrM3Ih
K6ROpR4QhWEgltPSkV1xWfenRlgliqbee1qt1OCwyA009qkaIRLII2GBUG5F
FRPbvD2h2/FIuvdiPBtcZsdzWzSjev1N+f/EG7H1NsrqDLFnp71MoWA70MnL
F15GyQNqvtzFwDpStt2oqZmJNjRGE66qyNga5qPjWO7jAtZwvThIWAnulsql
BxQt3Yb0uZwk1XMWWvxBM65FtdBaE8bE2l0vUilkMTkqjRWzrM24Aq4DpXCt
VNJcNideL0a5D4FVu/RoL1UmHf0JSsfStcqN+hYZqhwshhj4ItFhXMeZK9FU
+iDPNbQCAoQ3jgoCxXKAhioeF9BHiSeoolDEewgEbWbnwSeqtZCsPyBnJ/UM
s5yx3iHh1+nJF3/qPlbkxxGn/1herIwMjK2tUl7HQKaNbWBWb0G7xMW0oXI+
6OP+7kRcboWc2cz1MYnznu8XmI/+tYLrv4Nb79GZaldlXra+MB3nK8u+jgXv
HblmU2JbLyghogItpI5z3vOrhwZjd/78YevITmpc0ePvoIqITxX2DOifFNel
5jVWQNH372oz6AlXRQDWxBbxHZ7CWt+UJSraE7adkP0+gso0uh3Gr66vsNWA
KTYL1GBxUxqtcEPJXJ6gm9rCgvzd8KVY4rrsWZD50geKLFkhYb6/zfGou6KF
OFp10o/W0beLpbEZ7ZOonOcBPjFjJ4VHl1nipYpM2RtGJm1RUhGaW4nzVETl
rRDWFCaDBYTRcdjDuGoj6OIDZTaR1WKgCUDzvW4RwqZQMvOOpz7IRNNwbLbB
VutpfJdvD5Pw6Qz3mSoQRqdwIbBcO6p6y/mZex71jv9Z1IP6gOW1xsc3lcs8
LdBgi676K7Mo2TxcSZabf5XQYGV492WA58Xd+iGxvSmsc7RwVO5/s48tIocs
0cLHHt0LLYTQXCbSF1KdXLqUEBjK1k0rzXEiYdum2o9bn9Md+UhKkxnMp5G4
tp8ClTgcoXQ7UrZBclnAJ37Fwpm48iAVy0auqVMZAmpb4m4dceC9/YJf0bEJ
UbQ7MAI3giGBICsL5+X35e5sy5myjszKo9OYCiYyz+1yXE3rcsMgEiszRoE7
+335I3oP30eKCZFd02uOtX1AIoa3BgmPAmC0cpuxacJNC2u6e7uRhozBVF0q
NVPsamb06UiqoIiD621EZXzGthqKyTjd5xmSLl78UTZKiX5Km2rrKJNfVEcz
Ei5woZa5U75qCfPl5XrCTY+dNCJ7yDYAo9cJmRBiVugtc73fnfhuvtJB6Jqm
O7yYhmdPG6XIZDGfNLuWcyIpGT8Mqbkma1S1oFjk0ZJoEE3PD11uuT5UQbbr
0XUctyuNpJ6awHQsrP9WQD1+0FI5JQoZ1U7C/kZdfbc2XSx6XT1F8FlUde85
Plk1ef3v/0Nbex4Gq9xNmYxh5JcFBcNVID2S7RI8DVr72Ri2LYoHkhOjvgdT
5PIBGvuK/2W3G+80YrvdgDYhDj7Gg084rXdesRugiCP2GuL9c2e0efPfw/PT
M7H2OJ+TBUwjm+ICsqUkqzdk/9C5NyAr2dkngXOLxyyv2D+FCibViMNhqu1E
pWk5QztPQDGGzJbcnzHwpdVB+QIWe6UKdWL0iAyT+MHnzok9xSRckSrR4PSO
2zjsRYDbudSlDmgjTGF7dvWGRAjj9/fX08uwM7AlisP3XMPJGAKs8QdkklBm
pWQtTpInP+NaPbQ1JidWAyEPSwjgwHRHVisquKE+3V/Vbho1x6+5OOiOndz1
kJuqV6aU2uhpHiU3a6eWaStXTtYaoHM2LxjKMr+JjaLjr8YeylVBEgMAYrpL
QU4Vur1ierv+ygBQrD3h6ESL0fYi52dIhL5u3rnQRFvNl/BBMYa1yxqj9VBF
qJKRSeSyE/SM5Amjmbjtpv3fYL9pegctmBAu5TGrt+AhFuksuAA03b0zXcFo
zjvZNRvsyoAX8/foQx6/ljrZFmV3OMhrQoWkKwTrAkhJ+4GDAUQLwfQm951J
ysmKvEX7O/NX7VZcKkX9Wim4T+jhdTK8xYyul4Ea4Z7n4SwKM3k2MnucLyyT
wAebZduGnjGVEKcGNRRGX1XkERCROp6kF4boBI4j6i6D672B/mT9V3WZmcPr
PIR6hRom8FQ++1BkRtuvHlkqDZ1G1dACZLLwlLYoG3cp0r5hk5LuPc0ixhdu
UlSVXS6Om59sN8mqKv0OFBrwSJt979fIeDJ6CGfTbWAoEsSeUWaIbMQ9Rzwv
5CUfNU+XnG5sVbFfbMATE8aPGgVMCuxuH/NNbo5Lqj536EBcTaTK9RSuZCbM
zZni6X3NmrLUizALNF6izVCLPpUg4fk4EG7mpeQET5uKBGgJxyI47jlb2iKK
dIa83JO/MOri3LBawHINot7jakjs3GU/T+FoC0wrq72jLbMveDWX69gyfsmj
/yo7iKZsAsiel0+/rcLD1UszdJs+GwGFg8T4YyEcd3W8nAfEPDV72t2TeVkY
m+3ddNX2jt8jD3C8p3MRpZKgtnB4bq6ag0OnF/6gGKcK/RwbgJThaoPUXY7z
pVXdfTnwSVSIM8ZojAH7gE4r9oS4DhOydRJukKqlhdV6Hqk0Qzwat+991nIH
VMwd3GZnaxHxcu+wrBFg0EorycubgJMN+xSSazNYk0dsRML25qtywdIX4kp5
crXFYKxfObNxCk4YdAT4hwPfZQnplfLhILRAb1/amkx2kqOH7DvHMuYSakjb
E2AoYYenfnSx5Qytq7uJIen840WB470jjSO9wi6N8koOkJotZ7M4pN5lc97w
TRAddi0jtOhivSVJqp/22BdGMAiVMniIw0r11JB73NMDuaXfN1dkQqHkIGf/
1+/fVQcEyPEc5/vtLvHRR56C7q1PLtlU4miM0CE60WxUgRyZyZS56VNp3pMK
578O6UPLcR5bb6sZOfIVIu26RjuaPVJSUhBt9XZktQ5RdK6QoOBWiR0uzgqJ
Y8u91lL07tQDWLDfDqDglSpBmHccwYGbB5Qgx6FfzX/Xj3babsM0B5FQT+hV
GL04DaGy0MNdmIo4ZhMrIe8Fa8fYJH/omXH9bQXaAmOP1wuNIKOjy35RaRzU
TU/g86tZxjNr8/NWp9tC2zaE7fbpPF9DcdDs2OJx3WJ5Ys2SDqitPOQfRuZ+
0YGydIAh+kOAsXEw/Rzb/8VmKOtXC1hCwNBby3eVY5izjkl41ZAA1XOTMwkm
GfaPcA1QSQYZ7gTtR34tmlwzOfcI72910W+8kkezj0DIFhnseq+BMG1fXPDa
fXlHhjnPv4FeRwqCtjh/tO7dSig37EK413erRC2mghMM4Y77c3G63dIiF2ri
c2OhVKkVyeLrZeQxN3n0daaVzKSxoFnRoU29OURiNC6tLThofaBNjLtk+5Lb
m/lKFsRQrVAvevrp8D6Ss7+zCTSCQ4ZLKQc+4bIc+wlaMWLUqwtLTRazVhBN
uUDoVBGno2vA7pco7r3RGKHPEMdeNhriLy1CNWsvw2CsDwpyCSml8zrdo+ik
zHsYoidN2Kk/WjzO6EJAvd76GN8Sa3otu9G7ubzRIlqz7iDnMDTwOwHFn39m
+TJ+Wl/hIOJHiKSfdi5hjMDSDhkCsGPtBaZ7f5kzD6nPz2TOwvD0gdwT54CS
9YSY4JHf3jcE/tSZXAmFWrvJNWW2OUgO1fAoVavvpWBB43KZpTtoMUebTBRe
uSSUCp7rHCGcISLz12wfolPjmLWXPBKIhLUXd3bmlWu858eHKQhzyqUnM7pM
ST9zjXVV0bM6rgGS8T9+enl4ib006f+58GS9KI1NajfJ0mYYGlek9nYo9nCf
MhtIIHW7XCfrNglBIbxDigHFiBZLv9p5qf8/4+uvshQ5u9MuELPCdvWkKVKe
O7SE3NUcbq6w9BBEoN/qaZhOoVxp+R/NBAXw1uodc4vL9MyAhC84+Ul6uqub
ZJWeRIfJimOZ63aI1QeZtr5yjw8z/G0TOSlra0E25cyr52a2AwnB8sYB2dp6
6bThr4IpimFl4fnF9qYnjhBRzp6KaO5InBpiBglgA8Jr6xHxd8rLG9eLHnNc
NJ/7yFv1uob6r4t/SWV9uwFxtpQUDEpbpdtMFqJPSAXVRvkILENlDlC3+Bmy
EcTf28RwuzVffOeBi4QjYWoomAatUSaviReZTmSawaKJaxKNBY5BQiZ2tF5I
yapenmHeh9rS6lTo8Mj/0ecUCFwccrxri+FIXbWLuLXWTXCEEGTg57BIjVVg
jZxClN6PJTYINuChjlOqGBNVjwIVAAg+SdJ18/TEzIaQg7B6UIPb0Myi83Dq
KY9bxZOREcKRRhsn3zA7FLXTKcAN+/gZIK3CQpWgjhG2xJGUqPmAvVQ78Vrw
tbJkNYPo8MmAwoVUxZdZkSnWU6XrOVkEVNuZQmSo96l2gPs7I0tBbeWjqRmu
oijqLMjO+XS9PGgTYZlDrTF8v0OZjXlmlLfi7sXJjd6rEsk5RqYN8HC6Ey9S
IIvKzdp7LdNeAQ1Hg00Hgyde3oSFyzLK15xD2+fCDUzBgv0QLy5ORG0aH4eI
FSsgqnPN53QmtHa6E9duw+NJikkdygXBVI94qmjlF4j+Cn2mAqPFNiYJ0kd1
XA+RaoHRu/0lRhY19q9TowsWgZC3OUwF8LdyJJh4nU8GF2/PTdqaIh8ssmDK
4iRS/q2T63HXOOfBR5LNNvJ+2o0jYAhjTQdAeruJnxtvUF8CC7gDTNzQdIMT
LdYHWMwpkgqT/IVe8DUIAKNUOD3nRT37U7yH7qf1NozCV/SRqujpMhZFmroZ
3/eZYx6gp1vOqk7z3aM+D7dD4vY8OlfatZv32H5Y00JzM9NmB82vYx0cjm+F
USuJt2RfNYkj4k+WKw6iQM+KJ0RLJpxBI+hvj+odiLYbqrYpj2I1G0LDZIAw
shAeNufuhvJfarRm6hE/Jy3oq17jRZyVf8xekhhnVPn3gV2OEEnCG8u+tzU9
BiMm9QdKgHKiwQPjZ0guttV04WXkn+BuqN36wclXJGxGVKkkwsDv7fRTPC3J
IJOfyHHjCBKBjIYABjQ6zYCWT0cadNbJ21lW5fdvQ0xKhCUeR/2mw9dyqda1
L6FcnXcySgn78KpwO1f2RrxN7s6Ww+lzTBVSlGpS7D49hfkeZHHBuT3xHejC
4BQd/htxm6ZBwwnQhrGLHXejAWryrCIiTiN3V+vpsptOetAqYXoNgkPdk58D
pGZBOMgjt6c5opzxVxtUG0632z1xurXiwcnyPo4SxcJDjhEyxkoMzceFtxNJ
uHIKdCUYaeiqZiXdliBA9RB1WshrvlhX5GVPpTezNO+MO2wXHfX6nPTSiJxL
gsI6j8pqomcfBrgE4u4dvYcabQkeipe/ylixfpQxQNIx7AkS/vuW7Y0hRj6M
v8LLDVFb1tAqrQZCHk+ZmL+euYNu90wSlpk+ijWpn62i9x0ScX/5fBIH+GH0
kl9aGtS9mgVvjAt+db11hEHeKvQcCiXERIgyHYJfqcE7yiPx9dYdbITbP+ym
uXSLglhFOSvt8sn+nS3jDlc9o+q/WkhRNKtMBVtVANiMjvqFgKFVhNXIkr3l
3Y/JUyJ5sJ4T4SY5vBfeD6VURu6SjYRYbwp+V2X+mA1dsScaAol0WLhCPmkR
0cTqJjQggVZPmpx8BrYwa7T3cfA2WUoZVX+upxwxwa+cFrBJkFJe0P4tdY4p
I1gWyt7MoleDm42shOpzV7w+ncF59E7tFdW38F43WQQoMXJ60njd1STuE9Ke
mmk7Kmgwnsj+HTrbAjt80dzh4t/a9aE91JDTe2kzTqmDXVKr8PP1ds+zD7Is
U2yUqfQ2d6gOfWLT7RjL3DuGE3N8yHtHimPPfcjLofHcS0ciFrC+BN9Gvzbz
VqqfUvIxpjobblwbcA2ZDPUEyFBarsG+GVRNJbNo/wHPSQMoI12JnhiB55oX
XPrfT2FtHlilEi9mcqjgSCLZ1yVlLJA62YzLeAnmUxd6RNPebJxJTnbAdGvE
8fu3ygUt3ztfeO8YzqM23qZocckQC2pVnsOeeoYf3M8aQ4IkNlysg0w7pkLs
eLWxAwUl632aOcSggF3UONIkdv+5+TBuZPjFuU05v5fktZE2+YGwb4kke8as
3GwNqHJgYnXDQiFssc2+WwrZ5a6y6tZ1AdjLWrMVb2cqSgTKj7Y1+cB7TJB5
83Ivp0LhNm4qBM3Xuq/fr15mLtBDadLLvnvEjlcUgCzrbTIzKvpLF0tIlsZS
rlm4qvSMxBdsHkzshUmGPRvYpaou51UZ1+Oj7Ake+2QIuLFUWttG1t41JTLG
mUnsSvyHrrcG2558d2M6KBizD/KZUcvRejB+WRllZ6wnT7yaepOQozMEGDmE
40WX2yX20J+J/wq9bj2af/grtHcr9UlMa5T+lBsK85SIngtVkl2+vP8bp5Q8
xoeChcEKVGoj+BkNhbNtBN9gZOAEckBq04kS8K9ePfaNHyW+8ilRiTu2Gc+j
XgMBMcAh9jUntNNgc12RsPAWsxSyy2pcD+qDsX3T+LDMGLbcBQLkX3sbThj+
wCa7gUw5IMGQ5C6PoMxaS8B0wqkqzHjSb1GR8408VZe3ZJOKC2owHjCtULlR
EHcwlh7GyR0HqsA1f4ne47h8qRDJAQ2P6rVOaUCPlEi6yogb7SuQUiOezyqr
Qp+FmsSXbZzOlL3YcCGhy2xUWU83Ed+/vqWx44yTU/D8m3CdEgAZwBpzwgDY
SbzKD5wcJlqRtTY02fiRWY75ubvShC5vXWmojTuCIJXqwyKiv1MSXQMEZdyc
pstI654MnDWx/pc+jUi/617YzDydzEQokSSeyaD+rBPGhvtWdWC6l2GIiO2q
0gGCm1p3m70s48cAR7Zb/8+/O+npih1AUfqxUGCGRM8LfzZtaRUhjm9kcnkB
jfbfo2zeP/IpJuDs7jxVwnWteUEs1/xSMxlL/wqc0vZtS0sMW8flxY7HzpO4
5L/4E+Yk8/jjPCLWdISPhZo4v+uPC2eD6jB/9Nocbvdr3/21xg7WW+0Eq5fe
HUAReMkfsJ3LAYrfp/hZjOH5HkUH4noozNmd3CpHbV6hBnS1kLnNK6tw4j4f
Ibixf14xFThsqAiAGa/WoOKBWGXvOTx/E8CACRpqiIBGCnXvY48ho9SQ1mCp
m6fqRztA83rICUSst6T9AiRR1lm/V5xqPAKmydntS+nzFy0p23v7sHy/viVR
4LRIdeERv8f1MsSQM4VMH0tLkBEriSr6ieu+aqKjlF9hkTqf1onaibZ8y1AS
KA/K7gqmwOyAsBGF8bs0AE5CEDHiLQ4t1qp69z/+GSJtuisYg0MG8cd8M5x/
/kBCZAdSPuW2lIQZtzwojBi/X8XBc+fc2+EDbrOU+Rgv9+geYFrMimExipGl
1Y2Xdb0CECG1ZPiX4kaG69+HRlHpP4o7+wEH/2l9AeBTGn9//cm4iQSa1E+S
cWPZoK8M1D7lqxrRRErpwjyIxx0F0Ab2yF0g5f0Ev//loyzXD5zxVClq5AE2
XHv/wQw/Y2BlTUXsrouM2lDkPTMmR7sTepSUUVXdrBLD0iWA9uqEIg/4frVp
WEGCLRLtvV0BsJKgisnN5J1wTtE6oRsX/T/hbpPuFaquHYzrrev0xyaFzC8a
z+KF1DxyJj1Pca8LRw8QvwO0KDVNNk1XVjKLif/3UuIADjSdkSfB3hj7ctGz
+x8zOLTQmX72IT4ne85tbEwUI8tHa+DMxZwwEnnaDPJDUUvw7XRrqTjaVWlm
pGG78Ryz7b0rGG8YcfPsYD8O2K5fUUreVWBihK0O2y1kDN2QphiNZwhNMw8j
8OSAdFI3g8zivlWamao3la3o2jTmRYKXSqOTaeC3w0FRjOdEyWSCcgiKFgjt
eiDdJTuM+Iw9mAvMhksGjSdV14PO/uQfKW5wrT3vJROotcRiUCUjQt6CEqcR
LyKbbJlwzFzO+aCeTnKlhS6Oa0MLAxohbtcZJeEtD5ewFVNOlPMdU3hNxdkS
YC9ciFhI6I82nqX5d97mdLEWLPu2uEDMNBIJXFkLoYCUr4V3T/Re5+FqDQ8o
Hmh9i+genivzqYZMVnfgaJd+hU2QEf0FyfsrmwewQIYtxc6xi7s09/AGvXam
EtMfv+GUk8dEPQyIZ26QlySKqPbepLvpW6Kep7MBAxHq+aJ5etvMBq4dlSdO
EY8UCg7pA0DyTJNpgG+/UQK+MOMH8Otj55VgQlclyXY7eOdQPKaE5ojomOOt
3ZhyE3y2UYpBa/JxDMi9hL1ygyLvTdG609P7AdKm89SPap/EQCP55AJcSc2i
+3cx1hmGwuwz7A35DeG+ciORb4btdQTM2UpKncphHJ1F3XPB9stE9MOk8RYF
nZBE3USkwmM9842Ai+xwJf5Og1mQhI8yKqpIVD6/6Ga3Lekazj5Q7tAk2gsW
FCIRjHlceL6llZdr2B/KxUWNX7LhYDQL25+NDtbDvLbZWZuicMu7r2mTac1F
0MxIHMZHw8Ig16ramlg8oHYKqXnfDOmqd2UXVDV6U/EM1JwF8+pZVdKLc+L2
y0lIkYprB8kuHvf8Jj6S1emn1ypvZpMsKpEsmZvOVT057Ik+UBMD/xptMcsS
K0oyyH/AzaYdQAMwoiwfTK22SYAIJZV7KKiQfAemJ7gqYuRO+JzRiGSeB0t7
RUcwu99/aZAh6NNpQMva1pmo7Z3N0YVkvffh49tCe9EDiy0m7jCtKQs1R/C2
TCKFQSEtRGgRCxViFgBHAu1zGfa2GRJ/2IjfETOMf7oXNfb1NluU11z9qXbN
krnQhMKks0jQwh2jrnygmle4ylhWtmi7GpY8Irt3K07zcgQko4h+p6ShVpfr
iePZpbwESjOpm2loYWinNHuq/6sYLlghwlHAN4qWvVDvY6XI5RQXGOV1GgC6
ilu7lPeGkaTNzO9HRk8XNUfy0mcMj4osx1K9GiNMTgVf/OjFtcQaNJSMfV4P
D5J2uALrASvaxeXinN6tf7PqF0tVzTY06tbtl1BLpl9grr/BbbDeDVQ5Nd5z
M/vgPzzoyyKY84wDvx2MlWrnnfbucP+8ABST+suoJShMQ16iFtpmRyGNC7ec
/MPJ0eBuOkNQ4Ebpfs5oSLrmg1c6fnM3PTLOmHw2e5wDeuTiP1/NANWYApSO
HOK5Nt2wNejhTxKrYtFuAdNOb/KjooMleEq3evCKkhgM0P0RJRq4uonyK1v7
RCyfZFiGy7P76ad/hOLLXoeRdqQMaM2i0vzvuaEU/AYZfAXC8v7JaDtSeEuq
0KAHqMnpa5KWQ9cIy4i9icwQftwpCFNEP4fZH3jYSQHVvoULx8IRy8mLebD5
PMZUIHVo8O0k62yJQptJ8YIyPWxTkc3z27aMlVtFUSRzeb6miDXWBwwrGxLB
qvWc99e34SAJkiO8Y3IMLbTIkbM/aV6zA325Qr/zSacw594+8eqKXt1I2mY/
yq6qTJ3cmxM9GPqu4cyRCcPkz/1wdKuU3bd7MKp/l0zmm+uO9i4K46fcLZiA
ZFqeHbkMVB4qs96zQMEpHtz8eBIUdF/8ZQt9irPiQgtCntyD1Bjt8Dk0CzbJ
fx4IrUwLuzZEpoA66A2fBS4WV/JxBNAARllnyrKsQ2zh/8G+OCn8CpKYEzg1
RIuKnu8u8QlFLAiWWL/nM4sN3M5HblT1YeyCvWSyjzuDZ9uqiTyialtRB3Ur
7QrLjg1uhPLH+QdH001QA4/ULRFOvKwzhTRV9o92h+4kOMempY2ArBpRNJJa
xS/mBr/ZW80dCD26iRZPPP8wepH78c9uJrKdH9fUaS7Mjb5DOPUa6sKnZq7w
2bTsfbzHaJIipLo22mBb4EH6vqxHkd5wPnJpsekdifgRH0o2zEJjmxFcZCAm
5i5CniwFI8YD9h7LcCqoQOuPJITrfh8Xwl9XYbFSVjIS4HTNNHPBXUkOm39w
2jZvWbq5qslGnGqXnQzvq2c5mwMiKz2Khl5011cC1Aq8gtK2/Q+0h5gMSQm/
l8oPs/zJYPelckDp1CiRQKLvcMDCN7td//eREu4VGLnlFDQDzhjyjIaCdA9i
dH6hKqjMxsjsScofJQcEkGkMEV486DJQyrMJJ2LG21RtMMvICOKNoVOd7Dbm
Apm26EbK0Mxeso+k2L7XrZe3HgNzC/P8iqV4v5BpVP/eKM1Q7Ep5g0EgFbgj
TPEiDHG5MjS9PytPjbd8YO4UG1ZuqHNAiXoKf/UgUKdNJGEGUGBvCzpTiYqI
jcriItUPDFf4lUaXy0NNy9YDqiJnXkpEI3Q3u1eEY3DAdo7ag8D4YONTzKwg
S02rAGOd80E2Dvjt74T2wwFpx4PkG46S56hwqPFQ32JKPFrjV8O2sB0OQs/d
k9DLj6c65XDiI2PBygof0aVECn8NUTf2Xk6v2g/W+qEMn/gz18hRPadsBx1O
a3iFnYgjPc3uPC5/SxkA982zkBOGXvQEPnhA4nx71e/BwVd1mDNKyeEINW2a
9YrVa2pZR5T4y8glthCoHLr7B7LZgNFI5JzBfIJ18gfTKuLPNMr0qysPNIbr
Oc2fha1rXic6CWvVclXyw3BtUGWUrrIDTETBAAwb1+bnRL1apcBZwafQGkPb
45NZpjUbjsOjzMo4v/pcweSKrqYLhRuNICcdcw+U6DmgdabX7cTpvWkzJ+0p
mynZuNcRQ12xf9eCeKd61KH9N6u2Yu/uFvXb7x3XYj467II5ubZrWdZC+N+x
hOtstBG+oPsT//Xb5PBuWyDbPBHBFxNRlK9XEGsl6uRA9VywqxGpX7YTtMH7
GZ9fJ8nOA9RpnQbwy8FNhZhz+ZuTVVImc4UKEyV2bHUrLusaouguOnZGcKYi
H0SBrj0xcjudCN7XsnhabouH5rDK4T2BYR2AzUq3Ckhw2d4fwcI/BRAyYN+H
f+rgYAoXikJKx1JpbrOnDqecfhrRZyeEaIhKxVLIVyuwucGIVbmRsillz3Yp
51+jf6gqAD+MhJKz19pjhr8ayvkLIGRTthQe/yEa5Xoc60P+e4DI7S/hG5sQ
1EA07WWl3fJoKbcLz6iHW8J/QHL5rPSSOs3pjubscH2yBnfAQSiOHhI1kKgP
mwXG/NjWRa5utGXeG8s3SVATQDv5VX/LJAS0FsEMzYySKz464k/sSMTd8bV1
8Y0qWasNjNNANL0aV5LI7gsosG9yx4ZePAGd4ey+QIJa/tnglRmyseZt+2EY
T3tsogfbsUU7ueSIffUQ/CgJMJ7pgo3IloNyJT+mSgWfnH7Smy+IXlYbqLzk
9UofwpHlpZut9ReO5Ia7s0VKN2AtKNcwNf725C8pagayAvb5l0Q9obfzmuQn
j3RZ3mqDtWLHhdcAIAT3vr8HZplL4jMzi2ysLSeiIl3FpqAWjC8gc+TZSf+T
eRrR6c8CjrzQZltKMk7ir+pOlx7nLQaWXIU7CeymmTz4bU7inFW2SOsmlWHM
klDwPzI8Nil20JStRM+yAHsesidiVMmiiiwqA68tcMh0GNbMKZxhHX13Wxjz
lwSa30kThGPVvUDnd4yZ37aqTmi2ufKnBeGUURLAVBEtRAp9lrz5DQHdR9+U
PwFWeeT9iSl5Ihu+WiB5OdBfXnMOiTE48MQD4cxY92ylG42QckvbY44PNg6X
Invu3IqZ2hMxlPRdgl8OK5tKMFXjS9Wb29AYxqaiwXRWGT61XrTqOoY8G7NI
Da/yaY7GCFno94xBhfbuk4i74nfJru6isooKUm+3YAgYIN8qaAmGwNytB125
75tDcvhPKAEv2kJthk+ReELxeVmoa7wNyncYppfRUTuzuPYXjxLD6ng1E+Vc
WjXLdmPbOmHAU4d1lGlwVbST1EZTo6PxbgLv/PPlfwKXUcvp6GXymFlOKRgn
LUELVQoEMdY+OLRLXC8ehC20iUgaegz5v9NuQk8KevDa3X7LtEOXn4JXOuq5
lLeJ/YEV7Yh3OBWTrjmGgjQXpCUD1sFq1bwwPIx+YX+PUF+BUlFkYXrxSw5q
DdJ2X9Q0xSl6P5miHbCehqifUmQ3k+xhhQOKyg/va0eMM/PlRKV2u+LGhJRj
RMSAeUKRer70iof7qJIuWokTaBYezChSFwPyjbPrFFzYU6lU5fIJRDVqd/nJ
/waTiDnJtUN8919wjJmIekWuReCZGrNn8l9KYAjs1vi3fngSNnJfPuIUBBqx
4q9crDLYp7RNtkth94V3372VmZ4pko3cBsryM4/Fw8hBgTXy22t4DV4xP5Rq
J+8jy4lm0j98gyySjrYVuoEd/B7wRmroEUS4yI2f8+0WLhvsS0TFAIRpx2CZ
6VAkMZ+mbLw9bvoHWXaxjd6iTK292IYH4pfhsMEGPyEIu0O4y1WejfO7muUx
xRqTQqV929RczHGXlaCa8IAbX0fS4aiwP6YTMrri1GSmTWYsCLwFVemyZiEW
782bD0qZGc38qd4zNDMqbxFH6V/Al3voDV1m4CFojzOK2LmAs41XEHGfdhmC
3Zm3+4RqSSX1fKiCy+c2hC0CsmkFizhlQ6DxIvFTikFgVz/0MhVyJmn+fNDX
DRaubbQ6knE5SBhS4FMe781WRR/CkkDcUZ/ETdEnWmKjzkEFD3gtLsvxtIxY
aFsFV5ffp27VJsThYpmtiaD991D49ZCmalrFdg3vPVGyov5AkmZfWV8HnWHS
Yya0Y8d281CIH8h1GzGK6koY+7/tMsMj1wJyTDrEvEgKAn/1fOGAv8csUqiD
LmlwyAMWUrkdiQVuANTZZjYeauVBqLKoB+DCUTQqmP8MoJBsQIED4K9PtO6r
GLFzaVJd+TS7RX1nsyo5wSMXFMQ8egmb2AS0du3rqcWuOon2dGdRXHw5886x
ZGwf01i+EnKF2K8cxVGDjKXM2ksQqHEfBt67KP9uYYQS2J4rVb6UT3X52pdt
fLlP6YLWtVXOfsUpgGpFPVBOOXcMNIbWTTySXw41plOe3HyDbMMIf0YZDH74
LXZ4+1w6FV4Y8t56uzt9CUbs1D1hW7iJUQm9opFy9OK7LskRIumgm22wbc7G
4HVpuhLNZnGX+A4c5pnzL7xM9prkfDNs/XJ2OzbtRsJ/rekrnW+mhh+It4R3
dB/9dBLs1lF5m62SCmgz35rTofy3pLtckaHFjwv1V4him/nJm5mDBF0S6ByE
qM6QGgvUXi/WcuzrVDJMKlpVYBD0NlT+29orHFMhHr80WErnIMMhw5azPjWf
czToUodkfBJ2FNY4QmwjAyS7OtS29HdvcjcLDUxBsvo/R0e5jW2sz8KFpahg
n36l1Uyj7ZoqOxOXn1DzqOBjdIPtKpqyoKyQJrZs/yXSw5Fxbr/vv6GjgVyA
PIC94yggzAB5dUN3j8t5Z6Dw4x15xdSdEijuXdsRN7n4JjMAk9Y4oI9hl0dj
OGr7xA6giI8hqf0cuwS6I8KjRFsM2PU52EmXm9PYkeurI3bmGArrHdPfzYYs
DZbjD92FSoRV3BmlBC3X6prPjFvXdhhLo1gS6bOxEtr0/LLmBxqa2TS9WFIn
yw0GILiCw9GF03xKOcUKvsTRoKQVJZwenzZFcFLuleSTSjqw9tg9eTN1+2hx
sLwuHma7Qt4/IPHOwrAVWudjZLmTa/Lz8DKJQSGfi5eVkxrpTZB0vT4hn6Fl
t9OnlSaE6P5XXy0H7U9Gn9IHU3Ct8ym0fEIhJKE602c5xAX2aNtRi+fbFKcG
0CGsrNzI83AX6Y65rc0pBZ5SbL9lPIbJzTCdrOyJvl5XcUqm5TQzQG3x4cBY
VUqbXMwQnwjii/zfVdkO3E7YXi1BQGyrLzUmn4Gd/k8hCB8dfb7IBz1rze6f
F+RIvJfGRTvcF2PJ7PWh+3fk0rgg+7VqZ5F0B18zjOWMcK+7UAYyasvpoF6D
MKrtaCC2PBfbLvs3zpqZ+scvZnbPsGnR3c6KEizCLfANa6J8UGZXUv54WG27
J2MFdyAFVd1ocfNO2RJXLclNcVp4DYX1UMO3KG/IqmKYyiNOFS0C5fHlcsAg
Ojf5IbelkFCe1Kn61FJq/D/S9DErAXlfm5GHgtuWlNqKrFioCdZ3Yg2SdVkj
E3YtSra7nKjAHnLHaU21OKL1pI15ppsMF2jlc1O8Jw1n+islcaWMy/60PpL+
jd3N91SCt1EWgW4NrbNbBIyeuWoLrvRUG5mhz1Xzdb0+wLvei4+ZOEKDupb9
IaEIqN9q9uYRJPsqAbyIRZebK3yZvR7TWL1CZ3vBx0IhkQJk0XZMszm3KeZb
JrbD5w2VCOONdV/9MTKNt+DOVfRUQ931ZXL54kl82mxjUxFDU2ydWEQenBH9
TT2ghw2kO2MdRhJqO4Zc84qMN1nZFW8zxcaYlwimFSnvSoQVHDI5OB8KlDi4
5TIh57XglG2W2WLy9t3dVnEObnoBRu0HZ6KdID7/SopgTRKP6GEapA8T6VQ6
xQhEC+qglGMCxG95JDe6Z7Tj09RDkFGS9IwB1qaUcwb3hHm23LUjbLxUgzbu
p+S8+Qn3FH3G1k5VLh67ItiydxzZ4EfF+0JVzTx68R/QxpXwtp2gDCp5uubx
GkyzXK5DEqo6SOmFBvYCoSoTNC4RLCDU4kBG2cduiP0QzOUW9XELBr4ZaiG/
u2iol5g/YokIKOXkn3Pr2SRaUj/gOmSplzx1RSgU7G10Hl8bwbjdSlCC8lew
nmonA63D/h03Wtomohd4GFUXX9JpYDjPBPb+59tgbmD1LJfR8eVlned11ADz
yldTf4u/X5NRuL656x9rfRpbymg+sc7dZKjujiqqPhWFlqXXL1IAmesyVO5w
QsbMmiLASzWEjmzBIhQLDHWdV558fNOwS1+QOdmyzMA6fqevBX6hKTFTABvp
5kF7hImARkDYrBxHNCkW8le/T+X+3RzNeHP4R8btu1mOYWyE4b4/u0nbLSD7
Lu18F9vBPjJeFjJTEVh/pfrvFR0puU82PRuMhgBk5yFG5jIoJwvBkM13eAkI
YiDTKnRLHvcMqqwXz0K7Wif9HNTNBZw9aodF/1+fxZBUxDAAcUBQGCpazecp
ZNDJUC0W3CNO8N+vcOwKseUVsJsevxfHb6PupuyhtIy+fVBmCRDHLWBnr1J1
tFRQTJ/J6J6RGWgTE7jmS4kx3QVmY7tdUzX/W+/TgJgf44ZrzBC19DaBj6HE
tkCDYaOnsy8fPBtwckS/nyrli6sftY2IH7tx1UHkjC3yOI7masEUPBe8nW3u
DowqdrDGzUkuPn/bQskByb/TPq3e++4vpt0uiT+7I588fx2hZZ6wuMBG0i4E
+mSewN0tSg2GZ5Z/DySa61nJGk27bMlwZvZzrj0WvB9VpZSEgbOsAyVD5Ol+
oKLMs3/9xI9pTBQ9UoNMc6nsk+hHXrvzTdxShfbnRNgIHjUbgYdhOZbQyBPm
+zw9P78etxYJjpL64GVgNdJTKc0nsfeBSU+Zg2M7z68Yr64aYq70p748NiED
sBP00SgKAToHwQ6zqPR76+gkmunXECtABEvOVCZzHbXGAZRUo5QGYzSa2DaI
5EtZRQOtFpKze6cLwuA0yy5S1Kyij2i8y3hWJKXsaluVdwjXwd0nyq7Om40A
ERU4YsX7FVdEfy1AXbBXDmn+5qBIIQeA/WsvES2rN94qxFBlvOwLSEmKCXvb
CDTs068x3lh6yirF/7xOFna+M//Nrg7HGkL2VlyWiaCSAt1jsfhnSLkZJfvu
KV0u0ozI3ah8jUg+xakGh0oRT4866bpGC+jbiuocw6E5HA7AiQVgpqjHDIHt
HUoj25rIK0PHAtmN21HoVSK7hkn32gdPaoxDCZGZctPtIBeBl+rKkDe8IXP1
VZTjq+k0401upWeHwEr7BWgVtEV31sB5VwCqPVaK2aZQZ5ygrcc1OXxmoHkf
Bq934Lz0rs1UhYMZSIBP+OQdFYG3IiwfkxRSRFWxN6VPXf8cOAIJwwAND1AC
qXZiDx9jmCvHkd1fC03NB3K8hyvXIq2yZn3EuC/jVlDXWIg3dd/lops0Btjj
Yi4qin713lPGvGnQ9M9QGL80AKdPexidpa48ubiUsIMrB+sLstWbwLqWYCUS
0vNYngUrU5u15o2M0QspudEOEUdz+cjPTuzIBgwA55MalTUZ+xW+PFxQjypo
4EUwBnuclEeTXBYKfSU+0DXVC7lLIPnNzauVHZpEYY+NSdyejaww48rzJ4qF
LAow8PV1lQU94znIf3vUd1XOSd4HNz5U53rWZMLBUAVuh5BCsGIVwsyEDV4u
GWHHUQYwgud0I96ePFyZaTT2RRW/YWJiwyhkfGnmNrR3eQaYmmPPH0Uj7ir3
FfYaBtO67ELpBFbx+gwwRjIWZJQQPPDq6miye8CVtF3cNzIRYj+tDpLW1Lx1
x5sH6OuOh5c3zZ4gWCQblB2Cm4AZI4qcA5lKlHucoV1daMoq5z3cxvq95GBo
1O8s6RWxwsxwjvCZWubbdi2qRaAY6V7L+5GqbziVz82DFD3fTgGcUb3OiFi+
qYY4cWDl9BuUI1nyMJS9kLg7neaTIflCN0kwSK+AqzwiM3JA2vjCH2mugxXb
49VSKUi9Orz/uIYtRfcQ5mmfBXDZnioTpgSFHMbbExoUYCNkfaAt1arjjRUf
r0DfxwPXFSSyPXFXkqsZmoBABXDIhOR8/xOjShhsz8LPpxjyDBdnr+vwG02s
OIsFyIQJZfMO6YbAbYHQ+3T/Non7nQPLGHmPSdIwTWTggzH8nKPs7ri4UidA
y0Smy44RZX1y7KT4mUZx2YSTKim3NxPrlfpmef8vGS9yNkVa9E4Hza44OIPA
1zOa2VmRPm6aZjf4u7iQussA9VYCJADnqKlSu97b/MvqWuDTgrVGA4VEvAxb
W18Qagm4/p31wi2XyQOOou+GizcaELVhLmY2VoqAWisJ+Ab138KaDPAiJU6N
bHPOqdV/bh1umKYDCW6qqHNelWnp7NR82FQJM1m22s9NGe1rBkjbERJRk4y2
slkx5nSDDGhfwLlFORnbF7oQWHJKNS97Rmy+j/BFzffabjqsKidVTk5dOnOX
MgTTebx7JyM2Otv2p4R/fs1J8z3OgeF0qr5ea9fikjnfMtsyFIy2LtOQ0rzS
ceYTIGNv94qWfGCDhQWpTb3GNs/4KKbTOkuM0fRqQnFloaa2MWZdkMIKzca/
48fr6NwthP5e3Y3coLkCVvj+FghTVnatIO+ENPqVYcW/u+/JuSq3tgP6QTyj
Qit9rJxZKjuX5pwzw1Ntkgj6IMNydwGnbsi2geEeXPAKhI2sHzezVjLHpPij
sLMPb/6BA/tNgfkmxl50XTAA9huu+LrYIRTXMcXoO7/TqDnoTQMYgJrtEvi+
PD81ADf3k6TFomfLi3rNoCwqkBL6RhWbib+LFB54BL0PCJumHDRgHtspWd37
dygvl9LSma8/T0OrKfF4HJXPpfGwcXRc5H1OTlDheEJyZC4sJZ4T0lzslDK5
FmvWlGMkPi9deW+w9mYUMfRgvq51iztdVOtywMAbjrtQEAEMuQOD6j9tBxhb
Q0L2VPyPljQG4HuACuTnSJ2gA55uzrcT93Ut/EQs0cQ+pSdQL+hifoKvrskp
GjvDDOxl+pE4iWKzAMwC48eFCNr9Pc761FA8v8pBRROMm33yIceB1oSPbtLa
NJnltCZRl4csgnCZ1CsSY0gSvKp5zssMhrDjd3ivXIsCAvJavapzLevPh1nR
RZq6WBnt4OJDJprRpWm3P9LjQPsxf5fMyldWWe/7v14fahAMe/0g9gTHxkCS
H5MVixwZNlBHnmec3wjGwOQybb7phvSz1Oo0vk2RsFhKEtLnSz0cp8uN0ZIj
ErJVVPYu3vupenn5D9Vs3OZxX20G22C4Mqv3h5OEAhvEFLOyACH4kB3N+rQF
u5Pc+T6U9D0UuGsOoREGfa1zcBS2/WdKjZo9HRHaiY2q0SRu1uPasq/Ed8eo
VjT472uQR/C4qTHZJ5waHioLLc5cHB6qnm4mKoSN5TBhNkli+RfJXBCvaDgn
XStnAMtNEX7t+JyDgCEidxHZocechKxMQHqktFvFWHdPTvJUnE+8exi5pGiR
tG6IJk2C1FmUQqXbUYwJ7bLgT5wln6F3V0RtiLKbo7ioa/lqRxrmsHhm64bl
1V0lKWHqwZwKuji1c40AI2aNOIWUTXKhsToke64LGsvsAubzCji//BLIwFa7
P1V7ainZRNU7jekLDrS3IHFTrrgosNQ5FI0Xc+vCOTFjJnfgZxUNPiWHvhIr
5Xjg+dqRLYNqoA0Bt67VhaL+L1yYUy74meJ0v/FXFwG3nLtn6vN+hzIoYGbk
2gfidRrrpMrqi4YFbKYHd4ZcGe2xqmJqX1NcIGAiBny/Fbq79DE8C/88hr3x
5T+sGcapVeRATbDdtYViczrkRgJpBvmEH8zhSUXMLNdUGjrhED3lrHd5zyQW
Yz8kjjhy8xe0xSpRaJ/4bTvuP8fO/lP4SzqXkLYetMTgk9pOe4LW8Q8hkCFl
Azr2kqbGS/HrxD4L0X6rWjnATfW97xmtXJ+RkHovX8OA9D15GraKb3guFfpP
rJDROtUupzF2SMnsHgBiTX/E+5Gu46INl8LcE+xM5mnuz4ui7NhQdA+1NnVy
FuI1StEld3ocNRPFS1NAkaSRXsSjcTmCfeagvluI8B+nyvLvoePOZ/zFxUgC
4vqYByrGdsWo8NnoYuxDh5xLoFFlO91GoOMwCndfHq6bXlk5yO83mghRSRQO
2cFfuPIVsGfAapYByvtPrqj5CshbOKDQvySmW509AlDdgNiXEb2L+3Dl9SQc
ETH/n35hl0+GRcG3jnW/kr7vOxAx0rvtC2RwvvoZq4GWf3lB+r/T81ibDydH
8S0YTTdnDoWlF3Bo9yyZ2+pioddOT3msX/60W6oSPWaJ7oUeuUu4aSdLhcuh
hn5EwPAsbOKAzsEgPMnPnmNFO7PvtLbwIYict0Nl2SVqdFay0qJAslFSL+zT
04DjBeouTMcsJRVUCs1ZAIuIlVbbEOcSMpVTJBwJ3xY2vRHxTIm0twe3xlYD
jXj4f80L8FKuw8ord22j1MM28V/uBsmTnEX+7WxCziNYeb8KI7cSVSDyEv0h
ob0qyfFKb5fQXMNgCcI4UCQM0LtJruy2WqzEZdDxIrnUOBnES35kcz1srtnU
bvAIaeVCAjjo9vTNHzDxu2alRjhP4tkJXDV/e+VKP6mdnnqIzV//1nFqQIJe
dSZuZcvhDZRuZ31h3pPKPmiRZUQVxAL/j43U5+BMv+M0kQhmjxkwkPegW3vL
lTfpNUfRBlUFeTi8IX3n6k39x93JDpqnMFdcZvZPU8dIEFBcyK0vrxCCgF5u
4KczOsjubfC4m+Hsl11r2FihV9WVzurm6psK1IsP8scawcCQ7FEQm9HgnSdh
HprwmWESX7Hkrn0mZk7qOqcbzxQlFov0fCqI1yUMSaUcDfSNgBbib2OQ4GxA
l+wEiyirTcN7Kk2HLh1Z+2Hwwq2h9jTvz6lK3QKCwEx7ntDRbdTFqRyepMCS
UpF4QpMiIprRZKUH5TIU2TGk8TvmEAFQQ+rcPr4VJtFfsjFB+mgcUs2Dp97t
1Tqdeam/O7HaH3riBHLojFMSKVsyQgsgr0RE1Rr+6oA5a78En19qZxST9sGG
ZgsQqKs3zLHSeOOcVr8Qtrn2cZjsJoC97do86Lw3xCgKTdRFvL/X45CniRVg
JE72vH8ib9zpsWwQMzXC8ffBsUM8xdTL33n0glrWFI3l6CEahST5Ww1gtmR3
KzLXG6NaHmi9+ytpmPB7wLVgXOsFhcpmyXr/61us9BKOxaEb4B+XC4Wzwkc2
85m1opeaWhxRlD8hnQuAkabMwMVcCRnbELBrdCF2auAjwZDz1Rm4AHlAam2H
Fuk2d2pAO2H5eOOqXiHdZJnfWImuwrR7mLg44ZAOx19/1+fRXGokUKH2c26Y
RE3HeXCE06icTRW1AncVBshPe0lrqbwvpjlnE1xEnJCZj8yTQWXOjpoSXHs+
5wbGijISABfgdJtDbYiTVlv0srCL9JcMvwvR/Pe5kjNNulYCUldMq/om/SEE
W2dmxVZghjjzKMFm6DwLlDkgRh3t4nGZ0Ln2VX77ZQaXDMvadmBcrFD3ZSQS
AyVjikpJQg8llom+6R8EhViqxjPqXfSDpHS7LZe0oBvt/A9mLxMQq3emZAOi
JqXikIwL68PIsuROUnYeVmgWwMqHknxkbSfwJ66VAtWY1U+huOry6pXdkIdQ
WxwzBhdqY8FQ4zqxtLp0OSa3TASIBdeTOUDoQ1g5E7hz0fTodYn4QjcK/XyK
PH+LwlQ83wEtHMgoxQL+G65dutGv7M3vuW4cQWWo75YDzTrGS15628VUvXeo
QSSgBHvDzHUwLv+Z9dopjmmgzxSy4OK7cKcAPLQatVDbkN6w/tU3SJh11oF4
yaLGm0xMiGwiufejsn99iP9l8SrbOc2d7it6dhSfjThBadZc8X7NTgA+QEvh
7Y/hcbz/qirByZDA4uRZ646w6Sy0izoKgqglMMPitkBhH4MIWL3TgTYPHMWp
N76G4UU3vq4ZgjRFxxc2W4SUzrhdstp93oaFfojWgNbsKVNSiADMR8C4G0UX
20xSKwERW1x7Ltm/uQvYBpyynKEoTTSbVtASqXsfbZWLG27e1miOOWF4kzZl
lu2CDTUayOaNE6Rn/9xsJfHoTTb7FFm+1IS8PhGQac955qnybBoYTqX+Itix
hpJ0X9PME52BLyoSgoWNsz/xABNRvW9vsuYp0lu0M6R+ZmmnOPRcmh1WcNWE
EVz8awnj0L1fVqHXfM06s2a5sjtfakzODmuqwksPWOcCDW2+5hwQljTgJo9F
2Zjnvitl2oXaHDpift0ULAbvs/Ca4ENsBVjS6EcyZbf7V1Fciz/mtRTSykd5
jHgNlH1UhsBg+oB5P6tGmdALgJgTbYfoOQPUqeH0KaUQPtNSHRmQY26ziKNN
/Q+vO6MbpFOUthYtu3QrC9dgwegZZl8h0QpF24wyaOpOLQcyXHaSUioUStTj
UNyAZuG+CCBskLwYI6OmpYcyASjb5tn/vI0vHjK08ECQQWX/PkKRWRZDJtPd
adv/reXusPFcumR423+kgjjscmiTvaONX51TRxsKbm8EUUhGFzUEsIDzDAkf
MvedqGi+yGYK2p+XEYATSHTpelNjExfJcdn6XuQKZTn1HIHkNr4ii8XtOp29
6Wp2xt1VxrBq1xPdv1k9Ouo9DqnYeatW9+PuzK4qQCr1S5yx/Yh+eXfeU2yi
lSTTOAPtFaauGBkSNxJ2vUD30tV9RhDehBxpoaEa2sdIAjRFXRC9r0KvUfRR
LdluW87hru3tfNmnx+V43efYpduLCXfKvBMFaNRGngCp2xa2GSVU/0ioPFe2
r0bVXnVdGFpZZ2lCjWAN9xP5MP4KDxdvyMG31eqAx+P8YNYynKUg6NEhaHjH
PwcWs1Xe5p7o9IZBrqB5HZFdAeEmTHoRIH+/B7g+dmANQA+M+Uk/TqYrXaYH
+mDllO9Jfvih9NOrtV3kPEtzRn35LVKCwkJHrauEiDXva5dbE4awhaqQjDHe
GfI+i3qid0KZLVm/BE3/YvTU+9NLennwyPB3osou1Rj7NGGkL1NQxS8h9qdG
irhY4yp0bJFmG5/yt05vqiUXvTby+BTZY/xwOkIKxVXYFQ7EGnXD/Zx4u+eN
teBcs5dtcj0B8Yl8aTJopdbIeFWlfQhLqOOylA/htm3atvbK7rrhbwhKau3h
nWXTCekl7asRYhbVQO+XBh1NV83sJI5HxnVKbgmtf9M28aIhlVTxOsplTaSX
uCEBPjlmOmJ5Oy+iaNb3UuLc0oUze6ERGmxGdHppkBcXnBDrxW8/igvvq9Zz
lMeu/1NKkzFuVkJnfX3N7EE7aSJudWr7EwWcE++t4Sdik0+cVaSjgCWaCARH
U/MWfBvZhVaviAcK1+QmGZ0tmAPiGU3kHEqKz3L2hXh41uJqV834UKd5LxxG
dE9a0/WAf7Ym94dgQSj3nzqadb2H8NmDw1ZxroX9rE5bDhjUixor57GulBa8
1irMpyT98iSaer08oWmDOMaNaYk6YNKblwN97PbjrF3yf3/T45BfUnhZ+u2n
MIpBH8wRVpmbnvF8LfI3RNrlN7C5QR6qusrEbajnKrcPZwgrFqA3lTQmaLHp
zjPBv5tVsKLJf1u2TQEzC6bTxSdS5CG4zXQs3lyTdXObPZNYFCdSmQEEcc0K
dzl20nEYsoD0VcKst7mHnV4ez3WUo3lRE7dN8U2MjeABGRS9q31FAisYIl30
1sP+61VOF2zFWXs8uiv4GPoPUg43C7H956TCILjWBE260Wzg3Azv4wkpHXPg
0SvVFNaVrq4lDhn+tBmvuI0AEW7yOJEzsUGroD8LWneCr9DKMSnzrx/axLVg
CzFLVbwn6+rtCxuftWkO/x47cTSxlgkh7LjrXZzoI5XcLydNi7kpWRWJPkQL
DEi/lG3snZzKE0gFtoUMb/mCG1uX3kWe1wO5MwidnhZZBm6cFF1nzmWYB3jz
MlOEAerd877D/Q/2sAz+GR6EYdXtE9jApj0+2MVQPWrh0BuHduiG0SB6pVzy
lWWn5OpET3JBWp4JhZZVlCYoUGjGtw464JVsq+YmXpmM3nQcm+mVWP5QZzTm
FSZsVX6YQ+GXReBugNoBTEi+jiemHjCVtLk4DXZ4WIF4EjRqg0J2FZCQ8X/L
9DR3I4/lzplsG6MqUndm4JzWaAVFO0JisxLiQsFnLS7MSlRjdNkixsXnnMOn
1OivqqDis1RIIhdn76CaeRpExwKp3HFYOG3uAX7Slt1Nt0MdJRb5ml4hrGdZ
gZz5T6c2Ee/mpUX80o4jJ89/GcprQH7vUYNI3bmhbbw7mdhIIOexVbvQlPQm
AoG79TanSzkOMqn1kEq6JPMFpn95ZGeeUQIBQ36V9CmYV3epsYcZ66cxj4yO
YH64wPYD7i3gAJkRsNOdVwad84deIYQW+2xXVmZ1ZYjxvgDy7afpbHPzAvOq
f2TBSqwkwtn8J/HF3jZ+WW/Knl/R3QHGWQVNy8YMt6SoQMr4WKZujOVYk5x7
EaKpe+oBaXLYnbfY7deUACoOCIEFIJULqggI/mWsrJMHWJQbdCVPnZZlxwiJ
aOaFeadVtmfnrLXBMklxU3IFScnTW+9BsUWQV51ldEZWNpABmwBXrqI15z1F
emmiDfqgcBpNNow8lQa7qAr2CggXC9JRdndA1TSSzCfwBEV0BW5UNnBTClVn
M12cfQ7oAmEHoEzMwtQi5yZTjWzZv3HpsDaeJwPSwII+q9dnQA0jFopH8SMF
PyguppHQI+OiIzmAZ19bM2cKP7jcBSjpUznv9w8Rryub1RkKTV3Fh9oYhJKS
GU2UDlFzUv9V4sb+RP1dbAnB2lPZruJd5hCHVsWWzp4VkiGMKNWY6THb/IUz
GZjKxl2NMpirUEhRjVC0Xs7vCoMs2VTrHVVJhBswkP7MUQG5TXWdyK5zxwjJ
7zGs2qjO8GRKn4bOZanWLNhjjMVfcfrDtLqR8E8B5pEiumSdM4mGOtarLzDY
EBHNx71ZkuFBHae/soUEn0khsSUFFcwWHEvhUtxizdNZ5Mv6Rv/LLqBCK38n
Q6nACid5YUNpwRwjqKxlXOSkFWpxpwagMln5r1qdz4hnK/ufQ5M3X7eHaDsq
/X9+QBQxBsIwR+WrbNmizMR+wyYdZoZD81C1JwU85y6yvuw3eFmuyp4CKDUn
DWQaIuRWdVbTUy/1puP/wb3IrB/OAiaqebSB3jKA6GK1AyupKv+Ze7J3HCNK
PxbMFNyQh+wXkSbW+6ndfL849jIV1zeMHtaRA2wjcyeIMtEyyZPfDy6mOng/
LhCc6DlGzVMkgfT3FmZwNoDxxYjwvkUv50V87sCoXaG5FPu8cFiZdJi0T0Sa
Yzo44k55F2j6Yp2Vw9STahK7qK6VOY7hDelBAxnfbhqicgmZtMLWpJYW0XET
pwW76qozHr89fgUT7FSshvblGsZsbU9d/y85c3S9GBXMVsnn1+CBTmzCChE8
sH+3Buw1cnxtgecxGobeDpt59MsW/RBfr26LOz/klrWrDVQFn9LC0x5maIb2
xv1WX5k4X2D5dKWVrkWpMcmpzl1tYBJgN0VXeJBjYThgOYCaC7sGlz7ENJAS
CikhHeqTU/CnA7OR7xLX9tDfsCSFhCrQ/5xK+OjEGIOg1Ge9+FGlBqcZfBzS
cdNjMcyX9lORFApowzcVxMC4P+rAAC1rbdH35Z717YDCDlshJS/aG0+iFjJp
gw5bCuoXdmUv7vdzQFDVT24DGkJaD9YZpS7r9utQmp8Hu7k+0slhu8VXynNq
Bcp8DAkdemC73aqmQ3JXJg88maJxFS6CZ1H9XKAqA1g1k4O3hZDx6CXBqlHf
3TEjr+4uUo+arJ6A+1Ul3Bvs8kS+le0gSK4a/+wZtR8Tkt6aeQSvbCK2BvZJ
oTmrgNlZ/kxxtNFIBRnKOFgRpWwbprwIcnYTfnaHhGxJZInv6HJWKLy60yEx
3ntoOXj+5YnyXhfk0UCkAC3nJvWOkOspMdRfUL2P/EFq20G/bv14azlwpE8M
qTacCzJVnKQCeQLOeVO1pIz1kxvofY0EMyBECJckzpGg4E6k7uNjTiUNiCHm
iTqgh9HfyuKPWuTA/tTMaT5HffG3RsEYOnGIIh+Woc5JQYiZxWHpBmJrlJN5
kvOIQJU8Is+0/6bUaifhOulxysUcT6GP3b+ZwoJAIBtK3T1XQegbRvA2yNPr
SDon6nyFmBtaHuomlRd1ARxJa0LGwH66tcfeAkiiEh6HzziHLANVfO0RA7u3
LXqgM2c2FzzkB0ozaI+Hfsc8r9ydsIrSGYDzTTnUNRDHrUyaaHd48vpdHU7D
q52KQFvuKXogx704C2GjvpixQS9cGBseV/EPGNlnE7rECFzVk2imVDAbG8W1
jBVe/3ybEAucdRosUNJac1dbPIf5rrxbsUqfwP2TO6C/VAF9v/XfY4t6FwQ8
a4/X2RRo38IP8GoNPSsgnF87Jadf3HGSR1z3ZvuFxDVt8ecO5QTzI+eQTntE
MKUhP7RLe9x3xHVvKODhZAZreQ/dh/ELb4PqJqeyNuUYNGaFMohE66VfHoJp
/WALt6xOA5KGVDjbSU9EpLHB6AaFU056H0FVVtjvcF+Oco7trXkUg/FUtLoR
C5wdJHtod6G/d9dF0UQ/p7IlTReXyc7wLo+5bG9SQarx03cxz1mM4EJnhjjc
szq1oEkMQ1EcUkPATvmUU7jRr9imfJKph/paNsfdO2ef5op7PRG9yk2ppG+4
ABOQaVhs8qLLAtsv2Ss8C8PkudSlP8A81KLXPZPhzM6LvrCj40Djs3sHYiB6
aiUhkFdJQeevco0c2te+G7vPeA+VSwgd6dnhwx1iKod5gyyBh3KSwXGo71Um
ZF3xsNkBT2GD7awTXBX2KknG8TsqwV2mUnWCFXnfTKWQmHYrjoeU6sR/lBVZ
PJ8CqkAwL8ZUJRihW7Cs3mBiZvqjhnBjP5QsDyPikLrHuH6C/pKQwwYkIyIF
cRZj1+urohChraftYdikJxAiYa83lx8LMvum+MukXIH9cW+Kw1d231ETHv7k
qygNkNSWVi6ukd8hKqy7MMiZi2S4nDiTXL8iOY0YNrgdjNAXY8LZz33uLuPc
/5L1NtmbR1lmqqFEw5GAWmzCwHcsdrEzC052X5M5vtXcjQtlheiqEHR/v2M7
YuLqc2+tXllhD/HLPu7uk7ierCNu4nrqdYdpYI5yKZ1a37zhVJ5MDlXTplDK
+Ervyy6S7RjJTBEFbp6PqzUnkkWKFJvIcJASC3sbpqOspOjYyMNDwNkcJYqH
3iQdzokNF2K5VYX8hecmvOJ5T8Q2VtlZfK0hYb1ByDtr6D0JdNIP37s4UpT7
QgAHTATUrlpxUvZSB17S6nRGgeplwwMQ8+kH2/xC+R64vGDghJyoVqBrqg2E
vwKPygkYBoG1qIRQJYAAq7c6r76m6iYS5gw30Kw9QI4/GVfmH5TDi2Dmss3q
87M2T+3dwTbGk2FPF4X5IgzF9bkgb7zGg3FTP3ZVC1LZwXUA7RU29YPsVC/7
sTIWiHdcsOYdKVDBNdezcBOMz1ZPbnov0caBNrHDfGNj9PBk3NmP826S1JxH
2G0B73Vv1DdqrBvHZbENLYduzXnMwdwh+Y3F5Tzq0ia4tMoZbWX5qBQRjF2F
W+DNJqWomKfg1gFH8CU3k7h6COgNTZPmPO0tIffjb57aNRhjES21OcbjYbQp
Rvj7z7zkLRZYns3n1q05Q7ZgqKL/Flaohea/EpC6DVnlaKSXPFRrLffRqpNr
YLnCcam3ZChGANEGcrec9ER9fdbzflhMMgs07M+0YnFm8Ig7x7he954PDITp
Br5jXRNly1wCF/RlqiAQtBdu4V/5AObEtQvddUcm5jLxBijcpoNacUXBa3yJ
RgrF4nAhBNjj1NpH/+cTALAergX02meknBGGnLTmekz0YXvFgerVMya+ruhv
kAzojcKIWw2LIuN668t7+2ZLE39DKwceRn9OGOo0ysW+WRtdK9mckau56SOO
Ko/eEWtgRpCUI+xRJXr3lZ1ndz61GbncGhOfSfk1uRPKLtIgvi7d7xm8J5c6
FkN2XIDOyCpzj9rCCK3PVKAQH480qRozotfpSJYml52QKUFmIMLh+HKmn9lV
YtnRUFm5BR7IfdZnlQ0uTrOF+f+Fu8iAORSwFfsuFLqKVwh6cU4w3QftZyaI
Ty0B8Hygo2VoCpzQDLLd1DRulQFsgAtyuWXxt4tamskBFIMvP8Wb//XrFpC+
0b5HTBZcCFcH2EVgkzzn6N1dTujQD9vhpt81NKsrjOSKCZoXsKyovtZ6q3cz
uFw2FNhYHIt/BuaYgYowvJjIQfTLv0z2/clxsBrRb92BZFrnSKR7c4y7HPP7
DP8arjD4REVEdKItQFj26XPBo5PWPmRwQpxYVPA4uTwyhXUG4Z/ba46LgRbc
edhUX5Rj6UkaI8/B485q5cd5jEhiIPEzPl+qK8txvkdQtEbSjeKo9iriu0Nf
oJzBB8EW8/AZWidnegdIlDxBYyt6XQC2fdl7bojj7MqtmaB/g+PM8iLzABj7
2YkDdOUPShM/S7YnK4R4cr8Q4RVL7oDc4yMjsZgWHVsut9EpCpCu63OK3F6h
/PQou0sPze5Y6+8PyQoF210yiAIgVh7feQrkjDoswRmhtiiVeRBE44VLV2D2
d5lhFnXqbNYBeaEy7BxwyrWNg4CcSClWSWgXHd3iiVg3AHyeWIx8Rg6MOq2V
iiHFON7U89twANXwtRwDJxez0uotcImI5ynXr2iI/wYGtcHv98QgDkUHwDkL
Cj6i0EAnPD7L5FzmNlOv96oZJbcpvnTwL/1VzPa2xW+7TjV01mNorkXzBS8D
VVsma3xZytgaYbyAKzc6XCKstlcc5kQEK+9++HKz3iUCHm0kY5WmuNuuoSZS
ZleFUEwqikVdoC3doLnAmUj4A3G2dLnnZHMqc4umAs7i5+A3PdFVHieX/etU
wx5UmPtLDZ4OyP8D9kNVi4tbtVP68fj27OmWqCwGqHLnCq/ca1KM9PSUiwU7
Fcm6b6OKeEvXW1kTjlqzbnwd+Q2r9YBJtjNthsQfK/xrwGC/XS51ObGlat85
uJ9E03U/HRWGTInj4DMSZVtY3ziiyxUC70f020NdALOfxUoRLb0uK+r8DLP/
UhlDlqxut9G5r9Jxu6TfMle4yWZ/2Bf/WGtbiZTs3M6i4UFGolFxzXcHfNln
x+1ZeRgcNyuS9XyK2zY1kGgQuuEgoPAMoSzlEQC7qLE9U6NS5HqWekvAR5CN
AegQrfhAINVnxTY+Z9k2QNpSMBK66hMRYa2T00YJrp2+8ESlEg14BeDrN1mb
R9qJd3Iu1c6RTxVwH5GUZtjUYZNe7Q4s+a/umb/wUjI3qUQyX3lyWEIHf/Z2
AXFIqOzzywWqyPi5Zod6gMwKBi3cWxpCylBMXOmc8VCGw5us3bo1Ebdc3zSi
c9Wf6E4lmECMASttUfGn3ciCtP2eEe6mT4GDOTltV9npb5B8BgEKRdDbUnMi
42nPuK1x8s/BDXlBVrNnTVOr5rraumm2Smwl8+Djc7AC9NntnLqjFcKAXxSd
oBBfMCUnOO3uhajc4CRa1a5jWWDMfhMOBmAKx9TsiO+CidxBB+16wKLtO2Bk
TE5EvNUVGQWVmVs6GL3kV0g6D/9+ENnvuvdIXCn5N1abOQgkj33VPOiOJNlF
AIYXzEgYe/XC0Ce2sFwr+daF/lkgx1qdd0CjTN8G4BrLVepsyrEe03VwNdab
Jwja08wtjWWxDYbdMnXQWV25J28tmePeUjduoDyz8O7p8quu5qAc0qxFD4Rb
/VcEcD0UdrlEBDnDA/KLvVZ0peOoGDhkuH9t5sa46qv0knJu5+RHudVq6Ny5
ak+xDhljOiE/H7fpX2hV/T0/Ebz4nPkdWDEvYSRGl4Ih82dR3p6kG0r51jUx
Wyh/KBiI20T7ZphYvR1PKiMfYAzZyVvkaX1ghWeiH3mB4ez4Gp/RoAaEG6NS
SPLEffwMCgyMOioKpyVTBP0Ab3d1DmgCbO5X806iweppyqOymo1P4JDuOsQX
XMibreg7qgSaWZ3ZxAKZTVeUcciLrnxAX/0oTR8Qv6w3TAfE6cz1xVZ6YGqw
ZG6Z5xeZrlv2UZXI+M2h/1CIo+qSDKsGRVwI/v0nba6pEJ0+Fh4x+snPKQfG
c8NiGnfJLACxYX5R5BLBwa4LBqQhECs7jBZChEQ5OQXxpSE5GejsCXQQWs7H
pibHBynpvMEz7m1ONFyjQ29H4mI2P3OUCFoheR/Kpq3UdOI8UM6BqA8RCtQ1
f5SvrftRESx9n3Blj4pNb4oLjz6mZ6PxuLMq2CEzLFtZHaxPgEweTsSfDuHo
YTTYf0axUtrSerBWDs3QfhtrgbMy4tXznwACwQO6rRxjYj2eGbX2LYjPcrPl
AIs+8CxD5suHgfr5eTsna20AxxBdjg5GlX6wAzztf4ygpkaKXygYSn5YHjlL
6qzb8XMDir13p5/CPNqsTEGVesQXYOyRjKUHrg9nNszduetU9peWNTW/Lw6N
hq8kfHVsoDJIvGmWJyMJsL0DDt+O3RzGrtNqjm6wYcG+9lNcqYA8KsPf0VqB
EMpgJ0QWP8Fjm2geJAOtssw9nuqufAqBUKl7w63dcjozLtjdL0Ph83aBC53/
iK+24EHbeHaI5OA87QQngi768jwU1QQeiuzmLyKVbMf8k2uXbGGwADD2odsV
9L2/Y2gbICOtlKDD1E8cV+qbBaL2w3h46k9SF/aA02NVSO/4h3EHYXqmH/RC
oMIaIyFEO6XfbU7k9I/p7zwU3rNWJLfHg1hUsYFRzUMgOotZib+bphjDBo+6
xTopjYGcYg+nMH5faD9+ANtF7sqU5Az8G28fHMEAkrJygZ7zJPs5iqk1aSnh
JoAPJ/ENT7VRscVX7djAXVs+0qyjtKVmXV2GsxOlT8Qf0Zjyo4pM1Qb54WHa
SN2wdIq/kLZZleCJsymyh/TIGS3TjrF4DoTdVqMI15c+MR5rdzrqBj8wSXrx
11Uys3HX3aLMcDn88rj6j4rLPxIWgvTzt4vsdgXPK0UIFKVoosKE/slZVCfU
nxCYyv3pRh1MsotP5V3Ix0A/LH8/afnOt8NVjzt5k2ZuAGYuJFSW4HS02ip5
vcsuC8TgOVQUH3zvtkYuOmPnSItrHFf1qyOr3hFqcH2hszBnlQY+jz+Mtjls
Y541ElTADe/T6v0GylxYoVDya6ErZ5q2Fmtr9/les51T1c4SfgduceMv91NM
JJKGoJKKpx7wpWk7S/rEqB9WdjtZNXv8VJeGIUy55vZNan9UZvyiAQEXjpWa
qBSXYxsjW+5iTUNPAvqfDCn/+cD8inLjDccpeu4fN2xVMS5uo+RAPs3lVEYz
7n364XyXDHOpKeejCCqCb1ZPHVCJgwRY9Tl/0EgAt1/51RjJu88XwhFC9eFL
rR9XagiF5gUT+GlaAyXWeI9WVccomELxyWsC2Rs5mb2My48bWy71ZIuBYToM
2kVZ56PTwKft07mDJtnvAlwoMPRQ8/hJfVJ6ccs3lr3a1jMTdFe9OafNVM26
ztc4VrzFqcHL1jacrhDF3I0YXKPd2xjqWN22xAK2K4ZeoRwDgA2dMTsQGNX3
geagpGG33koWb9gwNldN+bjAYb8qZG/AuTdcj2/WQTsg+TnGXjoZau6NZCpf
kBietCAXVEEZT70lCgZPnJDFYBvd9kYs757oRRUseS2lrZFD7oqRIo5GUCKC
sCb6fjcsoRTTcOWsJavTR/zWyn3/+gy9eRP5AUpgVPxTaNQCncT+v5ZN5doS
wkerzSB12qZvBYh+MkK4Arm/Pbmqa/M7Mw/jORdhhPCMdvpmMFdgkX9VEi31
DSbZfo4VVbRXJ8OtDHi9x7NJlljA8eFDkOiBWvbHk2/BVDkompxMgVr322c1
5vJDWRkfVxDw+35+BL8Bd2bllx25OoaTAQWQS4eIqng54xo0BniU1Xy8v5Ft
YC2o9poUB3JoKCfjjCe2rMr4nNHQv9wXqfxAdAOq+mt3PkKVxtF0fp4KyXoK
S+RLv0ArhVsr2gpp3ftywhlHoOf8mY7CzawE0nz5RO/8R2jKKnTcHJTztbIO
kidkyPfttm0UJH1rWv6Et0u5luAIXC1afowvFLLfUyw/o4a/LSRx0xbwra/U
eEccvW8W9aRQKDKbcJycSf3iK6o40fuXnkSeTt4afpPBw9oeXdIbcdEgVAN+
3Wx9LsXCAhgRXo2+vSDwLQhlcjsZBZrZVk+629sZ+esJ2pnbrkKTgULCHzhn
p2mZ7r/h5a0shPqbFmWM9AeeQhhyQXwygTSnzqpID7tSUwGxUYFWAZvw6Ykg
0Rqrgy6aTB6sfkR808mCEbEk/2wGQrvJq5AzC6RK92tLKuhLqbKLERi5lnZq
hfs1iZcYxp0/BLTSlYNtwmPcalDwBU8bg7QZZt2xw+HgESSVQq37XYtIGXXg
k/GY7T8kmi1oWAbQyPuMjZRtU9BlgJTHUi/YFVXnDHySEylTnCVjtrXHubBx
1jGHjrq22QyDlfdk3JzQpxoNzuGENQ+/gEof3/ijyt3/JWLdcIOqLYVfqFbA
AHOKGCzgtHajAuMBmZCPwAG83wP2m3dV2nyB7bX9M0iSwQGSwN75BN1VtCnD
fy44fRLWDER2C46eOuTNgI/5NuPvKw1GRrLG9KBHPqDKhvUbNuHRMXRZzB4f
sfloYKN8pbnRvzamBU+VC9vkDDSkwSQ0PldPH7A9gNopKpTQzkL5B9iumB2S
nh6RkhL2CP1zRMFlNc282+7cvjRU5F78fBzYUAbWe6K0QCYH5QyE2euMW0z/
t5++Nne0dFjdlNSqZ9CfHxSvlhepSKakt7uXTOn3PCkzcatCcpefSpKAEJmj
z2PXxGhOgAdbJDyhkfgqPmI3EZYQiiaduAUXn9w51fuo5Ttq436b9SDGUUxA
na/dxlRSijy5nhlL23KPWVYV4Is8Ea5SWrS0FQqWMZHfic/kRsPFXgraJY+9
andek/aT//Y0OG60zIe8n19ALmclQODa8qpynRpc7R5c5eRKJolg+qbkYTnH
5qzlee6QMLIKHWRfxrWZijKvA8Xc/gdUsvxdtkahPtnfJn/7wQhtYhcza10Y
7DUP+/QaIjulVtTELk3hY1twvWMuDUncP2TQ3EaDbDNwL+npWv6F9Ory3AKG
96mKo9xAUAyR7dWtjhdgN4wNyjNUKyDjStmuAdj0ZJHdd65j2r1/xmuCJxaB
eBq/X+w3NkeeNTHdX8/CWFRjO+oymFCFE4PnRr82PmvC1yCblcmh41eh+sEA
AkS6/IB+OGDaRrBbh0FnEQdJ3PHx72LRfMou88btnjtRKbALcchHeAADFLd4
ovxZ+L34jwjdNYJydA93YP55nyE2ucwMk9KeI04oJI+13gEUzz4KMqiQ0KNA
XmHtfWLxERJw/wLEp18sowNvA9SWzrMWbYy5WL0I0drI+hfmXRymlWivXwKg
0XXSqVF3BadziIcnxSDzFGquggt8gqoWEzWdLAYuvj/FYMtmW1DwYtZnFlYx
676zFdmSsv5UfrJIGeaGHpCnbXEUhGxVrPKIETgakXbfkKtsSsCBxAPAv1wo
lH9JiTZL6gW2qJTt6YG1o4wTlfzfOEY1tW5S+USbrrzexTUPY1LYUOHCr1jK
ioe+6uJhL4vbHD3SXg2f9LpXwBJMtjyRG0HcuggZ2NKsRgFj312Mq96CBM1q
uu6Wg1fZfc1z3IYX2Gdnod+/E1urtkXwy9CUKt7PDK2PSdnmjX4/OSGWKxth
sVFUYjxPUXzaKt2AF8lEsNVB+/w+asSYibynuBQNG7QzTtXhSCRa4YEHREw+
hvSkWwXpEEUkGnfNQqOiEnVB5GpOXM4E9C75vzJs+e/q8lpTXIullTFOVYLD
fDT3Tsw58yli1B32thVIalTryVqjyMaAQYSMRjFvYEeOUKkPPJ4Q+vskYnUQ
y9c87REbPS09ezUS9Vgn4anAe1VwXmkNe2l/t3TB8bCqgrc2iNv4XIrJxpoy
YP1RPV8/PaozK+lGVIrnARD1BstAFB0bIMTdwCGR99dmekjNhQOp1Zr8nRFr
nBTyTb3xgA/i1NIHfsBq1SBNrYCUuSgN2d+4GhcJtjcpzjruuhxvYjuDqFyg
5FnNOcMwEasG6IbJm1jKv/eXq4j0pVkcKvGpy8CM7xLe5eUrSKxh7SPxClr/
6mqCd5lizAirVSiT1upWJpys0c0Nd5bfZWdnxBHqE9cZ9ASr5XdHN+FKDrPc
3IjiInx3OIHykKclydyXPDgC4wYc1ux32iqAnfAwm6pOC3ACCV9gwrJuYXWK
RzWeTU+7HAN+Toi2slXSEN2jqoy0JBppbOQuobZ91SpnRtaIAM+bSuiVc692
CpreUU2UOxspikBUGv7sxWC0pIi6dDvmjN5P4yB5NfP62JN7XZzcqU+i3egR
QsEpK7uO0/kzOyTpRf5HLy8XCfH0yxob6+Y9D5xn3uPOZfuK4k8gP9AOVWCU
nqY3plP3dxj+MaUImyHZcgXBHepUoBr6xojhxtcsg5k4e+/Y7la7FsqJckkL
gsSyHPcImteFILFkzYwKxeFDRQohtY6754cKJ3o92RGzmfBBuc0BjJCLQ/Zv
L64mYzqLEmst7rsbzO81+aF181/9jfb4mZhNFUEjYatnbaCO1045S/ZdPfxr
MAdKGMdfLeBuxP937DzDP7e5Ew0n/B8xpbySaX69qYIG1wA0qqd3iUzxRxTl
1dUKWNBValK6jneI4uA1OkECELKhgrhkOV8J8y0Zljf9cZ6DqdVar7unTSW4
cvEoIfC5AMZ3k2Ioii6Ye0gwWz74toLF1Q+wGXPRKH/z8dw0B0xFDF7v1dSp
mSQ2uWm99F1c5xUpdgImL5pDKvuTkuuJiSMbWqTa09OsonbsPmT1hQ8ZyS3n
6vrMCedOVODSlmNm8Ccf+e6fjKJfi5gx+ScEXzC+m3bXz1oxXHgdk+DVAFz+
ZHJK9dCc3NIyjJLHJWW0BbHuSCB4aBf2GQFO2BdbqqIVMY8vE398All1hGdA
//Y3jATNNaXikDRl1XELSj51YrX6ob0TOjXiuAINOztUmmXzbYvRj1WN9Ij0
IMCw70SQXdZGZmcd8Ii7ilgYjpiiFuajOhl7meqo1qHJSLw4bUXyMDNFToA8
S6hxqzfzheOvt+d+xwqSsnP7KLJskOBPFsOYcBdXFU+wYPFtcbOaeqrMePbU
BTcnEZxJlm/Slqj24EHtI2a4fEHEPnt2mKXHvmdnSv1gAa9fxDSBwwoq7FH0
QKzkEFALz6Ds5LQS9MT2ekdEvhhrlBZliam13SMKjDy87abS+qg7YDNsdNW3
0KEFMvX3iGbfDY80PQytPC5ACqBJGeAjeNwcWeFBuxQaPPhOAVhWjPMFFBMU
GRA1aCQiO7O0EljZSCNklGrApZ73HRi0XoVc/Tb+8mfEghF6ATSJiTQDGQ4E
I+nwgw5Bmls50E5GGDTlhijVdJe6lrL4f6BdSwfKZw6jARs9L6tYoNCXFd/Z
ldU5yGNAUtAhNacpfm7gxDcqzlTgry1T72Dm6XIm4I1mbawFKAyDIW6sEr3M
xGjjoYRq8X7MWgxLwWU/LPj8jDwm4bvt9XT6Z6M+nWS+kbGVaYDU5A9OpFq0
rO2H76EJhg/vYJhFR1XpCHVj3Mo1/TgkS9KsWzg0pBy6fDt1YBBpErYaiYE0
BJDkKIqcLdLbj7LDg1/fMu9jMTqkemqG0Nzn1zpjSFpE6C3uToXbjERovHEy
LkhtJzLbVyhMvyWF+pS/8J9MXDbgq+nG8Xf+Vifu7PqVHqVF44ijLUPrTEF7
M81SJ6c7EiYWYtafa5SbZ1gFQvyEDIxa4uwO4lAIMrX5f1fyPY60SJtBCnLt
qBfTkFqludhWeas/dUGsNdVkSyv8Xci8l5eQSTa44fCQL8rLJlwngMjDc+tn
SQM5Opxbk+TW1Sz9ONAXXoiMKRBYm6uAg5JeA8kq6OVs74VkBXrtfg2UOvM4
TWS7QdcoB0EFTwmbfzJqMGisVY3WPcFCVn6ZoDdhJKDDhWYx+aur9HAd/cw1
f0HCLuE3zYSvC+cPKEMOs+2UxOuPIg2i6k4LStlW5pJOYkPoRgvizlreh/j2
ZfceXXWJCFfsazNmvJ28bao5cNW8SlbdWZEPL/1+S1Kgv/sxryNfF90Hh3aL
ndBRrQ+rLsZngPfLOMzuuynjYwDIkYGhr7oYn+/uq1dE3suAM3i62Oc8qMyl
FqyxgDV2MoTc1Cncrx0aRrXUAIlsfelBJ3+yz6uBdjVAnmFpqdk2P52LjoDz
tH+HKJGjwLky6HBKjKsdwQw6ttutDoXCqmJLNGAZBDGRZ5zW6gJSWgInAQZs
VJrkrUBqZCbzcL+iZ6AOBW2XBhaMMhamV0LKGEM1taPbEI9Qh0Ww6e14jCm4
GZb0xsbpgf5oC8xw3BHAQn38FqKa+jRZgjGU10w3K2NI6yq79G4eQuwtWNQK
Pms6KUQWU/PORKoKSfO8r1fLBIvl05lwCknNqYS2oIguaNavP/6pyekasCy8
d7zscK7puGAwPYb1/Q/Z8h7U1jfuIWIWOx9gha22GDzLL1eA0U5fItRYrdBg
3Xxz4cjhZlwZw0Djth4qHYRpvzD9hlxfryPtJYZGTXPpXkuxbKZvHDLMPduc
sI7NrOU5Mmaa1ih0Iv4vBWT9ml2q4J1LKSGRxrXlB4pPJ+Cd7pHMq7zpUnPc
nwcAExSRtV8QGsQ/t2sd4N1gsvnytCsxTpP9fQ3BGaDyvmelmirkhSkzQEDH
bRoxHvcdg2VcFOzEwJMc4BWx9OwB30ta65tbny2FT64LM70Kz5fZNyvipkCX
2QBY0Twil0XjaZRVQ7hrhLaIpLYiucpxL+r2nrUVm5yujZOJoBrsKbhJSwr1
HbSgTr/U4pcf5CE+LUrV1ihwoK0z2AOGkLppPZszt34drV6pi92cirSy5PrA
iI5krF+q+HRjSTDrR/UFW3Y/HJ9Szvbk8IkZDqFopLuLEJcJuS48iB//8Cdm
BgYvfCCVzkoqRCQBFYK4zioW7ZS5dmr1p099qg5RbxbUEP7HYbMn6hpmqOfd
Y1bk6YPyMFSgaui6HcdMyz3+S2ttSaNW8SDaaOq9SMdtJmAzHERmKGEp9B2T
ioxqnePJmhDORMKfXV65b0qtZQuJXcrm1bqZL2lKf84yZgsxZKKVkaChoxMq
WPLK/ckLZPiLzowyggmlWjHSVy+WqhZ5u7AfPTYMfX8uWuI/uxXyobp0DnXx
bBuNDZVwO5WwZ4O/Xu3fWpQ83cULNoXL3d302EsYdJMwjJwcSfRW/6Pd1GJm
s8o5Ctl/RvsyHreKSCsxYWhfCe+zmxr2zNQnJdDrJ1gTWn3lvHrdwFZaxTHH
LipQd8TjAXZDnHgTSWQykVptaGyDefGxnyBbgys2QW0Qwt2wKZoQaN/eDh4D
mDTjVsc9VTfei+XLMHCmLygsbuvJ6J7WVkzKwrs+4ZNJeQqtuAIpRMg5lRST
w9Rv/cVH2oh5DStCuj63Ycb2HSzG4uoIYyWLdWnpMwR6+QgpQzEW9ywv4CA3
g/kpeHEsB5TcQwcEtJvRW3gic8PRtFTjn5IWtbzt2XlDD3ycSHNawEBBy/J9
HfjVaroxyXlcuN38Pi0GyP+fHVfc3IcECwKWQEhsVJvhnFgsudzLnaRkBjFy
7zkc2RS0rKE8Vqr586srcnsYDBVU86n9RJtkuun0nbTcSwS8zspUYhnT45SL
xpLyyKHtTGnJcByfqU08taHeXjozYCngOgL21OJPwvY0BZR7UurO7qyX+dR4
I6zZfY4tguNIIi1PBPfyxfURgk37pZ1xRbor14K/9BnpdCQ+uCHar/1mUYOT
HeQ8VhyMWi4lTzjC3vabgJpKTGngURzJSTQOjABpr/cyYQTndQK6BDGdGGIk
FHVgc+Y7+6psoEkrK7/94yPVj+O/1gbm1+JNoTiO7DZwnxKkShLr4vb1OXT+
mZBymFSJmPNq7UvyA9/DbCT5v9v16tVZM+7tDvedeXnWEezuPODoNjD/yhap
FsYTxzxxMxpQzR16bLsIv1zDeUrVpVdREABPYEdNknH9w3rYjaS+UAceAnbU
xTCMldfqEnE+bX18FKB8QpxDRxTKh0ymbQLxVD7kmG7IoEDpfbtJN5M+wNsR
cum9ZH1UFbIEKtN2XfLQoRiTEfNLs/dsZWB45cmbGcoVfjcB0khNjMZmQU8W
9o0Yyh6jP9mcZLnK69mDN/iQQ+Fkg4AJIOAa5Orhk/xR3MSBOGGMWijU4gc7
OM3DJF51u5U9I854o7bJ0fG9PAn3P5zX4m34Yl967Uz7zyOoljvoT2vQT4SO
tPvllh76t3XUfG8Pp+i6Oi3+C7fxVqS3U1iJSzCyjqIFv9hLY49o0WCpJXyf
/2WJbFK68CMCr3iqI4HbhOtD6E0d362UJTsbO+sI1aG+FlW4i7X0GVWsoBT3
z8EhpKR4nHknNHc0U8btBeaPStRm/xamR4uwjXzoHjuq9eERkWYoh9q8bAOd
4h9cjEZzeUaBLKlq1srghQWtHs9q5+B+1EEyYMLlN92E5SLcO//yrYe5c+Ry
yO9D7Sj7srBkzo/S8/LjLro5BF+4WlBOXjnbdjHJ7mDS1jofppdVSXmLMrUz
L1pCJK0kgFLpfeV5e2HArY3AqtMOggDbxpKEbMwD5+rt9y4Fh90SbkgZkd9m
mFtqzb9d9FZuMRcP0rhb21OYJ3h/belu26cQIe7CpIcLHvrOwl+QadNtGvJQ
dd0sHbTlwt566WVZAw8yYF+sDBfqsoFo6XXcz67rv/dneXp+CaZ5c60WLWrY
PMYdLdc08ab3b5SxrkEcIQK8kDtEQ+o1jhFgR83Xyq4uODvcxaHjR/SvuYkX
X/FV1IiNczijO0wbIqb2D/1AoW/CAIvD2cWkFjy4IP8CiDBsTjLh65+nTNug
leYJM9Tsx6OS+Xe+DkYzEw5hi/mHXwRr6a+qOWQU1/2EYU3lCXPvENVtGUiD
01ss96iMgBTKhzFysivJek/jzWjJI4VVJijmO9RTSBcUyqq6DMtEvaITJ9O5
yATI2watl7vQaAiPRtIHuE8HhCzHdG3z0wmaLhtwRxff1HiuFTFa0Wl8KmR9
uhuWW3HQZ/34VPyZyqh3U8KUrRgl3m/V4YtTYS9p2go+7pgJzdgQ+Gp5q/KD
tWH4OzQa24EE3eeP7p1oAmg/px+nNvz+BDfitpurL0kEN8FQUSIlhmQqgtK8
k42d63AS0qW/AMUmCyE5uIXUnUyk+D0FnU+XrOrIxaDDgqiHcO7q27fReDcK
mZ4/OkrpcKs91rz5qICecSxQEW/xDHusJNi6Yjv+nN4bnC+PN8lUn9gk/TIO
cRoNy4lVO/LktYp9wJfK1YMzIxNCuCR3FPBjzOc7/+EYnM+pLJjOpyDn/Eb6
1bm4KsVrZ4+u0gKKLe4EEu6Kx7EsFkKBY31En40WLOJRxsFhVHrP03Iu0wpY
A2iR4tpg5GisRbF5LrXC5668dkno50H/WXkDRKfah/e9aLE9rT8V3Ytz5aUN
ln55fFrjzegjvwKRVraGMnlB2iFBh+oe+iQc7PWUDEiseKZ8a010UwmL+WZt
GmvzPtci1TQ3i2UetPLQeZyOIRrL218/wJ5ib4xvsUxk5U1iZNX7VlTfyvy8
UoR2WNu+hZd60zmiComjWNfu2kgulzytSq1JxXD7Deew6eGpvZfB5QBKHwXw
q/x0aNHVqU+bjPf3Kdgmg5e5vKaO7qRYn2Q4/a2sngzk3pkTdjPq4Ya/w3np
fgpcgC9dy6lOtCGQDEfIMzJdmSlNybLHbZDP/O5RUtuUu9BB2lW0QJnk3qUA
83GzNISZ0/4hUuqIsitQXhKKhEZAGc8Qhm97SEJbgAYe+Lg+ABTfE1jlbWNs
7LeOLrlb/mpAqcSM+Jv86V8tZTHs7K9c7v2uCDTHhOQPoky3T6lMhpwn9nnu
rZLbr7QEcduWf5rIc3kcvEmtJf7N3i8ZCQf/JWStStAzOJCho5snIFMeDsGZ
ppSZEBEVQG1SoEHVP9emxzCpS6skp7kXLgm+wziJevp0HvNp+NNIo0cBC3z0
PBmkTsIwRRvOAebGKBhJz8ayXws0sxZ8FS9qMWUbO/UlYjWQHHuPBXy+3N3/
CFOsTE5zMuNb9v2CvYIm3mYQGKRbcRY89RCTLrpfBOLQwc4wH/ZeSp4LarPV
FxAlMT11AvDn15wzKgNHHspRJfaQQJ4YX1YCkjqkl65IXzo5fZ2/cEFrKwOI
GWRfbKftDJOdSn1faNQ3PHsFIDQPfEI75UqwMCS6/zxjTvMqsFHBAv9IiUa0
ADpZTfqnYNimz+/l2OTi30F9Gmm3c/D6SSZvFlM2iP92mvey2/KYQhvYrvxH
NZbc3RkyYuEPAMUiraGZpB9ewp9Us/6gYgIY51uy7t+6IKH8MpG0wKhMEgih
/uBsrX8wf9zOilCgbZx9SrknZYEFDJNfpsFXix1+awotwi7H8lWMJO5b1cOz
HOOTWZQ9c0h31/5XnmvDj09/PSjE5QSimFa8N/rASwDus66jm3DhNbnudm7u
3cgEU1E8qggGfvwcCEvbgwPCCPBS3Ezw5rgOKVc3wrH1rVBhDbra5u3tsSXF
A7Ye6iJULrO0/bItfmnOkW/0Sv2SYTiB7FTwAy4go6ORfCaGkJhWNX+C5Evf
j0d4VmBe3iFX5PrOl8V8WkqgUzFUR8CtvbBgEieuF2+L5gD0UWKFAC7U2n0s
xdVavoY+G+G53CT0jRZOcjKcOyClHONaGVWOQjwwTroQqMW3lGCz20bON9Zd
RdntQPZuRlL/jgYPK7gRl5J2/W0nlDdXyJzSqf+U/C63vnEHqHBukE/w2hzl
hjTESl3uH6JSQ/UlZ6dbnYBqc3nq5164/gMolnQzjMXOQ64ezbZMfsJSEMAs
TVYz6mc7oSAOe/aa0yI04IVj7C9MLjNLdLHUIRqxRXE6OysSPRfMnS0QKPal
VKrwbM8xCp5X4QbK52gy4cEuzGio/tV7zVTLzfaJIcTX1HmCAeyTpIef7UyJ
QWmN92F8gtEK8rJiZfOtaRKLc21PbAsFH9Sxlr+e4xbIkq77eV7fPVLXn8Tf
Ow/c63eaIJBftNf6OjPbrqR7Qvd722zz2+UTtQZZYTCJwaQxZZrbxs6Y6Oxj
FPMpIFip4XIOC7DOUwJwu0FJbL8Gdv+nGKnlZKsAut8XWjnEYVctfp9j3xG+
6ebKuOEOBQlL1uXY1x3+Dz0IkdPl6WZMzmBipsuSoazdwSQNTWUe9kCjKxvT
204IMwIWB63OJreIO9rVxOrV5+sqP7UHYR0b9A8RRYA2xhk/YglStX0exSR8
MWVTaD/UtDeGKmgFJl+z7AFHmnMEYvm+n7ugWTzDQMENQrcBHQlID80KyoRO
XaWpS2d7UbH/fJyUOZvGr34QsIqNM5hlHMKsqcOf84XDfJErSiQQGAydRuSl
kJceJLnK/bbSfpHW/lkTph2y0ZNXHQmoPtuFtDxpDqjxeZeNmw7JlKmkpe51
nM0/q/dPo2BK+AgKEVvDEVQ0R1Kx95CgWsQNtbt11pvrc8oyvkBILgWRlB2w
tZcg4TFlgOWZirjKqx/c0aEc99szl+q9OPp8cYAtPl3m/W3dvjDlND68AnCQ
WbT52gOMaUB0udL9zuQdUUPAqrwxRD5/S4cAB54w1iagBmUbrZCs9VyB74YM
5qxTnpP3x8SwrIYHLX45jZxCi1VVPm51edQFtFU0RxDI1SsRVbAw3uhvbCk0
NlZXO95fc6UsaO1lGVon3K67vfe9MqqZ9r1IIvscClcUPqoQnLiBObMEg8Og
qFG6d9YQ1TGRH9WDxNeVFF+1U99g6+C+7t78zkN8crsHVqyIJtImcAiA4H9U
EyxgCQzkNgIaQygJE1OJ0PuKuDShSwG7fjKxP9wGY+8moKTAnZq+iX7DVS0M
DoW+NJP+0C/9psGzH446dw77ga9e9cyHxFqo0j/GTq9DzC++I0FFyH0WwLEr
TmedM6WRu+ys/2eKXAIrFjxNNJYZk594W0TGXe4X4zfeLJXJwJW/vKTTyp55
dlApjCrwVn3HqRs0uuOJfkDYYpiPC3Vc/EuJ7uQTq3aeh9Yk4UDDa6wEHKLE
wcEt7xDb+zl7ZZ3bb1RlJvBxZomF2nIRY9UBLSrUVBheWFOV+QfO9rqgQ0Ys
FSlCZLu7ovmfc9iwCW2VN9qbZfFu2HjTuGw+L6FZkfbUUwZdJYjZsxRWDfKo
wc63WDpOWxoz50zQiDCDBfsWi7VcPGrkDbFj3SOdS3BFB7B7rq3tyxoU/pi6
0UIhjHKxUVPUFIwMQHY9SgVMAinyUJzOt81T/ma+tIBgcvS7VZhU5M8QAjuv
V+ZN5babwm/Fit5KFJmcupx1NOOMfELzwaPVbG2j8OBhmNB79HFNfDMJ9hmO
6RIEuCSyMiD6StjuQYKceKA9wBkJ9O4q20J956FetupGM7GuU+OgrxcYHpWe
lEPKR2QjkZ71/5VThm9nCsDu3qQUhICxfsE2NcjPx1nG6Re7bJx0Nqm5BF3p
ESI4kav7Udw37/0UK0R1L/w3mYlupNkJy1+yQ332opjmT1VGOyEr6Gb2Z7GF
TlRQqCMp6nzA90MFlyqVYFjQZ/K++MSQv6kuEyjearVeDyBzljkGh38qI4q4
pPf7TJOj5ATgRb3aPSREyM0lBo+/j6xSk+YR0E6NJln+deJiO36qNB+IR7Uv
4K2uYHGBdx6sUcpEc/rmB+wuDIIs7sHoB5gI/I2wraLeHQ0qf05sBub5dKpy
hhUv3Nr3yO3YYFFFlorarN3sXdHl11rP0B8pnOdZjeMX7q3r3J8lbz9EfrmX
+Jdrx1dTMQeNUkK6Clsm879niMiOtjZJTq99J43O+tLVZMbmqE0dCsU9BL13
UUwpiki1s2OktBCNxgGb2E9+LLGalxnTO9PLuDZrHjW+shfvnkUQ8/j4h9U4
qBhKHAZjnWyPNbZriABw1RLfyO4kW5Tlu3VbJP+cuTCqW5EenI9Qopy/Lf6X
cQK+Yy9jEp0EVpfkMRW2UYXf/tehf8q/eH+ldqrD0g9JcnG/OEBelf/r27JH
uBnAP3JXbdXLTeh9ZFum1aRMn3DRU/BEs+kycIxmx17nyJAuUNzkT3l7M0X4
StLpcTxWt/paYISC5K8hp9MN+D8qo/oxeF/aqEf9p+upoDjpBNLt2u+DxTJ6
6ZLYco4MqXZv/kvoyA6+mw9/WTXOUo35L8MCBux4cHu8foVdnXli3dbTD2Qy
Z5H1PL3wPSavr7uFWR/Ps1jEv9FmSNKnTpQ8+jLc++2JlQVbKXA8S/U04FnD
iEJUzu5f98s8ytF0PMlIdZmhi9oQlahoqD2ItMmkPb14XCgJHsg0Ld07iO2P
RcGpxq8qn8n/wvVTDI4shA3DG3Q84fgHCn48ACpADDTfeLYe4B6Q2AHLvQcr
6FU4ygPLL/2fgFfPHZ80R1mA1sPZ//Ud1JF1qQewR2Foj17O5YKuh2/GGX8q
UKDdbeLRUz/PaQVf/2bLAHTSiMfjyBk/Du9piujIXBMDTED/eQY8upoarxV6
0ghN9aDBR4t3v53HX1ZloyciKJhRnEvAnfkrzS7ux6Ic4GWOLJzvcF9n03Ma
X8Bp1W0HAZMCGOX21t6H9pYcCIcrZrFppJVhM1qyJfmm1pUEN4b4aWkZFYOk
nsDKBNJwxHqhcYNc1IoKqA6yKbO6QccAzPmoKArEdTllMg5cX37amQSpWrJE
MxN0+gFMrxKBgJJcVyWpxeH4i/dPqDz8Ie+q3sCOX41wyDm9j4zZ4A+R+V9z
Y1LS1mbxQYB0DYcFaZM+zVLbb4TsvoMHPCo606tMEdQ6q+PrC3Y9jafYLsyl
8+GVFBw0npKrgk3HkWbTH3YRHFYV+icJtcpt2dv+nC389DV8zU+wHhGhLiWR
0DluS8XrakPbNHDPKnJZxyEWS8YL4QZNyOzVhWrsCygTyMhOrpsH/6Ui8j87
1JAbs0zureDWtShZS4uGpY0ZHh54ZDTl9ZFe7CXXygxjFtshk/cMlQ76Kc4G
Q74lZ0UPEgHsZoL6qSs9Mzim6x0+9kduy9k6JGBd8y2yJrK2tSMd5mPxZtzH
1EaMPrPaimdwf6ZV8N9vUEO8cj04LgVn+xIQ2qWudRTST6IyXuHztO0xcY2a
vxBWzk6FC9P8dEh9gxHbDymlaJFFw4k333U2Uz3xTArWvGHmvAdVk47KC2TK
4V4x2gZpcdvhvvXHBlgSthla/yu7R1kGPIavULhAB/AmFMm6lCAVmRS4YZM6
mx7gkHrZq/dxBdfh0XtJ92I0Vp8NQ6J4tGL33nLGl34vPaw9VF27p8LFZ5Ke
ONg0W86T0A2zmBzCKDVm/uGvOmWK6jOZIbBdKTFGuAuF0zwqCglCoyX4thoh
YTRzz+N33oQbzya2lTYWOVap11KT/VXxR+/Z4S51n95lrCCD/k/kaibofz4s
KpNp37re5KiD4tXQRM9QoNY/sdkbtGn2mskYnZOFLPAtb6zWe/rBaLPB78eU
ItMnhWDju4d1yM679KbgPAnXkK9Y/+kADLX4+ekr/3Nn6rEc/IurEKZ5S5Lb
XrcH9EZ5lPzfqDyBVjc66Fgu+kEEkkYm2wpGVL1OfqT90zcE1xdabpt6f68D
ueoGtojhn5jzFv3CTVXbo+1A01XraeTHUQVZukiTTXLdeLAVK02f3DkDL6VL
OxZGohWP/vjeWPwXq06oBN5FR+kS/Bk91j+tXNnmwYCqNuQV3yijNY2sv5tA
x/y0mCJa0Pqy0sMMWrnSdx4KhOagwox+jfL3kRQpsTg6lFYVLvsJgw/9ZKr4
C2K4tVA2YWIF/311bzCiPydhI3LiXBRy5qNK93Na3UAnHU+VqxmmqmXzW4Lh
ljWnmanaVgxaNUTm6x+Nwra2VaUStDx1fcxa7MQNkO7OgXpqDSYwAK4If4Kv
MVy+UyXbEe4y9XAqw8Fw8/t8foX75TZVzGpuSduw8yL9y8mEd54cFB/28ING
a+JkDWEY+87fVbsGpciemADV3qluNRJafXWCt2in5qhu2re7fRRJdZbRE/sz
9zfYe9MOgcqbJ9w1c5Lva0BkWs8D5CrCsUlCRRdfAO/H7Z7c+WBspgzn4gJN
eSJg+prIgqzTNZ3pxIptF5dcTzCBneuSeNskwpSFedMk/FoWfluiTyTvjVUW
CYW3jpbieRucynyAD1g24lVkXikSwZmvfJ7K3JDhJ8fHnQUO5QedxsUm9P2u
0mpiaGWXt/9T79PSGZMAQRRevof970OAuDOKkWJarHtXFhLzI9cFaGp1fKRn
MhSlQnzNbcekaNpojkIubhNkfwihd3xTGxQg2x4fsJqPsB72Y3DZJlanOCD2
F8/9meACI9qEYEfEQQTWX6AZSNuaWpoeGGYCXBO4UksWqZ+eaaws11tvQYgs
sYXLaZnmjv40Kjijk8dGAlMooNhgMiigFwzUU+dPMPcBSaZqvdI6dzFTTkX4
JW13WgdDwOokCS0pEXVimALiv9aA+1LrNjFkEo247IDaraTdGdb7tloKdhx5
PV0TDUDbP9lz6TDttGHWBKi5631tZKbUZahpI5K6PoFYgqmDFnCt4cQlfWki
ojixAwDzMA9LXYX43xvRKAXZj+5BC04oSeC55R+/YOwZfCbHLg8XxqEWcVXW
m9YDDPqBGW9wx+KeOoPGOEtI7mS9Yd34gRSvm63KW+NU/4n68a7OQmSwhMBS
2I8S2eaDlDhWam12UrRr2X0k236zVTGzK20DnBJah/QEPw+Ciozut9a/qJJj
S7JH7P6qeM3V+chnwr5pJ1jXf3I/z+NfV5ygosvwUokqo3O/YmcwbU9ogscc
3zd+j0mkdcZkix4b1cX/WwZdZQ+pQW50NbN/v+YdhTAW+iKRjmiyunhqEGlc
qDZXCH7sZMAyqF+ZvsqWxtODuWYvwUr5c3A1EiEr0UNmrXdDPZTfhfBZX7W8
pWmUx3xhkctr/7GKQ6d/wOladSVWWkFlzP4U3yBcuz4h1p28uBW4rgCX3fDw
g5kAY5juofixIHKpxwdFUOp/OC2eY4DVvkzT7kJEhi8vU/c2AzpF/WuLoJPE
ol79xCye0eytUpjvyPwirzOqlTrIk4MQoNFDqNm7P5eVa/qkafmTMuMWOMPz
KM/mNePPfgWgd+ANBH8d07wmYnr2EZVzuy9WVnSaHunqgWZzjZlpiN/35ZPV
5IUg7jTKqe52UZt2ZVjakoN5jxJ6moQYGgCJMaS3nGY0zX7AX43mNRqrJ315
M3G6Jbc1qadLc6WlhK4sKkqNaGDeTE2gQ1GDiXBsaKyw6D9sMypev5Z4zfEN
r5UCLLrnpDkfDP7L9ZeSR8ZBt+ZsgbSUw9CXIn88tSMK+eOEgrF1PLR3nK8Y
RIXSvpNt7gIwf3vcdVBgEKZpf3MUQl88EGRYSw/NIDnjoE8xfZUqWPeGyD2v
2kHXD3g6MTga8/rXmOroF7qWYeudT7ljMjJOuUfvIlkciY83leKRIvl+pFqR
6IcTPEAchghDEIRv7Eq2AHceXMqVEQScUXzht+Bb/UJayGnNz1StQsM593Zj
CVi5tICTS+2I12UBk7gG8r6Y+Jzh7yGz/L6bmL7gdNLE4+eBmkStlEoX0jNI
fL5A2lf5z223Q7oUJbVXCmUicGpIGBpkAz6XjPSuJmOLEW+lhh068Iw75UhY
ZgdwuONjjjIep8py/nL/XjTaqUu55MYRu3EE65fkwCqFUJa+cCdMsADS2+Bj
37rAGTrbWZwpXTp/F+F5grYHIvS77mh4plcQBTcpovw6if0R73qURcV013GG
wHQT4hDYAIH4h2O5iixCljLOhgwAvYeG+pV7RER3xoRoJsfn+dIqDatsmoe/
WRNF0emhoS/MlFNd3S0o9S/Bhd6X2NNdpyEK+ifh/YM0C05Oktnx/lLqtf9l
j6GRD6w1iGTFh5TqdEx6OqPQu5L7+unYla9o5KjaewpeXS0LVCcS925LWmdE
xt+gXkIZVDZudRuFB/+wpPkN1sOxUd1D7XYat+bIprTTRBW9wA2Ttaisr4Ht
Ru93wsMTriRCVjZnbr/v7zXM/LhAZh/HxLgRpWt1dZqH51fs/HE4YjtJ5xqb
fNs9hIRh4aFIH+Gs+IA4uMwFw+srWLqhNjL+/Z6fjJAA/2CGdZ2FMkQDVZF8
cqb9e3e75WzOq7DIKh6O7ADPUUVxVR12vmtfr9YSAbnHK+2YTOKFK2kFOXnt
1wuJhjdHZgOeMHK6FDzWYZlMUWCma6r1uAs6v/Fml9kyxILeuNSgKRmZJQ2E
TnsKYwSS63NkdkSbY6Pub3380pJC1C8GHxMlUjHUViLv/te28Cq0QNFBbRMM
YcofUNNwndojePCOFRirsViMjLwpCETewMBwF4A+rEy+7rTZQ1oMUXAl6wsi
NKQwN6q+XkhDYSPcNhj9AI5AGyc9PbPOFNHFeGL4pJ1whvSC4dTqtyuozt86
A5T1CPgM2EalEkGomtRF0zJsY0rbjPW5+3h855v1JCo9pWjDgFpfs54NHFNi
kxaErFz3sAxAMJdE0bk/aECUsN2DS2JO7tcDQGTsdVN4KPeGi79qhW+nztGy
NnPZFhhtvqupVKbtmphAHp/Rpq1qBrMVRRfEGEvr5yLVf09+MaU5LGl4oI1J
Kv/XiOq+F6fm0Jh8vC8RxEAGiQTNeF/JSt8wqLfRND/v+HIjcMwPpU7YPkox
la0VKHcldK6ydSfmB9OIi6tnOmS60Ai+nf2vOz/mbra1DKjFyOIPEPta0ALg
7R120csx2y4jNXZOSO20vvNfwKbjeZKebDHY+x49dXvK2WjqY3+KuEZkMsrR
VmhSbvWvEnMicuxJuGciFnqCPOzDrEi5WRR0IaU2Lr26XvItvErx36sqS+TY
cCjDVOXJee69MhguLsfA05PAO/CerOakOPl5Mu/xNok9eharBhSeRkQ5BiXC
5Y/EN8AnKraW0NwzO+DAxlWf1ycbO9QTORG5ZjZpYYV11zhMktJuVubdZ7y/
YA9gAEJ2FC/y7T6N4LKN2rSFvC+AaZkRui2R9ur1jJASYY79b1xNIVYyPB8R
vhJQ0KATcSMVBSvPWZSPSdUSJZXN6VXPtqXFmd0Ci6r73GH2l9sNYjMq9oeb
UtbTyjG9sVUUtrt0y1xHb7SPBwwVCpu5p+yr2TUyThlEoTXYYJPKRMcnh+Gh
rfA6SY1TUIHdXFI81TIY1e2KXJfVU4Hf2PSCC8d2MTe4aKU/gSr81LyE8shV
o+JV4gHsyUZ3OTVW0c7EUu36u6itvt0fvz4NGkIFPuInxgk37JCdZyny6DgG
k99Ptoq1ibBplbhcOJzCeEJmgYlxFbibO5s8kX7SK5yDZ8ElNEnOhYownH7t
1n5nTZs7Qb8yJ+9qWUg+Fo2WzpJSFGlBfiKzbfdUQxhqon7eK9BpCITrq2Zl
w6bWhzUnaBOhhaIa1Ajx6SQsXu3odoyj0MNqHON/ymHotYCZaM5RhWWG3V58
FqxthZIatI2F5gMfgnc7oiGxRxWFy3wArDHiIClHFkQd7f8FwAHWaLCI4nrB
TDtafMK/3qi8mkar96/Y033sXpBZCwz4nrDr+yY2HDC3594Fj5h0ygBG7dw/
3d3zxIkL25QG2EyfYGAmUmupSWqo3UI0f0Vn9E4/IAc19tRLllEv3jv58/Dv
yq1QlllErJ6m5M5YK1HFmO/jGdWQ84LCpBLDEb/7auiuf/nuczOQrJMGcp1p
LBJOMEqFr0U7VOK0HipN4sC6fdo1ZpUXt5t62liMuHA7jB0ExgYDfP8ZAREr
ugrjSTgWC7lfzrEv6rB2vT3iRDMR6MzMQbJNJCl7LVwS0sxHKaNaw/nshKrS
fvnNZHPkJvmbcTAimt4svioOqn3sepjh+rkkCfuNsZRRYSynKx4mQmaYafyO
rOdWAIkjUgWanSvycWp48W5ktMk/A2OG5cqIYp1Lvgv2mvdIuu1oI++qdf0v
uyJvIBgC1VGZ+mhkNfjjetBvzUSx11vziJE2hEuHOJukoJeqP4YigXks2oBl
BiAAiiGL1lFObtKbRHL5GgLT8iFu9inKE6LDWUrVT/bjEjghAnvOdsyij5g4
Dd+nOfFCOAqtPk5+L7DKJc5VHff+t0WmI+uQY9HzOtxR8YNeaQhhnxvwvRea
+hA9eTMxoikQ23er1QPgAb5f9pI+OPgCuJpbH4BDKrKGSXuMaQqAdjr0rASf
z91NEPsD42lEAuCZufugWBPGEAAiVzjEcFiXuWf8cbW6HG9UIkBN1RtmoqOs
qg2RluDMFu7B+vk9cWOK7cafE0PH/agDKnrnGXFsLVHaJ+zxT3cnC41/ei3Q
BaZxSIpYtPXwY52tDuScH/XTbzZ/RIjC7dzIkKz5dDvK9m/Y4vfDfDJac/5R
kRWt4JLPu5tNwCKo4tuGZCJR8amng49kq3pKtxiMd0G+FGsHmdXMSykDv1dh
GDleHXX2fXYgGRkKeiX7PmLOUCc2CJrOa6BReULPI2+rLUQwHyIvneglwyym
lCeBdOd8LCjcLRFzvDyJtmjq0TYpP3SYl2ASalxjQg896olgMgspz6nK9zUG
tQCytrDR8VVqWeR5h+crNbok4n7Okd+y2m/WRFmIOrKkfXdRV1CRA/2G85ub
lvbkOzSAr9SfC0b13VySdPegOQfajRqp2TETyaVH9PwWg+9BDpAt/mIDi1S9
rPd4xQWuPQbPxKme/q7RiXedGEmTujna4QaDe5HgQ2dU25SbtTGpFZYDwq6o
EzSqsP3zZjFvhBNMYkCawTFmBmbdT1CB8ZGKVSb7fd9yqqNtgBN9tViJJoQG
pG966gizdtzSDbQRlkkW+mfdsSqG8P4AY1grFYJfKSegaGONSMOIcQI/kq4V
bQiu2MpFYVMFU/bqVPHU+CQpnsOIbaB/P9f2G6tUDs4urquh/RSM6oexR0IJ
eK1ZwerzWDEBXQpClyzn9+4J6SvE0tU9MrD5RvOxIe1EZguNQH+hLN7/OUMq
taIGadB6EtpJc9AyZl5m4IfsYU5v+BVKDO34UFi9R9sULLgRLSCUi44cz+lm
tjUM144WgMTtQWF1WQXBWngukrP4Gzp8VWMbz/APfS26DkfwPuo5/ixcD/A0
yjOIh9HCRfH6Vf4yKq/LVT2ChFjhPDsZjqB0iA48k8lMwYYS58Mlh7PcIza/
U+kk3fRowa3+Qq8WUcelKYJzpiId00UPqd8ygTBlG+y2uQDMq6P8y6kjVJSn
89jCkmHvfAAks/mjI6dUDMfUmMIBueStJbcB+RHqlikns/+dhrPOo669eehd
cY+LP41POVvSwJ+2mJGybhBewBmFNOUnoU/0IBivDAXGCBrE4hoyDvH7l0wg
B+uvigDG8oiOZfqmlHih/6o1QDvOUwxUVbjYCz/nss6asDqgQClN2OPvz5hK
bKOR1ZXGHrtpmgvz/W9sWLMy1t6hRpqh1Sj2kUNFisutTDG/DJGOpdQ+TcT/
x21LdNhHh5BxZemr32ejMiTXmIUZbdYVe6IxmuM/1Vp/M/hVYV6cW3c1Vdk7
elmMiaQotDcaFBEjWNlzyGpW75hmCiA39cniGT+IpGYm/3RuVUnX6RArFII8
skj1n4AmpxcZXpYlz/i/ScO9Ztfxg7guKGJHgxSpsk5fFEBa2jYBKyHZXklC
q8BRxVZ1RNUg3tGJ83UZUbKBIbenCPDL0sOZ99kL9qAOl+lYW5qyQmvJUmMH
d+Z9P7HCXKDUIskjQcg1deOSSefh0Tri8jScU8V9Zm4CP8iEOevy42ITMyXV
IiG9UXV+d3iYQxFxgOX0hL2+t4Li25u0iyzVN0fc9PSugHBnbCjrsUWh0HKo
0aUAPfmWJQtXNNuxLABpBxQ4/We0nFZmHW4nA3TIAUZnczz+lKFe3t5xSJcS
Nq/YlJXMdkVrycsAY+lVwVpRcesdWbM9cTh6N6PCuFWu+djPk9HTQsGU/Ot9
0jxBor40FYs1ToKePYPoi5hBfhJA/GhaIBaWWtgWbraN5Bwl/8/UbvCY/Awn
AG6349nXWDmD1D5m/SHg8K9cE/CQnTv3AKN/koUmN4cshP3YhYLi12GhC+gB
bIcTGcYiDYBJXx9kxL4zGYKji4UbDFqh9UMsUdwha7Ygg9VZis45QFSnJtgD
tra14zoAbILDvmP0/Q2o5JiZ63ABPyaLhUnAlfGzuylPSAK2AGT7Gve3rW4W
xKd4q3cP+EswJiNsK6XWNVQQUwYOogbTBYt8B9Yeu+mnYhT3kp8z8Z4g53i/
6D64e8BtFfjf/uJ7MnBxwBtou5WOHaU4BXzGUpa3TrRIjE0rL8h2nVESMx9O
yPUGzeZM8886OPrkJcFbfKDwfY8zRsUuwSLTpwg126q9hkSzHx9vWEaM1dS9
nHDryriCS/PXPIyft8shmL1bCYGplKmNhugv0NQFfK1Eb2A7zlepwkbQ6giC
J06sf6ChVmpS3FHtC987Bi0Rz/jhyc9887sdHQOjqyBTUYeqeodUNldVSNS6
pbc/PpZ0Hv8IuBSx3B/93DrwqoUfLCAascnb6G5mbN0ksPfg0Kb7kCxfZtEn
6hybwqLMyzhF4/NCVVoqntHGZ19HZgTs5WX1M3SNdrAGdT9LjYd5c1PJ4x/T
dhognFZAafn21IcvM4Fjkw6MIpdIbfVPnA8EWUdZpxxnM9oUYADi03f+innW
NUEIgJ5ZMvyITwGYECFGdkOFkcd8a3VcjopemOvY86x1pqgn9efkMnfSwnZn
jvXgPR0bWLZNPEb/8DzgogGtofESwDW/G/BoZ/+I87BNuXRwMDVshnht0CB2
KuxUjw3XAusvc4BkBvq5Jo5qWWC99SG4ZUOpVrQJCkn9eNfqqUt7DQT7Kwuc
7GeUJ3a3M86UGaQAxLCK5cqJpJ709gUKajISLumDEi0Xr1J+PPg7tAhtqAIq
6jve9yTaL/qxKfJVB2JP46uTU+B+ZqhxGAIHWtv0xapkTOIifaAix40kSMxV
6mUAXPTECglSwtM8lUkqPW867vDM+zLirUumxoJ29vl+lNx/ETpQIAI2MbQH
J9F4IsU4XbuTUb26O0gxhJrmcAYvWYkhY0PThRbCJ5sAW7gfqLKv2KnunDYK
65V/t3cH6wdfzDnCBOvjfpVcXdNRKANcRCCMZH7c8Mlkf02h0ow9Snu0nNvQ
51GeEN58+HdR56hnEDBlQQqXH2EXzE+C8Yww8GH/IDuOooH8aXX7pVmwRQXe
vfCQsrrDs2hoOeqf7475Sk4Z/gWfHs4p7XY9p/UUxLaoE0OwVdus0sgNFrV4
8BNQK2Dzu3rSaifwp+m+N565N3/K25VrAE38ao40Ongm3sVZYY2lfl16MYum
/3rGvZb/HdEd0kHZ6uI9oRjy4As6VFElUaYaLSRnU81Zmodkysj22gSAOTD1
Vo1k2B8OwQvoB2mYUM7kJpX0KS2Nhec87eLnmzC9q9c6MwrhRq+wCun5Sj0f
0N4wtApZ/WU+LBDOW2uSbcIVTufL/eqWgwkfXpXFWXQZpeQExozKbcT8YFms
HaQadtrMDLEmDv6ZAW7TPv6bJxGoCN+4bhk5NkJOh/P7MjQr7LtJqePzXdMO
gSbxYe1ZdWZrkZL6yY3ZCTaDNwgTc8vuB/X7ChlarFgBRSaSpugTU5xZO0I1
SRWANtz9UQuJ1Wnp8W6JyBQbSUgiwEU56ecXy++0I7dE3yYIThBMO4XD/tzO
uUFS/WFl+X4vLaGZWZMfdJfHClFtHS/yfS21msbdVcEHVjxb2WcBDXBLnucW
E/xTEAA9IUH/71vMXsGMM8SIlANOj8wMlyd77uSV/k2cyQyBLWFbQunt8KY7
d8YqV5XS/wlWjB1qBxPIio9wSXpi8KnHmsE9n1JfvP4rnpB/5lvLmsFoDypU
RToDYYPiL1aGuE012d5b7nrMDGyfDe3Ob4NrXLjqxYjOmB4b428PzDRHNnoC
4aJTvuM1g5mIVfOWzMTfO4uuHbby9F5LkvSqZ+0jLQRL7FYOfxpjch2ak/5B
hF/P2NfAPcbfT/pVXILKAAe+ylfmGhqs5X/us5skgcjoIdtGWtzfHU4+tE58
4PbuAp1Gtz3wO13v/YmNwPJM151BP2RrQIj+Fq+hxAgFVbPMmAK0ltztLwVq
HBaR8o17GJr6WBoqYePL+XOwYcP8YHjVErbwzNiC4H6keezsKgPoXYmLlz89
7lGJkrWr68tAuxzFCaHMbqQjrWtWZ7Q5hYsRjB177YSgdKGwjUWnhqWOa/xu
gUxxslVVM2cks+XcoBV7HXvJMjAsMDlGYf8k7mJpTk+D87pwp7ZgZbQEpB2G
I3L7fG8WxtyWGZlPzasJECKGSQD+YRGXt0KJ1rMBQm6WQ5esAO895Ey58V0N
6fuxiC66okjupf6BgdnzmO7r+Uw6Qtxo9Zyyl6osceIQ0c0eUQZIsyJAQXD9
1GHmJ24Xul/Q9E/wa+oAsYAEjM9cKA1LEeDdf3nUbqzXe4p9XUI9x0vPckn8
P6FNuOzGi3vhkNE5+9nRmipPMYHeCdKeUQlVTdq29f1mto+OPv5ZFVfE/fgo
9j6C5omJzzMWvdIl5VEK1eBAyAVdJznNgJEawQ8uveq6CTOCJQzZcFmgvV+e
46N1iuOyhE8krYCQC4lnaEya893sSosRfUmUW4mVqWHre6XfsbP/S0DOHGsg
zaoZh7fVRYk2ow5boEDDkK970RR04KCQDvwX0d/tRjA3MzdqIZv9WdQfAsQY
9FVj2v4a5d9UDxWlaM0yG4q/QbqJfuQ4uGk/+gO5R3dVszvNrxg1HyH0J2rR
NY47H2b1RJPeFANF5sbm/a4/treAQyWx7O/Dn979vpBVVDp/in+Cqo/gkEqm
vquOFYi2V0ww9Xe0h1kDEa6eJabGfjcQk0/T8lXMmHAippNk2hFyhbyfj8Gq
hF5VRcUdSvmIjG4uexVB2nSYPgx+tIT4eStMzW+SB0M8suetogmRJaS3/Pn1
nHQm6/mfxZxJtpP4AM3AANiH7ryj28RlrpwLPj7TNWt8M5mpGw+ZDoqnGZ2V
qetm7308Z/mKoMNw8PogC+Yj2aJUcLKvBWdbiV4kpJ+ALtgh/0P+aENdqcxg
4D+EPcBDbcgnTbvNumV9qqL+ZoYT+4sOsPPWvG/hoqIw9nxPWGViuVZMYrio
LlVpt3qL2o3BMs021eRinwxCsNuPbZa1v3EjsBYuqk76Z0HlYgZlWEE+kCqd
hogZDfX505B4marPX1DlwHXssUebz53IwyY2zBJrJQp9wuszk+LyEkQYLjsv
aryrJmmCIFdKxKktonILp0wpZXJ256UxmfKjoe/nDv7WoauYNXSoiNPnb4ML
/SDAlnYIlimn6GZxt2vCKOwjm3yuRhIwCDvMdmdGR3eaXGYBYXhXk8b+t5Ba
mKNFo2t+sKVjlopS+1KsjOfnCzg1+OD+ubOLAUCmTTTzOC7xe7HPbAiLwKll
7xITrPaHTjaA9k9+ew+D5iM1sYUz3kZJNvcSUuIUtt+FZPUW52s+m+YMSg4n
C18SuxqAZcypxfP7wAl6LR30Su40SnQuRAXlq/LdQGXQDEqCSmoE+/QAUDaC
TCFYDSfm+o0rTkvfniHDCVR/+igVbYXDB8tasULUhSO62RDZzmVwt/ETGKoR
uBhliU4YgE+UxzIGsw4QubGl821dJ7HgyLqUx5qccqoAWF3mmxAu+eGRRvqI
FuQE8pTTNqZJXt4o0gBsNSTZVsp1joO8ur+8iQwjjJQGifHhHQgSTJRPQ21U
sQXNTD17rd/ViytgJP2e2ao6U+Ez6KMuJP/2XWx4ey1rkC/v1l55cMpcGqNg
MJBEpTCDaFqnssFePmqtRfZbO6lDzXWU28eRT+CF50ket4r/y1+kyklAxZ0S
m5IkcAvUbYAgoWtAHm/1IAEbDhfWeSBOYkTu23pY1aTKf2C5kcDdK+/MNXel
88My5jj7CqU1jFueR1nMTjEBtneIJTy5Aunnvt1s1b69aMLm5c2QtWDdFR6V
NdxeBhSsiUuNZ3SrXMZ/ONihbdZ6PLUD1ikZ8NnTR1JBlRaEwuz6tXDHcC2a
0j/9E41mseULpHN8xH/aROixShTxKuRD8TlAa6pkudiracYynecX0FEvPHjn
QFwnVGOcYJN73+e6mTsi4LtYCmGXXfdAmC0tD1YhGtxU0lH8IVLPWTRuMpXu
OMXS9aKRTnVhw7FbDH7KZvddWohkzGOOXWJTbEA726oecxJsYYGGwbmcyMoM
Y6wadkbwY3VZjGmbSjHHhRA0NnVVw7q/2TQuNG1YD5yOQOLJkR2oGc2iXWeU
N6Q5kZ4Yu8yrhn6SFHQrQLa8WJCphIkzXbs1BCi7RQtP+QsKO6KVThTJZnQh
i6KztxmL8070daWBdR6oIe4xO9tXBXCZtE5qauk/SafrmAg+MmZ1e7AQ+8lX
yDiYAwko/1FSI47KROrL2kr+1hcQiAWV+pUda/lHhE2tZFmTplT/x84o8d25
MO4uLrGWLc144LToachWiuyzIiPKz3sRJ4BHOQEJRV08Qu0qDtBkkYInCw7N
rMPTUw1fwdIJzuyMy0S+ZEiWY1HMzeiBXnyhsQc3mjFRtjMmlYPH8f1OOHE1
sKvQczEZZHHX0waJT9/f4ayi5LzjQHCcwsR838VzxvjGEKrLijVgfXZlz2VU
n9UxuweVgfz4OJwWq9oUpvvApR2YYlUXJvhJL2i2M9ak2KvF+/7VlJh8O3Qa
S9NDek/xjs7VioKR91ho6E9A71RKTV4cjbVkI7S4+6WjYQnuQ8XGALsATPIf
QfUURbQ4VUILn+RkoKoamG6XzD8nmhWIPcZRrG9LWtTM8ECTXTnZzFAVgxW3
e+S1Ktan1DeSg52/OV4nziJkHxGpcIT2azAqEnY2dbXTfSt20bnIGKEqIkNK
BxTjZ4GBGlSO2Rjo57yXrtL6CwISDx3sfC5EJ69fPJeRdilwP2ObaWR2MEDl
Z/xy9ZvOKwNeLvoF0/ks71Z0hOC1Nrc+nLSIBsWYcsWUrZxMpxJFFTqBgYPz
hC8AxfCr8IjRZkpyXxC3g9n4ybUGQSl5SyZxsIoQeOgGsaUwvqI3+HoPTRPP
yqbNoalI0ly9zAhWiQoA23xXWtj9iIg6PrhJbGxfhoceMyA+OEq15NU/B9uV
1hNQ32c5v4K2mW54S+ZP6/Ciw6TX4ZvC18UPaRHBItdrtftDXBvyUJ2oVHBK
D2sV1DhtKLtJiDEAV0IQ5iXaJLqt0q6pphHHKAJidWZoULfoYN8b10tMDt2O
e7/stokXAnGF3VqDUojVGzCsd+ieRoMRdu+nwZkkZW8Z69jwXQEa6YUmbp5q
wqu8sBVv0b5MsEPlERbMkN/sL6iG8fYpd+D4+ZTUORSSpBZOmIE790LjkboY
SisbSBa6T7W0zivjSHyRWIrMqvFWzYLjhM1rq8pu2ObW62rw3jIXlZkM4CZu
0nTKb1cltOqQh3wlxOf5ECyLYSranwB0OmY/mPgAgi3xvZUMU7pITnFQskue
wBwFpnJzHwoIxcIIRC8Zy2FHQzc+HVUI7Gl0fe9VOuTE1f2+OnDJgHk4/DnE
ESe0MtdL1DykyzZO5JExV0uogBOAg0rdrCvedRaEB9rvUfsX9WpwVwcAcYcL
ozHdEGDPbeLNXxm4M034UFyusuH6pk1uonH8pBGZfM3S+VV1Wh3ks7kz6RS5
VoQpn4dAzDqrL76xp4+GaehZX2nmR2pnyFVaOrJBhfFnflU5aRZJwKsqH5XD
w0jvl0Wskr4+yV8SB+mMK6/F4QTNVIx77+EUxBORmO2zBr0zikDATZ5DGu5E
2633K882GzeiZk5w0bZIrlnk1U/QfuDbXfvPWtfw8oKONf3Xj19cxi5KaNa7
PogCr+mGT38cqW8T8XpXkKzDZ4GN9h9KWtg96s7lyLPejHdMqUE5Q10LdKJT
45v1dE7wQXsQz+ZmJfo8wtGofzWmTtRQMRMDORbzcWBZoM66W/LCYWzvUaRU
5OHo/UJ8tv6lYS9q9o0S1xacBxM51xcfsfGY0C3QmBpupJ/Kg70YN7Dro3q/
OmfeiSJpgtLoYYg4TeUK7VxPEDZp5DWMoY2Sxn1N3faypIFI/ACCvBQDosRn
VsbsxV5R5AMWErOVR2FOaQzW2q3FAPOJTvEsHpnetW1TrXxMC2iBgbx1tYZx
elYrE0oLIS9NzX3L0FJKqWVP9CW9GS2/wue0n0VYpHkOtoTWlK5ElfEykrA4
Yfuos79uAdX2IPvdna1AjfD+avw5T0b9XDpJW6oBrxpgnT3e1ooWUJHXNimA
hbjNsbxWltCR01NyDfLzvlLqXiS7n7sbfWMDdsWDqmG7Mr0P8bWxM3wO/9n0
xqZLavoXPXGI2cjg4B9GEm4Ju9SXn7rHpwsaZLDDSnX9oB6lC4kFqA0gsCra
kpebl0Vokw+T0Hna9SaaORl1YU8ISm58myU+ncJd8B28JcTeZnMA3U2Ctl+m
em4qpN8dHhosuuOIJU93/ivUSg+J3cNCrPWNmjbWCFI/yQccPAN374NCuI0V
O/iZ2El34Kwe5S+d5sgCbvZjj/MjBUtDIWIXPIclW3N1aXI7UlLDW6QKNJjz
4BgaZds6AWezsZz2okOTkrBZqbLmlU9byEh60s5REKv++RyfegxrXUvT21lo
j2vEgYS2/Mft8pP+8XN21SAW6cFf0lFwy/Ta9tXEzH61HYN4xNrYpX7C10EA
Yovhtl9GwQ2wsqwTWCOdncJ4yi/zAEZzZ6nBI5zle+HArX3qMy3WWs0n+bz9
6Grf2uSkxiXiXfPzFF4n5ehAn7NMhcCwsn1A4oL5YvDgRYtwxuWeqy1ZUqeH
TaDGkXd5MS0DCe/lBgT36xijb8M7wV8iV0RHpKVuu1h7CY+N0TuSsFpWI8G8
P+SdfsNQj3N4VeL6Yubxnb1RmmW/TZ9Fdbrtx47dvCY1jdbVopygPBhJaYMJ
Hd0sPtpJkPyTn2mmNGepkYgHTpUCiDAi/bDGfnIveGXLjxPPviMgsL0gF5FM
bZzkkZ46T8VnZay3hlakJjJ3OW0Ktb3h2apjRNbKIdUB4jwJrw9KPU1hcizD
Dbn2jFaEAUOwCKKqc21a07FYxty4N+jxk4eteU6ltS8N50BUWxdmePf/4Ovq
v5r0W9mdbvDXqifO+S5hqKg3KpfTIRnG3iSCO3ERR53+ESy21F28WtuATciL
3wcicHzz6epa/K8meocmmGtCit62pE/QXRfn51KqJmV3ab8UoggzFMj/DMF6
FsDhKmthLBUXlQqADhm1z3ER+VID5XCTLJMKsjg/nKyxGY/IeeqWD4MeCy5z
Vop29ICs6uqhp2+1NvL/662Qv7f29TIjfsNch+LPhfudUPGMJhg+lCRGidoS
WBLybZOEHXhzPMJEO+oOOKQ9iK4denAZ1S5ZWDqLdVbySUn0c897U2vmmjgi
CXMJg6eBQgNfUb0K+YEDnI2IS3aw73xVzZaQsDOu4SJRXFFsveS+taJcY5Yo
2mCnXgJzidDqfD6Dc3rFY5vgbAXQeRocm8jHP/u1QSWMYvjnYG/XJKacbxVm
oFGmdgtp5fwoWTuXfs6O9KdKzLp71EnQRBxXy3shsTgXh9Vhvz0OjDSXJYdD
arV3XjreK+j8zrhiPuaszBMShPl0YU3STwHAO0iT/ZKIgPfoHRfSuiJ8gLX9
4rNLMFybocBB3cNn6w+Dk0t0oXVO6PVT4lQy6h8/jizaniy5/FAEH+q0ctTn
BBbehqiH4Ww4dIPskJAqNW+xLg1n4Bgk67OE5KATRDJqyfT8bHnH3wZSSiZh
AutaY2bP9yRHSywYVIv9l0//aXC33Qee1pLAbP5OENDveDddFEgLtSImQHCt
1vx2Yo/42YeKVmSuOcNYcyUovkPW7wjaF5iWBqeWe/2xNwXq3jhehQQVpNZY
zqrlBLQkNoV6z9PStQ4J7oAenubNcmsLpzx+puomC/bBKTbcls2rtdv+nvTM
l1Jfl9RkZ6CMaj7vDXlowi3ffJxon6az88YrTlaj5ApiBozn95ZCLZJkOlQP
GvKkTpTbAiAPPzAYBNtHqfqAsSUynu+pvN+72THbtOr1UCeIm733t5x8dWAO
vxV+dOVX01piGpOtmBMKWww8w9BwqX0EKj9FLse8v4ViKVoErUculRHQeJHF
LjzJA/jCcpawcxsb/Noawa3/72dLmgQVvKpvgAXhCX+/PXoU1TDxw2xbVX+B
MBypaifDq+9QeugwDuuWHtP7fLLrkejz7rv/mfb/2o5UGy40CgErKj91ShGH
vUGWpPOXU+0PU19xuAHSTKMcAGIdoEUCcXOQSmICFOqdFP3dA6K6/4zMlA7L
Ju3B2Lx0+iWfQCugxrTwWBgkdgJuobGVYrhFRSQA2edPTB+hE79Dzp/e0l2v
VNWmblRmfkGUMHFV6ci/wVG/6WhET38oeuXGuHFkFuH84A76oXXCWMdLSNo8
ANu6n+MBqC0n2Vq9h/dgBKqein4bk/OHpVRxXk4rJL0uWgrH5EiXi4A3D+0e
KS+uWX1zSHxFSozIm34naJ0i0y74xFC+gdO6AF3a7VitPyx2+RN2ApvdUfis
hM948qP769TRux4qoSRF0ERKizF+jndQeI3RFuqvN3fRXY9ney4fkVAw0xA0
TNmgBcPx/bXB6wXnmn5JxX1rkzLoG9j8Ua1HrY/t4vXUeAShEwjdshEn3wYK
BaiL6l/aL4jAD5ukmni70YVwjMhb6TKAMuhvWsIzUE3lMw86oi9D/5+Z/KHr
F4QiFgAR+w1rMX8eDRXS6ErALOpqzig3JOjrXhc/l8YsuBSx84aVHV7dAjoP
mdEGuXJM1v5IbazXwNCwMsLjPkM9kvwFM6n87+Qujzp6F4VWjqQU5muygu4H
YIpUhZ0/h3DcZZic9pk1H9Og15ktLvOPAk6C+DDDxaUd3l37Bn7UK56clq91
JJ+lNO0ouLjbO0U+JDxTmxLXcPbsq7f6lC4FffvglqD9DCdmiobMsDIDFiEv
PEdFN14/+aNsea3KxeD5OoHW/M39szrwYEHr4yb8HzhMUxfnGiq00RK/z64b
SZO48aYS0A1eOCFvdTFQvwNbnznYzEfvz5WVWprDF8rFhc/vyz6JC0mab8y3
eJJUioQI6BWewqKhC5xXxnUCP8w7rqeqLIeyPvZdFi7aIk5VIcupvVn2g+7Z
CkoGrx7uq+nNjtRij3FdPzxh8RWbOniIwm15Qqg2OvNO+d7pMgYXeoRrqI/F
NOP2bPG85XWFog6NBXXTbJHoRPFXBJmyHwjOZ1ShPrEJb/GsSNoGVagGJvv3
/ZhBKHd/dIIZbqqL3j2lbiotezdwxVHecOEm2f3Ih5dxj+SE2YSoWQWJmqIK
CDUcbC7DTtan1qRhFCYavCA9ZDg3Khdu3LrKJquG2m2IAzf/t2Ly4uZTS+BN
6Tff+DQMNCZCUfP3qCEFudm6YuYVrGii56vUPtANnR1QTwolbrOdAHyI6zo+
QcEvjQvJAFfbWf52mqut4ZcEpE0hHwXxL1VFruvwsizfXL4Vz57lD9bESM6K
qeyG+P25UAtts5dE6+xbeIaRP8hF6KRzmZVnGRBPZJ0hQ2sf/kRXzTl1xAhk
ZW6mgsLynbaiDY2hJUFCrcmtkgaMHRuwQzhlNWHEiYZ5eiKwfssGJvTrYTHV
RFqSfg//hchziDd29VDWCpaSZKrTm73osQ0v7DKi2JXBcuA4NM5rGvPpvcWX
dK7L8hHZoU5hwwx3taRR4u2xsO78+A5nKEfemjYLYi7Qt2/Urdn4oAuqkQxx
qPQ7IYljlksc4xcHbEG0/N14HNWXF9bhUwTXYXgROz8zvZ63aHBIFo5VfMGP
iwt0CN88rY5cHFpI2Rve95weKCwFTugSDy/WEy5i2KDf5VqnV5Oh/qt56CT2
ouc+aQ24BH5x8A4vJpj+/6Tl8AZj346Ow9gnlgt6EgkEbEXW9cCfdhv8U4G/
KpvHim49BXPO1vxPKEptWVvB+7fi06fw12mQT0rbbZvGR+H8S/imnUqTvK5n
5+EL3Cjd1+TshSlXNFgrsFb46Q2oO76mLihDog2SDzhwY5jrS89UOzP+UuhB
GSl9plUU/qDpZiWroRbWnCgwhev9FYouYl3b7WmPCs4acciH1QkJtT8Nmt7t
zac/VN0YoHqYyGT4PTWNuCPpYikQo1+d11sxSW6S/E6SIzPjQe1clGUnTSWh
sTqQetFzBO8AM6It6zARMOblkfWLE4Nwhqt8/+toCKmeYv0fRSLOVJoBYyc2
F8Fl+kiv25qMae4nqgP7ydCznee0Rx/PGywkaUji29KLKBFZbVmV6Fo6LMYn
0MKgP9Zn7mHrnhI+ADtnHFi3FDLBMoNK+RH6wS1J2uH7ChKg+EfFttFbBFI+
x/EE/QoolmNOotz9Kza8oL1NZS0tNYjNsYcdrjIkFCrn0k1dD4o13CFYljnr
84pRjzynHz5CTT65YNaR06qt4vvzJLU2xHP4Vn+bStqTBnZmdAoAAXyQANkg
NV0kHbgT2l6GSCemXZRJOcim70vda8sGUqrm1QNRtbICBvIEgpODXCK0qmaU
c84++Y/R62BRWFNHtzxzgE2VQl9g2blAAO+PxMsE/X0yblCR6hFm2G8/+Mqo
F8SgRPliEbh00UH2WgevnsKfSSaKPU1/2DiwnEy9lyCHxVDoF4FV0JiJrCsH
5rBKJRW1ePuWredmJG47Eyu4HROFHac3FFpsB4+eK8XeQo14H/lp4/Vw8Cio
BzYJWZTnCKKA9CvUWcxg7kg2x/rKgCMQ9JZND0xkesHRSmkO9zDGR8YczbqT
kd1ZypPdSWlWhBQnw8pZtT9jHyh/zXNWmSkytTG+CtLjXt4BUnblie0KK5Zk
vn5HKiWlHD+VYUhVxCSKmwjhbueJgz3FRDopI5k/TZjQpgn4COg9uJEvL5W5
gqZEb9AVvu7zfssN/Uo0E0Rr+AYC8jhJ8RUd7UPasfidaLKPLU69FPAO3gcF
aEtNRM3Y8jXKI5yR1wdZZR8/92iIsielaetmDxRMZWsRgqRjR9+eACeFe+tI
kVa6hrxUpOR0INxGddG87ijXOhuucqKl16v2Uq+T5ephEgvnicClYUxWIot6
7XgUZOvzPh8R1sKS9pPrxd2+qwmnCE3c/2ONi3+OrygTaWm4h5lNz5Av5+hb
pdCl0/DjFOyncL6a3CZnGrJui74htfujkIaYH9u9gkvzRgJrSXT3GYIKWpEO
Yw3LR/1xeNBWHeJBiYyryeC++EpHIIcUuB/mQpomsFs+fu7CD4RUjbK1Gu+t
knLzlzVLiY3n07rWkcOk1q9vtG60e61pOMgxejOXffQGQDZdkwS7cQeoR0Vl
3l24XcRyKP8VRSwl5FjX+f9q6hbJttF8AkJNnsyT9XEStO0Z9bumyKt9l4W4
uIlBUrTx4M/ug371zBmpmE6TEw6luF+RZaH+Wqld0K4v4KkFfZ9uuWuOUITA
G6Ii0oPHLwqaa4WarpmRBbVVNV9Zj05ld8dVuwk98GqC/Ue3JiS+up0PBMxy
JSfj8TbPos9J3q7V14Q47VeRhJlTTQLqXEbaLbstMHuo4AmJC3U0HGkOd4r6
CHlrXp5QQFmSB7CkN0h76EcZ8+wP+pr/RoabfZ9XZ+iMFrEFyBuMPijeQ/MK
0q13nn1Ju5lmzJGUh8itGkBqU5lU1uXiJ2AEH8kpsY8I+VdLdzwbBQymW+nf
XI5QFVGPN7PnZ3LxX/MilAHeLRoCRJmGyW7CVUm5eRA90dqVjkOQq4XGsx5Z
6WOZKLKk8HFz/OLACntQ27SO4jKYQzmGSbDUBKp0XuescEytF+yJe0uXYTpI
1rkijI+lAofpScrZT5V7mSiuiCgZcZuPFiUwMVoXvPQg35uwFdPSyNkWuzQR
4wxs1fhEfN1HIRMeBh8U4uXT/TntRTQLdbDaNeTqFlMipM7h8NdxkqbXUi+F
cRby7q5hB1Uzng10B9qDBLD0oMmgPcNr8R+9Xg9y61GvC8YBF1MvsskskbYZ
OX5z2WBdaJGhCOaPR+QaiK2iagUnnuVBv1rXrk42iI9oYtgLZ+d/PZn9fFr4
AwJ26AsZfKjZr904rzHIYk+lmji2qstNjmxsHC4aXYIF5zxUjQiqe8D32P1n
/T0voKDJJJWW0LTPFZvX1OoO7ayzilalTu9FG0hCiJOLw8rEQ8F3CUu9zAKG
Xk4apTa+6YdhZ/2PRv1xS/qgPj0Xo3THvJ/XGESsCkeOp1JuHaNRL1gLelVC
/HKhMUkiNXfDawgZA8kK2vAgeikRtxERphUkg321JVcvqIoaqzWO/6UeqXGm
8JnvhqCwj4Sv3NRI99xIKwJh+PJI2vGDSnzoH3WowQ5yKtJbkUKg3WipA/Co
bmViWVk2HBhSVcOHgcZKiCfe0o8HR1wjbT3cx5tEdHDJVRQfp6JCl5Jk1AIe
VJMuWWvkM4ksRJJH24EC/K6K1PvmuPml3WWku0rsMEUILGW5cIM+7ZSvDFF6
hsEP23yzBZf7FpC2LKXAC+9BRyHfc6njR+HQz8TSFPeDqUK+9Gls6EPtraGO
BG0Izi9gEVJKpYFiEeAyzR1JBn14sRnZUlpZndxCPLcYiJjbwiTihKT7/31/
gesD5WAGDISljAXQ5InM56hkV0x3jYerM81iOToa0zT218H22+GJWeR8nUmw
MZtxlCtc9K6WlPtrou2r43OZ5QlbctUkz6CYyEjpigA5UBwG2Df7oaNdE8dA
IAuz8YpLaBgkg+4qK5BLwoEdRoMSbJEuemJ2f16xOaE8FQM+ALFELUpoLQjg
v94tpHaXw192JGLMq/uZLa70nDaoAiCHt3oQQrfR1sebe/HosArfOOJoQgre
17tGGxQ9Gvd/kVgVnrZCYK4ll5IvwCLCfR5bC/X89TKiMaBKFuD4oRAHaxbN
x1qHQ+SnWssh6gSOEv1pg3jKDc0zyYz0PsuWMZ5ZqCRFTC8zADDyXSS3jRQS
P+v0XqZINyQtbC5mkXr9wqp40lU2ungU+0jNerNmAdQh+XkSvqzZx+pEzT5O
0CQPgEVug/segWbSKIMafZXs2mKmqY6NmaNA1r2tqIj98UaM8F06iej3qyXg
3FuMXzj62tEVXx0lXVgl5QXd9LmNUTVB84BEnPznOjgHnScR62JRYviWdwYj
DuQytpECKrWRU47N+L/72I2YOraSA1SMwkHDJYJnsA3158rRc8psh1aTmt9Z
CAUTRGSmi0TdkTGYAPcq1NUbPCQeDSki43+mcIda2tvjuGXxX87mJ6NW+IyB
wOKsSFBru1EDMINipMFCfYpwwBVims71cxN6hSnsEemw+/X/BPkGe8s57lrE
5oKFyyN1t6ZG2FebDHhQRCgdQl4lPNh4oL2ZhRS6BOUbYe0826xpzMWYHQma
TbJcW9YiOUK5luO9eMvpA3U8UaxX4JfhmIzTcRmnUErarrRyHHf/YpIQfDe5
OTiXdL7+0154TXO5vP4KpGP7VYvyE/gAfS5mXTNekT9ooaCiEcvVKfTlcFi4
FFBUlBOF5xRloV0JO/zvNyUCc2TbiAFPgdT77p4+93727G78uFk5hI4sDmdY
IebWyrRgDLqbXqaVj2Pgu1WkFKd2IQ1jFfUtcRTaHp0P4ZknwoIsyUlvfM/r
RTHvMnnr0NgVP8qBHNyYuCAdlcvDR/T0mykx2Nou5hgJapwfceUQJ2qbAl4f
LDAeTa9QbO8FbNf++T3dvv+/hf5x1Y8Nc1hrpOdncdlXVbxTLw4dGgtUBwU4
6w+R5ZZ/FS9J7HBf6QUy3fPdp17xQXFHBAn0kDkMUDpj7RzHDOPVzVNyFeBc
8O/Ae8s6bmIhDQuNz2vzrfrOiEAZhRO9y2goiI7ek0w4RiIgZLNirqjLUXiK
aP+j4/1eRx1n+98QG+WEpR+fZt+/wtssSJJQ3AXvjIgzVHYhQxKEyj1apgOg
LxCPSZsrx7wBy8fzia4sHOYwlAcbhvHHL09fyLBY7WIUFvS4N4SC1Jel9rF7
ZWaLErNwjK9iKMg3Wwwu868JCfTGZFZ/WtCRDSFsKpD0bHIpZcAhOivI6pM+
lbqcpINulTpc+OAbttfXGXcw/mOUwdf74aEzmMuj0Uxuc2+Bn9G9dXR1ru+n
vRhahrN0aKwkPeAq0NLBE0voBEoqqC40wVBsevqlRxUQ2Z9snKlHhn4yZ/aO
1knAEca4L497TlcXwSjmFrq2JoRZKdmNj28UscyTa1AyuEl1ilqgkCuTsx7O
gIHZW4C8wW8DZ9MYcRKHO6k4s2XV2rpJioxtATndpOkoyBxqTamq6FbcBBuU
L/+FTjwJxxtJY7sdbtMceMmVW7f4ihvVZ29tu8VbaU+f6Ir+d3Tu9ivcV1Pp
kDGbfnKKpuVL6w4ndAxROmQaNFsgO8zSKzLAgPlTeKj5zSxap2l6TSKiYqqr
Fa4wGVYLtyZflqz7DBFX97ak9P/k4zXBtSuTH2M7svJE1rHG9xTOQJMzYBWu
I95ijAGTNtDVBj6j1N8eDYXlbFAemlODMhIfkfut2wb64Sd5bj2pHgapbvcs
VTS7gYUmZr2tHt2dfWqn5PVtRT6kh3eDzP6+C7eseYAEl4wD6BtLf1V/kujR
ZDAdS3pOWkLvYnAZ6xFe2KHsWMkr6JTKqiy+YAdhGUIlZRttnAnuVSEskfTA
szAgik0d8ZuZ6qODGmF5QleTELbqp01Dsm8JwFGFBtZbckCV88I1wR3QMcrn
WPRxXvqq6ijRCUXwjNBDdMNIcYQdfDsTLr8WWcVgSK8cYl426QKgRBgdbhME
JMZT+jo8mdYPkQedltSR0He/dJ9vxdwIbsIsz7CK10FmSCp0AKKiKkNZlkV/
GJzyn0BVLu/jAieR8NZgG4GDF5jBEmHYHJFubtnI89GaVRBIU5EysUviBmrl
sjafIMQQT635Jcu4zMN+4Z2nvsNfV9a5JAZgKl+5dfqFmbs6g+tzZPUUT2qx
0eN0cLX28EmxLNbhPEDWLmNJI7ZrTIl/9BBV9Oy20BBEcpqXAjlVPJxs7i+V
9LNK7tWpGXN89XATVC53IIb4zjJl32r09KheEoJvfb4WVlr4m+01KAwrleQ9
QQRCMLLY5v7zS1zUWIdAIzv5IOwlKHxPXhgFjz3gTm1WxR8W4010O/AjZrYj
0Ov3cxUek9cmMwrkv6jXB+KUMfcVx9IMWnw6LQr3ttWQl0ToF0CwhuVOVvFJ
rK0wREq5kwACwmeOAIIfyHsoIpNvHpAkHPleaG7ZtCkH4cD4laeUF+97VIfo
/xbBYIjj7uHkmSDwFCsJMJqRnnlDNH2jjn3sFORGg8opL6gcWQ6UD96gBJlE
5ke4HnukLdofFuwM5nxt1V1vl1PXvJEx8VgGv7OYBEIB27+GnzqKfQ/wNufu
vpJViP/vFVuWnBJAn6G6EETUe4E5U8vszA1fgYieGZbIMCGrtEupYwXvx5cv
2FPrY3GUIKvpKcctOdevjXjnVM9W1kF4bnTtgRxai6cwBOwVAr4I3w1u4qEG
LoyWzMzyYPxfbxLX8TKfSyA+k8F9DnhwdfQmc5Vk2hD/s+wB524NqSjQ7z9y
cqQQRKKdpdyvlUbcXfHoVtxkWPHbQJMekuq5/YQ1wCjS9e/J0l4GlPjBkBXm
GBhMZQIqY7rt+Qmm3NTf0uu6Js/6uavi/2co5HBLeABfeOIma5eDKlFUVJ4b
e+L4FeA9O1/cb8cAdKDfgkTCZ7XqdfqCaLh3l3fXr8O1kLyQmgeVlrK952LP
LQuESd9PEh1aQhyq8UtW7nXzN5zJWxmfKjWeX0iIxtKuyeZxkmcIKQa4SQyK
p3Pc0F/7cPvvvImkeaIdK6qsMy94eAOTR65UoJAJbHruHgq+QQ6Xxqzd0RE8
3e5u9Q9t0TZeoZ+emFWV4ekx32fkL/A7bVYOn7iE7XRW7bgRWKv5GEspFIDk
ZYNUdnh2euy7VCOvr5KblSGolzYKdx1GIhHGQpCLqVPXBWv1CwMo07Jj6zuM
MFwjGMnb2AOoXoVgLthX66WRw6AGmuvP08pg2khcwigOpenrV8U0WB+Av4rc
HdS+kbbUJ5jryiy4LYhlvdDHEoih7+EcgnGr9073AaaGdpClP6/r9ytVXXvo
IF38UjwdXpuPFDF0uY5y7LHxYe+Nuv/HHXhAdrFuUWdO5GfWYUCSCsOBGOpx
6YTxgDn+ygSUNuRP7KYpUSBVD9LJDHmxLmGy9R1M1oVpLSFYlv7mGMyNRZFW
lqVJc8PSMJ4tjnVxWqzsL84qzAomWfDwjOPFU9s9DYg04XvmH+ibym3Zzt6h
K1JS2BvNx/PbVkEJAWvX5QN9RjasaKg8vGjneizdRTPH3ubtUW3rzbADFeVb
YiV6xPZOSS6JAB7PajA6OkIxj1yupKjSgJC1LwSBPs0BHovOUTcW6bhGF6j6
2eNCD779HA+yxPIclrZH4VtbsF0fvy1eZaCUds3CvnjNPLhKntAA5eEO0WV9
RCzRvdsn3OukAkduO9a3VfOMVAajdLFkhPkWFhZXSYnK3r7fL2VvMMDbJICF
SoxrjZinAXcZOJqiIFxm9H5nn15KnrVEZkSG7tOXXW5erpZjCla8b9AuBHkV
IXx8mp1IO/tqH937Jf305xj7OS7fFJuaU7kC71VJmHgEsULyspP9eoHMT38p
dMVbBYwHpX+GiNyVUJed9DN3s9vjClmZnyFqDUpovFmbelGMpqjLv2NVgSBx
A1iMS2Rbo4DUIfBCFqJRVtiYTk5OwHcA1ogGVo4ddnhyZECcF80pFOuPQFHR
lGNwSe0CBHo0af19hJ9NoljqMcw=

`pragma protect end_protected
