// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YK8FeONx4BDdgm1YjuXCFTSoQBdu7jE5xCBNxjbzvbbkjGeMPlLUFYzgFqGr
eQJu2+XZS0tXUL8hKzPLmqnBg5n1FL9XZbiTUj6czMONlwzRBJVzgoO27GeV
OH9ng/Z7uw9xa1aVgsinEsGZVyrSb7S1F17ZSOMJzLteZyQdJOR2J8jXb0JB
mdjMqtbKwY6f7YpdCN+PH4VOdp0URgkBgUBxW/gx+Z/l11Cy0rMzUxRdic/N
2cAeGIpB9eFnChm7RXAONz4Wt5y8/jmE3YsQ7W903/FV8FlZeIpF3t8yiU9f
+2/gKmZ6hwRDvcvxfhgJrHzrjrWcwJl4xbLoW9r9nA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c0UT+GMvt0YT4e8NS21pCMLrg/eipftT6EL27YxRsShJKKmySnjThW0GQqri
jXClk3tHbBiuredQ4Rfj6VCQykSIP013v7esx7SKg0TabthipxZcRIhqzW0S
guaGxKtMVC5EPvlTq4izlo3QkGakrUA0zt3ooyVU/qDmiZGJ9+LvMb9aLnfj
H9DyQCkfldN/4PnLySUGtYFhAJGhryL+DwKIyzo+WcbjNEFZa4rX+3NuuNBK
mRKGFrob+JX97KuqFpeln/laIIlwBflf357Xw7VQEkqIwQNS5Yqy0/s0Yx8E
zYVLiCTvTUThsLgCNkC8PTJe7O0CQJJKc9PzoJqZGw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gNCLUkUePA8hGm4Vsije0DPsQpYj1BqwtL/EfkjuKnZaDwpVf02Zdx5Pd/eI
xcYvP9LyKfu1YqLt3MwnyuRGhs6FSe42OiaNpA02V2nbcyQtwwxNPP4rYyZc
/v0mffyedA4l4CYSiQ4Eg2VIZUPS4mmURebLiHAV4SZITpqJjrlqXtleP0cW
bYjMkX9Mgf4z0cdCZRbcgDil56e86WYfXQ9Dc2vi6OCOqLRXFxrgwngCqph2
cAbKc6o195xBJq2+5pL5BsqJ0RsJTAqA03ki6e8qQr/wfi1V99hQCj61TR+b
meDW4pObD8Y8CjMkXWbDhd7YxN9Pnf+uECqhUOTW0w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p0/zozpYJAVOg8H6HCaFRAqLn1V0OFTDgJuczJr0NEzf2zQu6JbFcix1sKIe
QRonB99Hz6LoEs5OsgxkCKq2ZpjQx4LohYasKMvNPBJt+8keI/dm6B6sWFLg
8zUHyaPNXmYy9TSfbKpzfsXu/4+WQkNjOfZWHek6lqgmSOUx2xA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HLGQDOCmTu6TS/VJVDhmzo+8krtGDQrMTKY/h7LpjJBftuItgqcA8ZD7Yo5C
E19AgoTLdCtNu1FIhlhAh/WMQ9Msq3tiQm+DUhwqydxhS+EfiYaww1M3tUzD
WtiAE/SP8v5k55xPnfH0bLaxcnjauA8F9vDGav5RC0NxIR6o0zK1xS4s9f/Q
jEXqSpKPpzgVWi34liq39dUXhS15WkmN75hRUzMrrSpQh4cbgC8iFNYOBsy7
Ft3wwE5ebVart3J51DF7NtC3Kq6rP/z1iJ5+2HK/mhsEAOSV4c4HAg0xEn63
pVdmhY0FTnnY8+JWIHvsLQ68WgF1DPptJAo5xQX+pDlEu1sszSGhhjKbA2lZ
9GIdygol11MTOKn+gfkO94snHETmR0Vjfgg8fvOh15JELcFEZY8ISnXulRYh
Eroqlq3/b3E4mo6xnlvdjdI5minhjVT5fdxJyjvjXBfz8WttwKjgkiPPuASl
sA89siPvoeLcLEYoLC7wABbx5HIx9vuy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FrpIyNCnFx9Mhgck2MGDcco7UHFeRp1hZHoLf9O3/gBIEG2o3Rpsduuc3KmQ
5M8apGZAQMDIoP2RlHHJH90hlYSGnmFMR04q6cahO6LRaM0k3Sjf+8OyGJXN
iQhmF0iDjScWctp5UE6ppMJqyB+L8uJdlA+e9way+Q5zzmXnmwA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FAgP+vNG3aWSb8YKrToYZv0Rz9+Jbgf0ccVd/MVuMRhlBVQVY0MrpjVOLtuX
7qYhOQTBY4OowmcjJuU2MXpNU+gEORjpxINW+PXIjJ/Fmd93SRSW309OzB81
MKoqwJlf2HNNpRanE0kk4kghie+U4SKA0OrIY6mb8RyIgXqPMyA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 27600)
`pragma protect data_block
Dm4r8YCik/+LclqQex95AO5II37Mhimv/aVkoKA71RKuVPjsnXRsrUhYxTAd
0E5hTBhh0l9CavpxnBv9SmMHCShINPdgXXbASdBPCMm+/3RBz2KN2VUOe+bl
9LBebsAu6F3oYYYoXW8n1jMBhvT8VzkfrSX4sZ2R/YQ+QK3RDOHRjvo+k/1M
KEGe0REgSY0bDHf/k3rN00PBzdo32IPUfEPYDUW6jQNJST4vooCK0DzViLOF
GyvC2+STUsJaFkzC/5dV47k1PJJOETe4an2cJrqQkdQ3/H0E6/MgsUU6/LQB
NACGkNc5kHdqrEq7fI73L5HUEAjCZAv/FL86OIeXwYY3Xz3Ce0bPCVgmsBlj
xt8pZEDCenc3+WuVTwxWPHGa8ulb+9MEoP3gQ8+P+idB6zn3a8GFVRfgTArB
+pxihWEj/+Q7pZ/K8kPV9XJkv9g1OSmRtQDWrCRVt4JXoZNnv6Pq9HQvcFzb
ihDSV9gsJf/3egPBmnem6dU42ePEBDlnbS9xHX1Iwi29xJl4IvD0J8BpDBq2
8dcwOTPCM/ZdzPiAWudOj3yUYmNSGH/8sp+Y8L788zoj05YI4KXGBZi/cskC
gozVSK35cncf71wW7RPR31Tx3TZseGSw5agXWz1n10PWTQruu9H1Hlx4yCmD
emAQkbBqSXM5bQ/CUnf8lyi/ZfmHBHu+FMtPlr6iNhz11b1NNAh/JotR25OI
dh+2+jdgvWxPi9yEhV/AaLb4VMduZ4iuoDeI0LEXxC+Ag/VrcKs05ACeUN3s
OMDRUts8PLy0sjOKOJGrb6L1sYFXcjXEjiB32f8mB1T+1Zo/Ntc7Hi6HefgU
Vr/+lwrB8iKSRst6Kzx+CZtD/uha2K8X/O/HmOpQFdFoy6+sbFY8ptWh/toY
IaRD0BByTDFZx4tEHcz+HBPzKcEWJbzuDDAh6Dv81egcOoaKCXW+yZ2jQmQH
FxmoBTrgoF8btu83hwcEhLAExR4Q+Owx2CR92YcOrUaOGqXNuaRO/s3GEhS6
C/hg0FlD2E3e/XTJtutdpv5uTGFK+/0XpQ81NC8WwXTqXwwgF6Qzs8R1yZvV
cQmnZjJwJpTS3mwwCY3Jwaew+zSyp2ZV7gv8QeDcy36SHHmtMfjXQK+eBHOL
Zf2OFwk452lTmlYyGuH3yKmuzh3KEzMtDpokqQ3Gh0Yu/vtaOtkqVhMGe78T
L56sPwoknCee2Se72Mn0dFg4yL5mE35bMw4xnx4cThrqzHW86gdaH98qKEEQ
LROfcIMKuOqsPp8TW5qrvG3JqYeSmI/8ffmD6yfJH06xp5W3KM+iJkiwTMX5
M34QQwhENKnUN7S2/NYam6S0XlweIdLZQ5K0OuyiVMssPPVtjuLKNIxYUFP2
BWC7qcLqg4JpvzcKs6krepWSblN8EyjdIRze2fynhclkAqCTFVX+LBnx6pV/
jumJek4rO4pNSA1pWDGkNkHsF5TRwaK6RfTdE5m6lUufYA4OHhlj4NEg42wu
OVrB8mbGqCKDh/h12uyl3b0oj/Ci23vDKb6ASgEBKJYXeOA+0Ip8HBRhBFRV
/FUMUZC3Nu7M1hj0+vor4WwVhVBGhhnuyxK0ZqQAYucy7vMKWh7gLRpGJaVG
kZMkl+gCJmfiWsmvPGwY4v7D/AUGkfDmAPP8eNP66PrZHe7DxQmoNWL+OlbK
qsHKmGzJuesX3zb6CZ4FKY3t8Cd1GBnP0rU49Q41wvVyNXsqwS3Vq4Cwc0NA
V5Fh5X/bTLoFGsx6X+maaC1CQKxof2lQ1GAsn/5RyI5+JZG3wQ+eqob9mW/r
bxXzHH9lpQ7fKMFvgI88qAevF57Ig3Or+7eWMCW24drZSk/G6vuxeVwxuvz8
liTRAPaZX7jo7XUKSn8Pa3e9Qqc3IcptmSAAyNMlcjtuEtVbYRX76TDePqAf
iJ2DP5a2GzGtWisPciSYvBx0y4FfZjZff28C7YZVWcVAJAmAhTZpFUKI9EVg
um6oFrWvtUHLzrfXRN9ZPjv8igXVXEXfYfpbpN9obDmCsNaoFvTpmStU6ccQ
D+0e2dEKrONalgd3ipHbas2BmBIC5U0xgpOCUSTu/rbfLkk+bErxD9d4VqUy
QVTNK5hXvLltjRxcbXTESIOF95v73inG0HAZa4EsKU/vxtdLZ2bEWYUbTyQL
VZZBVR4ZZaChAtdMzPC32tbezdKuT1FkzANSyVPPP4OetbSCRLM6+WVRvVlo
MUX/YFKZP2n0csReGnM3dOxhtcSBS66F4wvs0tubl0SUR3ym22jM2TCJZNLO
buEkrUQeOLqbgi04KZ6cLqUys0m82634Eg3l+Rj+KwzN5SerfA50/222/yZm
EQmTEzDGg+649+Ro8onPcMxca3L1efT/H0RJECYVDdmrhPdV/ornj9qp2Sr4
ysxLOv+2x+6OqOtI8i67ZA4zePoAxJne07U+EvLXrQbqF+kJn9biJK6YjUad
DI5Ub0PfP4tEVnLySC9dDVYfa7PS3TAS/6JZv/niQPkp7E7exUeTNn/CULbE
pbhukdO9u0F9FnIeuNSIeEGbuHwHXBAeTbbL7wj1MSoH8XdpBw0aHBzMAt0d
wCh+g/999j1qz/7ddJMXvRJk43QdGfHoCDa2xe7vUUgNV58bfrDmbaUe1Uwu
7dqj1EbNkGV+UM3lmJ5m0dfKjVshu+h7bDstUtZhBgO0LSat5MhVjlC2Nmyq
5m77qkSDU4LQeuoNm3Mn9Yt9YjMcjESfYg4c/UHpnF3XCbgLAychmnooImF1
vKtQIrCeR8VE1lo5y3cb7UlgnMiAqcnAhWbvNcXHggReIp/eWpNqG3szvpbP
ZWluufMA7xeiuBBrxTAIli1R2NjAnPsI7B3PT6v9qYd0BbcvQ5Pg3lj6qJRu
cJCjhNmllyxJcmnBjj/fGw2pSoEtQtIj4QJk/gU9v9wb/lQlPyrvFCpofDbH
al0YaZlx1NO31VGAsgktyetaSb+T+YN8FWph9ekV0tiK5n3BEo0+nunEB0yB
WNqy6noOsicCuZC+X4kP3TCkPAGQljCfDsiiUD754oNxVlA+2pR2Ie0Z7cV/
OlWL/BeMtNSZyYXeFEBk/TWdZgN0RzLZIJTChd+G7rJRZptmFfIXYXjsN1kU
jRVpN8exvyGCZxBb4v0NoBQWm8H7Gt8ns7dtNfu1E4oLgdIfdmxUBlcb/7Fb
IoJEOEPJru6MwbflrfyBwDsy1NT5DTkHVLojHOPCDaGcCNW8VUF/+omyQMlX
V+L+26VrxgrYo9p0NCohNs0MBZCz5JyDcrVQjUbcGxTd5IvDH3NgWnzwGMNV
Xd0LW/Rv8oc0a+Hc7jmV9jiGFfzzEFmM6Ype992kfwflrUKBZ4Tmwms38QPa
iS7yGc9T3PFpnABAjw46d9P2jY+aXdQn+0ISp9sUmE/dz0UyQKlrVR9FCed+
7B5N8T4aqLV/l0xW7szVSy5djt3JMXpYk8rWDaTymvWmOGqBSKHD+hsgOGya
LvygvwYnLiS/Ow567+tBQF0NTIFP3Q6ov4A7hXcaDLpfKnxzhPumBdoIcDej
BqT1vN0xsrozzLIVIwGefg2N4Ot1LDPLcHoAQKDzWrIxvKpfZeItWY3dNxYr
f99u9KC2tNTPrfH64IhoHcoAYyYcotHW/2oEuXcEz8WQkTMKsBFpvNekcCOb
7J0GUHscmtAO3/MVC8x/3qSgSkKCOlv01vaVl3cW0cY41IZ942wFE88dBZqA
nNpauT9f37o2qTdYh5FokiFbT3wbSjx5atNZ2efgJ3hgXsOrav8wyXoiCEKb
w2YznfremCG3hhHhJMpiH8jYruH45pU4xW2jbU3zz0/6rBtpddjjvSUYws4n
87IdV9lNKl/gbdqH+Pgoilr3+Fd/MY6TxZqVYwUHF94QbSDN7wK1ON9BHjts
gPnTlcZiKvCS9t3v4x+rt73thGz1Y+6f8fvl/S4GF/q7txG1Y9t0P9MJ87P1
Bs7KQpJge7ohj+IKbvc2mPyAx8WouVXddDqwBMfFJeR7H/Nds/CSxMYT38mP
2Yd9jhyKNBrMdPf7N8oVF85iQ8/LfRRw+RgAZtARfa+35Rx5zlbT57XFe572
MPvwd4/DPZwoBQLDIqE0TXyJs1u3D7QSG2QgZx4tgT1tbWDCj6P4+GWwwKRK
vdbnpKaLBJEtOn8bmN8XzTxmi8urP4mmVgQQrzgUJzT3nF3JnY/3ZQ8vV3wW
650i6KwCv6WRYtgyK2WUP0eSuN1IB/gO1C1teQpD7o2vR1TDBtbZtvbGmjCg
7QxHmrr3Eb2OlaasMeT0gIjOWlfGlNGpWkChIH0/imoW5oYXTtGVeSYMp5Is
r1kuGQQYoBnuNBPqSe6TnGSe0t9RXnYiuV/4xIWXIg3hb1zIBBgcat3dUaVQ
e500hMuLQBnPbJCUp6unkxfuX4KFDutTvskyKjmWfOFZBscKsYgS6+NZAa+X
z+kkzwm1Y4pMoWZe9y+62CTRYAKkWa2AFpNp9RSw4+/lKe3xlWzOJHLt+oiU
gJysa9URUtNcHFpz/Aha563LJPpz1KJ9bbncRbA1CeogLk4FbRFZQIzvxbYS
Q+90I1qlppG9vPz1ROUspduaeBse5y0OHbE4aS1kkJCP4Vtxjh1B/PQX199d
vEZjTvsMEtdlnj+d7pmcnNuzWSC0Bx2OymYD6zTH7Q0Gdc6TR6gN09Nb63rS
usxhaw9141hMu+ibhnauR1sMCA7nOO2ghUzvezvGyMDsbTyom4Ut5/EYG2AC
2z2ktLG9pHAUYG5ZJp+OKpZ93ciC3wTmaiFkockkMa5LHakC7PKthYTi7WhO
8o5w1gmMAtnuTsduqWoE2ZUS0V6XAW98X+mbLDHRKWPtxp1dcmSFYIrvMQkx
AlmDbrUZMZ3a+2i+ccixTOaxDf7W3coeUjZanNcDY6ikf2g0uNwKjoFXFYw2
iuKM0j+38ExiauaNPLD40d4ov02EtUbiaOCKtTgo8EPZuer7twjF4kcwGcEC
oX9nPoZ8kq9zVpAHaJSYGItg4ZldHqrvNvMwrZpedb/Hhoi3T2ZscxIDyVpc
8+50pjfeCOFQBMVwe3xBYacvwErUaMviM6ESh6fzIcT3YCUgDiiUYj8CF+tw
1kIdMganCsFYmYM4qk352nsAeg8GC8g1+Rda7Y23nLLVoZSoSSuqB6fuNaOD
yAa/JMuYZrSlZMRwtPwI/Yihxj+1GQyi7uVdKOnFiXoXxPdXgowgOvJMXr2X
9IkPtCUAjqxS5zr5/i824WQn0m/9pPVlzsBJ4lU5q+vUHE9nEPxZL5hhvDws
xfsUR1dgCFDjiTFOzdSmPntDxPDbHz/cIzohsmn92jCnP8g6VlxTKeI8afdD
z4XnXMRSkq64DlXcA4edqTpXR7ZViBMbIyipzqlqFKgUEPs48c7jdQPh50BB
fdJ3lu/b7ebskcrX3UtRkLD9EKzury+97lf0cmdBXxtF+/CXhNR1piFf0msO
thdaJo+qf9J1KfAf3z1zRKe3v/qHTmerl4VlK4EcSSqh+pZknue5CeZLftAk
wpVDlCOjfUKVnYlRPPPb2ufq8Ryc62CqEd2VmRK6MGI7f2yi7J7C2z/1vTks
i1AGqG1Jb2H6/RFhTOGElyW3nnd0+G0q2fj+z2Kv9nkI7IK3WuBsXoYnnDpO
bQ7tWIY8ce9dIll/0/atlcWfC/jyVEwvphiS3pJBu+kWYMx7sYicmfyuqwtP
ddKlCW+uWmq37D/hfbQ7CwqNQqRccbUrnbJaXH+fClGq4J5PkfaIAHCBUZPj
0AThF4dTN8qAVSuyFANj0+kJvog4thuGoqKOkfZW8+/VCvlou0uqpPouFOvM
6ne3aorIN6NpMDmwcS1+abYXgp/ceUqa21bpJMXZsxYfA/t3bJF5qXIufS9K
82TK4QMRnZlPQGRN7Ng0J5QoXg6+Wx3jElpOhzk6BNrG4btsIg2ummGNEpL2
L3UsqAzl6DMmQDkk69Icl4gt5iHLWAU5vFySrN9LoAlkg+bxc/5owcZRRKBp
XZVpN94hr5nMBTReReSRa6riVxsLOVaCBPfdoAGB3qvX+dT/sASNyKy0CjIo
Ya1ywn8c+ekGqJ7smhMXwOnFVLkv93ez7BUDL7xVt0wDxaYgMhIvCyt2fVKV
bs7NJYxF1F3rBSrpFDLu+poYjTWCEIctZ+oty48TNOQRe6YWm/CWBV22zOjc
M5/l6vzoOgeOR4+fm6CbfrPZDi43XapRSAccWmoJk8RLwAhxLFSELeMp8EbY
maLtyJNQODKrB5bax+Ikzr12fppo7x/o5qB633gWHKAMAjpFHTCbeD1eiIAW
f5JCEJNXJ99Pc+ScG62X24WKF4JT9YM/sVGHJ8FJvNrFgyX4k3dNZenW+6IH
CnvJfw1eRZgWd8x5yRj7LIywvKk/Gc5b6dyQdPVujhpM9ucPOomL4ho79yXA
B1E4gUo4ZB6ZXOhO/4i04f4Ni9Kn7dodl3DqgGTjm8fyb8MlhF6TCLojPCtk
jb7WBcMb/xGO0Miu8kKe7HaAdaI4iCUpm/1EEpPI3nSOi3s70KRLMlddk6gE
c9QaGtee6rJBoHzbV3AfmCxJNuv1L4eUBhVhyjO+Hr/VnUZHXKJRDio+4gDZ
0Ru4/cxsyq1VD5yq3M+uCjSz6B5u53rlUJ3kHn/ITOJiVjmV8rN6NEJkTO2O
8dGqXH54W1UHexA+MTQm7Lz3kkkdFqAQjcWWsLsR42WiixVl24gjAI8Vy4FU
BD0+h59VOMPiKdkoaUp2kriCB+cMQHINgbpKss+DKXcqOHLnWZNV7ODVk3r8
hwC/yZrgMeshaurGZl13C/Tr/6YC50Rz6ENkJ21mF7krfT4nCAHVpPxZfHJO
J4A1tnD9K5HjaCkFAe4aeG74sDspStUMCQqoIpND/sRNqG0MspbFLas87kRt
5rnS9+JiH6rGHucbIZUVCNd+gZYnUEuNXXE8QPkori3CNvHdAuPDKXNltxfe
b9+ddHFT9h+C94x4fjmwYmpWegyX8gOmR6xwKCZ+mVoBPLp7DjYZU7iEIbvP
cCqupr4SHuJehgXLZRvzwZ3MBz+FNsA+/nI9T7jMviOA8ZTxx3b7JOc59aZf
JoRGV72DXOYNixyj+6sAU4hZlujIXHHCcW/gTjzcZNyWnBQOxJdPfXGBIsVh
Y85ytvXDwAsCsxor/T/K41Fh9u3/aPz2rIBeo41GGrSAUCLSrpU67WTr3vfm
4g0Sy7PuD8Kp6sEFXy3ygybtg/k6x8biaSslpp8dSi3x9PdiEOz4JlKLQ3OB
jWkZmBxDV96TI9cTiXAQjm0jekAunq6pnuPcE8/b/Y6ZAAcORSdkWim0pwPs
NBgiD2RO+w5MPoJ8PpSlBFkBOiueHIJy5xoytqiZnTbJ1RomRHPvEQsHJAfK
4XRyWvI6ouhCCwyUjCD4S4jPi26ezo2GE3KANL+2Jmrt72Ns8kTKdeCpRSUz
IBJxhuvJ/kymnqXSbJwbeF8Mz4XBLQcgS3J0EQyazmegyzUpbo1NHf8Qh26C
L/UHxtuyxSnXPOoBijd4wDYX1rKHh5oCh3TjazaP2QK5u7fxzmYZe6QSwGAC
vw2P9Z64aqRsfTe3jL1d3C9hHAGZjsPUoFdJe6wWUOGHAJRXxLFXOsW8fCiI
pV/ejWJCsM1pLiqMNMM0HfmNrEXftxImMxo7mjrRIwrSbByVW6BXG+rWsYU5
pRMo++iYgnUzSbO/xmCKwPldq9B36e9qKHFYOAYpsoKDHoGgRSyx5lA59IOZ
xbtP5sz6Zu9Qw/KoqOjInTzDtn20fKeZnBKzUf4dlWPPuSv2F7D9s5xPrY6q
gS26lank1me9SYpcCdl3ebSAqk+RWNWCqc0F7nLKxVcqPciR73E7ig07KzVh
JOz4uFrLtUHp0EHQfVUXkV/ueCtBxUw8DE/yLLKNqW9nEJJMFIdoSb7AxpLu
V+hgQc8zDA2uUBad//7q1FxAFqTEoaeKi714Ck1b19vbjeVHar/SO7HyviKe
hVCNAFwBqG4FTeTpeSeorRFatmyVzPIKmpWV0tlin1bOIzYPTx09tZh/jlla
2iDcCrCrGLjZ0SmjmEmPQm5lI7sjiroQQZ4B8+eCVM+Xc6D+8jgTZdFn4yOj
1tFODW2DkBYW4lrybZmM+NSzmkVkFtzurzlexCpnkAP3sOIVoEbtR3ESFClh
BAPuDmWd3VcToV8vF2sGg+q/0lj3O/VE5jYp6LSXsmYjYn50B6KSjA7SF7qG
qpzSOL6J/B/y4BUscoBd1igjSb5y74GQ9kok7l0jg1fQMJV1HrCQWPuwAy7Y
K0cczxHPUO//6ITNg1xCo2HJ3iEkNbEF1bdofNpE2Y1lssCvWnmVz+GfOTwX
igTZOFvDXISXYCWTXMo2/YELhk21XOAXb3XsnAout4ii3HSPTaRAkU+2GBq4
QdXNgO8Md6losZuO2b5ohi8ACTmu24e+/ijxHYzeS1JPL6476COj8wc0X+KK
qoLGeN7IfafAHPbXQSINkXXQ5zz16eVX+z/dGk99bdtYDoJnzs8ZP5Pxyl8D
NCMMhoIYrwVprEFMyg7yhx8H30brFqP2yL4vI9K4bMXrzIfuaMK6TB4L5XK+
sYR204V4ZdLD+1ihqOwoaaNkbxIyKI8wHtDuZWz8BZlLbrIKKeqlEcpXV1hW
AQtwXTruDm+me9iWuzcK9WS64y9r49oCCZ0SCjPqcKA3CLbKELfSSQBoUwue
Zx/nfBkC7OA8uWqEFh+rxRzbAkM5G1KFUTgn7yygAN3AfO+C/kJzkGVWi9U7
EsRj5p37QmnCS1hChoiDKef4gyaM67WH01SX5t+DDedyxvGxY9VzkrqIKCDS
g/ihXhPIiYpJStPfiDta6I8o70TJHLWEcN2YwYQlf3ZLgUVTNkYdft/bmp+7
yaSwVgH7SCuDYRsrfNY4FssKJC+IhYjpZHc2un5x6ljIKWmM3CZxQEHzSDxh
yaE+q47//LMfMKfAj3uZTcZM46IHANxdIb6Er8k43Pn1xDGxzNd5eyN5pMkX
KCfokS7bM6ZvngyxQbXcifIn7xvSx0vg7MXMtY1hbonJA1x1WdOS96j2fGeg
DL5FpyuAkMYuxn1WoCvPzA5xv57BXNs0lSzYTek41/AlkjKeUi6cOwzdIn1G
zeLuHPeg5Et+3o1VteY2XL7bc6Kgv5FDoic0WfQJqH868L2VtXgmrMNEUJmv
qtL1olt5Y1Xj+3hBINpjEET8M7EF5iOvs35n2aT6d9yxLcMjp8O8ZDr7fr34
sFmipm15hfIOuFzLD9hSjWWJgzSrtwW6Q22c1ErOkxU6ESnWTRJAqdbXdoaF
EEUZSg0RywRrEfiZsnIVTVi1ZA/3lwUiZFdz43oz4POZblyV102ioUxjk1+0
k/7TyzyUL7qhoMwr+vk8ilXOZIRzcy3X8tdz6Tzyr2xRyVVQrD7SFUKPhQyS
QNZAiD+M7Zqp3Cd4DHQkyjnGsmCun6vPjX02RZaedU8MSDKChTtpdp+j6Qg3
mLOZ8V3NLOPXVFqB+ALT/gFXP8N9GTYgQ2vinbpHH6YlanZEn2PfmlhIk2hi
iREGMvkiDb1xelCDk8d2RC67an7ZWZTjvNAqjYlXZurL01t+SBTJ+sQObW+S
Nnh4BT3nyRj6HyK7vm1+CbcLABg0CT44aDBKPxyaL0ZjRWHS3KJxdNQcMNQ+
nqGcgMwvk+OgnRvQd+p60VOAbyvglVsLtD2Wv0EzVOoTKv0cAI+gCA2ozLU7
ddbIDKyGAnFU/U+bscIUQvUjMtHKcblydY9SForIV06j0EuMHLWxMOidMvRz
GOaYL5pXo+g25V3VO2gaefO3RgP6NMfjBuYCnpIJcbAg4YnQ6K0vxeKOoN8M
EufnF8E/D2YMJYLNVcKZ/yfw3n1CTnFgDnedTDyejjMw7DMUY2bCyW/Igjf5
lkEDqbSohH4OQb2DW+xdgfzlR5TOXxjJX9d64IwGX4qVoApl18sPrYPVZ2yO
yPAMMGaRtzdQMM9F1qKKlzpau8Qdtk1UaebTo08948lG3L9jBp+35dT+ajGY
LdrBXnqqU8bzjwVogNsVTD1nYpquZ4+XFx0ADBPJUbfa9zC45RKfe6bp20K+
aScy2zJgnDzUi5c0j2sT2q8RciCk1voRjL7yB7ZK5U7PESOsYkbPOnqw8H1+
H/S2qj/nq8vPCnwUrDuCGhAPD+2Zct9XQiiC8DM3Seda5LDEzWJnGVg/ICPt
1LykXCeFC4/KEKGxsCMsB6EHBofst69nFCZBimJVVaToiOOsjOdamjwbuu0X
DO4CILvkhhWueN6nor8E4BMZ2/NNpRskhekjYNHE3RsEUsq7x1Pzss0huhDn
vaoFirtMjVP6/TXdDc2vfjGgGOlYBeEsfGT7mD8nz32Q+zkNtZFcn3UrgjKM
a9X4q95q/Ro0ZRSffWRdeBPuMMRSW60vtmcVHq9Fk4hx3JqNr5QSqRQsduSa
AUUcvkhOqsNM3ysACifwByMn/FFZVezJtdspVy9kQDUNV48ItmDEyRRXsHpi
9OMpYHIG54XertRIbvKsC/r1R0KLW8yIiJVszF5IeLchYN3AqnbJCmXJkTqb
rxttG8lS633w44HoCchuoVcVr2iYyfk5fRCabzD5oDy6r3a+9gmUOb5pmJjZ
qpiWynDn4JCTmEruszO/8u3ekT6/rOnDk3rfe6lPZEG5MVlLYswjDB2IcP97
0zpJNa6LFBqMMdZJk6tyGN/sjQfNbbC7R6RiEBfJbi7DWl0jWb03JX1p8muT
R19hdOuOARNoFaqmNqB69egvzk2XvGpb/+VhNAwWKJTZoo3OjSIkZvQcqgyu
ZSHMmVuB55wyL77E1U+gMDg5KZk9T6e0EnLA6nLzrAiwGpJojcLSZEPztSK3
D5vJwvv/tkQ8j3Cc7sq/PsnyGZ0y8lrAwfJYr0nendrAPeJofsLgg8EslD/P
CWL2tT60xsy5wF9iCxzlCaRCcjRQxpz5+ZZ3Tsmrn8FLZlhIhEO8OQAdJUMI
FeBTcs3nzzv0b/Z0NRLhBcLaCyyYEH2oj9QDQXSLP4MVv/LNEoMp4J+YwhmF
l9wGg4DH07GvemEsiI9J/v6T29LAPlez9vQel0LUGVULxe9WMSvbIGmm4wOH
oLzF4J7scLaI2Tb6GnSRgFmn1a6aeOlcx17M0qE/HB63NaAbSjR+/BKEA5TY
dPbr6Af6JkaDl3DKzD1FocsEnB8ff2Hrekpw8OR2ZcaEW8FJB2lOAgas7cwo
OGVvtDSBLPenq1C5knEIdrL6G3UX1EqHfKAXnig7MIWdVtAZjp9mfb0Ha7gU
FY0RMAoJAH3IwlISPQjA63ycFjTMXLzcOivcPVgYv2X4+xC3p49i8VqX3Vqj
ZJHW5xWx8NZ+2gmY6h0uAxDhGJApz+UUAO9uXwgwMLcZN1Qw+fg7+e+vArOT
iQFuz51dGS06z4QLrik0Oh97hSzPpNMlIxiXpedLeUszCStoumzTvkURyZya
xx1+xpS7RN0mX7zpgJSBMxfHR5zF0DAZ1mvCyipCueYxsFPsWpKEPcz+QPW1
xwlNVCo6AhObTF8X26g5BBcniLWHGQvyE6LEUuZKW2xJe5w3Io1Qglqh2g+o
W8m3DiKc56eV8JKJr+6YnKJmAcE3NBJjNJTEu2PzoXIZxoSOo1ALUuNtffoJ
TjrDJqItRcPq7MQIQZKqfvH6k2ejlbS3zdK/1HFTg9DCLNfsN+54nQZimdPa
FXPx+eKLG2pK/Zh3sXUa6QdXpunFIisIICmYbq3ywuOVFWbKbzK6BvP4gOqu
L05/jnadVIkY35XEuYiAi4RSd+eGb+oU5sD5SwF3dU51uQe5rigXjTaSH9F9
QH1DrO/HHLB3J/9E3p8ZCoe8TNCEpVIxJxMLHJoN0PMAhgxr5QrcRJDqlFnY
nj8tiiqbCESCZTOENd6yrPIc0Sr0uQDh71tS/2LUn/CyI5dFTNkz3Nls/+V4
nAGWLCPFX8EglEbNmFY74h5494+opJrtvNWXOTGchP0hwEYUcAK5z+HeEna4
hTEiw/rKBNoUUwSOz/RKIWBlSDcDymtZeqPOCXJszNefACxt/wzyE8jskprr
2pNCq2j422aahEKYexARjOUyIwo3hLqV683LvQ9kc/3vyR7+6XSRW2pu8frs
wBHTSRY/r9LzvfZbE5vpEsHjPyZ+UdJlzotD3q08GtwJStkJlx1nSqn+Snym
slAEB5FmG+82WmjTldugneegrGXDGklu/ClCGMLZkDDDCPv7s2S+1I74ieLb
fr7z/eqFAA7A5pyWVZfawxhpOFbDcx0AQX/QxHHu/YDIsXChNZAJhigqcgrT
ezLOD6rv5d4MtFr6BtFD07nksbSzg6hWfDLAoFS9c4bAgFX1vQoLkR+0CgJC
6k2T1u9dvSQxvf/Ua+RnksaunWiJ9nLhxxIWb0GWud2PnVBYXxYxVEL3exw1
bCJWPCMlI6GqfTKWpUabaq4Se3CinKfSy7khVONOwAzTEkhXddS7A5/x4CYV
O8jqF9IvkYYFn1JHMhWWUF4V6276RyKrPGQ/9JmGpCT4urwuRt/25ZPXYg6k
dYgSVRlMEVLd71KN/nAvxuRnkkXPJNJIB8HC1rwgQJMEReAM/+jMxbN9Jy7x
1dTexn4EWBffUFi/llmO+mQGJarEFAuZN+InKSZP577v/kMUAnbuXnaa0nie
8J9e4ZncsapB00uVLPw1b2Vb8gZlvbc4udm5TaggDTPV7AlEBztCxSlFRbHA
xM6aUDBPZCSSk3RB1gcTGzzalA5E1y0i6Vf9gEw3gELH5RDbLnmghPWavpkD
ry1g1RjWKUL3CXckoK1YCi+8xsSNZHZvCWi/j3/aEgwX4QmDiLwOUO2FeOtJ
IVjDMIw9NfHDSBIHc4Nw7NqimlBcEN2AfNIL81uafkORt7NBAHz4xYyX9LNe
XNOY8IlAweN7ZLWeXUihg7exbAYE0ssF2OOGcpu4p0eghZP9fFHdRT1vr0j1
OREScQZk5F+fc35tHWLRPp89GVOACH9f8XNJPxaun9G1yNS4bNRCFWgp7gJV
20ynPFiCktsvl3ErGq0l3yb8Aw5VddDeYaP3LFaZOyCKhMiMVRDeWnnN+evF
FGvT0/ykX1nax8XiP7NanI8OXFfv+Qk/1GtDheG+sHPwD8KhscjJWjTgpgqd
kJ9x+XKoCnvbpz8iWjLh6XBViMWilbHOtCk15Y7E0c7z/XSHIWJ9KCudR1ch
+GPhIOef6VJu/bRnmiJTqsVHZlkAs7WzoDINmRTy/OPGcFaYWcTms9VjFG+2
bqpnbLutHwOT4Z6EXiozKMWN8fU8GOqsBFsSgSwQvcW67fuNEMPaAEM+z+uU
6KauyIz7x8derJhTsFmbns2s3u02n99D2lD5muJXXVzvnUhv0xx7MgnyyF0a
g36DNj38gSWzZ2D7x5Kyl1hcGPL8Eo7QKYHRND6xbHaEaf/z345uiBUKclfZ
RZZH6MzAuhC3jUZnfoTKfWgpVHWWzfbvJCM6bJI69Z4v0adiEqsxJzWI0b0v
TXwbxUfos5UCjfrjDJ6uZeUfaUpn8folCTM0EL3dFSaGq4p+NrKOQqaTTQHs
5XCbnejZydrmFX/+V6jTCHviUzEkFMYzU6jmQrhbmDmfP5wAb+y4v8qZPTfU
9D6sBHm6UYXZPFXoBYYBkqi+mu5wA+DE9iE6MK6UC6YPf68N4TaiMApq3AWe
2o2fuRKoX6to+uD3B5+IBcTcYGbDgOl2V0xZp+ztuqvWghbRL/GYN2lX00sG
J5asz/uqBB3Nl6cpOmM00ZUAaWkQroU41f3ejAG6uqnKDwkYbzmkA6c/hyvz
XLON3o5XOMJF3L1XRUq9SCVeUYCqwqGnTyvdY8PfZ3S7dmKkzmnFPWDBLO/o
tUbxavuYDOTsRVL5e3IwKcrUDSvcLnvseyAieJS+EWn335aTtw7ASbCI9zVY
7GVo4UCRsdaCd8mN/uSL6JTwZT70YBp6kLwBTMRi0ZEABg8uDZcsQJQoonRU
2PPqYSJULD7GPGKbRWPkRBnzsgpAN08fZziuxJRUK8B8fomAOdtsq9jZoevZ
xEaQRDkEvHSNFlp58e2kEfsqm6Y2O4qLigDmAT9ZiIeoB9hfAiwa7JFcQhz1
QM4yyrPol/KmlJhkm2hLDALyyKIWI6lYh5S1v+UhnMpgoif7YiIlYkiJJwSf
7WjzOILSF2mqb0ow9Ar18gnsI6o7msHs/fgYDXbREEeSOmpu73cFoTnwGq3P
/csSYOCKsJbNuHixw2HnMQU7cI998u/h/LXjJuApa18kuTTyItq9lROscnsz
rkWtYbiJh8or4bjwVB6NVKgAIcXjeFZOXrxAW2Vhb+SXv4yqeiTtegLmjT+a
cvYWqcBpCKwZb1dPXGSPul8YyMXLPoshgL1uxcluyBnGmKaTN9Lekqyuxw+8
XOHQpgrEnNo4DBqQMKfkU/dW05DzYeqKjvZiipkw1dA+GJYYpSJjdubO5rHT
Z5UQfX5W4jVHO6XcufL1sZvbnpz4uxX1shUxluZtA7i60nS4WeMsqj10BmMT
v7Z/5GoN5GsHLryEqSWxqL6jppt5oRn2d7M9rUBamaFnnSIHzqRyO1b1xCgP
3dy+WO0ZPsbA0l4EtfeaXdSk3Y+ea7p0n4R34/XOhq3uqDt5Jyb7eYp53S62
jDTKZjRBEgpHmJTzVmI758x9YzgmGGgoFjD2ADkOnePZGNIOf2TLphks28GO
8KWcXiIxclKYYYnSj0wx8PYEsWw9OPoq8ZJCXNqRBGWIH0PU1S5RJKYbqRcz
olsZ7geupYLSmLKjgtqM2/DwSUccaOVFdwZMCEHPYuyweF/0WwOSf6JTAK1E
r7AYzHtN4xPM86LUjFTNke5SxdR64rZLxhvs0a+cp9KUap7jLBzXcYIr5pK4
2bwnHeipV7CfjAdZ3r6ilBJ+z9w0p19pJwB3YXHAb8vp+O75D0CBdEcl1DRf
nsu9y+PBEe6g2fodj+A6YXKPEgX90UjuoQnd/+pVoI9SGaXNnnspuWFbKISD
EitsTE1evZLs9iyLhKpzEI2puXfRc23M95HcLxAO8wazJF5AWM5Fv7LO5NFN
AH71jq+W3gJQJpn5+HsEp2VE+uPsHtfM7ook+T3yWQtgdRZr1BFp2RqKw9c8
8p8PV21THtoVW+dAOOcmeOSbx7llNk0MbdSCt7cDEAzUz54QRxWlTo/TOyt/
xDQAaqJIXH0uipxfuA5KuenHqdbCDoJCylP56WW73w+QY3kJsi9Xc1+TDzZA
pVlef3QuHOyqMIMmEWeEq9HoGFfe8mHCxAnHnv9SJfxESXMqWlo6QGmvYwG9
eL5SXTbx/rxHoFj4T/KR2KXO1P0+pigoyXbF19ukLVNl0tl5/cfFOcZjywGl
rPXjQZhqiOzpkVWNtr96u/XJbLnOAZO1UW2XKY5vJNuBHC5wSyxJiy19WeEv
fVF4g2pG9/P8l1KUlJTzkJ6/kUijGXMKDvvLuvl7b2T6OmeKkvrDyIDQexEZ
wz3Gw4rEuLGh78FOHvnMEaWmE4rRb51Ib+prW84grzjVlvO6dOx6HrrKta3C
OvdF1pdwO9IlFgOQzilvTSOYGwLY5/yZX81ixYgPAqmzNU1bdCZ3APZGaICL
SSMIhA5n2/lQX27+NFpkTvKpKquiukVvzxgOeDGcRB6FuWw4rvi6xBey1ml4
z1WAqbgRjQ6mznpcqaCawZs15W4eie8xWPEt1/4/p+EMiPFmd6wTWLynnbED
/mLFEIrSba+d82MGfYRFLkvpFrw12IySQ2gwunHQtD9SVLzSmHXDBtFQXzVD
fpVQgZ744Vmo0neYrimOXM1cd/3RGZLW2CrUtY9NK1xO2IPMonpCBBTvWRMW
MRGFIa9GsdBh5HpwYihaK99F0CPRG/PXfnPljv3n3tTD5gWl8s6R0RuhwF7D
CGDGJ+9YAbB2LzAvd0XmX2zVUKlam3+U4DTbgEqKCoZVJ4naoO0tiUbmOCkL
FnIctp2HSKJZgpQehW0c56uHNaqj+HHQ91RaH7lc5R+gLqlloBdJ3hp3TKOa
SCKT5Xmy2WKo+pfbQ/ahgoYoYWdr2DRAAhlWwTPxFU73GAZU8VFEo0zpSZOe
tC8Lddz1WUCGfCNKpHVrsF7jY3J1yUz0lW/mgUqD4Jz3ZgDcEvChD9swezrx
8M8acUfi5zPVVD/ME5BxSVTTPNMLzkysh/GfzlLClWt7S7xgQcO4mB8vwbwx
6DqZwOWhtLMSWvqlzIHMoLAqmDHiueL0H9AgYhuO0WOuLjD6XXoNcfw6YAyB
BKHImGDLcXPTzvgiEiiWiw7VwX+10nt8LWanmMaWGvjwr+JKWlJiozAfgse/
odb4gksSWDJIfkreJ0/Jh3kJc5i584RENI09W6YCuqilXsvM8Jh1vgs9U1mN
fVZ570dBhJYLIZbbU9lwyayt0gHTtA5A4gGXA7WGMdsUeIEBM8/ohmPpMCWz
hfpiBSwlikQL+e0pfvBYckDC5fLMPNM05LrzQ637qaR2b2nZmXorfCZPMYWj
mcZegPvJiw5a9CMsn7MfcD6VEsx4V4VFSn7+XjDb4Qwxt4u7vfyD5Xu22JQa
Ow13/C6mCqsTN6aIQivG1b8nBY5z/B96SCfNu5xQTlCC2s4h1cCTvnmGMqXK
Dg/b/31yZL+JzBo+CcXjslXp1ZjbQO5XvESxiUsLphieZepwRR/qCcZnxCxx
vuHWE/7DCK27Tt/L651FgqzeoHYZCs3tf8p0ao6ppE0EDQDvlcYSwWXVK192
6+AZTaHYx6E7rne9LdZ+7m93sKC6H1gPIPZ15JjRakK3dpHzyYcFpQNoOn9c
PFtNvRI3WtF59f6FkV8Y3ZJSv6GTYXXXBATxADyvUejq/N2S9KFfjQsabLl6
QHEqJcxfDtDxshV9z3sJW3FGlqheEW8GB7wJzDZuHnfBXT0KvC/BCfUg1hPU
lon9THpAq3HQlT0uWP6/cB7E3OjvKVmvPQAUZodppVzUrd7KVCXjF3xvk9ki
oMOSQBZTpZETP+equEVroFTOlLS2OmzdIh4viYlMuMn49FEGjF/3c+CiMzBU
yatKdNz+h9mQGnw93pQW2UId+WLuwuakuHsh8xlDtx/MxyCTH/6CEzK8X9pR
SUeONrhvWv+PbM1O0w/Sqp97PnY1xGrba0WmvhbrsOz9i4Z79RgKDucJLCpl
5e2VQp/llezMcAwE1tcCMQUstmhYq7RXcgIbbZ1heu5pMyMyXX8VZVw4TJB+
efVX2e5LC75ckOj0UYo5Q537AJWg9pvxrXFuxrGW/HG2ca6PZUGoS6faloWk
iE9H/VGqaFRG/diNdpcN5sBLLtpjN8c4S82hu3FDJlCwTsGLGfkjJVdkt5VN
y4RCdFPyPuyHNPWIayay4KXC2DdIbsoKz0c06OxRWCX7xL0KUS+6teRRxg4C
Me7KewYL0AIafp3r0qv4oc3+bVeFswdAnY69RZseHHT4+j3BeOpnmgn7fYP6
kwiwFDj2+yE3zbn02LuEAixD2zEaQRxAUoIG4F6Y5Pl310xtnvm+cny+UM8r
hyUQZz5stEP6IIKulrS69l93S1R2tv5ddAhkAHpRYGJyA0Xb9L9LQ/ugWjDW
uZlA3t6BVk48ZGXFgIJW1vsks6/g9fWn+oyLLgfea05QjGUpqjMi5E1knz1G
5T7KLZK58WI8iD+7bwTITOO4v4zHUINzrIDqX5UOj5SDKqooT5TVuf2A+S4n
EZhoaWzTTwMBepCRgi99t+3XT4YBkcbJexxocHr9zJ1kyM4LaeGU2YEI1fB9
1m8FlTNprnjXj6qgTz7tsIcVTecoUBEsfmG4g001blxq6x0+F/bVGcGdGy6b
hCY52VXSaZEN72IwOspJNjRoyC/xx0itAYrH4b9yIE3PmrdMHiu9O1vNC7Bg
niKArt5JN54VKMiBrFCwN/ioebDI2/JyU0wMYgCDId/msRNOa2OPLQy6rTlM
gTVSbKh7y9itNNUPsuSoD/AuJsOKSSS88bHJnOL2A+vEk2m8M2xB1qG4pJEc
lNWPp/zv9RlSetOGV+Pa9mrh3t6/aKP67+TH4vL9RCmuUDLi6AKnQstC54kw
brRGgpjH3hj8yzmccDABdodihwk65KOPy2pCG8WDYIMutrNH1YlNDQ3ls+Gm
rA8sgStKiycnoxmwro3sbf8Xz+9oqn8H6mIxwAQkSZg5tOuC5owqtEnfcjXZ
qIylgBq7hGdY/jClnhJ8xUfdc0BurKT4dkqpKfEE1Whr36m3p2xc7BZk7Rfs
QXxKaCXRJbBH8vuCOUWKoFjAoPcD6VRC+RWhtdTpgxJpaw2M6kHBn46j9Pbc
gqp+o8I8KsCqKQDNHYi64K+HjjId8laiG+hq0mNJfLFbg9vVtCJokwyFuPh9
+W1LRV/UW73zOcprqHG0Wn/4KKjxUeiMklF58M11Bop6SHO+Awu+67klw63z
q43jEF9DdmTl7A6zN4Tt5M2pGhcv4/nX/rSQBxpFXPWbBRI/CyqOjDcDHlbP
ylYsYnffHMBuTtpwmHCgP4DItPGn6wBN+U9aTxTuQ5V8GfIxd5xqyiBFaFwF
siHxRngIKPuX7GKzTnLwSugemHkZ9RCV8gcumPwf0aalZp8bq3ran6Nr98MF
c68aUYmpmcySVxrKRlYcwPfR2NOhNqcUczRkpG4ljscCq32DA2hCS4+HySJy
BbvyX7LsbOxQbCD84XPDREMpDJpNBZd4GINr8egd8iU7Qu57duSUGutdSPM/
akwMdfYCTE0nIaWBWkGjeM8xrOJLK7SeXyUT++ezduZo6Ufv6+O9Q6aXAaYL
29fRozT0JI2SmZi+YnMJFeYHp6HcsCw1GTNf1mhkPs/+nd4bvVRgai/Ovx1G
Rv6kenav4RHki5buKw+G0c3OjcxyFSbrZgiVRtrDBfA9yJa1P3A5ixlRMxZw
X7zwBlpaBsFjsIunjRir1gvO9mFzUj1jnBeksI8NimeIIpK5UUrp7exs71ag
tirIvqvg9yjH1sdD52h9j4uFy8kJ8IovB3YC5t2LgPxy9ibFzWrFnwV6cJ4A
eYlRUutoYKgp0hN/ZKxjr87ymRIfgApCZXO55/EBni0DDhIq+OND5c3fQAai
N6eulUIofrtTqh2zxEUA/DpGkJCHY1qo1cxoq3Zo44vEicfPcjfhfNC2fj87
3I6QbZaQiaVXc83secT6zZI7Jurky8C7dqsE3sGNSix5TYIzhpF7qokQuJ0b
FpOQ3LMzlAElF71SAVg07KuSnXwV4pocRRNPzR9SgKkIOCLc3O/7aukY4vOA
BRMq51UA2onyM4C5Pl6TG4SZj3vQaPXZHtbqNAGbgV711Ezd4708Hm4r+tbx
8A2eixr99kqZowwlPOM9dJG8OFB8WU9Ozb2pKK9EQXxyi1dLJc6r8DcRPyPB
7ho8MSrZ7CIxEIMvr/2rvAIcryezUhrTBM1tp31zVAmxEJCEoveRNQiVVIGR
BTGyv0LGmVP+xZeS8lUmQOrV3OELpsnCxzxLRqcwzuX+XCweFavGYaJjPkjZ
pVnfwzesrKYjjlVUrK4hq5w6svZO6Y7LDNsj7flVXW0EHR7OWUL1qFnWmicI
6G8YFGajc9+RIVbdVy3usxcKfLRg3llM/LZarlKtZ16UuJ6g/bWecmHp8O0B
jopgLglS618n57iff0hJD5YpNGUec+sVxXSDlsywbKplA1xIjhd1SIxdzxwE
wx7DTBhH/bJEBszEqhSZ+C20k6gqPLoz5I7T5pRS5ng18QBm173OB8EHRsb7
HK1/OP9hVOvcJYKXqEeHyCpa2pbwu9KOwcQB2jEGnOs8WNmTzYGO/Rq3aIe+
Jsqzw1Dx33f/2PWi2mB1y7jvAakbmiUqmruc2b4EZIia61/KXZSTtkYkokP9
xrGq+P9oJdra6rh4IhXmHKsO1oaJHKoASOdLKc/Gf6fUV8kM9QxZ5qKGEccF
NDRcuMSx+wzmUdvR52gc2jU9Bv0ijOCRLtXIAv7uHq5A3Ve3EhD5Ct1HzloS
uhQY/Vc3Upg4hTFleGtO/iSacN5lZlFojhLjTYh8HWegSSdly7DypjZh5f6E
xhaQSkIV/pMI67prmgPtudPGCXo53gaIxxUdODLC8LhXoG2H7bpZfK2OP6xU
l+Hmp8uOoWH6I4g0Ez/gHO9qehbTsxJPzfvzngDA1MeCXabUr9aNiLSQha45
CmKD4mb4TfovMnzKWlDcn0/IG2IF66rIqn+V8Dau6UgW/jwjH0kQlQ3HFwxN
jWgg7dnVxWF3W5NZ7plzjwwdtetsh9r6mYsTta5d9/ANJ9eWH0+Hd2vhXcoh
JCvCu3YMCgrN0sHpLFXpRYjupy4sPTlD+K6pa7nbsy++IQ8wem0t9vSsSliN
v+bExOrZlaZjtIqCDA3hB/hMOlAn4mfvZFMb6EMApV4r4YP3YBXoh3RMg/pO
0ef9COlccAQmHVQ/5APNNscq18v7d3cDFVjLyONyTxl1ymtXMdv8YTrMA0Yv
+0guMCIO1i07pbV5ehW/1N1bwjDoNm99F6CD3aA4QMQg4bbur9/O7WyXYlN2
2H6xn/uFzFNC1SH+D6a0NBkN7vniyEgdTmScVnsMt/+OkVo84RUZgQbUvC1Z
f7WEcp+A4sFP8upc+Fdt1d/4/Vbbwo9EicHMNMD+w0s+XfomN9L/HUkApjD4
VEQTKBomvcxRJ2CkcnAgkX4X9w04xXk2CV6Pm8fQXV/fve2sQnMqA/lWaleY
aFYc0R4ox+AmTMS/1uyIiK4NmRF/k7wtttkJwpOC7rb4r1xA6Bx5OXYsbCz6
BdZtMtjdpA/c+OcJ61vj80n1Vo33o2HIImjZF9+zdSCQAjvW9DtxzpydX1Rl
DyZdmlNtKwuwxTCWJ0W6ojhygj8eY/GzteBBeNH3HZ2T6r0cSulajtf+aWhN
dUtMjeRKpgKDe2jfVl+LEe889sx+BiICTz5WurANk+lNWlMLFglFkFXx+nuQ
4K5zWymPY++XV0nHYnbz+VTTxiOMaWLXqwV/YceiEDGUINA2gjXmaHgRXLvc
8sdwa2/Q519liwqCNGU/TgRQUd4wuwXVxrZrw3vpvCLHzvuXOAhdQshvbINq
4V1p70FcusMtUVV2HuMgBrT71ZplpMAPO9ka+lORnYAnMK72+ZBLwbRbQDOO
9KNleNiy08ALdYS/fVMk7ElqpJVXsZUO2INJFq0fXB/lfdtGmmD2UNpM3fCz
v9dPad6BZuxzBrQ7WtztGE+HfigA3mqaKe4z0q0sK6bUUm+LWe0kbCCIcVRJ
UL/Aoy8YQucR4xlDwSc+CtCRpBGbpkHEzuCkPJY2EMQmw+yOwn0aoV96b6w2
jb9rGvgsQ5/lTezkEcBH+aEzlSicXq4nLQQERQOFuQWddHOapKqDjbUQPma4
o8KUnHxNnnrn8zmPdokWH+s0oKy+Qrp0KzKRrqW++AaxoXMGQg3C9PLIOgvI
PuY26ZIncx8dcCAd063lUhhnsAzfsTUKZTF5IWIIvPj1mbryf1XQhaCq/T1i
t73EOUE8tKNsLkv+jjwUJJIPW4h3EoIClNmMNQFeSOmGvsg4PLG0N5e3zQcS
M8WmM+Fcfl1M+rrkTnaRdgsBYWvfwcJyFGZalgNXiC1JNh+y1g9YIEMSnWvH
6J7BcjVPocgh82ka7/3QAn88FmJski4FLkQPbQn/9RvkwU75i8jMT8ZcMKNV
l2SlW2gt8CK1IIj/46ILe+EI93j47a4IdbirF0jQZ8AC2eOH3NJ7plwy20mO
MesytTtcxcmYbAorw9G7qMr9ZQkDPoq+0Duuu400rQTR13cmN5nsi+6iMmEw
4xI1c3McNdsnwGDWPDN0ZT6z37+AbUA9qDAN6Wg27UtIUwWsrkVVySW+ehEH
ATwi0tgb6XVNH9yLz0ST4v0Cc2FAOSF4TozwhzJpHh/vZtJjBxNZwRSUxhzV
ILis5n2TBi+5+N77v4pVITLKjMQMBfjBufSeseSYW1hv5nLKbP9w/SbXlj9P
wZHTTE7zwUn+aW9+PKEtpX7bVEexYvd3jj3pAsBrubBJ/MLO8KCp4dMxDPIM
yRj8DyPY/vJOeM664dEWFWUut72WVSaSRN9vbnXWg6Zwp9JqXz2L0JH1taaR
dATFknOflzXQFbwpt1GVgmM7rdQ9ygMWfo5jA+chQzl9au7J4a0bRm+QoMyb
sW5YwUlo+CKlwyw5r7jx8CcQS89kpspmLOmXu8qCI97EhmT4q2iKS8mJXomS
bunnQ8zVxMOL4STRZzWc92OYeDrbEkQ5X9T+cIugoesJGKn4UKqPmWj2P+OA
O74BPWQ6v0iZ6cmthpo3g4INt7DmIrCXYYkVO/1x2c1AsQfgGINvZAVwtbgh
mlr90igo0Qz6DUsqic6KOOeEjYnyQ0JChJ6pllZ6LX+aLIPAzPdXolXoJqQ5
1kpw72z7w+1cZFC5aIPMILBHS9ek7KsACoCVQwX9Cpj5u9IAxqZUdXqw5gwu
EQnr9gRXxJUHCOh35TKnFAfKEcSrZuAkrepaba1InbRZarFv0UF9HDNUFjPe
9kB9w6iKDZbnxyCc+MESzx59sDGCHmOGSNNtN08KfYnZze8x0tNJszIi+S1a
Tb4KfQh2PjBGnukA+DfEQPpoeAPuOhzti6kazSObCnNzNV6LhRCSPoseJc5R
YuH47idv6LJSAQ4vVLXZu9+enjZDlW32c77KlID9LtOl5HSfWaEvJpATDJxY
RD3UpzlHPB3j4IoXRH/UxUgeLo6sbyiYCvd/IXRe+OBVTYfQnutjxr67BJAw
sbIO9KsmQ5rG9vJeTVCXf2XuacRjcQHwOkMhN/3k+1FdPcEA89QHBXAgmrpI
NvZo/O8alSaKxqBxEiNE3394MM7VgwtjIBkXyJgHo11vC1dvRvToKgCRlQbH
+5SSD/eFQ0AoQpHRjcbxtgKM6JWqek69ijUAxxv2PtE5lg76ubUS7Hb7rFjY
8CTxterfB45zsD/Q2Q7cs2oBTC0jBSj9y7ERsJPGwj1Pt0CjuAzPwXC0+V6J
31DgkIsNggChRC/F0Xph6KyVdGhoEk8vXASHj665BtSCn/vx4aEv9+NrI7GJ
jgAtC2L1B2kEyGLUIH6sehPwdWyvOI+B8/keKUDKs7nGyX3e+SKXD5pUUJOJ
9wYGrTTkFsd8UuDL8yqnjaTEHrqUCYiNccLr46gZyeNKO1J+RbR1Ykd0p7pw
eO5Dli89d/INnZmMzbWxaHe+wrm9Um/8ugDULbkESjW2FPwt5YoqFJenqymo
Y4xa7IcCJ+WsdRPP69i6/fSvktw9LCl3NgzjCKzupaozQd1dNkEo4MBZm2vY
6NN/OoiOP3XbtVJpIjUhHqvpN/rHEDxWgl1KFMJUaYsxUmpP8VQkAGC5PlLL
+/o7ZzSwzYER/Oe3qSU3GrsR9+TcorAm5Dy3S40J9nuyYtW45pXPLuk2QSmg
w0vAYEhh+UTiRAPwSVfZkO3KRWVmtpexzO214y/dT4/seq2HlCQ9h909QJst
i5yPvsbX6OE4MxBWOGUliQjekTJt3Ht9HmrdmZPbeRFty/AkPlgt588bprMv
1gMiv9DokNE2IzJeevBv9mmZ5tHEnxRTY7XTvAhd7O9TP6mxlchqsG3U/LWr
bNJYpCwVHtN8v0XdQgVw73pEgJC+JhzcDD1ZagRuoLLA36fUWMG6PEGG4Jwu
Dd6+AlFWXhCdBPI58mc0LQRqXwI56t9x5Y8njw0i0WPMwQwrPJCKxaWbloK1
LgTN/mtEQEPlB59jpimJcLK7mFO364+PCvRoakjvex5DnLJsRqW1MLYpTPq6
5uxivdTSl3+EKM0TLBTGvON0J2sAssbLmgXPONXLwL0gIRn7Ca8zRtnN5HjK
u3j8JvjG6yizrHJzN1fYacqs9j5OoGTQL7jsS1cFDbFsBHAIKJ6BGzbTeXLE
WIgaZLGWlWU20+hK8e4iBmoEdBkY6useO6GhPZ5bFws/rMOZduH0TRyIudny
Cx6Ver8US7SfIoXLyUCA+p8TYLy445VCuCNAe813h1Sqs0G7Vx++KhZHpKlC
HyuQpZmu8vG4D4+jcm/Y/f+L6Mb8G953GAzcGMD8EyXSX02IvFOCOk0r7Rpf
tlzixwM1Wk8JB9qeNdEMt7qe8NHVvI/D814URP/4qMQmEjke5DXosZSpZkBi
p6eEDKLH+JShd+lRmN0/RbmIiqcyEMIK82xeijyb/tbXINDS4G1HuinC6bbr
vn89TojZ7wAyzxdAVmRLaN2RIxqMK4qjcFgzFZKBC5qaOy8d1epAHXiUlfUW
CkbcRrnAndPOEH5yHnolfbqDTWICHekjgtTHaun4cKi0vOgwJJ79qculX0FN
ilf9hQ++tWGY3XwNpsYiXSqfVFVqPLGJLIuvEpC5e5KdjIScbCMr7rXbezh6
8Dj0vDYAmzbiYMpUAg7p+n1E+rpTwJnzb4oREj5Qb5ILlbz29uVRvfJptWIT
269l1yFwEjldyENLeZ2eaBtqOvrk/bqWHhRBUjk9OfXGWY6Di0ErmJFIPiBS
JQFYnOAy/H7K2zoez8ZZCzjS6kpcyKm8xA3ihCcpR83INgCqlC/ryNX23QVn
Y6wfd+CuWumG1mYS6GQlWaKBa+8YPC6BENw4Rq6ehUJhXqYSltd7swpxCtYY
zH0wxukmNrK2Y45VvdQSyXP9syFvkjjsbVMaNvPP8pnKn/vHikaN4/6PsqDG
wuYLZynibMhlTSJTCqhfiHGz/yBpZ2kLzhc2f+oC+Koia0huzqo4rvLcR1EO
9lACTmel5+BUsfeWLj7wOD9IrOtQHXcuv07cQ2s81f901rwjadRv1tvNBar/
mN68iiXKnC+1YYYYuDhFiAbb+2289bMn4CyGlXvxE4Fpc63XG8pqbOh1sjnA
FpeXkIPJ3vp0RiXq+ohbuAkVuqffdwYdz6HdKCBpFijw3FeTXcs43WhaWYxG
9bakoGfO1cuqdYZzOJZmYDG1XOQIEv83Bzf7XEo+dCl0U7z1dY5GpS6QVVOv
mbDEcnKYYUqAovftoilqPtYWvfe82WbUKIVzJXpl24XQutJRZmyZnKqZYLh2
aYCzKjtvuY/prah2G6JLECATMNpFvqPYTVAQdSnFflZqE3cY3EHlFOryfXFb
cVl97nQAZq2iM7aqVgPYQKLCgGJj6mjsTlP8qe+146+DUKD5l+kOLG1bxnjy
xWRalM4RdGeO7ApHZcyVIg7FA9onnrGTN1mcL0V8hI7eL0nPmsF3FBUmwLBd
oeURcKL5UjMG6qPrqUj+o5cG3MA1dxqjw0r4BgSShYzofpB2z/7K46xFmS6i
7tW6TDvF3ShowzG3joJHkufFZ1PT2NT95Dx/75kmXKs3rmUQPDHF4BXuqB45
Wx8vxqKry7tyeEYokqIummS4w9iit3b/rTvLQ7xIwefLbZ3kUBcqgGpF5Ox1
HyAlaxecoskZqszWrNgk7FOfxBLVETDEk5PMoHYgNIntAMAMCNgVQ8fosXlT
2zmUyJfAXBGeaVXFB9oHk3+5VBK8g8e7SpANmoPJrq+rArEjLcsflTcw4ftY
/CPu5x8MHRcaVaUnJiCVTUVJVT1UJJVf0U1Df/nH6Mz3OydPseV1LJqUdnJT
iGtB657YAQhaeraYvnfyAcYBnduffxvDGQiddw4DSPDswnKOQZRoBXIRnP/8
GqQwKJjpzCQtEbvR7i9QMqQu1243JHMMhNe3YrjTmFQqCY19LL9/VaFAJs4L
eCKi3uTb2N0HyKmTIyQZb8BeAdQxbCLUFRJF0vN2kwU/zI7qE8/LyoJlqp6s
eElvo+1oI22Rzmj8tytkChPGMjZ42h65bhGojTR4Vf9RK08iGyA+c3SOQubX
agM1QMyCHoBCs+5DcZbsKCLQ+0/4irDuYILAZnUvERv4TFPz/mBdkJ+e7WLm
vOLURIe4zkIUYpECsN3RZ0ExR1IV2c+if5JeofH+8qqKet7LmksULEXFhhZJ
jnvDGvAu+j+0MWQ7jYwGxpRTynrgUbw3nqInMn5DrcLHgRJb+aadSVllZsNs
0B6r5v+hb7D12bR7yxnV2maxp1mNKsOFiDE7MuqlGYBMgph4Cn7ZbS/i/FhI
IJ/19QAIUMTq3Lcpm0msAz8F2FBqj7TZkNurxuVLwzCgADzh4Hwbar4tj6Se
Zyue/lryb8u6ZjiaSSKuNH7GUOzXsH/GZHoRsxXEG1wR3QDhpJCmkHUva+sH
ejbM4Rd4AB1HXgFCJNaxj1XCHjGxhaBjv+rzWa9S3m0hD8BRekVaXe3i8cvW
ADJXrVfNNahjRj9fb2xgW67HlJ5z5ggZMxFZF88CgnOt3tD86eKMZuHfNyjH
FZfNZinFV3JD2ktWN8Db+VprrIjVFyhgnc2wUXjLkR4VmTb8zHNtdxlgxf6s
devlfWxZAiFmQW9vHSXpejDvSP/eiwC4/f0vfqbFQ+l9bSQRLZ0+5aH23d3Q
4VSrofp7uTwgBG4uIQHrBxXyzeycKdOImiVagud6y0a/Gv7dBx4bWbcheLz/
ij9Nltz9sD0y9MjCSJDJPyOv20f4QMlFtWjakO9Xi6x1PwnfaICt5exA9HF9
x4Pi6/GCVVjc9FoHheKf9g1W9C/u/mOD0jpA1WoVuSVRI5MSeW3QhdaAaERl
Xfi+W0AREgENbDZftZWxahJio/ypm2RXl/4ZgXLuejw8yh0PqTIPEzr4F4SO
6dnvVNc2eEoXGvPuIpfmz++hIABxUp0V1WYYudlrppYz/XwtJhAHYwjgcH5o
2Z72rcrXr04SX5kdpac0daPuqX7rMcExDzZCxiMIYbNGJPlki8ARfCxE8l5g
2UQB/dIKO877u3yB+VDbTWKVF57XrzWSuEiAtvENP4hKR8UvkZDu8wS0NKGH
AKTAOWZzcPuztwFVQaPXhKRkrGb3aAoCIqmTSlQuAOgaQFwAqaJy/9iCIGyt
XnAsYGOV5aOzYG8pYgQ6RsCE3siWBtH/n6mx0mar5lXDiJ6n5EVsr+1kLnMf
uDWObQswibXezGJpcAKaPTrkkGKhKL2etnL0YcNxwlqwuclI4N/fraIQdude
dlUrDTRy0JQtH3BYxteR6+wyXqy6Z5YAd7ZCi3fb5bjQGFE5jxrquiDT4ZKw
Xb3eXlLtthVlJ6FW3ewAV4MmdvJS+8Bs5OSKXgCZVT5WFnvcPPVr6X6MwwUD
YTFGroFNI1gIeqSj7ucjpuXWp0UmQ9Kw9epkxPV0EJ79z4o+EhMUbvyzRIZG
TWYNqecVO4QHOxz4poaNyfLud8YTlsJAaSsksR84GPeoRqdgdl6LD4wG0qee
+/QOSJW23t+cZ4OVZG0ZA2EVFu5+Er2yRdus/Pni5w+QzVUyXyRn3t3qJ2GO
ecWaP3wmyM2Kl6378SVATuthxxv6eQ3PhirpOEgUaDhNTMqGV7oub+AP73+p
7mczOP0VPFYlgcPdL6uHrbfV6OP78vzp7wm1Gf6mM8c96Jopg5jQNPLDzbnh
wuMCvrgqhQxwJE6xbOpL1ei0+3itxvmEU+c1UgdiFW3Okgt+cAI9ucBMbQKP
BTC57DYzlcVgtIfgoAoPNMuiVEr91DseHtuB1VBHR+g8btoPBOu8YLbUmEXD
IWyYUVozQ9cUxnQF+7UzsxznrUHIgYdYKJ9lBqm9/jDXkaFyNYPC/uUXlvy5
Cki9HGQVTkpwnRvxO5X1w3FMMBKD2BTUI65hcrI7RG9SMILMHajstuUJjqEu
xioMyDAkW4DVDEgL8srjGa0z2inqs1F8rrY9v58Zioz3LOoZ+T0OvjZ9SiBC
vv7fMn+f/g2SJVfoSQfLA6y4EP1L+t2uMGmnaGWJigs+6Gwm3HnL/8vlZ/k+
SvQ4JVc9yGYJ77e2W3To0ktZMzRLy/9+5kAaZyF0VLariU49XnKe/Zp0VnvO
hSQ27sCEWtTlJ6EMOASbL9k42GEC9Qoesl04aJIX47++dfpNzEagibE94UbR
YdSqcBp1B3vNcGpbCHb4SHSwoPCKhlMjDR0F0TagpmRevttm3bm3DL0WQ902
gd3/xqkiKy68t7qA86RBdAkPKtFpN/TEfsvyoZxDBm2Kg5fgbTy7qvqmwwqw
On3y7FAcHLgJ3Mv3FrqytRI/dyibK29zz70FqA2zTBq9gXMtPIVAoKSVenjl
7ZIkLb2X2XPfCy0+ZQe0s/HZZVIlTJc8xOwqPsw03q9KcDLaThZlGYjN3gkS
4zo58/j942xjw9eN75UA1dEuwai8GnmuNcvKtmBrBcvpbgu/q8DMn6fbFEmf
aRQ3oHS8Sb3kKbDoV1qZqwjVYMLXn1IoizZO126R2P7i1ZhiP1WYDBu/OQBa
QO7EX6htjr0ShKOokacyBqhViptb6zc9SsJtb2ZEw53csjBbf+x92409iAW1
W4YXG+3+rszUsJjz1laNKnACHHqJHrbbOW9wmC90ZSscwQ2liEXABtef8kfh
N6ZYwaGQ+enFp3RCEmhq88CGlizx8mMv07cch8/VLt543rUwuiOvGIhYdKKd
Ae/IWtdOVYBHWdPpKb8VgobnSy/1X6S6JM66qE2q4M1jwAHvBqvpPLtRQSL4
0dfxr3Zi8dj6VYHDyRGlKfSeKXdefVIiXujskANs1KM4nimRLKgYg7uTt0aE
/VulptoxRPwSe8qxBJxjeb/boFGraIplw46f2WUIbrTQX28KkwTtyVfGnvY0
QFIj3Nm/h25ufdPHoi8jWPuNyYsRxv2mp7V4SHTpJveIAzOV1eO1+YGooYW+
OW5q/6CN3dQuFEniFJbvfAcSWsG/x58gPdaYMmmGZGJF3f2dxq+J/0gc1FAJ
CPIg2hFTnZKyP5O7UI3RY4bVD1x7+qXrvkGgCLi7Hm1ZyPt1htArCwgvFODa
C2id7+KKo+YsmTRwk0+OogqZNPEvWkJ/UK4fWc74JQvZVOrKF/X7vHBOuWe0
4BOE0EeNWurAKrOL5nyAxbQl0O3R26fkfeSM6iUAVQVxD7rM4dF5d+i4r8uG
ZQ0fyeLrBzcbW+zAGxJLgpJ4Ar7f8WqeUFZqKUdAPo87Iu9PVafUHva6fwG6
zYuns+pJJbd3u3DwDDyrMgqtyDFqryg1V5S8A/5qanb/nQcC1AoSAJyi2Da9
wlSaeLTSAdYoH/8H3sCEX+T0rZO76Uiu7VOj7KHw6RDo/E33dtUWt7t9sRha
3DNt7wIcKhl0U28JbZpgXtnIumVuo8gvuL1Ev1SNVZB4h8NRDrNMiYTn4/wq
wkgFu+D5MsWtV6PgLSGMzB0RKLNuMb0GCcs55ktBJSEua3bzvCRk5HzkLns+
/hmiUFbAP8ivUod8im4K+kV8VsT3jZIrVL5a+/swPUtVP3R8v6JGUgT3pa7/
HV4fIYaKyBDIt4HZ2bC8EFjhsjP5WAcIT0CQHNq5OYo+eG4E80cahYPFf+je
TBMk+wXKmNh5n76n0PEeMXOsH9pdH9w5hXq8WS2cuXLg2iJd7b/hTsHEY2K7
8meVpcab7lc1kBzaYJ+LpPKh1VCzeBY03TzYsBt9M1e0CfpJc3tSSjsrHBoK
WGMvk0aBw55qA86oruKm5tWBgR3kk/HQ0Y9XhS7ySFt7rbBWtRARTWOYdAjb
FSA1h2wS2JtDUJN6Sf1I8fvmcJjSH2CgKnvPjToKI3sS/J79itOVzeWcCKDC
1AlsnU/tjVcpbgSFPUV7Bge+qmDBlvlMn3rKr86MPq6KVcP7Yjq9BPWj92YS
PfO34TYh1uqlOid7mELbzb3gqdWyzIlzRE9aMiR/VU82XUQcFGrZ2bvfU3gz
Rg7v3CJgJJAGpe4Fxdd0wHdrLVbJMgGGYZAGwxH7ISiYgUhTyIC+WVOy6yz9
qdmvyMhYGI6xuZNxFp82gz9ULcOkYcBSke1D1ggguEUeurl9kgRmwyg53QE2
fkPjrZ8h2fgTwIQlLUSpBbsd8MjlQTUYxggopq/M6vZb11FxHQbjP32oZioP
+LpCRAGbazjHk/P8m1wW3yXv0xGLj5I9ymcM6Y+IhPgIXKlf5j/4OqM0I7v3
79sJ8j0dygNXDzR0Fs+j/3XD77TXvlKV7adyTqpClXyx0lpLzKdYN1B/j18Y
2jItbY6AFc52reYZv7CDeoUsFBInIG4B8Qgx4EyQb4GSSvDZIF+5OzRq+Mbh
5kx5klBO38Pmvo9wBjfQSUAucgy0GfHUVqGkBGby8MUcxpmy9gUv3mrrlPLq
c0TWoZ+Ep8QzIU1PQIV4WcQfMUcmIzseVYyHEQJTNTjCdni/N+hv7d0oHPY0
mj1Bu2aQbp8FyJBxiDLJirRCicBr69x8uHRJHQMp8YFb5OTqd6dB7irXnJ+O
5ox3rJami3vtkb/CC9QGJyohyRwrgLsYOba3OXvgw86kvSn9AZAFtQNtLhRK
aVOr5Qymqe22Me3cDw2TZiPz+UiZcgGTm9kcQMTyq1UWQZKs2wncQNWkMR7H
+kh4yrJpt1oHhZKRKjc6nx8IskU/42XzbAJdI3FRQkmJGTLW+Pxm0NvWEslE
uuD5e2PKUdzCQojiLPmg5at9aW4ewGwuAz1Wto870TSQEgeJd9VgXd33fIlJ
NTbbKNaQtuSH9/u5DF4oLrW4vnl0oKoNjrF1+ioEpnv5iZRcXMXLegf9Q336
uHjpzcZkEgHG8YpoQc+1efcLECBBBpW6tGiovSp3/mhNSAeMLVGa3Tihh3gc
x7kIEU70SxDAdeqXpBISSV9wNoAiqQwU0iya4jAbqmvd5VCH5a6iVmw8b8vo
59Tp2glmB/JbvMF0IFkixN5lMmXPx/dHR+/cIg1YXSbL/sPGkd0+3d9324EH
0qSu9jDubtcpJ0fgpaJLi4EnHO3ayHUDLOhJsWEzT7MTrC+kKrdnP+sJ0Wui
PDs+k4NgNv6iJWPriNvFJKNNqoKYr4R7yk7zwfJ0/1WNqcJuPXSxxy4TC2Kj
wzjlyR5u6QiwxGkLBlV1+DlceP4sgSp6knvSHNSGyzSyg+jIlFmg0Ekexskb
CUpHZpUTTUO5ksHgcDRmn6RI5+NMiWsUOLhJWyrtcAQZPjoPT+pCL/Kaz2Fd
LGtMeotMpqVFGtonVq7GU/O9JmrvGuK5O3jXCuNOkGZ7VBaz/p+Jesfl2xGE
ulz86B1xtwmKkmLA0YagRPQ/icIHvgk5AAQ64tXEPWFzN+2eomFXrgK0TSOw
l4lIR7iAjvtY+OHel26fn4Zq8Pf8PekC4ZGysMv9aEXEs25xioJPaEXSLpJT
Hze5M2F+oil+qb8azgl6weQMmO7QvbNieo8ZrvPTzYOWNVnss8kmq6UkLROD
sollYlNWAHWSYO0hAMg06gmhhcX1zL7kqdRbUolmn/glKe9Dxh5LjcsRVrCv
S7hQs5kU22hQ8CRGBUxT5imuXKGHBTufRXJOrqEoH5WcG8iEpLZ6IYQBveM4
YnmQddVx12oLhcFbdbNJkjryP4bdCa/htBDmqT6e2twJzZNsc6d+bdhdpX7A
M8XIBjVgS3EoAekdK93V+/KYx7aS42mMOez45rjy206PijMSkzyXfbsaWyD/
yCc3h0+qEERd1r14ydpNjwCrngShSdsqV3DySIEVcFvT3uyq9YqF/05bs/ZK
QZ8z9/vD73Cvox5T1WpgtDRmnPtmNTqIIuLiQRx+/KIMaDN40sCq5nW9AS3B
CTgaZqn7cPM2E0pzoEPJjMYzmeY6DTiFSIlkMF/RYdXWkfXLt9KHHh1tpRgW
KLcMOek90YYrzSVEEAYAaqfkCSSGvOX5OFhQiSzMF7jCnqZz4/vOzNkROSHm
rEZIXDXviSP9z7aAqEWBVrcnUAi4/9NIWNoyrUsVx5RCk+u2noxVvWqbbr6W
nH06kYhRjZw+2+rB3O2+32ju+T97Xjj4iRN1PMds+ULwh/jTRzkr6II1Xhbs
R81Kxk1PTk/idWi5rfnpVbJNFZ72M5e5aVPOrs4NpYSyuUDZG2F69pY2kC08
Kik1RpXMhtXdpfBc/qWh1aL8MUFvkhIHNhovLXfl58CAV4cFhE6Nd8MDoDKB
au+dlePaZkjGpSL2JpMZc6Th9dmMU8OldmFn6vLzXyQoxh5DBAuutLp0ugtC
kQxdv/WAGpiSFyE586Sifa4wN8K9UKiWqXLBWQVNYsFwbQrGLYwqHep+FUQ6
NyMuiS07/Cy6ItjYPzw8Vx6CkFugWvu0CDrfPpxTpsxYQlFp3MRsC5Uk9MOD
MEKScr2s6vnpUCIw+R5kI+O6QRSrbijde26PVF15Mdf2HBG8iVRYm1Jf5w58
PH2FCGDfh1GWVVR8PPqPIdLswAYwEUTAvNfFJg4UjqXe3bBhGRef5UrsRdzp
WMfwDCgXVUV8G1HHzBN0ZMcEgoL+d27OLHEw9g9S5A9IODi4l7MQT+FUycyq
yyzQuTmlsJsS00+Jo0m0FsETnvUHWXCOTsBCtUS3wYM2p1WiCiL/lvugfYCf
yHr/LEPoyCjBFe6WaubrvgC3gWdxU8Dr0KgInVQkZYaVYfzms7PA82qVrxh/
6C6WgxC7Da+CSZlaChj7mIIIErI8WNIrCzTwSDCNkBzOzJ1t6fs1laQ5oTqx
dYusrgHQ+GOi7ebfekVpfO86+L7Y97MY9YNAeqyVwbGjzET67mV4j72GSkqj
U+S0W2CdI7Pp0XvNB3ydT4U9p+2k99dPbyEOkKyFrlCcRoYxnEa8HRDHPnyU
3a0SpAcsc+CsehTpqpNXEnJW6uzWceB8qbYTveZ7Kh8hTDtYnii4UBRhjUeK
z/lzCwMG2l7JFksOV7MQDP5Otz3/s/ToNYC60ffwsm4/0x0Tjqqh/7PPq2+D
UDxr6cmiVVHEEcPvCQhvnZgEiWWh9XRy7IwBI9FE7dlLK1No1R3/spT3g/QF
zVdSYb/S4G2FjSAWCxrzBZzE/lASJbJ2Q12LuJU1vBlCWWovBjIJKW6UtbJQ
lDW9zpU+Fx4S7532rwdXgms+Q47/DamgllxwOU6XRq5Hzre1JE6Jcdj+HCPR
o2PWfh9toT8rqphU2nEQrArUngOEWiZ7PEH4DcL6BWxGLBi2Qpeqdsi1xMu5
rcjDnnsuhKWGFzbdHrffbDa7EXoOuuulXFm9jDTbVMMMHCz/Tuw7W0MoXums
k8yyI9VjwAsBMZ04p0oxYSv/YC9rbqWYT34dkPoSvx5Nq+GlNJ3zGt+8CtQA
sF+vgR59wc7j3BVVoUfD3blLQaaX8u1VU0teexdEKGQZAQS8HYwGOCzgYSaD
TsjpOBpGpeiJrFJtsVU6hv5LI7AMIQBVSF5gQCxr5L8Li4MZKcLun3nKGtEq
Cyq45QKhFmOxJHJlAD7jFr5ySsqP4PGq22A2t9MyOx6vAK0FXck/iIj/8niW
rzCcc+Hr0DRc2gREABfz3Ym9Wm97W74lT4wnsfNULpgA/Mwe05tgZzHbDkDZ
09mE+ljWRItZu0WJ9zDy0DFhm12oVLts/CIA0CcJex5nAHjc1wkWOXWlFoDr
+2d6qEsCZe5RkE/p/3GWArCZqLLS6G/69jXxkr4eaLEhN/busP7OiMjCEQwe
7Dpo7ODXAfQfpch155W1uVutOsxD1EGlXBLHMsiLCkfGkGYFNQrrzzwgikh+
lop3w0ODhM43D7pK34fO6C/1zypelaLcStqE1k6bPJ5kGiKIOe8ABF+KAQtN
cEG7seQeB9pTU7z6dLQp0czRn4x3Trw5SOxCSNyaxmh0+tR74ad4DuzG8uNw
Xk8b6Fkzk+CukVOfbTuyTp01l8RmIr2CaNbB9xrNNIFPARVnxsKG+vLPEVMU
iPbgj9HWy+xOagiOsSKJqn3y6j5MqJN8zkRtvwZuEY8+nFFOANjVJNyncNBO
+3mFhiPA4+M3plYs8y6tCsiJhYqkUquzwvU3DqaP7sOh5GkVjAQLfyb0Icah
cUN52EaWVWlpkBtrD3pcVi2lEFE0CAAJxcWi7i0QOhPbG0L3mQxH1cTsq7eq
LQqNgLycXqleytTONazStB1uJVzKiCBPc7J67bMDJVeKDHf0JOGPfQraClVf
pdD9tpEs8wS5N20xtd7f0mYJOvFuStmrCJaDPiz0GX8kxAOAOvcI26VsTRB7
9x9BkqzFR91y1gbCSWdZqalGVjKy7za48MM08mauS5M2npxFJ29auXS10uPX
5v6G6kX9ZB1+qvEzFP3b4x5/pC6rv6KgMw9FeakyIHuvG8PcA+UiiFMlqelh
lNw56XfpJkW4JF868IEvywc0DdtVBTy/GGmrY3K7Hh5QV9JFBI5qrTUQmM1V
Cyb+Xhr7yfo2aGVwpVA2WIY3deGKXM16TuTBt80ZdaGhb04XojIUJDY8M6hf
vuAgdtnAUGA/6IZs8Cm12tqBqWSx3jtHf/Nrw+GxL9E3Ji5oAiFPy4NqfLB0
9cuUScRS+haKngs5L5tv5yBAUB84PBTwjgK66a0+25Azy0+gBNeoK0Gmp03v
b9I8+cefaW2Hi9sMguiTPWBhxz4XojtkL6xrLGaXVhaSnFq2uz3Qycd9bL/F
yfmkrabKZ6Pys9q12yH0yPExbJdYFVw501Gc71DkngV0QtFIpvrL901HPK7e
psvVd/8rtF0CGv5kNTXFlzl0kyJvgXXGGlIkhTxTZzHBKWLJi14sqKg9gxe3
/dwCZRbmV7MGacoSHd2SFIpOh9TsbkdV9icZZiczNtj7EZcsdwXqoEUiOdBx
vaRLdY0+GYB4UGKmdq5ODhxO+DpaQOrYbW5vrGbVtajXjaJwEoSvQrFDVvDI
jXCTU1hdOX0fkxJjCAF/wcFYFQI54S8dxpolmW5jwIfu7p/tu+ffdcT/zE9e
1StPFm/Y8YNOHePwqZoZ6yCYIxpzvuV7lHrL5D8pyPeIGhImzAKN+7Dh58FP
bfoEOCohOx9r5JJ+EPAbQXotTOSUUp8Av+9qpGJeCTcYxFFLH1NcP8hmxgF5
Zz26FOWF7USBQG46PZFDNlM0On+j2z3B+zjRRvLQH3bvtezDBSukrv4/qV3b
QZOvZYH+QdMSYZdam8q8oyKx9T3SeDbbq3qR4Zx+Se3hIbv6b/wgclwfBx/N
R141HRDJK6zlZ4r3UUTcGCH/CL7Y0Uef4D/j6K8bicUzmu2fpvpLS6PsOiKJ
GVqExyy7YajbtXtF9dkRCsGPzTUarUXyak4K8KWsyV22M857BKeQfcl6am+U
yhFRwiuKDcrSmY1eZqVy6t0by30S0rsm+i9SHh4XNLXJvHvCTfYw2HfogIYo
HpDYpc1zHPp8+9aQdJdxxkbqFWJCNK+fsWdrvp5ArGHEwZvfgkcOZSUw6qzw
/AWHmNTePrRkxggQwgrBuwuiqJa6qz82ietKbxMldEtYFfrO9sLrwujefJ6O
1U/rqKHViKyIBVjLGDHqSSvLCwxar/LAPj4fwfnFCVJXRDHteFWc2r3crlqQ
Hxyb1FiDwLfJljaiM1WDrBKaOM60OqZaCilc7hRDoCGRmgyJfNavpGHyPwjk
8Kbt3xHKCzoaeuBAhccJb0b6zFLErTPMQVKSv/HnjYLqagwKNYGWyzSVhpp0
+qbkXW+EqsLR8VkRKq+jYkSg2g/lVaaRYGxdIpOR9fJ+7OiQNsa11jUnYM+s
gKFHOtMeWRgiAIal64jd+9XIRRaL7QicRnFHQjt+CEdVL+iQEHahBoT1ryWM
1Bw8O7Ppg5AXGQMPwpk0ZOg56nker868uTHVlybRuc4k48Zo3VLTaRJSI/Br
4M4GwiFABXYg0yivTEP7Wn97ambEcMg4obI0rBogs/Z8IdXHD1KHZiGPrcc4
qJxiNbzh4pnJlgnfJJrGM04O/skk2/lEDJNuL2/Elxl2fYhtPspbIyDFyR8Y
avnh3lf9e7F64KKRob0bSQWgyy4v0IJlEDrRa1Oul8nPTMOYjXHVMRjGMEIB
OWozM5JKS9MvRFt6t8PykD3NohFDl4h/I50A6qNaWM4X/r0Bvi6rH+YQMhfJ
Umi2Ip48S2W/ZyIJ0oVs1wXey5QZ6bJjPgf7GysAv0exwSv1SL1RjJPClMYC
ZHS38TpE0Aup6CmxoszJlLB38WOYf3CR4SBNfmOwnKDrnGg3GJJ1IgVvZny6
zNWOzxCec3dRHVB9Wm5hsoPPbAkfC/i0wc03rGwgusI/+VDDwct01R0jlI/t
3L2BxkNZ7BNNgklQ+HUeq3BJp0obaFG8oCnfL2SUaIxjZd/KHkXA24KdKuX7
5tNTCxayJtCd0ic4G+TWUz68Sb8xe9Ywzi2yWKJY0j//GJcIVNlWQWI+3O3R
hTKkJA0v/QPN+kKIsjkntgmvHZs5Mrsih770iKi1AsTH8fRnEUQBSI0mhNR6
wtEQ5PnuGwSfEmwHtff5qclu3e+9UloDJm9mLhXZZBOga3+lLB6+Dk/ZFTHr
sh+lz+vkLwP9ZdFCQwXX7VdCuVvkURfll5hc4QjdB21SCRK8c3XcCwyV+Lxr
67cWveitDlVl3HzoIQ40YZdts0ZAF7t1/9oT8cnCDQ0JY+FIVyDiIw/qnQYG
6lgLE/iGHmfZnhhRotBaOf5AT02AKCW7l3RTpRjDhzLcPLCuUQinO27dIdz7
JyfKUe9w7WagLLDc/z0DAOPFFBYriYFAHKCW2dKdQyvMWnDAxQ8lb89BZEKa
YtqlXroJQF5333wFXou4+7unzNTu3xM9cm9l+3O0DbLMDs62y+4vXKM3H4EX
U+vI1FiM0L2jvKnkHyr32QOcba9MxIT8Nwwv5Ecsxrx3FbhcdW11Idohf14x
2z36QiPdcGw2LZDoByESvSBhwTOSFy5ZjGW/W3dfQ/y7TdchzeC7UIvq4HmE
uzCUaEhyxOO7aCC7VB7zscwmmLtoMBLe/x7oiDSbALCWLC+RVa2ScO3sNeqS
Z+j+27p5RgGjzn2Lu94dGAJka9sffKoWQujjjdIZbmrf1H1uLR2waMPvm4OS
oJY12BDE6QepqqG9ZB32

`pragma protect end_protected
