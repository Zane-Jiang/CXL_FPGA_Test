// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dvIGOWcxJUL7P70kZ2/CsVqAOW2P0bJ1L3I/n06VseLxC+6RWWOyjBhYdozd
OnGPV/wTq6xYWHICwba1UdHs3t7FYBQYQmgHY2FtjmsfNluWISQT4jtGpCNs
y+YEi/uJ5gUAnATzXHezNQMOtD1RvBbQnbaBlyFXJ21nJF8S4yqL8hxQ/2+n
ONstttuXXjkyxu8YA3HBrOXS2D9VAZRxbAUNSK2yYTvt6TWGR/DtqT6xf76q
UZOrv5d+YJN1DeOpb+sVZkEbqbZCJJHT4YblrsuwAP6dThb8UgCQzC3CXHDG
bIJfTtzessB21rzLodNghq6GoNu5FXjmdx5TV9aXfw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NtU0HN4EyYYa7WoeTlqEF6ScVrgUs1qgY6f4WDCqUdRSe7s2e9sYCmFVTqgd
Z4FSTRVTqHjL+nBLobyseJWj86eEULNHf0wcRsSRNIltkTSPu14NOLMq2IMy
h2FYkhhROOuU47NfzMNM5nkIBO1g7Q0DTxzUL5jvkzzqnr9RUopQsA8VgjFv
uQDwQLYpCz1s7RcRb9IyA+GpSX1aJ3APNI9vW5Jrx9TBeDMBcCmFVI5tQIde
7zbIxy9kWW9J1WhaWzs/2zqfduqLSuscnUiPudujd52qsql4+M9BFZ3RRvOd
EQAvO/HRyRSE2vzFfmo/EkO/m3bl6UxvSy+leRNsjg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TpPwrd2S/xkq0iZtOowtbehEQpEVid9Td4j4S8X9D6fb+65+nggj01B714yl
ICRGpMv4ZXiFm+KWRipCNOGmdA4UJCt+//mTlv865OIEJS0lXpDiUb3J6om4
sr0ug3ehc/5wFuh+pftCjmbTbYZzU5VMx7IeNWpCskNVYEHvFv0Y8Vx3to3o
n6c4q4j/lvu2acOofymK9l0MDXDG6dxL15XzvzuWxSknCnUvgNirJW3s634E
sopomtkmjpFFU2R3unaRlOo2fkO4vyZG4rS8rIqxj30jeCz+6RIiZgaOs0fu
vpFfgM2YcmPHA0oawPNGO7Abjj1d91FzL3iY7RIksQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V7r9sik6tFYr9J7r/uvjnIIrQLJSBIZ0VJ8dVFD3MaekMtOv71WPwzuZCgC3
MbSEh19bi5G/cj5NCliguQ1TpDq5JxusKFuJKc8d0e/HzDhRZFzQMZI4aNWQ
OTRzl9D7zaEiHwGCUdXz4C4/WSgURdUYDXlUb9IlLm6shyJVIb8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VTtbtI7xg3PuMvkQKSZ79NiiitVYZqwbgFkl8ATukWHNehfjc7ZsRPdDqXNn
w82mrwbR/KFXnxOitY0lT0LSQ1lSsn/cY4dyuFHk30DFhL/0og4Lt+pM0aGa
aSYDs6F0abx5QeD2drNzHHXKAYFmorCYLQsgxFvWLtocrTvknuAwq6nUfvoX
tr4RaJo9BJFaHlKHhlZWz6yqO526C/j/6EONLaE9zSVQHshvhiAYbGaDVuZr
DT9V6wGeUBjbl3GDWemaFyFeJG+9QBL8by1PYfbfqcAC0mrUPDWrM7BnS/3V
e8mnduzCLskmhyxNqNp2+oErR39DU5+a8xn9n9llhsZmf4Eg18jF3vflCoi9
qqW12exaF6eKexWO6w3I7ARDYgSd0SGkM0EEPdTzv2gvQ/Wnj0h93lKsbcM5
iLPHczAz2G5tSUT7qW8GGl6aG5dPqSuO/Mq7nqBc9AybzYiaattAK5AtYQe6
BKsWmajfYyB9hOTLDdz3M4ai5um/dPUy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rRAMEKTO93ZEFubqXd9Ue6AgdBPIoJlVWovmtzUdzCUnqL5V1ovher9R2IBJ
n4FH5o+IfwU1ogwgdQS7oPeP0gmJjse3LB/kQHn4ZEfYbTDHIeTVPFTAFafH
lvUVGZ5Bs2s9qhABjsHCNryPcXIOcAOpoTnpvUYGpHw1s1FxsDY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sXdW7HchzGxXNNgbdmyONeoGp1phi5F/iFbOiGX/627mKkGFAcjki/MU2h9r
RE7hmIWsdDDa7PpTjk1OZ36LdLDwEpGDUE/2VVgFL/y7X8QXmHvTkB3nJMCT
S+WVzlx+b5HXhP3LhXuZJKc6p5/RHF/upWi/f5koby0z2ggZeFI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1296)
`pragma protect data_block
kdPxqOvOjG6tMJH2tD5nsCfylpVBdTIzlrQspDyr1uDq1f3j0wyUeURwWTAt
8V+acGnCc1aUa6j4zAvYVHopQNmvJ5fTjO26S3jPIp1Nr9x1lucX0WqkHmZB
9momavlJwjW+MCslEsDX+w6MfdFBuFCyJq9AKC+oLNKTwzSsA3jiQim+ySiU
TMl6d1wASz2E2wTm5Ld1u7dBUQ/Oehi5c0Rz6wr+epQsNCKsUocxFhFmbchv
oCDqODLc7Pok3oCQ3Es5soVqM++o52Np0R++QELlJf65Tf2Ias/t97LcuIpH
pe3YH+d+f/l4YdpJCBJPY8c4cPhGQ5z90sF1JpZnVZzXYMvmJTRcSPkk05om
eAt+M5tnWKPko+YTzn0GO2TI7i0jjLjmqvxND/viwDMuRYcHuBeoGSAcoN+T
K8IfLer2jIn4uv0mTZnYq43ZAktdGA4OHHGC+7yiDTTfwBiVgoPwrWyCWq1e
SUDKmPoPwtSSoM3tTzxaCasWFk3xp+gbkHM4sOHildyRfQRXHfBX2nf+RHEg
MuIndkiL+jvQUFcgOjReK87NjvJkHGi+2vmH4+5RHQYT7FjZ5O5HpRq52XwJ
xnQUHWFvMa7tByYk/XXHhwwgFWtrtH3i7Iudhl5waeob9irf2I7sI83ek1uk
FcUbbpCXoNb+JRU/FlS/TFmgpuJiIWYtop01PKfacHqcxykY343542QP60bb
gi89TCBXanPl3GXIZzar66CX1Fs5AwvUXVcxCodHNr1oZAfAOJTRQSu6N2G5
WoT+lbJ62eqJiiUaBsCPOYKNDamfhw5uUaBsAILt2pHFl4J4A5yJWOteqGU1
iWwRtijbzPkuKtDr8mrYLWhj7CKzAXNrNfg96CsYq6cRjVUgIOKu1OsfvJV9
AxUUd9uzcMZcoyrjvB4S9j2BKPpssUHmEibioXm0PgyKAEo9kUCIn//mmLey
3bANYkofLZOSw0yP1/khViIW6KWLOwa+RzA2dMOPGpkHUwXce2k2M2bGW84I
vVAwYJq9rq1HQG5MxjKwStIIMcRwH6rJhMo4AmwJH41Hv8d/YpZLWCb60z0V
XACzVuHiHI7/Q7gC3j3MkpTw5Z9WtJCW7llTjWtcm82JxFVVOes/R+zdVFKh
7LavnCKDKVtYaTJzVGsjImY7aMIwi7XE9/5E1uujeU9XDtOdMTLvIR4zEMO2
BQCXCMJLgicyIM4+6l5wZ6GdjYnmRDA967HXhuH3JaFSUZTjnHd/tucalcBA
d6gVpV6choP/mZJSGE8dhj19LyQ4roPvhS6ZTqTleDr/j3jEUD2zAShfMVZD
XYsB82Np3oiD8atnyWmec648/DiSfpvM0FrmD1HUdhSi3m4PtWGvSOfIlgPt
JiQwtuVi0lV8wz01s+sN+AONkxeLSFeKXOI5OV++MkyDLkGk3CjsnCCiUJ/q
akoxZyi+Zjb/+Rc+zUNO4IPaZikoF4de9tYrTPkTUkRL6iS+ZJ0Yp9ShO+2E
YunOSmo9CGHlgQ/aUY8Ki8oBglMCx2hLqIdNsgg93AREJ6eOGw6zhn2rwGg0
HizqyajXOBABbkn1pXLSQmYXhBigmIrKs5kTeSma+VVLwIvPrdZ2rKw+rx4f
gDsob9+/JgGuxyd+TC3fEzdlXknQRmem+NUrqqSZaTQigAoe2zbuoM85Y/nu
j/M8RCyBOF1MdllvfN4Hrx3UFMM1nVvFpJMAj4oxufksbtoA

`pragma protect end_protected
