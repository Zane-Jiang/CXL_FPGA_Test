// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fNrSaKDwQYN1BsFP/JWTmht8N9iuHBhuh/RTEM6UpfVnxC89bIr/XaKaFWna
1rb/25SmnTKLavTYEV3SgnGCxn+R23In2IfhSFMtbCwU0ljoIfJHEOxyMaIN
ri11s84J0+F7Hqq2e17XKdVJ1rwSAaeTPezoq8qcHhST0uuLuJdrMKFG6DkS
6+EQJpKgJo5XloTTRWTM9QFreCTdqd/T5+dzFe/MXyi82nzD0VBdQCuZfSIR
RygUuyKY+ILnC3AWadE8u9hjtpxpqYvqsAB1jUmu5mgVihX2eIGU/26IR+JM
GISS+wQnJy61W5YGz3jeU350ZldtagBbf+Wr71ONAQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VOhMLuWeXVYhU/ZdOAQTu8tTkG+qHDgQriIZ4449GuEUzcbXg/oFeMso5qQs
TkA+SJ0mzvjx6+s4xUv0ymHeOf0ViFO+iqFZeGqsZjzMEInk+6DfeFMNwzJU
X+JU/MCyV90i5mfL+9SmDwXZ60A/6WnxKJtmCGLvJgh4fZzR57NUxEvGbh0p
UiBv4r/UEGiyx2mx+KyTEIHuzuOzGK4ci1vWrc9sYER1RNJT8/MAX3iDywr/
CWVBWMo5nbP/RdWew3yjDMhGEY+do0uMXuoC85nh4mlamNQZB9mtJzLhGbZy
E5aH8BWpEQIdxAE7ezKsUsxCfj5i8NPn9czMmFnxNg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fUrNjKLho+RZGIEa2L5DwyXHidn29txHuByPCurYOwx22iBA/NjL0fOn+36d
2JT+He49ePjNbWPZymTmkaLfcW0aAJGkKUB71nGXqyPbQVWVUZrpILorLKsU
BpvtmRIEZJtiGsZpvp89BPmLgEnlmb7gOLqOdZvT7rfkzDI8De1w4Nlzic0t
Pc1RK/peFDOpbBbUJXWc4iDG8Ghjpm16GulhayeicO5ht1SxHPAPlJeHBRbx
xtkDf8yehpabp7DwjYQb82Zh9tXTR40Nv8kj6OH5JNrQ6znIDy32gF/5c2p5
zMgrsxEoc4u9WjJTsKXoLpJeSA1//sBrjGkcf/6tOg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bO/VGKQaOXh0CpJiX9OWAijWB7+xbYrcSWfRMDXYcetxi7GSIMl+syA66cJ2
sMJs84X32+RHsRnFAVslN9B8evWGRrr5Qpo/OyanGoYvWN3hJaAOjFwcrsGc
j3Qdo90YEdq9u8i/rebQGUDqgNeDRHsbAmuaD2d9Y0QglzNdQBE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SeAZAXS/aptR+G7LE71dumDL81aJVYN1GtKmGoI5b8bfYESWZufludHfKBnB
MWo+Oa/OtmKk0VjGoo1PtK9+sU+t5zNckESb9iw45Co83NChweWaUIiC6vjF
bXsl2KuV1aDA2lNCjirekEkgr/j1KJQj/qyGKX0KX6Pq1gM7US650GArhBWS
40IeY7vxoxbMXweSb2hfY0YEbBKkNfZmF6Ffqx6lhAP+4oG+g/PcenryAGz1
nhmJUY8xBNTdgWDPuj3AdM500JkezOzvwyton6VB8BEwGZFb2ej2u0d9bsMV
gh16Dmk7JRxXaA9UCtwR53ExPcMC86+pnkcfiXgBRud86eUIgiZuQqjJLG7K
3zSDULhDvkKZ631aH0IpdnVgX4Ga0LUTP68BxxP9jaQo+7QBAOvqXBykGyN1
JAmXsm9OAn/u3fq6hulX6uB4JHel8izLexjtB4gO5rQOwmzmPfJV//M3dohX
0AOM/xhkf1mGJgbbOCvKtCMrrLDjT9Ma


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FNp4E4pkUKxETfyexlOziIf3KG1w00/4ZcflPeyvnxuixPwXkYx6zVfVye5e
icEEJEltxgm4gwF3LgMrZ+QV/P9Gft4qHy4jZKk9duSIr4eGXSEyw7uesiBl
WyJZPeYUPFmBwzhcpA7ATOC81w/FWZVLib6gF2CUl4nWtzUE0KU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E0M18JknTCbySh2jMNWZpzxcgtuNjqNpC08g4l12If8zZFQZKGiYiMOOFMze
1wQHs9g/S6ZtDy5jpKjgZr9MgYMT/nYixpM9wGCM+Loe8Ztj9OaKTOB3cpPO
hifAXywjIsmgDhpDEY+aF4BTb5/n2oVucqfTbbaUXcJ+y5WagU4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 119040)
`pragma protect data_block
tdZKEaomrbBcccPTk1yrXyc8K+YaQR3xWkZflVErmE+ZPUkBAhSzXUZ/UZG9
pf337l7wzLeX0n+Fc5GvTSR4ipYspc1KhDtTWAL5t6ITZiHwmUnDVzt260nl
EKgYXrXSzYbE0iGRXaRRl4xb2o1yOBuQeYmwrf4ie2gxU5ydQoC7k1+/d+Ig
Bn+3f0pBaJHTAA8Zyl7q7oGZlVbM14i3tUZOK6AIj3rWHn+eHuGJKqDIX8Aq
tnxwOue3zbRFCRysQeidCiR61GmLcNfAqMbgwHsAQ3ovjyl4NY2ojuOlmG63
5HyFvfHeW+v9nLouoJT12T+Q58dP5e2H+V/vdgx+eQCyvnisgQ+sHa9j40cr
Gf3pc0V8ygVySTUAI7xKT+gXsoS44SDUz6zzZ4bOom/ounN+gdl6/s++0u2u
c+iddSuPcFDZHAVI3WX5JtdGVpeguPiJyM56zxVFB1MJXuhgci1cojKH5fcB
qbTIpH0BHta9JTn2wuobYqScDyG7+eb8HSzULEwVcAO2o75t5biI/PUzR/jL
ouexCadBO79cRgaax1+M3JHssdgUyE967rLkOmwrKHd68eYf6dDATFX0wuaY
22TaJ0yuQ3pqZfUMuUnp1HmzQEZVcq1XrbkI0vdGLit7KnVLjOxauecU+Q7b
DBMn1H22vwYLF5G9/zv4HjmqMkam80bKC5ITxKu2D5d4/ZGB8FbUbEP9OzQt
x1HXvayKgY+eFQKf0p+sasc6fMHqhICD0vlcCgUfJCyMl8c7bSpDDh92gdDe
TvADaMuNBGYxYv7LPJPN8mgqmOiJ5C7z5fjRj0GQwJYag8eLGSgeeuwLLawU
dCwudFM0b+Sdw6tsrfNsLYvu6DBz5nTahDw6GcE+OZpH4J5l0ShCL2UMPJ4K
ATMb9Aw8Rca5vPmy69aNNpiz/xmsvSyK8MDyST6j5kCVGXYZu5aQZeupyJ/x
DmHqXqifO7fjnkWWz+YXL15g0xNCip97dfhZ5EVwbjDywZma4mwrZu2f/OU9
oYx2Hjgvr3xwjsqzm2fBqdyUvPr3VweVu6Psj/g3yDV0b52x4QoNk+JcD6I/
YonJp+zSRLzvSSqnA+8CrA4UkoSGimzwRwNgd3EFrW9cKti1YrOkBjlcyGhQ
+IhrncUqdudvRPx+gd7IspojCYH0/TUS404gTKH8muZD9DJZsRXj44pya+Es
NK73Bvl0Q9HflfPBk8pIXZw4IjHYPgFkwMLbQQYS0k1u7AuNUSRalFwvd287
ctXOA+ZLLPUbtOoTfXs2Yd9v37M9BNbtlpNDU9FhAUVlErA/lp3DIviwrjvU
AH4F6cXtzqty3ADhnxShBwW+MhP+uf1gK1lZ5jPfzTHOktKiscv02nYxMr9q
0IFkLZyPYMY++h7WMZKhOi3GmJV/+PmI+Ci9IkzT235xGUihu/NLrGa3QJe6
eelLNetGXlWSRLhbq7gnlJANpO971b7FKUJYHqhLz6rHld3am1h0TEq5Fe07
qpOFpLe4Lu4lFKO/cXuBhOxfYe6GtbsEln/6l5ut9C4R5UnIrSI5gZRzvjib
2kLcyjPBPBkgOSIMNHQiQmBvqohpBvv3njchCjJhFylCmVyzk0Z6LWFTwc5H
wx5A36qqAJZesaUs4Nu1NCbl/JDlE+GE4e4Jlrqs3+SHvIw8hCro8P7rzn7L
4yJEG92+hmmHcBfc6tLasnl+J3waMj4HCtSsFlu3hsuaMDaPyGcfs0V4o/2s
yORhHAPIWFwSSfA1TieFIpKr7pAkwh4cxHZJBEYFzDUy4UIGkAGHmX8k5sE5
FRsQuwIm4Q9VpHz3x98vG5FNMpttV6PqcwndxTKTJz9xeewPLGpf+X351SqD
CwqldF/1nQ7hLz8UDw70sifdGjDQc+BAp84X0o7BBv9KK0GruO/LS3fv60AP
eBT6JXreVcrD1UMRWnvfNlGV4e6MB+xSPKC9WonCvedWrHjl6T7ConB0Udl7
TKTAMK5iPrYxP8sLWKzp+ie/7AtwA0Zg5+gZXxySs1YwmHjYOVoV8uXNd8AD
TWK/kPIyyQgZEM+nFmWOuV/yJedQlqeygjOwOQebTLeZ5sJSmtT8ejlufqza
etxqOGl/qHluaH77wlqECfjFH5OajyBoE3igAuA9aAW9IAI2sfSyJrIBq8Vr
VxvPlRCOiENwWW1EMUcFSZCuP+uWtn2sZ20lm5NzAtQOlkmKuzakgHl3LQTy
YExVqRAJ3rKwgXeyXQMYHpPOoeMlu7NHXFj3J94uDRVKTOsEmjKNlw+7CLNe
a3nzxRmiCz2S5u4tpkhSvWw3rtIY12Ahc6MhMvuz/xIh+L7XPv4ahak4YOK3
1Gj+wenSAMWenwT+DIwLALpTev7JjmjW/ipJqEaHPyrrAlp0sy+dF/DOz/Ia
7l63hlVPjIPqZivnHNpG2A0sgA9yt5ErWFVy4Zi02rawZ2qH/QS4ydPcrr4u
fdwJGondlPxFpEjQpWz+vglB50iP4hgt3xhTZfV9C6Q4KPieXp4T0PfD2t0H
NLe+zGGtLX8+TPQa11zzwNPmRfxw4NQust60ZOC7IL002hwBOQ7IqrPR/ZYr
TfS7k2ixFGP6Ne7ZiBo5o33je7tKbj3cqL4Gfk7kKeOzMx3LXCqn5sLHbOWZ
A+xyaGnn08F1tTkNBR0VuSyhAanvXA7OqOWwJyYYZhjc5ORBqjGSYUa6bnMN
Uj0arA7Z827W+hht76Rt2H+hNlwOlqFMsz9DF1EK/tgtRv7XrBNVBd42QA+F
wDjdSr3Yqs8z1Yx1qpE0xRnL3pWApLuUAZvrEbuAfqpZXkUnCsL4b1Y9PRk9
thHgbJTTff0LYQkgE/+lgA5luNxuo7rRV3Nrh1CZKOdj4u5JJSKNPmiX2gK0
dsWsIbB/0wxWRjBiYzWHD1O8Wk710dlqdi6oOGdGuZiNj/tuJH20rf6zADhM
aqgpQUqXu7+Svygp8dclz4LDijMjSVdNYRn4aJZmggGmnBMQRhHsULjzQCPd
oekTSJk0Olj+3U/w2qIuEWoaoSLtQ3nFXHfkZ71Zk3jUvaH4L+Lv6xV2i/xY
jca3zpA0bUHI7GasRCVQIOFveS9WhBHNfs/xa667Mz+qfqGXDu/HZC0K61OK
cseBO82OOh1UFnLn9KMlij0IZ3V0Wm59lPEuN9uAkp4Rti6x+WbZNAiZZTIr
xs1VwtV6fXsEQbC8iPMc1fJPpX+eoioK6h7iJHC5oW3AfFwGeQsp5C+vuqcM
oOo9o/KkV/F+jX+MQtoJG3DNZelZHM+tlJpzblxuiJFh8KLS2ddIa4WmNE/8
s7VDxjls9jbTeKGqmNt4rI7Wawab1OpAaboh/wz7Ul+RMDJh+Iu6kb1/Phrx
BzqrY/xRdGRA/Aaya1r7v7x51t7VdFiCNqVZqYPKJzdwXdM/b0uLS0AYp2u+
KiBb31q8NklZgpQCPROmrx5ZGb/LCYjKnEeKI1iBYgoBfsqG5gs9dvC4TATV
8S2TapnYi37EyMH5euCUbkdnOunmuoCx1dGRjnazZwDESJW8SbKBy+rAimBj
EPgFMOyHOq9cSnb3qlFoSmQZr8WwFpzrms/UOz7aPaT0F8eOWKOTD5Xa/Dzt
sh0oB+OWkt+TOJMPilOLPjYfZhs4XONtFT4HWj8rzWrd4xVKMbTQJgWe6rmw
Mwc3E1mCl2ItX9UMn6Nxz83YNzZqCG4cOj49glPbUBUcWbymUOAwWUckfEHI
1NS8YyfeCKJRlSLRaw4YD5a/j1Ne9oqMlfpIoKT3/K7IlqAUP3SVDLc1crdh
MQm0iJE/4YRpJAaoPQPQNG1nlX6imPET45QXWh66dkn/FLv2+nnHOHOWnG1B
yRsUhgA4O5zXhFm1D3xOgfcDB4xtXDqwJV+KEU5U2QT8sfr05kQX2gBCeOiw
0Ms+5BqtfWH8uXuJR3xeeFejiG2Rj2PVuHwOioEQVxdQKC5E5us9eL3ryyub
nc1eaTnUqdbUKrOzy5xfoeZFmEdtbMIG44WXTZ3umZA5L3wu7pvIEHm1cqC6
JNt57FaFEJoCkQ5L9d4fg+jbDAkk440xPXn7ESXa9KjtzLC5nBR2unP1/V+r
1nhPchkLgMA92k9pY6zC7PHs+QaqrZEcBWEwu9fNN+CjRnCcaIL6VkgnJPpH
k0yZCQc74QlLPR3lOGgGEKAZhzqEO2NWo+6eKXalad9brshXnaPQKN7zGt97
wViMbqS1c4B48VUC0TLMHKRjJNpiJIGgs6f3yRuq99XZmMClmt/4JN59f8Lj
1xnq6Ow9qu0EkTxEjnMOKfvFsBUEYY5IbkxsxWnOaIBj4GsFeCfaG5PdyTcN
kFJ/rYVVsO28rnAOvsir2pUB3DJoKpXxI8QkOLlMgqSQSsATxffySU6NS+8q
iKHqe1wf8ppXCTTBBOR1bYqv28DxL4Dwmerjs9CVpMW/2Locmp5QJPk1NtnQ
bEhXsyT4c26EvIJ5SLNGK3dGLbnaQC34nA/01+lVdhZBqPE3H8QbUiJNRiJH
vSqRjwfKLw3hFRmHq7i/oNlwZLFDeR25fzk9eOkoOvUhf9sue33CWJBcQppe
5938jX7uiY19jzibf8arPjKoEWjnl3NLoF+aHPx6JC0u0+Hv0x8NJXxkdmiJ
4frto3YCdf8GC5+XzNEFzk3f9hijcbRubJQTLy4hXuBgJToyYI7henadqR5t
eG5whgFi1ilXqmu1bNmDAFDDZ4ZJyrLommVTfciEnUPZHMIhREDKN50q5X4s
j295ggjhza6EWO7uE08r1k3JBeNw50+WceL+tkhGoTHvPHdU8QbRaNxAvkOi
CemvLzbySLnF0Wj5d8MOxrXoFyiWtmLXZsFvbV6CXLLBpao9pDNVrH9DIfht
jSV8kaQF049P+MSp4eNj4Mv4bs0V0vnu3bT0a4rFoow/TnijiHDIz/cOnHiO
e05wIsBPhHfjLfFZ3OM6TEooyrJnKfqNLVplA9+JBcDwWnXSQYzZp9as5ut1
suvahP6TJOg0jtKH9fvDzytjHN3ym9c8XQfE8I+E1qAcedXQmDmlwgWaDh/i
34feQyQdTpG7smAfCBMBh/vNg8KiOqdrD0XbvDVKFi1aoBdGc/2ZLkdnCP4X
nkuENP8otqywEBiHs8ujavWpKRB2Q4qy2FD6z+ja+iRNlD64duql8nFJ/10n
+V+I33xYC3E8JT/uFL/lbAZVAEA1QLmN4/o4BJx1VA4+lBw4wadbZkxUhEuf
T9V4n716VNXzRSfMSQyLCwNBf7/C291WmL13d0jOeyDx6dqhRB4/0m0YgIyy
mDvrHjDEpQeLAhLMyx9uit1tS6GS6uARvNULoDPtcL5/n9Qrta5qqbmojawM
EIae0jIakPEMKt2g24AxGR9x24OibtPsyRPn9uIPdz4GEVl0+P0NCiDwlLGE
s2LQuA8j3D4GazikBoVY06Ath7zW3TzgSSE1vDZ30hwre9OWnjc9uGgUhXkv
QghMnIFhzf0YV4EVsi5CjI/8oJW5r1cYAGQilo6sEXUlZcMsMGZtphfG7Ta9
k2X9YgyNXg8U3/B8lOUYCMvJqsuDQhMlp/dbOm7W5x+IpQA+Qr+9at5DtjCQ
i8qpcVbHT2cHovZgkR7xz09IQmvRkZSLBICgi2HLWt8GDK1kbM17BXfnpBkI
FHGltkeO07wZ00qj4lbhIiHEGNnY2CDL8YSEK0CO0IAJEP3+0jKqN4FYGBYS
co/7f8nASlJV+Er8laCWVIC6NoyAh6y2M/rI+5CztX0lZ/LUzAI6c5c6xaMs
vnB7dCPEkd0DZYbghQErpsG08Kkm+VNQ7hMseIzavAvYNks/TtDjVmMHXcr+
eo1//fi0UEMNRuVKFx0WBQ0lDLSFFFhd3pVJ5iid8esRqu5L0tX5FVJRcrtL
eNNMT9FknptP67Y7UwqlpcBcREDgGjnTcxz4fWY59Gl88hQVqWsoJReGYFpf
14S70xhMrOyEQqRc00TbZN/6ZFE32mUmRQA4ArN5jpyR+t2KaqH7tA65AWyR
B+fKVqqcgZhLOTKrUO1QMWzox6vZWwxf46W7kRlEXOrf/daDrQYprsJriHRb
rinDyBsHOM3kDnhftBN3PnlDo/r1I/LIVPQF3PXZByKKSm2nOmjKYs7NfAsS
+U6cyzRPe7LRgAUf+PRIOzMh2gzQQ/Rqt3y9SVBgdKbPmXtH8FlsQZlf8wuJ
IdgyPfQFycF/LNqAOrL9sEozx8fY+aUYnFT2mfbfv3wOpfhU1/7WaXYzfXm5
HaoEX0kENWHmtLyIz7VYurziPKc5bgpb80jgOWlK87cWUsgw2qx5AiaU0e5w
oTHgUALMauxyP8snDeL7dGT7Y5pfUxnk+TBwIe8WCLc2SUQACl5U9Tj6vq49
rtZNwJqwsUK9Nn/qfYOG1mN116zhUF23G5wV8r5OJ/puAXg2a5P/SesqJejU
RjOsht+u2LDmh+SZHTyup2Tm/nBUE7fU8X0zzMs5SSkbf/KXR4GZTs2c838C
pi5t/MlcnBdwhTPBPTrGeDY7vtdjnm1CxIJ/wuaJNaMPbnitmE3hztxZeQ4j
B9ya3SMDGbyorVHvLv28QwMZtQ/433FhEhyOxsFbIqQEXZgSh+72LNMmMOGV
XkM3MEuuXeOEL+w1mylgYivSoju4Swy34/6ydpqpAtsAUShAH0O2Qae8FobV
Ky/hLchfBUZQAdvpwR566XH9o/Eq2I7ahWSbqTrfxlr3haqbEqK5y0P99kKI
S7IVq1yklqzHwvV9eZsh4LtkB9f/mxmLadVgPwXkNmfNXVoyZYcMFaOCsTtl
sd/jmdSYaWmykPEWul9KYcxCI3rv+XVDJWhx1DJdaOuApQI/E/rj8e52YpcV
85Izwf5A23NHA2YuNAvFOYUkCNTcfsYH8U6OMgZwKZmOKroG3JeEDhTrfqgE
mVvBCAM4J3QH7Bjr1sIqA7ZGYymZtQBwevvM1Y8dXsSY9er0HAn8sxzarUnE
uAFwW9pDANguJDTXsFbne/WsshT0uQDut0qxOrESLHY+KdSskdttElSfPpOz
4UhzmKD9xaGK6usmulsWIvTeyqX1Gr2hN+qGIBs5qlouHbV6EohS57DEKiAS
CmWDdAjHgrNX/8XkhIjCIThC2qhrGIk9EMXkVsQlw66gIGE0+TBSffAiH8S9
L1V9bx/3XBH6DG5q48pRf9NhOHHDLEk5Hy+wBFSJju65dqvBWI0n8L9tM07s
8Dt20auz8BVvW7BSw+BqMIn/MgnJKbfDwZ348AeFDabA+LJehwwL9zCbZK1w
G66KOuUs9PoSsq+cW6WNAK2sOvJzigme1SDg6HOmaRHTtWHrpA+8TlXFFu0f
0urdWRqoj3wy/eK/Po/AXTWP+rjDZpBOJgE0k7HfWEjVm5bqwOM/Na1b//Cs
hEIqByq2HEzgXx1lKt4oOfCneeOsHlj8uKyv685/PTBgcKN3VvuwDdtSP/ZW
ia5YUb1KEFzfun6Pm37u+wZzGy8yR6QOFLXkkeYcpxvUrDikgV+po9N2Xu7f
NYz2KeovOTc15dQ5/WMWJIJWNDKXIwGeMvfcB3LiMurnzaWMfolMPYxlH3Dg
X8BCfgk2TiNAsb2y9CGWdkVp3ZaXV7TPYrbv+YeNXXucwa9qFqoGoQUpZnv0
ECKcKPt+OmNF3XK4O+RqB0RfyIgh6NEYo0NLqKUBiPDLISoa3yOCuYBXky5J
/qCVzYdYfdrBNKeOD1O+qZqS+MN/CViAu6+sLvvKfPy/v+x3u7jKOru39EmL
pEpii7v7sVbF2k+grZGdng1o+7IBfO8FiMWBHtsBD0o5ssQ26yBxs9FVH11W
hHymPGx7jBSSmZWDzocBS5GmYp1Y+CLjXsMkkSu23YbRHPuoh5Iuw7yCkLGJ
upac9ofhF3KsCwX0FWxCR8VW4vDerH++4HqPmgJNgWggkMPmengzbtcRJbpG
SoM3GbaMWLZwV1I3b/yEDFh276wBrQ8LMcH7FG8jnQGrjmowwYWFlbwUI3Fh
AczdQrVswowV2P6vXao9dcA7T67hLc6H8rXBwuMBb3g4V9CVnIhsb/SgbgdG
rljG5Qzp+nGVw1g64AGat/WPyAwWXJUqlpPk3yEbigL2rQIqmpuEV1gCIp4j
1WEFmxTWM+cNp5iZdnmNDfIiA0M8g9FkPZqflodnRX0lPhqHEMyIlqZVTBoj
IC0tWl9B0NUo1duJzr/2OJZfewl1ar6gJUZTR0IQzrm5+xpybSzKQYB8SRn4
1tpOMsckRlwe4mNdmviv2EuH79FvX8RJXXDfKZWFP7UBmVElaO1QC+NJGNBr
cYiY562Cl/DylSTBtWZDY/jn8Y/7kdmoBDUgjns4yrRWi1vQmYgNQdenTyvs
KexnGpCUcrLvyxZZ+rTpWCUmYWF/HTarNSYYJ3IijKzqvN/4z9UHyfYXyMvH
zX00y0dwjlAw2o+OspCHqtPBpA+uE1IDLL7PZkKMGAT5uFLhjggMNs1I320C
cN6KudLLfB6q0PwJX4cX2D3HPbUNgU20zD1aeMuEVGTcQGbkgDXS8mbFeSYH
p1Rdx4Xzao29NJUwlwxCYrj5YA50sOF5PpSKUjkreBfeOjkCb49dx3PUDC53
wC8uTuDZO4X6iNtePOAgYrFHch2Noq/UL1zLkXhi1r53feAHgHEyniExHQ7+
q5qSYwP4aN1hjWt1OsqLp1B7lJ6y8VmFU8cQ0pqCrW0n21rLbCUvljMbc0XC
Yu2qXS/N/FCDgx5D9YR7B8LCQGYzaXMq5zN/0/zs+Zzu66djWI400tgYpShx
t3ByA/rWwQqR/qOeeWOWyJQpFn2JTZ1GzthUx5QGmhpftCgzxtN9QbgIzHdC
nVUr62wBQXOiuSR88U6rPgiNUrGKSJ2GLMRzVyqlzrTcsJh+zpKELHVMHx3M
4+AJa9bDezfA5B/5GeToy4ws3F8fU8ITI37uT6o1SV8mzfAEufRmN+G6aPcV
FkPISnXBH2Zm7tpTbPctuHx/UKn36EdgeQAvoGJSyfU40PjGl8RUOKXwtl0F
F5Hj85psT46iZEVtfyd29GQh3Xj/tA1A3Ov4zgDhozYL/AG0ByX57QQgMGpL
G3dD97eeA27hdxYYnVVPYngllUR4Sc+Ba+HCRtLocptPSYQXkA06DcUTz3gn
E+p7/Wni/zvlsD/qQ0jR1TtPHoQ2iocxxWnuJbXIldo4ODpzNOPYZwMUgueF
dltPG5FSR0nqa3mVC3OhFAubSY3f7KDKGUnXLnk3vPBCC6XXvNhcJ/z1Jcq1
L59vXBqlazI25VyeLZXMtXmA0puIZgaqeu6Q2PwPJEP+0n78ezhvf/j52KnZ
ApH02nEtJi2p6M0SC0KVwIwLlQW6+vXMiuo9PLAmHzc4ZS5PLxnjHZY3Cbec
wF6F1HHg3wUfOKC4V6yhPym2idYSBQCH1zjSMlObN0loliqx6wBIGSO5IU6m
vGbV3K0NCR8iBFHgh3xIo5azRBu6PhUBm4/bFbilEtgCH3h4e2nKRNVRFyij
F8r7b9BDzznvaaB4f7kWsww+CAQqe+BaiHRLqD+CfI/sdAO86cET6LkIi9sN
s/iF+zjGciy3DFCevTgsbEnk3DQ0l243S1jEylCKZS6uiltUSOeYZwiFMWe6
fi68dOXJ+nbPfoSQ3QReenVUq07xwuIPrndV6a4Stlcnpc0EHm1NQdEttfj1
6tdyt3Xbvb4GrXp1JDdQZ/CKawttN8nzesJg5HE6YBXyIffXbADor5uOJw3j
KPVnFUCPYmpuNrnd2xCzs6z/R5rOXYh6Kaj/ORbb450ExpZr68OlYoVOS/cE
eqXUjNLxtks8ObnwDLbAhG0/ttOw0YBQj+ijh+EsMQyeykY90Q4OODoYckLU
T8fB9k4KlO+j79osf8woC86j3ZEutn0jOE4ESmg4jiyg5fanxpPgl9IEnT5X
NL5vjssgOGMFavVVAObonSnPzObidkqfWxwnhe2js44reGrLtZ4RjHbNjcuz
jV9gO/EmpCbXtF1EXHFeaKA8Di5/q+A736fYzBWk3+wggdZARQzAOEgpLXwB
TnfmwS1cjoN0/8HxciKgRfO9qx5F8hj823ZQSdhkOyMRbOHS7LVoF1131Pne
S6H8EDBV5KJpUUFWRsXs0a12cv1bx1+KUvWLZXJYArc3DvtthTNc1ircXXtK
QaO0T535cEuNL3yKxZaoq9YXi9GIZDh9ocat+Q+IjUXBuST3Dagb6Aj73ThE
wCYDYzMZ9VSxFHAFTtfjpnaK2GadV+KE5uDFIvGqnPND64zWEcOdJALaPSJa
aRb2SDJuOHn0Xr60GU+MArFKwEVhkBzKpTdX9GJUWyA9eQz3SEEJrmMXEPGi
gxqR9c+GGnf+Os6jKXoNa2+HmddTB40Go3i0eksIv/rd16IfF2fkV2FOh5sd
g6xVnMqGFi0RPvYNYPvQC9OlVbq9ETe2SP9/pVS2E/QdpbHNQQoSGdiFfNSc
KPOqNhmZ/vh//bfXeAnGeV/CWf/VO0YpgFWashPhe20LJwkcwK0lzf6atEqh
UA9T98UOjtaqmt8Wrs6baCiI/3678zucOr4Joa9n8OEGHIqtoaG0vkfIQYNr
Pl184oiSdBudyDyI+B48UpcaqHtEB6b0nH5zLq4RJ4XPpqpg8TgqbzYbbmTb
m8U7ENQm4I1DbvYwV4h5W7R+qO/jEOkFaIYOxLDLrnPXVD2bJjKbvn3Te8Cv
yHTJwrtBg5FSMGwzp2PqwM0N6eJupv8LPgEGc8bFieXuc8JWJAtrMbwY3h5R
W6a5Ber4M8JglONJ0orT7TiKny8nYp6UKoJnE8wSLYVf0/O0lWP6jb5u6Lrj
TQKA5hS4LuDVWsYO86alRUaHNTRFHMUniGtAErk/1vLk48f7ix1mbKiZKpfg
fg9IiknVBsYrRnrPWPOrIszxxy1kgZJurEbH7hox7TYm8r1J5IWYK3XbRCtD
8KhIBtycaA3FF8LqIwQrVdRBU3/ZF3FFwuGc1VPX0IDpOWXAINV/GDpA792s
nrkniwHyS2N3VW3lQRolD1Na2rXUV8SLgn/aT1MMoIRvrI85I0rJwzvw0UBV
YJb1zdaxGD/o5NmjyPKgF6RPldRxmNlVzZv+lfFnuTcdQlvGuHi/SXWKHqeC
XtKqX5FEVhVh2d2NUjkapXWRHLLg81lRwh0m9tzfyTJ3Qm9EvhNDPRJmJWQo
CbK/CfkLnO0JdcGqgm00ECnmnQqpsiIFZ9PlYjYDrGzHQdclQ+5HQUkeRyZB
cNgqyCH06wn80rx+2yE73vuHkXvbAnD1p4jdlRn70A8zqqMsXKdS+dq9PwEg
v1HcPspLU/YnlYCpue5dG6zar06BKx0zuBCa7t8+AjouJMb/HvAXf68q2TzI
87wIEqCdRuaU7ExGAl8U8SapcxPeX/QWNlNWvQlbnjdwreAyl64pXb9D7COW
twnuUCs1w32kRTXpjZEEwYjs5l6sdJFTrC4EkiEbB9wgVLbe9VQoPj6Qm7jr
F+/BWwRHrz30+DasaUu3PUbxloSGRCsEHMeaa1iETjY2vIQKVKgDmXPg4a0b
TmqwNqRijAZyLJqz4j6++FOPizLwPowj5relR+STbn80YaCzI1W1rgu8/39z
V39+8+B26KI7OW5RzoYqXKeQXy1Ev5RhsWjNUqTYZ9TzKgUh3dWtIXwL1yHi
7WtsH07zMRxu3Ot4C2Pf8KOr/8Eb9BZsk8d9IyGLPFHjaI8UWAol9O3u9lH5
vdLqqJy0hQ9bYyerxmHsl0TDwYgOOXDSPmxhsTg2wagJjuCKT+Y6kaGFcwEC
7N/hrddGu1re9VdnukOFCt7YGKT9HRcDnCAmJJg9ir5PcIiEiz4Z84By+9JJ
jFw+5Ww1Tob/i7DOgKqBgqOqqmrjXP/dOnnq3cczGCHVVi4OCQSZhY5mtbNH
63RS7RZTnluoyxxYxeUmihflDWFkW2/Q+gWWIqWF+7O5EPvbGd2PcONVOCNa
+3wMAwtQSWR6aar2WiMb05kgvExTxOg72AaF2yjC2B61rwGK7TPA2DAb7w2r
5UimQPLIdkbNSH6775baiksU9qTF171pSlHr5Ng2l0kqNVze0GYbXJVN+fLO
MBx6DnUOCe53BteFRoC5BFdHxIxHOfEDKbXOPS8F5xzjGpwoEA8iRtz7dNUA
l0KcKwlsp7U+Dn4vuAJwHukmhyJOUfgrFgJJWD90H6ZmOMtp/C7QXGNJfYh8
XbM6W4HIToSK5DQuEm4KASUgSa+xnztt1hnLD/vP2X09lZkcQubzUGTBidj5
FzZYi29+bhfTQR0LONDj+M0e3Uq7w47nX6nGW3CUOA46ghth7qb7XqW761vM
rjiWI6HjNX1y801nIyGjxAKX8Hyb8ItZCcyH8WJmIp1pdqzc/Ka8QzWTxbVW
k2s5IgXMWrJTSAkw7DmX1dsvuZD4y9/+4QqpQwJi8XLPnQhSMFIX9Wu6i23n
DzgxRAFovyqfNb7DAzE56OXk4XdgImsog1dZWkAXFqBg0C+IdPbvOYV9KEmf
/Kt8KYPNzZXHDAKtciXn3lYpRRsgX1DcUn9XLSdyO61iFU74EKn3PPfqFUgQ
sddsjJRltbq1xNS7zG5H6VFz+U+ySn6VEVeYcBtzyfHxLkt0B1+F4ANC7VP0
WPD8l5mv6VX7isFDJTaWIfB0HpSZQuHE36FcFSSDsqSKlZOuzIkqI5eCdnO5
s2fA2Ufa2ZY/4rV2wp3Ay4G5U8af8Xhke73E62iCP8ftPh0mvq9EVql4PnJH
u7U0lewjimaRqONsmmNJiQ1PE0C9cJGAcP0YYU1YyyMYu4i1GPOHVlAiYYjr
C9A9omSKUh5FehMIszRq8CIRjLv4/y0gmUS8NNe1kFg4DINAR1bciEeiR8Hz
iuTuV04VukrX1LboGIDFyrKAh8449AYC9NZJQy5d4RtH+le33pHRvOZS7hqN
/tjosI9n3j3D/Czx2JghzNJxZQQlAkNf5Y84wYu8Pggpa3fQx71eg32G55Ua
jfc8PznkkW5YuQvH0BzfLv2qU0VvgJxINSuzcGbxYoDc4uvBNcP3Ph5lKeG0
YBifCzldW8a4SkAmSbs2+u5VOp1pq1Gw7NtNxyPaA/xKs8F9+TFJNcwOMJV7
x8rgIAR75W3GpBgVg7C161NRQr0ZlWGczvO8KG/VBaDz0a2/lXbok/XhPbZt
5/UGEDmOnN/kzkE1jVNlRljVaciPx/FP6ehOeOPhIfp40lTCoXmLtHrVIZmQ
yxBHJRpx9eq1VTIlmp1LrLjYS9uqUHRpv58DsiOfpU9je1qcF+OFc06fpQoG
MWrojz6S893vU5K/brB4XeyorgqubVFVPjsJiuwHujXNklr4slrKy/WCXpS0
WtQ0T7j0ikmXsdEDht+rrVaqANEdmRDiRCXDnqhbPStCtODHoaUW2MLZIZrj
SLdySxUt9tlQ1JQCZmdxoN+Fa57qIpaUWlQSX49fL3ECeYdybaoiIkmc95rr
T+Qk9dxtwQs7aZ1AxRIlfWR6u+GUWnILy2ilRUcBvlD5Jwyr26brISkvBH2+
ZoFgqZhS7vjkOFzEDS2ekXNE78gtsYM7F44cCPyg2c3oYwxyCb3cF6flQJD4
zDsM4TSwDgSZi2rLubv4ZUUHv0rttMw9Ypey0YSjbO45xxO9+bMwnVSGiDe6
YRbAQ31JD/1jAFOKlbDSi6tA07qFO/MsLaI6HZ3X6csAWD5lWX9AWIEG+Ube
Y2rvqegxrZFqj9HxJDOMJD7b/44/8xLLUFAifdPsjTMAlh20rrz6lmridl8K
waxacY7rDxux2zNn9ztm9n4Fsm29Sud5OfoV+ZveAMvB3euTy8UI1I5NoX9d
9PfnMzCifxdQtAla3wHpQA4bKJv1fdo76KJNdKyDTv4vy7eq7/MtouP6PrF5
JJIp8NhCFyyQ7VJHqcgMy285xzUwJg9sg1qisl6eu9A8gHSkcmX5sGdQvql7
EDhd+CYw1rUJ3+IZOZGhV6hItS32IJqqJHjJiikbIgrbRUGZN2v153Qkv/jD
6JyQuAsOYn6fBa+ODcZ29M7o8kz4oncTyUmnYka5djmRJuBf3F/O+qZSDfdH
mmq8UiM6SWmx3C7OlF9KVRquHzBZ1biM8FqMgD/AZPF7CqlA4AkciYPJ27vq
hDhYYgyE/30YTWga5pXG/+5AtLS0vV6ZDlc2s52PJp2peFMiQ3cwTtun9nu6
O2gUNNq3/Qxgw57vGLI1KWarmp+2vOw1azYVkNORDxJbtA9bN9tnuNS8SlAX
fuJGIXdqVDtKlb4+hNW+9VUia3Bnvn8iHign6iGHQtzKQ/pk+rON+rDJrhyF
j8zVpATzWJOcB9Eo6WJJP5oq27Gjba6Nwddv0k1nK/N34IOxTIwUDFfJFRHV
XrMR5nHAwLYvS+SfbUxt+1MRfJNSw1BsGWFfwOEOncLfOl0g0GyLYHrDWV60
NMV8Dl3XaJdeluD3DRJhZBRBMYHi7mlg+gzNqlTbcAxd1wKjx9p6elUiP3sh
jPcxgEHNTqzFfPyxk8yL04SGFj5vTwQoy1zDjyeywtQVOQXSLTDAxhpbcjL6
wgkKOrElkrGHLgwpi//jsWa76OmpsnU2JZhnY711wl3UL26E6Y5ov3Quohs2
ZkDu1Y+G4W+1pCkRHTXCWNFOYaJ6rGSsmMHb85+ogwH0Lhq/gBLRHbSyyaAm
qZ54ysmqcJl/WrhIi7rvqwyj05qUMBCTQNPUFEGqYHIikUIwbingv4NJGwy3
ruJBPUYeVKIdaMYhb0npvkKO9k2Orio25ATHB1INrEnrkVYeFLW73jsfI2os
pkpopgyEXhvfZwDL7YoKd7KGrX12LSni+lzGA1ndU2TdwZ6azzbPRtsJycuD
xtRQ6eELXKuZ6JnYm3yol1NJiP8JRlD+ih0ch1c/gvFNxtRr1qzKQNnDRtCd
DinvrH42qliVVYHFmA1SctzWOYMmGKPXmWOgB/Jr6V9rj7kQNV48AA9kxYdA
7sqGSXnArCY1O2GqV8bV7MlJTeYZce9uFnrTSj8vu2PNPhOe5HhcvcrR2Wzb
lHtlJk3vsZ2FMxzoqfwfCphdlTq/9E+iAWQj4FRsbFpl2oURTLepVghHZQ3W
TfQVD12iyL2hUOhXbMPmgpAERQvqABn80AuZj/wWcBwaNnxp9UOhZ5eXML9R
uz6akHtBeaSrwEbyBD4PwN7OqTowm6S5+W1fzLF12iz3Bx1YYhm1P3J4F+9L
sGt1wa9M6/rkO251P1mM7Q4d2ek1WBcBLGpKyHX5Aku4HbwJBnH8wHq/jcP+
poJSACjjZSN3tVcHV6DQ3CDjMkAkkWYQcedDITsV/oeTSCrdZ3Iolg8qXOgt
84DyCWkVGptTsmYkD2J882nwkkAM0X7iPNaK96YlRecLjzew2mJ0gdCsLkhJ
7yz/22m7XVjOpN5bTASiopo1Iw+uSpB8V02fErV2PiN1UdTig+pbugEs++Q/
S0m396h8WIHmAf1aSkQm0bDdpnt58AetXaxmcv2cY2GqN0maZsG5y3m9FSY+
9QZr/tYvwB1NIvwd1WB3+gcAx2w7foKxicdru4oWSkSha8Pv3GEALf7ypiso
gz1Y4ViwU4QPdGKtWW08bboKbWGMiTLbmCZXLtbNRCb4eIYD2ZtPQsQkEk0Q
ZVskqvsJNfGQfNpGZGca4OkqCAkGz7cMygsKs+wABrd36v8kmke7GJP8m6KJ
pOQtoQgCI8fTtFjX9Gt4pg7D7w4p5daCMLBXl76zg7hg+oQcLC8IYDieDpIs
Y9yKXchoZyJfZfac8pGdTuL0t+6bsbaVM+KDFclzLZ7bcS/apiBzN6d0LMUL
CeGK9wb/Ch4j/spekP5P41y1BMX/G77Svu4Qqa0cvphnR/yf/+5ukFqkaI10
rNFSGU5LBKm5Z3PkpjG/2aQtbz0F+ubL6l7vDIG4dtKBQI4NZSvJn/LskH9l
BxtsfMd96d0fgB1vkDeM5j8wRZmkoHnpFjeG/5e1HCVJ7Vgv/KAVVG8T1kPz
iMgeV+SGwDYnl/ccP4LL/UUPxT9cV69sWO8An3loxnpx5BnSDUIv+o5IQkDN
hSa2Qk7oRd+mqthkKuEqXaHTlkI51cOwYcs1bZIEXlsTT8KSBMnRDKkbtn6J
+83Kh0x2u+3ip/GHvnQy1cVETTjpEjLeGWTGgHAnAuRqcqOBtlwQ8RDEbDZi
jfkFHJNQNANYa8sa/gNULQ0Am5JvRui0/3Qfc/A6pNGQvnuI4xcztPBQsb0u
0iXUv2I28Hu1KkZHZIlltouevtH3obwuud/HNuUBFPFrbBMZN3jbyTpoOoC7
WId7H3Wmz0slzS6fKv2aM1v+z347EEz6MJmhoHytEcfDhDnmfuoYh6zOIV7C
jYFic73FXa8ntSCQb+e5wYuRKZg4wx9dL3JiBTKujzDv4ykED/ZgFJkTwGHE
tJQKaTBLRt0g3n4ttjkZ+noJgCRskEN3x28VUUWFJ9X94SUe6UG4jna/48Rt
8QrnMvYfPybIyjSO9WyppKKB5iw5d3nNJIBgIECIWekNF1mjaOoN5CHSYWjW
3gVvWgkFOcOFCBd7Fe+QVAfG98UVJEpXS84Sz1GS1xIhnHn8TJR/uc+X0cYj
i2k1wR12ZLhP8g5AttsO8Fp9NjcNKQrfxNV1pG0cPMShtycZi9ZaMJkBdUfg
0ODF4boFoXTrVHh2WJS+JM6ZZhCVGPYTCuYwOnW/ts7QTCqrG95Jn7Jr0uaU
+z8IOGRDlQHjW2pLA7LsezyBGEpQFwrYU9/WHZkWWB1vvaT+pOk/ennEdJMk
13RMDfkkemE+fGp6XqzC3pkI6LdvzHZKjwOEFwz66/16GxJr5s6Iqr+AOJ8h
zQ8yWT5u/qJEbKeR+pTrR0GPqTGr+0OVrV9J89HCX/zlyD3kxK+BbNSJQXrn
2Hzd+9k/nnUp5lENbP5oDJ2wLS9WeFus4hVWiqbCRSh9QV0SQm7/5RxGafeT
lVkfEUSfKAmeFKG/DFa4sqDunw2R/jhpOUodTbkmfPYvhBoE3Bn3Zj0DL+Rb
DWVx+2keE0lJFc0tDGN/76XV3hCPbBkKcufriQa3xq/V49MvDTQ6d9otF2ME
BgIPxRvnrpxGIL0a6ZPB9Nu2DthItKIxa0OQ7vghL4P+6b0SADlGXev0OQv7
/6wym5xEt3+qBfQLRzu8lXtyOhmdoRqFtNG+r7cc6oKZTY6CqzU5oBtM3K7T
MVWObWKy9T8p2fNYkm3WI57y6iRcFJorBHGByIhUfmbsjkmqnUWQnTflNNN9
/qo5VtUZoIvuaAwoCVzZC6680z7Lfap1YDX/B5qLcTwVbszTknGpZgaQBIe5
nBB0bdF3k8WmQN5nBksibyfGe52vlIw5pU/3pYicLYaQSdxqRKnwiWNzyWao
yWH7t/IuhvF5Ng/221Z5VNPfo08LjU5oMRU2xee9nP5c64O+p3mP2vC6mVYl
hg7i+eRXoqkJiTG+kIMnEHNVeEhEvp/vCvfE6+YJmMp9abpCfsLzpHbC3gAs
Wnt03mNTH+oOY+p1DP0DspeMfCNJXYkmIGF/mzmFBw3QnI53oD58OhsABNCJ
H+bTDBlMaHuTvPkk5vmHCSULU7JLbXNf1IGBM+Sr1uO4wAK9NEElN43kVjRe
7cRvuqH7q5ntt8Ah5PeljW+REEj1XBeKWGM87X2yi6IAQzrzpgKIsuPlquTc
qVRYY6H7r3LZWQf/2ySVwHseAmr8+UTVe7QMEELCRwhRyBtjn3Jzu2T6OA0E
ejUZmmzSKJ68AOkNcd/+K35Hw4O5sSMvff8l9ulx3/TYVsMnHp+aEY0GGimm
CX7SkPeRa+xcDH1GK52feVpFlPZaAuaSrNBBwXI9CWh+zW2gn/wWed1BMg4v
3uwHODduCkjVF8gJfsVsjsXaFdNvX3eZuimDJIbeUsnfX5H9DpDX09cQ93Ln
fkvS3uPjrdjHPiuXG9SLcPICM+f0d7NgHxO4r2JW8ICTWgSxvvQ4NR+V5m91
pZWRqxHCH6Vj1EabWoBa4EOJIB78NF4y9vKZ4fc+kZmYweqGYCyPKf2pak8t
ovtSzG1BHlqUA4Z2363WJQ/bx6fPX1IkDg5zpvnYeKh2xtP8C6r1tA4wH0Rj
U5+s/gFhj/yiob9awtWa34NhtoGHbERWavWGUucIrmaKxOMuQn2hZH2FKxQT
xs6eV09HvGoCHMIoXS7/i58xcNH5AorZIqIn1y3DfA88DDqLS33GuwSUcRLD
24tXHktXF5lcP42uZ4fBUeXlpWBb+5UTcH4izYyg8oeV2RR7RKhgR97bgRNN
Mq2pCvPGE0wKpeO0cTnXH8vqJyVX96p2ma/k6CptC/x3T2S7Ox5ndUj39O16
x6lb6Ie6Btg1KWLOSWrJWCw/3mGxoE8n9TlOd3WO64jMnnAfjn5AFH0dKYs5
7MY2NMJ+tNV0W/o8AJlm+pYxhEnmRWsM8iOsB4g7c6SvTgbEmEJjLKodRiD2
x0wiTIyzr/ECqNfECYD75wpwJ67jNle9v1iYrnasMSt7juCZgwLLixLHa7fY
9+68+gJtFH3HOdhm4L9Kn5PTrRoxxORthtiDbdDFALqTpQCnA0CRe3vQm1+B
nszMaRrn/IPoZgB3A80ajXMAdC3eJvpXSx/eG6HP97x3GEi2ThtEiATqN+MB
Ur2NTFWr63HyHgcydKyzjlIquFUENwK+nyJD16UBbFZTB3kJLP5X+Kk2r4rD
bztOYsyG3u5aqR8cJD6by8J3hlxjVLtzy8bRgjRVe1Xlru6Ig+feGzNB2M61
bCy2bzcYwU/BNO+Hl70steD3ElU5XIACtAQOF0PGdPLSprWJtgP3secOhu4a
gsHcOlFa/QECU0b8s+sBvJumtPvn1TdF6tWiteH5GNcUDCvdhtjbXviGM+pI
kVKomL4KxyEdp7bm/RunW8e+VC2IPvwyXIlTxF/T6VuJNbxQJE3u7zqJAWkY
HWybjUKLpovpRFP19Xpd/AYNwKq0SzYgPSpP0JTYzwUPOCM32RPj5o2V1krt
KqZuiy2bplcT9Mf60hINk1gcy+Fij74MeqCUjDvi30BQ6U0vMsU/JIkHiR1T
L9jGeAfvtG2uDMbaBqyru482EyFYu6SS0oWV6Ey+5dcVbxAOiKxZQMfBNVxU
HDrY8zzzHaxSWVyECCtcB3HqFriY9A/2bRP3cA2b2qmFH7dLT8DVbJ62+ABT
Fz+cAtPAmE5OLHEcgvzZm31EoCB9HuvjBhZKsUEqIC/WV2DEFSzuSyr65L/3
wsDDOszIRM/JL8MWCoOiIkEMSqmTKqaqz+ioz3VTloBAzFsTugzEGYezx4ep
Naso7M61TF1fiT2NCslKwrJ99GIZ/8wcZQ/p9f3SL+CixQcmAhG/Wb9vv2wa
UFq2IEw6Ft+Cn+5ZMP3XGocKXMcCyyPjcGdp/lGhrSibsrJ1YG3/4mh/ZmUS
0eQGxGrfrHYBb+q+JuPEL4AIGoR77LFZZ6ov7ruPSMrI94SplFNmj3HFJ4YH
ArdLp27HeDeVOMLlY9W6/1n2+v2mwyecWqTr6koNoDkkTjlnigryHXiRDQjr
7Yzbkywa5ueMwynPtkLeunSMN7sgtljNTNByuuPIF4fSgcflQMVGz8Vjiw6M
kHvqh3h6aTyU+Bcgv36Se2iQ0gy0xmev371VeZBjmOSDDXelzHDIUaDzDjhK
zC6/NWfhPjFVrU9cIhhXqTb6LX/v7zNriJAx0pPsuA552N4oXgdKnGpHcFcT
YayRgUr2ObHRmnOw/7/4cHG3qSRQ6RA9O+T3/RqpTJrto17tymgxFVojyPQi
uS8XoIl6uF1iWrNmmGskbFeHgcRBTQeI3/QnOVwhI9l3soIksrqY4kfgvQjx
9Kta4VIdLk8NbmtneBYtxldclhhh7YBuBH1TgVFnxrSxxed4yHA7aI2Pcc6T
SG7H7TkSvVq3Px+9ljHi6pAAGBcW8BdHemJrcseWzuRKNDxLpnrwHCf+oSWK
4hFmUArkBJSpS34yZat3CjzaDmV1qUF2ZnAZVobprtQL+B4uv8jIoSZMyG3H
dUIxoRefN19P0jwSHnnkgM/Yoc+ZfpU7X6HaWUUOlGCMlM6r3b8EEQsVwL6r
G4dDZOzbRDDmEPcIpxyS+l42qFkpfqBMAxM30bABwJydXJJP7xEggwL6QECa
K9VQ4bYTxjdpVzaWpcA+RYAifQxABqkX9mCsaBtu7+jhoJHxaoICLlpqeCa2
3nXYh6sO8no0L6EZXphwL06xWUfqzQ1RzrrZJOKGA+dHllMOAys5nzoIzhhD
Pac/521fxT5fuIj1QCB9Uy3qtuKJv7zWbTzwHTGLoQsHArNYlp4ZeMF74ipZ
Dig3Tn2nqQesvB4VOTkENkChEoltfU9baO2/S7Mv69OYp1TEOAUJuHaxUFxA
XIs0TRdi1oPlisu692ooAsF6nycBRoqpVNryu48O258nM9OKNzD4f8vcNI+j
PC6u25HjyXUmUilbDG8wGZHWkpIGAUGjHXqdk5qEM8A0I6tx29ISpv84NumI
Y5HdtsfeLQI9miPOSBSHia94tWdCUybnPlojn5Ex3Yhok2cH5smriNSp56jv
KYVzXBMDew1mo5Br83NOlaFIcicdhQdcoSF4tPSV8lGlmVsQzSy2n74NulGP
+Fqvz4K3zg560WQ7MXMU1hxonjlA7rEd/dahhaD60wk1bn1E1Ubaxna1Rn5b
8jlfXFdMaS6muXmAcTKAwvnXGVTbs6SccrUYNNgumxFXwn4Jkl1NMcOQFYTi
7L8Pt7eO8QRc0ZEFdatYESyLDA/E06LdHaquUN4r6V1QVraMrUFta1zn/a2n
nYjGiaHu9xHso/veevFadlVIQqSeYv26gc7RoiV2jvd9Ryk0S1RJpinjq7fO
3bIz/kEgQbTaB6n2guYuGs1WcS/qd8FYI86u6YDO4cALyeT4Rw/LvSFhkgh7
/iJCFW2qCnYBnut4oWutV+iDDy9FgGuiT+eeFPDGB57/lNHPzwMRQQsovWib
vycTRl25vHapw1klOw14IURc7jdMUJryrUTBQeo/6yW6IMVdl5vMttiUl06P
pArvOhUbpIHUsVWmQCy6dYdDLFV0F+/a3G5JzC9FiTEOaGGzjox8TXVHsGzm
xtKhj4ZggpflHFK3t1h5isXwLpUCP/RmRkVnvUkG4k8hbnr7D16zHMP7uscW
pVYt0hNBOw/mN6hPTiiF61bySWZWMCdqY7kqFxevj07RtYAtuEqP6gjaxxYo
VFkY2RLeDFc8nB1JnUCbsCYAuoL3UkOIIVBw3Gu59sFny7/xKBuTlizvBkDA
D79MnVE20AG3IlM29E6HUd3SE6zVRNOG2qDGcSRqhPc7g9kGxJRWCjtuDmx4
QwKrrzl+xgd5BbRKUmQoMoI78VNoc6qa3tyDrHMjWiYzK80S2eOjkOC0QKBJ
Fl6yLQLcoiC6KlZllnX1B57N8VH9vyc8XR2A/umw47d/EM7AzGnPmImL9mSg
L8ydL3IfPTEtie4CsGJ8j17obhtv05yrsRCFqwr8SNgsC5dwGjFp2oSaqTn/
Iyrd2+74WWchSeaxTbNnJ3XBvcRH1C5uICYYDGQ/swsCajJ33+FCr4brc8/e
Jn6ze/dOZKSGb09e7CnHd9mV35dXn0p5G79DQAOC8W/QdgBnYYFl4adtf7Zx
A2977NEGY+gfSDF7/LlrPye2DaeOUEDi9/lxqoL/1wFprHr1FnCSU5XZL8pb
SjKLFCkpxw+J/bdwwFXBWoBXtGjh8/2V68zKHYs606/O0aG77YOW66ufoTQ/
mtNbf/9EFqrg0JBVo80sW564/CBqH/AB1f6Wk1Ae7N6g/s4p4pg+JxgBYmn0
UJoMDPnBgwJAtn0lups9XMn6lAsn1/DGmpvxBP+Odw92La97pOhnaB0X0k/N
LQy5oca6fRQ1oIPHePfE0KRR6RfgUX8Evdng1gYZ4K5jRIKH19XccP1Zj+zo
nT7qbRjYlekCxVkFDJfKUqVQFifGk2DVpQvGWQv1dq1sQL1Q3nGqZVeml9pQ
2ACp3opGBh7BQdFG6iRFE9u77bK92KxFrbHCWQlkF7KuBJCDd/9GgQn+G6Eg
YG+xxOSIjwLhDr2svltiyYGCU56pi+VnHjYFOQ3aRuOP5q3raFJGiZYwhV0V
+fEgjf5NU19EN/xt70GPoyBy7Qv4/7QkYgJtY1FmpI0Kof5RVYZ9JvwU1LBy
yL/eabW3Fg/ZKT+OwD6QMbJSc7hM6wIfQEo+b/mtjvr9JmbubgN7gHDd97Rg
l4GMEqhPvqrD/pQ/8NcZIj5MAS0IZQjf4kk7qPtvz4q32WUThREtIcSkiMaa
mQ2NeHR3Dym5ve3XoxLFtscVZeTxs8BFOiwFPUD2z1pGdIA1cHNZFTEQdU+m
K5HxmG74Q1QqGHKIQrtxszx9HpZF4Da9WGVB86MjyK1tEwvCcAG4T7Y3F3tP
6SiNG39GTIX847u+Ko47NMjw4CkF27R7djfGlWsgZI/h++Rehvqr9yWKZ0vW
zjfvR31N4nGS0KOLuXKVl4ALLRxUy3pBafpdixLIMqyE8E0YL0tBhdFMGzzZ
RJjdiGiWtw+2JYHMYuW2e5Ezmn4ssNaZLYWegyJPUvzJynIXZJZjOqeIj6+c
1WEl8mdD4Tu7eT8OSU3CML7GIcq+IMtw/4WCs4YWhbtwVvDBKrzERCVAmP2j
TmeGjJ37+ml7vWQOGAYH+rGnpGVtdjqiy7Q0SXRSoRaK5qStiAJVlOaypT4g
c1AKpwG0wXmq51orHUvv4zVyeqzynsWQA4jSWIw/ozu4onWzsb4+f5Ag+LPc
EmF19M0r0VvGRHwdkcETpOjeb3hUlwJiLiLmJKq/HxHrYwXG5do9dWTQiq5W
J3uIVqPuxP56VXf4cnZaK95oPQpA/4m1oQ8aSXOlUxdSvUrw6If6rLP6zMZH
FS9u+Y1JvG3Z5tLItdRHYqYHi26aJLDiXFRaNy0dBwbVhOzfGztyogzruYTu
DWO8LFsBrlDb7xE9ZXS/Jcqq/tfYTzJePQShKCTXb0Ye7iQ80Dzm+LWLruRX
w2KpQzAMaCfggMfsAffYWOgPxCw/1PgTuoDHAZlctArAboXoRl4f6jVo3NRa
Il0zW4vKWDclcdOo8C97k3Ae+JRKFAfqF0Bhzv9JjWEcmuzh8Cjous9CmDMA
WtWGO0GhfOrbNlLqwe6Ta1aNimDGm35Xuk3f8/J0kYGboHq49nuQH9S5supu
T7/3JNirZAh1hIUmKftH+DgZDsofulAZuV3TUMQD0OA94TW+7aGAnRpkbPjC
en9Th4MzjknHJisrRM96AujpsAk2oHpVejbmcHUGmmjKm8m0VI0SOM6y7TqU
cadEHHAcX9gyjXXkJnD7MR9GJfekCs8xiMjFg/kPez/Kfl+jToRimSoLaIO9
oGdNzLbSyostrna1NZurCftluD92BW0wdSuTAxo8yWe37zKbNoNEiQtbGGCC
nT/1E11dgfgCCTuv/cDJLlWsaZJshHOUfRsjw66zpoZusntWFmle6MA90z24
8NMYgZ/4eSVDRgahQIXckhhC9MQqOx8PoV8klbb1V1l5OAROfu9vRVIGue22
JlZIM0LhtD0tlpiS5sQkDtwqtXqpxBDlPuwQlWHydpKJJPSpyaGjhF75QaHk
V2kxPd18u15mi3+CqYkNo5nwqc1rWW1/SkHqcxGMsEIughuUTriwLMe7EcqF
SKqVrj3kvbT5Z4vQjsUSDUKH6qsqjWeqk2qP5wPA6BhcqE8ncZB5Ptu1/9nd
nmtGyewapekBes2RlVwGISYcDxMSBklvBvXBwNDo/m5e615ME/AeUMXi1rWM
XQDv6J6fh/TEjeCGsUgcTEnGuhODfR4F49zjO6GmaU+0a12cPuNm5f2u+LJ6
+r4Mp8WzuHqFzee/qnkbMz+kWBwAF8Op3yn064wnW0UJor9UjpJrPMyuKy5B
yfpd1cuFCKMaIB/LLwHJLbd6bN3G9teWGmblxoiAM3bR7exgxgGq8sIu41/Z
7yBbRgg+9MGEBXABMdojksx02qGWW9gvLnvzseO2ssFp1XUgHIxu5pPL46SD
FfJrtWM4eV6ennBP75kfwFGHw8oIXNaisYGw35V8US/UDHPhhiuFa9Pxb4gw
XVJocNahBjl0dFbUby7mHUSfh3LaIDS1nDPBLgLcztoCcC6Pob1YB3/RSXki
SxJhLPdCjzWfhdR5m/v+NK35c5ACYq/+NX9eKcfQTxcZRavElN1WNWjy+XUW
UV537jhAdK7ziV+TlQJ0zGD0JVA/z+2nRyWB9aoCbFBcXf9nhVyL36jzq81c
GNZaPfkY03ZtzlkvS8CyHm3UVTng0FMhhVZkGUiDPJsPTrnkeqPQ3SjlopnA
2KiBNB2Aok+c4HGzs2PR0zMQWXTxARlnQf0NJF5/EFi6u1hCAXlSS/v+Be0R
HvzElD04UVwdykXGwbyBA4+JJfepxQlbRMLsfPtrp2je3hPvrFWCO6ZCZtYv
X5y1qULRO8LR7+/RsY8vV08bb4kBEmmtukIDASfBcQaMJYRkmQgl0VpELZSl
aQo4vbmH9le3XowCE/iNioPPDD9asIMMCIhKrP2FBrOTtygkBZE1Pb7OXeZ3
z1ShkHsrzsHxrYO41rYi32KafT2EppntkKjjr5XVXM31Y7/fHYNWyHwamqa6
190pMCzVZGD3b4BdWa91qt6xhYZBhk85ZZWs7O9Z74VQB6zBX+84amcciKKQ
Kfh3AXmrYVQ+izJpfVRV0K/Ut4GqD6ADbjfvv3D2umoiCZ30SPobRSNkNyrP
KuhNkuBniKAWhdOg6dLBxL+2yY6FMkxoADnn2Hj5LIYdNiJNkMqBHD6ZDXjA
1bMnFybwyS1P6DJLOfSbI6KPTpA5DDKocXSvDzrDntJkLNINJmh6W1ex5Zmx
tsTXf+hS/DTTZpduhvEaXjYpONWGyoA4YQzc4qGcSahkz01LOAmnH6uidf8S
6gOIrpaWYh1jlM8F4l0GY2CP4Er0km9tixVA+jCGYWE+r9LjTek1yUtTBZDg
dMIz8Ahs4NX4pIeEW3+AYqIWxeukcpH0+ZF7BQlhG1xBEuAPtnCGO1lDo8xs
MO8Ns6oEBHQs0CWn/OnOG8r0ultxzdvfGs0msa8XBkTPOnxPf90RgQk8eq1D
l5vn7qFpvcmva8Dq2o8CGvrR8bUZs9bbPf+jtPfBgDzZ1ghFW1hmh9OKrZCi
rjSPXZY7Bea33bkYmQ1o+8M2C2Ws1DiYUE0yhK4bXa2TSbthtk1+y1oEUsbE
AGwA4StHTiYAtzjyE1Uqq+YUE6wzx2S3H5NSm+ZFBXgNRtUDl2WGT4o4vv13
F7jSTHOb6M+9WK0tkVtwDN4b9V+2CvdBRMV3yap/BAy/pvZ2HsNLRf/ukYHb
J1fui1C8doACpWKOV+BIeUZbMaHgVP1FEE5AC0GQfuod53vdRc6v7zai4Lpa
EsVib7aLpoLAR13bUqPPtEqFCMtUYcFeiwKC3yk2EPAUkDHc0xowyZfpX2C5
hf7T7KUDIlYvmCTDyEsiIuHKvcZPl33KnBA8eGzFe8JwDu6qLy86BLOuuBNg
H/o01nt9HgM2qPJHU2+D2jY+hglhxwrRgLqW5jQx4D7NmZJYzMDLFntV2Fps
vIhECVGEGgM3VMYxQuaOa+vUaugg+9JxQQFzEacoqhRkZq7j6ayWD2zRldX2
VyOey6Egj/NWM8qxZmLDiZnfY8fD7CVjwiaVKbtfI99OKRnKMLJoPjDvfKZL
hk/gwBKchFpfpnOKwUvKeWGDw0LnWhgNhBQVD14iTCZRljL+eGofMROmEMw6
s6ENfmlpvddlh21qLTXP7KyKS4CoGLSIj4uCRtzpjbc2H08kt9SbLgAd6ZGi
vN7gNx5LuSJhvjhLAi+vpw55hvngVPo5PYV7jfnslxZPr8nQ8pZ+dNbbkQCF
J/Yk02bzBn4CfApJtuMqQd7yJOUh2DKAp2q+qeAOk5AgnC/Bv8NPwE/BEktk
+kXR+YY4nEH73ecSOWU2B+EWBnJw6FDo7bdHBISwVFdyAcRAAJQy7eKCrTJS
8BWqz/rLukzygBvtQtoYn4QsbdlEUFN9V/kxIYjd3oDwp8WLg79H0fySPtEE
dTaJiF3L7AB/DglqCAiBLBcCCYSFea6RQeQq7ACUc5ZMuYvEPNNArYfhX/PC
PC5bII6ycyWV/K+YVyUU38KLLrLCIJrHm9Orzrs/hhNXwBd4bELhh+QtLvx0
lByg0foxBelVCfgx58mFKG94R/qj7FeYmuMJKaH51OLscmUeAP8iq6LAl1ju
oxAXK+hL4EMGSnqr5/4qgMKpy6a0VfnAYIdAS2TZeuvwXLStWjImb1EN/vtS
18z6dKa3GFVxGExBS+tJ4MfJsuWsLp1hIrYe3IQFzJUIg5uACpSsn9LZM0ml
zzFrkACgkrH6uiE6P8jsRF6esCw+VhtcXxfLT1HtXsphMJE5EbHm/YSJqQtb
t1+40D80iwHICVLRil+bRzjm4LLVmAh9wk9FRAuB426u1uFHcCr87gRN3qlY
jsRHAFEm41cyIKpivb2s5JtvalaYZA8bMCyyGXTwauLC/YlEQ2MqoPjKYrmj
9mgZBKFusRvgiVM251gwl+h+/lIVPy4mwefSSU2q+7Qo2Dz/+DfW/4jGRw4S
CTyf9KmpLQT9WUXdxr6lE4ym0cUSEE1qHQ5UYTh9RuqyVsSA+ew7YsW2GRse
rpCGyMpsTzUszeCrLK3QTWzp+nHSienAeGb4Fuv2X9NCd4Vd8cZUMIxItrqr
hMXQOxUoCMpWCumQnYVpE/2z1DAs3EC3cj+d1/RiP1ndT1CD5csM1zzMOYNM
bi29AZKXvXYNa/ca458pFvTJJrs/qO+BW4pBDlgmGRE5aedW6CBJbXGjf5JG
4cOIs03um1mBJ+/5bRJ85fU56Gwn6uUmbV9Z3JNttlAhWaoGd2jmrjVATuaF
8uoYktvW139imsHxwpAJ/0ViXVj0X1KPaukvcHq/LoHc00CX+CzsXo3tyiix
4teHqoMy6KfYGk0E7KeSDtuvZl6sckjguIzAZ+B2XMRP/DGeioKKpFEmLv/6
KHYOPoG+b86ZOJcCEkTbB1zgb7UuXM8ASyIfB2M5tjMRkyYdANZUZiHQM4Ha
DhSuSpzlDsvoubUxDSWik00UKRbhnoOvMq8poUE0DBXMIQ7UfEjNzf078AME
UC28JKaygYesiWtbm2pfIzi8DQaJri7vlbZIAKYQqUwIFAi2LRc2RGPN2qLT
qd+JMbLz9eKy+jZk6AdWXDGFZBOxYnStVOJqRDE18QxYZ0RZVJdngDaEOrX7
uSBV5HdFXo+is6V9uMCvogCIcYqwrLet/jj/Z0WP+VY1RZtIkWkFO+eg0hve
3+LyBPNxXOOAATH3VD27Czc6LYMFNv8JSbatfsMlcNOlkbUGANiqdv1aeLxc
Zjggm4XfR1RGDkRUEoxZ1rNptrWHBv99+CUD5TjwRoSsjAUSx3huuiuoRxNr
9WfGHowMLIRWCvKXGUhMtQt/K1ozecbxiUgpuHfdyIoqquCFrQg/O8ngY0iY
WxL14aPjpl505fTHsrNljOP2AsLHDFdbapE9U3ZfJ1eGRHlJiq1YwJBdPudk
4iASYLYFTavn0KOrzcpU/8BvB9bqSGAxJl8Ol/nX2PmfdC4VR66FiFQ/iJez
K68yOiksT67AD00tLo+wu/0DHGZAQ1aw/t7GOKmWPGUqtvgmM4AifCGh/df9
w68rGuoP5nRJ9MU+KAlEo5IZt5wnPT98hPplu/I+KL/bJNaLzIS+FNN6nHlt
g4bdQzoyS0gg/JUYoXdDUgFdrxRJafLnThMMtdxKlpo6FZ8vRir8XuYhrtkV
ydXBxnhFnNkDfpzocf8FE7pd3+RG/Qb5u6BfSbS2CD15H0eVtpWjrz+/V9hG
AwHvQwWVHEuepE6R2B+q9D6eHqCWHPhWcYXnyr6gcKM9sRE4MO/tZHW2H9+U
Z3XR+IcN4K/NAdyp8XLxr7nQy/kEkEexylmCE+bjpPYVTfo+vkEdiQlHZO4A
/XKZdfackrMTrZHOcCHi6APm+86Pgz3kp/pa9WgjSDmFypHSyg/cn4dCeN+2
8gNO6JmZ+MFoIrBWBWrnBrYen5y1ag6rQNzOqmuFv7Yrj1iqB3/OBfvdKM6L
2rOCV0JPPlkxEC7+GUNunSzP8eEVripbpb56WC6gKVuBUnnRYhm2QTqfPAW8
AZzWwIkP76D2DMlKFz3LfQv0Htm3gYsURwPyAEuxWMbasARCDcwuRLqaABWy
xhb70zR4ZHNbbEEzvNfb0Yn+i511terN1U7dlIxO8+xG7U+JTDQJa95KoBhD
76gTBYiwsjPf8MZfD5HZNtd+IqBbnlrjKppwx1rQMcrdNr59UAcNbTlpmCS3
qLlxQ1ptbcvRgogZhK7kwwyV/gJEZluD4ERUAV8bNUY79f32e0ayTRCjm0OI
ZXiUfBy7f5LvsaHEsrRkF8a/BqIaQuvu6Obh3wLIfMeAJ58Ka+xZaeHhq2pH
qswFkec6AyRLVdxpanlsB2gXxpvct95SuCO6+kK8s3Bup0gvSOHBWfrekFOR
buOPHzRqPztmWEQBTKYBTJ0vrF0afgJs/u2Mnjx6k5aHRQ7ov+BEIgkDnXHp
whZHl3T19jxmcaVBg8nILbNfc9bhkvR3wtXOBsUqs0VLUpT4pTI0BWgnftHH
QjcBZxd5ZP/LBsQdmxsqh6VJFgTvqf3xYorK8s8qc1chCjYcvkDlX2BbNq19
tuH7okadviEV/U4Pm20lRVZkDeiopGh1BsdhBb9zq8Fq1FoIVIfTzHcaK1cH
klNthbj7UPT5F1pDeYe8YsdJ78VthYHbnoOtOKZ6e1anmZWtTHnPOnsUt6ta
wHYtHENsCW3YKG88Aq7tH6b7SvrzFC6L8cPDb6VWpls7RIBb7Aiojqk+hZ+v
THN6dNuWxBYHzRX3MAT3qDTyDUOu0BTpN1AQAosB30De9HJPSOv2LbmKE4nu
UZ/RYTsyxMSsNcf5SnLQ0/25a54omvPUC8XXRjwCOQ5jF2n7Kn9TA//pP07N
POIclcy9SJfBdnuCMMqbRhCuqm3uMnAdHu5KhYlrOdbQNAh3UIp8R5sCnY0S
DnK3KsF+oyHLu8w3xrQh8PtioI0ioGnJ/Y0HiysqxGxzvGDYFJ9dTu7H1j1J
CEqd3DJJZrhpcttK36Wkycqysf9MJatDa1FZ26dpUeu13brbQFkfKhxUFUMW
h3YI4BnmVjlHil0Ku1tMspziicgV4x+m5pooBwErqTuIfQ3z8u3u1sCRcCfR
nf+wmmWEFYYnKfC12DtWT2bQ23kbw+UyFsbu2r0nU+ETFcrXC0/qKaweldqq
oj+AidpvShSyIF0vkwkGg7zT87b1gVBnvJEsyX2IgO1MOHMcwizwdchpP3ff
UB/xAY3hSTWB/n3JCIhug8TBpnsDz0uOBw+XuV6wsUGKEYdPrIHfcwH2g2zG
eo9Mp9wyJUnxX1fCuLQnfTvRcSQFVlB4O5Pp82/LJ4WgT7kuJP5GhZdaHtXw
bTTKnP7Cz3ZMmXs5tg71xWv8NmHE4LH7xPpWZ5DcHyYhMdpW9ydwja4OaDrE
MTTPddB2V90MVgJ/l7ql+GPD72JUOYGotyR4Mzbgx21267iZPtLEcRq0gu0J
qxUq8KS8GQbyKrITMnBb65uFAlbm1sH0c5Blnw0F9qxpM4dMksk7ngaC9cab
9m+0r2F0Gt1IcwqSM0GNLFUTC0fjbYd9KlTlY/k5gkWIBfLoICuHZGSUtkfe
uyeyQSuMaXnps3SvcYbTDBDvIzge5dnb01gsV35oDlbieO/xMnxipcC9OG+u
3nlI5WFFFPX7DZItnMPzLHDb8MJArZ2bh/4/ZlKm7i1TzCIO7r/9c9ZXkN7b
xysqqirsW+uuDrGfBnVbug291Mzi9eU5cXud+qhHUyK/e9dwgq39FWK5chQP
h3+fesyc22I0jocekxfgIYl8qNooM1emL3yv8JeAoVofmF8acSdBT3DwhIs5
rat6u6eK0RV/urAypH4p7G2GamCfsbvuAaZrG725Lb+SpB9dO1xjGrZiJUxf
c6q/FnKBOzzThthyBgE97lmrXZpUt4PgefvcAsEAbebiJ92MQd9qmanILHWX
Y8FW+BzPw/Rxj8BbOviSA7lFjRy64+WHPQJVJwQMMPvTQH9QNsjKO6rT8Yrq
PHBfBqJ3ehb54xAjnO0jiCyG8NZz7z6kMJ6ymFkcSoSYWc8D6FM5W1CAKXIB
caWzwLRUIyiks6zsbY6uVG4xwmpTewrBA0XvsRmBhDVl571CPxytyt+Qhzqv
cP1siFz9FrQWuCZ/Ly95QErxEwM3qT9XuLpkXbrUEZQlPLctv1IzcOqVf9se
Fp7tIUnfJHk0wBfVVBGWBcLNAP7sOkI4LVeRfx3FwDFb7AybGVE92JMoezkl
58MHHIs0Iy3drmqwhQmT5T/PtdcrAI88QIyyWXc+kmKBfUpVHs7cnK+qqe+q
8H0GE0x5BcrHjH2F0sBnLaHC/6KnXw5xxwbvgMvuTnYNgBNiPfmdQ7Q4nLhk
56uCD7eAhDQ+kwazYY8Zjjtu1y+ksEXdfJ4DepyUEQFVsn47uCUMMnLTyeKP
Vdj9aap3HxXHb28/OKTWDMftaTQ1nIjvCPB42K2kKYn1wkmcNFXSRbKS7Y5u
pr2FT3g8zARNgxvTx8Gm82OnJWhQQ6PqxIVHv7Dr7V9NanK6PPfhaL1t9mJy
dIeR609TmSFf5RuS3nUMg/Uz/YCtkNuwFzami2swWZ427G34ZziHnvKbGufo
fjxZzeBpQm4zVrPOogEkdsggzDJ71f33iwF7nXdzpANWeZ2LSXxX+C2mkf8H
NEq6v/L7La8JgdZduCP32VE4ANmCZb9IAhsfH+NwM/R9/3VWayW0PsgXsm3J
s4KrmNIlY43L3UXsmFJuQAetDG+lzXxKbvwbRtn8/RypZz5DbKDtEtKmMTMw
6cwOzaC0N2xUzxs0pVFzQsLpG78UmdYsajTQzHnmhaDVYaBLVKro5rS4jeA5
edodoMBWUreAHfEDc7v9ZiCw5yvUyPcU3foNAw+8QPDu3EMksZ5GpPwOMGSw
lUpaU/Zktvmsh79SF1+vykaSvKO+m3nC1cSM+cuM+i0trBPo0YsjNUWiu0z/
n8SsP77I/iGt6i2dDyxoLxl7CFwpBp7wcNrzCXS1g2SjxnoLBITTBfvZ1frB
gocvHEg08/2m3EO/jG4OFaKU+krjs6EVuYOj5vT0+wy482/82Co+o2Pb7Q6+
CE/unhY8DCkwnrajJj2hKnVL566+BfZXlApqV3Hp1mjqQHsob39vpNnzb0iu
WuAz2njSTqMPALRrSgJttt/zVukBXgGmAlTxYD9PoafU6l8rY1hWyE5A9RYw
7PVeoMOrrzf8MzmIeDu/NzCkn9HWJBPG11JEET7H9Qp4A+VTonFJ2hJkxjQN
RnhwZEzgmUXoUEdO0KuvrTzqVFkzt+WKJyFehRcqyZp0UY93FTQflwhG6PMX
eQ1bRDMTKrUmih+lclwuUvFLKntqhs+omQXm5u45kqjQYVLYAdFY8XrcRIbU
F2wmdMri3Kvm9u1WHDsiX0WNRNs8IAlbVuHsmp/9sk3Z5X8WpyoBJkq5XyaA
nfsi71s7biweWI1a7IgagYLnIgFGnLLIvBlq15E7M1U5WNH+LB503dyVdraj
DeOj+Qwtj2zXdvf8An0oppnGA7rbiFIM7qpIQZynoTB2tAisbiFYVx1gW5VC
hmQbZyjiQFsR4FiUo0adhCx5anguk/2X2z4nPUi7AyeLOqvBxL3+vo7eX5Hr
GLBbNxn3Zoii6eY5dogQ3OsxR9NJyLG6TmbgNWepleEhnVXOcAbtqFeqD7aY
VBC6Ztje5mXpjztSguB2RR93AwdmBvwdovp5D2xI1GEsjXCdyh9wUTp9o2VW
kb1BxHUHYU+6ORUSWZ7jGQHSq1VKdJTh9QaIOKlX1PLz7xpWhbFolUMNyI8u
RViNdj76B6zzuHbY6gfwbaHRGt6zF6yIMeFvqzKIZa1V32N2LTcgCXF0Apfx
8N5BvFhUrD4D94GogIiI7JfB54waEbcRPEcdbveLJF3thLDMc0hcVZbvkJIU
aRTDdpQee/JGY6eOPqPGKJJmGzdV0rIgwJlppqzWu2e8SE9zNGO9iNz2d9+o
gYG6ot5ICdx2KBc3beqaGq/3lC2UXaHy4hFUcQ6ArjVjbAD7yYGUxNXERT86
rHUP7cbNs//NSxHjhYEeWHw4Goj9RMmyQWb6IIHitpaWTUKyu4UIkun26L4d
rg2aJIwV69Z1gHciPPvfRZJnicc9vptFC0ycnHJfGdGud6UZeskuOB9B2bnB
eVPqB0mGlAGdJ+yLgXHXfD+qhPFRWb0ThpmMGpGVZSuGb3mngObuilSm4kkL
XyQgwtS9gdL+A4/QznbvLpMBlDO7WaVrhQxVQr6klqF67vYx3sE6NjalNZ4V
cbwip45LDMOe2kIlRqSF8gI8MvQjM4ToDnCdfIF+u77dS/LBrg9ik6KyVjFa
2seLXimKIQDqlGnIPNKWYY+JKzovlyoHnv4oeKrAv3FNH0LV6pqAe8DEAlmr
R653jwCkblqFOjZo7K7zMuqaKk+lImfDeecqM+HN6KlYAW8HmP+6ZqjOmJcq
kf33HoSeOdsTnJg8NlsHbaYj0Rr4C5hfaWOWuvGQEkbG+u8BKXugBrlLqRAl
dvVVIHALmYAVwaMI5AHYgHKWgFn/uvqOQHjs//g0XdjaOWDU7e6f+glAr1cs
TLFhlo81UkH8QhMv6785z/BuwEneoz1ilT51ZvEKlkG+W+Pmr6Wvbu0i+EbK
tY6QL1gpK6Oz922jfLqCpt685DiEyPG5INvV2iKNjlVN7mJIxgrvlQoNovSY
QanjQl4Kbf78++j77SBXSyv3PkJvTwmPAirrpyw5AccUe0vK8HfbPZTisAfk
5gJgaCjU9XlyW/u8BVRFj6I1BYJpsTNRFdyZn57GoATBSoUgocfC87EyVjen
EaEfDH9WvRKrCnMB+cQlEXU1Qm5SzYzXhqoBH2iMSPuBSgjhy65EI7+Xupu6
n/1VSLHfkL2dUfJOweHkwbjF2mgaRs7JIN2wqAgACpk0k40odSY36TiMSnOu
q2lvXS7Nls7QaDFh9vqHAf+ceBjvjfcc1/GxcSn4dZU8FExhfUc2P4YHuE9W
B+oVxY5hY6qBm9/P2XjUHs4X5ZTNY6V+bgZ25J9QpEgb9+cMc1fojalaLSp+
bAHhYkrIBUbAngZgPgXmAQo1vXuyQnN86XXECOUvmRrUcdxww+B+/8OOsrGL
44MtNUPw+P/w55t/kSc5j77LELlJ42GiHmfkvZaRYOur8mcGZdsxv0Le/knK
amAz/EcpFqMww0usbBdIInvmaTt9dkb0UeVqSerBRFOxGLPigMj0pA4D4ZF/
6EW+zt1L92c0sSc3tSg6ELNqy5Rfq313qT249tPV3JfBBXpuBI86TA610mVA
bBie8UjRG7zMUg/TtnNbtM3vrwdbhE6nn8ckyPnkOkk2B5PnezWQ6Wba2X90
cGvXkrV4bUdyjDC1uOJWGGpCHdDl5ipN8phPdQa5BQP6DYhP0hJlUjSNYRBQ
xSTlsuA4Z9JLFQPtp8M+ggqCjKmcGiGpTSUArbRKIg8DJ+NhffH5yTXrEUG9
tDIAC8dyI7HCKJ8krTl598nQG2aWZmKidBmDmNNYv3UQkunPVdd97+eiu8p/
+RRllL8xcXl0fc3/NnYf26OsZsByvmjH/jjU6GbDlbGidw/8Efw680bD2oJT
YSLS1IIOKmOKhOxfKGzdaiWKVi5wxVqcNW+CdrROx+kFBKSPCRuYNANxNF1C
prkLFgj/6N7Qaw9NzY3bydodouaxI669zolRccabp+7it3bD5JdWZOX/E1nD
xh1PK2tEsBQFbdoy9cP+wf3ynBTjLFcuQylNojJ3FZuzRzd/i1TM0thZgVJk
PF/BPqZzXh2PL/lgAQkXbiAXjzx+uk+cvZkBNBxFpNe2OPdTYQ3LZWE8Beug
DuH+ARO4Ut5wdIjDqSKovrccUYj545B/gnRtf8DNV5Tj4VQ+r7rVeVE0dL1Z
3ywkgiY5fntDG0pr8jmm0GnWhevZpODoLPYfEiFpF31LiffChmsNU8m44W8H
44m6MYX1REFvEVu2/k5XbRCT/AgSpljERRNa61LYOHNQTbMMzlM6VwCiHMU/
Bm+BA8M39JbJq0AWzpcNauQF+JIB1vDRsJGBkVvrXmrWoD2UTum1QluyoNGu
SAMd02MYsGYnVYU+/zZdLtjB29eoJiTOMSoP1b96YHpziL2obPvHnhd+oHqY
7pA+yb5nSpY5uA4zkxcr0t+zCTaEzddMO1aRKBajt58TRG3r11jN0TBf4Ex4
JvIoJ5PPvzCCw5el1mGZPfN4R5Nt4kYlDzK+sn5h12+KCcQAXqtf8xSpBrF/
OQciSDyS1ENnD9YyIzvPPQrAEKlS2knoifFGOMjLKsG4dljS3YBPAlbc2FQw
CM5KgMOve7VSpdWTn+6VRQ7rrF2F0G+pdllMiCUgQ6C0qEc3KgIO/gov2qz5
TOjS4CXHCLCV3x/qz/dvt1gS2DnJxLxioAe3AHv+DHZQFB8klkUuv1eiwNpp
IpAc5jGLYGsDMUMEMWJW9jmi8aXtQ9WtjCJx1HRChupl7XrWnZJN7z5vZ26G
VovmVrElbw5MAhJkdPVPqvLQ9gY1nbjpKovsGcaqfxq555ivP0iDo4mUJ2Q5
eDOsdwzxZ6VaTccLPXqm/S2oE8zwlnBWmtXFLkPO4aCa1GyQJv65ERe6eSVA
5vSIc1Dp17Po8p6vfPUdJCIENfFPnlnFraveJX1wIuox+poK9XvJ/a4I/fei
ZX5dBPAKhO4r09MC2QbErEKpFmiFLy/6wNHHYpfVXEuGqiZhPWwB0C3UBTDE
jN3Z25TQJMV61q3N2+biBY41N9U6qRVNkyHKbs6mVigTp20W8r/7Y5IjfYI/
b3+lL0fMeL0lwwC8Fj6M5Fbv8hyRaUl+u79yN3t4WpPzBFGQdlmPpS5RzCHR
9PeNggftFE7tceYt+Dwx+v49B5BfGdiqE/yfkqDoIxGPBnQpR2b/rxpCrrG8
IZTJgaHw1Nnz4WiuuOzf01teJSH1jY12WdvTgQnOeO9h92TVfqzgN8Rhhc7W
Id47+3h2NXqivdGeKe8VT67ZzJ7auRHTIPr1e/SXD04e1bqXCy37WybpmR9C
qDOAejn2xkUvVHG0eKEsJnFEIycVemjCq+Dr0Nh7Z9miz1MinVqo5d+WQVag
qO0ixOv9a9QQOXvpDFEhHgB+zD5cBtrccU3b3h7GsunF/Q2yELMqPamOb/zf
YkNacEXaAYM3MoYqe/O0mK29RfADi8VunF+AYl69TyABBfWclDpGKKF0IjmN
hjsfn2rhkLG5a3RWLBzlteRn1b2fuIGYblrouvXGbEzMPkyXqoPWQ1WSvVyD
WMz7iaGq5lJEtCqCTLtj53YiEt/XvQYV8XXXgQySsahJ/rTKNKwhb1RMEC1J
zS1rOPLK/LaRfILCvHJRwJlWbn5Gs/YWgUQDc6nioY16SpwzD5BlqC8PUVlQ
h0slTIq0J0HP9QY6H8KJJCXDml3Y5OpVDKhzUfWc++LME3fHwZwsfzSi5l4F
4sHGpswkSQ0bk5/8UgzVbvqanwrgV2+cDv6ue4IssKHYTO/t2LcimXVqN9qO
b1ByWjcPKDxqVxTlbnLg1Ge97/TZkSH0Mk9nDgsSioXZxCLiLX7l8SjE4IT7
z2VdCXxpp/u2rtqX1NZwE70yAE7WOAeXSkUdPUVWJ4BYS2g93chwV7anerlg
KzZeXTgofnWYTk2fO8LaZ+SFNAnXpyHtnTkPvgEPx/yUOrgnoofsdZPGMArT
rE0AcRIWz2enjkaezYZ+0odoQCBDJlO7mjVcKtH9DoS0pkKj/O4JJkE5werZ
3UuEmkc67GfSGshaGxMI00agiK2FIqGmregoJCZByMzbZerL/5iWAPaAVgX+
SRwXw67z/X7rYWUsjsRTakeFhYAnFKfrmpXxUXqudxGFlzo/Q56BweGGNxKQ
WP0dakYT+lJNCPrzjT8psUcFsS1DFvf6jOzIN/jA+qpr80La15rqXtdXe87U
5ahKE8SKBtWbb20eV2P8lYXtjMfSsJVlTCpgvAgGhamyaXUvROOfZ6u0ye6X
qHhsu3UrE7UEC5cWa98qL2KmoDClRGX3qwgG2CjLHnfae08W5bVSIMihiaB3
WhZoMRVp/ty67HwCNaJohxmG/ATM9d6kzMSw7UTh4V/10f93tJTfbWCXLcS6
Rn3wlhDJ8sb1nByI75o8S1J+4BKrYDR5NncvZgPVHuxdFRXfytJdHZQjHoW3
xClMD1bJSZ5ESod4zVFL4vNDUTAuVWP1opkg3LfBKqPeYjuMuKprHNQhGgnG
uMJEy7L/2fhjghpJssJV4OBlK+L8L/7BLFFqTV7XExA0HwX9RexCGh50m2NI
eCXeMF4UiWl2ZW5KoQRReJNqFrE/4lIlI9DGjHX6vT08sdu6lhGMBtHtY6L/
P4+NpTOso9ZGYYw29kXCYJf2z8bnH0lPC/phfrI9+VU+zcPo1gHumqm7sVt7
P/CgDlveneapnbkx7omN6ujvjOrje8Xyqrs0iA76Z1jiWaumRpfRJm8KWjN4
pJ8aTJY9pRLv0t+oWnAzRkzxhJvnAZB1/R/M7vJ8Csps2YfS29cqo5Wtu88K
JaDrGMdGe35bCbWrqAWstZCgO0l4R8WbneItPet4CyV5ehbldWeuDzHLjU6t
zn8XKXmdown/QRs6r2n1mjuznA1QsOzYFoO1V5D+hbNQkjPvXuJS41qsSYMz
ABXbKjIs5EqbMwSGa2pfILu9b3iUg5a50glGv/6mHUE3dl+9FECd7Ql/Bj5c
cjIB24kVJGgU+QAeQXW+tQEf4EkZq7JIwNFLcX+1+4hgn2GJqjnksDl0YWWy
pUZzBKejLlYRllwSTyf9qdJcLjzsc2jali1UGwZWme7AzQHRlyFSswwnuiif
8Zatp5eOcHV6Jc4XbRqI3lEYZ0Tq08PJ3OgkqjXEJV1G8EyGsyRE0X+OwKA9
cZKMoMBd630WSYK3gn1XLMM7/IssLI6r14NO3+wD+osuTKegty9XNyDaEzVc
Mua0IoufKb27XrHo93//84Q+M51ykWCEi+DnR/rLxqfaxuGa8rrLvzUP9tf3
6g9vY3fwRuZBJcz7WfCLiI7uWt7OH5OlsoGo28LRJVT9ZMS3wz6/Mxm4YfHa
/lDLb/4E6csCuzjAqc5c2rsog80ukJUW3bK231ZrFTj4gQ9dQMhSYzsPl5pD
d/47wtlwIoi4pYBtG1Cfxa75VNb58eSVgnfLB3LS5YLTi63E/hHCXW53fnv0
bmG+9ewoeS/0QU7i0ecRt1PO0f8WQL+vTxxEAYG8vr7pNZynaY50QvLc5lPh
0oqe0sz73LHfFq7GfwMg+CkLe86IekG9znEDxasyTfwzhRJ2bIQy6TA157xi
S6ASruzs7jLJ/kOVZSKUP4GU1SIuDqYrtFMEFInT4kKopSROXf3uKyf21sSY
QYPhL/XgOgfd74/JcWIemsyl5sjk8jbiHnN6rZ87ks+O7b06kCoeIwm7xw1y
UToMLa1EgDWaIlE5TxUapSeZ3brEcqFRxWUnk4V9Pa96kFLCv21oAnsVqCs8
ikPxMamo/nNHQ1BqM8eBsZYGIef8I4aLAUy5Z3roX3bXidGBxGQYggs3ki8w
e+EjKVXlCc3l+o+0zyDCwCzkPzFp94WjKeeNgvfI+QgVdWHuHmpwNsxIE+mO
/YNsAMh4WSTQel8a5crFVePWvhTnMYct68IxiWdpoXc27zeyKjrJZKrmDkHw
hmxkUYXVM/jl3if4sfpkxjGuSBj/WtBIbbZ0nEG66ZNqOfCcgpmRdt8MBL41
DcDOUK+Da68O/uLq3oT4EzZqksMl+OyfJ4zFkregrLJYhwjthfGjuRDop4UA
euc9QutjY7Yo0TEYEJoad31KwYNZoobNxtNk1MqUeIa2JvnIcne6d1/RnJnK
ohjY8j5J4ta7fonWBqHB6y0miTDiLhwXEsWO+whqvmMQUi8CMa07smVv4nGW
yf1P++Tfphu/VWX8dBBBqH5hjoAboPQfKJzI2nU4oe9l6OHzx57309B4DLSx
l+a5iGdr8Fijbl6hqAKWcPyvKtHDgly0atLo6zGSKQPsn2trN0fSH7HOU4S2
2M1noKxMKomtIJMF6pfGeYDrZJYRC7nlX7SyXqgfX5++GYAZ5PsLWp7C1PgO
KywVGkuKYSijfpmsxVGD9G/MwOGyQylCGQjjzKRTkljlGOM4ImiiM5S9Ue2l
7LkrAtF7CqMHjJ5W58dwKQqDpwiElgmmKyYSm2TG4sX2i1fpl5LQ15oBcEDx
mfYnoUitedtmeok2RKc6nRibQNOd4INdqQuQcgvKlX+85BKqLY/M8yAhQDQX
GnYTr7B5z1VhyTFej8nNJZAhdRI4jBsccvTunlAD6zMXDAByFf2HEaA3a2Zv
Nt2989U1UhesAm3M5f1S3e8S4eTwFtBsRySU4/6pA1ZecMtnJkkdf3fBobPv
Vq1RQPApg9APORC9HymfFdrqlUyS6QcIJoJxJW3ve/RYHGa3jMpIZozwUjBK
pKHNduwVNHrIIQLgNVgJL5Aaewi4ZqvmCEZLs7rr3ecPt2XNKV4sZABBoiLO
t91nsoPoBHBfKDeLLbZsrllEPZXG92v2kiWrr6wKsUKSToLLXK53aaaYJ+UP
zlliOKBZRAINHMo88dGnIqPMbnpA4cx9SuKmg/XRSmVfbu102VZKza+agPzM
E/Nm+/jhzO8yeZ3scKUyFksswjKOUojydbbi54oLsM88Ymx6QJdxoxiEAekg
doOcGdP4jDJMvFSCZrqQyorcLhHVxXL6Nxqsow5/FRUGjSrU6grimA0TrT9m
xOJB6wMapiAVXziM2ggiMRQhz4NKnubeVADc5Tni7A90YKVCzTRxCPVgJqn/
KZ5Bl3ExmvTg2lUuvWYd/VwC140o6KOrWKjTOpEzSH4fcRBgXvDMYIEE7nhi
m2ciVs/+PASG76F9jNNEZdvCBBSr89co9S8kFI6YjYWSpy0HgJU8z4LR8gwH
7Qs5GMtk/hotJCuVbzrl5Gv3E/VPBcItVLkxYfY2XXk4d6Jeuh6pTD6GdCst
vLgCZX9S27DZmMu1Rid2DvaEYmKWEJIzb/meNhPk0fAJuKOBQkdHokpNPVvw
aeuyh+ZvPc23Jxnvbfs1qNTCKKB5HUkPEGWjGqWj6epI8X7Pma+WLWZccaxi
YHDWzrIfvJlX13mTGCeud+nCM9H/vTIiA1t58qmSJtNMfSt2ZmXaDAXSRimV
V30llGNxUE4g0AW/NqGnNR+7FTpPIZP2l/UPitQXnwUQNwMcF63YdAmtOSIZ
ARlXq/98ir7sCm5tgEPg3nEml/yrc9HNuxgLjiBo5Czxtfw2vKV2RxfR0rax
6oNPk4xEfnPIeLdYBjPAQ7Lh3QUSMprwQ0c/2FIzs5zFDanUq/Y/otOxZBlQ
GzpeehkQJxbcy0m8zTKfl6wIQNgpF7bl4wj7XBUQiH69EO19UIHVXj6n/i58
NoNmRJtpy36hqnanaxAEm5u8V8GYqYhfdkWoPQIprqTrOjeu3izhma7r40Ts
Xj2YxOZS1b7uAmZHMoy3bS6F1C8m0dd5Yu4u/Z/OFyYFlFK3sks91IaHZsY/
+yIm2IZ4BXV5UGLWTVzokm32zPV//MJO8p/wyzrKbON0KYYOEYIpg4Nne/K3
hMBTd8sA9AHCny5gpS/xu3Oog6ZafPMT3Gpyvkj2GDCgFHFmG9erBkTQHP7o
AD+0dpxV+cnNHZpeOCbIHxt814vCaVq3GpUObYxfj1cLO30spRea/iOqbkGA
qBoyzMu5B1kl8gikqm6MG9ZarU2fFoXZtOpfC25l91yGi3Pm2vu5wKp1Rfiy
/7dlhiBULV6WZy2FsKGKLIpdSRKk9WDF+KSiLK9LiFDt695IWO482PKWRVPV
M9esOGBMInxNxydNRoTiIMKzeidUCm3Mfh2BaEwiIoKcyvlKEUdxfHLW/AnU
UtWc5fippemivtgPOZRRr9efqpVA/ctiRbHKOEogBMa0FM7uTnPIRjfUsQ5s
JaHC06oeUTQwfQQseq8CHsWuOP8yoB0mAsT4A/JMp4R0HMJgj8ALS8zwx89S
vJnFLR2NBKWbFftFo5ytTYlXdlj+7nV6CeovEh/JUgSJDN7DgggcyK3fVu/S
Y5kxJ6nOG24LXvh3sx9hyHEkS4WkuC2ow95yL6IDfhGukG5CF0AdMXjxziyB
axHYds6GbvXBhd7lokW+Chjccars+Udv/2TLpumliIgIngiv4S9YgDZ1BGZJ
g3xMeN7hOC0pT5ae1ZpHT201LHq8Eq6vCm6zVmQdhmOWI7r82Vcu08EQLejo
jrTX0k4eKnCxDhVkfJ9JXc4sHJqdCqZ6UKYN4BoGYPahy5d3PL3bgWLnkKRq
neZXGAj15I1Czaa5rLpcPhUPdGEPLYjJKSnuXXi4QNdD6cGEtMZ0A+HYgpF8
FNcFOtvZqlhsWkAE9556OrYB2iJO204H2guaM3X+J4wPToQwq3lYUmo93qRe
Ti7HKmsaPmfwSx1IaILGXX7phGeWsVSiq9hkODmjSZuB71KVdQV+NxLGwn5A
da9saZVxe3TCEtA+qlBswS4BwvXpHDNzASWRrPxo48DnCzqO54oN2ZZKEcsP
7tinjTFt+9fRoS+dP39x4VlLavO0KdnkBDzRqpwr+e7AqoURA9adjINuqzof
xfDuZHLYfX8dhYF7zfC/MCN+aclyQ6DcDuNugmLqc0a8htmOmkr11q39ZsfM
KpfBdT/XPq/0Fw0y59+Ww904lKJ44ChaKeV2XcBeXnkEEKrEIHMMp9uqBmW8
UtvItBBsdKipdFw50YHrsnoaQP5ne837n1/xPZcIcb4JZKlHMmsvncvfbCaY
Ss2xbMASKVeZvL0cxmTtBnNUvMBL3TojSo+uwwY80i6tqcNLUA2426BWMAev
Rf9UpMLvt1G79vwz/VKi9G1Kv7vNsCnQLNVKW348yS1e+VYE/j8ZmQZbqWCB
wf0YMu+Dri8jox8MA5+8FsZUGsnu8XBqJ3g3l2JkGPkS0GMQj4xg7uhj4Si9
uloNL+7VwUe4mW76vSrlNDEaJdWFZdzdwi+VvkudgvMCPBwSKoYq1lqw63xA
kJn5QKCOLLW3SPJ5IuL3C5xSU25kKfww8p3wQM1B+khMjBggvr8WEhHrF0qh
gwnPLMv+DH8cmyMSARPQrK/C+vf9aj12dJ94/ECR0BZnyL2IJndafVffGmMr
qPbw6b9X8kVHIxBURnYDHwxJU6A1QviY7Yy9dqheOvZxnnb7gZ5gQQF1/Sow
o/v8shWhPNcuRcLMDXuJ8KvzHTmFyIZFucUUL8b8SLwIm/dWE1tytHJe3inP
cQ5m2+IkQuD8L/IU+xTF/JKpy/+00zYpdysdKPjBs37N90RQz+iVeza9kIbv
S3VvO+DMu1kUSF5oF9MXIOZYMxYTv3rtO2qwTPdAh07OrVUf3tJc/uDd5WZ1
W/f9cRvI5F6/9kM7mZTFTvGl+6v5pndHH1tx/0GJSPJZorgTii7suMnLqSHU
Hk5INu2ZoDoEmKp0etEY9UXDLLsQDv6sE0W9i3guLblE26hWvNdWaThs77BL
hlpuonbmxNmy8el7Z2k9n3K4+yRvzevubfPRoKT9fkwnGfQ5aZW6gHUFTlBL
v3wNHF4/WRTlN4t0Lm6JZZVgCxrzYCsyEgvuFhOgABXHZozdFNERoKx6Hh2j
IvIkk508Pj6+FGH5U57TxLjJ8bYtVZ/dnaMfqfiv3KegXHTWMDa6DmpFdvXX
6sSujjwVvIllhmNLuqIO0WetkwuDBWksVAcbaCz59atzHWkfij2LSjeop/ZA
ZG7oyOsCZe+jyMXn/GTC47EK1ZUyItJRCIMDdU4bMTCbwMN6+qJSQYAHfWkx
zw2haFaERxZlFTxoRzf5ygiCTNOg+hrE7Zypo9EQ/nUOo2YQSz0uE0jsORUP
3q1dXbRTMLacWkXLUlBQMyLUySMU284d4ASlVMpTScrbO3w1+CP96iPKCFme
Vthl6PzrdP8T6f7C/U2xAiGaZb5XtMmvoMpt9zOyx/qfJsNkHjYKpGBXRdh4
Dmn6IFZ/8eUboq0D2y9FRZ4TgD2kT/FvrSOXVu2D8BuYQmiRJ3JYIexJqmmE
mC+H4DC2aVcx9ltQ/eFLv2aeHg4yMLHnJSWuQyH3gAujRuRuKQPmvBjFK9Ho
BN+udK2ux2sgsNUiOFjPYaLawTZjEcMflkKFjljeqYkqIa7l4gChCvTIk2Ax
ouxBaSHjuOlGWSr/CUi4vA475y2GIRLpE0+k8xysRhRpyMebYktLGK2Y2RCs
wnjRXYE5umi5P+N800280JiTtiXInw56fjinidZ85MFSpYTvFH6pn6Wg2+Co
xVbMwxjczBC1zwplsOuZ+VxEajnnE1J94r8ZRmmhc0VZSbcs/Qhv9C3c9Z7c
28R/i/44pFsTEspt81UGMwfL50pMbQHQ3+TThf1FO6l/XIKLw7UH0i/fKI0g
dO6yI1fELregQlrAMOo+JoCdoIqMhjcD1e6Rq8qF/IS8mMAXvN0+YM0wiXAI
Td2zMV6xSrMmBqjaDQt2ZcGszU/bIMCzGOwhqjKQkfT6AfLbdqLFDuAZhuwk
1sW81l/sgzM8zfFSAC2yg5hcxg4fmLC4SVXYKSDjcdMJ63vll6WGV/4vM1cm
D3F5wsQhgkMBIuyFTycnnGS7J6fzXXw3LrsRtwUo/Bhkp1zKg4BfzSxAi7jX
m/re78hslQpe73QSdnNjSeUTIpvn2kh4HE29s0/fHnOrXdDWRcAQLRqlXcap
bHQeL+JbPAXQWEX6xLu9LWf+4eaUo0E44yCg+H8xGdQNMfkip9nadnrIfu/F
US00FAZsVEcIV8gVJc2UuP04F6cML/3D848/g9BqYEXMakYlryXmQedJXGmS
zjgkSD0vtuTwu3zmXRdyIov2RcKhsY0MqxAjPPt4pYon9doMWtFJk0ZSAaO9
OG3rnkQ1EaqKslxmhfcaLAFpWlYOJ4tgCX2/AJkX2cEhe8+bAzdcC42SkRJD
loy+bd+KgadqCfb76u55mPkEJVY08CW7/96Q1B+npS35lKIoA1uB44OJ2aFs
sWyl6e1Czyxo4Lj83om5aiAsYrlnN0tBTJqTUL4VDSu+DBKskdfhn+02aWy1
5kNJpR/sf/+KQwlLHJlYlS+G6GSapHptRz8mdfvKVFKeNKKp5gIcTXz1Zylg
ozqiAAjPeSUKfJG6FDWo4deRGnHskHjA6naDqgGhgSz6U8l41eTpgAFUIvFK
FPPMl6Z+PuN3z2JsgASmYbKsNidU4KI5I6MEzYwVXaqJIdGwpxRYBLetTgut
z4hM7/pMgy1JbpBDzJwVAw+xM0RYtfAb70pb4UbZdvJWxc7qJD6nJx69YBcq
OHAJd0t/2/bcccGTRLkdhlyE5pjRSkWKNXa+MqTPscRDV/CCwJoGtNzy/2EM
2lv3PRvoh3t83vDR/voUYug+XBi1fYCjxwx0+vLJrqUAHq+FjaBYVt0KIkt8
EhJ9TRB15tYnNRnjAi4p+OhXPY9lgQyU1PZvGOTCUmNT2NQfO2vpHBVMOgxw
yMMiSYL+7PFzh8+XN+p+tflZSmMyPGDbFoFcABR8t4Q7VypcvTyuq8GV60BK
QFglX/iALdHUWAexCciUCTWWNYuAXmexKvVDd/nS274JvxnSOv3OcjaXWd3y
W718ek7GNfsc604uP5oT/4iNiD8JZsHfqeB2UCQ7Cbq8yzFBjzCizYRjLuq4
DM1emJ2efwQb2H6y+/fjutpOZIM18IELQQGxLukCgKzqg4SIgDQI0RQJGmM/
PDMfvSlGk+vpsylpBnZQLFw/fhOi5xHoVSgOmXeB6eHArwTqWvRNnOXuy8bp
Kaxjwm89EfVTdum4IO/Xzy5eLyYtSfL9OI+uki5bw2nQaRFVTpN/9BbMiH+7
/+fv4Hp18RW2HaftcU2gaZPR716CeYmVIdhbBCo5DHzBS2d/omGkRMjuhYTJ
odpJMEp6WBkK7OD3R3fFDkrFCWwfd4BUyya/Om5OoxDO2ODdTx3llTXwIBfE
zMhKwaKZubJ9e7DUl2NFGK801x6Qq/s7T03MwW/WH9IeDDOxlh4E1MfjGVlk
8b+Ys5AxXrqLgtR9LX0II3ua983XgwhEvPxrI9Vwskl7SGsh27W811jFB9CM
qsWbIGFC5GAe70X3HhyoVUSjDm7KP2pxqrZHFrzfMD7twYpesbmACuk8j0Wf
1XjzmJFif5egmCFhqyuVamDPkXDtYbxVCiG5qFwNidFXGf/EuxEMDLr4RnO5
KUGo04cwSNliX4LBYVOAwpyJsYc83sly7HqQFjN44AhOQXtP8DaYHk7eYvIX
mRoV7vmfxDKnrtf87zVjlkVWSXQPgQ4rBiPDX2SuFKzCHEEaU7x3t12WPy0D
hGRA4gkFyR+951Iw7SS6yfvqSBAylXrrrOdrNgzDDTnO5YhEOk0ScOsrHpT2
wsoiUi2hE1LnzXY6KADAZE3H56Aoo4ih51FIgHX1eDdImj/YAhNQw10ppBhz
0MH7OiqX8eNw2P/el3gKs42aSy3N8RR0pHtAiJTRzBkJOumXSdmwIN0so9tM
s5kQLyy2ghICLhi9ssMUGrdld3IH+cvcaUJvz+gV751YwXGdz7IuLI1LOsIZ
WZ7GlPgqAm90JOvuIUFsvq1QxWrAVlB4Dx8QGpumASK7SlMGhjt5qM3mlrfJ
n9xnQVQkkfPOsBkEBx8ob7p7jOaO9W9YtlR0uG5fIgtSm0gPzRK710rlL+UT
bgQW1ow7NuYfiFcNBwdy00PWXcV/PEE6foXaBp7hPcNKKfGH+PU+8Kujfnex
09MooUzpQhsy8bmUU8hZDa2GYLrMOkHUfIFEamwcTAzLgb5qgVAedM2BihLN
2k95uVx/CXoLkE6cGlkWyd++S/+lj/YhIWGfkaSa5B6dZSQzdA695npI8w1Z
zQa+8iKQGT9qlLJ+v2IIO+pUUOQgsmj4WwhTuoVsIQKxwWXPXrL37c7j1IdW
tDvCs62+xypoN7CzR1bf1lHEPsPR1suIo4xzu8RZ1dvrDi1aXycQ1lJG3aWx
NkOWYu+gRZgtnjxDrttXN8btmkNkFGHgb8A6C4KGLfMHxVhzJZbn8/YU+UwI
YgUjeVwRApgo2OCCdb9LIht1OBD7pf7hSO17nUfO5Q0UdJ+k1tfqxBnQ/i8O
ayfOnbBKXLrk1EByeKt12hmJLEX/Ke1/bkiR5ktX06VHxun5nX3Btk32A14q
d4RuqEqZJCiEAsi+QF6d+OQFVp/hWwRhL8Od8ADFWnYgUOlHG9XaBb0lesPX
dt12wCXPy1CUDa2KBG21vQWYwgV1gGOK1i7EeyyuqY7bN4pMKNxxjgtLR5EQ
NKS6ral10mo1fHwpev+1xvl9TBuxrSqlgT/azFgofjFmPWHHXEnfu8KofmPI
4VEVeaHaNtzvRoRfopwRytiQhk4PC6njiHQoWSGByfdtjTx4d7JrFskBhiVh
6s7kkrROUPiFDFKzFUNbIy7mxYLYzFJyyRzPxjpwChjEPAUJgVu1KU69baGK
1DIaG4e8rUMerlvLcGUrY4AketmMjp/IlcP98qv1NPB2MlzwlULWrBAfCiBr
et4z/XHDgcbMhwzIniQeOUMJJZobh8mWoTR9IGA5rg4QVyCFF10hp7jpoLAH
ZSpsIyjKS9Y9Vk6pkXy7tjmOG5ZTXCWMdSByr4P+/VRTjgeoEh/tcnbI8lnI
p32chgZq+6EpISJJsit8yfGYevplmDh128kH5Cukcdykj6fAh7ZS1h1qH0qM
2bFV/Ql0obHCrF+ENBdVY0ZZSbjX+hj1En8jug5u9q4IwQpfXylc+eVNumka
IqSDbTJ/GqrKqfABFOgiGGPbtSTrcoZgw6XVcFnIMtmyPUs/DbIY7RQWKS6W
BwGiHxtSHxH+GnT732q0bHiKMrrT9oqXDm+xcw63KvjEbKJN4aUhYtoUUdgq
Wv/p3Gjl9vJ9b0cNoLYyWBAg81mXZEZA5wcjAzXFP8ixW+3UZJJqJXkHtbWd
sj5cfTzF5fmjbEsaDu20ttE0A5mu1C923ul47MGIGrcA6QesYwQA8Q0lD5SY
SiQ5LpjbYsvzNV8p60qUFnkyU5kscOJmHtXCysLUqE87A2tAJcVmySvtUPs9
RHO4x1SWpye8fL4aGqKDUTdLqXn4h1sMgEBdh44aI1mBqQtObFm4lZURSo6x
P8pQTHIaJZL7gXXNC1zWJWuXNhbmOwPLsR255FxTtPwdIg+kd1W5gZtJIlmQ
FUNTR3W9vaIq31jtLobfFtSiiz4ZIkzwoDNIvrdgGG3NB6yxjJKtKLC0NXqV
ljpZ2+8BWGW2MltUoDD8Oh2WFti4BFmPPbJFoctwJHNIcZf+aB+7EhKJf+6Q
ietmwS1ioZ3+RWZfSJtOQIUKHuenZP5jnzS1peGfqdEpD0Wq+52Tj2nRJQ2P
K0+ZHztGJR+OefExqrw8kk4yrUnE7lI7Ak0G2Uabswx70ZVZRJ8kK0wyD2OE
UzGCWmbCpt9KHoGKx0Vcg/blWSQGoZasZJln+fnUurL6+STV9rf3TMf6+rua
5IvBhxLOXEWA7nTfuFgCseuEjvq815BkMq9g4R7NJJKlTxOEGmAtP9Ah8RK/
5F5ntlhJ05Yg08IfedXFhEbPvM/hg8PDxOTlbZzPu99PPTNhc3coA7d/1HPl
lrthMGvpHz6PUYOXPNqvqixnWJcz1qtwi1l69hC712x9g1EEqjV6JwMJl/t5
8Lm5b6FUY0zFVR/InlE3iFiJgAufuWQFLaBv6QL08o6aDxkGwTG5t+EocKCY
FLS51rKye0Gdnk9n93U5lo/OR1As3Pctlq/cgpkfZmb5caxbVX+rsteLWnD9
6p8L8PouYJf8+4du0i8pAT2HgdE0v7R+ZvwaXcRKHZa5cxl8pxtLyzC/FICZ
2XByKUo29Ob76Dhw0S7mG9Uz84GEQrxIrt24JuDHUJ1qhlCe7XE70DDEMpEa
4E0qK7UmNK/ZrGohz2LoijVuposbfHvsSEq1t2QZHAf7ckkK/IOpS0jCuPXE
tOC/+W/1C8j1ujR1ETIiQ0WV0xH0saSEaWXHfqdcqE3/QSI+LjNGZD0nMsGg
PGQihq8wAid229YvenFkV3Rb6nMHEQSFLgsjk3JF6sRQGZgSRdQxiFFlT8QA
qnOnXCkpE00HuGXBssu6GhbgsFvro4KnrLJNaVvodRs9yfPgXPkesKdkI+kr
5or4mct/rBajCm858afpZ78tRdwA3KvmkAnqMY0v5EnNsbFRNxV+u648o0Bq
gO4+Vz2jYwqHJzdbx4O4cxWEbfz5z/cmcX8Au97dIUtGFB/ShnqxX2MfO1c1
GVed3RulD9TZxOqJLD7A8e2wxzILO/amMWwgIZBxjt4QH99O1zk9jT0nqXBv
sDKLB4Td+pfPiEF/A6kosem9xaTnxcAgABOCRUibQyq/a3wKuqs4x/cYA3IS
BSMTVOtg4O0lr13Siu+rojgYSrrDa2fuyyUvfXHpHPqsVreX70FoixzMMbHl
Qj+o/f3PyZ7UzzLYXBG7X7V09JkjE3aKsZJY6W5PNzbXwuU3knSJJsFSkdFZ
uhKV5aH9anwSnPJLjryrjMfU9ttDR8DXPP/PnSOnf43t7tGY9pcSkLRTD5jZ
L96PHj/hYHtYeDFydvjxdxn6FFFpEA2EXy778Nx8rd+2gU8KXzSWcqA6S2ZE
48pD4lLkxY22BRBLwMH0gueTrbzDiKTbPjtIbpjmFojcv0MnLzTvhMLZcSSy
JHo4tFYL3XlGBjoeL5z5to79xcDSNnhewABU8DE6XOpJ78PYhanxbGauN96W
ZIOopMSlSlalbht1fePc05Kju3C5tMC+mi7B72K6EJsXTKKtnmvVHb040zL+
bKZOTUfjiKk0JezsDDcHRwnf1DOeCJP0viKd1VnCGU2WecQ1K+aCqFVGMc6m
VOa2Zvqg9xFpOBt6acxQItKICoFyaHMBKUijPA1rZr392DFXnwVMV8W48j6j
Q/PS+zs7TgkGJjG/n1LjzHWpyr8PdRp4+bxcayetxlYB8X5Rv5Showhh5UVq
bucfkbvd8JkFFSCmSI9DcX9uOusnDLsRBF12Aehvx6wutbYoyWsl6Uan9OF6
NUgYGI4AxwjB0wiKO8BrldYHdggyaZw+9LjGGNFQRvXsy9KdKnxJousTxmU6
YAr6h7yQMZT6u6b9Lx9wQi/VkjChYBEO51hvG00kuDYG8wVNCP/DyKl4Fnef
KYFPoGRGhTbvuNMAojVOgb+iutLgWbn9dPKUfMmnGdt2ARPm19P/sGjyG2km
nBOeDtdHdjL00KTZMXxnFn3mexIN2hQAh6mzlnRvE62ZUHJrIsmRGSmKeMhc
Jwc07OKliEX55FLBxcf9pXYGT6vr8raDrT2AUe95HogWqT1s781qzGNRjm6Q
y+YaKf+dXoKsh8aB6irzcFplDgXowVPg2f23LJxELlXtg+WmtGGubLr88DY4
D/rjtZVrbK4OXf+aSl4t6sHsJnT+jIzjroFiWmE0Lm4jYQRZ5jGMy1GR0nnT
BtACF2f/CW8s06xhhadQ0Y7kZzL+ztv8ULXkHMlfDSQLBMInmu1u4Hf8htBf
IBWtivDSUGhCT1dRerGaT3VFOJ5metGbOJg7Uk0swS+VrM43h0NUD0u63Gqj
Hyt4tqiCeB6qItCC6WqgifmA5E5r5KzhI+GRnL0b9HS+N29BR+9tN3NZym7P
hRd7dIXSmYB3MfntuzrfDvbrH8w0p8NGWu8VWoP0Mw0OI8kWv4gaFaMazHRT
5R8hYAbucJDDF/aDQLqEnDA8C7QsBMtN4tTLW0l7q0ej9hjmBqXPkZcHMpZd
zGv5kUST3s5Tqr591Bgf+oH4YvhlRPHpzyMbeQJO9Gn4SVUpSsQYhHo0zrwk
TVGg8KEcSN54AWn/jX9z+jw71G+k6SDSCuiSQEoXvUXbTaLJowjWy02csLRN
WG5eUrGUXlpT1jV8ZEErvSJFDu34O8EpkgryMJ7aY+svHagZJ42eA4AoBhpy
LgQBeOBI3Cm6uIgHsOJv+XtDyZrFuiVdIUNRAP335bC28/DOHADAK1+MmXtc
misnf8FwyyRnzIGULckR2IrSKbQFYuz0RpAb1T/tlOv3FqfsJDp8QRkm2nUR
ZMZhMK5timX1DW+wNr6JEMqQ+5GaS5oJ5gq35oHrSBmUgSXOd7evGwByHcI6
KK4Y2OfK4E+oxfaqeTefpz/mxgY6RYuUegPT6OS4D5K95vG4u7u4cjJiX4h5
hrd3VjPOBHjIlGDGMAxyCx72Vgk7PKhYZmpLJDPniff0ga/R+3Q5YnmvA82z
ZtLvJ4BTRFs5nbkyZWvMOYqWZIZou6p19K3ne4xcmVc4lkjYFXrwcqLnJLT7
wlFeYVDCfj9N18n5bbNeg8E07cSz+qFkOVZvzcXAGrQqXfHDGIigQbMzSVj4
po92DPctajC1ok26jN7SM5FcORuY5Setc+X2IS+qqqCqXoJS5iqDmcI0/4QE
l35BM9TtiNZAjPNkrn6qVBpr/BC7qH2kKIiLFGytEOoNKYISDSEVxUosTHVj
gekPfPQqa2NIwNmOq83RfF/Q0c+IThsiTN/ZWTunIsAQUSwqR6TkLpxC+5Oj
Y/ZNYxL4irgyNdwZbqy+2eNSQgp4btPiVrvgGmOsSFq43Ua1SqdfqJ4nAPi+
a7wSpaPudDejklgDWb+hJCre7b1qF2uEtcN0PiLBlNxI1ww+BhQG5lW0uzbd
kIXPC9ytuBVpcQWygK02oRkNnLKnsSybmpI4GWOWIatLeDNQM64+/YlDvBzc
9pkbvfBNOIoyP17MxYOdiaa9T444qZ5RdW1g0CMOEPeBjdovsUZPsw/jo+dN
pg0ElRuKRgvW9rElA3JbD0FVN2SL27ZV8mWhKtxqxoqFSHFyWzmKt2IlOMQZ
nrULE1rd5psFqrx9VTJrTK86epTYdh7gAKigobpfE0PFEZ+Kyv8iTASAajcD
93V0/O34C3J1FQxid1Ef4BUXfogFlmUjOo6PftYuPhulsH8CzO4KZidSCo1/
7CmZcxIIeGZqXVWsFFsr24DZNpnzrz8/rwk7n78I132aLoDCWi7P8EkUoMju
kYrhtvjQ+E1my7gtNvqPMfjv8PNUewEuNCAMVdrpMVDDRt6B3a4SndnfN1ws
UE+6gYORFM3CAzqU9/7hdEVlhfUzVn63+HHRYkO7144iXTfTW9DNMEFZ/njT
S7fMEX5eUZoHMM/PX/8u6VVSeADpdjabYTyAAaEIBmWHjiXVFRV0kwUwZdoH
5Jy8v+FIphbx7W+HIXdIJSalQxp91dZsb6VxM3HkmC0e0LbjYrHlCspuy/1h
1wrWH0ZM/20oUyN9VYCBIX1xvNWVkWKhH7x5Nsa5rCVANu5yIxOPjKkQ01DM
pRLG8+dsq7N2CM149aqA1peSEfYGVHPnrt5klFgx0DUvNTOCf3n0KVCPfZ42
quhhH/kSVceijWSBfIQ/ABCVJQAeMnbx5WWEo4AfN8cXSOJtJnU/Zz18+1WB
f3WeQ1Icbn4Cy/XPUmEOZju+MLM64kma7gMtcLlCJRwBL5HzAdN0pTMYo4K1
t5SoyTRmTxrK/1X/ixe8hoJmVVv0arOquZgOLme8MXS6S3OhHJ4AjKOoOEBI
3Bz9Gf8esHKp33+GUFe58xURfjkQwpBcCrGozsKOwDcmIIa/Goo078eaLFmQ
ZzSrhUTPtfVUZaWPUPKnrP+aVifRVCpC8jb17tsgDOtjrx4yRCKYaeHI/j+V
2uGLrQnPf9V6WV1VZ5uv3xGbkb23gL4Up60oO+YUBtjoCKoqGKXh9pPm69fb
1JTUIOfsC06T7+SL5oUKspQGrX0YOJX3iiWY2QoAiB1IsS2jl0dD0XCdlNIZ
TImk+LR3BT+Wr/EJ255+TECDD1VSFZQV1Oc5wC7yZBBeL7Gu/R+t1zV8U4GQ
gUZ1hV6qy1iBVzdQNKtGcGKMAiPb4w949MaZKwncpd91Lb4jrEbAwT8J3ZfM
EvhXt9tRues25M2tR/CducwNJQvaSN/Rlrptb8O4Ome++lkqvagBwnc4+zvQ
uJmw6pelGrMDZz5k9ZeAwZ+VELKDZYr+LDVDAlAvGmJ4qtMCYeinSf+VajV3
AhK63P2QqKDrcWbdvup8kAhfkqISZjtUwnIgm59NpERsItd2lGe0V3QGm7TS
MRimcjBvg75na1LLywTz+h0T1xG6raeVBONl3SiZknAahhYHdNftpaYJ77at
UGdte15dlo8XS1RyvuLYiKtdfTnmEuTtjDpTq6wNhcN1CvEPObspm0//hELR
AAIPlLpWdAAaRf+bYcRY0YYQjVbIdwk3lyJEEJLAoB5W4LXX7ghzmYcvCYQd
iRmsf6xI/PhoWW6S4n/o+jSfxZfkKq28wXt+hN6jOku2YX3qR0KCG+y2NqN2
uJT6Omb3/VMJ5JY6gWZJI8QjLnECswv+1pZp5G3s/RD+3eEcVuz3xHV8ICb5
HpninqLM3Uvl/nTdoTqKNpAWoibvQ6cO2YDf0jdS9dYcfkwe+CSvNKjbgOjh
nrp5OjwV+DtskT5/7y7xHHddcjh5g5J8GLRDO6uXhxYJisLSuLcDAlJIiN+b
Jkj/Pomufpl6gGLn/KdpSiMt+WMqoTmjg23W4bT5EpFsyDfXyhLYK2psEktt
lsrv4G4sUQX23qJ4Y20r42zlpNEaFWRBw2Ch2NGid5yBN1e6OikI0K4fQ7s9
C41R7LtZ4RxXFsF0Q53vW76xxs9MIoeTNjfF9lyuPFFfw0QzX/lQrbSnBqlm
V0hoA2/WEWBa0+36x/6RxTIvQmXzoBWZoVAXiA/L35IojbRxr1qNpoSIoZGc
8XleW4Hl2zJNFpLUSLmdMFqKyx/BAEmaxkJMhXnfHPq0JlgUSDD5jnch9GOC
YSnlc0Ke5ME9VECdUfBOeMuiJIYCGfyST/7gYhSkhe7m0ArJBt5HqsaNM+xx
WMrjNxAosgcDOUu56hSCZVSe5eKXDFhqfCnytA3BeXVolqr0yAdf+xH0SpbI
QQ163x4XvKECK7McTQvdO2+DLl+F25ENhxsiPkCIIMV7iFu38uWwTaSgEZWA
WlT95zfyEuNTtByNRmXNDYsI9LJ2l/i7drYdY2KC448/QtymUNKDv8QbzaHr
lSPe7pHIva6kv0euTbvzhhSrBe+CbQeWgniHdjPQeG92SkQ3uuCaV5oJDr4v
MUozGF0GCYw/zaKpg1tWcV82IDS8sp2aPAfKZj58wKnUGnoCDzTyf71BrTCS
uYuxzDte+Mbd3p5F/22kUkek1+DUM5+PWBreH2qy2qgX4Z6KCRP0IjNJp13s
WNfSl2Xk9wQOTsouUKASZDWvnf90O8pEbezJ4f/XS/SuvQwHfM4Btf08pUTY
NOjMqDSqPE31V+Shkx9vm9vXCraZhx1c024OZHSQuQr3aJ5iKsBKj0upPiMx
Cg4kiL3A7RXJ+rOZWjhghmLShT73/3O3opMfw9JuYh1jtG0oOsAQ+mdF/9cM
5Cu/4wqYH+9YQpKubNFj4S5iotLx98Crj7q/ilyGVuE9nXrtKx+VoVTDi5f0
YDOd0fU8N1D/vizBOtZylugCrPY2Iu7cT0PH4A2UE2AwjYV1CwZyBWswTN1N
1BS4PKPs9KSyl6bGOzOi/Nx2dmpCLMilzgRHO2w5vYDQtipvDKcMn9BiCwCZ
Ngz3RkiP4BRVuxwLmSJ3wCexKFNnmUaoSZ1TuvISXW3nVjAanK/5pTdP8kCI
uEy3qyb6wheXBAMENMkkn25gXxu2117lxr4AOJuwqk5/0jhhZB5XttHfoTBY
y3nHxIh3EG8DZBh8VESQmD29SXyE4+z2P6jTWlpFUveQwTxUO1GZRNXlxsIN
D+WBwLefA2c8vz/L9SrvLwBZMiFVprM6LBVYikua6M74AzkMzO4+wRWMu+dL
8pJvwHZX7xymyQctB5bHCojJZWkyo0Jlq13PjTDLR+gLAq0rYP8LoJoZpINm
Nlsp2FUngH46+ZT2QG2iQXVq2KNn0tKU84LUqfShXiSMiAENCcPFk6o8RonK
3kSdMsDc2wNz7nS6gmSQOm1FOsDLGBhu/kZDy8JifQyODVn97mDSnfmVGvHM
X7B1tzMWDyK2EEHQHMpLrxeaV9Yi9YN8Vzo2m8juGVGc9nrAl0g6QxZWLAzS
vsSzh+DQebS25UUqwQlz6BTr8/haxiXaSPoiKzDV01ng4RrgfAuj5ZlUz+nh
fy5/1nsziyKN9rkMCkHK4xFXdJL6s5SIiC+jdIIQBD9mRb/WwkNItfU6uYoy
dg8LO1g2lAUsRlQeSpR4I8sfE+/b6ErDzddJTEFi3uX9k5UbGkXK3wYUuCHF
8PAjl9ZIuGYPo3r+W24JqUiO4UD7Tc5bXH50i6sF4ptfvPRghB5lJVypRMLQ
bfRnIRtHWIQAYaAieqnQ9hsi1prLYFCEwIwfIvbnpnXlHvAB+MdnMQzhUhOh
9fPheI2kpPZbc3r8dU79e3TcovHEFK6eSSeyBSyKdduR46xfPBKG13EIrbmW
QxYWi1vd33bdRdztkXlX0L6OECa5pSyR5dmYxlIeihOGqKy3wZGsZG0bgQ2S
d3xSArmh587TeRGR7DLztyDvKbRvN6BQu/rkCTxZzc7FDflpS91KqRaG+WRa
PcISzvaKaSfDiURimSqB3VaOvtT0sdPIdhVuyaqJJ8bTQ3CH+sNeTFQA6XoQ
xs51kU5QpFkO0udCx7nTUQuI02sxQ4NM7KEObFzkr6PSlP+HCSwulC7jWuqW
gcHF3rE531h5xzXYiB/6Gi0SVAGXvfDxggMC4ZXQyHr73pEg0MKnprC0BBAx
CjC+gCJ+6rYQfLbKa+dWCF1ZVexM0/9H3204ckrlfzaEktkldqVW7zdcY+pZ
dJvM15HyqyxmlPVvHnJkVahnJU5Qp4GqDDpgijMPx52OwgY5vBN7Yw8rdOws
b5Ux+Wteutucu7nPkW1E0c7s802DvXdb67SezLkhmaSWX0insXUwhvrB1xzj
16Kj4IrbYddubQ5m8GqsoOniAylbHDwBb2NU9FqWYTzkKSsth1pQnmwYphpx
Tf17B+TNnfffM/jmR/qH1D0U/znrqfvIGalZ4v7APyB3j++XnsJoPdX2IOmo
vg+EOdSKWYNhlETtNyX7Lm7VHHtN7sXY986iZek4CRbTX4uei/sKo3tE7P7T
ToVyjFLMITfR/pmlGM5qpBd+4i6oqeFTnwTpFvIz9eE0OM/4lIT0CdXeFx8T
ruSyk0Nvlss7uWjFiYfFH7rGk0qgPVOCu22w8wQFCfSM/+3d+zwMDJeNWvwo
mNPridlSE02PJ/TV7ZXzjKyGtWW/kHX5/Y047HVof3XK9ShKagytb2RPuF/0
iASJDbTzYvhr0wVU0CmtY5bBkP8pHMFTRfeJU11w+7Bot2DB3N27uBDZH/l9
qNcIhj0O7ZTQzM6v9YoDJlSo8xsnlnmYJSGBjHFtPrlWvNW9+wfzIY54nYPm
h/vY02N5cN0ZT/iaCiBlUgQUzzJFxAcsl4hf+fe3NWR++LAnyQz3L5tn3aPb
Ki+wVUfrh3pnK0HYgnuGQyPYBKaORdGGUAqltYJ+0S+GikHscC6ZFWpaaGaW
wih0l7JnHwZSO4CPe/AC1TR+WqI7XLbl8Fwpjq9jq2WxUXcS3f7zNmewZJZV
NPAOJtKB0qMdo39ydcg7SRSzHCfr3wnj9xQjM319/DrlUEi4dnLm9Nfsn8f/
keUjcFs26Ta2tr1TIc+3h06bzHNfp3A3LrLtESy6Fq1DKHkrwurwCF8UuuhQ
gFDyjyLFBGVdd3ABZNRXm6vcHUuh9TWVBVap4KaOSRH6IjiwX5KhxzvFvaqP
jrsvzZgTeaPtVFRzjIGcHrk0T3UeeNyjhHWmwtv7AnlsJ+Yt4+QTQRFZhoE1
z9jIlRJgSxBv9ITF/+iWmGgquDE3XDpQHComC9xlSZbRL4svfyXPtIcmPzHA
Uz73P3fvLTLmw1+rc07AJ5/OcIWOCsnLubqZE7vWVkT2V/B9DZ6Mluirah2w
9PgRin/fK+rA6sBZ+KJrmTTKmMsvipq8aKr8Dn9kcOOV2tSZQwdhVZZBFM1O
iWja8j+4yL64ixGzj5RWlLSIYAHWEpoEzfjYBzqK76lZseOVtvJxjQZrW6HA
LE+pxZTm7sPkTLMBCT4ktOXLYecmzEUBzV1TSu/cgL5RP5LSjEKpu0Kqcmd7
NumXV1PHzo27U0c+Fwi1pwZOyUHF8+8+12vjIaPoMFA7qNTDn7pMZ7/OvWwe
EV2zDvnxInlKBi43mvhM8wI8Q0sDOmdw8GY3vkLjr6Z5BJIcgfTQfBHFennr
+7VgXzL0IsmyU7hR66N1a9do/NJHI/79lDiOYLjXU+3C6YdJLY6ZIDpLAKId
4MTlNsoOVZR4c4+DIH2UxI6uT5l2iJnivwU9mG65YrrHJ4vdV2YM6VK8degm
N5+s6weNePoaWMw0fGPlc50bGQCD4OSMXcq600nsj8lvGDWe+rHLKpwGbV5u
wx5JKasquCms8rrnjhyDJcenbQBHWNBbGM3HS6EthrCjk4T99aTHI6Lb+dt+
f/azu5AYiijCZAqsdzFhM0k0fzUSGuIJp2LS3bk2XTaQHF+GtZUW69NyctSx
iAyAoFHfuC4PGRPKhNNKs64W5bjNu3Taj84Ml5KpRbMNT13d32E0w97bcqV3
OwoIXqmtoCxMJzyz+guia7ntHpnO0EdTiGjzBd1pRJLdoZeTrllEyduyF6CP
mzuERx+dVJxIKI72eYdUxbU+9ZqQdTpC6k7QUR3o2DPNH6Ul2xL1M2635IHf
svLDEmUqAOEAMzDb+6rNKqaRzGhgpBCLSOV8S1RDDBAtnCvv+3+dNa2G+Hg/
4dU2b79jRPL+nVvzIJIUrbmD1lcXwmyk2wDLNSBio2YLvA7m1FrUT/Cy0fTB
wL+QfP8N7azTO8RNfN2VaxAdGD20qkDnsJWcoD8UVsoFxsz4Rf5ktq3JkAmi
sZJNDjz4MEEqlkjro/xTwqCzLcPJYBTbC+JL7ywBK+V2xuUd2CPQCYqX0j5Y
1OE5k4R51vI1Z6hE/GMPkHUaD0GtjPzvWPhneIAAfDLYObUzfJqN7PRhkxRI
YZ5eamkEm3//zP5oMoPGYmCDVk9Gv75v5nxIzVqILTCUxu3K93H5XwBM8yJ1
mR6y0xcc3ee4KLkvNKi7CutkC8lMtz21WcwWGGdPIaNdeYQP+Ate9gAdXBD8
pZSCRZelza65yebrR8zRzTHCSQ9MSxMwNeF7lAb3ULOABXI44ZAcJ3Woji92
gmbtZvcqyZBQM32WEhBOJuK3zCMsJdvHZGLOJKHqr0yed1mV4zDZwic0/3kH
hyKJ4p/8pu0WKJs6JcgWQwSgZKxOQ0PPnJGDPKvUXsb3mW7NajY2NR1oZ6Tr
hlKRmAQaKCTUN/zAKJ7o8MxShs4PDliKK6YIa+C4094h4zLGMsyV0GpT0FOh
9M/DhkoREp3fNbo1InhR71sJD5jDSLubgyYuVDAuQOe3r2LifnD+UKISdZDQ
4luPb7Z49lzuBoDUNVyFgXDpV9DdDjzQXg6erjZbs2eqQT6aSjphhBGXrs5M
KCC/g5AdR0f025lsC2C+hZMMTeFA0UtdU21NvbMdJ929PdMeeutcjb7j6u/w
hMrkVGmcIUTM0dtr0HnnrKbymcZyDmPGDGTNCEqUfhpxR95/5UDKQx0I175O
xqedUKTzFhgh1unVH/YpjrWL9fi1PmJAYCfN1JAxfPR0Dl6geQnX9LudSY/S
vngAEx4LlyaBi9b65OMMyeIaOBixE8w673Sf37kvIBZQG/N8QqPHWvAW/V5P
MJg4mxZHIABLmqcOzSSQPHA2CFWcep+ffgdHkiUMQFF8XJFEICQvCW79DlcW
pTcXf13Yf/tLkx0zpiu3NLkfifydblrRAZ2EbEZboD1HvUMDSet2NnakIRfa
h8nwjvv+JzjkBu/573V7MSpM/mXm1/78+oobJ6GUtjTxHV+Io6DFc3oeoF0H
fWUYD8Vl/zB5XzIepXoxT3LKdJRPqt9LdWcxQlf93oQDq+3qzrq4VLQUtfJm
BBmVY9GAhyqRL5OW9wENdlf4z+cXzBlBqE7LqcpT6A2dlmhVqI67bWBo2sMN
0qn1I/BIC5uXcrBXCnayViqCYpvPkwWPSTinmhqjw/GNtaIpBAQ7fcZqyM3P
Fqpw4dzLeZKzSk7xmplWmwekI3/IPTcnaCTS5Kh1A6JcQbzMysnsinDZJePN
ov8sBhdSaXx6TDzhBv6DFttLrGxGGWzQx+Ni0bXcfAYNketdI3TSzxw14kzY
FUY8QuyAW4bvJ2gEdX37IxEPGGXvPTAG8S+Y3b998KapucIN2Mc107ppWS3i
/FOyTrWlOtOjoK12NYvMNk8pU0q6mUZ3V5dAOuDTCI7FYSLNequWGtLqG1/s
ek417sIypBlw/G8oFb82ZXhY3fFhdWLUAwmtkZAnkBd/3BuxTg8H02CCXcoJ
mCWIRZ8anEat0KistFNDEOotFe/LA3Tn89Yv8j80enTmtipWdZjVBzTqagXa
5Y2TorptLgFkD4TEENdZQbIxgW1dVvFZ61JdvO8ZDO9M8Xf69O6zyfNTKXcr
EB9O8uLF4vl75YnFsjWhxU5aTLEAdsqkyZM8zjt3E52yNdf2R/MSc/k0aFVA
A4aOFgmqF8Xe/3DbBkOd21irxxVV43qjBVnLwS1wD8GtZy9CSRaoFxUL9/9K
Ljr/NqbjO0YgXJNMpgIAaDij2j8/vefEo3B3t5A3wKCc08H873/e9zzMLCie
YSLWi0Sqc3KRBMjsmV+iLhCxUEVcyXWh5JkmgOq1eorKBlcyPIRR83Acy/kR
jgY3r/3Jc2aDYcRmLE+qt27dVBZMCCu7Zz5limo8eGBEm6M7ua4lLvZfo6Hh
t0bEWocsAansW8EIyMuUMRLW9YPdeZP3UE+zsi/eJC5lGEgcJd4nXzDFVhMa
usSOmmehTIJpd4OH45fflKvpOi1cvhqqsHBE5Tv22Ik0vH0QVor5oIBJUDgM
zcW58eMvt4BvkpQLT3LYkyQfNVFYhCHWbbD7+iv9+Z3cB82DiHsBCvkd36a5
wO0Atar2jCgPSl0Dqgp9hdLll9oTsTNTMlA7qhksWL7iX1S3DG9mfXJl4A7Z
UpGQ2gni3//jHAdaK5lls8wib5NF5wfpxtbEQQdDf+CQ07J1WZDB/FOI2Nsy
cE/XaYX1CM8gWJl7f24P6Tv/qWeUcQdhp0WWnWadltTWqlPJ/9hNQ9hgccXq
ulwdGtVyDgl9ropaj9r39g335jcxP1Z6JlL1syRWHO4VZIZFHRQbwjkRS29E
8NO3kuB6DnLISDMxp616d1LaC0GlmnErX187Vf8PYdc+I9fZso/07rcoeAac
+d3cKbdQ93cRK+oUT5rt38Spm87vU6A8mruJXaG4YrcCfTAljiTtP27vklfL
02K4cqhaUfzWx1PS+SEsgo5lcdmhohli6QZ9eO3KaB8fmuww81O5f+RLC+VE
64QGFt+ZzTNMtMWUVcs4jgeqEmHttCSB/kBaY/0HtW48rRfbi9pCgJeLfBXQ
zJuexQBheKz7PGrJL50GPVJK8J6T9eefkWi649SoQK9IzWSUGr9KUGMWB8ym
kJy5Hw7edZKzromYhLu1fPpg8sefR0+5zjzqnOxT4GipK6BUAib9tp+4QUCk
8MaXJzVbnOBe9X/6bXjcMH6UC10RQhOHxIWMDNvlzXiKMzr9JgxQ1IIAtapG
b8GmGroSwzK268WfciArVxPCi+Ae7uBkn9qPdIQp+9MJw/AlOHl/Y1H8xhue
QM/PoGBFHHP0dzzP780nUTvEWoRuK+9gGkWDgMXFupNzt1UcPulXbUp15EY/
j9/FG1bFaDc0F3Fgoia4+d7ZT22UkI5sc2F6zSyreCMePQcRFmxG9jdW8QXp
7pZYR21oOWDzT7oiYFo8H0tU0mLZ78jrjujM7FG5SYa8wyYgq4HM5g34BKnx
FRpX07IiU0iVaJfwrEgxAIwAYXpvuSj8NUhdK08+sEyWEcBabrRivRFLXi5M
JQQskJjm/QO0p0giMVWZ/u9hjMe6+uKbODW8t+VIq4gMLrIc9wQPjt/nOaWS
W9uO3HG5XCjQxdGVBUE+dP1HJJUrM9gyOJJL9SoOUvw8EQuk1QpAXnUvqScp
flj0enBb1sVYVnZMoknvVk6Z8SpuqOjT3adhOTBVgQYzIVpPe4HyOWEW65HW
QYAE5mZopbPBAOb1XQET60JhiU31XFeOLLdbNmaB6/3yem5uKtGsw/vmmewU
L7T2QcwA4TXZ7DJJBq6By3QkpOHJnqenQC9t6z7wuImNT9hZt+LxVCZOdEv7
0dhPcBElYd/rvp8bD4l3UiKaitjNIN0PljKohxZGJGxGjEMYAi+fms6DAXVg
qGMjUqtAwhva5XWDhyFyvQKdaMNIPd87+OA6RNekXozqGR7iGmjYyGQqI5hw
oUDYThtcWpUSo+bPWI5+an1cD5cvFm0WCccgceKKDdVgCZgZPBp8LNV2sdnC
KeJgqEt0IFAJUO/IgLQe3eH8WcncTspjJlcFCgiG2gEdWn6OaAQ4nttdHOcw
bMS5lMnhs/EOLmprRVeJ743Y4P9XDi0vxvBERp5xqDu2RrIP5AsxCGASI1l4
iI2KfhnLxiLv5jnzx85vW7BlYk3bpxcuZTf8dyBXMpBgG0NrQ+1Hg2xyWOOP
ekFGPor1nE3UJKF7Acpuy7GJ0sEHxDU9ZA03ZrIXre1zojNE+R0oZJEbiqit
2Y5JXQLbHtYGrDIQ01YzofPl5r+vEYwkJr0Vx86oF9GcsLAO4YuCOeeYtZdM
9O+uXbMLfFCs/6Li8BoWMKRvv67WuOnIGR+kZmX4nT/i2hlmjcY65LTXS3nR
bo8CryacNxkFAk/DU7fcufDDNZtoqtaKXgaid5eekHpEtxTBpH35YHqOyIY6
AT7ukvUh/ifJQS7rRpLOZWiGrVdfXKX0EbtFD5r6NVRpE4OADsm8oHVqLVaF
rZ6OPAUg8GAcrMq3eted58zk50Em1aHNJw3GcJI1KQeeFMnAAkT+TXod7PDa
HaS8CB4Hww8nEx5JcPFVzRIxQBsFnB0zd4g9x8GPcy5wTELnrn8spiznYEGm
qvcVALDag0wDhMrtRP9zI9dA+RolVXAtxyZJDMlA+reHS0UNc7thEHvFvjBA
6t7iplIhgLZC5GlcdFm9LQG26irfid4D9x52Dn5G9/3DNNSPFhKn1yKW4934
K/8K2ll4iMpq5XanhBqecqKXXdD5/CjEdmIHlY8Qk08y1ID7tzbeNf1jEh0x
w+GVDE7P1pwTP2ntspak3Zm71f84iyOPiblxae/6zb9OmD52whXQEXlbVohB
+3Aw+e+UQ7Vb3GNE6Meq+DRfi5uIOdXNBxIMvaEMcsD0LVTQ2jOJHIvAx9ko
CzioKtvBJuon7YlFmQHFf7ZSpEfbmdrQoFWP3iLRDmhs/6sI89oZc4PQhob5
FZVqIyKSL0Z22IkfXFaOzyChmJo+r4OcHp2ErfG6u6A/9goWNPTXireb1bco
9dTRMOGpLKgs3ezvxXc7LtVI0XtDVfAJjpZ1qoGFziqDttRvFglv8Y++GkpT
jwf97tA/HcIH6M/ewiUlCd5n/2oLGyFa8DLLC3eGcrdIM0wQl58cYl6Vfz+D
OgVJ84HRR/hrGGMHL13cfCz6sc3CRonEdx92zQYO+HfYXXWHU3hNqUa8rn3g
DuCAH43mnvAKOdG579CS80kCchDDazgA2UK93B4OFjHKGom9o4qtzRFGV2D2
VnigWPVBeGRhSXWpGaM1C4EaKeCOtLhoD9U9K2oucn0Hw2ttbxzRZLKf1neP
lxHTUPju2TgL5+bzLwUDam+GckrcM0Uy0PME+qITRxBaLlEQr2zpstziNvGr
JfnJEQ8MbCw68dijToc4rtXaaDq4bhUIEIfo1hHuMibvoFzDFTCs+peQdUjq
wljdMTwMQmwu/DzF9gZ/4xRy2Gu7umbmQooE93hN34uQtaFkNgApmq0MN/tv
ZQbb7+K/sCHYykCFukkkppHlzlasrWHAZLyJUeWcP2LVeb43e/rF65wi+qn+
/63nnznOhqCPeaF5PCiFoBTgmUsYVRfmDqnCUaI0gv47NIgvrpMAaSpx+PMJ
o5ejXLRPk1RxXOmCeyS/43sf9RBJMOmHurLBnj0N6Pu85eVhbzGAHm+aCSjw
P8zyzRiEweJE+VLAu49v8CkBR6QKKvidPEq0RHyPezsnoaiYjiHO11OwFAXr
XmRrhVx1syoo4n7q2EAd7NRHRoJmR2lqBvp33w44jv+DPK8608QU3G6UZ9P/
TEHqRT97n5o0+qW1g74F/vO37a+IBRuPiYxlGgDAlYaRLmfLGyFWtn7voe6o
dMJtvuLXfYNLhQu2fp0Bq8oQwB3lrfotF3PQy+XLpRuYapS1LkChrxkj1kqT
ULSPFDfQ/0y03Iav90d8cbNuTHyYKC4+Mj2ha+kdhYmHuJtgmXmiVct/M6KD
SffVWe+/YY6tA6Cxw6yYgLF2QvetzcVzuuBKdIYavgnOHz/Rc0sXsqAiF85g
4ZS20kcDhb1V23RLBOgf9m3fTHPih2UFkc5GJf1QAb0jHZAQjQlrcGCjnlw5
QzNoDkW3J27I9NBO2dgpa1zNF8P2pSy5oSNIMchSR83FZHqg7+AjutNUGfvB
CLEgb8RazxovvQse3rGpsahkBQ8vpTvSbVwN3DQqJEvCxkJghI4WKUt6Ea+3
OMZuPGrinMLBr6zNR+0MEtTnMNIQjlt11lDjJRjVLKKtDHuwrY5QaR4oplU4
bWnrNfK9CSRaWk61OsdzKSAxsb6Lx5+CcxkjEMenK+n+F7pLeSjYBlNIfR0f
WRN77NqX1hnOCc5rhLyR6HX3NCux1nrTcMBlsB9LpDMQiu7B8nJgbB1Mgcor
EN+7JPzfRFXGQd+7EdZEjqY/Dm+n+w+kffVQWn6d6Ol0yqQ1RrKqmNVBulGz
SpIhM5IPmSFpfyW2+84vLJJvfPJcoyEU9G3FSx2mbDTXfyC4ueAPJ0Vktogz
dhaBvl5yvkXmLgxiYfMH++uPRm0w8TqeXds1BM7+uy0lZbYr3uWinVAlA4ti
wcGInHmh5uulZ0gkccljB577pfc0oavaEugXmbx4Gs+mO1D/GyOq63djPTXb
37R5fUu/lkQ8COwGR8628qKIfMJ6uD2VDJg2fM2Mbi8quJX32CUglvB8XOw0
HE45D8aDP9gFQjOso8qfqfhCOHzIvZ95PCPL3XY6ZqqsFjEpGHAVkg0cBZaW
ltfP3d4s1lGK7iD9fZLWCRNDDbDx+N9KltVtfGNasZ8D5F1PDnAGGSMpFodS
sMsIpvdyKt0jms7Q/rXojOEbeJI2cAV5yNZjCjOD/80x+RCkrQdD1x/su0Kf
15AmcEwAGChZrXS4WGDagV1lvkB6evMSxMehehmDD8tjtJERx/pUWe10FJEh
Cb3lsh0k9ItQa1bFg4gUn9+gF6xWT1dfP/SgViD2hl4STfqwczDKatwSDgYK
F4CZk8Ek7/Y9uxSoqbMBz3ohjyz1OWIypo5a1FM0n8rPYW2dtnXs8ApJZUon
WA/Gts9Pe/qejI/54qhVVHYDYJkVAD0hylOo5BwCaR5xQHzBiUGFpuOV6L42
sZZb7E4VqZ1G69PIvoWR3n0Gx7V7uFycGPu2J8iyuzlR75XUnExlZTo5GB8/
PT97j0IZDmSBw37iGfs0Q6SOtFznJNByT8UgYMvwvFJXwBNwLkBw7C1Gz8Mj
VTQlusoSrUtRCyl7kUzV68UVBM3dXnrLO/f1bOvgCEOWx6P48ot0NKbVlshk
HU+ghxq477jIxuS1244bKn2vUl/ZqqGHg/2KR2Ryr6tME140YTbGiv0E8jQG
HuWevJ3V3Dj4hkG8DZrnj2UGLw2HxnA/7F/HMOF07PQL5p3J8NIA27pQ4LYh
XdtxTdPGPwoIKfpoxdvMZswnakZOjANKf2vty2acXHEchart5h03Gnv94BnP
PKi81GnVdIEkzh9yNgVyHVKLOuCsiFNG4Lk628sxDehhIfxc+3vXMXAzLcHU
wlB+DilBv9AKcrfa57p/kWbt+i9VajYIPazBksOfTkEmza1UMz4JeYPNoZf4
BCehARyP/INWG1Apd43xDYr1G6ce0mcd4lYP3BNAJgXLnysWHWh/87n6fI/P
J4Daf+C0uImB9vqnmwCVoNBJ7HsMo9sEzAKaRIBmmPgx+B4G5B1FawR6k5or
y+/miq5mhm6sZl+SKc8nYVOLRqpu3zHRUH8wWeHwxsS9mD3u2K3FmpRQgvmY
GiynSf+1zLAJY8Ky1GIpA8tqZKqfZbtz4e1GeS8fW9DpgoKpoyQDdGBmQwKz
MJVUomqS0rrEEycTcr+1J4cnWofj2QgfOKJPgy/gOgD98GK+GHbYkGKZ16ER
DGWE15Er/Ec5wEWRxQNSihgMaAX6Lllwg0e6Kfr6hz1LriR0kkkvTyCTCMh5
YqyeyJKLg/LPNbVZBQYAohPQhOlS/VD/ZcccAYWDVex00pHG5l69DAWwWt5D
ZnUYU09fC6BtwmnLpg/aYuWyPQw9SqCmPcDqK8Ulz8y1ucAaREP5JrnJNlbG
3RKZW7P1uRvVacH68sc/8ret4trTfKlbWihsUj3ssC678bCaroj1LaGDKaMu
RBzd85DA5BEy+s45qtxWXPIgLxIKhIQk9sPMNWx7/LanDkJeuvM30kzCUxKM
HnDORO5C61HI+s+7w1d/1/GxHwNYgtmn9aMxm25UhAqwylvEzPzW4FjJJaB9
W/0GK6FN6B9RmPHgF3ctKw7LjMEkIz+YLA/IrlqoCKqealRY6qx3jMZGRnX2
1c09WPR0CDqZ6IHTYW78aaSkEU5GbDouXFWhBk8GvkGaaCnSChh0qDFbj8AH
3/DzEQMvMRbR/f11tA2EK19uldk9KjP3oWCiQQ6vG+rgMGB1hhU/PrRmGSdK
meYKCzy7o6MaFeUnUlCo2KX3OopJPKuXtl+LE9MceEtLzWA1//+wYWe5HrtS
TJwsfSS1iepKtu8hAoZxQ4yCbxUcMK6IUAsJZy6M9t6IGOqJnxU3GqY0DZ+V
5spyv0PONpQOKiFhGpwglXzaandCDUlGzFL8zgv5cTgbUA9WnQHa0WdrqQYw
q/4WBzPTwKMjmP18ZyK0uUEi4E/0IJt4t1eIjI6k19CnPD4RUnxcszSVQlI1
JnKOWLG/f1h5RVZTAQ0rUT6ZYgU2nmLmLdmStKTMcv07BionEpYlGyWfXZD/
omSn9OYQ+8Qk1yFnDRNojaypFGSgR0s2R1AK3EGAFz6bANG9HMPesIouI5Up
3sHBePbTgLmJaOMJPJ2bqwFNyLJzD974Gy1F/QtsEbd1XKTu3x02Zi/Dy5JH
jTJY6hAyPWTRr4XFr3ew2x6eBQ6RpPQpZOcMrYBz9ELk/8wMg54NCuddwDqI
3RMKphci5jJTpLflTj25WfB7lTZ3YTt8cndrT5yVSCzVYmzofZB8LoPctYvd
vPrZWhTc5MQ2Uuq7+Xqqsp7TVaQMISu4jcFunSazNnU0E0/JQGwdsCIZ4GBF
5EtNqOsYF9gGdpJ3+f/0fmg97aYfkk/2sx4NhIt3FOJLzA0VbRc+qkC0140G
GtKzdJEf5FekGqqD1iLwdNTPnfTG+QcIyibCo1RbwDNs/FuSYoNb7wxDOQzK
pIQTPgXkNsU9+ycg5A0u/rESi//uT7FqIAu99G898Q2j2xIIAH6dmidVoSK7
G3HTpA7hAJ13GVD5uJZPqJwB6jrp/uNTgNThCkCOIYaXAt5pqS6yEZ6fGrvi
n70/znvPrkvmOMGorPxbrgQZ6REOkcAneTjxzlDdL2eSyG2E3YEuLsA0Bw1x
cZZU37MyTRKrrrwXnutQuX2Bzh2fnEcEeo4W0TDiamJedzXvJk3PnhnSYoK5
bkvgMCPXvocCSs119CUeWmfByv1ztGOk9kA9mpSVFaZUfphEHrDgIKwFy0aF
Z0Y7yrVgSXsag5mEcO54Uz7AvBpxsngsl4MqYG+eRBw/JLzN4p/G/C/z58K3
MJuDjLHVddZDJukXDV+IrlPwThuEDkcSyS6DChr5GE9ZqSN1/WxsROmr8+iJ
R6NPtVk8+OTN5DRQNnlhat+wn3c7jYdtK2H4vOHnZTOkHDai1eQLBMD67BPL
cAddsSj9FgP9Lb9PaeiPDix7aS2FFVVTzHywIICvknpji9IiEc+JRsddo3EP
J65BBhZzJ6Bw9ETW6JOe6I2eg6fUQ59dDwM7ugwZmKE+LRM80xsSkCUTSvnN
8J8WDJClgnRPDdcZ0OrthxtnuVf5yfxlgSIMDwJt5venAexCLryiv+zW3tGY
oE/YLEwTOSEJlS+XkgvyT2cPXr5Qsvox86S6xJWDz5/y1SGB5hvzoyDoBmep
wV2Jfr+a1ZCXh72+nkBvuH811v+nG7vSaIYYMp1V8expn9UXj1lfO1YEDAzC
47KUK2QwFZyyIUcZyIkM/0tU8p6NFwK1FWxye7i5Z9dDC2x/QX7gFGcexsp8
926psQXFgRZbKnn4B3oF4GxUGPHpFsO1yO9/LJ1s+WUpTuMoYJwppvRIvzs4
f53rgJlXu5iyd4nQBgnK/oiv+8i+tTGtty1xZ7VLFa1/j1q+2ymwcki80bpi
OXBoBKEfy85GbojPI4+fwaGqa0HsprczH/iLqDZxUCKzT8qhPnzrF+o+vlgJ
i5qFTo7szd417nQqx/TQB128UZM+GQKggeDmdyttlLy1ILb86sN44KBTojK3
ZIDpuwjgD4j0OHlulTabEKfsgRbdkcNsI7m8kg0vX1vYyAjvj6paqypeYxqf
A1OZ8mgzEei89mV4x5CDhTWjVqFCh/sFctQBB5ntXodGaXxh4Rtq5Awa91MU
du2nyx4FAZXdRHeBf2iHAaWz8aAZ+xk/Zgl9GxVQJLL6TQSaIHTpT+aM3OXl
tjgcbUostKFYuityD8GUupu9prVFLiLz7m4oP0Crg0wXlQWhG13lrqiXu6Ip
E3E3IxbQJNZcNz0gMYxRvEN5mbn0VNT17/M1kSS6EghfiCym+HbyosxH4ZLG
gWdKUIF/t1oFr+lSr98dXH2mS9vy2CyGw2Q+if18zjCtv56nX/HIFHOj0oXA
e2Et02ZjhntiDaGjo7BLLvgK/YoE7ZPF1lzciA9tBn3xvCbGPo5a7qR5KKY9
gUQmdsiLRDBXFLGA/UxJU0rG5WTbNgad3P8g6e9qsh4L5Nvyfl+Pns7r/Fb6
sDFzXts6ipmMNGaAXYZHJo8/bLVHePyJ+yMJ2Y+9G9fo0ZDwbgE6q3MtJQDn
hR8BVxXrvpgLC0a5Z7Ff3lbOQ21GfCfK3vuhSguy+s/3nrWRG4s+nLSp9XLu
KMm2NhG7RYpLc8nGCnNeXDFTY0NyFUbCLCIId771RuJK4vu0dTWx2OOeEGdM
RfR0JIr3MDtVc/Ek13Ow/0f35U3vIwuiM4kWZZzjDuT1Kvz+y9jpL3jGOGL2
i7IeFR+V+X5V0vot8VmTolWgiJez4ZY80aAaLqeiKCDDfpMR3Ou8S3pJbmXR
/h3WA+p135fs0eHZL1gbKJJJxq0/aCe1WO5QaCj7b1Hy7Guj4VYg1Szz77BA
fdafVq1ghZmxLmJcFklwyU1A5yVVbrQpcny8+DqPxys+ZIHwbdEoPKGccEe8
nUJvuVyFjgqdRXa3DmeX7oevYU7Hi//SZRw04+jWAs2ea4voN8bVhjG75N79
pfadQ88o6Dft63/VmmHR/0nk1Uil6ppPqJE8IgrfKxGRyTOcLyUX0+PJKQct
ioi+Mxw5C2qNRXqf9FYQwjItq6Fy4PTIUm2we1IHQ3qPD2DyIQ4X5EsFeQD6
opLF2GihQxxWR8WEH2pXUjaj4+8b3QYoaOMRRHvWUJop0MOLjSs3CNOR2vlx
mQzIqmulwg6L2TQ43yEeevebMXf6bkD3c2/mtCYY0R9NefuJ8K3OXj/N95mR
Zh47hGTKkXrwkrMTCqL07PGFPy81VIX82SlAEncqUcmX3lo9Zr56UJedKy4L
Wu97nQtTcBg2rHP/4X85kHSfPmEXQO+7YLSWihJIlj6IS022TbPqjRRg7BoQ
Kn968ewM22kvTzxalTa09M4rYRw4bK4ycnOcC7WDQN9FKUV+WWFm8FlE5goR
DtpnYP6gg9ktyV3ke9F7qaKBImER+3lJeBQbS4tKzXIFdfelgLPKZR93sbQh
vnh8bQHOdOu3fpa/Gmw8RFAWJqEXGKNZ6kVZzta7W152oRguoFbE7lhIqDdn
K+fuwmF8BpuEfM5WWYSK2ebnGODPCBM7NQyzufAh91cc2u++7aS6oA/2At4s
VqtHpVRoWGNpLHy9qO8qWQyEhIzFk6ru9+P9zkMt2mlv1MJUwsjglj3vL73a
GmsvaFbffPy8A1Y2krNylLH3yz9rxqbKZ8hd5ky41Myz16OdAEWDJvfSZUt/
CpOzVZ0MR3TzSN5w2yIoz+dhGYFxR4KD+Ug3btXHrheH8K7txVqCEoM1Pm2j
zXXBi54NfW3hQnoI7C59p3iY7Fw3CqQa+uve4rGvcOPDtjddrYlI8yMk2ISK
zqyFRjTKYK5lNUQtlQoqS+UIpcPK7i/cz4lczR6TluJyRzd4UWv07mlObslD
AyDGkXxFzKVz3vCF7Crf5nVCGP/rIDoLOuLm3ykENb6CLt/dZGVouARbyP07
clC1H5c7VB6AJYKbSTPLfjLnaS8i6vu1/Hg1MJ0ZI3mDvUxWyjkwoC0flYQb
1bunH/HYHzS043eUoFQPAJ3VItkDGEt4ASeWxzUtmoVjc04pkz1yVmlQbuQY
rhq+kGxE8szKcrx3Go6oVsb6XrnCZjiUEHbu8cdLkejSqP6eBlQp2v38WuvF
0tD2Ojlv81+DmR6JgjleW67/MvbguUr+OMc13ehDgHQDI8XbVdMQHOe9ccwg
5FhLL+dsvOllBp/3aRLCRP49naXE+OiLdNC2KmO11AbFEe/FOfa7MmA0pJ7p
MR/U54HzyMHg9om87MNvaIPhsqKNty116KLXOGXroMZ/6+hYDpZdHRewwNKZ
peMBp606TUoBmhUbe+amgv7E1r/EBg9zS+fTf+vymXx4dV0V3IJHaUtSkidd
UvCy3rI4TcRWZ/iqsSsfGAj9FzJ2B7Ar45dC3A19k+3TPSgD/npE/iaw7hxC
7HdmsTZc/+DLWbLgzCwm6Q82c1DHpXG/krYlvxVUo3u8YvFZq4WHjzDOYzhO
ehCNar45Yqap3XqXC6mbPfzO+kM1SReUPIKMsKRoc4/ctKO/fbHKQXxA8mf9
cS/ITxgCde7vn0GKFqufl2navTkie/HzjfYENgAglW13ggTdDnn0p2Y0DFCB
x0WUwtz84seQEdnXYWbfkA8eMkFhypGfKY8+jJ/fzE4zvjQGnpjAS+t+NJaS
4kTisnnU+a6MjlKZo0It5v7NwhASvK5xG/2yBVC+hgqk7I/1LS0V52nQ0mYa
AFrXal6TsIf8Z0OfqejL29LeObaI6H7GFNzjHc35N4kS015+7wA5O6FZxoJe
Imvt8B+bCFSIQrL2BF/J6v0k0HUY1kVJL4sKSpcgtH+HJNYidirejK+Ru0B6
fr+/kl1Ju5Va8z/8CwwPcutRU0IKXz24o6LFCibGZE60PCcRdQGtpJCp5oIh
IXEmDUblUfTjLNoD5Ev4LyGxx6uwAD/L01Qa7ytWWV0QtrZAx/y17Rd9+v3y
fad85TGYfDd/2fIOlOw6Pjn/gUlU4D3YPaDtSo5ZteUlvZir0HVO/nUikxbS
xrVXoi+ULEomspYGlVpBT/OQ90JoyObFj9zgrAuxgbDQmBr5XP8skivcYaEG
mbDLUGwQH2Zkk9F3BBO+whEPCz6YFTU4O7CKHvE419ikZq2NjWPJvzrwCDeQ
vhqw1LlxoDWhfNMQdOeyUIBqwAb5bdJgWpWtK2uwEciQeRCy5LoA56R3xdPO
St8+UlLtKbEQl0a4w62Rj3djy2uEF4oHJGTxGClLKi/7RfojfNvh6qrV9Y1G
QTPEmpCM3pPt5fxlyvqhA9+wYZmG2lYngh2za2VCEH9IN4groi9xL6x5xipf
BWqbuHgVgwUKVs8rJclDY39yeJb5wefg8IC6jUDfWZOOf963llhHYm9eGINH
F0UCtVckBBkKkGHNEMS4+kTy1X1D5H1TRuawoslrsUOiZhY9kFewLxJByDsJ
I4cIB//Y+mszWPshzqoEPFQduloyBftElZg6bPI7smRBkAU1hcZa41SCOEPI
kckmvQCFVVkoVxhZPocqY+xFOK19uVWvhC0fVRwbC+C1olWvvJHPpjtX6WOU
6fjlv1UophA00IjZzG2FYtnNzqxVsenlG45yIV6fYfAmi+5KnLxcQs5Ti8VZ
WUPY/6xDhQ1/RKqDCB5Dt/cDlhpU99wHXqO4uf/bpE0ySL+I8/eIep8Ry7tS
APY0AmVrxfTOqgB8Zpn9fO/88rVM4dkZw+xjQGfZgbcA9lqpL9F91uCBnANq
gVOG4RHd4lqENm27jWwwB5HnPV49lFk6sqcRnRJEWEk9ZncIpfnvteWbBpaL
a3XxJ9HUGt7BBNWXsb885R04XQ9hJQFQb+zblOx+6bNu9Nu3bqszK0wgBIcu
rw3fk+ppjSfmarxfDsZ9VzuuR5Pq+rOCfaLmPMhV4/gSlgFSUw2P0lFoi3F2
uWvhLvRHgCxxoFIR0dLOILNJWbRdyDzO5eGbvqXrIH/daSusrAak4yg10Td1
VhmDq1UP2k3BrywvNGQZeWwKGbgA2nWwrlB9M4H0vz0VxOid60A3ZaeILKo5
XznblrUMzC5tCGxzFParjLWGDT9LQ5Yt94E4clp+ty4+FvBeAWEH6hRa/AL8
9Kk7gyAj6haVmRo+1Z4wsvImuWcgby5P65i5qghc89fXcwNZUkWhhhQZInfx
EzU+RfEo1Ai1l90Wa8UQECm0qo0VC8LVx1XIrxSYs7AoNkMhEMhLRrVezBoJ
dNWqo9JzvamiPfkeLYH0rOq+hobeulxrfn9+XA571SS7oa77xnXwJbwlBzJ4
cYLZmepjwirPZMocKUMnQBiRrmxtMOLSZ1OFaqCioMmXIEvt2t+nRrFhAOeY
cFuV+LAJdBU6tJViOJylsq5ZIc7igv0BO6RcfRANmfkCmxwtjYkUNBmHSgmI
AwmDjemzR1BM+nK9pQyRNSYrowb/w1ziMz6W0Jspe2m+1lDFAKqwyCbMFkvW
mkXlRuEayty7wFPut1h4exKXI1vppjwnK3rSXvnbcK8nMCYpwxxXLThna869
rGxzROEOez/TZBbzzSF4qeeaS7u34qgAvT4IeuerSmLipPgVl7NvQlP3CcWv
pBEwHb++ZRh8k7/YYo/knHK/vSwjpjXQ/guMLIOcIlGK57Puyx1rG3C0RQch
/5HEj7uuzkskvEoO4OD8EstW05ySqlZREvgpPujqcO7ULIMcWIuXCUclg2cU
MVzI43lMy9HasNlOxqjayKfo80HrqqlJKa5G6DPcS75lcFUaam9lMLa6v7dv
wPLo4znyND/2bvoTEKDGAYirt1g8GtScjPTfrQwQIiAR+U72Kyj+Es5+7H1t
SbAj0OgfNzpmVYu4lzgeLmXqzoD6rZJ4G0xqLhedrMZ1I0WdQGOP1MPuOQac
OGKetljOExCln/NwmkVMqaHtroegVdYb6jOlwOFLmVmoodTr6HMMaPMHnqaQ
x0tjDl09hjljHCGFBZD3+nl1hT/5DNGZ3xK3gkz/kXQoswiYfgzo2DE5wBxp
fTFl+KzQh7mP2doolKhaa49XNKgLsAAJD+ypmIvDgAFEA9bebdrHEwRXxEJN
Kx1Up1t6URK9+GaDFmp/DItesguP26N2ubFyT8Scx0jB0O2NsUp/vXTqOtRi
jNclDj5kH1eFdoLxpruhF726ulcFsyiA7dXTv9v4w7GMl69YzWPOK571egpj
t9bgfOkUIx+w/43UTJPYCpcfggK8vMAq3lNepy28EODOu//5JskECZSad1Tn
OX9fQ4btkH+35YJ0mxlpbtxk0vaUtPSmfUIqqZKoB/LIcJdaHjIwxgo7lWjr
Ldo8qrMdgP9x/nvGVdAxVOCKuAlViyBkBZK8vRCvYeCShMjTso9SrSYbidd/
7VWhdsW9FBfVT638IIfkxUn58dAqOF2va4rEPYwTQ6atpZnqIvJGlcW5CLHx
OKtibviR0ua/WsioFO6li8TgOoKhMRl/hB0jcDwEYHpBC0nqXSL27E/W+zBk
JiRf7zRuKmXaBcO2My0R2SKXwNjIJ6ccqorR5UgBchtowGXLRPkuRFZdqsW/
q/Nr+7ZbMfs8r3H2LbKY1ldLBvpf15+XVpDu9kmrjnpPuESeI4g0S96gRm4C
EkbCT9BHZBuOQcMOcEJIvFBBkNLbyjzkAb35W6M9v5ZXPaYt9FeuL7fuMhDB
sfWSZs1s6I6DOFwxjqpHPLVeqziiszRAe+mliXIi3JgkAzOoSj7es2/mj/jN
2ntlTTY2nQqztpHyCBpXSrg6+qRvrgiF4Y7uyqygxih1BtRJdJo12KlY9xub
gQ1c7/tG0QpYc3Tk0TjYa247JAMyy9CUCCf3kFGu3v6dwk/hmvVo2sX20MpZ
kBvVvd1qozEXS4cKvhY0SlOjqnLCQVRrGFByajnmIJ5vr4wjVUDn4udgxWsc
12tfNJ2DzbrcVwUct/lStew0lOaxzZl2ytzO0lRckgsStaMkW11IHnwXlykb
KcnP3pIxBAVZ461MYbMgl4Fw5W39Max9ArNpi7NcQrVTuokdfAqJcRHKNB1Z
/GwYKAi0KHyDDOIg5QB9jFqFNJe5JG9RS++UT9pMiEP0US7WDQBx7KVP+6iI
euf0Ew8Fab9bCi6quNVbjNuyST/N8OUK2hFAHo1xZsiqCvvTEpFwmH7fVd3J
jI/Qi6mVX8xvEyxbn+LxEIdkkrYuzjplkxL8HIAMJQcGYNTcR3a93U6HJlXy
g9v+xF1xOMisRIvMBtaWSVbBnj1zcu6i0rjU4OKn0q+fRaFeS4z+E4Mc0cuQ
CSl334iw0qJWnCQ7z9sg6yk6roAbrU9b/jf3NIYPrqg4TC5X9tMTTiXCdh35
IL+Vk5HWxEOz/BHeeBtYxrNOFdqumptsgIl2yuAVc/udjwZFQX+t/Krvmi8Q
J/ZZTSD4thilOiuqTj2CPRxi6fOMPolaZ/SEWqd6LgUbbHFsjmKHxs0oMcrl
17G4UCoViT8oZCza0zM2Jc7X9/jndnTD8qCxFGmudvdhyIy7WUsWErQUOpjz
ZC/ymYTlWoTe6VOPyhIFukTY3+UFtvUQx1rQvvNCLpFJ2RO9NSY+LzPNh7rf
miRwvIKsffFEspOYG6srIaVuGPWkFX09HiEHpEYncKClttWGtlE7TWmDOby6
M3E7iVmHKuz2a4LcT2AHOugY+arKFUaJ/wSi8578Y0MhBSiMBpjUiy7fwQT7
dsadoNo+S1Xa8f6uUztzCrQ1WEa+M4lLHvLe9c/mK7xiqP7HRVJG+1B6zcWX
xQTkmFw0gX78TVOhwYZorpyjalSP7bwzTivo5Uap0CRD8sYBdvlyG8tLlU4k
Hqxxq3j8C1T1uhYiDU6RVrK+6MDTE/e5VpPwLko/IjgqvOKnV/WvcnGLs/YU
NIPYCmS7g2q2syYwM2BrOmQJszVBRV26/cbQZdA5cSt+AGZAHAG+V3AqZ2Z9
xBVpnVCHnVwyRDTlQcjVX1zw1DNqDa6kkvAVBrP7biALnKDaDebnFtzgITLu
X1vhS5g/Il5sWTPijDtR3jPpsFHICB1Is79XKMk0vgMGimUSPH9xK+7/2gWP
Xnr2xqP6ItZg+J6rt3cBptj0lYDUOavjCFeCBhPwGHugMmp6avwYbv0m0Kbv
SwNlakVYUfOu17gVJbamVpSk/we0ZcJK0YMUEuR7vqQVZJjHlttWl96nabc2
sj5T2KItA4IFijboO7j5Wh8pBtbDKm4ntUwBrYPMnKA84kVj/2e0kUcsN8wn
+bUWyqyrYBgaQoz8E6JGnRqdOTBcK3H7xh6WBQqWK3+KDMkptNS+TY+gw402
I1xmyrZIa7CSjbju6rez4ZwB1etUehySwMgpCDS1BxtZHjZstgKz0t8ILQt/
3/SreSzUcValRWBuDv0CZUowUxVfrCjNyNVKy/0qUSEAR78lKsH5+LWWvwmf
95gc//bjoFgplPJxpNbJ5la/a+dXXHke5EP5aiUHO3ZTGw9clWAgYfkgkvCG
OrNfE1dT+KQ8M4/XjqH8qcyoYRJ7EYgqIfDx1x1M9Qccu4UnC66zYrI5wCPl
1h9HaFcjCFObCXcWgnFtOBNkWA/PR0Rp984JVNpWwHDiBsbEJYcglV2QUWDh
6Cs+CIJofcDahhPKVmHQt62fN4fSjhQXAMS9LdY+ZM7zmpybGs6fGqgPursr
t5JvszhDOPy9UPoKCAtd7ywoZM/wPkMT6DTz9sc2ksxNYrhbew3yS40jb6kR
/SGpi4/N36HUvUvMdEGx6HzLX1FDEin0iowxnSYRwWCp3nJYGRBAQl+m9O3o
bH7ss4EgkV0AhVoSA3XhTDGITJDiWcvhEZyVLe9GN+RoVdY9JREdWU+o+Mtq
flzkWQ4QfvOL46aka9rp8FhBASeeTQVsH4hc5s+vlikrwspee6yqfkKLutPR
Hca/LQzBU55083tjThlp2phMBs0jId4KNWhkhuWExsyDUFFjjp0gUlJOrW5J
RFpdWk0QGvPhRSkk9Dnbi+Zd+RZjpNzbuEkUHonYswrBt0CZhFl4uh0UUYXh
3SV8jskizaXplKuj79GLWIzfCT3iHxnP1NDiIlKE9hCvwrSNxvgM3RlTq0RU
Y1+RuIjM18hGK3RJZacBpao0v0ZN5x9OG5/hKUzZA/r/wjLJiOKb98OnjUqM
u0vT7AIYwqhnFpk88lTZIDW96Z0nftQFp5zZFueU+bT4dge+MNoQGX8XQkmq
HMHqpJ57/OVz5hMr/FWdnMb7TAIq7QG67kEZ+Pvv4oLpZjRmNY7JQSCiPBsA
3B8yD/LTy9vQdP+ro3Bh6Fg4Cd5UmTi+T1Jw6iaCxDSKKVHczLYXuUPEioMA
+Ui/OAZl4i0tT6nlrv6+N5v5yk0/6z6Tht4RRbIVUzpv/Mtcwk4zRpL68Cxm
GG33NP9nbyA1veylWxsEZaoB+GuvUEwanX1XUBZIZmGxhJ5XQntxyImBhLbb
HM0sneRNPEtK9NLM2z/UHpIyVrjvQUeWbeltLxyuQV9cTbsKQVoAa5lDl1ls
qzGcf5JvaVDCVKYPfh/Nx1r39LyB9z55cnNQqeBQWvSOn/nihxYALI0A+kFM
KFleYgwDKQJw7CKt4GtZPO23ZCAOIJJLFZmQvZjQILGsaH+q6k89whbJJx/U
npJhaYey357PywQqiuSAyyIDWEktUva1E4uWs9uqJHFGWGpF29+KeeMuaDVW
cSeONiTsl2nbd5z9B1K4dQNqFtftmUHMPuLet3NwEBPMEYJaI2rAJ8Vqb8Ls
EXVnjMXWx6W5YK9zerA9z316cGuM4kSu85TZA049Hswl5SD5cvE0JpWIdImc
LLQIdsSXSIrHqK/jhXTpV8j7+wUv6Nn7KPk1A6+ZCCpsLkRfaGtSG2GkVlTj
f8XOltRQhIOcLdsm0mpGCY72S17MojuQeG5t7WBkx5faKBtlo0+BPJG9//bO
ooGziQZ2V9A/FD7Tg139gznNfzXrzEjn1n2r5lrNF4WAcppXZMzEEpkir24U
gwSZbesBmBP8bdKBDwjFuTOddp/+BV7dj6kBeQRDEYUzlx0EC2uqPiYpc+3Q
RYmJrsyjZp5WFqzOH+2ix/x7xez7ZX8AWqi6pKLtViaTPcD+y5KVEuRv4RjN
ULBXK22GwJcG5tpMAjSdXQasiYcWcuYNVE34Yit5cCFjp03z7M92+D/QP8sf
uxhXTqEOhlhM0GMxOvAPuSGuoPV4ItcXIuxXaCRg3e/F4CrLMQetEAij9njC
TBlSK6R3XpSewLGOoK0ZU+/8CyoYuJ3z2d79UkxiVV9CgkdsnCIDkrNMtFbY
cnbH6LztVb95ra65EOkU/kOb+dE4lO+S6d925jtHI/04lTq/0VojqDSbwLMW
vZSHqN6BUfh9NV60gT/Nyr4EO8b/CVL6TOMR4vOUZFHS/TIDlnthVuCpR8F+
X8+UYqMWGruDHexjNkkTn19Pu6JpQ8fT15ERAtuMJxxX120/1u7hGgN4MKf5
NAu36sOMEMhCt/lAzccyo8Xf8cjn9NTwK25LJhlswEv55Z41yBpEc8JJK4lh
+uZf7cBuVbNtt24gjuOtr0N4Q0+OXmqQbT5cdo3AcPqaud6JfKDjrglrLXv9
aBXErwPta+fqUoQskMQJ8N4fU/kFAzj1X3YXhuoNNBqHFI8bYPvafNj3OSV5
MOEQMw1QLjUHu0yX3ccjQARXybf6K2THM/uTMZ1Y31HzvBL4V3cJRTUEqdm0
uxGw4UDnz2HT+Q5fHM2fOsbkaiBeITNsLTlW81TS66N9I/YYfZsyMGHuf2Fg
qo+0DIEbidandz3zbxkaPlwiYQR8zJLnAFXS9p1Y7VS1p2JHESNsIpQahzKk
DhUAwpaOSmdAnzQKa7RDjo9/wwMFf3DcbxrNP91E66Ziv/G1+2iXsNicUSA2
0rRVzZzNpAcoREI/hqs86ahhn+CK1VohJB0dlo7gb5k2w62EGLbQFXT+PJIF
YD5kUrNZIIKlTjYKQk1ZrPxL0AcPWn1rif8/ntJhZUmvwDqr6bIO1NSkGHWL
RX/DjaOr4gEzvlIMFjdfOYGqpHdoclRAnZUEexHldkRKOEE51PLQws/XCxsW
nfTvrDA53sg5/zzNV52bgxTfSOZ+Agis+81OJ253fr/BXvAA2aG57B5HNg7X
M23f3PQtmUjrZNGIrfRCtBrY2cwUl5SKXK9Rx2XQaujgcWOuf6CxdBMJxeEY
/JmIewD3k8dw6DjzsH2YIrxclPZu9OGkYkQNBL17jiYZ4XZlJFvkumzhyxO8
Iky4VMrlZtv82erbINIERbBpMGkTZ7NjutQLoe9Uce2xj5CqqLHL/1D0FXQ0
c9jdknj65mt40BIadHAOTFCyw7RNM7nn2Y4l3mcf9ldH4jPUPXXnEIlHX8V3
bpmbJDmX4YKZl7RL2seZNggoHojpM8mdIQ7+vzbA/OPecRn7mxvRlO7hixSw
5kS2rGWpUjkhnLXoHqVX0zo623p3veTj/nzf452sgSUcNbmigpZfF0kTidzZ
KZBVIYEGtRb20kOZzTPYZYZocrGFM+RkOFrtPwB4aUjvMBkJuhPjBcMRNrjo
FgWRBRzEtM3DMMuDG1mMZBSsd8csNMc+rv0uzBwU05k4M4QzqJj5p9jFbquG
1IRqsxIyvSzSzljxY3cEmUmetwQMZ5Nn+b138h1Q4FhWvtTuYpTAmNydd1Ib
KI8HCmi2t6f8Eq4A4rsHekyyZ7bxrLQqIGa/hDNRXf51karhESK1i6P0Yqu/
vVk8FsoQPVm5H4Jw1gWdfpMeBXLzY2FccMI/7kTphXCb8U6z41ZguyjqJXUM
SJSsfODWfHTOgb2i5BIEU2KZxCUMXh/aBEnlnsvv+ClislBgAL0VQUL063KD
/QV44d90nmHppKU8PKgUY6HprIMOPb++j+bMTy0/iDT3vwbIXRsuhq+mXhdZ
FiAv/AX+IQh3Y7x0fGoHamm/9JA/WF7nfbkwX9n3wMPdghTsMoZDXYEVeTdT
h7Y8moJQ4k7stKyzAT90duqGjylVtLhGOZ71j/d0lE4pZlVP3+N0c9GE5e4o
d4exk686eLvTjw9q+a6KI88se4Spht7t1+pbdfxDX5RezW5VdXXVrEijjQxl
OO24ZQ+ekkQeBxusvYPN7N21WaGx2NIYy9s92JB3fw+Zq3wMoGexpxSZCG5x
j5y5zlrExn0fu+eG3iXi5PSSbvX3JRqw1vQMHwtnm/7+WEv0/xHum3mKGPLc
fBPunZgGunf4b7JCEaVwFDeSsCJYwYvRs/zaEDkIp/TY2bfgozaRBDUs6KKU
WtHLNAPCvqNUXn8UxQrJbpHGeSe3U0pqiIqi0TBl/cLfGX7lNugNlSNawDED
367YS8x6lhPtcCIkMu8BMVy9OQ3NIYRbSPF7qsiVXWd05FYsdVRZYyvEZDvR
qBqbxERayRzahWPzB0pSH1zvpwqewTtZzfEjMs37FMy2jvRIf7bRYo1hoF+f
drQQXYh22xPBk3/672o/x2A8hS8kEJ3UVWnfV5eDfm40VcPk6pFHunXzP3ye
WunwJf1Bn5tmGVfrZkuZmcL/wDZQZrwMUZYqPAG69STFw7fKSoDASYR/47C4
A2M+BZtE2Udiw7Glf8BAHaN8btdvBZ54Xo6DI3dNFvMsJWCvIwrqhtk+8r3y
wGCr9jD3eo+KjDVMaOLQUWsj4ZflJDVWhCTBh9N3wRfO68fbFvEr/WZEzsbt
2oSHd0zQWKI5yqaVYlqsv2cavYmpGst18FuNYP222uVRYprv4OJUN463ZzSE
Ec7M1ri22JWjnsUpdHGdio+iRqk2479P9kzGg854iW3jibKHjsletjUecM2I
QwwfvI4urm0V32TZ1O8bFs/0MCoH18/YsSu7S71hjHWpuCgjsC28aY8fn6hz
xVP5MJw/phlJAloc7zIYT8BTbqFJkLP36kXvn5cn7BXbuqoImOfh1eq2N6T9
qks2muZoX0KybyXM8xPJQ5RZTLHpjusGUXcUl36uQZejAEcGGde7Cg9COOe8
kjCHyZQZtDfDM6UI7lsGm2yNhbkOnUkPN9vNiPJPr6rVV3aw0oMZtYQfRJ9/
SF+XZ3TPlI11MLxW3bbs80ag5WaiZHr1laa/jqhvBJJZuh+93fPNTkVaFb2P
keoUsW+ohJS8pmZ0Qk4nc2A1q95yEFGf6MLiCzfyo6CbWfsaIcdbHeFO0BEt
DwfUy5FoRFGuyupw6s7g13Pdw2OOS3ZompA+XHpAWzJwPfEdXNtV44Xl7rjq
L3mbv5b+VyWHk2mFW9uxZa+nYMUSdJv/1l+b6px1mnvQd68M7zXnYRWvdyId
gM9Etq4dVxQrReKu4n12ohZyLvf4YMg+JWpI4U0whCvhADZNo8E8YV8MFM6V
NcJye1oSFDA4lpON4BsHlbQ9QJsALzMTW/rzO1qostRJCbkX7m1gjg6eSVrE
fg/pgjCCayyE9aPp3mo7ZAixxXeBK09oJ2PyustVVXrjcUJfqH6iW5TbU7+/
KWezK1kdJIl4r9SdMmDVQoa6kcIL5HSYiPqpLnWeg56lTvgyNF9Eh3Rors7x
NIGjBSgWo5QqPfVcUSv0JhFO1Xd+R/cODAiy8+u96RVVcAUpiuz/tSbwHkuP
9ou6bICxebI4GGQjHRX2GU/33+EeOitXH4F1AVoAdbRg260HWFwEp+meJNx1
Clgl91SFQD+AOOoBs4M4VUFOQJJByvzZeK8sYvup35qIb9xqTpakTNXUGUsQ
ardJr/rszrHO7tG0S8aI2TwkDR3qG2kGlTGy61UZvdPN2EKnt6N44EIxngrM
CyXsJX8KyO8nyax/LUBjNhcJZhsbgI8Lq4sn21G2j9e2Qdgj3VzOrfKiqT8j
DELV850Dp5PI/+/wWJdxwsSvl+YOzTndnUQFAf+iYghvxPAwf3e6sfznIXUk
av0Y5ERnnRWOF71wjQITSVuaGNnd94w5w4lTNd5WjkX7CutxUqShLHxmN4Ok
jQ/xP55AicnAS5vLmEI6MY5nDhCqb88jlKx2oosGEKS5LpWW8+uHcvatNgnl
bkwty3XXZNfipWkZYfRV+3r78lltL3TtnZGEsrD2kN8gww30uCjpy0wzHVNY
6SJAS5TKG8JTFQW7yo25qgcuffMwQOErQVdbBeb032tKpALgJm7HRnvNsNo/
zOBTDPG8fEwitBhH5FiEuX0cgPV4RSIXaiqLMtuGA6XOJ48F2TmA3XyALs/E
K3LyjbEK0F3qK7V8k9VPqEf08iz6Be67UeD2P68nicvxFHB6cAK7oilFRth0
dpbHL2aqxbUAhbtKNfWIM8tCNhK4w8iVZchVXfLrMCm4SQHUd/hpZT4OKwRA
BhzSnZ4c1ZNXbrEfjRkUmb/pePYj8Rb3BjletzXqUeExU6LG1wpDHMw0Bn2M
GGHaLni07pQSUpYriZQPljeaSnMVNDctXo6/W2DABq8oQcPBOUNesiLc+2jn
XmyiX4OgyN9/ALApXhZeebWMJSECrtzsFWxjK+QKv2hgCzVY3N5lWpztVTW6
YaVYpGBqUQt5IZ1NPHBAB23OllIKnkKaW1BdtTCnEQVMrjc5LnCcepLoESSh
qVUlZum49itbkjjV26D3C/QPMPVg++tz8XrjOC6XnlKzlaoEtItbp5DHfq/W
5/o1z1RK6utJzBySPMVih3Ehb+f9vmhjnAEepdhewa7PgL99u9N+WXE4hiNc
0y12EmntWp0OgzzROmvyrRF61RHfBmQPczFmVoY1B5iuDHzzuuyv/DLoB7zO
gYZP3b1vjpCkR5uOWcLBTjxqBdimuD2glZjC3UFdxrd51q+GHtSRnkvbdAnW
LL5QVCVEPBE+XujPC+9zSlUfTZho2fyOoSCiVyEriihaOkZEDfj+K3K4nHA5
VSy5d5qGI7yTe4tzbLeleWyAEI1sIRI6y2CCThMVCR6wkhixQTkfLW8aqpOt
Zos08QBiMIsQkX9rhNr/vEVsXAY6CPYaRSlb6IW9oOi0BwTlJ2YQpupsDo/h
5pBv3yAzv1pcERt902UPUMdCvEEYUPbHTDWOQBqSYNQ4AicEH3bjkUNU5Lbk
LgYjavRvGaEgEmdMJr7RkQu7+J2PkJ8PSz31q7zqMtXWCigLoDZbdMgImO+J
HN5iYhm+wK2XSVu1WFN9+4IqqHXe3QW4BE85pIJG9794/gxInzLOHv9L62uS
lmIuOzzDxvSiUGohQq/E8f15BsRSYIkq5uqIotaSav4VE6/8+Phc/OL1yNkn
pEvlXV/TsmFfLm4bDPYQQgKiOxZSN22VjFbhI6iQGgPVCMHOznWlkdK9Oz2y
PdTZWZoFSm/Q/mIixNSAYAQaMWjaKcCPqJmHB0BYkyqmMjPN3TZgyFo7m5cl
ef+xYZ5htVOj7L0e2ZsNT8AGHweDtPR1zyplPnLD0hhvyDYdrVFl+43Zb3qf
exIY63dj2HHZkShFgYGJyhfMsCLt6xrkTQaR1uZbGZvv7GFQWB+nLqtAFXuH
Amp53etQzt6M5NBfcFi80qAFQHt4ARNMtHwUrOY5n3KgRK1fG4ICkejFVxiH
Kf5/S3O5GhNXbrz/85sEzHFTfTT20VfqeJOiktkWVTy5ZTWJxZxS8Nu8CQ0U
CF5vBSAkMGjE47rP3sFI61sLphnx5V9sGc2xuGMO2Ej/YLDUQbsa3RfpRznc
asWP4vbJNBDDQpKkMpSOsVBg8cPu+b6jMaMt/hE+XvwZw3tXgR40kqj4UOpg
0wXQoturDdHLUO1XdJoQ1zeEzyKHHCd9H+JStgDdvghb7OWd/rjePeVZYGrf
o8bp3LBHFIOFJoOzX06EakpbWPJtc39B7SQGgi9Eb1B/FKP/kZfmpzu6EgIF
ydWIqYdElxX5LPNOTPZEuFwbc0sQEePUx7AEj+KykfI2/2cWwd5Hj4Ud+2hQ
wSuLEEpchKl+TJwaXnoTJ0lS0os1n7hpbQgMUbxzs7C0rdix5/brPb/zZrYL
5xM4JwQ6jGj0jks4vv/W38Nlw0vAmGuWGj7f9/hlnLUlgjVMUkNgC/Vu/gKQ
AMOT9j0WplAT/4EoaAGolV5LxSCPHdzmF4QDCldmiqkcFBl6bMvSclwlFb7q
6sx8bGUPLYrfU313Og+Z8HgnUz1Y1hnEHtBpPTznw0ypioRGzmHw3xFNNM8w
mmKcOVWXOD9pOJngbrypTcCYLKQIn5fn2mdJ0FJ4uY4m8IKoMUtpZ9MH0bnH
V6otz6x1rj4EbGWfUcu4rgeuaDw8NjHDEb95zw62bDUJCgzUpvlj8l4lC1we
4BH+CYdbbqJJYB5/CksldwnWW/bXfzESEpxTXYj945WolgC5McBvkdUKNQD6
yTjxAp4ajHEw08JQ+QcaXV+wOdZ8avItD814lfo0BDYAZcttZmOYzZcas9MG
FPzw87lmcW4U3SL3W+He2LGVSP1cXhVyOtvK/uM8133nO94960Ijz8zme/oo
+p2SRvGwIkB3P4lazL+/qMMM/Db9NQv/yKCHsXBb873plRd+u5ivujBn39nJ
KejLP8cK4ylLsDaWp5a9u1PEFPPPldAyoLGbNwlaVD/bjk609sK23cyvCIsl
m987m6SeoHcKl2ow+hJXbtoKu55KSghwik8uUFUbWAHLdOMG8/MOJmMb8M2Q
82UUXkHa/ZdOlOm4PE1UTKBnYe7M7/pH5YH0HX+Okg/dCjzR0mqKnc5u4yTE
7njh67DEuJCCBHu5uIJ5CM/pov6aiTMPjYUuQq7Nzo6bbYNdtMC2Yq0Yj3Vu
k24OMNiel7kz/HUDSC90E0sbWC6egKepT4G3PDhNyXvDNSx1HjIb5YIyyiOq
KCjefdHXd2LVrYJBKB29aHvg6plwDJsfZ0+IdnfdaMoliiKUHO63OrkfYRFA
QyGucIo2SrrDaXVpToZprNK/qaKdufLenfYnBajxySKCaceiTsj40kGQX1BU
Au247LgN7VNd+c5cMa0uyxiJvZxhLz66RUVkcI69Afd8amE1Xwke8xlCwzJR
HnuYL+/c4iHjGLmy+ecj5izxCBpcRK/UzqSJ0i3W/p2wDCfwVhNJgCKcPQnX
f24tLxEQd4xtrzbQLaidK9tQknM9n7gNp8zuKlWLX9/IzP7aHQQYGaiJaZEX
Q8l32kNEjFxtS7Zg2Y518HImHCMMGt0PwHGHyi83+2imtADjRCurV2ym7Rhm
TxWKppN10HJIKOBXTA9VN9ZTqh0hP1mY+uDGtAXTgnblJjGxNnonYty3+ewn
4kpedKKJRCWzKUL7DMqlasxbzF7wyBvqNwZQMNoB1iocoSMJXhTAW9OOfv5u
cQjiogMBpLyQDe5JMn0At57whNwRfiLcWNoZhnDgCF8dVCd/v8+l0LmXqkjn
ruTfKq1jsqk7gokujiLHdCayAaf+YCd0UFlbequjnbnSCFZfhvmCMrtwVKM6
2khLmoth8FTp8PJGkn//iGsBuj42Zyx1AaNWNUz/uFAGaGjlswifE/qLD/by
6goKqXOSkl865/QYvpZNAHSygKGynUvETw80X+CBmL8rui3L6JjGydi/GPr9
zwFFFO4Fju84SPJDdAVmcZbVTDI1yfyBal3w5X/yf9Z/dSUedJPmGiTsAxuX
rlB2TEnXp8Bm5JTkgGZTOviFzvAD04IjN2bkek0DpeCHinD6b07fNMv43WOc
mKSng/8lsMc+mlNSknp4EtwlYbxuqJG4fpkN84fIRz1zCNqFaEsTSC/iA9OY
aIk4/xQV0yxbQJPh/Lpm6lhD52FBCuOKsCHW4TKZNXkjkcbHfUSBogpyKXe/
DT5ILHmi5wX/rTFxD72qn4CFiCPx0Um0ZW7yuMQgUdxruK7/DjVWNxfrSZfH
lcmaKEWdJz0GooUTz4Q19naa3Ha2CvLSxw1bdNTH34ogI1966QqR0cIX2HIA
xuBhYReKzXUceLN/BiNlPtBmDlDYIP3bNWNy2njTnxsx/eoFBs3Yi3CvAng3
Tx8ca3rlsVYsZ4IyxyyJBY2Mqb66yQGvmyry+ISyiswXp0TqM81Wp9VTHI/T
pme1vmZPUVluxv6KUS6a63qKE+iOpFnVar29uH0gqLAvQlmIpkc3NexjNGqj
IsElb89PU4WapF94KTt+SVXeclmFsGeAX5pQ+mZ+WJqA4aOms/W7Nrj4HYnc
Z3s1nmcgHG74slvo7YkH8p4OclG6AQ9Rr/LeFH3B2PGCCYr9mnDWONPDWEfH
9N8jX45mosAcdkYyaBlsYD3gMk7m8CBqZZBMLJW+VhCPNNuWy3NBVq6FRDkC
99N6grcl7e26ZudxnZ0ypF/bI8iTXyq7JL3XMGjKQL/K1MAI+bB5ew6PXhR7
/t5ld69FV4Repztijk3L2+aQJqXrSynIFEN6wfkexOuikLACtUDqcV4cyhpM
t57jaC9jryj7oRNy20PAAEEvvmuVy2qHERmI7gXxP6QQkKUFUjB9x63P6+P1
a55RJJD1QiF1lqpiBFZnPmrxB8N6e9ZFpunmGoxx4Cn47itME95bwxHF1mlm
X8hNYjMg7unkM6TAY/SQ8VN5rkFy8G69XzM4U4NhVtIWRWLkNPzZJDZrtsf+
9sGIpUC0IvuEuKWejyHBuYlauoc5NGmxlOjcrbwtFWW1ivMH1bsls6iooNsg
TJ3ZI3wHOV+jzHTJOVphi1L78imab3B+kJV0t+faF1+NsJVqr3WtwskOCHxA
jQAdBaJFBqTEmhKv3dtbHWQZbjlZlRSbP6zncdmf+q1FrZoPdu6j91bgNna4
PxMhPJto6nmv+MVpQgIfwt6zfaydUC76PURT8xwNUDiDrIRROOoLZOGsgDK2
ZtamD3dz5qad+gQWgbsvj+tEq7xmHqqo0rnWtmDFetc5+8RtFBITDex8JvO0
cq+PKIOaJ10QJhRxlP0rHpIGxu+nWPSPykjxpK33mCDCg+AplrixEsOFYRGY
pW9uq3byoeoxeE4LTD4l4+KR5tq93Cdp0CbBywKKiH7dD9Kuuh7pTVmiRt4x
Qg3GcmKF3wURfepLikhddsX1IYIsyLIp5z/iTb0zLURVryl1A3knoHyKevLH
z420746NjpVPdjsw9nT32oZlx1U5Qhx6IMSHOJCtW+NwIR0+yvcNYZFEKOYk
Gf6FKXqZ4xNqhubXcGorm3PSqTtvwwqBGzjQle344PEN3XtxkPsifpUYMA23
MKTSHRli8mytQm5SOl778tgn1aZXf05/ZoGQhBXVOu5IEh8G6hTp4il1L/n1
B2EEzaxB2UeKfok36cWoousqW+wtuuIo6wXmB3SBeerF2niXPYPHPAIEx2I1
xfXZ4HGTKHIskEGvMpxF9BsAGaI7PoOvIvcXehYf6GRSxe7X3Xcl0ehKlagM
s1/WgvJvIDtkkpzI5GSiDStT+T7qVNL2oSmeJ0XNPppk44vzXbQ3xUdvFst0
y3b69lQ8wRRkK+tXZHPLroGsHPRO4VKaWxvPgGW5YLuKPWtKGMY3eXyqO6SA
Vya8ajNV56fNDXWeNdpmuL1P0pWsrkQG1gXxCC6OtaBrBFtC+HdVyl7ymjvz
UvBV8NqlCcCNT3gil+b2ZZ3xVEm3kR7qDh9SaNlsDSkU9e2H3zV/RiKc6hjj
TdvsU7CJSgFGXYY3/QFokQwankpiTYpt2k4VDYOz9epk/XinqPAAUyWuV/as
mYFCi1O+Gq9W+vpX3abwjPis6v46pnjqnCrc8dTZcYU8HdltZ9wErmIfdDa6
/kGB+tjwfQ6wBI8NbO8QKd6kb4IAvcy4sBsaTAEwWoKrxk1k5qr9kmUvZWpv
K1mbyJaTlsRGNWsIySIuFQDoDD2Phhzr8yFBNJTJFznK9LgqrUpqw0+jTLRl
3H1UD25qPBUUnY4RSvlpZxf5t24ieXc/1MUlUJLhbD9JrvwrsNkG3AV/RmsU
lnlRl6y90YGa7iEJEy1iPP186YK0GYt+YYadGT2wS+5M/UvmS1eF/Nbb/AkU
s75RqGb+hTxaHIGjmEnYm/Yg+lO8SjrMXBbqhYNGv45x8vB+2MEc0u/2Bgpe
UL8pwFZJut8eM+u5bkvXnjoiK26H7ylMSvUx32OdFXwrSs0MbJjGpFlb5yz9
W5HovIVod8Xd4Wag5a7ndw0lptFYB+VYP5wYy6O9lNhZvtXbik1TyDv/xI/q
O/3I4oL7ud5p/YLuEMaTy3LY0uX5W0svkBW0L6TVdB5Byeory4CUKEYwJw4O
xrwvBDNnR2RjolO7Sz95vJBIq8Hutri4BrvJWCQ3K/GwSGWfTMaYRnaq2jF6
e7oa2grOX8flJIyrcEKIM53ToUOUfbnpggSK3TjLVqiQ6cLmRsutPuJzqr64
uJHzyt+EmC+x6F+o2nO9WL14NRkPAECJ2E5BXtlLprf0Lo9Wvn9qd9A0yAer
9qlSIeZ6VkGSAC4XOFO+qfQBYy+A1cjkZu5fHa2KtBWghVOFbeQLQpfYQ3iz
TKryNwmUYDgltMEjX7getscVK6JV//cWWpY30XRdFWVUVyArC8ZP2T3gDOkC
J76SzVMCwxAlRdpZAgDMijSHxC9ot+Qfhwwlps/G8LJbODmxtzaKpaLY2X1a
WkLMZaP1MZNI9DTKzjMrzepaJXgY3kwI8RMWFAZRb/K7W2japwgLqSnNmXVR
3fxdFXRQYGhqan39dBtowVfvTW34FcEbbrwyahHhvlk994X6/YfpTziDb5s/
mAJUaIeJBZFQqxL+X9FNuKHRJ5dwcAa9ftvNLQyvx/L91hKuqlGayXC5bUuj
myNi1VJR29PKFbAioFNHm3vkE7xOiZAUshYJRifHLj7rMhYnZ2EQ0HWylkJZ
2U/6ZdkErCzKNHhr1+ghqbqc8vv5cMvwwNmhu4sxTlQuXcCRP0WIFDq6Mls3
31ViGEirvlVl20E0C0ACft2vlWepq/ldnUtxjI8wRqhN1eZPZ4UIIZy2zBPO
BxSEth2WbFxEr2Gn9t4iiXzO+1EsjfxjSINZwqvQ3cZ7NLqv2ERMkdRFA24n
sXP3+Sie4LjqnFBEDmhZMn3AS4Gcgr0qfF9ZeDPhvQpJ5ePi+6+Hi4LHGln8
69tZ6fclXW5PN90zDReyybn3BSwamuNmGj1LMUY0uektko1CT+pAdlj0nujH
R+v/LVAT/oa5DSkTX2J2OFips4blYwf+N1q29OGcU51wuloDoNLC7Lqkv1oP
WgjWBWwF54CbNENd7fjdoyHToUe4bdnQ7DbYGRYGA/e4a+GszFSnFeYfGIlV
VpGFHmd1DSATM0Tbqcw4k8t4gmyLsNl1HDRn+ZbNIq0eWjLEDBvoiTS7qnK6
Ssb2tRJOaV9O/H27Dew7TVGx25qkaCMLAgrnx5NPNvRW5WR4SZU5EIPxcEIN
e7cVu7gVBE1OeMqc81Ec0cQd2K8LleNYvzKgwUbVIKg3e3V08hm72+QX07G5
AYdPhOc3uovkJqed99V1sUeZ+mjnQMMbunRKM/ekA5Lkm/4OqJ1MYPPgJ1EH
wVt5KMT5nabslWBK+BEOJP3YE3y9jal2/+aRreDgcbof1dhLRfCFgJR3ue9r
9AOZAevZ728gV8XRUvjSwQYuTS0UaOuwFMhSIR4IeiGcC/5dKTw5yt5GvE23
khkBReFBU+HYkY3WAPhO/xHYnYHITvR0UeHCSeOUXXaJJav7UOCsIQdKAwAA
IkhYlMDhV4Llp8huTd5/tpLoNu4Q3uo5Q5CaE/3PViRksD+azieGbKXSJqbj
G8UbMwa0VFqW1DHWU9SUEJnp/5fki4MAGcgMxtOa2y4pFr9Ty2+lm4y/ajn6
rmneqmAjMUUo9R3Q8rBoaNX49gBKh4zkMvVl5gzP3hBI++tOgvE9Of8CgHbW
pJo7VRg2ysb+S84/fj8VTAhiKhdP4g+DfGM59rfxBFwEC5Z8VTEtb12IzhT/
bFv3ShaZpJhJAiTG3hfyI9C1PIyO5YVg00gdA2irpFJWCEjyt19c1uFXT341
/NSIAGozGPw9WmY2+zJTQHaSzaGLMMju0Cy9imSYH4lkNku2qD8lMXFY9EgY
fU//bfgP4PD/XjvvylZzoNcl0JFfdaxXdF+o3RWs1faYZsI316ljKTFRWqmH
qON5YvNq9sBspN1Xrdtl8CmWCyiLCUzLeg9Er2ZMA+hGfG3Ah5aJ4PhUiySz
f1124B1l0PGRiymSCqwoDXMxNyMvhWhKYEIXIe9bq7brw0LbiTen1OV9eBlz
gmLqZ2xJVv/HqmBTtdMYMtLOMtCR2s8Ajsaxii/oPcjLkkxbAXAFZ26zBMsq
0WPVyGPuWd8QJYGcaDYjg0u41OAzLJnHn0KAbg2tWMdFnOzHJX3EOqG+BRGR
CmQ493Rk8OmaCOxIxuO5KGI1CA9tgPFpfMr+o27v9qBFxhHZbbBuBvWSpvNs
4GCDkZO5jHC0hpyTZ2VBXfK7Yg18+CT3+EF+AchegWJOtWgrrExgvbxF2qN1
E1M4kGb9frttmumd+X5cuWNn2nTpODnF442NC4KgHu+iHZedkBrS8Zwxubwh
ZcmvFwc4ZEcILDLv3HWm0GJMGtynaZIGzkV4ez6+TNkBF2pkWfb5hrzvPVmd
7m2PoKCJy2b+3xSfJbLCfixsfh61YbHKchBlf9nyqlM1H/oXhYTgvek+p6S6
izaWtC/rTmXWdhv0gZfu9Kdcy+c3xwi0qdWS8mEGXkv0FwFAZGDgvIGtWGIA
BAExoY0Kj7OgR0ghDL3E/bD20XDM+88nyZwzcnFj0DxwnQSyC1b5Zy9tjrBV
TLvGsXJv+1xXpMsKGvMD8PL9VkvqpU3lJHDLgMbarYm31Cy95LR+ipax4S/A
orJtqq+hAud82u5LSqmIpl/X2Ip1Uiet75yypjBlXtm7nj85b3b6jpSqpHtq
E0cVTSw0UbXSdFjH7KbNtXxsb5AKQuijeYrqCZV7FegHoYPucatRMo8uQP2z
odz6oF8xZRNV8ktUlomOnj4CYn+XFph5PofZ/J9BJPLzyyDujmr0yL1fBm/r
7iwrRN4ragP4oiDnGnwVMWupEKnxuwJIZylN3tCRYXwdTAjM6m70UI6pupH1
okAn5mvdPmp9DihgItLqdsA4FmqcuRWLzgTjADCH2+nTToKk++EYGnViGeX9
VjINfmGG3PZPHox7HSnnkLf7e//8DsTD/BZGCQ4DmQJ9R/YWlcHMnxXAe6LC
kmvhJji1ThG4WV2oiYBT1evPJbnhpKxJMP2BL9THIIpsFJQCHEzQK0BGirQA
3OsrV/nRb+U4W6Cwex620WX1wyIpubid8wG0qcyRaJTBYiA7f0aBmnkf3cop
LBdB6u0zv/OH9tFfZW/eZaJcCsZikFFUZmxy41sb4/2FWKeLhYIViR0Wj1QS
Pz9CRgzQXiO0jaCWmKVzwSlWHI8Xvrx0/MpHCQI01zuSKhJ1hIBsSjbSGFiC
jmczStQLxjaZUFeYVXORCB+dNhEObElwLsfkLcOKFbA1OYFpAzDKYOMm5hQX
ofh81iTxkGjQxXVMCnGV+t1sUtBN9iB1uJhhxGFD6tlVCTHVni8qZWbvAg8S
966G2MSbyPUkLk4hM9ZXjtw8oq5U0KWw+H/lW7if0uuL5xQBSPh/CZ4ZU0rd
03aqAmiY26AaU3CPIkRYn5px5dyPqIYUhx+LLEzYCxTSFBZBW8Tv2IWBcHCY
ATD6P5Z9lGF4zlAix/1s53VSDlB6CjvLE/HPLsupgRoOmGDV84nQ/PDWdAFv
lpGdoHFW1iMnZov9lp8glxxcgnhjmOvFvshqR3pXobRw0SdYsKqfPZN5DBF/
0vjGBCTDu1XD0aSG1SZK/oG1h8BeI90U3a8gqrd4GpywolhyJXeAKJ+wG81g
pz3LX5jyKdy37AUjj86w5MMoc6c8ToDYCPIoS0mHRICymljEcOlPUnGJcvvy
Ls3Pz7yHCCrmo2PPomJHK0LgRz4IirIKX9ziDfcsTqMHHKHlxFVj6LTw4FN7
V8x0zD4gJ6cDxMZELSAU7wGXBxtjvdm3zSz+z6bXCsyBDe4iUw4Ad1FIkqk4
Squr+8UTCJwRnyNQj/dLo4f1nTbziFPL5bQsxSWwOCOPLpVIqbhfq9oaMgju
TuhI7RioyXbeuM3dlEkFZCGDuxjzdmGo/by+0FU9otXoSe9GNFx2I/fNFRlo
NibONqa0G5leMUEwncvJVy/F8Tt4eMOtRVwvl9j5iW3ySYC4uAje46CvZD75
BWoNctI2qCvnoSOOtGtMyZHEWVQiJP2jo0eD8lfs+7HtW9j3ToI1hW4CLykG
//kI8Aju02gieeEiTvFI0He94Q65LcY2ckHB/3Nw93tOYJg5mYRTL8NU6tFK
4zi55/rSjxVmP2wg6eUXXD/MuH+bEI37tjILjY7vOMqJqyVWHuRcnmvq+4Ed
VvAA2uijJDx/zOVVCRRkA2ElavNZ5jcZK90RCQgJoSZdAV8UcSVznitvao9u
lZkZbL5VjIdq1mujBwDPPOw7YvHcyS5aU0hnEhvst9Zsm03hFXBkeox+3Sov
g7sBn/ymBKVa5eAoJJQYHHoPq2xYGia1Kpz+HmVOoKN6RZx9nS1UgqpJBrSI
YmZU3JPsOmKoRuF811JZNiAuETURf89vW8b1SZbvvoYrSI7YhnmNYqN8RilA
chXnP23GVkUx6FWe5fOmy485iVC67wLEKzewrAsx/ElUNTWq/NTu8GyXMgNv
9jK16WcfXVoHBF++pVqmNU8JIV/+oVHH7xPcSP7CI2b1/e2DS+lGdI7uUkS9
CgvCzKzoXqPRAeQ9oT4rmAE/ADsOL1C3yyst7ZV/iBSo+k9e+nCESy9zpGv9
47QhhmLf3EZYYIWFzNrpwxazgSGauHL7CEJ7E5P44rc+FucE8+nU2TEeuKf/
QwVtSwcdc7m79r6zwHUGUwO6oYSi9GvpIQcaww+PiNRLuuJCXnLgrv9A4brZ
sDzP2VfkHCGPsK55SR74mdBb0lDM/a1Inrlf/MKHg8XgoqKNOWVuYZZm0sSH
TOS+2WFNeCxsdRugGVR/fIwDyziFdrQXoY9GJausaDeetfc/ucLm/3fZiryx
oOuQJs1e17tzlu4xsW6BdLK4v/F9vy7IB4Fgg+6KovsJXdt19J8V2vzx11yJ
bhHYACxWAGg3RcjNrpkoqxMIEW9gBoNfeg2l5xLW4HHXIyl5Jp+ebhDXyheJ
FQ1nXKy83ocDP48twHFFYMXLXjgCW3qjr4K6QLO01ACT2mgswX2oFOLuUJml
L+g+dkGthDyHw9fSsNE7CJbEay7JMJbK4Zvg0ojm7+RvTtmp3v1DMRV4xxkG
99Hh1wT5YsCFrBg+CHY/KeGd6LGTfItGRbsV0LAZ/Eqccs/nkNZdIcL+aDv+
oHjQsHRNNrecjNh13kFSZmnL1sT2yhqicbPLApEVFi9xHrD0w4PMKR5vRpHI
7nPOPNLTQYvRZ3Ao92rarSnJwE7bBIYGdO/PU+Tp2qGHBsA/63RdjZRpwkrY
aFiFuSXveDNrg7MAa3ZC7hlekYSL1Ds+wtiBICQX5012VN6q60TKOdeYe9mI
TflhUu44riQJmejSwXElN9nVVb/EzkGE2eZQAgGZSqEv+Eg7ea1O/HFtk+Ll
3f0WSwRKz7HE9gGddym6/lS+oeVDjkbATh2KnNpOvy4JzaEBnY9MBR+7uKL4
j22f2ZGG7YGiAljHJA5Ol4CWLf2MZ1t0QYKFzABu0jgMjy2sdk+A4ZeBTjlx
l4JYF96OefkNWSlMTWd+K55CjCGq+FMjgMywE5CDkIiqjXX9wzLI2+hhTb9p
ylK7inxPik79NyJrdizCVM0Ju22lQVovts1Tjb+CEUh04Gy43SSBP0WhRiRw
nky+USSjCFnTaLznvxuZg4WKt15sVdMAq1rUfVHKvkizvADYwfNaa+vQBHID
lSXdN7IRZoOcDfQkcGYUjkGf99FIymcZSP29OkHLRTEnIRpFQqADJVPgd34k
7Kft3oLDfGEtisA8xEIqzGZYs5OWttCIDBK8aD7+GUsbZNLK6tHb4E/n7CR/
2gl9kgZiD/71l7EYa2ajmkMXrvCOhmk46JQN+PBJNUT7bMbizTpyLXQRH4Px
mgmTS+VKwbUd3dLhC1njB7fNSoAkjz2l7vdWRKEI/rpc2JtHTuQVAL7qKQlR
+6qRhSM+OJ84l492wsG7UlhtNMn/Coqrsb8k+ciO5fHYgxG5l9lAconqDRz2
xynX9n1AlgRfUsUzEAK6yUtPt28xciBdHKOA1OBLhvUx8Rttc7hPWftzlZMB
DCsQ3WKXJ24gGYGPdhMtcKeDkwxtUOuetrv7Zv/UMtPTKSxqV3XiIFY9e40x
9G026mAjy1Q6iwfTfiOUH0SWRaPdgMtayYg+vPY+UvT+kbfc1qbW7lFRhuJR
Ffmrt63ra2hQLBT/lg6lzkboYs1TH4chV3VaQpLVjGYy/KfWAYCTRg29fOhV
Fheraawr3SvWSQJXFJaiemASpvWo4fL+rBJpju9osc+3K8h8HBkiJABy4pQV
uhwhUffwPUX6QepXkf9Bi5IqNDMmVwsnMHe/hBQNvBbGR1ODuyTnv0zgCyn7
Lk9LAYjh34AnwVO3q/qToL/3w6hFTsHuYojaKEjB38DaUp4OiCGhpav1cD+G
hX9yIaxaZbra8sEjcFiEZPmuJgg9owPiM7FgHVHj7hJIIfBrSNSp0NaOqu2n
mu9ov/fPqS3O7UmY7MKIYchMl9WPE5neMuhoYCQIcKPiQGqPfAwq5sA6Tups
xkb2RGql6+scci5vpSHJW+VP/lfTJVO2nMaevfw30QaWxW6sMbGyLXfA9/e9
srolelq6AUHGFvR2eZf2meYILFBEBg6/RKJTAef3OS6VUQ7P6TqULN1tAAW9
ilSlrdQ8NjoDGgr5dhlkfnIz5nmvtkAvZ44Vb2I3nxuwk4lwm50+QynzHDNK
DonQoCVZWj6m8hTxZl3/u92m4JToPTEj0/CNvkeu3AK9s+9lteIKkIIRVs41
+7uJOHXbzht7raO4lmlAI0plFUe7VHn4/PmlDKNycOwzDtC61W3tQQkZg9Nt
xILdr0auy/3L/4jFABDTnDEEJy9O9zV8B/52Mnuj6OPeb11EdTlR21AkE7A0
Y8AOzVwG+CD2AMk5CObL6sPFcM37sqL89QYZX6On00f4vdhAR746cw1EMiIo
OHsXkDWPadFU5A8jYEu48FtN+iL9IBmgvNPKXLN7ylGBy93MzdOnrAm9SYH9
1E/bGfN+I4nW/C55F+3VcdqYiE1+XGXu3HQbUB4NKYVd/vX0Y5MYpHaMrCBq
BC4cKEA17+OKKlAAQiv9avChuFcaxvI7H6TfuKqetN8tuIWWoAP1UJIgsp9+
bXMPh70b37gff11/Um3iyWNOJ0yq8RXlp3wvcRCe9wAXGZ9mesAX5+bnq0Z6
ugUJT2A5fvb+VzXAmR+TQ1CDAR1qH2Wpj7uU6e3hCExC6yUCN2674vADI9oY
wzr2secXc2CT3oiBH1wQjGnNLm8N7xrRWkqVGfEtP3AZ7QuyuMCkI/bAjr2R
Z+hlNToMy/Ou/UMtY42pWX5iF/yfcmkETWqp2O0RzOCSjMVYGMdS3VhKyV0Y
xT+HtPgeIpExZs2A316cop+T8Z4ZtXpew3q0GBdgORBIaOOXLl5StuMMIpRL
ZbGRwzFAdgZ12kEdj/UHvN9keuEkRGzrM926cIOKf7Uec3sqT+zjz2CgT1m5
RU/SXnvLw5o8dll8aJaD8jTYpDcIt57kWScYrx/s9Nqi1b2a2Y7EMABmKKZ0
Z/khbe8L+dw+9D/HAYZsFyoxhCMoh9sq/KA05KDl9dPgt/TKfSeGCIbk1X6o
AUqCDF+nX3nOMslW6Jxwg3xFOMB4mBnVeiGfxbYGzKSoZ90181t4yHt0Z8Ox
8raTuHlDvE+buNN7RjN4/IM5Ry500ttV1bBjVa9nL3SRWJKZ1uYiyobrN0IC
htv6vAascD7mqi98kjpYD3FCmEGv3Os2qt0t/yk9ift11tNHEJvMBrDEcd8B
mxcPjy7edWK7bci2b0XbJXvj3+hxoJaA65azs+K/iM9AzVu1DLZQO4FBCyun
0SzMhzlynRq3aVyDVDOMGibAInaX1SHpISNn+7oOn9EpPgQgTmW5vr3pvSWo
B/tRN+h2Q0hrfwtqgv2OMrs0+WZkY03mptgnadUb/3Ar50qW4Lk5VIkM7nvh
wYUsnMFqZu3Q9E6gKNO4+YRA2FHUeQgoSWagPxpkmVVsgzyxmB2yzocohJsK
bl9faaQz426kpE0ENWe3n9MG3CTaYVzdBhdEaNs6peRBnvr4cOpVoeF1uoFE
Yl2hLpMqENUB2qaUbd60L4uiw/kq2rh2PSo4UJF+JWkUUJbmzvdK+PkfC+uW
CtQSW3rvQsM8S42aIPSchVEuqJKM+yl/mWxCwo6DRyn72pas06SCxWQWXflz
4rhOKzMnANw7+5RkMi++jACVaoVtfOP21Gzylcv2feJ3BTkl4iWL1773fZHN
R2mzvLcElL1zTQ4fHb2kWWhHAM17U3ITCaljG5w/LN5N1l8Bj+vvIOIkKo/J
FBk/bPVwGosTiXOybytD7YuROzSPIhLkTggMQFcOPj8wacGRYiwm/5NyVWMO
eb3QoONWiLXkeiHFGQS8U51US2NXnD6yNTR2GV9+kkoW/fY13PlpMGFEYwrZ
yze1/4J9MR3vDZ74uTQfkL3NPZixvhbEueqc3Q/XJ9EZEW8Dgk1KiJtHLYsy
oRFdOxhOBTPdPsBwXMgNBZuxB84My2w2N6Ov8Hn75WeYFASZajKCMgUCS/sG
/c+6jLXagGp+d4yi3tAZN/HVhsFuXcwjEQcftf9UZDEeJbtIkRAE+/5GG51/
lxIuZ2UiLBEXBlVEP8GynPsU2BO9fkeZpiI4Q3tiquKO6DalR2X6C/3T/b4P
4uFT3p7vtND6WvjA0zyRXRtgU+qmglt3iP+SsY7LcSOqY+rXAocwItb1CuIU
P+z8kcQS1SeMzRWgnKA1dGQFASfrNFQPeWFa1rSNunqq0Hj7h3Fy5sVFQY49
nUbQpATwH3bkeNZbTK6F15dCOt2jh/2ATqd3UJqEL3zgoJo4aRBUmVMXu67X
o2fWl/Fo09RCsaAVNURoR/46CXlrO7DjGnNqZlkx20XhmXx3rSaxlhErs8ke
qYzvnzm2pHUJj/uHk70usmSmezKBryF98wiYBMOFEluAO5+AFUIWba0TiCxE
hZHdMmUANDOTTao+aeeu3zz7/+8DSCfAexOEkC4ws7K6whq5ZKjxkEWM5TFY
rAAi/4J44Jx7bLkOvhsiKOKTNjNRUkHHS1Z4asToCHaZOvn7ochPeKlG+9c7
tbJ9WTx9EDGR/7DQ1sL5TNAK/paXXWePj4YhQaN4BA4PKNawi7mEQ+6D7XlM
BN57+EPFKtJlZASKq4uwoQ4mhqm1A4nFzmtWqZfAcntRWPRaJ+KOQ8qklZXN
k8ED31PDMbs4lQx1AEt85JFDOgll0QvtfC/lkVWJ6soP2gFxrSYT4M6vQxFE
crfrmzaCjxvYsTyMG0A/xv1PnmKTATqsZTS1aJXcrwp7Ku6+/e2+j0W9L4tg
NHry3lCsqGcgevWHuGBKCg8HdKBVOZrJ5RnawD54UaMUUB43B5ZsCSN9cPnx
xex8WBI4D9e7Io1eTWbbVY8pjBvkrQnGEeOMatEbkeAqpPI3E2tL1YGgVFGW
fCCIHD5Kt/RL6/ptiQmc4Gx6YPNbUxBsOxAj74+eZgFJ3xkIkjEcaCvwi+HK
Sy3nSmQp0C7k3eJWaJcIi3q2Y9PV9s151jLHX3QKhFioOl+j++pmd6Y4LoNk
b1IZ7BUtmUNvCUHSRx/ZFE5SiBukh00FqZpkDlHu+ifAJxIqd16ENuwUbTA+
pZL1ZknvBY4/t+Cqv0YupJqW74FOdTHMldMN2AdzMn53uoUdvOtQS+7g5OQs
bTIZAovNT0vYAUZA40isN58XG6CasiJYcnEE9Ma3jFoTlw2R+J4tG5NnIxs2
TZMOzrs0ds+EUfsFkRoyAhVZMAx0GtEdBr4W9XbwpNrgac6N1nZ6wSU17HR0
DxR7jOsrFT2uVkxh/wHOK/1REE6gvCqXmxjiXMslo4ugLPQJAlOak+2zxVQ4
WrCIV+uXZ/Vqoj9pgQTMoxjMDnGPYEytLyS+H46lK6s84wSGjBdu+5htFFrW
suiAcaElPEDI+FKbTOj1/cPmQ6XwidlmX2udqu6+4M2VPy9GpGUumeMGsG4L
1/ypUT01LPIFycIjygKzO2RuPN2I5fpdtByMmK4DT4/x4+vaMGavNX6kiXlX
IOLeAb8kstl/zmg039CRd0dM2o2Z7sCWA0eJU6R9/4ULwUzmyVT/zVeqFwAK
/HLUubOAGrVRvv/OM01hZIxo9uaukrHjizGg+x11v4BnGGnSOFzonuFE9TbJ
nVJ4E7jnpNIVnsMPIX5ok106WC5aactmj31N0+OxL+iwNXYZnH2W3glT8ias
KRi+UHxT1BNmetDbWANaLpGCChuBW/awvmE2xN28pR97CvdPv625aCNN9klC
IQvpYs820d0lT/1lBu/QZ+8AcnB7dicbyUC0vE9rOlwRu55I5QYDY8UCj1pW
7yjHkKORppAdDkHbrd8kotAuVMRQOYPpr3xqEmVJ+su6cMVeIQpHgPovaaK9
ohEclxe17PnQeT8qKsXdJ2CW1ITpg3olajEn+VeBLyMKgDqbiReoebJWFpKM
z3OX1z93X4ImTlSyIW6DtwNu8LdsELk792oWSYl0+XGltU1R1fOeXdISXy4V
SKpGM2s3W7u/HhNRRT9fzteZc69V4w/0YIzc2BKkD1RjNiRQUfD/0iDjvC1U
yVUn4daDRbANJT3KTdJsdGPGXqc0kH+r+m8leSBkKGegpptDaND6e9SZsEXJ
22JSeohNwjbWwc43ssvfoSd0gaywiby/Tjy43fPYnejBO6teIKIR4de0yNpt
KuKtubB536UANmqk1zRnYYFWPKVg+ZFsT7QiP4aOsgpuTE//uhoopcNoSsnu
VkLdS1hDhZiarTmJy/sYOK/SGbalgdIqojDZOrwmW/p0h8Nw89iuh6C5Eo3B
BntbPFhLLhrw0gCKta+NL154knh8BSjOf0AOE0Ebm7QsRiQYyIXEkmFlxV1i
1Un9DeCQgvRaCxBP1QrQxOl+zhUB1uCwSc7WqzO0eB5d0fXw1Yly26ZqqUDV
nwHMCLifnNRt1fnjtGs51muQsYABSIko+KI3cwn88SlH5TJLAjEeBDsi872p
+VLq/PdBlVIrgvzU+kieHKhkZdjydigzat4ud3MzEfnsG+nTxY9WeSdWM/Ij
djyG2nRjE20m9PN9QsT6OlaIqTpLwmc9LYa6mg+kJO3l4v2o2ILlTdbe4ZTE
AVakxJIIXFRy3JqK22T9FPHYF4OgRDAYtLYVFiTcZXycv55PNupZi3ieJz0I
KCHBwGbjmPUnyi02qnDRUbJMW9qZLImzzFiXj3AweGjgOPaFZD9K7fq/j4wi
QMI9hr/3cSLi8BKI2hdkJivkBBmMHL4LaN/lyu07GuvrtqfYDLi8DqWG/vXu
rZC6u86IAj9jk9AyssyOodlolA12Fhw1wwm5R2ozTVvAj+rm7VlLMLSKUUqi
w425j/fB2ODIkwyckFycecyqKDYOL6Knc1VKLklpMAf8pgWww6IlAzjZxWEn
Pmvu5VtCWkVI5daI6OogJLUd7OXT1s9EybPuN69QyEbp7VEGrsOlks/91ml+
sjGWxKPvoqWWB4JFmJ6oUUDPFDL6UDwuAVscR8R0Wrv2fFw3jpEeaL0j/UPg
+PFMqGzBMyz4WAmHsxszF5X+Ix3fw7wG/zxPSfVtUAneiGDTd3xMB+CMoKxi
NaZYpHf4HMjLQG+PZ6hOj9zvlTHdeEo9a2T9zF/fvXfulz2IWbmhrkJfRgRU
W5uj4LWrm60XhsKFe7ZzyGn2gNmHKjohPPoFX2FTQkp6upMuC6lPxLUoM/eE
JHYYgrL+6UAWlbmChugTcD8R2FoAZ/Xz6fOxe2tSCIfAgwNutm8qfKXeQWJ1
feMThYLnngrgKK9ld0sQLxYD5rtao2C3UkIipXlvMLjEM84nZmAMz1QtnG0i
933fVgSJyFTHAd/6iJy/+1NsiAAmqhcCA1YuncLaH+RNCTUbsNJE3pPMaJBj
94Ivp3h9/rFXvg/74nkSlweHYtWlPmiqRZ5Uethvo+9VAABsfiQXNTOUqiax
N/SUDRzruACMxnXPDSSI8ixRDmOM4Hl7XbSxnBUV6UdZ6+ICZ8ZuCsrc/YCp
aNv0w9yLXxOl82cngwXSgJZb7I1DB+DOwnhtz1/811f7DkcFggBl+JewdYPc
iKyZ6tYjxConX8AHlR/iq7+FzlEl5Devk6GW32fyLsAOFxfvKf8DytxCMfMN
LacaNDZbuCta7qsioY5X7yFOChTg7+5kiaCvOzryHdrYh1HwGYB6z+vf1BJL
FUOT5W7oLb5GwSZFUYo/5hz4XGLZWPkT597fWTazaXwOWLxM52krWWaoLAB0
+FvHSi+35JcWbs/hJjvEzW+9/4UsV7lV7EZu0pQsRkJEo2bTsWVbPrFa9CtR
0Y5av+2boB+MS8/z2+KI5Ah0qc8iqXQmilJU7Beho0vqr7Ib//Vv0PYCaaFU
eSJheMSjBPhcsC2lJfEmeeFMf55jten7v4jg23EISE+yWDheT4RqSybvAS3Q
TBXDoh36tmNLyRvDR59XJi7Pnr1pntoZ89SRB1j88rzD3G8vjmfGbssB/VQF
EwFiYqWOMZJQMmF/+nHTAdX/mLtRj7+JFlQHJzjPnydaAi6WiREz0SC25lDg
+hvijoao0hNZ1GolWmIr4r3XGimTF2sCjF9UVW8ObveSw4tmv1Gt/bJu5mkn
cSBmVXOiyrWBBr+QqmuN7tFg623hO5HTw2KJ3LF7lndHEP0nQPt4R3nh7B8j
StBaL9gjHTKi/RZEKKnOrYEqAmzjNBx5qoYiYecqyBjJtb0JtQ6ZPzBbBwLD
/ux0PRNSjh5aVS38faP+YLDeEMjCWwLNj6UGPlzL7l7rinXnITeojgj9X4+L
OBvSSIByLVgss4l5Jhk0LoBsQp9oPVv1tF2mp3o70Cbm2kUrtXeR2woKZwFe
emHizQErfsbATJwpwadWD2abDYFZtaX6IxiZ9SCZG68h8ud16ayVrar6Xa3q
AP/+kd20uVBGLoAIfl4QUNcjdhux6f/b23MsdkSTHDYkBYnpXnj/sqtD7+aE
rg8k1a7UESZ6trIIClFi5jJC5hW+++S4qfkjbrxDtJxKFePJnSMT6FcqJsnv
4D9dzGeuK4NVmyPxTN1+aBijg2eVlgdPO0dVUD1dzOBqshkuT6pz9JB8GoFJ
Cw1llLjzF0KNK/8RgA18B1CsmvZ9w7tKcFZmpoQ1T5KArJOdAFuWRHxlGb/W
zYDWb8wKy2xoAhymjfQVOU1kB1Jf032Eh/p/omoGkJS9uRabpKo+KiawPGNO
bSAJXQBkEAXVE7xEPXrwnBgcLMl1uHt2ht3XhcwdwmHZrSBAepjT+yvrMIIV
0H7Ue9ALDqFEdKbdTU4qt9l8u+k+LAtMNrBx6WrllU0lddcUvudIvjCrt7/p
cdkUBKrwiz+o4wde9YH8cmASE1BZAuuCgbxv4A3uXQO7s1a+r49BTZvG1ycv
SXeJUGvXLdLcxVSniHgNtv6Ib6Tec5cEodi5z9P/aadUbDwW2qiei081BZVw
U/uGTSYxxV6Rqvjtd5Ku74SP2NgjJuueUxW7na8kprSVKVRS9MNFDjVYBwDt
OLHCqfCB0mKwgi1lhzQ/3U1648rnSl9TLQUaU2dbUWxBnW51S4yZi9x4jdwj
OiGULkYNjW6ABCQQsNKyr6G2ncBR50Q65FLo1qzjdn587G0znQ/G5M+eNXeO
9YVj0bwIBWJM9abSvpcD4Dj0yggLbbs9/WHoeQCzwXscUTrIwUVRmiMf9mo9
p3WaUxsxA42uG638RJ3ItzeZPOLibZZoQhPwPpgx9oazGNG+Bh21LcvCT40A
LV+DrUgqmJBUB/SS8z/J6RLvpN5AR3GQXg7hfnYQiOBccDyvQ+f7zYWo2+rq
Ag1KLagKATm9HpH5Vna96bhcfgrYzIjIXzVRQIDHgUmhZ04rhhOmqo6/FQAy
Y+HqHJkZVa3FedMKdPwR4XEX6GRetGgJa5/6Yh07QGG90XrX+hCzacVi8+J7
qpBo4eMUu8mJbyBBoNty69d4LpQi0zAmcfVpghx8GBPZlV+DK7ttQHSi56od
cnhM0dEogSqt5tw78IVehlGo8j9hKALGQeo3yJ4nq1n7dS+/MUgI3VxbKKTy
Y7e3D422wXblPO9Whr5sxzuT2LVyqRy+VnKF6m1j/IF7ELWgfJG78B9aPoAy
gMkwCiRkGSxk9J0vBpmvjKvnrsGKWXgcqcWcgU/fsKhtIohD48LWxQ6Mr1zD
R9b3EnBuQPHOU1ahT/rnPF4GsxwHyzu1hFd0/R5jWHf69/yjqc0HE4l/L5eS
PpZ1znjmqxYoUtKFgUDsm/vknAJOP2+nIqEDYfYO9j0+qJQRgSgBlrcKWjJ6
5EwyD+wyjMjSWdkbujE0YIolN8NNIqXEO1LTnYc8aVgE6MqoqLprELFKwAXq
ZqDEFYpB+4vo5YvmLQ7YwlE0GI2JdgKU31g6Jsc8p41UeLD5sUWiVOIlpo8b
H7WsCoC1G0vC4lInIfTdGvE2dOoDIEyZguX5fpeEBIgmNtBxHSfuf++/H0e1
JX2ZFCBuqbG9rNFLs/QSZnffq9WlnpOEmSJoxIol3GrlUnRjXQ5csYVe/j85
nKhl/zadNmrQKtMn3BV5XShaWa9rCN37TOAmVreFIiGhxga7IOXfB0LCxCMe
XADFWjgakZsJYiwnkjo+ICrUdVjFvh6fTjQCeNZsV1WYsPuCtlWwcSLjK8ds
7RE2GN0cQ1FA4MU4yUHRadNTMidaJ/SXyVEf5WdjPqIHqH6wXqMq/HrdD/iV
IK/XZfOUjE2jh72tp9l5aflyV30clZPef02SR4PW+Xs3dMfA8jO/kUWmlGZ6
GgHONCsHFn+tH7LSBBkfxxeFQXJfgcUewjo2ZA6h9Ptygu6xgMYyaIFrvXex
PxaEvZZumy7tPAC3kQvNMiz88IcCPtb0O4i068sd7qJTH+mf1UvaLq/sg0dn
/eqL7D1IjJTCm/FXBvyOUHccxznHlGmqdrAtf712vaFA2W8hH6ifl8Ml/7sg
owU5SFKzWz77owbNDZrDTqJcH9kff6zLJWPwXl1VRY08/oCb8qZDfEHQ3G76
UgmDGEFdAXh78yEyfEVSuDoP2/sz1sTmUUfyb7dV0fLqvDFFNQj3atoEnnxq
UEuOn5CavozvlmWuhLvLhK5AVCR8Vscsf6Zi4qQpDFc7hUvdGFizOaW+2Z/M
7t4SGg0o41x3kHflbK+3kqDqQg7Um7kGWTeN3iqbDdqCRU8rKLR2GnUbx0W5
hpzUpnGy/968lVbx2Qpl08T1Gt+lub0ppJ/Rezf6I7LilK8VkPwsbv8Cg7Z2
qiv+nVxlJ7+Y0RzX+nQ+Pks2tWUWvofPchz0/d7BMcCCKFVKoaACc7EVLwQZ
QpPJwAZKoDkUSNFsa/kjFYF+2wEx2pOMd/MWRMHXNIxJ/7uG8V2qfizjj2z5
6BPwV0RwoqGUVuwYbBz+NFJWf1zLg7pHvVvCcf82x81cgkmsb0eSPGjeVzeS
yjZr6r1/WmKRlNJ9qyyp6bx0gKa3/PSEisKIyTPWiZECjQs6oGfknmoDu1y1
F6L8HoqYhtvY3DvmJl1IjZEdGwBgbGJcJrwdkw7TwTgwdLG3IyZz+4xP2r5F
AXdU501M5OuQfsXZl9ReVSpuCw0d9zeRW47l1HucFOXADywGezS6mj3sWeJ1
OzKrQMOeR2xDiDbiPsXRJaT3+YD5o/3U9m2UYI+nkNwX7ZDZ7hZkVNVTubac
x9qr+DVp3wRtwvPFPSdzZcgaWfxGKLjjjB2wjRQAXvlL9T/7LSOGk3qv/dKn
Fp2ZKHT9iaSx4jud1s1mXEAbyqQbSOI9d18Hw0I4h183i+kTBsGCW0/IfjfG
vNvUzx7B7pfjPL+0fmGFv60SwLozUOv2pRNslm4p+/quXZmw38vC8q1EMGj/
Ylo68OzpKwfMyqF1WC1n/7W8v2Yr9yw2kB3MXLlVJ4CNFm3Ccj30w5bWVohk
5AGIoFvlhSzDIr1lfwsqe6nyTsVB9CVbSly7kpTv5noCI/zVq21yvqb5L4Vm
wKWWoqN6B85Jd38qkoXGyuKIPwhyNQyieya6AYusv5OqGpOrRcL14oNIsm9v
o3ZEahLZjEMlvekNzzMOMwEdirutUtTc1a6+xYWjPQy+Gs5aLWQSIM3WfWBQ
eRYDrLMD1d77Gzld1kQXbitCOMy7NduGhKaJG5QJPurC2ngrsmmziTUujx0Y
DIGPOORtSsztSHmpCOuEs3xrZjhyXf1NTdzaLZl6YmASyAu8CREgQjlmHVR7
pe1cGBfy/Jxhk5gkdeLiNo7iSFeA8f05aNm+j8PVh4EGM3g9Weg0lSWl/6hk
e//mKyUwy8n2M4blxbWKrylfc67pykv38OcZhmO18J0XcREduY2UHKkVBFj/
QApylDGB/9XAwK6AwFiVVCi/KelPtjLXFPfwx28WoxpLY+voer4i1FHc7CDA
sf4Cbm30LP5C5jdmCjaDT93q1z7qWfluVjufw8cOBXUfU3jJKz8QNXr3mKz7
yeja2KDNk/lDxRR95/R6tQ7l7WGOY4s6XMCL2az5fHemXnkqcZs+6OZgmEfp
GE03oojChOJy2dP8oN9hjbjzdsmK8PT/HKnarGiGWdra99odk1flm+D5luI/
+r6WeLsbjbehXi7kpAJFlWGVcgoIHPUM1BFnM73fxRx6IH3SNzucCRgYRvHH
O++y817DvFrCClwEXeoT58giUyC5IMCu6IJ+TWRz9JdRgkmMVw22fzt2TUFv
mjbkkQ0OoZd3VGZ/pwIDrUgy/cBI4ozBrZyXFYYlCeysyDRrvcdS1YgNRMGW
dlkUpsihVl7HJz3ucN35I9vf0iH3NeH4p1BSaqY7cTExhD/obPqQ6ROd/gcy
hfl9YgAryIRZCKcYuCL5FPHatLW6jF6LxDSvtaUrp/Ofq3Qbkn3dgiJ4xPcc
Lk2OH3xzZ+Wx4y9T+Klw0SAT7mCoYOHq4tmpLmE5mCbiMQQICPUOtYAnE571
1w41wA5QsVEcs+nGQ/4SpZlMX06ktEn4guzwMUxQmNyYM/M2qyFLnUqO7GgJ
syy/Isa5NbaTUduPTYnawRyNCQ9I0bP3LeuEiou+7i2yvTL9ZTgbsJCsdq7y
aTgM81pvNnXD/VOgub/SAphj44Hh9jAynLWOStgo0z7Zk9mGJ2XplYS51XX0
TS6DHPGWbx0kBzwjWoVoq1DBnYnLYjvB8q28AiRL+PabS9ly1wsv1LZjm4F5
//Q0Vh2NuOYzBQeMMHjk6HyDwwJRpgtJQ8LNryPAzmN4+/YsINJiBZDZkRfH
KnvEH0V76V8K79nhy6bliFl0V8O0A+WhZ0avl90nS/eUgmKuQ2W6N5EULU/X
qtyK3AYRWnY+BOwiZZF7nQY0SjdsOXhO0NoZi2s0Exy7LbnIq8YmjSN5w9Lb
QtXeHsQdTmf9iTvR62Ajj8/N4s3u95wO9Uo0Gxj+QHDdzY7bYtht8Cz9ayVa
1DrLZGZlz3DNGFODVIT0BuZXwkpBOgjkh8/C3rmVWK8afu4wpYq1Y6JxG2KM
UmsYMuYlsFjTJvAaMXklrhIioCXaN4D18h3k0GfO33azftOWVWVC79QVsiyX
Llm4qd4Bv2Viwj9GIpoWUiVb1ET6QjvXiYucdxyvejmh7SuK6z4n6Ax+Ya34
K1QXV9a13dqLRW3H6OtnUOAjJ4q5ZNSS8bgDAnqol2+XVlTirg1r0/nOTCzd
MfkOFywDmydZmhRSqzb+xqHTU1COBrLwPKcpSxXxkNN6mnfvztuJAco3aqhK
XYfk16EX4iBGT2vSbGHcy5TEpTrPK27bOuO1Ijn65KhNoRVK28wTuH43nM9L
ymHhDwyaDJEa6HAnkLsa3wzZLHysJrDpOuMhwXkILUs8ysuaKQNOH2hVqR6V
AWhr4cFKSPpd/6jNbXrPITGygS+NB2teeQvluwTzH9KIu/nAEnpr+O8g6xED
/mYYMjYvYJ4l86muz7gGycfqPEHjxQ4ISqzSo5Q4ZfYtp3v5DMBGVhFd3ar8
hII9KTCcGCfn87Wb1GeL0NEPOxGUJk4micQy3PW+O5eUE4VXdVMBQPwjj3JO
NvYPI9WZTxUSIAiUcEzhIZY8QWd9zcOSDiaMF78ACTQV3k3WFP3E/m9v3OAJ
O633L/V6HqPdM2EBxGwSvs0mKqsSmRiXrcDWFguhpjFJ4kbjII33Me7CYqm+
poyDMJ5Vvmv8ABQ0lTPvCLb2/QzXvjVrghO9GIYcK5FWjF+KETRrEX+VxtxA
uG6aMEyxZojDj2l5R+L7rZORXWuboaH7pudTIS8hyEQme9BqGGR8P3NJnRKP
sZ9kR2ByvUkoV8k5JF076zd20ejY1TMTGerV2I3KHDtRPyN0nwPzkl9mvICX
sKPfQOCSm6JMypV11OOpjpIFPXCTDZjsmymOvoGlJoKuv07R+Heldy/ZFeoH
QOZbfoR5R3FqBuToKyOqG51PLZU+i+eBwLT8NPt6lWO2nQMo16AnbiL2FDM6
Mp6yAWseziW1Jn2y5SeK3f7AF17s9QjEOFo8eIeW82L8WeKVGSgA8TaxaB+A
g7HUYwdA+2P8ar3BWlwW8aMSMka4vDhs+hIJLiFhL7Wun/viHhRNJnXXZivH
o+xYwJPEZjaUFXqsZuLBYzaE8FkFDA9A/YzOuhX0DP446PazLq/lJRfDjBoA
5yRMCdFU6mHvakiH2lGkC/025xo3EnTXTTiHIHl/CPy7a0e1ziFNExGaEmDU
VmoHRg1I/Hd8hRbWLIb7QnoIQWICTAacT96GoXPIy21fNJa2dr9lbcUhk+4E
o3VGaU8ZhUE3FWpsQad0EWTrsalyUfXLjfCasQcX7a/bTCfQgedY+Qqu9ShP
+fNwhwMp4WbH3PkDLN5+iFVTY+XXT6lt0/tSL7skIdOqKCdwr5+RCn8nCeFm
nciqoU9OHWf6XhepqJUypFVETe1Upt7WkZ2113nCl3cDQXZM3pCfD6h1CopK
mt0CAYNQxlQ815y7YnkVxb8Xqetskas8CSjg18Ry7UcDAilZEC1qDd8HH+vU
rPErdTLjTBaae/I16EPkWe3vLIeeiPG3gFlTF2M3tw1cQvRJWsy+292so/q0
TIJe7jUenJ1L8CTCEwU92+4ToPkIvvYzwRA+03O70ef9QSM1F6bZlKw8TeWN
DVH2/jszbyZ5yO3wiJHubFSqU5VcsUVC7h7daKTx4AmWja5t5dAumx4QqNIJ
dKd7lnhvU25CMuAYPpDQeMWgR4axXx0LF4kCoQ358O3lOX8zcNFV7iZEUKE4
mgB6z1u1Df8TkbS4+f+MOesv2a9zhS0MZmfBSfTUu1SB2HfW53Wi6ArSv9cg
82Bl8QtLi834rF8wGndMrX8NMOsufHOKHDVWY6Zommz3rknwuxLklCLUlNoF
UIcEyFkmPbrGX/HEZ/zeVu1Hnj/lt9cLlmm4SVKecclXn6TSsa0Ayf0H23mq
VT5kVYqCiLQ6ojrGtZSi/d9h+w9BEke+LPdBvCI1rL8SbSJRWmAD6ekdWOJq
VnL9VFUwdVE17SXV6yx9aZa13r6cQjoDrvQJdAeK2dUsmjmuF4+akfgqkTUN
5gmkjJieWH8PhIn1qgsT60Yh5i28BSFyqzu7Oxrl0lenOCK4AuyvzAvJCeGR
biTgUbmjnEarW74eq3zhv63xhG3Wh0WJhmCX4BUPBR5RvM2aAr67ICd7Azpt
nFnruslLCBQDHWIXoKjTP2J370ClBVY4bKqKrN7UysxJVbye+DzBQAdkRFmI
uQVoDaa8CB/8p90ELEypn9ug0+ZX90NR2zwpZXDbqu3gKiDpHVpzN4h/pjWT
a4gCMwjEkL8vSQ3zRN4EXYhwE4bwsmUojUMyEC9KRURkR32l0ahAOmeiqvFt
lVjDIjKaeDF/hjJ3gcDYfKuFScLEjHEfP4FlT+ZRijFcALJPzJdKAWq1p/JR
pr/FG84yXdn0rDlyqq5i24hzOQZCdvYzE4mMS3nZ1UjeKnuqkOKRwig0QJjg
0XzyyZ4nLQ7eIj7sA6KS9dCjd3PuidGA/xUwR8WdqiDWIkZpFMW4FfhJ9y0a
GP5TjTzTyEdUfPysuN1Z1b/sn5DigZhpNnshPeqvWsE8VKtRuPt74Fd1Yxyg
7xQre6Ragq70B2R3ZPQYYKMcJpYCgTdHu8N70Cf166En2qo/qCkrZBr+3xsi
I2v1BWMr/YE/AxOzxsn9FSmmXh4+b6AKdVFcxIzovnORDfgptwAMtgyFdH7b
/it+AuzqU44GsxfCt0sTc+WZundJesAHgxuDaTidKMQ0oB8tSyUXkQxLZWfM
A1O1rDcuVbC1WhcUJcEvH7RFJggsFakiQUVd/PH5wqDiH/7QSYzPRf+0fLRG
GnyrD/EaTWVpzUUf75Z0WufjDbhlYS1eNn3nCwC/CRo6A+EyN4x4OexlkfKy
gakMTU/oTJ8seOVweRvlEHtEwH1G1Fq0ANcR794mbOWwkNIxTyO2pvAPX9fp
a8u86dNTLO+k3bsqftyLX7kT0WU8hEomK/4zJosrGSENmD9w4RDjO7hjc5d5
4E7ZnmYsJZuhxlwDpChboZoBPghi9yBPgf4ZVDz7iI7V0zkIx0cpB55+ad6O
9RT8Ug9xEmR42WLFLYv6hqpLyLs95yjb9tviUpVOxBKhUu2hRUq2otZy5aFM
ru1YA9hdBS8AWF1mHFCGBuSejLJ3ybCMXpJtDhx/dtICAUEKhHLcWBFDIYcp
obcsXCmD0QHdNMa3EP9WGMvZQhK9LY9zgODHz011lMofZZKpASlHtRWk6t8A
zZ9F3JlcK4q2u+3cNXoBhIeMNCnzsMBLzagVPJAGy7xqykvVLCn/B7qLvBMd
kN/dm5MEdk6gR23aC/oNfC6UgnklGmBmsXYDNMHAY08aqNQzzpjyVhbokB++
1vSnkd2VZpp+wlbqe09ty8OXc/5glY/zfwbjbc97SA+ZKo8CQt1sVnsxZO4U
v5+ByVSow0M5r28RFWN+5hVU8QtrOb7b+/Fv1x8/w+B7e81IMp1kdeir4U92
Zol+uYNXUOwql2ipcmuypa+Cvk+Lv/ybDlsk2nB5Vj8Vdo/kPNd+oqCskO27
FXLXSq9B+S8w8YfPQpdvxGWT8uxT4s2tSqNuH+7wBaKC0Re9wGFMzUNOe3A8
dg4IggoXQKzEkshsKk1QVl+n9nIrBimYD9b8ym8pf4pWNT7ruxI0i5+VdK0N
s2/GIyi1jki0ugDwhb8/96VEPSZ1lO955Ln3CwmVE9e2WUUtq3vHGZvbsrbl
MDcWJd9hJPN2BVEH00ZZS4LeyUNTVssMsncFdNbjhnmYKM9pzcML4x9vfid3
Sbv6lsyhI+kPfuCiyRCTryKTlqXavlKqkny9lNSOpZOty4XEbdBrYiaY11J7
6hyGiFFSvNG3Om9cn4ufXJLOGtcIXZh6jPa4338l6P6DIcsxayD/SWnQD6Y8
5/f7SHUhm3w5VM2ni4xGfhGrai/janv4wu8eJ+6GAb8PJuZDAhxTfWEwds89
OqroCY10jg4mhy1Ve33oqoYyz638LGvgyRgNTSnDI5hkbMrarPlhrPVnxfV+
VTn6kEgRPZRXAomBiP1l8EUbdBn3g+Rt6G2Ja/RfqHfEItUrgqUu8wsxhops
rXaYbwppI4PsXfTvsIJDt3IKuuJ8IKtuAiNQRSx4P9NbYE4GfQJiNcxPPrWR
hbSaccwJ7j1qwC4/Nf9dv+u1g33ixncCWvwBgkmlMfC3UGDbMHpZRUqhBBTF
4l+Jqur1Dlr8gDF9cx97oo+RT1U8Xeu5tJVdrluchViNvHH4qTakOfhtIrDr
zTBOK9NuIZIfyejEdEG3E+y2sNqBcsGHVA1GtCGUiQXjhY3CV8yt7CkgkdoX
o4QV1Dhhpzg/Pv1nGkaEBJc7m4U6JdIgISxd8RFAY/5hK2q0mHbQG8PJdBpw
3RntXuo5Ya4j/JtcyCh3ttFUOZkbBQ6QUP/ng+qxZ6xDxt0QMYqAaAR0akRW
xj0g3P8B3CdKrZ8moWWYVwVArvbEJLDHG6+NTeP5W8HT+lDNKwrELkCrLjpS
p7zZ0u8jgaLLpMAyod+CDxlf1SoPRxluqbIMWiqszkJyD6gQxWnVIXcPoQkP
UZSMsmgbn8Q+z37L3+sBi25EOENID1M1BZGJxf5Cjfwz16rEfoMae9hM/gfw
IcBqo7zY/V1WeWRNulYvdoovblYqwhinR7iiAeYSMiJfjVFoOjggPmIAsWb3
9StXPHXikwoAHMuCjwGikBZ9iFI8Wq/93hVZHesdjFXqbfSvMkN9ta+QzWY8
nhxQ/Gx0B2U7cpusIugxWBSpp3+JmZrjOFoNrexlSZ4K+rZyMYAdttPiVS48
2H8mzeLB3yq4On8oGuHyXZwU4fz1WJksf7IpMI4R0jJasXlPUfPHADbwqP4A
GwevrQ+yr3Dyt6SsuIxUNtRzqyg3oyxrQn3Vp2RRdqe3GeIW1Y6g9v95Xism
+QOOYuK8otmQtL5IKLBfg0TNIbL7VVNimAP6no7zTyra8FeoVUR16jr9dJjf
pJklRjMW0vyZu9zmIYG/TAR02PvAXVMPw2Btf76/TE+EF0QvjgZbEl9I4+sM
Uhgz4rpRwVwCp/xsBvoMklQOaoLHv2RlNkMebx87N/MBCSK15Su/cMildeYC
0ivSyLrZn5zY+tREdn/eFpBNMBd7BuBcguz8gKDlmtt3181z5XXOxNxSMGNK
wQMtK+LJ/hINZkcvEHUAavqg0Mqt/bVYlbNG/EaxBNi0K5Ua+OrMPnX8c/Po
wxGMOfcidVzLzPbQtwqnaP6sNyP0lDpte9cgeYS6VBpAmpiOv/MY8M0YXpGA
kQwlv/vWlSzSoEvq+KGHVAIKSHXsRDA4GJO3IYUZzQFxSc9u5Pmn75CAqLw2
7zT+gUF2tYEFOILMV7Z5nppRroIM3+51eYZ9W97xcpOorM5nNkATUVKRgxTx
Q56TxM1BQ/Ni7sbOKLkMhL4yXYOFlILATrXGE/bpweHaOdX432N0DjxAvyEv
K1jF0qs1Ff9/8JRVpR+6lsg9+K97iyxD4GEqaS5lIWq/8a9OKHuMEFNSAmZk
Q7JbRG5+17EzijJ0xM3aP3efbasFls0UAQ28DfetwvHgUZBjrD2H0zguqf7j
NVLgQfuD8336WS5KJrjUkRdALkC+UrfiKKXQGqVrrm75CoZ+j+P76W1/qjyT
GVzsm8B6ASAMZ2o7+jyPvOhGi+CaDuvNEAsut7m2xaS4Xlm2ZI8cqW4yrWKD
bwdk4J4vKJon+3UBlcM0CgYFkApXUKc6XLIE8Vrtx7ee3UwF8v7uIOZLrSHx
nLDcmlAqXVOVnwTYn1vNhw4QKlpWeaDuX1TK8g0+qlpenmNaoxNxA4NgiWjR
lcIzf2NsMXYnmP7h4jOOkQnhtMqH2yrgj34MX0tID6R2ET/ZxZsbOFg+XHvt
RCHxIZ4PMm2vVvIbQvyNds6j1+/1+7XIJxLLeOlkT+4bxRGpUn3a28iZx2CJ
UhFDkdwdys7EH6J0hSOSAu8Pv+l+/PzcXN2ZDvT3LF5YtvICM+U7IjVkbdkU
XKmLcsrA44OZJF/VqkpsmcX2vDr166pqg7LVZyFHr11NwPhpj8D9fJpcI4d7
DcQsAo7WUxYE0l/zpDX0Yurqv5MOswbbDxONbH43w2oM8LJ+tQ+zXn+8XC8d
x8aoTG0VunExCYnWg/cA73toMDct7j/Op7YWCBQoGfAmUZiD3J3bDMEo+S+A
z3rUCdVLbu/oQb6lY0Iu5GNezq9HCZKzcjSwQ4BtCn9ygaEqEIBFmNRZ7ld7
nJLXgLl7EQZujZ59KvGZb7pjg5S+rGS7kkpCiIkG2A8vP6LgHmRNvrd37NDu
DSAcJPTKYS08Zs4Bnkx9B/QrNKkXzAqMBsPnA2WCMV66DpIJIHQftmO+Msnf
p8vy16n7wtIfX7t3xvQIozjhZuVHt9vZMijkma4C5E7yXOgiie+vzI0ZtlN+
Fh7ujUL9R+WpO79MSXCKfe8+k0U02AHYRwG2rDrSehrPmPkpQdAs8QXn4IGe
LHI3jt9HnHamKgVccXV+QLlcMzZsIhNHNPsQ9bgsoMN6wLsruQHVZ4XRZRnP
uSb5kw+saERtlyiKQkkWn7fLOqVvSw2DhHNplUVtmxYO6bpDz17pz365NAq0
zUfDKiSLIQ7E9y1SH/EdrravfVYhyHJI1XKgnacuB6qgtx8S2mo1MAHlVv8I
kyU8jX3VU/tGveC30DMdBae9LPc1wQXz3z80mMJg/hxhhR63cMQCypx0VdMf
9dIl0MOqL5R41FvC/EQ9isbGngrTEIAyqIlL+MR8ymNuA+LViesevg2zDEha
/mUebKsfnJdunu77PQdMt/XnhWXcuz4V+K/4ToxQ4EoFQ5dGE1nezxQMgy4p
DywH4Jwdi8WkCkOIsm5zyqaqVVU3ZBdDrKcOT6boOXUC4MGYyMXnsPX2QYVL
zartfOm9IO5iL/gaalioYDt973Trj3gwX3xfhsaV8HC8gck3t8E93zYdgKUV
XUO0+BSyJUp2XURz0OtwF9WHjIvLT1WpqgkluehTLpGYuoP+DSpQZVx6ToWp
wIf5q7qSFpajKquGCkb3saBYCG/rxmEeMD5IV5hWcax+zLxzBvfRE35SEwTh
JZs1P6I4ZKHC5IUBgo3rrv+Biua7v1/6Yg+Q/TIwn7LYLwGqGJS3lZDgBvDE
GC3M+4iJpX5Uo/jJ7RrH3bqbvyO7pamVBgBPeuXki8nX9nNfWMiy8Y/X3yFw
Qe7RHONLmzBpInBHdOD2h1lBL9i/24rclW7c4PVK9Z5QhErmUCdMl/WXcISa
VATLII+NCvtnIoldALVDW+o8ti2NH4NhDfDtXEzTWm/7lEVghf3q8Va6JvKp
xSgZR6jxnBwBHrmqnATR3FgfMq+F8gO/X3Zgchz/ykTLEoAAVUWW8l29E7CJ
Ft5OjYXU47QXydp5F3+8FvqZUwG/WJw0Kw+AsJilFbWrA6Ob0VTR28ziNeDx
0usrzzZ4pl9zOB/DMbVduVi64fBLo8J9IaXSdOv98xUiGNYC/3cv+AetJX5G
CRujMNu8bszfzy5eV9E2U5fDyNAJofFwQ7SNmmsa+ATDA1qre/mqkFcvnlyi
qIbL4hN+xoVcc51fNWiLdhiGKsgdn//bv+NtpQNvpfgkdvCEhBmGOnCJvBB7
G3Nfa1nkCoebaua+fxMMOELL3WqN4jdj8YfeCKbGLzbYOVTrWMJ7EHdzDA++
B+6jnTcyo5IWmLw0SzZrVIGORf4bsFGGFvCwijE2xtoZp1jlwmO+yFrbS2A1
eYK6RJraM9+ZUxMTaEO0O3wJxk7b1J3EXarzV7t4xAFQ3ZNldgNbTSatzrX9
ZS6RJ6C7loIVnoEw2INnTfzbmZhM4B4ppLwQkjbG8oKq39sGlR/ISfps52oJ
3sL6SYEDUO8pvVz2db57eUyyuW7gMNuoSSGeD50DXQ9DCUVjvl3KS7EsNBNS
eV2a7JMJLlqT7PO2ScQF3KZ1TW7PUZ2emth0mplmusoJKmgHI0BwrKpm8jvn
WyW7euh0ON9E6AxGpTbpoqXRKwhM1iDYWhD8f+pC4lvMX7VW79NM+jiGHIFD
040Z9/XsiNOOqBIoXO3jO+9xNRKpccH5/k24anqssQUt81USLUgx9aoJy27I
VKYYcJmEfyvdG6Otn5hVB5fpuUvaYAwvK94yXSq2cuTK4IHmxqpkE7sKScMK
67ng0GUbtyh7RlX/z6q/f8yOVRGwabm+sj4ygVJTniW3mSgQN9T0LvE/v25G
3q037cr7a1Pn9Fqs6btFl/sjcXMoQOmtn4e+6CxUcGihpxidRvoyvWbMPa4s
OrJMLD4OY08VP4fPlFSovNLNBhe2mL3sTeAfUPRlU/AyktzN4GpdE8lzoHx8
/8MTPs6dJbD1RnKJIlNE5xgpB7g9teV9SVVqyvvKoa//b+FmeY7grCEHxa1x
irWqF9TGbGnW71YkoLUnbZcPzZV5Qmr2JaS1CNX2SPTABetlU9VRzXlEoCQT
0SmnG+dI3zmXsKFWtaimiQkMYYFMLBpz+WC76jat7FRwT92sDAc2oFjxSQQw
gfvPo/pgT1uU866TbUsMlC33bHSq+YPWkQ4YXGEnfFYCbf9fUe9HqDLk4XQA
IFVKzhNFaFGJTMLTHFL/x6nsclj+NKd+80fbu0C7csutYsChiq3S/YjgC5wS
C80qAptyd3tCi8T51rdp6qzVSqY6dMEaXqLcox6+JF8736avajqLbidy1p8U
Z5mW/trH8PehScpnTCQVB/KxxevYbvoT7NWncwDikEdtpIzUla3myeXLm/wb
dYqdL0saddQz7EQ8r8peuuOBKItfjKWQb9oUxoJrpztIYxzWq8v2antQb9ZO
pcY6Qk4UtMITW7asajLPj3pI3k0bARja8lqVLC2eiIdIPPqL+Y4NQhFSYySQ
wN/R90qJ9JwfEOujWtRt7e3Rf8V1aVNkqcfzDVY/JdFKtnAdFFgTzjo3c3Y8
wADKSALy9kh0jWTrl98CAzCrvarcRjWeJe1MX0WTaEkmm6APzkG6EZUgrVOm
4ExgOpgGJE3E6pBPINNUgiQc0YkfsXvXCjdG1j+bhvFOzoFb2hbUIvkj5v1m
9caUbrcAoQmhUp5Cik7ofarXn/IBKmzCtbugGS7THNMagJOebPfmXTiyn5t6
B6NXj3xygRCH/uGzq4yt5NxRKtWKmHxrOQ41yNR0qJMouMHvRTuQ+C2MD2b7
bBAftsE+gDJC8xVnK7UxyRF2rqvG2cLv13z1xGMmi8Uxstb7Jp2vWuvUDo7U
SciSqNlSbNhv/Bgi1aPB3/64HbheAlDayXBqxYpIWV8EdTlOLCo5Nmaf67xG
/QeQJZcfjORsFWYf2OplU8APLgxNNmuonPl0MHXM9i2J6RaK68ez/YtWUO6Y
RKPqb8ICBEb6GYqBn9KkA3LNHwf7MX6HPDx7cRqBNtKjt/XOzYIxZFtq7UtI
utEAgczEQuhWbKtItdQW78dUj7oQMtpLMZuLykRz5mumQ0VwUCIoQab4gAQ6
m0Nok5XhR86k8ePDaBqUJdfVHq1K9c63GYnFlj6Ngg2QgxH8kBRVrG70r5Iy
kKGKLgc9DLUh69AaHfzQjDTuqTmoLXkpQ0bI0Fpqn6tvHnVydyVgmacleYQB
EekTKqpDGtlRTS0pXHVuGTsiXJUs1OJbGUnZFsonntwcnROZW6By9lKqfP55
J8KUq1DVNrVzk0qYamm7AKmBbo12WgrEcpcCwk/plN+XPmNkd3pPglJS8kDs
0YNppXAuFMfmrgNMuyP5yWiKpeoJLuZUd+x3WIAsLgBm1+/qVw3VeBt3iZ89
EH6cZDLKY8T/irU3nZL72/GLjdjr9B3OozwYEUPBPbbKTr8Wq00QyTxrKVWV
21HjRm2MKgs1TCOAOs50z9RzIDtVAGzQlnLqfs5JmYEDh733PdhQGsW24NkB
YVtU9MvMGitz8znQUIEQWHDEeSyGELZIeIr4HhcWVcwkcQQjr9jbAozqmic2
15ewZYtgwvZEXxBYt9V5pD/Klr0Wo9ZOTGsZ/uaM+eJ/g/i9t9pd+s8qVzai
mEPP5rlxbvZ/lK5ekrN70W4z5OFk7qYXk40m5VQX7E18kALFPKOTrhX/C4ve
84Amq58QH39CMPcw2SCOhQ1O3pvTctgdid3VKFKP+w6WelQs6kFj+V+gPlnO
g5EYXGmE5+JxQ8fewlkVp7NTXq2ZtVTtZmqpLPAfb+aiB/4FNlLLb3yurUx6
lg02DERl4dq23KolWy9to4MxHda08j8EcN5R9CFD38fYRCQljhsHXfiXkjTk
E7o3VyMa94OqWnncTs/gkB9iAhaxtqZhoqSFAHNtRF7+x/tT4nz9R0jvTBiJ
iR/s8PN+sYR4bCorxm0mk7pFfZK+tb/A9NFz6an9/mnh9kaUYg2D8paWWDvR
eol/vYkJDYmA+0Aw3AtNaSk6tX859vm/NbPOOB4rBwthjQH7lQ+NPZZB6Rpz
/+o7cl3bnRHkQ9MWvzKoIGYALXVsdv0IakpZhfW+gCNDNdAMKuseUazGyyc8
IwvmD4li4ibK7OQv5YRLiTRdUlMkPN53FgMz3lYVOoaVC/IIduogYy3qf/iu
P2OM1IpSd9JuFjz0TDxIvbzf8Xh3vaqK/tRUWrY62KX+oxNTs2f5RLxcI/Mt
9jDgnM7KYRNzarTC4tsQrME5FqB1MFrmYPlVl+sv2iqom7zXSQvcKAs2XUG9
jzcCcsfdC/jaoJ21nj6di/0hzsi4TXI8xemvmxpjYg71hK31bxH4wiXYPJZa
HOKMxZkCwdxWdt8fzRr+lGpME/PUEEONl/DPlZfDrTBZx9990AjJXQL4n1d8
7paBB9lu3a1xw+m8mtvJxUm/xIplM2MEsT+9/XpDYF+U3Od4CDudP9UrbhLL
ROlgo06wiqXx5LyE8MpBnf+kTQdUCyUb7kkZc9U2TRqsv2kNeFDehZYn2awI
Kr1yoeIbW/jjqrlYZuykV8iSq6BeBMjvGJsBWJhAsjKMotea2XUt1mcqcSXy
XkslSvByY2hQLB1Gkrb9zK6XoYMo5yrtEmpeX8S09JtRAUEp16/tGP4f6IOf
UVhkr2eXcGsw8T7HqCEHUwu9x4ltumPevTbC/6bHYwcDqI1Bhn6JRj5/dkUI
VVOO/cv2PBiO97y48kaqDDdyetQ0f76hMAO/ni0Vb+qJpIPXYK5pdi4qWEhE
53i9Pr/8C+1ZlUvS0KpPuTVz/9WMrnFOnLQ02WDCGO3oYiFjN+e1pAzqdTzc
2JXSHEBj29M1n8zLqJ6HOcmxBX/nYcxAUWHwkACBG/YXceCKbpCl1r8dDPDB
E1l5ZPaktA21xfPC7HnQ57q3Wa2U0+kt/9/QRJieagw4WXdjW99wxWb0C3fi
THvlimsWoekLb4wOLrmTKl0JgvwscikEnhl4r9EQ671VH1Uo0aFdhZS80U7p
NuzXokqZN47b5dubFqavTRO+vXoKS5Hag1Y/C8nqr1UYB/nsi0Dz+fwMPsqZ
Zzbt+S9EzbPGSzXuCJ6E0Y9djcweEXKfdu3PTk4A6akoR7qmED7/hEKdwk9g
18Tw07pfeovLtmjxxo0QJOPesJ6ScrOoQgCa0cRVHbg0wJv0eLMKakPWnBiq
WdEIhxatesZ8obJfRkMtD/escGvW+42veeg34/3x+kcGuydX9zBej7Er+rMh
f1kw34S2CuIAPdHSK6Sm5wSzZEKaKyxgtS1LZW/JHjgE2izNU8UIeXjW7m10
XyAhCEc/dKC7x4vjEoLBaKhe2+bSkIKvmBLqYjRvIVLLNV9/enG2eAcnipqX
GHX+Jyxkd7wyUkp8BswhUDcUrhkzbdUqrBv7uj0ecQwHshDfvlJZY4N5L3P5
eKQmLHX46ptcpYlj4HgiIbgpy1IbLQ2Rd9wOV+BqZ1HZuBhNQdoXp3h40pmu
WirNh/+5afb6LZTIGSDvrESjXu8cFHj4L61sBHyTPM8BeUnOwVzrmxxfHkP7
/DymWT/m7STr/m2boKf4DhJE0oBByQy6CKKtuQq3FZp2vxTqoltASO4RM7/q
OhrqX9tiOL4bm9BhXpH0bKaF/J8zFKQWDk/QKlY2P3rNUp9AQI2m8TUG3q1p
5wcbv0vHltTIfNXpq9cjj6tVRFnHHWPRlVRhRGL7Vx44UfkooJkTBvCjnjgX
KZSbmZiPHKxp18jcJ+1U1Ue9RGrdb6U/c/P7SA9Rm1G5jswSqyANOIdJnFt1
7skw9qaKBZnr/dyv30ki3QRgDLbrCAN5s9PjQAyO46upbTu9upcqbU+E03bc
n9I/v/pDvP9HS2c9PICoIl59VbtYOMgI1ZPT5rkgdmhHbbRXHhXIwZOXE2Cn
BhQXj1gqesCONza7gCEtpYcM8+1RCsx2wd84DOO1pmgjA2RRtX+gze0Wlr3b
dvSNLJcgBf58S8lrWhFpEav1hVzwDz4GRydQaMmP1gZ+x7th1XYR4itPw2io
HIw+SwM2swwqX/qdIkOKkRaf2ZT63SZH4L1fcH3vV93ud1g2uXFm4jqRQ0Fb
V/Mtv6s8cvslFgEpxXCDdDspf4ENKej1Rgl4tWVHoI50Hq0EUAtvsXPIA0++
a5y6MT2ro4P4NY9QrhTysJd/jlxXP4yTHaHsJZz2uLd119l1d+EDUbgNJxeW
/8ttlOf603vx7S6UI9boKYNUcBjEOGiXAFJlmTCZT1cuCtwsYUtAE0dEnWzy
aatsDBFb+CCLdn9TqqKn0ztCxhaoR63aeHza63qnX+TgJE7VDSb4D1PBTgQL
9gWkvb9HQ8hT+3V/qQGqudl1aqez3lpLIynQaYUopw4YAE55UQsjkU1kG7Qs
DQb3UETNB9zYW/H3IgJSisyukwgUSwZNi1MUjYZZ0WgTmivoSo6gIant/1YM
yhTHp1Cef9ALZlSmdM13uBfMBCeZ+hlbCOIr1KjcT/O3Oao/UtN586bz+ujJ
GFqxySlW1AaypsONh86Xl1/Tz8ht7xtSoiZm0ZEkvq6r9LlYjimTHrrDPWv7
XZEp9YQJdq6GD3W8XN1Kdwbvv66VQi7TfMgNBCIm2P9E1hOlf2qx80hmvoIH
3CAMJxtB2lOLVaUgZYTEwgfXcBUSzmx/R9bhfErIEHa+PaQhS2QeP8vHTe1i
qmsB7qdSlAKyUxOEmXvVbJCxmNUQV8XuMJbSyCbg757GhqgMNkNQfkqCAj33
HV48nlHwhSD+GacFIzLy9OOhB3lbdr3GHMpYVLF7UjdOy5KVBKjqaHi/xmlv
468L5buTfGanYeleXu12wQxN4rGjZAX5ZbaB0JXiVQ/tUwT96jWrd72MxVZ3
glMdwgVRvAb+chHAllMjLaz5UaQ4w//dWd3CWGuAoJGpxvnpy9Rua3Y5rE9g
Rg2iTXW/PpTh8AUyVOCKPcWtwQzXr8w/bw4LfUAA7v637lTfbKkwzHHMBMUc
WZCRF1kPi6GBh9vWQg3tz/ittF4H2ARVsFCZ8ECHaR8WmA2WaJdXi2q0FHDg
SbNrEhFc1Up3v+5VvyJjhtN+KqwLyX4er8YvDgjaZeiKGOCTbG3+WiyMBtGk
2dkxu/cQw5m1n0QBivpwfb/HmTkdH6L8RjR6JLbx1SIhryG4axSln+r7OGJM
wgfGa3NjnH2l6fZqNYKC/s++r1KkpvCB4KYNlFpffepzctnLOStTP16Hf9hU
d1dw9//mi5jUz5V6rK0G9aj9WEaFMcBsAolqQsPJ+hGqnfwYYS06FVXS3fjr
6HNZT6D/8rKXTmyMolUNiwVmwNVqFsCTL7lq3HZ3PisoyHREnQFqaFkvfpGS
+xv91bXIsiASiO+VjzY2hVbPDCdyB7G0vMuNfGmd9a/oEQNjyOKlckRZOAsS
zYRzXNnjprh1lRQ6IlGa9sPPD0KNQJ6vkCE5KzvLJ1xnUSCbGv7DtkR4u+l2
a4J8FXmsdv6SL4FMv+rdHBbQVHvMy6O7oWMtr8nIV/DXdaeqF98GcXWK8Bt4
9Qtx3hmZLAV0gvsZoEhh1Axhcqlw19/0FSLGFGMOqj5DoT4qTL8pfrXxoNA+
BIzJHmOIBCIiVKS/OX6HiHvBuweof+Y+TkPEPkhJ/qjyIypfcvFsQhFLhQk+
aCt8HiqEUmPrGeOB8yhO5b62VGdefYK/9HOY21n5qvMHzOOxNVvnQq0FMH9P
JqFOAUqO0TgwlOt7Nn7St9y9SpHXIrfzT8JwwtPPKu9OZnXoPYBF5RgFbRcC
wqCGgCVY5dfRAPhEj4seoQkU7MZmekfNKbj6XK9aky1en/VgGUUszW8jzoKi
yuOMfLQvH+GCwNidEcjyopvgf4j8Rh8pkfh5f2P8eqlAQwzGJEMtZ8dF1BUb
13uMk3Z4lrAfdN5QGWGcrABK9TqKDVbTHyhuGoyzdzh7V067o62a9XhhYZ0d
1ncNM54zhF4AHl+1Juo7gjygwcLqUmGz2ACOhKZ8Iz0ddz/gr8ehD5dpQSbF
Ksqt7dhI8GvoyiCIxNvzDcOMJdCJ7+Lv4iDvYCNCO1RkRCAfPO8a+3LRXbQM
QfOZnTPKpjrAaj/ibmRsU8Kg0TYF1YObT03WJvEDC0cwXdX4mPFVGyXEh+II
WF1qV4ypyM0R+7kELnA44RHBbY2jg7uU24mjxYZ4hnal3u6kS7Tw2oIW5QIR
N6tmpGaURajUyAykR17H4JSu2oSLB432lEYC0eZzY3NFPaOsVjwkqCM3J1kJ
NrsCXMR7k9jfhvZKyfxaDI85wvE0xwjZT3HhgwcaMkeDM1w0s1e4nDuIt9ro
nKs/mTZ5QVmyzsyVbeb5kvfieI2rOyXuz4Gf6/yHsx7bDQD9Jox9hDxxNPrR
9+S6D1LmAsaev59DrWh9DySkovIOl5h2d2N3aAA6PyCl+1XSlzKcK0+sGnVz
ReIuibRKeL+ZLZ5pMqFMZdnD1zJ8eiIBPqfzskmG+66PsMmPHyU+Kjf07dj5
y6ASu0sosMHMbkfZuDer2/mp1grJPJrf9sOOpPOulNpdyl097uq/xbwp17rX
OcHpLoo6ES0DTDQGBeOfMFHtLv+1tUcFnIAgvyFbTAz+SJ4CSQX9RwexCulg
SWRnMZGCB7EQgmnyDReB77stncJXbG0aX5oHCAkl4a4J5yXyIEyN34t+OvtE
TQgsHTQmQwnnYGpwc5Z82aVy0jd2wyOvS+o8CN/n7jlycY0vzFEuW3LB/nOx
N8+xjMf/iqdabFPkVmKVKk3Ajbiv+Q0pYeeeVpaf7qFzo1KmipI6prbIQDrs
tEoC2J97TNCwDhl4yuYosib6V1cGC5GWVU+wNHM7rG3KyLSFKgBjx8F8QmUf
vLCDKEXlBRyGlYvHaxAUbzj081/PknNdvpW4xa0rvCK6LVhLNzy6ElclSMIV
8XoR2VrQQYFWLuc10b4CG1dtkQ9lCKL3LO6kKV7IkFejqRb+ALFfB0jEeyE4
NxT2jHJOKwRpHBKWXRudfiiFtJmrQY/0ZlB300D8IJXS3lXFsU0sa9hMiTFb
1MW1vL3Rm5Tuk9LXgCjJ/NegGlXPbrHl3jlV0uPlVHgBa7fSJ6PPccarUHkg
PW/jeg16SAPeT/zM40BoiGP4C41QvYegAPZ1Esvc776sP5hL88AauxxlQWGW
MpgJH8UI8X50IPi7vTxN+tpYjdU41vhzKCdXO9xK7AzdTLf4qX5BiAqIHGcF
YTXrtjoHI+O1lN+1F/feCCDHLdAplVjwvhmAZEmMri/ng6qM4DzdHXSx9ZYL
CsbzKY4e9pFuN+YhR8GvRJD4hqbVXTwWpbNVUqIDUn3TGvcSv8LkYGsPiCk9
yHzF6tB9gsxuu69ZPeMN8WTzuTBxO1wwekGw9Ez82cimS0CCnISynknR3MLm
l9VkhOwpYf8WigltWdqVMa6oEty7z4C94x00jztgeRE9XpBdjDpitf9JQW7y
3ErptwhZML4ZHPO3HWRqDs5IfL7GUFTc148PUZ8cYkTzNBMUPT6yFIWnFQ1/
yWXMeZjwdZ6tpxpBNNyaiYHP9avaBPeznpfkFNDIKt5FDFctk7mfbroA1es2
/zNOu5bRyqpAKSGN7j8pIFRBgOqmCvdN2Q/af2qxnt1mwPIa01hzlSOT6nVc
/8ZELxsc3fWg/XIsUhEZ5zpdWQMeQHdtoYBAyiFs0zNbNL3hCDd29Z5vhion
TJTRU9VBIZZcgEmi4WosIQjdOeThxgTUSA9dt75pEK3N9cDM7jmVKMfyDKSb
LYbh7sRfAaGVtb7uXg5J93b9BxHr8fwTjZfSEejNVVpOpcWyQA0tHdvs1acM
iHUFOZSh+uRJOghq2yry6fxsotK8MTw1b4fKgSLux93F5nFphJWkefN8fTEW
ZvaDkBp/2kuJvKtO8KI73NTrSghxTaZ2Atfj8E69fcbFKuoZyAiS5zRVw1t9
MzA4nG5S4QD2dsdK6e4uQ9BAKA95ptC400Ma0P1rqzMmyAHBUrMJ1GLCPx7W
rrPHQDK4Nlx7/+/Pk7bJ/eGxnUtwkghSUQJEsTj7ErBZvdjc93FrOdYsT0zw
tiuGsT/gRjU/rf943WYwjUecq+Uf6Vg4avwUmYWd2lN4vQp5PbNiCa/m/VDq
LtzYYh++YvD8j0XnAJVZ9X8HIfdj/kVjUTLF+/Nq1wmgved98jnRokN+GvuZ
5wpUkJzr+JAYuUFrEm9u33faM6ozoLysXMuD11+PluxGZnkFMDKirB/m5HX6
X0Kp6R2aKjOT45YJL6nOppWdLCAEp6scMCAv35sZDqIsC9MrLBTacQxDJJNA
cylBf+gI+aT/SYW+eqPQTpcFHJ/FibmkEf44hT3jxJ2nG5jMBYKGdLZNtCCA
SE9JrNm/dfaHLOKrUoBivTZ/wRga4NmstFcGx52N24yDSYFpSZAOAVI4JwUs
QdrGjFK5l2kTi2C+Bj38c2h+wcBpoANuLvs0gwBNHcpNq2ZA8Znvc3ibwE7B
KN5KlSdRDXek0fxa1/Z/WVLsRTHtp9A8l3aSM9WBbZNS7D0uS14JqbQQAF+2
H3derMdHlSnpLzI5U6c/NOvcx2SvF/dFQbUA6as4AiXUb915eKNqA7h1BR1j
PnDYvj6CYtj94YwFeLbGWF0+SHs7xhM0evUqQJ1IfnjTxKlIbwzmHA5LJnGU
8SNxkx2yIwcoxVl+K0iIJ3DZiNr8somhVTsNWN45DHzi07gtxD+JAnt+/Z/j
SxoTdGIwDbrXyqQuDlUCr6YJjYvF4sxwhrSWlCLF9Hr3zveTTQ/49cqAM52a
QGZFgb9Uuu6GKZHfP4HTX/Bu8px2V4cQ2jq64+f8kikALHnvqUOedQzBiT0s
K65JP4lWGxFoh7MaKF6HXXBJ9RDJQ9hPTaUKviQt7AYEhGjM2B0E5w5GddMS
0B7KuobvTNsBFCXN0/CfOCjS/8NTAgvSXl5zc/OgA+AFhEXUcGnRLpmVcJUM
QFa0FBVTBwu3XvdC/OK6i5w7fWN/zpBCOFO9wdhMXadSvViN1nfDhue+1l79
2wvn3i+RWWRMVcR4qFTkSFAkJ2s+EEc0R8VtquAJoYaLXev38EK/bR1QzRqy
wTSiNydl+uQRShazHOHKpydUsuAx2cQYkCDGsoeS+bCj+0ighYtmVv/fYSvv
jvVXmLoANui9nVhcoG2thpt6fSR/7vu1+WRBAOty1eP2Zxm8b68K0BWD8xYZ
iTOw2iRUPLOZ3W+qqTY1ae251IziysZqwBlan482x98WxNuvJKdD60wFlGFZ
52B5DHff96t577UQl1BDj45ZwH+0m6JBnMt+vUISGdJuCW9cY4i7yBYm1lfi
K36X9bgIVjw2nRJTrASLi/uI/iJgsHl0Cd/wWPFLbIpmE/tcAe/luGriBBFE
iTKVGCO+VzIOYAaCZSJUq2I977qh3s0Td3kucA2zIY88waV1jVuRy0HpPJ1j
Yiai5mcx48KtPTkIXLZ5WEtr0RCj3MvB+1WZ9QBHyh2gMwgrzRU+s46oymga
DOXfqPFpgC7fFtL+KPsWLcXYKvB9TPw4tiiMjmQLqAeLkwm4Pcmy/KLpDGoJ
UchINPY/p985sxQC6Mf5MYq5oXaCVO25+6Ve8bbURFCtHw+d84bhxLU1revu
SBytauVb9KceaqCK5adRekpgubDyx+SCTnLudjtwyRIgcWqrAgLSksCNPEEC
8bAkE/hWA5/gQuY1ThVyqDCO0FY/4dkJQdXB9uHfmk4RmU2cG+Fib8ooGhOI
7VsHHvtR9kMvZDXt5zftGNlG5hTKFS5gbWPDWFXpImGaJ8QpViCqlQp9uHiC
DkvFD/6SDhLMRc+ySidyNb2hdORcJYVic8v1QCOQWOdO6u6oQvLw0bfOTU+S
dieUHptf3tPz2XttHuqYovB06m0tYqDV+Cj0Dza5H6+rYvBHUeOSnBuRwgff
lz/Lt8ewdXMdrnmSZ9zVP32xO1Hv7u0vt01jwrh1WLMkly+JimjYn44C7VB0
hMTWMozNwYIuDgozMZ45Qh8PMg6eFs191qfr6T6y3e4D5Nhowigo8Gf2OdBK
OzUwBA+hJImo4mKB25Mbhsh966nx58Re19DrlFcHLROqWVh6HbmV9ebJ8XZn
jB8+WRDsY4qc1mqZhhUWsvTHqJEvASRczNf9w2qMc2FMeZW8MlmxSALOwJ8B
zWGMzm/KF/zkKNBPzGbJZgbxkPLAbpqDUxHp+HlbHdAx5B4I8bxtWYtI42QY
JgJBT/nNMOQQBluGAzeMSrFLuzCIlrPqmqAeKGWlRIZCvbq0lQcXwfJctyLv
NbsT2EjgN2uX9fO4cIbEPaxgFbWycWeT7x2Q4aFfHpaRq+6n29ftKx1hWNj9
q/nB2HnIRmSXuDZHTyU91vyj0QOGmWN3YH4ZOufQ6g76fXuG9ilcWpICg1rX
YQHLknV+GRFYZJwagTk5xObrX2TszL3Hr1TsZ+fqr5X5gVF2kOMLFqb3/YmZ
LvDooTRKe1GMGNf+DkaqAC8G2epL2MMlNRfgfClMqeRvpXBzowtRuR10FSuF
GxX2FztXcOJlXXEEqtXcAtyPr0kvYEj9NqgPI7xVFNlFuyC3L9AG7W934dgm
Br2xGtOgcxvXLFBAPBtWwEQJ4+GiXGzsO6+YJeOw1hMxaG3YrCcrD/Pwn/nW
KKtw1EuExFF0QulLFBWbxtBnS2hkzAXZRTy2E9xNxLtcbT35yiQmscIa/bmu
wel12dbR3YHRa7Xo/j6qEOyL6xeAkfG3bmma31fgcs30XUw14q9r2xxDtRC8
Ut5BtMyA70xWZIUyOWg5LjY7+iCJRXwpcPpusrL/nqE5oJyKmHQ547B/MMge
pQYNO351168t/D6eUE1C8Uz7jl9+XiJ3zsCrgDXeH1G7sNJbPpGkWeWBy8z1
iwlA+IyTIHmfmezL/ThbLU9uYgf5609nlp1S6yVLwZ25ThrYYLz3Ab/sKmOB
NAnPdJERF0+ZJVAeNzOQRVk49RJvhgXbJ1aVsxKvlVtBGqzU6MLhmevjDASx
HyF9NatpsQTsZXXH14zY9Lv3Ey3T8nJx55Leih1Vn7KOX/H77kI0amZSvnsj
Y86egdLjKtFAMIYt15OnRDLou66H1iDONjLNuH8QXOf/+bQ7UaIytvmT+xQG
07ZltFQrvHVJpNaf/Z7GKY7DbWNBTRojzJ3DDbjQJtT997Vn2qH/WHj80bhi
p6laDt04qtEWdZY2hMxBelUX49DjSMHVVgT7et4fIIzesYOAxGW6npFQDrRl
d2z9xJuaY6qYGSmz0OTg0oq4UoMgB4ayP0idDr9HYrEaOEWHEtD2KpfYmBFg
sf+2lg1o/tEeIwQiv5EjRHZ+7VCcwyiqF+sLEjZjBwUz+6aeKH2pAh9hqYai
Q8w2FXewpUCH/SJeCtBVXaBpovfTwXGp7vpC+z6BCyGs6l24w9nK7niVhsrL
hov/pJDZ7vqsWiUkyczdkU1DqMJIbtq9Hh4ZwyQ+Z/MZ6BI++4N8jiJz6bKG
QXd4nGMJjLlB/CmM87PE2wB47HOBfIJNHlZIajApu4LWwuylkBo6w5w1lj4C
hYte4CRzW9C7OlLwQf06IIe843KFoyrHcQB3ni1YfiXEdeDRMxi1LmKxduOw
Qs8N9a7Pb1W1b85SNOMhH6NLD1ilyFTy0lehCZVifGVUQs1qCvajEeEwM0EA
6xtrh34UzwXVNKzymM6UBGd4X6LWH2R6WvzAPvwMtP3VxmMXcduqgwgFEjJD
rrwV4fj5Xeu1H/KyfIedkwrSQKqSfV7712qyUfNq6oodyoWos4Jq8TgMgHmW
XKRmcUjdn0sc/8rOkICvdz1Joml5oNlvhw8B+kUZoxwR+gZRvdPLAcHRa9wC
q9D9/jhr+He6QTdfb8kBlgPBKuNO2E65Y3ZdHHmJ5AelSfZtJrYUHVs1C6+9
ANNNd6X4DMtHAsPH93fc/UoORN9KNPN7+M9bH8J3WfMHsJV25u09/yHiOX01
BfjSNs5/pD04+gJpxvBt/4n2IFbaZOtyz9H76caboKpY1Lpy8lo5b1K+ZJGy
AMdX7WxMoCtaAGXruzUsNdLYAvJbW6EimWiJu8kc509kuRu/PLwRhWruvmbE
vkcryffS4Kfn3F8GIAonk9E6U0n7fXJujnByAyXlpfi/c82nB5st3hvh/z/V
698hyfjPXYN2dt9BQLmZiIOZdsNrSpbRuAtco2tSA64cRalHUK/fWODk/B4N
bJr5fQh6I0czvuL8vszX7xyErRPj21Ud3Bo25Tnj0uQTvKS9D3IXmYiV+fQA
gqPwPwhpomvKxOVSJtypk71Qff1fg2DdkzOwb6Uuvfy6E18puL92a01KMRow
80nTm83Huo7M5iGSk8GOysQ2vXKXgfoJ1T4FPt9TIuzC3GEc81ZRRA6saM+j
A0x7qR736A96xdKcFIZugNgntQ1jax5QH59temfTkv1kOJDFZm9xwEcW9DJ1
im2RNAf3EhpitgKVFjMtzRMRpH2RN77+0MuQoq62Jjr/XiTehkjEyO6f/Ump
HPSj2JI+o40QrJdUVJfMx9If5ArQqnWNFFya74vdtS+TJPLPU/vG3Rt45cvP
NTwps74D4szUImO+RyoT0wREmDitwEbg0KHG61jloDOKPAgZ/VqKaRhvNV99
DZO7EZZ9fhYNu8U08Xis7zjitB2YYPnp+JynbwgAl+AkcXNR4gFLZag5ELUU
0xe5pQPVnqGVnPnlrLY1Jg8c3BdPHVF7mU+Aarf+zIfYRHvLmVmhJHiROzSA
l7ejefBCFoKbTwtVl1gn2mxcYa4CnrYU97EEd3hitgMnZMn2uLp7VtzF9QXr
w7J73FTeP6MiTe0jvAzxXAga9q7Q//wqqbOYVWULRMXBdPNWgcHTL4cXhoOB
tEfCb8sPF2bJ5KQkeRfDB6aIcyvbOWGulg4NKg1pFllkqxYHBoUIXIaKPXg2
S+KWZatNH6Uz/5P4VwA8WzDkoLIY9ayfMcEGfxdnweZ/KmC5/O9BWhLmhpZP
gkPHQrhyjo1+HdUQxSqwPMjW7ygtXfe51UHzZReDYbywBDqg4e9xBIYswspo
EO7LebnefktGPqHCenLXIG1vBS6ar2UlcZVGpMSOvTAzZatHAIBOwsm5VsRZ
gdcJ5YwPn9D0RnPGN1XITyuIK1GwMZqEIcnmDDPh+DvO5gwP7MBSt5WCKaot
xe+fdZ0e7oi/OkPC2Q7UOaobqES5X7DcIF97zJ5I4vCuE50Z3fbzqvB1vxH0
yCqn+OD34Iuuv1Nx15zJPSKCkADCIlmN777m+G5FPK39miqJ92ttAhPJe98P
uVtdGyKajzNet7t68CUWt8D8BXEsGCrxe4o5m0hvvBlMoNQDu5E1857xLbz6
OQxKkjayh4BmoxtEo40lSQOcg2n07QmbNOTi3oGNfU9Q+OUpWI9V9Z6mNZf6
ld+tPhLA6KFJlVueW6BFo8PHnch3P8C5AXSFikQ0iBkF+lI/PC8DxCN6E0dP
f59Ky+PFzurd1GavhzYWzBafkdvyXz1aJCVzEDFy748maAI8vcM7ISd3q67N
BtrYBoTqm1nxUFpu+uEO5Hp9TEy2/tliZf08u6DqdVWuVxsLoTq/IVaV8kwq
kOB4iGsQHGrIaqn0yKamcTZtf1Zh/maQeJR3yOLN2nr2DyJawkq0CH8iA1Zc
1FIEvaXU5eXYJm81os4t63JT7w7guP6iFVaTVbacutxZ37JnCKikLXm1l8FC
W3Um1K5/Fgdnt6G+TgnkCAh+08quhJpwkmY04UEn5ErQyGL/os4nj/gwj+It
u1b1vCB7IBbOblroLCEvzSxxbBXpbfW+omiWJ+xbFcFLms6JsHlfLVcAmMBW
bgZ7HWCOPsPjMKoA1ShZH1zRq+GTGOrGN9pby3sbwZ1uo8ZZm70909DRAbBk
GQmB6F6VVTZ1TXZChAwJAPcw40lWPBHCQPsLjTheo8SdAVLp7vAc6c7ED4Qi
1PULtN9u7yQXldJUchgmMLCLY2vzvXF6Yp3P2+KOfxTP23cq4hP8O09qSR9x
pG9nZY1jcm9vAhKT4bZVcpZZFrEYCuNELzrBn7F6iG8A95YQxv09sgHf3BHY
4lWNXbBaWeXMAtYVB13TylsqshzazrorjuLrT5PlGxF++tNRP+8EpWtMF0ju
DktvjQC1/51ubWwF08COMVRWzFVSNARNJOuM1+xVhziecKWmdHECWHpX9n0X
3a5UQkidOZSFN3pt08zzJ4Zdw58sScx5XnTu10jpapwDzm62MRpj00BYprN3
ichbg0qUfqUqPvPw+BmeY+WmPeGYTERKoB9OUP4tE9QSOYrtWvZ3nKHVHUyM
fQm+pEDIRvGPoR5cyoLydcEzag96GRmqBxLMENzohNi4xuTQ2nh78a6Gpw2l
dutUUQ/gYazvHl6JlzHtfiQ2W+NB7Knk8SGtFjUhc8vt9t25j5NDjZb7xiEU
0nEH1gmFPHTuRMkAlRMS6rZBesM4d3pMAtNv1f/mIxpgk7BwNulUB/lRSiHl
ZOYskpnRrhHHWGINVP03rYExEG6DBeuP9NfYEzwITShkbXy31HjgYIhNh5IF
Mt4uboYCnYiV4N0MypihZ2YiYXBDv34nOP56p3b6Yfmba4lix2tUwMTNHuod
NMhbjIdWhMGTbB42NuI1E7wwp6c/emua9BswKHM1vratcdt3GK9K3ElTP1bD
g1pNN+gXkAjCag7WJqARA9RfKi+/15lQ1fCNEpZkhHjoa8EEcMA7Q8sj65HM
6coRarsNC2hPp5RAo2MD9XvnpiObejnCNWt9RPEF5scE9f92yphfIgyMGLjm
7iF6nCitEnheLgAyQk/Bt66xvT6KLoj6tjCTC1qvb3H3Nb8nFLfOvKIy0Ns0
EnzquNtQ5aCr5e2S//w8Dltq5HQnvv3XguWXLOmCdMUoG8IZfxJnhwHTgllM
7vE7xUUVIZmVao4QQkslSuZe9cbxp3KQtuwFwjvE6rWlwMIxF3oj4nThIuKP
bQQpjfG8cX2uVOAcZwfqGEgQxapbszC5ALB0nU4bodLRxCJ8lbvkIre4AZS/
VYuvwSwHpV/us0KB7Q6nZdHUheK+ZklwAOEydiOInlvBM0vodOtgXJU40wW6
btv4oOl9LnxGUWzoprBHl9T9oETp9cNSzqdW2K1EidUYDyWjJaVXAbOryoY6
uT4ksPKuVyyE9HHtIUnAksX30DYafhIeRMVdAJfctMtDUA2P227ShlCLJBqv
U1BYr/L+79/QW4MlAH0c/8uP8c1Fr0zctiZL499Tvxy4STZzejCSZeCzGS9L
9l12kg5wyHNmeCTiO3vwGDml4pfRklDvh92f7LRTjmx6r9bIqy6I6NQ1VoeC
dQs5A/GPIzgcoS73Q1NtC95rNU3mMV+8Y73yks1XuwFYwTCtje92rJMe5mMf
20aI183AJ1QXAZsrjb2Ynt7fgFAXhm9yB/P2S/FfiKWa4ZrgEe2KWOuyk/S3
9/D3heNc38nNt4TkLNjhrO6zHRYCSD6K8RP02HnSf2uHNcdyUeHu98SMIeda
4l13iljtkNkIQEppRtdu9DmqPFxFHy8poL9TkVwJiip7pn8y+cRo7U7nSp89
4NLlspOjThnec9ZKIl1Fz8Ma/HEzY+/UFYUyACcefKKfNgGhCtqqP+l9wmUr
BMJZCGXSM0UjGULT5uZx0k5Ljgs4S/J7Gb8+eyuJkz9m9ymHsZqnXJgLVWBs
SqALC6atHZUNtg1ygaGpU3XeadTpZGY9qsoCjTWCoVNFqDafw77Z9Gsc6mMW
ao+EIz0d1e4Ga8lhYw2RWN5EsEJVx7tQps1FG5+gPSzL8hYRA/A/f4Ix55Uf
7Zb0rY2WNeQGOoaA4kVWrwERej7+hMHhqZ92u/P+ESYciRKFScVyZXC2Zd59
OEv4jrZeDfVRO2jp+OK+crr4eBBgG+hEL2moGDmheurvtPhc9XXr2DH032ZF
juCHa+lTJs927v5GxtXWgwVtSjCYzbFBVTqOaBJ/GwpdeFIwxCOhUznfcaBF
03xZmAwa+/GUzEl/CbseLD0jesa7CDyClgRw5ipx8gZcK83SNXIqVIKD0tI/
sJl9k1rbBeRiQGC8JFpKF2Rao4iJXzkHJZtFaUzGXzDd0FdJDtnAhb/pwRNM
jmoqliaH+JUFw3oyxStSms3Ra8pM28fqjYUkHlBd+8SX+fcGWJYG1Y/o9UGt
LIUdT9dMyF0ulRpkt8/CUQ6PHoBltkkp4sPTOKdguOTEXAkrXIF45HzfA/7x
7xh1vV+XTjakrLpy2NS00G73d33LaRDi2dxx0OnhM/pNhEW5APAT4EqBxjAx
Hu0i/nYuClxDd0khqquEs11GQc4aXiovSR5abaMNVns5CN5xQcQdIYKX0KWL
fAVzztluqYaInBf/W60L6Ad7zzcifZ38AKVd/JQoeAcyPiBrHAkiQYpIvM7q
fyAiPpVJyniQ45YpKryyfFwXaW2QKmC5/GAoKpfDLdYBuFwpJGoCKSvRMPEt
Tl0kijs3w87Ut+IVbcoXCLYEYFEROJos1tWohHdCtyTm3xObj8mfk9AGHtEd
J+N7+hL+I8+KVybTcqg3ppoK7X7UPSwH3H9YyjYW+zYxRXQlrcjK7aZqRTrR
7Ys2AI99kPV1W+EaATzRksa8yk8DLpBzbXdMOY2BcD1RHfHhFTWnNuykQ3z5
iHCffoSuzBLPwAbDJ/Wu3nOrBQsJRc230zrV+9iQEaE1s2cEy1WJv89qzLfs
HAEvsCLO/OBxKmqEvkyfqYiNineomLUDqeeNw+j8ftv6QSf64+eQrfub4ARF
cWDwqbCRrU5TlFPArKGGuPN25Pwvw/KuRXDfJW2LT/QUoyXfz3vPNc7lvURP
m6xGhXR/KX/T3ono7IPRhgfUwv5ptX2NKnA1cHDXC3CAMu3abFlg01oNRH02
ayFw6S/BUmo2gyD86IEsOY0zHnDsDs+TgWE0CbIxhxoAWHSPs1jbIVazQu5K
8QrBm42o3pdIxBP21QUZRsD3u15QiLd+hVZ04HwiaEQtp5vl4psWnPoYPeK3
dqsb0NkVvoKlW4RXkvkgvWcHJ5bcMOr3FlXwiwTkVxgQsowO5zvjEpVaYVKs
9hhdPSBMWFjzqTfBSMSP5ggOGT4i9jEeZXSJf970H1bZKzxWLCt5TINnK+Ep
hBdnVSR8taNYFqgjkOJ1VCx5fmcrY0l29yG7H3Mgpohoqj8qhv7QREjn6AIk
w5SVqaUU2xtyQbL5zPbHNP3muNbyvAc0s1cmwzTKFzXmZRD4SvXsSJT2wF+N
HgEnk4ECHuf/Rf2/5Fq07kDeQn4rjMXs9iol2asTRNSu5THzSczEd8Quw5pA
Kt43b/IztustOv1GvOcyNH3CXKWMzJGpsu6h7i7D9a1SlaQVvvr1M7wxRv0a
3cqoIZmuFxCX8sZgZtvT1JsOAApILmwLvJPTGe1GqSErdA2u5A4Tv7QgCPJd
VnMU2q1fe+xjD/DXGsrlw6AXfEVyT3iDgrSWiuglekTkZp+2669bc45k8ZAk
w7Z6vsH92oVndac346sH1fUe7UMpoG2PF/sKYmNka71F/x98SSeEKpiwMvli
LiVoS2x8z0YcjABa6RZTf8CyIhNNm+DpjrGqDaPNXdj55B0qPeguof4rsbHU
2xqUy2OdTGPpqOV+RR26oIsoA4oOj2DhqwmiFwKJJVqiF8SiER3Pk4gnofbY
bY64jX4gQtOarDMtAbVKM9VGg7iuejE5w4Y7bKWd6xNjuyB2Xe0u7A8sM016
u2zswQZ0Q1t0qvRV1fm4/Uw2CQvbzGJU2twXTTVBMccncAmkYVr/HhiBihGR
qO+41NtCjt8w/qu02GXk4LNBxSoPGZxE3g6pmjOBGCPWaewk3WQlLhWvBfw+
R4cKRNuVW5M5W8yrpxS9S8V437fjKWFP46b0n9dL1quqkoLb4wQwGskENv5J
8SUUCDD3vURanf7nx+LfK3/RqfZ0G0VV8hzFH3NIaFRXtowp/fE2/EmDSvip
jeVhfINOfmwSpT85xZPkThswpH5bBa1HBzmFZhHvS8uDzwx3XbOg7bZds7bW
Ldhz0h5Ti/80ziCi3RTiDmM24l9UC09OBum5tB711hMErCLDrhT3kCDtGu5q
ESprUYElZsjnSxyT60D9e69VblHgkTAXga+hghAydyTaxs7hlcz9JHkOVsmA
UADKvuKIIu/jh6ABS2N/rjdAREPGnanWPwCQL+x6kz31D16IYnlO8pl8xYBa
mYL5kmIOg9YKwUxxS/L8DlOKSOANDJcaBwtuQW/pEbhHqshfoI6dyR1O2XHI
Z+YQHwuZia6Y0kCVRdJuNVD5WBH23Rw3QdIFVLBf+gFGlTOFNNBTFCkcXveO
uUJKkYXQedcMD6BXH8XR2kCEj+KYqH/MM8NWyxmUEkplkuAMxUeI46FheMV2
uAtS9n708WYKt0/V7bSjOVfMJVXMtUrYdDfC9W6WtIhYMQOVhU7Znl3tzYXG
cyQv9rZgfcZ885fLNBcqx7IxWd98dvp3NV3K9/7UlFPCEz6fPfKdBLhq9g9T
0IyV8CZIerwuDEEPTr94Mkfs3cVtAQ0vHyjTJ+YQu6km9tr7l3k0dsCb60Sq
WW/sSY0RkiPr1R7AcCChQzwG7Us33JR9h3QhjTPOeI1ybbPSpQXDO2VLsBOW
ZcI6UGImTJzbmbJeZpXbeTCz6Lhsr9q6RUfRoe2EUul8kV+Rq/fi6iBd6xjM
1ZEzMHfEF8XIUl4lVUYpnUCH6AnuVaIAmbF1FpaExxxcG8wGhWKgx0jtY3M1
B6J/c1quINyxjBPOhoGwzZPrJg+Rbc/vgm9F9v3j/dsYMjZzFQgmCjgHGF09
EAyqk/chRAMzbkvqPQ+IXCKB5OOseyQQMj9ci/x5eCfMdsM6pWvygmPoyMu5
UDsRx9hdovrieUsZKUzykmM6WucGKT1KKYJ6yrzrKsg2CcsXThBf4iBvzhd4
WvEwUETjc5VMFSGQ/TMBm5eqJnUWWfOaa4Ncd3QdadwU9u9LaIVP+XITmjB/
jorZ/NsTzt6/m97dB1rh/YJXrQ3I5i8XxEttRMDNAJZJg5LLw3iRUcaOBdsH
nCZEZYkyTWgdAqIFsyJ5Z5Cf5B4VEvtDir9jPt8d5JvUkXVfzlHHYHJ2ctny
fURbxgAl8rsvdAC+reAOK+jzddZr4XjUwBmIS5tZDSyRhCZv5zIPP293CnT5
+fS6PvMyLMcPTA5e45PlH0Bst9JfUv4aXV01tiogjje9w5ZyYyPwHBeEQAT3
eVJLSRVQS+Zb3BUUXAQ6UKlYwdrTrkJVEj+qqAE+eRcRGqgH3wVEOtlI3dVH
TcVSo30JVFEKEuyrqvgfpIbIo8obMKaab4zlaSkwmzctDr/h3cI59YqKFEzu
u0gIKVT64ma5N6jwxOzYe6+QnQckOamX545B8k81FeOQgWBcgwHfP3In2QH6
9S/GhPNwCQvDjEWI1ofrl4+orZmhoFINtiZo0p9lN7dHPcxgokCZZPAQmUZe
DHWFY1g11N9pRM4d3y0vK2dj19MYkUPCNmIIDecJ9qv7XDgqMDwgkMNcYKTc
MVJv4UJUagOlFY9YIq8MdCqoI0cmFWcbgmeR4EV0MNq+u5xfKtCC8kHjhaTt
5ZiM1iCmQisAEpSg/fJRXmiQhNWsamvYJcGC/cu9wh2IGn/eeLSKC4M4NSQ8
bu2jj0wB02G2WrW7276AXvnD5WNHPishFVppIoiJQkv9An2FBLTfCwcXcsUV
vYr1FGTt62XQorv4b48fma5SC9fHGfPToKstf1sQVebruB1Y5jrQ2txVCoip
vCHPngKhVd4q4I9Uk/KvfbHkuoCJkjzzCkMptO4egcJ93YnpgwascAEEnBOH
FQmZ0A77aYC0dyg/vcV67eOiMEMgEl3Y3yC36DMGUniTyeXKtVvPrf51Ajh5
GABQQbFVaRuO2mm2J93zH+qEw3PZQVduc+DnI87sgiC+POkKKsQa9Rd76um9
Kci3h0tESYhpZ/ym9GaXW2Cp15tyKrdhAx1G9DMHSC0a6vKwR/D5xnRxwFlv
2+fqnnxiVcyM/zSTSMddS2o7B/dR1WT7c2gOgzencwwkUt9fZJ6qJMo7iW9s
JCX45BYmq0H0/CHJtU+vuILyQcL4v531t3xZcPMnxikCwoYT13Mz41u6unz9
3NL611pUsyycxJ0K5knTAUWWdqiu8wdc/9ADl9w+uNXEl6pPxUX1kRa+rHQh
1z5Z9yrNM19ZgnCFYu+CD8JEsCcTXvDhRYjn2j+LOHAySmVgxIOidqf+hQx+
7aWOdbOTMhfyVzlQTHVlD6AXAiow2kBLJxp0NAb0wt2cgj5nUCx1Mo8/Edkx
TfssOyZEOjIcaHF3y3AwkLGe/MoLjrA+PrCkR3afz7ox2k407Yr3vpS9ywdl
WdIDTXmDMatRZQ17Ys7hCeGlH2YQjsuvSS7/TLc4KxFBJ2q3uAr+5fXwpkGd
QXdkdfTexKzPCFDkx+CJj38/olfNfSoa/EWJ4dVZF27RBD+5MRDqgJqZKCUJ
NouqY6RMKp26CUhLnW/TGbl1V/ysCmfx0k1iETFIUobetl5Stz9GMq2r96Tz
/4s+bFdNM+TPhNLX9tGnMzi/JMmBAMlJQbRta7Rp7CBEUUc+KGOTIEqE7Yyo
YKoW1D+JomXRUSFsST7GfNBKfADAsBnhq29CSVjJnVB2RcdPJ/pW3QSn3dJn
spbxwsxPYCuSMwr2O36h77BJ8dMxI0eyzxqwetv0a8LrO7Q4PVBiPguJRbDO
uTzGzMHslMqzCzYyjPPBinyGOI8086QfTjrbUmkYqE3eGKzE8Q5gz3BK52Et
8wOb/NqgivrhfjLUOKKIPbL5uAuFpHxX/WDfTSRUPFLV3efLC8FCeqCln6ub
rFpSmZBpmSqzj6J/294Rawtxb4IxLbP9satQo81Qd6Bc8vVg58Zn8HQos3G0
p5wFku9UgEuhpyG+3BNxPws9KjFsFBjGCJaiFmDc1t2VGf2GxapBiMg1O6Fd
RDKiCSzukTgA8beFbBkAX0etgF1h2kKQQRpOtNvb+Idkc/iuUyJoHKXp/LyV
CIKy6g+01a3bC6+2nU7iGcVjW9uAKqxHvFxutEyTHw5/OjY5shX5wynjHC/v
82oEfkoqdI3WbcreYm7pNwUo8GMuugQOC8kvPw81/7vS3i7pgIYC/XkULSvz
fX0JCjvGtrxcPkU0iXYSPJCWl7bnXDYOnsYA6JnZiMlgHCKpDEnXQDRlcIUV
TPpGPkBQ9uLKrkKCCFUsIa8juu3bHEu/plOPaOQWXn4S6txyVbZCyjYQDiyv
AsAPutuuxE27aNTzoq2PKsmd/cIWir8d3zdIjx0jpT2mB5O8fsFSNGg0ZXd+
FUUteXeqezcFpV6y5k/QE1FP3TLEp3lmGc2u1JAr1xUz0/1q4rmCsnIxZOzW
8n/13wC4ktwFpyll9gVDqGZM7goiQvGGSy8x+B/eYdJ631jLXq9MeSvTxvUS
E4bpJ7AVmfzGCwNwGLXHhccPtRM2Uetel3HDm3OqjslVTzOB5ATXPHdI20gf
qGj5hnoDGDurWTwU1zFvN6d0UsE41VpiQydQ9N6+ZH7tSONDIZNQYjt/LwAS
gJuE1r+vIn9sJItpMCFbZzn1k/FZ4JX1BZs8KZZGHqyd+r6BrhaNaFTs9Tix
mUNyItjQVSJLRm4br3WTVKwLQLGHpXAq2j5p8aC10T1t9nVLMLSzwrloUJ/W
vI2J+DX0QONkJQ3nSY8hnhT9QKjGGv644qAN1Y4xahBJcR9ccmWrK59PEYnq
6Vo7ac70HUoEWrbfhzjsBPspD7mkk0xs98dmDNArX1B/2tEPpJV6q1xg1AUp
F6J5vfidTQ9V/MeGFlBZXMwXOmUDN17UpDvd36i30kIYVAZuN/3+mJ2NqquJ
DUxcbbmKR9EkpB8g+Holb3L7xpLJSu/oclPonBB1ZhJKL3AHlo5dQym18rn1
I+q4nIKYOpmlEBRyKrS+9pOLB6rrLHILvd5gekqzYp5n4TTuC14KQH/jBUgm
o4UwoQoAvkphEn9sE0r+ZalOYkng4IGKF2WrvSN23AW5xvvEpuelQOH4/hsN
cNjrLm6tv/J1V5TBcG3E1Cd7VDTvu2WWEgLd35FL/BN4VJ91Ia6UEL757hlr
hAll2RBcQUuVeCIgPjNTvhk900v57Hx7pbmRXW/wJzZG0RM9w5jjBI6EHXOn
SDLzf1pMIYX9SZElmq0oYMhwc6bSHTQQGmVwtXb8OjiFXVKqXdvXMDChYM9j
M4KSHjuo1OI4YUt1Aroig9Unqf88rlljhN084xogEx0LB5nSZC+evTTiJrE8
ZXrFRfpMV6RBcxVfC7NP3zynuHhs//64sqm2Ze4YRaurGAfjsP7zpyKQEGt4
X3eZuV5w1MF2qh5elrRHho4fVYzTgCQjuvW/b0kirYbnQA2XhvdnLQOI+eMP
b/QYiLZRjasYEM8fEefkZjosNpvcquBGDW/Sxz4ymBh5Kt6xxB6Iw/CXzyxQ
c5Zd2WMcaShgtshkntJkGDygc7L/YeibGyPEaA8gli6uk2zHINRM/y0EXpqk
pNB3dBF+km/OlFA7R7C7V3c2z/YAKCeYwlCxtNpHx7qucArfqsj9TvWExkGU
triczvjUo2VJhWdMIG7WY1ijrZf73Yq/AAQIa1k1pHwje538P1i0eBsSxY4D
Pwtxxvn1fLA7/u0AquL3uRQutrs+KWrTF93klf0LxN1vcA6Fk6NYAGbH1f8t
Gq6xfankXwnQ1DXYnyGMEoQLjQw2FVnAKybF15DVHWF/q7IMUXGu3xFGXOKV
DO0cQFn3EYjacygLe0IWtcg0cvBCFqGdkLuii2TUCsZQN7311Y/uWIj6cHyt
nJ7fXhkowhKpm4SHM5NZXDm79RXC3g6OF5Fe96UGGpE3TyaS5ijbAHA4Szf7
laSOAzr1nz8a4W2smARQEezoxwIRKBmAq0UyXN+gJNUDv2fsc7fDV6qXRka7
TA3Sc2Gud5/JagOFctfqMx/76xNZo+Cxr8b0UNUVJBeZtp7reUk3rdG1UXrT
VrtOo9fvOMPMPpQ58Cp7X63ALHVKjVNHX0elA2rECpZHriS1f+X4tU9tb4vk
VWEpfSDH0VMiWHMoa91pKX+sBoFMgHkoI4dUw/jVkN5S4Sc3DB1ZBQz042fU
VkQJ190v+ViFbumyJ3bEivT5/KnnWaZ1VTxbnVyVJlIR1ZAxy0LR3xeZvq1X
tLJe7ElA+ck52vjQD9GKGW3ufE/2Vss3m8aIeA0xY79OVZEShdxOvEDq6BfY
AYbPabnRPzghSjtgOpvkPUwBz5mj+gmNnDKG9gSi7QJtE8YRBRxf3f4jcelW
VsBbOtvqXBLdr3C1pQ/dv4SZNH42A2fxGwFaaxc1IYcSXyOcRpYSUNhjhC8Q
/GHLJojS81dp1mWnMj1cCDMPfGryIhjNpJ19C8Fwip05TgDE/hkgttif0EQc
TeBIUyWrF5oUSWx68Pj/j/GI0q6UgFECRJ502rw/sLAhOL8Hmtb3z9HU0ygk
8qzJ6TuAY45rJrMeRndcbQ4WApCKiQwyKKBaOFdhKCfZ/bqOJjTG1abovXBz
AnhQqco2Q9Cnzi7RceupsB7ZA63BwneMHMmMFiJFBXkdiEU6mGZncGFVBv46
+aCl6Cnz0DHNn9pRdUrh+UPZzr5Ldm+9rRLrX6SvTzBW91aEZzH0Ov2z369Y
zaAr+eLtq4IqwM/gGYKuhc1xUGV4i57XeFVCzk+gwI0bKafPjPxv5nokGRg4
Zcie1ZgqYwB/XO5/zTTL8wXK5stmS2NMUPk+equv63mFjnf9A3oMz2nwbC89
VxU4relaB6aLl5Yyy2OhNhKRH1YsBqa9wG0518IOsFkoAkK63hxeY1Snbdpn
ciAX4qm2stQZzY51oWYx0cDlVGPdYFf/YtyN/kTW4YTMFpVh6ODqPPXI+LEn
F4o11V9OhwL1PCVcj+1ATXCYl8F/lU0Q1W48g5H4nvR0V2IW12kJZWBmtDF2
MZUdBSOKrekLDCO2aHgWuQSp4nUX8jehyTUpgtNQbO+Ef3qAPhet1exRsCVW
bIauUNd0WpyzM+r1/+oeq9/mjGv2N7giUbtq8azVbcJW2LS66g3MPZW4eJWT
BU0sy7/z1C72wdOwFcQUE09lBIzFLTJWtBSfZPVLLaXxZuAp+iFY3B8WIkdB
K/qvCx7OTfU2pnXRpaA5hOtk3lq45O0OmiaPnQN7FTSTU67YEx2/i9bB3IBO
ayggbOpqYHHP/7cXWj/0NZnzdE1c2+cZWM8UiaSVZPnqLlhvNk69gvtrdHqL
IKirchDTKizr5adOSy7mI2MqfxKZKtWCLGlHajaVf7PmHCh4XWWDkefxsMB2
sv7UxQMPmU99NlHX2SzIHQC65Zli7HHhjHD1duLi6Jft88hx7OREpK2XSQJM
J6g0wwZgpcHN6wkoS1/N3cSWFEq5PXHHQImvLGigbXXP+p8pbQY2OYwKkqPz
wB/shrr5wA2m9XpFJYLRmhkITqd+3W0TmRvXEjzmIZgGKc9lveGVe2CZGxeN
192ITUs52ynA4VCO+nCvTInoH4pqCCyMuybaCkP1W/Tw5pfI6+J9uIKSS67P
c6jAR3flpjmMLaU6hb5+R/DcFuvMbZApxZYkipq1n7WZLS/7z2JnzBWHNWxs
3B/eQDgdP1/DN9BDQ5yv+JrpJ6iYER8QNkcOcOT1J/y/O4twlVbkT1k7ECWc
6KW1jQzKTsDDDlRQsLuQkrhw0sqefnhdYwsL+Z2D3D+Df3odfmYRFeW/SgCP
CAaDksAe+gQivw5oerbdKqgOySvEKBy5+CsXeM+X5zLpOHKc+lA+K/2vnkAq
tufZveJcXwKeV42XfkQ4yfA1ZEceLy/5DhI33e51mf3oM+4eOvIr/LSfUN3L
fKx6GubpOFBJQ1iptGyKHb2ZaQUt3hdsdWKhGcRcSWxJgWVsmlCgvsPfcGak
AwZyGVke6Dm206SiwkXdBsUL5fm+gK8peV7jEyRs1+FLlh2waLiKmAKmC/2o
+RACrsPqxah0VI5o2H1d5b3b5OnLahwZHyiq/6DBUByILypduFjvuhZWYU7O
uU2ZAKPfjN+BjEBK2r3UBsKz9iWQqZ99aizOl51fIXmyjo+4CBWc98rsOlXa
RsaTeL28B08JNM3tP4yS3/KEAu5NpegiQ5PIiVOy20GzQInqem+zYFuFRvdB
/KHk/L0jHMentnKhJRE65jRiWbJOIE2TiIzYCJNAIRYzGLOy5UDusFMZx95z
0lvAD8KTtDvTWdyJlef0HW2JEqraX2VsvpIr4NQcjrgM4CdahjA0wao+DRh+
OU4hy+9nqp7Kw/n9Vc4Ty0o2kIghHVfOhPVLsM2ViUFDZvCkU3xHsJygkCkg
98RtBIsndk1eFONFJJFmiFDnjpR+T5XLCSh6IiCnVn+YNh7X7tMYWN65HvPO
MiyV5BqECz8i25Nd+SCGEHgBuJ8pRhiY85lSizKk+v7kZjd7yMYWhQcpyzUj
WyBISVbJNxkA9JO/z/APhj8n0dDZu64+ZbxsdDvP0XIBjMuuBR5nYZ5JnGh7
GLtnF5XJDPjV/J0J44ouT8f5CO54cNCsh691UYh+yFJUoXndWIKXbxhI9Hkc
BZ5RUTeOsGOmApd/BSv1DPqKfnQS1leXE083Sgp4QnjpjreGtQJ41Zc/XY0i
4eC4fvt4AAX9WBP3WXIZO4RZNsr3xa2Mkse4AmRlokCtyuoHjYJTGBCS6iNZ
r3jR6zhm7ycZ3EKWp2EKboF+BpOTctY7h7nkpdzeO/DbUyocDXLjTQm9EFnc
6OsMBRHEmR3JR8vMI17FQ9WBjwHS9BM+hpkrlD8CrSe8KrS+SzDGdhwCNBU5
XjSSw3+X4h5q+ut9UH8r+h8gc7QPGua+JxpyBnVR7HHsNWIlfC8N1nE7CLqd
xqHSyabvJRW/z83gri9fRIJHpWulCPgsjsDzvLuSmKCH5AzoLinLOKpFeABf
wx0oD9wqkCrAXuM9uJBWkckD1iax3CXcGypTGAfEyHKYYD70EDud4bM+Sp6j
n0e6eYbrpJGWESdjUVhNErvBDLuuRYzPm2QCdobH4BYVUOLw/XJvVU5GaICP
7zdp3xbqTqwN+qH5EMvAHZJ8ldAkd+OQtdaYFzVAADwtwf/JmD5iYM895zl1
dEAmEN1h0f5Ytuc/rROlONTkxo9LpjH04vpUxr34HozaBrqDFl0ab+XJuIRg
NtBOvfi78yQbY7pTPYvEMNPESnVJTfeB8SKCMorVqh1SAHlMlVa9+aFK3inH
2O5RftkUB073yA2OxQw9DUT47XYphXfvCKqfCeN4xnA1BAah+E+Cbc2g9Czx
B1qwjZSM5qr1Xe22PkrOTEd1ImXwgYJo+bfLyK6yxzr+UeAmZ5je73pDDDEs
1BjeYoELOK4i5aB8Owvo3S+gXKoqB3jVueClJRgJ9Lj/mf65AqdZZIv4Ia28
2UoKbTYvFLZxRFYVFoGp/TD5iJbzGY52tY/PrjKxk+UyvbAtI4t/quvMPx9v
7dt196EyiFVodmGTuqq3S7vIiAT5WQeLTKMRsSKv8LcikdVEkRr0g86Yo2OW
XSODjPNpP5kTnMzFv/AMq0/y7PV9nPqxjfw6CE6d6cg3YFScjZLOVeMJ7vgS
3iLtFdHh+eeW3RwvgOQhGgMPsciW7Dl104+9imQiAh948Nh94VqwPbyzUEpH
3KAfC6mKgGpV7EdgJXAtD4Lh4jL9khy6pgZKBiz0lHXL/V3eteQhYVuZwz1g
iw6iJFZpnXM/LDZMJQGmBIkMXtVnN8Y8ftEczAqwpMcR6/KpdSKwf/msH2n3
uIK8hOptR8YUP0I1ocaXbdIOmNTBRt5giBw1aA+nmfkysqRV5SQoFXUabXHu
TGKlvrgVrGY8y5w0hu7R+iYqfiZ4ahG2v0KWvTnEX5N0JYlQ6sy3UvS1H45K
g4YeiNGVGoSZ0ixCeFXwhRwh41qzAz/GL8BbBTqQrJ5gzXLW++ORTEdfWZ1E
YfkveqQeVyKBiqZuGHTJz+/nrMOP0josAqW8LMjU8qMsH8Ipx1GpSYXRvaqi
J6K8v4gSo9xJHk+b1rziXpj7Gv5AsLP5xdfyUYDaoFeVhdmfp9noPTkbQ23P
hr+wL0ZOv+w6Rfv6H0bhSPbm6d8+e6FyNVAZY7GH4dSQkGNnRfYtV5vLPB5U
sBK09wODiQdRI1MlWTFECOJeeCtABvz1107DnYqQPJzMwY3RHLjBQNKlxCnr
igh61aiCAsjQsXB3YdTSWW5BoPXnazIavb6NDP6CmFAVi77evHrT7f6TUfMx
FUC7K+N8za/8P5srtCQ8RXqTw1/TvVzBg049iFpxa5HIpdhzF+7kJvHduzL8
80yFOhBv/qoHOY45hlgLv/SWi7CYSnfVOsG4O3JDD49Eer+7xHZJZHZyE0kA
JRw+m4hLoftHHle6A7rnEA3l35pS0nvs6JmDWGq4qJfmzoy27UC5kexVvXFB
L8Cp+sRNcjEOEro9vjzT8f1nCo15kUtpff9n61qflZDy4A0iXn2ZLVFqQcPO
JgjeiylVu0cicVleNj8wbpji6KuJCQy/2nA75qeivctLAx+44tUBoCboXghg
w8MYDyFtsaKk+eMaFMRtts5xK6RXqtEvkA1MFUMaub2PKQOG/GYCB6/xuf/D
Gk3K9xsosvMKyCl/oBtbb1SAfMeA5U1f5OPkPSrlMJhQmpI3CrEh3HiFmNtd
EiNYGNbnX/qJ+ryJJYsWT+26Wb1ppDTYMgcTDayElr9l/pVbMe0rLp1UowsF
1rLxLmK0hgM3AaIpAp5Sm0BQuq7LKVrS1qvW+lCJQu1iO2kHPfNUWdf3LDLT
Di+vbjTQczF10RFW10cw3NqvHEuM1BMGqO+Kfl9zI1slNRxPz99r79orZ6Ds
cVM+XYoYOJjy6JlYp8++reNYPWTbkmb++zFgursxuLCpvEfxEwUSAeBac3nh
pwRzdUTU/l7vE6ETTrVDzA4r9qHMXCed9wJIfNRKFB1DXLTYmTWJ994IpoIb
q+RPrCWqnFowtVuyhAXIw6fYkIvyepyBGkTH+49Cyrp2pc13e1FPqrAzjOV0
ee4DFXH7wDhhB12FewlxD6eXQksZXwhUgXxEErsTh89CpfAyEeWzLjRZM0TF
V+82V8/B4qG1d514LE3KsopNuTDGZvr/nEVhj1LNqJVHLdFB3PSTg4g6025V
IeP0sMTPdcatN6RJP+DvPnunkF5PIHGTk896wJwjH5i8DlAqSMXAqT2N1JVl
45/qRBO3Q4gNs4gb0bovqgmRzfbX2cvkErE+1uzw2GL3GBjJbDJcvgbpWMld
cz3IwtJLY7t/pFwebcWEQmNNcclkdmoCLLRF7A9wR67NwxNQSq5mt8C7HnI7
kiaDzVO+O+Zhb9/M7EMfU5rNtRWXGS5g7aqpvoCZ09iD3xzLeFDQUFKGGOgr
5e6558U+4ql2vEPKa3j43YR9+u8lUk0QV2wqYpdiycW8c7c9EXLJudQA9pF2
D6sSosQJKq6/x8TXVsgDcxNySO9bQxMJlZiW2deMaR5sPPcZAT6ojz/ByCbY
7wr67t36d5xLRiDWrJ9RHT1krl1RDcKJK3ieF5GxtmeXk1jp20epp3TdCCpJ
QglnLjhZA8LNR3KWmIA21yC2uhOT6XxGppXUrAIjrprvikURDawoyZdn8zRT
y831ZNrtFUwKuPIP+74eDV2QfhoS5O236S54IXSBg4Cn9YJ6ZDWI53CZRwub
0Rhz74BkCYPhjW4nM/mzLAh4sCJtxTLuVh/dM21y9DN7vj5h7XMq8nuChcy6
YFzufYWP41Ek3dSwxLvCoR9tgOIfzTQnLIA/fzb22eRIvwijr8nQIX2kKo4k
eoIVaAjMsvBfDMR8zavLpS2KIODsu0oIDr4HurLbujPRXG0UXEbu+xUpoJAP
L3DBtdoHyHUcz9tzemABiUF377fFMJB6u/a3OiD2NAzf3yG4eTOLSn9u4mK0
AaCEMko8cyoU3oAJ+FQ+3kdgPINaKeAkzjyv1gxccIeXg8MlRm+MQQPp4jwd
vQ7DwHYzTAMcXDhTQgIXyB7Vte6X8f+/zhBSrEVB0G0UmKHn+rm+v8eBgKoU
60C7V42KusP8Ciu+LbNDk4Dek53//fArr87x5ZrzjSAnn8THLzXyN0yYG8a4
fmWBehAlAUKH57yArD9bseZJiogTVw2tL6SmdciQAGwy99WeQ2UdTY1oxuA5
cq4U3bz34TWL2qipz/4wPi1bjQ4xW5HgQzaatA3FFTjY7x3bfc0Nr2TSfsEf
OPaikRunTbyCWR6izYQJ6oeh2dIi8cmtPH+ynRRXM3sbceUK/kaal+sIgzBC
NvlYesZLxTGuJZZuBsX1OXXlh6JySXh5IP1KTFWHGsJGBR+0tHE58NaiZSUW
wiADBfV68Dxona/m2i914I8isZbQDXd490Ld4j0mHlkjLJe1/2SBZb4prRle
hwKZi/pk6WTErTv/aGHCv6F0KreTqnQ+u2E8FeiX4BTaUm0vmOfSNq/OG8f3
nLPQvJvK+0ulJ9brcO1p4a1lyETfcMUDFGAbU/9EgNt0q6hAsfD29NiZHgzq
MayOnrFrxJdaZTqObxb4Qz1EeYDe/hVUsCEs0Wq+bV0t/DWPz0r2NXk3/Yml
iwaQfoQTpNc5GNYMiApRnF/7O+AgD8v8onUmW4Z9kKsrX/8n/xWuDin2DPsl
pZNjsrhLzkHUX84ZIeGlHEjcqSC6GsJ9F0LuFJgp4NOOx9JMrgKrYhqtJRUH
oLhMou9QSjNxZWt67BKP82wwnWbNAJiTIwvmDSKuYqqiZ0K7aRov4zeCUSMK
tHvacijWVjh1pyjaFDYkBI0GCfAjYYuA4Wiy/FT9W3KHA+cNVIoI9rVHrzXc
j3uHW1UDyiQBJ3HpF9Fv/DScyPiuCuGCgPxQhBxrUEQp4jTpE1RILJbUKnpG
tGwpdcyP8e4kzFRdFaQdOHvzITOMx7seMAN9DZ4LKyOdIc+fpmr+82ZdOJcQ
sOD+Ezcqvj1UOekFUK4Pj8d/+3sEXB0XM2GCmuhQhwGUGE8NhLf6NBrCDE2q
PWQdunhx03W2S0+jsIBqWYM7fY+Dc3da7zvA9bYVy1J9frjtdQdYkUyKzwYa
CdPu43gKnQuRvtG4bfZNIIvbnZwlnI30G2VwKnvy37D78qoYrMiRAcI8nDX4
34syUu8dyKqJIYpqLWO7o9YxuzD0VVM5di9IjL5ROtfYPbVC37Gg/D13U6cK
tVZgSMyQ8Mp/JhxcDOtM6XAepTuwRMqZm+g+mcdjZkxpTEGuWTSx4kWeuYm3
wOlkBYfPyorI1tlI+OFu22eS22D5u5NzFLE/qzkgWA0q0H75Ric8lBjNKF3N
yNbAtcV5LcnivMCsXXYf4ZSSuFJ2KYDxIVd7lkt6M4AEXd2K1r2x3Zcgi18k
daOtudeHu3QzRuuAFPUDd4hmpoPEUmFzfK+6vTHKutv+z+mGVnt19FVbYKrX
57WZq3NmcS6CjD1c4Wp/vue3if48OVo8PIM/5Spl2SDl+jpMjlmx1Vv/SyMe
vJmTfBbP14X08ALiBlufpalCA0KeXL3CbqEBv0MgcJq+Pb6N43kJkXgbQ6S5
mZXt4jlc/FQGMh701os7L6Ewc+6qpIXmY4dJp8z007RU6CW1Xw6NNcDa36bq
abBpk3MBvQ5bV3G1na5GwVStQgcV4AKe7q/M2ckIpIOC6v3Lng0ThOCwGVrV
2eyS5Ps3E2Y9Fu5CBXWQhN1kU1IXzQTShdP0ed0Azl6rXU8fadRPlDAFms1L
cUwd0Zyo0WwQ8kHD32civbpWzKs6wOfi6lyInuY3hCUsMT54HfjXhslHmizh
p4EOgRgc7lYRHcibJl+HJGX5+gTKE3DyHo6D2hVQMga1gk6sDkZSN1xPgTZq
XFD1ZEr/XOFF8M7I7FOZ9+SVOcq+7ph4ygv0VnuMsjVTlHLFUrPjRDrOk0gn
1SU/337qiCKtT+CfCRdcB6srkoiJ3n3letlrK33Ywr+8M/nSMbBTSXevum2X
D6uvmKmSIu5YEATt3opX36Z7Zcbmxk7SIbRMudzt6LGK5k3GHP9ay148wUJt
PI5srHmUoh5S6LN3GeL8TR/04hxhkpZuaLc/SaovsG3z+rXcYf+ZUYtcB577
panGpbvU+WcbCf3B2023vkNnVt01Cxzf+8R54u6JPaEiNimYI9kCgtXPm4OI
3WdHOuXSS/dbAafFJFPVpuFc0+QULarQCeKXer1/l3t7PaDcJRdUc9KWmWzd
QxoP7ACQ6SvaQvbQ28VGBU840lt8xpqp5oiGDNqJ6FPRg3qlaiqWmabwooBA
v708hiMYYLE2Fr0o1nCa1BsEe4WX2hnXIRCcrtOY9IJjtTQYjpdJrLR0GFN+
d+9pqVPSo9nQDDgtqotHta2VDbzQEvd/Fo9ILzFrf6Ury1KMZTfhnBi/POaP
mxq4Dc+niY1nhgxSNZdDAVjkvmU3I/SYt0y7NdjAW7BmSQgzFkKD8sebNWaE
SAUQMRyh0rBfejbwX07j1qyjGyJgkFDOw3FA46tRrpS4BoTFhxKUSCHzkcl/
GLa7p+JzPLsiIL5ECo9F8ujOh15t6uO46wZxP9tqi78CYWX/IEphzAzidiyi
YTEGGgCZ5KJmxaWy4F6H8eZXgJJeA2Qz+X67rdOe13Jgm6kpdb/0Zf8RlrZ0
zRlSwdrYI84bwAS5BYEDNXHHbjPSOD29V9X25aBoEiYL+4guUkPbe3984Fs/
3ZYgKZ6/EzYpHZHDgpF2i7C3+w5t1DxkkPL1ECrdHfXXDFAZUQNTTYlvNvP2
rIt57SYC3FrgueQgKmExkHxzlVSZV0fIn7fcQN1Q2RrJNy7rCJiJEn0nKKIf
gPNEzB8M4fAd1Yel0nStOlRpYhb/32h5Pepiyn3T2WZfkmR3OaK25f2+oUAV
qEJ/NsH+LB2oZpaRVqkqcA3isl95ul/F7mK0oddzENgs9yHd+Gl+EfqaY3YY
q8Uf9+rrxqPzHS6JmjliOFXp3+rBOdzmFceF7nb+Bl8/a31Kk7rbwkMglMeF
acdAhjF/XuPjTB/p1SnvGa3MCHIttNGPWkpggMExa2mtC5ofA+EEx/8cTIkt
GnZfuGbYaLxJEP2PA0nJNaetVF9VTxIdjmaNlN6HIxM9pb+B8mrlPI4du2oH
+l09SN34tiFtwIx4D2orCOG3xz1v2ZTgDr6JDUHQA7/1MN5YmJ8IwMbibdNw
pc5egtmICA6D9rOcZ3zWg3m8fyngvFhz7NjMHLwHE0vMBxO/27qv+PsRPKaA
PbJYOA+GIAq1zfspomOKW8BToOyUWbWP6kKRTHaqUq77lKnQwTUuODgRoSH/
A0KpqfziSJPrPwOFZ7vY9bjOF+tqZ9A1fqBMxMVzKYKzvSWbd63IkxPyulIY
JLeBhbdX2bjURu5P8tH/BAMCesRFLsELnYVzTg5QMoEWFBAho3dBUCJ9JfQp
uOxo41od/T/rbirELcags+iR1laZN/PhrGmtqDRp7/Uqh1k2C8VxTsMEQk2o
/t6ngIVhtHXy4YU1q7A/4/LwKzekcAxl//6z6JrtUvyaoITqWutq147A6Sn2
D867/BrfkBHmx5XuLw7ZoddW0kJksITcplvN5n2Ls6rPaLSH0znwUH/ROJ7K
0Lv26r5l0/IjjDOJC78TjGDHibdKRPhnz+0+sL2oHjueksllYz6FE33b6SAp
llTtc3Y2Bel/uEYoaHQaWWYsJjj5tA1e+grK1g1c5L1sbAYy5BZePQvt2E4L
2n0YRxqij8FP+4ZNVRN7j+rCBC7Tyw5htik9cOnJFA9+ZW+oY4jhwQ/HKjzP
ubtLQ5+LpSllT06WQKUEA0oguRHfErJnRXYmGDhw2WtuxusAQsMOgiATiebR
k3eyzcP10DzDPXS4t+1Qrokv9QGugkoGRNk+esELYzLBHYuMuiJi5gl9hKzd
RHxP8zVAK3XGlVevqs7My606F3FFKNO0HepJLzQBOrtkcel/8nMrXDjm96np
Ypg2edNVb/2gPVvYaz6iR36NS1VN/BEK3VIT1Bo+/0arXW/QaxyYyIm7dDEu
v/yyiUskWIF4P3JkovnhDzxgmq+hs9LdlJf6a4UOjbrTRujwwQ+x7bXQv2n9
HAkWYxlyvMoJ+p+ZKMGh3Do6gGDMiCAoTIbF7T0umvB/9uju9EjQYba4gRFz
iMR+leEIoCFlPIirVcd3082kYwe+wn47MP8t1i70jKgGhTBLXCYDQhD/HDYm
tYx4FCPF/C+vd3EjWaDj85RBGrVrPMMnRoyvQN2W3gN9bp0id+AH5EADVXFK
XRNbSZ+3Pj+agJ9+lFWB7D2zzyMf+MibR+TCw284x936Ev3DNgJhZsqfhunB
W9aVz9BnDfQDB2eboWaXPK/7z0J/nm1Yilf4yG2lVlhErI6fSBXezlbC+0Le
C+wGsUQ+WmDI8cWB0hP/lIVYv6b98pslqMTF7ipYWAas3ae8RWkvL3cYd0Fq
AfHueoGcqGboULEgFaYmjOy49/BMYq+7oRKzFyFqPbyRzh1IjZEPXIeIQFu0
WHLFrK22wSAr2DYccvUV6XQa2EXELj0M+iGLL98C/ahW3kbWIgAUmtEsag84
hV/myjTEgyfbhDTNsN/08NAP2klWxUMC8acol18ZkrCohxEbVov5hFXIFLDb
MGzfObmp4FSuIP/FJVHfSzL1msbRtblivX4hJz4FZEPbOYNUOyaw5pu556uG
ScJ9CYth7HLoj/cjsP4qB95Yq5QOWwV/ycIIAwA/68nhaiREQkpN/6OEAA+4
dfWYFQNdWEIqiXQUppXsQpDLlLPpA7ulFdjb9JoCbHtlloEbvCEf0xeUDTkD
tEvT2/TB5K19wUyTTGc/9lBvvLAysmVE4swvf+tKQzqAp0XC+Bav6zcJ+9GG
L3pdpsNPxbTpYjubb3OSLAXGxI8aEs9DTdLjNf/UBhwMNE/G/4dNsojPlRWh
y031C1bRgrZWxox54hWrdtaRRhXzQIbG7n9l0vaR4TD5Q3Ra/aKeHd+ReMwz
5KGgIfxpKKD+zZVter8F9Nz36RgWoDP6ihB9DTlQ7EnvMCBchaHYSbrO3/eO
3o2Vfs00seWsZo5bz5sXH4Aqgcg09JR/cCPzNVCuoZ9i2cInsL5G6YDTuC9g
S0h7l5muDG7YPMSMkYH6PoSN9u1Qa83Y3F8xmZekfv7LM8pttS2YxWE3402a
GsW96Dw6G+pdO9YQ88nZb+AEqEEZOHoLUjSnUYsDTnktaHxasBRd4a98pM3w
62yHvhkXo4r3tsS7I0erNPzCj0SVq1P0+dUTc+lmb/TUkBAPho3kQgcegJPM
nLqmIlf/rfc3/J8PzHmRpuy+ebFNFI0L4ywnodRWLzOQ99M2OmKFrLK2Q4kT
UEtTvFVQxl6UfUOTs85LKl52xHLeKyWibpe6oEopWNPGfUyanh3nDUpir/SG
goJjSXTLPMqvWd6JE7jzS5u5Vu92wbVk+ZSGJasqAAcdyPPb37UPUeaKdmom
DIPgI4vX534U3ikobPztcAfDXymlj5yBxNDxS9HY+qcKFYUOTBVUuJGeblLG
8cfic6tbcnT/QjREJSsxbzM7/deXwoRZgZ4c1LijC6/KJx2oIWr78b01YFHu
5jK9HVKngvSa0Pxkp77C98htMoGFBpwXf+4ky6R+5F8xyvECjRku6REY889u
iZ3XuURSbLDDZO2tg1qPWsrSmd55m+xTABZRQoQeB7c+iDrJpN4fnn5ZPsoh
IgHHRkY4DiY8Vyy+SxWFBtP/LlemSppOJzBJ+ouRsh87rgUuA03EBkjSch3x
IyHwshcDPJflhYkHWmK82s7LroHAeHFIkZRDWweffboHcE71iYIovybKol36
Gic/ncbK+1iVMeLdx2sIljklDI+H9+ITDfxwZvNJ40yWjTfpUoLZpFEuM9zs
juyRltOVwS7r1kdpWE2CsZt7tbCXQbx2Q7Dsil2VrFpymfreSklwRXb9/hcT
H8MCWY/OGChhUGKf+Kk1iz2U0saFYb40SvzzrLb0HpHcoxk5PNr4tO8PTW42
LKSTxbgrSq9jXsToZCF32hTlexFNGbsArqg2jU09PT37B/SR/CccL+k5Ckte
tFFVA/Sf6tczzed2XU73O2oDQVY2+jU7OrmN3OzDM/X/n9gA9DnSMWO2LoYN
oyyV+ghCsIiOLo6JoDIH7kfnYp2+VbXjNSV+dGNu1YcmXo82Ksj0fWHIvGK4
m9bpOVt8c+QpSn+2T2zHfrrQESOVj554r4Q1mvdkprOJuG4kKlw30WLs8Ul1
D2d8v4E+347VZYj8C0l5w+xJ4WtCXZC5UyYAqaDn+vg8DjU3jV+BsBvryzvI
wfcS/lXIHkljkjisnTINNoI6duj2tZN1FXeW6H81K5pbjmgFGV6nK4SudOGK
JctDDEAiZpuof9LV5+08rD9If1EGI/i2DExraWMb7/e9y2qp+deStwOGYrIB
Tw3+/m9wtCgIP/7e4QJrGuOOueVfHkvQPuyFyVatraQgLr+daMsVgDhvkERz
Nvj2gixtw7BLvbhUNIW0Eag8Ge4U+3CmpeHqlzbKuzIRmuulrIsT1tJO2CGZ
k/L2MGyuh/1guXoKAEPxPR5g/FPg6+9Xavk3kb5v7UtaHLd3H6PMKeIeBgGW
pckha2g8BY+ixXxxbhJx6X7Y3qWepcFDh6W8ub6vxf+qm24dUyv9VQoLlqTJ
OU0cVg7t1miwl/W6NM3XRwSEm7ujKxeNq+Jy3y+YbjlEZP/YJ4mbwwQgL2zY
V/538atdugFcoIYy7ANpXPVzkjY9qNuwUidbB8ozjJ3M+df9fykuYNlbEgmW
Xn0SnIbGfMzPp/aW/+if0qTCTanzDBjve3ALEHeSJ+6m8IAOWBwcfzdjvE51
QN5U8NdIojB+KP+MM5r2fpDXEw/xVBMXVh3k1F8oB7MAHtELhLPrmGVMogx3
nhoi8657AAhz6wI90lgJrjo4NVq6eKC6HFqqaIGYJOGAGTUoVNgWwq9zXxF7
KPbxEfeqtA58ZeQPIk429WPPrfFlqTDEHjH0w8Im7d43tG8omhh2lu/EbNJ0
ZkHz7h9GEVHEyfHkcGHklOruni+I3NslhfudA4xqDIONYBYevSF/aewCZ9M6
OLia1/CtaFnlGTQ1elg431OAlZqCTqZ3fikqzoki/OMkKirPvC2VrXPTvn+g
toEvHyiZO59bdEio8anQWJUqjbz3HYMfvyiXDjFsvyQc66e0Zoz92UmF95dU
A4HNSvqkUmRylvQgwmIym1P2ED5eb/fwHHKE6oY8QEdvmbmwxYlX29GNrpG/
0rh+qn6ZByRArjtAUYseLDpk0Ft4xz6S9rCPDudTm3kNYo0tEo4BHdy7IXij
Alv3/J7LzIx4X4DIgK0MbEuw+hSI72BNOxIchA1xx3we7ozDGIRu4o3PPAxe
mUtHJ/AD4HZAFFNTFVKenOF3W4VqL39X2Nh6UsQSrZFdMSfZiFzRCvntHrY8
9wQZxSw0x8yTLgMEr/G1+lFWhpWjqMoumEix0jmmR8LqKn1MOi4kE8E5Y3uT
0iL5vTR43gm4fk+iRskqS7d6h4jKxbv7mEO7oj9SCPMotDZ99iRZS/PuAIBS
sZhJBVM8zjJr5vkaI6EpZ/MohdH3uAUdgEGbdPH32iAylt67+5qHb7o+OILh
5gfSGQRa1Soermd8kLcQzKTDc/uCzefcuIkjOmUnMp6bFlyjxElCsHHP2Sdf
Eov2x0pmDyZWlr4KB9R9AWjD64irZGvN8n4hU4z1EuUM3nM7ooPs/TU1RfL8
GOSyWAMQziQVVRDq7o2wrZ36CkbdzypOdCM4I5RKEe5BmfkaT6BlLFGZAd6X
QCSK1y5Dg3mk5B6bVx4n6fufKi40Ld/hDo8wFiSMk04vppnsuE7eOnYWhqAM
Y5Vtl33gFEuon5tUqI0QtUy15Ny/OQw9wGU/41muRA8nj1Bj+RDCn9gZcG+O
L9v34XSgLuxfccbKscm6VZ85ejRouINczhSyI8teFHl5sAfB0YFCLixp5agy
nOXyQVo+QiY6CRrlNNlLQdUrkIZ66Oc4rpNfBwKq0NN3hSrSD+sj2kX4eiVW
ieFCbdU00pOmgnWcsbfh/ncYoFVv3Lt8IkXXb8owTFLLxHioyVpHoMMrFHDH
E6WBEWc0+9kPr6FLcb1/2w7FpHtJmC8uNiyNfrYxzhxUmSib8L0RBv0bUWxq
CMKXmvqa5MlT0hGTuf5Gg0/JlmLgOhHavUe8lvRe5DVN2/dLX4ah/m2omoB0
0edtRqwV1Bdjw8FLXUvnLuXJ+KG9qDvHtrxzJYGQd/BqGoYDpw5M833o/oqq
MbJmnW53jmyYS34tz0gABJ69rnJ10vhiZznrNBlQF0cJ6DocpLttzKZG8mra
USdLiaDN79KNQ9FvGFxz5SFpYvpXExjNMFYavgaGTn9Irlij+uvIxk+47mKx
vldlCOun1zz7LvpVHCyq3TX5SN0CZKLvenOXgFE6rfC/U3RWvpzQFSTFl/nw
KR+JOOr6badgCh+XxfBpUEV7h7Twdt1fv/RpaiSdAjQLtNZNJ0CsmkOICvEk
ZLXmAcOgkNxISIdaHZGAJiVhFOAAzU6URg9oqpM877iAzxQQ1TMof19uM57B
Beui38WetDcYZ5Bv5iPBj4ZThxXyRth3D9XsRhAAGOxGY06x4vccQr/VlKOI
tk2ir3T+TqJlqtM2PiJpW564WLQM11Wh5GlcZ/YZ/ppFnbT20KNQw3M88u+l
sVdh7HikaH0KrlrivayDmLIQyHL7o8Q/Vpf273c9RUvFAmr9HsIThi+mBXQm
+TtQa1yWQAwv8Ow/urQLX6c/ot2ABcyfKaLsdbuecPNA/fS573OUS8cw1+Ag
hTwj0OTMFC9XbxSLtyrl3J7Uwp09gjw/M5GOYJgyO1sL5b5s7Fq4AUdI43Tj
q5uz7yW2S0Qhgksdt/VWYITYyXFYvWyR62coPrWX4k2WI+lC7Kfj6ddAhmhY
N7y+J5RdB1JMZkbkCK22MQMNG3E8rA1W2RKKk8qJe6eHKd1px6pWJvulIAX2
X0GrrATLYDULJVrwM9VTxvMraBme0gtL5kuu6+OKnaLXDPvblpnheHQQ3PBA
AsZrmATxybw8GQjhb0uOagDX79ra57kDSxRFHwLeCdIuap1K8Xa5oBTXp3Dy
gRk2IxUFb3NVJGI3UfMpCAdl1P5wFBDn+xq9NXQL/fnErrjDJqvMalSDS0+f
Agz5AUE4vexXxj2N6Xd36aKdV6u9kFcbw+/4yDi3g1ohjxqR42RVuqftNf2X
0HL2yq/noPQseT4FSoEUa93zZeCj2djmmSsN5om8Du8S6B7cErC2vj8dKt4c
Jx3XXJjAf0WZGH4iC/Am98884QeMv77PcdFnm7Kp6adonk8HNSHWnXaSEiPj
WUnqEh02xqu69pLFcPWYDegzq72M2sAUCVaUoA44Ksr3Tp798sfw41CScQa8
BrSuRxZWlwXhWAappic0SBBFvXLNuxQjLKtlJj2yoyBLfTrhrmbEcZSnyxo4
UrdKTJvBuXDGpBb/aYK/tDU9PxLY9Oi/9HyFGZ9eivYrFp/8JfPzRqm7A1oC
SrIQu4Ji9WE6aIEcPwspIzluYgqDxSgzKrLKqiINjwCpzDcB1rT7FFYnxAz1
Cmc2VfZylxSfSRjAVp2fkeTzQ9kSGKQQycMuuQg8bfiKsV5hptsHU0aUZmIW
gekXNaLSBr90yMMBZq30e3BlDaLqntz/XKelF/d+XJNLtPH7z5iMC+L/ztfM
xVyUKG3VvBAottnaCKq5nEJnwTztmHW82PF4k610x2wJms9ViX+cDSFeg1xC
dBtTknU+43MwP3AV3/ORquhB160GtH/9iyeaOIsJYEBQcT25vraL/FKuRAzS
kJMG93JBfm5KGrWN7Qc3uFU1aai8woN9/dMd73YmSNBmaeoGI4PnrraiS4LQ
pc3+kf8dqpc6mkqQDwjqnp1CQymZ+875NIGTr+XZM50b0y7X+si0TaBMMgzm
5Ugq7lLx6YzoaMS4im7ln7ZRhLJwR6YMNkrg6cw9Pfr0Zyj/AFZcXe82slK3
bUZG+7he8L6PJd2R5JAD0J9v7aOAX7RcFkeozLmisguiFK+1V7AuK7khKi3i
vTx9jhmEUMsMmhyC5eISlLTYQXnHFkTwakCqUxn8I2Ie3IfHtK2Gu8wVUb6m
QRwMWG4zxnWjBlobBON2GbjsRwG87vtoFgR26iA3r3kktTb3MXPrOUzfe/zy
Feu7K0NlULNQK90sbWAuPwDXyeGfNwvEdai4nVZbAhpNMHly1QPY1I1PWXrC
Pcwp7kQ1jamvsYNN/adJbgf7NBT+2gU1pUf3bcufGPbzBpWBZcZFQ9TPCZAy
PJcM3k2dfslgzXgfpgNjGMSOpwDoaR036VHlqasdGF9YDmQh7ZJQG6ELRjUG
P/jr7e74m6yV5b/p4VCS4E9MgCXOdZYNp0+ZzT+Duv+MFYYCk6YcWHB6Ke1+
l5zOwak5NdqFdS7PICPhiNmQIRu6GwbNqHrTmSTkWcDFVMQPS1iAqMuhi27K
1KyAsvDwwhGEJeHz8BI0UMx9zGWTn09dsxG5THEMBCELlNamhWZ4bbNGmFeH
0ChEXromVOQ5liWOLWbbBpxUXCBQ63qhGpr5vbV2DhUgMfOYIgnV1DbEqva4
UKS/UcJOnplc/1OoHZ1Tg+gCQVEQUmDzG30FbneIFL8Xsz15d9c82RZMeLaT
o0p5LwZrFZcZ4L9e5FlLGlKO/QeyJ120A3EABFoSy+i47kBGozeUM5L7H9g6
efA2vIS6se4lqg/Ttqgs8k620CgfxKXR7PPeN47AUQkQzAAFDVDvicCt3hGI
z2m5jzs5usxxbOH9l7wGmOh15vE9b4eRuWxsvgGdKYOTTKm4H1h2PtKTojY3
HTjS8/ghC47XSFloiu3PwtmwOBABH+v/Sa4AHx2SiuRUrVdsUZlOhFpBJJiK
jdwaZLBt0w6VlwXeKxsTdE1j1Wg8C4j6GDddlRQvPUkk1ViDUs6k45Vchffa
30Sg1XqnOCK/7CLDGY1Z6AuFiUJ7tBkDKFiC82dwl18y7MbTH/lYzyJWkWe3
6umv94Jv+XNkoaLuzd4WxzJshyWp07EJL/5mu1l0gL2sYUNQ+DjcNSMsm9K/
nrB0DSPIC1Bp4LBhOKSQA+uJtpAGQoMewMUotru+wBDfMoGDpdjeB10sZxN3
NxgkFYEk3Mkwe7lx/Hj//SbBTEpw7ajBWqQ6e5rSRVSqgL/Tc0WENweTgn5o
q/WEZ3V8PltDC4wrZ8DDrr1wDOVwNLsz5POL8jg9hRH+yYMpJVeh5yOFLU7W
NCSK1Fsndv12/ik48USapVVlB2kc4J9VvZgNpo8Up4zniw4uz31CivAyIQ0A
OMUKZDYcKxrBHEk/ylmoxYBU+ZypqTgLlmW6FYEhqYzEg/9AMYxjGtyXT8sj
+X6xI2SFIpyunRj5rd8lyweBtyWG6BHuRe+3YkNs5Zq5iGmTJ732OGyxztNi
FOmV8BfeM9P/3wVPBdk/+rk6UIOO4FnFcyhzKGiYoNCqTtkmBo+TjGW3FF61
D+ZuklU0UYYCSeGQQgEUTbuBlZJ+ikHgHWp0zOkqRx+hv6Zkkr3fZYkKBhAL
NSIkdAGR+9KIsUBxPjSpYkt8mSmoFIJ1JCrHcrGrykzaaEDwMutBfJiiEytP
SKk1GNqm0m6f0Cs5JCm0ghOw9heVnQuT3yXjP/pSHxiusr1Wd4Vb+0O+t6ut
o4kohVMEf830x+irk4AjXynOZcBr6nIwf0w9BoyV9Wgk9yWHWT2DAjCuAPSw
zHRfxufvN71bi9A0dn9LvpxpI/9Guy0yM4DDqo49uJybykoRSHgWYhe8XTvB
qMe7KqPsJ2zkbFksUJbtz/CI/LnL6nhdTWVaoosxObeM1yvXQglhESFU3MNM
liwoxsvqSeEQlOz0IW4aVsso4hDOmo2q8+4MmmO7HNm99Gg2EaI2Er9r6MOy
i06M5xW/kDAOfIQsKTTDcm+z08MjIpzFX45HpmGld2+bW8zXx7BM72UKdhkx
ZWHKjt7iIXRmPRZ82EiObR4GVN0tU82Ha7wUC6jBIoI//BxADP8LLOb2/hdL
yBxUzCdCUTH7wwxrVQrFnLBGHnwuWconMgToRF46J263oMhMqJzbKN3+dXQg
9DUVGRmEG8yQLD/qIXtqjzIgi5XJLkkDCcv9S6YVCIe+vohMGb2Fj3oVEEuJ
7+ubUXujx4m87QkfH+1Njvk6MOqJVAPMBh48UgyGG5rXO8470/znS5JPwK39
dlr2MZq+uhjPdXEMhk6mV+v64ozkO2HPILRZJYakha0p+uFVT4AT8ijXL+nh
YlV533AJcGBZJJODWuc1o5Vjvj3mx3lPf/GPeJvFsiEid4vvXu6z+0fUche+
o73KyPTGrSSyM3yQW5Dwr62L3WNE1PM0Df/LAZb3g7R+jotAckR/OxnE+5bZ
CVogaI4nu6+/bGJ/Pp8erthet6XQWCsZI5HlFUm2N7frcs25G4N+zYC05WzU
WGnEVPoBEws5zeiyOiNmQOrri+knkNEme5n5hZjQW+x4880tN/Trc69TcyMF
26nzedT+2BgLcF2wTRZKlKuZnUWRKQpmyCzlmy/2C6/htI06Dwk+Bo8wxBf1
qFRzs4M+h6UR/O9FEIt2+fcTadsGxRuSRO4p6Kas0js0GPnTSs15VTdCVoE9
n443Vph9cNGY8aO6rjwT6jwZ+Esqfg/LrOrUC3t5C61bCFMKYfcN2a+7ryHg
6BH9yAar6JJWoLZSFcfEEEsXEs6hs0Kyqx7ZTk/t8iVPmCRCyCMabullt6Pc
X9lhe7MNEcHn6rqJBhibmOFRhJWCWeZFwitZnIbQCzPF7V7LQ17KaUetapta
4dsqFZIwCPgyUjP+w3hK5lOal1pPnfYxHjatU+uE37ESaYdnxpw9yLXduiPv
7mgV8uBuyKPlm7BodzJRZEj8fi7Xsybnbb4XxReWyly40xkr+DcXqY5e/4Yj
iyifUDY0OYXbPDg6u+k6PmnhEAUTfWn6uTgj2PtXObEVNyOsvNbZGLhjrs2Y
ZJtyAXKL4ACXh4zNFyuW9tTBGdY+NlRL5WcDAdLU4rBTtOEllArMhMiSJ3c4
tWo85A8Hy3mCGJavbpKwdGcPXJYvoFARKKHUyAxmV1uL+9tVwbo3COMpgbs9
bOfzEeQ+J1TPCkTnxRDkJYou/KI/F2Nl1Vf0fT9B4EHqNuLlWg64BqpNjtfi
hztRAj6P5iqDjIFADbOlwWLEszvLoBid5TtSlmofkcvVaqEyoOk4BP39xYEr
BB3e6CkZUmqeMU9Z5K6N+QJJLnc9gVPty4k3fa2sDpNAob4Tvqs2TePHuNlG
zea98EzoYxx6vmpkg5vcIeq4Ecxcfwetjb2cpQGYNYgMfhXDeNZeQFMu2kwH
L9+pgWhEy7NksHpJWt1pV5s16G/4dfRyoHUbu2p9VqXcOnPXOJrvIzbsrkym
n1pnLLsPhzilirq3wv+/o8QULl28qEO1KwYGJ9EdLh1VH1mLQohkJdK9Yfie
zc8BqEby94FbdveckH0VzvkW2ucHu9P/3OSRzEjcjNYGT3azQMYlu7V676I0
rpSgNUzr28f+TJSpzOvSuYhQaO4rGhcJmkx0OZkJbBHIdMGA593YyTIB5Si6
yG6iGNiHoVc2nliUIOzT+SJSShAQ14F9XlWPhLmczifddrRLM8Kkgqj4QHCm
2MEX4cfVVaYFqg/w+ds4VDM4xdAMSIoe8+HlwMAaxjGAMvgwPkqS6eZsRtb0
KSqnIYHqitTshyio2SnrTiMzOzqmxz8qJJFag6HlbKuckjin16bK0VCRD93S
XIv6YsNABgU3AEofYr2oRsZgQw1X1VGI/GNp7XRgZVg4ej1C+kxI4ToI2dvg
6RNglNYW1FUoHRHlK/4Nv8vyrfd3bV0HSDuxhWO2ODnMJamJhEOuxZlWogiG
Jf9eSU/5CCM04a2r6nJx56FfvAojhB0jjFxHAs5Jgpo0xsBxJ5/0D/qoIQnG
8lmmS9uueHJ7sXxOVp/X9Pdee8nd76goBjNXpE4M8Zoar6SHJBu5gsdRm1wX
P3Oi0TpxBmyEmTEJ225JqogLwfmG2lm+LhOOrSdcvjwj3uBsy4XbVvrylMAb
PAl5Wf5j+wGRdaI0cN7H6HHa9KQZqeTSBPFd8Zeljmb1jPXTdGX/2JDbGOP1
kBk6LRemgX7VNLOfTam2IKFH097fUFvcrPW7PdJEw3dtDW0fTxc+gB6nTax1
QOtKAteCsHqRfpInyA/FyaN1ZeQ4kIw+B5tnEwX49XzZT2akeUGqKH8DtaZh
wBjRFcP1xJGll6ylhz3wsq5lTXv0kvW8jcPDkWC40KBc/Z9M4ywLE4ogUo9E
D8MlxpKNKoBrJISj4QEU+YXsFEZ/uJ6ryWcrDDQmn6pqOTntIst2KPiTeQ36
p/XnFfRTbihNma/1C2rC4jasAcaIY9SPETgGkhETpZz2qJJT4XK5j42P1l4I
2pxNlmeWTcs+aCGzfZ98NGIjtpP2ytaOh2QPqM/j1Lqmdt4nW//hrrVWzEEy
9VeY9M9tLCJMYN1gYeEaegfPlNPRWuXpMF/o6pDZcvsh+bvvEyRnA97lGOjo
yyUBW9l02u5uc1vkDb1sXVSljle0aOh9CzgAsURYQVKjcZgvZslRl+hCPuJK
J0E8dXy0ESxYcOT2WZ1ej8bR6VUjv1Oxi8pcVSMF1Mi4aC2QdZzET0cG/kwK
zpB0wyJuYLagUUeq87tvPJ3jwDWk78s/IFJAmB261rQds/LLGiqKCALE5X5g
oC9lVt91854kRQKB5AV/uSDfpy2uCA6uWOl/Jt+3MVd/OR4ORWFS2boERC+v
7Qj1sjFcjHUi+3SQ0dlHJ2I2o/oYfFuA4CEjlq0LIokE+fFBd4uyouhHZQgH
X+kjOnYF52BsjpbGvfJWVVUceTEHhiGtnhyfKukfYYBZlDOE/zzkXZhBRtGW
wjbz7Zwa0HuuRMdXyJEk4RRR1fW2A2zpMDT3sQNC72l0+K7s36hRc4mCGxBI
3VEYm7sHHn+6EjCzvvmIl39npFJyYe0HynV+3Am7Mf3FvhxpUU8/wBlvNL1K
PTZ2QHc+D3biGSrB8tE0u9HdDw+MA0xCTdUH3H7qzKmtuUc23fe29XenByQh
WR5M+qSXxkfnEtmeoa4poHDQ61uNAEe5opwNThOSzQjmH2y9FMOc+2/NiVRP
SbYGeH7i+9nIcSue63b2eXfVDffESAePoKQICDF2v26D6WiDNjfvM10Pmzy9
GCeZiBYTsfkEjgsXK/o4DgKWzW2e4p9eY159TXo2vNquVNHVOVKQDIsrlOQd
SNLGm4Hx7l3VmBIz1D8kHm/uZ2n6/Bxrx5ftKM6GEoR6gndmnEynEHbTsPPW
QiAwC9WQ39Eo7/ujXseITYW9eFjw70APRDqzbRxk9WWxbmbQqvzczEu0m5Er
uQoyO7CZ3hFdxOPeq8dpjqaMh3uMkLJUlcJBNjeqZozlwMxSslZdayvzIR6h
55ddoE6MZazw3EDK7r+B6TIz6GBEUKrYQzPiTzqL3nDBKvKosi7vkMXfu9xs
/3sUvVPaqKxqfQPIqFxsYWQ/8jeeQYd6jFXXKs75OHPmOwTo0wAAkxCVNxgd
KsdLfxJDxxDNku1FUNtbzlR9mJXfdtcdg02aKP0EEVeypYRGcW+t6EdiwgI7
Ym8U4uz96G8lhD2r7qlGATn2nih3egMJlQ+uhoo/DafaK8RBuAfcAJzwqbdU
PNxHMmR955dGDsmBphatcvpzO6PMLFrtw5DnL6g4r/J89JYLQK9MpeqYVdeg
CUA/053gggEVwOlvxO05w72V9zqAoneuYmxzdo8ikVtjEuIoINU0vHEUWspc
+dfIBBBAfF2+jbQzRZeOWEIabpPQBqi/dK9xLWCD7qsj5EhVjsWa/Pv9EeMW
AneiktBVTKUSrcbfbCUY+YRJIt+ByXWjLHzh71+YunrNl5RJBCRd28O4h6OY
aoawRHavZY6E4knjT50SYaNdvkxsDXKGbCcOjYBKSlHlJkYDtgZ07tu+/ym+
k3vuENtnHeuQCFWWAatgJ+D0tQuw0/+sGy/zWPj46bZRlSYN2H9rsoISeTDK
6QdWqAll20dvcUL9/5ySVxzDQJ267yl1RBPMULdzNARWhIxSIwlvZVPRW+Az
lN3+kwryOID0o0agKV1EsNviA0JTwR1/2bXR/ZbbgYuecWmj6EOBdgctA2Xy
xa4pRYQEs7USHA4jlJb9Zg/Yt0QzN00uCVb0x4KxX0C7m+AzkFCxkeli9w4D
b6L7UMbsKgEQpIG0WtgUWZtyVw9HjHwqAmA7YABaFlSlKL79uyFAQs2IJrD/
cxaD7gMq1N7HI+ppvEUs3k5BKofHEIF3eJ/8kzzqsEUvh/TJ/x8G7gkz0I4l
wzvdY/0F5uT7WS+SxfrJBjDqsEwQeUX11FmNkpBXbOyrskGjkLqqYmXE7vTJ
nHN7xyz4hr8Fm9OXkM56QTDd/Qx6jVdUmzxKMLF+yMVoaYvsyFrVwoEPDabk
TxlafQRofFq/3VcZQtQTCMsi4WfsZpsa5cbQ2BRjqpEOSuyZabR/2CwegM7M
aqsmRo8QCNeiE2QownL5c6LE/bQSg5QwbaoO/SSQw7IHuTwN6+6MI8yXF3WE
dseyTgotJnVwAGyqd2YInDH0uBGRQryDWIAfN2KNapz40y80KXXxY/phtJCU
f/2bn4E/Z1y81YQkainibfXD8toIeZaU6TqiqYZ5uhUjNz/v1G8LgpMTfiZ6
10L6DBJIj87VvSff2ip26VThY3ESMTptp/kiXq4qq+Qtarc4W4cwNPzYG3qs
Nw7O3la6VNcutb6M+zfaCsuMQlKvVwiMKSLAwdU341CVhPsgk3wRH18ZXuJE
LFaMYvY8N6VBgzFkyyI5j6akjlx+8dvVtRnj4ISgU9k80dcBxYTZo3HneIzG
3uX2pT+hsKiOO3EqIiU/mQEpsQRkrOvjjbdyARxiOpvSt5jV4Awcie6spS0s
xslbU4eB+kzbGd3h+vg015+IqJvSIF/qDnQLQ4y9Q9/kGaJSjAh89WSfTHQ6
Wr16VgeG6M4XrGmssuW2o0MybAgg3PdCKoexpEB4xsfNOPKipn/x6XlVbXnT
kEXg7Hxqhzswm8UCN7jd0OjEpq6D8U6NELVhHXF1saKGkJMz4pXgdcZakMT7
UAXGenUM6aWOi105/AzqtAn7V5olDgzlP7w4iupZWVatTimr7IMOrE8GeUN1
SDJkl9of6m5Ois/BAzhHNfaP82KZKwXNameqfbksl3U519XuDKbYgdbRsjWu
OZCCmQu6tttgpdvSb4MoFr3vESwf97MByMX6+JgsU1NneC9KaAq7i/xFFO8v
IFJ7RnBmu1hlvhq+OD8E6zrqyOL/i6PPtBGMv2RHdAHAc+hymhbjQKpBOvYG
Lem3o3yD3jATAsoiHv5LlNZuZtuaJTrlcomxLEKtZazaHJmdUkhtLGRnezUZ
Izmu7QKq2r381ktQiV02VYIbYnZ7asDHegX9OdfYoAKDGaaW1qLmpLkfN00z
oeeejUy+HqQDUOY2/UlV5CsilVCCR19sXWo3edXQ+MKfEz14l06l/3c3cBq2
X0KsgFAMncGRJIxcfv8jPEDT5H65FDXu1AJxKzqVE3swcu6JpWJ+lb6ulzsA
39iFjKn0kVoiRHr191c43OZWgY84XNHzpInhaLBX5qZUvrWa0QEC3oe3NDdM
LaCEcmaEJbkre8nlI/lkwHafd0gHFeec+c5/v+uNG61zc94paRD2Ik0X4E2L
4fjZE8iyQU7xbCAbpYzSaJulOGlkGvMye9cHkeg2EI/PBJg7JF8XwoGIG4mF
iVaskDFEKtfio9Jn6VXLu9qAk0VWyJE0E5TDvSAaS+QIcxmVEnaN4Q5OUPVS
cm9ca0AU0FE1Ezklh44egAtj1tNHLLPPnFzsy6OF+OgEi3zdxuJdCTsZCF+T
s+P0kPNEo0QmISLFjGmt52gfgYY+2RLcjjDJpMaW6BQDO5XkTjEA4vEXb6YC
D7xKMrCPe/S3x+LCnvsC4X8VuqSx+3PaK8LOl/DvPQI/+7hv5HDt/VGVw06C
XLwKxe40ck8NEKgqhzp+gXlkUjqRxkZRgy2Zuc/R8PBZ72LckPGm8BrP+RD4
h0MNNt8JZ7M3xkMaBTu7BoE5QwCH2O5zB7u72RFMb0u4VbYfa6x5IAgQvaoB
DG0+CMYHP15xGXDzUkMgXkuVDtlPJognlTWtHm953k/HRTutszMqLTmBoJWA
uF9oTBfSTJnrxNK3sjMHjJOmL8mOCaGAMH/Bay/5Mbo6ZXAOIICc3lSfXWmX
r5Z2D8sbCxEroRUjgXiXAXFPGX/Yro99EKRYL5SOFHyP8wX8K0KphizE6Y3F
YKaIZbEqWQolGqEd/9X1G/aj1lCa+q89kI4rxvd+VvnlmHX3FU+DnyjQwwMs
7jyIVFRyRCs5Ai51mhbQPpZX5My/nZbJ4hbkGmEF8ddAWEGk0yFYA+cqa/ta
SGTYHN7xnvs7HLhRLLYvyBoKDXfXovvF+4k+gnviGISMmyebv98EeByXrj+y
ESje7E5X4yXR8j6d1zFTDqGQPUqFxDABROewWr6V8Q6ylimpywxdvCwAm/Pv
HJORTijZcgRqkdgUndhY7pC+pdgYD1s7c+aGkC3Jb+jMElOJqM3Qogdea5P+
ekd+CrfxbRDe3p6/b/1VREMPdiQM3YKjHCcpxdBt24JDAIHWYiAewYqk7B4o
d4yWCEgBOx+k8o4jS7spRB32njnP//kYETvLTkWuxsJUvJuIjkdYXqYfspu6
IEf7dxA6ZZocU+q/QlAbdm5eVFfnvOFiTO1fpnC3T0IN6gKJiOwSDYXxbSqU
7GldnMOBEWPISJwDYMeg3+fobyHCs5zAxSiLIFa8zwI4EyHfs1Cj/W2lz5ab
Ka2b7bD7LDjdD25W16hYFBSVwzJBKbVIYS4y0VkwN4KsqDMHjbFEI0kO9+Ok
/yDySsORBcuG/xCXpyqh

`pragma protect end_protected
