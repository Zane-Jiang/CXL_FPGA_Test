// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q4Zpq1mWdHMULRpCiHOQ/pUmcWCUteevn3W9fqSt928ri8LCuPAs8LIaEfUh
4dNdIvM9HgRFJgFmG+Ll1U9RlNZab/Dl4PHYSXyxioucdAD0Ecgy703SL+li
d/DziGh6JQFeFTqsE2bU4QODhgJkRfovk8Eya4rGSoVmjBjySr6GfijvkuVZ
fmvNMKbSl7LCzhTzSNy1gHoFXpHPw+SkOS0jFAAWZLi9Ugg080jWWLbw3V/H
vn+j+map/lX9TV9KmJ86LMRSMr2q9IaojOzC2CFxn4AaM46nDX4iU6L+ecp6
Vvm1NHEtnl1hfCZJC90Z92kudYchGBrY9RPQxZkSWw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kfpU6ZDtCk2XldTqNoGNIBmFNXHTocI1vh4dHD0MXVSGteNZvvm58sAHATiz
wrG8LteVexaF7Os4Fd0nawo8MUFROifCprBSno/h81+UW/V4DIdDlb92OcOu
0096v5/AxkeQ5LN58O35QpLlbDIbMYEm1lfL2X1Vg9zZMHXDuP+rQQgotrCr
1iENz6se+nmO0Q194fdVhbcPAUNLvKxyiK+oIO4LjogHwrpk/HxVogQtvcVj
spMpC5IYkrgQqJB4NCPkTLV47fMkqzhJKB1fC5EYrgkS/PyTwbMh1S5mWVP9
rdBt0M22svEr0hIjI8cXi7IKksdWTSP4pAhxNiKOiw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pAV0T7b7mTtqeWT8+Nlk39UJqbOK1HZt8IMansBS8EjZf0J7GakJeFh8DiLe
wV6/ibVRu6o/qVWH2egAWt2UkklxOlvwYg47r+fM7/L5kH6uOjhsjdITGzfQ
g9oLFdJ89zJSPhB162f0u+u4QtJ0helf9ApaogqgF8eziKPS/mdJclAlmWBe
16B8v1HoPYn2FwQnwbChI8AXJhiyTwP1FVvly5jkA9qfQo54dNqlGyD5UlbZ
xZ0gURzb7IZoiOid8oFgYD//71OdCXP5rRZb0PbNWFlsmtBUz/7OQT3wyHbK
78nQemHPjepI2kXr8TOnLt/xqEuwwQRhUet6fJzRTg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VbRNzZ2nAR5omwcAn5bn2Iidm/ltRB8nhnSJe6F1whDp02V3tcpR8vhT9RWc
JuJPgjoYNLQwQ0DI+X/YywhoHISgjgbX7WfyauNRuA9eIQLviW6hU463jvFe
HPDeXiNZRp6+gaBIg5KRcsuNr8MneK64QbrX9pDuJJymPXEauQQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wPv/oTWdUslhSR5g71F06l9oAQSih4cA97JcFP+Jrx/q4biBpg9OkPUZh46+
lpCWTDI8Ic+pvXYsrBOBqHxCg6lHq9CKtdSEvzNBvlvIHY2n1wDe8JtH/XwA
QfHXZ4wSFOoewFLAdZcqGoOQsyfA7CjM54ePB18L4+xuOZoeve2/FDZ+OKrl
vyWHXVNtZBjthhg/Dys7wtE4r0TU+yoKMTaw8GIJvaRd/7T5EIeRTJ1ZN/sW
DJPw4+qMalCRe3jQVP6caWDIzK8YUDnaQ1GYA4cCmtC3oyHzoPwcSMi5lIwm
e1AxpQHhmy6f3HE4F7E8+BkBqoD6cQv99lrjYX2XZQVuPS4LQ9fu9zswNKUj
+v31XNu/0YpUtJgZBR6RMSS5i0ABFtPmPCU30Puzus30lvg+XhO0bA/3mr4e
z6y62QA98X7iYCafrbUv5N5WeRTJ+yad4Sqv9Al72xrsUBcsT80/HjaVj0Ge
52I51mE2c8EZveuO7oC/zpgE1Slnmi4c


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RzCA3jpJA0v58bJu5UeBoaw/naNaTfhbGSt/wnORG3mGOMDlcvayD0z1E2W9
klyWYHezfaVmTKPIr+NLzveY2mN56OBnNYk5B1dt+/Uf/r/IeccmGFv6mH0d
u/TRW9jpS7Ez1Svh4GecKotkd5j/TOqibaxZqB74sR4ge6lExvo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ha8zS/QnGK9jnBTXAQqgtgyjxNIU3Km/TqYzryRmCOVOvhBOAvrsGFQj9Sk8
2tyN1kwoor6dflRpZAFD5JUfbGDj1JTXYMYsE6UNilpzYub16nW8dVZYrZzh
WjpNaGDj/IFx5ffA6XB1FfMynK5dpXkvSOcLEf3AuOuxID8/6xQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 466560)
`pragma protect data_block
nmq/3iQA7Rw8jIXR/N1vviMovhpRRogkq8pnbMJ+zV1/cEbNOar13CCOJOih
03jnUJ4UzKeVmapkP2wQq1c/DkYBDoD/BpuJ46UKzQkrDyV43+SUyzO7XZQc
341fviSTyhxEEfvbB66aXSvIlsHLlHFAENd1ahhPrJSeinGr8+PqiX5/4Sfy
PCBwwkpsLJwtufyE4S5aEucHTCjLw4wpZ/jiUXz1yJea5tvKeDMy2tRhbJxI
3puwSh3+PUqYabpBvmsJUAR2ZiKLXOh7tRenQ5FWoTClcx+QnAgDZuOKYEG4
z25iZHD81jVBy9ULQsPDFI0G9NtsuXP5rhe+p8pDa+h8NTeeL3Vi/0On7Bxf
lk+R1+puI3CQuBcvr8HPOBs1tcRa1PDquHi1EqyG1qS8YEYzFROyCI6CJTjE
V8ZUKOMQaa0WkZ37JenD4YbPslfeq7iunMXmI1gOcxTOQPmYqfeXWTlutmeB
scdctLxqTdCWdbA54Ru4sp/c00uHHv3ZNxhkD/XPrSzsD9w2svOX+EMX+fJE
1jOcCiFDyXHEHm+u/VrhjfeVNftDRSRdj+rrm4ZdKpTJTfDECiHaXgPL/A34
MTm63SCs5XDGrskpLAHItcwtNGBCkGl9UtiBujuhk8rKbHU+5U64nI/Tr35N
vF3F2n27p91NIZ0XBjRnhDhlPBlJzMzgtlJw1AqeEqVHrHLl9Mc4Ph79Q3dN
qRJ/lm07x1JbMg70aky1gpULKCQKOxva+T8p3f5ISy8szVrOJlvKAyDeNoj3
fjBGk1SdaF48bOROijZoO13wcO83x4m2EA3YQ9sqn5B/YrhajzGWko81ZZzY
Ut8sUD0BsHjE7rqNK7igSRODzdR1o6JioUGludswLWm9E9ZSq7rLB61w8ZsF
titDbmnXzbHPyjDnVF6NO3H2w6lh9FNJl2kJyOP5p5/bPm4zn12TEYrSx7nv
RDogn+LpoFAu5H+Otu9iltC0xOJ+5NdH8F9r70WG41TWccxHMbOv04350LV/
rVa5h6rtdaqXUb6BaTv8lHz6MYcR5frpoOnTIZDDa+GZNPxAFKamgNEzEXR4
i6P/9dOj0ObtTl/CGGH2BTsvd7kr1+2PrgO6U1defLY40Hm6w1hPM4vJvUMl
E4L4JKFTM8QKDiKZUc7y9BZFDN2Ym530c8s4xXYoaGP4D1+XkIBPLVsVuSq5
a9Qi3A4EXXqX5ebO++Aj1y9Fg1IlYAiowOF/64m70lZdITA1J8NR2PQMSim5
1eE1CTAAwOyPAX+N51d97i0hZu22wINVCSkMtmMcBofLycXqKhZuxJ20S9+t
no6T4JKZHPYMphUvINBNuOzRshwUYv8j+kdtFDhA5TESc6+nfpzq/g0Oqc0Z
p14UILC2p6mtZxuhEu82lhRAgGD3X6QD/6KXuySPHtaO4AiWlWHxgYUHQ4X1
T9QS3HTAJx8q0N7qtRO4cpGPqkwJqY0XWMv1bKjt6JxRf/2vSfuLzMiuenUX
psgY37wmmB568koJez0Hj+Gb9xV8lCxdjYi3LJ6ANy+MpOP97Ixhh+l+5CeV
dSkH0sehU4svIZwwRZX+yXbsjikIG8M6zZpfE01bDOSkbtnVjaEmoINVcZJT
XBT7Pl8c1+elrq0OLWJznIkFJIAv9QHgBR9Tz+elL+MWvPevwgyGf9mPFp8q
sg6TM4wJ7Ong9p3GZ7tcDI2oiVPStddrhfR8QR8lqVXAWAOH022bDq2I7j4n
UYycSHY+lj3qGdfrF2ZcdnRdA8Xn94y/HzFeAasABOeUFpax4qiuZjgjNtI9
nEe+IsHJf198CPs+aSYcq8j3PQSLbmbbUqigA7w64vxIzApXZ2LyCm1L3zOo
C1yOv0Ot0C/dEyD0jrq7LlKf12y/wZWRKRlgL1RIzdlvIsgi2Rxn2cHBXWMG
e9ztzcTnmdGU8Of4bLkCXAkq38N+jAryvgXyxUw5DNuTHPSCnTbHPbQ4HtYb
6PjejzsXijHkIUGx9fYYOM1Lmnxn2M/6MSD7mzLU+e7aTTsjyHsEi+NS3xpM
ToIYZbMN/xU/BoZaKzrW7v+TpL3eYCPT9RMQh7VN1bIcIUnJlilrIAtKaoSN
craVtDOvA1B7FSKXANqQ3lTkpmVPrNYRsr6bY6GVhA6POF3CsHDBABQqdjI9
5/7eOBfp6tn9p8Dccykg0k1pkd50dglIYsG2NOgdszxryr6NflwlR61tVppZ
W+TvWORS4tsQEpZugAKuOzP0cx6FmGi4Itb4UxEIXXgYAh7PnKpIe6tv6ZJj
6R5XsV76oeb030G7VXu+3y/BjpAItOg3nrmUkDBuOR8VEO/oW+hTNklZieJJ
fbVkq3yns4X9Dzp44lQvYIYkxse9heU+OIVoXsTntswy7IhG+jYLfOrFP1fk
q7ySt2UhYO9ucnXIYqhFqaCIRuu424pa7JEL9PpUz1kJVHEzD3rZnRgWRFs5
e1duikor+hkRxGceQhcSSYmrOzKmL8fpp63nAIA0Il4WT19PBBbmNV+syfxw
HC5NTQ977d+IcWdlNQyR/Bbx4TqbemroNMGBtx8X97EYlj7Ojqpqs/6UAH3w
fudDk4lBfJc6wh6Cwh447m/tre/XHhWdK1uIOL4KNIWc1BIVqeyN7xWwSETQ
VKQtKs+z9XEqCEFVHx2WYcySAhFwyR9tx5ZQdvn63lCyQdj5+iAzp5nWNgGJ
zDNzV2hlS9KRt5R079x9l8AfSsSnu+E8x8Mal8emO7LAVTyOOr4+opNo2oxb
JGrRqPwR/zbTcZdElsSCblrTe479/lZJK2WQUCtskZG220dBihhG2RTv4bSG
MIPbm6ad1gBfWBuTTHVGA8uy9f/alXWjt238+2bX/NUV62eQVCh56+nkj3uq
ec0W+jYCkyoXaJpFV2lx+kgKP/RCmu+ztNkc2h15AUVAu58Z6Y/hC23Xwx7g
+x2K+xAmCy8lvU4zgKpVH5Ngqi9hknOj6EjYKW274kx4w4x03zS18ad3aZ80
yp7N2GK7PpEsePdvzPe/N2RPG92bHy3tfcpWLI/c0tvcE0etQypaK4uC23VY
7hDNOLX+qKz9BBmwFf/6kK740o5ZNUsw1fEjWmqrD7p4NsoJ0sxs8mrAXn8f
NdxpUYeVjPr5T5TFZ2RU58VHkpn3Z6udDyZpvmGd3Oc2bMWp9HueiG92jWi2
Qtm5vZo/fTuF2EqSctvSnZZQaWPMPL3iWuEQV+CrSqzw8MlNYjAnTpwssoOo
AUKyxSHQDqMpKJMSdEay+SV9KgEWujk7kMv65IrHabrAL8lRY6ElpS0olBxp
aJMscnDbtBC4Bqn7IA0x/wQz7kw5AYoc2a5+J4PhjUHnscgS7eH3KgasS7+W
rm2HWbJi1IkdYi1RvQm8Gs0WUIyzDnXESCWkTvjSgdgmuh2UntsVwl3o0SGx
u1gyw6rMzQxYqD0Y57bE4YHaamW0ltbeVuHXHSbxcGM08OCbrUvxoZIB1K58
q+/VaE+CDam9WV9v3fDZsIqcafxPo7xHo3He/ovPajhjkW5LUNu9zMOoDmxR
ozKoip+LTD0XQ3WyMgoLZxWedPcd80jfJ2TJSxy+3RLzPpdvto90QiIm2C6r
HQc0HkcC36CAfaMNfMOJ2dD/1kuRHZDYTzwVnAH3F4LxBDyK/qgoIdcYvJTt
OBZrRusvgCb21kz9FEeSlPMyJ+M4R70REN+cKs470wZ3KUgEpN90dnoFtH9k
cI0N+KAczUlLsXSo7lFN8bDz37d0SYaRGPb6d1uBM7JpNSYjrzf8ETzQrzvF
ohNU6bL5+GDm26tqA/Xzq60qpU0UXNpUk9zD8tC9MXIUDU1R2c3HELZpMxgv
XlXho1IUuDU/qNPEQHH/UsNEj9p7ha++1e+KJt6g1lvDU0cEtUv04Fa8azxz
qvT/Mxe9c3/Fka1Gjb1YDuV34zlpTkr7ds+LBKe0imgFdd3bdfFYX7KaO4yO
yXJslKFfz87wxuVqjiioPXdMLaTeLwTJUSIEnkrkop+fLnknrzs3MkimAm7c
TNOT3go3Cp21sXYEe80tohtnR/d5sJiwW/eFlv1HGcU8zLwSDu/3sx1ANJCN
5pJSTVbMAebBXXYgrMXYB+4ysRDcAwiDqZaTWmR9XfhbBpo+KogQXe+mb7aQ
0DKwx+uVaDIoLaeBSmJNKM6mklhR7uAuPFYt5WnJ7aMAGbRCKVcXjkRXA8+V
uWhvwa9u+xijmm01dZlAA+K0Ez5sBmCOlM8ewy/u/hCmhrnh940jv1j2WcUk
yVvy5DX7zOOXkA/Hjw9iKu3U6l2gnZYr+gzrZ58hHN5iSJdVbKkF/qxz6uNq
AszC8UQuU5j1dGqc4ndv+KeZCZp3l7oReSthID8Chf36jzZ6icK6uFDyUJvI
sLLgza9bcI7KV1XymusREc/aQMgS26U56aBjy9SpBdxQjGTYUKlZsfHSY7E9
0NDBnpKy58b3TWSF2C3yGx7+5i8iMI5T3LsI93u1/e0U1uLSMFW0yybKkatY
cYM4zhY9sTQq1Gi//GXZC2srVtIU/B8FUTJSe2/Yr7n7BDqHK756Im0OPkCH
z0tsmXXxQ774Kp/b+VJ/wiPYEtJ9EWUdfvcr8Jhka5WLiL/FQE2k16bmfW+K
6tlUq/vKwsW0EDKAT63GvyMG1OKq7LIX8bao2wIBNBQkgmci17Say2j3Ekfv
WS3D5XDHWknIZX4sIb7jolwGmKohp+uM91giHbEEQG5hSOp77Y3NmHbgEXeB
OQiLb0KtmdJzp56YkUbf5WsefAorlApIAT4VrQwSREoXHqY2bjeLqHlussb8
wfpVcM5WgTxX6Y560oAsy7wwr/5wUgCJJDmYBSyDKfpl5ZlWCghUezod03Hm
leKEo5ai9MtX5uUf8fy8OFT9dFQwZKo47dZxdGV2SGIWzPOrLQ6F9/kWvhLQ
FiFj5aeHMVuAFsQg6qimeRFJ3eyuZNieAUKeDgiOf90FM0vbW8Ues3jRqv7w
VB1CboMlMmQpRRVtnsxPE/g7RcY+J3lMzLq1fEjY3RkkAp1/RBVBc7m1eC+I
mesbGkQ7TuIpsdnljxqYv+H8LE0/WaB6ncoTPmdYO+d2L72jC3Ln6FFInlgV
NvYcWVZT/e6vouO89wkFlS73W+Nq6y50cuMLLM6WHOMgxd8IobTu2MmJiaer
mb9gaLQQedJV/xc+QXrqIer+fjuc2Sngwj/ZhBIuekn0WEjcLjGO4n31PQMh
me1+UZnHMomdF9EJP25sBGXREheYEO0Ce72mJzWIzWq1uDL6E2x8E8bRvESx
M2Zg1b0ycqw3tk0SiO5300zwsa9hQ//0ZGVmhyZGrmp8fYYaDQ0n0VRucSqm
wU/X+ueZEv5pqH5+iRBVZoxGar7JMFBTciIrT25mikWHKLQ+UjIBEGcs90un
7w/V6V684F/RCWffUs+/PFW3yLfx+c61Awpt0oivuJ3tQ/YbrwKar49rJ560
/YEBRrrcGCuzQs/VUowduDlWlQIxnll2hT2y7en5GWPjxBuW9vYgrpyhWkgb
BfkULHz9IqsR1gLn1KGQIJ81jLa4uI+nvvERWAHLDWmchRyjz7fc1ItgJ+TE
7Hf2Mfio8/FC7dvpggHiMjcKeGIJv0FpvjHP1bySl/ZijgqM70+LSx0wpW0L
18mh7od7xMx1zd4KDyMkd8+AQqz810sIvzxp0PEQIILx0nBJPfo3qz+rUcPu
CDjnWvmMpIaJwwTIzzH0Js4xcQCENCiirZmnwlRzoVJNIack8V9zUDtc015r
AxWfK6uPyr/9MN7AH6oKItdzmc4gT09IRk/WNkBXtrvYEN6rOihKCgbUFvtw
FCPvZT0zjht/q0pHWxKL4+5NBqEZGfZOvu2RIT0T0LmO/WdNo0T4NEqZYJn2
Jyv/DDvu06/JnsAHEDNwS3aJ/istJOXz8oZbG47CsLYLozmn1s7XLe28V4d2
VnO5fC4vjYA4sVlyTpGAmH0hXcUiZ7wtjYSuRrxaVziWh6qjhd4RHOI2/w6+
utqq/GHEktRMZ0x/Y1CiK7PsEgNERRBxM/0Y7Y50ewIFGX9jMbjhzsI05Bnc
bowyQ8XG2gL5PuRMjO5mtfMGRlfCnZ+3JWxFgx0DBk2q3EXwkaFcf4INlxG0
1m13cHS1+lyGJVtTUecQa+eY1VGzSJ2EtMleA2gkkqO21bF3SFZPJQ3laMul
4afLj2aanHv/1FEMZon2DnqkGIj8EXG2VKv0UJKb0JAgOIfb9Jyzb+F80O0C
Bv1BXuEMXxf+9ZScyfMkLE+LOr8DUQontn1o/jmijYs/ZmXIZrgJgcY7oZga
JTYtIOV/ad5cAowG1zaj/USB0Wvtfet1hASxGtixyj4HjxOw/OaNS7B3Jage
0zlNqnC2YHErX6EzVaKTPECVvLTAEpzt35TYgQkJebb0oca1X7WydFpkEDcz
8yfUOvK8X1hujvrx0iPmzUEIrQ6k6S2npfJXxFOFGwm/SgSFsF3Yc5rq1uqG
Leo3alXhdc6j5JH+bhiYJwus0CPEOAgScnG3gtQN5byWr3GdAgFn+bsJMmHF
A5WNlUlGfcZ4gOiI3dXl6ws/n4np+a9IVgRPUnGNMMHdZ4PsB2fsbMMhrEFE
13zlEctaTT1S/9LVWxc2LU4FUPHwWArlX9RIuZLv+u87tRv5R2y/o81ODojS
LyZtNY8nSiuuTdBf6itR+9rfX0RMH3VxilzZxbOJKA0vcLRSZwVb25jlhweW
y+qj3OzEDQaFUhaNEPXvSfGaTMvPn9DxH0RGihyac4VLVW1xfiJIv36dN2CI
L+yexmCHjs+Bi2VuoT39KWtqTL9Dl/bo86fPqQLN3J2tExln7zPYmdJB0Uo6
hpewhLoCIjCwg4UrowQg0VA6iKqhFc33/++fMWtdWJbTZKVwdZX5NV8s25jT
cUXa2jMfX4CEfsSPxELu6QTdTIAPYNDP7sGmTFmqSsP5UQouZKUVX7gd7YHU
HkN9EiTO4kCoi4UNXDh0p+zKkBOqDfUHqTAmMraSmoDMuB5RN0d8/A0HLV+g
h0pj0P47JcIW4kwX7ijmcjZ8ODy3+MDqj2i6VUgI6Ca+lWqDd4n+sAfaPVs5
vDlptqm8OVDMB+SoSn/uL2hmhOIYAIcu8n1lRBN0jIQPRxv20d1G6ThHTp3s
BzRtyfeQcz5oGmxWpbdIeR3CKNEFW87w6xSRJEBU76SYLr/PE6ECy3EbYFfg
LSCuJ8S/UH7YmlB4GfTtO0Rz7rCdTRSQCoohTs6lM/YW1ID+oVxP/B36VKJ8
kjO2PZ2rHk7R3FNoklC37pC8C8DRLhQGELmUYXmO05ClLsnqefi15LpP1/AV
YsQPUYMr3d2QM8rubZoK2PXSRjvsPAoZ1nkocvMVwUcthdUd92w6Oo/3QH19
B0DqJu9aoqoNX5+Z7rqUjm2rRE4qB3uAqh90sdMZY5qZl8C3sy9jIztr5RLz
fTbPfUZ1YEgR7fq094DM+lt8J2bLBuvtdhXh9MXHYVPOIZ/3tHRpsrIjUJ7N
qPRAC+XKm1AotHyGlck0R6DLh8ytxypISJks9BMTirCTxM5bYO0bAuVZEzAW
u4R0GWqDr3vAEdsmPSCnNEL23DPgTTNpVczOhWNwqsxcMD0HbunOZcYlnD+f
yf9YrTxfLHjgk5vqrVNHUjpaMMCp+RCCxGRK7aS/Em+/rToIu0ofEntbd/3H
QV69YF4v5qPR/olHDvhF/XJ/55DI9VR615SetoF5AqwFs4b6EveH/440FeJe
v8+GKzcGkgN0yvDgtZ2qgF/4Xnt22hJY9sEsAKvQz/atGcDquJdkdge20uP6
zJvm0ZM6hgXJtHSZeK5onsxL6+j/dSLXRC1NcfopvkX0QptqC/GtEMC0QdVI
3W4Pg5KAPLT2nN8qjvBj/jBBzlDbh0Yh2NfX4xK5t8fM2QnXpxFCDDFHZwmr
COHc4fYygkKUxZBGX+FRbHRSF8O8QtbKk0lWo4p3H14Jh/UxAbIMXSXk7a6G
PTV2yG2h+Tb19chpmy1EZHLzAflqYe59rD8KJw0YyEYfSYsfRTJOpJttvYP+
vQfTMS7ohZaEw67hHnrEK5yHrqQoN5BcPxnSCOipGFSlKDOE5CzfMXSN750V
8EaoA9nPJzwdy4c/dLPKaOYM92urJFmnc+613rwmwBg903Vepo5Az1dcNrsH
Ya+VByeQlMxVI8yJCOHUw+ioFPPKtU+AD1BwNm/M6tVziSjTp1pTv0wF+uyp
RNaVUwYCvYQIWFybNXnLl2zmbXZaqdwyIrL/93zK8im6Z4iXaMqx5A4OE0+v
Ls5moswhXyod9Gtjsax9ILy4Yk5zakC50BM+aWC4BpJGyRYT2wnQJb+KMZ53
guThaQPQwSawYHWgLZe7Y7QfNGqwpUXpYB1Ie8dvyYIR9bUOL3baugUmzQR4
IslQf/cu3NbIb1qx1tCitPMH6HgmqNYEat5B19MjDf5LsxfJC6ll+2+dhE6h
NitE2h/dKZzDYuVoserskWaES8xpcW+dePN76Ho3Iw8lDR5VjdVgImMUwA7b
u4gKEvMfTjy+/JD/DjA0dafEI0NTXe2DtqGhM1fnXm6d/CySoM2fQh2HlFbp
qN4IS/Oz6k001JeROmO2/Vtp9MQAA76C839elJUpIFIMESQw/DChPekt1AsX
+zExKjSfzWy97kEHtcOVMEt6GWDlOYTO6vKsUaWath+jW5IEdMvSiW6hZf2V
004g33WNz16iQVpMHwm9gARysRy7b7lYbOYR67JCvZQP7YRJd4NEMqFVBoz3
hRA51nuApAWzzB1F3ICTz7phYLZ1hdpEwNwYm+oFnWRSNbuNEcb5phvkSgQW
8/HTOr3M36tRnD5zxNvTCHaBCZNAHRPww9C/zvaIEeGINgoTQ9vShatVysdx
+ODTdX7aVn8bFIeIknw9npXMK4I7KzjhraA+oGt7aSHNg0lqG0WI74X/SZUB
JE09FB4wQR2hvpkdbys8ySRA8AXQJ/RMSV5irM7tB0AKSKED7WC0mH67mJOs
CRNwgt4tWFC+gJZlk9D+qPsFqrbhNwsCADfbiYP+yf2GyA3CslsKm4Hi0I7Z
hi1e1dcnJkFjekFEeZBtQ4tdefs88KozEfrNqnOTNTaGdoOPRtI50uo3KlUW
2RfiD+Tf9hqyBdCLZtm4cAyBfAXNqavC8rvJlf1/we+8j/SxLVz33LphqO3z
qQ/LGRK1w4zeYyKZDrIHqvXWNgWsFeWFnIAsSSvmdBvbLgaXoZcmvO+I6GCx
hrtBdacxvYnqW4ReagSyZCJKOj0xyXM6aShK3lXdyg+2Mb7FCRZYorznS/Hs
BN2OSJ3BSWhxf+keSp5o8E9HR6jgZ5HWvI0bcKrMvZEnej9TdodafBWQt5PQ
IundDyNkbcdANSSpfUOmcUiQ8WEpyL7ZrMgaLcviqGOOa6chdjAavTlLiV7b
gIVY61/kTcm5luZtJAY+PE+qb84heu4phdIyj0qOK6WuDScxknaPoKlTIkhb
ZOh7U9pHLfK6vYUhOgWVtuEQZrBoWq5H+Mwd/UbCU+GFJ9DgZOX2yiC8gsls
OQJldYkbh+97lPC9fS8ktonFycahLcyDDF3iBzeB4CX5SeogGMf3YOnlCdgk
mYJ7ZLzJSGdemcoMkxX21YB/QUp8yx1dya2CfIkMQ+1ggPSBHaRnpbrAZGLo
igpJoKuGFMBMf8Z6LwLMXxfjU985Xjswo6jiRBlU7EsA43vgr43kHZ/Q5b0T
u/dIq3QdCSTsC0YbwcvP/xOCDIm46SgBhpnst7tdKhqevNUre5q64fdCSDyS
5hUoPRe3QXLGraJzYVMddPB75LadmhlhqC9EPgKBaXlFEjmo1gYCQFbC/Eg8
16bdDKl2fTKt1YcoMReZWKC79NZgO11iyFW/Aqzxva/moGVD9yEkCqL1PhRC
j+vLT2WMc+iHvUGyYOh7oQK/SF53ALPG4vqEn3+l639cyB7Mh5pIL7BZO1Te
S1/Wn0nDq0SQBdnFemt6kM3ObUGoR68369HwpUGAMo94JbB3lcT7zhg/gXY6
HuXkUyFtIcarbAjrc0zcOABRUsWMqZ6QeIgIU9p5DyXBRviBv180MAUMj9kM
ojNqDiGraEtIwrnE0JhUkJsCIEfxAAn7th+bpe85Gm5EJj9kEUAJ37dkXGF2
IMl+WnMV4Tl5nL/bpgXd12tll8uB169fY+Oe4PfkNTdgBaKOIiSjmIBqp9uB
dBCiFR5cf/+LX2NBec08CA26Fy/93OsovxKPga291mBUQHLDszx681YcQWGT
XqN0bqmsMu2TVJXRiTgrDH0Rs6DkNXYK/7ehXyh9nJgAUtMt0xVbA8L+XiDk
JnbGvRXLywPAuK1pkvJROuekWOErxPs+pBeZA7fDs2lfCt48p//PdCUlxWto
s4tFjCj8rAwDfLfl0EPt2lxAK/mbcZcIcTxbVCF7ZtcVwT7uFKuU1MkrwlPs
k56OaYAiQcZLMDzeklvXVCwAUXL7MnbJd1fb3eaalPVjvUuKB9/YWsyEBOaX
VNzoMCYAB3QEj+EQkajI0aI5Odm44GpExu/2stvIOyRr4/NXJPJAb7myxFHM
LtryExmjiWooAZv77jUlzyPjNT9KLousOaaaoPsiT9yrpy+PpuyUULG3gzUC
NyKDpcJkTl+Kcc7zE1G/1Vfn9Ejlg1ktbwvUadgurnK82YW5OPbooCPFIUJ8
3tPx+zgBWdLl5I23WX4Oi6Jr9u7mbQxEYBbRWQiOOBl/CPu5zLLAyIgodmnj
iSkX9DkMfKJFnV0ePRTRCsAjCdFzadfReB3+jeXbCF89iAH/QPVaGcNk+ft1
19fALcnsVnjdfDV8GaTDgLk47AOnDDRm8UdxuVDm1W1rG7Jk8F7aTaGlzMO9
VaPa7jH2+uYtHSn5RyBeFxTPe2RYje3+Cc6Z8uyVVI1RE6QtYU+NIL+gKzrd
uVrWrLztA2x9RmQ3Qi8DV1Di/EAzPd3Be6CrQfnMjWhBhWbXTnXdyfmFsYjZ
e3EoyfEX6jCygYOYpkB3ZrcQ6CvrYFFSntbKVI80d0SLmrox01z2NLkps37e
STMBd1sARaOWgAbUkqgPHmodNAJfyxXZ8pzPNdGtc1Ky1b9cihRLZeHvJcL3
JKOy9KsFENdWTk/YTqSrTDR6h2ZtI8g6qAFaWN6KtUA/XJ6dCGUOr4h82dRs
MKMFts/oQakgZ0ghb6o9X0n3MsgU9wRGVFs2zeMLt6A2zBzgmx5ME7qNhOK1
Hiaru/QI0cXRdcAmX0pvrbXSLLZqst3iRqJxXAkhjBiJn3bKWx4Yeta0eqMR
c4RnEEZ0IEfFEphIQ8BNWAk7L89MTyQ48NB52fFR3NagZx/NpXTkUtZ01pO5
71WUuIjGA2VO5n3Vxa1KiRRx2FtpIT2FyNcnNU/g8bXN3hY40qsz65WnQBG7
w7TksGQ/8LuCsLP+Ssn3H+nEOcBs4gVylKRNhoTemy0C0E6q3clWZPtCq4Lf
LtHiAyNZwLdED2z4ij5rU9rwpDUc82+f70YkjZb5y6ZUbhzDy60E6LPESEIm
4Sdij6BmhfLUGdHPnPL2J7S7rnZ9ASFibup5MHdZ/ABQ1lyssDDk8YzsrYLl
Kouj2thk+NKXqZmi8rEXcTogt30tsqM37SVbzECWP/VDGtkQNrYLjSGBpzx4
65DGgY1h1Fd6H3T7evMArW0xfNTr5IoXqAwaUNwCnW7EVzI4a90XOccJ7e0b
4x+FD6bh13X5ueWdKMgJnxSEnWd1jjImCmIttB32FtNpEiNYMOtJ4pMaRTgU
XBZ6WeQCtSVPtWyc0HPwC+XZD7MXcM2Tna5Xka6G+pXGiZpEv4eELy1JTFln
anyKFstc4xrlAIXdV3bHP4s7i1t3ZHPDO3QfvKpF0iLDZUsxO/eiyLZuhpNm
s3v77/cmRBQKju9UQz0vkNGkGbFIX9TagOWRvZvDxSG2o7XS/9OrTHqvMPTg
L+aBEYb+XJb+BgiAXi3b9gd7MhqBIdVHV4ZVYXfOpVMg7CwIPmEHUt+mn+sH
e05ESR2U1KvLWMObaaT96XKgeRGG7HMamaxAAnJoTLzQvykd2EB0AayWxYgg
8M2/MsjGE25a+ghigc0eJ2S53NCknmDZgGlqeyA+Qshc4kd8AD/uYIgSWHEC
r4/vP3rMLZC4c4OojYfrP/f/ujIyskX//WlStnaPtqFO4XMynmDkfHynSW5w
TFD6FXOTlZRO76nHVq4py1nNp9F8C1TthmnRbuO+1QI3ktdKQnzg2TxyyH4v
bfH5z9ppVJ0LKJ2IzzLr3kU5Kj50fgF8Tpc11n5ZF1VdzA5pZfghZo8MrcaP
zEViQhXl+7uU4xvASPtI2IJI6HWl46DMW6F14PNTUWMSp+g4jsuX8qPlxO0Z
87JGY592D1v8eiiGqg6IeKZLygUt64J7aUzdh+SN+TtnPoUaJLETPLrT8rSl
AzgDSAOKp1fRGSAVaQOjinTloUTIOLFUH/J4tAiZpTx06fpw1UyjgaMJg7l/
Pve3sD5M3K50NAab+fIQSN3u+7UgLS1oemqcSlnilEQNZ6ZN4Got6yOi+wXt
mQwYwbRVt55J9/YldP5bysl1Fmk7mVBMK53CjNgjGFHxW4ql3sH9aTWfYAzO
j9BvSfj6R7W61BUPIgQ30YBDUdEA2XAImVIrFFR+EzGG586snrDS6hXdHAo6
IIBu+wqbvXLhixXQgwrXPDr2qU35++DAiwYLfjP805JEkc25NjmzgDxJ2KGu
dyjsX3/jwIAGag610U3A9LpJb84XNyEOGnkHY6t2Re1Fwi4NIRN0LCkeutGx
HXs9kKEUDPvm71y9xQwnJizSL0H8Awjy9A1P7AyQTtjXY+8AX6KD5smdd45R
rQycO+JX6H4/bj84kzmjSBH4DmLku35m2BU3O83gyt3TqbMLmQnCclQGroEf
CP6chqEeOp8kgXqQR/n0v9v5k1R6UvrftVdbppmgrmguM4jlniuLN/o0ihkk
ukVRvaN96tM532tWxe4dobxS5/es/m50P+xb2zEKnyjGIsIbZnllZTHrF0Rc
OZMfxpJEm5t2cGio/Sq3gY4nQZ6tY8gwa9bianJ38c3uvC/1LxtezywKaHJe
SJXfd/psQg6l1Z92MNRA2VBcSrAO5IwMg5ayfoCtHg6TgzBcBZ1DYkE7cZtq
OhCEnFbnqqhEkI1Xmvzwmd0aVViJCeXsgsgB8EH6IBdF1g4hbn1jb9AW3EB6
WgDPo0gLBtIwhK3m0eqetubf5er4WQr1szo/euWpiO6g1cugQwzON/mMyHVZ
sFMD0yzzUEIz9mmSBUwPdp4nxcX/A7vro1+rwbRK12JNoQ9cEmQNQEMJZrwc
DzjBuRGoNXYRQ77For4YSW2FBpFRAXIdb+8dQPF5xqFyb7Iu9pTj2NKbgXoE
3wnE8lE+s2oA+PbfiCYoLs1GJwNhKs+i8qhjwTcgoVasCDcI6G8j71uAWgIj
xGhxAAkKVzWXnCdqlkdltks/jmBhl1AW1iOb2TTphZos5di8NnIxLsgpDCAN
N/QqRVRMgeH8rstkt7yoU6GmrLybwkNTxPl+o7LTs2MxNJc4YQzIZNjBVFRQ
4YhacMwl8bXD+BmKWK07fhN5Wy26m4ANYri8C+ccafl2wGtjtHFCRxNYGUpR
VzTo6zDeUAlPPvGdVEx/TGazLY9JPg0RpZe4BP1bpuUl9yf04+kHf89UYE00
w7WnyB9kG17+4q+KbJdHt8nXkJR6ScL9IV1VUO3tgAOvYeWoOcsokgBY1t8q
0bSRRDD/GHvvJfBu11QtbrC1I0JShgMaK+BtLWcHl0zQ7471t+8OE17WJON5
mMr7LN0qzFngPFoCyt1XyoaZjAd/MrfNRLG1WzgQe6qxQUtyPLeKhbF89SWp
ANXSEFKfF5Au7BwiLJRFljKZDzTG7Bbp34fJ/Htoc3ShAm/R7vpyQW0KGx5Q
iWXgHN/+qZ5+kfxpKGsGq6KHoKw6jxWcM2ZS/hVLOnyjF+RH0a/NwYeTzYRf
vKHaHAPXDyBoHkSq3O0hIWd2Ugf2326Y5q6pYoKna6hw+pfqDMH9KOi90Zuk
h7h6rnBAKA76QvckTR0ET02w/KuY6yPHshaVQccuCG4CO/Gu33rswMG6ofSM
jbWiA2gWk5uOLAKFmvcXjYa1n8hlIgqxI2do7a4kFGDRRfnwjNUQ58et0fy8
uwN0g0gI26u/gSmUCB+liVQ1wzWzY3m4WPWX/4LQgFxlJTDjJyban58OEMuY
ognwlUjSW1NU36XZ9rn2yiAXuVlheE0AUr8OlDQmEiZkxjdYqMo4rhColKKu
niVlFvGldVlBkpLQgoILVFBnWYaIs1JE7t0g79zyX6YZDJ8qhRe5Y2A85NSI
KDxbFoFXEKt35QjEoe1C70hFEw0unYM8OvLUxsAXIf5rBV512wu2rYHzE1vQ
cIHbB9aKcqhQKExkaAycNLOL+AW2zCvI85B43eFHwVya7Y7O2zeGD7sjzAnb
QXzOQSnRJ4W48Ly88/f7uscxIyn93z8NCX+eZw8eiCXr5h/H+awz1gzlW3vX
0XSlmiITC1XK55bDCiU5S+tAdjph/BFeHuWFo0YdRt9YVBeDkEoO2ZIwr3RB
RMy0vAMQSU2Vf5a/4yBOy1DwpH7I43INA+MsvEZRcIjjKT4El/DlKTQiZ+hf
3SaST+lq32iO6Q30oO4o143EnEbXnCXwkDBlaxYFnHAplSonD9I3gWTyZIC4
nasJTdnMLCC7eqLCq9VpxDX9mi6jTYnXmIbVmp5AxJe/vK8nFutNLzElTzz9
UA1GYBLVSEg44GJDWeozhn0ZTb3BbzwvivfEjHxWbApwUardkpeSzbJ3ECKC
RG4d2+WWKGC3JzHsy+SnOxqH2eXaLlsy+0VUKOv4ROBBmbLPrK5yvgcrCkVk
p3ra9yRqliAimd7xmsGatktkT5fUsFQp0O2+t6dklsqbGQ13ttA74/Jx6PrW
sN/xBaoyhpyjn4U46aKVbtfi2yLcFlOlsaaAjzOeWVkFi4v69vYPvRpEeNwM
oFd3hsYoIEktHnqma9dyub2KzWeCjRzggCt+f/AG5i/MmVPjj0jwBgtbws4J
qvRjJp7gO0QjOQU5cmL6UJ7b39bZncKdiPH/7eKJrtPdlQAE3+ZT8r4+yxDh
36plAKCI3qcvlCkDS5wHLdLLaNwtUZhfZXrQc3Cowv8CDShA465O9bLhEloX
MDO/GWGapBVlLT5llrN9wpse2WVmwZEDBk1xDlnKff9MFVtDTU2tELPVrfUj
nLzCRXP0xIJ7JPrNrrHNKPSwMHEsVmFvvam4EuJG1ayMVb5QlK8C0xa6KKyg
cj9TQFQ/h3TUkI6F+fIDDrWrJRUi7nbh2ViXzi5T3CjlpcI1vAXlBRMmx6wU
Z2acfNE0BMO0flAfL7dfU8cy8gGfjWVjPhVt8TfWFJ7HUFabAIgipRcQn/Hi
7iDuHEHjgGU9KZ0er0P8YSlH4isOYR1o9UtMpstRqvKUC2mXxoI3IAvjsWHc
yJC+G6J0mz5q2tTge1iL/3VxUB0cAeALFqbgUqyqOb50gxV6EROugojmLgq/
m3UZBNaqCeKldhEsprWbrpWrY+WfFCuo++WQnRnqBKGGf+aK7bmEuapG6c0n
3zYuCJjYi4ZR7ZSRmMOpjXaN0WFQdrF4dRBDkecZiVgCl4b16EGXUb736mEm
q6O+Cr1CMCbfIULMpkI3QNy53AMlYr7DZkxQmMCA8aP87FsbZIiTS7dPlx9N
wBqvoBBxrzF+1mw+MaRAFB24H2Fh0u6I5SKsj6N1Z9eDSZaNhjNSMcVaPZgI
LGE8O+HZ4Z3Mls5zwUT+tRBGxuPew4NEAT9KyAn5ylF0VsfBa7YrK3pYyex3
zRJH7F18n9681pJTFJ0bJj1RD7c5o+mpK1LmXwohEihKXgExl4cJFJ2Pr3Kv
Vl5lxV9L+QuaD78UHzYZ1js//GpZ5cqQn/gg39C+Ve+Ku9eJJJLYr+COGh9m
JTbcReOd9x61fHeiOJIbGpehae+CMdwLmBzDwNOs3E8/LASr3bUb3OFzvaos
SEQ8UF6uc8qZ1a9cX/Fvbp53uz0BLZSzLSNNbhmR7O016DF8MTAWreY36xi5
PK9ADJppHC89XJYXC2Cko2dyKKziYoLJzTa0duhbWrmayGDavk//TMeQsJNL
H+2QVScgAumREfoiZQj6vGKNMacLFOJUprdcEtKpJp4Y1SsuFcknV4Vwjq22
YTgaC4o774fNlhZjqd5YkkO5cMAPgotk2vqe3Qt7dmKTSIH04ePRFO4kZap2
w/4YwwqdUdDmhzZ4lLnQ/z7oud40daIW2R7snf01vuTUf+vCunjNwr0Uc1dm
GqzNEcLcX6ZM6wsIMHGDdm0/yWN1E0Z0uxeROqRw3mvc3gyA6KEAOl/x8lcq
namlnLwEkndFIrgyAO+xS99YMrMsbKLYk3lh2AWmKAJrIYzYmu8gJ40519Jt
+gXXFA6nuU8dgBNfsMvnIRiM7H0edFa07OJVDcSZu/smC5yZYvrm9T2or2R7
mC3SI+wT+POHGy9RuBxp/9a8KCg5rBZfg6quDm3SSNxCiRjz80aKkR+kBlqw
2NmxX8dWOI/86CYgdnuM0BIOIj9/cGOaJV1RYjUbBRLPrWb3YMbxZtZqEBit
2sNPrLm9N4GNp7yD3b6kxYPCA9KZ58u8ieB2ohkptL2lKRACDI34nHKQOxvF
KrCuywfZpgv49XyDsU3Wlw3sUK4R/Y1IEFPv9KvYUv5LgqcueSrHCJbXZPh9
0M6i2LP356TpXJj4+l5D+mmL8/tb5F4vN4UACwphCoM1nUOh6qgV1dgtZ/C6
bk5czNgbEDXjK7NbTGF6DzZdv/152lvAwLo7WHAwdf2kFIYubM6H0JXSzysO
6zbFy7IY9vtZa5beEjsi9rPo3SCW6ED31V7JPCh08SF7vqDCa0IazqMJNgIE
/w6SQWbUXqjHF+5GrUve4hgJ5QYX/Uxd/x/idU2AvuRmklSR60MyGfrXR2Jv
eu9XdxAvR7Cao4HDdNEU+NCinkXIU13G7he7h/GPUSbQjyfBt7yOnIv3FZ4B
epUnNoaRO5HVJzlls3I3nGvkB85RBT1EHB0UHM5aurr1k5MPTC3KFPZ/l3oh
SLti5duqtvsmV0r0qB/+Rma+MpLslZNbRmKE0qyPNytuoTeCFRIabt7n9m3/
Abo5qfX5BBOvcHhbZbTk4BlD4JQ/DRee7jV7cGXTezF8/6iwlNHQuv/hZ1zo
3ME7S5DI3eL3KasAs7HucsW4dEqQGjttdrVteYjCbYfHuhMUE66Pn45iVC1p
A+6pCkAWlLj7RsTma+rQk82BoWI+XxIXCkxL0IHQrACfuVN4lk0eY6S9wQFy
3IeCPPIjJfbsaVbbCH8mXB9q4fesHqqCC5hPKhTJ2xJwDCE9kQNGO36Lk6HA
iN/DXUTTP3thM6jcZKdZPHjicGOAkBO0viQlKgtKO+F0b8rYmyOXeGZxucSl
aNWsyj1/zvdnNs06FecVp5orkt9ARkAwuxbjmgWkUFo5wmhUxQlDeJ0+0W6T
yPPhia58rLUzUbRq6/wbX6rogcNH48Zn0GsQg1y1UZdzaLybHAWQEnPgJISu
R1Ss7OXaLiYTfwb5VEGqdii8RhP+gTMHl7nM9MlzJjhd8AfjcPfxQt5Z7M6x
rMdr3LPBnZw9HTQfpCHEWmY4ghpddlAfEDJKWScwXxS3/6RxmMEYpDsMpT1d
1kTQ5zewk78wF/KgOaiQkmTT2iSw8ATOTOS9NyP+9YTRtSjS7nfliDo7aiLC
Dsyga3TXbcraO8qMciPL06lzlr97xiQaup53RlpMwrcxUebQMlQHB0W6Q9lG
0yz5w2+YtPbwCsTMtv3SUlMv8xQbDFm2p+4/YK5Q4jSJaWXGw2AoQZWgDuOq
ynJdYxvpJ+2jT0/OGxbqZ7equcQ6Zy53SdB8lupjBZLG7eCGUnGYV82CEOBg
OWEoBLeGjyGS1llGLMo+KH8egUujsSbBFI7hcwFhdgsSO4/BV8RNWzAtCVhx
RzX2GZosvfp6H6S854nkdiAO0ZK7JuunG0asstS4i5is9Ty56SmtsoVd2pC+
DXekg6UimT+6QtvyWeFxVcLGFyFejbvmmRp4rFQZBeo8Fg8NDjEXfX2ugNkT
bY0O8A3v9Msz+BNJ7dkkes7/Tu5w37XGJbHYMcNiGV+fVQr9v21BLlcjHTrI
v6M68jli8qtz4bX1McORfojaAGAIMG2tfYuQwoaqmH/DZnxajCHQjrpocx6z
Bav2hkdAxq4hg4Mclr10Ast7seWIavZk56tV8z3ahwZulG2zsVcplEgU5Eue
4OKU3pbWMzxjOeqChLLLPjxeEbAKJcGVLVWES/db+HfS8AeUMgFzioSLMauj
e5v+r+z0sy1xHd7aX6pkYOSmFzBMfTVDaLqKGWAAbOVef43XvAi2E2gU0kcN
hMzR6zYFBKixLqwE3uoVSZoDawp9n1OlYdSAekJ5dg38hGqW1iaHQzHANRuF
LN9DacCBGrmRd1fuTOIZpXyKb3akk16DgNq24elumI6om+aMiK2SXEVzquEV
51ImpkkyMtVRjc3QYi6ZNpMqmOjGIrksA31JoE0jxiTw+Tg+m2zpqPW4ddHN
5FAH0kLihTSCw7/sOvnEtTxQTSjE6pys/+2f9hsHLe7f3YCf5KyPHV7qdqIq
cnOURBKYLrV5d7LfSOBz6owQsrpPPfJRuiCVqq0xPUYAsbQhrblqhYOugsaX
ZhO32VoKe8R2EDn5hStIaXnNcS8/PVQfRJKEMPBwFkxtKCPo9zDnYiTxLUwQ
IWd5xRIB7nj5XPCJ7oTDg2k2AuF326fdwVubMNK3J3OE7JqhIhBZkvsZ7C+t
Qf5sbndP1d/RSpabpsinon7BhANAXQquPtocqI50XzTEdn2OVgyuj0qYiwhO
rtZLG5Ej3x4oW0zM4HNvr3uVUIFlM94M8yZ+VBxPAQr6Wrtq4Fp1vM5QHnNE
R5M7EgKlmkrqMqGQMXgbrBh4xJDf9E0ys/ZHa8/g7Rfl/eS2VyZFZ1wjQK82
OJTsxfQo9dklhLIgCOvm+q7HlZ8NcMv1tSLqiXbv2Vwz7tFvTOPPp22MaLn4
h+hpn5npdIAGbmquMd/HXqVIteBp2oXTuENdDQ+9IpDiqK3tqoFcIwWNyQ56
muYj0lb90G8dH3M1XuA1pZC+3DqVV5KlJXWC6uy4gfeYGmlvy9NcBjFHWCS0
LCX+YgKAoxJqa3GqLeSn5wvT8ZA0kyD6A4yNk+RGgNpnRxnp9kHjxxw0Kwfy
vkPnzU+bMabDgUbTpgH3N4YVm1glHa12Y8r9aiM7/nrTKvt0G47Ta/0ftEkD
mOlU6uNvQzAqs5zFfHlhaMUhwYIO+fUOIePD5XZTZ68h3ShBWYfNRJxT6SAK
wR3XrA6Q2PJEZm83KTfX0919IiDz1T7a7IMbkkU61f+fXpF/S2Vc2ZeI2Lfu
Fo3/f3WwzNwVjifAWTqiwpnAv+KeCJK7oMkBuMRjH8jNwQleKx1yT+uG274i
DpYgER64J3eeBWXLv83r3e5mTtLDUvqoPtBW7AQjDDaxG6o+Sld/HSre5cOc
YELv+cI8AXInoWkqQnC9WxLtFgfhM4FE4hbedOOriiwlTZkIAcn7/6h7P+oA
XOHbFtTX4seazAsnsw+NU3N6ojMGFHH+1EOl/PkHXM/UAJAR9lCgagccpauw
4JSIJCh8ZLQZYnKLKaRsTvwnXlxYdf8kKE6eAGzRQvZQQVirYiyLJy9heM0G
HEPyxEfklBV+G51CPA3KhmwJpRw92N2F7VQ2Kc84oMPkV+Ikr0rTW3813mNl
fHK/ryr4eeFFnnB0FXq0dJsaTEeWhFr4/dhYBN1WerMVR7spAkjlELpUM7xb
jHBkkyXnZktfUw/ZMTGMzEUdcJQ04hRq8z0KS7SZ4XxPcysw3Bcj8iGLwTDh
lgOCHfS1XHoufobbzsxzq8LPsu6rhuHGtrdJ1oo2GhK/8INZPlGhe75wYkev
RE5sdYBFrGZSEe7J1g1do2YeDPiaeVO5Hn3Py71mE51yXuYyQQBSt39sa1Ov
OtNDQD9vliLfNsbveAoXs2CFo6BVeP9TveO2jBsaEmOLGmO8AwkQXFy42SJ7
z8jJO5ETBQnyr1qBURb8ZaXFqEFP2U6vm4MG8HkJwqHV8kFzDWqtxw25I2Fm
OQDL1uJaJbLj2ZMQDcpxGvAeG1tB731WJXM3ml+8jFH6+SqlO1dvK38b3cBy
yCO409eb9tdDf+dozb/XT/WAD5iaLMb05J8GoCUKYbO0GlTZKc9AKBVkYCcH
+u1C949sfnNWZ8DJPofTgNRYiI4MsOhoxeInWOMoOJK6ouo6g5MznGgSOfok
ph2A3zcMfLUsmJZraIE+V7LDNAmEUBq84ciWzwUm6k9jYpKxuuSIm2Xy8FFG
JlQzulFFITp/5rqdKo9oj7U/J/f+Cm1ZXOz8jMVXVjOroOdtXnsNuNrAhDFn
CqqucIrfjnc669lCsR/1w+pArJqd9OoVvrW0nB2wr7rh16uk93/bzYt4UOp0
NicRvxO47CevyOpaIoNI0NGw4G1vEGe3Ms/746UkH4fZuGc30ulXTKkL8iTa
obFw4Yt2RFwxOq6QfkLtF5lrnPH5N5NoYs63pp8V5sQ7oN6Ko+Vo4AAKfrbW
69ATeoo5vS9OzrDBFXKcxIPrSez3XlXlX6FeQuz/Jbyg2w7RbJC2GBWI2xPJ
cLqDnDtdx1nRzXeVg5skJw7xRllRKcT49OV7kjQBIsAnvf88vx1CrvBcZWcN
mBp7RSry2chYAYmZrqVUgfin+DbhuF+BhWbCaJyjy3ChGygt37gT47Z7hBa4
RhBD8RkqwFmzSdN8n8dLkg7Mntt8zSRAViXY2PvJNehGReerK+UCuk8upMpo
NORRp03cWMw3GChjEDGyITLNuGiB4a4vjDbRlpVGLGfMFBnDFmHv2ZnE2Kn4
ZPWGLDnbOwf6+zfsRnykLsRuJCiyo3+Cuxp6KumGXGvXEOrBXTvWb8hjifN9
AAbeu3+Wb+dXGs2b0q91UmEZXvv8D3iWD/U1t79c3q50Y+3D9bNa0axfT5D7
nUG9Uq6pDcAl830F7O3Tag3sPCtvJkt3mhRbWgo0ktwtXkRORTg5Aw1mn2Y5
Z2Q3QdKY2FogdCsCT8WuFRdln5CbRUkmvKUSiIYpbbdi7KXSHZ7sTHOb4tOH
TwkuMRot3SN4FnvAFwhwWYlZ8QpdY24Ox99csVh5FpurUZUR0OOJDcR+D1jI
tLug6PUSm2MJPvlNhcU0qYYu744laQ5gm8rSHhzyZrKG/KHCFO3TgSLEhI4j
XcTFKGZDlMxneZk+MPNrNANHeNDaGyo245YI8Hz0Q6WCdJO8fH/N0GA9RWeG
37EuEBbK21o9XPa61JzUTwFseC1cqUJc3HsvSH0Aa/MMjNKfgY3YwR9cDzAC
tONNaHJ0Yj1T7hpGmqwDkT2i3lqGLNQR7xlqEI1Fgo1nIQWEH6pE+K+KBszD
Pv4mP2NbkkV/jPIXhwUsCKFvh/y1pqPTnStb4YBd0cFwlf5FrCe7l2Pjrw5y
jOxN7pY+pSLG0tMtNMVvgMKZZLlYEnQyh4iXIHIqnGEeaWIhr/ENOgTm6ScE
gsuR6YY948M8AkyeaXa3FZ/pthK8kTTloYOT5tZ8tpQdheDuL62oYFVvdubD
SocQYfoAXgScnJLFh5rrqTQKfWuUjbz7S3Ldsx1Sgzd6WH05Vje6KrVf3iMF
6deGkN8zWkszA+LAt7B2M2BTlVq9h4/NWRql8CCjdyi6i4nx3+CzJkJdfOCJ
h6hRwL1yUrGuyscvZ+o1nc9oiozBWo8tnVKUx+oA2FUixwLjkl5KiXDAn9gQ
+uGL/Oiw591NyN9NUfolTara1uRHYDaiIs2BmmocBk4HItEHJ0ZmBE6Ki3HN
mPw77DXSeSYmHU0m+zuVIuI7fuMoXx1exToaiglegMaJoneQ+yjL4k7v/5sz
0bfik+Fua+vMYLAGtKTkul1HPh8nmYjY+iJNbwINtGAD0FhZgYUQ4jFKfItP
Lxt8ucs2Q5xghIN/VYCdWCoQUp3sADkyBX3f6ow+KReJY3ojt9I9w2f9TCC9
t+Znj1d96JQaurrE3D1mMpDGb6mnkpRSsiBi75kGOv2sLc2fr2JmLigNrzxD
4jDfvnEQBv6e+x/gUI/lJliHb7VCHf7ca9u3hheTNq7ZND+w1hTuTt3vOHJI
06rHCVcj/n6fN7BBaGlIGnWzgaoM8x0mkXmWVeP/ED8ni0iPgrYvqnjeAeB/
Zc2LWOHu04Hvo10IlIBXh12/NWsicDSCM6X1YL1qyXY2rcSzfLdwP6dCX3QW
KiRTtEd9o/OlDe4Qdkf2whaBquIQ31LMVL3amTmg8ZSXKwOrB0o6MrsWZwn6
KBIjrifhsj3G7wg0VKFW/tar2Vtr75de2WLtT3bdHQqfOWgS/tAvIg8WVeMZ
FWcvHOcflBJp0aQ8FBYefWdBcAZS/9tLysWddJHh3zZFsUl9/SW/WsaGoOcq
8+XYQcWn4sQ7BKq5geEpgGskFy7lt++sfVfYOIDlfwv90UmXm1rtSoOEsrTe
UIN1MtwDEAxCesFauklloAjU9lNzCEOqV9QkTVOp9NpOGq58kKRnhKR68T0w
cWaW6Sm4+4KiDOW4FPW5N4IfHCkEcRQN3XR2peYvDqDiHX80Xua38/R7/0Zx
XoJBIdMytzLoKCXDl8fBFwIr/ARjSMVmECp85KRaNjt2dayMfZyZ2yrdruAA
gst1QTLSYjXIyjYEL2f8/p0QQ4WPtGQNg+ZAavRN1SslZ9GM9/53GpeGt/VS
1NapLnfHIg5ek8AOAr/LyrOGQBro/IOo1CcnxiMsRiLdLVcUbnPUbgdT2aj+
3LtC6yy5q2DIfumG/iTt9KcfTPn3mg8u4PNiBlinavvpwedWGCzIvPcuvm6f
h/pK0Vl9UFnXTdVGkXuEohIbTS2M6YDmbZ1kbBT7+9JOmkiPrKWeE7fNu0Wh
NDgEmCqfyuGokE7X6pL4DmXf9ZG0HIDmhxLdiFrBH2c0qeOM3M5wCKWhiB4t
6F+W6vnSTdR07QPpHq4QxGKlJBJkXf3abGLqgcIUdQgxdvQLnKH8nlV3au6f
9c6GU7nV9HnBup9TOaduyv0pNCdYbsiWTTfEr6/Uo9L8sjG7j673CNHdZk4h
OnxMKNgr4eoMZBLdyGzxj6EsFeNg4I4a5KXcs9qVp4YiuwaD7aF/c3nwumh1
qYMIy40BqpzY0q5fAAsKqFCwUtzAGnPcSlv98Ai+VFv+JtG6cHaiDZuVqHx7
lOnz47C3fiftnawONrBrxMBx3ZwPFGdOrcSLe9RO6QJpZ1cpPkL3zuQAJuyH
JVCHZZ+bfknsF1OPL4eY6/sBznQgcAKcmd58XaTO5R+eoedqmzx7NpGlhzz0
fuSPMlVwQ3Ik9vOpWsccZwhcVNPKQA8AEY1tGLS6TMZaLywLAO/Xu2kRBqYf
HEJpd/3p08fma9tMmO1uO/bwosoMYbaqNRYTL3xlOXpdlPUa3qq+Xm93rFQd
Ftf2Dj2sMxuxDieYfLEQ4DoSYq1SJjISD8dsbE78fbHRZFSQA6L2QUWaGYMl
iEuq6xl5FkH5gJepfRoTHF50vLPoCfI4EPW0rFWFoXI5GD5hUoio032oY2V0
e7rD3mwTTmcFGztv33ukJ/5AuQrBQSQxZz0V5O5gUvrRrBqh3iEeGcUbv+Ay
vNpOwX7iXHk15PxO95jgo4iI8f5KY7ShHHKn/srmWEVnu1M3LXiClOYbFl1A
/UcghtFdCk1ICWiYxetXA1auPJfKAvtfLnsnu27Zj8Vk3Yke7reI1gWcKX50
OkS/EQi3ElrVcpLiRte2wSWUtVheex12sfbFfcRAr/fO3zzJTYJOuWWY+a5C
fjps/AkwsSBLAi6o+B+GUJ9yRBrfB/q0W8M9CC5m1a0bVRBG+cMVpuJVc3iL
oayCY7Bwp013QRZ86B8lOAbFvpS+CMhGEt0LBgHPDP75RZviWzUVqkO5DeVK
7EaMboYiFF5zHw+gzmLRnY57x8ba3blgDGp3rtV6Zg4600AAyzE7woJA8sCL
F75eCgKP+jqqMZ0wIX3Mduu1y3vd6wfUxvw+zJNrY1hspsPx4jUYj+dn+E7O
I3Vry/abSMfRDbJSbd2v1gRfXgXDpFc3cP4HG6Vz/TJ8gUFOr3b3tMdovoIt
aKbKptrM+E57yYFlhMu7sF7x4aizMqItdV38dgNs+zAE6jZCh/ksm/3SY/7E
Su4YjKGQ+2PR1d0w97gtHot2XN0ljkAtiMhbt/k4wsZhhuoYZadk63m4iqzh
h2eLLc3yAinFWmcJnV5Ryyu/AvVCK5AzYSXt1xeZCAOFr22yeHZB9aO73TRC
J0yoZ5UqwOCyGbPidYREVCVFfGRQTkNjL5nxpFrLdoRf9rpeffuv8Ke/oasz
tgtwSpiV1PFEtpRlLhGyx4MxMIALDStS+JT4/0rSNGMjfbndg4yLlR/gnczJ
yzz1T4YO6CBnfSYL4p7nVcuNt/mtMwmp+3h18Mis/hxd0BXsO/37YIgVEubr
AAVaWjgt2YtNkEk0hQzdOO/aFB6ymQ4imSO+31AtlCrxY33rMCw+EtF8OGHn
e6lFzMv47enXqIhMyMjoqFPDZxHRHlneWBtkUdgB+boPzRn6n7mxN0GbWL/q
Ddg0MF37j9+RlfRZeECeu2MBdLSp9rbvXYnkXFiqWJwyR/9QSAeOcpMX3qGL
Ehm/rClDnOE9bv1EHL+Vce14NvP708S6sUQOpdXcXSC8jzgaqyyXio5vU+Ir
yvJcNzcSN2IPewk5WsVC/efvevwO00BK6RAZzB87hCFqNf7DyIXvM4m5AlAR
LNN2/UzLiCwPDKPdWHfTXxmsRtyOCWtdMP7BEg93OWkn8a8c8fNuHnsXjkMK
Jgaah5uhvsBj2FnEycGXCZ3DBlP27eJJmL9g/uVtHeh2uMjsipZW4GiNcMKZ
ftEyrfxz2zQWkKUpHM/f3pmO0HUtqqtM+3nUEfZwKkMNQFUHkZXlX9IZYnYe
3CgXoCxIO2ugKYm6uyXJ/FmUNUSCHEK3L9IQP7c3Aus/3us1682c/bUbhgEM
1EJ6zdC3hcxUk3IUQgXOZ7vTvhacqUEiPIC98xgxmthkdSP1DXREcRmKTi5I
nzMoB0lH+EWL9ChQjupL44Oqd5pPKNVlXCQ+x1wRraPvwBahIBbYvudVs5q1
ZM3KJFBflG4sVEA/L4QAYbs+nDOS7IzDKEOcJfMnnUnneKCVvwOe9ejuSef9
fTqd4pOUWfvRaduJsHavoPwD/YHUqQBC64nTdwWKE7h26kU+IEmcKiPKyinx
E6qUkxHH75G2UHlO2w87jpcoIKfZU6+ocGxro07XrXbkUwbZ7MzLITZRLUI4
eAeWaDGrgrxbOgwKf/zB2pHs+eWec76qvkC+yiGN+qwHBnCGgAbC0MtNqH9G
FXq5ttrbQ32vZlL70fIx8XDehTsJJ8X3uMiqsujmU9CohH0XJS7DlXsMerDn
LaDpukOg83QBYH95ba6jV+h6xc20J9PiHeEvFMo7M/sdAB4cyHmed3IRq6A+
WGQchsVYLuMYV4U3ivEGsckDFJNzcv4aWh30zXPwSm0HHwIFtozY2h/hmwtm
t1bk0eIAM+KBbCLkdDatLVp+oZFYm7M0yPksDkJ9uptEbZMDJQCNkWF2zq/y
MNEUk9zzCUgW4/puE1UnGPU7/TXDborgl7QdZG1PjWI6yb6Cj+l+cBUzsc2Z
4cXoUEv5WtV8Sxn0s6sus/XVVOlzpUzKCPRICIhm5zSguW718PNkUrZNNgNo
wxth0u0OEDutiNc4wj+ipTKLo75kafACAnyWvnJ4P1JpMiqirPDvOdTphf3P
54EXuT6bNu9DAB3j4jggPrcOntj2GUHPBnBw9kpLioSZEOXbckFV2mxPU8ST
F2gKzfGbVkoj47uJlTW2Hn0NXSAW8fJnPHG3lBYa1B6iRW10EhXMk4jW5VeB
NUGHNjdJfWMQTsHqOAWMoSvsx+U3yWv+9g1G4RcuC6p19xejulnMHgPrjAa3
jEjuoGj1hzsd4ObaYKjlynEc4ASuj696eustbCN5OHluVjtR+2oFD1m0oMcG
5mqAvkz+fr/RiMtdquh0udxyfqarppu8V/S+lssqy/y8/p8lgOmqWojnMOrx
Z3QIEfAu/WzLOOp6CuP+J8Nogp14GRZ8BO9V8TGIaoIOPpYHthemOADWW0iI
s2JeDXHfziQV3BqgR+8KLcX5r0Wmlb1Q+QBFDavNA5Om1IviSbRsxkkM4rnq
CYvZEdkyxmoA9WF3oPLkexYEHYDjEbgqwA0BmNQurBmngDULrOOxUU9uX0/x
pl+bXaePS4773+QXnkWthACLJIqETdt/b35C1gwzNwJ9b9zfTGWrc3EzBFQ2
pEL7hKD+8V9kZUWPZxe2+3hUSBz83Y6QuOcOdrOnugtfRk3zLvbVb7ltolPP
N0Q7tECUOtvWQ8FbUkXJmBq4udDBQ0AF8bCPfRerCNUXHmrtagfnxXKKUH9w
RFvvaAkmJH8gkAMdvYSmAdRiNC+GAvuo1V47COOq2jWpE1neE433IgaC7JPc
UtsoI7dBs/sSQGIwI2aVdPyt4JEh2LDJycRDv4bXDYSxIrzst6fGc79AUcxR
uobijQ1edEKz6Hi4XzGaOSUynYjx2X0OfASywupIyftNn4ICAOpzVJ0RHUkV
vSPs4bh036PynCw71k4Urwvh+6HzlL1lXXoGVpitq/OVhPRGBBvnyZsEQmpe
0GbeNyXp9oKzfmjqSZG+i/iSb71nznrerxhC9iBn1UgWNUlvetI8qbG6rnPh
xdlsbOzZ78X25tYHnBjICVrZaUssZLAz6ojn+FLE+n+wtTBq3L5n8yMySaDu
YyOWlAj7V2xkq7FEjE0PoOW19tS1TQjcebRHV0a6bTHRn+P/c8CcCkDFonNo
tRfK6rFcJMsPZo2JTZBVuM4ouLaNrwoBRzyJ/nFJPrnUq63wbSLtXJatMwz8
pc7a3GWhgYSYZPfoUW509x9xNLdyJ9z8/kIomvRCIS7eK1y7czBYMHMoiFL/
BQlQCthGdtpSC1OSNL1nMNWkKr8EPwRckol0lM1dRfx7WvKgcvlRMB/9OfBy
/9Y5e8BsOknSEUyb6a9mrRGv9NJNMbh7Q3oVA58xTSn7DWcNxZ+rDxsrgch3
kLYcZBQLi72wy9+xZpQMNtAwAxzPfnJ5dKA/71oksEzI2bJxFBGXpDN0iUgf
IYrRP9djr84NTIMPGtjt+xEGI236j2ajw0vW6n+gQ8s7WMe8UodhF2iKlP3v
wznIFsCE8WmGlun7U3nfj79p/lfiN4WOptX8bbCxXhzJxCzasOq4KOf+Eu/F
6ZshIOiNNo/77yNfElPhX9/elO9A6Vm7Ib0e1YIOZi8wg2/1OJZAspfOM3sf
kNKINoU2EM85pBbBiBzzxOI36sGNBDSDkO6LDV0fz2m0L8xagepVZ8evTD8O
XMEo00wWbzrFLlZC5FxRJrB7JB2jb8VwDozZp11Pyn5FV4dVswWu0U09BQJM
/oURQJZSMnGHw2EMerRIn45bzRjACa2rj/Y2owmHSFdmDxFDGzoajRk9rQ/h
AUwF3ch5+IHWd42T792N9ClGM+QHqVce4hggLknz4g8sAFjLkAJSDzhT9oor
47JTWuCUWd0MmedZRDZTMLZQMSlXiwKR5f+EyApxWCW1ZpW2iTukmSczE5xX
0wCt+ESCEoPfftktPKA2DO6bHxdNHBM1/hHWeHU2pSlZBZmEGWN04X5HKPKu
CFcwQElES+8RfvDRb0XM3ycrIweixSpA1318TbqMpcE4pyLqrKaGcRAcRtiV
HP+VNpjgI+Y3Zz6FmJwHER8j1GDVaPybNQZnQ4RpkVZf12602AJsETHooHVM
dhzAeIf28E4L5JfMn87us7lRf+hzvnnfTwqSxMw8QAjVWj77+vc7nHidpdVG
Wic2GAgXcmsPW8bDN/RtEFAxBqXEBVxnRh/L14FMDNFja3luvBTmWwnc4D9G
67YRNelzyzXXzU1hiLOilk7jWSkFZVgQq1KP2FSUv4kmzIv/MR3n1lHJWR3U
LSUXcE6DR1IRGp1KcmofGqbzNHj/fx0ldl0YqFM+5H17UOYF31ncMBuN46zt
TVR17zqcdgqjrQbkcoEvOSjwze9fkQza1fsnlEDm9XlZESR/79BSvbUr62Nz
YGpcJhXWLiiS4NSAR0GwCYgX3jywGHszls3xOERQwVl1ehVgk1jL3+e8K5yv
/KutpO7r9O8SPOWUvuvmBXYtEq9kgvVkalCJOQepyaU+Y1jeJreWLrTJjEFv
5GiXv8kNUQ12ggv/3cBp0HZYYw9QafFWnGk0hxpfL8wizEeVHVG6/ECnUgfj
trHFm0/NTboBYZistdVPSNRYt/3vxsVktgwyEhHLJGTQea0bNHS1/0NWBTjA
jsdjx1VGdWHOU3jvHNZITQA3cdUrfiRiR5hT07v8llOzPt2XXKqlgMprM5Ov
i2XIP9lKpCXI8KJ52n5tVc9iPk9b+oWsM5Cn4yYGtTvsytdB49vQwIEttwZG
n3XiyP7SsNl1SYmHTVdznzPDbvxrRLleBCchC/iRxTsuMLZGwKqfjXO1um/h
oc6vJt7+Ds/JE/yzPF+nUmNgS9lmU1N6wuYvT2wnEoeMvDqt/tKy42ir9P3I
pFi4XgntMYCdHf8X9LRsHES6iYoYw6pAYV74uxcwAuHS1cRGvTwiE0EPVlVm
4VWSfTnipXlga7/RC0bG32ibGNZxBsbBxxFckrte3Ausj2Hk/IwZtcVKJuwQ
mG7PACrqvR6vQEFY4uinTZUhsAjO8449quce5O0ub2itvEsiuNaPSS8KWbiq
8jKb7/isUEmBXAwxzba8gUOCwm9tLFfeWU2D22sSD+ZgI3zcIhixeksHAqu4
I2vk0E2PP2QBLahlkwQb0cfdHIvb7YgZLL2AvH2fwH2iyZ+EfR5AwaLykrEf
tLKElDiMOTttvWF+3QuHIbcs5VzJbvu57YaGs3Ta8IknaTDZlVRDxCYPPB0c
oV9lYvUvQb2iWWLKbgAB4sz7Oc7/RuEde+T5lGTIhs19bnyXrm57TWEckFT1
3Vma2JcztFps7g5kyp14mpQSMMtVcLu2UhZ8eQVlxX/DcJJQzsX6eYUACUQM
k4wTtS977BVU6YheXGVGF1MxFw5FyoBC9tEPJOuAE6PlKXVVrF/r0UjtN8oh
LlT9xkw7YsnBzGtm9vWUNZsdN2ZGvtXnWOYlmi5HOgA08aSnhx1joiBaxIhk
P7y0/ZEgi6EcLcQPloUtdgqdHrkz4LBJtx09kDZ3LBI/IfjcKnjuhhe2yzhR
ip5g8rbENbDNQDgdzVaRKPBZYLfABWzWohvAv5bv5xUUIp8YsXHNuyQe7IGJ
UpK76wTCIjn6LEnZMRC0mI/MjdHvyf5eoHGr3WMAxdn2O5ol1euNbC9NZFVc
YEJ96kpgc37t9UZN8XzftZ5J9nkhRxJVU4n6a0yHlmyNMvolOP6SnRlxykse
vR2SsYp+T0aB9ucbpvAwdNmA89uXMck5uKH1FC9objj00KLkCVCPa//IPgOY
yCrjIKx862t8FCdtDmLN2OnGxP10fwa+8pNA0z5AOeb6w2HXavjs8hwh+FCq
rCh9rQOoZi/qTsJcT1Li7nkRKObr60dez9pyqWILxoX1zrJSJ/vM2umvw9rz
4hEw5upYiJ9J8BYniyzeQAB9EyS/aa/WpjwM6W6fMdnS7gvEnLBfeu4OxORu
9NBV43ekMtkitpaGaBKaYiqcH4dxAo4vf9aYFuakSAq1bTTCVHbkXqopTgyc
WCUhHfpvvnrv8sT+f9fJNivGNuONg/SfHbCaYcdode9yOfwwpnlca8cVBp7j
xup2xad2PiPJYoDGhQhN43jX4x9ydeGDdx3NEH6mQm0d//E6kZM8BTBlPOOw
8img22KN9sVwW+JYi0vO1hcyYpIPagdSRchpuhJTK4wG/64GesZ0Oi8fMsxV
oolr704ADQeCdT9dGIjqZjS0CRmqGkyJLyd5DT0tzr6614r1RcXQI5cfgWMp
rgYbPJ/tV3luqDn3Iy6y2okk8Dyx4hDLULaNj2DGxPwSDDs8rsAFPMk7ZCR/
5EK6jJfbyveIoWkqvAvBpN8Cya5iUJGk+N16KdtCC0ctSehsz+dH0cSKTy+I
woSY57sIxUFfqBqYunQrnRXM0f7JnOepD1hn4uVXNYH3zgeKb6+2ukG4xKWy
ASgoSGH63jbnLzHKCugUxRs7G/6GWlVmGMcSLOjv0obeKwbpJgN5AHjsh/W9
+x8mE9JVsGcYO/Dt0UhnU50q+upZF0cuI7jVPeruySUZOa5mlogqlebEwPcR
1+MRlCt1oOikZeeF8deo5vC3bMVxJ4dwLq0fwlxHJ8cIzMSbdOEur6GiZsic
J/qvkCRu9xPviz9D31MLmGCZIHN1EL84DU+je1DsZyM+DAPm+56nZoRbChJj
phy9UZeWJk/f0Bcjol3+d9bYccm0WCO0lMkiapswuv39oPoZt6MK7b1MtYVk
4llg2p84Fag+bIfaOPDQpgrXoEAZq7hM3S5kRNN8doeZ9GmT1mFVJnw3n7eC
4j478CshSBAR6GtzuSXwXjOxNJ5c9KsU+UEftaWWPvEbB3SQKa5eyZQCKVcr
MvT/dya56LFQbZk+h94KcpH4VhQOz/7JU3gndl17zuACjHElS8Nz+RYpK3/K
57KR72/LlHD7xb80dg55r8LdGlVUpMyyKaJ2IkdKs5D8Nc2rInLxZjiuftPb
b5XOzrkjzU0+ET0MpmfJdkmPeOK2qzkw05ErlXJOqnLhewEQUrMiPCFPSVYy
/295b5NnZvgcYqrBk8110m0mLJUb+wjUylfnALoN/UUFJrRxylVe4vt0L+3N
NQTJTXRSehmSta1/7jboMWrGjcHZMcz7Z+21q9X2vGiF/NQeocLwZTUeYjvR
OX7y8+IkggBG7xQ/bn14UuzVkS3QbbNXXILieVgIDEfEnuMTRh5P990YsTJG
Ou20eZFEuKsvuRsgpeNanUFWA+xtl9Rv2cLQBwS4bZN4PP379ExEhWZv0BgJ
Wmc3pClHRvcp83GEfs2ZEOSq3k+1lS9ZxfPgdmNQ/Brmwpy+Bn62ZsecKNP6
SoyYNqXUF8G2RJ5SU/PMR4xDkHZK3Z3AsuP80m9iHKj4g8sfhgzNocHQiC70
g6lK8HniHYW5IZABFCeYw72tOqiKWWuIieLKADPV0/NM5NUAMgG4IT8dedCf
Agz5TMjWMVOSLfZpE536IPdHYhkbXTI/UY1yGTqZ66vtNRKfsMSA44ILwkUR
xy0FOFF+C+nh21+dUOxR4nafWj1+DBnGkLOTEHhVsSTr7oHO+kaD2ViqlyFx
rCS/LPtWltn4rwcStnN8VyUoFzhzaaDZUTuF/7PZvpnIGru4q8aHYscS7OAO
GsazeKlqqJTQnsMiQ1cfDlFMMvsdeGOPXy0jtDS6a0CzLw2rbOAUgIHI7hfe
XoZUY4qxd6Df5YSDhY9ZVhJkta6siP61RRuwU04iWkKXaIYFq+z74ly5rqMw
yoddi9mDVTGn5l7HzBtFkCv8QfyrbhIkY06yaditfYNK6GqXyG1F1Uf/JahA
dhHBnIHtrF/pngf6NGInZTp+uEFiCbMpmmuxoyRkT2cZ9mgyIGnEhvjBzswH
b6SNC6b7eZ7IAAW82th6cfx+lthqyVopYuHM6UVMLNVBCSP4CsOSxoOMr3WP
Sng+rCWdA7Xhjh4RAkWrnDgT/2yvdI61fy1K6pLRvKNzbzZi0UtN9+FDqA0W
jJHGNLnVx5VovtrAWl4yGBSA0Tm7HkKONai57bMx/9LKfcMOnZi4HIp+jvQP
j0XHQwv3ncHAfVUK8+CddRiARFVQFaMKzyQyFXo0GkD1VV3+UBol3zaYRqfS
v90IrKm+zsYfIKdyz2C53wwKQpeHQZsOw+p0f5VeIuQWD8e/0qMYIdDI3j5d
ZAjVIm5lpM2gVa8oX3Ptz/Nm/JwiyWR7Ii4Ic3yRRFGFUPuv44rrmbaec5j6
nzC0xLM8hnrhU+aFkBmAEWmEEYOFDd/+djTD0XW4zq5dem4sRAyuGybleHuO
9Mz4/KDyOzGs7KE5xumnhGt12khyPjYwk0ZLnQKY45331pNRmbuDSbkjs3pQ
6CxU8aJZjuIpyYW5Xx1W7lsgKAXZdIQ84CUE0tmglsykHGOep9wFDb1kTIZM
X/EqZGvrsXx1VZn9mfJS6FOaSP0h0hUk4oQ5paaV8M1JODT91rDgz8+G5x8F
kp2a9ttxIBAc/x05op48F1zCP6XN6LaAXQV5kwcYTnrOG1YhtVx+EY4Be0M2
uK6I2oKO7LWAkuuefUkADu+EVpjxCMlV4bpHJZToLaz1/ZKBBT1MNFSxhOs+
aZzFRRPIssU/LUk4R1OPyWacQKUu1xUCGwtsbf/1Om3J+Fnq/JvUFR44Z74R
sEXXdCoZ0DxqAo2rUKOaMYjTXkH9p2Unubjw4z55+ueUUQ9IZ1g91bjEhu26
dhxxV0O8+7N0RyfF0CovJiTnxT1vZhy7mF0Qr+v316wIuzszJ2/CnDcOcIJc
H6nt6kBxe5YKWVLfpa4sGXdhrC3ShJnVF9us19QPtnpBhYAhCTB0CPkVLfan
lEwH+n1D1Fh/91G+W5M6bPgi7xhu8WH9fbj9VF6QgoidK1Jp2kwqMiaMifbZ
0ouw/PzCyPbQNLA93V1l87+2QroKWfoC94ELcCD+XHUgGw3py6LSPD/NUgWH
JV51VdPqgjwBDC4eLbP8f91qZXN83Q6bgjE1Mr5LRmPjoxbBeDw9YEbBDPn4
Xchuse9Pg5e3WF35s4XPqLTsoLzi3JYqLh+Di1dUtXgp444ckYZ8XelOCetc
ncYHjhCDCInGnhTilMtklVYuw081i5la7MThi7dgSs+CxUoDoektBPTKBoVM
EOCtN3qkrD/zH2GFcfW2izvmTssG+ZaBXQWhFCrJjlksF0YAPriQY0ycLls5
g69lvKmN6Oqe7iwq5sC8EEEL/5yDNDVkTbPR9JreLG+2Xb3d3DS84oqD66vn
PeAW6hf2oEaI5I4hbVbBcPhwrXjwjT6Th2O6AGSN060zXvmqHE5hdi+L116u
8Kal8Kb9OesyCLmF47Duj07RLH88Zn0WaAMZO9HzBH5mRKOlyVM34WNfHA7y
0bwMvG/R/vuiEZos1MSGOINBvw/po8pq+e5L7nFtum9GHh/6h5oWv0gQGHeW
gmoIoA1f4Bk1drfdPh0xgZ5yvtX8Tp6oxg+MezHqVY/Pl3D4BfoOyuDzVBOP
K5/9O+yiulSvRXkrhZmt2wkRP4h2as9Il0MuyIbtyvXXIPs6In+MsqadgHyk
Kqd1Fd9udFy0x6EtPt8nqnQY3/dPyzslNMbDPNEZGNb2wOQiCz9XZNlXn1lX
2aPwbpLPbn/719d7pMd9UPzLrN5soGK6omaE8AK9LBmDNbQigLifXaT+fODe
i5/i/Y/IEIYczSfo7JSGus46/wjCXY8hSRppDL4tbQqj20CGSxnPfD3xQTke
6yhXnCYI7ZOBwsWY65kHYEMyXT+fm0pWXi+5q0mvRZKzAiJeH8gZNG3QkGbz
1fmGsaHfTpX8dw5EoKnxV/fMcnEAd2K+jCn8mfkyDxcLG8M4DET+QjzJoyzq
ndpldMwJ8dFpH8DAoDRVBvq4+Wg+fkC0zlLSzeJhWc/YoqDYca/x1tUFdb2G
rYNdi+6qvIB52kXG/NfasB+V8r4HHSDBILC/73XW2SPBs80OW/H0cb/lAbpy
uCK1/DDc5OZkIgrCgQgEI6Tj190wfh3TE8gnLiebLwCulwj6ojpwh62gHD1b
ckY5o/RA2n7zkrqAgy63I4M691hQvjxNHEoOZG+67ITSRBPgsbsiNgyWK0Uw
2rvU5J0Vk3zmPwPWMksbRY+PULhojSHeOGAMhTxJ2vDKPINix9d8aEJRJiH/
B34vj07Z2WpThS5oKp46CF+Xhwywh3+SfdQUMp/px//QjLDqfJnvhKXX7h5O
g2WtMRQV2Ezk5DQaxNgxF3EWZ39lI9LsOg7BpB4lN/QPd0ZqaAm5Wkxt+aoj
Uc+7/hAkgwtY4pv9CQ4ZmNpkUIjZipgh06/1tS79VSSfJAPd9VoZMHqV7FLv
0sT31eILjyeNM2iBxSFBTeCNvQ34fwJzH01nJLHPR65ZXgCoKg56ze9mBzNN
hIu29oLWVQWXRKGnBOMrcV5qiGATL2GNK8FPxkhJfLsmN6i2u555tTQiomaT
Zkrnc5WDoBMFIeXpYEypdgFo5DtbGMbDVRvuTah85AdMm165KxK4h/T/SvE0
ORYCfey7+KyXKRyAzKBgLHE5CHR8FxRezS1gGAHjumC08fmCvVa7x0s4DimM
wiVX63y9+RTTO+BVO88SlTTtS2ARqkLuRfIinXtHUtnoYGLhZ82E0EnRryT0
JOMQSaxtVGevWXRtSafP+X7PFB7N8JzdZjNDLEK4Q5i+FMiSZWODAs2aXj/B
qwL8xd4BRJSkyvBUlvUN9wjhqW9FWOz20/F6JqLGLxTxBWyIg0wt6m+QHgL8
dXqaVxhX73TSuKVCk7oNzVd5+ssYTxEBlIgW4a6UTrvZVFNIxjXm90XI+HSP
Td9P31BOy7l0MFK0nNwS5p6c/SdnyAlwe8P/9yPRAwjQXPx1wccL1X8Xzd4z
N9FRHs21Yv81umg5+WNUc/S0BqjGuuUgrf4p1S+b+vaA8kmDgDa9DqEslCEq
v5mcad5YkThKlohj+W2XqVcawyMJThuosObifWy7Aqslc2n3Y6kNwULr15wP
JIDC7vGKHmZgmdU7SQXEw4Ax8FwnlotrOGx4SFYZBydlmVw5zAGkRC0UfTtp
Td1xP/3UOzTaGw6AOKfZTlUup3cQLcvMD1r24h8Kh9gOCs+TMZP2HWqA9bX8
cMUAGbVLAB6RaphW/ktCAkv5KdK3uQaHGoK3nbUotGX0gBXaqtFwiQ2yaRWY
TCdFZF9mTgVF8u+oDQdmWRDogKWN7E6+EQ1hh/9KxGwlagW43JWCbv8/GWfd
SGhCsYxHmG9Vn5IYRQMsSJgQo1W1LUGnx2ScksQ0nU2Y2PvGolY94FF1A7XL
83xAJIH9vOd1AuXJ6P93uAiXwIPu071lO9JJMKieawVfZ1pHBO9AUwkJunaA
czbq/HHJnOAz1LR75w5ZqdaL5U38+oEzjf3w44DYr6rXLTUvPHYDY+dqHg7z
t8vyH0fOdcFV7Lg9xj+Ou7K4usONRbEzUmBLDJ4YhspdHwQpPzaPM3zClvHJ
y9B38ix973woklDcl8ISKS168ZR7pE0xcD0VWi1baWQsk5eGuVuMmB5Kbaqg
d8rdS2TZBM5GO3jjqVSrCoa3XpDC8FcPYMoo1zj+dGaVhT1utYNgUkOMW/j3
aqa3qx9jlRnN3Jtq1w03aH82Gwee4S0E0k6rmzPl9WnOQ7O5MPsmi6c8Jh7V
4QQm9S6qlaXfwhSvBhPfnRBHE/AlViDrWi4r7eYee1d0EiNWa9AsGsl5yp+m
Xr6B5j7awFZpzY8iMr6boaVr+JZuTHHqUksX33uEDIIrvMafus2KjqYgvKus
QmBs+WrUKimLxRmOAK4YH3ZFSW/vUhp8Fs0EO3Jub11PK3VCrgiib5OvWzD4
ol8y/LTaFlxGBuvYaNc9CM+0NBBrphqqJ/6OX9oAft1cwDSRmjK94+hRFALk
KMahDdGaE+mxiWSmecPYRrKaS+OkwJ6zYyCSrgSPfmWcacNYfITaFn6oiBbI
sw5rKQwNVl9oo7tlcMyJUZQKUrvfFp2gPtKm1o9rDoMwgXgPneuavkM13OBl
QoyumVd5kW8MdjAxjsK7ZJq7c/NA07NlLI/BKS07ZPcDimoW7yHM59EKVSrS
uviq/PagHG6NfR+AaL17VKEqlUgm5zUmWihFCxujynsf2PnrLlTOK4qdl3BH
oV2hjtxngqlycczjrIzT9GA13f1VpECiUibH9ODt1mRZEsrDt8cvEs0wfiKE
GK3I7hm++TYvVjQY8LatNS3AEDEjhmVq9lXULJYPrdla2It48mdpw99ekKlT
MZUOu2+ZmCR5OrzG+1f20Pcl2K1S/SnCYxWR5LSgDK4ndgXZDX77/GAsiDJa
nNAdTC+wcEyAIlVqQSgOikY1I3OYqv7vzOAJlJeznI1d2jc+xtowUtnoKiAd
TgMLxuqfEtFAoloe+VZv4gpDWwEACSMU4FfvltducBKDiw69FBwhxjteS/JV
6wz7Ry80pAuhbczgoZ4S4Kk8yKSjDtgnIdbbBuJqE045t1t8J38F8R1gjIFL
BJSEyj20jvJZshkBTGm3oGz4tI3JmpookCVF+LFVbwcXxSttjeo0TWnwoBwq
abhcb8eXXZZ/XYbZzNA94yWRRVBXE9axAS/CCEdzq9MxZcCwoBs0UOQfhAcp
wq1mOjcnrB/7+GOHPLeg90xfqvePYm6zatWFtfmjU4YqMnsK0j8VNeiX96if
JxEnLF9S6usU082+/bu9WsaEgnes47Lcj+RuLk6+/dsmb8VGCdxTPQnH85rN
GCIpz4yuAU2Wpyl4gvVAFW5udYFLoSnSA5BIn0HqJ5e601weGCKq3hCy1z1p
U1gSbXhIujIDHFESdTux1tcHYWQfKQ/ZbYz49ezxBfH59DJcsTKteodsntig
9geoirEcnrFowHPAjlCgYCX+DfwhMPVes45/TcGTSdTVFLR5yDX1FNVF3az2
83Y1G5wwC2oe6TNQ/zQGicZgwbkfwbxgsyPfsQmHHS5sEFs6H1fhJ8v640rS
qfiL+m1jEOwKPojjfVC3NCJOSy+nILwReRnYoqspI9HPTjibBDq/DZLagj3j
OirW0SCtjcf0JhfzeirnKzti0mWyio9ifWLxl+WBf1LvrwuePLdDOIbQNeU+
voH11L4W+gOqN9J60Pps9jZMGShAZ6w4S6B33gcKH/QP6ewUCAuK3LBp7UsE
9AISwebeWsb4BaHUZupB+OXpsdp6k9WyOwPI5inlG9TJbZVjGhuZdffdK89m
1capvcDqO9eLnL+CN4tIG+WXPi9miTtXR7/nDcOJ4L32VbNpwIzjv71R19GS
tA/AhQWRoIczGZJc95FMLjaAXa92rHGMLe88w4Cyi1ejG6ougCm4U7ayMKL8
8oHugfFpCRk/JUyhR+sgWT2Gu4IjU//2tA6pRUs9FbWGKY4FOv0wdUjpsfat
4UdMvw10aeoB9oiNeBQtDUieppVJDYUrRatZadWzHx/HqFOjc73dZptY2e06
F4P+odleJEG63HIbLWnGmEO10EXAW/txISIhgg+x/YX+j9cpLoKT5+2oMHMq
6RGHB3VWOgXBUSVCveSJ+Z/5YHWDYt6oQo7A1Z9G+8L6M+YIK5Q+HiihzxFL
rYVnwPdwfo54iPj41dAlCQHpoZ7gUJ4fm9PPRzH6SYwU9J6rpZrJnxrK5GK9
LACaiF/NaYSq+lBb7EMqbKT3j1WxsHGyEwjgqZJu1rV49eTW+AqUoiVK0N8I
1TMubJpuLVhGjAXUHvcMb6s7UXgHy5Tzs7DimtncDicoU2v81CMp312lWAZT
f7heMXX/lDKQGyDvbdlthNE3nzuHTsM7XQI5keSHApn3SH+0v8T8p2pheOqn
RRwxJP5AzYRv8fBeLbmb/BghYrOE+e6pwwbBa8q5ImdQ2HIExftRZw27z8mJ
RmsQDGDpqm8K5RBpPYY9FL+Ycu90yCUiOYVAuDuCQ1WSBUVDfuGo8IO69tcm
FAvdxhUR/pko8nPczSJ+0LYG1Yb4jyW70oiKKunX6a9IjZG66wQBDWvIqr9H
KbJFGVmt2zle9u+/X8/hypzmWCafyupTYyXfeW2IMu7TlqezO2CeBHMlW5sd
UzmR27joFMNUSRh3D12hsamyBWX+/LbgeIFpQAkBxYVIb0KAY9HLAdDuSgvr
dF1hnvQ47Ry7pcoxKwJSnGDW4B85A3VKj2pHDocbgOg9Y73bKexQwC185uRj
k70y7LN/RFWcdIJ7tsPwj/5JFsjBb6JLeUHtzHb4+suMQev7GuZtDcPis1Ml
vXoDYAqEbym1c7L0fVwn/LCbK/iTCB57IVoW8XJ6xHbxI+Z4vzYwEWXt5YMC
vnYY5bXUmSVjszQMfruDpbgO54VOuCZXq2lKiL5BVpV4ocuRW/rQ7q+9S7bf
KXNdwnMM6rVuAWdWQJ0P7f3RELyLYK17IeYPrPeUc4b2w/rJKw3CPNpH+nIH
MIUAAAwL5wyJ6mYXzjx/TLemXRaRLcu5eHZo05HdWgFeMorHj6xZmO15BsLT
qGNgHqUMJkE4FyPj0nE1GXotEHr8JMCJXu6jYEC2NDqVYyhFsPKaNu5Mfgq6
MWIZt6iwCnNdZu23LtZdgR0eL5ZwoxyeppgrU55Bw6EfrIQ0qYNM5TYlBzuh
oZhtv3aKVqYMRQM1sfp6SK5ra3W/QUWv/Ro0Dd9uSp9lTDX2dpqHZaVFzk50
jkrToGe99h+sOna4eA1ijKPQRFkvZu5r5HsP8Eb1Usdo+W0lISl0is8t8NnX
hgq4KkahWFvbUgSwxww8fVNkulrqMfIGuPJbdgYtdXcnt9eb9DxdikX78xLz
2a7QDQeuphROWXCnWUWJfPmPG98671DcCVZSLqj4FLhnsz5mmhK0uiAjoFct
5Zai4jOGPKXlszqj3MVb8e1u4abtU+pQBwlG3m5azcVLUiA4NCdG9TrgoYi1
BoR0NWNAFqjy+k2aUsNouLUET5Y8d0s/Rgh2koqJ5dwdBRRBjuzu/xqO54gE
V7FV52p//MKbaJ0Yf8A4oAqkLgcePrlOAb5Ms1SPLHq4WxwhidXbVJh78kZ/
pjr2aaqxwf8yz8wHJpUpkIYmZS+q0mcni5MPl9+9nEIX5L8mRefz5/zdWYXo
g2JNqyOAUM0Ahtt5U2Tf18SSOHK/l9QaUFmFe3EDcKCl8mgTfmwJKUcYVfnO
4szLLx2K6ngJ42i/3R3jbfHv/mfjCuLyxvEunesqYnpPKHirJkz7aelc/ZLN
CEOBt5xEQKm3JjgA2u2y4cWGFEbyDuL+u13UInurDnBFY9dF73tUcdYcL18F
+ATNuZ8Q9gxvTpG78zkTmP5aY6u2zei4LVDh6yx3v6QKfxIUbxnOOwxjI7u5
Cw8MHWMRmqjvwymVKpI6/sizOFlsVKA2CwLiIcrwk+1N+UQGVbLouWgVwAwn
G/xs6TsHSA79AYQ71sopu5cCXpLecTSANlT4h55JwJ2yGPI48d2ZWbii+oAd
Gl8zlxLZ7eu+rBhi8eAqdwmRsovUHxRIEUrxXx0qs2BwxEIhdqV5msCTSfv2
MwjTAZgAXbGMJ7C/FF4Bd+GzOfkENMKPjGBYxuoOJddsU2aCT+7xAPlptBek
R9rTnHGePKOGpdcCzMoZg+lXgl1aPAwfU3bO8o2/7eos/p83b4L3uEfS3OIw
zBhYBibgHjw6zLi8xStGRw7Sk4qZtB6UEFav+Z9LpwM0PKGNwvq78KCy7K9O
WT8UUo+hwMNbkw/aLNilFBzdAksVLggn7K4TWEjrciT6bbkQXIAijB+jHCKi
h27M1JRQwwqL0xZBCg+u/21GANVtUt67xGqHpNPYCWz6J7FW0UkpET2FuEaX
ZWjDz94cxb05CMNEyCB+9P8CZg1MxikinFVxh5RJX65svK4QS6bGrpC6VY1E
dBq83OGz2vLNTGCk7/O1xmOMSwE+EL/aPIRZ+VSbzRxCxXfVJHHBC5qLw5KZ
hM1DWzSpH+pE3aiVGxmC8QtR6NOzDJ3IWl4wmK3bxNvLHbgSqVwx2NErzKlP
rJDy0dw8NM7fHMD/4NxMfnWZhNPjsxD/ihOLnUzOLBHqd5Ff48DLcYA/kkGy
hPlnVzbeDI9DiXkg9WYkDQUQLV1tjG7P8yIzmyJ6Z6Ixev/M4/qS9B3mcKn0
HnaKZPeCcXVEXJ7+13CZ2Ejyzga/jo19+uyP9zvofTpGatlBbv13Afir8MaZ
8c04s3IU7Ei5xC7arP2GuEt/m5QquFHLm2CZDnURaRVMXA/2SMy37jeHV99c
bQztBFQPxYX7Q0q7u+02aG52eJ+91phqlRLhHmeWZ2wuzVNt4Rr/VyiiiKH7
g1Swnb/AiE6SeAgdHkVsjcnGPklJPHlOH5YTvonv0ch7iSUnsDfKCMR0atqs
0sU+DcyzpAG2y7Qe0QqjdgcT7QkcFiXCVSauetvX19tepIRB6KlsX48VDw2f
EM6q4j5En4Fg/21t6R8SiR5j9r3JehO6OibytHKmj8AvQ6wAhALQ7st5DmvD
nnF2UH+vZ2x9xXAQwrwhVWu16yAuOUjcFfLzqieMfGuGu9LHy1IrFxxK91Ci
JwgEL6XFjI3LVlp5l+ghuucZN7ktumb1TZMzRoEiYX+f+jIsbwjT5gFWxvL/
udna8VThT0sN0FodZutlkGpQLR/blC1CpYQvI/u1e7mvzPdJabq7xjLx+mBn
jrAZ7/7VweY5oSTUegJuSUELV4A/LGL8esE+hOGF5pQQxFHQUDz3EjAmX8Eo
PYYDhK3sxKcZ8kfzE8V7JsminY0F6mTv1Xn1jtwn+xo/i+ImHHoqaz1/SoM9
Pr0yXhsjoDH6NPuPaSM6uVcx+NQZSBtMmTtXQjVjro0C/1d2BaoiV9NvlKja
KMgawQ5Mfogcr2ivXqwRoaP7U2rRvdncTeN+JoEcVrXmo5lRrrSgl5Nki7Om
AD7RpxJ7mEorfGEk4jFSwTYLD1OkL/IW1phq8xO+mbIn1XDWWAUU4+l5+0oK
OxUeef055Y9z9JKezTcGkRFDieNa30xCBwIL144E+KqU8BlzjhUnh3+dwPWU
aFXl1Ns2/Ye+t2iLbD7wRY0j2hYI3hcQ3rBATXtBrHL9PE5Dr8zM+FxGCDYI
2ezifgThhtG9innUQDcMRtSHnWdHRFPdGI+KrnIJyeyo+G9/zpmJU8fRcwLT
S9HDwym3yWB2/SHVkiN2V3uaXwKuYvZcuKbyUtwZMbLU+urHsy6LSFnmSBDZ
0R1/+yIOSpimCI7wdDb4mk9BLCd8uykPAtcmuCx+i7fWIN/9b6k9iy3+hwgp
zQ9bIi2M2hx4YrRNqtLxgyhQqyZSRpfMrQQxyf1xCFrENBs0CoqOL1Kt2KIN
CFpAOSy0iCGaGwy2FF72DCIURBPpWYVBYaQyJv+8/IwiTs5PQCfWPrCpHR9+
n/XXW7yXZvGCTsEKsTS5HGacvrcBARkylTEqkaL5y4tMnoRW8V76sKvfzDQJ
XscVnxi8JhNZ/qL4AeV+4Vyf52JjrzJBlvp+xGz+sTNLCaqs/f2qL7G+Ffos
YTUA5PYOch8e7TyHxyjRyJK6tk8tiSmgwoe3E1wSKi4CBhFbIwuGTkUUh3Hs
g4XSKj57V6+Z0IVH38ncDfpP+/5FzwJw4osKQ08W3RNsa1QmwMwnOBAK/caG
FOWBFcUsZ6yKh/8FBpjteapFhk2J1XD+jVRPS9t+6M8f1E6ZgmCenhI1vWPh
Z3U8KPB25LBcb5XKVdAehfAmyhC4dX6Sk4rR+/wgL8jkIgnGOrcDGs9qb0EV
9w2ZIwMapKk0Ih4MeTuLJ41r5oAE51J2+GcToL5/pt1cMrCI3mMmqLpPa2kj
7RJx5g+BIAYLSNSPH1RaeQFwMt/UtDKvxDovEAa7OxOOtmeknBihtl7iUZU0
xSPLqKag4rX/BqLD7hS3XAqH4k9DbJjMnMc0SU+3HxBuiLag4+K++wT4ZW9y
vyga3duyXT3J+rjNuLHMK1kqCYSds/eojIgzCLSt6DOcBLApoEqCZndV5D54
Nxe1BqB5SJkJ28DY+YEIkvpOvkfID3yEhyJvityAGi/zI9bINKACTbAvmQOz
dfNuECArW01f/9If7Ijzo0rBRQzukUCREdpxSTp3vqWchOtg30VC7GsEVl8m
Yb4flSRd3oqpYnIVX7HPW7dfhcxvJVaJNX9EXUJ26w/iCHDT/67lqswRgE1s
iNPThC3Tkhvub//eBoD+PTvwz7vF2ETW/onatN50YF1i/vccvGLRaUxRRzEz
tovENYuLseSX4/E42iQ5ccIWAFG8rX81B+B1PAU2ZRFyr8Tm/MX1dHcFoWCR
tROpJLDogDcrH7kmqt6vmRJ/fhdwzYFIIPKZ8ICYSrmjCgbXtAtI1yq+PaDN
OQ5oVTuX4h6ninU1rtMEjqUAmi8TP4O6SCCQkPMt1ss310UHzLo+qKQRb47x
qZbL9DVEdjcuDCBjFpAeJ1FWr5Rx8yYaqBD2dIpKbZjreUeGnALD1F382Y2d
6/gxcZo9se3ygdA/QZ3JI6ZFFyB5Yc3qo2I+Vj7/S+eCLZYUyKJnltt8PfsN
WNMmKc5/7GoGErAPCdTMeAqyr3oEo++r3HeUBVo9B25Z2EnkixrIps884kb3
EvXE3DFwL7hfcFaoMRv4tre5BPkimWrVL9s+8UDQPRSIT4z/iUuOYwTG1hku
dPOzjtPYMBEmIt87ol8k6tTNolho5uW9EdtcB330qzDCXKMLmEwMWNC26VrB
uaRZpONAe4pUNygwIOZejzcDmXUD/pjhWtmm3hqGjgap6sC9cMFv0D47Wn6C
+OsvuKbbGsIPueKY0KjDHEFcuqnKT56JPRLf5HaFNdYN+632jm3SEyEEVsUJ
8a+K3W9WNdONWlzwrNtTYFnNCk7oYJZGm6FPxldMSeGUHHaNGKnVksSpsU3F
UCJVhjD1Sy0oHMXkel9/FAS0XPAM17ltcJj3OGUh08+MKJQSQKMc7YfeKAh1
gaIemhjLloZvNckJXjpk2+68Uk6gLVF+RY16gdwealyNC9gZQPwZwaQEj+KF
aA48y81aT1DHQ+683bW4h647GeTxRxWb8Tkut+PrVg8v2mXU9TL0feI4NEHR
YK2v1oS/lOF8GByDWolBOkHVE/wNlcq+BErxyJpZq3qVMkGG51vaxxh1U9y5
+blxeHuDuOLzUWJWOx139gkMuK2h9zp50leTLTdoJcPrwqMe81y7u9X+ghQX
I8no7m6lKObm2J3yIe2EnHsvoa7n1+d4k4ps8+Mq7JShhJY4m/gTTRw8b3AU
6mlspETg6iZEa9YYjyznG34Wq2qxcy/uipp9D+spBXDz0YYCzaxZvQuVWH0y
nQiW2rEERwnoydQvVXpG8wilD5xDNXdEjpmEQlqXgEnDDD36XgqMRjcMuOa3
L9BsCjBAxvurtOxbZdzWOL3ejOf84P2HtC3LBIEd6RSlSlasWmj4Qejpzrxh
+VEGtqH2yC86VNQAa6SRcyl7a/qJXRQQPaqLQURqdrToy3hFCpxsfFi5IXMu
3fCl1VY7Jdd3gr0YiHWUmGa7QcDaySZw9sgcvBhv8EBdnhcn77Ycpg4hiK6O
zx7xBiH4pDrs0bOyfaImDsx6L0LslTPmP0iCKyDDqoRVpWHeFLP782M2q/2h
vc44DgxFYtswq1Ow5SlRqIPSs0a6qhdyaXwBmid+/NoKVGG7gmg1IIsl2KkM
GVeqIjPJ3S3J9VVF4yRGx/m2lZdCz5B2CS7FY3ZuBFZN7tgyy5EA9iyTkPLx
tKcm2LNkoSXAJSsMMuiK9kJ0OCFUM5xwmkTsSmtEUhjSwJQrcKHln+8muQH/
HagyXMoFPCZA16oFJuqpiUgPScKCCUlKKC3QxkE0Xboze10BU1ZBRDFQatz5
exoKZiujgpLr7fQ4UgKE/ywB9g81ese3K19rs+5ezQADCvZD8SbaQDQ/lvch
b+I8mxwYxyggbTSp6W55uyHj8kMbNAY7eGqKTrO0gaKIOhp8GV94pjwFOT/d
JWK2oIjSkYkOiXzxf8Iq5RAmit4fyA4sO/xwYKWJOsisd46qe/tcsBml1h31
n4G0F0maEIyHVDdBWQhDOpVoKWvzAUZSXq3KWuf/XL93k8V5aP7mdaqUmVyD
QfE4d0+QniSN1yIZMVKGOX6Gq1KwArK+/9b1Qb6DiJ6PKqRcgZGRTANtuQKL
ElfLYLPlvzGJflgGZvvYAjT1yTM1LhsWu8D36+XqGl1pcX7pdubUgsoCSGrp
ul5/Ov7RNecMn3RPR4la+CDX3B8hcpi9TUjaR2jT5vNFIPBsm6zA5JTe6AEe
Ezn0P1x+WNpUM8WhKmK+5C/6/oGqvTpOyep6XuP0kaeXjuIDyn9lhQ3NLdTG
F1E7Xe0BLPK6KBxWAig58OZw2xcFymQiEL1ACs6En4xcEOLGjGYEDdifLkJO
sJb24wiMN+qx+ajPKXGBqP3+uRKelLEjRm7MB4ZcgYUoQ0BH5Ae2KO/pYh3O
h+6RiuYUcmRSXmKLShYbxQIsHQNKDrCsE9WIECr8jXdclOGrPwG+Fh6OWqnE
92JxaKKQh2CJQSXzOP8casx4hE5kZGJwv3luNfF03zMvhwQYGNB5RD5OT16Y
Br7ZTa+vKp+gUdNCiA7R4OjDpeTJsBEv/aS/y3Nx/WOVSCtT7l4escrQ6PfF
H2qmT9wTfBi23CgwhntTx91hhxog161KJo+h3YtMMNx+TwVcPfbgTYIjRDo6
nJBmPCsemMsqG57+2ingItbtuFT1ImmJe0qHiocJGAo5y+2kOAP3XU9IXvPT
8SC9BgnQ43az3EtZDo3A7Yz8qiul6Xj2ylHhWrpI6zIBgdqU1oW1afrIUeHd
u4pyPoAzQXQowarbdVVUAhZ1F3Aez9zdcQvo8AmF25Q9kxosvoyXXNMi5mZH
Rz1BdwVFJ73W1RdNcRj7mHN/u7ZKA0jQCYJxuYb285uE+OZeKs7/NG2c4mvF
Fp+h4Zv2GFyydtwruWV3vbZgbLnL7h+AbVT6uyUcPCytVkyuvNYoy3u1dAJa
Q0k2LNoHXq+NJ4awZXRITqLMtsHZzn28MhyIjsLiwq6cZTSkHhbtPMZ9qqfX
iOywtGeSc4gEzJ3HbEk6bgN49hePhAh9JnarlPsCmYKjT7VScFk59fyOHpC6
k5J9ZZUyBHoAWZFB5Vau6htap90C0ULO/+tgPVErfjraLD+IdmPde+ZLIT5n
CXmvcH7u04VkTR9bljiReHsAvRYYxuSy5+OHk79jYTx15aMNpJeuigsjthCN
t+14MN0OtyVLKQUXH6KFTaaqnAV5RgAeC8BJUiOsZYOKFWGIoFkOKXwfWAc3
pqA2H6e23oBt8YU2LKXmonbI05qey35jUbTBeR7zGTQLe/lL1a2IQMeqAquY
7E6bdntSHDS1Ep09m99YiVK7fej7yy/ODiGfisz6j5tpkDRNsG2iZHL3TR6Z
0/MALlhsz20usU85yurmSJ912YxTxO5IUAPDbWu2gXxNtluXstbO7bIjD0vw
M95svlp7Y5qiT8CGsRTd0oaHBpBuS2rfdtTF2RrYP4NNHNvWL50t4VdzFZfG
Fzn+iip0CKIRv9SixgayWpeU+X+E6X/YWW5VR9nQMZNa1x2vf7nrS0kngXIL
eReVLAGuZWDPlFQkDnXc2bpNygk18hGzS0cxxG8QL7VJjAAWoN/Wf6hiXmSG
T3o7t5iO4HDdOxu/673UxgQerAU7fE5HnfkMCn4Iz0jb+KDxqCe8rZ/h4nxx
zeG6fu1cd0HriWxq9wI3y32MUqrWYysMldscErWiHOW79t/BF9HQ+GChkD9/
HJOJ9zzLNd73QRFKi+Pr6rqPzZALACYNgcHI1VL+39evH2CTsxdWbGMN1Ntm
6MbpvLvhX3BNRrWhl95WjUC/vGWcOdZPKb9pIvipCZyMyaLbLQU66n6XiQqg
jZkgYCsG+4glRhZbJl+pSqDc4BLeZb1QUsGM5VBIlasdaHSYx1eCnv5YDW7T
+C+Jbfk9OMH8tTC0YBvqbiYcZxpfEv1sLOBSv3n26XM0pS2p0iFZxQKBX2H6
KKBqUZz3tmoiZUPI6yxkneH4KUxo2Ya6bI0gwDTv/gCHz5vCyCfvE0Ysaf1I
7HLE5PU0FhKvAWtQmkeSXacXdHrkSSphpTeYbom7DLd62g7n8jgj4eN5RZFg
2SOkMLtEsybmUxv/+w22MoHVqlevx1yoOPUrvUTAJlAaWvNLv11oHhPl+jBa
aXmR4xqsy3dYSPkdAztj/Jn8+bqISb2B+isND7QWofDkHyPuinH/M/rgOIpl
ohejkecju83Fd+efP00HVklMohcsTfI3nBOofrXrrxHIuT1tpwaU/kkT2kPw
ypehyKQCFskYhEUe+w7Z2MMefyaBXOTX5w1wUP1UPQ866wKSnDk+lyCNuFYk
RLqSLSPnC0POekNpyV5Oce3A/ZdNT5QcSIFUrHVoWAsutJPHdwt7RbuWygXE
KBcj9pZ0P/KD9mrYP/GMfwY+362DkfhuQrqFWVfpnqJrs/tFhMu1opm0Ccyk
8w2Yq3gB3dej6A/19o0b2vUARoY/dPiCLQLv08gTQjqHNpuw/9PTW8wwlAiP
c58fUiS+fyRUp4xRaL3vvuMYhLJaYie5pb8zilaCVTV/6XEplJyi6HJtgUOT
cYzjAJfS/E1ZdUw4+wpY5udLb9lARq/oi9YbGVuMDYcKUXKpRbz+uK5eSmgl
ZQpD8P43sE8ZgiiOwuBt1JjPdEoCUDA2QhW5MWTbHyrA2dBNewRCTqbhkdYj
ICFN4LgyVBKT7KAE3rZPdIvMMBmNkwGhdyIeyjmUDdYBGIVdVtPlJ+WMhXkl
r8OBzFxDgBnh4n5bkwnVxAAp5+h6LrCH3nwOxfNpYc1Q1fYRlqNxowr3t0/4
Ge6Ue5CXUFsPhAegI3efP8Dj/EZ6vJG9UNRNzNhUPvn86E1g2nfVfWR3/kkK
UVzyCotPmySD1gUfo1RAgfXrBAEFvwUo5H7X4tcSfCFsNgpLcwMaHRVtdRFb
a9lfRhRdu9xbPVvXxCYAuy5NfEui36gOnOXA9z4aU27PexyJzxWITx227C0e
f7kieCfefaWAKuAEXVzWLhRmcJGeh0E6Cois/lsclMvpMVIGBohM+akDlno0
noeSPLx6VI1VNButHs975Dui+XHeZAVcomw4WRyziKuFzaV8reB/IsiXA7IV
CZqn2I34+Br2Vl1/M+3iZNn7GjWaPuRyetgkjVkuA2T1RVWT67O71ZEnKpyX
0OWiT0AYxqkJESI9DFV8jExk2PselA8R1QY+n0rBXImhmJbyMyNASTmJ2xyi
gV3NSNhJzRFdmMOqZ30465bfDtwGrypxKyL5uQfbdHck+SlWxoDhZg/KoJJy
u02Mqnca+r+k5+kxejYdwXgW15O+jqwhETcvSjTHBEkCLhPEwpyxcn5WSvi7
ugBRwABLEj0+vaHiMwO3EGl8spbdm5gtB3aTV9FfKMXYVeSr5LA8tcVP1jDD
eLk5Hdhfr0ZtiDUYN+yWPFy4JPAHPBzjy965vqyA3e8az5YW6nPRf+rec5ON
3dQJfBTPE9/j2s9lMAe+87d6Yga3p4FFpWc2hlUdnLW1IIrM7cqsSKwfXvua
u5ctIisaIHWkBDHkjq59kUKpm5BHQ71EEC+9oWVMO2THD29NVq8NvUVs1A9F
gDsvLYBseeIMW0Mwh77hbFui/KKbi41FEfA6IH/Gc1+T4+A0Tp71eMt9MEJE
cq2HOwzatOBMV8MDHuyS3LKxc2I1dhxPK3AbV2osxBPVFimGcqIQp0iORpp3
O7kOj/dcSawF0gzOxFGQQv5BEVl2xNsrjwGRpkhBizgRZA+cFC0QvxaY0F4T
Dy/MeOBfY9d+URmB6vmYNTqNlpJ7H0RYapRaWjHdSWPK3wr47y752/o5u0Yn
VEteL9LXjRJDLsh47OyYuuGqF5iofVDOKYhKKdDIO8GtXeFuCWxf1aXmUBb5
8+KkObcpxD0qxwdEkmXcYnUoLAYMT6fwo2fVdMSd0l6B4dGyAX7ZypR3m+r7
vjOGs+a487xnib9cIbejZNG+PDO7o3EZ3RhLSWu+p4tEh8V/tVbDKdCaZuky
eWVChINQGzE6yZayQCMzrfiUrZ8lk2wlQ2f3ViU1+Dd6U/ZXYMQr5/IAi7md
PrHx97ufLTranYKV0XjwvmXvov1tABFXu9moR9ys/4aDXHGmu/5K8d9Ofvk5
Z8leWiKBCUJjfPS32Bgf6FCLAPBP2Z3Y3e5R2kv8iGQoVIP9gjXd2SIviZcp
ih+DjqLN2ScRFOYD1jH1KPuIbE+Cs6SHr4/l5n5INCu5q8QlsV/l42H8qCkV
9/TZIYTAaJLrQfzuExtbN1Mes5YzicpbVnDoChXioHhcSwlWkdZjJX+qvwAq
9fsoe8C2MlucClZIZ54LYJawnnWw+QVkHCQA1OME86Ek+g6cQGj/fayQ0JmS
MX5VZVtiz/Q0Db7xgWFsZnE9MsL34dHJkI2/EU/8sNfVIwo5CUJn1uQ8jbEO
K2brIYUQ41fZgJwgwyfzzk9dX8zsOGT9l9Z/GwgQtHCq729xVKDqT9GxdTms
l5bu0ynFYyMNXMrs9A65xbkv6zsZiT3fp0YyH82brBYmdwbquaDgMYGzJEk5
3j2RunuhEEzw20oGUTsoCMls/bRkl4ZuvybdJri2jUfCKeYbznR/fT5uJFg4
WmcQ3JE/spezN6blYYI3OKvDD1xBa2kxHTM25p7RJn6MFlPt3LSYY1xrMkA1
OfZoqsCS4z1agEKbq3TPpZ3A5ax6sLPpRLUDsQ96uFmxkQecIgk0mT7defEO
ZydEFjf2Qun/s8vzngQJspDKqrmyc8Flcx9wGVkJA8s1+EF0TviXBzjwCrXW
2jJqMe2jBzEGG9sp5ghMp1YDVa2RNlJ5z3H71XpOcmPJMrkfMuCv51ZRv3lg
txcJIqddTkyEFFE7gJZEC+CekI7PVYjujQFXBzoedL6KDKxnJML5uGsjj035
fc1LZof1J7cdEhmYRKv+JDN+V7o9x+E2Un42paQ4xBllRvtRpBeg91JeAyrL
x3xi6XuCM7qzdnAsDjJcbFSMSiclZNkiItklZ4QP9OtOQ6ArZng7bNNs1VZu
HFN8k9MJhsB4bwDEcWuseICtqmPlIPX2GSAJqMrL4Pqmx9Bf9makgPPc+Yf3
98OSZLWKjSDgn6Lyt3wYwWuPjREmIYdaPUPNuSHxtEe2GoYCZb2eOogTbNHK
cuQiZGsMwR7kEZkuKnAzdJBpu0+cXermeWhPrL6JXlVhiTl+Ioxn9fwzsPcA
8/c30xqUiqXcD0ZOVpSUH1mhnC2qTQmsHSf9INp9qQayiarqE50coPyL97YU
GiStilLqICiFy1Ra7xUsKdoWxR+6ZKfej6XGycQogfZosyEBpdaIrgZovD9V
eChOEIg2umI/aPLMFYTpQ3dB9XUXbtP6m4SsgUGzVrfrgLU0bkc+PXmvBtiX
WjVhVulOioy9RsWunRcChOdLnxyGYYsIWEO3FlEHCMVgmpSxxHILIoGK501Z
j996WPuLKRWWsoQqHeSQoFAd+a/7TIpMf4YA51l3+oQEU93hAxj6FgctsQiW
EX7QAn7OWWJvQP0DI+QrLJ6dmZ0Itbbini2D2CxVu17QfRIl7NypMKc2BKBm
pW4oyCOogFVRd1ypNR6HQDPXElAx9FU7wkX1GxcaMNjZT5IrIpezoTgy1aEL
+Qr9aQJWAN8fWrrPr0HEa+qu7dqrca8Y9FRG7bZWcwXr3h2XEHGv1C3SI+Ur
KPT3elA6p54kA5p73AeVfyY4y/85+yuPB7CelujmE2fYqYHvLuu7eviBK1Ku
YheO//hrFcuk0BWGX3nhnG7c089Yx22voAHs7eIbbwvVigAn+7c/iNekwBjz
GDls1JNtC9E+3/ujnWmACdak1BGCiHSfFCg5WZ4LO5fPlBzUBydRjt8jzKc4
/PBvHJ69oqqTPerEU7ZomcZzwhv3Rh/GtwSJHquuiJ8E7trZ3iSiAwpiFHoL
J+mTF6Pb5flX23MT0rH3HM9o6PS0HzH8tVx+Fel640VkvH++5IeGR7dg6LNC
FM9bAPjWXrZjit6Cou482wOUCDwHbpEJtxrkIKXpEJ98bBRInyfiYL7WN48i
axADCfCfGXnxElUkVTZ9c6H07i31ZbcMG/9etanq1nB8mNbdbJo23kb4mfIS
RS7QyD56GG2uODda+rLUghNULbiCozunm/WqC612a8rxtw2jkH+KHtaCL8MC
uJKNk6OHSqrM+g7CO6+jO0YDVqIVCKmyRcPSrOt2e4a5rHVfG8C+OYwkroAu
X1Ez4Ru+PURjgrE6ng/5PAyzeLrQb7PwdKutBfFMdFegJOB/wO/jhr2zz6eH
WjcHAtK3rNUqgdOdqrij7j6XF6NJq9f5quAQQTkUti8P5aOMb/RWtk1dgIaK
WxPim8+Zfk1/TGoE8jTo+tlypO1QSqxtNynESb4cWOGMs5vayZ84ck/uGQDl
owW2yFP2h+/gsNzSRXqg2A1oIdl/hi2l+w8GoMJtMZDt1SlSVBf+DvhLF6Sr
fcTXY3vMvmfUh5auMUWtXODLgbLfWHB3LZOpQSngXscXJCWCEimTNYpPPbdY
izV6iIPAnZh+IOdHwm2QObTwkCZJJfDoFmMG+tTojH9/UY0Wv0CT8RhfL4n0
3onI9Gg59jlW59vO68A+Ok7kAQ0AwRB9qHnaU1psq20FU6tYdl2LXz+nKAAZ
9oOuQk/8aqyfcVO19B1COs/JaIJnsKvuafYMl4EBdlENPgBkF0K/55LeRmqx
x3uKn5SSranrCMLdvi53E11FMy0JsI43Xum4Qve19pjZ1lmUfosKU6uOsV4w
sxGS6dFSUJTay9uoRhJACpjCvtkdjiBpnsS/OSC7MhgGsmmXVAfZWsoorPHb
UJgYtkmvtl/o18enCcParhKUHQC/jiuyYCU9siRgbpBV+1ppH6cwuUqnKeyy
rNylwutQoC7KPr1qRD5laxNX8MPej2sOR3vHtwERjL1FFTE3LtgcEu5Jvfto
Brf/DpTDW5X+BNKEj+fZxzPOSFZC3XriP9yi4nt7mjk+zUTkPctywlar0s5b
r9WJRBi+aBZ9tk07KJK/EFgNEZRFhcz7gfdc8zl+0mBdeC/mRpfWNgaaYO/o
PnSe63h76VgbPk03sCBlM5jVp6lI9m1eNNIBYWpMZFRY6eFlE6TsB3KZp/Or
5bZjQL+VMgCZXw32BM5Lyylq+jNPNRdXqbgGSZyUQs7ynux8BfkIY6Bekp1B
tKFgRo6yHeGggeI73lgX6n/iOux5wOv/2y7ZIwqpO7YpKrKen2P+Vj/HKBSH
BtthO3jEu3eu2yIahkbWimCfpecFTvfIGwy0ehD4SGpKVGlxknfgIC6wP9n3
wFQnA+kxPzZJlxHLQ+e4gKFjATyQ/57+3oPtskCR7ckhZVDWZJT3nxD4L6YY
Z+7PdZvMer/i5PIPmAjhkBE1EwSCsItbLdCYeGTRh826d3r0AWIf5Ul6Uhdr
aO6UCoeToml7Mae3Yiu3iQ3dwvwFb0mloMu9ILWorsn2EH5LLXCJzXfCKH4Y
DUGW1I0UKcbAvoI8SUqyccdAaxw86Bb52S+gMRbHhrxGh/JIygoWn8GYIyHX
BSctlBHpKMQYWg9P7ubgm1Gyvn/OaLWwvHjz8nNPdqc6CKof04SqTa7b8VQb
COuMWTRGsoOHNvGmqkxj6wKuTxGDHMrQTN4by/rb+pmn5l3mOXRokWx5WXG+
4xc6t04UpDOLCN8ENlR9GjJT10aFMNf8hSnKWB5Q6AkZA62VdeYYZiK6NeTW
kcqQ8B7S8zqD7Uo9qcs1Bzz1IimHehoYUEk1KVMGED+SlSqPIFa3VNmlmq0X
RS0YmdoMKRP9vAR4bSJvTJIpPKFStjyQpRKkDMZrzsGxkn/gDRxr03NTBOU1
Zrrt+H25K4y/hCku5/2sWZjFWbE8Hpx+yG076YHzOSSpzmK+4FPSlDPY49uH
13Ho09RuLtb0kPCtGgnMBxvrgMUN1ZrCTtdfOvFko7LxwAZzOHGeeHC+AElW
6qQbX+R4kRaBjuBKwBqPL6HVYZsL6Px2rsWjk9m1+rOwynOpJbrRbV4Ci1k4
0l0sI4LDemUyGkN943yEG1ov62L3W9fjHEYruHrhzZoDst3IuAfiUDDwYJXW
bdTOK/zQMMpZd6ArP0jp0yH6xmoMZgKRI4UTU71ZPA/T+KA72M5NxVAx3vJh
1/t/S5Bqg+tWgJaxJdXOjU+9GNCIuXR8yAkPbKQEV0513Tq89T5Fh3eMOsmt
aq1BecjRu1NSGePWgzYlfbCjU+b97eWLInJsLiSy+nxpk0Z5pgRMs3dH587O
KnHiwRP0/LKzqRs3krP2MTmD14CHP2IHdVGdfdxdnMrtAIu/M//atj80TbY5
2djLnkqq6ot7ygLZ58L2AYzImMHOeozSnbubDwf/heqcU9PUz1uVsbQ/Anw2
qLoB8cP6oevn3NBklQEeEhYVR3dovRZLQ0BdMMKFBVYqVfpAjSTPzNBfi8kr
t5AAgTEcbBY8f+v0XUFGGRxrV1nfL1UH+SYb5y0fNq6EAvrYg4k3aGWExDKg
d7zObcoSAdnzlW1c6f3TmzEQ9pAmQ+x8UdQH5URT6aEaOKBJxXkyuQ9mhoHw
cmY6hRHPxPPCjCTHWjTe/M0RpQ8D2I4vXIjMUd19SMHCALy15p/BkFhbFv6g
+bH6Z3b6B+yyKb8zo+1eTmz/zOmyQOTd5wbVzja3M8uVUkGR/f6LSr7fjyh1
y7UXQT7ah9gMjqyZ/yd2qXIanLeUqLqJJdhJn2y23Fik3MiJZVVNr8OZQi78
XuSdAVn0fetJHtMZBI66rVn1GINtlruI764RbAdljgLK1Zis0O0U09S6TMEK
XrvmTHHJ7+cnNEfZjBjZboM154iECo2Ni503Go6xot+C54/jVbBMkdsnW7rp
/I8y+fH4lfgHOWUtzxeHlD6p4/SCD/LWbecmIK0EJ8LIKUYlsQpOihyLgTOS
KhTdtAY8p4PndylmcwLpA5v8JbEMDj+NjrGqASHbZL9wrxxd6kJrVL+K6Z9Z
WZl0NlKC2ZE8xj7BaofB/6O8PHEV2QPXCnbJDmC7AU7CKf1gNQ8VGW6zzXnm
yzlXApG3O30yZqKOhgL+WiyIXfcLimAmdd3LSXs1Q/BNVu+hdQ6oygp6dXkl
OkWE+uniOaFQBfTWcKPx+l+WER/10nhN6Mp7XWOxls13xKnUpIVIrJM5i7Jb
HPWTx9ylw0wf9jelX7fVPK7zjeN46rIPjiB/8u15pI5aV05tTHe9R7/mfQZ9
sNBrdNCiomT/yugQnJe8WRd3vikT2qzOMjlT8ed505cLx/Ub74P1JOzTOzKt
T+CkRlmO7YFVEB5rvbd310LWQ3mKPj1twfEGE3artDIa2H1mLyq/lo0GSc/4
XN7nc1yOfZq2SIntA67z/WI46UkeiWMLvrpqR7B5dgbsbN5qQwcZQoWTpzpe
jJhRgON48mukpmVZ9MwUpiaT6+xMAIkeOGbYN5mIxiloHUP9T3X7GdqIp2bX
psNpk6wsC0wMF6+LUnT2RGpRKqerxDyHw//N+6DtMyyda3tlTf6Vvy88o45+
YxxxTOb6HwPuRzd21plOrr7WhmvZMmCaNnml4n+0NsHXhp36phEGtH3lMmOi
26qKuxfkY5YNcrXInNEv9FUtKa7R4LkWbo8xGYgPZ211+Q2zO0CUW3PAjqhh
i0OI7bo9SgAsj3MXhj18WnC1IrxUEvcR9JcBs4wETNKSNDMWTmvlBFEHGf81
7FG/dJds6vCSVijJKnmqZPsIYm5iIhJllQZGSbt40a3wxROUb3OX4H62DnYF
fEnNHgvTcMuqA86ZHGb9cUAfMVNPGZEbeMnykdTnT6rRI2iyVSBJqcvNMGFU
wLG29wrAgjaNDAzaYTg/vCmhVB5aEkLkhqYJitGBHCmcDp+W865Sn6rgAs71
sY9wc1mUMYdppxgYwRozTp/hc4exHQjfX2lRIGVsEXbXg/quk9zpFtyOfELO
OGxx2DV97K64XeIdwHL5RTh05QgtojmOwDAdNAz5bKJA+Xy4owyN3kHL0ViE
mFob5m5EKdbPWeNBMOypyqPsotqldgcsc2SvA2Wy76FPNUEtsyz9csJDiK0r
VqeAeBNAV85TxlyiHlpzWn+feIImV2Q51N94+6V1zJn5ejh/SV/uWAZzbn9R
zwA8MI7eKlFo6uoT5leyL5gbcuoVhd8oYxHB2qihh9sw3wuZDs+dJ56BS0kZ
TzVrpflDS2mvTibQMOPm3CrthOfI5AOgRapaiBzF3kcTPpK9OBg2MeR/z83n
DTb3JDZvlNneGiBZuiG7z1PM8zveQ3ncPTlO3D+YcDHiiPaw5uawfU49xGqd
d7GQQrmTpxopxk9qKKy1IqeN3jT1i0TbOPQwsOX0Fkvyts6hdaTDLZygWV5d
W01qjzej8dbAo7x6HAeg1necXNmxxpyoYx812aT+NHxGNOsBMSuHLW1s0f7s
tJEo0P46bGk4JoPQfgrItt5iBu4huDeRpApKPpVFWSUvCVvRK4jx1c01fFit
O5Ui8KbJ36S/1IQ3hlFbOF/bmPBnZfJUXmAPR/rJrcxESLtVr/ORjsEzC32I
kFO2ok2oPJPMfiYyTKGyz64HMSAAhnzOSe+nQJ7jLy03xH1igLzFJ3KezhM/
oHbElLRqkL6ThaUPUrYkohtFy5Jg82Wrt+tD1SNw6T3m7WbHpOgxOi7cFdty
zmphR1YbMLbf+GH2QFGlmg6tAaXMSY1djwdMo7zIKUKpWuvhVnA77vpcj5wj
KxOdfWLFED6/GF/I9XdAC3tsNxMG/EgDwMHCo0bYJhnXWL0Ou+h2KUrAwN7x
ITDrnln1iOO+ZvOpKGB/qyjbsOPnlmCLxH+DxiONEDalDNZeP1hROlkrUeFl
9+xhBtPjF04LFiwJox/XKB5RkRvi08m1uJhT/40HQYkOEcpRR7mPAMUxrsiH
HvnlGGjV2MCnuNqO93hD11docTvOnoB1zFAOORGv2ih5hSdjj9MxgXuCVR7l
flo+vs9jYsD0MJMR7K80xnXEz1vadBiET4iD0NsY5jpx1KVtWe5O2dSmm/bX
dc6Se3Py+UN6ojS9/o0N4JGg7u50ZivrnxI6iFNNLn49lPH8QQnQth1HERGx
2Pk+YX8pSs0FCo1zpeAVxe7KOMxeIRkdFhE6iXIndSfWcBYwyQcjc9zCZ87e
yOelaP/OqCre9xhgL0tDvoj4At7juNo+dbbSdfh2LoD21AaFyFTZPCwUV75L
Rr78Yt5j8HpfG7eqxeH6PelZnSGbIkUSba6BFrl8rn/5R38wdF8t7s/WwFOW
qm3NgNkgrWZG3U/amtfr7j/dbX+wix7pPcHpHTXknWXhrPitfOEvGgpUaHlF
L4K9wHrBTNxjyjKOnVzWH470pK2e2TswW6KAMOpEUfsKbjve3mIXI60kihnp
caAb3xl1xEMSmZm5gp5dg3M9r/167O5XLO3UJWkB43fAyIXxNIQGvh7DP4Dc
+er+UxfMkSMjr1HrpTMrimWVDD5KL68JiPcxybdwXud8emLXsKAG/x91gfOr
6ln9McFHro0EGJISIrmWxUDpderEmP0xLcvNV/dKY6taoGoWiZuvA2VLF8xS
R/3rGnfSF+D83JDFesJWtYBIjR1BnYmtwyKPT0zIwxXX+CESt4f+nKQIdXEp
npa5aCbuXii8rqvNW9klijCfxlUtlFtjp6wxndBvn53x0KQe7ylcgYB2hmDk
dHVhT38pQ5mwikxzw7YqTj/dt+A6bKK3422sTG0PAQJ6O3+Keq9ClGKbG9kz
2MFkCTWuDduY7sk27fSoY6Ny6TLwTa+oajFNWHUT21pVspRNpQO5DREZXx+0
hPNLyVwYhvg/cMRhUbXEIrPoCGS1TAow+krFn7l/u9u6S9gVXjlAZwrRCFkM
GwkDYff407GtYk2lV/mA0AkJEYcmA8xp/dTd272kOUMH+Yo5YeXGW0tfVFy8
DCIlm9ydu0yY6zYUpno90qx7Dvsfrs7s/eZjP28iiskBGuzMlNPNExIViwBc
K9TO4F3w7/7NEjLD4e5pL+Beno8blkDIDUz6H/5tPOdBqCBMi/TcwhJHTJB2
hofcnatIDnwLXWiFAE7eqhP3vBgP8WL2Vsup5cR+hHDc5hhsoSMPFqI3cdt1
HtDzf8tYEL6Ddl2gQKmkjOsBwWRDPiJAV8vO12lxjFCTW1Z7tfw/0bIt41be
3BQdd90vjSBa6ZjI1CDwt/YlU9VSvlpQHfeNjUWf6nGkWm05T3DLG6nd0EMC
ZZDnHXxz4/LZR5KV/NDkpXYnJRy6cMruKoH8iJoeOngl8eZYQmmO3cgzhS2Q
Q2gepjp5swOTOFw8M040XpZK9vY75f4iz7mNQ4zszfs1cDBUL6atlz0dzdUD
9I69dxjmo7UTwd6Y05OFjzMrJTG4ACUCy9pmlQk0jrz7Whi2YjHh90+lcRh1
xnklxV6k+dSad7bVnZpU4Kmtc77H/ztgdSrO4zn2fW2AG9yvFg4GzH+mnMeH
0peV3xAhWm0C5Il9NhLpel5d8WB0VtcST8ePOwf1yFgx7WKgwPTik5IQc9ar
UnEqM3/udQRntnAZ69HYZvM1nJIkF3iGT49te+9sk6LxvLui5zuhnJ3LAuIO
etJdOfABKNxEgr1XU05Ya6toE4nuKV1aX7a6cgfzXKNCvhJ8+BKIog8q4tQi
yz/i5lS9KNbOuQ/i/aLvAXdOhiAduOdrvD7jPuAoWC7fNGvjtCpNnd0pmDCy
T+gpT9su4Jrz9e9rNhqv3465FpbGaQqbptnwPXaYVVXCfeHutZU414cnZBsp
ekOdFiWkH/4+5BfEusZLmFM8Khh+BF2NZEOjmN2oUw6hMS0FbY4K9bCawJvU
2m/gWuS2xCnSW5D9xKVIBiD20CLJUxdrbGrGI7SmFHgP8m4aVQGGgjdeFHXE
ZvV0Hao+yMwpINo1IF7amF837SVUdL4Jxgb8pC0gviCpu9VOBjuQ9ZjFjRJb
VUjg+Xt5+ua92q1MneHGcDFrb6hgsFt2m+NRVoIhV2mARtdhd1MQCHVXCAFu
7XwXWgOasFXEdCEqgWK6m/SNVoGxewO1WCjdnBhL5X1NJwBUL2qx2112CSAO
DMb0ErJp2y5H4iS0omrwEtdjyaJiCd/z7czfxJRATrHjd767kXhahCqma55n
dfJkrWfkcUI+ClK2WWZG+n1JL8ouzBsCK6yMyEYG0WAJ0+MvOYU8cNW9wrGI
C6FXbJz9DZaYa46DFkF+rFdDdNclCRp3J3L/7emeFm6GehiGqLLOjGtIzpoD
dDhwL0QdUVCqi4ddFRdwmyXPBhe2VtRxcMfPMVUMGOvmI4QUssuPF9Qs8meD
6kijpYrjvF4KmRQZKZ6zayevHXCEerYEFGqEA02FHolQkVy8ND/ltUci5Gwq
uk6QNrqdZ8tk6Q1FF9YDG7fONwNYBQj0CoDWjGWwY7xEnNZq0/1c/8XSrtLr
Ul/CUiQbQvwEhDTgRCBSBDGOA2rSQ6h+ndJZb0Hm+AwGRiFtrO/slVMexYNT
R4Blxq0u7+ZKISACVdDF618Eqc/QMrzPm+JN/jkpX0xluErcJC5RNthtRjcg
SCGJvETZdj1GdB0VyT3mgTfCr9SZAcNCkyx9zgeKcdDNjZo1AlA1UCwXu0yN
55JOivF9tHgh/InXkj6xTi5NL1svMtthWyUHvKES9FqQfN9zIQS4KmEEvxDy
Y5ts1I7SRWY567jUEuYeWeKQm0T1rPnE2RZmkhMKA6K1cY3AZJM7t4m9Jb3r
rA2UirSgwbtsBpv/C2t8jUdq0q71uM2DKmf445JnnBs7eelZnuq/Ym4CB1Hl
5COx9JIKiZ+hU8g7W/5wn9v4ISkvAU3eTcI6YJtQtsXYd7fXZ4mIx3r5lKrf
0bH+P7gXAPxniolAaP7L+/J0J7mzLpP/xG45DJd/EHI6y2QnJTMfAH08j2N0
TPDdmyTeYWk2AkETbmryH/fa98vmiz/6RNYipu6USdj4szUXRuwQHvHNh/nu
9Chw5JntbL4U9BIzPWaCNDBU93Xs2Ov+KXkjVinS+PcIstcMOyaTaCVAJNDb
8bDsQFALKF9RHGOAUeDptAylvKpH0ORArBvUjJyT9+Dij9uU0UBJMdJJzWiq
u05yD1KtOhvWn68cXiMtHUTwyRupMCudYbRW8JCxkyna5sE01vVneA+6P50A
t7ZjShdAPH+zzBIMcHLMOamKEjMgR5Y833azL7e3z/5rkgHgfa4EKc+C1tFu
dCmWCUaMA86jjizzbS9Wsh7oytt463NIjB5SnXDczBqZagZSh92ruCTnehjX
76T5wYdd0Fd4E+NyAg0OGS70xZR0UsCpCDlSZWbbQ5jQiOsl5/BfCnjwl54s
kokuCJMhiKi3M/Vty/7i+43P1sQBs5EuMu9+pNQi2hWdBLIWlXx4aYr1U0LT
gp3s9rWwsEDWEWq8ryQQeV2mB0mxMZwZxK6rLEWtHCzwQ4uEutrKy+MkbrfD
ksH0hNU4u6uOfet93DQQef/lkXlKofLnhGwfHEAdoydealLGAnFV4ZLT5COo
0YjreWxF3sUmcILTqVvzT2DdfjGneRmPitnRCuheXLpgne8TGgWkqUlCUDYg
gXhmOdnnBgKP4+S/6aioS8WNuOfTYBeLQIP+nnTw8aNZMw+/Zi1cawGBE7mu
bfrmnlSbCozltXvzTTKOU9KdscKro7byPnICf4gd2H93e8590kMA8rywgHys
XjSdx7DvCY+mfP6CmDvDE+j9qchsQ3TU1SBGGDL39k6hVSXZAhagj8vn6+xG
SoEs2QBGQTL0Q5fh5x0MqUW5+DJNuApe3P/0RjYYbwQWwMJCpz3NrlJK9tyh
6a1RkUfgLaDk29tuOj0sUZH56ReLvwg2vrMCxzMKwxpJW3bAd0a0WeSmtvFe
Ymbdprv6rJc1z/aTcwyWcgElFbxQEOzzqLcBcGTEHjVs/2jSwZog1qyd6WRX
QoiV8N0HT7RXbLzlsugqCjDIeqMRbrFhAhayHJboTntVmZ0vBmvNlqkpYcdM
04kM6/82o80ArvrM7vueveAv87tbOxRtQmrcgDN7ZLIMaphAAtEwHYjG/j31
vZwPovUHnhSPUk98J7AszVd/f+g8mWJrePyw7+kPaiS0F/P9RzpoN2Dvh6di
eR+FoRC16spq5tiPt0vV3XyW+Y4jXN4YNZ5vBwRKnGFNBLvDNMxcJ6W/MaBM
HwRM1L2NmkQMJkx8aRQ9e3yUN7keVlMKVqreUrRjMgiTeO4AMaaMFcbc4BlP
Y9HIRW4XL1nyiF3VjntV7KKafCxxyRviQlwupitDVI3Egpn4hrHfSijpn9xV
t1QfxlamUUAo97B/OZ5bev1BtXihic0llaZ62xJ735pGLtH8HaATYr86x3W5
XOFJ9/mmnP9PZdB03c8tN5Lqot6p+uuSYZ0FryqDyL7PpFnyJpGdo3uwJCXg
zwGA1s4yBaAEjuccT2jbWq4HgAqaY+WZ1XYZXz0RB/uHbqQj1vUen1ug5bPM
+x6T5t9zo/40OvgIIdHoFgnTBp7DYKap9IV/KMf878HN0iliRj9FRLCTz40v
y3eGNx2nB+S350ORele73W0Dyh+IN9/NKz2p+cR5fFS0+3meXMOcK8WutH/f
VfOQMqAdrkan1cQX6q9SpRN1q5HQP3gkYe2TTSb68uADaw4jt2oVdohvSbx4
xjY1XHv/p6W5PT7QzV7eXwk3yOW1Nch/wIH0N9RnFM2m2/lm4ZPX/i8AQUI2
vzJccvPqdIfSWH9iIlfhANkpeZjDGrXUEtDVW9IrMAEhYcWfuGoBZ5z1m+oS
z3RywBpVY7VkeS84/SzP1xmL3mqkgGeFOoxYcS+j+YOqjZ+IF1IUn6PpU2l0
12WHg4t5V7GUTSjKSglJ1XKNIXcWm+SB8CY8SmJAiYgNaayq4ASICQXkohn0
RpS6MonFUpELA6Lx2x5AG9utLqirYItITZ+zGQxaoJ3h4hr2IfyILlJz6RUv
DUUCCTkvpHwDST/ON3piDiOfqLkcI3bWVLu6q8FmuiJ3CzlVkWjPkhDK0WS4
wk0ADule5RgyWyGEpfukRpK/iD+z5tSog97IcYyPDPcyOwgftjgOrlTQry1L
mezlsfpvYo9bMFbvpp4ffKwrdHl3p6PJtQ+sEcNaK/ay86RJrl/wAihwkg4u
kITl3hqz215WauzT2uEYKBoU9uLC7+Zsw5pKNZ1W/Y2kgUQYs0IIy2vA7ChS
ki+75IiXWQJXYLf8jNO89hPFbAsIgXMOyehc+ZGM/Zi1AeeXUM4xqFubW+Dc
9y0yVqSiOE/bBj2M1LNFKCJIxL1sy/UCRRb6+VhXSNcFjkqvSEmv9cev1bpc
jlg196/4xmY5QQD8w3p6ciWkLXNvLqwkNj7JTgxAd1eQYRQQonAWXHt7k2t/
U5WB/olonyS6J2CyTFthmEOW1R7QuD5aOXsTnuLq0I5IOcx2K9nqutdRVfua
A/QXIth92Y6VmiMVjXuQT0NNaQitPk4VMXKF/ezjpJ0+KHsBPdT1HBjRrAU7
Wc8LftIvGbB8u+rITQEtSPUV5M2OdfE/ImDzCNBjCjqiIynm9P13DwLVXCfB
s4lnN5TD8CzrxUfyY5cx/2nRM3ye+ZnVKPopi0oS4KfqB2cOd4RUYnA/Ds8+
Snacl7VynAcF14+SbVRSJ4pMCoCwY9mHs6XMq4KZajgwFxwNFXkMYaS9cYQ8
EwsJKgoMHIemanuaCmymmREZcufx9Vy/itOirVHgIJzjRSNSNCIOZfs/O779
s5suoFGWkL1pOVwJOkKfa8c2pIitwkO4yTXDUjnPS+83QAmJoBjQF9TQNe2s
kMByL2EFAQ15VUkKolzVirduW5ZWJEn98eNEv1upqTVxu2z7Z2KluvV+FKDC
yqUgKPJyLScrm4AKuzEUT+fl8sK39wm3xbypO5hq6jnj/LhjReKudrx5Ajxl
OhSJTDISHWrD7uQosqwLlWSjT9E7WpVyOKZseSirpbMmQLw96O538GI1Vr89
BKCy00WWzG+2gC4PPjBgXf63anSXFyzWneK/nlqe6ZO0OOdrVN3HiGBGGNqY
ulcLrlitNNNZCarRvQ56wNvw5A8w455Af7/7YjbkYOzMmCy78Hl+Ho7gG6Ad
QWnfHLqfcpJ+ouP34jDE/kCisOwZcCvyHqSrsyhEAvUM0QJq81vVx+Hr0LjH
WF1CwFeFXms6ivLLzXPAB5l7dV13MYYxgyCSfhNTjidxZvl0kf4aQxt1bz/S
PiXsSDnkZhg7ijGgqIkepjX3ij5RVg2xGtyDuzE9RjhDIAchRJ9Yu79aZ3v4
fnz55F08a6osxwv1EH4hMr1MM8Cpi1wA145q3p+aoy7thMddhgtKBV4AkmZN
N6dWCEm6WquK9q+UKyu1XGN+mq+/GEOYHIO0dLRRRG2DdWWBQni9WhPJuWfA
q6wDoKoivgaC+0CKY/0IPRe70CaqoEXFbrYCnTErTh/1WQpLziXtsNFSfiy5
G/H2sphOEVkODJUdl03K2pCCprdVHUJCPiXLxd4/+xyVFhRuJZNwZuChluJV
irUTwiwAl0cNIIDZ5M+AtWjLYL3SCGfNHklJPpOUUdwltc7/M5VBlG3xn0Nm
m6dPF1k9rfyY8D/oNRwGjdRV32S5gj7qL5UUPNDCkXGW8MmWMOr6Vhiposln
apHFds3c4qMcDo0lqVRejkJG/V1Kzc4NUnLs7gxV/smigUMUcXmxQBPxyO9E
YJEtO8kC6WZChe9qWC37aPn69e32qpIlZOq9MiVUdZxamWEh+G2e4TL22GlN
IP2dhUFllZyrtzVSydC2MJr/aCFPatqJNGUwqgODO/jRc0t2AaDcybp+hfCx
4q6ljIje/zyefGntXnIt4gGoVlMkEp9z+W5Hsee7NeCufX8XZKfzC0Rs9WXH
YH8db+kDL2AUlEpdcz4KizQTZpvcVNgMj09+Xx3Vm5va+vNP/jotUrNDJdOW
OdtxJGnDGw6UOq4R8FkabwKp/8SoBLJWdTNhhYFlzrtpBilD3K+C9msCOAsz
L41T01Ei5PKXDedf3fOx7kAv7WWM6tzXXGAzGf7yDtcJrvftrRGHbyKVXHgZ
IrkC7uM0DQGEwP46C6KWGi2DkRhp2gURlWlBz+xoC6YbFklQUe0T0ctT76Ob
Ze+8toANRFf2ELrvjFV2XeCSQmqos+Wi1PLPa+1jTSDPNBXqsWYfgsTYlEZv
2jvSuDszSajqgSgcblmNmppIUTjveGQ51UZ4GW64/ZxFZj8ZBiAZjgkqvMx0
Vjmi6pC+qj94wfoXQmOt+02ezrQNjcHyrCdNd0NO6f18mDMftmZZScPNIs1v
ZPpVTyiWuFDUJdWO/PNfgHquZw1IPZwSTUWVk9hoNP5qwEQAz1RqtS9QGUmF
mGgE71GDzigR/+KAj2XrYKSeJQwuiycx4tUrG95SKkoPUA38v7Y7ilu2fERG
7LLGUe+Yt5ePSixn9UBhdyZUUY1+lAS4UH66Y9cOGg1grQr24XstLnddGhMo
N9HlbOJi7kg6/eYronfS1kkBA2clc9eabjoIUHr6D/J9p17fZp1LIxe1jte8
HUV4GXSGJfa65fxKuiyHYJ866aSyW0Tvr1uPKs7Movr/YTj95z6Vxn8JNU4B
VXmf68Jo70ViHV04Bd/NM40QdNC2HYFrXfG2nOB+nhx0fFzEs+r4QRwc5WOt
33wapWIAuf2ziC8sO6U7XfzSyGTkYCXDnJqlnkLBWMDWr7ftyMEgDRum7kJJ
1GAoMXS2vaOXb1hCjKbqss4e1ZwovsIztE7n34jCiywjaiq73pEf5Z/UNR21
tdWq+k+tgOBIvF6vmIL5gtcFbMIB5DU1/fY2qc0u/Nh6S4AWxzlClcDIzdwq
rFXjRxhUhYGRuzMxUmpXZfO50sCFAUpd+noHoOuO4oKqBdPfDRywBWnQX+AD
o8ZfBJwgRpYdTJzesuiSYDRZqugGaGE9RHZgoP8auLrxLFQR/W+5bkkCBAgG
J7k3MAz9g4Ide6VeVzjiwxKvWaP0NAgaYuNGuJjsGTpS/LYVbAGw4ZDGDQpW
WJbDRtHLErUus+PCVfv+3b+EwLsKqh0u6M1hw0fPbt4S06kKuNvSr700JM5w
LblCM4/5v3y/RSvFM8iX4baqpZvmtzQEoEZAHeHKYmnDY3p1qv4BU+bgcSAN
co6cJjoVplMbHvX5oPwSHx+5uD8cXD8YvCdCE/pv+MBzBED/rF1y0LPU0rSb
44Ygw7WpQvFOe0TSHJW8sSn2uNKMozuL3mdTc1bC4c0cmRTyXefBi2qeNDpY
TXqS6sMWtDiHPKZ79Gqhb4XgwUJjHLiGyp1Uw2NXSUpL/+RnKY7bHdG9oCgc
34eZBTEp7qE0Bhn0sYg0VqHV0g/o70uEvC+81M2hnCDdzeKPc5tP0HdvBO8v
rlTea5QUYPN3rM3+8jlnvstigbOR74ad87HpYCyLi5dt+ZkIWB9F/aRWhHLM
yehcAy9fdGLwomfNg40cJeiCT5B9SDlNhGiZb7yyeSkwBc2cMssUsveyZ8tA
bj7G9SxaEpB7wQfMa47zMybGGtR+IJFFAsjSeRytVLzB7R4kD7aOXVLi9SIH
UFdF6zlWYYKZJbrRYBnQRi9QJ3gDHK7j88wPKqzsQAARRyLg9+Q/OdOKLSQr
RcSu21SpAMkIFKxUSdavNNINQuvnwqHNduwwaSnN1ZfohT4nXzqDzhhnxQb8
RM1gnbv2DjpazhBI30j3PUhogsLUuo4eJesO6IvjslDRvpzbJDHSsHbduod5
WAKamk0nakdNyRkn1K9DyrmohGcmUEV6TH3zT5Ts+OEQpKBt4F3kQs22ehNd
Wp6yGtSGyQ7pavj5HHNkgPCpzniO4W9LVRRAClrW6OFzzO0EGWiYtSpPy4qX
Ozh4CG4N9dv6LLPfbBCJVacgBYDt6sBHktONhwqMGYPJ7N9oDP5vBLEnKi3A
yEpQLtbYxSCjR84yENbj4EEAyQMivnUGW6fIbawOfj1boLV3lhi/I/ssA814
AZUjbRNxX7H1xir9zeOLB9CKCvurgzhFpe1rWQlpJuOqnukYBiY4BItUKhXR
HsQHMZv6q/PbEMay89gP1jJo6IYLpM+1ix8oekeIV0hNTsX96e8SgCcqDtO0
d6vzM2u/nfZd36i8UsrwGSnTD97SsKa3XoVqLmFmJjd9xvvl7jmgEB19CBcS
lq/i3McH/OxZZf+Z1ERZbM5gs7ELcLUL7sawnfDQ7x8/gXwtACtAs2CemFT5
zfObhbll3KPXLS+8JheU/S+9MpBP9/PlrjcoQub53yne0xedTuttA8iBjVdt
3HzTH+86GA4T8y7VM1sE0wiBSrAsS7y+IjErPPaFXI2fA1g4SiIqCA1V5+2x
3TEVuA+EQhjNTJH9+8WTkc70FeUS4LoKtz4vQvEvIp2ziavUicVaBxppa+ih
xOfx6ZO57N+UNhYUk9zB3zvFPNkta7iQJQXiYPMqyphtPOpBMLEQRQw7sZm4
WIZqid5d7znx+6frsKcZkY7yuyBd7bFRw+d/CDxMov/aVlszZvLQcyca0usy
zVNaeURKR+eBOahmEzA+wMgire/nB6xroD3Pgdzj3QsHBahiej4FbVm7arrB
aqSiqyTOYOlrR5/CS45p9pc+n10lfw2djsQvUyjhvaqwwyUn2QIcaA8E0Ug9
G/KajV0GuFYirywhOSIHaFH1R0I+7Qb7hwjzOz4Y0qiJ2+pVLSdoZ/uZCINQ
XWI/5ergUNtCIOCE1YCsZ609006Heyj/Nk58IKxjyvLuzworI2Mnw1oJAEU1
9mZHD2KWuADYKaSbQ+6qRRWdY20IV7u9On/9cSqz8V4LPloKJAhaz7jJX/8c
w2WdM2Be7yokBXX93VS912Y4xFA0zxAoJne4k32OMDCr3dxD/AqsmXVDSnvg
dQRKMADIy9lhKQNyYfFuz1Zxx/yQ15Y/jRwdnuhb6tEtbN379Cuo0d1hGFpU
hZCqxwsHm6qnBuFUDLZHexo+HAB2UN+IcwhqF3WBTjQTheD7c7rPhKA/lZbb
AIRGGK8T3goT0RbR2dcTRpH9Sv77Yy7bNhJcZXbNyIKpEiyM3yoLMu6YnVs+
ZPv3oMhafMqrmeiKZuG9D0vzne2yTEsOnbPOzNK3biqVHv4CXNrliwmyXddi
dOunbeN9lyPs4tVFOPBCSu2YGYj0zCCbP+4bY2t75WNswcm0thyq2/gWxFtQ
L4Ypd1yODjUDSZ/C4cVA5BHdavNnhRnlPobwrgm0x60qRNPOlCfB7r9QQU7D
En++XRYoRwumaVq97QA4NS4ppe61gNB80JXJt0WoT9sNxabvi9vr8OzPLSzB
MgidNX7GmxubsYExZ0WxgI8ad5XNvxH9bA7bBpTEt38R2qJSvV04MfNK1pn7
V/n1UTqcWoBkbi3Ves3ltnWl7XkzxLGVOBH8wqXAJ55T6icrx0BkYBZ/kv7+
MGL4hqXcI2awBbM/L9JREvik+QV5z6swMJl+hq4JvBZ9NFoDQwQ3z757foXy
HyjvY+xV2koVS2Dgdfvc/juQh0zAdIW83CCUjQvC+YfPzvbl0o7ptjcpLagy
knfwA70RhL5Z/lErP4eXtm7sLgwSTPuZ0lNB/KH/dOzHGzDSWQK+4hzRNmxf
F/NQMSQyGJoFfrNyhkvHt3liqXQg+qTh2bSVpRtTUCL7c6sPhGMOyotf9E2Q
iGGZ4edZn3NBndy92wY6j3FR9AJIIS6f5zwn3mVveQHqWMk9RXE07YkaeEkH
a0KxD9GUdU3mYni5enVwJCOv0LpUWWwQARnkpnj8zIPnMziocvGGlCHYbTMt
Ew4uD7Ge6+gjlMSp5iRip6snev0GdzsckZlVKRKP845Ng8g8w3CUR90sB98C
nLbWYXBpBuw7wnx0ZELfEjgp/Hkz06jOyAfY+3017lqwT8uUn8MYfDmwvTuU
7gnFQSNm5N3nawBqcMjxV+EnFHrC0zNoTcNm6kKA1LfpbR8BqtLpBhxEn8GC
oAYAO/hErKafrrXTJ513dI7dznLE3XvXoEkch6eumFKw0eGVehWBnTm5+lfy
92vGPTuQH8oQp+3/9bx6nrvFOuNqaa6GvHl+J/DDF+liHLne4D/ks9qYnRFl
faBXD9pyGC40kQvyhDDto7kprZgxTYqLCEa+Ayekrn35HR49fmrqj2z9T656
pj1lmhblvqUYMG4ogp4QCpjk0QO0A8Qc3Wrl3pZaCiTNgagna8oWQxwKDOp1
ev6iLsSAtY100HSuZ5C6FTM4wd05LmGTaDSWJieTWm8l/7Og6lo0XBXI5n+1
nDiAOzHSO4ERqCxe8t3s6OVtUlwDT5VsmAT7Gx/T55KMUYniApyMk20epJ/o
9asWbzz7oPTc1qMoqx5TCq1YRh9bVn1PEyfTtzXuGFWbScafi1gcLAqJapdN
mQG7q6a2tNHrcp/0CMYinVreyCZW1ZYOx9A2sdwWbHivh6+DNNtSSM0z+pjY
vmFLAUhun7Sg+CmKAoOUrthOcPN5u1grIRUP1BakP7p47rQlni4a5ipiovQ7
5xFLo0uyjSf5/lNLsJq80zGk58OSKG4C/VpbDHrk7deTZw2lYzy0ks3afZ28
4V4AgsRvBMzqUaCWju8jv+/yGBnJCODc8OV/l/Bns8FdDBvzSMGctNo3U16d
I0yQIWxe9JDwlPfJklsYGoi14ZQAPakwre5sMgkqK6nwc+xX4FUZXGY/2qTn
f+BuiKmEseA9EH5jOHf+DvSWi183AxzY7R89ZdzZzMq5DFtuuOUjGz/4tCqa
JTR65OOMxIoJu6UEL+cbWP9J8elKJtFACzigSXAx+XpVwSj1EIArQshItlhH
bVmppEQDXy7kSRLkWToxXbgcWwZFBqYybkraXzUc1zbaneW0WSlRT+Bc1Tvo
VGfWGwaepqrItQ4S7Bb6BU+t/sdVEYzCuaeIKG47dAzkk434m+k1xuq3KiKO
1l9SKvOA7F6jUqJNMuIz3eNHamBIK6166I59RX/sGApcIgY/LzhCO2Zsmaw3
C+TDZH+ybP3QVII0r4OSrsl/8ygUCkKGk0NhKqN6tWQauGI5+U7pveH91w/I
Ek+9aEa8rNPu42R/YESLXeO9I+2u78dnYIHTSYZ0fsfgqMLcyjxJKbmNm0YF
pJiiI92vSeMqn5SSDAk/Tz0A30K27nTsfBsZg5UQT97J/+140tcbIFBG1Um9
XMDh7LPYwU390rcRV1vcxchnj/j7rCQUOEUYVUi5ciIv5jbadU6069QzHmIz
EjdSqdM9MTk0IdZP9z3CiLpm9LgFt2SlC33nG1usB6b99J58xOn6j7Uy/Wuc
AYABeZ5SCiQ1bi6O2tM9guAB9BogVz35mhblTdJ1d7jzgJ6stNDnVQ/lFBZ+
bDx0k9ec3rMO/4ceWo4PXCw00wGnVWp2ePx19N/s1d6Gs7oZYX0w7ecT8ha6
lkbBRDQDKiRKagZbM4ZjlZrnqIjdTKBtGgIL0ysPeoceieho6sGAbI+XhlSQ
RivcPTO0hnpV7+hLYMk8AmgBoLwZ8lD+nuD9OGFdotwtNuJSDUMA2YmKsR01
5dBJmtIXRa/JjwJBnOGUMMJ5DrucxZDITqtJquOLYbiP6NfQs3kny0ncAOUY
sx++OFTTCpVvdyskc0KAC8jwKSgy/8m5GC0q6iLCXyIXfPdJD2gy/mVkyQFT
yZcn2LpytnfDNJ35XdWmVRBiw15PO1xayP38oBH2EUDGuYyJqsbLObT7meWZ
lYlMf7P69MWklKMhqii6E9AsfQA1oY3b2xcGpPcbf0XXdhBqS1ldSLcVwa1x
XjhZmKnGbZSswIQkdXt7A7PLGRP7XpwRwifDQ07MCg5i9bHZ+x4qAMr0CrH9
oLcJm7M+ek+fj4crj8VoUzK8xK1Y6ZW4EuQbOwcHVl/VkeEvHKFhVsTsJ50m
S/+lt/DpeALaT513fP82LiBNjblbITN8IIpKFWvRIysatcQXaoVAwJOVExJp
YEh56kgMn+1HMppaesxTwUMa19n6AkCLHMf2HCH503PbyC5HSwZk4N8+cTdY
YyYWtd0HuOJTMAHe11sWOuKRaBSr38bTgyJ/TIRjHs+P0R1TGR2cqOtM7d8P
4Em1vadvl0JyuUaz7m87S35b9aIkXd5sHvIXhWH3f3ncmhJxjKYEDlvcSL0D
TkFOMUjoboY4y8n1dVcNBAFfJaSIjhMboscTiwmy487vUnCC9bXgvAvkHJYV
5s2Nl27EQ2zF2sHZX78vyTo/lt0QV5ddTvVWoHuvJs3jDETUOGYB/bfy6uF/
+rBeMq5e2fWHUsCP5xaYxJ2ASga/iwOhx1moi2BPGbqv0FEahO+I+KfmkXRs
KK6qnEh/ETt1VWt5Ok6zmzlvxVFH7t+2nwCLHupb8cUV7lHsoyLyKH31L3GD
wWEDJ7B+N3aqDMls3qDFZUjf+CLfohuhemu3bqhvF7xx20yeJYOocc2x2QzT
iZPCTgMlTy3a6Cvk2yq+441tq32YTy7Op/y8EiP6ExVp5Uj8ZBl/oBvjtKgl
0LJ2Xyes/4mHXM0F73+Mt8PAyWvQ3Dp1zInYTipdjzjwFVpEc86CTNWCpz+g
Ikn1uP/V+21wMDl04atXGWOJBW5vs55ouaP9QUBfjELwwWf8lh1GSmhhFZUs
1fe/ulxZLeT/OlslZWPI2jV9G0AU0ATAk+unt7ecSlhjDG0Qdhdv7jdWNIve
Iw/xGq2m8fZQAhpkTyHCYdpk+A7sDBqzrB0KQ7gls40naOrxEWd5tOMM6c0t
RDJ2XoCbRatZ2m7scP+cX73uIefSMAF27ofAvXwwaefLj9YquPhlmP9vOSCD
22Ia/8XE3hqs5JdM2/HnfJbqNxVz3E1ym7mxhW0laBgxbkUNf92sBbjko6aE
PvHTt2MJLwgte2E1CvOoOcZChtPPhTyD114snwUZC5Twk/ymcrBjrtKpyiD2
GRDhFRBGLsYX44eREK59yhH/iV4vbrjKPlQZFAJS3VPwycGKJ/A9+5YVR7w4
cunpxIYrm1+4gEXffbOaC9AwSCLO07u1E7at4Z4CFsEvY3dWBZiGDWO2KXsu
mZxWQiTgJa5PrZ5tP6Z9IJZkK6TXFQ9W3HcCqQJWyszbB1n6ht7FBawe+E6m
OHbmfekhd7l8M9PB6bxvlsrAbbUAYOCXne9HM1EEAwC9/Gdrx3MlRinQgYO6
6ILCk94eA6WfW4Co0tTFsfOhUDb/4r5Cn45UZXJRn3fktMSMBS0F3YzdqDuN
6iwc47Z0MyIZ0gw6XkxrJPLlMRqL5/45VdvDDYiRFGGPdWb5rtaEAlZAboeJ
ygYsX3766NrNXZB9WnHN92tv67ThEwvnyNwsck05aIYNH1P9jVVdO/67h1AB
FbR5HgXxd2y3Ms7TKa5SWA941s+Wzhh5uyol803P+h8hQ2F2+M8Sd/WM16al
i0yV767lQa9UkCBs/uWs54gtCdxd0qA+NP2PADaSmvxQ8XSc8vkbNNvjGh1I
lQ7gfYVlNzRh3FNK9nDqlUE/oagK/UtQvDjw/uZgDAOeJs26R8e7Ssge2Aj1
tN3pCgvBJSN4ZlUqojAz/0toifevZdNxWxxCI8gtUG6Csprc40tQnn+1+xxK
+TubJ45rfMqWydym5I2JA5zjHaPlyFUL6FmT8NXB/wrXpFMXQpX7LAV1Tk78
pHIBk6cxKW7hN41GTfy3RjnAgKw5vrHkzUukZqezUVeEt+TddL80I9fKoMvu
7i0jYbJReOeSK7+mZvA7Qm/cAasGIhb3nbr173V6MqxNCZ570AHwWqCB0BMg
B2JVxnbIIkvugpdNE7zukhBCrlXyXGN6PYFpinyAL/NMx39OeVag1iamu5v7
NLvYpbF0pw2PIuXozHMUukvHbD17P4ttbSg2QRqxux/MKEhx57bKfuN/wajk
NUNMAUCUBPOh1C8wL1rVseaVfHeQLEndpoIUAi2QH1HkOO5L5+w+aOZaqXX8
mMBJdLkAkGtAmyGnnDz4jmkSjKI+bqQ+AosDVLDJlaxgI/JgeqpP3OOxuPIP
p2qkmX+7SWKyXT3lNLnJA0PnFDehk7+CWc/opFWq4EeXd0MdKmyVQzcuTHCx
OwoWtG4hW7UdnPKrDuODM/2Q2jwQbjg5fcoCEdkaEkflYw8VWFphjLca20WE
I5zO2SknbsSa+thu/SuwTxCeqc3Ny5CVWtTJULVRAw5rRLp2ZtdXdGvPFbMn
rmbnaFcr72WqDtv7pRqqJvGt3FfJ7bFMkv2/E7gXR86PLJaH0xwbEwgk7nKA
hQZ14hCk/kBPR+T8VYEQ64sZSrYKAypQJ4BGcA3eST5lLCd8oKd2vTxSmCMV
4pN7yuC41ZLd7dhCOZAYGdutqWcXh2JDP/2RXE9zNf0peSoZgSlcdlvnzcRa
mv4upPEvZZlJx5dHlcl+KnnZ0qG3dEgrWFM3t6Q5oC1IBhu9PVwXNuIBWD30
Xe9HOS0780EmayLf3Ko/cVOqHNMkZr23tqldhCJscd5LsAusbKDwWA5LEQq9
twrz+2r8TF3fjBwNGj+owcOjY5iEwN27/irb99GneVGlqyljMSB2Dtk7sM88
uXiuwB6LTOb3o//b86t+/bbW9db6uIZlKoEu6hjICFcEHbQZk30P8iyOjoyF
HezseVb9SauiX3aReWfEGRn0YMaiO+us/GdkXHYvJaSVrbyE4g052IF5hYNB
Ye+6lUuwJ/PazanmvDflfcnDesb1dBRHvEAy5hYlX9cEkhT9JUSlCH+MMTEx
WZxBovWxLBONW7mSwxbzAAoxNJqBn3HQeyy6kUcoNlzwfNK4W2x74VkF/Sit
1vfJMPELJq3SFE0C2BLC7mN3Zsv9kTAxGEGF538zFKQ+b3RBgxlOsnB5+Y5a
TGNw2KnFF5e8Vzfv6DWrmWw1gkszTONPnexknnEXHO46jdpMxNUrRlpRNSgp
zgYmUt2Ntxj5WWopZQDit1KFU3N+hbpRJlfOz2hzVpXCMzTY1LwKPrIAbrAv
2pAreKJGjg299+6gD4LQgZnNL1vvVZqfGoXyYz60jcwUCg/O+vKZ7CwNnU87
Wf14McsqRagCm9OnDCna0FeFGRLUCJqBQTsHhz+qvbpQeh1JoWX5XGkYPu4d
r9HIe85PHKpd1IYhyqiQmIPySP3//fVPptfHGgExcbrL4aHHlMXjWWa4mOP5
CNlZlVscWdRJt9kroy22YYOINtZLcc3K2SpaBv4/eMccTtqlMEr4Qd90LBye
Wua1gD21/Gwm+WQP9QTRvAwGa6nCyqmmDGLMbHI52tvNJOTaS+w1l9m+PxQJ
Xv+mPZHKJDG0vQfc8xbLH5zzFa8tGqIGQm3RGQT0c3AIx0D3jRW1XscN9XAV
QpEBXZ+xu/do0G6NBb6mrQALqSwVAHZsDafL1/xQGvh57fACCOi1aIPciylT
7niUEQBuz/gTHkOD+H9ZQFfkXVKXqMW2WJEcJq8uIxAFJtMVgGH0wbOleUbx
pq+W5X3dhFSrXnUXLnzYNP1DImJMz6yj6l8vMWQkRtpHE0ZIw3V8c+7Ry7Fj
wUxQbRROnPok/gg/k7cMA8PZdd/OOFec7PbtPFYFwvigBTB0cvHI1B1u4v8a
L1Qxs0B1ALamtwUUJv0Zxg7T/yudcZyb/7nxb7im4Nx4YzRWzOAeDL5L6Grb
wYGsUp7gWcMgnjt7zLqqBCtU5peYBH+Rdp1r3XTFI05wBxeJpslxS21d0gQv
gnkeb+nfxHVnnqnmTpsRA7LhxPflgxcDLjRgWhEQO3FiEw2KpRsFLIn82oc+
JI2zKAgI7gfoEDwl5NNqf7VA8+OyQAMv7QEOnYPWxyd+xHsGj+PIg7DE0z9n
fuY6lmCMQYVNS2Qa8D5K7Gx2lHFviExNAau+Dzq7N7bMeZsY+wvUYLrVU7IE
MBQs4C4sxkGiwaitxW4bpEsH88QrwJEcuoMQn+msyhoPRniVqukdjedyhwGp
g6DeBPzTDu2jCD6DYobO2XJQBlJWe0FFuSM3Hi1Hp6CToCAKRLhMV/6GJo3S
sUyHHprSLB5wamp8vRFrV5VUwMWDRhq8PPD6/ev/mrkg0qvFWQA+yBQzcwpc
v8E1+d5EI9P5Oqe7EJiPyfa2CcGim93E45P2OR+iIDIx6RjTT4KGzPLVVfXj
X2MJxb3krKr060eOKjs1QMkgzUhcnPKumHFzRRUAwB2YmjNkjFOIV53e9MrD
sddR67p/Sli9s4MD62D+S8ahaHsRlGgnasJMzofJbDDkl6adBZeTZin4xXTp
AfkbP0SsIlH+tGeo+zpHqoZP9ZXMa1sONYGNs/u9GiaAjwWysv8zcm07UBB2
qkUnO4cistzqO+v87jYaP+cRtlQgxxzLpdlsWQzmY6tnsho7OkcXHTY9wjTU
ibwKkb8+6Tbc8w4vSTQVdwerNIe/CuKCw/FT1wvGRjrGFroSxGR1NR4m0WzH
thGYBklsvERzmbak+80BJPQzFNPb4AOy10IPvChMPAYYN9fLnOpsweDzKblI
oEH36IQ3Lbzd8C70hvYjXADz775HhePvsPJRNYlPAmBo2gKxxhvOWDOiTKkk
Nh/xWMtt6zGKdronnGVy1N4Vqc+h4cVvngs0b/QRiGaEqB7WmFCCUrNNAIT9
kRj5LHBneT8YPndpi8gM2KUO4D9xYjWxCgTjgKb00HvQwDRx9nG4RWEqo9ai
+fozIrOpr9g9qa9I14TUvHZ9PiVPG7qi07LHihcR8vpGoey+9HN1u1dJ1q54
9Hvu1kTFYEGn6ZsJE06h3m2S/OjjSEO2O5IJM5Jd7PIQnA7cSm0yN04WksRN
MO4heWW/ZDuzevysl+eRU6ThedA4jLdL4gg78WDkasi0h997FGLE36qbHqOX
I/VgvkLvmcsiPlGWFMjLCZ8lXPQ2+AHgwQ68/f/HyShBsgG19RmTcINdH4Oh
qpquv+bn2q8Dj1LuX7sClhd33WEiDe1nWP7VbI7BdhS6m3a35Kc9iQ30+Tsu
GyP48z5MxuAzgCBvxBkVwUwDPABOu4U8PUNieM4f+OMmH25EjTsmRlHi9hPd
c5dBjrCKzavUVEmhAeyEb6S09yIL2BpWJjfNXuF4CdLkcvamD0TEeEv8KK3t
PQOuo/mxZ6ttzNRxw1f/BH3e9VfOXAu5qx6IramlSJ6o5uh9bhhT1gb1mdFe
hUQ7wXigOlhUXGVXpT6LK1KVv7Y5Ny4vfdpwA1fuKWRhBA77l2vVLkiIzCrw
frrryCrhMV+ePUKzxAJEzENtD3qEce8ur/BpMW+iTWHGfn01mVSyNFMxbagh
1HnHX5b3v1nhz4wItetQJPNAEoZYzAdREuusk4JD86hCWVlSk8novNUO5Med
1sI94l07MLPz0HFw4B85hkk8x4ejRZ9tZtYE6ICCHQSShr7GMprLrvUTmQf6
28wNGXn2WJmZHolz9LnoS3TpiWtLErns/ahBt5x+dDcNiQukIcbb+IBNSBdI
borq3WNhK4vtWi/+WDQXzYH/dwc94SHMfao6TzgD5cYx//HJJOvZ+BWeQsgT
PuYusvZFznuOZ+TO+AdbTsewYng1Q4QMqWMJpiiEaybKxr0dlgbkAh0Ojdmd
ol8nCVBx1zC3nXk7HOPtz6PyFkIjs3BD60DvD4Yc3EQ1MRj3TProk7qq3YCq
7rn2mUldcTkFrgvWGDLKx7Nz9LKKLInM2KQ2k2qAKpioIYZmsvHqDbh+atVw
MMVUzxQv0foAI25tgskpRvCFV6GKDAtDhb/3d6h1Vvh2UGIhCcbJxH1FXc6R
AZwByvO2DagVbqpSrtOEFziexU36mxA+LsTIyZargEyP7B+cS17Qmg7eMv4e
KNkxZ49mpK8JhsHEar5EtK399S+T3zY4z0/Z+QguR7AbXhZT5LxTPwg5OC7w
VLRIRcInkgl/Cgve42QaTMd/WhWNcNo4VWkWwbmNUSqURinrx8KmWSq87aQK
e9uMAoriKVlRf7HwqdH8PZAEd/vTIjs0v1OqQC1Dk4wIfijGoEd3MxjVzxFJ
46tHbxGqwFsKu04rxZY3CpxFYJzmsitge8r2g/AC8Th7mmBtdhaL1CqjKcXy
r3+zJmx4HBOu4FdfHCCFD++g0iLcHq8+rkydtqgDylHiS0UQ/rBrL/Pl19fj
pL/S9I84RXmWdUaXsfU37ZSJXSiMY0tny+IKp+FdtkVDl9U0gbN2c3OZWgnW
7D7Ms4p3LIqpk42PzurpK1RjA2V6NGHQ7NE9EY5T9iTDU8/mElJwbA3/MX/7
V3esQAJ9VFNPzuBcc9RabE54Xz2fvQ2BTprdgC/i4ImR6nJmIfCUGPRnzsli
pyGib9IasCsWH+o6PuuEELd9dCLxw660C/jRZ424jjV4uOZ+nEcoK98Hgll2
zsN3qAuwWlE8IO4bIk0ZV9Zcp9DWo4AwrYSpV87wrSAqmSYPI/nsqSqfqSIl
eoo5NJqzfknyYapIBcSypDmUGePp/S9WdBVuX/dul85Qu/6Cq23Ap773UBfr
f2cljsEJ2bSxmJ2X6Y++p+40rH03JeDGSD5nwy8oYU9wCXe3gkhk35+CZ82Q
TSzLaf7nCusZSJ72wDZl1ReM0K6mkR0mgOC7V5M5xqAc5k/JA5GNvUfuEgsg
qzwE45eDoZtawjvD9u/dek+GqWi8hMf+SbBxOs6mfg00rL88GZ6wIT5sJ5N0
QX7zbOV4AEtNVsjPtQBI0qxPG0WC6cWSHREQv5EW1vK5NWk4GJli/M50k86M
YlBxbr3i7ORdPiXiNRCaYUcfH+0mi4x7mb4RoXwtdvlObJOA2d53H49x/Wls
1hw2jZKqFfyTNSQ7T5/N5Ke85K1Eao8014UVbi/5GQaFjPGQSuMWD/gJo0Dw
IT2utEXRMvN9WKaTJMoPiMO4gC2TCRE6DzErqAdXytMtt/XtYlKgPjfkUE30
qZqEW+mM6SxI1wZR2tSN1cJg8ESFzyIG5eAr35DioeDBP3VDpHfZI50I5k2j
UG8yqW/B4XTgmnpLvnbQPLI9raKg3N7NtsV1CskKKJ0FYbHEMG1Va8Ps7pcp
H1al8S7qhZfD+bCnMfVS+vyBsxBwWLEpRMrTcqE9nsnmEJDyvwKpbmke/8Bg
YNuSkg0GBA2PJEP3QsXKVq4khtXQxv9CNPb0z+Umu2k3aqMr/V70xFsVpJa+
kupPeQq4/DE68Os3E3CA/yBA5uVEzQzw0sK02pgw4oQa7opm1RspKD7O6ecn
wOV/wo06wlOkvWuVgV6WixCnpyLKdzv/O9MXC4qntgxvkVxGDM6mTYKPJIak
+YBiGSinMkYoAojUdILovofnVBASRZ1OEetr8DfbHytVKaRmwVG5eiM6fJb3
WMVkEml7fs+r+hId0OY5QPmoXlq2sEgWYtW7gGe6u/Hs4nX5d/iMT+DVm7kn
Q4wKfyldmKQNWu+VtOxGMmLe2LSlqai/i4osuvz68wR4dQ7pbJK4nqo2OCrM
K/XkMCWuG69yb4RkqtwTFQEq1tV8ysH4JZ3o167wrV0VHQhHMp5OyqyE15by
iRm37nFe/tzZ6WNb4xf/q7w9GcOwYWDhvUoq3GiybNwPStP5xCn25k/Ok9h4
wl2bWM1Y20Yn+JDrZuZrvZcxB9NY9BHuzhjX9EfhivMxc5CYKJcJJOARskix
g42gcdzdo3LxzcE6P7Icwcfmgpk4hdJeeIXIlgAfkSrF4OWLpgb4TGfozsQU
r5dTB3jE4KrNwtAUuDba4wqjOoXN6aNJR5S/PH1c2bAGOhTSmerW5heeB7Fh
NZQpAAINvQKxdGg7l3dH+6tLLNcTha8YEYTz690O5wbwcaSaYXp1IPgzYbMO
bpUBLAD51J+OpLcQJUsg+qETlbqhK8IQ+RMQ7IBjMMi2J79XmquGUivzasGz
Zc6RiRj8xTy+IE89/7bTXumA4/1J32rNW/0E4+H4N6Qal2eEMBZ1KgsFL5pn
jgbba6Zzcvgug89hUK8XqyYjXITozI2TMLWTpI2ddApbD3mN2T+nGDNHc0SN
RKeDMLRCE/tnQlM4ipchXICuhieEWaVMdBhNqORO387DsHgEDEbwku25ezgR
AjyPe3YYCVvgdojYNbbmh5Jpt3hjcP2F9prupuIOL32gSqK7iytekp8lv5cM
wFhXhxM50tR7B/UgVLSBk9LMIZ8zbYL9uz1BpHbFbPR+j5jjcInkeLRGSdxB
BKTBuY3FaQLPLobNiIo9ZRqhyXJh2Q9Yxeb9z6AIyFozDCLa9QlScVpJkgEw
XNV+mumq61U4gHliXL65x9KXnSkP9wzC1fJXBqiptpnMpcqIkuVxIPLQkK2U
EYkMlOOQCFi8HVXT714NTXoEWYKItBlkp/oFyDPDYNyTDXGMRVL8gj2yghKb
y3ithOqGdu66iLktHcmRyfq8LRg8YMrDlnk7pr9Q9IoIMLnqVJiieIk2bfKm
ZFVj1WhvUsXn8baowXuymj00hVhSa6FxqkuPFozP5Lqbhd/8ZSX+5y2MKDv+
nqShhMs3sg0d+uV2G3pcMg67QITV+Xjmwcxha/ssVhUaRP+eBnJCWtX0nE9U
mnC8R+q2SQhEKLQUGCkeiYNjY2umdL5n2+cmvFXnQYh/AEmzKIHJPfnNXXGD
sCgc/wNPEDQrQGYQwCusA/p2bk92voRZ2f70FYeZrX27Luyj5YJuvLfE/NhS
R+jJTn4y8ynm8Rpj2NS3guM1sO+WqCw38NsOxaIQ+SlJ/jL5oocfRS7n+C35
sijKDnNGpDnw19L6KB7Ov7VaJQljddP0+tDNWPFnlSeSV1S339ici6l+Uxax
pgieP+GACiNQg9WOCTUovX09ny990XGVrBAOMkQAFagO0gdFPSzlf9xLqKWz
luIaaqt6tcetxywFnnwkjVI+MZYXc4avEdM7r7AK1vbCvd9E6MRHGuXXyzXY
n8P++Sqr9fPMgISGn1RaXd6FR/Eo5id0Eq/xeAcXPDwuFDxwrRxnNtb8ulTL
855LqOHMfr3IWmVhI+1aQ/KbzADNxl0Wd7TZPIpgJrNa4YEWgV/LDpOrVq/P
n8PMmmZyZsXy0Oy/yv6eYq25MO+B4QfUZewAca0uQre4CPs/QZcW9h88y0bx
5ucVqMXHGEYWjgrdyPlMAKKw9bTh1IO236gVhCqMP1UuU2aI7RvlKibic1m3
5cs5v8D6WgDqt7izXnFL75bz4+OMEiS7TjpQgQdpC5fnoA7sVihjHHMjt95F
QxXMQhlHy4JNRHw3wrctf4gO71jOMteNEKpObikAynzXqK4nEjW94XWcr1YO
rarCkKpNZbi9GaORbxQIYZiFDLX+RREWXnOPjvwgmcIDnwtXBcsQHfz/lUeF
NC16MVFwedU0SdFwqb33+IZJL8h0DSc2qigHE2e1FvDuWV+jwJ/pg7Y+ajeY
OgbrAPmwCRkB7CzJZOw0iw6XOeAL/mbCP7cqV+WL4rdaEoqo4Cu46Kjf7OM/
YuStH/RcO/ggAp7IKKYEbkEQIf2kd3LW0rFSFI/d4QYn31bdKXmPIjh0ETTd
juHj1TPrpE8aOFtM5puyJJeLsK7cBTJbV8V8UZTPGPvG8V/eC+97aMYrBjil
T1e0ihA3Lgjd18PCAGq+vXstKlABkiKtPEp6qQA3R1F0slHXoYthIZApK/jQ
SVmnigFL8xpkT56DvF7KmToRYATT2zk4k6q/gc1rUNH9YFXpGZQD6+9G0HBv
HZ6A/8+uEJUBrfQy9CZBsrSCVwOb/w+sH8NabacOBkUPEUDtPPFmV2zuTl3C
fY+9jQn79on8uYEGJmbWCWtGJTBN7bQBPQJpSfmA1W8oS8cJrHGVFg/t4RlF
Z/i/NMimKq6b106N2DkO49g5VTvHoKNQpQlB2osO1rA1QBP/QlnxjazDBGzW
9XrZFonYeHr1zwNCdGS83fLKCTVr/GN1vfm+uXyZ7x47oZqsq3fmoiz7sccm
DM7y+ObpISAJEq1piLFHUe1tzC/ewv8pGKsAyeFP+zPHZ/NBqG9F+Vamte5O
JMqrwKjGSLM8j+CR3kZOmHOq2Nhe7l7wUbS8aZgDOFpfdu4NWPlYCNgvVLE+
+MqTZHGcpBkebusa6CQcyL6u4bQSWsc7RjYoajrupal5bi5dL2sdCWmYln5p
l97rcvTzSCOUrOAAlGshic9V+Vcx5e+BVAQTL7ddBi3fuwOh0iSvFvQ15i7g
aMneCVhTC5ew9rKlwADytbHWNZ67tPP7hgWZXPFEZU1JzHBwHUNzzkDJIvR6
4nZx6oEl4gRzSSh3SvRZNoy72EjYidKn36CIbM+VvPEuiCJ55ePomFZAgpqT
YEC9yAyowwhlQvqcvobLbU91IBjowLFULfyZ7ttWEvvtgJmK0b1tIV4KD4lc
V3fB/1mS77rpJ9iF87gNt+WRqcG4yNCTYMr7DT3k3RFLFjnIjH0VCWHYlMyO
YjmhKHAUg4MDjpb6TYxJgxidTafcn3y1Jn3vHMAkWzi66ewgkFRu+GTKTNQk
uOKjItwhgy1sOvVmOd1WRiEuQbxEKlyaPfQ2CJLpKMm5X5l0+D+ZVtfv4GOX
yhvxXJkdSTYesnw56PQEfEXH2i1bBSd0LRX/n5SUWto9BRoJVTvvtePvFTWL
tpFQBl898Y8U8TgpmjfbA0kv+ixpS67D/8+gZcJ6OWWREAz1UZP8KpLPjG7z
epv6VppXcl/bs3W/8svl18jIuopRCUMapmE5/v1YtHs/x0jqkv6NNoQq+n0O
BDp/vX3/EFoKdbfqi6nJ2stRlPHHIxEJanmgyQKvBG+CyRDOQnvjKEy9rG7s
LdNdxfuZVgRQDNvdW2FKJ14ax5qU9qYbtGAMy/CvJO5zGN7xaavLnWViskNZ
6kmAfsfZS9ru2W4vRQ5tUTyFSCVB7JPJwQNOF16avdKhDPjyXM7BdNsJgNVj
GPLpFfZPKyX3eoOG5e1ZULFAw8TRPFnny4tCAesb6LfOByu9LbaP684spghM
kNiTEqticb4cj/N22qNGuMBpSHwAcwdO26WZVKzccQxtEN4Hbvjw3MisrQMM
ZsayGtXujpZoZnho4lAIYy9lCGqwvuk8tsCyt+zpc8vtG+3Ir0BtZKbC6Nzp
SVSlgeJw5sU4KHo5zJjKoPX/UnjxmKhxQwW53JNQb19EKQURPoqhCpIPQeRz
GuX2qpnwCINGeRf2A9xytsBHY6gefG/r5r7MEJWLol2YK6lEoJiL3br5Wmiu
QEbaionmZY5x6YOgSblZnapa5EXwJXtfAa8XmdFVppV4CrbZ4//tDo0kRw9A
VixbTIKD4hcq5VYC56pkDXL0sLnflLkYxcymVYE7Xuc5mqHjZwbW50J/CF0i
+PD2XdxR8HzbyK4wXSFgYuXizFBQUG1pmettk96PTHmpTSzuC8oqi8hznoI8
nEj+9rAlafIVhoo1/s2IZBc+bTFCjxptT1V8j9WDKjRxUY1lZg0iHXLhIWwd
Jn6e2KmmRR0NNUrGJZGjkde1PEUB6CSuPB6w1JQJYLD8xX0HJPXIJQb3GCSi
2tU1nI6R31ht8WnPp4wIj6Ti2XwR1xdYya57+0TFNQpyiGkIoheA28CUHMWW
BvKrng3gp0enJHS6VPZ9XbHQtOZCYvR1mlddtB4j2YDI4nOYxUpW4IS6PMRL
wRLpCEjVxHXP/hIu55TVi0mXRJxqTz3jOsqlAkyTY3CP3otUyTrbhYK6OznJ
/42gp603n7AyNAWnbAK/P6aGflreFCWRVESF2y7O/8QzsRUQRyxmGqNbEUqz
9EZlTdcu4tSnco0FaRPnV9vjh0zMVVnpq/9efXfF1OvofisbiwNPljVV3odB
IR1tQ1x+NYN+7pbqZsGdPOHSEMGWUaqXF9O7W0nTXNKRkEhRD+bN6JIAGMbk
7msQleWFCgPdCQG47+6LyMIq9S+N7nudT2tgDRquaqRoR0mdA56m82442CJE
eHSHYMM896erZ/BDOVqV1XW9TyWBw5MzF8a6XvCKSokv4x82qIjvyJekGrNq
AE3xeoCLeOlJ9n8Tm0fwnQEOEjP0UFoOZwR3R+5yb3i99RmRYRAKgCfuoSz7
BPOVWkFkzNqSF36AX80JgYIEorh4XGBunufW3yp6yLcBUowU2PPkvoGaNl6G
+nRb2rB3bc8CoCxbXZ+zyrzsYQUF5vvFykKpm3W4UIqO9VC5j1a9AmI1Hnay
V7LXgr8zdq0CtocKq8033CUG2G+FYrwOqTYkX4woZgfdHnBLPe55BJ6XmJXl
vqMpr8gNNV9O7DmUCld+YdScV749Lo+QkItWlYdV9vE3GcABNcUbBlHPliYf
BOhrjf8GiqI+sczyx4fJ0xfAxlAoL1za5O1HiF6+ybHWmQgHEiWlLezDOoj9
fnVtS429+rU/Q14ZPFDzoZqny9SEE/I+y6JpTZgzBwgF3KL8Q/oWQHgov9b8
rlY8RSZqiqCnUc+Xcw2669kdoBKwOBqI5G+21Ko9uy2o4kTbUdvFYrMq7Z8i
A2OS/tYpZfSND41TizWKYatGpDwfiybYM+57a/u1y8o693e522m/cylaJQ8T
Ors9QaOOalClv+ShXTLSLgXsSgk1+Ttsi5PGANMyV3lpe0Uf1wy8vivEFH9B
GgQxjppIcmvHVopgILAIG0FuY8bJ/VuMjZL95JXIRTZjE7NN5kdgcYvVbB59
3bVbDfroBPwoXLLEqPXxZXHXNRo82mUIxbjRi11/p78RSUJ3zT5YA3+iPZ6Z
oRun0f/8oJYV7H5xoJ5uIiMRVrjX3Y+N07AQDeJ7n/KitoiNNC38VA8KC4bS
+YQ5YGZN/KOdevRBCzRV0DJGWUw2CLaxQa0cB3HoAqyTkqf+vGEpEGfRBmiM
VdqTFCZhNZyJ84V3TuryXZtc/4UoGloOdCPlz89Jqh6R+OcdSlhPPZC3d9lP
o6StflvQcAps7WjsuWuvpwjuZALYtED6VcSP+hddj0f82JkQdcjNrJzuPluk
cpBF/Acqwz+ZONCbMGtwud+Xw4mqAYHCw/Rp6Aoo/Lo1vYPbvp39O2Gi09JN
FkUFIudpERzTRfBM8UysSJosIkujBbFIgppPZF6panDh8otF/odhLUhQHYk1
By2fGSBvCJaeYN8lq+paiLCyoswNHdYlTw+i0PAFjh/6ZpX2q6gVFpgvKjsL
Xn8VekZdZIJUfHjRrkEj6LA6x5c4Z5J7BI06qN91nGOqgBI52eP0R861lv65
BhOrVjLdR0mr6OPY4cFPoaRE1e7ZfBqHp1R/Qa/AqpLDsIfJ2CFpiYCcJRbn
p5Bbivsu+ZP/GxPjA5usXCauG/kY8c3C2TnPQVnJCXYdGiNNqdVd4tOW1DFZ
V36I3N+Hoi1/26YlEtHIaQ6oFdkuKkJEyNaZOdh5aDHutNPZYypP2oozTRgb
+hlfQcucpmNcNLc5DmMg7epQGBUpU40DEPUhXEZ+lbWmSAxbh7mTLk23o6Pr
VIbfuyo0r2tnu1D2jBefDv1+9+F4wzUXVsVucKub4D24luE4z+N9kiqt0/U5
QLm575zu6jyMVsc624LEXcM8OmZoMMdPXwkXvejUWFb3BKwUR/Z2OJKjO0D1
6ZHdYlyKZV6MEJ7wev6SneNARi5HdPCuC9luxIQTI9B0/3CQz+YPFaO3zes6
ZC4vnwegOvttkQpFOwjsvqXNYyQ5lYNTxJ9RiHPe6U5jQWbUzvhgtykgEMnp
yTldaegQ+DJx32rMXeLyrBgN33THnuIdQInnOV/EFYfaA6cslSaoWOrTEJu+
Cd09UjEJe676FU9wBnYR/8RACDdcqHkYd92HH/U9cXGgV4mGtnSzhC6n0m9X
kx3PLb8nF9wejokpVZUTdwty9catjudLy/2bNEDZe3PL3W/pFyviO30jEhiG
7QiXWVfZF0wHVfBuwStz0WumLXE4Raq6hEl2so9P5TB6H6bI1ikagq19JmLc
H3PiXo3dyDO53kPF4KPLUm6QY43QafTwkWnQh7wcAt0rql1VUxZL4pDQZHWK
hYz0PdhnjNtwTsMKkqv8X0FEQ6GIZzud+Dz2hjoI15JKGQGJnucDjGfKFeJ5
kl50e+1gzG2Zx4VXkJiTR3jSmqr89dSYEO82HLmcFLcy52ppp/vO2597/crf
j7S7+62JQ8jztenNczYH12//EZ9ivKOQSY5ST89a+kb3ImhaG6gVU36OwmKl
mZGqAJkoELYr7h5tQ0YFSVjF3c7w2vyMxgIwxRi0PMJzNJDQ7ry9l/OWrAW6
WBl2leQc6s6rTQ2/LUfD2FnGF0Mx+c3Yxns+OgcvIm3oqAHcP18xyVRZbKjZ
K1krCnmeMsCtEOBtxBNGEMe36CZhSC7+jOcOWZ5TcIo8g0Wjh2oA7Y2x0fFS
ROo8P2TpMKP1qETKy14O1r6vL1dd2RBHV4DThpK4JLOo29OylazoTg9z8L2V
DW3NgvDxpGkPGfaX23Vu2UtHmtGJLrr+RTeDfv95gFC+qfErw3fujEXlVSsh
v/R+pc3ZiIiKLOVBHuTlXUHw+BClbTlnylDQLsbZuGlIi259SStFl4SAKnPe
5DkY//rhy1U11Q2SVTfCd2wtCzAKGfLxIsufB/Wn9gEWsLG5BnEI9OOuvQU2
hDubXXwHCDvhV2O71KFNR3cHq9O72MHx5dCggEmWf9pkRsvrHW9qKVCBSnjE
0liYVD9kNAiwsjrY3HzoKoxjviGLEW1ZNVcWNdFVmOkSuossZXZJVLZ8knWu
EMqaBNKYwzPPIVN5Qku1ARiIFQyYXcBgkgxKc7wyZmuAHxRoZdeIwb7uKc+l
3nsTC6UpnAc1NspiuoxZZj9hVXUatSc3LlC0+rbKynjKXfOAMQC0iI9z6kuv
4f42/okq8nGYg8jQRAnB03lpvI6/ITyoVgwjsY5RF0pYODkwrJ9QTwwUJ4vS
IchI6IuKszCzNh9Fm/Ec1d4tQKLGqvgFgF8KFHR2D3tE0BgZHwFl/GQm2jdr
L1ZsJSQbu8+6HnR1cr3bYGfL0k/VEDntPkGCDsJSwmQ8nsPjpGaUZ9jBCPOY
5DqY2JNqBJQHX9Me0vwWjOHZ72sJADelNblVLfcrDZe5vaY/wp+v5c0+Hkip
Npnv+iWdDRQHv/yCJHx1w2zvUHSHfoh5cxHvIxKYCeSPfQWVnnJIrnLIlcFz
hx5SNhvLFaXma5EB6P8aIUylHyfXR/w82boXXPlPSdWJJLK5WOmxcE64nsBf
gYF+S2uP4v7mq5P/bNar5xOEZ20GgWwfoQYTltTuyxPtnqkhiur7F/VOig/d
I03mCZZ56cBoUDoY31YOe//C1V7HzeirnCH4E2dtK0OvDNFQYHoYADmmHVXY
02KiIyNejMNDOt2Itq8WY+O3CpUkvBJJyX+jyL3VI9c6pGw55lgOlz2/OM1R
ncC/QCx+V/COgGlL3j9LuExslJxJtORc5VlX6fr0PBvJeEFSWKnY0bw+99m4
tOV5Z7WgcfieFgaHonZbEWtD72+ZnKGtlfIxznx4c6wD2KO3H19Qr6CSB0fg
9gC3PybiBH9fLb8O19fMvhx9WZ+bHkS9avpImqSpieeYSOHGmEPRZlJPfa6w
laBuN+cAcJMpxjYg/f/UV95bv8vpMvCI6zj+MVgJ9rn5x793z133VN+AvYQ+
V+6k0fVb6Lg8zqKaUIFcXlIFU8kc9qxTXAgw7cGm9CCg9+j/vzNpLPCw/YOL
jmYi33ByEtVwqSmEGEJvvoz9zXFrXFr7xJt2FvEzjTeteqZQMvbX2ueUjpfV
vaBI4mtrCObAn3/25O4f0KuILgDB/4+HCt5gkZrjpHkCPs53sFnpceggnc/J
DLLY2TwceXCWxVH3eN3ENEy49cRK1LyOAYqQX4aiMFCtPLS+tC41d2fW2n4K
kS/aldHS1AJGgMrqNyAL40LVcW+nT/ETk7OEWrUsKfcBJO+5VN0Ww3Y29jwm
qYRvNp04B6Km11dk3m7V1VtHBiTjOGknMh9qYWY9XoZ03zKg7qCcOJR+SFuQ
TRwIAUjjnkfk5B5Q2VP8e9pNcn4VmVSWo5Iq9J4Pzss2GZvRzcl79/lEppuy
DFCZBD8242GZ5aFwhWg3NVcAfLFBhIOYRDQIT9GSbMMM8IM3fyb+EJXp0WE/
kjpRVFUZJVWiJpZMPTpaE7tkNsXc2SP3AX7U7D0iCDmgPWDHQGpbZk6X/aQm
yRI8qtzv37yW8QEAaXw8hef2PKsGIbs+hEl06iR97zVtq/FeQhlT6IxglTh4
310p2Phg8Sf/ZVz8dTUyKph1pvXUsSfGkrlO5i2z/AaPfavDjj8sWzORnly2
vuEiYAW/Jza4/8lhCh/3Veo2rhwu+u0NCvPh8EiRAnanDKIBfBKmqk8GRamG
wJtGL99eioBXbl+5pgArQfsUniBYsuAZa+mnHhpq7j8bwbRNZCKKDEwJH0xB
BCpiJKbYGQh4MVcAAtbRnHFRUSebiNc/qkhhpT5Cy0NCA+Bdqqw/Qlzw0LhN
4ob/UYtcRu+WXIbiOl/aaPWAQZiyIJHiUz+c4SVQyc9wcsanOAvxOw+V9TUH
skw0Qy+vOA3D3L+bBfN3TYWu2bat+kla7O9w3x6H1EL9osBM3hwsx+386z4e
exezo2KJry5rwAHYNHA3+1UDZJkEy5f7VJuR68QuPs5Oc1NKssx4xlNzqt1m
B13pdTAqL459nGvrdAhhTkE9sLmFFpcubM0aGTQTPy+pacFiCb8QXgRY5uCB
WIUlCkjLwUxBFmb1HLYeFebDL4JyqmzpHzcuN/XNkXUE2B2AbUCsWUs32LKe
xyjSrMBwd47SO7bj6JBZ1c4K1NmGDxD49Da/hlf5TcyZVF+wrn3LA4rgxzWe
wZ+TVa5VFOry2d979GUb+MGu38SPfqJWfbaWGHAvlTmmNVaHhn+ESBxCPHbz
VgH5I1RZg5gTe6Napect2VraKrCXt3hEBMa1TK1xdXnB7rL4zKMHQKYogeNa
e7or8WyF27xv9ZdtVN/6fyGp3z5dLHov6+iE5DAKRz0BUw+tJ9N6q7JJ9Y1E
mjG+nzirik5mH9t4pR8Q2Z7bUb3pFZDN1SxrDR8GpGxFMrR31Qw4Jv5yxZD6
mUO4FDzZwjXTjjefVje8h2iAlPmDyYyryW4trZfN6xh3QziNag8FiDzJzhip
vNUTAj5gZfKPoRwJSUPRaJim6GRTfU1tdv7OQy4idj5HZzynslKq3dBOBlcZ
eY0E2IUjCGBApma9ZlFSOBNH4LX484OkyL5BauXrWR+zDQ9xQQ33Oy5sAjUx
pGlWL4gx8RxAhm4mgXxBLXf97aDXQ763ffAUoxYiHOuTZDZKQaK6aqv8UIAZ
ugUhj8NOZVMOQ8kxwuJ23XMFAQsaeJiG4FS10ZzIE8ro8srilvLVHBixQqjm
v8cewAtHU9B9xwRdIkbR/h0MLETw4lgM4/ybNtTVOiPPNx5V6cScTJigGsTA
56VUxCCD8k6IXRcJswJhVp4fuW9mCqLyglWefW4FtLCpLbstbDnWj5bIkiuV
BYNDjJhAu1JOaLwV26n7Q+6wiw8ghAXvjhUutNVRS672knnPH/aVYmq1Ik/n
9MNbrhGc1QJcyfaI188mAFpvFvIWj1LEzfvrZxROrW3aG67H9L2NSSJxpOIg
CkoZw5tL2dcJPwzTXF7hlYEi/PltDYbIc6AkgGaOPoVUrWWGTxx4GO8ASRNY
4TWyuU7MmCTeHdGuYASxDpoSh7Myav6574OPBlRpdV4tuq/xXJyeMaMfQWI7
2ZDPP80zjNz5T3mivXYg5pvB14UO1Tk/h/I0Mhim0zpkigezPBn3PHPJiLD0
icaZbu9VuvLh7/NPfpDr5CsZejvTrYP/KXYMTiHIUPFLckVKnrZ8rQuD+PrU
u4DHfoVtwId3Sax3ezcqEK/pZEcz4+aYEFFcAKwT0y+NelchCeRwTfuGwLej
z0itemDMlrM5X1tn03jFoGWGbYA4teNPVfUxLFBoqxX+JTCwjtqPIxrMkiZM
QmnYO25cnq6QJs3BwhfSPCQquivH4MvYm6saf26mmC4ZQRV+mE2/Pf+uQDar
tc+OA0Ueoe/jJtMTL1inG4VW7lL72TUdLCNvR6aBMJ8sMQoxo8Z5z85DxF1l
jJuJ++CFdORfaYFffoWTGZl9LK1sf3B0RBKZEWuHYUkJ6oOBv38LP1sqiADY
CRFoUG5pdr/kfpykih/L7C0w7xIAoiIq6i+IDeZV8UckewT4urXHeKqlQcu1
kAhgupHAW0muRHgnDAg4Zh01cG5U0UbZT4hQtXcIKGHF2KawWi5jft0dqk1d
dZYcrRkE9/ATEh3NYn31nET8vZeICC9Zj+RYm51B0hCnIMUE23iQ5H2vJkny
HfcpPiIA1eF9zik5N93pT6pzDeRGIKKOdaEWRO36KWdx81BIaqHT3HdPftDW
f23qFHpaM4aUJFRu6lybi5kKgcuxDqyu6OcfJa+3iRfmL10HqD/iT9mRJAKZ
88Cy5gkwKJEhahjk7ePtfMY2L34YtD2f4DcWinEv1DdZqU1n+SG+eKaZsG5S
q5/pPAM1fCthBer47AtQ1hcZCXfQobMw21CYaAkjzVMqLgEzckQVuaMVl8H1
8JqpMdxUp1cBP0yMvtWwk7krB/vXtAvMvJ7AcuSDW9luM4UoIW95L/EKSoPk
kPUCCGisNYyR2/lkM8t9vaxMcwR5S8k/PpN5VlbTxi+V4I1LQP/6xRl4wAxV
pFJM6wJfKY1ZoiveveGmkWNKBS9v2h6svOHOEPieAnHDBgZPItw9wRHgGwcO
AfPNnrO1CqmKdwZlwUccB6X6MOCer5uJPf+k1SE7NM8ikBSGZsr4MuAlFeIF
oeCKiIk87RcFXZ/GjK4mTivfm7O3ifvBLx5iVgOEg+qV/ODkErhSzmbIkN5P
zLC1R3sv9Ez9HxkY/ChyrHED3d0KeH9T4HKGrRxjpr73MSQYg0e/e/sigMVv
ENE7Oih/KpxgcLUoV0Fr5cF8zk12/C4qK462l8HRCghZL4JX+ma0yr+x7ZjJ
pX/f4xWhrTLTAgDAoVP13ojqJMSgo654di8OkYqTA5CzdQTeXuywLk5YGeyt
xW4UUoBSc7rAbDn4R6K9HsKoc/VUm1Q2P6FYmSHY8XsipNR+IIWD4TczE+Wa
6KovmC1IAfbuKP6dr1tHOoynD36iAinXaVderX953BBjzuNEu+oYA/mFFBh7
WosPcDbWvHvKelZerrRTCIIVNdoSOn0ulPvAxMIYekM/McDbY9TurOr9f44c
ylu19VRvIewST0LX+v2uq0qQP7KekaNZX2nen0r95GBdtft1fbfS36FwgPFk
IKRNyL3to9cqOYmD/ozeFAjTevjXu5gIjThX+wI5HoumPxlA1aifGJhGI/cc
RATszD8vC45C4VcdKu6ztEhqvPpfEuTQSx0BcozoOJqM7+sAuxf0SHGhwMhd
p9HCjwuXEOgsg7p+9EJwhxqe8eJMQXbHyuigTGGrPlJU1bC9y2+BKemF57bq
mwlM5GAfJgSZw4qj6tQFOUPuzGva2hfey3Oy0QlAbbUwbBEI6po66UpnjT6F
aE+CobIf7RZ3WjY6CxyNfOImdvgnmYN9DhGZ0Qd3JVdpdS11nULzAUa9/+x1
84noGuPLn9RqQJ+wuhOS9kbgB4dsbCFcIxemFU+Gz94jw+0Z9ttCROUI1YOV
Eknnq0CkYkTzL/wDwAIhhafMvv9IIV56t0neSiEe6GQ83VBbRU1FW3PvYVT3
Y5TdOey/eFtqnJT2GzLGr1hUn16T9ZBbPrxCSSvGfouoDcFB3a056BQtI0lk
xvDTncaGZbD8EG6x9Rx1xSBh4yJ6e/FYq0Tn+umHMh18naT9Idc3DIlRCsmz
bRzCqzDCBQlZaWw88bOSOm2z20x4eCfs72YJ7kBkDLQz8sDEvmvVE+iu8rbm
DjtE+HAKLFov9F6hbf2LuZxdQvlUUsNGqG2S55qa7ntuKbgcoaWZCfcfjW7v
zUJFZ5X14NCEaUiwyBec0ZK1GJMiNF/6kBShOFplcybsEcqJBAzObhUTBEmj
o7g7P/swAmy1iVTnDUbk/AhgFbnuccfwBVPOwBx6R8A8m46DXtbkuAhLl+dt
AtmuWw+OURj8Kwxj31TnSNwJkkvOUGiYEhlh3EfKHmPOL4ZXPJqnjHNIYmfX
xD6eTRi+ZdC+6/ix9ZL/TXw+TSAudZkOUB1GH0ZbfimlFfklWjdD+wVMxgSn
DzDDBmF1je6qMS+yX7KL3mNvAjELAG8ccf6YojhqxCCHyiaZDsjjTqMrWNJv
f0zRHvAnDDNgwbYztmYJQDU/WtUh9QPq7pi9NF8Y6mj9/KxL/1CEbAguvlNp
FBdARJbjKCLtMJioQuxJ+JfqNvyyAtfqhSG/OAHJZPxWXJtONhmPRA2ROVeQ
gm6ssVpwsFqmrj75fZNAzXQyavZ7SRnOcCv/QugLYBz8C1wWwZhg7sgxBKDD
zfK/TJVq3e+9KYqeFeQnxExI0ACIWA4dR3hG2WOZWMI9JifAz0SQlsQqRUlD
+QUGrSFUvadINcd2QuZT4wkzGS+MyhuTQrafpnWCOQVAjP8rz6xlm+6CWVIp
BsViI2ffYLhLDOJKKaz9jKNznZXp7HLPidU1geaeTFnUdMdTKNsjTjMkjrGu
j4NquBntWsfxIL6W2/wOyQNXN97yqwfVhwpD8wKHg/Kebnp+yWYhETK9ao4k
bGH1hclXkH5arM3NvIx33jBO6KUeiVFv44/xBJVZukPd8AtkDUCU7fV/gePG
JQ5WlHe7orbqSm5dwZR/oQ/3vX1RDT1cMRLMu5PFYGkM3UctfHO9KxZFdp4K
xTr7u+bRq8RaWlU9KR5UHjhf9+C/G99SLqnb38MaL/wZH3gH7btD9CvcQu2s
Kpbwv7BN4ZgSV3vR1HJDPFENmJgWA0jipScMaTYVuXHPx+knHoTtL0GAWtlc
2EFvQ4Lvn5UearbIRaQBN41sXLgPV6piy8JV/aiBp4Uxc/PE3gLD1MDCwGFY
Ete1rW1U7WMc6ps9gJ5aCxRI8n6m2oW4mG6cxKW+ukombD8FAGXrfL9yS8FL
PFuRXBvi12PbCWednPxGd7bQq3YBBmgZJoS6cpQFeNylfEvngSH9f9aQWpMb
eYaGXUVv45nHPWOp1VDBRXjnhcyXULO0hRBforfSPvMaYpJ3JBiCBcrtFlNE
EKIXgoiVb6KdOr+ED+58k2ul2QjiNdnt5yq5eTAaZv2yEwghiJj04CwBXxW4
F/eAMoxYrhsftcEI2cHgkdgLpchvorANJ4nOSD7QREOM4Gmsh/81ZbaZi6Wx
ni5wmXUK6EhIqY4aBw3atB36FjmipfmgL02UsVn3TtiUpLZ/AautLG3n8VSG
tte97LzrQ6jocVZfnqsCb9FzSDhC/3V05tDL0yrEGEteAy26zW52XegMvvf9
mpO7gVf3tL3dalaZ1pY0R5UQI1mVvOpNiJ5tu8AfYOtUd4+xmJdjRSDBpnLF
R+RuP9ESl3cOOlMzXQ34uecUjDToxZU/HUoOXqkztPzVP4dwFeyugq1LiMzu
MzptJ+wErQw9g2hDBLYU4ECXYSMMFayRasdgpGJjksCBRMcdeT2IXR1+zi4J
HVQmVq+C0hbC0eFz1Qx+WHWCHSuFUU9AQj0NQFUWDmZI0n2WbuCj+jryiTVy
FBl0agQ6nYsrgaNDa8PLyIhE+lUXG439o1j+06iJZEddAiGf0XY/2m661MR7
cOi2vsZjgo4yivjaSIiC4HsVk8RJkfgTM3k5AHP3fn6OMQz7DAITDvcQ30WK
38LxCKUORGDHibnYsvsS8IlInmCb+DSG4fm5KRa089DOzAtXAMyB88k33b3t
vS71sKwigdm+q11/4hAxpqmcg1zyNAoJHOsRt7/MS6yeMfdMu1dkDswNeA/v
sys1jb9lSQsLD5r9Wo4YO6COY/BL41bkMcKsx0PumyvVUpTjiSfe8Eiobtar
5yG2Jemd7pgxWOzQCv2BVb3SHiK+MAqPMg1WIwQiDvq3mVTjuCoY/1s5CW8/
7Qh/gDLYZU1l1/zJuQ+p8DBp31szd+F50IMrhLmD5z13Tlll1PfANwQknYjK
Z1/BtYG/gfu2WxjGQz7auaj1SfCGVszcIH9apqajazHTj6j0gVQZAoKGZy0Y
EJgzuYLvl+Zf2wSX0EzHSNQ0kXHtgZ8qarN41tjb12zX8pHGqSo5GMwSfNoW
RrJQUalFcWjoHU/z7NNsNbQFD6gX6KY/DEtWxgkw6I/Tr5WgRM1QLhh0k0fj
y476rVzaHZj10stoqbqCJdp83SjB97AIaBz+VPXs7+aeRbT2nuecc7ToYIb5
qP1bp/T9hhIxhhVZsBKdkBGhtSjtMALDQ4NLxfAe6r/B1Hn1oMbzJtBf+Yj1
3xL5CA5XCmeSc2eikP/6WED21YLoytb/hZqgrKJyZ/HsTbC68aw6w6J8oQVF
wsOwVXC9cB8/jnDbVe1lI928jhTkWv2tSl72Tz0XklevO9sKUCf7pMPhfBQC
cGSvkC3ugX+giMojXhXfKsNSmXpfdrZxk8h4fG8YHgOCbDAk+6oiuwdXpYnH
sBZB1TieKifdUxSCd0Xn4fYgzyg1nqtuispxKrRVRtRoH2DuQmqDjYU6o9j4
RSjX+YzsB9AYswJAb+l1ays5ih4B/t0Y1iy/614hOwtkDQyBE0Bv8Ix/t2Pe
UWY2Y3YMPKmYOL4qkQgnVmCq5bSP0r2LocxQrG7Y6LOrSsT5r/k2/H1uALnU
PRpqa5RHmP6UIYlqJ0lt5X7I44UsYa35HvM7Mn7q+qFCct6e62OMDq8Iqvjc
jMZM3Ksnkrs5ZTHgnMtjEYsI/Z9qf3eLHK4QXVot/IAXGQ/AMAfjSGRk27+G
yFVnEsLYeKIQsIxU0zA8Hbrb55qJ144vimqIPWr0XDlhrEyufMLFG8RZQqvx
gmn6B5vgLTqz/IzadcXehgmDohhjJgFLCfSKI8udiObq5aPYK7Pm+r3uQSbp
ToSXvVF1WJYp0HkH+VoWCYUsdkvQK6lXG6hBfMcdQCqTatrQMSgEgSePvvmF
A8tVhoACdAGX7rNiI614N6K7gFkItc3PQhwCFpP9FX3kAj3f9ImQA9zbNC0y
iOyZsEcEdK0HKVP2ya6fBhyFqZjDzDa5s1YMbOjkiD/4dWKnVmxKMNXeC09Z
tSq7nvpvGAHGMijgALXdcSlGHjv2GlyZt+KUHbR/3+Ec05RrE1YjGLMZuoo3
sB1oPc7my+RL8Zn+xQ3QsS4qY61NOLUqvQFSl+3RuMwqj1RdUpbzcYNeBl4D
pS/0H+lYxJA9uUaZ/3uIma2P5muEgxJIw+EU3NS0JxHV9oQw0LoDtspNhw36
q/tVcONNrdL/yDfgKArJqv+r1QCExusgSsbB83zl5eGQS6zUXWkUlB32wEF7
6xFyEfILufCtZXpDFvfrzLXLqq3Y8rUG2ThmO2XghHBnshSwtEixzBCWmRfn
Cu/MD1iwGHohr3Xeyg46wzWhekHS/agM2fSyXbyi3lhJjNOvM7jYqjH9LWq7
1JC6RAIq1aWHpT9Ynv2DhNhBsI8OXvLIVUq9fhDVoYkqKNZfg+nA+gqfYGvd
nFrf6FjspZXaj9AkqUGYKy/iTsunAw0IMw4ycbn3DB6Kde0z+FzvDE37LPv1
Asgr35PuJjQIi9WfpvddBaH2ZHk9bHF5YLANj1ljZadNsCF/nr9BxjJv8UUs
AxsdfGn3BcVe+Fttdf9F4TZ3Yg6i5zuesQqPauTg/ryv8YAjFI2g6N6GZN1n
cDFmChF5bgQaBAAyQl3Nkrg65Wx9Htoj26hrQP88JS1k2IypQt0qa35tPBCX
4HQDHK50UyWuW8Z/YKeV12GqAh7603UYziO9xA3DBM13b1IzSfcjKPAIt1Mo
khuwunMyakstMPaH1HUL4Z83XFGqkpBlS5j509BLf5yL74G53GUMeFkFDgp0
dhnm68GtYzGXMAfIx8kib0Gu2AhRSGEDEZgcs5XH3lXRFPPTAq8MF5993n/+
vZtFouWqATuYWCcLneGU6lXzokTwqEh6dmKtasXYTb6iYNtgKgz3q8bh/vif
Pu3vMVxgff3ML4Rn2/yK72jrsKtIpg1LDtRjtJPVKLm3iYP6x1A69BMKQ+Kg
zm0+lXkwGjInaUZUIOpwzqfu+DXbescH8DAoWg1sb4BvP8+PpiLsixkEDzuK
jKCj4IqFtmqdydhdcghKiMmuz0iLB28HQMVbyG5OTNPTPpdzqYL/5rOY4R2a
dBlB5Qsh+zhP36OTndX8H9CddfNFU1/negMJG8mll/8+5iad3FzI+sx9X9Xz
x58CYbH5lpKcFQiJ+NLz4wpwcqyZuoHXFOS+kCDgUrFY79ZeX8RMHFXugrUs
5fCtkJhDmWHzDDha1hbIkn9N2dWfZz6mKDDu6an/lF5Zo9lafDJ0nUjTfOKy
s8o8fwSNM2OVDa+MyW8q8Op45JV4FQE8YKu+jTQwOw+IYZI6Gvy4Euh5EoWS
gjR0+tj9aD4DA+fJR0fE9rBfc0rlEjmTAxLzIzZLzBYAVJx6cjCzwnqZl5RR
YGNx6q6LcqeM5f/chA2ciP+lSzz+d2ygXwMfryEmHdWLe5vmndU3+4v5EYuK
pj/ITKOgXTGy5M5nR3yMUqKlmx18TPWzCLOjGC78UEZ3kPBEtpinsIKS1U73
rgpJD6Z4tRM0GCHFh5+gzqWx3CThPQex7LXZj4e/4n98WZBm4ENLlJRyKqa6
t9UfFSY+3Xkf/RJ906cHInkFujFlVCRvQ1yqlyFzmp0t6GJl0WmNQw0W6SmS
RfCr36TqxjM3uRFKmn2mA713/hdNNCY0HGHkaktl7Do3xaYFtVYY7hcucxOY
nJBuG3Cs3uLvx//jtVapMkCxRH9J4NtDvjmvpucm44hyEceo6UlYIvhsHfl1
EXLSPC8RymAMj4m5J1qpAfc+444qOWcd+lSYgJ61TkIo9QVZEYE44PDTK3ny
1rd5kFPHPrgEcucZ3TcZLhbKq4EcHn3P8oqVFHaXfBAKw/xN3EeKzzA9FeBj
abybPsgm9ViAWQM5lS8RrOkqSJmLKTAe5Rp4ya0UOHRbx6e2ypSG3nkedidd
swlfUAJi8wwK8LPeCqaYc7cHDLj65zQd3DsE721xTRq4NPHXV9z7PjrRJtHJ
+ahGtDRwqPiOs0vch4FCB4gt7hz4MDhu7S6HNU1oMAMlR28Nfr05CtXm7gns
9Wxsxei+sM28sZmIiyOsghEdMwSJaQHw1K6rjZ6ggnQUGz8ngTO/EN8wqS4K
gZwIH+cA90NDA2pRpo4ZKb5uVH96RMzPAoe+zlxqF0jMDQFofDgBT8/NCX7k
ZliKOd15iMFB/swOXaHrbblK/aVgbORvZv/rWhmb7xSWp2RHv5HhnIIdQLM5
Vaf1D3FHyThz/9MAmCSbJOUN7GihDcVbBjSWHR5vbxW/gJBp9TrtBENw6GKk
3EYbVyjRI6Ab47toLFjaxFpYDXYOeql737LMKZzfmgbXnBAzzTwbKipD0z9i
UWodG57a+QnOobTjkthMotBn664gemE+OR/0pxhGJURsPO9BmYuKI+r/JB0e
FHR44vciiRQrdfB4SitL8EJYh+yWCbi1Bff0+zXx4qBLScCpNcFadGNcwkYE
Nalj1U+c0EkqcVoBaVAwEgMra80LYNlJZyveFjC/3OVx97fcHo+0ZQDTEo68
zxi3pJTG00DjrIOEK1TRwhcxpmQAiuHXHF2CTE1dB8tZaI+p/3xMQIOG/sQp
1c5o8LoO4gcif7y6n2GX3G1WiZ/zSHcHpMc+13qNW9uLL+J2T8SqtqsgTd+O
W3h7TSvu1VkPZ0J6PswmXJxkTZF34LO0jfSPwxjoQhjH30hd81G1ZuqfPkbZ
CmfUFTlP9/+PGSYo96KGz63OyWK3J/i7RaSE34kwDOJXPhTZHzcNp+4xE6gi
xYko7tXhwMuNWes/sojt/3gST9fe1v2DjfiuHlAwej94g6aMTmw2Uh5YVNmU
MppCJcc44vjn0kA9fube8Y6uqLq9rzXb8TT+fMct8zP4h7tRAbA5bnGY+GCH
VUicUUEhM/f6RpumMIFigcZkiOxIXpoLwwvP0k9gVOZ6eGO+B9YqGAJYoUUH
zBMEBt2n2cixZ8Pp0lRbNj/usZI9TIDZP4DnwCtGDl3AdxmtRKWYDfxDP9yD
eRtUmwHmH0eE+amfjWHg4shgrXhSqjyboetjZpPMlKi1IbP0cV7C492yxYsU
RW8O9/R0IVvkFOTEf309mbfjoi0dSjdOFzxztQcPQzkMA8Vs7N6zztbW15q/
CV0RgL0Ur79L0dsuPQXIjntIGLCqjld/NAC87cepQebigaBIoXV1swiB/aVb
STWYCdVHF13dNXu8zMi3z97Zlk5GqJ/YWhW4TDt55W8sLNC74cYUquqBeiQZ
gfvdmoVBa9JNpcTYdjM5IkwWG4A65NjhCpLJ7zNrGCKDJO0K+eHHdhsLlBG+
KtwGQdNfKQJDMuEaXgi2qEOeiGBRTgk2RFc+YdZTKtKoGo11CFyCBawNTI0w
HEbLC+VG5/0j+rXEkoWSted6R3yHf5yett2CQO46kms7WynOSsAez7kYL0As
KP0CMnfrKPsYWuFN/DCssmLhm14PCzPsdBFYvdo1gsmg2DEJK5DOcdsDeK/g
KOxLbGRmBohV+6tVg8nWy9RdbhyWLrqVeyVPHOycRaiwj/7grn3vmsQlMyMZ
wgJhGufFQpKnDPqHzc23LjCzA72WV2tzcLqdbnpKf4hpLRcdK7EOuSvMKNQP
QRAzVh1/TwBsagbXQatAoz2VleMe6LdfqBm78kxS5Ie2j6PoE00VpC6TTT3r
EUdkD+rfxmbrv93XOGso9kefpweC7YmchwzwC4i1Ib6Kw1qQQhmXhp55XBUr
5eQPRYyYqQ3j4IdphZKC1iSmSC7zzqVGrl5qyeWtKqL0GVm6p7Y20mkD+k/9
+SMx/Oa8A2kvVGWCfFOW9LYOCKQ1ovDhps+r9Myal1CUz7LO1Jo5tcywMaUw
TyeAkhq9kCu2zQhrKEpsjeOoGiOLyT/9AYmgqf44+DYXuCteMKP99rh5ZIBf
zAJm7/YOwNdXAWfu7lTlYN6e5r7plSOitlR4p+6BAnWnCzgL0Qw2gRD+kXio
GBfOiLhi4RG6nA023zijQ4V5/AxagjhGst1bwBe7mqkqMtrGat0VL/HaSCGy
CE/+MkFtdBkN+3L4OhUAPtVobq8Feo2Nj2Yc+A7Pe/czjjWaIC3aut1KXk1h
uauXhCrU22OQWa3w2ijlAkqmFnhYkrN9Y9h+w5OeMPtVKfWnrnGsGjYGPmPm
7xHhe2WD4z/505Jyrxzki54YP9qMTls/bH2IET8o8v69D3ndbKLWEDdiM85v
73eTFT1m4RaUR/9ngFSkEg1zLaX906t8J9ixc9z2Ttpw9aHvdLZaDS6X5vOu
D4f+PkUTz/muZeJzEmFx8MNT8qM1wJKfj6imR2W2Tw0FOnBqJiFJLQEpbXKC
CcJEQmL2k03B3ke+SsEECU1BiGgGHv8DpClvALNyFMvBKObK9JzbyOMsWDd+
q9/AWCkipVASDnQ/HBW5W6exlgHS5xJXh7Id/Rtnx7VWfYygWBvE+2VMzGL9
39kigu4iq6gSm7rLee6edahUHXttbqSwhp3TlG+ZtXHZZzvlWfz4S9vt38i0
l1hHLn0vTNnu9vf2q3cCrVrGy9x+THF1IHmrJu2IvkJLDEtilNtK3saTtkhY
6ARSb+BIrsdqEQkjL6vE4AJgfCTKxaBa4vsCIH6RtRj2N9CwAJMAQV9oq1Qm
n8pZzoypyRfVfhoRZhqdZdY0qBVAVv3FOZXPrtSwa5cbUN1GcaVsMhWq+KjI
xYnx2M/OpfOVIxOUDKlCPnwmSFsQyLXds6jNrJOX3SvvZh9fW8p8K+AaEnbN
DpXSy9GH0bXtKQYDxF7Fj62FRyz5g0a+/KJJ8tYPZXRLKqu5WLw9rLPil1Vm
2roPxKrv7OPK4jv5GSI+hi1nmoo1dVZwG+AJAE309mAVk55robUJoBU0iGVI
O/AUA90qZF5dK+b8brroiE29n0iDYyKdD/LOg0OWw9+1aOXeZZTg8jKMmBe3
7SonBQU7DXpEtGjTchNUhuBZHPNju/Pik/WpfE7RN03ph84YuqpFSokHogdF
Xo2qSpSqrxHpWdWBvALh6cD5QgFDCGAS60ejeQDTTCzY06ngDpjgYm1LjyHU
r3HJV0eZENxRoTmHjS0SoyLR9lGmjJcMR4TbUQD0t28cQkdZwR4ChAWtq5wk
WkhcNU2bbQe2QgMB3WkP8pG4BsGhbHbdXu/1zLJSScD1cp48ZWDMw6jRKxyo
0D7kD7Drcr+HU8q/ZYvNamYfpBswCp5XjHpOL6Q8DOc2ZlyyKHzJDVvSvQjf
HBtl03OkYHLYSwNcL/cUYJytSxVzp+N4gcIb/CnwPC1xwWsw4Q+MKsByJd5O
OcGSdVqKQx/64VrcvP5Pr490Dn0JhxGsztIhVG2lj1lg9SGG3poWVLDAeO96
epTEd+MSY22IEjo+mTFMLP/6W8V1csN8/oYBjYuMUoGYsWyfc/3H81KF9N2C
bBJHrtipQPucBJr4pH0gmy1bV9vKcvUiYj5vYx0FV1PrWq26JfhqFTvZ1Oa6
7BSp2mDZPCvyvSvVGxUfJQkoQD+LkoA2jZeFr8xOkm8rpr73z+zro3jRbBPN
UO0HR8bltHw63Xy4H+q72Ad95h5ZQ8MIWBKTJEDYstytPOn1S2N/icjRHwox
bB6ncNAzpVosdR9H0vc+OMSy7RHHZx9v2aLIe4XnU3tRlB+ws8VXQsxuN8mC
/a9SZaKUwZnGR2TOXQ0n8iXwD1XOlkWqQb1zOqTia2u7fuglOfTPbguq1rw0
K8W29wFgE01VCkmGGSXvP8alBtWrDHvGL24MzRku/RSaxP26LVpaX1hFdFdT
IeLZYOvjEJ8G8Rt+rJ14VJacGXCJAktreZOXtKhcpFaT1+WQ3+wxRaDRAS6Q
ZlruW/uL3eYijKwrtqaPm3ms4ABm94Mwm00pgR1dNHPPkPs8o+h025dLpm6+
3HF6IegLsNMI2WzNsQS6Wrc9aoe5RYxDJEfnzuQKrmITGcHMLVMvMB8qr+N+
FnOeAVMyuA853HxlEpPagwRA/+vFis9UWbdG1SIukv07/J7VMg6n/fJj3Kx3
9EdnarXqS1Gsgim+240xmLyzr7Bbd05yYHvUW6q6CEmHGobYvs6eiEfTNOLw
OHcdwb8ay+0DcK9KmYLwRRRsluMtbouIHGQBiNZu4abzA35+/MH1K8v6qjPl
3Fy1BF1WAe2//YY92kZg8kEzLmH4eflpZXYzy1ns0wBB5zywntOvKZHvod+z
iyk0VQhOnhP42LJUAubGZ/3NATA9mND0Lvgx8pAca62JiunskWPUDfZ+ktnb
CxbsLNMcxB4eN5MqM5dzTvVpPcNdH2bVb7PRrlq5pKAryfVHKqE+Entwi6Xc
AzLr7RqyU4P7evP6PQwevm/2huQx63EpO629RDrhNOWv1BsVS39dqjEWo0H6
ptOw8ZPBBOpnKYPW4DGOuVMynjuvGg6WBkBnTnWb4/6WDcwvGHbDxt1v0w96
y40GMI7Z8NCjRV9LmpDu12avx73l+b0D9XLVfp+dQAgXmRTuCNeuv0br1vX1
/9oGqSKnzj6PaZxvat4BdCBDhXBJqvq7Q3OdKWmbMh0FOHT1yGFkXE+F0kmZ
0rKjIytKgjH3NvL3k2h9JwT5uwv6FdDTKnzB96RTvAoET0si209N9PlxzHVo
tCSykTxcJYULlQDYihHLmqZz4COb6AGRGSTsDqxaf7cmNVVrUEq78S9FFQaj
bUoSirT8Vc4lOLw1LPegYQ7zbXmyT2KTn0pYHOH4Zuz01OKv5ghOrg7z2BTM
0BPkgd9psxgCKOS7C6T62QEDwA6ruKCtQCD44UaXWIajpC59jIlfpuk6VCzC
Hj8lvML7DimMVkBr/Lhww2BMtpq1/Ccqp51tbezbyQdyAGDU5MksDZHQRhGm
1As1zI6bvUAFDNmZbGEmh3N07lyiRM+v4tvLN/cilOevaHJEQApZLvvEDt04
15bKIc31fAucvR3i6MKKwQIoqGw2K2+V3j+MFjjxc2uSGYSjF5Zqj+96C6El
0iGsJyHNTUjVN1HD5wn/fRhaKTMGgP419DmPKGABlB1JE5w0vg5rpPWsoBqT
Rh88/8Cu5ht9Ic+LFdJGXdz9E7y6MsGmksVxnfEO/k2Ej3Taj9w1oG10vtcm
ZneXVdf25Cgwru9d8Kv2lUi8NAEetzO5NlkgvDtX5B5xsLCU4zgt2js0vDOH
8S5Ct8aiXZXqQwV+K5i6mAnMIGdo/l4LlOMMlE0TrUfBXkhhf0pgzJS/UeHC
Zx2EfcA0t8CGIMAXf2eEwQbSOQZ7KGk7N9YIEt+tAlaPcNCyozkO6377Wl/H
iqRVWoIgfjFho2C9ebPo1K6aVtPdZkl7Au9ic7F31gp5ctzqSLBrLxNgpPtA
5NH1wkuQVqaWTaroki2/Rhk+qQvvhxkLGnm1a6W4G7xP5vX3oCR5cIeBA/tI
TxiBZBSW0RC+lWUX6DAVv3iu47KJC8XeVcKLqjc1IYu185GFMoodoO5dnzZA
Ye4q9OcZk0hX8ENegMQxwpND7KjhnSEJwenLOXd/vM4P803KO5ZJJdXTClDS
it6KjGeYHlF9o4nBJmm7vJprLrO7kyxNYDsZrbBVz6l7DbL5U7v7EFR5w2Kw
DY/GkbyTnh9T2Ezi/UQSLhlwTfEitJIpqvp0u1aN/G4FPGSWmWet+kljML8Q
BB9YcAtIpFzHUb0VeHym4BnENWfh1VqjZAOJ9Nr8cwi2dYULl+YCJvPth2On
vErAhxGB2bw0THqJ2cMdx6wgX1nVhKPIjSmZDmtHSfNCzBYCROjE8RR3fogD
s76ve6Zbl0hPk5ciqiERCBaao3QdibcBTXGzWABjh/62HgXt1e8lgOwIFEXL
uq2Ohl54Nwaiyz9L8Gwx8bASnNPxzqDrdWZVqtIwDFh7s1b6AXVp31/h5cLE
z5smawB+wj2FS/kbDh6qJKFmdJjvIQsNaBiEa72tNOTpP8gYn+06yvN/+F+B
GpNOhlZrtztPMtqscMP2vai7myyAXPAFKGY+H8Gu5Nqn92RbKQoFb97gknEk
FZL+dA90H/+SwBcvpEzAP6pU2JHwSqW97466z4pMN+c0bkbaWan07XAqw9km
WsJ6IqKYdDuYlTzecGXa4qdQOsreMcupkiVJPFx9qZ7wPkB6oJQpN1lZEDWM
xXjplOl2yMPcg2EomVICidriQ6fRWPeW3HhnS61gq3EWqkQEpjHWgtrcsGGw
a6u/9KcdvI4/090mg2t9Z/Qd6Y4sy3ZpgiZ6RUPbvvnbCcN3wsU8oROzJ2mu
lZq3LHwohcdkzIDTREWUH75FUELbg7CPVJo1wetioZkKT5qJBe6cFddqFM3y
X4Q0tWmYQMXyk+Y0fXiuK9rDlEjkyIkmIrB6aBwsPt4VWJA7ZvQNk0L93k/7
qc/ZRjEfSFqYDhRm+8tvkpeokTs9JCctBNyBz+ESE/5EwhPdXsOG4MjAe+3x
Ln3bHde6HW6xdq0fV+nXm/VginX4bRebg2ia442CSmV+LH6iJ3+yyLA/HWnD
FtMRRpu5NnvPjt/Uvw8HgXxBGRSKyg4P0UlLSJkHQo4Hn6cR3VeKUR1FXg9x
E6oRutkH3WBNL+GQhXV4xS3u+0QReQmMo9VxokkCVS39pCn2oPepPSfyD3g7
B+TkwaYAELPtenLCl9WGkAg2YG7ygxwBMXSxceGgROZSxfO8n9ipKQZ5RBJK
Ou2dgcdvXEswEPG8E8CkvTkjA0lVFOK2P7PpqaE/H2WAv3WruzZkmMhezkJ+
24T8ufEA0dgRQFSQluvQlDi0sr84/fs4Vss1xO8VJcxxPnx+fWDYNk29fUIv
ExW6FmO5S9TTKWr4sLyI0kq+10prZ6IlBuMtbVYaWtbQ3MEZRPMPM9dFLeqN
HK1A7CTscA0f4uk2frBilkwqnaL2k7mkiWo4mPinkFEsrGOKJ2rRlLacoEfR
EaFVn+yFOJK6Y6OvUQa4u1PkDvENyDJqgohIOUnwt+Z6w22z8GApmlJ4SH9q
wxed18gTM8WeKldSPjbU7FTL0v+mWeI8zFe9cGS2P8A4aCINmbEJhspgsZbf
4a4WtqW96h2e8yufkNKLu+K+1tVVXcOUK7Emo1zIWGcouEWv7qcPyRCG2g1k
BqPFvHm2CidfsjZtd+oAp7emWncKyRCCSoQPcXe1OTfpUD9h7Q8aFi7wY22m
/fbPAdq1xQmt2v6Ej1UyXlwCs5Wj5RplbnQFvnQn4ZhD9rnvvHgxELC1H+nI
IYKW/yAgEduN26MMHO9U7+oTwM0fLuLakl/X82wYuGuEGMLNPKNhntqMv2jg
/8wW1QlbinKERi7uwTHF34Eyac0EkoMruDBI3dQ5zqMxA+8U1FixqUz+RQH0
EW1XbPFoh8Yeqcq/m47WNIit9vSEUjVDvRzSYscvH6jrSxcjFL47MPRrs+K8
T4PPK1rSHSRwndzyZsCruPrEvEmT7LxIg/Msht65/CfjV9c2yQUI2WTyine+
o9gOYY8vrW54AA/kyH1jewDOd4/8mNuTC4HQIP5GdvnG5NuWKGKh9MXSlrqE
zUwU9hzdoto52O9Hz1ZblfsCm/QS9urFks5VAh6KwAbsvyoFLCZWsa+jvQjm
u4qySksRy9fASGfiyHiyZwN2iOCdOiyqVwyM5fxddm+59neFFbExRdXdKgn9
qUqmduhqapOtxCKXzeh5zYt4kIwQUkrO+CnEKEDCIdyATHCKXg+eeS+lUsIK
Y6CbWUbI0ICmyl7zhfl/4KEPIE7LIS9jYAGjSb9u2x+WqEDh+YIBdxBROOGV
cJJn/F6R3Aqq6uicmkNfOyi3ryG8Cmz6yzKSch/wGRVBm+hA/9zgrdYp8m4+
7zFDGUenKyJce9mUIvHNBotyN/EhllINCPdLA+ohAemmZR5wBe/loURxQ6lC
7Wwxus7q1V/RO7PEPt38Hrsd4oCeosy8KYtyepOsBt4/z5C4U/X4HUpKg0uj
mvlSoOiDYTH0FDKyFatqn17ac6uk4atRCByxnRHr+admGWA+vbzMpjEff8QK
JPtiQNK040563TLeLymbBIOa3ZNinhXNfgpIkknMpFIzTVENv0+C+SF9TRtF
m/SvqLoM7dbmGNl4ZohBoIqZm4gxVALrbG0u3B2dEmsEXomXr0rCMhCtNX2/
Mn4UVBY4PKztJi8Ggi+w1V5gl4kt9KQLHHnBE1uVKYKKzYODJj7ktTEj0ILn
OUiw6ruAhYP/uKwyr22veGP4K3plOmxXg6Wck7bo17WfOGtXTBL9XelHC2FI
d5YEu+4v1/CltTKDRz5hCi9nB8Tuo/GrQBbBa65iQ1ipCFNoOeGMeAV1kgt+
jSmtGuAGq8XF6howUp6ITw908RQDdMEXa2o9PWmf+iYf1O9ZBkjigEI6tRHm
Djb/62NqrmBW8uDFLBIvMhZ4KbqLTNUk0zsh0Xt3XCsY/peIHKxRknVahlNV
vDxrqci4Q42MoqvQlzAi6UttPr4uNbTU0uOWgVm318fghYXs4etiYAz8dDd0
bXxau+BM1ykBZAFQBPzeT+v2QKnMlyIWLICIB866eUIImweYrIwRxgoFau4F
QPmThD10t18IqwObx0Vdx2qtnF2zuhTwRyGSKg9IbAh/Y41lqPMdjc9AEuNq
bWRHvHZ53CnVxy1qrmoLnJaBCf3a6Icig3Ww/Vn6CwLTGaDVXWgoe6pAQGcT
TrNhyDmdsUjos+ZPAn8e2Szx4MhGnjR2PS+khBVfHbiGErWbLLj3zhYlPO9/
hBVrXwtPpVESlvkPeBun1Xx+jZkrF++kk68YiPz7WojKt93F3Lyqp1T0Z5mV
+gvOhlz7VOko4ma6dlrNnNqTSHyOMompPO40qvGptK1jzRsAaoJLnLy/3KVP
NPYbT+mc2u8JP41qvxWI24KlZnpNDxPM5nYCCLEtblU3/K+J2x7nIPG6576D
fNe4G/UiaWdcVybw+7EvT2Lzo6jejO6I8i1k767BezBFT4NO7J4DEesySPxr
EnAxhqc97Fb6HCkr5r41IY+ZlJz6ObfJGewrBfTCCt1+s/lxqWQsNkmsocoM
2zn4oOrbv7NG1i4BIAvb2WAJ7MKTeqLSOo13Xi1rBRfIzCocdVg8NgnNnKui
LlmYr4rW5Sidx9xDSS18eTqWogM4sOoaeLJFfAaMU7230EJYbwanTerwGmOM
hiOd7QDQ/5Kgk7VFqRhE/+FTTL3UYBetJ4tq8oUZZi/DtTor+EfjY4e4Ww1w
xmuc4e6Zb2FzVE3yyMO09Ty7fOZndw5nt+GesVl8oE+LoEIMgZly+kywtNck
iV8zBg+YY5gtPy/kkzKcF88HFJ5lhhwr8KepOhhAl1deJICNw3jVe8inmxwj
U+58UKiC957Tz9KbadJwtMebAOjSb6e9Yhc5C6ykzXwRgAs1kxroDalbnX0r
XlwzOGvHGDBis1KTQ6DcAzzdWKCzB8XjpqpMQ/nT0GZ+GOZdL37C0vb5roYF
eXKf4fJnhUV8SyJkLXbFN/XzKaZ/bxZFOA+uNsdmSZLinalMrO7BTbQHXCCt
MNVH+W2IXj0jNCdiNlGBSSfmVzwgq4wb1BmwWe2Lpf+qPbNZLwXOXNmJAfJX
PVDuPIl7E4nEoyw6nQ6u1pLHcEWid1GRb40EYHuWOm4204lerkDjEQ2gzXYA
a3Xp6NW4hUTFC6W16seZorOL0dz9FjbTkle5XfNXUfDltSDvaZH3rneRPYs5
1d3X3gz9xeWoy6ePdEQDP/E3Zux+Bt4ZTiln1HkrSLOaptPC4+JVAizpjNUy
6iHlDz//YPhseIewBcfDCX7NDYk2DZPJeyf2a3i+HaZ/1okKusJ+qyF1KzfL
RO1fo0AeEnj8qsB2H6W+1/In0u742+v0FBkigNye2iLuTO+hwElihv7+iuIk
DkSB5jux+8exb/pXb1KJzEHzvN0KnqF75VwwAOCOq8OgurKacXAKgqvF1jzX
+JkE+BbkA5CspMwbu6kPbSFSPRNFVR5abH2W2ylfqDBPOfWrPWpDUd84srvi
K6P2R6nzt6BgPb819U7xL7w89h1mcrpNQglk7cOw0A7PlP9tcJbwx0MZD68c
XuGBVJOcViHnzDlC7P4v8tKV8HyPrxBMghNEqQbOGKY2TK+ebPxaRvF06cuS
HsRqp4cxr4K2eubX9dXkmgRaSt2Q8cPl2jr1+ffA8LvwfEOx9+disH9PpND9
UzbvnVioF/JaGF89GXJ2x1zcP61qToAUZfn6V+8L07VPs4WQFwFcBcWjggYF
H4TItw0J9b7rCBsmk68+cblw/TVyB2alUuAfAh6gKgtihDUnReqSOqNMHOae
RlxIPY2hIVxgHlH2Z/TZO8RJacmK6hrnY1ZGpzltgEtVVRzWIubWkCqoKsrR
C0xQfv1Z6vFxqenK5kmDc1MY9VOf7otYD8okx/mp08qwMI1DEHwx++UxogUM
2tujBInkwZibVeyx1vTyZdfiBZD3SAUYJ29ja/FkhAmUPPft1rz702mGQKdE
kbuyu8tTMgelYqC8amO3gks/9HW1RmbclUq3p+x/uJhE9QoX0XB9GmhGMm/1
VfQ9+8WwcQM+ZOVdsZ8tAkZXvX2eB+Z+i/E6a1+/ieTiZg1dQpUEQzkhFO3I
1WsK3inL7UwsORv5w0CEu2roag9mcC10EJuJcKryId6dNKh92TH4y31vOHiM
pXWjm6hVgcG3e7pnk6PX0l/Gnha7cu7SnlVQyIlvh4I7t7O81rQ9tpQpuhev
kh+Y4sxxPuxB7VpCfZ4MSN6YaGlJq7wDELCx+zKwjQWJHlJjrOYL8t8qd7ll
KcI9qkOAPXZ62n9ePLMkwMnf0WEQ518t/8ufehiB9rcXmlGILMUHhDZoSVqw
BnR4bgySux7IxZWiPi4ZEW5yQTkkYcIKFqBWYniu4fYqQLw2l2Gu7ruBB4t1
lXhfjwxWUSsZz0ABwFX6LbzRnVY9clD1n40dpB3eS1wWy57GNZ5t5tBzS+fz
90dXQ9UHhFIJK59WA2pSY/w0yYP0WXMCy6okF362EwuRpga+jD317jaLwp1Q
s569Ds4PHDTqrqLzYwC0xoLqCt3V/zCqUhzoT4xcCuzpdh9SJLEGLotalbc2
5/g3EvuYu91vNxN3aTc9j4K9ng2luE61nz9jg4bk2hPu/mFTSo5W5b/HjsQJ
cgUwuyvesq5/apQpItXAO4d6BZt9KQHNovYw5LkdT6OymcMjRkMzAY8n3SN7
XL9EHfTNUixOC5eVjzaB43jNbEFNLqeVSdKkXhNtxqD5LP2vTN5Ypyb0k6ba
sgNmJKkQLLZtbyNxEg4dfmMRiRq7B0Ixrcr76BK7RiwyhzbAColjBWfySKo6
XYFrOIprmyyO6s21NOEJTC9TrA4yXMoJmMCFGLvVxGKNPwRkuEj70WDOUil6
fcSXGxDZ3I6T3WrcI3V35QDiET9i4R8xzKzodX7/YpspVWozwI1Deg+qDx9A
aWSLHlxo0VfLL1bsNrbahKQCycACWUXSNg+3Em1E0Hb1zvyD/RBBB73dU+XV
3MzA+vdADANl3XALYJzbM3uF/Y5zPfkJUoixKl4vLYDLAtmbsDoVEOS2/gfM
p6AEzCiMYlZ0m0DjT0m05/1atgC8vyf0mWjnc6giLuXK5LtQP5urWWXMiltg
1NHPPKjdiBJ1LMoZo04qgarv7dd/L0M77ChVepZSxJggOg/fxaF/0VD1jgro
J3whEte8172tfHQYi9O1SfPlyG0aHvVw0M98MJ0dP8GLDd9yjmhYNmRVlgHk
jVZdKMqS7/bKm74GkXYI5Gq6vIne0m6ocaeTBqUG+anCnUL7Ii08Grxit7uq
b1Y0TjDsiNvI5AIaXKu1hsyLaxCIH0IkjtQ01AXzg5XR8mgDjIfK2cN8VAMy
IjTKF93VAPsljrFE70s+iKrTKxufHxYmScC7Sc248GNOWWQ88CDrXTAnzwDn
yAG4CfiHobhXYuJPEvA5QfeYE2n+8tkYAzPH2lA5aA6f4Sn6pFNtyZKnNPpI
76URLWxKuxmmPp7qxmmOgYE6rcg7PEPg9X/futluJhkxuSHymxiCZEnjHLKv
Nq9IqIt300ADBXz4OM0icJiHRDbdlSs69u9M9hQEg2hf3Rvjerk76g39lEgM
1RlyiN5ShJZAKzMaaDYNANKlmnbc/qBYcR7q/W9EomeZ88oGoyt88pMfWfu9
QUw8AYqw62+I3Pj37e/bsRRlvNJf+0v9AinNO4HXtL711fMJDYLOLt5oAaa3
9TXXRBN9nQ49CzNlSv1jsi2ON/55Z8p/5NU8ldpLLp4MhC/qQzk/+pDSvGq7
xsH1noSn2yC62tWaViwGwPM9HT6ak55d2OON77XA5XJJWX0zA3YlpUKqA7Rj
3rV6N0tzUqVqzQDLfJoi0q+rkQG/gLgOhz27kIVUUJszN/4zHZy7JrS5PwfV
ZpaG/iNEfDxCyCGR6vsxrzrIZCummo4l9ufu756vrQh9CmHi6I19dVpvGVnS
kHWyTOMfWXAt0CQ/6givesrQ6a0f/2fYHPncSMGPnrLW0wnHoPwtpKetm6Zs
JpMn3ZEaj+Eocgz8rXM1A0v7BsCQ9W4ndvNj0ztPDFsHJpHXz8vcK40WzE3A
PCVtA3VQfy4rMpNE9BHGJwrnOURPZutFGyslWFVHJeRRKlMbcoZ++7lpbZss
0dMubQD4i8vIZLvjaw4IjkOcCf0YyTrw9imG3QbdxNL3QpNOH579/JXPP5zE
j92NmZhwXqfLsmW8wRuv/LsKStGMOSWHW3yLIITtaLG3suc7iJMRFnCC3OiC
BpWG8El2YO0JcCFW1jdNK9X0uBRTHTAH+wpAQnVHZY3rSPN3R59jy6nqtZIH
CgEx3bYsgN+GUK+WzWENY2/AlRb7zeTaJ6mdbQzPJdHnPvib8zepJe3py2Cn
dJi06+EfNV7SKehARsBYfrecZ3VyE+Xg9crZxm2Yq3LPpeXBUBbU0icZ8n4v
kJN2YcGIJsYIzy4hFWsTJVyrJwpc+COTPWwvfkX6baff0VIQh9/6S/hVoTol
3aEo178leO+ANt6JZIfpHU7J7oapm0bPtLFlihNtGM1iJChdqYvc27ds04y2
G0Mb7dLivO47EEjCRnZziU6iA2T6Vzqy9u/52m6DBzQ7h18qTEeJE3G7sCYA
GpBvCpEiVOAHEArSZ7C7piGGc939egG8Q/MZyiLsCIaImMZsPiGzELcOZXmi
+qM0g21YuBr24kmaRjZ++Ar6jazfsPzojTcwDhJJrCRHQacKd6S3Dguomii4
U/533+bYroDF+E1pXYLDeGwUg2jH7GEogM7Dn4HzxhFocahWjL3pTygPPnev
VvB5Xlc3tVbWBK6f3r7XlxO8qMPGFvEx4okV151yJrsir6eW18romqW0IudT
bc8PKz0d40+4A/WN4jPw50vnoIjqmkPd2f9QKrNnhw5k7jAMFTkiTxAxpGg3
2dBTW6W7RyxyYh0jiEP4h5vkIaqLVS9/mIOdOPzGKOj+ZAiXgN2B3P0Y+WDG
s2jltmkI9jN+smo1AytTGrDzPJYPvX/HSpQ5BL75kiITk5JcVAqp12Y6aGyb
pNG7eCXUaXNwXiJuVaY3nR3H0650ABu9KfoITZBQ9KhOeLCKT9Vk1XIYNUiE
iCmbSokDGdbTcAJXo9iyAHSJxh7O2zrxr7zZgJT8k522a7nz/TGZyV7crSw8
sI/Lb+TjIMspep4012wL6TxoXq5mOCsqO/+Kroz1rqqXxrLbHmdgjTPq7LGi
+IDKIdQ1eq8TFlAcZsZFWNPv5AyVHu6ttsMX6z1kyJmQi8OWr+6axYNQ5/i9
YhiNoAUBcwAdsClGA1MM9lpLiDC801M6N9o7bNXLUTpqzCKfFBezonNSPAc6
suG0oUA9cY/eQxd9SIqdp7Ydxin5KXrKT07i2Y01rWHelJwXVHLIbaUw2c1U
zuPnKnRkIQjUWj08XoqeOrqxQaQJbbpC1dzz8FKC8+CX/ce0EuCcFFqlpVip
BiG0fX1dDOeSomnu6uxa7tOTI3fBChWH9KQTfmIX5p/B08jQYG8iKUofBl8g
nWgjDvlZPypLc9n5YDG7SEYqQG+ME9QP+ZCSEx9TXpo+Vhq67rUvhWjhA5zE
X0Xhx9vghwp0Bn6yD3HeIWxoBqBG1Lz4D43ODo6lRDX0QuFhkHmO09mHRfE5
WyUVOeISl2FGK28RogpI+i8T2rBKA6PMoQide/9hrqh/gVmByFRzVfWaYVBn
ZCaplRbKSRUAfFrI4tgDvWdHuX7RnQVf8tEj1AL+S5+p65qsEAJ0weFNNoV+
RnlMWpytXQRh4hbUYvTmGSkg88aWH4clOFCWf64My9B2El3xm56PvVkzmCho
I1qchEg54ZKGfy3+SBzSb5vdYVBwZDpN/4EW0M11rFInr3oOXBhZx42M3VRE
dHTYDvGZDQkGIBaXGB5kiRzqPbMvqwTA1XY8nj+A/t4sqNMfG8KAgkwjsI6e
ObBTee4GsEsxrOU5dagZKmEeaIyvvvwqKNUDgE8depnLSEPy8H+gkf0woHuj
I5ZP+KQqA6/CEJY6ff7OubTmEH9/cK5sG/jY9gmijt+ha1aKS0oR5wNUUsi2
z6BKCCuI14AYDYlBvYcD4Hzl0g1RboMLVzQOG/Xk9uQjtOcxfKyuLjAU69eP
eySKHKBn3DBUWj1xFlvuovH09cy386w4quMNbPQOF16V9Mkw4Rt8J10gx6zs
RlESVSnMhPdyxNzumY2DbL7277o0U2gLJIs04vmji5UTT5bYVbDGfX0QUSH+
fwVpaPefY2FWrYrm6tX8B8Dor8rIcq56agRddL8o8z7EhTmbwko21Dp8TTcB
j2siBrSWbQVh/7xLyW2ukJvUP6QRYIyTKgI6o5sNr8eId9JRpvJTWEJhnUB7
ivnP63ElTDIt9o6YVtkReOvNd2g+5ncslc90pQ27gyVvZGc807rP4Iif3pjJ
qc36Q1easEX0o9FDSpkbgUTwvKVl5jFFiSmPN6wzEADw5kPuP9xf0brJFSja
l+dE2Ix/YlnsGzH9IdwiV5ysHxLDA30eDWUsq3/xgB3z+aCmRi8Vt7B+8pE1
+iV91WnWoZLU2bdYrUFJR5rKIGKDjdbYUeA4fHpK7qib5AHTt+qSYKEvaa0E
fYY03q3G6iji958K+reBbOEU7+ViJQz0pz99/owtDcGBpEF7acMVtna7ysfu
ugyScNKkWCI4TeV5p/DdZqS/P4IZ5dE9gulurKDpT8DixFL/Qmd2kzhXpVA2
2qLCRVkrt5RqjmDDfqjFcy7QleZaMSx8vufW0zlMkjUwfnZWxdxStktBYPI1
nZabiqHJ0/+6dlVzgybpgR0Nl0lbnwpFeUzMFbjP4JxIDlbJh5Dl1IrdqcMY
gb2/IIgpWJFvmZeM3yGukdPR2VTl9EdvQiyeLxaAmkHpAdZclJk99vesKZpu
gyyaGJ2TfcHkTUnloGGP3UgJWdH8Ef8gBJJuYCh4gfAN5mXiG68AVPEqqLcA
b8IPlZ1pRYlih0lmPT4ymbc94zurpfiita3rHGN4pJB0PWl6ohhr87/rGdJJ
eG4EpeTzP7fiQpIwgE9WOamhYNbYJrDXpv60TijNLC6TqqaiUT0dXYnAxnJl
YQIbQ3/RBci87LuJfwFoLsy2lbjPMvdBFc+xinzyhxIJ3HgM2mWwRQVRh/av
IoVx2otpLMIsV1rB4URcz7Y/3c6OeTuu2OkrhzXNMI5FOwnHOwSPe3wVz/sM
vmnelmsYvGFuHSOsCE822g2taPv9OnS3p3vlRybRYzJ4zmglNagKrxzZLVTi
0+RmjGbP87QTneWaXuAZE1eQqDlRnCkLaoe4VxeZboszOPIFwT5vSpWYXoMN
tuJSSMcuzj5JyGithM/S2QUhDwNskfdnk7+UlknqOAbD0x8HNFaP50fN+amV
XUuHHfFSnWYoVSx0w1UeoQlQpG90VqB/hFF6mbbkwyLZUG31//OcAFs/LPvz
N7tmLV7gSxkZKO/d8nUrT87VL4WmQ1hw3pHLBOMT0ECXJnn+5HSuUAPqrplb
J1Nli9ew7BimQDixFJzkBPGf71Ub/vSl+acQP/oxRN4o25KpMQA2wC04Wlc9
sgQnOmDmmt05LoXgZvHkyxgUUdv4HyNX4IankRXjHttroCTESNU/zbDg86QM
h8k2YVDQhqadZcZIi0iGBZfDEGyK2GMqYPg29wTVeK2TIsyew3hz7dAWykNe
1ZqE4pOdbS8k8D0f+yxSemnMhAT2lTbjCTcJJzN8/hQ8Jy0fHdZUi9SmEGMz
IojVItilYi0sW+jmnubFoVGCedGupmp7Zn8WGaNljgr7HXmyGQcBRGwEg/17
VPlydbQg70J3qb0WiErbeuawCS0g0JOHrNgfmD2m1PJsCsELsH32bTS0zVYk
9fnVZwcDIQBIgyM4+XnU5r9QJkmS2JCetVzeVaYIMFYVCMq/8rxFc82Da4ql
VGZWM10ksf9UAuRORThSA5t8nW4mKF7TLo4LzbrD9gdGJaW2Xpi9Tzz8tORf
zXo73k345TPfvxjrXgj5KY4Rs048SZR1F/gtLzXIcdv3occCto7v+rQHSQPc
fJdnFsl97FGcgBprOtYiOzDoxuFiYZuhsCr4YgmLsKyqZUTj/KpXn4uSwVUd
9eSBASc5epWxI3zLosU1VB/5G6vz8ckkZx5hImYl/4jR29mNoINoIVb2Xkp5
SBGL/nYwqcR5BtsL6BYLeG0X69hIiGN0NK0WmCz93OB6ScyK26Zc0lzxsBNW
C4OL2nHzqf3fCJFBHcsysP0hDaWUxmtgT6CQmWaeJChNa2WDp8nsjoGYVMlO
PybxYGcKOT5FpXTrPS8FK0e0HT0F5A+I6bbYbMigwfRoxAVke7BEWLisilJM
7BKhVK6hkpPHTuK95CAtEOz8bERPLRHFtIsZ4ok8LjSxmCRHGsyu07fa8Ag5
AKZ0Bkfsk0HjoRLlSl6vbEb5HW/N0bTOmVQe7kGKXYuxK7NmYOriGm6zyj2T
gnE8vAkVVr23rGV3FI23XXx8iosuL+kptW+Dp1CyiantRaDe3Enrj+Lz+Mpi
S4Xgq2/hK6rq4YwIpwshWOgqYLWvHfNCxNPsonHcpU7GswUKRf+e2uILszSO
sers6oe68drWhSe5If2goBXILtoR1ta+08nQWleLPOpdcfKAxLng03d/vOVo
O1DnB08Fwys5Kos8hfxDPkaufEVygQnkwecr7Iy3xMmD93u5rrquimUtwz++
Bt2oNDPDumS6AXn8IxZWmry8azUCFhAZIoxotMr6/jeDccX69EcHs0q/nu3c
QqyOfWb7Y/zOxAKoeOrafP+gfgNCjoDJ4foIvghgypuOu5QzDwfbTcd4qZAb
ipJrGJh7l7gjH/zoafFbJ9SeiHjF+a+YglhJ+Cz/LwgZqbRsORx2fGPjGZBh
HkuNgkyO+JJ93ELgETpn8AJpMUa1lRId0LuILbRR+g9I4hUcrm6Nx3ntK82w
mNZQRH3iohyxvkJy5Q3jtg3IUsi6qbMjt20Ar4U9QyPLpNTjLGLAsDF+vC5K
FHBGHYPdaA4SKXSvUfKTj6ZRQLv2QVPpn5Xr4U5GuOp4/VECP+LofpV7nXBJ
M2hDkYc2vrTsxF21931Yk6PZrtFhaynpSZsWB/7kQ9Bp3jjcB7p3Fr23HSPP
71a9qM2DQKmiXO8vuLViuryl9KUEyYoSbjdG8Oh/XklLFUoZ5kt0hJr7YoFx
zow5JkvNzdKCr+3oci7s2FbWfN5QDVo/lheizBEHlNER+4WAppnztw6/5yjy
3btN9QfuVRb1Ppp+ydy7wEeop6itetsL2jiyilJsveA6bjLao49reDtdfu2K
qR2dpT5fYM5j8fipw7DLUG1lrUug0qQcEI5OOdgWDiIThNzVz/8rRbrQcCkr
1sbdBT9c7pfXQrt+s7VrqMFjRf2ExYoeKi55VtGK3Z4UVuvDUUyJSPzg8nFa
4T/FN/QDwkpdynF08quxmVZiKfeZnS59maj8k2ZKI/rV+XSYiUO1TabSwr6x
2Ftc12XGyLTnEzatBS1NbE6sc4NnR0HHtrqYxUzN5S4o4rpLxBPoomkz+Xg/
KKOCs/B42xgnQtgb2ch3QC7MksQSa4688HbasTaeqAqnudRMsl+OEy5HRqHt
BEqYXbopOMcyOBPnFrF3UENqYYy3uxpVyBqSZyocFqLVG8Srm3E0LGpMqnll
CVclp0sB3r8rCWIU4IvnRDcuyVdPJqxQEvEH/72tRWeIgNOvKJU8ga8j7mFJ
HotQC4KTILblW9XZSeh8nrlLGhLWwn+Of54mQg8HlRjbMoMjvUV/0ZNtJAdD
pjVQFhbPYcIJuag3bnCXv7YY1DThd3pHE7BAVqhpYfsu9+ktIQZY6jk06mG5
Hm8ZwU+FSeFw6F7w0nEcU5TkrJCmJhPIAfHYg44U1+jc7f/X2hs2yHqYCOtv
71P6khobhNLIJZZU2iO7fbNTNAIBnc3ns62b+jt+5vHOFYu/HP+umGly07Mu
lnpU+LXkaYF0VdWw51bEuSeyat1JxUlUUVNSPHsJ58PgCq9/vTxFfbtsz1O0
9F05p+YPGcVBT4kZjOjkio3o+P20/6nMnlpHVWReUV9gUmZ2JuMqhptxldyB
aMKzF2PPI7uIcvfNWQSK+Hxu/tkiNAlA8S5bheYfIVXUJDJ/+Cqn9gZVoVC9
tEoKlqJm6T5X+CZ6PLTn76sqMMi0sBL7EaQ+bTm131gnMbQOU9/NYnJY7q67
MJmleO1Pulc2TMZJD/4BnR769aj4X8M/3W+6xcoQgkRH/1it4Ai18iXUZLRu
lbieiTGx/Krvt4Q5o1B+iNuNLhNaX8vJCz1R+rcKwdraxSm99DceFhxvlo6C
sKEEhSgjzT+BKTayztKu1KAW6L5JAW7+IUETowg6gc9xTtdbzhlDlXzChB7M
VMV2MTUq8qs3gyy2L7Lbx8D19FUMQ5eoQd5W6nAsHksyWMII6GV4fXnoakCJ
/00Ru7kMWbU52VqJVihQvTRux//+nZtV+UFqXnkFZT75A8MEBmTSf6/YzBrV
kEzvkMS2cIqlmfevxZtC1x9TyFEpk0CYZuKRG/zswyGUFg/pqNzyjWgXtswN
qVkeJB4bY3AVvmFN3ShP9ZxnQopSN5lsl6l0qF8UeOyyUZZ8DnxhlGxXTQ+I
/5ac8edLblwoR0VQ0HJ5CdF2avuogd04+K0lNIpreo64j63qyLMDf4CyuXfg
CBVJhNTIHpF96eJWZpyklCJStv5xi4wT3EWioNf+qdpYVOANQNbJES36z2bu
Q31LOvg7BqAS58QkQFaF34Pc2IsOKPIi61mvxxxbnKcGXponou+kRQqn07Tw
37wbObEC/lr6qIf4mCsT/aQiv99SoCOcL4IRyFzOWto5rrGnHv1gr86tVPAq
5q+gbfIW0f28nGI5j9mvy4SMTkZbdvixPB2g1xkOV8l6jbj+3wI4aUGjla1D
lWUSVAF4jpkYXvlWA+ZAkAs2TSGusOsob9iLc5esxmCbibs6U6bCBAO1qZrh
YHIeSwdcrUCvD4dXhMhztmlEdwMFsMxh+1XwcrqU4//n5KckS2dT6NedEzzF
Z7/jp4guVGQcJN9zBFwX8kJnS/2s6NJneYIpwZh53gyEqfGbKXbip4xCNaeb
VRgZYJsMDa6uNhI0MyQSHkzqFzaupt80yddXMZ7E2si/Lygc64THqfByzkgg
oF2FVsed7x7LeUwKjFNhTuw5rSBll3Cm6et8wD3H+7nuN3uZYkAQD+5FZR8M
H71hVeOnHDGv8+4NUSltDIZii9iclNBN/sF79Q5v6fKw1nFUY+IbE49eq271
plYbSyomVhVYFpW+uQO7HcA9ti3xnu7sVMxeINdqw1BebEfFmbyBt5/+swMW
4rOYw7odxXPRSVLWa3KpFJthQf6cpFr0p8kSbfeAo7Y7119F7Ktkl1TU+hsp
znTS33xAPl+bABa4ozyLx+TtYLhNxAvOchGKmEsgpurev1dFzDiAtJcHjYQL
ByVfrebF9lsfrQ+7ZMVRwaS/r0/z1MT4PVASWXmjN9Q65iOVUlm6M9LgwjaQ
Hfr87rjP5u79N2xb/SggDgPVd0h/oGLLy8EiMcXYYErNIHS83RbTTF+REMww
ul5HzrNSEG5bm7q31C2uhmGFLA1omE0ji9/l8JDhhIsFGbvsYJuPazq7HQMZ
yFQpF/uOg/YlHcbxEI8VZxDMeAxvZaP8iMXV8WQ8mP66YFmJlm8AYakj/A9W
NxAyhlByQ706f0QHbr7UkDjwEDmEmdDxzFhFvqjK3tiPNUfUchyyKsfULg8Y
SzF5JmwS3+Ovt0PXZVmauob/i8xGJq7YF7IxDbzEBExcfi/eUj2j1+4Ggt1z
D1J2WmHnEI6VrBrSda0GXwCBtwLMJkNEcZcRi9NlrYS8mtXI7SG7eFsszC4L
xhTfgW1QjraQGhu8imwYb1m/KVv4GJsha3FnrRVlqky06mLMSmUhWNWicjRk
4TvaXY1Cj52dGAmAxunRZv1WCx88rDHFAp3uF+EFO7nzz1yODYBCq1U/Zh+K
/s+DPwfoQu/gNxxXpR+t36N+ViJAZ+XhE/1Q9qcu60yUMhnJARAantEpTA+Q
/Qltnaz0HKw9h/X89JY5Gxq2ruSMZAANWxWlL95gMDBkXJLO9eazfR2cIKKY
oc+4svh0ACbfy7PUejlKA7jo2Mofa/vsUFVDQRnfyfOQ/BlOvO8H2ApgRk3d
VqOKPBYfqEdYmLB15h+d1/vQQ2heDNpdPxmxA+LM4IjRkj5tZ+eY6nx87V3V
/h+fBPg+qneiH5TbsCPXs1Rm0zMFHPGRmuHISMJuxSh2Xy43AHSNuhegHR5b
aMBmfRADkL85g4ov1uFVFOh+y+lZ8yeUvmH7Ip9+CkaxuWV0Rq2bgBpvILiS
uN4MubInE159wISaO1T60XvLZ1XNJD/qhftLjkKGE4O/O5h8T1qOUXAuV2fw
TV+m0Bj+5cIfsgikMSrTnTewGE0m1Mh1ANVpySnEdgYdi3BZ2PaFBJXXEWoR
NCl26wZRNP9WHkBx1T9AqwsZwOUaRCriq+QimY/KxuXHaYoqQIl5dB6pNrnX
IBB1DiaPoAKZjvUb7kC0BhLL2AB/CnQ6Ond2BQA03E11itf/ZHRwujajNECS
f0FBWxINnEs6auNRSnIjatLLmtQPbFDKHLBX5qZHfvSG/ynzJe7jHh1bke+r
o/ux7v7meR732dUfc5cndMRwxuHLApcBj74AbJ3S2e28xwAUijtFvctbDT1p
svRxSs6SHpG8w7y5dXshEZWuRFT3soLvkHBbaZ2azqLHrIR4HIoYh/wa901G
bWVLSLToduZ0XCr/x0U9Lu3y8zVteScnQTW8Zydgo1PsjREFef2LJBGhP/eE
Me2gTWpqpjWynjPeWzOI+IjmLB/K0V8VjhBygf/NkMEZZXlxC/keLKzBTmYL
qb0/BQvQYO4mTx/zQcIJCN1OZaGR0Stmz9SWQHOh/BwMOiBTqrp9Rq1KleqA
5D29bJagUw6m49Y/81mN1d69BnCljuivVMCZdn7GN3F0Y/ENRZIcRcNjW43J
Uqk3DEDtdHIMNC0nHGs7BEv4sz9RNTsRQajvU3smGJl9ifLOGYvJIymBBOFB
qeTo7r7Ob0bbmuGFDJhxeQVtCzJ7uMelN40fWL3yAuaN8jZON0bzc0jXK9KZ
qOOIHqARUvVDK+lZvjkWsE3gIYyirsG0w9DBMDeXfEs1galkBGEtRs7OOAmI
oixGnw5Ezjl2yUxJz8VHrAO0YsziTD1HTs5o/N1SNi2KU1y0WM+XtV9JS2jr
iTEXy5LdK2qXE6PeqsjDWQVxyN9Bcy2RRhMPWbWdJAokOog3Is60ngcKacUv
takUdNvL5t1LwExiYXJ/bRVBHOzrY37vmQlHQaOJW0WV57wS1gz1B9J50/64
t4Ri6X+GKzGfZruwhndTksVe3NQdly+laASKaoOGDHe9Y97V8/wfc/SWlTxV
vKbU4RfypT6s8hrxC7yddEpvDVv1cPJAhnPCxp7ATJobSBnOf+AdwtHoWG5x
inHSw+nLp4V8AkHu6BqxIxbf7yUdPAW9R1YuBplwVzC96sTLNuA+Im/Sa/4+
yljaBSlqFfm/eaWh1QPu1+/pSPQLRYwB2ludd/QlgmtrPf71xSLSf7FZ5EYd
PyDCL7h4bjFYdNgXo7KxwZYT17Kh4JntKYzMP9i+3d7cIUV70DBQ5gSi6xOX
VAXt9aK9zV0bi4CvK1daOGaxXHrHYOyWyofqpSnsy64V2KhWdIsyi0G/eU5S
zvUWKSaIVkVuKFrPGIjRcVMaffdfi864DtvAQjd35E8Ea4gYJQWiV65q1EtF
4tOrJEzJ6KG2oIoJ80QxO+gnQdDeeEnzc9J3FueJBXvNBybkfcobTIcioFkq
ZwQw+myIfMLg6BOT6NUvmzrtXxmWJLYGVTJ6lAG5kCTWmZTYWTEIe/SP4Ja1
WMKM62mlN67g/N0x80gIpLUTsiCriWGanURqpzd7nulzQIrl05pvOb/3Rr2H
6AUFtm3N3LctSbH1v1gT/io99PNctT8qaELjlOp99KCbY8lEaevdR6WN9WQF
9WbKafNIsWCmMGScqibUzm5eyhYltgU48GHZStq/+G9wtP/pNefaKv5DEx+p
zeTVPzfi8PoPugVHmUjmKfAZutkMQ4Cg9+RCZiSrEF0ARXtIpGNDUYNwkt+a
GlP2ltpSq8iMEkMVIICCvQKsZsbQ/qiytGXawL3wbm5DHk3pdqEjIY/YPqGW
xenlJor9X3GQOuETKagqRwLU7J4HpdiKy9aE9JNMFMNoE6iF4tuGuU4XxTom
HDEUrrDgT6+VaDM4epMalmIeEL4TT7UTaemVtIN2r8xmB/qcek7AfObk+Oca
KqehkuZ54M2qjr9Q+scTBgO4/lAVBY/VFK+I/1n0lv5y6dnXc1Izq8OPozOG
Sm+SCZdMbuhFzp70rFnrAFvj2b5PcoKyQ4ddegqsVD6iGYPEten3XahrMfDr
5/9OgE258bY3/Wu7xeemxigEjKByI77TxxbZ4t85dGoH3HVfITKAMzFgGwDD
6j84zt8/gmsKMlFtzCmtM8024kL0eiAiZJ0rOJDqqi83eXyRynx/LqBYrfFw
+E8qQEjweD3dH702y/bSzCOx2SE+zikBF463atH9zbEiFMmvkPFwxzquxUrA
LYIqHrZ4gC+Oxsv3VjRNgBR7Q6wC4XgkFQgpg9aX75CZWdhfux0rC4VJUtOt
ztK1a5mDHMpRjLSS0zgzGlzWE+7fLQs9DHbc7fm5jK/MKsD2ICL3kETKRMQ0
5WNWqenlQjnWZOLsuMLsmHHC1Rj6YUQfOwWp9LqYI3OJD/cdyVtbowWP9DZ8
d2xcM/5Ty8q3v9owdL2pXT/MSY2hsRzf8jCnPkL3I2/YG3f5t9A2SYBa+31C
9svxx/FHin7QfI/VYtE9U7B43hmsrD0QtkfiBhC1fm4h5KDsAKjFZJQJ0ryH
qg8LOPwuljULL2uHiAs3bq/KttzxHsUaeM2IfdLizRWQMoAQYUkj4fBa5uxc
ejLZVvPhBBEebjXR8oLybttfiHjdzFSFMxyHTk47Ev83zgEuLZyFAb+Mdm7A
J6NsiFBZT1WS/AuI2ikS3clywtSm/5y//hIDd5cWmp7WWFaLeB1vaUxdVMu7
P4Q9uADaZqKPZNilTb5PFAG6SoJuClcHyTfknBDNEYEBNFCcPn+J6zgcTgy2
wnsIqs4m1ULVaIk2H/8jSC8AIcZfTOVHUT3wkyJD7DGXYshpc0QvUzQ7Hek1
4Nos/Xk4tbWZ6pjIqSrhP7WAhhAVEJKvJCodWTncOiVVZjhSrzaCldHg45/h
pDhPG8ohts+6i6PNyFL3siEQR/c9/h1zHdX5RGI1WoLvtgawId1ZsU6WJl0z
Y5zB3OnJPDWsZ1Q7P+Ctl8tX5t5r2f13DkrunpnSNTu0ZVdhbN0nmNS1Es4o
mJpy1sRzSag04ngT3AFobhDaEwFV/oPAsEfVAdCad0p+EUPIcCKMVQHWnGib
eMzUS4XBZg+nJ6BfmpJ7WLerYhdVoP4N0YGy9hBwxH/yNDyQjJTFIAyHW0Nq
WGJwaePz6W77g8djc3Q0ZF51IPqvLDpqiO4+R7vwFHMI8luNFgxOs0DOgI3q
BKChiDXu1CpAPmvhVxE8aM6aONvUvn4yb1rGEp8wsffvZygStQ2LnP/N2RKf
JrWFUeC0gJHOoWJZbmbX0cpXUoTlqUA0J92Oa8uF89OBpIgoO6aMwxcHAsm7
y+QSNVOTvi9p9QnEa4xbdpXCdZ9wIpqeL4pWl+GfmO09LDmq70JrcBsBOUkz
pQPoUjzXKQVBTDQqJD/vdtVcyYel08rAENzslNS47EEJHrsqfOVhHb6+rzrd
rKmvc6merMwHZAlX8Lt1iDJj3VYY6fyCUohdaqMuJx0iNN4wZTEaA8hHepns
djkNMA9rrVZfUIzGDTulegMH9DfyZU7V62ZxntB+wHepoyNhJ7BZ/qyXjhAY
I/eUMEoX8UudKYGxasj9Q2wLTN0SvwndPeNyUUKW9EahdjgcepEWXrcgL666
O/J8OePzHpwPrYa/cboRZq5/XOVph6H345WXoc601OXIs2XErGX1qPdgK9SB
4GnSEtAcrlZ/MGvJnKIBBKEwhRYA++xfI4OpbfldgziMj87SnJ+We3STnCDc
wnACgLTaXcWTPT6zIgwUKHfkN/M74yFfnSOvt4guEZuIIVY28+aCAiub99yT
S9tNqPtDzvWF9Y35uYlaoqAARy5e/Njsqpvv51hbrLJxFGCt8O/IwMlhD6Q5
uX8UTIZ0ANXzvd3BBMPCHzY+axUkW06HPNrhqHNh014d9srQkV6Rz+mxElva
QasUntthoRjvNjAnXlQrl/J0W2AyAnepfsFX8lymkM3yx1j2ltlVKC93yQea
bYDfkEIKYB+yH8/57maUiErXiZ8zdTQ+/fULp8OxGOB82FCRM2v6L2WykQDw
cyrHFI9ma1KIAwcxkrYG9cZR3AHPg2BKdyuBpoVME/Rz7d/cdN/7FEjg2IwK
ysXOS/vmeP3KBNOsNMtXORiPNSx2ZqPmvIvL4xCLnRjiX2jU4i816HQIjz0M
Kiept/j6IeWqsp1uYh4uzQZx7t1D6yGIak/d++ZKqozfZHe18RA5hJ+USZux
lBC55rnzRulZ+vE+XGAeC/pgPoj8OeDlKdG1xguCBMBAW8rbWSLLcL3CD2fq
i6ql/hdf5gQqlO7y5ga+AqUBLHrm9iuikM1g1hHtMHq/6NHBCW27Qi5dPVdh
/m6m4Rcyt2pcemhyZ4Y6yMx8L4vsiW8ZgsDwLki2p9Wp9pYKmt3Cz1QQeqMQ
q/8xTDVNUJcoWhpd/ujuWIwLMlTvUwhj5r7RnfrnSW3TvSkD4L0QTCtFxqIa
VIfyjiZO44LYTanuU8t5XsqhugeF70swHaKMf8fX29Fg0o+vvQlhau8GoMRp
FFVax7aV+tOliDQd1cVXjXgkYlnP/K6iQUrUNu/15DKd/7B6rGZiYrPHFLLQ
lh0JOEO7I7VL/9qqfhN6UX+A+aXGBJ/KWNEEKr/SgiplmzNhkEif0EHM7vCJ
9TwrSzlUlltMf4H7ETM6l80ZklVQAqc7fan4HEoEd77P9/NOv2SPNZYFLFIF
M1UmbQ8ijnQuTyenymoBV2X0F7VcDeB6xp5ey/9VpjCTLmNI+nArRNhnWZ0o
CzkO2dLTEzjbOA3YzIMvzIaqWEolnDq6Ghl2pcp8E+GCmDcPzMi6saa75KeM
5HrzZS1IutKb1ZA1bxfNdOoMTTEKkB6fbW/QsHeLSOIUIzJ/T0YroNJLljsq
MmN05g0yNSCrdICYgXLn8gCFocLFz+WE9Ussd2KgZe4+YE77kK1TckEoCm6U
IBpFCvxS3yEY7Z6IaIO9xiGmA74aNe4zbdAHHtzKopxJNQVVWQWP5ttK+MXh
VSgztjp9EtxLNa22BcK314wbfuxCe4tV5kppEZSO8jnzzk10w1KX9zDRdTfd
hnk2ea7JV5gZh1tVve9aSQjUyidchq0podBhuehoOA6QpyXs9eYgSptSo5Dd
tmDn8ISylhC/ib2IXhDn+7djZt538ElPAc7oEsqfPVm9IOqTDdPXdztszyG5
xm9bjdJhjQen6dZw+wnn4muh6ZAcbbKWS3IwWfqdMPV21PmFGOlsiFLoPCTG
pbIPG+0cYTLcqfamnaTvGFhQfparn9UJKWPWghq6G95B2R4Q8aPpwbWKPoFQ
YCHE166zIyEC7sgZwQp6zEEQogJAuaavJ/4w6XjqjXH2rgussvTBIYZZ0mFl
GkUMzDydPKm7Zsd8eFWQyYtHVhgjZft7wyHPG7BrRthQhAThqMCEKw9yGZtm
Hp8ZX3ZkZQqFxU/ktXKsF61A7uwpOMNT1Jl5fYVbDX0hJLDLwhRSEnWsold3
8b/Qn9q2CE03/QziC16H9WGGFr40ftZ/soSh6Fbgjf3+wIedYD6iqrVoAoKj
LA+/SyL3EqD/JvpV/tzfhtOQUJ2Jyz6mxA+qwl8c1SNBY6Hjzkj/h3S2WhD/
N1m0/H8NcFvlWjZL9lWfggqZj/zocKnQ6n+CwvWd/+bU+D+w5F+QkyskGLuT
OIdFbpyYeAhQf6RVzJCSaqYeS6cNGwLkNzmSy9LE3Ihj5IgWGOXHmRP+2HOF
veeaf5LZ6mytRMV7KfoOQPx4Gd11+JuUJdetIsZerwNj+V7Jqu/gkruDpNaU
cDGebs0luEKrsu2tgsBPH2swr5BReus/zuSwygz7beoAcyRKK21uKy01D4Lp
QwVATQPE1x9jI11vOeaFPOTWCRa1LHK+yeaI54uypfOo05iY6sYS6EFnC0yG
PI4t0bFzGlQ9yLbxPJdeDEPVrXrF9JF1dfby24KbmHVjPfzbYHw1+Xsg8T6D
ugi2uVcX+WpDeat5M39qlnpi+FLhR1o7ZK1VvxBV4o6GwDPnmUgusLfFTAj6
XNtBqEFuGsd34jmVXiru330Uhke6YTKnOAkgnBDsBapXtnHQuXR6aYLdji4k
scnccuLO2asqCX9sLzr/HZIh8nEpBTRgQPHD3YObyjHYjZUaQDZLGxKhYbHD
YQfivs78zS6rEsqZvyEjIHnuBu5kLlUrdhl8GTPQ1kwYv7peFL6xMKF8ymHm
q0vNpL39V1UyKzS2O8V3ZDF1rsSwmvijLvs8gYp9noUyMCFlhSGN5QdVHW04
cPKyXTtsl6yNlG6V43Ti5hASJZDc48zPWZ8mdoUapkoV/uPiQpa/DyMAzgKp
Q416tAMkmvpGcy/hN/itENct8/tU/wW2t8UD6mFzhLJY8FDlFRIuoKVmkIJ4
wAcpUad3XN+NC6TxaztBhKljq3ijoImshKyQTlCdO1jJkCMMofUpdbRf1h0K
KXITpB9EfP4KPP7l0z/uRVCe0hmKXi7kWY3hklWLdMI1hKpHUGoLJQ7Dbbwd
cGQOuMIs57PYtmSIlAhhQSLk/p8nMT4Ay+wg2RSsQvzWWS+wPLuz7EDwhkGE
6m1Pnlg/Q4hREfm4QphsuHRxjbbK2yW/7Iz/3EDwejSMf1EpZmPDWlPwwgGf
glOnSbSPwSzAJ1VR6rUPx2HgR3uCL3PMn1GTcAuV0VQF26rEzgLktqry1l/g
pUP4Bk2YEAogXrLv8K2csfQWNZRWz355nsKD8WlueJLd+SFof7S0XAJIZbIy
xuN2l6XfDE1lNOpQsUKW9ODxZOzIozvZ3eeeVFdoalpPkYqJnW/aEfdf2bTS
zrI5Ww2irT+OCkrJnnb4oV6jaYyLSZsagRBwJtNAQcA1YubiQREP8+evNhQb
yWLH0irCNKnorVO4fwui0zaBslh7Tmj7xUGR7p5kQlIjOveWbQgcPVrPrWgb
dD8NT8160+l06qFOnkXv+AT/8HqHmqZx8eeqOsfluKS/2A+j7l1xT7j83kTT
csnJeL1xTotmpM4DmDxZJv5UVHpr2jJSZPKJ5bR/HepPXwawH5Btxa2ATldS
6ZfP1rJYzpbTDuEjW3jrgShA8XZgxw+cWV/L/zz+RBoyLNUmV7eGq0GcEtll
0M/iqcbjOsJYjFHqVj3vMJ1bTSF/QYgL9h7vhvHBbEzUVTLi9HJ6agGvnVgG
rMuVSpFIceantvxHFvyaLMX6bZz01DmjeZnN/6xWx7dKSebanCwvsyZHKEtF
LKRJavSxI7RahKsA6s7wOiYT476+0NGs8zLe473fQdZfh84qP9hjnhIxQAlY
lNyt/hb9mbNcAz3VMnQfzRC9v8+hon0GymIE6ceivDrerXS+3fpKZuXIeElQ
do6lg+w6Lliq/1no0W7cc3ZrtBd+LmHkZ1dQ63KbOxsQ7O8RHkclGTJi66/A
rAfPWSTKcp9wD3++aoHjMNIwppF8plwOYH+fneOrFzgX+VRoE3zojjuE7BzU
2IytmtXFz3PNx0SKpbWu0DEl6qZy+mfCjS9SmiqpYZPkVrGdjQO6iSYp0dMd
C5t+pCvJPhSPgo6aPKf++4Cx48Mazp1VexE2EFwod5PukotOptqe5uvqodab
tSXVaX45s6Rr4cF3QyKHvw7pjCeDICy6iNL26TkvO3Km3xIpY3Hl3QH2uajx
0M6CjVzgpeBkihJL67wvP3rqnERi4NVn3nxX0oBBTzpbtGvBUM/8kZ65g2t3
S50Ue8MhSahocAC08vSLtteYz62ArPIQXtZbsE+XxtX5KwOmVe9jLYvX1dbw
wOZhK7qChBO8d/I1BXw+0RhbqXRROgEtdwXqCtnf/QsaMUeSOTjS3aGdIPyA
veoci8pfVxTDV/dbH/sJZWuf/+uL2cWMhow6zsEXpogk0ijBE415u1PBAzlN
iQY6pN/UtunQGn7AFZslkUIyozVOGWcP91wuxrl9HMb6ZhSN9Z/Lqs771IPM
lWmv6FpdJXp0YdI++r8NUCZe4UdKpKoeOjzjI2AmDNS+2iWEYdXMzA06Eg+C
kVIYtkVx8hxy2p+4S1BP5k1liXSfdC3be8vCZ3Ps962z3N0q91hgbn2K5QrN
g3s/sem7L7CvWzJGPM2+bYuLrOQIZYyYXVxG5tpKuNRLTLt1IbojGUj5EEO7
8XIiA6F5xs6pu+pvPluEXRuUJGeYebcXAz7owgZGWAhes/0vIzimGV0CXO8b
BWbcUyJsA29dhuna6c89rU91GlRoqjFoRjjKpYhYfcHWwCh6dp0nvvW8s5ue
HoceGD9vh5w3eZZxSTcrrirVPbEvSVh+HH2uqvP1XtfIDdGXPMH59ceiQ2L1
kPOP+60dM1Yi8u+ZLJD3nOaUpfJXKwLyL5pLJ9HpYsBrgL2RP9+kUhp4r7gN
g1RcNElLwV1oFTx1YOtTbkvZRaRt6iRLx4WZKPWhhgln8xRGOGqNQyqahWWT
mg7T/0JSt8EZEpehdgxBYRrnd8upzfbo+XGeT8dvbttihZFOQAZWoU0LplpB
PN3kQ/XKQDFg2lP92zN19/s9cNL/i0sqvXOHJJgxLvo37Gm3XvcynbShHrMz
W59qf9nFa82667afszxdCq6FROO5Q66NyZpV/KvRBG9jck3L0j0CA2lAINAy
r660Oa8NgyIGYqpSJkolcjrwEJGKnChlWzc8t7Wn2+BT/PXs8qnb5g8KH8S3
kSOPLX97PXOhLE9v+XIiahgVqfjLmq84vXj69sRKfLefZrOc6lU7LVIH4QGw
1fFF+CbhcGiDVdWFfib5f3nc5ixhQSQI2EtT0wAyVgq6zioKy3D7tURMWX62
ojx3hUJ/2YVU7hwzMDQdkF4yQlSb+FQkclf5MHvZSsmB/mLUnmrWUgcSf9Lw
uMRcwHhgvfHw0JNNqL+UrmrMV6YjXOBXI798SwYc8UuD3tb5VrGkQIRHtMvn
zUMSCe40FX+BZvvGvB27CUceZqWynXIuKxPeKsAbeeDTAXd+yXoE7f3H/fBg
txzNPLVlKC5o3siU5cEQpbAHd6XLXVfbnXNnQEA9RVS5S26v+OGDzF3lLIR7
+tQ5rUJjOrbx6YzGRIowO3yeDouKNMePoPxsQaJ5CRtR4oaDHgfmXlnoXbvo
6n3K1Cj+bE2KQQiZvNRkQwTYaMJyhy3pzhs4gSeaWw6GbcZTCs5rR8I9fIvq
NFdNeGm6tfwD2PaBh0e21dJ7VhjsyaXA3Ev39ssyLKstWAln3ykQiGP6/evF
sImh3oRFVV8t+asGMJ+FjSSVqQrjT1AvG+2USqdcY+YRE53jUOsdfEljOfWL
MxVIZELvHp5W9p8gpNWTwr3gJmc44wRX104IYjFv2cyU1tHwngPbfF5m58bU
qIcG+QEmn0S5SHM/CHiVD+oz1SEW5Rw9epadLa1VUDmHPHU1dIiuBF657p0P
519cvmpFF/ACxYKd4Qx1YO0tZPtGBm5G0fo56VT6cusnAFCXyN+rXU35W9kt
rfk+42eCJdAfxakmZqA5dPihQ2H7PWoBJBHVr1m76eyNggUf9sI/zlv6JQmM
piAM95aA3mu6QNnPGkXM4bJvigXVTudef7RkbsdwnnXcTUkPrKWKItWWzZi0
Svh4ivrni+ifVLVLp/E1Rl5GHv1rR8SWbTFfKdP6khE3NKWMxUX8G0dR0d1M
4G9N727cSkzTyFq92wX9Ps3SOgC2F7WXDHdPcTlo5E1n4drf6k/1kkv/NI/1
/rj9fHb0VGxLTm6Uvdpd6pAWk9WMKZKVAptSHte95X/rPNCO5j1B2SLbUD7h
msxOy65rVfQXMc4gMfANaBPCqHD8JbBH5JPhd9EiJyevXu3hS3ECl6DPlnlR
Kt7RzdvVfOji9921b3J+I9UT8WMals+7Bm54umd9nDAFtl2XUCFVygmEykBR
zDMTshgyK3R4A60lOMEQPQY80XkofqScEfKIJ7F9pzNst2D0+UsaYvZF13CX
pzaeiF49z+pv8sz+cpUo4x6RwM0c8z/btsWSDvUlywVUeqFJKZ5QpPMEayvp
uiT+frNeDb1W2A2WXKOtqAVO82ANUbKH5iMpLo1XEeAWUyJ430ceS+ks2wX9
lY3qAFatM3zz3WqrNXoCFC5g+sBQ4G9Rn0771K1J2vPNkIGnea6T02Hm+rRR
o4GF/aotC5e9WdIB6jvmwBjYtHlhr9oWKlMCHkJVNJmXzZasNLAX4m/SBPT2
oqbee9WOTGys8XjGlmndJL20mYYLXEU1PjPfb/Hk7zfwZE+VSuwc5PUYJE9+
iV+ig05MqT/JTXGjBkI0XsTUEXkc9tPiHg+LSffBRR70KSxsdRAWXRznd1DG
LBm0tQzNu5l69DeM0jdURovOKUoBzpDRIUNHJP4MqvS7azyFaV77lOZUHOek
sPe2dGlsf7jfUfiZAKWxSPI3tTQv2ZLqOVqhNbeoR+EYNYAl2m3n96IIMQzq
zqUiuOQgVY6P6WuQYjSEZBFuBX/eHM5g0cjFMlAWnRceuqItgfd6/WtrL0as
Qvv5eKQp/OUrq7Tb2pKSNXMN86XeG0iUd0KwrrzunrXufxVBaldyHWlCrz3D
Ncocixp8+j9sZRKNuXxtqLdPzqMnTjPj/dCqrtUu11YuH7Lb3EqH0R528FYW
jJZO75/6rEGAkn+tyYd8FVnevasDMsZ2ZSjTSjuq6kprttaSQA3wbM96JH6h
HrafOF+6D9px5+9IUIrLA5z7LfVA9YbmW/3e1E6VLzpRlHKX95pItzpXfC7k
zsLrRA29Pfw41LleGlWlC/UTjsvJrbixcdTtKHmxBQJNXhYlJYgWviT5lF6q
hdds4vAYBK4WdWfzaXMJAi9b4Vof1RXNxo1BNI7luPllJ6z8MvYcIR6hOWZk
iQcEMHU7rPdA0pK1i9eGRcRbAqrFjljs7IfWI5ti1hBPK7XXrX71qHFI8J57
u3AEg6Z+iTMDnGfflzCy9GEYhzSZIgS+F5+L2eoEO/hNHVK2QaNp/kJftlEA
bpkJC9lM2m53ExSiioWIULoxqGtLJyCUodhLNua3YyDB/6ONn1HP/xaxJeUU
z976t5X2hwqP9eE1eLoHc2H5BMeBgl/5wqGTHINL5wQ2ypshvUN+Nu619cKw
BBaZYkm4AVrj/DtULRZmbmSbewhw8FMUrI5UngPn8ZKFJD9tyoEZndnMgjRp
Mf2qmOaj7D8JEA7XWAp2OgBw95PAaCQ3rI/2D1Z7fQs31YuCOdiZtonnRrVn
6IcldHeZV1TAdPsoT5mMf/rPYnpSwxXPuLGQ8l84UaoiuZKL47XRY0aK38G0
qceogPWGdIwZIAHinpcGT0gi6lRtF4aCF0sd8RbD/7Qassw6DymX+kzT7Diz
3EWzSmyff8XRiAsag2VM0gR5AQQs8sz0NwUqMPeFsw/NzS68j//i+6lWNdFk
9ENo9vTsYc2tFykeW709NeTd3M62mBvc8vdyeIQU+SgOElOemr2mMvRaG2pB
LGuk9oIi0kDBURf2UsZcbk7Q+HrC+U9buBnGRtHySUFtb1gQfLPvUGzO+mYr
Toac+3rFjPEIy5ugG8zd62uA3MtEla1XioH4N4bZKzQRaUB7iKp0d5ylJyQx
yX0txLX0o+PwK746SfOLeV0r8F92jDCSx3CnrAgt65klsS1PHrSVGqvgHVWb
hAT+LduLXPUg8gKQtdqIiKlm07asczKaXGM0dlud876DpwJHEfRGmRKZmCrp
sd7lRVRso85sR2/oJcMzIfbLE7CnJQSFkzfmQ1cNYiFdwYquomMAdNJxUq59
5tO+Itd+oQp55cTeD0hfpa57IhjkQRMfaYUdUCLAjofgEPkMEc+3vCfKfPJu
8Id8op2zXfSlULE0uyCU0VDm7V7P89J43smbi6lCqml49QskpIw0cMklnKtE
sx5gfL5pgKQ/TP1YSPzjiUFIXekebZ8ZTCBEJyglO8HHxSH+42T+9+s1KWNx
cWZSkSCw02ozi9OCPKurRQpuSwm+IpIymIOtMLGexcib9tNDgWU0QB7BWYMH
7b06Bdl/9tVAC52cEZeCovk/rXUVcbAOUaHO2HUeV/izyGXI2Ma4sPEHE80Q
gaEEoZuB+cgR+6Og2w9CGOg5LXIqaL2lP/uxMpP+rMK9cSIEVUXIW8gzLgYq
Eplsh/3FxQrFOPM3ow7LBYyUvSoaXTJrKd+TZFzo35nn0jwrvO4lv6z3r8M0
LfZcoxIQfh1+MdfixvyM9MLUjSpwTIZ9WMhr6dH1lSPT+mbgSzPwjkTtYZUD
GKbB/SuF7wVQbV2lItlaztDvZxyZNtIhf+TGtuuFdTN63P7Bkvvv023XyFsJ
gp1o36tYAErw6KevKvhmFyzM+50LSuj6iNNCmZRLtC0wzS3FHY/xP1XcKkbz
/epNvEjneAYUWIkf61xrNRytN2VQ6ajghhpnCUSP75mIlXI2xgrlIxdjehhR
4FNIyHftxNMVRXfLZejAwl2O7rp2L6w4LFzDsXWmxcfem/uxY+YnGYcZJGcS
cY6lVbMiPziXWu9st1THk5P/z+/sxi3v2OXzZ5Ur1lC9sklqo5sGZHBkK/3L
ECm1IAb50xWHxs9CJt40pDKxf6cL9QMXon34ATmtbdwtNGyy8+WqMg4kz9Ot
qfCvnTj5EU/wmxTDl0KOI4NpKxzesZVXlC1WZefxLOicsk9ncasm7Ln0HlED
3TuEU2QGCJxnRbDeFyuQkNsF4mmZTXhgmwEWOBE9MT6ojxb5M4y83Aj6Trsq
xlwVDtYxBKyJWiVItxKUMHZj3UCxYvl7eK7C7lATc3Li8AYzzzxgebf/on6z
BNVV6TS35cpO/RYE+boMidUcvKh3Ea3DidhT9/ToHkOu39YhSM9TOScqehvp
1KjjylY9DLk44bj1EisYRr2J1NZRwdzgQlDo968PgCAlsY8n8N4/5rtsLtf0
sm6W88/bXddoP2IGv8H9sOAMylsq5e9HshDhBGVynrxDRWhTXEAYtY7VNyCI
f1Wai++P/XnIkmAE1W2KM+M0BfxhVZMnMl+Gl97/qVb87F9Cth0CU2J1Cc91
GJ+xDiKwA9fEVJQzAtanqauk+Gnkn/xkPqs43/24tEzl+nZogCL2EhVaZ9ON
2K9W/1TmCpx89pc9Yvbn8et9ASBi66Anp/DtAAVlAr3OmaIMDJt8ex+8mx+z
STa0gxeIP/ABgKCB/4XYWks0uZuW6p+b8udMgs13wC+X5NyYmu6/TZw8AqI3
YDRo3wpWGeT9sD4nsOQ0vnX2qEPCtupYmRdKpIPjRR6lU9UvutLA/3PLa5dn
pIcxWIzDZBJsFP4Mi2SLB18gaGHWfyusu8HVqKa4vFSGIqu/oagH79xH2IPD
RF9McYhlWPq8AgAZR8dZ5HwjJu2SkQ0y4+C49GrQdfW1IVtoh3hzmDGC2Fq6
y3T9WEsqyNSwOi++mpbCdGH1Np4T+rBchw4TPU+OxitVnE4LXKSpC3hrqJQb
P34Xj5ZNKGG8R9+FXuPPKuM6Yzcwgtup3jTCf6jUNG4PpRe+vcIP1/Zx2IZg
LWXEU7KioIvyR2qCLseEz60TDNe3Cevgv6FRHV+ar1wPZlh5i8XMslzqFBlt
LeXT16Wyq3G6E5keIZ0LMoLmBKHEkgEnSl0w+Cxvx5rx06f7/znGo36AN3AN
O36c+ZdM3hTz3qTziG/ixlg9wdWTe/g8swqGdz543s2q51ZfnAke2p9/mFaU
zc/00asvdR6pCVIVS6n7vdyC0g+ZaY6DC3b1zmgniQ0PqREwmCrq6Fc6B/Te
dJcesMytzDX45/6GmF7N8mhbbXPsN1X+EUbDHOwAe1Dje/ABuh75Wa5HI+Y4
XeKCxq+EzPO8qD2RmgFZBLPiLX3DXo+5Hvfb4vIvr15LK31JB1sLWuyc6B+4
snirw3BqEt9s1/MeFWddP2HKA/0/qH1nSeqZRh/C6dkWypvMeVknN4WeuKIZ
mPNNvxJH3tujSH7msQL7J3/G+EdCBRtLPGw6cND1whoaK7ZWOm8auxDkL0/f
omQ52hdQMR409flMgdjIWiHIOlPtt4zJBsyny1bdcF6yrUpHjZcpRNKPUJE9
Dtgpc2R1kNCn4UX+KLPopcK6F0Nhuw7jcXhaCg9+EMu5w0RyEk5TGI6WvkQv
WyjzjwWlIo5UkPznCL13qVnhj4f+41DtzLybUWXePfqnbDRNjB7LCGM96YH7
DKRW39LMwJWQCWQ3wxUXBPCmtmEPE79tPWmVxah1hR6WvY9ZRUhjsfXY4lX3
79hyDoJNrZHUN9Q4y4ZvNX0MFazhXUzucGEx04/Uc8zy+RJiHUNiHFwuNUnc
rWtVvxrPu8g9aUa3JeupYCqZgS0s3rbxxD0ZtgkBnh+/p4lmb7XybidfIRrZ
YcxNUQC3Cu26q2a3gBmzfyFAevNl+d2nCWZb7O0MeFaY/pwdC0mvusLm4Szh
WIqgp3m+pHIr4kfbz5ZO3Lfqir1FMI8aGxG6cvaa4vACXdV3s6u+N1oEnFiO
Q916Co1EWlHR4Vp84HPRkDW1/oQWta7aCOlKFkDpr9mKVQRnAPcDjl8xjmXG
a9Q9Z0e4lPXh8U2Fv2tHcxmz/COMe/tgJutufGNWYztqgq7LJaHeodAqcSSQ
TX/HA7xTCsZ6ulQwy3FXfXgbans1ZTXSCeutO0NNXZsBIgDlCDVuKV6P48mY
HxA8dUQ8w1rm9zT1GoMA4nsWVKsQoxuCsM4RVjIG4VNCZJwYFOTVDA4xQA+j
uGXYArNm9nSCNCEHQ0wBOX/VFbuQFeLIBvzg34uEPp5jz/9bYyHj7xl7ge/M
xRga85exqxUBzOgHlBsEYEyavDcKn5A0D/Mm++nmLgmLzJDAVvi3/NYRhafF
H5YsUTJDVSHFGuieuUqZ3WQ40LOD7lnmCgMWyPBEuxRVaJ9oLJJLmyRFknmV
Jz8HDeVkZ+4mvJ3fzFymrDXJnp4WsuaAPWkZ728/xeYrt3/kRSH1flSiQycy
ePOBt6dEQjB2Nw82ACxH9FWJHAIiRs1zKEkmDV2JabzGQB4PrTW/lQpmrHyi
72sNIcpF8BZ6h34jXzEvKCxgIHur7qyflyJ70c9eKDX+0M5OW2EcQDR74Rs2
5zniJPMVJpT2FFuevJNpLnNGgNsRQqf1QlhZRSNqZA+CfHzrM2/Ij6jCsu1v
IuE2z6PwiKeIJfUcio6/t2tIGIdTeQF8BfwC2fnWM5K8XD4faxgQkjTWlQR3
DL+oRVGTIy6CrTk4VUnTh0tFDYtO2rLJ/7jci5Hf9ybykL+1FPaJxOgrusA2
w9LX+XGJasVLLn0U9TjSjvjaYo1h6+qy9XjsHbcvMmcaEA33IvmFgj4va4Tc
BkUxmCwCJQozv80+n/0CWa4i0k5eS3bY4SPuSrBp7vbSurzLNi/5CFbzmVb9
APmNsUPYa5WoKr4REI1cm5cTgexW8a4XSAd/fLOdolYnqCjTthHnBzqwUlzA
Df8l991V34gawDzz7RsZiFaT/QS4AS8P3q7r8cgV6WeC5n+OSRSPZI6w3VJ4
nZAbZSiYeZ73TziIma74Xys0aIMWcIZd/zvL9f4nngJD6N2b3NF8AI+EH33p
L5EUzomXDLAyTc41hoEcD1A6HqBI0NA2tNSYZ+0fSs+nrnCJ1aUGLIttMzEz
MsypmiHBE735jdxZxsSVuf0TWVn74jVA12qoqIAlXoGx2KP/LnWJaRYHbIA6
QnAO71mqypgdQgtjkw34KbfYn+HsqFtwjzaxRFu3Dso0SPHXrOOl0eVWtTlj
6dvLZkC48u6HWHZO2AFU82jzXs9fPpWx4I77lklX3aSXzvzG4FctM7yCI0vH
vPhgX831wvHJd+QuvZ4JJzFWRQ8ZDtiDmOJNhjsDajzU+fm0ojoixpTnfsM/
dEh6JAUCA4mGUOmZo+GCEvNlCVprepgR0ypz9wmMApiw83QxdNZpG0KWdAHp
pe16ttQyyCIKYT4if5RduKzZVwPq2BVsJjSbnmj4v1tnGgaPzDVTn/cis+Nf
NH7TLZtMeJ84GY0lmo/eJ7YbtJfJNNPMmEB1VRav6FmD4bUrICOXNnVQkkfV
Q+UXjRlvVe32XvLZ+E3KFjVekpDAO6unJQ2WtY/+lC+/r7KacMEZxem1OA+R
0yMP+28yO3WcFgzSm5Cu51AKTfQu/g01R1vMOyHZ2AHZIn2YmJvnDDVm0B2a
NzV2ndU+4EjyHIAcE2xM5eviDj0Crk4pG5EFw3bRR5FITaRbTZJb5/rda4kK
QSSm2tl7RDg9aRc/gnDHvxudMesxzjXtxun28w7qkUiVoeSRl+Fzg3LKPxqu
agBZLgVMKv2K6ZUw2eSX+ztnj7Wok7BA6g1rLnJC03Szgn1q3Ps37q/EL/7L
oO4pCd4XlhwRjnZ+rdCMfVA4wlcokVG58kgJDtSCxaa97JxyLZg36CXHcJeJ
Z/TP+ZVDW+OkhpiUMqACsA5teB3EPSYJnIjWilooXemsuxrabraa955bYTRf
gsp/i0EadGWo2yDUfItmCH+Zri2CJS9bJvpkb56qyeGk+vKdTrGR3C67LyWq
WIsgk6Y27a+HxAaQmHo3CrsnRMWT18H2YS/8kf6hj+u6U335v2neJjFXK132
vEB6Xcw9pKKwKGniEnuAgVBA7iHDj8FgoPczXx3a4o4xvc3iEnG2xpXoVnXV
TYW2+bO5/eSbWMzmpezrz7+bGgFIodYUldViGAArEpK6HnJSpqCdWqSNJa1r
rG2XUu9jz2aAFhQxuurDsXpifR29AuDnCq8gJ5vXft57FkBtLBP1oInbBvgl
dAVAOTr4yIShK+bt/QDk/kR8AcdV3OSXLgPqch9aqLgrksVQ7oy12HZC9rW7
al7Dvg65VNU7q45Yp62By3KoGn/zhyburf1ecz2ureXq9cbuynGf90PaiMRl
HW3PDER7SZcWXdA65LXIpaFfK04/QixNc9QEs7dCXVVezyHNQtVKdak6jlGs
pHtTVM/JJQw2+WaBCMkTFqvgR3JQbw1PTV7qoZqxEyH8eeCVmby+7DKI1YM6
ayxhMRpNiYkr4kOqeBrnsoh64G5IlysZgG63O+qmwElmoP5l61cZM1yT5Soc
fR4uHOfreHpJilJe5MkGuUUd2neD8pW4aaIqH4cA+1KpCILB4tNFCek/oRwY
nGxSYVfOrcc3YflSEwJX/JsdJBsPRFg3KCIVYiRJajZCZ+2eT6t1nO7zqpzf
W0IA6iCneAfLAa02BtSC4Hs38hasU7tdm8GOIIORUrWZSdHjnp6iMLZoy0hG
xZB27B3PXLhmufrOkFHtBbvqbh1eMbWG9Xaa0cyn3NUUC4ltFUy5JjcjSY2y
3DYsrLcdh4Zc4KrSBYL5NLC1Y0/UnMd9tdPrkqycJeznGgatTiXpGAgo367w
k/LcaUBTCnQc41HH2ZZbCptcdHARhAJU/zyadimLr27IS+/wUZX/HLySNhV9
vXfmdXMSbBXfetGHUG+hfkHyLLzzoKO4RKbp7bU/tFARBiSRrRqvGwM85UhA
6Ne5d4eEo5PIXISqzMC0pC41ycYGYiDs6ZDWh+a8kVpJ+dEuvM/QDA9+Mnd3
Fxo3JmhXkZtsayFrsxMZ95hXit7lk2m8bHbrpXc+hjjHnxbq9lxTyRh4mg/g
oGo9PO/iF6MvDhkbTml0lODhg5aG2CghDRVUP2GWn8nVCU4HJ10YjVwSPssE
U3RWrslUPhh2YLxujcz+Su2novTibpI2Y7gFpKHzIi8OjRYjTASDFDXh3VB6
5nWZcXl5jldXxcPwVbS+MAAa31PZWg9rdiTDOA7aIo0jAava0gLlA6YJ0EKP
8urAM/UdhSx5qXxldyLkmEAbjVHSzJKwTVgTvytFO5G20ujKaodIpHlCaIsv
d4osxHc/u2oFHYOB0tkG0A9xCOdLhmDRTHsqoak2taMKT4UKnPVd+ZzwQifc
XozzNb4icxXUPrQqymp8Cqi8NPHQOHGGhnoQAQ4m2jfTDoDlvETxDBh+Ghdk
UBBh7fDmMw6/0hB6ux1djxbZX+f2X1tSidoyp8xlg1J4aXkqJX6dIpew3ztn
oTRSpEvweimwkfWtY3ysnPDmnWykkgVWYw68zOwQOrtVV/LwRn7LYHptlr7o
+JymtQAxGmWAJv3VkuaMO89yeDdkuKKh7Cd7iqSt4PihB+0Hkmcn/f45CoZw
7FU0AT8CgYbm6RnGSpTKPbga5ttuvAWNU8sTi4R7iThF9ZidKhBt+AEY+Xb2
H8qtax5haIMJfrQ1o7sd0Zn8YXcqf/gR69/bpfkRQcoeOHZIb09Ow4kFDYZZ
ffNbMF3Us2LQ4WJKwmoUEv9BhteyGXobITmG0L3AHltd4XQqZ9EvmXjTQ3fj
gVjIst3u1MwSmmGlAHKqMomtzdbYyRUD1nCr36yFI2eSIIj/YkT1kaAGJLUm
LM8dki0WbuBejyh+WLVvcjBDHWSRUI9I8yRrJIy0KZcSrvXJ328lNjaMPH7I
GR8PQi9yaypQSSogjcoKW5xmSEAQOJ0zLi0g9PFA6EaJ11kFZUPdT8pk2cVf
ObzCha3kns/LjzDeBTGApWu9+8kIfBfObuLWJxpZJhKCN+uqip5V1dgEP2Aw
4HwBm8xs5IYktNtvVMv7oV3M4KOqmUYeO6Sl7TdgLOoH8g1zKFZcSJQKfDfQ
IChXzRX72aJQjsMSEEu+50aukLOUeFgH7nOB5Fj1Wf80sTtaMLPr67ZKjmBJ
i83vfUYNLMtZaSf4LIaEy3K2Pm1jZ1uV42JYUk9mvaNZA3ZmtOsO4rsXwTkp
eBzfUBI/CN0FLZq7ifROlKoMU3LpyMGs84jc33Xjn1x3LFrufwqM/W4ADFzo
WOpPsVQozqhmPuVnemkAzTsmpyC8//Ea6fQfSF1HHq+JsA6dd7g8Ju6CLYIw
eH0IutkWL5bPG4tTlBI61dxR5N40545JKLCvday+WSj/92ZLoTMtg7pnMA9L
U24aFFy8MCA8paW3a1AT0UR7s9+6645ClhGYYVLMrGQyiE0EtoIjwTZfj2lg
erg8fpwS0jlgrCwsbe9+usde5JMdkv9GFEGRdGYc5lOHfKDJUS8qPFM8McAf
jlQGQtdEeKMCc7XLDLg3oUQIPXXFhbaFcec3nOnzuOeicFceBc64BQP6zQ3+
vnRYnUFTRh77F/h+sskTvTM154InGFui6dJAUEjS5B88IVqgC6Uo3Cwmqf36
4Ftd1VEwd7KO7ifkYm3aycVIGkXVf+agviA383sGbeHk/7dxbZ5SkJbWAD8s
xnxW3YaKXMI/ndX052YqbjcnylchbZGCWKG2uXIzMBD+iVMfcIAZnzFlQAAk
6koQVunHfIuRkQimyAA3OXCrT6ulSiVSnjEScfrtiVYYoE+pFrhE69sPZawV
z5bbVL0cs+E5qZgg12cvydvNskB83uR9sStQVYiZFcnwEy1M9McupaBaoyin
fFfE2rysFlX2JNVHI2r30ll8Uklvcy2ZJuViP7s6zC4Uh9NejzQVZywFjxHu
9vCZXhpuom5L1G0LEkPH9WBhvCVpvsFf+9n1OuPAFdrDSf3w/s4ruvPua2tk
yR+xjbnod4GwG50yWNo8IdT2nQuHPw1A8hzjX8PQxqpeyIPNxd/+kOw+zn16
LvRMiANmiHNtJMga+09PgBw+xqiL5OroLQ+VKKHohxFzpuaGG52Y6d4y711i
Tf5JadJvuHxtm2pAwNgnxTcZ70rUmVr+cfPzAUghqnpkeEXrbmBOeU7QBSxk
0Ku3bU5qtymkBOwT7VV8Wqn0oFCkBKT3LmDYLvNXIxvkSwuMZyP1rJNHICF+
yYtWCR+mo7bd7IgV9QuBPGgNr+lVe8rblAoDSifADc1oopyt7Bh/0ABUIqHX
NP7ebgfp1B03X8gCjCQ7FBRC7LaAuS23HwXhNT+rBrQuJH2qSoevZEsjRfKm
ySUHQkRNxwnHI+TpWtELrAzOf+iaZuISjyZkM9Krd5L4EM2He8Ac8KvvfOAm
SW3t5bddHRtSXhXSx86wkk5ZX8XA/Ez6T81QBjnHI4p0drsrGl5AKzWf8/jA
HHCIHLTN1lYSlIMzyrObe3wx6JzE7BogGeFkSHASgE9dAPHpadD18MDOEat0
aSk7CHVj9W51/qivAC2L1WFICAu5WOuOMz1IxpBEusH9u8O2F6qVKIZ6xds0
NS/TDbxGnd3W6mg4RcjGGbuCUu9ocdzKavh2/c5daJ1+F3mTKTYLzqm6S9vc
L7MKTfZw74ZiXoDgMWqipVthHEYb/rZLEVA61QttohmRGCAeeG9K2pzJ6lKq
SQ6ZOtanLL5i/4tdGMK1f1ltletzi1HgL9emy7IQl4mLfLqfQWhD+VmV6eWr
5gK3gCb7yEfh6JjnS+AJAMOGNYbpqp+MEMcLJ/6hx/22oNzB8BkZdlUOFoDL
9aOD7LUeoIii5of6FyUigyq8vv96i9fcknF/L3LNREpdbiXxFtN1kioyIwxD
NFJfKhNB4XA9zcpY+HQ28H3P7htUpneQt9t8GlHmZRHZwPwiEO1HOa1KVZOu
CTCZB0UcCzvmSJI1RUT7V8bMnqHXebGPaa9qeb6hVeFx5YOEl8N7N4wkPUcI
Zg4vDjVsyh9yLsj+DVErpoVq6UFms0RpNLAKM+NxodGSzFZkvcZEfNBFTn9u
LaCDTE/2njn1Ts3usCTiDg5/rgrf8P5UK6jO3k82fIizuuePFABvnpuGOmYT
NgWdBnWi1RW6JBNWqJ3H01nl/XDIEH7BsrInifSjzZ/8zvvY3Uj983KFPwAv
zNoWAxOGHQaqCw6/Cec51hdfthYnHZ+6lLOVCGY0c5h694rAdXrhr0PYUiEs
4lLcQhdZNjizRCRLkdKVxSw5XbF2TFaZEET/drMXidXN/ypVPUWbQvjHnpPF
o2snqAgdCtd7ZTPcP89IMBzK7W9tt5NG+K76xHCFcwzBfxChL7ugIoXVrrRT
25eDHnpNQpLFhdfIDHR7JLNeX1QgYTvT+aMveqZkrdw3MVX9DeSCit7qMhuF
iEFEP2QaxKwbzA+Z6h6YM0ad1CY6Q0X8Tt6dqiBT5tEK4Q6MlrC8v75xfR3y
RprADFHYo/xsYc5mfWg6ax/ecSha5UzHvPS26pkplw6GrWAqUsipx0D9RZcT
gYjP8TXQHNE8oDkU2jBeLLS6zOhP5+gPXJlFnJn1rav/NopBi0oSMNQ7dX2k
kX1jiH6XPAJi9GpwA7bmiINwpffkqI2VKyRhI+112VZ1eiLypi/3wqZyYYBh
YpuOQdjYDCmvqvUACFOVMxeIjioTaYOojCiqvUqiZpc/TyYSAgv8wcyjjc0x
uys9DEWDehoaYAQIbsPyoNaj24rtl9xSv7UkQ7Bo6UB8i3erkH+YdRxDv3VQ
ooi2vmnMA6hk6Qq+F7eWWgMt3noZT+hXCgoRgwqEHD1H97E15K95GziCkY28
DhDmWlt1OuWeyObDFaGl6EcqrkW77qYMaBr9+DrkISKZQGOkCEB5qQ3cQZYB
LMec4GTriIGwOrfpp/CHJcYIkAQmE+djDcXw1MRNXSIz/9sIJUIWnatDGF4g
n763XyTfTZ179wCqac+8LsECaYw8TJw1Byuy3pIdTF0XxuiInmSbok2G5loQ
Rd76sYwVgLP+vaIoNELm465kHOHgGlQay3SldNZ1CsZ3VFu0aFTYyxqAWEVL
34ow90of9fGfTnSOQZhBehGHF5qRZ1RzdfTMCQuZKPhMgjN1mYlCbzz+pCyR
/OQvld9gBaHHwbRHDxkVYAU20KnPzfaIoS2jLFhiwMX3UDeS0oq0bLdEUzcj
CDow0ej87lDpHtAOA8hcT7y8bc17sMRwKZ8lU7M/Dy+tCsRBPLQSoVotJSK6
JwWrV4QsofeEJWEUG/3wQEpR+0XE1yfbz2Pr/YTv1HkXtPow/9gfA0moPoQ/
uCTd4mtAoYDOaTg+Dvzs1fFLuDyKPM71pi5+wwhnXyXFwUb9sJ5j26BreSwE
PHxS2vWWXw6P2AowTVRi7ATVuXQJAabMbQ0IZLccoj3MFNOEch5srONXlyGr
MLpV0LuOLz1yNUQUy3MPb/qm9gt1CPx/Bqe0DnJaddmOZQ58ZyblOAKcMLMJ
kykx21wFSC4NahaYrBj5uuT8vuth6PFWBlzMyZFnvtNsG8++TyVgN1F6nyv8
FcEgjQrxRhA0aPxL2ERHesPV8MweNsKGUtx+9PtIbq+eimb0QSLrgiNZqDby
KmP3l4GlZHTlH9NCJQpYn5vQmSQ58SmbbtK+GdUdW52XOI1vcir+zxj09hk4
7F/O5T0Xm2i4pHQv2b1E0jwCUT3CZaZPstknZyO5SR9fmlMRjOOK3yjau+D8
Gm/AWqea6PPB32hZHw+i3vpdAkf6Ic0XVFGDE/yTusAn15Yop8Sn/i/7bM4Q
rc4HcLfvh+H1IRag0oKM3Z0SGY6B1OAFJpaG5sTIC4TV65KEd+vrQpK0/UB9
02DSz/H4O9zZGiyvlYftQ6dnNtTqKGT2rfqft2w2eQh+m9fc7DPFtmSEMaIT
zvlC0JbE7LUwDwJWuIhlIK1wWgrjKCJESgfjaWKKGzgewjOgxIQFOu1Wk7Gf
FPBsO2to/o51477Mp9mcSSyBMaTR+GJKZ/BRfg07YXW81j9LUhNDUjfRBBDZ
Z3sFZEt98s3PRoJujwyyY+zAndHKk20NQaRrsrSWbjiyOsY36s1G7xUtVPaz
7J4XEh8R6h+r0gPmOKMIA4QJKKmJktI9i3mJOmWZdun6AF1gL45+QMLxGVBg
b6af9yp6hLxgZtXzWY8ujIKsuTgD4ZHCLSDQBecOsMiYMFUjb+P3fkagRgL9
iER+EKHkC1jjhLrAjHpC3L+bLOyYwwlhPyrTOP+fPVt5W+lQLlIgCfacJgbc
ra3haxk4hnNKnCVDSyXqe87Ia59QLzWPFWdfLn7c3Ru9QO9Md8hl1rGInHdj
ekVdzYFbaIy2WFrAjoNJPzphgdb5BTS1sZF3pcu/sW3O/Xoa9SfOcoqxnNbK
9ItjmmM5ZGz9dgf3peEBR+0KClcH066I3OHaViUtQ7Doi3zgG2zQxNYN4/GM
zrzpB96UVwCfbO1uDw4fU6t97Fzb2ZFFhvFFbyh9kdKVNFV+8afiHQZPpnWM
/svh4crdeZEJ8pUF8cCjLQYVw9pQkIMqkVoCug4S1XrdDZtvoQp10AI43wPd
LfUlNQFKQzFlArb+XLEHMFVkMOMx/LJ0E7uNNiPoeiKCLJ2dJ4orvt2+7YAE
VVUB7xqC6QdGhtdJcPRyO99T8peH8ybAQzZd+wkgDycb6UGpMEtVuqgfWP2U
7QCVCp+/zqAw8Td2PPbXfBm32ri4ggCgGSrloRFsyAWFGVFngYs286rSgwHR
mnd1kgRXiAZGXkjqPbYz7Z2sAiDlQxoXpX9uLRISM2myJ4BP7vVjR626ZCSL
faSJtWHdRcOnoBLDbmMGFihTZOEeBt1eICrqpCasxDBBI0s0EriWIaqm3TNs
ZY4+KnnkSSGgHbwIawSbneZ4ITPPn6YU46jtcaZaBgLMFu5mRmLp92ccZ1uB
7k5NzYrJ3sjokH46apHoKenIqrcAlrhXQs8whYgQPx1zAM8+SSaQ9EGZ4NSN
dvoxj2cxtKcXd1onNKd4oW82KNZT7QRPVcBVkHMOabqR+mI4kbyhbtwY11el
NBpgZhum7YhdFY0FsmOzgvlloVNa/pE4Rcw54HtUSNPjC3aZtQ56pFXuBPbC
bGZ9hS02fsq1aPm1YgbW0u7FQz/gQQxFrgRDJ5yRq3FHqv1NRkzpj+scM4uZ
wK+jcwvLXzxxX4yml2b51aHDDtTj1TX8C2IHsjYf5OWgIeXl+ld/nE65jHAP
n5W1IU/jM07Ha1k9NNPvG/rEss+/tyqdnwWmGQ2FdBpb80d4RHBunXtLqxb+
FfC3XbF01LsveOQahsG0KmOTD5Male3C1uuVD8AwXHvyqM8Bq3OI7KytXlgV
o4CDGorYbCDDKOY5FuGcJ4whks3eNzoHaLiWel2sjCnqsyo9y/+vPp+gQyJz
ISWzDIcQWLXrfM3nlM5B1LXxNIsMtFR5FUiy4P2MboB3TSQTaGKithknM9kF
97W7DpyMEZfL69sXxv4EmrmoQpyrQeBGkfjjKToQE0C/bCRqcou/Fh7pdyoM
e3lJ9JN0jQThJZ1Ur9yZ/aeAkMunUjiTqZdppClbu4cTgBayIw4J3Jg4C0c2
lWZtCt9AXr+xqG/gzJHq/VDpV7f0/nka7EJd5I3xmZ0cBU1ftkm6MAfk3W/o
CBi4Hzm3QilkLIyuIuwtpygZ7umroxEYv+7duf3ylRjGxS+8mG4Wus5BMJvQ
H/8NRUtQ2XwGZYW5DfLuGYv8871dmHHDRHRXZUujxo1KMXtUiz8YsKH5xE/O
3S/lpqBFJ5cwbPCrHDLUJO6GE3AbhaXcgEj/cniJDbcdYVk09lBz5nv8tes/
p/y+vPjWFEgWo3fEZqXSJ9r/vvE1BTYJWH/fpAcAxnSDiG/MNDXfDLkkKfm5
WFVSBAuBWZdEI9G5OvkD7GQGvc8gZI1xPq7gfBTERBcrdj2SCDzHtQbW8peX
Gvyn6m8N5zd7DHoWnGzZoS92wv2Ub2dUPd0UP4XAORNerzMv/wO8WKvapMCr
DrbRYm6nNCr9LXCpsej4YJItVt7GcYSJq8/hQ/75bMp1IzCaLFY/YqLJhyzD
289JAV0kuDCj68wLCniTkBuFO0cmKyOdvs31nF9cbbmnTZwJpqvBjy2HJkJK
Bv9kBxycKD/i8OzhWADC6do5Jf0ZZuy/xDwy5/rrz7T2Wj/Eo3tQlkCCqNkN
suOQU6xoTWJMP5PHVe2/14zeAW/0a5kCJt3HXP3kl3ykJEmKi4oGFtvv5+Su
/vvVgYplYizoctOaKc0iBaPXsnXQtkaGufRXlsBpPWh1Q5PNoUaBjTjig0xC
snP+gAhjpff7tXJmrxLlGbrPKBkfUi6NJY2vI1X7+038wb3RnMNfAPMLnMxe
WgEvGYQuGjCIEusLu2HxLrsPNY+4ovgiTLzmvnKOLoMuLzyJdMejkI1M2kXX
MDfP2rXG8NaIRAO/RQKrtsz6oCMDFU1DWmi7o2RfW6m6ylMh9On35oe1K8AR
prvvK0L1fpnudWYz/QJcnRyFAcHPxRoWbK9CwiKVEUiNYAp3c4hmYpVB1NSL
9gs0er9fRV+ly2D5ZKRnR7ov2O6BYBSK8mPdxFx5fq3Tc3JDw6x6R+xhSkGI
A1G0AO9Yug4GTbUC6ZFlNoqcDEuxw+gjI4SuXmKzF1eLX/41xMJcIb2ATSmh
v8xr23b+zFutyU3qTLWatwcBO/AyOFqu5m6gR6IruwzgUc5eM1eK/dAc0utX
V+AXs4R3XbOiVMtgqpMr6wuIlbENQdG1cVPH64CrCkqaxXFE2jCh5IcTglnJ
HOxWYWYC08f0BjJAFNt3xmJm0xWRtYDlrHM/aQgBlDxeiReq2ZBoRI5GRwwv
EF3Dh1WTwccX3RWLvN2mzujaI2TU1ZkKeYCE5zs6rzcsHw8gGr0G4OztTekf
i0vUxLsVUKcVY5ywaHGxj/GEDMBILhTYHZ5n3eLTaNixVQN3qBu/WE5oF4fU
OPJDxWolVV2bPnAprTHI5xbLSPX7ccdRd9X4gV+saWFUvL9pXD0/1qV8Mnr6
jvrTtHC3I0G3kmwh0ZmTfb2qb+QK8bQYb313iJt00bp9v0L80AsbOfBuPXSt
R3snn3NqIWiU2gitdzBhjCFEVHt/Em9Sqr3i4XAZ7OAZueYmTzm4F9st9OHj
lCv7BxnfT/Gg+mWcH8tEMro7A5OVf8VfPZBsd2IAM68lira3vZTbXZUxsban
EyK15RlMBF6V/9Oq73CePjevSFHgOY2dCOr5bxK0UW9Lk/QiGF57rn/f8N12
wUN+yUnS6nP9DbvzyxkzN+GHPKmhj+PAfAnYFGk2t1e2jPki5BxdNcR+M7IC
vG40xrYilsGiWFyx86DBlX/cgvbtgtyaElEW1bdiFAcoX1kgkRCfYHd7IXQd
rnXhBeo6XFn6BF7Wipj56/hPFlmSAM4TT5NjyjLFFH7JhyIXAvwBIitMURdZ
IZgpK+R3hjfuOOAYYBHwrZyv8HPBCl/j3G1WsPvGNfG76ahII2htrkyWp18B
HGp1x6XXPzwahs2sbktuEQgY+tS5Z6dWGN15AU3kHz+NEVDBV2IgZvlcx+Np
8tNQqAqUYReEAcN9IuVmmICBu4UHgK09Re4tJ9LRVxznKnjwrTzqYm6wTpya
jTIDiOBS4e7fEqKT2fNqbcLLpejjZGFPgJ8zH6ESBtDgqFs4wKOY9zKJBeF8
u0f6T8GtNkVsb7VMlc6icd86I1nFAzgfaogFrJwQCUPWgTmH4W24l2mGbN5S
qHK1+zbU8119h1DEgYkeAUVWhKRFKQ/RqZOblFIFMQBfv3Gf/1mGdc6ERhBq
j0Ctj1txHtw+rHial0XLm18yD7wHh8h38t3OhS02BtM9IalalkxiZdKCTFiO
3YCpUQddJwRCSl1THgdew3JNy4Be8G1i3Pg0NlfB9hDeQiFonboQr9Zndxav
F2aL5+PAgcMsnq5T2FrGRympFdPVbJ78MQCZX/F0sjsgU5JF9l/qB/7t2VbA
sMZMigSMcbI/hVIkiJQzw/rtcrDE58xTPWsX7IgVHlPfDfZN+iSY+IE0AcNc
KvGp9YhncxMvvWMZWa11IHcFAYuZR8W8AwdRi77lMDoJKmvlwI0d5tq3z/Xw
xSCOvMYcNlW2C1dbEFEU1Ft2Wjbo2LKIOXJ/Wx45vtjPiaP+zFrUNv8Iwblg
FTqHhoqYKe9UnSeeE3oGAU8tBZVvWSR+FRB3VHDCh3hxkin7TtqYApQdLSCU
10VewDzzzIUEQbCxfqnLDg0in66lu2TCZh+Z6wST6SUSdhvJkuWfebao06Q3
tnoZ/htUIVjHj7zS+S6VawBJ1UXlz/jpDtcWESZsqKJr7DMeDyQhZVWPWbrc
MsZR7E74ea/xBYXXW6GQgCjgGA5eXvHr5QeUxk7XEL3xCF5HH3MHRfj368Gs
B7G+NuMeexyeuLLDR9pF+jfmx8/1gcZY2vGJGJaTCBbb842N6grvrYvUeR12
oR8oFT7DHitXkXazJl3vNV6eGgRsrxmjk53fClUkENts8o3V2sYSmMUNNXjY
/wWCgkvH//xSUcYrCyt66jz1ydT7gRsTDcJ8h2nLqvX87UVGwFZQ5MjPEfMw
KsqMVahWtmurudcchxDK1cAAgwhiNzZs6cuXAdeNbI1W0+xPE5b+KpAg5vTv
BtAMCSg9n8o3sw4zkQcpa8Gg7qQcLKlbYdTPDH1QJWns1I55o/qe5b+xyODH
moYFKnQIpmh+mZa8RRjoHUqJCWCXPge+Z/bbc7/kDge5+3o02GqecYdtAylD
zmNkgRZgDfxjevrgfhX43AK/+KaMTyp1zXKEI/VFV9i/wXbe4+yysVy8OFwz
68dTDW0gHMhKM9b4skdfH9UyWNRX0Z/HzdYRXzNfEHYnnhjzXlQP2TeoRfvj
pldpYcb0LuKljNgj047fc/xWXAuZibr2IPwXAi/AnuGRaPaUWyOOlrGVkwOA
RW4gcc+cFfoKWDnZMhNhIU56YWAUMGYvLWC1s+CtmZP0fK2uexHYVLO4b0pl
/dkQUhA4j9W8AgJ/uQ/h1xAftIDrP/2bWowkJ95PncyMH3IRMtKb6qj2EAxy
Bu2qdErvUBkbs1HRLbgmXMzufwXwijEDb2zh6pc80WDJXiXK597yfX4J7u5h
EVErsjfj+oaJr1MhXA+hfDz53rtJ8oPHUmp2fzcR1rwlQxBKJ4y8OunOsRwD
LHg3f5/SNAGdDI4WN+tpZFu0YLwc9Cv/C4s1I3mVQGk3tsgV5+F12kYZWgot
K7fSvs+MqJH1hPouCRuiYLGYpvh5iNBVT1wyJETVZnEqWrsBpgDXH8UEFmXX
uO/bsDsMkyMqks8uQI4A0PyJEzQ3hclU1c97oj+OzHccmYC/oU9P88MEKGfp
56ljtSqjbu/AsY9sir8FTzb11BIpkwksTUTLtdy7w68MHAfZsdw1o0klnF4P
Vq2bGrL1cXVNmm9WuS+EcqnVyHmFpIRaFsDW7kXt+lOOmXtoF2hs6Bv+XLye
+e7eqYI5QM7MjLi1oP4ho4g9lMY/8CKHcHVIQ6AbZf+jABmCdDl6+L0x9UOe
4Iit2D7fRzB0+pYRcQ8I/Xq43ZhoLfz0eqw0P9I5K7QSzfUL2FN62ulUTUMr
cqnpn4d3Lyu8RB84lMhOlD5cpqxcRFAUS2pHukr9gRF5VjHXH1dlR/iFA/kx
2T+fsURp5F8I5BV+UAXIdssFHRo4zaLI3cqFcCCaQHeegmu98tQ5Mkfqo66M
Gbvzt7PUH06/z5Ljof4Xtyr8j//52DaguPdWbrlyxAI13AtEQ3XhWgymMpox
QECT2hKQunZQLIL0IMCQ38N35PlcTnarzmmuEXmyUGu3Ad5eaDxyfP5PjM1j
UrEOjeQE01gQo9sMq1zdOwIZJE1S7kTYBhZQnDeCLn49gdMQMix5w7pCuElC
HmbDUKmDf7qEriLeAh66YRksVBv4llqMnlKijEa8RS+AWN38FPagziCEd0PS
D1Q/57GqF3meagxtDJJW5+JYFp+f21JI7uY1V7O8m1VFhDMYwy6MX5DIMXmd
v/tcGWalrFFPt56kU8J8c6p9mf/2C4usEf4ChZfJufyTrJw1SAdwBprYbX70
HJATeCbVSQ3CXz9baPSAemv57QSJa7liACRADkDRjcVrrVwVU20V/HWr9Pvh
Pv2AHXXQIK7hYCTlYLVaVXXns8yK7Ns3qYYL/WIZ7UnaT99S7xG3v1xPctjy
eEmDg/3QlVejBr4cmGT0Qd2hv+5ckxmJWhBgIiGPKdjFiP0ekSllYxuELT5a
IHdmwubwHKvJpTdgE/9fti3SInkG8qcIozEAby398ApkFEvwwGErSDTfOg1/
tA7MUm2bI699TsttwjbT+hUhBLwaC5hzSkSLNs3u4Eu41EWy3qSn48KakGR9
drhap0sEa0iD/apLJQF5XJV+LAX2T1zVC8YupiUljoeacuAUjQC3CX31hOrl
ddSoDDD0DUF7jzA7yLexLUobQMypF2XKdei7pt0uXqu+Cw+zz+PyhTO6x37J
DyqGgI/yyo4H1A2YHmCCyygbabySDGMr2RRSm1SZjm+QTBMJMC/PyDMbDmVu
xHKxNKDyvhc+UxucFlmHlXch72AS7bHxhyT18x3S+1mN8croNTyaXZu6wVMq
3rcBV+eStvg6iUMNVrcwAmo7qF4WbiVzb4+BKpGRgYnKrj00KoXZMeazMFsZ
/FWPRjBu1fZVS4bl0cFIzxih1pzwwn3Jk8PnSwTRP1+93dmJGxize3nd8gyp
spO4xZ8wXU5vIRB20UH3oZcIGYSaYq4R0k2j66Jc5XMCCPnO8b0Ep0uaR4TW
U6ym6ifFARnYGYOk8Pb4LTO5wodb7tqD6SAbAfo5sD6l2vVYf3XhSRLxiwHY
Mn8AHHr8OwGeZagro5QleyhEG2L8q/+sbKCmmBj+wNzLa2JOKCLOousSKwRd
ALnlX0/URulUMb9fopiDYpuBznaw6RfITLlWb0C3bB1lenMnKoJQuE7pOpYz
yAwbx7vEiJy1FuyjyED9ZjTo2JIxWYtqP0zbXQFYtJJl6fVv6RZmVPytlRi0
8IeGU+M5Neg3ofD4FqGOBPJMrkoaaQ3cLGTTghvlJxXOCdrhlwLBTeMmk4Y8
OdkHoqhe5nXyjpLmQgFOTQ+hIDa3w5nPpLBlUBPltbw6CUr7D6w7cPzehsrS
h0bBbomRpMLPrvMNAr34SMP9oTFDBe0y+LKrENjpAoC6gb1GECf8SKdTQP/D
kS6KeFzL9OB6JwTGjG+m3/S/uDR9visbQsXhCuXPMO8ca8dQtdYE22eQRNVp
OMW3FVIDR5fBKzcw5lQZBrLAjbeIiNDIVEDoE/mvmUZOA3k9ISA2cxf942eA
cqe1XK8wfCGXzAw2mkkSnha5Wd2Y9LK7AJ8/mNllN5DKap+RQjMOQi5fdzzk
BtBVzSB4VbuCMpoIKYNKcal4963UdrGslXLwQCKWBABGbkTyedZv6JtXcyZR
zFRGh0SNcj2/5whWewcQUdH0mWZPIGb/kjVsszpqUQvjcJJcI+TMjJN4Ga6b
4AACsNWxyQLEqIrQAcVriiY6STalZCAjRFUB9uHJoJQWbFq18B2ERawEwo6o
ApN4MNli15OkDzXCyZp7XKSnLxul9FiC4sbRw44T1olq9EPR7yXBQo406XoK
YzDixgi14wHxl3NQufi5F0KwueB4QhG/kdZVQFy2L5Q3pUy2sql6Q8hUcdSA
axgcrysIiebIOJMILJgwCqwV2UK7KeiBUq8esnrcwBRLWVr9/EBp77wOS9Eu
XS9p6NZY39qcfoADIshwBfRrMv77yOtrt6TgWDnk7uM6NX2HrMbcHRg42GbE
IdBTll406dM8Pp9lNEm//yrw4ZLuilbzYN8T+clqKJDs8zQDiTQG4TO8zW6p
qB0sp9HD/FzojL+AnCM56pqbxyAvqqduZP0DVGmpW8TfZ4lJ+RLNeIMXiuXe
Eo5iler1e7dJxn330IDetsQks4QjbtZMqLS/Xmy0EhPCEVInMxymkvgVba04
vW68nU8BEPn9Ac5rXSE8dfpX9lmwgopIGUk5EI1zqyCq/dD0uYjX1CO+ilQ0
8oK2jtRAoCqzlhuiwEg5dRCFyssPdrno9sfn4T8WFI19ZAtQkI6izWsYvTVV
KkBiP5EMQpDXR/YaLacACJFxUX0+ZdX8K2jDI/kE2w1lPD3Q908UFHSNI/iU
kSOBzSa4crMoMWLSR9o0yICgei/e6qKPEJA96/PEj2sGr6hm9zt+wbBkANx/
16qZbrIhqnaIZVUDuLXZGV0tU62yvb11TCoJkrsJJYF4hptuvRvhDx3ZPuq6
Jviu4q1fXw6IXfGUFdAuhJrwvN9uMX05vDUlqdDRPC9gXKnTocXnzor7A39U
iWvuG1aofgjZY2XAevnj1pJyckpLfEQQLZvmMTPLjLzfbdIjN/7wrDXSEizl
eSDtuhhYJWSaMoHDatJt7QynR+Ir5YJN+cZr+4NcZLoZiOBWHZZhNGJODmIX
74evGqHjTcOM5i9p0Vk7iUCEQb/0aKG36OSJo142DJPLR3dgWlmIBfbSI++v
ZtCpdHmHDcaVOeggBH4BNM6XZ1Ri2NJ6dIe8MdI2QWEgoWhkJ1VDbwAh/DDP
E0YLcACOsHRgqsVG1UNOcF42qQiTv9OqP3WO8X9nCZIYKXYtm/Mz/K1NLDWl
LTJbbzVhcji3TQcF36mrBPgOzrzmmLk1u4DCzM1tuv9OgzPc9boZUrvJtz+1
SugcuctnTJ+uSjWcm9GTpfh11qme+lB1UUVUB0ARZyzjt7zLIRQk2G8Fc6D6
xZQtYnW+RNQ/pOtTdweO8Hcthlvyhy/A7iKK9dXUqp2GPLF0SyN3VX3vSQzs
wyVCjzP+rWAD9gEawJBgbvCm3jNpF46/+217MCyL8Z+odnKlAKGgE7dCf5qu
2uyMTtca2uzKOKWhT0jO01I40HmVrmaVyHPzfIdrAd6GrTb8gw6aC2kNN9ZH
y3Ya1AG+f9BgLNEYXoCU5RYmxXb1Yi3b61eHb6ULXuA7OWqODDo+wmEGs/ck
dRbMGGLbEPfuu68zRN7Z3KOzFbOU306buwShQH+qpz8/ZNECjq1prYgkYnXD
IsPMWQm/To+eG76FbR0KK7TLMOo9nWHDX7opKctN3tw4nW4NsqQz/IKH+87y
/gESvVXxvhg5HhJHs6AAjVNsoPuf1zAxx6Q6Ahbw1k1FsdOS8EXyYl3FNVBW
jLAsMDoCaG3GIUEZShOo/8RJRsO08kTlgSWYV54fAQTK72NeEW60RVnWEz86
ibxLrLWOuvwwJ8NV2G9tHHZbQl7M30SXHjV/oDR5vHnSZ6jB+WDurpTD2lHv
+PuGJ3CIJp54K9WRYH4llnbkCU4uxnq8rxnt7ll5RDBF1QmeDSjnzmozmcoJ
P560eSwpNL7jcUuxHOVfhLTrN1JD5xfuadxXkcEWfE8MpBfMhgLD432iee/y
fDvv50DcjogfwJ0DX34fHf4yUxjC9t4hFsaU4/4LcS6huQTgpT6MYE4N/+fS
0YNSbi6tss5fhly96uLRBZ2OtCiZye1dF0Ec3j9moKY6BVILvqc0OkiiKGsx
ouir1vc6x+tN0OV57Os8iv/e9S+uC4e1CQyp/Qi++7wXqx4sOIgIb0wXwff3
kF0xM7hKVxzIB9OzWD/J2+/GpmVXh0F/2s+Hfv9U2gmr2yn1RlD8ui80WSkN
Y78klrN1bvuVzPhhC3yyLKJXF6Q5i9OJlfPuIlBs8MjHPw+j/9h6GEpO1yWT
9YR0f7MEKA7H3sjaRhgpzr2vJ6kZAylqc2nYPUkRxPD3GLg+i7CCZV4Vsg4b
fq7dl2hcIS6qlU0C+SFHCEMNv2KrcMtJXC9DQ2bC33wLIv9zJhsXTuyQ3y8r
vjsAtp8xR6C/6Mt4L+urDZMCvQVGBFWzgewxjv19KlpPnJItwXYnY7WX9EmB
c+Kmquqk67FrzCUhRs5qxGjcuwqWcnTD9I99DlIWwE158l2QmxLj2F+NdDKh
/qn4ZFC6RxSg9bKp06TMdH5B8l6z5Sy4AZEluSikW0vFtYwskRPfpyOkUuaO
wKnZeUnHnPd5Io6+5+314XeO1DSR167BBWL6rYlJcTUazLeMGQrdxEU7ypTc
KIIcbjFIgkWO5W2l1T21a1YHrna8nVp8Z4IOqR7+4v4pYiBKPt4GcQnRTy1C
UeOJD2xTTUGmH4jJblvzwob4S6f0rkIt9QKUrz98bAbqqtGX09aC75RhwFiq
2+KFBepoBl3k47bgkL6QjAHfQlyKMGkCgjQ4PM5RGCwMmPEj/lkkgUbHjoFf
06jQlebF650YOpikQb8ZZviYUXFs6MYfM5SgudvHTBx6ws8rTugcbpBbmXti
WIN7kgTraUieLk+E2K3rTQKl3tsetFzW9s61D8QOREmskGVrMLf96lo5NYgW
BZuNxEQhBItftc0ezNBqefKf/z6pxdkE9sCWbBJmRXqARraAy1q3ugJ5xgsd
jxbjlYBKRfzH7pZDn5DeD2cIbqiOO5obN7pGfYnTPc6z2lPb4K8CKqHEo3Lo
Gekx1KfzqMw8EISnS5GNtnzGphQwff4he2BeRKWFybF3E1yzYPrZuUS2wDU6
JvDRkomoAg4v2I6zMfxBpbjLFhvEnpVxqKWTWD2ePTWRi9Se+ZOdo7i8bJTP
IfgcrTzl5q6RqcDZ5mFKxLSZ3IdQzbswRO0qsaiLjyvJUqUGjCcAtLnX/+Rs
iVUT/LNSBvueykMku8K/a0ZhNYZ20y09pQSK/kC5ThuhiGUzw/TJFFJYdcVU
rjVO7OT3K81VTaEIqSEnMyNlYEXmG2HJggUB7PAL+4OIz3db/smuOfVL8SFK
LhuYHDDJJIFj7eT5xfE6deYccGN1At+CthnOzvC8+dHtWS5F1bK0iW8vWZvK
Yj2lVVakaxmYAmTd9aMm3NL0WNHTYoWHXdwalrcsQNDCjcjekDN1Y3QTWQd8
ogdCDnVXPkIP0T+t57J5NRiHbRv0/atJpS+Eb/RYJiGpbbknrqq9bo2UfLJk
Yf0OSK7658G20eC4H2abuo6S3d2Cpy04gOuMZnC9DBZ4DjyZV0RaAWKYNyXK
QFLpslaiQ3VxvpihY+TKnYP9TZPzRkOxo+NVUQxwfyWttewHwSq++0a9+JlN
uJqmwrQHE2qQhHlrgnMIeBhzltQejYiZeohUNMxcnVu+P1jMLYukuJqSabt/
VjC0RYfK9YErrlpPT56Nf95VSw27UUO/z3EpEbg964fg2jK8UEJ0CyQCD4NJ
d6lq7HUmMbcEoh9+K0W4B82C8r41xW5aiutfHUOcyciEhXSZUhjwyum6NrDk
wzxyH/22TZsz10C7lEGbc9dtkrjSaf3FXpBkX13kBbgbbKSjOXIKaGY5wYAJ
3pAzAVjrxprYdrIYJMm4HDbYcGOEALssB0DgwxegfJPI1u34dQH+Su+2x8a2
IBiefH0QtveFGgXeEhOJ0+qzNAcHUGxv3/s0++hzzf66H8gVvdx/kdLknXx8
R7ccV1p0Hv7137rYNlPEpniAS/d2nUnQ1U+A7E1ErAEjxkgC7sx1ELea5GXs
mXm0sgm4kemTRSv9Qy+zuMAB6fLvLkTLwMi0LYcQt2uSBRLPLs1up1KqtYjq
xMKZ5xO4TPG9We3j3QJpRXbLRkD9hpyxQf7WXKZlg+evV6eWqNq1/D0wuWCp
Pf7ph92ToREwUtAYtjb8xdG3zzp66l7IOgksb304cON99a3O6jr8oCzfq/7C
CwxPw4SIE8tkmgO16p+kI2KX9GODpwgw/yDX/HH+NGOq3Zj5YixFtVBdBKrt
eLlZp+Kz8IVLwWhBh63yENTk3n80YVWjmQCygVahEH3m386+rec5VL/vrT6Q
YrhrzS2FAIAODjt9I0mbrmYRq7KZxPkDrxb5LoUodV5/7bl6TMc1rZrc0eHF
piXGvUUoQfFokcweqdUl+2+3DfuUvX8qNKNO48ekTdtzB4fLPcLfb4Jw9OaZ
9ziAZUTjXCd2KiS0Dpc6TlTzBKKRdgNEhP9Zc8sbjf7dqaK/fFVygsPCCJaP
ML3MrJmmwXj3vywYBWFpm+tjzSIumPPWOXW7kvEXUt1tN0ayiEPZDt1VspXX
2uP9/mfLvBW3f5gkSmvnb17xYdH61hcFk6ncMO7kwhCfOSNYfTPAmeScFxJh
WkRyNzGrH9XelkHlYfA0v8WmHfz+Fq2WqhwOze8i1I7ubpURyRA3o2BN080y
b4HcS55Vj+Flw2jdR9UUDMwJEgcd8sBy7eWJoPpDSJlQ6WCHpHVAf0xBVpVJ
NMlDqUtvdX9KJt8rBwN5PrHPzm0EQpPQ6VtoKtk9dPEaIn96mmqdWXG2k8oN
RjkFPpU0dVrNA9rgixIWoLO08fAgLIlFiI5yCuZrKOvX3q+2G00Z04/ZDMSJ
v8eaEd98tZ5+cnNVSAgWg9m+L4eLHsa7V4tvIGjx8s9IfVhLRKQhpEDtsa8O
wdtovsnbEiHQwjLDaYpq31lMW+bLQ6X2TYskvia1AQmA82bxGgUMp767yrYA
TuqUpbTI9tMSx9slREe+8cu8eYDl7XGhLCIfqLnUZvviCbvkZ18igENC6w/q
jll85f5siFG5wzP2pB93jBZ7WaasEQVcdWSVV/lxAkQwlhvK9qhxeg8fO/vu
/VFq8PbQyCoH3C9k5IA41XIJ0aBwV49eaX3XPezl4V4noyCmQsGQ17oFti6B
fSrBaQ/lQt2ByQCWZdk+tKBe6sSXPUUTrNrIQ72z7HNBk8BgDDxMnmFdAfca
nO2wlzq6J8mJStwIYJDBPlQ0C8RKcT81l7sMZ9SHOiNE2hQDQ+UZKprTUxSZ
X9ULX3UNlUX6B629L0iIV0YzlbTocznUGGYzpGjSz/ZD19trIGol3JwqdAY6
k9ZHxPuYah/hwlov3gK+aYJTJipKyZyd+PJMUBuGS5x+QY+0pZBXnL4GTg9D
V9MADsPR30RWMuT2sM3YCN/GyMu6l2yUnT53J6USOnKQZxP8OgxZvqPZJKl5
PjIqDQ/YVU/2+Bo4bQ/cct+4atbhtb4GRukwey+pJABCT08bG+oqhI/gh6g1
82nLqls9GEip4jsVZGqeaN15b4v9kBqxB/BaWeQdCylCMw2idtIqb7MkyHju
I/fIFswRZQMYR4mFVp5wO+EkJ1n7hDikwu2upgjyVZ2CSxHoM37eDh+YAP2Z
US2vRuNfw3TiCCgCYC4UZ7heL7f6j/NRNGPQVWv6L3oQ0OXWGjb7XnpN7AJx
J0HNR9bA2Do80SwLj2+Zmy2Wvh1g95/lqV1KXES/IzQrspF8Xz3S38L+CF8N
tEsAGB6iOiVwvo1i3wCGDnuCDh6McqldptLBgsuvlGH7KNEMwB+aLnhPiCvC
IW0Ah4ZyqmTnpv/M6jhrh8uY7f3/g9Spd/+UkLLcZfwGawf6Rih86yirlkpO
s8+/e8qvq8967vZtLs1WqTKWDhLniqcko5Tup5wWD7Iy+zfuWsF3ZghRbb7Q
/uZq7y67DiyKcVMgS4EwdCWO1V3dkV7ZhohZzpiS7KSYu90/YBw8mFNsc9Iw
X7bNrYLs18oGc4UXQ12/tlVPxtwQYmZRuaneP5HBMPSpGeFnksVmcLWYcPlR
lBAO1Z59cNp550583HWghXwVhmcX9/6xJD58zhmpxAWzvKPVoqrIYVhOHcdB
7fZW6dN9kVEbzFSK0fVZNsyv99fhYj9R6Vl+C0KRF2luy98jWoG+xuUelQxZ
ZPunGdzH5vbapI3Hwk3tKxnlW8X9GSX7fbjk92prVOmb0LmSWqA+M12WhrJW
//yOsicNMtkFjUPNTHsiV0nlIjIBPevBAUkJ4J6LlPMGonjD4bg164IqCIXk
f65yVrGmu4QjiNnzup29wUa1jhLjSBkP5LQlpFBfwExRftGa5gIuAbV8Ua0S
apmNIILIIuf6ct4sngO8QId4CYjWIWYcnZddbR09y7NWLutd8ddHq2z5WFpT
Kcz+MPNVusqoc4Ez91tAJ3JItiP7UphyX0G72W49NOtD9RChc7lI7wz5W+my
TDFnIGNoGKNvI+Cl9SN3c4NmiKNxaHRD2vMkHJ/Mp9wqPW/A6TI4sMp/A+ne
f/Xfc6bnyxPes5I+kN78IbdKr6VUlzYS9qVqr7f5kUEmPYKJVfb0gEr1VUfz
skQSnMaG/Tk0P8uzPFB+6qL7ldepK7YkWhpofmid7f69STY5KPuKJYdhvZpN
vxR63yYtSmNk8VluveLNSaItbvPQYCUhw+CS6jRptvydh7DYyMbFeVRlH+KH
ZZ6+k9QnL/gqjYoJSBz3uRajDmmQ12tRF3nafcLDKGWO3cj3wS+nB7BdA2P7
oUQEtBNyYo8iGthKtdwNr1PtXt3ANnUwHvfZu1NKT/OHG6RAANtKs3n5hRKD
0jhUyJsNcpmaCuJVtIHoePvl05OE5a1iqhMCMtM43/4+2rvYYtD96uQTRraZ
8sMlqjxvpFF+kclB2ytoe5h7T7J72bIeJqKsaSVgSu342AMFHiWmGdJ3Bxmr
I5PEHjCEHtXTanEb34eJfmSLTaBSsqJNhv+wzd8jF8Er4aWYuggAiC8DAeQ+
p/fCwd6r0mlUdRiejpoT4knfUFUyZUpAJ/qHY1/Ir0TK9gmMUKnlBrm0suUj
R/uvlY8bevkxqlUsvqSdShdKWevI5rv1DncYTiKpvp5+sM5Ay9h59z4D0uSE
8hitsP9y3OC+h9WK4jOCIRM5rglASkWqMgR7mxrjg6EOdi+02PRW/HFsoVwl
nl6HX41wSpiv07rzfDtF2ZyIo8S4ATeIRnCJRs8HTKlMxDIk2EXJnwC3F+dc
rE30O/pwhDZRyoTw3P9xsKOTM+g2UpVxzAp+Yko8/Zj5JKflT4bmuohcT9fg
8uIkdgvmCbhkf6iCHXLEK3t1S4bTP/H98DuccgptJV6/7w38qnF9HDi+QCh+
NjSYPLC3s0oSwHJ26SRPugMQnfuI8NVTjXpgx8qDYED0UUJYrIQ+rJXLWrB2
ffNELhdUHvT8FZbhhavRsesc/vtk6X8TVEn27/q+IYcKELYPCd+GnY4RVB4Y
G8xKJy2Ov0kf0n/xl47UxMkq2cwvQpdkmBadTCA0wbu516mzWelJos3+Pmxn
Wr4dqRrrx9b2yGPILKJYuT46+oyvwBbGfo6IVTWEdY+KqGRAG5o9hH/0uuGy
DgDnZCPcTBU0be2xbiybVCjUYd5z8ooir2G4i71gEOpwWdT91GbAyAI9bnof
XejLiCSy3ViZHenTgtTWJF9a7nNLxq1+0GEt8Ux+yOvRsIz1iA5XkZUnGsTN
7beqJxkiTx1cHGMZMf3BCfBSIOuUE1gDdZx4XNlKidXUZZenrCUgAJG+SDF7
+usmSKH+tYHLrDYIo5GaM1dyzmuQPhfgKpopUZu3GfquU4DvEijAWdg0gcvH
KcdIiciXCFqqk8LXuYkGP2qSptdWCydWn3Mp72uisrMRmqHapud3Xvt3Y6FX
sXZOR7crqqZdqBPNRPM/KoRvLhmxgcSAJlTd/rQf6Hym4/vR5ZXavw7sJUq1
v53jgfLkXf1c+87RDc+0WpZXFGM5SduTGLm5wFR5FGqAJQfq1gMHd8PgBN1g
k1XwM0BbrdWn93rIqf/kpP8U0sRGznYphkKC/dewAASDuqHS0zqI7UdUhC7i
I4lj+ecJsWyeZFRF5bko/gQ5/Q6Vv8TtFtKsniFf7PJO6Xpc5ufRBsYuw4nn
R1EVfuKlgQzIXFEYNGrdHjlhx1yZ8bJziRBBCaLp2CGIuQINSxALrmn3WLDb
WATNSMHQyWBJHmeFP+LtcK7yzhfG1Qt3tZQrzaUw6wUfg3RsNgJHffEvBC2J
BNVXoWXGebP+V0USBW9/h+syBytzx+kyei2cAINL+Y7csei5AB2d4SE/LxrR
2yP4srbvJEVzryhij9bcqu2K9z8rlbXoEv1yJxsS3KBUghdoaI0/j3UOuDC/
5ik1q3VBFxErBAt2QE5tC8z3tIQ8qZM/sKYotmCFoJMsavKQ0ZpkaytzU0eG
fp1gbRPuowumzJC+kSjPbtNrNUDv33TQtFhlLHQfcS8atHFvw/MPMkkCqJKq
TWPgczCna6bmSZ4ESalndGGXzn/p5W/S8PiNQ5pEQoVxfXgsw2fl3bYjuqoI
AoLluig66AUeL7GFY8XrqUja6bAYALAnVDn8a+YunmPe9K/jK0e17gPxG9kK
Ws05tfGmyFeRL6vEGDi+dc/BF6wEJySGR5Tppe3psHxFxkGsFG7zkDBHaoGo
1gvuT914rATeoyTY3bfq0NZV8HBM7qr2vjc9KwAHuZH6Wha9QdHCN0u/1uRn
drJUQSJZJRUovO4xPpeyUtMff7d2KMiyIRL6UE+Lb5zSiu7gI7uFT97K/Dlu
7OVKBGlGkNaqw3wc3z2oi0qQsh+6cT+p/fgOlFSBNfloxe9QMGak3OSsX88K
uyfg3QZczxm3JV0XavYhrxaMBWxgmjOgjYZSw+xL3BBTFsblj5NmCn7YM/1l
aLZkHOliOyMiM4mT8dZPpreUV3MwXwSkDedJ/2+WLizR89MAX9Yq1C7m5Y9R
Ruj60SltfZO/nYjksbOmk3nH4vAFS1Ijq9MA1Hm+tVPUf1wRGHScvUIit7Yg
MO0Yw6pOWa+zZAhS5hoLwdvtYH7eWp/8zx63lk5nIABInZyFeiHzDJn0RhSV
iekDQV0q8RThUvYxU+Md4vwpR2Nfogpt71nQoj+UvMrsavq51KY9+vS5JJVB
k4G9SbzVN7768MrPbgEWpq2R7qNDaoeZm/pxiZnLC/wReermNx9K7StNNGXg
lP7lTeMqMtPZjxMotulAQZRLfc5yLsI86iE4VTw1tdea/upNfXjCn7WXOQY1
Eia8RWo8belOMZZQoCNoLc3W1QBZkgF1hlUdjeryPVCA+J1BCKa6E5+oBc38
oZBCyyckhEke7Nqlgg+oJj0mstllwUbePhyk8kfbD9yyOOZwiEiZEH3SuGbI
4UuXBQsrlM9Xxd5Tmlupdo63OseJTwpfAuuBvlMqWbIH3vxrLAoCnhDZ2UzS
wR3K4Snh8lWIqHCpl+aNDoLWx5WV7hlHMLfJzo+tgFbDeQMYjjHYXuP014z2
//YbjbZJZgUD2ADicive6D42bXS5/VdbJVXThhTZ3qKWyWd3CPht/Z75FTyP
kmsrWl0nBulaEV8M87JZP6BRGJ8n4rLfZaAIWSdDkC2vJ6YsNxJazv4g8V45
J5/Cpp42vQ9ROp4UPs1yoTxwStJCtvOogE8veV+hXiZdrCF1jCLzHwYmiuPT
BxaGdQRUORtTkTdtI7LgVR1Lx05YY15PBSsEPEU5mLYQm2AatywT0jen1yiU
aYjZ6GDcf7J6LMe80kcgmPv6X2/k0F1Y5n8buFjfcXcs+2TdHrB5o+0BVpWK
BZctdnSx+oMyHp9z8ChJSus/+T/+dgYe6Yv+69Kk2BGEQCwFSxovvXvK0q3/
Tz/rJRIlRgyMBo4mMgxCyvJXixIsyaOtEujbb1zUaCLq70g9blVAfcDT8Ehp
2ofLyxwfGW8OyNXF1DbZbSMr+SYbEN2GDqSJqCcwxqQZpDtF5tWh79ze8Unz
AqXkubzm5ZsCjNq6LLBwgqGs19KURKi5y1DQXTQdz2ASqrcJcYxXgk/uKT14
G3rsrwxnZ1fATJMA72HXcFXyiBn9pt5Tfv1upZi8mpQ/43+w1oXlBjolAmvn
ceugQbcXeDZvE8/Bcd+Qqtf94eeA8uhjwDUXnIwwQTIVUIs2EFwP978s/iru
zAH80K1N9LqGquzeTqKHoLlw6NnXc+XGeMaeN3CC2nu9YT91OFfl62bXnMxP
+N4yEa4hTyupBge3qFlYbh182Muz3foQjb0ULH4Wxqpn8maEViiEMKM+1JYl
+DJ45U6/GEqgQ5QRpAs4Ieiqv0PyPO500Aq0aR0DokTi3B4EbzSGsUxaezrW
8gwQOXYx/CMTBjbuL2FSeUEpAx1ZMRfDDRY70K1la37Y6PG4a2zHQIQDE1eP
LC7pOC6bbRnOT35IDS1l+CkHZZyy0nx6EMiC+BO/OBEhIZsUsWZTj+r+TiqC
bz57Nwi4inyqCTq+qF5roFuHu+tRg+vYVjgI7HWHRy/OvHJzA3inckFzpAhz
s3LVEqkT56GwL9+pn5UySwVlssz3xaBz1OyVrPXga5K4y4RDyWdvFabydvW/
fckyAAiWbZ89UBGIIDG700R4mwNleust1UxGIFJ53isKR7n8iOL9tXo3llRx
a+fQ140/ihKsHELrlivvjeRGgBx0U2EgiJBiD363J0qc+ipxK62vMB1Q+9nD
ZRjxuBXkf3KschqH21uieveyvQWjOS5Ox9ZSKxKEJ0ywzhSo/1Duz6WsJa1C
DCKyonMe+7r/HdcY01R9gP8lAFrqTgPGWsFJt2yKwEWBCk4/L2y/DyIFm8SF
rfMdZKHLMtO60nWBgjWHMJqbRi+k9yHQRieLJw92i9VE+ZytA86oNZ1FOkNN
LBJNTSgVGaBqJNXuRVHPJMusRrbvMChDYWxaTi7GHMejVHPbC+BJAOWO+68y
VuwpMx1FlzojcfLa178hVL54ZgPS8BNzklx+tpkiqpmLurAi1dnrGAkQLhZB
NKi/Czx0/S7oNVWnQGKNEquGYPoEHwxfKMWPy5yMEBqt671DCwjorBe5t3RM
ugCD7JGh/P10kezwu5e42hspgUjL2L6++3qDbRFJlmUQM3rYC1IfIEglgW3Q
CcbiKiFcMTKOTRibxeZt5FhEQb80ZJhpualbuq5k4ZooCrsgp28iLRJFzNLN
biyXeKiGdm6V9bcJLhVajeB5XZIOAUAcfKJoxEoq/Vvkw0x8elafMYJEjDZr
gCcdrOLaWsES/GZTuaLL6msZ/SP2LYzQNiAYKPmcRSakiDG2D6L1xfJGxk2e
tNGdcwUOPTIMHHvk6MUWTXg7lZozjAcbx8fhcRBnryfdcGxHN+j8SeKNBVNl
90KyXD7Jpavr955xsW2oox1gOps05PQCTffICWa16QhjQHtcU1WJpWxH6gaR
tFoDOEIrUqU0HaTtQ7kuiheevA2cUq31K9mhyadinWrrZX2fcQQO9BwE2G6L
l3JAd+BN2nPJbup2ZINkVIiy/WJHZIy/qDs6M/tRFsGX5TNIFNJyDhGkGzGe
G/3ssJ6sXnUkFj4VFhWsKdiHcZ2Lhu9A2MG+qxSwfmY28hBUDZ1F7PadyrLJ
/6jHfM8krWfF55cyL19nL9HqRyxJ/3ddWIyO5fsNBIfWZwKJR6Cn8fcqXUor
7DiCkHLE1MJ1KoqCHNV2znMdgKcTjExFdfIFtz6bFfzNb3d625n+jKb0hrdR
zDKvX44+U3Xa0NCLnGv1wAbEduxmsEWStgNjGySmnAlz41wJ+5w3OuaCMavN
B8cFXevksuuMtzaOhw7psdTiiFf8rfWa8p2qsX7qH2leWtLnWnqPC9yeQRqb
OkeC3rZzy66m4C7RRtSX1DULFVQs25NvyFVZQUeogmWiCnbaoET3wb29+6R0
YgLo74+IlRhZHMXgiYejgkP603p2vrKwBnEPHeXts37pfR0FMQQd4guCSb3R
TFm3Id8EIDHVMh8U24JXj7yiHI5KMTvlJ4o6y7es6a2tdcZQlcugAGQ7ap4I
WqPcmNdoc/FRE79wIX39YnaWHXlGGZl4RCqnsgRAYuBNeVzelsi1LAcGpHdi
rBUJjiQVleAfwCKxUSlgzIBb+SPk1tg7sIGrucL2r4A/VlOu9ANdabErCuER
aSndj3/A0DoTJPSNmHXJaDOF5bFb1iqFnPGx7JV34dvBGHVUvF5sq407u3xT
/h1nEcC2fG4j+BYRupHMygCXiRnNXmrOAgBs1GDSl58aAiSzWODQCAaazA38
qcj9gUuCQ7wZnzfPjsWmOPVWehHu2v4uU5S5SOfb6CDbHEi2m7c0MHlPOW1S
bOExRPKkfE7V82srDgfUqsMeV0S/r8BOiA1FfV2Qp8xxNNePSSVylpQuVWmo
GAsfMT9cnVGDQfxRRUVbpQ+DIg86fEHztyxZuyE+aUWNpPJ1d2Db0THCU6kW
tF0W9Z/tr2S6mri9hYYy43SnWpWB3XjqF1hEtlZodqwzl24juLeT0IGaOlaW
pQsOqEtYBZp1D3Zu+f38TP4W06EBxf6glpnb4WuVhlIMFazo9+U9vL0L/lfo
qm3e/WyDvOE5tJeDeqOYFIpY98o+4vsgXgZeC5AbrHztPxNVHnSr3GUUYb2i
Db1GNG/XlMgpaRGs0+dwAjKx/R/phReJKRRr5fE7OIIDSK+E86KouJRhQCoq
VRt+c79ZcMMY6hgQV82IkwXWChHCtVaDyLzeP7uTYB+GcvAOgsPg88BymKz+
2K6Nby/U3PEvZhtk4WJWKRLr4nS2Z9ZWlP9bmL0xKelpniWMJDQnLtagO5Z0
YEVvXIRod1Au8eM1Whtv4H8thmdP3NsgXxsfeogcUb6Cvr0cRVgrwMjB4O+a
UhwRVR+IiqAMNqohQDG5YGRKB3A2kfyxODEIxjSSyQpPzLdR3NT5oVj62GJP
c3oQFdbg0DDBibzobqfstFygnh3wKFsJht5GnVu6a1YwSUssUxeRu+OUQFKl
qoiVJufRjeTuV1U0UkaoMeqXHTPS9qx4VPiMKHkPY8IMB7SH5jr+9WGwRhpj
i2Ojox67QuhPCz6MZI3UvfQ/Kb0Xa5MWfLqIm4k5iydLoH7xHfi+5VQE1anQ
iUEMfiiC26+ltLfWQkvFyWqiAzPX9rKCcnWx2pzRi3cqLyv+TjftPX+mt+Bp
YBUu3xCUK2ZaiBgevepxTueF3OuvaLO6Egs4strjOeXOEV9PgL48iT+mOmrD
oVXN/GI5j1+vilytE4cZBqaUsA3On1UKmOT/aaaVj/Rd4bH2DSuBEMRUERmH
/0eGheSdXgrNNV2L17gn1JdKACvq6JL6/LLD+F8kcJNEbLXpUUVUmwgtLgzP
mSPCumvUO4T+Wl39/ocB4OQlmy+S69IEzCdhVV4rAbEj/zUNUIUGdJayjjW9
F/s0+KKHzaLGu0WdU/dZp6qLOmIXH5lC9iYCtMT+BasfSkl/lxO+dZ4azapc
3jIbGT373/NdfmCfr5DxSFioCuhc5YKZU2RN0TTePTIqs5VxdEsH9NKSFFuL
R4K3fmgUsrF8DmadyJokjarJfgho+SIjW50VHyjFs92Wsrd7uejHmy7zBF14
VO6MtahS0X5q9Do9+mXvC6g+hIQU6LdChFJHZ2Ce/YHRtfyOPYZBd12v1S0l
9aavQImWxThPDcE38GvzWlgKeiih57sxmRKTu2kpRJnRl36O7rBMbJRmtXnd
gqx0kLe4M+BxHGUmuyVcSHqVVQv+pPWYaDv/ki3keTQfkk/zB5C7KXFjCT75
jszEjfZQWj9gUwMj4Lgv+JAHPxM0n0KQtlAoPSh/s+LOkDlyqpTrSFStkiVV
LW2m1m/0OhdxfrivWhCqd+ccg5SAmoD7v8Dqvva7TYqSxW5sS/0oUbrTRiJ/
zcYXYGtU+eSchRzSepi9s9Ng4dH0s+vQinLrI1eWBNG2L/98qvLoO7djQHwO
fQefQVUCeRqQwsK38ZexwDvFwXD71znMylNAAHP9B9fx3kSIvPwuj1JA/E6Z
59RKdEwVVO43FxXFCSl5Bd9mt/Mm0WQMxA9azrY4X56cGoIOCQ5t/9y9q+Qf
BIe6WV2aGnTvK+ptWbJlmym8auMNLpHE4jHtgd/Fx3YIkVWK01wkP/v8RtXy
w+zWilD3IfPDl5SOyOlIUa+rZ/yrqNgo1Ob3DkwbEMPaH8MTekpjCsCh2oVZ
x6/0P43il2OBsCyUQqydP5LmUIqYCROk47DPKmJxhWzO1k6PUCoFUG8jPiW0
wl3sKJqFp9e2kxZNzAry37XRiNhqc8iZ3eOlsBqgc+cn/lai+1sJXWVJoXM8
U4qxkkljnGFklKJenbn7Gt4EJFI6/QoOvnQQlT7dU28qSZcHQRmSOOY2UhJp
tRvAl9QYpv7bSfC9SsIgaCpAsFFPCfnq6dFHMbf9jgzACdbt/0Y//Z7p2D8o
jIFQqSfHifNlb/uzQ4oo1cLNArM5FGxyG7+BXdkUG9gv8mvO6MXj/AfAc1w8
4Q/9N/55Ga8APs5AMYyJL8jC1vFIrxrWa9gmYIQKoMlECRcToAjEMQ96ggRH
v+w8do0h5cmqHDOAOYvFnnHVg9KAcAENlSsb0g+Y8SRluIWWtKUIxJYasVb+
WndHtOOIrP00Mfpub4SOeAUiX55wzHQtFVo3ULmNooDF2c9asjbf/ehtcZlr
Ht9ghtK7O6NvW5EVOog7S3UAMQZshkdlQwgNuJWoz35cmumCUbEmMjj9MnJV
OLost+1k3g15XCsf02TaDG0QnUJBa1qyRLzN6rbpt7amriPxr6EhX5uG4XGw
DfXjEH0FX/AIwUKNvfc2HXjZA+PRby23i7YYfXlKjkK/4Rf+EB0rOMylvg45
9mp3aQtmuuukuJS32mAlz8jdz+w0W+8wFSc/ItZjm8uywY9CSPmvgd0rWJc8
Cfz7C1SLtR6Hs6ifB6M4EmeaOkQ3Qxh+1sAdP0/onWcNpD4EGmnY9g6Dv5MQ
/1+bm+ALd3Its0eSkp0s6podwn55Q6c/EWgeqX6rW1mwBbpfI4sRi5BzEQwN
jwBvhFlsYN9CkVaCPvuFzOwpF386AHTMk3drmws7RhRWl0EyipU+yimtjvap
eONRoAmFJ4UtML12m85lgB4IY9DwTFGKot7RoGv4RId14Dnf2YbOZZg50oJH
rR25wxLjAqKpQIhLXEhaaBM61gF+24cibxnGKOR/O466JjVLNseCpy9K6gyh
Wf30EJxbq5t4JW2uNW3WdPVWOiEDZUrC7MfP1ICovvqOEkBndfLbOFRNFkZg
UEAqtNgD1Xg0j9DM8D7jTEh65SV7P5FArLKz5F6TMJxDGgu7bod5KVf3jrPV
kFSEBSXj4u/svhR8DkUC7lD0pOy+Q8YT+HVfooZY75EqerdFJLoTwXUESXIC
UeJnm5TVDLTQcEMclHzwJwjVfpEyMszr71fp1Ms9yfrCnT65V3M/Ta7koH4P
LfnheEYquwI3UV5Zv0IpUxtPC0DQeAPA29bZsBnbyYcH6Lo52q9huLMMqv2K
jT1OwjRQ/kqbuhjlQpPe86/hZHtgf/JviGOX9RXiZu9syoQhZts+5BApj1/L
jreppNSjK4wq3tsbC6RwKx8n4F3MBE0aPl0JIeEwfi99qfaaVMd7DyxcQXh+
J7j+fhKb8ZGjzZogUxBj9IqQz4VeqzJSkqA6bHf04dF9L7987nEoyeIyOGof
GWNLXLhUDHKoAe0H8Tn8Z/IZPUUk0MOxCIewv10lbO+GO9No7tL8Aypzu/gT
SWgXkVA4BaYXSCvtTEhQTtIL7qOUDLK2r34mKvDw6sUIUNRxaNh/Hc/EZ7E6
908iMawhTxzgNF7RF70wj64QF9/iIaFsriLCKpUUuwaw+Psxgx5N8uT0jJzU
VV2pkJC/OGOOkeKnQ72j37Az7UiFCWk9g1Ph+GvjfHJZaH+BhqiK8pFwSm86
NZZkTpri4XFNrwVs/9vec583vaICNMG8b+xdBpGnD/bHG24l4PgcYB6S8Cw3
kp89jg/H/qdfo0CizknFBjwRLJuhmELl8K1pGWhqDFERb3AVo3gsnDHoJ/AE
7FSxPw854q0q7lPXvmmauVH1TFxXYdYn4qCQTqlAuruNSbPo0zd4xznCv0G1
E1R23vqtIgJM8NkGtoOPszQ1WaOZRr4fJ4i3gg7UM81ATKJZn8wQ7S70tbJt
WzweNO4GPT1zuJrVNPx27FHDxeBSfUPWJc16fAAAuOtYnwiwHVSzQc2OZQzy
jPtHGvM39Cjd/nuURfyAalsnselcmekZNo7hGhudkWwAbu3LkwqbzgsQjyzM
OXSKOPPaOeBgwz9r3TzZeODnMpC4RsZs0auz9mqxTstN0hFkBRO8ylb/37ck
kIUKmq8f7F6+ssiYQmQ2RniO6R5eY9UhlEJ+PYq2F5XI77cEFnu+QeiP5pqA
Swn1oHucDgcw5FkhIwIEydkPUvVs14d9BSotv2PMhNELBasvnUWc605qXgwf
OOlmcAdwDw+pqXhltt1+l9ZpTEczEDYmpZPvUJJPHTvlElFx9jr/6moxIJ+O
1ckCXHNZWJgASJmSVAL+lkkDHDDYl9rCBCkDeDf6kI/xsX8iFOD2ZANwY0f/
3GAr4P8XAMHHf0sYGoyHE2gl5XwPpoi7tGF7+LA+DN7XQ2Crg0tsK7mWk0Pu
kTwCIPX8ijjrcHMo+4aggFC5zVfyvhKuqMRO83A43J0ORLG+3OxpCKS9nJ44
QVrmY9ejzi4dOpJ6O9yTp7rEGzAxZbl/7ErGfOdoiAmFD3CXxgd27vHr7A15
jzpWRoisuE+QpOrcXl/1MrhqNEgc9InAWm6vgW5e7gtOUXooy1hCtLJMOfrL
yhqecYS7LYvvMGs+nSSZviX3A1Gz1AVphx2/VNP4lJworlvz3+h09WmELcQv
QFzFjJwGzlzv4Ln3/HY3tpFA2eA3TcG3EbNOTkwllHQ3jqjUSXNgUhl2THt+
wHP90sgGUDEpj5w/dHxXJ+NNU9DHF2q3v/RximA8Av7U/0xg6yyDZiU0s2EM
z4Ae6EztH0OjfVKtNtqSGrWV1kJ5lrvga3UHZWDdwEUmYcrvRidQU+3cQfPP
eAROIrWCE7nb6Sur++7tkVyzG9ARkv5EstlxfPFQbcLwn6CJENB9v6JYWE+f
ZXmJkg+MkyAXF8ApQWfriNNQRUMZF7CO/yEK+WO+bpe9QkbcvNCwDGkmG+oQ
0gJXR8dnfyOW50+/WCBu9K/nDRY3r8fGdOuBbij8UTUlxFM4qUo9C9/VY1VI
xLqlQW8ZfXph1PnM0JzG9qS0Oj/dKfEriBDVbbL6fpCWKV4NGxZBnr6qXmX0
2xb8TqVZovN0lIj5XAReUYxBL7uQw+cq+MOsjhnyNnctJliC9hfyGndlglfw
RKG4hh5JenjVrnHaX3laVgWDssVwouSY3eTZdDgNJOBw2xkqs1QqnGOcf3xR
QRLCE271OIytgBuntS8EzA1Hlx9Wpbbfiut74AiA+lwZpOXCPYh70BjQO1ED
lMPMTH2xuQ/Csi6P+3YmAWybRxCg/4bfl9WWOdIk1ZOuQYrLub0/w2T4peWt
QrGpGDAzFJOOjebzospTQECdoLN5FCzCI1kkQq0MAB3bI0DrJB25dxnhiBD0
zQvvRKjJCuOX7LOe7OoyxnkKVmEjNM4cgRv7CQPYcO4wLSWQjvcdqubfIykV
k8v2BJzio8ZP2ZNz+/uv2TRGmAMmNBCQEuR4szLgLhCNHNd3pS8+/GF+rwBe
y/FR/trQianusYMkLdn0L2b14UquNnlERVjk1Zrcz7PuJCxk0iaK8Q5PbVLh
nDL6S1N8ZGiBXsqpiEVJIngD0wZY7IDl2t5Q69lAEQW40JmMdR5NBfUhzFUK
XT8x2Djac5s87nz4JAjxFR7JN221s7WaxAp3WU3yzDIF7ggXOb9+B0uaDfqW
OemNeC/i+m0wG+wZqlrz0BjZA+6rPoPCsLkI2lQOjgwNhPIYpx22DPvptn0h
OLI3JRWKFwD3Kd6M/vRtdLfsxKf2Hx/JMKQFGATMfqJXLauftud+ccqrviR0
JKxOkjM5/sbZGNsRCuDvmmmn0VK2RCC1sv7/LTxSH0yJGXIs+dwqIN0N53K4
s9/K9CkJTLRYW4qBVgj/JxapwV973n6+0TbS2lUPpegKDYuSwp/ecjpjtT9L
Bya32uDpMGxyxkyi1bT/NrmFoDsHa2DnG6psKMUPW0kZGb72eGoHl5n8IEFU
wf8pv1f3f2w8zyNQhDEmmQH5Yrus+8J8NusL15yzfl87/ef5vU2J0OPsWFm+
fUfTlVdHqTbcvk93RtGu2fm2ZCOsAe6mqwa8tQWW+83a/Zz89T/2swogixqP
T2sRLZfrzkfPAv/Pb7jRF+kvCZREi20IG7eaHxLZj6esJ2c4ymZA3iGEXnMx
FnpgomLo62t4/jSJj+Ec2UhkGccxb/njh1Wr59Il/H2yp1AKI3lqpCanCHvy
Abmw3xYgTX8BISIrIN3QCtrr63ZdR2aUqQ9DUHytgyLdAKblFQsQ4IQ2kIEi
CYkoB5JpaxLtzwvGHV+/DmaDoypmJpvAZp70j2IHcUFNXZNYL7visf3pSJM+
aOD63eW4ah9upZ9SDu0qfrjkLBeWYJrP8TtUzwjdhHKwhQ9DkC6C0wBaYiWn
3fc5eluxNtq881RW8I423StIBVMqqDxT3Ytz1f5OYhgUMHaBipy4cB5fdegK
WUQj9JbLGoJYoljPQJeuh3r9G1QStuMPvOE2hUCvcyA3ZLAKVrYSnq1vir/Z
89WKF+hXr3ShLRTjyyIaIrFMSvyJFZYtlVuNYmia+5YBaEEB8pVqsQQ4t1vI
xcanmbEn71RGbJdN6zqcW1VW0rBa9QPhtzTUM07ULUTUYAwW4ajiqrgAVEh6
oiLGmchhYteU4wPxLCEZ5tBdI4Y8k1cHpGMQJ35y0JEY/GTkXfQ1/te9bIN8
wPqeAVKr18+Fvvi8p6IgRkQsy46PDHTRuyrMGlgy3X8tUDByN4bGXT+W/bdd
+QC4xJAjrvyy4+8tLSiBgyly4LCxxyl/X7xHCNFIpHLhfUJsdqe3rqE1fy0h
zhim9tsdz+jkFd0cK6c3eR33SWprc2/Rf5uUEogafE6IxWV5B/d+q7FGMyyR
Tl8BOaEnf570FgoNHGCSjEyv+C0x5gJo1T59HNJPIlZ+40Y2zY4EDoO17nxg
b2xO1ZAlmXIs6yQ6NerL+tcgXxpVEPqEhOknJfcs85Hs9gQJFJTmUah5ls+R
Xdfgi93IO/P7JmCJFUexyobeKA/cGtxvh5eLg0DANhDL8rvjK1Q89jmC+e8Q
EBudnI2N78vwm3EhI7GSB28Srx64yLf5QFR0SEDUAnVHA3ZRZ1mcr+NWEcAA
BF+9cxt236YqePtkTOyPIjTh0gmgFqN7vTV/+HnQuZOd0rX7XpHVhKyCpCz+
uwlLU37WJnG4RtWbM4ZkfqhgnDSyGqoglL+1X3u2ClDeTsY0QGVwCxQUTRKY
8c6ioFlaolDOpzpILQdwR4IEEaL5gJkDtEzVkcW+1knFBJJj1/J2G5CHQa/L
RVqr/5ZVwlsw2LW7A+lEpdczBoRtH6BtZJYcDw4lIz2rY++ZkhYId8vau8u5
g9FK5n/A+F2ls9T5oOEBFDCSLqgMDv6LzNw/a0yraoqdgFTzNjkr+Xq8QE4A
HerSgSXIOJpV4Wewvg0wBy7DIfF9Xc4Zz1FtQ1/Nydg87TDT5er8r7cSKF5d
M0Ya1qvpzqdJA/yje1y4dlGGT753D3CEtBr6KCCN7Ne9DflIHOe1XN02Stw8
OlLrNBFxTagI3wBNQvH2BSlxfpsRgTngs3G07E2X2f97KY3xZt3dA7leGgXR
4431HdbpgFjHK8cgIOXOiC/T5BylijoM0CRH4xhZgTLtApI/hQFGjR0RzWXe
2MsctzPPfaVpOLnw1hOggDvs4jD528i256rPUEc2FJ2T/XHcglb+xYhNtn2j
D6LHGhcFr+zNZndePpFOPdXRUTje4Yarz66m+M9rDbVumJxaQxNn4SkEXSoH
Q9llVXX13hTyiFRXGXSJco/MNwowOeWMXiJMEbjb4pWViR7YKAVdyheLL3/m
p2CpXWzn2uUXtVhk+hcope1KCoMHJpnVUHloWzVxb54aJlW8LV/gbanmTi65
EWKfnRBqtHglyuqFHQ5ogVkQcuvb9pzvm0f37/m4feDZuHyUW3uVSKPt3SUz
MrB8MpOGHwNhk62s9cFapV+kFcZXzndD+IcmYXCs3hd1Ojk/R3Hsg7HISEmK
e2x4lP6vbbqGd6vvc9nFQna4jlCFzpamFTQ31ga9/l+uUAN++jcQsHwTA+am
KdufXsDr2EIGlpswZZ+K35rxIbTAopVUMhjtmU6UoXgYjw9EhokwxGHcSvyh
y59uxFEyQhScAPJ9HNO0NZSMctc+c4Mla0JAkc7iwlODgfyc6pi5TbEJmTsB
boyij0SUF8hS8btb3gTriVEOJzImwHaF8MckWgEeLYSq8UFkBKzl4I8efv89
188LPMzgzZP03VzLRzPGLJiEOTclgfYTHrSXOUoxOAvDzeeiIWNrLdnowEaY
gwmLGERJ6YrnGkb9AnQ6Clf1e8bt9WcqICgTW95TW3gX//Wf1AAbheemcaRs
j0iKj2JY+vqpkoZHXPdpWWq7w1Kzix0amc3d3nemrBdA1sd9Gdze9Zu+N3BW
FmV7k0CA780ZikLEW0NymdJNFexFQ8d+vbDA4VxoApyRo4OUs87erKyR2gxj
b+DASA9AJL4pnox3gR0piM+HRYuQkVuwhuOhZMycgwx3xnCYWCmcXmNOP+9y
Q3A7ilc0RnE43npr+YvIGLwTceVlxyhQr68wfdQhNOJVwGoCaB+NbSPDHPbL
AGQVDW5V200+4KI0SwcbiDkwk4fNQUDji54KBm5ztm29kEcG1uok/Q6yq5n/
x7jeYuC2+IBAN+LvGkhQLvNj6OXJboCj5xqAmbf8S5/M4FC011OyaZ4BkrGI
uhejyj4SefsShJCpURJTmxIK5WXgjN7kQ/4lTerNsVIjuyMQxz2Kh0BF9Q8K
bXHafWDHUKbPQk4UntyH/tpqKeogc+o84cXYDneK5kVGuRF25xL1Bmr39CAh
oxig8Kr76KaaUl2kO9WRHGC9EztmvIbP7K6j7sZiO5knfwX9sGV+/DnLRg/L
Rejf+RMLHW9G+nhp+YEiXVfxXzvsXyhPFnpa+ksOvH70Pp4uRhV5Z8II7tF6
SQa8QTao2bH4pplwZ4bLiMQtAwXoLxKRjwHt2H2zE4oAqbZGJepVtfu7owHJ
EKHT9LhLFsK412tfWkHgaridybQSqipTAnZzKKF+AaYleKmDycoh3AABtXNU
LGS7bMZOvZ/gCR8TnRh4Gayq5opPJLKD02bu3xGw2URNPt2oE7E/n1ImugFS
dpLfLjxjlSX4XrNl/Q7zveE+IrRt8UnM5+qu9/Ih5KTUglzc/7RX7PRvxljZ
fsIBV/dPPgD8KNhcci5W2n35zlA4HjCAbwgXlXQr55+gP4Uk/H+eOKBwu3+e
4GmOD071XJQaM4eq9nfVDBNFlxa88DKUiaUDH9RZBvVB/PoK+vPdBTuj2WZh
I++SRN5O81L5UbuqLP8Rp5+zw27cbIsrJgMHS/EjEdRFMkM8veDjAyo3f7IM
oWR2yK+nhLncUfdjPx9ul3S+Fd0qoG2KNqu61DQjSYRm3kr0bWlZqGewhJkf
VjRCuwHTIW1ocj/eEEiQr/WbYp8mTAlTotpx6odFS8+kwxpvCg5oXVK/jpxQ
RhH9utrGJNLHxLVjCrpLPjjovYf+PVY6C8qrH0F9/gIT0Hv+0lOKa8+LQK6T
X74s7s6xrK2WVO+bgAGuGQaXAypbdbPs2nxxgVgkGyS5uINETyoxJcPu+WE2
elyhTuCxk3yAWomGidrSO8WORaeX9t7MnGj2S2RHP6rNH1d7cJVJ8JtaKk0r
rmHautibvqpVQR8bMQw74maApZdBCNg84ONibIihR0Oeat00eWDqRPJT3GU9
BNliex72DqNPki4Xt2ovR3l8bUO3/qHyBtz4dtzuBk+ensE8MXDzXHtXZ9v9
PRajAfsBk0H+bHrW5El35JcNw9kvv3wkHo3fM7gVQdDizNvKKhCobwYAhay1
9bswtZEHhVzC6EBA+SYw91/G2uCy1VYgMfFnC/g6BWTikAi6lYqW8mE9lPLB
J6jpz7fgHjORBQNqVb7Cbha+z6hPdXhj5OWUSq1zvU2vtqXcP694tOnqTthF
N885ZeaEE2VfmjL4d/CX6hwiqfi0nu3nGg8MNrIz0TVINJp9MmNQrRqxcrQ1
ftTz5bDbk9j+GBBklNyA4cRvvkW1C3JU/utVcgfQ4ESFwj9jwO/BzAJcJthG
NMzlMeheTze9l4gvAPYYXYaJ4xjcR0r5px0UlM3R57mJt7i9B44GsURe2DUx
k8GaZtsoVLB7JCtC0oVL1jUi6klrnq5yHmhPyRMMd05JIdReqeZs1JQNxbUS
QHtLXKp6I8L7cQDWbUkrxJjMzvgaB0IEMOKVdKjsd7R8nrwHUE4Q0af5110k
R/e1FS4HU3Wl56Y8KVs+N9bbugv5mqduB0HYcf5akQJoBiFTs3ZdiQ96Nwwg
IxDkCQPMmDFBYPyCeILJEh7viBjyJPNDTIVVwH3e7XTxVggI0+z04KMZdEhJ
68Jn373Fxa9YMxpdXlFpQ+R/EiK4M24B8L6Rz3BW+ZX5V0knfsWLfLP/S8k7
8lCNK/Je9HcslfOOduWhP/2Xed9kddpIY6YVpxs9b37rnQpL9nIQK1vjM8Pz
xoamjZu/HylRJiLhUmqjXZknPe5nYUSB68BGodFabey5RYyAUI1/QO1ap1hF
/Lh1QQne+i4UPePyRu1JlZQxJqs+svTmFfDEPp2vuFF49HJ5k9lwVcZacw1z
/ydggY8YprJszKOfVysYiH6mXgrc7Yhxy+0MfLDalF21ZONZhpar4BUwnguu
JsRZ87xv6l9m0Acuz4OOiv/fVFMqdhNo2LhiFjRkiCPHxnUxilhnNPDkxEyN
I30I3Gd6DXx/FfvF2+Ccfu623J7NSrT31qc8wAx98tcFIxt2l6yN1s0Up3At
Y/ryJztb8jJbnOZ52HhLXuaNL/F2UvkHLescJ3Lhe0vfpVporIIaCCC3kcsR
IBtGG253Blg6r8Z24PmDiwpKvPBzSRe9Mq9Had7JgTzSywXtScZ7FffLkkpx
wJkHYd5OOZnADBOjNjiJ/RzJTZVQ51I4zLvqIc5nWwsGedcA5s/0KDvZ6VSH
hSRlFU3lRnkS9jBHO3636/jwd4lU5xtUrXG5OOgRRGAD03vj2dxs/N+3RlmD
+MOomzz4xkd8nWPBrRBYpchlWg0QYlx6TE+7XAAU9LAcF6dEjzFaVQIIbwAd
+bMMBJi5zP+i9epfdN4brcwmUNkbhuGC34nC0SqBUCcEzLGMkevp9sbeQPfO
q7A+9Z4dmIaM7RzyiepVKilCr9zB5XH+bII9mjsg2kQiRr/KVNC8jAtsC5MY
DR9njHbkJzBbFXnut5XGRKK4tNl3QAVYar2LeUTXnw6A8w6VOk+6doPGzZJ3
e7XWMp/gKBn2cMfMehaiq6PQAOS5Z1Owzc/xUfAloxrqucr6c7L+MTC6AFBW
6gJ4eaU3afFpzwGCLA/Q4KRpXMI9NtWLxpSVgI/MwbtnMNPlTSH8/AoLfgFk
L6zl1RUrGFbQZ0ISzVd7KH2TW3QshYuclk54wcuDRl4LT8WDTYTrazf1KGsW
u/eXZpCP0dYXjSVBjBro9G+MCdS+/p7qJghSpggv27RiUcJjuQSlAM5y/YiE
c0ViPl3WeyjyIac3LGfQzSn6FclNV9yiVxhK+jhYTpT+l+RkBM+3/AKugDbm
qYTRaoqxGj33Mqpbd25vO48rBxaVBgreKp7B8LX3fXs1Jo/Wvqd+ygOU5pAW
b8WIFhjb22X/x7xngsjSKuV2aNGVkuGddnaPDwKiyNLsp3HJHFhtdwVZzWOd
ngjCG8lgGqFnpjNEt0iNudgXU77Ga4KtTF+nWnnJNwoMB98WjV1Sd5v+78jL
GLX5YPKzcds3tgpd2uVsTi2gylXbxU/NupnheS0ujFGh3/5KsAoB4IPqq0GI
Q3a89KDH+uLOpb85gfpor+oESafy3lLTuNb8sKg8hanGe4rukY53R9KT1j70
oYiTuKzvWEuIDABqmIwIbgIacy3CXklA8zdCm45IsuSLJ+1s50zEQBsaDcS0
tdvnbfbFcYrwMLD8wyKCMMdkHxd0t8q/y4BGfJ9BHj4qvXC4dgMmlJoNbsqf
FE15UZW1xsbrv1YLtlhtAxMQ0QJG2xstlQhJfh+sHOlTKnKbco/9FEwv+Si/
SXMXV1ULSquL9xiavOkoVCXPGzhX4v1+SUmboXz20rMY/4VE2YHqlUiEAXWv
IrlLchDZRPr6bFuRcJl+3lfNZ0wTxvcPZO9bpkoX1B7LXMkbCmj23CpT8soR
OgDIlAXMqqLfW4yZxzFhhwfM+AuZEKpPV+24tXzSUh6EXlIbMCSYZnOkG7aN
WjVr4Y+nsGj8jcvLvqYgdbgbFURYe4I83/Pw7RrcIWMNGTM9ga+xfNMNooLl
gd8Ljgu6eMC3Jy3x1aFTfXz2l/VaZ7TVymelR0OmJlHVfu6q1/7al2QKLbfc
14WJXbkSRj+kGOQgGkf8eIH7WF9M1jhad+GBFNp30X5O85vqXq22eMsWeUJc
VmRlPJyQ0TqtRXgZdqb04xtSSuPDDA02+k86VnEUmcf96l0JGmX6N1E5CTYq
vekmP+gSCUD8rDD2Z0ag3pyP/jZZfDeBs8z2cnEpirlD9VVYcOiel4Ci7nDm
SdqYup1gU51tQ6m2Pt64nk/qxdhnYf28DvL9TXMBPyBi6Jywiyqe0h3/zLqy
pjhkVhOfA8fgpCCnnyhtLBdmJlzCnxN3d6yir1U7Bd7b8fSsoDURp7f6mvkn
k4qaLlqTCzyA9b0wooxSoMPMIk8udK2TX8TQtkyDTMG9UBoZkA6vihFWP5R7
D4E3Hf4d0YFyrk0dg0Zmr8r5TD9h9FH64KZ2RdGr3L6XJ8Wa78Rv90AnJty9
CBoFbu8tHLjcNq/M4vU3naDnDNJe9v61mLYlaqfvC9i90EkKqbyobqpV04b7
WyCxXb/g/4IPysNDHA7QD1jFsT18iLEemn52rB8fP6RpBqgwOVfXBRC47xXy
tYmPcZGIdZwFJYTQaVY2iMVWh72LTRsE1sCD4I9bWtSQOWKsx3kqHoSSXGUy
0CG7iAWAQ10h8tQq0k9JEYJL+sU219TQX2dLsp9tbHdu8OT05RThcRVP6zf6
d8lpqH5Gg1JIUdMOOwXjCfihyEx0oivMu35epiPpBdxoPcF9IXlb6Hk+BrHD
ukjMUEkcxJRWAtlX62nFmFtGACwIXHljuescv3uH8hsgBlinw/6wvxGVVfTm
WSptUWVValjvPdxUFVj4H/gjBaTA+QSie83uNUkCfwipzQt6IX2Mc5HpBiU8
+oD46XN+FOuKwao5WGCYajUaGW8FFA8P9hOCyUpgoIkjraO6uAV6ZnIqCZN/
3jnGd1ZZtAgnTWdjd8rJYPYjnjEYXHI23JSTjriVywvsC/5eiFyzFGCdAWSi
TAX1sNgFYK/IGypDfGyDTfURkbt7E1j5Vq24TAbRvwFoUOHpTelYL4pSRI1a
vPVeS2Yh1H+ZwaXMtZDvXWTq/5ZCsKu2Z8cMa34XU5C5TkM5fQgKja1VOgon
yNHn2hFLaM3lFVC8f1KqHL7vQ26t3MCQaLleYlr7ZLhA/zKXimo7gYhXA53r
/nchPWUuDcAUs9UrSNlgCadqkWW1iH7ijaW1aBIoTYJLEI69fq8+9jRJSRJS
3iM7haLBQnQXYiurG0zQiXIBhXfkElD59ggsvvNfYSaYlUvKNVZTgpiJgpPJ
7uOV8dlmGhV+Z/6qEEEo10QqbJzaMTcEfvw3qj5toHyiiV3vVPcU+4luM+Ej
jKQZfO+z52fY/dZixunl8xzpH3RkLU6xHfgNDcD+a5kK6GHOdIWZm4e5Do55
k9g6PHCfBUo2mDLxwIn7F8IEgpi5xo6gYJhCbsYTsRSDmuruosDy7A+aBcW6
3hXYRCJMZBZFYvkhBAv/p86pIUuKXmXlu/sHDbahLIXSE1upMR7LO6hvoWwH
4X3oR4BvTSxFKsA4aFBxTSSU5Se1fpTCchZPNMUbiQpYIcHgFjl3d17ZBpUW
vz5txkBBDvP/B9ckAe+JJSF5XYluggf7mR5jmUp9Z1bymVcqn0U2f1oaBzMg
jZoW2SMQisjF7IIV9Tvahgx+YpeQh5VHHEbVKjRvJjDeOGbJwgjK/RQWuhf9
mp9RR8ru1fNdyMogOKE4JAhTOzZkhj3sF1PbuxbbJuXKGLowLUWXSEVR7iEh
qX4vIL0pkRvweioVdgiTEHvnhQnMRTpt/LDm1RiBJUNR+0iRcnDUXDi7Nira
TVcpS8GIjUdBZAUc0144N9lbiLRZwQEXVXKdFgmZ7kjg6bu+9+pmYWyQeUx2
q4b0efN6JTNdVX57b9oum0QdcTteNQkv2q1PQPJLC6XyfvQMTQJPD3L7BgGo
LQ8HRiSfCDwyYfJr1v2c/3Wf9wtEq5/2H/LNkEUtrMvyTDBRCRNVbEUVzEZc
9/+/jj6ocEX9xTLS6zVlww0dUFQLhekU0i5SoPDaJScAZZhRbk9lEUEq5rEm
oxb0PeCKI4h56tkAHGYogKg8qRtvw4b1tYHkGnBV5wZoLg85wup2lEzfvnt8
01+C0VtGxWV2lm7JKw9B2lA2Sc2dyAg70jvVwGaEftbWEoQIAIT4lMLrkzEE
hCIlVVbMhvXeOIvJ1qJmcJi1RTSnwk2DCRoqVtEh5jssh5Z3DxSNaT0bpJET
k5y0zEH5nIRIaAT2EHKfpd5BzZA7Qhd4bbIodWRctpCxsLs0k6e8W63uB7QD
SsnFC+4drXNFr+zDnjh2gtlUXccSNkHte3cwwTQ7SlhedBr9tsjbfXIkzugr
OKOijmzpErtte+DNsePamDwFSNsbWkoBnx17ScKmMhjVPOBiLCBAb+kbrVyi
6yO2jlfX4s96YrIB++TmWcPr2vnkygAxlkfxkU9KQd5oJ0KteU83YkCjGbG5
aOEEebhxTdsMiOPtIe/0O2ox/JDq2kxUpOfZhEluny80UjmGfUU84mgRrphW
Zcq7mNTL8Vzfh8KGvZFvQgKG8IhD+5LlokzTX+e0NRRg2RWNyguTEoZQ6yFO
zH5xJf6Yvbi6f8tmtQqvB27nFeyQBlvo+DYWo2IXIfbFsgY3Ue/ngzYIh1QL
g78y9DBo4aG/6Pt4NUbvKL0Xo33sGavKh9QmIDDWDZ6+eJOXbKGkw1U5gmaK
Alb/8B7CpmMoWQrh4rd1JxJAw04vIXisOkVeYoDrI0rY3cmsji4IOnh3F3OJ
LA3FyCOsjHcmWARbTlTm85IM0aFdUzUENyj8wK72OZ/SkNBya+YcXPlK7Okn
nlEWrda86kp1kzIfwqL6sYuV46adN9p3el9WmU/O8HJuza7yvZlBGNTLl2TI
Y0mjzwMPBgN//KJKZFYrlhNoNMC2hOxisaFsh/4zjHzwSa/mttV+5od3YbzR
yYFdlfsE2R3buTmex43NUuFiBwoJe6xj8yEnKFhFGedbB/nzEIDUwpC2QPco
nctxh8eSkYM2T3gYJoI+bYSsP6LjtPMELpwFwNxUJeW1ymWLZuSJLJ2vCO/s
1S9ucXACPdcKYRRvL7HGYEkKXuAi5ouefBptfQMEsQ+Pk8xCC0v0i0D6MMac
PpuGrChXaXDxBSKcO0CctXv0eDayl6O5VXPbdCB66+WOe/DdlQ6E8/oozCIL
8LYCPr2fmIM+7E/ppBP4Riay+HHgVXxVMJ4Rk6lkp6saDIomfmPvPRDbO6+l
wtOaDL2wRlcgUVWHfvY98950TSl4mJQLB3zc66UioHbXKL7jg294wa7lYsJe
lrH7SVHFJb1Du3yanOGDaBdFpUiNn5DVNAvSJiMFMstf3UinXJkwOOtiLwjw
93OdJcGVfLMunlx6s/0IBGKuiM9c3bKRMsdq/KlO2tR/M5ppVXBUHJnNzBEG
toPH0AoZpuWTU/pKZxIW58qDSv6KG0Sdj38eU/YlwPKRFT8f0hu8rXNzSOFR
GehLswzf0/VUBKstcboDAQvuBa+cJV6uWq7QJ1qvJzj2f87Kq0MNklbbcsd+
tiPJl3CKmNnvVWRJ0jFaJOBbUCJaWG+HuGiX6gfdN45RmEIwTl13JKaQjZco
mboLqRnOTpRSOW18Nxd9C43eLc8ljM/c6QgZ1e3OKLxf4H/LsnSnj8EMnkoD
YsyvyjUYmwS/BbTldkuIaBZbuGK3iMWc15niTz2UNRteAPH5btQSoi8Y+rgz
zddWKnBWqF25iwIizwA9PbB+zXBDXytshgdlv7GVni5FcxsAaQ4Zvl+tn1ad
aZtoPo0MeMnY1vv7XJBZJkG5YKQCs2YhdiwYuuTpbK3RW4T03f6x1NA4Okty
DibOf2EQK/0KVrBTA9k3kJiGSz2WjLS0cGhZD55uCdM8PC5IOEAo0EKVI5PV
+rV1cA+vMtewtnOxvy8UY+pqWl2Tb6kCHqIJixcakLrjg04c1nxXXLAuDKdb
CVilBinIna1XpxwKKWyALcazC5ei5fnoSXW3luD1bFNRQLd1XLfg+ZtWvtSn
nkjc/iDPW4GcZURZwYQmwoQzwaD15CojymunBGi1ZLccAUdkiZdAlQcAnrhJ
C+exZTIdjeO4nFcqdroEdllRAbE7BfT2rO4dU6dNuB4BoGDno0DhT/Mbw37k
frO8luB4lYF5XDubWcsMKzJuwV6BWHTmAdMmVwEa4qNufWQJDyawmU+nbEUr
u5ADzRznuWuqA4lIZX7fJUlAdvvFvTQYRcXulAyVNTGlrQC8dMvKraSG71/G
Ku/Xf2WTMjrx8In9WQpkSiDpLgpMUxTLcEhfH8DFq1oKqZ5s5mJaoxcwRxD3
yUSqhaj57TbxMXGFJmSFlOqp0jsb3KSOjn9HnOWEeXTrHgswqmDzpadr1lsx
9Ewymry0k+fGkzI8DqWHm/bPP7ELAXTsbyHkNozvPDz77Q6HkHea31jCNHOH
ecCz2hr5Pw7BZ0GosCmsKWbiSTXIMLKH6DXoQILejCzzNWBZR917gOtA625P
hN57BnQYKFbxHnfgY6BM3/1ESNTY83A5hocAQ4zZjwznJ37l97DgOLRdU9uU
snophEfdQOCn8JomDwIFG2sM7lxlaVulNSm2lTlpNIlCg32Fmo5ncPIhmooV
MK/laKXXhF5JkVR/ujCww5VLQN3lzMA+JVNe89l0AZR/lcbUfkEnze+SMyP+
4wGR2b0iWvzfa7vJ1KiOl79rBvPlbVRKyWvQNuPTi4TVeas0XhOcmICcsT0A
Z7stB3D/638Ce2bQnCVsUZT10HeULzoZybGJrqRIkBzLoxgnrOJ3ufaSNgNQ
r2T/87uRw+YN1WB/LBCXozEPJX+IuDB7hQgB8Y4K9u1LYByJLQyo2kfCIbTH
o7yAAXqU90CFypWrn/1O9GIoBk7BHJHDCulI+xNL1yT6oGUXosXNLGbEURvz
GblZyVPg3RzG9vycMv8xo2laVPz2nEtO31+AwxZO2yTV+Yqe5/tMfparjtqr
kLQzIcHDs5s3vysoYb88/PGDzMn01IRKftG0aaOcVpQOENG6GZUxT7H9Tl5L
VxdPNX2OUThaWdQaZMFoTlX73Dygrekzz5Td+/RjDSlNV/hPmm7GDmFyecB7
fUcED6xlsTOQ4NFYYfBDMWHDn3dbogcsWD7EtNX/fufTztIJhHJbl+ScSGga
0RkNIdAsY4tB0CJWgse/aRgSF1h7E50nDWtsQvmgla1+YWe9+9C5lX6DGcqU
7+NoxZ5CjOs97R9tBrrYmPJE7Uklt9OhpY4zM0FKAwOYjScWFP7Tk/MqjkVk
1dJHYooIy/oxUA8ThF1dWZvvtUR4P8N0tPg/vaOhpFYHInP8+b2vwPHjrUmX
Awe/PsDbjCgHMBDsil1gVgEs744FL6S6aEEczsdAB8TtNKLh88sx+CFQWgTV
LHPSHkCVSC27fS7KtxIOtX9oVlUEXtuWXm01uCVVfBQy7We3dffPFkzpHXo3
aPI+aiAVTZyVOb6IGoDUWvTrGzwDaau4UtoJQ2Hw0FdQQDJttfZMgDkDUK+b
gzz7xjf9ElusudQySfM6Ufin/ZorV/MZIGctIVcCOAjOc8Na2AL1PBzH7cIa
I+NF79D5rdbZP6CrRBCm7PXvd96UVWIAcLUQO2Qp3HtbY9sO1uFVlND3l+4A
nDEdPdFc3DxAz7/KbZtotNYX2cqq8kJIAQHkMCsR3cdm8l7ivv3p7Fn17sjq
lBQYvwjfYLgr53uLDzDqheSIqSSPlzs7+ExYhYjhGaRaWVHs5FGA7LsjaVrT
uGKSgrez9Qaay2h9qTYb3elCvQu0Knq56uvhOYyNVvxGNTKlwkQS2HLQRzpu
2yKSDK6X588hstswqmDkwr9Z+1ADkEzFSBef3fhG7GeC8WbNwUlN2mbyRlrM
jP6aOHvqECdLRUuT7uSArIm/V34NL4vLksZWPsehvhkDHtQBTRM2RO3E5Cpu
CobyofuonBX64ZwUWu+kD0jEVhKrWuMvyBf6Q8Sd3xvAQ+EwPtAA04yl8pJ3
4ct8ruHV22zkCaZMIZePgNaIOZdM70o8afxjiMdC97hldwhzqp2X2gHK2IZA
uuJdNfVTzpUEGk2tFEq/82YDQPpXXDGBjC6NGSe02FEOnwIneuGRCwCJOHTV
CxbbrHp84hz9cYDTxfv36DShGHWtf+93AURxtDJ68BhJAmgR47+FjARFYsf3
T+gGihSDzVxvKKQGJpsVufBciyM1i+KyrMjEgwxwpeQJVYmQVkYE9zAG1cTj
zsCbR9eUDYbfzgWFrDN0dEizwYUtVtS7DB3dQh0N5X8IfF1Iaf4wJjWPHR4u
zf3ifZZtqbs9KzSqWlTqdPY8g59TOpUtFrNmfiHRdjpezCTcnmzx5nMUYME9
qSgyMLNhMpZ4ik60LsDw/CP4H9doabf3NRd0i7WZs5R/Dvl+Toi/Y5oUHtcb
DfQco4dhEuJ6aGo3fNI80dc6F+4lDFT0wM/YPD0eRHa3S/ZwanR5XbT9iEd8
3OCrb8iOY59jBM+VY7jtLexeDgll73WpODcfokH6CwoAonGKDO9g7yqS/Zz2
87qPKeWI5qKlmyXR7uVk8k/L1Md3lDYuOSyWvx2YhhrCxCLcYzs/6gG64bmI
IX/CzaKi2gE7b0ZP4CPUuAnTex5YSjDX22RzP9AiprFZ+CVcoNjQmtVC4om1
DekOQNPru0WKoqGglYqUJIxFePGlft0+DVOM/PfN/xiHERmU3iwgQmO3vVgu
2e+e+/XMX2U4m51a/DafsWBq+oCWb5HK9gbINHbM9vw+KXUPvz6b/CzLDDzQ
bAi66NoskmCTE9fF+aRc7iz0ofwAdAOFC1Du79dDIs/NVlWJrWbZVf4eF72d
NbOVNrfurSrhEmbXSkmJDfwboSv9bzSgnzibLKC7tFUD0XYSBllW+ufrgGum
tRcXaEljPso3G4WxesYFCLAcgb72rr5u2O0lV12RpphobtRFWdd+m2YuYv9o
+PS3ncdR46VNbcwcIce2yXT7J7PaxDVDgxZQ74Z60y27xeFFPTvJHY9mlymA
kQgAPDEjq0Ki7rhrQ7YRjNb7geterRroSoQDrrdW67fpnFcdwi3WqDlKRY4A
R9r9lkT40RrIBl6fJ9KjhOe1nFti6nQnzZEYXhOjqGLI6I7bzyu6s9G6K2BG
duxZtGnu5izfLZpKGpQ8Zt6yqPzEqp4HOW+nxTkzRnbWghRQYrtm2qUbGeJy
+JDbrLHR/4XUI4HkVSO3U85zX4G5w5lxH7dJWK/8J224hG4Cr7zqA/8xTn58
D5ywO38BPLMQlttNJMK/9AIw9HTerFLObTUygCuaWRrUFuQmkGD+dQllOWU6
qqONAAGJReXn9Nx+n0eS7TVknKCYbRQoGMfZ+MwwIINoiKpgj1mARD/q52AR
U2uuCHkJ1fxYw4AoQpHgQFXoN45toKuHUpw3ttGZfWrbUJta1lx/jBsUqjJx
7Kuod4DFgQga+LGf8HcHf//qbkwdsRjydVrsIPVdqOj85GOBUOWPXuupsei9
IuA4c+5IDlnEtT0AGXB+ibtJ8areRffXHb+dSkdzbPTmuyFe6uvfO+bY+WlL
4PbwbpvJpRsHxHzWCHcRvxdbFiWY51S/LVzqZCTJFjcHm5MexDSVhunn1/qH
pW+ncxXMSKMPWLdsQyVhiibmvP2cA3AzHm/zWTzOc8euq0Ihfr4hXKnzd5+8
Tsr/j5VLVcUSAqrX+RIgrbGiuGX9pxyKmCyBuN3vqFKrXqQjEO5rmVsPK4TX
NB9uia/Pjq00BGv8Te0vnkPjfuGdNrc2iebsPXHU4ExD31va1U+lsEXd7/5b
eoRX4TU/Cw+h7kQI6w/oRQm01uHgVHEa0Ruqjp6At8XQk6Cqw14FPSaBFvYA
n4zngG6OWV1ni8RYptrZ7V9p3cGbCzwGvlxxkpqeiboeFFrVaBCsB+HGkg6q
O2M/IIcW3ydX3/R2zqKTGUoL+3jnRn8rDXwAJUw9EYD2/joK7ZH50c2tTCAh
igLIH9Pp5wVEWJ48MJlgnJ/+P3n4TkvqXPSZhX+1Ut3Xakgbtfr1iebtzUFN
gfBh0jhjRj4iPjXRnlIIhiH1yR4RfZq5eiwr/kTcAe79KSZtJaak0uBM7sLb
KsFekY2p7PZElimyT0kSb46wUXpN9LS13+TLoVuyp4pq+ouhRTcIk6YEBLEv
aE8ppALLoAfPX1E5jdo0BS+cLfDfmm3n3V68T3jJyVPJlfOwiNqbrCUOvrO+
GpQEeagvkqgUE10/WTvTGTswDM8cbaqLnzXh1fDOATzDbA5wlwb//7HuzOZn
5mdMsoQn1gHU6fGYOCG2xxlf8ETl65mxdrX8nvfHsVd8l2rWz0MZbSg6KuBI
DwaPenIZf1wpOjO/8Hz18Pv9h5SEG1SHeYLGJlpijTEVdzV/quzsXQgzUnKX
nGBYVVcG5J8FWxQqyenSFemp30ShmLI4OuVgT7au3IwxSjsH5pXQVPIZfYHY
2V8q3mH0/WPEjosLeWwWduwAs7sCzi2wYpJo0TvzZODcSR9ckVBjPpO6uM2D
iZqT/1JYtz207+CxAzlbXj+tHqC1lLJ+X2YrDmN5AhOAF1O70SF+m21W4S0o
CFXzP0SfOUld676CEDVzNN84UOwgf6Sz53BWqL0aW+Rop8B11IegK3PBSSSC
Il03njoTQHecammSRFln7EFSjv98E6nCoXN5/Te3ML4Tgvq/kQRXx85OGT6y
FavQ6aVs9uBZUUSUiJdlNhqwt/dSWScxcxmtz8NLjvYX/256VEYPv8CZKHN3
R+NimiWWsfYjuFUh/mVwvYD8wwNzWUJupDMsscQQiOqKKduGWuT9d3ebm+kf
ERIOX4JvoYPalbMHd9Wms7DzVnFiyLhj9rFFeQOi17XZczeP7eZOf54zXUtp
3hAu7Fw3h9o1jwr/AJYhZ5mIAW7+OZAxSIHQSdNP8djDslTDMWdThgfKuqtW
oX4SfT4WHdXDy3vAn3ztYaXgfEbGzu0//I/0BA6aVyEQaYNyDpmMrSdns7px
qOj5z3m12WhkM55x6CBYNtmOaSagAE9zrLlFOtYmPj06wJ3RBupkY4Wk05wf
0jf9vt2aqRAjVj+Hr2jwqmHvuMGZHG3mJDfmm7//EXEIbJsdtQzdmIaMJsP/
4ugL+fQKepJOUbg9+bEzKW+0KnSuSpkmCa++SozEpMX5EG9hoYFva3IyuP6T
3HicT9jeMw4fKgtnGxo7xpGPQU0zk0D2+ksFuBLLXkhNvveKV2ItAk3s8y23
ONTdwzV5UiUPBBpi4bAX8MM/mQDITVgooYZptcK7W2aGtRODBkl+FBhQ77sa
23ybssN2wpV3rOe7wRAEohmhso3tkZPBAFMBiEpIakB34aYilkMiiM4dY8lG
id3CchBCgB/DaLawTndvBPv6KeMHd+Yxf7VaThjgx9TBaCo/ahn7wecyb21i
Q+kaegCClP6GugcrfAUJ+pi6DyuuPMQbNQbNj+NOIYyjko62xIkrNDnZ41iv
5H4PqUuntb0H4n1H1Osl0M1o8A8gs+VapD0RgbOGPZdLqiyLfhYykW7JNqse
pMmx/xLosK1FVxDRV7gLHzQBN3t/dpc0j68N+JbU9UKR60Cjvw4Pry9rIeeA
OrtmtOmuzMJtUt6V1TU87Czh0hByhIjm5r8n7BLa2nhT2TKIETluW/jWkoLe
pzEG5JFPr8ytcKfaJslYEQGUc6JoBbnSMok1gcciJpNclwde2xD0QKgEfqeR
Jhw9pWa0/zMuV2Zy5gf38HrFaQYxyVxlWWuV8vgAk2HJIRj0VKGuWdYv1ytD
vdMhYQkExMNsoIJd58G/oh5PCUkFs4Q0mP4+1cGzshGHkcbDR9En7d8ek3JX
GeY7HI0uBOXnM8hLC5DXsXHMEis1qsPLB67HtwtjCNIUhM4ntNcxOZuTamgI
7UiQzUv8lQty/2kA0gHXbiQRr2pIP7u3LTWo2mqi0r8PAi0Vh3BFms885Tss
p9gSPtB8SeW0K00Eaf1oElWgkG7a+hDeZ3gdgP10vymUKb3cZNW8wu0ueTmA
3Hn4oOA0kAWN7lx66oR19+nu1cMeZ6QHgudreZp3q86kD0lWgs5cqKBfWzrc
fxdJLQV9uy4hwZlQYquhDxNVyECfcMt4GjmO7HeHbG3mcDZgt9QrQZ5eu1mh
KhgdVBAPs9pH2BUFc1n6rFPG7VakC1Nqp+lC0hUVLI6Bbk25+q/r4HJq+c0l
I9yg7Jz/R/pRbbzCaI7VZzFBQVY9bnDdGDKsyHamZ8kxsWQCP3dufsGwE5/+
slw1HA5uN4ZzS3TyRx7GSJCPgclZTXmFOwZbXeUFKVfTqmi2uD7obmBdntek
ki4t9UdcgjCgokA+Cg24IbTEi+yTf1nDPw0Ip1Jdi3vWweKihnuJTVsOiva9
oFDn95EFs+bw06Ulc5/CCKQNnlGzTjL3m5lVOOfkxjNJ3R2if0N1o2ObAVrg
GgSDcWKsnElALi/ioLd7bCmTTR3hV2RhqaXqjLP0dYzK87LUi4Yqe+HBcAyb
lfq2fG9ikm4xaTXDnlHXuROGIrRDMVuIQV/8wDYqZ6K1CZFI3/I+hetsHbsK
kIznwrVNtX97D1IAYkWbtVzGQiwqDfLyomvsXOqPgv7H4nFxsC9CWO+sRJjZ
mtuD3G6kMNQrPHP4tVBlHWbIbRe0gUK1l9df++0gJC5Ryf7RUJdoF6nBHne/
JiZOwEZ2d+vuIi6yAAZMw/ecuAl8KZhMN8yYh7uxu/icmJqoyxviX7YvhcYV
rLGiWOMUD86qEenEY4pTOdQcR+uTqgEr0krHPXOzgeGgcGZXiPaGPsaVpbci
/x1IpCu6QCuPuQiSDR12z0XpOWOMWA+B255D3Uumu+KQh7gqke6myUA9hRXR
3jhVDUKjZJZEw5KLMDvK9aVpCVtzQOqtq4vCgMik43FgukTLQvJkYBMooe7N
3SW+nsWi0QIT+1PXBWQOnQjbfdn/F60tUlLbesOhSjbpFwIKdngXg/SSgO8T
t96yNqDVQABM9zfthOUrID+d1pRc+Hbg+OzBvx7QNCTTBSUoRMOOGvpCM6fU
0BD4m8STCXNYvD/UhNB0KW1Q85hvHhghzjGl7MLLkFlqoXfQviYyITgutms+
AD8WkDX0YYt+nQbmh43r8A1KdOa+YwBOGQ/c0xHZmO9J1ZxyZA5fqUEsjAOY
cyS5hlAfCuLuhUkmlgoHf9E7BBTg0I4syd2QIMRlbDOmBOmg25DbagqHFbV5
6vb+Lk8uoyu5zhgaT9XCT+L2i/vUTKgqu+/5lPD5Pen/YHdXevZqLBBQ9t6/
ZA0OWYm/a02ML0V/jeiN7rXvoPp0nCiLzg0WP1bdKOObj1inQagqMdXJy50S
tEIHbQLYVk+H+7JnfwANBtMa/lMB+g2b6PtyTbk91pNxrfA8xjr/EAG/MlcU
HtM1G+jYiyJPfb/NcyDclmx0/SXkSg2nJVu7P271cf1wOTVAKNDdIVWnqSo0
2xGznRPqzs1vCpTbNYOrLz+o0UBs8sEmDtbAo1qznsdzZBt2fgDSxWZgzuqE
5435kP6VJfQ8Nhvlh062EVssgt26aqngjXvgxflRYoBGafLpwScMlzEYYDxn
yDRdgbN5Z1EPWIGHDWVKGdcCwrOyEJEKy6SO2y/3MD8ncZVZRqeTx1rQIsms
jkES0+DDITRYpYp+ifviUz32r6t6e+gUaWpz1ay9up02cuEBk6SAoIvx4vzp
N6UW2S7CqsO3nAv7JCYT0vvfxJ28yL8tmkMbdlRwNEzFirdCeycT/7u9LHij
NE3C8LYsW1B/gjNAGHzqWcvD33nUH5WSx9azpYWo6FW0VF9ccC7EZk3orsRh
RLgIWTRZN6XNWaMcvH8KTNxfQZvQTSsGuL7MGSo8E+rR9rKCIF5shd7qFPzx
TZqOgxHcjLElnKOxjUlxwbkH55t8aITB8+NLBnIhVCBt4Heu73mrlbMvkJW8
EFr4PIGAAGMqHznPoO5+2KMXP8rynczGKbgtSQXRi1YiXui8AXlMbwtK3JFX
AZlY1+LmxL5E/5rYT2H+7Qeeczc0yymSxxtf1Xtjdt3qIxB2KPpiaBJu1WYn
YSBkkjKbkSWLuOLabkambT1wZtoOBGS76Ixd9lnOXCc4/e0aod+tdQiLvcXe
K7bzytCfyThS/DQsdSYqJde5yNQfpBC92/FZTYNKecGacEom2gVDITvspgnt
eflVxegooXq/Bs3cTMyF7Q0nEmFEX/IgQjOolHLscb1JdDf6tMkawnjFdA+8
0K7EZitV7FnFwx32NaPQSj7jJCYu7WOcT4Dyzf3J5l8jLUcnxe8iPrcKgNl6
EUyO0OpfUXrUTJK8dx5KWWFV23Z/llgYzsU5Dm4NTlL+M/jN7KD0ChFh9e+X
mL7QfjG0l2+qnNuY7Am/A5oLHlxWdb/ST2lj8cvva2FAOaoNkaZdtMv9DZPs
cgwDlJsDzFdnkEaypDpps1BQ1Jai8u7nj2p8hqgVSdjRaVLbauaHpr5bXxvc
IFk3sM1Y5HUxOJfkPTTIPV8gFu17ryWrs/PvlI8BN4SRJjztFGgLvIbT1Tf4
Fv/CKSETStqMqXsfxJ1ZIAxZdaR1nFxVIXI6GwtrFCDI9ecDTd40SQxFC0iI
7p7SqfJCrY0jlgfqx0KNSmZWSCov7Wm82YRwl2x1iseKTMr7+JYM48DD2BuX
a22DjqYHFWu7ieBnT0oIeipVfGcMZ8z4IURGwoAOF/JvOGDPDnIl0b7+F6ds
1hHddhz2zqWTb3P1J52XimqBRucrpqnL0J/bHq2S5FY4UH986XwNZSBGTOrO
hMD3SRb9JTsXxZnFhpx4CiMqpGHKqTnKPIq6/TdYsKcH8oOXRvm8Xb9BIL/9
odSRp7RslZf1o7qx+lGCegygk3Zds7YWS9h5tvhGGDQ2zOv4uIBqeIycQayC
a+AOaQw9pjtuBUCspIFumgnI5gwlpASN1rqI0nxLubkX/HROohq6/onYabZQ
ivnIG495bNRrp9m8Qwhp1C3Z0oKiM7lkmgGVe+jahCsdpemi4rNx7NRIvQic
Bg6dt/Bp+PI9dcfk+yO1O2jeCUzYgc0f7RJbzDcCFvSIdy19WP88K1RoTALw
qWiPOX1azfw8gs0GSIbA53y319AyiPNj0XgJF4PA2f1E9DP9L0BgEPcsky3N
7/SUkekYYEeVfAmY3ICUeT1EU+OIKZkQ5V+X32g0t8AnszmzucHddsTs0wiU
bk/QA5S2TzpoQD82SzUXjlu3dRYvaWPH71FFXruqMnliK5MdHtVeOWzwhuCA
6OWN7N5I2FPsib3aP3N3pmsshjE+8kgnK3Tkpzm4ouOwYfiS7KtFbiPsOYGv
Ff8toQHVwv64pLF07soTCRu+pvVVen+cCl7QwrIZqYlayMp3V0Pvkj2tmeGJ
GoAhv87mQErfkQWZ86dA67LFF5XjjzLedJNQjXLvzyPCTMJuLYvEz/LSXsc0
QQ4G06diysUDFGEVaYQCO8izjFJi4KCpfERfYNDz1fJjJyVSAgUv9vGf2foF
//PdWTCUY+l+M8+elmvmbnOn/rR+YVOXehDKLfM9I52/iM62lbM+EMJwGevK
4X2O/qjqK4BZkF3y5vn1w7o2wDgQXx2NOZvAE6CFG1vomjV1MDFBwP6UiABq
Ssa6m6PH74PaEc6bvXlsWSCRFOvwaHVP2OEdfXC/BwvkXeach5NiG645cs/Z
KHok3/J0q86AbpMIL+acpjn00w3Joz0z6vcXic3XaeT0YqFmxyuGdWSuq3tb
3qmG5AzuxwruzQwQFHj/m2YnBtP4+qPz6PripfGFV/4knp0dYSS85gZLgW7w
sUbqjZr0Z0RNwC8ZQxwGM/mnTVB+hhbLrlolG2hXO00s3EUhr5TSL8Ewrdu6
5Xpp3cJHSqW1XVNyNrpsx7jNfvQlCdFr5v3thmChGARqBS8RksMIVikfavc4
T+HjItZjrfQ8p7TTj7nqBbJEntWBiJX+IernFy6g8bVTPoP0Rx07upOvoL9j
IjsmM0gINCmI8kuZISRfBW/zV/J8T0sxAW8im29qtBWR0kd7AURj3lPmNDfj
qGoTVy45sUWA9BK+rMwY29Ljh7+VKPXlBv2H+5WAdHZU3/4POdP15HqqpwH3
vbKRUl7Ud+f9XbxeB+KdCOhBGFfx0URxI+x4vuuF82TfTf0ftriA08KFp6od
oj6S4b9fKLf3aAQezrDRVeFqZN5APZ01/bl02yamnvQg5Kir7roh8aT8oZQ8
kwnynKzijF+O0sPuZh3MrLrPFXTH/wDIU+GJsQ0zD+p8xVIIIPBZabT/lNAa
SnQ1fV1Jb5JZ1s8mx1jMJ3kLLQAanZW2KawftA+60HAhs5GVWO3HfZ9ySYmH
p1czLOLZnXQhTO/OFSjWDE0/BlJq0JeuM/cqfQAk3RTuSNjU8bMOzHskxHEp
Igl6agGx6w6ojWD4wn3CzsRRx5fYNKKETGrxJF4wdeoutZ/CeFbWKUzY5qeu
Ra078Vg+/9+l3DDz76mAUOY6fKDW4ynfPgqxxk+n62MUDyGPQzb1QA4eHQcv
GTDyCB6Bw+zuGXZkUidXZrqyRgwZk+0TiFmj+OcyIDufcyjHhkRVHo9ZWvH6
2LNxVSpZGbWqg8CA9esNgJsfgEZolLyZ+rRoVPWPa7UUB+ACp8GWiat30EAW
MPGGfnUFJd2MlyZKe6OSsvfl7S9g3CAsm8XAz0gH2xtl16SQHIv28FTqjtqS
JoXiZi7VPUKe29HLs3O9MxwYpfG+2VgnGdjk3CfHTMgGQTdcd9lmjT3CwHW1
N69oIJD+fGimijGJ/LgqhBi7SeysPeCpYG8PQsJNq0L7lOb33bfcwo6uHtj8
8RZSc3agAG3ENI7XIq2dDKrPcddQlua9xIpJXxedjmSwlRLm69QMI4yJJgQ+
FKOjbCOvdkHvzZUjby5C37epWmX/o/BdB7liA20jZShgT7NnTo6W+0Eyguh/
aEixg6y3T7SdKbLPhXKklB2dVeS9FJIQ6AipF6pgMFpr4qG69PWK7Cz4wB+a
x6eE/bbi1A8eg1UrPsCpmeGe4quzgyPL0l5aHbRXIfQ4vM/lq2ATU2t5+PvA
Iom4rIarujroeP8vYl5JO2kTYgzUNhvZPrwdZRYw+ZtGEwowTzE2Pxcv/2mR
nuRXIshY6aIte2Q9KaavnNGG4c6q11zjFX0gw09580wEIWl0XsEIs34DwCrV
SjZ3eig9W/wK0zelKad2ID8q+iF8rqCnwTbXCf7ZmFVHSZLnbGCS0V4cM19n
akN7d4s43Sw0doYPdwoK8EJg/H7Q5k/NP4pp5DrdKGa/HVDLDleSwG/s8V3W
F3VJ/IWwrjfx414IQZXaon+X+YnrY5yP83rllik9/bXqyy3qtygKohZOjkgR
LK6zgvkObKiCFRRWWXBYLKl2QYUwjwAtQwRPTTnNyhSfO34eMMB2oxZe0zQA
k1XtAXhy3KUE+uxKTcnjvV+zifO7MTmZyUmR4DvmE5Nl0gPdTO7tq3fgptSZ
uj61stQZ8FRDaGlpJFbsJN8gtTHIunQ2nEBlGRADrSgX4jBFkYxYTVqoDukF
rWrcNWEEcNMoxBqCM8uXK/jJ/LM9Jw7oevUzOj964tJ0lT+8kSC84kOSZ2js
A7Cl9H2EL+yFlNkURT2ejYIp1kVaqeOPd0ipd4cUU1beBB/tOzMwH7KvY+zS
KjNV7GBvr7I4M1q6xf8YFiq6+q/w4vqOHIdvTxUxmwYHDu0IeScBj/5NAsYV
7gpJemNqKenGNfuj4UkaYQtSHNBuedZDEaaoaoquXD2ET71927a3GS+Lzn3k
unUrrKxl7qebx9sBK7o8QMSBvmBDJny7hifH/nh8kTLbUSZGi2r+ixrz9Y2K
/x69VHxAZ7LycVOHujbIiYFXM7N178KLqN992lc1vznSjk3rc2HXNlhLsOI9
Egknb0FqngWu/UqtyhdgHHJjopBHCCWdy60Wm9dm0EJuLloiUx5/UKhxcpFd
Ja2CEcCieJnJoJeTZXzJ/ND+uS57Jwmia9YoSodpiG77qywgrglv+artMegS
ji2rylie7PYcDmkui/oBwiLS8JGXn63msBQN6PV8w27axJ2PKk1jVMjF2dCb
tOamg/l6nvcs6b415UEd/MhDestiqHpTCC6+jisysqcQ7Dd6qGCzKYcoqdDP
hYBR7EywDoBffxBCWJKZaPMGapTyaTOfeqk+121r1RA383GqQ1PALpaqpuXG
GGhCkuCoZDaVDguGMvkBHFQGB8GTieKBU/Nu9wIFgQpAiDvXECZHJssbT3dK
OFW27/R3IyjGkpAAJrtrpZrMH1LjNzUSQ5SO3Kg0r+kWvDxYW5fVdff+2ha9
6bULN1baIFFAzz7Wy6IKZoz3xxODoZyEvIiDlLffYkVjNcFE84UI+OG+XCSW
8S3unHLqKVoWdxvUKpCXK1IyAhwIQ3dpbzHi5Z6dXblx4ZsP15ZLyVSzpXwe
98V+xBJILswh7YeFfaK9MjVGavy2vSV/QDgXQOGpOC2ShYY74o16r53RXLju
JO4ZjtNW95oi5/713IgGzFF2ui1z5lFvy8ioVqdoonoIzQihMix07yQBQzfd
JjxDRKqonS143MN6TwLrDV70oggIf/DGUvhpt7Hbo6YunFLqw5LVV7uik9Qz
/bN5mcGCw6nNVRavCoX1BZo/P0EjvBSXxlPct2xvY/lTk7uwbVIh3wNHrxlD
weSm/RyogYDKW45u9ZhwmFTR8+e5Qnvf1BZL2ix0OdXGa3eioMNKS2f19Zck
zd6tVWvhNRUvW17TUibO2lmNW2lRyLLzAPnz4ECnL/ARRw7itowb1ld7aEaz
2vcLBI7aLS1xDrTNTqgnjbqu5mXn1giDBotYvvL0sJOILMrzpN9GUldllfjQ
npkZlcD1ZHrkQJ3SmU8s0xvNP9qEEob9EynO/3TqlbABiOO1jM7YCJwwcPXX
ZmEAQj0v7KAP4WXpTpsxN1refqzW+2B9pnwpZiNv837jnaYEIyQRMa28869V
pt4ZmRnSJxpqOCdqzqRp91fXjEzLRJk/AI20W3ls3pmdJQnovFCeCwrI0DVY
LB/ifdXqDRIao7zAPVbMSd2tsZXxLGlYVO1sg627eHKfcMuSy/yVciC1rw/N
v+5tCwuQwCBvfl9+1C2jI+LqQYzVq2YRXGDvT59oPM4zXAPdoLcjFILXvQsk
gmnUeFc2htAO6Ij5/Up0WX4UUjqgzmN0ug6KihEM1KIxvCfORii2TSbL3Gb1
s0Fdo+itIXHyKO4YMniHDJEG7trAme8GHVjxlXhzXGy4veFPENCRIBKAzJB6
28OqEQqQ2uASC6+zo+0fCQCYyPjEvpGHX2hDYvGdtSWEqgZHYA5/TwzMfilU
WpOZFiAbfk5nJIAXZr1of5FFVeW3RE/pgLUa5kjYjuqxOWUJfM6sCdOcRAVp
7sqYn8vBAxTUdkxbxcTUV7wE+FNMu3FXZjBAx6CUp3BfMA7dU/OClq4yRt3B
WlsCkIiOKlZFfjH+LjkFJAQZpgZkB2au3rK4aeCY3Y9qgSUFqcQwcvX1PUmI
tx6FFtEPP6RmXWY7PTddlGf4jL3vRqse6VRg5KoYXq5s2bL5e86gUgEjFUa7
FxaG6AYaaIRDoIkOUG7s2/vqH05nBcSFR0s0Wwmyku2FnZ4qLEkOf1WiznnQ
aldN42ZoiYkq5Fe2KtVqRErvs0TC0B42w456WHW3IMr7herNYkJF5I19U7DZ
3yt5U12glvbleyIHycA0AeJKs9FQEOnJGybmIO5fNpaqfJzA2trKhcUAxlwz
+PcrPxeZMbK0t70GkbvkxZEeIf9AnQ5YFCAOVwwN/7bQseopw0kpvVgA9VUR
VfRgH0MG438SDKGfgRgTR4J4cxsXXAz0Ywq2fq851A2Ae/YvJdH25qvJeqQK
m3ls2y5UgRXLSg/WJObD1F1/+q+gez4uXk1RBvhyDOMxCe1lsTGAwMwWuE14
UVoIUb5AzIFzo/Ij8q7Zs8TVy/zbzDxV0WqZF6cKelpj7p5V7g6spZowFsfY
Av+gi1Tr18iKnr+TP+ypkBtsUub3mypa4D/A/WtWOt0DTjFuwl3Akzr6MiiR
PwY/7MFcaGssDlm94LK9PQaDiYoNNY6OpbETdVQDaW/7RtZhKlk9dKx+vxEv
F5Uw0uV0m0aOrUybNNiThiaCdnQJpAjMlocaCanMa5L59SnCQYGYV823Xewt
cyLi2NbGG/O36TCzyrimsj3HSknf2Kr/gN2kZXR/MXEXPIoaP0P3ZfeFNjC+
B1KYvvnV1GtNHhQKhHKV8KoLsya83eNYvAhvMBQB1jltnNbSkaDH0ZRUlxPM
TlI6bJWr2RLMljV1GjJrF+ZHh7V3BEYWG7MtGnlVXvNUeQh2q1DjAdoMnLl6
BBgQeI19W2nHqcyBwYz8QU6sDjGlunmjNJSTwxgur0bNccEgj/GpdiZeozPn
qcqBEvrIvBbBMZFIRAmn+sOLJOabVGBwnZ3nLkaKtDPOdXilkYhE6ngiJT21
mrf/v8JLHpXrePx5KOfnpOuh3aFCPP1FHwgaRh9k8WHPzCTuv+XTCL0+2G05
355yMtzF+wJMMXXUsK0JPUGZ5fbw6iLEz8Kpdw6pYXRt2Ccmakudwq3yLlAJ
wDB64PVtzUv3lmslZkh4cpWHRJHjoQnEnpNvbQS+yMsUA3JXJ38mclU3oK8B
fjiuaHV8WYrOQVfRGMnQj92S7s6j+ZTobovxVmVKPMI6Pv3nw/xcLXFQ1LL1
RLncSZI7eKOyfr26nVUhJt6o9PZo7dZCZkZkKYP6yGTpdBvxhHXXXszC2ywn
xquO1xfo/czdFucl6+Wsj+2zJsBtEc5gX6q6QpDVterwK/Gd5sD7q1XAHXhm
buwXyiheQ7KXEnn+rjPICrRHh5OZ/0MvP9m4Zhz90w2LfGsRKgZyj+1p2+zK
a8m8+BmeC/MS1lvgV8ix2ti5+KIkWc5Gi82QcPV/JBSIdkNYM5MO2/iDKUzr
dXNuNOU062xvZ23H30JPldpQYKzbug+/0dRaenQs11kx7KCtux0du/IwNVRt
w5rVWKA93F28DKB+tOGPP7w+lryZvzqdENUDSYzyL0hQz3mCu+wJf1t1ri4w
6xXgiQMAz1plCA74emKA0GrMT5JEnKLMRH9iILoiF78AzwlHWpq8nCz/Bkou
Q0LFlBsu+9zZAGe7OeNlhiswEnSnCuXzi1WfxmdEkzVC93tubpYXnb9ryNx9
CkqdISJOnhTg1aYEAwMQX6tOx3BSoqRPanddYdQSTEFErTJMlQE7P0uSb1t4
X2FVoWb7cSdOAVHKBw0AoFIoHrZGaerSPE4oHIeGT0UOqhI5ZWAHuhp+HEWd
LRUdI07oCrAWftvG8D5r6yt06Ee1Z0FcFsFoJSPW3FVSETxVPIj2AxiC6jcu
nXQ2TtV++lCLZbVX2F7F0FKArjbzptjmJpu2Mt/ay26BmMR/SG3v7WUNsUSQ
WdfBp6SvqMxTj8UxEx1MiB5Ahp4LsvRNPv7uFfe5dbGUNmMyeHJn/Jm+RbvW
3jpbUpVnwcIMCVUZ2JEa+Fo2iqPa1bj32Bo3t1pu2/cDewckNVhrJ+uSkhnm
AWSQohNiMKeF87oR8OuyZNbJz/mc/4Crej8VDpY4wWtadE/PYiI1tPIBq4D6
er5rr9Yw9VNOrqLqM4D8ETyE6VS1R+sUmGgS3hl1EIKQoo8V9IDy5+N43qYt
tl34WclTY3WNM3cDYCZgULVIuOnkdg92I8HFslrThjZKZ22voI9QeVnBRfR3
SdQ31stxIHvl39lXxDWDzIdtf22Iq2YP8hLuWdxQJwREIB06njOOuPepK1Wv
kNjAe98ePZwOEJMnQd9PaMqACDSNUDU2PE7TbyV/tAJhjtTaA+YzV/TN3E0l
mClH7RYjnXD702/CpPZMqZvjs/G5pHD+AMKzg6+sz0htflqVmTTv6i8GDVwf
ykD+1IQDsamYyZjG90Ar5ea1TDwTZrpXSlTjKx4ov/MQYW4jldoWGVkh3hLM
3J0tIv8qg4REM9zgqWVor+4jbDNB+68xjXr2nU72QxDLHB7WLAkxGLsvD5Yk
PfGTr4Im5mgd5vGyjL+NHMUAe15LCVXi8GDLHY3M5QURVnssgA+WGABFceEH
24rgCEZs4GCeiWBoRk0X0hTKoUFuSewxUMXyu2AY35qY4OFUh3vjVbHr50hD
mp7A86NuJdKUy7sfR4O30lpwEmf2CcA9WE1xnE98SuzVEJpMBccTIudbI0iv
iGTuetM8gCQQJ16SZ+hzDWtv4ZQOWu1doBjyLpJ/2txoXapTnYvMc7Bot655
xrd7/qeiIt9jxZKDc6RoG47LvLeo4NSIK6EyivN6+vMHWEIPMvwfIF630mpO
v3Rfo7e33z9HHcacOeEbr7/MuZjCal7MeF9rh+Dwj9mKZfbI0eoN7N+9e+HE
DVSG0Qu/4wHV6LrW5SCwkBaYu+VvkACuI3cfCdhyGgRbL3yz8qaROo+opbdx
Q5Y254W/jl3oFrODUEIbTQQdGc209AxnFyzv3429rtnoKizAf79PPHuEhH3x
PWtMYSV7m56T/50kcIMZbiniFM0Lk83x0+lmbmiudNu2Vq3woQfi4XYaDyYC
cisvn3+yTjJNNQ5e7gbj1L1HOR+hdAxm4Ak4Ypr5wyRX5jCrDKXLz/4lPQA9
yuI44G8MPondRdwQp8D4CVve9XqEup2RkyVVphuIZTvk2qmvz9y7bwLi6Vzy
Zh/MQRbwuVJETd0OflTi7cgG3icveS9VVkqDjOqkFlZbJvMPpMagfrPVu+n0
gGiraKZbZ38EWeM/nuj67dCgiywiBVxgNOuLK0zOAP4no7yq24oa3O+juqRI
D8FE90ecpnvA75ik7fN8nwCn0lcEntkYXPcmxifbsEP7sINJobJ/14zPUWue
4ATshxteUBYe8lOMdF4uDvhO0a3qYEwL2zcyIXBSppFMQlEGwQ9KIPHIe2HO
Mxb7ZNv0fR2UKBfP8R7gqcgEYzeCghnU2Yy/oKlmcI1Ht+ChZD3wOdtIY8l6
TO+LeBWID9aR+fAJHgleoWbzkiSR/RmnTuuZ59X+8X2aKyeV1RaO0/4Ho7Yb
te/Gj0vVMLcyYSHVAtIqkN9WiCUkHL7jg42DbkxUgWYISIWcGUDs902WMc2+
U27wOVnI+7yxcSxJVSHPO78XXTwkyaw0RTjSFTukz7aa9l/04ZyAAhfqT4Me
Kvih7zv+1VPOeZEw5o8qrEYGWGvX0jVrq8rCt+6ZCeosxvg3OdhJtfKNbUob
JiUaHilePMoU1Vnd2lPWiEQA4TQWOHsqsjW6luC6V3BBD/GX9FQPqNEDP0nn
P7SpvaayYkolQ0M7dVXR2tMzrqev6dAt5bKzlR+RAssOAE9Oefj8WdyLcZH5
PdTYx/H2voVFY4zSowBH3MxmKF8E4klQRCHG9NgMYmsbMNi7q6o1pWfamtIr
ERN02IYWUbKkW+alRMTrKvQzVk5agW5JzdCKSIDh89GPrlGk3KltOtQUmubm
w4O0zJiwR2fRcbnxxSLU3e3Rxw/bINZaqdCEqURQizZgov7eyRpr2OJmn+13
EimiKV135YoiVfDoaHgpLrd01ZTjdtueKU6XI9niSsYMBcNtqzPcUp9A8f9u
9buPp/QgcPESORF+ImpWVeLfK9OdD7PbaZ5kgmCstWePZYuhsf1VPe5QQIP/
SYXPVBl4xHCdVej53TVjwbQqHFkhYy9hk6Lu0y/YicsrVmUJUpxbz08YRIWE
4YppFmXeoWRBWycF+FhUWD4JhI/76rjXRk2cJ4M0CvwSejxJcHubWcTS+17p
XcXdE6sdOJNQfBe8gFS6XE2OOW2qEjv8ZJzi6G2T9iFz+4+4PaoK/KmfTgES
mu6RL50yXz/vBGE1tytz7ZNzkXR9TGQReDE7MGgEK4fzzgBNxr9veJzIGGYP
Cw43YX4Zc1bYUXSS2NXGKBjj+sMdTt6D3G8PG/kU/Ytxsp9NNDRO5dc/cNXp
KbgAtsIK6OVqkqQYcQRDzlNYZJgZmUQPFcy7cOhbOA0AxNI4U4XeV5qYn0Jr
+yJ/em4SxRSjUdG02GIlRZX/TS6i8enp/Ap+YY/3QMpmBoJeRN7/vmS1IbTD
rOAR20fOgjL713pjVrp+gLY3CYTP1l15u82zLzIQjRKYDTlj1Ozpw0I+ZCIY
3TzAT3H2XOKaQV9eU3/CaRGNOmoNp3OsLStGmvF1TtX7r7Dxz+s0H95Of0Rf
dOgj7pqubOIqNCMX3UzhVyOE2s2ciQUdoSLLARArHtyobPDaDqQzyBmi25Om
sIfhD280I2XCzcsp5Olqve7BefmtTWw5k5faKetB6Aek7t8HRJNEHB435n1e
Dr2jAjm7uu5w8eeJGEz+XNOba4sVZ1udzD3WM9NreEd1Kcuj/6tjagRNneyQ
jb2C5zxuPwCZkkQYBHPsQNnGVGsqu/SKVcYyMIdqMUteOJuP0QuSVtOcY2Og
EWX8coR7QbMb88c42X/wpEtx7Un0mJGxIWEOT89OYnT3/+2N+Kp2vjW8pbGO
CA6qCy0Z8THJcRXdFheWuajJgADIWQTA2Abc+/47Nosk5uKpNTz7OsmwoMWo
lV4h0uEoMxFkWRen+0ooGh4ujjmNLnLpECPxTN4XHcxzdMWZxf8r2RXmMt+K
V6RcSnY1MnflCJE+ysvi1K7/obQSLKa4582bmyY8tdlfBVLLArIUgUQrL3NA
NQfIgVlP6j5FXDKv5slJCScnPGr2h36c75H2WSz9TR+GZRoWKNyFreBRF8hT
PQH6q/iONrQt0/F/YZQI/D66KZiMZgbYFw662ve3ZB3mgurGJFc01LTacdCL
/QQH3Z6IO+AsvUxn9XX1qT2C9pfN3hkevjYn35rSgN/j2CrTEon+ToOfESea
sJkzgEIxisCbmVrq09q6OOZUYcmeOLNmzVOsso+MRdq0zVBC3PTOBdCwZqHr
W7B2nYtzgnX+Ad0DF7Q0ZYDUu2cvAmZ1rf78UXoCJ0m0AXZh5Usb2oSyho+w
T1GC2VsIePzVcHr8uPVU+k/LJO9GBWq69H08U6ovdZvs/wvobw5iELhv9s7V
a78ARf6dz8kY7ksEY6XbC9gS87CGANyp8UpupxHfJ66nYCq1r+V8jW52h3qS
Bf9/er/Lb6ZRm+LMLYpFng0ruCkBUTGslgPXj4+xo80SkLWNePAIGzCj5xBo
SzGB+3BDJzK5BZkLFxM2sZbx+6n9oczOlAVSC3l7+cfTnYzo1TCUW6CT2znQ
gSDcLh9D10tu//4SsFZhc+I2D9//svKMkt09G2QuO9t4ADrqY5111PqSiDJm
LrsaIHwNz1MXEXosXTwf2n3pBulciuUUEeMMM0ndxgnBuDSD5KayZ2YSUNBX
X0L76JwFHRTcyfWucAdbjytFfPqApKI6SJ0gA5Z32gVevOkHkHfWI0K2uf+g
jU8e3EWZTcWDU463dFxzj4O8TwvXeh3ktvWDEBnZohShgp8hlSV5OWb8l2rE
LNtKNUSEDaPJifcMKjsJEPlLqfsfjshR1dywfS3aSw6cB3zEg3Y4Qwc8woaK
Muk9Oj6Niqx2l7pOlTUlUKrtKcBDNJkJBaPVzpjFg8LfZn5HeS5r9aQHwRO+
ZFvWzJoSay4Aj0JWl2NcRAoWN6YMDTupF6LU9cYM0rRenQRBtJhRf7GK/6K4
dncrWH7nFYTBb560GqskeIxEAxHwjGj155gylV5ArpK0LMi/9zJ9B4jnAgi3
botqXCejuAvuJ0yn2eMinUJDj5vlwT1kYOoTnV8RDhFSD3uoSCnDJgPy9Y+O
Ci7XDeOsYeHDTrIzaVnzvw3v/7N85S+B5uxDX6Y71A0nrBCAj3hSUb3jeZGu
BqhiXRf37UGurMqpJblm7pSoXK64eejBeqORFweBdQwiIbx8WeDhlpujCNSN
eFeaXWptEoHVaJFykvOy+lw2qL2kFK5Nrtd9EYRy/wyGknBQUyQqyVTWRsFA
8fbQDN1WuBla8P8nW/PmfwqKg6axRRZRqQPkxFDa+w25QZ/s4/ERv4cEpw0y
EG0cEz8ZhVNIOt/Ny5/d0YfYObgfVKpiSAVNpMXfkYkhn/b7dqLNfsBv3v1d
eQ/tagY9lpxSPhcpSd4hp+vdEb5die0G20aHQBlGCyrvbuma84dX0xxlNwAW
cxsrBNHkYh6CHkWQENJd6hMBJYcKLhQ85m6Qtdtbn4/ovWMSqW1E+nZunLQG
0MjeE2wXS+EUesDpT44Rkyqrwvh5jlDF36bJ6aCBJ6HY7i5o+Fpdq92cmZLN
4MHZTCh9EKhVRsgGC0Qy1P2yWFWgj0RJ8Qhg6E+pIyQeU7F0wS5Ex20oqafZ
ygpG04uRzTOLzWurKcNeSMmbjXAbB7rlNmOyEAa5vRkAMZ9JmGQjroLLz5vH
MaIswf0kr7aZBVSx/nF80s3s+Iuuqj/6kkX1EmkZKkoCb4blrA/2dnzXLTlZ
aAbQxaPfKNzSYhMovGNQXZPU9v+SuWxuxZvPcaRN2Fsorc+zKuRRKrrywYEH
9wFNBppa4CP0MJXn1WPH7vZZmNqeKrORe1OgX1iZXsu170srkI1qo5oAoaeD
1iZHsmio4OkDpTLFBcNXoeRh3I5+Hr0k9k/xZuf8rpR9hYfEcbZtqwgnYvJR
9F242sVM1bBKg8+mt72laLPa6cz4eFQDOO5xh3sOs+gdlSv/m8i8hmS3dqgX
Zv5+RhlgDrDG5L1un9Ucv/HRvT6iBoG/mJBz7qld8LhUOapmLJ9UmTZ0/1Ua
m/LuLcYY9h3WbRUOHdbGaQx2BWDcJPoZqDl/ipeBjYHug7ZEo+qWGnx5/Xoy
JnSfVob9+0ZbWA9fQrXSmtGEmjrfjxppXi9VdD4itBvgqca9+ygFutmgQwGB
qmFvvvMI2tgTLW8DQaT8hH+SSUk5yFzA4r/kCURPnlea2HpQuiz8DbqKo/jw
96mKVGFjU6DIfVzvUuxIUO1aBxQYGcrkWq8yR6X0LjeT2lpCvlG6Elw/r6VM
ZlSdqPm29S3CDmmbkkFDgVeNZAvFLu3/izC37FwAobUrvdovVz8NThYJA+8n
DiobiDKptDolY8H835FDeqkGg46Km/LxnhNSXAg/6NbbUrR4mvMo4ImOADQJ
AyIkmgOrpHzuG3iWqicV3Nkq2Zqix/SbHAw7MPbVxxxuwX+YVCMfid+ZAfyp
hvVJLi5gf1bXwmEiYfbzDfa9GM794I6xNrFr57eo43MjuVGbFBFUjIkhvCUS
/xBPP2uam4PXrHrrMIdfHF6a5QiEmsCNM6QmaQHozIahtZ+j0IyynFwNWRmU
3si1m2DtsRNKbAfbqtRA3VNUSG0WfAQDg5feZB6I2UYF4h7h2q4tmt7A2udI
vb3XMqfmv4ZdoyxN/ZHFs/6RBu75/k+aJlie4lt/F1l0j0Mb1/lMsdb7sYt+
aD+Ujmu/jFNGdK/qZ28wod+CscLkJb2PzcUFv5QESzvcRZIPEcugGo0+DcAw
J9/xNUUNPdz9lU7zPVQbVNVu3+atlMzo69uoTyj+R0D0JSX4YAfa6E4jjXPk
UicMRf/3ke9KVJ2I7IwdNItLVQnHzHxEdNzWPFfwtyagBy6GM31m67NEumTH
dGFu21NjVkvOmm2IlH3+yhHhNmUsiB4xPcBOWce9AR7zYHA/VPKyRp1dt7sC
3unnMWGUcjKo7jdY0lGJg1+csQGA4MAazPQBUbx3nYEEhD7Z07LP8Bw3L3sM
Jz9kxaivsfbbjZTG93ftYGgkM63napsulsNR0gRq4NqPBbIEwf/VIYeVyfiF
6V2msHVosvzX+CsbETlk5PjWyi4jbsKX+8qSoR+0dPi1817norGQsbqwberJ
7Dcrf8h4uix8NuEoSftORfd2hzwymEgJjcIjdYUfllImLVMIz9bJoaW2IqVc
EGSPTvVEjtOCvt44LHIV1VZw8D63nQIIHnatVXaEP85BUMVAIA+DYcCZ6tVu
oD1nXYfReyQHKUHwGFzOCgzDehWL3+TD+hFQP31KXK817/QFsUNDhhKElKM+
qwqz/wiyJ1dPxotbogH/QVoO1rgauCWAWbhvaYHynpS7IYtjxKVnR1pzfRxC
zLpBdx1+NZZkw/r9hwh3ulO2GePDVu+MlwgsW7M6nrNlyKYwcZi0lBQgWEIa
531klLdg845F4EzcYnVMNsT6O7UkWVNAjsaad3Uat4qeTOVqhzdeHpoB8yQx
jBrcuGgfXn1nGDei6iklb4olO2hMQET77IB4X214yn2JZrZ21wyai0oq3QmA
//yECQJKHGUlnQJNQn9wVBu+RxCKLPZEotPBEWHfaKp73PaLQUmNiQOyCDj/
qsiDQ6jBkdGe7G8uoCqjubJecrjd0h+YlPq6kgIyeYIb5F8KBeF+Z2dLe4iM
3Nr08muL0qNdsKN959Z9RKPEWtJ2d11LNPH4dEVwHdSRssz7yIIWwDfPlGXa
VaYgR15JBgsRzO3/PkZrLfA/p7oaU1cwpnZPXF0p1TCEH6Yq86J5Spxgw7rr
Yyv2FMK6wCbar65iFRe4TQCG9bPLbZt3MgJVWQ4Q6Uyo8j8ATLkBstgGqp1s
f8E+9rs40E8NvMILxKfb02x515mrmR+w3NPXh6i+9qL7VJC2FbD1nlD8vblQ
aCGoeSZspWA3xKyizaNtEJnf3zYQeE1PMBGj8p2uf4jvcacJe3Gm9Z7MBNoS
t5kFvvBm9OdaIPLy+CE9cx2/NXrvW1IXQLZ8hvhhLFnlfNZWDxlhhGpKHAiC
7gOaVtClU7BXTcabbdazuj0E5y6l7exID2Zvin6OZT8YFvg9MILmZre4KI5m
HPR4E9t6fF2cqKDtnEMu3qhiSXSl0CLNeKXHB8gfsAPLyegnHBNCOVAiQGvP
MzFuVKB/v3i2b6LqH8I4mm8zauVIYEfz+jHN6pukFJrf4F80a0Nz8r0nRQYW
+Yp6Cvz79hNeYJLQ8kTNGesyk/Vcxz8iLuu29FPwpz7xydHr+zjzomUDNGUM
+LkBQhYV/Kvh5x7Ygn4Be4zZ7dX7F+ET4K6pOnsHsmoHyH+3x6aB/gg8QYvu
1hBHW0Cq0JEsQgMcN2RjUUXi7Nt/JBO7nbk7V9sVde20eITsVEzQGIts3YVH
d8NJnM19cEqDhgn1wiSxaVQpPM/6viSd0xnKqXOtAAQDd4eDj057apGkJjw7
cFSnbjQ7Ywbevr3YejaHVDXbn0eXuNpAeDKp2oXX1tXI+701klJHrgnhhxid
qStvHceY93LZ+qAh+gH+4oXPbB0uCW0Qd/qhm7FHwK/lDor6RDXbAY+zyTqy
8mMSjFKTq3Kq2FsHen/LiJW1hlPAoRbb6x+u5Z3SBauQNbOuf5fpNh5OKrmk
IIE4fb9Hzmi6JWfnPB6TgNoPgGyN6w3+2AEh11L0Ghp29S2VjyBlaXzPBrd3
2giGHhTxrkmkEwtwGlAeNP4VI9F4/U27moDBjyC9KqTiJfqGf1hkxBJ8yp5o
3Q+HI88I0WZ6sdAATIcxxcSNxDCYnD6b2tIdEiNO7GTmDi9+N7HA4gcZizsI
lXASTdLLl9I9BD4hWy6z515GPFdBi3/kD2XKPgKnDb3mxDA9K5AxQ5fi0Qp2
ooza/FqrnqMZdI9rrIcKBxFLYCdy/UPUv6IGtTKBqCnF8vh40Q2qgs+NoZAQ
IRWqEyUrKvuu123FG475dqIEdEuU6oojRaZRapN9Q1UQsSNHeddL7Zfumuna
fedSYe2OQNzuteIr3myS/EXlS7/5TknI4DCb7pLEwTMulrVQdXuWagjsDmQk
/aFHr2xM48xdTUWDLdBrDdGysZNGtknzPD2+fZlI3LYvQKdMuqGkY6EWEEGA
1CEeqlHZuWVwJ2Tp1wAO++Xcop/mzwlN9vcPEIE+wlMiuL7TDTqM9koZ2SYN
lY+0XlUIc82Eupd40JFb2Kain33oiH6P5KgtJZSfDKwJ8exW/pf1F9qb+BmV
y0McAxNqeVoctXfBnXtn0hidZBzJm/ycgjC99ezzVoXcw2mTcZQw0GO1+1ut
wIsxaQV/ELbhRVdVlGMhXr0t9M+NI5vpOXlxIVcfFKsfUMkuTwdSmQHeIRvb
9bJ5pbkU5N2s3YUuYH0MJxN9VGGsRsebRCsiFRzlCNLLk9bJquQBMpVDAa1f
WWYnpIZzmYRN1PSJEPTAZaLXiJ2rG++J4dFlH1pRh5ClQSvZSdlg4Jer66cA
iNjDWyvEij9b1WEpZ2DA6+jjkBfMrKg1t/1CnumM+jiw1IG+FUbJW2rSsaC+
AdOyIPs1Pe1I1GFXXbJ9Rmlarong2QpFrv8IHbeuuxdg8UI2V/wACSvjSMHJ
MZg+vrDVbjkNMZXp43NlEtIqWfUh4cIxbmTJN+M7+huw53WqX6ZOxFsSOTRi
eAK/ghVYsqodHBK++AKS3ysGVjaHXCh206NURZBk58AZDXxC3FqZjGEIVnei
v7ahUhSCRcyQVXRxG06HAzNti5xveg0sJ5mzXYnI9Cs+Bu7ctC9pXJCjWCwr
RA01NCjY+NlG9+w5NVBVtpNaxGWeHhWSly9opvCmW85zPG4EPezxLMD/Y2pg
ME7POPiAFi5Bs35Xj1tOvcEaq8A6pDxGpkp9icPtlmvB2DcQ8ikTeHcFv6kf
835IZ1bGS6mMP8fJETzKGfvT114CU0MLOkpa7p0tccmD+V9M74t7VjT3mHaW
Trj95UGXiY8BcQ/eg4MoXhqYcoBx27qnvroZ/kVj8mrbWRyfjPg3z9IpaVbB
4VU+Di6OHTv+ECqT6R3TFGT5ophYDo4kEZDJBoEajkEsJdX9YLLpMM8KBuuK
sNWIljF+y2jqnciGBZKkbbWxuYlwswqyPoyD4oVbdE8ORP6q8R2UmJ5MsRaq
gVNpSQ8cE6GMPijx+yilbs/L/2dma2p0CCxz4dQHlUaQBtwxW8Z/uIhjdByO
OnNuHU0CAtzvs9U+ADbNErnNZRxYMRegGBkfMIsgq4vhvLkNFtDem8tQrXKA
GhCXK/PR7WDeu0INQSJeSPhhQE53jY6tRg73Xv3e6lK1eXb4upzwdN9SvRKX
/z9eKx/EOjDh7UOGC1sN+gtTqhhbnRCs0CKyQ7626Ul+q0QtBkpYfCuBnNuc
OgcjKnMOLMZRwUFFH4eAHbqF3XTOjsRdVT1yN41s9BuB4ZeFamLLCXHe2Jv1
4+6hIUlqwj/fve9w9xf2rMjJiPL5oNYQHlo1OAz2wX77g09u3+k0tO/DY11X
tlp1QSIu0fGB5ZlkRjVcaKTfOFSd1NL0dwAPPyfcC6RO1NmMsT+CF46Zq5hJ
8QLbVURS2aQ9bmcdW+D8kLYkzVVREmvj3g3VVYZKyC6+Nvk/jkYa6LuLqeD/
CsGTl640uufxmogTpK45A+6n6bqIptQ3V08WUiF9uvQR1GfvUBTkf/Nyu0TU
FV0jrauZjOgXSKTxsrOn8iRt8xNaJxQ0ICnQbalta4v2G7lkTEr5UE1uPKAf
aEEY0PRWUrJpEJ5frVrXWW0DkNojIxAKZKBy1MgzvoOv3xb6ZBQ+E6Bpve8e
mTmekJITUSqzb1jB0NXpIvU7QDm78cwrxFeJXQKGIAuBs1t+yxU4jkcVW17a
hA+qOVmZIBSD36mc+d3P8p7mG5HivzCWMCwRQPWg5G8lHjqpv8rEeRptST9j
ub4/YzzAX5/XpgFCSrPigOmRQ+YrZNz9IJqVDd6PZREWvqC2xWGF5ExUEnFj
uiNCiJJHcs1vC/y0jkrmNcoVNhLlp/d47hYuFsYXho2W1kzmQ7UMPwXMd0oW
BHcRth9lhmw5baaJyezbQ1CKjXYqk2q3YIc7q+yeACwAI0IhziP1XdHgEY1t
2nTHbox5Tr3z7NRSg7u3KrpRK+4dVGs2GbIscpFSimWZitXMFI4+NuW0Hzt+
JU5C8ec1PH4VtZjNF+wQEny2VY2iDD/esMU02TlvemnNZ1rikibDYr7GBbbk
xJISBjZvQ1aznvfYEd9ZUg6e8ZIjrFdvwfmattMJ1ZBEYlvUz0nUIoZhivlf
H48SUtz5NcnA4DrhyLOuEd/aGxn3r8QuDYocuJKjxd71RrOBitPYZUlXrhWn
SUWXAv8nkyVws1YWd301AyQEVxOr/TNJ9CMitUZ3AzCWF1lYM7eTS4s/8a8R
AcCSXB6T35BSDg2goYlCRG3A6jEuXpCxyPZ9/rltWEVxR/gP2w3PmXop0oSt
oMoVLajtqo0Cr1Pmga7yhXUBG0mWXzbmbpNPXs48UudhH5zMiayjmAqXBrWp
g1L7xu9dIj4nfco1Wvc0hsgGzDfY8LGwsw6LtxwWYuQW02YtnU3e5oTxesh7
BYk7ApKT2OAetyidH7K5gWiS+2FUUhSAlnf0RZX7nsrmR0E3AVZxdk5DZCVa
ZCYnqSVE9KIbo+ExWq+PixOuwITBhA39nl360jDXcLUfdru5fC86hOTDfr/1
vX2e83lkhiIQ6G2rBfcZ9BGtYsL5adn2zRMKxXcBPT8if4VN0RaJrS6H/CpL
k5kyBL2/RzxA+FELmFlmg0WT14xQxeuQpI2xkHPBHyrXnJbLj7vFbcu4q6sD
X2QUEAmNPTJil3a3iq8aWoteHNAvFmiQZb6/6gZfCB35rdnSHkg7xhtPL+tt
pt/v7/wnaTEWXgyegb4w74wiaQZ51xivtqrhgv6CJAQijKnWg8f9QSbRRDU0
/ExShy64nIVgJzaeKwKykhBgsv4lnrz36zF0zUZLjMOrGQnfBJ/+OWDvtcsJ
IeTiww35qoSOlQ9h/srN0afe2zGWl/JOoZFmjXNBJDHpSrvWFu0H7f9xpDhG
KsO4/Kd6Ufcy6vSNARV4+1BGvNGDkr6wDCC0XyxrI+ujiUYCSWF32s3AhBRw
mzZ9CSFndSa3Rza9MgigZN/3A2DQG0s8HUJfRdA6yVFF4y9gbyvZIg2EU6hB
/BJ2LFX5+l2/yqwM2dmZtnN5eJL7ZlpOadYOedgMixloJH3Y/MauwlK0JHoJ
XCb+FWKpl+jYWdW0dlIyZAXoS0ksHt9aIHdNy90KTgfM5pSG+y/x9tVraTal
1tOwtLtyIQZ6MeLW+Iw7sY7rxJJ5qnq50mNaYiEIV47PkGuAy3gcj1xNXpcg
nXYhXQ8Ab815es1kHg2x75Rq2Szug1gQ+5SCl9JAF1eUebsGIFYz3aIhg0P/
qp2ynnzA/YZlDdEyZXoHAFWW6ww3uYiJJqXmPbdapCTXKmCBNxznXk99w/qS
Fi+7qLf0KFnK2xPrHE1fvOoz/Jd0DROUVOEKvkpvuL4nKuJbvCNX4ytnGZvt
s1XLpKJjfr4z4b9jFf9DjvZoPoFdKM43uISm1QT6yuv87pMHrr4acrXVcSTE
AM33Xn5c1Tw/QY2WqP5EAw5gZiS6KSckK4oCNrkgtVpVd+NWoWzb2q9jjXhX
XGH4TnrZs1Dk9TMA/w5L9DmToptNHLQxycrCChFxJVEh00uL5bxWdCCRmUTb
kPBMGozn+6gmJvbvpXtdUN8CP3QX/1DWtDjM/Su3xyYA4tdVC3SlLLDt2xkU
l43jSF4UkwXFt11TrQfG4/qh1Cra3FvWyQaLMsXCMd6KyrO2eNcs8Q6xa+AY
9UgloNOWQ1NT31S9LtJROhunV81irs6KOFhFenyWqGxi+zNjiBiZPZdOTjVt
ed5aPowiKdbMbFaTdk2jaXnskWu+wjhH8Oock2M8X9a80RfQLYpbuxraGImy
gzZAiPVMsApTQ8Q+tsSG0iMuV7CfIIlQdxsRUVBbqyiO8n4z7TqEudwW3gnY
Qh1VWepJOSUqapVH6b46/dQo8XDKtdsAsDzSeJ5a8opH0uomrDDakAGL/uVl
fJpTwx2FYxdOStnMuePEOwH2/7G+CO1WBwe10upEThKR2/uLk44AVXAqhhjd
l2uMA6URv6DDD4ZYMztC7Y+OnoKvgVkrPE4Diig9CteW583gSwer9d5TCCLO
W5qFd582ZIZEPjFYuT4pC4wGqWkD+2dwKcmczroR6JZJIBcCNprb4U3VdTxK
QBoixjwuPU9IdyEN5YF1SVVycY0nI+4o/oXkUgKzgTrrUnsdIJ4UrTMZusz7
0Y9bgwVvIgS3FAUVBh/ltIW28a53xgD0kmi2l3kkS0/CZo3qDcVhp8zCO/kY
oP/NzPhFtt9NSwrR78pgaZyqxAjszpVJk5zg3LsoSjKUmOrAbGtrhdnzJ6ii
fgYItwVzMuxRcbnOInHFeMbcoVuSwXae00k063oku3csaiA1ksyXfaRzi/5V
98upiBpvJiLWMQCVm/th7wrZmuoVeMRg2bND0A0mw+N+2thr5yUOh2Dc0laC
g70D4CWzObZL/uZ1pcJpGHp/rZxEiEk4thVZ6Qjw1XmZZAx48kjE7lx0HO8v
Cfd2iNCa9Lo8FeKrzz9xdh37+ClOclCZg6jbZhjDQPSie7Q1fdRk+s3aERxR
NkeFDL+NH2/pr+RL0TK24NuFBC//ZDbeUm59AAujWNPfUL14scfcX5laX5PN
ENEngxfPKbINMClczXaR+lbZhNI+iu6K7amoTO0SnjNpB9uqFjw40XyNNCrT
yVXIvkvVXyqGYp/qd3kFt2iqeJC0/c1VwdvPkK/QNN9rjpe0uF2JwBZ9rZiQ
yuXksYkiD79AJqEqB5LPhUlGICDCo1m4Uh5DlDz+dw9RyrzHOVbCywypgB/C
PXEs9Miw4tde7EASZIVgN7TaKW+rFDeBacSiCW/7uJrjT6l643bDCRuM4gGi
CEc8HvpTbRBMpevcuE20Ln0eNWNfS/XNx0b2G9MQ12hqjfDy0OzAAd4ngLNY
mu21urbEzd8iBmqIim8ZnJw13HXNEy54omSlYz83avT24f9EOUPPFot/QccF
SmtUk6CoQPihls6MobL4DL9ghRA2luiAyl8DNXUaTEvPG/Bb2MCnqcDzkNLg
XV/1wmGvlUvfnXzcknNBatRyhBkyTlZGaJ8CI+rUqNn2QvkuQlIcFJd12m9k
7vozrry04M1epb01wY4XjDKmsu24XeuPqX1ZSikuBaFND4Z9aErCBd0J9ZaC
WD1KhV+GwXZIM7D59xmVa0sBao7r72SymZYWsQVV8VlBMCHhl7fWp9laRnMz
IBPBDWNhfi1MExK6d9wsxWO8IPK2a7pLPy1mjpTO4Dx7I97/BxPaDDseGkYQ
uw5kb7RLDRDXL92XiKZey5kfQRfBSpFrfmspalFl1r+tqgoTh0YKFBd4LI0O
ZiAJ9fmWbx7X9bu0e5PoppcyMNWli4mxUtGalcZr9RYZczjfmyDIzZcMpWtq
hraYfQmwdss8IpYUwvHVPGNgGU1PzwAcIY+OzDMPEuvvucXIizsq91H7OH5p
d/MGws5bOBhbM2lO+yCMBJa9k2dbUVACo+pljUbehLxZ6caiRDok71mIs++s
q8vub5oHgPDtznJpaeqxdXv7Z4gonMr+NjIDpO6VT7goGTRkY5t0eX3RCfAL
E7XngDWkZWDQ5f6B9mjnjxNSPeUlkxI3rjru9gAn42blDg+sgwqEnpgjjLAh
eLtIHcreS5qoqLlDnWXWy/sYBPAeXckpgJCy+owGkZweT0lmgYArYrw0gyiH
b4qqs03aTjeRdrlbqVyPldIMnIBKnpUeZrJ0DMv6+kz7LhfreL5qii9g+OxR
5qhR8h8BNI6n4TF5NhUnBeMbdsA4aIykClHJfThQPwQfl8ub9eYmIRyXi6Ar
liOSBnhRTFXSb3ldGzMJ7vktAxdguipJ+4hIr4PxaiL2PQgxS2ittvW8j+ca
4PyIDw3R1uI9iTLmnUWcsK0eRa8aa6R1A9cypKKUKAdt8PPYuprVutULEVtp
w1mRBFLK4J/4aFpIXs/CHhG9yanrx0ycee1QRczqoKhyImOT/QnuCYs+uL4p
xjMCNEjoVfwQ6tx/9gMV0s3uwYgDmzjx+WD9M/JD1smp4TZ1TqIUqiXcUBFh
2xGmvuW9YWipUfT9213E/sS40bGWbAtnugozbGoLDo4pSYkeOI4sgxwsVmjF
p82s0VA7hPPH/6iY3g/XeD/SJCIWpOJaC2Ily8qFuatSgGAndTNvVljgsWh9
tgoRmGbERAcGkCEi5SUyY0W9dDDgSkGpQo+6xTKNMMBC/weg5sCt/ycy4d/v
mlXJ+gjB8IHhEwJCi/b+aSE38ahs9e5LV2bwk3OndvYrKCbalbfWTg4GHSaj
cKXSn/0sawjuLJGEn8C/PAx4ivjkEU1GI0zj/wvR8hEoh82OBJVSWVBH3ppB
beLlUEWRgwsTShIdNi26/zCMOS8rYDpVNNSbU0rJSQhpX4RXkvFd+ZSosIlX
et/NlOXTmOj6NJDlZk6ZBc8jEWqsBEH/Wt6oJCKpBRXkWDfpLZVJ1r8tfcd+
tYlrnBNkdYg0Fw7FBVNvWhnccGEZ2jbqTXH7erEBt9yAEcUKV+OE5bHPuN7J
JaFWGJf5Gcvh06tTbz1t/zAYrFhrM0jfTHS6P3lGrLJYUhwI8HapfEdhKgDJ
qcS+oP0z2F2YdljXB2QdMmJXK/XX5NHknf60hIdjBerlp1X4PHoYKpkIQbXp
2K6k9d794uhQ1IXlmAF8HRMTOoDvdELnp0/VXrdNLgNq/tOl/tFp4xV/vro8
zAv2wMTTr62rI+o1qqYjkuxq2XcQSZiEQRBzE5g9B5DhMjh800MpSbCeEjmR
fT01nIFBRNbsUNFqEKCTP66CyOq5xOBp19P7gyGEPfCAKhvnPBpBOYvAGjcH
OICh/4WlgSXe4JgnEzSLFVL/lyz5jYRlG5AMMblJXBs5zyLcHOoHquVfJWyb
sSXJpA+0NIgDNkHKx8FisLvn+TapfJXiC18qBZM3XgPQh2iz6wM9AQd055JS
d7SKg0NnkEZAfmuBZ4+AbnfQOg0QBV6gudQTMY0oHyxaF/NIyBTcL+w0hlGo
IXRrxNTbrqDqrvKXk7E4VQsL+mtNRWalApE7G+UpFOVUOt99D4GP9483mE1R
l+jIflxVSATaUgzoMsJAH6weYI2ygxJr3oaz1RwbH0Z22wvJ5lQmIIhxlsVt
dMUp9Rv7fOxmqQtjA7lraEr170+Le/1xl1RMHEDKtQ2i39W/Y3XxoKpal5xh
7bCc/XYYK1JLynrHBb31qPCCFcDMbMBe9eynwPazcGNJ6rTTekW4Ve9dPwh1
sv8QzBDuui6aGPBTRlqxYhPcWIoopkFWdJYChv7PwqDEmhH0HisUUe2HCMen
LWdljAV3A+ueJIf7MpuMHdhwkaQjwrwNcKo5cLwYUa6EWdw5Zr+ezYWIzd1y
saC2ffZPUxtwg27bxiHfkNIiK6d2+FaDZOY6RHGWKMFoS9qO8jCRW7jS++eE
8I7Z43yMaW1sOefkRICQKWudnfGuK4gGg8W1EGAoD/YYbG8NT+JdOqHPtAYP
1cRjfzNP3Ifv2XjrFjvh6r4Ld8d6mStCKH4QoZXUi8XquQBvYIRfz+ZmH4xM
0ZR8K+PAtDG4Mno+Dprq+16sYzlkBKy7ZbhUb9c7yq4u9d6+LtnA01aDaA1c
qOe+srTsVdm1unhgF3lY/xAXA6rT3ir2WZo0BFPBe+Ypihut0j2MsbEfNRTI
hrfM0wGRwEAuAujGiyM5vur2SePXswl9dMIsVScADsRmSD13ALi0C+e6/odE
sblfv6b9j9McG015xAyBeHfowObVXpw+OHqGrqjFfCffE/GG3pMIXTUCJOyU
BuN6nrJ/d5XFqazfneAAdRCM6yibsoZtzr5VK1JrYKnRcflrHJTF0rf774pH
aUFapDE3lTpjgWoIg7ZE11rkz/cWDqTwEZxMUesSrT+e7HRQvtWXK9IBtYoS
PGAM279BMHZ6IMYz151PV/zR6fCmAhniYG8VFDKU4N996wNe3Sgmta0jsps2
iKsEPNI+mzGqF0WEZgW3zonphfiQtbB+lQop2ynt3WQY3V1qmY8WnTgH5zR6
/D8x8O7gyz0QZqT59KWdqFfDkTnCmcl/AxQdD05KDBgONPf+boq3gNYl2E1V
7pNRPgbVig7eIUQUzitDyIUL8AUexUCt0Nb0w7mYHkhSL87FywS9TEz3GGLA
eBiJbkIuKm9HgrIVrJ+jgMVmqLcDZ2i+OrIVVD4ASXVtFBantMQXDHjH9Bl/
YOVT11vsVDnX2NxR8lp+Z7wLh3H0CWV5kNGL2nWtsB3aj8amRlrQP2V7ZlhM
tNEM2nm6ig+ipb+w/MLhXp24o4RJIfC+ZswmyZrbqVTWUjvxgarzKW/xNyrb
EYXlhTqxQx8QRdvmIjXGKPE3WVLEJhhGt7eaD9ph/UDcOgf4sUrALsxZdG+J
bPEEwQT6bGap5cgzFIt7Vh9B5GeCuOiTUIjHuCc9Lf/yRgjuB9wRnLDLiZOb
iNk+mbiJ/D01fX0GXw4GkYXlN82lcW8gMjXsHh8uQL7f4icFQGUPbkyP2Rz9
zBKXRk7Vz+vu4U9+yvhyvrf8RXFqxJ8GwI8IofzLGuJAYNNq0NNpLBBi8vNI
9iKDmZASqelqhTCehFM/h8xVnNiwC6afu2umwECQEugQMXnlZSoHuxUSxKEb
lj7CvNUVSiVTxmdI8k4Q5iIefTyF/xli9uyTYZ9XMxjtiiJuJqiFfCt91TCt
0gNygSQqeI7CWxTEPSBqkVGcqX4bfPZ2S6PD4RUHmrYCLPZHXjGtdWM0zrUq
pm+9MLWdnivtawA57P9hdfLKFrOoxj4pQFpVvFakXoUX/Sf1FwYeLS/0rEGb
dpIj0JjT4+x7Ae8JdFNWsknoexJ6NfjnMovhrdcW7yxB+LTTmCX7JxhxM3P9
L054Z8kg70mJCMN/jaIQxJBXB6Xs6eIlzRxOsZxdqVkrw9L3BB3mpfHyISty
FuwEB6bVHaksKNxIjQI7VNACQziLinbjv8rTnLofn5yxfQUzpUx4CURPtClP
Lh/E5JgTb07dz+PQh7hLAthB4X6nU+KDkNqODVPwoM/fweRamkCF6Wb6N3KU
I0mhQiZjjSr623TP26mTDHlkM1FoJTlk1KAicqoerF19ciqI3GSrySyGjl89
Mxl9+nP9HoIjLvhRO13fQmG9y3Vpg1ORC702bNUZ3N8lTY2uYGvYICkIHqdy
99BTMaQxHjHC+gB1k6321SngIAZBUE8qWz3B5jQtVLvH/KAv5RdU4EELCpqy
2kO1VIntYIn42d6LJ7JGLYyDPTd7gVgUXufmGvOA04kmz2YHfyLmiLh6nQj9
LunjbigFWPJiQiISLgzogrZ2ALgRVLVYpWyzYFKjfcOGnIXLvMtW2K5D4/Px
r7xg8N0o49rSoS1G5rqr/CH+FF4qa59GtDDe1dRpC0l8y4q9TQw+2ymr3YO4
U30O7pKNGWM+la5kG0zHAh6ljPYwYqhPQnvF5LvboEToSHmANbWIxaJF1SLS
xwxkewaJto//FTuCxKn4sonokhNYyoHIavId83rT2SXJmFwyMCWGDYrh3F5s
C/BKQ7x3V80BUOAdsDzoVovATpHId8DUItdeCTJUGiGHlyR4PEOiPmCMKNr7
sV8Kf6UV1f4gQM6OPC/9jJoetzgvWWuRe2tZeEBj4nnXCj+G8Icj8FMktu3T
PhBC/xK3kOzJZu0sufhkHFSzk+g/7QennI7N9x6aovqattiQKK7WNqtbuAiu
A1itJSt1Rm4yiwx0nMLt0ATZZUdfDp1NJqzRnqfASEZtrWu1xKRRxuIdLLv5
CVlJTiwgYWjPOBu9a7ewWjIEyjcuiXaEhG4InMy8wtmSRMnbz/FayrYL2frj
FngpbcLGZ/chlMY/KY6fk+r8x0A6RZjb6sz0QfHfTWxy+Rel+2/DsSV9uHah
9UvNnQsADhEOVg2s0ag5pw60xylpV3rOcqaRnhVaxV2miUjRkPE1xJUQ0E55
2wquywww4LTE/CA3yL7vf2342fkvAXckZ5vUQ4kZ4eru8LoadvfPMWdF6rwL
tI1Ik7ZlyOZ0ToLaw8jO75A8IeBUGVfTkvstNqF6LOaUNkmdK0poKZFwTyh3
7iryOF0Cn7qiDAQf5qhxCMvna9XTdiqJN4Od54zKC8HHXBg9Zzew+VwJFj3K
utvHrVGAQIcfZpWVBTwq1ZIp4yGDSdiPBw4P565fh15b5MGF57RB9GQhsZM4
hqQ6fJEGl/5YIkic5L6ClkJK7a4OmSPYHwc0N1jtdx6+Q3irwcni58xwD04x
8w9BuxDHn9ojrSV59p5RhhYOCzoTxcYTkpo14E+Kp5N8lF9MjrwWoQY31c9I
2uQmfNoUR2xnb/cehsp/FhIIYWC0owVhuoMUMagX6DlJ+MyBDxo4CMgzME3b
Wtr2jZt0s2V3nw72PBPxI2vtiBgzsKuR/doIKVCco6WSsrHFdWTrgv9Rek7V
06M/bQwsYt32ed0Pgq5CYrjiyDnznc0BxGfBOzaItpc6eDsOrTVQDYbH0Vf+
Qq8t3mWMzlmU/cOIpgP+C8NKwscgLaj0RcmgoTeYF2SanA4dUU9FcGrQWZyy
peTkHTbUZ9rd9Fr2kMslk1JU0V8SChADzCu8Ccatl3j4+2+V6Dr5fkfzTVi0
uu/+41uJxVsJ1SZnnoe+fLRzD2xMDDWCgxTavVVd3L51UgU4vm8HS14BaVGI
KuWFbvcQAAQtjNXM63gWjCxGq6mg+QH0fMIPLB2wS23RaVJq99OMDWZ2DXec
DiUf/6eankOCtaGBFX4KVJ9w/ZT38J6I1wsU6KMDJLWxlWHksOiQFoPCUcgI
Rhw3C6SZAV9BB4c3EKaVaqqNsr8jZhqlzTzubykccvYoivc31O+58WRMgMGz
YPCZKZG5TpZ9LkdZRWgnemKTXZAtE/B1ibFo4uLs34xMl6jRDrmXmYiLgR8f
IZEmWI/NHol8DaZdGcXyZLoyP62xCjd9wemz2w6zYjHog4dzqfR2UN+bcmWD
K9wYLiWZylYF00caAWq9pGUasSt6Ciri5u325/ohLzDwXM/6qTL3uiGx+4M/
RAIJGAW6onJCRvAc8AfYpkGoO1UCR0/wDY1Aqvn06Hmzl9QoLO+JX+ZSQsoa
5gH+FIROo/n27DPjDB8sHN8xkVBpphjVRked/qMVRFPPzNm/gDubh2nBR6bL
utD8iUf9HiGt2HLai/wtfeW5cNRqWzXBDlxeta4bInglkYa0cYKH/DZQ/qdo
frfCRySZH935wMcOAS2rMf8GXB7TFLTqzgaJ9IqS21Etuv6YSJh/rhj3XV0k
omNrRf8UyDMsLmPEfv/1BlRo7COTvyNl+DlwOf3mU+im4xyvCyCT1auRoatv
l6NomD4JWWN9jKzQJ/0zEdJI/r17lpiiQ/Lc32H9VxLfeivq1PUubo67iR68
BXHHuOKDOJtv2z1fwPvhlTEaIPp/M6ozfVioQiK3mbXih86NyI7HxbLc4odb
rU25T0Du38cdADBadB+JazRpYz/pZj0cpEgsKYvoS3wIr52YanL1672CZRmt
P0k/ocwF0It2mPkhLo/DgKDqA+XxSpwW0k3lHLH3CSNXEaArOffSJ6av1+d2
IEGEsHWKL7YUzS2lbWRKZ+Eow2ZtTJsH9gPa6OabH4tL0hracvBCqi7kKnpV
jXaoaI91d0V4D+E3zOxWskTM3CY0+7BpqDyMRnlngPdBR7uchJYrvHppTGal
Vo3qEtSzEMrDLqvHuZTh9sOWiU1Z3RKGs62y6eOnkWG9RfgyX6SJKgbW+nVb
N3KSuNmU0YWbXiB5a52OjqKPCGkokMEMiRNYdw5C3qdZuXRy3vwL1rzuXV+O
MXdu0LujvT9kj+SCQ2TFJSLGbsS33vCwTUKebl7dJojVh+tBPMZFJPOkNiPp
Fnxcz68SXGKMsiYeS8xvKWcttyN3IIUMqhT4PytQ+oNudgV1LoiUgz0c8SRO
hT4/EpMdH4kLkgeHABb5OkbdY8C3HfBkhYunScH5dWIxXMjAOdJBEDgrLkiB
HwUKEgBmdbLnUB0fnL3noAyDHvGE6qQiy2jvnNE2yhpDW8Bt/b4BMeoKsYnB
M7oODRhIu9bz4r7RrFVAB9jITihwsKinzHrqY+lJYtYXruzxR7XxsfRpcZeA
4b05yy1clEByRaVYdpTdSsJXCpYsRvf519bjJ/3Tr1nEK2RYrDclop9S8Lbe
NGVj4gp7iJCvXlCXQGPip8dqxFx/SKzP+zVm8+BRMSk8qwmPVzGIBnf4aRZf
1i1q+IfRLdeUbIVJbd+UMkAE7lcShl3tf6qF0dfALiVqOR6abvp79E2o2ZyZ
eo/hTIaE6uKgLyV9JCNr1xrYGed1oqzuTWFKsS/mT7zgjt3kqqWv6sjm8kD2
mMbW2Bl+0Rj9MHFYStOL7+QOxsXM6Jq62HsuIPl2dJwSohYJ6ry4cwdSAHav
nIQAhkpr2fmTVj4zLqu0i3AxxQO4XLgIwNaynPS6Ch/4RTz34iVNXOKY/2ZA
5ZloZo7hRf04lNG5I2W1af1r7Kwmf2Qh1iGrnpBbCixdjcVIiShLrnKQ9bOM
OfLxPaBWsG/ThjiFPk1Bmh+qXvTJ/LegPNEiy5XF4GwWMXncHfs9wpVzgPIK
eEBFa4WCPoyHadocb7ejMQSMgc5dvHB8WUKqUC/yZOmjoOXjfSw4WxHOOIW4
qn63VEcqn6I99iuRz4BT6+pmbJ6Qfla65+X7yDHB4GeX4St3OigsR+0bu6/R
fVPZlkzWXQKrOoJxD5K+lk2NWdeB1UshAz1JEsdTaUmMl4/eqojQN1jsHuC4
jTWQUFPCLhv/NamGoEBVlSQGMFToSwlkKmJ4hBuzkBHTR+S0JQtKoDs7Po/e
f1szlaHKw7Qje0cgzJluBZbBNjQWcSa5lI1S/2VZxAuWOqNZByeCLTvU7qlW
rQ48ueKUanfk8rCGPV191jL20yHIAc7PM3v6BUAP04huJqGOaj4d71t+P4MK
ftIY9HopKI67hm7ALABAbffwfEyVXdxowyJEKgISz5GZ8ZJTA/OnELEnOzAA
mo0VamtSAokJnQmKYPJ5sDyLBYuWyzG8PYdwXrn0c7D9DUYErumgwbOA1Zq9
7y93iQzEzK4gMM/QcwuzWULUH/dwIbQAoZArGbw+3U/I57oQL7vFUrOl8nsX
lypnunTgU9cPur7jrWYVaeIi3nHzOFxdLotsKKaBghiIjZjkdIDEHiQ+ELXN
wv8IRKUWxLW6YAH1unmEFee5aALc80HvNnlTh8iEd32bBYm8Pjtm6+iwVj5Y
EuNixmlcsn9k5ycyulxoQv/CZ+Q0XY3riqPvjzhRUqdprr+ULJMTmsn8VFc/
/JDzdHU/I9KAhvlwyJ2B39YfuukTc1+T/TtTDFx2G0muHaRjoy0SRAMaEcYe
L612JBLFPaMosRFIWI2dqWDa77Swkq5fQlguSCb2IgU+xlKJo+8TyYA5MFw0
HBM+FOI17BxYuTpdrSswcJyTDBT2bS0TbgaQM1JwOhI6TAJIjF4gLSa9x9Cf
SQ9pGwilWjnju/Xlg+19rO4CG7qzks386X3h1zAaczHH4K1pO/GgwEfx2iIE
WMW+HOJgo4Vg+KNwWv0zOI10GKYd/rIQAEqprbf7SAxDdP9bjrc0FgfMeaBi
DlhpUuVc1i/H/KiVpBnY0FQcaXGEsxmB5gpsfCuOwI7ndAskNKilkAEL2gEm
WU41YELZsD/kCHhEpAAerQWUnSktca92WGGRY08TpxqgZNBMTVqnu/AejkEs
Cd5OH+ToZqnjs9F3AD3D0qkeBLoSFDWpoq1/wcoxc79O5WeHtwZVBSSPP+Ph
orH5Vj9ORP0OZdbYEUE+S1DIsCtEYtIBEPXG8NurO6fg0xpxfp5ND6uRjE7p
kKYQmMf1ckU/0J/ZR1ZuywQeF3qWaLcoq3epG0z6lyp4ke6XjdQXbYJ5v90d
8MxXi9HKCKKr57q27RCoIw46Y1+csOBHvBc3DDkWpGTJFno8nrMdxLzVapKl
+5LB+8o4mrrmxpSBL43Z8YdWqZ9TxUIOHFKgf7pTNwcIJRh8Rgh9w+yDZ1Qj
hxhRISWwYd5YIACn4Phi6Lsw3guBUoVjb2yVtYbgnIb1+JI17Vy0XWEZIGSc
j2EWrjGoqoSs2Tfyhoy9JM9e7IkSc2tvSlOcC1FzfjogaVYzfyIofHlkRwdz
KvzKOpZaU6uI8Wstk38rC8o0x3NbiaBEk3CILRv+0OiuXE3tVxrv8wELy0fN
EoqIbcAte6nY36QGi+Or53lGfDAHXMSxAIzjXLMLFAzt13Wkd5ODufLNoBRK
PVyGfQKSwt7TbHBvmAka44Aro0B3wk1G+DkVi4BOLy/HN8/COxZ4Tuzlom+R
Daqg9bmcEKWjrEgTyBz9jzxs4cn7GG03BthFH0bYBiAdi1ksgWh1c9HugVnm
AtCjplbriqKq6EHq11FgGShVVrfnpsdscYlMxb5anwJQ63xkd7Bv8ivg2EPo
vzgK8fDSpktu0y3u6b5kZoI5JupkfLgeyJSKgTCDb6asvyO1u68N81DxwcQd
aXdMxKERBtBgFM68xZg5fySZhNgqqws+JmUjGj+jmZg+uH2Q9LQvHvtWNVdi
8Y1LWLoNphSNhG6mHJ4jhblK+CTPHEKQ8bdWO96EUYyxn9Z2bv+DqAQwbgv9
yUOdf7RyFCi6Y1T0DDBeddn6N2rOg1NVhWuViXszo5LVS/UlF/tXVsnC1p9q
H0vkWVfSiakG6/6r4TlEWdb9C/gBaeyYDLE+CwXCKm2v9iqmIpAZcHfxm4rv
WCRZNWS7SWXswFizlHJlULqvjg/pNC/H9DJyNCYYMRJx4zRo6o6V5Es26vDN
hR3z/Orl4nBege+TaeDSpPAALjt0cRGf9onjooOk12uTJJ19vRTl8oWrmbMx
5sN7VyzpaC5fD/AIf0CSR/QjvKXxmaRfBOh7KnWGD6Dy2r0Oodj4L8KuEg4g
LOEtxGjD5GBar/a3JH+Bb+QXB9/Sq1Vw/TZ7UTLV0S3q7sNLRD/wXNKqFSMU
KMdwG7XgJkGjlpobLSX/qIuYWAeNN9mXnvk8KLcOYgiUwME2zsNYikWwXBqh
SlTDVIAE9XA7t+AWNwQxfmXEdwObfZC5ZHPZfoiTtieeRydtn08tZUVbkUmT
VyBoT16gtaSsvlNpsxjOmEeJw6/zkfu6PD5Ot4dMGiOagDoi2yQ6YTCYA1AV
wxEC4pAtMTU6ER2jNCUdGVRp9OtuwTdgXbss+BqTcx7/jEGjTTouPa0qIjDT
Pnp6XLcRZ7T8JSYk78Yt/MHrYxnU3s50BAsMJEr6CxurOyFmnwHRCMVF4tJr
vhKRcGoSQSd+M7LU6sdEYA8txwwWc/6qimVKAK4QXsep1cibxL3wPe1E5ve1
WKAyeQ9+mKK8sn+oJ0siHLgc7xGVzHZ5mY3gbMmldyc1ul/7EJqnKPIQrgrF
TW45iS8aHNQE2HgIHtRNpQCKl42eEZOsi4FbdDX586licIn+bbxNPikEIzyQ
oif5VZrNCEPSmz+wYG3OOZAG/N6pQu/kZChRyo2Pv1/EW72Z/RIcj5rq7G4s
w2lZVKOTH2eUx1EKiNarIsuD8/dsIOBaNHh/wIAMRlyBmmQzH84drJiwVWuk
8nM2M0BXVnQ/FxgxusjGP1caolLl8Un5wVjXoQnpsfLqumjtXjO1kRxYZoS/
E1Iqcwm9eXU6yOhVJszKAqOZBd0gwp+2zx/mq3AvnHeBqSYgVmIsV1lKMLP3
9yKJqNf/nNhi0WNxSsjScqaA6PjcKH+UxKsqeetQEr5KJeDcXZGVGoQp0Zty
ZDW3SCdHj1riE6aQeKhw9NwSzFHAOdGB8fbsv6R9hnSjrNaBHDg0obIvFuT6
n3cWcm2C+4GVvvnTHgMoJhC/Gm6LC9KbFdMOTGDkIc4Wazmc6m5AHyVDfdWS
qJY8rckWb+zt1E4MrCe9L2qzAAZJK60c/tmXi7VAFJDMHtG74/bULrffRiem
Fa5+01fddWWlne1OL4myTrGOwbQQ7gv9cEhFfPt0+z3Qm3HLXzsgsfxuyUdU
k2yXqycmOihCbw7//DF7jaleb0qUagMNUX0lJRb09p9DltrJCOdnpeUfGWHZ
hpx7Hly/vxzgupSvI4/uRSI1wMg+SuUmUlw61dzeoTdD4GmnzAAEpDpwE+Tb
3DjNP9F8aGB3rN2/ujAYia8XIELHtWT6uzs0YMJr2e08PfCNNU4iGxWLxy/1
arAMHC32irwjazqG4oNKkgBp8jyIHH0p/bMQ3xFrSFSimgZRPXV2ibhRyWa4
B/I+V4ERB3Qy6sm4u4/+cWKUO4XRm1pKTozQYbdVHdesCd2lnQUD3S2dSyhq
BLB3hOOPgMFpBSw7IBDEEDcrrelLXN0uBHXeOnfokYZ46ydVPObaMfQKW++9
djzOnleRg5WcLB1BrfhqaCVWFLOzzI7NAwLsi2PBoHWaVOq8W56An159eLhR
WXzdZ6RtY85r7F9TVl/PKY3BemNNpWbSYvLIj6lCmbf8shJdYhCZKeD11pVw
96It4YwKlKrYHGSRf3Aq2y6uKycQ1m9FVbQ05RQATUSr/XxkSqqmOduFJRhF
omPwSbV8DLHV/XMKsbo7hGdC/zITGs5xxSbN2MJcTB3SL9vZjo8IxwL7Xook
FkzJk6M4JkLPpddeKoEKhbIXU3z2mDIf2VYC03IFkD/Z580IKMGOt97WEkZ0
llxOgZAW8VQxqu7xKMMzK8tlKMbnNJ7H5098cyIOsxM1/6TaJSAxUjPg/07L
DTkOLGOo4gcWLY+7U7jp5jhzd7RyasCNCeWDTaZwGoCkz9w2Pp9OzNFMGnMY
3siNJjNjFl5D0dIn7n++L97/n/SpkPT0PtcEk4tfiVABKzKyJL6C9lXxTbVG
2rXZ0Z8kNgjPX+walqlzq5MmslqXaSxNqzycDLD15qRvCm1C0GcahLT9o7K7
pK/BwoapdQQALQwmK7Bgv85rEG4Vm7D+NFHXErLJCUOPXkavqDxUP8eCMVQM
Xt2R928jCwRjnAdxzIBfrJT4MKQuwx93TAjb703Q9VTeSXChmR+OKvJcO+sv
xKP5XI8hNndVZJFvxEff4yzeuh/Z5JUvi3IscT6j1wwJY+W+9hYDlMpeOhJ8
i0YID0+lOBfw/l3wIoXCPJm44wFt3SRWIHUPSYmNbw8NmUulDP6X8/ChP9Dj
PYSbptPRzTE+11Ldmo5WIM8UFBVWD0smOFdDq/p2nTlQsd1kkQeApBHO6Tcv
D3HKlI5G3wmQ7WuQ6zz3Q6AAA7bROVn5QnrsjoWQA0pW+MJO2rputLVKiz0/
XMuVNFv+SAberqR3GJc99zEdinNJufg+/MTcNGz1xsqefR6O+H2cug6RN7gs
/mrK1ydDluZPjBWSgbUJkZ6UGaszQxfJRfHsNC3fIjMQf5d33kLYj9wH6Hyy
rsVnOANm17cgjRokImM33g1BwxZ7K9WhsSnvBh9mtPeGx8WOGXv30RUnX1NM
TjcWpxc1OyIt4GSZYUurNBGc3KYq3Yla36V51KWIinpUDm0eivH+gDiAgU8v
yr0dvBJDskvLWp0bIZjnwDS9D0aODRr+M9lQScQQ0AHC57LGIG3FSM2juMOz
uDOsue1B6jOguztqQVYIZ5MCy3ukADxq6503zh6K8/5XDfWd3+JxWcOzD/qa
9u0X32cuNMctLDD3Ui1id/h7RxoeWQh/ocVjMxNEs2nU7cQj++8qE2BtWvat
VLRyzKfE6Fq+o8REdOeYuLDGbDi/3qNVnqFNGIwsL9Lg37IWnYFAAspxFzpg
jTGi/XYAZ6z1b7RiJy28ePsduxdxoY+W8p8o/Pnk5TkCDIdyFpjQhTIZy3YK
i7Lq434Bs+2cUo445yba8iM3sCtQAlrf40lzo18aGi/IoZNQ2fTcEgVWM6Gh
FndPKYW74695I0zBQsftWnCxjaOT1SIQMU2bW8p4tapPM32HcRSmwFESQgc2
0tJkfdWWxCYAPZN3Fh11KgWJFcw0XV/vCpyBTm8HYkecT7q7/4pboM0/aDwo
0+OCKNtJRuqFctJS3V/4tuN5FdWE7heweLJMkQjsS18dRJ6WDRQlBfzXoGC1
WtvUqDV8s3mPZ645yAEc/l/L+Q0O2SjGu07qbMqqTqzUweVLEbSC3aHEEPr+
2dG2TRrsTqFLvkJ9FG+7cD11CebZ3sc9eMZRHW78dJaomyGtAb4re6jnF0/o
gq7q31nvK8TypdkC1Jjt+k+QZZE/Tf9eBSoIG8VP96QyuJbum4+isQgS7N6u
l4A1nCeBK+l+xq+bBeGaCp9fhQSmoYVhNxoXPsQ7lAycteDnG2VQsaiTUcku
bXgMKssZ9ozwD9HdGBKNQooJw3+MAAElGNY7Y+EIngZGwucqj+rxFLQeLCdY
xq/uOD28AGNL+8eA8LPsLut9n+Kit/g1LOHMXIv3f5JPo6tVslJvv2BtxhQG
xnAUJjTXUKbsfiGgipjeVbjS5QS+QRlZDMA/hmwdKq96+XfBjJXGo8k03RS/
yvT0asVV7XY870DyLhRCYMN+FAC7jrBBCiiXJ3ZDRFnyl98UnzcJGG/ADAu/
O1+sssWiYLTXYhNDdhZRo+byJ4Sj0ukOUurmFB8/+vANiPuKMDD0o8ZNdMwO
FR1c7/8Er6gJrddVK9DtwujjyPwaqut5W0dQTFYWwBKME+KwL95G7hXSZCyq
SEKzXPc8+0P1FOsVtgNkYmSZeoNpiqVIwxfpcx3K8F+CUh7v/vxHIGwPIeB6
w12d8lEWobpB78fvHyIQ+nkXxYmIAKTtzq77FxXdEajIzwHD8v5UJQniDruk
7cF/QCFFY1JoN3wU1h4HjQVZcOdd8LRSZdiB6Jhg0AU+/HRaiZcnG+uULFeG
+m1o9Efe0RyJc8v3lF8CaIQAuHVWeIAF2Bd9pmtdtfyZ+Jji5iDnvDZ/oaYm
HMQ24PqLOQxcAhuFFQMJBljKDt2o4l1yrxB68amfWlqBCQdHNPqxrp0IJJ41
xYl8hguQTQUqmokfy+CkhhIVk53h4cys0PbGduL7DB8XPAvC77w5BFg512VG
UZpEEQAvpuAzXJlP1zpD3+d3OXs63R1oq+mDtVnLAJSjS4msXp3xPCoOsDkK
U/yavcVadxbtzHLQ3KhYzZJtYtU7Pzhh52GmfVJI5AKt3CDd0keP/xDWiGc3
TMDcQ7pF3Q2clZP6HMoOnRiihrLZN9SqyVbCRJE8IeX6Ajwa4sG6f38SsI0N
txlZ5zoQsFvB+sty95yJs4VOhhId9tQdbErWl936Yovuhaw4FUDfErRT4k+A
X8iVOoH1kIxE5ZnWqn5a3o0cjZE+rXM5JnJQ4ZJa4hV5tgWaSMRYUCInHuzj
r6MxtJ0w0I0a8o46VP+1U1Vcf4UXZcZfVONldWNRm6jFZSaOGpZ15/1ubwaa
aT3MikpPZ/JeOOjthgNYflJ6A855XB7CUyuUwZiN3HfJafYdFNobjTlhneYn
lno1/adKoWlSaH2JEFsnwPksBm4vgBc/OlDi2a18xHuvJRi2Ahx/NUX3J+t2
jOxXiKAMY9EzMG/gPNrsV+U+UYtzvX+eCLhl3i+2EC6Tzxp1P/lfaI5CndPD
/FCH2X5IrqTi3vzt8WGC3OW+rbmL5t9lCYdGw19e6GoyHRn7dotg+TPdPgnf
YEKZ1vc5aA/hm7jXm5o5gcAz5cgAYy2KBOluMSAmK2pvfkUtyEJLHA9XLJcH
LHsv01Sgk5daBpjF+KhJQAqUc2GEF8NlGPBtLKO0qcXDAeMZZS3X/lVOMNCn
gjUSGU7TMfnNdKqAUTBKpmP8f+/8Z3EsgFxZyuPLV2FmOyEKK0B9CDkMiA2t
5eq65SnPuyWJ772WkwPOD28o76LsTOC9LdQSM4BAZIfX2CsfZ1ifFyLxsEuK
FG4Ny4CIVynYSHl/ItGJ0fwvjkNdoz7eUUuqYRztrmQc2OF7d8/3skcduw7b
+BGsWmVw7N6he26Il6CApH8NeNUff36+3ZKF/o3cxPG/Kh9tJ/4PSOFDJg0V
0CgKhjT6KONpIYOk9sp/HV7GT9Jg8SQ1gWcXLvdDX3ByGLF3IyXDIB6rdnXX
moNRstTC4lPDDRxIUIiBc4fV9p8ZO04xo2LiSmVLaL/tsT1kkT7Nl+N5KgLv
maBM+3TGW+yn3E2fsAh/+MwyCsrh7EgHL3bDjbGnPk/ZACe2n6UJpTSIiG6e
7yJ1Tli7DQNUR8yC/QCg7r0lVOUatrUuN/aWZEOVZT3GklZpcEtoamlS06zK
g+0PYYPw62PGmRq6BEl4AXLH4BkKy2T+dMm7T/HhH4fmsN616dAcJU394AR8
YnpLKwJkzExoiwd7sjlV8LjEOlYYHBi24I4lLk2FpG9zx2N+gc0IY+xzqA2p
9wwKEa0g1GkEz5K+bCJt1FW4eUBMkVBdC4b1pOjsfdmdAaVbAM4NuED6x7Kc
rodHTKJJbzkMQQkl+kvxYsmtv1kDrnNQT5RU384hUy39UAy6VATk55FPIta1
DxPn8BWfEOdp0fmltuLwRgvaTUxIIQa0f2tnyvlr4UlCGz9ZgXqktpC3crCV
xSPz+OJYVLfUtxABQWTCyNX56dWkJio/fp9N1CIRsf6G//r0YX92N0AeJZzk
bJIDDaeyjZS9NzGKnQMo5GyDicPkW7DVr00BqapDwz7cifXmEwBOtdQvV8nF
Jw02C1aALprEOWcO5UZoijXaqbZyd26BKO+BBfunnqfycrAShrLmdcdwUv/e
oPqULsjWc2hTFwKXWmMutou22a7mpseYgxmOGCu3iOI/stlVDrA3jUebLfw+
9ThDYOZo9R8m9ZuGKogUVS3LupRZCPx5dTCXpp3rkxss/WMRsCZRIUjGxxRn
QRKwItbgAvZGjrTcYsA+1WJNEKBovBthMqb3abqVbz5wDvrxF9X2NMTlz2OB
hryKMZvZPzwmt+HRmRxQP8FAly4T3LbgdOPxgzlhH9DJY2pks5L4PLWNL9/8
2g/FCjj7fmv+M+SVLYPhuNdPzKOW3LW5y5dFpRBZvJ37d1tQ8yFmRSlBCdGj
4Szqzfsat6I3jT/+LNoYjg/sRjpWeirwqpZwQmS4Bvqx5Vst4jWB7upm2v0U
bvJl8ErLrUTaPmtuuWWiA088cHWJneS9Ca/y+0BsIjlHF2FjA7W9AzYFQAb2
20yAXx9QzjB90znFaT1o8xgS3quYDoiGqef9DdRlahM4FYCjD0MfZibG//p+
srROA1HONda89ytNbgW4KOosD+A1OUYOn9C+xruRO4sdH0h7W+qObbvJ2oTl
MLV/ZVKO/7vGXH85+mJ4OXE7jCKaZoLj6Zw7g8hi14gVcWbndeYTZQmTe5JF
Y1LS7n/CLYLqeseHHttDYuN2As4L064mvFh86DrxW873v7T4yhG5nfQOvhzE
HZmx2bDw2Ok7oHkMZuu+cAxDYacvCryI1mfJoxa2GhfoAyJnVUett75BLQIC
84t50WAaP7BkpIq3j1kx9ODy0e734fpwBu07QbB3Lh7DmcvE8g+6P4I9fyge
JSPfmgDcM/WzYMRZlGjw0Y3BTBPd+TGaWe8yMjgjAxhqS8FndQj4yK0hR6+U
qgV5G9DQtLtz5WSejB/dfJ0eiGG2kv5u7hijExg3W4usxoo6PvVkwOhWHhnl
jcUVVu2GCcmAHBdcT2JCVhsdAVfS9kyNfdR+wD8zVrNj6Rh3bWq5YYYz66X3
bXW/XBQAOFQM9FpVYvbIod8t+s+X6uft3vBc4sPaPotjJ3aXb3pHhdbFDhgh
bFbrt0IXmK2aGjo7xQW/nPlYHMNhASRgmZSp/yfYi58k3eTJSGNB+S83Xzt2
8Q5P3PoyfnofR4Rl1H5j9n6Hyx3ozPnKlphqpmi7La039Xjo85JUNARctcZw
VrCeJ1xAFOT17cTtPuRFthFv+dw/EJkhjabg0v40DUDymbVphCkVcG6fVlov
hhS5lmJiZrssx+RoTPeLQ7rQrui48il4bt3pGqkkqhNy7pGzFK6HvSgrSwsw
T+MZtqlUuyGl1YxVmgjmQMG6jtNTlwJVqPLas6DF8GZ9clKBS1Gg1i/CeK6F
mnIE2/nzMDqNhBTTu9Iy93JndxV9KvUOJoh78OMGbaSjb0K5TU5Mm9dtTJ/0
MvDmMmhiXvhBHESEPpctUpaOn9M4J2xpznPNj7fsgN31ngT9WJ5jE1vw0gfB
ChbIdeBOFnkF3p4/Z+fCvz3ojbutFgpdOSWnBRmB3VricmbOzFQPr8UsRB1r
vVsB17d8EjhNZUToUQ6OT5UsUkHfszzlk1DLNPZTIuOxHlZF35YQ+HWUrRc8
nirlssbAgvTToJ8YTmU1Ay8bnfjiUNbJzxJM0Zjbaztq2X+FmDsMnR99WJCi
FPIpHCrS7RbXcRuFK494KHHQO/ExfusCr1+wY07+Sy/jRUV9bCOf05kE2dXU
zhpPhfq/d1Ns9bz14viqbbzNjJURsq9istEX72C/opor/NHAXYJJyGQnu+lI
5S+oVb9cG5lvH17fION4Yjf7bQYx3BR9YGoFsei6rqcMQ6KBA1ITArDKIdmy
zc28mHOHbPGyGgxKL96zWz90vn/BLlnErkxqMQjlfnWgvaacydwpCpWsSfL6
7f7VyOKoV5dZv3d38W/4tY15tdvExnNn4RsiIjj6olbh4bUvCBu5rkW2LyNG
mUtvUvEblQzA294/ffuf+lHtX4g+BpaSoOOhet2XNUR+QbXy8Qod9BiZj6Bh
N1mvN+uKNK63dKJZ2lC2qY9BFE9Bcwmx/QaZS80CZYYcUw4u3nUK5gbQIIFT
/juZhUsymnj9a3VAHekBjltv9xzCmJTJ8ovMAQujBTPn7/V801Nj52Arg3lP
Fv4iqf5fsZQD7MyZ/l+lprbeR5/UPdxX3Q+s0Bb6IILbXMaAb5zt9VGj7+PG
8n7UzSsIQuLB4db08VhgFQvoY+cxWFVkAEWj9xr+clyoHpiRfn84kFSqzYVP
f41e0CavfPtxZQkT5xq6jcgCTiIgW66oELt+ir0VoauA/XMor7k1KOS2iEn1
VRHaWPy7z/pkx+m+8p8A6vMUtPjyohAEaqQWckzsDCnIRUHgLsDYn8cmpnXh
qMkPEVkeV4hqLawLR6VnLWzte2qcywNrBEZTLJxMTm1ZX6EaECKBW9a5PqzY
Yv9e2HeRexPzFHCQzX1OpM8g5lTL939qYcsLidSzu+fAt9ifSZhQn/cNbukp
OnxILqfrmzO7PDesdGQIyD/T7eBAL/4cNva7ett+ME6o8BhFkQwuAWl0yQQJ
FjW4OgAl2buK1LVPHcGwLMmGs5N0lTcFCNo9sJIAO089JNqGoC2CDcc9Hn30
8jrHrHN2bEqrKue+7KIYRE8kpeQeUheLy3B4nE1jv/7nrNEyu512vXMh91Qr
5VGkkl8ZCQFtZm06Tu7LtKcBdgkrej2jY7xuR0m4lXvf8W0jKoJUQYwPjMK9
XFpLooVULwh3oGvUHL1jxtydtg9h5ujuMS2G6mW0YUDVlz82AgFSD8QeMtwl
visPthRDLQFFlNNj9MvIqLrDSm0+aNFQOv/QxELwqGz0Zqb8rQp6ZQkZ5XpK
WdYtmtXUggv76joSUUNdNJjScJhDM1bUwnaO7U3csB71WcgtRBXVSEHHBeNN
nCDFSzlv6OjTx+SIQuZ2S6VPhGsD3ctK4nyTga3SyPd0le8tkmTBFgT0DD/i
81tJfAfSYfNIMms9UIBHaJzcq0MJZllYDxCxojrB5TWHA0gOO1gEqDFAUc84
UEANgDRPwsubDQrUEzRW/+e4hW8MkAkv0aLnN0sjh1R19iG5IBSMILzE/IZl
gOGlGFL/SzYgSOekB3o2yBDziqN1qMfMJiq3stYGDF5Tc3an7lBhSyGCpAGD
LKDGibDCHheN0Lo8oQWT5s6dnlGmLb/wJYIP4QrU+QUXNBuJuu5p5GTN9Vsk
LnGx5Qlugjkz1VkxgfMyFQcK/ogwfYSLsAEcoUdxkaI8FmLRMURtoYwtCa05
B/FIbdwfvfw5sG04vCt2lR76ADnjXkUzi0eLCNcJLxXqdNxTUYCt8e81TV2Q
0pOhFyJtn2gSM9T2GP97VyYq2zsFfWouF4lodntYUhtYC9leV4qACz8ItVxM
vGautlAqVyCFuJqGD5JaFuReELgSFipo1PxPqFXiYRGv7b+Ct12xkFsqPq7f
Q3Y9BQeq1oSCgQKCRE/T4pH1wJ/86XKYb/z6VTz+F5tRb53/8wMCSmRmccoH
jfRnhDLT6HhO/RnKW12wOTqLtI4mB7FElobSWnqE0oVStovhNeiFbSj9v5Xs
Ndo7ZyGnlCtDLZ2CuB9RT9AeQv/V/SkBqNeDm8M3H1Zb5oUcq9eWNbkaHJPa
XFxS0j0XQ9DyZQzahMEgZlmprptsVzcYo8zHfEGqQEED0b8Zua2TmIIKZ/GQ
sbBmRq9v/TRxdxLryZTI21NSc1NCg+NKDfcA+kLG/QnVOPuiHnMAmqZMuNlg
a2etF1nj8+jb+MlHuIITrkXH+YwwNJYK1lrLjQiacyPPQyYqMTFVQ4zZHIjj
yG1Mf47DdTu6Mvm38pzPLbkiNJXgwH3mHQ+421vMXdOqPgvm75tn/pWCpq2a
GVdihnwcO243RO6I0weZPaWi/X0SqzFme+/+d8s8t8A/tNun2W0tfwr5lnl4
FgjjxGzjcP05jmhpdY5FJArQCCe1XpQiY953DUKY4bqNg1HGcn0ftjKToTI4
Yv57QE9aqQwVkzxjPDkVaiqJgMwsAjcFEDobPQp1yF/slT415aJ5L7rw6EqR
hATAAL21cG8ORmmXkgX8wyfHKNrjsbWDUAPKRo+qm9NwDy6xiZfIB6ujRtMH
q4g9d1loREZYn+ojjEzeErfMz7INEw74pDftG7cCaPCiaAtHupaSnVYmz/qL
0G93SL7leralqa68XHwz1Q2/5P9KpxzNgVDYcBd3YOu8dctJfYXhP8Bk/ABH
8T6yxQXsZJxh32lLusQgqjm05RUBQaA3we+beLwS20Ry3Pxjpy/QNCnXqcld
xjFsMe4xBBYt2Q9CiwU6oOrE9NtEexRRHmoe7Sl1aIwEBR1vpiRX/eG6KG/C
tL/wE3ro1GvjcBa+jc1qfW9agyBIwxYlGeZS+vB6VQqgJ+jqAief3+ZoutVE
s4/KQ0whaArcJdcvaIA4Q2QmQhY0ib3H8F/B5Rz8AncYHHpO/QpizYhXP51v
Ywav8pGJHOCveVORDvYtY+K1Omm/ivLWs7N7/uibojNuvHParQdT0eRsmmIi
WIWd/wyp1TMAiT4VebFqHkYSHmkcvvrxK7Q2I/CE9UDbCgrco7M+Rd2XhgCz
0cQqs/txGzCAQRDPgOOV6Duqx0dqXldMRFUuhMhX5imx9I/lH+pC/pSbfgEN
743MydREghf5s04cdlwF9zb4geh2iPMDaLmvMe7b81QYw4N+LR2hstm/FAKb
tyPPDeVdBdLr+R3ahufpC1qg2PdBhaswpFk+X8vT6ktSmk7qp4cMPaRpUBU/
vpuzUzX7vcUsUGeSBG3b8NQhtzF9jLS0B+M5fH8SocY0FhYsdXRH2iUTySN1
odg9iiVIyEYeE/V5ROKksu7troJ51D2vU3NS6yuzctQf3+DrMiMgRDwpZ2oi
QcpUF9uhduX8HLwpmxjzj2aVEJS2h6S5UI43MI9geg+w72L//3ArgOw7cAAi
XYzIffqxrEEOf5lgIUzKldUmjVRakYasuS94ecTiZV2hdPYblz06dnIDwXLY
yafy0wEBbpuAg0Dxwyp45Qi+tTXBIX3f0Ts0GdUuR1kdpUkumNDm+elfupML
cj9i30B4ITNTpb2vbAvoUSfGojD/sWdVQJEsuoZSyrma0bVO3B0VUD2WNIsX
L0WHgY/T3WyGAka5EwsWKnPKrKIyRfYoXZu4s0h4gfqJ+3lyZCKjb9JPH4Gw
YifyG/0G48FnFQdqKVlO5VEpGVMx1XuPyDW4Nb22TuUAoIcy5fI7EVDq3sMi
0cwbj9QYqilTZZQeW4uXeVoVl6dyxFqw365AWnePI1lqiSTCK/GWmp/PrcIM
YN5CgW5Ecvmx5bOcH3GQ+PGq6JtFjBVjVFw2SDMRxAXBGdlJ8Ns53XbSKLb1
uT7C7J6E3FAX810RcNo3YpKn4NwyaXObgNkrufZPxCWXL7H8IShlMIO+Fjon
8IQTgMtgqFWBw447Q6iaX/0UaDHfC0yRS3TmcqnvTM5Eo46RIIZubZJ3AuAH
oez7eL4gAIImH+GqPCgzdrDGuF35wOkXpFUxllmLHA8w5/f4TFys17D1AsD9
IG0eek5OG3xMWDvy4FVFSGnf6cInUD0OfMBIeqaztkfSaGIGQzYCwDqp35U+
pNc4R2nmEAgS7jgzOEN+fe6rtzphntPNFE07oUIOyERgCiiQaWKNCC96kVb6
1JuVmbxpkCCdRrs2zMVSNQzlWp3c7s345vb1niScDIqSm5CCTuVL4hi75ODd
nTO9Lhowehz0coWrLD+a+J0IoEPSgLB/CV+0akJ3rLjUQQW7AOXj0/jacPBe
W5umdMoRyLusruVoULj1NVWnsZ2K6B5vBUCzLPi76FpGMYwzH8txG3Lvu9MU
iZMFgin/cn/iybYlMeP96mQ21hGXyWVykf6Qj4KyBZEWrbRJlxxxknvrrktu
bWTFfv+YmlqqOSsgTOSYRn9/Ykfj4qBW4f2KvWbgwU1lIXLpsQGj+JMY+g4G
pVeRkdXU5YUQ74g+r/XmcgtevYqlXyRcEz7JzqVMAtlnmTdp03QcIaXNrmfH
xwOObbVOxELhhpPQmBcOBZPFkDs78Mk0oxIox8fVaS6BWBvXA4/c5a9meug7
vZbAUSVIVhvKrvjl7AiztiJTZuoWkJE7noEKu2UJrzh4PIlFjEIPSqidlCs2
tHenRAec8FQZehvWph/vx968RjhzcQ5GXBPIP9NzesnRFf7V8vMXgbtvxT1p
8n/6U9Met8Fzm6/zUAmCyu6jSMCJi4BJtLA/pXybINv8nXn2A6iCwvJph/yp
wvHNDfdrVrMd66Pt10OsaITFjnNZF22l2H4tnty1Tcd4Kz5QBRZ+1UNbqYeo
yA/qy+wZ0iYeQD53zokG0FATFabiYLyohuG7AGz/uVacDyIh28r0uOhWk3y5
qxNSat15R3UxEuDjsPpWjADdmtOULDVQU9dv89naCxq8myEZnV0g5j7Cy5Ah
26R+2l3tWQT/wXF6ownTa0ICLanRxIS5wTfepJ7sniH0xfAiB7qiiaS8ZtjD
wWolwxgouf26ssA3ovpyhRrKSEhWHV1xbmoNSeAh4Y9XTHP0vf4ropBIlAEW
fxAXWU7rldC/VZZfJe3eBBdFMpBDsRPuztdWSlGT+huHYRcnTRcOQFPDUs4m
ywJb33XlZNsr3GBeiHqTqHL3mX5QHiWBwS9F5Tf+KtmaF10R3vwyCjnkN9we
7OXfDHgwHu8I70vr7nyNsE+Gtd18tdwWLM2OlrgyCkI7iFf5FVLMLOZdQKn5
Cmtpwj34mNReCDDZEHnE4b69eWV8vsFSsWQItC4FVCJQ1sKn1QK2rYMNNUm8
WHIGdhqRn0FksXcqwxh13U6Kf4UUk4irgI0vrIqoJJD1clzKigtioRU54lBc
C6WbFmMYLf293qWY7VyLQk1hOytlFSFPlTuSqRe9BZIAN8+pwr8tf+xrCEh+
Mo7JhRiOz+axHjdbu/b1c8fQvwpTmFXkDxnNZ2dzFoML0zOFIeuE1HK1bKjn
cPLDbZNjlCYS9YQgOIZek9lvfVGKkqV3cUTW3TSq3KCZk03mDz79qA5qIHuG
H8FimHTILydHDHyRIkCetw6xB8lcL8qcbT0K2hnh+6DJo+PqFwiHioZG1s1C
NSavL3WvNDlynO71Fp6qHHaW9kk6G8HdEaOsSLQg02vtzuzVMKaFfmN8mvA3
g5/su0QvpS0D36VVLhU/da/lH4sng8gjCfSMhyh0lgy1dSvapNCHLbF+pkjc
SIn3aOEQpDY575YzoYdonq5ES6aBLGjVbKuAm0wM4kYFj2AFQNEbh+OUJI9T
TlgOMtc6713ps6ANHYIUrfTqzDNjcQk1rjYS81AXnj4qNH6Gub+nLt+jzinZ
my+Hicq/Zf2TybWAyiec7N+sUQ98cgGaW4p9LIMhXDbwmapdfbxV5J7ePR30
F73VXXt1rUlcXWd6oNIf4NIhDPecMKr1AIqYovLVGeJvHE3zc4M/D9nzCSlZ
Ppq80Yelkoeqtp01l++m6Q2DO/GvAHmApxXU2V0GVul31SPDGtrh2Waf/eCv
fPGtJ0sXshFrLujNQ0rI5Fx0t8uikm0Ox1hTV9+XnmyUcCgQbviiHJWp6ERH
zeQAwCWXH3U0L4OtYDJ3VMebCvuCiO5YylwQILMR4+RDDxWrF7Zou6IWi7D0
JRzPMmA0GtXAhATcuiwa7cozKq+wmAPico9832aZ/sv84AufR95c4rqt4osR
n4LSzOn6zcego2OPYh8EuyFo/XGamE3EbBHkcrvoNPktw28iHrAUS8CDihHk
Iybc2/srLthhKuoHlS/EjD2YB/zIYNmJoJlGiLNWT5reGZ/JhNTGBRZdCFQt
G/G/HWgUvLDil/rJ+4YICwBLvnMzqoUATwACjtAgP8t2LQb0lwA2Vkc6abEy
4BsPzk5tKNG6dSYCPnUoO+nBFULPRIZEu217VC2q3gL3KUEJ27phIqLhCxyo
v/ncXTzmBhv0a6eqr8yTim4SBwKwUouiqG1DKayp2T/Ky5qZaSHCqBixKsto
Zl0NSXhOItnAJSngT3TPOYohoBNORibYTvGOLIVtvzwpB3FaXn1j6XqChF1N
YZ9xczX5HunJNBnMP/QATbbCslYziZzX/qOBUe43gGcvrjKb4acaAMgzmz4p
sphI2EMqw4fn2/SKOnhcRzdIIQk/Tha0Ljycy/GzMAqy5JNfXPrixEvCq1ge
ltS/4rkJlEsUR0RlYkUpasaejTJKQOz5e2FNUGuIu/2myYZzWE96tygEZCRO
jVNxwGDsYBx4w1B3QgfDXvTf09eiK6XgUqzFgy2VGgLtUwGzg1DQA6uuPTTb
RVl9xEy4SlCqixWOZtdiDjq/mnVpWSTHlRGb9rKBXY73GlUk6nNdcDjRovg+
kCUN/pXhBI29hjPiaa7GL7KUPJ5NodNYc9HeIpH6WZV1D6v8K2WW3ysQJtPX
YpCRhNNCurElw39I4Z1giDGu3FIHnh2Ep7+GJ+Jr+NPvfSxId8sEHJbO4kcG
U5UDJEgy6GwZ6p65jbotUh6r8yxCXLPvez5dFKdx3DAQzKbxAXuUDOqpDrBm
FsEgRRzOM9+Pmcr0P40M7zU1RsCBSimwUMc4nuBKFCe/rPFWmxf3Fz1db9EA
G2c6EOI6mUTbfKgaZ3mw75gO/EYAuT3u/GhmVcXeUcjtJC9tuPKFZrmBQ052
/BW+X/uwBvuMwgRBkulMWp9ZATSYUEEiO5LyDYLZ/4UyE8iy7SZ+35H3ubxc
JuYJv7RKu3GMvAxXSB7Z4cBujEHQkCPSOE4UQkEYMms9g/xQp08jn3f1QvkU
X9TMz2NmbL0c+f0mmq59lQKHkwV3criifev9xUJStB29wVSTml5RW9I6kbFx
Gh+Tokmv7Cczo61PAaB6Ge09yJCLFHlI60Ahth60N3JoyrtzQW1u2uicxR8t
vnXk+L+OruxFlDf+h7Jn5f6LFqJgWz1XGpOeypjFQv9jvKo71w8/joORMLhG
c98JCzeWamPJXLr8bmF3NCZMBW0rax5Aot7++wAovG2AMqfC6lZhYtqwwloO
iG3T4WTgn9KrbS8NTuYuIcTqc/hIKQN+fgLYnfgg0k0EodVu9UVB6S8Eljo1
MnR1IeY6pWfntT6CLcK/KreI6TEg9AJVMm1s0GEpI9JG46Nd6DzvgDhJaKn/
Kf8sKZ/Ov+lD63biFOT1u9vWmFK6m5nYs3Vak3PNEJ9uyFA+WgxODqlBJry6
IK9w4BGcD8wy68Ai0Av593NcvpCS3u3qMWUQO5LJG2hcR8lksfOgZnlIWU3M
SdGf+uYcm8NRtrdy62+ox+HySmU6DcqW4J9X+xmKTbV50X+T93XBVaJ7z0hv
VF5nacIyk9QpC8vGOqrppeqILBpuOGYydc6CYGMjxTpxrxPGEz4x+z6+q1a7
r1QrNEP1dcnQnPdbD+WD3cuq5Z1xkrLriec3suCvVH+40q99b6lInODBDMtm
7fFnIHg2Vjjjszzd7YGfWvsZyo5rvHTy2yu0DLletjiKmI8ou9cDUmYZjUhy
o5hPKIm2C4f7arhnOwkyXBzolC/pGf3PCnmkYk4+eFD+IYb3PqVyXYqPaAkW
yYyjFxlgJCJPt6fRogI0+jgtY25IFT2ybY3OmY7Z/Fe4L9i2eODCm/SImCyB
gW/nwaIYsEnLBEFc0vemTVN6Qc4h5VeI9ZJNEa9Cqdwrllt1eUEywt7xsWgI
EMZm3v6p+pq/q4L3/2kFjN+krvhk75V2oSh4ufL+zhaESbx81s7QKgBDV109
4wBDEhBYINeNXBlbZ6yR3tZfNb1X1cGpFaTahIamOzwbLWiQNeJ5hvc3wc+/
sv5a3txNXwEOptRsx6Jh9s6j4zF5SWyfpkSIOazNjW3HJyWBUGb0JrNvM+id
k7sQ3hYwS7cf77gebz3wfGPKvOit/5KJ9DRJHloG/tHoQW5RILKoXy9LAn6A
jWa2DilhAFPYinxG3dufIdZg93CG1U/QY2OxVcckjxn/wH3+oSzIhBSZ9o9H
3FM6//KIzBJKqpFzHNAZLj1r2ZNOQeJj1wemOlD0NRupjUfyXJb7rildKh+0
JWUEhNgbesa2UDC/P9B9kiHvpYcV2vpEePHn4Whx8u1lp4awFpOm5hU5SNFD
IsKssqr2jJNnzJw7OABkfJCUPKJMBuMa/ORQGVLMaCbv99cKmbAD0t1YW3Gr
/nv1Mr3chJRc2n5/vwnAn9+d3EOVgIyWVX3BnexhTWkQmbCRRVsG6Cu76IP0
3Gr45SQCSQD44Lj2norvVidyc9DXJSpkBmMD0EhLEvTMHw70Dsit+WQjJO59
oBCvMQYubaOFj29ZdZGalGPZFgQvwU9cMEGEFUCIAhOiLkBSQWik3juF1x/l
Skj+xn/2UUEVr7Hyilk0BpmsVIpgHCWKZ2Fxhf50MOMfGz/w2Dr9m8Qqzwwd
gPzW1t/PKyPNicLcqeLf8QBItyWdO9DUMf6w2Tf5LQBB3z9Bkhu/5P1m+rxm
d5Z4iE5ZckzJvFXWnEQxlZj/5paJtSjjyW+A0197J8nD54huqpOoiDdjWuAV
RbZ6pWu5siMd4qIFs7/mri151B8v+5fB6xFCKJqGk5BkXO+cuFBdYJZNnd/F
f2pgpVN8rcze6zD/S7joa8+eAalCkVilr/rOe5V0Ib8/m30UHG/9OhpzPRkR
ko2lyPnAu3kyS3C5NVo53+hG7TN1yxkjrZQDWc2D0iXwSfaMFOjUvBb3itSG
qpkLINHJoBdlYZCNHq7pyWfFWB23VcPB24pauRbXWh3rsvFDWVUkePKLiRRu
Y6HY+iWONHlUGe0YITkfkYkzvnU3CsKgnBLcYIJi957rAV6nwedCcFmNrT5O
2MI3THpeOyBTP6Q79T1sIP8Kl9YldpEUCaN0yNou+U8BCeoQ86V2pXdE9wS4
qKr8WXRtCJZHGnUHSA4XkQ8MpQrLn1zZZjO/IANUk9uL2FqZNPubI8rbuBSI
KJuPI012s0AgdPKTYD96BFk2x0ocLG+bkh1VoYq5QmHWsFuyy+rtTFdbwvKP
gIbJ8c7Xm2JawUxjHa8oJnvSqVdAbijXWZLOqJTdCmOIXJPwb4z1OXkBanfg
5IoZFdKJcl2eY8GZjc7BgBWxf1J8xdvRqRjuBa8ufAkUbkTPoYmmLrOt0JnA
bGkYktnmbDCVlCb2VjRqA5kTtTm0CkC8Q1LMwBRhp1wYcVsqVzQg0cm/dJ5/
rFZDAs9jKhVICc3ASPkMJC7XumKoP368zA2pdBgobhDbKgIYHfcUQcU9XaM4
+j4G88CqjT3uu2MRIhcA13x+lk10mE9fhrYfmee9Nfaa5XEvAwl3DF/z85d1
l0HuKs25q4dD3WjSay0O9N1t8qDLDrbS05wPXA34x6mOQZSP+LrjwZw9563O
uqdlVaYEonjncbKoBqPGgmmR1B7yalDfr3kjuYVgtDBz5nJFdji3cYu+kPvj
wkBbdSDxNbBPEhdmRziVrN1NJtf8hegTRRgpMPJnW82K3F1tLEX7SH43H966
onEhavAPFhAtDiaV8qHkGzUXVU/JVfRsxyDN8zJk+luXjSmud0nMQmB7EXwD
iiGWIaIy6KspH0Hr5mjWvvj4mGrw/yyviI/sGFpxBSoG2juBW3hr63wpCeuq
fWyU33fbGoLHQ/7NzDuyjpHQdpw5JfMsmGmRsPTviF6/AJehyqe+l0TAmkjZ
I4hMreLFMM6ro/bCqWfdSLdVgrfC+WcJh5LCwttZv6wTTMpup8k3aW/Wt82L
JQ35LC5R5l6EbQI5wHXGwwZ1c4QmrAP6oMB8OgdKLzin2BVIUOrdRX9SpPJa
YOyMUbG5wNn9iS3INP3owyIcm7+UXbDpmRKrFAp0hN3CsK6tAHxhQohQBAse
RzHyQg6lxznWrs50yJn+mVs0orjd8j63LBrQmMrfn+q2mxqjdbRJ4ZuM2EwS
sb3B8zh3huKYR9CCD6c50UTeRdwhM00y2nUJ4IQqS5Vci2VQn3lipfPL9Ig1
2S9UNTeZiVKAB56aOgEdfNFYSl2P9DTGJ92F1XikIfoAdWmZ0X3K3DBt+kub
tr1R2xGeLulmOCVb7WWNo+DLf2SDgAwG/M24OF4svGxwOhHqeq3N/4spws/+
BTq64yDipOPemhfUTuQUyiMoLWVSKJ2kejKA8A7GadIMeNMaC+HoRPCu/62a
8URmHh0k/NBnq/21c9vrqtTxWWF8foaY7InbhnUElJ0f+/KG1kr2SjhAaQXM
6sMRf5glsdoDAVXpz8wrJVi+d61FkDA+aMEjtW5PGBJFEELg5vN837cNODuC
c8kJzHJWcfOQp9mmy9YF8lnquJtAN7y27TevMZnFr+UFnUUHBLLWj4s+ckTG
WdHFyzFTZADmdiQk6qXrlMJgHf41SpalKaJ5iVxOUYZtozTpxA003tfEOpjn
z6RpzRfuTzY4WWZl6+kDzsf06gWUKE6xNkUitNF2UXS166Mx7WVKugLSvWhM
yFdeifx/1KirfSVN1/nfosWeXQed1Iauw4TSBz1e6H4taPtdjJq93qsTYA+4
P+jl4HxDbtTrTldknc4y0mEfBDLEPthKKZs1LhkB/fBXYDZ03acfr3lCYfBI
ILkZng4NVb5sb/RjXjRW5rslX/1Wdc+xkMgLFhPvZ+zVc3RbfbpyZsPeiHAA
58/7fq75DE/n5PFbGlF8xin9wbkxQuENVC7R+m75iUjz/zFk/MVW/fOC6hUZ
DD+E6d+aT1qzi3dM3m8MqmtNpn5f6w1ueqqw3ekJFmxYdbhX03PNYVeVqCI+
FnsGso6vunrcVMBL7forEA3hSbf0SMpEGJ85JvPGBgXxpPXOtB9/927mt1bz
gwKirT8vOwlKoTVNM/2lbRfqGF7Krp/UAI4cfYpLyx03pXnh4VKyuAJSydMc
kKX2sew6uHZtDeCvPtOll6amuxIAwGQ1vXg4T40itrCwvxGz5ZaCawYid6wZ
s8JHCTsZ4VgN1yaMe60Fm7vY5w9WkxDIgnskw0enCL10hNMPosDMAKIs+/eU
8H8IqTpEQMTR69VMARzfm/w3LYVsD/ZknM2rmHDQ1HM/D+zNa9llokq7ted+
BobQSWyVQ1kO21FfKouHWVslkOpbTN0xGp0zAR4TbVz/JXaNtZzIdlNI47sf
rwyZjwOtrkC42s/iafOXGVl4+b3JtzLbsJCElhG8iY9iRbFCLbc5coo+YlVv
gEEi8qPw0I38GF2Kwu/KWfx0VxTG5WYLD+/6R9aZC/bt40HahEw5vJcSKC5o
APSaUX4iRyuBsQRgXS5ly++aJtqdyhXLtMV/t24T4Eelp9yuHCS5S/s3Od25
pvT5yihcaeq9/9sIwckZruMYxGZQ/nsEzU+2NcyrA49mfqfxwmU+R8nau/Py
n0lC15kB2v/3ED0Re8Hb6ASD1qbXRgzdGpFZadi/IloAF2m6VDL6wDQSxtpC
mQudODpH22ruVsWajDGL/Z+yZ78nel4tKIvVKGXlQ2SYleblAHS1uT5hyGDK
vsVYNNmEa5UQocTxmipuwJWyois3UlNjdOuUW5HmiwM9OJk6TaomBwV81z4V
KQbMjhz2lTdUfl7Kgort0qFx9vhWJm7ZS5IWSMLtFEz4zzQKA4Eqx0XKeH+k
ERAO7cCCCRHoA1akTPBckyfjc5/j7AaJHcXTIff99J+Ru0dMncHJ0xn9qWN/
Qf065SBCuah5/PpLar7jQavX7GprKywrW1i2REutL14wlo9OUI0W//LvSQXJ
c466WF5ebGrFYy0eHTsULJUfP1xUMLundBVeL2UXW1Svh6p+aw/Uy9+mctLc
O/+1q5EkuE6XRT3CG00bYXuqG0WJ8ZkoRFpXTKXNfxcWhPEZ0ecLfMaQJwug
PDU+9u+/g30FxuJd2Er3zfvlXdIGDodyBoeSikfQOZXngdRA1715LwOqPvB9
7xuA2ixbClQemt8NVMZqdP4QsLeuypVQ17OwanGy9UDSOGw0yBHIsBPqeuKs
z0yzTcm2z14LVEHbGzn14R6bQX/MMqYx/fxjU3UmSrPz/Xw6SrldeZkbUBWG
oFtky7mzl90rJgXnsBvDL+MB+CD+IdcXlOYPBxwLTE8J0q1S2koMKDlUfk4q
v2rN9zYWgNCm4W2DbqeGk4+eIamj6eMspX/OLyvlBxvUFncts7THWdACjVHk
asJlosh7t24Z4/ARVvrW6v1EVP/9DRkyektXS2Z40jiK5NvCxEOXcRJeJtT7
HWqmL8LE3Bxlx1z0CgRUgMW4kcd9ZJa2n2yFvigOKCRClF+uqmxwqnundvQT
G2O++8/bQvL22O6wI10WaQAS13pY9zWHK1yQ455vIw3+Dgx7WbZDsEwOer0N
a5Z5MR2uPcxqNiLFzbryCjb9jDrBuBy7ZJezjCxUW+40h6NjnEY9YIyJZzVb
abx5aChRbImz58a3Ul+ipf6sEVp3QcRXZqfO4U3H+xp68eSTBN1KGcHrEqv3
VVbXVEKsRVA0GsG1BX7SKpBfUUiSEmAEiX2kJjs06BkHgRm7cobG/dEJxLCw
4QhRtOO9RtmolVZVaDItpw+te6mDLWjp6p1qRESlUlhdaVtZc1dR1G8rXPtd
MSZTbT+CdAxmCpEv2eU8jp2PilKk3mHmfHn0/KqZaTDKYzXwxLZS/LE9ooUT
ve01rxkEtC/4hVKPBa/rCSo19XSlqit5C5hFGucjxyV/dgj8OM0xJWq1wV4J
ug7qClwVu/XYGs6B5UQ2UobkIo4ClN1p6h5WkA10ZefE6mnlFwoskT103XGS
CF3VYWcRZ0AnKgaS5Ihg16SQqGfOhGmREDQGeDJRhbckp0YPTBvI08fUiAx0
96xsjHuh1iDzvwRlvghtEd/ITMJ5tkpDytJTzLBDzGGFfP8NMrVpWAsdjFf4
bDVRzigwzivRBJHNvpNgKIMQb1w9qc2ERg3k9vWzBt/fC9sYceZ9pjFtpxVt
MdaEgLUTr0qZcaOSWgm/2YTLKVoGkWIaOd4fT/fNAQn4QJUqF2a9+7cBI76U
zMvecFvool5rsf0aVBJFBwdnRh1LFwvDd0Ru2mOymSA6dBhRCPKPwT0SiYis
uhBelvWu6pbrjCb3ZGdFtTMqMFxBOaVy9dGV4kWxNrtMybE2SqVbEYBCmcJw
tKuNZakqy0voQs5ymQYLx9aJINxhCCtgBzZ4Qmvoiq/84ELh/w/7XOl+I2hE
fb8nhx0XKp+FF1+f3pkcC8XkAA1uBRQqRqL8sY56u/jQ5+yBXDk+AdURrNaZ
P2SJ9YEaPy01msK/HVP4hS3BWwgNb3q9eKaHl//Hxn0N8rP7HGRxTgHMJ37U
zOhV+4uNRPFz8GcrIZLlQZHZu21wJBP8vw4hERiGWailluVNS9iIMXak4cBM
4QVFKmThELa94+TjtNh1Jmndf7XxI39NDA1pbqsMN84LLBezRS7Y+Thkt55I
A7cl8I1XbYrITJ42DtDVpfbwrRzgRxPm3xvWPPZHlDjE46CoxLAGLW42EG3i
YocFO3CkGptliTeqQS6f1wkuLTyH5HjipI4cTLQ3QOy+/9hgtQeIV5SBULPr
h47iOAMlqoLGvH3YrTeNnXZxk3imcAhRE63MxSG4mHB+yhCOchMwAK5Oies/
xaDXWCA4kBH7JPQVokt87/Y9pkkvJuO/G3WFYFPpn2h6pf8fUiCV/qEOJ+ZB
uVRE/OHB0CFpUpheRD2CJEVYF7/fxmeaRVfkzlXOduJ4tnvOUcuekSpyD7ro
ujkhcgim66mx0+X18zOSO1ToZiV1kEceZrhxCDUe6fs8xoLpzuKOoAWWJq39
sv1rzndvM3HJm2qZ8sTjvbxspVJbiFV0GlqYN/DHxQW4qrM0OQW3aofOwjK5
rHy7XU9FArJpw6qFviMQAroNZuvrKHrDjPLQtyFk9zDmWH99B0/K4Vcqp6rf
BgOWOCzG5Xjo6pCIMfKik+cSpQhy8hRClV0+eqxTBazu1RkQsQ0jEG9R4G+4
36Nq0iGjuIgmO6rcClLqkcmUjApGv5q7/ouRzEKBSiisH95L82hhDMIElIPJ
IKbNHJmtUgwfaNligYsfW3udXKU+81h/j5LNsbbzC6wYlYuZMIs8jgr1n73T
RPAC3oPqLcXjDq5W9WBlGLQDJZAahEsXqm7leqP3wpBsAL4/4D0DpkBHdsj4
+UwDpvn0cWwrSWRL6Be7a4LnhZQi7JNbFib/M/6aPaXASTd5EHinacMBMI68
Zby31Fea9hBLmloiZTxr/9Fb7rI/Ov5VECCRJmbXXWZk+C23m/5aFsBAQVhL
RnohEEyiT7ytbDWorjeKFlTG6YtxOmia+jDmYs9wTXYIvLIv4bRmdSqJWbYj
yDtgRKBdvSlgl4BmrHVe3tdvZrDkU1tZ0EjX8ohZhXJI6MI4MWi0RMm8GkE0
nNnuiX1Y2YiNw/AkxOe3PbhScyUMv3+1F6IY4/pGLfHY+qopy4vvMDPAZ57v
+5pv1KYiv/m6gstxmpx1oiHFcIaJp87VMnuzcHLFKfiMxyPnirYSDONqYNGJ
gaPWqIdds9JXY6tgNFfdwqO8WXJp1mK4AhKE5RveouxYl5uh0yZFjrE2iTuz
6GUpGUr+krYexpkehtKdDZZaC2P1bXTJ0LgNpsXwi6ExN1fkSzAM4n6Amx1e
6eAT8+PesTlmVE3YejsJwGJTkulztM0qGmwlAxmCIW0KdoEOgEH+k6ccgwn5
qhGxnT4zy+aBrK1d8QsAkdV7PuS9NxDpu7uoNzXRviOLsB23GuU1HZU1Q2g/
pBcpYy26j7oIIhhK+sLV/pvEes3UuotcEHNMDZljRzsHzvrsK8e0Wya0WXyG
D14yKhjLkg6Hu2rwhYiPG9PkIa5tuKAhZTEGmWXvzAhmyamfWzpdbLO3VDUn
ycMtddsfl8vqbBfNPvkyKxBAUBMZDJrfzTXXsk1acnByFKp+gyzxtF0jWwPv
ae7xNMcQ8ZeZ5TFjwMDCND5d879y/5uufb2mhqXagTHtBnPS7CqYpJv2hnnV
wcf5JJUACXPdwoDArU/BjWshuNjMPihexYzQEY6ub4+lH0gsldH9LZxGfYm+
hgntsQzBWr5w3pY7ckwBwnFs7zC/YxT8MKuL9hHTccHD/wgi+Fk7GcICzSWc
0aPq8jIYBxe3IIRwlWOr18tSxvCoZ1qfRBZ3+2UnojblJeWyqf0JfYjZH/mS
QaeVxE4GekUvRZ0U85J8xGfpJusESRTfQujfjrer3Tey0EZHzxE3ukTdUv7G
LB5s+GYBxdUHhWyx4Qdhj/cwjqrX5b6hIYzDAYCDsJmNJPKgwohSVzy0Tk1o
KrIENQuLnf7BNKl2aGF6Uc/xFuFZ+X0goKoQN8C6coOGGV7B8sOqL/G7lL+C
4RD3Gy2VCta2+/VI4nVmFJv4knA2envqDOtxrBfpVMxRC+nNat1EABMkwVpn
jjtiPLJKrVN2xn9MZJOi9a3n8cF9EoWt3do5vHllHciABvArYe/AV6RM7e0M
JWYFc5nGu9exDdPfhkq4rOUSEUgpB9NkDCb/nCLAeUdBj3tX/SzlWsNsx/Aq
f1JoYvz+SQjtZa2ln7K7xs2Dgy3jFXlpEBJqhzfihSnx+37pPRWha+48OfTH
36P4XHbQogKbVsnUWG68mpAJNagTse7T9orDCk17M8GceaTTCnKJUbMfatUB
A6WKnVaQ7g9b7qQmQr5bqeZiCsUX7L22bFCV7OnUww7/CdvQUDGrbayU0zDf
BkDZPWcf7tC9/ARvmT7TUwurXWIrWtWA3/Buf+PWfmkHRsACTOCDLtqghgkN
mjj1ggoklVZ2M75qxUdunZK6YjwWC5fW4sf3+vvygC7C9m0dLU1LRant4kMY
orkP9BGSpRXqQOQ0zqfWn67PVFUXx+X36wWKyRptDbjMQQyl7ijFxXB48cnd
sisZhOQtvgLck46CgQwDTiMp7V5jWD/VIGNSw2H5DEJNQUeW2I5cK1WayP18
jYF0+LAHddZtQ4fPXMIauxgplwhejBztBuMdhQw2vKqgfX0Ma366CkJ+3eVR
6LuxA59IbDLI9EBfZewvW/58KuscbdzYu91BYTaGUIr5kHlgXIDKKz6vSoVD
edMp7mmmw91+tg+0cv56uNXui9CGJHKwbokbIOHo13kpqDRx26bblWo4ynJi
ZWzPgd2BQR6IMPBWrwab7l2LBNJJSkaHcLOXAsOwRmtws+dtO6AZgPVmt4Rj
/Aojs/kOThwuskF8spJNI1xCRM4M368EM8vFOwZkpo2xKJPjxSHW4fcH3bih
XZ1ZsA6fMwK3ZmBtP234oOpi0JKRAS63ivsUWErJyR5692s25h0HBUeC87Qr
XZASD0gbgv3fn0Xoe25pPpldPFrKk3d1dHVLKo/hX2yJY1/wEar+R8jUwz64
YRAWWNkZ1jNVJ46/t6yNviHIGVOJk3AdPBswzqTWDXoLynMygqXP1KNvHnFK
XlsGF26lD6MhhQMrRHWIj8qM57zMKdoTih54XCj3WOQyh/Uw7VWEomI/i2ZC
rRZ9MyhsNKfRHKrQTXt1UILqnezvGr1b2J28gj1EG+i7ld54UJaQDTotZEMn
9YQGkpDTGoc9OtaqET7SnWr22NwbTg/vMthGcM/L4yzku4af/QwLdu1kNheK
dEr0x9tA4v53kJISejDtqiSuP0NQl2U+mBSJK8KvYFEe0pd1iPeup6+7xeDN
0TG/L7uPqR2FHHv7DbCmJZogn/q++QH8Dm4XpeO+u7fFUGxxDvy610J3EIVP
xUUgv5oECrXS3rKnr1oTgj0ZXbmYbYIjlbFpixuucovULvRfnwxNjzsQIDxH
aK6V3Lx0e4JM26a72q+IXQbwNPhfX/5uE1bNfBle5P7xK93+sA9QtP3bNgyd
VbzYQTon0KU/KXxVTLTFSK+t2CDildKENxdRxZ0kPvF2TDuOw1JpOVgUJjf+
BkwIC9wcGRfk2cfHLIs1kT1RVZudpP+SHQroB8kPzpmJml0Z7WgoOq9bRrOE
yNNCg1qzOCY+sdcvG+KUD0MkO32kTpHQ0C9W3Y1jkUp3KzQRbA38y9UeSK5U
hT1aqsyvEm4psbm56+GZrZPTkgLNoD8dPdlVDdiHQbSBFmAFZ+kq1P+odHEm
5QnjA4dUWTeHKNju9WMaZW5qyNoJZQQctBgxzpkWbKm1b9m7jMgt+g63VR8m
VNujA9HnxNxRBdhG628g5YTDrq0ArONkcb7MzuxuUvy0BHSJPFiduGkWixua
EVlY9uhxCK1AK/Eg3n9HC7pgE6wuMrX2U8f8MLhoeyWyaQrWaTIrJVWjDbvf
7moMbYw0hBW2iEek31w+B3N9XX/mlVkJISGl9MPfxPOZPUVXjLeY7srRlb6j
idvBcCcjU1mkyBY9ibOqgpTPW/oHtI9TtSgF0lYD7jzDgLwrVa4E8vIILOwF
TmJrUdZVbwYvpGls/+Ws50wZWOuZkkLDsPHgEUPek3r+d5kdWDv5UXVxkLS4
dPGM7GyJgE8fYWWboCP3nfzWnz2IWtsoGxrI9fzkPqekiWMNPE+pHaUkCTMo
3Sqwg9t0WzwXBeC8Mj5Px8ToWBIi62w4pixtZV68Gc/GWd11t53YGlbpcTo/
hk5R9YAVn7m6jkDmo8h4tEHhZkbPYyejuD1pB8HLYKBX5t2PwGAkkY9AAg6p
STfz28oW4ul/m+jFK7zWnXFy1AaLcibcqoBtTFaaq6GvVYorfVkPcsb/qGI1
IVr6Cl/FwFzZvxmgR0yQQ4PQSmUTtRawZZSd7CNxKqXJBeqLRsL+ZpiNia5U
QewFQdzNrR5gNvX/NPwpKNkbLcc33iv16YgIgugsqmswbIycUifsSZa0RhtE
aj56wzayJJmn3KG7fPbB/Z9nQUCEPX6C0fb/UhDnhRq76sc7+9w3jrp9f8HI
tpITa3kBmHiOSgbrG5wWlmd2M7KFmjp/Xx/GTL4hrWwJjiElQcgxx1uFv6NI
lpzRgH7Nqzj9UKyMIefLH+lXcGn93I8WPAxdsPkm2nWgjWNIAYi6u5bAN0Jv
SP1WKcLX+wtia3fTJZa+em+vW9/IaPMF8Q2mP+IxTRkACLRK2dNUBv67VWye
gg4IWW8GtNwI+3ww/P7Pdi0P7z5waVSpxE0vEWAMNRADxJPV2v5m6h7JCgIi
BaI582UgYTorrxDWQ46iEgA2GylFQ881lIPKnCPeXnls0toyxP4EbqXJ7umM
nRFgazylzCfUROKADZCiyW4pb2Giqs/l8Hed5anKQdPHOrZxYS8WDrXj+dqa
nDJrPbTOOWOukMSYEXcUvxaKUiWXZ63mS1m7EVTsaRe76zcwpEwvTk3XijU4
IlnSsUXRHUompZwwOzUZ/KVLi/MRlKYBXE2weFSyDbG1VlgeiFSHpyjB1FMo
Hhj2LYU1rPJBvWi0WDvTexzYj80KPBhxUor4QgcNcK95BJVOD4xrNuf2x9Xw
h0tfFXzdUIavc5j4TjyN67x/A36AnJGUbdMFBR2KiJQFjOC3xId6R2bPRtpu
jO0tIemR0SsVda8if5xHGhplPAqx85Vp08xChH/s136ivRyGyoL3ds63AS8e
3TlIWs6HUEDJgaytlPQ6uVnzMl9Brfndn3muopXVTaH61Dh7gpOtezDdQPat
VQvPKZ+C0FTQVa3oP6jy+WspnZFGLTgTvmN0jZwA7tmc/OTpTYsrkj9XCKRN
yqmU17ukbAjlEmzFH0nxuyskglhM9VNVRrr7oaWMEXEN4MFc7Ipmxy0Vupp2
FCqcq3sHGTNTD8N8igrMrne8WwHWu1Uhcg162MtVcSHyiFWTB/zW/ZiCPniR
RWLFxivmk1BlrbE0lGR5Ns4ZCSgjknEw1Gkk4Ls87gsc0TzQduFZMOzcQvWP
WfOmMhTAe+8ajUcnCVRgNcnAiTXIMmeKv3dcsUStzHcaRcKvsTX3HA1g13yi
NaxxRHuiYJSRuLr30ORx6BBG5ZoLCweFVjb/534gi2RmoefZKJAcr3da6SBG
HcGdZG0a1Po7EmA1pKIFYOqJYo1TyQ/JhA9/Qf+WTBpfhhhK36Fb8OlTy7Qd
jToBdUKMtUEQfXu7WxT8Zh3hsQ/eyeSGYr10E8dAcQPq23Xk+yn1zswSoqmb
QLqeGy0Nz9DsbWtanZSfqQods4Hb8odOK6WWJfryS8fFEvfvfIlDn57BmcHS
sQ0TryKB5lqUpwoXgDvwgjOGJE3zqSbSI6Y7sUIuxn7jCWoCuz8GeRO2SNFx
Xm6GH6DhuWQT8I5lnnO3KRirgAGGKF+iykjiX9X+xsICZVVOIM2tPstAHjUj
W0nIPwCYy7Xqk/vrDi44+CbbZfe/9qtOChONjYy019agPErHGCQGwqjiGjwR
jbe/5mY2jVIwpsf/Kj6wHrvdMo5YkZRUjpsnFruwUsQDC693gEhP5uhuM3ey
a4Sch0gMNPZubD6j7ypEW9ZKzpNkFZg+3p6U3iRJaev3J/HZSW9D7/9HL6sp
EoIALymZSYGpjbOsul6zZ8Ntwjj9/tfXTDgXcVRYsOA41pj3jrorxcWXry6X
8BtgdjR7DwiMna8TD02Yh9xgsQtjaiQ9fxlqbMv0osDsCBL+D1vve5cchRKd
X2pyy8e+R2bmQA+zvsVOaM/h0q4XMoHFJqFZ1/UMOclbCCRe8M/TO2/S/bZ2
hNxTVdGuJYtczigFZ8P8/USDiyipqUtA81AagrQYK1pn4UYJwFa324QzESfR
Pj1Aj3cas5WwO5TPjBxH5/nyhqnxiyNmKQN0bJw5hX09zvrCtF6DoAOgx0eN
O9lIXmlqf4L3UgfmYO40zbuWbswxynHDxqt4YYi6TfkhCY2KLVhibGy5aGFP
9hFd+kYffa1qEIpGAWe+mi24tiky8P4fZzOAr8TCTFp4yu066YD5uWuoqdBa
O+y9cYItssUoosiamAZ4npC/E+iUq9Z8HTr5aTgLRFuZMGcbU96KZewnVDRD
uCEqRrtkCZlGVh0aKzmZF06mBbq0rACO0G2ZGwPrNhQVMIWsUG3jcCRKMeUC
Ra9DCsw1UPZ+Zcze3uelFdWARTxlCgPsVWr8bxIwc2CkXgsmInrRsz9+1L5I
/XE00c0GLOcnftj3/FGcuEe+3at8BmfwTaNV8sEtnX+x2LEzZ45R60vZqAma
pCEO1TOZOMFRRGISPz4O1ags8k+LWaWgFP4oypjOIAducTg2h+3+65JTwKb9
6+Nn+qiCzZrq+BKJdqsLg59V0LEDqIy4QxpxsiyG+DcAo5BpM3r3prEKHFNz
C++vLZX7XVztkOEYou3i3xUrK1uLf+JQFFiaKbQ25EDuOI3mqFGWoxXZqSYI
bO0W1Lzru5f6X5rT5PsajJ884a1OL2J3YKEeemKqGHA5b4F2csYV1boQme0a
dTsV/3bP3LGX1QAWgz9+e5yxLNncbUu4BngBy/Rkgb6neMr6nUbFfFuvTsa4
nkyGWDCriRZNRFDfgn0jD69i8v/Z4PIKcSaYsSa/iYjm1WxG/YU2Ai5t8kCj
1gy8FaL0ytqYFhjL5P4OnktO4YgtszozumLuU89RTt8CXnjL2XnMcFJxM/eo
gosjVqDSWZwx/pPcLSTDyyZIVEWcV3LmhwMJwrpr0K+Fv9NgAZQGWfeRjI1d
B6fb9pTiwaYKp5aDbblmdKuuPs3HzjWmLcxqPz7l9UQ3x4Ps2TYzd4yp3aBh
pFkEACUdt6r26VWklWKBy7bmLkafbFpc3RyLf8wSt6q4BeAefgjSU3XGQGm5
zZhuBQPS1zV4NwdbrW8bIfNL+KSaLS6NEu/RJ90TunLgG40Ue5Btcdsn264O
NRQFUd0EBdgN0la4/mHhCsAxbNv0D98qNEF+qhcyIwWbaaEc8nDIcJ4cfmun
0UujgfvzuhuXc7zOrpj+uS2L6p9R/PPmfTxggf5BPGo6Paz6O0HNPh6qdbHt
bUQqfykT6ekxpNGtZKzbSOee+3lcQdgpWzcTFwxJRV+ntifXoIzrE+DxWBUu
q/ja1Rtg/ChkEbRPFDkSAS265DTA1+tomwU17jMYV1L7LGPlPdl+WMpjfFHe
sUDgIK+VP6nqrXU5uptS+cET41cq7M/lAM4HtpZWDqS0g2TuKgvgV9aKZ74t
TzLwLppZJfhWqw1InSYMlTxCxTDF1yHHEJchF78uP0SILIYWFsOfkPQlUGOo
PNlKY1qdb/Sqekcis43CpB3Hg8NBYBBd6p4heCnB4dYK57Vj8RkRSZ9qxJk1
EgOe81XTpiSfeucCL+Q6T1HdglBV4OlFt486TQc+6XxzHSld6Ga4oXsE4tpO
nq3StJUfnJ7Tj8OyILj9U0x2uT+sCsYca6JMht2h0dXruZxJvH1GKcn9Ftz+
Tpvjp9dPnYGfzEYPJcIL/XmUa1/kj2+nkYhp0Qd1G0Vzw5Ttu/3OFxPBhC86
6YDtAlADk8Qq4lxM2UCldsSt7hZTF1J4+mgenmKuOp7huEXF+DnQkUCEE/EK
u1gcMrmTqFD3XQ7zggMV4LNZDbn7RWq61jYEdsLbPTM8vXGNQgyin0skMcrm
SjthMu3xa7IJYmbUcObh9QZYShYcdxomIZ2K+ENswvGpdPxKlDxmTpue1NG9
qC76Yl6p3dS0w3+1OlnrlMhpkBK4newAraxHsGZydAMAEhHzJuZzDIGrJpxQ
JZsoVnMUKMXfXcc4DAvOfNkKRaaCknicNbPf4OaAdlwP2b0WhQZAnR1NGQxu
fLIk1UdY5wAXYvnRpaFs4XQfQTTiVzpHpxOOKdIcsNQQkAtm84SgA1SGkNKc
sQbOMfKfDy1AZLf/Ik1uREMep0f/M+pIPYWDYswPeKIvCH+k3vrgITm3Zv6b
qY9w/uUkluDf/F7nuesGpFUAB52hdtnWXhezKoYDZrau2KgZktQQif7ZOQOi
qeJHtTSUopn6JVg8cW6QRK+lUdudhSRstO6S8VwCHGSaUfeB1oJ5r4e5Lh+y
6Xu7d9hmmc+96+YhUZQPGKIMN0hKrYALsV2xqIqZ/O9kMaOFkUIvTR/IrVOm
bcXwYfCTHdG0btqBq1EpxgGeDHA8dFJQW2V2XWZOGhqzIjxY99t4uWmWwMdW
TYKYYHZjJevoP5J6BOUogDdfsbYF9UMS5cSanw9dl9/CazlDBKQE8oia7vMi
/gq1GVh2AwxM9nKafAozJkDagmt0N6ovfUuhWlCJ3W9uQSN3SP+GIMOlrvOA
wSoLCaZMf+UQz8LfUjOzdPu4QDq4qHcbaqgCVCWjzjD/fHQkUNlngmQ0H4JF
ntjtvT+HI/szsiSncPKFFdOY57I0+gG7qV4L86+m0oGwzN4cEZRw3E+TVaZ6
uhexHOx6iNb9S9j9E4YChQcBesJfZehEC1HKTwfLvkryg3Vl/EUJNmz0fxqF
iOqnmBxQdqkVc5XGtQKpMQyzoGiQwkHtRO/y0v0oiTrOcxZDG5LEZKl/32RW
pS8LGZNMe2sCKP34iylAeVOUWdJH1kg5RTY8Ojyyy64FS+p/OkTXjaEU0kgV
yVbjOO64TFAdErhfD8Xl1cQDR+Pkn7xl1oghW0wGG363eYl1viUAJkJWnPNY
XVB2pZzWehWcePD4ecEnfORTBimB7Z66+wf0/QMrrZxpv87hLus9L+mB/t2r
8A7uCkBmtnII6xw9uRKMQ4s9kk2sqKQu9N1R5YE8B+cNonXZAA3HQBpb8Km5
aZYOUpuWoNoisrRt4H50HrCvI/cmH50pROwwlIsmPRxylEOp+uHVI268tZ46
Ts94BtZhMAqgZFhoNF6JZYKpWrPtFDltvwxcgQcASpKo6Wf9RasM0AR5K9qv
Z89MDOShka2xoywlu3IPs7xBbQiU1qJ9KH2Nf0RWPnmlDcMDlRXKzCpd+AOd
m87camsdejGKpWAtR3STV2ESWUW2WOYLqTMu7Seoim8koHCG/BT1spTzuLzx
euCmxNUnO1eYKzV5Yy+RHxJNpxFn0uCfTxLpMJSGKo0dZOmrqUrildum+/1L
CViN8cm1kw6TjPmL+t9j8JGyBGiuD9Q2FDAlMUWnbineErWHV1vk/+5Tq+RF
73BvB6Ym3PyTgC5KBl6IoSt90bne8TWwXbi1V5CP2Qzedhn9CkCzpVwegWKf
YamMaJhumn9iGIEtc7OwPymz1m7Qm8ZOgCKXn8K3p2KpK3pH6AEkRlSblsTO
zvxcxwqRiU92boUEBkQHsJMVuz3nYaJgQgbnkQ7xcw5RLDiAaHU60R+ZY3ZX
u4dHjkLRr7KRn1/vwhtSgtHbuW7KkEriNn1wAU+DIHac8fLH7h4+4BAMqDQa
/s4CqocCcxGwOvOKbVXZxGCl2Q3fXpwDdRVo0SkkAJ5mn6ETbS/AbQG6Y+J8
Pn5Agdv2VGQqkRtJltzBUaM/pWy6aKmsZ+Uayy/xm5gPbkk86Xp89PZFIL0R
7yaQs7rEZYkebIhHbzATYsSXktUxUa5cIyI5krNAE5dftmgIZkW3d6kthxFp
l8zY/zAoC6t/W/1cwJtKGBQIdfn16AEl0Dx8iE7+mdb24cwj32qToQkxbVaN
3yrvl3ZFwRZDaBeTH42shLHuOHHUpq5/lqivJwyo027+gMaK9MNvKtKxVbE5
eMxCFp9sQPirGdYI37D4j4AXvFZ56dmE0CPdeRq1KQHWxEX4CXPZlHdB81uB
4QfB69aYx33A4r2Vt9VMYJ05c3PLMU964cZ+oNBcfpY/WefhkC+6u2V6R7H7
rnp734H3PJaQYEZnjKFkuYaYKqlBqMurQ4e/dCAKNNg0KG1JHK6am32YJt2S
x9BfV9KoE3wnlszRvPbeHdVM+DHHMaHuiGPv9bGswH4m3VIvReq0A8IiQwbw
Ncy4a9BWVm0WKE3fKXKnvEBvu0Ued1ZwdC2XHk7xk9s6qyXiWodleqIyzcTR
+CSq81eqWIccVBpsXYluFNIJKhQsjEWfk+6rfVC5EM1C5cNogOWsg0EhE6Jr
TbxCU6e9JxDA3pApEhqmWAzO9AvTPHqz9msyOAemd+hyJyFtWymdnXePbxd2
/6EreFXUrS1zk7fx5NY+CIahDeBT6QAjbBG6kg+c2BTGAmPSeoCLjncC58Mg
VQDFb6aloqHBsSYc1NgnZwBYtNdGkwJrINpP/T1uCfkrer3p7TmO3WhERV2Y
E1Qpvtwk7Oy2L6slziqeKJZKW5sAErYldNHGmJ0Q0EbTIEIbkW0LWcXgqOhP
xzsBa7oT7sYW7zbff+hwMk23tGCjgRtb/SyddKq/UsluxzZIY7eoQgOWMyCY
mogB4qihUN0AjlfrB3zAoCmF2jmuWvhYMeCGT4L1PSpnfT8wxJa5N1ztzqGf
wSb2Zwe204M4F0JwMQgablL1Ir+PWuYK0O+IZ9U4iw5CawMR8X2yjPisfF+d
k84OwvpY6T3wRiXHzGEPKItF65Y84DvWNgXJfMItCBlfk5wHMJeB7kN0Dqeq
aseBIkc5U1UNXnP5qbhcg9jRRCNmOQetjQRjZti7mDce0u/R25zEekijoXT5
U4DeKxMjI+b5nesaAga3Q06A6zUxXVRnPP5vdMGMCE/oSp8HL//pgeR98J9z
ooGH59ctx98FiPQByY7PTytyc3rXGA5AzjXBo7cSbnVs0RoUjDJjE/5mu0m6
h561QVFbqMJs1E5FYUaICOiOWH39/RCB91d844Mdi74NnZtygNlYw+B9aoVw
WjWi7o7chnIeCehJYiEtQFELbIayAeYZKDXhdNTvExKJydpZKXMGnLgLHrOV
+knvCWPRPqRqKffLx5WaldXOj2nDZ70jAyhTUL1vMVp6lfwS719844QwIGrW
4GXa/YcPnMHVftJcbFykeqTw1yBo21aRYqeyfVfiV9Y0xTdRjPicvkLUQ3VT
dUZvl2nZDXxMQwDyZrZrLFLZSFL9fky7ZFqrCKMkrJ/1MeeLDjUw4Q9TLluo
yUOyVMA8Et3Et2IJzjJJ0I2/H7Zlto0iyBRHr2HxRbgkS1aU+q12HY/IXXU0
MlIizK9fho6CoHZu5DnCnKJ1FILS/yujmWv6Oflok3/4XibP9BRyqhjMxsm9
gWpApa1uTcky7UUnxttztSfJ9FhMmYXiIJ65tczd++/IKnDsp3AgAkUG1eET
96lidRsPXRNhJ+NsvuVtystSNtm+hHt+zoPmkQA3g6mDfEPEfvuZbfHBpeDW
tFyKs8eH3CuvuAwH3tx/xj6T5WKVI7mIVzSgNJIFsCg4CNvgp3UtAU+8e2ba
GkfXHowsfKg/F9cgnzq4qtMeEnZ9G0DV4uGRQ6l5EHZaze1LIxejDsQOw3ds
cIxfIqFO8V60TxDQbAUztcypXBBFujYuJSKNAZ36rurMcZfgLoqqfwLx72lB
0gPQ9a29FNF9ER/6bMY7kaKpSh0RIwMVPURDfWqo0uJd11Okn3tXvJhX6fEj
cwOHUia2+XH0P5e3smCWMyeD4jUN4pXwGqcAu3J06NYPGnWO/CEkVHzdYcAl
+hT5w842WgeSoEHp/joqLVSbZplfm4Wq7WpmhRPeR2IOIdNSJEUeDSXJZSHB
XH7DOlcBVC6HTD7l6wI0j6B6t87RL4hbkLMVc9EPDBfr98xalFVi7tUtxTjx
VpBLPNvDA/RpeGDOSSaYzk8c0uO3G28ooT0YHgggRPPkPuQXSdL17o76j5x8
8yDDbYm5J4fyLcLChC2OsWMw0Ka2o9D+LWS5ZwxmOGyZ1KtmuajCXQgHL/Er
8dJKUKlET8DjPDVh2dy99BtdDE2OE/TxPZ5lWmJDKBJ2GupcAzxdz098vF2u
wuMK9bfmI0h6WLjIF0M7GatnkXXeKVxLiD3Q/Oq6j9gIlIzUfQOsC4i+8HO1
XrewSJIIuyxV7xgMZLDHNeK7zJrBb8qyFtTpEvXcoYNGZwR5sVl6Qx3wl9de
tuXG30ZG/BGitEsgio77KBZe2aPOz4bxXJXO2F5zbpRY/yh8DWf+CytZseVJ
JqtgKpZVb2JGGhtN8iMErloIzyxl2TiSM2WprsT/ObDqyWWyVzrndnwFVjox
nsDvuNgNJfFVkFur2MLvxLFDtTBebdUp0kp510X9jJVLbqB5T6CBeP+dHIh1
qEVBXSa6vk/rEZrK4nIC8k3uZ4uBeWn0EDHmM/cb86Zn8JZt7VSYIkNIey/6
gHLfYabOO85DLLLoDKriGsqh6MywMIYIQxoPYqwdSTkEnRpj7ngQN2/19xEs
r1abrofj/1xrei7tBXx3JoFqXwvWF+tyCvKaf98j9A9qovTnO/tsahWYU5Xg
oRQEqSVG7krWApQBN3bytrz5Q9fMcBf1gpMHcZD3DXJOeB9Cvnk75wafJp7X
s0BOkKfUfAUq11xwQzs6HzytN0WWncDuj6z7hoTm+g5Ur9KHVh6DlFPQV0MF
kSkweSYVXsrC0/2BitAW9iXHuQvEJLfBJH7ZIYrGutbAB2p/SqjgBFICXlL7
skE29JkJ/DnPQ8NTfCW9V9kOInRdg1O9fmlwGHmkyrV/+4rkeJTrhShXimM/
J1dQhdj4BxZdtj4yqseOVQpgFav3cNfNMxIF5VhIOS+o3CaxlqNz2KTljmJ7
GXBOoWaTa1H4Xa/ENIz9uPs3reG4UdNqg+i+OfiOEfuH3vh7dHLDyT9yulCj
x6DTEEn71nQPKOx7Uz7MYRL4ttyUvHMkgL1SsF6yPruZ5f4r8SAhD9uDe+60
bLA4uN93+MFYTjg3p747fvgghmIILwmCSqYV6ZP5+B8TybkipkRt0sRnwnOS
Bvf4NtarXVBMoT9K24U8Hs2r9RsbTHaFDikC/21z00r7NEwkIYDx8JdNljG0
AaVnsu2qknrLRGqRbK5pysDlkTW9nxAxLzNDp56bBwjeqW27H4KsvuLcgKBo
TV4bwc0X9X4cBkjcY1q6Mld3xmirjmfYJYa6JrYdzVPb1Y+U8HezQ2tjMIPQ
JKqt/lQepK/ZBfxYBqR0Vwmc87jh0acG0+AePVjPxMkmQy+wy4HqnUeIJcKn
HVFAHMJ9B0TYBSL8JOohlVMjrIiH5IM8LEzoYnHcbMfccQT5H2emvB41WW4w
CqMvN4VrUxeXqLSOU0jCp2gCaY9F79Y3QmfPbRKKJAytG9tfjzos4MbsrcdK
PnF+9cGvr+iZINnq05dyCSPAgiIHlWkaP5utKH/gYAKVVOKWYsvOip2QyIyP
v5NdWHPwxoUjTj2OOjaUInh+6BK86P3ByTbSGXAQJ9y+XQp9ysbup8Nz+lbK
t0iU6EQp/Pu+JldpRYExCq/YJjU1GxKCzvmgNMphx3FjsFAFEyh7oN2tfLJ7
qgclpaHQM+P9X68CiuoYQmgalawNgAouFqSuXyq+8tgdEfmfHez+48oKnJZR
oMxrfIcHqiL10cm9ts3Jf/v5yJ3ap1V5rQZtKloSpqeQhlEQc15pGhR1HNwx
AD002Y0NfvZv9GRlKV+FqBL8/ZEocWsjPH/DzguILynoP7whglC7OFBFwlfF
I+RVICHK1WihkuAFCFxFGGXQOpFK+Dl7MafU08dQKq6OssOa+WvTuQ9AvHYy
zV7JZ3jWEhRgtzb/tFfVBNOeHVdiAJ81tu5+eUESBjCLm56szbL+AXO1nA7b
HBj3UZMWjs0Rfc3f/ynd5pVM3GAnLEG6GRrjY78U6CKTUH00YDoJXkU/3X5l
a5MftGBUttBR0OGvsK12xmlqizqi8yXd70HjhHFMPD+j2priIbnO6JKHH8pg
dc+fLlNxnxR7rfzvTUZHZg4SYzjwtUz0wudR90BrfmkGFSMC8G+T46x9EEt3
DxSYQsV6LDcnjFGgHkrehpnVPukTQRrvAdlYykIkpR3USsBtaxgkC5shSimp
xn9FGoZuM5xBqqDE1IENnq3sOPQ0H3FKcVuUMvDbf87dOpDGJDRB6r8TJpzA
80jB7Gac7mrEO5gctKdqyXVosuCz9vJJJAKro61d/gJh4vw/8/ss+L9EBHup
1ta5yF4CMyXi4Qm64DnS8Cc5Xk8S/lsujRrlzyAw0C0WlI6v6mRzbrjQH568
U2K/S1RwJpTUJZhKu+R6UJ6LQCyz+9k2gNeSdKzX20u/sXkKPfl+aJRboNED
QEs9I2TEYVlmTr2n9KIRtVutFMYDanA71ZzIwgOjzOZkZFIFXjRPXc7uP4gB
z9mU/rffOmAPCB/xRccEF/pIKVFNUqdyv2Yk/loPdKhxFpUk0OXpnE9g+gQz
2jGTaI7EFJk5Ifj+5uvXj57i7r39daaxKyWaZIdoXgPZ9mCTuhEQB4eLFJ7G
QJTbSVuOw8U+LcoGL5D+jMjnY78W7dU1dJm6ZE1zsEc8by7LcngKlKDxI2vI
90iS1q7XVOO6EajFs56EThpbRGP3/Is0A/ybP0WX6Vycnh//aKcpuxW2zZ74
ICtsfI6IjRZXikZG0Vkc2WBnQdElGvcyrkuoifISasWpqGGqaQ4r97cVHLfn
ReQPgXrW/ZUv8Fb7uWHIlxzF0EhP7+Qeus2xMm12Iws+R7YoKwUNif/R+DS5
r0CMLR8FrrM2TEQh2c3b60yIh9UDbZ4TA1lB2EjqJSJNsU2ELsRSJpxKq0OE
4bFi1ySXo2D4j7nhGZmBoA0pgEsacAYhkCSGQrsb2u6M4m/BJKYMmaNGlhMP
VRlDDC2ceYOD9e85KuDd+H/a2rI/vESMpi8WoeDPc5uWP5Q4YLcCdoBAvzxR
f5jczmrEZvBjUiCVfXmLh+jHseQ/EKp1/zjza1k+tN5OxF0OLiMRdrdq1+IB
AtUXhZrm8tfvAPCV00n8CVIbhPHaU77lfQBw6PsbFMi+hpbuA0cSplD8fXxs
BmoFGrsT7FsKaw9V+bzDQ1QDzN67OkPmyrEUjlmwr1zPiwWJxXOtTXlmwC6z
1trFldEBdJv3l2cMoVn+oOo4VQCGpFE6FmA575+a1JaIRCA4JOjE6K3K4zIb
6LleXLBDkcPTaPnyT69S2oykUnGO4YKYFX7w6dHS2pmCyYmrpZEr7oT14aEZ
z0PMxw1ppXkztlma+vSYcEsK7mWsHyK2Wn11al7jteN8Tio4gAq4BvkKao+i
JAJ9UCj2jaeKUjka+EDKVBGkQVu4vEVAy1Rud1xJzCQVaSqevkHOUUp6rvWt
U4Wid1U4FUH5idBneoFi8pqIlnN5xeu9icW0JZFYos5HBYay05W3FssjfZ3T
hmzhgm/UDwSuP3KZWJyFUOPLGYeYDXuSPepbsCidm5uXb+Rsq8kn1ur7Am3q
OhwhNMtYwoRsZ237FCm+4Vz71StRWq3SF38ajP/7KbnR2urvbtdZDm3HPhtZ
ESe87rSxZVToriYwuCPujnINibdU/ncu2Z0aAQvNoIIlbQCLD28sZ0fO//gi
+hDS9GcFiUhW4/AXFbvehBfIDOoxb4VQKVFEX3i4tcPcRYzOzSQ7UPXXG9yR
Qa9OBb7mDOtLCVtP7jlmPSMmrKaiAciV5VsFsDLflnkGrqi4U1+ISEg6ecWZ
7KbvbBGq+3xZ8m2Q9lP6BIggkE9pu9ulfVWPvRnXKNKnSWLZIXbWnbCXmIyR
xqpa+ZGM5Z7LUSZmDvjhL+jZijTZd5J/cU41gw9iUhPMw3VmQ211UJHUdML1
Q6aiWSQvGkHebbd7stXOwhZtvAd3VOz5uXXe/o7BCheFZssCVd4D5rq77p6L
FA43fCU9An+MynUFdjCGGB+so/XjPFK3NI+FoJm5cQDpErXqem2foWX/oVl7
POmzDplZpwDs5Z2bC/Q++10hUtNYuL/iJ9KwrtYxEkiXOEJAQrp6TSVMZIZu
Ht/OjWf+9VV3eekZKmCK7pT1mteIs2nK1WKP9scEPU2kDAqfrA7TXbuVYgWx
0dky/tLtm3E8oU19UaiQBayDRlT9NbhmBCd8Rd+GBIyf/ySdRGCuVWkpPCBQ
/8uO5Jp0dU+nDz68uyFctwoJRRM3x9xiqQuuojt5NmPxtcEX6XomNH5YDZ7Q
Xl8HnZ/dYdSjhEid+367KWkWuBEKuSNaGnr4Nk113C8f0URWjBVxsXcV/IKK
XRiettw3DpWEIzhVmUDdcsAP7o/V5C98dRl260ERQsqPH6YrtT9Fxpkxmw5O
oYCS/XnKTJwS+IgiSJ7nJEGwKhxidIoyPtGTlnmZXg1MYRqjDtJpjUb5DYJE
050uoZgEsKFkD0eSHuKr7vSU8Q7L9CoHpPcphugp2PU4hzCBaeNtpEgXhpX5
4eZcS9/R/2JMtNc5gYxHKf8CmfEN1+1jDv+SGrQFZ9ZiTmTONw8jSIK07LbQ
yBopfdQlLNhvJNzCvV0hBNb4b3jbyQnmBijCweSPDzI/kUZR/dQJfv4Jm4Vr
EQz1+uf+QyjkQb/rzhLg7F/2aPdq7zelj7WyvSq3q339Mfb+aSI8EjQvVGgb
SmSs5xsIzC8ioS593Ud+2S1SmH3HeNK0mIdAn9Ozr3DVqfpsnA2JJSw5Wv78
012jLpq7qQNZn/1SKJviYDpvWNUGHmXYeyl8vyXufVUXzO2S+P8w9vkvzwUO
bkVysX6d9uykwZzVovN2rhYVvpoMvvUvR9xnAtOew37CQaz97tGitlkA9hh4
Xn1rfBDs+en27i5N8nAdq2yd0Z+Nmdz1uIv9BklYYkJp+k8MRke9JsEPxLDV
eTFmxCUhx/NG2M4prMMqk0NS2SbUKXENTkCtBSelwmRyBZ3ZnDtVvWrbF4us
RDKX5BaVUcz0R/N1B22bdqbW2qfva5fSgBlW8YPVio5Q3chkPaZEkQy0fpmd
ft8tREO8PjFc7BW8JoIL+RTudvo7p6H3oiyqZoVIEeof03OtVfp9pMMTdS+w
FZQ0VU/3Q1tVnO4UG4BfpM1OJgZoDQfVeRAJIZGAdiCmQC/XdS1V3ejwf7AT
+dBF44i6bEeFN/keXNS5yn/pjbj8icKlNnCpwpsTCmkfrdfKZgkJSu5kLBHl
A6PRBiwNUOAOPG4KoA17pb3Qz0aBbT6Qy21syCRUg6PoeL9C6CMJ5fhnCpGh
MVuRhCFKjCmkKnbho8IOQv12MmyHtaJP4PVem6rYCcvYHhm2kInNDSluVqj8
04e8VIa62bHPQqpuO30jAWlqd2/5wODtFEBiOZxuivq5GrfDtOgjUMS7Skpx
KrAcLDy5kODXwTwJ5ZxLPR4oaZRFRm75mVzH6PWtzzFDBPH5XMxMuxC1Uiu3
hBmfrMDvLnR9MXSaUQf6CZofhlfLiaRpdp4DXyRryyBdnEFV2SdN9nH88wKT
84iMHfzj0vutENhKH0ZkyQU8WxoimePtCrHTeK4kRJ57FM2EwzSvSGfvFybk
cslDW9Huv7LoleYsNteuM8SA7YF8qXop42gF6Su9kVBnAKnHdB9F3I7EEwcw
cAPAmRn+lKHqUHzRTdqqqdqBC1sjmP5yqtkQweKQfd2Jl3fiyyumC8R4GVsH
33spoYukm9z2UI39ZNoMJmQCAL6dum+ehguZpPtXTS2usvNEphqHcSQc4zIn
RqtDlXFzHsrvrTQxR6gLV/UwlJvo+zsC9/fNCeMF74xfYdt306KtTjs+bnmo
zdLC8AvAnT9o4BYD0yhxp21/lt9GUM+e+DJ3N7oB7VrtVH7LmgjdL6GJeXhB
YXwyBMoUOylA1mbwHIzUDpHNfv4VWKkB/qEZ9J2p7OFPCEhjwngZJzhU9pzp
XEYmH0+2/KTufuSk0bzsm6997lrJPl/Bo/CbfnVVzAM4IXaZXMoMKT5I+4ON
tn/acpb1zcXQTK2FXBKGbHSiBkDHpp/RgeZBduaYnBGC8/SwW2HKA55DnoBx
IPkpWi/oJqvLPO7SBhznbBBmKlFWY2ATacMNVlcDz61Psgw+oKNgH0ZBD8s8
O/4mG0jTqiQ2on1FtYdiq28MGFX3qAHiEggve585i1af2q9IJeE5CYyYqkOw
d7gwz/SXSGm/DOO6mdvI0P5NTJgfMv1SideW1jLWsCKB+xz3jhIev3wnPEVf
SMAz1vXMbXpGPjkQUlA3d4ksDx1mB1CwmhrJK3lUuDQP10gehMHotNaO9CtJ
XZqqjYi4pE88dMeg77SrQLbnNuRm8kNf0tj0k7aYBk30hP2EvAY6Dj/v2wTV
35lmJciZkzGyU63m13XjNAGq2QeZ6fcuhERjItj5wjjjmIjhhlDgZSDiGIAG
Sl1poD8AS0X9MPyjV5LMI6Y6sEM1yXeRdw28QoJ2/u/PTexRApnpKD5alJiO
P5D8t6xDfWd4mTa0U0kdq3t1YMtUsx6tIrwKCU9VaKWdcqqYW4H/DoQwZrd8
NOLoMOmSoA7GZGvPMdQs5X/ShMrbBarerSDMO9Q04tdKm4W3hX/CBVMah0Hm
hhIz7YM7MUHuZUsDsbZhyUCzz3qdvWBOn+RyXfPZYKKtlK0EnLUfhLv/1MVd
PbKZQ+PPLrEmDIYkQGENWG/LwgZTOY6yxPusDwNhw7KPIN/n9WfIJ3pkeWoM
4JdvwOvBaN+eT58FZu0xObrr5xzHKn3nLV6nYc10/B112T3dcBJk8idPQdSv
Qw5uqBj/C7Q29RQz0hMirVs9BG7RRnIOUWjts7mA8O52Be6FOFULThfmGPYo
LXITlxP6zmDn5ljKpnY9FUbdNrwcVhNRaQe//N6zseqzU39Z0QiBp0fjzeud
Onw5sXC8nyqNSGpvgrlV/0PpyQBLtdEYLp6sKfjuiCujx6SaTinVYvasXK1E
zdxbs6Su/GJCsFsnFWMi53/Ly7KCW4GLEjF4f84gcywiMa1uBFM7EHchv7bF
fLNABI8uiIcnF4qLLZfbcbPa6Y06m3Lb0Xkc9OZwAKYvKYsr+KDjJ4jM+NI1
x7FVJ2QQD2x1fUOPXMEgBqmD6ZecnQjQazTa7YRfstUHTMeqfYPxUt0x4B1V
dWaVH/Ai+MuZl1e1oqG36yrj2phiiw3Uzbs3G3WBUWAGqzUe4V10DN/dwc99
pgrDgB2/XzYYpWRJKbMtfMgKGtY571W3E3oMkxxcOgMbszyzE0k/lqRnz4U3
rDWWYJ2wuGawifFwtgLp+kDXKleo4d5pSw5AeUj/wFcQ9KopHbIclAc3VqA1
il6neinPLNcPs4nhHpkYlpWZA/Tt3p8/3m50VA5uR/pXzR+QUpoE2PEjPWEM
7j0hX9EXaDuMlLMPB5Xmj9HbfgmFr1dUVs7hyE5joZqqYjVAWp52av3s23qD
s18DoWoZiD8bDgQmY+qufcgguaLQIhIa3IFo0Y5LjCzTkevaqOVKYcqdG6Fx
Hqf2Amf0OyHRzmbhrf1BH3CpQsBpF+fZHI95czW/nEI3XGHcbD5ubBR3d5Jl
Q2z/rSX74eWSRFHEiJcpgvYlRc6N6QkDenA6fHvFsdA5y/Y+fUSxxZS/WCY9
gbuQTswtN4VjlVcan+9CrfB6karsQXpzS4Xqm00fTflqgVdTMhn1xuwR223O
a0CxPhdX3npDn7xL6pKJCOEbCFf2l7fmbCFjVSWyg/9MfCNMve0g98shOrjX
WfYV4PSp99mjBpPbjIJCvYGPdWnl0werJ9KQYJY88ALqWUooq8WbZny9EXa4
Aug2yJCEsW5PwXgrt9ilRhs9ymPmtTNtru+MjUg2t7Ihc7Dmwu8dppofvwR0
qM7vh0wLdgCsGpXcSuWT45HcAT5UUpIcSg5DH03zIevPVvqQBdgoBw3iRoNX
vtw8IyLxGxuvULeLXelhmZw+p5Nj+HO6mPRGn62y9RyzdBuGgvb6v6/slWmx
04CeQKvHnSKo6RLcOUJCE/WwcgB4kGqdz7RrXEHoOpFUeK4qs34TyY5eS4Ip
ZrQoFhNg0gPrqOmQHHGVQKyGVU26Q2TRU/AuB7/Ez0ZZ1t1Gll0Hx4ll0GFu
TKfaRYoozS1jvlZl/JBkUREwzi+b8NLP0RXENOK5U8QDbvqUpXqksHe3gugO
I1KWVIEGk+Uq/zDx4lChJCzwHet4zZzHyAOUoi3II20PWqkFEwHSWeaQpOkD
oRZn5pW1INW4gHIlCgSeq860flXHoi4cSTYCdvL6bJ64WOYS6Y/Kb3LC7ikl
L/hQ30Ae0/USlzk+HkOTl54tNmzeAAYXvTB5yWJOr60flb7pes3Gej2Dg0KH
mQQbPRMXqbwckQKWzyJGWPT0PoR0W1n8ZWsPn7G1gLt2wsuq+VNIUkWcaS0c
2oSq/59C1goNAhCKy7Y+zE7xLkoqUN10xoLEqf43Vcvbur7P7qX9lkVBlVLg
FVoqFghDH1ukGkhdZuhpBAslInW1hmCJQvFwOmInnS8k7ce9tIbzl55KCjEw
Z6MRbaX0+B5bF1aEpTqULaigmCzL6mMp8cM+5KiWv8YmreWx+rCDzrcnA0/R
QmcB+GKyf3cwiDzMxqTmYHkN2fsrWoKsMqKAtICj9oRDKbF1OpwkpZ3vLRdL
XKGtgHEEGOcw7/snwjJS5TUubZgL6xtTFsiOWAttCRhnLkVjPMJ3a2egRFHb
KEkJeafpl+md1du6/EaKUec+y5a6kOC47krE8Dhclzpl9k+Us/+vw6tNuVNL
LWvJ+rgcQHovUPX6D6mGbQSb7Neo6hBP78FbTsUuldGfKMol5uoillFLlDc2
1Ar5fMgmliglmbhdEClSsY/gRcgUkz4pm52SqZMEd4CU6rFDTjSn5ugqPo5s
mh66nw88hWKzf4nW3ry5yatDeEGxHgfSIcIiTEefn38RDIoLDQQQFVdwAXfb
s6WXwtIhgNSKuxtpjKylB9//7kmii2QcduJhMnh6SBiosI66TZLPjIYvG4zs
GHJWtg4ecxSA4ASxtkxjz1na5QQCMVjnQh/0hg86TF9aOZQOfSDIVyWTcPAF
uXeUr5RYruHUn0d3lyQvNwd0a7Xck2iPv+tBn9EOlTei/B8S5xtwGxe3Hk7s
7VvroCWMRV5WMlm4WQzH3hKuJ2+weRerNV1w9g5l6GZol+RazuvnGGlHDXmS
bdDlJ+1PAzcB+PKR8/wCxuE6q8UoE1LafBLtNaT09CIMtMka5Kni6tz51qBE
CQ+XUpIpqrlxX1TEtLTl1v9+ilxo/+yv2PjNSmePrHgFA1BnCEO9+CyZuLct
dLHEsHkZlW6gPUKKZNzmQjm0PZ2nbZGkYTLQkE1j8tUrp0d+kFIihlMk/UsW
HiW+R+H9MkwaE7MrUSAp/upXTbnvToVGQlIjrC7yHil/sLDWV0wkLJdQvozR
zGCy9HEwzTi9YE9YDDv1qUDQf/G2IAylFxTARA3TIyi/E+R8pHxERjDEtGfh
gj8xcBqebfghMrWr7QhYD2qAiMHZdjYvXO396l5ndPBLboRg4iLzJ9Q26T2g
S5vhioIaApK3Ac7WTGzt0QE7eiZeKEmMpXqCOS0KhBW3J253dU1ukdrnDFV6
XoapTmyuYpHr1vzNlK9zoG3nZjL04tOMwAfYG49e+twh1RaBjWeZeB9fOdOC
9C00k+LTHFkCw9OsF+jXbe1PNTei3M9bQ5XNkshaPhOr8TkQ/gbRbm9ShFVY
+Ce13Ao1dZBaWyX22oudGOO5irEeSKwsG+3EH7GXKsuxCWjXI2I8e4kbFTXs
Bdo2QZVknjFXutxYqehNMZpmTQRmPDDHaOKb94Z+RGwMzZCtYsq7/LN9yCRR
3q+FLCHxVETX/K4CcBgQE1T6IDy5wUWZqS/pgSxA9FfIjxnI/CA4ddBVKg8A
vIt1epsP+8IKsE0TNUS9JAM+h7LYebLQLAdcfj+SuAZyt38nIHZmXN9MiXAq
PqLB/eVPKuoim2hR8pwktvThuUeXcnkguhetFYGIF+Waq+aoDQ6u4R3THoZn
wGemVSv6kPZ/XD7QhETlRCq8VONSB4carjRAUBQgzpmZaZagrTQ2hbwfGFRX
vaKwzEcotZecGFmnc8wvIJ9yLFtffzZjQU+/tFQUDVgbFqhn+7Hy3mpIbAoW
h2rHMjdbEoSo3vFTVs6750FfdYATOjPQ9NSsl/WqpphgeK0yistTolEzcztf
FZ2Z2olXWA834h4OKfqiKjOWWkkf/3CTHYCORHQPJJqFdCJBCWz2WemA9Dqu
Q8O95nfqwA6SHFLMGJeyb1HubeVdX3Jpys+XEFZXXc96uGIl95Xcj/RgDVg8
io8HZLa0XWYTRWybP94SxNCvq06u/qgExJk7viC6IroOVWeaHk8YmtvUkh7z
4LsAi/ZkPlUtVNdR7kmU2BR4lw/JDLKCBS2XlfYiUhU/X8W4+oLdLOR03pMK
WQLCeS3yikLEHxlCRoKq39tJDZ5WykvqAesjiGKa3+1u717JkxcrwbgOL448
+ogRZgz9PX9wxPt7hcOFknWUq9solD9OPH5VbsucE+fYVxkoXDEZ7Dw4RsS2
TAvAaWTrF8HR2gXH3Zdvwq01wJJnzLxIFznWgb+J2ClsNb/2u/Sku5z0Lnce
rrHMZ464jT0UUoG9kzdNqzbOHEO9ypVTtRGyjqqCejw4Sj3z3sn6VIROBmaA
6Q5Ne5YShHyXzoA1XfhAYrkx6vJsDnmF8EUKRkX1MvuWANuL/vgPYwuT7T0M
i3qV52i0h+oa1I8+XuPCE+YRogSN2v4qarwqUigVZs/eIn+N0MDm+zRynisQ
ZiMGdusAk3L69XTwDt8Db1890scHKCJ33cMunOkfqe/509iCew9ueJT6PvsU
vP4wfcvv1hue9FPFpUH5p80awkVq0WsaJ4gBvO67+wDG6pQQY+tAbrXv3X17
lgCibOsCTeuBiwcIKN+vZ1LLkkFm6/G56Z5IYtXX/wptTd4TZ1M/31kKFo5n
8ENdVewZoMmlsfFo382USGFBITNS6iplGCpDtkUiLh5rq9a6j28VejOgzS6t
sddvYCvqfKNg1HzUYUD+Vtzrt7ibb4Q1eWjs/9ZyoeyFGvblhpMt6nA0amHM
ZffXPcVN47roiGhpsTdUrRGq5IH/Oegswjh4SMlEfeM9Nw99GgMxn6FZFsEI
UwgaiXe4aXybzniThxJvrvbVcyJZsQbS2+MOQSmwF7VgyFrXcEgwOztbtm3c
/rjz3qp/Zj7JI+05ejFChLnwUj4HypKPZHeIMkCIFDzLMlT00RGxOEIMd3xh
D+0jPUQKfOhf7HgrwQniAgt5cFUBYqC+64SXJAusHgjqo0srdIzCVPnvzn1i
Xxz49fuCpgTJsQV+Jm2RlwWjh/RdrpQqkmOLU9rO/FGtS35CMgRgnlq75S0P
IdNk2+Bi4gy8frMkTqXhGhx96iOaz6XD18+VeU3+HviE9cZz94dyud3IXP5D
LvYpu07kHIm4yP/5qwBXyrHG99WXd34j0VvDcS//fZILVwP5KXUQKcyEyxWq
6f5BJgtzjnxOF04QGloeKV17mLhp1rOOVamJHduMw9zI7zeGTDfAZqM6VTSn
97+TYnkwWCJ1Vgzh42zCXkdMt/8z4bLWuLwGgCrr5IIct987dGCOl9YAEW4w
bW1qp00xZWycUuxKeS8VYiqfdnNVftjOFnnM9LV/lv3fWq3nv94+Odw33+EF
vvllDhGH+fv2H/llZYXrgGXvzaLnyLNqvunDeaNiif4AF0PhH2Swp70Y6f7N
hr2OwuraQO/kjqx0AvCzp70Tjry59mAs1VreNTFkGVeDBWUsS56eggaSYZF3
H4rqAdj76PAlYx4apoQK6tPb91gFZROUfY/sKFZ1wa+WrAzbE/oOGbhU6P9P
RUCpR/RVmLtZ6SBjrRsxvjij+jKNbSIX0p09jYM+KagUkLz6lb3m6QZfXS29
+4aAimI3bRxJaUmv5NW5B4AGhzltvoEHlF8W5uYHjt2Pb7J8lv503qSCmADd
5uJrm79purrsUHboTl0yBr+fA2GmAD+hrPTsvbMzQpLztXbAFdspCfpgUECA
ixHj4KUsCNtrCm7cygTjACwGaSjBmQmbO93OB67hDA49TRfsKtmz8ZoBpNap
KLIBTREAavE51dY25FUtfNsI+nbANQUMTmG7NLPKbRVoC3X21tF/3Hj3hvOi
zfrImzBlYvxf2nfN40ePFoGpm2lQ89mRqrvtFdCv8SKwGRaNL0ZayZOl08uF
L8RKlg3Ix5IpdL8uuu22wp4nA037vyJs1F1PJd5hdnYqMvY0KgX2ReyV8Gl+
1MdfA+2yYvhYCzPfTDpuqxRYWDQyUXkZkxCgW6xpev8Jw/o9xNykIuJMBp5B
9XZjn3/QTj+hbUXQuSdY/EHUmYPo1cY7McfAUZC5J0ooeDu9g/1xtPjuN46L
bMf5MBm2KhfjLdsjS3EdCAuQMKDgGMfxwShy4s5Iqhi3v0Nfj08XmiI0+LQM
E//mB2PaCPILOVW/qblYT3XR/VUr82t6qwpTbZChlWgkOghzeObSUY7Nk3r5
QED2yhQBJ8rCWluoIjrXfHt9UcMe/Aa0krS6DHHK0G4y04VkwLHlbOm7g82/
/+RAkNKjW2A6eRymhU5m2q0xkHHy53lQoQKEL/Lvi5tyEhkCpVb9to0tmGie
4mpv0N9s4pufLA2lY/Wxqp3E0c116D5KFQtVgL1V/Pvce0SzN+6pQ39IqkS0
cIVMNhQ0oW+3RfrtLqC8aZ35uOtKJJKZUCQR7osfCC2/G91cw8/vesGJVcpy
k6vhtlPoKz2wDyQ8lOmkSi6ar7EmyLeO88wKZzD94lm9w49QCiDcCuK2ynNk
HpzGmtp6re03mk/9vz5Ts7SaUGbZbXzGNtlOpNCfD0ETgl4PdMyloPG7De3C
zYY52bFcjHfDvZaj70cRlTxUH2wdOQ76vJqdN0HFSDGWYF3XgNjdRBrdRdd+
6emCJcojItB45Nh5MY5woehxaTRhFWmUB39Jy9P2AzUbe3AcA7IWLC2I2wnM
CZ3cElkAwtxfovorpY3EIkGUL1yOs+XvJzmE8KbsY/5KvrUdiVwcrX3Qfulh
NZQNZMAWOplq2KFtbIDrJiNdI7sRmQwCDXXqp26Cu8vo5j9TwLQtGA6Jfqiq
bcIzr+Y39ZYb68J3Kc5yIop65LdLW0ycxEFNiFIgzVnVYzG54kIg0q7atotQ
3ppEYJhZCrLSXLZJjMIR7c+UKW53gK5lzmxc2eykCDE2++Z/TDTNck+qkQS+
jViL8OL/rcs6ALQEKRxewMLNs2K+Ta6l8Rs+sKXuunm07W3aZ7S3zXfrK3Nn
dwehDB97yf/7qskttNQ9DKvDS0kdieP97F/R5e8kYCoBueCT2C96ZePwPf99
8Ih1/he0CvE9UVIOOMBmXfTNoCy08V2Soi2916E6aGf9X8UY0Y25qlH6DVrE
hiU/6nuhZ0QcS6TzMYQQ+hGplF5fce3Ti1VzVgCosVjSla1gTEylVU2ieEPt
COY49PQ11/KvotcQr+xZ6w0aCntL6/VHs20NYTuPVP/0Sp0BNNpaaJSWgh1a
wNSEpDucOdD8BwQ1pfn6V5Z4LUyNYv5wo6cUmFRHjXt1mC5vTBcI0uqOeYDk
vL15BxQ9B49RLkN8xvzu6QngVvvrZD7HS0cFmlnlJNIaRIEXZUd0cuN7G5GR
SWHIaoCBkgdbeOthQzUk70cd5Xv1sHs4xU8bK/+YH9iHkPRYrYQIOVxm7d67
UzDXfwSMPaqDFJTV6BcnG9CZadxpjTTVP3aGANqlTRgC5m4QUd6I4CEnOCkx
j6+lmzB+/0w8kjGDDuXeYz7AaZub5c2wPH+DePtegMIBGo076VZNGdGg+XBQ
cJeuicbb5KeC3WX+5CqfRLTQo2e6JWo4IYnBvuWsM9M4TMOJi1F4CvGdzrA6
jt7Qc+uOliuhwcMgXB/XK7h3gdVewWaM9JdJPwwMYYugYHLANd1fx7WZUfTS
zKf71D4C106Ljy4zNc46VFKhejJzC5J1m2m8TLVtmoWKVrhsa4/pOXnbrG+S
3lJtTtu0/cVReIoZzLR+MdvITohDQhFl35QE37hyLPaGVEj2WYDMMYuJXyGy
abMHVy4l9EMiEsL+9kApAfogrXbKTTdUWNdZHTrIPObzVqkNj1qlHf4CUCV/
LVad35KWKAR8Zop4xAqmW1dcnwcneLLnvQjxpi9ZAOsZrCl7FqNihHpujvVv
JUvOVlFAydfgbP2QeQkJ0k6ZIboNNtuH96KdO0FeGisqV84u5UY8hlN2ze+w
9UpTZglv+7Pi1+O8Jbv6vKqlGyXV0YuZdV8hpqNf03lQmwxesFglBuBzeV4P
vXAL0CbLz/G6LZF3OsmmrYa7a+xixS3s1zj5bj7RVYpeT6KQ3QKRxmH0FyQl
wTps3UV78wyNSGmb+F7J7jiOGT571GZm6ZqTTYTpeglDsryfNHP+8Ci6Qg0y
by+fNKEeLEqMG5fyQY8NDO+ybpMsuk/GimldiCXYAxek+KB2prMUeruLnjAU
xgeW3BT1/bEYEBud5EE1PDCUFC0AT9KRhXpGfRePzt+Ar3e/oG69P+oQ1GM8
iDLG7r9CRfKnk/O0eL6EpsdTcwfvXCveC6D0xpE4wMt2C6mfFPVdNxBl0Z9J
NJeYGuPtYRPjhH8zd4/RmlIFong7c6YeE6Xlp6LhZ1eYp/1JJ/bzKj49F+Bk
rFNT/i7fwzlVG3O93a6AZJF/5m8msJEK5dRfjQAJYogInFFCKCdyFPr2+Q9t
ldtQCpwr5z3vRr+qcto48irn1qQKIUYbQS2NZFvyLnzLk57j7f1vzU0jmdlB
Wja0//vALJZ0VeupyK4yMqFiHWs/4LAJ+mp3JPmotzzU03p5drdnqDzZPBvM
Qw6iXK3XwgBX+rNnBC55cGX7KXSig6Sd0zZGWEnowQfPEukopWb/oKWfUsA+
eFYXdd9hX4iXtaHR0iX6z5tY6C4qcG0H+gXya3WMRFg0UVSF1DAiNZGZH8fv
nwrxNh68mQkj3BHbcdvSh8H/yjNphJ29r6cVwUAGpKHlTFubQ75XE0cgi/wa
dH+DbcPNFUp5DteKHbim4f+LZdMQlVKpja1PIFdNdCHfHmw4lsTHclJkpP58
WAQMQvuk2tNgdLHFLtUPVcqO06Zk2jSe09Jgx16U/d7Z7W/S8QR4BzYT39OC
1I12Ys+1BfQuLfWqEWxowzxgmMW+JgQ4YNWz6nD4CfKllg9JlLB82IShUbB8
XJqFaTyPpg2T1dpwpKeAbJ6G2ugSqUfChufv1aWUCpGakDo2yBwtitKq2aKP
kav/odyTs7+fDS1hnKUO8FFF4YfbJ0uC9Nds9Z5I4Gvvu4bMPhWhcAK4Is2W
e1Rm4o0SKtnJ7ALDTfkUtnWTKNLn0nCAOLXT3USSoSEU3amF5/pcmEWfphrz
wAq8Qf1PZCmlCHOZl17pRRGiIqt9S5V70XSWayJOz50u9BSu3tZ1KTGSFUWn
vbT/DxeQt1LOuP4GWGxkJIDxbM4QzZCCLMVlbwsHgl1c9WhhqDwYPp0sGa4n
YxzUuJwbYxDTyjhpY1VMgNomA2+zR6OcK3fY46fTfNKCWfYPt1icXh79NbrB
vQrXXAQCMzc76ApJ76T5f6wqBg48LxAzTcEp/08HVMFcBi44xoSqaXT8GVfm
IObdV+4GU3hoUaUChpYEnDlbKuhemDNicilSlHwxHb5hM6gLEPsCBry/rKC9
3lovMkHXVApjyTwLC/5ymFwLUyHhJct2U2WB4kR01/TQ/DF02wyP0cX+Yx+5
YHepaNBVDuv8r9ndR/w0nSKVV0RCh3pphZsYPxxCkapf+Z6IQuu2O/r2wYGg
5P9HEHKvy4X0QVzWmna3tarWuMVlBGEEGi/QFH2Yw/xyoc6YRG1RXo5nXdzv
PnWwnhe0wM3AbUYHpIysW6LAiqiA6oV9wl1pIXrXaBRWSpft2rd8Q+F7jZDu
Yd7eVlRSxJNfIMwkhypxbev1nNGt+Pc7A12HEAOh6/NGNpwBKiwsr4pftnQK
TMQo8pnVpvl9SDMn1u4vdyNnc+5AlWpOOAWKk9mVt8W14jIzD/eSAoQ88wBe
HeVp2ron7djc8fxHQ3A0kxPpg2tZyeFdjH2YHHeeh+hecC39tKWk1kXiG4XV
9Dr4vhpSyCmTdaOiZ+B8QhbvqaxmY+NwXRLL5dIktY4Swp7f2noRFzO2pa7Q
1Y1UGrR/umPfpA7DUuRZe7Gb+HkfFNkPla084WRB9PM8WMmhI+t6ZfbNNs2t
GvrxMlkjIQ7k1ZypgnKFpXcKa8zvTn1VWHprB6v5zoZoZwlXNK/gWGZhfMMQ
Pk/DICWNB0KGz5BGpONMlLGvrVmWPLJBynFUSgm3e1QZ9f3YEx2wCRFAIoV5
UTYMk132E9uKB8o3lzHrTEMJ9IaAFSu6T0nRD8Hm9YlnlDp58KgR0d26zFqY
tc//dsFpWsmvAWk/iS4LQDwxst5dRIbZbtAw+TS8ZBldQhD4Dy+4LsxfgcWN
xztHfbvA8H0vke5u4Ei8e8mklqGruruavQIDmjsvS4vv9n88H24Gp6csVsPq
H+e4dzUTKrMyc76bd5YmrWkJO1O+7EZY+e0zUf2Jew04RgONfoAL8CA3Gxs9
SWQGC1qrBEeZsoq+ea0RvF0PeeUU+5eTVqX7vyRZfJ2T2SQvV82gZ+R7+oc2
ixfnPxDQeni0bIlan53+wYtT3AbnW/U7hQMTVGfHD44Yd2TreCXuEB5Nbbtu
TEqiXrdf56T5DJ0rspvLfNGxFHorrkSww7hg1LjXw3X53IXl1qwkVTSCzlJr
n0CutsfWv1hIh9RHIdOqJfotJxbBi0rTl2PaFb6andhOl+7TxP8yfYlI7i/K
LRGB81KEK2z4hkzzzFe3PUVfgyF437bGlCH4+Tv1gqzWoT1649ThPLjO2W/d
JsmfBR+loLeOLIViKM469doCyZFrZVvypWF2Nj84MWJm+xOPVjn/ow6/J0QL
VhLvCIbDib8yU3x5cdtI3iGJXsc3yvBiFRKjBX+TLvJALVHHisqUpJR5yiK+
Di9ZNfqX4Qh/zxnglwE1Afsbli2XawyZtQN2p4RRjT8HCXyGjtUx0fN1FPoc
b/CEg8BMZl2uJKCkfua+Mml/eiIZ00FADThi/GceSaB68XCPHgSlTNHyEcSp
pqn6DunuVpqP53SXKYR+JzpLjE84XObd3NIky33frQxLC/aAafO+e6WpIriv
9MGNl3hf17R3JX13mtMrI8Shi044xyOgqvSvC9OfaczDYRZuIwKVlzmsdkek
Wlib4JXmU7cWOjOLs1ctbmhVJREUCjTGUC/Fn/7hYwYs1vy2FLm4y0ZmZwMu
2gn3Z8I4JIxLwOKJp5OM7zBm81T8FjS0UXR4IyRoaMnG9ebZNKr6E7OWIs9u
XO9J3q6JfYZAnFZmW+2c/9P5prw9HIr9i6bdF+3uaUJAK4B0xv+3aqp2na0X
frN2v5otqZCVHFs1eVxRIf5xjy+9ddKE0ECQGfvub7221VCoSkCmQ7T3peOu
Cyg/hd8RjcnLdDd3CTPYtDimbCMhao4zgSn0QEQqW6MrJElgdMyWNlXT3qeJ
k5WEc7GHJazpp+UDOiwm9e53KABQ6ipxArwAlh915tGOQtYQ4pDISJLDilK3
xKljm3snNuiBTi6n8uhP0SKRoawhR206uGAZw/vaei+s40LtyBOMgpSlvKji
A1VCtWrzcZa/F2MYr7jsHfBCDSeWEOTywdl2EAAAHyQAFU9qG5bI+OvvGBdS
eOwdO6TzvckxlVow1LzZ6cnIVGi9lsHNJre8BIoifdW8yc+sFP8o4ebS9vVn
8szDskEL1xP4ol8wHPyh8WJX32f4Hh0rB/+iccOqpaUTB7U9G41SI2XHwvVo
sK2uh2q1UAZCgWKLI1N2oGT9zBcMZrO2mwfqnstVIOeBA4cx8A5SkhXG7bWd
1mCRgHh0N3xk+le4of63ZB7ksulFaSt/I0jfsfxac3HqGayKDTU4SLUkVe59
drr7oxtpiO4wPUIP2tJyiL5d4eCEoe567Hx+qwpLbimuMwVcHk95A5mz6TjD
H9GMOlWY/lEDZOJvsKnJY2aHY9rW9imLsleydVdKKCkjSCc1C1+CHJKVzkn5
bS8GUasoePmxUfy4nhVkuSWUOFFQDfxb4IbhCJcjyXN7OGpmux9h1FuOnX09
Hd1vnKwx93RKOjDK02BBZKvznSpycsKnRB+u5IOSYZ/NbDvufPl48HM0LI9V
JMPYjnFarbb37k8sPw7wltLT2ale+XKqKvXZhOXZ6JNIdsbb7ymSj+Dd7OUp
hGCSV8g9x0jr/nTiKsfis77W6YUXx9O4dKcMKDdlulkE5uaIXWIXznQav63/
5onRIA3cUoE4Tr2QYKhCVc/wPKN+FT7kftACwwKowS1NedsCSXUO5xNWeb2o
hj4mOiIOH1O45aqRh9Mlsz2rlajfh4YprS0VF7+6Xkm73wvYbXoKb6ZZMbLO
3fZKULeStuajhGmvGO+CNQC/NLamoMjVd7AmQ/SM09ED65shiwmVZ0dUwn4j
QmnGcqZm6puJ6/7JJqhl/s3MQ4saDy9mU2g6F2FVsWILhTtVzbRWcyLEt3Dh
YUSdeEG+VaJPM0R+SSxwSDyYp0z5iy4mxiJI+346YBtnWKkXsgFF+AKce3eq
FSp4ygLBFfg1kMUKf4GwgLNXMbjv2bOlkqMZJ4/14aonjAHjm0LkAZAz4jAP
SWz0MMJyTK+SKqF3xHqzGEw/KF/r/h75ZZtUnLkTzE2iO8ms+oKBmvYLbUVa
0egF3ZnZuLgCDUN7UWS0Kp4VT7cTy9r1xndXg6u376lZYIL6wNjXZuhsF+hd
UF4lyHLgcuw7vEmO2bFIdNTGSbRNtc2FN5wTAD4FCflBUocioiqsShyZ3EJp
rac4RPWPBTOG2KKU5GlF7sgLRhB6X1vkt75DwXXJHFYCQJ1Zj0n7yDi4Qkel
OISHfbVJUkv5tXbI1DFpOWzCq/uFnexOMzCFVdhi9xIsI2OWgP8MHIBwLyq/
+I5wm06J1KErcNf6IuesWMlHwlkLZCVYAO9gluUVbu8i+LwR/04Ms5lkkGjj
jnkA8AzHjh7kwtdjuvxv/VaDJl2FIdd74PWb99oKh0i0X00AFz0Cw5nAyo+X
ZcSavMYd4AZxqJk1t9JqBkBsvzemNyg7O1mkom3rUvmL2WrurNupWUqmaPLi
ZNoUMVPCTgl/q1uhPEZe01Ocjr/0c3dLTsVXRxYar28PkTgwtBsJbj0ABWb/
yZTo7U86D/e7U5jPFQrD9O+QChN7+HMm3xIedGQbENC7ovf9WhH0pzVvC23A
flZed36snEDAkFrqbnUyK3hXJ7y50NNxAQVVL9QIk1UzdVmiMHhlyhTVlHr9
IalXP+UdNt6PG/T0yVaUoKyOeHOCOo5gSA020biuQPeCxvAWFKX0s9UBMxYZ
brZUkcOk3r+zk1vVY1Ee4eapnpb+N9kvd0ZAAd4FPigYJYKZXzczr7x1sPBU
K5+8HjjMeEmzJm26LVyz8I9cXrlyeOsJ9jXzMg/V2gxKfxuowPqeExdpvq7G
CxNcYS2JJUX//3mZTUO00lFZiW7+IkkCnEiOKKGl5zkDOXU1raSKU55jpA/N
hRBMeY59r9MenDzUE5TmqectVlSPtPbyvUd9aPNPYorWMzzfErjoBRdXzoYv
KmcZ3zxG7MOTo65H5jZECNz5jj/aRE5yYXWKF8ZI+AAtF3+nQvGZOIVMyk6f
lWb9NdFcuX605uunugRM9gP3m17IeAWWHVNfHHSpz9u1m4UjFWwDynZa+id6
vdg5JH5ws+LBRlU5QRHc6OK5o5q2K//S4axdjqCdeMu8YX9ct1MTLtYXtaQv
8HPS+2EX5MMxWvU7RVIkcpWIHxqZpZJInf8Rp0QbyI8tDqPAXbGHL4NoHSDt
XGKr0q7HCSQc9DjdqtJcb0Ip1oNZLRjC2MD0mH12SMYcbyaM9Sh9blJAmN4z
p/o7i+m0VbRiQdQGJOJ0IudlEbIvE/1vqsXLOyQIepe7UthVpHBW23+rE/t8
h2zo/RanzsxsakS+EnfRPiQNESBjpy7xmYMbWLznlpAunBq6f4v9YU7TUlBN
rt0jD1Vq4wg5UBUBg+24lod6f2TcePodB7u0K6bx0mUSwQliXIbqzCQUWPlL
BJ55GRJTEFk59wHkCudxutA2qNY2Un33YywrkYvo8U6z+LsOuHim99eDYe7Z
ALiDPWMRYh6HbO0Dngwx4c/RYavtxDjdKGtzv8S8+FEZ5NBSR/hYY4tLM8c/
v3hevnkIDa4u9LCbqg2Qx1iHtz3+Wdmee2puXaH0EpUpyYDi6eHgq/EhZXwl
lH/LSSYbEiEdGhNQ4KXEdvY9+Zb1kEg8Z9PUeJyjEv5JrSxyEaPIgyfozK6V
FUnOfufI2dZ1cnxXcglTTwPfiIwxAY/kloZ6LPlQJ26VtSnKBQsW9kUTRq6/
jduP9/4XwY5Xi9O9nQr+N4qbpX6wPxAn0G9FbXGR9D67n9ZRk09Uls7LxXwL
Ql3R4aHBn0+2gy1mxy4h988ekR3e6tdK3UQ9nK45uWB1kJwR1ISRT3UC+ivs
9tsgWC+aulUzf/otwSQxgmqVZ2ar2uKuS/4U69+8wF8Bz7Polunlo0COdAZO
/4akwRgqXRowXmT/WkK36+9gAX8j/Cu3Xc9DZHPlqgMDSSjhnH6budAevqlg
+gJEuJzjL5eVWH9QlWD7AhvIZ8ufupVj93DgvMQ50gvIp8gJEx4rMN3HA3rB
wd4YAyFVQHqtW31gm6NC5xEWcpZJBX9f2SImRvDmLsA/+Ooh8SkFF9Wjgunp
N1GgimL1mysSRzNDR14Ko1NKUZxAO5YiVJPKH+Opk/rEaLJ8S49FtqXdFzOs
Ly4c9tYwcGcuGFdMePsAaU8N13uQcUR5PbJ5WJouISM8DFJtbT/KHMaW7LOk
XxL+8L6GLisEuqtRBSf/k055aG1Zo+wC6RiWh4xepxfBidXWxWXeZiBcHeem
YVpekZ3GqSeO9YuBdQ9AdXLq5dt5jl5uwU55P1OSAA7v6tBmD05ITYDuj3uv
L9xQqaMs0Taphb7SSMpHuUqjL48L4aU0ks3G3oXtTvfWpGLSgPKtIr5/nVGX
H5BeYsvDa7kZxkNEoKhPmRi3augPn15S1bVxd3yQmeDw3+AgFKDtgqvQrjdv
5EqImLJexweUF4CKpiT8H2uOfU6FnEY33gpEpTwCtVREh0D+zu46u+8fSYBK
DaR0N2rTOQyWmNNEIojrme95eDviIPy3w9TQRg6x7+ZwM72nrWMxteAKXSpz
OqYCHLZFq8Z8bDjhAtfq7fgypI5DxyLUobOVEKCEKWxhUBJUBQxWlvpsJEgz
yD+y4SjDjFmKxhBpIw/ZWXgr2jNiWGxh4Up9Abov9Re5f4De7/00Z+ocwHCS
0L75SoIj3FdvU8IwHtt2BwVUitKMBlakYalFkV19N3GMdE5LLRpYUpnSmDJ6
L8JZ+yCsXvLM9Unu6HDkECha7e5CUpVR5DuunW0acnGvZPTYy5v0uK1Q/SYp
+yUKmtM6q5syIBkcivzPvMv/nZI73GsNbOGWlH05L6ObHDSgUBVtyJbs6wMj
qJMX0W252WnVboNuL4zK2wQEL6aBE+qYTHCH3sabb3/2LxvEhhicwkL2co0h
RaUy5NJXWcAIAhOa+3U47UFJGWV+91xWm2kUheFJQDmcAFfvRDDPLMSnC8CS
bpVIRgIR3y6mMUBwkA7RoXIwXQ//+X0sK8KbmULTBlWiwzZDLX2BFoxxHdT2
HUP+h/Oi/Uzd3eR1Uc099tiV+tZws2NGpV1/E8y3NBRMuxgBzpFSEJIbULAd
UIIc/afPBjUhoGIBo65IzFg2RzYE0eEhO7+w+4URkwE+BBpQaO/KB/Hk2eK3
5bsSzhddfr5n4px6YPy1ghSRb6Jp5bnqm6/8GKgCc51FPCqoL9juM4UVxar+
CxecdPxd+vp5uwbAXpeczntWBVZAPEpACpyLvF4fDZppjJJITgCc8aNzjTsi
Fu1HtAKc8kZ4MbJ4ZROrdq9XMTcakOAKhp89NNBYwTJ09zcTvr1HscTLZQ3P
+uHVTwZFZOb+KTt7QhIS/njr7lSUDjGg53H71s83f9kItR7TFhWaScFQO4cS
hRY13BIqGk4RU28QDVfgVZfdICk9NXZIwHVZsBQKogPshBiH/teZiuTcYtiU
Gc8+031UIkO1gsY+529kV7zNiQyZCU0paEU9cyfF09RGd/H7InbfwPBMF6Fe
W85/2eaIIHIfA//Ik3fmPKIJWIENy7L4BHamWNHLq9sU8HS/91IB9Yk6Kj4v
yHYVx+PBr12Ul7IfaXvmAYFVplhUAsQis2hLTIUVtMmmWE6vGd17GFnJ2DXK
o7RkSX+TRbdvjQZVMBWHh9OfcVNJZYX8x8P9mZCcusDE9rGNH4BO8FSlk+EJ
iTvvwlOSiE8WnA6ZJ2zxfe0I5c1AwIqBi/ARND/UR5UpwA1JH0UQJ/67ZxRa
0XrnyQ2PVnJklVvw10JuBTKpu0RO5GbZYotlY7DMMiyQ7wJpBHVx8PsAgQin
gcm6olLk0CRD+jxMmGrzEGmx9DnwoSxz7EyKeKdeVHiC50sbte3SOqo+8HuJ
Z+udhgUfc1yjuqtMfok9Pgl7TQstUP6AqZns5w3hSlLCjoaGC7ZesR6i+pE+
iZ3UaNB4B75Q40VfutgpPhkOroTXB+UWdv0EwIKuQZSFsk8E2usKV/o+4yAE
X/ZENxg9ol3c8SqlMK5xx2B5kradEPaLSE0w+YajlaFfIAqPs8frmf/7dsxd
qnPvPKvDtsR14gwmTN0BuTEYibRPTqc54eC/YaqXbf9xIbqFSfF6KPT6bSSL
JamP9BBc+txU3AU3Nlb0N2jN10Oka07YCs6EQ3ilfKqC28zGrXKjiSxGGmjB
u8sCNTckZigkLkMsIm77qV5VD0iXxeKMq3eNWfOb+qCT/dkzkLSNxoGxGQG5
X5koj7W7e+HFBq509bUR3GiS6TloMyp56YGDh9WpO6b3qJFuuD62AHvzMb0P
WTMUK9+ZUZZdfL7SoEUDRUKekQY8q/VXU78a+DZ5w8qa3n9qlWQOIbxFb7+F
Kf+FVcecXEvW0lCzAcsasbCvtAmcMYBkWBZ0m2sCSJKlItLkXyPkzP/YTglA
zPu9SitKVI+ZRYENzZ09uOuIOUHMy52GURy976rYVdyscc/NbmwcwI8GzQh8
MVpo2lpjthHL8inDUY3OcF3leIm7WAIq60GSf6mlAKacekP6JpDtSceCfXqr
md4+DOXmljRSLTOJURRUsh84+Bar/5elgKpj+vPUI/E1hN+H3FAVSB7CCHVx
D10W8h9uiR1qq3yGSPGOz1O++PxKsoFbQYEwU/czTzArkdq3rb8+Nrx9clDL
wj9brFYRGizdHlKon0q7t+RiTfgrUnXJYdKXllD5qc/xN6dlvH/gOh4MTx45
c5HZzm6ZBjoBGUjof96xE7wHuJ4okAGvNUCdA1FDgNnZDyy99Rm/lsdzifR/
4RzWxBtcRzTYzuaCAcECxaVrAJoi5peKrhiy7h0+GqxdwXH+l8ctLzo8oW4/
E/Dru17PcT93HoAbuHUTUsT0WGRsTaNrBB2jktKS+nlr2DzVr4I1yAcIe81F
Zf7Ui36KiR6rbr4KtgaGOuA2NxtxAb6CsjR2Ed0Oy2QqL4xREjwsEMLHa+5/
VsoGpNnBSZWbZXgZVbqjfYZ2GlTRT9pKp0sOc5Q0GONqHS8bNQa3GI2CzPCB
Uqy2zBA4Gxooa3N+qfzPpedv7zYNRXw/W6m3r8tvbDHSfQUMHCLeD12GZWub
mdMiLwwW95R+la/KW/3AA7pDrZQ/2bks5gF2+iO86nPWCV1F8ank8USciRVM
oOsz4v5ho3UPRDK1/SHoXXdDeI9zsrsemLhf6o3VAxpQAwXo1dCOTGtxmJyS
zCxOoMlOP+x0ABv8LTcYQaeV+09VIs8fd8OYY4kjG/Uyfx34NPzTT0IY9VbA
fwuyEu19MSjYQLEfj2hLiqh9FA68UBwAgkNM+W83Azf6Rc9MfaFTQ1Hujxnj
1282fDlYNVFUOD+HMWLZWV9bXjus3tKey+lM1RxmcRdt5xIkEQzH3DnxY1K9
j6OLsVlQ90yJoVWs/uerw4X9sYa4rmvkAfQC28ernuaKil5rLu8kurOic7kn
Wo0bLil1jYkQknrP4bfm1ho6TNYNpbNwUXLsrQnSGGyi66XRS/BU66e6Cqq5
8ZmsDDYvuDJIcJD6GnHRNd8E6bqz59UXLAv5Xfv/woNz0VEvWCWIpnhOkUOJ
p20miL66GCkoo4TsKbIPwCzc2O1ndrGvL8NSgxD6RwUeSmwu79Mv6+K9gy6b
1lp4mzg2/8xOesIT8xiEmmCDBZtu+vbR/4bqRuZRkLkvOt4k+yVNV4VzbC7+
6S2cJLjg3ubIc5Wv7BuJ+JOUeO8aMvAjET5w5DEeN2wdr4+PopxJqsC53kon
7j9KC7ZwAVWw/4gQvayDMJBEP48MJS+fcm9BUiA/i+54NwF6DVMq78NIqQPm
CMhvCtf3p10CG3wTXR9KSUh06KSKaRxSMKKcFTTjrmxI0XtRIK+sk5fMXgT+
H7LMn/CzIxZBLhn9Vujcg58UcfZwZqhiSq5nT/ur7sgEXwpGccQ2n53agGwn
odNpHaJUD6rOjajsz7R1OXV1BfcEimG4uyyw395hLP7npOf+LcEv9j/W3SP/
46Cjm08wPIZNBewkmF+S4O0mOCfo8SacSBOe4M70GDqHo7TSSfpeKvMTBhzk
xB8DQy6IUFP+B+h6BIeQefNXS6zIB5cemy8SFuBNjNiDIhw7eoye3KFNLdcX
/OeNTF3Y2cIdaUBJYv1r4zWsbZ5LsnV9OvEmW2ofHAd+4D6SQh8qW/GfQrjt
jpXS0oTHWSh4nRQnEu6xkyLsrwhQyE/X9MdK6RwwNj4LSvEsUMFgvSv53Bax
4qHIWnQ3GAxywHGzmbNSATB/ebL1+UxhHg5FfX+hOmY9eW9/Pk7RE3eKxgGW
FF5nt9hfYOwp2W0uqr4itKvsU3Q0krMS8k+vBFaOYSvH/qz72DklS7TYySUb
X1v2BTLooGUWr90R8SG8YkAw0LaT/lnztfTDaCjXw5cQoVp2cJon3flCzd/M
DkfzOlPu4MweoSqQkIAdIC+NDtKCddRlQhWp6U+lPLTU7SAwR51fzjbmcWq6
yujUF1aqvkElv8js414aHOoQ9SzRErHAMJAGVOfLWadywB2Gp1tGjybOUXAT
olwRqbAUvxCTETntdBEiA9E/+fXpwSZrr6D5/Ctm1RKyZHt7Pk2sKPqP0dOM
TtYDGtg1SQGIqmyLmGOXLn0hAfunHqwSjAdGGtG37Pk79x/bT28MI9JUbl5M
gwhoxsJ8+4x0qblHtXMSwTYrU5VrrU7Uh36Qpb2X2Vr1r3izc2pLWLW0Jeqy
tlWlQ6SmLpAFuVSkeovPOAQVQB77TnQbq0LWib2+L7PUvJfylIpp84uszm/t
2wZT/Ab4Ey0cM2VLhbV8LO7u/AEhoXcrU0eWQgRvydfCRi7vKHL5sryGWSqk
0Hssn2Xwm0Ae+PiMz4terRscMN+CAPVoVbgem1XpGCbcOPXepBRKAdU8NTPA
1KZMcjwDc4TF2Y3gej0p/SGn5M9gwLfAUPyN0jr10/0my9MdL7qU6NHK0Ph6
8qVAja4a/JMpwcPpSHGYSzTFNTPSUBNDHUtu4zaU00DCc72ALs3OMn67QEbJ
VSMSVH7Zo1XoezZvHeuL0J/+n0GnDQYP4tS10Zdkto+USRYg1d6/5qTsW8kA
B3GasXErjoC576aLKdFBwMFGc/KAefOE8HCtbRN6wkzxbzC4FzINNQVfAFjG
lXpZsGYoGpO5gXPU+UB9pIkDbxFXvcT+QPldZAyggN2BjLh0esKfGrJDezhk
rQ7Q8m9wjoGDaA+s0/a4NlLHuLnKD8h0tePsMBAnVoRvfTowtZ7WaqT09QZw
8CYj2v98F/S+BQB48vIq3rDKmYOcfuV6zMCNCbReuODvUAhJeOofXpZ/pC5b
oAQogH6aHtRAll9Bh2Fj0dFHKXivM1cj08AYTnAVk0YueZN3MRiHYanwFqWY
d1XVG3CUepWvS8h1H8A9Xf0UPIBHemFi03tH0iXQoCveII/l5t8ArQi6dhgJ
whXELienyZueEXf8cT0Q5wZLJtJWwYO6VSYf9UKaRLCEwxzBQO4FiLpC2/A6
OHq5yPKfyME7YOf90+t+SXyCNxiJYJNR65qLJ4nIVl3WpgIIoVUtx3e6kOX+
UajXyHg0YNYoxRl2vFTOt7ZF2VM1DsDNq4P4cA9Dm08zc/Ra7+Tzeh+bJ1Yf
UMNsrlM+/sQ2PslHF+Yj3a12PmKMu53jar7irCJyxSEsfkVoRQkDDGfvSflc
p6hic+RUIuzj6/Ql8EBG7+HcCRO6kRFWilV3hCq0ZP789IwbAIWa853msSzN
Ylv5EYoglaDfCMyY4JAv2QpWlthOe/zo8/yRu9+OfQWqg2GgY31XW0sQg4YW
HDAIKRHNc4M2t/ERNDwCmjFPSSHKd5sIjDgTmaPYHhmScQv4PyP3pUW7BbfB
22QVrvawDKdIgT+J3KvBP2t+WBCzzI1v0fsRTlm+evSVl2W2WNGvk864jXFn
ttirpRm0coRrOPn7wSygKV0dt02+Vt4Hfsfu+8QbWktMssV6EIA3fqxYvdKc
hrwL38DyQGKwePKXU8uiCO3z8r7w6oAGAwvCq5y0w3mLZTSHqiRUvL1bVe2B
NuxTDBEzjpC/Wq5tD4OyjjfQeudNGNe9InmjqrdYzOHtgEhiR2MWzWQPZ4r+
FCK5BHhVHXpw5OufdOvIDVa/KzIwVxc85WazbByPYQkiLPYZcUjSyDJ6PPhi
4V2et1+hxBJAKNXtwmSPBYB0dxFdOADZguQceVNzarB7Jz3Pcnu8zvGHjqgo
1royHeBQMNy4COhUeWlqtHb6B7YrHDXjB70wOopsIywYypGgxVGiraquzrj0
iVoIAsZmTYAXUEplRW1ZmsLJG/9CZJGhvDSf63p63AVAjrwfOaJm3FQT9My0
Ew/NzVepB9xFc4s/y0HbzDu479EMaPYUbwS/tYGweEh8k/76+tbgFnxCxnLg
A0BqBsAk/Fd27h8wKhDeC/Zjjat1DxGOtfVpncNvxJ/f+lxCqoiwMG/dTHR6
pSaptZOqkSPErEytF56UYOT+aSToeS8auxDxzJWQvWvhGqF2seaLSTRBDHo0
Phuv96isXrx+hN4Mj56Oj7VFgIVr9i5pc7yKqDZqWe4u9oK+J+SZTrcGh3a1
t2k2TgbuiU3w7u8XtYJrf2imd8jRrHLLrcIrGyLhCif115wdXA5MZAycU//F
xw21JmWPBxbYqMo9/XKsRJBvjFRuGGl4zqqzMiCnCCoMF6kvRe2EMHYnoQbS
jBqJibRkjomxItrloSTEuYp9J29j9UY5BDLD6tFFKtRpbn3lDz9NPSjgmzNe
747oQ51wHADtAJQJUCuwq22pwMH+iW78zLwnMh6eV9TpbM1rDpwLjnEIJR3k
Z1X/wrgUUSgGfm1tmXtEIAKe9H1t+FGi+TF0QU/AOiFbgD3djZ43oM0RM5fW
Okjwo5gN/wxeEXfenkHDpyRMwX2Il/289DGlpJ8V7tHvfFEt87bsAqewRDYT
zdTlZ3V3nT2upH0iASgl88vorkGYY9N6xNcYpZlSAXDxrxznPBC3ryq3zDG4
L8JLP+LKGrjmpP0mqoY/YopcKoF1jIaeyg2qAUlVUKHM7PZM8vCx6RbHGawf
LIrNQkbUd6uC71vhpKPmxxae5vZJq6jd2KIHhAwtI1edSv9TxvjeCHAylWep
rm2VUb2ImYR2Wza4loa1iurlwK3im84wpFC74YCFLwfSnrtDZ3aAo5mERkED
1SqXjYgsQ0RcXaBUKqy9UZTlflYUE6Hfle/llTAqiM7+RSke1aLyQXNegnkn
ZqaLDKMzOoHeOt3/dHdB6Y7N6bHmr620Nwe4KntP7nvC7qQrL8M6EH1JatS8
LV9tbANAHyXhwQv3mou3Ebvub75C4xjua+AA1zo3rGevGoqad09emA4cUGQ9
JomjONnDPJ1gkQXE9tziXy/77pLSd6amslJElAzPnFtagWe05BwmxOYjWZ6T
P3SCsU8Y9zRUKLrIXfEAGhvehtcNvsu1P/89xRNFXz7ykqimyzhyrdSwiAuB
1skWAZVMynY0pErLJlsudnPiUYGUs8I9KVmMt3lWSpCV/RCBpYSzXlrIv3Le
E1OBhg5vY4A50dzrm1EHhk4cHdjrLI2Iq3Jp7q3l4nTWSlL2Ho6jDacU5dUn
c64zf28eaAU2yiQfmXZmiXKdNPDxlXUE9Uj6hr8Ke/MuslSYAl3yGtEKA9cA
Vt5e8jnSRtNGRMkSmg3SfbA4CUMK7cK1jVCkA5WgaYIqbLaT8iCVF2G+GxC6
QgobAt1iFq4kyJ4i7uqvDQu58UAcQCv36UByeBOf2Vo544WO/MNBG8xlpY7t
0ufIiTSoFIjshTFTe7lXglr2RtNkBj81Z286Dnw+aDj1hYsgjEG/ks0qbY3z
4Jr8VriQ/1knJN+qcBCwqFDvYf+Zfmo33ZP/rhMwMt0ZFz5ZEbh0A2UPWyeR
IRPEDk4OMhwPAd4QAjVZM2SsiUMc2uHv03e6VoX3fTrJWVnYWMNI+SCYq7Q0
H39kOMvD26Y7vQ2dZvNprcs8JhN8t2fTIglc8e0wrhESbS3+JiX5DSyytDzS
96KyWmgSp9cbXgqZylxyYw4uML2JTKlP4T9m15pBdtMQEMPMqbIZCQ7tPXLI
0EQnT5YNUhVprj9qiivUZ1b1r5ktZntaV+ZANCxV1FH4QSMjHJcUUawVgaFD
GaWa3VHZSxCvgq6F26QxwrVjF79E3F7c5kvIAgOPOZ7dyyJRfAZIjI0PLk/f
cYj3qi/itLNR0EruWSjFVqbOePRiqVdZK8nL6n6eXL7vRG7zGSXIbmdadI65
frvEYEeQ8ps4ICVsSHaJ6cyBrM84V+QGkbzs3xokAI8322oHDTf+33zS4yQG
WBdfXLamX07FqPWCk8s52cS58dJU4b+O5J8XufqyyG3x65+R04XrA8hzSieD
baxRmttE5+SJBdboLpvTHCG8/EWCJylwYf/ep6e9MBsPNjw42cNKUB2mUvWp
PkpEnpz+j3+ENxQZ2A0E/e1nl2QxZF9EsG3diGtvLhfuELTg7U29Ks2pyRct
P0hpEpaGrIrTUE4fIEhGA6mkd7O+Xq4tzBtrA9jeMTF5w3NiCeMla6WRQlhW
G5GKfhV9Vuv2rTLOjebVgjVf0PE9kraU51JYGIExFMrwJ1qp4wEy2mbHbyCb
YGm/nfTIn2bPCzORnXFU0aXFuYHJjxpakvqDsbGt/jiu4L4w2D33B8QDXJR9
1R1kZXXIS1B2j4p5CvAQ9nXMJLMbCv6iv89UMCsbwDogqO1QoGh/HSMgX3VP
Kih3tmwT5Cm5uVFfL4Tj4AydsqELtrxb3GKux2WHMy5+9Wxoclf0JbasR9wR
sbdysiEI+kBr4AHfbs89I7XkPIB1he69ZCljbNyVzRZTQKzze5b/Y5UJcMae
F1ndZbtFlLjb9h53M7a4w12/kfp5SBOmtPXwRU/pQWo/y94fS9p8WHSdeFQE
9cpF8xQOXFdBj1MtYx/98Rohj7DFOh/eEKSltGg3SE/fGZo+ewxB++g9YlcS
R8ztkEcF0hQWWABLDv9dTo6oBEipnf085LnqZi4wKP01IWw6SGIWnmITb9TK
ml+uaJqE/vdRGblzxRXarxwGBKASXIvAg1iKo1OUKD1mT2R015Xe8/z26Hc0
VmE1Va0moE63dgxdoyBlo+7B3ukE2LRvpQ35UpwfSEjkmaFXphCsdZLa6MPG
qRqG7JFxUTWA+Xz+oKUBtQadp9yrlV/7UIeBLUZR2czLoF8ybxRmv3ZTqj92
U/l5/gz9BpU15FnetH3G3ZnvyS3cWbWl/W/Pnl2a0jGWfNxnHu/U6VlBLupX
FMoKcmBu9z9aWCsfUYf0dtgVMH1U+q2oBlnpG/mEsBOrxa8tOTbq3t49atJK
e2ic2+syDyZOw0Kk8XL7AH2nvfPiRM+eV3v3H4Z99KDLw/YnHu2btl0iB6Ee
vmryFyxN+pEYx24GRRHI5syBu8Nrf5EZ5PiWzRyoLyAyLUwnB0Q6K8/8en6P
KKYQUq2QItAFzzM2AKF15G1ZI1wDRKSwZkbFjXZhiqM5mKzEPo+nYmpf0ezc
n20lepcme+nvLSpGZ7WXogklZbdLVj2fLFAkXXZWdoXxz0Y7qhU6KxbeXacr
c99BqKM5iCzoJDXl/e6Uy5emXeFJ5irMiH+WCkeqS/R8wraQf8a+f5HZqZN6
e/YBJLKJeGBgIXtec17D9WqTtxBZAyd99lFh4xET4G9ev2KS9rQ4suLiu125
lrnKbl0mapUS0yiyQNWpw2ys4iedviZL8xgYCzy8UBHHQwEqTTK5uFCwgQKI
bkdsLseNkZnv6Vo1MHfp1tt7KQ10JiwXv7d/ezSK0UctnvwXKeMp9sYGz6+w
Jk5DHfw4OKwWqqISqm4H64wAJTmlm4B2q6jyWFpMtomldOgodJePr8hpaXib
NSRZXNrMVltffUiz3soC/cmLrUcFa/W/0Ooo/nwl7hYEyxRGzTOLTkd9VK2V
vu7f1SAgQjY2rTLqyMhoEbLlVL1xFLMRBF8IGWJxfcMM0dXsUnACTXtbCXr9
D3N5XHl+ndt5e12Jl4+kxI2fxPQ60VlvWpdM2XplhrFq9Vplt0hDD0/KmoxT
kGmyJsEmGlRrUD+MDNfnyNgpjA7JONw8zqov/C8qvZGRKc0yffsldVi/xnAS
vrFXJV1UQcjm10O1r0B29kjUrXcsDhEVP0ZWCPQkvx5Kd119lzUXnG6Xsxyg
cGoptpoTjSdxSvzc3xlMgM5EmMyQpHRAkRl/anm38gdH2xGwYMAN+at7kocp
MpCvlV9SmXz98ioITpo+3W2MHIRXWpFvR15EDSgVWfIeIpESd20++JXpuGHl
trN8WSLzzVnyTy9XU1SLPmaygTq4SgO5suM1ySi2SL8ll03p4tOvyT81sG/T
eztJKIe+VLhEDQDpg/w5WGzLp9P1L4e+AoXO7sHAR5wwDHZq8BcmbzsAaAV0
QJe2/Sfo7ngANpu9ou6UnKvvCydtOW/SFOEMrGcQFhQQ2EMEpbP0aSiH0vHR
/rQnbsPqsS0JZJhIgStaiMQg5SbdwTnQLARKWdMeVjkRgCvWALWO2SGD6+WV
stOs696vakD75m+6+rAH/zVgUE7+LGzYK965kqG4XI+FcGL/9/aI12C2PeLV
RiEwmMjXb/aUcSMqI0NHxTKtuTIa+X9XK1Cc5U4CiuXlyZfBIHJNGyVQeQEa
CbpT9TEOvhV6QMpB9v/FCidmaposU2cijwjrwxIZ9oOTK/noH+7GG24+sT1I
lajMC9CJUz0yQ7Qua9eLQmc9Dhj1PX5zhFgA19T+axoqVMm72HufaBd/3MuG
O+ykRUQT0yyGPcRDLyLIW/YnRJp6L9U4z4GGeeS7zRz/ytfmbmEXZV4tl1rz
r5E9KI3cp3HxwKALOJcdpcYMaJVK0ZlwyPIqP96+1jFDN/ss0kLj7bYHW4hg
MXWO0gH5bBEzBuSVRZRpgiyrMuoXvf+wee2P8LzlX7UXMjkAZkYSBIf5QFHz
1PoFdZDrz74dIR1hOhKrUhdYpYnZ/7ryuGxZPwCjgBnMy5xU2+Ks1X66zb2p
sHoXfGTdtc+kRZVjsCnHyyNrwF6a8aoVK2IDOZiM4svYfhI2v2adi068q9if
KtcTpqP98Dq43hYzds87OV0oHpv2hNWvBsnVaikKQByGmH7SHarrtpJKjDvh
9EuIyi/LqrQzSIruPphOx6IMAbPw59JHiZ0Hv66+25lWBlxY0xzlKU0FWt0l
v5tpO7CUjRwqXJEjkgOJsOREhvcOX7KxE/musuo+BpKrztU2l1CSBZ/r9rGE
kFGv5c1JIFih918QwlNE+Huxa8g74Fi+HgvXEiezmk6W6yg9qjw6XTXMjLJd
KiMV4qY0jaUJwQHLKa/QplyQokZL39PuEEmtSIsXD/c55J4gzDdVgJA+XWjV
pi0G7ZHjFGfOeJ14FSthu+ICfC8e189RA16HzIU+JTncLv8Q7VtcRVuhLcTZ
fWhA+12PN4Qtk0QwknXKnm/ZXGd5rvviNrhlzvNJTGMfW1OAhUEKDbFJMed9
OZSyvxs1U1yL+C9WXb5ZqU6JfjQBYYNuknO0+ifOP5fQkrOhii92ycFpnMaZ
wSoO2huubKMSS5x2R8WDtRgS22DTZrr8IJqHKF0K9ZcGbFWdwInHnGbalU6o
i7AvwqUkHwfNKk7+JF03j1S88NgOqYw5bjvBG5u9d22ZqMaHaRTxMSuSEJ/i
ckNjGpOfIqe9HmjKLDgmH0UKbNVdS0NoifwaDJnknT7XxOES4/VOqooTyRNa
yJJSSm5ik/djAshb/doP9SCB0T6n37Jovt0Vu3TBz2mNf4loH+nZDdmr8LaF
FN+qkByAqNmN2mmgqL/0lsvQ/9I2QveeU4ADGxbrUUEo0f7wY2DW7zoq5Ivr
hU99/Wiywxtj98VqVTaHpZJawYHC1mpeo8ieJ/H3qWc0EedlT+Zr4V4y5p+m
u1arRRDqzC8R34KWWxhQNqaXnM1tN12mkc789TbEQjHKISjV2ENUHcrinxnq
i2l7b81C6ABh78r0eYtXcawIG/WX4psYz5GheMsaSqRWKNx9J/YKZbypiy1Z
mgaAuBoXbqXdy5hClYdOmupqu52pGMsI57//sL2i0kxxzbcKpVxbdspSeVr3
XuKgNV7FbrsmWZxXZjIC8cbqm0HCXsuFQKYL/kz8XsX6d8MkdFSdElx6cuDW
2ZsTHGw3ZkriC/upwK6uoK45t8n0lJS9jOZlLUWAvoquN4toHU50zaN5W0J0
Sv9COLexu8eHbiFZ5uw6QEcas5Jfmt/epBACsbXDpPMI9GjqV2985ZGkae4c
/k6URavTbVv15O6186uw1xqn73pOgTxx5Zeck2nHMh4s4HyLlBY1YxuFbfB+
qHFHhsCKePX4+HFQcoOwIk0QGHVz4SbqKpKTFua2j4qcxkjNqvZp0Rb17AjD
+VS+XKOI64OLIJxxlFnETQQHSUcwkEHHwwJ1uIA0OgOR/9nZO6eqivaUjX0n
FxT7GTruLEOaRQ8F431pyiqA0uclpcoIgA094Dy63r+kSXgSXbOUqHtQB8sN
BQxvtarkXVFx3yu0EQSlnGKHPAJtRXoM7XezvLKXOl98GJa+HhtGvJkm29Po
b+F3/dAUw+2fh3IzK67L69pHoetnHIZL0B0SIr51fJDuQDKMYJszNlJ12XyS
iwto7OIvhoOPMmu8A/NjKYFI/OxNtE9RAD2ekXsLSZKCW7UcUY+K54mvP0hu
P9T09fB/saLTIl60/yf/grd8mKpHf21PhjI2UMrp6Qb4gWYdQ+Mb36ZMP8Ve
Sa48dsYQ1Lm84O1QnesRoj57khJIkB/UcEwoiet2ReUhdHRtjpiJxIUrQCIN
xhRK292v1VyVYDAC2IF2KiDEZjGi3kf6Cf2HVEXhRTP0LNzPe1OMQRHdZTmR
N8XR0zS/JQBpGT6sUEAFsqbF9ZhTthnwgFXUu8Y9Lf5QUGniv9Qqf/iPpGpi
XLG1GsKiUS24qy+JdRUZe/eXnLBYV7Sy3xjh2L2MgNHPCbSvjjO7h/ucZoAi
rhyfZ/yvjuLwQr2X0mjadePQuwbB9Oj7o9qv4EpfcIQshhU0nV14tebe16Df
EiqS/IjjFAyd9o+Xx7bJ1upqQa6jVF9DvUtrbrvkoPP2xeBkBDH/yb9dNjaX
aJ8vtL6uWdiQyTmr5nxaO4kMnT3cSA607wHJBYyI5vfWp5hteNJ2LM/Ex3bk
ePtByIUDiUA3ijaNF+UbHjZHXtabtN7iDmPrVbn0IP1HTs/agn0r3nRnYK6/
yZdEWoqSCrI4GqUr7yXDX05kDrbr8ucyGIq5jfAA/TEfJqti44qoAuqQ8Lry
GHDqvWzOgCcuPgUXVYJYwxQilufEPkF04e3OTOcspXOaS7rDawOGjUl1hw8Y
i4x9qwtO4FPedTc3C6COSNDRRIiYzqhNTitZs1JMzfzn/A7P8vpfrf/uIUmY
dbvXUD19PTIGfaXjeAyDO9J35ebHRUD+JqhqhUpz0+98mwc2bzHYlmmT0FN0
EX6xNc0bOqQHUhYLRa7V7yhUHweXE1m7TN/0gqGgKep95U3MmfAQyPSnXNAF
o4SoSQSojZzW0h4jiRiX0BOl89rjwttpfeibBU7fsTF5SX5ENxCvx2NxWK9l
06F7YhWhdKS8XL4yIoKX34K8d5PZGi/ML2u3K96idL1VI4BFnAe/nfAhI5zJ
0/oEyGvm0rOGMYm+xjY56bVMVHmlUf0BxUzVmhyylO7y5poetg5qn96RI3/o
DOLXmdd3fkkKTdAEMCZectwfszGKjKQJRure7QH3uJYQZE3CDFVKz9hngcDO
L8d+cAn/PLDzmHJPaaNqy/mmec5mIPQLP5tAf5HA4somPOo2vJPQ6Nr5qDfa
cksZ5Nbh2ijw/aPkGj8KToqKnx73L5yt0OKbzhoxhpA0i4M0xDW4I/rC0+Db
1NkD9ihnSqF0XgmVsAdbJ5LQ3eBaGPr/Pjde1mEQZSdTYm1OJMmsSwiPM+nP
R6lde5Ga6LtPn2cx7Rmr8XU+va/N+nKJQxPROoiJtRvxhanhGadPin6SvJFc
wYKzKS5J0OpMTxeVeCoZ673rvybdG+SvdaaVTrG7wnNAqNFhX9ez1qdWhW5w
LW8oZXixAVmKnSClnbg8qLvQHCUotiBHigkAMtLPchQ2oTAicGvG5a0SVk/o
7jWm2+jrMlcM/FZl11HdMu/Z+O9M095VJzF61SFWMom9qhn+HanyRKlR24xI
wu3iJqwIjLBhKM0B6jKZ9fV3KIInICOPTISKjacyPaVejLAnPRNkjtq7tpoO
Y7tJogj6wt0LVVTN4x2fOcnSkJrxihihyy6cQ0yb/mJa12+JsmxHEkqWC0pN
j8LsirZG6Z6xKz8agODqj681WIXBSGDLnXL3b88V3cGco+yH0Sojyo5cHN4Y
gpZ+hmGE/PPo4h8YyS66S8ViFHEMLlWnqYem0p7axAUZrXYrVHmR5KGpuAcm
6cZl4gqxcAcMCA7jjaH4dpHN6SjdtsLanXIcejmairCy3Fih0fBWcun8yVN5
urDKR6/uCupHbOYPepzI0DxDm0gJ6JUIaH8LQybQhQWIHv85p/Rt4NT/soYS
G9S9Y5hqGDr0Vic/fbClUBqt6UWySVH8w0sTv1MoIoLOB3jcjA6UlRVdsHj7
AbQogr1vmkyjRXXbHn0h8ncmUJN55i0m3AyCgXgOO0IbwmHpDrujGRIMfmE+
OizNYf0PStrZFmWCLr48sM7jYwHf3KBcQsdYxZ7BInQbajsIetryX+xJpby1
VB98zyQGwLvE+KW/9CclxM1lLKl3LhgVqvLZzbaRNsPAlMUU+KxibRlDPbQx
pTqdWe7nJgRwTBNqFamtWj+oPzr6mGolbt8kNBsVdYIAYlapxIXZsnWBqwS7
v4F2B5ifLo8Sh4da+Js7RW3C68sBMOP0DGR+IvlRSS6mkrDiS2S3i9OH8iW0
GexIhWnUkrctxv7ukUNfNR6iioiOlFbYShDA6pH3/RT3CHKApXZeGWKQ8DMe
ceqhNb6qt4YeXVFRCE28LGJom4oDMbJyROg3XHl33tXQEEfXziZyxZsaVyYi
6nkJBkZUF5kgoYS78vRgsyAwBQVEE0bIKXGxT6+T8L8qJUR9lpSo4W6d8g0M
OdfcOqF4TlK2NjdBZJrdfFhTqP9zVKasMRdZKm+i8YR9EjZ3g9wjQdrnzoA3
L0Ge28mL8Zt0f7CUz/OtzEIKcNZcuUAV1RpKk7Qt64aUU7ACBh4FkBaQYKua
/QPOGfkfhcNtcWPBgg3ot8J3OWctXdq4vc5xYuNPqRAbknprOSZWfSawQO2A
XnP/r1pmArumYQhwEvM8VHFvlmWaSvdNTKDSm2eC/4AGl5+FO3sxKWxUi1pZ
do8xTd89HXjV+opUXrOCBwD5Jlncy/Z+GJh9flaZgWTKpEieKzXGo7hSbnyw
z5NHdGIZX+0nPGOFpZJRqUAOhRGcN4VJDiJM5h8MGhPQKEv2Ph+BofE6c5DA
UwoDOacquenOYKQBwJTCj+XD99KtStobaubtrz7T/VXxsBZgY6pGTNPv8aPO
WWvKgnhfKFzhWQMR+uO4G63gyKH22MeWWZMmubVsGpx2IzSjiB/JAlnZiK4z
euM4mTfaXfG8mT9vlCbGKYSytqiS5ED4/AFRSAOtP5SVZZIwDpVqKvCDH0IX
cJOmLYrLxCju760YoGQHNFBnoC2GXYFbvzF2eSxoxhtdSXmvibDUayBNvExD
BX2CQzu8o/Qpkjcv5jToTEgQ/UFFeYnnNIv1PLYzZtTMEJB5J0INs7z637OP
IcSn0PX2VMvHLNTKq48QlLIyzIc4tf1YwyiApsihfmGevC2+jIlD5d35aDvX
XR88J3lymR9fyFSXFkVq2SSO+E/Wt4qgQiZiMXSSFIsTNW3UeF4BKvQ2mNVl
VGluqVJlbTt3Mf8/dTGGIfva1nNLdhAQS0YNEf5dWVFmyhapIjg6g3bfcWXQ
9R5sHPH37LBNrzkQayullXAj+pjnAV6qR+zdgyE/Iaj1pWyG8o5kfC3FU/ax
k2CVxgQBGL9HlVqbPsm+Npl4l37mxMNOOXHgrAPS+ZRfmV3FBYn0T7sv2zZn
+XqGdg+KLL9I56+saUbclpAF9xLErp6W2lo8c5jTbTSJNNImdHldKIfcftSW
zxshUufpKKGJXw+3tk3f5MchEbJVtDsQYUYzJfbrf0FXcJgh8UC2TO4AUVML
QONCbofebwjgpbug9Eu42gCGUqyRt8+XJz0mRghUpEdWNoN4/OP/TGIWfXip
dSEMocxXN/QunhN01mvtIAUEY22WKdE1XHyqrkF9ZCnNnGPB8EllqMd2yzYG
Ld5SJpw087rYfNBj3JWIiyBGIsOuNkqH3cbAUYQwaz4bUWVFMigA1Ck8BLyN
lv2EDHmS40Z+LWhWh+OZ6pG0jJyhjx4hzC7CFP+4rwCE3Fg9zMDW4NLL2nfO
mTq/myW3oMHI80ZNOpKy8GpXA8ISEI/9XuvoZ+q3N90vKz6Dq7TsIUuOy7Y0
DGFWE9dPZXG4hJVye91NHXmltRQWc4Wo54VvDJp8vSgHgVGtDiF8Ii+erdF3
+1MKl6anCbNpxc4MeQa41S0qe+zFQn/+N2lzYmVql9sJ3f1goWKnh233Q+uo
egkhzU/6nxlDT78A7Y38zHITp/8DqCc8m2yBjW5s78EWYgasB1vwu19XXaor
MgqrGgVeLfq2/y0BxOWALU5sx/dsklVtZ5yyKGbgjuxm7IIpscnje3eoYVdz
5wqRDlXQIHfU4vxS5CT51DOUupNae9FU9BKvCO7I/pe6k6ec2kCbEyjMD+bi
8IsUcUVVNKGc2lVyCO8kroOGfLoJX0ElchBBejen6kF0Cw4+EtTZuS4Of6pa
8XjOx5f/iFW7ZJVbvAhtG9/qvDquZWxa2pFV4YI9lCSzxt2X3Ihs+Ll+ykF9
9OK6x39FTPvkMxA7xqtOuZx6O21xvn9H7smT2hRiv05kDYrMLmbqkaVf7aO5
y7ExX5L4aQ8XChTDSn5jlye6/JO7JpyuuTSt0Pv59wM+t/7omLZzm0wtW+by
Y+Nz9IkkMrfdeTAgl9J+SjlD//urFzS8yhSubm07Rbmwx8Fb3SX3Ki5h1unG
6bztpWnCGUelvItpV+4P6h5kp/akx99QShHHZhMrvItgm/nO1nWHcyJgALS8
h6t3D/7f2BJkgC7EtGCQGbjblddCXrfm1dB7/SQE0BR1ztqXZ2Zx2EROJfrJ
VyTZz5FnwgXJvaRQrGJw16wi1q1EMk/8pjxjGOc94ReEbES1ugBiE/woJ9E+
ewK1L/nfklfjvfZB5vtwEF7LY+vqajkvXyEFiQRttCAuZ1dVIrdqtZvAHJb+
Vyc+HTWaZIfi9w4LJTKtO2UM9S8qTqGcru83sitLOjUr3GOFBsIk5kr1/aC3
fS9wU6THJhZZ7dxxy3iybG1nPACkngTocQ0MSh2mO4Edfr06in6qenXZIwz1
2HXiUVVA+6mfNcNlx5k4ZiOnW9voi9z37ugvejdJ5/SLi8Wn7xgcptNXPc29
J2wxb8VZ+j6MvTMJ4Lrzp8OpsI4N2HTfJJQ5H2s83BTuLGPhzsLmqTr75rET
dA3MMDq0uazyzwxD5XfnKe4UG7Ny4oa1iZIGlxNEAzuAp/uljaI01LSHLpmq
+nx7/LA/WymKhWJUrn98AyzihmiT7yxtfsXVyZFqYAUof5BZLlGnQqnoi3CY
agxdADaTrZQVGS0EYJCy4AZpecF0fYt38nGuxVze8FL0ElwYbaIv6bXCmyug
kv3XeI5A6siTaLygI8/czl+fQYf7pAcKu3Z7EFodyg0sj5BNgLe7xoSN6hsA
/+iii5m/Wn9C39b5KX0DsY8r3Dd0GiO1iMuVBzhjadKRUe6Uz4CGigxCgByf
+3NAiOn5Q+5P54FWnkDDLqQkdkFMhg6YZAagcseIrFWXmXmDytObijj+BaFK
uqEOUTiU7GZGeLjt8RisERmhaYi4KtyYa1uko7oPT3uIkeTiiSa6jhmLK5G5
DWIECDrpvUW0ZJDmQV00DUsBINvxNEZgbMWe/S9Br26Tt6TpSQ4hGpczID9V
+mAQ7Ethp8F2ywTIePukpYUxGVfRhdAiQS512Aosw0xLVwkfnajXV1XQdVwu
pTlh8pPGchAY8A3iRwk22Y+SpBt8x35x71pDVxGDaoR0ow1rXmokVSwRq8Z4
1WcqdIFC5HPxKpXwnM1ylGdiazsVJxzBTpEY9q0mbS/1NVm5YLnZDobcjKZ9
ZWtjfQLXEkHJ8Mk94W/95kFG9OOZiiJU055r2RjW21sH2g7baCHg+fcy3GBZ
jyuhq7So5fuBhYGQnsnarVMOJRIlLFZPOTbzlRCwv79CT2lsViGCXwXsGcRi
HADZMBVdUpRg81fDJtduwV5IWNK2lrLi0qobUVgkfO9G+s27T6IwQHge/0k+
j9uodRpxlR+euAetZUJCX6TLePRSArsECgfFJh63+kxzoDAKgVFNgL1JH1uq
zv4jIqF9DJEfJOez+yoEBemmkO6m3ORIm/k9xsIMBzAHppzw3CT4Ya0bbDJx
w/TmzSp2bjyvvnm+Ds7eoHBTVncpwvXAuOEfIR4pIPTJQcwqKPFdeuSki6XO
06LZ7gH8rn9GB5nPaz10a9XvuCJSTWd70vB7On7HX2VUnSbZUJMgmOLA5jrZ
pjXGCvYkRvol8QyBvSu/57FYEf5nVMs+8OvsY+6P5txSg/GsMCV49PUOVNSu
5NvEMgVwYoKNwqK4/JjaO39HIIXffRMPhHHVOLWjXE7DWr4kmB/91nCZ/f/k
PRYmiOgQ7nhl2Zahq84em3xSHq4SzD9khZx9ETZ7R4DjQpeABsE9OHxcfQWP
MB6AdN0GyhBqb3ptxjMjezn900YBc8BN9VN0E5FT6DdZdrDhpdbtiG+MrhKF
LPswIIEeZ2S9ifBW5PR4cjtA2WkAeQvTbnzIebGnsZFdkZm2//A3SAn1hMQV
p6plDkQEcTYCmYW1iQYverfcJUbIRXuSCcgxfNfG+sgDh/x4tkhP3DsjXvsh
IdojyJ/V3DVa3oP0uv65dkOZ6tPIoXFP7Tod8wsi08KrdcHGnjyvaQTIMF/+
jQu5oX2k+/iZveCG+sGjDNxKukptXCSFWZu4XVxPClNL4LaPEgQw2CdHDuMv
S1Z2YhOts5fKcNa4vYJ/80qdskmv9S1zLgeqZo1iLRcyyt+g0KMuzA1Unutn
i385RMVuSWtd9mNukUe+r19uiBOv7v2rl/NYKl9D73BHxuiflKnbfSEWl+kq
mUfFubxsDZBFfDuptnUDsnBLawul4GtvP6Y+YgJTB4LkzCvBkSxhTcYrehje
VTlrfIMpJcWJZ55HjwFwd5bkQDPIxaBk6or1sd3sNWP8C3ajW2tdPmIB+wSi
Z5ZO12NWjRtQeFdxmQuZezTOJVqzbpPJMuK/E5Mseu4DDU15xDMRwZVTOCIm
ynbf+s7aw2Gw6Q6GhBUYN+eJkaDkSqdLerSWO28+G2sW1fR7xywlv4lhRo7f
a1xrCvDTJj1cH2pDJk9lSKGDkQ4kyY1ABlwAYb1TCpvxz1SWMJJ8L/GIkaLv
XQxy4/xg9T8kfI03piYrarZk6BgFrravaym+rEIcU1IACGCYAGt9ZqseE9YW
v0kb7KaatBI/kP4UNzryQTW5eCuTJ216SIKnBSkgm7W9LDqyhdazCKWSDvow
OXZvYzQN+KqhIPvsScvSHK5s8FJ512pfgjNblOSZ2WnfORretNtGPjVRjywK
TyqjVaECzwd7ampFgZypZ5Ir1C8Mqm55tOVG1whxEi6Izr1gI+C72/EGH4H2
TbLQAkuV4+MfFQ9mZra5BMPppP1LZParsHd1JHJIEOrpKoOsCGkSKy4XEmL9
4Eac5bN2wK/CWw87kxQIOgQYLi7G1HGmmIgGYleXxc3MXYYxemMPOpMIYZuW
5pePOtGtJdX0XSq5DztiVF+lH+h+xr/8EOtasSNDGzqH3wcUA2LDYIfdCJQl
tuJlQWZ5QpTS2addz0R0JLPkXRPgIKGuMGbzxzgdvHDm3oAS61JUhZCEaiXy
0dLomc2iqCKkKOMj8BrpTGz7JaeEAHlqzA5UnaieMXvyTnci0vPmFNF/uUTz
aYrJ1/Z2IichatWJhXB2fsLUYlB2zQwL1dFi5Rm8Kw8AhgxjW8PbKcgZYoqn
yjiftUFBAEkvcK4VfjxWqPXN3DfMkaoLRrSf9sQM+XRAY3ua/Gs/EMzG41YB
5vndZDQ8zOZbmzLFxO71N1LTIVwGYlCFP6qI9/l//dnwCQcAxqzitWqBXpOg
qxxewaGMplV+yQL36cZWIViryb1kDpYpIR4Dung6U+hsZ2hV+eSSqR1jpd2l
G1+L+fIujmm8m5WORlDfE7K50LzPG8mShjDNGT/ZBaoLUHQWkyjON48bztpO
XfELWZeDee7C1IoZBX10/q1z9sA+C11Jd/O9kUKg18lrETtN6kmXKMPn5pcg
6hle9pwxq1YMW3nrF6wELScHkbBiB+N9Sgihy1+qWgxDoHmmWthdPyyiNlXG
bWD+3WvxVx2v33ZNNVJgLouRiBcvZAM4mHwCtEb44a0uxkndTUl+uUv0qdp/
bKrv1RsoG3CA+0b02ZmDxsEnqAzN/Udcy3Ekg+5y2o56hZmfG/s4j3o4fd5p
93r4TAcIru+q34a9WEq1h88aP8UJsp7Bnb6GFRk4ogxDeCworTr8yGvbO0z2
wXbcL8UsRqT0Bz3E8j5+3KWddIGhY9A3ITcpaHLZbfXGn2/sfWmaLOb4VJG8
6EP5hyJXL+QMTbyW6zpZJ+lrfTQaXzL3fhPaCMx86CzZRYCLZJKS3iLafmuF
zSiKZqN1P1OpBHoiMraBcPjJ/3K1Rk8H3Q1CeiQxhPHtbQLbMgr90zIyl597
6uxvW/dArJYF3WxePf9ACWQzqeu49lpQE5yi/kw5biaYDE4YGjoXxrASvPZQ
zP6C/wxQKLzyEnb/F+S8gip3WIWRr6N+TvutVSSFfa7DkLFdDbHmdLqJyb7F
rzEnnlJPGcrYo/6D920vRXCkCf8iS1Cw59CeRWzG7nCn62noeouDzR2kukBn
xUJpxSbIaLEOwd+D1VTWBBOVLJmDeHI8naSykhSP1ZJfBiU9W5yhrMo2D4pF
xGYe55yrCGOoe6IpEX1kgHV9tvKejUOpV/Zi//YXenI1kKrxriR3FngJ0PuH
ZoIB92Fp4K9NUFKLT195WDYvjFlqdH1s+wz/Qm8ys/taYlOVbnibPsuGgnCB
W2OVEc74lWVSFkHs44QSEWvqNUBYWFBmbbdjO9sEykHZg61qYFaIMhLju6yZ
rXdEv9jCSb/nTTFAOlkHr8Zgzi7y1tiAVxDYV6LJwO0I9U0D9LlEyoCctrav
Gb2esk6Mf8ehbmdlsOVW0NFpQAsht203HN14XcYD2rtqhzEPXcnX8KI7+vhz
uD4D1T7TbW9dEQ2IFv4eXVkXzf3+caz5jh48aI6pZV7AGDRy41fBFlFX1AkB
K2VeoGs8gpH5aPa+Ve9tX9g7Jn3T/+NgLYjhyMwdomSIFebrV6gyLWxRyce3
Xfd7eIeVDCP1J1HVVAryxCxqcB1B7pCdc0OVGapFzFiT7wRF7ltAgR30OnDY
Tm8XSY+Kv6aYxof6pUongvH4k4vPgtDDHZgcw9nRRGEstUIBto3ztjR5KlCz
RLHbqEkN6YLUKtQB21MNSYnIEFPyBLKfDZ9yrkzaKzmRgT5KuQjU2RPG0qTE
jlUDzIIj1m5oy985Z3kFhmx9WQPQ4Lm399sTJmeDi4FayOiStchLHFPBEVVR
aK7xBiT1wb9n+SC91DiHGxBbVXGyXL77CiCEWD8PhEi43K01i5dh1eMGq/7v
KIFNEhyPZ/jIbHF48coFEpa85Sl4oDu49Mc4IbhvOqX896fU7YwVYP3nIcCo
U7Q+Q0oVqOAVOdq7EnyQPNbvzxBAxx/k/Sa29N9V2Nbmc7qkJ6Le2G/0zVvU
NHyUAV1ekaf8OOAvuHLG1Xpo+mDHoxkUfo3fz93eaYh9AFqGCrV/Cteu2/qc
dLfWaEK8BRqtXthEw+BELlFRG5GdVbXquOSbCld9FHofz+A1ImDPtQ5hiNtj
SjtxXu3DQAb576YnjIFGfVCs+MRxC2LkDAlxdLVeD1gj59y6qT45ucgSg3Mg
54v7Qbg0Zt6U218U4ZTDpk3BP2gXhrHJHDkzWnyO9b957m74vnbAMLEU763d
KODymiWDfCXNrXKBbNgpVXOvuyJEQfYJXDByWvdITwnt1dnX1eI8bXWyWlcI
L6AsfLEA4qdcnKWnaqAFRfn/nTJKVhyug2psCZ5c7A/0LJM1gSkist+koTRo
hW4Bbe2C0K0OR1Lp1G5+A6qiR+a4GGiC/ZzmlQuRQsQMQR83Aet71eIeQipz
zEW53hpGHAP/uya04Ojj6bKZv+eCMDNDfhx1k06uUdEzI/MOePny6eu1fmWk
QjCUJVpXRziADn7TmDD0d1xJDo8ModQ0L4JLNSEIEopBJd0P189xqleR3Ffe
b4u7QyRVERkwMIA98H6+CVBRhUydtXByMycIyzY7uiyCR9IJbazcJiUImHOP
0emCHVTl8xcw/DDwU5605IG+sw5DaU32xREQnehu53jlF7i4YADEOovDOCib
lEhB4ah5sEJ1zy2C9O87vqdCoUnVaBPA6eR4mwXh7xyLszwxVLP/FWagC5Fy
YPoFNcRTaiytunt4pNl8YvZovbSWzDnvF0q3JqM1nZ1VctqgTKHp6DddZw/Q
AD83TvV9eBOPJZeAH43KPAQmU83D/T1/eVahObtdPHMsDUFSVC2pzBnn/Id9
KQo5rGe8eofD1vhhupAIwP5lb0/dw3evw2VJJoPcRacRm4j3pODxUf4ITmJI
/5193swxRGbrmi+naRzSmSsUKMQkixCOoyhI+7Qnom6aiZBIJiGOSjXGgL+P
fkCdZLn/qCcTNjwmppPj/wGrEwxALq8HBYc9CaAoCECbN32RaFhPxDFteA+n
KkeW4X1wnKL5ALv9JBZDXD5CrDVX4+gYWGPT2oeiIBboHZBgHfolkz7ypTgy
9mM23dD955BwVjCJdrJ8Y+0UXAeQrLazd/+ckcV3iELpBHE4zr6+LeDJuyDM
JhOgYlpBFqS2osW1SDXBwQWeioqPUeUt+fpo2KRA2lavpPkW4MYTTpXMlzqx
/+xjrb0RyI3YBt4DP/hK4NlNbGFGEbV3uMM4PfV2oW9HSRZmZ9DdE79b4gSb
jlljslG4lL9e/00/cuamszNUQv0wbNiAYPqWMaq7Ry+GwLWYPiZyvLdSzNXE
kcua/+dxPIkFHdJ7nrR2tZHRdDzw73kNDb5c91jamVmuuf41D8ld/Vs/naUT
kHtKJwCEzqbKkscGJxixemThjdBT//8dwwVu3njISbsGmeYWiIcL7JI/yEYt
OuQ578yBIWCgLsngD9idR2/xAqMe3KR/8V7I/7moN7vq6mSebMY35fK3lxHA
77skHdkV3aEKlLAftX1ln7v0xpEAIeNmCEkxS2DS++IeU9eomyO7UIT6Xn4Y
mqqUZq/rYUhB6mR8gHpbbUZ0yi/TMhOUsvbycmFpHV7IQsOKoajyJBqPsFRp
HJ9dGyeaO30Pk29mmwSAfnoqAEwDI8oQz6A2DmDNycl6JaSKvHxEe+EogUtD
0TGOP/sSfDYP5cJJAFRWuVKEF15BFlqYtsMRZB/wiko0/jphEST0DwblP93V
vTz18LwQVwWQjfWVYve/zmAu1BwmiD0zVhRBoDClRpffGzmYROX/C2wAYQhi
cRmnemnrEg28e1H+EtupbWNHvYOldmbqp72l7XF0ZvUpSYUPmI5i4I6nssw+
tWbM3akCkc0lb7WyR7KmQRPzZjYZiUuINc2KMhFCTCB3XNJMelth9c6In26T
AtbTITX2+EpoI9333PKnwf6+jQIXjlzmLXLaXI0Ng3BEVPdgbgBMa24J7FhQ
ccbafo072ig0//Oxa3IGrBQWOh2xKtMk1lCoZLRkI2KjWp1oeEImPQ7rOSXN
ZkBalpm/K8v7UobV7xNOM557DeewBFIr81KjdezHK/RjZtsiaZBsbm7tHw1s
xgMHz5rnENAJ2zEOBopVZqGGF3EmHp7rsCZjY0JsqbvM+b2c/v6IozcHZhNo
2OPFdRLK2/V5qiu02fIKfZwP9RL7VCe9ZVcAK5GiswB5fXlcLugU7XMKvEPT
9/QG0BO8fTiQjDp+Ou31oq/3kncXHokgy66LJ+8kuuL9JCJAqAQXG+2M6TfL
yZ2JQq6QH4ENyhCqmlEO9sep2z/8X3T+6JE7KPjY6BYY1CWfzIdv/KDddqD4
65j5CMF5jp7/PtKkw0YvP9qFnNjVB+K1pTgkuoEh6CoyK/0s+uO2iKrqMv8M
myOt8+LIfkfZX+B8HtBs1MiUFGdfQOF/s5tjpI0QGeK8n15nNLifrjHhUp0o
qR8g8Y4lgu73SvUBQm/WvipBVxns2GMItyxrUQ/YBOSqg2+ZYsAT0h88UjPH
Vg0PnetUrvyE/BWMjxgBfg5pvlQUe3KZvFL7Yo+I2jTjrKXosGLOV1WIFY+o
5Um5JOz1yW1IRL+hSCabGIZaGUnJqrN2ejuwq0uQuefsm3uU/XXgM0/vyzxC
9VXmUO3xX7O9apkHuDHsroia9yi+9Yf7Nui/t2vnUS5OWynjpS6iW6ZasZOD
E8FtLArelXy2/yH7mIotaE2lUbvngtPT7VyEQkK2LwNdDwac/iwst5FgxYPb
dO8lkim9E+bEKaFyOel9bX3sznKfI1ucfdzKT9dwhOewAsQkl56Rp0XoTjuZ
akzmjD4cTr5IX3PLfzPmZLCChCBleD1DG/z9jaWcf9UJDtYY0OJCNt8XWj8f
2e4XqENPVf7ro5kT/okdXHal8q6B8ykWm9iLYi5dXhdV46DZROqfm95EHos8
zE9843EbpR2dOWYOnLNWrBud61JKdXeJ6OF3xCgPESufPaPOm7sbLTJyLBPq
gV4XhcB090WHomyr6oSqxgdmaJb2Ls16NrM1x8sotwN9phHB3t7ISkf3lUZN
vYKj73ze4V3SWxH9HSkUc8NLPI3jsFoh+8x74ejK1CmQsP7omj7J6IbSAHZ1
IQEgFo9Ww6569DAUqgcxeA0yZBGkJXbCoOBD/Llo9ZHsQbgLiBADnK+40tVD
jjom3y1xs2gB4PIaLyB8fbAZGpJ0RYmnrZNgYpKSCpONhwTn34hzWs+phutZ
aBndU0NoGy88qAqDnA4XRqUp97GqswVyXEV8hI1HsIPhSScUpYcBOxtyF8mh
+xwQVbFp97s9RhbFN4WD9yn2NiDC2E7aESinHPl8lt1UHNqCIwjQeXXBhC2K
T6uAFzMwcML69+4vd6shMHWZEqzbReZE8tfymCpkcBu44vsBYywM4W0obmx/
cd31uIrXJLHobJX6R1L/1IcGYoL7ozoG0iGIEYEpNXGwGQZm6WnwwAjAYnGt
8YTX4ePZjX9eW1kwkvcLurcFebr1WMLcQr780m1TyWoVCIu9fxhJJyQlEgr8
h0hqa6y/w4Xw2h+NruZL7pOfALybeWOpZAn1aJQuPwEUshk6iusnbQmVARzK
lp1AA+prMK14eEJmU4FqV90Bebaag8MYuyVf878L1TNELnuOIMxD4cyN8AMq
Hq4XIj+PnVYyEwoawa5jNvV9HIg3fgucri+1LhenQr/2Of5qRJmIgDfJDkAv
5r88Q8nOjWoPsCennPwfIwmRaG4gO2UHWDxjME054LBPwq01LbO47T/Qa06F
A5mpdFPiRjxmP+sl2ZkiwDadsY3y31kcuGkOnCZwZhXD6rJIkxvrLNbBxup1
XMsYfUbYJxZlFSZOYAXmtelQgxiWfQjXkVGv2RNEE8cfcqP0YZtZueU+/Mfj
SKjvunDYYSIRwLzWRsG5cLFq3vDzVEdt0CXwMpkX+daF4dRt+JGxmdZ3lovE
lqFKfqQY310SR+ipK5CLoUh8e0zosPU26kgtt95etQhPHA+fhYXASzzitwle
/vA6ieb80R+TExlYLo9TzO6D9glbIrYyV1UPBM4FVMIP7sVQJ5vc8dZLOPMN
6GeJYapUHp3hRsfed7rH7ZjIPioY7lWIQxrazSQD54jJ96CeUrdyXzb8uNcZ
3AK2wyqCkTQThC3i32cETb1nYfszEZZ227xJInaPzX+QhLuZRK+3/tJt+liq
qWFMwiasEFAZpKT7ImaN6m6hFrzMjcaH/SV6fx4WINgB8CANl8AmwebNxgDV
92M5IIgndIQ9p08TNBhtfrwr3lD+3E5AbaY4SaaFCYGIG8xQcVYxwqvO8+M/
svXYaBWfXqweDp7exGL6mZJkOZ4dt2yNS6Y8vwUKiu3WNxY0uXPLdhI2ipk0
iGPyXgGpfL3UE+BGlumv0fe36+UaBH+OL9kJI8M38uv+zaB/FjN5J+dmfpMj
u58gUkggVehLyTn6dOyZ7hx1Y+C99IstIMMHLAUnvsRWgUtqEHI66MDfnXWI
6HH16Rsgkb6V+RxlFITdXQEU6kzcWL8K8kpvdGJ12SI2lGrlJs+qMyw8RiaC
+Lhh1N2d8aL7LNWkV61rwdWZ9JIuQZOPrc+eevRzVk9x2i/jZRTCnUbCSS7/
uRm5poKGwffH52VC6wc9p1ilZd34YoOJEGsNvM/mNWvcsmTUGGcvgWevZ4Ao
QmrJFAVrl6HpwqXKPJUEcPzgnEi4Ui3sIqLjYqJyYS2u+JKbSeyfmoRJVKOE
HugRNDH+Rn+D1+heLkRFiNQoHnLPCU1/NmPkTwOvZbZGWVTtwTcM8fd2CA/c
n6n6i2NDcwUk47qogBmYhLj4k7Z3NsYpMsqQEeUvB+Fc+wZ1IfAHmjk8YYpU
y9+Ba5yClsATBv8Rsee66AtPDPgPRZfWTMeBQMqPmzokFE2QFclWCn33SeoS
bXoMAq8qEeAyms5MycKbKgbwDDPXsn/buTg5TaFtcGeqfJquJ6QigtaKeV4S
8ewDN0soi9FesAvaKJjlJjTf2KjpeqGYDuaEIxQBPpmBDOLAfM9DjcA+Dd34
n9erzeFvmXHOe94AGUVDRtcBw+nIrg7V3b/6kIN9hcb8JSR9S/J54dJrcg+P
Ixdm24GKMMn9Q9kHosZtr5+zuksWGGq+dZcnv8NhuSrY5+Hiva8QlvzlSXpr
qYOjwdxALZMOJosxHq15FbuzkStJb8HgJ4z8LLG5dBX0NfF/w38C7R/nz7gn
sqfzd1YHW+PleQwzfIi7HqgckS/TTHwiqd8Eb4D2UYd6DKrJIzSyc6Tv0HOp
Jfn6dk5G9ATdnnrmtHzt2VQCooko37W9dcy++Jk7HmmjMisqhphms/+IU48l
TdxCAKNL602Xf+5DRS8WkY8/srNRyC31EE0IH2mDvboVfRtR+H+XUsTfLA5R
pSmrYBjkHNDe3Few8Gbmd1yJn/rcx9ndbg6Bkla4dr2cMt95qH01oKhJelBF
lEHjScFhPp6BEWHHku5HB0XZXSsOx9Wy2NkS5jrKQ3XUWAkAAHtm2D8XKKzp
6T1UwlnRCTmfoeaQicZkgvrfPGgNlm3tgshsOigX9DIJLFhMsFm6HLlRmTGy
Z7dnPCBSJ7ICskf7GiUeyGIsLrRfwN05gOtyVw9mzxSH8Pg6voUxwA0HyGtM
s5TcsDapGOIIMqcO/VzkQGl54Mr64RKoVq/AvHdmc50Uhns8Bm7ILARAivrd
gVy1KT6Irh3vW8itj9Id8S/AWQRGJmy7k6IPIb4u7Mb25m8eWXs+Fo8R4yq4
/RUQ+XkRUTVoOYaOJT5SdpU4V8lJyEg4ZjYRmlHKht+jPoAmszf1SRBIEUiB
+8+Nr8r5xQQy766cakbYsJxSYNrVRpPssw8IIBV+yYlQME11NSSWXBOvFD1x
5uXiBS8BG1wBGawn44FV2F0rBpxxFIS8JvG8IUh5zsC9g4xoqENAivuXnxzJ
JBjJHOxminZFHcx4NKsWIValZiXAwzsSiE87cbiTHbyHkBe7YR4QjS7ITr/+
T6u55dVa3tS93S58KwFQLzN/8J03jpA/iMw74dENnkFx8kN8HeiGq64zIp0W
R32ubub6Gnr1JzA6XMFA8kYqD0JL/YRtnVEeMkf964yTDsFvYKePpY7oQoXf
IohSrTq9G+6YTxPxrcShiY4v3CNrQaXy6neFCEv2EepFrVyieZQ+/MJH5bTK
aVRjy7g+bgP1WwxwlC6dL8VQqscJmS1vxEX7dOLiA0smx+OSS8EYCiML67WA
tVFGaqSXhJQdd0eQ+ML+SkiTquYURi2dWpni2eesIJ6P+KZZ8HCpO7+XS9Sd
CEW5AU0Zgnr7jbpak5nQBpXVWsfrdGm6cctrJRUPivlRHWrjHyx2LuXgJcMK
E6AnS3YEbaLOD85g8e0s/NioTDyWbCUnQD5DCthE26eZdczeBOhRTk4zAmMJ
0SMGoDQcdMtLGuerH4VQgE0y+LFZF82iDbRvhBourlt58frWncqSQTQIZFvh
fQgo9d5BkMT8v0s7XPikCXB06LKRk2w6QNfg1S1MJv7a+neWtxD6Fn3a5lxB
VuvIvpHm1+1FPD+zYc0SI/H8U2nMhdC5JjQZHIecGNr/AglshX2OUeOey1RY
Gt59OVPq7aL54jgsPMZcQH35ItvtGGp1yExiNDjPQGhGzfgpuLzjIs0Zadcq
edyUJfqKYh76UtuwWvFZBj+Qd6oOs40zAPZnzNIi4DOkpY2Vb1COBTOI11Id
VtRfdqSpn13PAftsK//e2kCdB09vfjjsRcPZN95rHGIs7EJxMZM/w6dfPkyQ
n6PJJxhfppJaXPEeU+CALBuUVBg+rT/Hq+z9Md0GrQKJGzxviUdP5y8fncGU
bBKaaWTaUiFJCDzRD2YioVpv3Hxt4I/QUWqma+NYIb2zBmN6DZo5B+SfG5FP
Hw2rgNYp4nk+Y53vd8aZwM4KbJy86I+eXOD6V36rtJhm3lSZ3cziY9jLR0iN
Q/kSfFlbhu1RAsNux7/7oOQBnHrtX+mMLpLEZXewR1JVZ1X+w0QLPI8njsJ3
MQPBTgxj7oro+b8nE5N6yWG76EzIR1x04x6z2EAK5mfgoXHChDpt02yXEA9g
sxfAkFpAx3m3f8Mn5U2qkXgzom5XbPhlniYWHsrdtLmwfGK5rvAIU6VYRbZM
3oTGjbwtsVGuicUxQgD0AiEVvvg6ObOZGPYX9KfySx+rWX2h8rDECeUfGaxq
KsfuNDsFBNt1IG7M9L59zE9d1R+jVPWO1JIJ5Evh9s/RVKuVNHqc00Gb3zIs
ZVyulQxJEybXZES6cAzsU2FbipekWzrJJmk78IMOqV5PbN12dnDeMQpU1DSO
iY+QSebTKIRC+3RZo+dAo/YSgqFUU3JGOFVKJ8hjk5HD5mE+FNNbM9SkuaNg
6qN7S9Zppsy4uPESjvBvmpt46hnL3X5GrAHT2OllJVEr02949X5Hbbc1qj4h
rMHenCo0goNv2iNKcWvZM7BsxCKSU7KaLSeqywJdSfhVOyBGF2oTkV/zowP3
JSzMmxtuE9Yp3hlmrONnCJ5qG5QXvUSKv2aRTTJTenGypb30BRk9R7DaodzT
uOjEg1s0VRSV6hR1sZNUmKNu09ecYgApJmBMnODr4ENOBOmN7ph+zXgIZjRU
zWviL03Ip/s2nv+rd+E6hRVKdXTag0mcLsJqn8z+/v2OqFzf/qqgMrHc/Cia
fGzIWLMBeg3CRwK3MZo3nkYWaYXR8JtWm+magcwCvB3SEd/pT6il51wjKoub
2+wCF1bX100O3JMRACHeS4PsiJjQzYjg2TQVgeedbsprw+kxA8PZnNPJlzzZ
2tgVrEwqWttQ0I4tKDHCs6N/b9kERVjgetb0t8n7EkLvdyMq4wYJDjHlepT7
/85kJS5TapJ5CsmdQ33C6hj2V4cm0MMEMF9GQjqOxFbOTaF0NqKH5c3pyDzO
mB2J51k7MrH7cotId24F5GI8aZpUGswYsXMUE1OObnQRI79jIdcn8Uoi5Evl
VHiuRhHzYXQQTJi0b+8ZhnwyA3rsn51/eKOgojrxKfEVXY6RPHy2kB3HqSze
BHxPFPdZtpH6+H0WGvyso6cf3765z5OXCPT7fzaPBKBX3Vj8gTz7gIxSjiYb
ZINila+RGBy9MbdvMmuy/AqVKs1zrubF8uln3MlcdhbGhR9M7zbXFVo21SUl
HcK90TgQ/NjnaJp9tnGTFtygdLCIQEvw3EKYacDu2Oc6RQ4IkXZUa6yGrWRR
LcX/daNXG8DcEpW1hUnjBx+iqndBoipbrGcylTcsYoaAq6eC6yuLnZCGgroz
ZwFbZC4BFX6yBiWylUVFwqbaWEWLxYSYySg3KcpBHiVqZZc6zYW8059wLceV
ZLjCxmIDBuJZ/2VcBaR6HxX6QB2xE+Xgi3pjNgmYdRw5npvKB/J1HXxUK+2k
x7c0pken6rc75srmce1a3iJyZT/HIXBg2WCKjCiN4Yl29NrhD6gXbYo1+fFL
ysWuhytHwY2YCaAZROAFrYJ637onDikySYIqf5qwYAVS/Sk3lWMJi0UAniX9
WXzkoiSZhObJQBSzxETsbbzGmseYlpxQ2E8FXUiosKPC0s7wtm+S55PH8n9e
Jrw48YWeEI3jZDLkakgVdcGy+ky27newdAw0jUi8+x75uCBfWwWPA8ZZUeOH
0UMrVNp/naiEOFw0faDRFwe7i/LUxxY4ru5YYNLnw71mP1o0gUmhGSg80GJW
9VlWEkCUv5TSplcplkmLLn6YWht9+6u8jrl64JUXOKGR9VfiuM+pox4XPg+k
Ij85T/Dfxk66r25JcHOJMb7l01PLVK5I0K655Tei6vB9Z9adyw4lNrA15mci
28Nz7cwmtNqVUleuRTn10WupSNkRDpdS1t0HRJRDlsYYqW8xqKz/kDxpdfHV
a6I971dHYZroEqB8Z8qajHaPX45w0IYWhZBMaTv0I2bvkPG2AL0iwUUn1FPA
D3ZYX7vWoQ1251dxNnhWPWINNxcWb7748gxbeQjVuBkT12T3+8u1jw2Uqn1i
TR6xA6AzvVmhfsJjcrJPQC99dZPxhB+Ix76RCO2OV3K5aE+skwy9OVMWHeqN
O2Cd+L/aR50iZiBc4BuAewWk/CqEkkPvlWRK/+f+yIc4Bhe08jOsoC6O+Erj
5uOB7kXtr20RhcSXxWEXMVfCqq+B+4/pp+r8oqLJiPonzmVaSNwD6ZhYuKMj
hS/UvGgr+vCBBIAjQcVwtTOmvyZpZIYhh61cyiooGBuY0Vu6OXPvgZVD1KJe
mQ8OD8+9l52eoUPCq4AfPAMwZ1lwhdQlXg7tog0mqbLcGeGni7Hr7d6q5+cH
KyeC0X5PzCb1N0Wn1yDcrHAMF6qc4qpkoL2k0f/FbSsjLVFcbFbeLkzsfqJs
9kXT0QLgA0MmX8ks04Mxiyq7WW7AGCucwXDyr/Gck1j7MnKFAZwWt0DK3aRi
wEXyCoyN9iYy6WCk2/7l/kZBlpjgD1BhIBH/SrfaVoadRob6VE97afpM++Gf
LxS15+CwuYIDH0x8osAI91m73wP1t7t8733+aN//Xh6grtigscNXEoOWfVhm
EkcMWlK0HaoSe7ccdHoI5dSUw+FyC7RJn12zvAj0b3R1SgSuyn0yQ50I7D5o
1ok7cWTrwoERcsO/qA7Q8NA/u5l5P2OPB3KYd/O4xVmyewCEcHWDd2LWZ3nJ
tfJPeJFk336i037M9y5Fvn8vdseK7DqMwYFSNRCHWIEJ5+roFO+XCOc3stxR
5ZB6AK22qp4C/E+zdDr3smtNwkM7uhhXACWQ2dfxOFyeiJlgAtTAigtSVf/W
ekothS8MzeqTumUuMOMIfNiFVaQq+Ruz+sU37iAoSdvXBtlcUxucPQI15dOy
e3Z+61IY+EInDnzr6rLGSXqBXlY6JyHZEaI02aS0NAuWF1WUXi2i7XtNQZso
ytTFyb0jrb33wvZgXzqpfgZEo64t4xOq4ANcx1+KMFyTFo5ejlzkjMzHx71l
gY9qadJs+t9Ms0GvU453rn9Ipa+F+HD7xo9hkzlPZG/XK8AeKcMdSQmD/Lcl
Fd//QYR+RqzWx18RtqPCbfbyUaoHXQ+lTDL4RTMNXrI7k7OEOj2JRdo72kOo
AEyaXF6cprid3HZLzfRkG5bcXSUho6Whiy3Xf+UjjW/eEiBREVRnYKl3Oa+g
XbeHCJ535/kZDl9iVIC9i5owcDCq9SVXmUlOQOskn62Q9dveUDyIZKib+sAt
qFE6kY0o1QmA9hAzQHHWb4OLeGoKkLSudN6OwqyAwdW24h/6HYjSTgzA43CH
Ulf1ELVB3z3uRFDxTRB6bqauxtF7XOl2tssk4qz62hewVDFJcWzPie1vGTHS
yB+kB+GFJdBVZ28++9jJT8Aod7KQYzZpFLJqofiuPR0AXPLwWCNNv5TNSnrc
sN3b94as2zD9oG55f0iWaQeMdR69qpiRcLVTjxTha+xq98wCg9McTSChpKXk
1EfrH71nfaByETGEp1eRmIe6ynF5ayfkcvTj4cxWmMjsOLJhL1oG1Z0l9YYa
sqVAbZAickenOx7/jvqXVARqbS3rydictvkCC0StmGlaMSdDSRZsyGo6e0oh
rOQ3UD0VPoZPfZn7dYTtS5mXFPimuzdX4Unyd48XfyNafomuZkyYGTI2tMIK
oVEM21hPsODu+WQPDTvEj/fT624hTPKlT+3h84W+Ul1G5VYklwXTzNaY1cDk
3EnkxSBI0/3HrmJzk2HSfl8MxDxALmg9vY9hq6Ba7R44bcVnR2ven1bWfkQP
FU7MTIqw37J1mJyibhftU9SqWmeB7zXQi+lDWwarZ9rIT7qxRKdHI8sbTiAI
8UsVy5ejWe0/JMp/UB4ikDdNGq5lTmpyczgU/MdAguNnPE1STaFNOrTae1yS
qGJBYAhCwTS/+TTsPsWYchQawoRy8O3Up3us5+ctA64EjwVCuMTXamHVjFCr
Uakcm8PyauRK6sK7BpLX0kWAHvf0I9kJa9c3YAVRcao7D451Gjs+YjpuwOOn
+iQI8t+2c/rKMkIB+JQaUtUojv+J2KNKMwa0hAgL4ZcJmlWfEduFdFwlALhA
VAz15QW60qeOgnwNdFKyEVIwIbxhqncOp9YH3w6kFwEth/cnacT1A/LTdOLh
Lgprux23HwZyA+KQBT8q9gmWr9fsTFYijiBh+JzPPZgetOapO6UXUTii3wPY
NuicG03GnN1AVfcWS+wq1NRQwG3jVsM/g4YasD9zGcUyzDEMnXagnZ8xj2hi
RskKmMBQzsHYkw80GJYHtZ1csN9nIRGvS53Gkgm/LXvkxCTCGPEwukTuqIdq
c8KO00OeZVELeqvHlNqkqMYkXK0Ss2Kw7dvTnCe/mWTU3oLjWN0wIp+hdjDX
8KFv3HjZKYRZQM4alesyln6J8CID2pyfPMllar6vQJMkQwECyIwaL9+xkVb2
Cx+Wyc9bE7zrSvVTdFw64pTBIuK2Xm6iTwNzljq5f04FE54mivf3Eh7uxkoA
IlZQeqhDutxvV+ZHV8X/OY0dSgh39UGkC/GqsJ5nFlpP9cYy4lKUn2ZCbzPM
d9uBJ6lzfNNUMRWyVJ5zCTyxBrovD6uE/YrDX0N0v9rojscIo4T7MNvbgtq3
wo6c+G2CmkHBui2D2LzB5bS0xJ3JF84chAZjfK9Tp5zUbErMYz857Ns6IFUZ
VlHnoDuW8dBWHCUQOXaEY4L2lMs4MR/k1yIiylomUI4cp2ZuTgYNI+OdhYGL
wwtxwVI8DWIg9EMZxDVOmMQW2AMHUYKkDVDerxPs/PgJgoX1xUCDkq61UI4T
WSQNl/q8zRV6dzcjCy5ZFijxZjTKqHnfvccdIkbbbw3OJHnSEoN6grcMqGzR
nM9D46R7vxPTiPkxqMa2RcHMMA+MEf4rr1udsjYPCic7laGkmmzYg8v58o7X
pzz1OnNlUK1YwBVja8mMNRZnYRvm4xrSOE50S+2UFFmvzVygn9fHh21Zaoie
445dmvRBgHsChXTsUEz3y4qxLQ6vPHrZbAxJlG2D/VnzIMmg/xhgGa5hr740
OR429wffftCx5iMsDKNbOvgHrAcf2ULl6nvZwmxvak/TQWWHqFvnTutC5Paa
BrxZ5PtEVAGN5SSQGZdZjdGOfvZGOt3NjVybEcJWL14uZHA/idaKHJiu74EJ
QqVa+XcAzns7gLurbpCy4Pj/s3uFmZ3ydXEIVmIw5/Z1hHU6CHZJX2s4KJNx
Q+ryW3+fRQzW4rOWwZClCnQtOur6R4HSLsict/3HYSIY4PRs/d9pbbNdVaH8
TBaRXm92Alo5KO8P0SxF/ScXSBqEnV9SNlAhAS5sCD/Yy/DgCx5MRK7WFf18
4NViY+pva05NEov8SXjHJCWFmfuxCltx3cYGoNmlafoWdlCjcOQzLnSVX6+m
Wh7bIT0MV8iI/ReLcHT5WA0ygom/jjpb6lTLXleIjPL5YrVv7LRo2c9HfmID
WtNnPQFn2e7YZiuyscuMFGFHxK9ZKejVZmOgN87pX9pjDvcWhxEPccpqswQ+
RlBy1NutjbTpXhb55EWlBYguc1LXjBwRWDKsyE38FtpXhCbLz35MsKbZQagA
TAfW/HBCotsDgwgEETkzoQPxlC6dOsTusAGvFmP+2lEdpDo6//vR52d9lCvV
uJHU0E5zp9ydVHYa968bQoHC90blbPDihw4SQWXT1fel9NHBw29GNBakQJNv
PJwuE7eUJ76cWIouxQ1FfHFCsQIpR1QHR7AB7awig0hqwrlhUeeEGnGySss/
7jV4JpQyn6gt4hi9EEIKcwWGvnQI/Ju9/h5JPh+nCIApyQx8X0S0ozkBjlWb
UF9r++6MnqSC9AzhyAqDn/2oPVTz0dfRGJ73E3e8D3CF6MAn8gfIaunyiHGL
qW9YYnm+r22A03T8pGq8BR8Rx/tQbiGG5SAVuBCoakgetuXx3hp9CcXfi6Tm
ByuRQIiBDDfrB/loo99ZZPQaG5+bX/gjgtecv0uICZejyKRELKUZR1km4mnc
BPuPxmhBOblbA2UyM0LcpmnG9M35NxrTVelGiv0f+0kzFPVZkkLivc8vJilc
oUALLnWVpy+Y1bxM4es/bAQ9r2YW5OOyQ/SAibrLQxJS0z/lEa8RDa6qR7Um
gO4cLajAJGhGzOf7swOO57NepCgBH2tfsL+DdKH1gV6mdoA+1f60Xt63zjud
YbvN25JTB/jF0U97A3Hjp6MEbIXRcxrmocAgdmJ+lFjQjVtntqsWpWcBPITo
WmMKPCR64DZ/o1NRBy2AfJOMunwUA4M9b5MT+juErWJg+421t57tu6nAb+9m
LH2FTuTyG92kNKflGFbwX301o6l6R0EBILZ0fQZnksIKzVHqa+ZteMesl71Y
uKmhrUsNs6eKzjhPQIwLgC+j1sxIby50ixFEJamoOyxg/XDLH2YdjvPGq8Ij
0q+U0kq7W5H2FTek39REvTCv22Ct6sV34dr+5V9QBs+pcYIyShnOZvfLFvmh
nFWxOed+PFQoMcPlxzx1fiiuCMAkaJyhF8ReG6LEGaMHdExAEfnBePCTRpfy
1qSuNLqwBEaPOCi1QSs1YfPIw3a1+aBNx9VWcEh2INVPkQ7HHkNjKl8QEVSx
228Jsejb5tt2RtXenoc54SMHYEzFaOQczbkpi8lOanyJRVGv3yajrNHgNO2s
SnILBuMPgtJR3HsN1QbY3CqwNtMbVbodin3vzzK1qPYO6l2OOs4VPFIk9hS0
gZQdG+CVexOSBguYQEfYI++qjOiamHDxh3WH4TkzHeJh8pUwYaZlI90OoMs8
RIoezNSpOnSctkGViG2XgmkF4FFUhZLB1yKODPCoR9Ymahv+DQ01p3+nISZh
Fly64muaoizP4H+1BCHNhAKU1BV0SIBy+hIjbSrN/+/kBYAXDk77rnaJDMCG
wz/RqWcNJrwZPr67DSmnoFSi9A0LT/hM+Q8YnCI5Y4gBsV5upszq75h/Vxf0
hORgS4/+mXhFgjIKHj9pxhCUJZq1TFSfsSIkCQEm4WF5iRrIdJ7IBjvXQHtC
msEOyPtn59dNdN+uFJ0wmTzEH1bnrExe6kIn/UgwF3693h3jBKn3hyK+W13g
P8Hk75gt2ncDFLErNiaMI/okuo+8DjucSvxstr7kdlXsbF80k5jMVyqNKUpk
i/JMYgVrFguGi6vyFHJ/FSPQCjppYZ5I1T8y82eTdUfNVCdsZwvOWEt79ntx
At8xKpLD4z2korbobHU5ViikyA6Eunuh+ImXnnJCtJakmQ3x4LljvOwNmZVk
GWDpSsORAUee+jS/fMrKae8Wv0Qn3aCO9Rj/yw/V7/wKaLhqBuQjBrc5lb4/
nXEjYVmRaQNNrYd+QyLzTKd3cbBHc/ZEeGXdRE+1Y62sU9JmRo2gQhIufxVO
31RGPy5RGM3weHx2pKOHvN85eIgfoN3/PwK8JHq4jT4CnjQfhdj0mh+5unjq
IB//WGRVpEilctnsO0ZtnXUasQQharU/vyq3ZU0JGNrZltiAlSQpZp7r26g6
orLwTawfgK3sFex7cAm28x4lVUwpZ00HJJGBSXbVIWwJLcZtDfPAaNSB9acC
K/jsYGoQ31z2jq+xzzLuSjZm/JN+1TSp+DvKhQ4/cDlDzUlBCu+PGIuQgoTt
izd/+7uXt7YZtD28PywN5eL/TZIDMEC5h8ld2+k4hcxTdTeMt5FydgMd5Kun
IKNdhiR/pTKxRdhL/CqCRnDIFDpcqHeL1bwgNZ03yCsIvfKBoqUxW1MGPX4u
vVKqxwZqhAothZcgR2ofHX6Pp2PXy1Zs/vTRARag+QHa98HIj9E6DbVPAksy
oGjhyrcROaXbz1vFyA90q37OtQYhdZi7ODbptZATZUDxGyeRdo2bocmg5GPV
AzjikIVip5qGybL6LVCUInLg4JOwUHw+V5GcVAHJ+qNkmVHVv9MuhJkJwHgc
yjJUpR7OuvAUBL6bkD8n5HxI8vrDczBUkjfHO1yqVQ957GP8xqCdrvhhByrn
/x9Ogq10P6CaLlh/duR5d9TQP2jYou2h1wMlb1/AIJ05E2D7U83R9VLtLXMH
rdUN+3+5FTf57HIhXKfG8iSZs6OUO4uT44FW02crqh2ygJxg72li91Icd0Bx
RK+8K5FpiUTn+qavew+R9mnEN2wyNs8wHi73PAm1XsGLKYiMeMfMbEI+zDmP
gFNKtQokglqONLjHLXct2iSwPtu75MuhXuKgkQSIQUMTV4p03mKx3sP8Y9MR
Ygm61vuO03fNbkEtMzLxtYF3zLVqwqctODqZtq7Fp1ion5Dk/OLuBxl26bbR
Z8M2XX25jX4meSTZ8lKR4vJxpoHCkwZZRRxoSq5g4Lep9Sq4eXWkqbHFjAFi
YQmxAhP1iopPS6I9WaOWiYD5I8D+Z9E9MqBqQzljRRVEqymB3NmKqTyVcoRz
Q/IKlGR8KRksH0GvdsB8+mM2II790oyVJCnF3aQCcCVj3swTynitQxDWYTlT
V/QqnGWNMUqtEeiPguwK9aXLeANOD3i3SGRIkniYB1KUxK6DL4bPLRUWSh2P
oZf6UogmhWJB5BhiihSJzGt18VgX5cvbUzMm3cn+ct2a9eUAVR3ZnyKUF2Hi
jUKrN+LlD4ZtDWQJxzuoovTZgvnmVtEtY5fOI9JIOfHuYmtFvA9HyGWjrEQB
FZCcENMaOed/7DWXkM1xESH2Zd6rxVutpNl5DxvzjRZMa+i0ePWy/rb7NyII
aTk34pkv2diAq1wUszIQWzA5fISn8MhA81UgLR7xZfWc7i0KaOUrw4bYFDfX
eeapWs3400mSJjRBXeShfweFjwQP/QMpD1C1uJI6D6ORbtdnPsShvJ6by30C
j1CwcVKyXv3KnYavZt7+of7b/BlHENFypwMgSqvMgr1XCSgF9YlnM+te2zxL
I1uy2qg559H9DRwnI5HQXwtEdWVgW6WxCzvftIgossrsPTrwHRhRFXRfln4O
GLKbKxtjX6ZKfcp1fF/rq+/XBuzvi6W5nZsg5icA9x4NQXL6zsRqmSGXm1Ck
KLdOwPRbgubFlyBTlhDPBKyqRe+Sf/9Hzi+mqnmNlZKodP9gSpd50bf7TdYa
58kNdODNTRCgfdHchs1YVJaa3Sj3EFlHIofuHcqOsu8gCSEX9m429HtSLiQH
JqowxIqimYpbY0rtTidlhVehZL8hsnbadB2Fh5I8NTcM8W+3XVAz6AVGGtM5
SKiGMa6NJCCitfp5qNz+c2BpiNwPqOQE7MR0rf2y74VYpUk8rkNCgScFXVlb
riY/HLzlaiA2g7IX92n3pQWyG1H7uAeRQt1FcDvX5JWGyv+m/Ks8suZBVaZC
hzbTBKnlY+ka+o8uur9i2Dc73peQSmj5ItAvKHSxpdZoDwnbYije5Y6rY1hw
wDY54506x3l2vYmv5Vn5HTeaOiRNMD1wVq829exVfBtOu5jksWuqDkVo4Y8y
UrU0XXXM5qrNWnYa8840TGO+sUbZFZhYcjAtfsb3liu6Bc/ZRzM4kasteZ4R
w/vMf+3GEcO+wlPGQXqbIxRoH7YXlJQ/bTKg0NPVCGuOgYsxs3ESYRcrwFHO
xyk9Vj4a8qJfEhsTQLrxeRPfEbsjddzjP++cYiX5oVJuluS2CHDdEuRKuRra
d7IHlTc0qJpRO7/PY8pB+ZLBbyjHpsEwursCILGuSCQmjYVYeUCu3dvN/aIO
s9EEe4oJQZy6F5Zch0lvWcfxll0tN5cOfrHUNcy4WT2Hu0ixI/rvsfSaMakH
Qa3VxbT25ifwJYpsNJtB8Hvfr6Kc69mIowNr96E0Cj8zRPzXiEqnHa+jMqQf
4oi5VPAxHoZnXuBYiv0uH4f4gPipNcIj310rSvUZ6UoxmliMIIzusjiXjVpv
8WMebQH4kYI33tJrZ0AHJitXcBg5sVUOiuS6UkfgjNcXz5EaIxTbai6hRaOh
T2PEJaazgVZtKUdIvfi+sQzaWe2O1iERUheE6yBbjUE5GNQ2ah4zMxBu8eRy
O0d7VzZi8w1AwLtd8yaHNX+EB7ZqOsN+n2r7Z6Cru3lzkodEIPgykbp5wf/B
dGs3stXW7WM2gIu8nvDJc1LucSdllWk8XJ5PuPndpzHIaNDqi5EgcDXdnTbu
W1jf8YlQPbFjgsEBLOle3n8OeVH8SmeBSn+oRRIG7RPY84YpwZdQ5zZxojAK
FQxmAuDljI7JQYZwv4wEzi2oMDHqx/JtpC478w0DKfdiPOD0rDhr8pOTTwdz
AWxRA+eWSp4K+kSkqdUHEcmWlwfBdPeWSxwoL1EfN9X1C6dw1vCAeDmtcB5N
sE7EsxdBs2jzArbn9E3Fvf4KnVzW/io51Pmo9/VNnQc7VVQ/Dm3wpIFVCRHx
lnPrrwUPkEEfjautc30U2Oeo9/wIdLwS+W3j69yKsG0L7ejZp3BwxDuNIlWe
nxu6g3wDaTxsT9SArDHpP6ZYZtMD8BsUl3EwlETwDQkbJVq4VyhcBOKNHxDB
km8Cw1ee5M1+1VkKMaXbWjRx88aWM6tgZlgYOqu+FIEgT0Z+xmihK6vKOvtx
kGBaXiTOaHxjVR2y0ZSKB+dknpFzOUTs9/e3au9taEGIHx5S/+8m2ZQDqxZF
CGltItGtfAgT9hDoR24s1FpgsMrPJ6+OGWxkNx4v05HnrQl0mm6c7yzGsFwj
GfCy5CcyimVC4BxB/FQmq8hG8atu2TBzvEHwovb9kOF4RgtYrNwErefQ/nH4
bT/WhZCklvQo1fp48v+eX0alH4ccl4Zay6Rdth28D0tBhGsIXs4yZXXqnKqX
O0T7WmkpOTRrK/gUjAV3uwyijFLIHulx5ymia7TtWc6GNuHwK/PERoN2OyXL
2bxz+msDza+stdC06R0q9bZBN1+gOqnNi9aHD52wWjKNGQoPCvaeUlJmt+XP
TzWNxz482ZAldEgvYW8ojivLfTO8N0JB8bvTCBFQ9C7avL+Bg3ew9HlZHoqS
cEUoKEL+wD+rFi8y4rlMpgCoPjmA1WingmTdPV51VXm4QsOUv6FOjQRCQzGo
4xCqOXTK5nd8bsOyz+I22h65skvM1Rgg39PJaNgL8lz4IqpOL/eIGx4vEcrQ
rzwLippy7MSokTkGjAd+8SGfJkdPqQ1ZYFJaxMXH2eM6anl18O/BfGDRLp/q
+FAHvrjULTP3qjvDyM05UDM8EPvJmlgncotoxjXUDNnjtFTFNEGJIZHdFApq
wwd2YesZUI8tFsMybb24SwZIbjKeK7MXMKicZJv2CI4zzAT8+p2xXxxPnVQA
RzBrRTf/uaT77Y8iRa6nQ2UDB37iNxa7QTCUenzT0i+PyV0bqeCgvauyTLOD
+xG9UPcAm/miGXfOAs2cx9NGSJwi88iW/UVjtx3WDXyXffKfSKDcN+/toN+j
zNmzZtqTBSMUEXiyyLOWmcKiUnoP5gKGcvfiRLsnUfFMAJqbKXHheyruKv6C
WWbkJctK3lkzIU+ojVGkicdDLMP22AygfB4W8M1Ijbu392nFe8xSoCv2Sz8i
VLq/3VxiXNzZ3D5/jFEl0/LmrCXxqL5VmbNBRLMmM7Rir6dmPRRK8NwtgoVC
+F+52XXdBL8RfY4fwRtX9eBpBf8HBJUKjyH32GRxioLdM1UG7ofkUplbyUm+
eieIvYTbXwMXvYLkxMhzRIbpXToy3F7pSl5phc/NVmdVw2Alm3wJ8Kgc5A47
2CESDpxLGUOeixGL3lNqFPhkyDXDWdaB9y4RLauFO7f1Xvk7Q0C8r5buRb5F
WBQvt40zwzvhBExL6qLSD4zyzyQC66e8NPxpFw/owS1mcQcjhI4vjvdqPNld
IjsRWwF1/oDP78qmaNyz/sSSawyzVBQdbXyozfh3uFSRKRFvh4LN4+MCpXO0
QMwTZTLASU3iWRHV63aJV4Uq9ToC+1G63hBzhQsbiPsFPE3C35Hf6RXLDwVC
8fkJMmrNQYgtHD6t6dtRm+In5IrAkrQ4kGrkAlB05ZJm1M/hi/hTUA6l/tXu
5MTlGNGLsl/DnJJbPDeZsTmQYmDzY6xNKF/WZkfee/ec36FB92CfOnKfZleN
sUZPqs4ckIklCD+bC1L7TBgd100yRtAk/Bn/gmNx0cSJyijOI6pY0kVie9V3
Q1IwK86kC7MrUDslYyHUQnuckfqtn+M2+StBoW/Sr/xuacWPqLYre+rNyS6Z
cSLGngKhCzmDFj60aP0CBxVz8+/DeCtyYK+URYshLpB+omlLCc2cXw0u2/2r
hAGnA7xLhN4BQg2oPZOPi4nl3ris7HFZtoHHB4Jz3DUksuvyCAqAuuak0eG0
A13Npwiqh5yDpkwt3PpKHYeqOqkdqTary6P6rUN9HX2VK6IeiqWZmq6AC6Br
JcvKqMx4tOyTud9tqkInErz9jpGpfqk3nEFKbp8qr+qkAqh2SwgUh7sS5gJB
aDnHjFbDSB1iZRa55h0L7DqPgAKWg52TM9BI3Q9+yel/pvyJC4+PkLzkMJwG
NgKnP5eCdBSGQcCjBZUiJda764mXM7WIa3d9wBTxWl6+8bBJPu+B3TqTd5s9
8A7eZ+5H3Vb3+BP8P+xiv+y5Vp9oRDFDfDIEeeDvJMXE9ivhCyODS/3AHTNP
Sf9mzAS2JMR/UaVfH4x2uZMDcOYGykoHqDhKE68MqRkxufLcLef9M29HpXGW
RJvBy5bKw2MCSc+UiD0kGij//ZtdfW+w1XaD25A/tJsEMG0lbc8TRC334aDl
9dBxr0M0gWRChHaD9EMJ3fB6x/QsZI7hgCtqWbZwD7xXSD7qP/eohvjAgcyq
8wnHil71sQcN8xAGL4QBeWvei4CJU2rCGRvtPb3Agtcs0CySYLkgvNGMEqrE
piFQqKY7M3vbWbZvN6zWfQQiaQ8IXSTwoCkFQOADry4oAJvp3v1YOWruB2pg
MLiZoF34asmvGctBnO0arlbLi/aMtBSp2PGbjKZM4ctw3SA7DChXbvaEKCz7
ZHXH/+L2ouhVNDJSCV3fxAi3jlgDc3Y4rWGBwGox5/k1sSl87STB0r1Qdxw6
Jbuy4UM6N4IF+6+lAfPuubGi3dm0VsbqPPsh/bHnQZsN/1QXwGZopOjAxDsB
8qlmRVtx5Llu1V2IhX4Id2Qg2INlYGb3fLQNRTxPZXzpF8VFC9s1iALOkUwP
TpEYT7Jkpy7eSWHNlIJEkXNWFQ+k1MgnGZPwpxSVTKc+DWXO2EFuCCm2GqT+
uTRZGyrkfx3YL1UEOUfwORK56TWOsaL18fXjPzMxA8VTJ8vt/6Cr4kh009kC
YrxcJPuHMNjpcrrFtss8TPEUQSUSU+LwHeKBX52UPfmuvt5tWOV9umDVRTom
IeU7/xfHhs8ALwXM+64535GJCQgVOsuuaP3YIvf2k0cAB2NwDVvvrcCnuRyO
GRRSXr0BLIOsmyqLIIo158lb2ddCObuC0Lfj6GJCRWssx8Sba7cI2/k2F9D2
qI+SIYRG+IYX14U4VQAGQBbNu+BfjcBdMrfte27uXzakh1TmhTjWlzMS6aD5
sLNTS7HbldSicjU0Hl+osQxQiX5F4MP3DrfinCbq7oju5Vl6W0duPQEniUZo
cVu5fsDuG4X/esgCPOl5ApTnXyrEauuC8dNaFmqU80uo0U/lO9IJSQ+7mq93
uSY2AujIRGBqE+Y2Zd6H++VMq+qgBNCcgXn/SfPf7UosDBal8wjlFZgCYyDY
9b1gpXjxP90tvIJ1oGcG4LFLJanf0X63/OxHSPz5D+XZYBnUWPPAmaHwRmIA
b3QaXWIxOPT+wzYdRjjJczfU5nEvxAJgX/V3oNmF8Wz37rry9NquMmGKd5Dj
p6Pb5Gjx7a+7eCETSE62QXcYOzoscA7ejfGpdscRqi2swnj/xmK0YZRB01bk
SUPrUnM9FIkSwVSILvGfij+r2yH0D6SARasCTDrHVflA2z1XxP/1OCbtr/CB
48+J7PpVZPzuwLbpgEhnJNISSiYrQ6AJYIiSkK67a8togH6a5tXKydvPY9IY
UV9O/uRy8PAnXTqzJ8jQAPHdoEsBQVtGrTqdB6qkRlBqX/YYzoOpxbeelQVu
POecRgG63t6rJJgYdEnaZNSxdDhF6pqlXbdn9I3ZEAh+nCweP7ejLqt+ePCA
rL0K0hShMzaMDk/XLYfc2XnQJrSSlW8kCZKP6r6bPVb6eeQ8sX+5VoImjuxU
K9H7/qg7BR6ISNmSd+z/UGK8UPSb3xOHTNw9Orw//yLAayq8fQoVR8E7OUmv
DVegZWvKddCRqGX5jY2jRgo7uEuG2SE5qG+CRHs1HNJl+6zJj2XDrmVElnPB
kBqVte1ylRbHgMUu+XKY6Ke99D69c4eLkdLPZSvAHaPljvYiUblZmHCc1zQY
RU7E+YaWyWExlJYgsYKEkRxDIO7e0X9kSWsremP/QJ60erSY2HB50c6RhG6n
wTMaOiws1K4Jqy25Ny2qPpKE0K4KARK+4ES79zlIWBH1z23BrsNdEd1bBGSv
xMEpTF7+eUY5XlT8bUzyFfUdR0p8IEt2P2MpXMzmXZYoT2nhN7+P37Tf8YAc
WULcYjE56CQiZuqxBFT2QgF3u1I3yl1EDyd2v3sAWmayIVGSZkHPSVnfan9v
i6Y/33zm+MsJwNd9ERireet6c0oWGZRkRun7M3enKDlY02pBFXSOgFizrxTN
w/QarTXr6ZRMCVQlgMNrwrjohDA+rQzRgNDAIXB3WVCxA7r7KunVUrKU5pSq
/7pSSltfvD6uYEan/N/9Ew6vgBAF1emqj5EU7zqbSObbSMnLxHGNUWt4a+8x
W3j9E3qajHJWDXFSlA7fAt00NZb+Lw1JPpnNxSQgBkgqrOM5+mr+eeuXcC3I
Np/XgBCyFI/IicyOqyOCixDLKZRGMEggL1ZksxO9HjZ4aWjGm6Vt8kd+PVCC
8XTRp9qsKmYwv/SSdFQBOIp8xOD5eikGm3dbkn9XSCx6DPPL1wm1CFIc8Osf
AhSjkXT8dKBdHLeqXLZiLx2AyDtURcwJps2oV7gJWzf2Wf72EQZCJMOtD5k7
/BkxxYJXew3GR0oXbLTI+5jQyb/+P25kARAZk5JDo7Phsj7pnxZw8qJiUvZL
3sldmnXVwQtlvwo5SnfVpaOGIDnjZQi+2JE8TqNdhaLkAtYcdt4P367kVLBp
o9Kk+1u7UvOHjKzgslefWuSMLIt6BFiHLlWOHBbZ3VNIlynIV4ENK1PPscz5
1r1W6Ofaay/Xu8aCDzIt+UTM7MdM7GtEMsQsfesc/ZlIS7qSOMJbApPlpP0b
ALJK1s+ivlUo4OvNRJGAKqGn5jF7I5ihs3FxsrTaz3MGKtaTk+RlImULbMLB
GXxdXYkC0N3PrlIR6vkh7P6wlRfy8ib83eXJpa5sAvSZCOHZON6OUc6wXLe7
T46y4EUbfPJsIbGPgViLfTp9jtnY1UBFeYYMbFF3KcHPaw2OgV1wgdJ+Hq+7
LNKoLY0pLZVYSio9ENPH3ZlWl++rrJUT4MqWYnWkrw5RxmCxb2OrXSvDpp+S
96QevrRmeeNWKfQMJJevWlVjDxM2QOo9hHzSZVs1VTVF12LRoUtkmeiPQ3He
9D4ILoF9YtEDaJFo5syGwgDeUED06ncl4CDO+Fj45spgtennqXiLbe6eULHz
bvsYy7DNI5OXY1kO1fOCs/UDAqW2TtwoRZeUsbd+hH2w0lA5f0yufRj2vwJt
+ipWAGt9y2BiH06EDOzTCSovV5nK+wmddhaX6JvbnGXemN1OOZelS9i6vL+R
qcGCj/rGEBsoxHfZaV0g137Qm3AbhAMfjiv0ZTZrWZixxfLcnggewq7/YHXQ
YC2tu7aifr3X4PTiycy6TIBP/jTUn71aNM65tAmrCkzu+V4OUZMcqOw5toV8
+HVxYfWtOpWBvZKo9XHNCZrKW4VhV/vE/eEgzy5XR+5Yj1AKp/ARlK56eu74
AuSu8JsMLR+Pd9bYkaTeVC54fGvWm0GglMQZ7kAnKYwu6ZFRlKYBxgyJDcIo
FRVUhI5xTMLb7tCJ3oegZsdIDuzbjJku5RdSnbjY3zXwSIwfxZ03fhx0o7S3
7e8aS0rtCGuUPhmxdjGgPe1e7MPgfJnsvFrW5GqFWfnjfySZbyRYBTMhgGAv
XF6IAakPMAtTDrIyLfIDuSmY0RzzO1bSqwHO0ElKA8c9/gvXbagZIm9Y0OLl
TWluWBnuIYulEqn+u8b7UHXhwTxuIjAlwjtRhY+QwzyAbFs22l0oBOdJL2V7
iyKM6UfFDIvEAbr7D8g66Oo+poTaRR0tS7pMgfPalD3IilVco6JpL2ePT4Um
2WHxl35c4HbsyUV9ga4hc7i9GQjaIe1oAv3WvealovXUE3EPPV7bFfYbknWr
eaP6DMdrokFREChEznh9kPFCDCkGXxyGGZMHtbTbQwDWLlcckAbZ3TXZxI/h
wrTKL0cwRFlav51suhDWkhZUy5JX79Gf6hYNu9GSN7uhth31z3/b+t+YGcwb
NxYwLFy3E5Gosqjm+aM/1rOtuta/hDTwfyBlu5Zu3x+wnmhVeQXNSPjP2MJ4
7LAoICAMRm+4cBH03OKX5C61do/D07tSAEU/LK1mzATDPMj3doMbd3uGY9lq
7lVCqFI95jf6VfM3h7Ld4ULriPF7X6I3v9AGtgAT9hg7rYyTIyrDGCHQ4mKg
kiT0OA380wMuzGCUR1HhGnX/OH5xuYAJA4iwNnM+BnsBpLE3uSGJ7qoZ2TBy
ppAtt2oZGFvN08a3egtGAZ0aRkMyM7FwYeCcl50B3JX5WlxBZ5i7IEEXenup
0/gMAboeQFy4iOaA3imPoyuikiRs5tnjavs5ur++C8kaRDxT2sVyy8iJhBbZ
krsYBYPO6xg1UI6MKTsIUdlhNmH6WbKXsUA7WAxbne9kwE466U1EUC0EX2l1
HEkBMbhBMZE/kuTCtmKr3XABOzMXZSHttGCkgdBMrQZqaEfJvTiPnWG1SfQy
xaFAgkpNiM7TRbbike+mgbTjElze+4UMpI16mQR7BdDlMpUp1fbSHtXBrKaH
0CyUkrAOgMelijsF+GFXqr7SVRmrfB/ZB/oDyCdkHkmUgXeTLWZXfIbwy42I
nm7SZwUg41ujRpYgJyKYyLDgtiW9I22ZwnTAhF6YmCzITd5JgzNsVgeMihDu
yRN0QJ/T+MP7GRlXCQ7isbFGDKo31/MzHjqlggl4piJMYrOMmNGAOJjicAMJ
ME9TR+P0WxHBYgxGdCCA9HRyH8JheuqbjwIQB3/gtlZrGP1FXXQ23Ax0lfwr
KJYCY1KfIa/BoT0nVC5keWmiQdfQyf1RKloBi6eRWuSF3wfFMhC1R67ZzoYi
f8k+k+4D3L1XyZw52OokXq/5QCPxw3gR9kcw628i+NwwRs9P+EIkwDBpPmDP
rrY/HQMcl7IR4N8vBbFO7hzxAOx5WEJwa18is1rc/UH+eWCYKFH2m4tKGaYQ
GUxLw8mYnNYGo1oGVl3Nv0KHfc3tHRgtYqUY3R374qvCCoLXkqQlvTS+nVqW
yDmw/htiQPehUQPhTWgm6EyxW7qYfvxi34J0yRPnLFjNDBn37OxHAg2M+5/W
Uta9EHz0dFTSS5jQRKbkbmOVci+3krYoCXa8Us5jbxDGpAUtVUeW7l5JHEIL
4ZWXnK2hY1jYfhydlKab/yVASbux7dkIJ0NdfFBlxPdMvbCK8/KAsTFZMZp8
LQfBNwl4Sn/EusqWh5x4gnEayTg3NVlTq0xDeByajNjhXxSkFZeW4d+o8kxP
6WJr2WgBoJ7/G5XzTapL+gknQ0HOHxl0o/25OAWEueLCw0p4y0LR4PCdCRH5
8aJ6VDJXlcRrVu9fIDSp6k+OZ2m+2Dah3yMyrtQId6oDcrni3hL6lLVhHkI2
OA5dtZhC0tBYKJL6HlNM0+g2DO/J6PVJemX+pzFk8utuI10mzrvLbvAVAhB3
iuqw1sQ88nkEJW/opJj2jI4+Kt+tRILroNZHhPNyoWLZlhJaGQf0hPZn0A2o
ghSHIgCKi9Gg62aaaP7548Ssb695xS66aurdhJsfLOywNwizwaY7CKK4BahN
m9AWXOdSWEE7v+OGuHAHuKCYjJmQaUUIi1ZekaoFN2KHz/7xPVDft7eB6a69
i0KAvNjiWcL6L1/vmCdJINZntpE7dqV4W60GFEPgf1zrbnMfnD9naWMFNjaG
B1Wi4vNXIt5NBOxXxX1E4t+pkIs1yq5Ohf+ciTJVfw+lyAa8H4ryoRewxsKf
+9FNdjaJhuy+8SHh8MBwdepVnCiuEr+c037JvgTG2qnjmdVKyMcxwKoYg5IL
x/d4/X5oZoywPs6WEeq6qxGGbmmvM1gM0OBinZqms+GzMvtO+Hq5Yszf9VN4
mERuYzCLErBdJ/DfAAIJKKsD9Dbwpjrj9M4Wzvp/N/GVkz7H2WjTqCi5umW4
rUru5gnA12r1vFI9RfiwMxP57ckH/5l1fLa90C/4sUoKKld9LQV85XUXOVy7
pJ5L9MqQHVWbePSKHLA8ua+oHM0xravn7qSEBH5JTnyvrnRKSMJhOsARXYAL
3n+Aazqy4b1RBS/5McmfGgZJCYS7T1iMBl0YltIk0bEVIRuHXrJnO3k5t+Hs
jNQcAJqI+raDgfImRZeVxG9G82yRXZbqbSElyiT0aRfiuCXVsBBKOpvuKuJq
UvAUPvX8cbYoUhEMG0uQL5i5a3vnYaSzINsS9EsC/wPt/+6dQ57x54L67izU
5bXPVe9eOWKe32vSNwLGXI15A06UDya0kj3trymGDfFv1oAKpz8gchVhlJbI
JOb6rGM2ITrmOyFXZk0bTIrYSBGeXVYyTz/eThfqQC4U+YlPfyOEYfU64qvv
j2yUdm38ELIDqSre0Qv3L4DUVu4euNY24JGA1boDrHmBr7+5QgNCFF22hPyK
Lv8RM+Ue/hweVQf9vd6yclZYRs4DYGiZhud1DSz/n7qSI/6RqWfDiwCBPUgS
UJ59hAE/mfLBbciTANFrHloD0zuRqswhEYqICG1WuEtvkbwFJ459XQTBix7J
F6SfSq9jBgCdou8eSgqISEs172D6AxrDB3+JR1d71j9iCZCyX3PSCw4cm8XQ
yxPK++SCjh+/Gm0QI81hUbM4A20tZju+dOhBaJP6RqoKHb2s60/6HUrquXOO
CZHbHqdFoU+1LJRot7JJMboLBvI52pZ+dGGV11hdM1LNYfbdu5FoXLkNbW7D
BVGMfVG+/whveA/nHsuH2mlQQlplEns1skxM0kyciIqcvIKm4sHFZHC6BEsF
pcuoOWsIBp6QFKWhvAABMh9d19WlGBzguX0K98+DestoWuUkiHpIQ7J49rRX
ywNT3BNl9S8tJLG2dbBPtqvDOnLatASLVIMXYFnKd5wawIKGVVMrMU5ebvJ/
2bgjbJFSz5EPet4NqQBEuImyIpdQOcdQtC3/0lageebS2FNYMqOMJWaRXZ+f
xA6/Pv8J9mPsWYW2y6Jlx6rMVX6xfRuBi0OAZeBDJzJucJvkgODubUJf2s/C
j15Jez1lO5wFt0TZ/WSx+4kUJq4ay61HuVOfB7TScwt47+mqMH252rPJIALl
PB0y9ciE1xl1uFWwsQzkDBNBWpc78RKUzTQTO8KiEnr70YuCsEuiV0qdEPCs
ILdBS1iCfimvkMgBWVq6KuyFfinWjb7sbn5atOrlW0Q+yQL3xNT3AUX0ONn+
rmdOTLJCIivNLyiG9fwOEaZyUPAsbd4YpWGQ1ee2lFiJI7Wh0/FV+7a5cDmX
SlE/opT2ujkIXxNxu9Iy/PyXUrOkFB+sZt68mKV2RwTksSt1lK2q8ff96du5
pLBWDRCMdECnQlihYMJSGqO8vBy27pUz3MAgo+LQJ9//sweKh51//5EzK3pC
TzNJN12tToKmMXef2VnWZcGpwkyHl/aw3V1oszw3HitMoHVrgpxxfzpHRtP7
TkF5lSmz772xNzMH3VH81kl6HT7wKeaRmtdsouw5v/LRD2caHLZVXEI2VRId
+CB4Eej7VH5VnYw4YhFF8Xm6Ebm0FkVE149/IhwaXkTNg6ksviTgC5Mh/4L8
uz6pl6KXHaHp1DogTJwGd5ZzHUdl8vl/iyRlhE+BLABUXWEf1FOnBk2o9u0z
qiA3oSs3YzP/QBhhAALzwjoYxoKPyzGmYOr1LnwPuaciCwH12BZ64lyja1ij
hLb+cH7gLSnwBCInWj/gxTZeByLkpKCku4paNrjhh4fjCdA51cPKCkF0nPxe
TADduemonFKqJGn/pdHenFq2oANUyuRfkbMJoonWvOHQUkufaUJ1gp+C8SaK
5miXG2GiLtzQG2b+oPgWFTv4qJgwUH4Bdkpk0zDrk2xjTh10z2ZNwRgPJy/W
ILFMnSUpDeuzwQ80Z4Siayj/OspS301ixkiz/eWYfa7Zzh/pDWiMi8Hc8y4N
v0l4IXXdevRgbuIeBr5oIu1l3PT+t1dNtqsJicXmyewllGevTlpOyAoNWLS2
cmZ3IzI5lwASnMdcjKkGfLQNiMFB4o4UHuwzRbhfAOg7jGIpifYYawvKtLmd
QOYQvKBKsJI+bZ6tiowv6q494Lowzc5UDRzWd5QMDZ5VTbIYCXpaAIvw4jcF
zVGGsDKmteRQV77yUQ2XkQeESFhZpmhcSblgcCHVgl0f6X3FRIO6rgnVoMVX
IgTE4dzR5y2w6wsLDjRS8AbxxWYYr43lKuvSbn3lcjXJFv536fhJMjuYM2mr
4OGz/imWrqcTMlLy52re5pIJaENS/6wstIXVkfholPSW10Ie5aWtvBvaGBLL
PC1ko/D4/VjT7rybeXbaPEiRECs1F7gKvYBQlrt6rKZS4aEIQjN2DXMYwSZ5
zgfje2AF6QAJq6KvzJY86TkvxRCmC87Yi6u1swIfEexq6j6JD/nfqFnq5nIE
p4Yjab/1NDGuvUa1ab8PdSELZ31/5eLgFydAk8wIKUCjWi1bhaemlySvqMw0
0Kx94z40elJ5NQwyQOM/RvtIM+wdhY44FB0NXklu7gvfdFF1OJscKImep4F1
Y4hBkuYt6Ujvho6Qe6hBzclnGxUm4LqkSrrycQRIgsjdD6+BWd2BRfPz9UAC
yc5fH9YE/g4T/t6aEwaYH1BkpaOM3S7+vkCeArYbV1QX4dAjD4OE11IFXPhd
lOKgv3RTpREmsUKU+uQF+6dKO4yOfbkbCZcCHFUA8ydCA6NoDAbcbxgADGDY
CGhtyXYQlsA1jtLN0DP8Is2jCE9cjdPb9lP9BgKEv+OKcYhv9bazuxaunfrR
FjDQZwerglnWWOJTWju5cY0+OYs3WBC4TijHcDvxAK6/HZBDevv+XJFNwnZL
hzMI6ty6RwTf85tHVCdMwWUFBRTD5Vxuz8B80XoNgP5WK0YzRhlsJOYig1np
Aw7WgdEZvksy0Y9TVDwaIFr7CgD7ohbmSQTcZb2rDB+RCL+bWkoGYWtDiqxz
+HWCZOeVuR4aTuOvYtKoouBbDTJVVKhozxOspjtK89/Z6MlIYBQLBKyJPtxI
8RkmR/UAdSxEsneMP0x+G95WfoXrWdR4iFMvNuWkjFGYt2Azvh93dUKrVBSB
7Bk8z5X/nJXxXnV8xG4NHL5y1iUHfSKKDw2/64WdjLS9MrhZyClJ+f/90jDZ
PmlDAk3e0T3yIOa7S5EZZRcab/wWOogjLiJJUbS8Jf86pkuVlS91xycy4PCO
wohKVFA8Sk7ab93uml+6hPvf5jKhdjxBxX/1LuMFrpWQS37+wtQk0Co290lM
ZlCn/FGVHwIPL8WbygQQOvUA1i6qHN2lcECbDpIEkW3bCDHPfoNGPY4k9JLR
0lmmyOTI1CvhbdFyoWxBNfv0shZMdgvvAsEJxoqWf2gvjH3TJ/7OnrmOBsNA
N1N2bDK45BIN4CHapvm5DYVdtmrxyeZjD01FKWOBPvDaV2A6ds+H7iUnQxjt
tglQcqJiwg1dgyblCCv5uuPIODIekTyBmLY1Z4Vu7aoNkI/+dLvlAdgP9TNj
5wS7eOVS+Ml9eNmeXg9jtwRC36Qjpda6mi3cUAYI0hVbDna2FgrrKtizqsoY
kwje1Tlk+wcXC0YJnUMLPS2Iev0X3msuk+8PnH5CXA3AtJQlMoE/38YLgL6U
DzGMjt+hFQNNIWv06OhPIwNb0zJ2Yy7jXJyX36YKExKiHaYHNo1SouyGm9SV
zP5WDmH3Fft4nJa+uNK920icVA8oSDxirYN7IO6rTzUFtm3jrXfb2AZbUh7O
icxqOvBswM/TWE7V7cuFHlQMWRT5cy54EGEIwTaHmBCTqtZ1HYuBVowtCKbo
hTdD6pxUbLGM8BG9dG+UrPIBTEMSRI/Xh+3FZWBH9gt5+oj/+ZP9dIbUR/qZ
eq8mbWq6p7E0xEbitRl0H0/xnuwPd164AfgTQFKvvykKwTDLuItm2Hhg2wng
8MOHC4gp+xO/+M9osYse6ihBkBQCXH1dLD5NN6l6xyzXybCWoprHFR/8zg54
8U70jCvCwT6bCKBL9zMlCYxV/s6np2+iDFp5ntbWCi0sdMHzrM4fB3SM2Ra7
9yDUb32+96I3++3/P+gm4u56OQNmnb+OONBs8M2t9sIqEPp9o8eIFA2UAaAS
T8SrR5/S/pqMuCdQk8QbiMYrKhlpBnXNeC02kpYdhH8AVISVH5FKZ4m+XeUa
oRCAKCbHbxr0IITBkCDnHFPyWiyPuTYJz8fmOzO9FEbhrejzrXPLdxqNbuI3
fmi3UlpsspYQ7lcrCpktJAjuiYd05BJYKqy3WU0IXmYR/OxKa5w1x+IKRcGV
YO65N4IQNCyjrs6zqgIqZo4P0xmQjp/CrieG5G8XqYYAxUKse69vu9knLymY
hM3Qcx/FZNsiNAnoAdXzmAJww74/Sdh9o6Q4Q2htXpucyORM9e4/8npM9wjo
vH9tAYGnchM+4ySyxXjzzT/RW9P2ocrbTo2L+XIZD0Nmj2YQ6Sj0UjYdUjAO
zMAO3q2SPSRjUFd6mnaRaiFG71u04t5ub7giNfd1mjeFf229PmbXuu7tpv0x
R3UcZpTIikTpwRSHV0Ct2PKQs876avrXBHLfNxeMvK5d1XLyhCLKF530M+Bq
91jULNMAP9e+LvIo9NtRgjpdJYqg9HoBzZPWA3RD/Qh+kyJCIsZbhsMA2GW2
SFBkUewb8f1MqzaM81oXw99K5EsFgDIlzGgAaxlwcyqeoA7Lt8vXe81YiVyd
b4X9J+u8SwQk0o+7Fr4ggVmO/I1RC51YMPpM+3sGuoPdRItaCZnbwlTWQqtF
ZMQoCPBvsfzsv2wX51OS5cUXtQYOFJntpbAeFlSLwCBAcnezj5XaX4x/Z1LG
BA6Z0a8lzrPzmmTElGysaUOW9gPwij6nP3dvpAwUKjmJ72cMhtYPX9EJwdLe
+JxAD7ay9b9MGtoV0O683rvCHcuHp+tAEInIbasiBEdBxtRedzIHOniQB1op
/BuVaoYzZ1aPK9CSyUrfPQHWPhqKJyGhOM/hppAPd9zlN6LQLuEYZNwei08W
A9Ek9AXNeBGkVy91QirbYtQeTS1An64ddt1CMJTbX6wej9QIwTN1FGNkcPvJ
VaVlgAGkX1IChmIUxffVEED7BY1cOLl4c//AAW4g75J85nO+KVKm8xYKkFiC
/cvTcSlr9a/+fxzb1D0vStwvxAH5vvYEN3cweTdH4YBITx5EnYwf0vXgeMCh
1D1FG/30Xq1iMtYe+ubxfwz2E5G+n/Je5M5CkWBJUcUFHqjqW5lnJzNqfp8F
N4+UXI3TZ09KZLPW2ayFIJ7t5KNf/z2biiNiqdFjVvfqDNcf7aGsSoBq+yhX
jZBARIu79fOhcMRwWQIofBFUnbo50LVANF6z+J9/DBK9RsvghCeX9rah50jL
nMpPTBpaS/B1r4ECGW+VjNUp7nLioGfdQPaT0DTKUYihUZhklO7ZwHIzj28C
GFnjV+/p/yUJHCHbuPuVFhpbJrMpHJRn7iZPM8qpf6opFVyCQN+H/UqqEspv
S8hM0TjqNBYyi4pDb4lt68M3ttArolEzepp4522lz/eHdGQ8y87i8KjLCfRu
0JC2b/C34XRdQ3VIMZiV44jSIhXdLBuFIMI4WImdVTZD+2ax7Evw/VyoZypK
4V/joI2xrYmNcBHdAUQxPxfZJZdkV7Fd+AopqOt1lI88caDE/J/yfSTqtWWk
ZGCaI2JuF+K+aoz0bK4O7U/hrDRufXzGmj+/7uXd/oGdEpb1DnirLR0dWd9y
i6rvwxagH5frpSG9WFOFECrG1SigPleYl5P/ljTpIhCSPTkE8sR7AU+8QJn/
firDTOBEUpHW78aJJpAnj/kRlnRzkPeEzsBl8tWd08r3CIzN2MxHgBV6pKCm
snmTjxOLgrsVxZijsJF8bjYOi42z8B//sAKUC+KlDs0ZYCpx5h740H1r/at8
VKFUW9qUenZceahx0aKv9tXbq4WWJae4m1FxsOHDv0Nzwv1DkFpn+Dx5sOnS
wBB5Y/2j0Hz9WQYmbWqRRjlw6eHWfMEsZQlWfSux2QzmiW2SArvaqd/gehq5
/iDH6rovXcfMGJWasZX79L+aA89ZWnjNFmuXsic7uFgyFQslFeWMNmtL6QKP
u+gDinprrdReUYgM66Z47VPEUkX+Rmo/WaAVOpJZc/veWioSux+bFXzL22jm
/W1NXOEp8NjWLTU7uWwel4YK+XkVlxHEwda5ICuxn4Ej3EtW/uqeJ3/K0rZX
FO7sH4H+hvuegTgRx+mHz36/OqHmaD0+xOIADLHDGaygpmnH+vjdDp30zshU
+GWAuVHD/ngz0++7KhiGj/aPKbh1rxKHEHALC8QHulQS6pg/hmkcAu2wsS5N
NWtjr3uZdU2hfkMsbU2V+rf3J0cQbP83TG9mEDYAoq88fBcXpQUzMC56lXkx
3PJ+NWyVg/MI2H4CqNwNZzCbg1Rj/kuTrxDjR+8a7O8rZSnv/f9bRJDsz7ZC
TaNDtrOOpjpdN/gvTHZy1uR5FJrtuVVufRaLKHY3dJ4YWmdSCt+qUQTKFseE
4t7RwYHa7X7hauyBBRNCf0hW4FOlyCUIaEW/N2+S2ZdRgtfmg1ojncq5poGg
9Cb5UCVJKCMUj/e8VXUe5mA45w249Hc3p1jYfS6Tw/jQPSoVS40QztYr7HCQ
buqTvwzwZEtB3Ofkbp7uAUQxWIGWjAViMwZ1F+7OuOnNy9yu/84erVUu35gZ
a2/vQqjp1mWCcC6qINGW/mZi+kXqkEkozhUstLRyx3y080ZxNfVMP/AykLnL
n/9K5IbdjW0a6V9iFLoHW0JEj8XPT43Y6qRtmM1kiJcn/QSRVSSH3q9vokif
2NWd+Bprmyd9yAB2a7BcxczXzBXd73QCGEAM1aI1us3iDB2eKe9/bRu0nI45
Gf+xBGm/W5sHY692XGce92Cvzls/MREgT1irblRjRH0e1V0F+U3XHAX9mqnc
eoroGUqLaRt3rD2F7H6OEemQNH4W/s0YSgICPTpw3kPn3rN3MD1WPJ/zBy5p
H3sFfAUhZ835TzTBcVHlds+T/Q/KHPX7fXIOwXmSDN3QV33RQ5Q41bqHctEI
+sko/lWUWP8nEAnjH6qKlj7nVQLKJvwaB8lm7vsxwFGKz78rI5eUxPmSd2Fg
YWET5/txAOLCYiEqovRF42uxGwxGnIxJIi736ttCkPQCkI4w9nYdcFG50ebn
XzHeKtJNpRakst29IOldWT9E5QGIMVQ9ZG8LpYvoTnVgV+9on+8rj1vR3v19
ZFI25GJBRn5bSeUJ3fUSqF5KCIGp2CXkgXcbDSVuxGBTnCfL5eshGOjyMet5
IZFrHsL4Oxw28QR+i9xzFlFMWa7CTy7dN45NtmPp2hPCpI4YXn5pjJIIAiae
ftk4P5k27Shhh4D6bcJ9vNtr5xaCr3nFq3LVROJCtE6HvhOlNFjTTfCQG2QD
5FSFIfqtV2j67ldCQFLBsbRbEuZGBHCtJkvbuwIhYRAH3/MXHSzo7BImvxHQ
UHdNqhAhzvd7bWoMYHDLpyjoqe3Kvi4B662NH0wb/Vk1FIJdoTjg3UjWky7Q
HGInuS8Be1JQntOPTeGMkTrfZ1TrqSGf+sVe/uWSCkysNXIAS62PBev2K01f
shwNZMtFXCxriytv13u7HctBEVDsrodVrYwos+TvFegpYSxq4Vv5mjROEvGr
C94xcScbfjrSklSYGUdxTUyjFq3OWzbgfPpMWPEDmC/7jUT075E8qfFTfWje
vMUCo+Tux1QCzZdLkh4+zRFZ2qHAAHt+0u5iwplfb9OZBklxDKOJPmCXU0S1
szWe5ze5uTXzNKA2XLhfUziodajt38R57lD8aTI8EyH+eF3S8v9y+t8nG8Oa
ytFPIGbtNyi714DM2IA0QRJX84Ihkknz+OqnbaFtnvyLp3M+fSK8VT5cUtQe
ApYSJ+599/kods86d3n/6PzUi73C8aYuBoDj2EZMYjeeiPWN1s/KeEwiRBIN
cgRTdczoQgiz+dlZxcbHqWCZuOEPIn+zcUVNksniMBR2Ya6n3erJzc831R6J
XAgSuEINQYqdxEww3FNkKyyyFRgJVrap/PLbsT3H+rCrpiAnPqCl3sHQrh4K
4DTy4SLc9i6K5NjNd6Lr1sz02YYU/oR7iBhSoPUi9nbuhDakEWWxehFaIn8Q
ry4u1U8s6j6mqUUwIX3dOdxT3LBv5T2pNAbnRWkXH2OcQO/r0d090dV4Anmb
6vY4XEMxCpEwbjb8vQE2ydJ09CpHXqSPbRu9LdOCJGbizv+plxoIXkcqfwrP
5oNnXy4WqcFnhfzhX+ea1QDjFKGv4gWBYg23xbT9ocaAPLtE6mPXbbIU4pAM
P353ckrRLRt6c2icpXc1JxKjdi8DdQ8VYWTRy+d+Pch7GrFQgS5akf3/QDUY
iUqYAPU/knXnDKjhEdr96SQedINQ8I42FaV/oRCdW2intf9IVj5iKja9Kr/j
lfs1QhA0gZkjHUcGWMAk6LSe/BYYcEyS+2q7AKgsZ4wnrM8DCqBfuCQ1Y5cH
3f98SmKATbqAKS2S/YnMiUbvWVlen/6hp1phbQbMssCKFFNe5vQKXbbLUO2c
o+uN6a7GpcCHYS0GXF1v/lokz5ANrYslVbiX2cW4XfAHGvW5F4evhKzu8sYj
BHRBPbKkyCfvcmp8N7Bg+KpmLEEcv4MroZjRcTPWkVrlv8eaSXI+x1cnhooH
rxxX0B0NBOACDWXVsgtF8gA2PS/HlVI6WAFOjX3vw/cS3wrBA19CCd4S258j
5PoTLtn/nSMnNZ6ZjSfVaQi0FXqGPfY8DJg4rw6+8oL1hiJ9Uzne/viq/8LP
xtmAZfqsPUYZSwku3cj3g1tMbUieuWKCQ+9ttpozdXnaq6N+jsj2E4l88f+g
+SKJeOcBkpecc/wAQqtc3TZWjj+Sf1mMkSFyHRqffefPAAQx6+hVEpEmsYCH
+2yqSgds90xzZXDLVMJPJoKPNutuW2O/xJkEcqfYxQgUV50xgT+GTEcYF8uf
ydnQizKAIxkL8Dhc71pd07/Gr/nttae0reffMk1DqMQC7FMnuRwynVHcxNQG
+JG+t+k/Dc0trGEv5ZiNbzlIviLeZDuL1Nw1zqEqPi2b70RRP92dxsxwlrKA
mgV1M7dlRRnsgXno0lNJGfI+uGdf3JN4bPcCxglflDx22gMDqidwAofA/Wls
7cpbqt6Z1WWUBWCWpaPRF6p1JdwApO55uIIUxOB4BNXCUz0TMWVeYqKuR2z1
NL90Fj99uvijPFu9Bxkz5Eyi322ew0MDakbZSM52TToNRCjJ04g0ln9LzsdY
aflTM2mC15f26/VJFpilKIerm4unhD8y0LFDQ+T+/DffunfdDXLWjCa+W+j3
MC1RVnqcHcjAMttmpOzLlIQVKKM9btQFmp9zZav5Q/hm76NwTMHCfl1D++XV
hbbq+AOxcYGl1kkgBiPjzi6XqknqvJfBpLOZwybTRHIxiWNt3cWRDDO4twVK
1HPaPVop/zEjQcptEQivBpJr++hqzsaozH+jtFFwFDVwrH1v5UXB/M+/qbEd
qXsgwSSG7EJ/LDGjC1lI0mRe4KF2Ycqx6wdJwn9ssnffNWjvXC+eYA09MANu
SQz11yLBKjcJwgvonsOB9YhgTFBQplb1TDTCVXFkyn4hDcEWugkt71L78DSc
TfNl4amRoExJ5yLmjzPxMavFqiz8YzfNfDe0rQVfohhd5t0q9ur0ICHPFvF9
aw3ZlUqibkon5IXxqHgkZUgEn5M5AKCFANtm/HqUGMFeCFZIjmR0SmB0MBy8
HUqx3Kr0/NRkR0es5mlAnbvKavVozAq+4F3eOubkEXBWq4/ssx2lQuey44A8
X0x375adw8+Z8+KdHQVFOLNGyl+yq5jeUdQbVrt0GaJxwYgtsIf1m1v5+wqs
Jo8GKREVxhdIGWeDxX0WXHnXj8vAEfy7x00D+Y3x+c5z8xvxtaZ03luzueY1
SC2HdFaY9QZQ0x4W02d1SZkwKePpNy94p/IxMysCtVjhU5+FgObBhj8oPDae
Zv7vCkBgWr0ArxWejOtG5ba3I/Y1WBmJW4aA+AQiiEKHekhc9XvRAl826IoY
rqwZLq6iCUZmUVYKwYJy0bTe3SFLX/NkbHroKRpF9UIm2dxfsonaYNrtn79S
3WjFjDExAM8YF2nyPMwTc2/sdsReXFKABmqstWMgFH8EdGn9+i7mbDm9wO/Z
keUvjbCbZQTF2amIDyP7+Pa0qCAez7Sx8ZSil4D9WSxci4++CS83JpX4ufMb
aE2uV+4oGStQ7jKBLhcl5AHqXfvGolseiH78HtIilzpsXmau3ctOagw12jA1
1wUfJSYRf6c1C2khg8JwR05xcAwQuk3hnPwDRKmnP2nokjmtdSkOfcRaLyHf
q5syAinmjrQvCK/E3d+FQkrcdWuAdB6MJ7xOlF2V1X8+xnE97LLDz2jyk+48
8jhOUvtWt5qsJfG/lW5ywpqgJokC2IO/XFluOLPtMo4Y0FFUyZE1z5V/mKDO
THdDR9J56VqTKTdmn/v6jlZ+1imFggE9Rir9Jbk0x1n15YonLkRu+QI4fyiI
uJWKlrKfDInCMASf2GRTj5fxrXV7U5HkVj2xHMLkXXPyJTS+7x4HwWeqViCB
RkHCxdc6jB3d7COsmnbi2d/yvtufEuZryjrMJnxQucU8F1N4MJi74DLKg0Ku
OsxbkVZz6QAGh9zIvviA+GFhGtLF2xfHNiPYKCSfQOrEbWxOZ1OJOWhKAjPq
ln7XOC2/tEI/hcLFk4fnRcKwH2WY1XfcRy6hMo/02rV9Iwd28gjrK1MVn7et
p4OMBZrbBfa+L7+OdUwLIE3i67It3pWPrM4bSjW0MEF0Z9vPeS+8eDmjeW/s
0qyJBIBptgm+LFGtIBvaa+GKH6f15gL6LxorNyIaaaAhSJz2HvwFOzzbKYUv
Pd+wGx6WSqIc6VOptIUZm0cOrNRc44NX7m7Uj4VIsoi6WbZQDSVPhhshO4XT
EFf86GzdrLYbx4CfYyADuikixooOQdrZ5u+es+IgbGC5MiUSsLjsBGI2CLH+
RhRw0XfahUn6NA2Du+2CXa3yD1h5OriSyXXH4ndg9G0dUuf9EIwt8NxhO/Qu
cjcgBlQtV0H5xeogcMxJMAJxluiZbudE1QWokBkhrQv5jTZQfqmbilORrELU
81izhMuuKhR9wNrKYirNb4sZ6vbjl5+gc9paaP2vCrLYpFLAUQI9OLf8HZ5v
pfj/B1e8K3IAG1+tsoxzrkYIxLvMK+jaOZNvLtJz6TMjpY1TFFNTgwRlz/M8
wVYMDcpm9JdbxixNERX7o/2ZHENAw+s2nvEefO+D5DpYKfBLC8G6NMAzaObE
kaMrTvZVCcuiNpJleYuY3GtX9uMmkJPKrrpSBKq3yPq3TODucm3nhQOGk9v3
ED2E5BDzV0Ag/RNaY1ZB0W7pstzK3YV/Hpkithb1bEE84bKJZs5uGU8ds450
jSpmNIVyvGgVyhDy0W2bcCWZxOX7zFE1gl37l91i3f6V8OIPAyl2Nnl4JcKm
npcwunZz32i3lQdPjc/Td+RsNY8frAv6GNM0sPghxiioNTbivyUoKW4FjEkL
VwJjoiNhPkEDtjeFa5pZ1YmmV7cIDsh7QkusH2oXNicDyIV5EQ5vg/Sz9rkF
xWlNRj4BQpak7ASXY6LDUO3pWP7rfzM4lXeOJJbvfOzpt48kHyFYhWqPn5ra
RKXguf4oqjIvpYDdue2sE+iAoVp3ApGdtp2QkB4F8+a7tdkInTJn0yZtVIau
Zd6Kw95iiosWMoI6W30oqqbnTV25tufKb+V6p8KLga671STq4TZzjL5Mw2M1
Rb7H7HQL4TPnI6pT28wpyGzd4dcdV/zbqklY+KUhrtltGwyPX/nvy89lN0FG
xbsydR+bD9HMOzB2Rj1Smx6BtNnQ9nhEJVaAijym51waMwlwnjTkLPciKw7y
DP5E4bUeXwqKLmpZZFhlvbxrw2P10I/v1XrqPivMNVrSpkJBsk8TgBf+3uAQ
P1mwgbYUFJNayHehEX1Zi/M6qI3ni38AlyonXxB0UMw1PM6AxRwRuBp7pvKU
rwTD0EyCflg1uYYMlTXPBxTa4DIBf+77+yMf9FynmpwRw717s4wm5rcW3N6K
sHNOb7xAKCBZt6tj5K2h5ivibeKdr9uXz/ZegGSpYrB0zibfubuDitVC7tJZ
FAmzy7pUlmOljfuzGaKbjYvH+db7UtwhYUqmF+T3LpU8nzkjPvf6Ba9fIyFA
a1TZYjHwrdGphVGHRDeVmMFBvg7Sb9SxBT7wCqK64ZZrNRPnfiOHRojhezyA
An8qyb/w0zhMk8OO6bDen5Eavf+0uyP0CE9d/BfD/kdfTRqzA89eZIz9NrIy
cc0MMR0ixU6MTAaDdVHf8trTKQyQUOVfj+vJ+FUAOTdr0vuIJNE/HH1u1RLD
anr4AWSfS++rF0RmV/sEhb4znFpJ/3Au24sW/gcGR2H3XUsfaeyxidiy+6VZ
o0tFI2hA6Rd0TtJsBKuAzcbPkh7wIGfw8WO1D+tmOe4Xejghyn/HNy/HS3d+
nBfSj/TI/brCyD4V3NKKwsCLRryQU8YDUF5cD8IBMn2/TBu3QiDKZ+SLPOVj
uNS19K6fWwmCCIa/Z6BzxhbBshDTc7Svb1sF3unvpa5PYTRAN0ziCLwCDf2Y
MSEz+chy6Nb1chD7qSH/laXmB36I2diXobBoleu48nODvYtb4yKMcIRAv+cC
VbXJTQRnkMfo3w0m4RkZ1o9fPvCWMEv/480NP/kIEAqbkIuUBdx1UVKJ0xOB
diZHKAHdc5RbzXOijHgob8xhXuhiByr3ZWIvnVMf0ZLe/qpwdPQBUgDf45fJ
KtbuUwV0MmjGRZCOQP9TbPIPA9jF7fLqBdVYZ6xYFaNSSFlxOznENjei+Kc/
Yaq5Pvy9al8mwVXRo4oDiVyiS/7vDbBG9VW2vYwaUp2D/TXSIK93+Rzv8mY0
kFn22jj61tc36OJiHXeC6tJTVwZ1aJBo3DB0YLs6XVJc1I2yIkX8VbqTb5vG
7RASXR/1i5iwEQJnDkLJ1JHYt2CqfSnHdG9Cjos9j6lRPiXrqAekbd2w4hP8
c3s+8H/T6XiE0ps5JBWSknfo8IFkNmgBvfuU6qnw2hmWK4WvN0GiOPm+0+KY
0cKefmPm0UI2tjQNhvKF54W6NVM+JXEqhNqGvI3hPI4aBl30UxtSihERhbI7
o+B2aIsz//tNwjSvw2urPZoyZzlssQNhgYqlu+xO3rAYilDjeyzzuXjtGYs1
ZxQIgMLNHYL+qD8FECZ/wu1Z+lUkZX7iPrEQ4qj+sCu+DcCP2uO1AISsSGNv
7dCiprmMBzHMRl9fY4tyY5jjTmC6uOwdOXp7VuW5gHMbTzL9HMMFx3halHJ5
caAHZIACSaN+eQDSjXTvMeS8wMBMLhs9ai+dNDdP2cDvYqHMUCH7zHp4mKmT
Ln8BC9DC1Sdph9lxiEZyUXW/bNeKL6N9tycoWNz5e8j5Bjxusktd9kar//Lp
EWXcuozf+N/3GzXWrLtOy/5qyIMycpTpYcO+mBbJNGdBjWQ/JlDE8Fj4hfEw
hoqNTwm8nf47IH64i93vlUmt9lArtC8R7EJLU6smHDMaVTIG5yTrzzU9OrB7
qpKawL9RN12jGoa7qKPhpmHwVC+s8LwKmqULrPmpozmzvNsdziNmq75XbTpC
C0Vpt6HTwDL74cfwQkY4T/1KfgCoAm6Z64nQjO1dboNLk053whOfPSyvWFAU
qfVX2klq/9g6UL/TPRuU7TBnNge3KfidAKKtNy+3YSKCgrn0SNOo1nSV1ooR
60K0e1yNCcGQJZKAXaJed8povTfdgUZKFgUlPmihkmkYbABiFQyo0olRtS9R
4sjGcbvtoU2ZaNocoNOXZbGl8FnwsT8JihEPycJ9ncwMTL+g5XZyoCLIkLXz
ZFms2s2GzfoLO4Zvd4JV/rIYjE8m1ZZ1uWTMJNQA2M1iLQPAsl42IOTI0TY+
m4XheUyLFVcIkbnbWKFLwFpXEbCEQr0kyxlIdYlVCrn4FY2FgwdtL6rJY5B0
WjnzSTHzr8jDrk9JM37h43wZ8xWt+4UweKg0rDMjhqMBqQUvg/Di4U3PJNiz
87BZaohK7YFWc2Ut1z1Q9oDiLiYixwEXENlRctHepUdFD5s//8fDpahg/Hyg
EG1p/wyWdaxtl6hffb27pfM7BKSW1/PDKE5uqNc98eWPrDNZY+XLidLLU9in
1lPkqR9uC8Bk+xFJ6y5ix3a19zQeLI1rfpm4r489GkkBITTgz5U63TVrOwzp
d+sLB3D+mSkAqaiqVmoV9jHiQPnXRQRfvH9HwWA7xJMo54u8MVFbg2QVTGCe
tn4+z6cJNHy/EgT97/AB+WjPSIKjKADRTqJ+0Vixvy3SGq9aslDpx0jnaLVK
82IG8kVzRySju/H2Fv9Weu11i3njIfrWzatc+f75SRVRJhKYatAJ5H9oWI3J
Chu+LyK67OHIidXQ+o4f8rBLLUG3JBJyfIvBxKqVi5CSWHKECTXfpGeZjE0z
wCS+JeASyI1FF3O+lekLKlmVP1q0yu8ybyahwQy5i1oOzZ8n+FSQzGeGMEHH
fUEyIRsbagAToiZ7OCKLQWX9H4kOSzd5kNJGMwLFjmmPmg+GDpUHywdZxGDj
AafI3x4FWDplTBtIebWVFsPPYYfLv4hziWTWDLGrNve8eEqXL5YwZh7kHG/3
H2yosuLe/wA0j0eJIEl2r20LZDWEhTWZejimqmen3vTaAKdEc4Ratp33/Hnn
/gMVAyAxvd1qjWGAipUHcZ7WIKeWoYlTeckoxWl0X2Xspn8aNodVOPr3qNW1
zxTND+ssxnVlopeVZCWpb/uskB7DfkQ5w0apONrrQEAbqZuv3kb2lDzHYST0
BLISrAIXBy/ydE0znA9xypU8VgAjHl65XsVwT1V/wv6ldxOwLNW/1wFA/4fU
XE6zYtrg2HnkM56BmNntPfY1KoD9hSR3HjoFzX7+W+uEZd0j1X6C/EJL0wZR
LkwQ1DS8EYWWaSJAek1ftm6HmmWYYq76TfHvZ6o1yj6K/++cpINfpGCjnxeV
vnQ6H/eSnviRrZuBZ9WHrNrRZ2d+bQIezsGAdrEY9FLShr9Nvieo79Sp2mLO
+obrjGPY40Pr8GrhCn1tq0p48j4IjfCaE5lNbuwq3VK2Yu5qkhXQiS0aRm4+
Z8z1Uj0OsjckGjYdtOZxI8wau8QJXdiseHK3RC8sPMJ85HxBFkOCNfJD6zsh
zaGNwOep/Y3+owNGbUR1p0HjF/bgilrlG4szBPtikF/YJSkD2M8lgZXA+N9b
FhdEp9+HlAjB0DZK268nHSIVjvY0Ol0oJH9z99+zBeVGyvI84EzyhZsgPO/x
OAwA0TZppoPmc7WuiKz3X3hAzXu2fFICYffxcroAGxEcWsViiDF82ljCwH3G
EyIJJtiVn571xl/kmtYG1s0Tr7IyoIMrUpx0V2Dr8TacMvzQt2ltqVM7gY9c
xRTC6SngPFCDXf0eyhV0deO3sumyoABLFXKJpNmoJcAVCegbWF1BbtGiv/nl
g8W8tN6IsLnq+OUHXs2uCMErZvFpeXey4wNIIWvDPEBlKpxfINhgtI2ybAFg
TpX+t4wY9pRlB17FPHHsW0xQNww3f63hgV6HPYtHBBATr/clzpTJz4rxgD4z
yVUTu1qcAe7k0GQZOjghQtzd+9A8sGip5mBNV/a5MWu+nocREAVceRm0szIr
Cz7p1e1RkC2198JPWFroF3X6LbA/4M/DpJTUwKVzft0Yd1Qu4d8BbxQhv9XD
QqrPOSMnZm6+m4Hg2rtQnILKkzUtN2KJp4F6OCmCc+YuBcquRzdINS6hNp2M
iGR8HjG78UxBnoiFDD9WCFlpkgfZDa7OMIE8U3p9ejlPP+2dKdPfzGf35sQB
O2rqRPoHIk76NONZkcBQwoxbTLEco61eY9T9obA9uhKIdPSJtGSDYtQxiQIL
WEpS0rol58FOpUFblMFwmSVz4JZXw+he8W4/RUIEwV7qlxOG4PCTrKiDT2Wn
XooNA3Ul1+gsSXzaCOW2ivuedQNSFFxf9RLkMzFTbIfeaCvQJgl/GVFmTVT/
9qDIKf3x1RLSd4C99olxl+pKIkar3osaGSBj6Bc8Lvu60SIX74P4z28PTNEB
oMGJ8iEzjw+ZFDLd5ndp1pFw3+GWDMLknFiP+kpg7yHGRbD1SVx0k+TgfoEK
BrUEQdFcrvtH2FoeOmys32mCIZbcg4ePvDW+e6RWC04vVBLRcUR+OM2kvXHE
AjtKYiWrWbCzXB0dxnJWCAam7GdNpAdAT4SafpkabFHVByllK2SHYZqvz/0m
Toh8mxmya1y4P5PujCwXYx7Bct7D4S1/y2ecO7eA5DrqdwoiIKwaGx/RotFQ
JY4NmvnICSD8ziEgX5zLFLXh8l+SuFzbpoHFe/h6FjSc9r4jGZ+6jRPN5v3k
kEsNrdnoa+K+qKDCgVznBhRXIsCQ7IU731IWuFqpjeZ6zXRXMQq5aX5aPTRZ
5kNQq3ECwk2wpUPlq5XII8HppJOJ+mBqqAxNyXqQK1/oFYbdmTa4kjsP4w55
cDeVddBzl7YkEUlB1aQZiV0TEmIeSrNtN8E2egdgOFX9rhJ4Q0zDsFHaVO/3
3ebu2TvgA3WQyapfAyAon4xl2b1V5fVjpyhBRiNmm4Qrij+ZpQLviKPJ47ia
KUUW/oY5uDFIw0/9Lzrrq1xnbc4zytbVFGl8OgmZC6XkbvjikJ6bQXCZrs/2
iJyichF4zbJ+mV2mMe5GtUeFwMlMtS0BdOkekrkfCfJxpSfni6Ka6cLTLctb
k+9Pzwu1hQkgumtTq9Wkz/UFHO3jPBZGcyElREh/vdtasQD2ULygH0f83k/o
WvD2olnoEc6KOqW9Pdd6x+DJRQ9A76bsbvN5SW1i4PNwfX6xEO4e9HOs5fZB
o5dhFwCazc9U/sk6Hh4TcQkHUObKV0vyV+9pRO3jPVV3tkkK7yBt7eXppJaA
sdolnAcM4YBB1HnwPpqQWWx8sucbjg9EDH01yrHiE7CSAULTjuT2zmf9Oukm
0vhJb+3G/N5PekulerIuXkf5P17gozYTNPvvvsLS0Qe2ne1EQt53PbNEsTYy
AaQ7U+VCsu9d3oKA7ALiuH1z8KO4+Ex3LVUPgJQHQ0aRZuwtd+crI0Z4GAcg
WnG9F5ItyWh1Fr/7Q2iRwwA9gAI+Iy11ZiFAe4Z6R34H92L6Qwgs92D+VnrD
B0vZXPzZ5N9f8s3xV1j5nnycQsSHuuYSObN7dzP0/WHK2+lqELoRzmTR68Tm
Fba9Wx5CJTzD5EkzvW5lJcSUl+sVECyDovckjNwdLBnqTyhHEO4ltFndTvUC
hFDGk7w//QT1UYmoIV9aOUszgMSBXLSM131vv+SET/AOpyOMuPmrwhZ1Q3a9
uqDpkf++1Ow773sTjo25IEdKbHjT2O0+6AotmQMRoE8OYkhHi8To4xLWOKbQ
lwsCIU2yNygj8VphQ5wPa11YtGZHduNzFuiZJ8JhNgCtwz7nFWh+nsfZdh0v
eanr+6LYFpaEO3YVrSKZP1ekQh4UcfJAlM+xFJOG+cd46r/EmMojEL6CJxqI
CSoKdHSRitWPXeaTGyk9B5STLZ920r1VsBdpu0ylsOVrZo4fCD4nATffApAt
scMOfj44bTxq/AfEVCw34g1IHl+3Vu+zGX/Q6g60Gturn4Ml/TEmF89SHvtu
QopAFLOCkjwTOEDuKfIZWBEOWwC4A5loNXLE+bUzanuy9mjUbFM6BbA7c0YB
Ca29m0pQ5VUBLsa8lgiB/9T+dRc1mAp7jio8ygUzHpPfjaKl08cq2ooSIkpv
swDkyKbpZi+u1NS2HLBzHwm0Bkjj5/44j/JKni/oyIH1IHXEL4klXRSjtjCW
78Dib/YBYGyuyBMqmLZnLGTq4WvVya9qZhqxt/0zTdBFlRCtJPTOWmRN5mTv
F/+0F7GgEg6W4vrhH4zGiv0vjldNK8El21BOD+VjxxJJDvKi0e5+Ph5doZx1
17d/nSTYBDakHiTfPDeyupQ5LpStc5FmzlAPzFL4fzd27/CSdPRZIGxkbJt7
Mv/x6GJcNXqsVHZfARgvuvsxRl+fUgqXZj43F/AlkU9QmwWoDDLZrwP7c8Vk
f0w7kOLRg4oMm9xnD+8QEotYCqMrGbNzxjlPI6Q+Xgw25ha80zLKdCw8UQZ6
H4FqiJtpWB0JMkrgU5YQfnPYqChN5j89WPGYirU7xKPiMctbSNan8i5lE7Zm
+xR4o8UpesRkMoSdRGFV+lsjZqaOOWXrbIvToNx8taPyVoodbvXKW6RZAHUr
UqItPBhBntdhieiDVwPuODc5LA+rDP56rXrpXPkpGc7qsVa1fsJAhdTWLHZl
4gwpY0MRdjHayQlHC32SPSJNf2mCWo2viJ9tz5ZqqI5ts6T/yq62g0jCjDoM
Jr0QbCLIO5tY6EEajYN6MO0EmyVFhNBHLZRg1Vs9bXytO4/tZiVwJOv4GVF2
E+nn/wPJvLLg6hyB0aDco5qGic9CRyo1RmjIAJmMdO8hXAs3ERKuZ5j4msRo
y8YORsxKXgvVOsYDZH7Eosswjh6n0sxxQoYZ9u+liU9JbVG5n0XnW4oircXM
TEt8IwDaf6ftuT7fOC+Xc9X4aqppharqkdRLSO70LYix+pmh0OwvWZ39Xkde
SnzwOY945Czg5NeKJgGqjfE2G2aRkBz6kygcTtWTcdJwCXVCGc07WPLDIH2o
xzvXu2J/zvF7REM2jm4j5SPzGUilZG32v+rSatvz4viap1gzOjg/79Pi4kVr
8VYF/yD7RtYVYfsp6k7nAUf7mXfGVq3SAWZB8By0lyRyZauaX1kK+SS1ZUqv
RbdF6pafWNdp+udeGATzHFCTg2ttSlTNnJBPJ89+itvaml++WlaQGiqNatm3
05MUTIQ75myStVPlWLJJKYmg8booFEuGPYz8zuIqhZi+mL9uQaZSsri4/0B8
C+GRqVsTg5n9pW7j8psTereZ43gf7z6RpKDK9VDCw2Rkq5wsPN8CURF5Cebx
Sdg9YMc4Xgr8zIWCPIPNexjD+5x0Og2fsdheIhnefguRGR7ehTrZdw6fPIjr
gkv59Hv5QyfnUaypDvQLcQnEs3RHDI8ex/k9szdC/rC9xwguHPEmI0xOYPle
Y45wH0vDrcDauukPYlSINEpc0ZYVlIn50jaaKXMucozvbEDlqeP5ZLhgltnM
a9HLbtjbP+GQkwpxrGkQpsoO49ZSWwAw5Zc5xH2doqmXB2yQkCTAYN7tYIVr
BStb75vwbqxurV321jNoU5meFoe4CT2SW1i1/0c4OK3kLdi2lCAJOIrVZqpn
z9cz8IR63+v2Pue563qL05/Og94IxINdQEC3cw5jDKUWGwFryHWW+ktknwsG
/M8uXtYJDRBt4Ctqiu6JDIbuAC1yz9QKmR1ZX1ux4FiIntVnmI69tpv2VU+u
YrjoVrc8e+E7Wkb1T/d9GaxIl5YWx1Cm22kyTW/mKSeIhcZfbjUjDq3r5rm8
5vEYP0RGI+ijj4x279X6eEp+gJIKjDhh+LD408bVZQtr1NsWrHbSPKG/kTIr
io1EGFCoeDtbnlADC7iqIszdDeDy3NEBMCX4Iir2mUHSXxOEAFgbVqHZz3bJ
b1s4Q7L1iFT0dv69cVuVm42BF/KXlQ4iLgiMlKFEu4Tfp3AilJb5Mc8a7cbz
QL0EvJ3wVrM37oHKZLoYpNIbG3+heMyhmLI9X5yfVcNYVFBC6uN8N2H7h2uE
D5bJtaH2KVCAItWItnVPhDkpPkhP6kLIhUson7N7oqxATWnTJySWPV++XdMf
1yXzUFCPorQOnBmHIXvjB+N6f+fDLt3/BB1FiOMec3BLpX/bMJMCF5QqZkRr
j4sWrPdjcN4FOCcUySkKZTo7JNnx5ioM3WZI9Pvr6zlxvPAfnG6SYCAtp7tt
r+5/R0GWpiBxS+zU+3n6yXfwgPw+WLqc/HWILcNqXh75xoza69Z7q+KZq3F0
wh7SxWkX1HN1sLq9QbQKx+TC9KKSb6tDraUQXOAtajJ1E/DTlNnsAwwtGMQj
f59BUjxSjvT7h6Q2sh7o1qcoU8qsd7oi8zQV7t/BM6XF49HS1osEqR9ey3At
XOIp3p8ietsyrSh+Jmeq7ef5xqOEBdUfZOl7PW7ymjN+bk/6cElg4d1+4+oS
yDilkJ5S+vLXdU/2vtJwMvYXxH2ElPzpI2N/wV6d5S0sXyWGeZiCf2kKoHU1
8kwlxMt3YZphjBkyq3/x5StlUT+4R8ScuF00TL5w5dXhy9a9jljtNM6DZExu
DDeEFt0bc5KqhMEjHRz7pkdm4pThfLP9bnca7AtwOWH5rqkf3wMuUq7C+LPv
VBYPxI+RM2tG8nUb9BAHnj9cBBjeCtwBEbqbS1qmAuBeCgecEFgcO3lN7/CJ
Pay8bOJ+f4VnS95KbIFWj6ZTR0SmNj8EwodLqBCp/8lL+2eOln0zw8PcEzeS
LaHALmYBL4HRkTrQFh9AoRbnHkFCWilpnUQBV9gDcxoQNMUM3UO7dGyyXJ2d
37uTOyFvLEBhlFqbFeRnVIQrad6b0zIKr8amDVC78xhzIgjbpUth/wIAnriT
YAzi47wQG/9H9RcBKGqZiVOIUMmtX7DOms/NB+7P/k2ex+udR/eRj42zmGX2
d34WCs0TUOmf9YkEt8e02LYsM4ZLsir6ipFKEvD5e0BZ8eqYuG71kt0F/vUq
7hl48Izztk12GvU9E6sIqNShTAaO5CvPF9OgNE0sW+py9Ou4QITtjiliNNZw
7jyCIlnwvOxDh5R/y1mT7XvXQKeGqjuVw8D3NUk2ILxCZjCqIWLz43+TRF9J
SsIej6zRtikx+BvcTPeP/WZ9BCRNrF2aWaSuIvlu1cDEuZ7lyHPlEGSH9Ij2
baBHaLWKxusz8is108gbde7HBRB9pTBcZBF2mxF7RQog5+jq7bZYHCMpnNqw
q+B+l+RsDdBKiYlUDYlnpsFwN0ZmjoSBSb1cqKVsHCYQuN6YITLg5ObU4lKB
WQH7CGmKfo3xTumqQQSa3enqN8ETg01x+X0nfWdV8R1Ydi2GdirunkwNG82O
WsoaKpfk0oKBlcxM2Qk3nYWW6rlKvC/U/OW6inpRIrDHbgQDon6g7olc2Fdu
C6iRym6AmVePcapfcQxqyjmBSmVpFUsD3Fy3D+glMy04zbjoG3IBaD1hb29R
vz5F+xeAnn4/Uh/OMmtTn4+sfPIGNXCNXUjQYZEZtYIrT3T2CiP23UnwamBz
VRQbMnNV5FZ5YviS5oezmrbgIXQ37Ip9dA+j5xUYwUQt2Q706rvQ7ATgmuH4
inErX1o9zfGiCL0Gt/wx4WR2IZE8jGYqBNPLL8TJp8hmYdVHNNZmFY/mpkw3
Ah5MMpaboFB8k/4rp5/LFkSZpTJw6fwoEHgnPT+4kDxdFmtF1T5mde7KgJB6
U1/nx2UYSOogsbA0/6bHN2/GO4OmNbls3PhAdBeeQwYZDd0SBZ4Ztv/ayS8j
BWQo0YHYQcEzbqAiH+EhUSDQKmwlzNAoWLxtjlI2lR01w40yJnYCV8YLqubz
921QE76drHDcsHnWzQNnLOY4T0Ob8Ku/KCorvtHH5jA8eWFevSeM7EDuGDm1
cTx8HJ8pYupCTPe7am6gzlGiQJoVR75Av+KdMwQaE+Qvb8V0yns8IUUAK/Em
vF/SJdhup+xiBr3W/aiLAHO7ETvBrz9DNMoMcbqG6n4ZqfYIdy0A4aD4lRog
mXoPw1hNEun50Jk7vam9tmIgZO8uDRUfYBHnh5H0ZP8FCyi7BSTnR7mUeZDM
5UmdwGGnIw6thYeGesw/JTAbj1X3Si1yZVudiWKgYk4xhUYaDaLgCQD5z9sn
g6VdqNGg3F74x4z0vcSXAzG/pduDxGLRQ6U195EXTt3/xHGiYj3GcumjH7VY
VctuA9p9fn6+XN9+/Ymq6H5sr6UyRFPRSDQMMuIHz5bo3za48K/6nLwPYdqf
BhCDBwfs3OTOW+F8JVkbL+XHJ6ygl8QbLDWieSsLYAxVs1hdiAH6jHcHvhEe
1ky8XnAGdXt4xyW+qirC5ZR0MKemwSU5caCihi0tPKMvujrfuFmUkl0qSs1e
Y64iVXYb/ql7jbf0fQMOs7LfrFf1ycCtr+YTtWgVRLUarz20u18MqbZH/ZfA
Qr+fkKf8rsJ6twA0HTOHMlDuhArem50lLikFgG7/FeveJ1oQUZ+N+4AgszpL
CP4tUTcclGOBqj3F2BV87wJWsQnDFwLyXNuxkaXl2DU+tEMSSxK5jlzxfVgq
nDIzYzrwkgDZSTzpRcC97RQ1tJ+WAuemUEik6QQwCRtQfwfEoOS/VeM4tIzH
ObymQf4o5Nd9BVEmV+SxwRTBe7EdSPuH8a+1+gLbRIq0gropndsPH1zCQGHA
bO2+1wtrR7Se0d7EgtpL/g92wcubz858Kw0An7lPddJzoc7HYarmmw4fVooZ
7Q14j5vk22YkKpp1le6VoC3nV7AGDXC7a3ZYtVQltiyhunN1oeFpbSiospB6
p6Ljjd9aTtOQ/6hQiom8bvVwA9k0wfxJSgVS4lYQiek9v5jjB7WMyEFk4LnD
Z8eXAYMU99ySsj6vpZ9Uex0EnDfM9QRzhZRyddOQ6hKdZ5xP/DXt1EApqXAy
Wy8zvX9NW72bPqYWcHHv/XKchkui0qggylcuA/4JiZpHqtT+vNKBng+x0Q8p
47yYpH/h84tWOjIKORH14qiAo3noC7h6/bUfjOCVHqPhZzso0K6EfkIiNpVM
yzDeHY7vKswZa0Mzr261m3uFtjEPRx/ABao9XfmCYKPSdFd+w1Lx9u61/bKC
gomjMFp55SHWq40YaeHmTD/XQmKxyI6isYovMz3NsftxV6gwPc8OZCV0ov+6
/3SdeiJvp5cXU8V5tPcAOjlLulQVgEMntjBoYUhq3e3da9ELdaGVPz4jZ6eb
CO4Fs7IfLcb45dJoDEq22D5YlsB12s+yFPFVLbmSjehJInp3Xslup1tUBVcy
KLIkV4iSxbDVzGncK6z2OFqS/B3IyXdza6V6ckVQ/EQc+6gsp4dnOutFdqDR
xRt/OG0uNTNh8B/lNB85ZvGARzNUYps0LKoIdUTt3l3DlzlcMuoqfh2iaTzA
NGFRFywbY0zECwrtDmjKywz/+wph60P7t6ST73rHHnoWg86ju97qlab83new
+V6vbEC/2M8na0doU7H4VHGsm1XDvoY6q4+mM4MVHwkGoNnyREWr7TmDKECV
wEqrwjBcJ06mmwjM92hDQZquFm9TjhGoR4B+UKO6wsCPTqvklN9Hg45ux34q
+ydvOcFgtylRcpRPhEd/XgqaW/fEzYNZHYbHY7iNF1loTM1vRO1b9smSDZUA
5YQi84Q9fO79hpWbZnMYTlC6j3jbTWMSIptRkktVgtbLnCnXNNyh64aWH//+
LwKV0xs8RbX6QvhMekx7JZgcwt2by139tzR8kH/qYXI6rhExfhQ9cgonKdih
lahOTQ8dm4WbsiIVicj8WqEGy4dLAoFaik9MTjybCm1VF3ukMt1Vw6YVt8Ss
EMdhW/vUfLEl7Ic+XdQuSv8u6aVMFd20QLXPv5wrOC4GVrHHdPyprTUvRV+1
+A5DixKHcME3grYztCbe1tfUqW0ELxRxmEmLLLQe99ahSvI0rRb5HXKhdMKE
VoWGbW8aOssGQIom3beNNq3xE3Flxhw0C6VbpC5eYXWEs2rNTdjg8ei+URAy
r+36HtlpLCfQfcNzP8UluEfMzGGTWI9kO6I7+IeObdv27hUthTSK+CEvpnbv
6FbswojNjWWNQX3Vig1eZUjhe4Woe2Yd50OL2DvAk8+5xMTCidSzsy8ZSA9/
OMG3RYZ+LlDKLYHOW6s7OOkFphWTRhRA2pDP65ts/QL4HObDLD/n6GaAOSzl
Zvpy70FGzHqAME5TPtOF+ST/zSga9RKTZY30FrVw/GnBheafznum27S2N3aR
c/DuziH3xVlxay1v9AG4xxxlaWESCFisAgsEzW+dNAztl0uaMlTaUX8LCB+B
YOKpV+6GYc17pFL1bLTL943c57hwYMXTQdEIk2R2EKmHFW0p6cL4Jpzg6Nvy
Rkez9OVYiT0HEkR1zqbq4UKuezx5oRgGK53DoZ0gjHH3ZpSmr7hqiVQZMH3+
VAchYdzNZCYtDw6CcnZua0Z06oT9mcKB1DWOlFFWeWSpaqgYqD7DLAJTh13P
xUsjoifOo4UQM8YUUcz6Tlub5NDO459rcRGpReL/r0jAxRE5gjcfN+OiV4Yg
s8bkjko4xkNY1lKROZGs9rq/rMOAaBE//7kxNskqCp/Qkoo1Md0ueczzSkVs
ZboAd5v6Sqd6XZcVBPGlRMM4XfI6UNjN91KfuxFBD0qvb/gLmIDPldFyD3E2
I4fCnajA7L+t9GVBwPjhO8mtUC5+4DoWBwCcPts+IKy/Tmj86/trmXQdf64t
s99TVbj/oHiCpyzVD/cyQrxxZ8I0kYRjJrckyI0Ob4zJtOTYDgKCfr1PqDu2
+NJAn2SDS4mFEKkjyIDC4bN/QodE+gY5vseSs1Ze1AZIbcatuEd9ruVdKaIZ
/y4sgn8u1Q14KhxjdfFkwAQ8d6MSBLY3Ltk5dTYmhNYc/9KdW3g+vJ2b2iHp
G0qaU7fUkXaygtU/I1ET0XMa0g2+sRBK3Y76seQv0fo0OPDu8EHIAEUlMKz+
NnEWGLdPN0wCJQXVydrrSxSa6gLtV0MRF5OdzcYQ9MDimZlf0WaCJq3ETcrL
i5l1bBXuNuuBPb8zGDidnUNOsebr7JAmU17RxkROyh8lzoc+5M3L+yUQfweh
A3EUGDqXaHAWegPw31f7YQaIIauULcjb0hYShcf2c31y9oqd9d/vVAReWiO7
SdqTOWr0LebIxS6tMqQJwmLu3vugcU1tK1a6uEVNiwJU8sPNWzH+JVTXQzdf
iQgSriaeZvApTqZ2gZT5u2meHNf6j56txgFZ0W1e3NR5N9FAq1FxLXbIKyNc
o/g3x8+EUFOVywJvgIg+fuQrLrWXmwWxc45dKcRdlUKzf3K0Xj0cAC5XD0xR
VTVH0lwHdeE5j6iY2DPbRKuC81jsZJ1s2WhltJcJ1i/Ila0FmwqP74Nt2liF
ho2eSXxZ+Hy0ENt//1X49XhU2EjVCXHT3UWh/LXNMQGgNXrq4aPKYxamDdvh
0pT6gCXpwSkVjod7LgZsuPW8jVehhFT2s7SqKdM23ET63k41y+7YYrLB/zjV
3nxeoOg3N1T+fZiCUqBXKewIrozWXrhxscIjTE1x+9sGzTXvZDlOGiQM4qVk
x3hnu/mBBOX1VPTT7wyFGXnVBwtcDeSJgMCMOlWDa3H5xunO2T+mKMv6jng3
0mDzXXc/yImvJW+IBIPh6CZ9u0MOnjSBGTOpVyGTVKlFP4kYVBFIQcxmU5wf
vFMbxxi58rFwj6H8EoIqM7nFt4bLnmTNSv8auvraedWlflw4/zGkJTdhTTfG
HvPl6TrICH4qKqu0oa8ihbAH169lTtrLe0wjStRYbt8tqNCkmbr1Vzn4s7HH
Tq5OJXiyK6DnWXQafMT9az13lcPSu14TDr1EU4Win/bVIpDieG5sXWGr8/Jh
H7hVjmwmvLzSks58lf3N5NSeobSC46n/lkhwYY2CgfIHYL/celYSdoLIUtrJ
G7gQfvgKl6ajQZTda/o05a0dYPYOVdATO3Pi2DSAHaohEKk4/xLA3nUDK9iQ
7GXq70SDgrNUDo2CSIF0e+1T2D0iJM/eRlr0YGIQ7JgNINywWKCkPNs2xcGT
YBZV/c+qDYSq8j9TzKiqLg1TTT6ApLu9gEdLbnz+gTNbQMWNhjwbchQzjsGx
lV08fGS0B0HvyIeCuqbLMkU8N3qNZYR1cokPQH7NUJlwSX8NsGZZNC0Ndx0P
AP1pNC3Hkubui7dRFiQNkqoZYIED5ckZpzzkq5C5oJU2o5FPCI3SAmksWYYc
v53UB8MPrLjajGPkPH221kegNZh1IaiL5nwTiKiuzr7W7BMZ+c8Tm0WO3eSC
p1P6N4atQ/6c3QIePtT2+dkKNZMQ5YDF2x1eKfBjq3hL5Z1HZud7knv/ibiJ
yEkZDh2s75hu4b1VXZnz802hH8v3tra15WutgOktzW7/3r/4oZO2tgu3p38q
cLhBE5uenI6OarPI8JEY0AcWBRmP0yW3zij9a+tPHD0Rf2pM2ZaFVbn8GdnA
Uh4xm2pZRDb1gPn4JdIsxUR73FgHlQH9R4/huIUks76MQ/IfCWpo5gBgnb+y
S/ajV1Y+AmVneXK8mZ3jM66V0grb98NZJV9o2SdCuOIYFSuSpqVy9DZr/1VZ
cuA7dVNujJCNGN4w860ZhaDzunh7+pM1Oi9Z+CaOOmfGdiKhPwvHcNdlp0Cz
LIq2c2B0jnqCz1n2cGVO8qse1opNBOiYAHszy8xcIUbESsVYZ9u3rHwruGC5
TAcAmSh0RGU3FROkFO57ihExpazi6gwDU6Y8UvUuTnX6royuaa/NVaa2Lu49
8Y+nYMHtY6iGz3KDTdNo0drNY4lTon2BP/tO7ixQJfOgJL6C/JlJ2DFc7iau
vM/0rUvgYKlLi3ANE9Lkz+jz3BUSICaFMQUmVdsgRWayKGUKxZUyyy8QJshu
p9DhU06WkIRNB5+B41cojDXSFBHGOrCgBpkrsUSHR/cZN5xeZeug0SPoSLmv
g5oz3WKNPyYI4ACXeeHDkgNBAM44W6bNTDlwtdfWyuhQIgdqmwNXGkLmLk/6
b+usRhDavxEGhfiqYxyIg8uLGVW/GC0XJ6RLCErjNXD9DWF760n3h4XUYPma
aZsD9pBTmVECQ2frO1AJD+GXlOuH1DIcSBk+lNx+C+++BDNMG3vmVOdHqw3T
x8AzX3YXUViwM3KE99hlClCWrPPmwpSgMhHIzLp2TCUuFllayWCtTNrBRJho
yh2LeZeMne3V1qr7e1q1ZXaqj1jeJvsMJBKJEvZP1FYBwcqSkr4AK/zINPDn
75AZI0xJICVeNlA8x+gWDMsBPY9qDqIm4wQ1GglrtLAwZjdsMxcYKTi2U0TY
ijiffFbGoLthsIkb2YnSTCqCgFdPKlnxSGvowL653eopFWFsLtS9khkJLYrd
bV65FA8oBDVnjw+CdIJLVjawu0m5JD+DEQrTSoF9KOQH6Fy29yQ2Pfl8PYRT
u1vJzx+2fqFWj/EF+InER1jcbFu/GPALF/5lHLxz1YMJDZhQQbxDy9jRjIg9
oTVINrJIp/ZDyOH2l6dvnBe3c3YR0dNUJf/kHF3H/pPg8KeKaUvPfiseVDvg
D2wt0poG/2Rfj0Tuz7ZUR+JWJ5ko+kkQvoInviqAkltZtZZX0wPzkBg0OwEx
2773Zwn8dXyaFTGUGA7opQmpe0wz1Ui+UpK/kI8XOOudOzWVNs/cRiAjXOAZ
AZK44krFGaJH7p/eA42n3YiXBTbc7jmHxBnhHPdp+poA4LRpBVkwYTfQbuWR
3H+q9qvtXO4WmBzOIyhQg9cO5T3makIvH2jMBM189dhkmO7uf+DW06/RM27K
SczkLeSK+punmhkkjGXuOqRcYIoasO8bxJ4w8rdiGQl0zmWYaeFBhJ4dYz54
7tgq25KPwvjAePiSeRALKdChmJJeyHazzg7HV8TdG20mmB4/PHVp7o1N0yxd
tC9diwyPeDMS6DHLq4NPupebaMQDgjxKBiKL2oUsIjlrnnw+uc9vR135Bu2G
0dAM/TuwFC/z4ONXdnqiZeu8vYSTIEEFuvLEMoBGnP8c8kCBhaUjH8VdQ/iq
3sUKD7qnqgKvOF2XOrgYmhjy3QCv19mEWExKW6GIo2Gjo1zPHemztmdhG8HY
QDrR5yF8s1DUP5I93bUxwWgqQJw6jWbQdlruNl4IST5igyrhzmeMp45Uz+xA
6HOweD/TyLxUrg+wp4athXngYBArCkZEX/JEyvB5VBHqJhqEMu4+0r7H4S04
+ZeZ6fedGF2+0SqQaFV7Qb1OwldCxQlLkU/1pX+LMYfo+Cjzz8mbYznh2OAy
j5nutB0SOBA3EdHnY3x0yj+OgLRPo3M5p6hnDKdAm1n7FWDtdPDVpp2RwA7t
lsUil5ixbo+UZRu5aB9a7XVPoYfl/O6hy0XAK16ZhwPYSAfs44/mWb72u+Qy
gexMD3HFvpBozDOYmmyIfjQmlUybwV9uFwKkMkh2Ecjbnuw3JLrtZOIJzVte
2nJcjEREI5/o6u6VjG9dZS1bWfhHdhADtAulcmVEe1/w0+QKsHouHEEs23bA
o7G5EzRSvpYMlj90CNTQMRc0FIVcb7J1zKeqOSBTHH9jRxhMU2BiUH+X4BR6
jjGdtUSqnYWkg0ohkDm9sayuyv+LhCZOr85zxW2e1rLlwezCJ1blalPRgA+r
XQbMKYs7b5zhBNo3QycNniFQrOEM3pWkhY/TkNllsKSzJpEpgL7ijM/hVhoL
RbIkgKDE8Pj5Ij95w+ptKBs7F4LK14mZvXWOgfbu3aOeC37H/CyDw0LuUlBc
QrI0saLVAbKpgHdZOt3Ch0et+qOLMSHFUIa/67CDPIBgeOiBg/+jY2xHf5fW
t7YKxN1KumemdlGgRpRGo4LD+Y9v8PBpaohrkDifuZjqgbakf9U29P5AeFQO
n2V5HOKyMeb+fDvnOJY1wU3pUTKJv6t5u6TnU0o2NDPhRiwfsHxN0z3bkipm
vQZ+VVXu3hLX1NeMSzaFZw2MJ5geOpiJd/YLLPUcNZ1AwiVEhR4gmcSB+v1b
hNs8mMKnXzMmhfKeh1aakuTfln84+exEmj8TBrPtL/5XWPEW1wMQupsKwAZs
NNi8wMDOEhDhr8HN5qFmpo/DPb1delY8X8zq95UzHV0zvPl+JMNI6ktEkLGX
DonkyO5M/L3WMRZMjirCopDNyBz0ZKAtkGJZDfg4777AXZNOSPl31J+Gy5Yy
pRKv2L+5ZzZQhfxek6ZhEvL3em9zsd4PrYdGpocIw1GyjY/msRNNW5D81MXZ
3sw26FJjwZvhj3gazSg1/M5MZWB5jd0EybbB7IsAcpdb7L8H50i4M+kVfDoq
2bqDc7nFd3c89BYgTYhY7EET1HaSaRk1WRvJvtxzvvLruE/otY1iFfqTuZUv
7IaFp9L2mprapFo1IJizz2QvqH+CVwedrP05zmb5NgZpRloUe3lTFMklspcu
NcOxCXT4ZE6Qp7WXOD4BeuVbVS6rE3acJWVjylb5L8fJ5X8cx0LXLLmEn3dM
paSdPxq2vUFPpifURzr7npkHijXhyVAypFkOz+Yrd/QLtHdDQ+xvhPY72v/G
tWfQ7cCh4se0Zi1UI9+UE4ivLzkR92pp3i5z6sqqf35KFEGR7ryEcToTwc56
IK6R0GOJBTq5/R4YJVZKIMk22Rd6pWNf8dT+uUAMxwmadqo0+0vK6LrjWqPM
lAYjWEUDlQcriXI5+a8sjZO103yerWhZLgD0g+AbU4kIc0ms/1HqpMCwanN/
x12NxOXH8RkgsgXAMCFHW96InaAYJJMQBHSR6ks1z2q8ibHdGlmjPm56Xh9u
frr6q0bldldt0kUqw1m48vzzNukiVSLnC34H/cJfLXTX/xQrUkiYRXbw4hVg
Ul0FIfdQfW3g67iSz5D28VRYGZtjoLTamepfHAdNNYyrJ+AaHOY619CRvgC5
p53YcGWTOjTwJgQD7It8D5ggaFEn2D2vM0MNXHpME3pYyLE8hNQFhghv+zYJ
c79vYXfbYsaraAjHfVVDyLdj/Va2YaWMQOHEttCaSZEl0IqxE7s06YDdRpsx
UhJaEMrhgXqVRc3gnq8V86eBnwdyFQo230cx8P9L0FT3Y7abqTp46ouGF7N5
z45WhV3+mE6CWZrMCX9ceQQURNnSM8A7bMunUAUglNU3eVDNyqXksTOSgJAo
qwGVIpFq8/xwnEqr+1u3vXRTLHKkJzZ4gr/1issMtysET0UpQz5rmGI8F0zd
EB8mUyRpdQ+/WktqKFG5Z7EsIVtMk6H/Ck3gEnd/HnbsLKWt6G18zslNyvOn
vmbEFJEld0cH3eW4w6CqIVK7cIkoeB6dE+jJiitgE4g9U02VcuoKaoqYdGQt
tqXmq1DlwZdS06b90VVCN0BOqNM9vxLZENEfElebt3MDRfO/umBvLbvFjfwS
oSPHnAwLu1OOng1MSk6WcE3TRZbmRF+fJasfF9nU8aeF2C59m7vibKRssjKf
C7aAY4c5b0kUlNihz2nugWFoRebLMdH67EbmV2OCy2+4TIPYtgruB+XFGtHZ
BBjUkoyW80AO9WD88uv4VVDg+iME26Im3LE6xcJ+DKV/w54/+XdU4etEFTj1
c5NP+V5vy3u+8TXzFb69G69OyIjHGhl6++skH5jDDqt6kFuYUnEcWMWk+Q1y
dRwvyGx0cRyjOl6IHhQNFY861abmCDeNU44x1D83C+c2pzb7uHOiQnG3e664
69Qehe3sD1XiY9cIcsA87goZki8DDW85Zv7OM2I/RfRdeEM182laYfQbFAsy
1k1k61ohXGbe1FCK7mR96zCQids+tXqRl46Na684bqe7QXRDiLXD2+4KQy1t
ePS62+30jmGZkB2pN/ZhxykQO45ckcfyyXEl03C94xSid61OHjHHn5mZ2T6K
PPMm6+vvYH7oBJYi3jFGcIOPt2msyAV38t2F0A4om4Js7KPXJgBmL30aU86c
k5KDtukEBQNYV/6EB3k86yQfTC0CUu41bMBR0dhHs7V+k203lEfxIpcm2I43
SNiHC/zkgJVet/B5JLvBvsRpVqHNh8usks2CIDhTgaubY5zQGPS9HAP4JxPp
QgvD7H2Hw7iuQLq5TQ9VFQ1lFuccOM9fLzj/fbVjHibCooko6Q/eVTEseG5J
jLthh4DKqO0QjNwxiBiB2J/TSWDHjYvz+QOh7U7aIaYZry6luHi2t9gtW2iE
IA8bpE9/DUCoCcWk7owKXKOsi5XZw5+0q88E7JZWPt4kJk+ksZ9XAjQhFbVa
L8ra2L5IouW6lLClTWbxotTnp27y37ldXlKT6J7JuZ/PG8uufVgxfGRanyvO
wYrugFfYR4IMyjumCjHt29AiiwOSwWvrnHD2Ek7YsBd3Lm9i/YrSaUQwX519
WIPICGC7zkh5tqSSlpdG/3pFiCJhMHQe3lLE8i8IdrKr/FVmNrGCOCAP+r7g
I6Nj070fPVJeIMNPEzCYIFZlOG/Q8Yoi2u1q2Y0c8P2zdUYTV62HjQeMt71i
/roq3KHQYqOqaCb5ZfkAxN8Aed0Owu/UmUUZuTYZTB++kQS6NQ83gkaHNZgK
0jZtYsNf0JYetYlF2qavGia++5sNQWzMGmdC11lfwG6QUU2R1zYfgikqJkF2
bgRD8Ae6QV3TobFPCAlAzz2bMJn8MigluBTRlVJtbQnCMbnoqSDLJ2/vtK8q
a1vG9GP+Y39bSA6S2nOpZYi/CaTTjCNZkibcDy/bkYu0hAm2VI588NNRHTz0
l2VziKfj1Rzbbh7c9vHiOFJtjhXf552L+3ZzdUOVoNljRFrC7qDOUXeT3wqq
K4lVELqpfnyG3dLN/xi4v3TqjInJJg/nTTuSGSowH4BDP5oEAJCcFmy7YbDU
U+wJOkKSWX9+LAvcUgqGDiwcnJRr6ggjTDI02j1XfiERY8EQLa3G1iSM0o55
49X8+DoTdyfwkl5/eeIcahmtOLAmAQ77BSuEJzw4rhnCjjz7ydYZaMPobD++
NITy2Zhe3ItrZTqVr+ERbFJBkO/xLNwhRlrZGKj7glXRK5Aw7OWOfo6Uxlkx
peUIj7TapbgTWdaD0OhhgXh5du1ltkRxTbTcUwS9n0GWdwS0mz3X8NarGrMa
UD25LKZDboLRa3hUTtEhSjINY3SuaNn/An+FUWOE3abAYD6WHLPBgEr6JdQv
xa6sSqeZJ/vXC/vHAvUTGyGFj7rUfDBNk865c7WC3Qh1DrB4uY4WrqLhMk7k
6axYv7nksJP5/73mBH6LFZ2ohBcNvQ9BOJVvVurh2FSFxkelgCuslTSVgIkP
U0OsV5vTKUT4o98W4L8joomeGIor3dqFUYHq4EOQmnQaBLy9Y8te+h1TTGLL
HEyz/HjKbfhVRaMBhs1JOibicErbTMy34NCkVQTjeJmy74CPz36LvxTMJo7H
7RcyIj+yjpSvoYi0NJyhV/oM5pUJrgMts/KJXif2HfG0LEvjWoLGK2urNEHv
X9sdLDzkEmDYaPwfFyEfu2XsNW8x8ibmRm3zm4K75sAQiaVz//6qcmSQPekQ
Ms3zYZ0ua2tqnZzrQrvHl3aues1+WEbzquOKG+LJv2nuRHl1FAYPQ5WImuAd
UtPvcrBz1J8pTx0g0tgUGyh9IVSCBKDRERPVPrr8fQTUMwykEQEvg1wXcuAr
rbS1zX8bJ5Qzvzq5aJwKHGkgG3KbtCWY5QXTAyvnUnhhQEOyMTyheErSAYp6
dOboeFX1WE7IPTdEXTG0CQCSYg4ITANKUEvF8tqB+Yjq07Z0XZQ52m4msDqh
suRxEq2GD1fMOxwwpPotbDPNI7eASTdeAd3MVQe+ZQP20y2bc/CajuXkJlN3
Ft9+1JO2H126YCOhJEneVn85i9MflY4ULmt8c/DFtUbjyXkBUJJx1tZkmJ8Q
in5+uRSrjx1xwBHk63VTjAdQmmvt858BxKhwty/FOcVydSmKMUK9o6DyvxTz
IUbyVVo3AmxzO5hn5sRvc0srsLP+bZj11sOwqZ41JXixANMYCjecHNRul7ne
ddsnGIhfoCrU9LCgbO+zfZKiNYxQLW9YkWIKTubARc2YXaIx0iPPuC03ulmP
Kw3ALq57aj8OAkb/YTCc2uGcBtZxa0hFomv4maEoQpfDMr2GO9fv0dWA7RaG
Ik/GHHQHRhcmpmWTsxyKAjBJvuTSYyhGZfaQpzHniDboH+QV12OMXDEcnaFN
FL1wI4kKyI6lYE9duWu8jNnjWypirTee8zLZ1YAqDTqAuLgdVka/EiCwx2SQ
eA9Yt4Cr1Ps02wNgPP4sTfI0+dy44FENB3hcR6KDghhyK2cTdg34ou6EaBqk
jtcVlXLWnBxkHuk5tLofbN6PkAlxpn4Uc3lMkCmBd1YyqDcbC8Rb3Ku1W7Pt
9MRFrY7dSpsQz1R667tGCdm9RKd1iWEqpjb5+G3Rz9uArrpelHbU54YcQO5Q
jOFacmXWgnHRwdHcOVPJWsI6h2TTBPSe6MhufrMqtROLKYgRIah0OCBAdevg
ZdkfnrzHf/jy0uS199MP3F7HBMv2I/X3ZijBMWSh5+0Z4PkfwCsNboTeU06z
tJ4VF28VeX4OoXbThYhsJ8FLjT1nv/V7y0hg5ezUbLjCNOwgg0dSQXE5yx3S
/X5mOu0qbb+MscVJ1es2KAEibYkhzqVDay1o5C8m6gDV/mLPHfeHMVS+AuHA
6VuX89Gtgk3itW3npY7t2UnPXN7q1R+Co6OYx/Mxp8jkzqACmZ1BZncX4gMU
rllMI20GctfkHWnXLRYePMYSSqyqAp/c0dn7usuoblFNZoPRX4Mxx3FDiNt1
gRYOMHznHvd1gBIJKPjXVFtw/47wJPuE02GZnCW3NVzQpjKs/d+7tFt1vwPD
GO0EUCjcMrQ6B5LvqJszs+Yij2BTxcGmQypPwmJAQvo03BVpYFRN2kfWSX3t
8SiLT56r8GHI0Yd7LefTr6xgmMI1OcOl5nAk58VHlykBDH5wbWrELgkembea
u3vnar9n0eWBsXYJnrZJ0K1hVx8rGf64zRM3CfziTkp2084e9dWa10oRs7Sw
RS9YAtC+deaRQf+P++ocuKeuNYkZhXsuZBhqk3XKAzwG3mpxVSF/r2djyaB/
iytSahpFnaZ/PKoUMmYqZXhAsDz7srsd9tW9W79XpzNpraR9JrUmemERTLSA
2gJFeErP7gkUAdGz8kGgJEga2S813EFEgvJnX1H+sPLAAo0ZyL/OQrFQj1/3
O8PGDcV4ZXi9MENsJvqyOaFBBohog+mTifh5ncYq5Je/EI6lqzAoejibdjrg
OLNUyTkUyh2Igx4W6Nm0XpS/39mDDSteF5a8Q+0YVRk2mMH74XZmomqDIE13
hQLTyXBtWc291siv7BIYhQ0ztGz+yV4xH0FQBouYrKgG4YZm9pBylpz7i20m
OiL0/qFwiaHbxBx1mG6xKuPstspzZxB7QB+nGENhwSfRop277CJlpl2dwktd
Uv8OpFUPQGypQbi5hAiiOOC7Hi3g54tGMBTNPjklGDj7Uu3oyPYrR6BctB2F
sdHGGianxRDAS3I4xju8jQzhADDuya4xgKXVSplKc9a6QndUxefVYOoWYvRe
z+enQeD+N/AbCPzHlWZf7f2bKtxbDSl0Te8lIVmZlNLywVFncKpdukisXIGo
Ze2OZZ0qoLhirKEuT7Hz4vH6kraHDVK8Pqj1BTMDywARAGfptuRUWizEm6s6
BP2TypEL/pIlyQ6AK/L6/nQqxWE3EO6wPdkUFIclHhXu6a0MkoJbgAHWSoQC
ubN/8GZ6D6DeeLq6r9yahaA70nEwhXnZH9YdLr8wBu6vflM5pT25uQcK/WnJ
tDaGeUA9e39fFPSIGqWvDInlR5X3H/mrp4+U9nWUOg2SfR6maMoY7w2Ygp6A
xLmpzvCVE9L5J2RuFp0yvC04iFAHG5BS6a07645kdRxW7hYubmWNv8ZpYTde
8C3jZWAspf66wFgDvjGqVWnOaIAtlH1RpyLe4PiSlMGxoxoPQfVsd0pZ/TR7
aQx/1ywkS3iuw+tybvF8daQzl9AdogitHa/vy8fPmNt4xZXRHb0fGOfmD+3F
WUG/IfB3Dr69sWmrEVPGDOAXevdFTPXu79X3qnHnAiolHFAelfo3hhQpbMCf
Zm9Uhwk4fB4HEm+xtYYskp9xHj8c4/z9o9C0lFodut1qEsS4HxTBcqdXJCdC
ax/R3/lFvaLzh8io1yJVa6wo3gbwKYAdkofxUYDooGQqsw40RJP4r+v/iOMp
KUNU5OSmsgSACSQBd9usY4U6O0SxKTrUuB4y1tVmigTc4qOKux+ZrT4RNy+t
wwkZ5ul8lfaMtn4OO0vjLdRkvr0TgZyoHkdwoLO2o8AaA6wgskFYkjt6j9th
QPTQr4Nxy5N2o/GycGtCotvO+EOObGIQovXlRbYMrY8IwM1izfHYcfjr6jvj
/ZbpLMtRmlLZk5+kuBYC3na+MYQWcL7mP6Y0mb9urGrLp9Xd81d0sDEwk/as
jicnRPVg9Ao8AZhRP65TzZ+pd4yJDgg6v95/outXdxr+N9tztYjDKff0fZ+b
WCEx4F/jHzJBv8QzLxFc/FNx5AM7xU8s1HakAedDTJseskzAqNPM63o8yk48
zOiLWk7dYoOPSiYOZbfBfNQjNX+nYQc8GV0Y9viMpGSpV+bQt3WvTglHs3kE
pwefYk+mZOJLBv1NQ9iQmlS39oaFCHyAAYr5Ngc6ktGlm689Q0jcGGylcqNW
VZJQ8NjG+CXAd1HpLOKyF/t3vSKt2FTdMCIfkusUMl7feUpbzQjdjA7EpKLi
HSnwzFyuwib6WyDkUuUsEGDfTLLhvmyYeOCsJ2fByM9XNbB9jdXAsU1cbAAi
l6o2WDtljtSUWk0JSGJMthaUaysW1hd/8ShBsTOpQVxPQO2nfWO0NxnWga6R
0iJ15kk1QOHvPlr+FF9x4A4QZE4jSY2Gds+3Tt7K6BtrCV811EdRydlham3b
XN9a4UTqEdLKzMZbUCktoZPbwKm40m2M3cQeRLkjWf4yIUVywlhqeNGYNamg
TmIpi6gCL32+qCN2/cVoJEiXLdvvCvIxVrsQFuiJUNEFCfBf9dmcOL53VxlO
gOu38U2fwlXyzi+cuTrMguATW1eldbksdx90omCWfyU58mg4RPX1bMBH/TtB
nL8PaNMQQOqEN8T7+BzEbZd7urnYcvX4OAgnXLVfrNX/tNCfk+LTuBHmSp2v
LFhoVVJ7bWJPXoOP6IZ2bXXDyu0Nk5EhBSBIrWiQQDVDKqS53XTVyvSJEf9f
tCeO9EXcYDh5vkVgzowaim9sthJSJziZetDZP7prz2kcl+SDNu6MqITfIn3I
e23JldFcbMBRyBqND7ck5QnxtCXgIXRwKxOEJsi2Vb2WiHd+tzF7tYoc+qGG
W70JfjipoUkD+EdstwnrG0c8PxFV3C6mMBMKPa9JSK0cnz0dfjMYWPaZVQ4W
onGgMgmGxtVFOXmGguWrYwVnnNLJ52HDoNXk056AXZMDzr1Vxd37jIovcAOL
vz7O4QSo81ZfWBNjGVNsfrgOrswKkJXYV7omXcMfaoiT65FyWiM6l328S3VG
krs/4z1tDSk7Lr9qKMfHPLk5hgeQaYAz3WFE/H8VtTdR7khVhV4d4YzFpOMd
DE4/qEnwd0LNTip6Id3Wz8txNigSmi3Q6xMPztsxTzHOrYNxF3GR9WpQnIZv
FNNHjualIlL3utVNT3yuLRTxYiHxwd0NZMJ+iFgbTStKrpE3RMv0q7jUcDZf
G7r/s1NMDl6o/VrWYDMRSUHgvCpGeAz6ts1m2KZ4wTUQEUnJ9au8tf/pBTho
iR7G+r72F/+07m2CH+/KGsRDp/17iL6TQ/AN87VmgKZJb3+i8TrXZfaEx5ni
30eBZnCIds6IlgwMpBGGFI1QGUuErFYjlaHxQY9/Ye3LJq8uXA57t3g6lLMH
vj8QDo/hNQ1ID/qbUx1yHbAUq9vhDXKNBCcH4OGY/iSNAvNvc/rclFFD0Bs+
VFdJ0qz0NDsWxc5Tlf8tGfmQ9F7Qj/zTL57VcYOqyzPnflLPPyqAu/dtNLIv
AtBYUod6DkxdlVHNHcUmIiQD3KseiqPwjlbUMHxbphMdXJSOMPkdM5wTue3d
2Pva+/O7PvcUCPaiCkPFqdKfJt7D6OsLekmmuKjL9FLacxd6A6TbUwLXEDff
o1wdHiLdz9+muCBDZbToUlqLmMAxPvmU+crbJ1cqh8/bgvQi6KunTmwU4Ju8
YoX1RwHnEpRhimqGasEuAG/PVCZ7/49TuBQHjIeXl1fPnRX/vgNuI13naert
QT+wUvv4Xx628/bwlWAZVlzXII2B4xJ40+gHpyvCeh7VVLzl89DRhe2NCsmi
0n68by6ctjJB4PGHxiahXDAPXeLWeovetNZVqEtFvQcf6S38wzs9nAbYNgtT
mofAoaIc6wPOX+1s2vcSWKNsuHKcyfs+YgzjVGRHtrFjWHVrZXxPzz5jusC2
zO8oWssMJwcB5VsOI5MtNewpx7jEhZNA6CWHbbLg5cbFJeSs4ttbJ5MRdIfU
wccFwYmE+OskkUmGbd2MPyshMW54uYZCbDXjG1Xhuyv15BeZNEH6VHGZ9Xit
4eIbDGgKw99p3965DuXyoBM2T9oM0e93hM+o+qxIE+OvNSOvLvWcLd14fvnu
tI8NEPXf7sOfEbA7aPooBfCX9hXTX9gDfIUz4wPug0JA+MmTWfXDPHYFZB+y
+6h0i/dQ9XSZ7GDUYzhyYCi8H8l8+zgXwxdRtS7R5Uypoaw9EmdIEd45AYNE
SQzuavUx4p806gZprv6C/tafDgpvF9KzSjxbN5lw2U3DqCiLfHKqU6lt4lhP
2OX3TqgkHnO38QW1FSm4qatIK7Du2TGIHGA8c03DP6CR9VGwTDRNked3Upg4
+4zREU/vpJasVmzZi2cV9bivrV2bQAPE+94y98bjvC7xuxTq4eXp2HRqzgBB
fNOEz1DVV5OkujJ1cBr1qOiivu4TMluzMl5YtH55edix3fEfwU+9XlIfQwmi
2ojasKHdBCu11fz3PINi+9ESxnxEK2cVJSfCv5zbacaM172TYoTdABvk66n7
emZjqJEsiY3ZNa/5LOJZJCY+ftQuoKh7sqH8eMThmrloL960Pe+79qkTZ4/A
rWV1VrNGRs00ZCMMgz/sjq7L5KBvCZ8I3hWHOTMYwTE64P32pVnqIrt0qu5k
SOdVSoSjDJVkNzVZsoUUMBiug6jlqGEiHh7PawA70glLB80RPxCyfdB4zCkL
/1bKczxvt/ufcJ3bJtbaXNPpI67Jl5flJeA2oWWhqqI0p+bZoLUiyprMN1Ue
eI6ZzgrkUr8i9KdJ+z3ftsQBQnyG/bTDfat8xajduPrQsPK/fNFkvPXh0H+R
EatiQZeI0c4fhYSjIQLD0Oyx2QWrvTinInArm+cAeHp4dP5OMxS02Jw1HN0x
L69tk3y3n87H+jV7zUxVQpU1cn+xY2tygNgrlYU1B9lYOFRYW896ybreGF4p
2Xj8RAVPPUP4WbKZqHoP+JxQBnxltSC8F8W05+BErBPi1VXXzfjL/PsO3iKZ
HXJxjC38A/+1QXip17/G/erdvlp9B9spAlLM2HkB0RNK8sT4tWad29x0S7X2
x09AJqhCtCWX0ZGBYGprnrpOCWVs80Ov4fDviBtxUuJrDIJla5BqHRj6NuRs
kOD2VyvcCrjkvuEXDPLW+giqRCgSPC+arCDyrQGWeRJyFT07xwp7d8RI4rGz
P8vtbAoflcBE5WYlFHbi3BnrLD16hlLtIABcX8DGUWx6qGuBbsfVCB3GwOHm
T5weXZalGFdSWZhgg0xXn1TPvg9CRxpVEynx+kDLWP4osoE6J4mjzb0RJSef
XQld1CJ4qBCS5jEgPQT9M6BTVY/mXUXe/hz2Z/2aodG7GcOr5jd82K4m61u1
OnecI6ikFovOkmUUOUm9VTgFEA4G0WfP3f/UgrgfH9F50r/669N4kZQRL3aZ
KOJWpwDDzzLs0fE7O3vv/llvTU6kvGmwZqLo/AX5HVOdADPCBQ6QeOJ1xXpT
qYKl1zQJ8b8knpbcOMo1xSLdx7A65JR8yqsjVBthpzON129x48TbEbknnpuF
Gg9R0PGhubRC1HL52aSbqNjaTujCfkGle7nZZGOQMXpjptr8PrZRok1rxRWS
2pl8/BI6hv6p7yRHYqgPr+IhZB5WS1hJAcZJ0N2THsy/eXMVpiVNSi/yT2vs
KddeUcqroSW5ytlG6RaTjZC7Srt7pxglgHzp4aGWfYepz7FfyPNz75/MP56m
lHXICaHpL2oRG5yADjfD00CTQ+rCFIy5PTykVjg236E0zBQSzxuGvWB+89jQ
I2NOZMQvyAizZ+XW0K9cq4g3cgx6MOUJ7h9zoD/oJRLOLsplDvNG4kl6+0ze
EvbDGi8KgMsONsxBsk7MiXgGeZOI5oFNa2RDZ7GwQdK09HjuQlCFytRnQHnf
klMIrXLoEwQOmiLLDOzrv+ysKRJ/uRZvB6Ka9RdQC4xhx6VmKF2ltc4QAOXn
hLpIt0qgyCdyKUGhPe5DJ9MqDTX3xDhrrFs/k3ecx0xtZjCOjYhHVBc+n3J0
fAFfFRmAmHQPJWDEjKlBjedeoC9X+XBgl3L9o9Nz6jxdvTegL+2GuueYfNGc
JaWKF128MXuuIfchV98LItUz1xjPhfI5r5EChSWx2WO2vmiEeIkiFN2/FuaW
NZZ5VLthujPZdd7Fyge+Osw17xL5T71ob+dACN9zy69ueY9X4HyMsF/zYTDe
UEzhKrVtO2f8eudPeqvWKYKIS5Fo9f38Idmc7eoP+/XNON6gQn2skxs7D5i0
RvjWQBqAe5PcqS9ZDX4YO6F4cxcIir8uXk9CYPBnKJxKZN45E2TywUcHlSqI
Tb7xWOEOnZGiBMelAe8U53WZ2k0AF+ISwK58EooHUKnMebyJ/JjF5BYAIhR0
HffIyIfmdv2S1iGf3Z6UTKVYySQq0IEYayWVB9QTl8Uo1k+WHPvrA+SFAXnj
iQS+RcSpuzjzj/A/tmShTjiThikhW46Y3b46QihPvfMTGKGWjwTmHSFN5f2C
wwSqxpSVoEmxxsidkLsqgvaOE+SSBXIbs7peLOhPfAvfO950CRb/im1AIybN
V11zujZfpcQWbqXTIrBjZlCJIWQodVdtn1jlvVwKVosGbpC7QdCmrVtNhZit
lNUcza+qeQjkeih/Q3/oL0XNMr1upoJQDzGt71bjIqluZZqRrLkCw4YpDi8L
NFB2uRbziS0fn7ROzQmO8SodOOkZQWLYU/YG98IrXU+xe/UWAkNCN1KnU8p6
HuL2eA4fQrxEhN1/KMr6gYHw3yU7UBhellafTFQ7xJwlzM6U2p7H7Ju5/jmH
vuMaDu41OxsPLjDYxF+ltbjZ05R673YLd/GqVnrVDFGPIfjrA8z1j50hQKb7
YPVUGvHjyjVNnywquzobvxXaEsJr98PNC8JAa2oqzX1KxKgfz9eYPomJRhwq
liEX3RSK39HUG92JK4FsX++QBN5doIZuJe4y93CuVu8q5J978CYxkM3qpm+M
uQekD/4ywgUKTXzc1IgmHCdoWcNGytIqc6fky30rwj/vjDwK6rQaAtt7GSpT
rDqWtgtJ5nbpp/KXbY7ioQmBHWXBtqZwdgj56ivuP+F05n0OSi1WXXZRZdf/
z32fz7DVk6LfPtXXHSpP741HqnDYZqmPpzn1W/MKbzvBP3Zs3ir10pjCJjHD
jys1ZIA19RM42/+8OGsDHx7rWnRmBmPeYYT2BFuJft4bd/NDjfRGi4DfKivW
rnjaAfNreaM1J3KBtvOMXbyQSuTIiewJyaD+EpOykW7JPooVg93UceZMy/kK
VISunk4l0fWF+9AcAd5iZGtaqSBhUZB/W++Qk0F9F5MJy7SPEZeXmFXLApRL
ViS5HpAYDrj3ltqsiir+RZ+4skozXRp+ftA+7Rp7K1vrXiWlu4o1WEW/RkYR
9kjzpTA10o5jCClGPCL7EfH8H2TEgy+FVr6Cw4kGbmMQhlxzZHPeAtSgmcDK
bK6XtxPUqo8BBuuHtEqmcknflost2pZems3oOgVNIU8Zuiym7yPovZiD1Axs
mUlUIoKHnfpkyhVp9DEqwkL/Rnw2pDxnaJiMRfIlGWa5zTthcIyYh0txH3oa
Hi7fF113UZ5CUBwKB5S8HLA2CpJJg/xC9dhNcJ2AyaGAtOv15p7lBTBo3X3N
As7BfX8e9SRnjyaC9E5iYaViL6TuAD58uqedQ3kNQRadpbkHAoVQ8lsBMlmb
ViBVoqUQjl9+YSQ3IgFvQXf8AGIOBlaWcyKBAgAG88QlnDUKpmAPmu0lS2rp
wU9k/gp1E+UTpait2v7cnzB2ltKtCz88/+Zvrq4bZlRWYL2DZZiAQcTElnjf
VdJG+1BwbGdUbZbxwM5rkwqQT3kbmKE8JDE9urOFR340hrWHQOz8gRJ9pKh4
dSSpOWDHAe3+vhosvkH2Z8yzKqbdg5PxnJ+iqCgabBk7o+zlXWysCvVIAKgE
sC16bcdZahcVIfKIH9bfZxVFSNQ9gElhs2Y2hW+pu9//OnmhglYwmFddCKZj
spWqRN7u1TLbxODdE7QGbwz3dqhkcf6NksZLh123R/AFmrc8Wvstrp0abE2A
3B5BIwIgUZqh27m3EbM8b+Ye+PYhQM3tYoLq6TLbkFGOw7xX8G9g/dEfUoZI
FKXUZJqZgfDNrf335xvCNRP7Kp74RoRf44ejxtkFq6un39HciUEPzFBahJrV
QrWSjk3CYayoc6XBv6eDyIrqoeHwt//bd8Zotzoo0hi6yRiXBrlkOv1ledv5
C596CI+LxFfCV0veEI97Haq+KA+CbbCu34lzeyZX1htEiu1Om6k+hZK/W2nu
TxLjCHc6zIFdqDosjRsqF5NSua23PHIB/0/0BDNZnhV7YVBUGRahF2TzIP2p
fcZmemueIgmXne48wXq4V/vqP+0RvLkgwjJx8UTDa52AM1bj3oxwlLlAvRQA
3pzgyQhfFCHG7JWfyjvfE4W7ths7BJdtwh4hzH6hg6MAzJA5RCPDR/rigWHl
V44pIQH2/OSKO2NzMrr2/otnpdSPsl9DxEc7Ew/Uc9J2SoAG6VuMNdwGQqox
0bCnJVmIpgf3buCIwR6lr7wTZgVt41aIqBf7485vDJKZY2D8etGq2jlPlprw
adXZclkeED2q46QuUN6Bp7+23MrcJ2DQyKUTDov9fhu7iQ3MuCIzinJUhCOE
n2nWNsY3SRZMffFQuc3rfmEE3JpFQJj4UYDrtnZGRQdhhsiH1CHQofF6bNZm
KpScitqyTkNlXci+R8KozcwRJMRodrTQvp5gudxRO8SXIX/uDClmtTuHM/hD
uLhLp1LcTRByzjEIKEMSh0jIJ4zp/rC90z1tNqHMAmuKsks1FyLpsMc3iFgX
8ibPf55rsxcmgGc2JpMqXfix51/Ew9ohIDr6ggKJZUKyoQqeo3kjk83JMCx9
7zv/C25q1qqLloxVs3PRSVOO0OaA7Z3UbAWFdT1gSiKl2i4Hmih3a6M/cz4v
b8idsnqik2rsPi2q/EndGDj1sNsSmVtivJNrkcYa94Xq8LhijOtuHFMkpLPX
6RocfMo35glhlPS6pW3yfB7iDbmFsK0syjNIFGhGQz54QIi49fXG168XCt5r
uWJ8Fe8GA6Fy9phm9iCiXXX5eLXMRbkpaYrWTVnMTqFumev4liEs06xun5SD
mRwHZBLtjEqwMVYp9CuhRw6HJ3diRoZlBUGzkaiaeGQPBbh5Lj7vpbgubfOp
AsePYzgFnLf4hvCZzOklBeLtW/V1V0rLJ9KHd+l7ZPP1jqGhaicPfiWWjKwc
Zzf0ExmuKAd+SlK2Kbqijzh+ivyrgKw6s/SHeg8oFhOUN0f/+6BCl2/JQDDt
eC8UvMAtwzsJzqDnb8APkSnN6SLbSfWeE4IHp4gWa8rYUa2XsVGDFQZjnjX2
1+skDmdlVw0qaG/h8wmtdP3RrUvimPWOOk0LX/lcoq+eiOloKn2wmqCMYpVh
kDE9UI9yW0WOOded8WQEQtJMYUDruLeiHPwkNUwwxcGOBm71PENyfXVHBboK
UYV2iYC/7dlNzE/9TwrWkqwhdTatSDlEg/h5SHJehK59/1w6/cplqZnDYw+3
SKb+9OoHJeT+zgFEYcXHiaAIal+7QBplMXz1+PMC0LtggMH23Oa5voV9Q0VI
UyThaJny19Rn7X4IfjBff61n8bAvY2A4GyfMhmYtrPsAthxiZq/FcWTkLJ/f
FlzpYFE6v02E2U+v8Gsi5Thfboo3qePJ7FPUHT+PRqeLogcN0UFKh+MgASZU
QW162jOqdRrqE7a2Vf6BsPCqIfbI9WlwiaD5qn1gBCnrpY0kKIbjncuMNtuh
Xn+b7CUUrrPONeXrQOcInDjEqNCa1Ng47FzPnd99Z5j+ztDfj4cRr11xIt23
xC8vkXf1kKA0SSRI1Opas5jAFb1znAStMo8GlJXxsyjV7+ntig8HCR2opsoq
QonAtBFlT4CTpGFOcY62OEoQQLINAytEyYZ/EsfscGcfU5+b502KQNomUsyr
Net37YuurOyWElzccpPKOVl731sjvrEFkHth0u3HcaQ6ZvsQaa1rGMolDd2u
7WT284r+Jo1vDBGMPuW2IMVZTNpQDudgsKvQWfZbgtrgZpwHEeReyIDgoVVu
4ocqAb5rgdOkzsE2Q1a3vfVLtNBqWugsTR8Izf53x86euJ/fMSZXl1zYEQTp
H8EguBINEkBTQJ3pRs8qUY4CxoFMJ4zOVwXNL/cZXa2D4khpRRop1VJtCm3Q
D7+cwGGVYXfEld5/OFQIDzdgZjSuuxSVWS+KdBYyS9MD39BucNTkXW4e5JmK
Rd32PErAq/BQ15HFUkOUbGff+9socSQ3DUnJ15Xj9Vvw+L95auqVkzmmCqOf
3JUjSQ1bAk94aSNWXeeE08Wozo8prqh3Wat0yZAvRVoCJE1ZoH4Lw8SjVqGX
/Sw8U+N2mbuisQ4s0R5yhUxEbBxQF82IkhVXXi4xJNsgDo+FQweNKnjY2/T1
u2QwIilNyph8kTTV4H320pAQLjPmnI1cGL2pcDaX5SJGO8ejE7ATxwEgrQAk
xZmhsPloxWJ4jNCz/GDbNdmdGr40tJ4XKU/4e2yHMBiu4CluwTFBCGtAinUE
29QFP9IsupgtDURrdweBPgLsveeKYUQ/7i41mOSV0gVwwEpwlCsONYy9+/JL
oxg6J83tvx5hA9oSbx0vtl5BG9kvcGYG1Yg2nhJsmcDzbXThKu953C2QPFh3
6P+CFi4xv7FN33EKJHepJQieXkU3xIUAJoWw8gfAJnMWCYyiqutPU9nde6P0
0IeAAVy8xPybg+FaExOp4L0+LwGLUVpEUv/gQrHYFTiaiDFL/Zd+cKIsNqp+
Mw7J1xHO7Fny4ajvsgDXaFMe70Ezwa/a9IclkC/Y0fTXtYurQ8nHMX4kK5kN
+YiGEtrydNYMWadQRAdBumA87HHXmiEcnF4/O+f/D5vfaw1mqleILo4//uRJ
JBhrqyMQ8AH4ntXf6Iy5hWnla7aB6vkvNIdeV9qaTexa29oRXDDAjDvxS/z1
SPJDv1UqUwndIOx43TzglY/GeS9JdLDFDugQOTGMVWYEUrxxN/JNL90Rigow
B2J1g6qDwdFAXpoyI5G0hS4e2g45iv4ww8z11Ile4PPdXM45omlwd0n6eJVK
jEso6LWhETxE7mITwY8KA07y1qNig4YIrY+wTevScZE1yCWG5koeC5MJftbe
ir6HsBmvm4BHTo8OFtUFt+fg5rtGN2fFFp6F1u8jqrcS6QChcOZYhSwNb0tN
WU+0tpKjmeXjj+3TB0YUJhN3QxfW2dWNokbjWLdxp9AQX1QohoP3n80s3kYE
oogf7vVmxQ3tArbRcNXYFuWOw4EdGhs6cW1E9oxd1P1ZjWKdzNEKVyrPOPAn
kd1s74y1CZ1htCDXjQ7cPhcbQeS6McrwkoOvwT+w14NMgmEdQ8axThTMy+Q1
x5Ck0JjSXnGjCF0N7EFSE6xvFc11K330VRk7Pp1z0AQgh3jifB/nfs7c7zSi
/s9ARNEtS4NZ2cvxQDQz6zCWWCbTacS5DhLSxHPGs1wXqlnzOwaolRqSvS3B
f2WPRl8C712Dq4a/W0jjMJF5Cv2JtpcxcGVOhLD6P91fokgeWZSDrXkEF8L3
R5dej4hUzlQ4wuShxnYTzvBRGAScWFqLOCK+q/d4PW4nh8l7YiXdqGYi9V4u
Ie0ULZJF2kpgVkRzi1dlQxoBtLKOF/S4+HRNk4ItktVXrYgLrMy/ha9kj0Y3
gSmQiSHoEN1h5OViPRDrYn9qvmXLQjXNWh92RWnF/0sy+q5/fB723vU8SnVJ
yuVtNZA60zWaooGVmAdpQXFGKx3LPcbRRB0qzgMSmVqx/C8Nu2r6vJhbw2Qp
q6Diw2wj20+Do/SPqC160gMXsxEr7RPd6BUvW700T5lYUJ1W0PZOPjgHM6OT
kKsnolfOAjLvVp0eDbvjxmPuae39eW9w0Xt6rfR/f+t88+C1GMtBUDAJ7P7y
Zii9FioOhzFJHDRCHrZmohTawRaVLj2JELl/r/5jbHEQ0jA0H/W7VXjgvOHz
6oqccmuaQRk6ZH0xYMnrwalgL4LRhgNQCGnw4E4/nedBe9ETG0UY6roR/Xui
5BdYIoI8EwG0a+tk5qkjxaw+h4MdNqjf67cSQcdUQgCg+cGeCPvJ7NZV/VhF
FHAooAXdmhUD2g1Ogbz6ZCmmNqgGGJYMFyr/2g15gw+fjpNT/silmvBj7cSz
orwWwSpqMEt8kTwFRWu6iVyUAy727/rMJO73thTAsNZ30wFXEh23ueSIOosi
gxgEpdYIEaOcwQoqv78zlUpGC9SeWJNkAjagZgBUL6gh00dkiSW/ATCk3ssh
vgC6MKs52j/SPckA5XkPwIKpr8dZLVw5IpFHKJS2Z+z85PVF+A7fmNPb1Itb
QNlc7+QoCJM9IKY7brhV4cmwZ82o0vvq9FQGQTRhIoegQiotHOXfeSEh9EFA
GAmj9lq/1PLTjQCROHGNisu6jpNxUvWote5iitqXJ1uV094cSzYZBu7SHSws
0ZEPY76KLlO08gI0pr9wa0VVG6EWvgD4LtvYkjWgZUp4PTFR0hETVgVSS4nZ
3Vw2LzIztJoyjgPgvXHyZulieIVnGAiBFip+HjX7Gwu9RyYjnOn+ypXJPISO
P7o9DHYDbWAiUOCC0uFUykZHjdDD0wb/5UzXX/YCQC0Eu7yhnHeZkk94Y+IA
h+vA6eza1Aaz46fof2ZWF7aKQe7Oq4VfJ+IYvAArOcMfco/3ghzI9Oq2/EPP
ZorMb11UX3FFFDGGDqpy8Ncy5vodK6n2JzndNm6zX5wz6pcJsB98j+L4+as5
WemnQ850e7YAJcv7OJFNvQRfY4Xn+Fsojg8XXUIefStJoJ9LFP2HZUjrMXCQ
HllGgv1WBqCYSIyAS7vSCw3voBk8Luuxr2xSuBOmo3Zxj43l1aMpQPHKrXx8
UECDDXkJs5JImX3eIA89nrJVZmfJquTwF8fsNmIBlJSnuCkMYpFJ6Qwpg/WY
CtkrHSc8PPazccMdrw+iB+GlisijIGMoCQQAETlSkf2x0ukYbSAl3+5qD1D9
1NnsjKgqir1l6NmsYCvLr3j++XfkrojY8zYKK0dNVLzLZeC23zaNsk94wRc/
auFWQ6JG3H7R5dWSCzvvFdIlGKuJ/OeJVhtnkH1eu+OUSqYHRUvJz8xJ9u+E
PkWvTJVYECfuBXMjHTUdxJHojhP6dlHy/wIfhzXr+V2hkL99WGBI07Tu7Bvd
ibcjW6LVgR0pCLIqaF1a0k5oSe73vAy4PyM8SJdGSgSP7h3V9A4FOZmX4DKe
iJE7tA/2Llt7gUUqMS/gzaFne8KRkURz5eBQ6c8BI2JJApwmnyQKzxXMND3o
/vmS3y/e9A3tihXNHxTrPX2O5SHtUURfRsZGmQfTmGoabGFc8IgiDS8rmjpL
MNQvidWj89q1n0EYYQ8cgNmBP9l6M3gVXAU8cGBz1vAz5DHxrnMbpDyOAQax
roqUfiiDHU3Xnts1LJI5Nw/h/zyjXluuGcJY+IhX5Xr6hD62VU9275PYc/tS
MXSWmFE56K15Ow/67zV+w64tYwqEBLnQ4dj5RKckTcKf14+rbt14BwOtZWIH
syzM/F2e59CJBMDX4C3EEwpF16ZKEQaU5sLGjctIXK7Ozigwz70XEIekV9GL
TJjiKqsp9P6S4+Es5jK06daTGFtt33rylCD1OrdZ+CIOrbgxilSY/vLegeDA
QWllE6pvBMfWabtMeRwwvnegT7vpzssLt6eZlow5H+d9b4gugcz2ht1wQgCb
l76fc53yv1texrvmpwcc9Q3fszvqeBNWmxeTSShezCwlMmeBpGF+gRMvoF9F
8uRrjQRcOmo6MSwhvgu30fhuF3wELb0UNmzKJDkE4p73zSdu6YveWYPV5wcj
dTwCMwBKZd+8J1IzTNAIFBVv/+EB6zAF8uWx6MRHKY0IZK8phGABB1A05HPR
X1/gw7pp3TmsjLH7DwixpIieFOn9YF1fNeBREjw8G3PtY/vpC40WqlcMVGnh
zU363TXBnKTNGU9fWkwhSqDNdKCHCiGRpgGGSh5wzNRSwgyQcx4KR4yl6McO
uyewK1z+xDmMnLGyowyFbAuRd0dI+iqm9H8k0EOKbaEQkLBMEcrrPYNz269d
9L9xB/EdZFiHK5x6R1/3tD0y7rnqE5TMAeVInKSYVSnrd3UwosCTzDQB9mHi
UMFZC1W+UVfRbUA8UGJkZkeAoKvKyJlgBfYiucpvY25v1o4/ziS6HmjVlHAm
Qp7tWxpiRWMH3yv+cnnUHOG9TCBJ9K4W71leEtL0iJU8etFCa6lfCTjuH9Kh
CRoTPELNVJ+NFbI36FIXbWDmw4maGMTnU4QdPz9OFDvHW25Aumd2VDpT3ja6
j/uim3eYOxSo+KD5irQqRdqpRC7ncUTrlxwLEG981uG7L0zbOqYrbYQg0K5U
Li/RbiL9jmxYcPbOEwhw08NFve6dXoU6yFRkoGEGJezi6uWgGVUD89Q74Ejk
TSVkh4HzftOzyddapEi0ol1DgTpfKCnsWUe5CsXS95bzsC28Q6fIIQQhUSAF
yIlaPXRya9wbjBvPucnU1l1l/BOCq16mOmicrvuCpKxsmaXx92QqwtA7Orai
Lft0DIPpUC97LMVzaw4n4o0R0yg1NB3ZOUg3JPJqy1Y2stwKAjeyAlsd5LCQ
LAyGFOthBV3nowj31QVm8MV6ThraEutIauwepS6ALH9ToUd3yVEkU1mlKAIY
3tS5NX6oEz3bZzxHuLstE3aAeI4cfJfU7BfVEV1mpPth7vFayKa7sg+R4aFA
6wpS0qa+vBEKP7/hatXy6DpPVnnU18Kmgu9Vxoa0qAFsslZ6oIgtdY6N+wOx
XcahaACzUfRHYS2wJhT62vbR0cPrw7NNfOHot0WQfRPew4QA4c4RQVHH6JFm
PPI6shftMb88VehAfE67Q6EYc3BavGet4nYzfsQ2Fbca/N3uVQ7jHxg7eWzv
Z6CQ/Vwj7wtq+7ydi2Wnjkw+3UbVUBIAH3kbKzwoN3X0bgKjKc0gcBM8nnLB
+M4Q6iUdCuTxZhzWimzvKTQlvrQDXETv00dUsaRsVLhQP6ZcgoTrfn8jUo94
Xl0SUlBTqCmuhPKF6ZrriegvKqRqmnvyo8unXIlaYlSkvEe/lKV/YvOTDB1/
RiS271PpZtB05nO/dyfMMARkrIQHbqF/B+98xnzf7JbXgCqdXb5sLeWj0vMZ
/YDlhkOZiZJFXzxPA5m3GUkJrN1WH5ucfV17bufqL62Cm62vhNvHqBq3/owF
RJk1mYxij4EMldNi92u04Z3h1UNp38o0seCxwrFqKZxUbfSSx2f1qtYyJnmf
64auRbMTXRHkEoSCRhl50OkToGby6rAdH833hRXozfbF4F91mckfRWXfIoei
rYyz1az5FzDdiau4kf/fRfBg61saznKdnMBC6m+md+F34HBN6GNlJHmavtkX
q2X9Sky+B4YjP+kqU9gP1TD6QbeyVOAL/feR1HR9jl9HGM2+HwKwtXOmPXsm
S/2o1xB2pJeJodwCyv8E7+KxZq2UvSKkciUu8V9vDpx/umboKmK8uM3JHg0Z
6uZmpa39FXBKcRwE4/4XLcpg7kGWpOU43vo3sICHD2MF62tMT4GkgQS1mfXW
iut0nuWLFQZ+l+Zb/wBHNx1R/Z2aJLpiDbpAQUbStmQFRE3/6cJBzmjtFMOR
cmLILbJOStq9ywiJC5aXE9WEh977ID5tcoRewyx6JnNVcLWdNI6jICE+eb/W
GHAhV8UIlwqgkY38LK0FSHiPFn5cHbxQvQpdqZ2/aCrFiDMD70HgbgA7WiJV
TGVgnqE6hyKwZziKUh6Noi5yy6VTrV6Fup3nUWk/x6g68D10TkzXDN+/sF+Q
vZNn2lI0vmtCeKNu5j4Dq2NVAY830821pTpOVjvUNdiGtKVXwYtMS81X84Lq
E89NqkbwqPEPNDraF11sr9J/lT3ezDVVgkVbS36fOQ7KFs54OyYKRpnrKM2+
QF/nrqk3XxvYEixy1xEPQwNEYqqCX6u2lbJQMlvn+RLspMbj96rxG9CKGC+Q
Kio+XJBvuNr41uuE4sXMrtneXtNSZfW0J30vn50PPvRlx740uF1UO3vsBG2Q
D3BoeI/C2+EM13R0JqEVB2trwH3x0cVboaj3X+nVnPncqhTW10y0ArGM4lDw
jC6UoIBR7ZjyzNGVno5cjQuWa4Eb9JFN8aDKgEFLmpGhMLjLyq3FC8r+q07P
stjGDQfdxUItpsrdtvUdlw1SMTFKmqYDvWNOoBFR91RkdPvjZafurEmHx9fl
1RyLf33u/PcSIDNLvBevdVZUiX3+jO/HB2cv/1yFbkMxRbH9sFi1UqRTjbEP
q3HdYJ4JTsbiVxQCoXsORJNWq775a7AUMYdw/ILBENtXktiLbF4naUiBYpXP
F8sTgHX1M1J1FvVrCbq7924jK550ZkEdnrEg0h4770+sVhVJscUIy78thBtq
okJsK/slvBYTf9ro2sbS6KUojdr4wOUTEB7AOxjoufuM0p5SettTtqxUeDUV
vr4eExi5t6eUDTeStHeA7ztWgNHlJAfkZN2vxQPiX3r/myVHiPKpCHpKEGeO
4sb3SraOUzOqM1YPbHqn9qZc9IzT4qMFIXMPiOLYwky1Zqo84iOBR3gByxRQ
FCAkfe4bKUtVrX71Z80gzEPcdlmrZ51T+2f4zdDyQtkR6MoEVuYRc47AmcQu
0S965D5ckFozSIQZ2yuwMM5fcNfNgEU0LTGiqUr9SWt7qZakAGUE+U6+QpSM
6eJCmqDChuuFORqo6u4K+jiA0OncRIJyqcYLLtk40DXNJ1wxGSsr9lcKhlRw
tcSmKcf/++T6RuBRQQ9CUoh+N6OkjmBa0hDH5d8fXQzQxSK8BziX7/lmzQBV
j6sJbvbV8uYI/8JdVm/3gp55nBmIdzlOxbRa6AIXOGaysgQIBE9fsqt07e1X
KZIce3b599mL6PJlmNod9+U3VHJvsD1+e8acBlUMPRnfk0yliFFdRfPzV6Kz
Xl8xbx8vStfXRk+5UeEhWXuz3mCIlaAnLZf11iKo18aoHygrgJsDIUtv0S54
9t2w8lq6MwDZ61Q9EayTvWKtIs/TyBreEZzFZtc4CyWN8FaDmaTOgbrgIS2l
w1bVYeN8WzE7ltdTFA//ASSjyA8/GWtWqIdrxASqIiTBHYMc+SmSFLt+Xiag
mmC0qsudjan3qoy8IuDfKSIrFDSNK2XxJ6pbX1/AT1uqHuy8RKk3HhhaldMR
a5ZecnwFmq5CyxGO+yFxHE/wcdYpGl7C0H6vB7tk0j8qLoSvSAoqKZ6XRChN
oDk3Oyt9nnGhkobucrezKtQXfos2YyWduNcPcdGIo635nuZlVVrHD+J3+8Jx
G8AGh1MwAHWpZ4CaiHfK+sP0Sv9FPGfGWyvbHzugpYBgy8BtEH0xa0PalS+g
gdhT+kexd9Vxyt2g6ujK4F/L5zjnG1MOkRmcnysx8PDkqf7hn0lVyRXDIK1B
dYVjKkm/HwonUirM/RW1/tIY2otuQO9uY4Kbx/h1nhNgSvCGk9M9TG94uqTL
7jMoWAkwzYn2oD0fZJKl2mk0etcKXfLgiFYITIK+bkqmf9ADvJ31vaK1gNxq
tJkr+ZD2W3c5cw8Mth+vf8VWZ/+OeB0zzlyclD7BS++D1eq6JlxwRO0UcwlN
25HyHVVXZCtWBMKimaCpVFsiIERNpkkQcx6pux4/23AB/lKmZRGJvqvqBAxg
GGD9YQICg+PA/Q1Dvud4Y7DsMtHmxoY9qAUeyRmDDZ3lqiPxDz58tazjEVZa
efDYjfYAeMFZrENQoXlmeRQM+uV/AaV7pH1yN+JQhUfyeVxuemEpEqMMf/tP
UF+hQi9+xLyAOTgKF+kqnIKsbc22If+2l5q3ZkD06t2c1JoBsc7+iAplq2G9
s7GZ9ODuUlvV4lRzmqkGTfL6vdR/NtNQo0C+jL5626B8cSQ82AkdZpteSYJd
nPATMOR7T/PHV3Rs8RWCEWwhTt99ldbJnJ5lRRlQE+H1dpA4Nbi+P3VFmOxK
1/F/86csOXfvnJqJYH01LWxSZrudelPDggHS/B0+nSMEuaBeyfVSMfY8bOnf
ITCpyXGSVjZZB/6WcX/so2OQ2UC1gc82JLyE+uZvuzyRzVgV1zuUK4tHBL9D
xvPDrABNN28s13atH8DaXyhcvPpho/yiBKQHfDcyavT3/U+KDMGryWyISnOA
hYofj9w0ehu0nRAXPR91gNlCYRkjL8avotSkf/SiEEgPUralolFKV+G3hBOP
vzaVA/epxE51UjuDidhqJfsVcxJSh6yILiiA5K8YRC/MW9G24r62JzQkprPB
q/fLUkwGPY/KUT842Xt53qG8rR7U+4Tz7yZL6voBeMbEdHQEQlzv5hPkJqbS
fW5T3ujH87+KBYxr1aSoIr6V1b54tptiS+07oPWzK9VIw9mfH5msukjvv3iC
jYpdaVKz9H4E3RLBEkVGm+UsBDq83aSD55LcVxj2Lb5u/GGY0qft0wwpsM4B
+dBk1JlL/sr14o6snakyI3GboeFfa4UlFI8D1xbgfna5YG2VaurilnYDxwEx
wog9ohm/4GIwvPirtxpYYSh+RU0GrmCFpPX8j8TfpTXSvgh36VDDnX+rXX/N
w0oJtAejtFCgTRgvKucD+UGqSmMtbbxW6bo8yrW5+mdfhB9eFhzUQz85uYqL
KagQe0C2HZuoDot+fTNucbWKK2RfPvDh9VbcrOQWCc/NxA0+cYzAfztnkXci
rL5mg7s9a+VNcP5CMff+kCj8H46fhI1EatVQIVAZfQG+XWK7CDxdBJB7eZRz
+wu6OtNeyclotNPh4zh2oOkdm9B9DOne/jOrh2qiP4dFldsUKsCMoSmC1HGo
pVIRlXP1XuRrBKrCULb9Ar8WonX595bqyRNUNuZ62tL4lWpSydr/9zsa+FzB
s/9EKcv7lSxSk+4WrXscE/8KoOR92VozqzJrD6MkPQxZhPrBMB3d/LUk91yD
g5dJbtWBKmd7Dz9fdKKsm+DW/toWdHqrtkU5S5uOc/An54AE719rtRaYuSsp
2FWr2itx1n+Qs/8KOp/VvTb6mKspPIazXwDLPtODxajeT3UUznPurgfM1RKt
A34ayZhrUuyM46+MlIRKXeklziFgwc7pOM2E8uihTSZfWYMJY1S4dZ+mI8db
5nGKV9gVGURyFP3RFAfk9/ehd7nTlnKFL9uCicVrpVsbuKFbNUXdXjdTAM4U
7vXByjLm6nIpkthA8L+6KOL8Vrz8fmEd3WwH0jEEqAW9y5ckcGCFhcQQyWg+
HgbEct33BbRxjBafcZ6ItCcG7WUAcKzk2YXMzY+91z9NSCKJOqTTL7EycqYA
8RqQKHSTYrHULZB91Yr1dX0UY2XWRwXBkQRfsqLg1HSkv/pDCipFKFFBGgLo
1kVCa7QHVA86Uadt6z118QshIRxtXzdtN+M0uCXa4eWxzkHKuOXeMYQzTjcx
RZ8WGGvdt8+zzppm0yGQZTfRnLhXa2+37jKN+N37Q53AtHakke9UZoOEXowa
5H83MDkk+HEKCl6uNy5DuIK6OPRKHG6HDdpHrp/8o9MAsnQ7RKQulUkPKXiR
gEBC9CKmR6/+/fHImh1G147/IcsAxIGkMbAMbT/ZdEJ2BXGUuoASK+EjeI8k
VL0dEQq8crJNtMSIY38NNtHEQl7nLJF/Trmtbsfw/PESVaBmp77sxqQDV9dX
EdhYdaT0DDsZKqPV0MOhdZMI4fc93AlVNWTsFdfpiedEHLCb83ot5fcKx4cM
q/SRPGSFcHq9WM1lNUJw4zTzsF/jnDDiCoOE/Mr2/xdAAzKtFMVPlKW+YLuh
M+GK1EJlbyoqHYKhRW7N21UrN4vLXEprANn5/rIlMB24myQKWG3DLH4sJGFB
puXb5sw8XTaLFyUiPANLRN+uFZtW/pj9jvO4ZsfJnj0B+vA7MX9lPKExG/VK
ZQkXKze0Cv4gxfN4qNT5YLdeJJcxJnD8+oDVmGd32BC+h6dhMlF6EoQ5z9tc
kW/T+K4xLfOXmJW7cc9pNYRpt0WWZCbCzqVzwX8TmyHsD2psCTzgaDQ/KRbQ
dxGCxoE2zU+claTCcb9JQuvztH+3SCPesj4/9n3vYZZa0BZndHYWZl39GbZL
7IX//K15Et7Ow+O9CKGX0jjlYsibMH6uWga9xJByGjqISKTj+C8XGwfzR4mZ
YyuCMcsFIkQk2+OnlABArq97/TdVGkioYPAX4ZrRMG0K9etG7FrWTrqTneJR
o9Lc+tRqMn218TB76wzSA2LEzyIlXAerhSWrCH3h0zyle6QFfOoWzkO85Jh4
SZti+02MVdYCMrY8Aih4abTAfNaxi3QCmCR66kcYQ2gnv72P3hueWU7MOcs+
sG6Po4xKcXuX3trysFsINsC1dlVLFwoGsy1B9syxcxZSpfs3PTJbvqKNBC9d
FnVaAoDRcsSz4y19NClBZPnme/6rhPE85EWjGkcRF9diikkZEW3Q8jREcZHD
j7jIM/jN9+1moayw+TI1w+h1XkMppTRK70SGo8g2bCWWzH+BrPMxWpCQ4NY0
AMTxAGbRA2HhLmOlW4ir8pU0Y4GZ3S03uI/TZA28NXD4V0x4IcrTBgh6eH7j
jtgkfgyv+jMNNrLVWighlSNpUAFlVTVnvEHyWbHEtQL3roXc4OolPuqxcIk6
tItppaHOq1sk4WGb2PjlD+iQb8u3d/2/QshzUpPlnozDrErTYC0N1shMutUP
Zd8ZeZyfGtqKYpAiZqfz6fId5DsNdqu2UFPdsmMDV63xGbThjwGb5X2Mwcwl
I1w+lRYzaJWcXkc5xTXfaWZxAPbohUm4PD1ZJ/QcIm0EAOSMfHfpYcbkmE2W
UH1k6rEtM05zwPyfKmf+PESIZVnotlSUI97Iy3SbV4WN+9iQIunNU6hrnudT
1+juxbYYF1srnndvECxx1sN2OLHDDbHeePexPjar3CsdoMgKAcNUBnz5uC8Y
d/Q6YpZV8mWy93rgikxXSxhwXFpK+M2zJmHnyjDk8D+NzBKIWDrDIJ3HD5GE
N/B7wCPxWj/dYuSiBqNOa3GGfWDGQyiAUV/RSsNqSxBZOq34tgbvUKexbaA9
g/QPJD/lypNrusSKb4RwT04RNd4IHTXI2Mld+YZjgelfRBMRLFAa+KHnlYTl
OxYOObVwA0yA2wq6RMnlC0Ir+KDnwO9XdQ1ezZVV39bUmADr3MIVxaDJDcc1
MSttSf+6XHL5C+kISnoCyoB3BTf4tIyd6wy62t4cOSSAm3qIAsXefaEhSAK/
Q0i4llzByh1uYL7HzBeZhL8h/eeQgW6qECNrT1wOtq/mj/20l5uWuUgrGnG1
v0o2Xl76pXW3HJXc/tIU61KoqcQtYs4YaJxR8iqKQrUFC4eVHjdfT/INYTKO
pBe9svvWuLwIZeoDdfAgxx9T/IPBH19KQDhjC9dFYKvson68MWfiX3P2NVwg
4wdDqsfa1YHqx8esIM7QuVWMT+QitMfVRCaEiEk3AafOvUINNWQ3McwNvEJN
uLvwjlWS4fTSKh4b2drsZfCFlUnUhAg7mKZlKU15PZjGAgqxhBUH1c3hFmeL
VvaxvzE9OBR9FUcGi8qkMzCvDB7Iz5T8Nqq0hfMC3J4Ow8g4jn5y499CdhMu
ItQsCxJaS7X5ZMXnox3qN2rZJJK9gFWiWUUu9CpNlG98qmS39zCtqC/1QCmn
QwLsUrNtgngB02Lf8Du8N/ABfsqwem+AeHMMyRuaHVeGk36D6rhvPfbrr5Tu
91Cz1P6OaDwHrXJn558+Tv6UwnnbdgF6q5I+ljDkgh7Kbe0IHo0sjH8mnF1Y
/E3ietuC7FRE/vRuW6EFJD2nUcyw5anuMBju2l/mkO3VtaghLGgvXgIxJvCo
iiAot4iNsWkNzkCK2tpQ7SUODiu4o2C41f5s6RJ44UyYjDLn3NqMwC8d1EoL
iqrWIAOuECAes353ZIQHjga9j05QltxQFfBPjch/jwrHdxIm0q9VikH+NcZD
sSSv8maH7zP51TppPKBq5810d0aVZLIeHHbJD2IbC5ibaD78PM+cNV5LHGHi
RaCcpRcroM7ANkWvCJ0ys5OKPx1HvK8cCUYrh0vcOaBO/2qIi1PEjpKsWSSo
2zyiF315D34dR/ytp5pekik5X/md75uXIlxTY5YILQQx8NFfMfLqrgxqLp7Q
0lmq/od9GtrppvB5BAXyDdcMYCYleeuh2J2OT223FIYGDgu94BmBykXCx4ok
YQ6CCGdaKP497xz/GuUJmBNqtEEVJlPYv4gG9hVnTn+WjSojgk5aLneut3AP
I7mL3Z3A37SaPlxFxe71I5hO9/E98QwYiDBjMCwstFW26nvl+ZITGWLpm8ag
/RE3ppEGL398tmVmuzjxpJidcJVOPqhgVn9f/75K9m1SrQyio1BRqaJJ4Uzj
TEa+DkaH/p1BqZbNnougxDGKqpYtiqsdyZjoIFK57pA2Ms5Juzmf2tRIGfqI
h4nkm33Q9FMO5TV6OPa7IYb/fDL3jtT7GyMjpSGi4SK11aPvO2PVxyKc/SQS
HkpjPPiFNHKtxZDBVMpu2x0nkfOAZZOOoqMwtDzwWktVyUt1/hwmcc8lvsFB
wXZw/QvVpZp3bxVPh6w6mGeeFD+p/EZu4NL3Wq4hf2ndKF0SMgXyUfgeUgtc
rHpkAJlgXJRD8Et0VrQnReZN2orqC4wlux6hp2iwgT7xE5nUxTd/VkdsJPBs
Duok2E8i4QYQV+985C4Yw8gUdObhOHzp3V53w9fNnBhPjTxQzssWZ3tL4EBf
JVS8OXGPZFOylos+WzBcihGdALwDRKPeJGJvUYbHwsc1pmjTP5XJaTOZCMHj
e8Qm6fd3lZ1k/Bxm145DgUJKYNzLITz0cQQVZRm6oQvGomBmbLQIFe2qI1V1
XQAaUI0KcUGm8CuZ41fChvFhvaI168DTcjpKQYtwWgiTIsplv6yXZEeesiDz
nHumD5WvQOib1pRxIXrFvD3br01uflW03JEfSUEbBfs2Y0D/afRszldmnPyG
sao+oII5UUWkLhTPynplwGZjxh/rtTHvcY35Hs0AajzBHInIghW8Fny0WF+D
Ya/XevgDSFyTRnvwY7phN03aCzmjYZOsVCWCqAf/LgoVkQvbRAvKK/zQgJKt
4DqnFEHx+spivZDmqkhWX9c9y1qmjyxN6ce5Y5qtH9JvtGzQdUVZmOtSgLVy
3IveK9P/q0c2aR+nydPXgMK1zTVFIkl5GBxXN6aaxVP+1IYv34rpeFpYIs+H
P1GKRelzPf1kepan4GgQnNdO/WIcfhij1IM4bbz937zaARVaE721kIAvaaeU
UsRB0+CPhpYRMOtBkUUXIt8W+9/4LkjW141GE+0gpvIR+WJ2UKpHmMMqOhIK
ANkSfN93B+quVm37Edl5lpAV+RYAzF51pOOKF0RHbfi9vyQMzirLGJmzBphz
kEKpX+mm2FiJ5CYLyyilPpAX7kDiOC35TLpx+W5UKcCIotlwa3iUN9JvJvGS
SYYQOZqn7/qH2tGdnFXyLp+YFGaqAVJs/w7F7sxBDhalHMZ9UyCbXgzYCHLX
Y7ya4xlWuXiPHMPIzqEzsgwQv9db27KM04EaOfbIKxdzprsQg0m1NwsC9HFA
0lXGLpJ0JIiV5y2fSxTiMNXmDW4ru+76UPx06/KoTLFSqj3DvBP1Wco+z6NR
gTdSO13+7oj/kA2zqRgE4i7mOaouz6tHclbXVuitre7NcpbsG7zFCwBsu5W/
Jqs5Sh+muF7fU8w3knz4zzpWcdF9HjXN+6DTAB/NDiNUISUfiRU36yRjjfcF
Kd1OywfgxqwIoDocn3rHeSjdjVELg0/ixefN/vz1LPJKZCPI5LqwsJtu/fCw
MPiapUP6oQbYjMm53CamH9dqLCwU20Nteq2Dn42TNFLYNAju6Yj9Stmib63A
lFZwNLUtlSG9Ozy7fYyNKnfqaUvQlq4ekMOBoWf8fylJCkYJhxfG18FLxNmk
pDHC6JAX8LNuvanSJ0eOSD6UXHsMgZ9Ohl4kubVsLG7kNlKwPFE7gZGNRJ/w
bLw9FUTnMVrKlc1723tMBH25nblWroRvGir2hpetkmJqmx4b5Btj8vQAtixD
D54UHBJ7YmcKM9bqzVVzGMsO2r9GA66VmIzJpn2K6puvwtnsZb40gX4jiRCS
9rcjKCnGd3+9I2K5iDR+k1UpY8Gut0maMoQxwor14aT3cd8u/GlHGtpm2LhE
dmROijSuMjXJNcc+Tp+TO6x98BTmaYGLUj4/3ZQZnIPo+RC0gncLurAufjks
IV/mhh+tG1EBBp0gHQLNyngYca2Rf2lndT3mrkH3E3k3Td9vfR3PIjqVJuMT
nL7orDu2VLht/8knkq8n2yRa8Y735xAFPmf5oAEl4n2ERNHOoaXp87eI/iHv
lZ4SQgtzqHQlATmXIKo7fE3gkxAe0hXGb74hPe1KKTQrVK20QUsytwndQ1CM
CE7qN58uXKyuhSq2SIgUlSOhTMzQVdqqY7qQNVp1BF9nP1pn9bY7dzM+oIjl
yMTK1gPQxqv4k/2Q6iha2d3BoKa+bT5LC5ebKJbJV7lRCsUPuBa74xN2N1K4
6sTTzK/FXn5pBDOlxd7+eizYUpmKiloG5GsjrcQdFsam0DOpzXgRrDlMdOvT
G8zUlgLMi3awAegQtea9LD/9dedoCi2/u+eH3ol1D/HijG5Snm9W4I0EBmbq
QhKrkX1bp128gjWKwfjfAcqUddBxvxLr6UNu3Lw3dzSf5TFvej9tMx1I9pk9
VoyaO+p1ocN0UvmWIRyxs/QmaYYxHZGd6fRbBQGGVCjkZTMbeFKhC23DVV2P
tddRJ0MNK2jX6psVd8PveOXkvvWGmU4lWCqRTuHelYNo4oNQg7tPtyhfYiSy
xoPLzkodCXWGNuUjbzEAwGHBsplTcYO8TwkTzWg62g9hRya3wlfdlM0OF04J
KJO9NCLfdsurgUCZNk1VeAisfoTweSSKorSdx849niRYZnk/EE32dSNYPgof
fdnew4S+r16Obk/rdyMuTOV6Vtacfqb30wDL1qvFbYeFVPrRc82S0QZWMeE1
1Iv+sQnO6AZ3mhbWB6sZGjMQb7r6NZlI/+xN8Ha0tQbFCqGK50S6kCnLtlWY
MVroCIt/nqEPkPLWe7qwfl8vGRm4hMTJqW1+Une1cB0QsgtLqyNUAnsyoYt+
VJaKeVfGPlcKek/icmJavc1vT25416U6Aj1DezBeia5F70YpY3j3ne/ld+7y
awg1eMiHWkCSLAVuU51OWXsMQMYMEhA3za1+cRJHdudGGZ8OI8NJKFUtONcn
QSwDPhjA1ZQbHnG7OYZ0/4qqBlC8kUkRMlhIKsi8ETlOI6l2E6oOAxh0D8WE
zy2Vc3KR2cQx6gpUBPJ/oLY2p+ofHI+2zvEaV1wqCLyXYAAlVS22rUo3xf1U
vqz3eShFP4al1UPYICZz1d/BHOco7BFXNiFWAsba1kQ9bs/w8IqlmKwv//e4
iHsn17cykL5ygv3wtwLBKRbeBgdge7f0J9aFJnx40BRcrk/0ELJWQCr/tRSW
dpG/oyX2fgcgw2WxiSvghST0QaDr+rv8ZbIKyhH8YQ8b02W+L13QI/egA4cj
OMDw8PdpJI4KPAFbXeazN7pQKDe3jaDuTcuV76mjxQrC7h0vxYqY0Wkvm8R7
p8zYx6Ddyv90mPf7mpFukxeFPKKk7x/uqPe4LC5C/NAsnYWl8m4MVtE4BCAd
3KFzqx6Lj8M1RFwfumPxMPKt8fb+d6I9Ank+sTTO8Ixw+IcGpa4IwyPzhEcb
CoUlGkYpItl3BX84aO5rx1PYWwVrfo+rHJQMbtihpPq2DzFhVP3HZzxquxm3
ucfHY+Xl3nf8SQMZBvnpkojCohx/0ueky9ldyDxhzcAB78UlqH0FFYqBUY+b
B7/jriV9lH+OTg0dcaVti/QIOSfhqsF2dCXbnTotmK5cHl5/9H3qHCFE0q/i
ROu4EtACXNdqxlO6LbHLuOtZ6Kag3iJbKugksgFwTIs2QrL8Tf/IRA5OA1yQ
ssZepgDhVUrLVmMwHjiU+ARZcvHhaonDFnpoU39h5eD9DUimjoHG4/PQdi77
eQRBYrj1Df3+MtK/TgkrqnJeUmE8jK5n4nJZ8mqQeQEbfzkdJVE0MGo6SKnq
jpZiAVL0dTR0bKzGOSif9EWyoK5DqrOpDaFNwL3JCs3uAEUoWDDtxvVJDVCk
xbrbNBKEWHGFyTADrbvRePm47hemyInCRZnnkXOvQfycSOxM3EPPND8/5bHb
WDXGyZlnEs0emksFbc66gFzBdVv3dPGhzI3m0Ljrr0dw14Jp9LnOL9xu8VC/
9jinyDQQtoIGKLkp5RjZcPcru8J8mNl2g8NZIzJrIWZAftkp+sMdgMte/ykQ
JO/zWoAe/hRpQWI0d6TtIuwVGn/6moPKShTBlLOIfww9E6/yd2vqgYD295AI
S/IO0PhHpp6c257Unx9+NeNCsSab89ndai8Mu5sfW/rA5VtCQvjnbFlewefS
Wc4qgx4yPi/qVeShkQQmqPPTMnfmG9Njq4hkRBl4J3wU1QfFh5E9oPYUGE4Y
y7WvvmZi+dnly9VNr/gZ/icl2oEk/nwEjtpfcSMHjskx/SinUPUJTarKqVrW
jMqrP8cLAglxS4QsbDx9v58LJMhg0JEo7p7lHR+4m1Yq3SaHDt9fJOJ8+fXN
w0kj2Zhk6RKh+DfwlqcAH6zi0FHUWDAXE9jaKv1uCjw2/hD3qy7N5U5DG2Q6
8MZ/m8fC7rcOx3z4BhxOSuf5+WUM/SmUgbmgWP8RLJOqwAG9NQZOvNPRVw2k
fb8Ncyzx6jpsyclzpX0PyhGmbdgHemorxMHj7OLqwsVRGKhuyGa2V9QWRA/I
DCjqQKEWil/qgUvXyGDfH3e3YUkeWK7iVdaXvOjGKngExVxqjr3z5niA6ZHf
W1QiPMlMujXtax8yNljNxiuVYDZbCtv5Ox26G+BN/7uHOczcC+ILjZh8H0Ed
nLvu3UN7pRXwmMhSQFZc6RzfERIOSMaKrL08SbwBUvS/Cm/0nWb4No2yPtGR
MjJ8Rtwl44wRLXNi6vw7LtpT8r6bbRdRNHzFFHmoibmbea8S9ENLCRVYKC0i
r1qKwwbqDnVmB0kTY6IevHK864lOjedrexO7ZpHaijJW/lkGHfISmCqZPxLT
gmS9fNBkWwkMLv09fMS/MvYpe5DSe4xXpneJtuInw8IApWieytIYngf9ugmW
x2jqn1nMJuzBA9ZEVRToNJ23V1JCAJ9eiq+NdUzirdNasD7fnTXBYtbNDl57
jYQLoueDBHits78hHQiWC/lQJwwXYkMeOtIQ9zwvbzfuNY7nifEPcgAhWXLc
QYA/QAuGhyx66UfIhGpMIIgKbnGmnU2yKibVWnzY4Z4QyLI0rNSC4gBpkWLo
al0vshaDL5XTtWc5cFP0eBCbBwDtPuFLZBQkgEybyITleqv2fwyU/C0yVXch
bHciMdXRP0z4NwFvQ6asXBd73tGwAjjqDE5FajqKGb9LEIe3WtYxwDZiBgjW
DAtoBU4NjKnf8vOb71CZ3uU8V2av8fPlKAf9LQRJdyZAWfni7d1Dx8dq9LdY
Cj1KToSEFU5/3ggkbZCvC/FE6c5h/cdz2SkBYAiQA6dvEz/4Ar7IX0gCdgz6
yumsBul+HgoGanVTxMLSoQwIo5u9shyzcp80o+8J8kB8GXyPvZUugPRk3jdU
ynL8eV7Immlz2OxZD5UKzyJ5O9WKBs483NUeNQTI2dLlW0wJgLksIokxkuVa
eAoNXsh56tSoHheAgfCHPdXgqlGEaoSgyxRGRXEIVLYo7oylwXFT2nDHS7JT
4l8J5+z3ahv6HQekLi0rscWNdSIeHJ0qfs4w9sektEyXZQ2fS6+VxGsBF3Dp
zvvS4xMHCxYXssmWegevqhS5olcg+dfXqmKhU70zYUd4q/10GVaZbWxg0ilE
tKjGPOBCcwAqlI73gBX111rvGQ45HeJttBvOzAHojxcMnlAaqwC8eNGP06hG
Xmdnv+wlLz6/bxNjlPfNKYrijZDiEtkbPZnGZ0/s+R3jVL/mERpEkBZ1tGnU
M5PSkZcqBn8p03DzxGnsSFbhtw4H3N7O8N1wpdU+jnYd5Iv2dhH3XFl2C2Xg
OzBHrtPo5si+rbamGH+XyqeZLFWQyog1XCTC+AM9ezifEkK4FN5EtJ4/G0kj
QiTlddH6O5F84+ONVF3czWnzh5QpdaYUPWI4RTSV0/PcBTJ/efdLyGWN7doB
3TtlsZAnBXKzEvN0RXPcs+38Tg98OmInLnu6WPKg7I2AHpwOA4lFuiwgWjJc
SFK2SfhQ0kTIHBTJnidq7P5UN2b7vwhkyCt9eGOpA9yBIh4MW7yhdCsEoaUk
yH0ZAJG6jSDQCmOmuvW88oUXNhV2DdFQRG/nWRYXwRsmJSaNLMuU+vsJ2R/n
AMv7lKZnn3XoCepRkL5ElIz0HS1JDjdvMdDtQ19TeIIpGaxdDYAEo78KH0tJ
Gypt4fhcKPH6vnIYgw4531BS/0SFJ/jLa/Qcv94/wvXbizKlemynOivHjPwV
Wb6Q0ne9z/1nPQfn0kWhtEjpUmTjbVJsEju1/2ZoUY3NPDFP8WFu0c9vnZWw
NKpxy9o4OvP+QdyM63+e2R4Tl4I1hQDeFQ43vvylQ7zt7RDX4Dcv44iKmHFi
Il1JTJSc05KZV1lg8cfBNeP1mLF2v4hBJbUekJuoxlPQKhvmwmWRkZb8rWfA
wI9fRWlBN8CkDOe3GKH/FPEH//p5rqXp+NuXo9/oztxb5U6DvS54JsaA51ZX
5mIGSrx7stPK0MHOTX/i+kGNOkpQlQpbBbjL3JfgyadDYhwQa2ABPMDOd9fr
F3rnCGC7Di+a/7Sa7eL+XuxMZ+R1RpjkXIHI+ys6nLHd/Mhut5XCRcBuvT4J
L3DafsP+dDProzrU2OwDM+D2fEiNNVwbPDqEaC0Rpc3k9x0p4An7ooJDxrBr
ejWrxCgaTRzdfvwLWkXNoUQqjZ8KQK3C/ZvE92l+htMwJZgA325m1xBErCnE
l6ag3kjWqTVeXXfJwOwkwmsMME++tg18Z86HtY/NYeAzUF4g8ySre8sLOTmj
lCaYSoIkCjNEveItVE5A1inYZZbAv+tVEsW27CD609JyA5PrDDtI7Vvyva9Q
SsBYzk+mAs5ixcKoIJzujwBJ/KVSzdJ+f/JIkfUv77NwCf5dugTg3xYyjeo9
ulLVEKo0DzIxAO97ogiiDNrCJayfRe72paA0IpG9i8C4MBCsehpVMDglKCbo
B2yPa0t8qd3AK/QN7B+FwMvB6qsfS1ebQReO/gA+ioh0HNsDyyCAo9kivmlk
xMjrIoGI/Q2FqqXkxtTRDNqL5U+BlNDo5dhM+7BaLNJz1zfiDhHn8tQsEa14
Ce1pRiyA5ppKUgSTTYHJD/2ZFj5mgAHCpQ7rQic+HU0YuN9HuhpGSH2wgRKe
l0iXqvAW/bdM1PhyRX6qtSlKBWdAYwdLwk8nIRyZorqB1F1ixar0NB2+GcjE
O0tgcKcBogbS7c1+wm+nO92p/4fVcjOEy79gYLuFdLPK2Y7dtnypF+TBLl3N
unxyLNj8zfgX0axLPeXK8ddMvQLTHfBLPkVa1cOwA0nRyccIG0Qn89vzOpJV
sQPsJXLcFVZWFc+jbDiBFUrBAzwsg5e4hVv20RIOfN3IqdL/tQ9gBXp47XRf
KeLGXV3MUH1MuhiyM+G+OrCtpprSGnQL9PWU1pot65Iyc8QvnuEJAPKvtWlX
/+PKcakdniy5XZBSHN5QvGX3b7tyVWor66fiCaAoSZ16bQLhgU70sFHppvnD
/Qgy4PPpUAYl/w4ckxR5ywQ/h42M0zBvVXQPBJU6hJ8EXrvwrahwKWkTSvyy
FfKWgX2Qc6MGEeOr3heOB8NrJkffgB+RZpbYD+zIm7W8beXC9DRRNf63EQwi
iuMAp6PpfMZray4UOmWBKEAGcrXtuWD0o4YMJ3A1hldXnnqEYx80SJEXK56C
36JBqT+ZjCGnEvZlmqTfwT9HNh/yIo61CATji0Ln9dTQCvbL2ZpllnPV5FLR
GGAPLexyK0hjj9O116nJsga6EVMqsTrpISAno7r9lsfxrHNU6AdYcQR1CcSZ
d//I/Mpk1FQcPIgQ/c8MmNquoJeXv+gRLqUWbrGoxQB3Wy58rJSHsfcHUZAG
usNll+wgcCAxDJ8DRBfkaMBwFyrtF36nMjnrryZBUafun54ap/WHera/j0fN
s/Sfj0cw2SHWMWdc3mv1T5syIc8kzU3wqrZ2b4y42EUeCU0uDz8ankNMzprY
76Dm8WuNTJrEiDKvOwHzFwhIbX5vPoy5VzEAbzq5hyOX9elO/1+Y7Fd97oIA
SlXNPI2jr0wswkeOK1ULdYxo358gmofZAtEyFno5e4AE9kEUGhhZKpJdTbdl
XdKt9yVZ3CJ7+xSz57rNMET8+QagFhF5u4SJO9duczfyTLeoxsG2zAYsmAYN
4LtQ6l8DQPbOwOzuXW64vwNi/Ysris8G6N7FYbRJF9BxGJqvlH9J90txbPA/
miU9InGydrAFs+ujL3q14EHjxiwqS5qkdalMhEWKB94BTBt4sVln/emqceLK
mjugrgkiZZRz1SA9z2C46J+4Odw6b3TQ4hU3P/iBCZ87WIDCqhm2fa1thNLB
g2dLoME4zt5z8Xrk7XKktX8Q7EBQvrITVpmomvFIy4q1MU6YI3jeHjgM6dx2
PPidkXXRXQ9+Df1bcef31CEZSPn1hPwcZsOgR2f2SuudM2wsN1OuAgCm1qNm
VVIexjLLdF2vgVA9WoQ8upg5AM4tVxJT2ZYy85dmjS6aVfCYu04JMPh4BoWt
3mTqq+FtSaVXvlysM7cZ6EcvV3O272sXD/5i154d/+5DTyCBSWbdE4GlSorY
PtJLKQhFXMrT1JqZioVu37MuLPKtFRnmzXW6VQmZuXw8FJWMrS2BXm4z8ipy
LP7a3wjUR92ve0gdjAZiWoBE3GNhRkHOr1WcQ8NyzTeBo8WF4EPGohXJvv96
3FoBeFGS1oBzgInrJVy8VmPLzWUoZrBhuax6FElILNQifTMSAjISr3OWwI9K
DBYZYZBfP+cQE10/nVGFm3ZJv1M0bNf2tfswdOU2AL1KPKov9HSa+/uUkXaP
GEzTHLVYGBcob7Ls3SBxMi1Hwg0LQ9TWNoYe6P+yhM97ss2kJnsmyuIG2Cet
UTE5iiD9vLYkoGH2e8EKAhPIfTczWDpWAC1pW5hMe10GhGDLJMz5/onOEefb
TtIG/BKhwjrK0i1fmipgLElJwDDf1bkRxcvOVpsC2pYndFmB1k0GftuzHebK
e8etLrVluiuDbrDMyTzB6b+8fTRi+Lc8w6qVg3X7Dd/J4OS5z6vHkQLtWmAx
c3NF4iwcSmJvWWgxQPyjHoNEwtgv84yH5TCfqU9t3SaIzd7MP6NHPQLatcq2
1CcGN38v6wOeuA/HXDgZ0QTMaJuQ1RqToQp+AJH/e0qD/WCfROq4FHoeh84u
IDaEvSJxa0v/kMjMIC1Z35sApgmfra3LYZW9Oh76CGmFk5H9GcUDV/jlPkXj
Xtm0qOBs1tH/BTVTV4uyrgN59lnLxUAdDk7o5bPvx/vZmF9CyPEdyXoWKn/2
31VCEfIyHg4sI9ZhQOlxVx+uBcB3L1cTzXUVinDWBZPnNseJwKr2J0dnRo7r
HikZTmJ4jCtCUC7tTGvLHvH5FzjZHUYLtaaQyWYy/TreweEH6pK/yHMjPDoh
2GGM2/qY1gqQPdbWCo/mrgaaH14CwvSEyPwZmNP9I/K6w+hcglHd/sVXBB7h
4f6GW9nvWzrfCyDJ6518S7L78zYBMbGq4nDJRRRupYXvhlLgfzxj5E2Yyqx3
ReayMMaVaoyHvyVzfLYAPCEtDCF4Gm4+Kb0Jkpb7XWAI46rp4+/CfaYdWJCg
cRBjnds7tODbzrToHiYFiH6l/MPj3d63DPKdpySFGM8G5bnG2EViJ1vCzgHQ
k5ggX+ogJ5wpVDt93IgnG5BylN1aGbCuUF5hqZILNvnMVSTT6xqRmtrHhLNa
Ne4AYQ+dfhGoxZd/ctLEMjRKoCV7gmEixMVW9m8yNfbh79vFgio4r7IY90vO
0lM/ipRSTJBC146UvdtD8cMLOhr+63d4sXXsJrcGOGEaezm/+/SrLqeBkfRR
qKuOM/ttCtbBcdpwFgmJ67HjzpM/lgAnVCPe24fQtnGHy5wmCeT0wW3+SVDM
SQgQLEsqRo4wTUKLNV7pKswoaJgRMhqe7M7Pypm9vycHgi+L0cRYm1xcBO7E
ajSg2Yw+jf9JitkOMzxKSlk1znmjIwSreh5RfpJC5MhUmp/j3Z8aK2kLr14P
obChxC7dWTl6qakaOSzO0N9PUjXeEbIS4xl3rvqkEDxzdbK31cV9iWe1cu7v
wNMbYKCjwARi+5/au9fR65SYNFY6KzosWp/a4nSvqQHJ9dxmowknb8BCdbI/
pJsJ15V5VqPqVETB+ICQvEtsd1ChLKIohujSkSpsXtOTdJNJ56cyWTGQVy7R
Q6Y1xQzF01GidzBA1hHmx+Uf1dg7V36LiYJew9MqBdHW8EcAhjjAlQRzznq+
I67rDRgVAD6SG4jTJKTRB192GFw3G1z6paDAEgeB/54OV9pwrbMOO9B+t36K
2lUFQHZ641Y/k84dX3M36czmWeaLI0+7GS6zGyktF+u5+LeFQBqohXIPsFvz
5hLE6eFbfFRW84esb3oo8oSC/XCRbh0U05NqlrDCrbHmg95LHBF2rpyvCJl8
fscktOCcpj0z+kiMAZ4GNO2dYgCPPasoiLo/LDXWtgt0wBWPAUhKQoUlR8zy
TkSOewjDeXGZRr7/KRMVSk3aeM/fkhhUAHxBHEY1RPpcvYq+Fv33M5QRj/sd
AkkJWExffP5F9WSDsX5g9lVSdkLlrLF0kDDJCAONSmVVjDSkUo+GOa+URfBZ
IGWJOhs1uLJPzXQLopmnEQrsl0GWhcZSRDOQUsVwMrWyJKJFYM+oVrHwPXMt
m9y2x0yfS3E8WIx0ZI6g3ODYZNbDhaQo4yPfuvTzYTP3wop70i3o3cEh4Xhe
Dg1KEcIOzEvOumAcTxVr8t5j4ZyX7nbvuJwQ3wUpoyCckOPjY/ko/4MmOreM
6X8ZwA4flQYl7M3ZwjftUWogb2Ydhdf7+a7yn7+eqb74gbFuBDTHd4XBbs56
xGQ1zFk2pobDDHcNikjaqXdqa6tBbxLeZZHnrQmJ2uJyHq8wrc2ErkW8/MwP
4JDBMQHtQRBroUQrIeUlSLAa6j3mMygULtx4y1FFhuvevL8Yvof83wdXgDQC
jVp1d47x2XCF0mR0I5Ojh6YrS/mCWfsFG6tMAlCEkcs9mbLqOZHlRUAPXFvp
tMQ7TweRzjO7AW292UzOKfbe47+jwgRK8t+IjW+t91CKGqUSTNtqfG194WX3
bHwdTFDYrawSeinlJafu/ty2EngqGgXx6Z+nSnDJb43QUKFRoS4ioGbwXffB
J+HrsCjim87ExYOLGSXnqa+0WkxcFP1qjTeTdlvXK9mtu3XahIgSMp0mY+nz
itoj/zYLbQMWp4Hjrn/HE/Axl++77jPkWTvdiDEhq/2NrIKhgfOu55pZ+cJJ
xBJ34EwmO1UcEWn6k2EIvDiU+T5+Te1DF+OngduoElLgLtw5ZvfaK8Fry7KZ
mmYM6uycMzyMt8AbQ9aJk7AphIB+mIUex7AqpxHULdHyGo1OoLq5fUtHY+oM
ZbDIPO43N/+YTADQ/u+sAxPw4HqG8yfy9yYHjB7eU1jKojHql1hGcVWuvsbq
oOomiqD8S+EJn8611BlpJOjlPZ/IG3cJNNyT4LQlI0FnGN/MGGVR66w5k0WZ
nrLLrXvF/mKmlAsNORcJcK/BLV/AoVGhxXBbDkHLilz4atH4qpXfWwPjgERa
Z2DgB72Raw910GspdsBeQGFVTKjVXuC6AtogI2rheUhR6nW1EjTr6B5KgHM4
CZm9PGdUp1Yl1ed/CJymgSt79oVCaSRqNGFh//Y6sp7WhByPQ0XsXR7GOtL2
B4UFBTGd97NToI4ttoXp0xPnx4gXWkJFnCHWn7yeiPswmpOP/c8I1dB0rpLp
spY4LEZbjRy83TGkos/f2caYeIKA0Rw4rz9JlugjFdEqhLEU8VrJHdQayiLo
JWzoHPpaI3ojlq676Kl4fhYsvBw3JtkXmieFSQv+Ir3QnnWCDpMVxNBIctGW
l2uPnapxlYhSLK7DaOijUhUnLIk5kgG9jUY4FnKULc7vLUTRNpRrUjeMZidn
/XqIc34uvIV8iyHUCsKGt7Gva/5Ec/xyQSAsIHenBALaz9/qGUCTAgQjyX2f
nNPVOAdf6KSXj8DEC6QxkJhpi7SBuH0oEZ/wdwUFLT5ePDyyCbsbTYzd3t8N
ZV8QgXKcYwQxlmJHT7+0Airhax37RifgcnAGU/J83DGZlGBxd5OJU9VTn5kS
jL0jQd9AsFpmq39NY5Qd4HqcVLP0Fi99pQSJt7UgxiQ5p5RCVK2k/wHfBBos
Ygu+9RmhpohkSg/cy5kHlEHgvuIxs5X8I2oQ7+Nb0oCvxKMDKUwOF6tTmf8j
WbCUrEo1ZVsDP5s8DP/TAJyv+hocKEvEnQ4e2m7UbI7YKnkzHoXMHVnc3Eq3
OUSatCCsuFxKzX45WChbaD0E6Vc/ikkkGgYoyYYkpImvt+IJXiNqUz++np0j
Qj5yKza67yXNvlVWf63CrUqcOMJMVT0xRaIZCKrwiKbnzPV531hmis5AnAWL
g5CK+UPfkeSuzv/GN5/8LxU8juYIFzX7iHEZIxw1E9rfxCEtHBnCXazx58LI
vym6Pdf2uC+H4NIpouFd1zcSSwD+FIvWsEBmebF7D+tWv3JuNUG8uahst61f
g7dknBt+o/cKbwrdq4dkAtp/CIEfaZjUSL2rpBz7esDs9ty9JFRL+4yTqQNc
OCeNJaSZmUCCa2Ff45wLLnadd28TuL6wUV/b1P5wBxrFye1XikuPvete8fJ4
nRvZ0R9G2oX9R+RGMEM9ZozH4ejacvtJC03LNqXammpYdCx7srBVlPOlOQze
WMz5aFQLTZEi4FvLeAqhLNf+4ju9iaoF+OmGodQ+FuNoPuUC7aG+fsfFbGdQ
R2MwoooVJ1GBEgqGggwx4z6uxFS9P9VAk5Q0gs1TwtPyzSSguNZkPO04939D
4Ic3aFpDHXRdmfWXMsnFx33eTVOr2Iy4SkKgKuDEO4knxrOI8SiNeUkeWCNN
zolFSVjm1+Kjaq9qLQ5+SjY3mPdISflXw8xld1GLeW76lZxlMB3MGuvjdbtC
x3Z8hf071u8b+lcjbLHhYGznxKMdgqyOy0QhfDSBorj7D0ban8a/aaCVQDnd
QkXfWDhOdpG1d7RXZqBuo/NlQE5WMRAH3F3JoyXfUgU0SQX8pIfXkD8Fm+sf
7y88mHEFyJmUhs/Kxq5K/dDpeKRqmZeseO4BLHFadtqUUNCCazciwSd1TGoV
Ryr5UujlsdoSpwzMFH0/4EDe7XY8ohoVya/SttGjLt77flTvS4MHv+7TTN/C
imR5bEOueundwr+ieitsmRSw+99xDoO15I66OMj0Lw05b2TUSxqhItJDht2f
YWNSsmc5sI7mrAYViKtXECHbFIBIFnjl7sQnGXvhudmwekBOAz7jILlTLRNG
wq7iF1m/MgPJWmK9Ex2hiHOgSDXPR07FKpjwqFyJ8WSPz92jPlFOVBsHfeB2
HjgXshMkIsezXyQ0C5pIDvq8uF8ptSZjMalnboL7RecRhP6mSvhdtFN5UUpD
U2pa4AKRX/Xk68iXQbZmwPE6YndS3EIGtR+7sou+LW13YoVXgdwq4IzQ3TyF
/vTq6BPvU4jl3IZPeaY0IYwWvWOMD1ZwOYCx/kIaKOMzMGl+3+j8bXSBMCOk
Kw2mfslk83KviwrnG8gixJzKeQAdMNNNVttTCQ++mqJxkKxtoRvRTyUY/tvD
0EqtFqISd7Zu75OKTKMOY3A12VrzG6sKYTcbysyGyaDUZVQLEc0iTlsOOFFE
XdDRUs2Sc1gMHG1BRW3BBhVlCuRrG5jp/lAgxVkwdtRkG8LuBJgffIvLrYBv
cZ8pIyIwVS6R+yzdSCsrjfFsTR4lY9N83xzAcb+JhN41Tu8RvRnAVicmFA66
/EAbObTS02io16oBydtPgyu2qGFqFL+i6bUIq9pQHuvg6BakhfXIftLOD2tC
tfoTpppqft6sPrG7rVTYD4SO1poPKfEMhZjFWQ0htKMs92dutD/vrlyNssGu
q4AhfesnjZgXOdDnun7usNPX6v6IMSOC4c6TL1WHubrR5qZRNZaPdeF1XWs9
CvhWAN7c/7ILugDC0/WzGDTK8xkkVrR/iMn7hPPlOmzTmHI5t5zirpQAeP4o
yN5ziscESIqI6dyBkcK9p8cBwVSVj/mOiC4RsXhIKhTY0OT8EhTiDdNOeAcx
nq73oVlrstzhe6OWBEH7btmS4UQYtNadheXjpUGUQD76m0dT/MN6Ewr5xNui
ruMIcW1eE68/kqI9w6OIKhjHzTwNNQ27h+noCQcWPIH699d4pAzY411mTUZA
NgEUPHiTi4WKLg5xEomityUoNgarBi35NigSc5ITdMtRi/sANUAmqIG3thP2
bviZYXUY6zL3VFcE/2qs8lQ7z8J92bVfZWR4ByuTxRmrsjdNU75xqyLN4ugP
+AMNrvPxt+RytA4FaU4/mag5cVXhVe0ojfXLe2Rb7nuJML73vdghLKxKsqzr
K0QmItF9CylF3Y0PnXGp0+jTSmjI06+5Dce7Dd1Ua0uk1UMOndoMZEZiIpjM
KhlFGNEMemMKIjiceW4x7O6PvyxgqmHzzTJ2x1xuUJ2uIKtqQvaMUYELIpt9
ImZzwxUaBClVla6rUkOQsIFcDUwvOTaHGh3rewaky6DoG/9B+FQjxQxMWRW+
Wwg6ams3a/KwsiseBwoD6DNPm5dAz8GNOXGDS2YtLLI/eqpb7r7A/eKUHonp
XC05wa22Xp71InByPFgEXNYeQoeqEwrM1Kqkog5w3W/gWhM3epXwIg+g/7h7
aVIO5cRmjg6zJfQ+aA98ADpISSNajf583SjI3IslHbL0p0OsZVcmNMSM9F/y
Xp88nNt71xvvITOMU+GvLgd7ub8UT03VJ/nl2d7azPF9bhKFfZU+y0duiise
yyktALvam/9DULxGhIMZvc0jvRgSL8+96io5EKQEOQb060G2I2X98yrqA5m5
NuyvB38XFVzYb9HwKdQN8W8bOxDfXKFqXKyvuuOo+u7/q2fjs1s/kG0goxn1
I9oGz/lmDK7AEeze4EEZXiHd8CLSxES6D7hGIQtcyvd4l3MKD15hNCsPO9+2
BZDVolH9uGEB37L3Nt7NU1L3Hgur4xcGh/W2ErBU566RauHBPvDy/fm49mTe
mDU1qlESPWAGxnAH+4I3rqvVk//zM/QRTwzhfYsNguUVxK8XxSEZUGrR00OS
Asw/6GVSo0cdX9eWBbxIGMSrD9fNbRxqszA5dw4gHOJsL7+OoeNolrl5ttae
JR7ALxJdy38uofNSiIM6vpF+P/AYADD15I21rm9GGvb7QvYhOBmLgxxGLXiP
R+N8zTpPMl7Znb+/KBHJRocaRFOQcixgOgP9gF++KMa9RxWhAUza1rrwkN2R
UbYxf83CEfCyM4uM0dvL2r1XJDjupDlYn+i3xDFZM/nx1EN4SfVuPFd+iPzR
6D65O4I0+CvsGz8HnOq8oaNVtYP2IGmQD1HaAUpQJak8YhQxG7APrOf2qksb
xmelEBKGphwIQAj6pmZ88gZaFNg59+dWwXCdPap9b7qu/JEnayecWLEWvDrW
e+2w8PQwZu/eGwLkXP0/9NrIetsjLLtGZL3LMzcs9fTwL7ffeZ6RcoEdYCxq
eJVnwDesRR+tlqPgzfPNZGjnlMopc2usZ6te17hk65UQ969NVbJ5IpdPMnqc
dV16Y/ul4EhP3YwPbObHDQuzDls0Rz6A+kg4zdVjaAC6BXc19FO5/bXeUX1w
3jJX/7uRg1CQdmKfZ+9tLWwVVZUg99gu1LLtd5N0hfiTOKVg/DNM8UyvkYz4
SjhL05/B6Cqxu40saJmp/5AWdDfSlK57StTEQN1TdYJ9oe4bhCLpp//GIzsS
aWDR6MgF/gobiIm+/RdhTrjHktINIshfjG7LQnX6tTGaGbe0M9Ln8Hqk9yQM
av8Fp1uAr9PBDjnlvWuQy24vKe52QW0G8pCz/uPoztP5DD6/Nj192qRtd9O+
ScTOLc0JcCUStelrQSSZ6p4iECxE1ZkGXuLdJieAfRGLjOeeRNxRuMGHKW4u
yHgvlH1OpRPxkSWC5xu/1YbWpwdqcfUE/o/SL9djFNgeaMX6dU4RvlsIBCLV
5eD7y7pUBbfr9mMcAT4vi2O//zxVUJmXP1u4DLrtQASAaEHV1KLcXUJLgJrA
wjt+lZ8jYroqFMbTFrUoSZmQjOMyRtK1M04vMqcwksbhapTqt1LOCUSzFSIw
vNq19gpX8jAC1EB5xtG3KX3j0UVah2b+50afzSJ0/n4NXFNtv0cyufZWEeYo
nmfLMasZ1vqJSfbxPKCgF98R9GtpvBoCN7/yVqCR8OPB2IvNT9Hy4VaIWdmc
d6XYCrB5dd91v0/GFeROBJwNrEchlmM5dPK0/WafmwkMFu7idZiaby6W6djT
mEDYBq8iIQnq4SuDvjx0Y8ZQiwN/G7wpzh7A9rvX5DoVKUXzi2Yj5xqLuunG
cVlLOTI8PcW9kZ3cyvvZ5FcQ4hIU1q0MRa3+bSgNN8ZNI/aZD3ZonKuBn/9K
HeqS0Fgaw13MlkMskWlk+KAJgjAO0O/qWPEB623Aqt9/jhlQSKDZCVdH0PHF
roraA3Lg/aESivt90uUAiLAnTuqO0kzrZo0tLK9AKyPplXLWYhh4vJXKONDf
235w2rliKMd7AuplQGutZrn6sFDX1kWa5TIUc/40wUSk3thL3JvlfNjfTJRt
keMinIf1bIDX66kHyE/jdPXxPKjWywLp7+lJ1IiZrT562PZ9xxHGzUDBckLK
AzR4h12+NkPhRVnAx38+OHaYR6CtGkr3e2QbiM6NZTJ3TlfwxzErr8YiFhHs
WxYfUmPM0JTurfqDIcbZyWlfORFPjXUx7CluFCFXL/n4XaBqT1teBbQqjdp9
cr9KezYTE8C9gw0aiVWsd6z85zlvfLpZ3jR2jL5K3DhR9MsfsC41nPd2pDfy
S2HujKUg/A4cs6ryg5OEfjhrYOsCrlHHknp+AMYlzbPjgM2mqoWAx6Qw3zy0
S2jJm3/F3PX54bDhsLzDYHNM2oD7moxBhYY8cUhrCtw/pMMwRObStX6GpeMT
SmieEmbKZ/cgFFapNZuddGE7scwozmUU1enbfYBVxefLjcpcUE7Cdhj8ji5z
Q4x3QrkhIVstYSKeb2HKv03YVw2DVvCqFFigMeOv0XZicU3zd7XMt/tAUYHr
rFlbLSSmQwJHOjFcFPQrHouxe+0j8YJ8H7VbkFcDV09zaAAV/2l566Kb0Hls
to84WLItMCLut4ud89LEPIvixutF7Q7XzhYHOPC3xVirwZtMTirZaceuLpHM
Y/zo40nQbb8888UGxFwy7kmwyigvjEDJFNhb/bWFPj4k2CXgaHleZepCmzyJ
y9TXu+uCJ5k+RSBqO+1zCXWHcGoxcj1DJuShZMcD4yF4J2kktd1XciC0Gpke
S88BarXC+qZ9yZTrDF4Vta5OcEtz1j0PTjrBIjX+oGVSQ3IVa2DMMTwoUBWx
MWnAPcrCHpmuy+AOXQS7W895XhsHjnjSFK/+pqhuxuO5G21ewO9Wd2MucoUu
yRfRAaGbH1UBvc4g/+3GFi++KYJpqpG5hh5KMEYPSKlxWvBXTBmhx6QBBqE+
UjUgcu2bKZHEIc4gGTQmec0EB5cvjveke5Cp3NnxHYtEGcjI60fdEbFJadY/
7TKrvkuHwIAgrrKPY5a7z0Zrxm9KtdSl3v4P2j0st+Z/A6LoBB5gVIZKS7z9
uWUuFfxWC+Zr7BWy5tEsvsJLXgxarurlm6xlbq+dGxBoILYCB5BXd4yEcMHf
hHTJoDKPIHF12fa2WAj++ezdDmnB+ZyzqZc7Cm9pog6pqR9DWLskXBbFiwQS
zHp1ugFOZZUcaMaMpzoDT15KyuP71zAgrTVNMDFOSlnXF66PV3ynACx6L6sy
2tq07Eihtpjv6zUZ77LgSF87xZj7UfaTTIc4M3dRgjc8rAozzzWIOnADLxVf
PhhZZq/t7BoO7bJt0GNqkg/EsSFg9rcF5a3m5k+f6Q242z9S6QWjB/tprjkJ
wtlMztRD+5nxf4yARGftWagF7EuXfXTcWih4A3sNxzsDW6Hh4+gTD04Ymv6O
sddxnbU9IBQP+holbQW4jHbUrdN20vzFLmnOVkw6ocucAak7HwnIW/NxzUL4
d3HtDdpYbxF4cA2zlQCVpStaMz0vrbjvtt5zMX25uxSLPt5RL/JDAeGQWkXK
BxeW2deBLdLycvaMxCE6JMG06ctS6DokddnkjOH2AQRlMpvmR9IzXmgyi4m3
vDqxW3jAIaRCL18pX61lD9pEk3UwoymZTUg0HwVyhLJjWHZdkLXj8JvGPJrQ
ma9r/9pltsjW+drVJUL4lTCs9mkvFl9gXvVIIgHU6wNw95pdDV4TcM2QnHhz
cRGQdXbGOFtfUBbJ7ij7fY1FI6yTs06en6OM4MHoQR6SY6h8DV4Sz3agmhiK
L6cxPAnxu8V6NmZDhXRNBWUnCP3soVMBG/wHSy2hlQcwpOTJ1lp0/iXfiBIK
fr7T/zZOYlLkRgb6mkMplxpl3mJ69KLJTTWUcddL/USu4LkKoOCxHwr384a2
7j6eW+kapSlypqpxhPSWSEhAFt/r3BVGXIWhOgA1yz7L7V8NFuqqE1AoP9+u
a5RVfBmX038RNdf4T17R7ACFj102Ur8hluc6U/hmY81cR3ZMNqPEeZpROXdw
UodYd7dVPB00gZ4JmNZVJiuXCy46l8WBn9LmbgL0mfdflb6GJWq4/ngrdKtQ
P23F/l8+wIDrvVqhFgmgTFvoeZfgxjfBa9zh8846XYnB2QTPsX7pJqSOhtMO
e81+N+aGycNwm16AubruKdFjV1q9LzeOlJ7XSwsqW83ABlHb29CdH3a+hNt6
AW0YCLZg49VvZfVa/O1LTmVxQrEOJFfD0sCyNfyELfUCb2FWoeMYOZ4sgv3L
2PAcVEXVja6+4RJqrag3oZRzZmq1SD61c6fRicgOkbj7JAWE5en1Rg0TMPcw
wsHB/PeF5XPZwmb8Rp/lIR2WQNGDcdsBcTJCJT2sKHjg12XqNhrU94EpVWL2
di9LqSlJmwrilv/aUbxCQWlXEVUGBPB86Ua9zDsCmMU07EeShj8d0AH9Xlzr
eQ5mdPjvbZCT8N4sUhHdpE/0UeugFOZw7DxW3t+hdNJ69fjWIK0OxrvvQxcj
0D4sxKJwLffq02SQseCqFceIH3Mp+89xfC5uim+0jy0mWzegwRIzYUe9Xzsb
EzAbzFUHZEm18LTt0uKuGdy76uYLwuliSC9i9ol2LvF+AHZTSNJx77nBzBpi
sqr+qDldTn2oQGQfxkbivQwUr6CPYiWZnl/w+7Sk7fsh/MUBlM7U5561Srl3
Om5dVOq/2PpefrAyiQ4KTkeuLSc0L5xFUSZcdlhiZMt/wXomozRMj5TmPAm5
f+ffcMmuW2Zjvk7S8L1jm1Y1XDH5zMKNbzR3s+3Tfk5Ab3plLePwkFqY1Vzp
7uvjvLVRS7+iQGP1a1hUc/eXCO5bZedpLTDchepNJyNqNT9eTP3fEG5rop15
Ddvi3txSNR4S3dJ9/XgNAQlfkr70D640drLKsd1jcsh+/nexHgFzpl6vdOg/
w9tQkwAZLLk9MpCzqwL3g55zj9NziKirpzLoLNaK/DiZ4dZwxK3RONtb6+Xt
TMWlpe9keyWn90OlpPoMa94RHwLK0C2+XtJYKgNcmvhooPkSJe4TJUxD7zVd
Q0T1SwBDgnaZBckhcZGM/2wHLkAh9epy34VVfiiiQjljpPHV0s4qsPaedXqo
yhaomSvWQtvcsRsbtCVI3200evSmrCzzB8emCmPJW0VohvMcs33w2KeMXAj5
lDIpMuhamvnHN4Mgk1skX740OxohUJeFwvgKWgdbpu4LROAp+fj7Mp0Si5US
WJ5DTjmdw0aXH84pkV7AAts+pBYRBqiiJNdQx/051rCer82oWseaVgujA2zL
r707XDQy61h++4Lo98Qt2tZRudH8EIiZBLbdaYo26V6avdAZTLJ02qGs5G7p
IhgFSQaliPL42bCIF0bLbu0xXJnXgTxsivszdSzuTXQUl4HTS3Hjexrq0CIJ
53+17gW+iLVxe5ag1KHipossj5X01QQjPZm9VjrQRNSZQjSOte8/xusaihC6
bbfBJMO/6QynQlr6Cll6RmCqNiMrLTFBuwCRZ3odqrMkxe9k1EJje1y5PxER
Gdz7pm7ExEByFQbCOFI7P52pDaEI9oxAvNRyjjxPvmToJaDUVyWxf4tGzx9L
M25pNFpGm9ux71cnCE1qyy94eHXzo7P9HEBirx/0HC1US8L4QW6hj/GeYfVQ
MLONC7CZXXDYnBPhhi0ycqUaEWBCCG2MBp0PVkqd9M3QdHj2eFfW092skteZ
bcx5N+TqpTXEUaZJ6P0HOcEFMKxUzPKoIiengKTonXMDQQYt6+vltH+XjjyE
In4Q4jyvYoqcpDJ8KSQ/c8320kGeLFMoO3kLUNN3pgO84WHirVpV7yEHt2xr
IXXSJF1dKhIQrR++mwfebgLsivNEW6vsgMg/StCST8JoEj74SjVV4Hvz1/TX
LcH/lA+36WH4hVZ9Bi8MOaprXHn8cB54q1Idb+bBcY9IHCPZlrPEfwOUnm0B
AdI4x3sN61zc0y+ChTbMzAsKH2XKcn/WMX8DwCptNM/D78V4Dk5C01lGObF7
LvZokBda82hDTPKp4o67uOckIQMm4HZnEObZlSC8xKpcsAV7M7AQmPO4z0kI
NeXafC9ov0I+G7m1STib1c6JLgErZ7tBZmxQvBgqoibsSY4UdTAns8OgQxwV
A7+qb1OktDtKtGLXU1Wb8Zh8DBbja73NOTQQv4pVhOV1tvoSlBs/5+O49Qa7
/ejU2n5YE2VjZu9Qhc7A8fjXLTGeRZICNtneWDrXVK3uONw2NaO1+oQnHcdM
O07xwNXnmUK7LUIVEzFmDbZhODFSZhrcJOojm81lTQtfJdcsh7sAcweV+8Wl
VF3evg8EaqiEXxpX6Xhh2gvvp9J30OhfEAwdofidEeTYOGbLsdcADjf8ubnV
yhKR2O+NP6UW3Be4su9GfFJfMO8nghQihobZyXQQAyHDrDVV0MCIX8aoUS6G
ZEW0ZaMYMSb5kZ+n7thuU9OW9CzbznQQfhgyxBtb9xd8hmhbOR61u0dHkd2c
kaigq94h2zbimTLFRuLoRgzVC2PnBPuijysODOQpYJtdHsd5PODx1+oz8Bnw
h/gIOAIlqiltN2bYzvncfR3knPUmWVFZ5R9Wk4oYXGLzdKwP8naFjwb0JN6v
3Zhp82NSq0MkM1iyLFazIyx7x0PEisp0NRjccV+5fs6u7GaFKxzhMT02NPS8
MGCYG9Bry6N3s60qy0GSBqf3f3iG8WVbHlf3K9+t3SbYkGJI3nmQU0KIQuxB
iMIaiyA7W0CdtnZJjb2KQIkoa3ZhgCMdRGMdUxQ+CU0tQobHss/5T/lxVfV/
FDzqxKmSZ9JbzcO7Pnw3rSexaOntsI9YivJXn5Lzo9L61igzXaO9T3e6rrum
K1jJXScx17fOupOl7YjQEqFjJAHSG/RoonHQA27TRnyTSBGludtXEjBuayiL
y03iv4wVUt+QQ7H9VZ2NupscUL9EHVz4wgZXR/E+Xu7g+tLoUud4wSsIbz4w
RPUVkHkJBF/V/bzCdJNtIqvdEhCcXxRUJ7QIca5Rl8JpawaNJCnXI2wdS7SC
hWwNeL0kc8nwZ1dnmfxopcC5A84+feJBM0r2uTZOYv53wTOvLvx9ZFBuhRyw
Ikg6Oi7dEF5ZV9orU23nVc+DdiMq3OvEL5Xmk8y5aH1l95fji+vG5nyPuK4o
tX6LsQE6PK6J9z6S74hPS561ueGZNbvwafZncR4gqs3iSMn585h4oUIP6rLc
M701U3BOYpITWsi5iwFlsrhDf+zcFfUem4EPzMgxAk2VrpoJBFT5Pp8Yix7m
zPvpNv8v7LRCEJwgruPA9s3M2okMcCSt6Xuolt3BTHQ6V1hrXK362xznfujV
ue2GxkZwqNabN1xghDyjCmyZZE/yA1SiPiES3q6Uthr6pGKK1KTHrtq7togL
LpylUCof+t9H8PoAMrt7DZ/p6NkGF8TzVB9Iq9uLc4ddyrquBuYybyZ/bpu9
1z+5QIwZSHIAWhV+719YApvtBlEZ2Kd8Ox9AJwsnAF3KZCR/eeaZ/nAgaMy4
ewZahRFb8r3hkfkoy+kt6A2LyEtviH3cOBSRPH/X6AwlOGFM1G+KPY9uMZRr
M2Ql0y+c6u0rznw524uZA4C4ZgDefjA6bMzNAfzk6UtHa0nBFG/KfJbo8Vpb
rLEMpmdRMQFYXxphXACuxddhUdvzYDXh4VCfx9JdMfRH2pqaw+T7wrAE6hF+
WnE1bhHt8QlUsHWn099KAO8nHc9UnTP5Pht8ZuTjGdxhoZnpbZqHk2CZa8jk
9ciDWMMlbE6hAUCox5UIL8QL9WNtlwo785AlPYno86zVv0FbzKzQVBfEejpc
5EET7vUTaxKHzyuNcF2VAh0Ao3cDKpZpHHyfljH9JDqrSIFAI4hrltcSzLIv
7yLVIwC641DmkB1VFeJsngWi8tN34T9sN0+AQI5f/cuChi9sH0G6tcuimzwv
kKyM8qYQEFVxxDlHr+POQWk3OmK+nq5KR0qDAGRAh7bJLcBkzw/b5PBcW7dY
LLPAgawk2xXUiqxgk8bbKs047L9dXbYffXVwVIhpxADm2w+ObadRSJyu7rOT
iZpT/R8nPJiD1KSK/3rgtAM7Mh9pw9wizMihFFGXAJp4GSDtZUUeKjjkgLbL
k9UGJCVllsJGhOb8f7CEyKk+cdSwFhCBSNdQ5WxwaF51rWwS/X4cM5AksqwF
/8RKu6ZiTw2jmKy6kXyVeZCGcjCNTBJkzBFqGDPUMEWCKPcaJBX3WMj55lPI
WpP8/EzUnfniHjqrGFl+MDy8MOWEMqm73QUxJvODrZ2GYr4S02ouW3rU/LkL
0tPajfH90qUXkSDOjlNsqMGqKkh9an+ikG20ghlAp/31h/g85Ot5HAGet7g8
NdyNQwkt7se+FDTvrGZIl72yrT1YAQYj8SI0b59PAHFVYaKtW4rRhtRsHmIZ
SYhrQOt05a9cf9rrMJl6QAM/zh/IW43tQ43kF2QvVhtPaF1clep9Rji4MYBB
PzTRN1iWzVIqaxL5QzJzei4OxzslLQ78OQgOlW2gHYDbBYEhUoyzR/9f8o7N
48a3qtUfRB6mmcQivOht1DJkbPN191OxO8EXreHeDGNAs4GsbT00YGFS2DnI
nbySX67bhnU8geZjFg0CBc+zfCHGfV746xSn3FXjYXmQKYKOFRiPe/NwDSG9
pDaPUHYEOmebUZiKaGepvJyPq9w+yhVaWW/84vX/xBJKrmJMreQFHDoHD/S7
Uizfs2wDhOEqgYVyuAOfrUV9YJBb/Ly5guTDnj7RO+hstQFnwwzDqAH1gK+j
4wIIuGyyH1dyjUKt1xhHU6+gtgZyR8STQclAAx6qSJoJVfw5oxSeQnjOfgYO
RLruF1yMalvP9NYTg5cPmDyQEf1tBS+hQou5+FgriyKO+Pp1mdw1R2OmkqwR
bY4qwWLBlRKjXURlN0oGzSlfT7NXtBAEfj8bs8m8A09zfpk7OhzOcqwHzw4w
juBS34QHq38VDFgdjoOLg19iG1POflh1Qzhcmc2oLysqJuBdoGtsgw+LG84Z
azrgh0ObEF7s2IVF87IaCV2dyEPuVzEzdpKxDu4PxRbw/4YypsBGRWURtwdX
3zTvR/mVddk1f4S+XxJH3LCE0keazlDD+huUL/J2G8ldd25uht2zHNuTk08W
VKP3SnA4WT43sgNgZWByHpm54heQsonbM/xTwJjkSW8pgGxGllfHCaWKtvH8
xFSZjEUA4t9yTikI48KBwyW+AJy0+l/R0ObJE9GeA9BuTOUAfeEEMutc4AbG
+aZwR63LrBILcG/VrDrD4v8XAl3jn/r1yk26/uFzk4b8CQIQajGx277kRS2z
+RrY5rlw1koZD/GZSGi05sAq/PrOCXExutwtExje5x5BjX0g4QvAresBqfuX
4Oo7Vx/K1OQu0Nf+W2jtnvczgdOeCWv/UzjSDPG7S7fwS7T3VK8ShUC4a2IJ
ax1AqnBLEpdBt7eklrM1uMBXx/2/BWFhtHyDF4WOp8cXkTsXsphGP3ssAYnx
Jm8hljeuib2oeD3G2g5BR8HpYzKxcn1klTdlDsWRDcNuLctCFyLHyyPgDDHB
BFBnakEZOlXvr9bM7SYpcfSOnMEX7bI2bnwODNEI+5xoLZC2VigL3pbo3QdJ
JKjc/FDqTm9neMgi39QDZFco33hdxYpS93ouO5TiDgVgwgRxLsadJ5vJ7daa
A4z38d7svAcnmE+TwXOLo8Oa8YTTmr3udeCHsYn0ymddiP1MnqQW7852AOde
oq65l3/wO1W0he+ZuoHt+4QkuK+kecuMZAJZEMFvBfH780n13XTxs30fNoXU
EHYdL4qczDuU4r9AEMxf6/vGn0Y6xAcweNseHXwAUClyTgAegXZdkCy/Wv7Y
nlfW3NDoxUtc+j52f2qI+OcJyLGeFnEAP1uUAx7MF7C+/6pjQueKhnlIHUgF
a2mg6CBl5pe/4ikDZJkDl2u9L+O60DFOcEqE7swCqubAdOJ9uJ2plyQkxQXR
is7L5cIUElpYE0DEYD8v6NKIUDDsmK61TVnLuwY7p74xWi+FbOJ6ZxvL2679
tp3Uy8UGZp1Zy2vow4xUnTREyljfNU7/nTte31UHA9YYTpPgtPDQ5sk4jvwE
5/Gj6FHfgCuwC2EFU+CC2dbksAvnDjyAuR7M0xlXHKMgcx+rAbJ1+WyR2Arg
QoL4JbHWKmUqEs2/tRfK/6klSLzIHdxL/oj5o0Nw6vtT17kzTKRKK8LZqi0Q
PkOzpU3cehBVZSQWHZrn2YPtAk+8i0F89JpOXTu+gARZBBA2ox6lFe2PEoIb
j11gl3bBBbUcgWEao01+Zx6r9rQ5p01nRg6QDnhCK9k2S+gJ96ccVjQwnz/U
jQXPxZQLF3JDr2ksWYWINF9OMMk5VCq0RA8hOM9/xTqelA72bArcyAUX9vJX
5Dv5qWX51pWe8zAWvTzE+tbCX5uHt/bK8B1Yg0+ge1OKLOdqS5Spy4fdhjxp
FbCEpaqrwdQa9BGqLSMhPPvZgNtCMKJOopgk6jo7BV6wqJHwM7KGaz72GQjW
JAjV4YcVOFxyrYeQU5UJnNB+dkVGycgcfvArumoo/qVMi3R6dBpfNaa84A9/
XK4CbZYHUVF1JR9R9Vqnf+lDhDhNIg/SOvt1uGbIwuFBC4jn3rdYjtFq76YH
ExFf2PHs+YE0zETD1tjZgnicpxgICl/ap6MAQN5mUY3X/Uk2zStoOeLiJsdO
/jIqS0epUT2tfLtmkavZsPbM87BojYb5KsW3AB7jaj7uwVC6eKyATdn8yqG8
wP1bFoOO5sdT+qboIskJ2bYL8huNwrArq1XmFsPmJz0mzOd2WGxT5p/tgIC1
OFsksw8o8kG75NLxTIK6T0ceHBjFe2X32ZJKRHlQyr2WjvRfAe2+MOBvErNn
UE+dcDjn6XufmHCtNF5livWDUkfgomiYpJlvuvBVyPfY3Yg8CVGXfUgJJg6R
eAK740BfHyQpsyBB+W4FnSXiqPpBY31nJpkvRq/J6p3oqSrfNkkbm9CNH1Oo
0g4vwNTk5J9kUhiore/NDmVDFdVpe+AOBQVvnIlh9gsBDh7bBxj8UXBQjNh3
AWscnKUkSF7qpsN4LIt4mmH6yxR9q+rP4YP0XZMTyY1aDi4WZqIKLFAmq7YX
iZOhaJN+obsSIolaMHXIy4ltfLV+od3Zf5TpM3Qa5Ee7Zoz8Wf4mR3+xDmXV
h0Ah6QRr2fVYqVqZ1UJA0GELO//mSnl+Af1K55KhaP3eKDgIwyjC/X7dyxWU
S8mEtsbSpuP+ZJOKnIpr1QMf0wbszw4khqukMaHkw57w7Q/POYp8cenkmVqq
MRvH1pAtu1Ugz3u+s1Vs7VI5a8pUvG3H3acs0kqWcOT5FGhTtQUmojBbUE7p
8B6UdYwg8UhNJSgLl5GTqdieNkjVzg5pdoHDZJRCeQP433ifdf4uEmBJ4f3h
wfuxi1ECC+SPmgHlhuAdaa7ZzBH9Sy1jvqDEARYguixA05jQq6zo6b3pLaVJ
sntCqg8R0YNgIk2+PODy3bmJMJfIrHFKRzqo5svzxGp+B49I/z8bJKZFYuW3
s29dwH7MT05PgXroOUW7AGaob9WF6fiqKulEOtd3vEpFHzpPsbLHuejd8var
ByNzNzrPFKm5V5rdsaPAkm+4J/ppSKsOrZFFe5oSNAL5Xs3H3SNZCelcihor
TpTsyvfmX3rcF226c89X7KBHnK+bQne10VDWXxt7oMsqPEsDrGAsGhEMWj38
FQygXkxpokhZGHar2wG0VNKoWoWTM7iZxpsyxtHGZgHNUwvWYBmj2GlKUFTc
bWEzk85rM7F+Ffj4RyTe9pBsa0r3WhYhisdfXfGFNPktdjMduFoDA8awb5Tf
/z7R8gxlN4nOg3Oi0Ga6pkutVXrETu+LEUNuv+W+3urpJs314bUPddKxEuWw
6O7YASs8ivXm3aNW5UnPywWn5KCYnYOkrX09AlnAOIS73H5rtKKC/0ZdMK9k
JBS6KlqjWdkWzjMuWSb+54251Td1aNwF/xD2rJo7PLQZPOLhhh/sC8Bg+7bo
05s2lrJDncA2H3x0IdE8FuJ6o8qg8kBC5kyprgLInoNE/fmsGqofdNG3vz2B
Djc8unT/CF4fxQaYjVl6MCK0LLBaM6zd7riiO7F3QAyEU6hvzKS/4KR7Tjs6
t+eX+ArLFHLGf36dPQ3M0UKoOO9KWWBQHvfMgqd6p9EqD76aDKiSCLvA5Kc8
sdwaXqxyFtcyjfw24CN2UWK/pWcoVNCKWs14/vG8AsRHVCgs3jedWNC8qyLp
OtsY2Hau6sXd0Eiiik6oseeiGyjKsLkRc/GuNkfdficez4gbhyRKWab8xUjW
0IFlRRa23VWq3Eyn/8/MhQqUpIdQBlUlVCz2J3qety2KVC7c8ubGh8Q64cu0
PEr1vpTWeEi+/VaPjjRbor3pyFt+2CTlcFG1x0NWK+dN5PC0cuDZIiehRwm9
4cspPEhRD0oktdTgwjA85RJsZXvddfY/SuSBVpfDEsgiezJqohzH/le85RZi
qF38XyDWvcJsYBeb22cfwFFcuDncUNs5hw0PYOvt+gI4n8ZqmcVuO7K7Jj9X
ebmNpsxc3sogHLV310c37YVuminBYlocLgJrYzv+xuh6UB977zfjPaB9ws0M
37usMJQi1Q10h+2u78P1E/OkXSBPN8LBLYOuxyHG2pkm8626G7fAbrxs+kkH
JPNdClzgc5bjVCrmsybZMC6BDGjqOtizfPRqQ4N6T0hLj6JrvgC8pRo2Tc5c
wk3IP+2lVR7mH5NZ9tzhT93Uu1/dbJttowrjKopnCro+2gtkyRHio8dlT5wM
g/Q+CcCSDzBwAxLq7na6uK3HkcY0EmaDdHg1ysIINXzsE2+Yy6MlyUBKqSBg
LrQ5B9Vd3h163FmIrEnKsfmpt1agKg8+l5Brn3YRz1mSsp/3FRvHsu3WzS7M
MhEJR+qcPDgzeWNV50AaPoE9XEYpYWu9LU4/FxpEHNlBEXY1EnDGAb/XsvJ4
PlKxgZXm9OKvkROSvk/UQ6jfR4NOq0yKCtwx6u9ZxDOQuMZ5XLg5ZYH61VH6
i0pAQLBp5OnLE9N3hN8fkzBg7L8eEuZLMYFats8TGTEu/fT3a8TsDWVshAJV
8phIAO0vePnCaoE8odK81fifEauwWOEvoth+x9pkLFxX7AD7e9TOgoqBg6O/
kXp9ac/3eDUUqJHJeMlO8cpQo94fuAgeH7CaWJdsvzmZ//JqAe5L1Es5f9cK
jftrkWP4rd12ulsHhfWb2ZPk9OR2YmCo11eZB9791v824yIlekh/iLfmeiJb
k42awQDS3hjl9C44Y8z+x1OEXWtw20oNIqeSoFZ0QmJhzWJoln9vLwrd5NkE
SmnVhoLHECNHQirpxO6fRH56pAmHNs8zrYmvivBjwxd28gjlTWTS/ibdzb59
czqiT/l7YrnKKcZ4y0g92Qsz0xvKnXY+8GvIVOLgchD8PYWxu5mNZHkOWNzx
DOd9hMre7q4ZvUiHYf4x+LOi/srhEI3fWzraTWkrpzXB20RuzyxBVFlPTytl
1nBov9dsjNePcenzZ68bejOj7bUrujO/d1QHxS1ZANVQHjN4zMJig4U6KuAk
PWOIBvIgnAYPVXeUpDG6bT6wLlvim83bxqvkGPOIx+4LwZAkrBTM7cnEMyAo
+b8B1fHKS1Xid2cKEgXy3O9034M65Ac5KLJozsW17NIuj1LdPnQepUC2cMJ1
ZGZ54gfvAbuPDEtbsTWOwZFFHIKsA5MyU+deRbhQIwO9wVffovB5bjO8YDWB
NcabOdOiy2WQyPb9KTfZiO86ZUSBj9R7U6YL+Cyr/M4HGYlogeVzGdqJZXlk
vd4WevSPbCbs2dD0igBkWY1Aotqdj/ZPVEvX2jEjvKnGTx5j4mb5JX4Jxxpr
6xPEF43H/XUjTwfUzagtKM9M3e42TZQg8/hHSL0eH4oIl8ZMJ13bqLZ4OG+A
rD/f/tRzOzDU5t95Qqslrnxq4BMolQCQgstzwZhBJ95wLAMjqrkoWn3hh/YK
P25rR9zH4g+MtVHL+msvS354CEGqKdoyHGkabtoXAr6SxMkxHGLcfjFEfvOs
YVOGOdqjalhU3y0oeTH1rsDhpmOFEYP6NXd3OBZaOgv1S8AFjwa1KDKyBFIB
gvKmKoKRO6Fkzf9We5LYH6ZdYm8EmjphdAp1bMKgGMWFacHOdOe7rwgiOGoK
2CN6fFjf+cG/vJpzX2UYwFqfIgTHfbiAZgpbEzEZ5NUfLyHKXoWiwtn3OYsW
CoSHjgRnZIBryppTYna9ZhqLArmHIWlMDGEY7KTwstO6lyF3P2+RmpjqEXoH
G5xBqM+cLSE0apVlMOkNDHPN20ePN7RYOgcwIuKlWYxfQR7H9Z83vMEvehJV
UmUSu96U3m7E0Zl+BtAtaePXG3fyfnRxbeWe8w0i4y2fPpFHjVHlUrEbJc2z
LmJujfzzNl8siZJvLBhrxgCF/HCtP6UtEuJvIUknq6hYJUOHrGlUK+rOOg8P
7G7Tet2obYgRLgyY36N27JaARq3xzmHk1Rl6Zr/vCjK+CpfJouEuTWkdT5Xy
zu2/CVSO3loNz+ShD/0TsWnZzmgB8xKQFhJLoKdxZPBkPPZ09VTe89Ll4vvL
7zEU9rT5nqiNFo5fum0n/XtX1Gpda/mIFqNtTh2oWq3+hRSiQMotESv7WUf0
GGnLexnGv2A217M7tjnO/2NIAgRnm/+0S7gIvLGsvyrAtP+fwOAhLO06Q487
2/gg20miJMoLorQzwvVdKUSHVZt6iuu6kU5Vc78YTw+PgqB6IlOn9nmHxpCu
hhG5HbR5Gefu2+/W9WiCSnmLNVitK2RlIXpAmRRS6fB6GhDw/MBEJ00v4ys8
MAAHd4nw8GaZRc3EeokzVYHUOKd8d4aBX7RggzWwHbS2TR74qhfeV8NJEL7u
6zNzs/KyH/0Trm+JHROg5pBLqkM1lcx9geYdBdlqmXWk86Avzek/8Q5ZA8tQ
BSjPIAc5QWhxq2AUlH/lqQNPoA2M66So6ZV9QCB7e31WTcvIQzpWFgdOjGsI
XxopI8mbn3KAJ2RBTM/5Mv8LYvxu6O9bZ3yfzRe4+l7h95wOyMdE9zWbKfz3
QhQyKbtSOJhIiJxTcVL3LmkQAQk8nNs/6sPjxAjncI8Icz1zIHrGjURrKLpV
EW1wwJpawyCsrCgzjuQv0jZYMrHRciOyrbyB60S8TV5RW4tHFrCKrtvqKHqA
6ysy6vXj7lxmrOZxje7t6OIH3d0lEyaJzljZEXDWNfLFzgHL0foERDgBcz6/
nv2iW8/8OgjwXpIo1HxqBl9rV1H7i+bd19b1C+a/4O4ZOUpZBji/8IxrqYuJ
EC+t/W9hZXvV3LO07PdnzDf2DJGu7ai8avLoojAl6sJ8YCa55VBEctX/Min/
C92aUkdgXtSLoITKEcCxVfevDjHlWd+BBbu51KPP1o9OZkPCIEuXO4rcc521
xDEjpEV2F1d2wwAoHg+njZu4B4KKTQBjSY8T+lUMYCfiuJf7h+2IlzmPgaaG
q2ny749VDUySPKC90ZXAYDffR5Ze+A/vftHoR9I+UIZCycwf9DvnfC1hlARz
+H8Td+Ffy5i58YcWxoavuDtyaxOHwpSOeg7cID63HyYpcErQjbwm7n5e95iX
FlGfW5rmlpFAeneR/08Dte5SIfn+SzqdDGwaxPUMkcwH1EUAzMMIWlKLRSRs
V745zihs1r+0FGdzTUVODo3BC7BiNWLhB3/V0RefKKg0kIrXGlU+Q1lpIZRB
8SaUR82wH+lVcl41mak0gP9216oZS6aOhj6u8Y8jk8QhaySmM3WE34rIVoTM
9ewFZ2tFlp4O6suLmZ/OBBGP9tUuxXYVW5Llacy3Wjdrcf1X6zFgoS/AkssK
hIUy3emZdAggjyFqZ8vJUaUmPYzS2BjSI6aSE5T5c6ebgiAx+9NRw31umHKf
6UMVnQSIQicItBC5m0nmVh9tfocal+hMUJFUkL2iK9IPQeKQzR0mUN5Px/tV
c0iGQHOxTx1c/IiF9SICSsjz+7sjgUXvuCD+6Tuq30BLLTO97qWrFR7gH/Os
S20Jo6S0xm1Bm4PebsGkJPViq2r4jL6vzXLshF6DoaZMYmGqdjkPAKVQq7ZE
2Qf/Kw50YvG04r8dQRGdFu8RdZcni6jVcelfZA9TznR7AGeBW1usYX50hi6k
uZqms3YDRESjC+DvpPUAeYwpdsWpsssKJxy15PZcaOLx6V1G51ogFm9+hQ1R
nEmTdvQit6sR8/L7rYMJd8xGVi8N/uHQ9+fk2qXepf+fw4HmIHvsr9dJmNxL
BTqEeKvvN0CGmJ5UzFSJh4YP21yOjxwcyLWAnRkLY2gG3TZAhiz9FnjqXuFC
/j5ndq6RzdVWX4rkSd1DGaZarDXWh4fxOJaTsyrjOefAvfsY7KCbiD5aQZny
W+jd8/uGFxEgotuoYcMBWC/bbIEIfcKnmpMDq4OtHhW0MTqdI7GbSKNxgXF8
oHs9cACkYHhhj3RCrtEABLxNa+ulgFrmhpw/nOGbyv5pEMMkDaJYquuyUhvm
+JJTpQbvpbtfbK0Y8VREQ7V/CUNbn3d8ohPBfyhanklw4RfeBamVpDMhfS/k
kg87ymB70aVVKoGOjY81A9uRbcSOMJlvlLr1WjzuYFb0ShHNEymdzgY6Unu6
k4dw+y1wL9LTRQ3ZCRlD4sXsh1SiZgNhfoetvoXtAspqw+7I1kWfNML4bMxf
b8NWfdDX+dmNFYsKFKFLElbkfNUUayu7g3+0a4kUyaD75kEEC8WMYNvG2v2J
tTyCIK0ZNppBozL+L6qQwCqvBDzTu+8A9s3SmHvx/TuoHykNKoQq2MZgmmzN
is1K2/kIqOfAiqIwdw/VrkphPvf6UwdALZPuzEw8hrIBgU1ayIe80x4Cmfec
+zT4aTi0FgwBXmTgICwkbhrP8t4RnzAlogyCSPD5BA2HhELBbLfNO1k5SwOi
D1R/98MpU9GKmSfr+TKubV3V2/spRReYESUxnDBGaHMojttBAd4E4Su/IF5n
MZykD+LXqYV5XiBozWI2+WW10mdsUigB3GrA98z8KOUAS0JNh1npS9P8OVNV
FrevbW2p8JQO594Q+MU7DPwoXExBP7H8uDXL4pUZe24i0Rbq+2HlyzSalan/
L+i6XRu8EF7GObbJ6cmpeMzTjR0nRITFVDkQxQmjH9FxmKLMRxKK9xAGZ8Rq
eJkUTPbskU1QjrjPT1U4WNbWRbpEGHf6CLhnhupyqerqUxapUE/0WbINEQ8Q
+ErjNKG8FeHVHDohaxCsMU5DKeKjuy+Kbuftm7iTYY10RbF+P3G7VUU4wzeV
XXetrIaR4soI250VgL21I59uuAbjqcElhCY/c4S7HTycpPyhX5cZlDLFtLzP
M+Kth4cg2dZYWMtq7kXLxvJ9wQ4cdsRxWz2KhFicfmTUgBc3z+Xc/VIYjulh
dbUaRjVpK3h8dzUbQrbKCvxb0pY9CuzZSSVqA368TOIrO/XoCYtktJpL4YEl
DbcuDwXzHnR4S8+NV0JAw8TUrnT5/J+SFH61mIgaXUpERqx/iV4uHBNpkdf4
myw8oIPu4koVBFFGJHOnmAPvpzrkvbjDRILfS+1sUrVB7kbQhTUWSHQAjPvV
LwcXulU1BO6KXKKDXMR1HMRlq0k7xA3MFLEkrzBIkZ8Iq7ArVSJWVs7DrUt+
anDvQ8Jbtoz3joLHowBg7j/NmaAsM5rjNPfWCsPaDyw142W1zmgaAG0qLvM3
9KKZv3pmaOT+6ytNYovIKaRJpCMPQm6FL0fudHCQNWr0n90j6lW1pzibNmi0
cENPVRbzulCamZj6lYzwxzualz6tCXC21xDsS0tXKKkV1GqbKabuxIdUefpb
btTlGGm+lqgP14xXWrtwQe3UY3R2BLhNHIi6fDkJ4qESACTZ1DO/MopHK/Q6
lUi6eg5AKuF/A0qbKm2CJWCbWNdeLXHF1ozyRyZcqUd1X8t3hma0KpQFvdXB
5hqgrluJ26TDAbiN0Er+Ja1xTiQRKFIr3Orgf+zuA7uCcD2PqB2gNx1NHquL
tU78af2Ltpu69kJbD25H3sBev8JKveEHAcHzNG11DomqJC/r/Ogz3U9GfwyW
OQ9LdN/Mb166T9nO5CANV9b7snYvpGWF6sfSoKegMmDAPspWc1tflweeR7mX
cCxw66gm4GX0DgxUxX+0/gVRpemdntlSU/dDAJbPuFiaY7GzBqvUih06baO/
Vph/m25pUXYtc4DHDuhbJIvTenpTIan+2AVgVrNW/T3iVHKDQjRKXouIcLRZ
6A/sUQscqZKKdDemVqhj8JHazVblFyFwuT2Ab4Tksjaah1eGEB2ueqMddcVB
eUepTZVMXvMP4eAA4pMgme8+wUC8olQuLImyHGnqDnNR0oRyNzBVJXiRd2hJ
ChCrGqHYlkE0tOXv+2G1Jr8qcj9Sp7BmtEK5IF3jPZKcxVt/x4tNdtwwKGpj
+5ccook5jnMiAoZhBWrs+prreb/ogqd4m4vvKgW65Q9cXe26aqlsEe31ciNK
D3J8+qHwN+PjqZCP/5z83LiMITAUiD098MsxZjT5/3Z06/u8sMJDHBN9O8Vk
rsmZMF1T8gCc463QYGHKPk16NMBkDQegCWHPJslJV+bNM5u1QEMvrETYH6AJ
8E8CJT5gkATUruKzclVFiv0y1X47vlysO0efSWT3s/vL7n3BRjWPUOTsSUeH
YQqPuycK9nTFnN/192Cuj7RACPTpFUJKRdt1t/44cmFQQ/ReteCnr6a3YqGB
uSTwhjuPnXWQcA+GaTsoFc9VahCmzgA+BPSb3dxud/0sj0wDU/S4kNZTZc7V
VsL9s4GOgv7D4Irp+/nvUUolsAF0TlaT/EZaLq0kjk4ISnbzbwv2SL2GIcXe
tbtfcb/ICKTL/SpW0xM66eQplwCn4vCFs9Prpv8W38HsA2TQYf1dyRi9pt+S
YNJ0FymLgOsTo8b4a91SThXJndeeqi9ODeOxMk8vRyEOGPCCrHkCcRGgmx8N
xytWonWUo/6/GHZO+B6JMbelOJ0QrSi2loI9kEe8pv/93PyKPDis0KXSOpo8
MxP6RPHw7B3cqjXMoFxiPCVlhHEyiNPoZ9Nebkuufns6+z2DGAaLq36yRzFq
qla1hLricDVgCjtbmgV/jwTK9TA4N3CfCadEN3hYbhqiEBQVl+7spPqz1/s4
1Adlyal3G7eqURb4PLQ/AjswBsBRaJyw7QwpTxMTTCQPPoWymvcQ1FV7TK9L
9M5WxF7/blXJlPlR93UmvSpjncpsta+knApwzkNtQr3Phel/jRUnR8VvsVZm
awKR/LausUlu89tzLymkwv5wS4197Ww2YQ2kH6Ecmf3j1JLTVh7TTdzjRU4O
rr0g4WSu6Nmv57suEEK2GbLz8z8808FzqAg247q0TDPBzsY59gtqCM3bfLj/
nsRg0EcXJVQIslOWe8YWHzjiKB+5hY3pZEUkVmE1bzlw2JBm78WG6l9AWh/E
ifZ52sFJ1wERTsgdm9haPucb6tt5pDIb2U4AneAnJVgUGABLGZxiIvwo/O5H
/7OFshr62UHNYVW9WuWaOkLNH0OUgh0VP4jWCbqG+6toiCs+vbn1OGuhPtkq
bjAGVFmvnJDy1iaDaMs3qdsoS6qbF6ju1LU9gwkrySc3tcNaTvsG91CcImiK
Kijn6Xb0M1RRNsu00yLWz2IyJseeheTLg489Bpecl+UXn5qihiIqzQyXAGeJ
sqJvxZ6YyJiIpT7qc/lCWw5GhfOkNU7s1mDF6/x18uph0O1go4iJr8WsoL67
sBfSdiU0VIJgQ3zPxEmQ74yq1cJ9gM+B9KRQoqNFtuSlx5s72iRJDXeITsTJ
qcAU/w3M5jeUulrQo63Y5Ug2KOGVoBDQcJuVLbyGUpk3AEh2VOd+Mw0edw7V
LeJAa4ZKwW0FXP1RMtn7RWLmnR5au9Q5QQGP1kjKybGOgo+AtRnKmWMRWQNs
GR0lGELYmSuMEp8CMeoo74zhIwTS4cPaGPxRr/HkhLuXeNC3pbTDccRPyUO1
FdFhXVNju6Z2Aw6W4pUG7wheU+aRDG/NO9yXDOraw4KwiVgSSnlb6c8wwCDz
hc80YRG15HmGOQhdoFvuOx+kKuo++sIuDQiNTs1d9G7KwV9zsv7FotTZedk0
ReoSmbM4b3UUx81FFnmUr9BdrtUdsBfkfJMd4C/OLZ+DocAbyX+t3HbOHdfe
X5Pb9AABjl0ahrpgwostRXrBUnKrq4w/WeuUJo0p9HA3j4tUn5NnimHqkLxY
HqZeIeg7Z0IoCH96xFmNwqRDLGtMXICqacQShjo+X3g8g0xk6wAxLNOsFGxB
drrkWGq86+lrqeV+F/Gaj/qztjL8XPFD0eFb0lrrCsEtbeT8IXnD5E5jnMNc
ZxDqKwMs33ESg4JpqJZRMbru6e8RrFfYtfT+R4ydm7wXZEoPYtbuZnz+xEx8
6P1k6ukP+IWmYzQgGJ9LMUgRpS563+87S7kx7uT2My5f51wM56N9Ft1jrBvV
XbzNHWYUWRqtZhtLppAp2C5bBsqE7CkV689O9HafmV+lTFkHGR7GHpbys1qM
rqxXub831MEDWU/N8kox5y4LFbAM8i+dymQBtH7XWGA+onvfdE58XpwjWeFQ
dsQ7jaIc/isAw+X9vAix25r7oZu9UUNYWz7sABK5cX864o+H+Dfcn5s9aR8O
0G2UGIRnO7tF8PYZjWoeCiB37fPywkmP/hE0sHx8kWMLgBluKm8qK3LLEDF0
YL0ERdQA6CU+dtbpQkUM1Cx430tUMye54Unty9/ZJiCmtnvzR83QHXGLEU/d
rTsXPGS4gP9OiBrVlxDv3aK6p87OWutLdivsl4sVJ7jm5ZSPMmH/bHpL99aa
vjmx9iEvOJxwgtN+LKkA3V7j3wIMvRR/DxJEgVdJVvCxMuOVqrTVm8hI1eG0
aYyLevg2mhi5zehGfykFx3G6WK1KB8qm2rMXAcffxvBaLRt7+y4PrompP+JZ
4XnyyuZe4TpiJII693+TtsnuEjvu65Sq5N+LL9mE4/BmUJsxFVAL8UhF8djU
9B0rPGISQtEKdVFNSMWochAxjKGpwO1e3EDxt4Zya4VQ1aUgA9cVaaHe9DBS
QYcDFJvoJAJHON5OK6ItyYYJDpUYUicqLqJy3mDgSvEFsJ+QumO2W15Kp/Lz
Pi4vtTIH4llwWyoPWFMKN2cRMh2y+Z1lQrWYEnTQq7bSb+7HcfVBZHSQveMd
3Bucdz68iiVOEA/NH38pqOPSvIzfA6JQ3+S+MsZ7IiDlotJqH7RAGlE82GnI
ByEiDH6GoqTfl4Co3X6qYsMwsqQPUXcYitx5pcgtKo//eYG2pRprHn0Za4LG
lCoSWI1KQIj80zcYfSQ/kL2f6Q2iQNp9ldniQ+rmy9K8OMOl3HLR9QpNTSoO
GT9geBG3ym1QppYPSEJp3OyUgwPa4pcrea/baIM7qAe3W/XTH1OGBJy7fhK1
wLnNsDJcyZS0j5bjiMxO/LRDpwrXdE5rRjC0H06b3UFb2VkmpZjqfUeQ3fvI
esTd1vjzi5vR2hs1y4mN/K9rKCpjKe9lscuVMIqmkjzhUCBObJ7sKFnacSir
a4j6X9tPv0I6uDyvZJfd2HzNG/c8JLW+7tttCJKVLwV/btoxcmAYKJZznNGC
EjUARTwl5qOMTcMN2luZMqlA3ASU21z6uvaZqXXV4CIM33bpWJWAgRGy+j5Y
IaVXphd9La8RJsiNIvkrgMa5ozUIsetLRxJAukGXPj50VgcNsb6TaZWDkZaQ
tZH33QhF0wYv8va/HoVgbvocZ5dC4iuA9bbXoUWTGyJMAtMaJ1bNL1DL22s7
2ZqtvJezSBMaN+HZJhp9K121eiSISEpG6J9vlJNkjEd6LfL5U13XiTf6qtSZ
Bx0ZZFzDUu0mCZlFviHqBweLRk6PUQEUcCR8iaTus0S6oKsSmr0hqqKZhyx+
Ko6jQ8LrdWoiwXyQhqZZQl3lxu8b+umxmvGSdlaB0v5Lus2R8MvZ7wvf0EBB
hN0huDy0PisQX8GOz3ghiqIbgQ6SuNKQEnVkslfvJqNDJK8D04Gg4bEko4oz
yjxBK4/X/0coyNMm6sFL4JezCMn64oQciSunZBav7tOw/9nPb4Itw+DGkppF
j1EOoUmYh9NFzhkrVbIZV0kij2wbnSxNPCoptwXFLOUNKt9PcHRXoLFw2YtQ
fKKTCga9KX4gNY6MqsMxQjFhx3awlPVDrul/70kp3eTJt2vVVrWv164sYWF7
e1p+mCOWi2cdD8/5H84EyjYpoXk3v+d0LMQcftvdrJQs+RVBr6NfGgBNY/fb
tCxzcuLBADELcnu/mqZvZTMq+R15NjhliB+TIaSAeGN2IVu+p/acCMsfu3Xd
Eh5Mkf5MzquLMjRHozWCNSG+9e+8YH1nQVh6daSj0L3XK9oZXbBHTjud0Tvx
dyErlkXrZam7zFPMfYo4OYpja+A5f1+kwx6y57K41x/n7x0cGvJua6rUvib8
WYhL002P4XO/s6VFgjYFVbI0C0srwGRZdPUY+PKCaZfVX/ArZdNRNsRGUbGe
9UrYApvJ83ko+oInJOQYjs7ktk+VRLXxv193h8hEecHli0xa3kz07u0OzQ6/
ik9MvXRy6p91wwd6/XdqaSv3hx9tfUqWFpxfOa2rKdkk+EJclhWXC+lQ29vB
pcvctC6Nlp5zk21i8z9QWgZ0TpebAK0oxPosx4x7w9lXMcKzOaxtzeBkWPpJ
9qU2WnKwN73u7OrmSLPpOzEOwL7X78gfWRdu8xhVCfv5OjNsfEMg9n7EdwVu
ZXFmitDhlJoTImChySTV/4PQ2NTi7hLXcSEYZFC9HD+PTOoMLJy5md2m+xKJ
kf3MlxeFZPUFzogGOgY29rd39Tt7Cd/ZaXVKDpFv22JEkgOuqvlKMUIXqu8O
TFyhPxrTg1JWyTxwfvxCQdCs+mbsQcArBApegK6qNivnjrv/5z5Ee9UNMO36
It3SDxZodfTSIPtFDpc+TkvD57vcDIPVHCml/doPctdjOEz6TuDnp1NNZn/R
TtL06JDHRAXPneKc+wu7GDsJZYwj2ZdXum0JCvtWXx2e0B6Ni4tP/a/Pv/iY
E8iEeJ+AbfxrEuWACbbmI5HZr+R/sX4TaNTZILzTN06YbdkeVfNBgquRgVrk
1d0g1P17TR4UQb+NwqD37Oqr7S50BnrFbhC/Ygag6AwbAsh29Q1GQjR1MnSs
pD+omY3hj7Qk9Nia3qMMVGCF8jcv8ZIZX/zFhb5X+Jk1AXAQ5fAJ8zWIHn9X
zq64SDS8QJAu0nBISsHnt+p4jLGpjx77gyPgWZ+ZK9boDh2JJkpNL6/3Zezy
hRF5lKaWbgNRklcIlLH8Iro+fxFeq6gJYp1PAG9y+a0Ij4gt9qIGie+iDfzN
phXEG5k0K2TTamouDVlbIbXI1qJBvnTLqcvFtnlNnZrqpWXTk/kuOOz2o9Jy
gn+wiT0e22ADhDLXGPVRvo8kesCAixEPLfSBTz3Irf3u9nvYuhrkbJRrmPgU
4rDpHdhmGQpCR0vwGImr/1O4PbD1hoydHDUiNKi8WUIR0L1Uj+7ZbHMLy6fj
yj9NpaUiZ2HGA6iGKq7whRiU2LSHZ3bUDPd7Lh1lfyarhaRzptswwbdjl3zI
2IA/NKcrpCMJvSI5uI5Np+Fl24VI9871S/KnZlNkJa4dvov/GGVYUAweOGhR
a2Zij6YGa4JvkMrbtBfchFQOLzCok0yplaK+lkTATSAqVTU+ZTvpcia5ZIFZ
+8zfhELrQUidQOVtQ+aVCBWWBnTlTJIX68H5/kLJbegtGju6J/0lM9j/i79C
k2rmNI2RU2PvRPY3R72HilgH6twhVWNvbp97YX/QhvC8HASzVZcXSxr0YRZl
tIEdnFm6Ss6+V3S6ok1EtCQYzKD4FVBSlBOm8HoztJt3R9FgNp/4zclX86s+
qZgqb3swB7jim6GPLKEC0L9I9gGeVMrdSvxeoQlFCxDOQDdOzqI7eCNMuZi8
Jv6SUe2XoH9WQYWmxc8GskkA77YGw/EG5t4hEn5ZPoDYyRzVBscPMK4AkKpx
49SZZznjM6mumtkalwYwX4iTnkpykBVMPAuPuxagtukClgpn+r8PgyE0dNip
jzq7fGJpsTodFlvFU0u7rwVOWEOhrsdg3TyU7Rpd0FOLoQB5KrVHnrkg7qPf
Jpw/m+YTHJZBr+C6QTq4CYBKVYIRlyrk6mdvzHlgbyw0Z8f+BKYWRn3c6o71
Ur4sERPniencRNS7/A86yMZaCSxGuzplfxIRVt8M4scWYWczmP55o/b9Fo7e
OPN1qntIc3+AFAcdgXxfmbrS5QzkxxHTe413WtvsmZZe4pov9RzTLycW5ZKf
E+94Ui5kHP107JaU72CaW+BHdlADMVXkvWVa0qqgjTxT33WZNpf8gxC9p2n/
Jyy1jN5ekduisnfQABk3u7ae8TOmexvZc1Sw8448MPJ4upDQdUjNvQD9VvLT
uy1uv+jLGY4ZVQcqwTmZu8kPDDU/+XpkHNiRnorqiWhNsGDLxOvIaWCB9jxD
obTFtPs2plqK7YVKmcB7V3aA3cAz60p0T/SgiJrQpLMeAUPXKVIrBW4dqmVU
FNVYeJWwlxaVm7MuaXev571mO8C5bpEkOZQbkN7ZyJfv8yHTvrxwVknQfKT6
TlHSgzHIxLx0eiHztYxXuAv4H+n52RuP1CVIURugeJ9hTLceIc5Aaw6PzwOE
dqO0jYrWACnxdXS6Dr/xM/PVkKez+G+F/uVXu8PERXaO/OYmusqCWZez3ELG
qaPemLDAQJ4+YWp6c+k6aVSkeQAITkwhktNBpFBMsFy6ay8JCI2SWxVQG/Lm
ib2ZcEqtCU6hLvNIn/sqM+goAENPIl3pVnymm4g03ntbZsinFdgHMISm8pTN
A8zBXtoo9/lUn2t6qJ16e8VkIpY9+Mq4wwPJpRujNTo/BXHOisiC6ugodIcj
ct8KZsSBprnMGzyaoikGinGMTTnNr/nfkQ0EUn1rTDXQsC9k+VeEJjzi7Fch
x//vY+o0x88CUVjSGAQ+whu+eMteDzvfXm9PlRgz+rGhY5fm4P9xRsHlzx/4
viJs81xQUalG1na7PXz3FLMpt7zV4BeY8FFKAd92X0az6qh3iGWMtScGvsq7
pFWfWksKnKKTfWZ4Cy7l/EQF4utosFqVNvz0L+Yyg2rfA7I14cAFETs7Hqhq
1xjQ+VnKf9um+r1FJBgskcUSOW7NEu3e1TRldaPjJXeKV0/c5mYbIqPf4wcy
GodQQhWskssBX0Y3hLMI7qvIArvWG/2cWcCeQFNLAtwLQJ3qaS07DjdxTvmE
ZUBWvH0G3jhCEUNOml+0CuHNdBt2R4K6BU5LBui4OP0TJBjDvyplAjclBDOp
rwGTMHRtEqc0hrgCLU+Bnydm3R1Nb3Br3SiTUlnzwZ79L8jbSVGh8Acp+7bS
lblg9eQA6ytl9MCvamiknAJQsiLhQQ/jduckCU/h390QHn8kYPASGa3Vr8Na
PDcsOUv0hnvi0VyVT1HI4l7yy4cfa0sVpL2Co0af67CpjKLb6D72g/JaZvGH
dLWNDmXHIDWDA9KzfZ7Q0I9e9nulLy7qKDmGmyl77DuJnUQgFbPu4hCAdyYQ
YcW01y/DJE9h8FoCjorGSTaunBbHL5QwtqQNIU6T4rI11gue9N8cZDS0fTgk
gsu/i5i/gEB/E6uz7mEFNIsXld01XSAD0woejfxQwiFNAmekZ2C8J1XYXdBe
ySe2N6iqmNXW/P54R4FpXK2xi50I/vmh9fcgZHYtM1igUNb1rxf/A4QyAye6
nLzat72byWvcDc0XS5A18txYZd2axE8/acRbqhI4KCYEQgP1yL3Y0twk8TKo
TdSjcDQ/uBfT3CAIZoje8bTE8q/MzYxHU6niR7ppx83UQ5H08ytBW4Sf1j0h
S32JyBEmLb7iET7+w2BUUF2GY62c2fT21soH+B1ADN3/IG3ZHhGBpTrmbOk6
R80S6FB0VcixohGqRL0yXLmSlh9r6XRfJXqpyTgmUJuB7CZ2kOJczjVUcC58
GxklFJ9ZGQTphCZNnHaWpPzLm+Y7T8v2CdqZ5cCmGEy+wFu5AXoFSL46YCxy
JHnEhN3kTnHCpZqOTfZsBodnLg66G5KlrgL2jBA7RKDlBodRxQjzR52kZckm
lWtAHM3Vx+9L8pVTaevFnlBbatAAIGJsP1dO2NuOFKQu3gmoTTX/05+ttfUv
Q4Tkd3VWSdwwXkalJWi6BbxlSVV1idKsTFMWlwAFuK0OUq4DG25Zyi+5q1KB
GVPZlyP1nhzb+dzQ06DToP5+eCLCC91rN/dUrxghK7eA0xeXw0cM+5uVLPbo
Hyul6P5zgXW/PCcebl9qjoGKUGfCEfdBq6sMZSzf0L+UEel88jc3Lo3xJ3co
y5jkpx5e5rKA2fZqBGt1mKwePuX/6LOKRP2zaigXiulXWVQrKIDPSSSEp+Vh
DgiptLbV7soJ+8/u3lPAs109Qac9b47Wn9QC0kI1yCdE6FMaEFtnAtAQfvQc
Ws42xqrQFLCHghshCqH9YVBwF5MCsj2ygBr1JUsqhDUSSgBK22Tc6VN1ryLC
onRXBqTex+8fZk3Y9miuKt4TAvo7OPycdFQA/fszs3Rk01trWe2dnotA/RDt
2eea8Ooh+as7SRPsp7WWaifrOZTjGXoF3UN+NyyHYX9I3DMDDuzoieDrrPyq
Oj04vySR+Vv65itlTdXS89ZPEOAkTkx7aE7N3+1+RmS3cag/AWf6SKrYkkTo
ThRl2uY8Jd9gbE7Fz9CY3Gm5hGgFDdnSjK3CimNbm0Y3FLceHESsUO3Xv9wr
9kSH92lF08blnu1I/yWjRPljkITXs6HDrSg7x1wRoQQGsVxmZXt4BfLVFgcF
7G4qhCfeVMQF5PUZOVtCJJYumw3Ge6iF9KF/FPcSR3x1s0Per34ZVlzzqS10
L4zBNayIJxSRMJ5hfsz29sEX6XPZvhoj1WdCqtnG0HRFKDnIykHfeuBmCteg
D3feYHlQOP1vkgeqTtBFoytRWteWok+Zc3B5+IJMlvuKQKx+kGElyBWI8WJz
q3Wwf9OQVS2NysusLYSLmxdvEjSYn3838mh46NaIVROTXhSQRqu3qllv0dYy
kGAU3tlwuSssSCaD8p6HUwkKuLSCeKyatzbOsNmysfd3wFTep5Mby4w2K+lq
a2TIQRPzyj4d9ZAlsd4ntjJvBw0jXUjaFXxAFb/zEfBUTqR0mHa91B+Vqq46
sNzwW4gLtnm5yvGzriFg9QEm4XBt5Qa6N3kwOK9wS1+EpVwtBkiE76AWapfg
gOq6z7lBEkqk47yqg38tXUenfmRAzXCumaI53tQk/vGmV++YlhyqgKwyldXT
ntOT/boP108Qa9vFKSWUvReP3xgDxjjDzF38luxV+NLxJwRCavmSXz0T9Skm
gn7aMmSo9C9ETTmWl0Ic5eLJHwEL4Qm88xhu6OgPfA0o4uWOyrdFGYpw1grW
NRjOKahPvL2j2z8TUMDHd4RKKkOv6SomhqWmaUpZwdv5+K1pfS7sg144rYMq
Wa4Yr4G/WkOyakrx9imNVKq/ce0HHzeBuANR/nzp4xWLbv0A6w0w85WbLJUy
oS8EjmRTkQ/L9D+sLpWY7rMwlqSfFQDn7w4uXt5svuQlYyg72OkHz2WET9GA
+W7STJY/BrOnT0DSolKmRYaUa0HVRKI1PvcfACWTRyJTS6gx7vp4YvRQh6mY
YV1+M3E9MXBhPp9EdK6fr8No+IuEKRKQEOaOCpfc0tgFhKIAForbv2d+Fbt5
D2KS2FFSHI0hlmeEpESHNLOuOezaADq/aDkI/PDmrZRK3e/lJBvQKU96TBIf
R9BK+qY0BmAbuRvl5MQHBEFtn+UstBOI5KopVydC4qKOXRveToaO0D6Xdeyo
VPtW6QVOwVkFiI5bXZOlUXXwmYOQq1MMh5TaZzMaRKlVmJECO4U5cevxGxql
af/yfbZ0g5hGzHMjQP4XYkO97/WM+jqYn4gqUBvwpldqrmsqp4eY0JlVQ0TF
nl+2J8Fmvp1I2dc6/DGq1g6wwtV57Hh/erNBVJsDmhPeICMH7FxBycEqDcRH
HRkvUKbBOg+RH1dvGn0jhzxDTT2w3BPtb4Bfpu4YW4JLkiIOI8E9lomDbXbg
6SW22a3vL6cL+al3vUuhTIbEdRH8xL/U5nEYGTh1kd/GunvbcRmui+KBMHZu
jYjkSVlHMHdmX2ZnawNPwacSU3JFzf1DyVHtkzZz8ZCKcjA85h3gqphu2GJd
DZi3dbEy+O4TSPPldnetsqNLA6r1eFrUlXXITbssTZDzMOjXzPrsVpubvspT
j7F06aqNPFOsK7kl+zPs4ZDiV88+inrvqKYXE0WvObGTj9f4fXC6ANy6qctU
UT/s1HjRmX9oqYb20Lm3R7O/Tc2keKfQqiKMLg/Li5hQue8Hc1mu2ZpfrxPf
EpEeQ5ZnK6cWIU0uxGQ0CqxhTboxQGV/kiATeTfdg/ccblrYXLAwwKppwZkD
lFTwuj4mzBuqzXowZOdnwqryG/nPgh4L3QeRgGs1eUj0opr1iRZ7hZQIw/Al
X2ueVp/oSXIvDkYtCwICPQ2EA19iNOZ2QqNEXqQnAgVOgAcvRLCoRct9QQQ0
FWhvKlRg4/IWxCtZ1jO/u9KJomuhlk/A5/JbVa0eb+FZUHGSVgEOuvUjKztR
I9nhGMEjP5M9JRbfCz6sUVvMaWpzwaNvfrvHNkeFreHePPZKat/la6KtkjAq
SgdsCTQLo/GAHCom+9GK+JZO2y0MOIfVW+92cmnKBNlqCAcixitPF78sPyh0
IPpXXV88k52sRQBwzC/SRlFdq+SJsp4YjgesDsZ/2Qv78tW/wMDjiGPv0rWO
+mxfh7UcRWI2/RJi/9IYWJHqV8Kw+23Pdvsi83KvNQacs7Qu9GnXMZM/+nr+
pkijp86brpifxCG+85uFtKBRiPkiF2B9p3FKP3Tl5kxkRUn7tsbSXj03jsqy
+32yW5CmrPqZEII/aJDbSUgvrJQmgM4/8W/OnoA/UEYv5KItZTspOSRhYzhS
HTCSzd/xKYv7BSgV+BDPdZH70tdr0YvtL/uT24tfvm3nsp+WePLhXT9NsSYM
Yw1hVU0KsR+wIJEvixKYEXwGs9iA6U/EUo3xmYIyWHyS/R2ACpsQyHp94e59
3CHrluROZ7R2tGZZ5EAAP8MI89fiDp9LbYta3FwLYMIfLI8Ny6aObr+FqSzN
j7kfR/HvpVBaNJOMLZGggIbthyl/dYAAU+PjSFrVb6TZK8qqvcOlhow++xCB
ALv34++pFbeh7oXEcbdlm86cN8K9FMtr3XMYhphYL4LOu7QzV954D77haMY5
vbTcNyU6dWOE/qr9+EVgXdcR6njtyyc4dMrznteXLbClRLJMN4gwwFiIFyRo
S6aj4qh0CJmUibkzoabxQwz3CGFzmtdPJpEIVmL1f7eBHxbuhh0IgXjf+KQf
OTaY+lOJcFzKtZpcsWLG4HVywsi8o5VcXS7rMAsw18wnsOZy/qtxEb22x71Y
sNtl4ALPaOK9LrDMoNTEgEt3Osm2P7UtQe/I4ZpHA7SaCm8typqQ/FV3n1BH
XBuL6EmdZK/tRdEWUppo3irE+BXHSIhTucxN6R0mGhqZErOpOOm1RGkfRxRQ
3QjFAQ4jQhhYuAj9E0gUnNoRtjuso9823GBErFOqXsJ17yDkEKnYL8K1EFVW
hgSeEXNnJv04VNrNNBa7ys+WY1ocfvwKzxwB0M6VOxii1V/x7wel+33LR8uI
OWt50eIO9ncQNlPlmYfqhqymcKOBMnd7OtCnywE5s0eIQ4HBNPi14jZswTHP
jSrTkWgv/aG2DSmbPTilMeH+3AfSLITIaC6MRlWFckD2whgL7Svg7OkZjCMF
AoGIHlngan6l0kYpGWD4NIq8JAZLp2zoQ1xT0UD9s9u8WSx7a3o3UXK4H8uZ
jOcIoQ6lUvGIUjbI5fP2jDofNeK2Jh9R1BS8iGN0OAfITNI1na4QLFMnRAPj
/EZ89kqKH/eZW1B//lgEv2jbJ7uGpXgP1COafF1A7Cu0rpY03B7qy7gJvwrL
JGQsOjx/f6B0vVEu5S8fVFrd1o1UPMIw1df3CCGgpmLR2HamWW/7U5FYbpGn
EBWWkb17bUhhXjCnXPIs+ocEoOiTQyu3Gk5gLh+dxhk1J48i1Nw5q30f+6NP
9ZC3eJAMxSYiycBj9Sq41IKhZMNOtz5L+0zPZQgoy0l6E6t6NG5LzJ/QJjLg
uJsmH+3cISJtTbO6wu9OmzYsR20G9S3HVpWAXrmDK2pGn9qk/WHQ7FlFqaJP
ZRQeXTu4IfVask+L1/1pgEguT/0t99LwPNCgB5Vs/1VjpVYEGRxS2YEGEvNH
VsMn+ofNSLXCWnZPd5LSAPL9WABDoWqajZjdrekBdaUpVEzhSseYSAKuTLre
vp24KE8fQAY0hj2P9yIvdKyNhyT4DCF15QEAQ10itqNMxl+o1Wie7fvc6ZNz
xJLRqX5XLRgCn4wdiLa1PCFvfkvYgWGqG6d3lnekf7Lgo+P8FoKi3rqJydoB
Vp5cVmMKDS6TOSvIhCJ+bkMNju+cmPG2Qhcabrz67vwRq96VAY4Q7VTLtb8P
lGpkIoi14OJT0yzQ5ntsw6HRS0tNpFYsqETMXiL4XOp9mIh7ZtRny6Q3bjl5
+DPNjz7ZEpFDsdi32V1+y6Q++cH3DsDGg5LFpBGQZhfdRxUw+GydvUS/v8wN
bicwso6y9Oq8tMLdYMXbNSlKdvE2kR1WOMdqGGhYxKUhLHWgo6E6EX0UjrZn
t4WvLrNWfkULO0k4+7PLXnTLgrBQQWP+RNcTt3OcGdj8MGjBEq39t4reNbQ7
/KqDPOHUgq807cp1QsMfAOa10FoP34vNvAJrS5h1qMqZgs1SXn3Ed+MRdSHq
KIClKqosWjojlqgEtZJ1l2TdnEMoRu4M1QwVrBUe7bKiJp6rzdFCzC4DaZer
jQ1b94bAW7U09T9MG4PhOxHaTZT7SMn0ciH6C+oCwJLXSBpnDXt2R4MIrsWy
NuSC9waCTFNt25PDEE0TgeoYhz29zbUnz9bVc6mTgbycmF3s8pRUtb7UnRap
apovO9YzMEc5YCPhTqD3vvpwdS/AjDuRfVw0FjIga/5sdCiHTosVNRqpIKdd
na6OkCOkBMN/0A1ZHaqRnFUbpqhMhOObGdyeJz0XUnhySxhvyIaQE814fmXL
IcUfaSwmhiXc+ptivbu1WIw9Zp1E1xQzBc7SHxVcnKwi6+jTRj05WUOJg2vn
YLBk3mRLIp+Szn2ethHIG6SV6mlwKie2mIT3xVXRP82gBbydNLyRv+eMlt9S
uIIlHTKn16+/WW+xg6caJXEJ+bqO5i0+sFm+Sdmn6ccshqreSS2QBYY5PLBU
nGSehPAktohbPyRQmklidmqzaAmrTnPGd6swrkV0Bqnm0VSqbACrQDZCki+Z
ePaK+By1GbmgZJBqdLB3QtdAA6MUGJ3vbmOn+o3w8ZebSsKUf01/nrg555GH
SYIs5dW3STpSJGLyQTKHAyP7EPCfxNWlGxTthd5y8ZGCbkqcVlwpcx4P+plc
0n/BhHb0l/O2fm/sYuCReRG38A5+QAU7a9tUb9od0pIFE56cOuzk11D4oG2A
ISrQ9MeK1tYNYGeTKyJKj0ssDhlE0CbWijnpeFttufJHR7alSiwbyWV6cfIE
LRtDGevThpkHl9l9jM25s9fYvlzRu9hLbex11UVkqp6vAtJs/KKmsZdWpyNr
3xEl6WPv7P/lY4o4NXrL3eTI7rXW8pn7pkdjRZHuJXB2Gqq/sZGtCBqgIj6h
6AOtUkA/eEzUCXS3IA86ZvkgDkcPScqrME65vej6XwAt3zoVoGnsM3qNxFsy
NeVUgjp/qDudrJW56+62KVaKRBR5ceooLbT3hdm7k58riTIdQ2eP+6gpzgnH
m0B38jfrQ1KYb8peRHzrbDFfOfQPsqrO/2g1zwwP/aIsxje+zqAy4laQfwzG
R4hyMZYuI5zLj43BOaw1y4xDwrWnrOqJELe2ZiGYCkSlnU3xZgdcfY6ns9sm
XJVafW5c4T6HygD4k4+IOtXIb8QAMfzDF915HbBeBVG3PYU5KENe5ufB9urs
wO0ti9oInBL/2Zh61XmZ8POlxg+zqB0C5FBaKQam4FS2ZIFNM+rSazISu8OU
IOh7B3TsYRPi2p0VwUhZfHYyGdZnP1dWyIJZpB1HA8M/Jg6H6NqvTlntnCLq
JBUg628r147/QSd85wVGJvwSoS+/tVEwfQK5OG4UZwkXDFLmDHDWe0R8ohLE
rBtBdfgIqgsZKMDXt7P1Or5CAM3BZYfE4NR3fsWGiVN/y+vLQ6VivUeOmOlI
16TUmVQNqJan+BF8s2IqLBxGFvgoUsEstaU/dI9K47QveX5JpzgrLg8UUeyy
UtTjtIKBMIGoJV+ieNowMd6ueI8/vDpjIgF5hUgNbM+NMPYPGZ23Tt6s0ZxB
J1NaaTz27YNZJrcKjFrXpD7PZL09XRLEBfINnIN1nF8fUUrhXXxdBH9anA9+
0YB3EYqkhFgYRuTYvlz7VXYsb8D61QM7UvVgkaleX8jF5p7hqFlkkO3a4mIQ
EhA1GBIuJRtB9nn4Ur79NVKIve8OFxp6O3d7nnBMur/Sk34OLGti1kPncaz1
KdT3JOY+yc7ANHWImkaxCniaCpFWzBPb5ajPG3YAFI835LGzAFLtNCaIIhYJ
L6AgYAaoUMBGn5U/bZ5e93CtHEKQS8F5taJRcFitzd1hdIM3unZXl+H5XDns
8nBtdmYId15/z+QTg4Bd8F4v9I5iGcNXQfDzlT0ihMcTs2u6XMYuJ/fXGeFE
F5fkPNAn7ovHTp9AnABhZP0+yHf/tQZGIlpL1fQXUskX3plu27heuhPOKzC+
L1xiZMNKkiMtlWnsTRMf5fy8CwamIPGzGjPEvPSo+fGOQLL3bM5PgTAyJENG
sLi0pj8gfkXAJK7QLlOXQZonbqhFsf/5l/GZE7ksoeRLPXQj7GZVdwSdgBNW
vO6qRGKu5gWahliltZaOP7CjfO6/9SgflfIMmguBY6l7mmLk5DKAEisitFkc
awKnbIrywe1DtxfXELcm0jnJdDFJAwB7dz4gU9lImyIULKVJkBdnuD4CvviG
caG75CDas/MaUPGT1O5MqtVSv+hRyQ17pBbLhCXgdpKkvrq76O57zfAedN0r
vf+kWxgj18FIIhYTypoMsWYQ87czpfdUZA5BQYqYH1W6FYdcFhIkdKjC/WQf
ydM25Izs5kcjKYFMNplOOqcdAW9y4hewZskBx2KJXq0GtULhl4D5dRGwo5fl
+UDOHYxuPl4dx83tNqRBfZX5uWrXvitza/1KX2EIckbdDumpuHjLmxo0M1Dl
t9+WZMsVI59gv9UR2//IhtawqelBXzGzk7AyAHoqsgmT9tArkCQKeG2dDY6N
MXnWx3WacU/Ppwg/umeAmBW4gdr991G3faRtnDFixtuS0h2TC8u8a0BWAOUh
xFFs0/j+/Jx05NOPzihAs1nm/ujQD5rRtYv7rVaYZ5HpitadDtDqItPc6moN
5LKenf1KCEpvLLkoQg3A7uZHJpipeO/j6Zqo+t1drE3H2TCd6lloC87qCT28
kGt/BacbZ6l8IQGg7owM1Zvs0270HchOex9zgDw2pOlgqaUKtt0uXXmi4F9k
A0+feh2KvQICH627l030yFBSMlNpwhiGW4wPlQHoh4mAYOFxuRPhMeJWlV16
V2yvfyHo9Om8ZeIVcjIH/3a5Iw7TA0DKW2PmzuueLyCNhvc1ZaPH00s7gnVo
xoDT06Rg1WsVL/IzJcZRY/UDwcSGPpKWSisNSCec1lUgwHrCzj6LYoO1F1bM
tzV7TZJWaX2PcF0tCUNtpTKuzJE7fYUa+r2vbjV7II9fjQAeP2oN5GJoCYNc
ZD+rIvzJeEMKKiLi4MAZo5AfgM+aJza7k2rKDWKR1bX77nQjuzzTpdPh728h
a9Y+zqy/DmMfGOfXKrANqNW6NX91EBIItAKPyUaU106W5p2zIZ0dFRFCxr3o
4WBxBR3f7wCM9b2pudaOa0lJD46uZITsj/LA/PPGfKvtJ3PoGlJbeXhQfrms
PQQPwZxdQ77zVhZxibHWleVpdLh1Dz0xamLX72Kfg5vxKGznldE4/cko/DXy
Z0jCJmI09RwHvzlkt/DPA9JjdkFWEr7yZz39LoqQMdSJh49HdTDK7S6R9qSU
KfyrQO5u2cRHGQg4HYv8EvECD7/vQPk9KrkcysrdGfaBq9ady97eIDg7VTBz
aUOyouoq0t98Sbsyta1d/Zdn5BlTvHJR6NQHPWZzR5LMKYKrEq6XRIT2y0ga
ciC0kI6HnlK0Cvg7n3XotKNzPERkfaY+WkqHN4K0sOq22RMCnbtQS1X6v92n
ScGYBZyqhfHOYugxONut2JlJB4R/OQhbDdAvTRq75xPrQLqxmaz7Npt/AiRD
CBAuBpahJbdlCZBThYlMz8jlI0loeALRIWuzcIocyJQR8Z9LqyfC1aqcNbBQ
8pr4T/2K1NgAX9DjUlHNaZgPjC/DuafreM5pNF9yRIBZPnNPqZrfkqmjPdl1
rMRQIunT4RVY36894MJQGMg9yzGb4Ohf4aqCIGbXHN3pDUqSLSdMLkxYkjzP
tMdTXdFd0FR8rPtf6T5I2NOpKYXQ4k5rzoEbltw6QH9jPwgJviQghvzlK3tU
cA6alk62pxovXp56lTZHqWAQJtyMXXiVXt87FbyWjoNLxSoL4o7GxVNS1nfm
kzPigAViwnrUKg6rkEMAdBE3WXg4sNvDptpiqSV4r+L3Sdfrz2NTh8XPahjH
zZcx/F5a2z0xApfJMbFK0fnYOnFRhMovQReOV69+OGCJ6XFu53NHUrqgS4Jr
K9g0dCiRenxTaczfPChvkADzD9IHyDhEqhyCb33o164QrhcAsSv+xIWPmZ2I
qL0qrY+U0hSWTeX3uieNzdIopVwSofgcwYcfiaSPpZ1qzMQKxqdDCI0h3DN9
RxykhsRPlJw2NVFq/kOhjR/ljxrUIZ2dpauG/q4juZHsscESICDu78g/cpX1
rvqal3JFtklGzM4/zt/X9kQfzMGkSJZDGZ/juVHbNapjPqTNvOe2HCH9VfaL
oap6E/qPn3ALN1TZ25M5ksg3Oo7mzEeG8qAwiVSjWW1Zzj6KeFFeoQ/IyT4B
75D9EcWqt0229KrXuktkvVI0fRPP0qyA3MOzt66I5mjAEZMJsGQaKpI+zEOo
H1oJ/Of2z93cV6vX+6RC49HIRlpQThS+sEEgEkNyYpMn86kt9OB4x5cT6KOu
/4Iu4ibUmFG6x6BwicCi/QYR1/HGQ+cCJLexT+KI+SU/w0z8D1GisLwswDMr
VUA1tTqfK4YGOiQcm42zLAfQIdt4RWbT9B73JLipxiI/w90C55QGuAuTUag0
iBfTqlbsHGtDnNSavq/dsHYl/PlDL4UcFMEuqi2A6QJ75MU0CcJ/DK21z5Fn
KNFECPpeSvENP8nWnfzWikXcvmEqBcd0L0oAPlPgxSj68SXfX432x/AP1LeO
jgihcn3kaFFhMILbw0BRJDM/YXN7dCp2StlNUBIBCfXAV1mUhsOv88eWpNhD
CoGLc3glc9GyN7Z1sgZQO4k3UycrfElTk1B1WB6n5fQ9riWZ/e3AdJW7JPGh
3nvbvh9s4+dX61dlJCobgk3j/4G1uXHm71wDcmMq8nt+Lye13n5v48/GPvY7
A7JZ/Ys8coshPi50j+qZsoALwkcH4dBhjrHzcNon7Q5Oxai2LKHOIEk3wDFu
kQw/PW4aEMKMHXVphjvpbWMgNqE8ihVUGBB8laZzsC/l1guky5spK52jV5bJ
SjRMMl9xjhS3Ez+4nnKQCpsIXvI3fseynAtS4zxI1rKVUkIppURLf4uQ3fRv
akWX6haxvjfhyFIhlGKhPRJS4LQX3TFZW4b8jtBgW7nxAOXTzQs5WWhTpFae
cs5G5qSxcHIbZJ/fmFN8TU8sHuUQnoZfSs5hr3PPw+x6+DaXbhay+YVp76/C
eseqRHvuobMm52zwhdYUrIcDidUFqdxbF1tExYNzpxTi3CRtz/3rAumhdZSy
roNMuq3nPFGirMo0NE6K9yG61sd7mHWhX3HM7jrKuJA/D49BWOrIbNArF2SL
wNiYB8AEcl4hoC6D8+pNecVdkQ/aoG+eW9r8psDU+nd4GET5pHcKM606L+WR
vOwj/4ixpu96VkUqFHcNL68Pux5xOLzhrP3WF63huOZIBD/tjP9+NzDa5D/a
mcBAcSKDHq5HYN2iBIY7m0atSNuEwp21Pgz9vFHJe3eAu6ftmm9af6NjF7a8
DAEfaq/7f4aFlI/VNU25stDIJOkNRkI/WuGRzVcrEgzqNoO/wzf0u+dFEOeP
nttBiPQ/9qjMojmstIA50WFIm5R+SaiPHIpzx1NSErKsT88d5vPNNSu30LDA
FAtKI9esUO/MEQIPfNDVJg0VqwBJYRDzNlbcmLM7p0T9q1vKoVp3DNoRZqgE
fJWidZAWXkU6eGTTmh3u3RVfCtjmU8vnYGOERquDU5aavHMpuSc6Zc3lZ6Ce
rSRH8/qkyWhZD9+nOExuxQS1PtL25Lqrhu47zdFQxeoM+T/2PjRNqFF4Aexr
nnosdaRjSsqH+J/jsMIWxPsB1o5TKFEOxPegnN7mz687KSlmdRHbPGmYpZTe
tde8jPHEyCR1q8aET4Wri1dHMuWapT9LFyQZLMX7k/p0es+cnYYgag14NrQx
jpvJ4COdr3/S+RPcjzACPbWVcF8MbOsa3wGWb7t/AsdQ2nOrjM7RSF/VI7a2
DivwLuVxv+DrZ6koK3kscptwJqCAZI9dlhvxxMxhCH3Q0Cgosg/Eb9iWX+CB
83D6gnN459F6xb9jNKUnB4wipezVpAQivLMg8sWl6wHuwupkcqCZPkZNKCVZ
0uTaVY+/oPI9DkketivNwowFXXukHqtbiBYy8p2h3SlxA8Yr14foc/Wkt1JX
PQKe5xeLk5EBBp6+/b3hQKV2IjLXkTGwW7SzWtyKmVAyYWz7toRaSqJSftVf
QqTdKoBZ3WfUlGG01dFi7H0Kb4sxaXynh+CzdKWflPT2B+tIB2ZtcTtUTXR/
wj2CjCXV59RGYtHf88kRF9T1ZV8Fo4lF/KFU5QZWZrxH5CafTrNSV9Ox7a2Q
oPu+EYu9uLBLzGcqY9595ma28m4kRmtkP6OnJy8yB1ZlYpdYi4jacymE2i6Y
jOW/FulHf8AcAU4xw+q0jmVDiNKgdFZ2kPFHzRr22i8Fv8Om9kGbTgXLgBUs
212ka8P4eQwjzJUXeQOn0Hu12xkXoNB5OaU2RxWALf7MkJghhszba/N1rxlp
Gyd9nMcp7SzsGwafBxBrDZGtfEwJ5w5exufuXyqj1rQ/IuWUI44OZ/YIyoME
r8iQgm9F8qf7u46zvWprtybbeg7T2LwxLy63Gaq9+jrOPs+BHiDQnyXPZKel
g8lngoKBLcYDhpruJHZ8yK+wHMhVckkxAmdffwHzhoH1TZpxSz3a1Xhux37g
0p45O2+7qouwBlDDXlsqmIhWTWLmEW9e/QmImjdPmZE+naF5wL/Lju59xygp
qCDLrrs6p+85raVYOjo8madIqQ6E8PpkYCb6XHc4PKT9YFpzmlEIL3Nf7Ek5
/2f4w4v9ngbHSZEbRdtgOyrgYJ1pYv2XHtv/qOFv5biXK94teLCQkVAcoe+f
sOGUpcvsUJfgDFnLVjdU5HfDLruMkfIGLxyQyvKi7DSsBTdxHVaALbBblosE
Hy1/OJ2H7gv7W4p2RxvDTWJyAQr6V4qvevvpwC8uJAtOfXOScOZIZ5uIbmnO
bYgajt8JbftPzuuWgXqXPwBxUDoQSPa8RnjSgGTeEV/l9fxSPP04Lr/3dde7
UpAmGP2ZBK6i1ndMuJLtczzIUou+gbXBc7f3OC6IVsXaUFDpIYp1lk6BnPl0
AxohJSz5m8z3UmpPEqBXWUPcnJ5uObJl8Mzirz5yQPeMgGwIpcoTpz4MpBVe
IgiS2pwVvKhZYKM40t24Aqah+kx3jna6sxjqrt9SxOBWzL6mPHh4d6CBfPOm
ErcQuIvNXPV5FSNKs+JyaaBmwSYFtfgCKxT+3hMQSi4pRxoiC+mEtgl2/Pyv
slmiNzPO4vxvXWscJ7vZKBwfvUM5gYKAh3GOKX/HtfpJWhLExpJh/Ldh5rLY
b2eDOPq3UN5mAotEfqnIiZRLPv8CuB6AL/aBlzRdDNv0UD35mGgY6qOeOaER
JW6kG6dnVue8DSNAMYYY9Iv38sxQEqyiV08uphh8FUqXyNpT22fp7As8BFnM
Havqzb1B/kZc8RfwfSU+CVhdohlcNaWI+3igxk/TRJvK8lYEnoUer+6pMmKF
M7tICjxchFLLUmHRCQrmLO5TSXagyt8YzUXdSEBZ3nKwerKBgBNsrV0F3rUG
l+c62QHEd6G3/u43z81V4Y41LckRW1YvnNgNUEv5t3cOo5+rg31763T31gJw
Ir0drd1Kas+axU59ztdg8ElrGdK/MXaGG1kyOpVZaSZ9+uaDNokLLXxpWzKO
vb/QyRxcmk1ijhHZmaCeoxbUjefKoFhdd5IYb2D3ijge0i3jix9r0dcLi26Q
iOGy9hSQKn9gKELtrDbgM3JpGbDHts/j8zi1TQu1MoZ0LezOO/1b1wHiO75W
q85eOKqoJhIwqnu4rRYCLsT3g/fVV/2j6O/K65Fv5eLWi/Gm+mYl+kn65nrA
nUaOLibFBXPyCQLc0hTESVBSJkEOvmSGGUQMwN5dqRQqSNhyKhrA8Mytzz/i
KoGwRTw9BdO1m66aaR5CDWb2eVCe+Q6RSxWRl7B/aMrY4tfoWn2IZBut8wOq
NyIQuuyojqwNzJuKuc4elukUXYFBGPeLsB9KOrqZhPHHuslsdc3u9Myy94t1
df2ce8tAwy2/3EN/3HNx3/z6/ATgCHq4hHn/oiUs0C5nmq51j+OHL+Qoduba
ApP8dxqoyPv4rdJJ4hne8Vf1gtgPMmPOzedsDFkzX4qwf+PLnQNuH4KpdT+I
/TSXKoLzyLKZyZeyUZ60aiGL3x2TAVi1KCaQo60wm/mhXbl6iS66eFmH6b/k
kqwTQL3t4NF/v86Q5Djcn5Wrn+1mFBqWeX3JmRhMthgrwGYQwHtKWf3uvU7J
MnH0PzqYCAllMx3Mtai9xIE8DsO73nqw5bJSoG55Yl97euVNvlb4so/fKi03
AD1W3rbUrbNo//xk0fuWGH1bZx4qnd1rJIaNTD8WiuMiiVrQhn1XlpoFs4oR
Ohrl9zWLqFfG9LaT/QuOVuGkDbudMsmDwfCXRPCsSCmj5GmtdwU525d8FNp/
UbW1AQZClN8f5FEp7rL+yxoO5iyye9plk7BPcJFLxI2xQxSyEvOP02a8CqQb
VFVUQ2QunvsWggt7WplTlnJlr90bvS34yhqH8nAQ3iElDc2eY4NsfwyrsZuS
PLaKFmEOfhdUB6lvQvyuAYb4yXz+nK5B7o1mDjDDzyjnjztjEkzRyBWQ/gWL
gCEKk/rw0lzyNN2T4LYnLvwRZ8yocgD/SuNtWOUTu8WN/8+VVvD1VYnDVAPB
Z2hc/pk7gQmqH9PntgcFISTSnplt/cYPNxFTOB73GPlrEhLvMtPhIX3mG4+M
/CG8PcKZewgDRRlQbvWpnlGZgEY7HM2ZTonOOqk7+eGhA5g6U1R1dbTsLcJr
4gw936ShwTWG1vkQectBcfjMan3xonyjP8lCkZSRkfOitz8so5E/A++uNurb
GwvjNAnVUtBvx3pG/4Fc4ywKzvheLLI43gRN9mvAd+dukrPDLE58ZL8yswMT
Ki1DK3Dshvu/vpgb9ZQuHWM6Fr0DbVPW1Y3bCjl8j9H5MFUg+W2TzsxaRymK
PK7+f0evJy724yvPcRJQiJgoTyDVN6kq2d4Ou8tgKaJhPKy/IiArpVmsUCoN
OIS8mW2aHYO2k6x5LCER3dS/CyOmhRElxw4mArUNDAOKQD8R2aHU/fvS5V+E
IgiANDnjJeO+tvy3ppC+wLf7b8XRyT15PxSFYklbg9jq9XHpMdpdM6uNCHI5
pQjHT+pH0zaxT3NCioDgk35xXARkCTNP5Lkcn1HwzNQD6S6U7nFNCJdsTSEj
6p3PrDF7OkXT2qIG+TS7Jn8KLQ3SiVoAhOrz52BQtrh4iQQPsAQLkFQZek85
ZstCldS76Iinnmf/zQzYE+r2SvnoW/5Q2IZp4RFbspKj1pYSCU0ut5HbII21
5h7Igc5MHeH9N1TgmypUe2sBzwRARIoTPmU4zsme9Vnwwt+phRyYIBYjkySz
UGp9E/zTyPuLwe9xPJhY4FtLGESmA9l0LRJoiTjyjVmYLhCuEln9egi/rW4D
Zv6p5JLtiGDoW+oFb/tUTAhZmGZCbtsPOQbPZyi1Ykx5RvH0dgnGFdH41iXY
dZrmvgmMfW09NYd2OCZALamIp7YimUY4K41LqLbiX3LeV1vgvMJhA+K559kc
17NFJfo1sryPJt6z57hwH2pAMdCkWOS4RxwSx5Awgb0MFy01+EpS4384RCR9
x1mqzAkawrNXTH7RiNuTih3A0220qglnRTi2n+lhY9VKAA+oC8LF/kdnWRSb
zLjGQ4swjEmiLoC3T+LMayk9KuVYJRbGBTTy5AjGbdUBcInvfUDeguLCDGug
P2JsJW2h76ou4qgjRPWbNzCEVLPqQMy1df4eMWrKFDegUsGvDgNA0eVUbAQ7
nrlnwZ1K+SmOOA7wBQXgU8sp9PDt/w/m3Di/FSF0VnZnRqAdo68VkS2mJrEQ
fuDHit5JJWxoANWhxTTpLMf/CHucRfYkVnn3Ken8ptrWmY+0jqFC+chsD4RA
4woXYdqfkxUQJmLPcgoR2P/EZnh6h+eflTCpqpLuUKUVscD8ALpAcek8gxZs
wdI5CN0csJ515p9rvTYER83wf5s9ZKz4v5Ex62j3P3hKEseRX/2Esd2oWBTq
RbATOAmandUcyinILR57yh9e75q/XoYIa9osLfHbJOzyyyVi5XojQyQbL8ev
kAlZrlkNrwmXue6n11C00BLwd47/wXeNQ7NGlYcD1og+Pn/rozXy2DqqzF+v
87uuZilDitPtLmoe41/kSe5K0b8S16pYJfF4f+6T5LWffxazxCHUBB9Xg7mE
jo5d13f5pXnwlUFy/MyXA+O1NABj46fENPNFrKe62cxzHjYz1D6a33pqVfBZ
prsV6TiMzE4Khll3ULBryI+WmasG07bSSi6jO/A/s6FJMw8nHaZFwDDvWMEJ
6EuvZQhaVpuw4oLMnvUw/gjXTE0JW8tA3F1kqXxjcuITEXeOG+plWJzwrfh0
+BvVX/CPLq8g9OUngv3Wco2UU2iyiuV/jqLDRN8empKJfGV7JGSZiYgJ53EC
eeJEFXDcDZKX+KRR+VPuHA9pd1Is691jbt59GGQ+ITpYfG5LgoTEMRwyMtVw
tyjDYBz2kzHuV93dIc3hM6Na46GOMwfarEDnTui+Gpm6MRYmh/DbELX0ZLSu
QzXRMy2MvlIqXCxQSa7yeWYcWkuUSelA+7fv6Mvd26A6ZrypQfdA08nNLxxa
0WwVch8YlteUo4yqPKxxt53plZRZLHKBgHYOPOPvbmDKgPrerYAUiNB7+MlE
G7nAfIOliFgx9RSFFcOszYmx9xYuJuakZ6Vgockwqzgp/+WSEISeG+Dvaxyh
Ai7dwaESSJg9ZHDkPePos0SZJHbNHkuKw3Z31uX+yt5vKTpB9L3583jY/Bh/
13T6+ZD4dceEeQ6Czx8zNyxUaHVLaSHQ5cFFVCgFm6J3hVomx0zNfsAsKBgr
OjDCwKmYXWlfnTtvm+cyjEO18gZkoqTYapO+auc+/HudwW0+QMmvxfG6MGov
OJEzb10cIClPKEsFKJRjwl8s3Vp5R7FDcK7FVNvihFQ6MYX1aPgUdTwl7wf6
SnyxkKUPnbEseukYtkJdqgUYOBKkF2cd69siZ6Bi6sK9G2FKmMBFIxHzhbMK
fR8UhO/3CpRsOT8JXtaFEh9hRihcaTbOZBoHT5PkkXjSj9IqzpXGDPBh6Sld
Yv1qqDoLO9+h89or+udNC9mXNHDsxh+kxLzoy1FLFgwurrth/GMwcuiTO+XF
fJtWNdk/Fm/vlP6/IjBi7HDMR0HaH6nTInEejRc9ejWwF6sa5hd1kbfI5nzP
IfXfh+Qwcl007pBT5oVKpjyK4MvcCB5ahxtkpgcspemvwPLDxms/09rdJx9N
rw9krneVkUEKXbdInOV1Bm5ISHMA6B8kNasbwMR0+OR5PRLCgCNXtt0jfwt+
5y1m9TfsM275az+YZWLDEA8tUBxFkIbWjrgp9l7cjQagGNAr2+Om8DTv/gDG
nLRuufBZL3LeCtpyUMvJZu/HazBZ8+anyKPF6bvR5pJ2oJNjqWJA38987bXQ
uJT/t2p0AzUwUocktQgKuosXDsR2c1a69xpjB52GlMRR1twZA2z/bHwcy9MR
5gd1YKxC/tCDJPENszfrnoOjjIe5acZMzug1Elon1J4KWKYRdcTHpRaNuDKQ
TgS8QiZ6AceeDj5SXct7gYiLAeBg0E8L1wDbHhGDlJwsP+d/1j9eq7hj6utA
C0sUeipgihIHHu8jKz87AcxzsPCQkTBvEYeOSTqH6BqyS2nw+ciVIhybMA28
tz6sIeqw3oH75dI464DqehD5moIoCREBDGmsbyYoc9Cxf3A1Eol6xR4zs8oM
zkOPrJEAF4rwk/KAuLq/odMNPdryGZeZb76B7+ZF54bVbFqH0ETRjhQnUdPj
5hv2qe/wILzwCxB6BZgihk892M09u+Exj0qVD00FHbG9nO0lS8WDfxGg534t
3wXfLv+IaIAjeE5XbNZp9eAUPONI8su91r4f2U/gbRZquHOBjHk2tMYUePsb
in5fuoKGpKEZXMVP0b89lo32vTUrVQ+DeS/MJQNXIdx7IqITfsq+JD7WENnq
Zh2itwbwAGh/XDLzKwMZNnwWFB3j5/8l0Mwr8fJYvbB6ef2j4riEy+HRqmiC
O3cKmC10rJBURXMyyyrKXpkVwg9QhR67Qh0pLnx4bIPpFEAT1BYysmyhIaHh
HBtGs/EmUKAP5i1FvNlZfj3bWprRIJH271vMDBY9YHazpdaXHCSabjGJMaKw
Rlj1Wta3dUp65740M9GDtsGZlCxTbYahO61pYnU7CBKm+3SR4oTY0VBOobJw
nWANG6+rTrFeyQboGQ9gADvyLGt4+L0QqWjO/jTeqe/8o7v4MDAZah+/df1O
N778fFGhHgVqq+iXfcwrY0H18Rz0HyZg/aYAT17MLSwEtozAV11CGqGmDc7Z
1NbQRLmGDiqAomBPoqHqycFhtcUEqXOOJIgnDhtGd9FbFh2O2em9CKt1MBwg
xME40Y8PcbcfDz/STxVWoB24+KwVKGo6DY84vWlAscCifnnQtgV/S8DP8Ipv
YLvGdWm37VwrazUD/Ilc1v9KX9SnPEM5atPIPv471wsAFmkjr/w+Zt+xEhoS
HEoI9lBubMLaB8Fs60m0aQuwUq7USAjpUgQ1nPN4Bb7xY83J8LI9gb+krNcy
hXw7KTwg7kBaHVrcIv4B1O8vxfj8tkUuV8aGEa8G+CM8QnhT25M+/CMlfj+A
3AVA628ZdU70jxGnyYpU/dTZkth5qtjT5XwxMLt0yPFdTKMzx0hKqigwaWNH
br6JrUrK1UfstPru5IPcDqsi/N8MOVKbcDbhO5pshmMu2I3Lj3LbL0Kt4GEk
QYOhkoPtSM7xlkzD2VJEdvf4E5aQDZMQao8cnRSAWuhJQVg7RM2HkrL45y5A
Y2p5V7lebrJaZmfonRqWYidqgR8GT6a7sYA8P5NBFTLwZZKJWo3n3HHTC9ZQ
SP7d9a7qPTKMV3/jLlWCjF8MRg//FM0ot9d9cMaJ6872ofujqAZXl3Yu/Gle
tNsm6KiWEeOmyHYd7WHkwINhViULxHcl6ThKaHijQHzap9R3WLX4g7Ny/fLp
+n5nzQUDKgtjQ6AoqBnU/BZy47KYPi42QCzm23WcomEo4f3iUCyQNQdcKaV/
XCCOQFMFKfTRjKWxhZiMs7DO9SwopzMCxPx0idQ9P4G1Ma1drIagiu9G8PCP
+EJOOf8pLxuQMv3cRheiL9WpwXXKzpeLP0EKz6Rc9PYRDMKeaC5QldvzgYbN
jIKLqeMBvtkh+cAeITbG5g1vXfxUme6pttoNDnrmdlqAj7yholCEV04lwGLe
RZp69LcHsymTs/V9WoOBhba925RUAGU/0t2aRxGi/vn1d1tkQk1LOqimXUp9
Yq7YVCaSPrUBxBqaAf+4DUAJqE1bgUUCRhxYvIlO46YUsY+FVN6nS6s8flpY
efPGcaQUtrldg9n64cJWSvoRO2cCZHqYap3BCUqKMsJCnlgHLDe1ueoaLXW3
gkFNDwEwBhgvGBr8zNjFRejezyFMUGhfl/fbUVuErw/UrhKP66gY5GZlkzD4
bNDpMbk+c/QrBp6XO+g6MXGdkQ3WnaD4qCx3XRHCtMniygJKQxLNHNe1XSY2
kE1Kkqwub9IWRGXHN+b+P32GjfU1b7FMw/L73/6Mq6auCGHz8ZPzWbG1hD+T
y5VB2C7bC8oVZdshNSIFqE25bqDNVfg2ZSbnOcsm9UMbN4Hs76Dz/SirKcUZ
mpFp1LHEtFtCntd9prn4guPf2d+a1AsosWNSlSK/tR+0pU5r0X50PU8RQ93H
DfGdcUp3cKnqh+ocRjpX2906N+/jqU2GBfN32p55laD6kBBdXLDsKDvv3E4a
bHNWtaKEI3hjt9zG0Hl91bvFxb49z06HROwnk1ctxWadgCLVNc7LuiVgiubv
/wMdc7juJZqvNiX2jQIKqJZAACpaWLPsQ8+s1Drb2xRiXWT6a76HZtxfEboP
7c2r+wstDEX82RzjrorPFRz47qctU4PXmlDgBqPfvO/wvrigbsfx6mz+oXNA
jPzzEleGQ7MDLPseurUok7MsKMfWBAaOxwJCNa8+jqmxo5vk5Q27xMzj6UZr
S2MwBeXjgGHhr3CgI8z06iVO4VHE62yyj9Uz9kWAaoaG21e3TiGpDqDbYijd
FO7ubWSu09KDx5SgSQjy7ZO22WGO6yLmcFfWWd6JlodvcIdeqxAomAfmGUnw
gUiSyOohP2Fr2C3iiS+IIAzU8CSU8s90zn7borxn87cLaMygelU/iO6W1qVB
4bTk5v/pcnSgCHFFXAIsiqn2TcCdzJaKEZDnS/Wk69lydTOyt8cysS2JjSse
BVokDY2l0Rx3z42lxtiO5gJmO5eik/kCHhvtakQ09vJbq12QWXXxUEJUB4ST
YnUs5j33ZMv9aFdAkXDFCk4WHOb08couqPQsE/B/ci5ymLeMcf9LPgjaL+1k
1yxB66UsIpiDgrQ6WZhcJIHViJfXKCPqKaBYI5xXdvy3ui0ucy1fu9t59dSU
ErlmSPncxkjxg4sSEf3hH6rhRvlarIrS7yzw/t/bFCfXDZ/HkOC79ln3Mkbx
LG18EVdJ58pK0oGzXuxNAk0Urvj518YLuutZBFvsZRP4588h48OZEsqNfEkG
wbnQ7IcLNyg/sbi0fvBw8SRKeVNTUs476J1TbLyqwhNCqu/fZcAGxQUwD1pX
cyj8VAZqw9Zm0YZJTX72WUaGGK7EFnjunlplDFmeKY0rpn9KJY8R1t9u6kD6
07SAadL6qdqHQxKs9v0zM/rF5ZfvW22FjLLRk3lTE/MdDvCmq0v05IlHA4DH
D23lrs4sQmcQKOPxoo5kkw0cpApsgYgaDaynbh0Qg/LIksOZEAzvRVqVcWwR
HmAno3PdS5NnOpoXTGJbXB1+ue3BXwPCVi4qjykLhGwD8kIl9Jutgi+ExPmF
9wAbBEV0jYWqFVefM5ETc8tOW5cO4JVN+uRn1hHN4yqs6QK4y0sjF0a1/SaM
AGEr16Ct+PTY+JqjofAMWAuFbLHlTEmu81d/YDLOm4sRacp6JlOKlshHRHC6
0T/W9wezV8jZ+TIDQ3WkBeVFiuX4QqAE/WO/uPCf2/JhlGwUG9Wwb7gIMdzi
jx7FowQLwkWmjoB+fU5+Sl+NlnRW8hA8bDxu3CSljmy/ap/aUh4ipdqxEEvC
HOWOQFSf6SzaoGSvysJw3ZBCwtZzKtzID0rbCh0DxJHBlHwbc7aZ6D4+vXq2
uK4A6mOV1tVIpSKUUllAupSd9ihEoD11zXXAkGWB5W9jscBMOb6rBBTWSXA8
tMMptMu06wi13XijMUmh3cpNMLb500ICZ4/Vo0DtmACsYt6O7NXTKgcwKxWQ
zO4uY72r4vqRDB0meuZt1hGzAC/WCQK3QMlNVl2+6t+Fq2Q+W6DjEqMeGHN2
+JPi1ZM+3XHqKXox4jd+cz43NKgzMOls3v4iGie09sUSjhO8yM75n9kImMpm
fC56jjZ7CCKvaE/IZs1efU3KMUsOSTYEk6imPKJELX6yIZfiWRbstZKxwgDV
LzX0126xcW9heqHJCeDni83Yp4YB0fgS8v9nRttJQu9ir5fCo1tDGFelnsMA
CkUfUvovLtcjAzNegpc2jMYqJlp3qUWmomD1Rytf2tecgjhGqcmjKik3lCc8
MOg9liGx7sGETSk9PueMvDdLtoggTvI96Pl5BN1w3Zmn9uCUelNB2fR7Decq
+j7nQAIK0pciTOA4pSgXxQXGRADOPpNw67ZGWKAj+kjsUhqtQYUlXzxQMFRO
ls3V+NODNZLwvzZPpOzze40SW3g4BUHyxq/KHznHv8LnRy3Np2KSbH/5lA4F
fsVD2mOiqKCG9WcngfnNLgQY98DBO3Y3iG9u4+Zq/e6Nbc+bwLykqpbCzQ0e
3+0JU8dfKvhZA+qNctfhNjRko4YbR+tt3QxzxNOLM1ADMTFaN1duHQm3k/xv
2HzLeZqokuqucU5s55P+MnHdnwiD3gShT+BK9nejpS8quBArObL76BlBCP+c
sKrPRjevq0uF2aYrppYIv5u4E/Pdl4EKfUa/vTcQ7u8UF0ULI0E31fytaZsN
loVPFAcLu7WTjgveEeiCRnN3jZ2WmDebU4DQ4vQBiuhCEuK3bFH3xUQE5jzo
eY39cFfI++fAjo3EfpQnWXJUHO8Ibix5LR0pBQI9SwGaIzub7tMFo42H+CR+
0plk/DHbjVcRtdd1HgDBpbSz5aQ/IahKPDe2wYQjuqKTtRs/uzahVLjC+fm7
cLyTaZbHDECZtMNL/g9BKyqqsATpzPjsU8XY5Iyjm96X9HEWKevy0R4g+KMp
AxPbvojTN7wCS/FRllWDgB7UuH9LtUFxQnz4tQzXQpjH6P/ZNDbzkzbF9/gp
o4UwG538WSl0KplEGCKGdpKzt9HR/evBOfs7l6lodoVauAv2080YxSbrk0u9
Xnz+TUY2Sduv9gISJiVZdQ78NU8WetF3mkPfdpnmQCEfkJAFz8hVx9RhOW4I
DZZ14R7Gcm0Ev1swpiRW7qBCoYtPApRkzX9g8v2mo8nh0xJ7NQO2H2oYIvDs
MH8cYVbCgKmFukcEkvXFnOOn/2r9qBpq87ug/4uls5zb/zSNYW5RficSQZgC
1aTXmRihz5/XFnewFob3p66UPtxGzeeYh5liszn6ChCRQ23yQraLFFqDrQG7
xTjldbE+pfl4LfLpStrof5Zz/uFYv5gPQhQZ4+gLkPYziDL5NDlPwl8aAhjX
4BX+t8xNgWWcntYxYbV3ZkIHhj1Re78tVDn7fgszLwqWN+FYwQdoujlx2SxH
ViizAGFlWtZ/tNTf+4ByUTXkTu+OoIVvEez9rMRrz9XFYWtx1Ho1pcUnq/nt
T7OW3UJnAUQNBMpM/eUwapaZb7lq0dmrtweUAcrbmLWHEr609y70Nbzx9aXG
VFjtdIgbQLfXJa+3xPXoN2D0LiLvpH8piXeN5iB1L34Kxgn/HWYaRn2Yd6th
vfDYDZd5PQ+2VsJVtuhNJL2kJmgNy2/75VP/5bACIsNqoOgAArizuApMEor6
GO9QgoZGHvO73kZvR9vM71q8uGIbgFilL0FWFlaDP4N+gxhrt57NJ64C5DjP
PJIuiqRt88/9LW9PpP+5/t+pfEEyBdn5m8SMnWQbhdI3dTCFKhHzIFS4K4Nd
6DDNjiu2Ix3QyKcyfo2QC3t/snxgKB8S2hMEheqLOHTwtbnudjN6x3rAic8i
ilgg1v7ZzMnxvH3yDpdsQ4W4XF2QmY9VLwoAbkUO3EPvD1Su4b1FY2rvjPy8
i6pxMb4OvZRUNlNtUBorksxVS3UYzPo6wDRCJO4QO838TcPm05EIOdyZe+oZ
jjguy7Z3kFTnc8W/e2lz8jhmrhXm8IopgE7NRgTv7fX5gC5jffYrLqM3gtNp
yeZ0QgPbryVw3nIhLwjMziSKfDrETvr3KTzd+d+ZJxx3QFbzEDgQGOHdkzYV
8rxwzZ60ji+yShFWWUQl/eM70rQ1ztWoxMweSEdPJtdRRjWoBVMA2yJc9776
s0rdv2+BbogzRwnPYj1600b6noawRnNDXTge09QgcQA9FqAaY/V6gC6twveq
aAp2hF8hR1INXf8hLqwop+Hn7PsQXUWluojMHILnOzoBBB0gYcsintQ1upaP
7MBRMp7ifiKdOLlL86VKsy7QpDIPwOs8xGYS1unJyIekxtITGNwxfcW45xI2
8cKWLkm5efu5k/MjT3fFFBCbx59qtPScvXd5Y1hIsKlXPPts/a7uVnibpgri
a+ECVy/Sxg5/LjL/4hIN1Ha9WziTvSeG4WqPexiI/iFNScpe8nFEqxeiAkKi
qT0KRSph02HANKfh2ofxspUeEb3iAMd0zZ21nqDm8wsBp36vR89Wm6IVhY/f
OHUVR1n5bS7CuIe4QRyD9DaOSeeKDLjsNSiG05+ug/noRDZnFsuSbuyRzBoL
8s/e+OMjp22vAjAfLUNsyO6xp2ctpudjuysmsrGuh9Sxec5v3joaCSwha1eE
lVHwlib2F4KE1xZGo3EZ1cVJknfUWh/M+l5BFAR1dgsBbhtvllU//V66vtH2
fDvDAudKD6NrNPiwFGiyiuxbT3iVjIdUVQii9Tau/O+GeZYUINohqjGNQksj
i3pWZJoXlqzqESXfJEz9JdJqakm+t10eVoWpaKcRUPtsS/zeWkLxHnrJ+5VS
G3irqjecufgQyW4G2MLTmn2T588Wb0Mu5t1vh+J6Dtk0gIYKWyGu5Bfh7lsJ
QgH1QmEtwG4Kx5YPR4lFMQq8q00HO1nJP3576kVASGBPqHFJvrJ6jmwb882M
Sy+O7WC0Hg/cMDyIs5+iMVfXZx2dDEZuvnXIPUXtzj2afJLhkURSKBkHb999
ut5OEAwhABOGSw2poZxAwLuXtAoZXyfu5d/I0ilbol76FVBpYX1EIiC5bFQy
uxQEotG0boEcmBh4g56gPSSKA/QGhJP95P0XDFUiHFcFFpiWqnpWmZuQvIyJ
VvqzoJBM3MIc/TjGNjE4A2Xi01j9YAPxvFD8PA4JRqJ28GIiQcNPRjzf/5Jj
VCyGBYepnESXqoA/tWRhctHqgUfulgSjYPFxurCnurCSRhNZSFpoXlcUFo86
CBUDHHJfbeXzyG5x+LVPA7p3WXj0hqCjpTR7fysMBw7SAVd3FV+Wf50fVOaB
pEFrruf79ZVuejXqpzZRO3pWyYggJLutF/uI36SI0wc1CMYs1qcpX4bSJzO2
puB/6TYUmZitZpNWXDTqaV2YeTTq2fTOz+DnpE2BdezXWYLeQ+3W/N5OfO+l
2uD9+DSmVTKwx+B7RAGzB6/ZsvmS1jpH04SzOdNslEt5SP2+jeueBMqN07wy
N3FWrKDaPy9CY/tgvaNyLtDFne6e5UtsrkQkoAro1nd5ACTB3rcY7sYTGzaS
2W+2z/pOpOVaxpSUqPkIgC24hBTE0jGkNwY5TAnIV4NjJJgGQwf3vtKRkkzG
QLxcQsgmkK0rJpdNxWG9Wt3CV3ahKCB0ZAdx4SzTRN8Jr90aZTxXRaBqKEgO
I/b/+mGEySuatsdSqm25lz3S6YKHltV2wMKvvUQv9rsStr/JbBLPOobN9O0h
FzBm4CD8VVt3aPMFdeonUxnWuPbH8zX5HbESG8xW6CYL5x9Z9akIRnLLBPmm
aEz2Ak1rvFrBy/8nWJz6o8BQyzMq9omdUyS0jOZNZIhfyorMIa1Lacwp/qDZ
0dc3nGorueHQJ6AVFRFLeGahQoQ1yeQbpW0ddcP433Vil34ohWX9n873Rz6C
PBbAsKg5cMoTX/jo5Or5Yd/I+KmbMNaOXpwaDXgCFjRhPc/HWlknF6Mtcxnp
WIL4ZkcYsETD5imqXQjiThTqrpsXyzI7IvSE6VF4yJJNTjIiEs6j7aZhnYoU
DabExxs7uit85/owCqAvBqvvtlIvnh06vrGMienhERPonU3JQ96Zo0IaVhDt
76mYlhLOlM+J914FfDPi3rStWVCtTTJZTc17gf4K920cyYhLvGcOnSKOPIJh
voU7nqvummMB94WuYlo0Ho1jGr6G8XXt8wMKF+tsPvOkqoI0O2gQnKovNzvq
msANmUt0GlYfTRjdb7rvk7+RoPq+knqpmscmMYsy1BkT+UR9KyOD5gEbeb55
7OTcR1d7FXdSU6OP8z4q2Xq+5XuEJ45tTP8ATBtwDrhES4o+LflWmWP6noEp
M3umqZXE3OW1x2AVb8xnty10x0f0z0sX3s7LO+sp6E8WS/+jdzgol1ldACf7
FMCMIpDautjCZywHFLGE7zlSCFNwAKSte67XcxGZPxU5uSpmVZxYvYocaW3w
YPMMIPb3ZyGH4rORtrLrrdiU/jszzLSB5eLXBT26AtyOxYLUrvhKAVFa0e0b
ueAofNPW/fk54ugwjq3dNeTLrnV/NwIpXUISfSuNikbraFbGcVr6gMhz0T4p
wiQGJP2ahm1uI5XYXHHobkwn5xTjGnNxfDL1XGuTWlXm7am5XtLVuDlBjAmy
dvyyTnEkV3QNEe4geG9SXjnuH13S71+o/RtZ43eModN10Tfpi8RMJkGWdoLt
5kOE5bfK99Ael0gv+qN9thgroGEMvM+IpUZjqzDHNU4mgiMdq+C2rabGFalF
aWlFWo5nVpwITkHIhDIdT797Fgje0KILCew/Rn0TjQZXyV6YJDJywV7lgswz
IUvzz2h3D+GUyZpJeweirJyMqI5Aq4oxAA9WotCV4kXlarUaoWqLCYeuqvHe
2jGc4LFVmOVXyHA5vwtd4VmgrWDu7SR/7N8vR7Bg6UKiZHuI+h2dDQMVzx0A
qOkti/UVD1p7hXraO9DmZ/pvxRZSX/7dy0EBPgoLIQYG9U2bqRe1cHg7iqBx
bWfjgALDSPSf473M5oiA5lJ3yBquFEXAskbXZ9M672xoxJwjMSBeJ51MYbnv
M8yDpxwmnLP6VcXtSyNVOGbRR4E7PG24k2Si5Cy+x71xbsWhi2WKqv9yQBm4
htBOZGz1yZerw83nuNqkAymhSfAJrzR0dgzJ26UBUokzjciqq19wBBfE8Zew
uCwnqtFcmE3TTy0JmocmI+K65ROWcwS+K9PhcbtXP+ZNFMs4KOneJTjHNmJv
bJ6juSfx52CqbrDKXdZCwT77O/pzOAcyC/Xsw/10nVN/KWgCq2VTYTRaWeCM
XFkGx0CfuZSN7cneJLtcg00pMcB0CYNqV+Gs3+n5plgNcBKEQPVBhSHPLniQ
bGBnO8059CiLpjToIn5set3quOQ4ouXpqM9v1/lDUJQhb620IUu69oMWJDEe
hbooRGqEnwiZDvPJbHk1IiDKSKSGJ1QS7FhsA2uMid5IZougcgn7PK6+QHBF
U2GBAZlsowTjjjBwjuQl9/ziDZCzxichJt5Vzi8XGQ2+V1SyIzXOQBbWE8Nw
93Y1KcT5D8TbVTO6WjCmsP+46EiprDv+UHq+q+abC+M0EEfT6YKbp4mxPI72
KPH/JHXI/JOG3KsCeeoc67t28GgYPqJo05N8IINbfunmZiNkg9oJI0kYaUE9
+gt7ZF40mEzO2+DlgTLt6wpFHpqkI9qSHLbAMMGalbPIAC+Li5ZQ02c5u2ZV
cEFNDn+3aecRUriDXtfpMpzZ9s55AqAKo8uaamltVW4VmwT629kuby8DgoQj
M5erNzhD0nt7v1NBsyRZrkjIZ9JHgE5xx4dtofT+mWcvgiFGTHO7HHO+5olt
DnODfRfP+pDYZu5yl9qsO0W7yGukiL+4eYGeTsEIm3kvBQwgTqsEWCSocO0H
TpsogZM1tqKpiad6BHqhk0r8owwMSN57zVn1eSfpMj3BMEv1vpfPQXqgP1hh
6v37pKXwJSsu4LJYcC98Y1EIuAIA6EuBmAzbS9wGqPmHurMbyRuRqbZtlVat
Erc1rq5klv9GbayoUKYvvrsl0Ec2o57HXBA3+IYbFzfhrOGoSd6vwQTHvx7o
QBLiG81MwQatObc5IisBX/+k21DdjGLhAxmHZ/BWQiuPpYYFN2dmm01/uyCg
wx0EOKPvEQUVhXA6p7b9R5pMCNXNn4tLAP6chAbwx0dIYeNHn/NFYXkLwvjl
oYpQ8KvAT0Ja5u6RnHKdwgRm8GmzrMO6pXBGRLImchVJcALFqUvhP4NcLaKm
6Utf7JheYnb6vbdxeY2zKRKgwESeZAlSUzzscjOR0YuSNNZ38ZpE8gvVvc4h
Ir6luG83qmS9LbY8eM2mkJeLjra/AyUlNcIQposOQwJuUHfFlpbfGKNLTmAf
w6jpL4fxoZ0ySvaqy6HvvvMYzellKavGnCDnXwwM+dyEg+EqiEh1vSsPXaoK
pOMwA9DMoBk+dM/htocZBLB4oWeRMWiDd8uMGrc0laaH89V90GIkuBMlAAEl
ojKs2r4QnQF5K7IKGWDM4IE4Fu33Wb8Xtg+6zdNZ1U7dyM8NGRDysIGqz/IY
njkteTRmOd880lgnsN6yeeI4CmQMn7mN7aqHUp0P1abBkoxSTLaHCU5XMAHz
fJMFa77nAJgnhIQd4DrklwWW4MQki3zsnxlCNwWn0bWDbYoFdLC/rfYN0da9
qBzQASPkWNywpLfqhZBA+8f9MuLFtqKA1u271sQA/Efb3kdLIzebU2UUSAy/
nycaJZ18qPnZRxmz3Q9lJj5XWegpJ1zIyEFs1T7aShgkTUI2ggnPmpzLwAl6
n+eZObBdwgP6oUxVKgMOcX4UuzWf5Qe7sI5utop+M6KvTH7eu65QjZ2iZXqf
F00OURpyxPGR1Er15CjuGot6v6rmDZOqTumsissu80Z60oiu0SUuLG63VhAK
t/zFo1GOmvrj+AhXsEVTm1J9uEHBoYbvxtvngQil4SX2LHeoI4EZl2lk4pXi
HUMjrhhjOTZadipy8KVRSXSZIUT1MCLANxjG79xcklsbefjnqqi60rXjgmsZ
1BXB0oK2/lj+stpobSH07JtE+UYiYn1ck4PqX189/ZwcfUsVk7E3LSWQhWRg
rBNjqtCAwqwoiH4OX8IUv93bIImK9vd51xUNLajMPOL8bU0r4sIKLSKjNH/H
CsxN2KDax09Wsn/r+2SQeHaK6iCBqqFoYEdYeTG+M68kbckTGUwbI46sTqZM
czLiK4wSOurlXYZve8YMlyRpVTeklq2eH21iy5v705Z7TSuQM8QvvPlemnak
I+7VU+6EVn2g1XS4s9gJeVZa2vDq/Us1nCmLAq/MJBpiNMk64mclY/R5GayH
tMklsIRWRCI+f9CKP5Mi5097hwTREurUVW214wp4GqLfVw4YEDd2+0viZ91I
/mlUW5d3Ef9X4qloMyH/KVwMX49IaGfDionjkO8v8cyQ+HAWxLV1EDv6tMrk
KhABQ+tnOYC0qqNRPKAXFAIN9aR7RHUgIVmUSoKfTGGmNSra+cETwrcSqJup
8M6nj8lpkDELTuBA2wrvUGXCo8C0xC6GQnezWqfKkIvGjwqjzOGQmjDfTpkS
A9Yh1gzmmYTLmHQmvstJ0H/hClOoYDweq4i/hmtCBE9XwX2GdOo2F7Y5RgUW
OLOSc6Qhgy2XwoDgAbUaBWmBJVx6naaIf8TEs6n3JDMvcZmycciYRkx3bRML
CGMu1mN4+/zI93AFgPN8GOkKAEKESvUsqrRcUnVNWMS1REvAMQmePIix41gu
FXBGFJ3Ak0psa/ny/gCplicupQ3N287q+OOmEG/S7lCJLxidii45cmqqBlQ1
kfw3nnfKdSTtKyIUTcJO/8jZPg1BUYTEwGdFVzwRIgmseapEcNwOLOHPaLVr
ebVN85YVbo5PVi0nKgX4UuqgOarJRYnrCkMiINSJ2kD9xtoyRKS0JbJ2yW46
lH3DNYxKkJxgZsiimWMp2UKtvyl8I4mFmpgLiYZVkuCWF/+1l/dw0Sge+8Ua
Sv4DFC+sHaUYhUVsUDPdjq1f5BdHMby/p+m1z3wP51Uj1X2gPGUSw/toQRov
dPFHG0YiwHLlRqecAoEDa+iz5s2yEwf/QF6M/J34ETSP4xLIgjGv5sY+elwQ
n9fx3AljxaeR4/MEeIXBHrSO9uzhaEUyQq2N+m4KFaA9zrb/QNfZ/c/Y0EIP
Z2lKcrB5C+SRWEk9nmD93lVhE+32xkE587iZm66tBVBKnAdYbj0xJ+QEONQ+
kib7w2lU3H1Nbk+YezL2kb7wl7IAHSbWv9ATRu1nkc7G/x7svMs0yjq1KnDo
WUxnWIG2uny5y81V6+jeFQbOHnBmES8XRYYiRRdCnCTzWdI0+0HkBWUnH9K3
FekYC2HCxsrZpsbKgZLegBZ7zSS0qmaU0nd2gJbPq94DewdqPaqG4V5lexu4
4uALg0yarlnhzRhpJpczIJ7J/SvbBbOjrOPbpVFjU2u+2Zu/BWDMGeNes2A/
wlLpJSytFQ079tJY2qHVRqnceqhwlw7fegQVxe2ajeeowo6XB2jtyCkghwTf
jwjDA4VgHV+flKU6Tlov6eSAbnJC5H+Zb68CncA6XXslkQXdELa2qGQb+MTf
2WaFzg9A1v72rFdT60CvOrPdgC1JOVJBxMMA8Dpg/fptnGdaORGseF5Ff4h3
ElQoumVFUE4i89Lzr8LrBR9ju/Q0ozrdh9xGOkLLXt5uOiDxNHlSAuqPcQuS
ONISsGwAsuEKPtGTbm6WgYyvN4H4msPdKAzPr2U16TfNTkIGIVOgr+/tZIai
YSHd03vJ+UzbZxYpst++FD6N9H3wQWdu4fQ/m8ncWOA6qG7koL6CH+GFqKvQ
Wj9pDEfmScjsO75X2qm6onXvceoFCcOdqtYXi8KUdxlj0mKPi6LLiCQYYzEu
ACVBijWkSkf4kj1XvfWc6HUl+XFz4L2CU+k5Rhv1L54vTlTpUMnVbaUdF+Gv
OUVxqtwpXFYjB66hUkr2/mWvHkCblQk4avGHVV5QUZ3LGW633sGypYzD1D8X
Oj9ZWl2ETYYwkGs0FS0fHzLemXrcPRFDu+0DoQ+vwOEKNoHBr0LVMx2I8j7u
Ni5gDSTZU/9qihhhz+mVFdJJaKFawKr/7Cq65RAjqQbOv9fMJB/eNcWh8JnI
+jJrzgWmCTTE2juNJXjAMC/GqsNaPBgcjScRNbyVcpDAcd5FmxfvlZgOrqRq
2OijyCN5F3HJdScGiDvaMSFmNnE2I8+faNSvmSTfM6xJxy5rVVwD2RuszTyN
T31kyRnaqXC7szV60z0ZyUV5gs6gm/8fmIk4+QtZPlQhDPc0sz2WnaUq8g8w
X2W+G7dS/e07uog3oFSNTfY9DvGFe0qv+AHdoJCSsyTKY2vzh+/YKU64Ll5W
fLlrEpM7YFnA+9Ql7QRT3LrYtpRYWPkTUg6d8JbE4BWQFnfV4o5B39ta9Kd+
jdLHUwsX153/MTliciybI9glg0RCMqozJTn1w+8ob5cr4nf6CnLObeQvFs7u
d9GLCw4J2OVX+h1WMIlIxgVafOCN4VccMjzRZ5QahvUHRumsoVYVjCsiDcMu
69BiTYij4h8+NuXnK6XlllafId1k6l8TUnVwySk3JsMb9EUqFuWLsXCDVNyH
eiujrCNwzHGL9l8BGx8sjlkj4y30qFEKVEOM5xBgFsRgnQwan6qiacvbEQiz
wSjwuqsf/QWnS7XhA3x3FKsCCtZVpyjMG4ohS/TX22Iqv3L2c7F812ip37Qe
msy6dzxRfohmtH2gKYX9RPFKgZ6tHQpY64AR+/jZ8sq80oxe7VfBRX4au7KM
jPUFFnMqw1CKLV4AWRAUjskxyxs3cP8keMCnGqWG7marZqiVRyG/pJXh3uui
vsw5cqz5xwWP19k8idNv9NNoqhEcfLBywdOU8xh/wTyTK004VCVObIbeASCT
1W7PD7B9xRpV04/zN+mTpogTCYwI4kulWzjCsCvNrgasb1G02jzf3zQxxmZD
6XN6v6OYLtr4WsUEXC0+H1bhXHfoAQA5Hqtyw6JVgc8xwyVhiDsqoQMATfE3
1slvFnJNlXD3fc/k1ZVqYWoOsnid3vAFDXu1dYhqE7WDJfE0t9hdtpAlKtGB
bpzLy4lPsjugnUkYWtB8JOi1n61UmZGc7wcr7fZxlvWoQIQP/w9YyHwAZNp0
+e7Ic1MLBBu15r5tWxFtCDl+4at2fhbVwID/a+Grk9VhKJveOLM/bR8epDK8
krdKP5ERbyvd4efLwTSkkewK32qkOgJIPitKsvBixEF3wKQcVRCtc2CUd9EW
2EZRSt73ATQ4N/ZOJPU/LTP+SQe7ouwQHrkmZ7KbwqgiJGSmS9dwjrHYY2lu
OswvvolVFbBMfLlItpaFsT+pqDUT6uGdeTn4tR/j+TS5jERy1wYkyEaubucl
QLp/WVpsQ6ql8lWcWONUOpVuLGT793pwNa5rvfGRGR5/NTWrJSO/s9vGQ4W1
XvYi9cFRPoV1Jy9ELuBSyFU5f5R1il1/te7ZkEU1yutrwiCkiLphh2iBe0Wr
N8HqONGBJCD0Krnuj4Howm+LZ0MT803uyd5x8kyxYXxdWtg2RDd6OWouI+VS
7nkZZf5VLTX2aDrU0bMagRe6bgevMnPsmgIZHBqzQoR/sTKREsR+FgkWCpJm
t8xCmyqO4+6WTa4qR2G7YuQDkHcSRD65AnowpT0X8kwMCtmTAYO4HEOAMiFq
mJiwkaVIYt0iwF5ElQVW5vCIfIuoLfPcFjJSV7Q12cLpR1E+vNOTQzUyQo3c
Gf5wE1Y/Zt6vjhLVpsX5x9UjNXYz9oflGkzecPzhI0+p1SwIgOSg8VK28I7Q
qHNgS/6dEI3KVG3KtF7N5SzG/Bm8VCHiw1OlW+Xmnz6Ahf1eObOiECSHKoGE
4DV0XyqHMopcvgRhrRc/V4cTfuF2je6AFc8QH3WImt+EzkCDq3kKNk9BSbDn
5A/BwhXcpU8m5LJtwi1hSGAIaxxLQdE74m5f8h/UnbnPlA++ktFGVpAMtvfn
CU7UUq0Ttq+CJu+nVlOCHuTP5MwvGobqrmRy27ei9DGe1M1YhEmmISB0unjA
qdD5+0upAMRKmszv0jGAuPx7ebhrjDBNE/+DAEX8yOswBpNZJAvzarKtfnqP
Bls7BLhf0hHfv3Xnhg4TbwI5iYMw1Pn7JItmPgi/CnISU8KRtKP4hrL4NZMs
IMfnKy9RGhIioFwbHiNY2zUUVPEkcPlhttJ2EPTEYBQaJEwQu72MUXfBD5th
5FPCWbbfZ8wwoP6c5HEU8mWcZKW74WAwUsTBsglDpa5SEkkYcyrTXvQoc3Gw
UkyzM2KSw6SPT8Z4PGnhIMQT6L+gkZCN41pxAznyK0j0yKSfuXElUKuSXg9S
FMjGPm3XIyqRZpVdT6vHpdiEgojPe6UQ77mYgrLsLabmIAIyivaBGqydKtZl
rHODtrTLMCVBBp6ypRLY0E887XagR+c/TW9R57lTHoPihG9dlh88EC8U8b8e
yq//7pe+Ma94dr9PyoOpm400FHTtBFO211kCpgrCrGH+VVgAALrAQ9dKkiRn
L/52vC959/Qelpa2pSkxdsz0HjivVvEY6T0O0hmFAcuPoO2/CkrjMAz8dRF9
kNvb6bnfATTqSpNewa725NCUP+8CMFcHMcG7dSxOLOWKob4gqouNaZ0RgUJH
UHCRI56N2uThRfny0mCdgHll7Lrk2uuZXnsnQ8oedF4PfWlCYjUSrmSn/ve0
mHwlOusKbON8Q7s6cobiLjKxx96ll66XPQyQLOhFjvNEfDw3NjL1tXtFhHxr
vuoNSaU9VJEqg3ll9Npl+thllwSTDadp03d5lWyTyxIt/eNeiMCu6dwi2NcH
c8u0WMeuzzEMP+cU8scFYd6gbOM3xfU4r+ggizcrO8NsKoxem0Ze2NNOqeWR
hRCbQ+Tcmbt9d/Z8Q9weumb3y1nG5YDPGXmc7g65hS5l/H+fXf7knVS1+9TV
hQQL7WEYwjMdTTzGUobN2Wfa2aQNqjR/igI1Id4ckWxEnw88+PzCLU3l+gJe
oDeVthrnjssvTDlphOHn3GcGurlERT2f2kuSZH3JkfTTOk9oK9m0gW/AbhqP
U9/YQPlh9HEb9gCDhSsmLMm1N5b8sWpTz8zH+osJczjuoxbxY5LZYrVjQS1C
aSj41XtCfZOg8oPf8WZE5e/PiiWT8p9gc0JIQnUjXFH3K9F3t8o8/JUZPvFK
nCSXcjA/6tyQ3YjgWAhTUrkconXljxXfjLnb5Jkg3JQtAkj01AeBmK9VkCg0
VlJ3uqd2xihZ8OIi7XkaKpirpg/gluXtW2l1B3OdPxUnP6AyvR7r4BukliXm
S7rpyJbw+Xu3ILjUQieHknjER2+FBd6BT3qsgh0Ntq+3qOEECQzqNxNNFCRZ
oS3MEP2GzV79tkUyitC9hzOKvoHdpE4Z9kZTNPbdx4rB0+QYe/eyCTVKoHQW
/hzdf0pi8q0HR2RALAw54izz1NP4XEfrT3tGLdEHYLpnqB1+aUI9gNiMgbRU
GMvEAyZXhfi/tOcw3TlhDxnduHb61Db8tkZhnGgMaNWCd4MvsPTAKVWUYliZ
a+EyQ3ekjorCNRrI5eEE1rs+O8S8EgNthMObAiRz9YzqaSEAdh1bzlS/YCGh
RtZZExQrwg7hzKXEsMOJKFyCWIuMzjLA19Lj2jnA1cwScdKsnyUh03/cXkKI
v22vewelv5r/carxPzNhptX0J2mMQCCNLnWmG7Ko3f0XyYqH8XFahmBxr7zu
86cin6xCTW/XVWLKCF2IAzd0PNKorRwcpHGQ8EA75Wg2R9Cjr2wRqAQNZr+Z
XvDpv7hjvnut8vNKgxAzxG/dnjix9QpKdJgLqm6GTLsRX7i6MYEPGgLWFiZC
TOApYTynLTjOzGfAEs6Di5Qp2+RbRe3HP+R85M1XA/kB44jxkKf6+zb8ztnm
GnxZdC2lcNTgK4FlRPI6ug74Uagxp9dupAZ4GljS1KgdSsLu+JUWf7Xxj6vh
NTi/HyB3jHxnmYUmKU4lI+8p7wLij5by05wpM/GrLE3nZ+/4tgfMQAtst9En
L9PEN2GlEBfgEc6mUpVv/6ZoeBsgA6ieCff656fV0fDf0lrL5pJ0pELl8drx
YMunqVMAYTKuoNtdE2qG3PWU6r7jqikN+BImgbYftXV1tAG3G4/eUCbV83mB
KT95E3B1JPJmWG26+amcMIdv+MtDGqmOu6gZgiaboq1GKmzUTzE9jMXZW8/m
mxIDrZ8Cro0MT0Tv62TqAxpd5FPcX3+WrzoXFZ3KVLW0ulsMQWIcvSmfWHng
koDC+IcN8haFPkYBwOqeoQxs4OmhQaJ8XFKT/1/vmWyhQfZv3EHyEoWNibF6
951xqgUtgbpW1FDy4c9UOcphVeDXFHgsWNdzUlFDhH7+bKG1It5Ro+PVT3u6
UkgVe5AYZ6vl30lS/9HiTN6qXGAquYYkqHoTFtCkPFYFS6N73Fe6dGksvhR1
G8VNjpWbhrDvWPXbUjwJr1cPfPzfUdL0CU0BQqDyXOX3NEzjcCxXj1IaJrTj
cYT9ccCEn5UeGkLl+7H4wLMdtzz8bpL26bzzYHfhVWOTkQgnb+NYJ+hoTGFV
+k0F+rz5sOQCu1mkPiu8noxgO20XSfyVGv+4oyI+mlh8VuSbhc9+PD+NOjiH
wv8l8UD5owPzh/AJ1tNLAMoluch5RMGEOTg2gBGSP3e7qvcJI+JAN0dfGUho
hdUGPaKOJzrY+02J1iA0WuB4y8SzA0atCg5kwS3hmg090+pEGwY4tNk63sfB
C6MhPsMsPK8u/4edW9nDKT8tUTP3hjV6rRekfyjZOtknWw+o2XwGt1ICLEK/
u+oA5FfNEidpelJM8A9CuuIOTgKN0vWCaDqkRziEcUjdPLXy6oTewLxJhEbt
a9XSPfCL484yH0bBgci8rebLz9cFM5msPwJy6JQy9KV35lBqKP6lWQB+ruTI
wfzQzvXmu5rQd/o9OCNsBjrF3rMwrwx+1vrhB1c+PLecy3LNkOz8j7gktMEh
+Lto4BYU1V1yuvsS2VRV2UYYhM//2JNNSmVK5msagV6RLmi/61GsCEYgWTCr
DjShuu+ZrXR6T+D6Wgq0qa7/yyUFtUbTEOePYNIwTD80uuQJxsIkZ5hCHAxL
+M9TBAx30PyyYIgKdnqatIXokUVv91HOZRBl2C/YZ2J+E+kgV8weovdeauXj
FAcyadp0r4ZL75e3tTntJvUWKmWDdG3+PuqFOse+EZzVdlw6VW1qICBcovHn
yOc2+ncEC+NXSSLvGKtXYdVX/zbLXaqaJ/9l6o6Osnh7aLAVWzAezK5YAsfW
3DDyvCOe9bOyqOzlWyDpgzRBT7UNdFlQhbwOtDLOV/wssJdwteH4xAIFiX0L
HakmGjRhtT6j3Qs+vKJHLoe3dyGqkx36vqJ85S2Is8OW8hclG+JQZGYKAhhe
l1rrLhgpaoWxlt/zPFvIE4N4odwopdcdAFZ2oWIQVkChUKD9sSEe+XuO2wgk
3Xh5ynxh7iveaYfr2MEcmhv3UhpIRRHh8AvQLTnTs1BdYWkNBGAD4HVOb1ON
Ba6VpZG0xFJ13BmVBfrKYEOsZPLqpem7bS5unLBPMsna00S2S8d+DlCKPpMR
nMR5ZCuvHy5VzeALXIdilCRgSO8il2PY0boI0sNS/hnmrChYaCdEHGIh4Bai
y8LPkaE7ZRDJolM14PVi8ZkbHxNOEzl75wQBRDa8x28WKVX8Mr1dJPv4oyWR
5ftqCoHfIY4hKN8F6AWiXxeUcyQaLNm2D0m2UwTXz1jKeISKkOeDh3U2+cS8
FRJ/HJz0lF2xGJ0ROq1InjFkonQojX9QUzSDOA661CwCY2zEinDVOGpjMGdQ
zWlyFcIi4YS61cLp7veOyqn3Lmj7x5gOnxLO1tG18qo2s6eHht2ykUXjBlP+
9AH5o7P4PTERb4z1pr++2eTouihth+AVs+duSWvqLftoA1q2Jv2gENB032js
yIgQef5oE4DQnbESX0/G2sOGtArMbFvJjBVV+23zgtsiqhg2u70DswkAdIWy
YffOE4W4AKS2n28MWD2pUw6dL+qJmJ74d32ygJUMtLSkNT4cwUTI831nBeHD
AW4dEEbFRKHSYYuC/fd5rNqoDLxfxEPeTPhc4+US/nfSRb0c60kNr8TEL10Z
XhqU6r+gagovCwJWSCcByKLO4ZJz04quXO+KySJRShuqjrGZ+/JF2Gk0Hq9E
jXKFT3oia+dcMlN2QEelTOncUffHw1XJQbI4bidRnMwlZj9Em56Ed4ALfHWp
aXQjXR9JyxuNjTWphkEZLQRYKTr+XwVnsQ1OFLo0gvQQ/d7GI5vV/fIdtfzc
0jL5EJ+0WUkM+COB6AiZGo4ksJ0O31RXMnIl/zLlMsh+VF5b5rwPYSilRvUJ
nJO5EO5lkiTWYqmgUSiUEmXPyjjiDJfQubsdVLooaLiq51c0NRFZp9gztEvC
WwDsGbDFE1g0ywSD6ArL7pq2O/qKrX/PGXVMv+W7GkGxtbN1clAs5sHJ8bcq
vyodU5KEif7AbA0ibsXbX37baNTownGTfd2lYygbfzmP2HzYs8yG4ojAWhcg
mJ87Pq3apivYfTBLJ6EZj2op2V0C2ldLFRYZBrd84fEAP0pn64f89w2SqR2b
BmzlkH2EBQjrqTzmzTVo8z4PkQ23VQTq6qnclNt9hqZOWEKFIuMxktALnfLH
ebI//ttoZ03LJw7MENI63/gOWlG/JRHt5QkMqiF/HLS0gFO1opuKaVrNhmtt
cssGvnblozCRVmHiMA+BWIM1er2Og3y4hDzqD7rxDjwUhmLM5/ELb06AI0gy
NWuOv/24FLaWOGWQe+8SOqy3OlWw4JzowJWwu3zFuJChOC6qqAdVK1qtEEyI
yAqD/0hubRkR9eNFK8lBD8oRV7bJsqznzu28YYCGQYmTZ/pkajl71GkXWYtC
5P6MYWNmH1PBRSrM4oh2qoltF/8XEZbQtfaPcVwnxu4AETt5Mw484ccPDM9g
iuCYZYxOeCj2BFMFV6ApjlGGv5VcKp2Mmc+Gx0/Z9LH5P1QChvyB0mhz58RE
hH9yIzyjifONGJDN+o8pI29BlVCuO1RzD8FWWUhyYUN8ornOpQEs1ihKpHGd
R8j/9QmAQRjEAobKpknGYftx7pL+07QqvyB7LNDyDMzwATRCqcHRhZJYbyCE
tJkGY5w9qMmWPq+MSPqXLKb3INswk1XXjfRDe0bSzyGX1TguRJT6a1kfj+mH
8FvWCkELC1DKbnhGePqJ0ThHdJFRdwRwCOt+3KtA+9sdCyCx09IKhxFikCNX
I6eB/2oh0sri07NP0PWKKftOhq9rEZv3EvRdyjugVNEbOJA+HYwnJJujR3Xx
+SIgjaJs+NZOcCLOcJhgjsQP/qOvLHr4Iq/Wsqy13VO2HSeCwJ+K7TI8lYCr
iwwvHVkECkEGU1EN1lWjmiCT2LW0nD47h9p+q53rl76ryX944DakHDZAm3hF
tJluZvgzAq7S2dsLErDJxdTpih0mR+NLBWzH8n5/9GTlywOkfHfYnFuG1PXm
zhB2fWZF3c8xQMd6v5bQxUaDpcl32FddjuTjCJFcVdjS25gn/IzM0Qyh+AHm
sNSIGshrx1UkR4kK1ggaQLt1sWgkY6hfcRYBWx9U0wS162rrlEb6SA1pD1Rr
6q62GAWmxkEtykm05TbEDdARx3WTVtuiyRHeCCZB4a/8U749Sqp6LtyUIion
v72p4SXh0jGAY0xFsLaYqxr6zy/mgWawtkSCE7eX1o2KmadzNdw8gmEj8r59
1IPjq85K5SeDsnRkwd8n9bt6EAv/cWDHmSdwsAjOEGcGKfciAYTFAkRJGb4A
azA625BzlHyF50Dn4RyVybJ9f2IDREA91n3JI25hjp8OgxGGyMy7m2VPPM7R
sFprGXbSt0Kk/XqjlVOYi1FgsP8Tn0HnVP80jLPcd1FLcdYQdjKXWP80dVR1
h3lEToCucx0LCMUkIyQEJIj9p9DT9GRYdOEL6CK8AHD8DTEQ5nYT0nio/oNx
Kvdt2QpYVeKpugNQ1Y6yS884KQCzfjAD+rvCbgA4cliLFDt9jaccM2CnqznD
VOcLcgLfPkJVhQZ+QVmHTrxcsisJLQb40RUnXe/eXFGFxTI17tUrrL1KxKoL
WoXxRhlu2z9WGhm6Zb3PheXzTKJft5pUibDlbYCsMzGzKHTQDYnVSBzch6dv
aa0RU4LXZlI41NwHhmW/4m1gKNlpafLoBW9aDcXqRTAQUeAygnqI9A2zeuSx
IREK5TqlMc2C4fl3eQkdijfFHz30YFTQs7QUZGo0s1nYnUftuYDehqsI4u24
8QMU0p6Yj3hJyNg/0iurZJCne8cimT/g0FvP7fulobeCSIZanzJfmqOX3HJ8
UrKDUA9ISWkmgHQnwOTZfrjnARZuBsIz3NJUt+qNOPTc7ZueTJRVpyQ00roH
fX5gNkHhy0APgMo5Fd6S58DfWYEK0wjMqUzLBaI1fWXxPORuytxfCx0ijy/T
oroCQcD/63Y4Zipn8sWNZeG2QeqRofOSGgu4/enBESJE+sxyqIzyiK4eNiBb
3TybdFZkTUHNn1zZOsL2WIcHthepUL/4L8BMvZyv2znSAuFE7rMQig8W3FfO
FiS3iCEdMR7y9ZV4MkTOiu2ghAyoAJmWxZAeDZd9r0XyBReb3JoeY1oFbtSw
ENCCJZayelCft721ziKMVrkidG/JtZhCziKGdpyXjsC16MgizVkfsP7XafJB
ReqJkW9zgxMjkbeaXU6HfePGrXP9dt+WB5lDy5syt9T63aeLUFR+t4a6mwdm
XLnlWQrABiKabEu50mOFMweJ0K5HMNwTBAKzJMTTpuOjLawIRtcv52o6fN1c
aIZ+2RVSMDZBQwyMA/qJC2vFFH+3QYUUNn7qH6zpsX9UoOCNRvBrF3wK19n8
4ti8P8CuyrSh7/3ek2RbU8P3efjFJvWvJcrUDkmEFhA/bIj4wkCRqiEejO73
oiJDKA5397q7UM+9rl8mt/8LHbJBuLJVqWkLqvIcEAwjbJPEgVILg575ylUp
jPHqpfaLGax2kEzW8fNmWctYM2M3UypNYpy9Dj9pu33OASZd9miU1Wn7Z/o9
QZZ8M8bbt9L3HK6V/nRs4Sd28yl9jQyWy6t7OSKnUdHY3R7ifSsSvB2D7VHO
F0m53jct2Y88VzsgZj2jXMPxmyM8oyVvi3+hUALPGRAE/EO4Vms+HUn1WizJ
Lq6ggS5lr4KHAysaeHNSD8EBO+YTMA64UCozxD1M1n8NXd7TgWvRdD7xLaZI
TycH397wWWMkcmqrybzkUIovBbefJ8+en2uLxRe/tYghXGtRwECHMwzbhvjl
KsfAwqjpbWBLN6XbepDExFduSgnyDi05PT8Kp3mXj8xDHG8DiGyTVWVTftqa
9x3HtLXZc7u2nvv1O8EFbO/KGitWILGqc/2UqTwGb1qVi6YNkzqMOBnNVkZX
/4cNMxeDgPdSRzvO03lTRAR+ptBWz1CN5VgnhAQDeN52W6jBi2C+wmL82U3B
JQ3YJ63kMcK6U+eFwGnhPtMumxgxvLGKSL9KWTHz/O+8/gvjCKwsmfCW0jp9
TllRYiP1ibs9QvXWsD3wPXPSsbw+yv4Wb6TKAEK3xqKV21SV/UYEUuMZu+OV
+nxBe6lKtSNLM8zMZelX1/5TP0boGeIKXrbo6LWrvQ06oNoXXBvIOP80qBLp
akufAKW4FHGE5QRSXfnzX9oIKvLxO50WSlwI+XWhkpPtL1lNQ/HpY5fLO67Q
zSqTdnV1J7W300ZAepz/nWAGdEX1oGnDPKV8WSP7CpSIL3u9/Lw8CfYciaxu
Ir9/Q8hUKc0uFnpP55PbCPlvRPGijG8raX9+V6Nb1e03TLVqn7fCNNFYKTTF
EyMWbHxp1Sly3mHFvTV7V8VRYxbs9tMKjVbdxifx3wVNGM/E08TyN1eEFPoq
c+0R2INXg0GgKoHm5VVd+j8ALodxfGsNY8v45sKfEE+4GEuGCI9pFm7Io1+P
t+2iCvckjmw9ovYwofDjT3BXxlVuJA0Nt9oOa6qP++CExreaPOQM8kfIUnID
kgx41JXoxoF7ZKGHX9+wBmcna2q24/3TZunq2Kwcwfv8I+7FoGhyDQP7V7zq
tBDT5ydWMInMa68QbI2VJLAYhMDj+nt9CZRS8rdApwLPWBsxJFZ53p1HoMmf
If9wnAZsAhzTDIVntppVxfKNxApMOg9TYIg2uRa+Hi8mol5ZQoM4DaMZjTXn
WgIj/beIKAHOoWxwIJJpNy+Lo4FuR1ierfmpjLKFw/Q1L4ObJE5W8JptGTT4
BnF9YRO5bY0GJeCBD1/pINdgyNc5E/38UVX8OmizsjkTW7ktS36Lht3HfXQc
LbSiaz4PMRKgHe5cN0Ls9q7kiUw6AuW/ZHrwXgTp1wgjeGRGX57mhiA4J8Ip
f7d8MscipkppLAqMkhBdhp9wwnE05I6X/TsupxyODOcov8fpTSaoOYcH4hTI
Ed11T6gQaF0/k0E/ZTS8CnBGHM4F7RflWmQT++1/18WPrm6VWieMfeBzLgwd
2XI9MAQiIfjNT0XMMbtF7624EZWOVl8d1L42P77e2pUMrzeAlPSbufR9c73a
UGRVO5sdj7FgjRHVnVHl5zzaFWS0tkPzW+qnHVhnSHDYQh9MjrYHBohk6Gey
LAuskw5ZQdDGq4ocsWwUpD40EGvKt09ZIxSuieVU3c5H/Xu7deVHNluOf+s9
bFwph97xR+saIX8N2cHAA+yRqoVlEchV5wktr9PWNvyqdZv84vPh0vHfLZ6a
EdOOFtFvWndYip6vWyLc45Piz5yWTMooFLiSlAGXy/qtIax3Bz1Lcn6tBy2H
/Hx1jBOydMnx4Msv/MPyKlWh6PHHbW9cJVmRyjvMRt/NITh3noqAMB0XF9JV
k0Ad52YR98lV2ZHdmuTlz+DTi+kNwsM/od1+siqJa39Z2U3yMeJ2RUzFTJMs
9nHBf1P75Xj56EqdjniJH1WyNLYmJbO4EiisapZnFga3Yx/yGlEJRpIs8dhy
FrSvz62Ih/x19EgEA7Lj43200ZQUUQSAfS1Y0FoH6fKXzt9kUN9Qyv7/aAvL
b1wLzzNTSQH+8XKlFIG8EtOx6dYvZltPFmVBUi+lkh79FUrZ4x0AC/AZ7c7Y
WzE8rjiUc8r3TE0Wf4rxPWF6ksRoJAQQ9oe80nCXebj5XiXo3bt/TpfQIwOY
QUUeaLW3k66B4KRyx0T0eJAqIF0WGwNDCE1mNT4lRqSfK2qGzVYyMZStaEHu
q3fZyZTD/SMmMvXs0FVFHTgs/WmmFS7TNpUd5QZa4btuM3du0078RI/fQN3J
puAvmN6oLRzBY4Bwya7Nwqj0tK2fEdbqbqlKcmgDy4QzMU/kquLgdOESodFc
ikDKBSq9OyC6dVPRLT7IVA1wU2SXP5pWFj6TZ4yr+5gufPIugOPjxs+S5vHG
nLw10b0VWQoc2lH5HebuPclfYgUGBSS0oC/U6+AAKJ9xu+SoxI0kPCQuGntR
v7ozHBp3wVMb34Praxfwnnj0NgFNgpG94MrDVOOQHn/7RNjPTWNCsG13yYTQ
//Oni9a5dFpW+DSX4PAupdeQ/5pUKBKHhK0kVzoGx0Y9m8Sk0sBwCyU4+zbY
FP31cLwLMjHC+ktBZLBSh+Rql7ciBN6wLkqX5jRoA6hpAuVcjUhvGJ/j5aZy
qSGeE78H5vC+JzEvrX5XZ6IVJ0OWEXkGxJ/LFfTn4O1c8p/ulzQfdb1292oz
16tJvksTJXLPbrgTuMYp/1iFhlyxLYpiMvcaCwh2UvHeDN7WpOdips9Kmeia
dMCGDBEWDXjg5A7KQFbyP5sPSpBqfzosymwt7VRYYRRZ6G3peIUied2ZWd/K
MqmTbzASp3HlhV2HXFUuHnK/rg2mhybhSik+Nbhk4d38OHtkWDqRbj/GYrB9
4cAbIJSvacQ2n1gwG/S8OURKXRJlX1ZODXpei93rpgJ2ksWCvXNoSD/hTPXj
TEYnAF9kMct5yMISoT2xu6PDHksqsKANFEfRuTLb4YaaGr5eQE9dkNNsb4S2
Xl/1nWwzw1AU//py5SAsiY5QYxNsJyEixEvXF4sioS2EkUxnUEzNt6AtYpa9
lKxNxvLEkgQfmhg3O7ikVFkmrFsMT+XDuaGap5l5EVph0u2+DHVDgeUKpu+M
shirpCKtGgCWO0YlwtVsTvXHcUHEQc8v4CoXQ5moUy4OTCTHMi9SdDDj3zdM
ABYYO1L/pHvdIObFTM3nZ+im+C4Ux2KQ0LZeo6qhPZsHu6/ZKIFbCTmoJGIu
P2lYaP3hgHA9+tklkj7SdqW07n+veLFAxmizAtiK4D0brek7NrAJoyVkRTYM
6Q54u0t5bkUp5vEsyFp+44iQNwZiFZsdeSLai2NOvMVqEzpiyXSs6o4SILG7
9dA2ArxO5dEElumL3T8jWTJSRj7NzmxM9K55Dc/NVYAI7K8mkm93ug/BRoj+
Jji5VQ/pI0zXPrkhIY22EAy25xdOZ3fbnwEYxe7H7MueUPjPPSHb5BiMJXDA
NStpdlabp1UujPfgzoz33SJtuteKA4rfgy0yHhdHz9Fm6twoTC/6+6E3tjOD
ekE+3I5R1stG2yy17CSnZ9j76U78YmDqsSsudoVWZy+P6B2Pd2va8srrBHYQ
Kojxm3TpV58bkxqQUFMQ+1TV9yi7WHRP3xb0YOUAZ6SpcmsM3YgGJMQdjjMg
F4+vgvbzKf951aemZ/fZ1nPbE9akUdLaeoatpbtIQGnvaQRK548RmJL5V3qt
+OyeXUCB4BT5VZk4rwYOhWEbkFrWt6bM/k0k2H9kjdvna4xVOEq+aI1wZKWH
jnund1/VcmmMa2hPzsLXKg28VoYcl/i7z4r55hDKznYpRIeqIs6q/XlVQVUQ
Fh+hJf5VRDsKq/tjS1vLNV2C4OG1faR2mrxrkM/sm0gzoqfKnb+XA/jTzygA
7Npi3xrLLav3U0RxgIhJWs1cdVLjo/ydIeTJXmFu20pCtt018zS0l7ED3taE
A7xOVOQybm3+1Rkd0EWhCgZib9Rb+JWbSsvmCQNNksdsnfYL5m4tAyEHDoGf
AQ9K42Jm95afJGSy603R7e6Yol4darYzb2faE4oTDrWzNccz3BJRAwvwmBw1
26XfE4ghzUg2SNGdFhXLR/itw5mCNx6lc6VKoRxEcZiFaOiqkv25TIZfK7gI
xr8Cj62dY3hEL0ui8aVWMD7sR/3ztO4mYk1AKZwU18qb+8IHSA+NX0N5VBRz
EA8ANyZvDmiVY1RTSyCgFQbaclCwIuRvZ8zJxt4fJ4lnVbD0ghsnfh5i5U7F
cchVxlhaTlBX83YkSu/CXXba88aUXBd9bGc5CIXPgMfn50/NE44I4e8b5G1E
/b4pcxUGPPs5PVUKwKhNNjwnXEJWjjJhRuYd2Kl+ffWs8kryrz/8alFJC/NR
qDMCfWZ6YqFvG/2ugNYIAxKXC9qxtf9+RzWuzK2NJ9mThKkAkq/vD0kDRXEV
hKzUqBQslBZ6K4zuW0CcXYcdIeJ+PPKTp9vsPUfdAyBSkZXH6n6Jo7SNte9x
b8CxkYvKuMPu1iqw1lBKKdKmwOEhqk6vihelV7QbVQ7/Tuowgv3hthAwV2Y9
q0MVrzIyLI0ADWOib1sB4CrCy0CWEjOIRRPOJ2Qkh2FVdbfxunfDWmBCRk90
fvlSgaN8ahtxoThIpSRojyAp1wP8RqVkPabQPkBmTnBaIqShgVJhBaNW+K+V
+S5eWiaCop0HVksRjr4aOnWdTyGoOXFJPtYbsQOfyqDkdyD0CkShPSC/QuQR
yNX8F2LlBa2zCAXrdQ63oRPIP0z7lemnZxdscpja6zhyhHoAyn0wCG330aW1
fqUo+FK7L9fdO/edodzW15AGABeljQGoFQ+GXxd7VgHz1Wqd3g9FMvkdwT8W
RTkngqfZdXwDgzy7xTfH8XjwB/8pbHVsIo+1VOf2y/m0kHmKZs5wnJ1OuFvH
OPQIJP/2NKQDxTOH0ZEyA/QdH4oQaEBeGDapvsFhdQYDqkzN4GECQkmb9vEH
CFGAuftxpkRixM+06s+lD9Q3eh7FQmX1OwwH+v2i+pIews6mORQ1W3WTQzva
hi0MlSoQlHeI0Ko0J58Nj7rRDmisFLYcJZg39cWJx4h/5IrXGoMpnKc1vYgI
okhovubFEP92upN5oNQ5Jvx5dFRYUNiLbGtg7VdIgmnm6XTERXCldh4O5+Rt
shiiIHkYseq1tIyqSXeJUf8i5JIO0D6hMgwlAUmIVjvSD4DTCCMcSXOTQg5U
Z5eFnKXSxjPM0Z6O2HG8UK48icZMeTjKH7iigJESOGdHWVHHXUfGhKoe5Lyo
FdRus0C8XMj7A7KkxFjcho+e7i3l74PY/gbRc1a2a2UbWv7DVIghRSFO6L0/
UQr75WgFCpFOb6gJjl0knV1ZfNoRPmJ25xB9Tim70VnvIzZj0/TRk7zegeV9
iCHc3YeB/c64Y3zvCbkGSsHK3ZyxGub6sf2i5wNdX7HD0zLLuFl/KHD6AKD4
tlllxyf6GnKeIumI4aKYRb6tsMZzosu7gC0W4ybEfXfa/d61UbCH2ImosCWH
vZepG9QY/NdMblxCvhYG0MOBm2F3do19Pcf5V+/W91UAZ4d40DkFvAYpIGxE
Z2ZzaNUnWR9/ZsEAhWI9Oo32YL/PlE4cn4BR7bn4BzMoXAK0rsMjQTw+RJgG
YnYfSuVCI0nDLAuWoEjbxNu+NjVQBiAcHWqUMM+AVjyLldQUqn7OMwYhlZqe
yb7hX2PZymuzXKMUA/0KlxL4O/OjMnxXNu8TPNIolqImrer0TpYUHmnH7kxw
rV8kXN+Ub2MKgB4s/4k+O+3z7rlvjv7SmYzJesyhLXUvuBwr4mjy8u+0T1fq
Q0JKpomxT7TSfGgJd5QCmbZy6NaWIe/rKgeIHGuOBZypEPbEEsLB6bNOGekG
V0KFFfl6aor02I0vxqKgmtnh+RfefJ7AgAbCsaTRM0Asj6XQgAw4tsaOj/qy
T8tF5MdAltpHrirKi9NgTV4L1jstXqDFFDmv0JRO149RtigiTos1Oh15H2xR
5CW1YwFL7d7RutXCu45GNea0qgLxyVqcTGpGXDzt2PFWmL4tokUdtaba7NWt
vfSFc/RRG+fNwIEZRzrucu5MkbqDqm5VsPNn8KFb1hv+bl9ckyA4QufuXD/n
WtrLSy3SPePuWHddggLNX1hK0j3OKmvvl8JfKzEMesBTbCcRfjIG7Ds3wH92
lIOWVS3TmpU13x/xhu+L3WuCi1603kYX2JWqb9SPfhxRZ1nLNto0xlRzJ68a
ySBP4yCCNJRqCyKCQF9In8ItQWQ4pGWiDrUWBcw/CdUu6xu97dPdkxLq0LqH
Lnw0T16D+IPxe4edk+MUdcKQH7kL3N9BOHeMGbqEbyyFkarnjjBxM3ET/pZW
Q1TLhoCmGozN2fi8eJdKQd7qPcOQijH0I+RZERmyomKs/XHbo9p7qQpcWbH6
20rQuNvjqt2N8r0lnqTHnt6jj8gqX5tIC8PtGTWU5uTTdKXJlQq+b2v7K1vd
vaV9cVQVJZUjBALLvq7rmtdi9ntVQUChHmXAGtyvT+YPcXZsKZahbB34Jbwa
DgF4eGUHEWqMCmZ4BIpUitifT5nr5WLRAc7EnP3bDOlhyUJDniMECziJokut
tgcKe1S0E1UsZhitORQUPOlqmpmR9/oQiWslfQfIoRDLkgkooi1DocYzuGZT
ie5iQnR9yaZtUxDqjOeyuAWR2LAVyaxICXqomtIsmUywqzaxplPxyBNj4IXG
r79EfxPTgdWIGTv1ZJYBRpCFT+cHdifSCmJrkHSFZKk51SRU/xXtHQueQP1o
Bv14waePdOhOWOf21uZMwOVYZ22hmFeO4RPLi4M8siNtLmnX7uMh7nIcsMvv
bqGzNwAsvhpP4H4fi9AJlcUlripryU+IYRQxZVsfR3H6CBDNLDNqD5PYo8Cb
R7DSBcspE1q6lnJnZIe1izf2Ndqbughn0lfXxpY/M7XwBcAVd+7DN1MNctwi
u/r8EOlX8hJbEpK7A+Rhs9/NOP+FDIGSCXYcf6Qwwo882RXYt10GhYcy9aV1
D4V02LLXtnr8Fi4WlnSVpiCoKEydrgzXBRq6+6N8g3R/aXejDvOVPMkPq07d
MB0phi4IdzQwPpwl1rDj8gs7hQqMffUYDI0zBbGeRfdSZAVekyP5nncAburD
XkyXw7MVgMKZZw5R6LlA8Fmkanm3zavIoZTQrqsVz+XGJ1nP4569XkeHF8rZ
l3rSJ2HfWj/DXqkHlWfRDHJPoZsubqk5Z3cTWU7paug6ofvIvC9sE4WJIabz
Cr4S3EKmZ2Lt1ebj1U9nJzWXrEQ9BuMTFXQ2KfU/Pw4I+y7q0M4tGI+GVFSv
ip2Hoe7bFBi9uD9o3ecS1XfnEKhH4oBcfQ4s7dKmJey9y/OH/uyAop8TwclD
ADJJd9a2XkRjWuH5T7Dhd7sAa/8m8a5rfn1cHAf1Pn8PxiX8PI9YYELyClTP
QzkZgylb8/75d92yC1AI8WJAXSCZcLnawzG1+4qHehKAjlqo9zrKR+AlWgb4
mkKX1sMTn8tlDsR4PN8VQCVHZWV1SlDufWakXxnwimmUsOqrVIUtAvCTGBxp
amXjlw06aPDX7OFKf7OiN2upkaz50ah/L7ogpmF9wO6CKAKAI+ZxwbTEj8Zs
XrsxtRslC0zWNl7d5GRYzwA62uh5l4sE5zxt7urHqReB7WlMzaTxDkzPaq2X
EyCuNQvFf8CteesDIYtl3Cku+cKWhy4N/gmtKxrzWVUZe0WVnljFfi8bt+qh
GnTuesvtqIf5sYfRuVXo1ugam+kYLJ5E/f62YqOq4Yr5Y8PbuSyyzb08kTe6
SnLoJDEknFLQKOBq8XKGVhQSbvPiuJ/p8FCp0pIHdFrL1TXLQg0LAcAUagfd
pSd/6BRMCuPU+y42sv0byhBddAM3GwhecE5htiujrWMRC2NU3KfH5OnCugEH
4VHhk+MMgTNuUfF6mEXewrzqeRVyNc6OFYV75ah+66tVmsM314AxYDWuHV6F
HguZKo4prHLFwSxw34Hy7ma/kubAgdyYapD3WTM9qgyfa8oOmYTkX04tHQSK
MLPXQsFF6ArPuFHFUyWZEidXSzZotaByXFmLEx2w/+cJAFhlsRV7CHNraM8T
RKYZfGcb4pPMgCjQxRnyRCrCsKAEljSIhf9E3kl0ZwesiPK7L2IgDJvYfnm9
nY+nmILtxgNIacE2M5buerY1l0NHfuHZqTynwEVz90QY84/lrztx00kw5m6J
QMIFgVc9fVzgH4ARJHTKHYIgLLbxqdiDo+JQdCgyDTFm3J5AfDnYEnr65weD
/rV9ddVXuY3VIfaa52HU2/4AXQdXvGddZ8G4z4k6OLV+ZFAjdBj5h8G142Bz
cXKtI64ptZECUgBM1rObl8Iq77FV+3wA4/IBmi/GN9wzxHjLinnjFENqaeob
p0u2Qz1l6/xT4FwPJd/ehAIJZtFX6LtiXuPpGHV6Px0pxLLfHc1/dm4k0yWl
FQ7Phr1X7Rdbrwh1ByvrHij9gOZ9LEXiZwSWbJ/ODNyDS9nwMZV8PNKwFWNc
W9+Rnm6df213qd7ZzxhADiZUBPjl640XjGnglB/kDfG5IgoRAZva8Q/tkEqR
/XwqgOK6rB64oW/r2AJ77hzmoz+bMd0aTH0uXpYqAKj+sN+0dtKuBtRAov1R
0WDmePK82nvP54gqWgT2zhGstEpA8nr/oq/BYNCJN+N5Bo5rCIKxAYQT4WwH
NUPsCx1c3Yhy7lWA2O9iKsumWxy3Rt7JRZMlRZsZv+eQ+MluMCArXmMEK7ZA
cOnoAuYN9AnMq4X/tJO+Er3peNJZm3fcK4t8W7iLz70sIp53y3NM9nxtRcJ7
bjHd+SN+ocLEv+zBAoBwcbbkUhVll2//SJA5mjc+TT4xZexlWMtYBjx7SiPc
iJQmUkG2p+vVtD+vLA7ezxWzxXRz5yMWjUwSoMG23SdXIi1xzH7Bpv+MZHI9
y+kC45Jvp0yibZuG2OTeqMzp2AHWHF8Y9to/LSsPf13Q52uaQX0lM2YYT/vn
reZYmOX4wY9FxAwyfDq87auDhjSCUUkO/QplThEF3Xdcz8ewUnWmg+nYirxM
aH+o/IHxYy9QLLXxPRSgUgVjIEfymMMHr0mjQ4/SY0cq96536YO2HAfYI3WA
QqyG6hYOddsVQsMyvtvLLIR8OwlhIdW6wKLPp6EP3ue7kpHacz5Q3qnqzV3i
wACOuPrjr4bYkZDJ6lSvi6MfX+6wjER+5+iyJt5/7eH2f7F97OklV7KAbq5K
JMPBABv/HQC3zmoZP1jX4j7Ng14uJkFO4kqrLzFrOh3aYvRJfm7TZyf2QYnP
h+sRmYA6rETFQ8W8Vzs1N6GtebrTI1yk9TdmolazSCipRq3vC6McK88tFCoL
24FDN0tPiEH3yF0P/u2YkNvNwzpz+p1ljfqoqnKAaPM3hnyKQw3ULk01mpeH
BlW/ep/uP30AT6+OqxjnWWJ2IaFQ0ff6D7lsCA4KfOG7pnd5zauayxIbQuZ1
iQxgjxtZVqT2VVH7VheDv6Sz2uLQA3mu1nugQCWg1MyHnWlnI9phNoJQJVRk
hoYB1Pe4hBBEJ1FwPuZH+XvJ7e1Qhdx0Su3QTEDL4OKc3aU0TTdOVMdplMRD
5bsB9LvWzqZMiK7wU8klyiAdd7+qqWyDmn0EWNN8+1HX0BEDuK5Ucdp2J2hN
jNAHdTZqpmOgeWaor8D2MygfiIEAl9+STVAbBmkPP1kyCbfGT5a6GqgEfOOF
PbiqneNhYk8lsZ2wg/a4WawxamvuQrzOsuXGLL3rLB3iRIsj1Vq9zymqe76x
ghTsDCIwVGvvNXAi1cJQ+cVRVyM6exMDKqnXshzp7NJFlCPT3+Q6ugZrI+F0
7lrIfL7vHnIB5/CTdLVVb0gXhin1m7ZtRymCkK6QrryPn01g5Ob/c90hP5aK
3+h0RYR+hyxMDJklBvaWgJwEcaCCLV8MAYe5oT1TOD+PN96bp2tuaL/yn7Fm
DAYXNPfZ+YNId0RnU6/w3BUVaoOslcCpZHbHGFVv8m6KgWITTElt6A9LC9nx
1tTT1z0Gs/L1wGfIW5xTSg5A4tOxtFkWitgx5+gWI1bDoXIBWxSuB7PcEGKm
3u5Po7CwT/yhpoc1VPgdjh5wjHA7fMFCryVOtwXLlcpxlg6SGGIEGvjDDgOD
ADZfYOt6ZhV7TdtpF7cttdHwu8FN5vJku24qbH8IO0+0vZ4Q35D/qgL50gCt
W/I6ife97v/mzFXjlynRvULEOXk6n1bm6yuB7rDTlIY5eCs5lCcPy8xcOw3g
s0ur7ueAREPOOeGb7uEzFCvJx7J9mUgOP2hgCnshHPWQN/zllfvY8GfqrptC
sOVzKyz7gwZcoUw6wwxqfH0s9MxxjKtYXE5nJbGFvC1pJ9ny089JGwB1mVNj
9VxbJ43nypTCxl3ICCARBPLP6f7iVCo/agdV7O7btGrjc/71PmRVx8Ke5Qxb
FaQnVb6XdBh/VFectYIdqev6pHNXOYEgwnD7NrBJBhFlh0i5mM7U80OUW102
u/sz9TwRKzoVe69sZeTt885NwpUJzrZS4tlhli9W6eaAtvDu0Orgly4ZiWdi
PennrqIdf3BxNUEeuet7in9RyeqMkJURlbVnhUaAHIF6jTHcq/K8W3svcGiT
67isJaaIh/zhfrt4yc5L6lwqbf6SL7deGGwhiwJnUd3wPKPtpCcaZIVwX2H1
Nss8a/RWif05QaiOGmdNxMbXQhCv1om6vFCyRWGTfHCbltnUDT1GQPS9zy93
RXWIJQlN0qgSsOWOu+7B1+zjaK1HLaYKSSDVwDLmqQ/Gd8TKCzI8HQ5i4sy0
ZTG0ifn5eS3JIMhXdiWqr6iqw359L7bk9MnjK629j46GiJNlcIWBQZeYY7vn
h7LCCiioeOTU+fvm8ReWEDfbgvyfj/Vaiog9sfzI2+rF57u9vDnjNpfJv1mo
FkawlsptTnH2mb27AnpJelx088v74ExPJoZlRQALO3o+yVDlgfuCNx6FGGQv
1PJiKvfRj9fbbMpd8z5hTx3SA2DWwI/yzSQyjniSPmL1CeP3qcuKsKL6KPMP
HY1D/4dTrm0gUNOLG46RH7Jb13lYczIpOhg1FrzbYcvRRejT+zs45SyENsfz
BjrwV9JKnHMxtdXA6ezMxLz3XtZ/hNPrU0ks3AIe5mVUDSKga7RMXmSbwRfV
n3jv7+6g7fMboWKQXUgFhB0abXI9vxOOQq0JELPKYVxBcqf1D2CTWBShXok/
upUJ8OEuKeQ7JvaO2PVlWTgc5CaHir8ITa9j/vXwFFVg6hkOnjLaE6n4o4A5
pKnv6uUC+yrRFZYngyZJ7z05yasOYORAyaoetxTuSrBnuF+fZdGLBwIXYNcc
rr3nQCxOTCa2ZLP63ICoL0TJ9+vS/+iHDCwPxDzm9eDhyhh+7WMFvLHa1jDd
zuiuh/YjYBrHU7Xduv8zpS5xk0JqpthrXupuTHml7sNn0Upx9dtTsws/b+tu
ZXrwXREcCkV69a362Qi+p2PxbH5Nhtcb5Cq3aF/8F0a4RVfNg2dtV/Txwiiy
r6KDIh/ND0y/hVirnAGHxB+vXJREyj+Wq+eMxikpIDtJCBwyu6wMwDdSQiRs
apuiqo/m7egi9SQwmj7SqD5ojsf8OaYuuBwIKdPbh006r/ZbNIoWpEj1xGpu
J8CY6g81GTMVjkZg2KnkiczJIsDIy3KhoB6z7/rDkH2Df5x7G/x9BPOGZHDf
6hR0GOXZJOfjwYr7kdawxk94GC/78kzs979UIar4qnzlxgINpOLCKLfFyEku
MyWQb5vjWw2n6PejkezmWLvEmLepD1DPa+lVHvKPSDFsAbwHulm1sD/3cnJ1
gS/Q8ppVYKFpRDBvnFesA6mPQRPXEX8JpgiUdmpBRqPII8WuIA5I03d01Plv
9WKybGXQj1LsvqVXkTyED29bf9i35HIT4mPtR733BdEaDW77QwbL764sYruX
FtdP6zpoWTRm14A3DodruajooPkZ61vSWvpzCukw7Ggl6yTLLNSDsCeNTNmz
ebLHTcvpcC1qeqGuhUbWn3ScOwsJXtJYUJ0/ks2rGVVaQ5yB3RmGc3ZI9wvI
bIpvZwY30/ie/Upq0YMQFgtPVOLN3Qm+QgTlcBdMo18ZrvQJEYT64Tr+p4GN
Z3EZQ0R+QDEsAmC7br54vfwsbAUu/43Ru5GqhUNXmTRlGyVqhP0vVI6QWtm+
TObYeQBl8a1XZwoA6IzW18NCgLq/1ZsSEGW6tPQ4gfLdMu79uUdmzxuJUNWf
esUZLeFsrMYy2ICFclkVCqWOS0kE6QksiJUe/wIBHbc2xC7vioNFX4a0UVa/
MqqLk4f9yxQqKp39AiMlEHIOtAL77UmAENRZygaE1nXvcQur5BH3tSonrHiY
O6jzYKm2RzMNtUHlhzr5cMPjhnDmk+O85kEIgXx8m54l/uLLo6ag3E48+L+2
yFGKfWRxqBLfBGev/g91tgEqXOnUmf1HU2nGjDAeFwIbzueZmZKb3x1Gwz37
zWa8vevjjTfPz5UshWE1PmPYrD7gF7jzspEJ3KJow8Chk/GFdAPwkm7VYPNs
VliBJUDrIPdNyeXt6OKqYFxhrAFzrOYxmu9YNqN2ZFIBBSQPgIXM0t4F1f7Q
ISIO13+6uc0GdY82ndL0OfXHmJc2AQfDe+N9H22NRmpRXSL3y7GRSmrpUKC7
qH+3DMSf4qnIV30QRC8alDMoBoM/lF6sTGKsVdQf5/4dxaLlkLqF+QsnsW2G
7FE6a5C2MebBAz15XZnycaKFIC63SO8PN5R3FcPPeomVYq6n6TdEyxbYSk43
ieoA+DPEyyMVrFnv/yHLePP47SjzbkE3DIMVxWWZLbTqckrmrg3MJBZBPTnw
pmy1UD1G41O0LXTiDsM9az4MUQwtaKGEBSetwV4GswKJrZroOJrU6pf23FSJ
mezQ4mMLF6yI+N4jdQ3Ybz077Yd3IwYFotRblZjOVsryYqiIlwp8suw/Oz4a
9V5RHFeyEG5wb+LcFpWYf0mAyM8P6WQwIBRzwAMYqH5w0qywylhajWJb9iG/
VNHooMAL5azQ5TgQqeFFdkflBKQZy1xp3+jXY0fcvyJSDbeJl7lsA4ROIo1p
XgPh6s2/AFf0JeFdyL6gscFstCMW8K2K52PzZWNeRWSq5KhzknzIvmW/1/Sz
xv+OGFUoIYtAgV/R93mYQnPAThWvRNz13v6PzjB2ZB0RtBlsye+9yhx1ARqK
AscVD3hwwJaTx/b/hQnMECA473t3fCkU3z0gSxvPoy5+7bmHbxf4fOWyjeDf
xqps10f0pSEjSQ38CBYhMqZCwTCyStQj2BiqKCCVrw27PGqFt6cvFwYheNkP
mpO1vJpOok9pCnqgwan3w+jbZIxVObDVZ0rA8uaurpkgEYP1o2vCMKgaTa0Z
07bTmZmpRF/VsAPPI1kOQngiDvp8vgRUwxcF0nut5JiMUpNebRpjQy7ctWs2
rR7fOpUpLe2VyTeL6lL8HXsuAE9wEI4O26+bD466Xb7R5+RidRFwSbIDfNEm
BV06373jAGnjIgOUex9mf/fD96U+VINu9/AbdylWq9sjnQedTK3eIG8WSwJs
IwZtiqPYvV6k4xj+0/g7tkSnbx1qs6ksFOV5O+q/xCMh9+ddn804OcUpbiXx
fk7mRMhYLfOpG62UoIJ5A1TVxI4Bu7tB6lVLSf3Mgh+C7simEOF2m/yUWZCJ
XXXKQPwaZGH6eXTMGMdOgl85ToYb8Ds0nEkCMUNdj7enz4fV/Nv+1uLbozQT
q6VEpaEeRvgnjlSkjB5wmzM3Y2o2pZpWO3TNJqhdX3peXMHGalFVSfu9mnpZ
m9OnPNcZ478HD8IBTOhxY72Ol8IfkwirVN6TSiyTnW1bZnFiFSxSnmohMFmY
liSUYvEbSJ5qxtnapG8oATOmrXfbrtGZ+eBvykTigiNZmeK6wiirCuJOHN2W
be44J/EEiGbqWfQE7LzAyvAAA8q93Ob3ckO/LdFh9nfGGFIU6hkn1GYMdIP9
YbYuL7CBKnqYnSlKCG2pSn0jE2bx6d/RdX/Wo5w4D4Mz3JfGj6Fc6etBrXbz
CSOEWz1H7xB4WWG0Rkb+3uUTnnjU+3Cw3zkau1xDY7W0Hm57bTUnfuNxYx6v
1vBjfDnJXT+yC1MUfWW5PPgrYM+z8j+5HoWoxryMq7Ywu3c/ronYgMHGx218
39DQUCrhw9jeI7AKe4WnDOHjrTJsqVUCefyixYxx17SDpkXSURWS4cxsfHNm
08FvWxHjtkLvgpaUt33+W78oakc2vJAskob2MNln1gspCDMYWSPxshqFAgPv
hDGgJNO3rdYqrAV7r4FxA4c5RhpGCVFbty36s5Fi1/7zBl3sCY9hN0WsIJqH
sIaoZsWUFz+xiZrX7YAHS3tL55l2IsPrfbKo/OO7ubN7iU5SFREbnvJ0ZJpT
TuLVuuFFz+JKdjeWE+1A3Bl9Tzd5/MPFss+Mg/5ITYkbE25JebK9rxjPPR6b
PppY1FqG9PcDFob9N7QkDpTkebZCfzcwh+6iKcBy27RWo6cWNGM1ntu4tYLz
VzTpw/dUuNBlz0dWKEikL94ikl5foUtzQev09+pxyuMJ4S2k09NPrpOpylx3
DfuGAjRFgdzoChUw+txsO7CQj+/QzGy6OJPO5leBsVjRzS4vmQuHQzXbh+V+
T9aZO7TuEKrq2ZHZ3Vdzd+BOy4JfTWLesE6nIgJppR53uWWzY8YHQ/jJwRT+
lWTL9Wl9BQfIEO0vHgEM1sv3rhmifKrPhKKr7BFcWykgurIAVornQvNbMPKk
gDUtanqJ0zu+CEuAfIoItjsmSKVBAMC1gUoON0C+hcEsxosnFDrYBVgMrRmM
6e8vQ/jLBvt6JuJiK6KuWSlT9hoqqYT7zah/5UfjDSa4GZD4fEHgLxGJ8Zwh
j48KG2YLL5fgOPtTUcClTZ8FtueA4oKtX3r7vChrwx0nELrhGSllDUEymZyF
C4XOVdKIL9NUX8NeG64IR/QNbqm54CcFER6Ej/ht/AdQis016KZEE0LSZvk4
wktjponwPzi1HM3snJ7e5oR0ydpuDwJIO/TI09UAzPlBwOFLLDNuI0orbA6S
CL/wSDBwBUmgBv0W9nMwtYDpRGGJjgogPT2Ekekqoptw/LCkBJOuE7qPrniG
AJ/SS/Eu6NNjsRAQxVy4ghD4FU/SfjKFyaF5Mc/j7ghlxH9Dd+0R+ZFW/W2v
QAhrKjjzIXVBlc2PyyQHd/rDEHt9kHXynJaIdbTRu9rzHgJspEGIOjoOC6V5
qEsq4dSSbq2a1E9Y9O+bHT9aCcmmFFTUzQcLeOAE/8K+nSCMRlVBOxPh24LA
zrgsmJOv1ohrA9VxuV2yTRkZUp/d4apUenwk7b0zGBKVOO2T2xs2+EOr+P4C
GpLTBKQcdcBPEYukmRS5nCOMgvv+9zqHcEOk9waxIdxNesjBhb2PWXceqW9G
55+6zN0kpYfAId15SqCmm0j49PQLCS4iPr84PkWOPQ9xSZm3foPZxuQ++H5G
BxJrAK7boMSwyj5yfXJKqB2Npo5QupYJ+7/7jqLpvgmRPnJZNOol0kk3v5mG
YhaXAZ17Ukxt8SJXG1bw/XmOEbCo5R4fp4ZZxZyEMv/ZYY/f7sphkSpjvjmI
68jYASCpHS2g34GpWLxndtB8QEZthMNrKAShS1bqaXEzI5/U6Ma91gq+P1Ra
MKK0ZSko2KmFI5qD7ecr3C7Xq/Y28pOz2YYDKUYkqQdW8uqGRZDxM6a2/Tm1
N/8Z4Di+TOlKBkOg3WZ0awANlQdCKn3dWOu6Op3o+/YRajOzzlGw+wi6KAtn
HChilMH6Av8v+yKFqydYUR8T1XBtKlft52xx+qAxznwoeIDC23FwgkmVjG86
Iqdt1MYTADlSXdSUJNX962WkD6hXStwOdJXBqqmTa/ayBA93etYV4IceDBUC
SLw9MhNWpCDGk/TKg9VSgEl7NTC40K88XLirfqWSBv7bt3Pvug2pkviCnzd3
2BzIN5lA0Eg7kL45Jw2Jxqm9j8OOAijPUwdy/A8waehzzQeF+KqlvJRQMs/k
GjuqL5PiCtjxfYHVb1oodawFqG1cKsNjYFAUFABUfhkbjNQcs+s+iJBl/sNG
y7CJr2zCllTgKJWWaphHUl/EMsElbL2pAFgHf/1e66s11OWJmKplovpfr9RS
3T+j37sUvMjLwRi3ukvuHEXFMRAjaH9Ry/V/SsuMO9Y4HGTQfJ227yyGxgR6
s5TzSK/BIADoo2gfiuI32QqngwFYFQJ6OZsxd0WfLUL5S8a2Gg1txPivoCix
cXfWQ+/J5Gr05ZAvCTLWK+2v/jHWSFpYCjQ26l7V2/HZGjbrSUIYgI1+XYc4
AXFjXOQVx/FkYNHe8A0sAlCbo8kgjSUSMN5EBtNcAfvoWOd0iywVH6/B89qe
w7C/YLXGDrR+GiKHXv1EQCnVTBj+IU5e6zzgO8J5rG+D5dtA62oscU4AiFdM
PwHFZPeidc8A5pdjcY2NIrFbBNzFCjS0E27f5m4Ycz/BMFvSsXvbP/jbNlt4
ILt12AcN4U1bf1jfx/k34CqPEvdqqMbIJ58favlckKGIzJrCd+n9xB6BM5dj
hR0ya28XuhIikULamKP7JZl03JrAk4Nfbu4uCLeblxyG7v0o2vImn/TSe1VY
Kk7V+ZtVOyJf8DyCbxoXn0L6uJ6Yhe0WgHO4Ql4hYKp7LjgdWU/aOSOShLGL
JrQm94P0OcekXKi3FG1zGJNCimxQ+JvBWeyflhcowHU/VGjr+RYHRc7vM6Nq
US8I85LE+s85mvUKWUqEs87N5xVc66VwRItppwMilo7d4EcRYJi4lMh5qPVC
QGMELuAcwYswgmbnea6yGXRRcj431qOSs4ztuX0f3olZgn/HimDXr9texcpD
C3x6kk3Ka8+9CVsO5bIXZmx6N+WfXyMIxfDIJ3/70ym8pFUCePtoHg2Hg/Pa
ReerF/Ypm2DquPZjSP3Oc5nptBHk7Lu/Ye5DaUt7TGNzE9+b+H9yTLRFye7e
Cqp9V+fzr4ZbJ30r4Qj39lAUQQ9HLPwNhkmaz9RxGFdYIdYHkXmgrZnZRCwv
ILagQ5i9pB0/ttWAqe2OoyBgBPiyBLNKnmIQ++LvdP8mMvfiM+iCNk1BdITy
rEAXApN/0l0ZSr3c9k7ASxQrbiF0gPH88my9uM7fAyEObJmmVpe+KMZ5al4K
mhbDkVcRdhMrpo3Q1lwuQ8ERgUrQuj0YOFpza6Petx6QWWp7K1MKfCXeywix
TRNdF5UauHQ+4lZLwu+5upaum0LdLE+XAMeTjxqxh1OiJ9vqcHn9ARD9od+j
X6p4VqbAcdZvI7/aXhD1rDCumTbbzAhPDBbHMIZwIa2GARCZ1rDyNVsb3ugm
A9B6CcG465RcE4xVokZ72GDnKehHzu10IwiiNrwvihhMNZA2qTRtbNeJsBox
JBkpxkymsG3/bNXCeW1/uGge7vJs72n6kvPCAQ+3scqbZm+yswKkImVDla5u
lJVrkv3XPwDJ1BRRBsHsXV5mjO4CJo7/oh8aRyn/7VZK+hf5D/wjZDkKn/13
IMJq/vP1wtwWtdiA6fzZkVOEq8iERwqs3tVBrpnZdCYiEpsbhdf0V8r12iPa
fvMhyRx0V7lNQ46pKNW5vdX3Bvl5kVAPect7fQkIb335+xGyR8LqJuqLxXr5
Occ0w198fl1xJTQ3sNmgHEtyRuY6s9FWdBS9M3ggwPiZTJzxutHwDJ5aVB+7
g8PYxH0/QmH/pPe1FqT9SRPUAihvEL2rwIAlKPIsUboip50oxjO01nvm8Acm
tzU4yx8HiXjjmKfxbjntA7OxxJAtgTUJ2xQ8kRXSEPEyIHPtrNLy61png+jh
OBzEAV2j5H0uXsIK00b0saYBqSGS/FP+3uzKow1hJxZG4XUv5Ahxeldd341u
WFJV1hpGqkkGsxV8AJjY4MwSeByyv2/lCHcXwltUmE+DpB1MZCdtUA7cX8xv
T9TLt/u1g3fHfm5VRhiTXcuGDuVc7Q2q7TpW8n0G+44gUlr09Uxl2ZV2iLoe
hZRSgfphKYPcqOmyzzn0ezO+rJQSJNlgrPuht7VbLat30bRgdpeeHVjKCxFp
CbyoKA/xU7jZBnKKuUpxodNVP/oSX4uwkqnAy1y9To8MTb1qfB0R4mGCKOPM
C2kpTJ6Gf7/KyZo43Z6Rw1gx/JefBBcvvKj69bBONMf7m+HviU0aaag1kZkn
bfAqLwWp+TNGdRmnj3PnorR6B3x4cMAPejpp4zXsbVMc+GrrdzfeHocsxGlh
IF0xxxz3HkbTe98UF4Sut9FTLlG1h8UrAth9aqI89iatTlqQ2e1o6ucdHs2J
XA9dE13QN047vibPN16+eOlWpiAXqFxwRCNt841rA3XH7PemLnVsO373F1Ax
0qGMihenwK4rL9PeEV9BWrR5GzUuwz9aPnuvMxTWyXfU3iYy4aX1DqJ82MPt
j4PZOiSfSG2uz4vwGpOAklhXCxcEYLpLYUy+siXS31wIan3+s2lcR0cWoDZm
nmxyirQI7x/mPwpwuNGWdtN+zVzRO5DdRDjtj8AqN6hamVeUktyf3uwJM77z
DNMuxFChK4WHDcC1s8lKWbNs22uwXOrzJ9zvSXw0Q8S85M4oxp/tOMjJ0XET
C6toqXEqM31CKOi5161DoQegoO7XwQCvwpGCmDoVDmaGwpmcxL6es7DSsLsi
Hs32HO1XA0pr0vHFO4A/YypEY1MAAhldLhR/eboA+eRdCUHpJ9o7yl/PJftB
j55OCGj5zuPBJW9oLZhm7CCHVQJVFFKtPohwj5Rwkjc/SEJwsD/lFs+ivORf
Gw+G4xZZ5Ufip1v+MEAMHT5+G88l1tN0o/PNwEAsAh6NAkDm5yCm8cvTrnfe
6qWPIs7jOFYSQSBX+j6wrdLsu87ErKa5U3QIjpH+SZZkmJTNukHYXROazCaA
BArXZUp6G414ACO+TZDXjB/6R2hm1GR1v9TPSpM6L9qQ4VVMp/y3O2lkbslZ
L7YI4kGbwfr4K/jVyt10hfUqK278N6L9yRKDGfWOpsYOgvZ0QKBDv6eKOyP8
DqUhwUjQXWgxQNW9msijcUTF58tLdF7z7mgr8GBf/5aliSz/SOYIUAfoFTLb
Ye/A+XeRtxr61d5nEBgYcAuyefWjiR3os/ekWRtCKDoql+fF002TXDDWLvIt
8CLTGCFt2hRn5dDkpanHAbXLd4oHXwjYi/XPJsAtq7KO1ujraF2tuvR6n9v8
yBaVmFjD1/akDgwCyneDQFpFXvULQJrueVf/ix7ZfldmCTy0EmTdxt9EGez5
hQysyKTHqX9JcGfNwHgpad5hmDplOsw5aTMYiH1fkVWrdKMX28ejOQjsSgm7
2X+SRE7FmljPBuR/VSSEyMPlO3zjdlkGGxlRGG4EL1SB4bGYauTkJmgTNqCg
kEnC6aM6RJYTZMeiFJb/sNZkFIZ+eYwThKGFPC4YB38j+XOOC4exnehHcmTa
/WGnINP8qocDjPV+AemY4vowHFWRhQdN6f1h7CMqaoddAT+kiF4x45nWHir4
j4s3+ZYOSCuqAelcsegN0SA28b61kZm8M3YMmtH2godnejBOvMMZBTNs6Q4m
YGR1skI3sPxBS5cpas83aao4DknfUp2oM2N6O1InZOLVPSvqYcqpWE84a4R0
IfijSq04zTIl6gHTpQf1HSkSPjoaSgdZEbJv6paAt2ENZFze1xziqC/C4qtg
YePjB3szIfGJHFA5oktVGd+K2UgsdyJweuuZunL44RNAGdR9PWrfXj6ldzST
x+1zTQMAIY8B2C/gL3p87d0sY80zDYMeNfr0jSEoTCgyt6HwhPS6kZzSHL42
R1v75M5iBktzwkOHd/Ci+3WTvYG4SBO+r37XaOprcV+iULt7FzUUBicb+7q4
dx+n1ATHzIKX7AHEV1FvEWyVXT9g1cLg9+Pal9VKefg5bmZ3ZniO05Toe2Co
oxc18hXPRUWUaUen9msXglFW0jVwwhbCza4zhEMuwTtCBvzMEDrppLFvvmoP
gMCoksM4Y/96ms1Au4Q6vDnKYtSINwiHtK3gFjPq7/BZwHd6yWeMythVT643
53QrTnQNV+lORiWdI/02RURrZRHy6MoXS/eyFJ3NQ4Kl8cJfNj5Zveb65hXY
jivxjNG1oY4GXUCd4kfCJW/GH/gWAZ4hnO0mPYwx11GihcqU7/mVgRwQ0xPR
FduYOS3Nom0LKnb3aewainQIw32sRI/C5fpaqHh/Jrjg0PeuzoEqefzVzUxK
OO3Ijv2gcpzodFFidX00J4rP2EdZARyi9C4/VrYomh5LpjeF7LhxaWuMJt0k
3ZBFfGWTqKezsAy9XGVsUS5BosyMAqT60d+CSr1FcyBv4M780b7vFyNTsEgn
DpRvOJDO3oBJaN9m5ffrjh4NUJ/LFWkCC6iB6KqIl3Q+TWU6D/MehOvcvZT9
Q2sxFLg2y3AwdCV5k8iHLnk1aX14IcQpUCcgLIeCJh05Fk3eMSNkj05WqyXn
6UxFUYheoV7XR8x1k6YiFDLAL11JZraSJbTDxzwJjwD+Jj+qPZYV+ADFUt6w
mL3WnbQA6rUapk8J7lnp7+0CRemjBrwY8P/bM2N6kUUBndxeIQPI32yQQFum
zsV6gVyEtQcasMrGOHq0nycEZnpea4G/Q5SG4O6lAz03HNCLhpL0aCshFtdo
DVfzDKQ2EEQZMd7TjG+3MBIH2jHe9n/gHuQI6NujSRrGMQcvxuznTWO+CdkX
hDknG+28tC/fsflT9fGbmnWdi/wPuCoeg7cMYRf+fyqXnf3aGtYjKn/9so7T
lsh4Zw8odJ8gF2yA5GsJd7xPwfnafx7P/d2LdmnNbZsE3hOhpB9/vaZjopR7
v5wAVO4MN5+sX/OAN2bF62oxEuesY4lBFSxUAhL3CmdoaLD0W4UbERigo1iT
jtj8/fp1UPZERR1NlGA/P19h7J3WHLBsA5qBlGuwuh5SGHxurKt5KDGnnvWD
O9/DJPJvejoM6GraxUYuHWeSCPcLNssISwNK0+nv2fuW09CO38jx74Ac446P
XbEKMuBGRHh5IeCyI+yyXAF1qQXwZTVbdoNV0XRYWRWrVgk75ANe1NpksMoQ
f768bNIiG+OXAmLglE5NCXEVv7w6efO8o7ARZQFrLb41RZUPl26pcKR0nyea
qb70k+IwSkufvSwbHMXjzry8ky+uJx2JQBKilFrP32KVWnHXylElWflDSVz+
CfNHRpL+Eq+EsVLkwpnR7qug0wAbHgjO7DNPcCJbZU6DXteSP+lSkG1UxKQ3
qNau+NMde1bJMQccnfZkdwapVLv1nz9rI9UdLbUxxDNLBcwM9V7tmq5lcDJz
gputWVqUo0IouBaHpwtKzbZp1EkNJYIe7ejthO60vlcCaLMlw7h5PelVOYOu
QLJPe7pjfpXq3bcw69ESwHY/GEgEhoYLUZq9JgVliWY9j0eqic7xj6DecfLf
rmNfoBFFqHoWmAduwYgD9DfzDAAM6u7X9xKM0EYYpeVVf0PCgTsuanrNPp1X
t1UFt4qYRwxm1gyz4T3A+QR8vjsdXIPftpatJT9paEpnzPutiOAtYs4VoA6P
XOWoklZ+nHyMdg1/5CHV8a8DoFmGcW3jcHg9Sw/7beU8S6ISCgRfOhJsVdMC
PsQ/eylHOjLgOEJ46e7Tcy3yk5XFyQ3NOoTi/ueYhv+rq1N5OvWHhZsSQ6YF
RSowgV1HPaTHwt5t+eAfJNTreNzfwEUAzxGgUUpAIF3Ui74aBhY4SrQAOM/a
BVKxxXyK8QnZ4L4Gbd5PVbwGsRJq7V7aED0WVFojFJf/Z+elsgebnihJ6YDQ
pu1wLVQBYaqDug2B88GKq5VTlRGRP6ry70uT983KiUH86Vw/zNlW9VDKRwXF
zH+xPFNDCQ7IRPfd+Hp6xQX0J8S6gChnEOuMVqvR28wNk/0V6tggO4oNz2ab
AoH7JS7tc2mgSQ3EIrtuFq1luXYb3Ra9Qbdwd8gI7fr/hdpQiyUB8XK86MyC
hqeN0HBk+0SlS9vWeVLjeQLusLVlvf3Jxwd9xpf5roVfS9HL1ZjiYn71FkHz
JWoWDZAvLb2cW9fzexmlA+4juxfHJJxfWtb7aTn3jV/Mr+z4pWz51bE1qmCJ
sTwe42iwbTTVag5gH5H9wLykPfAJiGzsbdGMNG3JMgvzSJdMZbAJbnwfa9mt
/y/t/3iQtWTKWJy8ZLVI4Z4fMOrnuYmSGVac2marvHDGqSqhwC3gpV3fO0kJ
DWc4UFZfJB7caUeSWtEcpC0hi96Q2c1gYgVeGysXJjc08kN8UUMv9RlNkQP0
ZTEjwlC7sClqErrbfCCo1GPSDfMzHkgE3KC8ujjbj1xuXL24iB9mbnal+Ao/
s9foAkWE7M+31/EDxQt9sSgh87QVxNYSBawTboPvgjG9YaoYOCg+q39/9git
Kv7/Dmzb3YAB4gcfrW0eKyyvy3HNkLy6ymMEkrO48/94ThV9v8pmrCRUbiAx
OOEz0laGFLhzuStwt/SyeXbAPQSdnag3EjA0KrTT0TeKUwUcJAxznSOMkslT
APwjhXy5Rs9XFqkRxdZ321WzJ1cX5o1XAbEpidwB8uxGeRf57m7GAu6MLAo4
gGgqRT9cYLUEhqBX4scjaZQsMhZYF5D8k/Urtk81XdgOTZEAcBAemi+hhNYw
qmFQSPPQAkmfK/9udiJN4Y0fP4S8PbtIcy9VwjBBqMlzW0p3DOsvsNjBCIxf
mWtxSDDjuSx2K1qaWVYDxQ0+g7O+WIsfSheYnrrG9ihRzRXKE/laCrEGD0/5
GO1cf3QoNbVmRtoqm6Bv3y4NMzW7DEDDm1ch+d5YQl/JPA1a3UIq7lLkvY2s
N2ARlek4S7Gr4HO3zGrz+8IuGr+9ksyzVwYIg0uFuTheh3z0zha1Mh9TRPZK
0jbZRLROHOvR2sEoCBifjnc67rYUka863azl9XZsp/CmPB2YoFDJoZM26TPn
e0aHTB1X9prApOyT+8Ssemr9W3woUB1IVeUSJ3BarC4+8J4V+w/7uFQxryo3
8k9d4c0HWL+dKqcoiExjJh/HiHi4634YvIAY5NIVDcmgCBcE/YXQvWsW0xNk
itWtuLrXenl1BlZwREj5Fmpn0UPE5A09hHi90GpCLkM3VC0+TNejtivdLsSs
qOhRXF0/zWj3sihwAq86rQGvr6mKzSpLiiek5k8775w/WCb2Az8a/2MEKatN
CTvX9c5P1C579qZYczX+rfmCy7DpIflZLNK9jyjkhZMJccfQ3qVXG46Vi41V
IbiGZCRxGT7lT6CfX7omzDt4AJVH3eC3aOhD7GtIOWEA8c7UloXCvw8WNIyO
5bbJKPw9UWas2fcZcLQnP/rjh6q5t0NvhsX87vQ32USDaJKJhZJQp6fbElj9
BJF+/yeT0mnsmv6X9yjWLlgc5AU9tQQvptIj5+uY+mUfWBJfZtyW3Fr5HofS
u+vg57N01N7LhZ2o5tE9oMWU1t7ep0bfuJq8h208zu835ld6A7CBntWtkY2R
TciYn9vXxrm784VNtImGOEwKhncXzJoqnCPLm05ekYrR6kPA3HDsEYlN0MJi
gn0mtrvXTbS9vOG/DwCr+E6Ov2CUDdxJcDqI75DOL9bCwAHfkRIheaDhN7/q
s9SF4kUywe3SNnwlsQ5d9TxfDW2Isg/RZlGIwZ8QCX7lGFAivrR7Cxw57ETL
4GC4m7XKUD4TZjD8gI4ZAwE3HalJfXMzh9NPuDD67ExgpTHFdTsv6lE2Wgvz
sCk/4a7DWyWzdxe4619Jw/1QUSk8GLeXnTj4afIM77tRs219f3V+cgq3g1fI
yu6GdrfqEKYuK14opWVSL54DpurJ/i+viCiZzMOEMUlqv9LBX8qJDwsBNE/5
FmeukNdDsyvM0DVOBraDwAoS8sraqc9U6352A3Ch9XHdui4liHB4iPNPcN/x
EhxwxXKtfs3Y0FZpdYVzNPEYZW4LymvH40AngS7S5T9VzOv/Y4nxpx2QYa/n
mRfMVy+2D4fm7kO5VUvoXrdwWdhI/EkJqihVV+MsCLkjKZCWIMPGeOuM8G30
KDNyUPno8xJxSfSE10fFkr8WUaSyih+VYEM8sWppGgWk4sxIzVuFeoZYCalP
VLumhh8e+RD8rvuiNX9AglRQg8utPDv1yv2UI1LZ9m6Duy1Ez/l8nQLw2cqZ
i2nlUpTkaO3HtzPZSheZ9KMlHRTs351B/odGnYJio8sC6apbMKuvoZ62rrG6
bw29OFX8pYyKzY3Rk+2Biro4ritusvIR3/5V38zYZUGLaYc4+KMl98YJMoyW
j+ZRt9cGxtvy/PLpP0PsoPf3KQx/q6BBI6lKK/l1AWx9xAkGQ1A310R4+XsW
3M/tSUjwgvtz8PexMQTP45pHo6nYt3BqYSE7eJJK2ZivNMfZgkQ2Qc6Awc7K
IPkVAatA0Hqvyqys3OH8XCQ4cieXRX3sqcPCUWyG7jbILr1b5sdUcr9Nh1Z7
hzyFESwXgLmbj5FkPiDr4G4TMJZSnIgRG5g4GAsOYlP/caGJc/cpVCz5NC3Y
PRDiluo5fop+Fe/IBRX9q17HszGTj3gy9z+gBpVSmny3JmQAJdpj63cF6nUy
MyTl/k7UdNwvSJ9oApOcMKy0OtqnCJxCm6wWc/G7v/3Pf2LO8a0ljeCu4lDw
qw9CJ19Wd2zaKYDiCg+eZCl31kvyLAQXokweT57lV+BVM7toicUxb0XHa3l+
rZ0eMCFkV3SKhPtB5iwxJJEOm+J+pFBvkjOon6rZgd5E6Ciw8k9zMhEROenX
cEmueevc5f3QJ8/pxJG7xUp/uMFNeym92nCqZpIaqWhLhPAl6yuKloXXBCN9
50+oAf2pnwtGHwslfhXneLHhL7JBsj+3v36r2Rt+k+Ca2igNqrRVvwi+QwVo
xk3LC1+P70/kBjEPL6o3xdnJ8wMcHZEO+jIlbM8EzpqxTHZlmdnhz8UiuBEW
K11L75FeXfiV/glP1edHAuDwTzFmpzlFjRHy+8e6C968SALnURSKb5DGNC44
x17I6quqdlAdaAtxMDC/fG/3l06Avv1R162FsErx7eRGmL/4AGXKkO0bC8QQ
TLD4T0cr5cdoD5IKoaGgRC+vEjaMCKRPOm03yyZCSH1X42RTx7tfGoyCXi34
9DCHH7F+xJMBlsnvkDu0dAyXic3uwE1Iix9d7CfMxYmMwCC9M1wS/EG4TX6u
XrCe4kCAJCjh2HP46mfsNiMzgjTmcHzVy2vJXO40SHOPj2zam5/dE60tVTAS
wCkXQLx0NQ6OHu+XUotPpE618gjO1pCMRmgn9oXiW7AJ5feNnfOB34KxWpAl
mCV8kreWhpqzgKKDjP7psrILfYRQW2F7xlC1Ml/pGtDvXmWZFhPl4UUxRS8P
gyq4EGcx06eIF+EVqD6lMtfPddZZlBs6Oen/XvFAjqnahHCzEZorgi2puxW5
CXq3e5oAyd7RISjR8j9f6dx6ddoZZXAPFB61Sl+I1PKBvrm5tNnoQUqH5DzM
oi8DbMpgbS0Uq0APGiAgxk3V/LrLFJvLViO/6+fB+ppvw6Fq0NC+wnvKKsKI
puGYiXww6ahb4Kf30yGBbe6EDUqeWp+QDVwTMYJ8/74E7R3oQPAsQwQ5HflQ
cGdkHzQPp/UWV15zPDcAYU6spNYUs+4r7nBWU8fRanK1SnbaZYCBp1FSGzUE
1Xa7Ge2F/TUPgdvqfRn1x5cVCTPvTid2euqXRfsmNgwdEdMUn3Ed7OI6+R96
C2oytdFzFGmhZ7lNed1TXTXebd4Uvbl7cywWuFRfRM5r5deSbQr6seD7+SHi
coH/h/pdkXub/fWsLUecLdjB2CzR6R7pUwb5KHltGQP6tP3J+xgjPqIGaT50
568mtG55wFImqVYvVQGuG1u4g21rkEle764Fc5KlC3Po9AdYxYkY0sstkEgV
jDw0CSq9EX3S7mmYrgHvaaELBgeUsFBGFqZ/GIpzW66UgPWxEsrTaaSKNW6c
LnIdTSoESlZS5XDxKD7yO9+gUdR2Con5dAchdpXE4RunbUR+RSki6dBkto/3
mR1IzFARGvikXl0QRH4gECTgo3gTbYRtr56z9Unsb1EX17IxYBTKXkLZm9RD
tH2n7K1j0n5OgGPOTrI1MaiLTn4m60E95SubIs1KuTdiQy31wfK9gyzbCPP1
Y+ia5BNgK6Q2olRt4kCgl2/ooj09lNBFlEUft82nWu7KV70CAc4vKX+zQzWz
lS7NmtkRAiHYmligv5MC3eToI9Zxpy3eB7v327c1q0jZPd/6SnJjafpt6h/o
4mMdU81vATDh7rlgafjddYKBu/qimvN7d6/2veGcXWhtGQPW5uDC8M5iJFR+
Xx34g88eGw7xoVrCzUBhRf7ED42xLpQsH3W/GTOHDlsjtxEJvz0kVTWVaVIY
1nMXtyygCDWOCD2dO8qizgttVtm+CjfHFhrjMHjtk4oO2cJk90/qhN9/4+Pu
t+U74SS/Axo2TnOgGVgJ6HkivcM8vUUpT5R02COSUSrPn+aYxm3BbwlO8ML8
ky45AUNe6tY/Ndvqev1m7SPNhZre5hx7yolbFr9vqIDtsyxxNEPnKL59UWe7
lgfnabm/wOdQ5w4HQowfLvJHJ6KTbvWejavP3oBI4L4Mako/ES90g6M8lGDQ
9WEe7YwMSzGLErW3NC1FCfqP9scOdR36w85tAriifHf/yRdjqz8S5FYRfkWO
jnxXFb1yEpCmbEZbKWid7AyGJ2BafHWK8lXEvRqlapiqguSlaUCjss0LVpfW
sxgOpd+ZCH1HoXiworrJ1eqStbkZsCSxISsNvGVkb+P/Vqow514mzbAslswx
ShLK+NueWETSNrNIYiOC6ENQp8d7tYrMpQi+u/rSxrnq52wder8x+JuyST7c
DnbzmwI6hiYs35fRbL7w/6TCY9uxb74Vz+5w+PJ4jpM/rJqK64XNB3qpQGAd
dmRZa6SyiY1br9igxq4uoW3cfFAaFDYfargT/msAsH7S5jT/Mh56IiWFUIPT
z/K1+UM/DYda7RB8QmsGvkFK2/CD1ImknCe+/d1PMmB1z0KkZk6C0F8190AU
q4z0a7XybtY4jafJ10z2LJhfyAhTAlBbCHLzfqY9nBjZQCKM5Ait/NL1wLTu
/O68tIW/OmPI/JLrNzcjdu7/n4nN+8kxTOTbaYXH3vE8F5JrSTodPByQ5sua
h+17TGajXpo3w/hO6UXvYHAuS5aMDM4geSLtWrYf492AOn7N+X53I1OlueAE
ADd70pzUilheVe2ww2+tHRJkSqQ9HZppibI/p4ser67BovEgK+WXPcRSIlJ5
0FD5uFsQW1Rlswqy2lcczL9iJiaplJGnIwX12LENhEM2A+wy7LS4boS+5c1Y
AIzEfr2pFT4jSb0lW4IlX0Jy+3Bk9A30+upizNgoYv5THnnFv8L8o255DdNE
yuonYkiVji6LWwW2w34ohjJSAQfYfTGGpzhpdu/vkfJD1g8D8kWGQb6R0Pzm
+amxYRv0Z+J+N+YBGdLNRH2HPAnOgSwDgfFFbmurFndLMokX6ucfuH7G2vk8
H2s2AJVLuPPeekwrvtLv4RVMRQr6u4VkRRksyllgKP+I7CeevbikgyS4KK0O
557qU06ZSzZNVBNGSfhvQQQoddzd1pU6O4SkiMbf5gGf8Yyj1Bqlp1BuIHHm
MljlkEp5xCOYrjzgl+IajdHNoD6dlIzHluIhLydiY3/nDnFiYVSLqAJ3tAH1
BxaEHhMWjNNLX5jj9MAR5RfDvnnAJAgGCR4L3Y+oYAURKApQTENZ2IE4igUl
281SnoM/3rB+A9Zav3H56D+mNYm9Tx+aI4/g7/0cCgksCFLsyOr4BOerlTXN
KmMz2vIMiZBKn3tJWdvQb4Lg8qFxPc5gqj4XRTRGOlysrQQKyaRUSXMOh8cf
TXiuO30YGOccyvF0VmOCEkAaQlh7AmtamFEjoH+y7oIh/fGuPBwt9RtnMzmV
6qdzWzkfsqBxl42BgzpBrW4Q/dR34v+w5bfAB6QQd6ni+5rdE7+Rd5OSgRE9
f+KvKbtsdLRx71GNae8Q+Wj2Lhs++j5o9TiQ72IVWViBCeX6cEwyriRcg7sN
7Ggihn1U+qTpsfESri4ah3QVeQenpTCQKK4h510Ug+K2fQ2LjGycqbg24jT+
SUTAoCaR1wlckvaJqlSW8ZMlTMtHdJf4QfeZucCYuhS0yVvCWsWkBPnhqhd2
rOjhWrVeTVcJ4S629dJUb4pT41dl5aoF/1T13Uyj/NkByaloDmRhRcldOgqW
Le6q1TP9bMhZH6oRpf1Yd7fmar1DpXN9UGYblRZjuwfyXbE+sFjZny78gwK0
fY0ODArHtsBDywuT4mbdMV56F7aacYdEtN6qrBdlIlCz7NRF90ZheSjGVByn
kYBDw5dUxONAyLEROSZ54n9Cy/Zjt0thGBNROOOUaStQ2KP2sE4lSUI+kjQn
AfTq2NXULD5Nyy/ZFOp2U653VTmdq3+uIVaujanocLDOE+ABY0zciJEyVP9l
7yHsDYFRABu/x+qY1ekqKLJDGYP8crsdnQNdc++xvW/7yufjm+6J6h95yCFv
VwDklayIALiq/PIwRWpk5m1qXCyPIddQEMMqWCCpObGV2X9EaXSPjZueK0Ow
PQmyMtStNP4f/S6sjb5WV8+wjzty1xDT9Z7DVpMk5RlelzcuthFosXIeN+m5
12IBA7/J1BjCXdPI/HHJN4KvhQKahbKk4XVATbKzD5jpAHNdVZyH8rbP/X/7
o4/ZFr6FNc6Ne+ZQLBD7fvPFr3cLEuLyhFhtUGslhZWFMH0Qd7r9gYsw1PNE
oRf/0SsPbOUudKA8eqMphv4vtuyp7PLHsEpirEB650jIscZ8yMdvfftEmUma
ySoFsCQF80hBZlsm33lYvF484pu948Tn5M3cjA4q2jgSoVmeUA+p0SzJItbk
pat8ec/wKGKkMMgRXI4GANTYnQemwXGBDvHnj6CmZVOO/E1jWI9c/scmb2Rc
Sva8IVOfBGkzOLXjOmyWLVwZKg7RAzho/MHXgaUKhzoLgqy/hQR2+Q3w/xJB
U3s2nlBMnGa4uIMqUXsBAOePBYWwfrXcJx2N8ZuTqFxtpvMyRtfAtNOM+ojT
RlsG6J8o+xYXtxDujHxX3MfbxR+jK1fUAvDjeZ77zKmJbPGGlcIdY0RulX86
PqszL2srAOVqbvK5uzUNQ+JlWXq9+gK6m3ZpcySSFL1rfqug8JELJFcAAvx7
nxpPjDC5nPOEp0NaUMrUZL38S2ebWce3st2mTnxx7gjeShqUd9k1fOB4jmyu
A4QbSL6rT0zgU2uR3pVbON3t90gTHjt3jvUSw/HcqoOe+aEh7xtZ99h3GME5
uvee89a5qMx036I418hiLFqrgUOib4pddzXuubzOEQ/Y9FEk/aXzxkqj1Gwo
PIVjD2fxsL7tyX1W4jF8CaJ8WEc0TQKJuoVnlSdnfvG63IAeH5ybGe+nfl0i
j0IyLMEzR90cg1NXkfVh4SBBjSJqztQ0MidS7kjmAjAcGAjtHTSAeYtiyvK+
7w42r5ZZn+3ZRdh94ooxrwpqrSa3fEwyCFX6jH9BYJnvhDnEnOxVF8Gmif0l
ET96dZfY//PR0JywigGbBrfJC2iRfLWU8nMqLURE7OASBOAI0xbbt/X8aeTK
1kXqihcN8lP6VlEuIIikEEdjqH8w/MxQg8SkVKZx0kE3mWCa7JTE9awm1eCQ
QW02CtSIESJ3hxi9FLjNxo09xSUJRvF8KA/qRrxQOqSbcLg9R6+wuk9oUHI5
Zrb0msazd6lS11/HwcxuMgmuYl1l6WtlrzAA+PO74Naf2g1DdheBq94a5ksh
qPQGKqRPmv+PP/9l4RVBJ92e1BtJIURQCtIj0VBbhJoIqEz4prgjGTGZQUcO
oLWQkDOHZm3PREqJ7WHwmalfkObeWluU+lBYJkKBrfPVoFgJ9dzBW8Wlywbc
WRI9bj4XQ0h88DH2LyS3SX2Bfa/b3t56XiTJDCfuMjgZqKhFeySQ7sfMtJh/
1+w6dwvwsuBQRlC9bq5EbQqQyDj2Vv3lOAl89SmsKnvPQEhhGEcMRJ4BF/ml
t0GzbtqgqJ676Rdd14La+2EpsuiPTamFbZQHn4z/i5aLj831e0OWnHFK225F
D50dX9r4Omt7a2cqWKuCGUsQw4J+HzZYChsbEt6ZgRAhEvsnpXYVKToZWE6U
7eL+alsYySMUS7zCyLzvNTxSE1Sw9m67E4BroyVqRQlsZeae80XO+X76iOCM
0oYLqdUTJXUhCx3gvIwz9CYNp36fmsNnHMLaxhL7YQ3uBjpgBqYUo4fgVkYn
Gch9K5iPps+/swd9T/88ES0SJDYRGk/jc2tqCYuUoOKvoegkiElrq7Gi2Frn
VcW074425BZ0gFO4YxjAlZ7yz5sMGFThj26YwnZc7wYiP+rK42gra4ewabJB
MzxHG5GE6Sbxym7wyO6XMsxN/duvJtF47pKDxW+6KeGP8f6hw5zrOEAMSdAU
yxxcj+AIVcjDn+y1x2ZQMG92ev3A8oK1dMvjmJRGjfiWWMJAnhsc2mmoGOmI
MmFHsn99TRa6i5Q9xfU0rurPJ5xjUD406n8Eqt/Hzn0DA+Im6hedm+Ch134Z
BmE0ibxxpc42nMW43vJVz5C+Y2SxUmqIno1AeAjXKVouVbonhwv2L0KIL2pY
7/FaIdrKNlpoiTp0PNIzv9oUb8n81lpIQWIpuwojuVQCR3y3pB3p5x8mNKxO
mC+IVUtFrQCeh6K5PW6Qmkh9NNE1qwXuZXLmUk52BZ5w1zKIMiZTlraT+WZk
AlmFvRmEPJyal7jTjkY1mlSH/bLiqECV+Kvc8hB7p7n4dPCR4dq7GoABoQo5
x9v8G45Y1A0XcaeYmenra84tsSu1WK5AbxsB8p66hYPwmhDM6CxksbyozMiW
xub++RI7dkGTnuuVkX8FI50ya3KheDFc8QHDeBX8g4Uj9aj/CXIRydDGkY5L
Hpv5YB+sqM4H7/4jBpeL1S03e2Rh4jm0jze5Jha3DOAkiU6NtDiSdF2tM79/
oXrmOACzVEIs3bQEGwFJAsPmTh6TFZuciDSN/huc2npPt4z58myW/L6XFgYc
AYqDv73mi6WI9zxR60eoH/UsYeTpEYk7QeiSJp4Aej3aIwji3TWcQfFTolMy
eu6/1/dlH/roYelwjwO5AlyGSdwcFLbLi6Lf/8rbzBXZUJE9Ww9EKFHzCgCC
M9e5ZLqhh8v7kMlkV+yfCKfQgcC8CDGCGB36XetU3LFVqFOdbjybm6FZ3d01
zN9igbc+B8m5htAiHB2FbZy34uYVUnXWnd/0klf06NHmZby9LIwSaTnL5RqJ
M7HS++iRfLktbFPIquJnezKNsLgdse7JvAFWaHviQ1kM7LByRqdBTY4rCEuA
3hOKRDMwvNNumOqCx1ANEVTAi9Pq2WBOP52ul1LBfYuzA6sJW/VJKdxYW9b+
QiRhHD5Hlz+OGVUjJauoqIWjRndu2Ohfju45S0FbwvaTe2I6iNS933qQyPg4
gq9K0c0hCULtSEQx+jiwnvSBnOtr1JkEel1lzP02hmrpKED2hj99rVgM3+8M
mTuaopdkZGan2nOu7YLmEku13yj4amIq55iD/dkRXFQp62GVHBDG+XB0TcTY
2qCgPMYa8nXHeH0GXLrdNiGcL9fa6NZ3wvGd52Rd0NEOmmy6hszhAS+vPWE6
XYNFIvyp7FDtbRz6oEoq+xoWN7VV1m+35UUGmOpKt4ZDQhsFkPPn2T6XkOeY
yC4mQkF9flrV0WBlnwmC4FPeWZY7ywMVWP8mAvfNlbQuyIZ0fK9kbHCQ35Gx
MuG3chry1wUC7GfbdmoofTV+MMpOW74FsBtk5uOAQPXnd9zjCMZacKw0836B
bhNVsUxJ4Sn7p6UOgndJTobJ4e4cLvJkL7fwzkPbY/TOnNnCD/KLsap4oZW2
2tq3ME45acxmAhUZrAW73yhi/EiCXTR535HvBXAG93YyVixkoaFkvN57BxzF
7FBoT3gRIKIghM97Ui5KFeirzpchB/i0A09LA6PoxRerIYORpb1bYABsezQb
l8jcEwEq3HqdUEe2pPD/97RdOAnVDlznejsAbczXnpuM3mrAvJaGroa9Agvx
8mn3UJygF5FWPPRFVJMtbG5TjS1ANZyI9cGMIcAU0M5AtynyEhHVGH8+0gv1
1JLV0axeUvVlIDKU3KJ5MbiR02lYcXat1yrnWMJgqDoru2Wv9JssJcmh3qQx
tx+RsQjTAAudo/AuRPtr6fajZgsS4tXcDM7K+Cbo0NS7QdMk/0+QqB+hiKgA
SvMZfbLGSgMT29qsozcyM48xGNyJuQNYcNaiCjQQ8LAvnlowIHgy9kVqhO/I
ZXW86S2y2GMDjKsHT9EKXrlB71GUH6wWPi8A0reyTzbkmv4Whm+R4fGqlW3D
7z0N8o1bBFfwR0XLQbedD0553h+F4pP92gGixlXKkSTjvZkkvSRhfq07/0Kx
VhYujwgR0NprXsj6rSlpqNxcTiF/62wehOs2jHwobqiXjVHAy3eNbnQRA5SL
ioULli70dy1yF2rQgOkFQjpg7/+YyjJ6VbG5FvvD+1Rntl7EzJE9tmsKzQTO
pcPWehEta8cCBXA63gzYMiElKlA3no1sqHpIRYfZENn1SAca0Uz/sue2Egg6
VN8sVTESEtGJ9Li9igFw95aC6q3cG/0e0rQza1dwVVrvdIphYDiM+hYb6+/l
41vguj/6q1zBo/09EXiYITu87Tk9ynalKHANmgKU0/+hyVlrZ38lxzixiu0N
65npTl+IBIyIaVkCJ26R0vIVDPkSNXlar1xr6KDudlZgP7phBKEsRcqmUG+l
xc1VZZuGg5TqkKNH3yeJ8798os9xrg1g06kwVeLco4ksiKDVxvTGGTslqJn1
6Dtnrgo556mqvqolN5rqbjoc+RW1ycK6zlVWr3Qm0XIOx5FVVGepK+sIgJX7
IAwMB6CxcH2Zklj1Z4e449YjdyejQiKkwcHsQoRo4fRYfyJr4FttHVf4W3Lr
YO82CAR0yHu4soy/Oq4zaY1wwP5I5uSCDWIM7/Y5LnttneBsUNwV7zm67Qxz
n3N3qziRg4LyIUasMVWw8QP/eXCeHmqpMfnfnguVbs/g9us1EMhl+S+AXULi
1ZdXntRQaMNjm8F9C/ICMfGCYrb/A5Ta8IWphuhi43XoG/qR9l9YZfIY0BAC
la1ueeI+Qq3l6ySbCz96cgCTItAiHFhKXzT6ZlCaJ6FbVWzHERgAuzUnxjlf
giLuLoc3Z6mb4dg4TZYgTGDiTNcj3XDK4ih4rL3kL0LfnxoWoeMqP6h0IUSI
OZBmHownXnPbiHWANl8ymOYen6p+eQzkPebGO7pUdmJCGjdgYeaRihLJKb61
49ogT0iUTQKRjkSWvwmnwNFbnPJJZK8U2AN7cv9rF5ROmzRCH+SU0VqqSknE
aEOupt60MWmDt7MoXw0d/gee4yxfAvOkhYRjNQTtckTCPMLp+WFQhw20EqnC
4CYQb+VcBS2c/7fjp+9p3DgqsKFgbUk0oGEkxcWa3nqjOwymy12YoHnB2X6c
6+JuGHGFY8ctQAsdzSp43pHJzyLkF5XdrcKdiaJ64YROFpJ27YoVTMzJiz4v
FVOi57cp9iFPD/wwWIN70CDtXbkurNqbFxTcFDss2f/GpGzODG4xJJ+M9bcb
/HEQcGTLeFWKJDBdadfifYj2IjjIa3IiuUKbdqBhP8cHo3txjvAsVj32dhzr
/PivAoRkK92JRj1RXbE9gD2itQDv3fc+p9eEpUbwJw7kO35wtoQUvr7RYcTN
103EWDYtmXOz3kHpFXP7MQqHdzlofiJ5Ekas+jG2yRmc/FcTDnchfi9Y7V0A
uEk6eF/uE80RhIzjI8r8tB2mgnSmJ22KXZAABr8sp57OY3m48oOpoWOBYB1D
Tq5BeoUpwDy7qPZQWkxxsw0D4Prrns1INxsms9z39tP+iMOrryouVPMWWFv2
+lhLRnJTYBGziMVIYgcmLKOpCshGIdukpLmaIwP2QQbVSdBJf0apB7P6Mnok
skNgtvuY/rLQUvwz6Xu8LCDyA22FpGnuVb1Xkt5DRMtqw1SeFW1l6WHATLSz
YeKstMS2Cj3gYg/DpwhIPDDJrWaKLXCDsQGSHlooQYm/TCcdxlN2h7qtYTln
SK3UBp2B3ECUAUQA87CfTn6Z7MXHpQGhqHcnBGL4xAeWnSjjyxUF7zvmZH5E
fGDM55NWb920bax26ufXOfDNQwiSD+sJiWHxKNTLAXMC/jT5GYBkAx1ZwzyQ
U9ULN4llHJUSXGgEI9BdMR+GcOPZgbTG6Z0GMgX3fbrvy5MLrDqxQnnGgkm1
iMJqHrY2mweWUAwtBlAHetc4SLv47YBGkD20zHsk9XK/azYYhiuoaXxTJyFk
pJks2BVF1A7RAfGIP59BgewUbgb7bUoN4YCCN/xYxXzjFcv6pmZ9OCIeXEgb
fMc4uZKSxnR8LLQShyLN/m5GJIMqU3i3de/nBW1zt4TX4CpS6ybBVMDUl6Jn
UcSVhRAKSGQlLxkq29CitfB0RdvtqAxa0BaUYXHGd4ijXJ7pJDnwqlgJOk0l
8EMXIso9qFUn4Zv0dVfk6zU3VCRVe6sLU8npTcjhm+DahKCOwwhT8c6mPV+8
xC/+RQ4H0wAi6fPKWVAxuOREu22DuwTxkxuCCmugFXFV0zsjaDhRR2v7rtk5
Si0/g468daQe2vV2g/wbKIE0Yf8CcJ7LdOVRrwW5K3exSF8sAfKcP8dNnCBg
p/Rlow1cu/mRJbnLOc70mFOVjtP5bi9U6b2eI7plrWpwFh5/u8ongnfVvrVX
rfNghW536calAwLolKIrv5Doc/9BDKCpLe4xGPcJB7BgNOq4YdsNvCc59AsD
AvENHlObRQzFF7yEQZXTucfcQCE1IJ3JqBXFqjUw22eKTKsx3mlicIwZbd02
WlrZSLP4UwY/jnTDaQjp8Pl4l+gL2nTd3yTBZ/AgZmaffVHcRNKi9rUbHhkh
5s+8kuK6rgr+Hw3oxOYyxypuCdIVeM8c3G36JQbWAjvRZobI08c28p8pO/Y/
2gqn2lGaVU+WJ2Us5xwqKRyXvS9rEPoVSrL6QKuUuJOBm9cJIpVKEKKkD52T
H5lVmlb0bsbp/bJyGFCGYrwlcmNt+8xMMryvFGPNjDExxtbsoqRhUovyRSGC
oHSzg0Q1dGcLxLJVUnd7QYCGEvl5fGq1HJ+MDkW88v1w1//bD/BhsxG95Xh1
NKpxEeQ4GSiq4YKBM1t5eJ2upCTnhiZZyLQ715y0ngxKXVRbczoahByQt4kQ
VhRM8SjBit3AVoMamD0H2bph46ir924Ln2S7uqlaDA/yzXF0J3oRE5OUaEfp
5zsqJj61hQpH/3wng2u51xGKGTpqFxmXcFVDTkXWXDt1CfRW05chIUifBkoZ
NFQtbnQIjj72aC46yego89uJ0dF+Ha25jlLpKxYXXZx9fakat2LmawAM3XR8
Av53MPCcIQ+tVQ1FbGAJuRdrPvwk9CXFjewu1Y7wI8UQWZS4Yqp9kurofXfk
L/MX2xyJivomBKz4WZ4FDhtqR0cKmxUZ/68QRTHHyJTkJkjMPkqxL9DLCI8y
j0KqRGYdCYYSizMmzMTjkGUPPaAzv+f4pZKDOv8sNo6+rqVVEES2pJDTWM0s
HtfcHlF8U9+r83yoEAj5Hwzspt8+4yjL80ChtQjnIdxghPtKJAqCo35MfP7m
1O2XNMw43ogdbKlamS+71BFHFnlvoaTxWXqlMjNx3nmsUkNd0fP8aY/6hUYm
vwZx71bkA5PjcHLmt7wslAu/sPisCbSnyMObTXo4WREKzPUBxkobri/31wC4
xCI3lzKvDGjpJ3i1oGVEvA5l/DoQCIKagrD/9fq5ZD0oqzUGzu8PRsdVsxIM
QwDEW7denUkkwa9f6cjRbAegUVVOGIUVcTi+34d0jXa6g2RqAxE05aesEDlG
OGGc1XWyGMIG9lwAHtrkUkhrfBmSnfNaFZA+zd87DgEk5IZCnVBdMTmJNMQz
OvdFSoaQmjJbFAs4m+a50PhwBfVfPMAnT5F6rG5IPRdKJoJZ8MvRFVofsDOH
9j85ub0mN2gUlG13XjJesYJkNlGGHgEvkmZ5ieRCdTkczN8ICLdkN67FWiUt
s3paV55zFl6gLaXM6Upg6mol/znBNIKbXyLhAd/7JUi7zQwSjPnd7tQXpsdR
AzVeYNj+0xvgTNB8mWQ0+qm86xJ13UIhgKsCBnwWaXHMYepx/ezvZGxLWBv5
mJ9fK6zQjVmlgEMgKnDXS8c4AGjoFIrlIlu8f8TJOcUQeRfC6f7lKpjvb+HR
zqOlKx8JPvF1FZ8Hwv+wjzCBTBmilz4ucLgCp15XLh71uGkMnDD51IDeXDBA
3S9aeqiSIiIvRyudcmBUZM7N/rkW1MLm0nm3JzB3xUktewUkdtnbtJMTxZwp
0xoiBQzN1NZD8huXIjmhabnWL+PqiyYM2pmKFs0nWTkTNo7DI5a+9vY+xGR8
NevYHcKiytcKAJxZkwX2poBfuxwJ36rNDkaBlbyWTWPWH1cnYYA6pSoArull
mGGUqHaqqBSdFbUM+CzRUQ620RbT58lQv3b4q6KVBH7N2B5xEsyvVJ5ETtGD
teCrAYp8h7sNC7gZ/nL61w728pDOGZj+SoxtJFwWX3bVzPv69YOLalp1CE3H
YdsX3zWQcZfUEPrM6lEp/uwFnaTz7QIKee1e+sUTUOt9WWbNT+OqWSMJqpGM
WoajGiNuA2ecFHVeUjhl39UTap0VgIEFia9X4jn2H0LN2FxoTpFlOG1OskBB
J7WCcgxy8EFQUATXyMWP7z2C0vXz/Tbuzd6huZGMCFjVIaJF01NJVty5OtsC
v/bQ8tU8wZX5vWYj2l5uh3OWdo1x/88/4mz/harXhUFZ6fxcq6BD001MGvL9
ugeYYu66U8viJ0jV8+v6G2W+TsoaTS59W+dvRTpgtF8zYG2nDt8AT2vqxjrD
COJRwbES39L83OLCwwh+G/shwXnD0gAoK29Eq6NxRNibqSkb7/0nNnVnY2gX
g5RfIWzJVjYNV//p44pB6Bp99CDvX78HfVacdU1GuCd5nw9GhGG4gJyFYDrs
Jldrzz4W72ZBpGtfzgTc52cH5sBvLoM+gev7XK+JwnNQhliunH1rRbFWCDn/
I12SCi3+2X6fQDLNsT1s2NK1Llr6rBO2JEjTkkk/VUXEmV7ptUQ/ogVXLF7P
pZyQ0fCQKDitIxrBcA8+dbQNJ+C4VteqPkNYQHl2cipTJT86ezuMX7PeWEe1
TW/R5Jrr9Tpu4QUOvxwIKgmt+dfq+NFK1KORVM8FRjjwUTFqx5GU2fpslF8I
hpQZGqPL76rDvbqIqaLZo/0JZ6+Sxu6D5ise4UEe5VeLzSSsT28a4iQhb8kx
d67jU/sVaFF/UjVhzqUDpw/ww2Xxnl0tXPvHLdpn4vDEAQA1RmG/7TtlKHja
w3QOYXa4kWZK2k1N8aYc0YLUU+35pBvPr0VKOCXfmSSiqYiGq7I9Aqxhtb+B
ucOOTfE9g2i6F98tmbT2P2gM5WSXUqRrr05fy9gEoBITdKVkDQQMimYU9ow4
DKzbZSnKp1WDF5y0F97jLA/t1LKNXSVo2gj5H46YVKTFYNOyfh5cbQzbM6ez
nJAea6spcNTl77Qykt6hxY1eGFUfMPg1W0GWNlAo/M+lnT4bMYa+NpziRO10
8UxkZmvig8+Nyjx31bqeEwwGWUT1yaMAIbgYicIdzcFR3GslgEemqJFpelQO
2PXYLQlaYGCzD0Bp6vDtP1gU4PCtIDyp6qq6k8CHPtFe45Qc6TsovFf7iAgF
YQtXFMeYMM/YkX2ZFcHWww2PbWZQ+BKEcyu07Hglknw2ckKbzo3DEuBit8We
EQ+OWcZesc4MYDPIb9Nk8mLTwb8SBzdUVeE+XHgAOlqi+b70JFeKhZkRo8Ch
V4zuZnyI30n5VLSiHb+zFb691P0qfJ5ZE+dsHbC4S4iJFShCc8s5Gy1pwpk0
4qnJVSaF3uGZkq1bsauyC+Ccw4AK5aPz3es4PlzuSWcnIj+rK51IpyDRJhT9
/ksPehlurfGdKX+QQ/VUkLRYDrwd6bKLXTCBq54WTO+Hg5gZnI+wExyBlvNV
qcj1fLTtEiCSUzHMvKxpITsqzbGaLHDXq+NiGOKaihAtewxsxImIL4DZFrGR
uibnt1znePEh8vKqSlo71xIBVQijExwvQVRIweGfc+DD/0x2Dk/DNy++zxyF
5B/V5WAr8AA4f1UIKeCBZxw9sScxRCboDFlWfubgWDFcRuu7URFiHn7/Go1T
XAVsKQJiLSkggdhqsW5quN+QbFl/5uGG30rYEXcU/slCjFmUTNs4195kxM9f
iaFmy52V+Pr+EA2FSsbuegeSGxTAuH8nTQWiAp2XYOQonlXkmQwq6iQ/F5ba
vhvqTlmmuDr3d93drKpXwzI6xnbxwrbOlxkd1pFTfMTJtyQiTUHCZYoptUEt
2g9xzScIhx8XYkaacLs7c5cMT23W3jFNaKRMroRiztyQkFEnUVR20rWqtr8F
UXxAZZqv8SiUe962c/FP73JXLfd92eBcycMgmt4OpRBc/fx0abrsEFfWpCbg
VL99priiexoz5U4orxQpQprWzvbYXcy1VBK2moSPBlO0La9aFWZ0mEsyXbkO
rAtl7uWKpur4q45DTcBfSSYIFdFG9CVl+x1cgt1dufUC6/+sy8m5YsMfBWye
1CqQCbkuezbxvMT9N4QT1YTDcheIgrAf84zMWhSt26SyiFZVitL3EQYrQMOf
9JFPrq3Vgs3P6vGrhmjrZAIMXwiGUzYpH8MZi36SOmlkxjg0nWMGs7TOHIdR
5hM0+eUhc6uwMK1Ng9KNdNUei/9m9UamfvzrstbTHtDFpR7LzRxE4XJs21yt
8jAA7ufv08Sozn+5dADMV5ZmDNHeuSLCKpaz+dqJCJ2TpZI6vHd0LAZvlwu9
ybTaaMTTyvf38v52z2VUfcL+uFxa5DlJtvN7ZKEMLMaujm/Z2MfUCEeZzHAK
WGPAE2+Jqo81hHWkY2aQe8M5YTjGuix8/+i20eV3545FR8bJbZYhtsVeeDxl
HQ/gBYMxGdJW7eFVA57OzJcGcggMsQIJtrvY9tXSTgwFAmKPT8s4z/M39SXu
/z9j4g4aDBth5ZqbxWan16iDJEJC9mwIzglsZf50TKHufySutdQ4f+LhIfnt
xu3q272ePfOMqKU3ZeNG8IZj12nj8lPVgMQIdiEtnXX5otDW1bnUOflC+siT
ka/7s3rgGKj1aN3PD6iA7bHx5H4rUZ43yhfmtZbKhl7JSmriMTQc1XDDdUPR
tnoKCkGiMZx2kcA8CazCpQmDMcr9GCzUrs6w6UKGtJTW8B8sfXLeEUir67T8
uNdCpGEs0TMkAGefRIrIVzKSaFrjfhGUBX3n3d5tyFa9QHl9JTQUFN7ddQvG
Nc00W4P63oCTbNpl7NJlbEef2KpbBD+JEcca8k9qo6DCbboMnkV4UrqXfTI4
9ynHjaYfcH3WhS8uKnmEYDj0lk4Gq2BMz72w9jtk9/oNEs/K5AjPNKiV22QK
b7f9GkKA1XZZgN+IXnMZy3IYaeUgafEF2xYSaOtJtKgUHS5PlqrdJFjMkOJw
mbNnv4Cuqx+/NP8QGxDNnnQjmWNQ3WKyo5ywpWTC9Sjr5axg3tFe0iIqAWUP
MzUlulujKmz/v4p8dXGZEEJZU28y6JsGpzApco3PbSY5enNUUB3ok5oA1+Gr
u/hqUqj3MLscbdJxHrcO5hWrVFFjT3h8NAj9CzRY0DHbckyolrqyZm4ndano
e5O6Vg1teffgSFCY6VJ5eSZRyXRQ+cV4jV20GC3RNxD2LofeW8VwWwbJK1ck
QCtIN4oSU0mwX+nWCjBy6mWmlgczS8Ieqk0fKhPZ4QT6QaYkdEfSAkKpG10y
pwAtW0HRo42SGNW71kEdSBksJW32HYpS9XLC1sFidpQ9qJcN5GNaP+hr5eSo
PhkhosyZNFHJePa0NepLOXAimfYnBVewSnwh/RkKswf6zuSEVjaW+HEf5w2p
M+FxLk/HDUUR3rnbIZQuuVfcIY/p6hGidKD0Bd/aj8whh6hCor6umJs1mLJ5
vIrfr/dUCugjs4lE+I7glb1Venkq1A2adQuo5Iec3SyXUdHhRk0zgDMxeRQ4
sbB3Hp/a7o+l3eJg4Z8P9xKFHSmLwkAFZRZz7ZZn166dmy+YkrmcXY14naCR
4ymfYd6QiJQoDw7wg5TUEn99Rw+2WXciQJVNAtxyKgsFEmlOP28XlHc0vn3Z
xYjoyO/zC+XLxbDtDp1VTyiUHVliCsHaQI6zEcqa6ggBrucioRz52Dob8eY0
FcP9kQSXiccmHNt9jRPW21lQZXMpssV9e+YXxkD6/mJ3iYXrYftlioE13MSr
gua88sTN+ArfmXqgRMQskJv3b4ttWKSvHntcS4laj5CZ2Jg20NF6llU4qNfP
2GIRlx4a0zLo8EHjrNH/FIe14UgISx/OSdUIVebmxeZkE2P7C4UARwxQ6C9r
hfH5dRrbVzULMZFw/JVXebswQBkYtbiTARrMQn5/bfJzqIGGA5pMGWl4Rw0J
Zeupiu1VrfXjFlgv7sodd2UE6LoqgsRD4ofGV8lhYmSOEZpa+DA6Ng5Kan4u
9R6273sI/xvPZ6R8EuSJKKtsm7riL0lrLHYcT84EN5tHxNTDwPpZd1sBkKkj
xYTHOsT7e/tWSfkrPcskNxA2+7lWgmnBVBcqv3bXsFt8UgEKa8/Da/h0po+4
Ing1IC2B0NysNrsEAh+JoIWBCwV3C3Vc0t63WB5QeQw1TvOiMr8wjStqHTQS
J2MVnBOPMkwqYruIro8zenQ3j8ruceFE1bpNA78iTaBX54F5M2eYSWuExwRy
8shjaJBPLkcOUbrecJaa+2bMPGRGe11k7XuMIJmpWY9SG160/LKu5zsch2ib
QsLSB4iaqK5+NiR5QbRERAjNzG7dtuBxcmh03eeL9LRryedPv8Tn2QUCG74Q
87B0zBRFWcgw9y3u5lCoe/k0FBbIhNy3mbIui4YMZ9RqIBgFQ6UMmEAVXc8g
XAU9j4R0KDZsZ7D5XwBLuAm0DVFWWzOMsRAAaHTMyV8UgFVkkDwDABKbkeuI
FT/gcQWM687Q0oVXx7si4bgX59paZyUy8LQj8hI0npC0BQ4lJWcVEF3z3dWw
wSHkjOh1GrO/Vvvf4kzIOaPllWWJymnOfj8bBXeq3I3OhYS1Ppe0G2zkVzYe
mPtCZ61iH6MtC13bkCMihTEG+PDN8VXhZRYOa995oYuH4a3IPZiD5HoymF30
jAhk721ubgRRGoulXlHY/d5ezSrhVS77QuucjbZwDeKGZ89GtoPWN8VcrBp6
G35aNc+NGY8B58V56kDWWpiOxHmGM9EStLnDnhUwbcXWaNKx7i8cURl8s0P3
/xOV2dgxGHM8De05eeQ3Fmnn/+gndzjGtjGcrOURGGOnWM9+vhXZG3Yq7Wlt
bYwfoWxkfTN0LoChxUdZy/uc7HAyPbOy/WIxsbQ0P6n4lbhxP2W0Gd0zj/Ao
vhTjBP1jopjCrQ7XQlNWzC4i+mDhs5zF3DVeMgqMrN5upUM7s6KyyHSXQOXu
YcepScuonGUWAu5pY78l9xfNhbY+S+j9O+WFMNhsHMsdnjM2OKXeS/RtxFPj
DaiogEIdh+rtJUKQUAUZndia8Rg+Ip4kJAxu6QX6v3c2iu/d9h3weQVTUUTq
ZUNhVWUIQtiXzwz/NsdpdDqKQSnAytZkvFoN5ifMY6DBQHB+wMApCQFl4Rns
S2iASQ2F5YVf5AW6YBOqQfhuM6aXeH6G7hMGV1GvJbC8tTYQQE3QQrjoJgsz
/x6Pbk3wJNlN0hlQTjcXyI2jxbahOZbz2P5AuWdvafuT1+/LN82VtbP+qBYO
dxs51U6TyP5rSa5ZhIMYHQOkfor2J8JpVIHpoa8cbd6YpgAYGHdKyxTtkQdY
wpMdgt5I7VOacWZvJHw92O7sGXgXujOqM7QW0FFlWoVg33hPbCJkvtXpw7zu
NHoIkXFCyITT9OoGmn7V0ExyhY1PSQwPpDQelYK5FO9CzGlyD0ovLyZZntOO
atz3EdLZ0WDJr0OT/3zaXZR/3mduez+0YupR9Bk054qkgnlp3KdV8G6yN8xG
pYyKDMXZLajuRRpKka7l0sYlQlw0fcgqNUMyN4Y9b5Rn8zQntOg5aEegqROU
f5dQHVzbUmM3rLWFy7am7MHmyhkTuqKQweyh5UAL/ddSgQRdAK9PQOL4+D/o
hlOhHPLfdaNylsQandmGme+He6lvMxtu1fBFK8kIKeTeBTclWMlF1vH/PNA8
+nyDnvvnsiF3FzY1DMrShKBjZdnkqPiQQPTR5beRyZ1G661gKkVzFa6E/uiz
k0aDf8493zOJ/jJcrW1vTELpNt0A4gP3pJ2e2QmwH7r6hZCZ1fw+P1Q9JVkG
f6bZIjX01kMYYXZeEFaKrynRIPhcIXSUJNmBybOPssIpBXtZg18IBRPCbKND
LjYfU023UIxJMGdhEpv2HPrzB71EYkrvUiRmbTlHilx9ddF/1UUQ3F+kI6AI
SmrpCGE3gyayDI3E4a8ch0QQwPN5+5Dzrf6DJ/IgCEKvgzEsEohlIW9Q8+RL
nW6cK6MRtyaASSloIJFHd9xw97gfybH4MUiPJhKhLq1pJY2L7syZ3XUbKfZ6
VJrPPSHarxl0aFEcX0Wqq+RjdNza86JHFmbtlodxNCEmrhE7acXA2VcRFh2B
eZ83X40B2vkoaQn2/jvdt12tCyZWX/VLZd/mFVPHqkR0ZA2QANswZbb8w9lY
vSgzG8fGsf/q6sHnYk86IScd13PCreNX8MAPhAu42AQvQlVlz1x2EzkJ1a4z
VF3fjc7l5/8S8xFrDe2WFfeZlPL20qqzSUtbA29sSGKG6uJSQcbiepa21L5A
2YGJ80gQ4/L4s5lzL+qRxg/MR0niCPFVy/fAQ/+J2jK3Ji9QGX4fHK3aHjln
gPgYGYkP+R96RoehfUwSO8c1Sf9yVbjC9jqxba7airNbsU4KLWcIFy+TrbU6
YGgUTy7EPXClGAm3PvcOn99bFfb4eVf4VbyKBlmmmrsNB7WwJ6pxrBuoNeyW
a3NgkVOEzQ0LIblJJLpg84KLljbsM8FQ4yzWpR/SgUpX6kpEwzMzSLUIzZPG
NAMNqJBmEXdcKG4C6pzuXaBaKN2XtZKP2MMCkEhtIrkx6gxjgT9OGZOzuUzr
UP8FMUzH0eCG24iwD1iIbOhm5e/yu4UGBBeTBwX9peo2TlDJdWj2dKYtS+YL
Cq+NlmDi5U3EHMnwqqcuTq94dcahyltrbkkGsaCic7jpkgI6E1mS643PhUT5
6ua9AYqboVDhcYzZRDhnLAxv4YF9GqVaUP31o+GhCA2ZzrhWwv+9lD+O0CkR
AzOY2m3qapIF7g/xMWg/gKo0FMo7vDXABDgkHfpFAFA+hbEx9x8x2CUv/HQQ
0F0UvhcjykWs4Y3I2M23Wq3K8dKHbLZM3qvv0S4zfwHwTxEZskD/jEALPPCP
GpmZYzLFryot0y1TuogwMxNlNLgrj/BcGj5yLuicW2cVUwFOi4e5akEVMAXV
wQsEleCzjQftMis55jxWbXV1yF7V/RUAgq+FYofwI8OUvjJMhdC42P6R8Hnt
F1R/jMvdPpPp/0nH67Bbjc9czw5YZKdnl2B/CiwUj5sgmqC1sLmA1d0q0sZQ
ij8WoeZGj1SMScuryfA9+Wy3J/dW+iWpD38miZnMtXmN1mJ952yh8KgQxos9
e8ONQWyarlUuDHCrQOVKyU6J87n1hPdotO2ATd95iqyuqRGSwwy1xaEkvKLm
k5WhNoaOuaFW5AabxRmDuTSQBsw8MJQRmu6sf8A73sZyY0fVlqQmg+Y9QsK7
KECEyga2FrN4G8SJWSDF5mpxUy+GVGcB9YoofIj+2Wj5KBaplnc/76YnH40C
cfYA9YdGu7CX9w3jgKy7y1nugSoS+f/oDiZ+Cmo4BenVjTkqeuWSkVFA70TN
9nBI+F5s6PwqV3eMnPAafFCD9J5/mkgYVPTUmuG0nLDZy5c0BWiGOmI7z0Of
ETqtP59D2sh/LnldDDg6HdHXppeX5EiV6miVEe1g3NPJSLWgn8XionSx1X6V
NewkRYlQrWHcBJnsa8qdkxAx4skM8VeZPUwOtCjv5KVVvREtpsfFVE5WMWBV
v+kue4KmLKSObfPRUAnBoq/361RWULvSn5MWdGZbaX5Cob6vDrNfe8vDRpiF
od0X9D/oelkkpx74tiCBIUGHsi+HvOCQccYKz0bMmD01bS0lYOCWH2sVVd1N
3SwJGSlzE6yhwn5bd85GeiZgwlze4gn/Icap0FRfKNMkpk6WGZe9etHpoSbu
e27gcdVBbxOX/O2CG8lz/+QLfcjIbkPmGB5QQy13tE7bJqARKuAUnDQ6dlzl
4846TDRZTXsorxAIc+uUImViAIO1208YE63FZISaFddHAX6h47Nu7UZPsynK
9w7vjRHjE/5NGhJRhEW3LJOIBPc8P2tdCwfAp80tHVkS/IVUtqFp20rsww7N
I4j8RVONTGmgraIQ7in/GKSnRG4Eqx9hKnHIc+MbUIHlq98I7zOK4kp5fY+C
Xkfn7buhRVZLLtXLka6ntLOIHg8lyDMAnrv4k94vXNSy+w6fJ9zQuHDODejF
Tlsqnzeyv1HVqdFrPJVRhGKaUyq5rIlgCS8olhtQP8jCN0VxZ9d1gBkuAm4i
H4XeyiOfUhnLdGGefJ4OFFInswh3ICnyTrHW2BDobWsHmi1+ROA5x04moX5A
PLJno61j2Ji0oRoYTCsYGo19jJh9KHs8CUrB3nSBRKg9hUIerXg8knGM5oub
GVmTbsm5Di8toc8JAYUpcmchd+URQ0eW0Xyn+KLCCOBLanHw/EgB4lOmuDcC
IeRoCNh89u80xDM8BLn8jP904t0A5FWNcBzmAh1GfNVkhPITYxVdA+DpJCYa
bSsBjdBKQIZZxjNFzQ48AJ29dnXLK4gGaLaQB9FJ5oJ3zq+nrOTnbH+67jSa
y/MIxHonyuK9oTWABpPwfm3qHxNMjaeA61HnJ7exA5gcBfkxsOMlzNDWMe0b
bAjdpOQ/4ca9NhotLeFslM12BN94MRhTGfsaxxPEv7m7argd8J4z+fhJoIuZ
/PyVv0muyX7bNzFs/3pnHfeD/Nxk9YUb6oMXLMV4S/e66HytJrc8nXQQqueZ
Tpug27zFV0XZG5MVThBk8/U31Bdgf7SK7GuN3i89e9ZAcK+Mx69R8HAfY3+j
cE2S/OgTM67ebVrQbE5GsY9bqtxSFZjZ4kBh9JN2/SZxG6oD6IAxfxe4Jpfz
Jve+p+HRXGw5TXVRLZRz1DeBIF3iQ55RHkeNpwMIb465LvrBRb0RXgnHsDTg
vKJFn9siLOO9b6PirT6iKiQSbRP5zZd1uhyKmVsC8w4VtG8IbMxL3C0i3CKt
sFJtHStHGN5vsvb20wOd2xGoia4uOg0x7UjF0EigCm5Jy3keuIECeIbyT4yi
HA42h50xPCbTPYMYI+jTcpTdNhMcl0WZyxz0YPDyDRmq7LiZFw4znCrEUwYc
gWIxe6Hevj0zqYXGu+mOR7G5GA+i73/dUUFX80iHCoboctbY1EzVaJFuyAwv
wQKH2kYGcvrQuGi16856eMP5aWmjOPC/SjzQuHp4iQbDAfgBQxMVw5FQUnhE
blhCROzwrVaPoj72ykkOeyLurJst/Nqz5Rqd1xZQOA4peBtyB5krsRygqai9
Kg9srMF6fXDRzGJyuJjVT5r9eRsvEjq1xLJhmQ4z337vzX5/S54g1y34Y4EJ
kWxDoAGVW4z5PQBKcfTU4N5R+j04XjqVqFESD4jWsO4qgjXh5VJ8EeVgTuvM
TYBHV2pK7Tljj3Xy5U9SBTOR+GWqNywsTARe5NlnL/0fXDteqE5hs+cYitWV
yqvu4l6vASluY03JhhyQUpI5xevDAJJZpWd+9yHN/ZA+JGPfmdG5ui+4hDa6
/WvoZllfnIeitPc6GOZ7TLh6nad5rvIqbzEUfFVQY7dh1/Lo1fh9MuREMcDv
bvF0DHjHxc6B8+qZXurZHoSz18wimJuzIhFFOGBKl1OdTrMAFmExGspRNc+B
fbyKNtbFYfRZa1DLwnq97igagLgzz5ECXnXptRBUiVlKxe5/V8Urqg3S2If3
5UfS0aWVu6JthEhveWRk5XBTak1x2EJZzpYhzqZX9NTnnaHjAhXoj6ifDNeP
BprIHdJEbYjGRKW39Ws/MYMN/uU2V1ZuHVMk8O/bjDVHSxIgA4zSOYzsi0s9
gncp1xf39+wU94ORvOk6GbWbxDIk3ugCnYzbY/a1zPsl9YVOceZbnx71P9UX
ArXCYZiFWo1BVFXZoFvmjTPzHv3xowyBL923hVHuRSs7XqxDQauWC+tioPo/
ejzIGBjKnrzrKvcBBZVamLxZFDEwVLtQn1fvH42F3C22CTzM37QZoQY+l3gx
RoqiGmkvUiMtjzSNXeMvrhvZbrA4H/ylxfpxKjakhXmWWHgyK0NJ1cL4wlPu
ZASyo9v2vMmzJTyWXcsB9O9G8IhSrAHOhlRYGjUN+XIDb2wHhYjTmVgETjQc
8ETFSzqMdp3o0iQis/E/zEcbImB0dnraes2DFxLPSBbmmh7z6NZoFQN5NlQw
4Cum4sIW5ggtuNHvxCF0msTC6oetI+pDtL6zuL2fr+S0op2pxisllJW9ogny
8Wqw9wuz+wxxNL1H44o1QgU4d4tV+7bUqS3vFfv1Qwo4Lp5LWYBgQzD9UfF0
twAgD0g3BvLjGu+5Lj89eojp9yaDKyBLr6Q/29Pwy+LqeTw2lrBm0TjgGB31
bgzgqVc6Z3f17ewwcAR1uOABjLBgtkuM+JsGnh78BcCt8dbc2yzgn9EDQ6Kh
4p9VsAFoeX4WE+FqOUZ1WGcpOI4PqQt1Arn1EuCs6C9DM2LlTORbHt8g0ZxJ
YlKBEXvBjQgb3aaiK4IiQdzsL+BaPXCpk8I4amm9C0PJK/zVcY2xW9Xq5PAx
KFT1JXUn5a483YA0VfpRLTrbyu5HSfVI+anQeHac6Z8ou9geZ41Qls6ksX54
MwJQHj8UtmbWZNMdGVjXmrb4OSUyEMbkCp9wh4EFBgCfjsNIABsHisc7DyIV
2t34BjehYV1VrHrgI4h89Qrm/y1ODqv1+/V3XGscnEUKG6p8sZUVNJqxdvFu
tG2WCYNLuTbamSGy+76STTuwQyE7FKwQlAT3Eo8ayojXQxc0X6QKH5PCzY+b
j5LBnCkaTiWUSfEMFRGcVasJDcsHs5GTQ1MtrDSM2uMzDCmlwr6j4jb+QJTO
fmTcQ/ZG8hppKLeA/U+EWoISu4OtrT5vV3GPTlZ7itYfI0qH8wkynCw+hr20
iJpBujzDsArEii6xVcyFS9+0e5V31QKHgr8YxnLdqdB2/XudpVH6E9UTHbMM
AhO3iz4Muc7yt899dfwSWB07anZzKOduY3KcZx8o1rXgk8xrjjP/kaMcYzRY
iFHnt9Q/m131lMxM/8rVpFsjXUY7pyYZD4MwW9KbKMDpvdLoPKgWUXxQysbO
Geyi7eqZjRX9zgJl112Ler7lexs/BlxgxkstdHYIS422gpk67JubTWMDRZUS
nzip2lugRx9/TFsCP3wuODRhYS9rMAM4PKCoQvr8ejNKyHROQQGEHFlijU7A
wSbFngI1sxv/BWsPkator0PeHTa0+emPRzRLMmJ7+dSxTjsDkQ87uZiXM7p1
FsS6zKc2AAqMmKW3j18kOb0DdGtOlRhEGidK7e4iRrb3OAuEbrrnI2FzVnxK
8oaT2rMylgigmmb8ReVk7IDYKC7a5UuEE2bfUgz19ZZwia5Bz/aULXQ+6s4c
rDp7Kg5Vu0V2ECJafqeDF3atwugkSVQh2XTM+rlWwPlP44IwUavN7GiexGXi
VVz2RFdCLNYHiuEM5XD8BMEh1TBPZRxLHfH5KQ1Uy+Q+UtCtQc+Ew2eOKjlA
//+I64fLF9H/XWrEP78U0DlWTzfQVeBV1mM5xqSTNFQaR12uSk9wOQGjudbj
mkSENbFKi0340vYdfONhk8aGLaWtONK6L/bdpB7+9k9BnvvRNS+ORAap48co
s8FDANd3AA7cc6DfbSmuVdxdOWViEjB0ibGGXmMaP40k2pDQmOegURkLor0g
q5kZxye3tV4zHcLKnuUWB9BIqXAXE7ey0Jdq9pr2r9Ji2Anm1bAvO8WLAEL1
1rQB5PwkOTZHxAmgHPCPG0xkeef4Dve0X4WZtM15TjejjVU1cKh80LGgboqU
oyol9f657cxCT2ufbDfJFWQGCaQAuSxDnm10NSFHDal+DU1IFf5c4i8NNq+X
mTs5sF2cGxLYU6nlSWoA+18APM46mf1EgOhhyIGNyT+1u6ugGuImg6tV8iN4
3iGS2JPq7RPg42E+MrgvY9pROEQdRtsch30QqZNOmSuuxRYH3Wzoxa47PVCm
zWVLlsu2wtH+Se9CprRtucDEK7Mc57M2EFi/JNH2PpbRVFzkHsftDE10NeDI
GIGTZ8kyqysEDmoeVQwVBWQjy5EL2NYEXTUHMNovIhlI4rPV77X5M7BfFjct
czkIp96czZeGFC5jYq7eR4QPd9qXqc0nOlbYkMS8rqzGLAVV0Cr7vjN0M+uw
prpLNQX2Tq8Du0PLLz/YusFt+DR/CdhThoz7roZU4HPaY2afKCguKVLCP4wL
VXAAT5HnTqZOmfNyO41XFcIqIX4btYBwVheQ2ZNC7rteduf8PsRWw3SHB9e1
eaLCt5zRnRNtVG9A+A+ZqtLtbGK3mGpkBG9s4zup8dJ2QnNOGAZlcOgUs17B
TF7A5sLUg6Pa4NVDmC2Cde19/Y3LApXMZz7Yr8NqVJQCALabI3LuMFtQHXOP
uR11Dqae1n5bEJGirQSfy4RVDwhqmVMycSgM07kMNLTC3HZx67exWsj3ltpd
udhCH5r+zkpKSGI6zUUz//GZLbT31Yi2n7WURTCl0CyVnJiru9KWY6V72dsm
g3+4xuzlUTiELmxN/1TbHhmI/vsjzp14M7NFQcNHXEK2mFVL1Be+HnKDimp7
P5zp7wFgSveMgr3JoTvCVf4buy/O1odb0dPJnu8LRC3SqksSINyG9zlSC8M0
XdX0WrPkEfUZ+ZSX/n8e2OiTYyGPNxKMUv4V4yhFuLv/edmWZgQfwbdszSqL
rP844C0xjc9dC4l5sUhZbaj1/pYYYlavvxdtJBirvJYAeFk1qdDAd3+pUiOH
GE9kx+2V2S73CHKbAP5o294MvZse1UT48SM3vtSfSX/167NBaJgxslf5QE/q
h9YihInT3lTn6qUwjE7KZzCwAQMtKiMSfzp2+8/kab/uSwcBOCUG2mPpuzVL
6fPWWG39LconjJLg+boSVUb2WRnKc0rbgxune6JIpehjH3cQ1D51MH7fTJ5d
MNfSSGi64DLQXxJNMlf3JcNAs7kgoyzCzqfRGxsaIvAyI/BAilCIrfq43gNK
wgSUPh5LFL2iHcYe9K1hXDRlBdBcbBxSrjcXOdGccem2i7mGxi5BQhYkkkol
YD+D6wl/vkTU08V+eMGi9mOwLOq5BWTRadml/u7lZ+9qh2EDDwK0615YrOfI
YLxJMRzwqMnNWxrVsdkooZyOkmRvnRrLHRHz78gQiP0dcSLSjl/lg9ob9WVj
R9/P9jSRR8q3jKmvZMaxE9fvM3MI3GKuiWv37mnKykpSvDjqvhZZpb1hk/gd
WRirw2DwJkJo4nR+NMTDuvXXY2gAk7034ItUU+RW5jyqjsn9etkTJrH7LLE8
8oNnbq0NZP3YhlptdLysCdzmfjpPmgyqgdLcG/cKQ7LERK8UoaCpw3Tx5qAU
dCXIIiZRvaMK2GRY9q+QceiBihLRJnWPm0MfqwAc5eyT2UbjaPBZVXi/5CJO
z2VGQeP4iIDnlbSrgvHNTYlUpEQlwLprVufAoE11/OCbWpsEyh7lWSjpTWdZ
fFziATa2AHiTrv+42nYG3om3DIXEvr94UIrvTrzHpTyHvlpParDMapbRCMOT
stuptVOfVC9BNVNbnw7QOLgdNfBbaRJ7zpBWRzjhG5lWCZxrgMKppFNGFhL6
nikwrOe3Ab0SfEbrR+tjkTKQA1KUKuH6myaQJrHd3ybsDs7n++AYhZ8u9Cjs
PMDkoJFTN32qP749Yhr8AsMIM2MB8JyhfZuAsGXwr4pOQGdyXXojfKGnNiKc
98n9OBegB10bAGa4v08ybI3opmmkELZxfg4q+0uxp2V5KHh6QPSgHFJpW+cY
mrw76QP8veo/oCHA8AwALALU5FLNF8PL9QZ8PrIc6J3qJt3KFPtmIV9VD4Sf
pC6qQ8wbc9Y3D7/6zL3vzqISFYFi9w0WN4qki4tAMf3xdOg8+xoTEjtJcTdK
ehJBGX3RAwL59k5o/Jma8lmSJ7C3K/dRQyIaxiB/jiSX4iLFe7KerEACiGVP
WKZEdK4PJBUXWBkwivnnMzmWmqKx7SisyzbRZn1sbIC1llSk5UUeTn7Julf6
POubpdAGmuD5ZRobM3muvTxe9KW9JPD4xC5efn/fICncrxP+pzWtlsRpxCnB
nuE6BnEhJcbM1GEfp0sEJIiI8WZZC4ebw5slL/mwvg5EAs/OhXpJjCnh8vER
MbOMeF+fmVnw+ClU14wM+8mg5jyLsmlrqY1mqMOmqzaj55V7Ze+mVNnPWpc3
uSfJfzwoOXtwblRsjRtk0ImuvdnmuHSEjPCigPFczqqGIkOAxpuoRyaXHSm3
WudbKzsrSUzF908G2lh2zIvmYMIF/xBkHGDbrmRcsTPmRB8DFdDLJCNEkqLr
y7ULp5DsgkZDF9qw6uTaakNyQw/zaArp5EgOx6MFJUxNFBjlhJnbZf30Nr1D
RV7kBG+KA02UR3IoSAKdwO3IbviwT25Tw+TmUoy0wu2iBKrUlTDPZXQd6xi3
PyLZdiHz/PzCPTomXnekLKieHlOBDe71c+WG9XMKIu5j1ec0oNKGg2Z/JPaP
viFKEup+RAl/BiNiDEd9D/qnIAk70iqWzdZN3uv2dSrxBgY4pumRjkVty1S+
BX+0F3Kp/YgkyHJ+FvvEfNWoeFWnvlmRI4882gSiU7F7AB6bKMpr8Kim5ySq
+I03Hm4TYigtGLWaALS+Fcw2NLzVeVmzekL/Curj+OjKAGVeWy84Up0I7ii9
jxFCR+7C/6BuhzVpcBIeCMnFSr7fiJSd/OaN14cI3Kb9LGv7NwcuezQPpybo
wogaJTVo3qF+iuFSABWYlUMGDb9cCiANjuWLVoXUcQvp3sP7epEImFygzue4
rnI5RtqVGsNq0KLor5/C07P+duswviN9DW3HgFBYQy6JRn1YxOTHNI46yP1R
YnnnDP1kDiyHm3TtWMLp73qeZFyp2kkb/sQyPoM0uGiu/wX6IeEKL2FvTKUA
Ox5giLCHPuq4xTYO1UaFQlMREtq9Jx7zmagoQto7AXCAceDJCX6zDis08xxR
ZKy/yQm36R8xwhQFEtVBny8yaYmpVFCwJtN9mbzKcl3WSNr08lXLVArfI+u9
kOJP7OCL61u6dPJgsgW8MTeZO+isPjGoSV/T+A+hVtHWkI5LA1IMyPJjzdpS
K2X9xSXZ3Vl/u+xGJY+eB6/odtf8Fd+WiRGci4R5E1P5ejBhrYZZyNxyRSSI
QkNZaXJUkDlvzzg4Ozknz5xXXn/9BAtF2wh3B2uwbt4HFmIsPIK6LJ++WMjk
pWeOmStIZM7KqEisE+xBJhCDs6+ILJLdvfs9+3qIp2YMpq6XrCFB3EwFBqwt
5yi7Wotz6Ib9+4p/2tWIR4TKERP+M16Y/RLxBjTrhUm7K5rtiGhRyXbWrQ01
U5IZnNEGiP6jFlpohLcHY3i0jDc7RzXmrotCcJ81E+pfcGyq/i70T9QNwWWj
xIvKxpa6AMRXgYdnD2dxWp/6TEJvDESuacgNjj1SVlDcChRcbLoNu/Q7UYrt
QlbKWFqGJ2Yiuu621ybvTGMpJWoH7dWeJbEveYlnMPdqS8mh/O9UnAjMgt3f
T4H2m/v7PsdEeVmnwFnUaiYnm96EBSgsqXjwYihVk8TjEwENb2HLaQW2ZeTT
0SqDtyP44SqJPfHjjoICA54c3/A4CJxS30s+TEtmkIYlRZ4BjDhBaDkYZP1r
k0H6i9rHJx/TGO5w76aneLVeOu0ZwkUrP3RuPS5IslFyULkeOTQ/H6zFi+S2
miltUFTzP02ktGDEUZZ3GLK0HnwlrcYzmAiCJDi4Yz30+Bz78BuxcXnKKpQH
xVauuBHRiuWN6AIIgsSFwQAgTcWHQIwYxnbBtLh/rjsqxnTe8MGCwptyofKR
ZPbY8yvg57EVyrtwo9l6D2BKMzOmpvAhSUqmAkyvHW4FjGQ0T9eyZIGiZV0c
lbhyGX4JFnUeprytOAf54ueuzQtenax5iW21pSxnhKqjpd9vKg0yszpsNopC
NWkACDU2gz21LlOjWOZYUsxef+BYS3LhGuQwVCIdCTCZeL7P9U9xTyyQFwlm
Y02f9TliTXcAehO/PluUBuaSugplpUddVrz40XeWbrOz9+Y64i176V3Q3N1I
eF+z+H1Y6Z9p6d4N23rT9Is7oNx8kqaNSVkJvSL3QQ+DEP8vUrtvfteuf4Fg
3lH/SmlgokH0JZleZ2FkmY6c/P+9lMrn0GeoQ265A+WosLHfrOLEnTtGK1uI
WZOq0HrmrWUy5LND4AQi+l8RmqrZl8hzQh4ndLo7BYPd+UhLbS9a4+lWuvVk
yn1edb9b+b8Lb6764EtsY3pnYy/Dh4Llq5fS1TjcD7DawocDYl+1TTktUdzq
zWJclAolfWSDvTnFfNhq/n5vfIlRcSlYJID885GAg+WHc6OTqOldRo7cgev2
iylfDr5q5KN/aW1TCMigHhLPbUyNN6+7ghZTi9z2oLo1KEjfW3zqd3y5UxwV
Jtf9WT3UcP00aLNW+QKXme/fYxDAtRrvsQeDwFTJeSgrQFmUq4tr4vGgoUw8
Do7RF7JDK2DXVfxEVUocAAQW/M4hz5nco49NIcK9RLzptAVRHo1FSQDFfAPi
Zb3LDHIwYS6d2Ej7exd1z6giGTxsqL0BEjh5VOSN1H27EA7tCt38OwNvS8OV
cCL53bx7FrSPD+q46/eoHfSfRj/QCdhbZmlyOq2nB8Cxq4QGzJEG2cSxTdBj
JOvFO4OuLMXz+ChrtUflwmNDwgrRnkyShLKwi1FfTBRkg4YKXGZUd7TTtivV
bzTqibrPRi2Os4MPEcotDyWTP8qFpRjyVZR/WZsK4rjWlXQZqgLWcXvIqN3a
w56JqS4fzfdB+qkxdGJT6nBleIwxCORcTabkAZeFndMeN2j/PFzElM4vT4HN
Z9/xoKyDArhj1I6LdVgqe+kCx67nwLbhcacbbnu2+9n/heVstoUXKlDSHPp3
y4OllP6d7N1WgVLE1YQgU/jrRIK1UZ49w4idVEAgYrktKCZhw3jrN+pnXImq
omdFmRVbGgKHhTjC0HeO8+KMP/tBtSpSPucfbAeRdEUW1aYdGPj8rvWI9ucf
4LkzKlIzJNZbeouOai/nW6UJzi7H2iWshq61tB0CXCGYzElX9IaJErpMxJ9H
oHjj25elEFDXqhJWn2jbU6O0yWUqJNSGT9+Ef8Yug9gb1NHqyLg8UIfBZSvR
CVOUVPgBp5y7jYSaWT6sjPizD+47z6EgG+w+ruAF76+LJwEWNmQID0L09SXF
6fecOOKa7N1cbZdi1w2BpOaGVtVt2ZH5WTm5Gqug1dNcffD07xQRIgFQ1rfc
GV8iLprXYYKhtAUNn39cyg8UFffiIIxKdYbBbJqe2KZjeL3nY5HKFxGfsuAb
H8/3IHkjITHIn1beLrKnch5GTJcDd2WoTxfLUrFt84A4hX8pBGGTAJoImgqT
7HUhJkYL2covb+MC5IwV9EaBVn7CZ6ob+xwdl09/cBXoest5mHwp7SGA+1Kw
K6wVf/FasX+Ebb/w/qpPZr6xj5rV56JmumuhVJYSP0fLXfic3lKqV8YOUpXx
ANbCFFKEw7z6xdG7uKe/UNcqSnW7FBxy8bHK8Eo+bhizmyoXOvAYmzUWGQlb
UrW86eVnRvDA2aVIQ+27NlZ2X01Oxe+1eCpLEBt3iJfN4yzuKNG59lVIqElv
mINt7huIzdheGwjH4j6PVpjD2qOY9/kQ308oi6Ps48ht3Y8+dkYTPckNw5ZA
IkJ3NRWi2o/hBMBBXcdD1KSBw/ETa2NfUgzON1lx3OVkZD/F1qQeu+TfqG6f
a5Vt40iw84JM5KQODQgskOnlQbWlReDvEOxYRzhASEL93+IOsJPx6rRNlKo9
T+lCmx+HEBvdJWjvdwAzZxTFxIWzIwKCyU4V5jGa9dGsaNGgZF5t0cV92BpR
ITRG3kznlV/9e8wiSo1UgHvuvr9AAi6oF7Z4H2yiK1Y8TGbYK421Gxfsju3I
XIoEBEWeySZKS9DSYjwFRZX8WxtiS08QnaRAp+RhdzCLjElIE9Z0GcR4tHcm
BQtmo/HQloFv7OB896pKs/kGCDTi6XJjZetb+zanJxhfsefxJMdAddXR2jJn
23S8CE5EOqcaPptwSfQONBEOSsCvsnIW31x/JPA539tSYomLxUakdx5qWttA
HKDsdDMwPOLM9yggB0j9hlDHCpB6DCINXCcSafyNrt0Qr95bznYw3ggwNIRV
p4ijR7yCyDDP2eMhGGt8bn9bEFQce5m1Ymuo8bs1YEEfgxLF5G0ZEKVteRTW
HdWbqu5VB5PoFfJ7uEOTwo6cQWPj9ckf9p/7jyGPcs/FqLlpqzhpQGb0waBs
1zkLYiHhg2qakpz8xLDXU1NeRmLnmUoh7Yn10fyF4kchfdeFyMCkeLexjEUp
iRN7JfTCxQzh/eb464mFI6p3nNwyGXqYsMZK6Lx3KGU0WIp7PfJcafz5i67N
Kav/hHVeIpdvvkxPR+SkrjE9qFpxajIRLxQw1gHMME1aVy0WVJpBtnNTFA5S
NMXHtezhoOcT0GEkcUpcvYoK3gg4hjNERniO6XIrdcJUqLhwZIlcdwPsNSO2
RDyi8hq0finx81ShbVEIKIpprPaM9Y8WLro7fawrSVrxC7tILMBkCPebCmoR
6Mu4sgVxGOW31RUjubRU7jz6RcLGHlg/GQhWsuA5t0OzpwxTVC1gGkz+eRb3
f59M1jPA9bd073V8oU4uzFagW6WyPGxT3WYkL6CkR8zkM405qo+XF+GbAcS7
pgizkOUmQ1wy9PTPc4Q90QqRQ8WeCNuqc4pVMaXf4fMjGnMQtSwKBCfjufZg
t4sWwlo6qUulyT43sjSULrPizjNsrpc3zk2Qad98+Blu1nWXL9xm0hMVdtJW
3ug1nFDv/PO722vpzxqO51fC38y7uD0i/d8cZljt12Wa2LHD2QVjPn4iZvQx
R2bUsId2lxCnzI5G2gkev864+wjuWbPz9nwhU4tue5sDDAERNGX1ZRGaQ0C5
3jWj0NJX0mhrtU9ABkWqeo/6NnosFzakBVItiXmM4vU3zmHBIEIhDCwDndOC
Iyb10pQadPHn3vGAbTV89e0pHwKnweAzAuc1sT7DbdO2qxcD3doXOGzLrWYD
q1rQUibGVMybyupL0Wj0Jf8RyWqcAAQtD02o69zrwjT3MF3qVcmFAYatI0qg
ZchRomDcng/6EP4tECYAxyj3uJnx1wDxmx26gyNc1wrU/m/5uaCg/cjE6UQg
sZ+Ao2R23CAuXNJv+I4UIRY2KR4kWYnuzZzY7WKncA1qAtFvXtQyDsiNCufA
wsUf/QNJOAqtJGqmg2uQAFKiRb2EjGRkgbee+1DMrT8WnJgccvtaI+Oj0IYi
JZf8sIZuu2B73Sa0UorPnachPbGuNqblvvJknxmJ4tQzIhI3mkp0EtQsC4lf
H/xmVtYope2o2DR6UUIG9HvccalbNC1LScaqB3mbllGPgldKgI8mDFwShSJT
Xv/I4VvT8xDBTcUvyZm5GQJSyjviebedR9PfQKpxIak+VoBHqKpFw+XJK3og
icRn6CkWt8GXgZ5gBfSLiM+INxkiN9btyVXa8MfoDqlXHWrcPDNRTKVfi7h5
BzSmjSkMa7ZYPFpwxMVjwYmMWZnOm/8469tV3sUMo9e0zjxRt19OCXOwpSLr
5WD1mTxVE+ubhXb42Ig4udBRZYsuMUF/RiLz5ovJVypbcIkhwOmfKSaUikDn
szbFjMShNi0ZfWakD6mRjjOUEhbhAvi3B6jq31ypQDzFOw0EFSNGkLUIfva7
M7BVbwHudA+kzJzy4os+mnp17mhOs7YHQ8iL9QW9x+FWH3g3uuTWUVwgl4TV
nuvn3+gcaaYroksaIe6SAI03wb04GDnyD0FZ+inurvp1C+Rk8IOxAPHN9lsB
LI/T8I3rpLWJjAy/9H30yFYHuNTrjCbPUTrd1cRYRvsWZWEiDSL1PUilNf+U
SDZd4qNkfrz/f9cVjTc8IF4z4CJiPqhj4/8doYoWg+yEyucB8PufjQS/5bti
xj5PBfb4uj+Xb6t5SApAzJv49tiLQW11XCF9PrBRu5U9gWzfBJHjJa5/J54w
yEBwFlax4GQZyNEEVYktVwelpyXvI+D9rXsb5MXWYJKxcFkI/OUjj7VkEiY0
S+4RRSUgvRdU7Zg3yEnXskPk+QzpJ+UaVsvO8fwAl/EfxvcF0zHZ7PQG1uEX
P6Yk2s7UQ5RzXHjnMnHU/XKxdrADcbkl3eMVh/Q0upjR1Ghf7G970IeW3N0F
L5lLW9A4JTgOPRdpzRkxoMRdxVYJW5+7eJFGddN2zf6wTAk1ULQl1PkY5BlI
FygiIj2uZDYxHBx5qG3TPTHo1pJYXcAbbOrngqFj6y/rFtoWS3Fg/MB2z41g
7HA+AOZVPjzVsgZaAMXXyeJF7Zd1al4RQAcYj0lCGQuXipZC9D2vNGMTJy3C
ynaloyz1OOpZp5j7Kfu8cSQtRYGaZhzQ2Oa56xMVlePBw/E2ScfLQ7TujqfD
IvSD5hSVKVN3CnteZxjQcfXDnqpgrbCAeqKJLn4zpnsCgtnouGqi003NMTWg
LWhis7gsPvCkrfqvwXSqkRC8SYO3ACCTgtkyc6x5Qk2gJrGUjiNiLPrSdMpa
7rYnuxkMe9JEnvd/0Ppk1l8t8cWNXHd2dk1h03+gTN9nNvraJJ5tniBNBThu
Ye4HNGfxswLBd1fGcsxsX/gnXIYM5X5ykxqwER9OU/+n/kE+APETdaB8nsdH
KH4Vu7F2uNssThZZOFUkFADGD95F+iTlnbfzHdYpSuH96AfCjJVyx5cz0SA4
B2nVEghYhAgVXaEigbqhTT0PWclfX677n5Tf9WoB1U4CfbJ91OBV/xlmJCQH
2beQhLuqs6QC5dJ7iKrCf+ZCCgM0WdNMuefhLyCCXyVK9jzF+TOZKe9WWD6S
umJmN6kvBksJG3A/TLR0Spoh3KPCKW9INUx0GAcxtK74I4cAcgD4wtrGG6uE
UygR7jUj5fL80YxBOjwXn2fFdvDyQzlQv1iCWEzwCHTy3MvrqG+nNg7huE4d
OIBdM8n9/hkJZ1INi9GSaD2nbU791upSb+rKPhnt6a1waqVOFITXt8jaGqJS
Wn8d3jfQB4AtmorQTd/NFgmoJ+k8BxQzPHHeKXZFOSEb4EcHpzCRaqWaHfnA
tfV2/1JTWk7GzZpniZhjpgK3oRplG8MzSJseDv4ZKRDbX39ISdoqnH1i27tK
CQRpoJIA2QVT2shroiUU3RQf2ODh75OCLUMk+PwRyfyytSAUMjffKWhlsAuB
WLtQ/s3LNmsgV9wd3mLlBXdeiR/l5w5P3Uqcd34YGAmeL/19ohRe41ET3T4l
406sBuLgeFOUrArl3mgpYQLt/Huv19lIAziECOqhU3auw1WLgDd46NeWuEki
q2X8vGNTr4i7+rlxpY/bG9FgJrtBLthxgEEsYGHIz1ncfYtPMCxiP+7Z8tK6
JcyES+oSd/tPaKFn4NXKV5qJ/YbEGeuWDudzoh8wfhREaH0ZEJMjSxEH2fb5
6wyfxTBwbBY8N/U+p2TuP01mJP18K74IBPfH+uuXxgGASfKScBtgT7UjBIBB
uDXpbIAJHSGxSoP/TqOXE7QP4SH1ELkdYNj3zmkzFS+j6qyNDYzvNWexZri8
dCeM2x/c6R2Izee+TfPc5wH+YExElFf0oImPdz5jXGxD8oR6DoDo76wz45lT
yBfbGvE/emZBE3Epe2fYIXFxM1Ow8ALVaqfqXg2jx2OOEfEdz99l/3Sjd34r
VYqedq6EhrIjuWxg2LWdF1FuBCnBc1wSiX1j914AYvl/EcGjUUVK4r+0KM3a
9NV+n5AW+Zy7AIiWNM/WxrdqGHGppdEzZ7JNp1HuE7THcRslyAFI6UTA+QT5
l+RbfMKU2ONY4l/7AylHb0VQV56fPnjCqYuJohYPZIXnYad5wvuCknJHf6oq
2qtQKdAgKMnWNyTaiQGRcGNIuZVmaAfN2ShoFOxb5Eg18g2/k7TYVyJx3oVS
54dBtejfgAxugs+d7qY8cJthX3twmB/2NsrBoUzKkyj9b66KBoVnD2bueYh6
zNp0MwWzHk1XOw0DpP6Xcbmnzn1dWxVAI8TFd8xCdChsn+7NmXQsdZJlUj3g
1LbdUUqI5uWJQr9CY8q7LXOgTUp/50t6LFawc1vZEtHP1QZTX23e6f2R2YTZ
ULfTq8Qb7cXo3sRUjwz/eAIYlPBUpFsv87RPmyPx58PwHrxn8cc1JERrm13n
N85+YBOxcOmwCC2R6kFSk3Fr3Ib6iG3K9WOzClQVt7OM2QDqR1GJ1Gq8oPjZ
C8NJNjZSYtpemkoSliFfi8dFbl1einlxX9eylx630eryKYsPbtGz1sB7ii22
Wb0y6SyNQ+haaB0S4xnFx/TGpYPUZs7bve9VJkugbIIQkHMj5DWiQ1KGi5Zz
DVpIb+PsZI3J45R3/k3c5jD0XGj8V+OrlOP6VmPu/Sd+In+L80+o8AO3S8OW
XQu7sL7GXVmyVMs10eJJWPqNW5E0RwSgZX+Yqdo2K8V85KXY/G8TTAr6T+73
iW0jeS6pyqcXd7uxJ5rgfJYnjaZoAxXIjDOhY0B5BFAGnBhU2stylJ3TD8x9
CLSGiuhvLmkDimgCwelUr5Pe3KtjiPS3+MqA2wxpAOJpXBPeGsf1khIcUpal
qnyz/yDQqxCEv8/7dr+13Oi7vGKd+HjxiNMpdJiObB9UEM50Fl2ir8bWSXBV
mDDKIlEMlh+B+i5R50TdEuTO9GAe96F780Mz3YlKlyJF0WImRASJ3nRhmNdq
kisejPqdfjIuffldGYcBesFoSiENpVTUMmRu9J+2aoTR9KAmmULmPjjP5TIh
v5HZFyPuSzAzJPV7Z4el3OOiVTAAR/PrZA0HZIJW6uPsGjebYGgY5T8RzR5k
Y0Ffn7T0SuZd3g+hYhiO4moed+D5jalnLvixsQmsIiK71FyzXVd5habdx2xw
HLhD5xCXoxJyRNLAE2V0HmnPcZ1zNhPdTsgjiBb583nJlYOOIqFxTgRZIdpe
JtYWE1MID1hZZ0XfzZfjFwNYtEjifjAkmfY1MXDVbfrWnfllsOl1pUW4zD2i
mL2zBy8hjzjTpJSTheWfS9rJDUOcMYUOWKoNUHeAuGy57FjPS0HtR5zHfAfu
duoGJ6OqJTajBzJGYwmJX2h9Q4lrXv8hPbKCIxB8IJzZtfgJc7E21uBtSIJN
gnU+CoQn9I5bAWo4qxmWriTsqRLYRd47plPFiv5SPdF5ES2ILwEDMaTeGr9L
5blRLDLTfGZ+mhfhL7OxMy1+V62IFGau1/gUDMpxHputwW7x3l6IjE4fPlpp
frm0KruwgXZ4ux6V3uziQ7XIDb1XBD60c11MdX14DaYkCdm+vQe2Ae9jMxpA
sckYLu9NHpUgbvqKu0RPiM3u7q2zN+mDHiFh3Z+Avh0lU2j+cPdSGZXfdc0P
hKisBC73ipyO54fx0gKPaGF9PMEa+52tfPLxyQfWQKasoxNCVIw9U8LBuA9j
rjteWxuOwBO8nWvhdSoov8th/w+YVCibF75xISUOtSV5XeGZWhSkKKfNxtN0
atanuFQO2DG6d8J9zC3KcEGUSeM1YJkKrVqUidLZaXkzBADZIREYPMkOxwS+
F7ubbqnPTshoblJoqv/q1FLDf+IGyk6KRbXdXmIumTZSoz1ONyeY+A5tQxR+
zur2QdA6ANbHPkBm8RBd7gQeJXwmZsj93RxIbgpJxYPWQzO+jfmwixwglewY
qkxqAEZPnGS8UaRkeF17D53NNV37vEgwCQLMpIh0Afhr7/4f1jewTa/zSpn4
LI2LavA+aFnhwX+unPRhCu2QutdtUO09HX6oyEq/3go5Bc6vrN9fXwISGUpG
fW/w54gO/yjnAfoUTsODLgz+xkBCn+ywWl7+7Mpng5i5ZkYrRE7lv2u+Z/OJ
r734hZfThLipcoEtt8DBTaAfMZwtLUJXrL1znio8hu/lcqauy4+affSByN8v
fx1b5cnWGRmUmfDzSl+pC83UyiNnyGEQ+LMCFxlW1MG9lUyj4uSYzdrh5Lzo
9v9AaJWGWQtfxWlqbeZVPKNZo6Bp9PNp9gIn9zzgu6dx62WltQRpSZ/Ikmgr
anz10a9P9DGlY4sgBaIw3Dhx3fgnQUzK0MP36mAW+ute4DW1DjAqZwXHFIsA
M1UGkha2HfTWIkEAhScx7b+IB0iz4OFg0itHQQ5TmcG6oDJARvO/V/n6/KA9
GwReS33Ykikf0WVDCUQY9DEkazqBPc+ep/NCHIDeyxX8MxD8Nc4oV80p6tI9
QNAqTMyzDpJDrjxqroGsTnifggFLZ9RTQ5xxqARLAujuMS43ve7fQJshA1QD
jZtnqidyz8PFLJPaVF2mWpbGQzG1mANIiIUEB4rj+LEXbQuAyTYT66Ocjyo5
GnH62NL5r+5GvR7kBw5j5Khp5zOmKUVTOmhY7dBPTMk1vsA9kph7LMITFOgc
u/lBV5pWA75lsPpmcDey2YXB7yZxSuXQfsGiuVwCW4Mex3iBR2rpxbgfyLYd
Ml/mimBWYBBB3tnmyEwR1+1anZnFT5uRTxEHV2psn3o4QQdqeo7BP1u8O6pr
Z4zd2C1dQWSyJwbuIsxpgw2N8E9BJKnmEZrMDuRnYxuw3XLlRe0LjIwHfv64
tDww7nD3kUQPllMUqUm8jW+bNwUoTt46kiGEsZk1s2925b46tP/tTuJpElI2
3jJt8IM5F6HXnZiA1o2veegk7qmI/wf9LIPgJfAnYXfgJ+rLD+Y8KMR7PFKt
Blf8TvU4mGWLJbFW2YzA+zFfbJCG0W/6dPHROmQCv2Bt2VMnChYO5zVkwLOf
Y7saczofGsQsfEYs80z0PgV+qectBfkKvsDulXir1UhNoXN732lih3ZWzWCS
fg/byqprwZDPKY2VwhIxjEWVovk6Tcooo5AmGKKk++mJZeOTb4E86iWR63U6
sCC4A+TYwJ7lPX1J1HW/LgiJTI3PDImBC7ZIw8rvVtIYZk7kQqcUVPNCgoJT
xp63RCFqX2B3QMN4ZwEkSrf1sJhndv8eIaf9h7E9RYbpCi7o82MFUuSKsMJw
Xk3G5bMFFHsaympL7N5paMcOWAnWziVonk0tb8CPPjBYpdx9XMsFdaXYAqyE
TogvbnNMW4UScvlaQPYJMFc5xVKZTsnMCx0s4Y8OrQbIxSnyUs4e4/2aEz5F
sVkR6PGmzt4sM0OTKzn4euAC/YrgAUH8AjDVKnof9u9FwT2uz3l5N8xJNwpy
GAb/RxnNsAtWUIG8EVyE37JoTes2vKxFVbjASybFshiENdfTmQ1OgHw6PKtt
NnxTKr/A3PIaqfYnVOwm+rWM4dDNbZGPIwt7GQ1Zwde90Qpl5T6Cume5XCQM
CgUP+dXxBBFqy93UeizBfSY+xyKH1GR9ptse5i8IKjnnc1yUvEVXX83wj1l0
jFWbia0lvyFK6T++srCUYQ9Sg6QWCSgmlCa2aDf03fOK8Whji+giuTCx2Kiw
O7PSVjqL9eq4tJUDnUqE/M2GRD+DLZY7iD9clppoODRFTYfL/IV++e2WFUrj
PVgaqh5BOPd935dq3dvGnZkbNrm1pqdrztiPM3hg2Vaqdvcj77eNcI+q4ot7
Go8wL6sTluSDhmzYixxzAOy08HO1HcGGxodADhI6PQRe0LJJbA0+ckmdGHqI
aIKyEewmHTEjhwo9XIDXTde+oKJfJry62mZ5gEWcSnSDlPrMpIgR3uVkKFqY
VbxhaaO07XYGQ9+wdHN6INrP4H/4tWVpQ9Y+ZEvN4OHBmZoeMq49wkCdTRRa
1121Xaow7RxSQvn77hsqWTCbpi8iqOD6t3TxqGDPlW00rBcYuSa+H5vSsv8Q
x91Q8+im53qVD3ZzkKvCmqMlIoECHb0OmYN9+xO9k6K3Wh0LDKOhJDEu020U
weWni0G2WTwWweh0DSEFjGEndyx9dKPZG3XJ0DYsm9lUba7KJBP0gZ6V4GoH
WE541OIefCxUO/JfLv2rOS2Dym3lh2+LGxvZB+zJlBbR47EIeUp0SOfcKzpf
N+EE4f0IH8RuwIUOUrzuCQG9KpC4JKJRpgtjseVMSIZoU6wejUwrfKJFa4xZ
4S4/oKwNmq3LAM60xuu6s22FGt780t4MfM9Cwk1TCoHWtXl+JcsH9jIB8QDQ
fJff9ifJb3yDjkYXKgQ4UHXtwk7rUIQG/dkxosbc/k0YEasjUEi28qLJokTo
ofERXskeKl96OTVV7SKutMfCfU4hDI2Q4/OE/QWvSNAkRJ7OUy5k1sWerYYH
zZKLitrh/VLdSJgVDz0tHvtQhFCuEmW9G7AKbuTFSf8m8iq2MUZ8/5akugtc
6JCVJ3VjHt4PKxd25NBZtpJBso2Fl4MBr9jF3/NkgKhC/CKfiWPfehbChrOJ
6eWY+DZyObcOAi6FrPZsoCIE9XyZok9ieKOmPSLUncJnUUEMNGO9V2D3FwwG
A6/Q1+XvmmMhqvMzbhmrqNMxL0mRX1LDkTeoDrV9VO5wnszSHGIkNi/UGw1+
+y5DPP71Jcgtpvr+OltS2cS2/DHIUFkqDDhkCenqqF8RbzhMz91PPGXPhX7R
Gjyoo+bYDNI8FMopVQAV2c6B3PiETrBLNrZZI66i43YaxO38YigJ7PT2ENae
rVlI+PXX59qwtKOi5KJVaVyZbGZZFdpEDPCZaCvPj4xuv6HBQbUnh9g60/kF
LMykoZV0f9JrdZmc2AGNLDOzd+CIJ4QDA/wDF8v+9Wfbhvi7f6LRu62JaS7V
ZRuyQS75hGHsz7y44yFHiGQ9sqL2+M7+5NCwhtZ0AZBvUt+CbLej9YbViVd7
8VdrOl3ulPmvqx8Ewz8iWDjo8C1AQrh/xwbqspKPGeUxX4q/4jdlGiItMdMM
esR3sDilXKHcurTuAWOWOBaYV7yx4wkyqNrp/cjh3rJdqYzxAwenBpmJiRlR
vrPp95jg9ncABLkZcn0+tI5/uPRfUKRmfbAhf80hZy+Cq7QEWR8msqVrXwe5
9XssGYY5ym6fJJIxuPgcieoh4cQQmASFfdI1StrJJM2gUpUH6TRnQGy9bTHR
1kE6AWofZY8eKODkafEQdlD5YdIXB+Zb2vu9RVaxgQldPW93eiB4xXzEThGs
QBrAESdOIBGSUIdeTeIuRJTG/OTTwAPucFiwyPRl6M0DBO8Ozih8XAUk2WzF
cfWnsVS//tegNdNngtSbfg5t0AQzHaC+b5IpBGAQJ3S7CZFLF2FDXXiwJM8E
FVYVsHry5BFPVgSDLYh/Zo1KpdS7/wgQbqG9PPkXB9xbLcO7vY9OMe0oPtH/
59mbUiVBUy21eu1PAU5eHlJrwm11720CsHnjSg6kyyq31mQgsp2gtUvDxq6E
bsnFe5IYQdyT6XDzx7DN6vDUtdOxiKux2QHizP+JwHzGPYgC2Ov+tlepQ6nI
4ubXpUNgUaDke88MZRf1KSpxzyfwthgUcsd0iGluYmmQZ4qsohyqcIQKlZ27
+vZAMYcRhzDbbOzgmHgLMjM7J3aUe+nUquhUWCfh5hUsU13hWtc7fB3Rn6fV
BTauVdXT+L7rGNAReWf2jaC1iAebB7mMyHqcc1nV1oOpdqIPM+M2bWLWbjWl
Dt+KPnq/3UzP0dKc2ZqIiZbMkwKrzoBeO1qa2fYiwL3qPbWcZT2YfunkV0wq
wggPK7sgwyglcoy2LM6PrXqEbHCgawd1cMNLwoZSNEaRorVJamvv8d8n3cby
kFI5ewMkuUGI9RyFyI/ZFruUFgpr+jwZLYs1fKSiw7xceuIEqoZo51tYFUXd
kY+q0VXEiLaC781OZhxEMa4ov+k/KPi1Xl1oU+kKYWIQEJITAy5r5DCcW4KH
TW2pELQZyZ7psE6+L+43JSWEKPqANWF2oqVXI8vUtdDwxD3CNsZ+hV7z2U0L
cher+Jy01DWRDaRjw8qeblSaquurBi0mSibhXRTX7DcAZrRx18YwykaYgblt
764n6LxX6dAljzLr7jKpSL1EDGvmeL4F71DcTse8CnFIZX4npJw3OpnKxmFX
rFacXy3WyKJQUHHNA2FhQHN52CeUVXjebA74138bmQ/8axfxxgd01NVgcJXU
MipMiBABO3B2qV5vgZEJQXLRcfC0FVLlLAR9GZ154IsrD54bQL4MWIEo3qV1
CYkaos8jXsb38hwz+vJZ9stmh4mouSDnOwiB1pD0ButBUphChwv2l8DcYd9d
s20rJZpiAACT+LpMpVDjY6XeD4HotNM3BMoZFyhMjKEJMtk7yec6jaE2uy/g
7SsRzOOLEn2KP0sAmnSu5W3iS5LuW1uN8eMaVQdTg49lGcOmPP5dFxhhjuKW
Dk/0+k+0kH3XyqN0WIHsd7d4KjY05OAtxCtcOaZEsjX2Y83jhMUcjtzu3cFO
oBakVBUEVGNLfnGktBdMl2/Q1f89lQ1ZBPmGXztMr5KDTgkIlDu9MwP2uKXN
h5CUvn5vRCs5KKlRg053pZhPnQzz+F4+JjkDu+jxMwnAVjrI8W9mfPAsuMke
lVBkHNf/FtPEDbx2BeL1m5X8CEs3rK9SjMsTd2eFYAuJB4Tg3xEWjqZxGXHq
2Kiu4Ec/Xg0SLINJUtCnjwmpI3u2r/UFZmzlIfT1gtYFoj4BszPCDiY7OCrH
clCOkdlJkZNroW+BWB/We4HMCaUTS7kyJNKmXwfpDwL7ImeaIkys/FX030Ba
VJYJSnOLoMMhfQXBAva/2o8P9wLWCIBrerqFbwCqi0eKd+89FGIhuYG87Vr+
Hok3fl1BU1IW18sXyC9I2BY6tGkNQ0EOQJtkrpYaDCXpnVln6FyM5tknyLq4
DC9TIfdKKGY3MJ8UuLNniPhNeGINpW+65bediPtybBdYwvp/V6RGkzRxL6j3
II4UL+kh0BiV6R+xw4E3EnH0w2M5xNLK9Dmn6XpYmMrf2OBqo1lsBM2YYURN
BBrCn1SzwcA1U0yX7SgJ79riJ2qZhnYbXNGst5/fnAscReUXON3uHukfrpwb
74khXI6zRqAhJ4Jx5vA4UT/XUS4a9sUhY2XCCgpObzTT5xnLZ766NII2GRt2
go0BOJ5fnqDEC6XzNjsHvTjOfGiJmIFfhg4B08pxG6Vec5buuDK4Cex9Grq1
qpLfoCK75IG4FLoD1HVkj1w549WhWFqG5wqEY9Vk9Zxnv4nO/yRZZUTXswFT
hgl+C753o4T3YOkCweX6k7yNEoWQOl+GjEu4JBbX+WGMWdlLBM6wDAXnt1JP
TAtJwDtZjyASLvIVKUnHtLJZtFyidGnjsfQFuC8+7hS2QEoNC0JH9OwGmRTw
fG8Z71Wdd2BkCvRlvZ2I/NL+RrnqKLZMRZdqE6e2WKvmhjGIoYQXcnpH5umA
6SrQllkTupNlo4QfujoMF/qQvJhWrXZP9YYbTfjNX1jZxvq2IpNyb45JnHmO
bcqtD71jqND/x52YWnPRIW9amGdJd7GIVoIPQEUeDGWpTUM1uVf2vrdIUYZu
jUn3GEAZypuLxIrS/YfscolG+nxvuXT4szmOzu9DC+yFoLHMuu+/VOnU6YDd
bBhbS1w4v+r9tzxY2/s1TIftpUqSccvgIsJL+9dgX+Vq/oRPVyzmGAQC0THs
VPSPRCub0gWA5U2FWT9gn9gpyP7q/FQxz8xAXO8+IP4I+VpWxfJuGCSBHIeR
Pbnq2eLqO3tymsaDEFEAo+1LGdweNw8UDFKC5a2KOwUXXpByRLyGE/K/QLfx
VXHq8BvB+0DDhuNEuxj4Ko7W1XwlEfOxZZeOEZLI4UQv4HeLKDUJOQ0at4/J
R2sQE3hyQ6jFDPtr3QKwZQkZZ0WcIVkdHQxOiK7GiOlGCvMVquepc7E0Ijt+
AtBQcu4SPS2ygUFTNvp3Y5Y1swUM9vNGH3S2a3m3/WxpgYENf49U2Dujvzt+
BdpY0n2fZpdI81MtZcB4PmSORbTunMvlMX7EbulIQ6qtGiBpoRb00rt8O/2+
ELIhBxTI5XPoFN74COZb5cKjD6RU/v6gWwQZx/GZR925x3Ho4ay9PA/+WZQS
N3hxifWz9ThDyNHapZBMqzqwvl9vadpoQQJkLYJncmUDcdlTHYwdrG60K75B
DtvZwJR+RG5ZUj0S/E0wyK5latRTlshU7gVfxBHDaAjf31GNkl0mRQgDXkZv
u3ClKoWmypA1/cuan+AmI5I0SCUPi3bWLzuhL9qcrnssNk2unU7ej+b0xlvV
vCk15Gqi1pKBitSzvO2xX3rW8ix8d9UjSmNL4x9DC0ngyvgoARLSXp6S3v79
R7eZo+OfjNTOx+nlsNmWwn117+2V60SbFqAdQ2eyEE6p+dgyWTMpVdpRl03x
Q4LUZXiag8X6UbjQxj85k6C3aPTuAb09pazzPFJBY89c8b7BsFmYrbcQ3VO2
lnasI+lR/ZXqld/3Jn2V4cMyckYzhIpglPm0FCPS3CzsEXiyPfMbIedUAa3v
fhRlHvlQvbmskHl9ObmBlnWpZyIlsBQW5HoOOaL/44SvI/WIMMWl71DlWMZx
PHeQ4vPerSg703xU7YPIhjjzLLLBCA9B1oGxvGyrgVTjwDfa8uwOWHys12NW
F+OeGcxbO11x36ce+f8fiSJtoesVw5Lwqjdizdj/7kye5uadoRcF9z8NGf6K
vehTQagvB/1iS07yfSo6r7/10BSNni0IZ5AH1PiRBPtidxcJX0QDvH9LHMdx
DQSs433fHKK60w+sjGUOkn98hHJSBJ4qjwUEWZo3iwRaCkpap099bqBvTrG0
5WDUuICMZlBvPH1/CAXqhIP97LzidjXSMH/I9XU+9ocfSk6a0rjXNcTEt8+k
5H0IGOBofdZsNoMZX/2edmzW/ziDrS+slf5rMkxRshhtIm/MxC+44+VuisSA
xqCxlg3tkz3FlaKgmhG2ih1WRn70YSgs7TAWNhEjJxpugfpHUKEQd0NPZPdl
x8+fVsqsGBdFksLG/hntPzm+6LbPLnmLvoNyUXiilO3eOlOWanS4YWG/QSAA
2y81DDzUXG1f5qlTPtxpIrFz+9qcl5mxfexrHR5QOgDCSiQlb5E13hHM1K+e
a0mGUk+LSrjBBSkeifGryA03Vn7Hg7gP/G/6b9JbXG2h34C/nZ5zBTFigbgD
E+rcJ2+K3OA31LTVG0ytHLvsXD1ezsXjSyz3e5Nzmr0GtJ8dUNfva4u/Nx9L
im8ljFzZgWDnjyt96ElmjVCqvQoDTXPjxHztVowgxpBcB9QtMvMG/MRXkMVu
JBhbbTRuDM+H5HQoP+J7GxKG+m8wVOq18pSmwKmEw3B2qesRXoMxyZa1lPWk
EZDm01Sj1uay9cgcuHluUrvqeGapUkpBKJgpXCFqFaJWr7T7Y6lzf995V4N3
Ms6Mg9uH4aPLVvNUaG8HtvybYIIi7fDU6XfM5Cx/XQsT+AdeSH3FMBvoLNpy
EVDWDUiKsigpyfZPitD0jrpQQS1egGeo8e8ozugthtHXfWhTngGmHSjSbofC
KiJIu3xogIma55keTrtO0h4q8xr4Xh4tqtp70PhYhb4PmhJDR2+q2JiJJyij
f11pu9VLAuDX8aXFNvmUNe5cWjeBExW6Cz7wkqq5ROUj64LAUmLwbhtxFG/9
DZiqnl32zPi9rmABz1FBhsT/MSfEI8RKpL3Vno5lLoISE1U3C5idZnh6J1t7
Gooh9ZZ4OhhYBIUIvkrMaYYzIhg/p6Fp8hGxnfco4bpfhfmiKR3cyzrUQm25
OpVg8RSIgdollfJntvpK7mgONp2JOmjksIkecpjaTAjW3lljzZiNbUV4iTkH
sIwPZBCerrlzBV+4X/8ppsmNpzu6FAyPE1v0e6MLq3GXM+tnHj1nq7FjGdRu
qVHFi2P0FaTD5vEtrj4BNxS7E1V6H+Y0sPkA0TNveAgSlGd0zNaPd7TQhrMB
liL7+A/5tdj7/EXRnw4z335ZONVGdfWeV/6kc7WzbDMjk/5+WyPRg/P5e+PI
SJUO2VaqcpYqK33HZEb2LB55g6s/W9mxY2A3D4iEfmv27ztFJU2kb2LvtTG6
w7uj5bhkOAlxjTSz9NVG/SCwR9onj1rjHvA0UL8i8hCq/d1fK0bHatzpUtoc
tcdgWYuXTdKaOI5Axi3J3yJlRjEg4idRDFnvxs6vfnz+izEXVS0sSyK0o6cQ
3Lv/sUiQenOmJQ3cPaHay1fWx6FNrRb+wNDNGJhQZfh6Fv1XGDZloUVdErc5
6bjDe8q1fLEz+eTY3B0tXR/cdMBlnTLgwejzCrWK7U6FN05gueKx5Px9mj1/
L6WAVMq0pbeyN/t5xbDex61QgXSTe9oU9OS8WTxXfa4nHhxtOc8oZe1UuKeX
q/ZlKNhG7CqxYEhiO8OXALrdqNfbi55GKD4OF0Ue+rECsovdIF7SKfiVMJTN
e1nqFEOHkAAcIshYlt9ACQgxLzElBti/Sj7nwi55hE2dLdrT8z5kYPCQGccU
k0mcHyPWlSrQ2l0X5gx2LWY4r6vzgfSzg7ZV4GTOwzZKAI7ZyLjmAFQcRlyp
VJlKRW7+9XB0oulrw05IZQkkJGVreTsyS5puHKeeHzcbWG1B/KWHYVCkVhij
r/EnFFWSllJ5VS9wqZZOL1QznR4fmb7LxTiu++ltPowKI5gp71dZW/FbaJF7
HvVafAHwPhv+HwyythF/hX7DTF70HvoSWuW+U0os4BJSHAJlfOt3YvKHyEUS
gReIk16Hd9afYPR4I76/DFoivJFHpzsVGBN2wOLgBdVWOA7tbfo90caRoEEd
WpvFFg9S3jGH4qfXfUd7exY3G+zfl0yzF40eHURjF4RRziJQOfJMpIQnPvKk
Bqak69+QgOe6BEl8DRyQ933aJcuthQVcregU4qjEe4ARUC51nAEMu8fNGUcq
QKh3MOM+KVzOp8jLV+CMnM/s2dHwsg0O99O/gLzjSxGIM640aVXG5SrwFxPf
W5f5Fx8zOsdU+p2sG1R/IXAipqxJM8URAwJj9gOZ+y5k6+BwJw6HAx1W4PcI
0ohwTWCMO/yOuZcp5o/g6oMWI5kwt+mdP5xExKGhlfoMDIbxqE3K4iS68R+0
ejAGJGdeVGpLHH5muhWiDLqbFoAjoDeCG0yxIJWu3HgThpmM0QO1du3SqH6h
aDmq9MG4Xk7MNTKC4R4dCB1OXJTOJobRnwk8Mexyd376Z3N7pQx00CylETnZ
5TlF9I8FDrDCNHpqM4ZgGqCQVNfFvDz1g5YE/6+imOngCqsh4KL9K2KStzpo
0zXGReN0qMlm6vs45Kv3COjL6dRTO4GjF8E+V3iJrXKek8LY2OHjLv/cLblw
MMJ/otoPXEzjCvvO2W0f+z3nfxhqbGN9UxsGwTFo3cKIBUIAy7PUW+wKQvkc
B8kLLWF3a7JPOsqq5uvA3Sjs4xxlJj3A+CoAazZh7ReSIgZUv8uPFRhHrKUR
GIwZVOzEBnuMTlkGDZzNDs9Qp5Py1MLzvYuxr6QXyZC2Ddly5deaabK5a/aR
rJiBko4zOKdtQCgMUJwfSSB6/B+ixwgJI/6SKgWq/Amzt8dZWhusLiJRRrSq
iCX8ecVv1LSmXU3vnBtPlBTiXrpc3KcJ+dEvIXO6J5MZPTf/+vkRbq/MFaM4
JXuov+N0i04phS5Jv4v7VkpaZuafnxwLvWM9XiE4o69nLwpCmApNnPP9KGgg
u2PLq4TGZH1/UcRgErZ3sK9U+2K2al8MXNJ92HUahpnZeq9k+jh7Ey4j2VoF
wdwPjEniF2bbW+Y+bxlqFjwx87i9Veb0LBkrNQRwrYWXRk33i2RNtrqY78yU
N3sdki5P5kJkQz+s443rC416aWftwdx6LM8UNOQXaw46g9N0fKYmHkkI9HzG
ZGYctnwwE9Bwuc6fHvVfCmSF2eMlj63fbFP06ei6rdvjXikSKZbs8bNOrXQl
BW9yqX36OHGOBPZKkBYK+/9ymPfGgkaZcVWLIpe2UagqOHfBZQZqp4jSp7Ao
D3Rgw9x2wniDIFHaXrEBALc2wSBmKGQ810MS+0DGkpDfCbq5il5mu0xqlbxr
F6Oi8kdMgAJhnwY54+d9LhezgpodjdX1vpS8FraqXSPMwDvj781LoaNNJAL6
Ba3DOXNdZ2idtZoNG9aymCDjmq82f1kWBPZeknqbbFRG16y3CEZntDixi/FW
PQh8Gz60gZRd/jpzNBgYBId/OvzxiguvpAL6I+2eJ/VFtgWs2PF+3jyIISsO
DDM20hqN77nJRZbeQAniDivloW0YOBBitFOkPULv6NXv6nBZF8zkDPc8qTDo
/+lYYASPvJkEffM1mbGIlVmbo0D2+WCeMjccUo1jTHRjXu2aKHk2qThpmjrQ
JKABMVR1CDT/PwoxsjhVBAMnOL9/eCNqLnym4IyT7ttDWsfPNVFwnweFORoK
ycb5Fytuev/qHtnNaQDNfZHXW+ap/zq8ZQUCxjZu1BxfKJoekCDkHyFw7kiz
JlUnNFQj4o+Qj9fZ7PnekbTwqcbVKDis7a75Wxm23ipNLs57Ugha/py92+xE
RRQCTqHnNfyaLARKuUBPXpHH0Nr012S+oDvXEwufQ5Sxba65ck1JK0B3npqT
yvFxvUJdimay77shYw806QBdqCkfTJJnl7H8goRXfXEL7XnKz8zKeJCUw31b
VurxlEz06RLI0h927A7Qjv1dow9QfkcjGexIzgRDbaSRSElWwNao0+NAiOzX
WmRocegJIHO/Tp2jlC17x0MtlKok04mbEdJzkAdxhv61tHBPsn/5B+A9SzKw
0xlkcpxKZP7PIS6vkOHjHGbnxgnoJNHn8VEt8LJXHOtDhEhQBIqE1QRw0fsJ
hJ1D6O3ffLatTDVdkrTfeqN2XqnQjoFFlM6IhdiIH2AKqh+9B06bnY5qvBaP
qrsV6WQRkZ85jYarHNE0u7CdYPC0qLQ/L6rzITLpwE1+Y68z0vEo/1etzLZO
Gsldy1vSMdYBhWaE5OCDa0Mq/XpXuepiA2h9C/TiK7mUfbCs3IIwI9R6J7tJ
qtrXBpyFMUotcBzxnn3dc5PEgPM1RqwcqA2WgpFxkT0rFV6lsXVJn5yATpif
qRjv2cpUrP8msPkAPC3gFDHTlLCyXrJijQs1g0sKtyNbC5TJQ1mhCPRs+l8r
vVbdLfDdTe5C2bi48Q+mbnWU+kJ7bMxl0gRL9ykwApnrBYgt2XkG3nrPinPg
em5xeqXeFULp4709fYaUePca0tQ2nAOtZqyVdVFZewwFwsTojOjPbgAA8ZUi
O/CY/kqHlW+nOOmqntuf31SUqGIVC5MWfcpS5Cuv13RUqD3f2jqYbuLPgOBf
+GdtYQUqO12WcPGKKI8qR5ljBlxN4dL4DGKVWRKGuiuHylC3NkZPKtoG/Wg8
9c/ZFN5ypxpy02pHD7a/Qe8tIvFEufyNcQPXjHC7TchicJmnYGJT8m4WRsPO
qaPgaaaI8o+voy8PKeP0mHz87QiwcVyhZlp8aioZRQHjwpkIJyyKjsVRCTLy
HfhCbQqm0BjLtWTzkEiPMKfyqPn/Bz1MlbkwrQqBXHUCSb/0hxoYckGpJdIY
z7Nw7Mzcc4ryWEYoFjPzW1EPh4k4spznLaDe8nIbaJq2nkWwhBLR0pJx/tS5
sk+Bxxj5VV8aURrug+tvImLJLOMpLcGdznlItgoX1ZXZEzT1xxBDGDnLgE7T
gg7DKhB8I1gRKrmwae0yg+Kr0OzkApeI+UOwGMl3GgoSSmoY5SbbBtiJcMH0
lrm/uCUf5wnv1KZqPmk+vyfjvfiCJ11RsR+KGL8wyrqp6tSOwBuvekTwwHI7
pB8vPavoygbzroTCcHIPSv4XRNIpuPpUD9VkJuZ+d6zUHv71uid+qq4OAMF4
gZpEF05CKMmf+nZ5RSe/91681eqi3vkbRsWZVsbygP+q7JwQuH8UIxHvCXbN
sz4hzz8xFtJwXM/kB3EN9QoYnA3isKC1tpZycc2UXhFnr2ECBmOkUK8bvzE0
WGUJSwvz+owE4ICU9c+DqgxjPH50AavAmV7NMDU3QipmQ4pxEv9WPCH6mPo2
7lIT48wPZyiuZ2XrFXN3jHKFS1y1bdflMmY31tftADXyGkkS/TC7dhaui0iU
87fTJdR+XADIohWYiun1xg68le75LBLEs5EmI8euXsKBra/DcWK+L28+84zA
PsmECXHHFl5gn7Yh2WBEvBm1TnjnQCrEDH+osDQyN4whEvHTkWK0vD4tigQU
KErM7jPytVLDsRhJcE5/tA6tOYTKDqYOUZGfV19qkBqCmVvGPtme0M5CIADS
Ag28kX5coHmRGH6ikVGcxwKLDm+Xsj5m3EXWMqFrNpfant6Id5xrGUMXm1Ar
3RmKOfRdLzVinzAl1r3zP3WK11X7hsLxjbfsT6/9WeR+Q/fuXyTQYCZGHKlF
EZZxDUPacGHC/6+FIwQSY4b57bchM+JaNo0K5+ofWff3hSninLRwQ6lCkidF
VYd1UdXYBhtgLiXNfxYXlP0zMxKAT2MS0iu57evKnnr5Qb69HJF6SbvCRcqA
Q4IHbRoJz0zg9hqIUytvDVJP6ReS1zpbJNzvMB+UCYyYk+KcMkhFOeMwY0hH
y4BIjr3XVd4yrh5A09h+ZSTvOkqZ14y4aaAvs3Z8tjZ5L0qx4a3osdbIeuqf
NlK2Q0pvh191uAco7a8acCKbxjMmRoGBFmqZIh6wHLLAwXkRywUFwfDeFDYn
wMgD08OVaPx6Z4DWR21gmH5WWOLa7rRxTPcPOvDJC0zt++2IU1av4TDgQliH
n27gGNoQDRg2aL/BiE0s9G9fiNvfS0dB8rSClZBI3BDVd+Cy3Ut9ja8skHz8
y+ji04DEAgYTya4MysA7E7gvqQlDONwSl+jOrNwNGMD48tqqDvmrHT2HuBo0
CIGf5L6LwbMskv7Xs/oRnp6sQepqr25X3xj/nvc3sMtEst5tp6IYQJ+4d96P
9vu9+JG51oWp8s7Rl/6UugOrANmlSpj3r1T+wGRelwVfbUZQkRUg+MB+i97j
BFsBJPZUuEL1ryvq8GVgINegQatgGyqJIT9bw3afHmwcfvZ9JAIoLzo3l65p
weC0WDw50rPyb8v+bgtuKOHahLQc7H07yVs6dGsR4HSFff9KVzj2hz5XeubN
BxalM/URaRBtwUmsoMtr78sBcMTcz3jwsYnGtT+9n0p8M5CR9e+IEV0L7wcB
KPVq/RP/Mc6iMP/Jl3AFNqPP0EmH5E7EbZwanzniWez17H+55bKJoQUci/78
ryvZy9aDvQ0ySvGAMHI3RaO2v2L7shlQEXnIZNC1Tj2gmIXOijUUrZ6mRJ24
siu/cfmO6GrYWCbR87TVDHHuQmwnNgwAXC1qiktuKaR1gj6BtFGBR6X5y/Y/
EIFUH6T1tJ1MnTv1PxW1l1U0y1n9swk3iDmT/aga4zRBlD4cKbuXbU0AbDpE
IYsYrVRIprWs5qDXph2Yb4f0VMlokJaUEqC23KZSjEkeBKg7rMiX0Tild8yA
aXDlz5zEYWG5cTo+LleTBHZQE8VWPDjM3U57oJC3FZIE5SOXUUP+MsNeNI8B
z+DVv1t6705Mgh2NatO35cmWICgxkLlW62fwf5baCjclj196QNPpiISBethP
03wqotiVggnKAnaSfnrR1L0DH3uneOP6qK7ZxodFhxDczhWcWBewUvqSlpra
5kSm0lptSkkY1fK+AB2OXbBA1WrRjuMUCqyInxeXBJwR+nH3T1kmx5nzlpTo
873HhMLArcR1HRVMDELdv+nM6OHtiHib1LKADfFd0DnTuc6wbSNoNfHcMYUD
B1Q+OuMrY2C1GxF49zHKXZzEA6/HqhpVzlg6DH2tP7pqEjSe3Sn8vTpSvUCo
uC6fxxGQvNyvlEb9gxvyXbFGMY1X//osY/zbJJZH32LzV3L4sSDXiIa1Bjag
HdjD78t80lrvOBUXGjeQs1fJdeO6obOoOcgO3A/WrLUsqeYAIJMLFamaBRVH
5iPAV5GdbbclKNKQmHkN2jdo0LkM0JtPmIDJ2kPeyq63Oe+a6jKzIKeffBkP
fMKpJx3cW0iTEunghLaveuurHBIHTeGz8PDO6RIsC0rpklGWiUZHXQFda0pt
4fJkRkmPWoKUtvmvfk+AL5jIbAEG7r7ZsyzCYDu4i1IJMk5wefPayIzKSjAR
Q7IEtadQkyk3rePyScclfyGJtVSh4ZNeDJ5Qkk463Ga+PfnMwWyFGEAEIM+u
uUrHzVvEHwgcPs6jSy+eBQsMT0c3B5SXcaz+cDt1DmZntOlNjCDuPY0BZ48w
ezz1bAQLlA5xAyJKii70EI8B0Tx7m/UypKg/kcs2DndAz5mEWay2V78BJH1+
lFcc/TIz6vdJXgzSpSh2HCA/uFtNadNYCKV3wVgOyGPw68C7bUwlkw/HfI4j
TDlbeQXzo3qVJTcHziWov/Gx60VHoLoD+EAZ0qfFr3smhYju1aFYoWVBC/MY
3xE2pcMz1N3IBEAWScLLIq7HoxgoJLDJaM/G8PAMYBdqys7sg5IaFdwYQGIy
2CWKBYCPJKMKnDdHMe430l8v6LgmS3qGsfMJz162FhC1TF1Erv0AF9UMMypJ
sqK6l993p01wdt2uGp2pUWQRdfEWNdkuigQ7dbWerZ9hihuDnhRY2Ms3ajmA
DDmKZW0spPfq67FHhUk4alo1wBrVluamDsJBeM8cMpIRpqsMzeDQsZtFrDFh
ULaiRTeU+zLAVmfE+n5H9tCJUvShTdu9w1UO/v1BHMR8GaGYJOEkhxvMR/nE
a75ygF8i3v2MkJmILPXuywxQEsT89H6gN/Nb8/LyaVHDcuSL3C9l7NgTVCnC
ZPIxhrW5E63Zb3xyRmQM4yY9j05JQVb8BFTBwHl7EiuWdqIX7Y9Z/URXN1lG
UGUJdFGzPwA5i8prqDEQ83HRt29kePzkrc3LsTogkrC8D7k0asWDfXwxYwXN
6HbPdi8O3Di4YVC1kaLFa5jxljaDmMFC+vPyZhrseAdEFQQ3rvi8zNpb0/zo
ERrP8T+qYgysEjWc9WMa/kglcCVDkmjNYk4FagxelKR+3gBOQMhHT9+q7dUE
UccNoK5L1ILHHSiWmRj8mLHc3/hA9/A4Qw2v4uyJ35sdmQefuJWojyu7kfAC
20D2rlGSofahG0qKJXuXB9hcxX+F3ftnr81hnb5FlS2f8VvIdQZvPUTA+ejs
hEsKS948yue1SRCbt0CcFePFPeIt29tgsUhisURIDU8ES3qtfnxzRnJHW7bA
ijq9IbYnkFP9/EDcURDgqB5W2+GycvP+ncLNMBluTu67Q4cdXG+EjSdOAxmL
sLr8ql9K/T5pSKjYp/WulVXOBKm5GOh17eXQDl0/Jm9vz0CnNXG1ZQ2Y6Mwz
8BwxqCbp0dWKpe6GI4xD7FHsokOKXSdKgXo065dpdg+71PuQEXV+vS7mYk5H
fcpU69QsejFPw/qhJJji58z5q5wnxCbC90WFHELzLpgRqve+bPMYt1L+swBf
LMYtgbUjgbSb/qyTlTBRopGQdj8Rw7dCqDZ+npy2AKq+6rPDWwwUcb0kBH6w
DNVVYp2l0aeTJee3FgZe2bh9loi8PtAwGeNsnfn9tTwWui2qm8Lh69AaeX2X
WhB4O1Z/8KgpoNwlu0PKmbA/1/OyC1Y1T7Azaou0P3jBGJ1iXR/+g61MxnLp
5mmZvrxel26Y3IjVjauFQ0ignNKVoJ7HGHCWortfwgS73lGnqqWrZZ1RGzeM
ePFMZyc8YNWxLX5UjmAfeEH0LMNf3ZL1Lblzc1AyQ0Tle5S58X9V7GaOHY39
YSsUeB7tfTYZQjkN7HthI0VCEr6oG7L4H1S8ca2s8f5LU4KuYKqCGYH206fg
fKLNfS/XlF43a1VuXUx5Lagw7IMPSJ4mu/qpBdkabNdCrjn1GDF9geRQsNfw
Bjq3Iwse77loLS/Fg9oJnYeJ8IJMrwl0p3R6JHUsAl5qRPelSn+eh6zhBsl+
K0xdn++kHSGRIX2w0QbUMQC6nXFItsbcE9CK2EDVbcvgDiKh8rQyUd8T2gFK
DXNncpNUbxM98EHBW1wU+5fASc5WaKHIwHJGbJoyuoG8RgVD+3shC45ojQ39
aYGjNRVP6mRY7vZEdDZdxovmPh4mw3V61Dw1i65d+eyns4DaYdU4C30au7WU
X6E0ZhmJfD3CMdMDVD6AMUbnPc4kJ4eoq+ylz5AspzotlEvjXZbpB2IPBHe4
9qk2QK2R2N015FswCiR1X6AGaTyx6RsZPnbZ1EyuXQ930HibirYS3k8G8CeG
IBQRNfVGrJw6OSPWYCjT3GUTnnke8iHm+3WvDPqGKdoHvl2W2TNqD+uBn+pn
F+fzrj2OgTRarawIKsOjF4K39ZghD2MV4J8avGBbvTWEGeyETNYaAJINXSt4
H4l6QnsD5q/zb0wLFLUkS1kveA7hYcPMopePuiC3cR6bMaMAGHYxWkIyvwEV
JYk5w/QPUh9Pwh1bkIDYgm+zVZSzeIdCeRlikP8494J/s9adYWU+Co0WyFjR
pJmzzFHyANKyif/QMDm2yUk08aZnt7KlpeBMLY+n9rrAndsgxZRpmGY8fKnO
DZfo9lNddZ2vB6zowE1pNjFxZga1nKe0ETITg9rrkghd15vLeVHYcMQcLP8C
nwTvWNQM/9SL9PoGXlagZnzUhmLB06ytF90z+tAgwnZ650J97OorSzEGM3qq
uEvb0TpQyLKPtvv2NvxZmLSvwYu/z5r3+FTLNhez1OZSlA1iN0pDQK3x6MOK
/T61ruORlvd0iqCOu9ETAAZYTqAbnxJmQWOOtUQ/nr96mO8m/NlekKyKroKB
D9iJCNQywlM7isJUeWRSZeTkxo6jLZqn3zAX5drWARhVE9MBS7OZNU32TdpE
pEW25XY5fC+8ZMxnrRFGtYiGXe4VqmMBEOv2td77U82+LsXxhHiqpwuZMsfN
17cSG4n4VRg8BkRsIXxzmQ+uHDB7vwZltRVBnKeFbnHjIFdSOAVD2REVNt6u
LUdzdqYOrHOjugpjdB9KuBbs8dKlWrRM9/b1iu/k7Eo98Nb+fPgovHWMvujv
kbJgLqSNc6e94c/GFOa0InwMR4t/C68uwkaXbl4EV3c6SPPhnK5dcrhmzDAC
AXhpHnhtcAfpGSS2SfMp2FM0sC6Bm98MWOLS6ajstkeGkjppJSkBdanTXuip
ffXolGyFUEU+ChxUuPiNuqvlFSF7RyhH0kXoScC2hKQRpZTDtRSzQaHgCQaw
QbtqzehXRkVdqN3eAgXQrVeeNFSYSfk95ghqFTTqO6oyQJmsHyauqwruAfpR
eZ7058sOy/9YYusi9T134YeA8qBhi4Tynrxk6CUB3SWFbTR76neyPd6BH9hr
10NyBO1G21cIp0qmrz3gHx4XpFabcd9hcSE0BccAzQsmtLIMrz2PpANkS3iO
8tu/ACaSMTbRWeAb28iia0SGoCWL9q/0dYymjmYWMj2qzzN1rXZxAKeDDFzG
aiI9NQAeIlgW776EuoFelSnpvb0jttt/y2t9buvbBttwjc6ViqMhm4I+4WXN
xY9F28d3InJIjb6ouFI/Y1KRwaC7rNKgKVE/ExzonLHBrBJAHb3HF3aya+4I
l8V+lILbH3f0GHmMStqwizwdt+xe/2hkGEjV0v6lEYn0FKk+FBTgjE79G6XT
f54vLQA/eYdIa1HY5qDbYezSb41tsK2xzu5/YpPBppE0HqkclahXaLG4ETe5
tTNe9dd/GCD+6YRf92pm6/N9ezyh2T+vFNc+0a0q5VANqxKGfCwdDTs1yiAG
OKrlkAxsoN50kM6l/z6JQGJTCYAhP7G9uSH5caM35R25wtdMGNgod4PpN32h
1G4n8XP45GXla9h+8plFLeDzhsl0WQiO8IychuSo3j0USDZoB4bDcXL0tjbv
bm6s4kDi9aFiFo83cXCefX2W0lHfxzA8rYbZwLudXUdyv+BBVC3D7pL7Mom+
wZ8Ts3DibwCkI/Jb7kd7uaJ1fwsA48crSOc/4NKYGLEPdtNCsf00ujqDDv4h
rxFg+7WWJWjH6FYpBxEQDTEvaFVIJ3sq6oVhDWmFUwLU96MZzUynT6U6B6hB
S/IHRnvYt09QwtbiwuAKzWw8kcKwgD+Nft7ot+s4vRBXwq0e1zSw1UmMl4gA
ZHdB+QAE6fUBEP9AreJhUytI9D6q5KLopJUlixOY1lMFIooL77JWnDXL7e+S
00cUocWtkxT/lKE7DCTxaZgnAmQBTLQOhyb9DtnH3Y7QJ31kAjlZmzy/Edlk
u6EXx6cgpq61j31VKVbBbZb9G3X28VcXTmG9ldN9GBByjkdD2lX8YHdyzYmM
StRamvM3yq4UD0OnOyL7Ifd9cC2qg8Hznq/yQoEQiqE4gl66wC4MQVRJikau
ZctjXeiUKg7xXLNI/Z3YF4G2ZxNdypsfzB7PwMlMjo93w4oNshn3flLoHeF8
SFRlVnc8KsPYAJOM/s80QzJfDyCAdey+lUKfsUVdW08IO2o+wEPc2BWjN3hV
tH4I/3owseaSW5IKyvzPu/kVgHH8Fl3uO6MbXfjb7cHksw1PgZ20SCJpKuDJ
otl4R6CayzLv7lBApHunbG3kyK17GrvID7Fx0dw0hGMJYcqABwCCdWRO/ZWt
JFEjoNRcV2jRGWvOHx/NLQDI1iNzGP3BlUdGLBnCJk6gvCr0/XXJP2yYZsTw
q7JW/kdmFcDhT83t8bD/5C3z9zsTmra31OvETrhU8yjMTZP9PpL7mvUl2+wW
Gfo3exZeDMNWKZyY/DmbjJ31IktfDju5GZbr7/dxv46Kgjj/dgn4Xpzhp5mf
ooQfFmPZi2xq9c7IZ/J6NVoxVsvK0VxpRZm1q7vhSYdQWeQGpnQuwiFMdo+e
P0ZvtwUfbyxQ2KQVjf9YLTeklV332pNAYfrQcnqXzww/h3KlOuJ/5OtTh3md
B3GbsR77AC7bTRjjoLkldaS/Wlfyp6KihK2fb4mRk3T2O3UgN5a4WPsylV67
nXUYAbBJmmoz2+bt5KuDUYZRdcjv9N6YeWJEJg/nq/0FVWNiAws5Tdm+1cwE
IAw6jzCsX6N5MqQp4vHgPTKWtT/0xhHFrRNCsDaQz9SctnxvO0Nq5VHoSjrw
rcNVBQp4yuMVWLp1WjEnMUV+BGHLye0IEUORlmc6IbrrCfiLYZElduMF6Phj
PGg/Ssl7UjPqp+a+0Wawe4p9FW++qa5mdB+VnvjMaj2nGOP5KUj1D8YOCoW7
0/bgAU+MdY8EtN39rm11t5d9BtPdmWMU0joeKWzuFm8uRjUNe7FFUFwVcY+m
wPN71OoBBgJHesaVrmRk3TMPjCcPnYOo4q4GMslOReMdn/bXjGW4i/8oA4Ph
yMpRSXofJGQI3SF4/sAJFolQAyGgNOiiJxqikEIfD7/2s4Di/sEELxtFXUlV
58QlM1boH14m4aTPfQZbSeYi+1ZBCYHjzT7OeOz1YyWbQW3GxQ47OxQLyvtB
9b0oIicdDdrscaYT28d1ZAd2/3FMQLklB/F8bdAWIo715MeVxcl8NraL8nGb
lHVZjkXICpfP4HGH9NsrQHREUbF8K/1I0XcVpkn1HZrQ68iHmuFWlD6/+LGd
jp5dQf0kQ6Wf0PLdP1kET3TYCJZz/7cj6blYXO0vf14gMX9KlO2hkiIC0NbG
Myg70/wWwN+E2Ylr++zRY6Uu7YMIEaISauiaoDgEqXqBgeiPVwNWCIUm8gbv
xrO9f0RQi+sEkptFTBy+9Of7CMwIagzbqp+OY0rgSO7kdDCwfffYUYBJ3Cfa
1mqLP4ft1hpOUxENEePmbSeZ/hIxsObncqwn7fu2zDObzztM+n3KDMx4ZiQ+
cvRYl+T0xTLCHpYbnNGBgZrKKslnJlCqY8JC3kwZunLctTcU9B9Ip4mujATm
10eHg1v6dUL4OKvOcV8rOy04vZujtPw7vZMaTq1JMUJPCQVA0Fp3tM3v5HlU
7IwWvd+l/nTfIJuwvIMXROtCRAe0Q5D/dANIU6RDXZvBgtUIPxDZmdyWTf6H
aCdvupPLkAWP6SXbCjSu8bGf0XrTh6TFpvNB/xd0lWiuTi7F0XKXOv1obU47
0C5QR+Qazp24wOe7dN/ZEgbepbaqZj9kExxUKUhhD05Sq6hG1YGtzwbm7WKl
u35BrmTFwgYB0IOxVlSYGjNlUe7QMYB858Q+hp6lGj/vfkSg/XVyiP4hxQRd
FaDMMBaWsDdq/4VgFU7GClBA5zV2rCXygyiJNI/4SHWH26U538X8+A03MtYE
QfQIT29lsjqVpz8Fz7iQhxMolsRm4IdTcxzW/qRYAQKxA+PpGUKtchb1AdNu
DpCClJYmWfFMJz+XLBzfbICSTu83da2ydiLCMN225kI1vayyg3IHK6OAMNVv
XPCmF1gN5Fe8e06gUA37lLM5HjSRMnJ0E9CosNLQjwXaUYJtlHb4oDvf5N8V
37lhJA4kKRQn05rE1J3QcPF7RjB76Mlr59UnGbBDRKNKf6LynGgoHno1Rk99
TKqhPLOSImK5dgO424RH9a0odReXfEkK0J3ajt6sd+FSgRsxF4PKhmAk885l
hnkUv3Oxu/Itoa+NEpiFM4W6lxPvP6o+urIjLMaoTHbvHLu8M/dPmMaUHYt0
z7IWfoKJ8Y/O2uSIlXHvWyrXZUcMjcHBIY/28Aa8QAJEEPglWwHi9vs9jW+N
Ytki5AsCFgKqVXe6z8J7jaiAs30fX7Vueg5wfhY6IL6Duh5b+48IVqEo1+mV
g2jyZ0ZZptS8eA/zGMWaa2/nv4CKyWGqhjE3vPl7qg8o/UsuSQMADRx24zt/
7JzIUqtbZEQ52dd5lGPvZHotncFQJQfbl7sPrGRvZ8DI4sa0CIA0/dnX2AB5
FIcvXPsmEWAvgo61/Hyu0fOumpw9t5EDi9x/CoACfmdaUfGH+1PaoA4PJgXx
h6vMvq+p+gp5nKNSTiixNzMAUCtC31Sa/joOfiZGwEW7Xg1AfyS76Qmj41Zs
SMVFfokB2wSCpIgKHJb8/PObKCQXTjsyOu83PWGi3a3oY3I9vf8EPED8PvQI
otI07m7LjNL+absNiHFINX01NvAMPfitAjq1tQPt8M2evVToaOr3hP6M1c5t
2NxuK4Np3MvJMnTrXR/lEHVFW2jRylNIzngTspmE54yXUIgGa2YU8qKBFvt4
NQXe9F3i/fIBNLZpKmT8i3cAVLb6R0YR3rKTZF1lcwEdEdL8cIWw2bL2cui+
+SMitDlJRSlZHjsQ2hDPBW8F9fT9BnnPP2Hvfl9IdMMrOqDPrYu+rGzk7p8h
xPTsAIY2oL04/9Yf77DYDkRBkRzZ/A2ZkKtqnm63NJQI7bxlMCdbQzVx8mgS
eMbcuwnmf4JxwxA0J361M6jsM8pk3qXyFfpScIGQPtZFFyvdv8KsGwUGL+3h
R8yWF/EeuYyDz7NHOHnkb6Pax/k5BN+RnnfaOQI2UKWxznveqHkX+BFiu0BE
WC8JPTrCR7GP/YawKviuOtc9Or9vta99K7bWuUN4Rx/1O+5/2u0eig5xqXWG
fCAfyVnm2okwqugimbiiez633+wBmrIfR99aQ9G1VJbla7sA75gpkyVrJOCF
Qs1RJOoU1pSXzKEHFNddqQZb/19AAdHuetz/VeDpFBtKQnvo9INU5zn9tJ98
wl4u5iDIO9NxKRCjiFmnt7t+BIgm+rJIJdaafjPXSufSDGo+QFr7gAx3lEfe
B626wTfq/w0J79TaBogSXDgMLMDNGAqLM52LVfYZicsJqj11nfvy1tLZtnRg
1L4M1sHP+J0lT5SUwa+265ZG38FQ7Xf/L9VlrEwqx0ZlknW48zTUlMTUPvXt
z/7AFBDvVXLBp31N+d2jxsjKTJ5vpR0l0O3aXfIIQaIkTOl9VU0oIm1erQ4V
d1wqo+dq93zg6bFKQq6++5kULQwS9txh4unBULLS7gRaxmHvtE/l9Sgn1m0A
P5OpiegyDZj904noUh1MNrLjV+4IjqJvBpBmxHU9ykBtAu99/0NH4/W7fjFU
dqo+RfHl6FHquKfnHIEVE5Seom0+0aHB89ndcQXTfBfn4G8fYWE/GaUZRdM7
ykLesCowkL612qlOZ3lm6be4Qag4RdIZXVdVkwmUDpRqkGcy8oGkacWyk5SE
naPUn5wG7crGPVfhQjihKhNBPThFLJcC8akpfzk6p45+Gq/a7zXrUOKb0D2K
LY4pwQtxZVLhjfW9XdKmViYcoqfs8IMSjeNJAVmxUeQvFE2ooqCwq8cRb0Qv
xDIZtjLt5KBZQ8+Wrm1kvZwyyER0Z9+wZZZkJ9lUj/Wht1vLHwKDrxqawjFY
tMmJXq7CnQbQuAqllzJ8mZkqFPaTQFXto2aVKamm8387KNJmLeP5EBzLkmAk
AIez2lkGGMQ36Vmv5IpURyg+k+JEJpk4JgQfyqmnvt2yXe2Y1OzmxK04N+/2
myiiRIkwJoaUKS+2Equ9PPVBgkX9yDphvs2jLQplIlgWeVbmhPNu1J/l6atp
I7RIiW6StqMzl671TJRmOyndopk5cnH2bUMSvhZ5y4BL7IdCi2cIhfYskoRR
+FffLGl8+3EhnXEAlHtKyDkSDsv4JFijNEE75Gy1f2BrR/S7x/uz3g4gIV1m
Qtek0uYMYgzJELM4XQhEMAx2ijXkqa0LzLrhA2SG29MGaWwcTc3l1RGXyWbs
iDKj27D3vazCSSr5AWXKE2uNppu2uTnwxxWmpKGftNA66IKH0976ZZRh/qky
KPhIucvusCS5S6DIviGiMsxUZu6CnteX4zg6ivq2HzJtx/rzEj2uw1dmS7qG
gdiZO2Aiifz9AGRC4jOkm7ar2B7XUVD/XsTOl2xRaP8834GDN1JumlurTP0f
wGVcHUk840aQS0qtNRHUjw0vtox8BOUKPRW5/mZDHwrT0TVGVMc73zAa68wJ
Sg4Wf60TV4ce9oQoD1WtAkCgdwAM4kU3386pT+9ULRqZF8SY8GumdmezSMeV
zexo5tJKpn2yevmosNYU7yLSxTJ/Jo85oZ4OCq3ua3Um0iabsSan6cOsdARr
fhNKjHFclTMFSVfAwqBNJmUn0i3hZSH694wEO+GQR8qSJuhQjiZCqBvUT5Ta
pNJ/zW6uXkSc9dk0Ir8zvF/A8czKMwe+uA5G1d9l4ndEiqNU7sR8R6J6Ugrc
xhtpEz3qDRLQf+A7Y48R37y4E27gd5q+xNKOzWCcRwoy4nLI/hihwTASkj9Z
R6zKRMiTG8E7R0eF3JonuR8lhxGzimaVrS9fYbMeBNxlbNRSZH+aYn4ISjVE
PUSrmhbftzfLNOO+4U3nj8/ZMSo1BVRYjn2HLyz3zI418ceUSER+VBSAT3fK
5XL3c53VlXXk9zAyJqxuQpIuTxYl0C5kIY2yl/N6ZDwjDDV3KrBZ+5Fl4M4I
LPOCKAyys83XWMhJLSERlXTcVpkTvp7KgQKtHcF0Y4ANIhg3H4dvreR1Jsyz
hYUTmQWsNaRpIIr2lBmP4FSpnsRckCdGgQK88wJ8as4IKAHNAfvhLasCmB9U
JlaFzxMKVqG3ZSxnEj3oLB+hEZTtGPlikjfRDfCLpDA7B+mNy3S7j2neBuqm
9HN53K88eSspE5Kuq/xlhud+a0lgIhrQc/MGdiJlhY0ibrcGnAoWAaYHtiod
K/3yiJxZLcVL+j7c5pz34AImIQrmJbbHyUAQCH+H8XZQarzKLVsrObYSJ/tK
zi6BX3LynCVxJRBbFgtUqxAgwlSetkpNXzBtp0Hvt9R2MtNp7S/eJ8fjHJpw
U829ouxqzFTNlhNKsMi2mKdnxVhQ+fRNjhvhaYRz5eBFLdl2M+DNkm8dnrXh
GGY/A3lQhuDN4lp2IhNh1ZSO6D3qIj3PMY7PWtnKA8tU22kbMzLSd7VwpJin
ARaMLZSjWJY3FNByG4h+srrLBSqnsc76nuCgdxIN7d25jdXXuRcjGU3A4kj1
MxUCp3N7Fv4LrDXZCKRl/oldyMmDt7mbFZMchSg34yCrkEIS0jvwCk06pTt9
NWCCRytLrBDGIEf6/Y7ixhsM2HtojnkeT8yHV5/Owp/6vl+HwrbjN2fbZrep
OEF4s+IKv9C+hhF7xkcp/2S5oCjFNO1HEuGwA9K9Ib3OeOUv5/z2hCR/rcNT
9gVlO5rL6tGZTYh84s7lYfXbF/ghK5YvXQEa1+9/xNbCWJVpuBf7jirg1Qw5
eiCsdilMFa5qnCLRQj1n5mDezBRCXh1JJMmD2j1ec0tg1uZR4ES19Mo/XedG
ObPM62fl+YcNB0uzMgbcJfTs1Nbjm1YyTaZorQ3Du0eS5Lw1ZjP6O10tZYce
RKIyEcNYRgnhsr5zeHTmIAxw/jxJXVSAbvee84JrGC0EQIg6epbuGHP+pBpP
u40bphJgCv/7fyHP4BfQxqwlB2Uvb2EEmMymu7XmbB+/p12mS0znQ+9Zx+eO
ybDaIISfuCyyu04WKoYzar9ukwjttbM1vw8nmAaxbC6sgJiopf4nUVcWCRqP
+QwgcG1XagsInAboCOjGchO2EW5SIzAFHtXJ4/ge0Gj09JVQI0/aZQtdMjZk
coI0UPgpw4QXpbYSHi7gZW8TZ+NRFgrhz6lVAM2kt9h9UMZO88LVaXhtTqI0
dZ5mWFReD8EFhpcRcsfrJB68TO90CNH8Qfg9/IStpPt23v5wiUKHsObu+AlQ
3xxmd2w1VeJpmJP6+d05nm8t1kR6ahiPHz+v52lHREnG4DquGqBgY3B/nMvs
cxnXiceFpQ5sU2FoD4RriSPG01z+Wq2LJ6uyTXvUdC6wTzJa8lnt2gy9n/yJ
/P8Mysgd5qlVqOJIwituxKMDs4DzpeQqVCRh7IM9fR0nFfXPEgHNyATA52H5
yX5j4TlvXtMSedKpCDLXbzwh0lhWJFqh73Gc7bf87lRdg1C9D/avmY5nBkBp
hPhIwMqbgSUF32IwD4gBflzsz8THUWFlfEOjmEHukCKrpNUNazyu4MRGtrk2
vJ5e3mRHNOCVqtXd5JVISzd/IWPNUHTzvw+galNz3l5KBNEJUbzQy1HqEgPG
z8fEHS0P1SSX+CFWXXfhdhzF50a5KOYOAZCp01oqW0CO22r4+VimUTHWL/mH
TP4rDVbSdgWUPhlUKg36NaDNtXF4/M3APDKXSuva75Mly5yIGAILfssgmNEi
5HnTeHUOL7ehCef98mXQqv0v55g1T9Ktue7tyt1HJpLOXQp7f1eQfbQc8bMf
LKeIn7DFj5PEGWR1ClOdfcAFXyXYEyQsJHHDVSwrWkwE3Ht//zYYI213athr
6UztcgLXHSoHopNGJ4Dbc7+4gXSRvR+W2QKqkGhsjmQj4sNs550efdqsYqw+
6ByG+HlnuP4Ab5EMu960ZGbbDcUq738ZUE9d/zU+mYUagTcOJbsC0F6481+B
QMnsf7cn3WQREjx0KYncvCZfuJ109yzSjR1K6nC/cv+bjBkfq5Nm4lP6Afet
xvWyRZV5paBCF2Ni5xlVk0Deo1yiApB/bg93tDc360yVQ64Ah3aQymNEHdR4
T4edhGp988TfbwXLZWqoQaxDga2iP79aNHYipLSvep0GjdaQDwFm4kWtDcW+
8blzb5OOWoFds7SZQBFqOYpq7wEp4R0L1kd7bSwzq+2G4DipnGzKLjdner2h
Gt8MRAwXUFofv+O3d2cfoOuA+n7UG8eKnh/DQ7TCSwnrWb2SH5+OSbhI3Ydz
Isj8br46z5/F9QblMO/iiz9vQSHFEYo4P1LHSrr/mLWXth/huYPKNm4r67GY
Zw1draT6jKbDeG2EE0GGFlDHYSIQHExtFbSiy1ZHOv3woX3Ki8CYXN7yKmtA
/D3wYLkjatrxX6b6zXt8q1+Jl46b9WKWUMKZ0YLp2sFd/D+8ZCrZv0Z6Msgf
lrQhR1X99uV6DfwijjMETbQGk0oJbk6IpHGI8KCL7ChNAjPpdgJCqtl/RnJQ
4i1XndcvTqSrtsAEu20+20wxoy8DFNP8weP6kZYKBZAdrSHIYR906cVXIQgB
xTIPiYVyf7RMIuMpNL2M2So1KmUOd+2HQzc6sGkIqHZZ8WlAALE9iGO9jELL
mb2wx9ETQhLKygG0FV5j39SP+pohOVSjJ+8YVu4vxxJSZVXAWpmGJY+zzIME
N1v0r0Q1M1SDfp3ArLihSM/eS+3V+US7HJXX26AZnpfd0roNknCVIgH9IzWW
TIsb6Unx36877uL6gnFalTsILed0xE3MHqXh/mur1PcWkkOpD/SzGhXnkMmx
rFzl8d1OaS3h15xqEWoy3x8v95umBF2T1qeJh8SBG97lQ0iJCjZCqAs5DXVd
xLd7sGD9XZ7smRmvr3i7HVnqTc1V+skxGsTZZSvsxWVX5JGcGJykWmjtP39R
+MPhewcK+knu0lf1Dp/y0xck7VjzmbZxmyms5XwmgRk+GjmjciHOG7f9z309
b8LOJ3Rb4Gzhzeuk3IGLRNZ66AmTTuMaiSFbvFwXu3iU7xWvRf6SSjq3RUB8
U7NDHNc7UPTTgKPzKQvUhjlTd8ZEHm14zVSG0H0QyMVKfhhYW9aWcrPFBZFk
90Xb4eZCB5e66JETqBsk5vQEg6z9QaIZ0NMqZsJvdhY3pAzC/lv8WJP1SGZE
n1TXegYVTAlAUuhs1RdceN0X4Q/BWitxZvaurpDM9wJUj/1uQrh1hoK+PFtS
MM6kTcAvsReO++CxCXRJhkp5+4CdZgLNA8b0MV4rj/lLVmywX0hCDlfS0R93
757IqDce+NFbAjq1SLDMX1v2I4RgPJKSorbtoS5uGPCVd3W66+pJx9DvdKsz
Ae2MajRui/0GASYaoAbo2eftbIRRr9DampmBSyhUFh3j+HWVtXUyRzKcYgP1
rufMd6z1LhnSRV0wCm/kQMIYq8nQk0HMzh4ewHVokomzUDtZVocLhqOk0arg
E+ibcMOPpFP0IuhL//8RsGecJCKNiGWaR8vyveL7W0iSySS3MgXKDODshDy4
u5jWwYn/Zop3h9aZKgyKbOBDWNACT/T3tF1g1yfyD4V5xl8tIK2/tv2nh5rr
MBYGkjukBH4EYEgyeqw+9QxBui4wnE1uK1KmZQQeVugo6i6FgEOvFDPxVnBU
39SzmCAPHikw6JaibJZNCYe8eZIk/1b18uY5qSvLAC6/wWfUi4Oez+xgR3wA
IUFEK8kmg8FNf3aH1frByrRVsCIJE6kptCMQ8Gff2DYAsr4yG1IHwlcl1nSe
aJL3GW5YF291MKoUaR4QFBaaGtDx+EyXBnTdUB1g5eseo35eQLg0WihckRFD
8ZWIXTr9ISxVm2YnhIEf2DzciqrFvHvNm9RZc5xV+NWITRe2UH+YLL1GDagY
+Jx4DOVLZHXHqe8jMAEt2WB+57vzHEaWuNS2KfvAsRZPW+4Fqx1IeV5W7wDp
ZjUNnEX8jJvGLitQHgBhdiapOGT5PR0yuxv7mXty7K7l4vJp6XgljSPJmJSq
RbijuUGAnmYDLTsGVogbPzvNSKrkONVX0uvQoAh8bEUb5619nd0Ze7Ajrwft
bmVEz2t8WtHBWSkK1AhIaEDgxdM8sBpcBEgHtQ4hRs/ySYS5QY2Y+8aqsD6C
d8jLgZrGf77xVZ7zO3jzNZokJW8uhrq+3pwQ5rp5UeAwgs96wARQxRQK7F+1
kdBkTq2SET85X9rdd7zwxtnBoVNhX1yuRduCZJLQPmYD320mx1611cRdEjey
XXgG8kOLblHD4wd1jOnhcCsrkIB+sqMwhdnlCtBvxhhdIJwDMZiYzp9kb4rv
iSvYNH6uG2MdgCXDMUDxgfm72+NjFcXyfJJVvkK3KJ0YKdLa0nC23AKBk8bz
m3coXrtu0UQOOOSeOx/80B2/tFNa7ZJHftHTxnaZN1eS9ey2gZGm/ccz79iV
CiLYws82CAIQK89OIxthY3iej44wa3AA1yTKJKhaDu6Wsa0pfFJjMC3wSQb6
KLZqPSB/tEsaJuvQugqyoIt0Tgb1/1UqI9odxvIDZMAY6Kk9fyhg+6Yw/KbD
iZTjpPlq7wjgxfj4hz/zbTxQJCUnUJ905jLYsZ/RLl/Ns6AKyr5brMaG8fIg
EarvuVzGkD/5+1xT1o7XMTbX500r/vGUFEGuahQa60MpipEnnjF1tvVz688F
ny6OgcaiDA4h/xdT2M+o8tA0oeXybEFif5ox7VM07fMRnOg1qSX2YdEMuVjf
0e2Xlfo6TftYMvdcaokn8/EeTBAw5yNOA9RDgA8RVBPqrN7tf16JasRVPS1c
ghjS4gtYViYL4KaYPY6l8wM/nCGF4lqENcuEyxRCtPXLfVF66/Jw54Ja3Hbx
eBZKtaqmr0AXMV9E2aG93DXbl716+YCfn3eyJywoDK4n/3xzMFADQ1QYQYi5
NDBv1rvAS/f+/pRHNHRRBBxhRkFDYqmGPU2cr2LXkYyH1sU0vTD0lR/gLtap
pxgsM8j+MLJvbzvXuZfRAgFf8euSfTZXqRhkG498pHoQTStpai8Eg01yztFm
V/wg3g+X4q34UnhoWATsDITC7VFydqoWgD8BxrcQpzAm6+SHreV/4ch2u+1g
suj1LlnX9Wj+L5bupdONpmWMVM9eWoXHBOzVKTZCNU/mvVbwFU8Xo9rVEL89
K6fmdLDHOAmJ3W1lrjGQgHRULvbUk1qEqlRigUG7u1Drhi/hTx84pNX99ZIA
4mYIoT/JO/nZ/E7dZ0wuytjNhBPd4QqroXFv3ucOExbFj/hq3QzBizmhhqwF
ISlMXAeg4NDxxaJ3dzwFevgi50iF3UIWQNnK+Z+TVvwWH/yyVGYjPHaTAzu+
zLFoJ0ObeLlpgrqOcRlKalbXV9OnIe6eI+fu7TGSiFReNI6DI0DdqWY+pgnz
Lfxi6tX615XoKWQfFAEDmCU5vg064i4KJ89tEdbSEAp88MkWHhgX82zU6C3d
rX2JqREY9pj4DLaroiQnukJl2laDZ+J38U69jnpciUxwt0AOLY2HeiN8bhVt
mcec/k3v30viaPa5IYeoaGQI6aN8x3YotLecsUf96qlG2xQmGX7TJeqLxRef
gU3NaUJ2hsux3FUxXf0K3j2z/AipGx/smzGwRnp8QqW/INsMn2JLjMSX0Wrr
V6Lzya1viACVvfl+osIfRuPLpAUueoN0nF0n15lNrfW/P2uY0yVd4PkZXqoG
d2X3U/YrAUtrMEEtMJ1Q6nLgFx/j7DOTdR8JMY8sJVTOlJp8FW/YR13ZBt2Y
R92Eby1XTRdq3MbaslJZkylYAFGt08g3QHCULLY2pCK4G8j4Mw+J6uVpA3NK
mjwtfFz/V/JzI9XP/b8Ats5foFaxP0b/YZIQeUR+cj3Ru1ftYpnouVYKJUnD
V08Mwij2ywks6o8PZtzbFlQV3tzqtR+nvkn9tykl+ds8CbBzMQPJkuSVHO6E
E42lEM+Zx7ehmpa+eKDa9dmCF9bivsdmi/+qVCa7Z6NhwfaCHVNoRUeSIr7i
+kJpFI40bnUDWyABzxJl1cc4xxLoSMtAPVZ+4lpAuTF4DXaKmxG50gXACPww
k/6Ycmo+BUlNWPr3i6vUadTZ42canq+aS0itlkQ1UmOXbhM2FTdgiK78ZsUj
We65JyHzzJXHYXZNq+aaa1QeyLDkNT7FzFtlZGpEcwncF+jfMb2Z0R6xt7da
YqyEYawB/q61oJG4CNoekU+nK0Bfduogx4fbctY1LH99Sg/b4/I6HX3JKGl5
UOkTBVkbmcmNmRfRKXiMIHKNKyWu/qbKN8pJ8+MKlZ8D7M9uu47jW9+DOvbf
l5Kvjv53C6vzxgzGaXexNiBJMuflE7Fn8Ln8Q0bC5XUasxuuIGULCSrPmAkI
AYQ7XHlcUnLLt/r4iK4vWP8l4y4GTPwdWrGlM7GBTXFJr4/3Za1VlJ0xRtgA
IUuDa50wOBMhGX3LPtfcRktnMsIqan5gc499Y6425BCZxSLSwZo/EXgENRZb
q4/5wUhrVNaYeXE1ogv0ISFxsfuI2Wg3Kr2/Zdm53nInegQRKtYkAWRYqvia
NxWJ0mWislUVXylfbTrCLYlK1vlYfwyrKjU7apHH0RIRSvxS+1f2L6qYnPJq
BxdtlXGAPZW8G5XTk1JHlON6pbhmmJs0ac7KcymHcScQG4ENQX7l1ZmwIEzP
Zbdg4aH8WpSlE6chXsTyEWKU5e1DqsJj2IAVjKHE+9uJPuNT/cg/PcMRH1+V
MQ4v6JEA+R5XbmJthLhhoA+9+o6ObewnwQbZ7y7he/RJf01fBYueueXjx0eT
jweADo0+JBz7ZzHv0scBLxU6rjcOyHQ/l2LWvTIZfXQbkA/tlJds3pMyIs9E
Lgm9fyzw61yxrGqm3cNsN8Ja0/cQFHVYDWcbC8aytpcLxOCGeUxkxQAvX/pI
xkOr4wrd4yfEhSLGpZZ2C+58ip7qUgvp1vkdA8APbzXJNZUuPXzWBQaoefFY
OxgsZ9acT7sS+cXf3XD9xjyMPkKNmQ0H+9LLVDuhBOR2Nrbyqv7I5PMzeRAN
g3tI/O3VTBmvUMS0rEOfrotE5BtEN+j3YoYHZR299MLyECnnAnH8Uk8aEPB3
4eq33Hq2WVOsWq7/DtvNtdQlFfYOJuArwIiZaXPq/wbosMiD8DuUEF1n7+nk
oObsaWn4p8JH83DEuH8CCKD5BoJ91LMZ2/aP1guDSXf22TIVwAym1tiCx0t/
XF6qXALvlV4QB+unKLJc9YlsyK2Lqz9ohWAxd4h9wDtf/fDG8iRi0fQWY36E
Enq/4LrjCIERD4ASBOzpWZzk8hZ+8duaNElHhqH7htqXRGThmY49rBZAsSiz
QfkyWck7YnmCR0SlbFuYYdxCHz+gT+BNpnHaTGcXVxEpIvngbOJVIzG3Iv9F
V+Xuh8bAuQDrM9O5Qht7ETjPj3EZ49Wfbtdu/0HXRyT/wGkffMzaTQAJX2Rx
YhsU4+H+T3qk6uZhznEcif1706R0W7rJYM2yJ0vANLzG7/Fe8ruFzjcmlQZm
y2UowccymKrcCkuEmRoQYV7UPBjaSBySKy+HHjdbNEUQedORF67gdgCSnL02
dXAIj6UfBzcJOBTsQKEkI8HPlZ/bGx1O7s0ag9B0CMszG02AaE/cjQ/jdAzx
lSnClNSOtdchUBrADcFmxs+AkTMmmNaGaMx4Vbdl7NgiUoSjjZzPm+dQ0ORe
tz4DA4RtmYNDvL68XmptcKLDstzzBa7JZkQMQeSKHlFWWZhdB11V8JALwUmn
aj5xkREIPBSVhcY3z6iq9Z5lCzcgtSRT1KRwmzYUTnZ7p9Yn9mZ01SPs9xBK
PR7X4A115CBKyTxTelEJnWO6dguvEgaYS9vosYzN7xL5NQoKi2qS44dR63IY
S1onnV/4D3UbZJ2ApvG0Txxje+y3KeoJvj2nlOnAiEr9W8Bc9/SPJNUnz2Q/
6JjEZWtqdvZdSYbA807iG+V80tDgyS2E9S2JWVDHJqaqxhlim7QQA8K+TJFE
e09VnWNqP0/fMdY4chKkoDXYm7wodiGd/spfo5aS6Hsi6eO69NipGyzzS8dU
vGRBP3c9k4H3Svje4IOZOHfPhy29iFy9MHGrAqPy9JsA9tjLWU4Kp/cY/IZI
4Y1C3Op+V9GMZ5pRfdwnuQrcX8x7AaHSh8dRh/iuk9Xw9+IJT8K0PkpkQ6ah
TCXDFwVv46KOWdPGVB5orsAt8tj3vFdK5V2Inz4h+Mbk4bOxSd3niUpdslN4
epjBpq4or9EVrIS4PSv1x2CS/gHUcd89B9lRFK/8NSHiklI0fRU5dfBPp14f
42ND3zkoLXTNld74nmNS6XQg9ANESv1ts3DXqxptWoThGLGr0pidbj/lf1JH
v6gluum8z1iGo086ABfdEcGODcbxFZ04XADylThhnHQtXWekVQjeYNUouuFB
8ut6lKtYIN+JGCKGPyA/Ilr0HQ9+8ZHxEcrNEAQIr8HXpzZ01m1YAKxVDFB6
YTfVKT5QIVvlnnQgWQeCHxuKoFfpNCeFqP9Nw5zPhF0BeVDqKOdJTnUrrlcI
jGZKPO+CA6zKbADRLDJvyAaVBf/HwRLv2GkfR5Y+jQYctUmBs3j/FGMa2eW0
LZGR7cc4YMnqRzGGVqqjYLwTfad2JLZl2l1GL0bBwFjbeQDHIxwO9GZ5cHQz
JSQrKGhHsZlZZMm+eaidPfXZjCRV23wQyT4ak9D9b7VlN2LzPocPKtQb7DXz
Awj74wMaFO3+dTaZ9AMom3pnYsJr14liPCo2C9SqG2dNmNC5F77zRHuKZPHx
mHb6uZkOBzLrAjCPb0Lz7ti43IH6FiAGgYzM6OcAfJppY7cy7GjfbWJtpicg
jfULsusuzQf/EmzEK059+b8hEk85mG1TIiDCSo7/muN3moejRR9kAOAaMpPG
g3ZhRCnT8dP5H+uB9MhJFpGZtyko2IsK1psgWwkNCW1pZd+Li16e/2uiZZaR
zIg6UAUdUe8KR0T3lO54wAPwU4X7tYpuuh/n4z8mvRxZYCnjF78e/1Hwobtc
HNmwjrf8xuuxJtjowRJbirKvf4rXciFsTwSg8H/wlMkzf/vy0SBYlQt5Kpn1
0I9kj7CB4kPcO3PFQdFP3esLzCw4IcuWYxk7rs33LmNuEa/C5J5qozL495vM
FJvLjCJ1458YnnR1cbA8IzzXYdEdFfnL3rUPVJg+JxbfjkCS9B78CpcfPY30
v6pkylMUXStOEE1ZkYwMrJKybkVDlKVhOmYzzrv5DxcXeNDl0qxDFqz4Yd/N
lby22AOukWhKQbPAdxnvD639BQ9KY5tZekjo9lKSuu6/OXNL6QtPief50v0E
pfb5cfw/rrLDswOmy02466WvRsnse07jEDHn4iOulHkB6iD3slu0hj2t/Ckf
I4Ji2s0pdiOrNVglqDSAlK5HLsnt13Fj2sbkS/ZEEr4TdEaykrkU8OgW4s8u
/MY2Fz2b+njampD/id3+JsHNrG5+pPNXkX8mpRrp9bUx+bxN1OEiJ4cBx19H
QyTL6daY/Ux6PsM8dSKEICTr1/hFvnqWPCkx4HAkiSc3p63+jkObpTWMpGLZ
+zrD5cJvomBgn/lUd8v1R2xTiRJfBGcGpr74qZl38DCtsh0QQcB3m7xR5ECg
y61584uQtQvtcq7Lft5jIUGPT4TbyRwXr/4G3eHIoOo9j6Gd/BqU9xibellV
oh+SZFcM2NdrprOZXJcu8VWRGPVASZvmdXfemmuSRSENJ6zmFykA67yhRaq/
1yvFr/diRwW5wsmYdpEZZgynHgBF1XoykVmp6tydVY3gZwmnQxeJUECjw3fM
toeQO/J+xmbaZ+6zHE9q/SOo0hrJYEiQaYlWpHo0NInmo7pSmc2uvylOzDp+
KsYOiSnFTpyonj1yqkSihz5s/lcovMtgVYvVX8Sa3s+jqksEY0cWp5jAc8q1
DDubZXB6oTj0bE553tYkvQLCudj6N59xlFq0Pj73CLTc6RPQPqiUlwW94yyo
mI2s77HpaQQfYQ4XkWVpKjOlbrvK0ObIF0yIytuJsP4Z+dk/KnqmsNs0c1zg
Yrq8bnUmGWynjdHAmnsC7qIoaK/15TSsB2GO4VXlOaVdEg5lihnn4WoYPWxo
DEeyAZ6WfOfr5hv6Lb4SSwgcT38s8ZyD22aWcRoplVh9M2pYbjjMwWAcp2QS
wZ75Vv4lUoL11gY/6yNYZeVIYGGMC0uiNtTbCarC/iqy/q1KZ/t7e6GABgVr
71FWb7xo7o4YCXKl/fBjwJY5A4HFpX6W6oUZhhCga0XEtDPJJGY7HO4JM/Nz
qoHNdUiroJTWqSv3bwMbVqzLlBvZYX6fK9w5TyjZQSXMmmyp6RHqbLrr5kwm
eqqXYclm7304Ls1FcWPI0vF2ZIfH3tiCYhlaDPs1PaTYMo531ESQ4LMYu5nj
gIXB88kQTb+Vl+fP2zICXdRv7vztVkKmWs2lD5YPgXZkujMnMlMqP39IlkbA
I/+yEIyiC3u456b2K579bvzCnUw/LewC1pEbESV6swONt275W0rsXJBAB0Pn
A5rObiCFLzJsNJnrFh0zAbd2xGSLt8scEXYpR/3Ih+NdYVxYQjOrRv34AzBw
rFVrDDVowksfblL2+EClWqqx7CkZqlhpYWKKxXW0VsTX0v4przv81OCa7CsW
dveNSDHIKR+f2Tn6SEc8p3xhyZSZJ4j+CSb5+4x+xIux65B4JBiVn4rMuhUs
CGa+HY1eZ8+YYqSq133itjmkHeNOsFg6zPaEbS5a4AudBTTYTh2iD3U1LXQ2
9y59FM5tdtIW0K6GC+V0UpHNcZ2t8L5t5eVuse6FNrB85ciILCFjxlL+XsuP
W3JSV7XTdnOAxkcCv9EblgVnOlsQ8gf+cFicGDnmO9+/Uh1dYQjr5mVm3jTc
czaeIL0yt5ucX4y+4D1IKdLWuTEPV6h8HoImTx2n15dqV8RSO1L9kMMnHYRZ
ai14yUcHTFRXMQj5fWv1N8j4XVMjPFF3WRr0xUFjqnVI+S7xGq4F+XjOs167
uU45UojDzvRwXB3AWpA6OEityF1vSvQk96qKHuXMZ49ZkbZULqAkuwQYGguM
4MLkwjFbxo7yQvLyYHTiM+4kapeiAhLZEdCT+E/z6r/5iDQYLQC/a8DQVpgu
ZSevap9SiGGcF6e17UJijE18lz2EFPEyulyL7WQx2RvHg4aeUFGpzgdOXa/Y
E7Ti56zNYe1wasoEDt/upW674VaUZBTVlvArLKmKNeGrkMfTLBub/7B1p36+
a9X5GH69TpC7wPBGsezYuFjpl5u9G3ANtn+mkcqhEKjtjIgEjyGaJYRPjUH7
qAZjKU8vXtqS3akihEHXrAHeLjGObGvUN4+ye9CptKIOjOBYqs+Zk9bXW7Dy
xrLKlkQ23tjaYa8tnhnhZn8+oEvp/PQS61BUckD6jBAVuosezh7iziKOvblg
4tfHN1FITf6mOXw+xZ/AmeF2W6v5OQN5g9OIKuLJzEMjSO2sv0Pc/2ibyPfh
7ZQd++SNYX9EBfwNZPWbbA0hvz8CNsiHdvGyeHIiEMFAfTPWaAZEnECzh9wW
emNf2jdqDdpuaSeRipjtF/NNmdOU6mO7Kp3wm5CYuEdCNciMC24bWDVs4fUL
OKl+3idrfUN9Oa4DYNfr/FCZR0/ZlbpyZ0aJboZLgHwQhopwP8uinT5p9eQ8
7GO6qJyAVFo5t6ZOh4gydIIfzGpWS3gsajtG3wRRiUtiMtD2/XhG/SCQMnnp
dmco46xxb0pdP44/PLPAuJyR4+8gi/YweQfEm83aXn+XOVLBMRyyQP7GpfmV
02BroZ0QA+CazMuqmcJPVSUw0jUWJUEYsXnwTpGhcFVS2a9ugvcoTthP9F+/
Zmy/p6bOh0WugzbDcSD5GHpgylBk0Hnck5VDTpxBIWoDDTr2AMyADDptoof0
k/kXGq1m72Gsm+uTdqS3sld+FZI1vidv/V2CnLVPMWLTdWA/fP4R23+pmcri
+XAZKLPXDvajOHL01rgB5YjEcDmruXKxUOu20npYA/Lb5Zuno/yZU/YBe2IG
fud4eTuADXGIuA7Z1YLZzDvMV09YMWtZWa+pFL5MjI3UbOIg9NPSc9HppxL9
BodpVdm7/vzPqI8FmPQlT+e0s3nNV2+3OErgZPvCAsF9vCZVe0PrBGsdD9lE
O6m27TY2vlprRc70pdfr/wqMLaft6NpZhZ+D04OZOpkAgnk/VyIDF8X6Fa2K
RMhqyaYMfHVafjiEm/iZqlv7tjytcMrB76Op2N0Xg+9WWKABtG47vY/4uZDQ
6Agim1CyrztNYqCXRoXqNSHrKmIu4mVCw7bpNVHNLX5439B8awlmMsRM6SfI
pOc697NckAC/5cKM2LhYCTq3jPIRhxOfMk74O6JLEqqMZ5XtafYi43HyaiTV
LeC1ASh2gbYGUM5prUGJguLsmBhOAcxUshGw3TRFQkYF7j5LHokV2esdF31d
bY1fkI4UKVdp5JTcCwMx0zqI2FUJXbje4GASLt/LdLyt7um9LxebstRP2cyB
1hieWtf64JBURATngsbY5qK4MF428jlNABmSHpcRaBvdur5gsW6n3dDkQPGS
BJvv/NYU86f6m2+DhsbmKtYF+ky6w4Y+eynwH4iDLQpYLdbxQvng8MGZ+qcw
uuwl78P9vy0oLkFozYUDvyz1gMVBr3GRrRB2f6U3l3WcrDgvxmtw1FG24/fX
CvVrejYroVNPS/qiU5f+1zfsa7KPpDCuW7/t0Dj9/HUjW/aNpEE57/gVU7dl
Fu1CM//YAW2rG7Ob1j0YrDOKHQJAVih7Vs952H7VMqeM5289gQSVl1XoaBYT
VqPsYaJPlTL8peoB0ql4jA01yjk00tfnHeZxzxFx10xqUghBWvwPsXsq/eLd
VnJwV+a6dqj+I8oRSoiQE3bnKzI22rATrtZfoSeK1VdsCmK7+5ZpZyAr+24m
PTLm6g5xOuQwErBcuXz9k7rBqUsWzd0dv70psqGnAtDLRQRKsc8/3ZFBc6gN
YB1uYqzd3/MYQ711KYfG8AuclLQqjzPDG/XePNblgj1PVwky+jLyHhDmjGAh
QWMKyZhWCmfFzOfYP751VdGjdUwiPA2yqewbLpvcgnHr6ylbOyl0bj0TAC/a
bGsv5pELSN3oI7pqHkMsBs4zKKOfw8HrQej/QyFAlBwC4cHnqtH0b9IStCEO
8NgyyR4Q1nWa9HhIp2c7G60P2xqluWKq5vSjCud8dXK5Ocl2dTBiJdr6bxpu
XButi2pb464MFWDNB0euHEOLEGtKLOF0UMyWsWrCKbNZ3KkcdmI6xlIdyilr
p7lDHkOBENJmkM1lehq1w3hiWCZbfMoN+nthuwIZR9qwIWwouwG9DIeI+AY2
pDMz9Mgh2prR79UrzSMRaPVnaoyj3NTCY8clDlFvxTpkLuGUzxDhYpZ6c/1D
ttjaNqfFOFcKw2EUGdqVjROcrEtELrcBpyTPEZM/TciYcntOlstxtRs93R4m
QRYVjJsl/7qZRosqHTMUvWysc3PS2HNclpCEf23mjo7elwVe71Xxf78kl5km
KGnV5hmns/O2oCqQXgVGp/knW/PSlpZjzGS5f7cWuNNC6+VFi/xBXF3l/QTR
mNB+ZdC46hgkVpJBpXCBYOr+fXohXIXZZmRDe/J8HysDxtA1UzqfWUp1wuLS
PNfvciIEFH+lQwIYNFsGtoQN58LG0HgVK/Io9H8RGqfOnzUGfSHTPT11RPy7
BVCkp9aJiY/dwXKJ4OuPxV/BozuC1ggPOlrDx2cO30XUaHaPJ3FBxztkN5wO
uD6AYCMTp4auUSmNgHCN/Hj0eXDMbcJUlvFrqds7Aq2GLXMnAV3QQqu+7+13
zFOJJZYSPD11TZqZwgE6Y9oggV7S/FaVUoXa9IZ6lZ/irjzvay9GYR51O0xY
GP6V/vhrsvBhR7mwO/x0eZBr2XkwzUBvF6oT4ebxdjE8uOvxf5s87gZI13FL
bdFIbg5zvx26i9RTueaZn1BMTdSmVu7GVty3z6h7/r8xM7UtXGixdAWDowTO
fD2nQECW4kYQsDFVl+OMOm+CzEsW0G2YouQTNmB91mBmiUXP/S/eNyPLEHU5
nUKrejZotJ969+pl+06S6JI5Gi1j1qUs41tSGNZN//AnYVy4uKGeeuQ9gYyp
N+yejQoVFHyST4XjPjwr1QVM+atPK/kZ0BxU9ASYTPulhHRRh9G2ZFrD24rE
d7hKUHAATizVxFNXY+cGeJTSLYJOz6aKxVutlYnYgqZyMA6c00JE0+nCTZaJ
p5GVRyNEbzA73EycscVEWoFScsC7q9EuiN3iZp8t63gnGsSitTAfuRaSjIsq
dHIAf9Q4kPv6lXfFtkEQz5SPW4bdooMacu6HL73W/7aWleaNuFHjngXOny7N
HkHrW8V0nZiS+iyiLVznTfK4xRBnB6aRmycVQIWYBxGWHZCO+1zzpXfN5pIj
Y3OhbWwcs8M2RTMQzOjOK6z9r+6osnuZoSkD7dqgQNB5B0eYPIXnMZrBlsTK
cNa67ImBqiQueuEiett6QSlrM4i1vvczw7CCQy4TzH2Ub8lJpncBsx2IGRfP
unEfdHTDzwLJTY2dnox7fRKm7sG3v1Adq/yK1ZUTt1iJYceDMLy1q4+8Y17w
ACQu2Fb+rMQQp+YutLWkPYE0F5/LZ65mZrk0E/j26ERRPJJ4skAk8VIo/BoN
SHHm1OELfNCCqIXvKI0uDXBpAJRo4RB5fICbbZdRZ5TL7U9KNfhyTxsLMfpm
QW0beQydOSQ5aJjL7LndgTiqF9NN5rBrwSVWWGwwOj7KNE/IVVbfW0JEBxta
lWI8pEaO1SKwJoGTlihLw0yxSMKLK9xhq+4uYAvpE5wsc2sGrW3F6/P/3BaC
f4t+P4EBc/vl1oj8r1poes1h06xZP6rtHtme6JEE4qO+N6oIT2prCmW/OLR6
6e/IMUcJW8TV9kJpUqFBqOJG0UodTT//oyar/r5kYEj2N668kblFYscBSD3C
ogTACw7N5jT61dGECb0fzc5tm3ZvXg5HssapULjYFR1bzykQWtQCSkgLhAXQ
BE6U2x0rQE4/qLxcN0GI/PLYwL9CqzXTQdyn77QpY88OEr0v9zuH0aJOHWdv
rgrIOkEBZOS0aCZujVT+cNxVt6g6Mi1UetQynuhxzqHGq+w8oNssKV/yAaqq
PpXYrC19g49fNxGIe+hqxdV2CFEa8x8eNsfexaQ7cLMztU3if2Z5Idj6rPnz
hBFIFXzY2953bz4Q7eBQ57zjiI8UkoCbCjZaxqg1xLsfpbAkB99XiEZAW3i/
27Ee2/il2Eq6KUI60V11+KCtyMUVFyMpFYUA4iJ0yCcYeyGn8Q8uBmq3DM7N
VaGrp6q3FVA6dZpGoC07mOo0nTu7xmNY7nPbJgW+AJB6TjyXOwHz1K6g9xJW
CYy06ka7nJ8nUEmCx4VKOhVTPyBmMF2bqdJgm9JztQyF90UX5DF9Nm1CtElJ
8mdnomv8vKG+bedCDVz5Mo953iAaxVLdoc4wG0XbsO07STjX+Dk2/Xtjr65B
IlENXicOcSiIT3TUj4DjK9bi4M2teegeVji33hYiVE0U6IiJQoV827BRdu4u
kKMNoja4dgOkUYbTjW+XrP1kuLjySHdS6naMlzFpMTKHUwy22PXHaMjQjI1+
zDq8lK53klTnDLnxoJRwO0vEiX8b5KFA4LUSrOK3+8n1ZPzduy9DkZFPGGaj
DypSEeX6VfTSFOFbdt1ZeEoDaNLLMxARcFEzi2X3vmSywFsxs8Rlf01c7rb8
diLGnODQUMePIQw92kj8MxRSaRgDesIvixVxONL9BqUFKSJpSrOXISaV5rIL
wFlYxoY5QjzcCeCVxSUl7uRxK9dWbs5vJgmau4+3Ss02yQQcvzpV1byqv1E2
oEY09A1R1OXI5xuscM9guXfWd+RrkoT/ivWm5+3hfJXy9774CAGI5AIbe7wS
KVAKcBBSZwEX9e/sQsswv3OEQ6eycwB2N+CNw41FMMpGorcttYu07z2EXJVt
eshzDJofCUZ542uIJ6OnLuxF/pMJ5YcxBPySZo7EoKJAR5QbV9amcZLicKq+
aoBKBYyXiTNNnyrdKHWw+IQR8eO9S8edSprNF0Yd028x+WxLQ4ffciriFkGt
rFRKep+HHMvNIiLkQtJA/JhzguTGg5sJPjp0hiBa76NigF8qaKhS4YZfHosl
kAbASQ2na57zMBMHTUPLVn4Ctis89rE/ctPCxkqrBLANirnQXdl2o5L51Io5
AewIq6rdRklebd0xds+SKf4yldO95h5EITZo/2lJb/uuO7Gm/tVg6nubyyQS
d4sUQNj/qqTZJxt/9NHLpDmmg1Voi802WCmLtI2Sq3gA/Kr0ZbieCAzuLwRN
N9V1bqWwM/3NIljMb/AfFLAITvu6h62+taF0XA8dG8I3uMyTxYfCheSmTlAs
9ZqO9eAuZ2xlYHFy0EfS6Xfp/RhKnC2ZR2qsEhxRLJNfLcFQ/DN9NKL878j8
GzqX7hFWxhR6S7PIl6KcSVTxrlXyugRIsvFdnJp4JjguDvHo1y6W2mwKQnch
LI5r3smypOGB7mv3P0L1R4tjofIgamgK8mOYEWtOOlO9rULkLONsEXmXl7ub
ra7XUucfsD7lwldJntQUC3PNP3Q1LaOyMcmS5At1sLmwmrCPUxXIK5qrChP7
QxWIdNgd+fQ0DGZIXCRuyEhz9XS6i2QY3HRXvfFeP6mJaTyxv9dL0e7t+88X
ReJqyc8AYeM0RCXznyE+oq5JzGWGmJF7vzOpW2fO1WgnDDFqw2iRoUKHxjdw
k3xkZkPXbmVExU1LaB86MixCHcYlOla0OcN8qbU+0KG0VeL1p/KTyMy/tPLy
Nu7ZZ0tgj1XxLu+3a6kzyqH8uZ8VxRUFFPoFtfvTpPuiqWOQams0Ubwww5Ab
9couIppAQLLwiIej1eHF3nWKEJYfaIeYQdfT6fLDljBZeCdcf2U9Efq2VHmK
4mFVz3fXRFMCBhht1VdfaRitThqF3smgFOayeNsEWpKFNuPDHzHuiAdjCVau
QVzk+4h1Pm1zdpcaTbuNP2JjdXnrfVuJSFQAkcA8Eam5LauHjhz+k65VtF4a
DwUVAZv8ZXKmsXe8cR27eO8rZUpG40nq0vkIDmUUDbtUTWzg6fMr7bEpV7BL
y3o4IHXvdfiJoG0UckS7eUCZT54HEfK6RqxnDm88aFJcuBceDGALBzDAePoH
wYexj5YkTCOoMF0FK1aorOxxckpruPVkhE4aLoVvYnZBNWuucDCRfo7jyBor
dnSQxqJG9dVVf84RTA1u5Oar61U381ID77de5SWaBfRaHi7rbE8bBoJlQ3vl
iNM40WyUy3bkV4biwrbCyAx+ZTxLpWJJzL1pJ379Ti1VQchtIrj3Qm/qhohq
GUv4Z2du4H8LRBMxWPJiEfqUW8NmxO8Xf750mUzc3wBnJPHc1t8UEBmTzexE
oBuxGRvxd/WkhViyDu9XR9MIlEYo4FE75JJzY79uuVlkxTpJQcq3h4f6Jv8x
G1sV5oO2wnsB5/AgNeN1Zig/HXX6zlISbvvXqBpZsQWsmbyCwMOOKHOg22u0
JQ4mgyRK6MQi4hkTxZOXKooAqDn9VmMGZMVCg0TP3HJroyPSjzKMgV1ZuRlC
5pKa+B4sjF4iFU7zwv9ryLmlLiNvLYteTe91gMJyTqRImyNcTs+RmWGR4RUr
7xOHcEOqDasEf/y0+h5ca7Gqpnx8fHlnPDsJnX8Ph2WYSso1RpnaZIgnBuL6
G6rAhz8ba/jSApGRiGDyMlLty3KavSzRvQ91sWMLAeHY13gpb8t6rgeQxhzV
oxj25SZ58pWPNG2kCU6BUA74dPmo+mDxfyAF7bm631PWq6TmS+7lhUwbpuJj
Hfo4gQMncH2ZMAmO2g3ZzDPexAAi0OqIcUkvqdSL0QcbypnzbXZ+s0hJg6dY
DaMsYzwmeJFIFsmZTk3R++2lu4eQRJyfIjkABYGF51llPRMMx+cLl+P8EXuR
Zct+0bQsUP/8buwZNUU/go0pA4H/kIH3XJswSG63VeapXKm4XtzM1MuCZsR0
1RziRyG8UpK1AUOovWSpYfK9vALh/KhYTu5EihxY7jS14cNeW4gzdEVKE0B1
/x7TAquS8Hd/aoKMk7+tKG5d34DtzyymRRsURcp1D76epqz53kyWM7V2nPPa
71hjNvnNbVNPzB/kjfABLSo+B4FY41MP2TlkaAcRw+caUmMlWGeViorJaihV
Te/oydg53lBW0nlNtbw0BP9rLfzABIYgWxeApuKX4UKW9CKZ+ojF+IL4yp2E
HR9Shh3esC/deZMmz57Uia50miYHOh9DXsTtjkFzdPatNJ0c+QsM+XB68a2y
RKZR2f1pw+rS+mVGhGhy1VItuYA1AyrNcJ5N1GSIzrCmcD7aTQaqkTBNh+Ok
c22NwJXeUWFmsLi+FRG5ma5JiYDxgPN56Qx4E3PWKifOmNk7mQrSWkiMwbbv
R3G1cDxcitEzfYhVYjKiOabgwCQVLZ8S1nK2sySWBj/0tiSgdlrOSdITo+Gi
oV2kblXIPrrksS2dzSkBZGluNMYh1oLz7418x7T/yEsRhzy7zrdNMoPQ1Bi0
HaHKB1RrU8iJ9SEiua3ydMQfEPiusoSJT4Iqzq5GKXuYA/D+N+VXaetASGM6
EsX1jjvODh/0V9GPXpyW9JlI1C8bGLpJQjdeU8ErYBXNurjq+AiD6RMlm1NU
mAZOMHKmwmkNzEl7GbkMkhqz7NS2W3BZXtXYhRc9BhUDIg39W83Gi4RDFA5O
1BmVB5S5LeZteIwax/SWX8uIRDaui7AUN02aEzR3JnW+uPu+LGmVbu9cIeyL
RQ3sl6RuT1PFvaOXK03La4+v9hYN4ajd4D1eTqbgU+WX6EV2Raw6RZV4yHNX
gVvOCYVag/4+A5ICrEqvkks2kmOyq5hZyyhOgSVZPL7U7xonrTBj4O7UfIEX
+0uVv5FrTbJDBfAZmng6akVEOj6vNUyILhTdRobZ79EbS/mZV2/6JCSwhh8R
ESirJTeljtcIXW39gvif3Ue04zQu14k076tzOyqsZqkI9egc/yPGdkLJgDUo
Xsdl9wdsYd7UTh18SyLxo/wZKQ6DXUBdX+QwAHV5MSTg7pKR45uGt9VXl5Qv
zNro+SofMfs7d+95lunyCUSNT0HB7K7MTiEt3mFIEDZvt1SQlmrw5IqsmE19
/l514NO6aLzPM56Rc49Uwtg0a4bGYo0uozKYH7jCemQ5BsQkTgDgOTkFSP7X
cIa6MU33gnxC5uRY/UB/ESUSt7OW8jtvu/hezBbf9QII03h5WhTae8MPi4WY
5aofu6QeZ8qvt0gxv9qw7x0txDgg0dShjDPHVCZ8vay69Wkt+QdIawd0Nbb7
HmS+3cQxoY3QOkWDl6hJsCcfaDeBNiqAhqDZ6i8hde840eBJRJX+KYTMq+RM
JXWaXt6YOuvHSEBgJ2j9NAj/oOyVS3/sUlCF2at02BBemTjGPRhK6p5yV4KI
ypLtchgJan16gB1nHos7KK/rFljOBHk8INdXmUu/kp5FsL98hPvqJZ3SS4iM
UCkDp18o9QprnKrx4n3/uTEr9wt8euWhz1CiT0Pbb3whGzn1B7hlIKJHf+iR
BMjqiRwn+LL+c99NoBtRv66Z/ZzJwFG/G/XP6pep+vsSaGJTjEJT5cdtFFAh
+hiBYsF9lGH8+GCaRqYKXbpVtYyFK+jhM20R8351Gq+MPfrjS+bwiDeZm0wu
h2hv1VD1J4UgHbBZYV1TIUFXV0lQRba+yuCpu19ww5e1zolOhyuLo3FW/2MO
47AEUKfiI+iolTO1nO7jTCwr73JpgJptejP4o6X3/rDWquV9hMt4RjgCYmjy
u+qVcHBlNzxuEPDcIhklZYcTFFYGnW/rc6GoXc6zxN5qauCnV22+dtO5EbeX
oFH0xgUggg4iDN0M/fVcJ6HWE882i9G2xWTN+O6DD2OxMn6F0/7Y+k3E6hHG
HW0TrRPBPshjRJjBnmyRj09DyKEGbDMq5665krkouY9ANy7bgKKXqPlBYaYj
gs2PfuAbz1u5tPmTJ/kYymOJdT/WCYE3JdMaunxvW3muOPWmbVAxhY0BqvFk
6u+EmY9ewmLyYR0YVGWq90zkTUlM7Aa6ISTfcqZPkPkgZ/hfs2R8wrlygBjU
pdFUC+Wt7h6Q2xv0Qqbq3jbmkMKZtyCQLnvmPP3yTsseXmOIzBiI77P7l6DJ
WAM7kXya4yTimaN6QcuT6OfK8QhNaizrTGYhEr+EoEV1+ROxroFu+OW50/qS
GsRN3uAkCMKc0dicHqOukUkx2daunL6+ydRKDYDxzXIQn15NASLC+aoWMoBs
R3uHzEgU+i14eKwqTgmvQ3nCgrWzkGHXoQ2IfbenFhyp4s6O20G0naGVa/PB
IuYk5fbUg0RnnzIH1Q7vAP7I4REwjHUGYBpR71lTdYBelFMkIH9Q1HTxD0Ex
6ptn/W47mfHwvgNTwzncvlxTYFvK7XDdbzb6nd+c58gvNXMUp8mbswoonVVC
cowbeXW+S4GkoQoznn95aQKVjWLgw9LKOo17KGXHPzpR8ilhek9CFYG2KLi3
kD8dchv92ChaEVnzctmSLZQF5Ouw/3L/mcmcGaxKJjPTETr/imlD9t84N6jL
9TaQ50+UltmrfTWkxHGJ/xqQ22cSIuc0/1vI/WPEw9RgdZWlZ/IaOEu98JZZ
iBtENocZ7jlqwvD0vGpH7misvwhpz0GILBYrHvY7sIvab8/CbN7AqxI6r7+/
Ns9gmJHorD8C4qnXFGYePEa7AyZZe1mk2SJe0ID87ZOov8ij25YLKDlvq9kF
++Jo/CMAcddg5pcseHrhYHWW1+LNK0MHJ2DGjGMPUL8mvYEYO39li/u/5J8L
Gl5zoPkIL3K7+v6t2V90dq/IfMkO53AhCU6eh2jOVsXdxeaWDIiJIspJ7CFQ
o1hDT2aBLO8xxusGwFkkkF8jvhHu+8+BnR6H2JvZgwern4a9QugrvBwj5VFY
HcdRkNr2J+PzS5zFqaHPbXUonTuXCudRagnVBr0FXY7sRpY+G9J+mRV3ck+A
99XfNR/WiJ/LEIRHFf+Pwswrdzm5Zzx1eW98CVzBut9CcDttmC5ytv5e4mH4
Rv7ZJf4NnMNkwXxItzuWnaNCpjSFxBLHjcFlL2ya7Hc8mvZTf/lRlSGVJoJG
YV/PfpDT+IEfWLN63BGnMfesp2+OujlWU5d+gkY25KL0/zMBt/1oTFJ5Fh3j
6IchTVOihVi8EtNGVGKkt4TjqVXhEYtlcgwkdkhIyyRGaV6Az3p8unNvqzwn
zldBRy8KAhBPRtse0aNG1njOQ+LVCzBsPfBT4eaQ3HNF6AvLYPc58T9EG+f6
9TZiPB0TDv5ZtHynw967UQqD4rs2QFZ3ItbFoLi1m/4ysM88npizRItCksI2
90V3U1g4YybqgP22i3i3Q1DMfNE1Ca6ACiLTGPKwltMgypyHc+dLOkb2AKpj
tgX30tY1RjFGpi+uei2keihr7fx+QV1NUZI6iSHlV+unUOdw9VNPL78FExSj
OP6UsR8tbjJiJcTk5mUcqa5rrC/KUphmrDZcGNOiepS+GWqTPSwUhowNUX8o
nm0skH2b/gNhYu7PIdEIiuGppmrRfsTUpR1+sOEn95E/p59peaf3r/xE5hhQ
rGbJrS9uqr0HOKNtjZKzVdCUErpC7dX8tteVYQs0MAYvOfpsYSgzdnAkbXqM
joDUiPxfJvlFjL0SDCL/CBMkgohQAIJJiK0FfifeTHg22lV0CCu2Rq96bpfI
NP1de39t0OPZZ1DgyDPdLMNrWr/ehEfe3X+5k4KAwDSGSg19zjJnQjr4UkHg
FwLsuYH76jWkRART7YVPUnDa7XwZDrxs4nElYEmoW6/kvgySmUcUdsj2VAO5
ujDqbacVhRY/KdbFtdx/N/51K8txkl5hA4Ty7W+YsfrnLNE9dW0wuAY/VoGD
FEwmwAZDn/ucsYuFe7p5qvP0Gop0WBtA/gzHWKW/KUlZtqtiTJEdf4Q0jaC1
7bQTnxEblSRR354/UJQVFGPBUcQTAr7pyd/xZkOae0Dvc48JkTPo3PLLH0r6
9tmekTg6sGcprBh5Ku6h0hJMocQBMNJPBiXZ++AJiGzE6VxbOTEpH0LOzuLY
qo9b4aYjeKd9uSKf3pShzTpHzad7t3BewH3zgEycx/VHcA7YXjh1UfnWYyF2
qexto8Fab3We3Wv16anRHrzWgBez+ws+cn8MuZovQsv21KEU830X6rAxZhwD
RAab5iVRIeLFXEV+KTlwOTmDE2ojsKoSZm4x2TjHHrSyvtSb4iF5CmQL5ZQb
ZoW2DrmrNJ++yFbl11c4WXNcge1rL/SVEh23h0EP7a+f71fG8YCEXaQvlsQ4
gok6uv1yH6YUQKxhxVnW46nSliZX5AiLUkafffTsNiTIIRTxtJvxdl7uqbSf
cR2I0VRTVGd4uYPGgHQEHAaT480omJDf501VFwaVCQWND0NPMwOct03m7c2e
UzaLwYd8B7aRZbSbdwk/4FY/xGAlessyZWyTqeZRB8e3LbwkCc/GI7YI8uiZ
2WZ8bFeg1DAwdedjTRCpy7Gi/4h/WbNZG8Gs0uSKUK2Z+eTd4FWlbKwjTFPQ
nEod6xGbRTuMmAdI2rpseYPPrYM+ANKMmO9UCf//0UHAMGPhlxccMS4EjQ6M
rAHAGJp/JZY3cUcdzxBSn+FsoQUeu9aUn/+aXQMu0d/8CFlnzS3vVoYA7S3P
a8+kqLxTmpWV1NFP3qw2E2ln5klOzdT9Nal87aQl8mhEm3AZHlVxmuIET5O2
L/D6PJxqeKJR+Q84vldg4UVIadKv/NCH2SaNkB3BJ8Fif60DlmHKXavCOWyP
66srXGY5gloigK09Rs947y+dYmTRM/tjGk37wrsDVix8Y/II4twRAkU8VJbX
bwOqik3EIKvE/fGl1ZkJJ2wIq1FDvLKFEVnwOPyp0Uq87ajSFXZaE1ndc2Yd
QOjTTNidh+zHmKYyWFKsbm9740pzhblem9j8gfGVk8lmvBBwJNowwg4TLUMJ
9E4+yg6rqumYOG2wT4g57UbOXj+6OpoolGX8ybFo0fqqQxr1uZN+VAWYzaob
RmW403950AzjBCyZiBW6ATEfsUzwVLsDjE3jaFONFXLtqB6ZlHDXcIWtuJCp
A32MQS3cKw42bV56p0q2QI2V44Wi8IAivVzBTs4J8iK8vnFn1wawdGb2V/21
vAvnSaqQ/xvPcMVPa6bf5gvdcG3/rdYJ4awKtgyAelFlEOzl3TKzSQ93t5LX
bK4N/G/z3v9msSbtKpz51XYTyNVOtQp9mwLMvHsyyd13yYJK6qpzXHTjfPZv
esx4spl4XUbYY0gR+JlhG5Vkli3RBVROWRV/kSqQMvzmzvNWK16YO+FA3az2
1aJ7AlewQ8upAKuE0wRp3aigT8g60VWCiB9cbulGCfHZHU6/StWxhE25V5cN
JXZaR2A8qqc8Ag9ZnZWzApjErbw/DKDFi4ou9SqPWluVqET1gdsj0KdxG8qo
myqe2pycSCw9jFC2bya7KVVVURlBiyps8JO9PqyHbywiMBsU09u1CeIQkPnx
lVVQbZj19EzswuK5ecRFKai1PljiEhfrlHffQRaGnlaLepJqoPM5PXHODhA+
6l8ypvmPWEyOkhPT1yH309a3h42O9Er3zvBe013G7HbU3Mb7mqmj95Mt3+Wi
KxOECVcH782e3ulInOn0gjEbWGpnv1zEjJVCrcQILOky8CRZBRkAQRU1yS4Z
6dru6CDfkdOhQHJuZh6pZ2bSy0ZORH9sThElulV1SNwCxg9+9/LJ7X4hgput
4hp7//gBOY4O4hCJ0ShT7v/PdzH6CqfNgeON6tWl+DcV5a5WVWk7c4x+pn3C
n5rbrSejaflGS6j7DGYlQCQcJdcW+xfmaeE12znZb13Ij7Fbr2YCmMqIyF1r
T+qY73NRvMZFA4jweKwDmhG48PzkjR40F4ZqCwOrelYDn4E+8l+B2DYcbTmq
5hbhTvKT4/rtbz59M4bHx1Wbz/bfCY53cN9JT7ABJ4PjmMROG4U1y5l4jdIN
wr/dUA0d8fFAX2V3+63ve2ZwX3JYmTOyZxTezgUmraT5BeJ94z+9Yppz6iYC
sas7halu85YYl3wEKGDoKBge5nmXHmiJoRMeHdCUNuiARR4hiyaUp092SRZr
6rmPEvwho6vaa6R4kOI+DdkIv3Njn6NY3B1psOlhssmiE7MdQvc4Z5L2/bIS
qEp+m+ZOlZ6o+rDgJwhBXeXAqxrAgB6jFxL3OTzvgCGjEPwUqMwKAgUxwuIs
U+3KXHcc+cmGP2NJsSb8MEkNy2846RP5+vniMeeqx0CFiT6N5jqrI3p/kNjs
mly036w1FMSndH89Ujk3fptovGJFHjbFSZErNtBbUEsh2MO+KlfSWkiJ3JyN
PNuMvjzTN7RMR5Zn399dGcngPK2HS70IAW1a6uL8q3Cdx8r/YxexB3Gej8X8
7Xl9yzhNuZm2eHXXDLye2gCkMBMmaRRQsQBRuvWGqu61VvSarvqDBJmzAv+Q
qeISKFMLCW0QmpQ4cicLj19F5ywpc/8dDMRjpUa6B/NtzCNxW4wmE/V+B6L+
AMs1h/YLymsXWC8ej5HgS+CGe+EjUQAbyJ6H/3pnoVJE/S5attkmXiyi60Ff
yuZfYpbCeHWxQ/9yU1pI5GwryWQzAuUILbY7ejwX2Q0n9KTv8nUmojrdRYRq
EGr2BnWd5VHqhOQhWRcrLfqZLKjc+etT/635xjz+LAMAaFDVzq0BKVngKJIk
W/iXVcOQwaD1794hFjpsmiZz2El114DLIuKzjB+vNUfra+//JPB6jl9FPeCa
4BfvXSTC07Isqt7MaSjR3DuWN50GTWSrjQD+gzXhyegcPy4M/B2HNrChPk2o
0mwuVE5ySRvedbVJcy19wxAQQJNVGhTP0v5JF/GEFk1RvjlJpWj8KkvhFrJO
+4cPDbHzGZbjBGHdEW2V68sDyheIvj969mBEY62lBgSi2XDF2Ayn+XjIFDdG
vjPUEioHAYpamKJPVr9tlRzAnBC77g6LILWV7G+AMS6380fE4YixOVuq6NTD
c6Oe4mRP4xGbfzikwep2jBtiZr9zo8XlWxB6YrKGrXowbJiFYc7pVV2hcd43
Js/eKD9nEE8l7ceROX3b88Pdtu/fpmhP4M8LG0Kwjp1V5QxcFoZUkvrVFV8w
TrVKAoyrWXx4vPRk6N3isExw0PwPl9iK0l4PChZQowHV4q0Z0CgOoXICqNyu
hHd6ODJRWJHJZm8DDBReCt1elT0FxxnZI5PKv4ZdlWRFS03IHasSE6b27ao/
fj7anO35j4Vx8CYuLdL2+I1pRAOJTD/TSsjyLkxNcO11YzYZssV9ldMZV8NY
jz+Mn/HUiuXL9pCCXe1JiWCAaTkF1rFH80hV9vGbhyBvyXt1zMXe1at5niQY
33Ri1ZELJ6VjxDfYMdT+RdyHkqcxrRfN8x/RsG67+x0GRr+xZHthrXsXL3Jk
pPF8Bh1Ubnb7gqW/d68MjjggcPa4PyESMw3KODDo9XlNV15Yd9w59F6d1nyG
yKKhm1NeiJBogO55zrfz9RAovM389t2o+9ysdagQBKwBxtd01HwY/dZGUnvh
qjKhDshQRybh1nMfDrFMzPeYxu6sSEijgNKau2gyrEXVR4EHdFfKKXGz6K9x
4Ny63lkwbTnAMOW/jdbS36zNjngaONRny7kVjDEzTFWESW0UqdmcsSg/jHxD
KhC2pYKVYrlpapo58/swqMnFKuLodZfRZZawGREP/92H/KXiMErgYq2QvQjO
d7E/F4ogocwczvUNjq/X9vIfRWegjYiBVrSt7FA/5245SGKhBuYejHanW52M
wk8M6rD9kDp8DNIai4KJgva/wsHwF3cVjhjBmxl1juaQr8UaqCl5f8QMqbcm
jhYWqL0lv1V5y0Hogm9ZEBggkGIC2z2zkJncaApkGP+b94Ie50eWuTSO8RYe
+hQHTHVak0VzqLm8ac8V71lQqc91swjiRbwRwR6d7qY0kBQGN1AtNQXvMROX
uKbkEpYutNCEQWXw1icnxZ4oGI8sgDmq1XhyVS3w/u/EgBP4Kcd0vjw4ah58
UmqOEKhxafZdfdeEn+5jeHHlg501x4nbDSeF9aKRbXI36WlkCtWJ5WPiYMWh
sLu8RwfgXRev+Ax5/ayk/+v8pvGJ2azQzzkO5Y7mTKyAlk080kZnW0YM34x5
CivX2nyxvJ2jVmX3i5cDver4wo1EzHi5FccCFJI5+6uTgD9mCrIfBrEQS7sK
qOlMqnV2+X2AUjWd3uqhTIEjxpPMgKIHu0WJW2OqDPcE4LOow2EwVzAcEM9f
1vkvQ7LXX6HnulMPZyGtSZiZXlDhX/u6tFakE1T7V7EtL2WlKPNOh9ZGjl2H
6Rb+Fq2MBnz0WNb/MS/08EthBoejRnXuhCY9fRANME7xlwnJTz1sRIWdKijn
BvZoXZSUtZ+Qnn8pvdi0+NymB8gYOlC0LNQTJLlGL3k0yc5gLN7xsqMFneCf
GMsyms7CQU2T4wthcpeALezQ93W/+OiLqUefJD/s5MOk683oYqMOVKyEHsrX
zk+QR3X/11v+OVqD9nqPr+xC43MoT/DZkmfT962okrCrh5kdb6+t0ATG4I8u
b5MKygqmn26MFq+12mZMWrm84H18oh1Jg63o7HoTgrECRi4Pm+hfkKXfXKfY
bqPoKqbjZYBol9vCjJWuS5Fy83/qMGInC33v/9x4icYMdBYI4WACa/ky8vYL
GD+B1ATXAff1p/ccP14dWR3NpF50I3uk4tVC0G49wKNqSahj85lyW0eq8G30
6JkCEpYE1ol0quy12g3iN1f//Kzg8AZhyomlKXOlVOq9NuznLWKsh1pwx4Vg
ahXibFj8+KfFmmuCbx4kuOAZ8ymkro7rZao5IDHqw+BBH0Z6YMfy/Mavn0yh
f9haupGp43YI/yCJ7MeTN2FzEuL6f+Xi/67uWhHT7k/rDKrzsS0jIbR2aVAl
hM3Uw26j1/NeKvGZ87ompKVez5hTB64JA17sZ4Cral1Rt/KuMCVGXrxYQxqn
0bt9qYMMY5EOpimyTPneqnFZKMwUjRo4sy2gt5g57zYMu/JYAfDMg2GuCmWQ
0b+o9b2IWoCTB19YvnvuI5Ruh3VsooL/Um63xBjc81tSkyq7yykboW0kY5rG
T+g81EDvMHUiP00gQBOVCmivxU08ESPvH37gYcY2UOs2vhXBREvDoArBVx3e
Yuno8staBOQnlFqFVykHauERZagMjJ7FrJsNVJdPmFa1dVKtgn8pPR5HZ89a
x/0CwMZS577mUCjjyFHJHjVLhmaAnn7Rk4CAO5Zq3WPHR6y+z+904QqZOT8n
nPybbKRJjPv22Nx7yxxcmKEM+mjYjczjl9GJv5z1qsyVgyAzhMZjet2TtTJK
tdIJjuOECJsxbZzaBxy5Qo7gHrcObmTfd5i7vqgBncbjEfFx5FqSbvwSiFqm
EugT22gs+pcYLx9KKpZ6fUvaX4uKgGaqCd6MnWmt7VXwAZpp+Q7glCN/+Rzz
IZ0FAKGDxQdMDDJIlsLlS+4BzvmJeihrPcwambDjk62OUYZM66S5v8dRbHSo
92tacCJql0nVZQIkDkMuQ38eD5UZ0V3T+YJv+7rR+2pjZwwjszSWHjm4UYGH
zRrcaYUu1BeybEvGriu1Q10+gquaauz6VpCrHW8n6fLi7BYJZrcuHF5VPdRX
Sc1Utd7ORm4hWs1ocvGAtLPGaY1kv5je80Arsiyk4kTUepbGKADgIPqrUUJS
gU+1ZATMSCbt7XA4ZXmOiC29zYKz5kQkiHlePoVr9Z1FYt1XC/+EvAiGC63H
fhsMjPt2JkXi3Ld/YpWSawWhbZ07lMy2cYNHp+3SSyuB2X/vUzgEAUehs83B
Yf31arxUU5D+QVYB83V20or2mKVcZouKfBlQau3ISsf0oklfeEVZ/vxkUGNO
CJDW84d3IN5CJzNhnV+9QmpHwT3fEyXhuaJSJ5ZwX32j+xJloD/FRQm5FDCk
FM+OyPlYOEnpqXTbuqypVsGs1arZlyrO/BSCdJJCMmUVOcMkIl0OZz7PxGxH
poJh029zaj+V5yU6SQLlgUU7yAe7OjWVN6/3Ck/rHBxH90uyMxjjwWmkOAVn
AsQGhqXfowaoOrCZyHibEsXUVwTpu6Prm0u7LWeXGgytiMtjtHQSaWUshvKL
N9oKvYYfycUhY+jfay66fZxfPn8ikg4p0dzdSKYwRTmjafY3kM7ncJgvEDwj
nqhTvf/IpU3FCack0A5IIJLuyGh9QSlSQWAHyRXIYbhNLdP3plvGiSfe0vqF
y8ritZcODxDYWh4tVVxdSTDKLywY+KkaQw4HK7PSdJ21Crc5sIwDWHojoV0v
imyCtPC8lPQs/fymNetBE9oLsUd1Eki2dauOKxjRu5xeee/m37/IJfsXDJ7e
+QHqUAUvYoivSzbsHxkqyPaX+tTMcXfJbrzK4RmLWgydsYBI77VIJ0cNYgvx
VjPoEHEs5iS2Hcd4/0fT5uCw8CWM/3qWuidFohnNhH7dxRzRy18yhfd2bQLP
Tlu+frSYk34eVXdI1/PyT3pJsW8sG3Xauij989Ecub6bYsjv88n+AoQSaimx
sz0qHQdyY8bN9e1cAT2uhFqBA1YzR4FJ+V75G/z2STqRkkA5ysyW1BEXw9E3
GPK8PAdyOHf9c9gH27BFSxxcAfI5/yRomt/hbMaaYXErIIMF07PJ+/fRmFvQ
JSxv4AgxCRLZC32UorN/zxiOV+oNXv/vbYVGY0XSKsaNxU4isHYhDE8WstHL
6EvsqNslFkvOCNu4sCblTNxvFq+vbq4r7swcHI5p9ZMDN1PQ+VJJeXHzANJj
sjFEAu3zo4+/ed2q7pvykFlqpdVCFGe0vhcjK0DiWcEEyP/Hdd21izYTYvwe
2k7WZqaQyNTK3n6Z7jvJakLlxr9hIoBZhC7ekbO5fuZ+hX0XuALQZ0tcQ11/
mrH1Yr91xzsfoF4Ffi8SZEdWHvirBB/KIOceXHecPR/vADEhpvO6WGCTEHmR
R3bSYHDxAwip4PAKsi3bVudOFMMdcKc0Pwih6e4NBPPLd+s4hoWpGcEpsf98
STwJ1PpIz96ukAVQrQnPkA/iGrsNAOxbTlWoDiMNEM0r6ikWfOq4pJ5A5Ezg
RapONUYpUWU2Imim50gXCsrs7vvZbPLdnkr2ayWH6RO011vnqZ5RqPV7PZPc
IzFBqho6HV2UM2taYBdW+2dogvbMlax9Tg1mFg4tQ0CzcEMbbYstk5akwT5L
iNQTk+/3Jepnflylzq/sMCNeOP4aBLpizgXW7qYEU3Qg9mVUe3dOs6bKu/PY
STb46XVO6oT+oqiyu5ujKocANMUifXAwNoxeDFIG+IJmI6CTqCAxwFOidv1c
Mqr8oTxslErX6NDRTwWXiennJ80EoPEF0qOvMECvQLESaDeVaPNxcB4ZqbdL
aax3Sm/+AYXmKGflniGku5IMGr1MfBvdbbNgXA7KOK71VOIzpzAO47H4JsEd
sXH1JDb36yYCdZnqbF1HGxjKWdfZXjRD45g4rBfyme+5DfvzFKKuhKTDhpuS
l5/FkmAM5UxHzRsNTtH/EkQ/8QOspiKyGlXLNMAYEtoKfOtFtraNmYQkFZLP
aZw8rorHD+H90+QDiihr48i5j+FK9ZKwggtWoRFDQ9DIbnBMZ77Jk35VS2//
gopJpGY1WEwdiyoWyckXTrYJfmrgekmx8Z/Nflmoxi8X9cYTGrukCu7BeUQS
DQjqLzqp8tqbYwvazHXM15bBjtuYmSN/M1X2JNy3UYMCl/iJTnFbBwn8Gc3Z
zmlBBvrE3RApMp2dolewCOnv3v6G4mFiIfMgdv9LIV81YBiTwwLABWSb2+1n
32daB8P7VnQ5wXtkLvLfHs+KYM5IE0iR0ytRMmyf7MvtT9W3nWIraW4bv8Fj
aUUhhkO3akc7uPmCzRRdV/Vfg/ySZsQ0DcRM3cJ7Zo7HcgP4ld1sNVCKbN9o
40dyVgahzxCx7ptgPJrtpSx1mWzT2GfKrXr9aukllt8lNcKNmF0/ygCBLAdY
VyBFk5izq+CTXc7uWD3kviEkSt0WoJljdQyr7a0kkprNkomAltst0kDyroyp
BEGCyWI4rVWeDTWvG4Dfy2wmLNi5g7bgPGWOzGMqk662YECvrkvXI1635w4p
NQNvMAB67UA8bb1xVgLedF35d6Wv3x+sUIjmTmKwKP4WEWq+Sb0G00Og2dcw
oydN8CcOfTJllr7aeLJ/L6vPRzFgb9kjo6Ag7dVzScWoxz5Scjw/Wbbuhujd
4kMAc5RqdP5tCAQd9ehYIOI5CmhdE4/hJx7RoSVqptzywfix2hiKM6+IJ5LS
Q9xlFNL4Vf84ypaGzXZ1Y3U/jXkN3NFihHpFoLzNZ3ghRKwln4qU7kL8r1mF
sNWC/N+4vCjfvOAYtUx5hCrgcQjvC0K2nVzp5HBN3vSOVqmJbF7Elsnmlo+G
4MCr57U0rRLlqzXcjJ6pouwtzyZ2aEXfq/1u8cMi+nGCDW4lRqb8sKQfIMuX
QeXaLlYP/zDXScO3Lf51xa2hA/ns+ulZAX5KnyDd/B0GqAYj344zt89fR+D6
yUdORp5d+XtKH7cEqvnaJXjdKqA6vuLzP8abgCqKtVVp6n04WDzOysmgC/zV
csF69kP3lZFKukmYFBijXnMYRrJfIPZgBfeDjNlZU2rjERonvk2YX7tZdz8o
eDarCiatCZX8+hxa09GZsEifG0C4rwM4z9npITg8E/xgKdJ5k7a0eSyqUaf9
37lCYvxBQ4QHh0Llpo46XYGm0ewW+GpRzI7xjrkKNt0maLCEkGck/VQ6pfIg
pbORchJX2xs2CqVzDRJ+x8RjK/ASEn1rasw/8WPNfYH5WCElomte0j/HxbMv
LHaixNdHKnuxlrg6Zcwh328WsY5q151gOkgWfLysw9hU/cubIQIrOopHrXae
owyu69EiUahciu2N9x5OwvLFW6hxneab7TCkUGSUOhD7j5Iv3HkBbpjr4a5w
BckDtN1i1G5F7/Q75bC4QrEg1U3sW+qxnuw3YFf4naCMU53QvTD6e3IdnhzW
frssh+iw84AMEB2dQkA63sq2CtE0EjqaRmq3XU+IYQWOsJdqHa9mb61V7pxT
JWaKzlgUyLzKqx243l5MDtmHu6ib0enLM1hg7NrxD04m++xq+mL0KmgIogt4
+OMXNGmujpJ82sqV0Kx17YoJfKI0SiyfM9qLttqGpefqgocGFlSQaV35OChW
Ag/eQ7u/oWzIArx7nQpWndAHYyY8uVE+P4TpeKfhbLJGtBGFk0SjgsQ7jvis
QkPnpK6fqtK55gqlLJ2ug6ExRD6rXuZ/ET0wCHl53rwyu95W43qA4uNLnq4V
jftf3G7OjdJT4lvd/BPs9jxTqjkm3LqouX8fuNgelR/hIViVWyk9UutoEQtk
xsrw0tnxr0G71AH/hSAwwtnrW5rjeRealwC2hplai/f/M39DDACLMI60Q2Sx
mJR+ZkP/d2P6w5MxRQ8N+X/UEeNLufO7R3N8xevfBpqBpHSBNG7ElL6l1mwX
GhA1FobD0o14lXr5YHSI0uLG8KyyGEEORXjwlY1JH1YA2Yt/13ec4FqkeHps
SmkTI7MYzDHm+7I7zs4ndtOCvuaSpWtPEvd0imK2LixsmP8wEeIhTZDKGQyl
woUPnumY105a/gCwfbvB2EsCtWSkgG5T3QPhihcj7fULCkRRkTB9lEQrT6zD
HAGqTgc0KQrXlADoU4q7SwcsiKMPJzUfEfIJdWKJq49A/cop2+wg/nW0LWzn
Bk+Na9FvCZ645dbupe0ynsxsM+AmzaHNQiaYmVfBc60g3choOo7v7SzWAFRI
2EGq7hyGa4nM3jlAqZkiEVVGl2DQ8KkuJBaq6hyek4nHWq2Z+mS/XzkkZ8U7
BfF+W+69ORa2V41BfdD/T3kZecShQBghHToautAjnIXS6xIYB2mF6T9UoI9B
PkZTOcY1+EhGatSXNhubxVxnxhFY7LO6Ii0D218mdA3n0TSqb+dkcjb6H3Su
i5gSgCcuF7B3tnb3uI7bNlVWa+CAvHi5MXAI26oUhZv/ZNZHKN30pqoSCLe8
cCiIwjcYmbJGsakJPl0ZVAcCiydllhAG0Q0apJsD2S0IUHL1FnSAOq+ZZq3a
AK1j42ooAdt0ysx8mTvXwbF85OWP4AGzeGQL0XaFjjjvW5to4Ld7t1Qc/kol
iny4LHFONbHdhd8FlV+KMxhrmyjCxFYBjkSCa1guYfM45/Z/Gqu120dG42Mu
+mMXl3JpVgFaRCkjqPK+aGvWPl7BA3oWRBYxQJLq7v01H3X8LenNArt+nbgZ
sj0XfcKAg3Ggv8wzdveVxHK+HdlIyxD9/eIqPpfsaWbMdDNdpCIu3qQT3UMY
dxup7+YWRQZC5pm2cqu6269YmBQf5JURGKfwItjgDmYJMI2IsRURMtexMXDP
UD1954dbfYoct3YTlEveWuCOK0vRJj3E0+a0ZE3GGReMt3q5DWsX6IAGhP5k
IgXVkYjr71ZFc1y2afbStLkN0IJdU9RKIaHxEYadtk4MjsbdvjlTk70DMLpF
9BL7A5HUUU/nf5UuBcSF+ZEkanI9ilfBnY46LOPM3iJmQRT1oaIcI9CSDAR3
sa49cqdrr9Xu7t2DtMZOf3eXfyeOCFJmF0/qbwUQ82IbD4Y0xYWfzB1z+HDX
/lnDGy6Ep6RdJAkoiu8v4D25/OYBS4dwozKWREDH0XTMmxRaBXnEZbXCgwpb
bctAqNOrxYs87IU4SD+asUT461jj6N5VxP91Au9kbgUf+Uz7c1JlLUJUNquZ
PwUE2b7UPIhBFOuTEcRMjA//L/JVpKZAj6I3lOIS/OEqiQ0Z8kj1EGwyrbPy
rqbYbu9et40gSJeZKapiOoY9nFlIuzSGccro9SE3GeMr9saggK9k1P6FFgps
VhRYz3zPUoJKF21XbPpjszFlXdzE6swz+Zb+BFV2kRTRMSlpfxJQFQs6CVMB
xR7zhZd7YGf6s9I0Vf2MUVef6OmmNdqc5MqKXba99jhewDyFtW9TmcZlbc30
n+wONb7YObj61fi5yG4qu2TouxDl7wlV93UXDn07r5uWHMrUkcGi88VfQEQI
/Yq8IsEgh7yBT6Xs1COi+/ehI4DfTYsrGQ8b1BMM5JZGfPfRZqD1pX0Ct+v0
/wmNUTHi43dA0KlDSMDIzISWEzLFnwG+X3sW7PF1Nqz6MlQn31itCbJPycPc
jYzOInEyTYzA+BdStss9Tysl0yq1w0KEzwuIaWkdpac2CklxkWSTFW6z1hBI
7eD16IJWH2rNdWkDgnB6DFPfg0KASxgOqAko4J09BKuwi0TJBQxF9HTKad3s
q0BTaUpiwSv/sS9I0urgh6frK/V1cXpO2cLDcTZSRmxVTbTTHcE/t4OM4doH
6GlgsFclFnkylh4McRZFWvLVPM0vgC80/0AT52G0hsqI2+78M82uLfuwW/FO
9VeR3a8/ursCu41tq0Pwujrnn72v5nMveKsHbPNrgq3vHAkTkTLJTRG7bzhA
G1sYWMac7QaEjRb9CvXjszJQA3FMPIU83D3k/iZBOyz2ED+Gt5SdNjQzJ5CR
0snV6VY7bZsX7Z0Lc4f591LbEdNNxbz6tKfPQDkTe977KMQX4vfCFm+uL/Wv
5d8UEmH7nPMUBQwmW0ndhySPc4HB2hhbCmcfH7VI2Kp8qZotehOk4ziVX/HG
XJpgIJBzO40XPpo7VFXD/X6NkadQFqDTn2i4IUue3jblDw5okbvUnoEISEeH
e/qjzFMlMvB5e5OgOGOB/N5H+TQOLJU18GByjM+YjC9fY/tl3ix/X//SqrAq
850cw9KN7Im4b1+Mh3ntIiqKrjLgzY/dh5L10OiZYVsfGjUnE96IAva2Lngi
jiGMZiHsEQxZrkDeWkqdNspy0Y4ZfKVOVOaDcWGCnjQ08ohU2TWXw9aN5XqZ
JcVCaRDE5J+vrIS3iWabQf4QAL8yHrACwAOSD53pql0Ckfa5iC1KtVSo7b5R
XsbmP40Mt+rh4dbzw8hP8WFetUVIcjIwp/dVAbcHjoedtcRQZzeGIbmAT/PP
xH9VVXPoGnvWViAKb5dsYJkYBe5hrxKOLQon+9SvhhNvxxgTjTxarp4RYqkp
4TezNZafuq7SF7qTO+wwg+0rIMOX7nMDkrDObNIQ4HfGQ9xG+nzd+kVUXjOp
J/syef2s5fk9W/U2HLoTfhCFAr+gvjxUWNd4zr0xwhbXtkn0q9A+ixzNl/RD
raZcZ5ixF39KixtozuCRU9xW6HGjYCWwqBhyT7kDv8eSRBuhAiamt55oKAQN
3mjqci+BNMywpaVrPaCbY1Vw7KesMTrL1NRNENKxuVteXyUayKgKoHe7V8gw
KBZo3mZWsfCJObHPUNmUXkYTfYbufmkZ2D5CfapGDMoQHR43Yh4LTJKX6GRY
slS8Nk2kdNLEKe0OUF4HJamOCU3+xqy+nKPGiq8mh7ASHCIDpNjVN/V6EWjo
q91XoafgBhoas8rTXltByyG5PWIK46YRnSnE3jlBG14LDyjziOrKUcUa1UHo
XWRhCoZaMoEyJCU6gK0ZSLi0i+rP45BworT0jAA3227fNleznoUuiD/4N8qT
OPUiZ5bOCrcId6BWxa1dS9u0ykjYNQOzqSfVVk6jD0iK5FNCuA7+uj1jxJyN
tSKTl56tal42a/OTQvHCv47hyvVMrL2eeebQp4aCh5AoPuM00g9oJWkH1puY
7s/CdC3s2P8KpJ94nmld0O8hNMOwZIhtPM+LAVQU8vXzMI6JCEsMfHWg+dIq
y9HRjc4XnwnsqZB2VTwDudo5KElXs1XISUzxdXzyotrO7XcWy02cC6Du0Lz+
Hs5x3/gcxvfaNcpu+etK+5vuXOZsBSqwDjjyqnzU7QfU6l+O73BCJDlB5j9Q
I8pTtETvOKbSzLwxwfYcfulcLk5uijN+NW5jLvdATwGc72UVXSGUfp3rvOJl
K5hYkfzg0BPxQxZy7DYgi8v8oiXBQnRrSBrwNYO7E3q2+LNE7AAAbZtTOYJU
SkAG3xxqISNM3h3Ipyt01HSyefjSC2QxT5E9nOOp1IO/xzrLbkKax3pW3MW7
PPDIaImXLBudlSroiWbX9uN/OvEwKl5K8TmLFw1HCPKvs4GYUrIglvuCLsM3
QhXGXVI51sgI33WNThJMmbXvVlIVXJOF+i+NfU0pCXSL04q+c8mbDyPwdYHv
AkSAC/++kH2MNVnm2tt3a07hfoVJtJY4+xi2LsMnPcZg6WkupYvSR4IzaUhB
GAo32lpgo8RWxM0uWRq6QXSib6uuJ4nJAZ5ueBG8V8cz255UEBX3w3UNC4Ct
Ja9HKssedAWySBjsVf8PurPjc9oqbSDBBfw7TdKwfjaA3VS3jaLfCV5mhDXc
CVtzmObjNfhwnFM9k04uayIsiN4qHkhkrExPc6MKId6BAcRhNCzS+qFyfSQh
T/MTxYbdZRGQa4jyyXD5S8RKKFzUyeoWPH3tFmKcqJS30a4G6avcFz/0iIcL
JDgawnU0U6mty5qilLbkN6DXvae95YfvqFCxBmgWpxwaxNy2m6Fjta5guG4t
Va99sGK1/IAiZ/3LlHWe1j4jFJ5uXIqjofFy1/q8NwQIGV1SbME0go1QcNc4
/NAPylPJVaAmO1HzzUE5xkKt0q9uF9paOoNVrFTeucrd+x4eaULxiyI5gQli
fw0hUAPIaNZlkHwtGcSr6vnTlY6ieY1iUDwm+khXE/YFTXbPkc+ZgWc4ELub
PGqaHoDxpcNoozmKFZYXXDLCXsAUJWUk74uzyv/5xEzpRDAykPwrqCbLPea6
Qam8juR3AHzDc/DlfDnN7JjMl3FjEbdTn+0KfN3xc2/JmI+HioSjR6yh1nec
NS9nArbKOi83jEoFYZDPZTIamEisx8qlFncEBv6KefqjHU7LUkRLkmNyUjHj
KGPgDsUsY/qRJTHg9hxQrT2on5jFnAi81yXxIUV3EzR+exZMcWbU48atzAA3
F75ToEPX57/BC17vyrdjEcn9rOTVT6jf6QZukwR/4ZNU6vkd+29NpK7sBMhi
8xpEdix6BkMcxS96+96YCflIaAzsPCGXSkRdInQCx6fQ2oIJBtR7TIyG7abC
R7iMm1008G2qcHV1X2rP6bOLzyeW7b5vs+JmZRebaW/UEee/vPJaVg6ohgxs
Mgy3VVJbIRRkXwtSwkmvA7BMWpXKxsLluCdGrRDj1pw2mEhyhZrmKAsNUR1t
Ci6QGsPhdr3M5X2zBBmmEbZNeXG5herNZeNZpFkQbHQ2miOHe7FbA1dy1v55
eJvgWTwZWmCCGsnf3EbU7B2jcQau35SlCtKJSZhmQQk/Iegrm8IDfKoq+E9m
OzKDfQms2n7NtSlsmEAwqJXO8CZRGZ2zlqPRz/GT88wX4ykmYw+fyo3VCtkO
hXi5TyIuwUdFbItzsYHumFC8Ia/HRVhGD3dfy4+vnltdarXa9CUCGCVAlFtq
irO2zKf/l/otT4k6D2jLzvSIc54KTHL96+WeEk/V16i3tQIjt9V52WvfLXK/
sd6AyTwBTdCThrCFFx5S9M55+QOFvaQoz8UMrWGf4KgUHf5asEdUs4LxmlsX
95aCGWkyp7RTZFoflPbgO92EY5ZpBF78zwOjB3PHnHlAXOKoD2Kq1yLraeW9
EWLc67ubX9kphPox2DK82UP6m2f62zt6BruIn9chWNwN5o9694fWv1hkFgzb
PBYwa5oB7Mg7sCFBVgtcdvH0CyxmeBEjXyalMR/D77z8bPot9iT+7w2AuqFq
f45QH4DT9vung88A/ELFyyylDU0jB/5pzzaCyHG+I/4cBDY5wjVC2sdwYHxI
BPXneO91TwQroZ2jCIm6FZi4MlH7C7K94nU5XuoD0epB8r9VkjsEog6LNeCa
rwnA2ZQZ8Pq9uEwBEJiruefTc3FB8kxXGJrdw1LgPHTmK7Q5UuwX4W/BBy1m
SNaMUK7W44ljjXk2XAG9ZDzLCGahQkH/sZi+oCNsmn/WQBhBOJGxKsDFBdhf
bZuDx0yecHJmAlGaV40GsOkW08ufa5px5J8IgDEVFnL/1FUFhO5YSmDVq5rw
PAKloraFTUT8e0WrlQzjGLob1sYnCOOlizB9zF1+gOFl4jf8b6ZE+XnUP+hX
QJkOBhwuvjnDTUj7mhZYIMSuEu+hE/QlMOqhdZKStOgIdRxmV2qz1NtO7/eR
X4r4KzcqaxQNyXaCnvGFYvtLti3IUQ1Bi1hsJBr9x+UKtYY25LO95kKmCXIz
aGTyXXq8xBCc+K1teDgpKBpUFjaTYB/rLyeUIx0GMHHWdQwSYrzaaMU5C7P/
wGXdLotdcx1Eil3nGeVvWoRLXKl6g235XlI4K9aCuHH2/OhICEcaqpLoS6qM
G8w2G0CfRuBOyOzFNXiv7mZdDWxCQpztNEQaP2qt1rPMcyhXc2QFAZQr4kv2
ujr6/56LMvWo4S3SQS8XEv8hasBaP5E68aDTEP0ZH7AzGN65o3R/79dQpQmb
DW/+EDkJZ07TZgcLUlVAFd3pvGof7sppcm+tr5wLVGU3yLJZ9zLLj1lx2ZWb
hZB1REaL+O+XrkY2hiOa/DqE6wujZV8a008o7KGAm2O+nfJHXzw/iIJ9iQR6
QI7PDQrjCXiTeCQWey0eKkL4uD0xi3KBLpGGsbkNN1U8An28o6SWG2Tigcq/
+Bu9AGkQbeB1/mhiCO/pVKyax1hF1yMXK3buSRJkn/YE1x1I7smJ58xsq5+O
CgSXW78Jrh8BXeBkqORgfgvJAwDswHww+Y34O4xN7nLW2C0webfihFj8jF/A
UqXTg0kPDXBV6FrTr2FmJt2JKpal8v3JPwRFZITq7SYim+E28p0QjxY6wC/Y
8vFzogJ6fOfFPjbwmmO5azzxjMiBZyRlp39Qbv+Sp8MLvmKRqHk22SUYNTt+
TAvrNEMpKH1jV7fwC2PVrV4fSpKgaWjsfu7a3ULv4z57SHo7LE5PSzsIPXme
pc98TFWC6a8wUkrTY+GSRrI7szPII5ZwMHCSywLChiSN7OTqAJtmi0qkemH1
CUUlB7fWKevPVyOAyEVabO+h+77hzNxa142bxK2Lwe1FPm8H9Qi6Dw1N6ZLO
rTVSWSQ+mTaAQqlcy0DG54w09UL/90QKvby+c6jZNTUcHKt2A/LiyQnkVW6r
soiTj/rUZ8QQgoNcJh7HL9Pe8VMMv3Il0tftONMvGyG5xhd0/UafPO+3gJIQ
cE4rWfYO6cMFAmG6Y+SiERANiUgXRmzIz3zbN0SJSprYau8b8q/qI/pxSc4H
McnPXcj9+KOrEYM5SURkQi8cELg4pE5eYtMvHMcie5unCggUYVF3mdgqjzcD
jW6+N1Fk/snP1BrHYL+clH0uv2REBhbc5e1i+ZSwJpP2vUKzA16KpTNqx+eU
iNkYtWSQXUvwrT7PRx0t6zj6kEV5iDM9AF09omY1E0KtjPtJDRmzbtLgKndD
JdD/1ZWZRlcSVygVIyZZRiW5DPt9ONfI4ys6CtSFlY3/VWS/6plMKNK7nkP2
61DcIDauqyf6cSBw3UBHndB5WaLS1RZ7wDP/UR4Zftrh22WglllcBZ4LSj0d
kVm0Zqd3ifEPrPhxDDHCkqCpjbS4jRPr6epbPbm4aI6eKoAGuv3bjg5cfRFo
fJJU64b9/moqQ5/BHcbrPuYy+ZXdOpSp/OMyJoNPN6a43L4cG48xHXSPrzPn
VU42E7XmtUlmVbWxsmXoyreW92gFTtEHgOKLX1p3L3KhpAppkFW3AgsgnEag
0GahxHj7P0EGhP8Wri1KDWG2tS9XBuY8NCXSTgJkpFInS0jG99QqwPK3yMRX
LUgzkaJione5ujCXjV1HfD0Xhg1rYB9HzRNYLenZUNxJAxD9bJKX78cs9Tam
HaTFSPraSRpxupJDG8gMbLpO9xEMaMtC2kxGMgujtXEajKObSAZvMK201sr/
DaCDnH7wzqUsWuEaYO6GjHnkOiMQduB1fmboJeTgEpztfQPn3tR+WuvVVh9Q
JaErADxfhEkux84IZz9224azKA0gtH3qG6PoFAvlag9H0TfXbGJi32Ovnu+q
dI1KdD1vpII14/oX9pU2TKZwMqCtw6NXQ8C7lN/VQXZ4naQLd9oQRu0ej7mw
MdYyT0CwZy+21Rx+5SZjzY1KTxPk3LYFsyWQ4KMWmoTu+/Vhb3eblsQtOLsc
ELCQj3WQwzwS3MakMqIt/if0G1Pr19Z5z4sFs9uVqF242TyGK5aV69vectAx
J064BHyiiRQQlZB/PThlgBjjPerwKxX9Lma/ix7QabpBsCQbOYmCuOeUq3Xf
WY9uatC8D+xW31P87AzaqHja4J6nqvFMONFB54FWkOMcjgfC6xJgLodph7zZ
ilX8XcpUe0xeN/0VMJWV17gK4ZHkx4khg+bufA9xNdPVN4ffC/UqF5FSgOjU
6l8Z0O2rmlVgOb999M5Hox0b5LbGvrSAiX5BBMjLHQ5XMjp8S7bkVeGTH6Ei
962SLAFMuld6EcK5nU8OnCriR7dB6ow3nJXLk3katwnJCRVdqyaMR5swiq6Z
RaR7mRWwWDAK/rM7DIh2INJM5wsCLeud9eYHp7PDT5UhV2KI1uUQNc7uMkVV
ouYFmICpxzlDGBAbS+ijQ/mGrxrpppe6Cu+Bfb8vCNQALA3x2XBCUeHEDb9m
f+49BOLUvyaRz+7E7EIrS5PgEymOCMkHThIIL9qOlhBeeb854QgSe7CwD10j
SNjVz6LdUQgV3mJjuwSy74OTu7x5mL+XypbI1vsreeiNECWk9E4ZWUE98+CP
3sheFncileHtZVI3YX/OJ3Q7zOCrqkHkYNsqS4gH/xzl57UCzAovI7JIaZA7
yMa7TAkCwt1ZvaiJAps4a4ftSJm9D15yu/dXXwHD8pYa8pF2OyS9+3kne8jn
emFud9OOnTCgc+QuPqzJzoKIXwbHLFmx4ud+PYiCHhTI14A8JDlvgfgTZLrc
XrY+gQl4gCJCRZQeAlKn/G1bdNDdlRbA3xQGTyLOQw9pcCCZ29shvcPEDnng
sw4367KSxwDfyMGnPfQ2xBJ0HUwThdSMxLZ/43yavqkHlGgVHq1FqqxNf10W
YA01jRGJIfB95io+PoekCsFnFTbAieSdAjWgC5X/ZgdZwJdGDCuXikteHTDS
xxVP5GovC8NW5WbVS1z4/V13VBTL1LUkUxq5ZNxVF9swem2yjEaqhTjcFnk5
Bj8ZAqzd5VqAXVDqi7ot1GQHX8cT+AWhpvQi4/ueVFB3gT7CFRtzKlMTK12k
9+QcXfANPCW0Zuzh5OVZbTxWjFT8ZWLdp82h0PeCR3HA/mlnTDCCs0KpeEx0
ZeJQ6TtpuVo7rEMLsFdMheDXmGNWe9eP0tC/mx9GRXfQaOAkHXe/yk79xTbl
HSkgbMyGyuK1k7GM3V+WJz+YKKwd0ClXiLUAblMos5fygawrw+KGa+AgNi9o
I5DL4CEv0zHhbnWAge3T5HqGeGPkCOgushsXF60OzQ0Ipd+kcPj3gFLbBmob
gMxIRW5Gdsc61q4MTEP/Kc7vUmZCj5lAO8umLwwPJ8K7c6uMNRpaMXLyZO7q
rWE8Ga6c2x9P74MFIpE1QLOrBe601mvaBz5kNgVpomvzf7bD2WGNojXVkmHa
aqdj8KAfiPmAwa1RkUVk2ERzsCGfY4DyclGrw2HbsbaIxnwVr0FWDegNNQLr
0Grk7C0yUXNEUoppZ/J1Iw/5IVVr2h5NBX/9J4tv5phM6D6vgSG89q84XoJc
2zaeUz8PyyRD0i/l/Ms6n0jD5+HBGE/E0g1Sab5vTMS2qf6s5AYtEkazmHe7
+K8Vn4l6tQyLaOFU4PXIuQBwZ0hWVGR6RCd0w3i1oaFiZnJuV/TGOD/U4WFL
okfBauxW41JRaSUQDHGRvRGgdioQRAGZ20bPROXFioN/ueXydIG4Fp1OWxUM
hByHLyT0GWxO4AODiaC4/lFI0MPEzGHM4fwGuS96YuG8Pgb73qpMJGXK/9cZ
LzizdypIbsmLxiQINlFN49X6MVkwNiWeEclOsAnlJtp8U/+Bf+1wR+ZHAcB5
RlZhNmSFj+NMyExnidbiPFVLB2i5oKt6rH1hduLZ388YUhcrlnXbkGqLY4LZ
LTbItC4eg6T6k7ENO4vYGjFOcYRZHtU5+s3V5DMEXuOFJnuCyw9xcfcynhUO
xx/32Ibnsy1+E3kTwLre7uol9qizRcdO8yVhdp8KlHEOYTUEcg1xiAHtQqyG
5lGmLsxoP5Y/djq0QyZqhcCs843Tt/gLCk5txj6AKE9Ri7He0XWBoP8rlM/e
MFlip0joVEZg/K8z1KZo1nzzi1aP377N0EDxKFnk992f6s+odiNFoHMGtYq/
cSeVISHOdhQkBcfyl6QtsyNDJRuBSgybkUmc+OMHr2YSKYum+xzqNAZMpGRk
WFicb0v4+GEL01aXH0nBXsjnfmi5mc/2/jQAud4G1I7K6hFs7NoLtKwrtpur
ylIHOj1efRmwFxpRsQpLgBwzVzyRNi2FGImrXvJiKSeZyLwhtZhUi5uWMvA0
K5Yp4PNE7djf3n3mGzsZAS2Tsp9j3lGV24TOKS6PLysBwr+bMxoSKo2arZoH
ZI15ay3zaBpgTwR8DcJGK5ow7Cvq3w3GpaiABSRLzIIfwubFEiRW0FyAA8Xi
+2Z0QWMcLHytP6Xb7LzyXA4zBENRAqm8jDdnzjhdgS+ayfJCPrke1lMzISlK
etnXE10/9aLn2Ru6FfUpgZnBqzzAdW4oIWU3SpXJT/dakuLTChgqVUyr35tb
dsTt7iMv9x5fOa/NYfuhwXUZNW43ZtinFcgRfYBfFoXt52h6P35gWHwdDt25
5jeZpnphWqZbX7Xj6mRrG4OMCs3zOuGWJyS6MWm2+9Ne2WMncWO/B/xWr4AH
cmrcIcz7G50WiMKMgCERmGEROcGxZX5C874dSOsWdDjIoiLLar4X/AeIfeFf
44ijfmxn3yE5eWyC8yX5SGWbpnLJkVutff0XK9CDHNrxD4IjSt0TdM9KOleP
9Fvq1DOCdxt425KmQ++iei7plLvP9vGOa+0DfBi5A9oImkYr3AWb7rM6JiKq
AFCSZ+DEy1lcafXYhSwWY/wvduAg6Ua4iLmfatv/e8LRl3HhD45mOLlTxCR7
kvr3wqjTVSmA7G+2jQSF5P7YAi5S8H0+jzI9t/FGnjMPue+4NPzgPRfHgotJ
1FJkaULTWzrxgm2hZjOkM6zMqJVRMokxFVDPwliBNChduFokiRh3faIIxPBr
XptWKov+tr4+Eqs6ULNsFTxDamm13JuL7Fua7hNjqENN/kz8uAz/wJCljZq6
+0N2Trvc6aZkbUKSoIPuADIFMTO85TxbMRDcmyoH5MvjE4hBov5wstaorJYy
zbOYq8ExmKFcuLXzU402BnkBC+c8ZefnsN0zq6RdazSrBbrF3Rq2k8VJg4VU
a0h8o6Dn/295/Ydbwp0QSbIfX/UiTpkARe/HYRyUgd8Bs6sEtWsJiRsjqnnL
wPzw/kIPQnfkk9lG6nVr6t2kiCMy1VS5dwk0YUb8Gcfhkhl/9HtirZCZQqTL
YS5TuTPTZIuX8YnYOklIgWx4mPpYcNkpDpseX91yRS88oqYjLkkOfwhL8rSz
yZR+MJB4san9EdgYgcYumfzndYFaUBdGwpTGCVB/j3lycdQMInC8W4N1kFfQ
ehg27G03d5Ph6NzEy6JSVaQ5SHbRVqzKBz6ldJRABhlh/2rX3CwZT1xvRvcg
e04tMgCqkKWyZqN3dRo6mY3mqMlBEy8y5Yp6mQgSrFxlEXOGXm3vwHd2ZzI9
aCp/Xsh6+vp+qLnB6RGdQtEr0moTc67YDiNnHbaGNF3hiB5dnQjiYa3o4ubK
4428bJuuXpUKQAYNpbkknh6m1/Uill4AQQcI98IIAmdX7+Kwa2iaj0i2PRgG
AlFEXnybtDZdf/nH7jD9zwHaxlY/GZT0mbxxhKrDCNfOeXHI/9Qg9qTGCTo5
QLBeoEKr/EyE0UqjdJvjDozgG1bQFq2LcLi83loEKVKq3QBIN+MOOEL2emvB
YPEw8TwgZCBIeAoJMh9L6MKcSeVbcLr5ASd/ArO1Yir17lpvikXXH4GCdEwy
n/CuHgtNdqElQRE4AFQGciDwQX4WEERcW3hjLTIL8UkT2eNQ71QnA9OM9PzH
Yu4Ti5DocN9yuARIHxc3X9ajR0ezyI0SDOHo7yYAuIgkjAtNJzLCfzqvAy0Y
YCWio2G7YSi0O3uu95Y4IaHYnzwsv0iKHgVuEGtYDHa1RvlQrXy5sYKIC4CW
BOWRSsRt9rb3ZFvmjJNu2R2lF9Sn2WbpZgxwxaupq7xMZ6dIEcDvqXa+4pZe
TTlh76oqPKu3zX3qNX4+SqZjRru6nbG7EB5kpYpbOpUNQxdzTel8pydnvQgt
MvTXwJJuwZLhp5qoStAnTKalDZJrw/ZUM6raSWOvTl7l2NOt1MI+A7foWUj7
CSp/WVW/awYX+Mpjxm1/h07AVQ8IzQfCTOTeRiE1mDHK/J//4FYdczZbpSlE
GB6R+7dzfxOp4agssF3+4dItBz/otPSc2fL+FXZqeL50H/l6ZQVdgf5ai3R6
tdVOlro5uULHet6a9zk2qqsuHSHgDvQ6yCljNtNsB2rMFdgfSFA2z7j26WAo
uu9MVkxFqOEscN3jZ3oUKVS9v/NHgXJWf5hUrJVyJI3thJ1cP0r9LGGS15as
D7PDJm6WT+vScwy7MyZzFIWaAcpIW4wUfRFW04cUyGJlprgG/E6eYjjHUmiJ
LCovwZ8USlp1Eic+S/BaPIhdR1DssB6s9Ls32SDS3RUM9S2IyCCwUfZIul3A
SMqolBzO8RwJr8cuq7gfKGkOvFXtPRwbOBT6TTQ9vYTDEj0dJ9YS+tS9OcYY
LMj3BsKKrpWtKk3PWM4oCDSlMMcgMeHmZ8kFFKNxnLR6AvSyK0BHH2nSt7tx
6vQUJHuF+4Oc5+47xcvGtJE6rM2dF74uGCW/fMv2KXeM7NPkzMKHf5FzXbp+
NdsqP7G91bhgAi5F3hce1aRc2BpbzPxNylhJ5uKnnDEU+LX0EfSHnVlN1HvX
y0I1WZ3R4tB/iVdj6gspoN5lZZjHdAAALS3p+oM4Temo77gAIooTJy/8Gik3
LCNBc0i1LwzsE46vLBeZbeRnhQ2OskiLmTC6HzVqdUagFQ2YU505bprMK6st
6ud2dbPO2kRmYvLb3e/YwEXdIFgu7ZgjAjBY8eYo0yKlA111kCqpdy0JNzHz
NrIdUi37UBmdzvhPSQRUFg8JhS0GKyfNzDUEJEHzB+jt96jUezNxanMckizd
GuSEDmSr4+AtF5BySYWqQJnYt2VSK9pbIlBPWhrTBjmUr0a7cJkFKxkYY9qq
SHCRK2kb2ZdsdU17crRFwImPta1Gtb9V1DnLTFR7ZRrYk+7dTWjAJ7F2PpsG
iowSAOxAzFzCsUrjnxMG2nHlL52s+z/DkbWqtMrXp/1jK54aKwj9kMLVGh/Q
0ezVrjPnvvj8T3TXXWKaw7WEiin9ucxcT2UJVViLPHRGcpl9Dsmm9ug/4wVo
RQ0OwSQoVB4bb4OBHHH6lJy5eEa1fmo9eTC+wBZYbuP78J57wX6UMTH4hNEs
Cdhu5/St57vUv2XMPphGC4e9TEyK4omDb1IgPgpC2P9l9zKH4tgFE+Oryv2F
djhd6ybs+NsGvickUuFnEw0jHuJ45WjhcPf3wncAWPBA6gPwejGoVX908FlG
TeTubAOASfp2wdlOAgPWAJzJCQj+daBEjfHkbATC7dYC0gYPP4zKRNBBqhgd
NycXUKlLP54jL+zxZd627m+fX1e4URvltl8WZZKz35E2FF9zwmsCiu9HVS1m
Y1Fjj3lCo4QOFpkgQmwKOHKzs8yXWxA886E7wVKE3zU6msD5iXm3q1tRdhsq
38y1hybqNVjlEzupZuHAmjdr/HgSSoxxkOmvibwznavEJnNzxSCT4wfAUtdn
q7EyMIjlQ2cCMP0v5tn6CjbQlj5kXq5Y5Rgqy1fxBAS01jCAXYCIiWNueK+j
1pny6/rE441pG5+Zf84FN79YCPUPMSKwBRbz+2auP8gxfGvovvcRYTsm9P2e
MWDVF54StgoyiXTTLjFBi5pC89/zihVWMXUc3SnusHKZ0CUqgjTdWGCUtI3v
PjYuJDfkJeKs0e/m10nGDfCWRv035StxA7j3z0B/ynbYMr5KcN4gJXxzYJs3
2oupYQgsNO94NQt1F9pE1UhxCd0tWmZo3bqZ7xE+mV6ERrCQTt3qml4mkBbs
Q3vA/ta3mXoG7KP2ATpADKeUVZYhJUu0PRR9oq9OWrH9rLLFahZNnJdxPYJv
DfND1bnoYN613IPnOsDJlwnCmff9YPJTJnaHwPcc0emJrW+a4EbteyIW2uj7
Ej4l4M38J0wuSq5ECs2Ws5XGp3PE5XEyJIJj9aYF6SfdRxUqtRHja4LVw6U9
AnPUIjhCOGSiD4HCBQ5n0zmIEOCgfGCCILJ8qYqSfdtuXq87YFg7eCz67ufg
W42yUzShb+Y9iqAGpMwE7CLOx6AtcEb/VNNuPdJ5MNigqP+U99/F/ObPpidy
3cQ3xwdO33MYg0qlY4jpgaEDTpVSNOKnlmpX9kOHy8pVX5iBQTiAobfVLK2p
6He0lWebV/z1RQj74qD7qIKAgbdxBUqt+QTEByRtKECs48TCOrPuZdt2LI3l
utXk9HojmlV5wtvDZtayiv/b/3qUbz6UBduIo5ygV+FVEcDyuQVPIYcZmH8b
T6T6tv78CFDpKrJG2SuErVZx3XWzp0Mkg6OUmq7H27BRqj1hTrBYv38Y+6jV
TZ+aG351P+gIn/YE8ea90sUB+4Wz8JguekUh92bmbUJGWowYfSXL9kLc+On4
hrsr6ppXbb+DVbesrfann0Or80i6VyzzwRmSkd2rXt/reZgwyBACnIM+NlHK
kuoTCxAuezd5PCsf7BTClz5YoCmxqBO4CDp7MSKzANsjeijG2oXBjWOHu+0x
VJ+D2E2MtriFd3b8yNYzUlEqn86MvZDE+J0epxnCTRJDpbKM5SZliGvHdU8t
j2T8KxOAiRLNG5Dahn3AQSW2YfKVylpb80M8n64RuVzK5P/HzZD4hveT/6Gp
kj+BSdS2trdMxH76tVl/sdbIteWP3rK/Il9SQCPv1CMnNJO46fhPadEa7ZBu
qLDo2hsNTwdm5wDBTzG8fo9O/8hCuTLKasJamQVyKvPnOkO16ifTndzk5JYp
SHtVPv/AbgRzEaQTmScoByX+9J863G+HRGYJihuaoIw7ZsLbn8oewQ33jBfa
l5kNnoa1pVBvU55Makq2Rdc1PFDgN0QUA7mUfBCDSj/mx8FkzKkFbE0N3ffD
2ZK1NiTbXlznyOlpH3y1mJSyLYzFNk/4HjKH0fVb8VkTqLLzyo6r5LRMbPZo
O2v//z2G4Q88WU1JfATGZ4Wc6F5/tKAkV+IFz5TWcgsJnckneafVmZU+hV5f
8zDw/SRkDa9E3D/ACAM+Fr77xqciBrYa0SIoqlgBeHI2J4daeNlXhGfmJnec
WJOniWvICOfBw/XczC3+RYzK1SrChv9ARad1lngzLxlIeewg5aRkakI1t/09
FXp2f4cQa2lL1gossVEItw55zhI5ARDH4CMnd+cA0F1ZyXRsSzvcKyq+6nsa
yBENAVFK+/yIT1Y+98Clg3bjmU51a42rA6yJ4DE60M+0aRPAq+jM4Hjo1yK4
vbmMK1Omk3xD1ot4DsThdHXw96BFHEg+GapIRhzRtttdX4a8EX8B8ebNHFoE
ENSf37Ngw1kGGHuwWYFT+1xeG7ndB8ukevmP5OembnMUDbVLsuOcC3qYhHZo
q+R7nnnOkrfg1DrTA/BT214x6p9XwS1WhL1F2yM5JN6x6I+/sUjvrhU0c6nI
c7rTOfcNzIuoAjzuupgfwoXI8qMI4G744gqLuHrVjvwMPyf4KBm3jHZQM+L5
t6HDT+ZGk/1badG5bNoC3y5KFOV+jSCYkUZ8GoQABQceQj6F1NIuuRDaZgRP
SPb8v2+rNAapyAaZAofSb8i9ew/e2dCrn41J8ndE9WDdIBozvZIr5tNkxutK
Q62YkFSPIp15C3srjpfVZ9/tIAcelFP6+jLn1lEzfRrzqFi1yGjNKPVbFZhQ
wSigrZD42o2S5FVAaznexXd5OeR1Hxhkkk3zxE8mPrcrExREU0BRtSGLGQ6s
dSPHtMwBIpClu5GdbsYqRpQn8pEwWME+S3W3nyZJH/tX1x2tiVIMHO8xlWp7
5DGRHWzdcrq8oRyS1EsHvBf9dUZ9YSCy5TcSfZgdfMy36t3By8lbIEPmcsbs
cjBAU9HPDg7OdfQJdRLNoDcBBzMaA9lCRew4KI1kPNbMyjt7GWIeAOtHUioa
4jKs2TWAWrrA/DeZiNXoFW4d/HELinJGXmLclJMIqH7ogghUyBrnva09bkOX
tKTaDGvk8r6mU7OegW3U6BJch4mCNgLcuHp2oC6Vz216Or6wHJgw69qs+tv4
USbIziBHMj+qD2IsY68TRlSWwNfARIJ6IjGp11LBzVr9mMOxUmCd7I6LE3Yp
jbWEHgUa4/02v/Rz+e/ng8DRQEQ0KMJCYE8vP5gWG1Y2+rUQnPG9tY8YaxtV
ndOdexVZL28oYl3rhwa3zngqBQIaeS9frHEs+s66UJZCS6J7jbW0MgICHVe/
VzWh5TzZ0Hu8b6GQ7zA4+jAHKnPJaZKMTIWiyrD50yf9GIM2rgKDvCDAXKO6
lXCinM1kNFzTRgOkuOiM3vCJUxy28AHknK1vzRARduZVnvze85YckyxcG8gQ
ijqV3HVZJHoPTf8I3V15oCADilIuZLIgHzwzQG5QjrSfQkFdCY+b1jTKoTHY
6RLKHy95JpAoQM8MLkNWYkU2vXn3nn9Ca7vS1VIDYYk9bemzO2LumTV3LnC7
3aze14RPZPjYJ2X/P+CybdOUaiUeCpZGuMEZUd0+NOoD3KKMOsLxmDFIb7jl
uE6eidEmhNypGuN75zTrUJx3EQrMGwZL65Qkh0hDekiW95ImQog1o2RuyUXE
L6oWKUSZgMXL24c5Yjgpa7UlaeOrhuWOKi2Kll4c8zHHsqd9ICIXyLaMoTaw
jTzCMpIvfNtrHxTZmPP958vSvj3JUbgVjMWUEawoq6p2TN6bc9TQm3GJWHT4
i7NhMrKYgbfNOQdp1Cl9VSgxOgHSWIJaTeCQQUIsjzMPhweqAUWN2VsK6YgQ
4jCgLEYDq1ezz8UQUThLKot5Sow3SPlni9fhLVo9mZ644gy734j/Sq3Z/BCi
IHjeCn1Z0EBbgOPqe2tdYfm6bSgTClp6/8EMLTVwHWsDbeZLPnbv/4mU2Nlu
hF5YDncpb7WHJ/7owNNWInYeKoYYZxdsjkFGScQAAw3e8FylErYBQvibbASW
zDYBh9p0ugZ1NWnd9P7JQeEyrT561UXnwUjXY/FHyLxssj6x7x1u7hOru+0U
LQgq5h4hRdCEaqUvsLd7y7hbvN37w6CwezjDzT3sgCMriAKXKh6W5u4Abn0W
W+SkzBAwz6Fo290+V7D686uFDv27Rw9+wjpeVIDB8fvjUxvEXoFOOH1u2zcy
dqjezyQBAqC4GhWxC96jvDmbgSC19be3/skceTGLtYN6/RSzAGxbG9NnsnD/
dPLOp40cX6m4ayq8dNq5nD1nf6KvrJicIG65aQHvAH8d8f0DRow+2qXs+FJZ
sarROUq3K6yNgmsJsWcjUPVh+xZj04mIJHEQ9zCeIF78DAMmevffyu3HSFu9
jHZ0zmrgpmhrWADnLHLkCJlz/0mL8Xp23bh3vSrqYfjU5NbZI/7hVlpXuiBs
8JODNj8KQY0ysC7PY3DwHTN7nMD7NDyXQyHkZBK31yUJr2us2kjYzio4/DLd
4vpban+FixHfcL79neg4clrOIDtFQ1Fq46c/24KeAx/ibEUP6Bvm9/DH1vIl
eazAxNs68xsCrbUzPLzQZ5XrBO/ZF7PI1q8YWqWjnPJkf+6ipMUM4zepgG5O
nNRBt37KU2mk5eu/P7vsJ1N1uVznEG8o10gG/lo9vxSmq43kUZK4jUbEU0is
+r1B6nCualWGgh8YEcBZJMKZ8P8+DcOfZlvhOzpSzWWRBPOX0RN3jrgnxN1J
f971D9Y9jfgb5CIeLHnSZrbGBVi1zM+DEoXTk4ju9yPSzcEOxz4h7kJ8IWxR
AN3e7TH/38i+WmEW2NvMviVSX5+WKkmHZ56sY+ZHN/iV8v+VUDr3U92aPmLf
telD/gMlajkdE30Cahz5RoojjHI806J9KiHxqSYIHcoE3Uds9WtTA2fvam61
HtGEJ5u+JnUcJhMxroTWvFHGuthlIAI8LdV7XiX3T9eohvQTEV18qDSgJnqG
tXeobkJC3DqHJMszg+PgOVy5ulZdryV1U2iYH+Msx9yFDhWouIQhNfsA8QzN
xcGESlZ91q/y8KtX3TygySJhzog6yQfCKIEUCPEZ0S/CzPwlt/fTby+q0uUT
qSRnD6balgUnfbeyfFSRtUU96cgnZwq3G5OG5BIprD7RA/CO9zP8f/0Sz/g0
Lw00KPrxhKhYaE/2eZxhk5PgUyCA7+a3vxWqi+rL9DPM7//9H2Q4Qcg/23/7
Fwkry70n0Lu0J5eyU+z1aZPmo979Yb4iRVtPlBivS45cKwmGOlFBqNrwWpIj
X9Ue9Qe9awwd4vcaJmBiZlYTDLTvhe0rtlqwXrsELLeOPUg+z8Qxxv90gzRA
AljWDk1jk8YN5xqHtK7KffC0dZjmb16MoaICmpowtv+U/Ro9hbPGKnM7ElwW
2nzwwmGrpWTkSz+fnfb/AIo6zA+A/u/Y1Q0N6+W5IQ/ls1JQDlrwADxycj6j
7QC6ioaJ4gWXNeJ8bxbg5hyFQZfgwKka1I3OHZnw5cRV7TmbILsk/g1T+Aaf
S+KZpXOpABe9IZDqNtqPmTTBcsPwO5JumV0jQ9CkzjrNWFOIUWFBQdUbax6v
bvNmAAzgf3bXoXWmfLAJ64WEVecxnriTQqhi1PVMU9YTmvYV9bcC6jHLTaH+
ebZl5R5kuz3NiwOoG5N7yEnEet+JMAbAi47mKo1Urly4L33WVbV1642qa3ga
yZT6RNfsTYB8F/7Kz2asTBvdcKZXmi6+ba4LIN1smiQ2uRK/dep74RQkkGkd
9Fu8LWmea1lNc7lcQm/ehJR2MtxFy7jBVUzTger6S9F7UY9RQCGXxqyObXqS
gtWkvKHK0/GqxaOmLEleKZyswG6uzW8DEI3uefKNtv5R7Sf9RhrQCEMNwXBS
anqpRgSU/kdu75cFMJWMNMf7U826mp4lJuaoELB5va6yvldLUfuNf1NuDvEd
/nHKRATf+Lo0EwftsFdt0NlL9DdFrS4lZeLJJphzFB8csKZIpiL02faHGJqZ
rjbiOmnEDu8wTo1dVtYgkRh7haS609VPOZqnzVb9tlck8J75kOuNrX0yaoZS
V9kK1w3dKiS+4G/K1JzduEK0lXNKJtgBVL1W7fHjIoi2DzEnuOPg0ZYH46tv
K0Dou79eXSwsz/E3BNqJJeFTRvhJ5eFu8/tx085ogE656uLdXx0bNg9sNTmU
lXwlAxxkSsWoeVPnaJpiKZFPuI/ZoqPxlBhxoutUNI84oY4bA0WcAdvuEVi+
4rf11ZVWJhZNk2+Ne23Xswjk39/2MATKEM3F+JMhQxv0rwlXdiXF87TBwHiJ
0efblPiKzEfiI78+o5w4SmLguogApoAMWKmy/R54DJkcz++1j5s0m2By5NxO
5rPeOCAvU6jESbMjp1GqWzTVHHxuWCqqQHxhm/xOD5VpfJSui2IdCZmYUVYw
7GWav16ZQPqD+XoFpbXL9+x38b6C8gB2VzTXFNNO6Nb8jbkvXpbpDjixMCW/
yIU5YM+KUV5bQ+P2Aq/isHRGYGpfBwwuiyHNi6hZyTlLLv0kqm0NVOgVFr1Z
MJiR8fEpXBCkmmloVeinkAQn2BPiQVMC4K/L8DLx93WC+fwazZ2acdHbnfDC
HXYlRAcXreV9tr2lEHLfAIXCySr4ic1c3TQhE+Mx/FQzw03uADEGyME6jqOs
ll5AwsUFIsWYoQS4HZ+tXW0tJz1Asw9+Ck3Lw4MEzylM2MraSNfDuoaMXLhC
m+GXfZ7MTXSC1tAo/WZtuBWOKWBhjIePh3F9+g+YEDyyGK/8/FxUB+cDgwEr
a9OVfi3kjvB1XAtAWizS+//8i0KsjkR/YziG62XT3cgwAAAXcC2JFYqKQKbh
/UDdiXgTn6SLyTYeFzFKpcYB8/Ryo5IA7MN2sAKeboczMkZEw+P3HdEKf/Cb
5gtEb+rkqE0z5HaDmsBXaziJEFKY5od5dspuegZl89InzGfPmPRPIrEmdEyb
9iITmw6Rz1u91hrsNrU/9aDs5oW4Zdd6+OETnKXbGu9rPYo1sWjbpAiSpr86
3spaJLfOWGooVP2zSKEJsg/VZL7gn4pKdSrkv4urf0bc4NynNn1NUyWAzQ25
qGjMf9UUpIyYhX53zD1ueFJ9a/mz5WmCE75zHlPLwxcfVr5l39OX7Rqa2QG9
/vgGWlUUjrgBItpRGDXR/aVJkCV12zrkVtqz9W8Qe2wheQdCvV/UfZNH9Xa4
5+dtG/97h5OmGAe9iaDSukNCpXlP2dlWT40YPLYATyB+hDRLxEa2ZLFJIGCM
VjvUJwckWyJjh+0hdzcv7N3EWWllqAQabtEPc9xigbJsYZP+HDHySPFETCPC
h3so1BjpGoniY9qF8ocnk3xE6d/YGiDYEtp8ALaVE1lWCSnenC147j2ATcNl
DMaPH1MQKIJlrz0y/e8wauiNKdRgj1zvK6qDfH2Gc0GM1yxB6hPycHK4vOmW
xqsbEevwfowJocQxzCLbDKI7Wfssup8iI7qVm4fYon+JA+AnkDSyu6PaAuqA
SFSmUYBGrZwIvB8Qx1t7vdnxtEnTNxc1qWTkmF2m5zFJV7H/dTCxD1h85V4r
d/cSTuTMS+bfDfV/wHy0NZwQX27nFBScDZI8p2HXozR1i/evdkebY23WPOYQ
IlSm3kP0kzQUpdi/FKrQOyA09CFV7ogU4WCGEMGD+FPvZqS3vWcX0rNcmcAt
qopHrG/zu+3d3XN/VVr6cfku4Uc42NDrrAY+B6gLZBbAc+jTX0KjDeyIKW3I
ByaQHvhM9Wu6HKo+lEwpjyKnngAhgUYqLzz9NZoNyYF7N4g82Yxl9OyLkI6S
RvD0TbfA8JnqUwJgjVI4WBIaM9RX/uHtDz0cVhyb+U/S2lCU6sZAbIcizoCp
tk8FcaWLo8DSBHAt9nl/nrbYD0xWH9+mqeiqgfp8YkNzYKheZTr1dEkRjrFz
noZjC6Ty2OTQgzuUnMm6k5unmFQrrPG8KogeKyCbQgRJ7LJe80JI0ufhhk5n
BFTgvR9viNh30VYt1BDr4rHlUQi+WDJbXG7ytMdtYqQW/pw9jVG7nYgDo+ew
FGK9dxcf9SSqptc4daTVGNZlQymSXpvvXNmrkmudrDn/N84RaxKH9B/W+256
QRpLo0WLFTR/Nqc0jERlf89s6JkndDanIVTzQHK0NbxNS8R4An4tjW8cCI10
KDTWY04q2hVAFB4M7i2iWTb1Re75KvtZeppl00T0RQfzoccXXpFoFdaoUduH
o1oaj3IEOoVGMwgumsNfC7RUB3XB/BwlSrz9rK4vJRE1kh8MFdjW46u49hVx
bJIWliZPyRZZWClVSDKV1ohRGkNsgdBQnE7p4+/XQz3Ha1XSIQEzq+HObGUZ
5iryxhH2tzv51o7hh7lu0cq4hsWFYE6LZEXY7Fa4mbzw1aZuKk4gJ/y/Gg9C
U4U5Ognf9mwMuCIs5w9qcP03Q3G4Lm5dj62efHUHxBfwAD5pEMXerqG4D1/e
bCe1O4NqGQsFa5/c4P4/c4ypIxu1/qlCiNOHzc4wtqNihiDM4nTyh1VPglS/
dRJ+aL3/6q0WoqJV+LQ9mYG6WaquIumRw25LVdoxcjfxWU9kw005Ojh/B+/3
foRutRUimLHG9k4Cj5/3uWit2v+cc5ZPcBW8USDVksrLhpe8Bw+md7WYJBOB
JkVmSbg9c8atlYr7rLDzsdnWy0Zeo/f+wZdgfrCMOFf7QKNdJ4FEI/eelqGT
6cN717DeB5jvhoTA9gO08W7R0lQa7z0x/YcbDcp2ZIuVqZ++GFQ0nv4M36hC
+2o3V9i6e3tUvWJ4t28/v5nmnVCoIz6UJJm9jKrZxGoMruYL++fd2Unj72bW
k+4KnKacTwV229QVDabZExf/M3aWhGp2KG/xS6M/oEprsbEWUOodkzZFb+OV
1G+xO27o7vGxOvlbhxhtCPc6EmK23GzJORICV7B9P3YR+IJZjbAc/z8o6e1y
hD40AUa0+jN8QUInEyRZiKu68nNrcJ6rMbLMvnGFWTW+UM2b6WmM5tpCodRW
YMZh1C8koG6B8+tdrFVwyoI6zdecbUdxf6Nw4eiBHl8ZMrPoORzV+fJtdPnR
ggUoe+0IZvuapphHufcMgHiN8K1BKY4S7SwLqvLz8s4j2UuvijGBcYdHsMVB
2xwFnPOs72SzxMmX+jjFxaItHJg9/FOx78siDRtqYjs4uujsNga07lQ7sHTe
b8oAlmUewE5T/++gpm92Xls1q86xA1m2Mcz51bhUsO6ds5Qrl7Lmp5kaAYuR
L/hTCrgZB8cmVRVKJh/6YEGg6qGvlTWvCcbtQ5h5+sCtlTbng9IRXypHIXXD
oBO6hIBh6fkdchJPTqMpQy7HfI+F/fC/Uc5NLm7oXgD5Ny6PvNhW9N3da6Wp
tJtAsHrI8ZfI5U7SGYilFBTUWZcN0n47tPezDu5GRoY6uomdSfACqsiipS3L
zj3FZECapFGYySLb8rQMT8cG1p8OYIWxB0+G4ufv3kK6ifylPtpCYsyPOgf/
MncQVdv8DGK9Kl/G0beq1LcGblJA9fXR9Y1rIaVi8aYwes9wvFnPmv+kzLtG
iwHMa03YQUexC7HvfrEo6ziAAJPOmSaMR3OIqYWI2PnjkJFiZ3fr+ho3I0vv
pLp5dBL+Y+vIdpx9Xgcef4L2/0D5DgIjLoGoymHR4SRF3mP9D4Fcu5eSL2k5
c6OJl/zK6u+SP3WBCrMaoKVc5AXNn0I5lish/pggv5pWrj+/y5SXR09atL3s
BNdNuNUcxAvdhXW/hA5G4pfPZcwuXIoWc70UvvMZteQDF1t1ZZEMUnDnEzdF
24y0RZdk44+1e3olJ5XSq/a7lhioU18/tY4Aexjn/DqkGAfuypD26qoTubei
vgyI8povI3YVNT52tHVQdyqgnMViK8IHqaz+ab1PH5Ac9VGSKj8kqz0R/uVd
sORxad+beo1nrePi9NMM2JUzYRZFZiTAe+3Z+gZ8wPiSqV/BrTwHIe59Hdpi
BoXtUAAwEGNDQGHsnvBo76EQJa7viAjygw87n0JddBwiNJntmSN0Ll4AbU2x
5zpA7SWSYjTj6mTqocGTELJUjvhXE+aijuKw90WBK2pgl5U9LUz4+EA96RMr
G8xUIm/HmiDl0+zwHwMA4zLT2narKUOsILqoQjQ7+3z8gPxPRdaLTZPQUOqR
zXIpm6qymSfgH0Esg8nc1f/lvYKdOeOhGJ59Jt4fsOrJtyk4UHHXAMvKpZ7z
VK6koY8GaksAGWoNpqgDl8Vm4kRbBSaLFO7fZFIY+DvUyP2jA6MNuFNpQl4r
Kqn48UKPqO+8YvZfoJmwF1eRcspYwspi8O0AoGm9dGigeZOZLf3o4FxqqmrZ
FQWZ51HiDibidLuMEOE7/G/rkvOgiozWcRMCV0YlAxCwTkYlUHT4TyEbrabO
WvdoZ9T1ofY3Iph62JFbQ2urTLxh6c+USuicfb+rr0bKw0nKj/Corwz5GspY
9sl7H4VO1UGZBFPmuLQ2m7j6PiT0BDU2gmBC0/Y6hPFcGiW+FIxxfgDTGoEr
LygMSs3DZo+xfksjz+9aHSoSHPB8JYrdrXGffjISPYDgNqp0xs+2pJ21eZbU
hof4NCkkHmLe5CXN9X51lvlHdRM+507QABzVpYZlZiC5wK/4RGIOeCz4Lhev
MlI9BYGFdXgN4nYk3zJbKKKLoHYZAu0UuriSBthUP1/H0BGWnTEE4cpcelQ1
6JcWFvFVGE2dLdRyntdLJMu0bNHBfmF8G/l+IemTbw8eUSkesl/tqmSQjawy
ksNfy7zwoyzaYJozkY2je3XLa5q8Pek1CZ31t4EELcbc/iG+C7Lb4TfZGfdo
fpj5PM/mXOkgqpfncTtincZSy9dhSjANEnlMrDIdmE5E61qOVchtwC/4SHsb
GtI13wd6l/vicoCymfyVXvG/rIBgTbJBA8TaPpaGLeCNjcBQiq9EiCOwaWNt
g6qk7PGV9mXmYAaBpJxyP7auWkz01JEBAnxjJL8q3ZEOv6qcimQFZbsWnEue
Yj6DXSkpKpzPsxlSIrVUf+N/x2mrhuzngRLpolDvrA10+XBKOfeiqgbogLZb
h7HX0l4kiusJDItUIcWVW6wL1gpV/hjQqd9wt1LyWhnowIJfCxyIJmgQjzy6
uerO5JKDmGypzK0zCjPaynTT2lWMmWjbnJjm+ibEqjvsDm2JoZrPVcqCFuYG
b5OT7gRT5WQCFxjKHKneciwwx9nW33CFPZmLN00l6bUfcG3qcp3pki3nq72e
nyqA841K/yVHDPum6FtzPNJ8gnG+YBZagIikbGuzmnDfM+3Hlnzeoy5fFLdM
vw2TY14y7D8A5ZUVcez1T1ycWzr+5eWGESDUu2Den8YG/GqP12Z57kQWaGFm
tcn8LEkn5L8TBBvIr0F5XCsSLhf1p3Tn3/LOVzpT9C351XxjQ6P81tJyzwp+
YT+alcu62ezBcKg1RUi5JLN/BSZw9dXw24BeB294AwNJHugUb6wSOdHnOXat
vPUzNn3Gt9cVgmog3scv1xRGdF1+EuN29CXL8zl1y5SFWAfGBoC/dXHg9eTs
OqyeezNZ1gn1nbZ0m6xlvR8YPIiWfRSWGXlAGkZdbWE6CK4wgYW+ybd6LIaZ
KW0EiywV36NQgsIzydfN6EIgCJuHuAGrdh5/HXDx3tZr6ytW5X8LstHLf3Ii
l8aCJJ8S4fSTs5lc6STYi6ak4VJVvmDjc/WB+ZVWfgstCGiCs4IlN7EgFhB4
BtinxKWyROUUqZnuslmOgplEVrNDZ0Ms/pJowr5KFIuAhH7QJnYJb8gd8986
aq6jasmFJCVPbPAGgm5/iaYPnII91DpF7B7sTEYvOjTX9NzSkVt+Z8nmk43s
g0yv8RwMEzfqHMneQ2kCM8jxvug1xI5zRK0YTwGmRj9JqAuQgiZCzQfhzefg
Q5kNu+jeRFwviZYWWKT6AmGqleEcG1RjORPeJCx0Phv1gIQib/CFiumqYiTg
mvnxY1fkreuiSX2RVCMBAj+KRXL0/hGni+Z67da3Sb32AAiWHR9XJb+JhH2s
E+4v5vos1FAkki78wtYQOA4MFF8DfS6lIG2lLPpvZnWP395bdnYkQtdyBA5V
M7afzjiyyK2QhSOf8j1zdfeQmDJw6I9VrRWmvSAdG2Eo9r6M2wonTqAjpmyA
73QuZ+vMYoiVDYIZMvt2B3MZ+2q8flIPSsksXPnxRjfaqIoOvtz3QM75MZcv
MVqePKh0CPYSgsvqCLJJjkpWUMCSSvtYg3JjBOJWdDQTcsbRNpz0XcbciTg3
hDZcWQZrX6BlbMwFNFwSik6r6Io0sLGvwABl3UHx68rOAY9kgKMS8OQVbDlL
C3t+HCBrOjDjkWUnjziRp0Ffu8SfiXvGIJ15v36pBRl3c+pHiSdXW/IWlHgQ
2g2krJYq14qL7kCoP4Nwt/ICXNL8dInJyJg8m0JFmz3wnbL1/RoYWYqxS3if
2p1Eq6jEeFFjSpCt6j5CWhiglYxhDohsr4wCK6u8wtwneUcg5HHt5TrMhGXT
6qOCIK8N0T1LN9zeKJFlw57Sss0leS2cxW0MCgfT08HGy/pOaji+T3u705Jm
pg59dEl773oRWfInI8r2AGYGdJ1rChCUW24W9TXfzJnTZvP/LHKvA5xbGjgg
CarOgx2yTRJrZxKNrIrJy4oSJZCH7V2twmkSdnGg2sm120P8Jzf5L7DSxcIW
kgCdopf+CP4ZR9/CMhg+tJpHRlMwXW7pjtx5aGK4zyGCIn0uecS6IYzCumJc
ceDDEwrzaR8BZk9x1qtGxBML8EoYbUKSxjU+qrBLUbN3jCSxYFw1qJ9Ox2uW
/D0Y8LsPQw7yDNhoqicGPJi2il7w0d8fNDduE3h/l5oH9RK8JE4A/7O5jWIE
d+vF1BV7CsSMt37zCFXMGwtD299NnzaH+wDrp88VysfmhqEFbAv/mFMWXqDJ
ISItfsOaCH4feYHF8RIuYim/KgwXejIbek3ZWlW2CAvupwnRh+03H9yO8hvr
sCbZLlqo97ysB0JGOUZlIQSJW+1B4p1TSAis5Q7jIQHPEgIP0fWSFryqiBpK
yoAMFHIB338LrhqUK3mkPdzQzY6fJ0/z0E9eA6JeHYhdZ+W5rhq/n6IQMHPs
WfnraKDyf0sH2XKKtv65VF9C8RXNUr4Dgh9Tq1Mdkum4eJG2rw3To4BjcMqi
d00uzqGlvPw9w5rYWz1lsVhZEIdLYIITOCWWD93H7FLn1Q+miO44twzSp8qy
Tagf6pBRc9XncXOXGASgvxkaSQU1t3Rje271gWNW/m3ABmP7IWq34Fut8//8
5+C7rhL9BK9/m6iGGE8i1UCDb7Svup7ABC308J2zE0ziazk/hgh5hqlke/hB
rREv198XuGK/7kvXt77RBe64qLmw6Q1tXGsdficux5m2f5e3zoVcpQxU+9vG
apMk5u4OQVuIUQ6A0W1gQWur7s/CCWx6hKeKWurUYuKyWE+ChF6EXHmOfWA9
7FiW2XC+swunjyOgiskOWlGY4V2JZP40DwYjA4asgOlLkU7Z7zHnoQPDD8mV
+bw+aH0Gx1z+b0ZiXTUnXVQoc0UjmL5Jp45rHuI7N7vgGuFjOOTMnpEyo+Gz
P8fTxwYhLbPe9/z1xcPA4EkO0P/R2TLHs3W/ExFIH7mmiWkXCPHudXiIeto2
Ee92q3I7VPSp5wQ1kMb5KxlAEYuZNdMkm+vj665rsiqIIfPq98o1unbQFwAX
1wyEnl6iLiMmrQEaKYm8JP/Dpx+5lEXFnEZ5rU4e7uVFFiG+93UKp7bmalc6
+mv+dalKlSIfN0cPG0wjrYsY+qp/rtPo05MFu6+hD1xtOOd+iMqSwgyXRGA6
GmGfNjbTESGXyeL+gMP8O7CcnYLPsuneV70nDPYDgYPhN9QZuJaB+GvQWSn6
rla21iUBQ6O5xIHqFXPleZY5jDd5r+eXoTOimZ8F/o5onHEly1N9EJiPOwjO
B/oWlQSAsBO+ac0Mxu64ygBiioj+1ZkLU6cSv33iuAd9F65QFTldUfO6Whag
fHl4MZOUqEdhOFSp+vgEPJ+JecLjffZM/aIbVy3+pwK63MPjr92pZKAsFV/y
i+fVqsIivONeZqMocfb2GW0hfSlYeev2OjKFfktezlSBI3UjZme94xTaE9lH
h7fN+gvMQ/I51D4rY+yekepmWpgHT6oZ7Bl95opN2S+iNHPJ3T16S+28Y7TE
6lLHhUcsQFYCc7AJ8qdRLanL8H8bj4nRHukyd6bQio+VoHVt//pp5hgpsxwq
1ajQ9uacJd5JSSshV+r2XiyfOTkS2jShNEw4Elq6gZcg1P7WWdOJbiya/f7k
No+Me7+bqjxJKDUQ7D9Z2ok8JnUeqL/kr//aSCYlO4f5u5tu8j8pIrByk1lH
Dpxo+Af4MFpnGMFSmUT8zj8Mnmcb2wmozG2rtY7bPOLbvcfZ2hYNudqU4jZ1
Qcp9RUe36afvfeNDLfn/hhQ04qhWiPlKtlIHJFhgggsglp5u+2j2sCOSAxtf
XlMQ9YB5vIXvdqHf53raIRg4c9JmQwDAMCqTlq3Hfrs7xyz+6CfhScQ856NM
NytdhBQU94CYdRULnIYIC1aBDXYE+9ym5mqXFLcTpXU4pc4ktf49dy9XHPfU
zNS7j+AKf69X6pywtJmyIU6RGLmC/n1DxanfaffcoDNKRb6Du2eSSo199jlu
vVWE0Qe1NR1d2Z5nS3YKqSJD5D6hb34XiCCBSUnzAxIK87QifFhNGfmDdCo6
o/F3Oqhln1nRfoxT4DNDAEb0SgxlkTlvnb6kwsqdCL4F8w1wtiASt2MBAhAs
D4Npn4dEQ5sKESY4KjfNlv5M8dW050quNYJY9X640tie2hfTrd3roUTaGZY+
pQgTlPpAfQg0a+IW/E7rb8MAY7Hw/VDIqtE6yOV8HgnB9x4q/ytxt5prG5Ik
IyVByAKH4bBW3PcrQvQQxhTVKIpzzmpTrXQ8TDL3xI0zhp7nGZRtodPCogpy
EU1EPIJKJC6FGvY2V08werYAIM+xtXeVWlTdtg+hdd+2cn8fv1BEzA46yYYn
9Kn2OMbvyPhvMqsy5BQdnHQJ/DPKnviM1f35HKU9OD8Xi20p/BkW1tb6UFWQ
WgtYQeJ6qUC2JlpEJPmUKWPcqn28F8oDWDPSKnxUeiTU2FJmHJwltLUzaI53
3Tp9UN3ReWOztY8UbiaCkapekxr370fCd0XromIuzFxhF4DpVSF/xvP0uetJ
/O28WCeC+UPrpp18d7whK/Tz9BlLuRy/lSeO67QwMHgIixHBeQT59v+z04GL
qqogIJpq2I9xMQ2f26VwLtPbIaE2jFZzNapUlryQ7oeQ9jK2Jh4GaXh6OHJE
kUzSnBRhoBjP0uQ4ypOew3alZHfahePSh9s6HaPLmI9X9jXUfw2EL0oj/NDk
/2oJ1sRJCIRuyTPi9l/eopnuSshH/1AmweaM+fqWjtnCEyxfysuh0BBwIChM
im3OTyWGzOc49C0/+oHqDjNCJix+6MjPca4WQ8C2bo9WeyKaCTdoM3xUal1V
caW/8fUZPKeVjviJ7xjTCMAaFaB7YsrIaUB43VhLl5eCObC2MeQpQibHu2/c
MWYfM5FYUd8Do5s3ONk7y/nUGfmnElNFAKJU/G79lEtTgrqgvCN4qyH+WyJN
q4nRHhmeWhzzySoWzpAvxWsMsBmyysgLo6pkrNf67x8XXoXoFc/YOyCuCL8O
JOLs6myxr7SZZpLCJpmRrRR/PPLlhGWNelx5hbiGTxZMFp1BTigPz2uDxLB+
nMV5javwowGAp96WV8NtxS8E61zFnPHIqdwKfBhqav4kEWjsoUSzWyMpPDHS
6rMI0N+DWIu4bRFUXtMwsmOuftQGkD739lG05w8I7iZUcIcRoUkLF8yKxTwt
E7sxnDEC6M5m28uHpCqeHWxEQJSeONMm765vIJnmDqFqbEVF/t3UQ/AkX29O
U4FjqCY5vJKpxggCldOaunX8Bw3l/+bPK/kLhjeP+ZZE0RK/jkqLt/AMIOQx
zHhUENZiOi6LzysW3WPAovX4qBfIPTDHp5mTBQ1Qz+fuUhksVb0h26vX3kCA
XGqzVY7m/UcEJBKrdKNIYeaF7KaL2fwFgo3do2eV4lpAJfJOLYGiZMByBxEX
mVGOHr/JTZ3+un8kNW5xnlhBE8SXmis1CQq/wPCSjkqnCTM5Wes3i+CqSQkT
gY6eLBtoAhbxkAT9Z4F7ZjMQllanvI6yNTzeBuoYI5bheQvyzhURfv3ZBRQt
DWDvrLTO/5nVMNBEnoxO0NTRleoFwRSsBdzrsWvcK21//u6MLE+PJrzguw5q
1KDMNqf+gVscsvg8TSXzxgODm4WmyXd8/QB2YDakTHEozKkm+Oqymgb/QMtW
/OUTGapn2zg7Ohcx7DUdekCBk9q5sUKSGDysRYULWDbX/qdxgZ83pg5zEolI
g6gwlV4EdEm3SXLYqHxXpmve0Sl5rbYkUjIZ6Iy5uWdX3Xk/YK7/HpgguL0Q
OXc/3IHgM6ipUmg0xn4uu6q0HC3LFDlLlOv2BG9SyjHfPxTor1kTZZkoMGeB
i9pAoK+tKqjIlp/PNINQE1MPdW4vO7FP5gnzdwCnHa0sjNOSWZ2r99pJ58U4
Xg2PykmoDbmkfQX32K6A6/O/IGOLsK/d0ARXJ6JZSPPI8YAXmkaVwoyXmmA9
yJ4mfgVk5Zaldy/K6f4PwoSkOxfXmJZBAqvBGBIO9jwaPdGLEH6YvPCA3uW3
uLcoURSBWIQeoFxKDgoZVO4UuD9tpFR/G/d6+WvEJvzC8FI/fA+JW10y0BN2
cDD6M7IJYZalt+ZaxohbLJROSbsiXsvBV1fg5F4ulNJwWvMzHma85HvtetF5
2Whiit9+uWIZI0dpd4H4vrMXFiH4oPPZS6Eslw3JG11fYgRcKbEOGLFniqiL
5twj461jBjpa1Z+YBwcvCdvPmKrNgBmiXowKCeBoZjnRiKde88SzLElRqVzd
tZj5+FZ6nQWJAwTHxGrTADbXcQNo5s7jh+G9kL0zDLUoJdOdCm1FFs/16s8r
mAPltoekFKzyzR2A1KhOdcKOksuSyZpsJ5ARkLX+IzAkyHfGmhwXcN78wps2
/MnUGIUYpMdxMJCPAoqsG90kVWgD0SPIpASF5k1W5fD0V6uqE6vaNSZHzgO/
eOI9KF0X174GvKv7CRUX/rGeRKKoupSiL3FNchZOg1T0z/o5ECsFre8z0bXe
WId/SlEHZYQ9T1OznPMpLfFqqhlUVNPpBeUtm5WCcsfeZzUUTWfXOJH4nBqw
FSoDKRhWFAFY2xYgdk3EWaa9rAd0TsBd8aLxWRtgZULDqGXW0oRpzJ5ntPt/
ZMoRpO3U8r1u/B4k7GhMXPdxpjGrice+tNeQeDT1nB9ou8ZJ/+pZFDul+gzz
8C3rYBVSZe9wF/+i4XNCZ+B8agCxjbtOaLEPBYbhe4CO3FyntOQ+u8lPUN/7
9uhOctujPYawyOPKguS8oBZT9U/137p8MVwTIgDdFN8FggR09HZGVhzuwqhC
pyJYTR8JybYBaPZX6NuKFQgPCIvRAp83bGiwOzyPP/R2cZ8Bo0VzlgpQNBbd
yVqiMHHdJnsu0DqBFK0+nPSHSYlb6dFyaUT6xjgQh25/IFMfS3NcuJ0hp174
tnz7BiEX8QVTp5KX4d3+MQW8d9vz/yF+EqOhxUjZQXTs4u7BosnRpY9Y4i/v
fXd9wU4nkUWZWvgCYGLwYNmzO1f5TFBAQu9tD24d8WMAspWvyt1xBAYOEeuu
lcjl36wP0SBfYPsVXGEd1n+JhUE8xB/6ctUME9IdsKEa3fvXFF/tJWTT3JLe
G1sWxP8Z+5h+3w3bAziZAvzSfikrxicgtFUtBVt2Zdu9VO+cL5M+vsBTeXy4
KgRJ6Ja+yFVPuCYszp1IfIds8n9zDD+bakpQC28/+wXxC4QoDU1K30JQBJu+
rJMWEZNhguhhkHyINkN1zY5fcjcyuJND0DsbzG+Mv2Lq65awaGPnCGu0E7tN
3UV2rQOlnHE50qLMyrCnVChX5W+ULJPJ4rYnJf+PetnB1lDLInh8A1LlY3B6
luNlr4fo8wyOtRaFFwuKWmTjxmYiypq+EucN1A3g47dZnEENahvNX63LJJ9u
SXT2WXedMlaHk7R0L8R+/OWfWchGll+hnjZWFHsDeUwYcK/a3n5/V+NRQf0M
zSy8ZEO/PBvZ9Ohwx9v3j0chhvPgN7ZSxPBCGKFPQS0q2CyIG1XGXCkRzeks
cAnYaAgAKzpx83IYSD1iNc1/DPeg4me0rO5ae4uVRu2fWd/aHgCG7bz7RjFt
N/kwvpQ7aPGLtRc8f/nW8r5gscGLh96Ijt1L/CwIX5tbOodEm9oIXpsfu9OM
gqs/z0qZ7M2w8qfQvTX1K9SeiV3CoFh+h8FbUFxQQNzUtR100PbVMLkh+cGY
g7iQicxx6HwQUADVmmc/762ANQ9a6SVpTokEwfZ6vJAZ0jMjZiFyjqu5aDlT
W4AIFezz1+mJuOCsTDn/k0KVY606+RqgO2D7MxGqHld4aKOPRMxZVXk8lo1n
Pmx0pLY2dC0iDe+NZ2XxTwN4FlGw9jN9FpzdxqRRpAdDftZtNHW65gmARaPs
rnn+R7b13JCAfbBzSVpc5lBGcKxIZ+s6pyFtasQblC40opNScNSVTG0kgD1s
QMjOMGse3ClC/juZVLjxzoY0V4TnXC1ZoK9TAMMoEK3BbCfwGVNQOBQclTfY
3qllQoP6ha4FO344lYA0AA3g2fwj1GKhHevFH/7zTZreXOT9iVMyxLr6RW07
vJIzs3grktMEP2qjRq78HxR3SE5yU/rGRVRF7RdnxuQhv4/X7pkxSYiCeejP
A4nD8Yupb3VVBmw8ClYupYBh2PnKjtrrOD+rtVvFxui0/fyP0R4VWk8PBJEE
L7h2enOTIXg+9awZoDY9Mi4/7vri9EIXEhozrEefat+F+BgGi/yuxzYBu9kQ
nrRuslxRYEpUSC2dvzJujAFdHSxvsdcGCE6tNfklZidHxzbN3tKuTzpfvV6M
6266dkiGq4b4cUOncbSIIsiiXBok/WBS+QGOVvgwdoYEW2lvpkgZw0jhEMKb
jMy7hCGBhcNUoH9g8vmVMHsxynA7ltPXg48exvDiCGHgTDXjzPLLV66/tXbz
HCb/wHYzrbFvN0rLJL9M+9E6cTQ/tkqi3S9Nf4KCqhYeszg/fafzoS+eytnp
y5yH9crLnkVeHEgNIlcYuDfixbEsccD8XbNvTIu3c4k5Buyn3u2Ry2U8LzET
CTPtlnTZuiW5+AYIsvvrsoB7P9dapqmXbx0CfUI0YUJVQzLdgdVrXblDKpiE
d9KTQ0a3mt+CZzp8qTfLk5DaJq9sIjIL90D5qqH7FDv1d8Nh7NaO/H9oiMaB
JalSCPtNs7Ok1Umqx6mu7KYmxP/5XhNnJzYZGrZ2ZO/1M1+0H6+vC6Tygn4u
56AuWywF+y//KtwgdOnCjEqeQEttGp/w9d/ahSoxwxY5HeE1PZpzCgNXJXLG
keff2HO5UWyJyzN4CNOSCyEwJE/Uwbz3pMSxGQqitHjrl4eS1ExhzDMVn/4o
pK7CLwUnZyUgk4UHnbNP4/P/oHgNixPA5FQRC7D3qNa4FX2eV3BIR48Zk2N4
px4GeRms2sFPdsAy5np2uwRhTTcaajZelfo+TRHBkEJMiwlk32M28mc3VEvQ
m4LvocJpM+Ce9WOavKOKC0mF6WXFHWOPScuS2XZMro2RV3p6l4qfph5FY9VP
Y8pnbVzLnlih4RLzlhtg96Z39o00jeLD97xs2y8pf++T3cpQORuXtX+OIqx+
hEfzaO520kXPPeycjbq8Uf7XMtW0SWtWdMUCbowk1ibtbdApOJsF9tdrY7WZ
S/7B80av2+cNgB71TN8EevpwXqK6ANI8C0IKyZpYIGIz3QxKIprYEbCuw4fe
dB/0MSUi/MJOs7BghuQ8Wc81ERvpl6mUDNinIQ+NP/Oc0E/ag2ymD8hm2IGx
IxnKpoJZTFglA1dJKoLq1q0CMBdDZQ0jGtD7oVf6HEXq6TKpNkL0eg7jQMP2
GtIclz4i9EUxMBvUZjXV1y3wek3withw+SF8DX04rlbpeefE7vOYDKDa+iH7
a6es6u8odNVfAwlkR5bGsUr+BlcQuDQ8Mmvyp/CS/BfDa942tr3co8o/P1zZ
tlL3s2Kz159JBGQlwfHumSoB6rnVPX5jEw2b+PyfgS4/Phv5dV7dUxjJMwYR
NgsPQY1XqM6TD8jxB1a3H3dDgF7k5nfukZE6pr37DeNVjRA4tLYnhghzQ1SH
ALwNZ5A2a6VOliiBEzq2evqc7yE2GWKrgQ7WV/Ia7NG2UnaicbM5UUpyeul9
+AVNdPo1kOxvWiqYkWOsikaTxnqtUHXjKpW+ssXOf9ZP2daVDPeIYaxOBFdA
QLDpY4UjR468+dim9I+PXz8YEp4jVuatEkSCRRPvy4fW42MYstIijsbCMv8C
wtknqU2GHVUjkyJvX+UgR9EYVs0F+/8O5KyLaRmzVu1kXH1sSP89jExf4PVj
niMNipydmNsFOSXlT3OKeQrvGbxrkgPPB9EpfZKzLPWgWJLGK/c5ZpoR39th
fBwqLv+KJPwZzupvp6pcCX/E4H8LQZkLKZDN2v/j4xRbr91T1/216g3wmFu0
Hot0GM19vCBmjAcGQCC2ldU4NpFJTS1dCO9TvJlMQpwbqTG6gFAx69x1X/M0
rrUx/OQGx0nRTPYO3x8bIDedSO8CzeP8AGZaeXnGxxmVUhraWl0KIfl+BVDJ
Lczyl/G+bdmtbXPV6rp+g/NLLJM5ucQOegpcceuoKAK/hBCf6EQ4d2iy9u+p
2fL1zWIl4EKfCKReKBlS1Isd5RIEKpS5tVrGs8PoRc7+p1+s+0TU967Tkau2
GH/g8mgaITeCrFQhTU6UyaFxmYWnLwhYgokcbuK11TAgl2BWn5rNvZgSCY95
lgq82hv3V9n5st+c/o6FgpDdh43fg1RO5jpIsdREFSpXtAfr1MvTNy2gIRdM
614YvWTZsKSkq+gNgA9eWVBn/xTNBlgGLnZGsOW+PFlRaDwk2sjQmmR1ictk
MM0mmTtI2fbS4lcC+wHdY5k2A8fvy3UoA0q4Ro2+xtEBi/f6dCs3EmRP2Uoz
f38MLx4IQtxgk997ztrDe+ZEct5wBzUyb+QhnykGz8ApG5FvJYcNJVkXicMp
2H2Y5yCI84d+VIrWLttlhvPXyuox0/N7PIJH1y8tyF+cHjfmjIVVdxi3pk0/
wyyNW7Hk5IhllPmdC3S3hftOJsygpAj/3U6iT0AkcHlw0pE52CfOELYGyGZy
DtykZDlK7Oe0N1tw0Y8KHXWt6daXJagVNaBz7PeyUlgBl9jbbWEvLJWsAF5W
0Hw+CsO5wzNAQau6iXrtOt1g/AuIwcz1ihuNUfZ1Vu495Cpcw2vlue+ZoqAR
6F+bvTRpqTcwsc8K2ooyULTez5GDj3IzrpnU36DbfNlfOhx4ug6Vy3EP2xdv
KhvLgzxKWlJToyx0GeE/7MRdB43RC2oHthtlKUz+XzZcw6CbMIGCxQA2UpEP
AFnB1EUGAiUzxYqIVrAk38a4XpIDsglxUyc41gOn6V5dRlhYCjUZoyf3RN3s
A60D9Q60WmDmMsNlQDd5q5Nz+4UPHKZF2YULZrkDWzUKrR6TGkWmx8XZq3UV
E9nlktdb7eJId2LXdREEvbL5fZbfHYUgKJRe76o108Kx6RhpeY86ClZdsmJR
hLpjxHjqTccbzRKoK7SpueuKPF8IV8flFfjnKo3+vfv3Rvh0OgHl5ucWKJVN
YrODQ+lXJ9ncP8+Y5GEDdFu0wXpcqmAM47EtgXAZ6N9wmGvtkx8hW7qeiRzB
sk1a5b4P/abyrmtr9whglno65+ocvU5qc7kTwCwmn6/WaFzXMzRhVMGvrwXD
/oFgG/d0TE03pIRqPhs2mVYPBmHMzr0KDE8HJ4h/hmK5rnlKOs5Cyx1HtQ5z
+ll/0mDiWRb762JvyAP86b+ODlStgxPyWP5i+GXgkz/BBUSL1Jy0Kev8dc/k
uJloLMImPHE71/oaISaj0xQ5pQ8jD/sBP9BESZqbmyspcV2f96l9NzwnjSVh
r4UvVTDTy3HiBBRBF9gB62OUxhdbdfTX9r7+ody4bqgMK2bqA5zFY2xkQOyh
WvcMmf155OT/x7VyH/tCqdHMfeGkt+cRi9Rebjm58VdfRN2ZzNuxp/U1xViZ
oAom5D0rrB5iudAV0gNVvkn3hJihPcdrWALL5FweB3E75nvMT42KfgOLkTwP
En0htLSg1Iq4R+lXeTpxrAOQUtUt1pHCee13Oz1pk3e1UfzV+sCmlDzwIXOO
fVPyiF1qHs7zehuQjecnKkrk+2BTGhqZ+XcnjpvM8WzZy/nmwtAksM+A3u40
wNw33QmEaB5orPNco2N9KxyOLmc1yb7dfBqJRr9U77YO6oTch33pqUZm4xNX
DNAqkLVYV0opMat7fxKRjLNhmuZNrFIFhBdHuv5EHir5lPtGrHS0xx7Ut3yY
dj2QSYMzzgBpp8AR8qV10PXvqpiodH9bi8OLhrtX28O8kXQCh/Vm0hjTEOrE
ocSRekuzEP+7aXkbZV4i6soGRCAKbh7H0CYmUPyZt5UfpujWmibnhKFC1gGy
cCVJCx32D2DaXxraUnlCg/BrxGhYdVu+JgmVrKws65VPowTCiY6lwx9G0cRm
VDD0WSUUajiZ8KZf5tnYxmDbnXTZ3k7j0boch/FGdDuklDfCcpUXXRh3C6jd
JLLa9Jokg5cwFzavWW09ZOjAaxRZdpWEHx4q6NFUdr/nXfpzVgFcV55znvtO
HlWKLcOj5AAL7bRztbm6L4iElk8n95PfNFlb4vQVRWCGpRvZaPwx6SmDyoqp
1efqaTE3AMiqI7/XXkpiZKaYDECJxlxMjEHht+QTGJD0QHxWOoZlEPWjxv3/
XkBtAWwjwKgwdRNLPr1MKdcHcVdQGADR5Ghl+ClFXVYAn8P1tdH4Ile5JmKS
Q47/OybfdfJvO1uOv3rp2hsU0OzZWZs7xdbW1D77xqo7FwVWD4M55TN8BlYX
iWciBV3GNpwr9J23LHYTj0EK22CoDc3TWXl5FGQ6+Joup7EOwb/Z677vg1rH
9lzN30EXGDok4/HmFxwowCgngbb4kK23gFquIqWY/IYeaxU92a9Sl3C+JwMq
zVEotO1npo03E3C8clzJw4X4zKM4OpqTHwiiAK93CeLHCSWdHzdT8Llv6H1B
egbAUs/U8LHDeqHbb17FiGxx9sb428JPXpfEyalhHMURZj5rZnXiyTQXqPCY
lmTApiMxrMs3ITb3k+su202bqonGGH8O/2BvuRxvbYyNsS6oRBKLe8J4TBZn
GRJYCdmOU6XP2Yw65iJyEaLSHU9lsGo+WU82p5yJ+AnAKZ+oplT3QAuZG3N0
nwNkmS6+xMsI0fyKaTd+3Yz8Zz6oDbek7uKXy3YlV2DWzp30/5+GrycJap2b
CZu3pg+PlBtZ5dcWtIDKe3A4Mvk+TbWYQcdW6GJFoiSVw9bXqifsi6t/XLF6
k15RNazQV9whMClmL04OwzkC4LGjOlGMIgTYjqbySZkJQw51H4dmsq1WgnpI
Z2YPW1GIkau1C8A+TRZyBOpbrC6iUAH1tMsyBbjgXffEON4cEKGnLPicPK5L
iLdIAiCVVEW1FiUBbm/wV4xG1HMaJtqWDu+fik5FNdk0KuVfNJwgGQVVxtJ3
/DnfbmAlYf6tYZuxZb3V9BzX7P+meFm2isoeU3HaK3JEpepcyqVEiP1/SP0w
ME1+5TslyEDuotmnrLZp/bTxsAKyWQenc6/VSUU4V8ZPPiwO0pg/+4/lbFgD
5QAyRRz+agjea75/U4ceARtszOEjqhXv9toLdCU9JMWED5nFNuDKEyEIdVx5
aHVady2hM74McWrx8b/mJverM71m2AQ0yMEQuHETB4LTt8JfDPjf3fTxDivB
LoEoW58eNiJYY9ipfkmTyhEz0YL/V7OO07hUiKdEUE73C/8V+1eOZ9CVUz7Z
JjyVq+7xd3Z0QpwZ0LChJ2G9wKhzfWdM1oC92+UIF0xdRc8YCx1XjvXzJRNt
lVBJBH6lr3b9tTvfH81vYxjoVO0KHsVYJUyVtyEB0/Lm4shWwkzTuQhwoRJh
jo39DTRQAlw+PCWjtGXijsI9jDVOFBXRAmo9EFqROJoRoqk1mG0uIBOevKoh
JE2dEvrn1Gw3tDNzM+ANBUBq5njzjKTlhJmcZOKABW+vhkRv3D9xtAiBJdY0
BHPggBQ2w9mb8+mh3Z++YG9VdAaGSIh5L5/u7GtupQkemMN5pk4ujJOw4Q3/
RrUomHnCwT51XOyPGq4n686P3vkyb/i/FK4GLcq5NTJ5IBu6PnDyu87nHvq7
mGTKM8HvDl2za9FUpRnhshVOxnSG7gzA6tlJ/c301D2q+ucHHSVwYWHV53XL
B1i/f6iIfe3jBcHmUsEgqeIw3m3J8cR4A8BtOeyR1eyi76PcckijP+/qa1w0
Ekf0aDNFVZeAQjsXGToSJu/q97EKtuUv8PnlFop+LVOV5ZS+rM5TysXYh2z2
3H7dUflDIPlBbl7vkJ9W9d/no+DZ6aa87bRwl8MKKzvVnU+wMpxRKmiTBfl2
HS9koCvCb5U5OjFMWfM3/QKhRIIiQ2YmcRu2ZUpKeVoOtpRZM5xnvHhdojBZ
+v7znkmoHy/Sggi359hrKM7BLETAeZ1KI1T03elCV0pCkKcL7AeBWETQ/SFk
+jLBlrs+fNzf29+78sQW/KkAvY9WeXVfT3vM2/SL8hT9oWLfZggS/AhlWiYG
K9pEgA4UnWNE6qu1qZ2hp16zkUmYuGeDIXwqrx1XCaWoAlLfaAevumUR9t+7
1OBiRTF8r0NbBvZkP4ai+DGdwg6pu+XmnRR48FGRACo8ATvHApGuntymuYvE
9Wa8gi0Med6nvSbeh1RAfoLuCZUxhWl9rYXey0ZErirgKrRgt8Elm4qg3XFs
d2SUwQ/pVn30pwOpq3MZrcJmYTmwSm9bI9mZV2U2AIGWrnRD/YBeaRgfWB7r
yXdFk9xKJ6Rd77eP5vBKks4K0nmvH7NZdmDNVapPjsh+EwH+OcHU61RCJIdh
aubmP2ezXaN/FG6Q1I37lnZNZEsKTwcWOipiDUACmgRA9pvGvfVQtnfDniBu
isB7A5/VoZ5k4wUe+ghLsGi+yaHWcqItHQu1pdsWoDwrkEEckseaO3HuK0vY
URMYuILm/lwCO9+PUC6MqCIcvY3QjcZaMb+XUWx7oFjqkKiCO3rr1oBx/f9W
jh4wOBKuLZTLwRKmDTd2t+mmPADyQTkpUWFyOsLis6PcIcYJZD1KNPSgbEIK
QgWOrID6pjnUnNnChFITeMmhoEND2EwtIbHME/vnJgeOE8oiEvR1DnmLvLvZ
PHVN4UqJng5rG70V67OHhmz9wh8Fa7KGQdKeHWTN+PA4ZYC3nAIejp3DRMqd
L25Ne07CP1cckaufCHqdw6Xqz4Rf27Gypc5BKwwk0M0/Hs6sfPv3zchB1D68
afZev7V35zR8J0vJ00qHr0WGIvDNCMGc1iKGm6U2539QHyTwAi+uW3V2KBPo
TGCBSLy5+4T+pDvsT7Q0vPkNJDi7JsZc8h6OYgn7VzB9TIMkLc6G9SUjyKxZ
mB5HKdPnifW31GyONnbBfsCyms8dvWXYCRCrW41uBDFMZjRXV/AhTQuiYtmV
DeiFEZFVl+ln5LVxlmkdRAOzIhkYbv7uaRf+20hIlSDwh6BblmkrPZWntOv8
x0mayjC0mev4enbhDUzxaNXfQTIuyu5DfK0B6fC5qBVSBrrGbLOO8JhJhVND
E1LXkmfKIsWL1BrHTb7aIpz44iaLFIwuFQKHvyzcLkqOlxbRg+BynTyoZZmX
TjzxlQFtu2u5mGUKDkpZXfB8eT9RqVvce+ZN9NBWzPlXB4CWbAkmPZB8s/WX
I4zBf8N5U6N+grOii87HPoA6hnl3kTcPfb9n/H2V9GLmaflhPPfSKMzqi3eR
aRWDP9Cz7HQGj7V/qEM7et0piCxDQUK5jROOF6584T/0bIA3/zhJ9xknM99D
BJCxXAGICfOQVpux1oI5QbXOr6yjwdDCpzCgElFJfT9j3JKxMiY3Himcvm6c
mMbwwd3yCyD+NDKZxR3PGIDmJBEUR3x4+M++ZeLpUwW02PC6OTuipq+ayiet
P9Ak3+beu7cXOjBx3aZ6tQne3iCRqznFPBVocmlkt3rYBsJRzo62u1RPVkoU
KATtI56zxefhS+nevqLBhAvfu+1pffyQvLaroRz4e5HfuFy+oiq+W1HTCey9
3fY8VLzV1tEgxt2isTSZ9DHBIIZkghb8iJXj+wag1LVJsVUjAt8GU6aYTIdO
HqGEZGkTU4BbVkA1hFYBbbhoSzsHq7l7uqqEhyOmEaIxWjSoMRiGoP/fPs+s
Eq4FIBz+gOoCYL2tk02YsYH2e09cLgtlUKf6ZuwBl1kqqx+4qYN+RAbd/o4q
PYPq9qFnxn2+WOvwFnGkDtZuJnousys1OO+Qq+zSWJ+k8J7tPjXqadwYnf1b
ERAos+f1mw0UNCCvc3aHOazWWlpNswqAF+zwWTfsFSqI0lZgOg8gJXknM6MY
zVQYcRnIybzeRCrMOxPU+Wl4HdwKdXOcnLRgUCy3UQNODdNvMBbaqYTDHtCE
jrCv1verneaAUwWrkZdmUM2gOs3T3kzTBgTEom3g3OkKk8YIUTccc8zdyRMj
mV0tu8xgiELRvgfShu7VBtEsTeKQODNIASlhe41QOMUm5fTEP6LuE+yCnWLk
hDMqQHFcE5vGbNpUZFSIK0U1qnWOZwG3mLdKUsbMHn887hHLhJWT+17Y3iyl
fMGaolzYWjsUaCRS924+Dicx/CGIJX9Kp2fFyElxwAucBbl6uKnWzrwHj3LI
E1QVKeBiyQpV/VJYiqaJkeX1Qhpe6oIUan52+e+0d8vUZ+2ZEZnO44ql6uNA
Hr/+IfWkSUWAU6PV9wdhWTNlK01GpNJbIw7qWdt/LB8UyJJfzPXnRFp86seM
UvrSO7O8GLN+Fd/8EiDTeK4M46pPaz0pEvHj0kI8d0yEJOey1IHPJTgRFnJD
boUSpz2XAxg1YoNQfkSxszrIY/MMCMFWeuPEr7mxzxFU5wNF3Uv8Cq+h4Whd
kbnkVaxIHQ5OJBYx2HR+YH0EZHi4i6igF5gfaYKBOMGy5t/KY9+QCyw/9OuJ
ReUIZTiF3X3s8XUon8xhziY15K7SACloRJwNuGsf3uQCr4DrNJrX2TWKYWPD
TD0Z3Enz21tbfo9CkkML5Uhn2yimrILjgoEhR524xtaG1erxsUhviE0ZB2b9
pritRxP2CeTMR0IOM1MhXnp0eHPsmHVBdiOCQNRR5DBlM+oIwU71+HWQW5N/
9sIe2YO9KRJq9CdlJhtuaXmK2WBeC1sNjzVoSpQJiCN7nIqqPZt5PQaXCDLV
TFC5lUzVHqysAT8d+XB6C8vAWBaUWtuL66SQ9fyN4zipaj/0MmBWY9O2om2n
VcjNkkol9VJn/qxaXnRDby4wxg3VSxtZZj0i9RWn+SqsRLaOtT0oOrEFdsbm
OjYADdmP4m3Tn/XSkVI6DMzwPSWG+o4OFrNPAgR02OPjPy/Be/UYsEWiCGnD
4yEMgrjHk2WmU+N50t5kk7RvtCHKTwqoDkUPmPEw5f0Yw7lOU33EPVMC2yBk
0WvYiYqj7dIigXa2QAGcUBIhSBI25qEfCtZy5P2cY6DIyriLk8DmC49TOcSy
Jm+ebl/iVpC/nQaXVy9y7D1axld3NiqYTKNIISrzqgimJG2pHCU/5Yl2boi3
FciRxNAO61+m8ciMAQn1W1M4AM02oFUJ4bdzMY2bP22YB+XaQSjqFzgPQZaB
GkxmZpxDAqupbSfI7NsO6LDuwMc4VuY6WsJDHLrd4+9ep/P9oCVzQvPjHwy8
zq7haVV+Tdw6B4KPqjqgkTWrKxXLpnAWrRS6ekwA8jol3k4N1pjnQE2N3sx0
wx1GksISeTuYP5uCZI9W5sRx7PIPvc64pUa+3cpfaWVMJErKPlCjFS4oRoaL
3zQf7PiXibGiX0Qtl9SNK1KyJcFJK6LQNxYtXOxNuPCqqG9/VcffYGlZsUYj
fS/BnznX2UP8j1SXEzXDbGNBFUwfin2RuEm7cvoa+OzdkTwsjlGUfDe82y4L
Snplg8ThtNRFuFnXsMEcFQ2tyJl8vPU9yZB3gVO13w/8sb640yerfFqy18lB
fvcw2Du8mhYJGTUXf0A2kok+75orUPYR5zCHDrdqY/illjFTEcketMNFr3Lo
kPcERgCUoimwtQZDaIvBA5g6zJZAk9Y1/QvbcuEmfX36BkcmsLTSbDi+FTdB
HzoTdnzTxXLzzCfIp9MtPNgkv3pczwlODIMwkhIJ2XKljmqc643vyPFCEV1r
dsoHEqZyIiYpPYxK/P0as/nC1P8LFXbXREBPVGEk+zlCN7h0qJBNGV0GY0zq
wHdNqBbiA0pUp3wetLIFnLNdnRztmsWSUA1hb0hATNAJH+f9nvk7Vfp4xyEs
obodogA/aFbwSrxot6wr1+1fpOrn4PRYVE/3anba0wjuz7EtL6MkUZcugHsz
MTncdmOA5fUkGRzIOs2cX88KFkwF92eKrfgxl7nnBQaFnHcX/HL7Xx2RufwG
gum3fdeNdEZudxMJB7b6jMUMFOvj76gR2lSRNsawjK6AgoUZJPT6SbfVvByy
1pSnVBPVziGn/f+pMWh14oWaDkz/ls5aun9O9LdIf3wb2R4TLNOyhEU2eBJx
gu6irD+P0H94kMq7Z0Cz0stPSBsVzqhn9xF8KNLiInqMpHiwXgAgk5aRG+5u
aaIcgEdXkB/PRy6ke2Zi4YD4Cb5XCfctpTlR6sKCiaN6D2M86ROWlMsgsAPk
33wBM3TIZ7o7xEcjIHIeDNNmnmLy+GZ2fJSbc9fMQ5FrY1Iztt8qIOB+d69q
nJOQiXylsrdWqbK432dnaWrLg4q2PBRwO3UAWqBHrv+URMkwCOvbUl4tbHhq
gLVUfrARNoR2Yk/J483tqTXfU7qv9YekkrLy1ELA3PMnwlSyQgM/Ots+PptR
/GN3cWAKIkOpl+KXxUo5+q/2bN9vzfVfe3ua3/KD5kqFGRADUHn2t3h4N3Aw
NdU45o17D0VqOPdQzoKBH2epTVzHzEfXOwUsq1TXmamrttbTO3pQFT2Vuot7
YrMVx/F+vRId6zQFZFJAobwTYzZe/pTC6FUs4TxUFPL//KO3BshVSXH6+ehq
n51Ijc7qo74XMrzUpDl4Ov9Z9JsjYZpbWCl87vDpjDeJg5wiUOHhkVE7E1dd
THxdlFTz8mo0gqijHMkpqJGgx/RH3cG+YeM9VBzfpFvvZDs195ZAIBo/EeKZ
mK12YaoVd7pDREKfFEiZJGw3zf29R06yv72J3ULDyWdu+t67m07Repn08ozG
y8BePuZ4fF/WsvxnzNoiWabjYwnHptBcJjdOs/udGOK3VHJkqbaWA3VLuJEF
liVw7GwxKfM3HkZh155IujpZBeBBIOXM8Q+MaE+bkLGqIIq07/lzNiE70/mV
IMubkybTlkcAHOBF5s3wKB6k7EDbv3T8xGZCRalloskQLsjse5M24ohPSXIR
BsZxjg+gH/MAi19HBUmDTcczDJCk41oULZt2LLD45lhqiU+fNkuWr32KSGm8
mIVOW6szsQnqBxxygT91M9tPq7yKKbw4fPy1VE2t0FXqRb5rMtvdkgdOx9sE
5qvmt+z8omrgOwgcdshKJ5IYvJKeIjDcwq1/MIChMrA5DHHbJo0vScmyZyDb
o39+GNEi9BLNr6bxBIGwYdRR8zwNSMa2XZacvRt92/eji1Q2sfmykELujIwi
Q+tXTh7HFJeXVlCX8tf+Hw7jSPH8G3qlXRb5lnd+1dD+vT+nQhBfC27FNHqS
Sb3ikzhg9ZEa3mzhIF9E59ZHS7ty/XNiNB4NhQipFaCAZfDk27GXTJvKz42M
PGrL38MOeONcXg/ClY+mQEThsrR428GZ5d5wxdonIWpbeYqtVbGOzUuT0N90
cXGo3PLz6TE7U3QHyC4L3m0n62fFtqKTCq2941KL76X5EwfTVTzLTpzx1bKv
E00a1yww8R+CgACTMz7uXOSV5r+5tt5nPlcRaxzONA5uUnunor7NXhdPZihh
e5fevjtE4urIsHK6i1Pvt+4XvOT4tZpYHgVt5b5eOQtJhs4rgWyiSwqQh3qN
D5fVtv2Rrgnm4Srt/OZn5J4aZncTViwNU7cFRXk+zJBU7OawQGEVM5++DXkA
ME899JM20Qz3CxaBhfX9Zq417JFj35p8u74B43nvU008BvG9qhi/cfsUXMcZ
OuL5Om52HKI5WWuex/8YkbhgJ8p3QTlWRIhnjoRVJZVAQG/+Irr9KHd2JPdA
kGm5604yI06+xjwWKjf1mQWBWULl7mstrloI2p9+YjFyjrCnY4IpM8YTlfpI
Q8pKtveltMzp0XH4ldKWCcKzfSghCl8cFS13sCWf18Qyky9pr3GDnLUJ0uGG
PR+TPgWy4LXFLKwWXxdnq8yE76Jgoff0ZRo63fKlYp+po18Yn6UdkicW58Hq
JOd15SszemtKD77aHSQHdEh0XmcajOOG3Bp/MgSY0V97Wv89DRhbtJ5gaFke
wfkVLe3nU0sgr19B9ig+yPbr7huh25gaNmDobNKeHOYi1wqUOZX9zBgmBZdV
kfYOZqieVkKEwuVjb/q7jIYJ4WpRUocm0uBBeUf0b6neg8++s3l0rS79pnGD
mqENSEbTkwJ7R5Hn1jiZQ/JpcCVvP/SnQiFFAw+CsMctuflYodmbrMKxtmmx
SGfCVImW4uJDiBEPH/8I7x2Hx0NveRSl1zAZx82+n4cs4kX/qwufqSfrbWh0
tKCoWTjEX41SZYr4WEbGKh++Ex+2U9d31gD02PTq4rKlAUw/ybYkA1WfDAty
lK4ZDJpkZMwOfRD8lHY3k1qQ5UCdxYhQb34vU+EgCDyUHun6JfFvp+4F7Rto
cAcjKuZsIAm09NTQYXrltxl/7DeF5urk7rpz1HrI4JeFNhLxdjAh3Cn149aA
7FnxJ1bw43NvlRObr0AwDVrTZx7Cf0VK4HFOwbpw+VRWPQC4zvwvS6+lKnbq
7n6sAee66Pwi5WKUKXAZYwuF9y8oe3zLskQ3SM0KodoqaLDXr1ssuzzJYGt+
Bi4LpKvu9n6rpuPlOC9I0ZOEvMJogIYqoC0g2UW2uw6EmjIbJbDz0i0PQ0Hs
FWCCDUZEIe23VBrEnFQj4oPPwZkvnLTes91V1bhYq+LkzyC5egwrVZcIzQX5
UCMCoC6ozYWiUiRO082y0NyeZVhqiSmE/IS17AWGdfARhR0sz0Syp89u+gH4
CY1YqVt1CFqF52QkNPmdEwpMHa4htLSlCgxDPLNzSOKR0bj93M3Yl3VCZ9Qs
Y8zBo+k3+aOyfgXweYJA6RuU9l0V9kSPMcAbU5SaykKJWUkLVq4OSLxMpAOf
5XWXNZTq/AebhhjKrY0/bzhojzrMgRQ4xmp3HguY+38sF5HdZTpsun5NjFMm
UROXuXdVf/hkhs6zaMAmxXoxOYPWR24UgKKzA9jtSzUmZEeOIUPov07PUzT2
DSOZaD7j0NWHX6qzNXMMJiTXP1+XDZmQJM3VvdQ2VFrTnBXAEbHkzKIRUKWu
9gACrfGHtLp3Ec7DXL85Yl6pjxkA85G5ZTekRoE1/xPzfc/sCQr0xlUzTJPD
dDlH1DG66w3hVbiejAC1yIiQNiELI4jfi6/tJkch6/aTlBV7ABBl5JTzAPFo
OK9k46mN0ZfFendHQatPt4vPSOEM45aFiAmBWS0a0XZ5WZ/U5g3BDKpQxqpe
/GKKdO3kGKKEFM/nQLcFtdvi/G7+ie5XUu8/Td8+AdzOjTBxfy3bCfTKfMo2
KjxBpeYlx417KbnlvnHxYYq6P5QKRmY1Zywaio+vClC/OnqZHuSdZhC0aVHc
ZoCy0QoqCyaZUSujP6r86hs92vZsmwbtOGmErVfSd6/IeQl66GLWd9YpcQ60
XGkAf83qymuFJJT0wcp/Wo3pZYVngNGkg/+Q7rrNriEQvCOpveHPXygm9auG
MfK7X7nOtj5TIOJQUzJTVYoPKAse35OUuGVyvtXCT9s5vt0Mw7PrgG9JL9KG
6aKVQ1yf09rw4sxDXwH+HDD6jdyi1hIlr1a6pHi+pgZspY/6+5aixLJNAODo
VKS5KlGhrxVAiVFsS5eCPJ/z7Cu95fOUWzQWTfkkULg9meOPkmjll7ih25B3
dltr1MslfKdnZJok4E3tLVNaNQPm2CP796kR2s81w7JTVwSyYpd5LgPqJKU6
zrp2rjydWorP2ni+l0NIzauMB34wjEMPO0MiXRFafjMuMhHb6IKypYk5DRTO
ll9XfvXD8JT+LMtisY+Pl3Avn2zzsS5M1BdxCMGAZQqrNI8walh0E4z4U7LD
pzTVPdpPRjjhnpBWrt3K40HB9KPXMwRDsmiZDMoN7apHhyouERXu/K6XQmLx
lQLW7ZOStevJucQW0i1SbBNyUSGPHrjtoXbtYG9cHtH3TuYPAD4qp2LSt22H
/gNVFNXja+uokwvkyUh4a9cLpbK4PiruCnFrbhymxboxOj/hsEPmbuuMR6U5
V03HKq1i/ZoZuPIzH1xtTHz4UghNzMeAj4Qe66fpZxMo9s6HqJh6xWySsZCy
LHpBamoO3z7QDsjbpHniopwlYHWInFLUnkDyrvf+6NuSMnJJlGNpmO/Wpx+7
4Jtf+RBnwFKAbVNv0jdEEnnMxjmJvpP1/oOPYFMWnfX+wOk/OzqB8tzqErwQ
vLWMcKUktLuRiy1C0ATWfbObjctzIVbekJIaOeHf8jHF/fd702ROosXw87ZC
HyYtr3x1UcBNGJvAg6R3Cqqc1kNVULgjNO4IgWncTjK6JiT/vqZsYahwXcqS
LZLZSHfqVdOd3FdxF9ml6f1V3unNBeRc7uf8SaUpjy9z7VKbqzdxGyKy/T3I
KId35ecFkqsBl8MFlUfOkdvV9LJp+faC0EsfI5o5+5dQ/SnQuiHe1XokS0Zy
mhJbxN5YGTFUixZJRba7c+W/Wz6m0Hycb0cc7YSrAbKiwiFLG832F3YOWLR2
6Kgx66TqGLhWGSKOWZp/QJ2r9YgdT9Prgr+bjWvMAQdgl3I/Kl2V5Z/gm2M/
s2Hj8cXlyxy5HcHtlPZq2fWlv77IHZKYy3ueB119+ajNMWNvaDAzrsi0ik9u
kU/QCv6r/g9rUXaCUaPYpN47jW4wjBN6H2bS3HkhWvFH37yjMlVfAD9cnxaR
ktyj+1Tmt0Fr3puf6npNQ0a99rLxpW1WN830ElETYKF9tcGJc3aNu+R1eXu9
oMQqAi89PioZtLQBEb9PVFDOQPOA4iH7+l1NDt1v/LSS02dmmp0YRnCSSE15
WS4mAClhP/nuL6Cj6/dCL9Yvjc+1J2WzGzMovBZDLbUC0iRgo8aaSHVQUzce
diK5uq25R4IHoGt3ITaIaM+86zf/ueDYfwoxp6tQVKv2KlWsY55yrEEvV4Y2
l8vT5xGxXL1mnX/sc6pf1HL67kK9e5jRNRxdgX87nvSExjhZA7U4D4xd13QZ
rtNt89iZY8F4m+75wW8KmpjKktHPZaUdyTQMn6v3bCecv3YWumUQht1VCDpC
+pEaxAHUFVlcQ86d9K4fVJdmZfzDcQQCRjU1Hs30EmDN2ggSzS68X3ZcNH0w
aeolPvpKSyoPfUaoOiOHNBB8u8wVeXZ9IEcWUpXbiz/obiYoL0gT67YTuPvr
FO7S0r9x/Ze1cbdlx5FU/Z0zXSMD2L/Lq+cgB+0vzLUcUUzn12Y45TeO8GAl
xbzlbwQX8o3BXZbd+XiuSSPGWucEo2+KgrcRIbpor8+K3f8D0pWw0sC2YNnH
gQbQx/lm+xEeKfQ4y2nT0WTNbw3/ROACLI9rftwOZ2X/NXygaukf3+JG2TXY
G33jwDD63ro51vm11bSb8SL2vy6x3esJZxJZReo6lX3viqzy5VhDf0YoJQrH
uX5OjVyfmwfCLB+omTonkVWSbuYa0UB+WrsH1P1OvXkTFFZmWRHepQ0mq2rh
xpxPJqckwRKohqbYnDjchlNO32IObPqvNLugTg5wnSP7sra23Z4UPgrDxCKX
KkWMKdt0uk9ENJEUnhnNj/fcSr/Sxz1/szNGUq2pWFnpvJbqWgAjCTW1BXnx
1YIFog5X3TcDfhg2x1wZ7uGrh6V/LzIqbhnwCKU9ACscp7FJvtWm8te8PhSW
kAyhzW11KVismD+EmbNS6PynpsVn5IMViwP+vuI4NofHumG6h5AEb7sI5uie
UMcFYgHc/PGX+ei6VeKYsDQhTkBFr8LsHQ55iFe5zG8GAvMsSF50Nqx9pb4q
RgD3v2Lx3m2Uv7NnCUu9VFi3GDYHA7zpVrGhAN1Fgz9U/gXqFqRwN7JgcUEQ
78PuY+YbGe5RXOVmKU3UlAIkOgkJ9vj5ERlRfnymErpkSHyyjPzgNf0xvZeC
1czvxXqwG9JjkAlAbzmVw6778OpRkOfrtk1a3OUm79MwhFrOKWGxc98cettJ
vTf7rpO5hfTCDj7rZIY6ng/KjIDeIwaDypFZSWxYqm0yedyy5xJEnQoUSa50
gKT6vSqOau0JtObFGlKoq3Vcpn9QgFf4Oyu4uwfk8jxdleSjS5/ymyzySC5b
GrvwKATVjXGo1UtBG523gdyRmnd5VjOJnDX8tGqsgvN0qDwDA7VABj4V0xus
I+gx3ECts4UN7vBHpU3XFXJcCAk+4MQjZTOk9NTQYCdbrn3rTgssesmk4tn7
UgnhRbVO3bOZkonOjv+lEw/VTBSbjXDy1Q4fm9OW4nYJHKl8fdycfmlhTLt0
r3nAaSjAGIoMOJ5ygLViR2+kXSyRuFoN6WCp9N8YvJi/A6FKeDvgGNF8vlpI
H8nu0j2la4hJECVkDbzyruN08JV+L/H4jIRCWNU5XI2VwomSiYSNU3LGp5i1
Rgb+vkF+PtsOgHaf3jDjF71mGVlSKHQb4S967/tV6+HPIA2wBlX45V/rar9M
hRD4HbVwdjFEu61hKpcz25a553uKK9ummkLUfs5WattdH+KbaGRYJuWBTKNt
NaZvlUf4TlSIK9J55zQESDEQDbd1Ay/YRNJ20OrS0R/FgiE9D0vsFghUZv17
tTG0PUxlZYbGcXTO9wCuRsjrAdphaUJs8qzfpqlO5QTbXLiQfQBsKrOGVkLA
DMFufdbIhUo10Ika3cwPAvHBOtZQIuXQ/KJ49DN2i2HJGZeQl4m45tLKfhAy
agCOvM04u3pA0bYFTx8tXCp/Oz3dsPX7ERNuwADxDLsZOIZX0jVuBA/3V22d
vvk0lTa46PSAjz9CEeayn2JgRdKtTpb5xt5uvdBGiSNQOH6EBpssmaRJ6ubm
U0VWzZoxaNjYsp/3yNukzjL4tdouA+T5oemCZABSATNqHBJglFObY998GAe7
yLNex2mzLDPODeu7S6CqMgw6DiDlFgpVIFCUQIJWTKsXpLuAXvLMQ5dsPU56
iWioq8zwpiXJBY+goV0cI58YPyHqdWjl2feub0elXbJGzVa6CTMekkoQaIUB
rzJJZOQKtzBQRc17Zbyq4FXHs7HK5Xms1ZmdTkwnvRu/ejQ5PzMaitybktck
HZcmB4bvBm0JpNCNpc1dHM8OC2gPa+jyG5OC4LQ/uCA3OLybPLXuX4XbFgqf
1OAVsbAdKmsti9pmnRRskWrmM9GUTGZxT6AVe6yVbVL22OTel15A4cQTrxHv
KtiVq8W26tP680qfH3FEBxOJMrQ4Wngtq1DdT89uos712oAotWRGgDeapONa
98R8ztq2/hSFp6zQYmWlxDW8zGtgedOYi0SEAYR/5cWVuy9FN58R4mRP9DTn
lJQwmU9zw3NaUchgIXWBgxEuO2BPLaDUCNk3NRNBaMAzQjG2KvXEFbN6ZzYH
Uy6965lnGhrsCL+sxuhjjLhqUnOVhtr+xRGve8L4IrytBrM4omKktb8w+ysL
ekg3p9dYvEl+iwGfzh74KxgIjie/kGahpKMtwP0eMc5eoo4pUv4LRmb7mzgl
OcCnSlRHSa6nS8+N9Ci8EHGfkWbiP+VmuU6fpWerFaT5O+1YMJtFEZj9Kabf
R/UWHymiuNFzIq2FzLI8bqmejk+87n68z7Kw07kjLyHd/Qbh08u8IFvPG7Gj
YyyWtikD7nuRkOiI428RzMIQSF0xQxrwUV7hboMBSMMSGe3yT5ykX7bEAg39
pIu256QKk/zoIyz1AdaYIBAkTHb7ZnElhAkS+tMjI0nxVEnuAS/8XvT/WOkd
I0S7MqfcEXFWXUt4Cl/WjunD8Gm0UIrRrmEn9j+3UsvlRJlQhDk27TKUrv2T
cNNTEWe4wgf5KEu8f2rOl1PBFcRchos3T6IlMFfrQpWYYCvTUqSvWivGB/ER
AgZiq0k8jLSXdFjC1WMq6WhDTWToO2r77Pn8I5IPvUv7cpRbDtdzVHpXwW66
tkdwZr8At7utxAzgCgMmq7qofDb5MXsd+82XDvLyGtKmOlCpXRd/AjekinOT
wPZqniKQN3yV74nRxwDc/Q0M1NiPbN10KTfgyU13GFp1C97yBeuvKB/JmY2b
OthL7J5X0M3AaX6Pf9uB0UOEDfGGJcjD9Q3TDoEd0Yc56c2KAP9i3/pHcpVN
gL5XpFhxdDb/8k3BQjv8bNrhBBdLLRHJd0kcCdMKn2oJui/bMTUTBBr7M1bF
/EOaaQfbwW1gXGuFtqOTZNviqab0RtkRjqjem1Uh8nJJ+aGZTIkJRo3GbaGJ
n1DNP8Cwt0uws7nJGv3cDCnujQ2/RE462uXvBPMk8GexsQC221CNpzKhhf5J
47sDbB+sSQ1A5DduYwgCyjguGJ5ULXtbddYIvUmiyXN0lz9su2C0vCt247uj
JAh9FqlnrrrAEBlG2v5Wn+WR2hDHFiPFESipI3P68WzYJp3T9pN7h0WYz4q/
tC6pcg/QISIkGDpI7ue/f0yzZQe5YrR0w2avF2XJf73R1VO4HSX0KfIBlHjc
JuZMA3G6lAPZoi6pmXZwwYOAThOOX7wbOMOumFIw5q/HmbILRUbkC5G896GU
FaZfjJNP8EWRGbMpFf9l1woelpGkLIbaMuSzu8ZCDqQKwFvwMweigzUFJByh
sgEI11tjhzwNN3MUUsCLRYkp3fcinFurfJQLhOZENi8XYenbae9OmB9poJUt
qD0dFAmRzQJiUHVoo37mAJEM5h1Iw5N6VvgM2RwYzgb+dwHxXFr6Kke4hvCj
CAr+R42sp2AzzUXd19fsv0C2CIHoA7/PVbal1T2sg4JABW69jlH+7HKJkLG6
q/uAodp69xHkF+gppPVMBeQLF2/7MstOMssaSWJyiJvQeIblISH/C1jVb9D+
ipaWt03i5vt+oFHxFV5CiU+9HMzcc90SCcyYZWPLwK7wyZMUc5gpjLWMIB5X
24VD/QAERzGD8e0VWzm4XTPRrAG3nglhhCk9aBF38VxkveEhn1Skhm91plNu
qKvplXXAVfdl/33vHuPN69raNZ0WNlGTbmNc+Hajaq1v9kJNPaZGKfyU90wE
EP5GQPhHStrtbc+fKrNuMSOZ7qgRyPgJ/5xoUvWOC5XHYUYCUOfnYU4/TJEl
yEPm/qUdCEZfiF2fEwmrFkSfKn7CtmLx8wi5W03bQZmHeVeI4U94Wkk6G/Y5
1PPV8lY4ZeipRz5zj2rT6vXVHHldjh/m4570FHM+0sWrJ43wFbQP8f28Ut0V
MgVs8mKKOWCOTml0k39QAu01HUZ5ky2HO3fLmVUoC2Y4yrgd79pV8oqgE7gm
KFltKG/yuJkdJx0iGtBSrNVFMSNdBNHaB3Kjcuk0pI0wuNAZAcQpihvbJhjU
FFnlihe/6x/BD+KfzwqTHRLZHAQLu2BEu6d386Um9Qn+xdmUoepZ2DpOVYW0
eUaZeU6Ou8ZlW5khyUy1t94FhivIVEJsBhEl6kzXwDCaFrh0EEld4EpFJJeh
B+lDcw5XfqUXkIgmzVHaifurUUsiRnaPuu1uwuzOE1qilDr2Mekd55n50PfA
P3Ejlnsy6A3elFFduY8ItaRp98OBCloZb12Y2DsDKmK02yMdf8GAnDtv7cST
SW+gXIWJpS0rdjBNVEZIktRXSa9p19YdQ2irxqXnwEC1dxLae8Al+kLvS0/Y
oaGBIkQJVx8cgt5+2CCV8vkG1I0wFsfsO9Mi0aOUxrgAy2DRFByPeAZzuWx8
1Gww9j/DyIv8vlb4kILuk9/LyOrS+wB8h884VG3BJJs/3X1bGxMv6lzBSt9e
UCTZYAmHU2XjsL+9i1bNjAIDUlZwCV6DvsrvRLHFuRJcIR7ekHKIuIFULKB5
2sFdtPVgd/lIbEdj3BGHXQMvAzXlGtvh8TDX647Xs4hQJD0DA5/VdJNsmX3B
DdbUG5HjF92fSAiW3kcubctE2Tjz9HWTrZEixDPOtuaumJwRq8DEkBfdwPyK
IIiAX9vII5Wd93N0KpYaCVtir5mA5QP0aqpmxsJHhW0ZmM7kmeRIYr4KphQm
5OLsRsbBqDJ/gJ1b5jMvsW//LOzggcap87qEVooJCthxcYWllvjr6GCvc2+P
kT5LxyHAbR57uSwYJeSIHIh//Yyw5Ek1RQVRkJXiaOy+0RYcKQk1OgQXnNTz
56Yp6POPZwF2rgDb65IFuExyNUYYjzbTMLd27nWZkdYDd+UyuesBLgIC2dla
mEM38f8Aaw+4PWLry0fcznavLkSK8bNtyPDnV6LmdsCwCxAw/Z1MOn1P3J3M
1/sjddBfeevzui2TBqdYPIn/ZFCNYKpYawVgjBVdp6UW4n8sxQh1ziA5ij12
Z4ibvA3WV1KCdZH/ZZ4R6ZO8Zf8KFfh2iXZxwnpkP7EGrjErHZfDyXeUhG0W
PH1lRXWd35S+feIFg6ctierDL/HHd9z8p/MrFMzVF5UD7NqfsIgvD9ylj6O8
LWRbFHRN01IEP4082O8FQTyZfwJjDv4tPVogOA1yaoDJVuNTWv0x9tB5f7Dt
bhnsirKo1wAwJUEmqhA38XVLS5ZbZ6FrUQsQHjhWQ+r4yQbjhDSbKUKLLR+3
KE3z1M4OjIsG0LEtFr3sLNF61fvoHfcDk4DtoA2ybfXGUjhLJUVsulcaOquO
+ZtWNecjWN8q13RleuYLbUQ8wigzb87y6vvTvaGXvjfQ57VRE6BeOPSVx0S7
Pf06MSPOSmfjrm67ScxnVBtOrme5rFF8tCdktq/z5ewKNC1UxOmpzcpHEFeA
iUQWzONTTw4e+qvnpMkNtNoR4/h5dqg4RxJbYY6TlRW9RIrRmXSAUzOWLt/U
krS8VErLJhwIWX+b4wJ3oGSmxyb7iajZdXnj+v4p9cPQUxXngZea69JCJjKq
SCYChqqbMPVkpUd4ZlOO2C7pNNm4LCNIhLQPGYQLrtOVhtTaHah0dlK1GVYm
7GBF/3sSL4aIp39G5pIrPHMYJGNSlVSpOrXYPvY5TiQ5Wf+5GpiK7NRRK9oS
OGSqdHN5MATj2upXskd4S9UFeNghd8Xjf03c/xAqnGvRTMupeZXjdlxo23nn
dd2/pL08GKdiKWsjlA1eZAL1UuRv7aD6y98DG/gGKNAEW7nrAlFCwGsTMnk2
z89WHkcLuVLKwCAIlp+xGcw/8kvl2k9d2ByiU44ixbPRXRYzIjcLOzqLd8O0
tv83dzL9KVUbz64VauTkOe17Fnm6b2Ns1MF+l1lXPUp3SJJ64Zg+ktiXfEWu
iMFBopj2xElJBrsFzt582SsLbk7L7wC4D7NMYyN/hcM8URI1Oe9XCh7GMCTG
7xxjRXykSoYDyRQ8Qe+YxBGf7CRQpGLk2UPq1hvdhyrdIhdQ88lfxiI4qMZi
JTh8Uih1kXDZKzdTeTbOhDvpNIAmKCdjq4v2vI6/qvS2TWjGqNYsnDGJVBzb
AO6q1MLkXIDmamLU/x6hPHTUgWL6EeoGL6OuaLPEIh9/ETAh8fW7+5ko9ydE
uOq7UJnEFNsF+zdjw1MVNu3FNVoO9EaUkOswUnFPrd2tdWJQS6oT18rJDlPW
zUnHDncb+YGCxzmdYPv9rVUREIVI9h+yIntGyckmddbnnksFwWhm33HA4J+c
2PxwWPX8I3e6vuukSccUlJJoQSuu8mZcZAPrS4CVS7QzVg0gMfxt2Y1nm85A
QnJl8yh1KTUCgdo/nlFziSCtRRbPDxgybDIx06BcrUX65g18Le5KOxbiFp7Z
VOCjSdx4d+bqAole4+d2TFHVkvyhXQNh5KNQRHQwPZl9NpDK/QhveLoC4tyU
+rLy93xAE/UjVTef4sL3zDL0ENiWy7orXPZf3+VYb+vSiY1gHReNdJwXaYlc
6lLkzCQy85vZbraACvvkU988VR3Rn/CsQq6TQuAcs+h68ndsygpnmyr4QFzv
Eh6DzwAYdgUrYKa4IhUu3R7O1zjV0PmK73j4f1Nd7EzSMyOs9vLyyf6f1axt
dFI5ooAX8nhUDwZghV7vQ8arlSYyFpiaKIxBZ5b8DCHkXxrocoV7MFSzu4jt
9MLCvb4c0Er8da1vePIWF6vTQoDg4QL0Ucz4EhsIIpE+cW6TPPVvhYKJTlCH
sJuQ7OhxF9euevrABDWP/Cr7kf+mvVPTD/p1MHlQU9ds1gZpS32l49/zw5cj
lJdbXsGYVsxbJ0GEL50jXN6U01lWpMo4ShOZ5pMzLhvh+hiFHdoPd+ut7Sra
xDuw2MLybeJ2G2VflH8YZfyDoptI8p0jPY0jnuziFbbnndkws/XkLxI242PG
xz+j0HqnSKN+47UoprcFRqDD6TLk95cJg3BvaRtKXUPAhnhMNoIDiE7qndtq
ox8H/zPBdhlafat+YCbl442EJ903GNJSblrj8XS6HJe8LUWVFAd+CIziW8l3
bixclTFLeOp9rFbdEmw4h3gAKWcm4NFvcUedCozTeezh+v3oYlSxjeZQxh1u
LK/DtDandX6D7L/wHd+Q2jVD3jOlXSxmh0ZYEQC81PVurjvwmgX5DzYIObej
uVFCLI8BmLBv1UuJiGsFDvdoAUfLkv1+nABf1LUKV0XFWdXBikAOYlLCBpXo
HXpXL7MTqMh30Yvt9DeR32C+xjcROsa+sUweH4YFSbyb86dKjOmb3upMB8uH
cdKRTonYnTVyK3bgIBcfnkzhX7BRGs+lrnHQi22v3aHrFrtRz47ITYk8saYK
qehc2h9Xn8JbuGza9SAL1RnuHbGtL3sNBl/HP0aguqEkU9oiKVgINum0ucKR
YOfpSCpiilqURkkttlH99/XLJCFbQWDnTXS6S6h2N0e/3AUP3vHq31N7Shc7
QGzUnOouJh0tK02vJ9H0L8xX1atsbo1jSErdjCpTCMna6CbmI3m/5XEiMg3y
4D8eJ2AdHGnfP6DaKJ05OgMei2EKRH7KX3hL4hceyo++/2ytp3Z8niLTUQKh
AuHia05mdomGhB/20IwODLkYIens3zAeFyCvJFUQsR2sJnmt8hB1ZFtKJV9u
a/ueAbMKfNREK5UeDX2vBE7pH7PCrWJU+NUfbILe79FW8CDyIxhRRWwhOkCu
Vh6x15CFOiQ3tWnS9pmb7iu0FM5MeJr3kMCkpRwfXKG3jJl9sXGD2UE4m+91
KnIZtRKhqw1URwb+w31Ow4HwsB+XYZ6D7NZQNixpCMn/Of3Nw2rj8tql0tiL
gvgUBqyk5PRdfLgr68WyVISPmDaeLiqciqR223+sL/HhiNwMfPqNSxl9AmW+
zdexOIvoQGRntbr2DqTp9opxiu+chSO9gtGMeWwez1LyUeqJdjEFftpDreYo
6Vs7v6yq6DGVf17Gar+sZuXAC968PRxAFoXGrxyBEqgix0qY/oXJUK4ZAZwj
G43S0f16aoFNSoGvT3v1JgnAWLMSF9pfrwhWBttmyxtOQpa3xV8LAgLcQpvO
hN2dcWdnPGfIlDseqUZgfQdVVRkxeNJFUsIngKK2Wwgm7ikIPZJfIAy1sWGg
e+iVUlZdvthUDWbvw4yj58+SlodPzvuzz7h4KRcN+0J7ctI91m8GXkJ78EJu
NXBTG8QCLTfGzVCm3zzmONQbCqViYutAjO0TMvIkgr7rLYCOPJN0Eo8GEqX5
n6pUUayKGSx4rJ7ANaAA+D00fJr14JYKlMYuxrlzOoLuX7tE3PTwDz4jtQRx
ZMQr50487XQs7w2flI+eoOSqZaQ0shuwG2iW2HqYq0Tey1r8JoiErDP8mPxa
KsENsvDzXsFD6YbHIOEnPuCRN/Jg477pQ2YXX8dKuaFcC7zqKrptEajMEx3c
DJW+PkkbVd2dYKPd7kBE93FAItgsvnUYBu/fGii/AC+vspgT/NubmLNAZood
8QChuI2+HsTe/EWP0aKLTZC7rB/fYYzhbGOJZY78KIVOgZayJvybwhXqIn4x
8CgQRXTd2tPo70oyVSmnbsgr4i4p9OE/rUwLTCQtUFwLF3cNDhXsuevd5VwB
zIBOGh/pgTC6uNUEfaptgiRiSwPtvEWlSj2mQ4Apoi3e7SHl6FEE3FIIBRDy
64KMIc1UHG6k58kRcrOg6wnyVKwwkDUxDUYAArndcONE8h+KYnFySvysxKHz
GS4xhkJ3GvWMmeP5Z0XGMYp6uXmfH8jOA7Swk8KcCN4nqzdFzkGSOhrYG3Ok
F8vpBUUZEdhtAqW8YxhCnrhZ2Pg8lKQqjS6OLFhU5A4SzC0LwgKpg67Sjysc
4uDN3TGBRY/ryUNmOlhvVN5T7mHT1S6BgTcXGoZBvpTCHY+WXiH0nhNr4gRQ
rmOGsocUvjtWguWneBgtvgcKMfaivrKUtvVBDxYxVc9OZC9G0KO2n2EuhntS
CBIoPfBy8KyAeAfv+wOKm1+JEhkAjySLd2hACUuH1YWp4wRoARlg+KeI5fu0
XcuGwBIS2vF9pt1FrYnTHVzJfco6WjUsjEtswEEjOmuXLjpP4LaGOurmgVFc
9SMpmJETQkmF2qy+UDjb7gymAf3gL87mAAqGVbG0NhPvkwb0GPUlUaERAsFi
m8H4R5ty6F47sUxVkN/WXeLQKJz7nHrvfQdK74HoO3Y7CMP0wuwnucXWSEyE
pHfA1gkeCjvfr8bC7EW3rYMjJvH3Y9yGykHYhgMJwp2h2aVAI98R7yXAxbJB
D5zuyU6F9pHGmHkUKshnum6cJ4chWHmElhSnCJKQSSW3Drry+uaLtg9HeDWo
TZmmWa9vDW6nWnz5K933BE0wDPqc67Wl3qQtbB7XCDgfzLqPE1qvrOENOokY
m7DISZdtnH6IGMKQDfhaF6JrEjYFL0ijVPZhsrLzyIpZYnfqGoTpBIqnktH8
0aNjPYpdYmpNLW0KPFg/qCt9Sbawf9gRHr6esphyLTJ4pE7m2MT7AvXiKgDO
wG737+qkmGpfjE+U37JELWL5WbY8elik82utB2lddNfNSIP9p4jjj5Fn3qBk
2QROhQQk2bWHdfYs0xJlpnOWBOPerVevWGRRUhlbs0b2XAkOndaEpBYIMe87
bpUu5do5BwyVe20cGA/1XeQ2EIg043k+XhPIFOlPeuDUGHshLuvOI29p39Zw
fSJT3P1S1ynYOp65BNs9DXWPI2HZZ3IWL58IO5+6Idh+O3y5unI1EZfTULd+
7q6baxZ5PSTEOEt26evpj39KGVzwM+G635s4SyclNwRrzAActGdG5Zz7xQU6
eOutK9eBFBAkh/IIgC2q6YyFmeX97QLhjjbemC8iBzrHdq2Tgm2WAa/Zdrpp
JQPlTBkSCgImzjgUziWe/bIPSJ6q4W+0/Lk22+u9iyehYwMrGisQ+Jsebdwk
b7FOUasdQDWFMTRfP4OhKJtT9RmJiRrcifuBe7SL66haFtCOmrB7D8759jro
nwTQqLqlu37HzVUpZM2lwzE9bqJJWYB9RcrenHoIbfsEi4+dR7HVNraTQgfG
8XXeOxRbhKwP+ID348PBcOtMyKp/9pqtqpp+yf05wHcehFD/PAZcfGIbzS0M
j8sy23bowtqdMDafufbdMK28pYVA+CKDjqFZ7K8uXML9hk21H+/XEChEC5ot
0WO/89OqMQ0yEJxqm+Zig08lMZed0YUbsRC6lBdMum+K7d0nglQwNhdF8KZ+
UIiVZOwbjqkoqAxCVk7jbPKERG5H1d6jB32NKHzrB11dQU4/Eb+0DwxpH/Qe
CuvevEn//CzedTXFIcYraYcuWXiLCzDgUo4v4EsLE6/AfebFAMT92xrm1wXw
pgU8/SRM1fSL/U3VJJvJhLBM5dxIEnr5IjFf7V/wQRhRTeaAqYuJcME3GowR
m9XkRbCg3nxrfYGPYNcEmTesRfSXyj03qKhLxlJZ9bI5EdAWBCD6nR30Jq8d
cms9PSU5fKboFwr1n1Cc1Dl5+HzPuyyDXIZ5zmtYMT2UxguGuop4Vt1Klplr
z4DaFwevW4buQ0dvQRt2ifFN2u2Q7GKepTMTP8xmnIYh/st0kw6VErU32g6D
V8iv+B96WfkZNCmpWr+FunXQq3uaPy7G/Zkb2zFwiebzm5NRHWbv2oanNfCi
mB9MsHGJBmPok3bUiq8/oouh9crlpapcHsJC6EBJXI3SSkT1rFhizrk9Ef/k
S4qaa8mY+b8X1kUbNdkT+qemFJzGOIVVHSK+n/+FzkgqbHOdc7NVLBzO1MPd
ownRZLeiFVXsE55S7yrCUzsiu/dtJk2y+QPbWDdKXYCsUSoUxR/NTnAkmNnb
CDTcmKKVl/LHl8mn+beQQa/YfHOKtRYWZc4jCFWUmjMC654bXtJikDwIibWR
MqK2fNfRRWXjBFMwH17L41WISsA7jf8ZbocEl1+1qgBana83ynoK/GArcuwx
Of/EMiiukCb/zqaP4oTL43pdqg9R+ROe6HZpz5lHjgpupr0yihnOsh6uywi2
C8xNItgpKgOOv4OjpAOB7qkXM/l/zCYzEqkuqNDR8nNprk8Wg7cfvYgvA5Am
eJQZ5RQnCAT2++D79wa1Gu2cv6RSW7mp8abVzwY1pMFOONUNrfUBlMj7xG+X
2VLn92ypYS724L0ChSx+nqjssTb0WRulssXYTDPedBEtz9imV7ib8F5N0Qix
i+Kcir1e+0bvIcNj4IsvjaRi+POh5BWXTL7ylVKtElENRmQFEqkWH74LeVUR
8a+eJC2wQZGaq9p6LSaIJdwFwJFOj4zQxqhfJO7+tFTJbXEcQU+dtmuzP09H
FNK8x8zkPdK64t8nwDUIyF4QIkklvgldvw0qPz+kg/8jPfYwJJz5iTZ6nWmA
gHvpnH38DeeI8tiUwtastOfX+7kdbAEsejX4j0YiQpYw7J1VSsfPj0dhajWw
/2MHc0Zwuav++VhhLeLICpFp86t/xRceClj2BlUUW1nyLwHs4uCrl8+hERTt
eYynYs421YK8YiDbEPglUKrIZFQreHzkRxlvZUkECznvDa+1AkjLcuqxAxQk
+rOn2USHkICAhOfRgLrRFFg2EbKy7K1s89uF8menTCBCR58+JP6s3bnGriOJ
6SGxD18CDOXR6k6/t0NGC79m9rh0hIUGCfQSj/QQNxIdZbhRXTE4nrkuVP0Q
5McivrMzO5eUCdhox7WtAuM4rP9FFIoQCvKv7TjTYwL4MsYjUGZfcnv9b20b
J/g7oUAbTLa9w5CKwceIU4Qu50gDimdLWvefiwGe1MRZ9R3EO8hEwDwXrSdN
V082aGTHrDepFJn0Jqoh624/9PRUPzVNzGeGWJCvZm4YKx+ideqIvbOm/vVI
T68WKblIbCzhT5tbv8Jll9SB1naGNcEhj0pyIW0KdKZhRge4bQLpRnnJw80l
id8mIyicRQR1QDbXlkSmDdt3iCk2NcXt6u/D6yj8SsjygmJGLPeNx97BMN/U
N0CYPcHCzFiCPmk291f9eMgGwydK+F6UaAyRmNd/L4xR7636KMPfuzOlKs92
BOPilvfmjp12G+SGx5nsZTKdONlgqI86notsL30T//BWhbSN4p6YYB7GUONE
mPDXSBIVNwV+MhrRG/nC+PVYn3cR5UXVvUO0NGM7J2jtPJgML0TWYhBL+Xox
9QIyH4ctMBQUWReJZxdn8n6og6DUGRwhA2+2g0JCKWHfx00mgEuPRIalnIXC
i0DkJ5aOF+jdk0p9SXJXCD9kocsYjmyAFEYdDTmsl+hoIpNygQPofrQ3Jc+I
TzQLHO9XBOkZ2Ae6RuVwXmOVjfmuwkWBhGIOTd/bphXA0W5Sb1lFm186bWkY
9SNVa3xF4o1Tre2jeFoh3kLaw90AnpGNo/u9gp7nJhXto/qmJWPNYRAb0yt2
V2lDehLD3z/kW+ylkKdR3CKxWO7wu9To3rJYuklny/PjmAd8MTeO9E7R6o2a
w06Zao13aHBspPcgO5QuIps6qa/gE5/VsEGPtWDE3suvdgeJag2FPloPfgog
7T+k9cQohr33xEJbFu8jn9TH3QSehrLEAots5kzHwS0qooK2j+6in1kDxrKh
9U5O7wr6WJk1d9JLsnScAofSyk2JSla7QplhRjSyave/BnvbUQJReYmoPCie
DAs9RbOP0+ifV0HddERru6xUqmCDFy8BK79hDs3yWa91Rn2KvaupbyOy8BbX
DC7+fzzXIaWl7WGf9Yz1C/vgaaMN3cwHDrA2XkpjlseCgqrdFlf6Ab5ylNE7
kAsBtRKyClnaw0EpXSB9RXDZi6isku7GfHcw0Or82zYJ6bhlCFbONVXxKDS2
mcyaNMWOL39seU97pTSyq+noc8Pm9O2fFMCU4O1gDcu0rOqIUKRJOuxz0frp
LBGtRdEbqr6lca4T+Mb0ay+5l0GbLqnGuC667x+4rg4xTs+oLBMVkGS8ekrp
b2H7avP+FWzkiF2CUd5FoClNFTd0kctU+4XLmEiGfgUiy3zifiUvAEP/gFXk
bZO6JvG77jsxJldPUThTQFXK2EjO4lBNWrM4K31ZkrKSusyNXKlqnUk+2Zyy
E3oM1zERF3NN4l/iYnonUUP47L1Etb+bgTCpp/R6N9haKPLPDzcMoilD1ggW
5L7Ai9IV9F3xgrE3If7ImC82gpF1QLQOlBHyByEMnDQ5Mk4uzkQ31siOva+Z
TWBq11rApqTukrXPi7UcGBfGxKR4l6bxyahHFjP3V47ygRaNC9bNx+Q7399Q
ne48R5/inltzn9PCsEEKB7G9+AVig8T0NMIp+7Vdzi2jJKutzh3thVD1FRfp
cY92mIVufj9dIjTd6J+QDhi08Y+wefD6IOCmdf4V0t2a5/XAsB4jupTxJecQ
OW/Y2Df2NDIizuQdLhcWUG2eEgjt9ZsG8wvHcU6VbkVE9h6M2RQ3VlY1PZ0e
Gwd8ehyLGP73jSj9XRKDI/AkQC3x2BBe2JyG6BQc8zapcwNPOMtVu3VXpTZP
4HWVju0GBpbd97mJbCWTzQaA4+jdITa1FIfWSaXR1qvOPrMUV6INpvfL/tHt
QQCdSobXp4eMW3Ln2xVmGZWOgEdmn83Ou4/dmd6MoCvu60ZssVGu9dp6vPcU
Zv/fsjrbUw9QtWiSoa07ZRrQm4ZVbHmENW/j6bTL6kPcFYXU8mMVy7W8ye1+
JgTUUU7CzrPLmx8HW8kAVvI06+vwOXN4wzbZs8aV3utuGjmcKpyJaRw7Krku
KIsTOSbaFSW8GRlvGC3B7dGFssailiDRIPfBz+yMONtu4pEfGVqj1YhCRIGx
EuYfzMISBr8FfRKFC3jmHKbuoliW/My8rduNBn0YC+gEZW0eAjiWvV4zY6LM
qDgy9QkWvnHAwcv0xWW8gMb+HqUhvlWOOlbTU4A/cCCAViSwyTL6sHv/c86t
JWqsl89tqxCjTl4ETUiYtMOirxVxTSgEcqF4XjyOeD/fDwNGNXdeMWTzXGcX
4SscOircKZGj6gqTm/HQfVd98qHzV6qDE6w4miJuXqquILt6t9My8oq5VYlU
qsuVaCy3FdO1VLHUfdj7iEwa+QEhkwVv7urPiddKv8Ij85jC9YKCUdGlKQzt
+UBSCtrybLlefY7ZB5OwU+uU9G1zdSsKH4U8BxHZfZVQBErliJSg9zgb9xmL
cYVlXAfgx8AyD1/Bdcql3JbVyr4C7JHcxak1+kgE2YmHNV4sV+FYFvb/SdOr
oncLRUp9bE2fKOi6LPvEdloFGCnX0ztD38mUhhVQUgGV5J4Nm5QwnfAIwxSr

`pragma protect end_protected
