// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DMf7EUyCBngCK+hixsBe9p1C6vZhKgs4/zwiOeU74jN0ris58NZ2jKPZ5i/D
Ho3/yc/wPVL+L42eJVpfSSd1ce1H4jBU7xx6amRiZg3O2XLoj6312UfA7kmy
8sIVZCctNaAUuJ8wm1O/9ir36saO4zQhzcHElvN96IukKmkSfA31C5136sqb
M+4FYpD5Og8DpUjyzbQxRuDNyuiRLHFWriGzP6NCg4MnPr/T8V+7AKFIuWPL
8ixL9Qv4ftZL3kFG0J3WkvOaaxUvxx9mFHnRaR0ft8aBGQohHoHcwul19eVm
+arAaqTUBFmxvHcE/fQPUq0iO1iej7P7aWlc1typlw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o/vX7UIs4dDJSnh2t77N79Mzj1+a9Oim0SJPqcbfRxsU3m1yupBvQSosw4cV
NdPw6bqThMCH6mCMA4reGFgsKuPKz6DSx5ulCDRgmaCq4CGH9IiQNVGuLMNK
+suH0NDkNrTCRmzwxr9H1YfzCBZDMzAI/CBfFXWdbBP3IusOZmE/8qzMHOxi
iNbxjiLfwgdCtZCmMc0r1r652g9MQITrb04hA5z1sUxSXF/J80+fdHb9NvcI
BaP9B7pW60iJPlk1S3WYHH78EthRVP6RHHrb+Qi2PdJWGLJzdI+AD6NoWGQ2
/RQf3uSvMmI8u6nm1jD3Pbh5+EIDdo5nLQGFINK/5Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gxz6F03eJsSzYw0eJEakkSDATcLdnODiuUzSV7EqAewSmUFZyJI8qotIoxdP
vwPbMDyG/550rtOimGbG/B1Pgglp5orVCtD52xlMJdlQ5vr9f9grKoS1j+7K
fgV94YyUiNe4ZL6N4vfJLEPjbDCOUra9crJDh8s7FI+Z2Yd1lN7E9jLbVe3T
1qPgOPplUE/k4dkODJ40+s5n9tLN4qtfTLWhl/LQnwnVthZY+s9eJZWinujz
ObNm39jDvR0dr0ZT6kAxeYXVH9tSdvTX1RZ2vuysp/yrfDrKpR2gCQJ7ts9B
rurFLBnHauzfEIACLnMLAXI3bqh05XouGqCn9SrGAg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
es4W5MyILZRJpbOnieK3hbSB9eScDfdpc38wqrcDeufkfze3/Gog5SnUxjBX
qZTfxPHyBwY3NbwwiawARg+rXYquLHe80ElmrnUnrkRPR1APMHUAdTnbMJb2
H8wDOvys+JCMA4shG9uVL6uk8jxEWI9pgNSi/aGnQqUUcOFbWo8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ra0Qvq2yo420xwzBOaOjIhttGJAZneCdIAiSatOZwgBUNsm9yHp3vQ7tTbJt
CtHN0oXKCUoZZHLzI+4dpTaji0KEZG6t5B5NGs6q0gv82hURShewilbb+7Kq
rFtO2QQvcQIlmotp4B8SnXzGNM8Mdj/Yr972hnnimQICUtt82TcdnQUxzxej
qcrVeSQuvlGxvFVcgR27LhCL1afE8a0FRwPSUsDcokX/S5/GqAVel53Zo/+G
SD+Ngzb5O88L93XnyV/Hbcxoj5LRIYj8R8NFj5EUCVLjey9gO9eOeEIcG0Yg
PPngDMy2WU3DY/3r+POMOHTMN9zXSr3Mm4W4C2/GNmqh6DHhOqYaEyvIsTYN
QKKNHll/LAS1X0c1V8UckKMefMj7RThQxayKBAJ1VqGrCv+cTKk15BTg5WzA
bgD1fAE6CVHs51HqFF+tJmRDd26FwNzBg+bBtKEQAWm4L8qqGiwldYxWYcjW
oH3ac9budZb1d5yVj33dFoJ9WxDeJYWu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aiIt4ALy1aB22IbLoBtazsPN8yNRippHtc+ebTNCC8ioBj3OclXYiiHMO3Pp
2OA8FpCRbgD8XUUhRvEKKwC/I6gOPlwCHAXGtH9u5ynvxkcoyUaF0Hcu+zGm
ExadhNHOiAtQ2jwtYOXJV2/zvg9j07K1DdXkO7MVdKPGzvGUY60=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ncqs3Y0JuJit9JKNniJVPh2cMB2L3bWg7JAgpLmKVDpANsMqeizbtSoCwmG4
6CeTbrLiiHjEKXsR4+uhE+jj6o5ADaPa+763O9XHRPfNLnTsfVQ1VkRFJt8w
rks2Z4G+C+Fz1D2FrmzjIsCbRQrvMG7zhWfEfvhTYOCzUN9zJSg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9472)
`pragma protect data_block
0N1QMORMwL/WC8O40AjbDh4tthuoJdq2yaJMwuwCB6JxqD3VnjMjmYzDK1nB
yuHIMhhyL283IrLpqpGsvAY2hOxbCdZpuEvQXr6sqVnSzJWuOD4pH4zw5Yfu
o6UvavRUUlGc06kOr+CydPEHYhLZ+2ICDwn8OeJg1QmRVoXBl5CCIlMpRByj
+gXnmebAIRshtKPQdnRtevVZucX8Iq2X3FED20Phizlnc3t6Mrvpmcx4U4OF
YLiZoJcp/mVFsJX7DCP/1yotZQD6vpyI3RmScs/Gh0U5J52AX0L1sriN/Fkg
rDGIvDpcXHlkKg0e617nXX/BsjR8RQskW/UM2EEpC/eg3js/InRYhfGm6Vda
bQ3V+ezTmP5LERTqgyGbqOcVF946Y0xAdITiD8Yv0AEyzUzbK7d7PD/fW9lP
IXB4FvIto1CHKcH3e4NRu/HqZpdB3pMVdV8xveUhxD23LcEzlMM90L/8yixc
uqUVYwR5U6Rn4WvqYo8zb8qmjUzVcBWvWVHndA22lULyht4ttDbmR7lMIx7G
x1ClRzKx9Frbr9xmoYxbKv1xH298NaVv+yBUwAIch0NWcULK/yQFHplfQZZS
25UjK32C2uenfKRgBz0P1oHbwzk/InWYqtyKU+jfDgZ2C1SVgYE4DpEnFl2q
BOyObUjwWm8rhtIkbzlJ+o5Xy+4kEhQ1+9jMcIUGkVuQ/n2X6VDfPIWhcoSG
09uADHdlavF5qLF/Gi1ZOUFI5UsHFwtVuCJlqtf1GPbadNlr4hCAaad5e2xy
VqFzX7mnZqDKjtslzI0As7cabNH+ryq3kzs19U4WgsT7tOoFsPeEU58VP+8X
WWuSuO5372TWu+gtcCJWJCkgLbmo94lVag6o4IGt15V5SQIqeBR/jRVEl5bw
eNczQAyDM3jXzDBmkDF9H15l6eRZuR8OovejJyfpFLFbG1lKGloUgRg8OGFZ
LEGabyFqoMA3IDFzVZqPssig8hZ7kUS/TBMLEaD+Q52S95eJKBkVQEp3Mtqt
VK2SoSWgU9tYOnZoZA5LN0BRHDgVLU5jq/165UwnprbGnI2/Euyfy/Jy0GwA
S0kQNss4idtqUxB6uQ874+qMKGU68sgWZx5bU/bow8om7LGx7YuHLPmmDLfA
0NbUSBCui3CiDm/lzZfBn8phWmRhZM/G8djFolaH76CisWNvovRtAekAqS2J
xafh8q7VPXld2EDUGzRom5Ad1YYQsUfh0iDJYppU5VL/0oEFoHPSsW9zdBbm
YY8ld+n6AyIVWOG1RyKfAI25duwcpUtK6Q/VZqhs2IlEIN+qHUYijD70iBsO
ern6e8fR3+LvnGOpk3k/mCsaW3O7RAfpYoPRyleTKoAvDcxv8pgc6Cf7fFhZ
cSm7rKYCzB7jgCDNs0zYXMPbUERoMhFbRjDjtLEsI4csAVLsWoQTfs+xb18h
w7bfryxUruQx4pijuIbt7dO7LP25gCeQ+CXci1e1osqMnwN4wuylb88tg01j
KKL2czZHgNl5j+EORgBWk3ccwwwEu/ROkFQuKabsQRUMhY5+0olqmalpf7Ri
zoJ995dDqazHVPn7yNSOB9FAg5QFZA9KG3XOaO7L91kCUb7g8t1Id8PFfRCm
DC4SBJxO+O3n13DWr6xNE+Mvko0UbL+4Bp3GkTaOBkGSS03UeV66R47mAftw
Lywph0R3W2KMcHacDavItycUnMlDKra61XMb5n9NtnXoovWFmjej9XwAapj0
nEBh/O5s9qdYS3zQtLnFaXIpaNC44jR56grWmHp6i5+nPt2lTkkKw6FBhPuF
oRSV1oCYDETTHV8qwEzm/a+l5rzGUy9X7iU/BC2UAddL69mP7MU3spb0gi9+
vuP/2PvK8xcnzQNo0AsvgytUerdobWLSQnsmUvjvJ526N4OKP7KbJ0zCfqaQ
DzeLX8QnxnJOgX5Yvt52aNNo+D+4d7XUB5CrVoaHXDsJsIwnX8HrPRB4KxK0
QGHll/fSgW9E6AjJbnU+HnLvOKwtXFHHqFDhTlVP7Wv1WYCA1/S1OJ018kFz
tDK/okaj0XJg6k7SfrmS70MAs8gpD/SZSaWlmuN5uJX2tFDSVAPWsjkiKnF+
Gf+ycJl8FmrkuS265YVRSWXeiSk5hPWx7Tcx2Y306QCXR+7MLUBZmLK4aSfL
K4jeghXx3BOoZT4U21OEaZCpEt0152CpQd7LVl+eqgk+IUupYepULNLlxzlk
5Y8hwwel3SXYW3zDVB6qRjU2hnEw6nudEiU3yOHhHnksNmge2U1rOOeisLVQ
y1delCsTuvYcWVEIUQPH6yi3UtYRxBTto7E2GJzko29Jw3OPbaN/QZipImvp
vVFvy0x8M+gNYnfyMpTTceKqm2T0Y4cQMFg8yRX4cEx2b+ler4FZ+AyPYp29
1f+xW9X36Pky5SWDUbQa6pGiBAjmnmOYZaTmP1tYZFnsd++vsSqa5JMPbbW0
FEAQSDCnllKbq8NTbF4Pf+LjXO7DvnbkfXLeaOXZqewesB2IKjra+EjuOUwQ
c2J8Kqyi94zQVeYBJKKmMwoGngYE6irUqhES4N4QOF4RAKNqDN/Lbmy8gzp8
9WdxZHtCLrbd1KoOXSaFyaq6LRKWClMJLCMjQbIn5EwsDdcKypeUFQ6+raas
JyjMasij2GwBLrZL0AGuWdbH79JP0TrFCioO8BYyfVU2ttTAJNk7iJJOgyv+
vJR4CzwDWPINJ30Uv9jeqY3ApGhoS+XIIbfuY7o4GxThZ7ng8zTuQTMI5dPj
2oMYo8lO8yeZ7kvNsMivmT4FiE9XuA0bW6hEVm0n+snYi6cn34pDFIyD/Rk7
G9IA9rUysoUxPCytTAEKO8akFehR2wLwsY5sK0VMCVgnfBZVa77MBAVUIkYl
dJexvRugth9M5iwuQynB3JI4RCIQi21TgDMNag2oLOZCSqZ8IY26uXoCswhO
qG3lyjuAS9YN3SdIE0NI7P0BxRqnCidN6eLgHO40CkBU1WZIv2E1DSjCbmOJ
6cVWKR4cLL1sA3cz/QQLeROtxpXIh4ezDECxsYV93QyJL89A3TSrALqrt5cC
tIWfi70rqoUnU65x4RZ9xP8Ttqj1Vvc0T1ncLRgXnr+0gj1nL6fKx4skb70L
bJaQue+Dgmil8k9EWBtYq2yCatLeoJqrvU6cnmzYUxpdTX8xCQ5OhiB6YfPJ
rzv7rB/cvvcBWYHh8WU2LNbH6FCiGH1RnNeNKNMevxGKx0vMqcp6/JF2TrQA
5K48Zc6OofutpmyfH47grznGSBX5AMzadL3NU6G0uUvBXJZecjIotxVZpXi3
fhHI+M1y0WWOSD9cwyHvsR1076FeT7PusRX6yBuwP8aZWn+xg2eS4pwpjgr+
PyaJhW9XBSMkiDb3wVtSNltqczq9uapC1ujDikeOJBbZyy1eyJfrJVasY5lO
mQDQzW+j7NH0zMoEFFqwUdaT42ePLHibLEPO+gIEPj18ky+d+FBYFVkVOSV6
P78jnE8ZeAiXrwTDifxPyMYdULyGNmpBfNm4cReMmksKB+r3mkfUAO0DOJld
FFHDb/V/f+BU7g1RrEwGChpOFPCmQayhiSNsMYyc09cAZQseQ/7FOyXWvUbX
C4mCuxCDnoOP51kU811IUtnMxQVmPG1Rp3Bn0KJWlK8bK/FUm3gYI/7BRP3d
Z+QcInykhT3/57iPM/CHhPiTk5qwWEFAPxO24JssdHtgWwz7rXVYMUGilCdF
iEMuvFFBL9b+LB3YlUN8/wDpyj7NLvxG9dqury68T2jnnYMaOvj6i+yGBO9C
8NrDckEin6RsGLTlDkEcbaQzEZVNRh2/f5wgt1YOtALr/EZxRs8ZFyPdEBCB
mfrSuLFTsyyCBaWzrH0OA21p9jAVxtTgle0sjRIjHwoL1VeS7My+Dl3531HQ
Dxlt+iWPKr8ZBpp8OksbSgUSUjmV3JDW/gCL3dxALHzzbl+/4jkrEdNZAJUt
fUpLLfvc4mPeFsiw1VMml6wXQGKGEai+1IK62urxWPNtlEZxZW2l9PFSPmvX
xMR1rmADhaYCTBvHhQ82ZzWVkzS0fm3jMsrKhZQ4lWKWZLrWU5dhY54IKB53
KQzOd8Eo+eJY0lXt6qT1hc1TAtFoo7LFhONwGxO+a+tOBDgXb0iUTcBe/NbQ
U7U/44j0kzrvVboE1Kh0mmWgAGC552NwzIXl0QMgnx9XFdMAsTKN8a+cnVlr
1GVvqZh2ki3wSs22tHUEyyRksGcpu1Qs7b3wo10gpgoWCX5nsFrBgOy5M0/m
4fKdLa2Mn4q+WissPEJZ4w4miAjpOQAkysZLNUwHjE3ZwWraOQWMJAQB8LGi
1UZXkrJWgg3mzQUHvaPn/X0dzQZj8RmyeQqeuThLFccXGG+nFJrvA0BcKJDR
4rSdutpK01y6fQ85Mo7fUxyC2JRE/Uxrpyni0/HZaScxqAYtUmw+V5pKNdNP
aKgq00hI/pgzW+7GK7Y9gkssRbhZLw0L4VjBUSikhjle7y12ImNMnzpCdO9C
Lqh3xshAqOSrLHX+XtQC9brhx24p82WefVJx2OUAVVPsrDbZUurglzr9TXb5
6mYYkSFurBgNlIb1/vOIeBAhHUtHdm91oMSwIX+jji7L+F7TcTJgcefTz+SP
5HU2hqLRU8Iazl1LZ0NoQF4dJ2VOHLYBtrOrfL40YHL4UT/vgopVyMLAUp/Y
65YGIDy+5ooq1xfbcFli/gmXrYnK7E72/Vuxuw76ZgHJ1gg9tta01qsH7onp
z3DyjZcilGU8Au2+lb1tgQS4+nqS6xV4ey8MVdUGXG4lDlmlMfTxHNq6ekW7
Zxe8WUEkg2RdPE9mnlfNLQ9NlKv49k5KxftnxZN5mfvVBdQSpdk7T9ChPj7e
f1E+Uxndu8MT7QCQLSU3rniqtzBgo5ZbQVSuIsKypMuXmtNn0XMSn3Gz4ZVO
h5ICQ1q1Oa+bWmsqO+VRoZ9AJCQMbcWdEvQEyp6Fm71wM4EfLNIxnD8HZmC3
ziqAglmhj0WI2Yt4SNilX+A0DNMRVLhCPmnRNHds/zXxwMoXEfjSyUtM4tvk
WM4Y4jVCA0gt2/QiNKXOzbuqYDhdM0vlRveTu4RETcDUXFev++JkcfxZPhC1
tzQ5MlE1pOwnKyuNMsXLyBqBFFlhQ8cW/PU53XKe1curi7gIqWHMMdslaH1F
eUd32xupOkCRO28Rc6RG5xenoK0lJ/Sk+uqmaU7emqjqJcqgJxwgdjG7wrWk
Nzi7YqdzvHm6XwA4NDhezp48kGIm0U88gtcY3G+K0SX3O0eJnmoD+ucd4cL8
O1Ba5nise3WyWqx1JsRUvSajnc48KbcCDtk+uqGDegUbvGk+fh2Uy13LmH8e
nKB0cVFSyjuinhYKKG5zXYRkcTse1NvbGoiQjuoFfxWbUTgCHqEQsKny8Wru
9zSCCEGO85qNYxxt8JNzV9WGWAHJIHLkANBFEKLiZCx4Af2/vGlUM+YQaGt+
K3intWVVVrouWiilClodWSgUOstZTidD7H5PO1zpfAamt+lgVOWfzVLUd+I4
rfVZnCdbV5NTWUcXqIxydvUIVZdEvVuPH3mhNx0ACUPcAxZic5eFgBoC4Mfy
DWrJgCSXJsukvUfAUpqDPnaklqhX77+a18qtgRDZBffXUZA8us+3ajQ2b975
17NEC/RobNViqgeirHpofhxGoyWlv9PQHb+A9ATSvjGc5vK0ef8CfnhQQ8CA
q0FoAsQ0nTgr5lMDv2s+dkcmMmYKKvtXLUUmq4haR4hFhKxUYP68cvTdTaje
PlM1nwRhxStHKBHot5nIyCtfvdaUoRkIsYIsxNVXROcejIVDEWmsJF6bYhQe
e1jjmnGRUAeQccBnCxacT83feZ5zAr9LlmUlVAEkzGjsrWIFcrqAc96pMjUQ
dq7XSf5NvSn/tcvJGN/0wotXY3SAMmtF3BAkFPDEI+tXhyIcgS9zZRPbZu7j
HDzj+Pz47InbUOQ+tFgK2uJxDmveBuQxgLwrcIUcrLdlPIud+mEXAHfIIsNF
OREm9zkmSpQQUmk56XufbAjwVKCzCfKSb1LvLpN4kwvbArdHClHUXAIUjbG4
0d8NFWafqHlmHpdQ9EumgMVCQ8Bs10FYEAoAyl92UHE7+wb2LV5lkDNIoxR+
PxL2u+LqdcBDNSzbynQkx8P4JpJ3ZZFsERO1Vm8SjNucSpdq8fRDRG+a15Bz
/Hcr5BzCrdX8/mIlihFWUy4ZDVceSczeUGngwe+f2NZx+6MuxTd0w0ZwMQpj
D6qh4KsQt6d9hBD+FK9Y2xad2N+YOKjlEE7ZL8wCx4CC3upc2ZkK7deEv534
N11MIXCzbC3nrZqWYXS+EBvT7Kstqhwyh0KHBbYGMM/ODhVGjbRDKQLZKGm0
ONjz6Y+BbHyRBXyrh52aMNuI/eOYwOD/pIxj1MmSlF18TcQl0vhdz4DdeVz+
eWBtqSYy3tzifaachRe8R/W+PKnxVWeC/2RzEgmYf2kKhhRzGjnFdcWYPtbA
GVwOWG3hcGuNym9CI59fwfxyYr4XyxNF91xcEscETEuyzMpcjL01+I1Au7hB
8ysE+r7EH6punsOqoWc0XqfPQupQHWvZ9oRfjpWDNgjPrp9KioQ8QFHICRaL
r/tTfr4mBtz6Lv7QoxjR14zN99iO3wQQhHFSpdcdRREVkHnplVLq6WBNPaqK
JH05PpLjDNrr/FP4O1SOY7Z65wHJLUx1qknLMCdmyz/4ocRW2O8GJLh5sXxA
CrAI+HWi60RQs6o8LkWJIelMKrypwjCRjd7F65K4AqbPB8cBoH7Kf8e0AQH4
eaOg75Vymy971dVMmhrJ9iQK1b56SEOz82AlTNpxxAn+mV1hpHFL5caQpwNS
X86uN0eBA6MmlIudYepXSTBPZb05fCRYIptuxo/zDQO9FZerSN5b8mWeelhq
YVcrxqwhzYD5byPM9moJkaADzqdHRZFdf1hmFenqX68rakZgJZ1kRmYWRZ4y
GGLOtkP4hm5w3TcDchLalmLGZu4ekcoFogZI8+XI8rWGN3isnk1x5mUTaZr2
ltNrUxnXQYo+ki/mq5pEXVXoXZZrWTp449L6wF71a7zpenxcQ27OXfycEtXV
QxDPz8CeCRzLMzbaSqwj4G5Fx4DM3r8Lp1VwTlah5BZF/bxhb5ecl8Io77uN
nYHN7MfiASOtUqNe2NlfqB57rcY52BFIHGizatGojaGIhhNHPmvX2W3l2SGP
tFOHSii63+vczycVw4NvbiEMNfhH1hnEH7xZ+gZsxt5AijUaH8vWXiQpHlS8
nvctx3D/kYOU5CSLpYVMYLcSZOyQL0NtMdiV13Mmsmi+2NfDknTSC1+7D3E6
A6t79mmn7BzKfOY0Y//yfEGFsoAhrasYvH6wd8Nzl8vviv376jeeVe6I058W
pyfi9jFpawB/zb94X//zOl/QBRs9r7EcXmjC5ov00Xpxg4farQBbdCR67/am
3vvo9n/Vlg0av0ufGraNhn/DYmuUtBPU8Lc9VpYZ7JFfe8CBXR4Bm2R2kKmv
ONYiwDPTMUSCihOJ1f5QhgCX9BsGVbvlCZ0dasx92caDKuPs9Ha7nZfmtRgi
XpMq+dYPgAl63K9zH8Ks3h+2e2GNQaMUSmfeS9xagWKG5RAH9MtTNC9x8aOH
+f/VMvzUI4qphc0xJcZhvgc0bFdXdcEHbUycuiSQ3/F7qmr+r3iNK4BIiqgO
BLRco+s6ckzTWEO0IiONA3mpvE2YAA8KICRoZDN9Njudo1uJnNaZmkEjwgpu
rPVA6U2SpqN2FiZroW/Pa9+5l9Q5wAO9olqaIrH9VcUhXNk4He8QlLbULyRQ
Jl67TKGMG4vcynj5kD3e1par3JjtH8zhuzJzS6LMwIVHqLsIbpBtCmzIE76H
QtoURr2nL8xWbQvYfSOJe8o5gzwpgKVqdAj2sjuPe4qs8D1ThTUas8ppfQi7
4lrT0DeQ7ets4j5Ofm6HFC6NB8+YxF+IggvgQwACr7ijMGg5pR4qUy7ilWL9
tKuwTMhJhy0Qh48G40kbFPlZ/N8E/+mg+QN7KK3XNbuec8QEX2HtOSbHEVvL
4CU5tRb5LFZRPzQZRETDrlz9v/AsLAdHRudE+xm20DsTFr/DZlXtdaF8JdQv
kS/TEqBJ9TmdHt+Yj/Sq+th5yZA49are+VXRGUmd8450FwSQc6sSDKh+fs1K
RsUUYyOKR7KTi2yVBUP6oCkuTgi1SGSBkqUWBv7b0gzgY1BaCtgAJu4SrEI+
KpZrG8bgOZtz9aYH+duxVWgWHllEA/F3Dt91rnQTdEsc80zRuNLfASz32UhU
6M4JCaUuUXS5Vg1/qeQFqbwqdr2Qs5xVK0m4oQ6BZgzSOZr8+yX661j2iWHZ
a2P+SVSCOKuWhxFpr4IvzJsVnS0RC/6F+plIeR7ElGL1fK5nUMGINEB3ahJ4
/J4Aigm3iEht0k3aAhAvrB3WVrLJHUrpgUq3frIl3FnG5fTOZQwxfoOZ3fHj
ZoeE02XqmtAcvIPdSIctDWuors3P0r4Efx2/YLdZri10yYay6+d1u99QIuaG
6pXC75iBLsU/WXi4J890mvqcRC0VInOkPiDHGJdpDMp/NGVuH7yE1pt+GsZY
mTjTu9dSXl9HmKKf1w1ZI0nnXuboj5TYjib5euj7KPLf3N/QRN8dqOIOQaks
EdTiNJawh+XftYBR65xOsvTEL8afw+ditLDHmKyl7NFs6h4dykExcrPc8xvp
uwIzgQEWlN/SV4b182OU+Q4r3+xCmSOvmiPDbFA4lxGSOrq/JKzZTdFj+XNW
HsSfsCk8Tn0ozBoAwu4WzsaFh43YHZTO76gl14LBzt2IuBlIil8DwTM/poWI
+kKxkdo7ckYnOMCD6EAaCobGNAhNcM9C7aCS7AiCZCVBSDE03VEc+JNfTKc7
P0idPjDbtPMhIcD6syw8oVQR8MyBXHZb0LuOqI33w0bbMpMkUDTuz9lV+k6Y
qNV3dvASWGwTj54f7yxXbNt49CYZG1DgYMiTVWhIAAdTr9/6Tnt+uta21QDw
GqWCNDoOeo0z2IzX/5h8mqAL7PgLfOiDFAdCTrdZ315GRT1SMKHyFhbCgV9j
RgXdDZJnp13STWvxcglnIXoQKVPKNUiLRRnMvY5N4RPbcC+Wd4kOVG9Abu4/
p58uK4ECCtyk4tnF9XEHgiTEy1xg67l0obwLkZIQ9NzWzOLrsIajtcWxKaLb
YEi3sP593XOUQKMmrcbLugjYlhWhpPLN6Yubl39pTQEjeHQW4Kba6bu2qeNC
iGIipKq/Q9DDinNCpV3wLYSWlz1CWu63olHM/7HiuXdRFisqb3Nq8HexUkmA
uy95Qa5JbQAoUSWwWPeE/Y6sjdk8OTmT/aZUohW8l28VEnO1/oCCaRqNm1y3
0IE/C8NnQXRapTRsat7dKchs5/238jFBc1rlLk053LX9jIZkDQI0q5Omis8t
uux59b15b2Pz5YUu8xiAohsF3evqSMquJ2duckC/kZShJt/B6AId2P8vWkCz
5CJPyvz//nC675T5W//XAFRwTYs8qRVCzORFxOwcZZfb9J0n6I2UahEmHT8z
HcIARqmipGskiKXELdW4z140MyzCYKv0MocTyJCfchoQwt1E4yuHyOlXvGTr
Pd1ZHt+COGd6kDk7THpt9BgkBsn17M6FaaD/hMy07HgUVxTMUQjhmf3CAPK0
7O3pcYNAG5p78l3gcN9wgtM6EJLOWQdE85Bn7It69LjcX0jVDAwkercqeBF9
IMWpo0vr3nbTo4I26PKgAX+KEEsqtjYU7kPEmaaUeM0ksQdCobt2JQo+eMiV
3cmg17R4VNJuAK2LA7plvaMu2H1rPs4ffAlmYTEDuDu+BtGcV2MRP50shUKj
1W1HG9R1D8gZpYBp2dycUBOf9wB2xtwsF/8HA81IyH0uWnE1nsZwMoTxHFaf
+ZywHVvFkQ5qadL4XCFlgny7TUkFs2m3vc+0FDPGwWMG8QuCKVqBvs0O182q
6vrGo6JREyW/AE45v+BTDV3S0QdhbK6ZZI+TaVnqqNVHevH+ZrseoDYAcLVw
lZELqKPXENN9D1zHGfZs94OPg2tcq52uTr0E7fJ0wkHk0TmLNDqrjO586XbP
ZhSCLc8hpIwbdisqtH6gJG6TMpKlb30T+So7ARKay8biNdhR+VvDrPsAaDox
yMtm9ieUX//qdnyPPtCULW4LjcU5+CEDRZSx1G3u0isK0ttd53jh+kHeJK8v
+8zi2/BCxtd8RX2WtEoKn2lK7oX5NTzE0nDOsj/efc4CfUQi5rBmcS83za7r
rSqlnKhSeQ9B2EEZJQXjSqP6Ns1TlUhdGW1LasTUrlF6EmnwEu1pruPPgpKk
vTZHG4DUqPh5pgDNAAQ45gNmbJB8/NMMdpGXsBwIVI7Um4cdsCUwr/YScX4x
bY2tl25crQdmM3LraXZLoyA/Z9GYecTwJuwi/fi114lFHK7MBS9YoLT2vETB
2bLoifvFifNZ8CI2u8zpsjMWuecGvBDHIH0KC5zu6mfUzXlPlrONxUQChcR2
1oLHgPKAqYviTyzFhuzqHSG5ph4yJL367MWUpXCQkNMg/dl4A8UEhkVu37Yb
oxyBfDNpHLMHyF4O0fKXTpGu4Ufw/KkXaDbHStRNSJ74lWxkJZTary1tFTKV
SBVkKwVZEtFlpI31U2w6NKwxDWH2O5hUoiddZsVvDqcUfdt0JI5lGKv1EVDM
JiF91wpuC47IcvzvFle/6dHQ6eokUCwTTnHQLhoD7cs4M+ImX152hFfGdZJa
d67dXEpjhgvoL9W963IXtSdcpBZEPQYcOpQwCL7jSJcLx/wel6N0GMS+/bqT
L9kDZYitjQUXAINiHY/ez9SuCb8Pqw8l2EXSPPJ7FvSmwT5yDoSy0InyIV74
F+unzX2hH9Dk8gTFQsehTU2taE/3bX6IzsS+LyFLNkIjPjfsMlAC10VKw3Hd
liXLwtWNcIuZKlyS8VvvShNEHgz47aYRkrBsBoGXdF7JQ8rJYSElnVXyph99
yMOLTCGOi9/ht1YKDPyJRo45L88PNzuC+87kWA6VFFxQmIBFajnAe5uJm/8I
8J1Xg0LiwJA7jEcxSO/3NWYQuhw6c08B6O3LcM1482YMxjyWtrfgLwWCto0J
46l0zQ3Ftis8lUJ9XVrQtlG1wcLvBsvuIFExW18lqzswDpn6fM6p4pxyQtEA
G1kpcFGiX42dTEeLHOWryLUmqXpS6AYaiMe/x2C12zOdBT/M8g5hU9ah7ts9
F3tQg3KgmuBzZ0NkJMrk92vN1BXBOgwyy5qaaQFAz1wdA14pezx67iZ/iKAV
Ag8kYHkXcFuqPrqMsSQ/LSpoNaWEjgTuUEx3uUaLN12R7HawsH1+KX5pBqSh
pVkIRQVPbRZ7sm0AjHhvWplykgaUAXp3KWa5h7OfJcr9zoN6dn9B7Wo2ikmU
cMqelANNKLOAqH3nTpzLlkRLq+UeBolFM1Ei+C+vgndQblGrZQ+iNSeJUyTU
sGTk1NoObIeoT60XE3Yhib/MvZcbH7GEYmqxKYGzQmIQKnKiKMRLkn04+jUS
2GAWhuO7tE69R0vG1tjZB0LBMj4SUGbH/ADXjC633dRFdTuA6UkP6Wu/qyND
F2UJ8TWUGJO+hSu0hH8ru6OEVE8CRwZ/oSOs7aYpDRRqpSMyJIqh6H1GuK01
Sv5VbnqS6hZ49xgwTrozciqDap75vDHygecvTdBx3x9VwjLNC/8iEkFv92ip
kDORBi5EkrQ1Y+rPYftBHE8d0hfrhEwMQbldMnnhUxuYwE6iJ8K6XkpUqFaH
7ru2g0JU0ZQ+IF59VZCefjJBLlA1xYwQT4/WaKWVW9ARJQu9X5GUq2a+a+69
QpH2cFRzoFhdNfnJhLIpWbFnTxlUKl9S9ZRekLOZSeYy3BABd+RrD++GpsuU
MBvk6yjWDslEH7SGOoxJrwvWunzrByITZpwqd6qhH8GXD2vzgCdRM/e0gb8y
5eKkuB6CVJvIqt65I9P3jBuu/rJbftYfgaHf9cn50hwEg3JJD8UH0UYWpt0D
xvXWgU8LHrT0BUJgWPrriE8jw84thFCJALnETRmKTf5QvA3AudaRzEPR50fu
R2w3GAxJJSFYZHWabFNy3FsjHFl63qOtlmhtgolx1e/2Yu5u3jFqSR7+vGiz
3ISJo2GATQabl0gpxdESrfGZNVgyQBHyJ/h7WrPUc/oLrojmVI0YmAMctw7C
yUuaIaQterTY88eBf/MJnvADyTSlrIzrziseS7q4MegyQvxPGTf/YyyBAGI8
GFYoV/TF+v29vU6Uq4PONFS3DaUK+YFG70z8/uvEGfV8rQTQVzXb3BpbdiAS
3Jo5fuNGVUN11ytng8D669D/IExqj+TbBbkn1Ga3vf/md/PfGOKDBqZB1zcD
hRfBUrbj0aotFb1m6eh7oFXzGQvXLb9tjeLRFpxEZAgZf9jtedVzagdkYm4x
R6kG6tKRWNXMYoYtgx1+gffBjt9MVm26MPoDh6uc/NfSX0xy1BuflhzZBH8g
RNNdEFl+qU8a+zeeGviuKWYK+ardc1vC7gJdt72YLwY4MDHmvYXUyCtQtS1P
D4etMqjwCe+DN1GNhBqq7n0LVjVS/xkdcAvu0x4jip15Ie//oct3/MdoTuTR
m17Q35aggwxnt6wpsV9VfZTt6bsuvA==

`pragma protect end_protected
