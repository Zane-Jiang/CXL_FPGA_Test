// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f6qsmLhW2N5S8vepzGs1lT/Eesl+1EDCBVkyobmu8itivy3xyRmgLfbSp0la
OyozW6YDPhbk7wgRUDUycAhwUD2zExnJwAXM6rgzYa2SD0JsqhI1al8aKUKz
bPzLC9WPPDu82hVympiZy7areVBSkPEg+SUAsZsmc1bs2db0IleRut4X5W8h
fzfiRakD2VeeH4P100wbSz6zSxpZ075r5LVxMubnCy62ICndSXOEaXGEZr/p
M2z4UZTcNIrqkFl5HhL+zjUqFfX+FQTaxhr7eX47zLNXRRwjgzVFeAqr6g4k
/6QbyUMonhtQKABfa7PikhIN4C/EgerxFYOgoGO6pQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IHogYnv4k6zfueuaMcw2q5oa8+EmFkAfTC23PcMWGsPVxzlYeBHXMt5zRIPx
CJg0RJoLnphToUoN1pO+QWtHyxgybfVCfFRvL5E9bEt4tHFZQjNnvogHQfkW
suQ8mlq7nqxg6Qvr5F5H8ss/SZWKarTICq7TcWwETg7QCSUzcErpjvcRImIi
YicDk/f/3lby+FH5oFe36Stm6Qb9+Of62rUez5ZEm5JuraU2KSGIDceY2O5b
BtC6XKUeOp1gGetyxYLGirpJrn7gBFoJSkwB+l5aQJ+lZ7GHVpKHv8S9i0GL
EjQ5YdL/ZGo8lLwQVWh4b8JTy0mVaYFVR2BOtfhN9A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MdbiU/9rksnu5UVm5mNiQrgdwJy2LPYgQbP+eTCg38uUG6KqIeSkcfn5i8DG
fuW7IuTB5g/lUkZZdfwzBuKiQjkE1DAktJ8YhVQTPOU4YtB2yC30Xw20eTO+
0HtnPqBOf3uzMXaIrbYwX/BSIwCEndmYdFsm4RB2eOWbYUQTQHjmXJkQemtY
MrVjwbXaGTKzseSUx+B/WKrZIoISd4pEHRX/MU2RKu1a6omKLS5vJiGrdU8H
rARMddbkNh3kAcFh2zb52Qw/J1IiM6r+9GGTZtS6vXGP/8bC5kzRCGVbecNG
N1eTDV1pw3lEnpfwQKbfb2M6KxzXWd3m15FmocMDoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E/yiYDX+fqOXxlj3UhbqxHT3Wa3J47WUpFWWPffWsPAUZNchMTtpgnjAIKkn
xChfbPRY4nJ0WCxHHujICN3jEsfk3Sx5ZlkskPOdsNQ3QMVgh2LNSmabdvyO
R3AnZB54FCLMxuXp/vYA7bWTXpG9g3kkn+T/8T5R9WjOVYyk0UE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EkH0MdbETlMl6tOhsHqqN9Fj+zsQFiAIHfBu9Q+qBC0P5rYF3B7sttSNzGbO
HTCMgC3IiR6eoa4NVN3uNfzwyplMG3MLgJoy+RAHHJNBQtcCmqxFvCacLWqe
zXAyqqytPNPlHRbh5mK4yKRepaypeghgjzScnOEz8AI0vIQf4oM7IkhcyBuZ
pjN9CJ8apzucRvdecJ8vxU1NzM9Ne194mwha/A1uFH7/CDDzxY2clUV9qgEE
SZvOVvDZ7AwnvX4zVmNx/PNr40+oB3oNBNynQ0OXCQfKN3h6BbdXziE/DTYl
snqSJvmpelVzOvbzwd4OvVuhZVWiJH0iZN2oJ5x3RIG2518zUrNDZkJ1jB0j
29BIgLHA09fFVR8J2OAM1t8uaSBAsIdD4OJnRA2c3IPKzOMSikuU80DtlgxI
7tsURTind2GnRL+teq0MCedtd79bY8eoaUQhSsEjtrtbhrXgqELZoClMlvjo
JcTUA6zbOmu2V1eLA+W4iFk/0B7y4DAy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fUVMQMCsZcO2EssBYSri7oLDoLjEaHFWyh9RFSSLFMjONrAUH/Ia20lmHhNU
tGhp3zEE5x3gZkOcV/swtIjhfRvuBTnBgvbx/MGTsu15w5Dj/SQwaQLg2hpB
Q8FDU8Tr1Xu0RCNIPLcI1WN8K0x3ft/bExqa/ALlHJmQmH/TyR0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iNH7BoEDJPr2rVRMOc5Y1b5t5tc029WiQsP5ZGAJF+/BK1CflZesBPPuUxtF
janyM25pVLPJz6HBguJHrqXvcWPbDm9qj+PRy6SWL2CkfRsIpfEuOZE38Q/4
0stILK23tu7towzCF+AW+Jxc7ouZS5hnTP6hcM5tpI7IH4omQho=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
nvgLzsb6sYh2FCMv/MCQpmpVxtCZup5W59jURyXSEzQcIcmZi66XTALAOKcy
PHN724Lu+sS3NRYe3rKPb0ZqnfU/FvYhtJhRdZWDYAtFIuukS/WVzs5pHIsZ
VXSW1snb94XXfueW8Rgjs8DC0f/6bSRHxK5yMLP0eIVbHIBQh6Uu5cBJMi53
kVC4gw4cPPpRrls32jW0zPGYhUUZzUvWbCRwgWOghUQPWBAIZKlFNx+s+Nt3
XT2mmcHOWYcJzB2KMEtzTmG2dgKYBL3AnY1WPsBIct/vn4swxCBPimpGDNsj
Yzzrcc3RNt2zJwFOdDetBcdFD4IPu2T72/5gc0+s8CJQV1k3tbviWD/c2ebs
J3JMxYX+sRjJVlyUzUWIGcmhzwxRKqUHQcj/jwKQaXyCWfm94vMv4xX3Npgn
UkhdColHnKto9oAL4Dok/tjdf3H1nUJlP0noQEFakiJc7upFf05H+DA58A6+
deJwdFFga5KdKcLq2jOq/AgeKbBTkBVvANVjlXj2p/s1Erlr2kHRCToDkRBV
ztjYaxSO+yofM6PJfjGQet2vk7FbgGTtU9enVgxlt6XUdnMI3qI25ocDcSu1
RMgiAu+kn5KEX91AHPxaiF/zzvrjKxrgQq8S1LnY/uqQCFbFTIbl6+NXZttB
Alr2fDEhmM3q5NUyhfBtnpxph3rhAVXjEaEBr5lpR9rv8+vb1qHDx8SMCHp0
0YrqdkwQxODvOfL30R7HHXGG/RiplKcEbkGqmoNSfNLjtSXPBVY3+41odnbJ
G+t27xeelvmnWB13yyB3YI2efLw4Rr/I3yoIv/j1iBakGFsupKC6n4DVpIKd
RtsGr86fLg1IbWGNmzJmz2D0BJBNiMu6MSpGnENiHX5BD9DTLaFcJiU+3tdO
07WgMGTXmpLO9qX6QgFRQ3g9C6pyAwH9OJ771J5/qe95pHpNfWjQwCrA+KIr
raaG4u4bnuZONqfx1A/ER9r8g509ltjzZ8PcqIRGcYyEz2d50Rk8rIMv9sk5
1PKaI81S1gS1Q/tHCTuARC+D8hxrZMpZlwD/gHDTKlJfUslchdeAiqi+n48a
wAZIAyEAAFWzWUNsWvKOLqjX39jFSZ0g6rfCeqCRW5SCXCz8JOf4nEbiMWBJ
626slkTY2wu1bDAS71HPh+VJtbUO0/SJ7ws5RV8xUHRf8d4ov36A2qF7KZ0e
YOBUuVYyJGKMTVotvzdhWySK6hMw7WWT4wgY5wUziCXW9EegGKeCKMED4kJX
xyN0etDO26+PqiskFQ4ZlPWw/s6Bhdog8BHIiDSRDw==

`pragma protect end_protected
