// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AqR9hHZtUmF373Rcc1D71R61Z4ue6VLNNaE2QjrVCO7dgMmhIRDBN7USPkvs
xG0VQgThvE5JuNupKsnWtZhA30nIOWXQgF7bAQWMw3Z71lIrEq2eMj1IInTu
W5z/q0TjzpaD3cckicGOCD5qVmE/ZDwf7siSv1DtKyB/DcAyp3ZPEHtigDUD
Oz8MzR7ZKwygbvgB0t2MBExwhz6RTObzE+43XG7HPSkOXlIs8SAcu0tQx46U
QVi5+C2K3qhcx8DlEnwCckCBEBXK9LZyeVQtfg9dZTRoSYkQnW9whUtI1W9Y
HTPiCkMk+suGbSNMFQmNRxYijQMhdfzRSNfpFGIfDw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Z9gCw0Zu+mmBDcgJGUccaq2NsjR4wCMPCj+kzylYiR1J4CaFAERoviHhsuuz
cST5x6nao1qbM8kdpQ/Ki0gFenS6dkceJSNNjBMwWv+EC3iLGtHWcLPUac2v
7CKO9rDvoDoyuSgwaTmGTWfOTVRz+GzpearEpOAMMt0ac4VMjlq0JheZNw7F
A4/ihOCHbabFYLMoz6X7DK2Jnkekbl4zTaHTcsfshU+YJzma3yPxyGKSiJMx
wjhZTiUg0WUAgEZ4J9bgNCyWT95DxZ/kjFlbmRU4lqlHj1NrspJfXQDoaH/3
g78M6ZvSrOj+BSe7Tg9dnDtEQHMPH8nPkLlLY5xrag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MLjOJONPesNyJsElnkNrltj3nLRgpyzhkbQpfzfcunU4zoeATRT3RLXez/Nf
DPyRkdHmol4RxKwzwQ7Zr1jAp2IbXUiPKJi+/iTVbzgDSfuHJ++ktnQY1b6Y
uOvA/gEOfcO4Lk6d9zDXCHYc7jchpb3MV97Uq2tAEfd9/Uyr794RQVqgkF6t
z6DbeFWOjynIGNESuM7FAEfFDWMVuXysjr57HJt8iTyYpp+XwkFX9DbF2VBU
TAkqb/6VaH2Eht46w9A75I0m0KC6rU82itqYXiP8L1dRrpKfHFX68zr9QlJe
lJ823K1MpXJLT31izWeJAjsPklW4MGK+p75FYK77mQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GDQjyQLUnskQTKzIAQtnFWm41e0wBjvMkHFv6O+v2fHK/B1GJ8ypvMVferb8
lWw978j5lPCLnAkP4PE0QgYV/dH6+bifAYfQ7jnLE0y9O5yWz6jGYERvO153
tlg+/AXAGlgJZ+tRy4xXGOj9jZQgTpz9dncwNvRqSvmT0DmqSpw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NfopPfZpIeeYqTw1RrLJdEUL21tNrmQw6LS2vN3oJ0CO2cw60n8JWEQmi+qE
TV3467JQQyZvHTrJ05SI5UnhyKF3+3X2yvJovTQJE9XNIs+GqQBcqgpFQfL1
tXEVyF8YdxiWh2B/tcKr1VcBKPmNl4FTDeFNs+ON5qigflhtm/haTn/f9un1
gqQc6fEBLEbjUycebb0wtD4PYbd4TXktJvRl4E3JnYnVksT1HiL9WJmyc64w
4iOQMeEzJ8BQLWHs/QPnqpy24+js0m0HWdwmkizZL3EUjI5tOQ2Qkp/SOvpp
z3Ye0VBO04XDvKWIvBHahF5eMZgxrZoURlCxDZ+M79vF0I32cSK0X0lmDIzY
foXhQIhyREmzYbr/K1Apbj8IPrTVlTo1+6WP/3MAQHSBrj0f2Hb77fpE3P9M
3HCJt8I2wsK5CEGnk9TJf4J88cQ1bx71cOXr10HkrLA107YdQZMWoQFE0HHw
Ztrh0QnoLfXo1VHOF52jBYYTV9rBaZUl


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PLqFm1dlqDJb1DdVCYqiwyCRYjiv9WTQVtjr0Yfz5Xh85coF9hF6SLaG+BJy
3o+ce7L2xIezA3rDZUglERlRp69om4flWhVdYQGJUhxrZNAXsd4R5sGWrUaC
h1oHw7FY/hzlhKyla6q/kE8rgPzL7EtmfJosnN68OzagC//8C8Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eKYU3c6fF3CxGnJLpTtHMLXHnem+bZoPuEU8+6wncwziZjUG/V8tEN8X4i+N
rb0R0OMSjC/lvYI+jOeLUcocIFVkczfDQnrL98HsAgWCvjkA2rfsEhsPIHAM
DqIVF7EfksiapI9l4iHju7HIayAVs4tSnqyvSrV2pIySNH8EkAE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 196464)
`pragma protect data_block
z5HioESD2/X4UtRpBsxZEGYCNqePq1qcy/TnPv5XM4s8SLhNpFiDXqh/SSpv
WmtTBwXFA1vDpbIoX46/uWYXuLhoJvKfpm0EzfhTBd1aedqxTDzE77Mf8lEg
8ubytEFQY1R33A0sp8alk0TLvzyfJiiQ0T33QBLJaECdy5k9EOhWJFGYuePc
M9L+ofkYEklHa/LA4AW9yFIYhUVlmg95GD3oReT1L4/NGU5pyzECgIe98QZh
/5uJ66J1JuaW0xLWChRIVlSzEpYcdCJ3VgHytNCLj38K6kBGjHnQ8qvcwNwO
ey+kcWNa0MDxNE1GhD3XRYVpbeU59C7VOBDNTl85CaBB4lQNTSOCLUpU/ukK
5knsWb+J0Q3sE5+eoublo67Q2JFnDI7eRheU9AnKP+Z7K77f8H08fBoTe+oM
RAmYTSrB1q5R2J3QRxfYqAjGZTrqMQcId0n27WgtPpVhX2SYu5QV2yfLTL7U
LXiqDUEGEihZropR7ZB6nWbt9Ey2MxgYpedXX+rtJPjF2K0evbh1bzjDgmkP
xPBmvffJ/P3DdZgPa9oRgdkQvtgNUMv/VR62+s64uCsTRmfnpjgRg2b9YVl2
DGFBOmjOGteuNJ/gvNsOfVXVNK3q4tbM0fHhyMupWP0A9OLUkegR4C4ecy6X
KIZiK0tHoi9DLQ0ZPcKQ8FhVAAmr+rZbIQl9hL3ylBRnSHr25g14Uwzw1qLN
/iiB6nEN1GpGqsm/gWz9x3jQvR8ZLz+SbnPqiLxh4A9y5D2WXwqq2oQw/tdI
zGdLRzIBAxQgnDuFI7feRl9yNiydBkdxTSuNcmQ/b9NG7mcIwkolO5mAonyL
6k5sDJl5xtIT9wUYSrYBusKwf5gXALXVTgUaUUVTzUxNyH1O5IPS1RT+GTxd
qTxeVEyg1GM+GZg+WHoTgqO/7MsRMMD01l7Q033auXQgImBi53BFcCK1QCD+
xvsHAt2adprkt/UZNTo2phM+F1sq6DcpKIXsZ/HTxYtgCNGIW/3DKldWXnM/
z0ihGjhPFc7WA5iwEykvJpJVBZHwbpWFPIgWOsfBZagDz/7TSujuKlU6XUze
Rk6ACBalpQvL7mKQvzxFqs8FJaLUYUwrPZtYjpQ1Wo251E/nuHyvO+mM7nY4
SsfNbuhy0Voq+n1XYciRVpQ4YFAFQOuARijEZ2cbKfctRA8Q3TGCWLl7Nd9l
5X5qcGhfVR06J9n7I4BnA+KXUZvWP9xPrSvpqgBYHytmPcsZF+qKTBFxV7a5
KCuM6fYj4FQdwkAsh9oSeYAubQahF7/Qoj0VGNWoSuiVnXFEVtpyuACN905S
pJvBvCeVNv9B00CJyj03gaOVkQdETt3lqCn7YL46quLXjIfTjVcBgyfnsgNv
pzMlmVD8ESJE22IFC52Zt6RCs9Je2Gmgq/ZUSQpVJqdMAApySeR8Txekswmv
FB03cDEroJ+FQvWPt9urxKZ6To9gK1Jb0JXeVUJ/4s+uexn669iMxYxpblii
1WKuhA6pnKX6Yas2feeaejTzpRkEh46GzA+oWZnYU4uZgz+PWChfH2tZ/MhV
xxA1hsyHR+yRwqEQAMtyR+2aV5SK6tZjxbBet/c/ompZy6HqKQ5ZM2X46oC2
KAivhUA2qPYm0Ox52jSx5OJg8uThG5vF2r79qbVj13Q/K/oJDa1j7+Sd8jUC
YwALhZd1RaSgx6rXUtEelALDbar6Ej0b5YPwNaJLO2HkV4bT3Nwin4Ig9czG
kJt0EVBi3rYbnq2tUG1yHrlpIjE9UYbxtiokeEyeIXUTg6bFFhIe4j3KCjJV
kJss0CK2VBIspBgHVAAqbvFiGwitEVim0gdcxCKcqM/Iq89s2Pj+4zDIDTFZ
bnkG1T4xF7sWv6d+/V51nHLhTCXMcSliLEGEjmUR8Ujq8yfhxxwLtTjpgglr
m1WU3S6z2efRpr5OWxubTjN6IM/lDxW06yzz62r+Iwf0DxwqgKmfQ2FpwSaA
dPP65LccvbmyAhnYmVRP3uW18yzUoK810a9OF0Ek9t6ybDRLjCPMh/mi/MEy
F+bN7JvuntyZc1tKrzTJ3NmjR7XHCFLtSeBczMnvso/hmvq9IzzqUIt7bijN
VZb9ysZrIcNSWfN73+gg1WeX4N3HkEsgl4cpYPUOcjUdl05hTUhZPJ9eQP6y
NwgvTbXjWHH38jLDnQrxWr/H3RUyAbyaal+bPo97S/95nJEkQXce7hWdmeUv
bVcja6OpwVKYONXkhDD3uJtBa1yT9qcoaZ1wb7uUGObJI0YqfJaWAxwqrGK7
k6YBulvxtFeGd9sFnWnN7+8wGHYqAQs+cKHB7iwhboEialPv2m8kSbZNyaoq
00BBEGyv/kfG5mxMuemT/8oi+BZHlsineuD0Sd/j4alyzNs26+hWoVBmR/KP
YR+vjI4gjSZYhLMvvY1xlaVfehKkWcYbWtIIqPW2Kwezcs2z/hjgzd8/q3Yp
HlmMfVcUps3kul0wZ4AkwLcNOgYCNwlh807wY8ZTsGN9YV6EqHVxYaDqxlNw
99DCyISfoxgzSVLxfGIaar3dMD16qMfa1wiDDE3QvpHP/3CpXi9bI/c9V3Os
VThhAUqniL0CukUFG5fgBapMbCwaC7TKgD+LJYJE7NvMXyfdJp8p3nRP77qy
RufCcPgk8LC1c+wp4DCaA90GzmtN2tuhPXjxACgtS06FZqC9ocdVzCvd9rYy
ErVEfpVrysV4Wt3UrtfvwAz757ghOzziY409rrlo4RupS8/IG+eogd1uHt6G
VdTRH298DNo1EiAYcuGqbe+sNQM++1fCjtBxj3QO2j/Vq1lZ1hvDaJwrMkbE
r7rKSAI7JXf+OZuPR4rrACGuFyygPu9Fsatc8+mNA2yYwS8RT49TH/3Oni+f
KO+odgv/a6EtLNUa897YPXupE+HmxPT71PkKrOehhapH/xVdIE/CBt1YRRWF
UPam6RHka/LW9wdwyHVjJu+s6yG2oKGvvYpVK9HWyhBOCer/Pca9YlgdWClL
yYzYqbDUh4duAPPTCsqoRHVOBAU3Eq5t5nW94tQYHzfopeDgYRIvQoJpIpLy
Mdprog9nkfATYoIcrOeKd7sdrC9OJkE76bBMVRBQ7sGWs1ezDr/eQiXTkPHp
UqpiaES4A5WXCjZiUVlESkjT9+KSEZRcxh2irgrXt+u8nZ1N9fPqSeGqgqWf
ZK7hXybY7KpzVbfpzphfaQBJBwTSzkZYt4y2XUT/hVLTZm9hY7L1dtEMcfJR
PPFPaxN8w9ipkNIWQc5IPDLf2sf+AXprbhG5fMUZYTBsVFE3NKBpPy+BldTk
8gFNiVXOJLF+lEKJnlzZhG3Cjn6iU5r8fyv7MKE7BZmhCeCeBTiAHujQdJHV
xfMlHBbWbVYM0tuJB3NNAcz3Nv5smffmV9tf7s5e1vn3FlRtTSbgKXHV8Tvj
gIU5R41OZfdoFju5U7RTGSdOyHIFQgmuuGahHgG5uMC0Y5BZu4Q+h5KCOl3q
Aw7sCMXrKvnTE/VnMFmmmo7nIinwOKBeQg6a33/31D3jKoXqkpisJGRXWhaZ
y+wRbraDBjd2Jm85ZOYGhKMBtzemX5yNY4BsF3YChdURAH7Efmmxj/Nu+ENk
IewKRhLWlnoMlQl/+8NUuVu18Zl7H2LIXZD3yh6hyDZ51KyZ7H9ecDRgLnSh
RoxM17b42GgAKnhPQx3lCX7tYdqbCsQ4XRhBknBVAL9kDdzY7zLUtw4ybA5K
spPR+sk8Ly4bAQaQaHzHwnxhBidlta30gUqlnM26FG9rbnPCMP/8xevmKVBx
pLuDuW81H9pwAJtfhHd2PYorETKMjU1dui91uz1LCND5aK6doYnIhbEnTCuH
P1SyAp+OFnfYLhQ58PTrGk17JKEQBN/lh70elnas0YQnWNMqdOzNqKxsJC4N
KCAnjKbWNGe0yzMDLt25r2/gyLjn9rzg31yymbUul4VW460j3nBxgpPRLEMd
j8uh/ZimHx+fpckz5s6Mb17NoN0V6mcfGBDu/WB9qkBlnYsCkIDL4dt+TTW0
w2DaCQQ0Ak8jaa/46cFXOc+PHLCfzG6dXlLldYAagt2s37IOVlS8QS0H9JDw
QLDfdh36526BHay5OwTM+9A1EuTN/9fZCfyLuBC1Wi5PtXuWi09Wc2puHhUt
Hi8gl3ISOf9VzKdMS2bWWJYmIPWgABMAClcbIAHXOO/iXiUwKKUHWJ8ECEL9
/0rQdeAkdejz9zwDdYqlGl1fgRnm0EF8X57cXPcIvD+7U2mhXO1eAR+bR+1x
OUVnn+Wdr4TeVVrTmEVe5wmbwLnj0FsnDu7Dtv5I85oWyB5PffxpD+57Oxkw
p9rOp78yVMnjhOxWLQZckX4+qPrZNU398aOW4mWJ7dRT6rT6Z3mXao9upNGj
KEcHX9eq3xzEDz9mF7mlIs3l+URTtqxY1buTzzcwhar26njGhTS/Zeu4Tjaw
alBsTXb7gkdiA3a975NFuDxnGinRTe2wxKeehLQuAMj+f2rpr1NiCE/iNgbe
zJDu0094OEOf9CV6Gkh7o5+V1IPL+L6UlFyoCDUESOQalFRlUrktV95+QhfT
wzrOH1T/vg3nO13EvC0vcCx9dNdFmXNbjrpt9xwGJz1nBxP9iWhtRQkTZqGQ
B7DKs8VbZAW87VvAT1d4KWRG733pKl2oL0bW4kWivQjQtwO6dk3trn3+71Ot
YEKV7Eg/3DZi5prAOnpMXlVt0xBDXVTxpd2EqMr7RAQ+KH7KUbCpIN1PXng9
lEfBrKaI7PhjrujuGaaR4DnqAturgF7Edu+jrtH8YsnpQ1QiQcKDJslzq0tU
Uhk+DTlNOJKErVfldWVKyiUiSmdBkuPBPcm6cwQUhY14eAUwDSVMTv1Kwor5
zBFiHZi4EewHT+mufwNO6cJsSUIidpxNLQ4tDh4PmP6/4SYtSXdLZV5R3Shy
elUu6UhFkd2WnPDXSOjRl0bPnkqFPu8rS6ddGtpe5wjVrRIMd3kUHkNGEcnz
7gYRw9FeEpuG5obCrlbLQpM6JBdwkHKb7zLnhm3sHOJ6F0coc4KiBS2/cCMX
coL/x3FsCfhNu9o9eFYirgNx3AhSdbQ+Y/3R4NZN4ZlFfRMchubgYHKI9TPN
wj3HaKb84RIuS40abItxZC6DhZfkqYFPGsqC7mamfKO4ysL5P0JKwWOZlnne
nR1C4Aw3euXWbFenHlBgBfOYM7/SBA6+VPgGk3Km/F4ETkB+JH2xHw4s+tyT
9sxbyhNZ9aq2IFCC99ipJB4B/rU5pg97ri8rEk5b72vnt+2gtiS9GqM6KOwG
KLJ9wmrzoKBck8C7oYVunIotrOaGhibhrjbOnWwmbxaPle+jbtFl1+UJ/0d7
P3FCAyM0dKsX2K4H0Grn6NI36qx/QZeHEuS8v0WVKTjYiAiu4iYcPD1LBHRU
WoC5V9Rzl9MIDuCzLmWrxIgfJJfzeNqEoQa3RHUGTuJrtBz7R06/e5vzjH0J
eYk6T3YJeEpqS1IqiaMrdK0k8P11ELz2gQyOAQfwMRc42ScF2prZVZUsIj78
OUEaW3nGGlYKgdvQ5QexFg9tWG+uoeWpsBWQUal+vgL2Vjj0JBaJHfFqBKgn
Vhx8fPbtsX1MdnRUE0qrKybtyj8D16pfN5dHVpPo7yz4fMZQEd8j6RkLNpjG
ijAZQgabvpq9uwyAlpZ7rtX//3uSXbchrjImrRtIi54x1NZeO3/nCz8VXSN9
ZW+RQsIvQXaIeMAgPiswhA7Mk+s2JbGxi6sdxYtz5XhIKNvxKi/nPfX3BcSI
cgeY8I3i8MEi2/sSaskDMW+0szW3F4OIbkXZ23ZQ3VkKf2Nc9Zq0KyPuhgI8
xRIRXZDb4HgO9c94OPKOgmOVJHPhXvI6QpS1JvDnAXvYWdPpa8wu4DRu/bB5
+3M40WtgFkIw4jB6w8a5/u7wCKZWakL3Lsa6FChah4bvsMLtTkbXcFi96tPQ
0duj+Os141tqMShSyJoxTsX0TsdfjTm8yenHt5fMOkkeZ/EznmeWwdReT4I4
X4YmztJmcPRtzT1yZd7GAbsLgNjxPqFhIDZvmcbthpMOG9xVaxaMQQRGB0hq
d8+DCWd3IT2/5cDJGtHLGZxOoiYGeh1XVz6XKq8pPhPyq0WOF6VJc0gTkaxO
I9Gs+VIzbnVs6KS66/Jm8mKpDlHFzzRwi8vi5LL5dAUv95n/FkkE0aM20IIf
+GJTC31QqbovThi7F1OsGtnDnx9DeaCvv72q0H41SVz5E6nW65Te1OGB7XcN
oVFMNH+tq8UWOFPW6kYm3UmAQcic9BLlt9tD89Z4UAnDD/LfkDzvloxSrmSc
YX0jjDxAEsam5vQv9OanUxGGVOkuBtdusSWIUMlLBzykwVl9nE0SMC9iIN3V
MkZJpUQA8nYRd64RvrOMckBOhQd3hwLVMonvcgv+dfLUomDfKMVdQqqpKdpI
wfnfaE8XBiGM1ADvKn6IJLGwrS/ijOaMbJQy1xEam+FQthFRiYnhygEjeBLE
bexijeI84brKoSg6OP0CcXKicx4zZnl1fVR4l+VYj7Qc6BstxLi74yJXLTU7
rJOIl47/xxNmoQGQ7NBLMrMV2YvR5pKCKkifbHlKgkogvkPjbGHw4RmPWiDb
bjuOsHV16QOy6wvAaDcPK9JdWgWvFf+Q18tv4krUb7HKtsTvqu6vnm37FS2b
wsy8Yp1X1SakT4/YAzD7l18/YqsHgT5yOAfvup3QHln6pwEQJ9KduDG67Y/L
UrVirm/aJvlpepMYg/x5xNdGp3gPbljqC9+j1wetJ06cBenIIjZb7mGXZpfE
vXonKKDv6qDo0TaE+FJ/WI4wpfC6TQOb5XpeGWLW9W/VAHyoj8JrcwjdGC2G
qxEmeqAwZug8VYWL2kdmZw3kCvvHTMIol14sJNd/kv8haPfeAFHkYG4YLsiY
s5UloiUx77rerKk0PFz053KKMBPlOzDCKNVavp5C5ZJG6gqxcObpyUCiCV4A
BlYOPAjVmTHBwJAeRxS9XWpHayynoDKPOJTRkgnlvT94hQM5TJOV1xVMmT/h
McrbaFvbQc6pvMpWg4YemrQTSfrbzwg3YDch52nPImyju6cq3m1EPDN7w9Hn
eBUMBGNX1FvcJb1XopVx1ywDkj4aXtWulRzpaWXx975Qgq23iobmZaXLd3ZV
DbI9nUXYQZt+E32lLMMSqLOJduXbmWhTCSZgdPsF/v2Na1Kvxf4pjXPy92h6
XO9KjHs28C/s+wsWsyZfNVEnCoc1vPjAilmS9zazv3Wir2ZPc9UqqrCC5/as
Wnjw0k3nlllW1Fz/UxOqEoP/pCIJOoOkNEO8CVJlJYiggeQLCAIL0v9nkGTW
s0xNrTP+Wn7LOcMmcwOs4h03QAm0+pQ3vNARwSFvBu6Ogm5WA/4P3KnZb3m9
uWTOvB4g6laLhcshNioDYfbuY0IucN4EMNQpZMcnqLSGXaaTZHlerKOKPwNC
bp1ltcYH/KEstpQ4IzlFCaGtQwr/95PBRc80eq3NlWp98bJUW1COBXJcA6d+
tVVPOgb4OriWMbPIakDgWdhXWfUCuT7WYFFOhqPZgYfXu0jmLXFB0Jvy2o9G
GJTfn8F0gYNHTcZx/fS/v9iIRGZuF9FXrSztZ48rinSFvYkxfXv/VSPDYKHo
KHiasY8oAhpqfED1n7UukJgo4Qzc2yffxnXf6uq2CzYeO2655xtTUNzPopAV
/E0N+aQAn1ZlihPSeKr0NVLBr7DbzYn/RktXsxIboph4B1JfoG6/yVZ5iXOi
ZAs3xHZ4wKWFXJ6PEAy+Nq4SYgFe/f0nRYIGY/PLXP2SuhMlpVunSUKyZ2II
cVp79d6mxuXq2FkdwCVGdX3YCsuj3OxGE/PDO5S1JJSn4/iWD1huqTsAP/T5
VI/N7Tz6UubAY1fR4CJrOnrs2JavklAzdPsjepBomldBONNnSReHSeheEncf
Tirq/KVAO5yhYZEuDE+58YPR/1PeF3E5aN0aQrT3FygalNSfvxWghF9aXbnm
KKV4Kvk0wZ3950vaK5U1B3Z44MIZxGE5rZp3tP9QD92+vV3IOuQc2hPw3zN/
dE53bksQjf5hVgXHrv80AhcYMOaCUN2HTMo7toyIKdwaDryDtpAry/CosF8f
dVkyrrU/xVDdLv7GdeOGjQ1cihXZvA4UyzEDmjJb5qoyDLkqRDaLCP6OwzdB
q6dEbokPS1xXqf832w/2epp4Ly7nz+6Xi9Vli9n4HyYQdxeza5GT6C5IEIkB
Cl98HDq1TpvUW43wiOHosnU8VWefsylvOfpC83d0YWgmf86OqBuOabZjii5V
HeoFn8AidCjgtfb1VDAe41eric1THJQsDji9O/NsCqyJxAbUnjTlrbqIXfgu
Ro67aIoJdfG46WmNob4MzEOe7R4v1p4xpBjUvkzKGmI26y++uJP4+4E57Jll
GE9ntX2yS07DYe6VndprZ9TTb3/yVP3+USNoNzbCoB/3QSV6x2vbAn/xpw0p
mcZuRP1er3wygrA0Wpk9YACPWajlJJHHPFXk4iEtpAk0E1xt2cS/uTPoMuUf
mey6KdIad8rYkkamDMr7kLwoSHJPUkSE5U94omWUvIZ2yKeOfW7ZUUK5kvpI
euhCikrsNpVH+rDVIlJ4tL/IMbX7zPa+iCGFknmZoO26IAOmpuU0mvPWbTM+
3Rlj0HMey3VTiY47e0AKsQ8qkLCK9Lg/RMCONPBPCPC5Jz//b3CuLuv95IsA
iN7ODI7VOEjg7QpYdu98JDVU6Wqz5KzWVozOCyK4mbVoAQwI0900q5gScCLf
Fmi6xIb4Fueaj7okNxu/Thp3/4IqxRTcQjcU+vRWjnWIMO+h6mqfENFGkaS8
xaYmpKGZskCF5tuPhDqiM6Aj61FTfGsXZazUOzmUW3RnhBAIPWRvIZ1TW0D9
3hWpZfuJ/eWTJmKZySKq+BtjrP7D3KtGCgaprKlRf5TR1pAyAW43CqYwPv7J
UKgCOcco8Kej2J9X58/NumVWx2X6tL4hfzEItx2ByTcbWFyjHeRXmWHAkABx
KxcaqPP13+lQsNFCILsqxfC7JPWNJ4GGzZtaMYkknPHh36eIEmhqowQtclcw
fgymZ+EpUDvnlMKCzQYDrvybCypkpx71xnsK2duuU3qrSpoRKOXbC1Z9NyBu
GrlYgPG02rrqOHMVCoLn7F/2jc8GnawhMoRqnd+Apw1LHAgKaghaRiSMX+u6
tK6r/51dCuCLQaSquNAzcaERVLLJCDizaGQOlWnylWdhLNYhNjTJX0NZov7X
iDdTkDluyFlrfdMxPcFCccS3lwMq+W61icIv5skzL+7DGnK6Ql8x9NjKVod+
m81uPTZXXkz4ycA9Nx8ge0JL131/yZh1SyURESgXWyqpzycHEMrYHEvPKnR4
x7bZHuLtJ0HEwqhOct355ePpi7Ws/aR8zZiVrJkVd4ylrcVFf9nlzZ9eF8kF
pGoczwYIvxToInqiJeD7TaRmsCOzxuMbUmZMsG82q4MCojdytPx9g03arJcA
XrbDuymqQZ/mr6+XgQAm2fWFJXqUEXye13XdjohsAfj31YFtAJEWSD6P0xxd
tFL46ObbJEkhJmE0ID7/8lr/pHGRgectRl8mgZDYSpiX+SBggj7BY6APeQen
KMWAAg6rGvETsj2g3mSSbrGshH5wqSWElYl5K8XEBKJ3pf+qD9wMWuNUz1Nk
0ePgFx8AGPHAra0z2Nm2voFJf4+mkv82JxpWLy+u7q9s4wf+bbYM+qzNRjoP
vwXrdI+2xr++1+yOQQkWeOxER87uYRB3YZgD2POKcXFQHpfe8y1lV/WTHoMS
fM1VbgbwI84p54r7Klidd9iAs1lNgL8Xzi6uSRcrXk07ux/qKlLZv+hU/7a8
5BENIzTfE5wT5dC1tI1FTNTAPDxmGc75EHqVdeJ3BBc/mQLqPBAunSncZepN
zunlmFf8lyq6lBZx0wLlM9Laa3nA/9GSbm0YQdxnjPzZV5EWQD9o7smphSWV
HhAjKcTMW7pV9wxMM30jxp+g3n0odYgfkf/Rf++6Z2bgBdm86ByhPHLZ7mzN
IPDjkTyic8u/z0A4b8xcsiCYW7x6qI/MW7nbjr8Edq09d+llhM3444RO266Q
s3d9ON7roOW0Loa3fZX2PgA/P8uXcXm4sG7bOW4otsUbNAJUN7M57ZKkK6s5
KVf1PvkT07HR4GNPdZWCTSdzt7aPAQtTty42gWExAktZy00/qqzWoJYLchi1
wC+pcFGLHC/AsYCZFkIvAE1pBU50wZsIKQ2r7YgWbcZElEHO6q2Z+jlQ+tPj
P4L/N+cQSHdCaMRd2EG8ZxScTy2hDFqC4K2C6lm2jTlSMrjlColQIkMll+mS
LsvTJH8hYwItQ7VgeGdtGI72976eE2IZ0I3jiAichUdAb/IFClqosmg+tGps
7BR4nAC8fIeecSm/ggLuAKXhs3n+HuBT1gy7few7BUBSXhXWhHZ0HjW5qa+4
ZDAPXtlLS4FKF49/HobRZWn2YdQMnskq7Jx2JvWXfyxtxo9MOqPkR8jhpS9F
6xvxmwG9+vesSCb12QCZBH9LfyTmtNLbV1jLf07gFofSaixQBJ26VGBMEUhQ
dfR2pZOFKvsh4Yb3+Qp1UiUG9xA8lKuem/m+Cy4ObV+3UEp6vECfaW+6rs0S
zj81C6qWfGSpZa5zNVxwXWvZvo07mVc82xyifUocKViJSruy/YISW5yUpSJf
EBk7Thp2B6A3HMwtni5hWGmS6DG60tMPO2tY7ALrQr1v6uzUNgvzDNyUj75q
0yu9gv6UG8C+HCzXdzgZqWn2VlscJPZrN2Lr+58F0KOZqFAch0LqbqmWM4Ag
1NNjGGDLvyIlvgr+QvLdIfbYNTTx0wTTUKOzL0NYSfcpt/aT6HMDFWwnwxe1
iDqJCSoCrl1IhWXnYPsrrRHJkvh6kijLAJoGzRPSEbYVfFZghkCsAZ9/NrWA
YvVau8Cn6s+e/WHpn2DBtUXTXio7LGlTS5IwCC/eXB0YISphTykGrvvns0XS
YWrB9Wrov9ekyhxZGjdg35WYQNIS5n8+EIhjaiBlncuSb7FBrdwEiShtu/Ji
UKbi48vrWhuDwQaBdekOefbApqzKV1B21oCL7ZHKGnvnCxmylHPZea4VdbKO
OiIrQZXOO2K6LvWDvgcKHtC+63VHHbboyLBscCLUsaNI7Mf0cQIV/3oY7tQy
W7oc7AbR2NWATuFDUoi3ptF78LmfingPSjAYOliOXTOe5X5HLpDqRXthuYEy
2HWutOY8o4fuBWNRdDwf7VhH+nexC3U2shci3ZDcnyX0F0Kpc7Ex85l9mdGf
ASadFdwOgr50DmhrHpIriiesegGxx7JFh7s5ylfV7eBJflRGSCiyYngHVnxs
NTbtHt5yR2bFzVeFuMK9YimjyXtRx/CPF/LGNEzkLSOMoT7eC6EnTW9ZJHVW
gLsDBUEvlmLiF3TUw82kUpMjpC6yYsUgyrgSj4rUxcR5m4qxNYPjieifCdpk
TApFrcTfEuxzoYXf9rRMTmCNa5aSdGYWoaAosCnuzjpmJ4FTdAmgiol+c1tH
UvlriswrQ+SjD1YdqTq3wB5LLg1SwKt/l2KSECMK5yyzEfHffmh2eJ2JAFDM
iksP8TENFG6QgLMbGRdusSQBN2+WY/0u4MGgOzBmPEcztRzEuQ6DJEfBi2lp
hVfrFrTSmCYZ7guSs9P6wzP8e37FnBsRoFJn9EZH7Hu4jZMoh8pxlURB77A7
7fC/Q1SROSKkBECedEIn7PGFpudcxqGjvtq/1X/E3wXNf+IbN4uRwHIseoaI
W/InRy04oucs9eHORuv+o+GA/AgKRDff0nZMlU2XIdKXtY+tfN/1qNxD32/s
jyLxrt1gFFGR894+kSJ8KlFs7iyekptX/kSI2C+Re8fkQf27ws3ho93NoCig
b4u9rFHJTx91UhSG2wpQ/dB3IjmryTKB5oe6pIIFiVS2oqP055o1Vl3QSGma
Iw5O5BV04unM3eFNugFqR+7HoTpcXp6fbbSpZ8+NwP9tZLSEhG2nsq2ekaWM
nRjXdqVSaIsnjuehdpMnlfdjNQSAJ1QRatvYH48dCqxYDLPzNja0v2n98w0a
U1tIlCPXQdD+QAOuBqWTgupcqkT+ZC04GA56xqW5ufaPX0mAszrvmUFelbSA
nrFBZCE9RwV7RfEbgmH0fQPJxbsEr2yq6IBlvlN+YG5ENwYrnis8aPRGWZ9W
HXyk/r/w5kwjEqnDn1ABq/gKpvClZuN8Nnl3Q0/Z8FbTi3XH7jMn7b7x4vk7
3kvRzu9BRR17Q39gFdiGI0mfML/7MzMDTIlkQsFkxqD6tAsPSuD/Vlz10H8f
7GbtFGzcb1E7EwnikTK3oFwIwo7UqOAPI0CKEeJWSwD/WNbolOw4xEQLNHmb
dBwEryHhKSTt5y/zeIi5PAteQMf9CsyoX4N0nn6jePY0BRfd0ZZJas3Bb6CX
4eeyR1ybJ4hsWwk9d7CCBfF4bsdZlHRU2f4V1Y9ShC5XsLz/HR7WwNclx2Ej
3s7Y/8VdP3/6trfiUkPoHSIIQuJCK2OCrDkbEZQeyB7mnI+c8KikDuP4hcSo
9VMyZjcu+V/C4mgyF9vogwssdZqalsdJlUeS6wUvsTd7nsOjiLlB5onu32o5
x+qY07dYDiNIYB0AfCJGd1cv1HHnv4wFOfmFaR+iLyE+NjJ3sbm2i9n4J1EM
z3DthO0/R6Awcwjnp5E//U/P96lD1owo/rieaV3/5zolgqXX9Uylj45+aGEl
bBB/dLpuj4oVXtpkFWIg4+htk48z8k0YL3EqtzLZjRVc1jpdyHx3wik1whAn
dw1uznViD3sbxD/w7Oqe2bFyDjPdAo3w2/l5pfnq8haNaPZLZmq+G+TqFEAJ
ZRUBvholsfpoqpArWwVgm6ptmhIf18SNSi28+pjf5IQu6RKMtMcbaCWfS1vA
5ycKYXNmOWqyzzBivZ66UGj0XAUn9SNRhfzbT9noMz67k/cNNxL8E6X4T18s
Nkvag8MXih/FiCkj/2LkKIX4ID1kXsaeJkB9S4J8FIJYBWfZ7m7A4pL1GTxj
6D6d2g9EFS1/MvISzDDGNMb2ZP3TX/tZDpFPOBk+VkBA4L4B3wTKTn4OHCXJ
OShKcpx2jAKYYdNJggQZOiueBxtfzBlZDrQZuX4k9G5YkbsiluYb2QfZC/4A
THtztReycivI+G39iQzQ297JjrBDQF6E9GBlCQRGka6rT5es9bE/aoIJmvwA
wjbdKVbR/lRQLsP3NY/6EMePRmjNct9wnP/vsI5gSBuVSJBv0OepAoIXHnpz
axyzlvnf98Zlg5zVq2C3O78NjXDZk5nZiReqS6VMOdL3HzGGWPnVthQ1hfLY
DCw6Irl7CWKMRRzVodglgxvFYjVtznzfxWOg6/nre1ls6hySHmOmtxHZyOgQ
XPTv5d0g8rFMMrCYxIXmpk8K+ZWYOnRAp3KDiJ9vu/rBYXks6AlR/5GCvkg7
sf6o/3Mtu38w7/FylSxMEEGpuWn+EM0CPekKN+eeWsfay5tHaLEmVvPpwGvr
Yd1526xm+rcSSRQNc9077fKl9zw9dci0ogbLU2WdpL6yovbOvu4G9lkIs+mV
Du+kXkqhljh9BfzY7Pvn68v3MELVaSn0IhmtArWgPuejJ+ly7CE6OCIVI/CC
BoswC+UI4yKSj6k+04bJCDwHqEk28ZHftRB5d9cE/C4KuKdtHWQmWWVNefl4
hSbMU+aCsygMMahDBynTnSHsrdR9WRnJLYYZbLvI6gbPt49CeFKqL0XXW6Ct
tYi1180A44JUQxLx7VOBwD7ZqqnU1SwHxbLNKV9g/PRNhb1hY8LNgsYExJDm
ruNmQAg+RAeP3eZSnyIr830OGRMNHneIbqB/NcUTF5XWDRAt1vEt795bVgHl
ubc4f3qVA4P4JpGdqat/w+kJdty5933eiarFhrxsr2YCuGRHV7QqSGw39lRp
EYTrbiU2dRDlh3KkZ3iiH40qcOLPI30TJeXSOcOcpkpRfxbKT7tZGcTWX1DU
zEV5e9D+YCtpFKKlnYuJsCdevhJaWFdsH+hF87mKFtW0rOZpSmMDkkp6mo8k
EQACHgmM7oW8VsTudCE4cZ3HpO1b3MITYf2BdGuXKsFE7eImYSw5M8L7eeUZ
7tyEeVes79xrO76wWBTR6UBVUTAL9Fw9X46CGvnSB0EJMb3td6SWkdqy2sWw
PVupV4bQaE9ZLWjV0+IUzqPlOxp7HeSGdZ1OZZyxzUpAYbL9wZB87u+qaIof
U9HX88ove6/ueuSKy5kehcpoEJW5puHc+8V31HpzJrzRSupodJzejdD57PYE
yMxLrRYELOVuKwnOjFa67wVntYEHhXe9a4B5Nb7m3tjH4sGbMe20nJVy1y0f
A4HorEUl7cUv/FPK/xdbkAS8h3grPz7djkqbyAq950OR2L5flUOoDdbRCrGl
uSU7tlyYz8w5/VQ3yFw71cpm2aslye4e58vICD0VGbn1Eswn9IWaG3oacwO4
dMXxMSxR6nxR5FtPF5WiqGjB5bm1UvNrRMToQMyAyfNTBpnR0ZG/pmuvnftZ
yPQVUsc3gwlvzJWSLAD0/vUVODBLNcb10vFdJnGHWe13qqxQMjAiKSVlGRYr
VBX1KxkLNPaq5oU7oVSOC4H9svH2T3625KzzcFtecDSmHtkYFNr5tXKpLb87
PPw3MufCpO44DDRbyRaSv2L4r3jsIlcFQYtt6ksQZnMAlXBDk1fC9fCFwxnj
YkXWahKbCpfy53+r/AfolYZhXmz4SoUhM2Y88KEEZxvaa+BuX8ZaV1KUQ39/
bDIM+ZQEGbO2GT0gCxNPzfju9IkilJwudYWY2cyxaItSfIL65OINZzffSrDo
/fg8VZed6U/u7fikFE+mhKKXCSLb4MXnhPOlQ54iaoG4x4O+aozUmO0eRydz
OzXv7AF6ZOAn58IwlWkdFZg4I6Gsj91fPilyxFzHUm3d5EGh2AJgLybdjGvk
YYo2XseT2zAa6Rh/sh0r5YIGKjhCA5l5zl0sVpFzvvWlxazOw+O2Jp0gLRa1
BVIWq4TghtDwDUMV3NXGrUDO6ErWlcbn9hNvIRk7EzB07sNMNW7zFL466OZL
koMBCHguhcP+prZEeaCFNDDHey2HOfSd7+oY2mgP25YTFf4fVKVxv1cXFZX9
xzRtUZqulyi/5gFP7Wi2eYuqQlt/yR8f/aXUpnBM3+1rf+wtmAYk0++zwEb0
FULD+mIr20WbgkzBb2AYYVPkRbhxxJBxKyzpMk6NYCqDzP5r1P2zVJgF1Oxf
HmMIJLw4yrLeFWFktLcuxyX0s2ccoSLcbLqHBev0ntwaGVsy1R+qf0Sc+s0E
nisx9iTYwYt3F6BY1YMy8EYy/M0r9xdavaIUCLZflDCAwIplLyjNERVL5/i4
Mda3/4yGQDoSXOAR7hNBzK2wQfB4Tqir2e+xwI1WonzcaX+NC9sfSKpB3erD
YcV1cwK9yLTWSReY/UhYKt6V7rK4V9jFV7154rhYcESPkRSvgdlRffbN0iy5
4Ea3TqSoWZW5Dq44UHCGZ7urkrnDDYlArMLPNNjB7wgeXsg07XWRuwgwWjIJ
AmzmZ/904CwaruLfmH5iq+Tq4TTcusdyjXTXJpyzTJU02/StdR1Kx+9TfqwG
m0bqYD+nSJz/tiYwr3/QA5huB1KX/d13ERzam/2W3fdCK/af9eMi65VM3zwa
gUaumR04aHKijZxUlnuweqv1BvLsPUcYDmWrVnc0+EAupb4QRAaKH5LXXlrS
3IU/H6gHHij6rI14CKVfk/g/eVL9pG/FJEfgdwTouF4n+jY+SZQOCUg5IR39
XDZ5FY2IRu7uHhdQDC3oRd74pzh5eubswsRhNlm/3E+dfvln2d1HDA9gj2oQ
CLNM8WSfAee/NRr1Qmpx6jhZbLCufJmeForCO6IhqXiI+8ApGFBQaaCOvZtV
m+2LSGj69itq6cH6xd1HHeGfasSUMtCf8lB6+/n8bcgr3Uk8hm1LY6n7qDeF
56Y2S8EOueSZ59PUPMSwULEfHHC0qfAhsgdv2PSADxOXTqqIQKybNyO6vf33
a4jNpqjpvPuAX3YmGMcE4FP4IYJ5DdmK+lbfKQM4b/HbW8X9uxRqyg38sP+6
nhS17Rj42cJA2kLWYuE26t5wwBdQrGZ7WFWjYsB0PRNESrqPLGMw0OCBWtBA
ijgRIgA/XXaWHIVacp0L5KjhO47wezQBv2ZTYm43u8dmIWqjiCTHghTQ0v1o
0VyFaesSbqhkRFj5uydKlykDmZ8Mo/9NPAzRodSszWHs1TiEjfRmY7A81T+e
buasv3d/JUxw5HuABKfGGW0k3kAVJggzbeyT3zwhXn0eFeU1+GmztrHW3oni
oHb7hGmcQikfk8Mj/TVk0p/VQYqeOxawttDSe3H7iQQQrVbF/vY9i6C8nkvY
L9caxLs6cORVrABJDqt65YvdR8ins1IB5XXgkV51b/mkgtum7tv1GlpcgYKj
TxjrkZB+Q21PEBlRvwLcFcyr22yzYzRFyxAXxy2tkKdcR+P6YWQYW1Dg3b6A
G64k/Ebje/1UMyzcRKWOtp/t2lPa+2Rk7IL/TlnsbWirahh8ZLszdIrfJQbj
utLNnqXFNOEJcM0+QyOnRhK4jOaWqG8q7MSbDe2CvJtO95F4hxH2V0BvGeDf
OIbaPibBmNI7nvvS5+0P/jndpi23lzAjP+EGXaXAlCxtBNT2odsO/wVzvlDs
KASABywRoiYactM5y+55yUL4aRj14B4tqsgYTaoC/kaRVYZ6Dpq+xYf/fbOI
A1gcVGhrYx70dGjYhaK4RtvLsAZAijBu5i9vaztIKe7dA9gf0E14mYccqn7t
gE1qtrtI/ncqqs9LIJGupKTTyOVIbVcQx/R2DH4Eunq1n+3Nfhk6t6YO21DV
o1KUbHUMl4CoO/BBrJmsqk2p7pwpS9Ay2sOZnLzOEbYOtYhUyRp0uMY53zrW
Qi0VtLi4ofZzHuCT59aogshU7Yva8VhZpvo/NQw5qTupZTRZmwR7BBGtgVQq
II5B2wHal8rgf5APFW1JzhaR+iDTaZSTP0zigrA9wfCMFsLiWEZnfPsJMNQV
JdZFWsNuH4frgU7Ajt7ZzUourhZ6DDIEXhcAnmwMDjvfQOK7ADvajfHZ3uZ7
9WDnAD1HJfQvN3oOC67tIPDq1CiYeVjVKXmVYVIEU5h0m10DUHtG6Ex/7nMd
N129pD9bo7zb/oIA99kS9KstLdapi2YpyKWQKij9WrFPIalhg2zLJRc1sJq1
Ryj3NzABqym0sUhNVe5nzz6e2IYiTHIwPsuCJ1z46e9vthGZen0HLWEJPRP2
Ho8HHpXUoz8I+oAlB3qwPIED96QTV3eQHOfx7NCivpS8DY0xTObaVb6L00sp
FMePTBktoNDU0sPWZVrVZZCv26wO0dqYy2M60RzzXokv+4DpQgCRjA01GZ1D
4y1Efp3P7h0H2+rjyxWcXvASvI0lJE/kANWIXwhP7ZaEYKjKRPtH1qq2psLM
OMy3h3jutpdW9m3Yl6OFajRy8Vcqa1empKcehZ4I4VN1frihESdRmtkrpu2W
b8TJHL2qHmrJQ724WOq5Tu5todpA8k8XR9WNL5qBVDhQ46FFOn4w/8mAJdrc
beqnRDMmZV3vbXy1/JY3Q/iPsFHDffg9M4suEcRdHK3pJulCasJvzAqc35C8
W9ovU+Ko1IJfBOhDzyUUxV50qFas3WcMBd7HxXxWMJRzp1f3wB3dx5wcIizb
LDoK5tRHjssypA501Z8ZsdOOcERiWhbsu4QjR75PJ/NgAm8Vbzv/JOVMJU38
hH0h6zrmpY2x7a4xBh/Fl4q7sSpp8tCGiuzeubLgMYy/lNVuASenLbcdpYUZ
F2wsneylUN2XAe6h7EycSytuNQXFE3Mgt9A1KyNe3Onpdp1Wj3/e4hV60lC7
tTjymiblc4FH3MzE6Ookzb15o1LM2HbYwMHpZCa9bsZmRvq0oh1IYCHlyY4o
yTQlSVNGDNOYeWTYf7YABL61g/nO5DY2PEo59z3dkj1BlCGumGv1w2rv8tFm
JBIz5+bdBXBdolv33DIIH/X1mGYCQygmwtHqV8DKO+osLdVoOFz2RZ3dPdSs
Wq+CZzgKZmaqBfoG7qAlTiJ4GAwrZ0rQd3/D8Q3NxT2ei3528VkucV7afNFE
ZCsIM+UVPoanuECYvAQGwCvQdthvk4CAF7FFkeAwyOTgZYxzn5EipZolEigz
E+KFrS1hZIKeQ7a7B1CIxiJzPhVp8Wau57Gq8DhM//6E4/w+q32a/YQaUSet
NeEvW/xw7+N55/WxrTAOQGVr+0z8S9KlzYgacgkyi47h2H27X51vpm7qbDEo
EhJgNjt/L3A59tefjY43ELVq8hpWUmvnKB02suh3CX/CMO57X035dwF0Iv0r
VOhzwPD12pB22cJgUxxA8FOOkvJR2sBWCeuSaz6cypceiab6oYzPFH0N9pJL
luR+LXign6ul6impMviQu9ByQo+Z18RCKYc+tOYcV6ftdyFhoHhBXAvqBo+6
0GZB87bmFUG+VfFYcMqv8MnsJY2oYXeYkadn3/BpRvpp9gPN9rAz+lXXs2qP
SHnYlSctyB+enZldbsro36hVNE292UzdofYtua/AtK++txS56SRyE+5dtID5
31/i4q9DE44J8v6P50lp3y0e8KqJT2nBgDsbaLg60r9EILAOSicP46AHDfPU
HidmPQTQHUyH0mQrVfyTb0Aro0NBv4gKzWypwu+8MEAt36Plk2fomWnJFfJe
dimz9P/ihHwPElKClafSuSkUPMcgMDCz628dfkvMfnIZVDUrd4FjkYoTYEh4
Ry9YzFvp5pxNtW5BJxxx+aecd5V3guEduUJAwmRqxaOH1zSa/pCslXoJyBkY
T+H3jE4/av1XULaX/egUY9cvbcU4AxWfnCYoOUHheIQwnCTT5rD89X6mimNe
WarxBKG+6PtLN/+z8YRdpWwKh34c298F03LbkAo3er22hKiLd/rDK3REI9zS
NQy6iZ6T1PQ56wc7X7aql6E9OqyWeD8/ZfAwkZn7fxNOMJKMnFvJziyPSySM
rMsbzkj7taZJqBXw9qw7RKneXGxgCoZOHpobugq8XMydbEgO0lM/PTifqteu
j10TxLESDryb0go7OrxL88SzEgph0Vd3cwTMDvif0LAYJeWWjv936FUMX9qp
MPEHDYJeVqsKLjXBiHmGZOkHvBaa0P19JkLpY0lnzgXJM258G3QnrgVi2TuC
B9kbOksbCXwofjyCUFi9gg2xSkYW/TQwRaLCtz+L5cBvwCVxgjYBvo4NO6yR
LVRu1Y0nLSpm+MRRGTB5okRBZQOADM5Ji04igvwL1kEpKoKs48DKHSCLqdOK
3RZjaaQmbbOiKMaaK8ms2opPiy8zeUqQAV/zbhSWkgnYKftjOfalf4YyXde3
Gfqn/ZYh1Fr1VumTdNEtByfLQNdVaeTbyeP0bn+8sUg9xvJoaaXjP6Aufi7b
CTG3jVyhcFb8nojUoXKcQP27YhZoK2wdmijhWZmT2TNp2DIrOyPJls3SVODM
PXaTze4whOfNtHxkO6k0ru9POypeH2Po9wxtTHsFfl9joasWepeNKOgDzD/Z
21m2FY13ttyz1tsbbJPJgo6NglNU/o2QOTuCZTeWrKD0KbMgQ36P4Bu3r6no
PmAPbYm8AqsoJ3zrB7ipQn1Xvu8rr4IMEZ4VECkMaARP9noQuiWdxvKuvSd5
5aIqSJFO/zwnmoux5PutGRVPHDDIbU6kSgS3dxTZPeZUk01weU0qAixs8L2V
qA7fLEqe1jBH21RxrMa+4hZ8lE56CO7h51Ys+Fp9nO4ogWZZ18zlbO0GI0VU
kh8b0mx3CREp1JUG5m8RoskwGclbLAGlOT8lzw9C8cNxotWAupPn5LztoxQJ
aJHkCsk61L8IN4lc+6jZh6RwDzGU7SgEmaAwLh6hNZCBKBQS2R1dgyINyp+R
HORKFnrITjADbwYVOA01s/WrwVknzxw39qKFr6KhTZIlUhM0k7Gyv4C7ZojY
rNY5tM8W9Rb3Y3lJ6VYBFY63mTYMWk6LQxgpRB6Q/XnoEB41v5bJRn0JY3zr
yzxhNU7BO9W5/iMafFVhq+gTkLxDTJlSPbS/fLLsuhJmQBdo8NnOhxq95qR1
nANT9ctcJNpSTLW+Jbf34Q6e8klrE+INVOt1etmWwcSziC7IH2pXot6CZg4a
D2wQcYTVanFuGdn58x1bR6wW7pepzq4MNAJ+6/Srif4ScIvZUb8eDx0sLuCD
mQz/3BHh2HS46JHAkF2w22A7QGe/+zfASR/FgX14slDFL3E2RBj5Tywzm72L
g+mRmCRUsu93KM/stlos7yKWzCSpF58IXnuFBSglSgh+NY+/6V4vvh72eXi2
wT44KM9ELpvZYoK40l8zyRdfAIGr+0WurhmPh5covPRwylqX6MEs6vywlx9u
LBhPtnFh44W28QjG/XHB11x9BjNZPgWVacmGRE7PfA0/LIVfZgP2evn3Ntu8
QKe3vf+a8JoOJwPBjT+XqE4ZIN/HvLuzyU1kxcLunno+D5WCciVLQkGv2nQ0
qCLpXl5SRenTFkXfvMohNmRxG5/2g10rDAKZNoWdbidz0KwY9pEqc32Lim/1
m6J36lRhvANE4yV5MrVFJMf9oj5YKQArG+I/5R8/0zSDhcBwHc0leHjryvZH
7bS6RNYuY4hfmFzUv5pLhypGXIzlHN+cmpX4DXbPdVlcv5rzAVe3G6g2hDUc
jrLcZEd/VeCpCd/S6sVogDzw3dvYfJIv8lYmLMiTmCxbZ8Y0dsb3fyhMgDFK
LeRwTME5eS4c979nP2+Rd7MqYpxPBXKWfMtyUVaQR0Gp/i44BwbGrB6bohWl
Z2ca//gnGC/6id58QSFab5UwJPNuPfe+19itvTWKjlv9ZhwJGQMqoXL1wPQB
f7kp/xQnnkopH73F+fAdzof6LSWyPI+aD9IohFdkfePqjsAgBBGusNFi+LLC
EY4bSwnFLOPMcjT2UDYNnERmRLN7AOgH6aq4oiJbhk4FA34SGgU+hBTX6ryX
HULY4o2hOLubDpTNmxKBoqkpCl5sON2C1UbIOQnx2/FX+/zvYqGr0xXgxCYg
XsNxAHE8ffgucYRKOTKUDuJcaEMi6QqXOMqbemsi4Nlx6sYt7EfVISPFSXsa
baJPY12ZVePP9bYbI89d7SZfOYoWqb0reKEiXW3dwen3lOaj3kq6NkVxVcOJ
burCDDPzR8oJmqmWvQkX/yJZZzw3L+Lh8tW6FrPVaU1/N4OHGkUdMG/5woh/
pnJclo8AY3nF1Ebb/lZnMZOoS00iSY/e+cNo3cG3ib0st9CGX4sT2EoCQxOK
OYW37B/LN7B/wnsGWiSVM1kwVJiP4wI8dUUUCibxMFTWwVjGEeC3oGoJLLxu
/DHhwzcDef+7iCT72MggKxoMzZDaN32eLn+nqYeHyoA/LD5N2rOpgGT11YIH
VI/JZiUJsUOObfx7NZQ4LgW7DLbRxYO3znEVW6OCittdQ4CEdm5fuh7eiaGH
P7wh0mMF3PfyUDhoN2JJr1cN+WrTLTm3zIK+qLX0UrVFQJbdNF7DqFzCJqv9
ogi0fxhc3HYpi75A3mKO0C5kiVQthtqsXpw49ooE6T+7WI4mIasFONfmXR16
/+y0Xa6ohnIaPcGq6Y+L/zY9jLntjbt2iGjjCu84kz9sSLQFUC3mXTjfTV3Z
ThdEAzEIncCo6kqhNjbU6sOS3TXVcxmaZ6a+wk+kX2lGGi60HkjEdi5e1bJw
rNyr5xTLvfy0gYoCR4Ib74xSv1o3obl41AbN/CfuHpHiRlHheboBDGcGhZd0
55+Kmtx6WTg8azly2hQFG3/GWAloe5qOARrUtoui2J0mnm+TS+vI18zpBcl6
L+VvQnzADN6+ljyPiLnwZFqP6RcWT+sGbDjt7pRczDyePZ7rn0+k/AzcxcHJ
zK7305lnjRUaz0os7KoHoNdFvZfW5/rvmik/SY29olAAUA9YblrGiF/0uT6r
i/uk4e22C9IKfQA2f1775iNrSdyYiZfddeXnUTelp2xcGLOTFsgFjN4hhO/G
hjZy66k3vwUqifj/QumnkccZyLCbSVuXL3oMwkWdfkUdueob4jPAtzXHsXOY
oZpJoK5CmkeD5NX4xBkxQX8x3vPWWGOTHy3bxR/Bm8PCQvpg1qif45s0wxb4
mNfrvYYaQ2kjGfTfmFy7d4adj2U1pPJ1sZXtlBcUnsPKLc84/7OOlFErC1Ob
niqIXcP+LifjQzDbkvxC3cTsDiCfX7Fjl4iIp3gooHU2SadfZO9nzEo3Xgan
FjslruQv1acSjeqosCPh9wcT2CAKQAbemztj3ooIKzq+AQz8gx73r+JeQkfy
ap3BXkh7rV9HJdjJrbEGGcxbJwsk18duORWQAsq8eqW0iN+M2wB1mTQhqJWC
PPB31imSNQDWh+U/wlpGfjphs20sJuMB5N0ydflbyF0FDj9dGI/sBGEj7we2
gBzGoSJA8CEVUPmi6wn3VRwyoFEXuw4VFcfnmaeIbxu+QD6bYvgeFR5yjrN0
E3KwaMcYYVCWOA2HsnbU+2jjdZyLuX/yo65cbSgijsHCrGfjX2KheDHjfMdO
nZ5CrBFouJzXMHtkqTMJxJa+rduPPpgr4eAC6mpw2OeZ2P1KZzGS2PMvdOKp
5gNLowr2ZnvDqXAZB8P+HpLp+clEI7GzM44gIfx3X7N+MhwgAh8onHe8onZe
vEhLCTk6OAL3KY605zgRhmzMTbDTPEvIB/eNxbv58eJbLYh6s4znrAxiPn5+
8Ymyvi8LuoVWTTqGu1e678Wz2PuQ0GX4YmM0Ak02+mN936Mq1klClAROTRmb
IycZ6viwdVqUqM0IxaWtUjr3t88ArI2MXgzLBQFDUEQK84aBzGRO5UqQAeZz
0RrTcIiFrJy/ve5HOBqKjXjQm3Fa6lv52cOl5MgmDnUNgdYeFWsfvh7hwWTJ
D+Nsmm6iLDdtpTTYuPiy4qDNZXRdYGZagZTv4cgD09sMrkVyCrXbIU6KJSzY
kDH/u3e5RBLVuc+3vy+Lx1gJxlh5kpnb8pFVkc0teuEbq3rGsrV7ubRY9Fax
3zeGBaCOYA2Vdq2Jpl6nS5/oO1/S9zRQT2qgCJ0f2HUVKd007xvFwntjxCnC
vyl9mFME1rIIE9PipyarmIy7RxvqjseB/ZJDF4DmnBmXU1zLnpTc9ltdstFU
Fmm8A+H6CC7JZBhRdv7OZ+yAqIKTeo/5TyuhJp0r9VPlPJ8vlCElFS2rg5OR
xVpZH1hUPWXy6RQqLEOtZ3ioUbE6KlhAPKE1jb5EYzSUPprzF/07MfrYCPxK
r6DYR55+1sMw/BrRULmrzFKgvLFeLybyU0XrIDC71CWUHvL/G7CCDm9Scln/
9/Cln8Z/zYtOnGqS2EYqSHYcusXxmGZ0qL3ui2sn4a96xJzCwbDVKN9fL7n1
8bwfjUkPpIXQRgrB0D1IZ1BuV1TcyQ6kx0UwFhgHenPB6oojlEcxtNsh4H9L
9ykP8YKuJ1OaFVBxj4Ds08SrUdbwQKOMEsB5p7zkOzYsv9LtkLvCfffW0S5n
M1tM7Nt4zmqdJdP+DhUHvTAQAXATL1lbjscY0gPhQFiYPgSS86lGtE7tw0qU
sX7CthxNrxmqVrLie3eZxtdygf+Ik4zOgLoEogluM72b5jNDf2mb3xjAxLpi
yHZAvuSEMb+N8hE1QsI5pSVphW4wroQn8Kbp93odBZZFWAaAODXRyor/zaLK
jVZMlj50zRHE4zuyCG+y5EfiisMX6i/p+k4b38R8EaXa6SDGezo/3jvjxdHq
caBtW4a2zqYHJxsg+LCNOGB5pyxaPPO3wI6EpWzToWZmZrAGr1HGwJMepegS
JVRl9poEr14us7C5s5JVm0s58WysRrIR/4beVIRAmMJ8ubQZcmIYjb1OLwkp
HSKXubXLssVjTZ+4iJtzVDK5HNZnEAtkPhVn8weAJU4qUN741zqlqM4ewZlK
vFl5dsLrvfCLfv0OHaVH4OYylXitmLZ4xyswScNrCkwk5QxcEVlwU9AuNtdM
yuEvUOaOcVv3qKhSXIM0nswC9EZ53Mfi21pp2bXQh89cVOK3wL1HG+ate42P
MLhHwJtCPeyw7qXm2aZx/LKZTYQ6GP3VDht5KyBmqLK6xT7kWjFbaS7Q+d2P
/onxqnojiFi2acalhMvISMaqeGy6VH4HdbsJ71wHOYhsgc6Lu7FDwcHvEyO+
PEf7KzJZWUin+Kss9JUQBxzDGU7p2T1Vxy8j++xmuXF7bay6r13vgpKl1z50
uWIPdT+n/AIdh9lfEp/4wkoezNqzwlGYkbDSflMDM74ax66cy/Liy/WbzL8c
ozayizvulsfDbcL63sU1YbQQlXe8FLFmWreCmjCIA+X2al/FShSZTnVxyh4L
tBpEixNgsbu842mGwsdUumlBWIi7Nh0Z6ue65qv/uMPoFPyBhfWXSBEYw3en
AAfXasTNMwYxS0Jos+2uR/qqr3uerSvhqt2qTKXpAK6RdOzAK7x0RqGw15X6
PuE5EwhghW7bsSm6+1+5u2vYdn5LCXM4BvkAyk64D8NpBioeMahMF91KigYQ
V2M6EZuirPXDvHiZ5MoXJlBJliyW4bg4yaS5ntkisidX8GGMm1ZUGopYt8ey
XqGkSsTLQTzIgaswwQAyL4gakAJUlilFcjV80Z1mT9oCk7Gcpla1eD3gpg5M
O38hHPuGiGtPDlTOyHMgpLXNEYxs0xUkdLpeQv99G1RVSSyD5PKzZXCKJp6f
/v7csO2Mxc4lLpRX6ZnTOJJ7i8kauAFmwWEgVTZYvXzf2wCT2cnSbfoRK4qX
VHiOE9FwRvfq2dc/atIM9JQUsmsmMPCLCcq2BgMudIgGaH3KcQC6EXmVKEpB
P2TYdrSYLHd1PYqF+DVi8HONh2uPH0I3Y2vOKTsBkk2Ztzbd0o8r4wA6mou5
/XNfge0vgK3KxoMw195iaFyUYVYrWmvv9v0wUHMQLY6oTQNfc+hndj1eic6l
Q8g9GcaJetlRu6YSgXdb3L8wl9xYdEi3Abm59pZlmhTLPxgRYZtgdHXo6u73
o4CavUutNwGJJUCYT+avdOB+7UYIcmahYzDZtNM6i2JMPfHDaP7Zjgp4TN40
oFxBsWCoq1M3yApfbYU1eIeFLE5aBa7KSGUaYzEpQ3/kTGSAt4SqgV05z9/4
0oLYlhSl21b1SA7aNd+Mn+EPOIVUrSp+wKyQZPoPxC/8/DGYmhI9F+NMzJ3B
4uSZ13Um6hMgnC8zjZjWU5mQxw2pyR7uemlpZE8X8HvK8uupvXRx0C1rqc5D
R/LjJcn34FXCAxekdnOeHv41APa5XACgC9fdNOjMLyDuUFNQ1UHFmfd4M/es
J90OaCn/CGV4GkAmRQodSliJM81XD5AaynSy47gmKeuJ0XY1gfz3mWz2L/s0
VLhJDJSVWce7p+10dOEdFVKO5xKJLxmxIUmRaQfKyteDmcf/82aiqlGgrN1Z
Y43PrNtjyn5xyRJ1uUGP1kO/BmGf3ORdK6bgo4LNTAORBD+XYKZRkKQfv8v+
6QT+12azftwnlnmjPGxxWn7BJxwLOMrXVpRSjoKqGZt5WmgHJ978vofWCltE
yWmZQ/qTKGbmD+8wSpNuAhPYTcrQTl9XNouf2T9pUotjnlh/q2TpuHnH/hVN
yYMTltnKT6LtcvMdYRu3YwE0mU20CmH/MY1aaOEKDnShTJkvF5d8DXR8UGSB
S2R1OaUwRSsIdRYK+NNXfxguhfHkPiU7d31hJboSx7kFk8+THUrszP8OkqrR
Wbss7wI9Vr1wRKn8APDuWxhIpIBBb1cyoaBR4xoN17NSmL9/vB4x/PjegIkl
d8jXiybQYG9Js+XdntJrvFjItU/dsOSuGIU4vRhpFIA1L1aAHB1ZZ6n0wpmw
oIhGyFeFuaxSbgL2ZU3uBscH40k/zLmzKXV3Dd3pZK2j00iYYbTEucAY22Vp
/YNlzAzpb6Mhz6Km9wart2tIs6VQ9LnJLPwU9a7NRqtpvewGJmne37lgi2uY
9qkQihQmKjJ6Dc0mqpg0n6jtDAfnQbBjTcg129fD5vYA9lVkYBNy2k96PI7N
eADghn2Bq915t62Yo9tp00Z6YmD9j0SWikHhtj/7zEEyOgODUuSl0kW7PJd0
g9HgUGxnp0G0mUIs2EIIFFdItefNda1JmZ3+G9YqCxs8pJRg3IX1YA/a4pXw
ZC8dZYTmAj2BWzirjelfxZuHdKUhaaxSrzZwk1/wsSWdPZ+R1CDg5cVj89sm
g15BbCfIQmBuqwtzZs04+QrWPUbqDtOCRHr018DRi04mZYAc6ryF5L4JLxQI
Z03xQqNyxsk9Ehwxts+zO9FdGLbwiumcw7AzCvWCSiiQggUq2k8X1yQcbEi2
+ymNxt6Il7AB49kRI7P6PZZ5lBTWf4R+fx6Xz8ceKlmAxCBV5t/8gFN10S7t
+5TCg67X9YPOsuW1F1WuicIla6VHLCnJW2e3IrVcwyowG6wnWdCD5j4tWBtY
i+Jv8xzTqTKU5PG+lMV+HkZNTlfrctiT7XWYu9GgByJPz3Ve7qZkIBnrytCG
gF4JeCUJNybwgIfMDJFF0SQ4VmtOAXuRM+7y9kOhChWzT6H5yNO+NLeOzazk
TH2fnvZg9VHrdXOUwOZpPh/Z3hNDtacANUYZzvgAu+6/BDezEUB2pJuej6iI
RB2YdjLSUQpzt5K0wVI3/FirBfLVO0iEZtd6+WbTfCvDszn/HiOYv+6MVM/9
rHy1XhMrqxAiXYyi/OUno+6eqyDp2l3bRDcqqOUswLwsYHobNoT0aUiT4JwH
qOqos+nrCZfXZmLTFC6jAV9K6mIZ6mVJeLwTu4QFo4g+qbrtJR4qnR/r2e7m
7Ap7vQeQCkYoX/8NOKAJB1YyVS3Z/SS+S+Je4J+vBg4E+g+SknAmO3H0U6oW
gKNM/PcZU5knpMp3+YHtZJ0t6nKWtR290altNhNuY7EKjRR370LkRzMAfYuo
hwhj0oQEX1mGgnXyk2GeVknDckPu1mEpf6Dq/N9MbBkzCYB+Fz4n7I/s8rLE
sku3pdyFThkHOhVZXi8BwVZjuuZe6NULqBllWde19ajHQv2ssByVuTuLCDYM
tHvwWiVKUwkrVaM3LOnOZrXaeq9rK2DQ3i5bPoqy1ZoR1R3pP/2n0zqH3iZI
g5ZSdZnigUpN8DyyhoTEh0UG7FqJfVUYfkLCl+OJDQpJor9KDfsImNLwGHh3
TQA7JMe2qswUygKuI7/EF65fbmhwZsfeJRMPHz2RQGelRXjnzj7HCljfjMHb
d91dyuumvlYcRNxjOVPB4Ffx7BPECjanadZaNHnExf8pqiEf/ADGyfU4Z2PJ
1IIQ+r1GjyiZHqSW1PchSkboEBFwxfV86aaixQ48vmBxRiNX43XBifM5t792
+Dbc576ndPsctAQYG0CLjejmxRq+fhR4vOtRZFD+MAi/3GIPLl2YA8BH1nLE
oJgcMMJ6kI2JFicagYG4vhS0qqXadzUzR+qFiY1PuSb7gwoVw+40HyO024z7
AAKqUadnqszDwAeQoWtZKX/fa2XueNkSEOE32VROp8Fl3cm2PI6ZwoXNuHRi
Mzp1zDJaFpxIm7JB8+DgNZ8AZJ+kpCPe7E++cEslRq+51KWA3WeWonVK4HHV
0J+E0sD3+/d/2C9e279/Xe8oX/jAAWI3YImQKLuuP7wo9mZBecRFpLRgRiog
HuT0L4n8mS9XaHYUjyJNqC0JeMNm3aljcNOfpkU5NB6EAVIl85go6EIFhJ6N
k0Axmqhv9WZB/uqYnh9TvCUfmQyb+xZEdz/DwG3wYa4B4jjKjrDSx0w2IvSS
rJNJ8/1dOg0R/RroMXJnqkX7uzq+CvfbRl0hkMPPLtxgAFhHHWI47FypGLr1
K8cM19HNPZMZOg+ZJLqkgrwTTDtf5TW9xV8bhAcec9r/AH51iHWHrszfoL/B
47SEZEvH7IqIFiP3ghHskFMHqUzNwUBWttuedJhuaOFUX967ftb6IErkcUjG
fcmabAmXobgcK6FwG7fT6rHH/HvdoeAIwEH2FG7hv2/lZqiyXVv/eV/7IiX6
C5rN60UQiFpWmaP6Upv5ExGrufDmOFDWaK70s4Rj1RqZhafBR7GeexCMRpB/
hBest/k6641JCtfUFhsIV/v+atvSlglqXy0w3eGr1I2c8vaYZCGzUkb9OEC6
lrX7EOek0pGCkIPI880TDI8MwgMGRWsJ1UlfHVG/SfI55eBxDskkeS9pjY82
L1EfRYhjtm2rTx/tiJRBMQeHASV1kiQ96lIt30VN1InpWkqUFb/arowcea12
OHzOT9/hu6VthuGEdBwNTRQzws6CIr+YVlhSLW3aeHXwR5tHVLdU0wicGdrB
RKkomAFmuPt8zbEWBf+7NuIbTAnFp3whUQFG+0O2cYOKucsuMsrcsWsL9UN4
kPqmDqF8m0b8PUSQ+GMI3qpT1Fmy7lM8SeC3Y7dZZffvqckA1Hval+E36iYZ
R1UmuFGvKDn8Nk1+uUks3IDEQhKDw1lKfFTmOJy1qKeCWDxqBQ1HjR6y+6gP
MhYi5BkZRLOA+9feDPHdiGpUq13z/tnTMQwSkYmqBZWKlG3ztAUDL12vnGdJ
pJAynyrsNOI/59x4kZnw7Spg5RBEIQazCVRh1zsTu0KtLfQ8OU5StXvtffSD
XXkaZl/1fFRxOp8XF5ce8uHaf8pkQVeZt4ib0PY8tTqOnBXBQBXpjl1ihgQS
Y1i7HEEJCG4Y/yRHtAHGiax/9zkBCEEFjNwrIbpkUSpadgu4i0z51UGUg1r+
Ps8h/ua+644NibL8hvBMlHK4jqbFj9wgfECmT5wrXdW/66jwCB/1UgCHDQPG
FqnjuPw/7HLCSEgcDjlU3VACI6g/1RACug1TEl/BEXcA8IzLZi3XgI+e8Q7U
AuBqDLyypUi2zrEcq1FyvtvTkvczLlmKEyiB2tXuYv54Ejh2h+d5WWhVgUy/
cBszwYL56Lq+WyuMYJw5I6pjnPZhP7SDRMSbnBcWcIUQLr+kU4yryWFs6tDH
lh7hQXQV/wz8pS8P2wbW9LskGn+epE2kynRY/TADZAAaULAS3NpvybJy6nSH
TKTkjiZY7U2lP1drzWSqeHRo6BbEQmsJ9jpiwCQu72UJ76hA/QoMjl4LdBJT
foCS5xp/7YCdOQN+0kCwSg98/JgME+mgfs0YvFRlTotGw/BR6iaBdeTNkN+3
YBVQnWUVML96opOzFkMkiBNg6MF2+0Ph/ktcfeEbi02iElOYaj5H0dKRBEYW
r/OkA5/qDcpz8UzQhT39HvSSU1ZBnITB9LnWH127yv5KCOaNHBpn0xijyPKA
5G/zK3fV7El/JZb1cVwhqq/VyQ14nT1jkG77afpwkXsZ14SZiXfo8sPXatKt
YAAkUyR0B3fQZwEfnPJGQ8yTnjvBRKUbUPM7GAs6DlunelBBWPAWTSa7hEYW
sMiA8mtYM625Y4rOJeMRf4qm2b6KLz8glx5kfkAYD7BKLXp2r3IeSWuFM1Q7
OdJ3yGcj00BlkR+c+MrnXuuwFVV16UWRPXVhZO8vpP+LLuLTy65Cnq70Q+eT
1xBu2Ekr9vdFHwtUji7OByp/bxAGfeSx2IpmaNce/AecKhxLJu4yZSRSyX4n
rBKc3VNJ4d3iyqQkmIg1RipZdycvaU3UaZK1fhsYxDBGNb5KPDgYvowuyCn7
7LDffFfauora7ChbWtp9d4rLp1ZD+L21EM+KPk1kcJd/mBzX7xqrkLaHZyVO
06Y284U7rraQMUGOF20xbDLj4RwuBcJt7Sd7jYmZS0TPOQr7I3VfDXIy1mSj
v3dM0qpJnQni1JR56gNWf7xmS2KFC1EjTZPwT4DwBhmemF4QCdUufrUboMou
nIPafW9SaVhMhaIFwoqcRr0nbgiEtcClKNus5mjeaAJK/8xt+lfYMW+UaPMZ
2uwpCCscl9Iivkzl6tPLVtSN5EC9K1SDy3lgqJ/NsGMELHZP3NyQDCoo/gac
PO9Gv6Ad/atHsl9ftlYbjDI+lLujFTR0eXWiQzH5beGEmvcOCTzN0EAY4bMI
h8SPkArlJI6uIg+PEtZPVMu89FV/rXI/FCOMrd1datR2/nv+EwpENhT89+kf
+uAvsB3tG7kzSHoFzZwJThdltIT+6hX1/IuTRtoHES3RosVLLPUJMuVBifKF
Wa/EvxuMwRveqfKb84dU6iusAdt3VC3p6Sa+SSX31cURysDi9IUZKCTuP8Vg
29x1FIDjJC+zXB0pcwLeA36RjcvyhcFb/v/EjBkYKeDdyMdnb44/E4YhUSsT
MMIHWqGApKIt8DKNiktI3Nj1Xlielpej79hsP7mX21H/JUG5TAS8E2anbqzF
EhKzQdHODwIkO4/rLm/1mt84/N2WEzAN42Gy7xCJEOmrNskOdcXL0DkASMQL
wr6BifpPKoQTlou86DpTT/KjZ/5VZ++lE8Y96AYRUgJMt5WW0HMYgq1RA+Fq
CFMMGhX/39GLEMGeBDulyika99B+Ovq7AoCDPoUm+90DvHvO2vIZyFw3QPlu
2rJXiSr7xq+ADAqSesi3W1nIHMjnxGBXIEXLaOekewXp+ry1kzo9bzZfEqY4
MnoP5UMyoe89X/FAMrwQKSY1fqTg9gNNxRNwcBRySaGN07BC5CzBk4HLfWut
lSGUoyreW1OfS3I9UdsHrM2T52CcWI80CEBO9LZFO59ufs2P7HZeIUj9jC/H
cc970m7drES+bOZQTd87+NX4SQYl4RTDAtnbBIx9kfeCyujDYBtjWxneV36Q
EpDGL8EmELUjQbpjLEr25n2OhcL3TuYj2svo84TRkFY0NB9PYJkb5/Fso/Ur
qyw24IaMehKT8Psge/tViO6A7tpn63goFcP9tK6ah+zDuzC9P2iw/bidlwoR
s2aDrYWli+qqJBAencqEhvDHx4zznmyES76JCT7YH+vzb1FWgw0D37tQ9HE9
YbnGmHN9PdwqCb+NI7VmRSjYYGqOf9VpXguSZyeOHT00PJfJGfa9wONGV3yq
ri1EnMWOp06CrfGLeiOq6Y70SSjiOjPDtlY6aVQo9LPAYXv6lg5Jxcj9YYoD
1nUaTLt73BU4A8iMyz3Og9yiT9/mGrm9iHFHlDFqhIrf0kdx7aqCLO+tdpOv
LbFpdXDIxOILMo3IJmZC6V2aFQu0ykQlrHSI7K37LYgv9hWVKMPdadHgn5R9
lNY39ZDPTZwEMoxDFBW/VSKbBkKL+nBOsuqoTaUpFwDH/6fZWQMPdi1X+pT3
Wzynj0pSxW77A6VHbmBrgpTHz67kotodBvjeH2X9mgxa7pkPiSzaqgy+b7F8
8m1vbCzSk6LSJ80zQh1ifKJWPLYNgo+q3J4fyeqPMfTgsxpl+UppVLXjjzVY
+IS93AzJD2/OE/o8ER26SJ14/zPrr/+i97K/KfPb/cHYKwzhy4usaIHCdpK8
ZgZw5TUlQShheN1WjDDmRtIAtL53fbL9pLsIiEWUZ7Hz5N2zOIHrB2ae0v4P
rWyRK8gUAIVY9qBrFvOZsb9Y/xuPFet0/c3AcgCkE9LT/w7jfIXQv41XpFxs
pHzU+ucWETAi702+AeKrilbi3y5MUeD6XiQMeyxl8WoiquHzhm6lEvJyU26f
r/TUywhxCm/v6JoOH9SktIvcedNkUB8rpNmoSexyiMXQjoKFDg9a6rHhgkBj
1LVWc2b3UK0EVjycVRebhbPHCffpdoKZUkgQRR8swKgiO2cZxNfm5szQMCkh
K+sqB7g1QjpVeB9hRsi6JeEd7y2wXNrq/eGUFnTMXzvzXLqyKhEgbvQ0In/Q
8nzJ8O9mX8So74ElATfaLshrMgTF0vt9h9H7rbu1PkWaGH25n5N+RB72EzgB
eoIEZOok2TGLE5GICb0kzZvQwAP2ZCR4/VuKmDzvihVMJzJDQi45nfyKnIFf
x0AA2+P5pF3BMRoDau8J4wIkdvu7FlmmYOt3NccA+KRpLzznfOzBWgDPYWdg
U8TJEEizRFMofWs8M1Wvc1RyQ//6OXYVe/5ZUgA7L9zTrxbu9RJ9n8+DzG2t
ZNLmLk7FAUFZ0FL5VIU4tLAp9zpJ3xw6qTJP3Z7PXFA0+2wa1rv1ighvibfn
BxJs7rl67/zvregKaKKqlDf2L/Hkr49dPUSYbDg2oNDacJC1eYUFhQPHNw40
VqqmXg3LyoQwIlLNF1Mah0/iKfbNsCmzIG0y16Fy5LDWEnjne+4blo1DYWH+
Ka5ZF80ZNjHtdRnkA8ky/5akUzsOfWnrbG6gE3g4JdGoT2ZmsbXG8nKt/ntj
LDDJniErHyupDZSGDytG/pFTBZtNs7WpwaWLwaKPFcFiF4qbo/XzJKa8CmmF
4hEwKdQXsi59pjfRVWCfbHLTJhHmBo4LOkEwGLcnYnHECRFLYkfkgff0u2yn
HvHBLV+7HzrtbDcBSXyzxxm2Nhar+geYXcIZrZTmmcQtJs0pdVaG9w5eqP/2
pok8Lr7Rr0rV7dv8OlllzuBKdYMiN5BGG8yc77b+qAVGTwf4IYz4ZF32nA9L
Gx/kiUK0zCCjEvA0gP4F8oTbwvpv6E7p8HRm80xELxE86KCdaAlOqi/f1Ub0
+61+ob3tSzOiVv3AHWkJWMojvafkIkQzD5kNxEVHRSoWnrARkoC4wny7lvZm
MzJEKmi/vKerbgEam4HVqFfGpCcM6F+72naEgHWTUtG807RrmvB39AMtFDR7
TKImNqHFPFuI/IvDWlYDWHoNvBitbvpg9opi+qjR02CfSgCz4i6aPDo0nDKR
rbXUcRAs4Kmhg4P09jKZbHRdD2XyqQwqW1sHaRNM7w5eqGqI475r6HKcVril
6/3BQ/nncODYhSDkpZ0vjhmwnflXIZ7BnwvIzKmoLbY2F0pZTEcBrjViEEoZ
3A+9jAGGBMz3rMEouyaPCt9CsjvybqPvxnEgSPbOHddvJsJDT/IL9vZyIEHl
ufBWkKhccfR1B34RvTE7qIi2lFfx5uWNYKT7hHIWj75PuTfJiMmu6IJeGIxl
+yquzw3CvyL4nC25+d2FTwj1dBrlB7dg+fGdqBsAGQ0BsulYf/bfmAZ7uXCz
Kc3UYj9qpElFfE2+66OOFjmiVnB7HZ29gjEnWVc+lcwtLdDXXQAzC7T9/nX+
24hj+uumO2gpeXh7Dndd0P62Y+CdClAuTXR3XEjCAORPmJGAi0VHrR4oof5f
Od+v+2vBm0JinB5gqbeL//WBQSATd4XfXtTQ/fnXBJd2vxLEzET3PGdZ2Rqf
vTVhi+qN9G4O2XZ+CqOffS5k91knVz7grMw8ULyCEYuZFedbmDNdXPRANa1H
3KzcuXu814UK6x3lLw76qeRaHx2JFlajxB1vWwIRLOq01KLIvmJ2FLy6uZ8w
wOpSNPakjiIauAEZrijxBM9d/GBeayKH3wlQeT/iO1idTrJ7fbPqHcoswJIS
fS4p7vU+1/4RZUfQwj9B2q3BmEYL8QUoefNc8NJ2JUwGwcrnygERAvasNQU2
Xlq9LXnRzhGKeB5Lk6v9ovcvBPY7yzCjiN3dpi1K42M270ldbJn1JG5/Wq4A
uYF35/l6FGcoQtm93Kh1nXu4EFtFMkEB5FNYXgggwXaXuF+NCNP2l28p12Ms
ajSx67ESL0nFxhJ7i/2sCVEkPjw54n2ICDXGzPVCZSGgX+bqmHmZkTA/Q7O1
0E5sWCfqXfVgWIvsn8eVqdwg6TfQLwnLoHcDESEwG0LvzAnyhJWmAj+3uUOy
h+X3FRcq8fuqrZ98O9giQub+Z12EFeTYzit8i5pKQwPSGDoolXCaV1S2I0sa
F0WXJ0Weg6NyhWnSDYteSHG31+SxBwcoH7HrTCGuxsrAGL7Xs7OJDhw0VU/T
MI+Cr+CQUEww2eWPUDDOvTKkoPJtGecTk+sl9n3WhotkLEiDl41HiKlA4Cvc
/J/2hZNR4qCT9iP2Mapfadv4ShWTkgth2pOl0ryKkKR2Aq0BN8oMrn409LtO
0fd9KMSJtib60DpxLX0CTVN2tX/+3KSsO5qqHdEfX4AaTb1A8343kHTWv67v
q0JEhEdFG/SQ/NqLYLee1aAJympbQioedUMcl7TbnKxxgRGfuJs7aDQmP1M7
UdSQl4Cz+biZRYlLp2HWHi8fI5BrfDaqiUNOMiAUwgYn5Y+72Bn1y46Ava05
PVzpzxrGyJGC2zfnFgsaokiEI/s2EuBQ257t9kxJlIzwhOmAGc+NlgwwpgUT
X5H8SJTyAcRYBk+Sbk63EuOCarhFmN0CRV+wUAyGm/bFKGO3l97d7ImY8pdc
ys/StPj06CVx4x7vwpjbyD5QnxU/Q4zS9j1loqu8JMwZf8LhvFXt1atin2Un
Kgpj7byJxVCZxWkPOhSlHXUCiJ697aPMVHShYwBq0LO7iNpb1k3rSls4EgjC
v+m696sRo9Ox6Lfbj18XRFPYD8/o/jbrZ2LjXjLp4baGAeOwyYFUXYCwsBZ0
UXiBwg01bUScvrC852hfYbtCa0odcGxykspbNjZ56KVRtElZmVnkQRskd5Dv
OI0hEhhrDTAkISxs7jjstqZXuUKLhijg9E3/TW8morPkqlH5Mnq8nn7kVuv/
7fX+HStCmema0iM8sFOsAMiQW+D2Axi9WDywBU3yyLfZScFqO1ziDn+ytogI
MuRfbiY0c4zL0tTuC8KyL1x0UYfL3+QWc4VrpBRbbvI8zoW11xCU6e/X87Iu
NekIsMHo9J2eyQoWWEI0e3hi57ktlok6FfecLF617rtwby7Wiv+tll5dU/tb
VVu6KswXwI5kpfkxPf169RIoUw04ZUup80f6nqAaJhi7lIxJdDTaSJqcOxST
jiLRYuBYKzSr2JU9qBixjCjjuILYXoXRQL1uDiVpadQeC41b/zeCld+LKNP7
cL0lBY+mbyBrVdNscm8yf/IW7ALcRqIkrurEDUlBKAHakhpmYFrI8ksc/nT/
zMOb1D8RF2s0/WCbMlxj7OtfFhtfGrbi6BpwBbvu5lzk6YF8LYq1bQqYxNCD
vdnFJLHLm3bdyI+FuF1fgDEs0kUhklVSIA5rJ2FIDlzgjIOC8v3LeHJyReV+
0BihORLpYl0SoC0iXDesCMz9Uh7whYXrNaVauuo2jYKEhOKWtbFZKWgr79kI
1nPA9KTLx/EhnNoJXaA4cOeczr0eTNKmpQvtPfbFsTiiv+EXXm9YhZpg7q2+
LAkRXYM93uhv+rSqQqLpkAd8kcWABDF4u1YFSwZ1pyYxN8tDW8MJAoIHU7u/
TRiNK0jYY6M312dwfRpkep7ysbMsGQU0Id6ePMz5wPFjt4HEE8QP0EbVHFuQ
9HnS99uMB8N5x6PQHpF70DJy7kwTlhqEeOvv4Cthr4cCnFUIfdMppl208uSk
RgS9+XJ+oPDDvenost4nhglsA+CHoAxI+6HuIeB/BUTo4gr3UI/TyY+t30Ov
QfdfBbTn6XPvUTWd6l1+UXKfSbV6xZnAsJbV96NNB0qNJktXkyqotwhO/A/C
R4aM1elSZ67i1+o3yui9fr/Clp4Vu/6hxmkUR40RwH/tz8zWdpNzbGdSROcL
puIYusztOhrjc7oIIZeoaTTMVl4u9cyD190J9y+C0EUV7AVqVJ9J/SYrbfEm
X3pnUYSJN0K/VRiMO+RlKjhpFPMskChqx+S1Cm1+n63cH9jUcbAkyzoH6W4z
7ZFV/VLpjRflAHpG0OTizsPZXHCI5g6D1zdtFRzBJMp1u+SP5+wh87GPnzuo
sqCzbuCC7ocKEovL//aAbMVNbBWLOUU3kf4WDZsBM/iIvXxLjFQeU3C3v00T
taY8OnXt6OwWIHvQJlRhsikV3S4JAtzY21LU4+CxRjK7DtK6gRwf/LHBv6Rq
fJtX4YLG3iz5J82NPEEDx1kju1Dj20GNHwXcL/x+2rZWV+rGG8g3AmctZ+Ix
eIJ+lL5NDgiXBIahzgvghqv5TM8ovzSzUo22FUqYp9J5Pd0myVhj3y5eJN3A
zCB5yXVt0gyK9tKJGxvu/KkK6rUQpZsX+D2PjfB/oNKnSFAQAf215XirWHhO
QlAGbFcVlOB/eF5oEfa2r6ftFKZnNGYoulNXMERNtYjpPXjqovo4dw4xfoD8
lSsAKm2VuXOieF2icRChb0HlgNDa4jgSQ7+xbbxc97qehs+rh98iSdYl++hu
AHxqq5fM920e64cHenMTM4ZO4Gy2mxHGCvx7/GVd4WoM2eFTrjSAZ/5PZCK8
bc45w8HfU70xYRX3pyFOxhK5L6U6r/983ojIOOtKqquGDFJoDZt3fGVBdbZq
uQM/AkNVeo89H26diV8gD51wE6lTLtU/fyBMz3IM8pFoybwiMYAzH0Vck4x/
3nnc/WS6N2bCb1EW5NnqivT1B3kbZZeHTqQ/bZ95xWZv5ycDzeM1WbVyv4eV
j+06jgdxn44qclgZcDeBANDv7o86jP54IASdCOa8Q0EvOj02jBP13YPBj2Uk
Y5v77kI61ZRG2j4P1msShpIOmKHQ6VUXXO3ZApcCGSIjWqb1+DFTERzi6zRM
t2/hzy65rmK2lHrMacSHzuOHUIQ4sXVkio637+ShDoQ4E62kMdV1fBpmFIF+
walToIxBU5K4TkwdvYSVOymlCQKnZnKOQ+y8KvZNJi81S4x5ETTa50u5nvH2
k7g1GwyxVqo9E8NuZVxu6h0w1GyJtNhIz5toDqaj70f6+vN9ngbulpMohXrj
3KBB5gW7PBM+nJoq/bCXFNwKzXtVVVpLbiqLOvwgWEOn3N7K3HNltRBsZA6x
diRrny3eu8bbj0UK01vEZvNZhPGHIUcPw7BrfAzaPOl1CoGXJLqNy8tzjmHl
92TltIukfGd5F00ISwpUFPRkkCRuuQGKwFlpd7B2Q9gn5/ignDlrFRS960W4
Ng2Dogp4E9ZRVoE84G+YMZqIKQFXoG8FRxz0nYM75s8pdXzHpOBVT7R/PjZu
6q0jpGyXVBwTG9yJCXhU12CqIp705UTSbdc2mTymtTaMjeZEqMi5KSpeWYMC
jdkMClDa8/785jM7AuMoDeb7swzZGvz2jlm7wpBEZSdOXWrWy3R635rwnbBJ
NPnhF0yMD+4JVnPeIONusZqsvET/ZiFlbHn1dlw9cC1CT/thKxbyYNQS0Mvx
pS7ceGkb/4xAHy0+6sPfsDg3VlRkCtJXOyuk1BIb19m03zkheey6K+Y6Auhe
R0tCSkZQnb/6143YMx7AE74Gd6smHgKfUj+HUUhIojK4jFpla70qlsc0iPg7
r6KJgEznWmYBw3D8oZqT1PFLJr5Vo9siZ30DchxQlX6zFj4feO8sayD4whtn
rJTqxr37wY36zEdSFY16650NjbRw3+pBJHzZ1wKc177OntxGRWrAlt8debHQ
yU0Aa55BAmr7cHNCHbot9YnPLXkFs0MtbhUsLZPpubWDJPl5mRsd1msCgNpg
ZmzddYgilCvljRRS8Rp7R7LrhhlLzCg0wpLq/lkcCPT650UqMkv0TsV8O4FX
qzxuwTQaj9dppy8TcpiMHOdkm05Q+9j0klyo53BlcBV+iAgDRezYeMjEOZgY
R6Ky2wE3ilhYKhZzJ+sjmbJDrkxOSnaEna4lzfDatXI9Ovjo7kN5XseSghkQ
3AeByBwRHfO+lRJBg6dpHLNOraioPPH9gbCjdDDzb66mId2bNsWaCuLsO3n3
v+M29J/2Rv/64o96UfeLLy0Hql0DBYsPAd0DuAjEJtH7mBofbFrrz5INcYtC
Y7uoVNZU9K/0PAUeKPkaEoVdNW51eurT4jvJocdWDr8bcpaXN+xPhDlDRf+G
FG+DBIz1okniOJClsfHfR1XhNpBkRff3k3f1/iVys4A83AauqwT2oqijslsM
/7Er5u/OBnjEl/KX/9JZcEKVYwmaIfu9C3uSS0gr/b2zBWX8z0kXRsJW0klE
RDkjKMq2JgxNDDcKqSeDUkBsN2Par+MMd/E9LZ44bP6ajal2mJwGKaR0U6Q8
FwfvF8tyly+uN/qhqr8L0TF8jWefLfYqirly5nn8QX1yN+1WHWAgzOpD7vS8
XndvKxIosgnCm3DkWfZIX3IkH+W7cByHjvNLwcZcr21ivwTQQHDM9pDqoypZ
8VLnMMiMODBaCTQjNiHnBludjJU8LeOadUzQfkBDnvw1hMxuTb7lqjFukH3C
b3sz0/6rQwGgeVqbR9DLkypGHrwZyU1ZIlQvf9Ni41YnPX8EnbBz3qvLsmAz
PyV9c8qi2xAc9Wtz5KGIFezBE7x8K3NJkl4mMAs9FQjmvpNTbdfuIE9ukvm3
77EohQ1nYAcI9R30vzOY1XbZUWtu6kaQDS0xiQvCGfsU8JhnjIaeirpOk67Z
6Ezh05ab6GGArqJaI1NRz5V+q4m99wwzimEBs+aLAfjZVUazZvf2wtO6wAs1
FemZDgMSoC8NOswPYt+H4hEy8PGKRtPPul96lwXS3e3tNlfE0/zuI6jYozks
tu2w7lYIdvOHuJLCbxuaizKqgwcZT5lGorVYSUBDVO8CY0Qxg28Kf2lWiMU1
WB/Jp0vAbkO2+GXSxRN9AgiLBh4SOfc0ROdFQklsJIGxrdK28Iybp5nLBk6+
y4v+enSSczjoPnRa+NYf/V9aZ7lA5nlvSOAQl3kXzJJxHlLALijmPte2IeWI
De6p46hLocNsOftp7bHBF2Zc+u2RWSbUN1E+4x+KLbv4+0nFyBXpr43I+Zl+
hs9zAsAzh3Geq8T45zRXmhIh6WPGHFwz7KRJBa+9zo/QbzEfcxWRiCRzOKGo
AiJFWRj3/fddyhSnK0gY7UxwkazfZSsYWiVKDprZmh91Q/IiFGnsyZyCM0SN
/Fj2TeWcdwb6G6xP1oqblpF+RxgTX4qUdymCii3cETAAPwqDzzfJRhW6W5ne
TG1F22VzMRZvfQ/VpmaTqa1+LQAAkc9EW0I5l9HPMxTIPXKMkeZRXw7RNF3J
0UC3bICSr1jSg76bT6558I8LA4+OQOa6DZ6lkLsl8ba8602F8m7sNloW3gMd
Hp08QuFwhOU6nguobElYCdKsn5p8zMVdmDyQRSFz6x9AjmCziswC6i2oD5ot
OFs5IqeqUmBXLeMdEcG2BD29BcT0j++dR3cZLm43w17noaS7wIvszS7DRObk
X24D8+/lmBRK9++VN5KeTUdMU4nO4WndE4viZWss11BITPhGHwT/LZ134sfU
RKcpOCLmhDjDqzVbFIV75yaMfcYH+Fe8GdF16qekmcjhwZwlqB91swmGWo0h
RypS6+LlMAxfKAZ5cb2a3BCWgl0c7d3zKq96ueeh6bCgrccFBXt7x2RZWo+0
/fCzBlo377Pz4Qhl4QXy8lZpKfunHXWWZh/D/ySdsBFNdbc6b2RGRCV24mWV
FuO1UsS3WvANH9EKoOaGFCqz+G8mLizNZ/5PXE/EXwLMA3M+tNipTiOKoCS/
YcGbB+VFZB/n9OBTfZkQ6dQlPvDn4U77NrtapPZ7G6Zg7ArlDkl3vGpd3QZj
UAKdnX1G6CrNu+QhfavMkerXS0YmR7GjBhVbWp4gW+Z9ferXiI1g7PmPitNI
CTpSUMTcXfOv739/5wz8hB7nFMn57QvwoNK7nwwhTFeOqhP6JD4UPUMzQEtS
jVBz1jAjksO12Yu0DNdLpYfzmdWMyRwFvvhKkrsF04uijoZBsQy3zRz+aUXk
S+U4cRr9us/8g5o9/xux/VXwc5lkNxDfIKX0aIvYMN08TSNygAeRmn2b6Fnj
IAmErYzB4csjduedcsSG5BQcdeVHBeLcZ3wH4C+u7Jxv/Y4XJoGxrDPqYHt5
7BM0ADe+anTU9I5s09kD4RhpVRsU2991nqaRt37cPPXGbD3SNwLh4VZa8iOd
Xy3Ylp/a6THl1OQ3/1+oLWzPYmT+1diGHITqIBUGlA+5ajE65Tmpv60hhgOM
R9LpKxNzhf1IgWddtARxB7/kUZTaMX6JokkNfDZ7z5jq8bEypqeKYdbYi225
Fd/cfbCutN8B1ikShZFcyxI+vuq0VpRlOQDhYAmEP9ypmAIWVdDrZgaNQ4dp
WWtxevCXKRVW6Qxs2W2M3XFvpYuOURYoJRg10wg9kIwpEWE6YOfbYPyXuGFL
o/Va9pmhc09Em+FYkLaxT91o0E5DkTCnYXLLiSVWtqBL4QJ33NPtZJAMG7B9
x1EqTWQAfKtFSf3SazvBvA6i0JpUMF1mame0TKpBwgA4wV8we0Hiit6Z8j7Y
dIKja8EqcT7o+tu0e38cOE0Uhxjf39THfV5x4sHLxfcWlN6UupavjRVYGJEn
EJQk9xKi9pzTY10h4lY6ERSYXEFtAU4ipCzCoPEx7I+2KqOWPYEj/7BT5/Nq
Hftq7q5GfbX4NUauA4sZ0gJriPruiLhbTnydK0ctJ6vwHNAX/JliQ9QwmffV
h4U1W4yHDNI8+OKTx/o+YhDvBugKhaIa3djOJzoDy5aN4fkYva+IUAff19UC
wx6Ezr2LmGYn+RTk00o9VPWYgZ8WzcoGY7uV+pGNMNqGXsr748OSQAB0QGdp
lmsq54YSjqHWeb2uyxewenqU3laZz1ChsOoYAAKdex9H8NOVdQVRylFuF9sA
Pd7qRTSFPqG0UrWFqY92OP+V5unFMFRAk7qyowUwu7Ek3vly6PaIW3DzjhAu
hf05aMTPpUVA3z5NpA5s4m7/D8M1gmbVIpZbYQmGlovIs3jOY7b8Jl08A7aZ
FgvOykjnS4/5AB9AKmvQqzFs36SsjWP2470GV2OhNv6PWWK51dHJKvpN01VO
/voD6kWQBaaKsPvHvwKahA6ujCsgOPMtf4dDUrlYLWl6pFrCqjvPsgISAHIr
ThJ3FqZ8tzraumDvFnn7OMiXfEejoy3aVFQZoxlM9RTiiM6qAFuXJw1knlgQ
gBU40xXuqaREkfCD7Y+04mi+J/GbZcEe0YECBA3yhU74LF/ZsbrtP5C3JUdS
NgnOtCD0szQJ+i9G88d571XTz31fYQcpRwsRp48QmB93gZYjdzoePvQ13j9a
W1jeZzBAQuvoEjUgWoDR3WokQoEC64ub4rMH61ALMy+QW3VqBg/Je8+2Y1w5
7xowX8qSmOu8kkgkw8h+37C5Z28KdZQZGkshY0TJ2luZJ8yWayrr6MXsGqHg
HGjNC8xonFPK7uk0avRCle0YLJ8wXcqSukpLEtNBt11wnU4skhAXrT/hj1Me
Bb1j8o7ACZqyzb5POiT/qFRaDxxlvw9AY6Ctwi+7ArX+8El7uG/JU0k3hXDk
T9pIBcGIYx9WqgCL8OdfdKNQeMe18zbzDFlFZlj3Mfg9Ay6IDK6AobT8WS5y
XSYj4S53rToJ89tV9RHg0nPqErlOpk+i1NjjF25h+qQAvVNstBmbrhMAcgbH
pqpGAUT9GYWXXDA28HX6fM2D+ysPBdravKPfSmNiQdtD9rSzuTkjqWjD6aDN
MhipHBc+fjqFvxgNlYC1Kh8a9tE4buNC4f7rk5vnFdpuIt6pnx3C3apKjh0l
pmDEK+7K23AdnfQtvVy1D2+YTHzGlLkHG+n2MPnnWFPMR48QkU1eBuQNPmUW
OxIDvcspCHpYv37Z1YqC+duc2aQelwAry2RUXheTWikiIW8o+7RfTJ6uVaGl
ZLY3PJrpCMgQ+xB+3dm8ZrJZdtiIHtZ/ZfDDEPdCo5SZNySc1T82+3CAnAIq
OE1WcQl8cmf+AUVrezBMpCnv/vWH31Efd6d+TAG/bCHZU681QrZyav8Nn6Bc
VjCKO/RAHucb1NzH39TFvKbG+qWA/ZKJtc8YB+EGh9tcLJrsIeO6TzB1NC/P
EaZ3tQ0WqYWDflw3gFseiyEeEg4PlloFKA3Ji+ic5+hr6fGq6/ysldVlGd/R
BdOMqsJu574Ci9wekkk3F9DVok9BYZkXB06Y6PZS4WcBNgR4kZvbMDCnPEWf
kEB73PmM58flXOuld1qHAOJChY0sggn+epXt5RlkwguagIw893kh2VxbrTak
2p0o8iJZcFFAcIR+cwPzkDTlkH+Q6J7gsWNsz1PTxU2AHlGLNlFnYbMRwnZX
fgTbzjh8wNVMFgpR6iCOJwnZyAoetLJAdaIzO8F2NPuPmLW6TEebIOzGs+Jj
1UdhoBsizlMbweke+7cLzFeV48MRLxlW7CTMXwBUyhZ9pMMbjjtpsYvt1j1r
Jjki/gdSdQkFG51uDjhH8WlrEnLhPRGlESKG0SJQpGRfEZVddNIcS/vvAGf4
ewhZjHj+d+qbKxQgNT7Qd5mfLX3TTwAgTLc7CB4qB3afXkuOZhoT5UlGINVD
+M7zymwRGNu6a7zkdbFJqjqfCiTNDOweeeNMSXxEt4ufu8PS3x116giZvXIA
eyipumRkusc0h7F4eflQyw571tOPuVwnSuJJRSJTSJ12JwF1w7ufjGoYIo+D
v6+FkZ7ca21mudgMluK95IzKKWALbUM29Mol10QltM609bLhytimA6SdKwfd
ZtGvs9rvxhdAazk/X/NCkft2t+BlckGq9gy/bgnQBCxKTEmiE5fLSYWLpn5T
EEI1fwn7MbR/nd83fDre1KDnEWH5oHzHYtuHwTCT+SbO/kcMlWSKMXNK7p4l
c2TEx668fMvYuwlfdNA5XM8ycPSYmytyztQLFox9gGrji1X1QeyCGkSFBTAP
XRAA4PGIOyKDMAdu0MBSb+DFLDKcj7iBCfUZXLnhJXCfHjWAXWBO9vudI/ht
aXVodrVY1VcBdHrv/leUya8rLgz7WLZpWvowtB9A8Gzx5Oa++ijJU0yov6u0
QHOeptoWRyCq7tc6mVPcy//PBra6b+z94P4xoKVzZSbLmw7ALnTDI/837r7i
xed4cYlB83UW54cuchzyGhCjJ6elZ+26UZMXH7ShsS55VvSoZ125IOfO7pxn
t3XCqSPhjYSYmaBMKRxfwJDdskflVQIFIPS3sTYe6IPscACGkR5NGNPFRbHn
V6sMcUsQQRTjUMKw+qU0hsmEz/2CwlCecaMn2EshCYdM7RJKTgZZSmGy8ucb
S2dOAe8qoj66Luj7w8oM4qslH+ppHtp0IsAKsq/tkH9RumgziWQ4cV9HrfUo
6HYx6iOYD8UGyOy9B/6XlJxG8hCWw87EkCPV/pXldFAfNoHzjWuOwBVZqHFY
aZtCN9pPXCUc6SHYbXufUveWGKN3OjYww0BPXJQdesIZ1YAiPtysKnWl64XA
oPUyMsL+5j3sITZyIDnZFIJEi5/nlA+n44rFRZ9YvGnP6cuCt2YbS2OAWAJz
OaOoChtKcILwh0nozr19C90lFIA9VOm86UarsATE/0SDmhpJmAAd8kE7Ev5f
mKlcU8snTGGR4HKF/PTGbFJqg4QOpH5CE9TCFipkhibcHu9p2iUXqdJFzUwu
o6Fe/VqNwde07Ty0TkGlEnE8zxgW2phIjdctJEo6P675mp/oseGx/bF052rT
yfCquHXWkmND92TGNrPio7ye41Umf8Wue3JpI0fAhM8OEVAVUartUqOF6nqj
zoJJ5SGkAxWfRu8zNplKUxg69XNvPTG5ZhsOhxrQSQOXJAug6Gce6b4aFMd/
fyKBXrF/QPKZPyUPKjMLWKvbPxzzmtkQS/lcgQgkuqQJdKjogfgH4i7cChdE
SaSjvcjxmC5q7Ln7fI764xklxvKJimD1gEO5Hi2L7Luy0bDCbuJUlE/ls0+x
MLUk0XaWJ5GGQjAYHeUDAyyr/nx2e8YIflFcBOAuLL+AQdrLdx7N34CuPMn1
UCKoV4NuE0jEGGSHY0jA5qLdtG7JbMliPfthScLYSGlQAO4S3+3EY3UzvSTV
8SyEvf4PiYxWfHi2NWqnhZySP1Kx6TxkBNwESnHSXop7f0p8obaabrlt+Ue/
IvKL/0uwNFasnoazwLyoBfdNLOy7RMlE9X9ZUfCOHL5ptx2+qPnBbjlCiiAM
ojz3xQm8r72U+zfCL5gted/vCpIKCv+tVXAROjU67A5KIEiXbAQsZ6YuVack
tF3b4gEQQYsspu864QIn2l0OZ1LVKIaNTZ3nxmhvX/gxyQVr9IDNTK9n7bPz
SmpSP9OX026hGua3kcUohXxE8n+IP8d9mfe9AH16v+RKWx7WuDFxZHdRcUo1
h9pUloDU8sfuLyOTIhsblwSoTxI38/KXhNRJip32dr2rxWDW1Bp+RYvwOkHZ
g75ZfXgJbPODDYGEXp1UpTSoMbfwiQXRqkWBWJBGkovMg3k7lU1GRpUUHHZ3
o759xlF6kw+46o81QwyNMU6+kbqp1rs7EbCSu8X+VA1F03uK8yl9hr0jUwNK
lHgM3UUIVONmW2626Hh8hJf1R6sXF23GGSi0fF4YdkghKDQPYaAZLsE2CQoD
aJ518FNgqOHyWvng2TutUYdCPgGA64UdUWF0QHn5VmiIZs5ufGpYhAIL44XY
ZzuO8odNFjC7Y4hbDJtN8d0N0fVOHUR7PVUpvjtkdh+usxO4Y8jLyNavpm6a
oSh0DiZO5rye8cm7WDR3fuHyawAHDUvDd4qBFD0wDQ4YMLqL2WSC+6ea0TxB
CirJXdzPgUu8ndlCVMVYzOjTk3DOVDhHNkLB6kccE19oJa4R3Sz2ahYm4BfN
JWUCtxU2xOxnpLBj8a0DU59vQqRK4lR2vhCpOtl6uTXXS8Yg2kWDQgGZYEvA
0iBz+Z8EcEXp9BlBN5qWxUcIIQrBEMSGusyO/9faXkFGJYz3M/n1XLCAA3dr
iZ3rdMkOeFsVr+0xPP2hIeSGqG6nfzBIn8Lo0ac/B+7N28hKKMzpfXCz4617
VPwlhHSfnoUrNb4sCF4l1K3vLP05fGJ0Vr0omnxYvmRgKy1sQICEG1n/fxO8
mcWMrdTKWkr9st6FShoewuJpOkWMDHk8gCavyLaQDZICIvsDh/h1edpG9UYw
5AuQiaqbEfkqjoZ8Y1oNgZ5zW8TEOT/9P85ojd9RkRR8fjmIUXUZXXyZlulw
w+q83bu+vC9rVb7HZGlBQs1Pwuvva+/LpDNuWleKCVmixsNzvk2Y/qm5q++c
BYbzTCtdscTllwEcDcW2AmUVm90yAHIDMV/3fwbaaK9P8RPtbp4HN/5JWuI3
Byusee4ayc9gg80ZvTwZEN5lSuri5O9emGURMIhJ7HPblgvhHHg7dv9bGnOW
H2/1dQJs0WTu6i+GFbPWqXibg6VHrXWzZGvvWViczz1YqpMNXSYP3ejkxUkB
xZ1+TIUpSIPXDE+ug58OvOj5ONg6YVyhaOLfkksJa8XzrYNFBuAt1CTCyQQM
7fTVgB+BOMAXZ+LV40jve0KB+GzaBmc56OvjOmboBsMqKVmP7tgTcqjFMORZ
N5WzQA/a4eTMZBmJN9eFOJMTg2b3CDtWcKRTMy0VEjjcZ7fpPOeR2EJ+FRVX
GiM20NibpVReCjicvppmJgR0Be9jVm/FZ+z3gNzHyo/5Vg9oUXPtrwxv7/XC
T6juU4VhOj6CmflA7nOzdKKAstmHPTngeqG9cV1o7hQ4jSA7u38WYLC96y35
rAifNWeahlTgPdwmVArmgnAxgLA0nMg1LKapHp26y1jE76AXg+sM95EFjAXB
f0Ti3e6LW20A3vRGjskYVRnM5w20v40G8GLV0R8HNk+TiqaVnlDwK7BkHIJ9
TmhWCyraJg7ln4P3qY2Vgdf/S8usAJ6MPKrmGLfkG44PKMXa64SaK1veSzOT
HNbE5BIR2VR1KUZmyatxlFu+2TS/Y9yGrbMDTxUexG7Xi4b0BaOVD1Rw6rTT
851gBp9U2fwmQYKW1GdEdX6sBo/22e72MqJKpQly3SlGjhh7Y+/dqJKxsw/N
8zhwCIBy4xYql9xsSRjFnru/dwElHtA+Dq8OYNFa2eefo6JuWmD1qbL1GUt5
8pYgW9PrA+xU31NYeMi/qYLO3wGBDm2gESp5+iHAi4V6qi69Vwmk6quWVK1Q
l6sHr019SP5E4M8HbEKFvsv0cxi/cZucmMZwYpEYTwqmpfy6p8toSGy6UETU
PuskJAMz5gmmo8iwjAyzXQHmzJl0788jCyvanp94BrMaFZScBH37Avb0Oi+x
awa8hdbDTwaLOsL+xvqvVmco3zRAm3lYv+jWzpwObNl8LRqD4ohkCujBz5Qw
Kh8QTTA7qVvF0VGIO4JY1t/3XoVrg7fH8+WZHQfCPkNTe69GJmtSRRpnRAh8
C2JiXrdHG/x4bvlG0qiGSz746oecHS5kKL9Wniv6iMOpm6HoZRWa46ro09Vq
8YZhSmWza6YKcmutuq62MpKLfyUOAsj0LvSNsumr5YorSCEy1l3XD7ZGCJ6W
EAygRHCGOdfkbfiTwXJTxg/KMdSewFJAaGoA7Hlq94sLAHn9p1AxyGFTJWyF
PojUqea3o78ZkBCVf+XD7j+ggSFJPhwJ39RuIc/ChGHouQpYAyqDe0Y5LKX6
mL/dr5EyDR807XF6YMY9HA/OfVPPEfnJ71betPVqJy7FgFnUDmxMHE3nhGEe
Ok1W9d0j1t90C3XtkfGbooNAsjZCTRvLSPN5aFDDeyXkkCCkkmavuBr38klg
qrYsXf6mPYiQ+ptLuhPTmb2RSXBXVQuZ6i0cgHZiXQQmtmdZv2vt/Nl2EFih
g+09ZPGeswDjylMuQ/4oasfrei5WzMBJfgYbKifPSMfu7SAxR8hjJybvgNLM
OQPDSnE7wNb8mEzBkqzX5MqSKi5X8nPz7SfK0TK/tIoJaTgpJ2LOMXKId1V1
rY4tRximNPV6hzOM24lupJNQn8I+3LsiVR++eOqlrWENwg3DkgmBeNQrLCLl
3+np27MrNpK7sr97MUYSqhQMpR7XMnnBjf8c8ZTjHMYwPhiFTjZb+Rlm2MZp
9+akDL+RWM6WtewNheh6LajzYsO0Yq1I5UFfHbDhvc/3FZklfq++gJSyoY8r
gLXlfR1RcpizpR+lxaBxPwEWx7rEUnLEM5qCK6f7M63EgBAiIDTeKC4sK2wU
0NT4QhBqcTQA1RQsjQbJXa6srkTF3qEyFzIYkX8EWBpUauIMs+NUuA5AZ4Gg
vRfryGZp0nQnKh9ykrsUOmAbMrISyqbEm+Ytkms4WnuGlys/i7WsL/Xk5kGH
5VkKGUZRFI9n3ZJtH2RbhJmtN9jyGNl8HtY+8mt5+zHBYmxi0Yytu/4x8ISM
EGX6S/r85mVqvan7yGeGCIZtM4iEmN25T6DVABmY85RgFPvBqt5ccABEm9In
3TBxlzAe7v5viMKs+Ch/gXeqS78dT0AWunqX2H8tOttujznS901zV/Hblo0G
R0ZqflszDqTX3oMSEOV64oo8Ms+V1G2roLWI15wtj58AhDmlf8KNrydQTQPf
K7gSYspHtPCbcCP9NNDlxAFKrubFVZkHsUXyTHS+Cx2bUX4RV9rRSm5O7Ffq
9ep7Ypzg5bjuvEBDcwX/lrK2Cu4KksCSfMuv5ipOKMl82Rn84aWQVdLMr+Vi
lmYEmSu7aQ7D///qamG9fW/CAbMT4ub99LRzKCpDq2oXb6cgdc6P0hYeZCZJ
HtNvYLjyxwZmfIfnYFEVYQAkiUK6A/fvKaNdNLMiUpyDozUjaTjiXnAIiWv5
KHMUVE5W2r6mHs1XsmESrxBiQ1EAKLYQk4oHDXFBHNohnlXKkFZAHjE8qK4y
ltBO3SDVgmb7x6j4rtgPeGHnBC6S1JrAFhG26zcw9k04v9KWcrqNpXDFyrFl
qmQzB6uV8Rycsmy0HmaGJVEy6Wp2yxD6Yh9vZEVDooJBA5A2tb9oCv34+pUL
F7l/rYXXkJiiqItWwaxMw16Ml/CsXxrSFS0Avym6+qzIyUzmM0YRz32Zd1YB
QhvcjurLmBZnMUhbt0oTa1gmnKgmCkgEe2w/ZGvWmon84KXQiuDUXYg3RNjk
wgtgdEG1qkG5p3QN59bDqLCsAxSJjWQTnDBfE/xBoA9j0jMzJTcT8SliPjh0
avGGbKLiVj6UP9UmJIZg41JTdQ0Jz5G22m4gDAdSzoNrGMsLoAX4mJbd5SkR
MPoAnHBYmJq6K/bznv/s3Nf3cjJG+9fmdmvELIgU4ZkF6orZ3fMRAGWJlU14
5Yrp4inYYfCocJ6hIF6+cXt/WHgpqPB1+gv7i9Zl6id7+kFW8PuIO/v06wIY
wPXZI27SSDYj95zvZwC2zCmrU9WD2MkjhVWTrnOx8h/uvfVwpk8O/VeGE6ab
EG3vIl+6ervQgNnFH7jPTk7WG0HylZVcFP397tVQUbhZoQ1xGE/Wn33nFb8I
CT763eWexXmPJFT5YJTIe+zcRD1sanclQ0NNyRd9qj8eTB9zFd6MSRdHr6fM
BBTqf0R6Rs0ejf5Mu3MxbIHdp7Xc19Pe5mCu4nuclTSqszIzc6RxY1ahJsA2
qJDlIzGCZQTwZovK6gUp+QWtcqq8VW7mAp+Mfk2kqQM54DfJyHM6NQ/cInFz
RppFV2dgPxn6jbc2Dh+E5OBdK6cSwDV5jmAvlm32Tk5TV69E1/S6JJN27d4D
zJriSecm2a236ql0mFXc12lfnxTfPQhsPzyN3OZHdrwhKdvDIsrEPfEdIBt4
SWttBgNCOwVZEBTLGh/9C5xZm2RN+EWZyXR5evODnI/wF4kfwGHoefG/7uMs
Uf63FXvxzyRFsOZ2Zluz5cDAdIG4RlyubQ4VMJK9WDKDNwUWOrmWV/fDJmHg
lZ8rl15tEEkuGbet5z2q6e2iXG2DREjoFKxpBGUEJTrqNkwMocxJXisj1TAi
g7wckhrgVN8J9HnMgN6qlm+OO+axAY3mhsp5Pb6xKnONhiauLyE1HkEE7Lf+
uYKMIIpOwrc41/4tmzK1mxd5iu4+7w2AIXYuUTMvWM3qE6j9bk1WXAjp2AcN
lXCt59LZbhnblplkpbNVo5SCgWWP4v/UvgEyt5jtjpCV3MctUw0C2HCPPQdj
XFl3HvNoS/sl5BgYkLtWeKwmNNM0FvSySI0qOOsFN81FNZAptdSunMZbtB5d
n+h18BCh9UG/o6vC8x/NRjfIRfSHUXpicmxyXXgCD4oPBW6OQrzDcRkV2th0
/JlvVJ8jSdv8rdNpKdxlqxe9q2zNe0fldDLJJVYkBxLqMBJfB3JHwz3QaJjB
JTQXl1nefMQNiz0syM/P5ARIQ4sLpGVCdfNbSuQAF4+bsb7M1tESlDj6Sdwg
9EKXSYF1gd4WHln2ubNC2pIcMIpAfHNDltBJKNReA+pWFiuxMrMoqQ9lcKNU
+9GlGxSiFbA03uoBDUKcIXu0z3tpuQsGrRA+befJq+tFMOcCaYxpM9oyPKq5
NBD/Zb/EGsAjN200rZ6RH9uWUjcUHGe9g2iP+KzemJroa0TEQD2flGlVGU7I
Jp2Zh7AZxXjD7IZs/cAGTwdCYwwkjgS84dbPZ6KpmItP/JQUlgtfJ7JyFlxF
ZY2ULSLvt7QA3GOFE9CzImNiXny/Udjf8/eNiyE5xRyvj8/kdbytAnF3umQe
FNaYopp1EhTVF9EwsIC4WTW7RmsL5k2A4wY6dV2c0e2jRvypOeJrM5cF6ivP
0s+Qrz8M/XJTE0aDQOCdv1sC97WMx8uZKIqNNzakjJ6whprcJPHED7Cqh6Lo
EPt1+u9KBLrLY4f8f1/SXjJvalHjEQVm005PKvLcanvlPYQpsaZK+7MLuXjK
QgevOV5kLuYkLvVyrSbsNr16ilaYXbF8oBf8Rz/uts2j4Udo0xb0KlbujeYq
nrkVLhrzfE6ldYSg8D34ygV5FyAIGuI2zZd57OdIsLD4VsWJFw9EHsFBCxwe
+P+i0/EFI8VUiJ1AZdEehG72Cw6RBUW3LfQS/gcFkyO51P0ia6PuSJgf76R/
ZKtmtCS6II93qBPI1Pm84AHwhkUIrZ+3RVtG2ADr+0v67+GiwVho7HCm2v6+
wHuXbkj4UvFXQ4zTe2a51xFrNt7ussG5tuc8bkKZwVFA3yVkEV1++sBk2yp7
LMTdtB6BFM1rDspm7/sf1WO2rV720fozl72nk3D8Ob/CSqU0SS76GgskarR+
qzHtFL7S4YWJeczHTbd4+r+rNvkr3IcAN+8m8y9Ig3h7bMdzmf3MlzGHvNKb
QKmz8do3Qu04NnD7lsOtQ5SpgBzAA+BZgxaHDtrW5yebSQWprTfcv0c+poGs
MOVbpRaOI10Bi3NN2ZN0+2zMuzWklzcotD6HUK4QAhcV/k0dpMoAeIyq5DP6
5xbTwDlNrBGfbjeq31eVRMszpR4OmCYTXb2BMFWvcSLWfZe1vu88VKcQDFDg
xZISocoPJ1+Y8MJ8sZSbLindhzj42amnMO6tkeMfznlCXTklPgc8gUXHOVlO
G/Es+fhtE+LPzG7fPSZ9EGbTrroNONaRXckkytmJJu+9vKC9dyBDe4B3r991
Ax0VKf5495ML/KLvg23WXu0Xjvrz166pToti3Z5jo4IQWP57TVU4FRLaFFVn
8MNADODIzOOlkpXE4QRPpo636SJs+ZOAeduvn6ZyCdrsCDX6NKp+IXMpN5hp
yqd1OGOJNFx08ghpm7H+jXE5WO3AFYEUMkPcLmdv14F/yIW39Fe9YZnk0ena
sPqumOX0Q6u+A6Sstbg7Frd8S4Z57BXFw6phHPvRcJn6SUjwQzKwKUtm/WxK
QZ1EKl/+84exalr1kPwK40W9IpwSrFuBKslMcfpukGXLBzZo4W+vc+yqh4Pt
MYfYko0ar2A4t+hwb7INpyxv90EFApPJKzxOISY8G6siqa31lAOT1E/Ag9vR
Yy4MFHIJ3nA6P0sq1nZpJCYSqyrP29RC+eiOIxU60mOQTknm+uWnyeyxuojN
A3evnPsYddBvgGid6lQW4F+riGG+J6fxBrNeynb6r39HZfhAT2sHnZZ8kpea
0UJjpOqbBvGsj00x5XysYAL3ilUn9w7o3FQJoAhXp954cHJZsd/EkWhLvwFo
OV9luGuxfGgYSLm8j2wZRZJuAlNs7jcluZ92lRMlziJA3vJnGojXe3kgUkT5
GSUlpPPmflEi1l9nbXerFymyE7YAGDot0RySa+pVYcmy1z1bocCsDj662nxZ
Koq85SJp1u8ZShLHRKYeuIzu3DncOZGmCRSXJK2Vsh90h9uwauIT341G7voD
cKm9Py/WjaXZLrRXJrILyVsCU317UtTO3mATQgVU/TSEf9Vu25+2QFYaPbyT
BXusCK2Db8gm4TIQ0vo6R/Ti/RcbaWbRvVsgV/Jnb/NdgXt9JLUxq6PwX8W+
gGqPtWf7eZtbTmGjz4BtStmxfwCaEu5Wiaeukhvv9R7MH0YH7eISH/hHWigh
STTa7xE+x0W5GnEcMyn3gIqUEhuozK+Y9RD57PGWax2gsvKQquf6UmE2YPTV
Z4IRemb92XO0Q/1geunPfW2tiO8m1bwSjodtPv3pR8CSui7CqodcPtG/7Ali
Ph6it3eZYjJDtN5chYkQNuz3A7SR5TMti0iA3E3tA+uSpT94hBuw1hTyau/G
iSvXd/WAg5kEZ1jki6gqKMYPM456vUr+0jnXDiZ2iVvzt+COzoeEtLEoiKlY
YDRWs2lD3u1MOB2SN3a8za6eMVZU4TFaoB+AaaZU/R/v5HZyUnZN9mCTn8WZ
8pZOrOuPRSWuGCJdax7PhudFU2Qt32JRi7BXq2pKfNzC0//q8PKwxioymcO4
N1Mn7jmmzKMleN+fO2RsU0trSAEN6QZrP0Mp0jABQmC6ctkcDsxeBlLjTvX3
liCT7dP2oRpWedqGJmJ2E8VF//BX/olaR1Rropjcf7RaGacwAimxJsd5RZJa
UuYD2IxTSI96pc9efrHthQabcNB2/y4dXL/BrAxbNGsj3RmvJE18D+IUc8+W
4p8CznZ1HQP+kbbLAbvyY5Splc5dbOec+hv0fcDzEbKN/x+eOdCFdDLxFFEu
c6wJNVCYCHSd4eRgGOPr19XAVx4U8rhWXfRqgLpTLR8/Ipd55+Yq4jqPLrdY
ayvadwg+viKcqDR7hRIiMX0SxIvK/8TJnv9jtHU7y6lY2KC2lL5N/EEtI3V/
Gm2TDsNS/+OI8A/Ed7ygFSa7k36Tqnbf+K32M1e4Hqqk9fiacJ2S6AI6VsW7
ObPm/YzT4pW52Uk3DDtRLKbBp0/GzwxRdz0fLndJD1cw5cHPJks45Ejyj+F2
zHf8/mKWaw7yQS5r/zDlQAm1xrJF9NxMPr7AJrcpXdyMDpWyb5lY4n6WlAtU
NBYapvhssZIBLi6lGvkDQmO6qC8sSjSWfh/3jVBwu+Dp/P60VnSry85khwFV
jSWw5y25ETJwHe6gF3KTwbUGk8ejvYtHw5b6d8KtZziS5yBYlG/v4xbACsW7
H7VEqMYRXAj+PpNE80Lx1hRTHRFCdyYr6I1ONRPqN9p8FFlHdkGl3zRY6U3f
EKMFNHTZ7Q4QGN00xSlOdewkfW8qbcqG2LSVNaoGVkIzY9zW3zIi2+Cbj435
Q133UK8tnMH9w8HwLcQdhzad4eT/KbyIQ2tgK+s984j015NU8p1Wu9LTEeZ+
C+PbGu4Jun/YC7XxrYKBFODL8Kf9yhY70nerDtAAJ9to76GPq+GMKLVh7Rkl
+UjrgnoJyPniYDYYsBsw22UsmM+dVSiMl1/4jPzuUGvhiMrJKVx/jxf1OZr+
/YoMPRnnZvP3tg8hEvVtsM5ycDUF/7AmgHKCUXweYoiZvR1FAWXeEmdfpoPT
5JA/6t98xl/kP2F+qZQaiwAD/4C7gSr2/LYQbS9E06DHokYLnBglNcGiQlGB
ffUi08e4xtCOFSo8GbD0zoNwYt/KDwjpma590QaIQUiBI6hzf0fR24pw5e9B
Mm+sDleeW0lap/FxQ6nr+fGbow58Dv34ilWgWNvSU3FRMOXMX8Oy5ydibkuP
LkmjE7aIgjo+3f17QxxcJIYCOAc01BXF9FCMRZpHKkghvhBMlnDDJLGQilWv
c7vukmJm6VMozDVMb8w1u/CrCCgMVYjjs8kYMsygoVeqI7gSsA6tdSfflJaW
RYz902fCtMYGyjzELIg3n82kZbrN4BmW1uWBejAqfhKATcfZqeXc0TMuwvS+
1vCm9PGl1lanL8L7Rxw1LsLavKn1tKAgInCuQ2X0s92JrtgxN59S9Z1M816M
DTX3jkPzOQ51F0f3MkTPNwqb62tqM+FJcjtedQKSXDTXHbWx3aNpjDC3GsVE
AXy42fkLRS3tyzIy8E6qe44O888EcR/D85bbNXsP6s4N6u8JauVXL4TNgfX+
WpnZa+Q4Oehj8uz3Dya3FPRYFddsPG2Kk9HjPMU5dbIv4jx+UZeB04dC/OKR
8Lyoqaz0/0BPhmnMuXT78bBVLqBJ0aZjIN26d+jKl24/gaHSdm8emdl2aeiR
g4T34n/NXTYz6YKaMo0thTbEmsZew9EUO+NxCRgeuzmoR1RmxxoCCHp3DoJI
nOjGGBDc211dWXuDEykPnUJ+CU0EtwxxiJXsf2GWE4o2Y//Hev7hP4PxSAbp
XJVFsd84+wgpiUBtdGmDfdUOFjNGJMVvU/IChH0pA0ldqmWpxflpIE8XmRR5
QPWxBWXUJmYzmEnj3FW1ijjYzhNOkFvoDy4TBG3+P06/NDHChlqE1rN/2miq
HCIRwXO4EbxcCcfsdE9BKiYuppy5C6wd8Nu5kiEKpr8aAFYw3yHuRckBT/V+
VgP0+Bnb83hagV8YcWsot9s1RHTEAP194G/YRljtTieHrJRrqoDOo2O63/r4
aF6m+DdHO+yMu0XAby6iBiBEfrIyj2Z4EpKtWpe22TMg+SWkC6+bU7gFjk2X
2nXKx8wnOEK7Ets9Hzvzawen/3b7ah+d6QWN5vWrWzT4jSZpWAz7JElx1n1Q
hAPfZ31I7aZqlQu93Sq2uGeDXNZez/n/NSuKnjzWWAgOLsmtk3DV5K4MoKhl
EcvWgEsnV0vvCpcmtj/pUxJIPg/Lj5DnIzvIUW/oOVuXQnmi9FjeDNczrP9R
+XkUAUNlnRtEAZcTy8+71PSpH4sVyV0CV56HAIz+JIXy89jDH3q5axlIAiWe
ay3U5dSYssEl8Op606vGlrBPlHowCuGb3wAUlsoCDNY4LePYbnPDUsmfHz3u
A45FLCL9a9Jtfu2auaNhHkSnJjIs6KO+j9KJ1LpOdPjSyY/Ax9dV1HfrfwGX
DYJzjzoECq9XMfkLKIDVwt/+bME6baMXBBFY32mbQ56GWDnweSEy308IIOtb
mYDkuN2cAGTDFtahf6wZNQS3RrwvU0CevBFXu9MDEcaTCuOOTJ1J3nbJfkwU
bR4BtcfiANNadXPb4bvX+GrY+9P7wcempKlg2xv6pwpWPH/uHIskpkhqxQhj
OXLrWLr0maeBdtWzupslKOtYm+NFKlbOdrqZQsk1zVgxjiuUYxckkQ3opg4w
KJywZDqkMK81KSqIVn33lP1mznpUr/m2otFPj3X3qdAeeiofusKrEkDY7M70
7BNhxpKVc9hJDKGt0/+qexFhJrjUrMCurVc+i7fmIdJj2cwOUhUyruBtUahB
75qR3cTfJi1N0M467gyy0Ba7VGCFqhwD3vmZZVhFLwEzd3h07deapqpYRqMC
qQPGSLdMqIT7ZyV2M1P0SUnr200kDHZHr8S7y/XeuvxovGgTfY2wfJC6iRx/
UAuQxYM/JmtXpXrPbc4qj5LsxomOsbg6S9/B/08MIOA53ra1GVGV/xMus8Gu
f6vQ5ukwX8oce/kZfnTgf0ZoLny4PGvhKjAN/P8G2Uw6fPGCHGj4kswogoSS
E+vD37fKBzgo76DrqPl2xLY6wTNqE+6u8cggsk9lDNAd9+W04u2NVzmoVERT
Biwjhg9oVCYlpizdx0BwDRwbn55LAqOB8wYbIvZF4AFzkwdF7eqDP42P2YI0
nPupqeYqw94b2LXeh9rq0F3Q9RAyVztKHnF0x7nzxnLENEnzakor+FwXG3d/
aqMq4e3hKq093NqRyO/Kxd+59Ct89ViDJuCvl5xLF+aD0zDpGJdkcklPHGBA
I6V4SOvzOKfIQa+rRmQ5VEFKYmGIfYSie6vRw/p5maR/H+R0xauGgLbNyy4X
pQ2x0Koz4KPZeoW8ErhFJwlEWmAu9BQr/+D/WRZl+0QU4bxL0JCSxsRCrhLH
8lNXkpE7X5a6vq9xD2xfHMdUEisy8ojPkZGlxHjR1rBxLVDP3n/ZxeM8SrfJ
VfrlHbsP+1owy/bbA+uTcF2NHgf5+5gghx+G2wNbCQZWuEe3YS6AqbW/VI1e
xAOHp10T0JDohxXd8ZNvtb1CTNyZ/WTs4Je/PSUqyw294tsSNSAn23YVfxzd
d3Sbl1sEpfCQrz54aeI9OFbgo3HqkESgPi6HG8MtURiLbtbfuMfKghu6cH3g
4BgL/Kfik1d8QFMNTpw2ejWPw7zV8mkVpfidg4z0f3IK5W7e6rLrPoJaxvAS
CPvt+x1he8QjdKQKx9UCUwprhDKkGSBKf56/kasg7CGz6NjMcX9eB3O3j7nX
iX1tr4URE/F0YLVyzW3MQDFq0WBcJiVoqnTuTPVsJSKzwg48fZ8Ai6jyBLAu
fWAGjPwp3OXgCtn6poh0MIMcIPYXpFZYP8Npp+ILqCbvWPPjMbzMGutRxman
sT7drQupNghHwtLFuWVQeV2j/0k0YBzu06p7YHFIDCu8u8JciXuCcx935sJk
B0eePpNofIXPMfYPHnEKfJKCVp6i5NTnkU73SGUvSZHYd8f+2kezJUXP8MT3
3rl43fsIlrS1QQzGzaLl5/hXyhOxkbuMhElqpUSBzV/JYr0LixkQONUMY5I7
DChHt33evA+N1Xxz30A7Wj1eazW1b6N43kVh5vMqyWF7HxMuA11DZeLfw2j4
85lauhZlnKVU4HtXhi2bK2KSTQ29FRDt98CQQK4Q8MbeACf5/r8sf0OJxXLC
vWoos2ZAIdSKqP03ULaOUpa1WmqVhKdc+frVpscgA+3L3mCyWA48AcCrZLzD
ELX0Py2hq7J49G9MTOmqXtAbBCorrK1V44iScO4UvVIhAo2Qrw08KjtCiJNj
lTJT7NpvgAJ43BlT6VFwy10pzVFTlGbCtfnBKeGFfJVwvzmGfmIAFoD2Ym70
qKK98m8fvfGaOMuEK1nm4ITVpjt2bdJIJFvU9Qu0H4h+g4bUfB6dh/axq5ey
jYJwLdZF3otCaH2tf0hmqVoHvwWCCEYNnWOXVjkyDCZqQdln92nNrLhJB8G+
E3BhJ7rSNAQm+NlXESTvCXJHwjvGGNxTPQlLXwdL17igmBcOjaiYBArkeVie
VHBTUJAScGrsP2ND2bNS6sePPprrxTGHSehN7mH8yLhK/Y5nsGC95xSKP5+z
pzQsJnK+07LfQEX3g0ISyM491FjqFR0mRQHvnUptteLsVq0kWq1D9MuEUd9y
/n/3zNX2uZ1fesvjWLHBKy94ypry8C1kqFJWjwjdRWOQPpPAZN5vLkSpg93G
Vt5/KNK95nW8bE3Fr1JFjNszg8bQ6LfaOdH1Eaxn4fvFTwmep7rnjopHqE+l
Yn+9pDo611Dd7qWSoZEg5atD7lFodUOt0QulK91IasYUVKEmt9u3b3RYqMh3
giDZWrzJ5UE/3xlgkK4+8pVEzz9O0czUp2bM1u3UTurNRwUPDEXlR7bB2nC4
G5PWEM2qAbYY8YLE1g6Kj762svCvPhKONb7McgQsorapMaUqq+ULZ77FS+GZ
uczzRIfvvSj6/kUZn8vyZeGevvrAxj/REpWujFt7Cz2AUczjx14lZTP6f0HP
qBGdrQdMMwh899IyvdiAj9orp9UU9pI7eW19L5CXDZ3sbGPbXRTrC6SFKOzW
Ol6+6jeaIFGaCgwlF/LIkgqxE3E3LrBj04o970deXdhi93agjMV5q000g9et
meFJvCpu7T7jThEd9ky8Ll1fOkFqwORdppK4Ssj/oJa32TTUUtxT1zFGrpXS
WI+zva8FJe6lKXs3Gae4+fecZeb/aubGcN7Bc6vUyNUCecWIBZ9HfFZwC8PG
DFLEh38zKvAfBXHSzpXlN6iyusPe7oJw0PKr5df52hGKiDN7IrNPLrfrrDyv
eVlrhhb+NF5qPfdeoYeG6xgSSOv8ktRzcdHJflSILx51OqQd+qIiA8tZ66ju
0qjjB2ymtqm31fk17y19RPnFAp4BD1Ukbgs2b03h/y75hDaO7HLSCUbB4yqL
dD00VQBNShOYq+22FPEjXLevnkPvD0XvYumw7pOHH6D3UPFvuSbiRPxBy0bu
+BUFPRPL9C8rPJpxV93PWUPOyU3QQqUG5uWO1kOlFsFrzBARtKRp8Brcg83q
kz6Q9YWnjun3Bv+GMfbDHx1tGKUIGUz7lvV2dQLEscYkAZTVNKVQGXvTeGd9
zNA4v/RmOpbaCDuswZeSXtKHjHQ+FQ3PJU3C88aOw8USnMu4JUnUX8uFV83u
gzlRRcu4DQO5x5VTTlwMKwsTt2xd9bixWA1DuIM/VNuIP5fQ3g+ttdrDgZis
U2cqlvGaC6eTAJrSs87yQt58+a2RCZ+EtG+TGC3PMcd7jnIOKnKSAmQ5mRtc
d3FAKGXbisHVlpm5g9GFTned2cILA3O9W2YfY1O2zUC9WfImAo5aaU769R/X
IHhlfKdqt1H+Uo/F8331BWMMdqZMjWdcfdGZbL+kd6q4jPxhAtbXvEnz3So6
Dijcuq/GUOVCF7/po8htiRoL9xFAA2q9aNxQESTfuraYccrxPW37AkRsLfg3
iAvF8a1K7QZmqImgPezfEVWKXvf95MfT/IXjVc81z88rA6pSeLFIyMuqPww7
Ff6/Leri3EfVxWbTIPcf+xVBmtWzLKN656SDkZ9wsNY4Ma9l5hOiHY9NOube
7e3PXACctbUN/C7uGwswpOnNSgDWPEC1ZPpKTrn5Sft79YizWZTQQdXbceIG
QzDEEuVeSs5YXeu5jecSVuwntQ/LQnODkoJJlVIALe3XDslH22e1l1zY/grx
2ygo1EKfW2vUvPxZ7coduzrr6lLfYQa3xgbzU9ylM+S9CNoNYX1yjx2eHeCn
MhSt4AxbFShRCWF0tiZbNo5cpDnf4reY3akHJyMy0I+sEFWjlqLVxDPittal
eFQfjhhekxYe31L5gcp7rQuSkHZe9lpRK/fOng4xKT2tc9/SWX8D76Vlc9un
31dGkjsm3b7HkSm8wicD9K1sM8MUOf6lSXRTQ+s9kJvqWOUBOon3vlRamQsS
n+SfER2KBGfU4zWqXxJgBnQEQVn1rP675hTrv+PeVJr0X4JCVvGNqnBwx9BJ
yitcrhJEwvz/Aom6xvRfJZZX3IWMgshwnLSkSpjoFJ8H1/KldV6uiDAZ3G3m
mw1DYz35cnpsEHNvStGdMMM3lZgo2WmiT/pMuPFP2Za7QNFdfPzsoK5dvIl1
GuHu220DYVhplCFkD3SRRxKg89IWFgxcA1QlBeKTN8AGSl4XNZDFSm3pLP98
zLKM6MsHbz6fk7S2iiOLWnDJhY84QfPeclZOw1LSjAwvcrp2ZWLRcGLprh2c
1nc1R8IgAMvJ/LaD+TwMFDcYeZJ2s1ZLHM1IrKuspDcsXlqjNnfE/VuutjbX
S5ftYJj1LRwHDoJ3RFLzjsG4e6Xmmwzv7AzOCQWvldrKJjWjDVVymOZhoghR
3JoYpq7SY9QiTERHSgjXsEgiHVA5lMohiUJ1jzWIGiGWj80al+Ig3G3+b+49
MBmvM2wg5zFNwDW7BwT8tU+7lrCtXvd1M2gt5nn/HoAQnWhJnnQrL7qAeHU9
fpOo997oRLFWrC8L5QioSFveErz4Qfae2eN5/A1aHOvpuv1jSgQbWMHFd7aj
wJRO8FfSrWxzIOvV6uRPRvxPiUSlvQOOY6s13+ru8tCfvBGUcpvkXe/GmwOn
tazMRC/1JdFz+FRq6irVDkILOnvCyOiauUzz+VP7mxw2rjRaZ8JN2OwE4S6I
eJIr5mi1x4/92tJ/6GGDCQ0pWHxNfk4j+rftXaYHUm5LtgkF3FirFpqyEnAD
n5nNPCSndvH+iL0e4i+6wnS4AQ5G1KDrJ/9m8bHdPiYqvemMAiUzSmDB3Pxw
h8VkJhiKq/cybkiiHI8If50pse4axHYzs3+m+IEU/pvyrUINpTYhtFO9CVHK
J29rcdDoes0BU9IrqwvEB0NJjHkhv9IXwwVkgMUNeW3E1rI1gJu7QOdQAtiN
5yu/H8MHAykxdG8Z24qRna9GB2oc/Ek6biyGTmO+12WkYDFTXrvHpf6y1jiZ
fMG1szu0v9S/pyt4zbXKl0/fOptCQFo+Fr4oaYnLjaVdNotZ3kRY229B9vFw
yVtliASv5r8NmcCAe2NoFbjDo0t47I3Ci3m7pisudz1G7epwlniYGCZtVo4A
78w5of1b5SrIbTzBR8yZAs9DqwSQHVzhf2ZbE9OCkQZTCuCZzeASE65WhYJo
GOyVo20PsUvGxmRGEMG6FiCWS4yiBtXEiuud9Id4Mv4vX+InRkGBf6nWBqrM
RYJfrSIpqQPT/j7Q910rpGgv3VWornb+/wL+PtWIuaJXhGBX8MtZS4q8WBgx
zqUjClvKoPU+bUmcrozuDWzRnpKIVwh39SY7jw9yQue/v2uLdgQpEeB4oFLM
7Ws+PlhgQsPMn/bkH1xcN8PT9ZrIGpG7CKbDLAJZUdCuUdXQ7p2nFLOEmnfk
szFj3lDLqbFhVkU2XCMrI0/N7X6N9kxIQ1At4GekwhbTDm0VO6Pa7K0bC/hJ
IDD0vc/zOXzG2IaKdpeykkPa2K1tKAl7/4T4/mZq/9BHwyxXRZ2VClFhAiyV
puM2nN91zs+ld7TwnGKvCc33zoA6Ah98yj+DXSIPe6yHUqCZVidG11PoIoIv
aKeBoaKM1nBUkIF3Kk5zlmPxKAjUL2nEvHQoI9CcOi/wohNgt0BSRdOXijpr
cKVIXfsjYFeFxqcyq+VjLVScpwTjMzYyQxbuZ42GtnuIlx5mjtqDcsCWmLaX
Zb4cclwMnqGQOyeHQBpHQ9q3yNpodEjsvEDBZI9g9GyzhXPll3QdRWGzMWee
3gtUH7AEjwPAR63W2u1lHOZbF7kYcvWCfN3qC86cK2Z0YAHEtlsAu/7aJreg
di1pdo0yQDP0Sh0s3M2byE574ndFVlOvtyIXkemFhMM+gET9ZK9W/2wNUyKk
zTMIJdCPVczCl9NR8NKkIEPTVtgWwiqnRndpERxwuqTxx7u+/ndvtAHWHKxL
xU+IAXuCF9X6BFpMsFeiNNACZHHUkRKF9XG1RDJfR/Qku8pENL/oIFDpAk86
driEer63C0Kn2vY/XvevkBEUa9UHGIbOUTNv41YDgJPWjATKLj2+/jcsMgwT
Iy3YmLCKaaISG7DGa6ClFGDauEWDxXNWHa5Hb9bXdECL4ClItT8q4yPx0Yvs
k+SNTg424OA2E6Z6uIWU1FjHCv+uSox53RjuLx4oJTHq9y7JCyB2QNnmXsvn
eDrx3vYZT153YwSctmJd14OUPFCx/BXY2oMbkiID/8KfT4Ku0aLVPF3f8D1/
n43Vc2GMwxBoKZ7J70HEAeivDNcAGtQP/fMpaAKWn3Z17qDgO/Khfyf4q+pU
o/iRu4Ix8MWEi4WeP/GwbRtYVTnVbF+moMmG+y02QrbyRsp96tAmP4NkMhGa
9fdMipiV37bLFns+KzpsU9uSaa6uuBF4FnoI9W3fg3Skyl3Wg2eNaakXuhTO
V6Oum2TOwxbVNFt/CwtHUqLA7ZHcbRog2ENUUqSrf+ILz6hxDfcdtnz2cLg6
rIFKhs9yZF1yBlXSrBzo4bVncNbvVs1QoVR/AjxHbzvJymUpWcsdvFOcI4hi
Y3ABMP9JM/OgEn13JKF+sTX9yVI3xDEhpc9uPbEtCmAhwHkrA5Vk1oDZygDB
nC9WVJoxZRT7Kf5mxTgt79/H29hleiwXocT2mS2rk/tc2OSlZ4d50pnEkQVI
bmrAfpbdM5d5vPu+Mr+0xpVWhUiDkKWicOxzaEULdJEodmQQQsxtfMxMaup4
zOnck1ulv5Nj2SypxuYDhTtSeGbuTGYva7v7zlCRrnCrMb4TD9fBkIsXw2tS
o0lCksWlytEJ+I9t5b8oeUuE7fWZpYaKAtRAsYpDRUK2BeiMiCuB1lfs2/sK
168e80VU5dAuZ13r6zXA+EPzOFwiUQpV51J5Y5DiM0I1HpfauH+Rlqdmth3K
bFX1eVRdOC9SLnw9lrEjxYHSea9dLR+KEPhjjG1loHrTCUJ/s7pfRFATJ/mm
6On4OGXMmXFa+rm2wSrNcTu3Q8+VmB9VsOMVi915u1NkDnr8NTj9oS5m1DH1
SlRbBQpAs2MuSbc6aIWTUoIR6q47Q24uFJ5sEeGLKSdEvgzGYGATYqvARYhK
NIVQGscP0+IIyJfnIZu5RJjRlQyP9atIaPdAnobkMKvnrMehQi8aTCqC+Ex+
XjlEFGdxrU7VLpWErl29db3yIKtajifDOXJkiSal1xnLGu57Eulcd3lok9nw
NWZc+qAKfKxSQNgKUXb7yK3+GV63OTvmiqd2hHChVztvJjBOx2HXcTRz6VB0
YtraJ+wZnndURXbm8yMwNVFrPi+3QPXuKlPRDJ3QLI/VfBwYdQzp2we8vspL
C4ZuCJPAGjiDzfAk6AMPzoGva8HSmPCIXbvLpd0EODPsx3YbLijlKuO8Yx0g
jP1dcYBFD9Cu9DP8mSCJdZL3j8dLed5lfW9U97sOm37sRoXUB+rdXMEa6O1S
LdnScO7lYjLhdDc2L/Xfz7Ln4usN2Ej3aY9OB/zTbSdIlGgO7MWo5UeVPyB5
c4FNhzXEoUjKCxj4gzBOBBeio7gn2DaOw68zb030f7dmI5bs6Q+zNvfvTvaU
fk/ZJF6DyrzWA3a7my4+ZcWDBUouq2XFJNdm8YKQzJgTtVHh7j+s3PZYv0KV
zmq4ouRgiUUijU7aSWUdpIZrYPlFqI64Zc5B7s/962VUe+FwJqwuTjiXxY/U
GO3ggcQj2NYDAtzZCUy9FzlgsGkcYRNUADUkwE0qH3Ute9WXvht9FNJhsjre
nOe+SBZlNzS/ikqrbwjG0QpuiQ0LAKgQsNuhY4L9g3g7fXmh3t8iJiyYWnIG
Myc0+9s2d+wxZgSatn+plO67LVFqquconijQLoxmdZls7ceApPGtwgI4Mg7P
Nm2RSLBrL4q2pg8zF/yRzw/Y5AjTZkFDYbFFN1bJWv/wlyBC8/DOjNABFkU9
khYoMpVXPf+14bdyHhRuXEO4XfUveYhSeU0Bu3DxJ3nPwIalmXz74OgVr68X
PT+RfZl33Nsg1UNQJx8ig4vSA+7KUTo4I+TWaDf1dcUXt5T+UOO0hW8lZ2GC
mfINt1NtlhslcJ/+pSHbhBSpQTrp2Q+S5ID8p+V6S+NGNZ9JhAMMkfILgEk2
8EpRMMKJPj4ZfhTMiSKdV6+3TmkaQqPWT4COilwfUmzVM9AiEypP3jaz/4Ro
nKtUjfdcjIXdX0yoIs1Pm1bN/sXVOJX0ZxQUQPudWAfVVjwDZrNrfj4Mj6Z6
1FrndeSxIJ4KaF8SKy7hArWu7F8gL+PaLUb3f7NkbOLON18YXptiWeUiZHLr
sWa5qxKWQJRLwfk9GHoTl81rzIPlhQy34mZPQsHFbFQPz7hUCkDHin4dWpUa
zwTTl2U4ytZ/vu8TvTT1BDFwjse9Lne+txZX4If5uSls02OphcSKeG/0PC8U
tammKJFLhzpKIOEMHR1szTIHeTl6LHW5F2BLeTkCSzj4QWELvVcySSuCtmEP
mAGDbZ8Ymwr/qCjGu/uxRtBJeR8gWAtWl7nYnldTLjP/LB0laLlXyUaabbVq
A/Wh27tQaIQUDzXFtijxZgdLNKue+mmDBkUA1Kp9/Ic57pgujNgnfauM3AMO
L1neQiPKSrCmai1lRboilG3TZfUFlEa/vnhnbF0lOMYEj0OqMlcA7LlpBoHp
iaJUy2OrPRfAfOM+EQdZzAMjH1M0c4zTEP3az0ZVmV9G3vX+4mtTPRdYX/EI
K78PHYGZq1x4V06CSjqCOpoK9LLewZtlm6FLhgdORb6zqWDcPQ+UhDGLXgeI
XJedI9TMUgGxm4DaYo2aXS+UjGnHwqcf80flRpdkdMujqlslJc6PJaUlZbBo
v4Qbnj5JPElajFTCRPsYFRHz1ewEnBNBUN80aKgRnta4GOKFd6XTBtB85qQb
rXytVmzh9AuGwSWuR0Bxp4ee/sJ5aZMPP3/xgQwjZD/n3NRu/jgAuDZ4p2sj
yMw7WP+79nA0g75UXLOxwCaoU516hodkHjm9QV5HiboHeoc9e4L4j4E1HXQb
/pwehbd088sHofs0FyOkRYjosQQhHpJPuT7c/EEK8syfcdoJ9IO4rlYOv7E4
9KgfKM5qHrWWtk50+m+Ldbu0IXF44BkS5P3jVz2zRwyGcUiXCKFNSMOnVYOS
+BdqXvvjc5+Ib0RvXZq3+uR/KYNcWBKzt9L4O3KqTtMgGDUlzHUPzV43y8tb
dwWcnLghCGvf7t+Vkqu/4la+308oxDKnzCQNFuzgYBIQDNtdMvVSLdgf2UnM
Y2EU/u3aOTXR0oJblL0Z7lm3Bit6BwB29wlYYQ/hvqrRmcUUW4JFug7EgS5r
3CRWTT5OKuGctbPEdnGLegH/PLPmkC9phFCYBEoWqRyhtl/Yz91TcByjZfEL
WiJ35I0Y6TgdAahROka6OyLSAfnehR3AXYoJZMrrUMDTgDDvtIXx4CeT4Eef
KJ6Jc4eNwZuFUtVAjgsK5kuy5F6UGyjdQ6WlWB0P+OjiMFVjLgeVZRkDH9EL
6swII5pT+zaobe0ZcbjE+jtINTB2JbZ8TxjyiC/DoncNTg5cRpzC5ZReWNvI
+dyVtQmohwrZxOwS4FkR61dcfWzGBfwzBrnfExu0xViJOf6pv9CzEzpiaA/l
5AWmxKuPlleIakQN8TbQT5xZwy9YnKfDvZdblvMoa3ktx57OBCiZOooS1l6R
4c0amoQpMUL+hAlTQPQwvwVTYjwzcyKBXWW6h61lLAJM4KxhOckmot7zn+kW
E3VPKwp2xGXXhzNlXCNwFIUQNpLCaI9IxpvOI0YqQgBAbfnBIDBZVJCItkJH
0oeEnz1OV8Z+jSW7IDqhVD46tmgw7Zvxzl8hMlcsM//P77bDoP1sjJQbTmPX
hOKjiJYMQhAqleHcKFfjBC+baOhCbReihv5bwRRU/QFEatLmtnDQ8/GnKd/0
UuEaVzUHmC9XAoTzopb566yp+oWV1yJWm9nQS64vGQIyjFObCQOMDFAWArJp
EsXSknvRHY5x1DS9CqB1WZVZACJS/97o6U2+C0Mb/ufmS1iDQnbq7NJ6/01A
6G95aGk9CTykzkuZRVSfV5f4nVdXq1d5NBo5OR7p8HTBrINh7Q9QPwOv+RNJ
Qh7Tl709UwsUpaaLTno/Q1KQ9djb4Gnfpm3u1DZCo/ydR5r6khAp8996iCxM
WaqE4GuyvjVUY+F1NOl0+PxWc8WeqLMFIdpZUvXV+3JU5+yEMxTFRvcVmLEs
1rqJpWpLegOrKO0+IBVhYZCGx8OtGZvnCndSorn9ZRQ/rrwCdb9HDeVClwlh
soU1/8slwfUFd9gch/KlXv6FzT65edUPn+hdTrenklZSQBGf6vnGFYkCYljM
eAL7mdzGdp8cSnGCp+UXw8b87objnplQ7gCEm8wLiW+oFgRik78P+RAO+kxk
PQmV1Y2sPQQPZzGjQIB1Dv3l3wKY6lxZiZnfwvobF/KIeVGWx2Wv09M6ZrZD
FVEs4BSSU+l5p9AT4KR+3sS6T+8yBDVc8rY9Lg+jfuWQJUWN/7Xs1D6cPD1M
PNPD1373ozOG4W9CHhW3H1RBva54r8wi2nYePxt7Teoms0l2Wo2WxcJ98Ikk
4hr9EAkMhtmYuS5CcxqpftK8aG7pWeAN7HBnu1qYdqQ3VdY8Pdfl9aWQp9ww
Ha+l8O79henq/vRKfR4Xn2nM0mj0hiQRrmSE04kohpmfrb8UWhsLUpPtMECg
Br0y35GmB/H+FQanJIY59w9hXaERGQCrsXPIFPUprzssn8jGcNS8Jlt7vG3U
dKtEhCy9pRSje/WTPOGI2dIequoVrTzqUrq/IuEVLlfnLHVVLVVzGJ5mcJv+
/gqiT/UxWjEuI+OIFWLRZguKvhE9qneRGC9l3/TMDD4LP/kz6qLImC61BcSY
sbHJ+TfmE9vdrTtQCAf4S4YnJ1oD0IoGZiCWrZtYj2MqYnedIJIw3uEXojC/
H66evoBcG+nb8qNAwS8nmvi8AQ6FLZapMeA0qx6kMUX/vkxuLqgKfL53jLI/
vtJZbUa4UBYSfqf2HfJ/+FkmTgqAF+CIW5kIm2HtqcgXOKjBIb0/s+GxqOCT
Zxe9q25EjD8BF2H5MDQgNG+3+39ae3YrpnIXSmjWibPwNfpo2pqH0aNVb2JF
xC/jwNGOGw92ar5qWoZwA68+Vu0rC8abujjMr8TVcAzSYb+NQb97bW967eC1
J/FvmHf3N26WDXYzVALncu6Dbwo20HRmb/IYTCqX7mcB1/MuUakAMd4k8e/C
2+Db3wlczW/64pox5FtLREYbT8CEhAKzUlJgZibcdE0J5V0MbvEK8I2DLHO2
0ZOgqkq+E29Al+X8GxvdsZtNTiWZ0iefpgwAN5GKBR+mzcCwp9Wf/e6pv+mD
+7gUtU/NdypQiKPf1Yt4OZiXrfITwURIieWXw6g4jBwVVThYp2m4JAogvMbg
yrplzTUwep8xgVrUQFij07XTcYr9h3MotP1W8KcxfMx41lj+gR0Ydmx98lOq
3/6CFp4xbW22Ju0wVSSeLX/S0tyN6EQI+8LvP7fwvaWuR2PMJEfAxNs6Ovxi
FE+z1q4N8Ic0by+hIS0ZuiEowgWcUN4kEIzC4thFMqmg5CwcdgzyV54dqDJ9
LJIhuqeNfqFy3LVAs1wRThEor8VkFi3MXD3ydFwqOSnUjxTcMleTBVkehSyH
BYTumxA6fe+3rRzE2Yx2u2u81SxvfRMurXuuoqRQ1s68DxsoJfh5YfSvOZwm
96+cStmergOkMDOfpyo6oG/OW/iO000SgQug6dGJX1GmIikHvTvo/ONjOs88
IJHLGoF1bmSBgzE49vzvCJ/eVsLgQD6CWnEeS4v78bin7nZIY5KiKIvxJyTD
zcwtg2nrBrcNJMgVPCzFiIJHwza1QlPQvkcLkL9R1QqQY6RREyy5E8ST4le0
jPVdqrB82wgXGBTbnReryCuffxnbhDua5/8Ly5vjyhj6z1gZuf5FNbA+PIIj
rYG+UL7OtZU5j5gakCTRTtSnlI00Q9v2HghtWI2EI/Udwn2Gm1sFiLip2aeo
5KAn5pnyO5Ljtx73qjAjjFnTSz3izfa643ZaXtjG4jYtKWc7UWvD8ChYS9Cn
d9rksgDUniQrtVni2tMOkprv8uLVRMx6OrgFGfgoPCJ+yvmi8y5MAdmG0tmM
U+mxEyDZ9rsY0PVKmJQVidbvgIsdeKVKliJsn4LrG22HND/TH/3nIwxLVvYx
7bm/EaHyiCr3fcsmM1qXzbm1c398Vy6P8U4+Fn+UHEaHtBft6yY+Lb+NpobF
GeINxtXxLo68M6/swseOzMleCYetds3RVqCDDV10X7hTHBkTHnRjMsheoRgV
YNmT8rjuUuv4tmpT4XNlmUMr0BhqM28A1DOcs86rH/of3aSPAYe5JBnrPxad
KvxfbnczHvbZTR+6fhwmwt5/4ra5HZf7YrQJDrUjK5dRZ2Y6lVwP9250Y/tb
pB2Afjg8AD60nXE1gZZthCxyYxCcG/pOmAyfNMXmUrOw3S+pwazrSpwVFYkn
O6Kyrquz9Ov9mZOqY8ODBtKpuZo+LIC72oIQY1/iF+D8eRfZ1HBrigcWUMNA
yw8UiRH2kmSUVLZq45FOc8mN7WTuEnFKN9MvsLZGah7SxWjnfOnkD4mo2kfO
kH6i8go+evw4kIQp//LuB4pX52wjLdQOUTgNEH3nEWfrJxf/SBUr18hPGydy
voDVmwjoMH+1CYtSbYgZ3Jwbku2Z3+tsen2j3TohA2YOKlz1RMTLVYsbEI80
+m8C0h91naau3dy16I27Hr/Ya2gawH/jJ7Po9WrK5pd53/K0yP8jv8s0F/g/
qnNZsdxPJSllAOixRLcYUuZEnx0W3fSuz9rEn78bruvyFYAsvDvbVUBnNuXS
fM5v6X21u/AEg3dTBs5DmOu8nb34nmNTVF3bzsjYgaIY86c1WWrRixVnJgZq
ZV0e0NHCRFm5gSFFEBDp5mSnnbdI9hrZx4J+sfbcyOuDmqZTAZ8W8hwhLocU
LZFJtEQSJMqFvhXu+9WDGBJfOagyB2+//6zaM9vAeBE0/bYEN6UG54cJK7y/
HaR3x1FHcsLvJncXrceh94yI5gXQ+SQnek0iM6nUI/vP/ie9pDQ9NOKLl0Gr
F175kdsHt60Nm6PL4RA92v22qYkazRD2lNiMhnGsOI1Pncb1Q+RD5iCX1kmQ
6EO40fq0oURt/606UtKCQux7jYe3jsA0Z5SzfC3VhsoZb1q6umq0uqP0x6+x
SYJAiPp3JOPcFFLLJPLdDDU0KwLNwfyNcfIFH8oa8trI8NFn0bBpk9qlIXgx
jrdVBitl4MR7NkD8FIbdqvVUBEcO6AhYGjBGXmAS2qxGhzmv7EEHvuGd6D4g
jcFC7yagQy1yzO8UKN5ZBntWa+aUDlAAKrX8pnB0GvvgLdh8uX9RgOTt3wgU
P+wQMlWTwnarb7dHLDr+AsAXWUsmswvfcOjFnddv3TT3gRFtVi+1mMdiCib+
nxmKyrGG+9BwJI1+i6xMshNfFbWVh2v4pPU+Y9CfIRtirRVxwcBdNc2k6veG
tZD+GNuCCIcPtnq4BQ1ugQ5TsQCndf2Tw/GNQQAhgFQ0p1J5z83NeNoeCEBe
J4oLVWkqSVd854TKu1CEi+rVON9pk1bhQZZnzKDfzGPRVLfLqTIDUrQnqtA3
5bogrJT3DjrGOuAvZSrSHm/CY1rnik7SYKzkza8qVRdDNwZoMORsVyUQYE6l
ia2Eu6OrueL0JHetJss9R/p8jBiHHM5CjRw+lkrR3lLTf+hDLmIQH7XuS88b
HE4eUfz9X9eNZikT8srujyr3SD45Lw8AQq++PXVkVYoTkoBNRvOGYo1V0usV
mJ/h4mwtl9+vB5MyqRQqroLKQxWSMpVNnLrsqS90gsE90ZseXO/KjGOTUmVd
NR/P4C8fsMm9aNPwkm8+QuHxisy9oDE8SvPRKCc3u64AFlZJlCYFuW3gGXY4
IyFoTF6XK9VOREX4qdyQr0W+ZiM0ls8S+l0hBPb5t/dxfzYC4uLQRRD/wsjv
4+yDaPEj/WM+71dw4iMmTyyCQaQbVzPOk8DAUIPgt5TgyRCrAO0lD1hWc/ko
0FYwgy4FsM4tJsNVBu2GJCUiJAWGXWo0sH46X6FGzEizx01F7xyb0ZTR7TT2
NjjZ5DWDzrkSqIqBJSGkyE3pkdsPbO1Cj5n+4p8YRfdkCQLgvnwRZ/KsXelT
QYlO24nI+qlHA75g2Afk5IFDPoZvZ4exr9KUCg5WKYg6xZ/BEafNFX7GCq9n
fphhDf3izlF4Uija6YENPYvTRp3PXPP0i8ehfFJJAKhws/N0bEvqbracKN+O
AOeahne19TbqvTuk21aI8rWpEKvRYqxpGlOCeCiywaHoY+N3jCciCIVl9dGI
Ema5qbt+lZNczWGmqyUaL57bTfPMgPE/JW2uFRy8maowUEnexLrqPBs8Q+dl
tUdFIAlmYcTD3cVXJhx5mmF6sdFA+2FMMdQayow82QW2TPpgBZUh+Vx2qazF
1dYf9lvc7Ctz1X3Ow1SWVnRJFaldBMXPJ9nDGq6VFg+tIifa8DpKkW2etZFX
VwDMAC/wD/ta9BqJ0oJ9bFeUX27whJD7l9ar335K6Vg93M2F/JRNX71ORTJA
+z5i7DBP3CelhyspWAfEoUHvFCuXADbFkTm+wN98jQ+GaAsCkxtlZyC6t2Yb
fEBenYj1nhpNgyjkweVSfqUUcrvtv/rPFMxYsVn8woJOaqubhwqE9KNOHAJX
6NWPm2s77FWvzsz4WQgi0OKO2e5bm0BCh0zyN6XNzIw0NjkAupmnq8MZfF/6
JqM3pUe/eP7OCSaYWVskgjA6NWrMqivZyM9EA87VqVfqCLFHo/a+szLifqqI
tRi4ikreaVfQNLoD0b2prOjqx+09xt+hw9UwclAZBN+AT4huqH8aVfHGfEnP
SdN6PIMF1RgaXgZFpNy2Iy5QjO+x827CZFfi14bIuypAIjQG0YwJLfkyhdbF
k8zbPHQCdOkd6kjcjZPKj+up2fCt/VKsVhNLGL7Z4tcez8POzWNpj88JEhsa
CMXODhq/iteKOATpUtoBG+fdqrAtjaMYnpZI82YlLnECaZkGBlvSnNyclMWe
3ntuSR69Pj1KX2GzzFrXqUOcChvInAPyXiZyKy97cJgwT5owXbwjpoPVk+Ul
LveHT5BHyxlzFgRAdTHv6lfz8xaucnVGd3o5LUdvqa8vNluQ5TuQ9Dy8YDK2
uniR/YPr5gHOWtRjVDRGrTPxGvuRZoapJFCAa2KkJiSJnUgpkCp2dynHC32u
4ZdEuBpVuKFw8e91MTOxjUrrpsLglxo02w01Fitj+5yd+taOAV7bQvnAPhox
/ENwPRnAfkVpg0hpmBuuRx67YF+2EtneyybrLpzMVMQATl2/mNEroD5lBYgm
lsf9KLe+FLzkSb2KMBQSCU/EIlvyIMBk3Pu8tkxPo8Q0zFWsusok2Vy/XF8w
Ug0SW/ht3bzIiagQn++pj1aocnSNezlO9WCaC8i0JGtqV0j1md0Mc/aWJ/Y3
Jm0rMi8X4TVUcYvmummll7FOXMe6pYff7H+VMlxJuUzqJRKAcWbCgaQYgAfI
B8pJ9diRWlSwuDIPdaXVpOfgAcqZd1Q97xBKCHFevmSNHsS220wzOnJW3YCG
IMyBOoWoAxKGOLKfk3QwXRhccA0AozqIf4O0DMuNvh7j+oxWPzw6SCGLO5+m
Rj9DsNva4GnjwKnUAl0q7iQr9rCVxOxDFJwVF+wuCLZk6Yd5xiYeSNSSmB6W
NegNK64KvY6U/GB08w41/On+WelYrOeMpEgo4u/Z+GxDrRlV3tY4ExHjreAz
Yr3zS5FwSY1XpbpHoGkBQRS1IP7fBOol8MZ8FSfs4PzXGjDcWcy6EQ/bOEWE
qvhIp1+Di+RQQWgpIlEacDMsiifZlskVrWd+SpeoSAJikqm76xveWc8ak5/z
wnlxeHWvC7ORr07C0AFNS8Q10bnkcDgGjxeWpXmG/CmE2L1aGFc4UYgkmXND
0fKkDtvzlcXmraVXWTv3REmIgUbE4YLjkZkWoSsJ3hEnTXCGZZFPM/QWTSkq
yIXcRWfYZIALd08ZZcZHg7ggT7DgroQd5xqTyIG375jgVRYFJfLHNOYY5xPf
g5149/MQthE7LCGfC9vzvucJ9C4ugXx3QDM4T82S46dl3EK8MAOMDdl3FMHf
7DhufgUVpeLqob0bGh/vYIR7Fl7OVXOO0ZtKQgS7MN63HrNi3w0t9uRgQLLq
9qLRpg8Po0J3rDzF1+l31KthgFQ+K/uKfPDfErW+JWTZxtP4K8NYEfXm1C7l
RMgoyU23vHShJNbfHW35pyaS45K7rF95awa1X5TBH3Vm0K+6Wj3qmoy49Pfz
+zT3ZZ8dpt6jGwJ3+O/juOUatiLrrZp9eyiYfZ76IDfTDNjcj+wwxyfCMWqY
0/Xs327rnm4aUNjv8Mx2VqRLaCUCSMOjOEw5cTIJCEzNKp2fBQz3boiEHsXc
tO7KE8y/rGOVxOZPviYSRguFUuyHsYb92WSfikG1DqtthdKWjPrNnuHVIy3D
iFahdEH9bL5BinxO7WzodU9rBFzCnTqTer6rEAlTuhoPaTLq1LHf99DLNqfZ
WryAtQMXmU+ygtwJqodKXbYrSTiYXCRJkuxOlikA/vw2xhNlp39EoMQqtW3O
YocjBFQKNoB8Iw2TJxRNZyG6eIKXhYnq2jhiZY/QnUMv03jqHeCafQSAwpeW
LlvyncPG9sYe6qQp7w/CNfWMudwQWRto0lxKhMYix1Hr1s04izlLXU3DZspH
0EWuC8JwttJwcZ9ZZbPrztgmpBynhrHjXHTuvjrNXtFWR4azsM0O8HVLW7cJ
0Hj8/tSJp/3cU7lo9/tXrdW0WOkIvA87XUKbMwk+/RD4jT4FeFeNvUDa/ZeL
6pkzHMPKv8MRAxteQiDnGu0YkEJ8m7PUcSUUnrZEFqXh0aBVzWITjDZ2NQgq
UbC0Yvh+BL1xe2btyyQOo8PLcB3Of1cMhE1SuqLN3XFINXks4r2JV5kceUYC
TdV9UhEyTxu/afHrStrUosjSoWqvNSvozd3K821B6otqJYi34+gjXrv9EXxd
xd/r6/8SoXYJmvW/2NMwpUzl0tp5ly91bqZAVvcDtvU+ghDMYZZG2uFYDSeh
Q7YtpOAk7fwEKAV7c2NjccII4gb/xI1x4viets6M8+jlFbYf8UhPXwsM1UCv
i1v+72bk+Yo2Yjra+zJ5GO2w+i8ixYgtaGy+z6TKwoes/3yKwui9sePhWZf7
+kTWzY/B9+zUQsuIAYKnqMG+E8T8Sqzp7UySADxdSDXArzU7FFK2/8kP3YNz
FCxiP2LJXfaApqIKo/F5GRdC3Hm+bTenrg1UuW/OIoQf+z/5L6Edc8AkZK9w
bMkoWpT+lHCRAmj7t2fo6YCmayhsPPapvmj5iPDRrR5UGAPTDQXjCA/tz/jJ
4AF1lf7GTyiWFWYfNsXvx4od0dH+poQE+21uQFo3cgMLJVaXZ2wBAI4/rC3J
CwzIzrqhTJGAXKvxYsHNQBM4tWzxKSF8EdBi16MXZqQZ9RXcVccJDZC20Uza
Rn1jaiIxPyZPECB+0KdUHww5PL42LLwEyIr97ONgHPwjwh8gWUXwTtRoobeX
NEOjnYDmwikVh3RXssBphirp9xzoyFCf8rz19sw8A35+DOENitja9p64KPCW
7dbiERoC7eGIwIQwjA4ifmMjNnUSPQ1IBagKUaPSL4n57CLCizOyjvIDiosy
yUD9h15SkW13RfXMD4qbXt5Hnt+59Q67jh1pigZa8lOIMkHs0llkHXZpoXqm
9YfzI7sPjtaCg2GlZi+6GiSPmex3YbN6ilhQehlGVkw8EKxul2iVbDDP494X
nqP6Lcn+UiN1DOtZ+yf3zi8M9pzXXKYmBcpacTm4lehc9WYjXKg2t8cOBPQe
AvTOsboOXLtIRTlzAOlQbC/kiW8fehdmCwRLporZ84jYo8Wowu9XZ9N+Pf8x
2NL/nZls+Cz8DXd4YVMU2pLGVciHYQ2D9WpCZBTtBXxfnWnCVQnhjTw32/4U
puuhomthb6KEPRV8pZcQrsYHhBEERejEYMEj0qByl32w9sLviwDWPKhl+1jS
lfRegKxhmUlREMkALJxNKs9kK/nRpuEZwnwb+kjK2b4pfK4Dat6dqbxAgjgM
MbEJx0/z01V421Cqe3n38APQ0el5HziXlLqPIV0Wnc/eg7ybQXvQjgGmZJow
spLKoih+vuXfh5Zi7F5CitmQge5znypUxL8Zxh9w2lD6J1crWZaMt8vbtMsF
UzP5rsMeHh+Kl0Q60WqYV5pQsrhGFxE6MfPLGxJMxBRn8Xw4Eu2GUoxnOjBU
M/61Rjgl9hwhrHyEULiKgU9Z1DRtXV8MRg9yrTM7wZLePC1vmrxMwcIAYLHj
zKh04WKZ0Lqxq+claHFJ3wKM3w7IOoGJ2oNFfKqGoX0ZQvo2fLZtu88kW9r2
o7QLUvdzL3/YymTrOwvGA0fAXknUnpmGwHSrVme9TdGqDD7egPQYDe/g3b8W
lb1WDMz679iDH1gLQBK4MCENP7lhIsvnSiJpqs/MAXuLX/BOmwJHBqBbKpY9
ZRT5u3SsBk9yOJQSOJ3oDU4NYP+aOfQ4cpuI0Nx+5mH+OhxaxM4Rj2GQUi4e
fvVsRAndQQj6hU1/GWRjTX1U7HFVn0VEqb9MOQvZTNIh9ee/XaDILZxwX0/a
eRmvD+M4blbVC8tyT8K7Jl7/xjlJBqMY8UQrXFjNbp8MW3ERysRzzl/C6baJ
99hLR4hIhSBX7lvNEuH5mSJvsJFbCdpg6MK0t2ocbYvlvvnWf56O/FM6P3Jb
2/GWdTQeKShvySSe2/+AGK3GMYTakLRezhwGX9hI3o8ARcFCiziZciYUMIHF
MAPzTsNUsz5qOq/5NMh37wm9AEXnKSDEQbfN2X/HA0cVKT63fb54/GZojAaQ
0kQY6ymw+bMBk2iRPYU3lxnATgZlUvtIMC2ip7+ZXhovt7Di81Id4FT+9ggt
EpEKd/2v3M5SSzRQ0issvX+LV1dRGOJ6dEnJYGKaY/kVDWY66vKodbuCPxzd
TVv7hgf+0gE1JEEd+m4jgKUiMUGE9gtpB+1oNOxqoYWcH0NfFt/qC4v5UikR
eTvMFcbC71qEtpHECAfyoRS7EDKvIacnxcerWVe8V3XJvdhdq4c6eVR+GJ6o
p0YXjFZJMzLsg7kS1hxMaPSBN0MjkIPcc5kPz2doxtbkeXgMLwoJcMeEAj2x
Alfr+/V/ltku7zXsoLgHQ2M8tk/mfMlObETOM/PA7Nnk91rO6uy2NA2qKXxn
0wS8lbq1x2QKvWL0c1WpNpqssnEk2vd47ySxJW8w1cjKqDNOH4b1bFpo048J
sD0nkvH/GkH7gNAXzdZejXrGXABOsnYAPWNnNAPdyjivI0cInBW+eDO7jX2D
s2CFXjK6jCUAHrH48SGONk31wQobyp8IixsnzTc0flobkeBsKNWsptzS0wnJ
Bu+MUkxOvEe/ITk+EdxoOL8plzvnDykiFu6Kb8jOSyLGvhjKGhoWtxT0Zp2P
8OIKJ/0T5mlh6pgtbiGlSB+5e3PExhLuWZXrbZxAEvowOwQmpQdmtOkzMo2U
pBNeRXsX0Zr3mRDDPmcaYraEpvpH8M02VDKS4K79mkDm82jzxSOqHyHP7KuA
smyzaZzSE/i07oau1MNwkoDelUkePmTkuVxU5ECVuwVgfUHgbkoktWIJFFA5
zJHUjXlLAEC6Kuxk7ml+oDX6fBUVjsgXCE9iFvSF9m9YlZ64FH6Yn+VpWeRM
qE99MWqpfDvx88b9H7UkhYZLw+Yk5zkTAu3l+csyxPF4+dlw0Z0BVMMo8Pk1
J3no5hoBl30BY29SEOG4wijY25vhcB0jAJkEm9wsr/77TAUK8UTEQIhjZ1pc
r3qA/agyXbdWdDF9AUKmW9ws2AEzAzyVOFx9XpBgkN+4LBnVgTYmEsVxQD/K
b7rqEB5x3jBwaEc+X73bAY/O97tziG3Kjvjh5VmfgFKs5sHqsV8ziYpDKr3D
uFNcd0As2PMG90guVdImqWJAW1CTxl5PV1UCzWWpaExh7deZZ/fFudl2Tfnr
224yGbhI0D1FeqWs+OoTrzrhZ/viyHbkhqoJejTI4F17yMF3IoKRCFM1/PI/
Ow0fgw9ni2thBAt9q9lDXhlkO7Dn7XZkldypfyUgXZCX4LXixbeXTAQmpYza
fp1Pd8JcP/Ok1stPSHKcQRU00aR39f6SHQHVNE7GHhPmXDkSwNynVYXW3lRY
Je5EMEjDqrbyaqvK3cRapwr+qgQV7a/jHcP8hXqavsUtKbjEpvWGn8XQ56n8
JKMjG8s1XWzBDBVozyv619whP+uXBsqnY5j1Etv8tq0qkR4AFTgHam+CsJeC
OqoSTmZinTVUk7VDqtCTQMMgSxq1FOW9W4j7cgEDx9BT8btOWIRWqwDMY39L
5V3+DBj+Gt1HFj6oCm2XUoQo8IYq76RYlz/VVj41Hnw3XJaTDD9Ufh82l2/I
+c4kg/mPlJxzw7QKpUnLMnozMXoR07sDqoIOfzT9oWgJLjgSDfxCblW3DdCn
IHjS+TDhvIfS6/R9nf9M4RHjl9En7VApq8zGI4G7TcT9J9R1leiJPH2PdGpK
KoX+FYYX6KiWD4vvdDKG0JiG9bCivpdlUSMBGaSSOmphEz/r5TBeC0rjswRY
oXEi1y2Xcv+lQsQpjmFyV9TP7kvxrkLI0NG6d5u/syBes2xpbBmSNaT+nCik
WzEheOsz3YFC+1g8zzCfXptUNS3/EyyOrjjN2cAwPEthd04/SDSDTIK8WenM
ENSKfXhfgPsNYDGj9QgaVcfAPir8qduo3iaT1HreWWKU1FAvr1jeIH/J4V1l
l52HK3JZ0n9DiBFOYru6u/wPvSdK4xEwoFbunA2SnYFrkb90s1Y7Emu71Qti
xrjU4at8BvWm/vP+40y+TeqafWmlKixr/kmggkZCDlE0tkAR0HMoDS5961Wz
XLJfO+jVIsERWNAEH4t/pWC35VFWBAaGXR0MZttpw5KNhHU97RukZ300pFs6
HGdf64WXf6UpT9SezmXabqS7mWtNLyoGhKyjLf1C84sm2fWBZy6XRJYT5ps0
cCzwcNLSqnK9ji6A3o4eabYifHHHwkRvNxXohbITlySjluSZjkrnEtj+3csT
nyKaPiLZssLmxMp0ZLeomjbqFLlGmgWDcQL5GqLvXEHKbIp2hHH8bu3rvTWp
DvVj9bOmCjeZYwfWTpRZFkgtDwoI/o9c3WlzSHkNOxuoHggpyDS/OT8cHNvF
O9/2Xh4Hkx0eNX+40OyT886FRvqMu/zVD2l3AUzDtKHRQDXBvIfpJQFi7Ktt
3Zc9aL4R3TZCKt80m4m7rwbnFeO0SR1+wCZKNhACGlpzRUw061lNTHE7tGxq
4M7kQ/BGGA8dXLxy2amuEbo/p1xqXMPfbz4s2CU6pYOphpdN3eoCh8RwbsPD
GdYVxKLxSF3Dh+e32tnnMcGcVa9CEn21aBHjZKYHHivohSwdlnJT/Lt3GMGK
qniV2125o71lxdy2k/eY4Y4GPVp/na18tSkYyN7NK3mfG/WnhcTEHPHWrkrf
tlsasfiDfqh0QWhnqOeknSY8me23K4a5n734v4f0g/3h5/M+keVPwYWZwLZ+
TKmkAKIf9uJikZm9vLZB6BWJ4sBLJd9e/t4Zs9nODBemass82vHKl3hKvWlU
+TS7jvd/vopj9CxTMOgimsN/Oc6Rpva5DZc/svN/Kc64hyV3nTa9vSmmlPtE
NoRUYtMuiBhgLP4zypdNtDGqMAhZ2pZ9Mw92PMumRhWMCUP+cNANXqDKzsfo
AV6vOndjt7dSt50pnMftN881r4iv1GiQbBZ5mLbQlhs2CCucZnw3lhofxbqA
AnxQYFP17H5+Jxs43GUGi9w8KEpoCCdNrRxxssyQtraPJGCdTyWDunJvAQQV
fOLhN32kXLRkAVNxVoMTOLaHoiU4SwXV6RtmjDqVsyeON/dU3cK9uUOrcmrg
37kFKbcAGRmjY67zvQdjGluPXGdtpQtcV6GTdeKg9u9bQHINLh6RAHyQ30fS
hTI7ywsLdw2WcvmijCtjY28Nx8nXv0n0pn0MrYXeW0ANWU84yoQP9w082zya
/rAi0lvgrT21qOPdiBM7/0nuxPh9R3Od5w7LRLqpru3XiGT6X7sqLGwwYWA5
GBUN5Yvf9NC2+04n8bkEzDs++/JWV+a1q/wGamq/lR2qRktdPw0hUH9GLkaH
m/QkBhHhO3mURQFWqoKTN1wWXZBliSZ5DQWJlh9//h+34Oz7+uuEemo7RXE4
OgTXn/YIEzUakTaocoNn70OyHa8IvHNmU+52npodDyirUcQONGyn4FRKJtpn
1/azvOWXWi4infB1JMs131FQndhUsIITBJ0GtAxXFTmdE+CJuhEYm8aEe27z
OVuihfDWs3xycIJYvpJD9GUHDrhsRsiDrN5xlx8Vocbic1DY6PeDINjWSY07
JBie6XABW4fEhx1jtll76UeGSxTyv0LWs+YAInnTv94GlhH7Jnner0IBMZvF
hlvz1Yyj2EZg7SCiD/Hhwh2fGJncbS0mc6yFovRu6lYacJ0b8AxeAZ0+i8y/
pNvS3snoVXkfjt4iXgvs+/CeeLCv1auJMHt+NQnWNaF0LACKYMsWZKInHAyz
GYCHevVHrOLjq5bB3xKLJbYAfm5SPdEdWtka6VOZb2y0w3BGLCb5TH/AuL6b
voG0+EkHnbFTciydKWc+Xj50so/XwPQu5Of2Ssvh/9r/nn7clJuMDESVvy3M
geAlsxWQ3NMh3LTg6tyZ8WXU93L7fSKVksWzmAq/nW4uWFVvcVqtqxwLMZv8
R2bueekawqh7E5Fwnw8dWF1i1vk2pKLHz+NelZYQrgxG0ATSvBv6vf1W3Hzf
Cw9Db/vhm3F1AL8C4veIJWm8Lau4ynbcF1oSV33/mWtkCMmdEk3SjsHbFu5r
xxI1ubUZ+Sa7/3/T202k6skCnTBnLmzQKDCV3cXgFsQdIwNrbZiITrKcZVuM
dVhARAGzefAJwMfOfYdpAj/q0HZqeJRYpl/A2PXRcaMIRi9ZKaFlnpi733X/
+RjKTZeTnFnsremLp034uAzwGKTGSIFTC5IzF64NpoiHXv9LimCgugUroMXt
HesD6f6dooFkjkPXzoq2IUH01ZUhwA6wdcg6PaXWeEmcDcYb7I7EGMEWZZaj
88uWJ1n7ypUi6lep8sX+UAYPKkHy/b4u/Nd62JyUqD5wUSRsVKY4VnqpaK4w
Dy7mjFhw4hh2VAiN+8QqiREJ93XTr2nvpEM5mv6GbFQUI4EGFul8/ZhxTh+V
Qw3zlTKlyJg5FleYnyJoNVOqONTdzaf8gN7P4gixOHohiBO2G4wQsCfsVdr0
P4aX6Kj+vY6BzR6hLyghOTTJYuyxlY0OANUZghyIu2DAKSor53fGUhhh+lu7
ZNwa+spGBQbGH995w7IHhoc3sp9Cu1KoprzihGne3gZA3nViDDva/u857fq9
5YADYoHardA2/UIQ4hmgivZjGY34SH3gw11IzTq0V+31+Jrz6wKLEgUzySRS
Ly/sgRB+ox/1a7bDWloezAwA5WJH6g1jB35q5w80Om5f2cwjpBI7OJ1poEpK
bfDrND/hmnbaE17UcM41Ru8fx8cnHtUKDhAKAZsjsD6jQgWipPnybBnwyWDg
GyHoyA2jvYCjVxTacLKyLEoVYc2LirKP6EuFttETEAvZInFit31Uw/OPC2ED
e4uR2fMP3zB6IudFeAq/IUvyzjs8xtRZeI0KbtDWCodtw5peSR1IVk1Yf7JX
tJ17g0Oyw0tIvbD4YeRKpqH0jdq5wa3vDxE177sMKv38J/0Bmq/nP7IOE9pi
07WWxxHXExvMVHmw/+A0X0stVpQpG9ZyvUtNIFCSYzSjmmbbTZlguk+UwMzG
L4059nlMaF5v+uyi33rGOTjNHlGms30YF9tTQm1jk/H2DeQwFmRXIgKuun0p
ZwjEf6uZX7YJtkm/fiuuLHDJEkDsqGvS6/ysLvaijzLiSt1nbdiOe6iQ0WO/
ACNTlGRcHjMtMiNKsJ1SJJDb1aPLPX34E0IA0MCe5XbKQDePF/OQ9VnLKYoP
luOoEvRljQlIeray1KhniOar/vSoSrUlM0SMXayOKuM0tS+8P+vlvBwMGEMN
eBSmSY7h3Muy0yu767/NmD2bv4DOcCF+vcbW/KrxUXc5laI0B7Py79PtvaGJ
EaoqZbKskMGW64iKXOrQTIfmmXlHIOWHKL9OgAMbpAX6eeccOhu0i9RY1moW
mtbgDigAPK1wH2zFMTRCKorl5AqjPImzPaXllr2WANKAUI9OM38jeafYm6Xx
9KpzWqcnbMaZj23GnWHZdm7pPoyiOcRlPsGGEUZByg1zSKZbUV/MLwK5G2d9
zN9QaR3mSUnEMA0D5E9xfFuOU8P8rNiNBMZQM/oIHZEZ9mgaGWUNL3hju/r7
lM5RLz+bxu2l9Mhm4zoA1Sc+Bu8XVAvm4W42hJ3HeSHe1QHFY/FmTa7Uxee8
f8HlH4uS19Q9h9/c6RVNYHrRqh8hdOCSq6i2FLKmaTPOihImWEgEkfNYm6AE
/e0hdlNXslkeQ6vhGbWvRh3uuw//DK3mttD5DNQTNINJJg8NT8FdH+eiOOHw
CBd7WOTIR9VoAUouuM204EyT8Gqwkf+1yexhnAD01DSdoCpKBGre/MTi5LpU
deEZyjH0816SI2uORCaIhw1kp22/JqqiqHkhQTrxsjwz348VzDmq4DxOC1LU
KM2VqSeDOJWJx4Hk00QfGO3y9YD7A79X2S1pzBzjWxrghFyt9rr7t/lPUBZI
xmhQNNt1e61k/qyot2rWrVVuDaKkg2UzJfzbS20H8ZCdHner98G7nZtT56Ev
1ppWkOvzGOzd06n1oB9X0wF4AciddP4ekJZrr2JB82IwbhX818qyblwNaj6V
UT/9TIS3dbsP0v2VFolWmFBGp9M2v3EdebFeT7fvXnT6Rsb93nNIbV3OcRaS
qqFpRgw5viwUDKJVf+5q+/22HkkDPLL0OpQwzXw4oUlTbDL9FSlDACshyyGr
E3oo8b0N9S/fSNv+yfUKLQ0vTmadVtaZaMj7EcZOqOdfXkUy9nEgWYX0IeJ3
BO69LOcaV+OLBFnahWJzX1jhmgmb+5K6si0mED1jm0C7Aq1zDnTliBaWLYhh
DUqFL1LU8fSJPGjJG/m0vbtmdk3KbXLj+C2blEXvn/PHI8ByOLxFeyrSVs0+
n+jcDqw5N8e0HhKzaZz4NnqvfN1zJ9JFVMHCb72K/S1Z/EC8h2bBBr5gYREc
0/M5hsulwaI0/pzY7IIlVKsT1ZsDi0Nl/+d/xYwqyC6mIV/zPBNa1JThqsJD
PhE9rlaemiGg9PLqQudGWjkl0oUPJXLK+BtRbtVLpF+q7KjKq/s9+CAx8Kkw
h0UcU0tAV3OkPYTZ5waZxWHZZO8iDmrH3Y86Y/SlzHX89dTJn5FJAudMvZ0J
uCJ99OVrQIHRVKD+14DUVbhIgY1z/bEA3jcqhnSRFf43cZmjrJ54w/cJs8o/
srnVwjCLTIf8Jjpp1DTSjHQqjFPQAK+Z1w35+M+JwLCkKUPdEdjK5yPZelAP
cdD/HUFIiRytC2mRAEBRwtBc1vsd8B8jInhiStFz7EBhIaRSeG5oFqR3DOUC
FGsAyn4+CaRsCIXAIM7G3F7hcS6wMc7+c9UNwo7Wdj4ge45VvI9qViYCXqSA
rc65VpQTK408YaRpOWu8CMkfnyJMy4qBEjGb5mt4z7GBv6/7EfPRa5DH7qXS
nf7BvzrTLELKKp2xZzsZFjA/omPCpTtFwYVGQtRnLBpu/+34m4edw0OfAtIz
gvd0YLof4N61g3y51qznPNYu58KDW5L7FapmrclnSlCwwIWS5Z3Djfwp8ONU
soCvvNLb+s287Xj7+S9qojlXocTz9GswoW/Is1fQAvzGQ9Ir2cacNpo6DLGe
eK9mfJznWRcT5RPuewoRMke1C6qZV/fOXo64ZvIJDyzRKbT8Kx1r6LE/9q3P
1T/2bq+8DPqWMpOf53a1HLL2GMmlqohyclMG237jK4zYuwYM0x/oJvRrDV1h
SUBxCSnRZkAEHtLz7sPRYPSH/BUaIlASWJDNmq5AkIAfUnZ9rqRb+0Jicw9y
jDPLz0iH0INxH+diH35pscqnaUSICCQchVKQyAh+6o+yo+iS0KULmnIxG2Mc
PmtU6WAAZPrcSSgCN7dmfUlQuvXpA1r3idacXwXPJIAZBG3MGAWFMQELr/3W
uxdHjvEAY4OZJt0uJuqYlvI3rPnJkqCFutsBJGH1mEJ/WqMM0RzFi4tFYWdp
bOYCuDL5NRUV0spo5x4kmpPQEoJHD7zRHaIoR+3CvpvYM11kMhTSONZD5Qnc
/C5Trga4kznj6tUyyAGvsNSNIwquI5z7oWg4PkkE55Yyy1irDASFe3v8jQTU
nZxBIOqXIqjDStWSD/o98Kt5/X9HRcpL2q//1vGakPyOADOz4CUb4z1tHoHz
WhBeEOUjSPL5P2AwaJLSRZ3djwfDFfzJUOByssWMS+zgoYXlqs/I9IS8ARtE
sSH8zM1vZneuLAHNW95yuevDf1NvkcT/TX6Oq+l3IpTEP8MJJvVuYY7ZO3k2
+c124ILbKNpYHmrPlV8INzXreutExtXuNJ2RbCXg04PCEl1FWPoOYUGosnT2
+91+KeENvhCGC6dNgqp1qXXbcBC4UcHDlUL6m780Q9pGJafMlViIDY25gKQn
tQ7nJ6NYaBIFVc4fE5dkXgETyb7BpTTH/97Lp+k0XdjSZWAovEC+TRRB/fs/
VHTiK4vtEL8SXPOeILHNhZOa1tOxPXGQievSuyc2FrmriCW9FyM2Ib8eO9Ce
d+ow63oxEGkVRlp+qdHQhwhpN1UVxcqqgYJz71whw2DS6sn9mYhTbxV/o25d
XDi2WlyZypRMaTLBJZ4KPJsFjAYC+fqbf8xw7w1+lggV1Dlt6xdKe1Mwjk78
rurVAGGcSmojHB3/r7+cj10PRcMOv5wwDe8gzbVu39kwwn9MwLFApTNuW82k
F13h4McNfmBdgvWXmKuacbCAaOqFXN7SiT1ZzV967iYlcEMwI3TZY9yALVkZ
BN3sFhnRnYucxSgSN5K3/OmkJzbGGtEloob2az5AocucPA2yKuxfvty/+rOL
/N6qLyKjOI8QE0HpYan5NW8QWs6FNuEymXy8gu0N7tuLV7pI/2j0wToxtMQl
JJwsDeKu5ZPB0HBGl+GjpfHNZBp0vyGnxj7yC3zN5q2Qc39CvzIEtpbQvcC2
HjDrRp3FFghfEjGk3y7n1FxEbig76ic8lklJH0VA6K9LfxdUM6KkccGAoxhc
0fjeWK8dup2NPGSCUN5R180LdCVuK7Naz4hV+LyOxyzX/zpoOI23fcjxR3RK
5eQoW0zaAqi7XzztpM2RoWI7P+IZ1smxJC+4HI2EzCZjE44P/nocQfPpD7kS
GdpKs0fhiXOVTPom0SzZYO1LAb60xxcsA6zgcpPSHC3/UMYuPSU6CqW5xel6
RrRXVremTzAc2A+QSCClwWq7Z2ZXlsALQLvf+/W5Fi1rHEPOFBcfKBgUl7Va
OPW7hUcJi9KVldWtoC3d81FzosX6dlOvQqrdZEjZxH7tgyOJa/l/1j600iMo
AIKV++85YdbHqucmCRybRoEyQU1N1lrzRtgosFE5yIIGl/8lJQO4/fhXpK3K
1NsSdRkie2re0ECxkrPVXV1JpLTUvRERfRkHqH+0wg+TOq5GDtBi9DCQYs1h
9U9olP17gkLsEFjqMQu9DWC33F6xf8F7lJ9sv1WmtGFPX8W1iRlqocU04Pip
iJycJ9E9MieZmgjf6GNNZE4ALF6aXjgzgUspGDhs3YUu+EZJtk1ecTPoyol6
M7yss1vM62Qo9lN9vIIlWs5vYsF1SJPUq8O5aduL8iSrgjcSAWbGbKLyKRnc
WwBPRABBGPzUYyX+dd1MxoqPynqTJY7Dzo1zhbYe7SyLMNNcDzOvvXpI2XRk
Dh0Va5ijBcASc4W3c+p6rNGH4AFGkuDELAhcNtLRuaGKG+SzRst8RaoJcixA
SFGKT8u63RBAhAvXieIeFgFiqerJMS1pViiNaYpgUthiD1Elamd3hGu1nIoq
TbKVXagikc71HVduMEGjO0BXr8ELxCSgO9c5FV4QxnIDLKr5f/c1YyoX1MwS
DKSayMnrrj0fH2o81sb2fmo91RmRhCoyXa5C5coWSZObIL7tCLeJxHwQY1sn
Pv/nyF2EPzgWBGEIvT7793T1bD5OI5Dm/Nc1tyc00ahTdQ7hwtdIVDA6bXq0
iTStE6wYbRfxUEGFk1V8OqId17HO5nQ2hs0fzdd/z7Tqt++cQwVJ7j2UC+Ty
2mAHtWwKqy4OGoYYSIS3dY+JCMgP0nESIkAUEBz7HHWDgSLJjnW8nVD4pOvQ
Oy3zKcAT/Py1Wchb8dJchzQF4xCyhKjcAidmAES3+kQ/bvFK0UnSAQ2BWjAL
FogMK30axsDINxyf3Q44mw1omwv9qCQW/BYm7yrFtsaue3q3CpPbp2n27GET
XTbSfI2VIlNx6PzBXratQ/0k/AcmVetoQzxpoVaYEAFCgCFz6oSp0rW+yMa0
JGcwX2LYKr7jXFB9qNp8+xQ4Nh5eK4MZb+HEmsCY+Rq/TV1ircysHXdLsd6k
9o68IlenxzkvQS8zDKFAyUOTdiXF6WFT72OlSx0YE+fp6aYxJqVRUp2yW5OM
8WQTxa9AP7mNEEZcQozP6GD0lVLPUOm9w8pyt0W5pWCQoY41IEQhEDqM/O8O
ccn50zwlj05AQTDvMZYLnyreyZe06mAHMIHSC89G9bZCa58NvrBLvNrVwqHM
lhFRl+ajXG3HUsDBG2ciIhglYBT4uln6m9iV1nN/Nl68nyfbmKaZnR3sV0oX
98rD6X05i07HXtDqQz89wvwQfxjD9mu+VlD+9P+MaATdlZXu24X65DLGRNSc
bV1Ifeicg1oBgztPn3IgMXwn0vKCSFX6lZozPSWW6pbV0c83KU5yL8w8kgee
PjSsYz0LudBwHVzfETvg1g/vnw9x4e6RYhW8g0Fzuowb0NkYZVvdgGWfR7L6
s8fQzVo5NLtoOle0mddT5zusb10REWyVEmgAlLKFo3S2wT/Tie7vgW1RIHdT
iQ9mkCGS+NhJA4LphgDx4PlMVHlO3W2R92f1G5uLWhcu3Ndwz7gsLOFXWCgF
RKJ4Lq2egSwIqdwX8g9ZLafdUca1OMZwQHEAqc1Z5ejVKBHdnPv03YZMI04p
niqDgtlyDeyugyuF+SvEldnaODBL02PmL/K7KjcGEnTNCDnGIoByRAaH+0mZ
EXVjGbhUhj4zSi3RiHCEIdZncyN8iIe8KfkQgGruOcouWvte2ss20bk01Ibb
zgWGw4PEXlYzvA4slOczMQalSMw5q4znoAHzg6wJ0DOXcPmGn5qZE1PqPsBE
AH4YDI5HBVUeo0PZwOAk9XT7JsT+ru5I2o8lkB0/fXfAp9g/Uonm/JZa7NiY
ytp67cObAEIF/f1+hGLI23qBEsG3j0fw0TwPPem8BQI1CwpG2fcM0r9Z2UfM
2X84tKH5rCjdCs9xhWZX7rWQQLCzXQDWU0+EWIIuaPhtpK7A7ulAdu2M0Z/0
eoF5JWEbE9L0LCPnFdI26M/d4043b/T+dHzJVTzIC1OprWg4VYNzW5mYLtkU
dQ/lmSJIdjPmeXNJ4Ul70HAq5XaHehfD18QdAZRQcObovH11EecigJigh5sp
X9oeCcSzVMle43+iE0UpTkvrXf0sSTNf9twe1HPj1vPeQWj9KB0FVUpiVsdf
IpnJYkyeDtXJs3JaUUc2FFzINCATXWE6xk9gJPaKxHeSaBAOC9GIWXm6bQvE
wvIGHQQ9nXf+HAlC/ZAf77hdes2pjK0CKY/wGzy1nEXrX4QjNsodrhUM54kh
eiXh4PXZWzemNR4h+Fo6dyoFpuHK+qrDfE4gYvXT0TXOAU1mA2ur4XuuttCg
xuBmZRYGyIUUm5aPb2kvexxRyx78ok8H6PVRuLY92vOLKcCdibq7MHUh5a2w
HbOOWcBtcRab/ZulKEKeJDA0A3F7tK7sHLXs04SiF5hMs4nYWGndNMK97zWu
6UWIIxhu3F7y1tefIaPn7s+Hult9bHEkFiOVslgDOPLOcTrbTZt7UFv9veJl
DZzWbOkZWqd1O6YOVfmCAeuGv1Vi0JNko4MmQuGKx4HcM+wYGTCaVsXQCisZ
GUbRV0JbGIdH41+EACfWpD0aQrHywuNUQ9//sgV6daroaseB64dDtOlRCpwm
lv9Yh3ThgyXocI6ng01FCNW1VvTGObQGNVdd7TRKzY/HP2W6KWLiTc9L7+2Q
yFfNVp1aw0sEVD2n2RSv6TuOI1qrAhdy8qd69Z/DVp7mkQUmWUhisEdRVtNr
DrBrUruGGZ8FfJUGIpupiPwdtsDXhyxIrAcrZjq5hQlCPB9jSEHiLmSJhBoB
Qt/fKfpAA8YQno5BO55J15kbXu22UYa5B+g23F3cOuxKkYHjlgcOzodPyrv7
VlvYsfakS137Dsd3XfGt0IEQIVlXXGaUwc9NjCKVtNULlFXC9yYrxbm7enUz
nulD5GSRFdB2ToxRNEAmIA5oikZSW6trDh5AQNIZ2m4ZC229itNI60QGRYBZ
5izv1bshtnGRmlHA6E+onuLg2oKhq7i5PDA3Ryj/EEO2+G+pSkgFDNVwq23e
5wJCf4qgZb0531B+XYJdnJHjYUaA/uX/MaRU6Yy+W8FCtBitdD0aH51pB3YT
+izZXwR/pzzuqOYakSaaFCog6rk2UVZkWe7bmrUU1FFsLVtWjzn9Q/klITgx
YK8Ko1C1Rvh94e4HhwSZTpkWFX40ia0jMjD4zPFGJ6xdU+aHgUAt+/Y/hTxS
8t9aj0sqbRYHzOYVTufJJ/5TzOHwCaAQAFJz3G2Dqm7tdN8b6JROMCpFHoFL
k3gAkV/6/Mz+en9gM4R6z2GHVOJvgbVyMlUtsR5I/M5fKSlHVlbdO+l7y6+2
2+L7RhQxDXa/e3F0NZdkLkKRiNw5frf53LWqex4YYMBspclwnGAeJC56jj73
xWkEcIArdGuKgOka1Kq/6TqFDAn1eQ07Pihmevsd02X569Td3HJZoV/1lWOh
AvSigUHIhB9ke06ZwN1IhS3slUWCDxWawghEAVhW1EjrRx83haSqSqq4HBDo
mJdMUMeolzG1jbSAnj+kW+69CLxUZ5K2+2uEp0MnKS9LJxhVGc/wRYAsj00s
oTov4CFvv2F0x5LfVNRZiyWxwjPjnpiIsxTIDt+FODl9QVzrxUdzjhVj4VeC
KIRl9uEDiQJBXAHxBm+gwUjP3sBgEJDpqoNt7YbN3WcLQcvXccDrihE2ICqy
oTpgCH0A6TXa1j8gVKX8lc5sQeEmalXh3fIkYYfAU7DmJSKMnhADij+6BN76
ovtukTCQ0wb3hb+r1nDwHB8xEuhPuAJIrbX1rEjLbSW5MwQ8RRyp61RCF6WQ
SLe8yn7MfjSf2zKvc7IKhPSgoS8KLHljOK9/yzGvuk7WowWFFvgzyDar25Se
eBsivH33KAmZeBbAvjcYLkh66ib28b94q14JAbf9I+WsdIjJ7/L9R2YZ870r
ScYOKxvRLw01yK+jdf6aBRsSG3oeRXlESMi+Vy1mlzfJPKKObB5Qc88S7H8v
ZC4Fm+YfHZ+KN0eVVcLbd1tHlL5jy/VjH8UKyzDbTZqe09bJFkA16RZluAdv
FRwVxdvOq2/UO8wqUdWHSOIvKg4sWT0mf0AvOde9BwxoTSZx8pWeSxOu0jz6
fmrFy0M+mHjS/M6qgG3j4iUJkpIawOFufoVROOq0mBTN98qr3EB5Rq9d9uhr
cnuuMrsgRll0/4Iolp+Y3Pm74NicA0nDLXXWQ6ZI4c+aJccI5sMjdHVOCiov
hSLTi9cV/9eUrnePApcDqVicFrnebWb70gJhCLNTPCtjEHgARkRFzelmPVLQ
dgFbdFnI934rG/yfPsmBZTzTEbOxYtHynRBC9H06jy6eMC+NYSbf6gucB9OA
LVk5fBFxPCDcptB7WcnsDS/5eettVeCe+IwlR60+yU+r3uQPZZe3IVNaDrT8
uxmlBUCzlXe7bpqCxx1POeS1hQjgCXIjzsjX39sb2KG4MTKAHPe3SWGABtcZ
t/NTHGfnFkUCGJF6kVe+2C+zlowNNpoXoPZC6Aed8EQ9KIPwQ6DaqXnF2Ec+
ecgwOA2UaCxJgu5AZDzbirFqs+KcYLfMPPh+Zy+JVGxJVNTpiX6AA7HZdkJg
Jxm5C4wGJ5juzgQjpKI1Btkx9eW+oKr/PUhmrLDtckBaZ+Dom4a/VH3kfVJF
7tPBd8XMZ2FaJCtj3sfok4VAFhZSCF8mXBT2ntKLwVD8t/lMGhBySgt3w2WL
h2/Bj8sJ6yzrG4hq2FlOMVuMLcCbmkcxbepMyj3TY8U4jxEMhuJNzT1bIWST
OH5xQx9ybUOrHLFmWeA0mcNX0fcTTRoZujGsv97owLKJBz1X1iKf0K2HXnV9
EW/V9LRFlh6hHvUGlpkuQno4OcNGPN1+ewByywoMUm5L5VY+j2lSVvcrF+QK
qZ/i6G6nCQ3KpNmUu3I3dZKXvvvcKAceh4ygTlhMq6aCK0GUXVL/T1Nntu3p
LQm7Mrq4QeP5CwXmi8xN7IXM0XGb1lFFUwyt8NC5NHZPTxMgDQib0T+8BrEa
eDvWtUJczB6ENIPLXXrlWovVlTJLq6TxAb1K4Msm0GOZH6Fw0Gq01VWbdSPo
32Lkkha2UzURGdi2+F6IHazByVlaGXzvS0owpSLoLr2x+Q5QUkw6zr07Hcty
p//ltXGGfOC4E9C3zwuwThuixUd6vVjmjMnfwLnZfKCYzi7miUxDwzmSk9I0
ga1daii8N9XUwt8nBSDTtZFn+hWv87q2xL/HPPCOgEPCusaCdLEOfCCTIZD+
eFAwlwN7ne1mdabO1FDvq+roeNv7C2gtcZgtHWgUT/2L1bhjkQ4+Vwho/w34
28W4Wcm/eWyd3PKcHvNHIwV13qSJjAAgYvR1AAJdDlZBNwZniFIzbt71IvCs
m/HdKeIIfwrL2SQyQOLyzUFr61yoptDK2Inug8FOoXAWN7JgRVlnmR1ajXbu
WX3pA0qgIJ/PsExilVQvJ4BMD8+qM+yIHcdKn2Ij+u9247/HbhHECBzXE34Y
++odaiVuckpTJpruHzbQGFwZr/jwzL078H+jS2RQ+QWLeiu1yWKaKwoT3bf2
t11pVMOWQIOg+kExUnamIqXF49d5gl1J10bEGdzNnUkBVDX4ADHdPhol2/wK
DLUA/D64iSGMEw8r3241FEP/3PnsX7WROiOkMP0pmDxp7PoWyhNyI8tac9Cj
VnLrndbfEAN+PBpRTpzIFiIcS4fSclLa7SiTbQ7hywwmRjLauyl8kQJuWAzQ
BqF0gALhrYr58A8a2PJejUU0fCYeoUu5Tp2zNou997/yEZ+4iGlx3NQe2SNJ
9RUdQg9PlDV0yCmESrYTR+X7W+cowMuoNRMmGqNsXxeY1FNxrh0kKXniJwnV
e/mTu+K8sGiORqRgV54s2SleIhMVqUzk/43+tZEb/3q2kIOsL1sMgF0xTIov
/WgwHOmpaJ/FBq9K7R5WA4OlUGqNqj9K86c3HePnAkaZsoEoBO3jEd9MSVGH
fPg6BXnLu8X/Wx8uIBL9yA+13jnzLtipQ3ZEDFHIaA/4lQyGkS2oHATOezXb
8w3OJc89tACCPXirGNwcKSBk5cZL3KNpKD8VPVHH+34Li7mwbYBTYnzsgUnp
PmPEFiVUAl0blrff8yxNX215iKr34c9pNBGlcv4trFJw0/IpfwYilfImm5O0
w+3i5KDMaxHBTaX9ULM/+igI6SGPSoWGoF9fihkKHbfaTD21zFq+k7LBFINn
WvlZiwmHxaFMJnQW8TE/oTpqfjfikAWmHu753ty6Ce0g1sJov3F7yJ2dDEYt
q+naKv5Jv+87mE3AmeGaw0z43mK8NJCHEi/j19uZVj/oNb/V352bkeA/dzn3
4chP2NyjDwv+fosbrpnBNyJkP8bKiecxc51rQQXQfGesbuwinexnOrAfperd
9GSIvS+059B/6HDRc4CMVM1DdHcf+jTHvisdr11yHTDxibItCg9o7QVJSdpt
svNVMNOiv8vdgAryksKB82XeIv+ngGuVNv84CZ0i9Tecxh4fDohAu083/gpi
1NRS9bX3cvGP9grMvRVHHpu6KVTHBHgRIRXO8tK/5clAYPD0oWWJbZEsLKNh
kGOymSAPF3lnkscT0pGVn++RGuqlycJDdUAX5ewrHyV2tNYAfCVD13bQXgb0
Gvrk/uRyM8bXqzqeFyi8LrfmnZr5w7tMwf+aRQd62llG9uqH+afih6I37arn
vhvSbJUxQB5qt94AEUUC2MVstdZo9yGpT9ysSyiqPWwV7jk0nUXx82AQM9dZ
eMxX0xySGFC0qFA2G2lYoxTvuzn3zo+xTspca2QXphT5jvMJR5l8nxxuv/5l
H0QwmrqaJ8vu5s5wDE/SgycC2QnPUTV0QFGVMjtcTnnWxn4zOAsbnpMoBTEZ
SPITXsuUXtkPwkgRrKIhpYUPEfDn0wIjhfulh7kTikLZwQqXEnqhqkPrCGlo
NsvOVF+PhO2jNJEFhNo3atxQ1XK8P6IvXNfYsr4SyHgMv/JNT0ii4RPFcIdL
mF2W6p1ydGZaJjGpySWij3W/iZEiMUtmaNNtDuzf66XXFc7BbgbD1pZgVZ1l
IUs4Hjd6Qlml8PeH9kBg5dzXxOyQSwR0tN9ZWCIDKktzIy6cHO7Oco1m2PdX
BcGPr457jPiqHDK9BcJUZprlfxnUf6tGiIk/drbZXplvLbXRbeug6n/7ecgk
yr+p2RVeVd2yMen8KTVu3tKMzykMlXRzvwvEIOuglE2ThGN39H9R1Jm/PUvN
lWNkUeeYFHfl/CdtdNCVrPbrlX99sO9moqI2UYg2EF5AoEp5eXrbR9Lq6MTe
x2j/3trU/CNGdoLeU/SH+Zwxe5ivZq2GJ410YylDgdxMp5aiZolPfVe6G4J9
EFAz6k8+QKBexWf8w4hqrkkBzpqQl6tgL/Ism9A6rEsclLAt9Mqu1RgGPXVY
zsyMrcOHt81ONiwLIKbfQEgcQ7TRu1sepebuboniXczMhz7p6H/sIwi6W8HL
eiJFbDfUc6GVmPyEiQ0JSIRCp3TsfZYChLH8uMOFmIE8vRkziq8TUMXwZk8B
Y6p4LhfKtrqpwzOJp2aG4JvkqYs37cYIpNrmvGZFhgqqx45WilEXgi6yhXe/
dlWN4lK5AZr2S332pOzTE2OscEs2NUc+JZn4PT4JXboopWxaSbagD8hQTfe4
vGhPe1Lwb7hYEEpk0KmYyV5wf07TdTnnt4UvuauLDaha6vJTU1yHCBzlozbH
smDrJGPY5xKkByqDbwZiftRPcIS0nZkzlkkaeYPi5iM9YQaZCeQrmpZchkuq
aqm9VrlJXE8jb2RUCFGbAjtys3ppBgsDgp9mxxOdsEloRFCWhOA7XWa4JQah
SEZZ4HiSQ7efoxUruhVEUhSAs0ktHDkFK26TCF3+huiVZZ7Mr4zroqgl4oIK
mo2h596Zv2nwtsqYDjOpLYMh/+fH5rKs5J3ke0yY8pnMkBKj3VjixD4CazSv
/uuJo8q+p0Tka4aYp64bnA+B0DzyPYJFNHVO/swHIaQcABdlpl9cUnlgRvID
sg4xPEsTOFpdEfpQj6G+gG7zQyaZ2Jj1OLh+f6ceyvqkbCrSo08XJUBN2E7W
9QpU7qRfPKQoD9a8RC1zrexSabMLhdf50tD7SRfvzKArUFv+0YoAMxD3ejvu
9v4PafCmm+rde3FWhgQfSJir5TNwlNmgj/IgT6gPPiozpJTh4+GDYa4vbUl3
a7m9HIoqUvF85Xthbn8ohzzlUtynSyx3iqDVZz6Zws7KDWvnQfUhvjhhzgSe
8Go8qSGRXO3l8mbWevwzPO1IeI3h/sEc6shtkb3RowQxFol08wxkBTuuO/mp
qEgEd2QDoWIlXwOSBHClVOemuUa+I0LnOAWvjLLzzwnSEpaXDZOjrLjDjD+R
bcJZO8FBPjutg6CqMrEdNwaai83oT62kIrvhlbsi+3Ysf98NO8mOToEj28vr
DRSAuueFN6e0pH+fEJaRHht8Fk4p53tiF52P/KodMb1tMsmxnC6Sbfrd7TJK
ar79Sq8eXFc+Pq1tjHe9HYnBAYFPEKtg8Isk1K5kk0MxI5KQ2fbZeUMo0Mb6
3O+ma/4Q/RcYM02gEOrccvnkH9H/PQLJZyAS5zBLpph/UEWs7rk5zpxEOGdh
LV8PnE+anbob62HIWBCuLgWl1prOmhbm7CVsFPg9FYbEjSY0fgoQGpAXH5ty
b5cIFtYpuuMm0Z21VaZNgphrFVzANqWw1o+Z+EDptMzQ+KfYlYF5YDjNJWoB
9Q7vWzPeb2NOCjPhH17fLMgvj+AG2Rt6eABH5tsvEEFMWP5Lfa5Mi0fp5cle
bEIShr1Gi6Kk+NlrHzFDvPRhdb8MmRWijHWILBleTgqpPLfZmAbz2rmY4/iB
j5uUKYlSMUreKAUMMAylemeGUlkO/rxTnURvaVRg3bmzD6YXaZwGuraLcfpy
VDuWu08dGONcgrSm+qx9ZyWqH77iIYqwuMN3uCEQj5wctUVEoo1lqb2xVNrA
bzrzzuXOc043+rpgxi+eLMZUbUgi7b24IRw0vIEyNIbfJ+3V4YgGyYwlgEPj
6D2M37gDrZwgqtxCQFqoQypYrqiGrBWmeb+Mb1P9Fg/6EjPNpUC3F4eeZS0s
XLVSm/2tNfdVGBZS+WO8ugyXZyFcOkVxM8DgkhD+cWHu4GBp77garD/QVBDV
WNpDcM0e+0nDWXowaBQcDgR5glRDD8tUG0fNfEFQD7Ut/RBFNbTmbl8gqaSc
ddPpnYMl7rlsZHHcq6mTrNXFfDfgh6FHo4uoAHrdKvBj5CmQuQ6KQcGAzYjR
Wt1XWRtAnfolX0NfpmTaKNHew2OghIX21fCUQi9YlgV6C+waGKcCT84qnw+Q
oaXUreyTqlqpBFuFEvht35nVkRS+rEF7LyTR+8N0DgmF5cdKYt0b5Jbl5qOq
1exHeXyNG9Mq3Tt0SXRlJRqYyDrDOtK1qBAy/5wTFKOiwP5rRvT5v3krRq0P
JXwzFtXczjzoV2uIuKRkigcf58k4q6GuEUFqhwOUW4XJQ+HSLxIHE/lJy7aP
IfdSTNizEfUx7GcFOGLoZBKr3RDKfV7OZFlgdES9rgWRQQxmzpzsIS/Kn5hT
Wj4xoRnXZPnQ/8tIJZrq36x3NnFmjdKG9lkfrjryWhUtk/joAO4FU3rh8SgR
oQY1Ec5Z+R0P9oIEpWMv8EjE9JRNSQyNxCrab36JiWOaOIN13/XM+OGOBT2a
5633XmWE33YIDrrrahD2/m017RyL1ZKlZiuUeSNHum06Dc2TKBJ4yJJlmJ1p
b0tl+RLh22RgGr8YH0QDBDhmC0e2GdO+e4q3mO4VzUB3LVN/zy55of1seHE6
v44EiyFrMOm/gGpsW7ibl/gKRLvnR8FG2WbWQKIZnV5EIG+EgKSQHF6JxrVm
hd1FANjD3lVMQgmPlUCsPbW69/u3sslpWIbW9WTM0QESkKw8cmUNYWsxtEFY
Vy4HJeOujZoL3Vq2aWb8A/fnBsmQx369HlVUhNe6DOmydU9sdPuld/EdGa+l
UeEU4YCOidV0vT9PStAWoUGHWcBRTyEk6jMqvLKZ1eEODIVVKr/P27HXLqTh
CiWczGlJbm+xew1FZgs0QmI/SfNpbc5F6ZKvUZLv7K8Q2lo6HkGMau0B/xuW
+C4gpohT/FQ1ae9zZMJ+Zj1cMB+B522dKiKxQoBUUGvCnHeEdgBTYrpVxfT0
GnBkQvaue1xHPJXY/0Hd2jAWC58WMC2BFgj5yQ2w4OyUXLMhuqAVRA/w6f29
L8IQA3iX/boQBdkCjk+Yf13vOS+rXxSH8CkGwOQnE11AQ2MWNyfWiYG4pW9r
mCaFRy3r5OgLtc5Nuz39XBml3EE20EEceOuQUFaxUBeDYXW4qejfGB+P4bZ9
0Cm9zAc/GAQ2m3AGMxBAduJK9ReDa82IENnIcmle0bVidq0LJ8aNA+h+zJ+c
wWIJPiFntquN3Wz/65rdJ1hs69ePqKabutt0bQEU4I2/FlsiAGWvNRW6RSu1
ZjTdLeCNp7WP5W70LiXdjYmJ4iLVWYPCTzODhRjHxsWpg1+3aAvgUqguLexV
rwNJFOPoUvI0lupX6z3vgj0KyulBQ2IWYKeDRvkTnYKkvp8Rd/Occ+BK5vYe
da0+ZHpskBpBRdsuwAmE9iGBTHBI7xlmCPuBXmwNkkIhqkdc4Rj56B6IyM2s
iQF6myMQLTeArKNpvn582PxXxrLY79RyLyhajqXnj3znkqsXVBXqiQPkY8z9
du4pFJ+EPXYKhqjl8A2hf/0o6YBurVpXQSSjBPY992PWCWjP+MLiH97I4EOg
+7fhPc5R1P2b8MZWy0sDl1NMhSUCCAEoiCHR7Xlad8Bw3izY9ZJatHqU5MH9
fxvsxT8ztdZBxYEg3oQquWD1mMTRVfTe1BXTi20uCOc91uk1+DklSSXQP9kJ
jDCUEhgXN1LgVCq+vWaESVyYZPUqvlMH3wwOOPWH4PzRu/uca5Pkvr35nABb
7GotkqFbPpzBUG9x/cHv00xnhbwYN8tiZ50TGj6xvbwkaM6094HNt1ne1mOz
c8rZ7R0DNT30+JM2IeMqizwt1ob+E/YTK5b5nHN2wwGYUqMQIHexoQnyQ5up
25wERmOV2cDsIsDa1Oyb620e8iZksl57wtXFyhAtU9HaiW+S0mwoTqyDTCDM
D3JngHX+jP2MFO2cAng9Pl58or6h1jstGOGgA7AEkLtyh1vaBzGhEZBugQ3F
vpWQJv6bLhmhqMk9HLJSbrbWriIRTmA9sozfPA9d65X8SXTGeSYWXLbs3QII
S1bu/fqAEHs0dpKkT1hHWlG8Rc5FFPlsoLxe+nqaTVCQf4N6SxX5G7x0eP1n
NMxEbdCT0TyTT+QhXsWv3NSFyHZsedsiNml96F802FE1mAGr8cq3MHBucmwj
XL28MthznkU25oqjHvDbsaGjmp/dmo3eYj351hzSQg3wDFe9GYoSZxfx74Id
N1Q3NEew3ECRh4LMucOa1QSDw5/MbKE1kC0tl2OvvPSlMPbBbjAwFSr13Dar
ZZzz6pO0DFPLnlw3Ti0FdLwVyabEyEjDd/WCHEZp68ov/LXvMf47QFfqXzMR
FkydG/9g+vV9/IylybXlTueq6LMs6LV9LEczv7n9J2qiiua52nJh6Yg/4P7v
ws4fWTjoo1FBi9xpPW+O37xDcNmszPGhXdqGFtmbN0NqVkmLC14rSvyeFPuX
axuAPsACqRupX4dI5pS6Y8C4QPp3UcQZTaJrs1zT5AiVtiVB4O3PTou813s3
fS9sAFzw/5kTAm61Zpr+oaS2zziRSgntNK1nIFv80nsMnP4VnqflPIJ2ivwQ
StzjRf87n6t1sTNpqlwNWvb0uoCG7GCgZqzAQT6ncKMR992237ss3VBPFkHc
C4g0G4eBe1mGiMvOLKtuxSP1wQgfRFX0wVFqUSW2Zzwz7O/w6r34VI0GwMS8
WLqd86xtVDcQGSrwaQCjRCu37o5uZxyTv1xqSgb+gezxdSz29mHIB0RbY2Ld
aFQ5xb3Ma3nIpPcMEfUsC+d85Mxd7dd7UU/66pxUXriK6mrqh4gXUlpp40Lx
CHPyc+c9ObKA1fh9JPonvq052fuLrsRcsUcfEhvExWXN+1NaEwGdy+WpqlIo
JSXDd1xHpAAJfXXCjxAmGqVqcqawEbyvdWbpAIzySBRTVAPaD0+geYwZiVn5
5IdzP2dUAMYyXO4qI5bk9ugJBnK+l6R6sZNxwtaZLSY9RfDYMwTcEe6cLc8m
rritEgrJREqQTeUzhQjtWfnsz8ujP1hOs6MSXMGJvFiUjulr9C9LHEJsy5Mh
Jf5HEz/a67Y4+6i+CXRwO2fwQcNFF3r/CSHezohFjm7ta27XqAmMqvBjJtwi
61sJlElITuhSNSXTIjDvGNyyTZOISl+jIvt4OJVRZIPncU8if/GZTayZD+nN
QcIzgUd4ZwtGkGspJXFqVoWh5eX9HowcuipIKgjS6Iu0MWIf7BqJy9X9Lhj5
/Cm359DOALElNrs1eK3mHwo3cU3eQimL29OAJuqJSX8YNmDFR8Ki0qVxYMEQ
7igW17WWIxpJ7OoawaCJZiydsqVMeIbMW5+Vp4OFPFwwDUgCcf3D6d4vAAO0
6HpSif9Ioa3ZO8MUHc9Be0O0dfyjr/kT/kIct0THj5BM7cDtv8va8GSbW80B
Tpj0qC450t5os5tg05Z9R25XPf87K9qvep319IlBUb+RA13FPfDJp66I2AfB
EvafhclMQULmnlnmmK0mFkfvLj/C8EteWcCEHuRMEQk/xUbpCq8Ryem7ebXI
8ovOcHZ90ZEfYP9l67KcGeRl9o/qnBi/9EYGMGqW2NILYoKDW8gjZgKdzihd
sfopcXiqoXRvbC7ZQ3YoEDXGD/ifuFGGYlCBNWncdCUziF5wKzK3mrDmhN9D
k0bUEIqApdYTfWH99XaxOjBEAd4Q2RU5cnHZZJPPkLL8J17OaKZO5bfzw6ei
HlNrdkFY2nYuGXZ2RL3k9hcYD4QqM2gdBpj/FGQKumm86YXlJit8ozZKYsqK
CefSbYSGigw3FSZGEjzEo6FtQGlI4pUC9/HCN7O9IigQh3YcxrQCCRtMfWAI
wynEYEM+Dvdbu+hNDkbCQjEYJXo7UAyla/zPFyBVBJNfRczv+sWNWD2cIDYc
5VgjjyMjbOndzAVNb5oV/oq+YbRasTJNxtywcItn8qkSHY7VvwDH3SYuqZtP
RTm+1Uooc+uaum7r60PtnPOw3gOVp1iOP6/PzJQEi19Tgwr+Z+wZ/ydMy3DV
rAlqD/fPUZdJMuefvjqhwXDHoOd0pKhbawBfNSweyffHoztaVdXRyqp/g1uS
84arhsIPvolFf2hw0LyyfqQawqvLp455x6X0MuAkrk9aMmXOTFCs/Rr1vu+g
VrmAjdI9U2JnwG6x7AcR361UqVI52gBm+pVh+C6QBV8hae66wPxWmwP2/4vo
/lD5JhbzhQA4kkat9oWtkEP80+DgycTifs6fXQykoxoSr34J8JiqR2b4dlHm
MfmTw0meY9kMB0ox0lyq/5JSYJvKeF+a+NtftZVL1ydPAQhTNUCd6z5+wOtW
VZrkszAoNCcLDGzMZzvvd1kUrCua8TrMi5PgXH0P6qhg8dBe4a9jGhEHL773
tvEnjcX5BRaA6c9BmqfsdaU05C1jcjJH2Pt7uzDckJcrDXbYBM4atsOi7CSe
zbmbICHo+6J/ohfchYm9aIoqFVV7A2zQZXoTxBN8oY9rQxeBxHsGrH6bFvHq
H/3PTKILsklIy3WCIkJRaBc8aA8SDP3vwwZzKlwSOeXBxZLTvGgytwToDUdf
cqsKyPn7c8qMzarqAOna5YWNjwIXVgj9DFCufjCVec/InnHez6N6nCkvdf1i
Jccg3dxWzOx/gEC3m6Nb197DH4fYZD68LPYBf/IpLtBRKX/wQOvy79ds968G
CWua04e54+BXQVXR7JFnnHSMOTWczFd0xkTzpB1vCODK8uYFEjmTe4xGWnuV
R8EVL5CiqFADaUj/MGQ4VBd9FdHByfyL/w9qBdnZy/DAkaC3afvHrKUU9K+s
J7pjmHS12oOFjdYV45HvEz0vsZoDoTh+Ma1r+31gezsRtlyiiH67FX0exz4V
vtkJeOETeKwz7qnWzx+BodBkJVBk4w/FBX1xodbc9g6kkQXtQND1W4MsQWHs
KKWXLmUxjxDCgt3JRHblnwXGNXVnt+eyiv7gACw/pRwIIeOl5clS7P47lLeL
0cloRWwL3yApIsOKwbjerQgepF3BvgoRvlsdRsP3O42La8LVG1zs1cPn3MQY
wPHb3Y9C8Zy0Iqf3ZAzlTCGK4JKEWnpIGL3Pbx3FwMu8lC07lxJAGwsbXVfU
x+77di8wX9ADHwy4bC6P6T6zZPWQsSX5Tu9h3Dj4eNB+zBxdcTabADjxWUfP
OOLvXr763mF8e+hZoPRShGwTKGXLrQ93/PGFFmfPOSFW6wXuyVkyYWErmzYc
bur9wNEMmdx71AEQuVpGv6Co2v/jdEmoDYrbH7bVpRvDzFfQv17m68tEDUdC
8wLTsuN8s2Eliv5OKrRzLLfSgl4BevpERla8abY19yHgNRSfP5hb3hoZxVhB
9PgBHZJVPL0DIcS2wf5xx7e+yjITqGqsE4yWbSLpSuCWWABuIDcrb5OnMeU4
UmDVTd222KsUtycDDsRNsD2c1XZEYUcxsGmiPSiOGNWKyyl7oB4i11Ubjisr
hVs0fvASpxpugfVYAcKHbJ8tgFRSIYa8TymjNxB6hUjmrv+iej1DDXMdTnL2
dB+WMs+Kk9obSR/UBEiJ/O2dn9gb7a/PfhAmZw5jSTlqSLc1xGpujwXqyWdR
ZRLakbFsQpa9vK/34zTw3e6B5+KigdqwJ2SIDurvx2/1YHMSRXlT1k4T3hxq
9dDa2xzFPZYPd2WgsNcy4Eod1rTxrhHh6mS35TOF9Fz82Lf2QVRsKpmikmeO
5QPp/uGbs3vKYzbDdPV6TX7g+5gczDiwRWKkg8Uh2G23ly1U5Tibq5U/7WOF
j9WNNB9xH9V5iPvvWMLDd7IU0rrP4KsFZ1WNXngCtogRSlflDe1ofMwJVPhU
1ypX6edeEiRVMvyH9zKRIyZb2XzUDclSlBQav0y+a9qOIsjGFLvOoiEIDZpw
4q/TA/CVdhVcp25JuMccLOQtpiuglEOfvzr66t+2MlVaVk6naPhRrEfylbUJ
xm4HXC0xBKx/a/Z80IxGKkIER9u4PpSc0uMT3Q7WYypBNErBJgU+QVvzYG49
Aa3T9Lv/lDNuDvIjGplZPx6tEhVVsynWNQkSDeBfhd3bLoeiKkJDRI8Ab8HM
AgNZ43sPH60W1b64skjNJjxOnoAzGPjc4GnkVFCuWdU5LHoUUMGBsSsx3Z0K
ZOhWhYtxThUre3hllUx++HzoPBDFMAAl9/Jvmj0bOw9Tc0VnpV1T95CkdrL0
0fwGmVSpFgLbP5UBVIZaYl8jBBlwo6QK3dp+DElItWsKLy/x4Nf2ocGpCLf8
moV4yh78SYqX+5s36Nyj8xYIx1FOyfUvH9L/wiy8B0LNKjvEdY4pC0UJ4wrV
+sCfxARttARKpp/h2ur9/uxmpz1ciRV65O6diV+pqH4HkK/kw7SKq3b0PAK9
AgFjIgHCfO4/w5LS+dnRXwLpkM+KnnqwiAUvxY3Drixg+4xD3C2fZjXRRfPH
FxSy4Qp6/tSmCjWpDi3qnfCg1YO1qzG9B1Wr/uztj6pTDsuT6U7euzj2QTqQ
UPNdMTTL9sj6bgMRqdxfAwljyvn6KTWkBGq7jU2iiNB8VwxGSN1lndCoc9wF
TzJd6SiEohq2ZFrtLsaUsY8MiogMId7oyhOEfz0iYCJ20NohX++27y3sQbyt
iJjkDaGPUT1u7YNb//JpFLxFmmeoLz7bFU670dCL6QahRhrz8SQwhMNwNkii
H5iwoEkos/N4HOEgr8IENys5RvUoVll5l3yPWaW34EF93EbYPOsqdrAC6Wq/
R0wCdqPf0ddXI8b0MuhAfEgpC6HYWcHu6T/OBxxYzZm1DiD45fZ5pXEuWs7J
QZwGDRS8tTZ0ktZVsAqefjpssxhnJOsecEB6qht99V08z7uENfPxqTNL1y+S
i+HTYI4kRDdzW6mJiDydk0ZPUT3CxFHprssHbtxXBpBkjOB2CxCtOxhnfBmV
XZt4qJM0M8hYAX9HEwtTyRspyq2FMoOMBH8t7KNkjTS5nQEC1DeF6VKXoM9e
39vpy9H2d1q6Eo2rlzMpQ0mv5WyFnYGwI7YrFdJaZ6O8Gq6938kY9X2+CkF+
xUoLyx4u4FM48a6SM8WqN1VDqDCjjJ3h9I51GLeN0Wt70xm1cC9vUdLPZr+m
4S2VLeQCScjLz1OhnIQowBJxmDdOM6Tk5eUjf83lKQq1xj9Nsmh0eNry5UsE
qX5DLXiZoDA0royQ0t6JgmsjYBxTxU8KOHF4u51dYFmDX30sGJr6VpeytEMD
43KHan2WBBy7O0rh7I/SyiXXDFlx4w3tuGjsnoVDneJ4sX5V2MS7NwTtnC8f
JiOWstpCaHGugBTrQE/cCR4kQvSzqlTVISU3lyv4XlwN6JW6+/s1mboUjomU
4o92vIQaH9ulxL9PUXgS8w2TXpmbWlzlW6DlAMerqD6yGVYclwZjKyFAw+aj
C4eao5HP4hW2jD6YQWqjlIile7DVDCfSeH6/DE4Yr+GHM2UMjCKUxWGo1bU+
jFey1E4mu4THrZQozZaWpsPOvKSPEjUKWJ+MkHk2VLwm/3aWmKxdwC6zD4hW
rwc4DFgpa476RUtX2+LAZSp4lx0qcBBDengiw0XmFoHb9HQLxs9vnbggYsNV
sRU0Dgm5ZIyWH9ICvYPrpGt0R2dHe5p4Bhrt7vg53+5deYoFyttZzUqCPBea
6BPC4rI+YJrzOQ5/sEapzRVz0hk39vR91ThS/IrJwD74b+l9qdpKMv22N9ag
vVrLkJwBtUKFVvsD4lsFo8SGvZ2f67lkf2HCLMPOK2Os4KAWx3DfbAgu6FnY
9eV8QGGawK8CR6XNWnopS+bQ6pLGI/s8rJgvL1MbpAaGSlB7QQdaYZ4t3af0
9WH6MHkj78wg387MOuaA+eCAx/2TVOEyLJ3Bg5zu1a9bfSCe6aIpdGdITVDx
JEqS4Jdpw1wIbL3zudUpy3/qIcQI2b+y48XWaWMwvS6cn6JAMt0Pna9rlReP
vn+K76uoVaptQH7rMvLGcfw6hapZ6jRGgG8OTbSml07tCQpFW9O/rUz1SLsr
wRpMZ7xlKewoTdjvHsr9dXqPDiKWuOanPX6/CEKkJIKTiWgwCP9/pLJwXOko
C7GD4pF0qIN7vMjs36byHCDmkoFwml8yqNGyCl9X6CLlWY7J7rmin4v2Fx9t
2mvitt6rABH3dAlvQmHLh6SBRkdvcSLhy1z2JLn1dG+zNVfA4j7X/rDw55TX
zrh1DDGRPTLMpSHl0VT3MRsqEDpyioWHmHLZZUZeSF5mAB+Zkbp7nUE0mVxe
nO2ufwr8OhvwdcXf9LfWNAhkrHYeUv5iR+NGvLHw+Hc7jXckXXaqO95n3TuQ
IwAhJdViu9uZ4NpXNNU3TjlAPLYRIdBhRxl0pk/5ELJ8I9Z+3hbJrwCWIjMC
JFUElH6SLkmRZp664D6z/7pjZszBYNcX1Gd/htssY6qktmMeW0arXBnq6S17
s3s+O/N1RDCR4bt2kn6Uxn6CbW3m31hboBpiabehZnBGhBnTANVbygG9xc2v
meObTKtYQCbwwIielxPyfWFuB9GS1Dhn8qAQK5H8I3+XVSPApld9GLGcxRfN
oyF1XRhuuJFHpApOdNlN7e89z5DYk2kyfDoJQkH6ltDcWy9Em9j0sT9CuLss
NpKfaD5M5Tsq3HN1Adb9XAgSYuuCc2CV/ux8x0M+3GED+x9bNHIhtw2ba/xP
ZYpEUyyGKJcUYr1tTn2S4oMxKzk8GERYbHcZzM1dibk3N745THyrTf3Ucr31
xncyoD0e9OX2PZDIABn7GRzFn9hPVCJ0AJ5stMpNgKoWqIktPlb8X7pOa8hy
KB+h3ZZwMiJ8/LDPgy/a/Xeoeo3ubzgJHfUF/e+L2tf8ReYfMFz21QvjO+AF
coryYXHwYbn71RK/DmaBCOc3dafHkiVi0W2YmF8j5DYjYthx4d5Em8zsX6ZE
ZuT5MIg89V35yZ7Jwa3bZSa+SbPSx0mhOYr/anbFdjFi80BUMFx41bgUWStY
ksRZDRLVduKb+kI3Q9PIgsydFOaEZmkhNeFdeFa8sch8gXI0HblRC7ObiXj+
yfGNq7dlD7MnMxZcgFtrQaelHCXMTmq6vqbJQ5C3tEZGZec/Cu3h2UR6Vqxb
03BVFUkxaQkgrSBNkofVghxFCdR8f4cwot7UX1sz6rRRPHB5Jk/RDJB06++C
WexsLUkRANo8UNTKxQBUOSfp+D9vnnlzlVP2nY7zJkgy0xhAcbAb8ZIf7FO7
sq1t+vbnlHaFbE7rJV8HIEALy4iamUuwq4Lna4sOJKgvLZRZG76Mw1UibTBh
UDiz74FLdo6BAGpyPz/IvNCTueBcm4IWsQtoTXFzDThe61KctQe0k6MVN9FQ
fmxTlfOulz3VOE1bUD+aVPIbzBQcx8seWem10MMkUYww8HkXBg4UBF3nfZPp
HK4gFXAwqrZE2cgNgnwwmzIO8mfzCwvdXn+O+rJgeSQ2r3S2a/7H0QPK9mnN
UKIzJXNdPRqMlYuMSBo3yn78TWoidNaBvdBVYF6oPBCeDWVTuBba5GF7wzZK
KOfX/L3XS0kL/9qc8e9ZFhc/bNhcsOC3X/tBFsCD+hLfNiVd7pGHsAEsMbmd
j7Uv0mB/ldUuEiR0Rdp5v7ysJ2pVMb/ZvKW0ufQ79eQT4PMcEp94E/TMMKxz
0svAt9j739aOeXtkd8oPs+q5Dz7jk4SFkpeLz1c5p9CAljDBQPjST5+jC6zI
RhdM9wCO09SRZccgpZ+Zy0RKhVyd2KadUSgxOYU4jp+ZEsZtDbB9mJrjtr/D
QbUfSr0ckFZ0o7IxAghZaTemg1GqQVsaNQMVcuuDCsWoJwvme776b4/o1nky
LIYTwdi30heYzTdjyWBoWLVpT0J48a4gVF/3dbsSdr9u97OcOSoCnvQj6061
H0KoMCvWLF+LveHOqck0WngJVQ3WmBnJQ1DCQ2wDms+DAD5uLRI6fye5F0VP
ST0AgNaQtrRga7II1PQ2YlDlJvEnMZxE93SU+KZE4vxAWEig0y4l1uXDO29R
G751J1RgOrxyeCR/X0kFtswOGnlFuoPcxN4BNPT+DNl/2V6U17FhmlYqJtkV
0NTnbO3jzOMwrk7AO4pL2miAtUiR2oqaEBWZ7tCwHvcsAHV/a3FGQn4Uyo7U
ET0BW6NZLkv8ahqgonBRoXFZ/qbe7B/qPKycL8wv9ZSv9PsJEmDmpaFVNksn
+zEtQ2QIPNiOsyxWEGeNL7JLIlDsVBHkmcEaJl8LJZVfX579Ml0uauNGjMVX
MN4TFwzM860h2u0i14DB/ufQvcNIuesT4Y1HFB0idocaEIW/GzbTkbT7dBV5
RHV1DKMZVV3fsGjkBGVNGRcQ+rQguzST9H4++sU+Q4S4TgystsSyzYwweboG
iIeFDTamUhwP+3gZY6buL/ISreWdIgssUMSTx79B5y7yTPK/ha2b+xTgaquv
ZL131PSRKEUwMVMr80ydC35PaswrBYcAdeNgCtcnsssbHHZI1ngSm0zHiw/1
2x6gWKr9juSVcNO8GbD+KeJLH4/Bz2LIpv5FQwMGjqezaqwp38equ2dZhpwz
49O39V2QgLwec/EUYdkw7KdkfRJLc/0X6VCogheGAAVa4mYSkQ9H/pdxPgoP
lD2NH60KzywePDm6LAai/QXjBwhUVifwtDca+/1vRM1Vdu8xrm1JpCCPYUfN
iIN73U/4re5iE8LFB+13686nTF1dr7IrfiqGzUK1TasO4vNB2SzZdyMHrGX/
08KPdXlKhgJ9QZ1aaj5X934cJNKk7XjdcpDkwzT18YdEq6nkOY80Ze8y2JqM
z4PBjWOhUKBC3+notNP858tkaqRkLyrC3xNC2rSyHAbMBsZkvF5leGwxSF+s
fwpefu++Y+1QCcT0gr1lFNA0oZWdZddcuiL4r8L882jtAiiZNltfU39RTRye
xcp+HfGnBXAhFqdo2Ash1aHVo8u68R+35lS+IYouopEYUWeS9iW+4zHNXF4U
Fij6u3FxoVOiW/oAgDolZfYTtVh80nrYvyl1sj0KPet3AWUyrhaJa9DoWPsp
bENay7ul9M8WlQq4TZULqizb7ZzfcRW6K3jpHft2WCm1UrKUf5uKvsYTb9k1
XhLvgAK0BbksDC0IcG4YkxFxXrvEKZr4V/GcqE9KkGBxS8OaRRaW18C0oKgX
qOdwtU7KsInwofnOKMdSwF4kHIhHdC7U/H5pDXpEzxgytHXzTvTY6By+9VhU
sIfvWyhb1vUSxrY95Mo19HzzRPWZaziOv6HPQCgQvhp2gy8xm/beMejSeZWD
cIebOB5SpptecE0GHj4aG4rR1nJCziCtfjvYL0a0tmPXJSRM5Pj07joyr9kf
00LfoBUMDc0cAo4zaJLDbenBIsodrfla6UeirjyyzER/lGwqOpx0ox1MKR1L
CBucs4C8IrkVzzoE5O0L6PsxXQ1fULcZC5UTiYlBqEPAiGdz3t0yYR1zhPcW
ECKNL6jH7Z0oohRYV48fV2NbhETZp5JgbU3jyQ4RbwY8u9l9M2gHRA7f0VK1
BERx1zJASf9O1OTHs9+QQJ5PfGqkjR5gZrwM0pDH9RuLZnAezUHq8SsXcuWw
veZfMXkTp6EHVGVX9r0lHpvwC442aHeSaFONdZhzwkyS/M2wufmV1pmkmrUK
+RrOQQg8RztBpZ52DaljgYULciHEm4UQNVfhAQAhCUKNIVyD87hMFzVG0gFM
LHbR0kcoQEWsJHaLmDNeFOfBhTl+uHK7TbR8QyQcx06XyAKKamt2BmmqA//i
ex+1rh5H9boTSTg9SYSsPxiwBVVj6CL6NAElt08rP+U6SjIxZIfCQTkUe+K2
NV4KK/PdA51bPGecoXQtgT72/K6LQHKWP8yRt8DUWz0AZ0qmtVlIx62ow3Lt
e013ZrvaWolhnQz7xSQwsw6qOPEZw5RzH7uG7hXGSq3GRxcX+KmBVg1O273w
n7jAL+1rhB81TtKixhGuDs4lgy4NRLS7ZVuPgl2NEB8k8uqhaP6ozjRTDGsI
PYXDUefFDQ7uf2qzC6rqx3NPoSRLQXCw9Ef1BC9YPgM/1UIWj/zb/6N0mDcT
eRgBvjDm71Dh0MsXDK/F8KGIW70bgSK7kVgxdm0r2syVCVjcAy4VaJo7/LJ5
AYp9EFu8eZmdwarLhzdeSP41+ZCVPyCsOwDUKAqAi44lvQnfaJsbkUUFYjRU
5PTE3QGc9cM24DXec4fv6uCYJlg/+nRwE23M8IXNxji4I956MgFTJJBSjgI8
2zaAMw5miKLqH4nRAw13L2iSFyru34Y2duSk98l+a13fZIiSAfMF85N05RIH
RW5g0ZOvzDsKpqAaVhgdYHv6+EWfCznM68z/vqsgh+jbWHka39eNTma4E8xq
Y+10cqTqtWXaO9/QNyADrBldlZKtf2acYWRXbIecOwnSqd7siKF5OiR5kUAo
usl/lCe1wz+gg1XsZDNCjeNAirh3ygQ0pwlw5wSWJfMs8PB3u5NUZU2Uf8wg
AfMtiRHsylZgq8+FiPUkX7+5BclEtophBGvsDpgq24Qsnj/4FRgxIYGZTn0f
t0LtOMWTyOC6XfsklQCdiF+G7G1650NzCzMaeeBuVipxOm8A3cM9pFmEDLA7
VSxyxVOKgElI596magazu7RAsqS1yL5J4kD9STvIpF0wBTJV/hTy3r6HaK1S
XSMHIjwsCGtWZfcWVnGkp32kESeOfBVKJhbVYWItnoJr2dSU2J8eTjI5FZVA
srfWRyv5yzvPzILooVk3Z7BSw9P6nSinqTqDGch62NXoGG37F2LyZYZW9FdC
VlZpLzDMFXYX+zKl0KYlWBRxg8mseCAMfRfklhyHpweEU0ZFdWXfA0FSTKwg
pbhP41rJsXSzaDuEsP72kII4opG7n0TyGYg8Fc8ZnjSTq204XrYQ80GYlnwX
jg8BvK7RTkt/yrPhVfqs+NOnRTrVSJ1e4Hmu/s4rcNfK+MKHNPS5uMpD/jEs
hsJqjXCMqAg7tcm3Vqh+BpTeDgmTcFoFw6+GGQbKcWdGBd/r35Dek88DG9bC
Ml2WTYjpRVmhmYmA2Mwmz/KzNrXI7csRIISVv0dR5L8+tPSfLc3XPKMbKUdu
i7MKBrfXd/AwhbSHQ2hOz0cvmYN0S1ZpYiILuuuBCrthbzXLmUrPL1GybzbE
5gZJ7/8hLy/mof4v6k6T9ZnDefqYZ8lZghpwwxARe+YKzxDN15+czYAXfk/h
inQGpnzcjGw8im9E9essEozWNheh6ZpUiU/TfwOaY/uPeC5MALkF2dL6Et+S
WYalMtYaPqT0Xi06lAiH8WXTioY+dWfLVfeT2QRbR21z0Wk3K8wyW8XOwMAk
iHxz1ZQtZWsRT+0q+mgIE2shcvkjxJa35k1saOXyUmJxrGQXtYORaNmwd+fP
ocNq8TeV1wN3EVXZNYXp2ivUaGKTCgm+HZr6vMmQEi55zUinOA/KKIls7+JS
ihZT6+MTyiSo3gYWCawBDX37xPD3EI33QFOuip1+hxwzJ8lF4FImD1V/O5T1
lO+dKn9M1YlOPoBtrAb4UjmiQspGU5009DKTftR9Vg6NQHSLfPq9EAexq4A2
OUzXC0UxhqM+b05RB4L3YQftr9ZZ0P3sUcdTU3eSttO5cru9zk+4cP/LsK1S
PA69arOjpDu9Laf29zW+6iCRfitdA5+HDyXL12w7LMPBfonIK5VlQKq/KSpm
7Ku5ycVTxjnoYqsCSbFlA3+7HloTyQGyCVdT8nS3eUXX492AguWUfIai1v9L
M/nyNCpMdbLssYSOHjVhE6XvKuU2qYB/NotEhQnL4OI+tz1lYRh8KUEzPgJT
W+x3jOOj2CLtlMyXQNEL76DHadroKmcpFkxTWC/ZFqN/YaLhmqLe7JYeaFro
5Dy2SdpKX1NEb2Bejihzu9VftlHfhfuyHZnJgW6VyK7nHx0SZJeRLRCscFVU
WarGNAHWDGEgEpsps5delCM2qf2Im0bfHU/0ddzrwivztjLXBdkkIpeLwif3
Eh4G7Pub6o5yFlfYZbwDpnDW7+ef3l9iEnSuYOCH8ZQEQHGpqCJHyNQS78kk
MULRjPXtMSrb9YhPAY4d6aXHzBY5ANomnSf5CMBHExkpwxo0jCrQhflH+SAV
q8SENq46J20VSuXCAVc1DLHyF/byMIISjQlYt5lWIAXOChuNy37CTl/RjBjp
5V3KrVbh/fbktAWitstd0bFimQOCsAXAP8ZAzX7k2DDA+ZHGshiCRuLea85k
GgM62qWA+Us+CvpLEWJdzLSfAXBDZbi48zSy6FpsCN3aHTOOO+aT8605JCFI
xyRisz+47XzvYo32++7pSAD6vh+6uYASfdsYfoh3moIKvb0kNde/QjqlHcfn
8IUoJREwb2iTcxdBTp/7fsQf1+xLNpkSLR8S5U8tEDd1j5gEQZuK51s2KTbc
BMKYVc6aV3dVZWhXkbh8eTa1byqyjlgJdEtDqrK18ZKK0lRteRLhnAf6zLEA
e3wjtr5Bij+4XsxVeJreI2VF6phM/uhLpRhAxOgw3rzWhp1Oum4gO+ftKVTf
xo992VBK6jyUOvLViVt3OqfDQwnbUhPz98kPkBXqXJgrd+uxzeMIY/0FWE2i
rVdsPhXpZspxidfN+PZxjzwoIngMPIOIo9c0L4gaxr8G1rgcGX+68JCsU+6A
YVlpSJlSuFyRoJf/4vdX3xaLvoeZ9hxAZXOIGWS6fVZ/rndCCGhkEyhxVe3/
+KodfkqiL+qewAEU9FxrrDtrFeEcSeMr9hCANJR7WST3iehpcoc3j+s3X89m
KFux4l8IyJntal9pYYKjVyd8ltlxHMijbHm5513StXgUWI8Q6ZHMres5FHUf
lHZUCaAswYpvpJ40HU7khSBlLF087QcQRrnfs0dh53r6MaHiABE2H7sTfqpV
J623Ah4bQkiCZZpPVUzHfTraU/rRBPjRpCuPYLNwevnjmyxYC9DtWNMRVMN+
aRu42qIB5st7JuaKbeirffU4AQ9Tal63LzJ9I+TizexyCXW0lE1oF6lnathP
7Y7NL76L0LsR5EtYsd0F/hSAfbRrN/6Dsv2+UuuXLB+hOFW2tZMqEBdfSk9H
GzJ48Fi7PK166FMSRM56wcVgAiBsmJf0gamwvZ4F/LwPEhh/J+s6U9Ty3FmD
iuvfxqEeQynXiclWp9o5wpJjKhRRb5PF2tu5MVTJ/A+hNwB6trostzxDzNr0
ZeWD3SFsUiEnRE+0rQLzOUIkKIjmH7C58nGnabN6XJ5TD+8Gs4+u/znPXWlX
PFPeZZcdM/a7rjCpR0Upqou3VKXhmdmQ5d9EJcpabfKUob0bYAU7GAKWKy8q
rYJGSwvLiOzo6DvkKhDUiUaIGKOYREhQ0owcxm+pOKJHdPLdpTjoBZprXs28
6RLZgCGJWpN7NTBtfbNa/vpxJOyXwoewshlnuSatj65MUeDdfLAc5aOkwXqi
uKB4KqZQSO9pkOJcQSB69JM/hFDYOcMDDkblLTq9CHJGpDmcLJnNUSu4wn+w
Figtz6GTH1Jd2l0SRAH0a9CfDGKrVwNbvwVK2/J9xBtwhCEbiS2AGdmEc4+p
kS1s5dUHeApvua/Kc1OLh0CvLJUH6eDFmLp2fNaPbwj0UXp04+fuRAImhtbA
zxv59V7oXWVa2URf9ArU+K0+lgzl5wShFhHblzpfaCKGBd/6ajfs1QsyzAHL
XxTPsGaSnYbzsK9wJbASyLba6ft5g488I4bwIO0UtNres6EtkXvDSsCm6DfP
zlWPdFhVZXJ87xzxIpa9fsTfzTvPTdseueA8PVzmzD16dLM2LibwMJILdP8l
zu3VcSkSBFOcJrHx4cRObWfv2oiNLYgYKxtRUFXbVVkn+IdZRX+32N7Tdmeu
P60R81bPZGrCmu+5xvqa4HWdH7/P4FqMx2Ejtf3tUTJYXy155ZHT465FodAO
klHoG+4mxFBNDWHZ1jvTWZXNBp82E4UVsqTnyl3zzExmxJ/3hGWU6O3VDc5t
r0jo0fj9h1wu3g2bQGFKHIrX/WJ+d2wOVddnah1ynKdYmqe6WhMN7Y+gv/MD
KCxa/bOmEwoMn9r/uHdpAGTMKeLwyjQw/0p86v8uESd1q1U/pbboLZFYgGa1
PWT2EZjLtNqMdJU3T66pKv37vB4YBtja4DGtf+FdrcLnGUlE2qJVKCg/C2mC
VDb1EghRumVFHRyLALVNtU1a/zH790/GEmKKMKOrrLszVhzBTdVIFSUbm8ii
T3CApk3+R6iBaiO+2PGIlVCJxOR3Ij1JCML+FPkfirwrU6r3XumL/hA5dGjG
le1dkbTtCtMF7VfT5DicbdpBcSHsq8GrPl7yVllZsjtiCpaoav0V1zPuesDT
aLr8zMHLpbfFQHhLpUK/4mbbVfY1LnOqk8tJ1DBd/QqQ4GH4Z/wKLtxrRpFa
ncEQdoDTp4KjrcQNw9kGEfGEIkfclslq6GZrFikH//qx4cBFWKpMhr3KjEn9
BitRhG113xnp/JJ9PxeWxLLn/zvpZZvKMxqtrgu5Yy58HmRkSWiJV3TbSak2
nPxxF6szvr7Z2nJ17lw69dV5GQn+Mk3Jz46RpmcbJZ8Vg04yqsx1TX66zHlG
LM7Kl9NBLBvHDgrgvtD4G8DV12NcR5CJ/XFSOLnh+Q7gVokVitsczThpjDML
B1pno92HxukvSBmQCBLExTCBSBJBjhua4KDI6BE918QrSBbcVRxbDsspwbsI
DeZAdmDPn+HTetuFPwq1cXTl2GnWOWZVtSpEpXEX/crBqA1l/CGsw8LQlUkw
KUnBdDDL8ZAZ8PSyDSEWeg/sl1SupO/MGzfIt9cY3piOlINlZ7rZFvPYqh+R
C9YH25i/ksg/V2urYVwW53PoaJCh0gixN+lu6/uUOnRPEUeTP2IyEVxQDlkf
YJIS3PG5oZnx92MVuHjC3hatXsiethUNrM1Jt3jVC+k/ucklnz6aHmlj9sET
vxb+fE/laV55klAAzP243vWg4kIUMNSb6fbxDkV/U1fCAiST7/pT0FXasfRm
pFO2EK5tFsJ94/MYtKY+oyaDo4+0MAKPuhL113tNmXDZfXd8u9lnJ/VyN3xj
IYf4zdFBEsG3sMySwyt7Uu70RgXFxj+jaA2KLqaCSr0BfTKuPlIZmTugoDdj
NlGmSfx1fQ19fyE20Z59JfR+yEtE3oC7RS8RjIL6n62XtudZ35b+Bta3gFaz
5D25Sf3PdNK+G4JthuU8w4OXV407pHWGBPsz9dSasPa1Eh4pD2JoJMMvewwT
e+nUWMdisAbAwFmbc0PO6BlLt7ezoLQyost6LJrOyXLAPG17ybcdcCLCeaX7
oKqJ/mL84wo99TN1mfeN/FdNDCQ0SH0B5SA9BNnXyZKSAzPWkNO1JbBRpBZJ
65iT77BMZZGnFenjlplzmkNewnw4Fdh2DFpuXOkQW9YluRMwZh6Cp3Wi9X8/
FBN0eihxZGWzlidpLmLxPN25FT/qNATvixlcPm0ATE0MO7ybxy7PoxbWu9um
nXI28PjjsuQ4/ENM2lAsghKQuKXi9CJNjDvI/lJvoTVBRFNPv3eS+h8bFQek
UE6rUVGXGhDNBbAfe56kzIS1XxhXJLpGwiZq2S0FcAL7lDfWTZtIZ74Je6kt
bYtXfBenYkq4Uzc5xWq2+rsvZrorXUHtoUG4Ny/J1Zlxt6VcNadhc6eyf8XT
WvsO3ZGA8tenbsLlfRe8N7o6UvW4I5TbZ+YpbpDkFP9HXP9VrqwgKGLjxpMC
mx0oRIRCYe+BAp5hd3kYWccB8zfQ6Wr2J+deJP+65uxRWkSIoc/fvYmqd1+N
GTM8ADI4LDbXWuIfhIe39hy3SymUSmJ89ljraZGolaWNlm9oUZw732kKoINm
N2qu0XoIm5kTF1M7uCPeKfl5OwVkePPATNDBJI/6UFKDhf0PsbDgstz0Khgh
8/LhzSGQ+RzBPwIk7nT6IazU2W0dHPfDcWgVQXa2cFjzFW/d67v0OFfjawBI
m2LVcNGKuoD8pH2E6FDm2GKbekwE2pof1HRCYGmrQixJO2WDNCmQhf3wVR4f
m627KJyWx8oE64RNID5IQ5Nhjp3fshbfXQIv9V1dqm6ppVEh62pa8FTQr3fi
WZesu0n/GzJzBGSmYWT1lpfTIInt4cglrXlkHcIiYfsLrdfXWmkQfOHte3q5
5M96OQDdq9UGDOsVfPral3z99NzOGucKp08wEy1AASkYJ93AMUh19x6tYqPA
JKXk4EZOgmLmCjXfiqMjmUS2cACz4mbuyQnP7qDML7Et8eqSwwxV0yylL0D+
Iuxiur0C7KgC/3e84yUGbVvjTfwVOB9fjBnQQVZpKPfdMIHOSyu+Q7uh2PMc
UCGDHNQiQEQ663YvxFspUgo6kdAIxrl72k3jZkdLZzOHJ0o45rnFpkOQ66KN
b29OFg6FQ0bTMTveBBtPddfA3CXQXtz/i3rSPAqgIrmsa4LqsfOSU75rl+YI
1Vth73vVxyZLzTolmw7bRK8GWfrVAIVjJoN8M1EQQdbDY4fkGMjdwDohRXlr
XYPmYMAtfIh6OiTMLB9f6kpR4E/xind6hshSNFq10TXGemk1mzGDxOayJVhW
I97tMmGrx/1ChGZgvaJo8b/TfByqo4ze0DpRaSqY/azw98KClKSmdybx2Zo5
0pwQv4UlXhdIXgE/MyhxpZVPNeb8WEN0AOHESXmdELUgK6yzdJhpDQW5WPMt
W1tVDdV35BU32hFzYdQF+6/S4Y0ZP1pH+tUMMwYzoTpi6nlvPI1MU4zHEbsF
UFUCIUz8+7hu/nC8bkhLfuFBHr7DwfD4j4mwZFUKGSdOuN5t27JV8mW9ES5W
V4Lh3/HiGmNA15fnqKg8++DGXpB7FKnh0bwp+jIQezVzeC7r4ieIAUDY8Jut
JBNIe8ea374h+KmZIJdHcVuHDg8QTU5qR7sOwydpbDg+Klj/PyPD2MsNzOnb
PGFbpYpxClqqeQabyMFr4w6ClvzbeV7NELtm3NCIexnqUkJbsdySVYIKCkZw
uJF//vbj3GKyTcgLvBmfvm9BWmA2onFG8jeIJgR8pR1lAF+r/9JtZu3JQiSC
JFPL4Pz6bQ5x+/o+uDqWlMBDOUekZByx5nEaB/+ArgbhgitmKBKWZxisJjhW
mB188Jj3YwzsrWNM0l+2JXUkI4PsNtDff6YfvYyZn7Id1Hi26Yr627Arqrp3
tB3C+h70dLb0sm6z6YXNqLGIMo8VYq9lKMtzZNGvI6CXy9XWH2tGVmQkGy6l
sJlKzN+86+BAhPeDrTRqSeiOfTXl9hQ16zxGU+W6W03TINJVHTucjn4c10EV
NgEpYe5UPkg7/R9UAA376PQ4ghUMSZinQDxTFjthvoESvqeJoedghvnUupHY
4xUVvGPTY3GTYNsavxEiHdFZWSGNtfq7y13cF48s0ByFzj9ZBGlioOVxP/yW
M+flV1Aqgybarpwbnugjg3liOrkRI5D4twAYq0gl7p/rKs8STsutWJmZY7do
5qZzh+WbD5FtzmOCdrvy4QweLHS+ips7IMZXAOHJ/q3WbYIO9m58QbVEtQbK
Hg/juiKlKPYHsR+SAa73m2TNATvftBqYJrXLyIZtjoj0mM6vWERIeRoOZD5J
kydQNtsy+wWvHXDTgnTUMiD4CemOgewRW6ab3jN10AVM6IlKtQWPDqjvacEN
sF/ch+HElVIo71S7zenOkGKSwu+TY4kNdmH7IMDIpUqyJmU7kPYHmyuoOgvW
JWOXfMvXqIewodnwEEYy22xvjqf/U5damm/4jGNqXtfh/nzliuYDeWm2GgkO
rmkl1Zun2s36CtoIyu6jVsJukPuR/8yz8NO9cU9OI6JIy6n4fy+wq2LLxt/5
6mkhhBHvafJoIouNNL7qP8qn2iVatDvCS44qDB7xqY3nv9xEy+LYCHD47fXm
Jtr6HQOtsEBcnKlPofmmI5C1MHg2qTWlCdru2+OWW+n2JW1xBg2SF09rGdf1
c46ZQHSQ65wtL3ICcyg7z9HjJmsLSYFFq1KDA+TWbmyrqp+eqSs0WYROBu3p
9Ix+jjwh4kmvptMkOuDkhVAP+gph4/uP+SBRR7qtYyH88mO0QrRXEVGlOKSA
foN9WS8pjIjB+/4gv8V18tpDSLMp/ArK4juedAhjjLMUNboeanAFpM8Ti2uW
AIadLVRICZ7HpTOnDQ3w71mtyT8B7pZXZSyWJHlDR2colRR0YZATtgZjoQ3U
cmMOqMM6lRu82nS88wFvY5OBZ+sLcM2NXYo5wTD8KuYrQNxcPFpbuB6hc6+5
I/IWSDRGH7uZ+v3A/2dwYEp9a75VWSaZ6GEeiiA+YA9TO7ZYvTMBDXHcuh46
WJHoRjlk4GKlSRudsZFNXAmEcSZa1NtWbM9xeDP8Y5Ii5Rf4Czbr9KGBokx6
iGBQLEtjWxA1j5fyMzOA3TwqJzKCYLbYNmoGm7mjPoeVfWEV4SocN5OzdPST
b8mGQ7O6mRtXpexCF/W3vXdUy+cp6qr9OmfD+2W9oq0kjiMskhhVh36vxWbF
3JZTjsMzPN3oLBkH97PQImC9LMo9Wt4PUKN+nAMB483Ecjnrm5qkNs6Gog6d
FYi/sd7D5X6wFH6QX8tvQ1z9jyHwh2gpJz6Sia9QmL+rWkfYw5EEWTt8ogSC
FkRjBcNEzg2/O87fbAjGURWVmZX9PDo+0sFKvNMXTAXxrpyB94lqw/EGINNs
5G6JlUQzKWhDn5rf+94g/eV/gfaHfDYYKVtVicYFmy51m9yRa8Ks/kPfDPNJ
ACec1t50r4AZQtuQIEqjn9XB0CHhtjtN4ds2Gk+shNefyI0o9VfLjwpcBYy+
/3ePqTnl7jalW2T+xPcZZbXw/x9jyFIdsY5IWUlzwkYTvoKEKg3BScRGsO0b
mteRXHHFP14FCdG2oVnJTbM+SHLacuWzqmyJSauR0y9z47y6dQxQqMmueVIn
6psz3hIUHppZZ69NKWEXfIt1izH88/KDVnba824eyWoPcSX7p8GhzvtdPBqB
uYaSTYKhJUyX0OopuThlqyKEVt+oF1VJWOFvF9bHabX/hBeXFNnETcLtmxBM
08fsgfdAaIDUpZg8G23xBxUxhecfqHyHe2KwpzOkmZZdiDljvHX8rP86htMx
V4xpFgxQCEMDjCt9vRkHYbWtRo/gMaystfjoKxJlMSYX0qpnfFKNZzTqU6NB
VOarLprf8kGlYYWiiIZvdT3DK1QDOgm8zczvAGbAEy/1hkd0K0tsmHXXEOIU
ODbEdOUv59c450gUjd54teGkxCPWLxzGgGTCPZ0Cj51UP10DgjzNlo5vQxHI
5/4SGrSbL2le6HJb5YGED5g9BrJnnwYK1X5Jxx/4+vOyOAo7xwWRdCp6F4ON
odq5qwzx11Vg2/sgTB4MmXowghuDGQEyhe1Zy75PZ659gY2FFDzOYekMwL5X
LAFC9unOr/nncOYLKhPIXQ4l6Zc/Q9wFyNWvih9+AAhHJhjCSSpWerBDTiHD
08f8Vly3eJyhqJnWA0nVUoLS2Oa02luUBuZTLuRUqrreULdbjjq+dvrdhnXH
G2mCB4OqRhBoL1vYJ11i6UGAASqu/T4+QRWwGoqRLKrKS7bVtK9udRAPkaNq
xGbnEr2lDxOIpgDEWsz92UgCwrWs1Q9AflxXmzKLuLYMMICwnfoeHCDHEl9Q
JZpHvwryKNYEAPm0VON3Oxc1i5wNUzR/0IgEwFt2SBGUTquntHBon8WUGGLz
vfrD7K90AhUEGwx+sdUlpZp62CBH8HrfPOrDPnQl/5XD3azRSxJCNW1ik/3M
imEhpy12XPOIxZbsqH2pi3fL85Q2UTCXJS2RfV4uOFteB4orcMGqqqQVO4QA
RbuNUi7HWT516S0mQWBxAmm1IRvRJu2/chPEN6K7luQmdji1Xq2/wBBmZ6Mm
nyR7Hp2y/V2N3U26Czl8re/pwNghi4yXlK1FgaAsyoV0hoJeANHoriUrg7JM
FpKCJCkMUXMez60aA0KLTnW+wNRD2ZOCHv3sx/fV5n2Thnjp5aNTJpcatj4y
XNBYuoTKUsPmh3Ztt1GEXWbDhQFZ/K698hsgjQd2wNuqSs/YgdpEC1SzqM5J
H3XOttBx1dMxI/Cw9e5U0w8fQAtQ6TtYp+yd4lxYuOPaEsguerrsyLLRFxss
zei9Txg4LKQbb8bjGKDiMQNKPXuEEqaSUL6FolKCKMI4VAdSCNY/9zWi1vsg
QC7YmpHGEL8R6/n5a5Fg6zSPM2ultdZme7R+zpskcfcu7YIw+fkTJ4nQdeXS
i8XDQQsKQ0zPDSdpV5Mo7AKoK1VnNNdfA1H8j6zr0aBJlY7CM9hE4rMqx8Tt
8FRwCfcHl2t+u+q6leCZaPe4nQNpkGAtJY1k4mBDaCqqrnxd+QAwNVnLH0yD
7+Y79wd3C2Ni6RUWoQBooMFL6QLWOyhNvne/Ca9TaF6+djAEW6L1LcexRUOf
OBxu3lhijdjuK1Hbt1veFYZh55zTXBOt/34u2qtHny3DOxpIqG9pcMo04pXT
QByvhotRJWxB6YRO/2jwgrbkaPPULTM+gkVs3OTmnUepOjW69HbHc/n7dZeV
ILCKwqHza5cNc/9G6Wpn9CzfS2S6vY2EZp3Z0OCidIo0FxD62zi2wbYvR2P+
ekV3BY/Aee+yNLHY/Q4unPzDNGVLg+vjEtc1TEBzKrZeml8UP5BthCUNgOc3
j459HUhexTY2uzDu5RBdcInR8n3ogqsd62ShWjfH0NmIXEEAXZMYgXHT6ot3
MsOt9dKc2o/nySGCpEHDJxocHljGC+9UBGK9btRvZoD8nybR9Dl9j+ldfwbw
F50hcIetPMPSuW1ynqJhqPbTNxTHZABuR3gXXA6YcgAXfpvSsnTQclM9oLhj
nQxFLtfrheBmJmCrXV+caMgTkhHtoY2I8vptb3iWgJg8ry6HZmvlobiuHIxJ
pJB1rdf8YrTCpxBLz/EtM4P5ROrSrtUFvVhPckexbKTqbJ1np5T7bXQ/i5wM
Pqkgkm0pFyPFlmZboyai4lF4yv5AW5z+1Uq818LHccvw1whc6wpOSkGxFdIO
HtMknMREUB4mA8Xj25hgCzKfBE9O8wobrCXU70DnsF+j5rC5UgU9WR5mJ+Z+
wIovuQ3HqB9i/iOlpetnt/zhRij1ol8yy1D/xTCGF7lWamgB7mUPHseEhk2t
fDx5B8lXoVv5Lqsomvtz54Wt/ZKUtDZPaEba1YrVipX9aozQX6QT7NeZqaCT
iF3z6qMaVStf5XeXkLfAmId42kbffNLg5mAcWPk2egxDoWk4BvVjQ5yzCv+8
bOaLsVWKa39qQTHRPeoi6z+5tIuEjMHjz0dgiMWfNw1cfqxzlBZPui2S2ly3
dUlAIlemUPpURi87iLblpu+2Ng8vu3+fNVjeqC9CeREOnf0JgJUoyKmgqekq
cUwfx+qwnyhsm/xBbj0v2WgP/Ot8YCBBmJ9238LfyIM3eiCvRcgGYC+UCYvu
lZbig8+0tM6eIK7hol5KSvHEGhKglom2s/9yPM9JRaHOWwbscilbNncr2Tgc
iZ1/+3t13oHyYuMXwO5gIeqDWPoRKOTRzdohIVY17+WC/hYD8Db0NLpXUAar
6yZqM30yT6NlWhnSVcxPAAZtB7zb/Ev/gSAyDIxpFyYYS+6e0OmKJkhJceYe
uC3LmvtdQ0x5Bj0q5jWFfHTl3mvzbS4vXtDv1DP2KWisuiqqNfN0d1wivFGc
spUHGII+XH+L5mkcojeI96eW1MvLF8HTuI1/Tn3aP2U/ohhyhnHpz+TBAbo8
fvVUNqoHxXV7sxhPd3E7TkQdKAZ8NdzFYKiYGv31mTH87dbFtOBd4doxrPYg
zcD2tFJX89tBOIlQkrELpL5Gm7+DoxDKmckAg18DLUu5Rqy9INB/Gv3pk63H
PyPddkIxLWbrr4rDaqZdTVDSrT8R/AtoJhAles6kRynJp4D9sj43qEpfqiKK
tmU8zI+Jz7Zc3cUTlLRDZVxP1iisOcqqbqP+6htPxdSyp37JtVy749S7YrJj
PxCaln1RyhzocteE2Mb+ueACbQFtgiX19bfyckYeUHeC8T7YWLqxGeXWy2hp
LD2m28yTIif+Rsbb0+HZuOW/oE4o27LJODMuXDg+jEUSz2+itxfMJRYbnTDU
m9e/sUcEncNh7yDo60dMXII40TQqUe4FSlrRCR6owseMkJ6DEfIa0Y9cA+71
hdK+7g0mNA6utHh/cZpJTU1RBW4f+siuR6446baU4+WaUz+9ONnPidT0uwdJ
wIrU7OJtPr4Xk2eIZmFLGUMqmgLzW10POQPWx+9r/D/s1KonscJ+6+81plnr
cI2uJOIRq4jsiuGNtl/59Zn1WlPND4qoDHm1nXOpPgXbTohXDjyItcelxOsX
V+coDp25V5BFJh2Nuz506h6V0Fk6eN8stpxsbZZcnLSYmoN8SrTvVSfclnAP
rSDXkETVPwITT46xdCmzYTArUwF8uKhAFAdScTY772rZAC7ZG/ra/zv8iUOO
Tw2PvIWyMByVKFgCaOhif3ueOus5NdbR6Mz4jFB9omjHBQEeqQZJLB0IdeA3
0mTx3k6at2oda1jAU0cKnG/TuS2YjHAWatoyFdrGKJBAk0MoEzdvN72WJ+EJ
m+e/8q61aKCJUwpNBCFfR2JaWoVC6HyzPPJw8MxG65aqnMUSlymwnrmQA9Pk
A1tAdzo9vcs7sPhPLbnWc5wPzuRQEOqq9K3PTJJTsg+3/eCOrGT9qwE3j5LT
CXjHgBhPVdlBoYo60zz5vkmXyVB/hOCQ79qwrKfX6fI6AfUnj1tI13ESnkd6
/Jqw2nbbMQRLm0v3VPBLnfoFx5MRl4l5duSOyXfntR2q9j0X1UURcJCmaTUe
kohWH5E68qY2mDNTBg8BGehxfU3hoiKbeeM8JujWdIDWfdVUtcc5nPvT8NWl
MS9pUGjm+yPyrPIhLbwD2PKLP840Lb2jt3S3eBCMwNPP4030Z2hK6QuoPBqG
oH/Z0bPEaCWWC5+xoIwDVCjfZRgurcp5uUqKyrUaMyOkoqtkgI+1ltQYSuK6
hfVMIegB9bDxFQBnxNQbehH9Fj7pV5S7X2U04wk7HRWOWpJ3ARkj7LQCgRuO
Io5vBvQyuQmXb446DUtwoE0Kgft477t7rlm9mk91j1qIAF+V+xuMPOBNNU0Z
sz1C3U8wXo/QqF7LMFmhNJn0bogHQbtWe2x/dntJb8kEnoLHJVdurJGSnycu
ydPQtDXKCzh96hc9HFibvy1W6SqIhamrLZZDf29UH0LlAsxygGteTGCGzdcF
jJiQWQ7O4YDcob0g8r0KcXN3cdIVO0X5IoRXqGoeH8WrfGXX6wNz/6C1Q1EJ
S6HIdykx1EAHNW3Ua/WB0XqQvNSQnQlEG1HHavfjFfdIO0ypnf+cPBso6K2s
UkiIdi9wGF/c9OVqajB92mJkIsYlMXXJwRNdNxeDnbidZhkOGx7qshEIwZ/S
BcN/hHKrPJO42MKADJ6005nYPaklOieChFNLfK1cmN62Fa3njVqMh5YSYxI6
i48p2Wk7E04TO6P5IIRDxzM4PrZhkPlgKtos803pq6NuQYdtvZj5rDnkIb55
Opa5drckD5B2IRJw/ydJEIOGZzuPiO+8N8u0GHEXnqUDzQ88R+iVQ4/Q3vUk
9kAThufsWXyFmqSEya4nE1QDIWnbYxYlvL1lWg8e1djvmnr15NInbtf2TjRn
/6+4BRTnymoSo1Mt4fpUsZXXtl2x+UlaaRiJ4sSTipMUQqgKJpavrJvxsX/O
WVVUsGXUKUFLEgin5o7MurOgAxV5n+hBOG/02zrWM3dLcISGixisLAfN3SgR
JtYbEOZcQkm4arZfQBh8ZPL3NOtN/Cx5EIH3Y8k+PZL6ygAvN8RGehx9ao8J
jZkhMkZPkP4dd/7hmZychZZ2jzcW7Hkt6nZvSnDCazJd0GFppCQoIufpfI4w
4EppbBXD/wrHAO4gY7gNQp4diUDizm80sat/Opsvd3XVHOMAhgH6Cof91dUS
xcVraZy+MHH83Vep8F7/+RhnzObXPSq9CZJpW8QUIXEf5xiUf5hv+9+zujY0
DKjgiZ/lBFgbGr65/820wU5lM1HbqQKgR06TMYjsscLHjeVzzUy4pNVAszQK
klLik4nkc+TpTMEXsP2ziQDW3rq0GJVnyUltRVy2x0FRKMEtIQKpbit4Fdj6
j794+8/gc6CGZkf79HNDo6AkCHloUYKUFDfilxAHNrycjR3BxEKYJFsqI+VX
+X9YwVPIyB+7Z4LEvaGNYISentF+lqmPIn29ZakEe6X7E5aLOrt0hR/gtdNo
9S/GJcbUMl+ha5xGNj8vaOsCMioNLhsLYsvvdrXQVCA+eWe06YLkGy6JXz/b
AoeY2+V47hI0+I/ZX2oWo4/PxGR1ZXIrawtfmth0mYYPp3IEWr7IBNBODfDX
9BoptLXsSH0NTj1MN670oxH/c/VIbWGtCsJYVucYaLSmUoCyMXQXIrLfVFny
i0KrkjRm+hC+F5FrhvG2odwQUASilKmqeXjef0xAQutWMisXZD/Q7qKn6l+N
Cy4tSTeW+ukfjeAZSohZhGF7rBezAC6JJbvmPyGQjVUT7KC+8M6fT2MIBKxS
svQ2IKohCERj0CwHXP7vPOu0uuJmGAl9u9nn4Z6rsKdvqQmTtlE+NnZ0aRn2
ozGoSDaUmQ95R88R+W/F+/Uy5zcUSMLxwu7XQlakb34m0bqX9f8oBKinxkS7
YjzMnDJouOl4IYjbby/Jtkyd1AXaDXpGsa7XmXrM6d2CndKAmTplepBMTZsy
O6DhQll9Nbtfo2YqIiu0wyNovojEpBtU9a0TE48gFI5KKFbllYw4T3D3hDMJ
HqjRHzlylZN/MNAwNejTJrQFz5bIctcl/FEvn34sHymMce7YR4Micxi31RsP
C2No7wH1LBKUCq1ZI3dDxhRARvjY1G5D704pE8dTjgbQlEaVj8tZofB/Kdp9
IAXTdjQ+JVPxXUiPRW/vwgxOc5k9j4pfh2KO8SY0iM9vM6PbArZtA5vkCumN
ypRkb19aCTmVpcA46SUGkpraX4R0tcfX7uSPkCJJ3QEDTYNg/rltLAN4fGXW
MDH0FtbKm3DenTEDvQKEDHgOcr8e0o6lFacxtBsSpn4nfpV2+2eM4T1ZNzFN
RFavmh/6NLXDzkNyNl1pk5RfufqPumPhkB8+cl2KWCY+FSkt9Kwd9+r1FeZO
9Teic8kDYyIEwJIiG1yH2MwSE5l51I4rlvsv8rP33wRx1XWTXX93APzWdeHZ
0wYuwPdrpk1gmLf7dh8wjTPuQJrdQ8mso28L743xyiOr/pSxUqd6y4f+iWDx
t61FogVuxdNOhZfWD2nYR4nsX9tl/uMLJLQ+O1mxHsdaup4+8biXzEEGRbak
gbhREwpCd9+eEriBhWiyCE8hkyjRvdHP3JeFgca9rEWIdhqO3UkQNQ8e7Oai
8J0L05hSFhU6X3BG9zRJdncnIyXkpCBh4+3bdSnX42Vi5THzvdkw40RQ3hIS
IF+Vj71I/QsOoLZEtIy8/Yx3MKylpUOyNXdAv0dQ9BJqusRT6kEtSSDxB7D5
UYfmfrYXPIy9LHz5NdihrAHbM5vYYfIFQ3h6/zIjPViG5+swoSpD7Y00KUzO
AQnSn76ihSMJwEnbPF7OO6vX1riUhMwYhuYCsRB8ozhDWG3IgfqLPoLgVCL2
hyw8xTgTgUsxB4mUT4mYl2cyu5biAUAJ+F2tYWOj8MKc4ySFmw4rMMcfX0Fq
3feefRTy15sJvZ/UXBob/dvFBDCThriP5nUKVmixwo3ZO4KvNzAoYVd/4Vcr
w24ICWHj4M3wv3b9HK+utIKaXFFJa8Sg8p/BifxRLa7ZmDH0Cc404W+4bzp0
uRjLlCRa9zIlh9CsZTKCaaKirx06lzLRzfHNV0oZpr55RqEkzuo1TbM3LqF2
ZfBV9ZTAHqrG6vrJdNGaiue/7T0/r8edAAsZgNhW5CIdWOB+RNxSk9R33zoc
uWJZcCTIUQaR/Nz+GdkRbJuCPjnlIuZqf7IWZlLsVVCFuedLyS3heGAa8Kmx
qX/MPwD2r4nN/j1woVYUnH2v6HHW8fv4LieAqsHR0aaLn7KJQewZwnXsSClk
zS77QMLmeNTeJ8p3lD+AuCkllw+g0Llr1q9632fzLSlQ/M5Y+fRaitqXcY3L
KO+JwuhyZhMOlyG8kS8ECTo2/4x49rqcSM0E/Mw2ucZxjLaMV9lrWAmiEott
dVmRnwfOVE0uYJ+IVc8B7gJ/auBLonWi0O2ZPqoys8QTz/C5h96y/bFWFYeI
lX36fe2uvKNhYnkyFk4764UJidivkyqLYHQaBujjJ1ufXH2jXfAApfhAEAgw
NWEuJ1Pfbgx2rxGRxxTimUcL4kn13coGlsW2MeYRJz4sCo+G56rFmGaV/mQV
VecZILi7FxaU8jHT/viYOZLksCxC6W6DTIhbPPuOcmkdHuXWhi/0ws+Gw99M
S8h4lO7vP1Czhn59zpPLf3xtWVTx4RDleYPJr94Kc+qOOABq/tZiN3ip3Pjx
NtYkJSNyDoLWdm6kzQWbuf9KXoOxd752zYcoJmFWHk83Bpuw1hLrHlmioVji
Ek1StyqHTH6MJ4U3MWi7khLYVo2vUkba0t3rZpnPcu5rVZNO8WcKxOeB7ZdU
7UJGsoe10noO5f+zfWU7uga+UFPmE9UzP7LsQ1ygT+SYBnuTZ4guTGDbqmaD
+KTQsKUpxPjtHQXvtjrJBTkmLR2EwBkI1Xjiriygz9xWGMafObhKz2CEDxsA
o8FeNbMpP3aj/DUsiULZ0s6QncboRsMWNvD70fqwfHIvY2UpiTtBlkVB4ZYo
n8gmuj8UZlu+nNmdjWywCmVgPafc1NRheC8lb5XYcTGfx5OOOgs0GVcTW//C
pbLZX1yjGV0imWvh1OlLHnS7s7bWc7HSfduRx6AX81x2tK4rQqjuTyTtOfrz
LT0COlo98gjeibPK4GttBqwhLc1d9hYc0lgT++eN16rkOyvF44eBMW/Bbnw7
JAzltJgojD2QmJzIEuA0NNIfzWOua9gAHP2HrO/54UEd6gEqyiIJnfHeqW3U
iF+6ax9NylyCp1gNRW2AtjqRkbvuzG0yH5KRZ253/o+Sae+UQq7K+QY8fHJL
M2Ry8rl73PEpi69jELY47uLJlyUcxcLdCufzkECLK/7pCTUTsYZA+KKcCGvK
+3iB04DcK42sym9QALCg1OMnmsVRbud7OnNc3ZgA9qjI9ICCqdzsA4oxBBkN
M3bEOgssQOGvVMugjtablClnDANtRb6Kx+C8wqOFD3x7RVZknHU8APqsQpTk
OnJOjDUhGxkPlUzK0DbZt38ZmxVz/QMAph44Cz+zUR5gM36lguF1YyD9eFrK
NBjw2QDWow3A6yfuXZ3xzcZLp7NgWpNH39dW/3mg8c4B1JSdDC2YSfTOi8bZ
GqNETH/lRBEKT3yHPyhc9EnQup6pEUFzWzLvfhUvL2Vsv3dOQy1YaNWBRHd0
Hg8mML0RqL/d02KvbrSSdtjOLhwJ4FWz+B07q/K5sFzVlECPxqLwrKVAM9Ep
aMVLJd2Je9G7k9Yl19QqbpriEBZgmJM70APaPpzNRENlivlhKorH3FHeLmkI
7DU/i7hkaNaMTJdvP80J8nTUXGl/39Lr8Jl/Bs2SS5L2z+DYPCJ/mlSC37IQ
29H32O9A3XG7i0rN7y04FFvxmbJNHW/d0TC9kGt1tNUXpFVKISq4O0xHQ8IK
Jkv2uWVeZZdYSPmnOQGDwr+J0ajlpBYQs8d4hnrk16k78TWsISPKfK3VzkFi
30gWfDy7DAq6xSs0crTvkxqf4gfPXufoHRqlcyx+yv49Pk1+UBcom+8moqpe
9+PcADxnORnmxN6YfZEKrHjCTZrbZPA1ujsWLnWlH9We0Ma2MGIMkP0Cey2I
b7ePGXLmrikWH8S6zF9C2rDSzIh0HC5Q0bRsv6UfQQV2IVCxRFYqcq6a54Ci
UMeN2G7pxOlQrJcQQKp3encFJ9FwlnjneXLONGwsZwipYkha+K7hPH2CMbHY
PG8gRHCIGUHLJJKmsJzbm5gGk0a58yQSEMrO71P/o2hqv6VRRXdkvMbeW0Kc
jcgoRpn1E5ED+9haPchqZQiG63Uac9pDPpwYkctqUvWECVWJv4wppYFt5W2g
BFbitQjmaASLFO1TSmVVJG18h8P9zNsc4DF59yqibPCp64/aFPeTcQH5jbRe
2RGKqibt9PLY+4+ryjBbPZtPUc5QlcE0fm3m4T0uUtXs0d/LPnGLydHvu19z
iNuiTCeU/z4WgahML8aTOLT5jrnMJy50da0KyWfm84IthBLwtMxEUZ9gyHAe
iDIba+ahqR0EIrIWlGRTtjsiR1ifLibv1oKrLv1wGtzG7LO8yAgSDKIlYQdA
AXoO8cJoTmAR8uWsfMd2jnddyHhjc67eDE/HJFXk7b+lAhk68dheCpccz0dw
7rQAkPNqNSZYBm9ynAQRAbbDBeoACvAdNv7VauNA2YwGuqJNsv1aKNw7Xx2d
hMb8LlPTDf+MO8HRKoEoArhUhexeSIWrUDwZh7HVmm+4RY/cK3K4WnSFbB/u
p9mzCJOF7EOz6Pce+DylW4v7D6/8mWm2wzWK9VOVjOWirQPWo90SkSmjC62f
TeRUe1fgYe3SRx5hnvTHxqyJUL1Iizc3FPDDeJEy6bqSh4mt2I76wRZFmce+
yQiZOGt2Yf+e7f6B/EAQC5cPWvzRJtJUhYXjL9YNog3H7fYhacLAdMJL3/q7
8EjpbH30EH+aufaO+IwouNiB0JhgqvAUxp2HQ42JnKfMxMoUT8VI8Ak+UcCy
YK0UfBxZnHVx1i8Hkl4mhFrXt/Kq07cXFSu6eRxpOCJ7jStS/CgZOhPSBkWG
Nc6njinAgTr2byR5I+Zagi22CDfci5j2Ps2g167Nl9c4SoMpNdVe0KIx7Nez
Jy0PYZnmBQdHOvw2pl3S7HTRwgMMMA3B6Pg8QAJmeiY2WjiBygs/IAm/+9d3
HPMhxVM6UGQO39pQZpdm3hnuB/cfdVFDF7qk5oSgw4XDgiHF/JHn0Y8hn70O
AjvIgv1amygpE2DgncsPyyQScKwjr8GBnJIntElylmqmGnExyLgaWV+lGCbt
1Sb5viH/fpmG2Vcif8P82wbyFicMKsQFNHLUgHyHmlVzXM6YcuCsrojAeN+U
K9owtYSLRqcNWb4SybVphi0E4ylaJZguRZLwmGxxEK8Bdt8GQb1eiGYPxFEq
6adaRlSzcjOC7i/FHB4PY3XDy+DCVmagy8g3wpFzFJ1k1h+g3BMfLMYuUxwY
V4y2MwjDJdD6DW1Pbj4fgSd38f4tY1nhA21erh5YZPgtKT9qqKI4wGWvKi2w
oJagzVZMgohduYmQtH37YWkrRedT/uqywFlAI5E7Veq26fobmYsh95F3Jv4/
v4tsIRLlBwby+YJRtt4aIpEjF49JXbhgQ97da7//C516DawdVDBKWDSU0mH3
Npmn+Gu8PsQwbBlzESasuROk23ogh6UlRVVPNKQvPFZ/tXwXWmwRWE/dyril
Lx6UxNNwbYalVdgKjOsRkIlrGvCESrEF62GIpaKZrmI2LI/vNjquAJ5SLE8U
RdAAmYJvuaKwXdvLIVMK/tb7eqherVmCKP7SsLFPmOjMb9t4JbV5QRiqnL7A
odyFBsvvFPGReiny37LxHXwd8JXFdZjVw+2O7p4z2Ccag2YHLDbUEWNfExV7
Phizwiy1Ukdu31otZnTaNB8Vku/n8ELHFnK+JJTI2rvv19uZNlSdztuAQsrc
2iyP8wGim0Mp78L2iCP0Z6rw4fAD+Tiv+9ko4HYCKQ7MgdbUuRoVYpmuShOf
8dSNUodKB4Eo0K7x5EzCIG1xCOL9YRf/hph7w6Xz/lVgORMofo8qj2+69gqC
ogKoeCjt2mlhq1AnC2lSyb9f0xciQeSzJy9SQ/DA51crF7OkBZR3nfaVT2uO
gm6TwUr5aqohfCBNztLQCh8T+pcMTB+pHXUZvOc0icnqaCIqD8mcrz8A6ahv
Y1OksGI/6cVp0v30FSXm9fZphsC5A/2P8IiPARq7mKI1jMqddBFqgK1+FeBr
YDfSGqhlvkd8Ib+nwdPSbFEp81K4mErgdo4p39XWskfcbI2UD2EGAM2ezQWZ
c5uBuO1/VSCqocPBfQ6KL9os0paX5G34P8pOco8oaXOG1orITxbMnKPkBqop
FmfxaxLWqBkfzSXaEboPW7UNFFXuKEwNx4x3VHybWS1TluCcPMtnxzJfApF1
1vqdylsaIJceUp9oSlloPXJL8YfGm/yvHqK+7FHmvdKstVw6JnFXQdr9tC61
nfVPfKgqWlTHCjbrAo1lE/9LAUOUNKLDaMJzAfLthCJvWUlT4B20jKA/zQcV
gTIZFOP1/HHpa0TH0cO9z1TugicfBoalw83c1WhjOzQVGU/8StpOJcamfDZi
hKEwOoC8TDD9D7xgbcmbg7nf+ZhgVfkEGstlGsKxUXB08hk0JgjON7/ffQ2S
mZVtafGebC5sR7mEAawTrHX9FxTtO1D9SS8suxh6geyf/2HqJHyEu/BRWS4+
3gRO5KWSzGL55epk2I9OhjqwfPQoUPGpKIBEXpLsFA7FWef6pwcd/vMRmv2H
GlsUCnt7o6vQobBrMFNYKMMxDGCQxu0aTNfiavfyxoi8urCw6Jfjb/rYv0JZ
HpZqaRJ4DWLaewKZ9byT4DYMmNQ/5zJ81CXebBFhvzfOy5FmmEyZVsnRLIvL
1GPicdGqpEEF2OgZnYgktUrpnkWaAazR44E4kzl+i1iR+S9g1ALtBt9WiEMC
1aXRcLfa5wZJUKNcg4Kmtejw3mElv7xWvBIfrZKlM5adIXrTT7T3PLOxn9Dy
MJG5++objl2YfQPMqjAnHv2I12YEtpveIPQmWmEM/ZnxMbX8jzDG21qYUuEy
liNlFxr5IZUv2oY3p+TF+COeqgitO+XxFQKFDs9JV7WSqwrhvjIhAz9dz0K7
WcRUVER2WiAQrZAjgNfQy0+A9agdhKyTBMXaOJdL80XqSUmQAjJnKVr0N1E6
VEWhiwpwMbUO5uoQjUfLNEVKe8vtUgqJY7D8GuEGh1TBs+nzZwZ+uuJUVmnN
YMxijz6PZBtXGusEt1tj4zu6iAEhCHhUrQXQ739BPYPwRsxYhZS1kDNxRLt+
jA2bSzYqC7VUSZ18c49MIQnHvFbJdOQ/pTQ0dFruDaKnYCupBVXWUIgfdh1O
I5xsDG9CXKNSPCnCAI9emOggTQpD61hUvBczNRbfFwvbsYvtAzBv35ubpkoH
mOpMc16KtcuKsLqKs/lWllcAfZ/lY/TyOPEd8dGNbq9w5HOzqrUJMEPEpm3i
TWqzmyySkZffdfJztr6L8tlQF3sQM7I3yCWT9jVz+mnOqvdJYgkzwz4c6gKT
S2qd45PIlwcNt3o5HUwZLVdmWvXCgjlKPLJBlPR5qjhd6wOA0cTgrWWoejBl
lkvFeOFXvUl/eU0H/gn6jrjnQuim3RJjChH/2XYs2jkrnc3huZCd6EaVkeNZ
L3oA9BPF8YfO48EpSf5GQkh+bpXeqXYK914UOWwx2nUYNN1pDGyHpRDR9nG/
G5DawbrINrzyrVVWwu3GWhCK6ICGm2YSnh3xT6ZkZkdsXhIyi7uYy0aKUviB
3n+k3jC9/qAPlcjpEfmrRGuOSNVZmTL5JU/YMHk3w4dv8oae+xNbHI0MLT0D
FqEiX793K80xR0F4axLpBzndTFa1DyPB9Y23x2qsT9sEZKUxuEXOuT8WCBXH
vsdZJc3JOmnWdI3+Ff085nzM7u3udqgDJkJTMwDKAq9XyOB+Sv3ziclsQ8O6
KdmMO8y1obZj/noN2O2IcvZjmeDKsSrjcXRW8aAsjbg8+VcxCntwV4nCho4V
tmlxWx3EoYdiU3V18KECVX7pYCMdnv9QVazEkCVBJ4629VEc04CYfTfC6v8v
fdqoc0Du4wawrNYJ865VmJSd50DOJSb82exW/82zWdiFG3jVJE1pLBZXjDop
/s6OhlGFGq+aUPZWCc1leLTYPbrT1Dkjv3LtjAnodnh3NGpEZhgnrtzM5I1+
2T2OxLXfevzJRn0hKd0s16eWNrr0sVY789zIIi5i/U9iFoLC/YFbbdPN3aMw
+8dQ0GyStlODI2HHtgV9FUe0vLs2Ss5m6il0XbQLXBBxsykjL/zTSrTr4ByV
1gCCxehefoTA3FrQXBRQ8DAidiMsAX7xrVM8cnov15v8iekYu0uuM4cDalkI
Wrj2kkJEKqrHiSwry410YbcazuoFGsTMNcE5fiDkUAhbvnSB/FBGAP5Siee5
CbgiAoh8FMee03BHSJYKNv0v1/07zYyiZ/AdKvo3EWe7gfdMb6rLG/QGVC0/
3zhQXZAQf+68abS+qhGkswSj6bApPE5amrKaE62aJjMQeqnIElpxxL1fe0Bv
T8H5BYoJGXz+Z0whmmFY8KyYBo5K3aLf4Xk8BWUVk8S5eY4THtQEbR/rmXem
B/3iyt4JGmu3dzunm/IX6oQrXTd8eknLyYSI0S3QLEvoqPcfhmqc2WZqA+KJ
oRtu1JFZj0eOUeJXjb7Sp9yquotISHTcHBI45xMSspmetWVsVUeriZhbPYBD
98Z4tG7aInrtp/U7ez3lS8Azmmbh/kpY9QF5il1O6tqAvovUcxup2INlbxwP
RMkj/poIP8Ra6v7yyDDFUGpLNW1kgpNF7yYHs85oGVtmtrUlIuF6Q7ybybcn
v+4m+kT1IXf7iE1oRD2HQKrikeg0oH4LkhHZIOUKFVX6oQVUc87rCTlhBHiT
qWPTxWq25nChTHBg41Wqurb4XmQsE8Lj2DIDNh74eB8GEn6zDc5cZBnjiHdI
4WnKHfZ9yIfWAlQVqrxBz4xLn5rDD/ftuIgC6YgBC6K0QML17WXobe0QWjzS
XviVUXPE1nqkWfFpLsbF3uVttgR9PX7RiZol4pZNlkM3ynJR/Ww/GMfwsujc
QdOeQBbKegU82tFrT7LxSKhRAHEMTdg41dBMczHCkdM0FcpWUKSX3nGN94fu
fPGBvbMVaBaGOn8xibHHFWamUvV4n3zOPwJd3c7QU2byF9XInoAhZjhm7hdF
Y6O9pojOMiZorf2SEFdipvFO2+GAclogB0NMhydfOIFtl/EvXHMhRh/z7O/L
IKAdIjwFGJrcRbNTbxqix/l2xujq0bC3wxabl1kTG0rRwQ+TECXochNNV13z
r5ANz4GxqrilVZuzX04Rr+eOVbAnIn5930xPHSZe1up4m5bq2I0mi0NA9Ayp
Qj5ZhhjcijHb8BSAODeOlO2l5F0N1140IMkPDQflZmO/fNq3o3D+YJk1K1xn
0owrAZih5iyU6OWJzOdC+K25mbXdY9RqWfuipEBEcd46yZ9klNV7XGTr6W4R
hw7m2MTY/IZCtyFpNFbh+8cwpe6YwHadjof0+9I+cm+j1sL8b6XXtf4IedFn
ZNm1H/r/e35spf/H3pqwHW08nmHDbSwRzqOwWXUQfsWWvzjUoyQ58JtCwpmd
KI1hFntsIZO5NiIqc2dFLjIv6kFfnLmaUQKd/2KibVkKeb65LPZFJa9vYbj5
OmXLgz6JHSLJqDZ9zFvReqJ9fJVIVG4cmUEgIHGi48Nt4/y3kF9T6lA7GpNu
9t8Q9ekl7DnC+tViJWO2o/xMlPYuSlwnyZGKN336VMaj9wfIoQovdm3Srhu+
/jOsMxuVU84BTVr/DuxXcPA3GndM3rKP+hJ3JFdTEq1YDDuUO3UQN5pxXYcd
g9ESEmJY4q+XVn3QcBELDc4YrdF93b2amiFqI/IpkjQhJCfTxgg1DVHpJky6
LxG1AAzJNsrSENUhDgERIyssdhMx4aafXgRKqCUxjpJiKipn+krNKW0sDZZZ
L7gZbNLV+9jFGAsT632LHmpJyUvJYug0IUPTlupRT2JsZPtOamU+cUDoe1j7
3K4MllwNnBGjUfJT4rKdVG805KllLY7xiFxISLIMTP5GzHsRZzolduJbs/Ao
15ke6W938/cfZWCf245HXCuIgw5HTppE+jHIVig+aSSlLgY9wHtMI6/Xn/4z
CoahtkRsTHc4SluJtEDsAJ1C5iQx6/8f2LWraefL8V5oh9K7LGKkXEh9dFcN
v4Ql+xaXBmXpuOKAB3N0rsIjsMOCdG3TN/cBE7AjwD994l4NKRAcekAWXt4D
9pZ7Te5ZGWveZ2XiAIomNw8WSFxeKLzo81r5uprHGjIeBk2wHjEjBXHT39Tl
HaFdDHMBi6Y6qJgUugVIV5F7yx4PsGmhchdKyfKEQpB3ARJpHzfEzVk8goFj
nIZmyK/SWKCQ/LYSDSMPgVt1iwBGP5G9AYT2adlQGPzJZZF5XgG8oJlFEFFX
lYxoXt2MPQ8VtqLbtneHjiGySf7koLfhfyMRUVioGluAxbpSM2a20+xuvYGi
7/ew3UFm6S7MZeGGnW9U/TB2kZh7E3kADttOXCsQwXzHIOLBGUd87kQDB5Le
T0soylY1U5i5sdUroiQ4JgB/SjprnfyQoABL1knj5jkbn6ODeDBWLOsQ0af6
oHISrCkuZ2LtJ9Y1Cj3qMWtzczpY1/aCYZp7kNdJmyl0P9AAiwkvphJsi/hs
Lam8qvjIdzum/MZAL5ljT/CDDU4t7p95sVom23R8IYlNg9Ow3kr/938rXS1a
X/AHZmNcr4bdukQL3+Dm831c2fymYd/yDSTQw/pliO1J7UA4a/FptXgmbTRu
etYJap/KgkviKuwm4gwnLqjZEGzs9Pli+t2CNzKk4A8VsILMIE5yJurGMgod
NEDxJgnaciu0XsZjmkyOhbJkhuBhGnrFq59+ZPssSFrCVdkLH/6UvRY8QJbg
ftBL5F5R9w39CRRV8CFsTSZvRBg2hmybeH/LJlEYuyZunERhlytgB4dKAY1p
xTA+1DIj2FA5rZRWUySUTSAUXD8WIRoiTdgM6pjHQM/rQNd6LkJnuFhqsOgG
ix9mccjgSmqoqLy1HgDPfbUiy+3QguKzFXYkbMi8EVgNijocmJnCBlD8oLKv
9f5K3U34mT0JYEURkhCYol8+n+1NfzCixrffj7stJYQoidkfT9bWNoGMWZxW
tv2tkDbfif82M+EyfGy5XHrePpSy6CZLjduG0Gx9nfKFi2x4AizvLQ4nkWvg
pgSB8WgyMh/FXuMOIGmUBS1jHlS8n0mQyOdp3lxXgoj+EKshQD2lCTH/QSGS
lfrEe4CjjH4UGbK8D892/Z/OeCH+J4NyyFWSUwXvnor1G0HCadm4RB2nTxHs
fsmM1FUo202Q8Zbws60AihjvykcgKbMJyshRfy2AMCwQA/0NFVUS5qWqqhL9
5V0YNphGcEmP3azom8HsfngTDtUC1To/w7ewLHDJx9s/Pg3f03mjd7SOG6fp
dVX/jVjsztahq3me/erR9Uafkt22fmuWryHqA87/cMQkyZMCq4pMqMNtn4s4
FCwPUF9seGVEo8HgUuwKnRraxuTatmLMiLPm9819UJ9Xy4uEGKBOhPSppfR0
IDK99wwEuKkXPcUHiZ4kDOD3u7IU41+mMGI/cWFZmO00UD9b8mBDAy9VGOEI
4L/GHVBmXyPwqmbTUdRhFBg7i4ECMzF7uwcQexVrfY5VF2Zkx8WE8Xh4g1qT
wA0y233firYZZsVb3LbS5K9ESlG/iOEY1aujLo8p6NbNpGd+SotJsQbG/dUg
T4fHN4mpr0Tkv5sXuegN7cx9zxE/REv6ahMZHc3k4DvNmQTPDysb0rb08jz9
zKaw/IS+IFfRH5bQzu5Eqwhsa+TC0hson8KMxwtA7dPgTfFeAU7g9NI4czlp
tP6GRLPttaAir5j1p3dSCDOE8K4wyeuNb3lWkX2Yy365VPc8BJI5jgKiHf0K
FqIxEwZRgQUNVNHK/CsSHfmXO3tzqRd0VLqOjRGrAsIQ9J/kZRzfZ1usPxix
uhJ6xvHMggrRkbZxVBzpV2L9mHFNYU0p1Lre20AqEF3eGRaQCyyhQcVdFsxB
OM7ndd0hFQnwIm20fWJ4S7y3kKST4eImihmm0aDfROVYOEorVAfjdgFLQ82U
o+jEPuSrbfVnFWAkjgAfNoknUfHEx3SZ6BLjHp+H6Hud/SB58Wl/6cJwb8gi
Jx6kHvViBUCBCljqhXbknYlmZ9dXWCM33bh73Uq771msZmsUpDAa4TqKPFOV
G8fEdoQZE46qZd4gEKBP2FlQaFyZ70npX48EdbHIannmDTKHCjqs3kBqwmmx
EcZNLW6Np8Yr2x/EWq9C42fD42PSwJHXRGb7nhyjWgkz5W5kHFRBFhLa+9pL
iPyJ0jtnZm2nx/Jn9T18Z2YMgGeoZw+FoLjE/+aRFrbjBs1qzHuzM7JcwvIp
o0cfNxMnZGHcYTGvc62qCiuGrNxi4BRdXfN+Ct83eeKNavhWnvwLvRUNPAB4
svFVBaUHz9zZikt2YRPcjPgqPzRveJkq1gWkncmQh7fyhAROpM0z8Dve/CCz
aeaJr41Ha8gaiGwXorG8vdSly1fp9ZWEthXrXeuNHNyzP/x1nL43KhwqRY+L
hqH3MUf+AZrUnCdRZEccOY3x07mhMEl5TEBb685icLWZ6+aDXjgd3i4af02Z
i+zl0p0ezy/Tp+kwZ4X5faFOW1EL+seOgeiJT1o9RFCdRNpnRl4Q6FjEsFyp
Ox/2q9VQblk5RlUZN6nPXSnTAK7zmBwTH5x93G4LxI4D83thfiicWuDby1zg
oe6Q6N/L17Er+vkWxCGL2ekwkmr9pBl2q0mVudpH/vAxrZKkfKwAVt8c2j/P
vxbuONCH9asjRCtHB59zNZ2JfQYAj0H/NOXX5skGNKTKTY+Q/hpAzf6UwjF0
yWvqYw17FbWiCix6x8frZGqlhw0RH0Btg3GFmb7ofePmbw9oMzuafSv4xPEu
Um966VyLgP595+v3i1sxhwzCwhu+qytmRbJWIQpLwv25W+Xqb8/ft/N8GEfQ
19/rfb+qDVa5lYGVq3lrya/nhnDaNfymsO16Aa6AjnHIMQrJNIsDUzr62wz6
9i5tazii3Sfae2sAf9nUm8jzUkCaDlysCzOvRrHvc24Ol1KzzB42D5CW7nme
boMhxkRmnNctv4ab/NRYWfgwQnospqjyQhoLXpZ00st9/0iq/FRryA96ImOQ
2RAQkhcgbsogD57OmXGhmCQUVBnmeHs8w97RSJzHYdjF1TDTyuN68orLj8ib
aHODqraGUym3264I0ZLDbXn230RtcI8jlIi8lj4gITgcONfN9NMLFlnqBCL2
v96aQDSfOIl2LjLvzY/aJxx6DA8pj0COpo37A2mMpAkJspaROPwQxEBmzHeq
MoDQmzPoWPf7eYAubSVwEQ4LXkpZLvpdeJGRusERJ4jV9rrRGnRUPOLsl9Q6
rBEa0Tkb8l/gt6Om0Xf4cC2xXzuf+9OVJ/zkZkZU2VweCOU2te+KUA3YlR/C
E/xwg+hD2+jtfqrFcnHvfB6GYDn9A9NVcgiIjwYK22tfwJjI5jj1pvzbvRlp
EMJ0sM+K/J5pLlXppSVrPwAjgl0+ejr9sf0sl2ZTfa8UD804iAXIEnp0fd1p
HQhrF3SAy3YAnWKfrUBCCpWgoPhD5WqHN+gaxmVm1IXRYm1S6ART3cWbM+ij
U9Z1X9T5LiL8U+4mrddxWYlfkyivtjuseOoRhMXEoA/tK2SlIldmCBG85YT0
tZJPsvmVPaQTs9SzA6d9mVzoYY2SvQTeAQ/Yh2NIdYNjQDuCoeMD8gMsE1dj
oaKlStvLh7rDdBY6IgnMI2wy3knJ6a9/IdgXiFh4yTdhW5NdTGxTREK5nix4
s+oW3DKBdUiJQmw91ToeEGvoHdE2A6UxVh3I3F2CWjeQO9+fdmn94LBToATU
ueG85JHJlaelSuXvBp40gNFBJV5SMeeCtY+X0a/ZcrtTK2yzSBT2A3Es6WmO
MVg1702Xk5BYjW1j0jLGWLN/n543s4PyEft4DQPRAWEfl/Yk7Ett/dG40ylC
Krt3Tyheq9c2RRqiZPmDDUen8walEgthCZQ6I1R3174qbPeCMMSPCZBgxNke
QRHWXpuN0TgCQ3yX8N1wSTC4EYt4YosuOKCk322Yt5SrB+jXQKMgTIzZoT5p
ymaJEHCP7dv/Zd2QTJFtoidKx5l823vvc0B1xS4oylKirwlHOfy1dhW6bOTz
U4yfIHbmLmVIpM2NJCcGi7y2KhBvCjymiKzyrTHvdLVdyYZRlib71UEzEwR5
yH/5qOuS85EiKSA8j5kYyi34N5ecrLkOYI2jgp93nvanpkOIH4c7EfwO0TNy
+Et+1+52Y+aYjOBjo5+rWukqZ4dl9O07uBEifGQsH7lxwD5dvvqIWJeQWLdy
yoxU8Kxg/TLpzxvgGxpMVkZdciHu6/74KovRBFTYJwCcXZ0Nqv3wdVjRbsQ8
YWbho3IG+8RoFYZRRxqgpmp9hSeAx+2womRDRFsFtAdQpvq+xOWIdJWT4WrF
pPQzFz+VyzimwI1Jrr/DJfuHapXNFvh9w59fqplL+Cx4j+Qq4Iz2um4bFmW9
Q6trg2cr2jKMUrmd3GpxmumoENm6MlQDU0kIaSW/N/pC1dpUiwqfGo5D+yim
0aVtv/KGjYgaAZZNNA6IMBfXA+/dpHI1ovr+GIUFc5TJMt+jmGvFbB7am2JW
s1Ko5n9DChD7IMVNjrAV1WmjGb3Qj5SyGZquPTawk9G1kp9UWi4zxV97wIwz
JpGyQfH8zPp7OKoC/HNEyuBp/XDBc8cwNMlRsBMJu5eKEqzIKGmqpo6mM7WC
pyoNTEVT/dqkV5lFikD6Cxw64o3xTtdUtAYXRQL0IGim0ijMXHPkIfLgG+ZD
vMZb6En7Wt/vY/SEoaeVnd4a7usddpWfKFr/J/ra57Pn0EOnLY7MZMboZgHn
o1Z7J8LdfduXVXmWRMDUtzBY3ynjD3NCdiw9JW2p9J9Ojm6sV9+F+ioKCfq9
atbmtFVAXKkw9njFK/PO1arCT8pEZtskNbeGg2cX1IaUFx7mNJaqbmqB1VeY
H4Md4PMszUxLfH+RorHhWEbLLHP9PgbwYhgWgFr155c1zrqaWbRB3rsKQeJo
ym9IYtJ2WUvjPdDqLsiDnR6hSNOZneZQ+av+KTLq71PfkeYFpWI79HPpyYD3
ijHWsmtddmnUXRTZjnvjTTWKQVcbhVZnSabplMlTptJY1267fhE3fpmRYxKl
bRM3C8PBQsKdSlK0XnoVlLmDsOgY2w+ec08YgUY9BeutkW2p8MumcAhYCnyu
U80AiWZC88NPNKQUYtXZhEeAmW777FbMErLz02LmRckrb/Ph4rJQApWer+bG
ERmQHf8W5Oj0wgFiCL0sKRhl3li5gaUOwe2eg53EtUbe1xsD6VHzZtxarTXn
G0Y/Ez1ILZZlxLXi+g5YHRicuUHcz67G1kV0JrN41M3rKujoLbVS4KSEriAM
RqQdraIA5XKusimr2KmtKkkuxPpF6YHWrldQ41+tLLWy+Xik9FOz9O6Dvvnm
ZlgON0XndjciOqW9UtlIlx7lLrWnTOP2D7JY5Bx5gzvtUclDjXyeAk8J0fEh
gg4fEowlP6XDW27c1XrvvSaU+kf7XP8tzjn2m+zDMFJbjU38X9PtiO38eL0e
Rp23H6BWw7dmipNiM9nntjNBpt+ak++UC1046XthOcD9YPlxkgPqqk+nr65z
w2gnaFZmQK/wYPOqFJbe6Gb5shH+OWIK9lHcvIJD+arDbL7pz+w0cAicnKmN
ejb8Ev2jeulSf6V0mA8dgM3kPl2R7iDpSYP0lnO9aW15n8q/fZa5LCwLONp/
U8axZPwg1UqIDvNQ0pSojcxZxaUMw4wuHqGYcbOyUXFgKAQaG2ZaBJlSoOE1
+4VjC7at1CJlFsjh2sq4GAYmcYq19UWBlmk8kUe9aMmfmjGeEdlmzxEyZnFY
4LFp1Aubi3KVarzymI63qhoglEIhI2tj/Vp28tUh5x50yZkHk3DZpquTaGGJ
DeaV4awyz6fFrzUHGAHHeK/oueRZNQjUwFBqXpz8VcMnzUW8n+HLd0eNyro9
+bJl5D/4h/Ecufy5CAKvLExHlJGFyoGxbfbJtijdkQgrWcC1I60CODP509pJ
BSghnArR9cDR5Rf36GvtnJV5uQHUuidj8H3OvmgIkXv7cfee7ovv4KOK9kCx
ZsXkdpkc57Y6qv4cvtP+FvxnzY1rkVcMVR2iuIOKse40LAgFCZ+vIj3/DTuE
Q0tKqYt6bsumCmARSn6idjOSGkWnfVz9RQ5Wpt5Ruif18fri18d1XLzujaSN
5asGfwJFBOuzYiUskgds8a9C7vj/xsME1pxE/mu77PgYrv7vqsrFUSs5MpUN
ghhsaNhMvJqQYJhxCTq+qb3CwakThgOmMyZWcBZxFhXCjinbtkuT6uq1Vq/J
7B9PYEP7YIV3yjbAw11gGqkBRcmVvgTamRTDsv3PkrEu/eq/9m8D9PIF6Zl9
WKS0WtLde9vcbzRji8mdwSA7AC2CrY0pEt9RYM3HHbYVTNesv3GiqeE6yJUb
TIIbyX71U528Ef7q3f3aT/EPM5DTIBdIh8cIwwfLQVlCOGhwkBBwFjpNOemI
+QF8xILYJCi7r1T93fqptoxssNpfyMhBl1eeSuVxd5gzeggWiLIVDKqdWcQD
RRd4vTUdcYSDyOamYIGkTTR61maHmzALqfEoKkK02/lq9hzkVGV3RO8avFQW
DBhbbPN0soIsiBnMN6otBNp3xBS0dTtn3O2By1zv5E8h6zDihRpdOmGu0vtP
dbn+HoXRf/gaYzuMGk+6r7qthrYY2yw9meeOZlezeOl0d9YVIK2pskaKkEwo
hnU+99xdjoUk136+1x5vgqnPKuoVSoO1/DFoehh90QSECVtXpsv0XJRkhz9a
zA+6ZiX4GNCfqyVVUgK3DwjcrBuwLrZcFQOgsApkU1v1/C6tvrxcX9FKOVlR
ZEurlo9eKSzgrfAGMgMWRbB0IpPRQ+htlpP+IcvRLulEIfQasGRRPvEpsS4J
mMj0gOiiy/YS4CAzhsyjKACE2/vVwoOaJmP0guUSIXobhwqozURqSQRp9pyf
KCi0ZipOjrwk0/Et3Jt1bhUgBTJNwSjNxpk0hr+IXsjTKv6FiJYnIx/keqoP
QRh3o8mzAcEw4VLrsN8K+VbzGbOwYkX2p4ZxoW+swAVUo09yKKiWw+69cPbZ
Oq8VC0hBVp4tfBwTK1i1R1G5mDgCiudajT6j083XqYsSpqgsjXi60vkDVv5c
mpEw70Pp6fiYirUEf61R4xyfM7UUavKf9HhKRI4epSd7yggW+q6o2vxW18U1
x9lPKU0aTiXA97+/wQe8QvFPuKSq8spl7fDN3Spr1LL4pUjK+qeOQATnJhvq
x3eEZVkmKYwrkFSjUANViK+FgXJ+tPnIdA+calrVdbtT/M8vtcuwu9Se/XSJ
AqpCflLZGWAe1vkUS3QHTQZC84B/8QmLCAvF+r/fxsJuXJkTDCYjdHo177P2
K4WtpDLXUT2CcmR2LDKwZs5GEg0CoJWvaIx1hHJOvyIJE5u/BacQLdbgso7E
Pvptyrj3H2fbC7AgRQt/I2DmfGR/jLDOYYuAW51DaUh8UbZdsHXp5QjzAZ6s
6yLwb21lQJMCRzs7oVqW6csiH/+pOtRNVeqZl8K4i8w0LxY9tH14anaWBdhW
Owb4uA7HGkfwUCplh4YacVvRkbVTOBGuVik+MeN2cTPoLQF0E3ydHYbitlwu
Si0LvQOhGJFSnMGb7Xl4rBvG4cd579FHDV1Sc4JAV3V1p6hmMhi47NJNmqLF
GC0I9G0NxTHZI7FNhBsOqKLmurB8UO+4WagqWOllwXqvr/2gIvvGfBI/d3yk
bHUd8JHXeydHx6Bpwcu+bfmUFJwkzx8yhcguwXiREBL77qokyvnn9WImXtVE
l5+2NWs/YDBJCV5a2LZVjd2bxjPokfUXLAeBkIt2EUIVFffPSmZUQ+uJs18l
3pKY8mHe9QLPaJRITBuUaPvY90osC+PR0jIjdjc//ZXI7U21mLfeiLrvnJUO
xHRUcJTdr1l4hbw905j5gzlYAVZDxvgLm2tSMw52BNjbaw7YhqMWOo66xi1R
zBhoEM4gubBuQCGqA5RclYpaAopvQEtvz9UEeuC5DgpNe/MUSARzgnJvwEut
dP/LFZ3iplIzX2oXlVpF36vZgTYF5wZZbS8jcNAx83ooTFZgm1veJwBiBJRl
G0/e/uq16ztai4AJLTqrlS0CoKVuOgOgsIZJBYclm6F7i8Gl46tWrjFBfmBY
AuW1U1nUQNwGuenBO0oFDUS0AwSjyUV64bIvJr7oIGF/nUTep6UKvD2YVQzz
iqXQwwb0iu21xSY+ZrLjmElE7lplNzbJadruYY4QuoES4mWrr5AwuF6/LzM7
MaIFla/upBg7QYczHi9+KnYIiGTMkgfvs/56NhRHTSOEEYqh/1PU6IeTGK7V
qt4/M9OByLfxNo4X+PNPTeIBbJ6ED5PLySgYGTR8mFyo++Wgl78cjXeICXdj
tx7qgB9n4sb79mtTBT77ecikK+clpYArJUOXI4YxQlVgJxzQp/CMokFRxcyW
dqisgVY4QcNVapgGAwwBX94s4KNgR80t7LmvoJ15Fb8I0XzZfTxbhB/0FMP4
eEj9lKL4XJ6fHvPOVMnOZ9S3jQpvL3+ZjlLrtj0U7ujOhUu/XyUuJZKR4g1f
f30atsaClHxVj4eal5O6iBim2CajMNerM9QH8lLPkmFwQ9eSp9derylEElsd
O3QTqSQJUduc7l/hEwwu/fJ+p1/b8MD9h1lPXa/hA15j2fQarzijt7N2pPd2
CKoMRH/ZuPJN7Fx9gWMEo1dGidPdcrIFJ/ZjvJhwlm424jLETkm9fPyzQY3M
/AlrdFRzBCzzZXaWg6RgjQTSsmXTAIrev+4zcdcASIyIguTA5k7f7ZZ3p6nh
rfZCdIFrWHLCcE0jQb47kFskGGc1TO1TDkrES9WmyLUIQnKB9fqOOMQUceB/
VkSv54wgqWTVL6oPBEpnijnIWw20DgOU3pl9QlpItD4DKAMGeRnjcS5A3Q1u
6Zj+3a/gQV7YzVhz2nVZOGhnkCHVizGlF5yGdjDMT72q/ng3hdVUToPSrGPp
A7kDF7D90R+L6tMLr93twC0oYIVW0VG2UqikrWHncpXyp5TE5YrGwVlPfnNx
xkDJfem2PchpnTHeiV3QbsVkXFGiz5z6OyhxxiQaN8rYN35H+3LcIVSpVXuq
/uelcGWGIhG6Pq4kPdccM4z5+gN8uxyT5CFbd20o26YAkINHezfnHxxuVW0x
wseGzt6nzldMPvRI2YI0SN73rrZl/j//f55tQM45RleXM6L7uSIrk7eoHQTT
3I2LmBMmp2bBTMLk5KK1HynVZtbM0Lzhx8L+bnS54lPfWhr6qcjyLR8zKdXO
PWka+u/Tnl2/fDNosFsEHxgF6KWMU2KXznod/chU1Kyy3u8cFgrMCvbUtX0N
e4QJd3TpLtrHsDaUZSlS2SHzELZeyBandOc+mG8ZXFyQQ5u/teLLXhKmA2N2
MhnmUQeiI8vgIsWnts4w5Y3UQ8wlpjw1ukHuYMbE9NCPF2babSqgbcw1dd+Z
vxZjwS9bAfwxRDqZKEaApdr35ZmfVgf94BdSvd5Wi19PasgWr1QITFfOlyZq
vtb3uSRyPFRymuvstmyXdsYmGKYWZC/vbU8XxYsJDn0DO7kv2levk9pE25ki
GmfUDCuKlPMyVUHNVxkGnnmxQlNRaIjAO3DESa7Y/Wh8L6eqo9vOlGS7hmno
bT6qa3hCxnToPYHmp75he3IzAMrTXhwvtqPDEqzpj0nXF2T31t2jQXLAf1h/
ro9TfDXPpWM5YfSTkT3RFVBGkfdZp7WrgWeWVOQpje5AZbkGt/hOgqOfXPfH
gvX8IBEBWZmnc/Haj9XSHpenOUpggATTDxkPrhEWCoPq58m+OPRxSJ/Iq4PN
ejcSWYQfl2LOdCd8zKTT6gjkzCGSuxei/6/kvC8XhtbuO1qVUoQp4mwqGplB
8TxMDsOtJj3EB6/bgxRFfCcKzGIpjTEV5SJLhm4mY5yePvyIM4LCdRwOC89i
HRxTTnp/Pvt9XHYGftml7M2zddNE5jeOYUaZprz4A8XpYmEQuMPlE+9dPYSE
QPyAh1aTpGWEhPrN1uatfH8nRsUxU6Fi5rt3Bzzl+PHfSMCudIkibGjSeZYz
dnHJ3blL0m7OLe1Ad4dbmGA6S7KkFkaDinHa06whQ69LvJmpn0CX+3Dt6qal
lwtgdD6BnH4cZm5bru/wauDV5U7muDkRNxpUJuvW9HJe8JPcKZWMU3WI8SB6
jzGIl8B0pDnWKDSkeJyROMgrc9VbL0spGkPIQVK+81iySzJfsvYB+s7GHoDH
cyd/mcnMbEhmokA7cfAzNunGcoJTesxWCzZR75pqAlBAvCjVb2gJROCaNt3q
ymyd05TA88lmjGKWlJna8VOhoyCZEQhAZjXLB91WaiwHiTK8OVbgHLfMC5td
jA2TUl1KSXWWfy5ODtuwmBVcKjXSC3vMMYoLjKkLeXWM+XBnkDmmS6PkEe5h
XvCaCeRuMM6gmUIQzSM+/UBEmifeObVZyxgFGuRaP9g1QTRod9NTpm0pbbhh
zN4g9kc+KB1u28Sw9abQKHO5MxyL29EW+A+ngAvvhbNDKGQ/QPlrCVOvZCkG
DpGF9bCFQAkq/6m2GvXSqkMNK0SeBxHdyG3bT86QRH8wvs01EXan+3cXTHWB
L4SgoLkdRtnihwZZMwh2/BScSnnb5bVhqbUGYRJAQ57MxAj0Mn2Ek8Dzxzje
dFs396Zs3x6JQ7s7pLWk/kiZHbNf0MzLeWOV29jKKOrZ1RvjFCPnypj50Ei7
KTNzQBP8ZRvt8SNVWa8q3Gn5Dh4jbfCHDxBsrc4bfsJ8W9HUp1yfAFWZWCEC
NoA/GdkPRUjTsJ6OJnc2YLNXvhQmdAkwBPbwbeXLi6nDLLjyMsuSHuYQ6DuV
q2WUOhF3bTOnF3hh1RQlQFCEOQ1/st6Qzz+qPZX1FQCmeeg9wCp1VfaoSLKO
03588hra24outrTaRT4bQ5PUfjgAuO4dRE27FU6H29RPSHxqQTV/kTLzfNQJ
+/N7fbaRCca8zZ8hD9ZA8BawaklX1YdPeKyBcUDfEZ0vmQ2grj5QJWtZm1Bp
6KMde3u8VI2rUVnEB9Ddc9wdQ3fJ9Sqr6DL+/3rDHqIuxUysxp20btlXzVUH
NoPoq8Oqi1kVYExONVcxCpWn6PKOKHnJH/KV0huWvTxSp0g6bq4XSZ1eccwG
Pc6SGrFWNIeYrb+XM0g8Ykx7JUzlNF+FGcYcMjntlqXB36hp1yNudr8nyZSX
yJX08H//mZ1mXcWlPERHX2kyikOdkQpCGHpXLrnPeZQR300oxmD++wFRCY0u
Wxel8fQWO+X16tLKVac04YKpW0/Cjx6Y0fWtU5VtBbUK+CfZtqv1kFG1D5SH
7O+w/+OnV2S/PI6Vfu7OA5BMWfRCpsAyVd8UBobqkSiAi3uFEGeSzltJ5Hr3
afxdtDozVH2PRYXU0873FyuvGvhc76F/J/LZFaBjALTy95/V/vxPHjlt8HNa
2KGHXET9k7TNklYvERFd7nIiaSTrinIhpYWveaLcPo0oQSlQ4bHkYceYCWAx
UesTL5inazMG4WHJCx8UhHANQ6XW6+JCAkw5dR7SxJoeh+8PP8PvxhLPgh9Q
zSQXZrQW9mOWsPhWJ+viTOOhG1pK9LIpB+INmeO4ELGHTXL/xjzHih1p+4jU
8NYrlTRxzq1ekaipr4ruIN9ALsNmX755ZmOtdm47EtZTl444XpD/hAMROmsL
HTn8i3WF1hC1a9SeCX49OdhsADbhFyUNWfOEq+/tdzUa8uq6qEh03PnPIbhe
vSWFaWKqt9SnuFDi+lvG6lUCdpurcfijrHjiRZCw0vvyI0O9M78Dr1Ra5vdF
E1owME/8Dh7+tXIe/tUuBQcPr1h3/78nXiCvSlPr1HLRmwf9TG3kVy6/TQuo
13bwAsh7kScBs2GtbB1uJBdIWTvBjSSTcMx0iiAXvHEtRsAZWPZY/d/nB/nl
LXVl7tVDLu/VRpqI0F8hkAVHFpH0m0i6ujv2RH1Wt2ENrBq6WR60jWmqFT7x
FVNpNqFWGYE5AMr0X1SFGrlOr2SzZ3PMHbRa0dz0NkntcTWd6LOoS2hW90Vq
N7/lYOkjbOu/+0tQY4lTpu8md9GsUehJEibNCimw+KN2InhGv4skPSKF55n7
PHpA6iYO+YzNuql1SL4OhxIMc0DiM9hlTCGWGCp5+kRA9zWRbjgDtqd9Kq5X
V4WQEgiluy6rytICzS2vCcFtG6tHpsqbz1ldBXIlkiH2TtCWns3NTdFhrTWw
bKHm8Y7Khcp571Ir9SSmOoLOTJ6iKnj8W5rnrfdBAfFhjx3Xyx4fwZyvkbl6
474AneBErBvikGNtJFIxvGeRdSnyra8inh7lv4+xx/xgbeuIym58EoJbxjod
CZa7SQYhby01ZiUe2WcKTx1IMmept7owbEgy4oNCvA9LG8cdfw47JdCt8J3C
lKujbSdWLRmFQ3rZ6SyGhche0oEb7g38bG+tM/9t3Zrgo7zIoLgYxd7c1E7Y
6R2ZggZ7YBd/Z7z239LvaFKg/eO2a/SZmFmDVHvHTBF70SpB8g7IY56oRHzx
0VJu3SewWu7usMPS2VbVvM42y+kXop8ffMNNYjQTyMxxt4GB3a1Ck+Cnn7+F
P2jHVTyBmsiW/mt0j8WX8ovYCB7cnFybXMPhG7aoScABUH2bYQVqAPIeStJS
a02wsf162jHpH4qyzie26hTszBRkidEW3ftYR63mMT3LDHd7etSF2ldjj8wb
Y/nDabqAYLmpy4c14eMt0n29wWGR0ovwrGPX2HL7TMh/lDEyqV+2bZb22lpn
f8b2CyS6g+ApCUFZxx5GDZeJLq8ZUaD792SqWTaEreuIk5+eG+VzjPuuzhqc
4MmBobHBKRhXZMK4/5nhaWy8Ny0qWTnx4kTia52DopXRpLXCnDCp+iWU27uX
d7XA/5xQr86uYLkxzLhvK//jdOfk+dPOqmrGfvhK5x145S+R/I6dUU7j/Vpz
VTfTwoXzJvkAN0Qb2DbCrJftxGqKy1GyE9hkBqcWzIx3lLzE+0fh5Dz7VoD6
DuYS465fwqRlsRFHUrhU0RbFdyq9qM38HmknzZTyEgdfeHQjfpycJHZOv0lT
wkc3lZqcK/AjifsnaDFyHv0j74rIVXGAv/Ve3/OtdmV4WpR4awffNxupJrN5
7eUjmZo8hr3C/ARD3wU8/bduUN9fB35u3IERLV/hb+ftcIpol1L6H8T/3M0K
EhRUc4HYj11UFVgDkhh6XED8T037tVBpkp6O7ydl2hP0v95jNZCGx8e7gcpY
VEK5RuL8wfoSXGQAevpMM2hKYtQ7Cm0p/pp9E5rLt4kwcjbpwTaxEp80qsKV
JtZhV/3dA2NTrW1VwHUb/2G35Y/MuXNCRdRMD72g4MsU8I19l5SaXQLdFtfa
HSZzSvtLZ4wdEGwxCl3MwXAyj8w78MAr9HBTQ9NGDWZQ7pxAPWVyhqqagWUG
3VZnOAUSu6r25UUojlORgzO1HJ1GBAhEWdOdo/RRkRTcC9k/IpATazE96WNX
5+y1rX2qNN1wsfGZabdvQ/fBXkFw4q7zun+AFeA7b7xufYBPTS9+UGt6W9iY
mgJQex5zkL56hxBy0fGf6je84IiHib3VrQ7uWMnKe7sQWq1a2KSSLCJjg2iR
VJv68GfRuHE5KXzO5W1fc0Nek/I0EtsXjUYZr1WYisinpqwFeLLyL5qn3U8A
TaUkbwjXZ0QrZQGe+5Cc0t3ODP/o77ufh9Y8IB0JeQLymP+liHuN9f7YiYoM
Dox5a/OKlnrOxVfUM3V2c9ZsN3WhmAFD6jh0T2FixSYI8D8aq+siHTtnISvE
jAXm8KVnmSo5mGFpII9cluaxHJhGraJ8Z01XLKTq1e/GK5aAR+Fo23m6chWo
LJR1ZvbI47FNSVq5wBAmItdVcKNeo5iWRd7pvCF/Q5WVZw6ora4YAW70oDLr
1e9sPyf6CJBA14C6tvBptVmDSW/KDZZWtLmpL+eQXXd2yC3oEBckhDS+H68z
zHynxetzyDluz6fyWJjZUYWPcHB0kAJy7isYhG18Yr1CQ6RuU/SAdXIWUWtH
KUgSSvroZbfQrlzQ5EauOKIk08F4FBM+jfoErhYvgk/b4eSd9meB+eFMhauD
0zMjWkcBHI3nZ8IsqqMdJJpKQhBRg2GonqimdCscbS5+CrQuqN7IgLBneOxb
iKmUUCdqsVC9NTa0WyjlikOnBJClHSzC+jfil+OztHGs0EAVtp0XU7c1r5VF
BjU7L6kLn3jS53GZ4VPezfst6OrMkFH80vmw19E0xfqtOi/MUyU7JeK7fSh2
yjbsWkg25WSbkojkAuVq6+ALEdGklazjAOdO3ByT94b1TFnmzJrhfPYuCUoV
jFiFRwxghrhB7124CmrOomJ72JgpAq8tiLeHHl32Ak+Z6hDpfuF3OFvMcVkY
rLbXsec0lGO5KUYJYiISsGS83P75vkBTMwqEiIlkYbbiM8Xb/WHiDdnQZWtU
NlbyUnuttNEGbWT3eqTiV5CQdf3By2b09BHRcuo6wJSIDiBsUGvq42CwTuLp
yESomPiBABVmmMgFXr4eFpE0ZaEG4GLJl5xS/5KyCdqaLiZnA6D5Xwva81bG
KMlEuonTANeMyyOTD+a+6EtI9qKZICcjV6uXyAncbQ+pQRE9XEnUzh5IOFll
Z6BQayHJhkj91m7F9dy+3eWRjdbGkXfDbYSWoKm+0SqVNv8nmJlhXgXr/FX1
nLK03bd2C6Lib66g4iYBe15R5ca9q2R3yb3k3KqeEX9+Jtb6+eEffq06I+8N
2avzURDVJQPfdracRF1mN4b/Mf+gDSNT+vuI7EFTNVftLoQ/MBZdfM/1JYb2
uXNuJ2zvtqPoCvJ57FdOzwuuPATu+oGh5fWz/2wDd5kE8jlEr4VMWsVxWWum
4IIhJmnN1XJMJKSRxHTNndHnpeqZIfc8HcUDnpVgM0utQ2GW4FkKEGCpB4N7
kSLUjJKNH6N1Le4j2PORf6BdUv2F/jxN0wIIsjvgNnrF0/76wA56XDO7crFM
yU7LDrc8FhmOTTqo5OnSDcP5DdBPyvE1pZvUfGH5zl7okSukJXu4BH5QMQ55
5IUrItZ5aa31aCzBI4PrEMsNO078ZX4yKwn8nI2RO69Z45KFQz39kTWiiSD6
dYRCV86i67K1qQ1plKPEXModNazK+Y6QbP4FeOtflpjUh4bSm1MayND0zOrk
KUyTR4neCdWohalH5NFbEgnVFufTUskYWQ32lzoAxnCiqkOLC3ZCl/jgfnT+
0SB3iexBtucHwu4m7WNhLmDkA+E1vcWE/PmD8NhhHZG2R/2onCH0vi1p+Efa
OT9162KJ+Vscq9nFmRAwEYIUtfI/gvF9G42IDNEZNve13AbkjFrLZhHonsxf
Hpoh0yXVqaYe6pyhtfsxgSGGOuJ0TU7CDmw17Zty7y8KCgoGbCjxzfcz0cVN
LyGw1szyb9hL2QhPhMLs+z527B4YAFL0jglofClCNp7tdmnycPxj+3Vo4dvn
gPUrdY3+GNCDqJycjcmQ0TgC4QkHg13pRHKcPqFIs/aXlFbLoam4pQVvF6NP
a8vIUUkwA+/+zFofDe5KUpNKiyO9ijvCXgLglz56JiVCs0lr623CI8m9AkmL
CyZLZBbmc87ExazLh2561lFni9vCH3h6fcwlXLZpCzlvsro8pAoUh/XCqHtn
ytjXZaio2MCNPBHEUZM7YQbnSIDNXJWCBypDZwgKwY4JsuCefMrqsEOyK0Rn
oV3R02nt/FBADfM3oapOw244s2B9qNDGexJhlr15mjSoSk1EkIa2UfazOakQ
RDw4gs+2uZ4k073wRXtfu4+EyXSaMyIDfwZYHfkSAw+0ahLSfs648/3tLI4V
yqmAFuijXsNrfpw7KBUsXzxVh+zJSdRTeUEgagaOX+ytBzV9IE7s8K/eT85L
mIYrqEJg4XNeB6iA+kL+MdwfZnYNn1wju6YjKt/Tp6dI3UxnHl7747Exh0NE
Fg3SnUGLyPl5MysPVjHsV3l1E023MGFv5glRl61UF89dVM164kIO0N1YWTXB
Xrf1SmtQDIam0bvMgf9qQclsUbBgxAWwkqX4gQjVg9wTAPl2dGQQSEsdlQ2N
sy8ir2UmB6lI1/NxhZ+oPmrVoF2A1MQ0cxm+/m3YVQMnsKPbID35MHWQCIbv
VyXqckTJk1sB9l9smPqlgCiwQMM0mCgGriY2W8PyDt61EYJsUYQsCazTs7XB
HtUtZqzQIxNCneB4CFp2WEhCTGxFHI/QiuE/3vtlbGBBa2CXQtGrJKksVN9o
bc0VsQQWQeVoiyX8C1pdzoZexbl4g2zBrGvsoLbuvT8Mutg+UxZVu2zZmRMf
sQwYKuxsHjPAvoBGy76Y8N2La33tmUGRHJuXP6qq6qBL8j96OVNc1cKIgusg
nqvnO5syyWvAuIE3uw8t5lMKuXxSSqFcY1hxI2TY6EwCZYnG8eUERbjKaLx4
47UCrqTM6e81fzTE2gjI4VAFRk5hlARgRVH9JlXzbUgTdaAbuL5BAxanPTFs
8GBvU1bubHy7NCKH4WzqyCHv2/v5kTeoMKdd8KL0fjp0RzlTmnttpV5bkl7p
tZrLX6xxsjO8BGQiELAmokgDCdw6eB9QW/FiOZDKOfHBm/ZLoi5BbDpmMTPn
G4rI33mITVpJj5oTH6gX9tnk24gvx4CV5aGnVVcTWQ29BpkxDkqoLD0LMN0M
ObW2zEAHRPeLZTk4MDeqRlyhhkeCRbhGhx8gdM9A6+X/06PTARDpaxb8NQh2
shc+gRNJHnY2GJUGBgk6YSFSYcwV2TPSx7b1i2RgSvig1c8xHrbYUNuc0gbU
mdL5k61NJgmMUaZeanas4yJdIYGjOzw4ikVsrRD89wDIx2dXSavor/yXoPHh
IQ85QRyoABK9JpHlnprPkcEYv7l8RMDa0nVGa2qFDlt4sgruMMV5cG+u7IA2
t1vlz1q1Kn1pNi3Q4Ra9v5XFQ8VnB/hd37b4ZNnoObU8Mj/a+74kwjLkyLQy
1SfhBctPWaRnMUACpzUGGxHEM5RAC6jPUGmRmsbTv58S5iJvOx081o+utRys
VwKSk4sCdRyLJ6+HznLb3GQz5Ruc3Ba1q++VBwT6aT+WRvPT2U4X8CvUvoAP
lGLorEJLjH16dmVXVLKfrjvHAfBPXLQzgaeJT7MvWkg9IaiIQIaXZfu8B2N1
DgPIN/K6SNwATxkSXW8wYe7sde1vx5pdsRbkP0Gl51hIGMeVUD5GoQYQJpl4
6wR4YRxz/eKXgY1ioPnQN1E1nJjdw6iR57Dj4dQ78gqHSjo5qZtEA0WCzp4s
WsP/hvl4wjaHMEaM64qGzzn8XFqp7PkIBj5voSCS179H54GwIl02AsZclnJj
AVmocgmdh5gty/k0ze/roLqAFZI/78TNU2C2fPRQkchEbYaRlVqWt1GjmFMh
TyUQxqaNhhjxbS+jrVxqK4BmBzKK+SN6Isq8o0G0BAb61eNWqEe/NFkYAgTr
NanBiu8yLsF5XSI176V0oBWYGtqZHR7T/7iTIniAtG54O+yWVBtxqn2IgUmB
AWptzqF2sWpzDswskswkQ6PEXveIawKT3BzHTYQHu5wNWSrpc1/T4/BzO1XI
Sxxjr2Zm1pdRRvOqgTwm+lfeqj91GHIzzUP6sBzAGgn8EULK9nGwEKMl5g+H
Q+QawR5NmWKjs5e6THYxWnF3JMXgwX5sA7N0OkSlMgmJ2HoHx3ILgKMEYGVR
sz7eT79fZW+glWgTIO+XN7yPIzsRaeyDoFkozgviAnPCQpMqN7SX+KHyYr0+
6lMW76YNmSzZaNC+A1zO3UmGb5/mEegXn2oiK55EXKoVs9Bl3OLPe1b4AYDW
lv+Uf1VWYPp8ccZrFmSe0nFDhgO/CSoFySQOjUAd34TiVmZM3TgYhZQVMnz3
xv0zgV2c3yJihY3jrsrALPuzETmiAu4UTajwJI+4R+hh5/CBeeBZu0tQz6su
Swz5YEpLXebQgJHB6kXzeWIarfKkONpYF40Z+9JCzlUTQR5OsTX9dO2XZHFo
FhKgGxW1k3l+R5Si3KVoNwVrrJqAeg+0OEb/jXVNasROvMhyFEg2+dBIvm1S
uY8WKpMqQH1gegyxxj8a2FDuBRr3WAhCW90c9dFdbwBk4TX/NboSR34ztyP8
XWIhStOyL5O7OPACqy84YkzBuQxiSoxjwLJfZ0ypZMH87mV1U7ooEiOw2NQ4
zdLAuLauKWeyPejykaEtqNPzYKpAMGp8k+dvSpXYk22HFjkgRZdmsqSQCAjd
zd7judM9dOnc8ghT4nCWgMZ3tYY+nJbiN34Ikkp4pxXvXOMNY6QV2adurqLW
3+ZCYQwU5z3RZkJBKRgzmFEwosqOauVpJTsYL2ZCFxfJRKzy912WaoCqgg9f
e8x/c7EKTLw59wdL6XQGXeFUxuou985T/5e2H1TD/VZ5qlWLvDpqvhvj+NJ+
RVe7T7iVCSMKtU/GJ0vKKpd8Uahk/gBDKMinjQDrkLxiYfPXC6EfRv0h34Ao
yY1rqrwXEqJltou+l5//ZijFl0sGAj1e1wqmwz33Cd70gqgMI3IyWbzflxK4
Wyii46f4G1E1JP1Xsi6JMacx8OX4zE7w2bmtLNnId02DAjD7tolI1oCXthMd
mPctrcobie2kgeFxQQs6Z65tUIk2Q1aydhmEQAUhtqQJN6IESvHPbhbNtp9+
YzsiRd40pe56DgafqFhlT9isWEs3SUC30qelmTJh5IgCdmiZXYu73WwTnUKo
idiesT5C6rZfQdHrGWfb/kFZMnRNdLTnPRdZXDnceBjLTDbw9LPnkzbKKSwL
Tisd4iZ4ZS/6llugrNV4rpZxBsJCdnVfKnJugtSRJMR84BY6EHeKurUv2UvL
KGN9DsA0fCa/dpCn8gcXRPSfGvz8Me653q+6kOJaz/zRRz9IKbwS8MQSAO3t
/ul0ET0dxTFmo6rh/XqMt/3zYwONiAOYJAt8fxzThy39Tm5dmUEDcmREmRBP
CXRnrLD8PjD+1sJvlZtyhrvD1gjRsNUdmd1LY5+7iEKJb1zsFgHG7LqtumHs
j5jBUei+LlNUkl3Lg0KeTNEKMZVbf/hQ4EaToaLwHp+25c6ASYuYk5tzma/2
z2p9PjHb+C6lKtHQzIS/M1Nii+GGXpG8GeUCqVi0tgmgUJ1LbR7iWF3ULBWk
hjKqAIK9SGzUes36moA20oQb0LWM/kAPGD43CF5eGzNTtiVKMmrA3pnS1gkN
i7R345mvBKvmPpfl2MU128SbbYXLEfdRKwTUdvNwQcLV8bYsaZdtvRxVOd9k
z2/EEyWCKWvgjJN9KQcsis2v10dU67Lge9yVh7bnabnC5tKLqKYS4CcI3/sX
Do8xjaDCNgvCAtBzaOgQ+QA+ci2x+btDzwKlGu/eNKX7QpWiURljZHndm4Z7
7jwoG+vF8glS1yprIhTUppZ2kLt+qnjS/4eBuiIcEFpTYUvKLiDqkHAfFFOh
2EAwwkO0dfzv7vo3+NyMS/UkYvOM/oFaZU7pz2fFpb1WASWYtxG1LmLOH5Gl
1m4vLL8VmLHCDjCOo50UU413zr3Qs2Da5cijB0HzH76bn2a7Qc6JnSTt4939
PK+vot8wiql/8SplPIWv477qHQNJkh2yHNvtToL27w6Z5s7OdVLepvdO08b0
WylcGQ8OCeF61pXfu8N4/y1t21TEgOdVnxRnprnMNedJiwg31HbPw2/ncP61
xCmg0MekCewlAMa7iys56F1CmowHDZKupuD4mZU5c0pArqgbrqyY1CUM7zBJ
yxtibsbAYCV4FCZONsle3mviZGQkOBx0IPj1h/YH/Eusd68ForwhcCNvQvRY
qL591cCcvupU7aeWvdui2jDK/gHQ1se81RZjNr7jqFmkaawq+K/iGwDZcUF1
wK+yxU2hRLway95ji6wVGrXvgzWyg+V/h60PNew0Drif4lEO97ZB+HeuacGd
Cf6OsyCyJl4P07Io+n0imZeWeXmMPH+WxeIeWlmzNOUL78LBkP5wOuQGzMbX
GbH9ZuhKobiaOakn5XNSnrnfYEZ0Go8oO8Jx4+YoNM/N4/wLgZnLI4ibD9Tk
ROl6xo2Coscqy3dz6FpxTOsVRiUyVTTaiFl/vYf6g3W/emLvf+ibB2iMEKGs
KKAD/xWpSSFAFLXUqRRoOO45bYOxvilI2K/sRdm4gKxW3R9ema/ezcyIndDy
cFTT1OMNTQ5L0E/oKC+bckFqBRHWiO8Gw9+fKIKDKNVoyfBoM2QJJ8zCatih
8lTTeP7BetYOUZ1DDOc3TQMHWkF83LmVy1gOzdk9sotR4TQuTY9z5Qj+cDhC
aIe0SpAQdFRCEA5kRjvgcdkLkq5fYp/QzXkrnB6bAnF3BL/G1c1rrgFXK2Kw
K/08SNMhFhlRKUwY3Ronadzlu70G9KvHZD/9rlr7RhuZ1xq99xACcgkiQshA
Yq9p1JylX+IzLab+EdpUYoyRmzr1+4aloO3k3592hHQh8UmMpQmXk7i8twOw
aXW8CdJQagqn3kyc2fnEzaZ8OfkzhYOMpwjpeYKWHk/93jbUWnctzfS5iFpg
QxZJ287cc4Xc0/YzEGSO15a24Y3/useZA9d8iDDDTZA7cmZ3rfUZJQZXJem4
USqN426DazWVWYp4P1LCz6Z5HsO62+BE0oKGdjk7/VUat8EI1itDg42EfrZX
XVYxGQWGollGZaftGsLePqcHouL3GlvY8E0RPHAucXBKtYQgrg0U2xd9+WTZ
GyKOnRBmCdrww1BfpNC99xyvXZ4XGYr6k37+IXH7oC6gfZm1woBHgx3Dx2Sv
1AX17geK0WWqn8shQGQZrkPlQd7MuvYMxHq1o6FxvbvAwM3M2WpQTBCc1VtN
GAH8aOxwnOGy1BnjcjWewTw9LJ2lqc3J2e0hUUsrvks1VTiPWL0liCHN9pm3
GF+RcxsY0A7OFZHL127fobpUl0X9WhGjOmcKI33rMuGe31YS923FP8iAxHrN
8IB1faXpap/6nAfybZkw8BfWBRHk2fEnKbyV7bOgFnmX5HhB6sZiqqRV1LKZ
fF1NZFuIQyl6TFu3wA8ML7+mNX9i67t38fa0xsy40kxBDx0QrNfGy5jH3dg0
KvM7pfLvJAGTieZ3A+sTSuW9Etmc/+PImif3DZQ3KUeCSHO1ISrfWdSPZywP
0UOvwqLk8V9Uly8B4WMTygjOE+l/kpdV5DxTgNqpTiBxpJ9S6qGESkHE8IpY
C90Zx/UOD4iXkLgCBjQ7URVmp/407J0eKYAKcBrSKrBplwLd+16vVPsLGRom
Dwzgjw2TLPfeBq64RTLouNdII9D0/LZn1gMbiFrGrUczVnbPiC4pCOf5mAhj
QlbMOSF5EB1wMbxtZ2gus9WN56hASYUMKP1KzbNZj24wArQlU2sYUhmGIXzI
e1+sJW6Mkv+/c+IxfKY30pUe0Srz84i/wCv+jaE4YlD+AZoz8422mCRJPnSt
/UC34Xq8fnySB99ynLr/vRR6huzh865GisGDVERPg5F1L9uStOzsyV8soYCk
lx83NduXhZUzyfVz66xyF4xA9WULvHkYYASWqN1FJAto15NYf5VEAxLf6bVx
uhL8dhqmr5M5tBZUx7Hb8Baxuwxj7haCz6A30o0YagNqRgVCyYYGffSHiCVj
VZr1GwIUWCc9W12fC5gPpZhP6zX2JmDm4li43SeXpVhw+tg55RBzxgkWRvG6
00tBOV+0pmflEIGfUgAr67fAu5YHMXBFF5vox/Dqve2eZ0QepBKllc5sPlaL
Ezu+AVdh6jX2o/f8iqd45Dxz5ZR/G60ot8wlix0ttjbJIN/FgkiFu31+KFw+
iWc405/xoufCuKXZ42uUzlTQYBSWNX8TPiVUAzyqfHDeiCgSH9A6HJUQHaBb
IEFjWOWWy5mwjleOiDDs/7tI0Im6LTbFBtEGon93W93Yk53TQxQnkftMSwiB
USTsuIUTzI55wPnl/3KROerN3ZKACuVisOGcYzFeqp5iCJPuglnwCNZdpDD/
iN0HZGnk3EjK557w2RvkVTv3rP8zC+EoS4Xj6KrKNA8hgO0Zp8EdXY7oeSnf
Dq8B99pjwh4mmS0qhzue2EqQzTSJMxfQIcTIGYVqEGpnrlB7l4FUaG4VQNwD
DiMFjf8bwzbMkmJP4qtWQ4Dn0yMHCej03xHvlz31sbDYGG+vuTl1Dc6hwQTQ
sVbdrrB8YVPoIaADk3pjJmCBED6zxWxQqvcxwECRB3ywJd3/CKDXu7c/AoSe
IyrwOxUeODe/jh696o7B/4AXaqKqBri3zKKBODE2SkUi4x4vTkCliYGroWUo
sDP1y4jwA9PqecdiagoPS5kPatSkIRdkyxyOoPqN4v6A6EfpOkC8gzcQKCJ7
Cwm8us7Wm6qC3+XhS5jMyqlJ8+L34CquqMbjgF/YEH+9edWOaEcgCYZ/ZD4a
3ZrG376pfvoD3WZRprjvK1xEqiCw4cAGdHKcErBa0HW7aLtaV3UuDqndLLxu
F1L2gTIVColSc0mXZZEdaer2wTvE975lat2g2J676gworeGxlISSNkUmoTbT
tzF36OFsApSKeK0ce770hxE2ZY9EZgKAwevRCxad3c7QyhYjPrRBQO28pShc
uU4rUmwoYnirwXXXGAbT4f/0Zd9iYs9i51XO91P3GTPVbr2V+FQG65a8nd6R
Gdtznl/5ooRKiHB4hbD5fS4jv8gJfh0oXsRF+d5FpL8A1Hb1HIwacjVskarA
H5y3IY25Tm8QIsldZp5NIg9uCieb2y4s+/ZyCIC8jGnVZV8mrcf2D9KC6/AF
DoWyTjZbaGytcF1nX4GqUfA3FrA5Gnv6t+exfGYmsFsbkPSAV3eC+qP3eOSg
wYlsxCWN8Gy8HMgC/azRulS869WaZYlOA+FaOzWYxStQ26MU5R5AdnMCYoTP
FGQ1/PEVkHrY7TJRldMau4WfjURiQC1GSydHrw61l7HwCmHvfkh7LQdnWkSf
fQ30OWrzKAw0GxBzfG9isSY9FafXm8CxF5OdL3wyHj35mYdymxSHkTN1a++a
BFF0gQZMhrz8S6OYhvsYyT8xfIrOl2G1UJASGlU7o8B6kAZDOwAiKp23GWyY
9zR6MmS68/4XWoYEOozVF3BC4NZblz+vt/5xHiXv3PF1waOMTOHmVQodOlKd
ZQ1hi7U1rSueM94BiO73RQQPiANWUcccjHStbNoY3SSPxbG3XoR72eL1BqNP
lMYwx4h7BPLDTy00tyRSZXuMMBEdFeBm1bCo7OBaC0yMdyGsqgS92EfeUKmh
aMt3UbTgsYD3HNIuLtjjh8EXVI+Y3Z08ez18FFpTPTk2hfJfXHC4pW6EOHR2
w02NN+2OV0w6PPdXDI4B1rdahVtQJqe/kjx7TyOUvY7p00wzkHHjrwpsnf9H
WiBd9tK1PlHztAiDN/lvD/aXjL4VCANuhZFHE/7Jh5TvwR+r8+/XKXekwla5
AawlaqrJHUcPRBHq4oEyU5i9RDjkvT5WdJTgajD24BJZd0yRNUqMqOEm9mR1
m0hM/9tRkrdEmtkPuTkaRx3/K8RfnI3yr0pPC848riHAdQ/IBPgGMeVBIJiH
EyiPrWNBub0hcUoTCqZYNmoR064l+GVDKhYABfOVJHbU3KE651daecmr9j89
NwJz/zFin77zv0LjPH5XQhyxfa1EqizMHtheCqp5A8nGf4o00JMu1t08nGeb
yEczY5Hbhi3gx/ajHES+G/Eawx8YiGIK57Ody1ttEaAVgLMAnx2YILKVpmuy
YTt2Hgjf6257wdIEDEpluQsFH4rZmzyveVuZKGDIcqGRK8tsWpNwCod79j7A
jk3mtadkIg2rZoqywAybRNOFXvZDJBwQEWib6H6S0gXZKzEYCFk7YB32O41u
M2cl1f2vuR7HGWcJv1XEyjZxBEUIH3aBe1tOIdMNeO2N/WXSkDsGLlAGYI85
gbhs8fe/QHlZhp3TisbeC+2yNIQGj1eZt9ZgrB6bjsfqdKNC6wqAX5f8fcwa
9zYbFaTTYx+QFz+chkna0p5blPXTDI2oV/iVi3/K7iCGoyZh3swJBlVSO1hY
DjtF9Uf0e6fZv6+muYIHUZFadSTC4NXKh6Cq5cmrFfDTXNKsCzy12vRAwdff
jq/tJoSEskyZLk2M0uyAZgFjMs6vot2tax/tC4yNRLXasJtbP5WdJSFa/CsK
wgtlA1Xi+EJBmlM5C79MsxEHK3fXbj74aHe3k3RRTCQ6yfIyzdAqakwQ8KR8
fK52muOfIw9aQQZYjgN0Z6UhiNKGII3S0sLTqOU62bezq6Sur2ecPkgGZIp4
qrnlxtDl/KoBkD9+km7Xjr1Y7StwNFpn3vRyThB1fDvoG3fTaJR4aF+T0olv
AZI1GJQu4cJgdfV4UQXtkRI0CqkHCZcavIoSKuR4CzYXIoF1ewmpEdJD3e0C
l6i6FLXiSgend/UzZhLPtKEGrEgPe3L/NH4NeLbqMDrNf5nsWmBImGUOBITe
X/cDL8B1DGJmHf7DATSSXMZ6o4+r2mG2SLp2kWuxq+cXfQnHYCjaz6PQBwcC
dDAepwuJqrkEG8cN6DM2I2rsdfcCKBNY2ccM4Rb9Po0l7oCEiKWfRYi3cmr7
sgugzTQo4v7P5VrlK1d8OO3T0dV92xtRtYvNH20D/NwtNhHEh4eh1qK5NIxc
Hg4l9bn+mbGv4nO15JBA3BZVgyJKcwgZyRz+Z7lNnNwiu2YsM+rD2c3Fez5t
VvZbI2SakaWsP+66EVybIhmxfU5i+zjwDoNeDa9gOawxf8IZ1Kyogd4OpF92
WKsDeiCg5WKMn514hvk719ir7ilmmNMfk+4oYPUkmkG7g+oepT++z/evlk3L
27FWJ7XFQmXx8qEb5abQWJcwaJ/SZq61ZNY+BhDw9YHUrdDhj8IR1mly2TMu
cFzCv3cL+9KdHWBwf7dQnw5EXuwhhNK5U8DpnFasLj5oGe5ubB0XvSlEeEtF
cGyJuN5kwRYtJJZe6vHmfE7yUHCqM9ts/e1kbvjd2ju0OhWl8Q+40PhiN572
DdxAQhdGQewy4/TaWwFjyHEZzk4zQwpqcT5XcBXwl9HZIT3kQN+hzQACpsTt
IoqTwt34Luo9DPWrkcgK/l2+RYdAGtpsb+8k0qbi84SbDtW7pDYDEHY7cx7b
KB/TD7QI7rrI3xrMK2s/3JJedscPtH0HLLt1/T8DvrWcCIha3e20OSiR/jKy
eC/2yxR0YwyG46cwywDUizHxmVBdf3H0dTzYDCXQsOGKxF9MswraPRLzU5Lq
nk5/pYlZDyYN7Q3rdKlloTJhPMxXlIGBJQBQHZjIuUcLKaCTIlxsrfxto5IL
mDgkD+KW3STfH0x0Cw9i1+fUwaxoVVVGusXKVT3I2+KHPIXcIToAKPAkQ85I
fh3pSyiVgseI3nb0/cE8XzHzCAC1cLvrMZA4pZ9eP1C9noz5ZdChavLHPsjZ
S8xmWxXMwrLPN1fVwA8mnCn6zEc2ukWuJpRDAA/XmoBOCGCmWb0EhraQP55E
A6QwC71O0jrJhDbinKtAj1yyvN8tFwMfOnJdXvEC8zOAdGe/cC8rTsKXd6+M
5dxLO8wLMb0MregHaxdPPOlddpA2e6d1rgjjzk98hx0kPI60vfbLr+k85Daa
TIFMY5xN4lYqQ6G4I4/HH3L+dgI/XKfPU68Irq1wL5VNwXguci49xZeZRtpK
Vb6FTvQEwfES6DiVQBoLSeWlII/DAesg90ivK/y/GFCzgjpe94VQ3wnLKwTQ
a+Gd8aiaqrmE9TmpLm+9qyR0C/d3NCNCh0Nh+QMgP6NxRGeY9D4z1iSSzvHr
HMslMetL76DvmAl5qxGBEMn9sievyQHa4Oe/wFyJDQOeP90Ibsk1tJGGsoX9
1goLa0yRaZbL/lZCZZpUPQ/mGYQYxM7MGadSvpTLXQFi1omnRF30XPkCvE6w
020N3hEaaM6/35AmlYKHpYPIA2gFkhwZ4KWaZ90af9I4lAju3bC1hs609tzA
2HlFaNbOx9Dj/r18R0XlD3t7o6G3qNb2+JR1aqoKBhW7C/x/fKFs2ninm7ql
NkUanFTERPEOGB4D7OSsCNj66lKKB2hjstk4VIOJHhaeMFuASpXxeg+7hj+1
pfzYhA13OvNLqimqwEPT08WbTEnmAdko3ibkNq2Hqw3ra/P9bhN/+wOLDmoW
jYhLcPpWl2fxKTl32eiqrK4yBYrIMHAXisF0Yk5VyoqGiRvIwfhXS83voAQk
yqVtcCfZvLOnMBlWwOPbTDnTeNuVujslnf/tUxoXxqtbnwu5dL71crj4DNdc
wld2l3IA7etViHwlN7yj2qhcAmC3rwrsU71TkzSIAEViiotzIS5GdPwKA/kM
xQel0Pa6ygvs6UBxCoC56Yt9uZxfHcMeTnKot8eGbwYeqIU9PsvS6UWz2YYq
x9o5nkbMO6KiMBxNqTqn24Z/qE+7gOpn2lCipdzq8CFmqLqc5EHLAqYsGCMf
BJAqycS8QnP684DbbaM0H6mSe/1PBb8IVDYrzPDoI0cpvZGvUrYwTG9j4b7H
1SOLl1cKChJSDwwzGAYd8UH4+A9FA4FmpTwDAVcduYw5rHFr8jOJmchnfk8Q
voNqBxTFaPYSDeoebkwyNbXTmkmwtn5gPOmCrU0OC1EF1FYBn5nhHejx/RU1
3CCQMh7TpgSrRpqsov0aAJ2Vde0FuUzxp8LTJ24Uon9keJeZAz0ERkw1hoFi
DG2bD9NWyPPdQ+i2c4F2b4DixpzmvLhKOW5dxgwt19RLGVldswW58P3+jEd6
o2F8NpnByugR9V8mfFd9zL7z1eX+2uTlTK1oXr1PG0mVnM9cnJ+QEnFpLcp9
YEakdhH6H/SBw7fa33cTf7jXaI8vy5Oma0CSwrPTscZFEClt0I1xMzplS/68
1duJT18oKBmPmUBF6GW/J8yvPoL6p9VbboYwMBuo4DcEPyBTbDqv5rEdj5Is
hImqftgKIXap5/IQMWqK/6TykX/TVEyr64qZ7Rfw9L/XBEGIJPy/oBOpFLEN
pHpfW6bdhkXjNQQaPwpoTK7KeAXRY1jCB/NleTJ3B6GYe7Rzm3p3LBU7STaZ
yYFXv6NPOmXCljXvhzGFEfH3zjTyFCqjxEZMCq02+23E+37XiIFzgd6ov1Op
oe4g9rjbhUkfdV05uKkp8q1K60cPT2cVwqIDZ6IIhDYUeIzPvEVdOFrNWEj3
OFKSMOxe3crpf8ArLFBCOABARih3QonYViWvZgjaU8690F1XkjNdWgvAyPa7
SvKvgBSGpLSPFQ/d++Y2FXxDX/8BAlQOWB89V7UJJG0sPNBTf7+hF6is5jkB
EnWv4mPt2TWqSe+nbQTH4LmiyJgHSHh1gFy6mwB+CWh05LYhuoblRt5VmXxQ
JmTIht6yws9ND+j0fGBi6QOsxFjJgJWDNVrsZkhGZ0sB7vp3ErzC/RkosvZA
cvdepv1UtZrqwvCm6xf41BIHn1Y8VSHKga0geRh1RDpt+2skZVDG5lwRRgD3
xJzVska6fmrM0X46w1jeLjBfzPmO2cbIL+GmLFe87yO8AFR9shNwsFhcYqUB
d/jB81pjg8h5yzWEgAqRz1FOww4cBnJ9UrisIPZwRXEQkOMTSHWwPJXst4NZ
/B4PVT+CpDgGQjXFLBCcHFYYsxSzNMknSCax/xwHBjuynq8VvkGzuEhuLtpc
vT+y3LZzlULTwod5HIr8tD+F6MbUa4U9PuePNnv5EkWNrI1JiGuHwdm5lqxQ
3xYyzZsF7FgDNRKx5sjKCdDaGkylPItgV+8DgL8+rxv8SEmHvj5t8E/qve6v
S/FNv/5jPCeSBsz89L+QQ41nYHSDyA+sBU8vY8kHT/x+nTqU/Yk+3PZIZPeI
lnh5m7wwtSqpwrkP487i6wrHWp8ITL5jQHjDZ4qjVtO9C6OerggyIEEfl1Y/
MxDiEjbHGofqGgGyes5sHWnfvnPAV8bD0OHcI7G7SrdEMlGuVUCAgXMLCj7I
d7CEY5Oj+7C0ir92szvqtkXoTikzqtD6x25vuUJeO9jC+ET6w7qZ/9bDeV9J
LMOvDB8PQW+basBr7sXMhG0Rn1YJdTJrUyMfdaR1S9QM3v4R5h7+q2V3tcCP
eTO2vfUula4xj3iN6OoJ3XoyLNjLb0+Iv6xQJrbXa3cwSuHa0lqM00eHrzSu
TiKlhR496ReH2zvTgGLgee/2etarsPd9cid7d4CPwXCtTwoMhKXV9TRcWQqt
RnY5PUJom/lhO2dJTDLHrls1k7C8fm8zoqT8G+47Z0ujYKbAnA0qAqfdTnFi
XWu6HxXSNywTNGAyqTtIXqbcc/enxDwCGQ6mJa0yaG+j3aQxZcJy82kWnDEy
DYOwbMP+0e20hrXtcrE+GOMJecTdXTGemJ5zsd544wGemtjaQxMPkIgHx7H3
jm/5lE5nc4ZPGUx5LjygE4fmhoRMcifMhKw7LepBl0U9HhGdZJ6xXPF9BGPT
/8lUOBG4N9Twd/uLKKtSEJE/plFEZW8cuP7RqOj1scwZiac8V6XXi5A806w5
JzRl+RPM12umGWuk3t5cX/t/lMmYqAVSqAIqWf4HY/KowMZJb53Bhf4BBN7w
o1vGOEckPOxnBSoopjpq8pkMtwD1pq8i/wDDLwXgjRgxaKX3OsCOSqqPJB3M
KgTUclADLO8TSoje9HQuI4oUKmrbgahECzqT5Ytn26RycnxzZv/6wMbRA+R0
xf0pnG0yYjGEB3eMW7aN3RAqKWJwLFmToDgslq8agkTitaMzSASMpGLolPm1
lowbADtlJ6tUiHUgr7eBNnfKZ8FL1Yuygj1AiVln+vv9/lFnGyI1MlFb7LZR
dkqt2JERYS0jOmkcFbhHTqtF2Y/F3VE6+rDKJybxS3e6ABE+e4+LMWofnjOK
0RXMd9Z2u/nudWWbHpQBU2rpKK9Ee2hio7jImtuQGVYbQ6pDYSSbAYNZop4b
T1+4xi0mEnw1SY2CDRnpDvNTrryxBUi5k4cPTe+RxSmJn3L+zpEGJwJAlBG7
wM7+JB6V1AKKnEiQskoVzK0c/0jRj0AkK+BNtRB8jRPLz0Qhq3PZnL7LbspJ
2Sg5AQ57Otz0BKK9wPDvy7+3mB7Cpy/liZIlHH7B0728QThTb1MJwWIa1A/e
C7AezkyqH5nrDHIlXeyYiiOoDb4lykFf998D+tboCnILjvxjbr5aeAcvtPJd
zsRDemEkWEmnG9RGsDoM5lEhD5reXupPU62veZxtjuHV+g3dEtwOcBEbXDlG
5fnbO4ZRG1AYyXRioYon1BitnRJkOiv57KurAZRtvnaUSHwt+BYKftGy0ogH
aAsdA1IH+BwnOCgbY0mhbfieLmR74qCF8HrGsdBQh0Novha0xxdM4qIucuf4
EdpKtAjOi7mqvjn69oSWvuP4TNzSm7cmc5HtKqQcBJCcylEljbi9N51fdgp7
tjxyKjALzbIENdT8CG08vjVGhF78zY8mbZiiF9vXXssDRoUKvSF0lFLLQ0tl
F+DFPFr/T2HXpF5pHtumolkoNbaGcxKo7BJvqA63VzlRmdyH93ZJtV0QKtZp
GlObqYAMeGou1Tm3VTmZa0K8q/tt56j6pybLGxmdIUsgjNvMeE6yCQ6Uxio9
g7RPvyTuTMWdYLLeSjKEC5NvJFpWFgqaZlWlsVC5+TqztI8xZTDSIjvGMoO/
2dhokQPXkWiaXtYwS1AyXTxtebTaDc0pL0DYuUTNjbE3qu3QNFG3/Gv/GpnT
F71dd6TskOtjT9iPsjoqATjjh6uIjNmZ5Faq5rGlYTJnRNq02wNMEwodJwdz
Wb2jDx3WyWZkbylHqd40Xh1HMBc9YngUxR5WkrQjxQiNiqVrkT0wlOozVs7M
9HWRRft+NFgR+629BeWHukveOpCEE2WzSUBN3uAoC3tuBDaRcXOgzf9OWKCk
IcdNqAgcwUnBSKcUI9a/aC88CMKyDkvNgpIq/arD6y5SEiZp7nST8zQFiPQo
KAZmRRV57RDLB3gksukLYLOoWFAXIGFyp0mwNix8VW3OGktHHULsfbOXc5lW
f91INHH79pxlsPQmV7lkNNc+ab96H2RPHLvteiG6KTBUzNyRu8Q7LF4Fi00e
QYjnsJ/fgPPW/YETIi12jPvIs+cAQlADyiiaWOHjpQHOa3hluDjc31beRPmL
UJiy0VMgK5cF+2XuK25x2nLxzfgeosNfN15Alja4akdq/kSJMJiiNo83vFM4
1F39ZTdDElJXRW07uVGfF0ym/SsY8heGqqrgjGqlEou0f+wCda5FfNv4CxY+
9ZuyiSTGvlJAp4DGMMOXFes6m21rw5Vy5fuZdOAk9SrFt2WtQluvtdrOt9O5
idmJW1Z0qCbdpgWD07M60B+f8oBOwxfekYyNHqNr/xOPuewjB0LB3TfvmSCR
rm7gPv/lsuOh64UadvJ+JsHxWGDSjMMdlzvpaBJ/591qGhJW8iBSpGPjQ7XA
3b8neeA+7OV3q4q1NkmYIkEc8Pm2Hf1Kxu4CCvJtHTGc4yUF20eR1UYNqg2N
niJZBnFbC2ZDCifhs+HdP2U8ON0a7/m6si2P6Id47lYEB9M3kNPFtamtrIfo
v7SEciXXvvr2jKvqeQ2rEmh7ONzDZIQnbo0cCoespmacn6T+GQ5GvTpDf8B9
WnuuNCNRM5jNhypmmli18vUhJHZmqqBJUxZH2p++c/MtZAqzftV3kuK+6vzC
qRlbLiGhGcuuhvauaMcdVpE4xVyz9LfLyIQFtrPOFlIeV31MgXjxCk37e13i
U0bpMP0s3CH239vnaEUZ2Ta9+YAka9Pl70BbCg1UByuv5lA1SoIslQlfGh/F
I+DoDZczOPMIq8DhbY4ca+qwGoO1KNrmRb0rpi/ylKAzIti42JnA9PW2R04D
fCvb+MwczcxSB8rSNwH7FnwMFkt3RsvQ+eDM0xFvWSbdYCmGxx+WyPQuwvCh
oAZriT6dvAZtugtahGGomieO2FqV0Ewl+SKTn991yt/pmbPchV179F+cTPm+
bYUQqoHYkAFOt7k+6+k90JaN36d2kDwX+/kHQYcVaEGbgw0ZYE0cTO4S7CQJ
Ty8qllKf3h+Zsjvi/h9I9j6bcgCv6qKmBbYnl79cM5rzM0fifL0XWJdZ5p3C
CybSaxq6uhwByoBynRvOaRS9dQfe22oVU5s64gXZprH6VX+pNoXOdN4KPx3m
kxi5gzpap3yqijZLyai6Ej1vEoM1Pq0IrOkPWYVAPY7letG3E/oJ4P8RNnXQ
KGKOSXt3I8Jqx8+AxIPcIBroyuV21pewWqsV5k//vRk1Byd2LzPR0WoKVNOa
cV+juC8q36/N7OpNk8B1Bo23bHMon1pBVZjLI8hr+OsL7AdhhDcnv5a0wmRK
DP9TpNI+ZP780Zw6PkX8oCWragIU4YAnVIjcvceR8loKUb0YsKh8jg2uJOm5
8uIjUwQrm/aah6rijBQj6OSDZIYsroRnzvFuLyOGa+SmFGnPvLtn8gSqgHHS
lYlH1SXgo0BQnBs4EMjQkDtY/mXmWHIVu7kVpcPOSHbvRia+8I0OKVDlAQNz
WNueLw/2GQyrAyU1lvSsNx/nMGGAigSfCbU5P3A/dKSPWjQf/cA9k+I+M2s7
zr6706agd28Hn7ir/K+JtMnO9J8LkGmbhzUNvG93p42HQA+MktZp0ErBBI8F
lUArGHMA4LjbfY0vek0WPFFlnJ1Y0Nx5UCf3ZNHhLYMSvJtInnaqN5+/smi0
E8J3vP35MUBQNiaNP8a2RmR2JjU13q+plZCvEuYSvE4Fkl37ENyWLm6+ZKTX
82kx1J/vGerxfvomcM8+aLF2/cGHIuvQyXFdAJfrwigEuzdoepNQbyDdCoGg
wr85IHB4T0IutD2SjyclEHtfXUwhKDL4t/V7RlhUx7V9W7vrg3PLqdyPBeSz
2kHtAt0IJ9EzSLfYeEuxljKvmU94CTYBLiOz8LaehRYt9f0D7wKNPwIxplRe
Q3pSMppJgWq3L1Xi4OWzrx5+35bW/H3rpVRTtfmkwH2Vgju7S6vSKDhrZ/8D
SZPaFmYTLvgyUcoTjuKwEoycGOZny/2VOA2D++Y6zRYq9ky3Sq4yuXRL67Cp
Eyk0lkaT6DOiYgRRmZzibRyChACC2BmM+36E+GYuYSPIRJ0r9XBokczFMzmI
DcOrlEOVuuxe5v9VQ2463kG2mJDVi/CvoHIuHavlFLmSh3beY13aBsgm6eTk
plgX2T8CE211StWCN26bmhq1WWNyo272NcN4w/F7HgtWo1R54p4jHu4fYyvA
Ri3fIQwj1lFY7ynweYkN7al9M4CPSHQiDs0OG19zBw2KO+QjK+WICBzAaFDh
muE2TZdh1bQHT/nfPgiht9AorX82FaHNFxg3o0znE+Ma7NouFNuG4eAg1hiT
H0lJ1WzxtcPQA5ukZDIfKsAHAqmIxZjpbJsDkD9SXH4I09wOfpcKQG5zaxxO
avpfcGa/tYKKywU3+qoNNjflvTFfuVf448O//IWlUQdDUK9Niq4a3MztuGw2
PTb24O6tJSwytQUkIFCNlIrqZdc3PZcWadN9ls4kuqmFMwQNtQShLY/DfeYo
m+vO8IetDl+PgsGk0LPkUNqY7t8w7pNTuRS/RzdIJGAV3hQR6sKZvwLEnfW3
QnXr7bX7IByMGY/H1XVWcqfb4ltPfv79iUweaIbeW1Oje62H8Yvvghr5Mcwu
y+uGktea7AlUZg3IalTs9RrusEyUSPp+v+PyPveo043KIl7syB2oS5OG3b92
N0guhHIcc4ANstvknaGqpvmGb8TPpPM9E/l0+tiaTiLeC/WFxIXrC0ph3OV+
f5Q26Gro9r/Gw1WBqyxgHSqDfa53sKs1PJQjtf7mLKglDeEom5/v8vsNdxFA
qaDu7FmYu6RqW7kyDAA1dLG0UZD8Xu9zzOzk0ApSIcZKG1BDvpx3vFFJFj5y
bOmQ3JgwDwLaQ6JYC0ivIiR9xRcZmhum8RqtqKzuEyRUcHbkJD7ZJlgWGLi4
wUg6V0PNNQL2Fl8L/YwRviCB6MCj0AUcqk1ncq7Bh4BHGRo/HPHDhNYIf5Bg
DWhjS9qFZ/iCDw0Uy+JXmWqusq3rpDQOrYOhPt+5mTk8nZCPDkAF1Cu3NDjV
GxWUbdLN2gkIu5N1ljloSzjtjC6i4baGHrAyqsX/OuMdTY7h+PER1rhwztSq
4kTQ5Li2b7gYYBlEsM3f/0PUD+2CUcX7FYNwJEkggLA20bjiKVOSZEMbDxiG
6SWY/w+VTrjY6D95zQio91Nxpx37hvzLd67X0NF1Xv4h/WuqCAdsPKee5/ej
W6E9z1iIqKAUgE8LHVlTwtttlbKTiXvYIUwW4+yBamgSxy55uq3H1C3SfJeW
gQhaXXaNvqjgYNoK2XRsrnIPxRVZpXql7E/BnxDXNoF2NJH/b5shGN49I7Bm
tdmgSRC/I6ebaZi9npfgwaxaPWOLOC8/jF1ot8VJm67LdvF0mxYPhQg1tkBz
pbPBbGd0pG99BQYUCckdDkXS4G/i18ob6oAg+8QquXcus6Iv8y2yfvwMAJY4
8EaeYjz1/VPbDjUNZyDb5xMgiE/mGRA50UpITKxsdAf8RGStt6sv7HjVNDmv
pcxD6sBlt6AxWnpL+nYwXZPZ3Hmkkyk7MbKEknf5b6EPdE9GunoL8mwgfgns
5L+yfvduhXYRWJNPGSznpTqRVv/Rm7b6n4t0m3qFclgaSm8WWGS6cxKNet8U
MWx5Bex1M9/Ba6jA7OJ2TyijaEy0cmyD/aB7LXo8Yj+4nuc3+vWkqdrpb3zX
GMHORzMgyPaZw1WvE+wciEjpGn85zPlG2h43mPWpzglrP5x3HGLKkBxdI5Ez
hsSC/ZDTjYBqy5NGLjh/RkLZrSghiZws3Fjvlc9wxPslWLQ6V7NR1jvCKCvx
rRq/PrDRFRWI25VICysmZSsU6C30/pMMsSbhFjbMjRTNQWObH8y+9cOpVfT8
QdkgckbnVekP00EZjfSMa5MuE/qpwOa7U0AOR9LR+oyIb7Svqe0TzuqbDO1R
xt8xD7uS/AcNukR3IKWsrwPTK9kQhmtqVY+5Y660fDP4/pewZk5KlSXV952t
wwnkhUD0qA536oCg7WAXw/5vZZL3JUrMg2Apd/4oNYXlMrj868LiJOjH0pHz
qHijGn9Ue4FxdID2y2eJ4NEDRO3Tra+z5tsK5pOn7jlJetgZg6Cu6GDL64SM
A83hMCA/96UuMb6IlGsQDgwQ/C8FSKelq0HrqfYAVuM7GzpY7EyvWfJ4q/l/
tV8bbVvJt1YNdbLRtWjA8oTSB/OXxOxs6gnc5wPnh0W4t9qZBjKqlnxl7rNT
j3wp/RtmnfmtVY1pcwNs7g1/wyCDEp1aKaOXMldOpG9dhTB0BwXhDVEhI6W+
6MQpF+417teAsYjesEcnH4PYYmH3UjASwbVZl4R1B6/kShS48lda6wUaUoX2
CJPw0P+QsPCz6kuOTKWEGSV75URoupxMmcGC7W9Up8vQLc04wDjDkKoW0roe
oTuYDGR2ArgUaymWVkmHA8GZ6ZNWkb0xd60jrn+Qo5y0Rjr6VmHt0J88uh2D
WaqHCCyJW/ZMPFXUCRq66O+tMIJhPyDXbvoZVhqUSfmHCbEf1CfsFYSMMcoA
qbNhejTwh4bqw9cJOKb/eGaci9auDP3DaaxM8xTzFrZaJ0P9Kg49w6dSkjkB
GcJdKbZMX+9+UXtfXUQZHXNC8ri/rNb68aqB5ENxvDHsQv5aymMYeqAYi2YF
ihLz2egVT1PAnb8gMZ2Cn6a3+MkU7i6nt94gsbnrnNRbm1F4dibjWYAPreDN
xamqN5ywSr3W5NAi7vMGf0d2Do8BwfBiL10jACNX0YfsFNP+4eLRegGaVesi
yG3Ae5kWnpYpdxUQK43Ie8bSY/OytgTFY93kCYHd7m8cQIAO3QdBTwQfNQ7d
hKeaJNmsPoXDEo51OUbFK8tOt657jozg8JPWyxarl2nfL/qwt66OPzFDpt/n
/+xm8aEUwsv1CyXGkyrQVSpgr+Dx/LidBDYy3BfNkZSWbqKS0YW3vQ22dur1
6sxLDND50eIV2pRrzE0qoJy7ws9pzM3C1w6EHreAoJjwltqzRb1PNQNaBXwO
wKhrzQoJ+1MSbb9g+AYS4ccAstK/QEyO1UDPSQA2Dyjym7wt/QDQH4cop8vU
lqObOkFt/CFmflqC/H8hG0Ylwqfa7KE4VU3jtJjM37W7qQRpdYMY2J19hXcM
vqIv00e2IGTysUY2QuQ1YVT318l4LVBifwEpFQHwu2CRAWW+C5IKxZyLTyFb
CCsh+KLclSAWxez/QqQEaJNQGTr+fulfS7c7PeXvzWhBKQDUXIeAlK2wYB7Z
DLTGGok6va4NC+/JEdZc/IZH8gFMvQ04c95TBMxh9Gsxsejv31wLsX7msWSW
HlqXr5XYn/Ud9+6efgWOG6UjeMEjfJ5Pwak/8Pi9XR2qDCGfa8TZJHVHvcvt
rncpHryyr7QtLu64+4Mrex//QHwDvl0j1M/Bdoy03nFTjmv0qWWhoawxsKux
mmDrrB0e3a8YhcqOzh533sdwxbj3jl/OkB/AUsFBEwW3aQrY/2fMLvDnYlBK
dKHoYZaLp/afDy/YlNkAUZvsvsSDDlASvg1iL9XrY4lzbjXTOG3rrbuP26+B
lBBCPGBfOv1xPBSDZfH3tMLQq1DNPLVTmfRFfUVGc4L/euVqQB191vYsrw6S
+DwSEVd1u4kdy0tb1sQ7uy3U5C7x9p3plzKMVZmYcSD6mMw+QJ4LJHFhAbz6
9zHFxk/DDGumZkYMdAxBAdPy0ySt5aP91ejbjVxBtD78xiREYqMCiw9kvjdr
07gXHJeVZOG8aIFhsriReAAKbFFkPxgKBq0o53YOYUPe5GI3zS16suZXQMcf
P0v57VTUXUlbGbtFPQhH9i7uWCt00ynR926z1vSqecNuXNd6TImDgS7gz1On
HDFaDfiujSCrblNgs7DjR+3o+6xKRsDhmSKt52inKksqEhl8lsXjPesMQzsJ
+F48cv8lAQzevDXJ9rjbWvApevit9IKhkCFWVOF0t8DmXvXzDWnVh0MJsQhR
YunjExa+FOlRRRLt7wL+2RCAau9xf3Jo6vqQmlMNRjmi0fhKJcKURTK2mMU7
dv5NSaOznMCEvhdurhlRqcbrMGZR9CUVMljTTAwEdc9BxdVtcszTBgJsquvn
im+EFzjbV1/z4tjuMBae1gH/z11gNV/i8l9Qxogho52l9loXjOdDAWs0rrso
EoplrSHdLIC23o5d3NJD75G5yZf/189CqwngBbp1jH7OeO1wsPtdnvbHbkvk
5woLiVoqaQHEsFBmvmihc1uA6mpz/VjWizcYz+JIW+GtG4zw2xED2XceRAoF
MODY8J/0Mv7seswmy+o774VJX4Kx6VmKQhWmgWP0x1DtPaA47H2Elgbwehb+
rwkWjzQQD5OxvPc5ahue5/vzUhpMqgU6SST/11wCShzXzUg2jncoBbwy+V8i
WSt/1lbAp72mOXIfxSHNO/ogZcUCGyasmO2WShEDcj7wHBJwWUdV78x2zj0b
28voJtnDAAWFazbJFZLWESZOqXvNZwvjjW9fbmNFv+iB/yy8Rga4s8qh4yb1
ZFA9/ciOjpTd2RPOrxCdpahf2hfrOnmqinqsA53YMN1XuOnD1/IgKDNSPD0/
oOaOhEaScF2W93OwHv6tNXvOftIC34HmRUIMnG1qlSnRLzMgDYuNi/BE29G7
MZwt+Fzsx/tuewknr8KJbqmi4X0cln25MnAcQK1ZxpxKoTJ3EKwLwedQv8Vc
hfnEVWHxO9HTfExxaO5sJ0CBl0gIxzBwoGKR6ARCK2R+iK7nZ7FL/jUW6Zoj
aLwJBEyGd2E1Fh28CydKn6xSJv+Ei0g0WwAd2lGKfdnRa8321bJLAhmbuqW8
nNj6Q6YrwQD0KSO1nqRZI8ef7Hvkd3WoqeeP2oV6toGuBhsYw0weB4MZjcpp
n6gI6dDnGgphOocXRSvNVA+t0vVRXV4ycmtMU5M1j+J7F6S4wT2MRCUEzO0t
xlZGO3EfN+a1w+0Fgm+pNauiYE3oM+VMihntmM0PJ+rX8XZ6pE/LVhm/mqdO
lXj3tyOWy6riCHmnfgjT2HScnm9iyADfqTOAMKoHmhQRNbd7cJ4g+Kg9c1Hr
NRETyFLB/CXmja+CKsxgJ2YhDKTXlDGxhG4KpbjDPvdbjmU2UyfL0rgKmtD0
HMXZ8I4/T/fPDXpcQE0YQsBjokToDdU9UgTo3JlRYVdFzV+R1QYSNfL3ZlVo
ProyHZB//f8/Q7qL01w72l7ixjFHVWFKsvkh04ASEPtP3pn4oneqtUmW8EyD
RCQfdP5YVer8plvAuRPGUz97rk4Lnj+5ym0sgn9jxGmE808gpZAoeUtuvVDL
S/4K5D8KjmlvxxWm6w1BGOM3j0S5yomnCxNBYozAbNU/pvw7MQjMCKLNc880
PJbC6s7SwHP7jAaAnL+kh/lJYAZMPjyeEyozeiRpbNdsuE3wM6XZQ+n3HM2u
BwRYlP9+biBy3y7vDK5qOSfg58oPhWlRaA3/AMcBFh6EfD4MxkOyaD3u8LZz
QT+yrnKv5irkAj0Ukq+B63SHswrWTmdFYmCZReHPXz+cv12eiB2B1G6WCLh3
eKDqUjkcXvMoxsFxzXbrP/GF8HlGrbH3u3v/8wWnnfYNE/cIb/noPY4YzrwO
SBOcxjrcFgszyt5iS3nqJwop2U4ExDxiC3LHlUP7FykhHoD2IqkUCYdp94Jm
GaOBMQpWP4kCvu3qXo6het++lV2Hi7sVEHjIOLvMINdRtjl9vyjxmVLMQ4g1
KfG1t70H7DMxLL2dAf4wqjrhZwMVNlrIa4c+9V59x6dOB5SMCAFVklxAw8B5
Z8ZpJIq+39TdKtqjn725G6S+YfC3HIQmdUwx+VBuAaK0vdq7Rt43Mo1y/DqB
ASx03j4v0xpsJzGOvvjLzPyGIpeRXnE17y/5fuV34bhOlLpnHYC6JUylAoKw
WVGEalkuEfeQ1ZeSVK+B22dmH4bJm01qI+xa3sVQ6TtMhc1AzQqZU/pqGsjI
1ZZEaZbfVLhJ0S7VisUpUQAv2rcPHEW1/y1xNaefr48b9jkbb2Vbs9JncI6j
1wraDIDYuDi69bRCByWtJ0dY+eWAMSE8Kd6lh9EZMBZuI0CZpiJ4OVKKEn1t
LeR4AnKr2unSeQIzfj1z3vn6D+wmhqJba8I2/21yyzFEwkEhyiGB7x8JTB1U
Zg1+dpC0wfx3pxW0raKr+rQSdj19+TluT6bsZHMEulIANLJNQ2ZRtVj9IDgR
EPL9CR1ypDeWepz1yWYMPBudxl7LPtBbsEqrfsissuWV43x1H8WWLtjut9EL
DOIRqhx6Ur2xCufhgbqsMerQcbWpLJ+1AXSw4x0Dg3R17mnsUO7j62ATwESk
sAxZy86Q5doESpF6M8C5jzkHUIPDE5MwSNXfY4/oH7Cd87XTCFACHGDwcMMQ
D2z7qlEn+7dom8n6Bra1jLSi7bWua8sP0Hp+JGok1iOQxVnMKNJUPnK1tlwz
0ExBKDUpgsRCJYcq6+9rnvgxsCMlnury9R310diQl8OV2FqDHRoSr4398X68
ybmViQF9/3iFJfy7NAt3loYvL6Z50d1unqvC4pUp/2mWKfDauZ7xtlsJh5Uc
Y1Vs1kfTR58TyCh6lsz1aeGzqqS0flk2hmN4vhZgsEJz4xPYbHx0KW8E0Zw/
QcsU85ViX6yQg3SpAzU9Zt64OwzWNBCbtiJNgWX5n0k/Gf613teMFRQ94Q8r
YlR3P1J7J7R8pneaV8t2doGeXUSLoCe4VvEtyRl6kydLvK/2fPDE7hNKdZqn
9Z9eAJj22/+mvfXElgz59plUxx4/NGokQBcCg2II6dnZkQ7P0UMQs2ClIkkd
nzmQVIjN/UE+k04Jc+9qwTm6tcHKUnKQN0PP+6skEmUgab/YOKdNFRl5oqi/
vfTQA+tSaRZOPM/2wsmUhsJz7mEsVFk9xisyvzO4rwEGay/p481anSEZMrJN
vPeyMWNt0jNL8oS87M/MILFWQkctdC7aQRI/I67c1bc9MgSxnOqEfUaKp8dI
YqsFr3bfmnmWEYTBzuNQC8Vrh+FrN52qW4xteGinkxuwcsOZyZVPyD+pFRTW
zCRx4KBqGbWQpN7FikTcg2cf2Wr9LoAyA0X36jReX5Z2jo6RFDVCaqp7MZxa
/12XR4v7sbU3VQhrJU4FixfNWa7nqAYVmT1iujLb2reCMN7jYQ0lSsYrkU/+
ZgTGwsFIuP9pcgvT5ToVmOuihak2xJ6cCDYTcmFr8a11wRm1R5gwK8wkMQJC
Vhzm5wPHTysgaZDgJ4HS96/dv1E6kOLKJSi6y3Mrh7Fx46OwsfBALZu0Q4jF
qnpCXZmTMGJCpwJC4UvBVo1vF4opSPzl7I3Kga7rmVLn8gHvOWef72MA0XLI
3aVNyDUGDURyH1V5kJXEJQxbjjg/YjN4nEzRHLLkvTYkXZC/urJilzs4SEa+
O/3sKRZWcozPyhNSwSHJ91Y5ZcCEqd8VFU4qETqzY+ja4xrSTalCRuP8HoPN
OLBmQQU8xYT/LUOzXmjplapCdkgf+0QazqJDRiF1kfjZWutDizVj5+iRLMix
KIQ11IdLvOMhJUgvgdahofA0nCwGLXe0kIICWKjdtwTDZ8GgUkiBNsGP75ZE
6X4TmjlOqyhjJAoRLM+cQkN7wdKefdR/WgHD1OdhFa7DRwOwU1oWWk0+NJor
h9lzFNs2yqUP5Ugitr7jXRoolP7f7CFI99n+xHj+wfzye2nEyAXVBuM9syTZ
kXcHPvULiSyj+c+Vs/R+NhOyZWTsyTkpFp4QYU4uaofSUFXXxoxvFCTQg+5+
Fx2p7TFBpR8sTPdJgj2y/szxPBk9lSn41WpkEc9fvHJCl41HeQBO+3MGEk8K
5otmX3zESo92oP9S8/tLh0+b/VzV2nA7DoiPKZWCkiCPxbFx5yKr6E54r0Me
JlXO4t9SxeepENGhpX8N8L+0AixI3ecllX3BR+prkzSvlZQcdnqTlOsXVqup
T1OWGU3ukXLhUTtJ0SWE6KbO8rFGSE6ys3UF74u2kfR6u0BoUC9IR+dPAKBR
4ULjRM0p2OaG3bLVnHenMjgEXN4aaqJ/RIiNk14RCQoqpr4ATeuyg3Ls20h9
woUd38Lb+OQ69hu4IC/HizlcuvmNtrs4ITVd6Hfgf+uddTe8ZcGjvlSBmGMQ
z/31DEPy0+vraCR2q1EYnv3i9xUrLoU3Kit4vPL2UnuD5TmzMxFC8EAN08ip
5XhfHCvLrV0r2hzKHhlIb0xAFz11wYbmk0BGe3kP8xj2q3UvV3xPC6cxnEp4
o2MwzPg54B7XzSnbl2l9MwqK8ihdNsiDEw4tYQCpnuxGdmaAREDeov+2Ht7Y
bwLM+bJLwo7mT3b9XHEx1alAOf4/K4btrh+0RTiGUmy+dQckMpRxi+B7cuZA
/FhgjsnDrldyto7J/GY+lX6Gl9Kzc4a5FexLIVXkMDs774stY1NPWKsBSlxY
bruCFbAetZK8zxZlykgS1c2mXUKgEU+u+9Q1PELe4BEzeqzsWbujZ0mMx0OJ
WdocSz5hN5AAJIAzfgVrqWgMHoppD/M3WFgczSHKAapmmgv0ekUcgUSL/jDo
SU+ajoqA4nAS7k4DPV6Kxykzec1P7ZRfoJYROlcTW5gP1G+p8ISFjsQuiPP0
qJ6V4YU4Q0XEM8dkRsO/GQJIOldvXvj/Kg1R7xoyqxQXid+vT8bYCIg8jb6N
cjnPDN/29HnzaXsWm2lJTnWK2l5cc/yNUjp/sXr1dvdiWYmVU1VTEptA1EGJ
3T3gTZOE/1Xh6yZGev1PGRG1+UjYq0hx/Upvh4R51BnN/vS0ucNhKwmDuBzJ
jtMnauoH/7UkjZQBFM6UID6P68fBc4l2TCr32nZTAjOVHv9z/dLl0rA0/zGo
4w+T2n8kvUiV4i6ZSWvQZjzTA6m6/HcG6dx2VpZcmmMhGeygxgo5Iy6t2CuN
qiblPFtoGdAQ5Zw9MHN1RFrR6LpAKMoehFbiQweAhcm01tbEgEd+mU6SJIWS
VKxVKmu92QnC3aAbs6/tSWWQG/SX1BbWIjPgeyiDMuXM8cT6K3uwCUn/qNf/
VvrDWDYfuQfQFAae4GFwUBCwBARR2uiqjhcsGy14UACY9FAFJ0dpyXje2Cs+
9Fh3/yA+QlTnZRMfjOv0COXV/xKyGW9po+51u6wKkK74A329OoJAk+NxmDpw
hY0POoEoafMY38wMjwOfe6BN2xOnJDaCG3EYSW3bJaY6bYCtGy50tX7vqEkw
kQw2uYEnP6kjbyLlPAW0QZuWk/jwE7Vyvg/V3CdHydUS4Fs/1vL73xSaUOlb
gGRxk3ERGHc9cvwhaJAmr/XurvhxtjuxdtSF1RG/AUjTNN8k8LA+64I/MBwA
N9bF5tvAB7Yp9q6RIyujAAXFuP8dMf/a0w7j0IEnG4zvpUda1iPVPQXmL1LI
PY8pfGnPoiYL9+aboc+SQEPFeqwayADHx67l3MoCPKhcEmObNTE+rZs1cXaf
gsDlF/Osz8qvUJwxdVF88n2TJfjmyqbNNoxmL3VgcMHh47hgjk3h980zCcaa
5fwM4beMKgjAJ2/Ax+xpfem+jeM187fJMcnRgiVtWgaKRstsUHlFya5viro5
1OgjJ4QfZv/lp/D1AcreJh9hI3k8JaQDh6UElaJ5oUQaPQFYbE/oxNsctDly
1VB4vHphTSgOHfC0t/+1ahqvfrY5Xg+gfYOYhdDZ7DbD+ho548xRg9ISg6Oa
65NWy9GrF3K57YKN2BH4giQO4XWcWITCxFp13laugIiX0fWfDw8+JGtKNagz
N9x9R9a0fH2EgamlcYYUIbLsxxSn+AOpS9vOvAsP71Q6gYH4rkvfoF8B0ZC1
pcBnfC4jcG6UANgttD87jCFP1HoKNOgbEU+aIxbiW4sAeczLRxKOTWs05QaK
uakhepAP09VUnffwzNoq5pwdb4L/dkYCOiD9BzSNCj56iu2xCsF0iWojcFxP
tMO1CSe4NMKRVLb7kKa0TSpuEVauiTgVb25pNrMWJdSmX3W/GMPd+dfqgi+5
51i5WopTWJKZeVHEm2fhfbTVZyqJOGkTgoHz6a5TQtXgbJ6j1IeN+keCT5dJ
DZ+JKGlwZ8W0WcJCoWGlYsvLaYKpfjrN8erxiIlOO/dwswEgs9rUkPh1H4bJ
DhNh01ZNpHPFtYDG5JmP1JC0KY2/4Y3kEq7UJ+qOhQ0puMoA7Rd0JoO0jsrT
MLI57rRDgifcw6YK9D0JOanq+FOaTol3JsftTLAO7APVv2ajTAS/LZgyvfw7
poOhifY+LkwxcI3DGQ16rux+HekJC9Ihj0XFn3SqLzxv8yMWwq3733U+GKaf
MFQ1FBjBCS7bL06vkIcUXwxE0e2XrfP4A7Q7wyEQ55yPNKiCp94Urc6yM8Kf
tmJ9KNotsgqqvcD9DE+tPYTe+ja/qKMT1ZCX5xexIlindyPDgtgCBIB/PqIF
uP4lxX8Hd6hCYh5sCMTjUM42DBLjKQXEr+vCqWMgS+CS5D51zslcmJmttwyD
W0ZPbtopgyCREOUFV3gDkiJUsN2/zqP9j8vmsar03HPwLqzjws2DU8aNznCw
pANF1ni42V+DX3tw/Ocr1z9tdSZJN2KYVUJ10fKmkTrRaz0Hp237qhVLTqTl
0zr3AgZf7PWqw1LfFNd54vU+tW7iB4GrwTQXbsyUtCH8tu3aBfhZ5juxdXAf
B+MCk3M1iiJR7ofMPoNj1+U7ik8Ftg9I8cwU6Xgu54tf8VjON4niwtlkteUB
6ScsjwNlF2ab1QVPEW7rsRR+fLvFnsx/ysJUvXW6XbPxdSNna2w3v9zmeMMQ
wESPuxKjyaGpvs11RcAv1ckie3Phyweq4hredJa2muFqaLpdLvU5IMJKaQfa
mPJ9PZgI3Ryga8QfbOecKoz74Z5+wQpJTlmlDiIWdDVIQLy1dMWEtPjLOGN/
s5tBnE3gZgrOKxXpzXmEW+od9sB28lxTkwpleG6PnceF8ZakXmbZ6KD5LnFy
TemLB11rggs1xLNRoBxZnZuc5/fYewBCDv+XDvA8p6/DquQ14GEV8R9YikUH
YLrtU5SApkhWsLI6wmhyrCvY2MCfLA2tjAWOvlU6kY9J8FKuo0OYB4n8z59a
tMu6LbxvHERJmgl28qy879OzGO6joUb+epbrzrdHKF9xTkSCaOWkpdp736be
iKsdMij/jzGGwmi5s+9Dy7Bv4BCyKs1DrJC4+FYMvTnAS6I7nQgcTZO3bKb0
ICNGHxe8uKsmr/AUQMPgArdWqvjZqj7ec4xrPVHSwfc+c/V7WMG1Y9Swons8
2pRd2lYUF3Bu0xG1HCY970Bp7BNnl72blD6c+fxQDJyXg+6xwP3oKMRqCy+0
0VdKMadQnEJHM9e50LYjnGkK/hDGmDaRfAfh4EimfA4kOvWVkhVIpz1wQhUs
zazYZABpsTHLEoVuarfMwjj88PTciZ/7RFzO/d00PhxRt8dPuMpg+0IJ/0dy
nL6oYc1h8ud1D7PjHx6zti0wE55caQ911PqNK1ErwLBi2B/vXQa7xowMovuo
HxzCXWwJK8Xeci9584W4qm6fQIzor5jYCbK7ke3fMOZOEgnN9hT2+Y4iCxlx
XjGpLKI2akXgDcEowmJd+/VH9RlfKlsjw5undEpGckb6/hH3yXN+GOBrS4Xk
vzFYSOlnjRX5Edjtq0+8H83B34kWq3MWeuHSYbJxteocnV45Fi5wYI1AkCqf
psg02NhP47KwJhgPBnw7ktw299ETQMoQrbh+z24uQrqUg3hAPuY4+9mjJEhC
9fNe7z2OyOt3airrCcWsZUjd++9XyFw6HLXfKgIvnhmJ5hJn9d1mLVBDU9IA
PTYeTpdv8dFvtwQ0f7hHWdkEjQGiyOk8hkveP3X6NM4iyUvyuPpsmcY1gLZ9
SCBpKjkHu89MB3D0G55JzTMXg8kL3L1b0p+DQrvC5OTqkYPCpU3m/EZZ5+ul
+Y3rab1VQ6z8TXZEixQwGbAW0OBz5dbt5NEO37cnbonWP7VILT4YN/eLqYb1
Jh4Ld5vK2ZBbSy0K25Yu/u9anWhN+ijDuaLwqYnoka/bKYM40Mshniuz58Q8
EGDM3B9+Lff9KqT33BiaAhlTmW4GNcfuvjfRNC5Ea42LjeBi1EQxI0Pq0LAF
6KjMKHPuGLWH/tQj0MvafS8NQHqtg4h0bLYxbn55AT5Iqz0tYUeuuTtC2bI9
DhD2DcvGMULY/TQNNOnlIBeAwmxwXysTo8E+QmOsmb33YE5EO1fgcgsXOIGO
uto9ratTmTx8iOKau1gspk9mextwYDavZWXLqeLJc+gtL1KdtPbWbXyZ+1HB
PCGfpJkYo8QurTqSg/Oe8foZCn4UE5blEXX2jr6qsakxd5Bh2vtAKydBFTLF
FfOBAhIzkF3n5Rq3hD7HmLB58iPyL193qtFEBaVBrH/8pBbqPkxRrieSQ5xL
rCazX7hAawZbWni+vclJdA4+7EVSV0pIADmNBBCYezK//DY58zLoby4RK3wK
ck85It43NPpgTu46MyfX6Yq7ECu++AQCHF2buhlscIOoRqJ9fsjDUJylCO4v
17W6bry68NI63AaLbbGD/nQNuiGHJqNoJyIIPkT+j2XxrNQAm5XV1tIRRdRM
BbqVLpGW50LicYGdf3mE0ZWTjLeUMPo9GY2X3f6lR05p0w/4kiKCfUwld1ON
oeAU/6J6V8ZERuvYMwgKt/oRhwUh49rS+ywupbL9oCawTv9Wb4KoVU/zBmSV
R8HDZm0D4Cy9RCC1Z6pZoreDKYpM5wpAU55PZ9g6SJUfCsL+kec7tKHVI/qx
RLaWKdGH87uLSmR8qQ5pq7o+TYx/IbdWp7EjbR82Zdv+tHSu/RhI2ixa3uR3
GPhRSdaV8bOvkrm+CmLlmBMamNFWSqcYE4KHnbQj89oKZRkj/xCw7tAU2k/a
brP7y2aDIznWw03l+pxUDPJcrDZhOgHBIcHMu1J326iCwgtdBpEzf9q/vPek
fboH24winIG5Np19+OOUyjVIycl7f+Mr6cSCZFyIH2O8JFKib8fMGWdqwmtW
feLooA7VL1Fv4wvExG9oqu9AP3WUah1YFDYBGuD6CLkiKiKm1FAsBIKTGxvI
srNY/r1oOAFyxUw6gnk4wSxwDm0niW+4Wj/vhitQWIsdQzka3LZu9PXj3WhD
gssLS2rt4vGJt32pylIR7hPghqkT2pTlr7mQmiHQFj5Pz0Xb4cYEIg/yMOPF
8yHw/lKAVZP6h2P4xuKPRUFkReYKv9CXntZ4/3VPS67B9jX2B49Jf6YUOWPw
ygaTcYld1S+/x3cf7aSD78ToqHIsrlJB/5vgsSBP3mRYLwvmxe+6BNPt3QOQ
gPoPktXh2dkvQLfbN3qxFC+yx1GH+zswdtrfo8ubOysMPafQGaKb76PyXi1t
22cKsZCLseaGS6jIJ8dZuae9jtefwCJ007Yd3+NBYTM111Lm/gpDeHwRRUUf
pr30zuyG7SmJCUalm0bh9a3GobTtuOgMiqDfaWGgZ6T/c4XovxqOprvKgInk
87j+dCRCuJObCW1Ey32P5Hn6+GG83ugYhMp+7702QXYtfXq/wIMVhTAPlE9+
Hq9ZCAzvT0vtRCBLpCxl6/ZIxtA0oo07qsZ4RZXOb7MVbHeNuiX7z3mAby4n
ClCL9fKrADs40ecNIhYOm/19QEuL6gKN0gyS6Bi4m75+IxIAbWsMrDLpbzoT
WBVG4ZX3WJ8yTumtcvZYmlgEWLwqaO4Jk2LA+0Doo6PNocyDRLBTkG26OwrB
sg3mDxjbuXEq9FOOzwYDI7E9BjSh85oGTdf/C6tf9wuWFh6Wa/rbPy4cN5VZ
xZdVfY7lSeA9StICTkxJ0HDjzE48ZAg99UsOiK+RmzNfVMub5qTZd201c4H8
ReJFM5TNn95IUKuNOdeoMmrJK769Wuv/xJB7m9wmZeMjGw/2J4bltA/8jpKc
bqcYjU94kFI/Z7DXef2FIeUHmT1kPY/Qx0/6ov5nhg0bHTlWsbEmlIG5ZmAt
Yprb7cxXal9vlHPb2WO1Gov9mhHYYDL+ZaivVEcl4U1pKrANtnuAYSwFZtVg
aP4zcnX9fHm4mUs9rl6AuT9YJL/OBp82lI0KhMJaqlIsC0I5mRnepWYshM+c
Gn9+0FL4i7vn2Pg6dhxRYveI8xUEkxjg0V8BizGqIVyzYz00ij3YfQXww/BL
ShWmw9GUqqDt7L9OVG2224RBBhdDSYvz4kNrTvgA1LViivr9mIF7YDHl2b5+
UKKL5USVKpMHnRPZwBB2+nGKfcArY9MHnmp950D9oBVny9FJSbFkRPFPd8yv
mjZ/WkLwv/7NH2l96cNND7l3LHmdS6QWUOP9ZFBjEP6EaqgNJVkd8Sexy2p3
finItsu1XAdiQCsa/l41oRbsfxcCmlVmzPSC93XroTRurC+VVCg2cYhPysXT
C6dmEaRE5Xog5xHB+JDa5XUWA4hSitTetB72nT211aOJP2JtHepTsZ2fyiWQ
ym0tewHjFFXyJonYqxjQUz6m6zsxY9vg3NKNvw5wXOeLhg8Zq3bkmWu2PqCD
+S8E7Yc9pW7ZPsCLakz0sx4K7s0r7mwSJb+9W3LMxrs8vKjboV8fdaLNW22i
mRyrKPVRxndIr47PbepHPz2PLUbzkJcY99+qBTN9U+MW8uA79CdLAaggIg65
Iw/xW2KDqd9Sodzwo027cEU3oqPcynzS5W26TxaOPKelmhsCHqAKQqRhX2pP
Ra+Hv/NwDRIiLBhtvE54vwNm9Ft0ZYNgZEyXgk6FHm2wFfz2a0ig+PWJ4zmg
hWU1UPDU1doL2edok6vPs5FE41x6JSxnbtxVIs5mp+R99GNWnmcYDYfzy+Lo
Gv/CmyWSFLB+8F8O+sHpUpyF0bw9kryn+2VyV1M9sySe8RMrUrQeuRt7jTVB
I3iEMaE+FOPhJJQZWy8p2ttwRfKGLZIWNxZE1JOs3CNIBH5h5IoWtRKIsYAV
aA+RsgA9XcrqDd7EzrndlQvNKXRvPsFiIRbphVNoOaBZ9QQOQaPL/qSAxM95
PYJgn+tUy6AgRw3sqXDXQ66y9SX3FQnMyxyKPQIBVI5OAIChlIBnUaGgKoIG
3UEWnpSQTJMosnB23rYaDteslkD8bfFNxRFVBwLD9VD7DBC/XaqV/hCbTMdI
SXKNHl/Ed4R1+/wTlyzlwaMU6cJH7Uqk57dqDqyWNAChizVj5BGp0EfK4WiR
PqdCKySJiBfsxoO5VjhAeFs4YHx1zAtzmTsm55STumRt2oEEG8Rh29sNS28e
tWHVbtt8elecQP/A+3g0ou3N8Y3JoTIduMvzkDYTpl6CPu13Df80JNB/HGLj
xVg0lBowDdDVyMBayUy89y63HokLX+wvUOt/mzOKH2q6oeitfP0s0BCgA5cb
u9zvqVduKbx9SpcTEHDpaR6HFJGcNzsvpJItZfh/Vyy+ro6wBEz4Mm/eD7wV
nvVz2Dtsa2cQicjEeEjE+drqkIfKIKdql2UpylHKVKSLLAxMo/dwIJ0emGNF
TrudIMexmAfI3deuFKm0CYS3shDOvuSi33B2uTliatgAqZlbnpRABJBIY7Xx
DA8JlsEj1xYP/F7NJK2waBxmbd9DSq4+GCSAod1VA0NJuKCC8YW1+MAoiqk2
moOM9NxTk/mmqOA2bq90y1x0x9ck5BVEawv1CqgSnbFuxcmwrqXVo30wCc9g
74IMzaCPRiW0saeKi5ziRgNqMwc6TjlrFhe94dgI6Ww568/625nJbzAgScAC
WSnnWe5KrOf5MhqEwI4ZV7x2gsgtzmQcVgm+esCZBevhd7dz7E1AW7t076iX
r68GD6U+4Rnv4AQQGcyZVzJSvJ3VxE/XEWGktl6ANI44qn7cCraBX/+h/kUb
AduPBgtkCujA6PvpcPddYCZGlMaVCEZTu1kPpE+oGFqxX35Bz5Q/35aw0Q0N
B833iRacXH6I34xgwuPqtL7gDCSy4q7A1doBrzx6Pecd1r9AnivzQ1F/9QQ6
5tJ4dN1+CkhLYDQ/WasOykq+zYD2wf+Iclk42IPCGP8jAaa6FRU9FCFsMql4
O0JYnB+gmJnu8UgkQ0g/8GcXjGr1PByMmcj27K6Ho+huY3UZPdz05lK90qo3
XiY+m432xwH+lMkn4BLc5Oyg+TvEszD+wHy3rJClckEV98iEiEuvcDXY2wZc
rzQlW5C58UoSvgF9MT4DHdXa/L8S3tbOfQTkNiAAdhx5Y7RGJoTxqVFU+GuG
AArq+DWIr7KZprM3/ZtYjw+n/X8AL/AzWTzReGHHg5H1Ts03grysqohNqiiK
xq1XgtCuJT+X9TOwEo3OdP+NkJ+xRsE7ihwwrEkYE0tfQ+r9QJoOCPj54W7c
8qNJbmns9UiodOd+nCSYplUZQFEyMqSje7do/B3lYLTECTMsjrWcHvsHms6k
lwmr5Jvf7O6AxeG3HVTWvf8B+Co05rk1W1dm7ds//kpdDokI4msWsfwWviTL
ZCUcGM9EejboarCRJv+vbg2MScdBa2+zqikpNsUDsM8I4khActXtg0P0iILb
+aAv80eQRb+CfO6y/1/sL+nJ7+reWyQ0dSnmsAoS7WxsfSGuJzeRitpMf32m
tTZlPTzmgRfRjWAu6q32DwiJSjtZlFZfSvGvH6p8la0hVDOowNy9jR8S4CVf
ZawbueKw1vjL6B/gEjDUHZc1QDnQvSSn8hNtTy0P6tko4RGP7gre5bYxMDbn
XKYrt8GuyPLxcOslsn+XFCxwsOHJd3iaPRNF4HC86lukIrG7+e+NntC0JmN+
vaartgNlTfxDMdDRG8/ZoTx/tgbRoh8AyMLJ2VfPJ4B8M6lp2+kZvneda3n7
FjKxrMmGwmiAGtoeef7KurTz8Axattio5FRdW3BSeG9CVij3BsFJUo7U3m0L
zo+qJZ2ZoLfTDBEEkSUsF8yB4xM62AF+MizA/e3N9D4W4WeJojU9m1JnEY/x
x4Mb9dW0lRvwVGf+xxC+AHxW85MQrv4zGKKo7/qqjQ0OiGx1Y5g5NIkRWOL0
3cBkx1rqIzNJCedOYB/IQlIIHgp/DkJ1E8EF2BNwgVZSgWdfeai7oKpM3ciA
8Xp8zl8b072rNKVKeDKOcx2KnUGsWjAC6wHMS/CJ70W0hY+B6V66GrLWqwrP
uF19UFWiu1L2I9Sn/9b2JKDsFwOr1X+jxaaITcjJ+UQD1e2/7BvCPBYydWTz
BkB4DlHKr8ED5k1mSy6kuEv7s+OAdtuh2gd8C0Zq1eZM3kULfIlEuCr7rmFN
30aWjl3SH9ePAB37QOjyHoREoB8XmW+madka32OfHI3xztIfQrQZfS+5l0vD
ORNDn/02G6qxQUExIYkLsxw+K1mjyKcPZOL8VA2O+3nBOl0M5pI4+PPzF8BP
A0paPo1Rs99QtGEQ6HUHsTJ2msN7WsyH+gvG2a0y0CyJipmeeMFpzeDBfnR7
dPTLKB0+SQ2PV1JEi4jw8o9FcqhQd0xTGu3mUs/LdYzMVNf8lJC65izUpbRB
QC90c81FwGD2hTj3cN+T7j69/drhb72igUvmCecGoTNaj+8aIUlTEZvXOIRG
bOnDM0YUe4Ek5oJMMyE4tY5g0QXuFDhQ1uvEsO3iqzR/RKlxLNglHpwgFmAJ
frlJZt1Livyx0cYVUJYbnCeM+AxANM8NOkqYnIBjGRROg2FAKJW9rTnpX/CI
M981UA+nG0LBmLC693Eu81e0F1ytXCf5Y3DvKGLRbZVpkRQcnAwf9qABhTmZ
4OVSAKGdmJ8bAC05NuuOIfURw7lA53tuckjG9PYLGznOAfwaPelUeQO9A+YZ
Xhhf4HpB5QOv9BslkcPLFq0JD3tx77P5kiNBkvCseVincu7lkkOUuPYSr/Ie
JZPKO4RctROYBkh4dFNATkAGWcqDjFuGSQsuVl9LVzoyHdM+e8GZSx0UBGHg
n1QhM23p0IPjRsUGZT2jNGJ2hzhswEvsAY4sJbFgQiDLcm14/vswTc0l8sJB
xy+3M7zB6unJA/qWZPvoH3uShm3vAxozVw9zjp5sz93p3U5/okUFXf0gZtir
cRD1YbRYYMz2KLkfH2gF78quy0o3GneuZnDXxdQOGzbRln0kyECtPs6PK4cj
vVC2rV0U3hl4ObPfE6PyzzAiqJ1is+kI6QEdRYlwHqzHOpbej+L8PyMU6LAk
sFccldz6TxEhU9AnBu0odqyQXNdyk4QOkkHZZjoI6QGVBxHpxOOHYgLM8OnS
HmWaU5klt9ow0LpvGOn1DCa/PdhC1XS8HtwU5CkDmtSensG7THFg/cEoftf7
7n2PfXVz3suRUXApnJhP6bUsDSryQbOjJ6WqtD7E2Ot8l6nh7sR+ENvI3nZ5
8zY9bzD4PtxPGFLhErvk96F08ApkEOUNRp+4Clrw6ljJ+mPsDX3wD0AwGFJl
gp54HZIqeHyV6qcHkaME+2Rm+97RfxAJOkbchFeE8CzNa13pqWc4UIuwJsIz
jXa7NgZ0Nuc2CvcccU/dYBgQg08nFi7K+gfpuUwf+UUgFWOn7EhLDCpD1cLR
ccTAIFwxxSCt0ubbiDaqyck0qpVCYY+7z5LzUIBBItCa0DlQsNcaFhWyMoTa
m4YAJ9ATnHQ9Wzmilhe+SLP11e+bfvx4t70iV1IdzEXEEWbj2mUO/4MSOg74
5uqLS70gSsWRcLz0/0MAhSotz4gP8aqytDoz/Mc/URZeimXOA3R1l/G++MTH
dlKmxXRMlKOxxnL5gTWplLQMWwzlZlJozrGIUF+WBJn+a1Bo89PH5dk+5gCd
PIl7+vZ/NcyakpPgc0uPHFD6akHddezH+rbnZY33I9WPyts4s4e/Na3GRthM
NWb5zVibAZrKjBBpaPk4/0pfGG6QKkFx02uAU7a2szRubsUjyuzpwhT4ike8
ANSC7b6upeY8MWbK+hwV7ybVHK6NZzTkEdh/8cx3SFhpFkb9VX8V8P15QnEo
rnKSeYInKu36lu+3RoB/XG8cHr3aC4rrVtPh4WUV/W3y1QfVaf+uz1DQLZT5
y0VugH33rJTM5X2DfBSt3o5bIja2mqXoR+GBbtgppGNjPCAY9te1aL/0NPT0
rtcu9CdUSrG5T2rE2TD2/fC2s3UyiiuEIxTsx7onRCyU59ezrpHZfqkwGDat
tcoLYCpe9yogGiK3Y1/qgZ7gQ20kJBS1oZIsvyHO3mohqnxA/6eRHTx0/KQg
TGf8np14/qAzW5nXZeSWfJb1GfjilfGnppujUFTkWRjRvSc3Y8L+nXqr+Y0h
C+yelOLp+xwq3ebn3ffkF2nbS3avQ1mJOK0e9KNXvpftgDJQpPWojA5Rdez0
n7/XMvIXOYy/UTNE7AOeBKY94b0OqyqTLU82YrEaGPoNtPsqdfwZgalhGkB1
DNzPQxM19nfeC8HIDuRSSQEWaz1wPqMjiOz8rqvj5pK/97s3UG6S8sjZ0XoU
x9Ub+n+vC6cb3NHRmbU+Kpr2i7HMWXCQnr4rod+1Lf7xeoXNKiCo+BldPavs
F6HEnTnUwB6w/TPrwVTKZrvUPwqhH0Cna0ygN70uyfOGMLiPfWfBmJ+74ARU
fhaFG9bAPgUtudBl+upCqwLlgkpsUyRfhqyZJOqhR8HHi8r0pNiubCkrsXv/
Dv9zHa0yeCThtHXkJd0W1DXs6pnaEa+Ltk4POz2fM7Nf61E27lD+FOtlyxcM
YRfCaWOmY3/TrLEV6AcpcHdfT3oE3OXv2jnMF4kbiT1IiVLeZuWpOWL+6Rmb
HBNMApWWwddRVCGr8DfdnyNXEcTZ4rnL/bQowfqFq2zjEJDSd1zHndcY3/oE
qx9lxwe2N6YQtpLdb+/tedtWoL42aZPgJGcQGNSqL8+ychw/hjH+Ea0bBcMC
G21slA9VRZ6doeAhUNryl2IIub+6Vz+ih3qEfF2O9h6mdTEnCjkAEk3cWieg
yf1rKIP7mz+IpiBebnNcQf9g9XLucp54KQq1iKc59UeVipKhuoIUkgaBL3VY
f2BI+Wja/5RwUxx4xJkm0VapCEAZrfWlvBZZBzlhrCylRoytUjidiS4euQH8
BE2XEOTLAEvblVDFw8W/Szz/4CvlQnxlyVIvYMf0n56lVL2KizRI1/e4ZqoR
vE6WE0Wzkdj0D2ZlChqD+sP7WTI9l1phu3AO/NWGxAKFUMgP76islq8j8ZBt
Z9Z3s3P8gkP5CZVI/eNbHs2D0qGu8JItjaTeI0QXeqLqPlXSItjSI4SjXQgo
2i8MdooHgZDpNGrcHIvjLCN5tI3AwWGe7rnUoAUjboUKxD2c0EUBJ9gEhi9y
N+AsJL49I88wY8Oe6MUAcc4b2DK36pxAa29lADkhhZZaU7V0OCpdoD76LYIy
vJD8bH6NifWZ98sLKZBEdrYqtl3O3NzuAE6uvCWm6PAHavyX1XsApanYCMk9
mo+xL5o+vKt/nyIC8YaABLbYOsOOQkPvnTEUfmh0TgUHLoFZ5Emysjdwa4iQ
BTbY3y7W1RclPFDdejGPwbI9pTr45kpNkJz3Ff8YyHPSJHkpq5gDT96vafHp
RODNCRD/quYRY/cGM7e4blEnQl2J/Xz8TC2TFVd0+R1PaSjnU8YxZG+8CdXU
KTGQiR8z+bTc7HqGAxKKOz0WHl7GGxLASREkgOr8uR9qP3H+1EeURieCn6JN
yplpkVD2dtmJfYxWggWn2UoqzzN4BiWg8pk2PmN5LZBK9u8g37g5iCz7qlcz
t6zFhMHh1X1W6WvM5UzKoXPoqCJkkzjzQ+EECfyKoaoOUqgx6of3kCfs8Vin
4wIHrONoP196VDZSUe67K8T2d30fJ8s2XDH1t5uddWotSKFYypHGfdoVSnK5
ZtIvGc8WMgkHoxEy2x8q0Zd3WgJswuPFlAJuzIizmrYfdcaPCYICgWTp44/T
hK8DEZOtR/pcmJ5OUHSsrLODa7qnBVcGZmGwW4SQJb7+RkMnc9whVtGvDWsz
ddnouB5uNphZ4jJs0pjzctOe/KGK5YzPmlrEeL3gNkawFWDhzD5EBZGgjxXP
m/Sx3YaD78y1b47r0FYSewEEu4etuLaTiXSP4XM4Y2mPlXbucdfTdBVpQlZv
Kxu4NBIcez8b6KV+64rtlEudiNRn5kLXLsHK/MPAY8MpXS9E6OvJz4qKCucA
p/wjui+SSsE8+QSTjYH1cKSojZ+P+sYTn2N2de39mb+2LfJBu+zfQhj/SLL3
Xu77REpCOe2J7x/5sXClBoZ3dEfTaRJ6axVf26EB6zmT7syz3BqzXdnBZpBg
C/HZB1fhzxdzNKR6mTbjlVKizTRTGj/oXGep88kZo+2dGyhvPIEhBg94ppEZ
Fx8OQykbuM+m+GRHE4Llxcs9n0eXWX1OagAcwtvBBju2fPhV+wdolwwdz0tx
LnVfGi/7Qsly/FrDYq4D1ZzcbVNrPsRnmvj4lemUgM6nkIiD4VHQ60mRHaB9
s+ZoptWJs3GgPAPdB+HMEkbSQ3VICriXBsiZbMtgpTypiGHNdEKSgIbmf7jS
xq4c5Af18mtVgxY3rFIe0BpOaLfb1bbVpRaAfYBaUH5P3fPwEG+zMvhrkBYQ
tYXzgjUbnIXMJHI+3hSOwNlkB+r/6pIhmoTFz2N3QT19GUROuuQjIZZbsyHR
LgS/kPr1hynkPuiVt1gMmQL2TRSNc9FLL+ZK+1aFszlJEEkq8CTj4ecubm4W
om9UyBVjgSrcTIu9nHH8Cog0P14D0DfYLESb9uVh8iinZT/PUd0EhRR8XDyR
C+oDepBlgGMr1aRyISLvG545cQsCu7srTjPyVKt4vRubZU2Xx1QmFGcAXiiz
A59LJvizffpxyJgVqLiDUt5PCwYUroBcVk+OnaW/tk89l15KewwrcAwJCZXp
d4StMEWsyEiEaYiRQR01EYWsrUG+oEk7NbuYhNd82UDVISEROwA99f6HK1Qi
G2hTR5bT1cx7QCCxC8pUXyXttx3gGhMbibQV7/un2h/4A5bYBCWQitz0m6hU
zAyJ8mKC+s8mYbItlc0EgXoz5CyusugB9VvRTO8FEW0TQxq1i4Fax0Lh8UPW
xJ82ld5cBxQ5chixehZoWpgx4dZqKxTw/kJv0EEdz8lfSd6MC9ma0kHb2hjq
9tyErcK/d673bVJKItD5/uIOQIggvMfLSGVms56j60JQjRDRDNA4AUy0Ykrq
bkbni4jYztfmGdAaqqVX1HwRQFWW/Dmml6Zeh92+LEr6t+4u0Kdf0yVBqRBi
ypMCrgqNVnBFSpC6pkH6CWhsZf/v59/Rdoy8nryMAnmD/fy0tMOQTVpWcLMI
xk2ov3aobJRw+lqHGtClZ+yjCVGyNQVULCgTl7MDCwhY0Kw4uhdy4Wu0RveG
rDCNv2q27/5FY0fmL5tayeW31qiE1I3aaVXfC9ZXH4xfxc0Xrgluj5kpK1lE
kW3rjnQnSxdflTtMSSSQ/Fy45Xr4/QCQatQg/6GxfTwuHpLKaWsF11kxAZ15
2V+hEiZHIsneW2u35OlOupg/lBdqmmSmqCu/JdQaLqROYzyG9KeDEY35rOLq
JyXy0KtiuavPLakligP/8m1lk5uCRjA/b3FsrwO7/TB6c5en+rKyJiqauKE2
RX9JMzrcp/j1LGYX+fi8kMOKLOQZ07Bb+w/jFreazYaAQS7cFsU9iRCRkO2T
Q8ko86loBt16daCIeliHzxwuP17aLAYrNYVoM5oaCX39ouzcaA9DS3HK07cs
zgAzSnzBMjllHnNBGUueRrTgB6e//atgAnjxOW2XT2GPIoGiFCYP7CmlURB9
O+PZHKn/TEOXwlFGEvLjZ0mcfK5Zivcs18YpsLSvfbeid5cCzawzXJv9mm9G
bXe98gi5kyHyeU/4gMv6qmnba5Wrls5PjuoQl4Ihk11ZkHvK7+wH69Mid+PP
JiFpTZIPkWDMsQovpg+ryWRxPY3Nel0o9JBRkViE5OOCsqTsiF3/dUMxFJIm
gLFBc81dR52df6z/pPm1x3V5VqCZRnuj1qPlj2Ui1s0rtvxtNbdVaiegL7zp
PmQci2bHUDlY1lcY7+Q1GcKgQIyr+6cZAX0xo0Pd/SMN/4FkXRw2NDGWCHqv
/rUo2rCdLf6Jf5iacVNAMqjCjWmZ89vn4eL0TysRSgv8MKxrDGX8DL8adxzi
roTnP0koZ3fUuYuFuEfFMw/bttfGzGTZHR5D4CdNV0MjncQ+hdfLyRmls5Tk
qKkBmIuO0fJqeNv7RvnWL+GYCVmbCNULilBWuZ8Aj3trLbfx2dcKImF106r5
PMUkKIeUV9sFJWRrdijpPuSpbIqwj6fnQl/ibDPVCWwdxzLb2GYINUPsJy82
sWQYj/ufPT/9oBtbVDTBtlQFaI3SlUZyGnxf5XEGuf803QAZ4xqSBQIlOU7Q
6QIMjQuFaxboS6PZMHEy/rLvzU2MdCd+5CeUnWTinUxP6mY95/T10E9yco03
/1jNEzU77qLMMOhC52Zp4H8G4QhfEQZc9tD7gbTvpRh/TiIehIWj4zUQPM0u
sf/Kn2i7VxJ5oNqxJg6TbNIOdoGzef6Qx5Wk8pkyPrVW1zkmrHJko8rNRYvs
HWDNWYUousKbuKsVUfFf/auwz2IIbQ5Fiqm3UzP6BNWe+fGNyleC0jrK8qWB
yg6bv/yafD6Img1kmzuuU8iQ5PFfYum1OTfyFUMOmhON8aNNoGyxSfbARTGp
MG1dKHPAbKECQnzTdompjSetwwwNWAndQ8OfX4+pW26EVBqBhh1R6AmzSWhg
gkTAiweaEfQiPa83AST3uBJdhgpYlx/fpJ09c99sTeRBeD+r4PnWVyqfoxlu
1fX3qwjCIzUngkxnE8KqBbZiEu0al37nzdeDGqzTwqIiLy2JSsjSQeaxJVLo
5eWHy6x16F4HiA5fF5Qplg9miZ0NMcmcgtlkzTklA+J5Zsjev8cB61Q1kxRM
z70Fzz6CQ3YEdRhC6/ntOrAg/sTI+r8CdnqSyyOo0aePj3i5+iIzNNwYA6f7
srUHc0WLbSRE8BfgaBRr4LWOG23ACzREeNiYOuA8q5uoTY78Qs6ERbXB7sNo
JkdJAtemsPkTVuU8ladAB3/Om7SJTUg4WQT5FH/9esKLIkxEb5Kl3nA6VxyV
OkB0eDCFvR4IbV+JwZasoFMtXg4GGjypxucwhJJUOiSMaD+brJxpJurwX4+6
ohc4Nrh6j86PF/u9Qh1nCQjxOzA/XGULcBpKdDzKyCM9qwMZ/ckw3303hRQU
5YEr9/kulec6tLPztEzpU1FcT8+cwPv8ZGQKRGOu/N+P9Af2f13jc1gYjRbA
f7kXIy1yYkLY21NnrEQzHMic0U1Zeo8FLgo4ZAOKnxC8+FuMsLxMb0kU0dtm
r0i4DHvJZlUQOQ0/iphtwO1MnrHK6Ly+X0nrKZcWPhjJ1UKc6T/1TNabLkbs
lMXsFBT1+9LgCNmGayvUY8BBv9138IO85YcFt178vU37GGqcm+zkjdM8twiT
Fje7VC1r+lzZFeyuKiPNGLLr3da51CvezyBgQs8Yor20OLnSByS3Jum+vknO
469lGVrGyvnCSvS9wnt0eLAhZXqHIorSVn1GxagTP9EVtkg6qTPs3X6fLdPE
xdgf3bov+Q2KHG+XIjgNiA4h8neqAT3dzjK4UxEeK3VV0sIinasWRLlgF8g9
d95AAphSPJYBQBYrXrWf/qtnlRs+ZoyYWaKkl4MC5Yrdw95ai1QolKxvQNVB
ifskLU3iELRP40M9EQA9FCAcdgR6KqmDbUqZZYqwKSTwz4u8hZEM9by10/lC
nAq/xElmSGNJT5CN56QJotjChVLv8yU3ad31NWP8dQJkClcexDSyDX5iHBVa
ZM/S7thZg+ozoVgY/xx3El04BHY9fionxkHlRLynb43p+/+9gfu6Of9cpdNs
ViuchAeR/hHwhPhxVV9pP0sEm9Gw7WHxqKLB2Zmymw7BgKG6Cbz9K8qlAENd
Y83iflTzkbTAeDsNne5S77gcWlwvChrzvY8EQmV8dtow6QvwDCKEBeQ+r/qM
1+7wbp+nrd7QDdt+UFtWN1ylCM3R53HqTFXJx4J3S0twS9sOdOmJJgTjDsK7
izuOoaf6QG3Ie8BFlqqgSRVfDqEU0luiNn6C27T9pBah4FOXfbrnwZOhafv6
xPCGF8m15iUSwUXJ59g5FJeD84GWNBkg7tNy2vh56xGZJcCgpHautQjLTKg2
GPkyBdK3ZEH12gLZMbYMv6G4sQWO3g7mdGEmFFDK2O7CNEdKpK84a4dUQHQj
Ft3D6FpjhT5bHsmpcMOHapxqQ161Bjim46+W1jNqAKHE2gXhh20v/hoxOBcj
rX78l0/UvGtvq7/+C+1E6Wa1mWrsO57vcG8fVsQ/PmTwy6fBrcVMUn7wKXJq
/tKAQeLLnaZSRR03mCDwSH+ESdJNJKLSMaghDXNr1At7d6o6zCcQunhHSByG
PLFFekcz4zqjdvF3KxEdzYQbw/WuJhuwBYvWgqLMRWy3nO5GVe7klXjAdRC4
YoD88ZK8bUF4qTzZIE/vixAmEHgkc5dxHw49s9bbG5vCk9axgVkY1PtFl9BF
+y6oD4Qiqh+r9c4lA6dSEilcKNkzJ4hj9Evlk2zW0JwvOjYXQcDNOsVQGGFB
4vYqbU5MkkI4vELbopveTobbNa+afps9FxmLhqlqSymRodZ6PgwRlzoziI3/
Z4ZqvT7PznxUeTf3Ej+UY/kjsw1xabGfmDxx11BpRPl/kj9Zl5fN04pWO+Yq
wyJnWBhzrTHPaCaF2/xOu8mWWcQ1B1ZCmJ7a+NA157rqkprOxvtvZi/2D0Cu
LGWyGiCp7+y/OgJdaovCPvuHmXlLU3QmptnJZEv5aR/DMoMcKvE5fis/Ixw1
FLUkEYt+5TCFtFRK2saeRr0gt5FXPZzogIflty35qGuhSwFUS6hDyiYeLrv1
JBw5i4nydmUH4AhvUwd58CRFSedjA56iz1gPrzFuwNz40E16ZGIdDXZu25SD
NYIsbfdoK5yYQduLiHG5K7Iekq6/BmJPlGuV1HyqifkAYtOVuLNw1Vrn4mS7
wg0RkIa8cYmy2Pdqqz0mH80nrqnnv173oO+GmNWrGvv5E8sCIc1/ROCbJxaF
5XkEsJibRXon/bbfQRwfyIM4PxEwg1/hTF07q942y5XEhEONKYNzvhFHczkJ
irlvScacC620LB5fy6ke8HFudTPmRLAS8kFxPSfNFHI7aoib5QTmd7qtBjfw
gEOHRukqbDeB02Bbo3iJSkOvqksFIYe4Ez+SjqbrSj4yDoltEIfWMI8OfYyt
rKwrkDzkeBd6nA5XftYQeqxelCEWnvSwygseOWS4h+95Nlz9Uxd+mocjXWk8
M1J7uDlkyC8pzV1yvN6SUh+nCot5rdRIR5fbJAbtpcw+UQibCeTJvZRuGboD
st7xlahFwYDORfw14RKWZIauG1RxF8cYhkd/TCv0gIAa/JStFnCL/L9Yrwfi
hY32mxTwikcmwn3Bwny0GGQXIi9NGcEvB5G1JKxVt/GtRG0SykjgS7Cb5o3s
w5ax/et0fCqKbXhfSgyjk5Dai5ZtMnUcqj+fjFPSC1weAVialQiHHeGHK2cs
0/JEwZBwXJ6pZ7FkAEYBuv2h6GiABeXHbLvTANsdeiXX5XJ8Qkd6IG5jXv5B
Lx+GK6BghXsvMhduX9P007gEBHZR2BysSIMmqqAdYUuXCaOAF5TfrJIX5h/l
PSeus4NnVleBbmFlI2Gbo10bRUep6DMlYiGF2Q2sAVwY++Y/+qH/IjbAoCeF
toB/Zg9aSpqpRbyku4GkPESngjyiRaIk4hqEH1EM5/Q2Nak2xnyptEBRwF02
UZT4OX/EEgi1hiwvNBNLvFWybz3lj0ewEl5rSRZYEzYEoEpszFE2W6EhsTgC
RwlLPHs2RbuPY41c4ZWDcJN0L5mkcYRTTXrTbNLkmT2uuVxPsGnD/Q1feCQR
QlzVK60AuK0sQUAMLaL9aby+KXiMVUvBlR1F/+11FEVoOpxmNzyoQZ/+6FDW
m3O7Eld+IucKhmnhPfFAJzsbZRWmmZYGn2lyGUx/IrEvdlluQUOc+k6qo4xl
xOKbKJ31dx+cIixZd4diefg+D1eKPhxDQHiGPNHMHjT//Lqdyy1Pg+g5ui6Y
Bf1iJ9StNXLOuwavzWeWsHVLmufEpfT8euQ7Z9XXA/WvJejNojQSTXF8rMFw
djZqVcxGyFFvMVbhMtskMhhCxYF+Wr0lqXB0/YlZAYvEzdlOweJW47YCsdjU
MZVP8ogIwDXXW0WgL/iODMP2LumFcKlNRm8Mkskw11eBz9/HinlP7pVOP7YO
gCNJiAdNJCsX6b1EM4esDY+4TZt+k0ZIoyyP4JjUaA8eIMXBqy8wNSltJnh5
40IMZ17okVJcB2Qw+IJmsvSiWUOBY8ax2zAFcID1IR+PJVb5ZwEagX0+hveY
8ciuMFlyCji5GROK31hAaGLHS2ZmpeMsEgusTGYfQ+v1clf+QC5o4aWHbZzA
NLpDftPLPcUlMUT8T/i+x+CEx8t6SbNzvJ8KUK2BC8sXw10tUzpq7VShphIK
Sg5QiORCeE6Idkp80gCpe8U0X01wjEBz+/giszi/6WGhSj14FxIgRIeXge78
yiQmxFsWFvgKsBPuRb9F6VNtoaBs3ZuSoJNPgZNqER/NOLvKUnVwiMTQ+R6/
HULLdWCdP+53pErHksv8sQWBYv5rCThH9nn7xmPh3giD4p4SDB+nAaIup3B3
KDJsMhU/60J553VTHAFwFvOrzLvXu4XotL2o8szvNYn2O8P8IeUxEjL7y/Bx
KXn/HcOw/60YHM28ZzR5UklHVJ5O/vHDFAzE7BZRhOzqwlwjr3+wFolyIagQ
4y+DChwmnVF6Txn8ETCRldHJpOp9GGIhsBv8FIHIokkXkbTPxrLfSd1z6qx6
nTjFrtFQlbGcxqpyAnULZ4mmNeKkHqIJugtVSPwog9co3oJ/0E+uprojEhaZ
KJGC/LK1ME7djLquqXiWjVYPoix0NtYLl16B4cBaUzqlFX86Hkag2KHNlvqj
z0uDYMvxGw81WLsPUyPefsswZwhgFv8TqC6UlzHb6kpl+vnO2TycJlXoBLgi
oycAKperNkWQlDLWiS6/rsB3VREIhT49hicYLQEzveMAC4xdZBZUHRaglIBC
G3V/AS+qlyPkV42kgWZJCbuxASNUxs++uU416RKBT4Pj++ofGjm1sibWKmD2
y20U7ROA5p70iVAghCFjA20QvVjYVDLdjD6SMdrsGcpUXyweN78WK2/vB8qs
4vZr5UrRWRQI2Lhr3rDxb7aR8UtH4fw9y10T2EnInO3g+hPxhAF994IcYO59
t8qG3J5A/pWZLpJ/BsC7J+qPmwL2nSWuhKSl81eXwYGCNb0s3a1kFPLlKBHT
9p51Gv870VSOfbvdSWYqVr7M6GMJZO4DsvEuS5A0SdmEPRHoYEhnEipFDCHH
fTVktgSTefMunRr8jceqv1orU6mFx590WhwMkkDjOvg7B3nGmzizrU9VfsWM
5EtS6UETddOSOOETDIY7rZ8ZfyI1wAFaT/4XEd2lXu/F2sNSaPRLi9sh/Ijm
hq27U+qDGfauUmT0V9plPGzw4xhZwNloKSEDmPXGBO6v9gB6xTzERLgKiPp3
wINbwpEXSw8986Lkdt7khUzHcdeJv9wvXgFAgUXM6/5qpydJWRagM4UREpod
XtcEsSil1PmO4MV8RPj2A2eYAwHedZk5vQ3PVdHQsROjc9gDgJZlTI2k/oU6
NDoVHv1f8RnH1X5zfYH6p77bLYJkcOwY0H9cfPTWycsFCrDA1VRTDMxnZA6m
LkcP3IcfGa9hJUu+HceSY88qpsmBt4XgkctoPgLx+wrrC/lJG8+J27BmWa+y
apsBFJGt43pL2L17QwOSYsyE8jBX0oQicIhEP2p7AsRRFXHxFh7kzijvxjEz
dWLd5QH2K2t15BhH03HUP3CoecomtJiOL+J9W5KQWPAQFQEYFDCkzmZRlOtz
6LujbGKStddZ2KuZhgeJsQyIUzDe/1AGsnfDChDWjqrTn6VfKPCwk7Gu6bRz
Y3jOS4FZyf2zXeiI0ETdyuEtFpOE7frMY7/MMxJLwMf18G293bTAHZX7s2mn
rGmmBfEIr4kpx+4LLNwZrWVCt7UBj+Z2mCxEx5cls4L3oBVLdht6mUNp8/uW
hbyDj9Mqg03N9N6qv3LkgB/YVVw4FSovBFaerQgB6lFXXCLF1NLKt7Q9POdF
CHvpdPu0gYi1Pa3q+DFOSjbz7HOK8V2ARDPwtFDHQcEwy0uU/y9hclyDfpT2
5Fw0fmRMi+/9/a9fliRkWvmIuxmZR60W/5m2AQMH2CBOM6Z88ioUSWDVllpx
SNsu8Vy6Yq1VMhWYRGLtR5FlSYIVoFwZkW/LAeJ1gyBOO1aVivzuHIGVdh+d
DC1CFzSp9pT9msO43xbmi9vjvEbCEjc/Z/sE9RYQOvEYjynSqhvfRSAMfjES
yYhOEzaed7Ffx5sUO0mPMyzdu76lhZc0BoDbz5W6NNCwihn+LAGMc8HNVlb8
zkiysn8U7Szxm+xlDUTqd15MScPLUwkrbebZaKyLMnde37r2K5mC51Mcng18
P2SSRS74wPUgI/HxrL+oyfBFTN2OfG3xVwpwW7iC06xLeE01wWNkvKH78psR
ejRF5b1xKWvuBoUFmFHyidBjST40mnQmtc88cl9Aheo8APXs7/BorY6b803i
Aq3cs//CC9PwLCOllYZeIAhTegMWZ2Tt+4pSxWBij1x4vYQ+1yaxUXbpLvpj
hVMvGlaS8CQ5hS/aYLvbKXc/W9XHHv7DDfzj9aUVZvTZz4CUxbLr0Xg46j2k
5svvob3dH7mvQe67PJl92GzMPSuQFFK7I/NkPq8PgKiULIhNoUjJPPLigzhG
2jjTQ0tuu345JwNxGq8jlyFF0oFDMKMSclm+IQUDi1qlGuqXq8cORpNwc0+I
0TOCTsQBp86IBksITgC4FXbJPTjRMXnf7esg7+lE7pqgDgpJ/ivtf2omh9kL
K0MIACOBPedtlWGM1FkLY+rVo6qUOjinMPUcUSMM88HHXcuFBJq+iwxVUZMo
Z17Dui/DuZ6nxT7dgYub0a7pa4kAlojCKU5svMUlZzcqaUzSxuJTnZEedCaW
UeDHFyP+6Kmrod34nvM+OKBNeCXILjrOUHG00GKQ9sue6uZ+2go/BKFI/9rT
2V1sRqeTuLQiy0ds6+P13ZmCTLTXmEbQiSsvOrh5CGXZC8rL0ILeOoz/bOAF
YfvRGfD383+TGAAcKFAJeBVwMbWrHBnQu4/DCtO6nWCshX2XDW4TRongENPJ
wMHmDZgDH3KGvqZPxT829dCtOhDf7x72rWbhKZp62zWmR0Zrnk7kQSEBhs36
4Ye1XJ+knBOPv5bxA5oPn4ekh7T1qTDqEKmfz1bA3clVKBz8WQuM+mcQk9du
2JvwikYA4QImFjP86pGXRslQMwTL7cKWdSpOpPSU9LQu1uqzEVZgUtP7pCag
c0uHmel8DfrVeF2QeH3wFz3XNo6x5bQzVNx18ofDXMIJwmPQh5N/vrEWTdvZ
CVrlzsHfxiGY65ioaNyFn1QNJpPdayK6z6zue+ZqdsUMfcbjtiX+4q5y/Iu1
LuNykGkKWMISdyLVSrRZxki0u5NRMtf6x5KvzaOuQBfLOL/c6Ptld2RcAwLw
pcZGUOC9exVIGiQzjcQcKN/TtDrm05nerxSlUwruKaUhU1sougJGTeIsGAsx
5fQiY1Fac9Qp3q7dparEIEgd8lekaxp0BvcZDwISVx612kfPs+dlkgCrwfDl
EKyS+ScYQ3A1c5WpfCrtwsb/W43gVn7zfLrmbmp8vdxegxGCZj/m69SvYHiv
shKVLr6ZyOro6df6Mdj9liOzu7F6Z2/U2uz+NzLRPhXde70HVFNjX2b7QF3y
e0BUuIbD6MzbYvyUgiWuAltBiyXq6m3QH7Ve+13hzZtg5+h7ZPcXW0MKINpZ
+6Tqs0vj3/eGjk9rX58hHUxfYo+dBayBhBfNuUm0+eojHqR4PVirPK/1Lw0Y
iPkukmwlbpC/7Re+poR6/Is3yiv3nQW/fnHDrwEXVE8z8rUTOgB7GzTuV4pb
M/12tboVuIjD2oNO85DzTK052/oolX6xYZmmWc2KkHTbM6ah/jGtOWso4cvZ
lHzoWHo/ZJoSkbPxdJTpV4wtnn9gBtfdqSAXFwaOaB6wHsnCs598NJzgTZKv
Nxs3GprQ8MkFFm/cm09PfiC3PqCmJ7FutJQvu+mV/7DsWhlgZmiyOnMRZuwT
Slvn/0VgTTQgvWgKM617O0wGIUy3mVCwMytJvnyIPtIVckYsgyOmMb/I8JJq
nVv8Q05phZ1NecKYj0qjjvMfxCk0DLPjbMCgIqMQhblfvVnF3/V56qTb7m33
BoCvHGrRdvP+v60OqvxXQijRlg3U+HFYSVoWu7p+2w8juSOPInWWUTMfGiEI
8KLLFwcD88t64OFWJkOUyKX9+Wtb0cAHTofpe5RnhPiK1KwF97LgqASeEcTZ
wynggdsdhcAn/RE8+dmGaaT6UFhL93PQN1lKuJKk1LMeSQ5WtjnovhpbkcsB
wiov7PHORDQFyHRnW5f+P98xAsrqRS3sNVO1yZKOJAo65GbXadY4ekfrB2dO
7wOE6qq4WtBgOQhG3R8j8sHS13QC0OmYO4sYlv/EStxtH0NPALvubr6ys//B
rQTeZHHRlpINpkUbF2pWfC4U7zmKtMMoel1NdxuraLtR4mSAF6rAzAXUFZ+w
QGNEsz7jz3apiqhTHOu3Wu3vyZohwUMQrgCYJYyrehXQh4PYziJf/WNN9W2L
O2nU73xB31zVzJaSZKfbAZa8xUzlbEkekUUnlJJMwyUNZEG+U8H+6RK6SkDO
XRgaiC5uzVTV6kki+mDsRDrHanwRgyCDgf/eJ6cshBWCxbzF8M3IN12BazUQ
vO4r6sX7Ypeno2A+KdCNqEMq9px4xalMP4Uf5MlEFeRXCxyDDQtIBkQwzn7+
p2W0sluOn1+96OvIdd3okDj3oTeLrmTTWEr4TK92PIu+C8tYJNZ6WD+AQjGP
Yju9FQZcrmnVLuIPwqshthrvbm1YG9yLEDYZYcQHLWT4NU0rnstCWqMJzwcR
No/3wWOXrjxPxL+oWHxnTDA2+FJLDqonE3eMg8VhXYIMQu9dbGUvVwjRKgUS
YHitQlAQpEuzruEYFBRB4Bu26s6BeokYpk0xzT+yKk/JUzgAGl9O+pdzuS4+
oMD2rEWpQJ+CIoFk8GwUWz2pY1UCO0AV3/jZ8tqgWhQxqntjHKGFIQszVc4j
IjbIGiTTChJ2Lw9LuX7O+/34v0MnuiQi2heloVBJ4MFtp16dC+QafM8m4Uls
3FXiKayFdlt10OoYeCLXUXPJfmX29mg6LyHtLtDDjZOdX3JGeuOKxItf33O2
34EV2NyGeQCX9my11MPePUm5qk1gdupWf+KtYux3vX/Zimo2XpGdnLT2hh3/
70S9rvc3T6D6cX+t8NCoi5UOlIKBcJPw+IHhTmzhfduxBc/3XILzNG1deSls
aAMBi4dIv2FB8XyK0zlXE+Ibb//xqOhyh5qjFHhSiuPUHP30XP3i7QHal9jK
aoQ96/qOIINyN7r20cTb9m6NM2Klo9Hl0eKmr3umDHnnJ4A/O0qlt86FVsJq
5nBI3mj3JE004a7nBdbCXOgpWVMSVcRH8oxeWRCzQlqmDrOXJzVyIOERYS4K
XqrLHFwd3GCJ6V+wMgAzIf0yfxnQ6cb12cwd98LoppoHTzl7uprMpN61b2p3
UFjmkbyB4qtDEsY+rxz7a3yqT4DK/OJ46t+GnTIc5nVzCwM6+oixmJZa86QR
eLGgbrDo5RUtiB3L4gMtTBJrmja9zK0z8jQuE0V3kCwOWlrdRQI4jJDCQEwr
yjF3N7Ik2Gl0dncPJZrxPsopa8UVRJDe5LjU10PwnvJmVrNqNBFs9gx9KNfv
HRP6TjnFRIwOeQ2Hlz3wbPI8xsuGRgFbAVvtTZ6aUnIp88GH7BEQBLNxph4M
MoD2Px3Nv6orbIPJGE+OXVboAlcNtetI/zBBQtCqlHhJrVOMP17RtmPdYkCn
3DCNYnwOXYQN/3T2dJ2RKfDwMhdE68Y33XgwBPkEOd7BroQOc3oLmX/k2rWR
HPNTJ6F7NyTdUhFzd3KeBOTU0Trq9+5myq6CeY0TT9hFtNSIVdZvzNdgMsCe
obC3vMdoPJKFlwFbouTKWr9ISkfnHqc6Jn64QIDftjxe3sb3KCFxgwGuRmZY
VaukmoZeyLeuwoDt+6sSy9SYvhYyCeC6ecs8BUuiMJay4vhHs37YodkUs4EI
Qr5g+4QorZu6gnk++Z8cW2wXIQt68vhRUTVIU7gmZUvO8HVHub+1N81eacPg
lvwVbxezHkcE/cmLyZvzbclj0JAraeMQEhRV0uHWHU0068czJ9US6aTILkeL
P12RKR2urZ1M9zb+Jf75uWS/oeFZXDO5TQO5U5+YKyYVbZlwwxPcYG1b1mnj
BLIXgJ1fFwxvLQFNapcOjwxBVXgN3QUeinGaCdHQKN1U4Y1UpIb8HR6Z9JTa
U74i0XXvi/7m+yP5TQrQ7vDiUc+3O8RXkYLfRDTmpBC8xrLJDDGlv+xuvOej
Ien+NRcjc+RMDFf/rat8uwohqSBmb8kybIoqDPhl5zX8Epxn2nGl6Ytjzb/2
H+oGXcnfMPsOwz3CZrYtl6ZAI0XXxlFvM7xBkimV9SZlK+T4XRTKjp0NTAOi
Ol62hjeSW0EO8Ef2GP/Z2QEnWv8gHaoM22Qtq3OXNXnSosCITGcWbGsY8DM2
q9UvZGFqZRx4sGCAj1fYjuvsP+ElL9xINz64evyAOcAmKvcfbRrPTIRsgwqy
FpwON3D6+2mxMCEUktk4corIZMypIv9wNHJKkgt6g1lZZV7RZ/ziWsPkHHyM
KRqaKBEEFXn99xbuCFUeJ1t5T5hFrvggOhUBV0XOecLOGYuTSQmh2uBpQzEQ
YLJiMqaz1zyKWZ5MtBwUGud68Mra/dA1FlprJQfVd78mgbGPi2+MgKPPz5FT
H2eWyvkODJdF4agB1Bfe7ZlL8mpkIErjXhoJJzrwY0QXNLtnwIUdmi94v/1r
Oazl2tVmlog3TgCqqNOIuEn+wa28xSP9V7hqn/sanV8trVrmrgqhCEEXzTFK
qtLhg8uCXKF4Gt5KfwiKCQNJHUZmAeoJYHAh9FZNU7ILGzHC+p265ocp+H4g
pGlCKVJrueMOAnRjLXU+miQ/KqrVpJtvVe8zFIHG9tV5DImF+RWHtIkZ6kyZ
I8tyd47q3B409iiCsznfFJK2z1sv9mTWxhYFCbUuXk+fHvF7FFWb81UbPcYz
b8VYCOePeTa7WDo+5bgF2ejtsje8YdGu3bJzhj+53KC4QnnnhBnz2BrhTrrV
KvnrAcGGjwkytYpJXzCYe1zu/8ydphMqn04svfYpg6pNznpw6cM6mxirEuqB
8ZGB+cwIU7xcpGuVam4xQld7XYBpzdy6l2nVUe9N0RommwihSjqgTokSUSDK
4/XMMZnU8FkeIJx0fUqkcI+Rn66JcKzQ3NwNRtrX0d0PEmvn0ecMbekq3Fb6
kneOQ7iURhI9d1QEq6d3mxDSyy63jVbSH7U7t5zf4Whav+6cW+Gz0GNaXrMD
cjDySSyCG3pdT6FMhz9lmG9F8PTz2u/LZWd7HgcqdOB0FGw1npft0oSP+FLk
MggZiIIBOMLLbFXaSWxGRSMCs+olmNoMM/446oQDP8+2sw5p6Quu3xpWUKLF
l1B+v9HpdiXISnBQdXv5S0Ze7RgPOMm9XQr8dsqpGmioQFp8r3RcWxzsGKbl
bUrLPEm8ZPOIElR6Jid+OVijSLm4UuubzaCL5ACAI62Ujs6xnl4NDsIoYPSs
6G5f1HHcv3AZhqdYGquK3nKqv8Q2OcB79vLOTUeM2dMzUxUCWgXbmISbLr7g
mC7ijCDKOxSeTItJ0TlVrHR/0Tz1jvGNTGs5UySaTXx+5QpbnFU9qxLyuyhP
KA/E+xzsCj4Gc0uDf09fpur706nzL7ewqSilNNOJZqZAnWRHesDlN7DTAHw6
dhYk9Nq+WhtzQSdNnbB2Hx2i9LavRg5d5SZElUkIRzf7rEjSkjIdgEDWsuIh
qc0l5EsWncKEeV3zxbUc7ej3Qt5D7zwFEsz2RsedFTLqtAy1i6e/eJ6B8vEt
mqD83i5BMUPiOkvOvsjCN5zSiJAh8cRUxu+FeHZ7oAW6jHnmcLIqfeBJTFnl
gqPJDc9fbY5dMs2ix638OevUIwrRbtbX7EaYz8MivFXZgvADUwZo382CFACB
D5nPkjDgAmSIrlN7Eu/8Dl2BG0bhloPMCbdi8w+i8ln/go3E2G3VkoWyJ1yf
/fTw0odwNbwsyVCl5sUUxprB2U+ej2E+OP/Vk/t3Up9sJGU8HvdpgB1FNE3O
CLy2ZufyhGtBFOyDGZoceYcyy3gJHdGJLqbOLo6Q3OmqQxYkI/bu8fJq4iXG
1QikgFW7hL0l8oKOHYa0suxnU3rbRAkmCVjI7bSuo2FcN66v/HMyoZdJw/Wo
EwfOIuixWw81GkTLMTX4wObh9QqQYR+FuS417u0HAv5hDJKu3LKvkt26k9Vo
zaA4D6+pbF+npRtl4Q/F/ZQpH/YYYSzb74y02+H0vh0j6liI5YuR/rg/HKlT
bXSZk6UvPFrYDKolzwo+XZ023f6btVtPUOEqXtfu3b0hqdS9vln2gbk/E2W5
nx5momXNb1LOtpcjEfg7GEGVCXN0c4Pfob2ZqVr4X94acN3M8G01q+FFdlxl
rU2BzHP1nYFxwpM0fSCsgeGPZdjt9yzDSB88vcMUNtXIid2tiUKQDodFYI4d
sBDraln/YZot0NGHKT5rifYKMNTr+ra4imA5yo2eBpmtKrEyHMLwvgfVY7re
pEztGuxnwoYLu2SoSv3Xu6Or57cCPsfcO8GyyzfTiXSTejxl0zEJGleaEfWr
5DOWNPjws+KYZ6MJCcyidaZWyuK2Y7R74UTq1pYNW6Wo4euP8Tc6FcK4u6QK
mV0iMxfahx9sG3oHr5/mymk/+EnoJePHNWwxPgdhfBWRXOsd2rTxEN3pP5W5
pel7h98uXkXWskKzWTtztbxD0WFC5jNKODKEXkDnFrl4Llb48W/4tZTHOkTd
clNxf7ALdklwVNSXeyo0MjRlOGkqBxgr67/DLaIPDgfREm55XZ9DSM9WR2BT
2hfGHDpfBX7hksgG34zLJfclkoG6cnahSDRcBIY/RnmPPhiU+BJJtcwI115R
0ABA0Aq3K6/crs7VvCq094MsL7+AYfYAx/0t+dMi9IyV4/sVdNM1KULWXWyM
8hh0pXtTluiS4NPbbxFQ8egvOtzUOUaM4ueGV+vmWC7s4moEXx86aV1yyv9X
DjYnecRbZJKFC0up28b5UhWUo5EyBWa+6oXDXD9k1Xt0woBJBR1KHPuuD0ad
7fcpss37aXM8DSvAIjzOS79Mf4Q9VMreTsHjbJH6oyvYlpO7azT0raDPbrHw
HMa3L0JlwCwoKclsK/CJQbdBI3Ouiagos54R+f3FMJ1tM6D+A6SnbJHGSTMM
omQBvpqvRxSB/ZC2Rj45U0Ua545c3wkuojQRl30cfHfI3Up8CFc32j5cJKfq
JHbQfLDFCjajd/yAHHeP3SiElYT0t0uxC3kpxP1phWSVOzn2KIewQXKsJEvb
MYC7hRxAA3MpZxEz3p/fHwfQXwANkhYgtS1rkNXxfr06agjzIaeFfv9is5BQ
wURRKxnHY1k1XYdBwnHBPYYbLVAFKBJyY3vGKPMxqXP0yQP4PYP2UuETovbp
pf7EziPpfViAdW/mxJFyoNFSXL8USCLOkqJxRz4sOJ5I9Q3+CmXZM3nZqeoU
gXX45STAlHPSafTGfTgYS6zwXBEGRYqfNuECggGRJ9SwOCiUaoPY5Db7PFCt
biMxI0rUlkgnn5CNs6rp4PuzPEmVbw1f8w5ev+uWrlhlHfp2xyWjklDkPNc6
b9aRK83RHZlHFyCJzvoFryc1dJDvukhuawS0nO5Rsr0ytVj3C22jF0oUDRGN
N2qfP+0S6ojglH9qIrpOLJdU0+DWT2zzlo7nvLEXASZGQ8PVcaGSrH1SJmGe
VzV5DtLeUV7E05UzLuzAXBqnsQe3nfQdxeyBRIME+F0Ckv654uQcpVVA/nEQ
a++ZS8VMXBMyOS4O1Y+thZJxmds7yfid3AdQPeOD6Q216LCNy4xs+Gw5U2oO
gma/NXpgyuh8TTQHY5gui8QJw8sBzohzsoXuQk9/3yz1Im+D+FxkyV8B6H4t
MRpHXT8q/8ylLIgmeWfu8ExJxZ7/V2nTwNQH1CcvQVgEQYERuklV7pNxRY4f
Wx2hlwQ61CJgIVlc1W41oNmQ6NYnEITjTycXxc12Cujw58plfjFJatKFuAfx
iWrFCBe471qc7Fh8aaRONdBTYfFm8XwIVsUA2xOlPHgjKTqJ8fmlj/VeSAU7
CjvNj8w5uBhjrySHCfor3GdeHGv400wN7dpkZqWyFo09u8mASfCUTGQdb4C9
EwgA8f4Y5K7VEoFh1G738ebGbCe1sY+X8wbXnJcD7jyhT8B1fc/FBo4Xh8GY
A40jWIWIWZ3MHj8Fxh+8kwAQnvdzZtp1tPCn/ry4LLrHZzNTWcPIALdIP52G
lPHa0qxmweU+eQxtLc4oLUelcmTv65Wcy/e8P7dK7gkEBxoja77LZxKrCaXm
Can68lA06Q9JhLo05d5L4b7l/4drGB9S8wGZATTdiBpttvsP5aXLlAgZaiS2
/l3mXCrTtelFcheM36bOdNEqoDLU3f4RHOVXz7XwDyllqy+ER8bfj6YGQDrw
Q0juf2f4lmigWJy7yweLWqSuh+eWC0q825HEWdtRjj/bT+4Ci1pYVHB6Airk
431nvVZdK4b+Rr2hVFNqRu0B1m26HNG/bvdIatSxib5PHyQ0U5GWLEaXoLIJ
LNYy+r8QtLH+Sj8do4KEeplRUNY+fZr6FQ9a4Cx2tO4nZWvTPSiXwPxpn2I9
8RCpW5ZcjQTrkvvE3H/9FPy8ht6bygWeWT5vy0ovypFxzg6cR2M/DskMTEB+
eHYqAzDEa90fVr3D6a6XrdOkia4ZtIojLsyNMF/wTONBhBf01sPZwDm8Cd55
LhESGsW15BzT9Hlc45o9FaFVEWLDq0QzRyCp0QLaNfYTqKlKV54RFRtjO8EL
CsHuCiGIPXhXCDkpAovYvO+7qyGnkbE5yFyMxBhWRt5jKBEZDDPi6Jxcg28s
sgbYcrmL6AurFxB37PImfksrlSoXLZVxb/K811KGEwdWgpqHs1l6G9L+VJzM
HljTNEpGxMNJ/f9/+IWiHjEcXohhHV2Wq7GhXq/yoF4zfvd9DR4Hbqy/LYQH
UazzWxG12KjTQtBV5ckmqTRu2/HGBGv7Qh0D7CuWXIxeJjZMFkm2DJXqvp84
uWFk68Qy2d0AcFdkyjFJ6e+VuzboP/dl+ztNZ0XRga3zpH735zaX91Xiv5dz
GTKzYirQ06YvznY9ghjpIOvNYBFt1jI8d8ijdvxvczGHdxwLfTexLHv63ZGM
KeRCsJ1bDlnuPqFZ695PM6AOwb1SFPxnhZKIbDBNJJI0+qqheqlh8WB11dJl
ebTHo9ESiE90UO51xLbHrkDuCqOveKwGrek6Z8rT3mriHQBc5H3wXjBn1gS6
SYx7MFcFvyAFp2OWXqHVLzT6TMkDtXYj00XP0isKFQRKOS8tkV3rY52887q3
m72exVCZ6HJQhyCZNp8hhDJ67QkM8d4YRJ8lRNZ3wpnNPZ7ZRY6WWpaCkYzp
mbmVNP0zbWMO18wJIiSzNFMkCP1mH2XyJ+hcY8vgPK2cv5Nm6Bj4S6uoqA4+
l9STT+xug4yC92cgiSO/3XohfGrTTVHl1nHhVXWImolWEDuKkJd0p7K3APO6
Y+wJqSCaCC2X/0v7QJYDuOHiTxvXsCo9J/6wfUEYHOGvD99zyb4+LT1xSZi2
FQEuX/lNd10yrqny9lzc2mMFWwbIwmzrRaO0pcabh0g9hVxBGsatYAtHM3Xm
hDT2QaglS/aD285rzHjsgOmbm7Z/JfaH1mfyZBY2ea0nMSOoy0NcHftbp5Ck
Ji7azz5ak6TXIQkrfIHKN7s+vblHzC08gFptcg6bypg63e/nlbkPKZD023KW
+1dayeQBVkQdxf+J7aW0YnEiGBPANZZN7KdiEkXo/bD3O/I9xLRxLg75mqHD
T3grLaZvgk6d9le79eREfQHff7S38DPcXMaBrq+RBAp8DdyKbw0ROUOb3lZs
nDxvm60BIJCwxlME1KrKAzNDHU/s8H1F85p1EoF+qxkyJVQom42MNPn+H0Ks
HaqJRMtKoEsitFHSPPh138fIkRVS2xZSFdJ8lUMaagtqCHSl34NwkIVXjs/v
aCoI4YgqS1VxAX7Zd4+zILXlh36kif8oERSFnTjPVyjtbXA9gyMQYRyCbAv/
7Ww29klI+M2p72ICN3wSbtItQGk9ZgZGsupMipby4rPwU4aHM0Z0j8jmRxN3
tg6BEgu/5L7FctG+PpCbzZN5+aovo9wBwUlWwyN6u1hUlVAX/dJdx/3N9bD5
wByCmIVvUo6ovaSnN0xQXzr59fle6YHFARGKQPjo9Q9h0XnMlKjCFf03XoAF
gZWWPst48DpA2r6May2kdlF3gzA4FvZoW+4+GLswApmCT1ysNeODfBwiB1Gk
l742X2YCLATMPbbK8FwCUC2h2+aHRPVW0t03elQiItThOGcuYy91ZyqO60Eb
eN/x1Ng8Ds6sK8Ze69EH/n7So1EBw4dHVgT6lX6nLLW+Pwi5cIcaFV/YHSCv
ySfyfJ0wJCD9s0wpugoYPDOHAha1H6+oNqDPNc0GX5rj+Na+dKL9D4ZVPDXe
lUXzFw4uiB/fmKTOvT/bEJKZXU5Xl3rK+5cz+6trUdyuJVggtV3wp40c48m/
WT7JndyryDrs9fj3LcIvaycEjNRI/HQ+FNEzpKAe9jxG4hiKf+akq9m79POH
GJNr/u7wS4uxBcxwJD8gWVdsJkrndUI5QaeSEjjzb8cHgMFYpOIhoTN7KLoG
UuaGMtlFfs4s8kxKyZshIekX7x90YzIrQ1npwYfHyz2X8VnTbqL3NIERrxjt
VvqkMznfDlunSz1NddLmAGChzQs9NbudYYNcm5Y4yIM0AW3OBEjzI8mVGIdm
ibpKd4pSfTBhrRcr3TLA/RXwdMWieeevUkIWNn0uWbeexehM8Vev6gWaHQeE
7eIaWZxAdMv1vdDSnbvqPKD+KRXpdukWuh5dmTTq/6U4+EXn6dii0G7E4Zpq
Rfa9+XilN+ktTOcjvSuftqUblZ0YrEkW50oI6HU5bmd+51Jjek2j+OJpnv8L
22h0AvOLfkWH3zasiRkn7nFYABcpltFvtScnA3jO+G5YA6/0XoAMr+KaLzvM
QUa9qHpirtrOGVKzyXpc8TC7awZS/WlNIhHuNjwQvYotQ1uFNhFwKtt15uTN
0B2ilO6J3RO4gcKkmiPUjXS/4wm/iJkvT46ay39G1eXvRZjJL05EYo8VZVhT
j1Vaq0YVH7uJRic45uldmTpC8CPz0Yi6CcTPxo6uHB//VXXr7ECnvkI4a4Hv
zSrJ5S+W0ZJyiybdwvr14cgLpklGGBhbe/44lvyzIWOQGhoqMuAtjfDX3q1/
kAjxq4Q/kDbG5E93qbBcCgXacTrH0qJMnU0+wAQGqOIxDqKP7LWUxU8c0hIm
KQ+/7e0XtCNVZI2mi9pwnDDiwd7vQNcSpE5yI3JMKCcyvM1a9kL1sa81myWq
wxNY7FRrnZc2wxAcZs9BvLr8jYZaXa3/ZzuUDZC8iCtWNkktA5Gi9pBOWcF0
n7ALGRk8wWJEBhrOoAUiI7ezeARR1yu7i9mG2Jp6GMil/VfuV3Xd5NBYdAwG
ghJYEg6gpTUW1ylFZ3Ib+sdlp0us9g8DJzntMvHpGbQQusySCJsqfHxctP0Z
QOdtPD7Kuge+VtibgU95LzCwHJgVWZ5TOt0MiOFPMWJ3ckn1ARnvyLZo4ppN
RQNenHfyAE8RC+0z2q4noLx6s2if6493oQigDyBSeG/l6PeaqfIS5HRX7n5d
tyJYhwrShHXaq8cVuoxFef5ni20IVrAcaBqJah/X1p7IbFGw1j4ga2GXShsA
d899htGB2AeKgjsd34QX+qb6F2TYk67eTTWkPrTJcdY+AWUPNTq2rNLG3/js
VYlaLT3uRF8ZUqfuh7z9NBWWem2h6qTCwNGmcs+/ubDkEtn0/dUnE4ht/2xk
Nk5FGQSkb/53COajfUGOgJmOl7GmXpXidbiULVYXm7/zpWiVs3Tav2RtkOxP
y6mqCZjasAb9C8DluUQLPCmmHXkFwmJjqUlLO+RLB/WZ+7x4hDyikBowIuyF
zLhJwbqNfiSHmD33nmdTDB193CT28crjIvp2fpMWXJIVRB8V1f7Rb9CvJ4Kh
t9E2RhwYE7aebyUR6Zgl9/2Hzu/WoBy6Tbifd7RYVFvHInpm8XEhlirE/oG0
fiejnv+BMmjqN77CbV9L4ZTo/h+Drd2PVOQhePKyuhFAgFPTcPZH1tBhj9Ki
VUUa15QKRYh92QR5CrBhhfxGgIcpgzcVrykvjE2xJFehmCVh/yapQCnsb8l4
BGLcCxktl042TVTnpNOY0UUrL4WnsIVA1jcOnswo4Kh4wTpRw/Aele+q+jbJ
EpywUAj8QKYfK5CxGDyJCp2RXxr7LWrAUByYVVCrTpcJgPqoaiZM/hcLSemV
4o9rqkiREA6DG5+LRKKw71wfddZvApS1GOhiwqie9PBm30DVNMD5u6FsgIzl
ZLZsohe2sc1ulrwRPvMDVir0HjUlk0Pr0K3ug1Wht5eX/JBEj53Y6S/EuU1L
vgGxnIRg9BFK8ADQKYUPFAgmNg83mx4urSEJTowgwfYoi2q4mN+xbDQzANnb
7c36k9klYNiD3BnOJezDzP9q7+Th9GHqc3hsOYbzE+pZ3BpVNEu1CHhw2Wbq
oUjQWscK+CsND0CTOZGIoz/kSgLyXbtG1L6yiHW+gC6aumXStls0te30E6FK
V69QIWbPHPOrNXzValm77uH99vKP12rXyDAi4I8JjDGInwn7JYZaD6+T20Tw
LH9dKx3FDXam4tgFhjOaR//yzA5Y4Q9pqfLI3Ji7sGNFiGmyNZhrGc+hmsiL
4lndUAZrPnZvgtu0wcfnHAyNP2Q0lOq1LI0mDIKfumAKZYAEWvi8ZUQL6B1C
he8iLttRxAD1NM5+o0Fp3o+kf1SYy8UF7NR4N9lyT71ZLMy0ZGZhNzu4MGCu
YXgCl/RXaSTKgmGdPbY+YdsnLmXKndTYJd3ydhn6empSOSa07Qlie1k5LzYU
oFd6Do4KljhSjTt7YqYDamQzVlYM4Q/b3SQRDoh06tdWUCTlm09S0HpMP3cK
nJWY5UPFG73tU9sjzouFARtxK1hht9n8tnQG0VoYqs3oOKyDC2sgCFlpBC9M
I4SbEICnaHYRk9Js57idAQG5rLGTjrWrwFgPANIj2MmX3htnO4sdfGMpJlEp
Lh/rk0UhVBsbwIgwupxasuhjyoRxoo5mwBmOWn1f5Kwutx+pJsCO3eIJSq2E
1tOExXGf5gO1K4XD9kPl6gngoNg1X+oXJB/N3BcmlqdF/I8nAV97DT3LlbpB
4YGE2cP4+ZCv68MEHkvdmUCInpS1NiuLaDMUWhpDcEMfu4/DAWk+evuOfTup
6+BpxeOH4KTmWSwC0QC7IazwzOSLK1IYq8PKEMF82qnYDiVb4ZUgayfzI4rC
sMdLSf/BwDmS6sAX3wu5pxmFeL+DAXCqLTyKICSIx41eKDjnTov2Nmn8uNvE
cmVBk+aZ2w15hFsmbP1MNG9/oV5ducXEb5ca1BXM1w9bPknNVp+/z6zgT430
/ef1Rk4a0nXjUuri0rvm4h2ayh+quQDQ/uAbPh7RXJYIQy8+dGTZY4jILw17
R2pVcVsQYUeMQH6w7O2+tmH3KcaLNsV7hiLvI2iThAPXItmhml4Ee03wZGIJ
8E2++YSxxOyHX5z+7ENFo9Tc9vYi9FLdlK0nGwZv33wEYyrEru8IzsY5cIQC
vCv6cMBa/lPfnKAdidQZ4E7oPL5+r+agn8o7VuxipYRiOtOlYVRugESPj/3K
HQwQxkU3l995hR8c+e/vWOp7j9SRGwoX9tfQ62a15dBaHpJSbF6EGkubXOI0
Ibu+QBGLaT8ihEz/tZ60n6cGIQA+Vk6I/fMOtY4OPX44nAWBXbaDE6s3EDO2
GTCu/O3UdO9G4hAbf5HN+b8H38hxsMxREyr5HcM/a9ReoXmpoWrBHNuA+mqA
LCGFcYe5biUkpzGZW8xovpug+feQoHtJZmFh+KEv8kQTe2tWuWdmx7hklO65
4nq5j4JH4wWEEVQvAr/7T8RyGJLj3kxN9cZiNbjRXKmWLXErQZw0Yg5Aavgp
XhUhbJdA27+19P5kljiagPLcRlzsT/eDyfWP1nZHwHRqyu35J3deiv2kwCxq
IXvCvnbs4HZyjOY1pphVfc/uktNBVqV1QL1Ch+oiMKjJIAxf+TFDtq39n89E
vHwKqKy4IAdqo6BvymKDGwtAijkiLCKbyM8jtz/ep522Go6Jq+2BS1ubpvMi
+TOCt6u1Z4hkVjBE7gcRpqVBWmYle92blVGbbKwIVctjDJPdmvrdSVZ/dBF0
Nis6yXsZkuEOseLpEyCr2paYG23aVWxorhx5IuA8CzxiY6D9iQa5s4qixlso
l5C4paU2YpRzuPG3TP0DNappICG98pgckrpLb8ZGwBKX8BkKlAIuScoXiFNL
UVSrmamIIY18lZJzdbwFIyuz7YJH+oJ2YSPhLFPMg1tMAfEDPIfK81OWL7vi
IRz3ebFpuOa9SLwJGARyB1hdXLkdx8NoPrzvcKkHY/FeHHVxyRBBndHQcuTZ
nWBoUQXk7rmMt02c0NT8N+O2d3x1cPagd3T6X9BfoXS6Lh8IFe62okRQC6Zt
maZY/WeNKNcjtR7S1XvJSAVm6A4qZ+Xw8Sjwk0e6YmD3kwDnj910wzt+VHcr
XIlnqxK4kLRqWZBVYc/VEiFEfwGfr0ZYi6gejpTlQJs4uRO9+9Ay91wOHnWo
hTPW+EIRmIB7Izb9f490XNirSZZIXKVAm/SIq1tz4Sqw732q5J6I/f0M8X/k
MxoykJLZfzRLnmTXi3lOzGVvABgkGKJH4aEA5jxh1kHgKzKPlOnJ8eGYEN1f
nNwtJAH+HtuwnwFeGEODVgv5cskoqbkp4JfoWlLbrqQ+yqBIKovAgUfAak2U
WGJkgHeGdqWu85Rbgm6jelW6pW543/De3GTk70ahex+U9OD73jIUNcEOJEpn
+oGP+5df4+gu4v0CspWHux57MzrKePORo0g+iJ8oE/FR9fVHsG1m6E+xqtol
b17XBTKQXNutYdq2qioDpqU3y4JeBgVJ6sfu3l+PwtVvoNlM3x275Zsf5R52
uQK9rClYMi2T5pdm6HbFUInozn9SLi4/0yvZ6mdJcnsuXwvkyGRwkhbrW7t+
6Kdf8ctjeawtLtHQ7H9UC4tn3yaONQBPxmqxk1zZ8s4sj3BZfitwgMhTiaPT
QTlZwKngpg44lHPSR4bmafpUQg20Hs+rYZ72NwbEv1ptJ8frl3dxxLVaO09F
Htr7AHw+NMf/IgMZFLvHzy/uWhwyUGVhPnvo6T6QOplN9HHIfpZA41Riovwl
b3fmYLF3X2hVMYbeDGxsFScRbf3Zjf3Wg6xfX2LKKAJc4NzxrkKX1UhFkpAy
EY66WXSfWW7HRfFdob9V4s4Ny1CvVGYfinX7Q9pdcr74+kqBlYDRSZrghQOp
0HqNHAmMJANBgNeZMpsYeyMqM568j87SWfl/FrfBs0pTyZGzXc6iLapwEtlr
ZhqvxlUP0jVWoojD12NxNnFvygX+KxdoKej8CnPThMlqPx1RRvC6JJjwq8H8
HexqWcQh0PcDJQCDgeCb07MnKrEQjJJ/HMW2O+85b5aF+z2R88sLQ1Ec2OOC
YS+WlGZq+mKkZHF+pfmG2m9vmv8Snr1oqKwodo3F2AwhITKPZd/OD/TSD1w2
OomXBvJMb8XF1H0yAe+k6SDb1kxO07hwbmlYFjlmWGAUyQxu9abvjMnAzX0y
VdudR07bPz6oupOHjUkY/DBWdC9Iz7JxHvsBcjYZi2EEQKlNaxas5vGP1/xk
fCq/q46e+Gg5RZOJvSWVOb6LhOagCuii3abjzV/c4Z+kOrxgcE9Ge0lbqxHK
UrmddVX6YO0+3YgvwOmc16Vzkj30XL5IIvF0JdkYg8uwl5YQ4paD3wbiZdK1
bSLHjI3lCScIZezWTpAJUPZH0SL5bmeBxb3sgAd3iit8ZS3CIAQIVxBlzw/p
YHQUZ6c/3o9zt4lyyeRWq4rHjhsYO7TFQchgA6F3BIXBrRhp88f2EGJ2zkLL
hmDX3Pgay7oOm0asFpv2BW0zlVvt0znMle7vqUlvnct5RVI8G8z+zMkit1G9
PbvwuR281BwbGLEh1u6IS7KFEG8jx5swGoTAafDm8xryNWyCZOgDH6vaTyK4
xCijcGhHETL3GYa7cLpnEqXSrcgpplfI+VIWHNO8HkRASy/+pifXx8J6hsLL
s1OiV4RG8hTH2yjZH4NatVj3Ss9+CcLsH9G0zadcAfW5/hmG+eziupsIEGWA
lFmLj7Lduoznijk7j9PcE800IiqWPmlzUHuUXZj8j4Hj4XsCf/xdxnNk/Xk9
cp3k7j05Bphl3/8ZzhUObGQ83Wxr7Bzgjkf6aGbY+mBPFX3YqW9foKhjp+yo
qbZfwI2gRYcWbnpCuYipn73IIOKJJGA1f6IQSm28ocl/hYMst4vGX4/KERwx
4AdlmNyQdWDvUlMtwEaQJpQqIM7iIZVUj+AyT0Wqm8Qb0xTeHhX/9v5HSwyn
YK+HFooYtKU7bamLHPIixJuNc8GT9ZH18ypTA16M3PzUqWpr8JNNY/X3XxFZ
g63Xvgda4w5LKadhJBNsSgybFs+S+9WLk+h46BVykN+8KDb/7k1AEv/oOvz+
2GJn0zJJd5JkPOd51xbOZILHFwG3u+UvgkCIk+LCdCd6hZFs5pSLYddkduuE
oHyunPu7z1r9/tSlUSvyIJtvMJiPeyF071auLVHm4FaWJD9N8gFgxV8WwBW+
o/GygMFLWXToo3CIbfYESl0KQjZKcGyvEaWQjcQAYWpvwWXPyP7rK663pQQn
0dPeTPw3hSwluqk1UWcB5A/2A/POE10wEEIvSywG0j/8hPieblLFx3aX/udi
pUY3mu5fxJJ4CSISVfSU+UCJZxtzTc0UpR0pfXxbyz251ACbdHITWreay/Sf
3lu6auGh/XuLN6TTL2Yy8ItaKlm9yHJ4qXrJJOYRVQo2Jd1sTrfbA3eqO5UA
74IBkfWr/DxMo5ewTqHzwZ+EQUrjTgyBPQrWv/VFUes1XVzut0lluMeZACMT
K9XY6z1BZ9VTPrfucHcEJZHzwLZEpFG/igiNMhrOlp22JEJToj2slq7j1lfG
nzCQQ9BEVVtDenDUqQc7ZFONvZ1OuwA4BYSZSjqy20kD2r040QuCz1x5C6Ge
hABHcyhFi2tXd1f7zGv1NTv9n0AEsK6OeCDv5NjQHqfMpdiu4IX7ILNJN/F7
mrLzbyvM/W4L9ub9bi4ODIc6QuwOFELzzoaYRrFFDfRJiv3f5TgmxO4QCF8+
7ooxR1mBPuH3aInGuo3EUvOKGTD5TXiFnp/7ZS8hWk6reRsRKnj6GA4hvlQo
5pQRqg/OBSis4G/frXduUdGzgTlxaMQt7sOvYFxGuqGLdVJfb7KN/ei3p2WG
4yybHAUnOJLxNj6yIdZqeJ/tjI7REpmdaHnkn1/oy3/+PJRMMqEBSek6CmEm
lxsA711QvlKnkkyViqQJ4k6SzYpzCivcriciyoDqAqr5rE9IKWkNdH6CmoR+
EFXx2/we1G+3MuotERgmJnSRy9Ri2mkmrCHM8VkKdL6py6YgPRQJn2INO7sA
xoK/usufW+jy7zzSB4DxL+qlDf4T7yvfpUBBHo80qtK0oxAsg0TwG4qcNGzV
AgDwQMaAYyk7TnrgUqRLYMFULL2UWbHqx84o2psfDUWgza9MUBb+oBNxURwC
wv7Z5QDmzJZvLBKMlZ+0ZIfQRrUumRUWvJdoq6mmzkdIJ8LglWQMbdmbbs5T
vZuTeziRaHvl8F/aEmYHYVO+LiOV9O7v60tsKE3tJlBePHXeftO9gWzOnDYT
NAK6ncdddIRmfJPuj0QFiyZAWpFxmSKTnducrEo8HX6UahSoy/7aDurhMrlr
gVkT3TsumVrOHle4NPzYG4fUMMoo4I6E1tvg06AvVG11/2kzNB5iSY6waBwe
jGeSD3jauoddyrqHrYTs5vRK8D1PGnFgS6Zfn053hvCBLCeX83PIFTsYDMCP
fJ60z/0ymMWCuLk487PG+x1fEr36/p3sSK8PyuFn5oQIh3CYo/N0cr4cWoOB
UZOErJjbS7GAwV6LowLFPpNdo6iVmduq8yyH/SO6zFIMkv/KUeIw9vOt4B1D
KTU3vJ8Qg/YJpvi0+IwfavFCpoPQ+LyKNNuC3xI2bINvm1se7d3kuSUFSvx8
bmzKjsRtaP4R0npY6tknwYhC5USKzRUoZdD/j0YGNsHOPBtkhV98efkMQAqG
jbbCvjaU82gN6g90z8eqazrcr2h58GnFiAoHBGFDsRAYabEO1b10JRqppsjs
7r0GXZ1H+aWFWgnRk1efURkEF16+Vx4CZvq0ShcmImVdonp9VRktGxLQoyus
6iXcaxYyxDLJ0uFDJJjeBwom/06+/4CPxBbftykYZz+K0Tw1MDnLctKY2yuB
vuktZLyrNrikC9xisjZBXlmeKVIIFytTwecs9fQS4AwlYb0M03pfOHpeVpdh
yvtos66M0diymcjHszwurMsW08wTNU7DNnrsnQItM+wL6zH7KSV6Vp6JQn+t
mqKt/JGelKcsJ3/WH532QExbhfbIkiOC4duIBy3JgN6h5iTYaiWFbPT/QubO
Dojd2wVCo+yfD2ZBukuzsApK3dasx3fgwqN3gXzhU+F6qDQz+1uSxW9AoWqA
OtFiCz170T57Q5T51qMzY6HXtQHt2AY1Cq3RM+OBdlyq/adXSBp2ucMISYlQ
lY8U0fh+/MADrSnlMIwlRvw1Av9K0LPD+Nz/egbE0EeEKoQnpZbD/8LlNoUO
u960no7wlDryxkdSPXHNm6YjTde+LCGvS0/eDyynVJp+y4K/GvJkyZSZMCmR
DrZM77ekiAVgXc7MRAAW6DcFeGU8qTgyr7XnjEBn0GSbaF+eP1yFVMNSjETR
+vyfXbheCOLBjZzBDq04idWiq+O4KzmkCnSd2rsyGElmcYKFNALwhsF/kw0d
GBLPvgsMjOMGRHF/RRZJd6ep8klue96VGdSMyimyZ3Gw3qk3jQIF/6mfEDht
7m6ddK11HhKAsX9D0l4diyZoO6AKBk0QmGKui0Rsy4H6UoFtPJFir3J36/gl
jzMhq2MdSg66CB2k6fXC0jDPCYwEUPRfCxBvG+XzI7ikQhY7DrZhNgSsmoKn
kNCU7YyUZTef9joc/iTo2fK823ZsG9RpMPySuv4apIr85x7Ve9US+yJZM6+7
u0eyWLnt//1gMjmdAdie2r8RKVsv7VtCa2RnGqw05xVtNr/RbKT0t8XLaLb1
+IaDTAcn76h0TdXgLjfElcRgEWGX36JcN+kzL7eXo/t9ekvZ1oNcw4SCxaGO
ECmJPdxx478OkKJx52PZWORW9HtijOVqQy7451xLsEnx0XWgfvowEP2H0SYf
AXIQryLjMxfXC7K81nPdebXHiDEQERqGDNgEwfe1FqqJIoC47/JxLkmX8RCv
tpqfcX4gxAQZYxHYKKKbDJadkRpB4lsvxvqGSE1EiQRxJHnzyY5V98WxsbXj
4x3xFNkmJhcmTfbjCmKgnik+r9GdvvQOee/2lTvIchz6lkCVDPX75ydECTf7
+ED2pgIEzPufsVKBtBYVBhz4ZRMtHGXCTBV+4S6Fjdm1en8dWzJAtlPlyLHt
wwleLJtes3Lb2ZNwoyksdCIDOFE4gfDAItqKMEtlHhC8yr6SnE8VxAOCKuZ0
kovKZLbekd0RpPz8zPiz1TLBrl9mowZSHPSKjuAusidH/uPLtZO7EA9W90cQ
9DRTeTTXFBfTZxD4xTl5cyj8MdhVwyGLkW+ejJvQv+ZJ03VCBJpvhQEymTm0
L14EqHaVZDxmKRtbsSXwhWAqj1c7CUfxjDmjAdMxCMZ3AG/No6ehACyXoyWq
eB7v6eBE8wChxKg5Q8p8UVDdxETQ8wmbEKV/+EcxIh/HMeJQ5c39bzh14+Xz
9uTCsc4SaHQkv8D0G7ANnUkA5FYAG5dj0G5aquyM0K8hbwJpxHrE+FRgKqtT
qUiiNz8/oNZP2GbqdSRbVWqVJIWHG7MhaimV5MIdU+FG//pYkI9NZ9Tf9UKa
8z1VT5bYiY7ihaKSpLO5Is6faE8NkYscOwMD0sqsXvTG9ixcI8Jncgc8cdz9
049YIamdmlMcsTZDtDMpjiilVgNBOcABXO7Y1TDAFualxLiYd+zsNJ4YIZLU
1DDdqTzW61wghKxyElLc/pTseLdFzncXSacVKnGgi/v26+5W0PYV10PKmeou
EiLxYs/+fbh5nKWGjChJPoWYvig7LRSE4LkxkZr4iIf/ddAwL7hQAQ+kKxkC
1Ioaiz6HNYqN5UEggQzEFKkmSPDYWA2IHmw05Nr3cqE3hnCelYlxFsbW0FfK
xQSR9nRfOXd02uBfRzpfysw9wlZEfhU0cifjccruW9l9xdXu8WfD64Z8e4o7
kgOyT+2IljF2gqatDY22NmmzlZYUV2yRoDccdxamceuDIKbDGSXS8i++5J0M
3dB/FfZG2g38OBheUYASrK/yGJ/Ql7OcsSyG/uLs61xN47pqxLXwyM/iwTEs
671KEgzSw4w6ZnC9VYfyjw80IMLmaMGrUWWNP0Lrtj7yXPeFST9RR0opmi0F
BxyW/xV+T3oetruAdUm4x/XA7uMP0hGPAmVGdtC0kOmLmPpRdAVXyDbdD6ZS
8DlSJ35nVmtYsPi8kDUHYneOAJpIn+pqGzrFThch7bjwAQs/GoQMor9NixFc
6Bih3zm3rmgu/hhTfgnF8czocfBknxQRcGjFdx20Cn3mfCShTLE0XEQYLagM
PBU0lRxpMUDdFHmNTJ+WasbqOPi48vyIexdahhUnMjsisv/ntILGO6b0P7vj
gFCebUj3Cy/t5nyaEz5yrfSGCGk1hgdh2nxH1N0E+2n9p65pkFdeX6SLzo3c
77nor3VFA9iozAOYgV+VtkIc+M11SeB/tnD1ThfQAyNAxbb/jYNizBb7bFSf
zb8ALx5FVz+h9hiZexs7j92LXfSWP9yk8W2N6xuyst50Y3exW90gSlWAOPrR
6pvndBH1FTsfq0EJh3GyLZMN7HNRUk+pfGJf8BvtB4xkTDJ0/Q6P6QPQDk5W
98ru/2id8FI+BHMaA4gCi1IGEEWFUmTnX25j/BBJiXf9sVrcdw9IyEowW5rf
S+dApQJI0yklcigipb5V7kTzy1tZ+l6t0PbZaEZKWZW90KE3aoYWBOS2EDcR
e3paGRCX+tq74w2Qid67ghZpA2XD6sGaTQTX2CNvh8KpF+LODABcJLCN67tE
rmd2GGr6qFuTB0oDJga0uHAJ+7/a+N2txqW8tVn2fIArWrC8uC8OcYvxy1lO
k4ibROSrzNSbOkXYjwlk7QnKk/kr8sYMXCI0a+/3FD3qla5gaYBfH1uyl5Qd
+d3LrQawSLzqXBRlVx3lW2gAGMF8QNGebZxE5qSQFE4hATiPan4DW1fJS3ih
9hBVBHP4Tk8dv//VmnvbmY1xAlb740rxwasdIAsXq7tD3182vPqKOxVL21xD
lQDpCwBu5UPFXtJChkfKAbZilbtC1SR610wyrfVRUsm+UQxwPy0kBIgrZa7O
ZVsWa/E+c6z9wILuy2T2l3My+mp/aLculo4iil/VagZhkTEtLoLiqTqzxL7a
NeQ6GkY3qPc2MM7mK/I5IjltgW4BqB9DoOGiBbYaMF4bEwhqqL87nnu9gHA8
IH1Tbq2SkAu7DeiZLPZcCJCoHo+z0Eue91AxGF3IZhGQUXcKI2sn2YGFyOPP
QL22mhZZ8lqf0C/D++ls0g0I5Trcmey0PnVhYewaH1OyJuJCp376j4HbvRQ+
WCpMcwuimXbudgiCK96CX+P509UY6jI4afJEvgg8EvAqejNmkqvM4kxwfzyO
K/hhrTNc5jy7OKU8kYKOG/C3+CjmnWP8rj1/ZmDg9TCvUdMmCdrP/T3A+5aM
KXDAtOj5UUdmFEi8kNgMAtvB0FhScZSfjnZxcZNnht2WBa3G7pW5Zldx++G0
olBSEbKtCKWSznahlDwqI+zoq9rST2mr9Ph0zwZ8GqtxMXwJ0BB4EryIlcZ9
k02fmdo3Um2nYa2Hyg/m+75GnnZfXyFJ7vQCGZKFZdxt2t0olBGC1CRvYRFs
ebQs9BoW+aQ869x+BsuJmPI3ETU5kAu/Con1hf26hU1L3LDUHk46pPrxfk76
0rf9iN292RJZzA3yQJK/PqOMaAy0eRKQ+1HN4Uv4UnbD0sZnXYXOPLgnglOZ
ygdhs9EiI2yDUOT2Lu9h21BnlJ/mDJJ+jrgjNx7gModtROWUxfUNj7U/ArMm
SlzPT+9I3dA7pHpiOheHq/4gd+/42jwBMSv/3B9S4cy7qDoN+GZXUP1M4jli
lJM4C35238CE/UfdF3lr/DqN4x/TJSSnXMDdVUoKG0l0QaeduExr2+uDs58P
nCbxMmAD43IDubVBCAYA2ToBwAbsCjXrUVgb20fLXPI+XJyUrEAlkXXIG02H
ytcLOXwuTcQ5LAiPXE3C3zaZuFaT2pJD6eWvsKeKw6bnqLbTw/TVXTaNc0wt
S/5ytKs7TZVkIMOilaNO3+BeNIK9uRLO12vK0f20dhLy43yUq86QBv4gZQJE
571neqssZk/yfH4v7TcxErhpVB8++Bw7MQVuEqVmnwb3mGU5QAhvRjWyLVRm
B0FnuRplgpBukS1KCRPLKpJ/mCOAgsH3PC9igN7bgDuDQTzDlD0AC0/wvXpW
GcF5VYXVKRdoBWSA8QiRG+FvHOR+RFgAaOGPIY9rbJ3DCMOwA+o6rNytsv5D
DzaKvVvUOZSqMASIbfVMW+IjtUGpWnSENgl9Both6ngHOHSzNe/ujkbGjPSI
9XvYLlElgQ7e6NyPOD6ed16xZmj2EZwpsbsEpWCsEUHGVrjZtxvw3nsCrOXU
FaH0Z1aXK0maiCDdtboDYkMNyy+g6gQAQ/fDpaOkXUAr9Wxj8g6vu8cVkRAj
lvKcalR8/kUYOJTA/Ho+LYAuKYqzy08JhcPS+1hMPlVIMEO3t3W7fxDq1T7p
Eg0JMz8cZdUr1exrAoZeZVOvmrl4oI3aQbAODvwnbUPmfs4Ost6a7fOghRIM
huQ2QO9rUTNaGiWyffoAFVRooJmGWsVLj3wfRmBL+nQP24xg+Y7zXqp+SC61
q/vZTJnZnU3uf17mxoryWLTB99S0Wr5hAbf8hTXKiAAI5i5rz7XnuhIBA65G
WNXZhLNg3gAkWjA7aJayFDQLl0JSTYt2ZOFE05JVjwTxj6KebWvosvVoMWmn
GxSg2AUSNU8Cj14+n0jXJMASkBjzckJxDSzT7Fc49WQ649aozqITSbjMn88R
t9bBN1E0/U0WHx7DQI5kMp8D5GciKVsXATMQ2KPGg3bHGBM2FGaU5rIEY6UJ
tKCkxNw8AGX2E+7K4yNeEBVkHVUTTUsQzSnAP7txteiRu/KvSMvOrQdt+EMK
PP1rZuEUG2UHipchpFoVB8P4i7+ZUu17szDFGpbIHMdP1Ig62yDNuRcS0tyV
klgc0YhOkq4UKfxc/Mf2QjBkeykEgi8xwqartZNr9kEgRjpwsukYFbm55DkJ
4V8+FjLAk0eJN8jen3sEFpVhpAKi1Te/NAWEvbCJaO7d+/ERlNbrob/6Y6bD
Zp/7Bs/8BWjy9qXd7WVC+SohBh9Ru0tIDgliEgwmAbskIyFI+AO4h44LoaSb
K24yC23KNU9qhHFUFNyPB7M3ykG3kSgbuIMzUXf3HMaDKWXfoWyzBCs9qMyE
iv0NBT1h7w2KbZwQpMMkYd5kVcqY++19ZKCtQqtZXwomyUmKUfbofWsAzGqK
QmlMVfiuABdIJl5CTuiTWh32r8BtJgcmXp3lqj8U+QvGg5NeU+AY9MxwIXUg
cFm0wZuada3LgLsyY539tfkaYwGOb67aDSWEZKpQ0lCBZ5yi+feVE2ZefP9i
GkiYiJHopy05EeBUKh9Xa6jYoOJxqaJJ12Wq1vRdnxq+ZAHeiTFrZqoTabIv
AoOlOhQwK+cRTvD8BGiFpEHyaboH6w+7wgKBZ44WwZ9aMSb/T7QwRP7ml6S8
XSDjx4qJCRzlfB48ep8+t8tGdrnbpj2eX9MGFNPN9QpAfo6V1Xanh94x5lst
sPOXgA5JmUZnMEtZiuy+KyjyRnXRHMqQxsPBy1enzTwnhvwtbcqa/BxaaHlA
OU9XdwkHdi5sGWTVgTNpeBM1Yf4cFyprrTuivDlRUYOHNBwmQA6rnlOBBkiT
Sjfw8KpwSqHVENgbr7sqf5Q3zcbAxpKqz33dA9lN3zlpaXeOW2CWC9RMy8Bg
75Yf9nBsw+5++yy1hodskUMZEs5BtQufwhs/zpoFis0GK3XUcj25gH1kYme4
GBwQ+YJxnpp93QYmeebsBuhWjyGbF5TTVTovvCw0t9/2yOUGOBsEeb1zHmca
YuKYhII/m3ldff63QSvlLGLGC4N0NkT1XUPYS/KqMLdR4oFgTKSq6t0eItS3
q4y7Sjdr4nfw63zTii1fqFvqq8XDcDclpf7gef7tfd6LkUxUkJJI1K/pVEMa
P/Ov0MnG/q7yzRVVNzvJqPRef7gYjSVcdvZUOSIqZZx4Tl5v43k+ZeplLxNg
O9ioIqyV0ODjI9YRlFs9GNEa/BdQzmy6mEsEjt1SbbryMs0Xk7zI6UPF9MvP
Bv7sid9pJzKq9/pB+6loy/HoZCwawuHjOJR+AcRXUm8Ni08Q4u/uB6YUUiJq
5wkcbk4A/jyeqPd8RFTC0KuMV3A8gx7tP6ZxHaTuIhjzfblwDSGxTPfNL9tu
m76lnUtEufqfGTC7E5UY3MAEHwfho8VrbtHjp4mOV6fxfieOPNHLbAweimj1
gJ0phvF4Y23mv2YoV+TylMs2lec2WnGcscFq35CeIWz4aX5YZrzfWQZX5nMT
HCpec+8Il0fVsJjFzHZgTNOSL/ZyqycrxGPs9gAdOmbys7prPoxzwYuUdrQz
32ilMHO6tu+2aj0da2DVdiU/scigL8NVUXyOdofsqjvx7WaRNsucovgyQn+A
kga0WFFusR70ehyRXtPudidACXO/ZvIJAZ7FlNPi7hRRRHpX0gCynYZGU91P
ycVT72KOErimEbyME5OLHp+RFKnbMLw2LMQLeWEqX50Q2GlRfHixOUFRngmB
f/Jh4UFwjgdxvE8N7D9r9JhfqRQLKSI6qxt9erDCj9hzHz3/vOBDlOE5sFdN
x19gySc+F/tKZTGSlbP6uiDE5+fCHPukyphiGMOwmf06E/nfdlvWchPPV4y1
M9xKgDoacdi01gw2HG1eMLaOXhUZN0gq5488dT94AdMf/5JLZdjmI6593GZ2
26Rvh3KoRMo3RpM0oCTehbRzPrbMu924Je/C15V30g5o8pXu3RZMTmqp0Ydi
SdYKuiEO+unXC7ZKiElLlbpXtsEMqLMRB2T4NnOVnzUHCSKVR+Kmi9AbyYPc
23r6grQYqDvNeUOnhUtLCc7t95Bl7RoxREKb4V76rAVynQ8n1CaKTuwK7mVJ
mwfNxUjfrToA/FsGd/38a79M6s1g3joPLXMk88Wn92spKyKQBilSeqgAW6qF
yE+tCTsIjPcXrqOoK0UXsfZK2SRPZwYCIVTCiRH+bSqWnuwf3tBJ71oVsyzn
8/KGoizNo/OxHLXcXcgSLjkwPqSRdklKW7etdC2g68dIGJ/PUc7A9DfV22LU
5m3ylStCDlHSeM5epeCJqe0ZdQyRnh5jqLh4hyIq1JdNEEJKvstyziRYygkw
z9Qd+uWmK9J+fcuZGBsMpIRkqtPKryu6mjjGOjbunGNY42xU1qHKIJLZD4Mj
l+B+Hw5ZSws8IFrrPEuBLV1Un4PaTbgdW52IobQ/LAgq6qdFfQLfJkSDSS38
oVlDcQwaiEwOF2t8NwuJhphz7nmmuR1E+rBX+uM2/wR0/ITqWrBl+ZagKiHR
LKRQiUaapjEBtEM9cZwtTH+//gMlrqTCFtxRz0gAVSUwZLAC8lY6NBVXbkc1
Ac5TqMJEqY/qECWPwj+5fkSae+g6HDfSv8Lwee4c+lTOov2H0qtNpuFn3KZ5
aorjtSHREHbFs6q2TaMY8euTw/XXq+mArl/RnfGw0GwPer0mWDptPIY/Co/A
PWGrqtoWZf99tQ5JlRTZbzFkMvsR3utsLOZB1JOXst4n+xZ/RwVveXBEN2ro
iOLvmvmCXXF1DB6g/5NzNeEbslva+RHm1Yx/eQCRDQqEZxNxr0kI3VpcmCYC
7ZDod2fe7B/OL3Z9ErLQI3YKuX5r6zXIW4jPC1bPasBYBVAi3Vy5LQ0a0hfT
dGgytCQTlNWcEGdTOr6AJDD+K0xuLiJVX6RtoDig6uC7LjoY9SgbsDb5CTcv
cNiEipA6VjSulNkeAED+OyKSl/2hh/VVJdA1Ul4zu52frKP6xEO00BJm9Kx3
4dqbLzsts7bse8WfKeFl77qGMe42SkLxAFPjCARSFl9GSY76IW74br0MG7tC
MWZkJQUXijUTaxgGumrM7b1CWmykClKuJjKKOJ74oCRAjw/WKxWCo1ZmpJaO
mPmeKpcRgcLZEHirZ335H8ZcHIxgIA77EOqfFaHe1dYyMdW62MzMzMNbTAt5
MmDvoxRS3pcORx+CNLp0NW9oBVmLfRG2FRXm+z3BAf6vSbmAsic8SQEVXTlC
bCEdle/U6SmnUo+z6z6zX07SyBqFS7n5ApTmnEEvpUee2e1iT6b4IFFc5gZK
KOgUzleWiOnu18nrth/5pZjjvsP7zgBlsXG2ZvdR0uQCrUNy95cacv1eE2RU
c8rifi52QcEGRUxcgCFVK10+kNsPF0KP3x2Ov3PECnxmL0qF/WYGdx0asw39
dXgjrSCt0L5OZMzWkwnlC615iDwDNnk2WW5P/9udO0kvLK/zDChFgdhvBUjZ
sGvtL5wW861Po+Bchd/gje3oIfK+EdAs/bpAnU5SxfpKGRcURFczexaRZ7V5
zVh2ISFQwVFYJioHdErzbXlJDVLUBY4kKntkuOztEl+Ltdwaeg4AhXztBWb3
jr/m1SRJiBOaHTz1AUaREaSUvGmfUkv1CdMhhCvWj8SPwWrCCBwPLLa//dBH
biyYRsiozHFGyd1BzSRG7oadXEGdGXBp7nZJzdllLbuIwMc5XSxExzxEik8D
bHgunXJowJHDfdPdLciZ1fmESGZp/iUHvVWpA+Olc2az1CteN6rG/zkgMpWR
13Vwf/jBpQEHASj7nYSyqjkggNOVI9gE5V861ZHYMoawSaFXbDjpMccYwUXx
ffChhCwK5B8zDXuD9dhxajmjTZBzDs/KOBxZb//Amu0x2FZxKIs2mhQRyZYj
KNg2Pk1oc3NHVQ16oE8GizmOoA/KhIKTC1llfP0mzEc5mOzPy7pVsbS7B+pf
rt9u8tFGsKUmKx+Hq4RXqkyf/8FozHj+OpsqOhRUJgdPOhadVSJBFviE7/kc
V6jXCvpKXdhfsWtd/uIBKtToXdGm8twPw6uV3F8FDbObt/bmtS+haO5ONoik
Pqk7bsTn6z0Rs8k0foWNltStCJ0H0KjJpU/UyLienQICbIfyZTnxt8/M5RwN
Y4absGjem8rbYQhWumUOPtoAgl9TTjxPfRd1jHkxhvGCq5f2m5bR9N4reKRN
CxfdcsCnsoqx6FwORm1w2vVW/2lQBSzuuV8UYK+HSyYPP3KL9ONhTIdM4dS5
+27gNvbNA6m5EBP0gnsvXozaTuSoAhRVPj/JGsJLDIfrYE+WgxOwn4f63iQ5
kdg90NfTlp0+iZO48LkUj74XCIhup1Tpe+wlDSJ301OFij8zrBtxSt0EvXU0
wvKtRESx1WH1PfFg5sT345l0Xf8VMPzFDO1laOXdto+66/SjfmtsFzMKrv64
Xm4WKtrR2NDdNet+wu4/P+OpeUH5TkM2h29OGDfcI84sb1bTRUVggEzFlbPc
38qGAkNNaOlQ0rZnDxRnexGX2nc3/8BBgj5uVcES/wWv6Nh4OR91ZX0FfbJ0
BJ069NDeQfnwG7pWtJPYlsuq8K/jb2BdBuyL/kxwtf7E98xV0gAOa6s1aWWe
IGlcvWPxuF4k+MKYb5KbqMEcroXNCvR/u8ZLxUtKjUQaultAbnODVfZsuyul
3AtlwS2IvG6ZYIA5knbjz3Lp9mtxjmV1unAgwSK/kUSVR1q7DE03Gl6nrH3f
QHA2GGdwN+JkW/boor2rHpUoC8zBiGBDtFXVMCBmSEhKh/TPgwKSzRNE59lw
9KfDQVBwO2ai/kFZEsdiL/APFV8yVJDMgF34tVKsYVLALAPx0MXaZwWqTA+x
knI2BdZaKKg1wsdhxyOkRBEWcYPaV07lOeraCcURdZNGHqCWOt9bX/F8XvHZ
0ENR8IwwVLqvhMCna3FyqWDvuHua6nqVY6tExvuz7n0a5ZKPaqV7gT3EFTh/
JR8X+Lob4kedDarPYs5zrlEH+dQaFpSCuI5kyM+vauvnrnnOKUq9+93iapsl
ATDLcKj+f8pLDZaSC5abJQmz2F4bvHxvzEgr6wfawYjcYBKTUPZVJ+tq41l9
Tnh06xd4ONMbGAPvwhz0kZpx1QgTL1lZaRuj6hKH2b1oMg0FiYJYwwYHPPj7
HMKnfTk3/HsdEWqSIa/pDmXVU8SAPwtfVrhqP5K68UFSxC/tHmJ6FyTZ7qDi
JiCjoBNd/Vos/PpQDbqf7tIlxx2NvyZ5pGuDUStq+se69I8F/4yyKjC+pcxe
w/89uxJgq3NR3Pljh6f7SqTfpSo/8QWVX3b0a94Ew/+oDt14D/ATu0Bifex6
EbYNvt/xgR5aXbY8oON217QKtHoNdRAvot7yRwfU7ZG8VFGLzGJg/fnk5hX6
MTOrWLX9eFlm3MD1eLhrK2ebKiAiOXswTL7Nx8efSFjr/kjOsH20SiORO9yo
GojIj1CDLG6agCJYCBSWBfQsz9cvoUJKM3ulkIfJ8LLCZ4EjOT6nBqk/coWp
S6UMCROX9QjkQuO19O0nHMdBXY87VMbTluCDKRDGkttsEFjUWA7LsqXfnJzQ
jnagU8koMW8K3gYalPg/ICmAmZcuQ6jEwSb+iqKRunikM65WvWNL622UiO7G
E+mHuCRhyHx2+Qf4sQriSppaIs9AewBCuXw0ulUdeddqi2NAl48IJ2Z/RXsX
I0RCi5othqF3dp2rMci4/r2AhU2qpBzIAuF4nFrsz0zIzF1EkPa3kFceluUH
TzZzNhyzt0SYE+7o0qdgsZlJC3Acp9oBJaHCxXg5AD7BE2KtZo96x8ajifYT
++zZvbLsmQIyQKfyZxfSvxHumsPNYxZTDYNaCfmLKXk8AMyScY6rYukO7jUd
73GWrG+FNeXCpevP/TY1pLtxYUQwfLFjIfveL4Mq4T5Ul1X0/0Q13UqHRhnv
ijJLuyAthF4yvEoDxbQOp9p2tQcO5Mdq1dltEDEFKt4RiHlbBSksz2pD+kdz
YYrnlaNXP/Q6R5rB+ucvpbQPTlIpEH+2fWzAacQaLHeYsvKsF1wpOkbTFPlK
OfQVhqDopK0ZAnU0RBzRl0FI8S7MXqI45aUHWkbFo+aQYbdM1741pTIayUcF
fz+BC9gCB2K5UHaaoU+1NVBGieSf1VBlyL90igsBE1RzRBEGONw3/JfQfkdu
QCxTFEIr9dVQlLlS/9Rd9ixRJZ8spdWgXKVfBcGdh94AafVpPbZqhE4jksPD
SYWOr9lH5MRZ9w+Kdun1yHVRtptIA1VhpHxuJfRRMEDaHPhbVerNXI5l0jpc
P7laqy+Ry0n4cHUX8BcAL/OX4zDUt0uWbt+BqiNUCvvtVTJRQfyq2hdYDpE3
Od7p3fzsD7jXIWWo5M6ArXMvC4rwKhmZO219P+05e8w9m4QSOmfxCSEJaJ75
nJ7YfN1tCb0rBN6l4AQiabc5bj8G91LHw6BLqZXv9PFjuEJOmedqogbZr33H
f8/gbAZwKsJqAGPRNsXOqaGsLM479M0zT2GvYoGkqs9SF03AfQ7M8N5bXl7r
5toNq7v4NJ9GA+0euuoBRn2zK15WpkJyJugzactCwuEXab7F2Qy1EnmHOjGr
S0vSTFvdVwkQYjYiq3QJHSyoDDLex1ipmYkRnZuwN5lGS5xae3idurjGWaDn
NeEPu3hl0+JXm5Vym2fm7oXExe9mWMu9TW+q3AEE1YG2ONDiq+7nKrH4T5Tf
j2ysvanL42p2vkQUeY2cWkRzPMA1ASe1reTpEj65NNWXDVFZW4de11U42RKo
Mn38lkSVM4fvw5vEbpHpmDfKAyh1rWlkpoNyInbMMd5PhR7vmqkxbyglDqd7
acdLWf6mNszu94zxD/pU2Rp4UzIGTPacIOS8kkYu1JuzWixo7g+seFcJ82YO
jGpsS7/FeY9IYXKf4QLZvcIfKawu+qEGg6jimyKvc5+bt9EkioEGU7BEvZTb
4tUxCFQfY3XUzWts8HqLFGzVpXHW6WN+/pwtI3pqodxqnHHTCacbEpf29Bml
nBUThEUxtcJt6r2MhpmRx1WaUqrHrLD3wvL0nLxml8IPqhs6ILxoG8+WF3Jg
gWNt+hwRlM/reWxV2CP/UfDVAv6M0hV6fZ0vFjDAaN46hrWwEa9bzkY3Ltiy
mPFq38sAwnmdGHgKRA68ot3VhjYfdyFjPXhfTvsJkL82EGMRiJ1dOwXc2Ly8
DldR9NXzNRHRcaJWqI9TmT72g4QlJoMmV/iaQoGMcQb5PQ3ft2PvwiMSvWOQ
wFa0g55sETntg6uYTHNua9MpJpdoHycoJSQUuB1ZFgDFlXUUSLXuhUJs5/do
v5476vuuu6ZH9zXq1U78TNz5kWFrlzYRNuINBLDjXQ4BnWtcsT2E4aJpzlSK
NOLcz8qOP6YUDYkQIUTpg0geMyKm4/+l8FfLNKue+9N5YEhqOH+pE7Rtc3sL
DRE4uSW32texuZ2v9i6e6ycfFC91R/oz486n91tGfIaHRCjuI5i3q37RxRht
ojTDLTFjrQOJ4yTaKqNqZkzBvYf2QZm4sVFqcJ2V+rmW0oCo5BUthuPPJs9D
/SwafUN0UgKeos2X7JOHG22/wSUOgIlwtxgefcZpvvEdb3nOPnayDtECv7Cq
PuA9n6mFRfxjNeX4b2R0tJyS2ShAXqHg6nPBRSDRvE0ypHxx+5O0B3bfuRUC
pKAj495Nzs2t73EBDuluokAILNg+PX5Jc2UPMG7wGk09tV9vnN3p69XZRtdJ
7EfB5iQeMFDWpJhcXfGg+1rQ97FIJC5Fa7MlcyCn5eyA/ujhHzmL8bMMFZ0/
rhsUW2RaFFbnFycTMaOlxtxVxDjYOX711SznD+ALlsKG08m7xzF5kx60ruDQ
5dSghCzkILR2XTcUmnbMjhubG6by9bCWBEAKXoY4EZT6GTJCuYEfCDNl2QOh
q9NExgEeJeinNns57wO9OIuoIO8l3QXH5eww77M7ckvquS3pxwUw9YF87rTa
Mj1TO2uJOsR9pMPfC+BlQpIQNvEvpiDPSFu/M25EUh60RUA1NdyX/orrreNu
xc+P6QpxNhhlnvShqxxiIUfCmTwSuD5+sjiPMISHosRsCfNub2cjFXeRjRJ9
RhQEwcweGjcgSer+iqIcEP6Z9oeddJ74bnm0n0EkCgkXtPv+LiOPipkvrB77
sgqPxnZKjCVgXjfMzkPpTMC+/CL1RmugMqpbqodhsUSqFWsn01vTAWWzna+G
4Y/y0rX0onUuArJ2y8E34qR/uv2WfxAScSStQR0x/beHHU88kODXxxe9UeqC
BYZ/6M5f7krQ+L4xAyaZFsA+aHwqpjN6BAb4XsBUfCKWsXK40QR5QhO0x8zP
kmUR2Mk94XsjBBgWzokKx/Y9qdgVc+dzjfI4t7jeWIelEl1KFACxF/CAnUki
OB8rNoFMBZcaCnTIU5cJgA4R3ud8IzW5pOJrIykfrSHDtxZ0VWuZBYP1xGRh
MWelHqDkthxWXHYCGIyqZFgdYDBbOqSNP2AgdWVG1jPjYan3LlM+QMD6m1cZ
7TTq5QiHLEMy9fc6etYC6vS8SqhfdHhiQlpoGZqYnAXLdCJPVQzqjMKGOoet
gpKeEXTC6SFjnKWKdmzoMk9Z+aH2AimX5YFnTEOaDCBeHtkghzu1nBPa0yy8
UAQhjUaV5EpIWEtQdiQavwZkz3kIx9inKyUia//0Q0rEHGoqMNi2VqAIAHdB
V9CzB+GW851VzNAk/tB1ncjQDAejOf8iX5ETtYfeKVGvLvCqYEP3Nk+EHmEw
Xi4GZD/SjfRPQiq+pa20LXC1jwO5oka63PwdrUveQtNQd80kyieqq3kb8vq/
43o01VgFnYDplhJD/0QLIeDJSkQfYW+DPBsObzgFuFtmw5cf1WEMvQReO2MG
UNCJ1FxKr9qPai5iIl5kJdZIRxIscKN9d47zxeAJ90l9S/naww8dEyy4eoFN
LtuFJftGxa9vLiNTJScT/X/7JiaYBN3zlqCK43I3qT3f+bnZbtQJTYvqmRXb
iRlPCSIo2MIciMxTqeacs4aX777ZFqrTh6CPa2lkgNxgBzi2mfAom/pJiLck
vbJ9VTBOyFolLJKeXb4c09IAStwHs74RE4uKXB5FqkbyiCsucKq28ktXGiLn
vqmaEz5St/OB0Usk2IlRNwAK4YHPsKkomvOffO589ImxTv7nStcEkyVAimlP
InFpj/bwv6rqfa/28bIhGfmE5Y9iYa8xhZ0YMeGU/BGfMi0dfo6Iclzm62NM
sal/T6Bz0YsyfXzHnTiiKfCnQHcFidsRsC38/N9kVkAYRP0QTQ+svhddImV1
5EpxYrokm2gHFHEY1NayufrwD/EXVe8T4z2u7mixX/6cQHPKS1mQRNcwQaPi
M9rCfvTFSfenwdKIsCkSdF5Rx7xPD/pWO03276pThIt+P9IzB4CZYGJbahUU
StW7q4xXfK4boUA4KXjU9+4iM3bJfE4l8+/70r8sgIc32bed26s4F479F30g
CwmbIOlAQWqx2JdUlqXrCQ6HTqoQsJgfDAs8jsPncwtGVuy4oXxWM3PDtYt2
mRIjTdHsCQmmEI1C1e8fR4w3JHWV6AUJNyEW5cW4qdCBN2khQ9OrMqlbPmvL
Za7dALBHPM0dch9haRUf2ynuBpcwjgQH3Fe0uxJlSEVG2HZBoXtSSkyINlJD
A4AEqlJSl1IjQQm2F+sn8EdXosEzIXAPWTh+q3ews2kfh19HmwcJUeGl8OMq
2PhJmpKf6PKgaBRQhPS2JPL7UR+fHMENfIJFAHbe88p7mzK3aDqw510tlRaY
DVakU6YNFrzRKB7SdqbncJtB+Pt6Q1u/Ovql8Qi2BJNGEWJb1OjACcomkEeC
YsZ5b/AY4CdIRZD0VPJw7In0uE8S04GapTFSWFvJ3gNJLF19s3KMyN9Zz+qk
vX011dnIaCn2Gd8ZkAZcpPmSVqXxCEEAxgMQkJDmKRrZ3Cy+GNSnntEdifav
7v8oLhQTXAc3PsDhAMgsTQCDUGqqdTRqIbb7R4LZiNsCZIebdCJ+2giKFvwS
RjfVnfLBWnR/7kobi29MbVDT00MAl8Qcexrzifdlkj7FEfrPO+sXnu9VXmXE
cQbQS4HqwCmfb/LpR7nyTR/koxNnJxlLSznBfhKZ73qvz6fe224AUC15bTSL
tDxAFqZ7S0bETaWv+922Risloi/m8pTLRxwHooiONWv1fnDK6gVCMSfaY9tT
SN8DTwXFltebUwB+e82y5CXrZiMIDHlkZ3Rn9/EtJyBmj+E7KWqHhMS9wkmD
IKXvHGqNxP+MCUObbsgPYqIFdWBsxyYAk0uD/MeJ4U952EcbdFi4mCJghUBx
lPg//HpsSEw9FbrOhVrLBlOpafhaIbIK/FEfZ5CXxaA8DZXcnpQZ+E9mWcGB
GNkCm1OWmf864QnXYF67xf8k5ux+QVMQ90FWjPKgU54u0orPG0siW/MlHE1e
4eUruDh6ggMKHo60qmMsd7c6rpz+TMPAHpshR12dw4dK8OZDpXP13Y3rKcNz
u2AGOVVIbInhBtPlqeyiIOcoT2DPipHl0noGEvQACXynmFaCVt6WyvGB67Ax
KwL7n8Cg9TJI0nA0UYEJtW4LjUQVdkm/3opbzoivR3C6QaxVI1KZKynP7G32
560m2reM8jk7qeYSIOPi0Z0VHJwPPQ2quQtpBZF35jr1rgr2k2J6yELUXpeq
HgShYGlqSqfgpKnY2bajkohHK2U9lwGxeVPS4UH5/HXytnIrXLoiHptXsC4h
cfOB/E/eg7FkQaPUwpnFdtRn8MgSe5cc63MU2LzQUxhr6yMUflU99aLCbKWJ
2Kth2NaBNz2BAAijb8l2JTVko9NQVx3OOuWB2g2dOvQ3EhDP9BKoSSRgPpZz
jTjjV4VytSFbM1ZGEW0jLrKMDGNW5ZQ2+zmx8H3jT1ydR14Kd3oFhWUow6um
iGHBhVSBtQqljS0GWBBpTEj09Cln0sZd4V3XRxKMz9gX9Pdlo7jDBkbLVfGd
3gr/v8myFlgGgbj1R96IiCctP4V1JO3lyyA3ic107+JZbL0NsX7ibt4ohHWt
Aa4f+/cTil1r8NHxP3Wusq9ZYWS/ymJwWN9/eyINNgifWsKaik5kd21NfNb0
3p+vDMk8Ktv50KmyuFm7oHKBtI+wx3KrnkaGk8RM0Ak0KcdwDaVUxSKvsHMv
ytAQguEwFpXhqRaTAcjYqWMJF4IieCxHu6lf4xk6sq/xtKc5VYgDpGmT3BEl
sSP1fJ7TEC7VnjUDo4CV6vvdqlm7V7VdV+QD9vK3TaqVVclERM2PwVS5ZAnO
Q59ZnuyWva89q5bnUMw5wYIylzrLYZyAwbKEN6r9+vfhf3u8KH8F4R+2hEmn
U1rN8HjT+po3i9OmossNlR9yY0tHZjnbBXIR8NOiIMNlymFFy0QHuCLHtUYQ
ObQ+7g8ydGyV1S2zqusnqTqdqpF9ak9NKPXUQh0fMunbEytwxgar3SaoTUW0
VrQEhNtFLxMFurpVj16RaQWQWVRRzuWvdFVYtA6i+8qlkCMbKVy7meY/oPEq
GWOfz9gUbgh8/ba1aSsrbgydqk0aoyHOnaASMEI2eE4avnv99OnA1VgVoPlm
wJQ111yiVLV3z+fqySC5c5N1+/oniUdbZCjBS5p/3910GjvA0QZqfO9EEXcD
P6QwTG1MeA9WNl/i5DiBWO6WTLnUVj2BVs3OpTV8evrkn0eQI9lIfsS7IcFn
SYTlJphy6aHHwpBKiQD+Hf+hL8ZSBG+bbhmByHzZw32CDBPHnb/2MwPtW2aN
lHSzz+3Hp6CEEGIGCVDOyoRCds5L66u9sTEkGQ+jjacO8XYFQM13350OFonP
H8UTOvkpCWurp8iqfqOhiqK7Y20C82MZCAPw/Et37qJlVrN5fkuhYqv8vnd1
Ovk2K7vqzRoefviedCW2zvbAZZUik1NSundy9YJEgiJFBXXE0wEMQoV2KPHG
wBpYfA2Q7BI5CBDpWpzOJBLqo1kgKQkP+OMmYQRPi/Wz1C3hS75I+y7wqJ3s
b/RoDAK0byRzvoQPBhR4f3eJSCR4IhH7P4MAcg2UEqNkNuRhPVL0D0SXAsQT
bhLpz2gb+rartqv6G8o6uTLqPdBVUSphlj2Gdfh/IjJ7cwaQJsIGXnVnRu53
+NR3c0uV3MXrDOWP31q18tW9H1t3QIjTzRaWFiAgpD543BTA848a2zmt2SNh
jxL534TbFqTLOS5eeI66PuHosxIGlfFElRiPdA758TYCvVryKjwffUuno3Xm
HO1mMLBsjYx09pV1hi2MMVJ2A5KS5vmiKEixM1h5G2lkle9rOvph5wobu7AN
v/JCg/y4MS/nn7//I5yIJ5OnU0SUJ5wiAdTnpyX22467O5W234Xf/x6gwOY0
MSk4L/poa65H90I21uStzSCwkJrIgnotVbgBj4W/pSsXdH+X2smrIlylYnEn
hBEsBGJJgLOonA79PwZoT1a1I/jpBr8fHp2WeTrJdf/I673VTX9ZfR51bvRe
JdlL3FDgm9LSZIlrgzI44ErTUunTGxxSjTMHHo55+p/EcxRNTyfH/hPocHih
dZXJ7zl7RhsSdSLoDGAX9Hob2JO9zF8UEmO4x522TNSTMwdiGG1veW57Z9VB
z6kS659UyB1QNIpOPASMREtJU7umKlPfIIjRFnbQkj39o+mgz328DiUIPrxj
kY9dNSBumUJnukUg6+IIzlUlptqvcevtj35BszJqqoem02ss9D3s8t8JVDgF
WKWD7Q+TDQkDA2pogoonzjzHvn/ad2dRP3T7QZP3130te/zUIIhIbEHHjV2j
ALv8gahKBLC8gch884VotA/gKJ3RsyAK6H+vRPgT1c5tgItGEirGEWD4l+cB
bYJ8pCgDcTFVVO7rT2k4dp59icNL9kWvj3F9LlwRHRuWKgbJg6yUcvQeEj9X
PTPGsjmnZ4ZmuT3sFatFr2SMDfraXkBMSpGZuBPQdAcceDxu3YReUiWVi/C2
qIZb26p00PsyC1tvEqN7olwAhv+gCGZ9I92ARG68gP6ivAjFBlv+9ZwNeuj5
M5LtjLEr+pvTIb+v/OsdrAVzl0f1kYjCZHqGRa/4fxXbdgYAJLKGt3EtpFO4
mfFUGMzjRwOrm+/cHKrZrJnOgghAX1CxBVZt6FYnKqd73kRrIEo7iDYhyEnf
1VA0s4VgAEFpnj1ZFR/tAWAgP+yPq7RG8iRTq5p1A6KpUglTSnmPtswyp9R2
2JJjkE6gLApIVACZw3Pgvp+1dp+sOePkOFccSGoEwTsP2XDztnZCW/L1+VP1
6d1NEB64A8upUK23JUsbZUw+pWBGBRKN9H38qXskwqbZQRZ08krO750ir+3o
5Q0ITGDbQkxYES2Fqw1XCxGZ0uQRe7SqGCn2Z++u2Y3OBTEu1GmS5LFOTEk0
UqjBfZ/m/c9vrdE0M2ls8xmw9NFVWcFrkgsPXDUBkJ/lIOXcMyw22BLt8TH4
n/iKWhHM4HOgewr+MTDcDd5cdmLzD9q4zpKIP7Y9tHRIcXa9szhxgja5ryMp
CG1MR1BaPg+j769uesPiD3veWibRDIkdeoqIWUELK2rfc5wMWFgO4vOlOtXQ
75q3OMT6T0605J+PCOnSz0VSgOuNhopwsxe564jjVTGuLSF1fjDVJhVpDWEO
DdaC+SMBxh16w7SLlT97VUgU+sOpk186yU/CGY32BGIVEUo7NmvRw72x3Eb0
UZvFROHl7dZP0BFTC9PAqB8w8YaOdDnU64+5K9SshiBnF/m/Zp3y5YsehG33
zOhqJx6yk1K/J93Etd58aeUY6tt27PJOhp4/JWODqHODaEhcu/G5z0FaiEMs
maa61pHOZCAu1CWz8PCzab9d+QcFtryiBw2Oi/djn/UngZQaqNl5pfMBVbjl
p/QSTzgLlf95GEpLtf/4CRyB0baya5djakmRlxmMDXNGzODnUlRh2Oq2eB4h
zAq8qs+MchTygnvvdMOqPbOx3km+J2+Vp8KhLRGXaDPndlcv2Gn92IpjIqez
9GyM7T3dDyZy5fekCtdEHAgXvcyNSThkbW5BUYu33wGIVXI7SYn9Ct4eqzOO
4y9nfG5skYArRGLNbx2+kZnxsqsAXAihoMPwJE9aK3TTTjxmS1N3NLIcu4vP
94+/ENecRKIk8SqYk+HGLBGjg1oZOrLC0zf7pYOP9zVElF9t9yML/K+zeUFc
1z9cFld+RNEMYZLI1Z+JSLhkzzQJGMt3I9JKfkUpNsOiqPBYyggVECPcsVb7
bGG+8APZBendXaaGglIpS2nSLUZ9TX+0DW8XERjLRJD4V2eAbJqztYVMUvlP
Hpbhu4drVVGJ4zcep1lUef7eB90uWJ8F0kXOYA+idUShAVA8ZFberABY7POn
vYVioI9qLwRbtYG7rwg0ipsxdjUywzesxGp9gCwcx1qYO0qYiHVY0mg83gIn
GTs94PIBiYydfb5tHuHvB8UPeU5RipiTa9QtmtoYfUtqbs+7TVKNWLnFTU6V
JIjs1AW90Vp8fR4ov9HG9vaDsGOHaNyTknCzYE9yI7z8NUOmr7D+zXOROE4u
TOmylcmkMPJ92jMK0H5z1UN2667u25Bf4whenJBh8l5AZNSkE3powzN/Lv87
JcMld9/AGE3OSS4eadW5usbnZbO+/aanvw68q91wgwrIZ8t37xjVKg9Q65PD
ZPattdQ8exSpUZrYceo4sdi62bEgO8NC16jz9WzPRoYm+Cw5QP5GLzd9SzVa
s1CilhoB3cBuXlrzGueGXOoFmzWcxNt/RYk84Xl5h/kH1JPfFYVJzbW5FVvj
+Ev1Ej1kL7QkdTIKb70h+LCe8ryj4SlW514fVbLTpFl2iPTO+dxWtA1DF3qq
AXTGocfNfdlCFKdeQZUoDrR6CqLN9PZaBmoAG3IApn7YmWlq6qDmlmKKZdye
H1ObqmJd4TmkCD/JwFcJsvpN5ipx3QEhTsMF3Gmh724OFgWuoVVfqI8febkN
/KP9mmJy2y+hU7B6zyzWhGOn1hLJOLXZ8twE7HVPR7SVPGTwCrL/8DaP3MH0
JJVPsUypFOjz7gbUVRedyvG6gfdq0YrAhzf3jToO5Lm2c5rvQMHp9L8cN+UD
cKpIEGPpxPAbdkuPDOBRY3EGc/Nlc6LBKq2OrQyepKnht1fl0NBCOTg7VTHO
PejHJUPQz8wk7/vP97UcTD2pJEYNmepFkp5LKx8Bh6C/CjhOZTgHuefwFy3a
hg6DRJyMpuLuWZOpJn9ZPAXreIHjcnuUpJancaPJrrWqQSGSV0y3ZWpJmT0t
PTbrx8R0idzq1++BzOqDWIY6Dgcr9YpPMrG48B5jofdfZserTRzwthysPyVs
DzW6YL+9+t92k/bUNEAOAC3zQA6iiIIK/clt5YP1uuJ9bfHyXgmlQyLFwsar
bqFwfIS26NJyonSiaf4esmKxXO0d/WhmoeUO2wLxUILCciXRcW/JJxWp9Zd3
WHpJhHSRghURfTzDFRuGbFTUXWaxCOuyhk9NV2EtJuxpw/Vmknf+3KDj9msO
8vN1925pHS7FTNrsmeipKmBlTaUHFWZ1BLTByKzGjaSU7NxsR+MNagIgLg5d
1TFS3qp7jJNR+Dcast5auy5UgmgSwQ7ExKZZK9EY3yY0YXO2drkgYlt0MPI5
j3AAx8OCLZYVhA2CYXuOPSz1laA/QcJMqDqVue2lmS+/8QJlOfGbN1yGw/WV
LNpBW0wjUm/+aab4VGFKrdtnf1rMkZyY3Ni67gTftWn28D9tuFA5+yrxpTWE
KyHiGGk13KI3yhbiUUAub64uva2a8eyJt06DETJ0ti40qB/rPpRtNVaNYJMY
gUMSMaEuTH5J78rCOe8zOoJVdSGOjjhOXx6Giz6/50alN6+aYkiUozjGb+cK
O3FUdw8rbWqUGI9KEM2F/YObWFLPLowz8WVEB2OsNa3+re7MRXDOKJtbPtxC
fN5BlNFircZA7Z4+LFp4L9DdNyp6XXwBw47IVq4tRJyXE7hh+CGgyWJQgs7g
0N1PBNUqGPbabcpLNzKcJS9VKFEgfIpmUR1sRFiMXitGirTSLG6IsiVdHjeO
prvYcUg6b4y4BkjgPEjeMx73bLlJMkLY2DBlL01kRKdZhggo+KucJveeTdit
0HIXm/+RNBDY1A1AsAmauBBySLQvGvbltG7rbcZoOTbCs/aB2qWQggTOC41Q
xyy+Cv5jzTfUl1RVrtQXDMbwOTCyyx2QPaHjiP+nSKrzAGqpbCfrs/22ez6A
N5ekrcvFWGqufu1OTJmcqY6JpitZYu51cfhWjBZwttdqS+Wpz5ibvq/QiG6C
6erRU0EnKZa6WPfq6an69SN1AYaRu306uu+Se5ECajGAqU0d7ypRjycb5XxK
4jNUhf1rD+nJZdPgQ4W9U5gj6oE3AiwBmsO5cqZ1AicBLFq2DPwZDCFfnJhk
HRXnUzMDMvoLAGZ8b2AjLcEjeK6mBoHwfZFa6/PA67Rwyy+z090Vm+OwgTSY
qnJ8eSXig/DwlyX0nPUP/iq2AA9HI5+LC4xDWyfhpxJ+KTmP8WoDLCI+nMNS
sQrrxRbaH6GYADNJFEmp1KqcFLmH/xAA1TPbr5fLpqD/cg3XeAVu7Dce+d+J
1zrrG8q/Evp/IY2j5I64r7rQfydI/R+wSTAcTDH0mCX0MWQF7lYbnI/LaIft
zJYIiphUX6tbohO3GXM5wukGDDztqmCKm9x9GkRmbUh3JZ6seL91wl74/f2p
vs6Vv8erbvj56i8L1I3rGgI5tm49v8j4FDxHO1Y2T9nLfebLGBixtCJ6o6e/
DLFrPABI+oFuJ3H/OoNUW9/7li+7iJoL+FRjgrezZz+DMstDO6vjPIAX84aF
p7cdff5xRra5Nx6Fny8GCo0S4v8CvYly2PVBHZJDYjrY92upyI5ZgyYlcwyZ
Fo+4FkjyuxECo0LWAoai1YakhEI0hLEHgyz3DzgzMNwLZf4SbKL/LC7Bfvhj
hKt4kX/T+z05de0PqnGaTxUwsJiJfEH6AL9ZZp2aEjMIK29EzaSjAEHLcajE
5wYFudAQPyAESLP98+x1Rm8OyUkLb/tbLDBjnXsVjk45muWPaIAHBYhSrkxB
s6XNDrmIpMc5eVkg0kSJgS5UCjbxfluFuuBAz6GyGyDjNcwEa/rLJ2sParuk
/9FnHbHFypnWJjrWkzRjM8gBrM/MKuuiaVclIA+94P330bPmVHfsRUJia9LM
Nr2dbrrHw7jro51xR5luyeCKVvC2PUeymbb+FTgorqCmCxhTtLE0tNCwfp//
VFOJjjyGfI2Y/A7YZAEp+PzCt+3MG5L7lTLyHQWH6QC+S8Chx12vWEG7L5Ek
zH57pfHdfr7Cyvt10vczhEkt70mi0kP0psjsFh58c4ynuf3NIfdREwzr0Zk9
V8I/EHK8fbOaavGKykacbU+ycAPQky5GGKnFltwsHP4ue/kRmdFqN6ltaY9J
Wrqp7eB3JrBUfc7KCGhgVoBgF4t4kr0ICqBvVFgRSmbEEDxmroJ0jUy2SdnC
hsnO/ePyxRA0bnNUKKZwznC700k/DqVbGYlrLtZl1eMDVl7y3Eevai9j8Ujj
qYOcxeRI10+T0UgnXIZwH9676QlM5Z839emKUQisl6z2S60h3q+whC9DgQVO
G26Kd7Ck+B3y6q0P7KUplAHtsNMMqKOKlVW3CoTjiGH8NrbskxAgWsOcFq8w
dZFEZAbtaIWhS+FN+9VikjIFVzgE+5BnwdTzdp8iHWOetDZxqexTygNkX9xw
jJ6mReL43qJWEICGphBS94W4+OwwksyZzIHGUcSdI1BhECaF4/NlFHV9epbM
kp2H4yVUnw81S3dth8CMPYK9oG3DtDxHHtcFa/jdT+PoPjmzMx9UIZst/pxM
0lj076dbjhnoxr5W8sPCxDPE1Vs/JVkGbYWH04O9Tq+ukpZCjfZ5m3j/yu0F
bymvC+gcP1b5WHCKE/ihI1oFE0n/Lv3Xbeq1JXujULQUvsyLkndw39xY16kO
4T9lKmFZXCd+fpRNgJ7PR9+nLqavgWAoFQdF5fhz2/tGdnok++YrccT3qg3r
fDhUXEgkH31/biN5G47Nt49Jt406c/rZAQORooNUCH59eb2OoGZqH6M0Vi5y
jq7yjY0f1//M6+M7qQYTeSOnykdLf3W/zse1c80u+lCZK9WqPbEhzA8YRkEZ
aHvBlZqCP3m0+jSzUEt+n9ejJKWn/8qEI3ohBVWIRgn9P4xgRy/+eWOWhP+p
rIN2NEdD8xxmDRxHN1W5wZ1rev9TlyBP1oLPaPtikpNHYl8pAD5HY2oHuX4S
gCAcgcRQGFRRlayHHAKKMimKwOIY0NTx2doLmcCg0TMobZ/DLPFaxAWfLSeH
V19HcIiGAacMLfiRFA3nZyM1534yW8tLOznfThukGN7i3U/Wt2bdDXDfwCLL
9eGQO04t4YmRNfiRmeL03KquFU0FWiM+Nc0TR78tSA4Se1KSqrkgsGlovRJU
2cbmuR1Up22i6GXGNC16F/jJd3GijlBuUSoBoIRInJrgDeyCu2zMUAilxoff
YFDkZiOU5VtrXQl4IgPY87XZzO7k65FPQT6Owp91cuPZdi2huOdyh+120myb
OX0KYZk/sNv7m4gWP/SHnUPN2PtE8CAvlRUIYJmYuX87r4eXhGf2xO6+JK1T
ttQNks8Cfesu+IXHSWJZNXj3CV/1d2hW5I0ZHbZ2SGzgWu1ql7BOK3jBYEHL
evNJg4aM0BVLTn2wiUjPjGNHfc8uahvu6rQfKnEvzqjsmwBFZQUBlZPFx8BA
+1sqvr3yMBiyF2lgvUOulLw3Bwh9J03iBpw0y05SRIIINZaSacqBlwOHx4rA
i8NnyJ2VWVkqYnS/gqkao0aqHklETHl20gmMZdQHGPmEvV8GSxFpUGPe7DF0
5B82+U2+7PVZ3ek6bDzXsmFQFu+VYkB9qQpqKL40CrTQRF0x5NXohb5fUbO0
suiI5G95E6sJ9R+o4+QOLlDBg5LtHC4U8DztTelKHFEndGM00+YjI47i9mQx
bYKq+8zMmuemfkpfb5nWAveSYgEjrRnibkO1DPiJQ0y4yVIjy0kdCuJ6g9TG
3lQEJk49kTEINAhDcK37ewyU3SUud7e/Ukr+/9WEjf3QuYp9JXDjLWEvlE01
p78MLrwRDir/aA5zM7yTBzgS/6JJT010EpvBPUAO+fDhgAo471JFTIGszXTM
sB8vA6vCc+lIDn5iiA0mReeEv0DVgFwjdHbqtc2qg8TuqeVyzJRPnJvN+K9I
OdSF54mV4xuI/uuELC1+qvrci4Fp/V47fBs9TlWnT/aL9vJLjAmvpf0We7yC
0zkmfCRBp79qOR81wbB1Hhdhgor4sG45RNZdRZ65oVccSeuf/nlvXUOjg+kv
/BfzGn9QbIEEmihoXSU7AYITUhAib8fzKhvwYpL5mqIeBlqu3dLfp6Thg/XD
CzsjgQs0aOFN8RDYn0YArmsB5SVeyucYZ1o4TV+KSfatJ0SG4GuEH3olbJwx
DFsEz0T0OYA340aNPUwtSGao7IhzCKjfN1ewBZT4Hykp7P0YN22rSEaDquwS
Yo3nA7P9tECkBpkRH2SLYy9e6if0r+gN42g1dSPwLifUdWSbfnh6pFgU71KX
ze34h+dkRY7Yrnld2JyM/CkrcC6kr4tjDlLWKrpNq5RTM+BE1Njl4GfjMOcY
Oiqx4Ld3F3myOJ5mx+PSMvmWOYMGpHwgz4xyQpzMF9kNvuvQnkvZ1clB+bQd
RTauGxpw/jN+NVlWsWM8qxkNyVixdZk4cdmz9X4PbGjmHqPGHGx/b7vaivKj
xwVtdgNxxcNPF3EYmCI3fg79Uq8NXtDV0MnQFfKCmtaLu2i33Suah+econj8
uxnyqvSbh6IrFfZFCRmATZWjowicMMfa846so/ddtlU8xQUw6mgCs/mpQZCi
ZB/E+lDoAkDX5ScOeQKAAxxLWDOuEUmi6aPhzxPV7BPZeRB9c2i4gd4faeB1
G2JQcoLmiGIzYPsUCefgkxjxWL9IfepAZaYF2Dn+8cgRoZuDMjDg7ArBU3z8
xZOsC1XQ9TrTxzBKoE9MXx/05gzelC2liv0CkYJZCGqF6mZnmfzCKK1al39h
Mv7IOQqKBSTBoZv4Mfl4XTFUZ8Yof95WSj3Yxwm1D25/p3Ky5v4cTtxaEc52
6iioNZL3y2j+DcWnZ8zB3YR4zZDHkSv5fyw9w1MiYwDqVBnXrQRpFYUoX1sb
8BqPZ+Yft63u/m6Pq7i7ugYXEyaoBxKsyeFjk+KsHoZoYG4nm4Q63AiYJyoH
KvDkr5OgV11bx8/0Zt6VHTFv89oAZKWLryjoiSYf55upei/rGTXNys7y7TSb
KzglBH2BTIuwGiGRKWAPYjtN00PcHPtrWN7Pi6U781qIuHwo3QMRgHg+hGX8
GgNA1Fkxblf2D46Uk48L6kZtwfhqkY+qvIoX8TAdpt7sTP/EF+bml2OwSgHE
cij6qOwN0Z1FzlRcsLOj3X4V4Gwp0eGYcZ3BcIxLoiAcwM1MjMDiRsCnBSG+
fBsVizFqEqsgkYJwxV6RHLWa2Rfcl5f6syyIhcHU7dTea0ulB1qNx0FwrEXE
g8TWn+livonk4lgGoRbb0diCLQaONeWZMKXCexct+FssnIisdCDXhgr41y5z
BQ/f07K7aXum6TeZ7QfO1596HJOkLUjrJ+rGjyxtjonD7wG0YY/o3Ce5UATr
rK3jjX35DTDdiOBIsL8RgF7eQoWuk6gdorSbVBZxHG7swY3rn8s0mcxtGUb7
W7vtRwipT3oaEzPdxbIjRoosVPtdYz0r3uOqbCaDNKlfkjHS2py6klMil6Ar
3y+EOcVUj/gCqMl21+Kxz8PUXS1FwnFaKENcYhuIHC4P9ARsnHv+wd7M7Zaf
fUsQkKzrRvaXmqGJJNwruOuQcZk/WNZLF+PUtHas/P9mAgZgGO/NuOH0rle/
FFeo5m6qekmp1vQO2G8wNsFQ6L1iGRKMQmXT4On/y/CaG8htMK8jDSjel08C
hlD+fv29kVJzHLXDJOCrBt9NQmKf3+UrEQWlOBkWAEJfvXVuvowREGxY5wEE
YVRsqXTYzk+/+/V3pmX+UY6F1I5EIGd2AweII4P8tAej/dOMUWa5DfeElm97
CY0bquUJYUKOfBjGdmcYflbGc60QSIQ2TIEPE47acGqGjgX1c/9RxjGSc/iT
0/Bba6WrwHbwTEfRrVxdpwcY0c+Y9UTLOiyfxrYaSdwlcEvYozAGMsBlDrPg
46yzdr7/73TyYJSpJCMZG1Eym4lsXLUSKtpUVhWS1e5Bwpj4E2ASmRYyFsxM
GJC1K+Yy/cSh8Gz1rMzoCqQqiv47NTfJV3EM2vT5yqJkIThTgB4o9WMbtWZ9
IY5HJJmOmE3R2S3D2HmX0a3zK6xDCzst05qz5+OSMqk3CAH5Lrdize9yjex1
gOwLAijKkJz0X+iduaMP4hNBQjIwZgt8xdaPxllBL5dV+fK2BwNon5UV32ra
pv+m3OLHlud5f2CUrlzpDUaCiplbvLfA+KtvOl8IRfRxyWNMHu1vob4qVpPa
1VMs6lB82PdsPkjpR8a9+WdVbmptlVIj7GnyRn20aHnkhTHKJHaQSIUK4kC8
riNO6vLiEWW00axgs5jWPsT/DySlezVp0d0dbISAu15XODhSXoeSFemPjk/O
Y/laBSut3Ccpmqj0BQbDmrcJ8j28iRGDP8psBVrQWTsBtdoC4kPzhbGPT9ta
QhVRcT6CPAPfIt1qioqwXIhb0f+LxT+BwIcMbY6jTRWBfX98or1YtSNTVTQ+
g6hegcD6ixcl85wgXdRFHWrLKYIyqJJyetPMwxUckIlbPNWVOX9GtOC0iXUo
iPx5k6fjhDTC1MxLH+62CB9EkKi06PNzlJZ1JAa+mVmtPFbesLyc3wsnLwSK
iLa7SD2ztv2YnmGQ0ILjNNqZrbrvMtD1lgdqo3n6DEVIbTCqzJNCZLImMKTk
1vvAqNeis87fHGOTvX5ZtRCYlMRTHMruI8nxo7HHocIyQTuTA3/llfymiXPs
pc4W0FXx+iC2hV3g7gGklbV1APIG6fWrucE5e2PVaXu0RcgRYuD6mQKOBkoK
h3DkaZIiDr++28azyKKt9fT3u9zcFrXhbfxdgc9DMDZuvvsVZdEkyZVAz7EN
4ZPeN3KXARD/DS7e9OmsUpokMggxo8bDDZzrx1u5qBe/waSUpHMcGdkX4l61
+1PZ79cFPfLH2YfStNOgcPQwV46Ai7JeeLx/auSVyZNdjKuU1YxPzdIkKYm4
ID2RjegyZTzhV2Y6q0L6Gg+dgBQ+h4pPHuKKohwxHyGRwZn8ff8SQqTiD3Lc
lDkiy0MaTrip/I1scHnCsXqO72tplo3no6Hb4cJceY8kz9bWY5deZcFf2UTb
m97cDaGhR/DrvhHXc7mBRbywQsyXZue7R5tkuL4U2KzMgv3t0cR3JQTNTdPk
6kc+6xlXh5GpJjwG45/9KqnAmx4HlW1S3w6TMfoQk7zwKeeM3rODsEhineQE
wbA8SCVHfQO23/S7wSb5zRnr4nz/fsQ0MZLgsoFIR724J8lHVkx6DKBpmYpV
TwZsdTwS7J5fCLMMv3uZGySrbA8Z1EuU0nSsK2IqAFA9MHNeFeba7n5JhXbV
5yEpnkDraKogTJ2JiP/fWYvCkfPcXhagIz0dVQTtsz80g/eQHoFlXWvI//IU
4dPaWx9P10cvZG9BrCm30NeyPEMNrjEvesaPeyidJmAEcpmWlP0VshrFtwJY
gVX+vUJlXW46BN1ULW8Mi6PV6eoKO3vT2M3m371SSjzotPIjJXnxiby/9fhB
UtF4sYmzxzED/waYsSHjFuKhpXmdrAmkk3l/644b2MHpO99csWc8On+oEiv9
S7EhEnaL1lztSe1W1oT1cJTo099Q2/DFKognRJ52t5bNvni8jwzyKAdBpNlY
nt67Ys5xDo9yxK2u4WvnjJMhFZ3xjU3MiaSfJkqS/7rW1mEFH9karPWTj9cT
ddtRqH4uYCFea4EcqRoX51ggwHr5/jiRbtmNxKU4zvDrHcWGPauYlFyrctvG
aPla0OayDoU0/qtAitguBdSdqgokPr0XC/EsafQERumr4hRrMbuJxUmo4WIH
1NUQ146CmKr05afSUdwYtZ/ppKUvVqNf/Ppms3ffKGj+B5MlEgVaSC1wownY
tUqIoWZzzHooLuPjkO4czLcX6JLh1P9qDdJwz2fC0LG8s5hdj9KFwqGZg55L
KYwGLbZHNrKEpL32fM1plk/z14EZtSHYO4r+Ky2T494rdl6XW+D+nEoWPdIN
Btgzje0jpoJj3EWZ2X4NCmLF28v/gflBxhdQ/0FwiD7bK+gJlfQy0g73pqzv
F3E6fFQ0vI6ANILIlWgNQuzaiS60w0HzA9nc1im5UzlvHTkKcBhdkJCChbBe
ZPhsGHfl/qlG1cpPddVmEqaECMYldp93HhUUsp4zzYVx5g17PZeLdR5yxNWQ
ol2RDj9h8fRcao6hpUOOxDhq2zOyV71JprmxeAlITdQ47E1aIDFQhpiiKZD6
s9ZIvTZZwlKwxTis3V+19ZwK12mFec6zCAe59dgPaLwpC0cjCTXl17PLcPPJ
jLn2jixPpFSlPF2Zo+6ihKheu1/1P5bTQMxfUG36orbAtsQxeLhXKWWW//I9
SiGAvF7SVLpzepejL2uZTOzBPKwWXP84KAQ03g/h6kAvwp99RNHwUYMgV3KP
DuhCO6wlTv5BUiQ8Y5hqhG9j1iW9tXJnPVBFYvNuUVeVnjLDlJFTimI5Rh1l
fE13EOmHnwMn9TNVz2Uv0Fd5Aq/kRVyAv9/4W4mOuJZAOqgiBE1MSKnMpiEI
b2M/GDJq+w0VmYd209zbl4vcC5bWmqrGfxzgOjE9NCsf5pvdCIJh98LpPtRz
unaLWiQIq1ckaN2CHX22tBiy9Sz1IO4PS2otBFTdSH9HD67XH3QhCKQHpsPK
33Py08s7l6lLQZsKIA+53w/rlPZO8j4R+nEtJ3vo7XmBdDLxXPj9QIocDUYv
sr6ICR1RzgMJzPS4VfQn53ukbtkz82R2wDnFywnlRhicmnotCx+YizLGRVNN
ANr4+i5B/NzEzIJNgEEtiae1bLJZtvwsB3NgA5xc86OqE1AaY6WwKVDzW7Z6
eceSAeX+uUOxUzMueBMIcwVVxp730/DMfScCBQTgkzHXbv7efQ3jwJFy123Q
sPuVBUtiGFz1/aWFfZIt32Kcxl8InXQk4Tl9YFusngkaW0sNzmdDk2IRvF0D
BEiiclWeTeKbrTKmxOenQeCy0Ts9KkvEk+2/u6o03N/eMMk6NmLyAdTF/9ns
1FRXM/BZD+wABXhKoP+Vhj4dMxiJBdMytlVfkaZiyQKvNO2xl7QrSycgbspB
iol9GLE2tPV086VZq5ozuSjSsiLAqvk0hmoszpaEayKbXLg3JD0QJvrO8kLz
WbpZNeB4qW81zMPsFecYNyuAOwA+7ZdDf3igv2aWVJz12lTJUIoChW9bKkaR
Fo3TI5+KTZuPkEoNANRUEvCJ4PdpbS1Fv4I0vPm/wxir/B2+grtUchvzPan0
mw5TXlZOXYvRWsd+bmRZhZVIZtCUmuwDofA+3SeLNaJBFz4TgqYtgjFayJ6a
XrOD8lcAzceZbnB+cGo8KG8gulhPBSoykoQao0hX3FVtAQuWTQ6h+nCldCzS
FzYJDAsMK4PNvgnidOPizIaJGxibqIdNNpBvUnvLg/YZs1WPJuWoEXdn4f8V
2FHRAZQokZZu9NFbUKC81UOyED4ZMilVUMjlqlEnbs4U1CfD97adX7c835KE
pN59YgeGEp8QvNI6DUIl+RMUs8wCpTAQc00ANO7+kcVbMPBKm5qcqwuUo+5F
wkkIYAhpk8ea3kX8b7D55R4/uoy7WG1HaJlOBgMkhZumqjbPOP6XEAy2Figx
dJKXx5jxCHncrlVnlcT2tn5yPxS2RNdWyhAEj9+frfPHFcMLo/AWGKuVBIjz
6CqDu0cTCmcuYTOlsGe8s53lcwtxkZYTnTsvnRx58KpkLINHB11GrN5Av/fR
qDAWLBkXCxaDD8FjydJ/EXRoIiyJyTfDXkRTb23+CQo1Kx6i7OSdIB30Dj2o
jEJ+uJtVdyMsd6QZ3v1crvkdQweOPF+wU7FOLlsS7HaWKK8wZdN9RMa83eqM
Hv4Uy/WDqE7W42/ck+RoN+fe5oHQ6rVhDRvxGIUNG7fk1KiP2jIG/L98Kqwt
T3+eb+hjfzeYohFP1/XZO7wcJC48M1ElRVSCAWEWvCF0/4wz6BgiLBSNuQl1
35CgckOIgD54vcLBRDv0hw2e4gIon0kksbG7kEKGVp8thKbOGFJKC2gfdl3h
NxlrtbpakI4geRbuPBPxzkjxAYvjyi2yoYb5wgkBbBjT/QOnHWIhNQM7Pytg
57j8QGhpg1y/oR4KbSgBoWkaMwEnEleKP2JGfsSUWZWrEDg194doUsEhDyBe
sPOZNUbM16GExbUAL0+UKEa6Ezt5nzBwzxsQRprQ4zRtsYIWW48nFCHO24AJ
WB38HtWuMs0LWAygX/hUFLOXlwJHtml4I55EOu94jwG+LQ24T2zXDGxGfhaI
XBQW1tEOW6QFF6ZWwprwRu4ynzcWSewfqyE6MqMVdOR4D6beVWZSP9wgBGxo
zjpN5p2JeNi45L/gxA/risJWYytF7w2Um81L4DIOBgZtjzrbq12PHPks4xZD
yTtoES1cwi/VdYCSGockF2clj+NUmqNdUvqeiYnBFFA/IMrZxwcOoPAbYxaz
SQt0wNYwHqyCoZJtA2R0fkF909oI/jCD9/OGDXGIaS8IrkC7qHM1jMIVcJTC
/a5VI26cDBw0MPd6C6kvTVLWNLji7ja+cC2y4etGgQCojDRG+I+s9m2R1sbi
g7sPxPILv+sG1nSe3QQGbTHXechpRDrBhiNL4WOPV/KTNzwGcxI9I7HQ29f1
bUPb5ZsM8K3g3fsofDHQgT+cn3uUk0rf9N4GpIgad3t1APkMC1kKEZcBUr+M
/RTrYvwm7xkeIGNQLRVYRkRkixu7cL/mTUAxtRduYnNrRrvat3oXUkK0nNw3
S6d2kMgdaE5foA6HOewXGhkgeZqA0P70IgWjAvDFfrOErIm7J/4tpnxIZQdQ
RksoiOwut8TTlXv95YQMcsLZdwQnvQGR7RDABSjILHQnuoVyQryIalx4NqHf
OTrrIrzppt12s0u8BnN75G4uVy/fFDs0RKI8l0FaBiL0YoVrpjbJwe6Phd0F
o4S7kxrsmSa7zmXQYcXkYEiz+YEafvqOPS9CjlsbbRrjbVsV1ciuYfVGETC/
UKSxBIxjIkYiktPXfR4LNSkyfCwVFc1SlFBHFyD/b7voXkl+scmSAK6pWb2K
HYyBPgxexq+FAkS7ARP+gQt5S0ZTyOqm02Kw8OcNOD+zPOe5RjEjLPinUV66
9aYtT9UufW9zuxqC5KauoQEc2HK4Ixmm017k8SbTyRrXcxkMXj4JIyWt+fUQ
L2Qh+WnxrwrlcvFXwUHCQbI52YfphET5uNHP2i53HbXLaM/29O/ePSXpNhdo
8rXI2lN/0Glnzhnez7YMLUoNj/2mvmUPn4O02MhOIop59+0rO1dV8ZMPLzBH
yEeEifCuQfy3ssgNHHqNN3t3Gtd+qwsc/iPxEKHvsu9J3Dr9OgitF4ACsF+5
0MjyOdr05rgIajkQPiJEOvr2gUEGvfnTMNavDYEdgbQHuLNncRRNJUE0vTrV
/v+Om91uY8tFVI20EdjIK/toPmHGb4hJmAmDrdoT17Md5EMsKspiQELx5uEL
N2YrWP61iovp0OZX+W+2yjlWz8IQZ/LxV6gAANwuAbwjW+KDjjx6i1rKHaor
8i2e48ESjKbuSF3yr3V0xcqhjVpghEcXXKAh0HdFFT3t21dCDD5V1/ZmN68N
rQGxNdgwi3x8RalFkOytrOKtRjZjytg4d/e/VBBbjCsgafpSAnhcahhseWVC
9zwvkM3Knm1xZEQvDO9XZd4DrZqxhJYbKyju51kvqXkAy5oodjWOuFTL5U4h
XmHsdNZzaZNM+4FbQ9Y6ovKornwBnz+fdYADeznNMTAc+hHttF0jsaiIyd2J
r56dxUMyRrFSdQwi1W0pKnD9cjZcQer75sthniGFEFvk0pA1zogxAmVB99Wk
cPicJsobmLsunZyg33AHf5tTWwOc+mxAdWigfXZRkrxd5L8LZMju8HwHZU7T
FB33A7ntxLr/2sO+N+nLWCAl2EjME465cTcSCRw7mUf69nWFYWKZ3BZvoSPf
/1dNQF6qkPizw77yC/858Z4tay5vV4wvv8PYzhyaNEO4qCPTxe+Ip0uR/RnL
e6V85Rr7l/3n/Hl4/hnNerOF7zaWLAOAQFd/7epW1tGNEQVEHdnyiRM5LMwl
CrygaG6+GfcsuqkuKNjoZzCfKmKKkeRHBwcNCGMdAcDfLQEw9zxRwiwMn2tU
/lnBpInfVkGWqYHS7CWOTjActPeThGZ3p5l8GGk9wBK3iyoNtmvhX9Y5z2L0
taRUxPXoG7p/QLnK240/iFH6igVnnx9yzOnZEXcJrJpj/sITh3OQOKEfLS5F
6lJaPISt+VzlLu/fV/7f4V66u79cecUqMq1kxKxVT1o9RYtJZwE+x3Yw8L8s
6L/cM2moOL3IjPu3m4voRtThXXOUHwgz1H6bcHQRaLR4NKeuDcsuvY4YSAbW
2dcqGKgQFglUypzA/9rvxZNkNgSnusBWHmtv0rixBrfiS43SVKshhkRQscrj
cqIdado0kBhuLkBggukHz6aAfdciH8y3221RzYe2djrHenW34evVdyzZi8XV
C1qndvYdWUMQwUgjjyvyiqszZgS3WvoZrWKNNzadohNh7+VyGWAxnFwYCmk5
T/R2mWWabr1+UJX6aXK18Fa4N7UGlIZDtYuQlG3BQhT/Bud6TgZRfckWDeDb
UL9eV3u3F/cVDrAdimXkePf0rJn3rcG0F+x830tImseJzX+y3Ajyk6Yy3ZR+
RUxjsuteZs4e+sITF3+M8T5FXvKDaFjVmAinWAoWRTdTNH5kBudz4Cp1VUAB
B2XIUAO/oQt5ox4+B0ueRVKEeLiK8183UjpKjsFjg4kLnhD915EJrUQ3p0kH
cS8B3vmk/UtVztgDdrvKX7cm3mPoqzRtb0zbd+nJg4ront30MneU7HsWpokM
R/hpdp5mPTENWXuszP5mRoiCOB+GnW/W0NqsWqOYtCWDXrmpi0VA9dp/r7fw
rswTH5JA/7Rx/j7aWF8Q8+D2Q0DRBM4T9u3jlMMYCPJEaKoOdT7NXGg5nnwy
wnss8rBnmzNzpzJzJ5EMl4772Pae+H5Np1kmlB+S/0nmA7o910yqFBulJGtW
Zmg3qSoL9clN5sS9rYZARzhjZ6MFliS1mVZ0YFYB1fRF6FYSw7lHR91Xdvl5
QyUEYklKtFloK7Q6JpN1b/IVQLs96W0gX2a77z1630GKqU5xQEcP7mEoKEy1
exQwdNeG6GIukJfNGDruBJdWnSGGb6Nl0DCnVugrjMEWeJlxqpZbNqxDAcWG
18tGFYxP3MQF7vSnNHKyrkd9UT9owO4dl8reln+rCK69aZYIYOwJCIL0qNMl
QmSzgzgT+XgaGYR4wF4uEhrysdrn9uu/0o7REfsBstjSpPRMc3fK50zWGkSz
XWijDefmIPD7HpKk9ZvlF2fYkLQZJTiqyK8eVGB37rkWabhDikcQXbiBdad7
BnnLyPQhglmHnGQtAOckuKJxxXtmicb2ODwAwEe2ESTr012Cm+ELW+avOu7q
bm+V5jNfaN8VSIFCAtW1cu4pm0/vGGaqHjdZspX2pHjXD3PtA3jT+BgvIveC
8byCiS+N7R2tq0f1lrIokR5fVHUnQnoyavfrwOOUYtY3L+g68oGVyXONfHnQ
fGJR9/5om90jItTxAkvxBqWtG3DnFZ6EWZcyTxEyGfEwbfFvoZhNIK0r3hTd
rvzZfN1V/zicCK5o6cs2woO2riKvRAY+jatM6t0U/gPqWuIs3FC/hDuURk8B
yRt97R0lJJlWANVw/IkDz5AvsIH2t0XHUwt8gbbhkUhKC3pJ1zXGQQ/3QYoz
vFEnuPznCIbMB2uyZ+PXGhWf6w4umG6EboeU+kMKJdw1zDvbjNPYCNvs8pKV
1uVfV5gpgrqbA6aoX8/+T+eGDMOjM+SJ3R1/AkKTFtADMMl7CPQSxVXd/TeF
KwRY6qLimn8ZeCRkcSqIoxDLT0QawD/cyQDd3Itzz3qmylZN5S3KUIUmu8WW
eGzc2EL5yWrTWNNGh8kVJcZ8RdTkOvUhWe/BSv1uz3OVNLvks+RhXEDSo30A
0H/neMMpsMmodX2WGNErHfIHybzzNns+IALr4kRX4jDl1zDUCfhK9w2eAv2v
VK7TiC/jvLmw6n8Zwzc2wFvEe+AtbiMYyqm9RLTShENOIkU5yPy6F1j8CuWG
+tYWdJGAcOEeihn+DDHphAEDzHDfPj73crQU8UUDaxtuN3MRpdP5RkIWQ/rf
58Y/x0mdeIIKpeXdcBD/qWNVKLQ2yDaUInr11vFPaGfiHGVPaOVZ8iA+I86+
MHqI9c+yBjJG8BWkPyNGmiGoQZzC1RTCxq5vToD95RRIk0p+31ZwZIBNxdAt
D0OXsu4SGFDaPhy8t5DSv92MukqSmMKn/VkoiS8Q3p5RpLfFdSkphVTbNHi/
eeG2UtFb8xuyi7DukWoNAV7cgxPoCa6baGIwQ84cJbEMxKNwM2hlj9kahh76
9HdbEWLxYc26NLcN+PbIX+rjdah+3RIL0S57sbmyueUBMOoG3M494jWMngUk
i1tE/aJ0LCQlOEE8mPOWW7Y2qnmpuO74Z+G+DyUpYLWCUS9abqIURcgpOUmb
vgywScLvmX44Irq9PFoIA1lcDvN6AR0aWs9DE53ndAPXU+UbpJLQVEpm3wgY
lbOmRsCkj+djBuBuqd2EoeuB9dspguLzF4kavF2GLJfMXPrRKGClyZBPq9JE
EHLMrbG7mq7Prt0HmsqGA+uQQeeGAs+zebqg6o3Wy8iOQxNGUYnbJBOLuF/W
j5uW86CnpoI1+t78QaUsA0m3yb7slFwM6sLwm2VBxxa24R/pBSgQw10u7TuW
gi7sJLWpRzsIDmoIbRI/YbpeB2DS9sQHcvGSt7XdmNgsChdcRb1/MJ0gqqzx
msqZ88iQDjikFVAcT1hqWi6NY6fKCQCpFsuRIZxaiaFasyaITR/YHd7NRZCq
ZSVcKvaDTzqio/2pv+szj0fElB+8PXTQ1sgK5XVye/iCViKs2N6e3qNA4gbG
zRJnhZr6xfN+k7KKAgecqlRAcQPGBrGyNBYs9XwMbBW3gdlGPU1ccKVcXzoF
Aj+O4/9/k8sukSSn18nejF1rXp6BO8Hd3Qh7+HP1kcGoa8MV5fXfAGZJm9Pn
QWHasjpBl8YRjcryzkT6oJVmRWpIBaLH5h7xotaxAh9veFdmMwBkAE3BYzRv
/GCAc+Vc9hLXQh2LoRKrpF+WlMHVSJXp5Q6MW5j4DCxUmHv4LCJGTMyjeyyk
Kx0XGrZiH1I5DmSPwBdWdQepD2R6BUd7AyPg7B1wxvPJF/QZOCh6tWymJLSg
M15kQshJ1S9Gguscx+YzDRkA8ijfFVJ8rDpddwkEj0C6l6QgdisDI/yAVmD5
b82MqAQOaHOG8u8b7wNDeCgnzLErI1qR26CtHZGCLpq6ChuJKvfmPxdd2tpe
gh0yEvSc6ZqLUESsPvIIsqypPZ+M9u7G9ToAI/ih/xELqlPlpPBcwWNlFPPY
CW9PdwcFFDDQEimR7Q6Ew1Cp5/WniAqJfLngrhQzSYY5xwPY0x8Qn0OO75FT
Ypmi5MEgvFpTQ2QGtOb5YVGAxt9PpD0l33RVK/CHD1HWJ8Pne3iDOt7QerVF
26/DBe1GRRt3OwuOeaAnUJiq58yW/Rb5pA1nxJLKKCXG9yf6ed6pHbLVdqts
lHbUgFS3NIyLN+KpSN4JNe6UigdbqbTENLbNpDAjtvv5OTLVuGokw3wHyJQP
jSd68iDE90Juj883Hsi73ifm63G8P+jDQK2iJQxOFEGPwcHFYTAH1NDxR8Mz
g44AcWHk9C1+fD1pNYdD/Q5loQT7J3S5+jP8Qejse/ZacnSLzKFRhvcVRfNC
NmpfxZ0efrQvoDTfGMnegYCvDG0A07OHGd6RIgJWZiJ659rpSfKgrmcGl8nM
PjE5rawKeZOTq9VC6mNgUSIDFG9BmUzsZQ7kW6Mc85/6f1/GvDSjgEVEnYGG
0X/2hPOjVOlBFiE02pi2dOK9t3v2XRtMTfXLyZWZr6ZXaDb4ULisiTx1Js4T
hI2nE/KcTnpKLvCobEyvcdUB+df3Ua5cwPvtl6SwcP5mv/dF1qGsmO0eWqu5
4jNWPRXavLTXziIxaD3kSS5sVXU7m9x6tkoAZIXLHkdUUTa/TAAMAZa1DToN
LKJN5AMWB8yfV5s8VywHomHiex9sSt3F48CjqtCXwW8UIBrdxDs5CYzxjaSv
JY0sA9tgXmGUe219epG8D6UzVs46rIZK3DkSAVoYpBwloAS5YQm6h0dyidN1
m98PeZh2qzqZCzKJePbU6+KcTd+er9GErWdAW8buaq351rH3MneK+RMUy38P
fOwBbvKNunGLYghi/l+Z2vZ798/oEsGb7Tptd8vMiVTNsjwOgMGy3Ba2u810
iPmneJuU0MXT6LHf05HxKf8hMjukYl6UiZQ9DUjm8PBUnAsdRhK26gIDRJR+
JdDaCJVG/taHHKifyK/33DGQuH6ExFe3qhWCWogQXUysySWK1OLEb21MujvL
0lfWomK5S/FqAbAjhNYkA4Wc8z0FiYgFyRx7XvNIgSGfHTDQR2VFzy8Qe+Ol
K0PiUuHyE8itoNhhAk/d+skiCBjM216RoR7GLiV9UvTqETeyfbLBLXthZXR1
9QVGxs3IKHloMiZI6h4XfVW1As4qQBcML2LLhLtEQEMXpDwxz2/Qiievk7XX
+JQSRnGZtVoG7qvcgyYVtUZAXMQnYgg8kPHb1fU6SEoAkU6wWwu8zM96h/lx
+0ILPywNBMm2QNc5YjD8cso9XMP7n1k0DPTes/CHMb7cyk9Yk1FLB1BHP6eu
rwVjIxKKeEd8QZxZ6IY7Z04kkqNRO9T1x29IfhObOcJqcUBreeMjyA8J7CS7
xwO79B33SlCN93HZO5jcxI2JECn0KuDj+ZiM2+qae86Mn0z1OWRhh1pQKXfS
316gAOGFYbuCyeG4ZKJqAlVJKJMTG/rDyN45ytC4DSe1DsHnLRWSX87F+49E
com5PCzkG1AS8g3p/wtMRhAFEDJ15fU2q5fjH5+sycF3xqJ0S3Ft2wvdC4Hz
2D0Ej8HQJM7pom5kSUSSd1Mp484d4LMhI1vi7dWLjPBxIhThR6l90mIb6snm
gMT4xofwSeLblthShN0QQ/HgQDRaFHbtcC0IQGuiRgkEi4t8NYOQNGa/rF/8
LW1zYHWWEq9vwtPhepmB2d02SsCATGb0XTcwDi0nBtmvBXdOKkUXnkqNy6IE
/Om6tcVFQcJ4G5QoGXrwm/j3vqgQFaUre40bXkMHxIewp/ZrYxocs286WElI
1Stntkh/i3mmEu5MtQL+8pCPONxO+Mox9PhAOd3EPUhN4V5p9iEvgcVSWs6T
za54p6O/FU38aoogGWUpzC3n/19i3j6rJyMFJWFYeS5YN2KPwQenFQK0uupl
U3RSI+GB0Vi4zOZOtk1e/xLXgrqDYywQ9QA8Z+jiERyFkCmExLHNESCu7GHO
6YCcSFjoeVJhse+MmvWESa33Awvp2RQ46DJz0O0ONdTQbKWYdwXUbAu/ggot
pVnVnxg5nJjRdxVxZX4Hlhwa5pmnM0Bw1qTHVyQJ3G8rUrOl3qRuI+mb96vX
DBFLQF6nSudl31ABa12cV5xdU1sVVAovrGAns7x5igRLBTPPeOsgvVDThQEw
5YdSTmvfmOrgwhOqoL9kBfEV64RGhvP7X7KEY/BODyXUzj2WoLow+9XSDzNH
mzfQqMjXrKLQ7om4oTelPwXm95CdR/Tsi1669dGZ7iM/w4Jxz5volDusJ5ge
tJxhjqS5ibJH1L1fpyCN4gm19onNfNmyWzL81OhjgHJIC+tt6SWza8727X96
bkCMsjWmeo8DUxfqhNTEl0F8rckvEWF7p+fn6bFTovlwh/JiWmiG41qPlEUs
+wgqaZJVvplv2Lz+jmfyfUvB0CNoou/cWpzSL6+a58UNdrzaiuUApKq98nTZ
/T45BaE8mapRV2eaV3n14L6eqziQYsimOMTpflC4DcxO5RIrDXWbY2ejIjeo
JrdBzRXi358O1LqK3R6l5PlJ4cdO0lhMp8azkqf15HSord96cQdiSbh9Xpk2
0D5UXhrUGtkNZPH3oL46XcUy0l1zTl2CfAHc+BxBPH8M1PtNPATLkiw9Wmos
vx4tEWenY4qRVg6w/xg8eKZxlDnCTUA6542h7hCvzNyy339q54fkt+dK43pX
tlUGo/FmiEQ9z4jk/7XABYq4j4+J4lxAYTU3eolbCN7XnuA0N0UXVOu9g6vC
yzQDkquLv722XgAViBLQjBCB2HldU6KtHyZfKtszZl+fMOUWhBCD9SiqeVk6
BpMppZ5Zf50AQrsArAtvj7B5hQpOsXIlQigR33YCvo/ht2KvIejtKJ2yezzN
lUPxrpak+C+jDl8QcAUvkdUFtNc/xU+aqW+8iFR6wgYGQlJkCfsl0f5fvZIH
1Y6WnH/r+9eG3hivT2GYpv0SMsXPgOw9LRn+FZDvUT1XqsWFidfOLgzDprCe
mhvKiZ7y9nTT8XCvnptumg7ORYHfmNjmGVoSJz/njGbMrsjda2kbvoUOIwG/
J+aFFVXPXcMVRiITqR4X4/fk2EDjLMutrV+ZsGU10JcrXFSDTMfZViP+xqbk
I8fAFuCSR6g5xkbFYlJxtJVqS+HBj0M3oxAe7IgA2anqDA3XOiVl7OZjRkBF
obQJSMzP1ycu3MZJEzlfPW07hqy03Cc7QbQKuaeYd6m+3cbDG/y0frCUDNnX
rpxJMT5MWrMZD8OVrkwKb5+jx2HQosWdee6r2kvTDLRCpcWQTLf3GYZSm1lE
0BztH4vAmq6DddzFZkQYUdSgnEnRbnha39h1JyKBrIPTz1D6m3jTxcAowoAN
I8vI9NRCeFBN8GijiEuWxzHmY9xqp4Ouj08mq1lrROCCs6I/lqzC9kbPer0s
TbLiji723Uu+HdwAd8xjUb/HAJJG4UbN2e49aH1r1Fay9YvMolKjrFDPkomU
SGhOqUQrcI/GUZgE3RGBPTbNnhA2fEPK9MKRUic+EnqLDFnCXw2gsPxbZr1e
DHk1yTS17hCYdAoPfbxeZyhNBTctljKJzai+oAQWFtoAP8t0ntdIAZ5yOj0t
aC+vJyVVdZZXZvCjB6XnmLTbVz0gY0fa8uWWgIBAafRPh9GWAG6ftfnh6r7d
RahReYrXESomoYlI+zmGWR82auO4L7fUjCW1OINPs8RxHQ0wSW/+xqRP+wUw
sIUHCjscihWg0iFqcbBxkBr4ldk140n8/owNwK6cgpYg0PjsPomnpIPMGu4c
LQY2K6q5IVAm0j1dtdQcyVP4OTL8mdWNJ89j1QW/ILkr0ojzTWdL1Ckltb5s
7dNhDjiCbTntwbvHECzuzWwmTV82v21PcYicmy1uURuGq3H2yiKYPbrlhG3B
X87HFf/s3Ri0mK7Y1BgxaGqA8/hIjX635YspD1R7njS+/BF0YwK9i0PitLJ1
0Epqnh6QXVWSRCjgY9kN0Wu9JG0eIbUE6vKTEGeHr9bzmOD41pQReOzUKBAj
7UalynwYU7+Ub0mUaMbIk+cXYZ0Q+4qBLv6b1eGgDzmyldQSy50/PbaT23b9
hcrb1J5E/WycBe2rUgGdpuW80fKREPe0Kmjj3zyj7ZKFo+qdQ/yKkkGCaJn8
mlau+P7lO/ZHS1D7jU7QgZ2qPYAinFkalg4YSLdXh7gjO7PCLUx3dmPUZ5+t
K9JPZudM5faOUtbQkYcHLwGOiBajMxpzno/wszYPotXszJNczmU0/y0Fsazy
Zmsj68zJkqVZRNjbnb6Vo8/jtoM8GJxyjiD3gKdMBDpoi8+VAsSVKsLTSOWD
BckTcg/t6RZO/cvB3ASBDpKslEsyGVDiJ4gYgOkXEs8mCOtfyJsqOL3OYbxk
QRkHFqneYujc2KvPQRDIKxMqjLysY6suYby5Lp9AueNYSEjpIV1UsJB3BXto
IFcH2S3RT1BUODVM8PIoRI9+3kZmjnCQgLhYJdDSwQ8VK0xuBvY4F4onA8Gn
286jvA+Y3CgvItZwIECoS+zaS76oUZ0i8YmFhSo3syrmrGJZxImseEPslqxm
M/ETjhKBSjPMmqwSxksiT97tVatNcqpuBCyN6ddQQQII1URC+hlB1/Epp8qx
lzYveArMtWLgpMEqb3N9qEZnkWT92CV8LVbf+icTvO5ntGqV+zNjR5nu/Hav
1thilvS5yVdLIjGPEanD9vcW5iXv6fY/5tOiytOy/GfLwYyF15DuQSuro8Pl
MNPOUqKjX4fQ8a2mhtwG3qR8W4xiN+UQ3IP1PaZndMsSYdvtTs5UvwgrATEa
qeHP+ylSg6hJ7bB1stB1DNGm23n/qz7o0gOldR148u4tuNIz8xG9H5gYMxeO
sJ7v4pBntpo9oLXmbaCMDLdTKGqkmZt32BTQE3AWk04OyT7JsndGXUM409Qm
z1TJrywR+HKgjwP2sNKd2zuEN2qpoeM0uhFfldgVf4EG64fO15ep54YGbWG1
7Vg9lCGj9+nv1TuJWYuehQf3i6HvJuDwiHt1QwK79qnEQvueFC8qgm4LZLdY
tbXVxz/woknzU+B22StnMjmeUPoN57ymYYBXpTFcAJ2RNcitg9uetBuh4ZFe
ck5N4ynbrhJICa6B9JfCK1fglya5hqmt948L+qdd9ZAZLfaJNOm1PaMgPNRu
9iUjo4mFI/RDYYiLkWq1pCPtbc9b5EQwDpb75iO0mhYX1hv0Lpq2jV++YHeP
JZMKZXvj3P0O6fFAz7vHUuW8yAzbXecCwTWmOvEdwD9b+SUeOIOxrDZdqzFd
fTFfPwqt4TUfICbpp2q3jnD2JfGK5v94zFhCneKj6qnguBjRgtUsDVPpd3PR
56gSOGYF/rtF7OQwQabgNYmBLyqB8Zu3TwBwVB6DnfJqFX+p2Jcn58xdMmj7
ZNTOklFgvELqLGI2cDutnjvWbDbPxyDGiiTxcciYMRqZzSaS2ZpwLN5vIf6f
5Mx16gBXErdiuHwf8xhpcxob5D46TYdeW3VQaqwwsmH9idP5ZUcc5WAcUoua
nldSuQExANNekiuoCau0fTEM8C2CpzwnXdP6A7rxFJASQsdz8HUi9bsomtOn
qGXfE9F3T+o2uqyzq0rs+FiZ49cXmNH6CDmlZGHGpAQNwcVe9I1/9dk2wMeB
gBOBsqQaU36by8rLMlDloFvqmclpay7tJk5Nuqp5KowZ8DTweMjStuvhba4F
NBkc+iwBqLo6r2AezHBMnb0a/DlH6hXf8f2iQ2tk7NSAjvOlj/5iq9retiXr
W/A6qUj9ZAaAs0QcK9g7tZzIxuqJlAW+sav8i2RSUuXffY9OrRx+XmE5QLwS
s7hhy13zACjHitL6sLiFJvfMwiXw/uBE7IS4CBGZScobZj2C/8ZvrxgDiA1l
ELA1KKpvkdo9od3eeSoSKVnVyPgsoNvAe/T0esXMTmugf6DG0jt1jhDtvb+6
m1BWh0e1D7IxhzsVALfKAVMRVg0EVpo4N9vvewJiHAm6YUg/zg6aCzQxAYaa
4aGGdcMA3W8o70qQTHY2S0eN2vSa9FUAWkBKSn6rT01h4HiFYwcUL1VfweMf
kawYWsD4XVJAnw6E5tiuZ3EmPJNo3KSIyj19P0YUB1QXPlkB0FUQLD6ws66R
FWsLE5AKSXJLvuK8+8QrA/2FYiN4bsfNIzg8BTDi4/QSGkPy1sjpIP9aI0ZA
uygLj1RACB5Bdoh9I6u/LXt46/8oClBQCdgCvSTezPMOL6INxzvjrOkcQNcM
4uBp50NElDNTtAGkFRDrbPk/lZMzl0VwsXJ9FDCX8f3gz0So2Ggo6HtbAPlU
vQ/eAsPRlbDB3icfmaBPNKeifmqa2F5eyNgciG0vauHaz0ZiDZqN258cD0e+
FH/nAtWqO6Wfzcy9KlqO1hdjf0aO/XjS9GH+nnvrdGR3gCvZ/Dy1I5OJjzLx
jf8emLKqNd6WTqn7OjzAGNrjyTXPmoDoP1AHjdAHNYuFcmNRDV4VG/yAkxdo
jQFIf+AfmqgvVwtBDQA/ZVWCRmFFUwZs8m4P31Zwyd7djwW67r9xjf1IBWSy
vFgsgJ0KX/5ilVLQRLVlYT2z81i3q4ZU2nmUoXQbq43En77CFchSWlVDT9Jc
00mnVlddp6287726KGMIHbB4NotiUdaf4T7hB+pzqtVnXSlcN+L5+gByYU/q
PzoKQJMwRk7RCBGOQ0lfNJDwCwjA3UxALuK0Hlk4CzTPT7kwJvw8Kw7gGkIe
nF70zzNwDPHnYA0Qu3H6GhW1XhxTuNyZFy++NldEXA5Ec21Ij2Nur1OLF7HU
eBmV6fSRj2JxgfKBNdnBdkwvFEt9HDlv5ZGc28TdokkGtmfmtahrGtbbhDPC
3YWVa0Vd818keKScroCAgt2LjYJT+YRbg39wG3ZbBx87dZ9a27AMCkzZlo9p
OeMOOYKMLM8Zxia0u7c7ydDZxFkwkTC89wMnhkSMD8Ri8uGX1KHKozj+wnbd
PxTiBkIcqZqb99jQvldQUjEsUoxz0yABx12FBEridyc3WkguoGPWAfAVXhsi
6Vjk+fhLYc15yCH87573CKyFnmtnI9nsewZVULXd5Jin725303QHfZLoWlWb
W/yppkFyVx2hvDpTbshcFNgBBTHCcT6/XNEag21Fej3Qg4pJEjo3ipiL4j73
kaOljWaFY8qtrRD08oQwGeyR5JANzSipOs/G7ltSUlTPh9oSaECca4VubVD1
NOgyPwgAbaJCsTnmmYvg4EVbiq2dSaIieDY9BO1g8dbzk3eJckfaXuCtIZXa
kRrAd2IXXTU4Q5oeqWn3Anvk8LiylksWQqNcn+mH22v1kLLM3LFYyJYXuFmw
sajuirru8UHlKjr+FtWOlGybr06Yswqt7vP1rsg3sGeo4+bbbj79rTvUjVVj
2mpqSmhO7lYL6um6SZZ38bK8joI02ons7tz9ZFF3/JF2Hxw20XFrZ+pdpKgV
jRx9MWFnA/+I4nkoR2KjQ2m4IRQYHyWRI4uqBtdaEAek5vGzCQRB0JmD2xOK
EIsfZ0q/9Tp/OOvC51LaNyL4Pwg48vIk+GbCJvq6p4TtKvdDC7kQ5yf52E9S
2MosBr2EfnaN0buyNaBYifjTczJoRzSvjC72SpBropdM3qHfjajqIiF3oDpY
1RenfMiGh4Dk5MiyyKw5/PC7DYvzYFHLMEzQklxrABeXqezEodywRDs/E+Ud
m/9VLBz2Y7L//8ZdtdKVLK8s7FiJMfYnsJ42H1QsHrrfu5v86NP0PVKDFkUJ
+cdBQUwgGoHkugVEbLsiASZKAfvVmSgLkQ137m2saV883unZpbwy2/TrBrS7
ca9uzLYu5+1wMneemJOx/g4oW/hHw16BCe/u8ZCd4Uarwv3Jr/6gVfB2dhj1
ABmXFiJparMu9EEtPIaHTIGAxS1e8+IHisNkjb5N6Z8jb4O+fWzDX5COR3ka
r5naziOzZxWrfyb0VL2WpYfs9Te/B460QS+JNqEoay/TTqxi6g2Ai4tCGgOE
I+oE7DLM8M/WP1RSq9WgocpqwFCeDWhOZ4ZXB9gfOtEDFvF1pjzxMKcrXq8Q
DLCd2B4qFj32r6l8XBFsMDJCifF7ZHMANLan3Slw/S6OHHIgQEeaDHfjRiJP
WSbi8vPH3kF9AE4tOQk/ey0L8vUF71C0sm1V6ooVFTzv+PEE13e4wis2YQCV
k/Z0zjAYppeu/IHeJOX8EkUCbH0XSgCNXSE2pBDhGak7pC5mqz2QTT5njVIX
ibfuV6BVS6ljK/9BBXmNbFmXsgFa101lfNubEkiGqbjhKrl3+jiMKGcWrwx0
qf8e8Cngx/q9Ld6AcmtbW9xWwR0iAXmwwLCXoZIYFRmo8bSYHxqiamA/8OYi
ujz+IQei0vlbXW9SMZ7Q6WnBrmXtVab1DgWKI5nrQ3H2Uwn3M5KgOYIAIn89
wmrK3+TFxHgX8tg64uClg5Zza5BROYHXnC4cq2Z3GB9ZPvKBJWMtxtVJ3zm4
Iyx9W6As4cVW6IVtqj09yHcQRONkEt7hN8sx5W4/Q8Rg+vsme5vJ8avHaaX9
ORV+/jEgv++fqvoVHduTK536cc3ZqxyWZcV5UbwRRINNeaFYotHEpG3pUoQW
IkMbSyqR0AHxECR/I5PPnP7IqdfVOrp4Og3JKvEqyqA4hV1eWzhZ2R8Jcj45
Or8ejZSavgaQV2kthNVeUR1wlqHA7IF65kYiIB3Q4n6CIvKw4+i1tdvfsFM/
SjkzGiSgn0X5TmQPFOpwtTqPNlsi4Lv4qTyuc+zOcYnNQklLpCBc0XVrcHdb
exscT1doMpMidJDBx6m9y+3zf0hiI4PuLm0q0rcvPGl0rBayMSnjrLGIqMWD
p5XxZ5Sxhmto8gPTkmHer4n0fJ74/0klYK9YhnLdWqmOwjFYcsieOXpRsdUd
dlvqr1qZYAh1h9VF9OsjSSGretW2yc6c0+XJjmJJk3Bjz/NRd2CsH1dbLcEp
etGohboiP5zk/MhvbAa8BC4xyaQs6f33JpVGHxau6y1IgixsmG7gbghD9VCk
HkhDPIEZ0llTiFqegcVK9BAZWVN0rIOsb0kzynRXtaAAiLDwPg6kb1M1M4k8
jOj/Bh4VVBY+HTNutXWtGPYwXxlhrzuZbgRX6AWsxrb/tR4+EP+8+pwcJRFn
dT3VUl4OAXUvu5/D75CCRjgSq4mtjlvCQOUY7v1NcagUNxDBZy0hVL0IaWxl
Frg3EzZQHB7zgJ9pqURn/KohjSqpn/SIwAZwRLyk4t2ulJsSGCQg7K9o3BMJ
WX7AytBgp6l/RxN41jeLsQphryoe/gcknsF2nJVxoBdyJfoAbQc7pEdbNAF5
+O8PD56qVi54VWDu+CT1rjnfIfNTegN/FjDDpOMoY9PZsudX4iox2dk09XdE
I9Ckl8ZWZGeKkSLT4r3NiBiS1TzyjLOqTeTX0+7CgZeXi2WIm8nBLbEWjHcL
G43Owzffz8QeykZtW2H7oxWbT7tEWeIIGVJAYLua3CAsng1p9UQQkbez4ZJU
BBOOJx9YNCGNRDM+X912kHZyGJyS1TsttrNNdhw0ZBcphNk/hgX6NvNU/Jbz
PHxXvsVlJ9qIpFoYx1/56hdb3WTp/BQjxKQybNO8U/+uVQAdGBrO9AIKyt2L
OmhICUg1w+OTRsUOI4VPCxxqWBrdopvFwILijC2o+DC7FhqPHC2HT0brnmGP
X49nawoIS8n+pFuy94NujckXjNasZdd1KPwHCUprM/70+iWV9AXOhyigGBN/
r6wpGM54lh4W+mqH9QrPj7/xJCMPaG3+0EqNWl/z+Zoe4DBOz0/dEwDMwvYu
nMs7XuJoJUAL0QuKnFTAweCI0+dMHRS+VHf7Z2NDSSrlPMO7nVO8dZtlMMBB
CtVQlpEGLK1sxMP6tt+esWGUsOcgX9PLgpcS+yYrV2XV6D8CTzeYzTxbjbY3
AZ4JsS3KzawSwaNa7zHQCVq0NBraFicayYGoN7VTdiZx25N17qvLXM8S67zm
PTwMbobap7xOIyvrWJU3menBPPunF9zLyOay5hTJRPOv5QJnwY5EdkO6bli3
Pst/1tKtg1r/cp7QUNLfMXU+p03ppLPwN9wJ87zYU8Xr1bounjhN6Ze6uLRI
HdhERc84tnXcVcYvG4BPBoGyQpYzqQXIP01UkjujqhLrA4mfWS37yR5Dzp7e
vt9V+RbEpqENHPET5RdkjW1Ll0pmvkBGzUn87Xtb80LLVP8urFb/2v1/IKU+
l6y3hOXlqPGKPYJCeGB6f3VGfZqrQooXrJy6G1Or9EZEimwr83Xlp56UVYZw
8eg38PSZNmInfO6E4gTUW4ekVBXvXTRr6fU30A03YPNOSAroXh1Bk/h1T733
yC/fevnwYHtYGLGRRx+qWON4rFtYKrvroFJqGIMuHIz6O9L+z+6KTMV6GpEf
lkTasCh9BzUgVEudXXOFfbN8jxpQcpOjt3RIuO7Floc/SRrmDth5sOEyY8H3
R0NXd9m9+xuJSQU/hM0MgSlScVqpV/LMUR67gWKx8zux7Kw8j9DGVTtx4+7i
+O/RiFlgVoCotgF5a0e1vwcGrNBfR12KCDQ6ebPpQWNgDH8pzMc0i5Yku1Td
br29P/S00R8c6CsaaAzUmukmiYiM6tu59i1+MzN5u2LUxGlfB7Wjyq5+P5wd
/HMGxxoZ4J+ki3/JUsj8CWCi1O4JIERcTbhYk5lCh+KlnITQWM08Ng3IVSfZ
ZKBv0m0Pw77zBCo+guA1d9udsOknAJr3hzERtXVpkSFnsX8KHlwrha/v+C+4
MB2Yl7Li7fZxN+Sh1nR62eYarBasp8MNWnWWKC96iSmOouDlJMsk9gnQglat
vZLW9BTt06GBi1R9aPAw0Xqb4HCELXQF+lOenG8GfG4iojDD2Q3W8El7BTNe
D2WagOU25UvBdUgWlaiQHmlwCGxG3rQgVYmxSjUwDfHd7boiosOMiSDBImo1
mRtXCzDNP9JHaHiIF+A7Wjbf8H8m7PFlC2rQqxnrFG18zSYx+O3b7j0GZGS4
84O5H7oY3I3vrOac9YEsdpb5CMsEbpOsD/efqM8L1eSZEK9wZqxjrBnPgp5F
qEd+bTcYPnyW3wcNoh8MJfusCTU75emW16lqPR1iyv/Lr0sTRYKjVySRbnQL
7C54qvdgCt2vFFvZNPREO8vu6RyNUDZp1WyJRljchgH0Z3hXLX/ybdWdvUBX
GSW9g+y+SM3yyephWvlDf3E6DAOryJ/J8OUaZYU+W47Ap4GU6ZGKFlxgNA+l
0hJd/1Bdblg/+x96CKz88ulJQIyXMpQ/cXv1FbJfh/HQvGuFudX6T4fsC97w
Ym1mD3mDlPalE9sOMH+GCwxHj+KI2kaowEPiozutsL8QlvhMAH7YUvxmNJ0X
pQoobinQftq6A1pb4hZ3g96xlZ+eHdKI/8fOZTfRWwgi4dtok/zIjeqbn6sH
NWhOxpfYXC6j0OfmTYPIM6pCm8FadwNxF0/64Gjfi8NWRNXRosYaeSxqf34G
JPx6Ryo8Sq0DeIF7gkzZHLdSDo44SzKVOkj4ZsnVbGoPaZK8pxQWIUZkcTri
IsfeGUOWpiyGTWygHJkqDHF9zfUIxfCIWy7CQQjzCRFJBlhWY2q0bTfXWSHs
yZg6wonEb7QMIM1rkr5L6JferVE44+s4UiYlMN2NTXr5QJc6+S1JB/ZUlObX
sqsZwwM4rDg6298p/98224TxuHiW9yfe/1H31OfqeNs6+xDrysDSFact+0Yp
IVVhcXDduEc/+1Die+yotC909wXmNUrt0kn7jXKEbdrCeukAPG+GjVT/HN5N
Fj2is0c2Ss4toDFo+rMPcs3e55/qdvonyt4QB1pFJeqCtSOc+CXUtNhW7NND
I/TL5s30r+4dqzESYOkDJ8sLYcBPA8XCye//7Y6XS8M6olmA6KYtarN6iP5H
d1Vs15bf5YhM7pCfIPxBl6A0qg/18Y+WszHAbfZWTX0PwgKfvM1OEg20caqU
jiQJh0h4Ohg09+/LA8uoh/OZBpUTlle+0BMpLYb9gnNe09MTou29qDiLLPS1
+3z8LT1eKVbZOEiZuA4ig343F01dY5b91ixtpRJkrhL6z/zwvoB+BcDLTEg6
s7t0tyj5xuKT1cdCBeWh1CS2D6zYkeyWIpAyGN87SSBYG2uegr3jtZ67/ZPH
jot8MAqK1lWWkqXAtppRQt471g5Yi8ZqTS4C5chw6tI0dqE0jnsEFHe6QWHh
aMdamCiigGXyAprHQH5PKAK0Nd03GaXsitzFisURJns5CSoN/5lI2vz/ae/l
FGxey5TnTUk3mQ2MHewGQtF99LqTWlkQD3+X/Nsu9d6KlhjNu5FANDj/Puf2
wToaq35XqAJ24TO6MqvMWz3gDy5ZeO+BeDflPteb6xzzTWJ6GrQx/ZQbZKMz
chjt6pNgMnruKdul09baQE5sHeUywagX8XZCHoUvUDR9hkyUQ8OvPamD3nxT
/rjvdoBFydSwzxl0l5ttHQZCO7u4OXSVEuE3Cczb5w5gtvw7Rcc2/t0Z55Df
kzMNXiQMA7SDIwq4oKWlkWW1zEwxbe+6Bg+3lzsifh6dQA4E/97d526N3H7B
c7apkh1yy6QZhTEt5qAIAjgAgJEJ9TauLd9xpXm3yH82uZV45VCcqzCz8yYn
FFztliC723TRFdBFRi5P+ikE0SJR3Nb9wHJ24I9uwOto0UjLjfkojDnNgVkp
k8cx9mmm8N6zjNP5JVb9R2nIZ2CJstgP6U3V/4kEs/3hUgCn//8m4us974Fs
zfM5PW8YCMpUNzJAL/kBjGT7GcMUi6HNPhxQscNfucKeo3u0j4E9QHFlnnNZ
8lW1ooI+yypiHawvdmQEF9q6WsgrxVtHy5RH+Aho8S+aOgpBxUGvvpcVnvhM
drxcOSoyvkknA6lP6mViMyh6Yma+dUFmTn9auUhBUt3N99WFiHdYF27eLO2T
xhfgTex/QbSqk+1lZrdhdTilnJYX8yKFUKfzpO4TgZOLlTYvDUoiWi7lDZr5
rQYGq0E9txfp4rFAEwaosl20vBhqnx5fs5WWxPcdgb5JwLhoUhcdO/jGHhLv
zPwu4zbN8+t13xeR8VyuCwoO5ezye6AE5iuI9bGgg+5xDlBURpVdQOBPWYU2
YkpfHq5OeR6fshpowExlyxM777+/4D7Cbp10CiskdZzMxRbuUrQ8J+FlDYZf
dhQIdGEL5IkcQKlA9mUtwFO5uip7xRAjZVb1guDjvTZ4ENuoOWdvgeIoUQKK
BCsqawpQtTrmrb4+fZfv41ttJU9FillXqmZoiP/FVVSXcRr27sUH53tNEny/
zHSqJ3QwyOd9iwZrvq0Qx2QnJ8QLLwp+W5sLgRYDNfLCbrF7mYTZfWTZhIcG
NmEayuP9JC1f22whKPeyxfg5ew0LLkC5lzPkDO5EQy1aI8QnQfS/4iN++L4v
MqdMEQBi+ju5kL+0wWQQBwDs1teBwTpebM5yISzwYujJQcw7IdMuYWETpsxz
Tc8F0A63BmMRLZwIlULCEnJhMsB+BFPayo6vdLz3q405H5DwnFRj09HyJG0k
TXnFhGPuwI+j3edX4qoiC4eLdm+SxBcDvKjXlGcMgCu/2acLB0smvl3bVRyS
T2KkudBLwnLTY0sz/gsX+4laeQTWNCMSzYlSER67ecvd0er8WhFdvT6ZRRRq
vL5VK3i+Tsrx0SbpuUCJa5LdpVKQJPAz+PJgfUg/5KtMUsKH77hMNIpHWBH5
KSqNjEHjkVp839CLR147P8nKRZfzp3rgvDTfOW4VBKpHCsBU8kBphNWXjSIs
XEXgqvPMoIw7Ae1DYxG1OceDYy2yg8puOZKRRwLjAyKAECT9DUcH5mEZOTNa
zgZ1hLDIhWCp0q8NAsxmLUmNb+E0aXFPVGqFJVMjEaj0VmOrQCpxEhliPuEg
ss+nIanvgYEYv3NexVRYenV0b1Pujpf2T/ia6s7Lisj/KwTxWJfGbwFnpRrM
T8v9U89jF44E1Y1KiCyCN3q0JB1Y5jIE/iDybLiNcPwgsdeg0yeCQ3r8J0Sh
De5KkB96uxscgMLs3OhFHzNMVOaU0G2mFJ4+s4F9Sfc2FUYjBYYYYw/qrpM1
Q+toXnjPZI+0z6o1nGJpWM8go571ROnInpkWGfzs5+BiaKJbhyXx0JSvjWY9
22zhAxhnKN7ywHpZs1GNmkFkXYxVUaz+Vi38QPtIJcVjyq+iIlnMolfkZgpO
Qo9yjGVL+wb6XcfWCU9tbogT9bjToXbvCX44hDdO8oCHFGbXVWunXJIzn0cU
/ZckkossyBq2+DwpiMHx32ZuD5nCU75wTH6QLuA5kIVSq02jvMyZl2ohqYsy
P1479cC6DmKfkloT+ZlMrAXKfQIALrjmSGOPdfZTJApfUj5Q8YfWxCsdAmiV
u/v5esEbX6vwRyLFVJqmL8XIhw0mhFKXh5ARc1JiZW5skOv9Hfl2LT5+nrRn
tdj/6ymxm7l+TBgvHYGCntVPN+fSbYXEzw66HnYYYLPrB0VFriaPm8fkWnoM
S54BW6fRQSUX22sVXxi04fPQOpuDHZ2HdV9nBLKozoqA1pvSi0y9U1yv9sS+
eFo2hRjGo4xDfXnCN8ZJgDfIsaHH33kaU6q9pCx4F+WeYqhFkMY1GWD2hcQX
90E/3lo5PP2UlSsH4wquGyUfz1lKJ7ud2Pen7KcUOYDdRBsrtzzAHmDpnMi7
KAPsG5MRPdOrzpqucl0Kfdj4iFmT6DtAzghjRGQl3BqEaiSy/yrDmHhb4ye9
FlFOLedMdNb/KoqYvYNuCdnelVjgNm9MDzSvmhGUgKhPvjTXBx0uF6nfiVoh
nXLhmoFSODWMPSfMAvGbnyUaGw7m4P4RtLiT/1IPsVSFfKQWDrmdhOclkUuG
Lz10xmKpKS2tiSowYW1aZC1RK2yb84DDJ2a2hD7VOU69q6DS/Cl4sMNtwcz6
V+Gc51SP2kFalYSHfuhGX1IpXBKRhBbEW/efcxImcqIqj/6CAaxLxkRjyFpm
rybZYrggkccAdcXnlpShCsUEjmfLrgRI9F0+t3WaufLBV1w7MZ3ECsb2oSeG
94OaW6Vwu8/sAvo07FquQthRSDzqGxmJUZ42vvo/mwBcuUviHRt1E+GkafWg
JwINHO6ggrWF/EDLFmb9SY1qnS9HnqUlK+mv6wtjNf6gmqjhCFdF8zgFUYZI
xMJOEL4vOePyffMq8tYVTbOoEW2tbxXDQXd2yhirklaVS/ybnXNYVVEZ12YH
bN4IEfFOlAb0LoClYujwJYOcmDqAg0pj+qXE5xyqsAN4BYVopRupyiq6xDCP
LQqRu0lHdZtH5G7WcnXV+R1j7thi27QalaWlTop56qWBxgraQ24LQIhs8Gvu
7qJc3HI+JxaUsLf0j4T/0LEjFX+Otw7noEBupzjXMSLe95WLP3sU3ghjhosM
/EELlIX4cbIFIbH2gtCKtxQS/3Atz7qijtStwLXTnE6UxBoBGZnYXD0c6v39
CcaObXbLy8PwNT7C0QtzlhKkQN+VT82b27CxIWUg5/0v/8T/6QuNgZjY82Ar
gpNJiCeQA6LuiE1UrkTZZNFGUwE1UMdDXwF+WEkzDC7sau7DkHTSYzFJrDmv
V7ss0mSmw0o7V1i/4Z3HY+PWEdY/nZE4iFMX97qwbcbY/Jg2I1Do7kVajqVp
F+Pj6iE0wrSgaWzAuDS2yL3crZhAqcPykVfbvZjhPDhbb9jUVQZrsc2Idw01
JtinU+ZtgSfG+09w+gPe6b/17lwO52/dVeKjQc33XUcI6qsjaApDhay4GqxT
nyuuePG5hEsZ2BEw1Zwi2/TNFelEYfT1ycD51/TzIQuHzLs1BB8St4p0I/JE
zMEqU/EjzT/k5OUZq4Ky71hUsB3zE2F1uIw+wDFHydSj6QILOzLMoq/6b6b8
cMftbZY4EddCh5IJrT4O5jxVYJonFQyFbC5HsxItixMkFIMKEXDO8SAurw34
21vo1sxaI68aa/TZ/NbEsUmFSte0E/wco6rU5ORJKutDPC4rraSqXDvMkbNB
kqvY2EWDlXMmNuK98FGTYNWWZ57LT4VBIGw4w3cKb2OpHQi2Q2gfMLu7q9Q8
98yY3MomGX1wKEpRf8JsS0djAUWrShF6u2xFFdTvLBnovWUeGeDlvpNpNITi
yhq2JzNUtZk9cB304ggh1Eo8ngbohPUlw5rAI9nWlkuQhGOXozctip7geh2/
G4q/3673xvL7gfc2J6omUYiKWLtv6VpYfcWJHf04HsY71pUvnOWn4t4eKHEJ
2GI3KCP6Vp+ZDCCTXGn6OoSn3DMUR93pSU4vNf+pYZkGX53D/43/zaFhAXb3
BJGsp+PIQuMZumxGg4HvOBChhztXmlKmuc8bX8hKdh//jRVzWfbHY8/dHcME
uLIPaAs7lNGr/fRYfdxCQYlCoyl6BhCuHaGQNoRB5VuvaW4c0c3aafC7T+QH
Z6AeEDRKtS/XHISo/ajxjQqUfFuw2gs3H4/8m+Irxojkw5agdv60NXTQEqpI
P5k/Xa9OCeUOjG61erXMSdQNujGESaNQS8nskMrebdjgsAWBoV42/0x3PCWu
HdbGKyaeX6GOQmYXSirjqAzPselKRHSRYCof/wDuQ4BOvz4Q475hFH7SwJR4
+Yv16vzCaxPbBpVVSsJ0nclTqPwtKR14PSSCOO19snoJoGJbODawcQrWvQPZ
4wzRf6n+L6Fj8ECQ/MyJCP7bGRSEKKc6kpe06IHLixJ22ipXgvMheewqKjlt
3yLuNal8yxuo1BzKkQXiQ+lDOcYr8j6u6Ry99oGZRqBeO/jLou6O0i/Jl+Sh
XvSziAzp+DAhhuecLunXnXEthvu+4S2RjN7befmEqBhqlsteGcC+MJCiH498
xCNDtGkcB1+aSAQik0zPeQ/l0npio81vNsIZi1hbr3G7VCAm+Iyw5Gyceill
BZmV82/hYrUoIMvfUsTFkSdGttAm7gat4Ae/NJMJuAPp/he/NHYppTGtQkB+
D+HeqpIErUV3A/Gw+xt3eo8GFagAvcsJqe6zAI+iVFzivotVaZubL2xwD7NO
4oFf4WABFapWj47JD0ImfSQ5p6OgweJ3GJUNnQiiCx1zEyh/FFwBiztKAnCV
K9Ukt3AhxsmT8hYOfQpFBQ4qg4WrZA0w/n4VYXM4mP3U6xzr/r6ug6+kmc+M
a9MphH4+YYVJ7Eb1wNUg47+2jeFVBOWxm2lMCRWJ9JGsUq/Y5CbK91g0Jzw+
+DAjre/lnE6u8QaYyEDRQ3PvXyBc0JJDBZNnCs2OBgkBGo4D2ykEwbtFIjJg
/u7FTS+8UXEpB34VqhBKR0kqc4t126Ojaj95x7lN4kXlKU425UCabDLCVAly
LxPJUji7SZU7tKFSxXZA99DGVMx3x7rm7ApZbrlfAiqTnYIetyTvFAnwRSn7
VIzOvvHxteIIS1kNbnEPtalZdygwvA0bW3HBsnC9+ADSgWX6p80uPw6lAIeH
be0iAr+Q268JSdV6dct7blPXJ4E0pQas5zlNyoKZF1u1ijjXO1Txm7AuC9Gp
X9/Suef/1Kyyhs3FV1j+VlhWXAxYsYLeDjV1VWZz0GIGwNGtwbhMsdu8b/8N
ku5oC1qMGHq4nG+OGHauRUcMtiIIj6AU+Nrfi81rPcmBWS3WC34dHKEBgKkS
kmDvRi1C9T626FMP7huFmuqedU3wAAx0PbfpZ6o3JWH5cfJvCjK1M/t3wDEb
IHDIvQUcpnuaL28ZmoS+g4r+7Z9vJth7zNVd6cpn3EeDe3paE/LJ+W1JuV/c
KkByNekjpEOuUqPMuqP93ggzZaBMdel86JrwSWzzGWHyVM2wg+gvtn5rXCr6
/6pMJl2trx9mWYR6tumQK5FlElAROmwBqCE1Dax10wbHRh7H4kEv6BoH19Bf
0wKyFiTpAjTeYi/nR1jG6PcEvYTt88CW2HuohQb1ykiEo5WrfOH3AFrk/Vnd
UptVl5XKUmHE05+JUZbNkT+NeOs67qev2dkezBkT8/Zkmdwp7HwG6WWmJNPo
+fyaEZit2tvOcdh77izB0dP4dSS3o5ue2ccf+r/DcWdZFfYOgMgxEPdd0+Ua
1oeXRLYVHfbvu1kdnzOHZofvCIQjVuKeTqKoRkdYYREEhKDhXGHinwXP74Hk
mFlZI/a/ZXPZHWrUAnz2TQOKVgjw2vmjhlbohZJO1ci6Z0j0siQ0ufmMJhOJ
30adzQdnk+QwhFcrAtisSSGXIEWDQCcvqOIcoRFNE/BlqVfar5ZvCB5LP36x
1remv/WuSg1o+gbKuteZfP03iS2qHTVcHAJwLX2B833nlJtQAUhSSqOyouXg
SLp66zFSTR252nAojuKxJ1nZGvBBauD5Mg9cDfbNeYMCf+mywXKZx3MK1OH3
rTZHmZHPIYzhZoDAhN/p8lDuKNLRn2JwimThLQR9WlojimZ48uxTHklSQZZP
lJbEBTilRvSJKIJ9FwqikG68mynT1Uq4x0oy1ooWAvltEa1d3KlAGAEZT7R1
unlfW9poudZtxkUsaMCA0aPB3wzBTn1mTPIuoe5qdXOEjioEe1bU7me5ip15
2Y7fjX7DyiXyKEXg2tU2+go8q8fRCDnSGShw7LaDfk2XbjGDGM/AI5LidQSB
R31ThSKcfOXyplsdw85ThJXZJW77AbpcP4cM3l9cpfomZnPXtMMm3+MqB0hf
Msfpv3tt2IJCl95yAUCh/T5yNYLhiO5fYi3uo7I+BgEzlIgSdpG/KwZIsTnp
xZ0a3l3uUEOtLE0hQWwkIgr0VBosxO2YfDQ5qM/sT9JiFfo4t5dxIN7uqjiC
J4ewWBGYnRQWAOxeCmdVWyRq2DBiUg4M42O4ulqRl9y7+NHjT2DxNL39255+
25Rs9J8eKO+Pn2sCjJCH3RKgbBelGr3u/gqysz/xR4EPBsGLBVk+hiyK5ObF
2fQ6V03hzEWQboGgROWvBis/5qHqRyUQqU7OPGRvPocXIfSXrhPQv8oTLJfA
YeXy2cZe08/vnkGNKnNZTI0zQm0UXUxHhSfw7X0oRF7DyzOK56/YxE45kIJa
OVy6eE5nTEeo88BsrBZLjeV+ap1dFbuCuWm8OsNWBj6NBkh/JJ7BRuYLCuc2
SBXTPCrAxNAEasOALora8Ln2URjKSUlsIc/FPBbmxJYFdL0pfCQ6rerePRRK
xcC5AkJtYqLeRPVDy6zCbgHYidaeFsC3TXSlyMfmVy5bJTNmHrfbJFRC1NDP
ITVifzlL8g7itHUOk08FufJh1w9UzzWtF/Kko2Qlir37trhd1EobJ7kYONt9
Qvw7Jvcx96WSpjrLu/B5H6uBwASi9V5Lx4XnRv7ubhNvHQ3Vy84NZRgAJsnP
owGepHUu/V1CrXVW19YJKsMUBfmI3drJiXuom+Wu3QDKXXKBpMX5JRdHuqcW
t1VLxuAd/WRV8magV+iv6i8zSZER0gFE32ngu1lVSAGl3rhD63QhkrNkBhU7
IChyVn9Ei4DZArW2lY02BCQ3V4Ou/WaGHHKsv3aplwnMuamgs0340lOBPMEk
hqP2d+9O8A8NQtCMdqNKDAh9XyKjZjbiNr/JPRmwIQKppD/Jq8oOI/NaQHyW
AH49ix5HuYFSTe68fTqq2S6vbnsVGiIFZBwOV1LrL8pyW+VZ9uUyCAMLCMWL
7On55lbu+XorQoCEErrGkuEGqBJz63UDGa7QoGx/L5k2On+TNk4M7UdI/i7K
oihqTFCxNoibF7zYbhmaA4kFnPDij0ZSEn1xbIO8ugXw6fONWujfDaIYvfwQ
/qxdEOfMcH0HVQG42S36HF+5Q26q7iQG1XpHkStjap6O8iPhP7RjH34BPGDv
ebEKYuimUgK/DhjsaEPHRRm5ZJoivCD50qaKQY54zW0KvtrlD2OM2JV1GCc/
mSC2Ge+AyGjhWYGn/OpsGSR2QdAfAdrQz88i0Wchh0YDCfc4OKi7CbjM8rY/
RUuaWqs8OSrwd7QqD2p/9kfsDlmX0NdE5nDr4Dpj0APF8lVjGlAoc4E2psXl
s12ONFrtEB1f6F7u0jXEME5BzHsYGDTg3kW5v7FwTIDnWma2c7b1v5gdkrJY
NMPU8rndszuVMNF7DBiJTmxb1moSTzqrwDO/IXCp9yshw0lLMtl/3uItFe8v
dcN+O0G0g2NyG2zoDM54QtFkiM9aAqdDvnxinj2BzGGrEdvO6k9j+BfD5LC4
SfFdJhaU2HFJ9MZwgdvH7aHpePxyKupE429BO8yLnM4L94/eltb7kz68jI8S
+KXs2+fcHWxgNpS9lE0Sasb5tfVR2vwjFWeVzWVenqHSVRnFj43J

`pragma protect end_protected
