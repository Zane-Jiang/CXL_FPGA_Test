// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
n39npMplT8P/VyDqFeD6rMgARpeeVQImkrk3n6mcmQN6zZdNSmgIlQHvka0+vTOb
Jmt/kSY+mU2s7wsjlWMx2WdeTbIcLbTyYdTrRmsFxL7pxRN2uC7CQxG6joRn6h/P
OVa7ozZx5oaIQgt1u6O8LsP2BHcHn02rR4WkRfr2eMw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
zQ/XEyXz2j59h+VyAn9xh/kaSrTkgmlXqehCsxT1LK4iJfheks9La6d/+tbTpAN2
C+eIRUmxclEfKaVpqnHOuQUpM6dWrVa7UgnmvaTPp5d+kwT23t0/cCcgiETLjmS3
52JE+JJMPNFRG0g+AIVsCKU1F5RU5u6UbkntqIOkgTwmwA4Gig4FKVwpsMTJ0Znx
nZItld8jEmsxodvAXw0aX/ppskUXq3zLmvr/gzbLPcoHExy2H60Go4ucg/6plsi1
Or5eOfHtCCZWMubTgeNhSlCVv+BurRmoTTs9pM7QbuWM7qsCRg2lOKVpTineIIz6
EydbZG0JxDAfkzR4HYG18lRgY87AbrHB5dS8n7SK8vhTthKzEhuAW4sksKSMWVMx
/gss18CXytwKEsdXHzWziG2YPM5yQQ9xRi+OWI4SYfL/KPvI9511XqPIk0eNEOE+
JmQS1qU25Omm/TZxWNxusjMD/VW9aaxjQ9c+GL6FBM3NCSoiv66IlpQPJsNJCUzK
H7y3OEWjeJlDJ0aMka/67ZUDJIUxaXwpy4JZ+qr/GuN42M+9d++F6uS2OeH9YCS2
BV9xKhFO3aMhlgWVN5tHHwHu/+euXEVX5Sr2P0skOnxoyUdyu1FFCwv9TXGXdeUV
wvSOAijnuIspIXMLSZyAnrUk2qkhYTI7tOBA5KjE+RkV1Q07bdjFqKpqAEmNpNrM
R4X9blkCHGMLMQzvc1f3OQYoQeV0jYks6kJKY5a7UjVaIJntuAfNZjNNrdg8CYU4
LsoZ3R9n6/5jH9DyK2HTzroBSihC0P8myq39j9TvpNxIA5tQrSOyYx5pkC+iMLRy
g1iYuNvxstzB+m8mxoP9PpkV1pMdrxQxU2+5gx/Y8Fd+jIGIh3BSV6QLGmYrpNCT
lDdgmuWxGVF66g92S9aFlYfXVTULQO6YuWxBegUZwuErfJGoZhtam23XH+CLUaYj
jphf13YTeu5MwafXOD6uAaZfQHujIxd9lgvg9key2BFskaFjCM+unMDdr93BIXyC
5oD7lwWUfCt3wJAdCMOLqESzmw/heZ+dcW/FYqWvBwN37s0lSjPNj6r/GHIGyTBs
+JAaYnPo4vgbMLCNQ7LahuvcWWw219RG7DWJZDfMEyfvmSBkZQAzEUzvWyybKd6y
oJ/Kp+YN9lzoHnZor5PMe6GVGaC7SS6wj1+9wtwjtJe8SxxDGtsEsoR6RVgpud+V
wlwmFjoPrlWFwGLd4A9nA8YygeejdgjyoQ62SvjTQwfhvLqgoA6HboSD8VYwwJ7w
SceHoRlrdteOwD7DQSsmXi3rqp+UVI3E1se4uEBwAjRVPVj/BGkoa7OV2DMqLjAZ
ZK3CE8hBx1t3UhJp8Q4T65ffCQ2PfwU8iRmzWDCh1FCR0Wju79dieTTwtqpspsJW
VGO3v/85bW6DquDs3on8/NEnDfLgJj/HOptzVEVDoI6q5ESUKX2HmWMNgahXPNC7
amlospn/+gSAlzwZc6/YQsXH0l5wthPEtC7wnsrJdjq/Ndq/H1XNI68lmkRCyxo0
Uh5/znaibGCFVn+ZI2FpwGERmI50pD7q+s2A8idWHSwbBngjPrBcVby7J26c5TJB
muWo/1p4RZRs0mJ7zyxgMrGQRXDRspVkvP4npFZI9AzaDEjOUlkLYFIGWBSc0llQ
ZfN5FWwAPQljqnvH7Y9XHR/JJ/kVcByI9Tr76+8XnW9GrksGusG42SZmB4mBWAvw
QfuUPgUIZd99A0fApPmQqBwZtIGwhzbKkoZvhYs6VzpfLHjCdd5yA8A5Bb9045l3
plVkjrFMHAwdYBAgJJPiVMn82yCNGqZ3qzidQvZ/wIqi7CcyKVYoBFh9Eq8LFFie
YKGR00q6KvuWWIaPXDPsYqHA9TPVoIE4ceu2NBDyCNLGnZVcTRZhLRFPG3f6UjKs
P+XiKOIqx8aMwniDvuopIsAfKOfuN2w80B+ePicm+UJBc5IL9xmAdSW99KDQW2Su
cLUEY8yGYUj93f3LgSFtK0sfdOOiP8sosZ4CNFzjPoKq4ueZoBSxQ7IwgivkX/u9
T0peV6obDIi60x4T/vdhfREjB6NjNu1Ny31VIHk234MBz4q6cw/+7Y+4l+jTpzzD
Ds7OURQYf0VbO3QDCQnIi82czMqp00mcRiyRSezS3HfefWRhOA+EDbIRvdI6x9G5
mS+cIrPyNtfSjLdvODUbo0ob/APY0dtcjtL9jQ8WAKDx6cWbKofwNie2RvTZcOTs
uYLoGLM7PnHK1230Z2vYwXAEzdQ+rxng2oaAgkicX1cy+GAWy5jfed+XuW3MqMTW
hyVtEeCPmkfrWd1Dsh/SiHIWxsvwjLzJAj7Mzzy6yQJUu71r0BL1PZwzXMrYMgy6
dTCRqF0sq4RV0PnBkQzJAhHz/re5p6bW+lKC+mpMRpiVxGUS9VmuCrf08cTMhyWa
eYXBPefDdsiEN0nMdtUb99C82SiVtacAP72vNJkPFVEn3EPDcySbr7UBlgORuZHb
Qx5JOumm+aUa5UTVBnKbYbkJQOHdoV38by96IMBhWrK11X6yjzX47Ks1PhmwGNvC
TholAI770Yc6E5worjNsu4ngonbImhRJ2a0bwAILpap3FB3qkAXe6N3D1GAQ9ex6
BXQAmBqvHj7KHirRQ576lzBOh9sCN56QoLUGADUOnNQVgmqOHlKaVlnsXvQ9fr0f
B07dQMQ0MT7ZHdfAv5KJO8xbdO882Rd0bAIBoXYLFhN+50vifNhmDFDvU/A+Uu//
isW+dp6cl6RPytQ6s2z+NNJg4tayQEUoP6YmCU68XOlv2z6PeEFYtk/FXMDauFkt
BF1RadxWFnMv60/ABzPpCx2p6o27VwrTb9furp4/tTSkzuCv9WqlMVTJsvNEbKD+
lLOQHJfepykEmz/PpiHFC16lPWtQcG/tN6SmH6TdnuudqhLJeKzjJq0+U1HTLl9K
5C9FKYnM6GsiwMysTSMydMJQcqf4UEEe0RVa6IqE+Df/uU6JI/xqFBK7kQuLpOl1
NNeagOeWolJEokFbNX4+oLtjqpFkePnfSXngBtcEG7Ix+yU+siyZudx8ItrLSVHj
H5P/wgQJn/7uQonlvugtuvLe79Hop3qILpk1EIuJhM9CZAO6dUuQJUfGGgPMRAm2
oqWJoewcCOU415xUFe56KNTPNUrcF9FPxhxJ4Ppdjoti4aLEDb19gYXEpc6GFGk5
AaiuZsAiuYg0z9zVxOU9a70wsK0xcXLIQ5b//Xrp30UMid0P7I9UpxmHQX3uIMsm
8ktIqcr6qFL6rEr7fpQ9ffsKR1VA9BViDDuSV5qlL4YyaYMvLknOSBFkeBLhzJLt
6nQW0AO4OiK42tXMJpF75/2LOBE837r+pHOX5aY1rnW3Ot9u3Yy+6MnHTt76udnN
u87rC1nnsVCjdJaKTsLLPW1CHdjfgfKFIFL6FYrbxufIWGfTFRMvunzT5FzgT9Y7
VhbAYSYmX5wkrDl51dAB3tLYiZDak6vyp5RhzyvUhlsSlC3nh3oCMBZ+l74tB81p
87JXI3FvxxkfNTG1sCsnMQw2liveHvoRO5rVTcbxqhMCGJoce/P9KbmTWh5Y2TvN
sqmN5WUXnsN2vRUOU/+7mSkvS9S5NjID00FtS09c61kAmLalZ4IL86DWA5zHsRnO
ru8l0khi9ntP7iL0cGfkfESq+WitpfzKsdOt46SyTtZe/8jiLR/G5cIgNv9Zl5mm
g6F8Ldwq2ELGf7Sbo1jYDnqatRpZUCm0IV2P1UdwT6Jv2anMAo1caUWHNS/sviL+
rfrE+UuUOmjhg6XTsjka1VCLupY/XtI/yTlieNSj1plg43IO4KKh03CcOJyQBD6o
S2GwjVZPG2WJDJH6jAUZCVifTlPVmg9gzVa+zA21g1HYd6TUT/I730e+/zQQB3Ip
OmnaSte1Z3GfRjy2wgWqVHWjgUxWqH1pMp6BajaAMK3o0F1vPVsr7qHI6As7M5SG
8DnHKF103SAjicdORSo+egTlvrAnRUY7jlYIZmkRCEsBo+djXhfgGHZXGqEmKlON
AcU4rrQICbq6lUegZ0+EeRZMmQOuvjRHHy2Ck4yKWHGaG/94tAP7kAN47+jPjgNi
ujZmK0h1lLcx1IY9QJSEBk40TolB3x8gNXb1T0vClY9pX668BDLQv6qDMsGYj4RK
Xvb0X+3s2HCPqA5hPdNa5SrWOOlEdCepE3MGMuA70Qnqz8ywNEKqWVo/96uYG/+m
286O7aWcksLCKlhhjjnmVh3oYcdO+he0ooPueY9eFk/UXlby8vIj+h5rISx/67Ok
H9XcRj/0eam500GPXhMMCEVFjxrMPF8MiZ7uvO1bqBYVrxiF3TuZoqsil09YpH2H
VA9grsfBEchnny1MyPGCGqRZvN+ySRkIVCfDr6wNKI5jIQGz/ngkxzfD6fxG7Aik
yAx+IOkGtNI0Of5AJzzwASkGKKLyPi+veVWSg90SywT45W27j0H3eIoMShMgIofb
xJNaB6VRUbxjHtaisXVQJymLRJZ7kiF0htXx87kqxdQ6WG6p7LN08Fhht8y3vx7M
Bw0ZkvHQE9oP2/qs3yf7zkjTfZUJVPmhHPL5IaJLC4/6lLv053/7Gre8rVWumxT/
BdpmaEobwmr30ZVssMw3ZaqbULW8UD1UlQp9dRurxxIm11kpeP5Chux931WTcYBR
U8LktytVHZpUD89boDk7MdOUiZ62Vihhx+CyKwGNwe0L72B9C7lMw/VgTIMSw8A9
Gry62JsnvWuMN+dejDVi+LOEma18E1sgD4e3G7FG2rEUqRAAIMalL38B4tzBe4Nt
6YqRLvG8ASc8rNTXx3496tTWh+igspEMuIjiJXv2KK+3ZwV/qGNpPkgpLLGd1svc
Q7T+04HRm+VReaW6Xc7NuueY6HOJSMFrqZtZ0Hj0RQu4RFqHi2roNJUqIKrbOA1h
0DUKN5t+l/L+uB7jS5B1mKsMW5Dzhdea9b2AZ5JcbDxiCS96PAd9TxpE5H976HjS
yHNTpcy/nJ5pkRqfUoIaCMHcVHYI7aOcTuEY+tGc/lxw5B/XLcgsJO1Nn7STBdpi
vGt+SZEvLpGS/hTqh39kWTV0DpdAFwYvqLweYBVK+1lENNYx3XgKjADzJnAgLfjU
xRlfFnQ0+rPjIV9pqXW5d2VvFrtizLWvKwwOW92G7mhqhGNiaAdPatlSlUb5IiV2
tYtn3MiFHpyF1OL9PM3D9y5JZkT0tSXF188AbNVdMiNESEnl37vbJG/uSzpfzpnX
vGJHuUmDO5lsehLEexRhvMUltF9LxM+GsWI9UvCuMth30+8xOEx6b+MbdZCym4mk
gjFSnYB976iiElwjdfqp5/pjESThufzjE8MffVk/GTTdQ5R4WcZzVZfJNpgj22Kb
waRj1+JIQ0HdLy3ZKxbNxWT4/QTcVMIFFsLSERGJGHyupBvf8MBc5ZSvLTl93pMs
35o7xZkyM76VuZd0s7O1rC9/7w5W3xeuJVkz9PuEs4zevcYrINbm0KUmSj6JN6JB
CJEqOzKGFAIYJiRWKz9Mq7+WXCpleB8wRdrxDMaGP9bp9xt/Cp4ZxQZrvXC0L2D7
s/WpCnQ4ksNCUwbwI3B485E9v/L1XlGbMubxDyzSSnsW7Xxv91Xr1eBUZhCH3dlU
98k8pwRsOS/72p9SobcXStliOky4xB9y7iylKIda9iaHuvmZmaDZTJXwbOzQN8WZ
SXc+OQEGr7rF/73kBNo/CT7mJUMdN5hEY8VJMDy3S0f6QTbtyF7KbNO6WWyhXEZF
XwzUKvwiUAuniqr+B0/amPbYonxlTtjEnMorwUObBPiDLCP6vRfEy5sfqdgJXjXw
tsYH7JJYjGx6poK7eSPWWd32zkfPVmlFz2mpxUKIw58fTiemu/5GpzmJYB7K1udQ
TLl+nCg5nFZt1WlpS3Eequ8T/Fy6ewPu24KTcFeBPVfLXxPd8FdJZ0eZA+Vb0T8I
gK8dumXGqaxKsW0hXm1vXu1j/h9OWTwHWt4GpoqxODWAWgxOTUC3mTaUXKlmZZmz
QqJWm3n4DwxtzX3TjHkGQy8/xinn72rljxqd3/VmLbdlQEGVMSlUKSIgnLLxgxo6
h8t4OX6TgJybVL/MGQTEBy3XldIQiKv7EFDEBVPRCw5u20opsu4mE66FQNfXVM64
M/B7nbruJOvCIkxtRgsMFIwnhXvsufaQwU63F8ikiP0HzdFl/aV2eLHxma13qW61
I6jCx+hCnEPBE+NZH0ormGjcsPHrDx2ZjPaDQ5lf/FzWtiI01DTm8NT/UMxLWdXr
Q9KA750/wpUkjxvIWRYBgL/aENG6rm7ekAqt5IjZp6RWtUZcKX/9423D9YDRlDW2
FjGh2NMpQhlbgEyx5TaZYdsvF+6GemkVrrSxxieRV9ZsKN10zWQtxGub3WC2mU28
2wWgR8ig7toubkm3bOUoU2JTETZ4d8Yx/dCZ6C2HbfYBWUydyBx06zMrFWgZGjTJ
yIy4NrXZKNszuO/UabVVZ2S7Ri6c2gEPnIKFaF/kmHdxojuMGwoaXZ/5xWd8OeDk
uhlPdZVoe9s8IhGM20nDUBl3pugZsenLiaIDTy0S5FPcBI/LLcrD1TAX0i1gw/iA
eHGUGSI93HWRc17TRT5WhwXxmsvFuVqd8+djm7M7g0AJYiiY9a58UJWsvAPNepAS
CL0J8iUpuTcj2H480RMc5lnrgzZ2PffQuJJqZHL8+RfpuKPq4vJOmo3z57UfWzov
+FP09cLSsPJIheC2Gwz7SAG6hqqEkeIMgARiw7bQb8d99njGw02Goe0LWm+wTBZC
QxNiOut6sbb+8DpKSBA8TNyqc5o3wWqol9Ct9zz+6R3CSG/u+Z4rebMfiWj0TIue
/FSHb4AFEmmH3pfYu7u1yeTUKl7BNlOpTO8wNa1uRr6MP/gHfM0jExUfnRKQGhwm
sO/J/3Jn8D2d3qmN2XcIiQcYXK6D8hRNQeypAKA2Mbju0fHs+kQdhwJF9X4b9haa
Xz1EOXyxio4jZLufAlv1pQN9tl7wE+x3Mv7wtXLWA+rsB0kkgJJwb/whjVE/YhFk
hVNBMRcnkPCFYsQvvVVN0spy0VoThTkjfyS1vhlqyBf4E1xZ1gosomPz5ltJH6tK
pGWeJ3UGyXvVzycUxrcRUT5R9+E768b8dQdIXvLoCxZxKeNYMPHVQdSmfMKliGNA
ROb3lqAnb/MrvRvjInlDlIO+er93yP+tY9Pk/VUHW+0hzIFzkMpjkGYnGgTA7mif
QnK/m3n1NR+8Xj22zoSz7JxiylBXrHkxxPIlOYG0gsh+SKGe/hEHhfWJaxbWdp1h
pPTFuW1WaFMn1qYo76Mro0W0MgyyoBa0/MKUy9NeLf3gTlnaZAqfa9H7vNW1+A49
1w+RgEyJS0ohW6yyKjuk6pOf6tCHEMWJoVKuFhfSTGWjX7noJXGMOGUmRaUSBfGp
GjyU/Eo1xJU5u4Y1VJdzjGRkbQiLay7CWytBIesJ8SRFw/Jmc/89YrEGrvXjcjgO
LoFWBkDthg1dYJIKqDORBpzv79lo7E03AV1TGbjSeMAI0bvv7Hswc5eHPA7XjAbD
sXp6wcN0NYFqkoQLCdNf6TLXpUEKY+eBSihJWzSEjwwaKWmC7MK/YnhovNSc59Tx
RiPCTLuHQ3aMVUD8y9khx5leqtiwvhSdl3zkSQ4RTvmAnaMXk3JiDkkIWA25Blr1
doj9uGfI5Sp70k4+vwgH78WUBCx9J6pBau3MQ2ShBF+hBHUhb4adPe5NHgeweft7
yUz0d3pxuGYvqIACT8HpSYwgJeUZmvf0mMIInBVCYFFUuvL3gly3MuBP9oHNA9mt
7PBXItxB3I0aqEsyuxrlmgwCU3pzr/axEhGrvSTjycU71s43NwxAuTsADxt/fybz
FjTMa/3hFUx4DmaYnzP14S8s6ifLHUY6a17bBW2up2kg81+G7IA06XQASuEO1Saz
WIoAp2/en6oyolKBogx+qTUjxxKEGUabZptKUPaaMR7LzGA+oOfSvFNmIF6Fmfl+
WGUezMLXYgZ4izi0tazK81x21JXYr1sfTxX4/ZYtk2ou9i4IRQCgPLEJTx33S/Dh
XFTnkZJ0gov0DJib46L4EKFUjpZ4KbZdoFxu60TVnhjpbhcXj8N+4hHvd0Dbyo6z
jftL+6qghNrjS1fGTG0McoP67v//6DjedCOxfJvqf5RgwwpZ0m6iulncR7iHlEM3
0RhzacZpHc3h1yy/qV036866LspmUsNRamei/v6R+xg3Yfqpm7oN9uCwtRmjJpFW
KUox1gM09rLjkYwYgMbXJHr/GshtHpe+F2hnvK5bUUrXSzROTIoZMD7k57wmgjeZ
6a8ZlFfB1Al5qpZLmNQ9x4FS6WzjOx5zZcSVwo0QfBVQQzBgLjXJPVtoSbJEAARN
JohzC2SOa2ZM7eoa0U06TgwhFjvzME5gpHiEpeQx7qK1xo7x93obEZez+lPbW/SW
zjeMgM9vFqUpSWYAjARs2s5E/DCI3JISuDSQ8NyWnYiRFWqRnBx1yP16la0XOrex
JLtxVloX3J5m818Oo8ra7cW55BaNhKYJlOyE6tC94RXE6B2ePa5+ONIXDkGlCE2F
jthrDHCPvIotX3iWRrNiTZASgGP8ZVsg7LI4TvM2RLOQ2YUHv6LRXRscp1aTlsfs
TnjuqaD36J7IAd71SUaFHeMIOddf2TKlW8mi1wxR4Scg40p+zar91TKwlxNSARYX
ncnZvk8Rtn9RY4B51J3aRe0OIKGp0B3peezc8D8SfpWYjuTI1mJXGnqEudSmEhBt
DmttjD6Efgu0xhn6IOwTELj4skzs/Zy8nBaBE8TdInYG40/6a/ZGJlO1vGY7YZNN
0BPMpo77iBTaOsaT7s2pcsIJ8ByqQKdMbgSExjWb1Jvy3u7f0gI31QQqmigy4Y6r
UyZlpO9iXnk/Ivnhegrr5si2K8hxRuVfWSZQlA/Uiq4JzUtWOOHgD7IOI6OBjDQy
8G0T2HdWSoO2doQ6HGgMy6u+u928pOoUpjPH2i6zxRzZTQJ0vqeEliTaa+N0QyIZ
5NCrZS6I0aixvshFSXTC/BzSq2QmH5xXSp5hD8pwI2tSzyqvsOMz9GxOrN13+LQj
jnIeqnDYjPpYj/BSbtuFzPhP1eOPTG3GYT0q5RLkFafsqmjyRKWX18mlio94MsgA
WqO38ZhUAJrooRsGkNSndDJOiWm5nkVCB5qlK417MsXLvYodVnd8tUDa6kAwBzvX
R7OZUBnEqKOPuud+852fU6DxjOln1Wq1gzBpCFNR6sVcszA6Jyg5Egz04A6JE1k2
+b4Me5y92++j8Acj7qnkx2DFF/3RaRtQmlw8GrWNkfp6oC/hulJQurH+ZRVwcn9P
iMSgO5blLkilcMHSHtCTmWXmSZLuUVbQ6lfD6MoiRIMnxUER3i2JxKIAoq7CATaY
WCDi/6OuU2WJiqKbNCbLMdrAB/9jZTl1Dyn/+zDgjidTmFigC8gr5nJgVUX2rbCz
jpbPFTFc5gp3OR1/aayQfuQ8+Ycn7ZS8AdcjcLcp7IXa4ap0sROUr0NHnq2kVnTn
i1bEh/exV2Lg1cZ27zaTWSnoJl2Mth8hEOrrOe1enWjCIA/S25X5zZfjTVPExe0q
QBYAbfI9CCCicZvMtccY3E9+WRRnRWEFBOlaK3GUTv8jN5bspSJRRK+Bkc4oFMJw
1Ibr5f1YXMZeE207t3ZQaDJRjmghdMuGXDVwdYPTt2iDzonqpQtmUUeI0Al0OukA
K0OPvxCndlmS061RolnKH+YWp8j52Dv0jIFY2dyu8xT+YedDsANqu5K20WyIohks
5EOHjZyq2RR04L/TSTfd/bnHbsu9PHoNhHk7TXidqeojihbUm8InZ4xWl8b0jIJp
fYh27XpBdU30MizOArPgNzVHthDt+RLNI2NfZMh1mk049kx387S4j+SMXX18CM7Q
e6UbTD9LmHwbi5KFeVWeqJm0H6Ow0hnmDyRWVnV8SwmSvv8/VodMRMdV7yEblRVf
a/UNLwVN9hzTlYroTpqhIr4nct02to/VvPUTg4tA/M34rRCGLUYXF0IUagRtT8i3
CMkHtBEIOFwFZZ3AFymrwmzqcSnlrczONTh7IvhHX3vMQnqjkeTTbd+/BDTfBV1S
cgbgghF+0iZaVr1lPLQfViY2JmqZavBTYl1M3SGEdZ4ke8s3pmA6qgkqpy+yrfSN
opEkBV8hXK9VSZQx45bc2tJUNSbCyaUKAeHBCAPzZpLgJcgrFty6koJiifVIr0HM
dTOZs4UJw6utMyC+IddPSd1efflKjj62V3o3t0tD1kWuDsbRFzDxQgLARqjuvcrA
lZ4OP6Dx5MDXCAhQVLdK/o1HXo1Cz8ftqYrRkd9fTNplattOkbl0wUOXv1Eq0XBa
Y3msxcfLhL7Bcy9tOWTe0JoauoQxInEi5ySAR1LwpGSjkL4pj3B/qjHYDxL6GDPS
SdH34c6T1A9ZfwZK5AVQXxeEER7nqZ9/Oo5afnYDJ1Wsgiw50BCOvJIcHt4P2k79
eQPCHbCeI1baOgnlpwjenaekA/sW/lN7Rw4uzUb4qHVn6n+iMqICPZn5X4mkU+F3
HR38PtVIglQw1sWnbFrh5VfFJnPMonAOknrKaXxZFBsUWMhRuo1fE7Zyvhrqyw5k
XJuuszMCYJzqdJ0JaeAy095wAkNk2Q9K4PRncOCuBRh1nSvRmbme0zhY7Y9tUn+2
4ny3EYoZmQ0kvhz1ZvI1DoxvCpj/lSiOyzFc0e8i0k7ihvVAWpc0i1azDEEIdOb7
dJdqGBcd2NhExNl6TrInuOzqjAqQccO1QQ22zmIb3kaonaaToPqTDqe+wyA0IZjt
SIRs9d8Siuq4nzvLPqq+5XKLilMwvq/eJGDWedqii+OMFMyRWTfGvZJP8FyuwYcP
vZ1T7WmmgWQdb8/oaCxvuvqGzpAfn4mNepchthPUGXGVdaS/mKAdJPK6CFaXVoGQ
3aB/3jrvPY0yW9DHyBSPUvXPTHkxGNQyFu3SHHx6Z1vCoTBLHLHQolBm8uqQeFpi
ou1q0rqe/jW9LbBdUIFCGY7sgBH1IR9Hmy/oobdqx2ypPgVsYpySpmhJNr4SN/Co
MTumR6cmlhjyIzGPvrlWkZepSxrvFeTgyQU0HlSKebtKsuvf/5Te1MUwLasbNTDK
PABsGSZ4wfrjyI2Pb4rWlITpK1pFQN1aM6kLbaUSi7leYeF7oyeruUTwPv8WzrMu
RIEapFKez9fVzSXKebA+qJeZBoUEB3bJ9n3KY2ESabQe+dEokq//TmP+iYlTdWBi
gXAD83jvM6IloTsEmlD0yieS3QFsaF5reDgtsH+o0hvB5TR+STOKYN4oKeLeG4a+

`pragma protect end_protected
