// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W499j9tHKh3qFEJ8Skzg7SJQ5dKBJoLaUoOJOD/5iyxMXTxwGqYPwH2hZSdD
KFBUE/SaCdHWOstPTXumjA9TnQNTqtyTzP0nXAlH7DQgHzi7TMy7yehgHft4
H66D5kK7caZ62jlzFfMmsTXJkvKa4npyOI6az1+PpOVYrnqE+fk0XLcLv749
sTCJcqxBPM4KsvhVbkXX3TtDthsaZ6j8UoKh9RC3PTk7dW9K/iel0/E8Pi4U
M2A5oVn5+qrVoemS2yR2i6Gf117758eTMmQzPer2e/MJJj9T2kG27tnCfzNh
Nn5EqvpU4wO/N+n7havdmhH0o+NfUX4Et6+bRoY9rA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DYkpRAsxeGJJx69jALUTDORMIxjMwdbPDUifFXRM4nerMaQMVARTBn6q7jCr
7GSdvlbuupoE+4x0AvuxgQiGeiOh/M6NP0PKGYmMPKpPTvof/tI3nJB9OnUn
yRLvwOH2Gx60d7gRJyG3wqYgN5iVbmXVyktSlx5dVgIMGoHkh0UzzQ+sYYbw
2q1+vulYEMWVuEflaxRForh7WU/8ZUItBIYYPoQrb7NaeyDDMCc7C5R1cKFy
5sRwscAg1LfATCaf7eiwY2WMYhXrf/Lao42bciI1w4ooJ1TBZ94Ywkwosf9l
SwXbagi7P8ip/8Dbg/6iz2UuogOJwNsbcrCUrD0PSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E4QvYV2rPWfeSjOeY1jIXDPnTS3uwvmWLlSHy5LGtS+Vfa6G5kpeGmVlnJM9
VtNI7SjJ5CL1ViBJTInC7bq7NI0a3pw4tlgOWFKHwthHTtBJ4WaLZYG6/GrE
dmp+C5l+PROdVGD3IUIjseDdg2tatpdAVN8+5+D4Lz+JuQFKYrEsXCp/vdkB
ytRQUImg+MOZ1SR2aDrt3ntkTZuEOzr1EuKfMgNisLwOtcBUHLIjNp/X9wL4
im6FyU9a0uLQbGd12VszlyOX7O/6E35Rya/bCpTS0Bsom6qBLU21G8rd8r+Y
fGTKujYjXfPHNbXgkZwQOSFvpa2fVa+wOky7DRkKRA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mcnwXFycV3bcR0W90blFZn8Sh6aA380+1ppCibEPLGWC0AWKA/4SkL1jTyu0
uLRANDYyWrzf3gBXJl+Jnx70oLIwUfjNcq4mKVloyt3wUJXGIKdKsFk83Q2b
0ZqpcloF4KygQYb1mX2pBwON2US+XL2hWzjxYT2gv16H10fx8jI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rBRuaiKSOy37VAObxbrsTvmNUTYyU5mzadk7RvRB4Hc6ly+95PYdKZ4YLUPJ
B1QWbiUy/u2n7wHhjnNNgnQP+4CXT+1KsYNlR7Zi1UWmhtaLwCAV2LBLxxv5
nFP8Ps2mNGVPSw7U49xNoWK4a72m4tP/JgH7yoEoOz8ZCyeQ+yzWKNfg5+01
BHw+OzxN0Cf7Fss3NTXhHpirU4I11Iofmz1FyJjZfMSl0pGbdDm6AgYJ9cyw
ei9LGdMhC16QCDl7KPMfNOntdsqeyH1GDAMI4oIbxZ+9SOi8FKJDhGx+9Zf7
XcfjWDp2y562PNNMz5HVnPhzhIlnfPaVDR0H2nv9bkjLYAW8WbRSdQFOc5TK
YhVGpPZOp9G3h3zKinKsU6ZC95SKtuOmvBD3QW/0TgzMzHBmVBcbBDBcpYgw
FYJDNvnYOVyokraPJfxCwHhMoGkUyMIyXYMTSdSSGoduF0sntZGBuwMhVzlU
eNCU5Y9FUC381BPwJ/EU5ry0QBh97jjT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZLTbN8ZL0dkPdQOVnY8iObuj4ivbzEEg5zBAOCUGcD2jQkQAAVZ8KxB8V4o7
dwBZGg/pAaFj3z81kBnbWSVN4AiUUk6hNRPzsQM1ZYIaS2QuB8PGoqabEiSq
FzGQqfRxNtr2zXcYN4EypLw+LIE9GGt0n/vh8td+3xG5zM0mUv8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Eb4MI2s9J0TVAY0QLjo7FVYUwmFqSdQChxhTkUIYDyr1GlD2OtYQ4E15DLAv
SST3m/eTix4/BNLcF6dLL4hFrtzwZgei95OzKRcRha8FVScLjr5xNWLosw18
MhrX7hUXh6JBohe3N3/QU9Temscymxx15yIHmzZ0A8544sWdCzI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 30800)
`pragma protect data_block
S4F4hNaMPtiWwehjb1ZQwPZ6cy8oDZQ6wKtUbQVR8d2+xgKjhFdIAtiGcs3q
oIilI9XTzkDx9u0bgBmzsHEYI3il7iaNunt2QAh23f2pGUSF5vZS2GAWs0V1
xMX3kY8nVEoil+HPNheVysBrICXip8zhSfXKYaBW5y4rstR+9rkzhWkwr8Y3
CPWReFmKZizJ0GyIRZbufo5Mgwj3cuC1bxPcOCpGwow4qHWh7j1xUKrK9R4a
nVQ73sDCUqCHLtE6OuFja0VAOcVuZ0dbggeBwKYf3MKF0AYFTHsF8qmRHtlB
gWUSmDLwLzH8qKwyXcgNOoWStscNmUVhow4IxKKuFXU4vftGWEO8QIDYNWJk
vwNYCf/g7J+9cCHgatIcLC6XZ53N3xWKWKPh4uVJOnhtq+Nhu2O/bXNrqJdt
NPNtA4JwSjO/Ch27bRTIHKkzmv+Fcz9S4ExojAgeAuv8aX/p9orVculRUhF4
BZynHmRroSCrkr2eggT3PCWoHWS8uDuBtzjdavkaYOp5QyE42OwWFBgpKOjU
JG5Z4O7uRiH8dBOLquDwcRmsIZ3vtWoF24t3LrkbN/bZxDe5vkfbHGADFj12
S7TwYCSBK+YOq6Es/LmMgJAKbJBKRicIi6pTJJsmlkjO4+IHxxXAwGRYk1ma
neX9gvI8AlOg5lovAzgdPBpioDvai1Q67STOozvnAWvw68/3+Xsa7Y9kUqZn
bQ7Z5ycQ0x08gsY3pPFE8OB2lT3LCOLl19MgUY5OkEzb+m3xVe/nFWjlBtiZ
RWawhroQUmAeDMcVUmqDpk9soEj7LIuN4WBRpisfbQwtMhSdEWHPZfuu2dSC
sCW3KJ8njnQ9JdPl4uVasr3GWO5DGtYB5umK9s0fEkoA73xL3V2EfCeD+Muy
m+QFk9eH8TgGEmcuk8Kv96P8om6NVy2j0YRcPhYLPHDpMShKHQZbPVBYm0S1
JSsyxkIempqH+6au+2c3UkhgnhmjX7f2eoll5p+xfdIf8RETSnofqs3zy0x0
Za9jCN+7DO8FwZhxdWn/r1MWS67Li7eODz5UaFs3HQudd8Qu0c/SU5INfGtB
2FO4ArG8ml7aWVULAXdA7wvmLBIBn33glZUz9HmC94zpLu1Kda7u57fSd5Nt
/LxGFrhwq0pn8bn4+KX23TNGhuokmuXNjVnE6MsHTtnKVXe6aJ/JfpyOzG4u
zrZjvSOGJO8N+7ku/cBD0Vo62HTVUrwTp93yQ43GGKHGAUkb64H1b9+5TSen
ruNnl7eW+zd2JGRoyNQQ1ZXD6nC6uEVX/TUoqNbF9OxJWFj73OR1SGT5e/Bh
2rHTJvot1OztgM6i+A4dhVsGyLEl3cq6fde3+RhI7Rw66jF4AuNXrVmxrmRF
CTB3g1JwQBcQqBrvO6GWLs/YwauQO3Gd8kKeEQrqLt+Q/ZtkS6ljnEFGEA/e
1PypbQq/BfReeAxSXIr3TFmGDvNrcAfV/JqyL//Aflzm/9u8C9Uq/5Mqxgxy
y1Y4B1QG6MIHBhZwCeMFBTItJXhGn507SSdRNbhb8wA1IE0I0OCW6JuRIbeb
0M3+pn0yb55O2DPdgi59ulFNzOI87BH7JbhXJn4uBoY2vLA9Unkb6HkwKeRs
cYb0UCJsyVJcWry/kydPfohJOHGXWJ+lpmxNhwq0M/B8rV7OsPXgohudsqMn
BQQte7rmdr0i3nSNzKqlNNQFwoU9onFKwtH7eE+eq5YAWGbG3pQJ+E5GM1fz
rUd8KU/OwGVdMHrvPMak1t/LJaopNimTbcgNvc7Sa0L7GxLoMLa4SDQjcb1o
2zfflSePwJ4o3KGMXv4GlJ5x2vpTWxQQSMRu6EUmam+kvTDDGscOdZ4QkhSh
9QQ3IkTWQ6B3v0epvm/qa4j1Z9OFWRhI8CbWqwYKkFJx6Tdem3K5hE4ao2tm
G7A8PchH/p8eU6qZA8kke7r9ixNV3YvAscEUUfQgsKwxDDgm7+qsLhg87tlv
8tVdfQ2C7DgTwgV1SyTRddWfH73IeVKzKQ4MG4c9arhJoWfLBK7Woec5oueL
GTOVJADic5ScMTzbGrhojuraznH+Pb43uWF8gNSPE28mJ99U6WtgLgeHdN4/
ZZ+Kj1G/0fdgXPhxrg7wH7sSPo1jVU+cktwmxodep4L9dfrfSDbt9kvLYTYN
WhQ0EaLYc0b3t2dntXm8XU4c8+2dxcIdGGNn/nf96UrW4t3cXlaf5OlmXNjK
ILxR7KhaeFGWnRqnVrA5YrcMRxri2pzGFn/r0Z8CAh28Rsqqwum0EwCZJGQi
onQNcspJXOIn9pyhSNzRL4uQg9fq7uRC1hhIeeAXh0v/AXUEEsYEqfQdA/29
4a2ghoUBZ5BJJ+Zzoh23SCga3UwwE4eb4p9uagkP4t78l24Z1vmowIHbchI4
c8mo9na2hxt8wNEYkYsXIFdYYBOfzKVOBB6ICEIylNkG6m1Uy4EXC3cGL91A
zhLJ4fW9R//3h7v1SCJPFPKmMI2rOVpRLQ6EgH3Xzpjkbt2JhjbPeLO8aY+2
buROx7PJ7yf8a/7TKtVJXmWL1jwRrzqz4CVRvCSNMp1xcu8PfpU5bcfGLocO
3sMmlIs6YomG3JjyN9h3kgaTZMeraPiJ5NZSi0E22N7FfCwNqOPaVLEcrpF8
AEbkixso2XwJTGVB87MGPv3muzxetqA094bg4C11M3ndiH6IqHvCgK39bSxW
QlhSSMnpdeKLwyNn+okQaOJIE77PQrFWK1e1l4LTLRdl6krafWewvqD2EJfT
94B1UoCKyEVHp2UtGKJ7wUJW6HBkr0vqVU5de/bnkPuA35M6CKSGDJZ8MUka
qHcGmEGmicOkDd9otS1+xKRFmU+me9IZleAVaNO7ynJR5ZZ4JIZ5hp004edj
lSI5uHAhx1bRHqFdiVzL5nk/DGmOvg4F57E0Zn0htGjqaI1W1DjRddHlpyxB
wMd4bpjC9YfcKLvn3AIx71NShjIxWJgQu/QpnDk6PPk4m+GWrjYXmcMZbIK+
yp0q0LRAfE+gPLrzrkcm7wEEnjfJHMWro1oCktTPMn3tx59kEZcwkqg/BetB
sbF/XnRPzDE9aHDyWrPVaNKOcj6jVMpBxvIDR33rCMuGCk4qeoCgWk6wAxTc
BFjy2oDC5sqvvDJauMCY50HTyM/rXWwy9TAtgYDpIDoVcevhT/LOgz8+u50S
sIvGdLr1ZXVpwYKQ2lrmkilKbRRbpHJO3dCGrEYRRzGBJc9/6FdnamzLuIgX
fo10bYBKsBfRC71tdKvnCvqGXPtOa4j7cVerhSIaW4MZkgqMSXtPqJHGiE0I
4YHCN8IoUJg8ywV4olmJT4DF4a/wPQ4YN7b5mPZmh7amlX3kif/y4KtC66EE
xZKP4QgBKClVMHRI7ZIUChzmiukKJk1BqEEYcHHIzRhN6aHfmWUhCnipvjS0
+kkBpvmhVcSxHzbCX+tIX8ztqOhSXPU7niM4BUCvFJr53VDDa+HVC31O36jr
wvGur/TBqj7AmBxeltLHg2ByK45/Dy4rmWR6GVXoYzXPRpxTFbj+vKSX/oNv
GWKDT1VSQEvkA4Vwrq3GWt8pbxRCiYqYyY+WTY3yq+PYPhfjUBELkJLfIkhr
9hCb3EypZ9fq28JDo1dUTLkVg2/ojU5bRmvnX4MRrnH7jqVGGwEIXpV6Z9Bd
jy5WaLp/GFBw6Yc5or7svYpQTFlyl/NQzPWivGsapYKPEftthrxMf706zrex
hEGwIL0jV4RlqMskjGDWp1PXEbgO4Sd4dzFTVbXffbJUj1fnTY3S4PUX/NoM
fFDDmwN4FhoPowQXolwotSPYpk2MAXr7U5Y087wii75yAXOzYhyjcyqSNCc9
0qncYFFUOYxYG9vGOsfHdZz/+R0qkmO9MeeNmFoCe6HHqk23/2eKoczUIyF4
9Jw0O5FjuR/jv9Wzwm8CLZEt4gU+8cnKO014fzHSByvbuJxnnW/PipvR3vIT
vy4fbx9yTFCv5/W16+o9bs3uILVjlQzuXOjdqgU/4E+RUdqJy6DSYPo59h6l
LuceJt3Noqf52UK4DSnfC/vpx/PHNz+OQXnjRnY0pjDR56j+h5gua99oQc8F
1q7mSd1tYEa6h4ulS9AnsGYNPiIoqic2NWT4DJNFJqhXzkLFCq34tU/OUQko
Ty+K01nLSLSjmASMQsAiDo27OZigVO0/AaCqRVXc2Z/3WPzfXkE4sImGA8Sg
1uWfhW0mhgWU4F4HTQE+ITkfQssNgvORLuoBqAsGgU++fKWK/tE1ubV9h3Kb
2mlW+pJ32jSGm+MPSfGGt1GhYob3AZZ0zB6pfabgkp8Nd4Gt+O80bFZEY4aS
jZtq1S4AUc7Gc4ukbMRyD3Dm1Ql0Ur66My/9NNUqCeZ2CLyhwoDelRmBxobQ
nDUl2q/4Y3ruxOB85Mfa6l1Xg1mQYbUbhZDPPFvM9W/929uiQ4y64Opq7VVu
NnanFDOw9ZUhrPTRs6PVs6puvvy2+UoMtJgr6fLIEjiwxbN/XoWC4MkpUrxH
846u6L2pih86yScJSQQD3VRUuoB3bhOhzHxPbp/tAUdMtRQN/slNwY7NGsQq
IPur02hAg/jqqPaWfInA3rnHPeke/bQWXc/WQbyc4HBXe8DZH1MvMGH8UOms
yGDd7/Gq+ttDfwYCx2A7/TAHzehE3k8KDd+csa1VRc4KaRwtF3QWYlmCFkVp
jPx2Nh09lwOF/AuPwrjSd88EklKLl05N5SDqLhBkaJVGS2TjzKWahhHYtk10
9oT/H454GtY77Iak51ATFIwD8oCNoGJ6aV3txcLfx+Otd86gP2tP52qFXp97
iMmv3CIbArlABeNSBknsi3iOWS+QmOBIn6ZK7YjfanFHNKelYcySvGcTdXP8
46VBGROurAqjgntIzKUCxaywZs4YQhFP8czpdIEnCOOgMLngugVfI4zSzdyC
aF0zmeMNIxJiwFQb4TmQKwqV6AMfYDuuwzVw7EuPAVo00UzdUpQvhEC7mwYW
w2ChcYdz0+3bQO2iIPGBWYoJBkZ/i4FGrqrXgBXfYI0hG4I37aaLphnpZILF
AKP5nNvIdQMjk1QL1QO6/1P2/THbuCLLqCLhVwYYJf3VH4Ej/v4QwDeOJbwv
joYeTsA0PbNTgerF+m5XXtKuV1dR/VEk7zoCMD+w/LyFKD92JjmKnSDFuzHu
UKW4wEGgFidLQZiD/jGDEaPqycgpnz18O5Ada4Yj1EiixWoITC+VVjOMUBkt
ircEVCZJAP39yaPWhfIDFeD2YUsWmdVUzM8khdHi4xxxVnICJu0ZyblvG+nn
m47Gemscdr1vCnzh48mhQ2Vx6urQMYpxXnuC8HlshVmVr3GOC1UPkmW7rCms
guyXH5jcGs/Oh2CjzK1ywwqvl2bEac451W4ZwDT1xfJqwRcR3DpzJnyybjzl
UgBBtb/+agbCXCijKRr+hfr8bI1QLC/7jeCgljnaTA2gd+K6gnLT20p18iXd
lAd1QUS7Sg5X2ibwPkB5Mr9PedDDp52WQkt43cqAlbDjHkLiUYUOkJx37aKk
pj0EpnfVx1cpb2BgxAPQj4ORgRWdJ50m7cLaQc7vk4e3D7NB8ZYb4SbsysRh
vfKS0rppa6cLfOw/laHMSmBLOjaQ+f2BF8rtKHqONZEUFw+IYw73ztEdj+0J
0u+sU++OM+Zg8H2ZiCfiRQPtbfG5U1qK+4YtrCor25b3vsOPQ+wlVqHI1ryi
fISjHGa/Eq8VfZouCvzwNBbynZ1wnK8bETHIW/aelf1LvfQP0LKOMP/U+ne3
UrdW69V5LMkQLGCsBzpiGvEaH7h+v5gAv39y1kvOfsbhN8OsPZOoycP3Sp0C
kFi33u+8y5IWpG5xwAN4C8i211BQyHivRywXlSxqNbeE4my7FfZ8QNNXOo70
lPThVtvorsw7hxIAvUt9EAZMhH9Usjd5yk7yXx9TMw3Pqeb9MKG9lzh3VGSQ
mN9U9pDWwefL1iFxVUaKPbKAnqzkQ8DLc/Xf33GVdNWXwuCtHQ5PBONbFXgo
N4kSkqRHG3fbthoFw/EPdMOO7wmUgJzqLRcIVMHOzhuAPVBtsZZjqyi7X+tQ
6DakxLXCC+KvDvA8aAdqUjgXgxiXdd4F59MkM/xRGeAjcvkdVr6r5zTXrNFy
+EnkEpRXKoKBwjudUldJ7IazAOiOCUypGkySR+ME9ogQ40wlP8XXmPSw43k7
vOY1vaXFx2co9ZyqPtPtDQS1EFCrmzCiZpSafzDwvO6mgXV0Cv/jhd7vKx12
pds1+A/wqI7yQNahaKXK0sM8qcYFxz8yW/km9jDyv44QRtEHfEZUprAKUq2j
mgkOAqOW5VhO138DhCoVflBvg/jNGYLweM3ey0LDB9d4MSHUnHQsxuXNNpwj
z6+7j4K9++UmnA5YLz/oErpkzTlEsCW+7Ivkrx2hrM4uEFaf0btNjh/vaCdW
9J2+8UIkBJA4KKBUIDuftHJ+ZzAPR0xJGuFYNFMlpl7zqniz5jr1JPRumRU5
RaYohJ/Y2QJ1KPwFEU3Wg4k64ZWLlPUS4miuEISysuVTP/iIZinon4XF9zi2
YfjZ6rw7nWOZW8MHzuVMKw9yjVeE1FUY4Kk+wl80oKoS2HTix/UXeE6OsJI5
vG+Fx3hsNqi1sk6sICIyvk40UWwNQ4XTp2eH1CsdXRBNg5cciC09LZai2HJy
sedXwCrc+GPwOH8WqxAfnDxcqxZ/0xv9q1+jp9ihcOgprGzMuB8jbBinZ3SD
shYvIL8vGvG6pwSE2b4e7mHv3hNmbulml9Xmmp627eyzzoyiF/9ywM2U3sV2
pYXUwQYDPpilWR1It5ZmBfk9XG+6+NZ6rax6vpKOEbY1ETawDzXIVwp3KALI
ivLZl5sFrhn5mauga7ZxxfiDlCjvrJF1bbiOKsD7MXva7xuU5KLS09+fRsUc
UlHI0tZVoT6pxpxcGtPXUSDXlnVw39bdvEUzcJ4z42iyW61zvqG/CpJcLhtS
Dvp8rwuhr/EHWcVRViewNIgfck3lZwUHGUX4N1wWTtMfdhgp3u6RAcVMA+Fg
2UwuK+rCOWIDSTILflijlbjdy4/2A2YT6LAxByg1uCSknsJ4FcFya/xi6f0Q
gwSqd4qLe84sQpnQ3jfYdDD8jlvX26x7p796t7z7qb5ztNS4BF47tbRatUES
qhrkp2+wOtFxTs0D4R3D+Z5+5lPyHhRu6ZyWLtsZEEH0wrU3ru//zzCafalp
34LNoqRYQflquZZFBELgCnpcqpCAENNsd48vsJu49mgwSfPxsYjsOpedNwG4
aw37FAvsVEwkbpidNoP3NoKlco+g1WUmCcMM0Q0RsDMZv2D2XIIR0nhQrsW9
dOKuqcYid5C9JbmZNWfoBkaDQMQuA4nicXZ2T9cvZlQrWJmodUt9WQhAmn1W
97R9WdmJgwxFVURuZJ8uGNZvNzEtsrWqtoCSAzso+WTsubgqCx6yud1dzQbR
Exz4PoNTFHBgGvt8KufKieiPc53SuFnBLZdu8dGpellQy/MyWynBt7Wt841w
K9q42oioC/j7HOnNp7P8qKWbsnkiknK9wVRnn4wjVuaN7oORSjrr34qyi+Lk
q7vFrkuxUWrgdzmLZffHLQcXTg4zJd6XZlEwrjuk2Z4eVy1oQvAiIVdMfM+a
ePw2n4B/q0dcYhTp5cC9/hS1I89PzxU5WxxDdTh0Dfskc1pS4IddaIT395BW
4hyGsbw+NXz/wQDy8p7H0lUXdyQdJQvznCdJ4yauKuJd60cazDG2bszxAbIx
xLZFr+VZIWkWGmKe5Y6uoJvV0H5ytUsfq543qAUUQ+gRTGGodc15VxWUop7D
TLZdMPWMGuA8n1XeV1t/myo3AlQ1Z6CTBM6jroWRTsC42l6sRIgv2IdU/qgh
3UzPP9MxWpTsp+vCK0/fez+47cx/86aNGYNSo0LfpAFfPlSetTz5CcHMy5hO
oMsGIwHa87Jh54JX3LPlF/oatIieRa3nVjPo2Cs2mJVL5ZvEw6epKx25TT/+
RXwHATVwY5P30+r8pPvHJZY/I5GKMVfdn6k8cFfiV60zVzmFXH5csXB02qJ8
BWXt/B1r2/UQVMRo6cduLAo/b+FjfkoYbQtmv4I/KOhyF/iYpe560A6WC/1P
NQ+GnBulJjymbxftPO5YcztLKucfUYX6GG70eOFUrvULYxRO7CLZ6i7JH88P
UuMY6biykvgBibPoxbC2CkrxZyozbXeUEXHq6y3VOIdlLsV6lYvzeNhLVaez
nYQ6fBOEzkftfkSuUJAnLfLh7RZTMD6xKLXVuHU6lqEFfXQU9jkPTtpN85VG
UO7dpQZjZNBeM7xru7/xF0H2VCaIyKnLAsLg5fLM1RZH64HDIBzN/4uSlJcO
rzDOaO0bR0Tc/yDCTKN5TL+OBZXyToTrRAexWDTJJB8p0nT00nT299ZWXbbY
c3giptu0u4P9SMMCs2TVDjfmWaKvtC32tjgiGYaphM0ib+bMkSKe7JQxZHwd
HB0zhqH8jWpnbVdCw4EpcKcCyv6LrVDR7t7UX1JonduYMxGWrnsILCJb4Y+5
zfo5WS4wHllLUb4wgTYo14vHiZN/fYr8GpD+h0koXn8xIp3UIqw1X8R7Tnsb
he6LHcBEU9m3GT4L3R2+/kEFw12n74JkFByyQSlhP5LtP3jW1iFYOxRkEe+s
7V6a73S7JscynkvV2sLQwW2jIQhlM4jbUiHp/wtag635aAIyAGIrkKTEKFk5
Ne7RVTLqX/XaHAZ1k+R9HoFyOKrXzAyeGC1zddNTrQX0B4pD3sI9C2hB1Pup
UTLmWJvb5nyRv5RoGXgsoyUSR+PNivWFHfS+qXPFvT6GnImLD27UZB86XTlq
Jubv68R+BIwoe1xcXdLHcrpJX26rZAXLNtei6ZLS4I9ZglDCn6P/6yC14H1V
hN3bCtGRfGYzT5A6zkNmVtKvRZ3OpBB/PBya1AJMOMQyEggRqiwNsiBXRAsY
RoJ3TGD3UU0UV47WDifTS/cCFil6zKTMRGHlfqJ0RNLmw8xXguAZyrqrKjsC
8sNAE+ONdeqcf5d9VWMB249WjVMumY38C8aePPdQn4wRZRLBO6n8UbGV0G3j
dD6jiqXA9yuN+EbdsEAaCjEiqAhqulshUKWNhTNVr6feEyQx9q0w7r9Hwuoz
CbSJl5yDf1uj/yXzV1ZKO6/B7nHYVnjicuboqccaZcXW9YPnfwtjtn7SD6I1
Tf4glwIM4yFeaCqODddNpvs3i3Heq8/AYfphoWTa/6d9+kRt/AbgrDrSC+k3
hPdXOHDLxvue9KQpiMJ9B2hy82HAO8pLVC8YKKpAGbKHjy6/Sxx/pr2/QF4K
urhUGjJYbIZVybcu+5145ufxIa9O0RtAMXtLfZwxBQ4AfMUvWpL6eNGEi9LF
hFDISbEmoHG1joQZKGhRdFqigU7AKh/auhyNg65CVrU7hh1sujaImXbYRLCj
gqcjhPNpKD/4zZ4nt0POygvnCYHk0Z9+Gv7xdIk0tTjPWl/GkOQkVFZdAOoq
gBJUNSJ/sq5vJjRm9+hrfFjD7SSimrFE2CDD5ldYfz9ehrGC39PW1L0tOdvT
HhUTAO/6wL0m8gVbVLJ2v1VLDeqDIO9qDR9EAAfxFUAHYgqSNAPpkPNedM27
bhuOZJaoEjJfb6Uv8e4SyH0oGMKu+41DK0dCFzIpdR/yFSvB54Xau/ALWMSG
MUWD5ps225OHehYh7lTwsIRIQK3eg5zTyHvILSPrxbf5fmGZuymT30SmhZKg
F257b5ZSSm7VHxOy3BUkRZf1BqLD+xqbeFYX1PmwBIyrW9fK0pLsB4xnn+U5
KJQoxz13Nlfxi0PqGOH30/d/epHJCzscIa52xu5yjYcGJZbI253lj8wfMft9
vxwqq4cRyYoHnJbednDBY8P6fRi29Q7RKEY/58tafthKQ1rNr8ab3KEhRR5m
YluEbudHpq8H3PiOv/9gLarOJL7isM1g+jE9KkS5s7y4Duopndme11AlCIgp
2svQF+FfvwSICUcsI/NmwaFPFpcvUjVn3ysrGmuYUrtlQ4gnmrdiAdkO+BfF
7Urh3psK/oYH+p7C+St9Sgp87+woffcPx00ENSsBDkCI4U6jDNsBVL2e7I26
N2bav/zRScp2qfGR69pYNPfU6ztJBkZnbI8PplT6j/QIcU0vYCXq/HmJik/J
5RVFdtfli5ZFFRjJVW4/2EnMBUddKLZ11m+2Ci+XEesVmhd6Mk8F6t7wbOCX
LJiGUUe2Enm0K3Qp2UyFDBJfMuORfZMMLsL0y0I7mLPIJh0527OKVXLZtizj
Zsu6Hzj0j/LrZZKgOR98D4Ahp3aeaI+yfOZ9PrI0NK8Mls9Zz20g4JK0knuo
Ae5LAJI2d0htGOjuojNKwf6X9cjwUnZ2mX+Z1fJaZxgJz0TJ/ItQXFqtfiir
k4BqvczgfrbfOrrBs5olsJ20HzdH8fHFlnCnTbqpQ9G8zulTC08y8nt/sJOq
/vJsvraye1WQ/jZeLB26BZiEfDENb1uWSIpaUz3ykMTbznjSS2IGlVSmaZm1
bUKSQbwC84p9J07E2alWINxKKc/lPWQIfhcg2Y9i2NEtT/YL6CZeJaXnPfuC
SVMSPFQhxUN/EQQBope78tSE/vBkskoKM0NMMFMAqliwadPNB7c/3CumjbGx
edX1LLF6fXZNuXth0XaIr3hKmKTsEFLYBeYM8dJb9ZY89tGKJgPMLR3QjaQA
hoAODwzFOne0cB+vwNZ4vuTD3gXKanEagOIaT5172twHQ8YjJhB4ThmLOVxW
EuBm/OB7htGrhOfhP5LgYwJe27LsjOLdFSol7oosciMAKlhTh0LrOkoMO8Ws
GQ7XuZtmzLdDSSLbr/dlGV0Dl8hH2RpDWxwT0Gj1WoVcWvEVeVj/LRV4ln8n
kVIWmvuI4zgz1okf5JghZLGdjAY486cvU/tM6OTz4E4Ggs3QO4sx+CW7ArbZ
wU/rdzod+69DpORRkVlEYwtBw7o1TA+5kga4SKlLqfwbeH84r9AmXyRyPlhM
uVpCmOCH79bdeD3RXqPBggVo3AFhQaJL5iSDy2gM451P1d3o6aN73YvWKIq7
Dxk2UzzQq4xti4q3NwVEeXPUL3HmEBxeLXlDcrIBUDjjzGx7fh9RUGfXuCWs
8AWZylbqPpxTqNHvEwZlz6LG4fMt9y1JTPvAXRIoqqKWRP3J5kbuwTFO4ch1
xLTjT+lQPys59FAGe0Tju4oJLiVu+eeWr4TGUW+eMbRSpqbFkOCU9rd9mKio
4t80ZkaYS37sWb5JkGhPwLNiAoiRwT3MI841Pj7GcENissx7uiZJaq8F73Ap
rgPTgeoPrW1MT/Chf+bwTICPICKR3g6ItjmmWqmcSr411OgFCdyhE8FPb2zw
Q4YCsvGYpKdbRh20QYgDQusFDqnYPlAzeXNBScrgHZ/PLts/TR6WLTq6oeSD
rRrg51YyYm9gZesz0UnkPseB17EuUZkPXwedexAS9bec5GygbfvAvcHVkGvM
eig5LrN1UV5wcO6KjPJCfNAhVRAj8dEQ/B50+iQHxnNgfJ59S5J5ocEZS8Ra
MCVS5RwyrmJK2UaOx3lCNavmtKLyiku5hG2eUxCKIhm/MnqJN4vOoPK/tBid
jucb1CzwdcH0RD817tJpkQEm0vrXvkFS6Q9rwW5IpyeNeS0FNLIP1ttR97Nm
ked+iH6O4lgV4lkQET9ReKMkiOE1GAP5axMFtWcqFHwBZsmg5VeVUn+TQ+zG
2TWoBkQUO1x9Arqbh2wh+uYDY14nQxpyppdcjrriPcNSGhhbZtLDXuXnRMmC
CRGCn48lCH+1C5szjxx/0VlvQgMkzOYmXUKCUWF4BMm36SAc8WLd6sXeoKu7
0gpz7yNzOqCcR6V9ScBDZRH3+ADT9EWOFsdlmHwT+LCVTbukPomrHcqvvkE+
XbMJ8VqOSCvohkdPihhORB1CM48Dx5ebrWww69jX8Ksnn/eud/cY6BJx/K8U
bMXHFhW44yWICUn9/+1GqXToy3A78C4syq5xwW7CNvcUm9h7Cour/DXw3uhs
tSHjZrX1o/XDEejMqVeD4Er/kstUvRAUG69E3Mk+5xa7vmo7OyIeecXZ0/60
P9NpsUH2H7PQBLwbk2PfAFX2HbQNQl701PZPsZw/kMwCyav5999OcSWagjvq
+M/FVuhn2AfYHXusPi/OaXR7a2DmC/eFkJEA6HX51BUNgp+jlwXVqDtrVtpH
vCil80sPt0PRN4tEzvIq7B67e5kvgjjDeN5fPUQaVzSpCxTFKnNsSWk76lMM
dgUJXYJFmJpIjXsHyQUNr76fbXVSVxbobywHQyYhARPbokv+hvzMvDgFnSCL
23uMAyPnqGtO9MXrghM3ldjOj+2/9XcHxpat4hzQzpW5P014r+Io/wEV7LiT
5Hh0s1gTJIeqyXDIIDxvMNx6m18lzgi8FE+YLhtjLwsOVMYE/RZ8YqF/SJxn
NMIa4BChmRnnwUH03LIz4Iu18q+mteb5pLtNeuV1zGqsnBOO/Kupp8SIVkKM
F2cymvt2L6sR6QN4DF/ptU7FVK2NmFLXBcYog9+W4bqQuVG1c4tD29aa5344
bcZyMZXR2WsdcJoCrCMYS7bTk1a6O29WwiJdUvxW2ScAs267HDFyJRUslVmP
Wgwg/utqOYXMxM9el7+Sz+7yCgk0zPC1jx24qRQ8heuFsWVR+4kWjFUAiHHh
hJjU/3N9yHHILNcgyEwCEurirXlg1s82IvTgcmh+R7d8IOqTp99dgdyZgUoy
2QfUwzD21e4EqK+Vm0qPbScT5/bzQSC+cyy7XBFBpTtre/PB84zR1AQ4vqWU
LRZwvfuL2EGRHDvtRuHjweySAckkwlETbp5LqZyu9WvFBd7snbIB9Uf4Va+7
mABeKIvBdIknHMBSer0gDwh+9MLvuub8yupJarscDGyXpvm4T3SMK7qOV816
cCJRBQG1421UXLTLcz6g5F8zigEKiqUT6OxmVUMZ527Sb2Ez6nVInoieUrzr
H6Lf3oMoulSGoqnGh8+VmYoCpPqep53OOTOIRocfIESrBuxoxNC4Ip7WpEiN
BPF+Gq7cZy+RRj4hAtp2lBhLitpsUz7wKFrnGkIyKxvQUU5S8+FJ15ryON/X
ntApZ2kMuZBbJVCwQ3xmAVNttHOy6OmuCQuN1msYI2k3t2WP/wYRNlofRXcj
dwzP615LyGW5AuxmTHq1XbOVBkocri7oca+t67R+tesy1YxftcfHelPb+yQe
3IzseV3xyEF/v1H04DPPvkDays2Qa2EaqJDgI+Lr6fwE/oWocrcX8H+qFyZf
JBbVn/jlneXHgleXVqmAbkwQLC5D7FjeCealN23e4f/FYu0eVSP+28LDkZCv
8RKGJMo3HdGJQibyqXdBUYXhlj/m0w3myX4njmTkiBquoyn0qHtCuEaCjtyv
8zxlZOB1IcyPYGZFuoNgXV4EflS7iaBwRVV540RGv4X+cr9itPX+OSJJl9DC
v5pAbjkmvSaqQA86zUZFeMUMyDwsAD1PYG4RzXsGLJ0fg37tiAzcpm00ljzV
I3YOh4aT+uj+EY6+POnI1tqeuA06w/HpcRZsLqyUUM2e8p+29ys3Uce+f4z5
YD1En+dmJVNknnDnoZ1B+DEDLvPB+YNRgNORZyMQrTM/sOeFOunXy+KGC/+c
mBBa8NK2UrxCcGzjHGPkWFn9ue06UWPNqnDXFjJMKmzpv9FR5p+C7nlJMl9l
Vay3yvkxZOyaiIIa3g9/Ar3df+d6OUPiaJ7Ea+eSajcpK/Ko8ycq93onQTew
qDGisdPlH/OYabmiR6xwRrPgFdZV9XVfwpHLGkeMYBBYe9BETxuKVSWkhjod
AIJ2ETIDpfYY58cl6BB9vXoiS8z3o+JhkDd5cwAytnMcTwAxCaGRZU3SC2ti
WHyXRAdW26eIGmBwccSjKrl7wzOVHC7SWTDAErsm7/liOiXgd6tjxsAt2PuP
1zswbY2ONd2oXrZePfly6ST5TBlp/MsNzNuXKjKYRwULyXuSH7xsfBl6Wcev
9iPQxd+Z5Q2m6ThT/+SBQwekuPzBFKXyaQIhybmop2TCvF5d3RamDs5Pipgt
MBahUX0yOYJ3BpvLACvNlyiTBh6mEO0tfrGkuH1t3gDdY212fnl4edX/HGQ0
23EH9HYGeXAmL1r4UMQ16NJAuoIr4LRxRqi3jJNnRUJZexaKpWuw7E+VHHUp
4cXpjAOZHpHpPQNpaFoyzRYdzqBuBYOUP+bZ/egO3TBYA9ZE7ra03rNH6GA9
3/bDXbR+oSLKMMUjI0EdnJZ1s01lNHrezvREe2/PtRoVKSxSJVaSvW1+5Tg3
oiH8oKkblJuCB2xtH2x+pUYJ8F6u7buEAs28M4izgLST0HlYpQiUw0fHbT8o
TPqwV8fAdUDHD8jXyPMxmp1WaNyVNPRu5CSiwY8stVzc1LyiAYdHRFB1t1DN
90SYZ65bF7SazFFOt0x1wiFyPsrdHfJX4Ffzk5AZHN04uyGRENYUeHJ6MbBL
CvP/MgUdUShW0oq2M1mUx2ZOzWd8SwqNOlIqrG8vWmwf06F7U0NToWNH0RwF
A4vUS5QsfeJUcii+W3C+CK1nzmyLpwtO7QgAXyPUa2IS080+0VeITg+w1kuW
3iA7fisHvLJOeVcf/c7H3qeyRduUgFZiPD85Kh9g+jn+LO3JeZGKP2gtw7w6
x+Gk3t+rCGv4h3fpzgUfRXd0Yu4x+Vw9CmNTvC4u0pjHVv198k9u9Ge8pHzP
AFwn9y60sHPW6aZTr2UtB0SB1v4AmKD9pHGqcwQoCV054NsRlOysv8fjdqMP
fMtUVtxxrL+9slOPqP6s6uHn4i7YVUnISZG6XXmqMZCb+eLd1ypMviDEb4MM
Y4oU6D1qpgmc7z1UrRAPewjPLnCYQOm2LX8t0Cw0MahxZGpo4YUmoA4ooMpg
MDbaQF5H9vabgONivITmi/9b4PgEAK5O4fih1AtVaejqqquuT2KrpN8QzSJU
gGhI50cteYLe4+fLMHV2/LEaLDr7VISjlsYcrJM1lTBECIFXzioO494dILle
TdfhFpuA6xgLDSTQO1niNJsgb8gPEAjYMQdFsDe3c3j4NLdstuIRc6V53cyM
zyKl3Wa+RmRiISQoQyaf/Vck+N6pn4YAxRA9RcAqPgul41By2sNNimzyOAAc
GlLT4kEiFtkY3ziKay86LjPp2uuqyfezpSCJdhb0yhi22qTeajq9yFGMzs3Z
2w/CSnx7hlZAKi4KpHMrewAtcg6crbftDKqVD1+rTDpkxFL1kbBr0eAjPA2E
cTaQf0KBfxa52ijG/xoGWEv6TMtM0jlR52gNnopjPHtHVs085QtpHWmk8KKP
NRhTg2G9CIIHTbUHxfCFyMbMCuHEXoi9Lc3w+GHyJfPNYnr8OH6aZO6n57d0
t74VUgdY203E1hPY1pKQho1z+aRer5uDeZk/5dWrsqB849hGmfylnhH3m577
ADbmS1MDkKtN/flKGWiRlC7ieAGIL9+2ki8SThIqsruMQcYbHY62yDp4C/Mc
X+BJ/EaO8kIsMVUHek0H047rUoGszuXvsVbV8Y/iajSEew9tMp4IMYJRoOoy
XWuxtSeRpemaHc4A46ZbwErVsZURcJyf0bHpTs9d1LZog4s8bxPoof7KSvIQ
/OKAsheM8LYKOokoCSNjf3H4wJheIVR8tHkuAz4QNFIDxkxctDFvRqCOeu0x
z2UQbIXMEUTk+lpLIUuSZqtY4KPSL3oJWS2HnbFyhEm2AtaoigDosrEKMGd8
x/FVll/hhv4dsIv50Y6vddK5uuRkADzwiCZNa7v+hohd5UXrDSq8mGvA8wcF
0nCMmTVqJXMYuQWzBlO2UzO3nLTRGeSeQ8wKE7MwoYpLvkANeeExLqMoWZoO
bVZTxbvyKpLvgr+YgdTV6DtR0oMB8fJnVVLkdFRAjxTktGJQXfNJla/Jped8
8VmQFiWgu/WoehfXDi/wYgGUV9NHdyZB5VLm8yX9RCOJJCMda0qZUDa/Q1bR
MlllO6qyXBMw+2B92QoRIpiTlTcbRxxsRYMW7kH0n+U9ujkq5cQj+hHUaohJ
ukPZ5DSb5PpOIVfGR8TehhnK62/NV3rldRxXj1kfreppbt1iUClCTcAmGDo2
RutoPSUyLorGmJsflq9gyX708qxmzHodSctsqtwuNwgYDIcqFV7zxy2Od7mQ
E7CB+9uftGtMTEQIK0sqPY6TeOGb0gP2Jtj3lOzScnsSNMfhchgLlq4fRR82
Y2kVCPDhwiOzqMf6pCkNI7hTjlyXn+fU2m1e933GNKKaVzqKoCA/nz7X9eNI
digUFGFeeiflMstzgmYhIfvScGSR2Ul7TOAaj9fcaB/2CI6jiesLkfeIdPgZ
cDIC1JYUzMAA01xNtn8TYISWYFDtywRhUo+xDc/eUpjAXWc7IBNYhYPwcMLa
5rpO659gHnHFrqBVq2T6fGtmsDdXIbpCVl2N0D1pU0rgPjtcslq4nQN3rbRn
JY1EyI3WZji5Vf6s9RVnEO8SzsIBOlWg7TIaKxtanMjuKetukoUBB2j5DJE8
GwF3s6Nljwvj0/tT65Q7fsI7854WxmhjOCeDyLdUsJqAyhAS6LP7kT+juyQH
HGcTUnxf9qkrZH9aS5zAxT9X24gzz3zidB8BuX5sUZGgOfXUvCfJ353QU1fS
wqKU9SX2Dv8koYJVoPPt2Z2Qqs0UAjwyHmJWCtAA7C/jd/jRddKR5AU8tYmt
QZOyKLJfmPxMVXPsWz0IdHLO1wrSbcnoYK9Yor0703S0A6ywy74xWev19TT3
VbLdSyYNb1JJI3595Di/cl/gG1tRbE4jiSBM0T9ZEX2e6KzAjFuvzYvXlKju
CsfQqVtObqV/6np4JCHp1fDc9C9IOmRbFPw6FCXXAF5UfvS0Pyf95an++oLR
vAhrZBP7yBnn2eGNJtK5/jW1kUv2EzrV3QjLqwjBKCQ4Iy+iiBiqbjxk/YU1
uy+RJP4J3FOFIvoCUdARo4p8HLrxqWpbhVA7OcjQ7T6YLbKVN7qpNoGcKrQm
QmKtsBmTaxaH/aJ6Vn5WRikjlzATrj2JzyI8KictmyVXYOwuQYTDp8ieWiuV
lSTOtFJgEBTtbDKnJKcYK97hgAyC0kZajunZmhX2tUoHSyTjo+n8yFPJPmpx
fX6UjkiL2w1D7SCwbmNozjHA7dJjPw2+5u3tl0Ods09OaunjJqI5p0/GncVn
P0Y5ZyMKt1H4f+R+xcw35TLHjQDxncO+SaXnSaDcR9Ct8v4g0RmMZuRyhUfy
/fi+9UPokuIp9UFKvN/wzT2O6ifH0hrQRfeiyApyDU0tJcnZOxV+ygYpek17
todPpLEpckqa+zK/jLh7M7Ya3mnEeh86j8UXOFTMC/MTfJriSsbo8cRpsrl/
ahYmBV7b70HEUsqwrsNC9ZL1hov1oOIsFCbM9RocfeeX9/4Omaw2/QmTwnSq
FinkCFBDmbpTaRJlsNL/JlFP8jHoaysb1uV4a8kLpnTYUn65ydm69+MKzg2c
S+PMZKpzjrs2pPQ6d3TC9q8M15vCy+Opeyu/Q27GVGnfy6YUWRSQACeFgfDe
SaosZ7EOPQsidGrMH7dz2gpVx3bpCp4L1fBUJjpd/SE90faX05SIWjzsp/Rp
A5LZvaF/K0Z07zwqLIvR5nUbmAC8+ZF136y9tpARXAz0h37Cw1FxDLSaS7QB
6ZZF4+fBhVBu+3NhXbp7roua0EHBcFOWT29XtpDOJI2l0VtPqCoaDj+PScYq
i28h5wArJk4+BjXIC5QBKdlV11B8I6pvIQVrPt6758eoaOf7mRO3tbRD1HoY
1D/i61T/t9xHWuzDqWHAWp51zHfX3XgrsO9TyD1XXuiy6QAmC+37Kxqf6caq
oNJf+J8jyGu9YcGN7miajZrZjLMKx6QbWO17Fjybe7ENqpkCaDwg0cvkH9kt
RYD44lE51FNIIBld+e6vceP/iqX5i4ODq68bwxZv6BE2Xh1N92jSK4Ipu2EP
rRMrc/7YwvvCl9y8tmXftVEB9AapDiB1XE0CyCDHBRjYY721AIyvSMQkPxnf
Zt7GoDK3BDOT4tHgRAWsxSSz4X9f8VBUaWJQ8h8tGORfmrVWrasjZ70Iw06u
qLYB0YGsqLIOzhnl/zUrOFIBdgodmDxob/GxI9GnKy95kMoceIXq2bO6OfHu
mG2TUkucFtBFQD9CR2b4/dzht5Y1xZJnsQH/gNBDCfbvwmI1t3m+A/+0BiHB
hxyBcYlMM8c53RvHqhf3APpHfJwxsS4va+9n6sxRdaFFHRF9s6m23NU47Qgc
NwHUNlnnYbHQiTJuLA5aQ+ufly+1aQey9B0R1uYS9qxupwN+w3ojLbr2LUn9
h80w9kQ2rjk1vCTTYeeXDj6Qh8r/bdSDs3NH3P9+CB4HGrEhdDUgJMnAxjuD
Wbrnb3978731O2LmnfrghIgRz08ftjXOp4cbQ+6ZcT71ZH98dm22/7xcIa9j
5qGv3+Otfk41b6G4GtQcG3S3wdJVZGJoncsyIs0KNsaSdvdqhS7I2UpkRR7/
EfdihqJIcbmqYcZeSc9dfhhKwW48wNjqy8543WLAmiithoFUuHst9Xkw0Tm5
7oJ90QF7kUFZhq/KkrJXTAEIKlbvHy0bRJZLwk87NK266rxqmG4gjaOeryr1
1Hy9nZGCBLJCQXtboCEOf4rF5ghY6adyANwDIcjMUif0PqEyfMsi8vXRD0j+
uOsDYE64UJCY+q661EWt/gAOdhUG8yqEvmBI4nwyK13F1E/6ibv0vuxJhysn
atg5Yu60zze+pV4m2/2jdveRaWr6Ekdfjwgv+GN5OSw/nUNbaibR+pBmoyPP
ooTPkmCbn4dJeZMsOGzrd8ETcPZWYEqOzpO7uShvMgrDoemzC1zyySi8Bmm8
WIK40uDze9IHehxfASvvnMy5LBzib/23gPkTKvgFtV4Iy1ZoJXI7M/SSU3To
Q8QxBWSuQl2SVKitDX4yKxb3WgDFv9LvlV6VyBI4Z5BspLDflIzLSfoGMjJ5
V5z+4g9aRKFEdMJYf+u6QUH8wwuRMoRPCwtbtBDira7J/vGnwVGGCziuCgJq
wHYRFaTXKWcv/U9h/VOAn4z5Q+SWTEdJ2BtMW5gOICQm30eosbnpGjRJvzAq
2G+AS/+md/LY8fdeC8Y1pncPQ9cXAlvG4NfWHTEZP9cblDAp0wBYJKFN0xDL
KXxcu4O1cRE52EW1xAjAzL2JSboj2MKdSpVU2gU14fcswq4W7BUtP/kktluj
CBTIiZKT9pyY+QzpxXn84McSbB4UeRuM5ahkRd12FVfIEDHWokgxXF+1Id53
1GV4UtFgG9LieDajbbSJ6+frwbt6f4q7GbInZb/qD3F5ZEo1XNIcJR8q5Jyx
pMvWhAoWLotKMiBGb0K6aOsnSmXtGlYijbVMjCZ/t+lmZkfxzjkZ9XU+zBHs
LSSpV2AIXEPwSmM6yTDumhQcluWHIro4mCnP042VXnWOL5n8fNxRa2z59Ylv
GAl9UCwP4yVhNW62dxgnQ2B1l30ddLl68aD2Q+ZBF8I8Yi4cB9GQ7b/+CTAe
CRnxaycmqDNLbFHitEkpOtGno0MgbUth9+Nt1KbLWDMdNHi1jnOiOrO5o5TF
k6/ja070pFwlfqk3hcuYoOpv20ZDqHQExp8X+dAq6wCvUxl5peQBvHENWD+L
bNt6poRoG5ZrMBEzjiodJpA/byWTVkEGoUxpZ5oRaktTnUiWMVn9JpIIQ8OE
37JulnVk8rcRdvHOQ84Hsn1Eezi5JNzD/jAtVQjOb6eYjqwThSiF2sFsCXnn
o0z9bvo9UP/Ooh4xhVEjtfOhNqq1p5LEfpCwNj98+uD6FjQqWLpN9NaxL/Wo
IxSysBFF2UoXzYNZ25nu9Bxak7tp4mU0eJ88zkOFjZ0w2WQ/hUxK6BUX9HB1
8j+0M+T/vnsjW+GIdtcX7Gs9azEM8otjGIx2saKb82ONJsCTBpYRfI6ZKpO9
O/9hgMIM1EU9aY6fxbA95omkGCsV1yxtAi2Xdu6YVlW6u1LefMkH6c4MyCN2
rah3Mf14C+PYFQpHO3Tl5N7oNVUNcq7i6KeXSf5nT4Maw7X34iMSurqxiU7h
ci6BJWvZEbVeGzm8SD/df4vznzRWw0gbdZ149I3991H7Ye3o8W6kZsDEbIiv
CWxHXUGpqcFSkPbQgLIurySb/eXDolQc1M86g52vVrF/Fpk3uAj6YJFOe77z
E6aI3tJy1eKfewpO0tzPQf22BfD8dDDke8dsvedHegAHqf1RTFYju5Tb4Ao7
TZgLBtg+DslIjCFOHk4/DdjGbFmDo/h75v68tAimBVpBK0KOpUuGWm55JvSL
Gj+PWuQGmbxGzu2+aV4GfXXoEEMnvEy96VJet3RqqNqRcnHXQajv+at7l/ur
mSiMTQwgDLOrO3FlE/9fD5Un2/i6Rm+sky7xlNWRRUGvAGl3nNkwz+hlvFnb
MKnXjMoC5gW6VoHF3T9t2i7TZd8kgdcKh2m6qGEXk9e/2+DZIFOwQv6JGa1i
owgpeXKSPsfee1yI7u9kFU5cFelmJ9eeDpoMIvQfdRBCyMk1nvzfyKwrkUD9
HQnD4IQG7Y0P97FbTsTePWPhsJ53T1cjJroMzbwEoAusUbcpyH3vDhPg1x1u
RFa2PQeBDUyV/VrQKGNvaHI8W0z4BpkBPd0VzTo/qglInkTlfKDLSoOJ0T3S
oOavksYlleDwpqHPmdjULTe6q6nm9mBYMRs/kDGUlfy4OCq/wGOesx/TwUxR
Er/ja622PQV8WivJZiloFyHVs8AqLRMyU/CnNsdllc++y1hh9jtq0hdUhEfO
v7pO0ijXh8ZKqkUpZ7/zGjVowXL15NrcDO8MYxEQ3/6aErhmRap2hoJPx4HE
DJgToW0Y3+AGGeevYKFNijuatLc9vO6qIFswWbw1izVX0dgNJSpqi6Lq6CM9
QQl4utd6w/kmS3RMiuERdc7FjqdilYVQJYGVr68OnpZeqiComseTnT/6sbTR
MMPs6XWrCA1sRK7J7h/gFRa+yUixY7E35jXFSlHQFNYVUax6AuwXArttdhBg
NZ7DFhWlXjxw1GQrv3BZPIZryZn6yvr5qp55FaNQuq9Y9bRmJbEFATqs8+tS
6v11bjUMCyt/SpCi/4BrzlU07b93zs2MBUIUFo1u5p6jE9uQcBRPE2xr+9e/
l1jEWlMqonZ6L7SYsnR7kDuxtHP3HKPL7zytvjtkuUWzAMrIETUGErsP7Yiu
BqXb8IDqcdbOFaO/mP4ecM8RVJVjWgAl3NzDxuRYyWw/G4tiHZdCc+twNBsZ
QOfksa3bsx6gso04tmCisg0BDe9JcyUZm4v1M15t0vSzgxvh1WW7suMkx+hW
l5uIlJjXOWdvD02ga7UgmLVJfcMZ2sxLaerx658MXQi7i8AnWOW5sr3JtWUa
iz1b1XbXacdl42pobBc4qrvPLhDT6wXh7YeAWp7uiCLjiotywZfcN+FLeF9q
uJWXw3zWrrV60aYLTtYePvbGiFucgLOIK7NoCfde9gYzA78FVKt3Dv498Jgz
Yh9xEJiC6OfnHeoeepVjbpAY42Bcm9MzawoWx4Yuj0LHraNs95FrfhzdKb8Q
BtFrh8B/YEdj687jqwcFsi39aZ4TYjZ6hSw0DdRzTz2buDPWWwwkv6bq0lZ6
JjsATZeUwx4J2v0X6OO96sfiUayfb9W+6/qI+rhOgVSI6kquMzetCseji8Ha
RZIvPTZ8KYXDY0IzHfioXSh6BUvVR/qSWQFFTcyr7XTUHvwkxzX5z6Kuzp6c
ch3LZBtbe0xKoc0D2FugEREK/ZGTb4ALtl1PYB34zntvmXWMiuO7P/Qjewfd
+7SdW3xzEGP6gRH6PIpoz17NVQAXkdfwtjGjkdkw/dREbPq0Y9AFFlT7DChw
3MMRNWk6jU48n7rNADHpyCnGMIQqXx9j4E2Pk+QEee1Dljrs1Je0mAilLgmy
0B0Glyy6eisHgJrTowV5KYGcuDDTfK3BJscevTHfWde4t120DbIs8EFUd5Mx
cBeyYSUClsUlR99vfulU8N1fjgR2sPm6M/h+1leLJ4nWI7XiB6jLH+050KMB
oH7u1gWcpgYsGwizBbo7Vw+dXf6MZ9Vr7AbpLpmyYfxi8PH+6KINFqmnFN+L
aTfcYT2dgu8tNHIsf13AKUDrULPTfn+/DKUMhlqQrxzC2diAWZyu+fTCs3qQ
ayomOkRM9b17dqYX29sm4aHlSxKqB+Tn7vaLaSEfFaB/E5ZdzTlFAT1qOqNH
HnfhKm9AhIg/XlDk2FHChetZvogs6/Y7zFyDSxJfjAAPzaJwvlX1qrSXxoXK
D/nTrMmEbWTDMLA4YAvh6Na5uSNRbvxs+LVJMsZhGr5dB35OogGJeJc5JjEB
9ssACLM4HPQwHvXO1cIJkqTs44CXiYza4EnooecsK2hGOzEPnSOinGS81RJS
hZcUdLrO3CNJfRMbih6fG/x1IuLa/pw+4TvF2SjSUoAxBHT/YwPcpuLU8Jvm
Slr2bv67hdT/D/I+yaTJ2G7baWvivqIyeOOQyvUVSLjZ4VmJg2OSCALzPjdr
RL0rUUL8Lv/fDrQOyp0LJUK3HVoxRVWn9N/lbxFcpLIpiF1ZZAQ8nZh5PMIk
P6wpCFvdE2uF8k70OuuYcInaUIZPHlUcmYu425As6EIiugikdvpKweP+kIgm
od4Wwr+JrcnBqGSh/YdIVYNVJwAotsJxFwsnSYQYM7xwciqki7gWJk9B5Hi1
WFTECmcyqskYe2PBhlXiV4l2jMRUbRhd+vTn0OdtMaxIMc6uAbv/DeTPMDkW
rEgEaR/J/CQf4KjOJBdLkdrxue9Uj5gulHHUemdwwb2BywCmp2yJQSiroDD7
LhvhUDF6UK6STHRTls8ZL0Ojxjvy1wamEZrZ9f677dz2AcjZjXs4G/h2laJw
RA8X5Pi1lB1SDpZSV9KFm0JP1gvdn+C3L0Y+1dFi6kVqgzah2SauM6Fh8RHW
oeKuHVr8CmymSyt2tHdm5uqWKc+2QzrbbAByoEIBALCSilt5gndQIcpV+C6V
pj8uWEGwxuUxWGa5tcCtlnvfjRNEeiH7F6N6LCCT4vFZV6J9HxCs8OllmJGv
yQXGMtW0xhExroagRER8ifpu92IbhK2kAsfvIYWrA/wC5jzMbFMUA+eXDWVc
QcrAdVWpsSUDAzXn3VBcS/aUrUPAA5ZmHObKi60MSejr7WpZ2ZF0Zd8VNAPy
71IaCU7TIyRRK2JoK5jJw70AGlytlMWEs3KFROfMAjU/Otqx/RP1UNe0q7RD
YDUXiGKiWtKwEABKpVom9SUCezGNklphfcMXSqa0OGLrHpsqx/IIuQsBSj31
0UKR5Fb5Xujt9WMXxpe3t1CN9XJuVLJihsFAeKDav2nDPpZtKZLFEqOLy2Gf
hB2ZJs6g/YpiXqOgI7NQzWGS/1vzFMa+4wMLdpjGG31YlAaUx4mamSYEvSB8
2ugW+NyFAXVxt9ACcQHoVLQDWg+oQtrIB9d2GMyXX0jFWfTlxaACZ1yYZmr3
7WbfpxSedfKGE74jwSwcKVXrLenr/0hv3NZOdyllDG17zTMj1dB/elPv7E32
fyamuDkZwzzeZPRSO9rhYsfPE0eF212VDF/7DFIclqoXn0Xn2l6ubleWyZq0
peLPBzpKZQEGxxAVNQIO1nnaX+sACb/kYxFUFPmkhFSnKor5TmnOR5bhJunr
/ecaQ/YWnyPQgu1PKQPzKasxMsG71P2chDjvlcZz3tr3bSFBn2p57h+6QyCo
N8UmAeWbzzjo+Q1wkeBaGV7MbeRFAsFW62dSDKe6G0EBk0igV6/lcvyuUxMb
SrAkj9ZjE/ncQh7u2p1mkTV7bY7wZp3QQV3cIJj7g3Hf6hMB8RHhEyLh5oPF
rDT659Utwm45xHkdWHx8De7h0j2L8bhn78LVMKQQokziI67VQuBH9RmVDAAK
73qg0wNunHzk5S1OZEinYDHmVfGG/2CUkb3/uNneH1TwvXhcH5hJCptwhHYC
bSuYEdvrJpw598NL1U9RwSA/gvwVGVRBNMqjVDfFuNqV6IYQale3nflS7GX3
Hj497Jd6Gf9qJGzrwlWUCppnuPX7DV6/2igWOn9giu+H52HZ1mHosNVdYrlk
z4QLR7RQ3E8tlvDVY+FAzLiWPLAYnD+Nf7WACl+pvXcfZnNpw4hrsDuJev4o
B1vYgSbjYbmja+lflzCAOggzVioBoWqFEOgev1xeCHtcxDZs1GCKONq+A+N8
aKbNui+pdPFI7/wpJeNHi3Pc4Gh3chbqdpTSbeQ7/SJJbQrQfiW3pFlCMEWJ
JaYEsF++P+7bya4Mlwv9jh3NKjAbJVSEyhMzTkIwnHb+qOmn/RmqAR0coR9L
NGmj4wGppYts1VxbvLJSQ1te12JqEYFXwZ1asLqhd5tRkTstPpdnZMROZpie
7mu8faZlgybuc6Y6NwkGgWUgjLn0Ah08wkwQVR3wfpuBRFLS6oSwIKqZ1hCP
CcFu6U9mMtHqB3M8qj51hqBMHyOorX1ZfZ4eu/nQEOLWQpQcTuBGnjrokjb7
7S8u1dBXdjRORZiHh25VgQQQ/+o2bIWU7MfBgLJ8ZJWARTI5oEcgzET/6u4E
BP/K2751wf9Gdqt5Zll81fS589CYjRLgOUMSajO7C8MZbgDiHbX1zOL7GOnF
PogwnY/o+TB2oWuYvoT22QL7WGEsAbItwm2+Jn6/myJTLwlcGj2beeJJZBQ+
VDHRzrv3t3jDc9nc8byPNpyA6+ho7faiewsqhYG0f7T53VXf5jPl0JWwlG3Z
xnbyKz3wk8BC53un+HwXPxH7nv2AUVwSlQ/qWIxSZQsCtkaNvXRzdJfxr3xX
g/wcsizRT/Sar5c4nO6p8z2JSNUlaourUqr8Q1zjuAsa/nJ9XdmqLGPJpo9l
vK+Tbmtyxr/JteT8A9B22+mu67elPewQKkLQ29BFYvb1S4OrK7S37mYwiuKJ
fPeDTeFdrvBiKTmBxVt2t1YlnDBlpDODem3CJuUfB8VbtCejJvO65s/RNu9Z
tqUTgeh278NWR/qa9FPntdWLup0LZ+Ni4EG2WJMBHgb0hu1yjrEzoJEWTZbl
3DxJJ14P2vXKZUdWc7EZAOofStqLDt2RTvH3UhwXIdPrluf0UgALObYyklnj
bIM4f0lhEyXm4RBim4cfX4TGI0XgkE59hKciDOjMBwVm5Ush+jqWZEGVUsRY
+cU+RMaif84sKtLBMRD+5QC+hMtmcRUBTFaJaAmhnR7XcpAFE/EsPg+TKZoW
O8tX5uscVYrHkeewTOQoC5h1+/8orWoB6hcpv5G2uUvZPyUMVN+MilPDL6IE
zFi1panutKEFsmCZvNm7qpT6XrVVxbVsSAB5iMP8JPQsSexT8P7txPmlkwsM
PmksI8Kh9mVB8jQMQgpVEyGipMdnqInH+JuHY8qb76gBUVu5L7VsFvGqnf6N
IvDOYlOHpwiv59fnHapPHicb/Axte6ZCOTpz5Um9QbTgqyZkj3yLHNKDugK4
/h1En/9pjdH9ameY732UqsC3j628gcMpzcQevYkQOi9l75ptBJraVVkFuoRX
yExB+5qkN9wiSNlnh8N7ifYrMlvDqDla9br1Xh//N9mYOLN1ZO47oxrmMjF2
SYj/JPs0fwbsyIBnJx2HXe40Koqt+HoRdksCYOyvKQ65H0+haqViXldiG0IX
KRcoL2QEuZzzyANBd3Z4FGMC9pgvkNda/JEUjjEQJuFChwuQjFPAmIS91E5s
bDt3dY3MnQPyTD6Gw2WlVEUP/Hp6VoJ23ZoyiUvSoxPtRieZ2KD3goN5hx4o
HfNXJcwDHsBrJ0uQk6G4PudUYc9OZyF/bw3r/AVEnapmqAHMcgFXvzIpmNRf
FqR3xO6dQwBxV5ac1f/0G/C7x+ueQy0Zg9zhN6l945ZU69X9iTi8WiA9zOmT
lU9uxalgzSlSL2+gxloQj6aAf0+jWuxN5TBYW1YQZ7cofMoX2e6609oCXfzS
a1O1oGiUg88wphFwy4oygSvHzNLA2Xsw1xYHppGmtkiF6ePlvZrCJVAABzU4
Gt1SN+Jzvk6GQL+2byLN9+XO5dPdl2MrPRZ1YUJi8CUVNDKUV/pN8CGYIWqR
hqArVIF59GDFtmzaEuvtI5ALoBhMxtumMyuxNRZhB3Y+pQ+xLb7BPcQ0/jMp
UIH2IL7GFbvXWOSqXV6KCKuM7dsLJhfkkhG3fDiqgNLxL+8O74PREuSDCOwU
4+YCbfitv4jJJ8EjiJfAUtfQD+NX8pG2VHeR9QmVWYn/MPcZKIIw1bLKlXXn
aNcTKfjHE5hlQF1ws5LPADZOWGx4QL/BTr0AJW+xfeVKyUZ+/xulZo+1UgRy
ajBmCWPUSohISdan0X9w9j+IXX64+gON590ZMdycp/YTFcFG7klOZoWxxmPg
7pAuy627cdremireGii5/y0Kb83s5tKhgIjXBuf/v5N+J//Ry+fUofltLqLh
tnHv43/Swm+xnPLa0RlXILpLmXYG/d7vGh/Il/etgOROGclCuSB5lCxmxD7/
CSUiZ6crmwOgnYR2yhtEaGpslx8O+ItG9cMNMT0YTZUI9eMmH6MH4XaVuPqC
W8t+SeK8orFE7Nzn8te1SH8ZdBVCHY2nUmzdnjEwSvz1HdS9wIaPBlAQOjPu
hbOfGxAcOl9Q/wF11M/IuZOLF+OjUmTW39/aaJ4pofYc2yF2QLMCumMoO5P9
SX8CpngP5QGl+DdBsUlpoR3zGSYnuJNMSQEq5OXkO1aNMT4NEkTeRziYijPn
LqXr5v4YhgWrej3pW+rnwsaZ6dcBQBDu4jBbLD25FsETvyySxLOBx7wuyR8U
YwWww+9yMkd0v/zfP/Oljdi+Ri4HbIKF0I1TAfnGX92pZ5LYWEUzQlHCDIF3
JIjE1eEDfeejXNZ4azyQ2p8viHqPnMwCu/mQFWoVLzBjF5vFzXszU+Vbzm15
3cl0aBOxbOJuDxfdZvIf2RM2CVy4vi0SdqWG8exlnpIM/Y9JOkD6wJDsvuAc
VHRNPY4swsAjfwYSl1LIuuQ5CiCGqDzI1Hy1O+YkLw2g/7t5xXK2h3BOj/tQ
SpCwSpy3bcgF4fjV39qpjqBra1CeASMtojeWDkZLbZhTXqHduLKyXwOvOC0J
Dxu0Qdh6oFuhtt+TL3b7kEzyZ2DTHa9E5AlTaL+XDutlevsd34rvqgbOhmtW
+XNX9bQOVkZ6M6saTHZydc8mx4ByldL8SB/31VIILMLFzMuB3aB1R7fVe7A6
ftcw68f1TASX8dqgDmBiHrwV7FlD+plHfwGBo6fYrkvO/dKyu0hR5Gpwfcoa
3yMrtfnw7edjPrWNGpMhJp+O/m3gk7caEsGy0SfE4AfrodfEe1wpmshar8O8
5o5128l2ruLpCkvxsdyh9Aw3AGff700HITV/h9ODmBDMzqhcdzwoDl/jq7zs
J7NEaAuOGPZK3Lq+C4BEsuerP77GD1dNd6uAH5DylnvGcnku5suvI2xrNJoH
mNRJ+BO9P0yyG+BBA54zMyhiGmcnnNVzdmD3rsd8qL6qLoIjRfzxNaL3ILCM
593/rGMuUXe45n0b1ufVkm4hlEbmzKdKNM++dhWR7HY5Zh7nN+LJWiXv8O1D
npsBbyhrypLInnfrbrryhhGwPUuRRogGo+xt5S0p1pnbq4y4yPntJRCj06FQ
4QzUF+MVIpAVEqf42CjgJa4XxIGHig95qSPaxavW9LIbGMBuJUeVWf267zmN
KAfy7plIMa7r8rPbLvqb/7KxnYXgjN7/0grkD6nTW4czZ/pEi7/yOgQjnaz7
A8lep2pn2SsMVCbQLmB/6q8vlHpOnJcytq1F7HUbvwlJnnaZsRilORJk5eSW
ftwBSGJ+JNHSZww5uNOV89sbYZjigW/hijFSp/Rjb0dQ+48T8QsfBYj+clAM
HxEwiroc8YNjXyKvQZkdwZHs7+o/Uayuq/0sGyI/SS9N5BRIZk8zfhMCdStm
MzfiT+LrMAZUjvgOtshSOa5LhhnksOxg0AYB7zESHZ0ya1xy1PvOVSla1QyJ
tQyXFTcenFEHL8nBliMcHeqBLdSjnu4w2UFqH9Tzr8m+08GPe3AblG/w/zJB
oIn0VVM7tDWyRWK0AbYoaEo4p0yeswZVPTIJ4aHPz4k4XWKBP8VMTLNjKmpr
BiZBn2c8stzuktGxJeRfRdTDxV7t1xjLeGF29KgNvuGVHOhFSQRA9b/GGD8G
CJpkAwp/3CyWouSQG35OIupp2MeYm2AvT/U0lbSAi05E1H/owNVoyRlOoXGH
VfUAIS6lLnMgFPQq7V+vB8LX1QebcKYoH2Oj9lV9Lp3F/VCXeyxZaXh2Ff84
2Map0b2/n2j+mSJ8bBGoYqLBGDQCkp88zpBhXjV/xiei9VFC+7qRzsNjbVte
FMA0rZk0rJLeLrNpcG7UmlaYNo7v2adm8iJxRSbA6A6xOMSM2Uyng8ytYLwM
BTaNuuYOGi3GFucQw15OLPmLe2wsIPfT4MiM0o4Ypox91bRnK1dXobMAWVe3
Gzr13H5QBF0s65T7sTjP1grfFCw5adHVoUr8tTMGdCwUn+6boSDRe6qfcFxK
Fun8Yp4gcDLoG/47JwcggjySi4DAt2e5DN4oj7pPxk+XTlYguh639tLw2AN2
bKDKt3F+/dVVDx3+VrodKwMPa47Rv4ZtZhtY7Xvw3vrsVEMy7jWr2WbHFmma
1JrhtReJp6z+0cRfStiKU1s6C1jK28sJ4qBBUKDgfrpPqun9fTdrFepMbI0d
eweCiMsRfPcDgF7frT6d87r/QygssXb5xquYYNWnX79cAf35lgzLdQm4Om8s
aYsGg4hnI9krWDeeZKLoDQt+bc+Mud0TNt2Mmda9hiKoriOd8fizO9YKmmgg
Ej+XZvgbdbCtR0u5WrAoE8U899wSq57t26DqVyE6JrXjC/CCJaumvQKhTDVw
tNLpx7UeUJN9l1u+VUepcJtD5/4PJnPdsv8Z/edIkiyt91Gy/T6DEQDNS1Ti
22BncgqY+rxKZfPrY8IHEvLL/63nBNKExP4tcKm1uqJlg6wG8DS3M3jONQ/j
VTlcqdJn4KKyoKiDH9eR+PV9Pp9xBM0BFOIi0x841UHM9HLJ2Dbtj7upqQIa
hnimqa1yG3fkVHNeCZ2IJFMLMonKH+p+flWHoxfpk/xPw+pHeQPyNHLgpHnd
jEO7EAQp4I4xkrJXmNUqlxWgdo9plExxT0h9+yrPYO9cw49pQzxRE+oeCY1j
w2Rb0apsCYUJfSnuhdvSJK6pxupZBmYpO/8E081lW7WySicmG/rSZKUOiJto
qb+6lHACjFJfGHleiXpr1YIW0+qsue60xY1xCkTJLCNA6hZrpagnV8UN8cgV
CC/QA76UyiOmPmFcpaI3no2NhWlK9tO5l5c4IzU0tvpqaSuMX5aJmsOy2RXh
Uz4mI3pH1F3UPjez7+IXnzEgJUMZf9xourKarKuw8/0ZSEO2QMuZhFuA3aUw
GzeNIw34pwCquq0199fhuwOxZg3x29gAFk9Qp0a5mSyTRSHKih8dJIpz1t1Z
yVfTT6nekoeX/oiAHGdajs5zydyE3W38VK8gMR3PhqzQMPauJDXTd/JwuBp8
qqT88+RGXdLzOkKgHf3WcHlXDBrRlMCmKdnfch4fNFMH26yOg7OkhjWq9uH2
WFwkuZc2yxvdNm33fOer6sgBaq9eqQ+IFLWJfy/ClllCvxK3slvt3Q52s2hX
+tc9zzedOZIoIfPwe1iaUMxL11AWgC54fvu/Mo/UWRaP3o+pymipsJ5gb5cm
UpZvEfEYP2xIm/m1WhJFTKXAsbeX5RdEQY3dVq0Cb2GslO9jzp1rnCwd+Qrb
58jMDpgs9Vjiv8OTHjc12Cvhh8XtD0QP9iRIOr3zAJb2mXwUjrfFM02iLFZm
7cMKr3BKJCbamE5/x/u6je4BJhajI7FzYbHZoxsOS8LSVBbZkbG1RajPn6vM
m1mWSCqjCBYifIU9DpmcxTJuuYzsIxfN+rxlWSFPJEYWuT0rRMJcbe+2WG2m
1Bp22fyNltflnlQED1DLVFqeWAXdBrU/wY1X9HRJG2z+muzjzfM0bQcP06yn
RFSzcQQKAL3j5Py4t03ebKlS94MjQmZ8LzJua7bAG2UmNAfuRD5ppJtVNtkt
JiRlZBx5+ki8iX+Zgq0w2CdDVUp+zZNjGo73dbFaGAJ4KvtXfZTePnmn2/RZ
ZKTQNrDuYbsoC1Uj5x7FwpCRDmOYHDpRomqVC6R5Bzx9dd/IobvuJyaw4/K6
DJfYJXT5jheFGUnYigS9rgtt60j2VLAH9DWSQI3MAp/d9UOXEUvdNoBgDEFq
WTLC5xNoN8RlEFKw7dsCm23M8ZGgP4igUy/g5tEiGmQk1f6mbhlSnjcgH1Xj
wg8hHrzfyT2naRPEPZXGqpIay3nKHbpe3ecGrVwRqGnwpN3YxTE+gPAZpERG
N7+WESv+n/RcrtCZX7+vAXOCQNpVZ/0XSTkWJpn2mAjixCY/yUmDSYXxOWrs
9JtyLK+ArYEiICqCGrDUX2elmXeyp4Gaut+pqoIqgzOF2tqDylbQdhULgi7N
t2oWB4KqazIxx+bUfz8y0oWzCjycAWe96dPqKPCV67PeYXqoaEw0seehAXNm
yT7mdAq1sg+BfOg4KKFy01FJBYXON+m9Hy2/W0x4ZZgm2dxGRGrBth5z155I
I/1vOD7BVeeFZ8OhIT+ZbD13J2mL0W/kXHkRm1RzWLfnzBz47Guu7mYWer6K
6pvmKYSW8InhcP2j25jmSAdFmFEyJpcK1xy2EJ4WY1UP76IlUD9/uRtVFW+F
FdXUh+NIyKiRT7kpAJduIrwqLqte556s+0rd/atp9P/Vi6o2tN/9WNpdxdcw
LUwlY18p4EnqVljKqh6XzgjyEDY3LDY/3dxZDfRG2SOiG2o6d/LGVE2Awgli
771iSBqg6jDUgIHh6jCPLvlLWjqj7swNU6JFC1ICGFY3j4aMjZYI1ZIrdPwM
Z1HHq6Lt32Vbp5b4UBPcwTj8k90RGcdKI2uJhC/MBbWZhAvQf76UnrtOFVFo
1F5tN/9R71TzsRtgFLbJA1LjCvhfwR+umQ9cjVcgiYDg6+Ff4oE3RODk0c5j
RfA0yCrwInYl3tl/VcQhamLAypmR8355+Y/wEQqwW/AxHx+1rqR+qixvrzrS
kPYz3p8808SirY7IQadULtySke4jWtArG/NL+hGHFScvbYGDTKEF5XRP+esa
+n65o383GvbvSHhCffkgLCe5GplPuMM6Z7RPo7juxVe/YHi3dnF93+zDiLXu
hB68icDTMdA1EvwVv7YdqOa6obYEPdTy0J+ilRo9iZev9j5QRrFypCyacenx
hHMBF7+B78ZoL2ZH/m0o1ZjXv6y7nlOjGJG/Sl90CBxXylLhRQYVIPA4pyD6
QX0r4+fg0Pbd86zw7zpfjsS1DIGZh5NyhvNAzo5fLEEpIk9HnxCHDjnsN3Ob
wxQJ2Quk2WWWvj7njURPT5mp1jjJoFy6PN4DSraaYzw7D7/0cUt6vkHG2e3U
p8WXjkoDVY0RLl9419PxGhD+0tMJm9XN78+fY06Xrvk8QSa9e31tpMMYI4lB
HyVsz+knT9puNBVFQLqS+wCBL6F/n6WWdyOPey3nhJgQoxiEiLSs2dvg6y5S
Ofxp6hxzh6CfevjVW8bXhCZKk86PPG286Z2kR9aTG8RvgZj0tZIJTHnDQ0X5
gfiJZh9S5bE5SLjy41v0X5PEKX9/7Pdmo+zmIbr29ruLn2Ie97xGKmcIlwee
v5IQEXSIU2eyN5kGc/ycM8trFOaYIYej3P3lrdpvJjCqFcConMsB9iFBdKNJ
rV8DHt4rLmhl413B/Wxy2W11a3DrQjrHU3mq7XmyGUuz6x+xHYG4sUuVLdEh
zjtvmqPy4I3BUUrBpJ10R8q118h+SEqryX7+EvauPerxLwu7DBIMK0L9fLpS
DiLmj8pO+kOsxtOLYPktduqdhZZRzcjK9UCvhN62y+s374R0uOau8LyMLfFn
2krmVOde4NALFmGjVXsoBXatSd6yb1PhLDyHF9SkJZxj9NqV/3GkD5VcCpzD
dPrzq8o5WofLhuCHFh9mlOcDcbyu6Sp/l3NOrA9Pipg9sFucEjXzUksyfzOc
GGnoTW1gsFcVgODrzVGE8k7U0HF1k+VD0DSjnGSVrN6Q2b8QLorq9lpnrmjC
IaegjileZpIrEcgpcPVs9kiPNn3R8XatCvU9T8BB9LX6Cd4QDZdKHZPQZRa4
xFd5ql7UUjTL5qYK1WLK0vtT5rR8QXxu9qW/lwZ5CkWhaHmQFYPq96aIqL+v
y2m+08Xt46NgKg4XCWVckQP6xcUVHb4jA3ibJmsU549AzhG/Jwa6OwljB5Qu
tKWit6lA32U45FN9zjZTdtsRnCp3hniJqFRCH/7CnPXV6ORFnHVlUnzDmk3F
R1r8qfF0qC41ZUmPc1ptoLS0wbEN2Xnxo21FYeYC1FJ+dWay9DOyLxbjS2jY
xGaynu3Q2uRiWbXs7teo15cdyQCyN8XPjUZtgMWKglYXxTEmcsCq/eqacRXO
8ROMrHl0Lz9rjmcTFetBg1sxycZ+62D8tCDIh9dARlMyl123GdY2ciTjff6c
wixec3O25zlJfaevG9TK6ozrQlLu5N+OO5rL1b1tjtH67KLLEWdDWfNGv1jj
J9l9faxl56mlrZqK7jltPSV5QisKcZjaxCu6Qxaf9yqb+LyCG3w8cOVKAFyT
xbRFQZCmrh9qeyYZKzyKsZPvwjeG8hXRPik396WwXrvuO0DTy728su1coM/T
LhN0HJeIdhzD+Xm2FQPDWQmZGVZ1onxGfs1EgiqkP7ggkMpITkUI9+yWu3PN
DQLr+DFwBotugxoImEtOMmSQuxCAOHoL8WauwTcd31B0CjnnS4zd7NVLx3/d
yQAaWPJ8aDVt1Q0gdJeR1LEvjr+Y6KfYhYRrC6pqhWFwXXYENiZoIzJ4ZAka
7Dsucnz9DG3d9FZbk+Wtyv4TndXxcKuDsCYEvzuqtrrB1asEpPdf2TQWFgrr
q9llH6XIdkNzKW0R05o07uHodRWUitDCNfOy6ylSYlFvRGPUPQsbS2A8cwqk
jzmT8EDarE6/FpFL02W7r18DKNRVmZLR8WnYUwWuiiYEL4+LoYNgZbJmuKRB
ATFXNMV7rZX1VwWVTxwBu1FMK+ZK3RoZkwBZgw1++BEYqCcN2M1pdwBgs163
ArygyEiGtv6QiYZ5y6wFWq9i3vcC85pLi4cD/HIIau7rk2c/pF1M0ot+FbUi
/3zUkPQip0mKkLtf2a4OafQ4lpCA5Mp0EAcJQCsSNd6qhaEHHyMHRMSWC33+
mOQ/yBG9NpaUMHMfPhuBYcdoHuQeslOkm4IjPYzEyMd8Rer1i7aDO+Im2gI1
3EINIB1N97y27/DPTt5ksT56oc/1wyN7QJi8fQWHNsJZquCK+ZgMAJsvlK0S
PMlhFpoiEoap6T85h7MPMqsilzQu+cSsq5s6p+fdnCnSv3KKgRFpiv0w2Q2o
CSbb2+oN/729/m5xtJs5rqb9M4yiU+wTibqxDOCO/V9G64mClo6VsIMYjVPX
WBAJAINyQnj+eWzF24Z/5CrY7IfrRf+0hd6RvLrmipFZWrN4rPFKWRN3LW68
l7mBIHrX2gx0nz2cfEKLnle3yuJky/tM7KSfvhcsdevMTBMZB/qZUhO3jYdU
R17LqMGsVRXpm4sAppQeXkvbJRAMSo/g6F751nPG9M9DYdtg38wGRqXkBHGd
tbGJVhvybn9p+ZfHCQqKqHBSYOexxKW4A5Btmu2aRJddX3LtkU7BHeJm71qm
HzT/HzL6lZdd9cvVqsBknbqeVXXm4Ka6To0vAxRTY5OluP738kWW1AzMGg6q
Ag3ZBy6tEP4E5c5WaOHOREydlEV/LVlxcSd785yAd/QTMx6WqAPbZRP/FR+y
Kd4HYhvrNsnbyZ96Vw/Ui/cjZ6yg6PNYCzg1CVXfueSFY5iL4Sr0eo++jEtA
Mc4fMcXrK3A02ARZf+xEUpTyqTcYi+9vk+EsINTLBScHNqef/fBk8oX7/TT1
on10AyRTNjHG9/FdtjTpvnh619kqDxlo71kvBD8fZ7awzyvcDIs0K/y6fSiG
Ke9VA2oU/HR30FoYDpibKg8rbJLfW6/1OAZW8LUaSSoWAlOTWRXU3mijDmoW
tedTe90Fu9VnwYX3pOceCDIZpWeylXp+ee14kL+0OF+fnenxdVIrG0Vcmp05
TC8dMWgJIsBuR8QI93RBWYUxBBxZ5O7lQgwahxdVEA3NA7Io24R8FzEGuqCZ
25zW7r6mwm7BuN+Ygtcxn/YbkAel3bMlV9PY8Ngqzkb6sSxOESIfTL/iVkuf
49hBQhoZY2pS3PYiMiH72A/UNFwfzyowOf3SbrgqaKjZ2iRmXl1qxklx67TT
+xxjB1RKSalYIAI3s52VWmKjYYKZkSPIvG7DEsBVxsSAl0ZRerX5MJvxmhCy
7kBMwpFv2G0m3o+aQuMmKXPyO+p49LLrx51tlTgQkGZhKBhrb2P5LsRs0hjM
v59KJY1yHsmnjGmJLtUdc3t1V2MI4oDFpzxqIlO5hX6OT1UxcUJTudpP3xaI
ypyaw2Fz9r1q4X0ZeXvGzlfU4k0g+rdD8ZXshRjgug+Q0o21er2Xk1mLby5x
e1bxumA+hI6lbL7USIT4S0b5I+D0L9WHNJ3uwegpEsYrgcog+mO8HtzNREsM
RjN8rxrbH9px3xdUHluxKcSeZKMLNl6gE4DIQoKATmogzTzsJ8V7rmEoNAbs
3VLX/Wr6G5tNATQwvh71TyWLZYuw+HDaebvonEcxALuZNdYXQh8Gn/iBxWES
SIYBVsh4s/9tkbwXr+QDjkU7n7MfTdJRD8QHlnNX43vFR3ihNWwICs7qMkCL
HX1ENJvgjTqnwGeONsn2Cz2YcwQtdi02kpz44KGlBEt3/Pf6ObSyvYU/uEUo
w9iDSdXYwyqFCo/jVshW4lNMEkXfzpY8mIV6TdwAS9Dnx+Ivfbwjm906rtBL
lmXUPa9EZOxq9Ml15xVrfE7A4bxHQAzNvBXVhhlGgU2ayjjcMfSnA7mzTXG8
ekIzXlCdX1ko5Ssst/25BKTYmBg+h+jDLuzbWk0bXhYyLeHoKCvveI12LYYE
NHtJb4BF8WQfgZrDOX+ygscp5oNiod+60c7FhfIc9c08wGauUw0xMOLQIcii
SThl47PlkCnd4C1dp60Nipc49j+Pd/1aBYEIgF/TwQ9kokaJpVy6E4JcnRw9
02hah5TcKFTP+Y2ZHyPiM0oaaDotziNLlq8kbDRxoFaA6/v/VlykU0/61Z78
OH/2xIf9MStw5Fq9njjYCC+m0PM4RMpdtvbunhCm+5eEXWWttWl2VdktMraS
xXhRz4qNlYcWVK99XU5jbl06W61Jqzc0Utc92pm2sNnuEtG8bopv7CIAIdqa
Mi+pSAVcsrUi3WUcRhiSvCab4kcbpjBHJlUxMIQZDGIq4mVgqlimndFHOMxJ
qEzGrk8z97siSnUIB7PglS4nVlD4RtLWaGhEBkJXdDO1fy0X7Izst00WEUXo
5OLiJVvX76HeA+Sm8uL1FajEr685Imx0TVmFb/+CE8GS/hONhFCZCdhCKFQf
2pVNc2COJziO1SZCsrF8Y+jDKyFHHKxpkpym92IqnBwt+YgycEFy2RLbdD1+
wARCaEra4RgTLcbzaFXVpovo+H4TsDXGHbJvskVNV4/zLbHutfQWHMUYHv7i
sNGRX3cLF8UmMfiJxX+vfii7+44kPKZxweSCPrQTV8PQELOAgFM1uYyqqRAq
J25TWTVUy7kZIrTcQQqT9FAW3EK6xqh6M3l0vrdlYJDWHZ8W63edCHTyoOsg
ebN632GzcbEZwAxljZMPjb1wp1wp1pVAr3eCJ3EHp3huan6ZaanHWIZ4bmnM
nbrRdlOopQD2iAfhmaFHqNAZuRc1qRMELXNqIW4YVWXexZc5h4ZxOqKdHfku
B5AnDmc15hB/pMv+sTmwwenCO1GpToSV/H+RR41eh9OykAavJ3m4KGOF/fqX
GIUs0FVc7oOdpO+2wDOtDUVLhPiof/xAcAbSiwA67/rZqZPKhX4ACDqjlCM+
HNMAqNF9M09tpavXQMUsNERtGY9xIcKBmXo0y06BB3X82xE1u3Evo0BxJox8
fvQPqu4RFVZjxW2ni564kAxfBHSqUKj7bzN6NyLaKcShGOT/YfhHhwQdX+hh
Bg42vFVBBj3KwcOZL76pIq7I+h5kCr9GfBMVrqgMcfFtDg5sPT++woKCcfJN
qqs9khx39MCcHOKJczSrW+lO2gM65u1RA7PIf8KjvBO8zLLiSbvebUbBSEqT
M3nSOB3tRAs1bSvVj6ROWOaYpSZZoMJYdhOf6YJCn7K7rc0vtlmtUsWKq54m
s6fM76OoF21CRf1QsPo+McukUTmidpJ6x0f8er02F39Af7gEy31dB79C0pLB
KqYCQKGFoJeaiqOc/EOQquA7YEpPM85feIdIkWtkvtjuxtcTQPNqH5lruVlW
EqxJTBbbOPQUqEKaCGpI/hPnZKVpkyNvCtpsQLq2/bQ69/ldY/qSGFDQ8//i
Uui4InV+cIv1bTRDopar/hJt7PUH0ZXx42bfUAO/B/MiQ6wt/QeZwh3oU0uO
8m+ob9NMo+ZRGY6jrv9yhC09IGNrYYxMi38sgUHnhNHvVX92SIk5jGTB1yN5
82kOSNfC9o29kIu0hK3Vg+9Z+AhO1xYWm191xwjgXTALrZ8+wq1ICp4j9DtQ
Pdfx5ppk9SkVPKpQQNKzJAHNXwaJTC/QBj3FOLpPzDzhBBAJZyQ8xaPRCUyN
E/ApmumKk9rp10ou8g00Ysb/HoPfm7E1qL2N8tBNqikr0x5gf6S3pSuK/d5/
uWzxuZJUMul072tM8fidIt9mRTmTC7jWIyVngau6Gqi2XQrffXT694qiDTie
YmIvajszGguLM0plFnEVsQ8z7WvQj+uQ7oGdm90foW1jDvHZlP8cMDPKyJ81
VCfwQdCwgFXbddiRkoIKA+IDwPRVoU5c8+w4bps82/9UixtDrUImnBzFXGap
H+QutixnocrU9nExzNxBT3unugKE41qqocBq7o7rMUCdfrDhBEVufQipCizI
4vE8y9E7o1Cuwp2/QoYNxrD836oAbq932mSqxr4fGvAjecQO6Yld4uiRZ3jw
RQA0w3jbeOzfL7HU3rAzTAGttQDKmYLhtPS2KtcbxVDGRD12OtvgHl9Kd/j8
F6Y/kebAQMbtkEAHhfIiZ/vi9JuuDLCgcalVzJXlwA8DvYGTxPLG+qBjNKjL
i/75ITU4RLK/wEo2IF327kC34CaiXM0Ng8qLJYi2nnQR3RwZ0WHllJXKcKPv
KpyJBne2PPpmCrwVrqveTBNUtfLtO9RCbFXwCQo1/j3Gpfkn02+TGZLtQoEy
bttIPXn/riOxhgciQ81zfdqPLKxWnntZlogE6XnkufjrU63gwQ6RgMjFDRQC
7Nz1lWB+xrx8jqqxYh2U5RuFPcsPipx52qOkyS51JSqN4HkUByH/eoUBIk9w
2ZiANfHqQRj7ao15GcCpRLHZQfNa68pt8zTTXvb3kulZLKMpZ+6ecRrRwmEI
YxEu1ECMCcita1Be+oJZXi9dOnsjIEAwsvbcWN2yGgwapfjmSIvEodWBOXk0
7VSNWyf9LgzVHcs/yQ5dwpwoukjJjvGD54DMRBNF0veTIz8PQqIUbfAp6TGA
hZ/2j25HXTSKwCWzY4ROumHwrYDQ9lJN8Fz3myeRWk8lt6d8STshE3NvEp+c
8pjkFp+yFJejc//qrtVGACOxLFnQRUfhMJZwh2iiTswTmwZhMxUk/Kd18sB7
EUfczzNH0z4MUK8d4krvRzJsgPgYDngxiqik+KqjVWA9oyZ1xvFzhuyJGc+7
xIwwzd+veCD60iz9d2jcyOpD/Rxkmo8L9Qx85JAvS+Kqk2C0j+JI79PpACbH
UQAGs4KcFYlFVEMQPVEjOzkuCWpTR/OeffNGCf0aoWcfr5Cc9/xfcoxGtWpV
mjNL33wAqV5Aab0HkD3I23jiYz8tbP8JA1oIMRo3Gg9xwTxdKD8SL1pgar1I
tgLOJa9RsWcMxpcVV/s0a76YRfyVtWb2fRlj4eXpjuHomtjwtQvNLOl3O8aV
JJxO+19hE4oeExakV1Bgbw8pPB80IJW5x4B51sEi/yNObUYRcluppwAlxSf/
I6SFhz/SBBNuXgPM/n2ttxbbeXnMA11jnwnvj3ZIrPvLhLCfQoTRwnplCy4Q
1KRGM4fGfr4eRn2TFeY8NtmJ7mO7x/Ha1gvSawBmPtnJf/DU46xScf+aqV5S
oFZPP0Lh3gPaHxsFgazygJMC76lj2uRYyJarT0GdXJgGmqolrEE7BlyQwm3Y
lOJdRh6hE050OyypJjrckifP6edzdHiCKyVIt6eexL3njEln5omoMPCRhMqJ
Tffa/WtrqEpbttKM0j873MkUsHpC1lv0yCIB4Bsi7HT6Nr+ST6dpVfnK7ehC
/WYQSXryBunCR8H3RTaNuZmDgT2B4I5XFO00Z5RoKP1ehauI2Cq2TivV0zU4
rCNrFPC+Fl5+C/YfyGaY0LtKR2R+UzTZGoggh8qTPeCc73mGEh6w2alzQT5Z
2FD9i8s3NHVzIgUXeGq7S97rMTYX3UrCg//smYKE/rpPgYyk+T08ObjpLCs9
heylUA6gaLd+afStgOC7l5I0PhYQr/0zInxJXlisZQDurY2ThSHRgAIA1vOh
4cfJpgyyJTTxQNW8JqD7JEOjYs+FKPYTE1XQed/gCfYEXtJPt+LMDHNB/tUG
5f59KLvsZbSOSrWYXYhMTzImlU/UINVOhMEW2hr4ABF74m1/7b22CVn+VVRQ
3SVNp9jJUigbUXzFc3+bFNPNalt67nLsNqPPkVQuGOUJT/JBvWN7mrvdwSVq
QjBmbHm2HqZ44LetRVeGUXRIs2GlYvhX+njdrsIYwM+A8NQP1vfX+jMjnHvl
2AqffyaowUmohKiUKFUh+CXprd0VwtrK4ZROVPAMGSx/bZT69s00WSKHJ+Tq
PneWV8ljevr8Q3nsuRoVedliJR730whuvjns4yD9Sk5dUPL9UXpulxVAYwIa
C2r7HljEVOOI0PTYWE8/iV++4Av3eGZPk/6YF/DRXhbIODGmtJBvKD9GJp08
gbPnrNhputBXWMHlheDRebG669foQC0j3AxgLb+YDFORYCEv4Av8/JmW+qwA
ijQYnevm4gvF4qvD4BbO2TC2/3zIonUi1kW4PGkGncV2U+Z0PPIpydOJ71Ud
bot8r6H11D9U/IPq2zR12l11WYInPh5o4Vd2VxuHV3Ha02GCDaHou8nx5iDH
aim5isAZ5sZntA+YFbji+sB4EjxfDAVPPKzjudTqSaFz7pOzXheqgeh1c1I9
AOrZ6X0naW2KYgjXfSJzqAH6HJ+OnOc6mW/SH7p9bJOxzyY+g+cpl8aHTm3+
bJ7+VXBeNaeblfVuKf8Qu9NY43WA0NBTzbZ+nnZEDxG/sURQ0ekcJ5xuxaR5
+HytmPXfLyIaFBY63BXt1SWHe7n2iX30V/v8G0xhENgACOiRsS7NXpEpKypO
80jnj6FMoxAleuE4hJNXfNUPs6fCPQyVt+dqznOG8+FNXtnPEnBmrist8Eo2
LoMMyD9k2RE643SaibtEf94xPOVNaWoeUjUIyMATvYvun1SJVfCytJiQVXW9
pLCHZpQXj9zubxLrjkovb3JgHApip65BCeP2OqoQbvSylhTxX284WiBmjRw0
SKBdSaNT+abbSv0EZyPrjaYZWDNfAa/u8Dgmd9b7gVyU3zVdUTvVGs1de8rU
OfcM51rkHre/9ynAaZWSXaFCas2RUnoKN8O7itInsdY2IwNikXJjf+/WO5NQ
PWq6SDrNl+iy8ZXl4pBUF375W1bw52sTc9yS/tJi2KxH9AI6jdnesfXeXr8Z
DMj7VJsrCK+Q3Zn67EyeZQjwkEfeUM0a2W5A0bnkUZm4ZPrcvqBDK5yCIAiT
xteYzYPACIX1klvH/m5qDLsK/QdnF9XTfNS9OLwQb/u3YMoFz3rWWqZy+9Cy
cpDJ+hmeniuZ4oQwrAyg+SYCg9KaxZBbxOzLmfwAKs9mfxAPsSb+5K/SKlAd
MnkIeunKxeBjBM0jIAoJeIgJbcN05NETYUuVtuH8uQ+a3+MzJaqiFuEPyOSe
mhjncdwT7UNJsOqTZYslOZleRC7qZt6eL2V0+yiIQKGscTajfR8DRJSyTKIu
5UwYar+7KshqqPkNll64o2uBkww9Q+ZfyP7AJgn3mAcpaORwheSy8d5dZOvr
Oizi/7rPeD4PNNMt/Q0p4K94LdxoZndjyuiulLBtuihEHcoJNTVdahSzOW4j
6lCh6ZJAHuJAr8uv+npERiEPH0KpYsLGrkgPm97oqpGm5MRlGYmsIOZt98Yg
elKAYcEUoU8xPvxe6ag7glBFwXAGDyzUt7PaQU7UvRDg3+GlvIVv6O9N3DpB
tpdauUK0Grqjb7Oitliqdsyuo1IzsUhmw5BVjLNxJEMAtovVKmGZQqtulozA
EaQotmZvko6u8w2UC5YCXQC6MGfK0QF0g3SJ/Fsj1HA1DSvqA5HC7q62o9EO
LBX5ZKVvk2AisZrVMT2F3VFDfVsGxGiakvY3P+FK2W2PnhWSTVg+X/ECeIcG
mfJHiFIlcHoxom9/qRb2GPVtdLKjS+QeJbVXWIVn4+sJtReTQp9MKw3Z5hzg
v+cROl1DrImXHARcoIBk5CQZ9RV+yJkCnsKAi/T8DpZuxyFptFhjed4AJ6k4
aPlFBGehpwEGl12ZyN293sj15V1wrvezktKQREik6D3dcmEl9Df+hIom7hQ0
TfjFR1Fv4RiVcNTxqnJ1i/EWWjEYqm9469vG7IIko6yVwCCfa6JP4G57JJ5D
/ZtgsI3Q7DiXIrWGVdziezcHthso3wMgs6kU1otdYITHRFo6TB9MJ7MBowva
4lD6HqWm7jxzQctCuVj1LYzlm/WkXf/tdcwRL4idc7GCDVUCElRk4T+NdolP
2Dr5CqHyLyGwVUbk2kHydZ7HLPlthCMc5cFz++3fqke3RYOh6ANvm09D99qy
1k76lxzzGurLFAy8JyzZepdz7JlxQs96K5LrSeD8uSjnoq3IIdQK2ZHZHBqC
1Lk9ufosDbamk5wO7Gr+rDxmzks=

`pragma protect end_protected
