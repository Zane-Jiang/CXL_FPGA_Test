// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qnDSkVJvOVZFZnHNmoBiiJbFUNkI4d94PLHCpmchumdnZoBbKdv2Errn52h6
CZMU3865n37HTr40jMNOYrRyk4MrmJvYemtcUKnyTkH0DO8OKsuhfQoesfd2
TUZPTbUcwWDlq/9+7iqKESHUSRfkB4nXRHNpJfyy1gOEzh6M1ujaXncWr6eO
bXvpBAnHAHcrKUVVLDcLgsCW/G4baaJ5a7clKmhN5VTp9Rk8+aEi7PUMKl3J
+UjaElp+myU1CehZL5x5tPccmIX2V6n4ilWPK9A+2qPNqYAqoA/sTpW6WQRG
3aGocmaKPehPpx1LXEaYQYt/FVYMCFRSAyQw/CPCBQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZGkfRjZHLt4OTwnxW2WGnpq+tFv4B1Tv0N0P73BMQ3aPC1N17l6YOIge78Z/
Ebh362YHliBwSn4ZWUGPeC6Ov61+meeqBwpzuQqTPC8nZVVRqlhKerk1xxIX
MrF4IVhPGrawSfQaUYmcep0ArUq73smD46CWYMlQeUzKharBgGPCjmVxWJPq
LQ8omIMpBDcbc4E1sMa831pBgqMzPls3QXe0w+jqaDLS+ZWLU5jY26Lgd0SI
SpxQ/AZmb9/KOa1cVyqwjRhv9bgv3UQUmrc8H+Vk4XlUA8uGNyRIvaiHmk1f
dmMhq7EWyuP3+BRmFNn7YS/mBX4uizPHKlVirzMQQg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QTxOmVFiaLctVA0yVifA5Zx2fTH/eroaqy4rx8YEG3M9E1ADzOHr/eVLBPQp
nV3HsWOB2+2Vk7sg+yJ0Om8sKNPYU8Dz8LDrPfnrA7cq51MHDgZMJ2bnoUch
ON8c+XJVjfIxrj+NIQYjkAFvt+iUyNwndTVZEZoh/8QDkCuSHtydl5MWe4+2
3CalvEddE/uo7BoaDcvc9QOOkuPu9qZ1fOZpiGYgNegZHTKFXjBRYoy32zRy
qTQRKhhlLYroXkQqqTP2WLh5TJvdDmW32s+/LsbyHAWgRdgQ6diNVZMSZKRZ
FeCugD8Y4MBvq3fGuLxb+fZvt2YBQJpRXV8LTXMbaw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KXqrwncK4CxgM0GGIJl2avBiibTzzhSJcAuhzbuTJs0I0h4hufj1C5BlWhYW
0Eywuf18Cj62EnllcX2zmYzJJYFFn3JKAYDYam1DI1NjuyRrBRtKrhNTI80F
EIyRstZcTKAkDH/8QO0fWDjakb5qRw9jjdX5FTWOEpZVdUdDyVg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
koSBi80FPos1di6NbfDWgFf8o4kitVGQI8YcluULnFE1sPASwilpB5oeQJ+D
qbEBjkm4gXzaGMsaAQTRbHxjw1PYJ7aNC2XAyPiOtf45CkNOM78tT7orDhj2
FB2RVu5DV0exsFHeCc0jONptIR5Z9M32V5m0LWmv3tCt4v+wMLIfifa18Zx4
U2EVbP5TQJZEWqaiFUhpaGO55PDMGJ2iilwmvUc+Su9q2rz14A5R2KpDeFEj
G6ge3hCM74dUnBSNChb3SlPRBnf5eaVnVWCKPtoA7kuisKNXlswwhSl9NInF
zVDrZ9eFNAXtkP1BHFG9BzAHP2R1UicikBtqMXSDB+7TwLgPEdniT48hq/mU
PKP3wqZWW6KoyMlgXPrRk5zRmfrEuhP77rLAslUbqIN1CCAt+6lZ+QBS+Lor
a4msNMzkk1lo+G12mo6jyyoNtGGgGE9I996yr5YNbbbGHeMdRiIUR84pYHiG
cYs6bTnsCr4IQnKeQHTKFHOf7Yqgm5p3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FSZCVegLikH79FO6v9xPWDTxbiiYxYrQkT4/RXjBkU49ybwA0yo7gqE8yjPj
p91BKqRo2Oe2NEETceJWwj1clOLYy50by90/BFyUlsIz+H7Fkp05T3hefajg
f5tbhy4+acnB0TWTEecx6aIRU+ZYYeDETrCrlMvevAX14fovzlU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lk7R8KRX3JTdx4K3KTRDDVjfy4bckr8actSMbEkGQOGw4SAxapIlD1OT76fC
kBau/s/9+NjEYHsMdvbJ5kN/4faqlIy9BVymB4u2nveYu777i7nj6sf3yCc7
XWw9LJDjfQlOF7y+vkReIR0NwvErLzOmshXAHA7cFV4oK4FXeIA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8688)
`pragma protect data_block
VJNpbyXHHQoIj1ZXeaopxPMWgMxscqRm0yM/eY2r4c6dRpjCBlEu11zI3tzE
sb09HnLsKulX0rKBxxLIOJ+iPb7550/bSPQgzMC7ZrLaAhAmdaejtMgRYmjD
yM4A6RqU6T18Hj4UZXE727Je48xVDn3sXKQogqIBBK/xpTXVTkf92XRLUHYw
qwsnkLkKniwLnw70ePGUXS2vZhXbSB5gZNGz/FKgV6RUiOS/wkjSe9hpbxM2
fnSSAzuK0sMPCERl9ZJQupBdJjBKS4Jp7kqxeG6ZOJw28q3tJ9TUpnswKjVz
LMKcbpOEKn+O19+0B8D/RBCU4KSxEPScvhj593wH8mHio7om/l+Z6AcwMqib
6/ABQ/Xi3t6LY7MRYWzyG0rBm6MfObrfSyPhieyFQVEOry1sj3eJrR0ecqtf
bcTC4EN1nB1JalT9zUbB3JYcO9PS0ur2J5NLWC43gEnTw7s370mM9QbQdPGP
ue22CfUT1U4BxKY5ki4X63xMg7ZABdu7/PCPt94cHsjo/DvDq7sDc/AMMQR+
b40U1sgb16nvR7AxXvqbatB46jil+LFYsijTB9mlfHb9flqwRCFhxY0zvVIo
YMeNmrD9iVshhT4K91Y6GggP8Xr9OD5OJ8wXyhey9KDPZGE6I0nGcDUj2oVQ
lRRrMnDNHPh/Y2KkBOSwUjWs5LF3PNz7CGtYUNwpiEeCOZ5+rQNPz7sEsNxe
lu2xWMm5zPBMwoIN+x/D3ch9uDmip8iQ+fd8p5sBmOsAo3dy6ImpxunkGTPY
K9kPsp9KpcP/j5S2AdcmmPl35cFsGh7/fmpUd5bZgGsIJczd/bie7yfsz2DM
IBKpDEPzK4KAn5u2CAFrhS/RRBa0yU7Mn7JJBevaOvO/hrIOzUGasqH2v8La
Ih/4jmpDemj2+wYcfrT6yoALRlPkPplBpKU8JiCxsG4JXGRTaCAV31jpcTpq
gGmrhlIhVLshGn+1hOwoAV7bszK/r73gGU5H6Qdxo/Zhoxdy/JEz+Xy1FaD2
kBQGiShrJBRbQx3K8fERc1Caq6ucZFn+7r2gJ/bmICZXvfE0cUpWabgLHmmX
M1MuXNZsqFamqjIW1myMpP0ZB7PgqEz68zdkJ+pnQmgAzl4ipVM0VtOlBrue
ldR4BXN+GWo20nyYmj3Tslunth0x8ehxE6exAdiaVskUFYg6+UdwoGVyjg4X
d763HMiVCnATtjkFnLWwvUT0Lt4/pHTYAcu53H0zu7y1tSvF2ETw/9iSm603
E5B/nYzANrMV16U6Q6395eJgY7fWOOHkdRseTA4vYueho++dUihBDSpikmfa
s85zmYeg+EhrBFWkIf15IlX/JkGZBzR4Z3vaE8/oRU7kceUA7faSGSal84Xg
eEyamj+epvKb1U4YXxiSU/UzT7tHBsl2oGgpL14VahxV5rzj7GaUIqtyfczL
mq25jqRpTfB5g28vVTGlNUgfLuBvy3zANP9BzJ5Pwe3RsbLufhnLUbcHpHBw
KQqFTnoN1hgv4Svd5eP9kcH2EU1/a0yNr/0yxYqBKI+3WCcpBtO3D9OSKQC4
5nQDJb6kr7yVqPG3XyPFo6eilLibvmFRvNBh3ZI9W0WQkt1ERnpZO0LF6z1f
C1SApMb5FR6ChsnyVLAi1w8tXfr+z4IgrZGhqmXDf30Q1rP00KHg+hM0lgR3
wu5roO8kcPu/skeKRo0nwUKvE5Pl55jAT/fZxq+7vWG9uy1OmIVXJ1cPTZye
1mccNeJXwdhaE8Ls3P2eJzL1EW53mo54G0A5H6oNAb2lBVU9PZ/bwXv1fvle
cj2wgeNfAC4Kl1NPi57z2RBlDW/uGVD1q9OT8h7tg3w6XPsBzDhTOd6G8245
2WW3MuQt8/x98IbbaQyjbPbNU9Ckq3qZFvKi+8GnVKtxV0nYwFqgr60ct9xo
xfEej3J9Wpqa9waO+IWeFoEQ323tu8lXJReJyeEpvnnkzuv6RVcTnyMzULf0
MHU6yZmI26EuhKXNNgWX9dPdMfI8Xf/1Ci26mfng4t40UaTQziM20LbL4FUL
O7ITdIJdlRHdFe2R86fgSumtRob2oR5B+YLW9P+2yDUzFtZJubhJCJBSv0Do
1ebr/pmvHayttNwIyEg3U0eZ1E44NDn/MlIswORMm+XS8M1Iup0I2YEvfPC3
L3J/Q4CxIPmgfMoXWosj8hFQTNSVR10mjQsDgjxM5A6xakKebpwReWRjNIcE
CU3OL4xaOrpzZv5nt1FO4BWYKPCh8Xc5tweNX245m+oOcl/cN1NzZlpJVC81
Wj/Typbev3oMMtMpE4OG7g4xAohAdKCx8Y60gm5RBEZhvmdxE/VLkqOQsOLq
scqBP5dE4inhcc3X1NPdId/PPLddVUX1QSlTWXO5SX0MRhIgWuwzK0Wowo0W
YFLxblU2nv4SVrBlhAvhJcICE5enQZzjA2d0V/jcTnCxc9Z+V5rSyvcet8BY
ItSfc55c8hNnaZ147vehr0uXt60w4JkTWYgoHrohyKnELFNPpHCJQgKyjE72
bMbuEW1bgbxNFNvSUiQItHMTrB3lUDhpqxSMZ8GKquapXn9sy3bONZQiv6l0
PFwTph0Y9kdSRME2NnOgUw8ijZa/KkO8f7zjgtNjuQhNtwgvwiGgR7D6G3G3
L6OF68hcuTUTqAsRhAks0ofBfFgsOAttm12yBGP/jeQM8/yDsc/EzxFwFk8n
7Dhl+f2QYN0SX482XZn527u+KWkny4BUHsQEIufBLljIhyoUeO59rIUoVzcS
lVYnWxkU7s71W/aiyRFlv6qDqz16q9NiD2gHnSURDzdH9aJYvFrPPrRDmmTC
QRSnGNo/pLHBw6z7TvqK+I+iX9GLKnDtpNVYcZTpJbbNyCdr69mhmLT5EVwe
x7J6W8Q2ypMyW3AzJMywGYIBwvGeAfmS9Txrq5gwAJSDlu/Ql28i04m2AsO2
3aB4vu2ge3r+ZTmFod7NSWVG3LlXmyRB7KlfzABQpLmZ9mm37GGAFi2ri86o
9gcd80lT26SkgFfcOGm6a+WGVvdCRP+zzZZkSdrwo1759FrcFfcT0B+pM/to
+08imVczoSJKU/hZit8VEaAL9BquECrGtb3x+UPYuS5ilGrU1C3E6wD+eeXC
ruOQ6zkbUgR2NE7aklCkkCfjT6HQFzDuQ1dy04vzDqerkKlx6uQLKxqTcIew
KlPPC0nkPu86k3+W8ZyBNbD6JvqoYoOnZzLmPnT9bJthIOR0h37mKCZQoy3/
d80+crWQ+McUzpLIdYtjwMPzCKKBNeKI5i/JvM+WhUquq6JQolLlbqKv3xHP
YyZuc+a4ciskEMwSuK7wa5HtimAL/v+Xl6XiN99qsqGac1DLd6uIcBKsNL65
cLv43rlnTwtQ+vu9fuj6NEUm0YIedV/Nqr/DSIwFdRiFLUikqbwcRYvDZJ47
Xt14jN6KC8jg1gN4Q/lOPauaFliyKIrQWRf4jye+MtxDbd5/y/q2bkIhaSqe
bTTakjcKz+9TVRwb5EHzswJ7AGQqvP149uY+0dBgAiZQeefSQ4/L1c3N5Svh
BdKU84lvWcUdmMIFj4JOVA+MoKl90GyXixK5fDQ+tipixefHcijWp/HvLHRA
tq2CLhLmG/6K1ylaXZJpxfGwolxS2Et7Ocq8qk2PAiJ4pCJRFhR+GzHu5Q8b
asOLoQjTAuo9y3f8f6PPqWybCe/2OUkUZH6xSGTGh/7bNXbYvNmJJE6jzSSL
8J9uqqasjPAErhCT+1JPCRpiStmhYH/Q+KaYiB8AEJEqL2rZNio11aWj2wvR
NahD4kqyfA234KQ4ZOL6AgAVZUrrdtdD7G6gJfN1sAidhmyyWDI5dAnJZZ+p
q/gTXYN3rbQEbGJv5Mg+QhOU+MZVkh3uBKYoDhq9mb2kYjgDTIo9FqS033Ir
qxlhwQDo9o09RAtNXlH5PaFXKqbrrSa/x/rxhAEwN2ZHAcf5yJBQjyeJ7AY9
lVGF65WVlybYKXVpvDBUa5mxRohIG9CPUyTNe/Zo+Ehm0lmj15jPO6R43V+U
M5hR/NXj54vvD1Fmphdh7PvpFT+Y9qlbzlJRp8EXxgGodujJC3jhk7WWE6ov
Io5MUyFyUlddOh+oQiBq0vn3Nk4fosykW27Uh6RuA5utiEFxoiSJiXdEn1Oo
0OkZghT6OVXRiDh9molEAl/0FIXgjajohI64pJ6mCRD/tSALUjT6uqSsZRi1
BEWDR8+5V0VcsR9Z0gj4jPk3NFvvjhRA3LblcQHlH0B/9BGIe8OhKwY51Tsd
Dv++wxxVtQWIth6sCwEKBMmsQ63p4k9dj2jSjCdCPdoBn1hvyVsrHON+mE27
DBd4Y08kHsUmYSKDQuVaV7NNK3Wodq5o4ismSsA+WgBLcuAfAKWBLecjcF80
/oQFQa+UYpqrxJdlvGhBqCZ96p1DQonuuGzvPi1/zjljiy8660c1hiNge0Sr
RRcS5mN03/iy82fMTV0JrdNbJR8U1Dwx0D2/ACb7xJuzHPfDJWVEfnxu9B04
SovG8MlXTjxvPOWV0YNG3H9jWGRIvQDNci/VpJDZiZgDuxWEuzO1uWmQcF0z
PmvalLN1JbnSA4KIonIvopbaWM2RXSaQqG+ngI2l/AZLJ7vKPtb5RsA4aPyF
YRe4Q5vQPiTBdPZxG8VQR95FTcoViarQFlG3XdZM+2qu/PSJ/HriTrLKTEmz
kzw3gdrNmCcK3gI0VUNgZP6JiWr16RYfflPtFHoawIDqYJBCnZlBMdEhLVRw
aFxpXrZq5Ui44vskQKZ4B+Wsn/LwcmF8eT/W9o1sFCW1xrg/La+ka2v1nrAL
YbrCkgDiHs3VhwbfBh+ErQHyAGpOkod97u0UWEgwL6HVvtQsLWjWJH17OYRT
7gE07Dm3bfxDI1CHM6k8EE8L3RIPyW+fDnoSQMXj55Lr8nZMtZv+1E6GcLid
Ft2ScnsEMU2SdtQgmFhFfSh6Tu8uWXl/4ixcJ7FxyfkQ0Nyrw82f5rxw1f9q
YfAFixyEQD93G7lC0B5dKD5xSWlkGODoA0PANP7UkDYabmmRuATLQfdcdZNP
RNPiHTzIpbpP8LFrLnxgbQvgLBrSTO4k+Q+pcqwZmIH+PMy+dH54ud0v+xVr
wAjtd1YquZOFdkfETvs5lzYLgpiO9QU3l6jlDDXka4f9dul8L2zeq4UktdVs
YWP78LZD+rLs0v7YN0BRN4QGgN0I3LLGqkXxmDHGDCFWyD4Zos7VlasDlzxr
ILgIduPixPk4zt4RnPqasrpCaD8UZM9GyCsFXVtA3ABW1BjZinGX7MmcNmG4
NtwrimK6MjfeWsqMQLJs2+8zfrziakeCV6biTquyobS8qbBYDNf3dbbuAOYX
Hj4vcB55ThnbNYG2nkAMcy95DeEwX/EOE0aB4npj93PY98L8LYImi0sBxnkj
uMyaX+clUHNAsb5D5CnpHNEtYApUcoIeL5TQCGgF/DZcIxUYjCUIi/N/yip6
rdMflM/LAUEWGt/GNMNNIpztOLU01IuQkjlriNNveZUGXz8WDkakIk5OwhPw
OjCTI+kMo0KbPWVnyAZdFDcJcUa0sDD3QnR5OoVzX+nKqPpdwObj9+zTTMb+
h8q+XwfRB5q8pqVRq3WHL/RygpQalECotK+T/K3TgDbGu0df3T1dOMwNYgdA
/zZgL6zDtJSjeVWitswbwMW2oPBNqRORAIyFZfL5vweUU4M9/da9t6buUv4u
BeRFSaDxX7Q7nY+8u458fgCQfdAynFd8yoQYFqqjTYQ76dCmH+5jCAd1HKn6
oxvnbZYFFBXiKyNFu9sI7mF52r+mnILcZOJsj6KxzLwrYT5KjoL+/li5nYYs
hXYF5G9McY0XG3uXGl0XK5sl/pezXOTubnXa3AKZ7h2YEvAbOuyMuJZ5GrNM
CLF50Dwp9AGb1JgErlwqjydFiWgw+0bcNfeqTnBpasSKdexd1e1xBYlmaZyz
LlAFu8MFMoQUdccOy4FTu6AbZp/GwvN56rZpCJIp1l/OiD9xcIdcp2PuMxt6
yB+MSGzKRoUQrDl0+OxuBTR5uRpfNZjg7M7aQk/U86O91RLXWJJh5Y3eaunA
JIekHrMfMiOAwRtGtfgw/179XIgM6JaeQPi57kUNGgy0oMFdL+F0Iym/qy3A
Khr5/dEDpeDGQfue3hIXDcs1kHMAf+gpzXDhIVbmDU6eQHif5RWVZdvIq+NH
dJ0PT3QJkL+qBY6JN/mJq5MQMISvyUTdu80nAoqMYRFNCKMJQl9/MmGvsx9M
KhhEvOhQK6+WWEFqr/HRQiHK240L3mXFSpbT7i1fKrxEhMZeFdeKk8jyJCB6
MVlGnz/5usRYI8UYlFZkIlDiGBpMR8pDaMI7yu+jxn5S2zmbLa35Ach98pp9
b5zfcG5F6pI1uhdBg3zkndfH5oJDwCG8HFjyjKCqn0wr5i4DGjGmR/c3V5zk
qfyD6XzDkLGhwIIRryWXQ/w+A/o5vfK8klVzqN9kGoqUQolpyCJmHYtqZOau
dhTiz323CVMkpu6gjI5Ic/03+5aNuwsUkOMjjfY9jcyVLYo+vv3FWykgzlDq
zttzoSWprZ20Hl+uHjZr5AgTEsuGLzo14fg/PDWJJ/jQUdK043zY3BPPkYaG
YhUSFllObVajdWQORiMKSjNsnhAov7KfWsU5T/VzC+C8ZEEX37dCsuf8Xjt6
NEAEVJizTQktmnw6YXwkXUQ9aM6YXFOU8YmnaVegkCHR5njQWHW1j3dCo5Y7
QrZve5WojkzfNwlMsXFzA/4ZNHQGkRVxO1CnLAMu9ZalctI81nlLeW2ixMTP
uuiCfLuahLgCffIfHUTslrLwnguT5DPInjscN7xFSWg9Vjx2wpg7xBs1YBAu
09M+Eo3ka9r2AD16DPuuR+jiZGS/GMYN3um8LGcKs6EN3/VRFT12AaCE4RUc
M18bpoa/MvORKkNbdyb43IHkyTYX8G01oH/Q6VEQ722UDgpwucEiFQ5ViN6/
9dCrwgpen7tNgLsnCnsCmaoqhuLJzCRA0oATuFtflObUhF1z5EMR+VcutCRJ
ugReD8wo0TrIJhqpziLw0iU1rx8tCCpA3dIneYGCwJnSMvr/6/ksuAs6XXSJ
kg08/qqsLxQIG4tQSS+sRpGAKUzT5jvg7NM1DHycb+yDNxZmqTR/VZvO5i/Q
n4JZjuoFRjhmisfYgeeqyCWJ1kj7YeXHbfLFmpym/LwKxw/GhKNcZIKsG8TX
pzciwnsfEbh/Fw9Y7oz+L0HFXXjEzeJGA/3QdUnqlRPcQw4bL4ab5L1dkzVs
q+02prmGJBOYqtr11bDSLKptu5QPVZInDVytjInOLZambzQmvr+SzKI6erIA
IOaf95cGDxIJ9/qvLTmdPbgSSY2i5pf6ZSgFmWQL+jvxBVBV4C8i3K05rLKQ
qQDdcDFKc/F+BC1UkNwefvb62kKVeAtNnjSxlkBVFsHbZ2KZdzXFhvOypRLP
Q6VFiFKT4eTfmKzsz8mXVDPtys6gw5VFhcT4w71MWiDpSQV8+mMBgFU96Vlu
3tbsQKsHyjll9rZo7hBlKHCq2HA2AAHhHwggH+Q1Do+n0MpymBxhcXATV2jM
ivHkip8E94WISD6nwjL8RPqUwuWURqP37LSA8N8N6cHOZ7Pc00AHmQkHlq7D
t+lZB9TJiu1OIyOTeQN9V7XzViVTDiQ8EIYPqUN7G7ARrCQe1kim2SmMgb+w
/g96URBmpCAfnhCpc4OV7vmdeYd9nZt1fwypxiBEGPh7byNNYqpADNeKOWuD
H3JYQKddxoYQxpOLtrutT0ss/SVb5uWGnlCi7M2TbnwHeMWTcwKjS5LBp9GA
iTMKM3SWLBh4DKFYu5wJx7azaG/JXeeQm1skDqpfxct2TLPyjhLf8w0VBrq1
/j6umg+TjkFOr498GYPeZUrPx4ykz88fAaK3cZoD1utGMvKc4j20cEcwcoMu
SLTUB93M4814G0DpE43JzetjlE/rR/3+FevsFThNir3H+tBh4J3SFiUxGJ4o
okE5CCtPL2r/Qcx/gjBVjqzLR35h5rHA6il5hoTV1ZIjoouuwjgmatNwyxvl
Iik3i4Wmc5ybYZ8QU8+CccfeSFacp0YuSwXx0PC05Yru+8Z02tfXDVpL8uUb
GWUiUcSZJhTQBDzYb3Zk1kLVog604/U3qrOYM/X7TAUjaXQ+W2BmGZuSzkyH
6W5dATwrFZbp8uZAX38EIg0oLQjmyXqNdfXDZEHG7pbh69ELSE1sH+cuhDBX
fV5rnHqqzIoBCr8ymSfgcc4KAgQKIcRdTma16qvFxYfNZQJixN8bgZl6eaCv
kMUJtUmr6dgLi0+qgC31KSBLn/OlBx2hVfcD1xqytucqnokBFJydVIre22BX
PhF8qXTNosC5MOFcHW/FdyK8DMMS0QqvnaioYvVNEano7yFORzdeuxg8kCwX
qsDEsT9wHcdm0/Hdd1iG9gHucMLYkOV2ZJ/oni/qQtKURohbX7efI6rvzLRf
WHUPJkFqOqs4FJx7KkGnNQeXrVSpAXEHhTMycmt8XJw8/JxvnM5qjqWst+Qf
qX+D539tIpxduULMc0M+Q4z0Sidl1yJIOjXOskc0nOjOoCBVZuHtKskHfd0q
nussvSLUL6dBDuIRxhpwIXZsGss0VIs8DCR/peyuxKBOGDjRPoZ2QBek8aAQ
1UJNeGCeAP0J73bGjgrGUtzXVISITqzEckQ+8ApY5NXZfl3MyYb8QCasSdJu
7iHmSzaGekDcC+8v40QxlERRR1UGB7iAWdoXVyxfQQ9T+xvj7zJrMTc1+3Ry
lPS3pj2gLcUF5U+Z+CiYxAT0OtucTfKnzh/b11SjUkTKmm2FybbrnA0wALAG
TbyvKFsodfe7EQxK7ES5xXrGtNpdYGf06wnlwQoEGEB+reCZw9kiH+agm5mG
Pc2U1C1CjNqWvrO5SX0ghNF5v5xP4PfW/qwbFusbv3RtRqqINBl+l2b7CEo/
RMs3EfLtAzcAlFudOkcL7X5350GnxXeSTE4CxuM/+YeoBlxzp995vNiokSmD
e+8Aevd1cvwNG3tbM2cP5huco3sbhmrHudsHSgsCcng6RoKA553ctyZcjb+L
cGGrYEwuvlBmFUDY9UEcv8lzMZ30Jf1aJOpUDA09kQiBovh5wTcNcC+HJ09+
x545MgGfMNMeJRMeogSnlhC88TLY+rPQkLeRcdsx/uQmv8AxLyGaYm4HEIxm
a95FCgwEs8tFb5CStQvGXq8RlIB8ict+FpqPaQk5Er81nMzAUsyQaqQ7hJOS
MQ81FqiRIIUYu9B/4pEc/hESwvsrYzWssupOdn8S+OBrTeMwQLoegYJp9EOr
cDqaC3byBvWgaeb+PM8qbxOGZ67kHeQZZObQVDdNtr41xnc/1PSCwtpJLrNh
gHxPQeiUenv2lnV4UKb5GHFP6N1OWNrRQS3dythFLikUfoWCdLYcl1xYQGwL
F3e0VrEAMwrnaU4/jW1umwUCeDry7xSnbLY4otSajCLP5unzJezDmOoPGWSP
l8uY+Q7vbwIR5KriNvNBnvS+jEmlivbT0v2F4HuVki1FYfpqH+G29ByRUnYV
x53VRQQx3pPvZiVul2TaHWGgmCcop6TiilOxV+aCTeQvnq8F7vrBdD7TL53Y
VK+Rysu9WKDqyNdKfgbTvZ+lAtczwkICPDfOALluyYDXvZjGhZ66h24HnNSR
S51N6zJnVxDu7phTIa47diMQRLBuZPcdkD/t+jlD/ekulwSy4ehTST9Z0x0g
ZHmPdfNoPqf28c7urNFnz8gJYF5LcSSOQL5Qprx8WNw/Uipkoj05/WGpGZ9Z
uMaGvIQVipLJPW2YPLz1t3v2Rkv3Wl/e8y0saY4/1mKaC3UIx8/wT6O7rj8i
JA7iz6wbXPI9o+CVyKbi2t3UZC/zrVHJFuWmhVUAnnixkiyiQ5R3M2E0JHJe
kzNrToeUQa1F3m0kp6nSaWYWnqD2YXJL2MGWdd/mMxqaIfcuHkvHWXg6gq7d
Vt5xhCC/0t4Prm+RQtReztD9Bfk2anltuV6/dT3cArFTSVhu+3t4WRYBXwqQ
GojJP3vbTO8USErjFQNwpF/EhmRcJpFteBboYy8MeAg3UBxbH9nUWcf5ahO4
mvotCcqrB8yObHq4ly3kN0GiMdZmKWMv1nBYy4/mtFcbDObXf2ZHU8+zlz2R
Ksov+hYFHc2uBgW5kEMQB+QsP4KQYh3TbZOejyX04v0jT4qtkkqUPH3v9Jqd
45c6q66RGI61PN052F50LsuyyVcSKom94YGDphgLbf+X2ctAo08DA4oGuHgq
K1k05RGyzfcJkIbKXNR3Ni2c7z4yE6NLDImvhQQvUwmUwT2UFjE6FqByF2a1
1xB1Ag/53W6Yc4ZUnpH0EUqFNRncfL/EuWYzGHubW9r5i8cKl8MCL9a1UrI+
6bRd+qKNqCq6MrYOsYvAtznmx8vwgT2pTZMlZxRVU117TallWvXMnsyVj3R7
7DmblRSOA0NMUxVXySBvvu1O7oXXO2+t3AoIajdGxWUqM8SrW+wfxIdV6cUe
0A3i76bKNoqmn4WvjAP0SZDXws7satKX5OJTNV+imu/73rGCBr1D5e1QwIx0
4hzaUHc76FRzqIrfsRVzIDdh5JTGM8ViyCHC+x+KPiAzeQvxOzvcEYI5NQpJ
RxRQGIaY48z1cyJSUmDrHwIeNlqL+dfMRk8T8mHbmQOK/7V3Nbsm2K6f4Yz0
cP7Oeyn3TQD0FuVoI7L8Fjkfg/aTX1K79SKX3VDIF5uBabC++WSs8rcWBy4h
jXIAMSImnN5XHReOo7HZsKtJoq8CyKf4jSeFWhqecjre9ux8ugyuB7kP1AKZ
hJy4ngiIwLihIULq+BVYzc2VshbBLoaS9tJVUaJuCNRbTUR7f7YbhGAas486
9L7NACbJxgsWL1AifyemrdWU825xv9uSpRUM5A7oXVS1AAJVz1jZQmfvDuAX
1/7Qaumai+2fX95iGb4uXmlc/370XIVP7pMwlkDlrK5D/u6HASKvY4/zENM+
4mmAZo7XcRQdcmbxNNe8wm8j4eh3/cYODK74fruNXnLBmZ1UBDj5UPiHJWsH
Gqtn9YNAMygOqG6UCA4bDUhFKjrMeaH1PY4EoBpuUm7AcnNgL9tK1Mj1hrMu
YEMAFbmbHedL85olnIBA53NGb3w+LDYDKsZHa4ko1OXUJwplu9E061yh2y/t
u0vc/zac/N2QwJI5/4eVcIr9ImmpprZ/odw1JN8y4mJMpAsad97hCnbvm6kx
uGSJUtOIL5A25/Aug59RlMUb0S7SXE0O00/We49urzvK2LRMY9HGoJeeykT2
KGc84TZey5iooHbXFYCtv+Unt0+fDldmqEh+qIJ/wPX+0gi9++Yj3jtkXlzk
qkV7q8mIjgZhvXWYD2AGVjEsPUh+hzFcW1P/GdcklxbuuyR6sz7270F4nTry
Gt1JC13mggHE2ofZiJ0YGXxS7HRguvTTFNDsafiAgeqnn0pRpbCiFFWQpZNU
rI6PY/cBQVTzf8BGWg8A9mezkgUPghFPdFhnxQmKBB9Hr1mZcbtEn8fMpm8S
BdSePxME1NSqm2XBcpIKxxwTTxrudIACPlI/FAPF8ELAQPGN794TB3eP7pAA
B+M0

`pragma protect end_protected
