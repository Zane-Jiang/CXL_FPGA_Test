`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
nDlFM0zNHz2+ccj7sqAS4OcGGdSusAaIQoh2zHLs3IPIupX0GonnSVELcrxsngn5
ni/KsBqMV2e9m156UOjV6YjJwixAMUDwOIZUfKe5Wc4J+zHvz8qlwaU44gOp+hZO
XEcQkyWaRYeGQ3IWevjNZKOA7BbPFdQ8OG8gO4kP3Io=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10080), data_block
R+cxwQJJRkYJaTHlMrybbYe78WD/QUKNqlklB4C2GLravoRRE+vojAKksHgnO09C
/dsJGr9AMz608GpZp6YslI6OUJ0ShzJLVZ+y7cdhnjvNvNwnukm+MkOLgvS14Z8M
4vgv8Yx4zpOoWiTiGK9WJWcEjK+7mOI3dFfYGw5dv5ha64djYn/EMtmajTgVpuYC
geqjsufFuo19jVXv9GZDNk/tmTRUuNgHL3jVkmCd/qiYn81BZFN1Gp/4wyAR4av/
agZWOcdEhSiCLAgmj4WLd7HIC4GJKt8mllAg26JkZKZ80HNtpn09PBWdTfJlCSps
fYKKLmDSunQjamuoQvEIsfAl1SxezFHUyNow2rBwnKA1/kGDwN4nLbvwZqm2FWxq
aZuIurst7ps6NhvZvO+St1Ocf2aCQ6dc/xYQn1u+ue9S+5+ssno5qNHGcQCjU+lh
A1Rk8iV5vGCFzK3u9DNFTKcSLLeB5eF4UceBYE/K0CmOGYVaK+OPTNZoTIpR5kiE
JcwE96iT2co/wnwmRspOLOjTM/1SACnpNe1Q9JdF1XNMrZTpo0gVy03ByAcm6UMn
xUQDGKuKQsyMAHTV4NF1qLe430KpC6rIy7E5HIG7NqNVDNHEK6tOSI2J+FWECpSG
A2DKRvo7W6MLVPVbOBDUV+iEF1nTUl+ipJMsL/6gPPFotvczsaYuiVzffV7R5R8N
cwKPGbLB6wON6xep52Qauvkw7mm3UkVycyUVTHsnM6q4mLsRZ4On8TqZVAZmBs5K
uWDH75Nv63aThjGdGU4kZ208/XMh9htC6eahPSFuwIZVLhYyk+dt56pifWSC9z8c
RpQ67yR+t6NvidfkgiAUxJ0nuHU7tXPGZlv8nDD6EdG6RBQxgM5tHkknw/j+v2fe
mmlMqDB3T8ByUZim9mUNnlMtTUdAF3tLco6OE1KENsF+Mxuf180lSqziH/lTdT6d
ZEe9bdIqMeyEIULPj/me2a305pHu+VRRe7sMp3YxD84sBe3KQeBNdq+lPJHd+f9r
VQk2WNlIcqYwaOtt6WpV2k8QiaNnRtuZgi+gJGuWHFWJqJtZp9QbxrJkcd0Xjcbz
KGW8UVhbdzdvfEWzfMKvNNtjOxFAN3CQ0fAzjc1PvPZKXJqDOh8O33mMv/5xv3ts
N8lHXh2QMOJoS1t5ZGXlvmPHLZPnoFgID1knw6uRMJ0uYbOSPJE9PGpJypnhWrBT
+H8aPmVBmTL9cN1OKcU1KVdSxFj4L3HeCnZip5qesl4Bb/PmmmvGIZ4eUn/K+1Va
Se9Bbt690yyfAzwGO88HU0jYdySzgeUSSuezj3DVsayHjpERyrPYKetH3d1KT9E1
HADJjybTRPXnZbzY3uzQY8wSL2/g0b4/tsCWU5jqnbAemvBF/fASLowyF/R66iFv
UdV70vadnBuvTPZoxjqgQ7HEJ/wY9aCBLI5Qdmp3WqzX4UKh25zPg9F7t6IvKLxG
h76U0ctMCtM0aMWUuUHHyKLAcvZPdd4Xp/Dl6UY/P0ooqH2ZpRHWv0uaA6zhuCW5
j0xbxt/2XdXpiV3/WMMf5fktISYcuaO8arM2NJuBitHaKfxzhHFPJer7ecIHr+A4
lEwl6HO6AoN7Zfu/73/oDr8/F4Dd2/QDBPiKSRp69R2AcLy/NNn6fOadqB6PVwEC
8sjMMXNVVjTyaPvl9FGooOxybwZzUwRO48f+wjUfk/EC7PRkxEjlfoZL6sU0Qdiy
1V1lokv0i/p0MbJBFsNGbxsbJJrWCkOv3PMh7SWjw45+xw4ugZqwUYIQDxHbB3RH
OB42EcHoUY2/6o7k1WaDwYnGfd9LYKTMmTdDTqkg75uPiiz6xSLqoAc8CURLP8Sp
d51/DBlOAT497kN+6biK6KvHU1g81GVh3dareNph46tQsAvJiDfWzKODYF7mzpbX
HDkXtFJdXgufSkevILQerkQblRYqSp9m1WNJAZqypO0g9ykd0av/WqglT+JYtXG8
44kOl/I6ljC0CK8sKjk1M/M/APvdOkUZn+SDBH7criDscy4rsi6Aj5OzNTZoayyM
3lQhPMSvHrUllTs7wg2MtIGsY2idQIKtOzpKtk4PhdSz3e5ZjLUhX9AhKP+NO5cA
dlkyAfmcE+b0ApfnrCrhxR/XGhz2yKxAJ7wp5EMcQ8E2q0RRrgdboe6wMQUmif2m
miEFH64SI4cXAmeHUv1M73Pu3TzkSAyGy7FmTS/md+OQbnWAxKBfKFUbU7lkCzZ0
vhbebBwChCIHotDP766CdtCnx5tWEqLXigBOiX/UpRgPIQpoc4vt/tZR+6aCfqxn
2d5lxNHb1gqyAvL03tBFzGLbfo1OIAP+MOwT15sPV3MMyW8WjFxXHdFsa6OXZ5kq
GJvJWHyfznT76KVwESLHYmNVm8krXnrXYiE5jDx9uEt0abWQZZsrTSqwk3JU2Dy8
hLBQiGO3KA+nt/PSK+6SSr46Ljs9J2y3odCsFbK5zpY84Ran31EiHH/usd1m8mNO
4wo2cIcNbY8GBt8NLp1YrHhHC9JCOdUWTa+1n6GKXG6QdQWifur3V1Vz4OpbfaLh
N89MUTPD9vjg/oqTgIO0czt97IuUZqgIKtsVNvQ8ViLrKYfunuC0wQBoeYBb8dwu
MCzOYOAKEa+rJ9o4GejmAFil7J1vT0vuQrfzRD+x8srvrfCmDI3VY2UyRmwt9ZVv
D+5tcLhHXRHYE9TX4/HSm7No6EfBqvl1Nv+sT9HkokbzrOSrlvuVTm8xnAghSo+O
yLyhvnejFPQXSW9y36RnbVxHQDl2YLaid4QqdL9v3WrIgWGwptDRC1l8XkSHlAYM
ppEwUYjTpGMzeRltAIqNwUaFQH7NjAv8fPSuk7R+tFj82Civ6V7WgcaQ6Sn8srDa
cn9UFH5GO/+8VXTThg32N7OUFFbg2ovaS2cHL9jelKPsyljN9LvatArx1YsnvLfz
AGPD63wio3j3OPG7ZeVQ0nRcbNDi2RfGhBhOuHk+5TyRhyL+dx4Z/oWEJS8Yhu4U
2QRCpB4GXWR+pIxS9BcBn1wG+hSL9j+O1pUluyM+do1cxKP0VaSHq/yehwP1mk4g
e9yb6IO8ZJGiIaUAuw6O3QRI7fopLtvsyuIJs88Cm+XCOZdondGhNjidI8EdymSw
zKs0ChoFEQYcHKmF/ToR+WtsRA51Z/epMv7IxPV+e0quvulUFDQCEwknzaMF2cEU
WB5XfZJCI2U0+71GUT+HgGvNa0e8dWtVhb6a8xZ7Tt5tTJUzucFKFxjbvDELa1xZ
ItMNb70TbYjygMBuBhgjWwJp0w+fjJjKb2dHLAzN84rGhtXLzaweI7eTA7QIdxTF
j4oSX90wBd+bgz59m+URq6vOpNaivMrcm4OrvgkVmn5B7tvjwtcTUZWjDwfyv5Iq
GRM4WTSEb4Tcm1eWPYRBgkaELTugsAT2gwp3XAq9zHhdYbPneUEp7DLY3tl9U0R4
04BTJLg3QmOZ6+kXOJXsoinirJyCFq9Eh0go/wqdFxp7CbinZ+uEeWtWva45Wtz1
Z+Jl4PIsO+B455dINeLIa9wiXQrxMrtAq1MGtNuGeXaZ0R1KCalF89aAcVKXtho7
4ZfChbYnm9y2M0hI0W4oL9C+GpJegiNLTFHRwTRjwve5lraYGTxPfQyVwM1L8Z12
xLOeLU7j5WXW9Z9S6FZREQINbgdxB4cyQPsreV2azjYf1PMg3k4bOrra42mqlDEE
FSXEDi/o6UKEH2po/cTVq5rM8LOFpoNYiXkAIjy0IOke45JaSHIsRMA+64StzHaV
F8//ILkxr6Xo7SheQd7WFULp237RkXoc1tP3F5I1jATgIsFk0X+VJK2fWelP6o+z
kgIv0w4E34sndtNqhgV14ap+ktr3kaCUxaPhfAO9yhcxASLME7ig66/bGsVnsyvb
Se4vhAfU8jXbV5nfkPS4qf8db4VuIPYXIvwTAAvQBr1epDxPeMbc34FKJ1vUpARM
k2FeavKtMq2INuVMYLXjFmlc0JAzGnKFGC7+IGJp1V5eU3lvW487gErhnrxMCjX0
Yc3xEdmTBOn7HnYkj63wvRdkFxpg/fOC5cyeunuFz0vazy05McgsAdk58sbqWQSi
Qvp3FpyAyGh83WKiin/Lgy2psVw2wPb1cq6Qe+ot+dE9QPr2Z2+a03ZjjmZDXad+
pBylSC0qAuE4iGIrqUQUFH0VYSRe7UZ2EQduxffjlJRrmYz1uGtHGMfDiXoaftrY
0w99SN4hgYqH4Q0CYmOTXd0bc+lTFJGf0i6uIuQcJSGSueWv1RVrYUZ62EAnMc4d
5TXhEzg1Gl+V3M3Fcz7jk5zHKuoM5voBIL6rfpr565cBz4LL/cFFnWfvtxMMe6JQ
7oZNAg/RWq9WA6Paz/J+sp4AEONL9xvlnMEw1HNSF76VBR2JZdj1qJDVy48ZiQdM
8hHR3x5tzIZhh4TI/Ncaeu4Do/3ST2ejxMru8yjigc+4QaYoMGSdtDK3lA3ebEJ7
fGZYGMkK0zn3qBULf3V0Ddtt0XfHYTl5XfZdQnnyHYx3EYKnAmPTJ1a0r0y8zpjA
L2CrI0xttzSXqtq6h4LBhwywEluFRYKgxdSkMLkHlhuHhFmFjP71WyFIN+8KxKD5
lQXOuE15/5SMZxNBNlvukNyj+obrTBRiEn54tvoOLl8d6RofVvGqYRqiUsFkJaJa
2/KTLMRsXpib3mOPSkk1K0h3b3loDGqfJHjprZiGTMuSYOiE5aHZs+IM9OLcmhXN
HdcY1VNhQhaEfHPSzzeA613sWHl3CkJRjwTZwXLf193er34kayyEPZQmniClovQt
86GdS3RPrageuX3lG3ziQT0fQd6kKKjwhjKoFSQYsW/vN6RU3QSTrpFJJcyb6Pwe
0BKyL0xfcFXI/QVmzxGB3NFIMYkyKFJhujjAcSEmNFtj3Wa4bnhQGEPrST9nW3EH
62L2TLp7uz1LU6VGX1ghy8NU03WWSStbCiZCl3mTeyDV8UXRkNBg96IqLDnw3Scp
h3/41+h+xY0SDyqaECLImpCeK1+cafIPu+7H5ObdRlTvpOudpCn76+h3GB7kGAIl
Wj8FNejMdbvuoq3eIdVAQyau6vVmN9XyOoAQISG/FevBhR9lGaw6VlRzkq3zUmHG
Z+TluLek2/0hHJJaQMDAYUs1nAPJCSKoms9AvU9cDdti9tE0CmN9wdxq/TFY0Axd
ExxLyDkL6ywGt8RPSatNqT6GxP985rUpz6gataFxuc/G0+MAjY7A6r0aBRKSkC0l
eQN0/em7Mm6cFnjbTpVu5+BiLD3a8R/XJoLAYOPioQHf6ccO/Nk1Fr3Z/JAcsJXa
tC8TrPGtOtTX3nVXxmfchtC0i+mh+/YfoKM3zEo9OHTaH/I2BDFF3y65Y5Av1l08
klipOuUFzCHlP24cU21dryoKA6JaiWOwgbu/PcAgVy3XT0SmiK5bgX1trNjgsk2Y
XQ6z92yOtgwKIMkhOTK6bOdDPaTXMwZw5PPCkvH6Z2hKpXMyqoBU+4tT8MZm38rn
Q/NbS2u4mdgegypFlZZnN7bBBtr8Tj4qg7popwlw9Vf9A8ngFBVSWCSGHwKVx1J8
0wCsWElpEsUvDI3Lr1SvlljWizRA5MOXNQJ6OdZ1ohQRluE5GVdiGKKedG4sXI6a
t77R7IphkfAryj1p2XNylsq0z73Uo+NLQBSVXTib3K1DwCw3A9xmGWvjV9lKAyO4
ZX787BCDvlhetKxUfJI+gpuMvkaz9jCTPnNeaA3LoUkoiQT67z9ctzs4+iR7pKA0
dwunAlCWHBa/hHBlbxXkdBIzs5Xa5Yc1odptCSiz5f5iHbkPFFJ71BADFoGV4yjw
azHYbSe9gvjadckK4sLqn0su4eX/G8RxBW3nJG4yhpjB8WMqnfGq9eQtTqbziU/a
lXTHl59siSboISiXH3mOEUMz98uCahhKe2jJH8+Z6uWlsooe0QD3OLXAyX0Xq2C1
495jlqwisa2fnBOq3ll3eZqHeTjwa207isFyQlvaiudMuTIMmPiloErdGhFnzKhG
tN+3YlRRsuAiYaq7dkw7KB8bp7aBPIYBgQr6HX5SuHkHd0mkNnCV462XYJKfdu3C
jZevszMbtceqInw4XrBLFuZytD7BWo8BsHo03CVZ7v02O+a5rOuosk61+I/TZWx0
lEbwbFPKCyfcAI2G26e4KJctqkrl8JHxENcZNmT6ZKbZP/UpsMbaT2tUZp5IR3iV
B9qSERYDdyC/PDXV78wVqhehJBvnwxtoRhAudNwdwaF9CPwYwlqN6sWDN0RzCLob
sso10PJRSVFKRAok6pumR3yYuOrwYEQaqAXGAUXJvUPxcEWjz0SyXvrpGJi4Xknf
/RB8pTXeS566S0WCjBJ1KlAuEFOLSTD2yI+Kxo0OIM4wZVAEG8+aAIRAFH/NHBDz
2msqBc2gumtdvMymxariz+5ducsnnOvvTYZJqFNtA8A9XQaCKMmJE2uSG4UbwQg5
jADt7aGrvTuto8cVlT4srbtttslWB9zzQisJ40JVSAgRCCLWtfQ3LxmGfx7Sjcfz
rZun9j1zDRemmgqL+LX62iFaRoMinGjM7+3ZSFRlxbgMtuRvaKQM/d3Kqw1RiBKs
EC2JuVoEc6bi+tZ92Yrn1IHhFm/Wi7UCB4DCGJ6K1JjgISIoT/WHx8uxtNwJT/hq
aB+dwkANdhD8+ZScwVcghayVNQq1i9Uf90zX+IfV1fjzx6xm4TC+by2jxeigati4
ENPRutYHONP67FZVUzHXFTj7XkkCf9NeoWzP81+nLCT0FVEoI0ZhdRG2CmSZp2Pv
gnvaAC1G66V54+HMTG4Pdj3Wli3ptU6OU02BdEqjzl8mmhwVRObNXHTaoYLrwT5Z
Azq6vGEY1Vwn7sejVJ+WRANn/AW1Lc8bDQUT9cYq8tKxavfoEP02w/u8YC2arlLA
E/76l+E091SvfhCNFzOWmuNylDT1ozxo6fm5eWhVc7GguI4hqRMbxf5ED1AVdBwO
MMmP4T8gaBWTNUtLxKImhCKDoZmcxOofNNuBYuY/0TuCEozrrLX0jfSkS+ZTT9aw
+armyWIy1qNMOhbKBvOXMku8s6M7zS5v7pzoq+H72NrrNoZqWqN25sGXnfUhl5S2
rOBpk6VIXSbebli4ER3QYXJ142aytFXUKuKHQXMZ872sKC/ZkKjlTXNGFdTZ15uq
5J4sfOKMSVFuWdPkruBuKKsYK8OH5UWE7uob+69bDHUVe2mxrE02tRExCo/tHlGd
0+R4XmvLrQTZKGoe5LM5qa/SR3gt8HpD0D3PxjGhkkp228p6NkCi0xJ2Wv2ytBpE
2FMnXZ+8qSMgEPCME2dXE4Z09iDmkmSxF4CWDiz3QJq4urUBQEFJH7JEUATM/xUf
i57Mw5iSjMvtSObEEOiIsqxULOQKumOOXf08JCyT8UTbxGFRQvZ1sE3JzlV6+NS6
VIWNeqWadqd0vNEXdK0eWwBRI3J5W4bBALzWUVL7QS1n9dqZsuZr61dIPjWEggoa
My3n0r3e+IAjZvRfaVLu1IUXRJfinKJU++ujNL2pCdydr1cvpftnLjTh2k0CndnG
bsTr6W/DlqJtxa01URKgwiTvNVQAUuelnuDmB4oQ4NIy0erYJYY41cAfMFBdnNRN
OAfdDx5mHd6k3M8cDOqlycFaCw6tZDu4JtO+sh4OtEHQ5qiV+ftFlLBw5wx/kI0S
EVzK20YmAlswVeT0mS8GoiShzypvPZitz3Y4kr95lnIlNkplybh0CzLySi/BrYPy
91atvVG+Pwy+rPkQcphStGn6vR7meu6yxaec35+WG0um5NERWmNlaisWaM2pQ/tD
vaz56ZsNXK5iMq98x1DFTJ+IEISftg0Zt3/pPRao+K4z9AOJY9KUrmGGUkg0h7S6
GHXB5QrPyLvaHuqX/fCQHGcEYWxVg2YB9I4rkRml3FpeztQnVlD2l9ehgzA3uEZp
gq0qWuCJCsXOUSfM7DNg5mYbs6mnLwca2AFGIU/gusM1yumplB1GUouQ26Uz4gFs
juGdXN7f/2h5gsS/PX6HTvG5zj115kh9OBdXvbTBUodm1CDL3n5I0oj0zcPdXUOU
3rDujDgwrwuP20x3/4YUHUJFoxfBxx8qMWwgIjxLyIFASK9zaqbMrCJZ1dzPI5Ue
TTM1sOvOX70cSnx/szSRV5xNt1Wn+r3zAUsUE3m52ctM/m0LnyH98o4BLlAMbtkk
Sb0qu90FcnXTvAv9wEb+fyTiNf0ByIsDehLEVOvvSVNc3qxfboP7ZszXv/CXERy5
GlhSBzc9UuXBm6FPrjN9/sfF+YHJB181Fk24IrA/zvX0IBxIPQn7xcQGZvYEYUCi
wdexZ3ja79Sy5icxIDYkXMmTPYAmoYh8NA/HajyrJTx/+4exgZtQ4QbWFAdjtJow
2tb7FBby6p/GiQJVIcxBcZk4h2/SjFbqe3YOoM/4Cimgasq7ocxNZVLKI2/lOIUk
fZ/NPEDCOfnUJzFA1XVN6CQgJUWNl+YYxyqiMeAqoyeyvnJuN9GVz18gzvCkqHpw
K+dWYs6cv/nqDZsCVSsaaErspvhI1tkIfdmvEtQV2dAk3wKa7y38It5EE/+xN0Le
xrB2lWEdmztiKJUwhfd5b5PF6cCkQx7XCgHVRLeCUBzXvOBR+wbl3xsqO+csMEWr
jBpmTie/F0imAXIVjjW4pKl3pCylpmOToY8xr965ZMcJAyFjaY7B0lKH1Gbogk3/
BPlMOSjHjl7nrtXsGeQT3FsKzYVzbSZG+e2YJLl6k3UiXC1JYt1zO3q+BMkcJGm/
rqQKlX2szGkR/wBj8+9pp725saseNsqsnKmtM34MxxAzsGoTQuh8bHpHPfksnHw7
xlmcVsh/wXZqPGnE2WFiHKG5xdM86zH6Zy403MpuwFb8+gR+Xfn/wMF/2o5IP81a
h7uWeSFAJDQuIcBpKFZPKx49KowiVhoqTUv6jcD8Kv7T8kpBXPboEr1gQ/wnTB2f
GkKffz4xIjjA6s/HMFHqrn7NbzFxLSSGuU26aKb3ZP7Djb+F48udNO1JlOkwCn+q
XuYuVLl6fJX712k6KHjAScXQHuMX1AhxIjfDCxWxThUYvZleap9bW7QTFw5nBWXc
d68sZRetXwhYUs8hWBfyA/kCRV+AvUC3v8cl9radN+5OxR6S5uwjS5jwCKO+LPKh
j/Li0KP3w3K/5+eqzF1Lo5ca6mBOnUIew1KWbZRV1S/HxenVAJtM/ysTULJ+5Z45
rmiyXn3anAjoBhUaE5eNNbvSmi8eVApbSeC9qvgGIUJrjSOB6udGP93ACpUOpnhQ
pXwmhyFdjKg0+rV9C3WytRNflrTIzH0WqfPyCTbT2+Sgiml8IYH4coWjP+uCxjc+
B2f0RafeSvA5Q1H+XrHH6ugFgbLqq0FFKe+LwKXo512dtSB9c35YhJr2FCaWZU97
3mRsQp59cosCRWiE5ZbZMQn8ywwU0UziH3dgF1Kchr4QxzQAPzGH/dDA5JlzxZmh
CWRWfhJ3A+k4g93iSc1hFsyHBpCDpqvwhhJIWT+TrVfNs8KIBM5t3uClEq5rAdse
dhaw4ECbNzNNHuQ6JsBOZt8zSxAndez0BYQY32z2p3K8qTeGlB0huVzAEXsMemhX
qKauu7BQLuNPgmz5iYa2PU/BlVY+rAwYWv2aB3O60aoRUCYoo5G2Y/Ox9jvy3txE
uGYRp4PSzQrJls4V7ozprrmQ5FftZm/Y72vv4jl3fViabiZDMrYsX87RyKv4oJDW
KQZlzS/3Uum+UTwAM6+xRezeOTMlOU77GsYIF+pLHhWa2aupRvnmlAAy8cvCNg6z
UAjbRR8ExAnUSS1kSfa6PCKXfGblhUSAlIYgGR+Q6EV1p486CwjwUatFQ4roKHWc
DVNUowcClg5nzkArIFbu2IBb+Tl2TCsrrUzF904X9qRM63id9URu5rO43tBxd/EH
VbafUqbfeP5O5L4s1Wg9JwxqgGiPnZCMPR1hlV8J5SQAsPhtOdvM0NDBccDfhL25
ZGyYeOsAtGvDTclwMJ9hQNffIl12W6ceSYYq3jK+iAbNBuUw6iHCcr8Ce12Ptt2d
Mg/UYMQAL7FK0m0oSU7e4AkyYJ1C8zBs3h4dSw/yn9MWr3jRVga48j39c0EOPgAj
setrJGAavtpQpIyyTTn7AQHIK6HZlXBBa0ZmRSTAYQthEq0uXJoNR5/y/CcOdGrJ
ZUNH/SYjchzcArh/xecxYkAoM8xnhS4IHplyQhdxYKCEhDg9FA0xJNpUjeFNdyVQ
IK3MCgCEXrvBQRJ1sHyAGZBqyCOzZrKXZOr2PEDWVEOnzjdk5VEtMhWsgpkgReIy
0JBsLrABYDDN9hUv2YfzvhfSSA89xpsfSJ59DSgSvSaPkBRGpBF2KcylgKbPM9/n
itJQgC+I8b2xOczPtRX2iRbhgfO8OP5bx5T/Na/aW2UdBwZ+7Fl84qZQPc+aEnsJ
DgorflHTHxUbMnQONjHXgjmGLi7EvAFcEovP0EVSh0yzoMjhcSeQsAa68CPq8FHv
4vxltBZgl5gd6uASJHi5z5mFlhvYTCV5BPgWHvI7Wwemx3Lq/nZmRFtKD/qL87oE
IF/xRfCl/Z+l1WTj9+AD9XaOhIPnYxr1c/ru1H5OiTGJMA52E/fyKdQJxQZ5xI+4
2Hya5fIf2JwrEG00QaCl2ht4N5hZXNdj1p2cm7H0Ke8cC2jzDBizkY8PmqNn6dOR
EQbDmOrmgamFw2RrqTrkbvrBUheKXCeAk/2WS4mKl6Llv90Zwoi98TmMWVT4uW7M
TOGhSqzMhLNl94mmzlqurLbSl8/AusPZlbaKRa/MOmOAI7W3FnGRxJVO3PecC40T
Qxa6guEWMqDrHxfNToJoCBMmCj0wYRgQbwgqYkx8YpIolP7ri1p/B4iBjI4jdIz3
VpExFbxUTbmKBjywetpfN5A91DJ+fSdLcZqDg1NwSZhJWEnsjqHdZC8tA3kQHQYe
3O3ScOWe1ViNf+sdIHXyPldfQxpADF4TjdSxiMWKjC0DTMQ/71mnzB3mROT4Me55
/qgmzErc0kZ+Dzl38m6v6IS6PDlYGTaeHtD5QYiB/5PFPKaVU03T0j9EYqGo/c2t
gA1fk8Nw4lARHbuyfE7Rt+X+psQiC6RwmpqZrDTVoCho9v7SmsTy4vrYIUGh4Jyg
w7j915+Zr/0qXcXZoT6C1JP9IMpKVy5Sxqx8hp4Mtpzw8FwbiWoKipJ/VRJ3OcZW
y4YnY6VqAEP2N00JZ2xOsmnIye2tDxqonPLyRUrfIePijSEqIIsCQXbhE5GXAr9c
qeJVsxgyved8e0f+DAh4jAkRHVTkeL8ks+Ts6deHWmdEEO9JRqLV6jYxoYhNCyMC
66wB0q1wJoXhgWT+L/C22xNzIHNUKNySbOp8a1WkOW7paOlQD1KioUyUqeopUVku
nWKWiqwByJcmxrCszxI51IDViz1nTY6Ufg6B2QVrOq3xv4zuXZPYw/SZdMLQeGQx
QbO4j0YFE1+QjhSRrAWlMPmkFVVqFEEspKOm1JqXhGrF5MTrzvYYCkFCigGKmWa8
s1JSnJ5sddFtqnJLKoPt6GWcHuDXyWyhoZUS/VpdSNIRVv7EpWppg2nNwo/NBnit
meJQ2f2Z/yJ/aAQ2sGe1kvz3vJf6scGLYyPe7G5Bif0Lo7Iq2zGEFmmkNE1XDHgc
kdWPFLmiOaLlS24rvhGkIKSIsWl9UGN2rmLDnpWc4lnONKL0REzKkNwVzX50XbE3
OkWl5S+0Lt/uLX+98eFT8gjnaJbtB2KdgMgynSuDPQejpX5XqxOxu0+AOpFw5Z7z
VdsPWR61RkIeDG+J88G7kFQKYZLsiHrlLp/a4LK2eVXVKLi57o06+wstTBg5ZfZ6
xh0pEeUmBcf7qUgg29xI0sSRNRQmMegcTNMWR7q9L9f7S5SElxWzzTTNzbKJfwQ6
NZMmXVJoAa4rMfSEKLH6uxoCTosdrT284Qox1/OvtT07ckoMUn5zVrn9RSJQ7qTa
Luqo5Rf8R8wEDP4ASO1wE5dUpvAghk5h4fskBgL4VwDoUZtNwwxj5/TnhQ4UYoe5
whDbv+jIosD7aU64sinDS6kHDO9IjXZ493On9GFZgmyKZ0xlRHcANPfhocHE8ZJ0
DOieU8fK8/PkX1sD/lgmuQarEtRA55aWcwr+HtF/UFVkaLO25JClYSQHvypO6REQ
72jSWol9eb0Ux5CmIA0qMfIx38ctLIndwKLxtgVPg6avCE4vuxr0EjDRzT4Ar+h8
4hrrJUJ00Uctgj6FSLrT0Ibb1/nDSx3Ux1Wo7EdeABLz0TIOMWbvouISDTa5HHtP
uCaj5kyzHi8jSvyMlQ6qigbFFU1CtiNKl3GVHbSW3Sxh2MQZQgioCEj1X91Y1L98
9SqpTov4JRcoghihc6kaE78aBgBXGpvsuKObedg3Z7hwAimLocbjBYdUcsQT9OoN
xXrt02PXGtHOAaeGfrfLhKg3X0dYmD+bxLqUaV/MaLfIgrarh4XkHIjjNjbLToQl
hwJ77ehvaLg7ZeIm+uqwjijW1cG3zRW4Hu2g6oxe+vvjmQq3rasjDyNp0j+B3O+3
CmW6zNj5qb/oIOuv3zAsycG3kBPI8slMc2CQDjSxHIzcTNK7wu9GuL/9mMDGvXtV
kwRxwnODLG5xFC7//kTEk6CY7aOI3Teq1Tda4o0/bW9aguDsGf0YDmoiqSgYa+SD
U9JvI/WMdHxPlltzedlde3DtW58/zcf5KS8pY88tj3V9lX2E3rF7jLTWAZLnv1pb
IIKVbSbw82eRSMuyQZzSDWtsJcU1hH97s9dBv8YKnRsnygZ7gcJjqgC4AkihnQSi
1ALjwsMd8X3OJ8h1Og/mBN9nHwMwQx3YSs1X0ctJGE+7wCQR5KintB2eblrY3i4n
8IxcICeP3N0sYC6/+JnNZeSt+bvoNbL8jkAHQSdKebmT4Zf4rAYanMDXqPJ7PefJ
okgXByrITZHvbrlWtZK7JdwR9TohS8fijdH404vxyHAWVm3/5xNv72o+S5FT3A1I
IxscIp8MqHj/70EHSEkoMUEaxKw6EDflZGcO7z2n4308WX2BKdgbnxFEjMtG7aec
akOjjoyZadN4jNX9bVQLtlBjPADweZ0G8cN5IFFBcHLlli9oM3xKeKbFGMUzCJI9
FePeyMPiNlUFo1mOFiJ4HMqI4o2I0otdJhZbnKdRLayM8Nx8DuVYEpSRKLHycK36
XNrOTC+F3K3dgeI5nsnrzXSzQdmGKokx4ShDaGUn3qjTt25q4YolfT+9s7q5MHUL
Bt1ZV/AOO7GkHiZlhTNDELcyZPLHbfP7+ACxzwAuQ7hABlUngYSbpvNbR1Q1UGFM
OWi451lOZ7EXm5HGjdIYPyG/r38FNNy4JklHn30utJnj4LEPN1bxZmkLyHhMopUM
03Ej/UJ6P9Rq1BDm6J4i4olmpePlRCtZL/trIjxkqkcxEJ0POaLKIzhG+G8UOPhK
`pragma protect end_protected
