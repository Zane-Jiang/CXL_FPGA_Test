// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
WLl1VPfpZrlG0hO2oNmD8UeyB3rQCEGwjjEFOM112QkFJH+lyT9qvUf5OxFN1YpA
xnpTS0x4g8GBgq+7ZGZvpW4rrkc4qPC/0vIpR0LwHxkNUbYeZsjW5BoRNjuudBHk
FdhB2vPJ6Uml4KNjBGCXkSPYvSwb1XOLt3thHQSN52q9lwCDUljJwg==
//pragma protect end_key_block
//pragma protect digest_block
6EatfkJ66LUZThDldv8arZwtOVk=
//pragma protect end_digest_block
//pragma protect data_block
16SqZ9dTsqsQxx9DTOZ5ba+rbZ7tSXCXRjZnD7QZMpV7IIpsIl86obQXFjPvDIR4
mxAIykoKvdNLL9KGTqfuMEz363x1c0DFD45gKnbihSOaE1vFN0U8QEASxEXR7OJs
3MD1jlsy5f0jr88ru+k/VDuO9yQunjUSm767KSdecC4al04nXqxgAvG4WLhTeYqI
BzczEGKFmTM5lBliEvl8kQzcRydTbUVArj2dsqkZPg8QskSFf699UhZz1MQqEPik
jLN2O2/Xvj1YzCgqiKWSTONqpQbOSqBhPHzeq6DnnvoexzPsIC9ZsnPuIzsajE4P
waWW7TZXlhDytIonBslBgvABQ0LLY8qT0kdC/+yfXVEGBhCBctWyBdCh1oy/HcgA
poFOOdAQ8bbjxbzVOp9EK5NsvLelYhnWGj1KtRYGzW1uYt5Kh//3RZ+zgHch51dR
TaGqsYYMmNuWPvwouev7stLFXQsqDjNw1ThfV0V2Mf4yfuu1CkXa8RohJfJfgioH
7SW5uYQjLkYWMPV8H8aH1ocL4cWtNErXerQFNFA3uqoXxmAo9eZ9S7A/nLcMKVHu
1F36PJhxq+wGuacG2ktHWGk0VKIi1lt/52rx1XpZ1qJLaTD9s9/rTjZ33chOW1km
BsF6fh1SZ74LJL9PvbKvtnAlvBNuvKSBkMbYnYJEppFXLfmUgFY+PzvEvZ0EPHHg
iq1LCi1J4kI0mxgWgtPXQLrFO0RNEtO3aAIxdYkQBb909uzSQTjvzpiXrFgba4ld
Lo9/EAhcUJyMM2yUioBLCmS2YO9qYJl6BNp/6b+6ONd8uIjBBDTztAhwlHmcT4S7
kklmJtrd1QFW0tpgP4CgFD7Tgdbr6C95qeySBa7H/h6NMvU6AC3mrM+dJz0rD+RH
ivrOPXiu4cQsFbm65qCiCl6IqadWRXK5tFW7XNRRWZEoZCVnsPGqjIp2vULKNOCB
mj36KaoP2wT/eL8CzJDV1CbjliG//FfhAK0WHGBc+//I9c2abNggEYfosZgRCdi6
rzE9u2mrSZUQJJfpTL7JLuuLx5P0mpYyyYULAXsx8TAFINWf7uuQMSEqMde0AdH1
oWF9yHA4RFZksxGj8qO728vJP13yQtts4WfOVKKWnDAPr3t7+t5RqXHeSw+hL+1u
DGj4oOi1RF8Lap6BH9688IJZS0gp3yqeQQVomW74js11sCYLHJcDc8Wx8WizObFe
offy/+pLa/xAlJTkdY88M7q6726vTERJgTLjdcvOXy2VEf7M2ZIeOV2Wi+yTQ1Kz
3o3nvQn7tm6Y+YNVmQP7GJyZwfl5yfXlr4dNZXliueoEdV2rM7IVyNNmi7u2jCHs
LZAodvmO4z8pgydpG7BW7AJ4PMv3vYhG0XDnXhUo0DfN3+/i4PbSzROxVHvB/1cI
mUBoqy7MOYLDDRyuqWlT9UDl88pgcYfmAswZ+8OsrYTVqGYLV3M/yq9M/DprGqIo
q0lSoSw1jWjilH959KB9aUgEKcySIdnUuAx090gNJcadhrBJU/cBIKr/n441AITg
tiEpeIL2eOvBxjPjsBZSVhUfJYu6QTiabObgmWurJYQjB14XDW8dY6Yd+iS4nac8
PpEFvSX20FCV2djjDLxbgvzKNAdhqRoc82Dn1xgH6TAxKxpEMd7Ps8vEpfE3WIIj
niYfnXChOdERAZ+DgFtujr/m1Cq9yZDn4hAIQJ6etZTo6GEkh+1qDw94nGEYyqeu
T0BfQSX51aX4gDc9HE/xbgjCAmGBL3laqQQM/6W9QpxTkBMPLsrun/tinvFGjXXU
3WyCy4TW4ZBBZhLDpxvywGxLztBCaxuP33FN7jyBNooxQd70iqOxTfLGvuHcJNav
pDPP0Gf2GPqpq16m5vBy49dD2ubZ40wsj7QvoiVsmFzXdPvsJ1PsFpyp1hyCo7mL
g6o6Mv7QR8wEdhJ6wJciATsr87WHYcKVZPT5Hl6Hgq+d7/8qIhCQ5lRrFYepiXU/
DBAN1zRRREo9aGumN6sIY+isEZnCJIFaNYlpfFpnJf2FN3/ohKXvWhjhkbHYjDO3
Xp4r1Wd69kYq5SPUwyMYWF0Amj+Oknjn8zn5KmfyY4tHOJFEkNFRxexJhY305Ilz
wVpFqJYuoteH/4AZ5EpOmEGPQeAaFRjDfvJXjed0eIB0KZmKJ+OSzB4s1/Y81bgI
LOeOic5gD1bFjzZB1VPIvW8Trr+yq32l2a0AUwwiV9M3bUGZ10oNSCytpJecY4yF
1GKqOj6oHZBHp2NJE8MrwqA26B4lUKX6NjOJlr+z/ueeuYQjamjKj/KEVKdhFCpW
KhWAJyhHs5lwOPZR/2eRwUJ+LQ/Qzvw0gjiYj72un1+ed30YGr9YdfgHV7NalfEJ
C7uMW1gcNOQqNnP2O5ZYGjv6pGfxZw1DKH1EIRO6yKeZjOqYSIJptlorbeCawZJc
BEc1XyCMQyzrTc9EmQOvILiv/Qtcw389Igdy6vt8EtZZ191D0a/wMB1HkZdv1GwH
GYREvseX+n8H0N7HmhgmaIGW1FADjmkoK1vbS/Rf9jqd0IHCrg42pK7KIM5MFCn6
apgNyO44MVZ8DMW9yMUqFb3OvxLFXYh3GkA4/XJHvajVgSutLpn3UUdg92i2UnRM
GXyY69yMFBN8yIkZW23ud4UunwMohPKqHNL0MN7gU6MvM8Vb56uS3dW7TFIM3wJb
KWYvdYV3ogoN6al5r5UEBw7nFTeYbUXp9la5RG4OAsrE2pmXR795j/5hUELcY+Du
XLMDyh6iP99mpNsincR+9GTO7yW7C9s0dGBai7WTnAI0AAf5XwnfiBWm+jf6Mo09
YfPwSTPjH+UjLlyZoKY5gGZ+VP1xq9W/q6i+taPWUNpJe559kmhs/jf28dWS4n91
BDToktBu520sHInAJy6LoJWdVxXWO8B9yCJobfqTVd2V049KaRkV27rHjlSoQC7l
WJvq2IOWrjCm++qi/LpZIFP1ujdFovMZfpfbc5yzfisFJtzA25YRg3QUT80x47G1
q3OMn1iqZASaBPx6x5Ffzhsvkq3on00yjRtxmdJWt9ceZI8w/T/GZIJi87wvb+SF
qgH3VQnAFljJ9zc7MsmszbbqZZojjEjPAncW/DZPVEizXiXgeUwmGQLrVzmBq2HR
QDfA2sHuF1r1n9v6z3G4uvyhQFCuPmP/0V/UfxM1XBf+aG7O9NytzOy05EAi+sd3
0fuz4G0exp1l+l2InYYqsxYjm64UhbLgYDo0kRvzgKLkDcUQZoKO2VY8nD4KQ8mK
mHpw5yLvOwUUYHvIqnBwt1UA6ZknKRyF1e59hljKlXMq1ncLArGFZKoJ8HF49BLg
NS7SBIOiyvODWm9EcMA+UkIs43CeYB8ajnMv0rmb/5LwXbVEtfotlrLZ04ABbmN1
DAZtNe5q6UKTuetikBikbsw8waebpNYMqyvFcdL4fByvAEi5p4IZ0lItyomVl8xY
JurYf2xwbLk5nfJipa7QO6EszqZhJjiPVa74jzXHZBZLKI96FHNUK1R67vqwP3ws
H4wcNgNd5E5VkwbJz0/NiMlkt6nPv7/6fIiEbpOW8/3mjjPGDWHaSki91r0gbxea
ReSNU7G8jqPt8wC3BIbd7PQXYhCwnVZfPligplULqekBQTzrxTT9pCIRBssXgUgg
tMsrUV0HKPc9U2PBDPaI9wL/oGisUZgq6I7415lWt8IDsEy5CkuwpU7EZPiFlR0v
W4JsX4f0QBfaCWltJEvMSUjGy/PjfPERRFBHEjNkC7fwdy20I2FF5RIke3tYW8KU
Z4/S5Py0NdwCe3SRpXlVcrR6nDUaE5NB406rubVpYjnbDcn11XBu8wAajEy/Chpj
XcYH86tiERodYDt9FRttmn/HXClEJ/mBIqnqWRUHHzxvp5opQ996Ma55BDv9RjGb
1Crg3ph5LFRBpU94hr7p012JJjtdIZAJu9emQEUjMJHsqQ5PSV9tb7SI3FRDLTWx
aYCRzH+xnmKhCNavc14rugYm3DQNa9/yj9zZNt69WT0tq/k3l8XveOLogJd/Mnl+
Rh5zGXWIMTZSGcYjk28YDg3lGvXO6xyRoK3FGP+vEg3EjIfmsPLOxjgFZnI57V/p
UdCEcVuOvRRGs79CBtdiHtDpUhsyPkRaxc0I4ilxPICpdxTCT/78Ish51sMbGkWO
MrVvu42lrcXEjUBirTTSniI3w0Bgu37i2cCddEA4qWig/vyzdPo84d+HGG7S/0yy
7YIoiSD2lPXzf555Pp75bhwk20V4zITDsBlp5GWg3YbOCy/UMtg6rB2D9oA7Z75R
PwoO3Tf54a6SBaRJiQxHojXGoIZIBYgb8Sr7J3a9GhDpRCX46dCT4+Yu+8RIVVsm
qZhFfVqyjjrtD+0J1JGRSvKrQsV7mm1qW8dur5ZaNOWdvMbxiLfdk6qIYUplCuF1
TDB0Y6CQO1oQzt6QuK26gJCytTF/7nyhihU57FYdNHhGrat02MeNwf/2o21U7Exd
c73ImjichEB3FJa8ly/SssX9SaWK/HHChiDneHX/WwoG4rufBipY6SW/53+jqh91
GImvXUUsN8FadCVfK80LD3BSNL2+oqsprFzXzcH1O1tyOJnGGIAUrlQLPf8zxdxA
bx3kvZV9f1jXiI2ybGgwEuxNupBIms5hkNZhXcMHi2sjxxqpSMZm/tcM8qqhD1Jj
m1rNh0BvKZ5WGXks6hyArEZTl5QbV07GQhlOvLWMdZcB0/WG0MA99pn5FqZwGG8j
ZVhgn5p9JIVkj7udTU8JCPSf2Bq3aEUcX9LcYoPyDu7xa14fJDJ4/YSU9JmuPuPy
3x22KIJFw0yJicbajCKkvujZ+jzqIOP19hXRRZ31lsQbdgwkLGdMcaaskk0xkA3P
O1M9DnMcuE8fMOnz3sDB5LkgyiJ/xThCTwJVXvlK2lRjAaQDlR6EpBcuymQL+VH3
nhwWAA1nRqreb4VJerJ5JwKuh60PDJiuIWYjXTCCXGEuNAlk4c9U0ty+UPdgbv/e
cOno5GnTzn3g+r/YWZfd8T+x5smB9Zfdu3LPMjhvTLnGrT2MWyer70nLJaMx3Mrc
CG7tRatLy1SPUT9+707fCvVSqg43Lw9ZGyjzszI0PXIw5SMpcl2y/rZZw/q67kHC
qsDkRjf9WBXMdovT2do9dhMvREH8WN4Ei43R4j/bUhZSWuIglBTF9Q7mTQzZqXlL
8diIyBoHGnvURadFjDa9byxQ5UavcTsxQHf1YxBSYlJ4nH54g3gFOO1jn9XZSX5d
lmPqiizeNVH2bJXIA29SIZyroy/ThBPhz+axp1IJwrQASV/uB0VN/PWMMGkcC90G
xa6PzN1wFk0ipsXlEj0lenh0ZGvrE7x5RuqhaXrU27oLEJrUNZHHOo6qdpUkTNAW
vjq/0mZFAxeAImyBXVI4Khi040TxdVXJ3zj4rrbP4va09FNgSmI7WUxlv26ZgHii
9PQJk20kkeHi4EjJo3bNF7gcxlelw9riJHaPydIhBLDUubTkv40Z2FrO5kId91UV
smNYMCRkM9G49fJXRDC0k11E9iP4911zbAs2/U4YFAyBnte1Ii9bd06GiV0Ar3p4
Bohmjdm6bvstFPs2XuUP5SQVMdoCGFoyXJv0rqHFtxIt8IhIv/tw2Q94NKfPv9V8
7wsMGWb8nT2m6THNa5NBPvLmUIpEeUV4eRF9FuKTIBKnbpJLtsnft8b5HWWePQou
aMBI2twicDn44LLlSj+8tgbfpdPzdcBpzFXDYtfJUgDBqKxYg7in+EGaDRJK2yH2
9GiM0zacDhv0GMqWPeXuRnA6Iwv29d/0H2K+S3FlQW+ir0LLlTUNAm5j05rK/jAe
hpBvddXY5MG0cy5ah9LS7otrc8JtiPu1QJUVIZgkqvNThgyyTAuTQBtnpVn8pXFo
4H/1QOkEm9UBjx7pZXnyqSyBiiY810/fBuF5WKJP9fSlSAnBsY89xUaGx9z+V1c7
TMt+sIrvhQHqYdbr4hw+5foq1/NuUKZa/fKyr21ciBiG0h05Kp3Ystn1U5T0Q17j
InSn720wjY8XlaG5z2Mloccg/hw2kndpplThyWUbKFkJR/F3vHwBLS3E6V+vUUrA
jBkwdeXgKNw1CbNmJKash0Ioscq9p4catcUWwz9mrQipyoKTXUd5qCTf7qR7ch+z
isL9jCok2zcGhEVTAANuky+PZcOHrm5VzfNmnNlPb+z6Wbw43NoXeDfuq2ZQs7VZ
WNtVlcAFS7+A0Dxenlxe2Jerdnqbo3hxDU4OpJ350xjlnsFvsa5HeaiLnnH+NhFe
H8x6+88PiPbsqAoK+wrRs1W8UjqZkjgMbRYRBt39eCpYLbiSDTil570/tblLeLPr
FLb2jgqtijR2RMw1MhxIkC1vMJcNu5WS7xPat6a/I8vwotKWEc//bikfm61M6P9/
R6UVepjdBIKZrbvPhaZC2iXxkh3w27MchkkddsNKciJX2grIxRUsnbkLJDtkmBBW
aC6J5OY19+0kvocQDhJqyr8QrirB8Pv7H5fAIvEM4beSFfn443WSEdsPGeHVKTZ2
2znFMMKUlJonWdHWdSN5rMhJd2npw0stuNhkfR/i5tBGOI5u31QaxmzHNUy0PLFo
8blztUvyFb4uvQ+C2XMAU3ScqUk7yOFl14PVM5y7mNdwC0w1RdnQ/jAKod1gtdGh
9gccdSV6ene96CEJI9g2jaSDKJP52BuuvjjXvSd5mf2820vetvXMgJBNx6clMYN8
pHvP5B2F1cXmM9iyxvaALhzzdxCroZQ8vOyaR+krPLdJtXxc+LpjZ7UDQlyiYfRC
GNwi6+F8jBhVb2AkoRC4xEL4088vj7i5WLaWdMtSZZjTcThlkQodiMHzBVl3AMxN
KRSrgjaQcZuDZzHmd9CrNbZ/clw0lcGgW6Das96dh8GuUitUDcMWtEH/O+LJuzin
Q+aAhTm3BCyMLOdFMiuGmouYp1YQYfIDw3phr1VPEM34ox3q48OVXp5Mt6+ZCeQ8
X6pzDdUiDdwFHwiU8RCeYMnKaOVH7OmclaCtIhwX5sq2Io+1Ec2DYs+Pn+jQVpKH
EhMKlsP0Y2Ast8Ve3SrkMGFIGFHgdVqDStsHbKTSxpbw7HZbgSzg8vM2X5dJdFC4
aSCNPFddiRuNUJGv/lSAR8en204xloCKPsc2M2dduPv5FEk+LNdCI0aRt2CdnDsT
QBNBofZDiH4e8qsZHaVAZvNRaFf6pN5GULZX2mFyzIKy+Ewh2S0JgAqGuPZ1imBf
jOf4/mYWmYEMOeKb9lNtLEpbqW5mYEtyKVuHNarBqGItT1kCr1ocrK4+IECYkfgm
OyJj91jMhVMiHQiTnVFiP/EvdRADO6D729nwmhgfPZYT/CVjzpWU8QBQj4ytkV3Y
fwMCmIkHL+hzX9YBjLutgfjQ6s3y/EAanPXuoHZcoWZJA0tw1EPW+zqvJnQQbmDw
73F2Ppaq8G4ZmP0Ldzv+q7Tb4x7+9BNydahU2CpuIoGLvs+Hmlc3TG3ofVT3+Z0y
kc7lrNo5T33RVrPsU4CMrNJaKI7oXe/MMRicd/F9YDecASnl1xq+y4dVboURziQO
HkH7BL4hvYMolqNs638BZjDgj9se8sCPtKpqctik2zRSDtxbYYYb2y6Fq1iYpXcx
l+ytPP0f6lP4ah7Ygg89KvDAPhTUe2dfJ4smhCXb2/pK5svxYJyY3rQqbXArtnnw
udKXWgBus1fKEIO7361PRisRl8z3eWF84sGH/kFSyuhoWdgcH2fx8p3Y8EJA7CuU
8QRKzCEhDDYY9zP5AGH/WA4BPyooydxqFSMujI7l86KH5u6zFgUKJ/fUxdX2FBBh
CtwWtIV70fXQIU70tn/Fk0nCz1V11snfD5Wwo2OJGZqYPEvI6xZrm66LgysNrQpq
DFxbd5BfYGT6NhyTjdx0zm+0VWJzr+FIe/kY/X2otavrJPz/2uBVv6h6W0suiwh1
HNKFnBcQlTDHmG7VR6t9aElVVRePkZ9qUO+ZPhPSyDMJnytUDtncKSdt1m5cqiwW
zRA3SwoKIiMvtMmtCWxtlUii91wTGxCxWfXrKsZJmJFLTUIhsMEdNCGPs5GZO/we
De4TSZe4SeX2B25RPGMM/MJPx7oZTDyZhYmny6v2TCRUFJEGNpriRybMRZAHuPuF
v8duP9XpRN9y0gzToWEUDlIjTtpJcJeHS8SJAvdGeB79pViKfkKWGuC5I905na4j
4fWxILtGziHtYGiJf376xdhvlm9pLE7wLsZhC1iKeATRcdj3dIo63qQkUXck9cer
/31y/jhwd+FR36K/Bz7zTRuFO9JvDmZ9wRDvIb16ZjWZqQuDuYXokFK/70rBO6OB
sH+nMx9RUn5hqCd+Ho4Txo19NjNQTLrbQdsAi2TzMalrVAT49GuqEWZdDStoVp/m
eEwyivaVCmbvWSAkQw93Ivloz3vTr0LP61IkXIAeb4WDYFFIgFe+GKIXAjYVELfC
0nrwswg97eg3VnoOZcKDA9EveJS3t+YfFh3E10HREHM73fG3m1Lze1gaWVfG0Pe0
F9xP4NulrvpYdKO4Ahlx0I46aem8zNdKtquIo7ZBH2jF68qWrvbndgD7SCbyN/zK
04fgOjJatVQUD24/OVJ0Qc5jrhe9x4EVcrdo4mwN6LxKXUywIlnmyLhkh95+fe3y
F+vNNgBZz7XSKqZzWHWYLbnq47weeTeUcRES1AeuD17BaAVtlALcStvlns1hEoTU
EsA5Kqt3Jj2pVkWRDiCvu6XXOA7On0HPtUqFjbQUkEkJszzj+CtMlYy4AlYpxHcK
FoRQI1qrVvSaoAgumURUau4zIJIcMMybYzVA0KgoNnMyRVYEeCJceOKyelXlLvgv
FyWKy8dLH6NZVRRIfIWnry5qOYFPiVXQdlqPxKNoB5SIqaJpRRSNtX4f8+wn4l4O
RyfdyHHQOiXi2dDrz7sg7GpMP6w3T+E61gNCKh1nTpx5MaflUT7i9TWNQGHCEEO8
cFqhXf2HiVjYbvnqBbacNvWGzZ3HHX5m311KZdp0ghfDyf3pJ1a3OWP0Yjsqhkgr
txoKUdYTC1pUAOBbOt3VXf6a249ZeqaCj6swl6Cxqtf2tpiYh80N90Xcdk7QJk07
ZjgssmNm5sDWkZed3DRB84p3iGz3aV9Kmenzt5HNc8SFpnB7b+bbnz6Mskwmr48y
PgXCzZnnemXayUFlly7uNflpkEKYyfaFHmF5RXgvs3gHQ7yXHhkLKJdFMJOsIgGs
WphAeJMz5txqmiuBiOhALSTUYHCPur8UwtmEL05VSQ667jIQUtZD7k+RVe3/FZdx
Wh20FDwhjF0/7GfAWOsOtfzQQlqskI91LD63c+MjPc4ZkjfIYjpLDAorrPJsv4Tf
JhuaC12Q7z5Xg+CdLHBD5xD8heuNu6L6sciK4pzvqL094ckd6ZaL6SsVhL6lxs3K
jK7YDKZH6Fnm75fOfdvTWBB6Zd9/j2V4aZeenJUxUJzz6AYkMIWytXk90fkZYt88
PVprAXOGP1TL+kxisnFwFQ==
//pragma protect end_data_block
//pragma protect digest_block
WO6CQxihBC++Pgy/W3ftzPET0YI=
//pragma protect end_digest_block
//pragma protect end_protected
