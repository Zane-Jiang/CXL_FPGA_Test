// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
TYjxlYqiFYOJ+Bkfai/zpVHCPFtlv4zZ4Sb3EvrIX6nD98tk3PgHb+ZoBPidAYFf
liIYSWdQhwI/WTlv1CaUivPwN+ZEboDRm/GYf1R0j7FVA1FCuNVGnprxodCdpKcr
8BYIMw06Sl7O9OuP2uU192EJjhGj4FjrUZNfxgExsEs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8464 )
`pragma protect data_block
sGqDlItZDgPP1JkBjbaht0IMQEWcAkvKnSihBq0D0bcoJJUFE4zN81Zwam9UQqkq
lldxR6Jjuqr6AQsq7F9x7Z1KhV625NHEkoUtS/wuZza+4hpZ8uMbaru1seTpbApa
gup9OhMsyIrpah9pLM+p+Rwyb0Ga4VJan/dYX93jAKqJcJRAyjw+Yg5RSd/YKZzs
sdY+3opQp/Aidl/lxgUnZjfj8fHVrp0SJJCgNWuYBL/tKDYF0riG4wMqC4PXyMF7
QSFzYE9yH019iDcEaXCFBHZELHu6fHcdVYKSqFxFIjm5DmYFLePFyjJwn309VeB+
+Wx8E9+mQ+dzSpVYYzZEBDJ8B13mlcMDFG79TLGsTEnAlLBedN/8Wbxpdgos8dRT
3v32NkgJobVgw/4qUjvYuzA9pBalXmPZLKvozduL0P+9IfdBb2co9KWMGcKtHH4O
+7VD2JHfHS57nr/Zhu5kATL/fJbIbxgRWR+jWaiivuTAPtzSHBvlMW/AkDjXiERC
/qh4gdNQd5516uncrMqUyZgwSVXp3dKx5xKgMLOyJDSb1Qf5RDclrw2N5/hsxlIF
aX6e0YSObm23AVX6Xgpnco6Jj1anuWf5UHLxAVbE5DDHuehqlaSvR206bN0h+byt
RCnF/YC9T7Arde0rpCGkF396EaJChkTkBBIouFDw7nG2Fk1D0wlNRNG2ktWZFVSN
e9OKJ9JzVAVkQlazEMAIFEgF182lESC9xcUAEYJq9li+Mil2PqUM2Eu3fS/O91r3
oR0b6rOCtt+8t4badeHgk/Co3CN/ZOIVFcZv6FzuafvBLLeLzE5Q4Ot/FSjSwTui
hFuslD//EUamHoMcQ0JWC0godEvR6d75T/W2/5j9u5+A6kMppfIshFIBWquYPUFS
aHhPRBS+cTMfeGQpKzAzA6Dae/LCUAvcQm05lkqRQbwsdf9Og5Cq0U+FLvyyqAw+
w14hjK1Dzg7Mci3fdTRe3b9InmRZqg745vBFcBezQk7MnwlD0EQXEvMSL6BZOxbc
dd1WQjcm3HePAz/AWt+b0dMbnhc66CU6OtUi35CmKdA8uHcF8HWm1iNxlw+ky3mN
N/0tT7d/soMjn+H32QndZCEeeRBtkjHxAvRi4DPHxjivdPXIQgEjM5H0qTVcHTpP
0FWqS2dwtCUxcF4gZGB0aIBk3JDuX0OBuVzm20hHGHc4wqxGMGPqCD3sX3K6hdE9
ighPKUzTE+4MbfkyS95KG/P3ukQV6ewXBBtG7T3wjfC+SA+QkxVB28EDv/lR8l+Q
Gs7LcdSCr1R/79DZSLRbi8Sl3yXRx1GvqFBhPzmsJJf+v0yOvJUhaCgmJQZsyJhr
cEMFQWLL125QZYOJPUhOiVNg8P/B+XzwHXtbMbT3KVNxpZ+J+VFE5caSVu5005Jn
QLRhrymr2l2Khd5sPMqPGZzVCB58OnncRovTnxbqAPbQB7Ahdq1c1m9dxR6Hrpiz
1zewVJqitszvhDr2MyfhYQvWGVh/Z9wkODABTd8ebEaZdf+/T/UIfG5YcasveE3B
KIfT5RkSz0wzYiTfJtHE5xmAI4dkyY/C1LJF2S44B00eSxgbm+QkD4AJeH9MXGNt
d1ZuAA8ycq7QBMlHqnd58KeLVmYRPLs7egTnkEGnh0+uXdiL1j0uinvA5bjkc9Cb
cSzcKZwYpSI/9LiFRXobX5jWdyEXTlQI/wLlI6m6bsye8Y4s7bc4eNK4hlorV2sO
b6nEoLKMJtSGIU3uugypp8ow9F1GHWy5yZIVyYikG0sm6uNfd/FoHCAulZ5Mcc9h
9ZtM7XokTA7kJ3gdiAvvVaHYqu0fbxE5TIsYR3W2p2vIQ967w/PbWR9y4BPRDnBq
Kg3L0jmdsQfc101wInoe344NMQ2tzWuJiLHV5F9Uqnsm6C2gvSbVRDwghPbhIRQY
7lRoozGQgvEuicbng6m5MZdjLwKfQ9sccfwG74jgA2YHuRbqzlqsdn+gqClv6lmS
Ho+pZmZvDHiapxfOoG6qVfbdOru2Bhu7SF4kIhOU3u2Nx4o4sf8q39ka0184CIlM
uQ0W6KfEtfRW1UnGuenBCwOWymvDunEXK9Eqt2HWPup96obtflPI9R4Yg0d7ThsJ
JlAVHfoJSL9e4ufqKR8zcpVlm1FYJkJallsXHrieEmm5wK3yTGrb18h7HYoD2Zcp
YC5AesdK+Umb3Z8Z5ttlGiHD+/h9UzUcCfkQRKHUIBRf4x39DPK5RcHbBdgCC5BH
BRWNcnI7a9GufZPSHyBe90yHOQXS/+9PDeJK7cIRtIffou1ILfTRr6kqzFa07yFS
cWYXPsOzA74NkYvxGdoxflYT6oxTMcZgiJFendsXEpRl8DjDN4kD5Cv4DkyOnXcz
1ixJ2VtMqCsVpiJARtoqitqswil8NLT822Ns3ijyE1wE0APgYeNi3n6OqRlv/1bl
ph4ewVZ1S/jmvkQFcNab/vGWa4yuq/lm+Q8JTQPmA2OuAJ/OIL97IFvVVFAiO2Fn
sRrrTOg8EG9MjT/niN/65/PJzn3I/COD4ZfcKoLD7LbBvyHh7XILWCZ4ElNJAyLy
61zzcA05HRqkubVzlly9kRk66iMH3zQoM4onIvC4dn5iChm2JeBGFFXpqK3F3E0K
VlNALvCIX97m+A7+jR23SY0zYp6Uwzt6B7HBqyLSKvcfsw+OsyQ6JY1xcJbbNAgi
tc85dDF5NTOLWW0y26QMh19Tk63L6ZLSVnUQQ1InjThXf9qGRfagmBsnRbrUtVxb
TIuAIEFHJaK1zLgBTof9u/TKrGJOS4LHOODdMYFf01+sXOdhb+XluKqIczE5JjqD
aLCx350ZB2AzxNmvesz31BY9kzEMvUdVRQ05cZY/XcrC2ejzGA4lrilMj17+OKrE
7RayK2aUaf39/YIcmuE8alO9A17CNskDwh8a6Z5Z1emnhc/kxSiYb09yBwN58BAd
L41w3Ga3OIAArdqxo87kR5G3PmG/dNbAF0+ttLp/qSQLGihIVfDk0Uc/pDxeDBAe
gagPPOSDAPmu0E+H55+oTHVcfv1v5YzTPda9w5bxigz1IBKagSfkbZR61dh4B98c
PlKmNCFbVPIXwngN1NE1AIXjrGGPbXOxFZSqfAfGczQB4GG0w6OZrklI58rXGI0R
n74knwt0YS9vUn8A3xBh+wNiqRdDm+a8pyL9JoPvSBQtgHd06hsUc0c8Pw5dl7fQ
mBSRtjmjmuKkBfU+atdN2WgUBqYRKeZRkZUwS9ngaePI42ngPgZePPa7FZ/j0Tg4
O+FoASH5G6q8fagx2vW4FQ4msagvvQGrkVQKnwh+3o5kuAfYZbdWETF4ZHjMLTZH
UIbUNObsPdLhy0N1Xsr49mAHEOjz2zu8f68+Ojrq2UCKhUJCWRxiKfLy0wTEr9RJ
dKYwvmN0PnUyHpXVYmjnfLToNHTDBtRwZJ0XmPr0stMFssKFleW5ah+PQJ8HYABE
SPmJuaxvQhHzhhzmmm1tEgyDUNFxWbQqtP5E/B20glM/osWH6hNrHevQhaD/hTpJ
76542wGrpo1HrkpyuUVJ77qyz4WU0rZlI2gvBO8+Uq6pHfWLpo+crUzuxbwE88Os
7UpK2KTnuTa6w7+IeqB51B2caXIaQHsF67WtiyhE728FHOiWX6eJglWHw3MHe3wg
/668dy9DCo4zl8IE/l3sD1CSR3eUHFKtU6vNvWminSkjCWYpvMC0J1VpI8CtytSW
1KRnAy8nyBlxhc47CNPFSXFbx0szNebijPUVBjqAAKix6CwYXBwFr/zbQMP3jw5h
wIWYAIWvjAG3yL9t7gppyMCRp3tHt+sQDG8PJF0FHZmdADA8/kQuOHyaPZMh/vSe
lPHbbuSEKHeX4WKC7WQ3o39cAuY9XINmAfuP9m8d+s6fi5Xt2cdAjAhuHyXfM12L
GA8unmuKF+6WmxvKocIIyVQyt2keWXCNuYyAY7kqrRjFmEpa4Clr2a6oHuPEgxSJ
W02JKNpZZvh3dOufnzsACutZc/C7vBO8UrfGwFwXoLAl4d4BBUbiL/6uLJYd0XxC
kotm9KBNmHDKaRYvoVpohrz7AAesxOSfYMU+oolQaHjKH719Hrp89cYHmlWdMY82
7QbihvZ1qqvViJ3r/wjwkl2O6WsYKpeTVEgZvbHcM5OGv/e3fSCPjXH4FpFaO5uI
1wPjSPtckhFNNi66wcH59A03c2BQI9IPHprruIfvexTc3y3bHhK7J3FzeVRfWwPZ
sJPEO7ENzU9u0Kh6O757yjagLBECwqs1HuuPPubOxT0Z+qPOXNwIdZFxN7OtsP4c
dex1UeRDWp45X2XZwUMtAID3WSmasmVtzH81Yz6h7fFp/vtj0wE1s9zPI1OAjTEb
kYbVby7FC5DNL0xBgwR4kJXAk+4kBYK/qTHaqazkhY9HjZOTWYA3OrjZZ+0C+iqT
YVGxqRHNprMOMxB8NBqaWrwi4Tw0/aae+OYYbynX66bKU+YQP1ZHpVAILrDYCAf3
jKheg9ZNo28zkEtOQ2zPaRE38XuO1vhRaiRwLSio66wicwZYJEW5xJi4WDHMeisz
396HzWPnNXBQteZNIPE5ZMQrYUMLyV4UFjQoobdfahnQxyeyvW9ddDjSI2zHnIqA
bAx2IYX/BODmsCKkbb7riQc30XkYJsdZTUyelng1NRhDZJSdHE/TCcARYwmmZYsy
mKoa36ila9j29i4r+FCVaBmRwev5QXjNPhpk85ywpGfwrHQBz3WVx0wOgm2OQOy9
586NyAfU73MvARILtZokQcRULF6DLgF8SMEfKtQLUE5ahQqHhfFi8Hb5mCDHbaPl
AqevZ4c10PgjrRr3WLGuiKgRXGWXpnP2JTvrKHJMMebrXX++9QQqeZsSOR8Rx07Z
5WQU0qgUUqmSQhm2uMrM7tcJO7VRxWiMPBdIyAoO+KemH9+fcgLVgsUC58YLyq7y
kt7Fj/Yif/RMDqPzUYQLvC5z/c0faV9Rs2kayKpZIj0xLDon3hmAetv8YuRGIAvp
tH7RivWq/PPT4y4OozQPIW3ZnBPcuCm87GO0uH6fhw+2lNyQ1IUxF3Rp5LYFgKP3
ADXTJAb7mgdYAKIw0j+AF98ToeOTT3lyxNran8op5yRP3An1SFJoExa4aykfVEhu
ioopTVRTHmQmsguT04zlXJcBVHI3bEYx1cZiAnWIr8+pv7TiSOLzYhVxNnuDJ/wb
57QXBU+CJxcicKj9UILxqieN/sMfg4m9FMKw6Y9I/MASysLjNYd1c8V05rPnTh3E
2/M4tNJuBOHz7OUCZFkmOfR4YiBVr6AzAth6LZEHn8cRk8SZ4uxHh5txholWzSQb
Jxt5cysstxs7D7TGn0vkCHWD/cjGIvLSGOsjyArayxL2L53J89hpaaMhtZoaPH1A
Lk+Hj3PGpFCh/W7dNEEeVLZImJjZp+54+rBX23bpciWfc3eMJF84jp77an9iWs+D
+iufjX08ge/DBqHj2Z6Rebr6nJvnYgE+uDL8xae05AP2ekdxk7SppUklrhsrnw/X
J4LJ5wtT8kJj5FU1mh3Ci3YG7/2cV35rzEpEIPDfY2whWrrjUy36zd1VFwBSdETe
1Jc37KkdzizNX7fdvC3n7oQwTnZ7VvCa4JCCbb4sSKe4XjRAfLnJGM7SW/fYa+nk
lUNyQx1BIGWjlL0BrCwKWgT35yEev8JkpD7OqLQ0GcRlRWqsHa3+PyX/6zDAxKTE
NjrpT86TqOD1yUDDiniXIGxgVEJn78jrOOOEUKEMDNxFZNBUqlkc1R5PivBPRnVP
JQPInG6WbX3nrBBGliQv9ZvOR+mut3xFtx6ezViftGoIaer35yIHAxMCLTkIH5eR
+apXZrUE5aPXWX6GHQNeWo0/YpqKphVtmyB7O/p6CroFMJnkMfQ6lrWFV+v9Uwzc
VbVk/s82kKJYw/I4hMbz1ir6TusH2m8Nvn52PviyGHGmpDND8RsAuUkZ8ZMNO6pO
H24BqHIrHW2exr1Sju1lzLSRNjOkiXTsP3z6YLJLy4Hx7ipR6+nju9uGf/UTYTew
V99YEB5bvzungYlGK7xEI8to11sX6rR/jWuVXVonDGGlRXrWbqyj/9seaYW8MluF
luUVPA8XNGGNviNyDxFYbj5dq48K6Xga0sKxiLm7QLJ455Rzb6xh8Jdw9+iDliR/
jtNQUFbFuKrVonIHPMM/+amgVXj0EEQ2rHsyl8ZxrltWs1at5+ER3c0RiOmHbsOU
4IQ7w6HKMdNT268BDkFcLnvhjz56B4wqKNP1yeGu7GIXInvqrsMuXB208fNd9FKZ
EPnLFXMpa/mkYrrw2rRuf27LzSStPMVYfAdl0AKKwa6OHyJ4FroLQXGLuKFeY10i
CTrYHdY3qlETESyEGt9k5ZjVDb5w22qAzPEhpu+PSgDfpmbOuvJRdYsxSmB7Geg0
P97XgKx7KX1ixL92uklNFFdT6cpnXgK9kD6x9DPfF+pqy4u615orCPXvxYVABU4d
l9q38cITv4G6aqiCwr4fY+L8iwK88Xxiq4DrggNm/99M4N1l8496cEXTXB3hTEgE
GHzvQ4b5HZMPjzPHqMYytuP8aGryiA4VYyGgbPFyFEzUZBuBuPJM8RYUozy0GK1E
iltgn/aExP17dlvkahBks37mxjdmcxNZwHFBIsv2dNL3E+WrVBLk2zRNJjZI0N9Q
Nxhy+gbUrrefyFf1AgesepFa7tCf0J6WMw8nFW0EikwWcNIOBeugZW8/ET2o9j2W
fZ+6LTMRE/fhNlIetRFyQqx0urHgM/5hoFOHIYNFgGbADL3/S8tuYB2OwXQHDeMY
G3pTYfs4nj3crjsrQy63FrHxqx7I+itKvNzACzZmbnM4RALTokjWehOzV6zVdrhJ
33yzOWo3f3PW6ZD1+c1BzpQPQjdxfwDD6u8tC9dmogpUD0dqPCDXBLaKOqcBIbIo
z+RwsqU2lU85NOlaTpB8AgK/y0VsT07Nedb7p4jthzDVf5G0+vkOnICWpnUKUlWS
wWHwx+y/6CLHaOgodroQf8e69E9azQw9Yo1VqwEnVmg8uhiK3fB5M+aIGmQw6bTu
HnTX5jGaA+p1PZrJKONGsBqlGw4m6Lo6HuGINt7uONefWcaZKWuhM45j9vya9JqV
E2ih3ZBoB/YoXohkLpmLg/8UiFucItiJWBARSgo1cPYnaGVBe81BTs4YXsOlbzo8
J8K0c9l59jkbn2cWtP16wNR3J3VpA7cplPq+08DDpZS7Wp4dBNeqNUUCCI7MPfQE
V5xDg+2j2nWKYrebP6pNaM8lHpZ80RUrUH0g+bt0AXqz0OE3j88UPUMwR8y0CBLz
HhuPzM0px8i1DdGjYyDHnDIa9C/yJ/m8AdFkaaLKzIujTEUONVml+JUk7yGJBI2G
4+k0KQbzFfPlQSL/Zd68KgeA2vrJuheWm+b6mOI4aKeYKnn2YjcbbC4n6WlzxMki
7wCawTNPd5r5+jGLyt5u2uAQi6mRYG/2h/TeCUNxjYj5UvMnJG/ZuLUkEZbad81S
I3chs8dhXossD/IBTk66znj0CMspCy3pAHfkovQGSKQtetLYdUhUIqW/+TEIImFr
1jIFrpRDqbaOO5yg0T5Kt7OZFOYSGM7ZSkuvM1bIC/0JEdqoQSIF37WBflTEVXSE
eQIs9itRPVoF4XdkiHrmAK6wb/6L5PB0VTjOhjOaS5fc0dHbPDsc+Nh8ealaVH71
gg7BNm5XgU00ag/0hhvx3DlkBQq400HSXrezTnRdpOH+wrbIpXZv2NXzScHpIWbs
AL6Sj9NJ9+IBMuukC9006czhr59UyCBnz2ZIFnlu0qSjSygUi2Vm5IVcRJWHCG6l
quPIPiWG1WwiQZJLBcE9QPYVLMrd4jJ3jKSqSNabsQ4L3QI7/6/bYVbp8xTctyKJ
XOVtIzWRduKwfMbMaLgnUupCS5UuIzM9W2pwa1oWLZZ0JSRT6u7NoNV1q1NvgRsb
RwWFJO9Z86k4q8r6zpMyOWzyih+UDmAig5GWhQukf8ZUr/LHjmvrvDAPKt7C9N6k
uwWzfp75JiR8oidcVl4XbxDBpc6e10z58zhYVkSRj7GVLkWpjALx7iA1TvMj4sqY
uemGilMMpbms7BWIWbaqRuFjoQsvBtUGPGPfekBynzm9x/lZPRNvNlQYXfsCubvt
vR5//ABKU3dLP8TgsTJuuXzxKi/ahAJAM0CJ4jQOXFCBqJMMYoypLonq7NO8zOsd
vOgDiBPJFbLpVl8tYhGkEJQzN+2iZGZ8fu0EYAjiUIMVhcAig/uvxdMSMSf0910l
mCQrQQwDImtw8/oTSK79B+jL2svz6Bxog8cUadWoJ174OXg7KZ8j67eJMM59yL3r
ZwjNNb5xAF3yGXriylkrTNbq9KS+lg3BzGe3hp+o5Lb4J03E2CbMiOewEyOr4N/e
XsHeokcwu4VWnbq0QhV769JSg8F8KJrjEUv3ezlPOA+yXGxu7M31OgU9YeL17srY
n9fjHoNnyv264XwUFtNh8H1S/DmWFvOgC0ndpK87gyS5te57hJPeP2gHuWtKRmUS
3izyPde8ljO63zWZNRnfUezQidts7gy5NAvuz/rPSTqUjSNpcxzKbes4Jp1UTJRq
ckg+3wPYfSNmQu5RtsdbxpR6hdej+QRJPCs2Hk4UREFvoPA2sCxKVkRTWcyHttbU
AdQC9Av8ZhnXILQ2ScoEoVt5NCb0sA1qXHbfUFAMSogecRn4u6alyv8DzfCodhkb
UeXz/0b7EGL7jRdWeuLy3APjdrN8TarTTU0zYOXVLpxAfdIMbW1kneMMj365uDME
+j+kktRSH8okJnuDDvEATCifDv9EKzbWHOlKDmGt9l0ZTeC4ZJt8gC2njUHJ31g0
FTRfQP6Dd/PLnOgene2ert6gb8z0qRt8sZDnH9e9tQrZOddaXrY5XlJE6ErxnD3P
l5r8SgF5NDAluV7oZCg11y/QsH265PGWfj/E/7z7dAfUtFpzai1QpOUjY7++OpF/
qF1RDu7Wt+VEMaanSc4+MhiEuqmMfurv/1qD0PTX5gf9/VAdKY1AgIuBb2Q5MZJi
rT4SAlYzj+ZNzU51kC11fWvoVQqnTgCq11X25qc6o1dCZOMcZHicQ8DG8qeNNKXS
Le0LtdhHMK1jAwGpVJ6bjyWBKZMS3M7qjdOfgnKBTEmKp+kMcdmXf4iMFstqxeEH
IXxTT4bZ/xKDMwSAvMAc+yIz3PQuj8D9GXMAfvjy5+BMBvVTuDlHjDJGhHaRY5Aa
70FIW6cQ2AYqC2CVljFDRHA1i34LLfA4zv5svoszow2N9DNSHr1H0/VAPCVDwBjx
uEAGU+sqewQGL9FeCeWSrhwM5GIq6zncrBoANmsmXVGOtfSAi6ENGtmNl45MihUT
EQhfDrO3SFPMhOagSOg0Lmasz2U2J6hFFi1CMfTzcQlSYge9ujVm/ngc2Hxbf9Xq
bUpNpyuqQ1oB7KHYaslrNmdZYv8ChNrVtNIV3xAYK5dbbmYSBerGrDCT9TMkF6OZ
DkfqwV1IaTlBJcikrc4rZ+IIAzLsyaLWB8zyC7Am1T3VrJuiIlEoKshZ9f08wgnA
M7Fp/t4Dqg773r3PcATm6OvrhAsfmcJQSxRfQMLQgnO1E4yPjRGg17g6Gy1fe4N2
KqjAh3gbVS4NQ+Wx1tjJl83DXi3RgpDV2dhucTuqy1c3IEQw1b9XfFkm8VRpk7rK
OogBLqeSEcLA2/af635KSj+GFtWR7Aj7UlyPEvez9n3ezxZLmIutSJHkUgHjn+KJ
hnaTqIOBSPE+x10FfxWtgDs7vTemCYZgHWG2zJpubx/Np1mIs4BJkWIcB8+zEE1o
zdHucEVpifncHcWbJaca3kn1rAxp4wdQxJbK3ymju4PKU3io+eqfFmDkhFBudI59
rvLIlIST56d2hPZVcKGq3mRl5c7QPhufpX2zQNabKoSDL362ZxawwXY59GBSnS+C
v75CppTcX0pzveIpKGk7FIHcRNozVXKcdeUaIYnebFjonXkd/1uQ+tLz6utGFUz0
BsAb6bG35YyLh/6Uo3YlvHMFgS7mB6kLQpUqnCtbk0/dQ7OYtCECnvXXSU4lXyl6
iLKKPCR08nB3ywKhP4FTMdYXSmQ95WonfGl+YIr8K5woyVrmXclOJI6q1V8wEf6h
lsdeXXQdgu5rGm7JzjD01S/fd1XO6tCqj2GMHXOII0CL0s/5MBNQ21B/f4BQsfGO
0FGJoKQonzA+pOjPzvGumg2c1KrCn39VQOvWqQmNqNZpSHTaJX/NsRIgIgBoQdWb
wLI7F7vcDc8ZRkysnJNrfq/vZLY0wbWD0DHiiEU/500VKdj21ituium0BzU/mRrI
50vFUVboz0X5cHgGfpZuCqHsXInqx8pFGLd36SSqIfv89xyjVyKRj0mXuqWWqB/R
NNFr4NIko4EWapCE/zk7x4/iv65vfAMvAHRVbS4wLYHWj720XmDM1U9eO/YRbTxR
bo5ypuTCN/oTQgFV2KOxCaCmi7iP5gj98tb4pXDO85KRD4TGxvfw44F09Y2To9F3
XHeX8N2ntD8vkUtWSfTq3BXBHzlp+Q4/mYyP+65Ga6pTHrRPq8GwBpYQgIzC8vGl
AKJkJXYLfjEYdHpL4g+XbBvOHXOa+m3Y100xUTY4Nny6L7EM6ax2gEcfklJEO7hU
pceMPRJ/z87s0zlSwjKnbPlOZ2D8m065s/d/Xhi1QF2XXG7ofDekcCFbkJ6R4CM/
DYvve03EW3J9+6hqadTIfEpqbGP0hEt8pczpoKx3/Mvg10Jx2FExvtbQHAkqd7cs
zUznsYiPmqsro3XtZCqbGKTgm5ancdjxIud4jKr+MTquV/DUITrYx7Ld72iFE6XY
qjO5wmxnjhIPGHRy1pxiA0s/MHBHAEnwYzmC4aF1eAaI6HlJQRBL/sCbMuk6GkwR
znQMifscYRGWZTTX+2ih8sIrhEyPy0mSM2hPYrSZGso+dUXVvsUfuEAlcdfweZOw
sKJbNzuAX/azD924y2kIAPHXCFrAYwTk1v0RBNVPl+oimOvT/bcH79YnepnzyXCI
wOxcbJOSGmQ5WcaeJhjxf2uUQL5585ZOy6UcW8DZUlqsz0WwK66rUtMoSwW7IiUP
Z4waALn+/3EuPL2zqxIksEfPVbxktXLiKAjw8+GIUFg71VeelTBcFeEiFnTmaaQz
OAp8DENlqq1BHobJpSMQ4HGbExQwJycl39Juf6zJ0tXzoXwOK88JDOUTiSxjX1qQ
tOsbm0n7df1JmGmFd8h83uMCccQ2xSvV7NK/+3VrO6552UNfvWDheSw1h5Ok+fXe
1i1Q6/kYoAni0aQfZUvPcQ==

`pragma protect end_protected
