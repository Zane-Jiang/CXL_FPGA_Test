// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S5hHqRUmO2QeW37mh9IB63EY4zFkxGUdvNE2hq4LV2r349SkHk+n2Lz2xQl4
2zj8e5Yc04nM7tNCVLBIWbdqsAscLuJ6C77n3RW0nE/wmuKh/V5A8ptHP61v
RHkgQEEZHEf+xtQnrDidKyEQNMQatyz7de7aSQf2vzoBs778AzgJB/kXvJrw
VNe1dmRZaBa6MD0HLpP10SRAGnTtNx7r/s5lwCTYoDlMXJRCNXMRIjaRd4mP
B8DZ+nmw6Bc3rIyHyUJpc8FW7IHPzikKmIymG+H+PiIgvCPMHad1ehLFhulv
h7E4A6XPia0eF3VFbvBG1VYjHGMUmd6LLwqXgzr6jg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AGBSsUT0cK2z/2QGtCEBDgRhwHGLeuGnLcjQDz/57fozO1q0U/qo1YF6q5Ww
21bGuVbD1D9wdaJGFwnbeYPWmwWfqe+XhOCVOjCH7OQT5dntbrLoM/k4qbNK
9RFCsFJFBnxfLKdtJCrZ3omHdk+SzDt9iP/SEXDMfkfnY5ODuk1kFYRPsfTF
uK8So2W3WnNUBHoEJkhpYYiICs2tOL65uExVCFmrYeIbDRBRaaIOm2sNF/Uh
Ah+GQ4ajTde4VzR/Ly+CKmob9bipxubZW+LWhR4Dp8kK/ValRV7WTJJmqie/
Vtfnut8CR6vhDN+vUBQgoFU5PvJxvGerMk4hXe4Gfw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iPNN4Lk9UOy0Wd75X5FaAnTez0edozES+1LAaLU9BP+TcRC2N4Sg2QN4beNF
iePumpgK+LTc2difHNiZk8OFdBRqPBYujY1/+enNBv/xc1jiKBsdgOtD6Flb
4QZ8PkSQl/HoRQdgRzmjQVFYT+DPePSF8I0ERdYe5r7i7xyjPZIKKNjAgMq7
gDKvVqN3aQKNHl7cSYPA4BxSDdyC/kvj45bPUnaMomJGIk/NEy99LcSFuZ9W
MW1A9+cmUEh5RtOWfV7vHMMeZlEDD62XqE1VLqfFgXVbpPHq3S9jYUXd1zi5
730r+0ED4RUEpTzu42okabF7GeC5cpaZE9KArWMFcg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q+X+NxWGaXSFd2LghLhUz1UGm+2q5kDnqoTjkeVtbO6TqcV7TUb108soX5GV
kwycVfiusC8Yo/eTlHFe4IIpfko9aRifPCBq/fJ1OoFQ13eOMMpgox2Fnx0H
Yc0eMrQOOTyh04J/dKJjRLm5rK9UDDE7JPdGogyeYsudxOiz0AQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GcnbZu6T8ASokZhOX50opEfX1WyAS3dL5bndQKy4ByXFzQMVF0zdaPYupCUv
Ckr1hfXBvgT4xfRywyfVWH/VvDzMyle5UjXOHw1mXlXwRx6qeZxG+NbXdBqw
AHE9LHl8wNKa2Q14Cut/Tmn7AX12Q8izY3xf5JsN/OIktHBvcU/0m3Tu8T+C
85lI/Sh62sXHsyzfrdUEy2BKix9Aj6oEo7QdFpSkMqXVbOErV3YF2TCJfNYi
TB1I9zgzKFG+fos+syi7w4i6pW6aHbdZdC/2gQjFBkF5LXrqAvM3wWm5dvJQ
gjaiil8XJ5OR+3YsRdmtv8e5NHTuJLYTgby/fFTOBRfuPZmu0kt6urKPL62/
jPy+KSCxWqbqTBsYsY2m/eBLdiLi9zlTez0DP5eVsj37LaWV6s1PShW9Rwtd
s/UPqPouZrJ7cKWrG6+U0TIJV7HWqY/T6JmDteXn6l/K6KA/4GE8OiflWNdi
HBP9zEPSgduuB7Kiv5psEXsDlaiLqE8I


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vb8EUGs8tHBirKSp34di4RpoPIBUf6bA9CWpM9QtMj7UmOVhnG4zWfW1TACk
3l1Fy9U7cr6NWdHL0FxAd5KsJfDHP7DeCYP5xAafTLeE8lhU7cD+kn81qlhv
AJlZCw1nsqLv7RiHXqVz+46MAbrqQCAlaOqVqRHWSafA9F+YOnk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Iwy+OVCRiu7AEHYl4jleh5x13y7uPG3idPuZaxpHm2K84CMkD067NmVwn9ij
Jnwm5es2Ug+Pwq4QpLhnQtMG8Bqt+u9VRsmVh7GruLtDnKKwlT7WUz5EDnNt
FmpXURz4glQW6XxKA4SosC0GGIqeJH8ETYUvBaqEityAvjmUez0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
91n+QhuRM+g6ksTWcIhMHpUmrnsEZWiY8dkzDSNb+Rcl4xL/P/qD5GVNG73P
uZ7FDnRGT9YqW3WreXpafJMcPdBz3LlXgg4ZH4cnnN65TBdUAFQ+Cl/uF6sA
4yCwDY2aKIiGFr7/+PAu7paEKAwfzgAA6sjjfbCODKIFoej+Q7eZGrDv962L
FU0r0o1Yw2gG8bYo7RTxR1zqFwbWxL+g9vnz1Lgl1dmF3xzNpWLGGoAyB+sm
pcazimuyzTQsh7ooKXUQF2IsM3uMHxi/xKAibqXC4JWVi7XtileADq/nlYEO
F+sygJyN1c6+0/0kyDqiebOG7Rw5asCqhXA5j+6N65ha+Oy4wxt8bo6fUqYf
GjNnEVm3ksf+fSdylQYSGctqybktKs5Lk8zARYFkPDjAVd9+tzQJ+bVhWnb3
K8yGyMIKN346GHZ9LX+Ki8nhWgAeVC9cqCZnOD0rQbtrpI/6lZV2vtSQdapf
NUPiw+5dI+MAcHod3Q/6V533aawmIwzc5qymQNCLZkcBpITQjG8+Cl6ih8bg
dmfrmj+JJl5S1mW6ZOo9GSx3fyQJwoFylVQbcGrJqPTN5jpkUxZkB6drLzog
GBB2aZowVsJjsEy15jkXU1qC0we34MwR6uwGRrdAk9z3EislwPKZX1DA3nhn
BkxPRP+JWmBnpjZhHqpbxKeeBte2pdLiCmEu+UlyTVtMG0WFh6YfNMpqGuNa
39Jus4TmZyMJafpHyeOncKzaLJbj8OUVRQOIW94iPB1Kk/pYxY4nNrKyEuMr
/1C/GiF+d33kn78+HeicVPJnHVoAMnYTflKucPP9XUU5E/qOcwG6tfGp/6BF
UzKvArQorQUwfyZb/+lqBHN/5PEkoNUhw9j5DVCQQkwtmTZKlCzbNFiZyL86
Tao4KiazmiOagvEF5iSnRMHQVaii7LHPBwmUoWOX62wJ8QL6dVtv+rmW+nTn
jzw2RMDaHv0dGXO6uM4WygevSepFR30PpTrzHyPUlr9i8gIwq4arcxeZ/pjM
x3ZvNaopSTglrGSgMWrs8Ei/SbLRka5JZMPgd0YaafvXvazJm3gjd4+xLRS3
ttWVFo9D44UHIajoso/JAoqThzQ1B+QV5vXK7xQGUlYC/ucaIQ0A6C530PHB
+qMYy9x7CZ0KYoa3o9OoXO1vkpD4+B1ceeN8cJ/sXYvCiJE60n5RlGGKDDaA
pyf502cBXaNn7TCBDub0jPa3DXmfAFUPRJCgvo7gtSihIutLOv7H+qNCbQ2+
UMZEN30VwG81V+DxAcNG3TJm/4L99r+G65gJcNUq1md1c/SjOduNcANC9gyq
iUfc8zgaR3EUk4dzawKnR15Lb25DD3U9fk8DiPhmSJT6wJwUT5R0BhjDCvGk
/w4tRLNCCspXh+dcETPSLMo8J14HMTxZuPIdUSbfts9CVzL3Ni3n1rJRgabt
enhBNRZGV0UG3Przf4HCTZbYvj7P5do1U25ImKjskR259r9O1Yohsy30PWVq
hYCZOJrMnCOd7TfQLDHKM/WzuVlBeFg+d3RWNCrLOd+2ykmufUEMufYnUkA9
tfZfEEr8Qfv2ARiZt63GFcT4TruFK9zw6JhfLB8sMKTi8x46qaTuingAQ7HW
9E5NezOauRlQrqOBP0cvHRT+muA5fUs4+xAous/kIO88Z+62b5EUev1YCmiX
ah/cmPHKjHBM3Pwgy6FEG/j9sRFJdCJnxRF9C0R9SGE8m7OnoxMyWLnIDaZA
mfgUa8QubudEhMV3zjyGEZD/0ZyYv+VmZZCxqbwJmFND8sVEg2U1qi00XFwB
36qd6HFhRGppzLTX9shmy0vhaFjcUNMkT/4=

`pragma protect end_protected
