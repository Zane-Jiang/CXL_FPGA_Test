// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
FmpLQNF1LAlI68Jk3C/xPyR72dh2xvaDjCOLwFt+YqgUpMUpEBaC6W/Ic/pegglg
PyM7PBRLbzLqcoAEPBBXS70wgZ1cgEJDUOtsHbAfNlr8Y1nmShxB7L2nJii1yZpn
ABp+9E3aL6SkRwz+degX0oZdXCXJz/9q2s8veNLB3n8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6688 )
`pragma protect data_block
z4zP9GQK3cA6Xg+CK23OUKCLy1qbC2FwYz5cVEb32Iu+o2v74f8/otSnryQOo0yx
rd4YcmBuH7fgHQEEqD43zExBEIGC+8RerOv34ejLiPT0oFOezZbaZDzK8ZRgFk4j
AFApiDheO90DReRBuJy8xFsAPH5APof1k9gh4y+C9FCiOxZU5fXYA3uS1AnY3fwO
93ldKcnBionHoWbNiq2UBK45OyG7rkbJCnlmbb9gaHX7iOetgyAdZICL0royyXmZ
dCRj3NRH2AI66UFIU1asxpZbQTC4Pipmcl4n8csT0zRk8QYxgSSYiuGQLS18XTIo
bJObj2qTA2gsj/aZdUFLZG1riPy/5GH3xlsMJfGCiP3kqSOYRKSd+5D9YTtKH5Io
QryIwPnuylpU1vzngE3IZxNlOHRqTjfvmudQIbP8wNQ0J5VzFgxzxC30UEo/RnIZ
0bKTxpeiSfECPlnQ/X4E3C/3hEFPSqb85tYB+oiOnyf0GeRpkGU+OEQzQHCfTEqY
LJvVn9RnrNkSUolqVDcIhuItDCi7Ag+TMUIslh8ParmSZGQ6wXZOpNBWx+6pXqtm
B4NYVt7jkyzagmsVGQTWtDg8j75YfGBE5znFHmRFeHUFBmyGBAwIa8IzJ0ct7xYV
25jUqnieLKPHCO/0FvE32Vq2NkuEBo31CeThZRZUaCRlx1/l8T4yH0pI3O3c4DU2
slseMPPF2hXnEBCLDoLNOF/z4n+YXXIBNOaSE+lJtC5f0ocTJEYYMlRqe5cSxnUv
k0LR35SDZoxZT1nfSrpT+eFN5CEmaMJTQxE3JHyb/4RUH5F+8EO5MNJogT7nfejt
/miNoC6cRdKbOvYLIl0mj4Qh+mNOdGgqNtsz/RRQdLtZg+7cHeOFLe0Ysyha5E9l
rt4aMjhUacKWwEYouXAC8KBhZxPCiYDomqSFDopz3psIXEyKN0huW2kn60lkixFZ
yUc2jWq8rfathAwO4xz4MEl52ryMhE6uk7FLlO8LJ+qmqlFB8hHRrUbL+jsUEgyu
YOjx5iyQli6zU+FEdss/OHOlhAFrZr0raWww+g05aZe8Edje6U9Wc+1BxhlzWKIL
/qsmri/jFt0LXcT/6ezR6cieKOyZhneshX9otsvTO/0fgd0S//MQwUnaTG7kXcpi
NaYO8GeVaJ1y3XvqOmFspJEI0pF9+5sTYOQlKAQBG6X3CJR//ZR28pJMx48/mwZG
+xBFUAHbINPHOsC42o7vijcX4hVu1mk7O3fudAD8dO4tJXGHB9u3MZe+edNCwE2q
nypIsxew/2HmCLnrZ9wgLJr2GvPvJWrRoK96uqg2aTcclB90XMYm5Y8OObX+5ttV
Lad6L3GX5XiLU4Bgb6wVIFfWy38om/hkxhF/Vs+jmo1UCYmMtNCfRPndgDzlBdlU
mt0AoZ50WAXvvMnXhRjs8FbsF2DkyNydJnC8b++I4vqj2rnBJm+AxFw6z3Q1u/8w
Dtz/KGqm72unAAs2gg1K8O8c+G7DglUDJBzp45tjXLgB2EfU1RlgKzRqpLUlGyJa
BoQvIQODSER56Yd64XA3Zg6f5k5L6fuZlqRmDmmRE2ffjDNzxJEBm0pyMMO1vRie
Jsd+0BJUo2VPYnUeQbVqSEb5CD9Nz/Ba5/tP5UTxtf2sQReqgjF9CXW/tCZBq3MG
nYVCQab0TAyWqcgzc3QLyLDxIJmT60FZsPhMo80RZcghOQFw4CzUTGVDWedz5wkf
briNM1q88AH1lPYrnguKMsyhpURPYee2YBYe0rUfSMKvN8zwF3Pb2gQcGeOVIHz4
qsHmDGMCdoRDl34zteVpgD6nYiDxQ1yOWSUJOZo14fQiRIF4iS+ad3xDicwuU+di
QDWkADKU5h/bBVNIktFi1toKHBtiEp6zcj5hdYf11T+P5OkhvnpZBT4i0rWcnsEE
3cVOttFSQS80Y+lEN8ohhHsu7N/0b6MrWjmMhoff5MHrlTFI1YqkFf03wbyoNjzZ
BWKTzuIpB5LW0Wq52SIAmYXnRlwyg9vyIW1gPPYqY55YipdrDpE/ICO5vnm+HOQU
Hhn/tdxU+ZwS9hryz7eYafBqDhwcR1MxUK4SSFHcpES93ZvbglG2QWYtzMsmO90V
Qbz0BGGxkULZ+GAHHOcxkSf1gyvXPTb0F0KykAzsn+lyvwOGF21ywGBo55U+HiO2
tnvfHw0jxbJbqCHS8EftjxBGz4d6nn6GDopilrY4BKbkFPqvoqklenT/dM/cVzSv
UYAQelujvQ5zOhDWhV7TiyNQNnv0bmKk2wYgPtI6M1e3AVLpA8spOFmiigzTYUSf
U0gWx2ANlsKBqnLiIKSfpH2G/iZ0Erfm6y1jh9Y5uX/GRQ7RqYNrwvj3162F+vPy
08n+Txcuoy86QKN2lfzYAxX1n6lvvGm3ZCT9ByVA3dRzjfvfO5CB60k3xYxOO3oq
xRMWGSdHfWIoxoJvFYYmYBls6ogiUItH3WcpRBcpx3A6HKfzhhyGEIAg06kitAsg
Px3zLmpBvgK2IwDkWCATfmjmlcQBtUOCL2WrQ1ph1OsMcRYlPUeLtKsanKcV1tp9
3nXs/8UaCmLWDh7W8rrJWSEkZeiyfMgvPDHTzub7R8CXAQzW4OmVE+nuhkcS4MBe
Wud7saZkiLLFvzockg34/WARwIJSyyz373rOoYPw7DeliAUPsYYNauWU0/+wvvxb
vdNas6TJ6Qxpgh/ZaAJ8vVqPykirqMfs7xjSc/AXihMGMSQoECTVFJkg7Air7gJT
j4Mbx5ys7yLj6Z0b7wp6oGsabCCVBM2HEqSYANKvTKqMVESaX2RM+eyQDet66M3w
YYw3cnwAet/Y9sMlvTTURt1gxae42GxI8/ApPKUacgL/qm7T2Q5TntYgSRBdIkUO
9Uc7azNzBU96heffyfDhBabTW5AkDLiqafLtDbj265n1fmr9aSsom5bE6IBSANhD
QJbkrxX+LZkaj8341kpodxydF9po12GEeId58TfNlZyZ/30UEA5NqhsneFcWf/2U
D3NXFoMO3y8NHbwvDlfAQ3ZenehXIf4IuSK4jrznKEwIg/XBiOrsVmcckKH2i3UN
NdyIunIRKn4bi/pRBAzEeJvPgH6nr7glAmbvrrfVzXqBqXOHkFWEdJ4E70EAxds0
NIGEzCvVEEssIJD62ZlZdEcT/E+yD1W6jYwbNCKeDmoXQ8Vk1eGeBJNYByW3qAbC
2y9Q+d6rwRyL1VN9Oaa5GXGxpnY26BEYsMraPa2IPWl1miANI+h7S322wpRnLqRF
hLZRQUG45aN7DYxxdEncG6jLd476uqfDh2mE0FkiDNFfPkcyiH5XjOKj74RySJIS
M6UUyimsDvthJEf1EuT73sswNtno3A4T2PVXtMlr/UHuULXPqpP93gMPqBEg0sPS
GCCBZAtBBAbrVlJ7Rrq1iJrzXjH7hgON/zNc6Od+M2R1TkHOrgQ+5a43YWxQkhtd
5/ss5lGcfU0cctZ5E7MN4etM5ZryTquqyj0ePWY8rsc/4YvqbbkToqiWjQsyoJkc
fg3jT0vWZvwpRlC45nzK+WY3sGHRhLDjmRdOb0FEea+KGCirgUyQNxtS7NFGnJWk
yOhQ/W8khafwjycYOyaszmxvvb/4TkNJLcNYBysihpFhINdZ/OwLMnx1t4y3HPjN
1wqdjBlQzDqzDCJVsga/cV9Je/geGlPMJ6ZN8ZtNmeg+TE5SuO5Zcl2nW6WUAGfs
Mb3cJbsx0pX3tdFMEt2IDx8LZBi1bUpXBXnUjVqX0wSlyE4b7ox1J/K7PPuQyBhm
aRb2gF6lkX9i80JrmDOaLdO4cForcK8cypQSwZErESoJdprGD4x/hDI4oxnGBQFX
yqGw0Nmo2FcmbbxbNFB4dWbReaqfdSkNGpq514BiDB1xrgiHwLcJZvkzkrQPDIJW
GOphKQFbBy7IJWcx7gUcnshSHfK6KC/U/TDP7Q4BXXhsb1wDUWgT1t1guaGYrEvF
Xof8lWp5aEc6yEejrI6WvF1m4k3HHENlnrGGvH/n+N4hAJ/1H5mbInCS4+UMl5jH
jnmKJhNr/S/2LLHWHSptIckIxkH0dVbov8jd3wYh0v0633/AommCZdKBsDgrDJdt
KFwJCqLKMbKEx1sGJqf31R0tnB+kpOFA/kVoNn6r42mh+KnNZg7/+vYb2BgVRd/e
TZaR1r0t6F7Gi1Bcmf5ttLJsFZw+4QNPU7bz3KUnOYQOd95Yny3R2Sx+ptNJczNU
QP5zNwe0wKnBBQrifAKI/YwBeeFrS6DyuuGGQ5+QfUsbu1a4/sUzZoYXfO8A0O1h
C7AgkA8ys/tuWoz1AfPsoz10L1CGhSU8mlIgFk2hx3id9B+k8wNms68mOOP2pL/u
TV44LMTVzmctyr5ddUozgFL2RyKLR+nk6JYHo3tCFNuy4rBDfcedAwDQQHC0mcG/
HRy+JXEJKB1be28fq9HI+qQrhcxnkOJ2tpjmQCWS4v+9OB9k2G5LtktRIZPMQDiu
Cz6chVCQctCewfMB71LZH1E0Q2OCrVw9jlTpPldEty8/Eqw3ZtfdwCi9Wq5/jMyU
p8gPGw3Mi7G+pkqwt/YIZWdjOCBVLFKy4IaV30uSzRzaFEKrZGFK719yIZyhzGCS
64h1O88Uu4TUduiWb/Xb98WeNHBgAzSmQ8ycGZbJNhwRl/LFhLKZebdjB/GIJ7g5
HgG4a91G2G9Ji2LCnWgxGhRiirRLRmmnsGqz3kCezY50bQKDFv7Xs9Iws6mAIaJN
J1o3mgIpDg36DFqWvnWRZjz+hDAPRu9it2602l6gbKCIimQ2lY/uuf5N6SWwzNdf
5StYSa/o/xfQZOyj5nOleZGb8yTTZV63kHQkICUnBPY3KRL8b0YW3KCQUmvZKYJ/
H33I70s/HrTU0YfO4Tcl4u9Pbi/mMU0kHQQ6sxyDrTOKz6IpRS05GQ+UyeV3yUIH
OxWAWwaZujFIRJS6p6c+njfPRBAFDOs+jqisI9sGWKhlkkxIfO8RhOq3x4WoGkbM
383x7VoVRCzyiWOKyxX8HhAoLWBBj/fyPE97feZlvsRyGPzy6RrDANXUEDV2puzk
DhZgTEL14aISINishvnfuoRDqO+r6VZtK0KesTbW4dZfQoBDYQI3iyISpaUIOaWg
vnX8aaKqJhhJyn5/67K38/fWKVkVltw6+pgHmq+Ko1TCbJ4qyBwwgdvNzH0l0Tt0
vrWuRrcLCoePKEz47akdn8BnPwsp9+SO7KQ0b6UEwV7WsZy6GB73Su/Y67t20DU6
yl0VCRZWncgOtAdSfGa+zPDE6aVjBuYC1OWXJ9j5pRg5USUU9EwJzRNNmA1EeIeC
DZpYKkbtKb4yenfkmD/CVQhAugmwebrI+qoiu9KuLJftYhzwIPQu+gPRKCsjZ4CR
bRIqF8r2YIqiNhQc01eMNv+0fLNlaqWEHyBWiU4xUYBM87ueqU9RHE8NcqoFpnaK
9mqdU8qn3jBOtdihpxLgZAHqhjV+OvHOvLHYfJzEJGG1eD4Ddm0P0WQXSpeQnTE6
ivAliFphjq5X/3RjNIJZAZ+ThLwfnYIKgJE8dA+zhP68vV6xf3zbAWi4hHgTllSp
yjP+6Z4QGPS/YcqST4VX0RbOEthVKcdwxiZrmFNvy2Y/w+EVh4082bB2vMtIIDyV
D+Ed83fIUL0X8XzITe6xmKsH2rgOLxr4q00MIn8eh3mvDQTy4b/YHjwmnQuk1W2g
EdxQlnurKqjROU+H79DwE6V5L4kxw0ztf9VpUmhB8lgSvFQ7cVkpwYSwN1Q3RGcH
Ngt3QFPvSpbpld2UqFE7MjEyymvds/F0HPZfZDnUpatZ5eYbBsBxc1pe1sVZNVMI
052VjhEK8QdC0UIy7UqQL1CECXtl0TPGD58oksdSPwiqckAT3Rgv9uCbbANVzuKn
6NoNzkezjBN7PcqCFbm0JcTbH3dhNfdIRLaVr3axwA7yx5wBl9vEKLeqZbxQm/C5
ZnWjA1lMXHeNVksQ2wQrxVLF9uimgPtHayvWW67jYp3wc7jhVYGxxgUMYaRY3DBA
BEn79P53PA1UGp1wxT1THj5fjGACAQprDdWo3TKEVOYaNTELRKsAURDX333/Z2OR
UAhAIByIVihUuQRfg/pcz5Tz2a4wjf8O+8wUNLcW4ZY1koQhlSd+jX52Wq37+G/W
wTeM4L4hyJ+9VDuZa9fIvd34IwyPsob/Q+BxP5V2zri4F6mlS1J9E3tYN8GQEXFJ
GEIpSdLnvX2bsuOmN2xCAZVGJllik3aRQi3FhAdpczJh1KVNatWKEW1cTZ5pNWVi
ozmv43v1gqGpG21vYA8FndG6QfX3OIKbak10rUr3o0ZLWpxBZH8JJsOlfqINIU9M
mSx1FvpVsLx9LNmdyclxpmkX3OThZLIsoRk0yX+dHWxHpICAIiQBIuBalWSl17z1
QP6dXd/kQm4idgJYCB0Q5RuTIMR4V8275+P5MXduPlFT3nZRZ1tp3H6Lb3iyDgcE
AxDsEFtWEl4liT4PPqBBTinakGwje11MVP2wqWQ0lHeIKJSlHu+4sSpSFNq1FKbB
VsfPDwxNijBlrarLIr3yY+5ekh/E12Y6NY1lGSeOrpMTQD0KXdHbjnmD/Q89ghD2
dmEaBQnb92LLXsROwUxOMw1fNqqAbkHHe6WuGpO5OLVS53AzYG7MQm9j4aZMzOz1
pDrxFdrm0Siy/EbtPpEyIivKwE6cR2EEQUpVUZIQWcOBI1Z2kg+dGHI8Y8q1QvPk
SHNEgKN7sHM4CEDsVrGOZz9j7+li9NBc256Hdi6N2WfCs0mq4JXISzkZSNqvTAmk
vDC3Yg7VxR+O2PX1THbeL6oc5k9vwqJvrC/ZTIdV++PTi+Ax+qKX9ItvlbZc5snl
PmLwGgAhOYkhv8hDvcBA4NJCcYNzq58VCdiXfpc02BgjHdu97RQilCnLVilu8zh9
s92eoPxZy2VmBIJ0mLMsuomSyrXT1EQpEOPP66C8GnDqdqQcwgmkEH6FUVCu1FdM
paRUc+DqPrnYMmvlUxX/IOlm0xRbC8zb5Xv4thGdoLNP3pEdgrs0blTGR2FR6ofN
Mqb51yjXhqqLen2YIG4eSt7Fhn9ph/lAz1JVGpoArYG3/9/EuFPyEHoRGU4HX9qA
SVO7tH8O1V3OVvm7IRkHQTeCFl6Bj4oK2QAD1R7ND6HTMTKWVy6NJ520+l8p4sB7
/jDduSH9zKEuTeL0DCIJFEiaIgQ4hAKkAQI4Jcc4ovSq3znl6M7vfgbbkbJntTM7
zJICjOSgtaHUIHzxyrblg6ul3vIN0a14xItA6p/EpIuuqAHWU1ADOp8d+yjxVF3G
eVR8GN2FeAchYxiZNeiyRbIrAhCSErERwXWuZD0JLaw0mGLYsQqe1iuSyvngZQja
gwLlAJo2eG/tk1vZPG1xh9MoO2q0fkP/O50iAplhAse87CFm+jBlxOUn9kKU7G0x
nNMg9bHHVHn4GppHvIVcwaUzAnS1G/KlEQgGK+BOXDbA5yEIiO80tgqXi11TJ6sB
GX+uBBcuWbN0BVz6ZZ398NFMlkJfTVK9yadll5WWQNQWGK3W9YaY4v9C4Mr6Mdk8
nJVUiZaT+RrRmt5Msav/X8avJz8h4pHDo4sPdkhtGg8dasJ2tnnQT9YXIj+ajqcg
rYqfOxKyjjIeU+EsNKZdI2Kgc2hj7fWFN5KMyZlK8sOwCNhwqY/KXR+a3UTAGlXr
g2wNfL26LIc5StKXBZlK8R75nCxZ3bmw0ifyQXkORFcJvc3S/I3EDMjYo1Jc45+c
mcnjjD0v/zcN1BxZF0K2zmKxPF0U+vV0CtMFhZmxzXKdpZsdZfDTfTgReguGkzNx
RE1leO7dAPT/GFoK4A+OhZ8KNL+zwUOAPfTosJZNvq+FDqV+0X4rik9f7gR6R5Lo
SgWaQNvGXwxJta2akHTLxN4lzwANh8swOx5IgwG3qedsngFzoknwf/Zf5tvCinnJ
nSHonXoeoHa3lYq8CKn9Gguj1Dmab3tZW92Q0qRlTSDC9jLQJL7SW88jEO+JdcNt
uxbEXgrgrBFkjQGGQQYQ4XgGCFvay1NLLkzwgbkkEmxLoYp/AHvLVJyyru9JgCZ2
CpdYXD70QmpkmYGnxE9lLJZGUSIJetG/v3S5+/jN9bZPpv1vMogNMjbtX8zsAyGO
SCmNQg3W1GFXRI9DPZIM3tXrXKyNVAKui1+8V1BAIcMVnRhARGWKI7cVG/SWzDDz
68Qc4i9EII4Z6H71vCWSrREhjuhAaoN4ndBj9qBgq3SXMKVt/6cnMxUf91PeQKQj
JtD1IvBJPDMekWs8xulP3IhLGfXmYWZ3nisra/k8yA4DZhOZ3rYsZc15wmhM9QBR
kGjwvznN7oNeRJy3VV42wms57XS5BO5OWscfBcGfhQ++pWNLzydRxPTDkZOAbjE8
cGRfBLGif+QEI6DtDH3SZJjvz6llzQwW5NYMSWQsAwfdWeY0xQQr1kJkIZHiEJN/
GhCUmgec315m/TlMRip03fBd5uSYZefdUJdtHdgf4Qlz9EXSOmIFZ6Qkp97dCy3M
uwo6LIWso9/9wjzrLep3rZ9hmZ2a0HupbvczFzb7ur70+eI2TqoSst13lDIPKKfY
T/yb67hJPUL2SxS8Owmo/chYhug725GkOi7yGxTThG9AZ8TLiZHWaQkD+XGXodAq
pQL3BuU5PNO2fDP+BHWy+pRf5BkObmu2awLbD3Jiu2RYNQ6ZnzEuYCB/rp73YMP/
DP1TMaLGX2JQCiP/IKY3YL+4zPIM9Jl+7nlaNLsHDLeOXmnW92sNxFK1WH5CAUG/
oboHhVl4+PoqtUQ+Of40oEntbNMNy3Hgl8W9MGOEM9AfMlplqjp+lfamjPLEcym/
Y/4/0eVIZVe4DJqJuyxwSOrXqeOtJ4AWQw0S3edl3OuRU43gOh7QEekzpZ1UrqlI
udBlYBRXJrFk3QA5VaVj/g==

`pragma protect end_protected
