`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
P3MjCpUZlCCjwGHV84H19oQvvXCyAhlUXNNh5kP1b94Ul3rLdp8yTP9tomNFLB99
RROMfgvbg+6z3WDoEcPNHYO61FSpxzxnb0P80kM6i2VkuPxr6h4fJCK4zrnoQdUJ
QYNspwDeo03OMstXTtEzFelQ2uUdlJuFCrjxHX0uM+s=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 14912), data_block
wnL1aZp6oi3B9ipR2nTiATVp6sEcPeUqFEmaJrbj5F7gsIcwjWi75pvSqXr6FZbF
KoO6FPQKbDGz6rqxkP4VxWayqMmGAb4xZxDcWFAjlDcs6jSoe6umPZTpJkM90axX
rBbve24GJhQvjFj5cUs+HWs7WZpNkrXoZjm4Lf5VjVYSs8n7+ASkAufWfgI+bh+C
leHRzlDIVHJQClfJh9Y9P1FeeK52QuEtggN66Jf5g+9rH6dDIWl+D4WxadkPZbfb
hFpABJBcFANUKu9cEheYvqjonaCBB4m846RYLNpVFhkF1J7kD0Rdgn2hOv9MkSdr
Y+SNGfX2eMmypulO66QpSnr37372fIOL5Xl8/HaBh0lyzPAa5QZqJnDGGi0TmWQS
Tk9w2DuNPbLRxhCQAAAMuxmP49IEpEKk1Mxw6CPVUYXuvCSX60mKmOAnSzJlohRp
mnISEnr2LXVfPjDCgwlg14bK3pHrBHWCKVDQ7zjHfGEtiO1U7ogd5KW4ZeJ0Lly0
h5galh+P6l+tYDzzsdmtQMw1UqPB4Cuj8BmzqNfTXQiVFj3AdjOeBREK8PBAzPjg
wST6ivNsZM8L9tqANdw3CG3KHq1dJY27wJu2vVICkQ/sVIvnkAgDMxFHzcB/NcdW
2BNKSqtXadoN9n0SaWzTYjIBic18DRwyYvSMqWrd+lhLN6QYCL64wIOMy/Yix4uc
wi9vFHtT4I4AWXVDQA6BLs2ZjZMy29Lfcu8vihitoheh7pJZepBhp6fxc6ZWcooj
GA07GBjb9JbMtDeEqBk7TTQRdGIjEqeOKJOWzAVu0ibyc/K/+R4qyNwfS8ncs2gH
gaXTcmw8lTuDiOBEHHpp6pCRciYzqY7Z7jCsOgOwtcw4MHkbLEv/Bq5Vn03eNvi3
/VeNCMs1bOrc9TgbIy+OEvvJNsMOKNSxmqgqz7s7SzLwH2snlRqlFPyf5PIWchiw
8XEJA9oq+Q0BIMbhSyJr343qFu9ewG9GHERHT1QU7jTW4IHDqBLRvjCuW2JIMYHF
qbYR61xYU1ca8UKygXe7Pn8l1/tkOlMcYr0Zp55on2Jqzd/9tukXIxBpe2OBq+Me
ggroOTinUNfdBLrgr7g4kiZ8FRiUApwyldB5t5G4HnxrTtZwZtsdyUt3xxdtji1A
MkR65ojayIrluhTpFVZHHeYmKI/+noRzDFuI2LOdBqTNIvCtT7tCINibOAD9UXKx
E+prtcLTuCQZIfCAmPDeyQ5y/vV3edKegzkHBhYJE4QYg4tufilFx/0CWWYxI4qC
y3Vb2jQa4NsKli8GW+RmTQvefjojbryL7X+DycgwS6geUFZ17Uo4XvxViXoR4Ej1
2m8A83KTUCLCY5nxcDyhDladKZIYhIjzSONp4bbxqcZmWhvveH8PgOpYmJMwXJUz
fdSIuE6TI0Ij0ws3QgrMAE0hk6iWHL64Ebdsx/a7dgGD740MtmoQBuw8Z0RffxKE
8Z9CkzQgZr7ir55kEBwtFCJ9l1sX1PUItuDKf5rWxNitL7b6slsX9nGWPWy+Utza
B2r1hMnjOS+CXhRm5Chrf8SbKMj5/NjQPgSdRG3XfbTDmr84RoboudqnN2VswOPj
8gkwymlPGSJ+0a4T40opWUsbnC1BQTWM2gZMBigla+PtSkZTEoBiUTzdNG7tTYsI
rpYRy1kokjObh+jBjoZIR9VTUuBuW+hxViOUkiYbIA1TmiFKivltBBDlKOFEpMux
kfC4gxEsSmfQ36BGbuohYh9JShVbGWpEalsd/p3z61z9XCVJhjn0EoOAAgHYlC2E
DWKvi+e9QSzUvony3xkvS+RWNP76+lZClgUIrV58bUasMLBFmubTUs1YvzizkBQM
F9n1CWHFaSpnImQn0qz/LH6SnfidBeCifbABcx+McPfXkSnlgHIrBQOo+9T/Q7za
q2sFklhj5mQQhYZ/IwOpdu/IA5xn8DOFfrsf9NQLkALO0s9UOpuCUGghPhAw/y90
W36IMsHrqNkyKD3Dk8q6xkfpXsH3y8Sdbjzm6mQBh5RhLxFcEbFKQ6NVMnrrfCiX
nqrF4LvBaBrQLcNR3fcPqq1rellivemfGNGYE4jAX/pGm6FTN7vXo0DS4hQM8O6Y
W58F1lq3sljjE5Er4HXCV+kmy1EsGg0k4Hp8JDTDH2vkW4PQAnNaEfJMscuyhAIM
Cs8OyDXaHCPOGubWl4M5mEFSjIRFtBxnLa6CRrM4SqhpRRVktJ4zprDC8VczQzJH
BxlbvzgfZJm/rjVErizlb8JIW4TjPDgBtKBoSKDv4CqdoqPw3Yo2hUlWsZ9T5UZz
opdkcuTn4qTn5j2mPjjZVEiRUgBeZhU/7p+xYqJDVp5XzFWVbzvkvV7M+PovdVrJ
rGG5tUyM2rhb+0a1pQZSmMgnr+8fJMxU+cBGPUOFMGofML85NDyNMGd7ooy72V81
OAAsfQkSM+/oqh7jl1XVfIXVU8meW8uS/aEwA7urQZ31wyJMbzYwP8Cb1On2StVi
c0SwZm2X37HqrfOSu/+RbpaI7JcVzoOKAVqlGJlhM7+pcReD8H3Oo17SvMwq8Ooz
NK9EjijNJeTARDvyPV9viIb+9t0c6uj8jOHdln+QNHbVj5SQgp9GlAujlRAzXubz
qcYLSHX0957efNDJZhuYZGNXleDG09ct6fr2CdpJdW1Bm8dmZn6v54HR3H8QVV+S
GePsSrBUfnOso54Pt1HaaorwZwK11a7057A757WKeVnmycnfCReb9hHjNOyjtZDc
HYBYougA/8hlLe9bT4cIcKXIUazi8uhAw/mWAh41yw2pojz5pRGH6Lf50Ye/BjEK
NAazSJbCoGnjP7prDfasumBI1novQG5I9QiBd4GZwm0gKqJzEgoPnQ/s++R5sBRx
O1J28byxgh5RTcpdJwXL0P5xr86XOyMmjrWLG72UrRUg1p/5F45Mg3HrY836yOVI
SAeQRhE8KfajUb0TfijnL3JGTtjILJRG27oBzRZWqNZ3Egf8RI0Pc9rfUr5SYL+Y
Mu6AXL46AWpQKO2eOo6hjNuLm9lamBhgSFEFQ9YhCACS/f08ot3GQgWAORbwH9U9
To12+4KAnbHmhaLNkaG4G13ZDWjHYtSqkQEc3W9LU0e4lkdC4K6jnBxytqmGeW+v
YpnzwQ9IDi1lTMhNiZ9uCa13vI7+sHcpuoFBwo72d9f0idQeczKbcM9k9HoR5p4S
U3lDUuNzWK6bWnpAaQ0C4Wdn89hgB9l4R8fDGsN61bOEYZdfmYrzCmO29Y5QkAoL
i/jJ0VRDCyqf1BZ2ihB1z5FgQ0tPP3Ki9cpNUAZqoDulnvbdIjpzVr6VHmoKXSyK
gjKv1/8IsG7zROROfjXyOYnVLeubq5Oru2q7lXCp1azdmW/xYAk7Fzp0JEDGXxbL
x25ZCUthMViM/nZAsf3912Vt7ko2OD7vm3DxZYBjeGjfBPTfiTj+qsm/3RcjXJKc
m3vyZ4e/E/kI9i9oQ/e+k5el18/HJO/rs76zf2oFsbiUclSVHuIgygMhA+ZGmc7C
aivR/C1SSaL4+Xy3EwhpnoFDm2e+QTbk39VqX3FY+FVp99kKXzLyYzRgcAApZNi1
mNm+JqS5OQesMGn4Y1rXZBEV7FlxGgv6uXMqCTqhLUVyFLGaFbhQbKF6uTJKNCgr
GgIUoM07+p1TydHi9+H81Y5jAPx6MuvxsNHPnZVcCaEibJ+g8pzwcmBshTymaRRn
Zm1pHFw32QbZDUujrUxiW/gjFuTI4UOOqQKg/eQB4kZuVHSEJriNA9cbEzpBK0L1
yK+RFRxVWvcQen6Ns5EpNzxsUOfF24IIkH3e9Anl0g21qrCGcsuR2TI3mORy14ka
taV6klY9/n1u2psWzYA99m54b9nIjipQNTEvqBT2rX+MCK2tOM26IcqxLza32qZz
fGYLu6lB57whKbgXS1jWeV7xQnc/Mi2RdyXj6ZEr1MQMOoqpRJrKhurs28W8JWOn
KeCMZqxNJUNIy2iOOJfygZe+8n+KFUZZNf9LBwAZ6KRlf/afdU9KYAMcpWZ6/y0R
rK8gKpSqLFUvc2rubg6dlYuhcieQJsWnpM5UzQP3nacHj0TnXFK7Z3AVtHtCXmCJ
wcghFaLc2tgxeJ9bF2ZShkEOf0wRyf2k0gK5N3cT3f8XTSzMfSEtO+k8AFq36VvN
JqmoUuGD41k+DyszBqGV/olVP6PkOAQKepoHHD5oLQEAKZx6EMF5mAGsfL5Xtv/b
9FVzSQanPv/RICcVm22hrJWLSFLhvGdue6xkJ1Pa6eoAmi1ps3cRv5F2wL37+uAb
DoxnxSWa0VOjgj/Ty9w7JZHbgQpog5CzARDkPF/0LDVMf4TMyJaR+Nahx5XjryL9
EZ6SJYrRZWUC1K5y2fagt5f2g8hV3qFT3qigkQWzsMHBMrPMOYEMsnlV43SZIDH0
Zl3JawM9lIgY23Rro6nhC6ST2m6OZxFAQl1vswtRbB8kUrsDnxPf61k28+kGETpC
quM4JhIY4oPTZC9Y5tByr8MrCOTdApK5iaNVe9SxMfcwgbvHbxSg5zF/JF+L5t0i
L0HTgjPQd3DFfxtDk61q/W9hhq6vlNKBMCet8rkBlpYK5ULuIby032I3qCdkxcti
dbWmy1K8OPUbhl28sDyASe3YP6e8QD0pKPVax2L5axQ1db0FlXcbpEV4hz2coa8Z
r8iafpXmttysHgR4lMTwHvUY8IeRpUTF2L2rnM4GVNnWkfT/hOSMgn6MADdGClY/
W5w8k+YxH9+IkMbAsN10sVHTHD+nYO4ZCY1/2QBBoXoOrpR5TIlfYpIgFLqPPuvl
oJI5pI2B3m1gUffMlEDmO0AMdK6+eBMEB+H8tVbWfyrMJx4dUkUPt240CB8LAQLF
QZEFWrZDEa0BpmDQbfi7OhQ368Q6BAgT9KvNh8DaeCY8XroBcce3AcaHIAzBVcuT
/a2bXjnNhTecfk40fz2ZfOXQeK4JeSAWqQbY8sO3FNuVbvVbp+Us/cyGsxvBucTY
dM+C3tQXbK92cV5F/p5Hvt1rTedNHsF6u7q6Ex7ylGJDIAE5GNgWVbtDLUzamIKI
EjahJuvPqrvwIPbC9GS6M39+LBYSRrICbvfLWNRecMqJ8KeEVCR8FfKbH+NZmuee
Y2xyJu9BfW8jC57geU2l9avMHsf6PRV0/15dUuUWZNZEi634vkJvbShl9F81b0FN
wn/HEQ8Bo8ZRhQtxgGiU5+d5tdAeMO75oy9C+Qeiilc38/lTe5YyaxgFABSXRGFf
/HG9zi97PC8Gv+KjvlTRAusIls0mFPySV9l27OuDq1fYvMyXueFHihRSOnp6+0kw
fqLV55n7YalkKdUd8M6UScTflGTknpV2/wADZ522/me+nCuyYlWON43BCfAWVkw5
H/79Nuq5sZ45uDC7UJ0Odtd47JP47buKioI/uSAA5bFbeABrv8Zc9sT+o9wgBChh
aOYEUw5X708y5xzNFIObAo0uyOfAetBlEhzpAjy8g32+8/EqOQRuG72374jlF6pi
1/GEojaeq+Hzsd+j/MZKgqqA9/Uhrvm+HeWl8O6BXM3Sy70GU9cL7HJr8pWRIy6p
78abMucl37FYfP36Nri8Rz01PtmHCcj3C+bsNOMQAzMh7slPiUrVaAQ88xbzd3Yb
lZMUBGXUgkmk1eoZXl9XHgxOBlaMcROW3TA47DztUGD1FQcSS9gfRAkeJncu/PAg
YjRfm2lfFJR0547cDAFH/eoVJqxP0i7yGmLR04p9x67UnKnqV6lUC+5a6qUVGaXf
5gzVGfO4IJOHEmf8JTyvFE3TxJKXViL5Qpnl2yIHe3ivRVgufhRYLMOtYRxPjKDa
zdRQbkkpP3ufm7dE0dOlYe5ieDj5sLlbPuxJPdEqjQ/2t3d35Ji5mkDG+jTS/XTV
pXnKY9eVoBEBy5ikOpSkpn0HfpiIrkyVN4wmlLH3Mw61utp+pvts0V4QTg+H18Sw
6VIwh/hLpkceiavThUe8yPtFntGyJpR8KNK5SLaHdIKq/1sHC5/Q9COgsY8O5Oiz
ObuWCVFKBe18JTOzkB/aBQGcaQzhRE2x37Ir8stcRtnj8g/VumdWb2z/rDpOHfcD
p9iuGk+GmrTy/MG0WQLD2OfhPcVVZ12ZgPTmiPi8LUgBNtpTyAIQCCWjvmuKgpDI
5nstiT9xIVyqfZ3chgUp/tTiqlo3wbcq+PjuJT1FlxeqO5jEUOs/4S7YEL3/Jnfh
+Z3gDbaMu6GsjfDrtUiDH4uT642OWLBnoVXzG+nN9/bIRuHHfVRT3ya+ia7dt+pD
7tQf5zyAEx28+FoH8fFpGLX9d7AOasalBTz4stgjwlaOk8Y/W4WimvIQkWa4GhXY
L7tj/uAA1NznRzw/Utl74KAmkVYTeYCikxJs2Bok8b2Zyo4rTD6N7HiSXTyoMyqZ
bHrT6OYcvKTfUnHktFMNltVtOlaNLx2dZrxlwXUzlDY0i38CVAIuoyuqTjwU7wcF
LP7gFg4mZSZKQSlMekep1mSg4RpDr0JgY1udlF0xt1vCR5O98FdWEVZ+VyAXMNO2
RSLg1yl+OEUDpUQ5gFGvKM8LDeu3tKdNg9cWjPaId0O+5I+oIKOPAxe08ppasDCm
G1huwGrNkstQLWJ+YsDqlgrvMdysGGhQV8BWiP3/xoiwqgKlnEg+e0h4DC7i8a+3
IF+04zoq3X3pnHMIIHBV0R/9a3yPakXntWsz2hfAX6XPpF8WOVNprYIYtVoKMBxQ
XsmunDGeS9emXoWI9ILctInSTA71VsDZ5q8S4FkUsSJp89xT33LpA9AjQ2b8t+Uu
G/Qcu2ei2LYGHC8hbuYreI09v6PHXNcukU9onK6NsxPvy5dytIPVNIq23WLSRDbC
rHJixG2EQ4w2m21itxH10+J7uy2wPU/w8vNyB2ri2DusQ913jxCLg2Hf12xOQM2p
wCRUIItLUCHnJcQztLg/JZpvextMRRiVNwM/upleax7Gz+MNnGtxijtaFtApRz4P
QBn4JeWxwX1U1IZbYKQSQr4NsT3zgU8EiSguL7b/YelF9709TuH7UzVvv7Mxyoos
CyAaTY5sqWS22u+G37zNIEuhJ5thJyg+z4xQKxhzNotg48Iw9iNQNwA8VnFaryUD
SzNKMigR0NJPtminW3jElXndY194KHuNb3lcaz1m1dfEpBvin5F7mmkgnKd2Xfpu
1Rd3hx2wo9BeK5m39Eat9SNZz2lBZUtm8b9qtDzh1JQ+9fPW092dz2TYHIkL59fw
j+aXcqp9D2My/UdhJotmYSDA8rGr+bLm2wgFQWMx7MVTAGkeW5sZXf4IV/VK7Qbg
ueXnKOYYYShyooQ4R6j2gb9CwY5HbvM56l5skkhPh7S5Izb8oFQZxH49dhSwX4Qd
LfHAT4UHYtD4lP6/YSYzGxLd7yl/yUPO0dCoBc6FQQgNzTs5EFPRiNdeiFypy9rh
Nro6fFmmt5ZMdMXudX6GtPx5x/0Q+CgDlQiKnMx+VWsBWDQo97OXi+MqkaY+7T5+
F2RpU3L3avs3cEAfDdaIm6zzVgw4i9qgDUj0cHDG/vPwRZiga1HWT6IB7x1TyXdY
eK3wA6DyyrJ0/z/HCiGPW/c+pJVzku0TMre2dZiyEUWWpeR/FKolO9x13l0Cu8u9
b4/TH5DaaD1rtFueQdRee5edJtc25Y/rirODlw/Dz+3rdA5lg50wq2llHovATUc7
GN9uTDs7Dszz/KH/rUJDREg2QaSo8tGbQuN45mFnO2DRIa2c0vOqKz/apjxehraw
P79nT31qcMB14xlLGV/UahR7OYZSvlCfBxF1UmzBobsJrxlGtU26oIO6SpwN9vYD
Z0V7pfSGQToT9FMzXJG3Maxv+9QT6DzjXU9REzac5QekqMQUAe5NepjKZELtFw5P
WqGLojmLc8DLJTj3YkdaeDcZTw4DFabjTlm+WeDAudoMXFi/NAczYMPUIy3GoT3S
4I5E9DGV7t5wYrwsiD2EaMH/sMfXZPoy04o4WKfSYWKqxIcAN3RXgYNk4wIggGg3
9pP9z5VmyxFIMlGeOPq7j7nroovTpO0OfV+RinoNgLXPdZALK+Y3l2dlgqO93/Jc
w2stR5jsXtVJgYIkUYJAsERkk+Ebx7NamJiNh0H4sH7sc0zTKTSqN5lwTxnyx/5+
/9xfbPkUbrpbDLp+QRrJdwb6mprKlx/mvsW9NFevSRlFnPExsqYktF4NrtbTzK6x
avcgsJhKQB7OBKsJeK3NLTBDvOFQsWfCocppiLTZKyprtZTIQDrkdfOUOq7lxB9V
26MQZ06irVyh7jey7eixUckDFRdbpYIYw2bTkSugExAG0NolUT1hFvb1X9jj1M+g
GTbx94M5wwY255ki22bhEZEPSLKpkumV+KSkEFmwoe71FwPKjm0grIYsXEt98OLU
1e3be0QNyqOEhTBG9iZWbIt1rTWNYa7AAHFun9SDcXs32ekRyay+nR7KAcOXZmAU
lw+HuL2AU+wVe0snKV7Cc8M/jiFwgmniNZ2R0Zc32eaCRZVsMallueUBk1t3n5WH
E7+dIB6uxeFg1wIE93ufuHGBXJYrGuEMowjDu0jJZp04T5TgixxPRQZ/d6Ny1tf+
dhFPCEajhQbWBGVe54XZCW693/AjvEeQtvqhSqMARbVAayvmm2Nu6reL0G+z/4N7
E267pD3KehegalMQHDOLLeamM8bqV0C1kbyniG4DWlUXqYZVR3yD6iq7NfF5PCul
wC//OSmei8yVXBNyiBLI73QvL9aKCsE3DTComBFW1c72Qfd2UcIh8N2E3q7PGelS
OFFZoqGXWqPD1RJ+fAPmgGO2DeUKvwsIWo1Y6tvHVriFCFK36EYufQ/A85lc8pYh
L4i9fkzUBoBdrnP/8ivYdPzOW7yx1fVA8pfyw3SY8rhPiH3365C9k7bAdd+V9+ak
T/DdrY3Szi3dvB3nPZY4rpLaMCbYL4NqfU4zoS+KaCgDCOCsTyVx6RhkYmbe1d0r
5lneH+PbNbfwKc4fVEVGkWduW555NYlB7ZjwEm1aKB2a4n5WtzU//uJSyQb5rmPB
IQy38cDhYy2S/75LW0iguxOyYnA1QEvayE5Fv6FIEK8Sm/rEKcvmr4K2BYEC1Dol
PlFNZrbslS7pWxMlybN0uz0Ym9HLpVZdYTxMEG5kBivaJwoCmMsGAkneykibYE9z
+LJs7WhDRe9D3K75naODtUc1dpcahJQjFa7amre4xSuvSB+FuafxoM/grfmVCU82
ekl3o2aAn1VggjRPq5rmSheM0xuVLooHtvW3XiL3/EeYOlFJrZX3o5dFq5LVE3ck
hK3P9jHRp07ZM4FWPtZsGXmidrxsBZlmAu4Mk4vRAmekJ1yBui41UM0yy0lkNLE1
OPGOcG02YiArSdAJCvNEyr/Yp9q8ZY7M0w0v5p7foWPrDd5Nrly+QMugeeRK2xbp
AKF0xLssjbRBybuScr6UOT5cHZhsDL72TQiuiPq60nSJBmWLPeoJ5MsRhcI154Ll
/4LbZH2au/HI6H4jzrHMEdpsUBnqgamiCEnKkZQPJPpcg7g6myEQ/lo9MltTFlWr
wX9xmQIF6laUBf6vSTbOPVim7TiMdgTRJ/Bbvf/TPqhHQIvqQE70KdaGcHYRLYNc
d0MFC1TvvOgzxViOT+q0JjK+0n7zx8a47PkW28DULza50lXUKF32TqAswteVLjyK
tujYr0WHHGi/Qmc+KrChqb3wyA0JFrSafdfqIvKLVLQs+1oGCUGcK3iMGALKTuo4
eShX/09TV00kXRx/N+QGWGCp7C1+ccALT/5ThKnpLs3q0xAwsrsx15Ce0JD/r/Uy
56iDzuhHjVX+QSfsgHPG18XgYS7xFmcz96rySiSq1z0Tr8Jpj9hLwuzZNCtqHyZU
udE8S+xnw0XZu0rNXig15XpN9MeCSXS/sWnXS4jYGgvdYm0MKsICQtRMdxQgl/9D
cT8nQLRLMMEObC+sF75+6GW9yeTFg/n7QuvRKy7UNaPvjoNNgGbknMr2eH5OPSkD
kKRm4jGwXt1mXtWLi/sN7+Ic9U68zzaL1JkS0FcG8p8AdErHSotFEydJ4hSvHMtP
0tPLYudPCmt4G8lZEBQOxcnxOOg5uTQLCZjf5oHs3adOoPrheDcj+g9h0tA8Eb60
nRw9vTEGvL80vmLk0qEAmGFqs0OK59J/DblNixqPTC7A8TNGdcgIUmLNMqKrBqdD
K1PjOAUz56tOxI2gEeo8FxoHLAPWyzom7OJYiUhPkUTgoL9IO4K2WHyz4HOw+YIJ
3NbfmJMGA5s23YgiS4YPoub//SWMdoNDzzH6DTN2gRW/hGSHBKsTl4QI7DHKY+r7
7HDdfvgUv4gTv7nAFwZErgmtKaj+kYlFWAe4SUxYyuYn0m/uxaXi5vky9NWdqtRv
pjrM3pIJFM2q+4gPdzH7ImwWZvdni2cdU719cIK5c967z41f+YReLpDfXWgaNmYy
W7tAqq9dzHVFRKvabIZkIntB3BSwEp5JWR36BsPsnwVAfKEZkZvntxrSJRAcukaG
KkxzC4GiaboJ2c81/BTm5FQlcz3q6X93iys5qvaqdvmr+J/RGPQQ5Iz3be1Z0QSv
EtoOv8UIT9kZpfL/u0mg791YaaNFDBqqvHDx0BdLa3KyvySBKXVc8nwQuhQNNoDY
yQLs42w2nd3hxzDNRkLIa85lHj8xdWO6QWlnzXzX0G3NhxgaC8dhrVKCQIa7+KB+
5Zizf9LEypmtBiwuCMlvVFt83Tjruu74L6Hx4SiQB3O6itVw26s8hZKoIKJEQ36S
xgJGIG+NlbIjFwCyKnVMRnicTZi2BeLC30Gb34hYg/1Ai2e+cn/6KueS9IbzL/mC
JC7ImH7lTfW2qNyt38vFYHHc5fP1TTTDgnapS76Wa9sYnIBSjOTq7iEu9o+hfN6p
uM7+g5ZD/q2FXXbvAyksPRDQgZvh4vKN83XRzz6DnL8EUSgIq3EBITLbeFWh/fVW
QphSIf4ND9Up4KM/dA7xCScqbo0+fBt0UvW3bAdl+H6nVCaXP8NzKXz80bisrmbH
48eIdyE76epSIlViQj08S+EgxiQgqwTZ/7wSvXSeZ4tlULi25ZVbilE8ANQ3zysN
KwciKI0T6gxe/5yfbBSWW+IF/25uifvuBKFMuPcl9iVYLoT06ukbKkceJNajkKQK
tSehc7D62AiESPIfALzKblG7k5l82Io3P5CWuAfSrP/mBdliCthAnd1riC+hP71j
HNl1GkZkK2342zAkgLwCPFj9cYKV0DK1+gs3WBHFb66qnq5shEbKSM9zkRCd3iPv
znMS5/we5gYnv8/mDJMJHAa2F47rh2We4tc/g3PGzUpR73GhNQuyyx8AlkoYs6HV
dpj+U+GcXW2ESOV+zB5auPxHjABZtLmTBchuFnOMY4C9vNzGIQ4wuSVxK64DnDxT
iQ6VisdYB7q8CPxKOhVXsZbcyCy9YBg0wOG4h2VOCm1hQdn31DpbzMAyVn1Y/Xga
ff1d0E8Va4dWvkLolgAMZJWYyHog05iqsls9Hl+ELko1AfGJiraouyBy73y2V4r6
EfkNJQwoMUNZmXqanPxbw5iwNbP/YioCYkBIEh55DQ4JeXuRUlICiFE2jI8NZizC
UCw91C4i9UhYeAqit8uwXi/7gjQq7X6DUK/DeiY246fox5Xgh1YqM38n+EicRJgG
/9DUpI0VSHD5cZ17qUlF7znWAlo1OyPEL3oZ95s8cH5clmIXdAvpUouI/eH5KCY2
S9yBKfn/5/C/0hAakSX/SeLgPOnA9ILz67bQJd9ynGQSOOepfqBY3tzK/oi95SQe
asVKs1babgU0kvxLKSK1dyKUmi5c1mN41mUwZ+PW7kRw/D6I1tlUcKzqcBHuDtA6
PLFc4CPrIFq9frc5hpewoDAHqOHUxxMOBFWxI3GyQhS+Yya+Qwahnz40LjqSMHz6
Tu8K45h2ABrgiVhWR1AgEuoP8ERyBAbT/B9TPPKAeSFFwU82nEClzmV5jaAh2Aex
IYxGa/gCNqCBCJtLrVf5A9t7JFu9/U7zXh/Se7fGjCc5C64WomidKKhSvRmmAqy5
gTnDTpkfBDo3UgB7NMvCegaPWif4hs9SwA7Rea2anTJxACzjB0wrzSXBQJf+Phyr
PL7LD5IYB460PMoE57+f0EvgV85bbV6ABY1Mw/6uoebekthAypCqD9NkLeKiKevI
8j/5/HQCQy3V4LUYPXhoFXSBMwC1L/PcZplunNJ/OX6NuRnSVud7JPEj/1zqhe0P
vgNQH9p44Jr9wXEGDFYA/8IjlR2noHc6qSwZCXt7veoxWptRIdfTliAjAjuRKUZY
iUFM1KtUhGlymCr9/4CCYa8XQ5na5o/7sh7omEWXTuuaIKbszfFrx92eYaIPZNDN
9o8bWaLckoArnDiW3z23sc7k7gkKYwtN/qeUU3GbierPUN8wI1f2jig59AxJUqBA
UkLkJYtaHMRCA/5Mdu3zu3Np2a6zr9LV0sb6nACl49EpcQCx2EJIkbJVY+7SDVQ8
djn5h8LZcSlK8lxR1SgsPmyzB0ADu/GUy2bMPgaFkwQB/AIdx6eiyb9yL31P7uFI
n63/NEeFyJb7L/C+PppsZvEn4DcE8LlUUf6TQzelNj5qFOFZXfHpxsVr0SBUslJg
XBeBjmaaFYUbswRV/64Ik9No/I0w6czHne68F+ut860KJpdAjWX6Wb0cFSynYJUZ
4aItDo32h7IDQj3mtiRLn9p+erd4qz/BsUhfSvHMjUIELedDusM8GJN+3CBHXkcp
Ab9uS1LRQWZaVoXq6ZHn+eZj4D9cDhJdKQifr06rI+nQ/l2RCEmtuAAiTa7LKfZC
ypV5juAmdeXvbO8IIZbcAjrDzt4pdP20qYOptl6jNviP9Z4nTK+m25VvDs/KmOfh
eSivU+pREKL1yScme7+Mwi3/tMjZW7SC2d5JWgJIv0wnToUm3Y7IBVfKfGOoUDi8
SeDNDTo2hVclRVqN0KmB3w1yJuGqSJOjl1N6SZE0JaM+9L4+7cmHCXYeAx8+qs/B
hWON+IdOI9JccoQQpgQ3twuXt69B89FsqkR7uaVJH6bAowl+jzl7VOV9Ihf5/r4V
ANGj0xWy10DBy37efXvfcFNZFcdNb27/3neo38uEUl5TNKcELgx5GUT2bYIepDq5
vhf5yW5XEARj/vk+iyP0gcmrw4FWKVtTNhh/7HZL6hjFhYsFVgYWCbQWIg2Vjv9a
SL0WsRSgNpDwug+PT6WB226GVCKozCvsYAbl8uPIFFtHtqXGz7QAsCgEZ2umC6cU
yq1gUvK/pE3BirHAtuQBEaW/LaSUyJoQ/rn3Z1TZXB7hgtnAe41C2riMELNFC7yM
N2PzejztCekq+zZ1TR7Wdx7LSGzPPOxNOcONYojnpXlOt1H/hu0IIVb9EO1s87AF
L4gu9JRD/4i2tTnh2CSlqCn2nuk/TVs9cWha8yYFynikwEDpimL+eDj61j1eEkS4
yPyGpouG7WTWQ+Cpqr+6309DWKDJOFKaTLTIBW1SEE0HrATyKQKsUfH/ZHQNFzBF
/QNWF6Vl/pMd5RcU0j95E1KXcaHieNI5kCodaErjjgMDa7/L3HiE5t87WCRBVCj3
X0zEIy50L0TqZ6fzGvtnEmRHUXYD33mz3zLt+50nMTNrp9XMJxFrw9OV0Z/saZdZ
aUqGZiB4J4EUbU+E7bd7CriS7so1pBpSUU2CqN5pWL1kRP/Xt4Cg4NB6UaNNdEgZ
5I2Voi6sesgqUbi7rL6+U8C6MR3XfNfzbygtjlFWEoRObno3bI8hm4QSeuODBE8q
9pMb1RQOxAjxjhzKxJ5ugpRzPuYOWbMmiApEUhfSkjUGz31mwo02Nl9h6QJYJ1L5
v7RZqp7IMuzNF0GmO1ymvbhvynyIQqGTq2kn/ujPlaJmc/P9MTWRxonvrZBLyxHR
z9nALFduSBVPqu5s1xr721ALhaXS2amqoPlxktGu3wAaxWUcX6An57wDrFJlUjjI
CtG2EAlUnTaPFDBJdb0nTVL+lYeCo/AOYDpT58TGyWkYDxOOi+fSE1vfI5uNOch+
Bq1td+ZXxSNA0kQwnQrtZ6geuP/Szzy58MUqKqnT1/D2zmzAEZqWahy80CEhaGqV
9ooyk2MSzarMREcxeoEnj58gy+KPe/CYVL28hgBgQ3XP8suL3/lR5AtXCmpOFSiW
kInOx0PIMxUMWFesMOCaL0yo06cZ6bmOhJltT+78ZQBUNoFRgZ5UlY4fMAlDCy0Q
PaU1p3f5e79oIu1kKOydQprvNFD9L9LzG0tiV1KH1Q6S1IeYEm9XKg2aXjiHyc9Z
vv1pdPZe4vfeDuCsRh4xGCUxi1P8vBkzhcCGFLO5kxaREZHlkbjPL4TRcmPhl8Bn
BfVEbOzOiRqEvSl596J555pVfLeVacBkXqfDBUEtEoYnc44ITHP9Vnyqh+IThMMe
mJEmQgoWqLWuXkhptDK7WCzQMvI3F5po0idXbIGnPvTkWVKYuaGs2kO1ZoRIdQ4R
zKNb7WzgoeIt+FasvaUSneJLaBC9GWiJNjDE9ZbDsOSAHtmp2C0f4YciRGwun1Li
VvzYJ7NkXBLjmunIP/UT3eMDbc/VPNCKnh/dknn2zAQxS3xz1Unyll0yd41OE5ZR
+arxfSM/DR7rtTnwLXtNdT4xiFth31Ga+we1q5+xt6M8bKA/XylbFiTDYaQT9lKb
mj7/TjoWfl7kZqFAfHTZ0hoPoo+1BYNfsh6HTtdiuC10xY/zp3zFk+Ev3ubop5Nu
b+D1z667qLrluQVdkrmTYtWmuB2+YzQe/4XK79CBOfeCwEulSeZCUkis2s9harp7
sJl33ZuKa6V8cMbiJbNPA2kv5p9LSvjQfjPDh57RFZx5S2u1E2PKHAP5uvhUsuAl
4r2GVt0R/uvjBva4Rba3jWmbNdY4a+EBFYoJOY0TNFaoxpd76eW5Hb+rxrtr7/OU
MesLLn1+SJR62j4M9rhvaX2sKtli1FcAOAIeRAe/y7gXCBPzBZkQ31mMseH0eH0L
oFSfjlu4g34fJbGfzg/W2lIeUkvXjQB1zJWna7bErKdRemWX/FyDTxVzNmcvdOxK
lzGIq4lV8I5jQbHl8LOE+UjP94PGP/f3BfhZqJuz6iSnHskWB4M+oUdvDdpvzgHx
9kwbkrbgzArBkMRmdab9ZgLG2DIzUxKsNEkGBjzSCHZiIOr2OuoyfRtNtK9YCh4c
8mVHXGwahcR+hmfhcUKcTJEwBFXX08xvnzsmrI82c3do3eVjdNl/asEbe2u94W/f
mx8k3t8wYyXOV0QoVfHAGRBe0TeifShJQP8I8tBgNqZU6LnDtUKwHyPbSZVz/U1i
4BRTQOHxrrffSozXnmtJrVPQPDS1qLzvubjDsmIoa2IN+7jkNYtFstAszTd/EvR/
58QD53hhAyZzL0u4oL10iZ9j33oUwoeAhhZvzfypJNQZpe7UqWPRr1s1o2ApNkCc
3QtrJb2APR7zul5W0aN1ruluWHFoQp2OIPns+WHFLlxlo8y0Uws9wldIwvWTp4sj
6ILJ4jEizARBiTXk1FzeKWUYXEU3HFVKN5ErZZA0EiGWyeGLyCnMEhXU42LYFL9X
i09bOy0Ps5qE/yP3H+sFRerphFLQKRCTVO0WciFsOXnn4G4DcYb47a+daOVV2nUN
XlPn+9eyXHG6K41sM23PIKglQ4VPisy92NHCNI5e49hKCbjNQddL+QFRdoXmWJ9D
VMM8TGA2WK/OHfDnVWao4fZ792o+ZF9+i0szgIT4EN35GSHDOQh8KO4sE9QGMso9
aq1olxFh6BmzG1yC4F56fVbEd2AF/PcnMID4HDeXCR14oLkieA3OOWoSxTxqBht3
ZSB7X3h4U5eV5nHzynqaSkVm5nU3pXWU/h7gSDXgF9ddN0CZktAZPJst/yRxJRvh
U5O8AQvW4h7zzKlmbPyvsPqcGDX8tUitBdeEztW5NFYjYdgmATSCiMvNgclrPBZp
H4xcV0f2lDIlgnhEeEv6juA4tZl/GkWlr1APp8gQSW12s6RhNGgWaVVnImQR/1SJ
DCSewDmaKGQGU7fgddKfvemzjsAZ44VA7H31eMnD1Qm3ZnEqhSEKq1D3oto7xE26
/orSXoN4fpZWpauHq4PrWbdWoCjPRxzri3Zqcsv0JqvQ3nV6SSIVkpv7FVBUkko2
Gh2IcHlASGnscKuguWMJwajVY7IEdzIiiXrYl1YrhHDBjzKU9K2PYX3HmFSCRC8Y
6NC2qUhQ+0g6bpMfsWfgODdX0sP7y2w/dU2LEVL14iWh21ARQh2MV+Cy22BrUyap
RgOlce5r9gjlhYshe2I1WY2cyGsIAAx6uwP7Hsg0YmCNfDOI8Uyn8XRcwp7ReT+6
bsj6Hf/ZOm8i+oEytQ50eg5cteGwoicmFQNJsOP4SzalD+79wLKdwZbdvEPnK8te
V/Ca3/bHh2zCX1F5sQTKEykx3eQjYmbmFE7GhB4cW9oSLr+lctQqogwE0cPEwTV6
8lP+62pNN9isEWCCeFdGmEcnE6Z5emQaFWOgucAAN28VafrKYROjBGQySuA9QWyC
z4F8VpFVmGyv2cqgESiX3h6UPVkLtExAntYB2fgnKmbQPDcxD2i70lVbEJPjUWy4
71U1NvXuNXdrQLIxUWMNafeCyCZgsRYZ5qzcyYOEomSm+qHlKBbOSHjYe74NQ7nW
KRGspE9qnjvPH8ZZQASdYLGnkysc1e7qgVWQup7xq5LWrZ9iY7zT9MjWizEkVmb8
i4JT2B1HiI+6KoKXBYScr6zayK7UF3UVeEMXv7Rjxx1KDVrWVaD/GwRWf2wNLOsZ
1l+RX+Fl8LiDDCkuaHzq+OzWPvlzW5d9GNA1bj5bC+osNXR9eAbsCGkT5Wg6xZR+
bw1rQil11eye1bZ3EPS2A+5i9lN88k8+ScG60ob8KidWT9jUoTvhsY+Mhnm+ewvT
7jxyzzVK5Db0iDizEMO1J3iXeGK0/IvwU1J5TSw/di5qiF64MUH3ynZbbK/K6TH1
6wvW33HkDMVnKXbyZem7trSsHMFh7wgYEa1JgNZSEpUNYWWibqfCokxbTDrn3I3y
ZSAvca1Z+9MBQIp8Z2r0dyZhsEsMiuY1NBX29vCjhw81eknXnG70WxigbJLm6Fof
12VjBzMNTju7k7hWyiy9SUoKv0Dzgx3vWq8PoP2BLWGqB9WIOno8UyE2QMkVXwXz
azlG2Ysbl/VbBFQWeWqGDQ3QLm/Y+Q+H5OZnNvCFBCkQoFG5lHn1LOKdC06vW9MQ
A9cVlkmR/2A1KsfN6h/yTK0sz7ubYCGxHLuSKPKc1rziJOO6msBPt9hSnCp/Qb0e
LOlG23N+5hmsm2M9nRv5ePcNWfJ/iyxPjuryVsUpJmxQk1yzHzLoY5cLOcbXYkFH
M1xeU2AMTS18CG6ALPVuKC7eo5UuJABsRrqvKn8x8pGnQ83iJr4mw+EIHc1z7xsv
BRIjUdy3CtJ+TMna2KIsIMdYnK6ImhqmLHRd8yUZmQ/i+eevdIsiRkPw5zfDWQId
0VWgGIdG9q3jo+9b4ZcXsg4ZMYCMlm0tikDNLxIxjYLelhku+tc3mcL3mn0p0/sD
TffJ56N2ue2HE1yCc5Dk5FQwl/mWrC7P3Fb1bUYVY0P2Hg9BF676wTyWqrVLKhin
Jttsit0FgPU3fZYrL5kEN0S/NROYhukgLO+Tkt9Tvxy+BC4d+QqNYqlkLU8VNdEu
sLFbKskK3y1XH7rZmXFWfuNyql7JZXHIH81CP00hbnrkn9PUcFoaJRAcW9nL/CYq
AOPzxHmWTjh1RFTDiZ2j21OtsB8vZ6yDQ7xKQmSCkGrqBbi8d9pqDH9qIOq0JBRN
AM9gkIYyURjYwTbfPV7sU2TCWcFaupS0TWlGfRnuBa4Gke+JC6qm/MV/HjZ7dXtA
c/l3Sl5oAv8VVME7zAYsAnHQPSSHVZfRl1q3/sYxce8CkVNlA4q5XQn5IG5dVY1s
tXHqCtGWUh+E3HaVkuKs0QMoMxt4MtWwIKZr+jOOL6DSxpOS1Xuv/XuuoVcO/M8a
ZY8Zw/qQZ2WAlXAKSOoh/jrFfOCLjWFLx6TIQdyI12UP/bVlbL45Aru6VjVyO6Id
fQFVmCCiugBZ4r9hYDBYHELpdfDk/1HrMNEnUYj25g/w7IRzMiTVIHmMZC1FGRZ1
rhfJ6tMyIzGaS1vmQ8iEm8FHVQewWMX8tw+7IP2vpMP9WmLryBQylxP1kFMiDrn5
UrsC+22mpWt8XzrkBGvT2IUwGrQ0oVbz0UwiVAIJ+3iOWP1xY6FyEuekZskF0ZAr
d40NuO+mU724K4bOX7Tb/GY7/qjMkzFDcFA/RwDFyBzip0/HeCgaYuFuOHL2DJuz
togRMc68FEflS6iIymAVTfitfMBTksPYPfllZE6SZTgxrRmRYvDW236RTgfj3Jp7
9hOg4Xq/SVGVRKFBosdnySyzI6mc9SR2P6hsobWapwd56BM6C50raKW1hOXOp+gO
XlUR4etxmqb1rgzwczb4iDdY7nJma0cI6CfTXRyE2I3PetbIZ8tytZpZPqNPabuK
tunzg9h3QMy5wPqS6++RduvDkhBbbZsleL0py9GkGdwCTODIsszKInb5K+2eICj/
8NMUmjgAw9yLjU+xSGrIwQ0OLvqmTTW98sjYajNphxDI7KC0KZprrJ3VApVxzpu8
0+lui2lTJaQQiaOHbd3rzuM1CZYLnxqz+ENlcqbkURFY7bJmDrObxrJgNb4PVkll
HAhIOIQxH1oSzppYHRFV61DFE3DOaHMpenvdRJ2EqKehRRmpWrv3jCWFcwlaH9DZ
E5xZKTLlY96J1HJptb0CrhrtH/Jt9XhhJ8vR08ZsxrrRfIjyY5pzonW8dbVfnrw7
n5ebENCMIqzJ65vsnkcqdAAy9WVoIWIU0Koh/PQx30Uog/4/Av1CMSajiReSXNcV
Ph3bhq8Q8oW0hDS/MRi19e74XHl3oC/WLrZ/0AzKeykJkf154iZ6hLlSAsd66NAN
q9FVCgjOynYGsSSCDH+lyJ7rBf0v1G6Y+0JP/klcC4LNi113MB9t6sdL1i11BTlC
zzu+VThoAP2m06LIxnyFVDztwaMb/AJ7K7KvCE69oxDKVL8R/T5z6hD9oYBN/tk7
s8yhv6bKHi2MYTZPmh0QFx/h82I/lV9VsGvHUEsiy0iqm62VWUKLMOS49kO13GQd
ePJyRf+gLpLVS78HErFxThITZcccYgIh4c+lhSAQyqOrVjzb167FvTNVx9bB1OHA
eGmAGdCLAG5jy7uURFHdaQ5mbyVfPDkTYoDEUcpRBc26L+Za4zhlYM+xnIXBbiHG
2mQAtVtSEl4UhfCoV7IG+kxLQAue6xFLXZwmgmV0IwH8uyqWGySHzWgaSQ3d0QKM
ID9L+mlCDGdFDE9OmAcaTvkX0RcMJJIc70yzAtuHmEFFPeROcwSzfUy6mNpbw869
K39EAXFdOsKPqFj/hFO7Gf5/tOSk3KsytycBxZ0D/FdGOpxuzhjaRjmdqzcjB0dP
9v1L1Uo4FGIO41ahiW1EyEi2idcd7YzkcjuEc+bCuwCF1msqnyGjinxD26gwdeOj
sqE+S0mda1qXZ7jE2KlOvvrGA1nZfWeiLwg4EZfz1EGeRNbR37wloSIlwucUWHPg
QQcERG0LSwgvF9Dp6iV4/idwUYbg/6iQJMXGVA4PBSR0kzg7GOxp+zotwrXfjQXR
s5vv1CmwXObaPYHu+nQ3/xI9LjNZD1XjGD0gI+Vso5nH7xZqQvr1jfA3VHTADs7+
smouAAhVDAByL7jcx4oX9SZ0J9joxA/BNZsZuWtSI00P9FxI/vwd+Roekr3r5J+s
QxafmBQHi+yhB+bJnL4asNKnPfereRwxHyg23vEsR/EydJTHdtTl572iGp6nXhlf
HQdiVNWuSInQCM53Ac5TEOxu1FCs0oIr8VnX1vUvZNM=
`pragma protect end_protected
