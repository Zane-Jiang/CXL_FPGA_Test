// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hZeZBNAJcn5o+HBGPM1sLAMJiFWulvcf5nrcibXWYTaiZ1i41lVCrDagO8ab
gUgmmCBEttbO22Hrlh5y9Kv4YCKbe9QaXFa96IWUWo8Sw4fRkcUlOxePlVvn
fYghJafyw5CK0FFV6o8G7dNS/HJLEN9Mwg+touXFivmSY/wB0og9w6n6Uist
YCY/qnAkHQoPeNwCsdCCDAK8a/Hwh4svrQgpMfX8b/JROb1A/QbQfMWljfID
QqMRRuTXkX5MpGoVO5wuLgOYnYLDlA6nUnpXSKKBspmdGbl7Kev0+N2ge3bM
yC7U7jhTH3ViTXaBn4jLd4PryrWgLXwD1iXmfzbTZg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OxyDPNb3Qqg5v7M83NPV5U3C9WgSdmP4tPJt+IQzUpqV1MhfgRP8rba5bQJ6
A7PRqSs7cNjDjIWt6S3KAfnLiz0Vd4nEkAjAl9zQQrC8CD0rgnw2VLNt/1hV
Dl8WAAZDN//n7zbrjKizqsWp0Ss6XPVfD7Kyz+1e0cRHy5FpSebcfaIyxjdR
xIjQwsyQlE+nqrcAS0C2CEoR/PLehLqqg4JxJQ2SbESq467qiYgtiJ8RlHw7
06LNygAwoUa2gsyqUoaBnGjRh+gPAoMpwskswE9+obRuL6A1ZZLHR5h3Bv33
0Il2B9X8u1lizeexbncdhe7P4AAiL3jMOiShm9tjGg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VcYu1PTnVz9PoMXB30ZVmtC1Y+b/lcEMbjwcJoNAGxXSGHTEnSDcCYMSdu6n
BdPLi+ChnXO/7bZanz3TW3WWcVkHRk6uFNvFC25XrI0YNTClGs1LCys36YA8
MdV8ZawgXLTAvfhcdOylNLnTux7EK7g5cfaPQYLnUWUzGeLikMl0LCnr4dik
gbfRllbeXO/AymANYQsEn3sjI9PgbPDqVL7egiNQbIEUUWUmdZtHl1elEqPR
95zmBGvwroMF06Ay+yVHhDJvzIYnhU2Lb3nUhLntW1ipFi5My5tSwIsfnWNb
cCIf0SxW2FndaMxBT+Qtfj2+NNiQ0GEPB8+AN6cK9A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d4YhJ5w3gFvzR/xgiDshFWnjEkNxhd0ZKbsAu+5UmHJsXw1yx+eyhckdTryB
oFZpiI7pw5lWl9y4yvf/bgQW/zh8ZhnEXLtDXciNv7vDnbclCzz8RwS7PF18
v00ZbDRgEekHXYGCAPLg7d6eFmp8xJAaBkaI6sLwhmfFU2zl6yc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
H38kGfOhYNsiOqETxmWC+PBeKFKdtdIKr8P9wRVHPBVb0YjNBm1m04Hq5bzZ
PwNgQ2U5EsNLfFUeDqZIL8jyGKTQ6VYTqWnZnc+c8Qm/lCyOlGgTupPsVI0s
81lsSB2GEk0SR8evp7O5fw5BywEUfc2GvVOAihjAZdqCnzsE6tDQAHXLCqxz
HfuGKYjvqDP7P9UIlVwh8l/iPm8ovz+TGkLLLrkiJyaG+TNs930jQA6W2/sx
qyL2Pj0yrtLRep6WXIsjlOw4lPTnT1h/NuRt/dbKl8pbO0GGEGYmN/9ox4fl
aORHnQ6f3BnCwfFkY8EKW/3j4ZSoJ/a3jk3LyGHjMSTlCyHP8VBKObkCTX9n
DJtvpMeldarBkLpOvA6MBly7cepVpB/A6koVJJhRFqijKyahrVTbIih/WVKH
BjgcimoUXax5Ql8ZQFPQ7zD3b7RKgMl9KWfIFFzR0Tbr2sefOX1reiF2c0vt
i0tt7Yuv8jtDeiZSA8iDDMIXYUd/OSpF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
geXrulwrqoK0glnwO62GO2gZSyKQlJsi7OUeRpOuEYpyievCf/DRqpBeuvN1
7eWMGm4FP+BvH1SHEC4BJoHPOk4Uck1K3G1j5h8saFA2koeb+G5U9Gidqa+h
xe9z4oMPwQWzn0jnjAuNx2ALd12FAY2tfebWWsY+8Er6RT6K3wU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VIho+PhxlzlmMhY5J+G1hj7iPELRFjJaUiHgWbZv8ynJRvCK07HCKn7vv3yX
m5yuXU1mUX+9anJ4IMEWR8EYEPGxauq46cGPqULbVXa6wxxiNa/B1xaWHS4O
4XDQKhvJRbqkaSLrZQw3JL/BrxJQF3kjB3VpYfmOfB7i62M1rA8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1152)
`pragma protect data_block
R238LVr8XeCaI46adoW5KakHuZjsgOM3+IuHuCmF8wFy8+P60Nr+pN+FIyX4
kvMDpedo9aiRHU/sGQrA6yKoQGubR8oCQ+8LHNM6+PS0BkIpAWAda1pr2ki9
nYUyTRjRSBuT94/PmsfVa7xAY1lAc+O2yCVmwW3PSNrY/gbhOpuTTFXlrbg8
LJJ5IAcKrw3+BJepuDLKXw/I8G9jF6qeK0zaZVLrQ7NOwKvLosMzxvD/ztlO
idIeb7lzg8AdKDUZvzQ4e/7VR4HdcxtCudI2O0WabCTLyX+LHc1fwPoOIp4F
Mxam4gygKfwL8Vl3RzPCsKwAmERkZgNWEbI9BzDnpodEjNit5H1K4nCcOPOX
AIBrHGJtjCS1qR/T/Z8MsqoSVcf3NYZz1amPUyrdDreD0+Hqn1mtsXhmm3yo
4IbQtOm1/tz7TXnFk46965LyPIQPbKGUWqRcGycKNw1JHnBxYQJWPtguDgar
3W4dd9zNvaIfp1kHdFWyvZtpdD45dWaK9lXUtQEvvtZMu5ik9/aYl1Bp4Ka9
1NOJG0k6w/3bmZDa8Ko2zJVSFHxsxfKUPEzev7Ya4lsQZ+HKyZ+5AK3nHYE6
t70eE81Lg+FEA6QNW6coBzoMicIjBsfQjVl6NjTMysEC3yW5FkrhCUWjSC/6
OpOOIg+90OVVe/baZh2LYsJmQYdmYoAIWUXC160v7A8cNlyVTtU94dlZzJUy
YFGxi52RUwj2uBssu6Frnebal4VDPCiR+s3+f0bvRHK2+mW8pVazkLXY2wqo
vXz/McMqoUNtV+sdzwWoGdZMNvrPzbm3r8pYN0L4xw3MwXLYVQpELsO7TbbD
4kWIiXPncDJ+DePixVbd6tRpAfgtHINxwFFJMi/U0VA/Q6nCcRXGTzvrIYRQ
lfrzqek73ntVwvqrxQNF6hjntci8ntYf7YmWEbHMaOmToWdicjATju9qcFFV
+k6VTuHNhbebkVZjVZ34hbBbjDzBxqjDUDo3+9L4x20XtrkrzqrKBe4j0THl
o+/0ZVWIGuVB9RI7d/sCkfX7jny3thRnpD6/iskDD+qhJ7FjIQp8cMvTKx6G
45FKt/lQUEqjh+m60AVb2M2NgxOBfWTP9exorfwRjg91A7hbOwXsv2I3GBFD
tZmb4UkYDl5FafXxe2rSpuZXEfwMnQlBTEA4d9PaMYeyFc+3NW4xNMP4x0+C
fD3YojyUjm+vUw0t1A5vc4ZacPcu22rt33J3wBfIChXTGX4f0JldGDCdJt+L
c8Cdh2m85CdvvgfzVd8W0mc6hKRCIJbLzKiAjlNabFUwvAzCIs1UBbCaDpSB
FXZenfQnRqYHNlConJzGULpB67jS6qtw77ZX7FzptHwYUOA1bkLDijLplMI/
QBTLthhxyBPxcscYm9m9uUjqYd6dfxlkNCUxTYvcQpvY/cgkacinZILWHLKj
WzU0epTXo3WJwxZGtvhNIFjituZg10if5IQlrOVLwEQS5LFcTeKxsbjjkqKZ
VPyaQIUKeMjHDqlypwQBpGVuHVnwPeA35DES

`pragma protect end_protected
