// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r8O4i4LxH/zvRCjpHVpOM2aikajSHcbStSLKmBF5pzLVW1oZlAkmfcbCDp6h
QzaFpBr3545/eQIzOniGHX8XqErFLd09JbsjQ0cDdqQ3+aqCNxKIdmS6yIBo
9Y8TVuZGul0CbPafnxv7R7/PmTZJJrrPspZfqPhygFJE/42InDf+N/R/NNkR
uQLpH/Tv2T9Iyq/wWmjVgYon59e+ItxqvSVDK7iSPqqcbKoYynlYmOH3bUcm
aLfhxXkC57ol0xJgy7nFAnIDlKyEevef7tgw1Ws70F7mqc+U6vMQ8U/6Xz+j
EXV2nnUKNhXesKk62657tCD4LkpLTPdi8CDhaMJFGA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BtPYlqErjgFb98W99/dwsqmlk4MCpGjvdOjt53osD09y2Fsg829xjRLx1BvD
m3wpr44Z0JxNiAXYT86smjV8a+Uz0b3sxdKXoxM7nePFIh259nPcsMT9ZQLi
expzkl4oCVarRPbE/S+wrPdWk15oWgbwyNRZt+O39HDD9gLl/9Gc7IjMcUEh
OvBOJAVx2IxRFX7Wbe8+O/GFJwGY415B3AAZyUmDhElnBD/MHQqIrx5N1J3d
U3oPVmGGnJryCSKh7PcS7A9ucCEPVuy+BOKBOHyX0S2JCY/gJAijCiTLjcHH
ZzlpQRNX6KPUqqx73/TwlcSvFBaov9ZKOljjcF9rIg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K9jJYBQg5szkTDbmai/Ms1jv118XM1ynQd5wqIsVfKF24LDwwtxkCR8jugS/
YZlzt/4SrTn+28lLjlGiOgwuBieoqpxd7Ymk62uvYBkFIB6BIFfpNRVlYsDX
R+uLUoGXdNTcFDlB6nHkEjTmxGMNQ48UDmENd5wCdo5+KwRy5rxVrReok5BW
zm05+jAWiq7exWv9lah5F6qlzv9gfZ5FOOf+b/QqzgR/efOneiEy03Ehw0bL
eO4M94E49QSdKYVhT9C9LGBdMtXqeYLxg1nJ/d8o70lkpXDrzbTw68h10G2h
+Imw7UC4IUq9wpkASwTUeRViayijX12VkNQc0h6bow==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nlh8vJyak0mj6eEu0o52g5Xvnhw3u7h8Ek1Q6jBbTmmDIQKpZdyOHmsJ38fV
2JmwLqbbtwUGbevlMPdUrbqZNbEoaevEWPmAVUjxIbLnY+U8cimwBDTNHW4T
QJHbuS3MJJsCuCnYIyyQKJ0fz/0Aw/pOg346v/U2fCDAwkQmi/g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SbkC+89H+jcfpNp1L9lRNY0Mqfn5gm9wqyYVUjFBwTRiTq+2jbQGOaz569s2
2toXUY6e1bzl0IN6lwiOsHPfC10zUq5b7Lfddxy8kjpAg8sbzfYrGhq5d6kn
NL///g/T10SddYguttQH1MsfWBUerddfSFwLmrafmXXcoahLNXIlvVcUwWfq
zD6dznBT+0n9EHjr2oSZp5JcmXb3c6wCIiX4+yTWDYT+y+JCAqg0hD8wS0yi
EYcdD2aKWp0mTXFnVhk0Ee393H2BT+6K7yW/87xMeVJSNsTKQYv/tZfikfQY
qSv4aBsB8k3M23CgxEwaxm58+TEbzFI7xpIPp8wAgQlBDu0rNP+By4J8dc6G
5t+EK3zRTQiuXWmhHwYBIyxmiJcF+VuhEcQuNnAjrEB254w9DQUdjUtzilIB
u7ySHLVWoJ4l+ZrZxPXaDLuUJ0skeCoNefXwksMgV7bH+ZQ3/hWcdCsUl+29
4Bu/nV+++x8PP8wLUzoj4UsN0y74z2im


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QIsWo5qvEXYkf4V9d/xklLINIa7sbhiQ4IwD3U+PoreIHKo8ocl3J9kQ9Dld
+xgS1gLP/NttRPqAPfQvETrPXc0RiLul/L07Vd4D4msmOZz19R8Wl3eThHdD
UxUlsLRt1qQfeAkF5oi2GmpY/znvBpYCQY3jsyCJGqf2zqTpnyY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DvqAIFFpS6lPMm1vHgSFUrmGFYoTM7OY1QRPjr6kYL+2bxhueHcQNaxUusY4
nvhE88rOBpsRQu3qZyn4qSuR3k1F2n7lIq8MAEuRZbEXzA8FBwdr7AaVQ4VZ
QvMokWRyxOnyCRcVfPT+ZEqR56TithihMxfHR6M2GIU/GcrBcwY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 421024)
`pragma protect data_block
q0E+si/FFBEANnXMTB0nf1ZXy2HcWxRe2GLpyAPpHuZk8xsq/yA0mo8V5BjJ
rI0+H0smQA6O0CM0QloK9KmTl4+iHuHaR2WnIo5c81zmZ/fvvebCcm7KudBJ
kuOA3feHW52eWKvNbIY446uwFWhgWF0jy6oKH4tDdohAnqZUBlEi/Db+wK7I
o0Y3z2eAB1rd78rqCP1dpU1uWgnbn2zG+yoxpQZgvoQcUHERsxZiYBwJwa+O
zqMFtMOZFNOCN9dBr33xaxwRxDxw8dondLB5AySFi9t0c71KZbvmS8T4yH5q
41/fc0Rrc7QuLaK3RgNgn6SbtMExst7mbgHLGfnfmK2KBt70LIeK6+aDzQsN
SI8FC+AUehvFa3AL6/qXm/MY11PYFKNol1YzI8+OlhMCuMJ6rS68M7JReWeH
RIOaT+pJD0IuvqkiJqsWVPHzMsLUGhQaZxbT9JkEFZXpjo8QgFudx2jSJDUb
rK0W0FvsuDHMdEe0x/53OUHrjjxVaj7B3kDFY0eaDd4P84An0zYj9E5Hy5lB
bGg3Dda/FObOnXjH5orKNlZdCTVw3Ewj+JxFymaZzsUIachR8hwYlFWVMzcz
aP1p/D2CZCeK+BoKQ9JIBkotbfXtxarJt4kMQomK5nRniRRrW58+B6tExknd
bwUygObOnUsXbpY4wK94uT/8rpD6gf51jDDf/3WlQ/RiXUXT3Le2RsHuRcaC
QvVz1QoNyCc9l0DfyqrSCkJ0ksON3aykObcwp3HmVjTsKd4OCK9UuH0PcNCA
xt7KmXMTEOec4BkhuyaJWKHKU45iJAA/Z8EfpkuSHNstu0TH6iqBMpJ7lRE4
u/g+7Y2IwO/sBzSUH/0gJ5u45WM1rkPwoAPUOEohG7hFfvzcTTAbxNNvm5fA
0cVBBtuJEWVEnafdRYgYFBi6SvQR97+w+hms6gNc9FJCbQJiOyG/ycwvF1iK
YL6k/ipmeMh5JsqnUl6yQpbkPZQDxDt+SCazGB2ySSgakqGDjaqt7fZYr8pX
g8ApeEfiJXgbJJ0WEodaKetHc0sUIqEE5Ooc5AarLUzaQ1zV4XKNRTLN5K//
InZStvXfvaO0kL16hbCXoP7TLwLeHFRY9742grghP0P7UdaPZyyOXTEx2z31
UnMVweM+GsU0G3imL8449/eFDMdRkL0h75L2d50zQW0fCSWw/3rAxglU2jfN
Pzn73wgoUo1xbNJgN1dGT7tKJvEXSO/Y0chXe15HK6nrb0HRGdyUjDFIoCej
UUMsU6ute6fl/EnYSLeSjNKaPUhmWuIPF2lQ561AqJ8/7Ve8P+0hkuhj7/WA
/fsQZRXxTS3OCCFRUHhbU2EUfHZdj6iTBR27OIVxekLXbrrH8Syhi4Acd6K1
d8gcceKURvW3L3WcMRld1NZNtzCk3c9yv8DZ+fKz3es8leVQfQXQ5XLJ7oPX
cYYTbANbRbXgkAV7+oVnRRtstF9tLq1HaSPEPOmZkckWDQqnMP1WNnIE7O3C
ucJM8dZQRjj7/82wm1thlT7k2cPlTloU09/wsfuRD+FiAN/U9wxjQwfS2swj
mX/JT+czMQ0M/r5Czs568jgODD5ayEc6jhAGFu1e1v1wx0sUzq+f4YDYTYmM
l/3f05IzF6NTUA9L1JWe4VbhsjjoOmZYW+WHY6iX/55+4oW64tG/GMibuJP9
88K/KX3bs/tLZUydCiNtzEvwpUibF3zLJ+++gjEbek0sE18mwrXWKK9aEksV
5CBaNrq29d27GfldgyagBLcJbWq2ievWatoKcTkb27q+VgEsklLyfs5nrwSM
owaPOrauc8JRp4HUngwCtXmo+9XIVlC+x5C+b3cojO0d4l99o6U1QqlXkyPt
ObDoqxzgljCHnWFvXqlMdztXaDbjf+GYmIifli4Ki3pSjgMzvdhTWKPdCX/R
mzEXZGjf9Fd7gFnK67QfxX/OemYO9oH4TTWZALDDb+JA1vaf2KLf39PnoMcw
Pzd/iIjR6ZrHtVImHjdOxbja14CjIDG7nJFHpbMt/NSJATa2/6mIwvONdOCf
eySisrhQtshJ+aAhUooj99PBLblsL/2nqqsvD5YutpaSmrUk4m048Gsp8Cva
rTemTsTk5zmFIl5Jd04kJ6KRg+enXcGuF0nfO7HIceZnhJROFJbLAvwcwS7D
5EpO9tR33J9vfQiZo1y1kOx+esARACllDYDRdgqlm6333xbE95HulhTmxW7W
VqpCyGv8o0JsnnwZtj+1gYq+hSJQNag4YsxGRmVJpPyZ3HQjvJs39zr8j8x6
z4FWQG6jOHbFRuKzIlRCYg4AoaLmK/PHbQQvhbJyvmRX9LkQk6fuC11tYSRM
o0VtL3XCbsV8qhe12p4LOVXfcu8oguczqijTT950TWC8gwQHDQSs9sETW3ng
xwLxyCiDGdd8Jc4YL8U7VNIvZ3La14ZcVULu658rppMAG1XFZZGCbct3WRdI
l31h+tdnnEe09kjrT+ef8AwywD3ZW6hNeyEctMarO2qfTCxlAGZOF9cBoWtC
ZpHmfKWX9ksBLL/ij/kylwhW31kjQ9BYY3gCNNjkA9Jh53wsoc2An4h4O5Oc
EulKpg3K3IG0OSnQ3GzVwenPwYsqep0IyKnezYtGhPy9JLJqMilJGEEgUDMq
1KTQZUosOugM7QCZUDwhJi40VCPyD9DAxcGkUehhCeMt3XhVRygFRzORNpEd
SmFvjJzB2NBl16ebOEWrU9hsGdF0G5YLqsRthG2YKlWrqEzLapoNZRQqhVJR
WRsEjse7d/t6SSEOoM3gFLJyNWeRDRe4UK8dpDn1FzE4ZXLAMGGVruDdYX6V
x0YaiPQT79/jl7rvOsEqcrwGAiRarDpyyVm+Hp6ETQzzmUS7/WMW1J3eFJJg
VOVYByctZ3XGsjS8wcCMSYoYN7QtOYWeRpScXteAPQCwuA8ySQIcPUKfovAq
Qn1L1rYbTQj8wOvha3rHnbX/KM4hnfB4kaQkHAEU87KzVGM63fAuwU27PZHQ
2P1pkZBuJ6d5H+Gkhkn4BK5T146vibJWJTlzthF5wCTdIhrAN243Ee7lJKJt
Td8wDeKdpEa2hWjS9a1k7JPHRwKFgAUp2Z5MaQzK590HT91sfxRU7UhCpEq/
vv6cASR+zscrGyT3kEau59IctrYW9fHDHqM01iwvyoqy6xDhta3CcHQMiQqy
9spGYseyKdA8LOsWzD4zbI3EUI9XWwqmr+WHOPyKM/9L/QK2E0RMI1OzSnKL
cNrnEpnroOvR6kG/GWQQk32+2qVGUabuEb7Okz5nET4Q9G45ftOGpmk1p/wx
4+hNsnHN3TCUfhnJGdd6NXhFTLjXBZnl4eTOxXP/L1HDGSeSnZOQGPdZ0mVo
/9VnKZWuVLHmAZ/lE8EUc8Gi5wRHsbJBL+6aiJn21G/fAJIiAEeTX36xtPxb
Zfc2pcQ2ETpyNGbFQeOs+nD5ZVde5c5xWjDGw33clihsWmuTWySew18mSI/Z
MY1MQOFoI2EJX8m1cMRPu8biJtcG5NdrXc20n5fpkH9rSOEwYEfE7YL31xzF
2oVxh6ZuvJeZCMPYZAlZe2ctvSInpfKH8ghHNyDzy1/R+sP50nrpSrTd6MhY
Bt2S8jMbj2msDhV3NIcZI3124qzdVV+1m+9XtS0o9waYxYgO9sJjedPugTGV
dDyEdxq4PWBc0mA4WGeNymRcPoWZ8JkyweIKi+SOdGUwaCJZjrD9K9WHa4TY
UBdYHH8mhAlPLaRizte61icV2EHb1JRL0oj/96Wox8ZrDNLrk+edY1KK7UJl
hKwTtwkNoml2lUH2giholYjSqJkXrxd1j64q1/2S9lk310t2itmOGOwSJfQt
duOrlw/+DK/1R3veBY5uqzRlFeUbJWwXgHflK0WnsxQZrrn5/VOgm7ckKtPt
piNWwzuqL7+DLRhzQIJJL1hwIDzLOnhdsBP/A3nk5+bRsxqCk+dt7tOZbJNN
X4ULZ8aNhMqZ1fGkuwNJxzlwqtDU8//c5runauYx+9Iy8WK9U+JkI0TqNI4O
bHVcnFOqMO8raXmt5GiZdAsMKOuFLt/43qawa2hgeRVxc37+i+XDv0BRrg3k
J6SNcbGSarx4SVBCC8HvJJionZrUtZ0wtv6dHEcYQotLEkpUJ5Aqz2nIdTHB
fuUNY95ZQa9ubGkpntaaDVXYgtRZWiu/SDX6mKh8jzktp+Z3eAiIkdtC+1wo
y5fSrg+unEz3mqnNqREPiGFADvZl93RkDYm6jtQipbVDnUIjYCIoJ1qm7zCt
eM226hzs/Tg4gqMNhPTKkj1H4m+QpbM5yRISQc1U4M3pK4XkttHQ0z+7OPqM
PKf4TrZebqYoBLm423TEHUSU3Jn0LLfGTZZH71EQzw8kHf+ehKm0TLtYCato
4rPkjrtmfHVUVFHuLL6hq40Hauf9bak/aLqbqV1JdZRchWwnG+yAU+wuA5oe
qwLvPIvOhOL8+aGE+bCY5WApdDAQ73NqjcEws1WcvUSHZiVIJp5Gv40bdh1F
mPfwhe0DmnNkf2+9IP37l8E8VekInirxb8+RerLCWbDCgyc4mHqjns9pmOf1
T33YIcgJk7fsc2h4Xtg4tdpl9fgEZkZT217e5W1MbaVCSp0L1JVmnfoInvGc
trNlcuvHFNz6bL4Ej53Vg8Qt0M5czj+HIN6ZjZlBTNi4eiEIyhbi0H9dL69y
WLuRHw/Ry60o9a5lnUXKYm7nxBtIkFaHi/WGG4YIpYnpfkLZudui+JZPz0fo
LESnaj0Mnk4Yq1+1pOJJwM/INLBAbKzpd/RR9WyZgObGCW7u+Kw+RctNGtka
6Ol+RPhnuUAo5XYqsgxYPhjUgf7R8kELRHd7wmChS4OuXRjz8XZOaGZnfqYL
XBQSwq1Tntu4u0gl6ciISQrPnCvfTejWZUoDdmYd5UJA7mIi0qEMMZS0bARX
BjU+f74hi0LtmfOb0s2G1zHgC6T9Rg/QZzzeyv3iE2geNSzGaJ0K37qMA4lw
FsGujD33l8eX87p0esEZLRecuBeEImAjkPyV/RPUvTA7CvF36L5gZX8/suyY
owPm822S7/HLRK5gGe17q2vDoKP0cp1ZwGI8eJM76dNOv5fSG6xmB0zQkFMO
zNP+oww5MJIWqnoNdkUVWSkWH6Rro+BLkHK3jhjhA7uG+in6h14BapngD0ju
y5+Mo1p4ZeKwmphrIvGtINady1EFAAyxabDT2DNxSs2YUUtat5Ol7piw8dBP
y7H0Apu3cUrL9Hz4yow9n60N99bTdlJgLsLDU2ZASMKkDo1lk/jVKv8CCySM
S0TLIW1wUsF3BIZWy/Awjh+Zrzb0hQ/hk3d3ANGYONxW0yRLYVjXCLJ+dR/5
ohkBCL9sacvI6zbExQJIbExcN6mHFT0rCK1bW35GCYEjk7OwihfKhgkXK8Az
WW8NTzZ/HU9isGkhvIYWtQqGAMHxmpN2l4iEpkU33BczFUYIMwt3QkeOZgGr
vTMU5s2RIN92XOXOl9hjw8bQM6vlfwFlaa/JqYdT5ar7kc9RSDwx+dv/62zM
ysvibc2PnP3zaWURo4VjSThmyqz1D8Ffb7caPxg4Zeko1XZtARMxJiNrxANi
M0vcK6vmNXzcy7feScLJOWa5fGoP7w/TVdz8UGjnO6IdKk7kuWk6Fp5UkDin
w20GdNgkBWvGB6gaxI0I+yGvPAIpe1Xps3Zr6HcgiF9ZaOY/oK44UM4tDG32
8YIc9hLwamZJCpFte7mcUpOb4asA52lOj5QHem1BfbJDLQWpvQqHvKd8+ehg
K6MyUvIWh+BpbdN/lGfisrWxaNMcIAuP/TO6tqxX881aBxMRA7Ee1ldVSJ/i
6GG9j56hrLUFArklWpYZF9EOUCePADw6qnRz/A4ATHNzVZ06G92yQtxfBRKw
siRvT/3oMgQB+QTyzHpDeKG09GnajO6UJ5kaD+C/yK/laN3CagjuYFBGhyG5
tJb3ev0dRl+ZvjBp1moAZpR9ecilgwgzbdf84I+6Kewq0kTp6Hf0dax0hqN8
V3BgoPSPUXrGaWiD6ShI9C5nWoOHoDpMirvmdU+u6prRbqQnzfi+o6l81NfL
fKzISOprjRpSwnCE3GQOFAZV4lwIRYSOdORbKAIyvMbWS2D8vHIMChrSTrhi
YdvJ+zU9L8ALrZS3wfoB3+TAE0cO1W3GqPjPiXgYHDWMs4lf9wPTGKrm4y34
xZgyFX7Ctvs5b4Xfs/PWVV5FvWmrVr7z0uRhOqvKdE0AJk6u5gLY1Irea9MK
1jd2te7kR0Bvl854o1cMHR33t3t64Qai+97SOPyOLz7R59imqq1GnqZHGa3F
TLHYUp2VCX8hmgdEELinTsWzhYf/lwHZLg6jjTM35PzAJukPvSpNHR1ui63X
fRiaRRO/+xEQgx7mgUOQTQhAHU13AlX7cyceWBqomKaPGmThVBFR+WJzL+dE
dCgJSzDDvvYYhDTOk8zr5hfP7c7KsD8WLevEEML5gp2RLQH8R03sAx1zWmzF
wloHN/b5xJc9wlLG7iJs3O6dxjNP4s+/xY9fSe0cTq6jdg8etlnBFqpWOP44
rYpQsCnwhl1TZ2ZjOpXIgLn8t/8n1UHW6rgqXfqc/tWkqtxaGfKIK5CVFed1
e4SjTGcS2BZXUE6poZtgoOIenDFZU96AJXo0uDl9zgd7JIg8eagVW6o8P9UF
vV4+u5IugBP1oclnt9In/C/CxlK80HlETj5IR3uElUVez3qq7HOKHkKpU38K
cELXBLP+CSytz/9hBOpYwuGdqSBK0RUhqvA9FB+F5/pJdIO0N6hXxB3Pzkqq
0qvYXgrP5v9RCj/XXVHKCMxsy/X/ZogBermWXBG7C1ORDk/fpyyCtIlsVz5J
yroExWoOd2rwnXsO33+tqYEm+7KXNlNeMOOzDoaJ9EYbLrgE8ORUh+MBCzfv
U3flA/FyaEd8GzE3K3Z+KT5mYkkOya4+E6kMsteJHF1eMgCmIL8vEZMxFZ0B
fSU8XYK3D2egdy9i8SVv8K/axkUXj/B4dq2akC/n2HvySD3qOzZiPQUMN14B
CY5RsBlScKDEkLI5TSun/DcRpVOLnioCLStQ2RmBE71TFsSZv0vgMJgwuLLX
8wpYg5M71viOOTI9QhobypCV/oWWnPHoFQN8MvSCjxAJiN1fD/jpf8T+8JtW
cf26gmhhHGdLIbJNBBh0TAAMixdExJRn9+1mOddnjWnxBXmJXn+tvUgbdUHg
5Z+DGkOK7BrOjHJytzKjMJ7ViYbfER9soh279sj6obLmIzQMpJ9/tiC172Fz
w2ToBbsC597Cn8YOYSyOvgSzK5HbvpM+VUZ6NzwZ0jS+Bc6qnzG0ST5zhy6/
BNzNwLIr5xOPeIlAlkRYRbiTmoBtiYbhr2Uwj2+t3JsCLD3l3vpGLj9MQGCd
wADVPFR2Z8ipfhQq07exMqXUpt5pLZtwrJVT4lA/f2kSf+48hsXuxMz8PfFo
yNVc+oztesKBpL4ozWOMwOVUdIe/OOgDLwrqHxKp6N49P/nB3/kzHq+NN3Du
d4yKkbXEDEKmaB1Zu3u+TmpiNxD4T6OkAXjAR6QisBncCnC8vwjuVvfSxQy7
fMX6lN6OwwRH/T32qjeRWn2/6/8rCs8i1Bo7nPPXPPZSg1u8RuiJa37a76WJ
7NoV0ifTTo10RWGWKxccIk7H4WgjFdgKLgXfFVhyeMiSuliSXpx3tt/RF1fq
zlZaay6FP6wSg6ugoYxBvo/A7zngh7NlEwghvYkd499IxV3WS+5On/Jzb2OI
vlE6+lfjMvyThGhcWCUKvFs+4M0Pcc4soP/kPZYjL1pjIycLSAq6CvIpVDwZ
IijcLgTotrgeVkj/3T84Oo0c1ifaKHg31+9wWsWKLXzZxn57sL8HW3gKYeyP
7Hd5MxbNZQZM8yv2QpYzguhBskgb5m/qfuOd762F5XBNxaqPtEOddrL1I87D
c2NK6W7n7l9D96egTsFxk0IK/sDO1StXyyFMm5bdgHza1WHADq1RTN60BIU0
mmmBgA25F9KoJgJIqKhHvEHv9o97ckLLD7hBCB2m8a1EvQvgxJOzmxa3YCcq
IbY6+Bu8ntkULoPHNGVfm8P1+ARf+QahEK2wEBzNEN6MCVBYAysEGHw9dUWs
GQTVDeOiuaAKdHzCHhq++b/EBPjw24ugWBLyWFKBytxMdU+pvVDa5yyDafsR
0Hzln80FSIqqlnvt0J8SALAE23rXlSkYafrVtZydLXNuJxIKgQG9mSMQGmlx
8QJ44L6zNRa4qcF+23CxU7b14FkXrZImoPQAnf9L2DlYcKpjJRZdhrMfyOFi
4q8ortUyX9YniBflGPhbaTgBJaRD9oRv+Qawam5UC6HbJE+Izm8mhpfXTb42
Nml5oCZMZoZpeKvGR50ghfC3UYT4iateuCpehE+umMhOacPSR6VpyGt22vBT
HvnUAqddMyOMrs41EJcoO8+5M+rWn6rQ1RAJRc7TLv/5lgMtUuJ4kwquGzbj
08+ZfNaUXkdfovljrKHfRBezYeqgmGyBVi8p1OtIze0E+YeXaK/NgdfBl1Ex
fSKxwAeZ9+ABKoL7WTahRgA8NKp/5Mb5kTgdKOmxWa0ziME0xmVa9POkVwMd
n6lo8UoJpRZlilbKui65vZ91JVDPdp11XAXBd1oZBro39X6erZttauR365Mb
0y/1Y04LL3rgvhjfslNXTYlnfluIrOtB1zww0xMvkbtVrthUDiKXzMIhPk3k
tgQapxzNtYbWIAtTqr2eE3NBmefr3U9YGTpvCmIM65ikIrYJBE9DB6FTkILV
LjrDawNWrABa4SWqr9WFNJw1F6gweL0oUCgn45CtvhsuGe4pn9v6T1Xg7D38
pG9BFirCGlH3byI0gn5lEK6SqVVySMERLOw1SWAh3kJBrQaJEplIV3cB7hoa
jPZciLhuI4cMjVHc0uP29rbAZHV/MIdDlN7hyrWPstFpgJbiGQmmgMEdkZTM
TK3ZeWORndHCR4zy7IEZPbHH59tN2EjpBuw604ucTXvJLhnEdicl57CnUiEQ
cssQbG1xLbIM7Uc8+YhN4LRPBbcS2FE1UiAkAvGJAdeSpwHX1Vmg9lTBuYR/
Lgust+9mfU8bcT8YCcbvk27aXuX1gFGTmLVTKWiSpdCL+EWDFa/zeSc9YNKd
1iRSQWxgHMrG2H44oyZmWxMpsy0ELYg173zP66nQdobwokfhNFxYDmfBiGGJ
G6WC3GXBKhrkWRunKgBepR0P0CfNksMFJafb5iW7CIw+D48LuuPYfMJYINzj
DvqEBjgtupnFmB+PwLy0TSAz45eme0nBbp6W71YBrX4nROpiQVWMcgTZNvhI
Q5ksgFSHRwy4K2ICL5YFATNUG+h0XalQLgQu8/Ce4CuLGhrjU81QrSY5NRbW
IbQixfQqg3DBPuzp6OkGYSVhj2ih+G2D97M2BSOHdo79hFucbYbnI0pulyWL
GmkZa83DgjEgA1ZpvULwW8DQ998U19+lbWLdzO2SYDPhcZVCE5XWbyBEq4/h
L0NWCIouABsK+HltfJJl+FfsSIoX44sy99VLJRq3G71BrOeRs1OWmbev6l1o
5eJ2OeIZtWX2jdELbYmsSvxaYJShn/AlQ8KySUonoFnnbEQpSxuufiNwonyT
/tO6dahmOKuzK8YKeDWJPGPUWppnhkE+ytFzOQl8J5kRFxEXrhltoBo7m9a/
QlJDPVPFXtSmOx2iFoieMJJp+w8vC447zXEehQeKBzv06lI0BoEw6OI2LzS3
W+rMJc5Cnz7W5bxiRY/HJn+vbS+j9IsAH9eN8Hw8tIb09PMfjky+YBfGMw9N
eVoqkxX5lh8/q7c0zmFppRDp7FjNpb145K8dYGLV9T9vAq0J3z+TPxKaE5Bp
LLUqCRkxaKhj01IGK9HiNE0Slg6NlHUD4a42/Ncr2V4MgKGoaaAbzfuhh1K+
KB9C5Cx4+HFYaLNVL4l96YusGeNpRDfpaWcMjTbacXmCawud6ccQfpx753ot
QokBV2w5t8e1KrNzNkE/IMcvuTlxR+ryn2sZtPvHefOz8QxSar+cpOFgb0OW
6A0LdmLGsJzFFkAnv+Kki2JHz4f5e2pY77uR18cgf1gl18HqITsdtE8x11rh
YmuTrRuYpXA4GizXmCmW0NiL7imoAENXI16ZOPdg8pEPCGra3RRJNPB43kU4
dZ0aUJQGNCbCitV6Eg5NNlh1WObYw4S394xxx9UlTfh2f/+27BqaKhMpU3p/
4YFFxfGUC3X2lOilb/JgN+637e1Y7mZDNTExiXV/Qj5BL+zm68nbO2l3Txui
ZZWr4HfGqVgsdp0fNLbbtOVxxYO1xH8H+pxhB18yS3SJbKk/AIUZ0cosY0VH
DcthPNU0VDpV3/5DQfTA0ZLCqL2MiKAfF+NwyiGG6g1PMpGtvFlz4PgSCgxb
hLrNSmLm+3NohVGDwQLk1gzZiRdSOXlTSxsV8UEwPTENPvMo3XHhwfUaKrgx
ZhiZOoSYrVEsKMnbzQ9f+UGli7MBjyf+IUA2FJjpQGB8hmiiHiK9FB/pUZGu
dRqRzh4guUXl1/DgHQsAz5wq1wf9WJYKgyTj0bnB0RFkdr/Or4Fp69cmNt8U
+pjclrZs+b5EBovy8akQ2QWsBJctb0FJjhqk8JQ/Q8Nm6kBUpPcc+1/iVcw1
sRs0Zih7b+Uiz4HVxeNh5Hy24mhPDQjNO3i6tczep96EzzLh3+SSi8BS//dH
f6mXEk3knPeebfS171HsKcVxaEo/JkKDTgXC2yqhdlhdZT/dsmCLyGKNJs7o
LvwIoHgnO4L7EDr9Li2Ipz667md2qxGXtfqVT3U+6moNWd0QAxymt7Hg7UUO
qgvNfQf+/psbcLXWfPa649evhc2xCpAwkZeGj26Cr7pffY898aeJ78yBaKaH
xniTYNuqRqeDY4FAS2sQonpIdr+BpPDx0ysTl5EEa/EmGWkAaSGMbybNrE20
WvueKo+MO/5ktdEI/vUzCDqGNs8kIC8PADGo5K6qCPuuZ5lKcoi5mv9rjQZr
BiYgupxBFRbO59oIfkS2pDiTKNOak99RmK+e7qmUdHkEXp5s5IGujB143z+d
fabNr+nfvuFgrn7fDs/x3DLhgjJBfh8+xV70iluxYJbGg4FLMq3Pe9jVat8o
a6IpGkiFoJ9v4/O7DziMv4BehZi/buwQ2vxMoFuf4DOY0/CoZTTqUeuJrbY+
81jgoFqDKuFAyh/97pPGuGyzrdC8H9Dv8EEUVROt7oBPvPJN9D1Bp3JbEpbX
rq/XtCa3o3yZKo1SxLj43TVQGBFgq7eI+z477Gss0KVaY2gFrXczGSCXUuCe
/ICECBV3AdLA71MWZxeYOHj3FbTRZKk8EVkQO30I8DuwcFwwL7j8yd0G4kbQ
NMokRLtJRdIU8ZztmqKglTZalb1e/txwfqEjEB0FXRxJtiJ8tmCOmV9pQV2G
vyzicdbB95tsQGHq8Pm8SvRRr7Xup6oyjYz0uyiNUBFBiTnF6pGfzDbM+kmv
L9wJFFDRI7e1IUWbd/kSR3TYg+usL57IS3LCE6lbz9aveMzVcjACzxwvgAGT
wxPmDpTPwx0v8KOiMqOJ2P/k2LBFJZflAEi7WOpO96nG7+5qQFWsqsE+n0Hm
Nv8/+o+r6yHYvZObo7e+XrvioxvoFm2ZxuBPGlYuuY585izJpwNnQHW5IdkP
eiXkVouBTsOAeeqIbTNAe2hoFWNb4xO6esxN0yFAyE2gV2j+SXZeoLczOu4B
lyfNtGK0bxb8Bhf6cM0lgqWsgu0LZkwQT3kC9bqIhRagzJzMqD0iyceYcAuf
OyKSMJhGjlQGpb9xw1+U/fyi9ZJyRwlw4YhDcGseGU+rP1bI8LJ0caxUvFai
iAiZ2Pe0z6CYw0UoXGJLaTcbLBfZ2HNta/x7xI05U1JWHL9ILmM9ZQlErMgX
LfaJUyYtENcwLBZhb7LdH7FsrtVRjzk52z74M8JxtSxCmIfP1jMY6UtHcJ8u
PhulYNvaK/7qomHmjtaR2rbsaUg/smZ1q7W9IlQ7bKZYSGeUQodfzpxkcWM/
+sUUYAcoHUdxSBiCHbufeKHeyte2zeHu5YdIUjLZl6UIPG/iUJXBVoW8PPex
srq5B583Ia+DrUpOeMgPLdLD6R3S3c35TJRrjwMaEwh6oi/Eh71X6PKe+VaG
U/mgV7AvcQVdKbma/hqjcOyKin2RwWRT8YGJtPvb8oMepEvifj56BwZ8qmul
jERfp5TbN/KI/sKkfH9j0DfDSf6dri8tmK5R2hWmG9Y02iZhdSSuRg46l6f4
G6boegdNYq+gfikk43gVNUKH6Gno0c1t/VlsGbtPs1EX+YixMjtyaZmeHncR
fyuDH0ShzeVlK8n5sy7+dko2Wy/ZrtMRCg5dr876OwZKOSVJ4gvGsuJrqTFK
2epGaU7dJ0mtISoDGsWiam/W8qPZUnmkzpUV/G5txaYeYpyIvVgxJkoGDnUd
LeWhZwQogSnt8kIVOsay2vIwUJ9F0Y8w/05fN7h224hdDuhJsDP8zuxZHB85
ymsEXYRnZ0rHp8rXBHpKsrtRStAMHVSW/v9UWsUUa3/l+pGsJMwjm9TW/Xva
nRN/BXHsM0Q00xfkvNDwHsW5U0O58qPNFi7cxFBSl6H8BdWC76ThzCgDC9tl
RZkkXjoUoPtB+gxA2vdL7uoKEpvuQcLklbvzvwTGpDJ+8wwvHIDJCN/4OvRf
biSBPV+SCWsGPyqQRmrk2g51wmdauCtSzH+NBVCAlKBK663fCPCXbV01J3O/
rKSDto8Lc2I+C66HEBLreN1AE2RDB5C4PJOPBjJZNMwY1utCOkba3BP5PSOY
wTzYNrOpZa0Zqjvru1/WhxR3dxt5d+40ejeZYU1brNua7en54a3fsoJ3gPkP
2f64CjqV2w0zEsTDBuXZaKOzSXPz8JH758t29mS/xw6VvXSjKmXyS2zwFHMe
59oUIOVwHh0sTCcyqcceiLRsz6hIKXGkPYf573HXML6PrXAzl1VhGXZLFP/b
8yBilAUwmRHhlIWTNQX6NBtpo1ctBxoXklr7vgrJiyg8tKqDfWLu93GLKhOG
7B5zoYtFzTMzL69JPiqI31+HwjVX4u2FTYiLv99/uY1aHFCGJwWMWDqnXV+P
9+nbcTTLESMSYgIxnlacPtZ4o/MdbhcfvR1/rFCwOe4cn7vQ4cXJhplBw7pa
0KNaBA1hC6rBnB/VydKdhFkndiup5lkWo0Q3jmhaTTQId+uUhpLmaqwvNELs
TrEv4VnJ3R3JOX1WaHBV1Utd18ne2QRrCuwRLDWN7TX4daYCoggbymo1gdfK
RJV0IHU7LBM1ddXV2gvuQr1T5LoGrqbfogDcqUEkpGvpvoJ31v0Y7W/nmZOQ
VZpVyZBKKe/7sQA2nkbBhjxzbzGL6xkH6lMim8hjkiy/dbx3Wvhoktoy+uc6
ou+pYiQEH/a0ZdYhJjD9fX0FlLh4/VrBJQe73raNpuAJIVGo81n8E91L5B+5
GHXHVwY7AjzWyFBF6ERL8bbIwrItqrTqMt2x9WUrjhLvSkW66gq0LOOGPkhL
60pX7exw8JNEJE7gHpjVi6E0j45sFqfXvHuh6wMSxp+rn5Z5LF6zs8TqiMLc
ahWbnaoHmC6j3Z0CCKFoDx1KA1GIMS3FUyzrxOgTgyqZhndPjuiOmVKSzk27
4lp2EqwZ+gy+wVX7catMPxSNPeW/dRFwyiXiTDrxQEPjaheAdv8y817luMI9
g++9NVJYpoutW0zh0MAjV92rUMyC36UpM+ZxMZjkqUDbkwKy+5WVAyjeLrYx
5uANsq2lqKr5VVPy3EQAoloGpmGxkYvTo9zYxAf/eWt7696K7Mi7AG3elVMU
AYZw/tUVG4thv3p6GcBkg0oUHX7rwMvqdVeyhRG6Wr5kD5fHYAx1n+5uA2pY
p7CXl6p027N217mdLLkRZyZHo+xV6OS7a6zXyOM1NPKk6k5zCWGYPYnSUZMY
K3UcxM+0kurx03eF+M2f+Y9AR3Y0onWuicAiQZcMCwKW/cF0OJwokA7d6bgc
LSnj1cnsh5vpLDa3bAd5jiNdLbwExe5iYoYcQjDgzsElJ4cJrZoe7ySn7hFZ
P0rpQcm5LWd36kJlQNz4to7IxF+ot81Ql6rH4AO9faSJ2G+s8Swh2jURgiOr
ASaj+GuDt2TJEoS3Qk90SgeSr8U1VcT59KDPLWhIRLF1R/lzsW5CgPuh8kUv
eyxPHiB97OZXNomc9xx9oouhrg1BMP/Rv3JD/Vbc9kYWjF4qqwoN6CzK5HPI
43JiBJ7mdrelxA1tVPD2Ox4oJixytEUVVMp0fEQKuYUGyqX9qemCCe54fUCh
Zrz12hDFuSGNP3ShFSJxPctyyqilfJ1zYfgIHZ6mEwKDci1Gq4CGXaCVzFGd
+eV5JlHTleLOniFdGz71mAKQfPx+0H9V2rPtvpPCRUMd5xFrN9PdffnkaN7c
X0UWumWa3IcX7QO4lQIMSo8cmDr2qeQA8igBZ7HJ7vzM1sVy5ZV4xSp3GlJE
0DXwpsa6a/YBK5A+jCojtF5CVV8wH2Yf0qTYbvcriiiwVRx0XxEIZBwfd/ys
AiC6ExgNZXeqzOmlAY4TOLs+rx0FOn8tA7UoNTziCKfS23ONTr7Ks2T60WAa
Gm5fmcWGbq5BoTkfp7QgrVMVLJZmBIyYxxbuNCnzrKXTjMOHbYAyUx2p0wAi
UCmgeqUg11vQ3xDGWF5lC7XAMqcvNF9awh3eV2hUd+2JtnXU4w9ekVCG1JQH
842rby2x4GJR5vhXVwW9EW9i3UxNdlZTFIdC/ujD7iAYJu+Slv4a84/YP448
9FZR1Doooxe+gXQkZy0sO5UcGa2UTVqD4ZNLfuQ4ANGIhqeuKX6uiv1bThIV
eKo+PEytrogjsO2sgQP7f4VzX9V1WJOBTq2nR9GfuxmXVNTsQojggJvOmVQV
LsvzdaV3dDT9alOJEZyCBePDxEa/ZqhBrwhLycst09Mv+hLCN7hcxLVFLsR0
MnkoqKQEZwICyAuHS9z1tRdlVCiM/oI3uwF5O9rlrDh6foSOoPQ/vlyyL+qj
uqxaJYQzObp8LTKLz8jeIQPgwlTRg9s8/Dp/1uX1olmjlKRcsgXHxeS5mNQk
PxYxL7HTlnS6Tkj/cfCeYmzu/bNR2t5a0layoyhjLTIYpL+KXoAT5CkxFjr9
0QsScsrdomYV8/5YkDv0qDodP2Hak/a2ihkYjvNNQTYNxtAxDXGRcxJ/pYTr
RbSdwDyaGXhMGAgPGjAQOum7oPTUoowfBApbPlT5Soq42H/qEzy8V5qy0YJC
scGd+GIpaaEXr5je/NJodkyfxWM2eJ/iWVOi4DluYwa7dbH0rOBjI/JAegE0
YF3YUKwGeG2VGnsXeM2WYQYy89aKB47NvTKCpHp7xloWH8RD7ASihMNELrWR
OmQCDQIFavl9YDJe2haV/rdhrtYb+CMfVTWV5g5BIsQCMjIZZMzMkokN5zuI
zGI9A0rZV88tvWEuXCwNp1C28CqEdul677Ay2QTVajNEKH4Nnu3kdL5V/Ba8
DVj8P3/S10GzAO2xhjg51ve5390Uc38FBLjsNhxFYfH4L20ka5Hbf6mi2VN7
5edAk8Vaj12yqSCQw6PI8yWIxRKiIcRi2PpLFmWZ+x3TQ8qaxVBINWcZolvV
xzC9PedWbKYScUL4DuZxIdzusbXO0qsb1k34Mb/UvfO+UrX+imaE9alY+bph
YsEg5Ni154oPvUOd1flYQ/re54XuvIJtMiyEDwXV42pvilsg0dZc3V+rUJJB
uuubiZ8L/S4+TRB8IZUUnEyluKZ78/2/EOnYneOK6+2qTl1IxE9lmbhouCyp
xeYqiXvjWtyMxU1rng8gEUmiXo8HXgHf5zdGmnMbPOUC9sQn7vlc/5QSq+0L
oyWQGVryR/mZ9WGsc5TJdhKde1cxKiXyIntzW8YLfvhOe15jW7zIW3v3zr3E
ZBFVrz+yg34Je2TywN6PioYFS5w56Ey8AWaqQEnAAmTJgbEcBQwzeQAMwRJx
V+uynkQePfCZzZ+S7AtRTgHDJ4Dbh6YaH2OMJWY2joC/vdfigiK3X95iHiFF
t9AlYM2zdh6559mccdAAhJoY2VJxn1BMScaddvAghygnSadog8CBX83k0Qnb
IFgDELz28Ys23ierxz9P0qyrFnNmhQJ4bi1i3wGfyoPYSmEBXMKHwotq0K3k
pEWULyUJtbwgB0XwOOhACGvoIbjz8u0TVmyMQarfz+GareQaUrwXq7zUPpM2
BsPO9V1ELDlypdrzNmcuJBV5lBPbJjjPzBZyE6obdzXnFhsmr3HCMp4jQjpZ
si9TMaVMQ+1RDRcFPMkotbCSRn3saI3MLq/1WFT30Qe4vw+aQbtNyPN9Exi/
kbj4vJF1vQnF8tKxMHvEIDLx5qRfLE2HzVrcEsu5rEikiZ/0WkYjEO/eeoIY
ROsG1Uz6pq88QxjFSuGK6z1QdgXVn3odwqQyUr5/+TgDDR23X4gARgJKYmch
0VfuDF5zc1yBcGDc9bCtEHPboM9ZviZFDded/FBf+5p0JgyP2DQQz5gkeXIk
18/LJT3Qb2bIRvHNBP10sM2FSeBfRYqaYMgGmHQJnLceki8WpT0o21l+IYH7
DEMHHgbAY4ODE9YtPIrpA41XBHB2RMj3SwoqaOASsl9fx1/DdfTOX1ecGuhB
/AEvuW0OYYgdu5eNWTaq15RwUtYsCqb7uAc4bjnuKHibim5tUZYE3916rplh
HBX+olxFjlFXxGTbNfYK251ziglC2Coq4a+vdM5DBnIepedt8k3W7Mcbjg/B
AxYL7jgjgGZ/JEcxWNKLNueTAkC7rjM+C3ibYOeQq5wGSiii8IHWN+7wpgFx
6qwAxQvM/mexaKWO2fACl9Y1FIIiuZFf3R1juKbc6ILlYpUTsCqyfYO/I2mx
IyN4O8wrUmUdhKGuGSM8ilmocRdpcXihq5scYaFs9JO207XvjihEU6p4gddh
6tS4EOxx128ZYf7Zlf+5q0eOnK9mfkei8Mn0N2ENtZFz0AoRSkO1MpuKmyme
nVvNs0ndqZ4zUPViaIrDyz7LKlWDqJS6o8abfa6lS2/P91YjVtBxFLpT8ZXo
PA2t0vLNt9acbHNVHwO+ckjX5Ej/A8OCpUdXkcRNzCBrXKbjgNnCuB4vEhu3
Y7x5jJHZfKIGwyjatSWum/MVRLJQfx5HB9/SyCUlp3SOG6czLme7fFeVxQ+Y
Mw8a8GxZwWbmTNg7FEsjs3QvguV5hwBUvPEbZkA6zRgDGYy3H+Ap2eTq63Aj
2GrwLLISI4rTC6lHRmzmRE8/txOoY6mYP6FTl9vsIqKZW6p4ebGz+ELnYXf/
JdpuEhCwErzUIdVmu1zd1tq1iPxgP78lqy92a39IYDG7DqW1bJICV4PvU9g8
DRxKvxoiu57EBA0ZfIWXTohK8nsjpl/xSu2P4PQE1QtbJW/EV87YKnMn9oNu
W5g1yCAB2jjbGdNM+9weXdkLGhK5hd9gqt8lYNSO94d85AWTuWghjyPcNzHi
rj7liSbp5KFi9ygoLsJz+KogRqfYHQBpr5BpNlDDnOabeCnHIccJ7fVt/gv5
S8mq8k0Fdo8PBOtXR362U6dgciZVo3vUa/tTyt9yTbwUXrC8xpZt/BoVyFZz
ll1QZoZIrd59FebJT6yz3BTi03w4DjlWMSYudCHXhH6qgzq5Y++Lrp8FELo7
942zO1Cp8pTTg1tm6jWPbkNmXwVY51Pmckeu1u6/fQdclCVJSSWqQ07gslNA
I/eR+SLJdJe/cxrJEEyKqZyarYUHfxjFgW79ufJxYkI+EpwlUlxOF3XSUoso
ZnxiZk2ujPSW/Nudjwo2ZNnKqFg3dDqZIMr382OwEREHAJneAj1Oeemyq1AS
QBphp2jsk6SrQQFvH9zEDGmRndB/MFsAq8uCNUieQDCDajbfIS6OzDV5Filb
LiIng2beUB9kFIDsE6VtuZpQMmsUS0kw9KFsrFAgiFqe+yHpd6ddc3gq28Cg
KRxOUEOQZOtxHMASGXKoRdn3CWXnsBVyX/q/MLRFvQUZD4/Ma3KNq3L+xrz2
z1ZaWV2zNRLMg3SVx5W7rsy0Th6PSQl0j+lBbssA8/PJYdvGNrsi+fJKC+Za
mHnDHfGk+QwLm2jZg4fzjbXzhkpruSkStzSCxZ1UDhMmFxxESVyXR/7uEJA6
XAWEzt5anqsMrDgrtCduzxVPn40w3c4M7m5ewt0YxunK1FjaD7x/HT2aFoYs
K0GPMKDwWWPZqHXUGtL9kcZ3x01krqruKk5rVMqDQqC16xu2/SBUVwx2pXN7
9XC2cGSZ+SJTRpA48licAuUCUA4CrzjgXslBNn9q6OuOkS3Z6J1TzW3+erPx
9ISbaporMbbbm1ws6G+W7PUc77uuDy4lNlIJAFm4kpACc1FOjPfrkI1dNFRc
aWejZz32bS/chLj2Kp86Dhb0tvc61475+4AMZjZTkG/pJ8T6TgzjyZzKQkdS
e/6L+iJaDfwss4oJVxv+uWW4U9lCG1gwLrPha4fJ01UgHDJMbyzTivQoQWNc
KmDq4H+UsTM4XAPXQBf5gm7oRuoARQv2nGbs60/0J7Hm8ekKTeDnEeHJd0KS
XOXvMP63CS9UztU9MZb94AHSSao2RAUWcDmTv4brziZlRdGKyUpZX3J77gVT
oxs0Kow23MycOynfhz7qiJaZnwj1FcWS1Z34nVsZpeKvfvj6CXf09yiE8FFg
29aDZVNScfc0eJCm6HcTkQWiUPiOuqUgqwbehMTJDI/YHunV9oYNuI/1EyrW
UeUc/j412omllJSUropeiNhvpFLf6xnpDt+6LDkSOtO7NoNbWbGi1v8VueIt
HAajexyRhvUnAa12lESWM3Fm1nCzZjT03pA8azuWqH2irIaH6J9ooGscSN8S
WwVOfNi2D8LVy0cT3Qu2bOd6sPaC8DQ2LDIaxgAa9OdqoJHBteaYTp5uD3u2
4QfY3+XQVCOUOugJuv669CdpwuOX4v+ebwHg7ma3oiSLuG+Xp0kxy7qZxPwP
4r36hfYzEGyzGIwoR7HxQ49Rw0WJx1NayXHXUPW3pqTMTN0oE1+OAktxzTqr
5mnaq4mMO4gLgt6DImMOuMH00aaIb/lumnf0w1wdL6qoktTmkcQA/M1t2WDj
/CN87H5l+uxG3MapAmGYXxxSfop1S0eEs3MmiDg3B/AMsDG8B6lMpmAxijxK
//tcpUMDl+WaLjDJiGxPUw7zxIELxDBS0EyowhbqTvFyAAZWtYCoxJbxko0V
KIi9Wu/cnC3Im7ccjDJFRMCrGF6X47mtIL/gV3/5vYkzuUmjCLDTyFIkJ5AJ
geFk4AYxswtezcteR9xQizGd07gl/jlmwkQjKvFtLF4OaBC4QHY3ccJyAy7P
jtwdcId8KH6Nl9K0spZ/kEdIi7/vzeJxan8zvNQzOawcjAMkKlsGLFaZpBaD
D3mSj0d2nJa3j8IzzXOwmGByOWYOLoQ+AldPgSMy0ev+HFoZXfItIixhzddi
XdAzD51tfnJAZV9OSftHyFYfW873otyqJJ2bAEB2PU1X3ey2tjzBAOxL7YWd
Nb+SVUuWskxM6YA9pR5BiMQ8gCEZBIad2icxQcegNXRhF2NocLhX44fFTg6r
1uBU7UFkRXs4qT28hV32lWDxpjZFnmaLlkGynSpoZpZRg423CKzVI6GUcI7K
qiEA7POP7DS2QLW68Sc6/rzF2EPH8iq+iLhuHtQ/KpHcXG5hN/FSs8lPgCbB
0zn7G+ordybc/GEjk5pZcsYIP9P5+xLZYe6IVE7cZBYUG9OkJVOrqOrLHTAy
yDBduYvc5fxRKhW82dOLjBVv3WXOfuj+H+w+0wQgH3ctGsqmHa5flCp9PKvu
zMjGNE98C/gaBRlwtmNM+9YOrW9DhHiKWFBfHoFg4tXOKjCJaU8G6TAKAwUD
mV9sNmaKrGGbm+8/DjCehtBKCiC/uT3BfWyEGdoV9PLA3kWV/EqN96N8P72f
nY+n5ylmvM+/kZ9pxVpCGCktYQUlPRgozfSl1mHKfY3DwdCh6sinEs1jbqSf
cDCTJOdNRzSm1haDEKPwlmoqCkOOSp5EeXWaJaSBT4Ui0NyhWpZus+WFI/Zy
b0Us1rq8GF/KNN71i6JBkc4pyHNurDb22AEczhFF3i7TnhkyaPKTeiC0e34/
mRKckWd8L8a84AexO18lCsK2wiNpDFK//gfcwaAO5EBHpGOsOEwoWOlNhMCb
YkVGZPNeXqBd5rC37mf7Z+36BPsujx3bUSweEBsuhwEOZKh9sivEi5pGB04C
+T2F+7CxyrcViG31C5FiafdGvNte4GpAT4CJmNqSgg6SpYSRVlZ48xu2pL7U
RoYHGwW+138z56bAnXLnPnrqa21SdzvND+OpHeL/HJldyfLE2Pnv7tPPc/TK
nI4WVOSiIym5FZHIxyG297O48zHU8T0pduYAThFfcuQNhJAZdZOD4NjGAy+h
6xmYFK2dgPBHFNvXVG6sNzHnrRxDDKDhn+g1qnbZVhLRsezo3uJ9XivmYBR9
kfGR0ZCfieB/jtgofW681V8vqTvZ0DMuCWFTg2lH3EDqje0byuiUgZhU6wbg
YF0wwgVCICsb8v00crw5JdsSlBabQYpO82Td7iD1+/pvNo3u1DAy6nVRYmck
dp9r/+HPKOe4NDcNIZiAYv/S2rNvw7onOz5mZO/D6sIICvdpdiOM/gkBeQBt
Dp50EX3LZ9faQKZBCzNSgzFRsvuakWXRK3lTzBaxvtWmC+lauyUnuzL3ToOQ
9uAsG9Dr0XP+Jftt9zD4LdPjwQN+FsMJr1NmHDU72fvkU//Ypniue2YXCnAm
uFJKH89QDRGiF3c9hOndtAUTa+N4pQTdt6ftry9zDIHhtHlaKgFLayVXvlUa
O5XBe3Al4c/reGBsJ7qOBlc1Eyb609gVzC9nhoI5NBPcNvEFEHXhDFN8hoPD
sBO38r4VJB+Pt+9GxzD97I38I2R6B41qgkflkQcYKaHkIfcZ3fDxPKTuWQ3E
6dPrNFBgZgIQd2PAfXbh6Uy7lOtYgu1UxUNLcoGNDtDDAKnvV7HcN4cmooYD
7a/Q1iq2ErukCdJwOFO9JU7nlHsGbJmZlZwMUJS2xYmdebnHFyvKL0im/jfR
Fz7oXDhcswlXnGwjPZ5n/3ulcGrp7kEi0RExmtqYLyFbniZrTkH50nt2J1mZ
Goa9xjdHfxX7IbZA+6OcrvBjYo6aJJABe8KB2hFyZ4k8ttJR2MFwopD3LgAr
j4Ns5eZ1GhMN+XtNFbhZWWTY2JnF0fIuieBbs33SaPdvyHr7doJBBdJs9Mne
iUEPR994zMFZsqXSGclTU8nR0HjdSwlTClIW3kW1CVPthAkBcNh5gMFK3gG4
MgGmx+DoOBBjuZfcvttT0gNAKk/unUe5ZlxEUbKqa8e6rIeXxpNKk5k7o8gF
c4MK0ksOA2CPz9M36oQNF9ESzsSTaL38tMotTq3ZNRDoMHRX2BD4OgOn3r01
EdoZ8B5Gzv7FvlRzEJ9G+/c15cXQ2id1Z4z5s04ist+6zWj6uuYGfrsH1PxA
1ayA41eTx+OsNzVmodY44ouqt9GTF4v9nIFCljBcVDExPjfryozkUfGStziC
dlQH0wJ9ssuj5qUXAIJWMGOzWAL026tzuZFNwBijNZ2qDYNEOL8TO1h6PqZ7
GIjxtCzSR/RwPwLL434+bEfZj5peT8PSRw0/Gn4Sx5PVuaKGzjcxu1uPqcWT
1/EzE1WVElAa9TNzlhBkwmYKvYVJ8w2I0ViG0wKp+uZT/lGTouDXYr9pmitX
MS126x/IUFEPW1p2QuXDkKLChj5JtVjI1MGgq98PSMLDdiaTbN7Miy+6yjVd
mpRp0hCIvt7Z5u6GDtyBqO6Yy4Kcc0ZaDe9sRCuBYyjjp19XWP/AFqNaqSF/
K4/pgB7Fht4r8pVPG/C+O6t1kLZODrsO5XuxbCmMa5ShnwJvhgTzuW2hFE4e
AIGfCRoqiXh+QT3c9DSAyHMXg0JZ4vPezEKRVuLHiiJ9JbIEnjc0/7TBlpj3
e1F8XCzYQUlmHxhBo88ybvkfC4f3WnL/8rRdUArrxOHEBrcG92qI333cxwVa
C8RvO/HIA7VupCI/4rXdchTJraQpWgIGpRiN9ryD9vAT1GRtKA8pW++uPEt4
XTw78V6cEgr8UDNU8k8SB1vVVLxvDrfan6YFCIJL02rouNinyRekbVQgp9WF
1c/mDh4MmL8WpCMuHalN576a/8kQW0UYPel0pESVk1n39bz1z13tV+2tT5Bl
TPzLEATjkmzC+FCwa3WnbMzk92p8Zg/LBz91pfQizjVq9+ZcH9o6bd81oUNb
Kx7Ni/VCLP77BMZ6K4XIaBsYwWantwxe4WfHW63cv6R/x4+NoQeKAsLcS5bP
PavmBO/qsnD6gZt+GAuOkiYMpLmSf4KRg9DtQR03ikJrcu2XjZXNZDV1dZHL
0gYQFL7WD0zzYrXNhv42cOWxYur9cze1g+G97QMmF8qUIvc0UC9r7LgobFOM
zmda1RevkGawSR0Xqfg3EtPsH7uZVxrRVDVTYBkvT4tlsZBvUyk1wjRuCP1F
q5UQP0t/LfYRx8I5qn37RXxqJp2NX0dUlrwTvJr8javlWNM5JD60LS+ssWfQ
WPmYY3lbn4CMCYo4y2Ag593+ovKT5B46P57XrdW0wcTPD0q/XC8L64ix3ncz
HozTbQjdkgap5j511ejVF3jwFcyg2KLN3K8wb+/1AlbeX7Gtx+cmAj18/2zB
l6DyxVceXXX51nIMe6hFgOrh98Ievnpb51fpAaWA9a8b60oEh2UbgXoBQMHi
+DLG3TUyzFXo8zVgfTga4K4XAfWm6SuRPBvtW7N7T3kaPWEokVz6BCXXBmdB
lKcY11qnnKmbU+ydKE0SfTZPzVcAKeacjAS9MoQHSvSkQXrwTVHbFPMEajLJ
3VtNWI+ccfp8KubsyQDSHY/Ynpm2hNi7KwpRRxXl39IuMiWJO4UVYKUExXxW
hwn3kuT/jvobHRwpGxTrx4+G/ZFFQZMrowFyfq6wMS2Ec0TdFnI6nZxD98P5
CjZxBi2LMEG+fZPwtEOSX3C+/DFrU9TfUhVyZeSusTeXNoxZu6irNFFCaFGD
gf1TdYqmJqunzIm9Xzmagf6V8s3sWehOB15rblzd2o/7+7HztTKxFyxtmmV1
OZe1a1QPvAbrqlX9Q8XSVeGUqfQ2+KpN2SaJFwXNcBGpswR61QYwpITmK9Sk
ASpWhGzBHGH3ZVn8GX3rJsUNz7W05Y9/TSTmuqxeRqWL8p11ArcB5FvrH7eM
PdOe5X4khydfTUGrZ6l/HFGGNBrgyzBDfu6iaH0p8zF/6GiBCUPQCcn1/OzL
3Nt5GiB0ndgLPYkVxXtWjxmitq6WMUTdP7CQwXWvGWqM1NZHGI6xyn9lecO5
vdlXvkueZih0Aee+QuT24h+GPbv78ZlVqXljQb9y5GS5femATmskKNaV8Ll+
sfSZ2jWhXaUNQs8ZM094lEzKqM1ok6eaAMpfnjOVU7OlO1dCIfnvxhaIQ+rC
vh+dItEhZhIwC/IY4O8FxlpuyGiwlevcvZRquRrjs4TBcRGlhz4N8O+GKHwr
3nhGetQMmaIl+lEbTWoKQx1O9tUt6mvs/mW/vrrMvLXFETd3WYbi/vGahGMx
T717iwez4mjTPnz1gYcem9MEftL/oFxfnrl6ixO9OXt+wX7Bqsl7oHhWc2hA
7qloKSJ9YHu5sEO2COP4hZ5ybU8wXXgJDCuHKeatMj/UB2ZoHH3Af7TAHSkj
N1VnBOOe1ODSCo6xZHvx0yVjyqmMRbwX6EBFGZ5Fx2z/LZ5ZpPX0sQ+8Swyf
Ml5sxw3oR1GIeJ4MMFQLFv/KpNUN5AOR74VbxlBUWC5KQruOnNP+9bBX5a43
FZp3fcEbw/iZnMM0da+IB1WygbYdXkiYvKONdRVDxl2GnAL3kmp9cQzHC82F
AlkebjTqrCl61EBIFrXKZ2w0LtwDmRpAB+KQxs7ba96wdtY/7mbgU8ZTb7Fk
VYwBK1ICagyXCL/uvutAR27PQ8imqxXBRaf+mXNplZMS4Ez4U+NR57qgSYCv
zHJKTYpfYIaKHgDeBVeuoxWm3bNZP2dGvLKlqc4FO/VQ7hqLXhlWjR6wUMEy
48Aw4HGrOle2D9vNboJtP1UbpEBhWUzsx6s9XViaoxJOq5yVurxX4aBlbLZY
N711bni9l4jMtyI0zvrD7AWdgqYLnJMys1SUl9s0lm0HimfWbgKrWprHBh+y
oDKPZOlszzQXlr4BFslyodOYCBzCPcAaQou7BJ5ADHpSrthcQO9aQlx9s7Z4
Bts4R/eI0XMidhdcBDMs4nWTtoQDhO97rBng1MDZJnGAkbwZo1vDL0Rh3rgA
sCnNueXf3Q0w9rqlZprrItodb+36Hbst0X42qLi/oKuqDQi16OcjygRkm8s3
0iyxm1oaTAtqnoc7vPB+Tqt3kUQqQ/pCdf2ioyGZiXpS1frrOMY/D7kzcLVc
j0CntqpOAIJqlHha5YI2axGY5Nd7Pt89edw4+Ch9VakXAP795FTY7/a1hwf7
qxlxV+HUna6LqLwwlO0nkd1FNlHnXjiIkXfdt8vg9yHSdMQY/BhY6jf2ONMt
qCvgInfWQ8y7fMn/jk0oSpta29dtgZSZxuGsCPtLHMZ2SRokFIbMau23CBXy
epu2Wqf5DomPbJkrN7ETgcS9CGvkpKkiguzczGS0jx/1Vp2zonEnC4hqXdmd
P4aMHZbI66PiABn/DBvJ/0yGtzQmEJL77PmT4pDnpX6YOrLCDqLEguQmHnGK
xlDTWknUKi/kfwkj8zP03KUmED/42rLn8pRkBHJm4mFVKRrePbJql4MdPH/n
ARCA4ZmXACroqhtFKC6i4LY15JFU5k5cs2YtpPTwUavVtI4CVT1SPszszztw
SOmo/RnK0mC3fLlzko5JyKy2sC8sWNrlQynhD1E3tg58ex2qISZdSax7kG7I
RCUUrFI+8X4vzXdIVVCaZGghNaXGMAAv0ovC+67IIx49DYg1+sF0bpoXeWUS
ii6tJ7o1ktBuAsZ1EfzhGq7sSF7gkgcsSlspf8ey4nD/OvmL0M/JliUtcP+6
rlblXIzUD9Wdv2Wh8Xl/hiGixkygipYNAvja1KSI9PUXovffkAxoRkBSo/pc
XZGj9AqfOaAiPruX3wHBtuFUIN9nMtEVN9HRp5DK/IWm7HD9Lyavcb59SNlw
u+nfDIlDNM7SI78SQOi2xEk1kEwqCoFgF+lfoxccGzSTkPk5TNhg/MBTW21U
FCPJDanHnDYquRs1bpwoaEjeEavF52IqBjJkyQoyhrBB/FJa/6LvFSxC5nxk
s7bTNUbKT0LA7h34rYkrsHsEiNeVqQwd4U55rkJmArbpH02VaUo82VX07Rjw
GccAIDqL2wbXTcu4zOW7SLjeIdwpRQqqvBqQ9nhpjdMV6zIWXVqwcDwmRGkF
CNxbRFM+5EqEhworjqPX6iX76YFa8umeCwl+4syryltX+HJgDdLINDD1LxzP
AVOSLXbupRg3Yu6XegxWsdADQilrJ/a/NiKj7KgZj/SUZ8GKDc7fXfCjIotU
NlSpe5rlkgb+yqdy4FiHlUEgbeH2pzm/8s/KLOfE3PWKUilYnkzCnNCqo8FB
LfirbdXszFLqB8y/IfDxR7cu0z3Zm6yMDRHn/cRJGAnuOLsn+x5vI41SBUvf
0SOscrUX4erCLZpmon64c2K+wza5UFq+o8F7sxxE0piwY1KwtTwzQjU8DwID
ds+US3zBG70LLPot6ATMVFfenfJIOGN51NV03WCKlGZcBm3bHn2aPQo3tkaU
CExytZ5OfEeYAsWUgbB1ULLG3GodLZy+U6cFT6dnnOFPbQ+YNaK5smYKmB2j
SEb7iW7V8pykaZgIuX56uZo5ZG5ewYBIUSGa4eXwNWadsrXWPGDjfCYC5K+h
dz/lephZJa7p8MumvCxKYGYoUfW7BfwHDhn7YMy05ySLZQOGESLAB7Mlmjpa
Nfh+XXFI/JWkOwCUMxhcON9UFxVOmOMck5cUnS5AY0snn5N1eE4CLV0nsxZ7
c9+GsgojJ5NiPt2gr9qkwnU2BbMYOZQtRpNsiOu9NAekqw6YxSdIYHiJZqOU
tuxPS8xlWGtoz+yrEvjXoQaOcpWZL4mumxjkeCqn/sbNPt7u7A4xAa2zr/ny
ym74mWAkV4b9ITbwHZthR6WuYamICnPZt3W4TNU7c8BoWFeTBz0v8WC/GA+r
JYb6osubNce8k59Myn7IWcna3kM9tZCnf5gh/LQzzuC1BcfRL6wlDQK+GSS1
Q/5sSaC0kRFEvcNmPM1Uwtw9nqWA/sTlZv0GTnNv35M17Pxw9YaV+RQ4ewCf
EB8CD6c5FtRHHcS55o/5OJyunxrzMOHi1OJX2k/5zbe1QG0uuMlA7F5p2sRG
lxEbCmIeYxLGf+hT/pYjXlXjG3rxgzHB0wikvuMTChNGbquxR/1eunBn2tXr
w94C0nHTll6EExgSw+J/dWFMJ+mb3jrwaSjHBtY/GhOXo2ThjDG65tVTrbJU
agy8vI7oTrLFv3jRyJVhEG8cMwkiqGaq5kWBnEPaxZ2na8IfQ0CFsn/xR/s9
XuQHvsr4MjTlfTo9XqYIcDmcH+mU7GWZQ/+ih/soYSuXg0icV5CSC6QQsbw9
ZfWpyJVbreSlpBEPlKHVgV55VJAFOsWVe8k1gspwBrpk4BJ4NvYkPbkFqHP2
sVJRN9JDLB1oGqq1bwzB06qxT8/uPeOFiLg3NxHG5o8F8oLdfL5EBLuLD5N7
jrtp01prH1gVmfDeMn7v42VG0qkeSHHj98ee0DCrunJLUiXqis+nzOlFDBoC
Yvq5NFjtTFpQX6QBkk32ItDVkXuEo/iC2eTjva22peMsGmlSNxviSs9EwDD9
/589sl1KifFhcSIW5SahNBY1ieo5HGFPOXZOsryPpR19po2FmId+mXU4VRqf
CKIhbdVNPabXOb6CMANpZUU5gP/LXi0gPqX8aQNTvXvNrmxCeqdjJNM5A8DE
TmA6yNTnR6ZfllbR22vr1bFzsx7+6N2A8bvBeQKg0LCV6hYpY5sZCz9wGICs
qaxnqYD+0XYt6h+qUshMNuTgytv3Lii1O0b8rgjzJNGISq0QiDTM5Fmapm2R
i8KjdcN6WPK1v/DkdAcOYa/kLdq7h7Aj2wqRmR6g7/46QXEtVTAU3ATpxOUQ
FPpIiRdzPV0OxpUtsM2omxSLRG0fr8zFA3ALNtiLcvUlRoMr/Yhn8NQTAL+Z
PHlims/pRCf/3/bUDpKKPwZz+FFAiI5y4H+G/dw+Bd6Xncn1cGIJ0tbaGww5
PgDkrON88+xE5NYgnUXuttqAaZRAui4xFIlf5ZGvDAh24mMsOjiMKcyHOkVC
oMQa7mTs2yeTHgS9s39c2jmzNzaa7uL3MyOa7vfhz3okcDM5lrP/40RUsBwb
jWx/rgT4gTlSFYTcu/t/f2/o6TK1IBb6x1ZfF23H+3nYtyjoft+okRFEFE5D
l6HJ52X5X7UM40qvxtZh+m+XgCTHZFBaXFVY6iCniSudo1nongi259X00eVq
wqoSuBYBq5znnOG/YqfF6xdjvSSQPkMF+2xeP6EoGkc2q6RKLxjcK4xmgvrq
fEUYLDFqxu8QjXcHeXuslpEQ11bfFhK3sKhMZpO9t1seMxPmMjNbTZRL64kq
DplwUguFkhn+sy0MVgPaWy9TNaprjk5daywogNAR6cMlNAUu0KDKn/Cpk03n
d29ZTdPJ4orL1a1sDXDNZ6IKN6W6P3ebKCQWmC9Em3CncYwbbUb1prC6dZS9
IuOUHgb3s7pSRdK+O55qH1MU7S4VSycYiPEisCPFC5/+Ews+G+Kb4xyj4mpK
0xP5zopcrCTChMWL0xdAAS1WVTNNKkIxYe8IYNQ74R4DCqLGadOU0eNsCgbJ
YFQUdstjaswqsYvh4zdwt+Zuv/oXW+Ubn8T6Ln30BcvmBUHPo79ZxB6P8vz2
TMK350tXOJ7A5RKzKUGLE7YSwi1PLAOFSA/AAOsPjCbPqopBBfkgouAXa2jk
rwDVSlZUYzgyBZflHpXJ2GViJz4b2DJqAxvbBBjDSBpu5dukTHBkNxQDZmd8
aR+EzsqW3YV88kksl/LIW73xwAMP5Ql+ed7M6kVlksD04gNwTWvXXn6htPve
HcsJBD8byTg0EQY9fZ8JyCg45oGAzQhF5jyD+UkcbVByyFooh8uJ1yZeCGsQ
3DW9ipo8UDyoiW8xQPv9Vt2xL3FOdc03z6SeZPQv4neqVKs6vupY6hHN2Qhc
M13B3ej4h047RNB9MYCCv4H7OGH8C4qdxsylQJprjxM18tTaDsPhCDZ35NP6
bVxAYp6IXyebImZMie6xo3+Px2RaBGA+mwbmwqB+fpZEX5nUrTkvs3mRQrPc
LZ2PjocBs7/JLgnvr2dPJG8i9YUwHgAa31y1m9oE3AgUmFF9ffsKPpEbg3dQ
EvvtEVJkIkkdRPqc5NziyfkzKmZvXtIipXUzZgq8gaTifRi/Z1gCs63GfI9f
3wC29XXLEqQQ0+NiQ+YHVT0t7dSfpZHiqbqwD1qkphQt3RM/m+NviPqSP/Rm
KHy/Tn79/FG8KyZ4mvc9PlrhmlXVhAnwzrPo2IUNwgcoR5tvWdx8YYOV9PQO
zw2ihqoXZzscEPbXlzFKMtETgXX5ZtCwmlUNI4kb7NqoIXASBP86gerySAHF
xsq52DsQc6FEZxLX07L16Dtu/SDYIL3sl8e4JeJ2N9m0ddfn2PV4MJgOzerp
JAj8lbuSb3o/Cetl24dV93EMUqxSI563VslGx4C7xIwXR2H7TF/Hkj6BDQhj
5gAdaNaJISvqSKLz8r4b+QRf1wuq73oH/zcPm9sLifBaeelEw6lwJz9M/L+s
k5E6kr81Ufwe3oNNnJMy0qcJ+jdd1zlnFrIpzmLRsKuLoBWjiW8zEblPxu6L
bNTioy6vcqNysf6nGjoyT3FSDFXTjF+hmgwW0ICe/BAKxrk4F1rJTqPfLoIq
ELJa/vjWMgZF9b0Vq+uxULM+Sx+Rw3B4ookkVbdVbMBQhkdyA6TWkODy9Zvw
doEvR1mH5+KPk8agWrJA99kate05n8vxsnLJjj7njOQKlouYevaknFwWtTTE
g05DZ49HaxOz2eeRLZIkCr6qVFTihDPitcEsZdQ3gmFCP1i5IV1bm1tK1YDR
MmKz6wkoxJwzviFCCZRNiZ5VnLV8ru2OOG5WpVi9bpo0h35HKtZ4bKi6dkf+
Xvm4J9KMI8woui1xL/4ALY2BVAYsmq6lYi+XgWehXx9410UoXmpxG7HEPLft
d2MR+qIOKE+5ICbhXOK/4R+k0mrpKo7oYG0vAjeOgMAhzuTIfxfLa6D1cWB2
edxKoYItyRY5WSF0N8AB/xwm3u7ggl2o4li4MDCH2V5y8eFYuLo0PFExtA1y
qNr9Y78U1IcPZCG5h+MRwSl8HUIcau8BbGQ0O7flK/k8P8szrJdVuj5xzVXq
06Hu8Tf4PHDXtlKE6k6Ioje22ZNnx4CXcD5X7ng4V3KLTm2pwma4y6o0TMuB
CQuwPILE/cYWH7CmfRB3knNXvpH3sK6O89Q9WRIcuO7DXRWfkQg/lY/I7qNj
sMnCiPIcARPtLCLdOzDB06mlOHloMmzja4J/OJ6ItCz1xnSgSWa4n9FRjjtA
YUxMlltcMOTNIVu4ORsVdx0Ww7L2hgqXyBxwvbz/5LrGY0Mhj88ZrXIUkvlo
LMDwLxeG9AV3JdOj86XjgQnNb9MrdmfhRtlX5RGPKxXUGFzZ2VUvOGeT7E7y
0afo4X8DD0Bh73MvPivIuu57orKUnAhYh7fr3EDyxuWHklWrG/ZePW64hBEM
YSfqszDx8Qwxu7SlMOuCXUK98wnLWnoLuYfUyyi9drvuw9usAIrAvlmaB1LQ
2jbwbmAbzFPg3VmMfPL2/I0m6Y2deM6K8FuIQx+yVHjjf8NRqDjN738gyubV
x8/2TU5ZrCpRy4BYiwOGxgwnhqbGF0gdB58gD0dJczFaj8RRyomuoUtty/yo
knx3ViE3GW0ho7z1+TfwXHE/QMx3iHyTxx3gC82cytOQNua9zItL68cl1Dg4
YYPzrd/6RceyHv1T40svTVQJXDSOoU8W0HDxRq+0Qc27fLqqOvhiyIEJ9JRi
YZ3Lb8tIv34hGv7Rpfj503K14FHfmx6Qz+dXprMiE72kQlOxQdHJtikTup61
CbMxo9uxUXampp9feppD+FdBPJTtlPdqbx31xzsrW2c4OZeMZ+M6mssJd0Z8
LRtc1T4lMhZpyoq2UoXSzr6gLDDncDQyPwAQjzdeLHXREWFHVNnpjjnjyvNC
2oePzGkd6fc0DvfZLHSO6DDqUI6j1OyOTY6KlRjzelHACMkHyOq0fI1I4DUX
iyIuWQ3CmkoprOewFkv3koVcrQXHjxKswfo/loLGlsZuCdekvRBSDK10ZlG9
FpqOls+H3+zoywzLxWCO0VBVOl2mbBhEO4uEd2Ig1/StFdyrg9NDiXTBPbkD
AwVNpxLtJS8w6M+xFH8ph+zznlCB6ubL84kZU8gE8rX3HgBJu8jaNs06OzLS
KBurWF6eaGFGwJKSa1ZfbMHRfTB+XPiu4YE1r1jNwEJ9tdcndySmTHSBHFPE
ywlqHmoW0+WRzrnfUD4x1gszQ/31e/el2G8/OC/6vSyKlu8vycjNEV8Vd9in
ciF/xp9pWhCIl6KJWpNKDvcq5/G+JGUu0VqesTbqrHmpqFAziBUUxfYU4k1M
rpEdVT+gzwSbU+ef+8JCDI3dHhg++qiMY6V2g5kdHvbStaRkE1WakGdH+J1Y
3mJ1GYCR8O7w7vRtmC47tO1xpq88nwzOG73fTooXA6mRqZUF4udJnODinuXz
f5MoWfVuodzNympzu4+nR+1f1GqnAHv3iGq8QryuRefceEDa/YINbFfw2DVN
3VzyRHke1QuuwwIAA+2OQQglglgX8M3VuYAChZ+EAqvmjMtu9UNmpHmXdGfa
E0/aIF5FaIKF4eb6T1hJDZb3Z/DXDIVabdT/15R9aMMN8FWTpMw3Hd05G5F5
Ct/Eo4RRyGXTTt7Flymu3EtOcRvDKqA9BJ/NVRDdj1kThUXZnE5ASitRtDL8
GB1xX3HZ17otH1xJUQV0toX0efv+qsgr8/F5lRQGcJBCJGof/Aqcxjins6Nk
Wg8/d/ZfrIVYcGv8GR0Evr6D24SDyZmvDuCYbHNdfiuRUcAu+0LiP+FqykOx
dnRVT5JIWHccf1CIyCUbJ4RayBBvj081ZVGqSOAcTt+Ik7wjp0w05j72VzCV
JNwaKPd1RVoCt9YBwipLRZCMBBh+mFEqg2/d0zcgAgfXVliI5y6hShmd9evL
6xkLDJDiBntI3wuN6TEOMhYeNyGeuZKobG8haIefO15cJAAanBO8V3gZSr9q
51TyoH3EKpzfzT8KACImWmHzj/X2/saG6+EPDPW+6sTBZbyeUcJEhLyT3FSH
XA4ArXHmkWQNn2sZCJ5gwg7tTBLahf9YFrBzmDQQb3jTeRi/040XY0Xl+5B+
HN7KU8v+36rhgUTLIgiLUrZhFSxsOJWKazgQf3S5aYeBtC7duFLOIzlJfoay
y+6N+ON09QDvXTnaiKuZ1tggOEV++nEhMhQ1KdW7UZzsbiUMsdbpySKCPsXc
5xHyx0GFzbpbCemZMLOwTZ2fGR+eXRSWPwgfX9l7M8gXr41UGU4PffDx5/ze
fK5JWWDhRwPJqfv1ilrv+xqmPQLO7cx+Q7CxfsmtRVtS+HpDvKDa3KbuyxFK
pusbI3ywUmgEKp0+kixP1dbf4zOAWWTjNXweVOHed89ID4w4w/OOmgp5N3OD
i1gMBlTOt7rMBJoUEmPcfRq7FvsVRo1L5gcR0GHvBr13P0/7myevCPZ7O9MS
Z0mQn2Mqbz/wPpeF6rJHw4r3bmwGajS5Jcj9uH9tTJrlZVyYoToXOI9Xf+1w
Q/IxW5SxViibKMRSqx1N/I8j5hwoeIG/23bipIFmgNev6ZUVV9j1bppNPr/h
uhJyJekOmxAXaOEeb2vdeW6R1pc/a3ynkg34D+orhxpPawGsBMg6Xd7shYhb
6JRHPVk+kIqtc/uqA5QUGXpzREN9RSIh5Eq8B01JcKZegO/aD9pa6lNo/MeP
iX7Jb0DMWz0cFyYUag2ZP2CJ6omE27mhnanj8iaDWDD5Oh4iVYiuMZ662lxg
2TxnFF2lOpYSMnIA2zE0zCOqoyac5/kw/HAD72PWxwlsI0xD+L5ch2PPAjCC
gw/JClASEYBLrpBvm7wopfnYhMckq9n3JWFUcN1AZoCQ83hgrUj6TFtQyli1
GQ/eh9cclnam9+EobtcayTw767aXMMG2G1Jj/WISvkpo+Fa6Dos7Ct0pOom2
CzwpNFxGH1bjg/Gzuw8e6YMtEqIPjbOj96BQuzp0a12CG0eRTjzGfLwY6SvH
RNVC2R5ePuMusNwFhf6a2Uwxvp+F1/ySNowDNQwuRRIyFdF412LC9dIqrwyZ
IUE26jwalYEcdCHkbhmZAYQfULPXicsp+ktPDrxTCANRpnsfHur5eGTs7Tcv
UfSLcaiM1xI4pw2NjlcM47FB6fQIBEBSCPLGop1XXMUcHhEk7Y2tbPsTQXO2
Aro5ER3VidEQyMVoN8k4U1m7H8r2aT+gq87mYnkFdHz3lR75vJi9k6sMrhua
5C0VxC66oog6slw8g5XsEXwSQqqf0yRNaArk6OrXE9nsftN6mJ71FrI9IYRz
Xz6EjWivKXVTeUX7NxqqfSEvNxLoE3WudNw/FvRCnKXT8N4M9WLYmWoIkAnJ
37VNji+uQwb4h/Xphbw622+0NL+UT1MssaktIdSoSp/G9xr6EyijZXE2/ja6
LAhJQ7hLZWzM8s1PIADeSfNcZbcY4QyS3NK4bwR/e06KmlFwzRxETa13bc1o
lUvGrYNzqIHFCko7rWI1B995aG70AeRneJKeHq7alOf+BBT4owwhLtRDazzU
bC9QBB37bTYcoiAqJiICVfadJxS7bXikOb0kL6+uLVlp4Q3NWC7J5+i0tAs7
XcaU+lrwFJDKPErj2YF6M+vccaVp9ReiNJS3CsjZmCV3UCJGIBbbyg+KKPDu
AL5Tbl+1dEvUzGAXfZ3CqnC+dCU6PwhWBGMr1DFkjsz3rBb4MHYLsNCF+zi3
1E8YXyxEA+qJPIs7QSLL6TRyA4WyjgPecsTF7P2kjZWXxy4j1ZKQ2tv6Glns
tzEh+UZggWuSfmSxdia9y83MkXs8wbQzWRMFBgQRAmKiq4ozzXJ77E1KaPFV
bJQ7YCxvoqdI/MmWrvz4hFH17lwHYfmMS006hFADryxt7T5UOWJLcQlOkdCW
A7HwXLZqy76K+OJeZJQktbKWQ+jbytKSEq+sZpgFyLZCUBxzklDueJbR+YCz
/FLtrtGK6oCJxdmYiC4RmWxOayg5dGyUYtRiz9oAe8q9ZIQuPjs2sgaCbIth
5rLz1JbWSdGBhUvWM5dQSMDNroKPHepEDxO8XtW/1Udlw9UxDvjHphmW2wkx
2Q6UueSWdXUVOst1S+vzoECYMwHxXI80UUa3tHZe/4yRQlKLnrMth1qxek9D
SKcB5ikrkryYAkMSy7Ap/XDNfZIsmurYuzJTLE6RyHij3HHjko0oDxybSLr6
19+n12yLYqRdQuMZp6AtNdJQOzo4l7bbGthkIFHiDZhdFnAUa+LqYMomTRC1
R/KlWET47ghKw6ZKWJIBHuj8A7NPuioM7eYnBdn5amUq3zSc/InXfFm61z8p
yPKx+Vn1lquTKwZR2LMoJzDN6hYVVKG4NGdGzashKRhKsLUE6adbIfb+QQqs
TGJAbvUbuS1ksCPEpRyGT4PB8h+tUyNxCIsDaR1e77rSebGlxibjKgC0k1VA
IddCDyoOshxbDjTMthmcs6CMlLRHT3hRCv6AfpNruxGMf6S+NXNIpCb5oDoj
ui6CmStlAzfHZjirQ25jpL9YE7C1nIyh7SGfr7nYN/Pj2Xx72sns9Adk0pnC
/geeD2U7dytZYHzm8OLcf+QyxeQIpOP8qO1gNIJoxafTrIZhnTU4rcv308oV
TxQm/36aKtYU/SQANcxpXzsKJjLdh4zOVO15E7FWuSpQu2UpoCL+RJfQ0Pk1
/gsTawy9ocimuQSJ2W2c/oUSJv7EpVU6ruWksuBuQ4aOlmE2UhpPqOXBb4n5
ByNc7fkBpw2O2mLU//36O/+eEk8LJq3vsciPFbc+IJRSSUxlyb6oXT6mhXqU
6GB+2VUe528VlFMwzri9snqPOeRWZ47IK20racXCUpyTCagN1bh57As6vjVK
BUGAGBLHCaAp2GVx9rQJqyHTfWuru2wUz7fQmwEBQ/3dulqFmSOkdKEhpSHN
kqePU9RTs15usN80jTxNAK1vny5YYeamuMaaKdPPRXbvVB/O0fNd4/XodS0+
O02F2LPq1NehEzT+acSDeCt9jHRmYD9RH7hdvxY0whw8gl5Ue9IANHPtVfUA
HySNTPbhYrqhl3UF/Zmo5eJDZ35WobW3TIWtd/3dj0yo5T2OlPdxg6Vh9YB9
C1d667XDBSQLTvE3DqpBb5kIGR/urftd9JMrX9vlyQcoOsQqqQT2JHSlT+Id
v8EsbIr2ObmhS5KZeZShGlA01tOYcjlvfEAeEgfjhMA+YntRRPF/7J/Q52qx
13nrvu5DBuEgFcrE6+MX9W5xhY47l/wSRBEgP/fuVTE0v/gnOOYVzUf67wuD
HO3iruM8xP693h5dpJg1B2iHnU13b0IHi2uTvjhJNg1+lBHN64MJIcS/ENvG
HeBQT+ShDg8mpwRm/SUwX954IQmhzMU8MHBhoXQ/MmBv+lFqrj2rIw76Xg1T
+hhHc7LV+hWl0q42BjzBND1lvtoAxTUKMGU+Lxge1xuV8JeMpHdxJj0AliuH
05ZbVmu0LbuCr+93UInqoBwPMn8lW6DKn5Lh/b20vluESTJfc0LDz7FEKZGt
zL2WOEPQlV8yaji6FT8sEJJMEmArxagBYqJZ8AIWDTrWWcSeL4bKfTfBsJHR
rhHyKAnbmwARsXEJCEUc/vuhS35K85GTPshqxUv4KwcoSzCxT4I6jvu4GOMu
kkXxCTyPmtTPbyUZR3dUJ0dwFWiAc2yJp8JOWrt7T48GNHh/mh4Ba/yE82mZ
0mDjIcqtTepawD/Hj1dANtwTYorNKlrHMJyor/ZC221k/pn0szuDdp38EAHz
r9n8Q8ZsmZBkOIuD+HPweT3wOWmYDGUSOae9AHV10SBDHkZLJ9EFE8QINhoD
db8RLIZiu/vdAXU1lSxN+7emGuLyO8DNzDqv64VC0QpwT8/OkUeo1Gb8+3dI
ZUVCsKXmbB2phrVPyeUDeKwWcrvfgyYBZpuToQNFTnWl4RsVZPYAYyD2EgsZ
xc7MIDXepZ6LO/Ecf8h9zdRhfKS9YwEWgiUOhXR5N9M1irzEYmQZDYsJLaPl
0SRY+LHOZKsxzRySMH+K3O1isXxzDWDz+jBWAHMRSTv466s9W6BsmjH1fyID
9yVBRCr1mGtbUo6FEKjvxragZGbmx41JV1B+0jkJsufQrUN7yNuRcUaKgafj
lGG4o5hKlPIojVnaFhznJYMiRloFyhv1IbGpQRAEkYh6hZA/2yE3c7wMBkTo
BWh3gRddmCoy4XrZJPSQPmirx6tPuCGthz09aVaZyThbYn8kufVatemkjq36
dXQnuKh6wxjIaJPzPBtmwRMDToaKsWFcYnTjqro/fkNIRiUyv53hhioZW6Uz
pblccmKB5iZgQvDyF6GE4zfxWVwvZEdiZx6lHt/AQIve7yRAiIdRSnXVDfH8
QZJk/Kt/dg4HFNjy2nvNTtEVrBLirdAmlx3K8HQrSvKNIMxD7+aLribi+c7d
W+dGlsn0VkDPIKn3BoiikjUHgOZLGeWMXPSIecEO5/XIVRvKFZmXQ1TAwKEX
P5CJKx8oMefO1QP48R7ILZDWuw7PXyZMzRWs3oCWZzzlHfsHg0AFpvl+k+iX
M+pnGWydAepy9CZUsoeniyZOdfXOiF+/RaIlog9uNeptLhM+32dsQlFnthZd
uEzuDDKoun2BRXu50Jk0ll1MX/AL3fq5G585ZwWrQXLii6lJ73AxOPOUKvnl
mU4TIoiAGgzPFK/nJrCraVB2AjOvleDVU3mfpg8es+bhOenOgu2ntEj9Y49d
aPyQtkUnuckOSA39ql2dkS8WQrTBfwDsXmJpE3tfzf5daAkbxnxVSddbK4iE
mvUdnIr7TqfFAkuJBgFR6Nec+nrqwRk523oiQ370uUfsFYQA8nYugT6DJA/Y
2l+aOndRwkfDwrpUWCGPKEHUw68qYejWSc/Yj9Hfc/0IaJMV3d0GsXi7xSrG
5LLwTcnH0sFjflrjN073Xt2adq6awK5Ijg+yAf+Kj0uKKWwTlf9LXo+XGBuB
YJXIwFJeL3WLyCkzgbK7w2CN0N6uBSirDy/xpiJ0eoED4M4ar6guPUh/PTAO
gpyuZ+8/LsT0vc1NvqYl8tAS/aaQePy1tdSlmHIRPC2yE/0DugUU0qYg3ieC
y5zzZMOThhW0HZ5/4ayOPbY8WQ9GkNram0vKc85rXGL7oXySKccg/hB4W8Xg
EDEMjB+2CIPULCTpHLU7nMsZ0sQNcY1wYB/7rIoXwg2I49Jt9CNLaPMeSfz+
HIOLaiV93ykFULj3dvOcnqktTVcEoBSur2PEWSX8ebJYB+OcO8JoybsqXUrK
lMWKcINfs6ThM4xxnFRqzF4xXOxFhYAXiefVDqHdleq19kwHQ8akuBDAmo5C
23Rywn+lYIRb8+FK0JabC4gNIZCfhSwXaov4oqPOvfV86Iz4D56E9tP8PELp
55/6Tq2b5GI/Ev3A/cSkkr2gECp8chbqA8pxFOZCwG9XtRxNV0GGxT94wfvX
Vc88qGkz7oqEhLQer7JM5PR8rLBGvPzO+7TDfzT/lu7cKxliDEKBzp+LPQCx
5/LJDz8fy/l0UWVQBknpfLCQVRDSyZz/7PTsAryOEawHylvMF4bIthFmo/YI
AnBZKAeOV3ppGA7PbPxD+DoLu6WwWHutKehGwFy0OI/RHkltx6IYn2l86QFH
uJyzaBYtOzymUemvp2MD+SZNsPY+60FqrRtlDnvCsJLhTawd/Pia/4erkDHB
EsC2Yjd8nNVcOzy2yliBZ5IsgBoFnFDo11lqb6whDgGd9+ZOL1M1xkk35BA/
PzcDZSo4s9g0G7IPbLt6IvP87/OHNHyyLCjJB99h/wR2yDPuSownIJNvh9Hw
Z7uVT14GAkhiWm2sR9olA4uaD2yCpHQM8i5w3yRbq8NWsC4RtFUv27l3CnQN
ONJM8XaLLOOzGyBxLIKLyctGe/B8mguN87JDx8M7JTJ9SJqggentGGkwfZel
57Aw6bZw5vCODKINxa/TPYbZezbQXTT5JZLNXwhKT/2RSTH7VCd/WYy4yDnz
F5jZr+lEZkmAMEv3cgmb1DuI5uVCNb1w2w2shmRoF+QWZiqTF+sz33WVAV16
aQhgRKa8ln2L2xYhspXzJT6u7kl0fjX2lqnsX8+xz5dxeUJJoq1UTYzF/UrV
1wk+gs7qThi6UOvaB7dgxKUwP++WkN0FvkK8UOBlI1GI8gSPSyGDZeBKe1hu
bR0+j6A+8hYllu6urKNonVF70KEKai3hBeQFU6nIyk+3O3wsxNrcpSZxGJSb
eVBbH/vKFOPPC7CGMmpgIt06wvWgwB5YTMaGTScWgH4uWO6f+Ub5tGQuG6kq
bDMRIvuSj5Z+evFCGA2mBxmH7nmYSbcaTce1bbsmyAku5VbxzWiP6MHZbXW+
QM8esbSVqdxJO9+DdsCDnhRYnqxQGfTGQFlMRq7aEiWTbGkHx2WOC0ne1qA9
iTFYP0y9N5VcK0VwzNdZBRyE3WNJSD3bhSgXC1NhXaAQSZhRBNGmPk5A6OHS
jQ341WVI0ebLnHGi2reAvp7xggH5PWi58fwG50ddRMShzcsSdWf0kmnKDsmM
SruDouNlolkvZA2FWqzIJ7IBx6q1mCXy+g7L3CsMD5Pbd6T0MjnoEVU7JvLF
WNUs7ccMUGn1ldJU0zs08I6vo0NwyXRDCumZrbEMdoNilOcx37yFtDm1Vgk9
p4sR8BXjBR5rO+r8T/rAYQ7YOYC2eG0j2iRxkxw1QFFM/D7doXGDWzsqFfAq
nCNPZ3h2tVnwg0lSXB4GSqKzGFEe0K2qBcgh+9zN37380/KM+1rL55meOk7I
4gwb8sUoEbDlQEYTvOwuEP1Iw7PWkojx7pN5wVKH57P3OZ+Uk63BqnlXEzaq
nmc7sWl49yAZkM8KtN0bMwCTZ9eKZNG0LIhdmtk74bAMILvL/zp3Trz4TFc2
4DtfgJqFjBT5xWFeBWeVcZo8xhs6x+ImU+V57I7pN4yf3NMGynzN3N5+v728
gPuyV37LP48uJ7HZvMm+5mWSyiwg93ggcQPZKvgdC48mwFru+giOx1hCznTG
oD29b6ckrfM6I9/ZUe6Di+2bw9JZAFzIKpek4vp6aPK32ro48yPE2uozGXD+
m66EZhFbA8KU/jvJcJbaURRKD8VXz2cOESJyx8ib1VS4lSN0XMuO6wJEw3Pg
PqsFZLQWbDscJCkT0yThlq9z4rl0u/lKxU3S0M3CHsCzWH9gMUVyxdgNbokM
HQlsLCywH3n5iZJCa0DOGZW6UmSO6LyXnbAvv4B4ga2XtcMs9ZW+WpYT1AVm
t/ig8RYNdmh2BEJvxk3MYNnQVRJmehPEgBfuwCUBSudW6bhUb3CCwB1wMKBZ
7tdGX3GkZgmKdyodUI2U7GfJb4rzynWa7CVCr+CPHo/U4qYe82M67BsI2WfP
AximOHOpr9XJccLCmQ8bwS77q5KFLBexzcSQ0eTjndsDfmsb/L3a3KckOAnw
9o+59aF8gfVq5cXJi+RMZdD2Ru/8cfaUlaPm/lrPHgUxKe/tJJSiSQiIcaob
c3VVUAe8fX0Lp/nq1aC9VPmpAUFwyVPliG+A7SmQgM8lQ8uvXU3v11nao3k0
HHOr/iATkkXnYISDyOpNUCbGEs7H0WizhqKObc/D21xgAbGaHJwQstVXadJ1
ck02bIruKMtA+UQfZ7pQSKqYzvyq8f1NaAx+oMLzi0mGTrGFIWNJaduB45ws
wYxu4JZiM/WNhl5AFJEOk/kO959VQNqsm9N+xUAeznlm6Xv6/9Q1mrbG/SXK
0GzMiwR293oJfB0bQ6c1aT36baqnYIP+l1q8G9rDVN0Rpyvfb+FrOzy45Rgb
tVLq7GhhHg/UTrpeAulS8H2YV8enrv6cJ1B2BeyF9LgeX6U774+SJ4JSprJ4
AcaogI5zWdIEPS1pMjmdRF/i3UR0h3RAAMWLE7sxuFCcp4ebsWIdP0Br3P17
b5KSWFx5wNpjt8CwySNHKlFbJ745wfW/DqICns/ObtiO4uLjjdkF9FiH8MEE
nKxr7RVMlQ5wJX8hzzv1Y8RLr6BuqPknycxLk+SpNHZyTng0guQWl/a0SvCt
BgJhW9pIG3eAZxla0RhPAMx/7PfvowH9e1l65tJoM4l5pFDMZVpIz+UArplr
5NeALkc8O4s7CKPnEn/n9/wt4knqNbitgdK8mtAQ4TErDm3u7itocR06zrxQ
c7L5d1bwxxpw0ahrZVQ/wnikk7KnWPKvPX5WMHLsbFckxvMRCUSWjhNL0gzq
5cJSWC04njabqTDOPaKfqfHlR3XK7Ki2fHcFxdIViJP/lhSV6qdS5Ui4H7uU
yu4xxzLUmgnShNqYAhEeYmBKoAyxl2rGlDncMaIxSedHWD+b9/m1Mla0dR97
h97GLM2mfInsse6ksBstZk94LO0O4iSNcvRXN4ZU8E5Tvnqt7IX3PrcZLSnf
kdJBWGAP3nmKxeKE3HXNhSiM7hq+qhUSuBCSbfbYB//H6DVHJMhQzgbRBmUy
qWq/pn1vecI1j3JghNA48tG5dDQz1uiIRqvofnkvlDJAkrUqc8dT0iHewH2W
RXeDbarqc1bEyjCm+DqELcvsux9sBmDvtpd6gJsrnNp/YPhIKpSCrYyk0tFL
i7rbqRquEpdNDwIOPrb5vmeBBEfs+275FecgI8DF/9KqRI1DXTcUPTS5IC0B
BDxmd4oSY0/bB7Z0NNcLP/cnOaGmtccEEPbAIhaz/Bf8WpRFkMp8536ockyB
Qd6Cao8XmzVq0pERiO3boPu3jJwMcvknRsTn3P/CzvPp7cSUTP2dHlenHC2y
HMH/uq/G+NFz7Muzs6Hb3YA6lYRP9EYGQX9XUG0/rZuO7UpXarhd8uWDYIDE
YRaq7CBY/7ezoxEbke97nNxcS0btY5Gxz4eGguF4MaAtASUH41C/xxzq46CG
4B6AGdP+gvY/MRllOO+FWa95qcsM4080eGa8kaIbeireZmFxovHgLnB8pNPr
S6XBjuMpgSbhkW/qFmqPSbGTvyd6zNgfI8cYmz8UCP2tfj2Zp/5302n5B+eJ
cgLUr+q4y4qTRWbAlFZKjoOuoPorQsCHJSfdkxGqSzsFzPWDZdakvfUthh/s
Rf7zIX1GYZY8r49gOWZUJ+kdBoLpb0/WL7zRQ7PMvKeP1E/9wlc8Mb3KM8CT
CHPNGFrOxdt+ivQOd1NkKGWeGUvSxH9PkBhnqSciQasRvey+zTjyfiUDZunb
W1locYJNfNZvGT4MIJLj6eiZJ9FYgBTr+TyNGYBiSK8RvzgN+QCh6hRywIWi
cRdxITaOv4ew/LDw20vfRg3R3edPbrQbGk5+3v7NvnHzk7wNhi5K6BKBLUn+
n1JtakFIm11ZhSxZ5w+8p440+I+2LuU+JWAqajXmuGiQn0hatHbR1T8T3jRB
aBAbhP4dc1Vq1p0yyJIRpUe9TpkA5NYzuvx0i+bwd1K62yaIKsl9U+/MxoRJ
bwm39t2iUknoJpbLnxafd5Y+KWsmh5+Ex8Gxs02bpBeklp3G+xr3ynVvq1nO
LLN1ltFODLr3cugumuuMuLOCe70GIknuzE/NiwYfrybbgk8VmKczDNxs37Pi
qgiIJpoghK385lkatOhZwxlUUsZgWw//EluP2g5m2OUFJ5mBsxS7THSb83pK
fObzoDXiMsae9XCmXx4Avg1F10tIml4wuxjs5raNBT1rqkNQ70YaLlruUsqr
6TlCsE7wvFbBz0Tr/jxRfiGjCXaE7+NbJpk2r2tA1Fu5W8SrmWasFClkEw6K
dsqClPEl+MtGXzfSUgSfXgAIWSyTCnaslrV235c9C129M4Gz7NYRMAW3LGMH
+MXW5mAAcj9YCMMTrI6xNqn87uopSmAKNWkZmOJD26wo+oP1j3YHWWrU05Is
nIbUx8G2G3v4/SAXL4nyei4PrOmaVCK96UJETNSDRm8Ji/3BakO7i1Q3eiRR
Oz8zhpe3ebq4+mtMzQuZvW6zktf2dlcfdyVLIaKrSH4rYZzdQVax373gINhI
TcnyqYCGSCdouG7bRnLLUiuN2AyklBxzRxG1J6PI02n9eYh7rXTLX2BMnxFF
a7w7Z7tFkmBUL6FPJgLsWNTHo/OVqO07Xf63kYdNcn22C3DBepEa5JPypCiI
5KwahAxxqADz0S7rKousNsxp+lyLi+/afJ8ikGgAuWmSodh/ZFgAx3SlhCqt
/IaP/65R5LDpyPwHfTV6FsrJAD3xM5c7Ww/XWVmIaXcXKbS0lITHYQnEwWDr
QbR/4oKjAb/MIEDmZC8GJ57jDaGFK+mhjHOH7CJqtzZsb24DkY2eVUxo/DfP
PtIMi5HVHP6d40u/MePEzDxUWd4sK5jphcrUeNM9gSd9Qf5gcQd/+GLg2dr8
J0GAxX8sIry2fVIMG8l1Den5R9gi0OEfm97bbQC0bpX+4RxRpu6bM3Vbfhp5
ykuYrV1hGa++xXtv3sf1kinExaOQG734ttI8z87CwcxhoGoDRqTRagWGG2x3
2M49+zE/YkZTjalwXACAS541DwTmXEYCh9YwlwH1G8y2dahZ5na48Kdl0QIF
CzW80SbQLxMKSyX4BKzwH3I+Qdbca6XLU6XJhMn8aVAACuFN8yxA1Z7gUvLV
QIgo7YqzNb1SoQU3BFbIulrSdsS2HlSvhviaXE0pJe0d4Np7TR3slRiuRNKN
UD7uRw54ZXCEaBw307ZuskzuoOxJMZehb9WTVX+HrJIddg6ulflcg7AY1vLF
Uw6y18zAPJ5qvFK293NSK45EFP4kly3DYrxKj9ivbjOyW/IOl01ZIy1RWD3r
bg0w06ZJplPqd4B6h/IjzFrJ3TaEXJ652NnLx+7bZFtsEua+p9wB37szoGtN
bOM7Gea9k5YeTtJJXwSGBmqajpZHWDjJaSuN5Wda7AadGdLPvd0bZ5QGUu5l
TsXwfyw0uHswGX1MLEeeeeXeSRVNkMNKLjzahoE8wfJRqOXkOdQFHK2EzhC1
3YndEuysA2nd0MVJ9Ya66s6acY1C9vt5Vc2JttdKLM1obwtJ2iXncnphfRi+
VihtnAcYqnTTOOriioAO9qDxx3zFgB8QmrQPD+RqIOwFcRKQCj0QPlw8EDcT
q5dQ15NDrUGJur2x/Pl7R4hWlfpoYDbFOnDej0XR+IiWnIVYftMNREiGWJcV
kxPuIjPYrTNPu7NTUEh7l94e3q5/P74hx40N9/qH1skCWDEXgyx7kp0cDICc
SHYeeBV4cDdppby0r/bIADOjb72nGCQuVID8A0fe9+nxD1hwpW3Sxvt4XrdY
oMW0w181VKppp1+H/M0aK1Qwg4fIMhOKAw2tip8JLT8MI6eyl+sNg3i3JMPm
1OIE5SnAK5TgDhAzxy38hyIUIWCeiwXBxQ9MPsesqtABanwVCALv3jEiA738
hJuFVVcaFJ2jVDBc7IZtjPqZSLJuNa7ZiTeZZ34+SZwb+nvIncrobbDe9LzI
xk+rA2mDQx8CcoCtsVJwgLIZCz4c6fvcyCxl/w9hp3TY1MfV+zE8/rT1bhfL
qzYA2SZ5ONBKi5/LFGVIcjSZLUhoQUYRZM0sxFTUuSZQdtS59NyB0m6mqhpZ
JMjYZwKV7Be3Z+2AwWgBho6d6mj1wk+xlNxOqyl9Kni3AYcMByEJn6i28uLi
eHaFaAYQTUmIS9h5J69TZOclpTtXDIfh4eiaiNRCU5S6SCAs1hy+3NVNlfPH
BhpZjUm6i34/oDidgPp/Kr46KtTkJuFWxJ0GTdDUxJsUY3ouASZ0462mZG/w
GGbkF/QHVbNKYu1CKYLaK2xvXruLoV2T0qVvkBFKUcUNbl6icfFUgQWup3uR
3l0fEL2fp4owgooM4ZnwPZEQR7jexBpRZX64S8NcGNwCEullQvYvZNEAVaej
6M0AICxX3EB2AwEgHXo50XXWxFVx7h8Dk59jiWvRg6/cmSb0w6O5D4xqOSei
LN/y/wiWX9nkG0K42xl2G028ZCDV4qQCMiG8Aar9NrmeDT7+FIFFSfUnWaM7
PyOmcofYRWLCIwGOIsqeyLNVs3jFxCnnZLkonIeDufwU2gSmrXlboRaC2R7b
/MQyATGHvRS+Yn20ebcEcNVwsoMVuzU+MLTu6A/fq/bZssL7LqYfxkMoG0Zs
TAHM3z5QCfED60NwcgUpAqLp6e7XjiIMorr2r3NvBBgzYoGxz3bQF0xWkFAd
xRdqgFxlwaA2Gj/Ylpzuxoa9X2mgvixmTSR309Pvtg5IGKN51LdInh/YL5AE
sWKlAQBaqfUoK+McE6rtYtvrbij5DyHHlSjDvN9aDF/agPsBMmKuk/JOyLqJ
R2KAikKhHe2KumP5lCPxicdliocmfJ8zLdRflZ3v8q0Og21M2PpUXG16mXoP
wkmOogYOsXvzg9Jxj8KnoiSMo3bEhac43poq1mSJR6aMbM8MmajQ1SywdZUf
b0/vPA8ERMmk0Yk5w88Dr6/sN+pVStUaEF/bTVwq6BLNd5m8LDgZhhFjSeZt
upVMcHl/Pyx5u0Eg9ZfYHbHkK4TadvMMeAHr08cL7i3By78s9eUKk5m2sr6A
nxbxFFDzZwDEwGsQz3VcPc0c7UnQHZtGr0TALlccQbxmzRTdmTSRRKM7uLhb
1t4gJhx4jkwYi6BIHnBqh8izUaSc1cKYJ4VRiE4G8EtoK+n31zEC70hzFoH+
81Y8oz68hmCXGkzJIQMqIJmsmMaI4BbJd8hF75B4SVETSVle3WYNgl+DW0Om
/llV5/2EcN7u+JC9PeM2+6OP+lyBFO7KftAGa0ZmKVrAweoXWa3C7n2MjiCn
MbpsIdXjmcM9izhhvd2a+4Wp7rNgHXbdiddQ1sU/VMwELLMz84h9ROkgKCzd
+P6IbX57k0yOPhG9zXxNIKdWgycoJZVwIb3zz7zKYFwbJUDs2Cme8xuTIlAj
+n9gCtz3E4ZWPa0XA1DrfK1tuFATmqGji+jBIDb3fBYvDjfjy4P1hgcD/nnt
3atZge+JeabDjywrDnPGExehc0xEHGJ8WODPUSvzoQ+uWbCqpIVPsghPLuyd
DcTyKecamlOMgLhVFcK51R1Ke2BQR38MCgo0vTrlQpmX52rvefuHTjB9Hkru
j6owiUj5MvFW7xNVOeW+NxSQMA3kg7P5/hjtGMabTpx4mV3VaZGrrxLjR5Va
MVmOFrCt1H/P6mvuqG8Qo7MnbcV+E74eu/jDJQ9yj96n38xM9T9Az+qnFLtQ
u0gKUJfkEGXpmbL+9OfcXKqLzRdSbfAipGIB0sMfT9mLkvkb9hOXBoFeNrM6
o9K+OOeZEFPvI8UYxULf7cX6388zgqfAe9rOFYiqEafzsMal/CWs1dEOfvor
ZVNGDJMUS9TqUuJD0oFVexAiA360fQ2pdge5vYGhOi71gxImVbj1rk6un8Y1
YMDUlGvChNy08m6Ket01zNlUnbGrl3NdX0X1gQjww2lDZJe2IKcFlg8RI9rg
9pCG8E6GBjSRarUnIJ2ghtYVNejEQG231eYEJbrnAzxhkIv3139jg+BpHueS
cThJQ0C2Jop8VXLjRcO7C9k5jQ/qereI6/n2LwYuKSAn6e42dxeibcK8LNz/
cdoyMdlud+/TxirnABbwkSPO0WlDK3IsGPhGHOH38hCyV5S9gHskGljV3pDY
TNEFURWne4ms+QCPi1SIbMtFGrS6J/dIDJt/GdjIEFAgKhHF+Jvu4Nmybmwk
NWEopDL6JYPtmK5H9p3W5dad2K8Y+89x+QwJ/c/OXxvLiIxRm5VmrJDDvQRy
tHb8TTyLq7E9EbNoIrf0EyBGaXdh+TUBadr2qpkGYiMhAkI/El8IeBwHBPhB
eTgLGC/8EFjFLgcYd+PrAzGObUyk2HIXHYLyCN+4hqvGRO+K5fmgA3BRw27P
UrGHlbKNvOVq3CcEpXEeXzVvn+TsQMOkeg3wcWnkMSXJNr7GHGtFBzmetYJ/
pRPf96uIkEB1obG0RVBnhJwgykdupKuB5OnW1ONpQEp1GioDxqiql5tMepPB
VJw3+/bUl2GnnfnTSLVhCgc3JVlub8GFRHUapKLa8I47P6ZYykwGmaiFvHge
usCyKdeXzJSGqzFphzH7x302FrElgzAD64Dypj0blIUDa8i4vVLvAOQ1etOz
fxgg1cRbJe7+aSb8GKBe2BMpTKHs5br3MWhixLKQtDSLKFUIsR3qwKUvobNU
P5v8iYNoobtFuqLzV3jzyTws9t0cR6sV8uWy2F7ZW3QfZzcjH8pvgS/0KBZe
I1D/RXCOeFA+8c67CkMODm/aIz4ejcEhhiPnHzz3wcptiJJWMCUqHm+Y4xQp
viIJdL5uhmFbskOMhHUorsrYhgS3kNttkU6mDqbDQOlO0PpcU+/hSKmj8k+v
FHi9QrU9QIJ+qhp/l43NUqwkWRnzNzM3nb0Bxt3oCCEFqjvWHxic1ptTtu+6
gd89WJm/yWpJYJ454D9ekvA8Mo+3MRDmBs8XETsIMqJTV1wqIdTON6AU7zOE
tpDRmNHXeD+AImXjgIpJvcNXxg+Hl+TUpKI97pNx+KMpTZ9wTDmVR7I8MT5R
TQFaudpLOxodAE+ifcfz23ZJt/XNRs/g8oWOMLAuQ457uGNvhR1EBb/fM0Pb
UedXowa4u9MCeLaWH0uXCF3jlqHUvyHIoFEwtzJIqGv72A4VaDDAAJXFBmi0
0GZpRifd126esQ3DzQOVNIsTw4LUgNZoH+4jcQ3h+3c0io+4o8tkXU5EdGSD
1BBTi5xX5aRDhE/zGxmq7PAfvA8DLHOCXyXEZUVfwtw86SV9kTbQx8z8yGmS
DLmi0+RMeRyB+twNUCUIHWcJWNWY++IjKWUUtbf5jMhx816v0AhM8V/eBJLi
Y/NN4avZCE5ljdToNXffjDGAzWgrNrUR/lp9vjXx/8/0BYLkGPyzE6zDGLBz
iO+MjmoYDtY0ESTYYBEFfB9lepXoIX58eAdPOd23aZEwgFB5TzdsaeVhWGiW
qgjouIdatQOkilNxYjCu3XxdYHFLgEnzo+wrU4pcfs37BNcp9MeNgc/dhR+v
N4kBFlsnDZMZDtLUOLHsHLogViKu7X0qyslFvKEpk7cQIjkJJqwYPqM+RM2H
7ZzDg7toKBzAYkFFezbwkUCw1Gw88/gKuouQE9dQbkllfPudbJ2egfw9j7h9
6tnbFi8Gq98Kp6DrMFZR8QrrQHTUYNf5PduqFfXuxPZLuFt8hlHK24pqOzjd
pdGXzHwVCPbWlVlMI0ERfU6eXoO0Gc/58iHBQpcxTmnx0scTaunwGo/J8chP
WqWFdO/K2yxCS/NJIws+11kecBIvG6V1XzlJp5dv67VEGYQWavaEnJ7uPw67
gXqC6fSpvb3Atm9/D+zarYdBGFTNzJ1P61Y5oFYYsMLb+MSF8OVNcLQxBEk6
MyF7yyJZhtXJrDkRrVakc3hvKT3ezVBn3r9GwEpfKkHXeAMx+B+OgQEuA3ti
SEDd93z6Ss2YcgovCvjwqEmC7sjwRJC38pgariIOwT6i/Kg7ImFUIc8Lwkt5
m0OhZjCtqMgMV9uiY3pKxb2JtOfCUbbIB6sSMlxl09LOzT/4EgEInY/+/9Kv
L49dYXGZQL7r+v82cbmaf3yMMLS4ANzxA8MlGZXesXSjbAaj+sTGeqTtUbDX
bWCVjnjwMoN8E91owY1Xgkh/oKv7bcMfrDTfxaXl6raY4riPW9x4jhhlNBMV
0dkUTHyLRiPqdUCgPPCmUVROLKCcxMGsmhVeZa0x1TiVN2GjjcZ437UFG6Bt
0wAqkK8qZg6ktY3dUHLc3ru0vfRwbORduLfMNx/sik4sBioreOJr2/oz1Gn5
b15BWsnc7mdWGaxxiVqnNnr3PqSYNNQRMLFVZjIYMr99v3ZXH2IdxDG0HWuy
AtsttxhzTzvEc5Fc6lUY6IKQYhvCD1mXslTslr6iiyRD+8xFFRV51Q3Vimsv
0NZE9iHkayQQUtdyRx2sOumhkLD/gbxkuf+n+JslG/5oa//jFrsIZl0ABDKN
/rNFlajuvv1wO3bxZvVt5kofU5+l0khVmraYgBerdIDOFf8b6ICg2R2OxE4A
0fSPgiOLxV54x8cT3VzbCA9e+XuXup3dcRlVSB6grY4B7LxHw9PRsdYee7Xu
KgeTYvf/Tgo2HFqWIqMhHgXgQ6mE7ggSBlZbq9Ce8jPsHJBFnqwA6aKTAN6Y
vDghma4EHbvj58PA3hHPkM+sY/iYMdHXwB3Y9uRwvTPF9MFkVHZIPugfhL9T
nT7Dt29QEa66m2ls/vSRbY9Ve4A5I9Rn4vateKqwYS4oEuev1krWwTAKEpIq
nKZdgu/GrevTGuVwMp6nXlESzFDk0wG9eG1kqeEYPx4rGV7Py/8uQJBkXSvS
uuABdCf7YsHb/20P3t3riqSgILtyZAetEkmICsErLxLY9tAkmXkk++04EbYl
Ioz0UuoU+dZdU1fowZCNIrcfV7dIMXnz66nuQwuL8rUquL2bQ30315pvDPPq
zIM04GqPFsZMQuVPnJWOhM52g/8Z+kcB8T0XJMm4NCpztUlmL8Bx+0Fg5ULL
QScz//9eBoDPXPG4GF93xYYxE/z9fhFVce+Eytk/8UxS3uj6Crj9Ad7UGgfh
U6xyELn4ZcGcTmoMnJ5Pe1Lo0GLrARN32YXD+8Vr1bvsTL9N29Byc3PNFSq3
N61OrH59PIhuzVZQOSzPFN4/M8mNc3lIlDP4gvYej7I0v7koCmT+UpPCA50L
Wm40gLm+6qT+hpkeFYFEjgU5BFTGg/zurrpdMOXaH8wEdIvZzGbzjfN767JH
UvMgfJFXKvkf1rmiXt4uQh8OL/H0EFIC/j5rJU0yW7qBfAxiY+WWEb4gjX89
sFNe3imNi6nT4RdK3zW1uqR6lZOO6bnoU7KAhcRaqGnR3+FHvdhDbIItV0Kx
KgvxFFl2pPEqXqWSxb2LwwlQ/Sq4/vEstA3ZwCzaiU3qiescucgj9fqHaadH
oSr/Ryrj+BqMSKPg0mKcFJg9Fn4xqu2Xm48bu4YXovIxlQBRZthxvwFElnqL
RFvLHvsnafa9zHA8U7SDTfdlTV/aUGR27Y9kHo94aP381WNoS2XX5WHxtGte
vuIifDdkM+YRofHpwlrVkSOyBASlcOGwkKwLEG8yaRcgi5Y1h0yWHKcLJNcG
o6i4khlcsjjL8/H7+Z3VifIwopiLBBgdCxx+RJNxu4EuPQ/HcwTN6su7xFH0
i0X1YBMb2ATjnUZUZK1G/4Xx1HT31DJClNhraDE491pWPEMyWti6hPbLT6aD
PjhyeqOGVjV5BVbBo1730yIKcYXYToRysasmI+OTiJqHZcgdVzVIv+cYxOWP
d1XBma9t7qoSEcmHn0egqZcNz3cdq0jVGTBRGK+XQX7+HM32gEToQmD/wd1X
8arxCxSUwxpNigBdkmjiEoDxT5VltW2o5YDyYR1R2x2KwIoUv9S4eTqpNOyw
LxN+90EK2+ks8sUEilyF63Bc9Z6HcYDZ+H4q0yuOlVXDJXFRXSS47CJiQpZq
+cYb4s7xmO3SJDKvtFwyiVGuK6Ay/wZvtVrefgEOpv5hVHj8QazK1VpO0V6J
LyhKiTcP/r/+Ppd0vQa8D2Q8Lr45wlmEhnSuQCyzhDbl3Lke1c6D7g7G3Qdj
wE+WibQ3/2SZIrXNIhhMYAhIAboapWxD5QpBJahUW6yxaxMU7+gd69PlZmQ6
ogG+4fFkC6J7ChBMt61hYZxIvk//OMd839AnWKGLdabu+ENAYiKa9ZHTj/6k
nSSZleWXJY+WJvKO6KnQHHlmnVzQq9M80SPWEKpcVU/xDO/Xf+m2PrNfEBot
dIxNkuKm4+xR84ySqHmprnwidB9r171/HYChsFsnJ+Bc9pdrg13O6qMS56lr
YlkCqiUCxanu4maLVj3BLe9fvGogXqs9vDt2YBPLzsd4ILQEbioavbm/0xYX
Fw/Njg8USBgFVGezMfg0SiCkhvTsnHmSANkSEQZfisPwseC70hF+P61Vh98E
hIcvYYPLtLCZMctmehjqoaGcLdQD+0c7jV0fDHAeCsvNkAe7R/mQYYnEzZFL
f4hQYhnFqLSNV6Qw2RUT/jBdhk5GkDmGX2sXzHk8ptFmPI5YWnfNa6JHG1X5
nJK8W8cz1JNjh6TZuEbKJdFRzgZVE5Ju3bhL7voTiRMfnBcs5lDIwUkGHg1Z
il+LZjQEq5qZWbIb+AzPv+hXm0Xwf8yvHY2IKmdYdvXYdc4QNtGmjdv3si2T
TQ+0m3FT7UJui1GdZR4NcPKz+NM0ZgYl9/vQflJAiJUkkJRL8JyaH4TQmu1S
U+racnZn/Bmo5+4l7ho4ZydaIlEDYGJ9SjCMODOrvXDq4J3TjE5RO2OXtfFW
5PqRCIJFLJA6wv/Bp/5+3nAWG/++mKss3KYLdpE08D6GcZczakYqW2mad+j9
epp/aUaGUjlyi+k6zj7rXpaqISlEn/aCbNB25nrvk4Gkwk1Vo/A3zFU7RNpm
MOyHpeeugKuUcUvk8tlZmG+rb57CvYINe0iD6he5KfJP8ixigqs1p3Z2Mr0z
dnYJ7bWe+dAuxsE0CxMF5wVL2natqDI7ZYtBokeUoKqi9MnqZeqzANEEW12r
8mTF2eeD1ScvoFPX6O4ZJCeTxyhhEX4yWTzGsOL93rHb8C6Mv4bGygPlQhpH
ykdscf/c4t++hKXLT+fL0PbAAnmYiXxy2gTVmdx/tu8pw3AC6UtM7DlTKSMk
ZiSBw2UqdU9YFL9kHW7+DJzatUbLklPE2VZ5+zZ+/mgyXE1u1JiE9q3T3BC1
pwW9Y1o12JlNHx3yzjMGNyepHqgizHSAbEYiym7voCmD7grOJd0OJrt55PbB
vlAJITtPF9mISQUVOmf9r98snS/jCnOCNPqX5FQbQCBxGucCWMXXDDr6IKbV
+MTgggluLhP67LDPoFIJ/GeevXKUt3R8N64K4qZzpDgaaPNjrA1VPTtxDrk1
t6P61f0S6WxLKNPn+TRHALxjRNcBvRHTSJCbfvOWfMGK33idCVURruGGAJv9
84xYEfO7j3RUYAoCc7JctNST7QODoImFQIzGcuDtI526UDG+vYcXYHrvBe+2
sprZwLW1iwrvCUdjwZiL5cLEIx0tMr6YE5Vku8Srpx2ashyiegkX/6eZ7fye
mIu+j275DkGYCJ5aodYOFEcJrSq0L/4C3ZAYyOFLu6f5MexBD6g1KNGcQbjI
Ao/2ZkJvNglj39LdwT4W7lKKSqxa1VnT8sdzY+QH9koWrNkC2Fn3Knd9pdIu
tLgm4T8DYTVp6OQz/8YUipH9Rx3M2A2+asP11IYmwjdjZQnAceDDKY7HWN0l
6Trqx7FgTxJjKFo7Be3+94nxixf9D8eMJ8vrITRvXRFKyJVSzHxWbWVaINDQ
BzT50mNQDrZoix1P+s9sCdDU9UdJ9UhJc7VUPfK5Xowsiw13y0X006vmNXiZ
1REbO0/xbQNfIha1Ek1DJ90qp/EDFzjDlxnedcqAThBbccr7NomRZQ/mwFI5
rOedsjzDwOH2uAL1B+BHyKDlly5pHElPJOrKmr50sK62heRmJS0fAdux0gqx
6uHuLdJtdIfOzspTSgjctU7idfgJrLFvu8se2flBnKi+N+Unc8AYW6Qp7uNo
iyfk8TW0D9TEXeKnZgHgRhJ6oBxn1uWKt3q/SQUVWXeAXX/IT7RZcNmDjX18
YDp8scVN9PXqVqdKufs4CkOVgu1TBI246PthYkWYmlqV9qj1IOOmve67oJo8
9+KEzsVt1CuxfPA6zNL9A9MoLgo8we3i+zrlzfNdV5ZUjiFL5kQ9E3hjx0e7
o4aGZT55rI0onIITEheskhyppEAOz5oFCAxicmrY5+ggtNmAhYa1siuEaunv
plohvLPQh7y30EfUTminlIPo3ZpMn658gI9Ap6cO9zNp8JKQeRXFooHq6bRk
dpIj+6U7R1ujCaVcjlQd8lvI50At5sEt5efVPoyKRYq0/xc/bUChH8QLvRWd
S4xMYMvR+FNbMLh7bDslpHjpBj4IyXTHY9swrai4/7goKpDLJby9l10vsoY4
Q+L2YFzFg0eIOREFbzOPv7SVveP/kSQuVVaKKiZpnsYOlzoByqtRdX9yV7Iv
cIzLVvQaBK9K2xAT+3u0zaBQZr68vp8eYzCGLXk/eOVVn0clVQsAYnrQbydb
3c+jbIn5HH3ewiy6Zk8WRbHY5iV5CxBTDRCM3KwRdrdX8OATrirvd63kE0Oi
jtgN7A6M9kTEv6doxHOakCKiCJ0tIFmabmdtTjcxrVSlNiyWOM0dSVSOI2xV
rc4I9pvQkyyHPCri1+ABdMNKP6OlxyfbU5rr/ScZKEROhxRj++NrEjdFOe4B
m72rAxSnHgJ8k5GuwGcb8aElIWiT4ZJ4g0oGWAuhXNGw7pH0ZiWIeDTNZ8VP
qI7okn4c4FJFQnJLuFzu5I5ezZ+qvsG4rR4pyzb1B7tq99VuXzaMuFBq9U1Y
fH2qtlAwy2vLYAE1FcgYoEFidOI7X4ANl1orjXALyL26TUi8dynxrMThhIBP
Iupn28Fq05uOl08ankVAozi/1KS8sa11dUC50QLcchliK9knkVgKoJBP/92F
I1KOJJV3AXKe/l7/QpNnwaQKmD6FV9u0H39o4zDRWH84aGCDyiQLqtnRBDLm
WkOrtg0Ar3b4EQp8lmwepT7xb12JERsOEoXd65OPXO1WPzzZqGYbBZdocCJj
h9UoJkF/lIbwU6fAJ57mXSQCBoa/irO5DNNIS1l1ZOzUMXrRNWjtzxmZGJDH
37Jr9QIkylxzLaXtQCU+eATZi63nLhkNl0tNtRwsHJsJKvbyPsKVZcyEeetf
76Z23L/8UbmSKJWzwqiSq3xCaBm1p+opI3i78S/wRxBA0+KkLqlKLKh7NbAr
2mgBKsbCrD6SodRRoFBkhZwlToALS4pFcMzxtRn7NvuTqERDgdbiiRpD99M0
zVSh237UF3t7KoF3Ehfbtt1lSiaON1o2BFK/RrAn25g06Gky6JOgjFnIPUU7
zVA9c1BgO0wToIjp+Tx0y/3oMKb19A+nGKDRjYewen/gk8xgZWc4ekmagUxM
XY+KP6YpoVlVvGijPyQBmtF5wRdK9uRsxpwbh1u5b7F1os6LqqH09+10Nt7H
59xN1gSkG068wmo/8AuF8GbBhjZfMSOM/Sa5b1rDGkx75cD6HcqE4klt4J1C
9tnCFWgdVfRTa6h71Zv2eRlRmBvKMZk4NLkrZ4riHsetuTiP7xK0djbsS1vG
nzGW909uXJkA5swhdWc8S+sFEkZnCIZXsi/W1MA8QefWrEpYFj99vUEL6ggx
H6Cd/7tlwuWlFggjKKnh4qHvK6OKobR4ofCDggk6ciftlZvztImrhbuQs9VX
MwQ+h+Vt8MT0Xr+NNvpVsHWqwnU8UHdX7LQCDykZvH4EetrFIVXkQbmjN8/u
bpV3FBHJpaD8CFF2iG+ngwRKATGQV5dmMySXtNXXKeqxNTfDMtwRKoeikdXk
42sUJtG14YwtxQOl33t0Ktx18Hhn3CkYW3oVfHo2XlZggZ2KLsXk0nfwNkOT
7Bu8bKX3XGpIOTB8J2kl2JEvZpyIYVKxtLm75eU8ME6yCUr9k6onyql/eNQQ
IN0dZnuK0g1oUrnL33YfFbFpLPUCCbcFZwnLvDO4D90EKluLbl1AENoh6uBc
SmOA4heaiKz8z+MWdqiDHa1DdLYTsLZNs3JIJi/nIN9oN8UpkLKc47wCGybH
kqgCY7IlkVkGNgoudx7+FqchvfLmcRYloKuzqSQlJBsbRc7yDjZL6ZY4Agns
wsNdhKage6MReuNW4pOZ2UNOYOQ3+usVWAdv2JS1dFUztk5sY26vI6xAcyyJ
Ycwu3bWk9Yr5eac79MjLySpJ+IYdc2hZrRWQDT2NadiyxIeRQCzOBCILkoN6
Gpd4XdZL7boyXbvTEFL7K//zuABZoCbXlG0xR1Am9Bn2B3bugMDZs0pKRyGr
9mrAZBWj0BIfexr3yqKRnFMBhzocEf7za90EQKkFMM6vmPoucH1G0geJ++Tj
Q80PZB06acL8Jj1LakoCmhrczd+saqN2b25qNFuGyKy3xbpKkN/tkTlULHGe
Ij/gwE04v1bXqfeEcYT153KY/K99m5IiYMOptbvyco3xV8eHZzudJzfWrpc7
XFgrabMWvigV81LhJOwHVhE7r+r/x2qa9HCU83f3zYQ/ni4DRTUqrhNkMMKv
0tQMBMNMdA5YnyV28gto21JWL/yD/NVpxfFSmY2jbklOiDQRea/koMRIdW+k
zfl5LcCmXOrdeUmdshChBZ4AqpELOPPvjssYxvx8E/AJOyD/WNQP+gSyi4xH
Jr8yrX58L2ea7WaU4SFk/6k45FvHZrs++xOkHhc/M2kMr7aAnaVLe2mUjK9G
wmfRy02kve2dFGNSviRqZqXtoOyAbMRbybeB+q4vBgbAy1BhJC4pO3uG8lKR
f4OJ9da5dll+CxvsgNtXyPCF5DWGZDA1Psx9JegndbqxiASgHt/lrP8AxHVS
McINj381Z1UCRdO35FF7kXAfCcx/GIsJXsRKm/MB7ZD1+3vtmAWZzU0WB84Y
vTbZsd61AKp66ed8DuGbUuVIDun01GorlM4vlqGJvrfbum2pb/DRCGGNl3bo
ZrAj6Q2zR8/img+/EM9Kc+8892RHSJtqWh3abyF+JvPFV4kdfVX1K0I3pC4+
tfsQHj1jfgXJ3Dzdx/PCv1vDKMzm35I5hGaWZn0cZRiJn+T0MeAdKiu5N/d3
bCvIZiWK4zLbezSQFWjmU/N5Zn9WulzMC95b9v6z44YoeakX1wNGLJ+AynJj
pQ8dHW7ZVm1q99U2TOxUpjRDLIVw2a9ebFRBE9nttJNYaPXTsn59/JpJ+gwR
/cgNrXtyS8uzNBABSF50+wT7qxIAOtH8xZ1Q/tA3gYhEs7Wf6L3TaXWHb1rc
ogQ9l40w6Ve6L+l2VpM3ML8zuc6KhGguk5OCQoS1sV51iLvCmaACCzSRmDFv
OolGI0LyV0mwJhhTJvLVC5jW8Yq7WqZ+bNxFmM6A8phohnP5mQRJnGZcKF4G
ShXgmVH8vkMspUZC5scToM8Z3+1TOy+ulIbgtWNQtkB/k+P2PWjo6KFMeHXD
FdRQoGUytW1SHOj7GstjM4aJVtKYeNnJjVupb7HVXig/MWu+IAPhQxA45HCl
MxE/PIfMcI1GyiFwwEBoPHLB8K4flKcTopRvddNqfMPixXm0uTYbWaWS7w0n
Nymbp+0skK5KUU8VevW+yNdcasuOasi1raOPROPGTF6/FENG4atIGfr1k4sY
VN76p2Vkw/RfysIQ8m+th/RedHVbrmEFWfQaIKtu4hqR1p9ad2GQDg/KVfgz
+6LRpb4cBSO+zYiYVkgL+Ar5JIenyTGqWC3nvyfPIicIw6qIjfE42T0LdA5O
VvWGd7/C8o4tYKmB46FoMIsgaZyHfLtvmU/Y6jrJ8UIjlOHUOL3MDUmJZIne
dXll7hvDd07fJqKn7szdDk6YrKKO8eQFRO/kKGQWuXOnP4Jb3QJT/Wx72qgq
363h+mThYStu5LQRHuS5bhqYW3SGcPqhBkYPf2Evw5EcqPjv3KsuX1BCGCmW
AqjfXuJWXfa+Dg+CwdXhpOEwS/yKCw9zcXeR/eVRU6PI81fsMFG1TSo1pIzO
R+aUGWrq8esnVQ/c8N9EJr0ERJDWLx9uVRHGQnmI2I6FlBeJJY5Pj0CKXEBR
WBYv8UWYlXDkdbu4vTf7h4MAWA9Cgl1dki8dARE7nrngSEhrtMq8eLENEpqv
9SLe9/7BTm6XDq5ZwxHNllt9Sm7b7cHQmDUmZ7hJT7L9yyqGM+TL6K92P+86
ZdR/YWTU88fft6ufMpqExUf3KTNUuKwRpefH+csxMZqdWpCb/hTiBHrzI+Zw
NRhIYphbdND/l0pqKIwZhbfTFhSk7nWHnXLKHsrYtuIWcCIiAs5js6o82Ykx
R4Kug4MKnBnaSCVKVZJeebqtDUD/3Shfpy2htcrg/xVGg1vzc/FNjfZ1m9bD
u2haRTWtf6UZuMjItaImKTLyE9oJ3h8Ooa3C2QmuYaHAxAnjgpFG7DVQuJSv
btmfaNt07iEzuPPEkvS843dTeXOmpLgGCSo0GToJY5lLc4Q0QfIIC/QxTg/H
rfOIdUFFsLs7d/5WSpB3tPXvlDJpCbO6cbJEcxqUg81EbNMPyQeEsl7ky6Go
vG6v/f6abNhLT35R0fxnZ9myTiQ2ljHy/lJ5Kob/wn+RsaVuBIYhPB2qAYYp
VK+e8hqS4JJPf75mjP9LHiXBz5HVrev7PrTxz/U0EvfaUkfRw7YMjnKu9eN5
8erpbks3gGg/PqXflw8DTnufcTHZ1JmIKLolTtIIddmXB6oOojXCKNUuBBNQ
nofTBNnkcKNC00tiuo6KGd2BYPy6LyLzwgzMrZV2YPoxnjBHkdST/3mbGX13
FkeamyR/AHnd5VKejEg9q6NT4L/eNE8HoXJtcjhKQp8EjJjdV5VbAzGgNmhB
/NAvFSZ3YYoJmHmj1kWUIWUjqmX7MHRqYIGLYcMSORJFe8gZUn23dN8zdy0+
g34GkV7LNIqIATiZvDfscyBfeeuTk0jYZQZBKgdKtxf651EM0IS+zN1CN03Q
qKLZveEEOTPaOwQrWFtEmCI4NgKcojCUmFwUFOoXuak6u4X0ZhR2ZgedYrI8
YWXIbokKg+nFBjCXcCGrhqdzzV/KrUlcNuftOMuPq7BqACg7kZXvJwiRGf8w
kHQ9ghzEFocKn9LfA9Zn2OmW6Lx9IEdx20+UW5Dq1YwAFXTS+DAsM04sBoQ9
Qynm13Xxl53CcPhuUNL9mQP0om4eW7cVdh6GurUKky4Iz0yGi/H56uLqIIAG
Yb28y5/vUQYc4qQxnnk2X8OIQiTj24C8eryRJZXLbIKW1MDLqzi+HlA/nIwE
zwu9H6t0gd9TL95Kfo1acUiGQoPoGSzfsWr1lNvu8FY4R5CDFr3AsRpIR5mp
H6NAz4Ig2lEo6N2RwGrNB2W+biE3BlU7xx8TG+J8ISEQsoZ2eF660TF2NKQm
2yrNs6Uyk+UgVANuFuYUP3kxHnpKJDi7HIHeis2obQlRTcVRdsNxclWEIKhL
CwrOFv30Q69mn5dikVuFGKYRm0M1nVUoAdJfNZc/A8eRLmYX5Ogy0+iPX1KR
CMOZziBjDguhd6X9nNmVtNu9zhvNRYQwzxqoO23XTqBc/dT1Z7S2yK/kYH6m
lC88aND7hTAql0+WmnF4LxFA/44uKzi5o+xkwioXkNFUpS8+1JkMK84MDuPX
NfyfMVYSK1GgfOCRH+BjmDcWc3wm6+gfK0uo5kpQT90AA9cOLEu2OrZyRylk
W7kL/h7R+7XAkt6LIki0INfSjQCYfqCKXMkFvRottkI7nWhR6/W2yik72bIh
kskA7fwIcvfX7T+kdvCDzFavBdwOYLVh4EruS6p5s+IVZnXUp66np/sORdiF
KhFi8Z41lpMZ3TQ3CWtAoROncaeA7Nd0p+COZhWE/AkPduD7NPUQb5FpEj7Q
wg0e9PTzgI8y9Vx+MDlL7RRd/jylHUDFp5IcrksaCYnfGKn9uAb1JtFv+J8A
R+SxU89xInblgRffm0e/y1rsQqILJbialDVvcs3OCkJ+q39BuBkHMhJNVPLo
SfcYfRLNE8qqEsk4N6Pi30h6K4yhGff6lchF8OaAzq8vby7Gi0zP5NnB0Ald
g3dAX6n/H8vMdqVYX2NkSOENWeLVVU/uwf5rrIg8btY2LtNOsvj8qvbQo5SY
+yy6RfqTd4MpgRzazGjcvpfEIcuSXPZNXodVVTEClQAO3/XWCj9BPIg8/QOw
68QN/NNC2sJaAJMrMg0x2rqL6z/as0tRtZJ5n3VTOmIn/gELXmbka5Ya21xS
kUK0rNrdUQjRAlWFn43Hk+ifrsdoF1T17GXgUyWBg0OcOZmuKZvhCCW3Zsge
l2+nMIrXMZ6Ns3YR7WqzKymZDzqATflqzQBcvoH+k4EAdgRh/DB85upfSff7
Igh/EzRWO64tMzOFtZhdREzmbchYMXSTJPhqZaZ3w0rGDDLSWngYFpGbTD79
7qWV2d0ztr/RX/xYvt216agucG+XjBUi99RvHBQRI/YjsChTsH6GkPGW8ZhN
c963B2aNS6akhT/5BwRTK8maVVuxSDI48bbPCehDGN9de3Hg3PUp2sERWe9X
5Wv88F5wQkECLa/cfV1dgxlzqr/7M9TEuqR8YGNCJG0D6YgSx+x7BSvi0DR1
wpGobQsiiChxhBtrTTVxNG87YHTjdTpxsRBVan7glrt1L+RCUxcVLftIybGN
tYmTTLpo9Od5NZHM9K5qME4wedH8Gci3//d9zhEuluiUgFIRNVrwHV+7li8M
jJp9RmxhgyqY6FY8G0G6zcZl4pqQk4rm7WtSg+NCkq4MU6asAjMg/w4pdzSO
cHSHtMUk+Sadoad0wKP63Nv3No37WTStQ86BTYISjis6datV4Xvix1gDSTNi
0baxGnTg3hWbGvup7hQ2WVFvvvbjZzA26odLHBXUfNivO4CDpD4YwmUP0ueS
0HNDTAh1F6D9c0/v5b7LiacPK5At3/vHIO4rldCMywOre73Htqh7tQrD+mMi
mveyVFb0eSIFd+se5CYiYg6SzMuFaS07p6Fo8XCONzy3eoK6myS9D3fXNDHi
TvaRcpxJRv5cpemp3ekfYq7VtOsfagN/B+WQO09aqlNTMgOkxoczsQa0Ce6x
rAvWnqELz2nSQgu29e6UbmlZecRHPHl/+dhSmvzUsGQy+YUIrjyN9LVG0fVF
Y0oEmb+DTKLrrKUPF8JvmEiVoQBv0WQHB1WwavZRu6jyoCtNW51MdU5DsGmD
kcBPOx4e52tt+k/aMZXt2p6bIA+oXT8cjy6CGd4zvx0IYiodEmgs4yVBX7TY
zeHNf8q9+broVYexgPqav5S3iq+xcp5d7NwOrVVmzelwMntzH1XRQoZ11mwr
fecgZHYyDf6+7vf5TF3q7wCEMz2ZTbM9iFGNugECEQ9DOgihj/gVlavyXbVV
Qn9alvFWTt1FCFWbfuS0FQdWUMntw0NX3dSHLMgv0wE246+RFFTP+MXY7vgO
IIO0I8A5VEfDFmnWKmzc7Cm+FTr4ekRMom8kXOEntWGrGQBZkY0hL/NjRwAP
wO4BTYNoHCC6x2Mev+j7v011odKyccbqR08gz0BrTRMhpblDvj8HaIOOosM+
40xFyDW0ee+RSa1YkWpK90gp04zRwg0pW2MyYf4sO1UF1pD6/EYnM6c589fn
o5lJSHjElTTLjSjas6eZf9mURKEveMVB+U78MWm9KxpVoZagIFxMjsXvWAI/
Qsgn1LLAP8Bq6qeE86hcQUqu1aSBgzbuijapyBtnJSXHwjSP4txfDvthex8/
H8z90zHGMYSdBpKt6mf8qzXlALe8i6j/kXlSxTIahPDtTwrCy91m83ERvYhb
lFORXmAXIbZVcTMeey68X6SJzz6spNESdwufJCZsAUfu9b2KFyYfoxHjVpjo
pdVla9F0a2AfXty1aA+43M5TerfAfCJl7Wh4TcukymyFDEhLG7eMg4GDz8xQ
29F+iyNiiIXwLNnNP7teYxeeb9+BylI56WGuWiJcLcZIoBaH99r8K5WBDw/j
sujZ0f0kywAz9+Zy+JnJp1z4EWol6JguSjMKLgyax+eTyldBmLR+5kkAl26e
14z09PrKCB0/bh4gjrnlZsYkSYMS1EvtEdX40D5af4mi5me94OkBBxBakRDE
IInKuwVEyzUPGuUonk26WQETeCc0TecPSkLSaHoEkz0YevTu8qQGVRAWAqAR
lSpP2FhrBJEpckaoCqGfurxKZYkrSn3dL6KyEbobdO8+LwczMJwGx90D5GQS
PSI4pH7CkXqG32elWjl4A02FOIcMp20h7pAmMKon/SKOqlRzfXxHSYefF/pJ
pBdJvZg9YhOt3CjhoVxPjZRy04f0jJ8ugfBHFg/Wlxg/fqjFAWR9GUSTXrCl
OC8A0uxbUu+Ro6KqR4yPqpOyE5Zy17/aCsqE6tKXBNY45zdgK+otk7MUhhtu
BPDAbUS62LU1HidffIn/5Jz5/FgdcgFwxnNcelt5O/nHQeRxZF1bxdRpY4DE
QIBi1Ih2kxfL65Ra4KZAKDdrvVkBuRvUvYmzj7L5S9Hy2LxXLisseQetue2p
UEwT9geSIEI9v6qAVJOBM18tVeset/5IPMgb2PwLKgf9Iz1cLACIo/fACYoy
o2Cjx5g/PH/GB3bDLDZ0zn5aa6Mrw9LSoVsby9s7Al/CbvpFmXt5Qkl9hdLf
pyP/GUsZetkrJmhbWy5ipPscN0o7AkiBBzOCyldSP854dYCd5oQvJGNeU4t4
HP8GGXdVARYSNusspNaUcTTm8TCnktzlU41GLMfR7ypx5MaBF8E4K3CRW/+a
kCC0WrCiQ+FUzs5ieEyD9/jHs8siSlH0cTuZozc8CZr5mOhESryMF47H+Y1Y
sH/+BAl3t+gl4t8Wjtx6aoJVuLWvQYyn6WQZuxDWH/2bKkLz+ki+OPt48vh1
gFCzatRE1aWCGtKmHyJCDqvAMqKYcibL3N5c1zkOxVDrMxQ7+XbcYSUwH8ZD
0NrExaM+lcQtU14XNWsgeZP+PdNFlh7vGnNZ/Bjd9MpOVUhj66C8U6CpY7s9
7YmrbCOZ8W5rL4rkhaxwCzTqz7/aJ3rKLnTIqCfZLgHbmW8+WMbPnqAW+qYd
PXTLXerlv/TkjKeD4YEziFHZh4bKnrr3R0CXii3/eMRMNuKWtj94i9t95//3
n1NWaZba8iCGS4noA0OdU8bjCu2OlEcotd9F9GCsmPV/0+qCN/PfUviplRFX
uUtGKLQB5yV+zaykuRFJkloBS5vhDIez5L/9y7BS32Q3eoAWsvevS83Ide8U
nnGT0K72m2nPUz/r++jDs9oM5cDSA1zBZNmalrxv6Xo/jhSxLfh58TaYz7dC
IH5yc3CncG+7DyWHDlBGxOuxtOp+2GFHlE4EhY81Hiae/Gw9tUu//dD120t0
okkOAAv7XLaaifW9UqKxZ3VIAp2jb2EU/eFWWk1RJyxaE0tu98q767OWCGVr
PvtBw6b3hIrZmCb7kOiDuWlZOFB6pbAfEblbMZdBGdv1iA1TLoM5BFz/Y9v0
IjcDyRSh4uCfKOA0gHUsVNsLkfRsiWgH4CPyj0loPsuxmj+YCTudznL0PQDI
0rJ7qI5XZXq3zYRdQHZSjqjM2iXnMVP4iR9ZfRwaY48wnhJEdrZ6GmTmvNeH
zpHjsiu8MUf4QoNqEDn4LR/h3ybeYqUtO3b+kG8yFwCi1ffax13w2ykt4l1A
XJfns67n/HxZxMGojurHFdSOnP/AyaizT8ytRebmGif8MDYTVESJoGpAXuVA
LPG+0OZTWCLG6SKAcChabrI26k2weeviIJ1vq11oP9CEnmuO3Psh3P0CZrey
sgvL8KeB5ZCy5gwiVOPxVExTtjhzThlZpOAgEq20ZJeJOc2kCbnjLJSzbYuu
+oUlDR3hmfgtc7z76ruyhK5j+S6E8Y3OlYkGrWgOBCh51+nM9S59i7rEyteH
RyxjASB6mnX2JpfHPLQT7uojNYtbibzn3jqHZgsqz4A0QyjWXsRuPGiW90lW
BHIDiDVljsiqez+PMLimEogP1UjjU37018mVA+QzS68xkmpn5W3splm+gfZx
SjGbP0IHKoqrtlAiXnA5RIEoVmfdZdGViEbwjOY6MGbI7cPXMJ506EjwsZuG
CZyH6CkxbMz9DkRxd+2eLK1ZY7zSwx+NcOGfVL7cjwZAXhAWb3js+oGFlcOM
w4IFSBryJ4riL748T1/BeluMsZErA8xs7PM3GzJAJItFnFJdCHlaxkNogyP7
JWIqKHsY4KTHRqlLECdW9zhA6/XWpTp8VXXcio0qvnXeFoe8Qzl/oBoPoLiJ
FFBR2xfrWa8cN1fdYMH1KtNIkQ0JH6jtRvrugJfvDyxFiGrAksVNu+/NYsQW
yUtciVkZxfsU6WQFcDJfM7A6SSx7U20o+TH5p5lxvRm1FIEvgnrKT7+9l0jt
DDqgARcSU2CqmEmHkuS6qHr64+u04IhPR4oXZyqNT2Ow2hAhXMj6oP/5G7+G
SvUDuqgfezRM2C7vcHIAsuTGpDif8/8F8eygX26rNIdIxCpoYbUNyoA2jb/7
LAl82YA3mLeBT68G5357YhY/MSx5zcmU7O80EszkhsbznoRrM4FvPB3BQD2x
sMdwonLt53FtBfmzw5Oq9lBla8nZMlLZw4IY9uO+BEImvsJRuVG3pmISPC15
bNSof8pKvLatvpc6r0AVGzkDG7qr4odxEU+F1sGMFZLOtibM5rYIAMrZAUIO
Sto9NU8gZIPS0qD+PWThp+6sfON0PK93w3Q8VEmrfoV070BVKmI7N5mtt2Sy
RA90rCBDjgP2xyNfGkeMHa90g++SwdKJf5aCuzcmjwftpQVWA0k0+nLToe+3
nYEm/3TwL8Y4Htfvok4WbebQJaW8O4hpxS5RV/qN3fp7xoFk8tSAA1LT8oIS
ePdM2w6kusdnAFAfvJYukVUE4k+mKTgD1nxNW5ZhS4OnXrYSCcPGFVzYbQrp
7ACAJilDgkL0fy+qcQDZLtELELIZNENdcjEIKss4Ax5+OW6YMBEn3lZqt3nc
7R2Dk8DW0LVbqs70/J3p/+12hMOjv/64DhzQrtYaix32QX882kZtXCMR4/b8
rLRQ6L0gqSm36O/tUGHqTW4XXr4PwUyznLpaD5f4f9cmjLHgKEF9U5HZ6CxZ
pHP7Y9nY3T2cKrs1cQOOxEyMp5hGygnCIBGYccmvN8kKR/Va2kzgq0+qBQ+g
ZD49DwOV82ox3PSE3+Rx06L7GXN/y0FM3T57wThE4DrYA9vRi+6JdlO4PW1g
YWi6JbgYiKGuCl62kNsQnau6GPS4xk9iHFIx+JP59QIr0LoU3s1w6DGrGvcj
JCtlQ9N+PyUlGLTGF2lcnbkjJqeuAcMV7J5r/wUyir/IaHptWLTv0ifKl9nj
XhZyqpW1Zfvbu+dworLQtmwxrfER7vJ4HZsl4dlTb35tEGwfQanDgZDXg71V
LGA7YCkobgYVynh0hh2Yhli68OhHGEtuHo8Wk1p6TajKHeRGCrzwP6BhFOnY
9G3z4wf7kFzMMVYqIKCwwFXNfoAlw5W5cdjICb81j4cXMPafP+jV+VHX+duD
IbeWanwIYs8x4VVsRx9huPtL75DHa42QOmjBXfkWJjRVZS2VmVNb9X1o2rgM
W7SmlDoMuCAKae9B1XhlH3dcFPa6CsG1TyMTZJQcC3jRdX+Pkyoc7j9QOYzz
VeMEb/bSzPJRMZyIzrMksiwV0+8m4V4IKui2CqlMdPKV7SMEngziVJSSNxAv
O5+zUaqDP+y3MyXgo0ZpB0mN9Y5xkx0m6wWf5TypaBJs8DSdkIm2FjX+iPW2
MbmedY6ywlZrvIySTDuZlRMrlvuirBn/9A8mLmxgwHq58NBDPu6KRn1Lt80W
xxXM/H0Zjy3NbyRqZymZq813AnwNc/l4H7wGxipXs2aaNXrpzEOhlYbMOtYs
5uAbYMtk+ouub7X+lN7pdH0NE++26HIUu3xQ94DS4mUyAcKLb+jTSMkJnMP7
havUJPbs+i1zV63/KpPgim3ACnAbv6zLOR7prP52hBsA3pmeTVc9RC7Mu3FF
0UsC8DGM1kBWE3QhDZwHJr795COq5dA5gkykdREvH/rvy5KU7EucW4G2FMqD
RCUn+VdHu2SmAGmG9dDFHsfn+Z3pIsLCXeCojqvuoZEfY490pw90slVvhNZR
Js9fSiavQ+DmQJyMBtbuJTzCOsz05jC00MDS2euPcLvjhXQOYKiuellbi7Pw
Lxxxjp7DrG8OvLVpOm+TDHhvIyRocg8uTAS7Tg+gSfU1FpTyB5wIIbRLx/yS
lCgTcv1F/HAxK9uuL/RV/4s7jWQpAZ3xlIGX2jTK7kFzLeSY2jx1xY10fpps
s/CC7oll3+rKviDmhxl/0zsLFXUMy/21tUCZwbuY7E5csJBrmSZ+2yW+LGqX
Gfyp7CajEy21L1oh8dOZI0hOayey9atecuSj2zvSFxaI2lMndx0QJdtMjSoL
BlkCkuj4gy6IDug0wrhgkHUjh7FH1duTZIMTHXZE6xyugfDr6/2H7x5NmPGl
UBa0RxMLNrDgvcYQXcdeYrkQ7ES+69/yeS4HjJN7Wsnyah5Cw1j9CjSlh5Yk
SX++G6QjFtJtIQb/b0qij9CdwGlb0A4kWGoPVf3VUOv/r9akHUEgJGaR3dDA
sas5oWNf8+kW7/+/Xugt593dLShrCzMs3A3MmNm8o4V1vcRY9JtAcRNC187U
IjgoLi143RY4umlIrUlOOFFiujGjSuBndydK4z93nvwo+VAFy65DNZCuzfs/
6msgKaYJG8jw3MVf+Bu81qJioBluZ6wbpI093BvB3pGgsQA5WacDgZD4mc51
7hi76ET9uI/3Po75IqEd1GSV9KMQkqnu+xbN3F2sQhAJ02GERUHPed0QQZ/D
jT1SIMMTFGv95g0H4Wt9KkZOzikzlctO5q12zHZ686RRuiAuIDuGgTD5Wv46
BEeyEDp/xC1OEi3551qk8G8MtJ7eYYqitI3+YG8XNVK+1eg1U3L+5DUa69TX
Ncv3cHBYcEYpJO5tjZiMK1Pgp60IpxaapQaOfuzxrK+A+l/Qn8Fly+C2nfMY
aERJgmE5jVzBpxY8Bdk7yHkZE+eoBSISuaHlt3s88fcwZg2qmODJSgh6GGVP
vY5QCwHc+evRgIDO22yECHzjirjMxqTix1J+WQsVzKQGquiIVU0yX3isNunV
qGf1TDf0b+GNQFYceJiXsPWXRtE+roXC4zmzKBrKXBbilafQghQSTsOEPW5L
7+0Bda9aDrZuwc4FXW1uIGuJbQyaRPhTCSlV2YH3qwJUl5LkhWhZjOHoasga
WqsqFIwrOGtpqP+D96aBwA/L4LJaj747CX9KmjJOBhdWLxNalG/EQzQ9GEtx
ypC4PENty3h2PaG72mMlFS3G5VV0QGsPA7Pga/rK846benspqKL7VI3TxR5r
khIWdYMVotZqZU/K9xcTHoWT08tqH3D2VvWNGpP0f86ev2ic0Ohwd19NEAze
afjDp8+BvWmIYsQmMP9ZI70hVZrzmJhpzTlluOT339+AhPqbYo7HOtu9r6A3
MZONhtoYeQ4kP0g3wXDdCyARGiLGyAvAiQOT696D3MaJQGaSwYhwkJrE0qHb
C61681wHIFil38GiBQVPI3c2HIKJFcpA4xq/56WhrLn8e4Ru4hPeu/t4Lh2R
qY91UTxu1FYHi7l+CylrxdSRGko1wHyVGR5IHcEtkg6JblSPopU2klX2wktK
Ot0l0Q05nQd7z0VQzAJho2ef1R9Ps62xrwT7Dq7ka0OqGzn5qZQYZEu5ND33
lNFrrkI/hpH50N10Rxyne5OqE1xeo2bQRt88r8sJrHWuuHaGsj5Ax3mvXl5A
ektPXmteWB/tyBUiwCUsogQ3546kceGONC7RrZT4giIFXcFXboGUuDsUFL/n
DSXKPvu20qrpxDGhSZ6bilwed7cwJXSU1V90O0SKKvegHAKW+HdwQsosgC64
MyHrjjqkzeThyF/nls0lAqvXvw/0CEEWUTnCctC+mc4D77nH5uXK7CUt2vIm
aK/1x8RHgTtMq/yo+z5c9asYT1gq4bp6q3aXaT1aK13SjlRVwGKPNcPP2MvH
mSFSGlahCdoe30s7zPfEYWgAEcRc4fOyTqgIo9qrL+2AP3FaOKqvKdN81fa1
UFJ2z6FUC6JCiHDQlQ3IOXnPXl2spKnMOCocdIKV1ZBTpdhPehXdDrbUFTam
YoXSuGo/oPckhE7SQVsuUeDnrP6iidQFQ8STQuJECA5g/tZ/sNuO+9r+rZMx
98+9BXrDNmyGs7GHvRYaNOBq8hYlrZkQE/5Jg+zTZzyrmHdA40STweMY0APA
6EE9n96xucRoEjAmh91/TGai2PpzHR2FF5reBgLIBP3k5Bqhr6qAmr/GdF8P
EDz3IKVkOM/jtKheG3z4ICcuyVr0jjhe5eTF+RdPQ2eB8+lREjyNYd5oo0u8
Gb9rQAZus8blQsDrtH/PuSVEmHOfZ2wMG4D0cNU8uX3PaTYXv+qE4L362tJ8
8pZCgfoEreapJBiD56fzmJquREZZd+K4uI0MqgV74mFw0YpSLIsMgW5b5omQ
HySbcvaJHRwFm1ZnkEM7J6X29xCw81dhSFSMMuqH22fBSjeyrPmnycKbHoas
3q0CuvN23OwvH5ffpVaPRVgX25aPV8ETNmbO6mTPSnwhuOgB95kzfOHLLPFx
sjzMCDWCpV6TZ1gPCNCQQ9HchI6OGW7YTZREwih34oZvJReykZOOSGsyf+t0
JRM2/ZwmPKEy692imdIIZMd3Mn3pw0AqtVRmxZIqSGWQPNVUYllKBxKBNEot
oSFW3qPNE5BX1vJ4+tB+8pAg3lNVebW3Cke4yCg5Ipo/Hwf79y4jJnUdNoCC
M0rM/wXPUGaGN1fJevwbbtXzVKz43Na//7KIm7SRPE4CSIH+T7qQ4Mtyhl7r
xEtg0zyliZcVrm8DuNUSetR0xlmYM3WZehYKWiLJnfUbwDwPJ+6gTI4IZ66F
Bn4TwVBqEp3x4xWmq+st6vVvkdxIR5MGJJsEkOfLeFEzpLAWegN6dr70HT23
FJx3Fl9JMl29Jt5/GxUVnS6eJy2faKgbLenmGkcCZ9gpVdcSAw8TH2WoIWSo
o4CwcajbNfKXavaOMOlH+318qoHGlaBJVqFHRSviaXiCnzZKO/0nbz8aOyno
8YYBd9xEYpyBJWGMH0YNFdwppeLLVfzywGlJEZGKrgupfn2sEULvofqfzZ3g
avB1xPhsNpcf+gBcJDkUz/JtDgOKfDDZp6FSQZUFLWlTfs8VhMI0eRZL9CPD
1u7eoUqC1SvyZ1m4S2JHy1hcSy3rM21lo88lmeqKPEHc7N4/hHvXWccLlOFZ
FWHlEU1rtvklNyjtpgr7IbB3uj8oD4ruLUxJjiSkD7JcXPU28tButx7FR9Mz
ySnC773eBzxYL1PDvTQKaFjteSdcENZ+/dTdIMSB+fSAYGhlz1T9K5wt/uSI
rvPou3nvz8OVKkpT9DbhOX11lHSX9+I0pwg4vkqDOL4TCd9gBk12Wqgv5Zdm
02qVBYw+q9vopSZNx4Mt2gPRwIlf1jeEn3PqE1vAtjTtIl5KiyXnc4LAFX3v
d0SbskxWtCBaVK5Nr4wWzZsdaO4ztVujG6tHc155DfZIS+4qRbrqeaGf6CJI
zNdyI+hzPwkVGxyTMH+0eMcGwZluh7TWCPsm9RIj06RG7gcNA/b9NjasQXp2
e7YyUkwMEVd39ZkkVlIzL+fYQec1DQZWIEIt3TLmpArQyz/U/VCqp7pmDTSc
VjuE7mbsXTic4YKdLg/Z4qvGplJz2u7CQmvjcC6kltRtAzj+ZYHca8N4n40+
z25PSVBStlC9mHPA+3IvGKRUXxfUvq+qlQCto/ebWEyQCBpZKdVkl7UmSAYd
7rgS5RIIglAKSNRVZWqrSlJwItcetUejN+nBjPmZGZw2LtxXjX+wCHZfW2R5
RuWilwG3e6pkLWn9mVdNfqbG6dFWr0a6nT7rXyDZinsMY2+IHdtKFhofSzyc
GkVK00gPQ/caOknyizO2o3A/L35vaAIDAniCBXSDbph5zjjQSZihiodF6tLF
vziHR744SD5oCYobBNi/GHa0syQri7+GhppMERBZdEsqlcqMh8rG0Si2TF+Q
2XMyV5Zs9gTTWiyE5RnK5Zi3EwF+Er4kug+QP3lvwdmvg9B218F06RJYRWSE
7wDQ8n2Jd1aZDvmkxhNG8eZOe9KmVdcOyQkgxKtqy6cdCSWsKGsotgufhQRL
HoyPK/mNeNwpy+ia6YSRj63CfxXZq8mz1TcnSgcsX2133HDKjsH1mmPCHwdo
3Q2c98NaaNUMumLoL1Kiaeqv8FNbqnpCkasv+BPJjifmzjuR3lEKRGAuScLY
lYhXVMhIP+N0EdtHOJqFNGn3dgazcs7xLdPMcm4znH2sdXqouaUZYJEaEiZp
CNGbG2ULSm9ksE+1GB61WxaRIFI/0FBULFGHfn0VHCpTnoFxdN8ucVZuE4Hw
z/3uZw9rLzGzykzj+A/6ZAkASdS56YrJ/6UxpKECafrGEhaCbzLP/+WG2CjJ
KI8pFlq3nINFIIzt1J1ERZxuqUwfX1HvluOyTwlRmhQcH897iPrz8OYneHJ5
F5Z1TAVCH7RKNCTi+miCWw4mVgnB/in0VibYMAo0w775NI1xzh5uFxcZBPje
0/OWQ+4olpqlflujDIHsThIBcHCibfX59VFMUfRivyygRsn54MDpZVIP5/kW
RLkzF5Irg/14XU0FTGHCI5Er7s2GpINGcg7MfTpMl68q1vFOauhbtzb5qnCq
qu2xzkM/Qm8hq566O5p6W7aOO3Je+8xgkrmGDwZkWP2KIJchDQLFmcI9hQiw
UCesqPxpuFEv/idO2DNnvTi1Q4Ccr2nuZQDhkDsP7vkaZd1HTJXvM23HOb+F
eDpkmk5PoHIdSSTJM3xkP1UTcBElTaeR1tncjKVR0NE5L4BtNYqYygeMYssy
PbEwPUCpAmn9lntMjJnjpbx84TSrhmNd/N2WyLWELop6lwth4ymclny+aGyY
XH0axzLR6eDJWCbwTH7krnfvnMQfta9b9YJ4LTvw31lqEawXNB7yvJuQo/Nr
hprRv+w7Ww74u8pKJEf4qkVZHD2gjZMOImEdMlpJr7R0Bn7zIh5+I+HeYZ33
PaIdpXAR101lDXxiXWdGq7mLaLUT4JakoYdPelsj/4auATZwOOGQH2vkHPPe
g4d8qjbOMiJzZVaITte2/R1nsSMf78g7Bf7vw6Ikvy9adJrXbHrP+78Z/BqO
0JLeWoPsXD1DgVQqq34PGJ3gYY9lCiD4fNdynXn98/+npHcpHjEpT+P+Tf3D
h/l8zf3qM3AVNjN6ZkBXKCdASEnatqAcpejbxtxiz2+lMraWA0NLH8QZzHiG
Kij4LxLxQUf7rRQy1yTNCbKQO4XoRjOiH2+C5vX2K/dzWrtVkPWqfGJh6jC8
4O7ARugVDIZZJEk6AYBf1HRF2uLNtNqkEk5PRdDJgJsNC7S9CaoFk/jgPfYA
nXdwOEPwBN4VHhZLcoLqAK95ViZyGWjoZNlMJAy147z2+yDXhpNJz/zfBpyH
nGRs2UbOFY7Z6t4Aqtz9Z34BV0xoPCapz6JgtZN/pASDThXT5tf40PypwjSa
phOtUafM4OI72LIaKGPsrCjjCoQssFAojo9sGvmsho1kUsUBlj8FGjXcANV/
RLV5ScyQ6VMvNo9P7Gb6n30TDqMJG8HaeQxJKzWajKBDz7oDM/8r+IMM/goi
73eIV4Z239N0w/Yv8w3nCgOPsg1KA2lvPTmSHE35gxk121TT5BbLABMhqeLa
6jqbvLdMkvEP14M91fzO1xGCqLDOik8oi4MeNhkOoc60fCVDTkJ55nIUbAxL
J/FdTLDd2bTjAihdM1uYPSAhVfKbF6iyl60Pv6Xr2N9pzWeN7HUORAd5AMh6
bzr7w4cPLZ6AtMVZF0YaF4rQyGeyGdylXemn0RK2Hrxx4MEv0GZz8itDutDc
IiSqRx9xCSw0KF1FStROWrqXUMoHQbDz7XtflmK1WyHAQjJLMui8tt6b0F+V
DckiYnn6xYHh9eqFycPNZlbUaLefElxWC7Q/pzYWPoEnyMqvzpdIu6HCMatQ
Yq8y6z2NV8EPNAfD6PnBpX8ujiBhwnoSnFdE4oYBd+LLGH/DCl6eFkf79p1D
P/hfP6i9V8y90CPy6UhIAVHzsHqDJj+n0jpkBqIwKGm8iUKmAw9MvTn+b2g3
9c/V2sZ51Qx7OMHJE2USxOhv+plcEh3/YuUflL+PydDi2t9sa0kNBhBKyUBx
6oqmjhjTBSxt/25d1Wkivkv6xUuCkET4Zat5OLrfxZhwNfjZlgj8sB6hYO+H
b2cib7R7vrgh5fqGfOp7+69Pg7uNOoB6E67nKL1FiT0wKKxBhaHKFaTcLoQf
oQi5KyxnZ+J2zYXRs243ik9BwwzIS1iNfHf+HgsB+MFwvRYlnWFfOv0iTNt7
tfKsj0WsxXVjRSHlsfeJTdzXVCSb8Qmlxn9fty9ubBak05ucp1MLZveATUiL
QSR8JsJPqjm0FU0QmPgOC0FxQIKZQ44JVTD276C3K8StM/we0++iwtn1lwED
w/uN70uF2Df7DSYlDFBoY5gaDgthenw6pmYe4fjf6jBioHn92Ab3MkYfj2Dc
ag8nf0n4GmKtzs/iAaUl7+45ox/4cOEUMR3EhETJI3y28maF89EZMcBjo06P
oacGL8OWoyOZNWJTeshMQWr60GbbxsHai02tejItcW9zWu+G4KKy2cwPenVs
iRQG84qknGJjn5E3zuSsZ9UQi6XuhrtqsJ4WqHJCEn1FAB5zo4JsYZC6FfyU
KX64C+//BLmMPbOL0VX1ls2qSzWMHOi9JknhqfKg9QW3xG5hdrV1OfAHj6Ws
ZFwvVTXLkGpZ6OGODXE7ynT0grL5P0zfR0Cc0xupsZByzabzDxd9VwiUk6qj
SS+QjSdearoVNomG3SbvWXvZ5LO8fACPlBO+l5JftjNV+AX6pNngZV4+Ausj
52oBpTyGvrTt1/G2QW36tbcp+8AN+ZZd9B2ItpUhHBwMIOwqjt8swNJ+1xVV
SD7jmf01uWrQtEwlqxUqkekcP6/vvM+ShH4l5v/yb9yHqbOw/KRBZBv7FWWZ
9kYOpQjWtAbe+75fwl/pnVSgDIPldee5+UJXhauH9M7PJouCmaTs4J1wlpkn
jYsPti4FXwRCJydnhsK/jQMAUrJUXGyrayVhhvmvJpA757ANxJkvEWNw6z5t
wI7fR/TSUuyyN1ZwIilYF5cR2bboNYzdkBw6tv7yL7km984+wIujhzO0AsgW
G63g5Wv2N11dFzfgLFNAwhcCijOM/KZsjJ2CYIanct3gYPz5sXBMVnGL64aR
OooD/Dxbc7i9HdbCueltS8uzr9TZcx3v9YolwCr5vIa3G0GB4UIzA4/X1pPO
UBLNRR4eSXVEkX4n25ejlWCyUpvqwqaJ7CqYRc9NX7dXrWRTg7ze7QCM36rv
ccyGOmYpreGI0FfzBDcAAW0yCnP2PRsOizzb8J7yHoo7k3XZHOGV89vSfiby
PgZ+WuXaa36wV7b0FojBXaDbfwzinG9nq6KhYqzQf5DLNhF4KcBc5FQIFjFt
erbWI6SZa6hEgO6LAGN8bxJtjSBToq7KkhdQYbHnn+/gyZkVZaVOpvrXPe7G
jkTm7sB4n9tegzsuWBLsNOcQGE31Xis6m+DANcfgDPB8J5hvXW27j8y9dHqf
HECu3BXNVS/duwu8mOLXavZ+dzjBjTc6O+1BfcXSe8sbtki46cmDnzBFZ9/C
8Z/JzOmiVvOlFUt/pojVMxCqJeqABtGCy6CyUeUpISLWXFpzYlprQB5qoHkc
zwL/twg7T7WBXx4ImmNNzyXDYb01EaQsbzsipfTONdkB0L3A8LvR5mhCXMXZ
Xdg5nyphs+gJ7i5mlU6BAkl+AE6jEhaDaB2xPCTbZ6w5QWVQJDtvlrOziFxl
DnUlCF8Y34QGDveu2kjFabynR9Lrq+xHyqtoVS0cTJ+AZPdktOh37r9Mwaua
YtdejkaP5A7Gb/THekXGFrGNFYjCg8FBV7Fy2DcHx4ZpI1tl2WGEtrNyAVCx
Ir1nNCAP93e5ByUN2xhwsoqrSAuSblGZSycAGviYSWrHn0dEhDo4riEuN25R
dLAARIIw/Uxjfmki37DvTWPC2x/hRtzKyqEJ4iTA0GCiXF4hmVCitSt/fold
Ph7vNolb5oLoXGQM4AxJewenmCXzDDkarrY2A+a4wPPpsDeVdoq3/1ZISVXU
wjXCAx/6av0RRTxWO7XR/6Ky2y5uAr6xlHGsVmSahJCkth0i+HK2/LuCVNWp
mWT6yCEsrfSFTbWRpSgx4+0Aj18dGI5iRfaV3xnjFV1sYFQGQNCghzNSlnX8
VoDLCGzreP6lughFYQj/gzMdma4wQN+eyfMlFa95ngfe6gXJyS8lfU/sNCZg
9A0dn1lIkhhaGHKuQdyK58jPFtuLxlvcGc0IEVr6ovo7l6pebQ/QbMr9v7Q5
RynDGeMDQt0hLNZ4CICyJDlqdhDdtZ0pU6xrixsklFUjy+Achw6Jvz1aSeZL
W3BoKrTTaeibtLZFyS3Nr8RrRe8KQ5iNUQn161eYJkifXGPxNo1mHVe9CUGN
SrONQVpmFyWLg46wIfe2onIOIqrf5PhdUaH2jyNn9FiGhNOD6qXyiig7xOAZ
jAP+OCN5kbnrPQgRYSEBSk8QpHyrCht78/r5uAVoASwpfCUv1Yma6KhO/5ul
xAXKtc0Q7GQmfM82kAJWO6n8ozHsIIUSBVNMDYVYWq5XVEHkGPylWYISE+XY
yIVYG7i+Fl3df1tn65nPvrhE4+J4EUfI4PFBmBuwTJapUfg+jZ67DANHpsIR
R2+KVq5LZEYF3QQFl/k2r1+DGwraAfdaC9YljR14BVTPUyz/z8gkt2rZXB7a
SgG6LC0jriyy4ygkvWx4fzszNZfD9NTyOdC4WG3+l1XtNKHChgJQbsSjCyOg
Q1ZSsdsrau5oVWCv8XN6ZPTzObpY09MGHW9gM426gzd48Z6aedDKHty5X5oD
q/HUuCmkZP9gy0aNjPfLKueNoVL4+T078L8xAx7rFggGG6JdzW8ThLx9LG8x
Rp028a7zN8IK5QS8dh/XjC91xA4+xe7cxWP10WlPtNdY41hgu5G1yvO4qOlh
0QWrF+oMzhFYeycX28fVG5dnuXCRGhvrMTp9TTS/h//vQYN3Hze9YfT9quQo
nBYgFZLvQG2YthEe2SKa6VsEMfr5O0oVSQ8hj4ZIb3sdH6byVK6oDcwbclr7
2EEdSgfcutcE46Z07OXqQe4fn2tdSGKk1i46bsoeeTKXzAbRnQOGO5/pzclN
54V8KxElqI6Uwa/iKh7kk/M0UFf7kqtjFJL3Cg1JAdewNFxOxhG645Q5J8xy
uoPZWS1rhEPa33aCifKjMGvJg46/GIjnZOKSjnfYesvQOC8kl6vb1Zf7+2Lz
d6EVpoLkrk8+mpO1EwuzX8i2KJTw5AdA//yB/KS9vr6gDLjOCdAqUe4sIC3J
gvZ0oNE9I0Bc/S/FwLnCkNU0Y+si9V8EcGs6X/OgYX0p0Ni2zesbrN4A/0WT
BPBE5AEplTZ2DMEe9ahgU8Y00udXv0/WRlJAtq/Fopuon58nVnR1PeXXEMU4
/Op3Intumc5iEWFKHCxCS26OMDxB12SSvqSVmq+UFOCEGncXOCDnGt3a2JtM
bhmtwTTU0w8SeLIkMHOdIIiejV+E2PVaNzHdWbSzakqcqMArvw54Y0zaBiKV
QcFJEfxa+V0+2wkJFshD4RJVQlf4vT2ZDhS5y1dbWXWGFKe1Rl10StljUFn3
5Z5VWk+3wLARenaB4UoWK+gxI/mUy+tAhSz+2dkXrDVobIObT6dljhoRXCpk
c1URmlvIRPIXPWHGY5dQffQz8kRlHeo/O6zMQmovIFqvdswHkDMKy8xvq3a2
lWClG5Ydoc1aYjSEGNmUPtsG6GrnZhcmhlFVLlVCj9NXr/+NNxTfr9LERH10
Hl57ANaryCDQGqtwbOasB0DHjvZU+5CjHjrEQNBeri1XRAzQKFuH+6XwaT6b
LeC4x0GGPxZTSfXZ6RFNryVo5+h/nxE1g3cMdOCyIRbklYkn/x7ScghXJkqa
LC2CzzkwWKG9UZHZRBxwOQQSW5EtBYXgbCgio8p/5v00vhD+1DTlpFSczEd/
6V97U0cOwWPC133l1WPBxfiWXJhxauUSX2yLpFPt0XIsp7vYY6Y41WlfaBnQ
CEkAHijVFnRidy54SgSm/m7e4kQQwDeHiDUdHyTFWrksgb0ERkt8TJB4vzgb
hNNresG6URa9AYterfywYjmsPg18knB1ZYmrhZX/9xABqepXTQWr9h4xsSoN
Gk1LoC6e8WB841ieH239Wp4x0LYRcyF3RWKSE2EPhh9g8FV7B7kJ6AbfG43e
hqe4t0dd5NKY5/PzpxpQ6sEBuKSl92NX0Lo3QU7/jEIvA89JiT88cPXssJEP
I3N7iXXYiADijtPe2ppQcgWyEHDa0GF0y6yimC5kwHyAE3ffh3H85l5C6PFa
d1TX8zVg6FARa5BULWK63pbr/ZMX/dudE0R+MgeXy5jDaEdfqKTk+WC2RZ9u
qbaNPceAyw/+TNTgBeuO0GoJdrX/ozPHELSdHhP3ElQBJS56FNT2b9IUXVVc
uPFf18Rz8S8Bsk3rYAsIkkaRrTFQMz2yQFvt6inJB7lPWOmmCjpkAryLsxXu
AhlrC3FJK3W9/iHzNU/Ewm7cy5DBmjYDDXjr3Fpc27X0e86kzBx3BTxnI0s4
9RfJPCc9KSjmFW4+fvPHTH95snj2MRyLWWBFjpAQVo48wpjB7PFpTowwk5up
xnfR8w5akZYL4arYFcXNE7wgC4fk3lzarIiJKR7oGEYywampWMfontlj2huk
1m4rEAZNtSd1T+ZFfF4t4KwHgd9sZLtrcWev79eVt/GsdxfgRh023Ty10BNR
geGFQ+28AvMS5GskrjNGltHTs7WxLx9XQFLNmo3613LrW/OcJvgBkPK221tF
XvZqTAaWabVWIVJQNzxlD7TXdPmNAJZLAgvLnreNBaUDgbqMPgqGvnPYah3M
UkolDk0jOXfjcie1DMyIDanfU8HZ2mPmYD77T6jwLnQ5ekgiMOFl9YRfc6xv
5QL5ruF23G25Ozj5p2WL1hhtGPrpPosllnrvZeXVCgTxZCF5l4eaQRsGRF+F
rmwakHF6/nfh/aC386dj15PO8mxjHCmfGebkXL62okWKPXSigFweaF6vbBfI
P/Rx2RY2xkErzS8iDvVwGZw0PGY/Esga1b0/+jtL+ElilEpKprfDwPFyYNlx
wxdjYTANJdxNUCp/2T+B3s928JxPd7kCPQFISByFYbb2sK/RmveR+EivVOaE
xa/ThDIn3brh4nH8UYAP8xFhuh43mRkGSvtX7kHevbpqY3z2QP83ToNAGoBC
cOjOTL1D59ADeFgbuiJiF7/PBkY5L1fEwmSK1qd8ae9HlczlOyqIN8FovmBu
+LQsoTWvGwtMdypYOxr9s9zzbyKbA4gEWx4+WVEuJBzkNdza+ETuRcp432kB
UHIzS7Af2ZfoPQLJnwzjF+YjAy4ANgcml3rrz850LOUQqIdaXfHixawsX2cG
GfplvnUEPzLbygDUlR3VeDlfq16250a9IITGcBoyqU7QCh+cHl2gScxOeeN/
LM+fnl+FGs4+u36UTV9iqkXW8WuX2Ou3cRAXE4Hph7bsp9glFGU5cZaIWO8n
Arkca96S/XKrBJ9p3VEGc0dsfVDQxOC4mp3bGlwmG+YZl0kkKGVR/4Pq1ZvV
J0qiFo7C0Zzq85Y/5+8D9k2gKZAl4tbWnOAGSSQb+iwYtR3/AbR0jsg4mt4A
LXqFNIVYNwv/Mod2iTqRMB8DrMEeytd0ud6LdqOedu/ZHW/cfHRkwzZ+8kT6
wVfCNFuuJ4tArF17GtrfP8pJtee1dYNFJ55z9cQ+UBdbd6vrE4okvoN6UoeA
fxUtU+aHrrixmrFhn11c8gIrctITbBcBowpxzXcBBSaETSLosvOBk3q/vaj+
5pwMRSCqczxK95vfrsevfjNX+SQ3IXyU+uezt5UJS2x73z/nhsu6h6VvzlY+
9n/vcRxrr/O+Kd1R1GSKQvZ56L3b/BEp5ktMMwh/oLbi/LCgDETt5r7Go9GB
6/maxf3lqlVvrYoOW/XmohTdT7Gpjg/JReb55jwXAbE1lEzVlSjadMJ70ETA
zVzGQNontkGCBTa1rflJ9rsHgDJuhyyt0z0/eBt/2hHn3QLYZOfgUGNKjdTu
LWHomjA73YH94Ldj5JYLsX/NFjcgTOvWkK6a3YgYoku9vu41o47QzXsGHjcn
IRrbNvACGDRdgGh3W4+EI+2VWmb2XikFPMCCYGWZW1EylhyzyzO5eGFdeHZd
6c9dKFGO+e8NbQrAQH3yTcFBS5GuJYi6A/rhRRzV3ApJ7BxXZHQQhAZ2MGnk
XWOkAXu086e0chaEfbxOOdKWbNU6IShcnpO7IyvZPaDInyUoJdFSY8Qgh+Gb
oxQlUrRjxK/1NiJ4t3jT+sOkoLmNqgZVoDLBH3VvCIESSJs8nJue7ZsVyrPK
0FYM313mi+SBO1yOSW2dn0SWLUGADT4buoZjR899143eI15n4sIsixijTtBg
/CYdM4QymxXjQprtWmSc0IgkPsasJOIgVbCJ+gRlVsNUXnPruw4x7boA0Shj
cFU4PiI/J1dBDrv/AQ5OEDweaUULyerIJc7YgZdOsH2oWxhcN8PzMULg4A+D
o+iJ+wiyX0fJmkodLMamY8PXjzGE7u3MwdPbJdnUvCmphZrKMyd0XzWnGCyp
lAjd9CoxlodRlPcxYhwZAdUcBgS54pXI1r15F3AmdjV3/QBptMYxCEgN1tn2
NpJeKZ3NDaHnGn+7sgBptOv+YxXQvZb2VqX3p5yHrKTmV4Z0iq6b1t4k/Cr/
iD4zFi+tRkzv2WzS68sFk4OToW2v0+eqqxYDF4pO4kPew0TvBLBtfXdjPbeT
FC8uqNQ2TVgDN5StsUGPoHBrFgGnfPa3amMhs87uiL8iKkd+Zeghh4EHLv69
L85MtjMiHTtkH08kbcl/RKEKJABkAXyUu5klJFiC5LO/P6JUHWKtvQ+Gj6to
sU8QsZVUZ2NSJTxiadXhsSYZn61Lv37euLZcFaRizwStFy3ABrbjMFAFIeiq
CyWQJaAOiCeObBbq0SoltYFImJ31JfxAkJF15oGP6TLcOjIUVMa63wolha5l
rfeZFnWYNFojpDMSqktZhJTQrBlxWST2/eLzupjT0a+rj0EgFMtfQqE2lzsH
GJRHnWwnzB3Miz8l12x4kKs4nw3wxYciS6I1X1eApZrwj8BewjuDrXI4QJWR
n/zT8OF3nebDfoEjUl0vNNv3XhOOiSQhqI94f+bcCy2k+/NKwj7CnBkvqxh8
bFWtgGVoU3cTNDLxQ1FkQ/CHFJzZeioTY+2Ea+9VHPPYtiNRztgBOBQqHxP1
/+CVz/5QgZLa4sTCCQmCd8vACPrpoC+c4qO4/abn61KaSVZEGbFPfwlPOZEB
iKidslFLVs817bHlShdOvOdHlmJOtwE34wm22PfCz2oK2k6NmXihYhw26B9i
j9VopwGPC4zSSFR/j283hSfgdVOti41nUOl6WlqyWpXRVMLcPxieoAJAqPYU
sd+mFuHlJeZtM3ynlkHPL9tyhcpAAR0DGyzGfqXy4G2qSHK/oBB2oLjYaqSZ
qaQE3nHpwF/UEfSlg9c4+hMNcwAke95DZWT5xuqgOl3FVOsi211uZ7pCSSli
RgDYXxcgitSTf+dweL4pRN/6I+o8cFf/z1xh2mCZ964+vJvfuSOy22R5nONf
PMxEkvi5x1C43Ke6fmXasiGJQY0pjXekXc+uf4JT9S1kLCQljVyzTUAc7IsE
xv0Vf6cd+jFYHNwXZMju5oaK7ZCYgCioX/CHHCpq7SvT3ar8/FxQZV/4zmRC
peAvN1+hOH7UKKu+a9CZzVcTfQlmAq4I4LuTqie0a+UpAzsYIky9RkCoEAjY
thQUSFCantWgy66Arv2g2mYjydg9+IBjGTypneAIHRo5UNYDcvG+rZtulDz4
VRQILxzcaGgqu5aQy+vmoNf7qLeZqvjmjKcGptqMNetFTAS70w/PzltAdXhy
72DDFVOYanCDdisFdbB4+imoinAH0+WEIZggTlsZ96LBqMWdGqyWek2rvCIm
BMT6Cg9DvLDRim+eQa9N7fod7L3DYziy5oTiHAf42YJItIVyVvfcVu5tQLrV
pOUiUzzJ91iQRkeHOA1UDGbVO3x8Ack553nPwcoWYmKNAjhby+AyBQsFWki1
wiAkF4Ro3FAhbtMuponqW+C+BCQBIFVjz77fEZ7/oabNiW7PX2ySMc2QD1sy
LtxS8j77II6ormnH5OTp3wQRlV3F4VFxnWZ+3S7lvbNRte2bVkaj5tqKyI7c
Mp8V66VvXUvsnQhBZgRYjuxULWEbUzNG+qkzedkeFw85SdJUM18/H4V8+sx2
/uJIz6wy2ORlHVVjmbMAknEjKU3buvW4SC2ZaQbQZzZsQ8oR1oR//f2chVmC
dMSP091ZgsUY3mG15D/T99FK0DY6X4CchwlAO4Dg98wmUQ7yf2spZW4fNwO5
82Uc3qIzCgEoYPOiljkzDL868zIXGBjykEaWp9yrGxKFjrWaMG6h8j5wwH6W
UDKTzTZZMEqhGQyrsrnk3rwMUnUac3yVdM3KktcOkLjJKfgYGeIjZgsW/2qr
e4dG3eQSmOwZMVf2tccy99oJ9Cfs7AE7uTbT8enliFCJA4KIiqfMdwa1SW6d
fEY9ecjVR/ObKmI1BDv4b+3zT566Zt5v+D9oPe2gzPxI62VdlK1prprtW2d9
GCt2KmogPhYXr3f9fdFxHLRgPqHsDalIakyCa3vP2O7F8p3PLAmc+B0ATXQD
1jSPof6wRxyj//AwebgikEdu644k7bvxPGiFL53iLklBHUzJPkrEEtb3lwRi
iYRfnSemCkbNgkrenQNRyl7GCyhwIdXC0X6KRT6CppC+EpjUJrAmbIVaSO7u
IjiLVnaIsL7kuJHJIKmAsc8Wr0lb+HOWEV6GnjamlaDF47EToH/PUzXeS8wL
aJmqd4+ZJkyNR6FBjFw21obed9zrDeIMfZW2CD1nTYeGTfaMwZCF2+utOgLl
Nk0IiWsIMMuE4XkOep8BvLyBVTaXTU++ir5I3ej8vdDrypf/apKYy2fGBfK7
2EKalaxT6q3alpBULnYSUYnvr+elWcXvuNSa4qPsm/UFMeCa7edoxfPzp+m6
0mfRIj5p81ZuXzDcvvymNgHhSpb6KsIPgSAxwTxlLrQ8FZ5AnoC6Q5CnDyF0
JFbhd8IRV+FcNFQgJdMTQFgXtvngxKiUVhCaT6WljdG6b09TTnr/B654BXS0
UElmU0KV5n9PNdOGZ8+hbzo7NRUam/85gcZdwL/VQStxprsQYOpm/nAMT8O7
+ywwJTiSVsl7OjaDd7E9ZD0N0RXK1sBoids/yoShh6CqEjQ2xhr4bophJSzu
wrKnXCaj+QzwCvZV2a0ytlxqIB+H/lFqiOCVSn03HW21R2tf2LX1xxgjdu2D
x0j1B4iSWth0VkH7VWuI9pp+ABA8qgUqwmK7ITlVsDDmqm138eatWubDo0s7
Ab/KyWzL4r3++wyO/jgoph4z5xqQAIUz3O6Ua8JA2H6hlECtKObIptbZTFRd
6WGXdBsSrq9AKvkqhDiY4uhtQSa6+OUOUQIgkoYwQPAroElonE3PeRtYCeCt
QbiGqYbsr6edEUf3C7G2f9jm+ioGV/AHCuetm5fEZcHrKe/4Tv4ZW4Pmaqyk
E3YL528FyVubC5XmgHKHCjqVhwfcseRE1Y8gZb6JjlqHLTAX7Ansk1cDU5XN
wrwRIv5/3isibtvOF3bvSbrtfrkN134SaChBYsesrQRldLeEOkhu42A4rp8p
LNc/BXZgR5kvbNa6TySi+FwM9UxW104QdM17Wat4ChEWvH28vBK9uYWpWpY0
PcgqC8uux9lPrMkIS6DLW1hVFqb7S0mTqmvdnuHi8LxByUweMM4bOGpNEqUq
7j7ZzjJgtMXxTulCXpnWXUr/fXBE1NeQroCfcVzLbQy9pXtwz77iCk4ypugc
8UlYOvsY2GQJWsqvuppiuuya7PWsGe4jTLcOXCu3VtgEw0cKqPcrx1cBaqLb
6kQIhplvImp+thjrMHdaBRTwzC0mYnch5ZhSJjlPYiuPWh/6FYuqLuazyjiM
LZ7YupsfXBEge/rYGIoUE06k55GQNoTjClFuH2+1Od1pP7y+4bVYZ/0PhXTQ
NM2dskts82wIbYHgSdPSsitT9h3kEslEgWiAbazq9YAVARDjywKelQpcaVM1
wXPdN58w0AuuOYXtY58kIMmaeQVjhSavvIwABCr9VzqPRMuxOhocASU8X24w
ZU6PrODVQu4P5v8BhPIU7Z+CKlzFkyqvKPJvAPrSj4y8gVcLujilh1PL5cq0
EhkH7NU9rjeF4AmRVKspG2fDSMbFgO4jsy43r5dLqByC7xizfwA1FnIWoPsv
yjd3xtJXC2QgUkNBuvNX0isYyx2BZ4jpFqKvYd2Wn0DZ8AxhPfSE7AyxyaNn
QPcc5kJScmLg6SSQ0wftI+ym7Il2PGhGi7FY0R8eUo0NxjV2v18ZaMzkg8Xy
rV0OCTxoANB9RSX2HILM2MXIhveDoLVspl5NRykbQ3/wzexZ3vy+HjuZzyOS
bsEHwdLvbACklx2TBdHQO4lu3yyU72pRZ4UrCeII7a6hVVqI8kaXJk7OD+4k
JGGDweDG7NW9+rx2e56RyMs4jmRUZ19jYLDjLS4w6JQ6gAXdU9Hk1rYTu4Q8
U8NqwNPcy5VcIwmIJVXLtDGJ5eWVk38eR2zghT/F3vFw04jvDVldnfLxmZST
9615iDUEgNu4i9g4KXYhj3wlvMySd9nK6UlvAA35TVyNvE2CzJGP6W76cRxR
Ls7IHfRMVyf+i9k742jMb/0jG3DAPA31g4Ecr/iyRJ5wE8g07N5Knt+8qop1
H6ZYirW7zspu0COMhifRxg4351QcR2IacSNfVNa/8JiRgn9u08EEGFe3F2fj
PWUvPGs4ZHzixYDKedgX6oZcIlGkX3OTbkH7PA6ToH8JUc7sepD/N3ObFLLg
j6o+SdhYkAj+D9HVAOSW5zWfx5ICodNBAseYtoOmSbtJdyLteCOxj3ltsolx
3/L9CUQZSqTo7WhtN5787ubFu6mxj8bSRXEVTTaAI3y3UTF8ZUraeSLb5+u7
Di7fbl7W0GU6HvbX0DK3ZbpQGVoOow9Idj/VA3UG5/A7ThN421ek+eDNe3y6
08gxItCK5MlTTBOUPflNwQHJVslmzqlJF1Nt8AWOX72m0CMoa3JdokP7mJo5
jRORFEWqYp8uc2ueej8tkqShCKXwZh6Pnatj2GfhcJYFdDL7PDHV5oFiYxsG
6s/kw8oFs+Ju3mjoNAzQ+w9jj762/0RO7jjE2LsxaW4ng1u+sqTf5SlYowma
o8lIxKGE74fW4fm9z3y91iB9MFIIf28eaN6StLkNBsTbmtoFbcFN5+NhU4Zc
aJfY9hdfFauB0CFAdkbz39wb8EEC9/rD/L5hbVJSQQ+QrK3VCNE4FO3ksDV6
QxpQZIqYDGmpygowX9A45uG3g2li33IkGTO2soPNPf825NXaG4nuNXZHYxZV
4y6XQhpiioa3CTU4sBGc5/U7Ejid70/iOrQS/L4KUykPZ6qyUY9oCfzaEDFz
IbNI9oek5lJXCEVqGpdN8s/ieuAy02fscMvmrjPgaXtxxfDvLwKmttWBGs34
R03QbW1vsm7i0jyPskvQH5lIsZadGGvUlx7XdTnXif3+bDsWk8uBwSFfU9V5
9axd7B5nYwiHb09gt9VIOwDQCoLPQhmVhfjzJcIflOp9HYA05qYbmnnlI+f0
sSXuebAd1QGwKj4zCJMMeIJhdgXVl5EmFN9SEgxHz/Wfd2RVua9lJsmclD+F
SGiUGtPPchhNw3TmZrVUMYTCuj+vC6J/B1Ik0z8ncu7NvgXxNf1YFxGsZEuh
GAg5ER02zTtCKjEEr8AXNYEAUnlCkbFFAemJ+0jVc4ymvKqDNlxXJaQG+V3r
HZZ7DjNVDNdh91n0BgSxTDOoKcqE9oyGfAc4bRDJMzZza8j1WMNQfxNUWY98
yld0IObH6QAwpYTlQAZJs2sRMxLAlYhiWx7yGZSwgO+JIr183k64jaxalUKt
nv1LuhdWmMVGItt423N4qw2VAPW1M1MaluWQgV/pqMCx5CfP3htI7uxrJbVQ
P/kIuAN34AYMnNZES/3nZ9nGpWQ3cNX0NLW1VNmuaZWC7ajShngPJ5UbwYlw
1fGHUpfO9vmKb/dt8nh+uHHBlr/uNFjA+1lFvUsuBi8n4U+FhbIWBj92Ry8k
b+E4A07fX5wob4PqDEjZG1w2MzzpVW3VPE4ngCQYJsLytF4T7pkYJW2Q7TpI
ivmYI0Vug+wnyzQ7RXrSvOO6TKfSn2gP3wwe9Qh57Mtou1WKFdXZY3wMqBEP
fLh2qD54rFWV3k1b/BML6iggXD0ej+ataDIFaPewsm2uVvVfO4livka3Zj09
PBjbHyrfxuRZnspudLJ0174KW52FTAlhVE2zYGn5XI69aWTd+YrX9jXQXBIY
O6QGTYZZXz5ihMFSvMSFfz+v7jRjt26Z2L6N8BssiY+t0LC4rPnu+MdBU567
UgPO74smnZLH8yP9LbLy77Uj4B+2U+WGa3237sqgHC5Gpd4REdtwRqZKjbpd
B/Jbg1Tc2/P5un6K4M6wxG9YaIzZs1w9Ccb5Q8oBsL21K241uQ80feVxbNUt
0IM3iBD1ZDGSJQgOXHjaHLciSCPG0Zhp44CWtvwcsWkJtXUKcOJlyD7hG/Ry
y14k8ZrUQM96+ClRAjbQHxgxx4Jeyn1IYkfME7fV7HLbExmV1xaBf0Ome84v
FC6OE99yeeacPDYi7SFDGCu7j6pB7B1shfzfUugjRb2IDgjV+10GqKBkf51L
quXGfCA3k/nFNPg8det6Q44rdbWc/BB20MU/e3hlgBJpGUCR3Kz05nV8YSqr
o4PNJB3dLxdykmY/8B+FnJeS6it+4vCxaYPIU+pokYLVjWwfeavlUmo3uqYa
r9Z0FPJw5ICgHlVqw98iublf4UAIBEETSZvW8866OTZ3JwVSRctomTa8PEvX
nLVPWv6znFsMwdXv4F0UsoaI7RKdpi4u60OTq6rL1U7WTj1nRV4fY8JMvqlv
RFC3Dv3KYPFqtHMuxHgxUmZjqMVzp3MHU95rYRw5FtlL7vm4ub5yuaLBVokT
bwDInCfFbEK4O6NWe4qPueFIOz5JxwXeQvgEGYMfkSTw+9oE5UxCfssPP7eP
q9386w6TmI3iGtOLnO6LL2hj10Nyi873sywyRMbjJiG1TOTvFQp5N6as+F45
zvlDbC+W/iRl55OTQ3yodE2xx13GfVWKsLSjSi9UPftpV35ghG29EjC/dMPO
g2h9NmGb7zB/YdJeGNwzYNHlhLQ5vzSDBgaDpWLHfwH7gqknczI4F0jpVGcl
ZkxElMvPtAQURXdS5xlN/s83SghcNxhwZnHYLFil7kCk4XkzKys7CvcGfr2q
Kq57Xt3u/FcNaSeVdj7I4xvlk19NsEIPo03XAjBI7qGWSFem4GbH7aWcPkB1
0OQEKC1Fey9jhJIy+7mtAMjPEuT8H3zP3wOiS2mfvk08ollmntsZVxvdWEjy
bvjcWoGZKLkL77cf0DNc+9WGIg3v16tRoeLGU/pjBhDwB/W1dr6V/2FyQa4D
l7mORAp7agrS0yxr3MxSXyH8eMsABnTAbY5sr+pXfE776hwZtapJFFynNidM
q9Ixv7SsPEU1iMx5bx4SdzN5HOMQvbum/txU3wT9yJdz2nHD1K+iS2Mo1HyL
b1WA+u9dNeFACwwg3LkwxoShoIjxAxnmJubDEzOpwEFdxwa9v9gjhnTPdgKT
wx798lo1eZZK0d7WK6P/hdjp7CMFhlZsfm/e9exoxv7WRBdPuCI4+ME1l2gr
J7GMrdB21NwiBeoELkjoAQL3sH7nNSbhSYd6CyhUxsS6d6zwI7rd/fp8DPl3
UotFKJBzqOV+GTbrRbYisLM1jYbEDg1ntVtz90x+Wd7MqdwhzFRPDHrdN+i0
TRVC6CK6YCuMa+kMHjOdO5rV8srLkRSPgv8wbwc/tyHUn0yC6c8rI46bBenu
eYAKoff4AGl8Dh2ZDvdLFDL7tr1a1ynVKafWutoXKY1cVx5puZbpGQMEILPD
bUEIITJWmaD2wBpuoN5idAJl/6ER9JdctGUkSWEAfofDRXCegjZcNGT0eoLf
PUQBDJncFluDl33zTluYz2ftUu2mWjgLm1SxARyhK0Yh3h6c1aHLBxpDGfBG
hbMgOw/KPtys2fob+cuaiZi9eK1u9sUzWDoczEhvjgzhLQ4WXVDlTYBdMuuc
aOZZGfj/OeErUc1C/dQzZBsd/+mo+AM5VieHzoyx9KMxgO0Z7U/9U32ykdui
vrQtoYF/v6dHglnq7PNj7W8SqHdbtQjlIQcZ/7HCahwNiCdlElVU1jBv4ANq
bduo8cRVQf+aoLZSvzGTUNn04xpRza/7MmTYxU6//tW+oQTLV7OCIs8ZfIXn
yHSJtGCnz2Gp13mDRgOntz0/XfJcEcs2CRjUJCHX8uJN7zBBLoW8sceqBGVv
9xF+oZiGByjYxn4u7rUFLxpO8FJ+DLJDE40WrTRxAOmF9iJKlfJO8GYWIkcU
ZVftQtDN+D4AQVom9zM1kr6fhixhyZEAqaVgOOLKoT4uvHxKSOLXOe6zIey6
3A5SIt52jw7gSR7OnXGXZBspT0QZu5BmoWVb6f+kiPjJ9bhBlFxBxL0xUuGC
3Vni66MSt1FLKnoFSFCBmLVFy2moq3PNEDjRX2gNVcGWTKc09NtAR4M/zazI
fxfGJyQKaDmtwjKTuNABuLhv2otgciZUxZUZQHnnhdxGKB/mddfB00lokoyT
7CgA19BX2787A0VSlisbIJ962eaNHOq2141y7nGiTDcD7oppWSKIyhmSHgdj
DH92sdbaOR/CYI6OqOLy4tFnllHSpQ1DqUga/tuCj3FWYjVqvm9cJbSeNFDv
Y3xH6eUMGIUC8/l8sthXob+OgqXHriHu3wMORsGW1aFMB3eca/X4x8pCIvqA
eErqLGgS7L7CMhteZ2a1rpU4j3uIQRJuiQUZgVMqRrWLb8HAar+/fsM+rlmG
ylAO9wDuFeDxa3p+PoJy23xCh/yWpfPkQPm+5AsMwkKOhoEw1C921vf6+gtp
jVR70bWZaKdP9xIZTmZJvf2j4B4WU6eRxhVBjWU9CMvz53ZaAIQ5dLobTOXD
AZr8swj7g2/hb276WisThckJ5KhROHIcG5/0SiYMYZi69R5xKm/2i7/MLmlm
vhBgbiwn3QrIrxYHgKod4qMgf+unCwwfs9s3MgJV7gU4YAScdQEYCOc7suQ4
kzEfofssqcd2j5FywksQVtmVCnKBDpj98a+VA5bBnYsLcPjBUwnZ3LqfdIiO
owOBcj5mGaeajJ5jzHXBs0fV+P7S9gXGBydY4Mb+nDarRUAH1o8h3vO7Svvj
OVTuVL5tucP4GhwNhnF/3hROQPqRFWfbuTftFPaeomtgyj8vJYIo4mHSj/Ql
cLJskFVPXGN2LSV2jj1lg6sJXbUWV90usJi+COid9yjY84RPFnMn3gUzLL0A
VcUIMQp1Eri+Btk9QXtX//ode23K0d1HhkbLiP6S38B0y6cSowJVW0w+542Q
bLARqHyNSmJ9d5EDMEmfcCcxaNZM+uocvQsLbuus7FTGkabA7DvYL51iiL/1
DSGjxcggaORU5s2Hzh1s0ENhbk2K/CCR7lmQeqEPoSGjtjTE1EFQi3VyJxuI
zWSiMj3KvVS7nj/A1gbbyelFSKyERHv7alEUZQ6dn+HbADGU4CgxALnEyU3J
jJGEAdo/BU+dyea52QIg5Xx9xejSX1qaeLMlLvrLaCu4KGAdQWD/77t9yt6c
wHNQ5DoGSLPtWe6WDiyXtDejVsRIw3TqNgQsW0c4qB2ywxllyAVuNypnTd0i
myhaudMNopKoZlg7h+RbPNIyd1Eca+mkMUqunOJU6NyEBRCdJOfDx3hmW3tu
4YmaQTv5VS0VIboki2IFoczQIzw/2Gd7yXMlLxozDrFcHFeKXUHiEvEkUgm8
qOIWw8WTK7F6KDIAXRH+uAIec00ebX2hZP8X/071aj9BWdV0eq+5XCVC4M1x
hc7y6F0QKBqwJ+6y597Qq36IGH4qUyBXqrLoJVk3VmBNHzDOfggFraYzr2k2
qMO1FoEl9FsKQBRTEj02f697B0TZX0MjBP1d9dnmbWCaoR2ZN58c6PKAQdvS
sE3xiuUZfEGVa3EBSLcJrKhLY9QR2o3AWcWccr7RNFp4HFAdHjnIAcCJvl0w
gkQzRbqlSSxNCK0sUHLuQQRtUwHDesfbTZmhnNt3/zw4G7CumovTsRmw2RG0
KTO7IP2H1GbljgKGt3QQcGgoqPjRr8CoGGYms+86IHUTHEYid01mfNAyTuIk
IdmoXrJvvWt90H6LrHANIkEXuTNq7UQLjRUGczHBeQkDpmt2vHHLAKKjt8NQ
bOYvMupqjHL41upVU1tDlaqYLfritaxdfAtr1ps9DyKPtLF81liqmVPoF6R/
jUf5aPQkPeCo+QmHqCsHY/EjwJxkQ8C6B8NoFbpheatjYcBug2ksVtcezdYK
T9uYf956R3EnajEUZVXVAta9Bbcdvxa5u+6FVhAHO1iE/v0SGTo9iHoCzZgM
ilDNE62oeEDvgh1kxEkFlilqHMCyCl7NAXiwBAu+JG9owNibDgGbPZBx8935
GjMk6GNO4YAVb7esVjFlGfU+DV9ytoi2DDxSCHL/5v6368WV0E4/fdIv1fF3
mVB3jqERVe/vaJKb0M3Jo4Y5hvOHKXJ10zZ61Audy7xQKFtgcY3DdSKI2Vzo
GZllnOLN6m84ncskvjvhD9xZ12sfrOhJpbUptPsSsQ2sy948G1rsWfkq587i
6UIc2n6IhrW38TzjdYZAuGUTEe157djNQxd00g1iJUu7g9AuY6rQtDHOvks9
7AanSPeMygqBFCxzT9dk7UUP+qLC3x42Xh/t/Yfu3Bli9ZzOHRJlDbAo7JfR
/jAzwBTID/ng+zuayrw4LU3RF0P42K8MljSllxIUFjjWW6lBVBWegajiyS/J
R4VaSYP6xxwK7FoFx9PNLCP0Y7b+gKebV7zD4KjNFXR0BVkp8vH0zcj6R8LO
QlyI7KEpMj1TcuInS3ni5RNZDunhSEWPTNXvuesxyzy5OymvCpCK3dUMvs3b
5EXdAMpW0IuonGHrv/m96punDkcjaao8MFlQrReT7yVu67kg7AvVeqHz9bsT
fxOX1i+R4M+DCqVrfrB1A4eNM4cmSeqwvtIcH7jsZLFTvwh9UkiqUbH+GpGR
2anFEd1ZxnRLmhXGYusUvaTvRH6C1DTF2+nJhIM7v/JEnOER+ZYaSJNetL1w
BeVGzvtN7wCgG3YojAiIb1c0IvsacP9WTVCJqRWb1dgoT3JO4xEBLAweL4mx
YKD0eGJ6cKhPnY8i/KcEfHW6Z8P9r418vnl5dFHD47Mc5PrbbbQbv+Z3x2pH
1aAoIj8BWC3b8vQUxu2SEDDZ78HRFMDzYunjXKfFFeA4sdLFbqz/9xQGWHC7
jGOeNCIO5fbTlVPHgNITBm6Dx3ggVWhyaiWdLqGr6S8tIuI4/IDisnom/qwE
u5TZS5dUa83LcBiONA8tmcDzuc2WvOdTYWu1jo/fncUu5GGMx2AKldECC/tY
YMUZ2Ynux65O3p4SizlblfiY0QBix928Tl6O6Vi4+prXU6ZhAGSa/BrzEGqD
t2IhIebFO7ufCvD9sAHvPKPBkcAJ2BETFM4iiIrO7zN1BP87VTaukMeN5FXt
e9jZ2lUypPhdObMwAvjP8wQBUsVyOZd3/C3EvHK0YwPH6o/YOUHtacLJaN7j
Q1WaAhIfIweWKCHpg0d610hzA1Sb8dgvJxfkCfFFckw5bvn7RRd8/2ozAaeD
/DV4y16kZQSAVcQTgpZ+2Q8HU1GxyLSeAZjpDHYGgZrdchdvZB0Nm5xYM73b
lszrsm3IPCrv9bfhAK3UYSr30Xwt4xsICheERYSvmPzjNEBpIiwWsXnffxUV
Ze3pFyOCAkHf2TNjjrRneQMgCiOcjRs75rA9n+gWR+FB9RZ7p/HAGbd3BA1A
mrtz0372b7osuvAsuyeSd10DzQgHWEGJ8BFttAZcaZ5QW0I1MFSZ6AsPRrlV
lNgtEK4D+wOk1n3XnJB5qjd/F+IRTZpbGO/WkqudU3Qm5TIhdm03+OZ/dMVu
2bmDdNKMjW8iIhRVqKCPfTardlOdtjuxDl7Rk7abG27AkrNS/RbW6fZoAvyX
1dnFsoMygu/i5skpA6SiXYH2HdWGr6VjUIqN3+OCw0ngGA5u6XvKQYLkIiC9
OLX5pEOPoJMTq9IyseKnhycyKEaZsaFPnHqifqbBwyj4MBhY922TFMKeEKBE
iuxHcwFW0fnRoTpgxbsDEOnl5EGQCYdafvLFG+FPbqR/p1Y0DQBXFkJ1tZgE
8c/0WyS0co1cmT8ntBNcKtzjAWsLQPUsppy7CvIfqd11yKPFq4+7mIVsEvDS
TQQq0gycvGOQhHF7UAuzY+pGZzOEHRaE3OLdP0wnUS7iiy+hN2Efvs5cVCOn
9UTVnDvctpDfigboKy1OqI9mq5d5LSx1a5+ZdMRdhq3hLpYPt8vUrf7zGCdk
P76yfWu+v5lhjqtRNLjmZqmBFUyu0oIPBMQo9xe5nNyUTA5WgY/0uOndDCmW
K9f8/z7pCZXsxD+eNASyNv5INQOIntfyaF0177ZeJ4MvNkN6zbKZWZvAzeOT
gr5SBTAY+keEoLunKtOge6nK9QuUMOBCPXT29bDnkOvuoIFEbSdGnrdF6b0G
cRG+ldw6EjyHvgUEnlUQHBYjtdla/Lbmbj2wwm4NpQPKSyYZ8CKJkP11JYYK
gjBBKzcztbc/UR4GnSD/AfMch11fphe+VQkHZBv9xDGAZA840ttGX0IEfHCZ
t92u0VHuOBo79v8vovgIuM7AWwlgfd630GFLIYScdErtHuerRy+/T5hf2SAU
2jiEvoXqDLvfMpKGMtJCc+tuW2K2qZFFNMYyx2fDWx0Bi3APXDj/+L5PckW+
kgGDXF4VB1spCX1KYMxlTJcJuh5PdmZUfM4jvx+KpWS54cI78RI7HYy+LEXo
QyjxX2oN0gjC3x0L5y58tewWtAhm7pYADNxdNpl8wWwY9dRWZeJmLHMrg2dG
2Duv6LEI8dtRavFF4VOJ0yXxARnE3Lahh2Fq5WPfeGJPkzx2oey9cPcQIOws
a7GfyQp6UJ9Wv7ovhWNCDCyNXAr3k6fV+2pFc9OhAM1nS9FBLYBieDJWJYt0
wwdQePnR3X4BrHLUVtgVqDT5h5O0939IQJZJ4WRz3pNOOymRdEfZmtgh3LU1
Lkh4otB5rXPH0eTMimKwcHKddFsRKtjQeQBGN0RZUgYmjkeVAQvzZZXe7daV
NVdArjV7KDdLKY0Hjp4wONApQ2c6Ok2XzBDhn3yu4k+xQMyNLhZXrcVV1eQM
M37npMJRoIDSy8RXx8LcwtfWfC/LE97nJWAY6/2DF0LJxrauNHcM6EHVW3rc
VzbHGyUYQisd/+Knv5Eiv5l3NLVp3dpGxDOcg2KAQqB33G7JdBSLxQ+j3teD
7QcJZNbK2VY/0dvAHpRoq3iihNivEB0FJDou4F3q6Z9U2TTyQela2/Uwhhr2
ibGFzL7Dn4t9ezxPW6rFvkouwN9Qhfjeepg/52dT+xfLq49L5m6bX1kkNocp
HF9xtj4BodEmvC4nub68l9HuZg8la5KjpL/zyJH1iCB/uhiTWfgGTeuvg5sl
uL24TKefreL60D1oib7OMRWXQc+lbHUugPZKV2ihyVZM1jSMIe9Yz+9hrvQO
sdIv10ooCaIG/VJNKB4aDUSUM9TW6/BMKC6cnGsI5xX4cAliJLaN2PJjxjv4
tDR0H2XCZpa35QQ4HYs0UhlMpdPlkfE9CX7V3Xy9+npYiE5RKRF+oj/iLRRV
o9ZwNyj2MDU0rgk3hjE1T3vxRBvcCgMKeQuezCM67x/YBlHltIeBVm9ikCc7
Vtru5droHJ5EkhKQPQ+iCxN9nNTUfweYuzdUBvYcTb/dV1bE5Am2ELvhrx0y
oHH/tEOprxtHD8xQsKV69+SnhGPny0lRZ8GWFvFNSHhMRprW3SQnwo4g2dTq
mn6yvTOZoCLOA3rUZ3ockFuWussWm80JSMocOcKxdctzb+cH4ZvAmFyIcdlA
3UezbqPysqjVJh7vCaTihSiR33hHGr/VwP2/J8TqcvQ3peuIpvvQ3VSfyVJ/
0rLemP++25Lzb40nr9FGvi94k0BW879coR5n5TOAWw2RaAuM0yAG72CcGXph
6ZvqH8vYxk38U5iB5uW8n6gIFfCGXhaA2iCmzUwXMJZKmIlz7I9EWzHdFWw5
Igl1Ze7gQPePGkp2B0JHIpoAwkzyctul5Lufald87lEFKXOICePipR9rppx8
C1R5KREUgd1f4rpynE2Jb8G4qcGHhzoOyZe3565cPZyRjSyk4olbKyiAPPgD
iL1OnWv4RmdpPkAOXiFa5sHBw/GQ2CJX78aMSjzqs+J5vfw3HANwECil4YU0
wkm1f6QZY8P74u+5pOnF4Aixwww1WMWCFFf+XiCOG2cMAnIK0JaYQti5x6Ln
Z0166BpaJo4kq6sdBn5nMk77obMqODnQfl8xDYyXv8vDX9RjNJynpjhfDKP1
WtkRqAhPSITCn5P2cvg7VO+ePuP48zhzDz4HWKvCMFW6JIqNRZ5wWHvpKUKL
57byAyYMRNMCRgNizGGWegD4IVjybWriO1X60H5TGJ1SH39i1KG7FdejKG2B
Kz11ds/U0eZGIeYINlzlfNaxMBxB5bWZ2Qc0C8GWw1QvrWUcegI2gccNu6I1
qxBRkg5PHKsC9eHOZ3Su5nqSRzN2LNSgYOkGt3cP1x1Mp3hSgJpkRFwOzgK3
KWG+SSoQvyIUo0ytNKMd+G/O8iNq6YYsHGI2Gm6zlL/bTLOJMWlirQTrQ8uP
d+aCT4v6anAPfCQLF4/AwV/pJ0/djP/qEGEeGEIGfSc/xxaviFAIRXL6dc7Z
QDIy9uGFEg+rViUqkU2b+mN09DNABEjmTIolEcWSomxCjFL6nPBro1ZHwz4Y
TTuZFZV3OYs4Pa3KKw4YDmDUrnsttHH/kgXqvtWjahIcjGBYYJ/dgVzPfwqu
S7RGFrSnwE1fYeQ1Se/pvn79RRgVCDJVD/Tyz4+M7Im17Fho1Rqx40nbP+nv
FArMlRwAUgxGcriZdaoQXdcFlzSH/mfRyMk44sULhezhkJFMohX6/StI+EhV
QQUm5VUxhVNL0V+X/Dxks7yL6ZAbIoQA07qe/xQFWUdoHiPrnXirHnJuFizP
F1wMVTmqkBQBd7KH6gvyjQRWEmbcs6RrHUOr/SG7/qZrDeevVshHm1HEQGZB
bbgWwjd1Jpq1njY5bgjlovFxbQ594QYk6A3KDZmQirK0sWQJbwWp9chgeVqO
w6xwUpsQA9BsWf/atRacyiOumoxdenQK1E9LosofRoUu0FFSrxwPZC76Ee2w
kDcX3OhiEbO7SnWdJMcdfuBo4JrKt51ueFMwSUef3qWRHs9EdnKDkoOqdJPn
PW//apJ+ESbQiRwRUhSOicrBY663+tWjF2nExIH0W+wU2eBHmTiKSUgYPvKe
uPSZolV0QEUiHPcHeBTrG2EOA6EKuFQQYxKC78NTojkWM6MnK57c1kQ5p1Td
V02Lk0sJZmS3k5iwe2d3ha60AOZwz2nRBF9Tx/cKK4xWR7TVszTV3miMI0HR
VHC9bdoQFl72C00iR5zRk6m7cfLIqaDJ8JrwppRcFGbXVywaZvUquwfohJAr
e2b1z3KqUIXy8VIrQKurvhJ3F1i6GlXDl6yfXoth6YxEKrdVn7m8aBLF8AT0
RY0HoTYgB8TbvY9Vl2KdzNUblEb8ztF58W7bR/rkEMsSM4JO5ewA0B1/2jdc
dmYwaN6t7aatGQ2BfUXpQeuUU06IJFVuwcNiQsYRxwcMI0K8YtdhGYLJAMqt
wL7Ni2zz5oCuvsZLMG4mmcwcajilD1Yk8Ld7hmLr22xoySHPQ54rph2RPsXi
T2OEnRI+csyDH0kZfsKDKqGF0O123+7TgZN9N6d6uQZBmxVgVWVPZC2quoq8
lApWSoOH3Mbef/1ncPfoBSZ43Rm1GNdIUN7YI+fa6BKpCZmkCTDgt2z+s4Kr
XSifg18A4IwfN7CJSbW3A8FhT46VmRZN5pK7KO7CdvLCbIyPQIXksGqIEBoN
wZvvSjN0fwt01gBp0OIr/BBx0E9oqF0r22gaGTIYTjjB6MTxtS+KMxFsKlBC
yAbvbj8dLVsqhZBw7pDcIHhFU6///LjHRmblq6+9qXlrxuh9G0aWzd5Ha9LU
0ZYbm/GH1EYuDYXw2h9J7addrpwkOY998+aPdBPLDbwRO28iKoeAAjfJY/ih
EhvvT9UFxibHTkKzrcTe8KWTEOhHpkDYLXu+d2SGi5kpsyfgEOrs7zMWdYMb
n8NzT28rPwAuf8uSW5KAUB9EaA/NtU1nEr/KPLgFtyLRhLFbDNXIl1w2GFdE
/m6pS3cCbWXpqG+4x7IM5W2Jw4/T7erqkB1y0EPzLkBuamQuJHE7I+e0oGqj
A1JijCCpcrsa3ttP62aMYogCZBte8FuS9eE/uNr4svzGGFEf7TLZhSUmFZMB
DXBtGmU2o/Wu/L+PDTBg6XmkdBlzY81gppGkg5jOnt4eYj6yXa/FFRcVr4uB
glnigcB4GvIDxy8KhcMeYgHAg/V+u0FHAy4fod9m+Hy5fP7TPIqUXT35N7+x
tzKubK0BPUcgqq/knDbqBsWfA3222gaztMxU0KHdB5QDzEbOgCMouJ++zqUs
Z9f6ZQQ1SSQ6ivtmBE33bhzIRyuPwnh+gwodILumRMP2VGJPWb1FWAzXgLBq
05DKJrtFQhr9VJfMyppyXIr8K+xXJ/1fumAvbwfcspbui6M2oRncz1N5dBrf
7fSeqcIRH4ZDes3Q8mkm5/FP1/E+zJvnkBUhKgha+9j7eFQYM82WhacP7Cjt
8KCh4Guc/mhs6C0G5FZoMxQoNDqLjk/ybWNrZyoAHArSE5hq/p9LPDZ3EWA7
j7uQDbKMkFnXvGea0BD7+BJ+FsZGi8EAG3WaGfbAd1Ou3av0dWKBeScReReX
vUXTVfAlewmM+DdhxVIOcI6ElCYRTgx7vxS8YBHwpi09h0ov+RGmefgtE+R1
Cbjx3FJdqcL4dGpIJLlfaXDLe9m/SLBbwnVNHj34g2URmrIkHdM6TXQrJBQy
5jqvBnL86oGb0aQtkcqEP91cSrHlzqS7XU+9BFXIU12JgleN9xnFz46ie0qO
+kQW1EPnyS13TGqwMhELiCEwuWEW7EuqxWaJm+DGn3ylXb1LG2nQVkEKzX+Y
6doBSkmHMhkqprhpjgHhOkY5w6iZm4sogDItCwj2ZXxGlriXLVk1X1bjpfU7
s4nasa+leCcQmyt1tuYHcQgipvTfUxvVT6muDJ4l5pituWqMlakaReUuyi6L
EqFbTSB/e0XbHXWF4Ip5gE/fVX94Z0eYjQ1xOrtV77brcuaFlSwe2Wyq5gvO
CkJCjf7QxSZFzkey5wQQ9G9NPkBacEb8yyS0M/o1bCt2kNVGPKx3jjKsvRrz
JiQxyYAlNKJq82ZpjXb1vSeHDABxD8Zmfrw1k0iXLSx7Wyva//+fXVgvjuzb
yyCOZWOm9WUK97jMabKlAd770zDbTdsSe2KJl8ZedrpMpWNZ85NHPtRkZZTo
E/PPX/dPStZe8tEzZtDz33CG5jt7KSfN9Kai/DLNjk72sVrlFKkiavPAr00L
xKTguiPuq/seZ/qxVRC6McIr/7NsMvX5i2i7sH+Q5EHG570bp8WSOZUaRBDb
/Y9Fv05OGEWZOMU/FMuxtyeqoZ//x36F5ZxgodLw0vpKRkycPmXxis4p83Dv
ursVrC1lyrrHDqdtnBckkLfyY07a6dh/OxetygUCT9nF7DwpmTxBTnZ9/KGg
YkldYTKqYDI3QKFd2pRIKKZJH8y2a0oYjk6Jcol48E86pk7M/Y7yFcbZJ7Ru
nGuj/SOQjuudWjdLjDYBGT1evWEkiDq/2oVTRRbbt1AcfIjMjB3hbf0OKCeh
pY8scFctyqb2PXtxRp1KaYsaJQG82hp2Kzp3fCU9yhvKKmwWtSQDM9qgx/3J
p7ChU8ely1CyOshmitw2x4AKjGX2PHJeqqxPr7WBlnvDhpS92BzHkqDygsS1
bHTePdadm/gyMhoi6VG86lF1JgbEpzoA21D7mh71Wb++vPNZS8+dRqPyjeUk
3Xny1PV0KWN2lFto2wWJ2Vg71y5v5qpmxnCGKpuslwYaEz2JA9GBh4TggPS7
5BXN2Oe6UUDZ1UVm7aO+ukxLWYMv+alZOgIIA8EDOnHqNmMLt5OkeXl2BoCb
kLGEnERIgX1Wxzfbl1eC2HK2GewbUPNGEuZjGg3XLwWGEjjRzrugdFqYAgT7
ZiKbAfQFGrzCXno/2m3wPnria72GDDpHCajuZE/Apx0JdJKKpflgZe+rb2Xw
hkCuf3ZcMlwkFVMvkHs4NmuzHp88dX11u+QYPb4PGqp1oVYClfrsLiui5bGV
5BGKzgT3smU41JbP8/XP7Kk9JV3+BGAp0vqcCVlP72yPCuL8IH2jdeRmTokL
ny2eBTFtRHJ8LNwPCjzDyaYiSMKsKQqZ7dwVyjWbH57Lf6BVGk0PsAplGs8k
KywyLoryezf3voGQ8Wzn+j6Fn3AyCE9cZwMANSLjIv5YWIPinzZZcMd60pcj
/ukyosmmjKR0eevaiYscC1yFH/3NzESkzW/4mSW7Fr7V3HU3G8a6SN3K35yk
k3hdm+fMtmiq5f1cW0rJ04A8JRGj6VyZIxwxDvMJ/Ht8QR0Tezz4xPL2fzhR
K5MKH0H5HOjw1+h2wm+p8AFUFTB/HbDVHZRIIn2IS/VC+7e6RFWpi1OiCmRu
OSvye1eGI/mdKmWlCbk+CZAvtEVFuSYr95dl7UIn/1oUfJYOKPopYcqNlEc4
o1xakVYLppgCQVY/FV1dWF+3jqJCrJtC4835BNco1EEcmln7NY4UTnFxXvTT
IEwXTkIk7ZcwxOsz2AQ4QWZeIgGKkEvPVaSdB/DmPUophMjAZ6LJy+mpRHM+
36SWf2MlbQ3EWYYeaQe2MKN0JRd88LfjISmMdXv1r1mz93bnjrZh2wbrYwXq
yKxMsXkZ0x8bgjL2a3pukEpH6Fcgy+ZP7S7mz7G1Yf7AEA+LdJBde+CRcNPU
MkxSW9feMz5fYvpzyZo1zeycHdm21PpGuGcK5cm+0PeE+mUKskuPGAzSTIvh
7vWUf5hVWQHTTXZBfrcWOU+DbARCFCyVle1vFtuV8CYkh4pI0L4n+y8BXRJs
hC0QLcFu04qUJcYUTPuZJi1Lz+FXma6MNLRCC4rLDaWNhOPMyKWoYFo2x+5x
2xHFay20V9rBh+CPPvfrimzASHxP4hZCQfkzM++dlTdLwUlP/xfFa1DlCZTP
d9jDDwD9uG3tPqeiY6eZhguSsGJucWgffmm8tu0fFDDnasrLOOYGgImi4cgj
mNMfJlSiLzvLADn8TI6KEEMdGW7PO/fAq5M8IC29AVAPIPLK+yAl1b6WLO5+
zYFQELYNk+hfFL96AQaXwYh+HRfQ1vGTgCoyTXnSIY2iwJnM5AOlK0wC/ku5
iVYZSF0PjBwhA3K76Xzl+Zi5bgB8KmM2bIODTWVQExhMk5rFs/a7kyIXQyiO
iiuC9l5oG0mydjjeEvAx4nxXIbDQgetattrm5YkZ9Y27xC2c6tYVzewYz18m
utOBOJrfJORkGF6op5xw+K1wE9Xs7jybt5RyRF+jTdIn0y44zaDGJD0LmZ1n
UI9dYjVvX6eS6e4ALqoBaI4+etU9r0Uq0jCfinYXb7xvUCsgRMiXnZ8UUE+b
FT9uUrpvRTMJeWZIRagnTb0IpCX7ZOxZcQSrOC83JhpU+/LtoC/tDQzig0Uf
WsHj++YCRwYZ3Eut0uia6Fq2gN5cXcl/S7DqLuCxnS4K1Yx1TQqkFZWyHVnf
NZzXqEccnMMNjJE7mCXi5Y0PSj26lXp3TnXjQsqSI92CyGdLbFg5x6B+6O2X
DZFfw+Gqg3YOBv98/PXqQJBba3cfVuwn1+bFvxx2yU4Rp1YrQMN/1vkqae9K
JbdF2yiQZVdZ1OeNnfXd9yXMh5fXWZOD4q6aiTGhqeUu6OoohLlTR9+Fy6mP
gJ64yk9r5+45IAkJK80dzKLHwR2NfW55jzs1BYowYiY1lvwfuFItlGYLde2A
pbPsdtsxcttLNmkdSVcQSXjP2fux6qYYAdP8KZwrO5W/VNNVpNLDOjUpbBjA
vaymz4JD00dQZuiKgw5mToGgAM/r2S9FQMsOAxJSMdw0XlVW599kz4PVoeRn
/VzK7y04cNOS5O4Qf+eoIvMWtmb/7hZdLJNOhcZWQmcVeaGHY+Xd+fU3d1Q6
ejELEtLKV04D6GkH/joBoivM32E3jjDhFAOhv/ey1CgGtvdDmYtPMoCtJQjc
Ty5Z/uoAfPia5OB4aP1Hzx4v4Jado9OkXne0xnatneL6RINtz63U45pybffv
foUmjRbqrhw1I+71Dwt23LkGoeOaq/EWrBqW35C8IpPF7gn+LAlv2elUA9tc
xgDUGBC5EaEY0K9DhbUqPrrADzk5sIOIf240dfuwpHrpQ6P+GdJyGTmS75e0
xZmg1UJpCyEstxiS9ybcuc3YEiE3wZsyglx2TTS1iLHzsFomfoAt/l7+V43D
ernve0rZMog55N9BUqKDZjjwcDRMWxX8nrmCTiHYMsFlfEf0CbLG44b7Ue8k
w9KvmEhWietYMgJx5wd5myahty9klw78v3fgp6wWO5e/4EMD1qItyaNRW9kh
XHSKpP0yaCeJw4g6cbu5y48jPM4IDL56nVY51dTTqx+ecPEaN6xb/0/Y4TgO
o9RELpCV3vvDeVL+lBE707/nf3/FwSojvzVqGJx9dnx/u9Gb3AiRnzPrA1ZF
TH3gxb/EPhUS84vk81ArPCKSq3/j3Odm1L5rpKftr8yFvly5JZGaCl8s75ZA
uEvaytqC9O2wT+tDDZNZV12r4lDmsoQanhIw+iPjCio0N47cWwEn5VaE1PAO
H1kDEMrWo0EOl6XXRIPo9G93mEiF6wZFg5vbEwHyMD3s+WRWmzMMHCRlwGqu
HvrZXgDq/JJiLTZye6HBeqtbnpz78Wk5BTQf0ZDVxc6cce3j4vO5kppX9V8L
9q3trwXhpUvf07h1XA7VnxnZQqsjCQ4HHpfXilIpQ0CBcqI6m4X6jKAv/dSX
LhSsSJMVsprWnK4B5tPt0d+wVg+DP13F0o8cxSKW2qLykFpxVoz9vWXzhcLf
R7YoXHrBvwqllN2KeiS773ocAxv2tBEJY+Af1zjR+bxZ5NCi365eJJzG1+V0
Z+dnpH0dcWI2nJTs2tC23BIRJNDIC4yECREL9K/Itu0acG4HX+QB4uP1117j
d9NFal7pf1cXwbWNoNJFMZfrNrdjUfwyBIl1fOOPubotBF1zyHbiIIqCC8AT
cIZnXo9KCdLlUNRk16dgL3F6ToIy8APOhQXI8OPIvYe27ky6thk0a2Ota2Li
ZI9AaNzUGIoy9WNNtlDnQek71nyF49X2Z9zLl4x8OVtW12MLps+p3e+DtaDW
FJIe0awNMBKAP5qemADEXI4eilmAlhXktzDJtstKIAhsdBROal8LNCTrPJ3W
UfFBQczM8tOiUMDscKraL8qboiszQa39/IdyJa/MOBfq8zrKiVoZc2OQbGaU
WCWgNOwELqD5CYNjEQAEAl6nxx+paOjuPBvzAIEHUHjcHxE1Ux1P7SqcWQOj
bgpVkizMDi1c851r6uu9uMIvY/0Sq7SN4id0VDhHeRaWH6d9JDOcmHYE8+m6
gIRTCj5rG+H08K1ddWr/wlHUM7G/jxGmf+EuMP0kmmzFZF1qG79u22OBN6VS
ENOsFPTcowb8GR/DKNTXEHjmoeI8qvqZfUiFQWTtRulKY60uA3MprzX/YQ5b
IFouJKJOPH3UNtIvDt8zZXlVFSU24pLyrwpcU61Kb6QJKZHWKEEBFnnM/l7e
UsnB1W/LYqWrYssO+AfU6tNtOHsoiHOo+WteQ+nUN0ounohgCOUT1+Iq7wwU
cO3COELbdzQv29kbn8G6wJHkqf2oTVPGttAju4JTVodyQZnMver/r2sUidjT
RQrnUhr+ZnK5tFpIpm8AVdk7XGfW/ITC8LIhuNGDfvyhPgqwecDDNuo+an37
UTg/cMNXEUJe1zN8eYVOMyd3daaUArxfs3BCVXk+adjHDCCnkwWzXfm8RNcD
Ah2zE5JzXK6U7WtFfq9D/KxntDgguGx8NpgBPhPfFX2TMmUU23nz2nrD5ib9
l8ePEfJwhphJ0SBf5TvhPhnaqNo7dSE7L2vX+x0fXPtqJP/zm3KHUKv5HUZ3
YZNGaOYKjEGgsMDy7UtcA0mHR0UODHCimpxSqkLjmnwMpApmNz1LcuB3SeBe
WbOX5Ed6evrG+WPRYQGOEkB7fLOrK5EozPVLvqmh0WYj9lPKt0OkI8wKUA9e
XK9TADFJGXO23YdpQ3Ex+XKcb2R8Ps9RBbLZUTz6qug1Y1j9RQg+ljueG8BF
1mC6xdGvFM24j9lvC34DQf1wVWeLpLoIfsKespaYXWoOeNKz6XVQyehVT3gS
nocpho10tk+/gm+y/PHjLenJjKWb3bs8zJCVap4QXx8FlMoj7NiaeXksT2Wi
CbXFnIEUIsrjTKURyArAzKUbImsS9lfMnlziR5V3QFkrtQ/48e7tddjI+TP+
Y58h6cMevvKZ0efxbOR5BXOfk31he1ABOuIIcJZOHO/o+/Y0u0DHrmit5ClW
me0dWHZvZLqqPAmaBO5E4edxNhHCmGi9vxVkx2olbYFWcqC1VHqw+0cfMC3b
9wUWLMOYfSVrCDnigp40hPnLAEsZS3fJWin0cksseu5cCwtmxYXnirjFuG17
LmHfDZVWyjCLPgXsmUcTAN6RFXAyVbVZgkn+95i50YEMmiX3igpPqJJeFzUr
KD+dRJU+L97Kr3J3sJG1y/GxhPcqXBuVMWiuMhvwfKILWh3emynpCW/guatP
ArG+Ytnb6W3El5JOejNjmlxrrAQpvnZlyzJDnnyR1Wa/wNTwbKwjmvHmPs3P
VM/Pa0K2VVCQIgExV3A/tmeOqDdjdPJLdRTC+YMeHXlNJTsKDpvFgeWhALRL
1hcan6V8y7/q3OilWqZXpxOW/+nBnWu0vXfG8ZeA69NmIVMrBghtrw2AqoFi
bU0P3NGEkDhLJMUyjuQ/nEqJDTsOBHA7jnegBPIlzJuyf0mDDoedP3mLSiEu
EGhAPcgA+387Vo9AFksHLEh05u4JTKiAEQ5APg6wN0eLibRpsbsIVB0SKLIq
bpFo8f1dwSk9+9dn+RqBF0bFT8MyYc5qXO/9lvXjBKJ83WwlkK/E4Gr0SVbx
lV2IpVkZNfr0iP+LNcEprtnWUXyWBQfJgpsHAayUvKu4emMajAUdPTO7WfPa
ES/blwGbuJEmAUMGJ/QhK+G4p/WvM/IaOqx13nAxpQOLycEcMFZsEgSs20ZM
aizuAYN1BlC9OwCAPBd/1GwEv8HEOJIy3q4qiSk5i8o2yUCqF7kmt2tGLfxi
b1ZjbgFJatrrG65Qu65r9M9VWe4lsOVTp1wMq/IVWHl5E6Drod298YaA4kmC
BR5ZrQQfQAlsqncUytrK7epN/k1VL/I2i75wBdTzoRNHwGn8a/MQmpFDV3/J
txtwuWVs1QcCAR3GaAKYd7ASABMfYCp8Ti/UfAG7n/bOocT9V14qauJeuCP1
jOGnr7fliWBt8T3FwshizaJtrRe023ixxTQ+cz8MKr83M5vCI5h4neZB60Z5
/RO91vEIQqXNPcqHvn3FlZx7TCN8WaNE90uvlopDlXWGujnx7RCr6Mb7Cp2C
zHTA5kzGg3yrUejkO3+P+hilSzlwa7TlpZjyp5JV3GbOkJTDtA4uo8AYb4YL
Z3P2KT313ES3rid5q6OseuRph+iV6lkdFfF3BVV6KB/lmKJCSTvdWpNLCYDr
b3IQrmdObLMh1iSJzUtjzzC1Vtxn+3uMoP7FTO4uKqO48CQm7J+pC3lFm3ly
p2Q5if43NJIEMJSSTkAbdGku8eZM5JJyOeqOaatXvwE/pygVWe/p8oevAB/Q
o6BReR4gz74CnzLAgttcRlDXPFoYf2MUBdWTG902cWWpVJJv6C8gbvTsPnsZ
rS7MEb0oa5VnfGSYT92Zxh/fZ/GDaYyonlYZm+Mc820N/gGZw7IaEqyA8idF
UNCKtSYZugpqkBsUOjl0TMLn1lI0KeLeaKvkzfJPXr9fvzzSoB64w7/rGrUg
DFXm9lGOymSaZ6BvW+E9DKaoMArRo9QPvu2ssW2NTyiAOX6AT45v/2Dm27lU
wK8TuiJ7rKsgygbnd7c5ePw4Gn0AwDXvAG0Dl0kIUsw3g3tv738+nktN+gPy
aI62C/2MJA1UeEu/EsOsmXo/qOhH3oOe1Ao78MLZmsMTd6w4TphEkh9S51tC
ZycfvzoJnx4P5OGaENo0ZkibcI2dfyH9STlhy3h4jZP3w3Fe/hb6mor0/2nb
RVTxNogOIV8vUmqH6/+aPY2PAjvxdc59hQYgP6u3RVnm13vNpkiX7vbhiNXI
6HV62QhnDw1i3qjPCTqvLVqeyRQqzbbPPSOBylf4YcIc1yHMEXHeG2Ws7nc7
8riY5Zau0Z8BFpnr4V0qX3E2a/M2Py/VgFiXU1Ek+aSA5V3xtKdjiPWWDSUQ
blmsCa6l3bT7b9QiFmsESfQOaYRerpSQcBLOpn4OMjdYele5hvmA8jRMzXKa
f8LQICnkpzhWaFpvchBeiUFoFavlCM7HMgKiTrNs39tZ+shPnDC3Zh6pm0Sh
qX3/2HKcOTJOFpaL5g/3ZpV1gCnxkynIM/kO/qylG2WHbW4HzKuUaJrwxTSW
9TUPXFPtIhGt315BwDAPWQD+QpfPyQ7sYMV1P7VTWLdNyMGPjHuvmmi5oUce
2KzSCeBuVQuQFVZKWRsReGG9rPBDYzTukW25A5JUBN78AJV0/m5lYnxs8X76
RtOOKHNsXKZB3ZGJtjbKCcGkj/xY9ZcrTXQbLbrQYT7SotttuXw+yJ8jPxnw
QO/UwxEdb7OTtyxFmSsNEvLJflDHCwan8uk9WOn0dfyQvfcLRS6WBsGWypm1
s6wggw0qkUs3Fjm8Cy7fMNlKZvSk1XWlosOjeCEsnsBNnYwJKmcmN7v4/oD+
JEUgpp9pEYPToOPP/LB2Ut15pZZ9E0thpiSzF6tmVHxng3aBD43BMm28sPSN
/1fSjPS5a8OsNlD4VOA53F6LSCdlZcC8yTfoDz9qBEcJxYwx/NRLYSPDKi1w
GJfDZ/wZEYPs0Tz+TPGfGXMySalHll9mp9fS7IC1pO53n37GWjrqLNF7qoBw
Hsc1PPjtzRORLllCACdxJQybC9aEUsZ0H67CQadNPdj/nAyvdzGAKj1ZBXML
0lL3RVVsa+Yn3VZtbQZ39mphfoLZSYwcBKlmpTrL3SbxB1bfcke1vYoLU1Vv
bp7/wGnQAu+JHlgCfIMhZj3zLHuCVUDg5pMJ4GKlyfkxcKwCrXxkN1tvD4TG
6xAGg/01erj9D6byoNa/w1MN5GIi2+FJeetx5vMibte71XUck2ZkuBTJxsaP
vH2BknBCc9Hv4/KpLinytoisSfIIkC0A8FAghVCscbFHAdUjcjWQg9Rk3AAt
JIHQBwRs3kehdMSI7jKwwrTMr59yGnYDZA+BBQUo2lHMGHZZktMt1jJmQ6oq
Rrxr6Vx000ol4cDgfxfg9qrOGOFQWwyAXgz0wYmhMPq9zoJgcn+acr4FCeJ3
tdIDjQw3Ca2wQ+XJY0iK+d+rIuq1YQwTKk2uK4dUA3ik0Z4NwUW0Wcsn1j7R
lVAZtMtXAfJmWK1BkjlFO2JhFz+fiOrZzQr77zWYqEnZpFyVz20tQIcWYv4K
d/U7sUImt91Uq1R+rcyOt78WhjplnFEo/qa0bPcvMyQNLcSRrbgTrhqQuP2L
5OPEggZl7icLaIwlSuSyPY9kTmImR3Tqrhj3S4fDpUnygOOaqhu1H2o0nLK7
sLwt4kZ4/audtYMzAlIybsoJawdAItOJOSY1XBsyn4i/grwGposkMPtqWTab
Z0HtiPUqXVwEJstOlYRWMdi8Ixv2nwZNnoVN74NVIJ9bxwbTBVUqcrGUeraR
FFaEJinwS6y9sDG6vD6YKyReq4Q912CW54JCZjcqprKF8zg9zUwaA4crcByl
wsDjVnq54CamQzM9RkUt8VpYc51+uoYEUbslv6X1CZbEG7cNVqqkDqrCPmeB
+zMOgL7uzrVA6NXQikgmKXc1B71WhuEuJRFSq7NccIil0Sp81301ufkQH8WD
X3wrkOkbzrSmXykVi3P3av7G9IZ/FC3vPLZYWQKS+Y/bjMz1ScARpJvTI0wn
HMer5EKOgoX7tx0BIWdmttvjAEVOhPfyK8/u+7rJ7fMOoOCddMW3vHXW/iT7
ww3paCZwIIojuqNkrGPcYqMh/ib51NdvpB6x43gEHBRJ4hIICmt5qTf4Iu6G
HT7+t+51LIvMkwmT6qmc26zKsRMufSX3H99mSQ2zl7n5gidzbYXJs/IciH9L
7py+u69gpTbfHvqSYOurrewzZsYjBt08PPmsZv7xKvfdTB5VQNk7ko3ARcjM
iOeaadvwY2CwWYZ8Y3dWsAsEB2Kk8y81505rc3XdVICPfI3nYLaxRqxKvGpV
+t0OTYIUR8E+9fpU7F+zIJx79LvuEvuSnm9OJwavGk25ofbnushFzrCDYRk3
k/vbiYSeOdASZMFLOf/hsDcjQjR+S0XXSVQ+Z8YrBu/lMsa2e5vwjGawa/DC
c/AOU5Vqv48XYF5j9XadSxGONYsgkzwTEM21S3QO0R2dcLpnJm4jDfME/p+T
Lx8gDqiKeoELQdlw0tpJSL1hxYKf1HMqzbKBalqLVPmyEfzJc15cKsXsTV+y
WId2ueLPX2qAGOKsFCfDz1xGS8M0hVP3gm/OM6H4blcvk6xAsnjSs8JV49nU
IL68x+U01RnBSLzTZ2BDYNsEo+Dg+y6E5jrI+38R+x+IuiGtozX7Wkg+0zz5
I3ka60+oGRxM/9TFW3YiSUXRR2i9B+XHFkzNL69uRxiW2/nj/ZGULLShDYMM
HWliZYRnCs+IxY0TB3c9taBhSFUGDtAkp20llrJ4dHWe7LEFIkQeb++d2rOd
qzqn0AgKKbeLdo3K43y/XDViS+ieCASG48LWlN5pDcwYCfCJI0A/OwjHoQUQ
70iHIJNkdY/qVl1/Ca4hpoMuzjO//y8pR/cJWy+uti/iUiady5u+QUQ+aWkA
K4QeuTHtMsdEnHMwzW9F9I6Iclo9AVbJcNwWCl9PqOxpvBeUE7Kk2Qg9b2Ne
/iOZzUPnvb5gu7nFfQdJ8cR7/pyQND3SKl4rwlXkkBoGOTjCjshiVLDmdpCU
sjAkRBkgJIdLo2ChhjxBrbKDHMQqD4HvRWT0HaQugu+6458dy5zlEiWC/tfY
z543FG/Ynfk0T7HLJDe4IkrVY4JL2icI2qOJ/LSVypdilLWGaXrOWungTDE4
O2UbDafNJ7//g+AYGxgrJkkIgoWMjjkGwpdn3pdfoYFfLCXL6mwvluyytbC5
t5YMehfrz34ebpkkC7tEN+u6cAEkApq5gQkgxRRuGtPHBWRTCPW5iiIFniP6
cPDWigk9AdOLgr7LekKSQIbULS+/ZLeMZXFyxsUE/Wz0mHA5hHnevuHyhCnW
P7hI2QyHa8CulxFJPJq0Gl+Ezzg6D5Xnjz6h9f0p1znTRBUtXjkj+L/oc1o0
XXk+/LeB0IijFrRJ176l9Erjj1ABFPeM8Dm1sGb7ZVw9iwuqzxMZ6mrU17aW
QijpxbpNYLkm+EBpKfAC3GIDvToPmsNQhiGpm9FlKvrqKKwfcC4+h4fMgthT
ue/pfdeioVPj3lcrwnu+wdULzLy/IzQrUEV9/EQv8UtqtGfip3+sSjO7SUQp
QuGq7iUibLs5iqfqGpRUEpUiLV0LSY6Gc9r0aZsRrLEYkKkhB/62xD0if96Y
NPyNqz9xaYWdau3udaiGNq5pAdsWZyK8WDkOQwldjutqXPPZwNoqMEH95FnU
n4jNzO9EAEzpYwns3xGYxE3G4peL1SBZ4SEn0hzYk/6phslVnDeyuU0sAA25
lb5glT8x7xg3nr5YEbub1gSSxIrdkXjJGRWtlM6Oi4y/ei8gRDvpKTk8Je2F
7jINHfGE5Asl/zh4cThav/X1Pvs9wCd/JuG8soeJ0dJ6Inc3VC2A5MB/fwAi
4qFdTsTF83Mh6fF45tPi2qFouxWSi5P42k2OatwXCYxnO78ebrMwCBhKT5Ut
r83LkEh+79fqEt+vbc+Ny+8luuhuew3lZzhVFRee6y9TYw3Xal27yJxnu40a
BoUlt0Yq8saf56kKvXlgylFIaJwr5nZ4CRE2p3KICG/FIpUZlgRG2xWy92XL
SV7mujhQ+0F+IyknYVu2jAtfBU+20hPPg2/WITB5iuLu+Q7lNH1kdIFWNtZX
2YTL/bhXzw450pMQOr1bJ63iWf8OYu1SEKCbjXKRBxuIV++sZ4o6M5Wm4iMQ
Hqs3oB/TwSZ8nUDu9eoqb/0nJ15urUx1VM1jYMWUa9bAcr+oB6TTya5ycvyI
4iTOqliVpbhSy3JdbSXaVrM0XSa7A06zEqVVBB+yA4INrXrHtfbqbW4qHxCR
GEHCvI5zSv7neymoQa1ryT2rbhYNt4C2Ww7STgEFJWgmjAviNpcUiQBxND+F
Vhgmikql8c/OJHkFCk/asMTcE7laWGNLyuvbMRA6DgsxgP4gwaF7w0kBc/ot
Wb3e8PhpAMVJN1HZJ1Tv63o+erxV6ZL+CqwBayfJe7jAHdWeBNzWg7tfv4kg
07ZDIvtXlUMoJ/KWN6yV22DOqmZVd/tC9TKocbexQ9c2zXC4g05xecgD9bLG
N/kOOqrs2cVEOMrzXbQrPjs0vRvYGAFLx++T4T8sttDqC9MHwFJGmaYyHkX6
tuVW5WFV1SWyDJN1fmLZ8sw/wamhkcLtd3lH85IZay3iHhZPf1bvezKfjpWd
frx5+6oFOr6PptvWiTuinsEN0ehetCmuUekvm1hvN0ZhfEUGh3IjZJ7w3i+i
cZwyr/AcgxvcRy+n1E1xNhK8D5xYHOQzsOjSCKjPF+gLZj7kKW3w46P3Q1c2
wjaUM8UhgWQGE6KdN83z/Na4EDBGXFnFd0Hxnp1LXxOwjVI65zOeCRygjG02
/qvkEDrEcBhx7u3271NN+Y3SYP1Q2c2eLqsxbJkz6bZ9vtl0f9CTS+Yv5XXT
uS9bZgZZQDNX+iYMDF2e/y2qewAWlBleQIJjwBWaIoLKS4uUv81mm3ZA8aD5
2C6+MKVxD7gHsYU/5muA+KdFRz0bhPR+I3hsK6D1F/60pEnp65B+8Rk0BaeV
2IohdK1liugRdlOgBb265qeyVx6LEpKSEINkVLbDoMChaRC4cYMWKpkdwr70
9fAwv5GvfZMboCqQI2PtTghcSwvAuKEzn25AXgAIjlsggxVgWkg0egGGqMUu
PEaT6s4ojlzZIHF1Ls4eYtyhMZ5Lf50rMmunApYx3YSswj9FKY8k678GH5ua
w67skNk/YtP+F326QJDVamo80TF8OQtFinFNbJ05N23sIaUbltb2tzIzmJnx
vhOklBm3VR+Tw3rVoM2+xR40rEI9Fb/C6/BEjsCypg1JDbgTZfDo1YqSLBZU
pUFjD4qDM0yhNJnq79Ky7Z85T/AItQi3i97luxOV9E0PwFdnIGkQIdBLl66i
4B9oLKX1gd0oBFg1zq0HWIuFyVfsTbpQmAAdSlm1wSAezyjuPc512Gl8Gkh2
pm6GO0NsCoub96xTYqiP+AJxKRrj1zoYpHKJYZaP8mJSzeu3rXM0EkanrvsL
CLyLMkFPmHRlm/ScqZIXt3kW9a3gYs/D5LWVDw8Z7M2pY88B2h5VzJGSXe6Z
K3MO3Fc2l9GQu851s0dSpzTK0+zKq7G7JN06MY+6jUF2iwa25A3sgZfM53oT
tBaLe2fpzuudTjPojDLPsh+dMBjylMhAaz5UyFEbll+oTFg9NYzeLvTe4Y/n
Bsp0E8VuaXoQCdu1PbHzydH5OQA/SAemJSCX6/UuSbSqp5HzEBs+riyRSNte
S6dlRN3Lk/UZmpzrDdlpNgRhRd2/Z5sQlnT28UveqhgmwE4RLQ1gIULvHrFZ
BC3nn5Ts7Op5lceIBLQQL3zg2TD6XrU0LprNdk1iyfvtCTOeyENfP6JJ+jST
0M+OVPOdbYuz6SYL5g6leD0y2/WlGPNfNG/06H6RAd5TN/PamuzIc3UKbQgw
YvopQLK3cyXuzg4rvR4L5iCuOK0i7CpkpzpQCFi1NXnf5BpnxVzy6KEctGa7
W44ktOVHVAA32lwavY1TXRgzH7BZ5HmA02aUkQ0eLP1RN39R8uNtbHlVl3M7
mqqHE11YdG4yDqG5/aZFZvIOxI9NDKztBlbqV+bBsvBLqLbjqSK9V8NkoJvA
k4iepcMRN9mhQ5RDMBYWRtbv61Kdavun1ZlkK8C/onH2JS8DoXr32v3GY7Nl
vgkLQOV075ONsEQvnmYizv0dGrzsmAw4+DtBKMs6Zp9iULDFPnihf1z9hwsL
xOsyIWqJr7Eboq+VYNIs8gWx+5u8R05qExBXnEEuP48JJMFRGa2quFfVEl1h
h8Dl/PzJaQIkC9lbtCqpWr9GUmfg7vqpj/kLsningWxT+REGqJe5Yol6BUkw
FKaJ5EHtNWR8GvSaRebT003RnB/CvtvCOg/o65Bk+AA1QtDVWUkgaOjUH96l
s1fsUlBPlz8OJ9NYUzdZTqzqx8xb47uX4EfXgbxjKJT9TvNa3USYOlCCifpA
uCE/Tn3iKApvVb2n4avckkcdeMwwW9Ia+t6y9FiJh4aJnd6Gkr2x0RI1U6g5
y9WCuodBmq95oOYCrdEu9OopYVgH7lJ2QhxLpF28nqCdNmSGqCpEjW2zt/Dt
udK1ZIRFfhR/TAYzAqfs4I1USKwH0rjCE0Uu1KvH3ZRPkvxU7fV0pkJ6ZysO
2LEzZPt3N8KI8Z4pdn+/EmjxRado42QpUlR4xG82GWwv1BSbbz1wG6pDoKVC
mbefONkr67MzfRGsR1K8iyjEWwcIudlw9wrv9bUDpuHv0e9MjCrXPhvynW1p
Wj5nJaa8eOFXLCsNkcF8rcSL418fSUYpOkNnJE9a/AB3Sah7T46mHltczI9j
5SNiZRLZBFI7cBfCnuSteL9Hh1A9hJFj83N266iWJFTkpAsthNeUj0Yw1/uL
tY12D/GxBg38+Gky98qNjFrUtw2TvvnuYN09f63uJWmVhH1QSDJNB8Nc5gcB
XPuWkgb5xtncwQBW1PgQ6qWYFPqT1aS75d2C35JNYkL9L/Qw0Ik+DfJ25UG4
5Swr6PwbYRRQI4vDh31SmAlS+CfylFevgDchOc3SjfWFws6OgRsI9RzKZbNg
A7l9+ZObnpOQnvAPjWb9Cn0QA4+wi51R3KzWmocysRHq2sPOTSS1GXC3F5JT
m+OTVVK5sCqQzb5bGiB/c/Dx6b1BhBs9FbDVvGpQ/WuPZPrZPAFvaQw0SmJs
zzqsIeeATPFUugDjWQsvXCqNsLq+3s1+jxtNejGwrZ/5eY2PKyO6jWx9t4ah
LdRmyf3WohMvdrwGmo5d/NhgFUYFX5vBsV8jvSsByZr7ONq/LIuU/94x18LK
gQgJDDsEs/U4O3FC+eU73FQkarFWvhmCdR1njjEsSjLSNhiRSe5k8U0sVrVn
2LYNOGfKg3h5it0QgTgaoM/B+hFxqarhTWkvofPH7rv7vRJC3WQordYc+XDZ
+vmwgH+Tsljt/jcHcX9T07G7BFEypHpu1HWVFLC++PWxn3CfIAUYv1TBdW27
vZlPhC9RWPwwGBsKgnHNlMDCMvWu4HvQYg+tTFWG7/rzHKv6eyD3uaKIlRvs
dp+vomcS20qOxA9Hr8QuHpBTQgmZB+Ew6Ama1z0NhMmiMn9616p8PYFbw8Qp
H/NE2cfEVEN2O8zdMC0ZSwPdqIZ5dl6aAJTzJupKXYT9kACTPYvYTGJ/eXSu
mQTBHSfPhZ2xUW6cW9+KHJ6Yixp+b3TLP7N/0m+DJLK7XWZZITeBk9A9YgO0
PpeSmdf/m1v2wNsKv+X8i8r4tZOShS2d0pXZ8v8s9nr8t931WoPq6OqZGCxf
MolmcsZP1ShSdtdF7bJv5G6sUUtpy5hd8iqlHQdTyxKWKDepCImVeMbli1T3
e6fijYVp/k7uZpsUPWQBU75NLUILpFtMzfmyxygFGk1SR5azB3SvN5k9DSHS
6lkgf5z3Q4GMD5ZvbmsOn+0wFZDgoq4/F7LwmU/jABgmt6qE2jJ6voYqfeqy
9sKecJognmLGoTrFQEGnsCxqQO2Y4fxcYRbtghcGtlB+DnUA+3buPT2QLabV
gcTPz4Qil+ub8KMp5YP5GpVps/e/j2li1AJ0+XAwAfwDKoVKp8/0EJTg9LOo
KcAVhm5zAzKzNvhQaScqXItpT5Sp+aBHmyVbkh3R+K0XmHgch9KzPEjWZl8c
pZQYbnllvkmOVD5vFDtYhJaNv4srDzt6EALnG/24ZinfVhzfsZWarpOa4cnD
PNTovx0V66BwL+9BMIwenSD2zeVdEbRWFV4g+AUieRg7GB7Lf9Od6a7I1tPO
CD3cKfLnAbCnTt+n5atUbGDeMEJw6epIXYPMYALM8xcFrsUipkG219+G4rJc
jv0lPr4UZhcCHDQPBCHFZy+J3nlledTpHi69eP84+Mf3Af0Rwu069JRN25as
JyK/M/le5+CdYSTaabWPyRzVjXh38Ykhfx3iNpZ6dNTcVGRVfdSaCeBSmtKX
Wy2v/qtcWQI2zGnRLqpFi6Mgz/gm9VMvFRRJQOf9Lr/+2Oog7yFKAP0daVZB
qCVUDZ/VvGum8nSDlSXIcIkLipod+4acr4uGvkNumwCrblg2pOcbg4jDwEHQ
YFgLBk7U8EDiOw/yN7CboioZ3Rc/i7lEFWix0canI3RaDcmrqob2R2v9c4rD
5PrMCpkdSNSAzaS1y9NITfRfPdHaMdS/M2nd3+dGkItIg2ht7g89n28WRn0c
HYQgenvj4hyM+4U7Ssgtxgrzkf1CcVWyrFcvX2eYVy9nr02PiDfWUtwt4K22
vc14LI3cwhw6e0v26rpqE76a8ewyzpcre5gp5QoF3pmiSpTCeqoa9TcrqQwk
VWjLLkwaxSG3DuWq4J6pnT8Ajxk8KjXBfkmtJoSLfGjuXf83V09/P7yUrsTB
EmPZzMlhu485ErMO56BRxlqxyjjuCHiFcF+WW2h1B9V4ujrVmdawTqJfsBiq
lknWijQWAFLhfb2qMLzdgy/EentXNtqExf1qmUZA9AFQYNIE+0LoOAopCL09
V8DnX5ANAz+Z6P0ryR1dTOenqeYLRSAbgVAUGafRzFRHKZNjEfmtboJnPpjW
3guWFAipy4FKHqvvt/woIpzivXjvZAMl/KiZa8YIquQ9v9/d0ZoEidFxUsr8
wvekUrWkrqDv3gjPGcFUbr3Hbr0LnBx3Z72cgO/3tOrtF6QFwJKJLkM7tMJ6
5CrCMOIRstlXbBQUg+B7/mrd+yRuidkCBBbAVNiOmRV4YBs8BiMvTNP5x2EN
X9x19LnQShyZF1e6JSeMmYtwrmx9IfvA3viLuM9wZ1rAEXOExtHyTFwIIuLd
X43ZJsPIO5ay2kjHd1/7vaaYwOAPGqVFvLpZIiiO1yfURuhHw6pVCL3zoIbC
HefJXz2v5Z9iYSkViUP9Uk0mQxD2PjoCWPihAKeBoZc/pdo+72TPBmUd8Tt8
Irhh/M/cOo+t+Y39AePNZzzs6m7KilYxEtDo+qakHK9ljg4E2D7hh1VwzK3S
PD7tpOVp1PPwu9MgDzkR5J2NOJerUPTff19MK0sakQQl+RcAi8LhnSEx4Hyt
yQhFsQ+/TWbZuZAsvfZFq5n9XhPNPY+9QgBSNYtF2MRFR37y2+r1ksDNSAVv
PSpivYZjWw7WHvZK9T6GzLZ+MuxMes0Ym5m+N7XxDgmAGxAL1zrSCWLiXU8l
8Y65jzRzK3Hi95O/AXSDR08L2iHZQ9xeQ7jk4lFy2x/k2WyjEs8Z+6YayRCr
nbFMicUev3NBeZN+OOLEmKn2Ug+bxpW/dG3Ya49KrfLzSNaR3NTwRfQzmwGm
BNMbUiYvoRlhNL4yThsvzBDtkD5XFC6FRVyZdf0rIhgkKPmuzD+Suy2lQSnd
cIW6aWgb8rz/nXdyb8kRbgJhXb5bibLrYYe4YRbADGUzdp74Q74f2+dU9wxA
T5WPJK0qFSKmUGt0FlJu2nPY5GbofvWGP8ZwsO55Wjd5uKoB0g/yoVeRihYP
m0VMDH+3TVbEIDRumvi+7V7mszzfMGKmkO377IZKLsQeTlKthzUQKvYrEv0Q
UT78s0VA8zN6p9DplyoFMXK/UkkjcMW1vmtSnygzRT/d1eblDxx4bviRTu0S
OECMBIC3mkbnQFHD+H7zLAwuVJIVSqwvlsn0uTnU5aF9J1QSS1Q9k+wjs6xX
nY0VXxPDJUkLpLTYVI2mDgunwlBKwMN3rL+OmFftesFaB+Z4wYuMw/H32l4+
syUo6ZxW1tUGV3KoyrofeXrzQl5EgwDehvH76tXZWG7212wnNSdXRob/CdE2
DRYkW/qBk/rfuKxMlXNtIYN1EM51WD/wHhzNZHkOuDFkg1ETNVStzRJBC8P9
T13va9QlakMVNKdjCcc7NM4MXi/9W8Ag2fYosKkbAaPe6HMLwquxATX5Zt/z
b5e63svJHQC+UKjQP37sAE3PQVkwS0l7Zvudpp5k2UYZSJXSuYwspLedBNK8
PipYljZPxuoqVrVP6A9foZotrVFtTEiJNm0EuWMH2Gfnc0PlNikghgFj+Fxi
QeiKG7ZoKlOrHm2NAGzkZsltEv8geBIvYFSGVGdhw3C3sFNQhbr8YKROQRzJ
b62+1pqn+cU/YrOVWqQ7RbOHb5lkkBeGIop5uVCx6XomMl/Z+klqLEq8pHgn
BJwMyBAQaAYIUOrYQoUqVJ1O/HS6WSac94aws7Z0f/8J/Hii9Rv6sVtlShJ+
oYLVLKr4IIWPVhGFh9GbkEC8DHtjHVAPfdn2WyMX5PzQ0F5m4DRADrCqepI2
Vok2Euj8UHc81/qvs6+cW6XzksPPJjkhWZAljzfHIJ62HoObR8GxmzDYpuN0
dvI08OrI96uPJAnRvQe0Ei/0B2rN+Rw6yhkvuirSgtbAHQIhBZ09WeCovNsb
mP7ySgiqtgDvJThwEkuG8lztwIgsbKgpVzkfCQd9nKM/cpx8vRcFffs9n6Un
Lad5g0IZlz5GLSOFZcFsZja7q6JKA1/Sp25jI4CY+39RoY3iMD6m5qcCjc1Y
1fXgeyQRlIscdEOe37g7YCtbthKhaXGYveC7Zn6dBNwmLvYFT3jKI2UY5WPL
zPrNZd1+CZ7YtmihtROW833UxciswoYgMRn5/xBP14wK6WJ/D9zQAtxXrIXu
szzRVFDjuH7rAb8pC/TiWfalAWjYOSceo16kbJeK0V3Xky/YbS4Et1/rHSn5
nAnSg7o7D4PhT8bfmFiDx2O4eHV1a/WnAbVvjUGTr4gXPhXykbgeAiN+UVZn
3ijcs8V9+Ah9lfjYYpWalsaeA4ik0zAnkpdKXEY0BKuQC7t9+dPorKilXdlJ
945TgaGk1k+Ei288K+DXYJ98AKz3YUXFuvX5v1HgxHvN9y0E5AC8uwLnZDTi
ulIsLsPZYMN8J5gHeLxBLLibjHOAoA2dK9Qu0UaWhyabvA27KoNizaRVz6yX
R9VT9g+1YHb9pMcFYq94NRCdUW237CmdOeKOlou5SaHDyuQTZ1Pbp9y01Uuv
KqjaInVpmFR889q3jTs6BHgB/xZp3iG7BySmZ87QaG++0M9hcGZfHSBWfFab
BcUsf8tD1A80vHNGFDUHSmw71V+AWLzCBLAq/FfNipl2K5ELl2/gjIOCaB83
C2/Ok9B91DoUxMg3/TbNB0ecviJLVgd++ozAK+W2jbpgmgiCct6VrSBFhXX/
CxkzYzCmFGtuq1i/65xMHX9xGsWO7CpcfdUNu5eYVBwu+6VK/wx/UYWy6aU7
a6U69m60rn2iXNeIcD9DsPw9oHpV0UAdlsvEhsIoMtayhhOjrCKBdKXQdETD
+Xd4n9XXchVdNO778IvlZBQtB/iFe9AgsmbgqIncd5FMA7LGUUjz0XquMXPd
evJOAHWkFTwtEK4sQRhOS5XP4FsIzrWKYTo5TWNxGLj3F2oSAG79194aQYJG
XxPldrbWqr+mpfDfsrSioCgzIBU2GeD9zzqoeOnD6jLK/srdUeycXVFXIjdz
yZpucqRlfUP3QsEI9QqjBoI3aAHMbExzlwtx+dGUj94GXNE7qExNE6vRJQ0P
ZjhH5OXZpCsFw0z35lzuOLpNPZScWq0zZH/rtN/oKwY5s3p2iJXNyqL0KEG0
+bUQR8LvsqfdEZK7PJrFR0Ft/c52L8OPm+t5b9+eMQHT39JXssVVSNLy/Z17
S+4oSjJNoWxzRdPYJmie4XUSwe4//qgWBOh6InSG1aPMve7qqNl9hDzQJdvP
RHmgm2jyu5RYwL9sjo6FUcER4XXkuAetcbwZsjrHlvkFH4XlCuBRJF3ehhZX
nT9oMSIBKmDRZAXDz2cMMvQK5vGvVY8FHg+MMit6hSqFE8GI70PChttrFeVM
IsmOWItoak6IYwdcSpP/DwM569VT66wVBz5BNTQyU2BGxHKT2uKu9De7PWYp
D9HehkpzAcBwnPwwSNQBX7zmw9anUkRBvYhZv922ydXL+fEbZEN93mt8PxRX
NElnZXAb2w0SMCN+SxXtjLwWU4ZgFCt3WdtO3A/BIkBz/eJfEZP7P3lUehYT
VyVVPMlLpd9m2TMjpQN2ZgiqJPDMJTmhL6vKRImDm5dwjVDexRLJi1rmi7LY
cENjFWC5JK+ZRnpovqUjehN7WHrpGTPey4/xWNipUeah4tVub47y+SUtSZUt
ricxoFsX/iYrdXI31HEICXVOXwPggjwVCPoR8W/bh5AOoyylfOTQB4yg7O0y
3Z69ckST9PqJM+OGxyWUPPgdNKrBUFJAhQynNfRGYIMkV9Iekx9G+Q1NZrb5
lBjrrH4T9R9nGanQ8DZesFiOd4gh0mkyH9x41ASUMEQJsdcELvjKJw5HOvUr
+veu1GHxgEi6VjRctRBBcCUXRbMLGoVbQRhi4BxbC0feqN2UbKnutHQWoLoe
LuDXuQtM379xDLyiqDB+BJ/I/9qBsExvdSLi6LdibTH4u0ajGB9ucaHtd7sh
jGk/1bQEqK5390UmUCiQ2g9T1NNVXi1ioajW/GV4pSQFikk2JlnujMdzqJWD
6dzNT4Z3RBRvELa5JGMkdU7hhLkDX0rdxtUv6OR2jnFZhX176TI7l6YQQcYf
2CjjsAwOduPsUi0pW5ytaT9tohEEeF8B4BQxBjFDyFFMASguD6V2GJRyQ6in
7b7OAxmxg/FqUf5/LKK5iql8FI1R2ibKC6EzNaX1BE5d53AACXK+nJGFKQMw
aDBOQyqWdHvUslko14iVsq/7bEIoR5IIqkMPAdumRolsQlOdvPZYXl5FKfEH
OhRwhARr38nhoBU/ktKu5jKp38tZxtnmr7wF+ewhw+01UE1KYkjtRct6nxbD
s4/2hOQAU8znWWmQ+3WkeoDOdDP0GOVXPYTylA9aDer6O7jLveXEh+a6Z6QN
81Cic1pL3EYsU3aWwiGwEiv2Hv1oqVJdkoiTVggK8S0PBbIaAfFmNkBt1Y9c
bJN4uBClW1vCCmCIhGTCYplPgow+mrd2qhI33P3uzr76BF5fBeDCErxwGmoP
DPh3B4NbCYxrH8XMkCiMXAmJMHpmw6WVLpWCiSM/o/Q7ukFqACgLWsJGMfvG
dUmZBvGGJ70N+cbOPYf8i5RJi1lXLrYGsDte3zAjw0e6GvWID239iOgMtDWW
IATzFM2ba54H2n2vOBB0fI59Lb/NMgiaKIVPa74eHHurINDM9vyt/k0C79Hr
bhUgSDMfJBT+btHZLdJR/6yVRDgTH8NN5/RIUI/xM8iP+2XIjN8b7WVc/Bu7
Wxe6nYAVCJnyKkmoAJf8wkjJtBF7cHs8dHsCHNj5j7s2c6I9tk3lf2Np6LX8
GP9nAKuRjTnlZEPCj1XaaIrBfD5L6LGDahgDMOUIf2x76FZRn6aoR67Ud9iw
HHLNgtaEf6SDbzKDHzneI5UQbJcAv2dM4XuQZ2+0FJvY4+jRzqgPFtkFd3N8
JWO1h+dlzxC0W5pefR8fZC+vQmIXW+HXI4ZCa+phn38EpSMmKL9wn6m4nkEG
W2e6b9DsLij2xfERBTZF623ooEXMDjgph1oWZG1jP7NtG8h2t7sOeFAJTzgE
wyA1tsMUqg7Lnt/DCfY8/yy8bMksgVP3GTntrz2ver6/bZTLJegRt/88B0C0
FDYNMVWibfC4E9zrvfAmQ51UR0gWRT9mu+pDiaihbGn3QZxnETBfGQFp0Y21
30izQPZGwHo9WRU5RUAYx87UCsE1Zb8EfdG1GZqBMj3dPzM1lRdxELa2biiU
YxdMtDd0uu6mCE+WGo0I29PnJ94Sfshtx15mh4qrYh+eCZoyLya0T9MzeTc+
eLC/GWcgJDCDRmbDvrzkTVIusPgeKh8ieLxvktlG22TOL5OuQ56/h3dZNkCl
WXmPL8wAM2Qa2P2bLR0NR3NxSpFchodZrpgWpJgb154hEEulSz46rGUEzGH4
2zxuHYpgP2Rnfe4xlhuwM6SxvqcZiNvDWO3tBtnvu3uBWIiQ53gDVnLsktBE
1Tru6BCNWZa8Z04WHn37oCjDKGgA+8LW3dW4OhVhc6ZM8nXFJLK8vwihhIhs
1KD6XAyh6nZ9LnRNMMyTxNXj+NVBOcjH8mJmle0C1wjQ6JbrCvkNBQgpsd0A
T2xgUoFCPadNSXXpZGMzFKfTtw150UlFBQxVuVSunPf6X4Xi9/ED4KKVoutm
rRKhyK0eB0cmVTy1tZUHIoFw1z4hpEmMq2b+cemLKcucn2Sg2BKHExMXJ/i6
Uucr/FKHZcsKMwv5Wr992z2fgheERdo1nQjPHQb+moPNlD8hnNGUjA/kESIl
JdBMIgzCRHwM0Iy+Zfq+qnY6FesfCI0wkf67HhHAwkv3wcyQF6103Tlsc0cB
9p/Stq6TOqYuYHoGNonMtBd+aeM12T4t4xgSGm6XFnOAfna8pJQNlPWP3vIK
6yfqttjFjUosKvoUpsXUlTpDrWfFWDJoKVYnXsSUisVAHAM4+zfd3R3O4Vh/
VX64+BbvuViTkusylb+GW1De4QPeZa4Cv/oG+JNWgn3mWaUeiMeO5tA5Qkz3
pupz55ql+R9fYFB8WkgEjzoPpOxBymCl18a01J+Zbgj+I9/39Ingq3BE42XM
j8ZlR120lKxm3y3y8JJydM06fWTX6ytV7fUhOWQBM2KtMGAWmV9wuTK2E80Z
9edWXAi4x/OuM2w5Euzb5qATd79/K1OOPu2MMLOErtdABFVPJJ4MyBh6gXVi
Obp1whf917zAFpAQClbnnczH+cn8Jd549JnbK0PQ8Z5rYDqUorYRatD4PNDK
c2iek1KsnEl03sj8o5f3E+L/xvS2AQizocD08l5gvVSmT4ps1e2ItA8svzjl
kG3nV+IMOSiVTdF8uYtkBGcEj5US9wCRtoevrCx5sEDEwt3xOMzyJWyt3i7Z
MQLeHxXLS4lsWUdRFk+8eEtv0bP4HW8FbigMfBySGHVl50iDweEM6sG9F9qi
ZSxjK3uJzPEhyKCk3k3VJSf95l5mld28Cg4gZI0gFMWG8CM2/5jms+eWDm/2
cFrUT80hT1Y/IM4BagNIK6nr0liB0A3/sHe0qZXVz50HDYcyIf4Fgs7/tjsr
XSeEocDp1OrsCg25d8dLIThKP3cJQb70QaWl3EiSqzSKJLcb7BV9SvG55lf9
53OEUOMD+YHkycgazkmgql+YFWCDpbYc1t4Ww5VLfEmY/YezipPNZ3CaiueY
bRzLp1x3fgTWquMzw/JQ+Cyl5VSgB/e2fUcggj3UATK6KVM1yI9dYQdE1JjN
Jud2eA8dstw1E7BZh71ZvjcWymi4LJr5v0QGxxOo89+YrqygrDflf2VMr472
dFebFlRq0q+NCYm1DAMBhD8v9/0Z81pI5dnglSfldoIeX5U1Fa/GS0k4klJu
EIMXrzfwb22sFcr51GssV90Gd5gsCz+YXSn9o12XglMBX8TGC2U2W1hg0M0g
TvmzWNuD4t6yHxC3/R2O/euB/fArqP5qklBP+XcHdGUWn5zoPrnSczTw3fSa
93XmpxVP7EXdjSS87W9UlGQLKjUQ2lj57YL7eMLO7PALzpcmrjZi2FnzVkLY
QjUvo6S3G9nCIBEPFKisRA6KOV0C9xGW0KUDLdnD23GhBFYkkmqndKgg3rMp
peALP058/04MhR4Ounp4uBg74Pt9ddSILnrp2qHuG+PD/1x5kn4YghCFXqwP
+I9607ztWmGEj1bjpZXK3R11oy8WrnDiy14JIqNvkIVslVOEGr1HzgAXO1ZS
s+IsFU5GHswtTRPYYUDFvAyfw3yiWxHquvAx8u3fttOhH9nWdkIN0fUO0nAd
AQmzNZojQtP4NhynqgFCbu2UnQ41npImAwJo/xAsVw7Qw1kxx40ZeNpXviat
YVDtyq4oprm2ll9/yqehHXiRJG230oo2SUWCSGttoOhSjkpQGXfFQdBRjWVU
lVIkrkwkZ4FYQDQFJ2DKl9i2wkf8M8gtFZ0EKWF8BpE9cv03EAplEXxxI0ib
WfHNpD521fCsbeGe6ttvj0D6r9RrjNF3FokAt6JZs7OQNyvenueDjIWxDIrb
UAmgQmg5uKFa0kf1/dbDXQOMVVrNiuPEOHAjoZqhb9Y8+bc2q+7CXW0Ab+CV
3b/rG1fRp4OoppwsxGgyuodT8Kw1P30hi4TsXU8Biqabjweeg1wG7l7WzeS5
x2adDJGqgr1xdu1RJsYNDrm7fGdaNqUdeUNfS3s8mxLFFQ5z/Dg4HPEnhUjN
jPcyY5IHz2dBVA4vYI525LLvXGd6P51bCLfJnfAcawtHjl5pY5PE5LcMti17
STvZZn1clVy3VyhyI7WyQewRXsSgaj+l66ZfdREACm7rQ798vWjJkc0aaAB/
Gdy52PwsVmkJeNHbLwk5eE5OhhFK2NP23KYg+Kh8YI9p6AxxHWLHCQYhvSJU
Ovto3V59sW02Ly207Uvq7nf90bGDq60rFhEH3+QEvb6TK7Au81U/BSbeD2CE
u8uippeLNPsMnLEj/Y7KPHWZ2Ui31cl6WPtOKlEMKsjPGIu8LTaBK00xZpHe
RdNKmU18jvUGutokZf/b9Wei4O3oBBF0T1qKKd0vuXL8aRihHSviGGpVRUHJ
rqNGu1gZSgYRg/h/AAR4ROaC22pj8qSi0KLdezuOZUbT+5MViGs0dHIZOYV3
YPznJnU5LnjiyHwlsoHhmvL2/arS3W0d5NRd2EWotFbiedsvp/zyX1Uby3+b
U6aZ8MDLDKuvQ0bTvw3mMJ//CaPl66CsOZSyNPO4Gc/tZ7PBtJGB+hd6+uOz
zqkSIqZ/9ykOIdgkvtMV5PCuBHhy0PiSJddkDVIc7BmmkZ3B3W3HQvGpTebS
odR8IDrKW6DZdE+oIjQPWCRr94kPAGwa+61ISg86111Xi2LXcesCz8vL1dYN
oSZ7FXhWZXmETD57baHIgIRXLMMYPCf+Rwu4AXBqvUNg90lYY85/ByoiAbQU
SlTCIAUgww6Q28MhGjdA5KJ6LcUh2LfcShCPrOI3nnbniO1/FoAAuMzj0njn
ROg2jsTYbEarKt2MzDhGALC6gyzgAhsxvsCVrYh+GpILtXoSU2HItooGBQiY
4Xz/8RRiWmSNTNC18DNwn47QwQ/xK63iKauZ4hWqqFSGTBlqlrkyAo/CVD1l
wmbe/4hPUkdr3BthVQMn52/amdo44pAB4wNnKaWvPKjzkRSLS6j/feIfg/MC
+h9M1t+oSIk548kZC8izfAApmEXDYRMshAYbAnUk3rfQtcMhf72ntOboA3VV
QjBapqqie8IRdDJ0uXCvgdSiIAC/rScsSIQ8fgvqPKbE3+vkLQ1fWx5N8l3r
xBll4KFoG9t7MiJ6PFWgL89MIytlVPDS97bPq6ivTK9ukGujfW9hxEa6eeGR
1sXaRnAhtK7MNAGidxyZN7gt4iVKV2n64lFceYmKoBZ72Ny8MguEK+tPuhEe
tx57B2IDYm8imvomGe028k+MJTg+3G0OhEDco1Tc18B2gADMkWnMlxqLgGyd
jSukaJ6Jd8owvwI3tVMTxJvCFxFUkxTpoYzLTZ+HvwyPLgzwbdzhmJw6lZ3I
VTLO798amCu4gv5SK3Pi66MLTwfg8Eu4dlwmX3Bfmh92mBEY8MnD+TD3d5hC
TZhDOOhFj9P4M6FaL6+OWC7RFKjBs1GvYThFzFTneOHpWkup6iy/fwIczSAA
IJiP33+KVd+QYikdwbPdvxalEYmS1RAu8x6xgfyHDFtm//sXMar7p82OoLI/
BiqfZuSncq1ws4bMFaZWianBk1FS61aF87+thaPn1kuiJdYUqXaAEVxf/hKE
TnEtYxJ+rQ21jmSQqnHzHUrQyAu1d/qMzY9i2KphL4QXmN8tgEKz0mgzD+JT
Sh7pZseoovIUU2g5TEEXJA0EK3DzsWFHfDGz2nmX3TGK6e04K/DkXPntxlr9
lNGdXPsawzc1T4S5FHrCNcECAaCIkKvCsqtdRjj1f9w35MOvJr/s541fVLPw
arPMapiR651CHARTd0rC41ObFCwyGyfCx4Ql87VeBsYGQ39GBNBTy7eIRLDk
HAA2JW6errqEPooTReJKulNNjCL3fZZzUYTcsRCd29dPmRNeTnA9btnaI6RX
FuglNo/aDjc1XjPboAVpbd6fzjONJCSWA95j8gdFxk7E01KbqdesW8WmME25
5Lh2+S8dz776Q30psRqHY79N0eV+U8wEs5RWZLc5OB49Znx7ywl1r8AmvJDJ
L8s2VbVt1qkkIuothhIIW3ipBwzWTQcLdRlAf3H5nu8p8HE5WzQNdaoXTk/C
6zs4UwVp6+D6U8fdeU124ag8vUp8Bq+Szvy8o13fzbR9LEw4rIoBnT4FAo0K
ETayeAuEA52+G+FD7SP69oU/ddCDZ3NpFQnmFxXq6lChKGM0O9TKtlyyvNz5
9h8KoKHchUqZTUVEQFPZRUwwSsU5AATfnuWgnRtb88p1J6G8cqre6cIL+ssP
5bx7N6dwWWpoUfs8g6fMom4DRuPlpcQ7aGnIX+xeziPQYq5A3N/oKr2Loian
RMzJcDWH7C3puiSOpDaXXXzuQiNDAoeDbySfOKWCL4pw07Mepyc+wsNVUs+N
QdvM67vzXhdasA8fPCyREfQQOD9HJo6N88U13h7nWWv6inbd5DsxEV83uJkc
y+9infia8bsM04mm4ZLOuyBzNKpacG3OCG/NBogjVMkX0XRaIrfZxJ01Cyou
eD4e4G1DlBpxS3cWL+9lJY2PXhZC6ozu33V+nW4MXo0vHpGbzvtWIDoR6fkb
nYXMWwZxA6bYnARXU+lYU9zC2iJL9eTfXimm7v4YisZ2ckIu9YF1SbW+2yiE
PSr2HkUut3B4n+4iQTC4IsmaK0enHLbdf0LP/mqasHN22/LBpor+KanxL3sg
oMDX5L3kt6bin4gvfeOfwehFPfU3+PZC4ff/aqwoFznxXXwwYJz7ysgRETiY
mYwU3ZMRXFJXdKpx1AOuATrEogtjqP2ZvgAY8eJr2Gw+Cxi58J5yG3cUwgKS
FLkvxJtFMrKr+CE3DTGKMuGBJ5m5GN33C6H0UbrLIUceZQPE0TLsrWGU6x6M
BpteOskoehFETfHbJnEtp7lNUzrG7Ptt+dbBVU1GxWMh33Io1Ti0e1kurne8
lStgOuh4it6IYPQX4Q33W6FQfG74OB9HASGLcXFxnkRJxJgAb1Hu9ekX9jFk
Ka8iMit7xiYIyNk7ey+3UxNfkNe39HPH+zx/xxCM+JkdTryQ3krFmuHXkVA1
NqA6DfDaXOOoE47+TqQr1UAX2Nx4RwQEfrZlXOAe1Crv6PY2neOyG5ow40HU
K/25+l4aRizQYWiqY0KkFPEECKN4WP/2DpVXEQ7zqHR8GoYiWvdLS5oiQWcF
A/liO1OlZjcYTgV6Fq/RkZv0NwFBOM2zbPdZGgv9EO00jFjk+bXDhQD1laT7
4Kq8FY8Q/KTPb20zFv3aduUa+1bxFMGSQ1Joz9nb6qzHFYVE/IpUbZi0Ur61
MoBOjSKRU4NY3fYFtV8KI9HYamRHURZiv7+L4nXe9TA2tXkALZJ98QFTLuJ3
b+d2zBtZqTQANCofwx9QEEawg6oFy6VAQgrwnhsmQTONUKebw7Mz+XJ0ShWz
zy8SL+/gNQGdxBmYjvjDzWbgMGrweIrlL1AGNgIsol0pa25MsVtmwlp2D7ey
K+ugrkwhO5QCWK6i3Qv/yv8OIS3SuzqEDazDOPlQHY8mPt2D6v8FhOcsspSM
00ZjlH91wnppTOmXON3SB5IhhjuzevHjDjacKQpnfuvXKBX65d9UMzRPEb1Z
DlJtoegziDWoP3VlOWnzzuYjUqywWJpAmm7g/xOj7rjl/UOd5O7lDKXih3ps
VbVXqtVfwbiScduiREPsm6skhKHW9jqZKbP6OKRmuQklqKBTQZ5h5u6H/Px9
UvLfhwj4OCposOBUNuoiRo5/nhA5kW/D9XNGLCY8zK+9Mf6VZPqZSEenR94i
y7Qf964n8i7LUrvQP8E+3zEkBvrZdzwjSrrQF/fV3ZJqQn+E7jtyrzip/oli
HkM/wyvea6TzeplAbOkFi2TxD72DDxHUPBbL2oIfvjOS6PXAMov71C8f7VJl
UYIFAk8xYjUba+le5agOsn3M/4iTWXxl5LxcbLexeq7zGTp4AIE9qn2hSsdh
JYUOlqCtnYbfj3Mfow4YrntqN/dQwr7b66wzqlZROyMzrJinCDmlSwNwlnlu
V5fJjl4lDmc3jlraRupIUW+P1wsjG/EA8XD+VcBdoXKcKVSCEVAeC9ICXO0R
PbgahrigSDm3GaRszLZTUEdbvHtrzuStKFsCEVBli7WFdZRckH4S1FyFsD8g
FwV9kvUompd9xZHl18DLY85UWLuWgQTBFyUgfJigq1VkBP9NF6zGNCPJvlSf
Dr/9PHXpLrGoh27f527OeucKTeNCGa6j1prJIW4ByTIhMcUgT5hZcTcSYstK
Ce+655b/Iq5vPB2bTWYihBT/qSRLv8o4krb8/EzRtqxGFPO8GWwD8QFOIfeT
Ii0sOmQujpOfdH4zkPOEM8K+6+Z+6m0aAhEiG1MSZyQXhE/6s1LcAqpLxvRZ
Qk3oiHyleLLqgqBgz3eiH2yhtO47po6pG2GRC/J/2yA9EzvBo5dy98tX+iOk
Iu+ocERCP2DUGa7W4+AzUtBJUEb9mGPvUOXJAQQM+KQyZJCyPhkjoGWwgkeZ
SUVV178qnR9EleiEFEH338dtRKnJWBMt+gC/DQ3hEKJAcMDLsuEc2hDfD2MS
IexCtzy6ZEhcPxar0hASt69suT3kXz6vRrQ5ioWKMRv25W0aFIKzGB8lh8bR
lIXgjC7V+c1srD52vihp24b5hQ9pxPmFwLpNwHRqzJL5bEZwgAnuyxpFP6XY
7lCw3Yl1Txwm4q0G2oRVF62HnvtFTMtGkB+phx8IFqi4lKWQsF2eeoX4T056
xRTJG2voE9s53eYDT+lMe4pRpb0iJa2XqPV7RSIJrdp6WVo1Q5Ct5b7Rsq2A
rCbQkNtx19470AX627d8T2Qn2Mnc+40VB3B/2S47fH+h4c+LfiaWgJS0PVZU
M16mqcG+hFaFl2ixowt7z4M6D6O8GEzLbAhiXLQsikon3e2oR+RzK+S/m+zp
L5TUV4ecmlBneC6b8S9HkHn+SBqvj4hCar4KXOuHrfmOwRYVvy2P/DeNBJXr
GM3BaXC5v3YH/0LxJ7lXcShZWTfWaqZSSjKfVZtacOXzAlfg1OIDdyK9M/Sd
ck7PsFuIh2E6kiLPDf+ncjuH/tQxrz6A84OcKIwFuQsDFrRxzQTJL7OZ0STR
tX8DJbXcCDd4TjhVwPLY/NGA4rqal4OpQ8A2UweM+TXB9zP2DvlEvZoHPZzy
aL5C0Wl4IEeRQgOMo1RgQaYa+hi8SuaCtqx6nHQtUJvSZ+M9YIAVvNT6Pc67
P+3Ws3pobQxLwLyZuOR75DCDBioW8EoCfTrhAzVWFm7AJimCUKFG/CZPorEn
8wT+/VE/iAaqjH5BbWbIdvNldwcahWsaua/akrHm6Vt+9zrRURtkGtslaLz2
02gcD3WbwmvKE5MWkTSavbJTzOJSaWV6Ecjgpsi0enGNypsAKKbN5F8hnpQO
1uOzKNpwugLEne+kaJzPKQqzWQsTMhLxYQPoTbkCYuG2RaGnzBfz045zSLJ1
a9ivbXxkIN+GiiJH25EJH8qDv8TOPF/qfCzW4R4/77EcRmmK/Ahmyk33i7YB
VX5R3+jDzmNe1KBAv8qXzYJeF7eftXLZHkj6+TiSIB4s9zuTpVN2g47/W+WJ
CSA6TNfKXSAhRhmvwtqcD8Qk1mpqhwJ69E/qAzwa0YgHQUBDRT23L0IZHrwm
/SSoSsSXPSptaxfb9x/fR1Sgb+BB7VVOXK1mFL+V3IyJVb2ZsEGJaLgGs/Fj
nFOcawCO3SQWMTkFp5C4xooq3t9fw93AOuO3ybabZ3KAE1ub9konQxj1DfCU
H6MoqzjAnN5aubzIfwq4aALcPO9ouFZ8//KSnER3RsEXLlnIl6495URLjYzI
accimlXJOHb+VUYhQepjRtMJB3PJ22tWVshA4OJsbt4lZsYlWDntvLm9vfS8
cEdqWd3XcrQ59L7DIj/aPOSf1sBrE5A5es4wK4kjThn8EhZv+GiqOwW5HPwL
HuU+osiRzYrc9DPVMCB127PCTkQ99cJSY0Qp+dW3eb/4HRBNBUBaE4kkK465
heOIMGi6VpFCZiZb5tKem+eTdXtwabsZnoysyzzdFEU2z/LKL9MGF0EkSwoR
v9Kt+dU1GnW4uoD+8xTSs/9tzFt/2PR0e+vytET6CTQ/Z4it2ITg39VBv4Sh
z0uupIl5NKW7gHhZQGTjEA3EphwkdOQ4vSxr6JWUwXMnEi/8mQbYhOEcVAII
h8e/ATubav/hJsuqzqGTgw5unndK/u1yvN21AKXmzw07luHLSDtlGCEBSi8w
yER0iI63AIgyOBJrsF32mPx/beuoLVnlh1K7QUxQ8tSp+WR0AB8uQc3CRsS6
A5x/Exa7CfG5UJzsTiiJDvILuxmCU1jhpMccq6G68QzODmCFpddRdmT9okMF
DXjwyi6bFjAFZmZOsBeLvXhsxNm1F25ofXhoYPzP0f6mn3DtXNpU3ChKDgGi
ngBay3mq6pPl9RqV/MZlSz+UkWgTkY767Nbzb4zIMwt3r9CRaFuWfohvdMAj
JM9iuf6ahNgBpKD2BBUwKiRQxD0NcMWgutbzlZveLzBcM/7KFQx9PSPqLt9a
V1b0v0upMgvHjYt/zM4wWAK18AkJYxrrNg0jWuN3mUH3GQz68WBcOckCrLpw
T/X5TZn5mBptFVm3VGnElR7G+79qTAGP1bNDecSDPP4fa/IlqYtQt5E42vCl
tuXmzGyv2HAAPIOpKF2PuEM7CN7blg6qq7fPmIX5FTnA7SZcIJ21HsCcYIK8
SvIuhqTXL8Hhga/sWTwwpk0u/TpLXEDJZcfmqNFi+Si+vaB5JgtuwMFrkkEg
YerTxPSgVFZJB5r7oKPD8/ODICrwnD0zKrPm2/MLweDk1T6HRbpdlRaDnrsN
B+8sGwaiDvLcNzFVTKFJ8kxhucXMUfsz++EvmMVpEuPFMKeS6QgFuE6cSPqr
e60TVB6XxpLaoX6HAagkN/ucikej+I5jMgSilIE5aLgGurrQbf5kkROadp9E
2AP693ZrSm0xsIviOMHo5hsyq1CaqA3jNoiPhf5yUCdKmGkNp2l4+lq63PMh
LH2bYjocx9ODWhBzeq/IN+5UN2Pu2GL8dkkKwgbMdXZUoT3ScSFMZmKedBj9
EoI8SnOcVdwMT3tmDaX96c1W8meW58YmHho44K73KtHTd3QYcMdNoDM4rS42
07A5TTnN0ywpRVC965I+yU1PU7ohTgChK1Ra0f09C5AxHtcxpYJS11s5W0Op
z3qRy7dMOP2H2ajYZoG0OPPObHGRcjpmJ5BmfQyPZ7fLAbNTIHeWaqM5HOqc
Z5RB48Abwc3kXubGi++NhoIWPwo04VBkJHlqAQVolMTZBJaqSp90XLkV/Doa
JPgXp6GM7+JwbA/zaeROp0HP0JpuaPJZPTzwcaQeUikp/N/ZUNZzPCDY4kfb
pnt7uR7+hxLYw1YQ/7Ue9+BsqzZElLAswAyU4B6WbyiG//gybcf3RFdIvJgr
VPYImwEJ7wDeeXh73p5yn9PtkbgvJHgtzHl1qDzSDs4JvZjm5scYb701AtTF
QDgMbg4goYcdWq4uQ9JS+JACxQQyMaBvEi5xFwQQRfBfdtViUAgJtygXxIBL
DQONYVFPrj8SEkHRetv7JKRAyYgWK4dN3K2Kg7ssKEQA+gDPO5kVwS7+oJni
2Ec13fjI2Q4nQaPwno/WaFrTPbcH9tmzMOyLSZxGnuUr6IXz30cvdtRzqv4J
7UF2ZB1ylvzADhIZmzfOVWcwAgdoXZgXsZ0O3+KbOAHObJfkGgc3q2VX7qRy
FW20JYn1NL58/ExouAEGLScytCh2H+Eb2wF9hJnxDSIGqnXqMTqJMSak4Oug
4ivh5GhJJqSGlR2vNZ+vNAihipVDpzm5zVOfFKecv3JyRHc5en1D0HlF0iwg
pqNNAKoYNdD/dvqg14NeJ3Tfy8P+Oph+QEU7+1xqksXJpIYCFDvrF9Yki6Cw
LR7iFWQ7vPuxFDmauGpn3Yp9yF65OkScSiApiGc56NrmNqL8lqn97s7dQn9A
bWX+C+bq6p8PNkBHfwzLP1kdkElXqAH3/LN4BfzXA2EWc4b48Y7HDsU6sQxq
t4Xj1LsPZEY29yir6yC/GntYFDfFr91SiiGFmlk3j6q4VeCOUS+2lUZw/Ovc
tVb5KKOUrcXoyVSHe1uNqXGb2dTf4OUfirlVcBct0Blacki3C9bPgSGOfXFH
fReTSiYPTPW5gZhhBWI3Z9xYDDUF19V1xtZHF1+Buvqw0SO4ksNv8Q85cs7d
I2wZTdHNhbmxw5UTymVcrN4c9IgPCbxz9AD9lMuRTND0ZjghVB0mjERieCA8
NQNJ5zHpD23bRkEGmUjuifYxwnpgtKyuvdV8H0fYJCOB9E56t8Js6P5Z01j8
ssVSmW68WHisj22WcYkwrARfgwgGYlWeMhutQRUAb8pZRJfEXO65ZySYzu1C
MlzozwOGxnhNd0SxjOIkqPfYmVbCWUS0YwVNL163Sf0a5Mwm8GOEl4UYZNGB
LKSVKYiu+ulSX7YW06+SV3Y/+2KMN4p5CQmPmxdzpok9d61qZUXW/K7EOEzz
KlsS0bDFEymaBCZKMFCbexJThX4Q21QwOJ269EeNPIWgvgSYHqQsKkFc/M4b
ULqXFRZBl7kbZryyq5Yhh85HjhvZcyM44zjlCL4lXg11QY77NnqnJhgRjTYt
dATj5ln4049gSkz/1uOGSwqLAOiBbnto0eU9Qjk+EYehtf1Nx21Sdmdv91Jl
It/dSQiwps//aKRQd7C8tuibrlnwLNAmrronnUeF0HG/DPjW3hLfV85uBxGO
Gr8xlRivT3qRa6BG9ewxTVHbdQtKVxY1Dw/oT9U9wsk+U9UWErAx7PxSzNRj
CwaVtHiybX+vH6tLRCPrgor1FmpdWgRthRvoWPc7tJ8WrBVQrVvI2C8MTiZ+
0X/PfJ45hExsTAEMwYKXdNm0BmNFYlG3yO2WVmfWNgGOoSmDcxbMbxlOqG4c
qR2HxjpS0GFqTCoEEpfLLSCMjG4oic3OmILSNAYfVsJaPb/Ada0arWyq2wwc
vLnWsGAl28WM3PIZ9/+bn0PVLvWBcHPH0Gt10AYwSTNZUColCaKqtgS/6N9E
4i0XQAexkQdI6tnQb2CsK7J7PevrSt1Px4Aa2NzDMGlb1iHIpLTcbO5zRdzo
I2TEZesNgTYfAhRvEYDW0CRB0zxuV0ZtEhG/ksfzlsVihGLfXS1gtkE1pBJR
EMxIEg9Pc1RH407RG5LV8ZIDpbUz12wcZ+cU7Kdj6lrsdOMpOSoUp+NjIKlS
EjspDMztfbKkOV/fGm8gE04+iIEoCaUhHQnkKA6/zPJtSh/tv9s9N4kCBt2Z
PbGkKom/TL4fngQ194IENwwoz54k3iesVAvase/qKN7rjowrh5VWof81lQ7A
hanKaZg5zfZXrJEtvvAQs7037qAVYJztDjXhpBr53aOsef+ME6MLOzUhN9LL
bVATR9svXV/5OlLAs5pGUc9EZc3xMqpgCjgf2qbvEgEnbLFURDSnOEIOmnJW
K/gVJA2BZ6b0Glm0A8cLLObiOyW+kV52OxPpVhHr3MuorRkwlJbIKZEpXe7z
9NujwBmdFM0oGIPVA4abCrhGAJ559SnVwxQR1lfFZGofCkgRefEXfyeC4oCg
I3617Gf9O02NdR+82ahorJCaw8GGt7dMyhF0ZUZrn13kGw8VaY6ssIchQko3
dwK5WuNvl8T61E03kT7SJBFGB+2oEogOgvqYFObmY9kElSshkZHWdQWDLY0x
RgLQv6JCMz13cqX+b9YB8cn0Ia0a0GL6e75nEQOQJGpt/SEEYlTL7Ca32Tr+
15XLMWNKAEbiuktHKWUEKWPDqO9Y1YH+2nEPBPMO7Gm9KJvxHF6ivJgdrsLB
2nF3GP0yQ7814CPcz19e1l0s46RJYR3bMiqwYg2tZtqpiPT/B2N/A+EgWih1
YQqABXYRB7VQL/fHyNt9hjUehz+O0nP6BZDucLYj5DO8IcI1KgBbqUVyX1fd
b1gPzKTXtxOEFJqVOOEPdTm2OHqL1kARRa81GrgIbyaseYNiZB4GEZAu0W+z
LPbyreH0GoJPFw6zAEisx843s/qbLW6pm1jkgxvoUga9CuJBIoqu1TrqzZS1
9kPDntMhQIFaa1mujIYezftQptCaX5VMj1U4ZCQcSqtlnc7sleJJ57igGLKQ
QyWuY0s9yRolwJ0sE35C4Ztp+cuN1DuRbbuVIx2ARxolwAo5zsPucuXUimpO
C22D/XDnSj+XYwRg5nfARzSBFGXErExJ8ISSNlI5lm7JKlkTYByFe6KfsJyl
bjLjSI4WjLVw9Uw4LVB+Yt4TX+5ogwiY71jy0GEvAvLHkx6nMTM6k3Ut7ix1
9jlJsnEu6DNc3D7aWDbnz1j4mRQaxJtup/HCsiWX2H43qwwBuVqLR43hJuVU
hi1H7zEMwVhqHKGSfuzNapI5PsF4HqIRTRtfLz5wi9oKI7GKKe7/8uE5iSs1
0GCVbVJXg0dD9KvOuTet9Tc7e+XQCcW1nnm/MRIaHzq5q4zSBx+/ESDrtUmx
CyazWEEbiYHSSbkcVv0iO1wtcxZ5DQN3poGL1uOyTt7/RJpeDjygrPt5tTDy
aEVjDNw/9/NtUURI8lg+Sz2NLlx4CbP7JKppcLZtZcYdG3xUN7LSfHXSjMG+
LImJFb7PQ1JAiBTgtTgL+ShmIAe8fO+sm9zXBObmmIrikkVqMpiWxBLnM0Ee
DYqCBQ8j2LKD3f1NFVcTqXom3kf9DOvnInS3Mz1Mxv6TRvSHqo2JCPf/AXMz
bfPsrRabRZ6jvyy0zS33AIccppTO1pGQOrqEqGYlnFGfYN92KsIlLJZarUCr
6bmBOPY+0jF/+X8CCgNRAt1gDWewVr7PtQHryRDPwqihYvpQn0JCrDgc9Nbn
XVkjwZ5pJuoNP28jsYndVsplYATsxgQn2FtPJe/UlncouN6QP0JBsBP6kWm0
69PUmKbpMI5SUgnKthAnKIgPNjKq0KitOUUNSfmbpAP/5wgxzpQ+CDkOT3Fz
GfMdzKPok316acG0iiIqAa5S0CN1RSd1qahRdI1wtSqJ8cvJ3pkneA7CZk56
u2LiQc5pb9xZ7kjPs7Lr+QTbngAYbtkLU7W2iEn06uWJIoZaBxjjS4QgZAty
L+80n72vNnyTCrpbQfw7XQOnrnLvRah93hBCWeSrZr7EVIoUH9Kf44ogvB1m
Bxtpk4wGFqXceQkRWFwgg3Ss4B3Kp1CCl+y//D23qbouioQfqylY8hdyWgVb
z7Ur4k+Izm7n2f7uTXKcuV1oQf0GydYv32MvbYikxYoWkUYJvBCEFKzaP2rf
r8xNi3THeVpBXWrqsKR6bPWHA/d4tk8VEjQi3rXF2OXIHXO3Aawr2uR/3Q24
77jhM4+pP1HAWexoHScXSLeAgl2S2tT1ax6zT8+hn7I9DgywLZ2O5OMe5COE
jrG9pGKLoLBNH64kQK+6W22YsJ0SRKfBBdjCoglc89OFE4nYWNGsVKLy5DGB
FVh++R45DA2hiRT4BDsM9GgKieZ9fTlGlegGL3Wb5qtUyY4NDKjqIC2/+19+
YSyMiM+minZ1f1SRjD6wC0/YuLS1bjgtBJnw2+enX8mb6j1ahS1qIK3iyEzL
LaVuDHhZST+fiP6M70lGsZT7fR1YbyrQH6RzWNnXn9eJfaL3JpHKC3oXSZAD
ebYUKfszn8vtnMdziXFCXdDe5snz50B8vTHTIvPFjOuUYSpgfkZ4ZVx4i/5S
fMFTEv08EGgFFkpu0VmCPFXHJvw51oW4f0gwzlabTl+obnaiNFAz3dZFUjZI
Y/SvQJlbr+/dz6UmGce7uSk4B8Yhb0pDEU6m5D6h3q5EDP9hDCHqWIvnk0Dr
n4WEtLyNmX/keY/j3ehKl8/Kh1en4F5wZUOCYslQzjLLAHT3GGoP/WIyyhGP
ybM9VWhoWN6PVFHbtCYYn2+reOFGi4YtWx7cZNpxmn3rpgQpzIkWyaof58Hh
PWIGsDEiAuMNc1DWNfevb6vKK0aIzV4oLOi/RnU8PitCywymxnFujyFhjC32
PKqCI7MAYUltSNVBk7j23pzdW738nUDiyPAHIoy6akTd9NliBQVb8hQtnfSu
oN4p9mFJJ5qMmBM77xpexP03GpNrQj+xM6oLUrHGr4XbEnWLb577rkoDyoK9
rQxxEcHoor83RehVAKta6CCENyammlUInrJlh+ZvSefQzl9wCdVjfagAb0Ug
+miVqMWToTDr+SbVvl4o7qOCmS8CLVJy8rTiHRSskLal/aOMQ3KzYp8NV73b
Xl+7hVfuzBf14CLaMIqk9pUErCAgz+rY+fh1Vo1MW9sByE3WRtqLl2XZUSwO
dpLiIT56I7wXEO7/vLEyKyJRWvw6ABVwkM5oaS0cd8A1F1PZzC8UwnwtIgdE
IM+NVZ2Fai6WqnXN6EwSwHyrY3/KBmBGguYrDwaB5WfRAj2yHgV3sTp5EYFW
KW9gSglOp7LAjc7YyzGualaCX1CEbr3Rqa36LhgKsJEcPK1WqwjK9DY6Hsnp
wUJRoeWjJzeGD45jIPIV2ERhq9PFF1XKuPTkSnwbYrHC8gb/4OgHAIcpLpLb
Px7qJSwlB2tNaE7xvlr5I+st/Mgk6RIUwu7jg+z/BJ6VwZfMiWLyVhmKdVBU
2dDb2U38ntwJfYUz2AmCctG/2thVlsRjWtg+BeGEBXZNOtc/8GRmTwPXjNwS
/kIhabU2a+6x0lEAh+ocbNdmU6KN989jN0Y9cQHAg0Xe719E45TQWARk2HPV
U2hcak1JhrT5Myq+Ys1dM92B/LqWZ7vyWG3llddcYswXLwGEgb+03oWT10zS
9i2qhY5A6EB//vSrX5WFTbr0Gpf8f91z8G7TyrwLDmaFMU75ey2ukeeUgwB7
TIoygBf/NvJOTZA8vMoVCl3SguR0fh8wpMwuADZn9HidP2sompFpCJXjDCAB
Zh6rAAREAvyhEeUH7WElExllQOnF4f8EAmZryMKeRcdk2z5SMO+zGNYH8pO7
/fP2LhP6ZyqsvDV/3vvxUIugSm7L4RbOdVAOHK+VRASA1CSws/6IObHPJpmQ
3a8ArGQ7mGezbwryIqoEmvo/r80hQ0vzAQB/GTVEB5biBTbsUPTplq2jwdfl
UICC1qAEnxxzNrvFJtigAno9jFas/iICUX2K57dqQDlxwMTDQkyWImx29FHs
D5pOZEfqrkJJRYGFwv7n9F8TswpraxHfaq5AgraGrdMrbm1pp9NU8yYUPz06
6gobuj0DlwiAMRqkgM112badBKAmPdiEEs0kB5DhrbwPtwj85p99alOYXgMC
l7rvzc1R+t61my3aAF3hR2qEvF5Ykg6ig4fz4ifStC9VIUCevR2eD8RSnvCG
hXDBS3w3Ta2eO5mPBtTQgrfvXkG7yCjv3r8ODsTg82LG/Ddd8bitA/0gkeJT
p4VbHrETV4kjd1U+pqcZS2ouhCDkVittuomw5QhCe+IMQ+z4311WMx3duCB7
0a99/dDlAynEnUaM+YyYji4G9u+YQUb48+0rOJ4dK5nsLO00ks7zWHorb18+
KuKHGBfLrdVwYe1xAaVaeTY3OJy+9L+grViS35NFExcjlfLAybn7sHGcNtux
aK6zExiEakzd7b9K6WggiMfLPLUw1pbPzpiuX5QB0T7nzyKoq1uxqnWR3C78
hoLTXk1W8e8HD/jRElXzB54u14ibOkaXdJ0R9Zzd2wkX5bpExPD0p9vXj/07
smtKsn1pTGreDOEOU76pIYbci7sNQYbdCHdX28wnrW5RSUduE8HLViegnuIF
ZDYhV4loTSrWrY26wvCuWSKhphqsLGiI3z8MA8IJOR8Afkd18E3QTvBDe2vZ
DUyQOl6VBdrZrOQ+74ZE1TJXZKUQJa/nfU/ZpsUxMqucXDaxWlGX11rIP1pX
cKMEzJOaFJpxMuM55yFLKNrnO4SxPOcwxOmmQVSZhivPWFZ1Y4TOuxLD+ABg
EsdWG6+eERAec7Xl4OcfQKhLJdzNYQZA0MOs/VuSkA46dg68OrhNkaDppVN1
9I93f9DNViYrdeWhbJU2pZixfv1g8dcNHvdEePe2A7n9cdthZ5b65+seBfV4
NTacFOFL3PRyEHsLbESaDgnCgIXcijXl3CeHVrT59ORkih2Fq2iOxYt191XL
oBAnbgxfVd04lLiyHgSAjtILujIDm72ywah5poLG3xNpE0U8WBOUnpFX1qtu
ApZBbijeDOjb6Eb2TyfQkYwjs41kdkZMI8/rzOZIDLaRgWW7GFYOIpE+kuHP
bvCGndDclsxKQNIXKJYEzx74V5PlBAmRb560ZzI374bmYtVCMjnsoCodwj2m
9mirkt1BtvJrrBV38a7O4fjZqe01MP9bH8y4fZq1CGJwMgmr3T1bB87nq6H4
35E+eR2JiGFOSzGcY07ZzVZdgA4snhS9tyY1VxZvzplGklTYC6ji4tXIUyc7
EzeLlGOIdXeQAZ/i+WtLMSopuLpvIq1wav7ogPIWZwgNpzQZKE4g84UMHjUv
91q/wYIjRdpG4K7uW4NQOs0YUxiU0CeebnCtDG1lqj5iwiGNMEzhQ+KWjDPA
vgRIsY4txiVWh6QZlB81SGSLnBq0cFB86lsGIMP/bdWfkqRfzP9Hs4oCSRJ4
QJhRVMDgHBMmsOjI74qZYkjmjflbpTLQ9D/0EsUls85skx0FDwuzlKbDGWZb
LrHkls4hEP40fk5Vpg2+XMKRAG+HjrJ3K4ESGOzlg/yuz1lEK4ZIcZtbOrGn
0lETZGVSq5ZePuPCxHiLq4+Jd22k/jVp4PGa10FTUqy5JMK48+1685vkB5mH
UefpZXf7Pw4Pc08HT+tZzoA2mNWrYqe2+GzQhG9Si5KnFQ9dFDC6ktORpjYa
onjwQXtwgXpYqmVkcZUBrTGEx8UyfSGkq/LPqqyn/kAS8YFa0DB52i5j7bUr
VS7vunrxFgDS4LxoJ1jUB6Xb3x+wlj+8irbeVsdpMqNvStGz1nsUGhqQsHae
Rku5o6737y6tTTqKxvRMjoxyAkViUtn393CzqUB23s1H/o6HnJSJtku3lhqg
YsENI/POhU7tcxANPLWqJqUb6q548TGkpZAM5Gj5voRbVqTz2XAZgrWDez13
lchv6/IkJqElJjXwQFV3ggNHb3UGOgrVhQzyLc6PT8iZvGoFx1gD6MCoLdah
F1GdyFMr/gNE7C0F1+B9imGAHPeAhRgkSj7l5CfI+vfaxws1EY08K1Eg6dA2
2kT/Xb++t+55de7dthAZyIPXTrNUkAupu4S8rZTmqgA6Ne7nj3bmQ+WMkcUc
LywSCw2ItpodxIZsSmkIHFMB49c+Hxl1596buNoOETYPculXVsjoCjRz3g2M
AXwBFtpqsefCZjcJkJtrqYtF2OY/K7bY2DybHR2xvR4a+yxEYw0a16IczovC
AbCooPbVSFFCk7SdzU39P35QvUrNzOpkQytz6MxVqFJMpEPL3B4WogeP5CCw
FgcazRcd3fQSdcxU90k+bWyoGYkmz6psUxLBz6xywaoHn2HOtN032UOPsszd
ICXtmg/lnvtdqUIOAW11y/3yC+yTbeNoVci9rbQkPm4g0Tm9yfNx/mUlYYDk
EO9VeUujoJXWS/2slgTxqL70JZ5rBABGsqovDrlaGB0reRMC1xL29NbaREE2
70mpiW5efG4vKUGmWS1V/4Es4x7BZ01X+S0ROat7MH8EOMxxWYGqzPhvblAd
q+VUSnJF0Tiohh8oPuSh8R5MoCXy2h8NxQWW+QyvP4ijZg9LQ+GOSU1MV8mS
Nx1xdLsExVR48dlqYz6Pu/Qpk6NQSYSwTYzsOTgOQ5y3lM17jlcP1wt4o4O0
lJjn/O5rQuSFOKeBI5flVpZJicChPVVxP9zpwEVCdO1S7p1NyC8S3DmVXW8Z
EiETxlSmnJNTwGYNp6+1JrSLM+Sr0cS4I/qNSopgXbM43/HQB56DZKLwgMBm
OpnxUg1Ji3e2Wh9G4DvGiKDsF/QPwvpRsZBJccJxSJP//MRc2MIdf8kP8n1y
4Q94spxbrBeMHwiC1nemnponOpUNNbs8YSyHwomCmlunMlzeDFUr0MBseDs2
c3vXxhRM0ZxqeL47NeKqI1Kg5H7HIiupV+9qfC6TH2+/rI4aPz/oGQbgE0mw
WqgPJJQyU62nu+3MtYk8Ll8/fwAXBfSC9XUZIUmvLtNdS6VTmkXxUSi9Tn5h
cIARVefQ55LM2uKCgmxadYrwjSLD5nkhu/fAAkxYSztuYyd9TD4o2L+DuOpk
g4EhSXhURp63lIOMdTO/o5y7OA08nLdUK1Cyfito31f6gL03Zv9NI30KRfT/
Ux0u4lRN6FRlnQZRpz3p7DeQ/yIFUiQJmKSVN7GUiW4VRcHfyPhdFI+L2ZKx
HqCA/g+YusGr5v/HFnVvmauk8zp8+MsALqgkS0qBExO/z/l5uJyD6WxqjHxt
0HloCKGPYc6eDEZ+WvzHBLUjJSMRjbjc1uv06XB48uJ9nt9tOeHU73tT4+e1
WZ8csjAGZ+SFzAHv2QzWAQ7u8Gg1DiTs+4AVthjBlpvKzdiE1VAGm8zUB8/O
PQAnJEFjuyXt88c/wsgZ91UQdCdnvWn4FrYTp5lD8nixZEeVDzKoRSQwvgld
5biAPHq6m005R12kZIeditdm5gV1MY7SMYiY8jOphSu4uqqhNiYz59KGRFbD
RMDnTUlL518jUWe7PBtMLj6CwIxVmZIpzLEd81uJnGu3mC2i78T16MAD/o6C
wgB9DPZ6kY4NNTyH5euxFpQ7WkUjO/tyQQzZJxvAchvtvgMLmxonxIkEytGT
BJEI4+Jfex8f4a5inSZGBWW622KL79txBRlVYzFiRRkj64+1GtWZ4f2GUIDx
Sw8iBV28OYNThGFlM0YpgTcO4XsVdBPJftLOlUZXmw5KAeHalsbRKKXe8X7p
PmkvzhwfttabgaooGeQiaunEsPJgga/J8Hr0wzruPiqupKsmu5NiXkAnpwEM
GzozuJdceQp9WdYEPlzOPzCgWU0X0MOPaflpQvdBV8+H2U5v/NiAvb79dDkj
j5JuSI4Xb8mc06Cs1oDWwkoaLn0fIH1oGEvE/M2Mou1FJli+u1jSOCnjhTXz
ul1JkFkuosnQ4bp/OnvHoDTV/w1lk2EsURLHg3i9oIb+n4YvC5xeGeX0o5v9
MpJR8UshmjFeUdfEBREGWqq8gMjelSTmhVXr6AHLSY4Qvd2KNlo2Pp/XmAUF
206G/T6VXcZZ6g9xl/2fYrgkTGYNfrJYr6hv5U4ZAT/JzPqdLhVPo4hg3wOx
qAmU9Ki+9n5Vawnq0DPzfsYAZ5SbsnyBfBXbZxUksLT9a3CK8byiak4VzOok
SAd33QYcEvVqdOi61KlLP5cJ+oVyVMSrWUm9YDi6Qh7hdUPFYlOeqA8XWL+Z
JRby/6PrYn2K0wISDGIi3Lx06gAxOa2WjVkH7TgvhmGvfB3+BHJoXsAZ6PYI
QJXvFYiqr6vc2ZXZbgya4C4OP53XXznhtgsSG7MuW3SE0XgxWpXvWSy3mJSx
2cE/e7LotnurWtsXdituD3+imrNgUSoi2dbhyDGo7HMbhatS4aDrHE44QcXo
6sJXgsJKo+fS28GA9f+jN2LstOoi/pC0Jl/byuznTyFlk+nJjD/IEHT1FtFS
gaiuEURzRKybMkR5qzyRU3zyXfJuKiN1S9HGeuD3uARmYDmEOVUSLiU4K60R
5GpOtlFlm9B/fNVJaS6Cq3/yTlAmHuUITikdJ5opLMuXwHtZ8/0LAeqaacym
fWAaztX3RMParsY1R1zOqsnPFXJzziMONIt/UbMrhJFX8XPRpDASDDraD6lR
/AaIGAJs+SyjvEPBlkunpm84lk2JKos4siDF2BlJwyHLxPtGLqO23OVAWWmz
em/QIIQ9wtsW+Yox6E91NwsA9eA9XroZlUYehUZhsavATyNyNp0edx68os1o
RdD6TaNsOn8UqFZvpMGUtN8CUG1OXLxhyWp3gKqbipX7UaR9qBpXt8ZpffI7
Me46ryNatEwwTUgJfRn3sp35jHbGctndUCOOPha8GjvfKPGiPz6mxH8oLqaz
Ve2qtkyTK7cqtScIPW3jc1HSDWozFWgxhdoBwPsjixLc5Xgmrq+nWYO7MxCo
OTEcSlBVY1cmi5ScrFUsTu10sb6P2Fdv3UE0tE08D5dzKPLPWiKAUMobrnGq
kTEswppUCw8rfP3hOed8brWprZJpgfx6BDPfJLE6UdcrIUUxOqv/tUkGNEHg
7FISFXM702NNe6sUWmxtwKaSm1YTx0tSkfjjNb1zZEvoeH+HrG+ximsBoAyw
PcCtBqvcpPjgy8N53Mq2vt2GshTSpxJmdCcQBfuinKiaVPGb6Ju6CFxROyP5
UrVWnOa9eIW7qKme2QidxMPKND13CAjY09xQqeTGI+T/2GtwQ72FB0zsPkGj
T3E0Bv7KD854UcSzRA38Mcx/QoOvHIeEfDa0KSd+ZHBQJxM6T0R/hADuKw83
ynD8YPJCYDDEAc26x1MSH1ZTIdKWnV04w0nSIKfplw2n8FAwUIrJV4lXrPl+
Pj+jCi7lFQAugzEN/PZf9qxSFUMao0PEjG1pkp+EKWa0sRZP50PS4IZYLnrL
m3YIRltRA9kw/QaNZeDNHAP5L5J+YvQokQMaNbrzeuOMLe6GV8E97IA+F3Yd
GHpHEzd45H5MbDMeq2IRsdfCL9ak/obEVfKx20Rdkeqd1QMcFdyYbYN7j+Xa
yNl0oUcZEKdykxrnbucKH9jp+06WrorW7/3SHMyMz70tV3DsypAnrCwQVm9A
Wp9R3PhUOdyTyos2wGVXUiW6M/GtVV/5eKVSZ1P7BM6/dftfSGuib0UtsNdZ
MKnxDDNsxx3o7Pr9HjhQoPOMKuVmWX1II8v+LAL2kf5WpqJE0o6ucTr9J3Ch
qJxnyWaahAjIRsghu0RxQ9psx5LhxutKl8dbm86DBc2BOYUdrUwUgqmLz0y9
JLn5Rs6eLSUMSaunBEejXOD7MeHHIn8vODNZ6B7Ap+tgrRu10dwYGRoFEyHk
FXSvi4w6V7Fnbd2S4vTMfavSmekONgqyvb0k+hO/Z4I0BLmRaGulYYZNxzn7
zHFJquWqqmQ9hi8Z4JrZfp1s4IHIHK5UcM+8VslKZCnQiv25Fd9DzpHk+pKZ
CD5v4Zzk8KydpjnKLRwWmSPZjo5UnaJAJVFed4IKiNjwoKqhaY2WSf3Kky9A
Y/vTevtwI0Er5ScDVOK99o0RSJzzDQ9ieJ7DfJKWx7KzYFxPNrNtgEObUbS0
bLcAYj7sURunvG33QXIbsP/rUL5hG11sygl2sVqhaYTWTOPdFo54BbyKGeIU
WCEdhCWm1SPbrseVz1GXIIYTOZbufe6TFKm0lY/NXM6W7TgyMRwTKDnJ6Ktn
Qdu6UFZJDCJiOjTl/CtDr/6DDYRfTaxU3V/iIVtCsjXmM9uWPqSQ5wwNqltW
PBD8T9MoOD0LbKjMl8pwjoNY6kpxcCD6tHcgR3DEvfbzg/pymfASx10Q7hVn
rIWe0w8VfSbIwHuJFKq8+x8WHLqIqeSF4BhMZQTuNK+tnyVkOW7uMmsSlzhM
jdtxXpiPK8Guhg3n4ny3QnqDfyDL1gqcIIQHxCFHQUlli9hgWg/JWZY4DqJz
etzZ7hqEH8us/gVk+1liHwZe90nCKkM8x5UrOxKuOjIaOnDZFFQC0hKC2q9Y
WZKrSLWGKJQFMO39vaWCHr1XShZQzLeo2gNYifMT0rmHfBovDyATGtIsN97s
hw9pofQiKJYMpmlsUdfgzYm4M92C0XKg1OIweP0Zgwb2mlOJaHSzpqlGsg4i
5Cz0qg4f8NR1KswC9Vpmpjw9mWy0E4t+VRPq2Frh/ERGErCvQx9H2Pskj/Wy
gDCGVLxkg3YQDWY7a9suRMpk/PbIHsrfv5BBpo5TRjmyGuEi5ytYxg8/wE2j
FDARumsgBo7Qy2iaBHqW1V6eBAbEvrue9vo5bykgy1M8qUNl/UfvyVgOPPu6
034Wv8n0BCkYitmftnmimjy1+tVCX+JvXgJ2tHR02X94UNIntbE0skd/csO2
4zujPgmkDm4OPS6a+OIfjYf4yt2Ryte98a5rGWViThNJI10arrzT2b9D/WXW
cE6x7O97WSaL/QK2LZW/qmavXVXeA2ovayIhzUDzNh1iikwC4EYvhI3RFc5i
++5CFM0fIejNXgzZhosOyxHl6aPQJ59O2x7lH5mJGm1BPK59mRUMORNnZ6fI
Fj4XmBOAB/QLOsGFkQ8nxaVjOTB733pm0SufjtcAmK62LhUpkO0PJz8OPwoQ
dEwunwvAFRl3u8MkFLUkERxUz8zUAZw/OnK6Xfo/J2ymF5Bzt75La3zQkHRx
65rGRngUpTTi/+w/X6kTYtLoSCr9D3jlEz6AjdfiSiFd1Qv5wKSkZLRtiqU5
1YrWrVzwHi90y26A5rulQswHSlDRhHUMgQSrlPnvtfsa93Xg62Q99w1ddVrJ
Fe/T5EqvCOCFr0EieA2TRUvCAejEM6uN041A4DOjp2yu1ZghuXGd3135KjHP
BeEndxklcsSBRtEzc0kiVZQrVwtSoFqcAjyptZG3RNhW8LQQxn3rsURZ6g/z
Z+WuKmEBacrr5kHSrII//SGiakq0rCQa3kauLkyPY4xBthFnFbCZCQIshIck
bpckdU4bjUhBpiV8m+9ym9t4YoY/Dh5pfBLUOAyNFu7S52j2WB/QEaZG0vhf
HPxtTQruwlItEVrA+TH4gJsY41NDvwnU9O7askxH552meVM4VKFaHwV0QgKW
+AuU7DxI2qnAGMpGZUoMXN2UAgBLrvzXQW8WwQXLjWSvp7k3IMOPiIsvSyak
dZ5wec5wgAyU0OKVFVZXqV3wpBbtsG//fINP+IDwG5Kos/hRCuJD+VjXC4u6
GdFPvg3SAMYTtk+konIwi5SqnOB0Fr2DHViO4kDCPuFwlij1bu0qble+iw39
i73G9M9/YA+EN2OaAWHQcPyVwW+VbWjO0NCc9NccFSZQ/7Slr1SP3In5KOTr
9C3Jh4dYGu9FRneUhqXvWRrAhMBfETdG4BobVoRIpwi+IXrfIDP7UPci+rKA
vR+83PjQagOzlJM3wawUAP2ERT6tK9r0VpxoJ1AiA15YT95t7Xw7lv/MuAXy
DTcHjVBMmqrLb7qjqwRx2UXJ7aHhcdfRaF6QT5TFKHoD9+NWcsrh68ryZ/H0
kYmQiZlNxYeNqJGzcgnGxThh779ukeOuNoZtGaX/6Mgv8liUGtVwjNbF6NuD
sFkYnUNZh9lnfmO27fVkh07aBrypvif621K5JCh/jFnOHHs5WYtieCTMbSVR
XLNY/CMtGbDkTmB+HK7b7Hfj9YZW5ygdFthZsQyH3Tclmqp+ZJV3ymAN/Bv6
31I2hxxr8tWLBr6jZaugnHEmD5rF6avwSCm0aw5yt+9cNjI0c6vsPl16UQxD
94JXbVSZJq2kfNS2afMFWCQMWDeceHcp8E8ZDPaXRhY496G9dxedUWoW4Qc+
dZ3hUwwNbl9EYn2CPrcE4QYYMAdfW8CoJexxTcu6GifhNvI1SF2cCe3TUPqz
EctuGxxL2dM8djkbC7k0LllFrt07PuH7mxPWjEaSBiUfGI6xS1xAuknTkAji
sR6NCdfCqaYoE56phwgTPhnbbSe/iGEMdxDNFssh9OzHA4+pQsEFIsgfr8BO
fFh+Z6+MrCG5u0Gp1PBAsyOJp9Yk642Bq+vr5OAVEoKWW+HbWWL7yVijWCv1
TYdcgT/WX6CDTtcRb5hfBd7dBlgMEhZaf8LYvSxzZj8eCTBfNRKLS7eQ/lWl
fi/Qj0Z5/nUp5RrYWzOdwl8FGfSj4MZqbEHGkPIG42kIXDo8fjrPXkqwc6UM
5ourRiwQFc2/TyxhFK+uDkcsRtljbc7K79579drrQRRgKK5OfJw9WzIaKuNH
KlFFd+EhifNqoG2UootMdPVfQIAFUE38VuCa0ahFuRQjaZAEu9ufiBpt2MyC
5oqsTm7EDsooX1qRjBh3NSLWLm9CCSuNbKS28Oskrs2shnQaX8RVSPNlpDUZ
xOXwvm6tbGkDs/WboIVdH0sD4074FLpBQyUhh812quE6hRlv66G5INfvCazL
O3+ylBiDcZ7zYpVqMzF1ZmhppSt1zKi+36Jc5rXyawt+qP4pP5+uX8xVH3cY
rjmyAIeU504FrcJKSfQGwz1hq/H9tBQWaAkM9ju79q9B8xNQOiira9Z6sK+Q
jYRDYlHNHH5q1B4TeQRjLbvWhQ0NbZBIQ5ceuceWn5kwo/GaO0pXAu+YFIY6
5d4dfonlNJh0IFYwpVbEcUs1hRng/Uimq8mrspFYMdQXe1phfJIXXLKg203d
8Nr2Sb6acD4h08d5dLw9GHVMa87D29s6rouUoYmLqlKUIIbltnAZv5bB7k9S
ocWIid/iGZK1HhaOmDOhv9b1jkLQngorncQATvcRUfusz/Moao9xaq2TfG0L
mdyxrKC6gbvLtGS7ebMiwqqyqLRvZJWyqao67Z9OvQnJhwE1zjm1IeiupIGO
sR8/scc94fpiiaxbqMxRdcViEv2Khr8ul46CaRNAmsqdyfSiWVUvE/lwYSn+
CY1ochGEwpuC95gLR+2QUI1+zQBJec7pHGUFOZpnC1JZwy44agJn3XzvNc5m
6o8Bc40NJy32gX7cZ6XFv0k7mbrD+EjaFz+9PIQmitz/VRwOmHNhNIAIW2k1
3vjiTMW0CnVVUVE4ovymxFHO4213dViWuVg5bUgLzaJvA9x71qzmdOi1SF2+
vTipGDvyl8YNdxXYPG1POGSSFD1GTgjSpaGoRwa9cTKJ5J/HBqeuVvyGsXoC
Pexiyq2YPZTn70M/0TOjz89nblcEZaHtUsm1ZEj4ymRCJSbadjye9CO8f33m
N5oeAPGmyNqIHnaTOmc3LKF6FlX/KjpCtAH/auyZGmIdDS9kXoZZ/+X8lZD5
oEJAUK893Iu1478oBy/ybshHkioBq5QtX2/8ognc3O0A/kaviLuuM+EdMSiq
8Cr4O1DKbyFe8x9JJ8v2EP1/gdeIkuT73LTL/LbcJMf8vqLj6jJLYB5AZeZZ
XIHk0n0aB+JYm9YQRZAkPn80K5aedQJPfWy9WzJ6rCBGKxKW0PcVFNj4AMCv
x7PaGJT9HREa7UyrCWmr7ScKK2+3z6DNXr/JRoUvUvMcaNdgNvMONeIQh35h
s7FNpZVcVVBLZQmpuuBrPZPS3Zk6aZUuvKGB2g4RPPKx/wusP6iVnEDRgBhI
7hpe1BeTgwv2REzLsVsaDaGX+TYRPSXG9/iWeeWNTX5xb7PJnsv5T6Jf/fnp
OKptqnm2i/Vq/Dzd1QLfGen4hQ4tB6IPlzvqTi4oFZXwxW7DItkLWE4zE45V
HSOX/IyYtpp13Fl9CGztHOQ8LhKecE4D97v9r8inpcoaNnECCckZZjTxL5Xw
ya2TmIu89kleNARy+8j2GmDa+CZbu4FL+/S2xmWAho4r/WeXPrY2qEe827vm
Jequ2S6q8dLtwVIX38Az90pc+El4XbGH0sEb4WlzOvD7BUZlr+bTWjSDOZQ+
pjiYo91LqP3A3pC01yOOHjdQcl2tJ7lsnxPuwm3Xw18PKnnStemJOi0SfPIy
58xgv9jKwKkKqYNXOIp2VP7KrPSREm9fqgYRk6EO8TU6rwjhAfv5RF0GIT9D
cQ+VTkKUX9aEWisPyqa9Ah98eaLQYSK23jAuDpGJqV3Jv2KMRMcObiVKNI5E
EeSgFE7lsjtZxZh8EPNRsdvfv9MuEj470baXCqaXekA5gAoHQMBYH8KWGFxm
xam9wk45aD6FmKUE5fW3E2OMbZDUVgzdM4RceoblwxuQx2R75tGB3pCizOOt
jL2UTVpLxe/zts6jgbzGlPJOI5hyRT8c2Q1cFxW6EIkCCSv942tFyiis5LX6
23HbS6YNIwkybqUj6lDohQ/jTUPrSnczWZtw/Lgby97Lf1lFF1nTVTCS27TB
1tbcbCxWtvsWegV1Rc6IbAhbTt/UYTB9y98eyHb6coTdvarMH74tuj5yX3fm
2BsX1pKCvl4fSmcdknsgW5iaWUxe9PJ8Nnm++0Nl4HVAyjXNWaBKHwkw7K0b
pKlHHkutP4EzeVwVzgXP0j2D6F7S8Uiyv7XLR3wGgCSYfafsrdpIW1BcSfsO
IBcKYcfWvnaN845k8OWmVmzgRQF5WXymr+qfS58k8rajrbMsL8rCjbhVc2gX
KUetIUBX49///npNvYZtysdf6gSnNqnntMSgXAecRrs2Gme5QMcJEwYci5kx
cLYg9feI8sePtdxSUB2E4IhcG3M2nhRy7/BKaemWZ9wb4HefCfFY2DhcMSPK
R8rrdnHl8T8XBRaWOz7F9S/zaRr6c7IgihVMMOb53XZaCkKCNS+OnmiPAbgF
51fvpMJ6rD+oarNH4qS2iRoQss4L5YLY544RJFaG86KUYpc6ISK2HMfgRL/N
YXFi4QJh/hjwULbEeET3XIejhv8A1ukViRUXSwoF6NqO89ZGKiUHPt3Mwrfx
VPUjuc+Z8c8wHJ3bnEAgj8qlQDEOtRW/r6xFe/wrXxzAiyTk20yJ2YVDUd49
K/5In7ociBFulmCAMHEGJITAutYrFm1cDycDcB2gcFBEbD8h6871f7bNtMGI
Mm0D/T3+iHSSzkvdWyrA5kNyrQPBxViXn8l0VodbcX/QRVgsqT2PBcUjFc93
WNCztVxWNsT+0V6qg4QCQFv442P4bEovmlww345TziQ7VJ3y56fq5ooWoiPc
cjXEohEpO1BE+7vXjJfpPoolQ64k8/v3zD7Zvp+Km6SKxHCnnBpVl5a3NWch
smliFdz+yGq1HUhVQ35QEkrKUXrjIqRPDBItkdrvXHY6v4aIjjZf0M5yyhGz
Nge2L+riiSLGGfgxYwzRAlnmG/meGA6/ReMlf4nwsiHvyR1aTefMNlc5JnpX
ENEeMT45vfHxar2MIuUfQPbjBx2niRnmLk4fBKMsRAUs3E0z7LSpL/KsLP7n
D6Dfs2a5w8lm9ijhgxz82DZfhg/ET1wRfMxiciNJbmJilutfV/wJD7XkkhnV
NzaHVM/XNWi8UXu2t7jqgVwnFpjkV3IA22shgQ3CpwlOQ2dxtSdKzGoM1pWW
iB8sAh9RG50SrdnqviFacl+ksuD4newwp/geJ1jx9sLUrMTq3UtiYg6Oe1rG
V3hhPfUzuTBOb1ZdRAu0/vpocUUK0FTB5KYbYQhscvpqZ0ax2e6qbzeyzAF2
Jq4ucsIeD3dQAd9YAC/lg7T0bZLr/BVghNw4KKE94i2sJmYn8j4KZJDtBa5o
yExj0nkUE0tVO1BGzlkeN88f4FxM+xtazH6EBxE6r2iIkNz2VyjQWD1JcfBm
/uH4C3AWB1/9cns2Fan+9caipDsqy8fAwv/Xzi+oBOIlUhQmb2VKHrpLfuqX
y2GEY5n5F7TJ3wiYmJFOQj7CZgDT1cx6tlKGhe9TciXwhbA8tz39ZHoFTa1I
Unl9FpoOgKV749XSS+sqVvNmtr+RRNF0l6K26eR2LH/3AIg7MOQmRhCtNTju
kztQReSCndBloYcZ13Ec3e3Ric1vpSpqifmR+9C2HmS4KcUoHCy1XcYA3WdH
3nZMwOZvC1lMiVpLsaBiPUWEEqo5KepBoiz0mpwYyuaXfhbDBKQz/koBlLDY
dUS6XAGh3rAWUZQxszF49Ig8bxV+NYMF/qLM4DWERP6thEUNqXNHNMB1upWB
qjdU0kIGMOUbIjDjNeYPq+CzPMM+o3CttRKU3ngYElAlfvJtrqIz7XA/8JNM
3Xi1yGdU/TehasrJsgSyXN2RKjgmHOTH++E/1iOd4u+rZiG0xeseNvLT12kI
fANml2om8KcQ6JgeJTvRUUrOdtntvJQ7XdoOwqHNS+fCdXlUfSSQ2KfEohUK
bX0l9PttWXVSJPXQaETl2BneCQP9zJP3Y1XYAf3sTnvKjDpawWazAeb9Vaa2
cqVs2chUoDZKNAy0vmlP+bN+9MV1fdbSvcuwBxifgY9ujMlsRmqJkFrDMzVU
Y1VJjs9PfPWWeRvIzrFcwWz+A5vGWGPnmY2XVOv2/biNefTEtJH+xNpF277z
79qOZXvXL+ZldEkhOHFHMq2AqrQhSElUGbRv2Btb2B1Hpf6os6OYQ55Zxb+R
fCNR7REsLC31YQX1Sm4EkRcvHcBl3H97a4E4NAlhIxRyah53cflv+wb6saAl
qoZ8igX/GIiMkYGGA0634GFJdGSBErgVsmFh65IJhIkR8zj8PzcET5a0jizH
xMLVxqPyshYBm47JqNg3rYdH3P0fNKSoPc+byQdIJG8XEGg9TEWJl3V9BIii
HArij0kVRYYBIsWeEpzNWYeaAjapp2V/rVhaMaqTKu9KDP5RqO574s9nOcP8
Nd6CmVeTXy7xl6/546eVuC088B35rcOoW5uoqXMsTGTxxUAFj3GNDA3LSZXy
OBkT8ybXTP0dzdlKc1e3/dj5aKaQYleS/OWPU6TRtaggpQOX2eeMMAEanWDW
JbVp5sptS3+SSo+QqZqDXnF3ePQf8eTFnt3CF8mt6PF8YxRwIbYEZkBorC1m
NMQtXAKMXqDy04bOEnW/+BLjf/ODZMePFNDQw06dyT9onOvgdHo9DCJ4VAKL
2N8fuDTIzHvXzwxRM1DZscc/fO2WCUK0hd+ofN0lgXdYCEU6hCg1mB9hhTp1
ntB7RkmouLhk04VgiF0Xp48yIu4EniCsIdv56z9J0V3fBnUmUAPPcFQKiZn6
q2RRTiTl3HIcoQg6ByF/2ZML26x+00nvcW/85MVL284b/Xx1xTwyJWD5iA6S
6iTxLkQronvjd+lVt2QnMRSnc9Idj6BmeC6L4bdrZBh7YD6iYD21TF3860Ah
9CExTcN09F+ccftPF6kDi5aVpKlrxC/NfJ3W/HDnc86CU9cqbC7NJlecrGOG
Wnoagf5VnUcdB/OV2VbpdFdjMq8CBvx57CaiM+eyuyJujNAcw8tKQCrcDwQ+
tZh5wflQckzCXfcvwnLHC1jbpXbMQP3sjWVQIUIwk6E5XarEZ8oxHJnokGkt
qb8qCRbMIJpTlci6WNWKohZfaUO774jzF7ImwKlzuu2/jKjXXopl4pyKax9i
aKLq+ywfM2jKx0DZlb6m1DwTz2X25JmA0TLtlx8pLywkBiOSn6KaN0nh6KSD
K1sVDm9w+didKpBoPSZwY8r+lRKoTK1qXKAYZqvXj+V/WIgGpXFUx+88i+Mi
FEfbkiyG2y5mXKuQAH98qa+D23z/KxaO8Jun/7f/faXNL4jzRzkEqbRBv2Bf
aTtNw5Zsli0S8XF0D4oT++58ZXLj0VrJvPSzDi2/03ip2jZcurkXjolxzN/T
wWLH9NVBknyXbn8vlrzsZ4dMksOBHIn+0UXS5iEG5TXDItnX8UP7P2Th/sZh
xi3qDgUvJpA+II5thQRgDxr0yOhjYlPShMS4zA0KH0vTzbPg8y/Rkt37I6yf
4GnWmgWTcbHJ4FxXrJLdiK3wSGmgeYE8ZZE05aFcCd62A8JaI9e3Xjfht2pH
0MDlISW0V/w9lWew7eYPWTq/8pd772vXuElcZRMrFFI5p2A1rUYsyd4V7h58
JDdG6s4GRS3HvriUuNB7hKqlccYoQRA1uP4V7Hi4MuT6LaSFc7EJZHoVVTbo
0xl+WmoA7Ql7IQf4nan4+2omla+Ptth21pEIAZvUG9yYyArTpVYD3V6DXF0E
YaUD3wEppNeiKLy9UErQGd8ofimlG/+sqWyuqV30UZjpb0eliytQzU9KklK6
SMDft7Q1h7r4RaFehgDNOEupyOa/9rjBqRf2/f4FvEt5fIv8gZtMpZeKi1r3
fZD3NoO4EJ4jA8doFhcTFo+nrHTHmAhk+IGb0B0+Qz6igDgxhBaigl42Cvol
/OjOUL/SFOR41fFOvZYWTgMfWglL+4tX/6qZskAYCD7M6Ove5vBl6K/34jNN
X+o9PnimS6jSuKzREBht2knugDfhfb0GVnr3K5T8a4gG996Q6hO3Bi1gTnBM
nmKgh1iijZZVSzYbS466I0F0fsSY1HDj5LK0eO70jNMD1FMLTYBR9ITFvQeu
51RbHTbO7jjSIiFXTjnGntIGGySa5XJrjeBa3QaQg90euZcuAx/OjaXk0RLY
wLA0mIBYGFuHmar7f8nnndKtrWgCJ8N8eAgwl4mkZhD6l5d4ppxt2R4EtKsW
QlVmii3zSLJcU0Viqa6Z9GwYCm+HA3u4h34Dec27Dhkj3TMuwyP27KV6u/Kl
4q/gDtXBFG+rtXl/l29hagTzPXrBFnBvK8FVw928vIIpkk4F40WxyFssxeCX
vHb/d6G+IGQ1Zh60bL0L57uD0w04cYsjh4XW9DwMgx5alDJ6ZtTMQ0vfGIUS
xRhzH/FYGlvxqMufgLCZxS/iXDfv1Ct2pxqDWapjDF1plkyhupcnw56ilb3N
aJX/RQF0wZuYaMl4F1hSjygIhCd6C6Y+gSakRRnTVAsST6qDjCWEXVy3eBxu
vak/seKwxYGhU7u+SGaZd58kvg1zJfZSID/CE+Uk69Y6x7ZSTJD2M/IS5P6a
7UkBmRjmo5p/6ZlVRVksoSeUqeaoUBic/o9hVRQHeXUu91XwQOLV8zS2oRAw
rzj8uIL5UP47dS83ddJjb0aj6/siZkGKzCWQ1VCF56Uo/X1K7GZHewhInQg6
OSZFJsMyo7dFxsoDXtQSXQ1DP6JG1K6Dpb+QbYfzaYoE4J2jcUUqFMBJcUkk
+pAH7nY6zlO3l3bL8cgV4YyOmhdN2ET/4Fktpa9x17j2OAQ+f+GxnkER7FFZ
aByciYFZfV8GLJlqZlGAwNkLDtvxJ2GQf2jtamQvfY933G3KOHWuJbuOvhhO
VzxJSH1RhlE/SZnD3R6ba0CIywQyk7dIj1zjhrMM2nudS8y4dlc5mBQegu3O
CtROBK7WPxAtm5DKOR2xtHIltQ8ohqENJyixxoksmKV0TskOkjYxVW6HHjjN
SoO0oQCyojntcvTJxTphQoCGPtUYqf4dBZHpp/jxK/UaCSfgTp6UzBB3KVRN
6lTSZdgLz0YKDGDO9/ke8iY2i6WxFtf/zLOkeu+wn2d7VFckdcCflZYoKTRv
HF3prueRp6NTfmKRCkqbM5n6Yn8kQICjWXPpAh7gOcn1/EWz161pBTJ/PNsG
jEt2/9ModZVgV/dSWqf+G3WdlIt/l2ZKrQhrKxJ8GzGogm1jRtc1p3BY4oOv
QSXTb9c+ilxmI6wn2oHl417OzviTUPFwp2IeG9zCQXeA9CN9tGSbx2R+cG7y
gZMWPx5tGXM5qtv5dtp+XIcB2Q/X+WOVFZhMW97Rd94WSgY/Efutzp6MjV+u
ykHIBj3TJcY7mnVP5OEEjmsn24KV2uyLPx+tM06qvARdPwDVBNdT1dFqETkl
PdpGQ1H7L/W8IaD/AhSpi5HSEVtsap+iGnxLwkmxOgfS+Gv1QraxFaEKCJMv
Pd5jySsyjjBjDubHkk5V2/uR5IKCgK9JexV72/rlifpLTsxn9iC94eMBwqBW
lh7eM3WlFgj7u28S2hrY7ToOcoJ6/fJEBAM43VgmedM8NcMNUPOrtRX0Uz1S
dcfRrx5bjteYnxaas6XiiuzRA+Rqhak6wqL/NDCz6h+VLRFSL6MzcJ9Edk8I
CtTW93rO38kGLfsmTWfEmE9zghN9ETkAtgQ6+TSdAOp3P6pxirGnvZPo70ev
SE68WA4t5UlMMRn1SkkIPSC8dOJdrJHaE1//l6ipDy47lngn8J9JwzCMz/20
wyQKDbA6D4AhO8/SaIE0tz9munY3Ukgq4NCKkVkSEcssZ2TcPSgifmW31xVA
B43hQIUsQ9MpT790WJsrX1kHep+9ICIpH6skSLQp30Eg+z8t6RxkB4weAfnN
V17WvtUGslIAAdUEN6vB459uMQPGUik0qUYyyC+4Slal6AeH57VbhqHhxRjs
AecaLfIx3FM6w3TFdYPGfDMpUH33uiMocPP+1/m0E/q+jhfctgadvAKpXMgd
V9EJA5MTwa8D/GtfoiQdD/4AtfqKoRq6FSjZWNd1qOtW4QlMFxUgqWPg9VYD
hWY0730Zo2mqAij3H11RtsiJbTAd3BCpvwxRgnO6b+u/Du8Kr4b4AZ4tUZxr
O1p8T1xaxvJbszP7Lnu2akYlv48qb+P2MjNUYgmnJtXopJcnU5+MTpIYebUC
u5RAKZwpj0sjEDF+lrN3DIjLjk2xesH098p3bKoST5vXC0oqNsX4LxgojFd6
x+jCCZV3dstzZCm5SF5ZGZl6mwvcU5ORfD3eQRghJSDSxiBpesh6nrh/Uogt
f9rbfr0AfPKXi3B38AvRvLaYR56p8FGHZkvXHd7qxp8k6RZQrmAjfAe8kn3f
C/Zk1kHezlDLMWCOLUiHMxSXdqMyLuA0YCg5WOX54V2HQOGsitppqWj8vx0s
HIg6uflJIL2TO2O57eelUFHFisqBvWgqWqHgIkfxy6YUOrvsvOB4APBuM00+
sYJLki8060Q9ipktKLWA8JbcDg9uDl8SqyKqTGk12HXVmP+ZlDNUsy2XUe3a
uiQyRJycImTtXGaY/naWtGzxRZmrNS8XqTWCL+JI+bjnUNsEzo7mFArifAxK
D2lhd2vjJyVibylGU4Nars1osjI07f5g1AcUQzHg46D0KIF4v+nuqHb+Lh1W
r1GwnZqFc7qemmzWAI3zQpSzuWrrzXkIl5oLLnQytGKkU9DjEQR+N6V/Ivnd
7m71PsKsq/6GkhKM9jmrmZLsKXvxXBDU+ykUiQgKRkDosmGHxvvLTngb8nJJ
8iLNTE34ctogINIwpVXQmxcFvs/dEn2YkA1Ng44G3tQvJ3652VpbQrshx3jO
stm/7pYLqErgvff1+HNRB9zwDvLSgjz0C/Tqxc+rO69QvtkjTiGxYb8dahSn
hqlqfFivxo7Vro8apYSTX/qV3upTbpafUWilt6C+ziu6V3P8Xx0y0CPuqnqv
B87dH5EvFip/Xo+PgKm/dkFZa/N9WpnwathMjsNMnO/hHrN4tqwr9ATwWU2y
tM1cErcvmGwbPWspj0+I5n806Jo85N3nsZPsxCv21ArVJlcwqSgGft+gyOX9
L2EtsCC/NFARsY+osLLvTYCcURbYPPAWtuguPFzdM1E/9luEwPS3TcIN+sVw
ucPMIAfG9uMtS8O0pIdskkmUKa8713BnQtuvsJtvMGxDoJN3UN6/KNvgDaQu
zoUrMB/B8YE0K1yRMMm7uEPIUAaqq2bbzOAQw7FCKzoAEdyypWTxOvYk5EDv
hqH7M1Rl6acPAlVqQHhUKgfqz+WbD5+zUjY+u3oEiJdSmH5cBV+NJWdhYqvR
gc9u/VspnOw3CtvEmW7+t6HxC0CLaKBi3cpdy7K94xIs8Kh1QsYoiwjlTG2U
9QqlAjrKVpq/oc1pNuTzt2kxp1dTKM5RUZ/6RElpYKBQBADzzEsA1o0eaQHs
4zKr/tzeIlfbIq0ERHgVN5M4K4DZRICL+Ytq0Q1dqQgLVNk15uqEGEebONmm
NX63955phPvIrRQw0GPBGoDqHE4w/xOxz6xtijTeLEHvtW27/v5qelhZ5vEM
rbAskgULY93zaL8BDRr5hrYfkS4li4PmfacZ8nvx3ReXmtTVqiwTRx9CBERS
3N4YPvCrrYSDo8gSxovaqURbMUaDj7IN6HkXcKJPX3xi25uT2osJGFQdnW0D
H2gShf7+IvFkmO+nyuwD7bzKd6l9vNr2w1/7wr22rAEQTFD/RfwmppACuX4e
XPf2se8Hi5D64rmtAqSW+q20tBEP+dKpjOfeqB8mOaJpzQkyo6HdGif0uzZT
za5+DmhFunrd4YnqHfTMdj3CFVK4ZV1cXvkKJ4ylmfIa8dEwThgbgKp4qHKh
xvwSgr173dT/i+c4lImdHPNqLP9mcDFgZL3GhkbzbABgThKL0Vm4ASW5itL9
hLoPNHVoiTI87V7IGX1uVLRAg8wI3xnY+JNncswWr0wrnsWV7BgFArydqPPd
ROSmmSjSGBqgJEvJq1Pvu2f4+Gio3OXKOlPcS7mLmEUhGaSsxf1qwffxmeh3
Flkwk3b2dw5Qj06mIZ5kXwb0HN06C0gtsFFzr0to6bx1d/Rn8fkOHAx4Tg4F
FTDTN4bsNuC1/a1nyByqgCPQJc2zdtpJq7RkcTZK81muSfTqBuPt3Mbeghf0
cNkMQcnLv1p9a68yK0qAxI+i3h7zEEqWA+D458E/6OrSwbyWFERTPoeN7zwO
SZNvTjIth2M8WGSdgs0D4kAvvNORwPLLQ4kLXWqLTDxMc+kSKqjVCRGa2b/a
WgP9fHOmYJcgGObVaEEVfs9Q5e6HBwv/x7yd7eN7vNPj0e4UjDCHrbPmGQgF
KWyJCOIrgxKeCE97B3HIWIcb5JG9idIM+zfqdQIpWFOaaFAJqz3WdtX7y+XX
lVIAJMGr83jnSl2rYAAgUwSc3GTlYsAlmwlCBfPzETsK3PcjDPAt2uXsLtkh
Fv9SC63BUQwXaFjs8JaEc1Wigbbty9yFsXwMW9yipPCWpPpBCE3TnXLoLl0o
orWdgOUW3JD8n4jpXqlaTuewf3Q1dvFZspzQfClT9oq7AlxtRMK3MKQ3hb47
YU0ang9wqpUnplA1T76nCNZ4ImF6oQfAwjpfuhNLc2VXH6Y8CySlyPpWIISG
ji16UpxSWoXaDn0+da08LHzWP8xvo2ovMngSUxnRbb2tWI9EXIdOiJxjE2qx
b2SghvzqFG8pmaH/ZKdiMz/E7Fk8VbMwlrnNBhpbXUtmNW/hvfqL5GwAal/Z
/9f5uAZmHZpoNXRURNVptPBSkRYx53phOqA3kRhq5G5HXXEPPDxVA3qefdr8
YsOCSePlPRNin4DOtbztHHwPox5edaGBg+fashD7BckAZJkv4lrFqT/mP4PZ
/tLeD3m4JFKIIzfW3rdD+yYHfwFECUzMvV9zulgrFdUBLvWLxA5mNrn2itNy
WYKapCFFxPVzG0MeW8aPlp4pnQAhd3RyvhFDtp7p+DorSrs2DxkUx6Fuw+AT
sxrGp5jRIIkiqV5/1JS1t0x9oHiRSTAJY5QHzLB0oq6qw19BnvpUyNiCiU+k
wPRXXFdySIqn7rJozn7zNz8IrJgAA2p2OHeqQIXhZ389gTrbvTQWRxWsiNDL
MykjqojKcX+Zm6n8h89LIAo7Mleo0Qr711oeHrHQF9RzQRiTXIsv4WIy1ZWL
2kcgFNq4ihs6rOXH2CE/af2NE+CmWhR2LectxL3lEJvWvg5ZCB/vlKqk8RXI
dyNs1lpPgs2UJ/cjxKhZrp4oZsSn0kEM1ybI0reSjFmDouaZpJjir0PrB0Ga
YyjLA5IqThiARvCdEwbyFfx2pIIKNAKXNaZB5IGGlVD9lfhkyxnwc43ygluG
d2F0w7kawwVryK/tTPzLuwB6NRUf0j6MBmuLeS5Zk+VGqmB//caQ2sg6udZZ
a1AzwJ169oSvee2qfMTB1V+yRzoDglIMH2mNzMuEoNTYPMr+iYT8vWe3FNNj
kmKUBtom+65LGwFCiydZ0JVgWx/ofwdx31OIJLx0PZaUiNT7+4jAEDRMFMP2
bpXXL9WfM0fyk11i3mAA2OCfn8G771ZEFdD/+g0WENjKXN/IukIelMaAd43u
Xmw4LV95r1tJa5h+S/sZnVUH9+pHg9I+rDvKPzIX3JaSzaXWPFpW1D81s44+
SQJwkdIuSj5DeSrbOSTGwGKXewAVpCTUqKTcS06JlEWgE6oH62lx4T8JqExx
aaBux/0SqXhp/ZnxbqCOtCsPR7ZdrCWlrHyqXszaBJdeZm7ZMRJwNxqfxQ6k
oeKNYBahgkZPHVxnkZa+r13xP7S2s+tqtKfg0sUxpkVC3ASjLuZw+56RzJ3O
cF2ZyEX1oJzvQzmTrBDi/6BzivAuJHwySxmrs/T3nd9dP1OBm3XUAJdtKJOg
T8ke3Uc/1+WkHQbhClrU9IHGmAwXCrhH+21LXCwUUldTa1qesZvuH4Yf/vzg
d5KSwr4R7yWMTdtpai6WVPKyrWbUOUlqiuJFEjXOIMnLCFrcVyVHfonb0AYN
bZWRDPjFdUyisQbXjPnqorE8ssMHSUqFvURKZWNwDEEvLmBO32HWwdw5XDmq
2/gOgeAJAF+EoViqctvzTl0b3SKp6Ns62CMsT7rJzcuEkt1hDfq4o1aTtSWP
DTbVukPbQ0QBxPUnuJfd7l86koVos/IzIiUQy2TvSyyZNOgkWa3QlE7R3AXe
T1lHkfMR065b0ujeqJDgcNCMfYBE42bYQwz0lYkcjKlOITfixRtNh/YB0ZLM
xPmg4xzBGwGRNuOpLV0zeOtvAVWADqNcJjXNy7OkyxXPO9LnMitU8//YDqBU
um5H+b4Sxi9HxsMYD6CP5Ml3xZX8gUSRHI51a5NxigiBxWY2ZuPeIVMI7BST
+3nGEVU3PQPZb/5tH7mEvOmEraBwVBipvOtjH/usT0wcjmxEOpmD2Rm+3QR7
hC/otMqlJsv/TP3h/CGOrNuV2N3jMhSXixMHHapQVBS+++omZazc0nfaF0J1
3CgwzB8Hh39hpkm0FRl1w7Wwx/4J9fKxefT/Ex6JxohXXbgGz29bC1JNNzjm
ZSoHzAg3iRZ++g+vTgp0iA2TdCsagBMYLUHDDiytvLaVdFC+IOAK/2BSOS7y
k3XT/AWchbxbQbq2C/4Reg7qufKPuaIbzM02C7xdbC9PPfKpAiYC0TdtgZ0Q
4QVnO1oUuhtFVlBeO25zyb4hCCB+WLe95C0bjSDXAKQHBG6Bk+USsrQqQ4hw
vfoodQOe3kW5brvtxuxk1CLv0qUUWCBsDt8M7VbiemD5y2OlknlTq65wtNBu
DrI7RlUD1vZVLnNQwDFSLWsKr9Ey4apLHdwC157Qhoa3b3qlBKL43S2PtQaf
lml+g/RbqJ+7sNpRdeD760tNmO7c5f+Kl7L5UZEmBIeQU65glLTO9+y8Kxan
djI1PcjwTZuAHNIii8smpTHDyca0c45naAwMIS26+rxDkCIWzTA0TW4nBsyI
qAhbaCHA9rlLFBI5SoGMo4OvuSQsTBYYVltWK0D08pxMB3VaS7WGFdwYfCGl
eNA/YA7CQ+WEsY1uSN3jvWGKEEcm98vG4jk5gjIup6vQvsd1xkTl/l8p48xs
GftiQblP3zJKKTgE7INVNxWXn6//Vej5dWlQ+DK+2fRmGnH4DQ4OE3E7jivM
GhXk4+LuVoiPBDzG3mEOD+a+o5NzpLG9sP20pQyzEaYhVrLuPtVQMz0eg0hZ
HIVnRPwVaogLtInc/R5iKacad+W2N7nYA6s83RCUfpY+cbcnoVbJiYELmCjM
Jab8KbuEM8aL8nZv+4qp5P0RB5cet61m+hyQAjIkU8LKzIp1VwJkSu93CZt9
9NCJF16U8N0BlfFpjy/ZcZ1ZwnXtTvHhLzI8jAXcpr/wdt1mNLIL3A/KTtWb
8Do2S8zDX8nUuB4yTUNh+NJ9jeLSbZeRes56z/oYErfe2DqvBfa8BQHsMbX1
qDFvHmOI70vVhLy/QZpod7tHxzBA/h4zYSaqOx7kerEKL2MQ34dPOhy94/IT
aekeC8GD1a+fDS7bQT5Fa5RcbmuLkYXPaXpYqRLdQy65LQb2kkWq5BLYoMJI
wDwDr4JppXER7i/fMh1N7AomgVsrOdf8DRQf9q5yzrCCpmBKSZiyJVcpneHq
yMoPbOwv0n45aLMJ0uLvlQtWooe+gls6Dsw/XiejY//uULX8oHJ+D7kEMlsJ
uDKNogU96v1ebevZleAvC+53ejR5ijIknXH5mhsi2xPam2JYdW7k6U1IXLBy
pxF/u8yRhJ/PCOKJU4BoFq23xGjspFBGqsrZ2jADvGfjRmDkZ+tqTBmlD27k
MictYu8EwT++NAR9c4PMxcH1UeF6Euw7PmPMLLSifpTDQ4aLnDCx1Ugs4w1t
F8ZQs7BbumCn+6NWkO3AJQyvs0AKQoa+Dvw/Dj/J2WYHOInPrFd0pL22ii3D
/+x5L5UnZf453PZ28YcVApFgjjeQb5HLP3mkCCEUj4ouxCmIGoUiQUH+Z7x6
xkFLeQe3juwA/Fpto+7tP8lfvkvC9uO+1gT3H9OaDwrTN/rFDrKaikfZpGiN
klYZBl0S1+1uRymYVgxCAH6B/ZLxZYeh72BRseQkTYXCVmYAf+Zrhz0AdS1H
xpH77kmeUt3JIOWzvdnqkKluwFc2n7ITk00FDP2FWkYYujxZXhE2ISSB8Y96
dTo2BEPK8E4iEONjfHUFF6YTJqUrmMIZz86VP6C9f6/ehrlzBfyqO5DzdwMd
Ju082Kmfo19ItyDBdsfybhgI2EVoyiz/VaCXBR7R4DgU9m3fRzLCYH/WW2cv
WpgmoS51KkCgHuqOZWWUm91rAzHcGmG/BIoV3tIjtMVdVM6l6gx9FyOHyFYd
INPaoJrH6hkiAhEZWxOQSziRrYIHx5jEclrjMKOCTJM9FRSf2t5Hzf1qGYUI
RgoZOdvtAUPAMs+8mKyYSqiBmCCvQxMi/Eu+iM42+Pm3V18zB7Bx3TCajiL5
ojIgB/SzV49zLIyxerNfQ8uI6ayTIZJI4duGMAfPV/S8rHGW2MpGDcOsZ7Xe
RQbJh/VqIXi7Ix6SmzV6xbbzf+K17igj+ngfl2FNqLP0d+6BoID7/mLrjbxX
ENNmSnassyzIs4K7Dxhp/df75eYlNaRrcZOOE5hXzlOLblchBm11UJGHgn4B
gxdNjyRI+3Lfr9W4jlFUNhc2xk4Nn8gqhCXCB4IEnqKRA/+qHGfNqsx4yYZG
Jk056kzI3p7htXzkUmdOVW4kSbxUIh8qcJZVxku66dPQrOTjCejbZ1BH0ICI
OTI6i5qQHMnqsSbs9xVlYkbrF/77f8wPmX1+dG7wXbkkOzMLDWFuy/CzCbQ5
McFiH4WAbMEwLSfEPZCGJfpZggScEtv9i6fW+a2LJx5bhIRCxU6x5su+nTdl
25jmRuYbau2WDLB6u92FW15QwzWu1pNB1wbyskq7+22Zr/mCJY8NDE1RhwW0
gvy09PT/qG4yJpV27ZBxQkgGZj/A9QVUh68m4K4PhmDN7+JGMXiJv4yfRzP9
qFVTtufKftC0cJQI+t0jUCCFvGKeDf+DVT0S6Q7BvZM3/cBbcUYdKXcwZUq7
TGsCouqcygsb3C2szOA39QL4EY9gRdweoqZ6JP6mBYqCfq2mvthbFyDNSKZW
9Cffy1Vfmsi3Pr6xOq+aO0HclMT/Z3W5QVhxon7svUmslJC4uo6nCudhPk+1
cbhzD0sXnZg4Nm+V67HtqMcYbE5zAXXhnUXurPqvbT1QmwEAvGqyOf59gA2M
7AYcHHDIHjLvf/i6KbozM5QVhN9rW8ygbKpZnaPkDZsN629Gq3yWcsefIe09
CKgct+NbZDPZSKF8S/pAoAFk9Tk5CAPkfhgy7runcjiAt7s8AIFlCU/vf+Bq
6wMkYYVCk91LVITAxtMUH/WOznLp7qudYzELYAlIsu0AOhoFr7dEO9pYaN07
kui/y+VegmQierckNj39mwNiAAgmH//yNtfOMuejdBrT57IK9g1L/q2KljD7
y15JLhcx9pc3cr3lvwdteXLwpfm1beEzEVE2xfA0bv0hGGvF4Mtu1cDO3jBK
uTKSE+NmOLFslPmC94pYxO6U0N/jW0ya5a4MjIy6S7aUjHfkyNVo0Ndr7aNT
hTYwwGiG6EGtCs0RCEY+PXQjhtfagaXX29anT3UQzaPs+hYbbBtrbphNVi7+
k/SuKa8bO5U7hs3U7GMkB8dRo90emoLGCpW7W1d6uXejp9hM0yHR5DIFJzUK
G0TJaLmXDzmI3pF07JjlJbl28B4YyghP9e00zKwM+tq/ikzPnYtk3mSr0ggU
pku57lrHTjXbwTUNbTOO7TbhmU71rC0xQS6srLf3yi0n81TuUh3qGZTSHgwP
UhUvoBelDWaoOvdhjJYUXHKGvjfs/txKQvEbAsXnRRecffSElJiJK44U5g+n
ZWP5KoC5qqShayaZ+G3oR4gmC/OZDnPQGhaSGGxveW1V9LhX1wugrd6ApD3S
Mf8q2n9sN12gRv726LiuEZhL0cky3VJk3H+wvVz85mEb9cxVzSeFXHVspq3Q
V6a6OfLU2CAAOJn24aYj6zDdPF4BPJn6q2BzL2cJ1sRWDfvvubWyxbTedoK8
29f01AZ3n4jyLPJIiGRxP3LFD9KFZqNAjL5/nXq5ov0XhbAbqbm4glkQQ1mz
lWohrEqFN1oXOehc3+/20I6lbhr92/3pCpboutEfo0BSORO/+gkDZQQH0yrO
vLSp2D1rkx8ATbrEMPoY79Hn/zgvQZHT3m3FMgpO/lM7cNmtnbjL3TqS5EEj
FG+XAihU+DiuKMCXrU/zf/oTxq6J2bBpplvmkmN8kHjA+mimRdvTHiDrkk13
3O+8MKIh1Jhfs3LVZ320ZrXd19gzIZ14MS5dG6BbbXkClC9Sqxi6280ky6Hx
rdIZx2DWhWd8nJDaYesGTUZpbd2EURz0XjcsrpiP4nagtD53LKpl5rP6KxKB
T/wbBaD0pWHNOdZDMPkXfAdG/ACylTTZ876y+sZ4GWMJjaiA82vp7KjiL8We
cb/L8Gc7DtxmfUnwq6xqW3HcTWuY0SHlVFecCcAO8WRomBdRnVQ+wd2iifXC
e9U4YwHsGMm5lIjDtAVSlz9MsIXFTqbCqPXW1s/oaBIAJSyz3Om0Zkadc7wb
OGVJoEijAL7qNMTu1PDjU2j2iibpaBMP6EpATTwI2sUmDI0vaHA07FIHNTwP
C3fql9boDAIc+JcZ/lOSCOsmFZMv/cl3jcfRrAzimiybQ6P226mZkOET5jwf
vSutFsJfqkmtEzA6hqsFissvZeoeDkRBXCJ1JjJmyB0Klq8WfkQWZ2GLxBnU
tmBVojdKLEXO26U4ltVpNv3v8o9V85kdmRzV3OzFwNsy1GF5Pwj9++JQXnEt
bqot3AtT86Hr0vYSVJOOF1zJ6SqUoBeVBLmJx0NYpgnU1IgVSNmVntkjXU/x
SjMFn1wr6wDwroh9ut0jJnGXDt9kHVsrgaHqVzM8pwtq3yfHUAEsyLpjO2U9
NeMohZCOdhSI4JeFHMLZ9sHs+ed4pCU9+ME2AbvYnYcYw29te+RJ4iOhMZJ3
vmzxtVEgGHRX+DyBpWRLkYsZ+wce6t93p+sjT9UxnJNnyOjGKiXPiP26QQpS
dFJgEDFdkzGjQHFq3Pdv5UdpGjluHjoxDdTfCKNy8aJOQ56EWMp1djqAu8Ay
Gt5kg2orcSkbbD+iz89ag4cNWHDt+HePfkf5hQfV8L3mWzaogIQFqyVTvERu
5dKt/n14eo381kra6fgc+DBinOvL3NQkx/pKuEzCO0Ra8Q7jWR9do/pl9V3n
DSI2fyKE4Ij7b+FRAfM9XuKLvnSpLg1h+BOSS8RmnOERbqUfT+6Fn8xZtpfp
UpLqRr1lihFebgKNnA07NP/HT37lgv/abeONGlR/tOo2nGqdN9OFLRZQ0dvK
W+k3nSzAkcOPcnHmmzKmB0BrsjD33QfUzYsW52myE5Mg0df2y2ymWQq9LRLA
AcNDXQPgJH1YGivf66Xqp3fpbHXoRBiJhga98b4IwFfD7IvzeSIbsKrLq9tC
BCDgPmUbH7OQqbBk03ElSP/o0YIARQGg/k31Y/RYsRhVzMAev+j5rZtFbdxm
sKGGPhlIOMFA+TI2PAW0nVz2RS/IAQeyxTZhGta1MlB3SFvSDg61cxWaJeeE
IKW+vHWnolVB02oR7oNEhAypVXk4RWDgufsEUkn9OeEtv3K/aE1m1KABi/Kd
v7ICycMab336K+zogLfLcdamqYowgiBtjpR7nBVJrEAl8yPe09rC9UlnMzi4
DVko+IDhi3tQtmqaUKG5O9M8b9rnFNzvHnp0r1VZC9cmQFUmL5+iqdGntpbW
YTBLN+levMHZkrY8feXXt0pRqG8yxOxbwd12Lj5OUkhiukwJKsCRiu453+qT
h9sPkGzKqUfQNjaLCTaso0OC8rIhd6sZkJ3sIztHozwlGy+BBZynsoLTlUsh
xYRRrad1d2CaMCCPuJAY1zPMqqEfKVuhJSeMcY9Tr+DHLJyXlwk09l2nuLie
IcRzZn2fM+dbpnIqKP3iQ11TEBdLtcXEhCiQ7zkCy+jfBsdcljrYNFHh9TnG
nnhqngI9O8zx98dCenMJciB8Mv0lcQ4c04T6E4KbGLU0ZFSzglCWgOggSN+D
XrwBLKWmOY/ZKP/lRg1EHuvcBSBzVCPiRpKS6+4X+AVgDgiDTwWtQ/NG9nKQ
YFJPowvz4r9Da7y8ntMqGuwAdqj6xcGtcwQaVr03AQKRoOOJl9LynZd3NEKx
gMPOINQLZYhjk0LjW+CzhVQY+LBXgj1dqqqYa8tqgcbRlTW1tqVq0jtP0FR1
FD1GQ9KT4HHo5B6tUnsCv2tenT7FqfFHIJaLZdjuL7A8OdqeHbR8eyWM8oEc
vD/QbZ46zWTs1TcNByxKF1YPRW7a9OO9fO7MBIRV/goHV8K7dUCCQyj7ZIpc
U0eiXx4B8l50bJM7Qn/GaPmSDXQVWFJEd7Z6pzYTWDEEeziFNLxOJ5JsdUDr
LjO0OXbIWUo7XO7VJ1OqB/rkTPXRtEugz4MpPJOAObU2CaR/SJ8QFeIpkSe5
zlWlCSv7R09VJlN6DR7f8PjPxMBhG4JB65Ri4NibOCsGrB5Q3r5be4KOqxpV
z+xzJeB4zqhV7ON3y+G9tzsQBjn7KYxQToa9PCPXYpM60e8G48HlJkDIHas4
KGWwbvDmQULub1brZEltuTQ34CR6HC77GvJlBnRbdRKrsoWAgvSP+vitB9p7
/PnhtVee1pzxS/CM/F/Dah2h4UweA/tfev4m4g7y18QWtbw02dgot7sGWY1a
+IlMEM+yw4imknapw6GBQO5kyzhamrKftmeFN+K9gfE1/+RonmhH+m5JSVeW
ML/w8xIhw5mxKWO0hJgeLeHnLPtj/EQMc0ZhAEK6WYrgnAfW2Fy0lYyMNuGA
Sy/nvXMNexnJpr7DyWO/wKmofaNLAhWCutreY05Nnhvd7kVfsYNXRz2++ViA
lkIRI8K0yRU5D8Y2a1YTbwI6dAsf5W9ck+PRjjxmPSdfwegq3O4rlmdRzRXN
JtUsnoGLPqRjp3naNCRRJgVd1ExCIuckG8mfjRx/UH//Fh0v3g5A2yo8t+Ck
Oi4f318ZMkPio+e9J1uKZIVBYSbJUGkjoaBMiVIl3sb7hmB9aH4ZVNbuMs+3
t82TsVW70Pj5p277aEUWIBr+QotR0w5SmhsRtbGvOMISY+M+CvtvgJvcoNlq
rS8Un5eYVYxksx+HrYzJQTovEiQ3b2dU8ewQZLehCOAdzjZc40RVOA2VAbI9
izW2ke0CCVfINOSemv2n4F7pcFHpVOAL/iNwEEtSYk91c6VBrIR6CvEWJBOs
S/G3zCFYCduKenGiCdCKoyaAQ1Lf+6VnEoOC5aBIOgG+nQE5OXBf0oqTRdNN
xuDcNxYkJnAQ4EpYWiCe3NTdzPL70mFIBnhcGKAx+/GJ2bZs/7Tzeljwci9C
9UmxL6FAu5tB2oBemGprgDvXyKE6IJt08z6xWQmLsgpTRgrwj5La+u1LG1cl
BBTBMv2jBcKUFxwerZPF2lN5H1NPwoOqJUE7WGFPhqMSPbtuEUsaQZqEztLv
wON1M42hHFbj7Y4lsdlG+2MOvluWYYZ0ov6eFlVwwJRAN4BbcCsLo67Ff2x7
VZlfO/lzNutdYvlHBRr35eddHOYW4o07rNLWe3M+7HF1hVUoUir76gE0OdyL
qtLU/WmLnpxxgquMf+82k+VVH1Kkf7YD5lh5FHIx3SwqFOevS6UJFDBloJeO
VeC14gthVPaUTzjy9NLdaGv0ZCQtNJOQBXLJlMr3phh3NmiZixKpKkmK/8ww
lXljn4WvF05VL8EZlInAwsx4gyB7yC0fJqYgCpeler+xqwCx0Osivypx0zYU
tPbO8qpb2K8H4F26yKtDlaFlm1E4DsMNR9NB+1TzEd9YqJLcjTj7IN6DBubl
ZemAt9lopoRD1EuT8/1iH3jRZSDkOytRhLm5HxClLcil8c/8cGe4jme8UIf2
D7V5Ceu3h8HNsCuEkeDvuzXRAneBH4aTdK8oiSPXfsKBl+eGfq6Rjec9twTL
QFKAkVzL3RWxEvQZuTQtmNQhqP3E5Lsjl5MAyNXiC18k9HEfIWUAXrrSomPX
E+6SkzYWbHb7p0OUyACsEUPQeW4StQo2YMAe5qYKX+kiF48HnOWc1/ApNEAM
n7gd20cZxfDTunqnQPi9PiJG8iz7VYdVae+eNi8p2GEl5joPk1/sVQM4grN9
5ZEGncabZ4hL5oH70+d3oiHNN8Am2hdRlvWoaCR9VtX2w2mDKrroR5jSsF71
cxEohY5jK8n0RkZ8wNCzqmQCf5QKEz6mlSnsH3HgEfOJFTXXQSg/tGa56iDw
hNOMcBMrUCu+IfQV/A/+8t6DPLyzAfR6ujMCLagvc7Lyg64yHDKbLkSOoyxE
hAtDM8r5IfTI47gnmr6U/e8S5XnGjK8jpNaEla34nVA5iKHCWzH1FJqR2Z8m
QYUTFjSJobI+DbqH36wywhQoRH/8xgsHAh8x0wJsbmI7/dutb201Ca8URb+8
TneUPtY7Rm2fJ8I8qUugMz4n6WQAEKrf2qDnaSJT/fj+FFPSc/amHZeySXrD
jgM3ft9d1N9fWN1EMnJEpj8gxpoUzZ6+oEuKcYYpUOQbXP3KaYyqTu4fGLxE
gA6bYfr6SebOQLjLAwD+cmz7sIwocrhEG3VnqQFYMLsGOmsE6cU3v1dD8mnA
srDCDM0aCV8ho4JvhihXbUYWXu0kBhL0pxospdoUzr6R3SHbuAvH/rAiZj1t
cn2cG0R4cn0zXVsW9HCHhklB6hdWWuVvS6e+dgSG+sfNxQ0hgUKXn/7eb8GA
9JoUaCTcla3ROholgc6x/wsNoprWYfR2Ybhe7zHPe31hLvp3mUUodODBECDM
vqvb8B9ztx1TFLDCWS+/y506l/7o5FbhbkLax9eAJsL0eXJFI8Xw/X5YlL8W
otxHQnkGhVbVgq8+9qwk1Svo2DkwPMeSTdZzD5IqLvlepzTq9UIQIM4dy0g5
1qBKWiF1deph2+lZ4CprS3PFzX4QghRZNLmYrYxAAHuuBOidgxj78UQnKEeo
j3hAz5Yb2iTvhaafjFNPL4UXxMARh9lCIAUH1TmzDlN7BqrR8NTZ1AL8uqF7
oe9keJ/6eikEuUoPR2M4B/oJJUn6BBPnRFBAs93ZGSNP3iQ6WA1YYZc6n83H
M3Q0ivmmBVnPkFqrlPh7JD7hfDJuZZK7zKZhfgvq6XCzk2+al7u7pdxgEX97
+7eTyqWgF9tCl4j9GTSJaRIIsfIo0gmZbWuqG4ENwQACmGi1HnNbPvd7gkYh
EWEbWRvL74lmkv9ITlgv7BOzvC74YKiAO8ElL6BZdJ1MiOYAy468tVsUBOvB
CvgiwHv8ttMOSov0N1bhnTva/037a72AGrkwypOVB083N2N22QInytn2SgH5
do02EJJVBcPwNLzMw5vShAr+Y8deJ7gBJ/pwxqTyvhDfiSTP6wVmb/qgBCsk
H4gmrTSnXUk9YNgXtJgvLcxOuw7FIUr0vGIjkE+bBVMGD3Smidiegp161T2J
iVmN4nrouYZZipx20q4huhFTnyMZJ4WqqGFQ9je8ZBRKknYvgdw5DtN12rLL
W0MsLwi0I2qz+4xjzXgjRiIOCy4S+s9DTzOH4sxX9K0cplXMscbV/YeXqvoj
g9pz/SzHtQMsNU7y0fPX0Zgh76K9UsO8BixMLnXv64LEqgNrGh1PwPvjmYxv
cTVAUkNxWAR/SArTVGrwJX3d2ZHvozzpSIBx5ac6NxECKwC+P4Uk7RGr8kqp
TF1gi3zhLDYrZd6WmlqFroK3HVjuSwoTmx+R6B97kj/mcZP7DUoV/OnNKonJ
pe8XWS6h0B86GCp3uMf9LSEcGO4PhWi7xDJSfhsvnzEbBvcTU4a2khXkQ/xi
FMP8alqB7A9CtUPgHG7uAKHSj+eCJtCzMUmaj7aFjxIeWKULNwu2tkbDKjde
ijkjm2jI/hyjTRYVm6UfByK4vxjVRAMfPtdDmkCzQVb06Svmvy0GRiK7tWE8
J0VwLgDvuxW4I5mFGw14mIi7XRAdA82nSuEsJsV+JxBTyLaJ9/Iz7u8JPVk5
zc4CHTGKBrkMHYQWmb6Z8Q/6m1s6/tcCoKmUA5s5BcSdNIGwh7srU9G30eKc
xlKRcBmpf7+uYOHw/amKBPKo6zkYoqh2ywEljFwASLfhYMJsm3hXsKbEqKUx
poHoU3RevfQH/gHGne86/TH1ZvfRdrnzPfkqL3H4HyO5kisDVu1GTYeLIsxo
ifJR1+Vs9qeax2WmWOzL7FBxhdkAA2obXOm9GunB6dUDYCz/t3YSXDXIZXEf
3wcl6IHhXfpe3piKWB6GDCYy28xjtzZ2bnZFQ80Jg/MlPWz4OHQNO3Wigk2C
R+6dnKwahxmoh9PYTM7VxA+0P0g8ciEWT+vGnW2qwvx1FIlgc/d00XJ/MUFJ
v8CtDkvDM/NkaopGskHgo3v2KSNeHo+prk/fhjVsPyQF/whRQPlRKFf83M46
DgAqqP+WAo8nKgj184/J/6BZwyC+r3oj5mMNM8Zc8kUmzkH+0QgJ//UGFoMU
/4c/U8Z8/jd1j89qcN39lmwF6VhpP4lFyQ7TYmbwLB6N3EpPLvSdYH8n7h9e
okX7aI+JJT4DlEGHK1xJk1mzhlQpX/4FlnG38qDbiS0435c9QeKGCNv+lsoH
OUZRX8UDwqbvS/WUbeVRox2HIve4IIwpNCK98PBnz/4iEUbVo+ixRSYH1fW1
5H6VqwIaj92MH9qD83IxRsEUwqbtpanFrTKFdq8nbp+m7YIxASd5jRrMimjx
lfVqgoaUMnJL7JcPJzQNaDqacKYAvrkslCY1kX+iVgvFCCVVq54ruPZiRUPk
jv+LJ8158tMYtlY5939ccf3yuJPmS1QS/o+p695VemiRRQiqCYOr6tPISqvD
LpkMwRFABu9QJ6N3uNPOfPgFSG+EJV6XFhgZ8wOg0YnO0QqAt/Ea4ayJD4aF
ANpK6LQWRyQbbL9WHz81FsuHo8WiynYUwxFLVVdVh7kf0kb8GKKYdeOa9qVW
2MoKbiNDVHFzTYTVqWnsayIk5VAAxDEnpdKVa+HaPfvnLYWVOuGfv0magI/E
S8JgE8hQj0lWVVJhkZc8/BXEyzZ2llxuDKTuLSqNN9qZcwHSOBqXdIObzbp4
0zxEHslkV9P6A62doGP661FeRA7N0Ori2EH01JarJk9Jb9OKVDQzl12I1hSz
+Hc/z7rvsOfq1qfDYtRSpTnnG5F3eB4sI7r8+fhFYTo4Mdyf0wrc1w7pldX3
zD3Tei9bcEjSpHvnsfFlRfK6IlKn5AcZfRN60XSgvPblvIoUHOm5lgUoH4+e
Jb5A0Vi/44DObHnuOe4RAiayq9ji+BqbwUq2UV9q3joDaMTsVVU6SJ4Q/phe
6ZDScOgJ9bqNd4otIIUDUP4YWQ95veluxzr9Iv8gwuDOrWpLFsiv5lzccpet
xsgw8y8WI64nI/2pY8iYHFFkapJDSoPNoS/quEHi2+7box2pxyv/i+y24pBS
8TPP9nN68tmcEynkKHruVLrP2PlWAgpCqqlTbYdPPHUcZjBqQ+kv6BC012ya
vRo2YDtqjweb/uwcWsyRx1YNBWRJ0sfm/juQCcKbmtK0ocjFXvYj38c0fnFu
16YMsPvRmSmbslBkV69N49+Hob6PRg7X79OfP64mXNjrKa3ejRNzTt89z1wk
JUmIQFKxMpt6ACxzjW8WP0ioSS9/a/xRuBYLr7RKJU4g3sYqXrFWwfBuAlBu
J666uPKyjTDHTOQMbhO/4kpnVub8tuCh1L9syQWUEJ/sqzQ78Yw5iHTUw0sa
ZoriMDTKeSf6IAE1m/HTeV0A58gOofJSb6updZ1+dloYSkEDFzaDSYd51Xjq
fURNVqKYPdpCPh0ypXhpuwsW+cuY2/aNhhGXJ85sIwlWVHV3a8jkrGZKhtJ4
yjexCQVrIKAU0UOIgAjircPtjc025TQE3J4J/jZZqAmxhirRubfNptSzKHbd
BrfkYP7dz1KvA095kCXHj4vgfChlqNDRNs6zJPInZ3aD4o764IRrvKKZ1eP2
AEIAF0NiJAi4Lrjmsh5Z2KoqT3CUOcFAIsEquEEmO+VBW21/cF5LcALdfOft
ACqD7SDmOZpiI60sd+KdtDFeZHTVw4kyK8OScIra1KubnPoxwKUb3TKvBusg
tKNsXsYyfIemcO3/DwXwdiI9Rlvg/jUHWhlc1VTwsj+ca8VYpTPTc5/kNCUz
TAav+oHZLw4xfyMEaeTXVuCZVPnXTvcgAjSjqpjrRTZJTUktGODgjYUAF7IS
sdBRlv/gbwctGoyNEcKHYVABJphMFFu4Lb0s6NXG5zjy6EQ/sza/Egs2oQq0
+Nbb+SG7rblpjJ34j1cb9IW0rnSGUZrIIXn/d5SqLaU4hEZmNxJgMYspb+lo
sut9TnfPrZZzsEKnxNe6YiGv4U6Zd6VoSabJyhrstMwFKhUyhcDxeNf3xqTS
+VzsEArOKooy2g6tY5y+THAJXRtcBExao+JMRIIfQwBP5qM84HU24Xfj7+3y
7vFEfl9lO9Duxqmoe4Nc91m39Sr7NLK44cEy8SV5jftfpzco3xSQaMol+RPm
ujVdmu+Rn4ZnQkhVLsHUMOE0y0jo1ANJjpJ+IfnthpF0+jNhhKuCUy3hM8w6
Ap/d/svV/7oCnoCYzSDIt0Ey1Z/QUTJju7r4qy4/FLj+u5gpB7SLlS6Ph6WC
HrdSsx/DUmalvdYASSk9JLaP+j2ll9L691rZwY7eV1xBKmwc4QR6uX314fz+
9Lj4ezmMCpUOT9H9PFviBJ6t+ljMRxV7fEHAEN6bCsxS6uPVfUctpsV16AZu
S3bDuYYDdoj1np33I1GwTTbLH831KQ0O0Mx2m8IjtbOzA/Xi02Na++Tl1ivG
FZMyCxOmSBQGkRlbtFzEp3BoP1iL0Tt62GnijvnJTw9EnYzBPje9D7ryqFso
MX5lymYPzAttzSQhJtsj/6G2L7lMpgvOwj+pdVXYL6U6o+O73ZOc9us/n+Ei
ODF32cFEFbAdnpDbvOJZxAutqJr75o4y2weAeNMFJl+ULBBUNfUSuDHXZLij
XyWZOJKV/lSpV31PpRFGf7iPFAuu7R64jglbf9ToYD62VpYSXIGhEiLEbRox
9NLri9aCB2oCmNwFgit//xX3g1w29cxYLO2ezhANNrGbf/kwgRtQOoVeBceS
Li9eKfOhaV4/j+vewwQHCAbsNMpYwQ03hB9ljF6t2Qxh3QzegmujwhxD+qZe
q4g+M3vg809VFOcUwSsvy+t52OU00B9Uxb08mwom0UHueaMglg+Qll/62tpB
YjFckc1GR+U49yh4DO1Ouv70OTyaCfCQyTGKaIJF7/jZaduA1KVFWDEpTWXd
mJV6/FlR8EvukPiWX8LwNUVLnCdwpvTq2Q3Qc6qLT5H8vVypBZL1vqYeUbrh
Hqs1FJzA+0hiHSEUpeKNd053DGcECSEEG87B5hxXjDDRlf+fgmXg8EVlbJsO
2vwN+0w7ClciANAhO1cOrnN9oSttmJv151qoG8zKno7xK+b4Mjs0ojcQhTsd
cG4ecAQLsstn5wNEO50GwperbdxWJwDEew4LEsIsv0eWZYTXLLmhnsfWMSSh
qPREYhn8uFPVeZ02k5rE/WpLzrrQjTNdZjfwOXCf8mPjtJDVPZ+VlLXJI2pw
UMxfEhwc0F0cufOGXs4ztrNn17/CpSW9TnBbtUNobKT1DtJATOTouYUfQ6pA
vuaBYsYDTKnpYuEMQt2V1neV88n73RMjqiq0DVz6aCW5vzBt9Aw9nkKeUgU0
eE+7+yjb5dy8GEpDCew6NFp3MjX/SDIYAkqjyWmDIvSbhjj5F+RAJA2SilsH
7UAZrvIMqNx5frQKnaLv2vNWJp33I423iZy3jBk2tK38mh61YMdydJkRuUF+
uix+FpkfqUZWifUWA8WjQJlGxcpqm+kYsLCZrlrskZPiwsU2WV4CBgpLPT5v
P5Ktj+9ldH5DsvYubHiWGzBMNuPlTp826/ewrnvJFP0aCswqbktxzOOpq90G
3h6cM0o1o4FiUeM5FoSwXxIwfxRAKqEbKwG60wjt/k/Bs/c37OFG1h6qEYKR
1kiMp/Y2ZmZL++0fd+JH1clU8JAcSLgx3CTfh7vTODH8moF0u6SWV5vjFFMJ
6CxQolwBByvIXu6sHxdmwdX/SwzwNI1ufufHlBasK0OoglQ3gRCONl1vc4Eg
Q5CbSQK8EfSo8d0F9IudvFSX4PLulaMyZ4pt+GxqD7xAj90G2eGYOTeYMS6U
Iynw95chr26BszNemGuyITAtFwFrVdjdOMDEpykNqVZEDuzH4i1ZwO/0Urcm
vEm2LU++8VEavJsApDiJkRS+jW0Dyu7uKFGxptbdRx5tNX/CPrKttwiZ5xQ8
wcMKTyf9lNj9PiqW6++gzPTpm4idN24QUfgRx14mZ6FCxhswSZhwAbhM4Y4L
rzR904flFoSsxA0aMBVONzUGlLKVYWASh1gNMHght2soHvw0mgzz7jPqkOBJ
rYT6B5hRTFkTcqunzdzV9fAtZ+gjxbUNyHRCLL01hzEv/qVka/iGjY4x57g8
9kpEDEPEKOCwN8ASsfsJEzW4ZRWxKcY283w4zbJywzEpGxIrS04o1QAGilQo
sQYUDD6j+dAMoHZzX3lWqEzwGksW6b9lDBkKFuyRXXkqjKJnCN00TMOpR5Q+
R38gKyltu000Pbqbp6n4J6+61g0vkcBdi9j4x1evz8ZvPmovg4OZX78cGGbD
tnWjEJ0uJ8bMEPKth7Q/jHHEtMLyAdnzQRBVWFiefnogq6i/AEKbG9cQZcRy
GhCt2lCPK7Gb/CN2AWtK4IY8TdmYP4rMQ//0w5NcFs5B8uBQ1rEq/sLSJi24
88b0Tw7MF6pIx7HKJQbvL0CCp204mU9l2cfTjyDmUmO7S2CVqsVH2Q56f2Dy
5Mj9gu7gWiD+4SaEMHqSNBRJlFHKIxJ3nTKiqGo9qQYaHk6HvakRdzmmBYnq
gdC4VL4r2GQxmAsLwtm0NNn2d1TQvMK56cQKh8KWIG7sIbdTHtIxIJNxutUt
YjOHHNh0intPVjCMh9yRKvdXXnkmpq3CZe5738PGg6vr33yv2iyYvzWX21KB
CJQ5IUQVRZ+Nw98x6TSAqdHEBV2CA+ls00qb8Ah7ykbcmIylzmz/EHjlVPAm
gYgNQ8EUiP37AYKWt7/HhumzUYk6tiZ7dUtnyhkc9l466l2OCPyN0p04csKt
hyRObfyi6totGQKGyM3wmuwtbD9q6F23wHouUg0ZNl7FGBo/vj3YQmotDZqK
1l/1Lfh0pKglQbWJ5f1bT7O7mmi2CNTJh7ajU1qGbG1oXxQC1UPPMFNqfJsY
oOdbMJSy80cbf4USqRQe6SvYlH2/PMNwOHzzEDK9duWUQ/TMgtr7w9YxMDND
MZ4taxtC6D0v5FobV7kJG+ez8Pcvw9Uke0LMCVFYd6GAdLOdr9sfccQZFCA9
SF2xfa7OyisaqiK+in24O40UfuS3MBrPkS587GszWy6e2Jasp8QdFswKzJO4
LJKV5OFFa48Zxz93JAZDCUzCzFn50L9VtZTmw4V3iwGOq7zs6aPwJChUNlBx
Xy8E8qP7+sBhHsC4aVlME+rdmZja5sjhNLS3QhkC0+g5TcCvi4zsguEJILYv
tyXebKVvV1gAjOYf577ff3spSrlCiH9vGJjaeuU6z1swRHfkF8xMmcm+OgHb
Z1z2bxgyoyp3r5w4x5b0tlIK2aXeTqRN4Xhh/3kDfrLRIkzYQfpJmamGLF+Y
cJgyu6i73bPZLSsh9+mJ9Iy5Qf+1DYhGZW2bX0D+B0POkyUNz6FZ2QlnPHbk
El5W+lf3VyRgp39yhkFljaWj5TzsXui7mJy9AFYMVNTiaiyGK2mlpc+ZqDhI
4kbDC1N96ORtyFEfjmQyIHmNWyoqtCGyGt8yUOe5ZAo2dq2MbEmU1ScOatnY
YwFN1g4bB6WGAbS1F0BaftpzGhxXqB2mNQgtR9qv++DueglUCkSKWuR44UHI
X8U4yR/Ie69ZC/L4su3rKWHY9VQp6t9AjGIboSB2IbsWt8l0YkhOt/8WBkMz
KfUnnGnaafPQ2LrLiTTKfSBAUNQBFE/l9aqCOaMGShnGQz/dj9hFsYhi0R12
lA+H70KLZEdDfMLJH004I3mizzqQIdarFIyJNcha02N9m7tQfFKMlwjKoZJt
J31BQNsFF85bGnfUgJ48dhUGRCBcfQYWnVhmlOXd5iaOOU8iMr84Ja1hMuYY
2BjY5XHPn6kc8QkFTb5vn+Dd/4jOQ273Ovf1tVh87ptW3dmo/Wc4WfPswQWi
4GgQh7rrbKQUGSvXulN02Y0pMl65ho88KFBhc9HeAfn+kgwqgc4cNZjFXGC4
f2Fe4CHrmsybXt9nk/ULHnlPnnqsjQJaYguHb5jOw+IVA32PmmltGQsnx4JY
ngJSSdPYV/+QAlgbHMAnOznj1yvKzTxYv+VmOlKtB6zV+YIH20aIwHgBQX3L
n9U3WbT6dtr3kBvjSn4wsn/nXR5RkyB+wRzCrEmZCMpCZLOR2sW+8fwz/keb
hJaZA2NSJyMBCb8jmf6K7SxIo2fQiVT5YiMv/ptPg5XVm8OTKUJ4M9PbFVWf
pIO/Ut5Wr+roJlb1AWRpemlXtoZPH+CAeUBQHHcmjmzEF39bXYFrfjjCTyc3
yxXlE9oZhzbIib0YxjGo6ENCW/U0SIW5lm919t6WcM09JtR8oSpdks+9V4Mr
DHhdL6RRyJCouADjrCnpcxkX5DLGpnB+wGDo4a2iknhsHvrPTIVRM96uKlCV
HirnvNxSSHoA66mHcdroKT+TP1MzHof2EcUfbR+vc/hUwZ/eWHq9uCtEDLsf
1ZfPT7D2XwbJpvyjEd2dOQhTnqZHeOO120ESryYt0hpwT4ZVLi2guOhwjKiw
FQsBM0SYWSAjxDTUcJyWEgL1jWfgpSgVkhI1N+NShCbj74r+JNHC4D4kA9bj
V90QQkvXdnJl0x3+BxFeMiKAaM4s9QG8GOBc/TuvmiagWaGB7gZl/+gZxWrn
RXxK2FLVn0C1EnXMaH++TQBV8kxhrlOkSBb8trlr6PB92YUWbQbY7zoXBWrZ
7OitBRmS4Z6Gcetm+nOYeC6KgR/XZ7EGtw3QlSUipSk2vgVbt5TqrwVOOEJR
yhHLdOEs8z9lIr4rMHP8AoLwFBZguCcXDp36I8OOg5Kl0MDfBsPf0DhWS7GL
aap7g9VJYvXKxvh370vB8gCkB7rit1CnFx0sOfp2iAgvl0kLO/BGJ+g+8aa8
6Q9nNlbYYfgYXBCshmPwyYVeFt1S9BzAlkNx5UeLggiW2E+gkRGxru4AE7/+
YTN54rEx7kqdN71dGUDX1fpx/8MffRyHGFswhnXJH4bLV4+lAojPXI6Q0bYe
/QCsTRJMJzANJjOp/Gw7Cr69ad3ICRPv7StdWTKrdiH2OBa2K8QRGecC91Ot
Htnbgjo5k/sFMr2sIjygnW1NJZKPHpWlJxVdawvLKwRfUkjCH5nU5QI8+pA4
6e+1GbRz2MCY4rYLFzsnClRcQ40E6JgmYzbtKN81IiXHFC6MTs422V5oBlHF
OzrW8mqg7fm+NTQigoba864bHUEWKEb05OxJOIcwQOxHLA+n1DhpPOfHhs6A
/FFegZz1HyXSYNbrUzO4ReqJLvpfF99nRwCyzPPpTFKsSf2g2FWLW2JkroRw
IyDZdj2baSoNvhdmsxfsqzvSETg53Dqjo/hb6r3EXqkSHUJjEpXsQbH2SicN
nNgnRk3N+AK7VXD4MyF1Qr+sqDFjwqy6tOYcIcbnW0EqfWjdj1BGz71rINAL
+YWuF3+pTewcYO5ptf3MvTErtdszGaQCVuifK5rJR1hCyae2WhdGb+ZYE1BN
pi9CTdG/suBLuSMCMFxaYPrQQ3/t3u/u5Sxga05b6dkIGl9YCf1rSpke16B2
qAaAlmsk9J/WvthNDfkD/s/lCMuSHfdaVIGajNutpC9okgGDD5i57J7j4gTU
TarOfHIcaH+hSDjVPblSiQUXO5hzpzavz27ry6xqi79GhCigRuRziDmjj/+C
hZuOqCdnzh9sxSLBR+Ys/Jg/UKQRCYqopb6UNlS+joDCP4QxCIP/gWGLinHY
kGx1YBfQSDqq4RKMxoHGa5AIpHG3CbZFYlHGxMP/N9QAx1vz8QXiHkDZKAcz
yhfw7a3xe6Pie47IdevH55Kh+5ZJQIhlh8Xip/xMp8hDPaDnE4t1HSl3/Ab2
1Z03DyBIR7/4TKf3g192Bk3rWLI9/ydDTKLo0cJC/Oj9WFvHrzXj06ken2M+
gF1k73fdUjlJzqSdMAq4A0MjgXA12v6si9ZKUfjej4ZftcKYF/h9cpbI5Bsb
4FOArlYCZlLzbC6NJzjlvy8uHbV9JRRk7VE7vamyEZAgYqVSJubadp1mR3VU
kGLzOSt33yEMekbRKe3it8trBwInvCUPVrsZj6+ZRtMjQb7GaIi9q0QJ9Yhm
02STP7J1zJ49Kap0Pya5U1m54NBFn5Xyhl3USW0kfimuutsRI3oNcNYJ25/G
dVY+3T98G7lopGnXCFh1Q6s4Pi890twJS+CtHPoqbPfAxSutTfjqB7Tjj08/
jAcfdk38bXMZE7W0Ehk6DZx+v8QuWNcE1mggu529DfyqADYOkoyhA4A+7SQX
VO5Gy8iVrPTfVMbE7LcoswyZR8/qwfnldoSGlrWyS011JhflCaF1PGsL8YgR
3gy85Sc064cyrQw+G0JKJOhX7pf5IAl9tcT5APCIaNQfHxTHVgPwbGwkPS2d
sUOPk1T5oRsTZqB7QaOj5/B4SdDg17UtDsiy30fXJkDflkkZeC1BC+HaSjQu
XYu/cRe7RgFWLoRDLBrCoyLbpnDZ/uyAbs/pl1gx0yuKviko4ZAs0gTPO2Sw
aWRTTrWCVNJa3mjqK2S93LJCyoHfSIwX2L8OjH1QlNkjo9mhyVMuWRspEG+l
QmlKfVPyj0MEULJRiRT/FjmjIr+XijeHuoTaTa7Is+AodmkCT68f92ZEkh2C
4vy/OgdkhoPuq9G6o7BR7YybgvbtRbkLps3AlDGCaEogCsjyy3mx0YjccPYx
ZUGM9e8cdKe4GOhjrZt/NCj1TDwAUgWcZ1pNeENILO8K1P64k9np672O6vYr
GyjNXC3jWZw8meyWMl9oPQRvp1iOk4Wt4Dvog8uJ2LhVcrjSCzDKJrE6pYew
ZTWUD4bk/OJpPCqRaxYnD7I6zDjtilaSVK0tqoDXSd2Rf3Uf1kit0YaRtLel
upx8TZdJg8AFuXrB0cTT25KFyIlQhTwTI0arm+lMpHMcHMfx8SfAlTPXlOqg
k4Jnbz2pJqsVTugvc1uZ9Fl0FrLf48Hu4Et7cLjW6OPPQGHm2C0RNYeBD7kQ
5rpCvgJbxeH/S0JYSLg169OZg7GvpffAg8SKKDMbMrDrZFe3Wvd1B9Fu7lSb
T7/T/5NivxA+o3tpnyy2kUqTXIRwNLPmnobhSs2+wcCwzYW85gL6imIocHYT
kJrsmXb0w3ktj48xhXPOUGE3wlb13CMxRqAcSnTimbLMFIfHur3drdiOu5XX
CGRstyATUQ8Q1Tg/DMLGVAWGY0LYLjCTXaGp2KhxV9+b+V/wNBl7+BlMncdn
3XwxFmNkeX1BsPYU9vVbVhKEKNr+TBxn6CrsqdO4iXQLU+SDi7ak9YkRudEK
CO/CMfe47ckAh0/AekeyWokesTfMGH6l9QJ5HGc1L8JcSUYdqtx6pRRVmRht
5/DG4U9nSY9PG0FgYq2sl1xP01LPK6rL00K9mLOurXqvk0fuKgi4LbA4b4M7
duBJZXEvHoBqs9cZwhVUhgdiP9Izw8rrQuOZ9QM4FyDAXe6qnxHT+/xTYNTt
37ibdfIpJ0+xWWV/Aku+rcsOUQqs1g7sYUlgmdTdvgvPxKOXmlx60FiXm8Mn
MsMmnNIWQLZQuShtJpoWrtdMWimNSkLMGi1rFX4maKI1ycwAoDO136wWwNNd
r9FXXKHydAFLjsDSib8UULHHVEFcmQUzI2MqvcNsLImoxlrdA4uHpfuAI4G3
+NFBOREJM1IYbWRG1hrWEO9lclWXBRUZXPiGawL9DV0/lT57IjLMQloUaUDB
V7G9gQ0DktmPuHLpTPXnVb9YeYlsDqq7+53O3p8KXed5wNqFR7aOVnxq5HDd
gR69xEQicfrx9EeXKpC3XC0nU+imikh89Gt9vAIXilS64qOWcK71UaTuCvUf
bmJzEchcnb1FKHk3kjq2Zy1JJ/RleZr7Y4HLCOMnbD4rMBq/DhjlJWolclAc
Ah99qXnIgvxO6d7T7pP2gfsriPCa9iQwrrWKiZ5ZZuN4OtxjEsvyy9Kb87cd
/+fnmAPk85fe2ooQ17HCjeqynUJye1CrSJBw/wxECIFx1CRyt7aSm259l6OE
VSY1frWEii3/SXsnp5T4PzVMRJ4xJwtGC6bDGCvGYPHXxSbhNRoQYgYHjR1S
9Bo1XOgJwSMIqT0LgwTqphzUNtbTKyMq7kssSjZnDLwBnutZ5u6Q97ix9n9X
Uqr0ssVeajKa4iW8epKN93It3/Klo3Yv+5Ked7NXtcoEjvqFWI7agUteApFc
QJoXvhcckspL1e9cY3zPa4j9U6uabHSG0JsUUFtrgvZJlhBPdTZQnB842p/e
xes0lkOohE7h52HOSDGO699U+0gBeEZ896aguDG/0BGN8RXIHx40Pe5IvywE
BH8YxCkqpHE/UKRhxefMwXVQiG47vYerlmMazqHpVGUcpt35lqxWaLbw9BXe
p1j5CXPNdVynw6neq8363kf8d6nyAUdbbAbrELt3r/w5f4zfT3Szrmt/wRca
b1mlYMeCatZRCVCcowHfG2IOB3KDsOo4i5E5XZUaRTgh+30jd5k5Ty/JXy8f
/cqmZ5/j4EBuJ5cAwDXIY/ADfA9Kl7jYiGEx0dEshXFuHitomMy3nHhH7UAU
xREistxKx1td49vNFU/8WPnh1LaH5YFuK+X+vN6X4TBBYlihgPuq7No1pM6r
EQr2QZyS/RU4Bl3Ouq89LQMNNOOsQH6kTK1cjUyBf3tRyZPJ2ehO/Dp/xiaz
YyJ/nq1TuKkeS4QiMWL0xekKOWkZEFHrSypHMAyDo7EyuB6hPIDaqWAbfzbc
eXSFvJhAwY2a5dIWSt72keOu96hasiMsvT72R2LJu/iasB97st4k3MDR4bcG
MAa39FCzLBJGS7KWMJoxSS9+ChbNkm9fiJxzXSZYIA0unC68JYLhd+pPnJNd
5auAgvTsseYNf9VckaBJpvuNC6s0L3FVifhgh/Im3l/3gkddEi/VfWRezz2U
+v2E+w9pCNKDHkJkeCGi2TMcyIQexUMI2X5F9IIdNSHhLNrFtk+HWUm2xr5x
fu04LU0rO/mSCVVXroLPiqkdmi/k+ErfCxMvmKoMTR4CcILB7CKe+V1wsin/
f71TI5/kSp2tfoLSPkzfpWA7Zg9ptKTsaZOOmio0efbpTZ7/6mWGOpvD9z5N
GzXagZZI15DZplYndLpoyxb7my0q8pI95A2hh5nczY3bnmh89qgk2g/O5qU7
g9BioQp49FUfnKlnAmNwEy/yol+fUVVvsAyE1E2wHns3A+ljuNJTYzb0oH5y
qJsSg+GDdFsI7fWeIC/MrbPGOrPa+xoJC4V0SPp6uKzoVZO8OCdjfk/k2StI
KgAr/kiFUkx6hP21Gu+a1cwjSonFkaKEU8M5gNdOwC4brsUwaYU+WF8+DoG3
pTRn/xnAJPCKOWK1jS+ZjEXLFEG4W3LjKGxH7T5wF0/jDT8Yh2WjVxNd8rdO
1hL6XgPxidLJ7q0aJ4FfdLZv83mISL5D3Rscj8K3vzYR9zl0Gqr092zIdmqs
hJe9cY/b6ppvqCT3X5TbwmZnTV2toOgeMm1q64DR0XOVvQRkigHpYlnGoga8
xT3dlKLe/JwMRfvSAsqGGko7ElupgtOTydnC/A6WDQOxaVQYfv/6hHIUubRv
d7e0ER92X0DGJxu559VpUL4FHlw/SGaM8LiOMc3xArvPGWuxrnVY5QK4X9Aj
/XEVX/I5u89K8+BcGSe1CrJB8N24OwruOP5ORnsHKpZo+SY4L9oDM3S6tzwT
AtEeBpN08PHfFo1jEd8lT9xlJ9qZOWZ/+LiErW2droxgYflvbJBEDCZTEAOl
j6ajpcbOcNsqn4SUy2SDgiB+GeKcxc07zjZGkx5j/x1BmCy5cRCfMyFRP+yp
DpoDCPrMOa1fUoW+2fnTPplyD5MuqTSFTn0YwqGYczljztdFwssQbymJjbQK
+3JfDlaOgtLn5k5IJl8VjlbxfGtg/ng5j63aShS615GaY+panpazToTJi4nA
zdKIGNea+uOL6Y+6YC0DhLO8e3TGlOCNdyDcgt5IRbOkpWIaBmE3BHThxSbh
C+EbqkPpNgXKbfNCgxq3iIPLaHJbeSYDnrnpRPBX8M9ne5r7Scz5Uj6jU/Fo
6+DKuSX5+xRN3NQyOMOeCWC1mrTrTj6B/xBelPzuXWS655XBoo9osMvBMUvS
72hyLNsQtFs65ZfjGpb7asJHZlNCGLc/pYz/fOtrtO2VN0pQ/NgYhHOvL4uF
4os1XHfw3XWP9hOJgoNMUP1doIPAq6xoJdcNpBxPetoEuao1YmlEYA7OsWZQ
b7JyyR82MV8KSi++Ad2dnVtxHQG2kFOoR9UBKIs2Tu8NLOvZQ6p6ARctGzUW
NOALktjhF/Vfa+AHtAHpyntfJlxxSYz12ZYeiKZuTmZYZKE8G1kfU01CWZ3P
w9l7IQC7bN5Al1Nn17hbGfO6gNomjAbJmOaDcLpgwPQN2FWgB0Vb+9sYjVIR
czYJDcQDoLqgl1y87SIgJoby+H69fFI+9bc8xR0o7zeZSyvjOJNs2tBaIfug
t5UecXSebPUwu0n9huBe/FdGF9PrbbYJwoLvMWIPkuIIdODwlQ/dmmK/15Mc
dIUEbPkgOxsnmrQDw76RAQTk3fypkeMgdRDA671jll8MBwUHMr3UPPp8WZqG
ZQuPlUF7TF210XY/ChOjgx04mezXorEDyf3YL4vWjLBAjoGjdPZJ1eShHAx2
slPWGO59Z8AQE3DzUv/sevUSmaQ4gEhGQWrtPPC/u7NdqbSPFVvpGoCexgBZ
U85/ANq6nukJTKD+t1rxPJjox4SAxv61SWbyFVx3gATQk3zi8ULpL8QJdVo8
uSJfAUTgZ6AhInNI1kr7feXZHM8ejRi/PRvVgT8HYeBYWYIZFY/ZjQwKtoSg
D8j2hN7YRC5qaBq7W+whOpW2Ul87yQKoIIXMd6tL92bga05KlaaBeIl9RLfw
eRIvAv6ZEKMIzoHPO3inOsVsmj1pAkrqyc4MkAzYTmibEoqZpP3cs60hF004
k5CIJ3m8V768n3G/gatScNaEQt/+J+nAtehBGAVN3++6oGvb4tTbgNuS7IrO
8xhZvS2sJ4DkBjTYzzK4MdIQB3hXG6WIZoOI7EwNFFIZVe9mo0kO2VgEs7YD
bnSQyhid6N8szYZrplWFlyDPT5+4hARR3F9UvD5VL4H+NgxALnI5D5lYgom1
X2ku0krT/NV7Fx9uu1FwcwsPlj03W+endVbV9uIb8uwerZs2Ju37mZVKrjDC
haQdgORC8VAe44bczTDqWpwVyXZta113Kx44SdwJdfHbVmD8sW1fuNb3Tzqt
ACk9Th65mYFnteNogifiXqK0VV2T1LAjnhHhJ9imLqwy708r3CSaQN9vc50z
5dlN7W6kc71SY6x9fbTj3VG97qlASDubO66jdCBKidfJ07RyNBeqLDztYlop
aZterUmI0wjyQ27KCXNME1ChVAn3qRyGzLImZmG3dMrRiwbyDPj1nQAArIdZ
F9EwxxKY9vXmlck3o2GlXhdKIMdM9ImsvUQs7H4MThOF618zZufslJ/DANAY
8ZOl2O2KTbzFTF4Uom4vMADHIGq9WNrRGizlHyLqBneiZuL9OpjhCevV6q/H
Uj7/7IlgULJFXzypYsz/CsiMpum3XV/kvbz1oEjAu3Qr6sYkkkU511oER9tL
urnRKV3LAUcBC+CMFP7zFEmn3S/4wf2y2dCStfWHDDHvUM8L1VqxeC6U2aiv
c6VmNaG+38BHFg7UbYuWOJLk+raDfqJPkxlCc11BCtSZH/I25IjAeTxkPBac
W0U5YnY8UFVJ2Xg5jbduNa73kHyRSfskLyek9CYzjZOylsbBqSt2E+a61J/+
biUiG2/VRYmk9C5l3NT7iNNSBgvUP1E2Ifkn8BKiYsq443WIoydMRQpp4L2U
s20DxMh0aI6bMueJZ+Fj4APFJo/IjZEmGw+6B87MNs6/xCYWtJeWkw42x6ky
DujAuowgshO+ztZk9RQg4oHZgdiq8TEy3RIdCOQQ1tz5TSWnYUJTW6GchdyN
XjfEUENRn2AC6QcB4uuCdAPFeegguFS+NAdNlTF5Mr/XDvlyZdWV29o4BwkF
/ndksXqrE+/sLAnyJlkLyy5hzI6xDvkrM5cR2ven7jxYdTWCbl9256PuurqT
ULk0nz60rKLp6nSQ2cOpWja1KqQoX6MsVnfHyeMgV/lKfwzCfUgmpOUIzdQL
lMoBVMWw538ww8koH5ep6aqbb4mHOPrElEuY51JiLc6/0WEQnSENSxCJJvZQ
OudX3I9Ctj9Enjs9Sa2P6xlr0wWBviL4ruNZru1ZQG+q1YnBjLgRub9qGg64
pNewTPG4VI+b5IZhCksiFj9qx3LJ13mxKpk67QumMqVwOV/PcEkp+wq56GNZ
8AxZ9Mte47M4KqdhY8vCbbxk+UnC28hhVsJbIRbzmd5YXsQX0McPFlNSzhvj
Mha+TfiKu+1mEtRxXJfycaQLLOO2Y+BgxEWwg9+dDlPAZ2uVnJP6qrZ4foIh
w3EWt1ty0wRElElGP5YfVH9lsti3+x1FNsgbCwhL0ARs0vD8VDeBnJkk32q+
K6p9NrRz90NIevC/aVtl1Cp6hizONZ4/6U/9QO82xcwv9Uk+sWerq+RU8caa
cx73HIZFOjgrlIUeFsBrdgaRDYw1aG2fC364gFw6W0HL/L6kQ4tSZEY+A0ex
jB57W77kokUg/MvK5fdvux82ApcdjDWzafDHFAj2zIEBVr7rOxRgfZt/nsl4
4xvQf97I/v4nxvCvNweM7sj/ETRWN5XSewOdBshhj30QtwNw94dUptzMnLLs
rX6swSmnEsG3FhEHT/PG+yjhTFD8QO5T3JYVAk/8iryxR1H+MQ64YupgQnke
NZeU7Z8+5jpzzLjNdGu1Ll7z76H8JLGhvu37Td3N4j81HVqCKPdJLprdJx/E
lnmXWFxJDWa9mgGmf6b/1M0CLOrCWvUCxdWK1qOVR8L9FVSspMrwA72raVVV
aloL0wRJDPGvfOX+AboGIh05lYzyYVZ9NUVKOdd5gxUH+eDyUPuCPTnKfsp/
xdsdwqaLZw5jzszupHlKWnPUgcm4veGUWerBj5sF6ABrkTGbbuI0XfNkpiDb
0XchOgfRlqaAy+dG3mqgpZ/EbsELDaOAvokLMCCHt6qBdqll/k8J3Xllwflp
A1IYYB8i3iztu40sy9XHRz+I1hxSQ+fYt5cP8ZJPnBs/9hUaX0ODphqLrdqI
+V5v/BYx+d6PAwQjKcMWtfkbCsiVBIFm++kGNjpMmduW59fjUXMyYjIerUuf
qQBcbB6hNYt7iydxDeGbdff6Fk01ZwnotaRSLdNw4i1GfItzFIrCw5Z3NpfP
glp8LzvH3lP9McFXDhh/+fDE5poq4g4YMpUszPFsYIQsWmCLPOfMOK4qn9fv
I0nIw9sspZBR3G/U3nCUcSfNB17xQYSFximjNvp/606Z2tpcbyzUtuztqw7q
vlnRFd6+s/r2MrhEydwH1a8IgFHZ5sZkW5Rjeh2zeJ/ZvlNptWVOjBkvX6Le
F1MjA+7MS3cnG6dosAV+mkqTFMaBudzViAQS/ymnMIzSorztRepqmxuEMW2f
0iEfQ0Jo4HoB1yTwtzaE004heUh5DfaU44cv8JsNMfbqpE+LJBT0c4GF9bBW
x3VQ2TwHC9PCSES1PajEZMbbM0N1Mm/cC5riswfcePQZll50VYe+bwPaO5ZQ
fjMJYGtnsAwxtYxLVvPz0oeD8JrBWhxFYlu1++Y1LtPuflxOJSM5xfSMiq9A
JJppWP69mQX/YeG2iOv8CnA/SxrWV59tbsip9ibvjZ28eExzKPUktUE8SLTv
SVI+8fvG4f2EZ0v6XKyNlj99NHbB0wyPEYhHwLqb7upDsM3Cwxmt1HeiJV0X
HLT5cxsmrWCsaxrmAHDmZdhpi9ECDAwk4v3kyGXKbcgO526wtYnKI6hNidQq
MNvVlgXYxyvr/hBgTb5YtPgKT5hwtbc1KmUvOGn9VA0Z3qfT/E/Jbtd86Q4r
AWm9regZsMjeQ1ayDB1nhqcF+Wg4T3sJIGw3L4KYxFLinxIuFWY5Kpm5G1re
fcP+vTF+wdBZMGqlWiGVnKxTUrAPBEE4egr0VxtlEjb8XFv6cz1Cb4sAwhUK
cQy+zHZ6zBb9Ki0orY2r8e1GzUMwEsThTErtsJEI+AiSgVJriK9lcyqdZVEb
qHAJUsVZNFCuic8yHpyvIAbV23ne4VGSrN54vGC9UqY+5swNoemC/yKUOzro
dIto+iOqZM9yYeA8jnMp5nQ8kxsbkPV8VwPjdaXfLeI6GDSeE6JDTKRNJR2C
aOv2CZE5P1aAY9UvvTyUAiQ6r7DS2t4uCimV9AUBVLgXrkV5zWt00WZUIHY7
kPpgNI0Sl9k2vduxaExT2UROFKBqJ/m0g3GptfO+GUErOLtWoKL5tr3arYQd
SIDjA6dgrDz5+e+M154rnb5H+wpU1xZNgXvttr0acV8bnq4t0FF10Z0N64nO
MZTHVug0NGtvxq+/f1sYzK5nhRPYiS3Ecabo8vWflle/fLmtkSmmajaI+YRY
2ArqYsDCwd1m2I1QcZrIxtO2PSp+EHfKjtzVtZZk7LDJZNTBlfFoflzVr1/D
eA4h3ctF5rVIsiXO8Nk8YQCnRyBqm6RpcxwcXPBov0rwguIvR8FFPrpNvlGn
MN1qNxg2kPK7womcK4RWxri6UJvYJ8o7cSPeZI3NMxpMD3xqoGkiGHxKV2F9
Eh3yljrN/dYbR/aBTWE3yedkoE94XxHRYHEFkAz+ntXXDt2yjEqQxTV14/OC
asZNpkLpEu2Ij8me6MrGBJyMEry13M8uPTkWcq0i9EpAitXqnsVaMjdNiFyr
r9OYUQ2y3iYLsOlFjlImthxa5jkx7ZWH47qvBdSQfb7BEgKEHutqLK1aKBBD
PwHLBNF1993iGX2apEAiG2bPjmjyIvXLmgOTcBGcn2sQ0zll/lxZOLzKNqhO
oaBoO7vfcCk3R/awAk8IwTz4hLS/N6PGW6LY6Je0fcm1QwVi9TgJmiYGQvXa
5yg5iiWFP23ssEeXCY1EywlvLgiDU1gx2dSsCAvwRbP7XDjjuInzQrXzDARa
dQ9U4YnhzL2h6jzs1CfEWtDVPklahGThQTrhrvM4c/bWlSlrHxxavBWawoZy
hgy4ftmvtQvHgJVv+Y5gYP0XpzA/OrPD2MXcoB1u1Wjqk5AgLzgFwERMHDFQ
Mbx4RtxTwvXSIG7t3zSFjnolrfzPyk+Jn+l3odop2jNrz3V0n+bo0X25XBGI
+GtCxsKIQZ31SP9fclP9PbVX/FQrIdTJ/BZUAmKrPQ29INg8Rblw76yugBpD
sLowfV4xO/pxNVxD6tQC76rfU5/EWC0JCQhq6g3JN6EZFeV5IHVgkMp003jW
RiJlHHSGWhchZ5YQBk5MPvIwxsRsPBGmGiSAxXixYoQynycdfvYuXXa19raW
Gdf9bM115SeO5CRqDHtlczTjSL/iQmWB7G35Q8DCIXSuFbRWVXjpMRpv9xsb
LQ9L99TX7tBEUKpEqBiy51ZSI6dj5+r5Y3VuPnDg53pSRk98YL8dWGerUg6f
+pVMoe1dE1k+2/OOla4qg6teW4heMNzya6ffwAgpT4/CdFzinvI7xmpPUEt2
ddoQyAZaznvVUx1lIhGl4vr6RzagFkwDMraXX6YUPJR0TTowwC/81d/31V1R
MPrzZra+FoDecGYl0BXpnoylz9Dh8OZDuyW3L/tJgSXc/GjzQ5DMPv4hdydI
TqUgq065uwn8pXTAa6kZRW7cRvqull+qZOhahBIeDSYbNixL/GL2pxG6SxkS
RGoLtHSldmFDTfgIlDNCOWAsczYENIYHHwb/ELTrA6xil8GPKyCypFIIjNFQ
JsxR00KD6/kzQynLtSFNySx2iVLn38bBh4TCo5b7UmPWZqZWMUC39kNjjEKs
5r21X8oX/HWsaZ/sj/e99HVEiTxQQkC2vsdsLjAQZTHaSgfYzqwX+MV0M+X6
Tr7va4gGPVID2diZ/R+T63Xm2Av1gqelEO0iiHxOOBvaw3t2cPYZzWi7KE/D
xGos8zFaDEbmuyj+EeXCMXSNawwqH6lLasYhk99+kikouIJ1QyKJTyi0xDgJ
J86fCQYeuBbvV3BE1bPfppZ6bx9OIF5uyQtQZjKc6750WGMg6lhSO+A6SA07
+Mk1Eg0JACTQHF7g2ndxzCWyof1eHAugi8kgIbmLfR+yr/WFKjUu2pdNMHL5
mNh+iL4RTDdKk+jVGtuwuV9+97z8vGWs+DNGZ+eVWm3DVitXfQOkU53pJIjN
1Jy2viLw/w6DGTWy77Qp9zxIPzo+wPCtBvpoDCn5kb1sEGGIWuoW96ZvUXp8
cp5ZPW+mDSDEhCZjNPf9RwgufZsAB48MRH7yXMTPI3pNhDGQg7YZaC8khsY2
qgUkMNoUh/ZhkpYsTNvFp3+O1Rh7MSTFlOprgUUlr0isZB/psUdsMEnswfeW
04QGSQ6VXPoJycKpP50AjpGQJ6cZZXuu6uBORiLjbCuIyY5sy0YJkctfmfYd
9m/RiCjwF7T0dmgu3U+F5KULBiP3Dmf8nDGMLK6ojF7DvJvvhQqPKP1Q1dGv
DOlkCwMCIPFgokUPOQldlYMyVpsIUXIw1D25c7xUMgHR6nIx3HvdPR/CWcXr
1wPgMTBMaUO/VoRspRrrJLEAxwu420DZAoG0ktIlzGz4fNu1m+W7PvGrvmVQ
2qQBT5GDCIQhXryAFOIPyDaVOppQ/SY8iewLIeOrqKVRXSn9s6+Xw8Th5OfH
GPH/Y8PxNwdgex6/uQZdit+mSx5uYhnujGCvJ6XhkFUxYo2NgxwGKHxPh17z
zs10LD/i/6uz2rrbcLt/n+6T/4cvih5YHHBw8159NS5SzT9VztFeKxTAzDs8
orfoIy9mWY1isQqxw/euZecMnRDWv4iNy0AG+l2afwfLnp/47Gu5rWcgbtiz
n6vvT5YEXlY/SvtJ95zSWklYs3sKSMCZdz3iKhGFEDIkZrvNto/MdYLhKMkA
+ddCjDDe50J0r3NBzAaK/pN8/LFdAdK+LA6PGmWZNagW7hBcTu8C1q9K2EJ3
8uIJQNPWYzs7i63d1AF+Le6wLrPXN0cg0WFNOcLIaE77pNn4xP9sNrfZoqq7
cK4EQraweCAnHVuXDbv0/pm35t5Ec7dgV1r1AfsNTMlaQqq9Tt0awwHR4y+t
KMRSY/krm5G8gVlVVXv6o5FXCrcgDgRjXzpd3s78zuj6XsV1JUNyQE40NLVU
DaKhEe9vwdlFrJ6mf6lOS5iL4dTM1wlWbz4AiIK8yiH2BQMULF65P9pe1Xfo
26Jfw2OmbDKYRYzxGMzG9MobSVBh/SqAwgj92fkjU9/efafQOslbVY7GCIsw
H2sn2+yY9tq6uOxRP8hl6lXUEA6bG1v73QUsc5GpnU2OVpc/0jZScqPz+SSl
ongnEpvhZwpJJtyKBfV1v6SNcGdNf+mQP3ENcgRQaaNrgJsz2HnIRCq1/1P2
DiexgAh9q0AE4UXZKus8pHSNUNEzJQrl4xJYqEnuzVc+2lQVBE/7/HlRUsvP
3uZcv7BeiguIyhZesw/LK9VfgeXjrV3ayIq+8ceEM/IhOuHTTWt3zkogx//w
WBX5v14RycMr7GrQp/efQ699oRnb1wi/ScHBiJj8uQlUZClcuRH1OxT3ajuT
8fYwF33KM+ZAR2K+vCmV9YCOiCoqp5gHX0kF2s77bnUIf1FPvSZpz4DvZ/9K
++zz38/so4x0z8n+5B/XGI2t5jsOiFh0px9VEWNjuYr+W/HLfcXQSNYfz3GO
MsRVm1y+xpM7utPbbZfGaylkj9oKGrqgLwML/kCLupNTRdahkoVrbMaFVzZR
VcFEDIi9zF7kqthMLeB/m8qi0i2FF7sjYrYsHoBuknFTRYhMd7SJMIMN3/yh
tkLIQ7iY6cC7mPSFxKJQu+JHSl4X1xsr9alw6JMVAG5TCqMYtWBGJoMt+JOy
tqO37Lr+7X2eyJEmp+nVFD4aR9Fv0onNpsAT5fiZ4E1Prc5TPP/ZnbAu+eRR
ys2Ka5Z+Qz5u2ItKBtxYy8bGa3gWbvPcZT8VDJr2rWWEvngQvytul0ksrvbp
NBaHV6QxxM8i1Mr1V6tjCKqy0O1PJ4viRXcFOSPpUfzpSDoRyRXi08LTmEDc
1fMIJzAv2uCG5zyyxfp0ABLvJE4bos/w5nhph1rTr9Llsq49oU5cAJ8rlOeq
K98OtExYiOCfjMH7+y/+TufQNtWjZaT6wSdrJu0mkQiO+x4wJVd9erq9dDoW
XFGJPm7hYVCcW/7cx2WwIesHeCH2P3GlXe9cTiZxmeDPvntHn1ZGkM3UjTRO
vfr/nZx0ZGX+26sO0Dq3ivNXEEFRfiVC1R0KACofW4vp9ukMQB6mgFyy3J4H
TQaU4A9Z+NIVIQf/IHlKjvF5Cx9X+yzMP6oZTQrGsXcwWu0eJFt0ZttVj+yZ
InsleWEz0Zootre8XIZOi5u4WZbDSmN/XdkZEHqrULTESg3PLFOU/PsxVHiU
D8nsQsvGB+VXK54RbBkVvP+LGEax18ddwQX4Yqfu4iBjhCiDlojRC8fUXwwj
YwJegEs572L0gdv2NmiXSsTLItQ212tRAmIHkImCGPKZLsfu+fguIISFyydH
xdZjPHCq4ejypWO2WTeaWmx+UYGuxMMSLhSM07tMoekntgWdCTpmVT89DkFz
5Ex6OO0J3X5zRKiR5J0RSNxS/JOVZuVzey5NFSeB0cUaMHRAuocpqISWOYOc
/T9mc6JsCWm7LlpB5KJX98adOyDO8XU60Prv2rzNrcrFe/jPlkR3skjydNN7
Bcj9ZUxNZAYw4l75gsWYyhF4sXw5jLAqaGjRRzYth2SEPbFNi5Eua1+watYF
n5pBOxZyeaua07eFiI1M8Ol59VVeLGjsuxLdtoLcjmhYZ0aZ0TrmKEyCSkXR
+RpHiZOq8+hsLZZBGarOv/3s59ckiIAsEOwWsl354X3b5tl6nWG1gyctCAnc
Vds7/M8PSFsQl4OCyQUAaoi5Zr/dinEtd2dXzuX2++vk8W1thfYKavcwz0y5
q1SSw4/cGsln46O0w8uTMP7lFUNMuhv5PhS3wSAqrQv/m09sqaitLBXI7nZN
xq/aY8DjPmXEn+GGpsJz5VA2EkIdGS0Kv6yaHQZefqyeNQ7LI22zTTUSRBdc
tRuGHapb78M/lJbq6wyLTXNAVATrKajETCUcVKl44AqJLfSaPhtbdMM1Eqre
e6ISg/4IAoOf2XlMan+hx5RJYhSvZRN3+uHoLZN8zVpOgKke6jrC+fHp9JWE
zY7DKVZ5pO+DwBNS9sJhmOFjiNX1r2IgZ5fbASHF6RO92BOF0vkT9jVYClQN
5h88kBt5byZGbtsZO1BCrt8pU74+gO54sD/6FEveLuKE8ffdC8szUTNrOKjZ
ezRHx68kbD5ke/pOdNgZbes7U6+IhmRd2bLpH0kP7YD/UitMlAO6RYYbZjKh
EghnVv5C5nyYHQU+S6LDaKaZMhEBPM/vl7zqJ3snQ8l+0DK5CTjUJBtmp/2z
g5Yh5mb0DVoHwX5OKDSbHybMf0bT5hPApOurJNwMJ36EY1IKsCkMCFyfVswL
HdTwYhGw0Z7igbMaNn6otmP0qR1f5VhAGA5ncDr7M5D1jCUlygF4PB7jwaNs
ZUYjafLAcwzn6oe7e1G/wBruR2GnfoEMYaouUiv8FjXU5OkJHESBejLjAs4T
DhqrTHnlR9z1BJNMODYQACdXuN0md7EvI1U8TcOR/gJ606I99n+mygjZg9lr
Lof3RoMTcog8xNUc8tkHbBxK6QT+xsjgjcrejUDOEsTDV2ThXvQFnuckGorx
8ExGnI7iZCNP1IJ0aqqsmxNgJEJp2SuqVdo+QAgm5SXtYEXYnYaCZxvLArFc
nbkNdqxyb07n/kMKXXfItwlmIPT+cuJaGsjXqR7lDBM87LZd/wvOZ5+CJ34L
R54fhJml7S14+ubreeLWpf1texgEC9eNLkkBqT0CxXB59TaXkbVx/j/Empvy
m3H2MhLEz6mfMM6SaVLi9bgwcK1l1l0sqn1edZIc8/79oB5BsykThfxZauNH
RCUgZMBT8dyyU/GEDlubpnajJSPzBBfUYC6sgPQ6efH9MOk7Jd6T1/w+hWKJ
9gQx0Ubg0auhGjjZFBgqjuRfNfiyYpeh6E//TvWERPMvDVc41GgIxLI5zBT/
DSvdTZecgbvZnuMHMIw6e0vU5Ouuv05XuG9/5SFiTFEu0iZlXzu3BI2cI8Ba
q/B3L0r+2jaW+4//yeP9P2MZO5SFBhUBLxvorMkeYbO+wGtdJFiT8gkgAcJq
S6d9aRGw8Av0bCszbaM3N3IMGjQqx/vWT6QsC0QmQ0yqzscOMzEjT+YcVC7R
k6jZzYUg4RgK/2HMjdgwFpgs3eU7fhN8fkE1fIp5acBm7PzGjc3SrKc3JZog
mEx9J+RhiAO/v8/loonJF6PCyOdwoT096vNDdgr3s8+4DDX/BppTJ8RJz3Vq
ctEFz+anwK9zxScjoeeBjpzDJRljCmYd8MubSOb/LLB3TUzYAk1uHWFM2s8K
ot7RaoLdf3PluWsq8j6d0v1MFtRUUZ7Lfn8pUY2BCmUuW8QO5xVLRy1p4c3O
ll91iHWXEMGFnlzaS1N+4M8zGCk+FHoaSayMfmT28YLlsk11myFlFWIvY6Ok
crbUTF1baZWj1F3GWYPzbjfdclgF56oABYi+ztWQcpJiYO44YCYIE6uaTfbP
Sl9RzwAQXDiKJ+QwvBBN/elGc/N1BCVziyOkLvlNobCvJoAkw2J1gAu2urjt
/45fD3j5MlWgmYGZFSXh0izJ0VxI3zVg0m8kOQp1SY7HoF6ko4A7aYWefqkm
cTqBEI+TVcFOnJBQeWjreoYYRyPkSOJybgyueQyBI5PwAwynFfYqkNMw8rLC
4o/zfS64ljsQZU500Vr3UxpLjlENIzikuw6bVK1abMX5I1RslbFs8Hg5n5zD
o+irZsa0MD6siV09dqVbteZwpdjZTcppJK8qp1XQ4ujsSiztxT62YRwNwz2L
fNjMNiNseFsQTHrVZstlVCVbiAJiZKiU9Z/1rpwT1kMIZ5vwOcbpuGc3Zn26
xujJ5zbE9V4h3xD+J+gwkos21CHmuBQFBknoCAXe/G+1+rutpgyi6UIGWbba
Thm9NzYCqX+rAGII/BXxIOfXWTu8ZdMn/woiN/UcStL0fAPYHx70+3PeRItt
YIhjj3rZ+28BNbJwS41sOtQk7oaKDgbThhgzZ0Cd1ijAXXuyUN9hv2KaVloe
Ck57W+j5ka8Iwz9Ibc6kqUwLkNEDYidbqhB+PfU9JnFDZaIhZqmYqJk51uIK
o2weMPKT7XxMij4YDpwbwPURkoXLhVZ3NoUcqU76XvQ7uSUvn0FfLr3cFNcz
LxaGb7vFfWmr5/VekgsKxKXyrQs3k/ZufN/NBXt+JkAkDd+SlfkiUsSGevh7
CgBbsLQ1qCbygEBq9nD+4TY/u/VQ07Xb4ztuVJgB7i51EDfnr5TGVsr9WeAa
LD6YqsuXjtQ2AGsgEHUNBPbSde4L5AVDLmzhXcJU4+ZCrhGH1l3xt2DEqtVN
AryceK2CGI0VLYioEf9EfFqKQQwNEcAFlPAXZKt+Q127E6P4ik4ERQAViqJb
QM8ikzKchk8beeijtqY7ec98kG+O/DLScW7HRu4PvSHTsh53d5eXQeiauM4/
DbrqcNR7VHjR0Uzf9NklC0YBaT1KupKvCe7nsv1dkaoX4k+CfFAbLEHGktAu
noAHX4fM38WNJk4lHNca3ckj2S869+CfZG1tMYIRuRqNzf3pkLr/8moKlo7E
+frwm739D7MXmN8yq4OpuMZ0amLzE34BxSe9U+bzpQoPkSixc7Hcotpz2wrR
bVX3gkA5ZcKtQO9eTeXB0fo4j++90vcyNgh7vYd+udukyGaTCo72tvLdErNy
g68gLtdcIhFRlGc3ENeXrpKw5hR7BTbL72dx8cn+MQb+1dXPET8soPdSKLGX
4BGhxLUmOFdYTwPPZbPGB/Dkal+oOo+lQ9Th2vk3RWPSShgljR6uvz+i+YOE
ytstWsdl4MQqnL2VLk12FCrCWv3NkKXNCKZL+vTF9A5t0DFu7dIaE8UnMnXy
8Yg7UngUWchQ+d++AmZRhQwIBCHP9E4rW20xffP8af70p16oHYleYLv1I+cK
1ZDKwvGSEo2u3rfwNR6nf1BA9wxqVPNmMHtpgfWbvtRVvDrLX3Xqwnih42En
ml4lIESRarH6bRlAR9k01UiXmXwduRaGFGQN6TNsQ2+TFtgMvojnbO6hAviO
NcFm4PcyoAklzzQUbaIRXQOHG7usBLr0Gc9IvbPlP5GlHdp1NDJhPyPEwbPj
02d9xsJrM5/wiNX7EBpmLLzECK56IB9FTQc5JS8VpCcivjMSqydnOEA3d3MH
DKStXGECOGFzZJ2pa7Ed0y17ulW6kWo0nfinU2MQR4PzJUIc6ho06Nk0ATR9
97pN8KQDhZqSGMrstSvkMpCxzPOV/dLXu3jYgtsblcdNQ0pw4notpSE3ApYz
Ha0Jj4zTkTFZ9ic1gvdYV84Fa2/ArwnayU3P7ntCzYMUckxa+IAwkPbrepaC
KuwOpmz3yReVPiKlKhd6IJh2J1DuWgNkPN2myzN2Fw8MUrw7+uIIr2IlBDJF
vtidTmdLRSD9ldpo2nypJ2r8s0pfWwshX1KGt+yOjNd0AvFU95Jo/LETlSLp
qOrR90ehUQuWnbbKpQUbn/886sx6uKC2ebT9AhbIOtUv2VTYBwypoArJs6nT
RkUaef3wvcpeiYhBatebnBHyySkQQIihpMotSPafNgF0T5AGPIOLr9wUTaPP
ApalQ/UMQ2+HBvxhfYYeUIsR5csXcvuQkom5fMhBHgXojdf86SKPpo0oF3j8
099lg321OEt8YpHSqTsmHe6s2l8FNikusLYuXs22jNlF5f85U1VzNz1ge8h2
s/6LvL3oDtOtPb4eq7pf8v1eNUb1ly6nxoeZSPnVP3mbbIWqqoH0yYosUm/T
yXTmyNkgIDZwmLtNzb+OakIfJ6/lnbkb0EgqMOKjSFvPC3htc9DuLF168MT+
2++Bzt2g46gnihRJVT44+LKZOPXye/shG9IICrz+kT4U8kkEIt0CVatuVyq3
k/6IHuDfW0yNLXy2R8gnLR71JUipGLqkDBIxv/b15iMbWpP8YA9vRk5+QF1Q
p1FRyKhm2EvOlx6a6sbAXmfAFd8PaScMusmaCX2/JTVANfVXJuAeKZe+nXDU
tk++L4wVKutV3jSHcv0YTR6PIJ9hUpvK/khjh/yg2xQXpBq38lgOyq8xBWMh
qmkk2PUZHLiW2emvjf/rpkuBMCDwReo1THeYMLuLB4HJnrsBa9bpuAH+xzKT
MXoJfV7z9aQLPlcSrU9M8mtm96ZlnwvlSLtCEADMTTQyPHl5CW1WIXL1dVwD
4N/+gNpQgBVE9z4EulpuY/xKA/fG6OLJNqabqQKmYVibpAgoQ4UHsRT88BUV
Yl/h3OaQW8/+g7W7KRmReHwX7i2FvtCy5daCTz2UdCW1qJdNRLra7Bjmzqn/
DjQCoinbxedYu/i8M0wTUOTmfVAqJH1XsdPO2VTSH3pU8fH1sohqDj2rcFxp
r0i1C9Y02jIA8LCp0T6sfGcR+FT4VaL0wAki6Rjt9/ghurj7BOoBqFoin8K0
wjxpb78kSEgNyq1UKuTrhpdxMe0+axseyv4CaPCDVLjSr3gd14HmtTXkEhOK
cK+Sp2bCS2GgFliPi7kftXV6TU/8RiYuAzRHxCH/bKLcG64/tqaLnmxcocXm
vYL9s2eDOaureKlFI/hirtnUO82p2j6JbgmB7KZiccK/Pd4RlWvfU+wfXv/T
HR6dyeZtqvwbX1CVOTAADLpQxZaka418kvNual+2sRjqXXh6UdcNvQ0dz2Dy
lP46W/8T6ee2iCZHLAsAR3vIUPVuIVQuH/V4YNAg222IPfFZSk3Bmzgpffiv
FWEcezV6vDmvRPCIhjQ1EhUR864WWwWmp2XeNQZuzFdoZK6SosEgWoRpSjOQ
br1ttUhlYhce2KPq/amPqZOwvIrTlL3toIIv7uWlu+V6HSjqfi+xSOVDxAKD
uLB2UrQFS1GC6LCavAgTjZYiFLLfpqprJ7rS9ylWymboHtlFPlkmGD41hHpV
yfV7355U2YGx7gdLsNOZqz0An1G0vmi/OqxlsP9PxRf4eXEKABjYnRwDDfvL
vTLvrx8j0vku7u+eVEyUIckP9V8ZPJ1jNwEqdELKsnPoYBzKuunFdeNKzh6Y
hbhAe3ehx62JW1PQBYMsGdV7tUrg3ErL9WqHS7RqztIQVlZAuyPgF0zIvDjh
0LyWqzIYD4DvtSAysF0LJlwXf2ZFrykTir9Xdghi7t5riBu7EmLPwAKUZaOm
knZz7gtPDBXGfgGuqIbZJG94CpcJ1Lqo6nCjKEb7y7iRxsvgyuVFJdH7vcqU
UDATnY/jlS5AmmYuopU8v/Si5LGwigfYlpA6YPKOLUHW9E0/taAt/jghWOk2
9r8Tq7SZjQrlE25JYf0fyRiq7xuk7X9jW8TkUVQAe3KAQY9r1+IgGG17z4KH
UI18Z/jdXql/SJh7kqdorTP7T4yqtGkx4fgFdo7WwLQODPLjngctHnfce8nu
iRbmMj3V+wOGo7E7eNsYRNou2PiFDwQ7WZ799LCxpn0zbRmWf1Mk5b58xzH1
gMqbL9L+pNx+jsrBvonNLwLW6RCs/d3XIui1JLg6euG2G42FmoWof6+sDxB6
VUIi+DR3DfMUN3MQtiLKqRlrQJ0K+CaHY1vtqOGK4vnwuN9wIabcxHoPfZ+h
4HwjgzAGucX2tlC1bAYx5/iMZVOz6Izlc1Y/GbW8Ow/ms0B95lEKY7qdpf54
IHws3eqsjOty7I2vhBvdAX3VTP7RuYjJQkY9MIjOFUj7tg3oPnzJIdWpEiKb
CSo0m2/XbpfFiKpk8HsbjcJxNxMcMc1yHXxtG0EVuyWBB4TBW1waUj0/zdQg
mUXRZgiR6HC5B78tzTaEDHYwsj7pHn7rMSRsbb4AK2mTIlZGpEdFoC2iVnxD
FZRHxStHWA18TsFEziheVdZShNzhn4X6SpV9pHTLhs579jFt3Vj0RVeI9DWo
G4kT2EbJOB3F8RtPMwVLOPgGg1GDlrEuBJHxdka8GFB5DkwAuOeRpv2H9CJ/
wq6tdbqdzbBMeHiT5M7aQoNJDbCyUyeBpmhj4j3AACa5Vt9K88FxtlF65GyJ
Zcj9bhwOV4mO6jUZelmZDwYUHDAGvn0oMvmU0UyOJIjg4/QgtnYBzMllauKY
gkS8CUZ0tYrk5/nYlpLjdfdL/JmzWeKfheWEQPpy/GO0SfUa+FzbeY+HAFa6
IQzBnptDoXEob0bGt7RQf1Dtj4mXBnXfW/HBgWAXd0bH0LDmdxb3YaGRV2bq
VrqYJuOCrceirHfpPlxA2Xui77PX/+1n9fRcso+6jsdXi6PvxKUgX5i6cMfM
0VAhnxoa80S/NisugLZ34zO7aqySju1Z5dWn7WxdTcwNXKqnp9/GbcKe+hP8
+g8Lc6c9dFVq6wzme5paSToVP0btRxov0th07BgDiNGn6w2jBUi6bZ9XNsYM
Zzzn93BeE5zMpI77e7cEviZpR4WFZpeotCKsn1xY0BMN9dbHqU0Yz4sTDxYv
Ix/ls/Fl0mmsOXstxNMIdYZPVu7fXFkcc9V8VapRty2jZi+yVpE12bSnUfl5
6T8RkmWCj+XBu2PJd0J8IcMTJtamcaNb52UPfwIJ+6OvsBGKobF9V/pkUBwT
NLbE0iixxYAqBJZkcqkn445uZdgq1I9vocy+m8W8jd5cOrmpXun6KGidUkQ/
JnD2aG0i1GDyY03cwribaCiXrKHt4k1cuaYanTZPut+0kRbv0uP+6q/IK7oy
7L++2KdoEwhdjByoAa+jgsdzT92/8VwkkpRfVZBDTiRBwgfGHcaIB4s8gjmm
DYqrC2ix4M7wlSFec/NMFa9+p+qt1nUf9fDXqtl19RPEotaIZzjF/7htqZvJ
mR6CMj7qv6sYaqao0BtmhRE+xdLpJBtGZtrgRE+iow+RTgpiyDa1nTYf6G6J
onibyUDiIrkmScQ9l1g8gaBmNgMpLYTQryvkpLSdNXSmhfz1XoA4YhT8iEwC
GvrDv2FuxdK1Dt5p3NT0BNAP2fcJyHWXXrFJtzarzTU/UoWsJjoJHZSfTlq/
LeBopJD22ugkIj6b/TL9rGwObbG3noak8AYVxvo0RnMFk0W1Lev0oubbedwX
DoFWu0XiKzF0T02SKi9y2eiEygd/37eK8icjYciNSynTD1Q2BPTkR3Iy6MZ6
JB80nDmIeVNPAIWQn6TaQBPkO4zQ1Pp/S6OsKWBMpxgW09wivxScgx7X3stx
zWKeLVzdwe3P41ALFkovpKk4M5iqAmkZU7bct5HhflgfNz6+DMiW3dyKfJEi
9NVwoMkgxY1ocwU5py9nFAKLwzIUkvfsIYPtVv40ooHmznrOvizWP0Yaekc4
S88+CLqZ8zLDKR/Oc2T9rjng7ZcwU8EeGd7ZtYJG+Hwkn4HEqsPGF1CVdfkI
T2jYz6QLPS7FPzk0HyVe6pIDBFrR7VI3Gl1bsDqp8lmtdOgWVtAwdE8ZVpaf
XJvw4wzgJR99mc9B2LMb5zcrHkjSqXLi5KdJh7zlxEGdEsExj3w7TDNAcJhg
Ab+p0EfLUOYfUX4rso1SZ0ZpwRe2/AjyswVWdG2syfOTupn2Nn33dxeVblpc
Q2NOvwn8ZSf91OYmBbfw8hGgGArmo4DRbeOYMm6tVTyepnJh7lxZ2xkd5wSD
7/xyfUWRrvGoSh9XXtZAxaE0CNEUxwql8yjidiI3B04nVd+OQ3YSpc7nvzfl
lXLolDwfzEmUmAzLlJiYaNAVkJQjpLXbVAULceZJd/xK9BFoUc8WXBfTU1pM
Dn3dKXw9XykHXYFRo3zsjPmdVsfXSOabK5cmz1W9mbgDxVH80Bfu77UMQTcq
Nq4DAiXkbWobAXyGdLtt/fW3bbb1yXfgokgatqKWBlhX7qEsdqnt3yafY3+l
GKU5NkQkg3OPEdlytP5/Av8w4rgK8+oLH6fz7cm4jskM4dxXkkjoT5Mrhrl3
rVMQOpvJe4YbO9Kaz0SDywYvBNhTENlZbFsk5EW9kHwLTACHbI4I8Aeztmjl
USLVQHlyisZsoQLVO0WLZU2r34NfZAm/8LjhM+UDQlwZxFoNYM/PC6RxHI9S
5HqlWUsK0YFZl2ATnMLWesKTJsibFmiFXFt1LDkYH5s7/BlN3cNU6PPOPgkn
bMpVecCqXyQQI9lVS/WGaSmnTS04jpmk26mpi4VT8H0x4+uG6nscDsKH+Q/t
koSyQeA3owLZL0n+DiuRTshCN/CgIlbsF9GqOTtFNr2SYy77XiB2cjGyKmGg
ohkNyJkkvJ8jy21aXcNaoW/zTOWu7+tBz3jc4ArN52jQ4hzXQ9EwcZ9UKwg6
+yuBAcFBoI5PK5mvJqKyiQZuqrgq33HZc5W5zExSc1PuETzKTd3pnMPqkMWc
D0uMZdE0/vErompHalIcnd+lWab474/Db4SH6YbSgOodwLEIMJiOKjdtDNPo
1K4DIZ1IYM861e7EfETr4wSILl4399kidxdtBc9am+Yw4t7Y5aEvKMt1s2Ao
x4DOJWO3OdcfyE7heFmg25cXNTp8Zz+6U9eK8w65jNfJA4BUkfg4ZPNMC25S
fCGYGO6cYINa3rOSwqdmpDyIo+r3UxhLfVK/c7BC4Hhh0/PGRvQWPBElZapz
n9QCZfAhlKZSKFPGCEHW+wKDeIRFUa9a0oN3kZ5Q+tx6Ezj7CmN9lPzd0iuc
p5PvQm/tLpc/uyqaFDNpyIr3RXwDIc6FXvz9jlFpM8Zv2LVLQuJGS/KSRXV+
94SrSQjuH5ACdhtEWZzgj0oPX94hPuABmFDxwXeLX1PFx5hojixjxRswNbos
bj+eOrXMuayQKrhkaWfhiWr/VlnMlYrDKPuQJWEy2qgta71ovTtn5KCtWlwl
lZ9rXwG+iqbvUJGwFKg0inybFFK79WXpfw3iuv6rPg1SDGrEK+Ay12/X7l9k
tKWwT2L/WgYB+X1VM1SLgutkHatRERnwMQfZcknrExVABdi8XSJoWH2t8NZZ
hlyhaMQnnuL66ddSF3QFMKDB1Vu2BBVGPvHXhFmQGlpoFkIQ/Dy65C/6KzHx
3occxZpQ0SV3E3tycGwXeDSvAEjRLSkoHxR8vnJZcV7t7EW2LnM8HqXHBEx0
2VpjuR+esLWU36kpyTQsGPZZ4KhS2J7Abab8zkqpboTajW5q1QvVAg383tOZ
Ssv5CCswnQqu/srRZH1SAMRYmlLR5+mm6k+dZOjaJE1wjirdGJzAQ8BjtCLI
ZHq6Vp6B7fO7paFeCEdkd1X3VtYtF4uva+P9kxCGuKBw4gwhmOqrdk4Y4Ums
Vws8Fvd3hi98jBBVlQ/RJNZaT3myV+zu+Va4UHkrclUiow/tMW6RXFY4iwnA
w1s+n8xSQaRUWGnefqLhWrMo8VVkQFSKdpGwheapd9hqSpdTryd4Ee63iFCg
8jPgW9dtc5qTiKMoGnaRVRNEnuWc1B7d/qStha+VNxr3F2rVb6emrC9gba3X
EzR7fQjQAP+t16lvHPio7FhnNUlLyDRJNWR5pZJNG5KUj7H9ftgoI8x5/2JB
1BmZuinuVialEgNzuhdGPs+Amz5cj3Owi/9VEqE0gi1SdRb5GG+AhlHNDgNr
m0KkKgR28AzqhQmTt9EHoRjjGWZc8jMo5z/G2WPij0OqHCkfkgoJNJMfaTuB
vi/ntubGDFRiGz35EBxBTMplSEo1xBrDgWf1Yc7x/5c98PbbOyU+3xm07r3A
t7un8nvkSpi+HCO4ZZ1P5aF1moG1doMRHAi54H0HgNBk8gkjlvgMyvWdGo9o
FkF9KwNEnL+vVEnvDujxD1POiZOUMBP7uIwruH/TKJRpR52yleLoQLolgJ45
IYaTqpX2t3EoHO/L55LW0S12gbuXt675chkP/FEBikUN9o44OdfpRxH2QaKb
Ti01w7vOGf9YOrbbdkoGaTc/rVbqSh12HW81pucDeUxRP2abC1UuEYhFRBa+
lAOQrjxNvf+DduN0XwK13didWEueyBI6W4RiVbwfxPmnL0XfCHM4RoegEc4O
DuB8DqgIgaSv/nyV3qaTdWuyxvdI1SRoBRkPlrxykN7kBCME5O0WmwqWJqAt
kwqd2JfJw8KgVgaKTZdvDYtMhLoQhuAF3HKDzebzRH5a3www7xpvbGfiU27I
w7b8ZMUzqylHXWMD0qJI7NpfcnTX/s+6Og7FYO9WCQjgVAF132Ajypq2ZhrG
mlAmpaLWNKz8X1XIm5/Uja6H19IUh4mJz3pd9ZitFSzHrK2DCLlWNtCVSCaT
cvPd8IDdiiW4mTfePL7UsUsTGWZSTLnoWZLywVbyznMQx0QvetC4cdpMwemt
0dsGnwyrQJcTjk2ddYw+6AUo0XMK1adiKXheJI6hOVV9GC9Sqh+1YjblMKUN
HnebE9eLLC845YPpYrBQReVyNUIfIPXfG7RGqAHVWIxqax2VTj4TMasBpvGI
IOgGG+3a2SkwE6+UVMVj44q/octzARKsnL52zdPcoFODEVt6IEvREkp3+rht
NL2POuxs+xOk0ggpK2aEp4iY9uaprFlDew5FzhBwKEBS6Mc7GrNrXVjvGaSL
I+ngZTONMU8slS201R1RUzDN0wgKxMHNIzikdNbsEQ/yWyizPSbecxbS7vse
Ccr23+Jq2Q/WSvvobKM/u5Xx0Uf1PGtGy+W/VokKPSCD4rPjfBYY/N9r80Ic
azZOu0r6f71oGzPuOE0/V62hLutQBplfGovuSCfU/MzF0e6T0DroTBm294Yz
v8yJKEb6aFGqa6a7GWnbFfdb5BRxq2twORVo/0uu5VQAoF4FKs/+URC4tiIW
jaEGLDUxkbW7eWitSPDqSOzhY0FzFwrWuvnUiccxWPjE6OILBhaH0Umcqapa
ToqcofuXF+SRjIgfwl08rsmKAYmY0ZDYq5U78bjIgOVIYfZRpbgYS07RqGIx
xyp9bJM3VuTyv2YF5kGbX4mq+NTeJ/H16VuJ3dvprkFMkW+eIHLyKPSiThQp
MaYZFD3I1TQyNl5m14L1ryy2hDJmvMc2JSyoolelIyLQ+Fl+gB3WTyDvssXu
CIO+LRAg6zuEf+IYW9jVT8STbxiqqLo34vAWrcX3Kn4HnGLiHmkMdBikBSvu
dutYPdu3UItTb80pePVHHIIDD2/cTskJ2GoulJJ9karq1Jy/K0MNxPxwr5if
l8wyKiXdImNhRMZ6xPIhZbc/uDKzm4mhbhiZGZmc+9S4vcHVsdFPkpiAqBT/
pvCx6POgBc8f1VwzPtUwJVa6PFp0pFkqP9bokGGQYKNaqeEW389+zZfBglkm
KqUGRT49C7+2F6F7fzWgJtjlnjNp0JjgJHX/nF9UxVPkWVBz/U3ngsICOiOG
jmRrJ90XAB/e0UhERKD7IkFOf+m2WWS0mwzL4BzElMDu9sr0OZ5imaPOZAWg
Ulae8r1aWw9V1fW7vanCUtoaiX12cSkQeR2QxQLoWtb7Zz7VUsWA2B764MGh
Fyy/IvnBaed794SZOieMlyvD5+7S/VM2IRTSja13IjmhZPbMRUbGTTWSkwVK
P1s4oDBA1DSaRQALU4y84ziGW30TqOQdnfar0E7/lJ55Kc3x7tV4qJ3QxDCK
K+QwzHEjJ99WdLTSnEwP/qjExSqocQ0W3+1ZLbPcg4pAzNvPUNZNFp0Yv568
XU+Un5WzedpqTUqbt39p0KVsF4+2I55lo+KYTDRNvRB+egqBLyUD8y6Wkw2p
ebOdnKd8p8q0nIihiXCmxdWDyDmPb7zvYw5+6hEgFviz1/bOQ2dLAfc/c0nj
TwF7c+8NJhSNiOt+ShDaVBmitF/EwO8l0VkldjJ/S2KadD06kNyfCvn43KzQ
/Yr4xHDrQpdtqF17SontvwdnIMKhVQY8mmWCsYQeZe9Cr3vYqPQGE6EnWBcn
evqlTl0BZNRIUDcFRGZiOLcgmRQEawotURRvDZ/FhE5mvQX98mN43XM0YdUe
nDjP4ZO+V/kB6aQ8PtiNIgDj6DVNxvo6B3vtbNqDihCU38K4guWQOEGbzT2B
SzDE3a31ErQ1slBtdYtVMQ9vD0pa1R/bvwMO9EuBY8RpVnlaLrycyBTZJ4je
CyeA/U7gqZFrxtlDjfVcH4i7Y1zkyELjaBBRYHNwa1pcGIkL1YrnUQBuCIUy
XpYYSAbsXymdZ3waam0QDmL7iNwCO8wDqCP0NTHiUfrNB+AoBG5HZeQfBG6K
1W+urPF9hEli8ZNNoEyCNSQJZyXPSjam7onkdzVJAx6oeOvSIgp89GIb6ocF
eSfAUPPJ3NRysGi8jJfCCvmX+7+BbWQrvUpfsdPx5FpqEvI1gGGBSDR77hew
THXrxLvRh5TRch6ZLMxFM/tWrFjvMx/pPbG54Pa/US2O1wPlbn3/q0Lw/8s5
UtSM2w2kRWJmBo+zrQLHxiiwiApc6Z5w8ejNH2OATZlSwqedJJ6ND25p2KaS
m6vQJbf00qg6AxqAWsaLSVHUHsaxmiJWXufVGONIYu6q3OaQdUaA7vqR8jC/
XGHmUxw7sj9kfh9TZIUmHmVdAWQNIF7EY2xRShverzgcMHa2hy+IqP4B3ctm
/U5x49vBevmLdTA6vg9hHFIa5OzBTmIPsjTF0NK6gKN8dIKw8CmpOWJVIXgg
O2sgnw388C32LHT0F3b0AH7ayWW0xHyaskMKwIRgeMwnxkGEs7C7Ld9ssaE3
1FSCpexLafzCsgzy0bM10U+59fEWzV1oOdfgEkBea3AMXCWyUMA95mhd+sZf
cQhyHBOo/KSxSnFR8myNoCoS+DXEcVNK1EnYvA/P65HoobTLNbXQnag2Nx5r
ygT9dwvNBJnbfWRDerPaS9mSqBVRwQe8JYMhxek8Qy0JptSOBXlu7Q9/MZC4
t5wnAfq0+6LdA+nrua+wMI9CtrprQFr1Qgz6Uh+LvR8li9gB/UBGxuiW8DGN
IhvNibm4VZ6IFvWi9M6KspWgIohkfqXSOJspHFh0VAkIECq8QtuSbAA6/PEz
TShTDFBBgy5tVER7iZX16mxVQNjOFomAMPJ2ot5Kpd/JU5pLDslzMTWCxYl8
5DXtxGwvXzd7HQyEnMAUedWk21Y+UGFQa4xLzXrBmjR5zKzveGdfLhzoYkTg
40H4Vdltsyqrs5zM3fjwLdpMpFIXYngu27BtTAprzcqNeoLQATmucdYVykY7
UUws+zpnQe1tx65YqYn0Jz2caTvYAubl9yRd9RocawfMNDQVkbaKXQxk2FmA
jA21crCW7m3qGR4P8wR22YIcdd+/7rMOOlsEithaae0ryWTBiv2LGgT8MFAe
yzLaZway2q0CNeXLGd04LMKOodGo51A+D3z2r6ZoONF8utayZtVSfINIDrL3
Y6nPiCP7H/XYcbVVWgzwFgg+41ZuLnfqQbPmNeUjRwd0857c8Zd6kcaM2Mi7
0wZe1xU314f/fKayjUPXkB0QQ0nyRKucGaPnq7F82pXr5Dv4lrJvo9BlimDB
b7tkTNhG15aQszdoBDqRaL/ODB+D0sVf8t68FHU7JjK7edHjdLmGykbq0PbJ
ytM6PsY8ZjdMLPMxkIY87JdMTvoagGUIRlbHwFWhAtpWNqebfp2WFqmxstmQ
QIaNwW+kATvLwCN0ck4fc9baVknYgjsdSW/Y/YZ06GedD7szTegT2ELhgQfs
DZMNX9fjzk+wT69X7Y0Yg6bJ3jpDtR+E55hj9vnhqfYI8rcklY+mOy0w/aGY
8FwjLKe/Gycn4AOccaM/JQGN/StO2VIDNGOvZRrk4E7MdoVNfcdhmlexwoJA
Jl4cPqu4AooORrONmN+16WQJ5iM593D3sRrshEy0mecrWXGO1tVrrgxcs8JP
HpXR1zgjOB1OArgksQUndIaWY0HLGUHk33GIChFs3bxGFMBG9Bnl5iDPHCbB
cHGIJD9ikH9xAE9YqWnu6weiPJlMr8PRR34JDSsubJA0MGNC2OmlRCr6W9cR
z4lazYyT7weQcjpJcED+aCV7tk2a/GOMe9gDJDnsSklmH1r4+1uQd4rRudne
SG1cly8rUCIJWbHHSqe7S9RI79M5ZHDfAKDqCGoBNgkRNtt/dv4En+Ogx3dI
K4tDKQFcUgragvE1ZXmt6AZUsVY0fo+vO50B3OHktUJudzK4fPm8qstf6fTm
WidNGbvbXQfCujX0VuXHa6IcK4ZM3MH4M8xukvj2dzPQDsdNJj0+rv9jADFU
CSxXLtByJVDRB5TEukApFGGksqEV+ggnMdmu54yQsB2xtwhxpAfGyzxK1bFv
J2fPQeZqjIab1gJr5cXck/pCewojtct7P5S60W3fz4tpmg7Dww6cLjwrm42H
z7Axfp28ZwdT7BPFPn/nz1v/EdQpNyzULdwNObzcY960vCTXhWA0t3pJX7wZ
2EWeQtbJbPVTAuDY9ynxWdN0QoN4NXEAZl7BUzUNVL8MKO/DTBTrzXyCPHPV
Kly/60ZziC/QDNLBPXnGBSeiagYb4QoAq2neBWBl5PciAQ0azceSg+LHQa79
peCeM5LLBWrSpJnUEpxwtKE/veNvm+YbmrUmT8sBiLLQAGxCz5GXi9vHX6en
d4Exr6uncpRXBQUAfBZ/ESaiZNi9AwC9IFUaEcN3vHGcvpg586EicAAIBYmm
Pv6czrr9j0zB2pNPPI/3nGIHnRGAYYTsg+1qXSjM9fUkZmMAZfM5Ka1oeZIB
Z7gozf29XmEJWLHGqP3FEyT2ZHAszD8saj+KvIw8lsdQeLX2KaoVSaLQvsO3
E6N2cAgHTYLjPp3XZ0I51kWdy6+fpES20CfMX0TPxB7IkbmrA3IKpYEJyecT
JjJGCCGantEOr9SkCSUPNgqnmxwRo4qNk2fCzmWPEYVA/Lpq2fO9G77TSMUS
zmeBKDg+BbbcS/JmiPlnGumXn4L0T7aD5joo9qnDYGqAJ3nJZpKHQCdFF7as
mKImYIlJbjQ98D8gOAn6FjHPPfCvwMQ9+BkX/n2hiwytiikXuEaVQgJ/XMg3
0HYqE7OWJz31Y5IRUwtV8r2ir8MyPKFYvuFLGHymG7rgh0v86RF+HB0irxKk
zqeQEmJeCjhLC/YvhF4ggUhBn+fzYZU0jwGDkZKA0LHMCh7O7n1d8UhIOPLv
EY5Q2nDqzWQm1icOAQE7ZC52rDj1Li8AOL8ZrMH9Xn2/iYdicHh3GEF8XvA+
DH6Q7/FMVHfFvwt2pJNqDaySC4DPaHC8yonkGcg4e4cVpsl5aGfCe5X2CVvI
E28IJunYWdaduRVlOE8G4b2mWaIc4AZesZmzQV+RB8opKF1NrR3w4AvWz+E2
8XKUkGQrQX1/2HjQwC70RlHZjoon47MkNhBZFyXheYbljtkYddwL6hWL3DWb
rX60b3R7kyXs9dNd2tEh23ftDWwJLZmCqTxI+H+vuZqp9t5SBnDhWdOwwuVY
joxIHDi8C9rd7MV8cV/qxY3QTzuFsDybJc5mLmQTKPqto54YhNdijMD9JBjB
7HdKiwd7NSr/qILYnUIJwKHgTieUTEZCSIjfZ0n+Tp73BPloYr+T0bxUm2Qu
Zp1ZMqQlXpR0rqRzBaxqk8O3wZLs5kxMFyrBhCkdNd94/fAiLt8DUnSNUq28
lyrhrbN3pbF3Gel/9vGUmeJx/bVLToEjkRaN6g0uebxo2cuATUGZbHVqFEt0
sc/ggxFWGTXQnW36OqgjMA5X99U+JEx3zhLvn0ORO5C2Iv2bIsWBDxyqBzFY
PIzJPA6Vw480rvvG5NbA32eyKbrXRtydD8o8+k/iVl6JYAlwOtyMtQVVoSXQ
7uZ5cYuFEtICyzX098LUcivnEv7LGga++8PEC+bvl683Dr8Hdf1WSWG1jwKa
VDXeHdksCyzmH9LmqV56HqoNftNsSqNJAf5jrQQo7DG4NGWR87pNcgoWfbFH
OEkG06izvi9iynWQTC5AAMRnX9YGyP3bpVmGnTp1uSkN+zBB9IQPjux+a38B
QQHGodSo9ASnQdqzNaaU1e3dLIJAGmypr5mHkjHzpomqOtmoT4Z17vxVL61D
PTgdGhFAxQPYpb38C0ycPXW5SclU47TP3bwGJo3KgEFQ31brWYELJoJFyKbI
/WQpBER9tD7LbQ3W3NCLwsimwO35ElafwG+mijzlCFaISH7Re/GoYfEHNnCp
D/QkxaIWvmRbZio3uT0H8d+n27pZqkSuK2v+5U3f9HxswXsoP1Sc5c2Ia8Bv
xAhNoDqEqy/rR9Ve0ZXUXQ0nhD6gS+hCDgVMFSkw+Suus8q92KwKY/1Afqed
/l6bzt1/GSLqnZ/xVxgeSR3UFvR/UwzXoYF6gEEL0c7ALf8u+/ICofHX/nca
kwUiu+MsjqyzYWpYmc67OdI5eC36E1z3mxbrn1M+IcGXSrcy9pD3TjruEAZi
W/D433CsUZEgJkfYU6tnihYHHF4JRnyZ8X3aGpaScQghXmIcNZpylPQpw9AT
l0WU9Ik2t07aXoGT9qawTcNGatX9jg5E2A+9lfwPJl3nS1fgpfybvvGioN2O
BPvIxTxmB5cLN6wlRZV2HlqOFUPb+eRk/ZU3Jrv796inyIQ+ch+Zd15hVmdN
SfUAKmiBp/ACJs70O6S4mTgyrJgIfgF5IVhSisiCYb2DcngioRFUI8OqQg8o
u+y4MYhR+XjFPAncBqYxrUssk0nae82sX5d4ePSJGx4ze5Wf4vqsRnmLruoZ
4Nbtxm1Pcl+GthSWIGYVfkecWGs3QRtHaI3CH6xbAZpVrAUslHs1RTAwVSqJ
M/fE039/iNoHKXawX/KniIfNvG+WVR9k64cs9GjbJ8nON9bc2B/6CdiqCNc4
bLXxoBFzkpfvZF+lBsyDRahpsV2eQZEb0xIJCBfp3tbaB9P5MlOt42x9ly/p
2jMZxL0qWNub5mTH+g0nmKIEzT85EAmynRQ1vGF7hhpEHK/mockFpLPCvFeQ
kzn1SEUTqAXdVFsVedmENb7qQxenABS5GwcYqJQ2I84qc1rTagiQuZhVqo8H
Zk0eAoWIR3EcH/5K5ozdmLV4BKOX3Fvrq3vmaGHuqQUiUHDrlCp20FaMi67D
/Eu4FPU1z5nETQGoyFkl8pppK9OSvzTaXJJD6F0ZzsqqVkKxMEpSiAJhQfrk
efXYKpPKLZ5IL3wORTtkGGQm7EMABaK1YDZ5YYO2Pe3fbMuKHWTLPS2uDxAp
LRZo/GSLcjPuvGL8+SegiQU8pJMxA5iDpwd7v7crGgSSFAur/6YWuV4z5GyB
GZcV06za+M3PatkWbb0ovrIuyzxP+JMXOIaw0/plhcLNehuGhU12viRwlLLJ
dblQkccjlO/W716Olexe2C5dEF+FUI1R56plObx/qPakeE5NXTrQ/6+lCjFd
HQMPysmPsIHBeRYfwOKFdTRLyIEU+UTkriYHW6H8ue3p4zdPCDb59YfCe6Z9
W6Vyly5MhTbQ0ea22Ijf0ASj/uFbz9O4cG1tJVfOGEcmi9QLxJRhCx+LWiEg
8mV3uYRA6Vz3T5xm5zopJ8ZWEsRU2tbupGRzdHhLu7w3Uu90+YyD66haG3te
K24D1IdRwwVxrpYaupUv0cV6Rm8NepCywmLqQoAKHp2hh7MPXuoRBkyFOCzV
/80fwedY5My8OC5J0z0ZMkRaQbfVL3GLpgrqmTbH/nK9tMZ4WuSDPrF3CW4/
ktKfgJJ/K6UegM2LCeVJ9bwrNanSsM3Gg/raqY9Sxo044oP7Y4U0A0X1iN7v
CCX7I93ZliJ0GhEVsTtvBGRUQUkKFf52VO6wgrv577bS/B9z4jtPgADaOecd
VZRLFhTIieyxtGShn9XFVlJyID6hqrFWhV3lRen8vAf28TeNs0VIZOB3c5VY
16WFXYKQjIu9+Yl3vGbqhj9yLpg0NfWFpP2l0OOhA+YzfTHJY6sfKPY7d2JL
YiW+0Ls80sFpsg+X6sieaakMZsROGBvqwKS1zXkVS3Y1oI0uaFSzqTf9BfxO
wXrMeJw5IYLRQW6lZ4l4vlFxxW0AGYSwB+0zsHjilOPUJSg41lMVDJmtx8qM
g6j44I5Uu3lY99fensySJD4HsMuomgRUWwV4DoGkO8Z3JattbFosauF1zf7P
cTsyhlMBWqQRbCAPuU14epI5BOTi7Fo8W12JdOksH8cojT7ENCTNzd2LrkH7
HO+PVF4H9+QaHUbzqLpAZ4gUkjIR6tWVgTjyHCAHLK8PmXNBmCikulhjQKlV
OJ3XRn05Gx7AvhzXDC7uMJRqTY7ZG+ffOXx6cHHuVNCWFa4I5tnUna/lp7OP
UgeAwZwVE+y9AWeGqLmgOJ6vVHCgkdbIg/NQBgjaTa5BpoLj6HTzllPuLhJl
UbS4yR3v/2BVPyf61XTREA3878umafKlHOC3pfOE3nIFKXwMXMsFuDwBOux7
75amDerNrjBh6P+y4uVjaWvR819Y8gCbWr3eg0NRDeFH2CVX9MNJOpt2rSft
U1eMq9hCjPfnawkU8zhGaIWWfIC8u0khUASQkwFlZTOsytJMFHTyzKOIanLK
cljGfJVNhaE8ItGApMbeJB4+Y9nehZSwBu7xkJsPFiDVCWWYfRfG1ONqqY2u
t7NflipMEvMy12SvrNk2hILX72ktnu439yjjDmri1cWo226DEH+tvIac7C53
ss0O83+cFbiwWBfFkA9Jf14AJZALXrWOkJQNi2pJuhHWgNap2BNGue4O6pmS
MdzviWXJsok9NoU1nh0OQOIse2u2nUJ/DjcIooa8HtUSVOC5ZgQ0U7SJ4m16
dxj9Q3ae3utVPBke8LZ9qtawAp4AxKULcu9MW9gploMepgw1F/YKJXb/Rn44
5hDQ8YGXtcp7dFiaQbIt/PWx0ZRXlZZO+Ql/AFZX9q0h3StXbYVe6ziw37Xr
hHvHpgN+Wo+Vsw/3i/8F9NzCD14c9oitql0igzvVMm6HR4YFVkpd2niVMLbR
P/xlYHTjv58z/WAGCh7aUVBPDacFYsyyuPRfsqU32N0kqp/AY3LHoY3HNFqB
3SsOmsmchsd+edaEJfLGnpjBs25zqOLf+mNIMPGvVfzy/fl7BVtFJ6Q57iFi
tGdlf5AnrFoF2T90RFhPMnRFpYstL3o5i9hbL273vObnkSSds1oK3cbllefu
d8SUw+HJcyrKnQI82OWMtqMlGvd5m1Xhgo49NlLMpFaEFxSbEgonIm7Sl6GM
U5cIpxnupcFAOmoGWXLO+ZQQrXYFtWNSJ8mmToD+kQlJWPBDbf/J+QG7QiF5
Ohble6fOLQu/6H8k9uxgijqYMWi+pIBSjhEfCK/CRXAggQPyeWU2wWj/zXry
PFSYHxbcNg91ER+uBHj+UqcT0Vk81S6VBomXZSHC+s4kIQSlfRFtjI8en1NX
4CgjDkBq2MUGwYSLcBqSs5LnB+ycvi1BGB0pmg73/tMoAFYSNUQ3O4pefrey
WlLJgMAkZMa6qf5iOueEqyobS8XvGSZdip010DWiWybetgZ/UmoBvxuhOLXN
NRydghivA1a0tJgvsFqOMrjMysm1RpEwz6PWCXnSqod6XAdSTtEAUoEUnfa3
xGfg/5TvHAELXVj0BMDPFJETSoJccGDW2/iha/LC2a2Je18N40tuG+/PAA5C
4n4nJQ39m8bFEr/L5z9Daou5UfFPoALeHYoEfCrP+sQ3F8yfK0dA1W63LxQF
CXyvjxC8ZceRxwbtUzxJctXsXOmRwrOa8xlRW/LFXams/i8HfSfGW8MbyFd2
DwWx/I0VfCFAdgydy2WW3CEpQ4wkTbN2BOawYJ5ZkQWDFbBqYasi1aKQhDNt
mINqdfbTp6AcZaC5bKPwEEMuUulMcQYckVxdqwV2tB7gAjVbdBXlhGkhgf4K
Cz5/xikqFekeSY8V9QFWhO5tYR8F5yB9bt0tO3fZ8l0XAH2qLA6WNP3pzYf8
dB/cGUmDf79z+g31drxABDG3Wy0sO3dDtsia5+CLxtHW5Dzir2Nco/p2+hQt
zg5F9AYCRhaDIkeq3uz7qtBgaphArJt2B8kM6M1491MGGLpvhE7U2/vAEvVu
xHs7K9yI3tx5pC0tAtpS/bitZSzTleighqlhaa7j/PpD+MsvMaY2/VPvQ7Qo
KPHDqojBsUvZcNPY/Xpdub/Guq8WadAEcsKipjsHswRShsAaoyhLFJ7zR+WX
Co5F14mZV/sXGTrh917TpDRO5b/SYWA4twVgyEhYSx0CA8CNuuMM28+B5cJM
R6tAjV4QlzgjlFZ2ezglaykXrq/MvEzk37AX9n0g+UzD6XvfogTPD2ijnh08
kDbrzE75Wnj76WSk+4lNZ8vWgZ+GJUc5feVdyNliooE065IKQ5YI7l9hHUPp
VTsTk9MTWZWJvKSgxShR2te7IKi1lul7n6N0qV+U96Q3XmAIWwMlPBMe+5Yu
U5BhdC//sGvM/bGuQ1fLQ2316KS2vJ0IDhW7YUrJsL7Fb/vQCQPytFaPDoDR
36uHmgdqwfvrHZTXsu7JzRVaZrK+h0BbWeoHnisbX9r3q6cVntDbcpkVzPvv
Nfvg7KLo7oU2lOAMJKBN1e/LETDP1clFGf1+xpzuUdoXtUtRLzzTLbD+VWPy
lm5XNhVNL2sFijXC1e80YodaduVA4XMmgt2LzP9b0bM5KQKO58ej6x7kfM++
Ga81akNRtiVYuf3OQ86Qf8/EOwsNPrXzoZLhRMkqQ5oO4Fmz5e/j+taP7eH2
fhtKotzVSa+2BYCSOjzoVI27HJuQc2SQj88h0NLYKOUAslqNZoZTLdDBowfO
PI4dQOnOo9Vczrp19OlgHTYz2BmpTnl/BHWuvRIBLsIFQrkvTHrKwYBJKR7E
7Ld7R6YrNYnEkaDxXx8SsQtWABU6ly0pMqlE6LjWxdquVMIV7zSsmv8MHkTa
Qu1xIq/pdQHijzgEY8VeKmgfCtkWzFbNk1NTXMrgCBmfMo4lPot5/Ua5GIX1
GWX7NgKQjWbdDxNKqA7U3qKPOXwoPBSTOBRb/jlXv3U5h5ND2mzuYvHqEWmY
UmcuEpgNYPg8chELO1FuLlKzZKvhT2bRKpj4X+H5aKbWWWiFwrK2XpjqO0Ke
QVzBpK52phffOnhploOa5IAFWlkGGj+kBlthLnporq8ADh4ZgD+OMP7soGNs
0WZxsEG0eVZ3mjqjezgyIbHptTNLbL7KDqCwejsOki9c5FZjwRL1GfLfffZm
kk/p5GjYdat7OvMXlm2P0zzDL03oT6dVl1IIofQLvwvWUNa0vQy//XQanNYb
WIQ0rMDZjs8mvAcL+nVc6XKzB1pBORXyUwA+o+ywFvdYPtFmGpvRhUOG0lSp
xDmuGjcqSlDNw8bD4fVpFOT5iwVzv6O353NSqj5GRIV0gJjTzmvrmWBucYc0
s8iUFA8ca0J3hgefWOuq1kbt8Hq8pOiZ5zmRdp+Y0rB8F3N3IF+NM7LAp4Nh
j+d1S1epWZfkCUXxupnKAU8RPqmRR/tbttPs2JGHPRH8Uh3xmIlrmdCSnPIO
QWKkJ7ZG3/PRp0sXGEKIqM5sF3n7R7FhAzja8WKSUf2FhD5gOwGn/WaqpMiK
mZyEKM9uHkoLddFZOeJw0tz0xML5YIoowbv+CZ34QhaPKOu0+l446J92vlvY
0eWPpiDGjN/e/wxs6PKWJV5vT7LuTsD3th+jNuiVzaUOqPtpso6UlSQpibSp
fQSC2zsY4H2XNdzxFDbAnC/gKQ401Ze/2fqrJzPGxTjk5phdySmNMvUHSeJI
+HUosfUW41++pZ1bmNyESdhmn8uLEANZOfQxAlL40V5oWk8MhV3b2RO8wlfn
Hff++HD3lUTAmlZonI0jCErw0pyChgpm7wBnBGHiwycCfUmJ4FhxNlJdHk0A
8EcEEOxAP34WS4tomd9P9C5Rgz/o2Q1SQAH2Fo4L+dYg/Fs1Mg8IjCzzmUwv
5IngmhqtLFnIuFPFVKvVRgvOxTUvoD47N2xiib9ra8jimGTBX9bdZZ1RhbKF
Dhh4ggGOEQxPiiRqkwoUrucyyii9Zr3wgOEdkumnsnmtWTW6LEU+5uITkWmi
DuydcsVRa/7qJTSnj7yJqXSSzhc3rK6td9qd4MpAZTYUE0pZFcZs8OrVRgpP
AuRrDOeerV5yTd2SqZiKJ5kSPzHwna6rkuW2WXkZCyitE8+BmcLG7a6tRjFW
EK1TFnDOIrwGYaB6VH2ysIcBIZCQ8WmKWcsnRHdsBmUT/D9kHGC/bom4QOSL
kKCNbKLU7WhgAiD6QcCIn7aIO5V5OJ4v7byAg8lFUXuNRsUSjBhBAI9NXrvS
D0Ppecb1TdmmDSofWlQtcVn2i8RGavmcszylkjiyxVbA4uLtKw8P0GZo+sVa
GoaHKT/RXG2H5GW2j90bUsN8uoEnX2sRjk8T4mVMPpjkXrja984XkjlEWBj/
tpWMXRLY+AjG0anvzQ0SVN3AvzX3o5n9U7tQek9ed4GfSn+3kxn8xNV/4pyz
5dTjETzbYdtmy/kdyBWSi2evyJDQe2BtXWOvltW3vMa5ovdhZhQJVFbVnEzc
/RdMatw7SZu06e/ajBlVBuUa7H6LIzQwgrfWPQHTCZddhRDKFe4da5HKaoi6
ohfQkWWN4GsJNEb2rL9fbNl5yQsK8r8zfVJvh42DtKoFGEBFyDV8f/MlRYha
+mr/oCYTqRV27TovjhMf5llFrvNQywA6oLj5p7BJydGnH3EpweI2JgEKe2/5
oVBBmirXyxWn+m5gMpLrFaZ5s/VvEUqziF7qmE05m8lmmKZpKsnHgpRHGwhu
PhsDmI5G4vt0+jZvaDa673mxLFDMePyzWsb0hEdlNwnKGwJOuBcwVeLBe8rR
RM66s2L/wDGkElABB44iUB9ogNFEV3GL4+NXfnzDydpanCN0c5rvL7LsH42g
I3kebUoOp8sAQJe9F2kpKWk4lnQhPZ42gU2FnRCdXVlOtjEmjsjbxp5BnSA/
Cc0HC5jb4jPZjsEm1ZG6DYAsjvPfeE7GVLDuyVEptlV0WCtwL4oE1fyfY960
zKKQPygc2zWgkBTsCWC6nXygCKnLCP3uI7/WsfmtRqwOsJdko7TWB0oDe73I
d1UwrH8NiGwPFwG77KP8uPyUlDdryvpTnOklDCLwa0yQRti2cbsITza0COb6
6umPlHiRJV3XrIMXt6Prd+sQ10dAfZa2rfp5VonU1+vEWgH+3Cavu86GXCw8
PbGT83i1vDEzRn5oeuMiFPnpOuSXkUsQ8uHyiErvDzYuhVdtjr+AizvFwG+e
bVYzLHmgs9ZRBX/W0OmqUxVd9YTIB6g1ppzwOoMjKofhcDaumXgrCXsbVyo6
q6uOKfZXGqaWhlba+UC93FH/UuEu3kspc1jolcSPouV9qhuHF9D/BvMeMi2j
G901ZVuuk7xXPgb6DTeoDxqP6lbqEuMMhMc/TW8THm58U5C9UOCeMFsF++nA
/VFfDs5SV4OqH4ro/eKxQBHvxYWlW1V8V9U1eLHAYrt0m+FKHdQ7tLsaKtg+
0PzLVgLqeBdac9kMHLMc/UVYWWioHmGR3+dA9AEtV+DOTC/2/9x+mf8tdmWE
fhcdoffBRZG6c9EQ3kVRsVJ+dTX+vhCPj4DPEme6oolxvJI0HNeUFdp2xcS6
T+W7XVGrQczk1nwuFYViLCK+QmwJ8wURl5vT0SjmXCHITwTcAr7LiZRMkVp1
UgcSAMBoe3pdxw6RtzE5CnO2MYMtyGQLutSPZe8sm2vscRoae12UpJoJvlr1
IyQ4jOFclYptL8gTgCG+l3L28Vd6qYSKOJSsctrd8lDxXPi9XWuEM2dsHKAh
XYVR2s8WQG8r1eGbjZYKh8hPD8Ad2af3U8K5X/mRWT2OaoRBIzbebQMmj6iN
EoHO+SZ5trg+o4e5u90pv7A943db/jpXeSgjLUW7u6cLivC2DSrO4yZPFIIO
iJY2YP8HdtDMAyOnNqMCajmoTFD8IxFbMBGGu+3xQxhFCkzuI2QpwJYj9M6B
AKllpmYrwz2b3rmFyEn6Sxwm6ywPUb+L6yckwAtf5ObMPMN1qlVPhy3jqq2y
TaMuaPhWP80evZifdWWSlsnpDqHJwV67u2wXMuJYnZ+PsfvLe3evPUAltKWk
+pQQgWL4jXDK1X/0V3lQWgIrp++OIQntYau+2kSJ7U3Tk6X0jnQfFGLXmWbR
+erDSMvzlUDNcpRVuM+JJj5IQdl0sVlxh+1lSsw5Jru31EXdrzg7LcMbZgt+
a+lN/ahckWK1UITQ1nUwwQt3W31vN88CPk0hLY4b+QLcB2Owk6wCNleIPNZK
s/nja6ujlgLbwoT+4LVec7qgF7KuBTCIBsJwX1w7f2GTeLquiiH7nzJU0vGW
Bh5NYpf+2mM9uY12D5PgbaCphLqgfcUtZ6cf+nNJbw84BGIhGOAtgIk9nxuS
/jHOiCDm3M1fTCDuFFDju6nyX4/+aCMOx0iG5GvbrBSNFrm3P6G+zODHiCp4
PpyuFrzh0tJHdBhDfPa2WypHu2A7GQxR2qh1WIam5Y5GZM3GEyKGgrURlNo1
DqWeNaYk8rlg/V2d+0COVc/kH9u/CnrsUicZwwu58CxpjHFN03xWYp5ZrkyY
6OJrCxDu/xTldqzQiYAIx+1tdiVdlM0axkxRGbLTvbnZM3CFQgXnGMeczQoc
6+tg50N0TwN0alb1HkM3MuUWvJgedQNNCbv+uCLUsY8JxEDD7Zh5VgN1Y961
O6n+7QH/IYjNbYNXTlDsrSkq75u6hsQGgvVcUsVoiwkxxvO8DPW/efX6JrUL
7/ejm24voyfAzQ2Hng8aGMEQp683xbviKBu1v8phL0zaF6L5PyDkHVEHOFI0
GiHLxcxINrLD6CnVS4eIfDh/3+ylnlWfV2lZ4Hkcc2TOBuqkk2XmOu4owm1u
PPbxcxmmCp2icZGHwc6++7BVtm9As44mMek5UY8RN1URF9MH3WbsQ1v3tO13
JGXa3lP4hnjdGGfp0wPe0EYevpxIRdfJenv/hR8gqte3m86sEB65pE1l2A41
o70dN9e4PEVELc/IqzVgSKgJpJyWt2mgJ7P7TaB2B4Y02iQeY0A1WWzC3oCT
PGrumpIVlah/fOWBCljotw6RmEbTcY/zMgxH5OFGHpY4ypR1WmzIH641yxa7
JFxNveJogrIaN30vjTBtHncYgT5v5St1Av5jFLnVoHlahnHp0fh9VqvhLqwA
lvMgFj62Oiemb4AROo6eZ8alXuWZNiqe7Xh3oVC2/2EWWE78z7hy/vPn9JDJ
H5oDDOa4bpqIu8dWPpoY2471wFj1Hkk2rb5s7yrsDk9Og8Mc4TtXRa5zGcrZ
Fxz35xby9HW6HcByt0ZJmsserknTNBIv9XBmv4uqpw4Chu0sfioIMNrfsCI/
KDi7LYCJa/T8DiGPDc6kLtt7MhvNKqN7/2j4eKG7diy65k4JOKRNn8hjJpxg
kZ6VJFT6zyC4hAcP2C7tBX3oqaoLCZhpqHFUvkxLY0DaqdykWsUl/PKCO5JA
dYBteFCLcd9m4JBPVC1jOS50bVUA4EXH3GYBDlIegUk4sN4duC1GrwVL1Fil
XxDle0DeVSbZyzjXVoa/zjSDbgTcvO6YfgxNudXUYtiuFdyBLS5pqyFodRdL
xYzdOFVacXFVxYOzRlk2EDVmq+Wjv1TO+X4LwP8qj0qZE3cARrtu+EjmFQsv
wyoyhcuKHxqiKL/1PO/fBzzN3xJ+MeAzEYlvj9Fql87OieZZNIDKqya2q2zx
1Vtmy8TnTs8E3z3cL3v8G0yEnkoxS/kpSJbTLKkeZKU+rmv3aXBi0DCArdpn
Qn7d0tGZGJUDY+Swcg97J8nf5OXFH6vjFL0X7SSQZG9/mRIQRkHIrTMsdKL7
UfiVpgoJ6qPCcwg8/UiWr3vUHGh82nrdnZM/tXNuCPyGX/BxpHVbAFHnjeLF
Q5bicWiEwJTGHai5kv8Tp/aWshK/mb/o9EAFR+W3tuS0Gno9nqB+qGHgQpkx
AUffDaaAAAqFwH7w+B09xwyasMVh8pF3sV8Skj/FhAGGDZkN+wtUtgN5cZil
Q5kZT8De1tqvfu9dKzbNTg7WkuUQvFEtUl1Oq8TdtpEZRd5g7NjoWxMkzDkU
tevk1YCQxV34AJNXqqstrgMV4wIdVtjJc3khV0mxRxd2GrMkwKTG3exqsuzw
BcQwwvqXJcgnI6HNmOC3z6g2VBla8rRSVkoqd6e/hrQ1ADGJGygODDi5j26R
cwFjnYiQr2LwB3+e8IDk8vsPU0H1N0oB6ByYxy8Zz0rAC7ZusewE5iLKFmlv
8UUwgu4J/pwFwDBTkQJOiSww2cHZznaLqHyDoIqZP73jh/zU41goVBdNVV9e
jks/vnB9YbKEpSPjkOmWSEIqCngBQbdFN/v003VqhBytj92EJzccaLWCvx1S
5BQWwDlJEgJm8trBrtFhCSz+mV+6lJMllWI/FIngkX9bA9YdJCfb6CQQKuj5
QuajGjlIJBcmMye96B1kmD/Z9Vtqx9+0dIv0WDRUBfXmpmjPoDkmLekaogOz
ILTU402OnrTWeC4EX/1et8kMSSFE4YmKN9DrN579uFfPqPKaYEIbGe6JVn5p
9j1Alof/OCrT7YOxshLl16ZCCk5TRccBavPvhEQLfaiXKbCk469W2JQBMEZW
8W57bbHbaPN4guCISXOwMJNY60036sPnVpNS+M5kaJPZlgdB44vsZzgrkXm1
MR5IY2XEeuhl0LOJzN/vilrTO7TE5PONa4W3yuxxVcVvvNAXkQZm5xnFL/Bx
aQzHJcLAVX85tx5hGNm3Oyu2O675AJgL7tnATI9UiT2hzvHHbOAEb55Pyfbb
ZzBcrY5KchkId/CMhWxXeT5bx/FFSDi/FUKSdYU00QRxyeP7eMFFcXrumvLg
wYmH0PlnuuHYeXz/J6ZqFg2rhslibrWK0WvtvAKgXx+X/l06HamZLqOktXjI
uVgCK2zg2AI7uyyGSb3BLQz5MfZHW683XubQzvtuK7dzExtML3hQjxyigxM/
JcutFfSBLBPXisgCUiAx8qA+1SJIs0oTYzUAMIsBrEYtyEuJ2NLJnnDXvoFZ
caIwRNdiKoDfjIGMLqu0MZ17Na3cI0ZahvQBAjjuto6hOIJS99sVm7cEuZaj
rw6/mKPPLZcnqC8RuZILnrb9shWAi5dGX20X52afSdfB/JCPfNi9M7fgOy7v
Iln+fSam/uuzfz+EdIpf2EL153fT2IfNS0yhfPVKaImFsnGSzXFaEHLmJdFF
VKQmlloKLQkg+enQJR++13so845u3IvLNdV+qHSuOQAJL3G2+mgBWF2RMCtA
WSqyxSQOJT1/2ENTZKZzPfJSKDw16Ou9LIerzoxSD8Ja1w5lxQw7wGbc0OV7
uxOON4L1U20VKYkRkXKx8Tv4CHO3ppsTiKG29ORx8y15n6TrW8chKXYFhq8K
JBd4WzXu/v8pIvZMbmrjPym0dk6Ua5x48p2rs2IMqvrCN8YdgGeC2Z8P6GQB
dD1JJmuoN+Dfwnor78boYm2mIFVnMiIgRHnA0nYfdYJ8aUpfC4oWfklmRpCK
jFWD3HzZ4xhgsvzxJ81u6iwMvrr5HgR0UdzDLlwZ7gb/9/ElGbeQsas1T7ZA
VkJiRWAyZfRCPCn7h23SK5MDlwO2ezl3eII1rXbzgqZPCiVw9fPRjI2glluD
TOjMuO8FyHtShSm90yXAJLkSynT7vKuJmahG81JWX6VSZQQUH2y0G/JLFq1W
5PtLit99qVlG4vi2YD3o4AOFcHoPe0GEUE/SDAcraeZmgtBu35dr+xuXwOpw
wykVQ8U6c981F8h5pX0b5oEOo3IuVlZuccXcfh3tnN1Z54lv6RG/tdAUvYs3
zlJeo2aRjn8E2U0RVmRvDoFycY8vZdatratrPjXt/VCikI1UilX/K9DAWfEL
RapRcwaX8j1I2Aq0OKFTFA4EpQ5rmMQhK3s/F+FnbDaM9hV7422i7MYVWIAs
45O+oA0e3W004GRH1AJ3mdnKuRHdF092mku3GXScb+ej1eh+xg3s40f2bHME
d4VYtsES7DSh1FVOX79rxsljsmBQKd+qt237wD27w799ZjoYoGGP1SrVHyRA
IjFzOeYPj2qjvj5PRSFm6NnBHWsxs/YBhoGNxek2ymsKvonNslV/+upd9A+/
4uRucqC6zy7xlyDgYNEjZ7jaUXgxrwitq6Zf4C8L7oVyCIyBi5Wh7fvQfsno
Lz6nDJdAK38aWCmae7rZewAmu1/T75Kwe4tvyxZAXfB6uDXP0wBCS924IHBk
NRcqFWhyZaPUJIwRJDkv1WtPISzod1g73r4aR9/Rv4/krzW4zs7Ie+7g/P+K
LmMgf1F2GzZozj7hZhj55KUUVz3bUglrnuQnKgUd7fGZSjPUOUmqFHiXFpUh
qcYIyCFaFW+Xv3gme/B41IQsVmng+SRSRUqVebqogE40/4FCKpYI7670svWH
MX6Sc6Ch7AnBtNzFyAaMOXtqLRi/RZl1cHFatgD0SD/9YJQvVC1D1iNT6wDv
uGOJmidl/U50Ra2lCnt92XoCC5KURGS3uaSYlM9BbiX0QPR13kpCzqglbM3f
2VoU/coVgtkfFiluy2HgKcZYxrW0Jy/XIYQ9xjDUJtV15YAB8MW+U8bLJQb+
9wt4cvTCojyoAUQPqgKXT3yXYY+i/EXVtQ+5dsR0Tb9m+CW9hbtS0BPFjX81
l2gewkvDBGsRKuSeokGHyxad5c/0SaB7jht33TQCLFsyHBXueE7Z2P1+6d1o
ewGc+aPGtDnjDnAUl7qcTldA/f+y7zuo80Bxf/5j/lWJ1oOjigD1bbtUxODl
owr/EHfbAStWmUBezB4jQtJXQpwzsQxMLzDrw5yvN1ozSL0HBYlIcFdcrfBj
hZYLz++7JYoMGosIN59mnv8rJ5vNpUWwT3+ZeU4qvaLJIb9/kdQSXnz9LLUj
GUERIkg3EozwxzTQM20weSTzHAXD2psoNOv1N/9FPyyIVC/qL0nChH6389u0
paoPmjaumzEsj7YcUYGuvtdZCLdxBFeOIslM0Y4vaD0UVOdudHv3P1UmSle9
O1FMP6eGWIaqqPSPbrNBc2lOigXzLf00n5J1OFWANFb777D8qTdvCUtuoamB
UhtEtX7hlVX6HIyXE4NRX7+bw056d6FG2qXgJZ2i/gARifUqHcbQK5cZ7xGg
kW4CrmSwT2n8C+zB5f/PIknm7qPeoSI2ywXrH9tpdzef6f+tMWMOBnD1eCUj
99M61wR8NGAoad4uQwTvIbfEWsvFo/fRAn6TrjMU1vFj6CQJosZjsrJ0PcTA
+97Fpst+QVUaq+NIDmLpRPX1LwmRiEfJyj0dQAhMNVPmBavYm0JJZj+cebC7
lSw96rFdaoeozzsKmhfy0iLrSCYVD6pZGSIX9IJG6erCxBuo+LPIra78Zqmm
Rsk9tT/mgGW3fuipXOTLpr31NK7tE1tFp+8FkiJZE0KtN0IO86aP/yXCaVqj
FWWu5h3NuPNllZ4MeNtG/tywUD/kJsAYFHRpRPOaYDQ/5Pe0RCTaWTr+DZYW
Q4gs55qRNipGaMljEW/QTlh1Ahb1psXVKPLzHUCPLnE27RMavd2QnwlDrFNK
NPsPxbwac7offgLZRCMGmxdyI8IJHgRlaw7vUtamZ26QsVyqyvT0+AU/SB1n
YqvkgACDfejBgNODFhTrVXpSYLZTbdqQRVpXH61s9P3N/Bj+JIHKVCfo/C/Z
JBXZgHkgNBSt9Xzj0hYNBc7NDm//dzA+VlEEWdNrir/sOBKJ15MmCvj3PBKe
ahgM0eWyli34MAU6gfuAf/l9K5CmO+CrdDp1L5Hy+jR53INBi4UVKxejPSTU
jB8knQ590/ODyOGiv4K9z8ARctPjKiCbrJwoorxW5KfmpgJGE23hvNUVbBHz
vh8+doNA2vGBODFJj4iaZyLgWgjjcxSiu5QKDzK0QNwbFjq77Xps6aqb+p6I
p7ZrpO9VN66djPLQX57HIvVJ29L7hw74BPt2NA19TR4RXidUO98f2+bZmhNT
5aXvLo6v5VsVYDEJqcBYSPVk5adAR6SuqmGwTc6ECqha1C2QItDWSL33pGKO
cXDNjClZaM1c2YGP1rbKPdrFdKVd/Bw4esEmrMbFA/iffU87vS2fa+F7MjKt
x2SN+8WEQ8w41Cm0+v9d7qDo3+ZQXxlOqHS5cESRofpepGUKLu4THLfgNG7/
Bzv5I5qpKuC8FWCvnCF6Yshxd5ninQ26vhlVooabw9KrTCygArEvHL3d1ljs
ZekbvF5xcEku9i9M4qa8Qcdh5xoQIeIAds/Oe2ABo0VnLmfFc9K7ES/nAzBt
dNfUKLPS82Lh9iD9iD/LoFE+75RXf43EEY73bI5591ZnpkunuGS+8xDZmg9w
r+/nw3FYOShLgwWUiZPbPffRWhF1GRYBiOo5zf/oUPpIKMW/7XpHnyWxGoqp
RIksbc5CujTjB+BsdZyGehYX0qL9FN5dME8liNcZRZ743M7Uqg+zyWpGOV95
atEYRaFBu17kzzdFQCm59jszWpInrLzZjXu8TzRhaY2cywLbN/vXhvZbX8yg
LPY6kE/jyeWQB0Fb883CfllVXfUOiy0kbLPbGNujvUaXWDo1yXJsd65NS6EG
+TEdEbKVmEP1yNmN8IFXT/DvrCxD1HrREfgfFfdRGGrvAh7XSzDVrCHHugRS
zKhNV+wnGNG2Fy3G7FYMPnwuHlIc4kn2Eb87ksDI0rgiSlM4taXgIvmzI5x8
crlr4ZR8A539gyg/nG1RWqBeBMXExr7tiQti9ODn5E6r2UWZzKjliZdUjA1z
hH5GX76WqlnsnQUUMZXHThPvjWjqKtwGhjfA9G2XuD+cQrEfjzOQauC89E1W
7UKbGXWohL32khD95oBMNU1KjZAP6qT23GESriP5MxK47Swq7VM5Vn//n0nX
PEzOHriLyepiRzA0FGzvHmVVHcaGUt5/H+b4eohgjgBbuMZnDLY19i4W2Alr
cdeAuN4RFTYjErp+7pP10/d8/M8SR0Yapu/i3UyMVpt3ggphr9gLq32ILriZ
8/pcnAgmx6TpCJAP+BbAVru2K2aONBiOAwa4SEMttoe7K77/aGzcNC3LhsBw
HQx3hBYsXdF9NupUZP7Lg994PQlmQyEvSYoQAWR+eMQaOPFAfEpMTMfOIzNG
ZkHK8KIYhyK767hcVIpSvxKEa2gE3PlqChJ9AwwBDqOLe1UOA051xobFHz5r
01WOgcg5/DxAAOhpTX/Ksvow4BG9UWB4Q1e9QpuZCUXKdkQ21pygWVeLV1cw
kyZJ0iWXZ1WB7LjcPf/sSW54dFqLm1GUoHZTVaX3bnoBzhro5AfBiJXtZLuX
i0Uh0VEAnLXrco9unFUbPZI2nRMABtazQSlYDwAUYYEQ8PnUPlHb6KSz9l4Z
+viDt9a+BYMXfxGYPvCnmcUCl9+Jikxbtf84KJ6JCZBexFIVmz7xl0Mnafmj
iPBPZj2RkigswgvUXl9iauZjlDPDyDM4Dsqve/eddYpbf5mw+rnrvPUscK3w
gIBsj2cZqcyfNN7SPUFHpMbg//N6fvvH89vuzo9RFCwxeEANTqpFZ3I5WJvJ
hafzbgiQ7wMRDotu37Kf4uL0JMKALtci8PFuKmOe0VOsofCou6Rrj2Nvre0e
vqtTKbur5e2t28jmNjqcRDqgPLdD2hmZJPrdGCa0Dqo9i7ttsg8rZoQpDjWX
PkS4pZsl/OevFG6PZa3nQZlzlhB9fS65dF/aUw2tjeutkgNWqAMPyoQ2pGoo
Pyp502GnTXovVLwNrXlWrsLEEkzB6KE+DOPyAjwO9cDrKhB7wxoAE1rhhyPA
vhXJ5hBAmbcUivglwyUUWepGNEbYS3DN2xzckQ5YT8Z9+22F4I6C5b/f59NA
yLo0zyQ9RVhe4RwDB3suZqgUvk0t2tfiyv9ClJhtTr48pcP+XisoiZe6VtSB
qnqKAgm91wIoKArApU7HXm26JRwsTui/L9/EP/uC3FXK2rOhVmko0dzPbVpR
r0eFvlaJwV0I+G8J8iH5ZIhrFO8c2VRNID5YtZcz3TeVdWCDlnFnO6GtUeeI
9SJ04BGFK2aqrAWmYf/EYsakb30PHV4BioaX/maJLGihsosfY5nIS1AXAvNz
a+reJ3XX8w4yZIPXJTKf0R6i2CoOAyfFiFPeXAESbXpdf/FjRREtN2ukwka0
pQo+7byoChxhK/thJRhkXYxafc/uf8BEqaId6lPQy18KUww1SVbvuXcMX/2E
EgVWZOKqhble5pYQj2mLtYQjc8G+xM70/cwsH+ro/gwze1hGcMUlzJK4pDqa
erMOy2uqb5xRyKuif3qXQDia9FjPreBfMYVSddzNvEl0To13P3QqW6LnI+Jg
g3+39Mft3AlvUAigXCbQuCVX5K8zgU3x2Et6mKoeCEcsK+eqtYB8ouYI7P3s
5GecCthHaVfd7oL6w8ogwkOMpbc8QsLKvbYlsk/ttAeVg4zBAVUF2FTPhLDt
ab0eITdWDMVGPPiqfKBwIelFnbVHu9wGaD4Ai8PSOxUKvSG8sYszdXq2VyB6
b19O10NaZJyXhp1ZOZ93zno4geY6CjF2B4IR2rmHQBnh/+h69fJA6Ub3vrv6
fx1fRtXA0uVAwUL7iRMc0ouuT0s4HDEob2D51SpZbZTY8+GwAiqqHpSRCBmx
7EmV+OblPuu38VlwGm2qBJpPhtku7oeM8QwaP4t0uL8SeIA97KQMnQZRMT3q
c77/nJyRDYHth1CBku8oTYt/EFZ1YB+ZOHx2sjmtquL7WqSEs29LfhYIbpbZ
QOkgpUrO9Dt+2IxcSbU5uRhyiuy3VZKg22PFnmZ7r5IkwwbXFuaehFZLP+Z8
OIlYwhECcExqA8p9DEAKxPFlNwQ1Yshvdhu+NM7O/HNeRPtzD9LmfeJs0zmS
FgR9+TJ/aICczaQFHi1f43/q/fcmOMIVx2cK47AAQF11OCldEIa2C9HtQvB0
xSJvmbzjV13NXN3lmXb1dC/7cwi5uhTWcr+rJXfGxtCR8ArwdgQiDpjqMk3Q
g3kAvT2CbtWXps4lcl1oLeRWBL0rJeIJ5wrv0eNDn/rwKOUA3ohvPRhdwMrE
zRrrW3UzVX94kJBHIwLrNRux+yRwNOKM1ju8YVMLVnonV2eMnzIESrD3UXiB
bcAo5f2cyaBeP+19LorlIGK36NH2Hm28NX200JCzDPJs79sPG1GBsOjgINN7
fba+0enE+xFt7MBv+gcN36ni1ZWPmgD7Rvva27lCNIw0aYl5W+r2kBL+fo2d
7nIoZ8yppedcwTQUraLx8pnzbvKpvof/W+NyOvuH5EafuX6P1Cy9G1gExFsv
yc9AQH6i2dEZuKChM1+bHa+1+7oSc+UiILjhaySOvW1dpUenNFPCaixLEe09
X82ngz7xm32dN/2YqRJ4yknNfswUNQKlyP0VFoFRbQXUm2qt+pOUC81lLvqB
PsKwtKEmyLY+Rvqvc/b4Hk6xceeVukOA9hIsTmlziKmIgLRnhRBaIOMODdcd
vLLKOGHXAtnq3yi64On5Ev35BW9tLZCBciesboLbJWVmVh1mhlgnD2fmSnPz
VfRpLitJsz47CbC83HRxK0dnyUhug0P7XV647z83qNAeujTSHQvbkLjDhSfZ
9VqPDQcoXArbKpE86Z4k/lEWubTfQt4q/gF/M80UpWMJ9OZT+UJ7AOg7FxtI
Sa6BKJ8WotHLzFOFRviEUBOUoN60KPZKYjA9rArd/aVe28+MGa5bdooSwJ6b
rjo82GQcxJdXL3wuQ4fN36qDjCGLMKDZ4Ha1k6Q96zpWK9Gtoc+0nrH4hSjz
mHcqAMAUzctqTdZAdk31/QcTg99XGZUxVg7gi5nyZT8vHOst7mU7Fjl7Rkdq
FHW/G9cIrFjxOB8LJx41aUeWE+5XRtESHAgOYQu8O8u2U8KbdWaxDhUkXugW
J+FcPNpM9jeLl6JnBVSQJw315ugFRRpkeYPzCSEewa/Q5KX6QCBKxtxbzkZh
u/OHn3Jxr8vxzsuBpOEBo6N5Jc9S+fE2HfPKK+yz+2ZZJtRExpFjIzlkeRLy
SyHTGTA/jpSE5ks3iuGx5dNrYW0ifYDF4a7uIB1uZQkghGKFw9vOFcNdWe7l
nLuXaQAA4AWe3JDz0yi2zt2Il97TPPW2Y50vwFPNC7Jwxwjtg7cRXIUGDCpj
JE/0PM058dBsi4wVEvg+eFKTo4ye/YGQ2QgMZmRTJ6r06QMIWDXhsHr4EFZZ
HcSBhFj1cBsOIArnw4pVDJWDo6jZ0JuidalxMZR7i/pJdeyIES2VUO8e92LS
JgZyIxtP0W4kaZqYRfWoeBplwgRY1IKmuhOF0bQXfffKPDw6i7rJzCsyU2S9
f5y1tE6ToaUT6R1jabSm7PbEQqZGKetXNeeQ5vfN6rQ1DSu5SRnQzUppqEpG
vH9WEI3xGUxxc+c6HgAEn4mmUXwl1ehjVcBQQJQ5Tl3bUTinZ4sE+v+5Vtzm
1Kwsike/o0oYpOIfnrzOT/FdpedKV6ObFpx+jV7IQZAsbRvcrES+cn9EOHoa
vjfqPtA+t/IVN2I7B9ED/RDBZFHTOSsyzs1UQ391m8QCRPucXMUEmNXWbnwy
ei53yw+vpncUjmrfGEq2czpNcBz3zA2205vqPg9WCBytH6I7RH7m4wgR9rYs
6w/bQbUefAwVfw3Hcm3chkkW5PFZ8QnVq1Dbmd3SMmNEOZThkv2Q25ZpqAOS
OUiAoA+pD6WtSQT+vDkX0P/SuEQYV4XHrCgA7sYhU0jW1py5sh4/A8LWKhSh
9tGF4JJnrdmbK9WSsDOrEvOIJuMsdni/iEYPfK1kS8CsfS6P1tjCjM3eiZVD
Zin4Swf7IH/wu2GGl3c/xiivR88Y0i/I0Y1x89WqcmffIkIS5AhplcjQyVF3
INw2NZivAgxT03BgLlcO38U0qS5rRFSDchwxrQupKdEvd5Ca+DqYSUeCOdij
9cVNAtkGsmZJc/WgdyX7BWse5A7QPNpWGT8yMPXtE2g2NjRNAg4GTx4n0bbX
jDgnvDd4oGx0xFR0Igx+51ubEZAfbJzEiRCvJQPa7/h/NdPqWM2vp0MXg7Lx
bUmfRkHSyv8ko+vmGzRMhD1L2eLceE/Y4UoReNDHomhXjxKJsIq2j96+P0Au
dr9KGKhI37EMS3eXfmPD2oS4QEqXwmB3d2dj+RmF3CWFfjONk0ATFkkURyxx
L3utoEAtCaye19+1Mb0eWuy35gu7JWyBiXG9Erh6DCGTSBrotDimN3vQRpHS
nPzKEYHvs4M5NXjJKGWzz8dEFZWbid0VupsnyNEv5GxJRZUAmnejl8Xl3sT4
pmJC9cOcX0RFbCJ90d/ZGbw9t3Y3jw8AGsBdEKfOjqLpc96U4er2pih5DEeJ
zSAJ4tjvTio7Ab0d2zQSu2QKEiqsgKIbNNK7NADuIOZSt6i0XM5ch5HJWfxU
UesSgvXKX2mdJ8vz9GWaWa+pc+VwNZwdHTW8uV/2OC+lanT7vMnZQuxGwhjF
/z3a0+/Y0TWwRhJD0S8zKGI8yxZiU1fvCoVvsRG2d9cRAe1jXt2gsbFX6Sav
Dv63NKC37IEmEPMxBQbIGWe2IWDCTuQnAcKFsWdodCUw85ByUg3KfDIHOlxF
gtbQvLkjkN4csX3ePNGwpjRu6zi8gQGbsUZBZTX4686sFsU+6i70C3gY2huh
cCyt26+0ocPDUMVxKd3h6kt8bGFYKNgkaC3yALjXzwq7pMfWevFVYs+aCeNy
it91jK3lmdXwgbrTSDqWiSvuaseyk22L+KReFEWLEqGi7ybauSWPp/Ufb/fw
MJTCUd54SJqFHN/YY7rFrIqIxHfltldvLh/bDeMxpvBHn7We8U0i2Dnc1jc5
s1e/eQf8a5/f2abr9xPzHAkCF+9QqOuEuvhGbGdpgV1HGPk5D4V6kPoutPgo
47cEDmfo+ywxJZVtk78dz2LFqDG2QMtV/hbyqnfpjmmfCGj4pGiKZqHajoVK
YidonwunZVrt0x8GZHFI5f01BmohzxjdXgNPUGjEG854Z6LzMEjNkB1VUyh4
M/zFC0/EE2BIZVj/vFPrhJ6Ttrt7qIhChX/xhetwFzIjyWxRFE2nRboIk0b9
mb4gEhH/+7C2Ad2HXkxOrRUkPs69k1nWy1qm9Xy1zSDGNqZP8I0JBcBckNa3
9r+xcJIymtuVGOd3TnTXnUdYDtsGZbUXntdMSvipFhd0KjnhbZGxqTXZiPvX
a53zrtFa8YxoLzm/sEypFqVn9lypWLbxzcWtVgwks4Y4QVYHlLnZ8E7G4OE3
RbFGVuzLBJAZp1U8h1q8AGVEhQ54vY5HJy/1ue4DhUq7KWaL7alKqP62Gx5p
H6gF1gmul3VY3JMPsMqkiCuyu1aP3/lmqShLwlMI2wESQG7wGQHakGoj8uR6
BL551jf2sfWsFey8zIh1nMPgzNDyUZg7MKEAv6NxGa+SzFJmEYWm6v1Bmzb9
8pS688jW2MvEX+t/4yBWnzOamKIPly2nY2fI2CqyeyTVGA3iBxYct/NdBCQ1
jCPTweaqyxRpx2yyxaRAxJEzoqo5noJ5rPww1Ux+PRUJi6We9tNkYf/o2Br8
Q0ua77rShUBp4Nce5bs4/7XY7NfQcEyN2WnV+Z0Sebo5tPPI3bf33DGVM4hK
x/KSJen0ykbIZL4FEWdL9sJ5pVDVzUCQvzAo630435J7CWjxThzxFcgbiBhb
0uZVqsf8996X9jj6z80UAsgy39RMaYoljR0KXsGkHAK2AcBDKyKNSO674Ogt
nMyqXn9jq/OBmgR/lu9K1ylOFccFBstp2K3TtvEXQBGYaTqOUDe5xawfz68r
dbXzaAkKyUBPzpgjTZmRoUq7G3XhlG1SsfjKR7b6FGJidbhTlRvYbDD5TNQ5
24PR+BCkhtUNHtQv3UXZEhwUf9pQBsTfVFE6x09tDIbjp3+gpgTZiwg7Aknh
8iqMysYXAlspDraO39Md43tgUWwiUOMf/xXbr79a8D0RTavyQHLRU6Goe/Gl
VJkOxSYoXfGqsxDaLEx3QLeOdM2kvhCROihruzBeLStSFijAVaz9gfDd7kDL
INHwsZAI/ou9ifj8Gs9UI61bqwv35kQ5iyFuO2xOZFCtpcixmgC/cFXVVMQs
dY/EsOHz35k7y5PYUvjIjcGfNCsDYo1aRoXSkc6AdXHoDPkbfOGu8MguXkkr
X+k19mQgOVw4TfRLpMbNateMMRUm7RmO4hnsBK71dZVD8w/jHpHlG+hJout+
bpVWY2l4AsmlAOJAppP2l8PUboJ55DYrGzA2/7CIjKlSjgdjm3NYyt7Vayyr
iN9S/3Re0eg2nhgK0xXwJ6tZlEcW55QCX/kqkUc3Pt75PDO0FK3G73YDmtTA
jSqAatsc5ljEmec9RQImT1cL9hTG75bxCU8nPqRi6ilrK9M2OMymZzjWCjMB
bXTWtItc/kjlosejcZt/TAj4/U0MguYi1Qxbtw4SpBI4AqdrfnvsbwuukB8z
yrKlnEaiAI5/Ap34V5Qd1D+M2E8waQvrlqehyEh4CxvyXCIO61vyHfwoT5ll
84QUWkfcSzJvE3VgtQlb+5UxgKZJRzxl2MVFxYJTqJAYguZxJT9NnkTocizm
S2XwZZSHXStK2qyECtS++0xLFUkUJO29zlFFd6DPq86ru86XDSPW6NK+9fOd
gVTAlUI8QETpWeUMvYjUgjeymsAL8F7h6fwarwZioLj9la+ICnXRZczpvolB
HHZ8Av7iH2K/9XPTx0NOi+uvk9//9JRe3AiXtmsof1QPceoD3qLGoKE6P4s5
BTBGsPw7XjcFrFMDs5Go5tr2BO3TUMvmMzjD+g3CxTJHYYGqVNt6r9Bt5nbY
rqq0yP62G88cBi0tkjcMbfEcbQmDLVt6NdC1FGMgIq7O1C702GP7ZCj0kXw2
kWfTH+akLE919MUx94l8lck83OM31rkPXEBdve8qoUcNC+Ay4bdY1V/W5V2b
7y26m8QYs7Jy/y0CeqqAF2ZwPDs3XSKA+F53QYIto0zrIeUiU2ttg59irihx
gGi9J32ywWTHC/+dr6qhDxjoJssEFe/KJr+o/hRDPuzMUumhAgQjCSlmXJzE
b5ZAnAuS2+4tTA0wR5ECby9vadDO6i0FUT4zsANtTHknPFQLgDSnM9iMHhWh
f46D72s8g/DcG3/dpHtxsXiN1rm7Q9IFLDYmn3LrKyPYPAciu1vwjwWkJrO5
lqK2dQnQOpOw8bq3/+X/PkdN2gSz+rm52wmM0x5u2yEY9wQVvEAAFXHk7XMM
oZ2y9IW/kVVnBqf7RPvKUt49HvrhYmLAjo2pT+FsPLnOWT26pHaRzOyitYkK
L36q/XMElJXJ07deLrz952b8ij5/4yQjozVPSgYy29tj9fUADfYVkkomtsNy
/nTogViS339Z1vF93qtJbBRzWpP4sS126s2rObX5Feq2A9u/8MKLvf/hH5g0
fF9+WHdeHPvmZEHOGSqYb9WTzBNu8ChVR+V6J6m35Ua4+nsUDSFodiCwgWpE
UU1rQlNNhKH05oDjaHHPHU1oR4EXEzM39bUUaZCFflSFR/PrAdykqlN3MPoV
4kCOnqX7sFa5wYAoNi82stKmcRg90YnWCcGomQLbAMllSRO5MHef2xQLtqY0
WTgQ6R4ISRD9YlzMQfHVQ5FSoZOofBJabxajWK1IioL2PwdwJNYv6x+FxoyK
7KyRKq5QRe7V9WP61SusITmyn5YW5e1UeZP660449k1/FSLA1CACdf+tTwZl
KCwLbpOX/l3AX9S8pRpGFnfXL3T7Au2jc1k5b3dvsQpo0sKTVvC6WiynqMZj
JtzsPvn5q4j/xd60OSsZ7AwE0aSWfDccisLHAd5XcKUM8BOTLUYUj5G5pv7G
MUWXto2qLSZINJM5nO2fZiVPTrwX8Vdv/hLJvMKHxV1XY5KfV1BJSVojzLcP
0W4fddEbgMASbm+GJWj1taEyUcwHXYuc29RKwWxHKubVcLSHMDLTR9RB7/JQ
XZC4qYjjaZcSws6Bp02iGHd0TMGomjqOTs1lxu7KsNsbpCDFW/KJhBXVFUzh
0KPOwSneUrcAaOHrv20+zHntkYN11aiUyQFp6WoKGF5Zxq4Her9l6IrQKJct
SrWFpGI2B/rgxHjgwnmzByhkRtvvCsW9LaGjhjU4NXcLuNGu5EFcqEoaUSdj
Cb0DYYGf8oxyqHg3IjrfURMc1hyqb8cOBExW6CeCRB4tZ6LaUyNU9vb080M4
BZdVUNEO14YguG5BcPdIJPWUFRd1fY+/UByNZa9FljZ/UgTUAIFm4mZt80iq
bTKUXMMWtNxNKpSND9SjNoVubgUK6gM46Lf3b77QOTn4vmwqFXCM7m+yMNXK
PwDYHUk0v2rvdE6LBZAHpxkCN6h5L1YzHeixFFMHBXwGKDzhrwZwRPXUGKr4
QctbsbDfnsWw0kdesDeDHJB8nWxshhDp0KrvzANPsZz8OhpPtEwEkDu5HuTO
fW5G3XGakGWO/wvKa/VdNAidHceiJ9ZRVgzE5R/D5nVZqm9Omz73SvgrArzx
eieFE3CAbOMhdhkkXhx3WaZGLejzaNDQrVNcFdlIAvkrVDyXIeQAG1CuvNx4
zA9ETdzevjYXy7nVR5VsCezFWbX2uY4Xnt/chDRrA1A53gfUQ8yc8Eg3MYbx
K1ipV0/ozIzPhMzzMlK8duO/3IYNmPWCLgX/mI6u4938pdiyvZdJrvaJnR2a
NfL71LQXMA2hUFlnWJ+bx1sGflvEP2YlCcNVP7SZrhERP9DcAfc/sf1D+pDr
GvnM6Es3GYwsbVTsnO1u8tosfKl932oRKpcCBOJgsf1UCxHVSsu7hpNom829
W8Q50YG6Oo8x2mqaDDf7A/UUiJ1q5YHktIKF51YiqvOunAj9o/ILu2k5s+BE
7c5gmBcnuoKQ247LblML0BPNiHUJwGE3DhyDu3BTBCiMIPzCZIu9vMo90xhq
vLPXrkAn1R/QtkMLLO8SPQ7pHHB49auwgwj6Qtf/uhsJJjcUIzJHc70KLQfw
wFGiEUp8mBLOzJqcs14SQJjzWUbnUS5yhiiyFsCytpKjmx2EYpq7m6vawRaL
dbbSAEY0LwvT9O1MhVMysWvnXWHv+sOMIMFRfN9wg41RClGQXjNFo9e9NCzX
eqoatSPR5BOUN+YKToh+Bs7B+sOnnERg/Fp46CkdZxYfpc1tCESPSsXSWZ5T
RLt6zC6YP1Alcdr0wz0ga8jduPXVGWeGQShD2e6Ebj8x/Dpp0Sp+VC83RH4G
w+KXxZ8FfJ+vANP8gcUpfva7+pdVkdywklApSMEAC7F6fl4KTkfwoPDKb6XA
K3Ylz13NIoCIYJ58dIWO5iVS4hhWv9rDhv3mT5ZYHrw9orMdM4X5urawGQP9
QzaKQzzoXbPX1RGTY2X0pptPrXZvtkeIKxjNXLJwFIer2hTtg/gyXsEdzqon
UXVgtuOLTDPR9Civ4NnmgRWPC7GZyg1NKSaI52MVYeZY0fxKmxBE3QWqe7d2
BxIyIVwVdpOIBb9fM79lUkGG0Iyg27+ykXh8DWaNBcyh3Httm6+UNASG2OzN
Dn6iaPTPFIKFdUuX6Hn0UUj7daeWiXq50MC6qwvWpG71S2IDoapqjmetMur1
mq8TASn9uMl/G2LnrigTyhBnvqQg4Fki7LsJbul+RNaFe9jqC9ngKS0qJVPY
gYuYuoGy1hYrtsAb33XsA2Ix2wOgi4Rkf7pwk1vY66nDehGxSkcnkQ+BG4ft
A9ikXqaXNeY9aFhUwPrk2lwhluSGysMDyrYkEYnesWPHq5jdlV8jk+K2cuFn
ZJmItQWdveicpI2B44KHEwKJfaTevE6TOblrutTgG1DKNiZid1M0C7QAcLvV
EFrwAIQveRK4ro4r4YEklAVtRQgIbaxucaxiieumR0cE5fgbjqJQXkGCG4T3
ozJSsOGdQthdbSpB7m/6cjAh9wg6oMkkGzK68HmmFsq8EZcGNTeZ69HW6ENW
qFr0Dl7coDPNS5lSIwc/49dFu0YZfDfw09bF3ulFSh8fOt0FFafjLqCSY79K
6JFT4CISg26ORor6wQY/tqtzNGoF+IeN+XZYT2RiIc2FG6VanKbtzIW3AJbm
v1OxiAO+ExFtfIewVxqpgcW1FAXFACyr4a74qzRm24MV/ztGa/OIiwpXHLL8
xLxRX28c+q8F3Az+K7lu1deJro9jCYfVQdF2QMBhztD+bV5UNe2I8VqxqtOu
jiiL3mWadhYuh4PB7KuxCYMUSo+2CTlfa2UvdVHayursUqXuRkc1ACOJpb0a
qTe3GGs3ZrydOZMEt7tLj36KD5duQYo7M8j6j6ZU1rIoXDVEokSlZlAIEOA8
bS5vSF5ElR98xiq6OexFYxHmnfTu31Ajgxv4nh2/zkTlXzgzcIoLplewn5SH
UdI9GUJFkIFQ8rHpxqQWHtk9i3cmy1D97tpUxQSFFqW+EtGslnjLSc5f0599
vSXnay/sRkmvpcCCe78zHcsKJBu4/Qhfs/D09/eQVi2pxB0G1Oew5VDYWVJz
pM01ias62Loby/3vn0FReP/a/jLh5aOVK+Bh7x20YpTxPdJDWvwYPcuRw/TH
3qlkaeSIl0E3HiF1a9P4xFRrf0RMjpdHrDcW6VrqqgrgVARM3Q75OEw/Wy73
+0botsBwfV9aaBtY8bDKtHLSfQieHj7F4aaKXfzbmQnHleLD/vgtvBKvnNmU
7C8qapJCy1Ox8JfeoGPoqqb+GjksfVuNiDH0XDWSPa6ep82ltTVjLuiQtEMm
OCS8zgt5Lvxhg1WLI2C1guPtKvHItchkaQvyweHk0g0wADa4Y/EOiIZQ638z
93pXPpZn5JzlTaftdoz5gHcBBuYynQFjEiLKRCPG48NantzDnhtmk+PoelvT
xm2yXiEkfsGgIKGRJ8STX1KO65fZLbu2Lxs5TESbU1s+kQ+u2Mkhkb9o91ca
/HN5En2w5QBg87QlMZR4Vfa4dLkVJtIKSHOiLzyDZ22lxZIyuCWtMq/JH91G
WNv0NEz9NE90hL4le/xHOYkxcDVEouZFrahxmJN9+ZTNKGx7xPYC1K6GOVcy
k13vwBguKaPUw0WTyT64XepZd14o+XkTnzDOvK+sKHv1O54gPNAx9Yij6m5p
MjTSXP3eCsytamHTweYWZfH4vio+nsG5+2axzGtGL9wXiHSxWoX1EzSp2vvQ
j4NS677Pp+egQDAxsJavDkpWbEguafEtODeGpNHOiatEPT+dcgvZQBfYeyET
UZdRssurTqvNvjskPqtyMxJyCymd8UIvDtMz8feYPFYAWMReKtgg/4GnwLbW
dybYv436smPE+yVAYeHfVdP6U1ycKChk+GveMdS6SCvo+1OcyS95NxxA4gs3
dXPXh2sreawvFaODHJhX2J76QhCTyrySzNVE57TEGFK+XJzBA55DAjvq2VQm
yOYss0jZr1UJPvXBEWGS8Is9Jb3LfDdvgr5iU2MsvC4nb0tv5USccMFXpUvs
VNThVd+sFyaVAMpjZ6pWxSmdoxvPr7Oxy/zJ07MUY/3aYnl5g80xkTQhz6Fp
W5oZbBq15ugMzoRHkjf1xNgAa5OWt3ks0Zp0XDGQvRwMshqAbKJ+7GpYKSny
LWToWn7SEPAN10KusIDOAifd8KZVq0yquEEaTOIQxzk9AxY+fY4hJCwfYShf
uA1NQsIK+W1pVXe77jO0Ak/MVCZ7XGaXK9+vIqn4RidqocIS/3jr62NfN3lY
Id4LZ5CQMpr05caQYG9jr1uDWjRvUxwhYzEt3dC6jGzY7M4nKDRCO96r79rN
wzt9jKzP5SOqPwH+qfgIT0m+NbC8lfuLgiPGRgQ9+8YHd4Yf68TuMfsjS7lH
unjNcLBv1/rlmRH7XPeka1nSFerbUVqF7q9cw2xnYKtpq/wmTaqUHPrqb2QV
hFAFwPxy4HHZkGw7+6o8vcP7Js3F0gnxO+Gf8P4qsqB1xEUtW4XdJ+tant4K
v5l0otyv4ILN56WYjCE3AMOTgHDuYfdTAMqq2LzrIApvee5E/jUXGOigX8sx
w/UA5ICQXcV9jt14LcyrD7ArmOOi7Z4frH8OLqStaq7vyco9j9RNJG/ZoiUd
RDvXXob0VTQ7tU18wsT3nvDLkmcLLmkO/muRcSaBkI4Cr8GJ5QRTOJG/dcOO
YPECNaBPBFzGzF6ZmKGZh6sgdY8JUZ6swaUR34qglAK+ETyTZqhKLj3/2plA
91c2uF7OcljWr2LFKEJi3wY5msdqfZ9YO7GV+hbRw0Z7pTFV7xWvFKs0wlIi
YHw16SOFT6CBp+Egjf+UIPJOEetCecZxXUiu+u4iVaA1+6fnk4qDjhdFa00c
T3q7oMD1EQDPZjwJ4yiTj4Irl1HwXcKHk0hWSBZ17l7r/4dzZVywg3Uipe9A
m97BHpewE34V6O7Jqma1H00s/qRTxcCe00h/rKdDAneAEOzydllsBlsU/lb3
wiSleLy9mYycVIvFU50igCTPreRElewSz4UePcViOjiISL21Xtl8eyZfJRKp
1Gwge0/KiJaPQWuyyJMLi/vO/vA0+RmIMdT2xMNunn5O1A8hMGncgkwk8qmd
r39aI5ut9XQA73kK4iud3aSnoGmvkfmZcFMyK8XwnjdoniCYzYI+e8FEgWp+
KLWT658bpzBre+dAefT6l8oQcGO0kFh/qF4rMEFa9ayziWw1rhjHW5Lz1hg/
l4cTCe8LVPQwJhVEITiNBygZjj0Nj15HxPCrJZVqc3BCH/CVg10qmxGMqDZh
ZAL/ObhLWfhaznQaSsIfwKsqffsYSsVIqEqwiYrXkmsXjur52AU5n7yccMIN
EIehXbMJhaYOJwM2/Dw7S6jbEI0M08B4xYPk8BOB1s6LNn02tGQw+eeVY5Ux
543I2l94Oeym5ibxreYSxZAj1qeSu8JYiyn62yBozIyj90sbtQykLXhEQv5N
a0FRfFrcsDShb19chl03faBSXK8hNTNaVDxC/uEDW+zkJkmObSeILtMfGsX5
2kWnR/paXh40LMGgw2L4XsvUEhLMSlpt3ExgY7bftzBATkII3uBuxsRNUGgW
yOhppMBaLDdww7OZDBd4B+xw8SuDTj+z6X5tq8IpldST8yDP1aaHQQKbxzal
K2UQlOx8jCMq/mdIGnEsvAL48jn1ls1lGb9gd9CyaWfucknq8YuxjP0y6zJU
8V3TZ3Vm2LbnoI4gJVx4E9S2p6ln1aZ2B9s/ejjkBGVEwzy+m9ovu5IpPPNr
ZQbbV+BmbQt+yQwT3caCrrYgnrRo/r5YUBqiDzh1GemrIuj1I66v+rBQPJ5A
kZqc01j51+SkMJFGQ4HTBTDGkajajRQpwAwJhyPBmsasXnsLEqfaV6sw88q0
y8/W8pncSfBq2yMSBAImdYuPjRDrjdhMWpjeZHyWE2ozbVWDVIPGdfNDGqIR
65h1sa7xvahOKTNwjRSmuCwqv+cuTMHPx0+O9rD04tmThW8l4e/buSb/bmZy
v56RiEXRYwNV83eJxBgKT+4U/2roIJBQuL3xM6cMmnpJbdiNAskQi2E9Oxb+
esCNXH+PSwf2WKZvy3sUzXoE4lVSFRABjVlSwPam/RXWr8osSO308ILWMfOt
9bsqHSqamB19qH4LRwqfMvJP7xOMzMO7Y1pRV+P8whY+Vw1F07XA+eLk/9Kk
ue7bqAqCGyoE0GBUD+xb1b7urcTx3JA7CTCKgN1djl5mGmQW8oGNwWym975Y
DJDomMtWQL2uMFDe8xJ23ZT85KtFNCFz2SAglRLC8KzEkjYotn2e1R9pEf89
HCjRjYRZZGqt76yrvITvHYzN8bZ0bhaUxus/fV/a92cmYQYFAIBnr/8xtOMP
LMn9SnTmXay2aka3iObWXBMjVIQNpMdeq/qoVZ/dRhF0FleNbLRNTGp/+0BM
kCZp70D8TcK0y4O2OE0uE6W4x7h1gA9ZNSx5jVIp6fgJZrV6lDQLbdobbxNG
MZnnJ9pDO5pNUpIz+wg9kiz03dLgoMU64uqx023PmJO/FKeikt4QTYhyhgo/
U9mlrUAxbPewwM76i5DyzrcYYnTme5C7qfJ40hoJlpa0NAl9Ovjy3O7zGpro
2VYfCm6hd/q8Osq4Y8JwQe9GDfWni9GaD2ABx1l476fC/wgN7M6ehNcNSu7c
l/KsbzDVOHarauiASOVp5F/g3oRKtAnOvZdHAreSsMheFUtm1XkKdrkNS88N
ebzeLJMibrE+MRs4U838TVW7tlRb9BYuuny3Kv0/YB+u8dcLWP51Ixshrx0d
TrOt6duXFEr7JQqYBrf7DEbRmJjwfXFEEntQabP3ZlnykePhrqlhVNdyt4JU
iAvoo/NCx4bxiSuk/6JNov/rEzDgHLqe2KdqefAvoMEq7lIhPk6VckGch+eW
hGcOjBztieeNM3ZvsaC/n/mM+43Oiy+E3gL91jyaggkQPVQoMiqOJeF67EZJ
cDP2leygH7S+DOyY5xJyxh6pg4Gxq512iyQ3Ae11KZMFvtleAOeRQWtu4hAS
WFLZyHjAtnMFg8alJUD5hhCJt60sOfQcOUgRArgDurhvisJGs6OjbSo4ZO3g
ss+bWP7hwp4MFa5T4QC4fhDLnZozXt9r7R3f83YO7fhr98MOul/pLZ733cRK
YZoAWbU3g7pRDcQtWNLd22gdZjZ4oPD/+vQ/YHE233Ew1OuVU9EJ0lZOz8TX
D5BoJhgefCQOEx+IXjnGoWF4aEFqN/ErkbMphIMMPR8zn8T+K5QlA64acnZN
Q+FDeuMG6N1EZCzcQyLAnAwtcF8Qiilqgaavout1pJQ0cXQKgcuuWEfZe7a2
IJt7cDVnBqDfRx5a4BRkxlK176u1kdedM4fZQTDHQFELJv5uHxmvKRKVHf6K
yWe/Z5ztWjcTCZ1p4hOn4N0tWm52F9CgtK2DroiXifGhTVaXrWg24KovQCKH
oAicrT9Zfuf79jwdSnVOi9nXugi8j74m/XnVQaIW4mmNpAbN1Yh5/XS5SNCF
uZ/fpztKlmByr1pNaRvATIe9H8Jwo+wYFqKeezwFyTOvn2pri51M7roDYCd7
3Ya8K8QnKph8pacO3IK6xPqn7ibnRYXVaReTFbko/GGhS4lQ7p4TRimVjsrc
ttBpLnZ2cU1OwAQX9sMfceSzB2WMzW+f8zaaf19ViC65FY+Fs6IlbFSUJ1vi
2/1VQqkOHeHL7MAPlUIK8YsIFeq5Xb3QqxhiCCCjzuD+c60sMn9YJzQU9Mgl
NDiGsHkjVOTaVy63ms+fsyI9M+wkYzsK4bxFoXjKLIe0BD0eFHt0kY5gFbYV
XT+HspARhe52/r/mTSAuvPJs2lOlSRnGn+z7XbpNXQUxQYhGZe0rZshsbmL/
qVSFlS39lGK1ewJF8s9NGNkjIUpqcloV4HeamTDaDlflpOhDntoq1jWVvMGt
T+iwljjntCS3BLd7OpjLGLKuPTO9HW6h7E1JdAKwEkfY7pHWmowlXDjykC6E
arOuSSg+vgjM+LeALbmdbjcel09HXHhaHwGMtsloyEs6cLRxL1VHIAZ+TGuf
uqqYIzz+fVRacuBvUyVRi6/a1BfQDRLu0wvn/zndoUqRjVl8qrOno+wWWkeL
d49LMVkgsXCU1OGVvVELUvxOYYbpOI4HJTqNC37d3F2bdMTyw8cuhGLskeGn
qrWydReP39klU5QyE5Pykz/iV+gZY2rdfKDO/rxwVY0zDJdmXGgMwl6eqJa6
v5m37bX1B9rIqJcP1zgbr7vfAZfgp1kH9IynFgS5Q4QzoGE8RCXksRa07Pjh
6monvr63bPE+MH1/aEM6MF7Cl6iuVEkTlVtYExBHa0abQmCtZyg2l0s7+3sb
UTHCdwjlPn0bcqzvhDQaQHIHMcss2OrbAIA27PXEk9nexJBg5+e18ADud9PL
ksJsVa8PIVTuD2cKgjE+KNPOJHLZkUqp2RhGxAZEscosuObVXPGbNfKGcM0x
pQhE3LqVfh9qmV3fSKOxKke7IvW+FPx+0RdbJeeCYoMMW0JzsvIgQTKFUTbJ
1pfDKUzo3rRKqeipIi7whYh0S29/sV9+1caJEUhUsko53YxDA2ABzAWxcNpF
7t6julKssS3Q9mhHudKxRILVTM/ulneyfbSe2FC4vt1v5S2TLjS49rTTRxFI
Wth2nyq1GShd0LClNJ6o23R5zduZp06X5dJ91FGmuUP/yhG+w0s7xdyt8nyc
xmWaddFFxjwyhxhfkNYO5oLR2/cHRpnQXCiQAsVkRWLIeVUJkfYn4PniD3Xu
YLISjepKm5t5Fu+mNUyj4wJszBV82cKFqVBDR64DkVj794VFumrkQ+CD9CO+
nGrdet5sOJPcONQsh4a2oWhKmckjbNC4AHXhj8MSTq0spr7ZDveK6y5Pl07o
B/ZfqHh2UZVtP3lCKISvoztB188jVN/079SFgQrEnLuNIo6kjdOwdseHLQPA
xxuwA0W1BXleUTjrzT5zDVgde2R4/3YHU3rd05LT6wiaFOv+S8bEL8yzg5yS
lb723w9sMst1D7fgAD3VvfGJn7rVClcZb7FRjUL1MumaO1Fjs/sQYQuZzb7l
rTqxPAUSMTrlYyLEYtAqIjaMtuXI7861ODofjOXjxrIvBlehppO4lpDAytSw
6CQ6C5rqTbyobfSQspwek9c7LIoGAe2g5i5oQn7J7S04t1uIQUmBE+t852NX
Dm+14V2L+7H+x8z+ysrXp5m/+XCQjDxgWAKmCo3Grd/t34k4CTCRIyMWDXSp
8/MIOCyd5ILqKjwxaMBXthIeKhm/MAOSUlAVZAZdJgOW4Zjp/cxegOvNA3Fs
inSyFCssNAJD2xu/bLBudyQoOOyBrn2nNW7DEMpm42wVG9N4G8IRnhc0/gPO
m6sJ122+QxXO92oAsJ+x9D9AjR9A4SE43bfvgbaoEIf+xiFUczCIwi6GpBe0
wkix7uNPn0VnIdPhEo2/W+vBgQtN9WrCupbYNDIBxWMtdJZ6fbgBGLkm1EkU
5JFoz5J64QIAAI+g+oJ0QoIYbj7tbwSuewTWlY0f1iH1GNp6BeQkiTlao1W7
t8rSie/NOmMuRzJXZjzz2QYZdA6lQgtV4IlaGV25RyRJfml4EeDdPE+eNUS3
WnIWMbVUc35ZxZ1y19RWTYMNecSyTGuo6Dtjw1MoC+0Q/r5rOK9mxz2oLdlF
/8VKWFP0bzxA4WVIHRznssXRLQzsEqN+6KSTtr33FCW367vDJe/6WRUMd5a5
yJV+YtLgZ+x8OqP3GyORLi4ABqXIe80/UBX4ziMPV4HTaEJ4b60rj4T8Elxn
vgEZxSCdrZ20FpHW5urbsCRpfwTZrrmPrb5C0dMxoPlu10xIYo6QxDNmBB7t
VcEi32/ZFKgBHQY1zjq+RmjDCkEH0fOYNsVUkzS2v17NY6h73GfUh2lQwt6h
7DSRaEjFKVhV/c7w8fR8+kFpINfniB7zuOpx//yh3jFy8a5NeiX5xwaf+zuM
mAcyuFyxNDfLi+b9ettMDRwT+H3e9NnCz7MjrfjGk1WVZcx6cHYQ6wr5kAig
do5J3LvQiKI7YFkgR6FOGDT+LDaTkxlB8xczYJzuRm3fVvJcgeLuNrmj55in
s8M1leFxJCymzrX2/j05Q47ZyOa/d/1WlcSeNVySnY5qKzEVJVfIItRWhRNt
1PEdi3aoc2j+fKxC1fykRn83LR1U+vOoXiEFpXFjOVm7P2uiY1q114Tb4+UP
BrhXCcdNRJYHoJJUABWaOPYaPzR6MN+wb1FldBE2xb3Mti062x9xIVCIIb2j
e8KsMzQ0Emr37PIiOl1WDa13pX5o3s6OCR78x5EYvhY8sm14+Vge5JSjwD01
SCs3gbI9IqhCPtSumzp7HFppSpsZnWQn7DO+Rvdhlzqf/c4mCDPQYF9WSS1W
AblwsnyorcHnE9Cm9n6n0YqbRfoH5X6V03KYR+Q0IRhSwV2HIPWd6lAvAKN3
qS+BqcvNikiKFhz0Bo9Om3adMR/UPslFoJSLn3GQnHpEj1qD77tpx/PUMazh
yljQ6DOyFtneINUc3GvJjf5bMMvhZ4c9vvgDVUTLQW7asQCYi7JVqVhr3dd7
95Rmyxg3LjBCOaw9mc3cj3pEc3XjGVGbyZwGYi5bldwo5jmEsnnJ6AI5G4Lt
bgjgrC60xWevWH/MnmfZ1Ytfu2rMQZrcUrAfB2bLutq3cl7oUF2CJzmq5imk
6uMzWKAyoY+mNsV3gC/1vH/2S3grZfbkHWFV7r52yquCNpY5kApkq/CFrHbB
k/+ktslA3AbmHY9f5MgmIsurBASjwaXYkxWKyzTyIcKJLejbnHglLaGh0ACI
wei8n4I06Z4QK644GLy3pk0eBAVPm0nMUwUCJqExPJHnq0yv/kEIUEPsBXKd
bB3U682baa7tvsvh7MJBktfEMMyG3japKX4Cu5YtM85ugvOQw10/vbBtY3Q0
XEVPsPWbYbTkOfd0kucD/673YtC6DQIZC6pbAQEIhWOpriOtoksoK9ZfXGcH
ptBIbxMXIwN58BhrXHlJsS9caSzhvUIHqepYCucLfZP4OPsMRKqeRXZri5Vq
k6SwIwbbmjGzM15DlWV65R/pSwc5rnCCVpDE1r6YOMJqjsXNGdKCkp9UJS3o
XvvvwdCl7iZwVLtA5cT61hKXXND2+ANXNjPRjgDfOT/hihn8vcoLCaUr7A4t
AnVhkeDXeWQrAcU060pm2yIWyyWn/5tZmE398MWb8hcl9IHG9UNDzGQbAgzv
27Wrp8BQ0NOoia8ITflQQ5xdudLs7B0QYBbO38eixEpyNWYkAMjVh+MZUO3/
02h8LZSVA9rEHkLaV24IYDFu/6T6rJeVZAMWp+v/QkhdV1yz97XxBvOQ9FSc
o8ksxWKK7ly3t44Np+5FKV1Fs9TEaO2snlj7aqCZEWOqRIXk6lZs4GKN8LgV
zuA8GzM7sQSQliVvV93H9tYJ+Gj42UMMhthL0s2jzEqTNeDKxjMUbFB8snNU
l4gloLq1YEI+uosILT1nzj63sp1hQ+ZKjZLx51dFk4H0RhgdTN2SpWUjLveJ
+7qox2pdBFbFHVGup7070y7sIRMgSlP4kBSfcTjI8fBorYp9OP3k8ZR+uifX
sYpUIlIT/79J0NXvKQnUQ/dfFYvGIayDW2WZBG9HVpHvNPtoe6RRyHRKO5MO
FVSV71fKSfen1bZMvppXQAbDLDwrj+wuo0YYTeo8OtlRQ1Wky65pjtX/wfep
nwChGYn6Z/OkcWDyjktSZZNHQUt5cFkYkA3MPHdJp3ZHDf89MnagrQIS/nqW
blzPTy9FKJ8imIkLnct9Wi8KPl0TuISnjk2KFLM3HNLHG4qmRM0IbeEw5JtO
sjf/d69xePrEA7ZTMKTBz1G3kdWBv8p27oGBgip30RakWlKih3cErYUpEyST
m6nisTiWQ9072P0Gno0P8sSHeZgSmLowxRk+Z8zgF2aAmnZc2yVRLlY3Bk2T
g0n60DuUhpTED3qaqRyOnorf2X80R7nQJGPPwq9znm/7CKIuyLRnwrcnb9Wx
qyRPLZ3A9/BNYYQhkhd/JFcnPQ2NLtFYgr10byc8d1HYeY30HC8nTSNgS0N5
gppc7RJj8w27rVxu9xek30AvTW5B1gNdU6M1dXlrWcrVJvFdJ5HNBFbZS59x
kJA2dEL/9M8lOnvGK9JimrdxdfEH5F7PlwLJrV+Ew/Xe11BWYTXJNnxVz5Y3
4U7Fltt8AFKmtUluSVzcztW4/sTaIVlWeWcOHHIVzVECATNurUlZMc8laYM5
nfE6hJ/c3uwaNpy7Sxbk+HB1iGsrbX2OJG108qHng73L6Gjq4TMBp0og8b38
+MkLmqsUb9IOb7+5fMNixFDWZDPBR93PztWz53W9RtwLMVg8NTH1A3VdqiuL
gJprId6LmljBmDr/r9AmsW3uITbHYNCp6qNedqbzGymIxYJeiMGfpbEnbjBi
df491avmowtWKimJC5g/pR7wZ0hBG8hIUjenPzW7Fx+bSAKe3aAsJ2RQ0z19
Azzz8CWXzhxqEHxFR4oW2wBOKeBjfxOgIDea27UKMfCVyx04aU6brV+2DThd
DOsyzbLsutRVIjwoMoUXK/yQwKAaAp6tYC32sYLJ5rmCjPo2DP6SM+YHBUDn
wHXng9uqhZ4qdBPMTgt9lA+gG1wXHFBAbfc1E6HnccfK1Zye5o69Q047rQs6
ouOGMjPEnSJtEGM70UcMirorNiCWtfhYKvewje1RG0HqFEFZPv3qwDtA5Ht+
jHF2yRIhg8Ylmz38W1BEzza/Bt7OZ7ZnK941SP2v9aFMpeTwRnlDlbv+G1+P
Yul+anK3XyrWgU+09NNWb8ZjdnI+uFzbVKlpfAIG6IYuiBWFu3+aFgiAdlqI
ul+8+wIiPokAEfuvyhIIE7Ws3C7HiAQg8MnS2EnXi7t+lNms+Mo4jrxbRxOq
oHKv0mphrDA5gbpHjL/YBTvA3tgAuBweXy3HOrH0+sR5io9otO4A5CuzZCk8
WpnqWMasZO/NjnQl+1IPLXUlqWPa1K5KeZS0ECxTfDRa5t1POAAna+7uAIdy
MWlsiV3Qn3of1xU9+JptBrFNITgoG72FIqyZMuMdASwtEdnCXIIil4dZB1tG
O5VQsw/gXldjWImH71IFHWIxqQ22WDWRY67YLcZ2SKypxP0fZjvDSvOPuyCU
9J1/9oWzAtXZVxoskpJCkjbTSjX1wPj3l8QA6rmBV4ZKcs25H386rMk3ukBe
o3R6zNOHbmGS92CwWDomiFFL7+LyOQg43PmfWZ224xnpG3TdO55g/IiyscRv
hNXm3k7Nb6pCktgdLWylJ+ScTLb/7cX3T3i2bif7IZbWXoMnhwcf/B16jJWq
xrg3gbS4tl06BhvWrIBXzcunalTXZ/5NStH8z3BP9LZnZUqMGSVIuluIjWQJ
cMGWk0tND0nBBkAjSuNHlHZXn3Xd1UsdynmO2zKWuvwUtyqptWrezS6eA6fR
sG7/grskYI+SmBBzPgoZfPJJMg6uAOhR7hYVrkSf43faKdOTWsDxvS3UEMrz
FZRWGcdBMHBJMge0yr5AXaJfYFXW9WQxu76HkTZe3Q4566qEAUU1t9xX5NeY
ob+DO0g8t5lbSfLi43Fk3kZLUEaoOOK0zrBLtAlVcZxDfWC4MV1Il8meF3Yk
SBeAhGb0oMAjoDM1hd0HgAavL56oyhnQML07Lh7TicgF0JnJpw+SpiMZqNJy
02x4gvG//1y71FvTBteISGBwnUUAstz0hgBG2Rar14VzXo8yJpZNdNeH7gdt
zIkeEkY4v8vopS8f2F4nQ9JJXnE9q4ju8yIfMBQYfwOpl0JTTbl36+WCLCFJ
WHtEDYEJFHt9Hl3tFViedUA4BBKXLqu84J63ePwvtNSr8E6ACri3D1Tk864A
7Kj3mQPaCvu6mnkUmMlOyHNKhdJBN/ohB3zehFzO/gfi+95nah2U+bw+eM7p
K16PTeZXrow1Bs77FBxHLBF6A1Dle26GNW1n6Y2yShkE1q8WH4Tl1HfbdJn0
syzzPoQBHmCdaRU41sbUYU0wL13XT5I2XAYCqg6ZzseWhTtLarVv0R24qcAk
b//ESfXBc3CyrYI2BwN0ZLSVDDc8ho3GBp4Yi5UvheN6mTbr+oY0D6nB71LG
zbwr/QRd84FAeuaBvxezWBSg4LCID8ww7i7YRzkUj4XGz2C1kIdxalQNxPmE
5qQ6Ms/bAJ6OBslOIG3FGUg/3p3RZ2uBO9Ft6HMWhZ2qth8AEPNrQJG9Dd6u
xjWB6z3WQyqhGSdpuGlxcYfoMicuIzu6URh76GfnC1hamCGagEPRL12jBFNc
7ivYQG9jm0NDkk0Ba7Fm5mlD1is2ZcgHLlGrUd2NT0lwdGI411Nj4JJyU5EI
2I+AGRt0lP9DiqCgtddAum6VyTepJ0Jh+Wnf4bbn2EcaWFqeSRSJVPvXzwjx
o0roMxD+TTtDpoISgXEC+3tb4bZuA9Zr7nr+mykpavbLrVItsvDxw/mSHXhV
JgO22LswDlT5byec9d0QaSLnjflx7KhpHJD/s1C+jJTP9aRzvrw63WUZa2+k
WEz8PdxodJss5aiwZ+KxzIOHweHhllcLEDDjKUDgL0CKqJLhHGGPlNQnTdzZ
JB3zqatfbI8zCX0o1QqT68WfwwqBmTjjlg8wk4Sxzd+dO+U92uOPaMkUJUA0
mtzjHmnC7LtaCWz/ogucQERkKwVkGPrJV0rYmf46GqxSIdaZKmjx7WLRibEr
BRz90P++g23K3Y6tzTb0bOmV7XeNQphCQK0KOtN0UeqxmPTF7LB555xdhc10
eqVA6Gor29aoMPjsrlMeUl3iksXjsC1R/VWaptOt/QXpCkfqKjGLZlw4TfFg
K/YbObs0dPHSY8I8sFNaKaSB7FmjxIJDroT9RQgimpPZVf71ZpIwmgx+10gc
aWbiw+y3EaXgNgZeuou43BMq1en/h0FxpIZu4Cgg9BHsEmjLrXwK7yFCs5F/
KxKvGlIy8p0TI5ct+k0JVjP1HImCy+3GtMJ/0M0ev1BW7JeNirT2x2VzJFGq
AhfWGxfKUPgrBIZWA+1FbN8qlcICOoEGPheopUQIOy2PwUgU0BuK+3CHIf2m
NxXeeeFD40WjXGvNFfjcZoIc+2ByR9mNDZibGhUYG8+QYdqTsYzmLA/M1c61
FgWhF9ue0w5s/jGohK48c3c0t7gBfYIXisIFs7vaOQuFK8LTURZdH0XRnlTn
7uq6QUFnpbiKxzQO8PKZqVT+x2yiJXqWpnkBPnNhTOCrN9Fyr+AH3/alscsQ
zQtvMAVA3UXSYZpU4xGz7gpFXrh4OIIFjmSMngjxCaXn4acYppnDzpNw66CI
IP0Z3in4ct2mMt2QWQNVJDwtEn3s9OVF+LWXbqdsgZ2JVq2/OVc9zIcbfBr8
UB/BtYk8EXbWS+32KQpbSSH9O/IzxDCLksSy3cU5wQRz/pi18Q/c3zaXUAQo
/h5xop4+s+Ew3HSN6BmtVXtXbSrikbQSJAhFAm8JJDVtOKp88FVGUKl27DtS
9aFpJppjOaSK1bTP+1kI79m8gNgq0rDT5Wic9Uc0wQ/lduadqIrKRDNJsf3U
soz341Xp74imxK6aaf51LqD4e1nhMpTJMHFZ5ybaGUFgEWh6SDI+R84r/cEf
y1d6MIgpyoTKNgnqiykNpR4c0JwwPERGUand/vbLijMrccIOwGwRNbTp2Mt7
DGLTqKG0pKoyRSe6vlDD1WbJKBHsfxx9/3rbbYLDLvs9kIYS4uQFkZskGUM0
QAzuBLRAJ06HVKg5pBdzKTIlLoAEr54neyY8gEXN5mBX56dLk0jSJlNg/03P
vjpyHiuHnVyMTJZ6j6fn6+b1Gdub4qpGKKOYsMhwWSIIOjyUSGH26FnRIstv
rAoYjRQ1MaKwnzAu7hvj5gBwvwBo/HC3iCjTI7jmVdtUZHXu8tJ2DiFjOMLV
clc1giu7xqwUGszJb0f35umw7ME2iNYBeW8ua3M/EQLy+WiRiOJDbxUdiV6H
SfwjBb1iZvZNlivF055RkNHeodHKEneDrd9jPVnCBH8YO0YKTF/6S2ximfe7
vRLutJazwpW8stsE1nJmoWxFBPZ00DH9R3aBYQDHqj+amdykn62NtU/c2qdw
81niZcfhSvO/Jd1zi1ztJVUkA0DiXUct8pmkuLOH0iYDavd2G36Apfukktch
q5NzgLQsmwhKb43sqQihL07EgoFg4nbp1XKSsdXyCQZTk+o5v1RUJJ3SgMjL
UD9WgRkkF2QFkUDBLqfK3HdpNnkggdaLBitX+jbTy3XsxSSshH0vqe0O9DEy
yfuRSSwwqJbuUAYWUkv5EnIarjDrInFfzSg2nvE5Sx9VSNoBanPd4R5A53Qz
NmJ4rkhGbEwGELDuitAjbUuFk0nzRe6KaCnsgeXnzTN4IwdWUvbsqjAr3HSp
sTCn0/WANKRLyBPZyl9lF+sHGe0r5VLtToBV7YFP64/M2Tpv8T/4LyvOeSLN
wg8oWfPINIllUFUlxgppCvUzWSMF/X+1hNWPk9ZBXKv1ZRBt249kmM/jpuMy
/lz1t0lgz3K0mavDIyeDJDkVfXkzzMHMR4l2M9ZQUdv40u5QYxu/4KU+BhBS
mDkLqhJ9gSnKLKoDz0FfVSRlGDyvYg9Ps3PDBs4dqvGr05yxEvR/1JcORb51
qQgsbMgZgk8AXGn62prp1qLzfXYoORo8rqR1FFq3RGiSZ8xddz6QoSEB49TI
Ci1ZxwfIMZSlxvviR3rnS8SVgp8KpKimPHzrzFod5EWQVgoJo84n99jf+d25
9Dmmwf2UEGkdJ+Rq6+7MN2nfUgCAm5OHPk6dctkQZNR2yC1AzYEB4BA2N5O6
KhassKsPUSQlyFSl/rXzeFtgLcS+x14yt7hi3TvHihby0Okp4f6sJPVfnWZS
p3vItt+2U+P7ZQT90uro2kz+U0iLKakDIW01jC9yN/8llVC7yDTUDgRNvN3O
hqX7cNfshc/4I+2A1HYXGbcSsHP1/5NDiMxcCncDLX6C+kWnegOf1Ot9vNda
iBR+7a6hqhsyH/+UCANf30D/l0TxVESFfbYIyJ9S4rkbuoEdC7QMrsyzFojd
alx0xHpUcgIZZu06UGnW94GSAvVv/M/iZy3oa6/znQlMOiU5Ta15RL2x0+ob
mTWZnt+IXn0a77cE52Zplju2V+24Lbld0txrmXbLVhtZj+u1MfBufJmmSKeX
qDv2ey6svmr1fPwuzQSTzTDXdv0hU16Xj7XLxBeoJECda9aBwhAgWU+OrLQX
2g+p0AsOTomvFts6JCStzCs8REWcJgDazKAKvNiru5LiAooOh/rrk6ecgmr2
5ZQS3yAveDiqLSA5C11c+5Y4pmAtqJiP5RgzkmosXcqttenyved8jFQAg4AD
e+Yu9PJHRcSTTTrJSfJdWGNf+oYtNUIUvBFjhCxbb6Q1ej+kYu1G7u75LO3Y
UHPpytB8FHOdD8+tQMtU3p1ij61bE9TSOL+Z66SeQlUvXYZ7xaAVsj/5Igkb
8bIWPUAmcgesDUXLvYWaNoXfUBO7KzXryTcf6g0iG+ikt2yirNwHZymCPDZf
E4K/Ti4MaLbgzTt6YF4Kji3to9pzrmz1rgEoJfPjCRINLKFo9iZviTe/6JNt
Uhb8AqM4ZXrLI5if58oFw0g27dR4djPvUHNzczlKINEJ/AK5WxgRdx/5vHrM
bwnWLTsJ7Gv9BpTArHwuwUcvZ46b3Rl5FIbUZn4WPCvguJRQ92ktE+bTmaUE
jWa8QzJhAtmFZ2sDTxehHhdLFCZL9f5g7TgUMBoWgv8drRe7+iL7VraA7iYA
ZwFovoR0X44uji0d82AxaYSbheRiKv3rLVsNOfiS6Vy6OAAh74UfmCSVozb8
x7pus+wYchlZg26f4BXYvjFGH/QFXR9F/b+9draVIecWLcwNU763zQVGQfum
SAgETVYaWxfoEolru2nJnsR3NNlbflWxl3lMZPOe0O+M+qe1oMrNqc8zmtY3
tfWQVJeTu1xDhLG/JLGd7tQgrjFfxw3c14dxBhoyFOdPg4dgCaFo2pvDGgfW
g7RrYVcM+A6AWHY2sO9KdHDE7L744yLUDeGHDtd14Niu9y7rc3aXbcqqIkji
TEKrDMOUiz5wvplFBeBTv0UosbaxvKv46mWNOyrZjdtS9dAml+4dgkcR8s2e
cgwo6ybUabQYKt9rn/9UxPCs6Ssw0BVxzmFmMk49jAek4suOHT1uIsm62gZr
1r93nh9WglYuLwGF0U+cnQhZ6qmHo5O6juLGh8A7DwdoEVgDRmhire24C+lH
siiQA5Fd1ZsF38OVQsSR6Y9d4XLX+bstrlmKMQEOWZEnMKNiN+Ews2K3evzs
b4Mw0qL2njrfGBqxNn/B7okjGICFbRU6tZuxQIk0ojoAj0KRw3dn7R2Df3li
q7esHSnQUK042wy+D0j8pPObdj9YxAm1SdK/STgxrXmY6jjQXCszVZEH5UVL
0UqrCFLDAiU5/MjCygS3sRNd9eYdqazpxtn62B73OaIf6gG58p83vNlwxUd4
oqoPcrb8GgFXstCI2CJHZl4ed8tIvr9YSXODm6YRDEXJoLUpV7uQfGKqAIQe
0usEVkePy/XiLkMMQamkioMVox4CR4beV/+SI8QJnO9xWrSahWoig2EHOI7X
eazBXEJqDRuadf9bUjumWpdonrXiz78lkXkl5RYZX/J3ovg+vgnoLDZAPK8Z
bU0f8spYmdBf1vtmZmNqryKGWLq8qefclo/FYwidtyGPdqD57uULYEZQotN0
Dwt0EshIKlY6Dvsr1IqctFuaXvpNxLQs/syjTe2r9H/kzvhURHSiF9uXSvSt
PgtOIPXerXmrU2s5+iEEtk5tPNlAut5ogH/R2sYRYmVZptLhxLuB74Z+StWV
9ZCWCyB5zureix8sgojUo//LcAnFBk/YL6JvPlQ+GXkSiIY9rhOQvn0EFNei
ccFl10nK1Hs/+HmQqIMADawUmd2hFwgPgHYj/7201K64ZjZ2Q9ULNVtvnQck
zkQrIfCT3N19VkdiM9h8KTnEVr5IsqL7cUOr/Jh9xXeOUrYa8dXgpRx2vR4A
OGBRk/hB3PQEsQBOr23opsMtkND0H+6ah1krJoeHiqcR+3+bwfS7gajIvMzM
cGMC5LWkbonaOT7ix13NODbwtopnUTcNxWXLr3ftPYIwI8hWpUjdJ4RSyDcL
wzII+vzpSOReqdsLTZ9guCvrj4LyjNB61YGj/zLrQ8SvsjxDtK+X9LWPAe27
1BZG/l7LXy5znvXwwGtnfVySAT960NRd9Wp+/5TziL1wc+RDUERhD/f5W3Kv
98l4yrL063Pp/OwK8AoKsV0XWw69LG+NwK8AQcuaplYWuEbcCXi3FSL1uevM
ZL9xsbgZPa+VRAK2ZYMZ7awJ4seJ3SW9Ll1QIW94ZkVIsEzTzOBlyqtfJzov
pb8fjnpYllVm8/+7Qe+CbjqxxxAC645JLvs5fLe1zNlhjcpyOPUgYISqspXM
pIvLDH7/Wq6hvoM8db/Lt/G4s1HOjaCeqyyEvdoSC8ysIBQUBbt32HD5xQRy
qEA+6s0MNjKhjqL1EJMxnFZGuBo9F9ekkfEoB5kpA9DX15CKfgRvg9y1et3Z
7u93KZzU4o3zLLz1MF5snch0Isc47JQqSTSLGZ8ykYbX2RRcFtHreJfFbUh3
KxkIxwQwzH3pYPtMC/Srv62yJXX857H9Ljr5tmYNM+V2zUyBx6b4uHpP4eGc
NZsnad6hAPYGVwmDfPPhTEAy2EVUNp6ERa5bE7N4iNN4hV6kYIq5RvDQCIsK
MHqJg//2CrROxkBAD5ItPKl+0P/YFLSCxyjxXLLVzrAan0i4qdRiP5B4dshw
D2m2hOyBTTW0r2jf6X2lNdJmtF02mGnM1X47DrlyAWkO6CjeSC5Ul/3DG36w
t/rj+j4h42uYK0QHYqQxwm1Z00r9hZxFOS82rPQUhhqg8Z+ccLxpeuK/NGjg
nXemN2rKuuXiXc5EZssk6LNYtWH1sxIU+PKMlVtjdDfe41FU/RpnxXGbJnxT
MVXOCnRmeKAOd7IHrw/yfTYmhqiadD9q3GwXf3+Bb8DSufCtP3cMPnyJ1nf3
/e5COwJlpFSuDuZ7lujNJZ6W6Pfb9bQNZkooyLtuyXHpSqFg4fKkfZcei3G0
94tkvUH/5/FNmjjwLxWA68pXGBytN4Zy4rZK84fdypkiI1EOQn+7jJdGQxgr
TRnu/0aFs5KvFcjfovGmFJBrebdO0il84++v4XkXz/lfP2yBZ8VTc/UQi38q
/Shc44wqwXyjpJMah9xryaxGqRMe2Q68QHvVXbSZTPx90kFmxlafnJYtZBiW
xKFh0G6+/eO3+k80USPYFNSPKVqlJ+ZPoYnwXH+As9fPUrtxDbkTr6eP2RSf
mZXbPEFTto2xdUrkhnkGSBrFp1WibZYyyL/W+SvCGHUGT8RoSZU8XC9do4lk
Dv6rNvkamg/MsHctPqguMHqxnV8i3+1N+lQ5pf1sJxsUlZw+T4LSaS0EVU/X
eo+/jNWbk/STD4D6UtOLQkUhnmP1Bk42mFv2evqUFusj02FAMM8MNpCevFcQ
Dmc5Q5gTRXfqXnWsAwwj0vCSo+DUVyUPM2uC23GIAaX2YkUhunULJiK0w0e3
oA8A/QzW/jq9M5rDweMbAxJjsfVTiezHCoj3yNWSL6MCHOb+BIX4yOczK6LV
l9s+bTmQ+1qaF3CZBjXuh+5T0tse48vf1lqeRARcfBtPYJMI+OBIRStfm5KH
1bpgjog3+dKpyhxg+WAFbsz9pnYIMaZFM9+odmMvu+A+CNnae00Osx+fB5Qo
v58XXyQoOfpK23Rrky0R39o7glkn9SDUILZyuuRgpOHSI5H6F1hLanlYI8vD
S+I/kQGTyAGaINJ8O5OXppOmbAihQ3qfJxLwyF+CNgpxNYLJzqvOm89AJCjg
/lmux7Y8HQ7bM2RqomuYhuh9Z7DpF75tAcO5pfDlIwF4BWU+S5MfnlwciqAr
3WhrIVjdZPdNIGCbWVf9TRn13vC5bwBGHZEtsr6qIIJkFgJfyFEKILFtx0wu
CUMHYOJhHYHv15PQ2JM2b0q0cOd91ZecjRStLTOkPEyfDraN/lP2iOgoWLqf
A+w0QjGbHGyzJmyIxrLAqe1pAD+O/PR8X/JfIYjHONXxwuPpx0Zeia9md89g
Uec9/LByxX1yhdCz0GHcJW+OAMFigCpIEbQVvfDLuVFleWpd9fEoTRjYQGl+
2vdHogdAV26W8DLYx7Yg+537gHHTZ5jwJrRyHt8wBnUkBvGVf7xfyCJ9N9hD
sUjMiqrN80p0nGUVEAgH7twwJh3wSWqwxPfA50eQ+Yqs+1/MSNnBNLKWvhxJ
eD3cOclsDer0oRjZpCowQ7eeTQBoEitrpvjbtPBRVPmZw0DL6vwoUU9Ug+OQ
fFE7gjoBxsg0P2XDYYOgW64GkGA8DlUeoGmNzSAvGIYANYCxA4Z8NQ8WhjMN
zb7ynAmjvADP39brtjL+6JAbGYF3ZfSpeAQUcvcuXsMXCivJWPDCIpWJI37f
hl4Qy0yISe7z6doQaujkSZBpWFHD/Z6Ivtm9LCguV2vnlAt/8vdYeNSjEfB1
AwqLIHAnymN2XQ8XEfFJQIsosZ2/1+eBJEsKTsh21BhUeWyx9uPYqesm4YsV
yqx8hhZHsSmMYIIYnolBJzf1EOEPnx4sKZsgJ5Xi0pTWKDlrjE7v5oQq+g4U
Gil3yS9pdIjH0XsQemS0pXrLUqqiLleoAJ9FXny/VhEOeviTkQ+5tmh8kAZh
9390Xve5dqZN6oUYXH2ioeghGqxcSK8HPFaMp2FOYA4yzsbHhgPc/x6Kh9xG
iDQw8kGOVg97GKyCLCptyJbWA5W32MY1UIeM0DWtk+TDMyLZUjiFRnyo9+Uu
k4RUP2ax0ELZGSDmvt7X3zjK7LVO918fWO0ZIPAYS+HjqecxMPxue+lE/DC6
e+X+c4dUFWlEFGI241AZRFEJmpi5c8Y7XBEBm8+fcR17GMWglXxyZmJk8ayK
7CAJyjPjDQUv+opzePffc63xcaUPbytdQQHV5wp6wOLTTt1fWCwjSHwf8wLu
49kI5HvDW4OSb+YjacH1LiHm0HI0aLaOwdmx5qHiQkJ1vUnR7iXFOlbgXaNk
mGI1iGhurHFOXTjVqlBF+OenV0Qp12iUoxgAuoZ6TkYZWmCzzaaJlYtPOVYE
Yvq05ezQt1e2sy3gQ8wLfjRhbUSgSdkwqYm0D4Qr/rBUTtL624pAcnM+4yd2
tfU2uLyu8ZRnJ1STqfktldtnNpnRnd1AHb7d7hD6obfrGiEXs436nfrgEAeJ
LsRUkFznSrJjRLl5KVDFh0QFNdUfGOuEWF92EsP4Toxh8yWT267CSx2OojYH
IC3R6j9XSJRURnOgUGLgs82xVBnibBo2LSzUN/2/nR9eKR7HM5HrL8WlOHeP
fyRXlHpGSfRJDQiLk3pLGj/4OBYiNfIbIDZBfPZzkk0xxm4PCD3RgpeAzJaJ
iQcB57uc39hs/xKVclvxCUvgweL9iN6kOOVdK1BxKSanqY2QQ7Lnmm1nd/Na
R1C5kiWbggcmUk/rzrgD4iE/q78puJ7EDWW8qKzszA6GxZKvdzk+bWIfrCCo
c8ozo22XkFVJqIMSqNj34sIthsSfB3ZlbCpHYc7tl+F1iYWL/qzwWFC+lowO
35gnlGmzHLc1pv5QkYljLfv3KYbKofSEhBgI65k/bu5C14MhtYbwEv/Brst2
jirKgm6mdkGUGfbKeMCGcT6iQD73irzS9L0cKYizlVT1VAZZUvVY8NjQHkal
78jlulYwWxU2A2NmeY1KHNxSDJLMmRO14zd+GXqN70qPIixAkexJ22cAYVrb
SzO/yyRY5BP3rNeKaNpbdB1rBoT8rlC+xDCBWXO2N2uctsQxEsRdcZzl9NR4
IAtsWqot39M29C7pHK42Wm0QjH/6zQ3GmQAD7wQqM6CNPf7vsFwDC+xD9mr5
SPlpfMd2VBk5V/web8MD1RLIQO+tz/+DvfwiOS8kpCpCbAvkI0l7sAMKwt9H
wMMELmkHewL+QUY0RcB9T4jlDCdhLV1No7iAJ7izrEtYrNM7KgrQmKzzamDh
Q7z+FNxK5LJLDKa6kAp0khjSKt+sygYQjNR4NRcxC6zNqTvrRnfqPYMqnaNR
JPMz1zSB6t35R9FMwTWaYQCssljg4Mkq2p4mKcixtuCZtmdbtFXy95+ruIEB
mlZofur5psAnR1rm58nZv7cohwk//z/15hIO5SVaAPn7xuXOLpXw1H8oCKxn
U2IIPp7TVYQ1oIZNBvgCaTV8lhRsDWfUAwliNhTgll0Qo1MXW6Gw2TJhcpLM
h29RencuK7OVy5kzeDpUONywm6f4p47Ky5rLN2kpS+EXKrWWTENFsPifwND7
E4awcYx5VMe4TsmOTZ/GRQeIvfuyhp/tseXEE0hEZfFWk17XV1PgSLn67Zo1
gjEZ1QYJaHi+GZOiCut364mz0BbfmC+I7Qe7+ODLqFpBIzDHtXp4IX1XN1mz
I6025qUR7bmvhHzlvD+Iu/nnWa9AMj/j/ZBY9Ilc3uUkd8trXJXDlty+74VU
MHkT4kx+83Gq7b1/WtsYJHsLK9bxFc/XSydLTV5JGobfHDyeqhkhdvMN1e5F
E1VOPAOACUw/JbJfS3/HvdDVwTi0RPpDDA0jPMbWs5O6ZFw9XnhFi+1w60QF
80Pk6t9073OGnfgqiYyJEl6Chzi5PKUvAE3b+fZgo1N5lNpLe3h41kYmoEkJ
kh2Qrx+RQsVxiX4UhFNSjx4MnVGscozOx4KTXzszaQXjLdcdVv6icTohQS99
rld59M6tFchFiC/wCF8VgS155po2oY1unSLpUg+FK3szKxJx13B9QsRogJcN
Jli0tuJ1AvjlH7/XVQpXRqybD6tZkYkjqkFK2F18iGGtFA1a29uovDdqAFZw
lEMT4hIUr7DIoY0h6aSl4aiO+rmBJ5pfq8ABCJA7Ubb6ZDgvVr2P5v47xz1i
BexCa6kF0xh3ILtQS6WncQtwiXtldEHRBuOi5jVECDOUJX7cufZZOTOzWEFS
grdOk6npLIlkgGRY6NTcPqo6fqNsJd4msRNZJC7n+BrN89wqYjfoCdJol5Gg
DziaFbekJ7RnYuB3h3m54EJgzqIJuPSJb69MI0Yx3zP1/LJacGsmL1XMkCNf
FVwCJXtwDeVN8n1UoWK8dwafeIuWFQdx1UJ7WgqmPl4gqgfd7t/LWA3+hnNJ
iwexFwqHZMLCvF3cEoRVDOIZ2xXivmQxHtNN3XVdKPZOnZCQIWiAasNDX97S
Fb9yn6FVADYWl/HsEl/cIZp5N1nLtM3UKw9HDryvQTJ+Fwil8sgjU9jOxQsi
zjSZ+nAFBJfhX4h3gOVZadtEcDg5DGNw/lCIEFbLjrLh8a963PygUoqlf4qu
DIJJbtUARreXMAe6rs4E0euNOpDkUrQkYr2Vsk2rJ5kGmDafpQ7Nnh3YiplV
fZ2uaqLO01rHqemdq/+W/3cLF/0NLuGbB2Jr9niYQYmutbK7p1MXc1QJx8+z
9txTfDlLo2Zljt+TA4H98zwZCVkdUUda3eSUqX2g5wOUSwCuGuI+AH30D+HD
+pLvr/DkffHjtjQJj9IJGMjd8uhg4b67x8DTNkAOmIVYysRx1DDJN0vNTz64
PkmIM/f6nxmunSjsSvzaq+ptuKNnvbYMkV98j7Qx17EqYtRcob7iMtpIPlw/
OiXHynw1m3BsT2ONZ/+m3WCDaFF3/eXrKvJBg0hkUvDAkIYDL4RXFyS7msz0
By3eksoDrhxYMt3P3moeCj8BbEYJTCd+iJFKER3mj9AmRj5O6duIPAeLCh7+
jr3BSYOPdau9Qoll/uPhNvBx1z6/Bom5OaQ+7NfaWrdmvwMan1UGTY1740Zp
AgfIQPJJUO1Zqrp9XK1WYAmoIO5w0ZGaUB0cEJ5h3x/K4u549HKK4nca0HoD
jXQdbX3G38HNSf8UkNrfbUMO5KjbfD9Z9RRSDeH9vEk17Z2ZLBfn79SgyWDA
D6eEnZhKAtHn4RSTj+7nB6axKQkppIeLzxkZeZPKPR+7F9Zv660xiBBifmwE
6yAxCFddRnd0lnODUxuCB8OMK22xxzKy1rKNg1re8nbwS+6hIP2tCAcPTx2O
FS+dBZlaZmPHzUKF1HcesH7VPNUEqdES2g5wGLF/eFebccyLHYTS5k/S8JRt
5ZCAFLC2i1ERvV2Jkhr8IS6EeGKagRlt6gtEM+9V88fwRxYFjkTxjbP9mrjZ
ZECvqQhR9mY2qmVYlBNE5yXFb8u3G1TJtiOb6EsgtuWdKEfjXKzlPXYH4xHL
sdc1PPsEX5o7NOLcmvhJmbajPtuQN0BN/tNe+kOXu7rt/sn/GEx7MvOjrt4Q
7eZ0uWBZCcGIY7NUhX8/Qt+PWj5JkynB+JkfPQnoaTWVXW6MJnjx5ZzznNi4
H3xXB/VADCMcXX9GlriFxA39fz35jz8X9grlogc4ai+F28Caecym3VbsiUci
HP/tBeOsG313oCGDuHNUCgEIi9rZeb9Rfbl2P1yyXGE8YGPq++HJg9hFZKKF
Dc8UTu7WZGIg4gg2BKneAyY3OJWWERAWV1GLkaTBm3Q8sJbOhanTgmkLwgLY
QM1b1HyOdJ8RVmMa7lCur4DmWtmwZUE+RJ6HpKAlWcOayHzpYLepExUC5Y3d
SDrljpSITW0fUkydFbncp6hXi12I6Fek0df6ElkaSXHqfGqn6NDW37maxB6g
qgNyfoGte2vUiKs6YRwDBTCOxtUtQQ9ZgLwwVH8UQeo7hzmi+oLc98z+YcLF
b14e8Yw1bLNlmSqnHXz9QyJ5dQ4wuZm4OpSHrodSIsDrO15WXw5pN3Pbkk+4
Dxz87WrrwcajVSisaf7PuKpSaUKSMUTbs1oM2WKgJ4EOnrX2l6g15/CPeCov
87AeodGC8CT0ldrfOWtlL/kWG4iALDDpOxSXfE5AjNb/gG8gxqcPdPskx5w3
pY2Na5vzghvZc4qufEf47Ekln2xURvFdnCXOp3VIYW8KQDgBbWq+Ng+0+iP8
biBrxHB4b3fqQVLSIBaIiZZffVpkn7U401muIkZveGuFmov11qPvxSl2vyWv
rXT5slv0Cimjjk1eGgQ3CmF2G+0mMyEG4Osf8Wwqf1BBn6KySW44BU9k6mv2
a+Zr+GtUbr95sMLyeC63tjeaBs0G2WKB8Cc00y3r0bdvkZQTEYz7QBphLzZ5
gWdoxZJcNjn3Gf6TFUAYhtW75ltwuMt+UD/dYfZfoJZRLubl5Lvcw5oF3Iut
D3Vtd3ale3+BK3G/KYxd/6sIqqIjBOz2Xo9i9SVjBFMrD6VbDfxl+nt/HIEk
Rhf8k89kfYYam22WXKF5xq67FJNkAKzMw1KjlMGWfM2qjtrqaq17rFo9OzLS
rQocZ7VaikfwapBc+sReqZqqIDrvvu+0AUh441O/ekGOBs+U7tWC1tU42TZv
g/R8aS9jkg90AOvXYv+DUc4IebAye8sYQ9PD4aMEEFF3mK7ks3yOTQMWoUnl
XcWnwE96ovjFodxmJO3K3J5gIdue8LV96dUlacTBGy8VHnYXu4D7i0kczNSw
jckpfiIoFglDFmijx6+izBPhJvoZduhJo9Rs5uNnyC41XZvDH1naMKOqb4p+
CrOScTkpGraiqp+RhktLOypltKdr/qtHNpJcYCEoC2xj1AmKFwlzGdo7meLe
/DiP0pc+Kr0lBCsz6cj4JsPdERDUWQ31DAz2+jdhPL44Wj4i7fY0tWdLDPgT
CDmdjgoiNGV2dWCzrhd2MmlVMMPnB9bdboEos0fYJ/2oC9TG1tAZsHPZ9ror
qyWDP6GCOrFfrR005mxx0mlMlaAI+DiIrtZsrv46YrQaUYWP2MeFK4zvJBjz
17VPCx5jf28ogIjimr6JP9sCyj3NnofUiT+/zb4z9AffiLstsKyZrINKxDcV
5wsUzri9YC7upEuPFin8lz95VrrXI/sKvIuWJI5coYtrc77GRFBGT0F7PJvj
twyNkJEBya8RS/hebi2GoslnLD5AcWjxVf/F2VHIC1lxUoOgEKkBNxek2KLV
j/GcPH+r+kGuE0OJtamemKEHs85bkuv9+PR07fcyFJ77N80zfrG1lpxLf7Tk
2qOZDKaGFjdQ4mVBBM5Vk2vb5fYz5oHdnoRytYFnWsjfg1QqEw5ZsiMUyRgF
kQ5M6yjzcOWvR3oBSIezW7fJ3vt3nOadjamQ8Z2lOvSfw+zAH670NBirY307
wF8KFlsJB2cNh7jYzMAf6RUJpWkCOAgZ9cxhGnJkgnvwEDf4vxs7KR7Xfp69
bUpZ/MQnjf5R3UvY0Jxej4Kc4+p+QVAILQATdC+7UCLYoGjujapzqH0AKvM2
lKsd0WwPHA8fdnO/Oz7shiirY3f0JjCPJBZTaoGz/ZVwnqJJW6oIie6QV+UD
5Fmly10vzk3hR4/ILHfsjlk4dt+qrfLsJSCCUxpa27TjCrJgLkweqU2dPPH3
sT0O4DoC7xUfJ/TN95io22enxTJnOKP6vazkCd8jebd01LPVcqFFrV+x/zT2
uXCvkqG8IwGvan8Snnv2Oqi9NN60/ysRGliXiJEFalYlNGJvcopeGDKwEdlg
Q5JeYFnIUm8Chyt65a+qEotZGd7zJNkA0JuJVF6hPoVIcqjGUOGuBBPJOCV8
ptTQN3Dnoiu1mm/VirplOVCIgwy5BAJMr1yx+Y2Pryy7kFYID2PAF6i4hzma
/CNiky5zJcmVaRTJf96MK+qk7AihBCvRmwQxWrvqBWnRgedbNuLsFltjA793
QDkPZ/zno/DFJxQ0nSElqoitFEHd8bFPU3HxwONM/4zU7Ya4RT99lsq7Yldq
xQXtGvKb81ia5bxDWKqAtDbGMrRD8ofCecKwU1GpaovKpuUlUQfqFaKJsTTY
rKnAvcE7C3lWVaEU4YjcPBt7rMTtOikI4EpQzs9Q+G0N4bx/+f7u3XT2UJJj
huWQObAzcvPMjGUy545wF1HP5EQSNWY2FOjFVqo+nOfv1v+3TPxBl1oTXjto
IOSUnCqSrnLjJha4KLH99TqVfIr/UzdL9caGLsTimomFBjFfF8nw62Sx1fKL
YyxTEl0zNTYWWXHC2VglR6oFfHWY/NpU308WAkSKsmRpjaoXalxDLY+P7UZL
4UuBEMCYM5MTGwSytOiD9lyj40Dq6JJHsKipuTOrHb7JLHIRY7Ku19moz/w5
xz2/ueeMBvvZ+Qv54WYGJ0cQukj/6kt5Mhd6afgGtqqJMCcJ3LMCfoTQ1xtQ
eVMwH7eVrBtLu7BUxz3S+muYF9B37FMjQxW7GhzHUvCPOB8GfgMenEtgoaDt
AO+DFqQ2idq1ubqqs/WAs2XF6+oGXL72IlPpGAV6g+D3BJHPFwnOiz67NFwA
AQYvwFg9mItDewbm9mVp+p644SOvw7rcjRo51X5UWQkoF9gK+PogvMYT0R1l
Uj+wpmrRN5Xz6rVk1HOiWiv0bTyewXW7UE2v+KVEIJ6BafNfnYXB0nqwlz0y
C0ZGzzC79ZQbXRvmBhd8OtvCNDDnfbqc9S2m7DeKMiN7oIKFP7/Wc4AU/6dZ
GD3L0fsHGsMVUQtqyDjdcZt4z65f19pXqwBGl2V0ClXro/JH1AohRmIRhJuX
qpGmSiLKlznAtt9Db5XQ0ZWld14DPDCV82lssidTOteh/twcuI9kYXYlIWQi
oWDl7XX/aMe2pnpJ7M1I1dS+TrmiNrAdp60Uqwr1+dhcnUkpBTbzfOOghq1h
8vov02UequJWj9JiwILheLN/98+GFANjhjn7rwXLET724iIviZS9q0aB5dPP
dojxgBOE/3/JVkqTas6xniObF9FZsJSnGpsD7XRb3s6KySHjTvnvx/GLle6x
S33tCqVLPgrr/1GlJbGOpp030P6oDtfS+kt53qGbfDhSYNlD85RiHzF3bz6d
vTkBkaHx/JAaSFuLV+mukK1HBc+sbVGA+tTD/kPRkrn6UEJoBGdMvN1EeuN+
Ucg+eLSyi+/cDgGMLZjOThLqv6LWa4Xfv8UXJJJHh6SyI7b9PedlCDr8NrIL
H9Wm7NSnl+o64PBuFVT0TrPS2KjfXoudX2qoKxQjaGr5BETVjht+OL9PM4Zj
jtRE/NRnWJl4GYd+TUCpEEXYwD8+pBA/cd0m+LVMH07qxfymsP9d9gMMBorb
CbTAJxDCeik0inJRCJh+1OILNka5JrP7HmGoD1ZNFIlmnSF+jVHoHoVv7G4i
ixWC32Jjho0ff6YFA+hUK/9ZLVPqJVy5CmhIe4iEvV/NSkcEO7l4GkplLkti
/yClxWaRvNoEmGC7hcaiKE/qasH37d7IyQlsPbOBbfmOhdAxesXEGzOMvKrg
yUCJuLUQCd1tKH7w6eWDZB70Mdl3T6bFj46YfTBBYdLAn2YvkLbzJ7q4dT+4
6pEE6eEJ+EnS4s04mP+Ri6Q/Lh0IB+/H/eJkyO/Uij3769PHZr92EZ33lgZp
fbcnPqG2g/tRPyuxXXABhwPP95lq/UDsg9eW+eBE9P36seRFJRQczf07Y3Au
kYEfgy1r3nvU7NMKsNZWPu5iKmqHhLpJKiC4foIEUqwkqlUe1XWKK6BDSq5a
0h7op8RYgJ6PqyCK/xGpsFcIuA3jen9KiuERLi/ngapstt87X8IkLiEacXPO
RjvMpOgrn1UpcvTtasGVEOh0os5KdHSjFTmrLqFp50dMnDOf9r2h4DRmrJHn
0w8oK6/f8Ua97c8ObFfnHYZugswNWYRi4h04CZz/6/07NJPr+YMNr4YXQ7Yo
603lDhrMh+Yp/WGe2HWiNAR/1DvNrZ7/qPZr3UG1r+4DmjpV9QPlEmo8vMbj
M9LuqtE2sf86MaRA2/rZAi+0yd+v8mSdX3wERyRZhh+tj7QGprgBFAqAWR0v
kBSBuggFukD1gnyrhg7TX3HKHmIg+Q/WcA2YoXsuiJ9oRtl5s2I06GK9MFDu
f6SRZj/mIaSo4s4fglsfKqyo27/wJ1H9bWddoOBxUnY07BwP8zc6kOZpM+sR
umWTLUETzJtyJNI4ETRGFmjVq1Fkq+CDYKNqhUM2b9s7IGOw1ju+XVC6R6a8
T+CZUv7Y0brW1LC/lbmMHi3VS1MPtpYWECi9JP25+BrO7cCJDUMXQ76k1XsW
rNpmnOkGzrrAzpkRyh3/FRp7htPkGwBuuqzAkasAveFrZX88cmMJIva0OgS3
1AiHNaaq2nYWRBri+ireCeB0pIxQg9v1Zanro86GSs4mQmwwhVgLkJIyFF9X
aXR0lwiHAuthbNuP/TeZ4LF5OHbYpcWynRmjB+gUlSYu+jVEjExcVMnhzkOf
03UfXGo6M4VhAuHjBVf+7iiYRJNcywicMNrmY7KHSCNZxt6hSoUJu6t3Cp4R
iIoNoUMmJyH1Si+DHfZaCWx5FLJuLqC97FbNCJOWcPhFpZWgTgAiCTFw2nZF
5f/F837MvKcxriII2nd1D9B+GKKE8J76cjeId1X1kv8amJVsDPcmVz5zF1Ak
yLzYpnRBTuh6qrAC/nGzM23cnJVQ+yxL7ZiDaVKea6UVXpzib1VRVg8WknhB
IY8acO5V31CgBRexrWsZurj+2QGwrwOKv1j5cnJO2GEtIiRbpC+UosIfNCgn
Bsg0e2OZpVbD+dappQPc+vzSTHzQnwUFeYPv+mX5XgM63pcLXgZ3h2o5e0mY
4+rHx2c6YrLrHhclQIeQMDogEaMyTuYsTQqrYolExvD0SMha4zlMR/80Movy
eRzr4vvA9/wr9sGc7ajgUE13wFPFet1kpAq6oXYaESjKSsnA8PWGO6sSk8jo
l36iJAyzc6cCP9YRvBHb+oJs09Q3BNUicDIAQIfUkTtdrw9aS+307hbOEZBu
7fpDRreB7/60YggmyegcmfbX0GHCcSk3WZ3UDg+gimSlVwxxVasFGblwOdyB
loQoOhZTH1ZCpdCzY8+agIyn9rx76F3eTCglj43/77VRSCbpVGYdqRMXFD3s
0YP8Uw0jojm3FmcfpFOMRBalwbMI/L8FJUC1Il/U3T4yOM1H2pbnXAqkFLKi
tB/ZOElSHLBvwiNM/85o7Spxv7o94xxbsXYXwqVUmqnFKRQpz0LNWwCTlGik
PfJ+xD9+4K23K5pffONP2AtzEv4l6d2BdsKAuCvlv3ywerwxxK6A5DkOkBnN
W6RdCqUtybhbVSAcwRK6b1aBdJgKqiZuRGtVZzaZ9tX/HekqLnTxWxcSuLQ4
6+CqMY6vikBidISSodUs2tMGwFEpcrP+ZyfkA1XRJcIVCWWpVc2iUxqf+uQi
4e3YhutkqbeFqVCVLqA8zVQxw4XAJqWrrJWVCbSL5SnladuQfHlDmDEO4mry
VXmRN/uWuSfL/4brWDQLf7zfTxodSnYZWccftT9AhQjFWNFVNOXIPHgZU9Hb
irWIHXaTakyM5Ixjwlk5QyfEXu0y1D8uqBwP0wM+uYh8jdLBRmMO/PCL3LpJ
/obYogh7VrLEzrACDjEJitRu1MHRM1nXiMknM1JC8VnQazffdS6fp/fM0sv3
3l+0oVWA0hU1hXAuv9NrHfF6fkJAUvHosYn1L8u0BnH6uo//btgsdpNlfHoh
xa9hpLxhq3T3pWQ8sAgCkMbzpFGBxvxQzMi6rRoxYOYB+knrYUiXnZjntde2
odIcMYK7GoL4GDgl9B0rODdpUTMGpZwE8PmS22SeIyg0zFzRXmFjGukCJAsG
E3UnHT0apAaIo8UhGVVwboOq3DPWe2DaMoqUTT7E4VJ8aNDG6IrkHhGblpHb
DwN8lb2iLEYl/hSn0oad9rGt/q4R6jTWTPtWwaoxS1FOOwrlqO38o8laoYgL
eeLT5IBONOSpH76E6ykZ0Xw9f7n4v6ZQbO3BepGRb0C2KpM6bnvN7JT2yFHh
QMbOYEzedqdeDy6IZmFZLzL/6PxKcD/0pyU18g87rttqQIBxLXOlzkrVksu0
P8Gv7RPIDENjYE8EQtAeyGIjT6C++bEZAyd3/QNg3y8IlXtptltLbeuY6+0A
31UsQTabRIgoochxD959lv4a0qP0Bp88S+McP/VQzv5dIfD/DXyBnGJk81Y7
BsMAddS2Q4k2ntkxiddEcHDLQMdTIoFOCYa2N0W+PkT/lQoRnLMl4mbjcGfC
195gtFlFTl5TJcJdOdgU2ZEI3C8fCy4gaptQta5+a39tALjxs7tBPxoy+7pF
8jy35W6Tv1XsqUpub9eXZDw8/HWes/LtOzmB/8AwcYwLb+2P+gMR5Ix7b1Zy
g5N2Vx7vc1FQxA/62+eKwHMzwjtpF7pUTwypopCfy7fIiDEvsO6FiikCyDkX
XcNWpA4mtIJAh7fw3gFmKZNyoXkucasQoQzovCeVLHTcxfL7jEg8HrehQsha
GDZFFddp3RyBGcD50GWY9dE3oRIhcrmFfsRsNmirrEwqvbH/XwlGXtFyoMdU
DcdnwsVc4SUC3lro+aSoPfSIywzyq8yOhjsdJOm9MCJJ6Yl+KBsuqrG8T3jd
gOzfif9IErwujUV6P2eq163eK//fVNMhdrWMWMfE4FKZH02eFryRqomP7Pwd
Fyhik9wZYlg6H4YTfLDetAvxKToqpkiRZnfBZpU6K541zLW1f37qqs4lyPaO
J5qxawIRkMSsARZGwbA6+lrsdFXoNP/HMV1KyQkpJ/0iNkAOB9uRyP3eHUjb
MaRweGqyI3qhBt9B/LFiq/yHUjuIR+s3DIquOIpkNFLFiRBT0AGgHOPO6sFx
oxz+HVP5wbiywHzIVHCvDrBfCIjukSGLI/oJe7+X8NxgNBNPyJDRWfTszPTv
InyO34eBBFHZxAHNpCLQ4D5JuS+4LGQeDksZnpXV7iOFYM0MJcOK0xeMcY9w
Ea6EahL27Subro05gaONYdWLhLhcXSI0hoywSusWgyX0P5UtePtWUPqQXX0r
aPDUWaRLE9AdVdI+UKxY1EQKOuJwAWgHhQM0Pg1Y9lB94fRRQkGPqotMCF7g
stCvod4l2tyHbKbjgiMvwgbLoExd3WxUdnu30GPv3f7o9NFXV4XO0B3yytqe
hOuY+kCY0MFYp4A0jWDsv+bIOVesa74F/gT/6koZg+xFrsEV07PJZxcjN4ec
S9aDatDr5V4o4HAY6Rv+L1wlTPaAKT+h62cZFN2jkPEP6pAqQIekC8gzeGLJ
t0ZdLRjQJKlzKNuo5SAZzoUSy9Z5PmmFFCN2Bay/kCdmJZ2c21cTC+JdEMdY
cVQwV+ecmTgZv8z/aHNmpmoRrn0RiuN71u19aa1by5Qn04BPD+YyWNZmsJ3y
mrZ0DBENDDpqzDsUwbVQZubBh7SDjvQhs0pwVNmVK1nVJtEgJqCAZoLdMwGr
R+xr0RbxPi7ZFoYMlF8DqzeCWkrUy7T8hv2X9eVO4T38YiDZRRO4FV6+vT/A
GktFwS2hja7XgWJLtbIEF5fmQV5Khc5gPVt/BODy9qcnFvIzS53fSjG2LzKY
512kkpYNEQhhDLcKGY+pICdl04kpQOyTlw2VWhtrnYbTqAg2FAiZzcLagPlI
2qWsNztEUqBTha62a5ZE+lbMxSq//gmBWa/01wuGk+WWqx5UA18wLAq+w6a1
s0leETDADR0rRj5XLj8NoNoYUCMQlmkYiDA+a3Lg4yYJfdAXZ1H0fFujnRwT
I9JyoinK/hIkXdlrg/3/f9BYLOAazQrXjRKFA/T3eRRVAr0u+/YNUxYxIeda
xrUzk2mjOdg9xLxPrTs0J6g9sjGCR2HLc536ORIGA5U7ukibaIsmlSg4e+a2
qUz7ISpI9VJAcmUsqETqpyeePRNcPNcQEIQ3AF4pCM8xoH/DVy+lFtw2dZ5i
bSyP3tuFq0goSH6KzwfKTAnBKE8R2foTJZdhBsNjX/8WqnfE8v/WawihRJAt
FnIl0fWsfF02GbIPvhTqMdnJsjg/u5SfdPwTIOZ3mkLqftt6f3mKmLcYn8j7
KJedH/p2a0xJJfpx26zJwlcGfMofLaxmB9dBi6SQpP//go/0lPLkgCuktFJ6
AC69le38ORslnspymg6K1raijkrH57hn2cEieOzcbe5b8FpoIZ9zWymMepSS
54poAICSH4YiXFcQtLrK4CIdu8UzJGhFVbGIKJoTht8D65LaW3l4E08s6UAX
Yy38ymyamFWwI4nCeH46KTh3Hqy20uJ+nB8YmkZ+JJqlHD0KIQ4934SVlYuX
6Za+Q8Z7usD9d4N8x2vaLqzyqVNtvPyFUKmBCJNx0qC7I6fY3P3Loy1Focpc
i+h2X2DWsZiaOvoyLzo3hpHJ/tqXC13ISSGNpdnYOZ3MtT1KsFGF4LBxuc+7
ZybREUKRgjhb5cHQi/fAhfDVLPeh6S0EcdQU3iuY8JDrV+oJ/jpS3uBthPM1
raK6MATgJN3BdYCqHH8JfgT0ClUo737GVclkgmCLphXw7sGDlBebT3fGcTTr
KtMFf709dLRhiPcE4UjtwR6yD5PcSTJp6Q/RyuycgkOpIhpyKv7zPMROsfAY
0375Zh+APcWQ4ypd51Etgp18PTDGgfibVmdRzwKXbk2HEkEwARJNBChlwCTg
4Ns+m37I4ZHwYNFFSD9ykiWnps5+qntMH3WioSNTc/PnlSRb1dS+RDvrGRY3
oIukjE5dybLtUdNVmZDJja3hplOSMOiyC8Vgh1d/mBUFREEWzRV2Wq3mC81s
DnM+i+XJOKzo4ZmTAFGXWwnTDMIsM8QM9dfS+fVuRqYifd6iN9uljVZgOLIz
r2HjQyWv43Yb4lk4aKAd9dovAfpnQe1bnTvqFlTQZk3aIy4z2rYTmi1jKuSA
y04TgzYZBcpEqArjv8RmVrCtiCN+HPKcRVHmdBuVTKSXOUdDgUxh3MODqeUb
lLkN+gm/e4PAXgnUSi9/C/iVJBFyQi5waVB4DU1hP9Nbwv4iMja4R7K5rTKU
e6QKk48VJ5CrEVxvA0C7zT56ztiB2LmnWmxI2rOwZLo+e3BNab6xCRnE51+i
z80E71hZo0noFDql35MzXTT6ZgMoAtUiYTkPk50OafAWUv5LqQHh6ZE+llyu
Mmd22L85cjKsgs6kGQUhzhH/YpxvzjgN507hNwSRTn39dbGrN1xwiUPEOiaJ
Wv+ZFwvIB8SiWvWN9OjS3XG04TgFqtuRQo643MWPlR37WvawvkSk2+qOZL7I
iXC8tqSVnYaO4ub7zCLmQobJLe4odUbch1y9TXQaHJnNuLW5H8sTRaDCYyc4
d9MYLCbERhSwXglm7q9Z6PvcoZLhUwREXbKgJBwFZ0N30zBTzz89/Yfnd7QP
mDo6tU6wdQlPGc/unrv3hER8UOmaZOI8iS/QfjCRDUo7SZ7wb2fNxCONuET+
NnmNAvFkB28bCQQr2x8wwC1FZ/v4NYQMjAOsB6Aj2EoKGgWLzpMp2W+c3IE+
Vso8hVcmzlaY8Jr61pryLBr+QzUYocCcflYFkkOSueWWjSY84M2/42cQKwL1
L4wk+8Zr4zbCdi8cyAsUlp5YpmDXZ+wPr2dtxufjGef7bG8bc4mvSJrof3+0
UJtfL32N9FgzYRSS1oO/3oTb9PoAZDMJEGkhiXZiUCvyZ7jHFo9CTDeg3HMD
QDwP2ZAi/BnJT1kbnESsGLPm2KQBtoFTGTJHKWLaweSSidJYA/umbWPL65Iw
7qY0cwfnu5eYJWnrAUp6xSNxt9a5KkBOpvxWQrIK9PmgGc1gEWEoE9cq7TTu
Nl9D3FNhphiQFpFVYVXD1jI5umHYi5WLrh6/akE42DwUEwpd2TX4FUK0J91Q
CeBwl9N6iWgP3IARGecDi1viSQl0cPSuz1w9xe+cz0xXbUMcOGbvLhahD2TJ
T/3TU3j6cTZrlxn5n6nsUTcXrQKxtL11Vpcqdl4bUc+lRgupUFvbQOhZZcj9
bIpC5YMNJ2gR4nPj8oYQNIFNIvmnH4ddNWZ95HR3XJGdE9YYjsDCv2K9ysei
whNuPwOMbY3zVgVrmltyc+U1S08jllhTRXt3xdvjKa1YWBu+nKSQCsZX+pZ0
nGIh2kwhIpq0FmYP6JwLa1d4HMVZ+LSKPEuIl4LGyhuKwu5/wFoZaS3c/JQR
azjqW8aRcnt47Ui7pZOp3lY6kWXLTNb1gCFuLFO7IrClDSBAYQr4HGD7yPqN
AvIbNJfXpzHtBbSp7iVyZ80Gabjhos6g7MaKva5kF4zBqQWx7bh2idVUoOiD
NDhQjYF5rDvbA4oizhrA6y8df6tebO/QFYPY9hEFrO53CnkV3c2SnUZc4eAN
md5MgB69EbN/gM64v7QuqDXlCaxFixyUzR+86rG4Mqu3SdbFPiy5xjVn7uwp
55Ar/7qnYDfqdzTsbLh2wF5h3MPgoJ3Ztd04z5iO1rwxpmkR3C0d6MaQkSLc
vdyiZf5L/G7mpnUKClpG7ZppBZhApQM/+Vh/GsVGM6vlP8joRGU7DR8NpVUW
IPKvMsMoEA1ZFPfj+xLsCbV07TttxtA50es7C78f3qt3KTN/fucLOJcEn4qu
qA1dO08q/37P7hXqsmUF4Gd8BVdYmeoHauAXn4QPHVbHKVTAwFB7ar5qa8Hw
mImYCs+8J3Tl7RZqFiAghzCNoVDng3Yrnnd4MqY3pw9GAXMNLSFs0QkMojgX
nzc2d9WjPoi9rTs79uLh0SYAGqFf7U7Ac7VOL3JMDgd1okMndbZ+esbQuWAz
FT+MKHYEHYE3MBusiqRcIuiC7qVMbgpe05zdglW2mH7fVD5OzdOVsVs8/jjr
Em0SRlh1BZuBccthlVuWMjAeVB5kMwIu1KGoudIQBHaHeKD1tdTuVW0lBJIf
/qDENecC3biKaBDRwjU/OLBEeWGWY1DGHyzLj8dHhWxD5GtvJbimss5eCOou
CAmob6dfpaLd2P0fTCQFDD5wt8sFhZIHhrGl20bHBKJVRAJFUygkUe6be/2h
/ZzossgzLY0sKdUEOzAnkaooapRvJKm0UmNwNLXe52XGM6n6ZmMazOSPoX3p
7T7O5zUapwHUvCXW8yKwKXvANKOz9ticJd6Ew2O92Cmcy8E08gRtFowbPzrc
RdvK+zqbWLcmEqUL+p5BxbyKucxWgAKIYWHjRsMn1uxEIFOs+AZd0XOvIV5s
Gpdxn/1KAOnIUjnp+IQE3A/8tOPxDDGQvp9qO1SWp6l7xcwGU3MjiHhun8uI
BeWObfiQ67GF+uXSV0bRptUkRtAWtlusQQv/6LyZZFIQpGvJ4XzPnQFLYwqf
0/DD9D96xqiFMRySoySCaajln5goh2B1lQEWVPU/Ud2PorzL3pXC8wImQbD0
Z1pR3TITZ30KkedTglrJMJ4MlDBeqB4FtS/vZ8C3Wv+/HSBxrxCLI0mZ29LT
rXRBiAOoehZm4gjzCPOs65O0Tnxrv660BpG3uHvUasdScFBiGSs5Ia92VWH+
aqk/lMmF30mk+Mr7MUO8jSDAX4TINLkmbsH9Y0gmbb2l6i7ZLrUsHPH+4N3c
LK3BXJBKVY4q65m67EknjZcLo5EyYTcv/XjXT8nIVq1OUaWR9SKyTPAGGs6/
Yl0WJaJ3VBNRMnOk1t2zjO6jvQMgFOywJrkTKo9qeJeQRIrKZoDK7yR3liVg
/xMUsLnmMaN8xnpGIRYktal1DFnop5W0MJZDketJqXp/+BIPBE2HMj9V1GMS
Q0rSd8CaAWTMB0e/jXQyllRSL5gHdjaPdIJ1V4ayk4asfQQpxgf1Nt+lfm6c
vkeuGuNQK8BIRgBDoSFRS/PkkaN0eGnfM5tKCgpcU9708aDc4Nhak0elRqmr
dw9qMxqEUHwTjnmWC0Cd1n6/yHWArWDGwNeewoEW73xuwo0ro9Vy0zd8fPMD
Qwm7tgtX2ypsLWopDi19xt88G80VpXmJ2tfJ7EKI6sABoaf/YRXSXKLcW9V8
MRQc9aF7kQZi852DwKSN/U76MePLKwzAgqEzlFc/suQbhvn1rTfL+BYkeT0a
mmySsBBF9ZF2f+BmG0vkVfZ7e6AqlWzi71Qjwt4SDh8jAeEzm7zJE/bSrGiN
9NDCtqjoaMARkF7TOwADu6sDMkOFa7C3Uc0vdKxotjU8IWhb2XBx1c3aWBsq
8V27+96gYCJnIZIVrY6p5uhW7+2Fe6eXt93XAvUDF8ts9LQ3za76zB1mB+rT
gGkEl+EkMHsZ7UAuKnnEIIiO/RJdywn6tPqTTFUFDqPVEF7A66vjH/YuwrsO
M7FgVgq95PiWp7y+ZMZ9etjgcdf3oLrw+MwLTaQwoF2hiZHOykPq638EEsdn
oXTiZN9Az4ytVC7EWbhUQBgUL3bYU4CEGr9gESRaLCXr4u4HMgPAJeKwBss/
cG24DN3llB1lT8a/+rplAHxoL4pEobPLf9tbO2LUq3y/O7kkW9D/wnnsR7pz
yfeUKKQxD5S6R0vDknDsKjdQFSoGCXBzXUYYtQjNjrE/WFrlIQWXvmAfdKNP
fwFu5SvzVX+HFQWiHaJpjgWU37HGFyEyrbMqahPgdIcblvQj7KgfyboNTgEN
d4BkUIeXqLkiA4az/UJhYwwkxLGpppl9/bdIGmi4dLsPjRyQt0RjwQu/iM3P
I7biBRxLDO4slXZsCvBuDJ6I5AfMLlvc8rlzYJy1H/P/TtY6W6X6P6NXiTk8
uvymUZeWINPxx2+iI39EOrWsnFimzv6uMQQHAuhsuU5iMnLX8NmZYK947MlY
3nk+KUDBq8gNnlYSLitQ+nob7YvbdOEfDi9COHpiBjzZZZNuQd9qsb47JJNp
hy3Gkm9AzHJVVF2iUGaNwNOP1iGT10FRzi7E3P4IPlpqr0dY+KtEYKT+j44X
ZLs/0G+aK0aIGY6gsHZYDO5SxSv0kQviNxPnjrWE5I378v3WAyaHHVt4ndzV
s+ub4W1hyQz/BvlzjPeXu+f4Tf7RywJ2EAMp9f5nuiQl+/e/ANqXhQl5SJjH
CLrUgDsr9c7QUa2VzIt09LjOdVUO39T1uC3EWGEMsz/OeI+N+Bjp61WmhMUz
WcvdFkIlLknVZcm9BA84B3mLCJ9WnnCTzNNByk6v0IApaww1lD8T4is3eH/H
e6QyR/CbJYXSHaEM1VEerSTg/HH9VSz+jFGTkt/KKIZ/WUgnnHzGlbbIRVKr
+5pi6U2kXSu1N1KERiztSTS5oyxUtQkz+yNR2nFmwTSlXW5JpBvtWCry52jK
B0BiKz37sH+ND2ZT9SkJkGRBxsMDzhJNIZneUyfVWoiiKiQLJcQGQudx6ppr
BsifEtkU7GKAOqPM9GF7KQQfkynpvLumCul33ZO6ENffQzG/P0TNo/9lrM5e
+Mi7qW1GoO/mpULzsk323gYpFhwgrfjvpaIBUUPi2sXCRodzTrGl8vi0uANP
nNb87WAode4ofVO4D7XTuzpmQEs7+8+JjjXZZ6jLU+EkwEVjavcVeNznv6KR
5f7ABIYWYalASdJ19oeyYs7dradH+KYfr0M8VPgYe+gp6//WqrniwGry7rew
p5PX5/Sa9N23Rdvbc+slF6GCSnAUyI6iAXA1zZSHDlW86Kjh9BCQQYW4uXRf
BTbZtW/KhCnCwsws4B/2EXmeq+2Fvz5hZG8EeIXYyEQ9zvmEQOVSg6iaVUfW
UAe/fz+/BApn0xR38btRC3PH4H3h3OOeWbam/fMSKriVsWMgdTcNpxWzqEFn
HkmI7XzSGcilhJsBM3/Zk4W/ZHBPEpO28cR8toxD9BlMxp/YQnaGn9jzFHIq
K8LhfSMc+q4ARor/VVtp7hPQjCbUoAx3FoTiCwSZwVXjkk6HP7hqgDe0DHHW
R3iuZ+w82l20kSTQIPmvTVOIfZuuI0dV9EzxeDHaDo1wbKTe9BBdkRURgV+g
6bxgo3+kpbkTQwm+8DshBxh6Yiqj0WQkYGDPW0ahx7kFuQ1aTapTh55R2R+r
61k+kW9Jb8oqEdyRnikOPBQxQQfulBJZEohTLO5WAjxHobFh4XKHjgiPA8X3
nVK7Qs0bUcikftYDJdYgXVyKo1aiIfc31aJgO3CKijPty3bBr9VPP2/l0DKx
cxfra6ZnWGpzokROc5NySq9K9+e+Fesk4/iMB+pOQuqQjGZg4kRmKpDZKsjj
bYIEXL5125f/iMxcaib1EEIscTme1a5pCxjWLmYSaEzBN7b7e3ftKr7XBP8x
u9BoYP7ZhPowpeKdY7G91swDbIPee1PSCKKEPigK4i3ZFqr77c3AnfTsZavz
l3hkvidY7rh2tXG1vfaUfmxwhBftDdHYCtOK0hCL74WeWQwDp6ADzKqn4OvF
JJ8FMsvqPOkijE2EPIr80aqtol5Xn8tsdUxy2BpvoDhyps2/VaRlApFmrb9X
KGzoO7KFi7+jI3oJ08bnYmjYZ+QbFlo7t51aRmqYROfX3teNp1fA/GxnT/5C
3tAi+Ok4Tci8VkWgAkkPtyGZq0/TJ2LUocWuNc6lXVDfjNdtdnw+s2CqohzE
u+MsLkVD2RdXzaMO89ADiJLCRokro/0v9GCfHVXwAD2V8aD1GI+cKPdZtENz
3E0lyhqcZ5XbGYQS07fIp8QG+dC+frIxNX5Wdq4R92svoO4SQzU1yqBuzv98
lSvpCgfMqrh0jgysQfJnJBQnbEAVgxnd6U3WBcKr0quWUqF6xoMqXCooPVcd
+5sj/O7tN2v4TMWGwe3zVtxYke6cxDrxwLUGoiwM7YrK5qLNXDaaKgCG8qvk
NEyDLdjvNpnJsbmXSW+BvOnKkc/VIWDOOtazTl/F+zqwoY7o/X5VF4H4zNwV
tjPFjqKchim3ZuyqNIqVb4L8+MRT4zgsNPIfyOD6cIyzPPc9Rl7tm3uz0BpO
jpRpIqIPNA/TX3zfWWrJaF+JX0fQSZo2nYv+r4hzDALLl/igYnq6TI35KxGF
pChIa3c523PcmM1PDvFSxxhd5OTTpqE5z84ORI8P1D+dOpj6n9K9D2F3uh8X
luYJRfgH6+dl+Grf0ILcTx7nRjIHUDN5wFE2sbMRRUbNtWhbt2ZyP6/7/hz8
ew85incueR9gv85QY73iB/o9HNNtQMik2YC//fiCoQr/GkwwK4/OQ4ARC/G7
ova4ULgbvDY322uMb73TwxCfJkkTkw4bOlmr910ugGFqo/J7QEyJ8pfSylxK
lb75qlzYr8Pqnfqi3CW9wLqKt/LxDKRgKPec2HgutS9NU7P6d35VPH8QeMYV
o3XIqtDdEmahCPUDSh3SyRePoTRS3RjOOwIJspY8E5jGmrTdTv2jIxydvkNo
jMLQb+qpZejfz2oHrXOUriiysiZ0loxuC0gSmb1RSwt2xPo0FBsKVuIPEAH5
eakDJFFPYlgKMQFESHb9sanfaZPqmq57zCMf9QMY0Skj/y4NRRZgiV5oyvCs
YCZqidyox6AjNehsGhxHgGsuH4DOS+aDfPGGS9TmB2MayYWN5bVukkYGfITD
//rkfdwxnx8UZDTuQr5ce9j8wYk6I/3mD2/LWfnMkUfdhygGrcFVXebKRCQ+
JmN2z/KHZWN/juEWswjNjmHaa7luJWD1gkrS+zIrBojyYhZaZLJy3QzUk3Eg
tK8vW435+KLF6CbtoD4S+kRhfiACgRALFWCFSrOphFvr/uVG2YNc4uc4Gbo2
tutwNfLtNpjPzcJJPbDUrQq6TN9P+GoJykJRDn3hchOZJtEyPh00QNtIDHSa
F4W+V8fT0+LB6DyMv+WW7Ao03a5+AuvANslPc4Xe0QN1V2pME/mQtqLO37RG
qlxmvBpNQF05nHpfOtHCp3WILyuzRKmOlIV6c/q4gMm51rBxEFBg2smmiuJq
mBa6a9Ikr/K2hUQvTTDrjaRHqKQQCCqdfh8xhOha7MNcp0SNc2RLUe7UOXRe
Pvxe4SAslQk+UPh+5D5cQ5YMMMldU11CGvTYIj3lFFLsMNKbJUDnKYNQ5n7K
oxqAOufJ9+YRbP1eO4i7rWRe8gyFegeQxRx5ZOATOxSI3LMLQLJh1XbvBq7v
KVG0Fvl9sORj1KiUpAtvaMTXsbva4WsHO3nbaJ1B53VTII+YSQtpn/vCVxIv
ZIqumyFnyi4U1g2BaZVExXG+6cL6AuH4ikqA8LSx5Q/HKRI8QDVKgoX6K/eG
h4E0STSTJnfy+IWV/XQnAVHVfCsvSTDMsnk0s5LTJAxHtUyo8S1UNupDMhNg
Q70MEbhxIEJftKL2E6afPhQiEaAMihFV4hTG+X/yNOWnQk0ZTuosGvpyvTFl
GzlLBd6sIWxn/YzGYxKuTLdmUpb7EdST1uAhYTc5O37I6DeB87fNFuIpCrP+
a5sy8z59Fqr/UUE51dnBBGg6gK49RD03vG7z76PdeRt/4EZKrXLJKX48luqY
STyvZBNeG7TvFKdO7Gl2/q9c10+OyGfkF8CgFqhWKra7pcBTlIsWQecl/TXG
Drgc1dHyoRv5VLZlcc1eQknJugEMrf881PPSGh9+RrxqN/7yLcQo5r1zLbgw
AVQpZfrJUycbAetEkwu509LI9GsQtUWFODR+B3Z3Ydf/CAtstull0WFgkLw9
xOcg61X8c2pljsl0C0YuDCYGzD++hjhNQNwGO3DKpNTMj9yfhRr7ZAKfxLLd
h5SWIJ8TfMKm2RLd4az0Y3Qj5PAnX3/IuJ2+9wVIucHzCUXMIr9M3CO5oakc
CwOYerPLxyIOntX5TNICP8CNxxdDqNh/zsEySo2d5F7N5eoA60S3fpGeE80a
efqakWgB8ibQIzszWEGQi4WK9uvvbHUpLrB1DHXqpjhTTveQqrffNPySHCKr
8Dv4KUBNUGBg44RGm2blfrAmyOUH1Jm/AxEk5AAhKyM+uK3s64hT3AKstDmA
VHvNp752+DUK8ChPv4Nvy/qMd10S2sBrGzQ8MQVf7qCvNPFtmgETEpsgKo+e
rJrqmW4fzYYJTeROYpFcIW+bCrXnYXa7Tg0BgGXich0QO8+xKJjx/iexUpQ/
Z3SsCtvPPDiQzqpe7w/+/8KIioOBolZsKTDZSYELnVkLkyW1SQRo4I+5fYOp
UOXp2+rocscTCYIFT/thISA0VQ9fW9LfVdYqdtRLCLhw3HXTte5VQYPIaWQj
yWrMZnzTghQOyzKTWn5v2wKBVefaNi7CnGkHSI9yXYZagW5RTICW5ruK0d3l
ZMDJk5slFJW4qoAle45ny43etDgzdLKRsn8CN1KTMi0OykzsZxOty8lywrmF
aUxnKtu/jZ2r/DAD8Z0sn8AIK+8oEOfTjjUN7eLw2/XQnmOWQgzf/UiggmhO
QOj1Xajp3X8F5Kvp0Go3wN7mwZONZd/8pYf5RYGWfW+vH/d5MW6JxpQBzlpu
IWhAn9126BPmqHKVBVGQNCDLn0pqtVJDaYi6NV1MUefZ1bw2VwGZyn3C2XiZ
6OkPQtG/PUrw1osZfbLrbkTU9vbBO8NL9Nvk35eimIwTVN/jSLegnMAvFvt6
StoEnFoe0pa84vTN3XGdd326KC5YlvDYNRvYw5JAh2DjZu/ZHSt1tqgteMeR
eOsTNzedibkNvPmZK92ilWfLq/mshaU6gBd2GUwP6pjOsCIHza8G+rPtD000
dFdxQHlG07+EOLlvfcf/UZB6P0Fa7xdfGNAnqOOTEaP3qy86+6nYZ3wg19iv
8jaacEYZYRLNP1FsuMauO6M5CEzDPWWrhBHjgELOkjaxCY0oj/LIkFvwEllS
kPWIICghfSowOkEQZmv4MKElK22LrV8Yjapa8GmuqCub8IRBRXwUP18qVUoi
i2iib9iHuPhlR/v14mXGsLyCmCh5bIyft93hObvvuqjybgkCpEJmPBEeGcxp
gXzzh5tkhXS/4LMxYZWLr55qkGd85lRKdcEX3r/X0lLR5VvE0o3dDmtFVH8B
ba0V0SHunz+Q31xmz+qT0MpRQF2znOi8+UvPUs6wwzjLyvSi63JFGUFhaKiz
ntrY7dC6pgH5I0xqQceTdZD4sRmPL25YDgPWmDqGY461/TwQbhK+a8Krh4F7
qvKWvNIxsy5iMR6URcz5xFKhyIAd6/5E1acYIOzl+X3o79CxylFWKkzJq/r4
tAoFeIAzsuuAv1gh1M0z1O+7BcoiwF8Xl+goR8+kueMP+CwB5sDEISJbhdu4
y6xkbRH4Nc+DszwSnRC/eKcHtKBbiJRuogvSfHPfPRd5kBfcF3pW8Q5Fy4Go
1hdb9uDETI2Ia+qK7gP3qKk8Y1ow9yLX18IQ6rsWS5tkryynPAvq1EmpILid
v6DNsqkr3fuFTsKPXkKGx1g+2PyAOeTXh1WyDgfayc5J3KYAoAvnTUy5uzz7
c1a9q501/pXy6AC5+nEq7iMB9dVvv+PPYlvDRl6m/5G5c1AFGI38XnY95NrW
S/aN4p6pw4W3+sAVlZND0ozV4OiHHbUv/MOc5VO3VxELnn6Wb2M29n7ek/x9
BZXn1skFpVt1z01pCvcJMRXdQ2sv3RwAx7XFm2mg8PCQ0PjouuG6cZbfrSoi
EznVSkW8NI93GzGPC2uS5e1TOYHOr+9+0w1XfOV7hp+BrLyphGRtOoP0nq2l
Ox8dqeTP4hPtaxhwauA4VVIOXE1rv2kc92jlDR7zZQViCc95gd8TKmKS/Grb
oeSV+dxSC1VE0zsRy80Auk2FJSs+OHZGvv0+aiSNNWc9cx71DTE9NZihKLpJ
FlgiedNueUbnoH5Zd/h/PWCxOOImp2glehtteDfPbZZvYynqIikcWCCPiITn
pAL/ieQjpaCBWo1StL+0m4TkW0ld2UTdAq29TXM5cTc3gBfLX4lDfbpk12b2
DQyvvIlY3xJ3L6t3gdwtQ5f4340DO31xbk/cMji1I3dncwqWujGi7w/Qi0Qe
KnVJwMCkjfWB4JQNPjRu0dVwVNk9us/0mOSuCBHNj0M1v5OUk4mdzRj3wF0/
A70tW8q/ouQuBff/7BQxDUIeAfPFVqqS1eQgJOMqBKzkid6nD/1MWDvb95+p
LJHPn2VRTsv+w+oxdP/SOuOPOxtdjM+hp1bhbihLMxt+wQ7hR0gw4U0sCHqi
/hktyjTissVLWuyk8dKUxXXSxiGhQAMqdDV2A1wRqbyDGwMIns54cSsxyKQH
NEiLrW/eMCF8ZZTwYRw3WyJQFIo9vpKV1rw3c95y/08JyFXTKHJzmMuwYuE1
5FYgWmTbdYm6Qc7BHdWhkbOs8+RQoBA2FdleKR7mWnVeS0aM5NylKJeCPQa4
KsT7Q/0vInxSKQu6/N2bliOadaJZt5U7COkKzr1FHSUdgWNRF/puovVxcebS
OPmWpg8twKKvpJihQcA5d26BV7mkx9Ls36vfzBFVFIyPsj+CjqZF36Z5oQb/
zbDI7IfmWZItRyyqzxqvl4hMSwnklJ6RcvTIqojD6LBljfUPeAvyyvq1rW25
HKOnKTbOheDIrefme7rBb83JTKgE5JIexNQ+uz044cVhrOi9BywlEHWsZ9rN
LlAZcM9ZGeCebxwMIyS/O4fnabygOTmHR9Sa38vVnCUo1km2KmsEg7FT9eyF
dCpD89szjuLF+hPchoSEbRMj16hw/9kg5siQgCU43/+8xcyEqQCtzIYA7QPo
VRZ1N3L6D8iJiAdLX2ymCRQSVfWm0wDaI0EtuoMQB9biGOBIlL/kv44Q6BSd
9jsk/D3fCYLdsdDx/OApCb7AT3H48CHBL9kAcOnzFd21002BpiLmNgZwFN85
HFYwx3IVCuN5UKbMcTZugO6+Lyry0NgPdxfbPgSwpHrrXU0+SzJjJ6v3yTXp
jTN5COgd4lX/Un81lkCMiBLXbq9o1zETO43ufTS1kvRLt3gevreOPMdvaDeL
wHqCRJf4iy719UtdibOxyONlChE61mTcAHwYEqP2UU1cYfrSQl5qeJuy12aB
UN4bmum5zabCLdK5SpygxnzDwxjjB9P83GCpAp6e0P4mAlL1LCs4vakdfSN8
yqMTI/pJ4FWaASeUqdtDGeufZEYenUrhB3AQZFjpjKh5YxiYkHuS6Aumk6Vo
XPhbdKDc5KMD0F6CWrVw2/3DEcpa/KX6U37QHyby7IC7zWlxpBxqmAYoE9Ey
Q6xDMfL6NZLCbJiR3b/uL+rbzfGgtE8ZNyffNjzxUAoRfXFcxnGlVN5TNjXK
K6TZpyHERatXV72lz/H15fYbamJlHu1Sd3BBluwfM966iOL4sz4KK79eL4/P
7KiobUFezsSlO7UFjrMQVCFTSjJv+c2AZ/rt9M4CP4gpNfTcj/WPMbT3c9sh
1vXhh4VKoMbElFeS+bcOYUf5SjNI7ewi4I0X3LxLrSL456Mvcw/lVRKwSGHo
b3YuBBlDs3rIBUd4a9CbJzsT0Rk7vmcc59d5D+0N/SqktlJ0+fYoHDFwGaWC
UiagfDiHITKyZeCmzEBn4gmG5NCdf9RNuJ8YcZQneT6xvcbmDzqDx8TJ7Xfa
2nsUoaWkuitXSoj8jZFNMrXyGyYaKNne2RK8GYGXhFTgvLefJDzpe8YbctiF
eGF24e9EnjwCq+/JlKMsb+S1Vp6I54joJ6+Ggt6ko0eCIA9nfwwy1/DkC76Z
WOQdeCpBxJEi1H06j5Jb8iOl980FulVAA0yt+v7JL374R+K3Yo8iRw0OOYXR
irxHbr7Mkx7U+TI6zejpUv+4mRA2voenn7ayVBzNL1LLUr46pbA43TsaangE
EiLJVFBIRUOPNyZcgex907uITyt81Llz878y7ZsGLLILGo/gXB52Dw7tnqrz
c2p6emNOqLrVTLwEqJjmtH0coM/ZpUHWbAepYoaZ6rUHCYtrIaAmoHtV7CFd
M1oWHGIHvLlkY4YDnsIFJq9raYBAJL/RW3UritVrX5xN2J2lQpGlZTZkKaq+
tJ+PEnuWPId5Lk09i/nFVPqZ7+u4au7lDuJXRZJnLpssL8c6PuJel6KV7X+L
iD1EKzDPzMIZwGSfHtUFye1AaG2f48WALJlk9xiJMEYOsz/XE24mRr6bVebZ
q2AWtpICmXXitCeSy5zpgJ9LAHtW7u7Jxi3h9l4zHc095XHFFheQmMctR5sR
NukyKVpJKC/KskLnKohhSUuJShlW0gxUx5U3W+Ct6HSaSAh7avSQ7uKihAIJ
oz5UcU+gayuiPeMI0c7+Mx41VFQdCDOi1YNhNqGrl18Y8x5Q/p1GqVRdb03g
sYo3P7SJBmMz07F15Kh8rQzVZu70Std5pzMQQxWZOgAurdsnW7vp2qoV9hNG
2LA7P8iiu18gR/JWKHZcJfxCZGPbjxqWbDlugmQlyfYWvUyboWD3F2By98nm
UiBOv44jlK4iR7owkN2kfcxOLYAAZZSUc74jxeK2fyedAxDdSpUz4xqAC9N7
yk4DgouOYjUcv8jRAGLjiywcyRcbzn4Qc5PFmG9A3vLPf44a5OUUtIt6tLSp
2YbImrsxgQYbVu2RXUaLnWGPtT+Ql6jWWMsHObe5VGVx+8+grQiUDtSgUU+g
innfzZG3JGNIFA3Dbot59PK5y3vwVvVXlrskrg+eeSU2c+wNEYqG1m41q24Q
2m8qQ+b41JI271VIJnBmLXNoi7LejKT/7j/7z8cR1nfho9JzXU7iO+aPFiBj
tK4hogL4spb3+CD26vFRU6Q4VPHJfJpP8GDws+jQxX2h2saOadzbG6LXUXrI
dSBLmDetPQUfrViRUb4WehboV9FOHMuftBBYdEe+0ufC/fH+6uE5Zga3x8Ba
qbGnhq3ZR2l/JquJNn9eA5C6+RWKgBaSdxWL7E0ykyq7TIP6OjC1TxkWqoK/
nCym/ecMqzdfXBIzeoiuMDrgGYZ7xVs3fqILeIkzBB0LkjWW5lo9RjwxGHRH
eUQpYglc+4T7CO4UNuy0MiGHjsUwAvqG9NfMrT9fAOpdqZFz3ZekLsBlm35P
KOYidPN2PtGm9A3dvUkMewhAK+neuPGoKfGO2Yky9zZt5pHT73knjVSoc2AY
epfNfUnhe0OTjBcMbFT7ChzWV2RlpV5Kq/ZIyEKrN3TPc0NeImhweag9eNLf
SJVTPTu4zpj+a3gEnCeR4dU8MgHui++CJheYJP1eboo7nW6Bj/6OyL7+If4v
VsgmmHm5X5t6j9vKhLWk2NSjioB81p2tM74bqLyGPU0hY8XCq1OvE3c3uBnG
sIXBCJ9OUO4niRrRd3IivCJpoV0WiFtUBE2xDtgBmsLaoNW5L/F4q7DIx9Dy
1CMsSUDtR9GNcoZ7oPole8lbvSuaCYTw+iPS/0JxzHjjM6CAwP9htm38X+7o
c3gvJ9cvxKojZbR9RN56hw09L4qZd8qk18irLSdZZJxvziMKzq0t5I4F5hSU
oCXu59aUJmo3r3wHWKddDjWxQAQ5PWuiwWlGnZwPmUzxlsX1Spi/R+YOKd6D
B3Mf8jgzPG/RnpJ7L2RbFKxo5tCgzvls5bZkZ+QTv+vpITzSDLYjcDWg9S+g
J9B8NefuvosLePMaprsgZKcZJDb5e7GsuOPUIeNpbpk85kkkUjtK4fN2euP0
Cb5dXcVImUyS994v6PBV47SxBhxSd9yo4ayLJTEU7j0wIOu4Q5M6HdzD3GhQ
QHxJPuUJg+wpJiimO5sHv09r4YH82UpVATq/1PpptL9rOSN8G/g74F6xN1fF
vMr+Pv9NKpIuFjfstOSmqGM3UXox5UqyJ7jHcG6mYX7afmH3VXo7jhfrGTpD
o/GVYseVf8Ofo890uy2YeHGf9uuS+gnvsGm6NpfmakUupshSKyJ0p2RxhYTj
kqVvC8e/lJZb0g3b4u2iKNxkjhFzmJgzW4R1s6K3iNXLkqqBscjKTWz4KfDn
fy5H8v4GhY45y+ofPLgVSguuJzC2rlty+5k9VqO6eNv7pqMbslF+Ru+EBxEv
Ko0TVcY8YEF79Rh+3Q3L6qYTXSXsjxQo9R/l83b5azN7/Ap0vKbYZf7jFYRh
WJB7J7eqbjx7TsU3QSF45CAMHvSnaYv00sMJfPJdMFDUZy/EX7r5MS8dX2FI
eSI/9uVG40kZdfPK4qpuK3RjJ43TRAxtlDwpF+D3NDvjOddUo+/eyZw6hE8f
hZ5JvtJ2FnilrfBneZS7gdpxm1d9OptNr2J7vaiwLsJLNHPZZemTvk9FXJFy
t6JOcFcmUGpilyaa7g1+vbOgkDFHwEb2fjZc6x9OB/+L6f/Khgf3ot5mdff/
NMWlYwF1Q3vPuLYkunIekk4X74LIZQUgeKcKYEcRr4uXeDd9eXlsRt5ZN3W9
08VwctFvE6nHNSHPTOmpcjTLgKMuW3vm+jby2njF1w1OA9ViKpTxlDaN1xGm
f5ltvAZcZQP4fEdhc4aN6NjEdqG06vo642KyOVUT17ZVhqAQPVk7S7DWYZtx
otqDHlB3FAPbShqSbuGCKZtrFaErgpWYSpT3ltv6i5Oj/t+eqauXW6afZZ7O
WrVkcsbMNeRo9ceLSrPuCOafi8rdcpHcgqzGUWhvSolmMNWQFFHSf2CPIX73
v7JwAao/YztsNQLL1JzNb0yyTvFX8pHnM3l+JuUAO6+iK4TTKyahDPxJbXPX
EOOk+g2RPLcCnkoJqmASBakwT13rCJCS0Ceh26uJLIsJ4k0QIKVgcC+7RFUo
9t2LGOo9mXlXtTjLUmckKs/7UGJqLF7Z2dZlfBjFjHrmSGYtgbkpb/XI7pov
d9Ej7mSWOVbpVu56SIdpRjM1o/inJqZr8GK0sEl29iSmtbyV9OfbcwuzBlq3
OuewDk/Jo2SMdUHuD7y7yx4ZBSiTcq25lO/S1kslUbZ0rR0CqaZYfXr0Qbpa
S6VoWwbuujTbYRRaLo6Zdu8RlEfHLgSu0mt98fvuYfC6PNBpVq1/EBMO+HkN
h3eIU6gGbajix9adBM/q0yi7TJGp9nRG66fOu0ou/wgerwg4/jgOjPPGcKHs
Wdu/FwnwbZ7Xs6aPPzOTS7RrbQJex3eBVeJ3wVBwdgmQWKkxq+Bhl18tPucB
RzNh9L3PRsDbgF6D21I0c4ZfevV1bnCnzLXyede20YVdvwi0YmXxWC8ltRB1
zs2WYEhAV8FrEjtGs08M7niUnB0hOKr+gZ5rA/pxFWWHp//vGbsgp8NyXNNh
MSM2HKgr8cPKfEE8XOH+HT7GH2P6IwaNP0N9SbGEJSyPnUuqWkkq5LQrdvSH
d2K2wCDcsUJITYsf/qFiUy+n+5h3SO5ctnVEhP6aQjjQtiDYbFyP51TcXsDt
fDyT8z3/i/PpMVPDodvxXaSNmDLePURI54RRmYkG6/+RRiZGlmI6v5ZkZPr/
obBckyMT4tttOt7HxHkKn4VKZlQgbQh/co9thX7NpnOyQ3/gXZXRX4YlKbaI
sYjAWiZTTDYPecpGAGsmADTOJXyQWAdezalGtJYVwYgXmWsOw7e9qoAVnEe2
QVDtNGlo+Z2fD1d/wbQtLgLIBjom7F8fJnVJu7fKyH/+d7/dhbCQlw7T68qX
YVxkun1cgQePy1ViZDzaRYmipYVxc19pONw0scE+MZh8HPw0Fi8wnqO2Ik3V
W0XAXUtAOa76GGCSh5ZarucnBWQQQ4lRisA3Y5rj1I38k5oFHepfH3dqPf7x
D7u0v6BavnbN1T/5jGovXWqTcrceC6IszhLdTP5e4f5YGxNzOa+4O/UbcOVF
4/hIB9ZyihU3wJ+aw8knCTiAf2gQXw7FS4dG+Z8IJZb+8na3of28tsOUcZ/4
slBmQQ3c/sEU0Cdl4vHmiCH0nR/NxcR28fRNhtu+NMzxcUqfD1bOkvnXCpED
T+41ksl/DVeU7L9Tgnqhzezjtzghxusr2bt6g+BnBMsb0+rF5MRq6XbfQxRo
MT/ADIINTgdFKF8ifez803z5PdbVyk8FP9ulSx1ed7Lc0YKYTd7K8qt6k0Jv
u9+WldbPDxqbpBFsMlcXp6brJ0NmVVpXiJmGB0wruch6zjVhTDAjJp9UmU5r
4G+IXHcRckK4RwF/TmFqfywsZbAAGXxIhTxmTXA7aJO39dGuTeYfnZF5/jgt
5auF/6d0ozFPiaa7qg/m5Rc53vqK13i/MpWffZX/52GaXhoAtGBqZZXyvlSV
XZ8b12n0mr5I4kMIQZ0FFDpLrFGFFKhZ5S70eQ7fauEXYS/bydi7/PjtyJuY
bbQqwEZR34aKIZ0MRMvu3ta7BIUeavfuq4zot3FMLEi2LeIKkn9kj4vTDabw
vu92JC83Ajsa6qhIxLhncPzmfMOsSaGl0YvDvDgB08dMK9OvB7PKBZT2KT9q
Els+cvbsKa50XcT6OVgTIF5pBlKTl0UnKvRuFiJlZrAGKNi4ilLNZrc+Ov9Q
R1O3LsmqEY6xy5aEd+1rZtjV4j2zAF+d3p/Q+mGyfQA4pZ0S9zEncWw8dcUu
8wROwpxFKzmp09/D9V91zwg/VIzMGuAOs9cUUJIVSeSpKq+FVQ7T1q6QKQ+S
enomkI2CCyM/yQE8doGKyJEdyAsZ06QSiIynW6aPSxIsUYFhB7QzD1kkAusv
T5tP5JUeMmDXi/DxKcwkS72c4eZQt+b+VtvYzf/t3AKKO80HxPMmp+lEfykK
Z9Rwix3Q2stRNnlo+YdDez3SfHS5HboS/DUA9Xf9MAcOrOwjIGcOqg+gL+QT
d+Nmom0gpyPwV4DTn2PXuHgzzrC/SYm1AYBVOanh2U3FuHBJUkpDlXE3L27c
yKsPwol0m280VGdc6WrK1WBmofZ1bFNFPVkqce9Y3Bwfj063HyVPUXM+CY3D
r250wbKsf2hwC1MClzZ5d0mwJ1Jo+LsjwF4JkLbo0rFBYiT9h4yxSfTCDTZr
dKBUfYmRvyuDDyFRVhXWqRh6M9tkycJtHIEcog2RqQ6PSgDLPQJbPuk5QObF
8zL6idIPpe6VeXz4BfM2pJ3TccJ2JveEo/TeDrHhZKv4kPhvGpIk/+WIxC/v
ouxV+MU4iK2HG75u1fPK6JHxXAy6brpOaIclEnFDuQjGZeEabF0kMUMsRG/m
5SJcXrpmE5uCX3LK0087fv/kF7MKa1HJI42C84xuHC2dqBlGiq551cmaSM/9
BvLE7A+MOVC8/6YnA88TRFFKTK7tHPSO5xfwJuiHNi095FPi+1wSgIkx77OF
NUFO9SFU+qg+IDmKIEmEIZgXAyEalEswzirva+TZbpZdVghTBHpyLMwA3Ut+
7sFj/EV4NXVPgX/zZio6p2J/K40Ob96kD92SCx9GvuLdz5sP5RvwGtcY1R4p
PWw3ZDvIbDs5UK3dggAY+BWZlZ8SXuJDbwaevJbTQB4di1eSFirjmv+fmt/S
z2oDY2Tn2nagtYfTgITmZr1CQ5+wEFqPKLhTxblNZ5nKoZV+r0HqoxO8bZH5
XCaS4i14vUx/QEoacyVC+FYV7eIoTo1sf0sXkGJqJ7r99AHIlB9xWV2C1DLF
Q/QoNj90fzb8+Yj47FwvkAkMGZUn0gyo2ZgcaP7TDEt+2K4xrOgQwWeMODCg
7fJ5QQhBwqUFukFo/bvgjF18aeVaE4nbzYXx/QwSJTFFJHsYrTPgB7Y5GTCL
ahoKZLT059FMMptNjD37IBVWaLbIjnHpYV4loXTuVsYqGdHxXC9fF5xaboh8
MlzKsIgG+SaI3+CSlPtIDXcYzxOh7b3+V021Lhzjbi+ZjuQi8HgjYREDjYbD
GECMmijNs28AJVtoQWMqj8t1Cr2u1eYi+oczwsHupNzINWmUGAs9vbA+U0tM
ChpLPIIgYIBw94Mqi2C1uC2ksDlQe1Zuwtr1s2A6eiRu0Su9pXW+wA6qKXN2
J/m03kPbZYhFnSM5yVjQErnAJ7K4uGVooWiJOdnhbgYhpUHlaxcxT1FXfWxj
taYsXKxO5BxE5WUmn/jTbN1Ish05VkZW/h8adNMrO/Dh4ooiLTELILkezE4C
BDuotg9ZEzEj9XF02awS9BShqhp6whJcuk1vT7zI0QDS2Ay/RKrb0SDVR7S/
yeR9AaoFjz7ldLTKn6JspryK3KO5J44ajQPgw1dc/FW4zLbrKzVUIn3+9cGn
GNCCu2DcE7H7ddiKatOVa5PSonJ0J9X7KeTkOR1+4N8FJJARCq5JiMR9WVWT
hMaAOWCaZ3l3itMP0zHmeO9NOKhY21BLXZavt89EpwGJ/0AL0hxKnylRczjP
bZStFz6W98pJ9EP0qG+B+h7YDBcCLEVHCRFD8BHuc8fu+FaG0LGGaG9rtNlD
0TEJoL+OOX2HFi/V1Ogf+PqjxWKjme+ZCD49C2b81wvICdoR5P1O4uAzNoYV
wScqeIlKOj1Qw6JlXrKAYCMBZlp1SqaBLMMQIcvnuduwv2ROFi2/t/QeoVzL
lYLg7uhhkvHTlwGM225VlQv68iG1/93p3/gJY1OSO8Ij/9W2heMWowOeZi0O
xuuqL1ZNmo6doAF4Ky38UdbPJGaGg0eC5vs96QVqcsX35AEbmZJyCUVcbcFs
qwIx5qki6c3FnUelWAnXLNY/8VEMdNoimcl+exPJ1h1P+KMo4zBsNR/Gau7o
Ov38md2Qpx9aWht7kiBb37TMp/HmyBBWqjXYgnV9/5vUAevtzt9mrQ0vbnGN
Hv+OVrCEunUFuDst65oF+8UKi9vHf40ceCci+rmZ0sBuS84ci50ZEW+AQRoF
iJ3Tla4Nxla0DPwD0dlzYdEJhDp/2ohPNXof/ft38vb9fvuTctlIxlnC7JOU
HNKM0zj0hYgI0tc6N3FhR5Ga38CPHD0xDhxmsaCWVBCGkLloSjePn3gsv7nH
jB75e+bRExOsHjB/OWNUl+zpTR4yZ3HRee/E0otlceAIypnOziqcelyfboev
7Zqq7Cc3sT8QDgve7WEKK0PR90+4noauUdwywpSGUFIXy4TvoJxdRVKQX6R0
utJMIoEQI4R/D7vjy4MMFJr5wN8WvtNqO+5PjP4X6s0U0Mx/xCLnQe1h5i9R
IxrtiF9gVpqIOPqLw/rZgX3uWocyWqPiVgLyZgree9lNUQq8Uv1GwfTTcjZM
/v6ZFKWedktuLuu3+/5wm91SFuaUO58p7jckAVrRxgUE663GYQg5/jSS0CBg
d6SnRCQkeJM7rshKgdVLjWHHmLDpY2kxev0TXNlYycah69GsfXYM+YLq3CNc
0UmqoQOoCwLVPCdFAHpumc9Bo4KJS1+MtCj6FBey4XV7lCHwuklPSjHtdOZD
Xvu8SEST8PqnTIR6RQgK4tVg8QuidH4msFfWN9uypIiMyznrHxcy/XzOkF77
uis7811iuA5m03dgDe8c99GXK8XEfgwfEjP4GkRfn14DokUS1/P9+2IMQM1p
vCXYWqZKerF/NwjWUY/UnpuP+quEAWuhha7Wbj6vXDp+zRCzLLaXobSTCwAi
O87iMytsCEgT92smvxrhU1atnNeo04MjBcICw0zQLzqtPZetB7iKjvYSy0wK
pvY+kR/DXtUyobA4QUWvG06XtpcfgiEBgi2z1GT54LnXbw7/OkwoPIbSuudM
o6tfZ+YLG0zhInVugQGdwtXWpPlCNnCKzSuKaxhxYhFPwaqfMH4AP3nXaCiw
RCsO8pyJ7yys+PYlqhOTpMWuWxBS221B96aFHxgwngJCO/puGSetZMWWStOv
37CLwwttsUrAG/iSkY3JB/B7XwaQZ798A5sC68eyG3UjNE/0606jcRXpk0k6
1vMZ8vlsLoUputVCL+gsEXWOrzyBi6cHre5sNhvoud3zuEYQUI7uxKb7AegD
zvLCzgo2ds7jystrUgqlLNtP+W4f+CmspuQDM6UHasIRoScsarvzi9bki1lY
2jt9K0gRHoElNVX5sbWAL34idtrDk5/xvcOahrBKeVXIaovY6xOBruV6rLp6
t5P17qFoxQb1DA+aZq86sWydJsdi0mFiF+wjX7jWgeoQP6r8k/medFJGSu70
sMv570ihHzMY6crlLe2fSnlbpysd177lOil8SyPlf+VwRNJdgeMILFmuAuI1
rOoQrGc+PLfNE4ac16D/l32GQfkci8fVYfAqSZCGm/K9JFTTP0qhmNvcicEl
LsqsOn04OYaT+NqdFx1OhYUWAvfdHbWJK+CVo+RHZdoNcJqoxoucS3JVdm0I
hCZb6bRmrCZpa74X8Pco2qOxAvnzeLIfQdD3umRr/FtZ6vwxzS4h/e8oi+Kj
Mud53m/Q2/1DHCQZ5xPW8kAcs/50qlcWhPqWD5/CfTgwsm4phXQqCfgUs/Uv
wdHTAVXxL+ZAVAD4NFCCX2/I4rx21wkThlF/Nu+2hYKrImOWAuKyZbbRUnS7
PnoWK3XZ2MRH8tPSy8/Kpu7qpQ/IwodPjyS8+sutctLlx7CxrubRc1IhI84v
rfJtoCESr9Zr0UJao4FMv7YIkMfgQYiE2y0MMcQyKSnG/Q67hknc1VhyVXYF
IUmSSdu+ssh5cmdkx8DC6DVoFS6mx6MnX6f7h9jjlfhJezGORaVV79XRj0r9
YN5VkcekxVlpN/kyGJPI02tzbgXKkgu0Jbpm1dYMy56y9I0eCCnpQyz32pMD
CYq277jJZdX5mdrQWPQ6HjNGQgZpvnhtwi8SaFZWJ8MZik9f2AA8yh3i0jeK
9OZ5/X+kacR7GgmvLDm0qhv2nnrCQ5lb26yPZmRl9R9iMLVILsNP9DSYNakJ
zqTTxmWoC1PITBp8TBJ+NFi9moiwbIN+7TIyRShtZ5SfXlb4BTrz9Lwf/lbm
V6BBFRizhm3X1wRLMDQ/Dt6WliRkVdig8aR93/o6EtEAgpRNNiPjjPXxDmln
GJcFHIVVj5q+U0yAPBkMN/HldjrNfrM+xyHp+AcCPUOVp5MST+A9u4NzrB6I
ZMTqWvBpFBGxwXchM/ZyjC06rC8OYD/Mr0US6/Pu0CCv+9UYO73k39M1kWYF
Zf7if4y6L02xEbUp56LKSZrvnbI3T02a0l52AI9zKgzqKkoSqJ3/ikcCGSiV
u+iJzgYIyacUYcUxVeGHwfzbrFuARrKHetJ5ENmb8wGM7KpvsAStNpLOMrFO
IA1tqkMJYFkw54E7X7FAPbB8tAd0G4usJygW3vFI52zXTBUsffaOtCo9P3Ux
kYWZqRmA621+v43InKZqfOOAJiwWQrhWOZUGcKEAcceYp2Gbahw663wdwFCF
9uAEPauKvRww0hbMbFuPo9LnZNnGPRX75vjwi6yxelARbWd+x6UIIJWsW2o3
n/t5i7DnlMlOve3lnjwSXM5OyLo8cGsLbxtTNGhQP7KMZeBFjY7dUmTwxyPw
Fa7WdGR34En6fsjG5Zucj22HM2bI9HvUrx6rALGY9erH+WLOrUtUDJmlqgCE
kT6JKfXUyrkru1ctz/mbeYqiS5B/bcf7+/Uw+K6N9bBqm/PvZWcxmsB7nuWx
FeKMBC7bjp4RG2UREE4t0lu0G1A/7yjxclxmG/5xmhHoyx6M1maGednLs+b8
miGiS+btyOQd2uMjaV9RELr4Ik1x5p/MnttJDzrwnu6ztw9OMueLFjqE1T3i
x1HegvsfpaxPI4MbFRKyuGKVUG6xut4ZSsXTPVgj883aFyrCroS453tSZSkU
YXIBvjYjbNf0tmCzd9ppaEoOjpjpnxzTwnaWrI/rZVssjy1YyvlBuraT5oAH
i9ZY8bG/bMDD7VDVDxY7qkukNQlh7vzHMvpKtz5smhMQRoFMgCYcRp9jCnOG
iRghFItBTjpurYkX+k5RqGmZUP9G1kywqVnvL9Bh7R63i40TsSlJCBcDjJqS
dHRHJp4IHy3WEhDFdnC4g8MTrix2ItxVp3cXt+nhYNUrIhb94E0LY4L3aFAU
qljo6yaLXhw7A5o9ab7pUTjypt6jjiV0qIRlddZXqNla8sMbiEiWSbB1nH5a
dqA0hB/9jtoeNZj6pTPb29a2WdWLXZrgW1MK8V9TOodbOHVtISxrtHj664ty
IUtbhwlitkHx9Kc7h92IOaI4+lW8XX9GHJKl4GZbzIyo01JR923yPFc7nQWN
HZmoAdyuy2flS+usUxkyiYLlekhLjli6gIRDEABLboLDyQoE6opWMICMi8cz
6MGbIRIXB5qNgA1sTA3PggKQ+5/XpYsR7GnP2MwFAWd6PO6TzRNUA9sdpzkF
8yanKM6zZhkys+Way4U8SjKLlTQkbIIwBf0ErSM+BXUVeTUWqz3JrY+ps7KM
FLh/X4C2BVrzmK591K1VAtPPP/Av9RYKDQ90yO2DMv6f4Q8FtLRRmnDSDbsS
SC4JH9We6aEjgBI23FwGZhfM/ACkpBqqjZxlOjJjSb5IZQytWpflo7L9aEat
Nm3Q31NTj30OBFx4HNl/psx+K5vvHe3O0xDlAP2ldH0TaiFN51SamYqni8Au
5EYB3ggaBimifS6yJu+0KF6SKwv6G0S41z2EGKln1gvz9cvhDKmFJVRTRpOF
xx6/gf1okmmbDe2NuIVYjEOb3VQh2zQ1OIFZ2UwfuUtnPdaNT1Eu/DQ648Rj
XycwY4L+8+7fvJWJLkSVwY8wfS6Qz/0j3q8RmKFrCJ1Zn+SrsPyMMkZRo4Ri
8OtWRcr2Eo6IBpcSpEwDechTYpnV2+1lNa+M0c4ZF1QLwT+fqYCZee8jej7N
tZvZgIG/01ymJSDn99+g5dGhfvxqP3iOZPWOEh/fVUTu2XtBRrJsaE4Ucnm7
TMMNRvoZeU76q66TREwf7M/PB2g8q6CRqS1e7czAJZ41uK/MZTVVXh138U9G
y8cjlT+0acvNGfRnOmsw2g+2IT2YE6BwIYu4KuLYsCSIgxh5+C39Hhzu1fcY
XwdbWC5D2XYgnE1pacc8A37ODfTk08ogNJTh0x2SIUPFwqlx2tbR8sTyKML+
vQlNBhO7U6gGg0ZBxh2BX8fLC/FJffM5+7A1vYZz378Gns2AByUIIw71VJiz
ONshj1CKlQJo7H5fzxr02N3gGRvcsi4384ge3azbo+rjdTHYBkFLRtvcb6h5
Vs7wi8Re+thJILZ1I0g81z45ziM8BJ3PBNsZhOGiS5EzL1L1I5bRHJgg2+YL
8Mefa13Ve2QpXksjudiY95Fa13AehyLORA1hP+jbQC/ywHB3pe1rbL65Jaju
EYFkqxyZ6bmwVj5559e1S48K7DSowqLJxIQuaYfS+aglYLQXk9TqIgAt2RO6
FpByqN5Afq+gpqK3Y0/tZaalJBhejO5xo8wlfaNgcrtpRWtkJ08DiiPK+7Jh
/qSQxTgf7TBPktHIptcpMEmPQs1LdNNFKpUee46HvN2pwLvrRSnJekl4whCQ
eZFyIw2VXbbbAYUb+Yl5icpkhgHbkPmLaFtXgDhKC9vtIKFA5i53T2nfr7P/
JRxwr14DQoSr2b2fFfDXT4rIDEgVAls+c4xCwtV2GCpBxC5heHp8181ZKY/B
tJr30ZD/YrHx1h4WOBd3OreneGQqufiXjAqVQ4xRy317eyI1Tiu3zDlTXeYT
q9uqFKfpD/NX9XudxAQdjOX29VhS8+tU5NCw27AnKkX+jce/2Hg722U43TM1
fwj9lEXS0Hp49adqzHIsLrln8s1K+RHmGcFgyLcaJPskB0JJO0hN/AlzLawu
MBwxrmDE99pYcCn7XppjieUPOliMijjmA+Y7EZkqZIE322mpQep4NjUrv7yj
yoVqdMZkuSYCEuSJ2Uudl7hdO45EgCUZogCsclB6dHktPfJyxC7zwciJ6Vy6
mA4N0uu+fW3p4rg9EoyAQXgvP1bXA2dgTbmridPaC3CELuXmftAbB2xBf2IS
9l4jnIOepayCz0UIcclxQaGrwVpJFAUc8T7Zk11Z3MCCQNr+iBIgKmu0x7dM
0+i+tr4D5OU/aF5DPuKHYTiMWUqrHSS7gxrWZ2zpYEQlQNLTrwIdzGrINNnV
igeqJxlmlypI10jz1Vc8fymUYHXZXjz+PRCvWeG+GHm6vHcsgFeM1wB3rHSD
xQJo5GrYG2tN2p9Fl+Ef21ghs99P1hgZ1GAfyat5SpqZw2e8JYrNeYywe46m
EJrjjsAf/pBRS4eqo6zhWAqc2QFudSjzmtF3juvHzZbTukDXme3c5Lg4R5n2
PD8IWjZKIzshstkCFKR4t7ToTMPyZoarOPqSyLtkh0llMAHho6MY8UNiyzwq
VcULHWl6Og1tQozh0IuO/+oxgLLn/HYISiMYGX5XkvK2oqVUeiT/WPsDi1ri
CB+TJm9/i1lOZkUra/EK9rJWt3EM7psJtFHnV9Vi4tsZdZ7tQgy3W6EcLynC
ukOtIvEhABxFXBBWykY1ELd0ntCUB0Hjc74oU+qG3e5jX7LgsLGloCFN+/GM
qDDV9dUbtDlMtTBOc5014hy1aRmtcCsDh9fqfFp/hgl7zFbLZmXCw/fdGKoK
Pb76/yLtVK7++9Xt3qY8DE3OFWI90nqTdOxvo9P+ZeyeMGg2oEsi3oiGREbp
EF+bk/B1dbW7MxdeLWmTvAzJCpb3cKrRoMr6U0PdI/uQCTgiNLurotIsQouD
hX8g3gl9ZKu1lo6kMoEXoFVpMkbBjGQcXOeR37GxXAHS3o8c6By6k59yJNpD
bIYTBVBslo0yltVRREZIWonSAkYqBLiWA+IvPich5XO8Rp1z39j61RaoPPuG
Mo4RKIEn9a5HN+qODfogTrDMPFOrxYr92eAGGmk34YOFFp4qfGYp6mfJ0puI
domRdHAdfMACM71v9gDtD6hMR5X/WDBMtduqCIQh0Mk48F4ewXwxjAD0O8cv
oub+15jic+A8CpAY8L+vSiDbMGUAfhknLfFoVbeGnoJhpAo4/3L/M9nImCi2
PIX1yu5pdlE5KNPOdgqXDRqZG7kvMFxGIslo9N2vXqj7p6YY32tdT720RjnZ
Z0MtBSxkM7LxVM8S3rKTzlpadwauxuHPwwINCc+h4pwB/1guJbihCskW3H8s
xJwxxProLfEsaDRa8ZVl6G2g8BU9KP1jdqAZjjjdqh6ssbA5H0W3pSK2DEOn
zgxtyC1u578w8vTA0dgTC0avP7VaZwc930EO4/9Ea2IYwKpD2A3vqXaJsCKb
V4w0W+U6lhRBI+CaOj9BYs/ryd3QkY0oybzwh2Yt1YG8TXFdgkBmq8ttSvHP
tYrmS0zXyxuyHXwnw0gLa/D0Rj+UnqJkAvDIQMLNR37MiZ+vUY0KeLE/A5A9
VpHoMp8FCCtcbKlgzUIAG5SiMR9wa5IJFX1DCXskwMlRSTsRw9+k34be12kO
2hvKFdkavdiP0DuPGOo64ebZHxyKSnrGR8ZYncKedgPyVxiq5dyascH+daqO
IHphU+TTSLUvjvL2HRYISHu5u9SK7r+8XwQwUBIVoYuY+plKxaXwT4YLPuKd
VmpBlc0k45aM7UWqAHrlw7jBDbWgK0iDNr7PPIAGeJkoVRmdRPcfuCztW/Ze
uxDG/uCDZuOalq9Gk3rmwasLrOgO5tp5GT99H9zCNZl25aBKQSLmHXxAQafN
BIVPC0ofc/Ebt6TaLC+krFCj20XIQG1zfY92JdaQ6Ef8+jCETLf859ArQWEg
WxFwZ/XvHWrwd56XjeQvXqkbIhAzF5lclAPBm9LhU4/47774wEJM4YKKJozf
21uwyaeVyEEXa0L2xR8Cqnw1AQCM8XCJ3BoF4EFKkMZtogVFRo/pBKr5FXPM
xUQaF01P98CUqsoZCxD1mhBaK8wI2YHJrV9CJniifq6N2H/frJIVokEC1Wxr
kaB2VR+TTdMZOa3L9HQs6GApKG4B38rU5Iwb3SgnMPaM88OGnPp97tG4LLIX
/4SxNLSmjSk742KsXIZucxqs1UO5jRZF6z7IgbfhPs9mOaOZqp9F/l4u3g2Z
Faro1tsR6f7zI1EuX+axtUIMdPgbnAaFCE3jaT9FLNKxwKH/Bo8mXv+b0YuK
wkT41Jlwd+mCm+QhIdehmg/oQo/1RetCR6qevlnDBjJgO4rLGNHKu/7cWGMU
5sT5uld7H2roDf7/48pG/qGB0yzhLctpIKSowvIVNjrKHMf4HeZHfocKdxJw
nZUbIHh4d61q1aT2UkC8bz90ugb8Khbjwp6BMTJGFlan7W5FkGnEou0OU2OM
u8EBFdM3MNImHIXr/+NkR6rSO0W2m9VF0fg3W1LibEPvDx5OoFxSvU1f1eQ9
ehD5r+tZxdkHslqW7fo6ri8wUWXp/WAtTfrQsWHzelPgblA17t5ex9EARb8l
fW0in05QH7hMILr+nM97NItdkpv0a//zPcK3XJE3LL+nky0LY/P2NnO4FZVE
9I+oF8DcbyD24eNX1i76HwO7JnVe9V67DuZh1lAqrJFx0eGuLPeE0eUXqnfg
pfT8XG6KUG4Kvxd928n0ItxuVONGGNJoN1KlkSl01eoF29clAqELgBa47HzT
AqNTP8ZEA5phtT1SVDLUUTd+OMy0MIU0ombBVBFL9ZGfEvHfnn/0ZXFAXLDq
bEUJqY0RZgC250kgK2ieZnXboh/EOoqe7QWNeOJ5wn8f+UgTLsWmpAM7Ji0/
Js83Gx6FjaE2lLWBuboakThmO05hRm2S+tMrHiCCdyqqNMRaoxvyEForqXNK
APrXnnOHTtufxt7yGaOoJJJuP0rmyTK7+ppleiGDs2VysQlT73GLcXFCCdU8
lDoIXHj/y0GvQ+GFoRR8My/ViDs+OsKL2Ds4viTCg0nJnqX5RokdDdlfKxiW
SQQbL20eIEIWUcs9hbzrahZiexjn3BSbMxfI+zXsQNzaSaP/fAzYDc3D6AQb
g9DBJc3+6dAfleY/JufvjEsZDfwvQSBTFJ+sySSp95/+ZFHfyuy+/vV546oU
IQxRmx9jB8LkzfOlN270Q4O3fDBj8eKgOffYKyKHKW8uVyb+w9BopYaQ5fsX
7LO0C1cKzyKSVB0RC/Ydki8MBItqQqRWjtV00YXrFCgn6s70CY/hIPDEamdo
HF8jPWE1pJGxze0rbnTj+xkUUG+7YgB3+3E+OOo8RWZQOdZjDzTiQFdibn1V
LjbYcZ6UQpIRgWMbY0TmOfeV2afE8QevAXER2GePluVsAv+pHKFu5r04c3b4
K1P0BlacexlrFjhxb0qcJkHecg8HTKTCpKAKb5UcomTQDorMGRd81l9mBMhV
sQZFMh4g3ptJsS+eztsGVwWyqwBOLgo/vYj4U7UTbRPL/Qi/04cl0sgB32SV
ebUYn3n0OvHfzJN1tXslQRzYhGB611m7kkHZ7XDYcupRAKhzUieglmfrJPsF
qwsMhsWfUXlznV8mPIDRXLWuAj8wnhzKI8KD0usGwhMVy/DnYhHmVurw6dFi
oCAa+dpm+E3BHZU6aewGcrjQn1C0XdUBDDXP9OPQt+iUEOcmFMmtE0hKQZbi
pmIYC9zG6E3VL9U8/Pj+JSNhOXEiesPy7ZF5AiITh2u7DQpK2JvARbYeL8Hx
pGLtgjhtzXfdjTLH/MvzakMP4vgQsBnvrnhU1DgoyWvftBsaYxiKKmtu9JVx
IifknpTBMj4evn2CyeMttVV/IatMahiklPB2hypequm6MPX8ppIUvFViV2eo
zN6A+qBxtqXtap3flWz9p/dTvkjCSxQ0H1HWBdIW4sBAGAhkosDVto9CEOIF
yEJFMySZqHFDJ/Kmat8lHSce28kjprf33sZMwuGmZ+7nExMYtgpgAq8w2wOu
GsCYxJzstFpFoCiOJGU03VwfkhJx72fE6xHjwnDk/YE7TUYwfU08kguRu7tK
Vyecg9y239UKOxeFNNg0wg1Xz/q/RbVG2bssPYQ83ZKbAjvWqheLXpxTMN61
cyxry6vE2cNvXnqXaQJNAABtIIXKwfbO8UfE52x7JwY5/ph3JHfhHSCAQwrj
JD/gH2AQMbs6djvvoMGQv0vMyEyTmoNkEwzlW3ODZaEHz72DmmXzwbEmEJL8
72sI08DNAwpqZP0Hd/ZEZ8OoKgWpjfFOa57ghpFwio+iBmwWy6kxbmhXjLAu
kf8thTjwmAYCngs2P1vR+sp95itv0nkfIFmlu4ZyehF+JolVSGo8np+h3GIW
yoz3s4vKgbmI+4l1bUxggjezwvMYaKM2XF+iKq/NEtvhuW/CUOHMWfk0c3RM
5F8lXToHPyY25Wy5rmkdIGWcsAfXS1b5gtQhw0shorm+4mkVWQSVBwGKkqBt
gRvDuJw30Qm5ASL7bweK9//BcvLx55nd7+RCALMl6WRJFBAP/XIQQSqUIYDn
5Pnp7mfXilM+VOyFM3ZIhXDChLXGiA54uhkG23iePhdXF8323rs1bg4nricY
bBElktT3NM+rcuezJAAuDEVdn8juEgAkvfsWVzN31eEYhHpVPZWylKEP7nv8
EeE4u8V9R+vRAJTykD+HodBOJeaLb+IlXF9aJAM40Ww7gFAaLXnqzDow4dNg
HGO8kcwLmYkEaufCxXElbvJmNJkvBuFwDRjQSO8b0B2jx+zvMiyvITmLQHoq
ivGLB1u3ma+UgS6yu/pdLZKCRtoFwvel2bFwazZERLgYemQSgXWxCOeHT0x2
zRC+/OU4urveVYaLpcWWXyM2C2ml2ZD8Ng1UCSWBFn5rzWEXmod131NxTE0H
QImbxfro4NXb5SOM4hjY8AhLUBoQb/LlBKsNN2tHlFeizyVgpuBDXyDOXUG/
G66A1bAtxyk5sKiHYZjn4Hppy6FoUm2xuG9oiSMZ5v40q0nWCdju+zVnabbo
N6eEEj1hgsEHm1Xv9OaAnOdS8LhL8Dam+D+FmcPIVgL1wF97H+ZEhSspDDbz
3gkN6zuz9qnz3VtgqGcbSmNjqc94RU8t3POuTVY71fVg7oiGs6DKDwEuWpen
QQlH3x7dmtusn5bVUxfS3hOpqWFpPEaNvYsid1DJ5PuswARlvr/Doo0NpqN9
rEqJwLRYrfHj0lVdwwpNM6QFUzNxyHPPAt0tTTXlyrju5lMDLy2O+cPISGsF
RObtLik/IG82d7w4xVJNctLiZGssbUFRj05eiliJvajht0rUMC93fpxAuKHA
E2wA3y6xGlsdbWRLJUrVdC5ZxfKuMpf/W4ivOOsXzNXStYn97i79q3mmwU3w
W1/8h0S6Bn4Ua8EvvHS+Rz14821jLmJNv1Mz2d/lOAXX+UnWB9cpMdEhPWyy
a8uW+Pnr+gVHXiDuFQfDs3+WwhPA4MZNsfh4Xw6CjSxOaqegO9BSmTUU2Zrw
QnzS+vmZxyTIAknceqwdZIUEGMwP0xRDuqVLNAPS8bYLJWbxaq0tAlAGiQgd
yoNKS90yVn/0HwLISfI5lZXZOumCr1aOTwC+jjT+wQFINojbrOo6rUwDePwI
9aJlWXBLAg85yLH0Y46MQBn8wod4781tiOAFE3PPtaWeyLZjVvUy56UDwd9f
vn5rTMn64rWwrl2ViwVBAlhzmiKeiowKD+cNisKdnsWn4PYKxkgGc4xlom5a
v05juc8fvCzhSJJnokwkYRUkVH0OEiFKRYm1fZC5sTjvL3t6LWO4N1TET7gZ
LYyBLcETbG7ZMrYwnDuQJI2FLlKENryLm7TPa+rjG2mnSEvTnwq7Rj1gNDTh
3/6vhXAjgELQv/PICkWJxTmUrrfo6YI12m2XST4GeKFZLMm72AQ7bnyuEEys
G5DMruPrTfqtNQgzR78fDYHPCVoX9Gi7WlKRMhpmAfOQ0WETPtv0DnewWtwm
UFPlMo9s/s9sTLfZuVaZ/9vkfgljzomCDzF7sTETRBO5ToqP/w0Vdo287jSm
ggwLRq0BY3jm7hRj1qXFJS6LKmH5vNdrnxIpbwFqagqGXErf6L7IpvTdC8Kj
1F9q13T1pLKlCKxV/oBPOVuJDjbS7LTsKeoVRQRh4cNBCVSMra8RfRkv4ZLp
hm8kKjdvnqp4/29wCDjzzADPyQXx1OQ3zcgV2EN0hBb6GOh+qsKI0c4GVfSM
ZDjMFNz2N0wq+hbx6r8awaXIaahOMeQWHOqh4871As/5KvKLHm2BJaV+wkCd
r6W44lEqP3TJGZSk5rOPfz9hwLFhbtkzkuFwL2JIMMH8IWieH0Pnz4ga0srj
cev+HPEyiv336y0b5K/37QdUexitnAgpeqpmSLOtE49PpappG/qk6FW3/i46
y2OV/PBh9HfjQlvRtrkk4UWXAA1iuHHac4UMxeP2nfLJRV5q32oVtWQ1d8KN
gSIEXHasqDa8MRUAMlp0KIvTE4fwDnirMVaNuwON7GtVPJBRgc5VA9Z7bZCu
fGjxMRNV6f1Jvc9mfk0Cm9NKAcTP7KPIyirDAUKrwGLQ+fuR5LOOE/tGnAJ0
tzfoF59mqC22h6Xce9AR5x4N4w9YL/XBzE3ddERS55LU4T/19gXkszR1RVkF
MUZdJLaRGtGEUDlA+pSOPBz0nf0HyYy5asfKUgbn7wE20isjwN/+jQhTr5Sf
gkcmpxn0as4ND5u2C72W8Ba73EYbp2ugOzMHy7OOnmaGqZXfF/OL9ElczdBL
eVKr8BylPGYEKuOCnKaBp4S5rpKE/HGjXgVle2GdhSae5zX3gLgOkNei+L4H
SM7ju1lbtpwcF7+175WcLwDB7pX2fqjQJ3aQn8XPhumTfxxyzyO/MoKkt0wG
bN0nK/kR9A7tMpzu+d84mb9WrUx5iCEO6x/Nhpb2jW6wHO++7zqhdAeN084V
6YLT/RGYUCpK5PhpH3Xr+L8sQEAltqH6YUWCwZkSlOcEqeBmoa0jBTWNZfCF
9NU4iWFL9CxuI7OUYWAWSgP4kcPdQNtKVw6haw6NINEOgqqck1u/xO9vjZyX
j4rR7E9PRMddYa/QsoVzzAkZXr5ZjUMld8Qggxj5YI5sBicyv+H6FwHiims/
sL10nla/VBYjJLUt7oHe0JxCQUUgjcYVMFTuZ5QIEf3NFa8/b39aLrhgPn6z
UNdPXR7zc3EMTqIvuMWI5I6zoq2sFQW0319zHoBseLe5FiWqW4p+FcFa686K
o48JrkV+jTUIjddos49dgYn/h4mCZVPeuISo+FNFLSdtk0IDCh8nQUVtTLG5
8Z1BCpaVtuLpQtnjVabQShotksjTiP2EY2hYCEbCbE+YBRB5eLq2AfyhAHcc
KxefPj9ig4a3lPJyqHgrnGdDzJYZ3HfqnZMTIINCdJS6JnOViUQ1O5LfSQL0
41J+t5kCs6CJI0EAAoWQe6tl4YkhgPEg8K3/IUvRo+VdBe3ADkFBB//Kv2VI
axdUH58V0erFlc5T6TOCvoqrE6l3QlXCdsyj7kaLXPDr0DBhXkbG5x1tn4F1
pOZWugNc5kEVhvjNTGyXvGVgUau7rHgSwtv/btqjjXzjU1UKwTiNRBbGDRI5
Qh0oZCSArrtlrd23XVlvLd0ZHY8LT0ALOes2n/NntMFKnpEMwSPOGi6T3Pay
0stqHnDyg8ZHSukxwoCF16Pg3sk3pDdmOipJTjP/DTgu1nFzvCznlzHvJjj6
z87K2Ao3YhdSes+1fljo6zQosR73qiDmySk/me3ucX6xwMTMAdMx//LvxgL8
RuRZoF1ATPXNu+vACG3nQ5iUO9OmcRv9DZYZIMCvD8JNI6TT0lGynUvnuEyV
xLSaJJACSPp0zLm2ojR63V3GHOKGGJyVsxGKFIJqmnv9zr96GnQuD9bkbvGv
odriJL4w+B6ADtbid+QMDjIzypM8GBLmiOGU4XaDptBoG+fjmib4yD8x6XVy
df/OOFC1vsYJt2BbjfElKAh5DOv1EWvkbyT7f+Oa1CRAvZPzHwCCdhPRU1lA
i093Yjbqk57U1rf6CLAldSRfin1KJ+EM1ZHDHNudF/5NdbvGPWrYNYWalSaL
tcPXjNN5UhvjNOt7lJ7P3o8aPKvp4TGqDwFappQ/5mdFLhRqb0sEQ/GRfJQN
oShIXt5vghNcIU1BJkxUkCh7R+gHrkPdfNL9GhcoJ1Q9acsWbeUZDsAqTaTu
JLPdvsbnlo2cKdH9t2uEmPMGQJE1SYeGa6XtGLxbW9C/basdCgkwNcm4ocmU
o1nsyr+OZyWLkO4iF/qoX5BeYiTPI0PtU4SniexdI+ZCYINOxKZ10hqNIn58
GnILupelzPf2/EGUi1HmwkgxXHOIjR4hlWYxRoyODPIPjjKkO0JfjTEcCPCj
umvQ54Cdeo0PdlQvhkYKJbHu6bafJXVPahdNZBpmTFq6FNFaVAyT/YEPQSDI
/rzInpLxkTY1lqwIsFGuXKdqrbnjjPeiSRfmhPn6OreJMfWLm+oprdygNLIf
zJdrzywYIBo7sm/sZFHjcK+dkGAI43GArTXBPTYnEYO9dRk1T39+tbpGaZhM
lfWtYAP77fVmzG29757NWp8e51YyYVhD0e6dbxuqCxSb2Y2vtOjd2Gscwkyn
kkjW0g9ZOmA4+JaTDHVIa2ecOQnjkJzjLmWob1muwrckyoHphsmY64GX0iCX
zkBC5giordD218auxWg3guGkDaFHcZTrATzvw5BWsHhVvZaEvfQNrfBAHqPd
MXI1HpusjA01pJqM/hRqTbBLU7msQJP+GN0zDSwHmHjn7wER6MNPWJfzZrPK
bIfbVwRghRpKcdO3FQydoU33/Z2b0yLx7jPMosaRvHZ3Zk39hgW31ibEOAVm
1gDSCsdlMME72FVM0v7mL78GTNphyphgW3FZR8EoXun8HPbP7+YKE08OxY6d
QtEeOMHrNZ4DAv6EheM7sqv868DwhF61NstWSEIdGuH/nIkqMo4c3ttK1omd
7KQycnN/Y6aDY1MjQEuuBK28dwzBzX7zYM8k96acYApy0A5t6CUgrMM2bxwc
JVdZniTlzoUGL0x+6RoC0/kcAcfJ4UZ7lKnqiv0HjMjIbpmUDvECU7NCRl4k
Snoq4Jybf3UPbgH43/Tt6YPTQ1sgQ9vzzoo/1ta1IedEHN6rin831BszW2nc
1R+l3JY1XtIqEcljq3nOyuDlpx47sy8pUngShB8Ern+zCNEG92GnQHmeu5Wn
EhOZH7DhpllF4wIWAFslkxum1ufDbSLLY0nJdibk1yFW5juYBNrHDdfEfcDl
h9DHVRuBSmmTnlSCk4mj1/4bcrsewgeh1DkAr16LuxCBOETxRgRaDehub8xO
i33dOMzEjRUBi23vs16SFJ4mE88SXPGisjOvVFxK//EFpGGrpVYeYMnKJDf3
jMUR4zuqV8Za5snZAi8FIv23ccBDfVzEBGMDUxQlPDk9Nch/sOwKpGYvnD3B
M8XI6XLNA4CvXBxyC7eRWYZx5w5gcoQFqHG+pdHHAjIOn4po16+T05T80U3+
41+IwtXx3zdKaLMxtkGiAnga+Mt82IoAD+lE5OhsznYA/2iInaYIu1EnceHx
3wXsHb0m5dzLJmSZybTCnKs24SBxMeuxKtStUYYQk/ihw6+ywBdrWLiiL5Ts
onH/xKdzjzMyaCJh7WXWSG+v/tPbrHMsYbAav3hvb2lRhP8V21Sieye34oWc
88IhC+9dbU9LZENsteFHEugBMpbQchBHfWViVgS0gAAtWbpN7W7pP+4mKAjW
P1e1QC8LsoH1PIlRPRu9bglXID5eR7dpUSn0iYilQy7J2n6f5a2cyyOQifCK
lVL8/IeBwRxNwJGysrenLwgV7NVVTLMzTiFypSZXwh0fWopw2uqviYjkwsdd
gbpxqnP78vgb/aLA62Q9/rwk1JkQz6Xz25klw0+0w1rApTwBmdXoRs4WP1yV
zYpwXwpGDCj6ahs2ecw5Pt5msTABocrjySRZH2OviR+9SJCEIR56eZV0aW6R
gYdzfYxxWqmGD6xugfG67qAy6dg5c2iSRG/y8S+QqS7Vb1w+hZi2EJwIGzI3
vpfVK+lTNAQGMO7f35JdwSvSvjAy6XzJ/L7XapL8ma5wnHYl/pfml2qVFb+W
NI2RkILFlc/fL8HXqYm4ZeiP2jNRfjgmQXJRNH7UQ3lLbpBnnv5B2YWIsfOJ
57xnQ2JesInXy8jzU17iAfOwjqjMtXtyJ3eckbchKfq3pDaseAcFIFDlAVKi
7fNeXWcDpxTdKOeDa7m5dIr8KUMHk2gggxMoqcfyNexWy7ytrluM0JKgZGfk
wV6CJDs+zTzKFIARBsdjBczhT8v4a4X43Qv82vmv+atcXCYVmIsr9MfH6zWn
j9XbjCCPGg7PoZTaCT/Fpyx5vVmEDpj20FxBMp8kiguVzQByOALVjp9SgGBn
eJ8wFxHegjLpDHLEwXqYc3ucUX0BlgSHR2030fRplAtWHuLiG08AcRBAw52+
iuWGl0EMLO2+IGvs57DeOrY/Oyy7yKIA+3x0r3RwsVs49157dzbMJ3BDjzQl
Yn3TMQMUj+DjJV8TblJ/nrVYiBYn/p1QyeC/G3By4VURNbnGL80voyy4x1At
BgjsTyNqvZ7lWD1SIa5AMQs6vzxW5JPXTrKBTi5Y2UClYMH2+IZG+0G1RlWQ
umV1UwiDdUCQX96DUMyjG5pNrq8sQ02S/4aUSefrvu0bcY8v4e2RhAAjjsHr
1XTEtNMfC8bdh0EvLAbRNzDcY8H++eEiWJv6+aj5dP9Y8tT86pRLfUXAGP1n
dJoW0eOkaBdqVIYsWzDZ8VFugmVp+Ab3WdpU5aBq7SUijPyKMJg0yz0Ie51a
KAciTsR2fhw4TDKSR2W4UzZMgTX6OC294f74Qc50SDfn59l/g+4gHXf8n8fH
M/Gca3kEMxqBt+0ELSiKDz3p6RyeS6RIoK6CUj/4wm9Tf6KDXOqzTV2CpEtA
hM1STy5OL/58qxAdITd2X6gsBUi/QBzr/5BF20/braxwki1iFt3HgNkulwVC
UMoafZuLmqVb02rwlFtxM5O/RWusDBEdiaWHY1WtP6lXlPNbYHWk2xppznZl
nOg+5F2WYQS/MUspkHapMOIvJa92F5WccDJTHkwHMN9vyL3/SdfGq2IEzKpB
cj8O6enB1I329rLyork5W7/ouLUV8HXunKjlDnuk1rYkSMQ7PnTRSFRFUmXL
sGJWkqVP0rsGXu0ysfL+mj5Uq2JWElSc/Ou3R8ZH/sMhd1tQGADOvm8eHJog
yyC11I9DKg540OhQ65oILScYambVe2qKPrZHrpEKbdaP7uNMOK1SZv2/PhRc
OysN6tIenC7I+FczkGYC037f6rmRKr2zBtXcfVOtxVK10yIAKPLIYI8yp/Ye
3yDyx5VFz3XX0vVTCniw/NUe3G+WeNjGUIJ2/3eTbRDmTyEp4Wc4zZ8CjNRX
zFtY4ZGCYJHlcluahcbXeYkqvNkzyr6taXMBZnGQ6Ya5nAQslmg11Y+TdYo4
WLUD2b6xAJoZDjZ5m3NCOQUjawp5mygpdwqp3UkiptargVRG/Fv7hqFYjvyg
f0KUvun1tTRTRbe3Wva/DxwQ8pLH3bPPOZESAHY1cCKTWnFDcdz3e7gbaUo0
AEGpAw5rPoTFeiJ0/VIf+C6s7bLKTv6gl4VQs7Nd5oADHDG1w8yi4xf9fL6i
HYWTv0onqwAgDjxw4rOWjPpe1qU8S6cTuFKS6MR33EHiyYHynqktE1bkJ4xZ
xj/T54V0bpayzwDVPMwBxO8Qa24ZzG/uoGVmEQe6rBtn40IsuVDa96PA3CII
qtxdDaTmuTDHzPDX4pLrikRroHV2cancwfkWmk9VND/4DPyK5OlWeUn8XGWf
Bxqxa+IbhSqKxSBkYES5YvU1QFFrjJLA9tcrsl/1AwRcqF60ABsCF2u2JBKn
WuTA5US8prh717eydWhrMY9pSWUZCwFv5JPiOvILSrCMC0dseYjHpMlB1ixb
1PGDi0AVy3g6lLU3h2h6/+erkUyBqlfYNHOaP8BCVW1zcDDOvXD8PUcxT0Dt
Pb/K5wIXcwZn/Vdb+74DqO3k1AbvWjAtkFZBQssWwBX6DYZp2QZQnWom75iw
+iJIX/ICwffRx0q8N4ok1uOSit/pUYvLIpbLk8Ra5xyeE63Mq0wPZqeUCHSu
F85PvOY69LmlPuUVhIkzLmj0uRAyYpjUOiiPTg3D9lX9wIYkCaOwkmQJ2n8t
QQXdCK5UAljbQITF07K2H1TwQEz8IpX48m9r4SkWwSIeCju/KMoE8ImxcZlK
TZBt8lBXg9EbAoQrt+n72uGoNYO7eVPfLdW3Wh27aBv12kHVtLFB06NdxSjt
lrbHd+/gmVtb+2sSAHXQTmn2154Lpj87OZCNynC4m8OyjgTy+wf6INUVZfUT
bRANs4v2e15L2him8NkyktU+Q0j+SCEXEiROxUHVukU5LJsgJZ60kiTQEBeq
jRsTzhAdEFM+iPr2io9LjIgFiqSvPUPw5LvHMGMfJFanCF0lcvwuOeuQT+QZ
SMpccIg/iuyhkeHZPqFzhZ7iQycX3VBg9RL9RvLcs/2mNGYM+00K+h8K1M3u
IEkVQTT9zn+iSg1YHhqT+1AeJrFvH2fgByrCMZtWfKn4OG/DFMTFaa3yY5VX
tGzUqB7cTyzDicsHcqFxkql9WoaR3wyOcAAXkPuNrkV/x6JIKCvrdj6C2l6J
LX4gTUqgwcZ6u2o2oIK1UQlDgnw+ZFfFJbHaJoVfMbXW+TEUDEAUOyH1t9ce
5xmVpudXudbIxCwFj+QirR2lVgRB+KrZlHflEpLHBP58nT4fXSbh7OHmco18
C0D6kLFJKhER0a6fBPV3BnvkPW2nbqOAQcSu0CdyB9Da6BHZdzZVo0mOQKtE
3S07Y+8ZTgy5TyyRtdBM+DkI3JVu35wV0qCvu5RhEnV37u/o+UPU4WIKe47x
8rOJxBv0eeqlMB+Voio9tOMkaEHqH6jb/i9wZhpyGkHJDN2inO8EbIOzF6HB
qILm0kommBV/nc1inOz4Sq3dGYZAOHYPEumnZBBqEYGqhmshAjoT09F6nDkW
UtVxh1hrxgQTXmNhK5YqaEiLbOrBQzMEdpu7W8ex/r2Kl0NylJ1KgQ4WOvIQ
pAZ4Vzg1bDMhyM6YLClAGXVghRFAc8ofSLF7cy+cmBkYzf+hIRb85xPOMgpx
YB0Kecr7YFYL7XsPT6FoWF3SIA5kr6CBt9xpoyKClvwE9uoIOfXXVXyx8l+2
karZRf5N8nolRsXmWFKxwmA6bQs5I3us5v9Y59yTLDOeGeLkHPV5oaxcZ1XN
GCVYsft8DLmuujSeFCSAn8Odq2S/3u9WzucdEUv0ALaulnX25rdOqiraZ6PR
KrBarZZnqOz4TmU19SzDlNmCHb1V7c3n3xJ5oHqnOoe8ky8/8F1fNLQ5Yv8i
e1cC8DVlR6swyCCf+e8AfEsYo449GBgJ5q1l6Nqays+i+9F5gl1vPtk3Ro5d
orQ0m3e7IDr/P0zCl2SAR0UXSomEmrfCX771IuPnxBeVTJsR1G6myAcpSp9O
9e1dkJsNCVvzUvWF9wm+erNLJRNU+mlhSSFzfKcMRzSwaWURK/B7k/6PLjRf
7shRDlcvPS6gkJ/KegPqcmohCCixTjMGPqHfUA0iFTK/noLGOwZ5Vd7piu+7
cMNdWP3ZSIyr5dwNeyE4D41vcycnJ1y3A4pqZ0hMtdFOF4g93NsSttZpudWM
A21SikkfsKheOEuaUqB51NkXJP+JM7Vtxvjg0APoT4b1Sp+F5x6Y+4ylC2pr
gJqMed8rt+Bj3o5XwxWqL2kVVGwMF1Spr38X9pVBhwXG0NET10f+y9qJHRSY
M3mei6LkcAHmB6L6X8fojtUNev6hM3GrpVu9tZKjP0lc5bwdaf/16sAu+bEs
LU7lMvQkvg3DXpNJGVsc/hE+I1juByI58t/p9gz5pEFLovR8+dVIem/Wtp//
TT9pkyDzaGNOUYJQYJm9ASxtfuUuplyviX7leK6i2r0frTV0g4EmAYRJ5cP9
uVQFMmgCoNby2U++olCHz6PYaZSBhqCHiufli6WC3Y26RfsGcG2Cgo84UeHh
Ppls4rDUsBZbWvKFVSMX9otzCB+l1zEyaWIXhjrguLDSucOfN955bET09Unq
KvA2tt4WNfRBnE0BiCjDxCZ/VLe25bjVbLC2OieO+8FMb22UBCJMd/rUDLaO
XGs6UHjANlnORLmdvUngF3bW0Mc7f3qkBu7UyAQhBIBTwNWuI7tvkEX5kdgV
rlGNNiofath9rKK4OfkqUFgkG+V03773oW3gS9sPsvlP66r8ISU7y76YsppJ
wL1q0Eqs6rb++cDIG+xX7uwshhV65VYryFy1RPIBIisXSRljZb8yGdo8kxni
/uPbzJ0eGBRjm5aECQbMK/IgOw7w4wxa3UO+D6lkhLmXR+l0MPd8AM2nZNxE
fqzYu4U54d1tlZuW++rUP7xPUZKZW1woOCnlTmJtqSitJZWTQXvScqOnkFCz
m0TeDHiBlJI9pd4oQ0d6MrSJGUmYEVXEIVfsAXIjhWGrlRFZYonvihoL8xjl
TFL+inVrEWt4NA1I4bPCI0cr1Y7k5BcnQ/3X45Udpyl30KIaFtttomhX7OIf
vV0Mo1OB/8aU4rGn8TQpRzV1wGEdUVxXlK5yOAdvMrM16GzytUuEPBa+wtgg
hfJdUiKAD4Q0ULQ7Yc8+kIcFlDugi1RnAQb3ek57soqKux4Rx6MqxyIdmkcI
cXiMm7zXqg1VpNNBNANaQsFc97sh1JdBy6nu7iVfhC262PQHMXRdsi7VXbe7
auVfAo/c30gW/ENmNNeTEoIPIY1644jkcLxkLasydXdmxE6FY1L5VmwLp8CU
Dds2C6M80wzItHOc8H+fSUr4GaOD5Br/l37xVsQjoO8nbZCu8dggT/M2C6iP
lyixY8+Jztlj2ovMSOGvf6Ei/2qDHZl9wYF2Pdd8q+737kUXqqbH9HpsaiOd
xQMrfBF1W7RpBmcAJf5+CmWp3YQTwf21eKA3cjRq1V8vt75+ujWlOfOGuatU
4HmbJetCqqEr5JTOb2hRbwXjU1y93VCxKv2oqwuCYK0oZcC8lULrqHosuDT8
8vbfz8wTXdDS1uKGmoh2csR9BPA/w0s32aMo77/IhgRnkWSf8voV0U0gbM+n
+RxXmbzWCvN0n6Jc2fQbNkPXNh5Pt+WLt3tnhD+WRRno2IOdfDQAIxnExFW6
RPdQiGvM6RPCegVLqL8ozeI1KUQU1yLhN1xXAtNhv+VYEp1pFSxc4I+YdHUC
ENi1zAbChzlZ193o7DD/TXCUY6nzlmrbTa4E0lPfLE9Rjmoek6pZBy06UIEt
0FHybeaww8lxYP8TXAgZgydSnWujdMFXvdQDjSKnUkJBRE1eu5tyszvrN8nS
FD3cViWIBvYXrAbV+ugPHtS6ADvHvBhZCb9EoIbRaOTWg1FSE/18Zn2pm5Pv
otviOny1Na8DRE8ixhQCNusivzM3PqD/PqdfP6Nic4zjJHsUx0FHJsYqa46w
MrMiTEZVv9/z5XmmEKPAIwh27nucPgQtUe2EXbH1sDeqJg4PpRddDK3f4Ita
Ow195C/9TyYj9We9pYlG5YxApY2SLf9OnmmZs8700Mk/driUgNylGfPGDf5c
3p0HLgm43pZr4oy3XHyamiW7BXm+QDTqoR2rXYe0pDwL1IACA5OGEEt+g546
hbFLh6H9ItYC3y11cddQ/uwPJxwe9CnziNQn6oE5cr3y6Mj5svEZowCiG8vf
A7W2pd5nYodUc18NrUoWDzGUVDE8usHl92YgVv14d5F6CCKG3T3GxOU70vtw
cSWO2UnsQVl7pRCh/vy7dH0VYNahigGxmHwf/85iqAvhnm43t8P9j3CR3V4F
nuWU7y4xjfPL0Faql43sxsQ4TnRpNc7ZBE/lKW/nvkHdy0WKaXOJY49x3jx+
2pKBkhFoKQ8ndhdUkTD+C6Y/S715000cMvMnkF23ATpMkoX3Pu/DOlDWwsV1
Ev8rmLlhpeGwTdqE9ZZF6/l5NvKr2r4EgWvlEulFx06uclNvSBK8ikkt6gty
UXhtkN6LWx+bJYJmsX+k2XqjoDAgBt8rgGH7JuHqAdUslI3OoD3asF7xiTby
8KSXaH+VikD5eodggAfABJwFtgJ8TM3SQQoRk1oE4ep6UVRziEpF9pEVtToE
TTPOPM8VwKLwSqso5WdFIn66MYeIGm7n5j8BMPP+8DwDUYV2+dAwxKMYvzC1
bbHc2U3CJV9YpCFNspyOR4tOgtUarA/jq885gM1+7WFeNSVlL4oTrAYQdDa7
7yzSvKjg3eRJd6bVuRQtP9cnWTuVRMjqnxu6DieUvxJG4bL6MKCab/EKlZaS
4III9gmAs5kBYPY92CPXlRXhGWFiZm91ZLXSVOJlH+mrJR8EgYDccI9arBsP
R0BZrtFaA+H4fV/13zKQ/6yzJpHSmLIMyNtPbi9S9lfQsSLTk3RnWkTdVENR
FiivWYT7aoI/mGt3ZN/lxKDMXY0YhQOHiG+XLbEM53vGeutg5jhqf7OuP0vh
DXEu5v/Mm5qtPYYXwLjpeBgK0giasoci3+UeWVPWOVtiuZlpEntdJhmOlpLi
XE4GxlbIjKNr/yxIJSdeB4uStnA6PRIdp9f+wj9YheygCPuvWCVm18m30YU7
dxUDbLd3duWy+DR6HwnbnJpJKkurg+0S3jVjxYokXaKzI6bLOwjMmKfCYdIS
QFceE5GUK3XF5sVJxqPlgO4/8U4ufSggBOYmzLU9b7w1+qb8inhccVQ+b/OX
JhQ08UH/mkHuSK1SwO0pKEPpTqR+wPaBwcs/YDGR0J46nNHF4ytHFQVDrs3t
P8SAXTVhEfVrIWWpZ8X4ixv8eRHAmXnpXhUzNqH3v/OXZ+SCcnrEdqn9wBpo
ggyQEo+/5qyG7jhvMNoDBckXGBgRRA/uo4g3Hd3v9g9ltWhjFjJSEnm4bOS4
D9M6CBCUC6HX/82WSzD/kH2w6J9a1askOAuzFCeBI+zKwhnPUMLg31V7sFMk
HXQbGEQZoQVBq9C8Q2eI1PsBPw0ZfwPeayglYyWfButypLBUZzKaO7hMm1iN
ywci9zLZngzR+FTUZ/36GwJBuzWiFVAUEzt0QTGQD+wDes+QcDzO1OhHlRB7
1gLwVHP8xhYVG/Qr7lTVTC46wTE2NHw2YUjpR6YJwU/OX/X+xcBuJnv7nl4C
70DpvMFZGBoVMJAGUdjiXw1BJnHF5tyiljdupMn7wW8GH+aov29itz0zyE70
kg+dVuwQAxp915ZHeHcWXfnflw/BXOwUxpqlu7k0PVNzCZon3WgOhHkqxvaH
CgXst6f1/dkFOiX6bLEP9nveEZRWxEm0pOuRn/XtmpqQWtApmdjd2PAKoDuG
2Me78QlTbfVPewQcjxVqHFKhWxISBjhjkJFrpOeniCxUdhThWm593PVTGhaP
O2x1aLA1iYiMWAklBzUYTCmije5SGqbFej+6kAYJJQ4kMIqbw1Padl9jg0QM
jUzySv3+NdLkbDqI+d0xaW+5TSJFyD1YUCUkbZ5Ax83utCEXpnUkVKX0NNwD
PAGX/FNpQVPHMRUu8qaNERZqCdhUtoGB7gvzaT9yzK5lo3ZDSGN4Ua4hDiaf
ntHFngy+imJIwJfhPK4ZBiR2z8854rkOWDWQUKpqHYllNc0QkfxKLXnKRlpm
LYpdxnH/ixbZFwlUhHUCq7reGv1nLYmVVxeHrqPaw69Qml8LE5kkqI4JB6yL
NLHzzDUHm6oVhyNrquBaGK324MFDW7vIchUObzTAfqMzgHnsPK/HiVmxt2jW
a/5/k76s1g9KTswKXWxajn582eHGEKoKwbMWVp6kiOsjyI3FF5UGZoZ3FY3I
E+Ru1SxWIcGvyplSEJilrr/iu3wMwD22OWQi7coQsnk8zlDT8lpLQOSyysuk
Oxzp8I+tvz1I9CohZhD2E33or9dTtrbafP8c0tXkSac4DgZD/7sjOhc1+vmu
QG0F9WXHUeKZ0VzwMjXr2Q+SwyOK4uEbkexz/B5G6O5W+tLqD+IW2S+ruMC+
sZ6w2IR08uoK928DMMFvdc3W191hHBXmWeB9NgF8tPRQRVgGWMGChFL9aVge
z5C8RwWtrpV158cioTX8iyo3o9AWZsELnUXYt8HfXrq4XP/+zfhhR+mpHjR8
Vp/WFVlzeAE1DHGXSzESJYob2vrCodHfBIXXq76yXhpRpcP7KE7gD6JcG6Js
jiKw/1I6pnfBfMt7rqc/yYfcTbzMcrrncX3Vc8xVMriyK91vZ8GuWwigQ8ab
amqxsZtfkHh8InwnYlZu8Rcz2qDEarvL+aU+qverIHsf9gEUcm1GbM8q0BCK
fNpH0OdaNgnhvk6kuZL862j0vFtC8/L33m69kYYvlRDWH+7nl1mhTnQ0YLYp
70HQfGqakue8Sk9LuGG4gvgQSh5IUtIxwAkpi3f3k4jFoby5bcBw3j/7LuOZ
Y5LpwbrppQsBg6wdmCIz52v0Lq/mQ0l5612HRgxnMmkP9m120vqGYHYcBGi5
bJnHPtM4TgSuqEIIsFHYZ/GJMmz1Sr5aEyCVeYHQCxB8kbKo8SK2nMuOiEtl
hnEFCeY6tjCVtA0slrAQl8Aekhv+/rlVvLYRV8lfBj97Gmsb8V1PldhUGP55
lvt0ZrO+ah7upIbLtiVlzgclo+/jP1eu7Y+QIvCQ4XGCoPv7hfa3cKwVQvvE
0FAG/47ONIVEpERXfsB9sey7ix/O1SJY0R1IbtiuZTUqHSqsupCgonMzBc9n
qLc21qUCvAfbfeyoRuRWdg8NdbpeMBouAyAXGjmJGG0pQC7A+EzeF8PXOO2A
k4WRoUYh3/GwKQlDqwQq+s2Dt0AjqbWPSW0kMnhthLpEQRzlYoXunkJIXLNZ
/8uYtiYiKOnuml+kCZT/GngL3RFboe3Fj+5YEasnD3tQ7vJ2xRAc9XFUwpPD
6Cbyu5IVGGOvRnk+dH8Lc9RixQHM7cGHc7C1MdbJlGH3n+kcaDxq+fmuZ5VW
RW3L6FYGU02y1yJg65chpCqa67uoW2ndohf9emvPvGVLY7o1wqhwRlKTbuUH
GJPe23PRVxlP84yGrdgYju+CrCMhN7H4lVdcrWAUpzaUgUil8V+uVvHWg8XZ
GaCsE4fuv8RCJYsNST13NRerAp4mgAFxhA3/NzAzlZLvhPZW0B0DPX1iS2l9
ecgnoX9lM/cTRGH17+Pp/+chV99r9qK/LvpVwzP5KoOGrJ/9ZtLcjsoBJWgz
UjyjC/X76l0ulQQgszzVCXtAEg36EmVh7RJ1PFy+l2yvhHNRz2dXikdR8rJ5
vAFDXxFbDmOxhTfU7HuMe6YhcqXsQNxeyNCE4BiDGzkWxVeEP5BLzyEGITlu
SBC1ViuIS0IXolYG/0XxuaaE1YbLLIgOkWgeZ8DV+aTxshLMWdlUGLqqmRA+
2xLR9lMFVLZKCXwrUpLFw5wZFliqIxcCBd9KIvQQMpHDP0HBKTgndCO5eXcn
gRJ+uPRP0l9ovevO7ilMqX5CIistqGG0btw1l8KJcV3IsaJZixDJU8GXzR2I
QqU8Ory+JC6erg6nwRz53+PuJ/aV61KTtuL9lchfBYFHcIJlx1vOKlf8PRCh
7Q7T9jZF1fn1imHfBVKkv4JFhw1ls/2tjUZ6l2SLauTHD2fE9TpflCa1bcdY
u5AVGU9d8gSi787YjMX2BN+06J+VKnlEl2700LV4ruhFYm2alBMUk1v3CyRg
lyxfrha5xiYKTFSUkb3kjQ+PSLpFdV+HEIInyq4K7lf/3D097XXigY5ilomj
tWBjGRKGQMGqYrGuI9dJoLXB9ge6pk2Wq1U8I4mWGG5fb0Ip+s9V/Y75B1+r
WsRY7zNN3g62Wmz2SqoinlbKoEjJ/rtf3qC5Ygss9cEsmbcjkGm5ZGMeOcIK
x/3dN48oNuBSbfwb59U/Zo/GE7zhgTpIud8UXZnISk0eUc7KxHCzoI1h4vxu
x0y7euZsq0XYoCDL3QycCEdSUg08PdNkKApSwbW8CxylSLU7NriA/43JyX7I
oPEBKc4XiV81flz3Kbao1GPE30mW7+U1KN10oVXinVjRKCU23cNMOkxH++VH
ZPSsm7BCapr69hFl0+C2hH9lrYpwNfy+d4+dIu8zwSRGFzTa47gr8hMdKEf4
XfZBZl8RPiBgJg+RpMybUEikufEmoLV9JQ5EgqeZJS+zGWOEj3ZlWJJwtYRV
QLEoFvQBv+pcwdcVZvcY+0vm6+iz+Tbbyo1Rdl8TsvoumRy5/HVW1uXwYGXu
TBXUJ1fHUwjjP/WEilSIZ5UwiYNCFhhIIiwtzYjOUnBJQ/pHyzOqd1owcR+g
xfZAtDOb4LevvTBrDDpKU/pJyrM4U5PF/ekY0Tv9mU45oLJ0U1WzmtkgX/iH
bAyghaesbzpZiAlymk5lZKhy53nkozAOoFm0wyP8MI2ZgUBlqTcCWBHJfEh6
cj//OOMJdNOL3jQl83pXXKRw9M1/y3wwHcDPMTtQ/ZlKw0LrHZSU9sC+IH/o
sgkCe65NeHqgjXa0S6xxZShZ4IG36XqdEX41yIBYBFMhfd2ZA0WpRTq5TPJG
3uQZ65zgEbGgHmRxuPJT8YJ/H39ZN/GrRJmhw9xGrEncJg5oGO5pOdLSyMZF
m8v2t0UI9GV/vcM4AiZ6/Z5ae0/3wZKJ/+flnmZGywVZgctS36CRZIF5eZMC
kvzSF6A/4bkw4PIjAL+mIui+zglbq8V426QqSFsPPSqk9jnPeDflnvGyrH+d
dkwt+2LToWqbw8GnynqfFP1r4HyeElJUAxpexgBH61cKUUFdoFH/kzcejq2c
F7+2L1Drv5J06SSu8BMWbKdzhWCKmWavhS3KNPoXO5/8pVBcv3AO1tGMwm8p
6TQ7b27X2v3flCVd/yT3p1swnIk3pF2uY48Ev1cZg2SFNxcQR4hTp9d7bF8U
aWD85z9hP/ySIG+HYj2DgOQvp+tXAu0aBzw8KKrzh1kYF0WTDYRaRMWfX+p5
1mYg150U8WR7BUHqjzUTe5fyDsakvDlBSXaY7ih1G5RWE79CU4GfdDoaGgJN
nbJFWI4szJ45cr2KE3JaK+XKyzCHS5E0GwISLhMfy4UOqO4UCaYJSGFSnJf0
WEo5+JnVzG5lAupl1xR076BEtzxBY7ZjSR8vNy5WDi4U0o9w/k1X6OThu5ZE
2lx635YcV21w2PNhx52T7+L/vmrekA1sWN5vewvy3T1872K+8OHWb3EBGXJW
uii4oxssVscndanlq+KiWcRrz5jIRSWOUqaZj85nkaRNHSpSpxWfvn21SmSv
0A3AVGux2UaXjrF73V7Ibfl/WO+Kxhsf9nBpp8Ez64cLmb+g6cEonmMTOuPh
iQZCJe3e04MMNmZW/UcFKg+mUHHWSXm0YLlsDVjHJGvnjxcStmL68lodbIBx
lJ7Btd4duIMBPnvLH07dVvrQtyN/GtbFz2R0hrJZ746r9AeCqc0FkcYHG1MZ
LIV8w+CQVk2RM8665u08+4yfzbxjZUo+FTkSfRr2VIGMaybh+qbDDAQXqDMh
Y1GKp6sUVkUeDJmnxfljSteDFDfxuiqsZgAzCVUYJ6SnlPqWxsBnqaeoa6/s
H8C0znwhAxdvWfj9Omc+N8MpnEmPTtJi5BOugRBEkpBWVRvkxMGYkkkUZ2IF
hAznuYC7r/yZN4gveoIFhdWNeAKLa9npC9fa4UFOrAzuHPqx2pVBWQruHIDs
tE65a2Xp9Cnh/lZOTc/1rQEMR65uI0m0h2GfXfA1xxgCHJWaaFHq/jqNYcUd
yZ5GaECKaCB98EzbFJzImpFmK0tY5MFd7DwpiIQKdKoQxTz4Nqt3k7MWw9Ia
ve2i0xF3uKpSAWJVr/txbwIO5Dv0mI1fIG+fsZ+KTBBAsYxk04GIAbgA4dfB
dx2RBGHtdEaRC9m3w5u6bEwcxC41EaCRsguwvXqQCO4CwGXCkSfHTG6psBZy
2F7qJ0pLZkg5w4SjOquagyfKYvG8fMyqEUQDl4ljvMrEFXV0fVYWMZyjRw9u
JvVDhZCSh6ijWjlBWzn+HEUAQ71KipG+DOUm/qFHN4xeXXHhQT4J1eNkGO/i
55qXTFGaAQtZNfIaHWU6dLK/F5HeA3vb+9bUL6XOhPJL7hjBsCbtrG/BRhWW
fZjkdc70RIH0HaVtfrV8xengSv0ZWLGik8lUyaj6s8FzPB4s2FSCpMXz+6fc
dUCHNanoaAnBueL5kWa1lg5Z0P2wkpWNHfjZqdw1ouHIc27EoWVe22EBO8dx
2vauXSWuvM2x2xy/U3S+t+PWk4E80PAd8gOlOX0pUotFmXGtjSKwfJsDY1As
C25w8i1vmVFDIXS5PKnvPNMRd6fOOpaM+EKfIBrVpmvpk9ZErP4yubOQtIEW
fgxIq6dmpSTVScGMSuqxS1G5wG/lQlUrsUZ64axiuc/KFhSTfUZ9eerjFTx3
ZmERHmU+LwivOPO7SgJXC7u41OSvCrU/smvTF1UiXRegeRFh6y22nIRlNAXm
ccwiHW9LHPpQlzio72epga3G8dF42osJPvPiDUu7wqZBJfMOLeNKwWlHGcdb
CJDRLrN5zeGC1zap5nT5Fv6JZozth852z7ZP9WfoG4bzkO9QVXeQotNblFxC
hMCfT5j0fRvyNzf8HSfUeHr4wC3UO69xtrtdpCwoQZGTQAn9pNShkE+4HOdk
eF8msD7v2Q50Mofe4wyKmISNCHqiH1QX0sGyVnsiQLA8zhPU3UYpxGjvJCgT
gJHv26IdJ1yWDnvATpDvhjUIwIbKAj+z1SqJvFz8C6qYzVv/jT8ijqyxvv1n
NXK+fHhfxyBlIEGiEP/qVrwaAmG+LTW/fWZThSUZ/QZcaLUbEaM2Jf2KjhvV
K8aDlbwXEMbaIDbNb+qtw0IsJdHpbhEHRbD8vXW9lSBE+wUhps1gMuaQYBrs
Ej+/igFJC0q85e4xG82ADW6ZtjKKbPbpIrTxp9T17kLhK/1R1JSJs+MQ4olJ
VHOK85pIJEoMSkc7KEt7bJnjwWp3eASyURT+/Q80tMsu49wg1Mkd6GSYukKk
8VJDrSQMrfb+wcG+iz3hj91HZaj6jwTArFr9YRGzIVaeDOnpKfaMTPES/Uj2
WQsMwGOM3wd9lNvSwDUvAqZYlrxbEXXiE/qGK3NcinxHlMTt3fOeJQ60IOe2
44Q+AmlgptdIN1WIOErX59aOu2x93X3sy9ZgNZ08MR3gjuJMA5z7I/CUDWkF
4/P9oLXruJWqN2QVidzjkTXRyLBvlp/5dKg0Fe5Z9aNmRVsE+RwPCZmziQR2
salJHB2zqp2RRNMAsX3Jc1RAMVBU0cImQV+x7iSITtX9HQo3x/ac/PjQu+hz
y2HP8vhekkNeDO83Rntsmg7rddKpiuMFUfmOMtn4sGgkQV+o6LMYOdo7mwYX
KEBYfW8WpyxRWLC+nil1NIFCp5Ldk2a0XWrAkybIjE2JCL1nRFTJGlISFMph
RLjHn+H1kGm6cwaI+exQpK+C3H0sbb/q+cVjAP1jwQ5pNJSRgVatZugbHaHU
7GDb4fp0+cyrtk8ky6M//xrV+jRWHGwcUp6Lr0s5ASfN3N8n1uIBGxMuxtIu
o9+6pcW/hZmiaYXMrx/pdOED6bCY/lAW24duajKO/ogOoheSAzYfRpjOjKGK
EN9sn12wWP0GM4i/a1rP2hE8t1aFUvPLcI78gwb2WP0ouJZKC1PT+ufG0m3I
P9ZkyKdnoPEyJBavMFXaNBUIMfrXtxRg+EnRRQirEsS8ski0JQSM+4VnjxVm
KvRopYiBBjXE/D7ekxtYAkVtbLFSeYIp9QkASdWKGNUj226jIBdvzmVArsuY
1qpaFO6K/FAiZBy6DWrr4bMALh5TngewuVj3YhOCkbFXPCA7h8c+rOSaeun9
GddTj37mpd/R1uvgCh7d9PLqUZ52aqkxrJKQT3yVWalJu2NjPxWsC3PQjJY9
v1S0AzCsWO9/3ZL6Xl+qEsluO42+02w8AeEsDwimazFm4Col94NO02vzum53
wqFRdo8wLOLJU5UyCtXxlhHjo6cKzJTr4pygSkjwq9Y0U77eQrGHDgT3OwMx
nQ8E3xt7gcwubNLTSoUV9squTsGDeYTQmEpne7ov2uZMfNogN0G/iK4PwG45
iben/OANbdUI49LCGUKZ2btsC59sUajZIqiSA+dvNLOhNHrQSAyVtOH23tyg
5c1+81ud9ig+Jl/J9Xidr4NaoiUUz09ieZsPrcbXcOezE+xi+K9ofwRNaC5q
xk/qmtCqwkqdQaYXiJiAV0RL9iTCjkGCZrlt7GksUqDkmr+R2ebYtTb99mLX
1SQK0nW4PXW0lGQF4cMjmQg7hi5QqMPJWAsMzFx3kbH3eV5VVhXOehIotkTg
f3av8FxeZ1OuV5rbgrz7+yx6BJcs2LUW1g+Fe6ctQoKH9zXQ/xobpJ1l+iHm
jsO7zkqT5wZwRv9ecsThZWLoXxjLWQZLVHnbFpr78acCF41pSSoJgN+utxb8
wB34sVzZrwV6OgGmWfOdgQe8qK1Em7WaOwQuBc6vzn0wO+C6D1BzZwB0GvXO
Z+aCUNDBfo3aw6kWp2fS0gG1Jv+rAR2EQ4jP0D/PwKK1zcTBC4OKZLsYyZ+a
RvEBEFqGdxVQXiy8/LKYISVCQDa9pooW6aF9qFuC+v5xEcfzzz0G5WQ6BbQw
cgWssOKEIeAo5KaJdmL06HWelPcQfzQwwwEniu+OGu/VW/ImnwM3p1CpkuuV
Dz2mxnBXFIw25u4ZtmMEjgVJQdOFtZ9x5aQq/nda3MDUCTR3Mg5bmdDJOO9W
NXSWBP5D87tTkDls7klfsDSh3S8rwYKOen1BWPzTsHqGVeGgh7Un+KMklLzA
R/sg4uOxFrCp7fPtncGfWW3TZfo3M8W3j0kNi25yQraFpuUJtSK+/PAFqrKe
HKkGrxnmmHP/zxrvHtRTHLa2gy7BuN1zN9jGwP51hR+0mbQNHiKUfNbht0P1
7deESXMFY3wjf4TLg+dnk6AOCMtMvImtP4Qhgi1ASaZsJPYVugMxkug5dcpG
MFW16DnCsqbmzRgLniJhG+Yhh6yHpOljrAmySk0duDWFkSAh4uTQx4wB65/v
RXgNFNBeU29p7kwoQMcc7lPpORg6WSrCjM19+YMrtLHcNgM9zR2bm1DPNsFK
IqrhkAIynd2NMjVeETYqB9e0oic05N/izVQqGhwL++7xFw3g8NZYmOJ1nhqv
cl5TH6j0+wzN/c+rMg7P72/olhy3AgJLll5AanmFIwFhaOS4uHEZkg/1wEtl
MJ2U/fBE/3ZiSYWF+pOICZMZCmudQGiPV9emAph7sB/dZgqJAFTPkf8LGQSw
Dm5tNJI5QDln9XptEZFxxt7dg15ncgPWOVrOFPgkPT0Wz/YfIgHyvutit7+h
L4+ylzIaHD5T5rJip561j8UFtNHp36NMpIBiEOO7ol8VjCH4A9sGhRFE7xot
KgBzUMQgkFCWmSrZhaiLHvQlgGN1AWW75bIJF/MnSIgrmzRSsagBqwEDCofQ
v0SObMPXIxd0Dbe/gVOlYcgzIKG7hCYdxyNru+hce1ZA2rssYI5K6Ty+dF58
4ig9t10+SPu2XzaiaKqKuoaooUPXn4+1v34eARgAjsUlGPB8b/VLrwQVdkXd
7AkJydtiyiiSKe7fGc41OWgkBSWQYlJB247PwL4/MKxdtiJTn32vmeQuT84y
zpiiTDpDL6U/45lnNy88pppC6+RNRvVh4dnE1+HsF7vQ+ys9W/CWk4QQdpTM
1dVo9c8L/PZoSFm3RvdDgdHD5g6HdKNtIN2PuYPTjpeQ4iKaWutFhGzuOhJ5
Wj8ulp1KRtvL7QwX6amQPeufZF7YLXw4iPHpoyTsYBBqyqMGoMm+mM5hbnRW
98TmS6s74s4nhn4kP14zdX+FrbccaqLwQCdF+8v2CY04nurTBtCOuWmAJ9Ux
6bIIE2KCd10zK7k4LYYD1pHZugRZ1AcHad3YbLQq27F+axpea/lKQQc0f6zk
u3Z1XEm7S/F8ImfI+PhSETznwbv/R03G8Vv8g6+OvlIu8FGnzcdLJwbcbWar
PT30l13yv5zX6jwX5U5c/TsHIEqtLMt6M+H4ND0gDinhc8s4VgntYvjj5MOn
ckSalkGBZ1s7vkjrHmq7XkKbjbwCvmH0R4CzQG/XSfHty4Xzm4oe3h6VQRte
9oXqLjnMms59/1qrFQLHJclm6CVOLYdzNYH7PxIkXuUqW2+Gxp3cbBej4eZO
0IdF+kJMAr01/i2z1+W3HJ8nKFnutFEFOGInhQv0g/NFaOrh/Vb8Md6gvI8i
SZT62o5cwgx/OFYtmWwDcHZ3yZZXThG9l9xqDU1Sx6D6ZuqUIJ3F52PfhApr
C10cyWbwRnoSXUNUQF87RC6cAEhJR3iDh9APY/g8dDTdY/nlvntNdltRxrXQ
3YdOilMq0gTHarnscrZpHjownKEkvYm0SKqaTz5H4teibZ84N9/RKIcgAMab
qjtLHO+B/4nwNnx4E4IFyrPCupje3QXgKgggbYzgkfyEippyPyCsrmCGwN3I
6Yif4UtPu5I4pvktj8XkpV3zSDJSyfCvYIdmnrR7PvbSg2uoIcZjOUKj/OED
P1WhKCbTtlOfE7sikZVOmvcmTDj8ZGqGYxe5ayYAZWxJswU/itoqs0tLtXEZ
UoajBUsKVrZgd4DCh/tkETEkBAKbE8jEukoRspNFhxczsNUyt/EKtpwRjKkk
RmUn5SV0Pf0ygXaiuRNjYoms2IthpNHPciTurU8R3d6QG7WUe5Gu5CuKgmfu
xUIup1kQoSPMPGS1VMEwTa6zsYOF6pq72gX1GVuLRom8pevfuYrhzUWdR3jB
g23feu7k/RjfWFJPs3dOH5H5P9KlviUi8fLtWu6AvMGYJRupt6WhiIlPPi+p
XDRJ+/QO/pkG/aFnYEV9v1aun+tfF6AuZ/p+xSbw+My5tNyUlmLfoqZ+Ag+I
kV7eY/b0+0YlybziidgmzmjCHka0xaxOie9qZHhzbg2GbgAXycGrlhbU74dC
vf6uNwpfNzj73mZ6cruw5qGrtKlqSl8+uvOGbAPxiABF2kadOSaHNpUHk8yM
JqH0jFVl92uDWu83eCLzbg+yOsubgBzKvogLTl+D+OYmVM5JkTOFm5WnBb08
BkxRzBhyOmAWm4ibEGSyeG5V248v4zF4EaU/swfoXtb7eXkjbX4hjhcOZL9m
ECXQohbj4D4yHNMBvJ1JXOckdsQUV4CEgrgm568PVufVbqx++Y2Q0Sc2Ys7y
tFl+6THKyG7U24MttEt6TSLO3HdRhJlRfIsdLcO1skEpLlCC7hZjAFDQyeR4
dNL0vbL2zE7DqkIJBWBCnpE10wBWUuMsanPGT8N/SIvzgEzpnEI0Don9OiY9
rRdJDAZ26f/MT984m1HM6QSLKfxrOcb78PjQkLhbLucnpLi+lgcUuoDUjt2/
hCdlMdp9rs3ej1vz+iIEneEhcdAtbBLtKLT3NT05xmYofcjNPEdI07oEHQGu
rI0ZjEeLsW4rVa/61+pCKo+h54CWwvHi9aTrswJm1rwlrTsKoLUnyfXKxP3m
EkZvkK6TtVhlCcHv+bmM/u+IMH8Ufrihd4VuFjpFnAUkE5bd6iojkRK0pZ5E
SXPzxVSa3ZCeSU20UHnJ3u5OGTirB2g2Z6CL/tBO/JjnTLFiO881QV5cAyZk
F+k5ew3Je5WsoeVarIIdhm4c3hZMNQiYQuDoGIuBX7+M9dHiLIhl6lbARxfQ
NB93iSeJ92HBAGYLtyStyASG8/tKCtw8BPn8HXwv/70Rp70KB6Pyc+daVY/l
SHe4wcGFHM0cF3+/KczKGjhpicncRn+YvZWENmty6wuZO0jqR9RvH8z/XaAv
j7IecNepLJmCc9CroYAR9ig9EPnkrsC9SMLEn+TEloYCQbNtjzer0DaQEGfS
Cpu9afaoAUJuR9zy6ZUtq7xWx0mQFiTvhOfb1zqqMsMW04gpcE0MIGLf9esm
muvccXN4SC1FuuYqFi67lquWP974Ax9IjgEbRxhhnQT+N0sDbCIyprG6Hhj7
ILsCtB/whoNAmn1RMl8C+0ky5bs5hQIY1+x3v6j24i9zvKvNYlLSeWKU7LMC
+V7mdDkyfyhMoRoE++J5bEB09D8um3CXGemASYFgjfubO0OniMWMNSQK2o+g
tVMwtuGMvPxrOMdEWZw7AO0UMQmmhn144mkgoYX6X9jIcCb4FLd7iaQsVdrt
c47IsyiFh/wA13s/+xyY6IRyXW2itGEHwib9V9e9nmJUz7bVBE5wrkRRE8/N
jTHl8PVgl6oB5knYYtrC1/6CTuzGcfdvgdlZR9AVY+clKx1aSUgoeQUnhyuI
wuzKhF+gZQXFdTsI+ndj4+GvN4GpQCQICpDHCrjcBIB4zvqocxuw04xUMSTw
v2DGLbvVHlBDsJTHf0zBaNgqAFIYaEn+BAU4VkZkPaC85R7PkXKxfKrJbEXA
OWzXXlwk+ucj+ue0YQJiGXgJP0VOzWPPdn4dKP1XWe3jd5HnDd6a0Mr1VMhk
RjoR8Bq9Nz29minwzo5m25pihnNpg2MMFjUo6HRfQOyUA9NtoyeAwxhLTLBg
HPvLRyvoEM9XDCnBuMlg8JC0ZdySyhkBTNLGkkZj9Zr2A6YKygXe86qcop8O
YAX/eBGsq7A7SZZxyS4uUbdUodkaaxkNPJqQTCuAtme5osByghO+iAW8dHlQ
mOp+ovlGRhpi5CmAlV/Z14qeUlPh7R+orViGZt9zmy5LRPsZDy9krJcuPYAv
MlWq4QPq3ikTZabAi1JwcpEeRo3r347SG7ztfMsPtVBExO7tQyhBmTCHXgjD
R9sOsra91Xdcw8y8jLmS3Nf1brxkwytN1GOhTlsd8kUubzyJjYVjIweNin65
FcHEgmqeumOXggiqWheViJtoF3+YtqUt+u0a5xai3qmvdd2wpeOUGzpCDQdW
LetSTIYPuevm1pi91jPoyAjTXKax7nVJR7Zzyor0g9PaCdsvtv2xeIGw0tdC
4gjDDrYDuaDnQleJ1sByQMss5kLFpuClxdaTHo3d9T68p2DbnLlgUApDSf7m
DasWzmbYUxoe0bro/iFH6RszsK09JsGw9lfVhhu77fQCUULMEzf5XRtDmIJk
lU8Z6qMYgqgf9WEHjIVUBK55xWKtuzdD5EYs78sMstCYQsRlhhR63QTEitJ3
M1Be3rkUVE0c/E8/Mw4xSJxrj3tYLIkUC5kL1/FvtOno92M+wm4OH1WuL4n6
6SZiZVkdtEZdn+pB0YBmQ8uyC6N7PvLGUA/f8VNdQBD4TWQP28ipzOHQHxY+
4TTjlQsrpOZ/7q3lh0sCav7NG5EtYAfjSu4LX1ybrAN90D8RffQgc1DvGlOB
WuAFSRS0oIfiVrd7gelbhu5csDdTxn/JWokwGKIdNI0A54m+TN/Df9q1ziQe
rkcZeevahvsdnfbWeiK1fMMn0L7CF2zV6QFUXISK/yldWzd5KEG06shi2JXT
aMF7vI0RO4eqU2nA6nK28Ufx09vam2Iw4HFGoqAFtfclGh6eYixbRf/iu4re
hOeOX16UmXVkdXxrHmrb1lEieQCKiV8E0MC4K3ng6n4zuDMS8L4MCn2L6euc
jyHuZj+OekWbu3sVzD4mZCqe+gMskl8HoSK7Ek/2SWA/ALZnxIuULvZBC6lH
ML2ib5x+zGs9eS31nmlJdUe78P6bVpY9P6M3Vnl8uBuecOcdoHO4YDoEXMzt
DIUiUDJqzd0w5ueMTQig8wPaCf5PSUIXvAJOK4d8hrmsEUQQRw+SlEsaVgIl
wH3sd/xQygklUs01e34UgbX+FmRxzU+gcxy5RTgpi9acGgJNYz3Yj4JA/QZM
I2pEiKgwgq/Pje/W3jfysWpk88XcNf48KBPZcMekhBAlfQ9F4qsbKwdz2iKg
OIphLBVRTmDHVkvKJVA+xYmzI7hW1h5aXV7T6Yl3Uah1AFYnbOLgUR6gMlig
2VYJJaHaM27EDnOXNUjkA/wSlVzO+uVyJv68kfhzK2nl57zi2boECJqrd+gY
1xuv4rqs+9cbts2xuKV3nl1fjEownwugcDeE8YBh5tlNhJ7a1QkU1KNT/pUF
zNH2mcVHzToCkq3ere7KHJs7gPIJBZhaP6piXRUirTdy0q2BxUeDcNmm2arm
onQS9iChPoKTudnXDWW7Oeh8uIU/hCAKYN2lai30GdidHF7G76ywRDKS8yRD
7sdU9kUj/uuEcw9JsepCIO7nEdFYLtVdDkB+vOzRx+LY+sOZ4ango+G82XsT
3At9SExl7Y3awlkiDugPqOfEclmH9gp8HvKeRehPC1jSgT0bWVLowtszg2Zc
3gmTXFFYcVa7BCZFju7sihVzaU7IEscJajfSvt8VLrXeReR6yo/mQeHsg4Jj
HJjEkfXUoNwRvLjewgXj1w7wxv1D4kbutudZAFZcpSX98b8L+NAXqehnuuWg
n+wqrxVOmTmbv+9MGsyS08uvE2H8RVndDyAXj6nUQp0+V+DDYlc8gFwbgG5i
4HxZgQ9ebgMbpts1xkeWAFVdH8+7vz0liPM540av93wPHAnnCZ5pzChcQGD+
5Vem3lI5P8VF+ISn1YG//f3CpH2cxZTgOgLHcuSHqYJmMSO6iwEiScfsxM76
HRuGeOwyt2R/LJ9Cei2xj1gC9fqN1Fo9YqTLrqPBwF7e4E5glPYQOJg0DAup
ZuBYPUE/mv7nUe9zMjXC3HIJjQlPEO7T4P608e1ToqCuXbxozLlzlyL/ksYc
tk8U1acsuU8eZxXUgCOct7W7tQK3VyZVagpIiFXXKb8oPMmVfa3E7tecNR86
r7w/dOCAZScD4hPKzfipOK2bXinFwBgN+t2lxsyXrrYe2EgmQlgp1O8zh5Im
yPIQIdEwOuccJHnAE6opij5BJ8syaj9y2soDl3JaVQ0NrSp0Paz05jyd/Vj3
VoX+IXuKLcbVRsOJSmyjw805hFSg6LYe4EMf0mRONNvoGJqpfx+SFGiFy4oH
X07iNN3v5QXU5DzCt5wwBdUsk8Qh+Oe+Erm4fyvVRmledZzKdmfMCn4/IBOR
ur9XyJpEFqdFkAgJYCGqGMecIM7RhMDv4n5cUcWNQFF0uky70BEicxcOH0Tv
yAqTst4BXX8DE5L+vz3Wa2atQTrGEBoVDCrgUfk9aJCpc1pSebP/zn4EqBUQ
krSnoFdlVx8A4EYzAgI9/MhSVS1U00CxcS0UyreuIIBYh9KN1yKmXN7oZuqP
YYKrsNIQEVSbio8owhy5mlG4IammIT5w73iiHsmkYO8zmS/qVboxpx7KwmJm
VQ4vqCbBZIe8bTWyGERri7me375BrR6CRnVCavDd4u7CzEXNFNp5XOCKG/Qb
2eOpk5uU9j3BnkRkPh28gdjpt0Obj1ogvrXtNDbvLqbmyscB1o8m+Fq5pQpi
xhovWRFGN8Gpbbe+EvaWXyUSXuOl+vVLLY1Snp4lIgNqoeB5p4nPS+0P4u5k
JYIbYwHvVmeocltfboJZXfb+r0dVootY4Q9cRjd4wNNjvvq+tjnM1neKpBhE
Rhii/koNRpQx0htWAMLl+9Jj2q84DV6YbsdmedymV8w48ZOg1kgbvQHXCUGL
aLSbIshWUt2a75ll2TvkOK8C3otj5EgEF+mkZDcdqvXY4FxhHYeFDCkDfDpo
Bwjaq42JflbLOjCRLQKlwXrUnt3NC5f2Vx8KXMwePLbnQJ1UYXsyWLvA3MGX
ZSXx0WYysAkGxsIcB+OOtX0jXKPVKIeN4E8tlupJDq27xg0p/lLy93wG0vca
PiEczssFWv76k69VP/sOa6IOMUabO8Ezi4OE8fqqNri3Epy4vfp7+uALCcGP
PB5YZZaebff5Z322mf0N8gmhwTenCaFvVgZu/Ymm3ZSbGMZJ4dkkZb6WLhDQ
J6TpJ1v0s6BY0txkfTCwVZa3t785Jtu7j4AJTKNXN7JahTkZ7vVmS0kDCyVQ
iHJLap8/Prux9DHVUnoUr6+V7bOKacKHCCReYHFXGDlycGxlefvs56vZTwC/
uKN8ZWcveevJB7flQaywZVt6LvDZfRt7xos0w/pCI1HdHuLebfvHyy+t5nrR
+JJ5ICCW/4TMvKE8WjbJkjrhs1nvaY4y+FH3vQK4R+0y8wCKVhg2JOkTWOCo
CA7+HtavqowV63bV/t1HwuZkF3IgnM0XGOSCi72PbM8XieGnkTOqDUOW8uSU
RcM3Y5lJ0Gj47p4mpjMSkZmXlJMUHGTnGuaM+hhx16xG5UnxKwXI4TJGypMx
veagAylSSjDSk4tdwZs52w2RpY7xErw9zilr/XnOAyBdGvBCvSlhrkgVzj49
XvbEvf+BWjJR6atKBLFfC3vVw9JiVpHBG7i8EK20O8GCHPSzjsxYsZcBy4Rg
MSIxkXFsab04GprQq3mBUl2sGzKH3NeyzQYHNWa4s9edzl1ZGRdkVvPa1l8M
tn6+UoLSy/VNbR21HFt8lldriTNhGL+0j3YAVRLSzKv8PKz3krdeX1N0sGJm
iFs0TL9EtTvJXgaz6CZhVWrcd7KdFGVHsO2bOAbcy0497JzWJ/ZqPSXmLAV9
w6/EMYCH0qQYlaW0Prm44phZhSAoSIycMTRruxUDyBx/QbaymhJTHZ7cqKRI
n5KJZPcvnYQEajak82i02S1fq3xvdZ3wIyTh1RtxuBrT14j7nWkdnpXgNKZG
VovR6k9nykCDGsUYspPAJdReph/f9YSnBx6ojdzmyUGoKPDrxxgQchDWyoaA
tv34TAqkO85jAyZ2WA3fEQj0sIO/CHcfSDl8ybS6AwfmDoqt3oHEaMBHf759
eEMJGFZIH+oiv+oV6AooWCrpkvN/SpsNYddNvRF/0+PjEU7T1mkaZzE3fStN
fqab24LhHkRxahQiKXTcjBmk9kLUvseeMKCVeAZosNT30lavBa3UjuD70aPC
yQgiYXV7FmVzAUxEbYOwmPts3W5fSnaUGMQufdIr3KhcPWxkjlbhYszHoyxY
qkORDkdLLqVbFJn+B01NazrJcUrfqPhciR4Wh/CYVIzpY7Cr9OEtG7jWfAyz
4WVWqnowPQ9k1vXghYS0o6Lu4eOPPJOJKhS79JM9wTIVzBJCmlymI92c/btv
Ekl49uWPbVy1v6bprRzwlwkLTrjT7B0ApHzptpm2AZkSiT86x9EcDiJjISKB
9UVYYpkijw71BZCmkOhx53IXjPdRphARtelY5OW0Z3Dx8KTfLkhSdZzlgVVB
z00Hv3MH5KLOCUM2cXooNVt0jTTHexu1H9P6Sqjr3VqL6ouTSu5psfFw3L0W
UTZTI3fw5ax34qYxFEpS4HWLOVGch4/58ldGgJJ3MpOldc5v7aq7SIJkkyXS
54GRrlfAAIqcn6A8Q0WXiBv0CAji4/dSVpPWK4aVFGGtt+LPHK+4ZC1bZ1R2
rDVJQ87sNGr8+cvr8RxBrRSUTUOC9NrwISe0Fkbeunrejla9f0rrjJyYavtM
F8yu0MH7T9znTNtxcVatAHWmDhHgfhmM6ANFs3AQJ0bEhcUwxJJ49eSQfFAo
EgVCRPfLhWRF8jJXGKrHlJThPQEJCLTqYhR9/eKnHsK9/+GTQl0xsoKzZUoX
gjkng+a+VRngIh90ieMwnL+6mwGzZb/nbEEr5BIrdISrSp3UH9l5bYnn2rEH
C1RSgGh9TMlwol03PHzPBdFqb9kuBWpHBIGjQaURAddTPqNdb2cXjAazcadv
A9F7nTUMXpel6x+EZxNsrMgY2PtvsQiGT4PsSmuwB0svZ+Z0439xS/3Uahxk
uT74gc4z/vPNAs6zKICXD+Bq+sFJnt3cpqDPghNhuaBK6OHAFGwQ0be4b+xc
GDkz+psToMn3E0yX3ivK9fmosH7trPB9bRRJ2En8hCvINHrOQtFVADo14jku
wkmMcrxkUcrP4uSmq+U6Ek6w3eSX/bDHkM0ygFsDoM8BdFFP3X7WEeaKe9zh
LUGS9EWHrVe+u5ijpEoF7SL4U3CpUmjEo1xxYg+fVnygALxoven8L14CWlA3
XJBwWejxfySWYtA1/K/E1Yrs88ddcEpLUGGX7kOf4yJQjwUPaLCz6mbtkpEg
jaaGbiZyVzjSRuTsYseDYnlwsR7CYtqSpE771vFdmC9Bq24AH8mVmEWr9s1m
ipifJmv34jzvxIhpZHuwChMoR2jj7/LiJ/dAx2VW5gIIeVXqw1X8n3QrlSfT
oDNs1FIJWpNKNzNAXH8H374T3yoAhncB3zbwN6iZXA+jyA3pC4GWMvBxgI9g
okV50o1dwi+uCI1blWEs7PWAK2xwT9o7fperOkNQc4t6TM0oOZwWPQFZkzB3
N4Ph0zzlJcznTJxmXls2xEuqZZw/dfo8ZSfvgxxoBjjvjd6ToWZR7vXZRmt1
S/oDOfOku52iBXVx1OczBhEX4WJ0kzUH382GLQb7YYZsd6dD1g0gNspHdNqe
BkEeuRGud7Zrb19ir2nQejBY0vhMDbLgW7Jpsh5ai2IJFbfNwm1psbSpY78I
QnMJb4CPmaCxjTLn23wbV/EtwG6Xjmkk4xB++nGsAuzq+y0EY+aTuEyq3E/b
2R/QwBPnx+QV5yxxw+69T47zKk4nBVYI/BT5V7ojB0pleSI2WR2YG2REQ+NP
MTVb1wLdGyaV1yldS4KrrX92Xc8ndlahuTIDK+HNt65BvTuEU0tGsE7y53D3
8MIDH6c7hUSBaNJKI1K488cMmQMiC39dMHudllvtDFJuLUz63rgNItDJFR5E
gw74t0M3JOs2r62/NzWU1hekS6oJl5AdfpQ/kHkoW1i7xywwdATjYa2S4VUf
QHLBVm1KLXEaFKHTdEp/rIqsmtoV5mKv+RpYnvV9VFhiNdoazTJLBvb8CN+f
tSyXZrrBDG6SC/mshqlFSai8ys9Lwm8o7NyMY+Z0tl+dOz4vTwS0pbGbCejA
+7UhtzQysuqgdoIEmkp+N9xqNBoV9Van9+Y5xYdwBPqIF61pJDWpfic1NQa9
WkIDY6jlbGkiLgjIkPZdidHA1S5RvgJO7jpZey9NnRJgNhGtZOzpXw3FBLtK
+gAGv+Vva7Pl3OtAZTp5W8RKLXfgzhxBsAkU4YqVO4R63gfr+RWasGFyFRRt
WixMtPnvvMAmMzBIUZQbBM5SqjRZqIcGAylOtWqEVo0Ch95tLVls1HtlrQUZ
QFIyWcqlh3tNYpbFlAGFQSdgfkxvh1cSeuH8AP0naoFHzFu+biq2ni/+hvIn
WQbHFP2KiO0We5CtVfiGfLId5TPdquVkI4ObGs0wHMKldQ1e4ExOBfoPV5Jk
hCYtejK3qOBflryjlJOhalkzV1t8tLxlMIJHg7p5i/UcO0RBuShsDtymtyB5
U/fmXZ9yc1xJItHobDps3bhB1APCvRleLTMw+0EOeHLtP3MEx9faICYB88La
QvKTlt9NUf27lcUhURewUp0BH9PFmngqOr+fy5JU3G00n3nD2R0Nsrakraa4
BlDbHlk5YXI2yzODS9gUpqPKFbhaMzTUO94LN5iBBjfKXZ5dMynndNAHdula
BK5gB3bgNptwpsoaoZkbcZRJTmtD3kATURTvoXcCydATZP1SS1IK6QkK47uV
sn40aq8/ucB6lImDufQjWNjEAx7mCM6q14vQvfS7IL9/aL+La8EyhvQnMvnj
R2qsdmDUkMp5tcilD6X4NY4Pxtju+fpJuPzXYoHaYkxQIV2qnJ/cO3ndSmyQ
oI6IpMAI32n8lOSFXDzKBhFt46AvZlKoh2rzOp0pFCPRBTViLUT3Bsd30sKT
E0iqjwOMUPW2GGiuLT8FuGt3Tz+pl10CMSsSP5PCNOP6PfTqY4eHj0OQlDa+
NjXEOrDhypCmY4HJQOiN8x8vzuIBGO3FfbaQEROzrJcjZsIHpI2LGjHu206s
stSfQ1oX0yOQL8lfqmbz3jo6EaEWwetuN+03LwC2JYN3g5qV8m990wDv2lSx
CIDORbYNIeMUTQAFxNN87w2+yGnJp8eqIjM69WrcIroweaOrnw2TmuWI1EMN
mCDQH1veG8CQb/QbuoJvl80VMU1623naLJ5DFUqaalmKmppPlVvgg+TRTnJK
gai0I+M9MeLiGDxOc1XuEeTnDOmUyzgWL+kEHnOwJ2wXM9xlfC5egkDor2WF
OFlxuDCQelWC2edJu1+Hkucqtg6bcTHd9V1hup9x1LO40NtEOnoz4C4rPHOa
qG2v1zekiKP/sskMejFETlOBcO4ixbCmxRVdCxqqeHh8P5iDJ6fZmaFSKjDW
q0XSf8MS8xxfW3g2zFlBhOEazPTrQ27rLvnWRoMLLThuUJjpfUBHqeDiBebA
883aG6zhwRSXs4XQwCLusttiapY7uw0uhmHPg6Qa29jdEqOqTORBYiqAnpLt
1MbFLMQn9aZc6Pt5r0t2NuQjNmgdQohGJFmgXxxJ5rScyCXeD2KLW52LMA0n
Dy/0m5G/5SwqGJ9Yj6UVJvgwizzApQ3TK+2jf7l0lOkUioDtm1NtiSU9cJ0U
yFXnJa2PlOwBZN26Y6S6RJ+o92vjI3cTxJSCjZyunaWe9MSA+suV4xeo3IL6
7QIC9BFnap8OCfdqhSZCc7OlDZ9KKPuSEfWDqJRmqlQjT7A43xbEUbDjf+bJ
/vaRlTKJxbPLHENN46j45l69gr543JCGP3E3jz+q+ElKRpECC8jLjkxYcxnT
uHQ5ODvSP8TacaoRmWSCry13bzqD/vEqa3GnHYVQOKeeNg8UF7J/L7spxBAX
PYygrwjCSHXXV9rb3+eh2swjJ0W4xK4ysQrU8FztXST0xIoArN98frnAvrAI
e64e6VAoiVysXNxJbotD+88WN9NJCkgE4kpt62Y1285BikxhNOm0bfiYYa6i
fPXOND216l6puWJiYjd6lRARmnZ11z49YSot8WehJR9B5z6WH69J5Dlyiz7m
VzMUUA90M+1gpjNDTjM79eOcwiFoyKlQvGVFzK34TCU/zVsvfp36bhCaDTsN
XTQ2egUIHrT7wZ+8Q3Q7oJs88+P65Gp+oF0Bk8ciY9zwkFM/BpbBbxWlU6ue
rPleGdzygnlG+EozeTio+vbL7jcO/PSRugaITuydq3JBKq14LHiHquJu/tvE
+M3Q7+TY80GlryaBv7GMW+4STA2mfblawMDAY6v1510H5j+i5mJtvrj4s1R5
Ku5HisGT4G0ahJDxS4Voz7xBBln3JKo2dwZSwO5JHZe5JssMF0bM8vZtvs/6
cUE2mZlAb9t4ZJ+6Wo5Y+Ajkr8l+rl+GVLBvLthYd+nsj/wFcCxBuwZm7rNQ
VaHds8Iclq878L7b8WSm2KkiEbDuRcsUCaMUnDyewLJFMr0tsVPv3/EGaJCF
JWEWc1JlfPxzHhf+iNDZoxs30Xmsqt29qNlAaKtrr7KGXM5KsKZydZH3SiUb
iPY0WiRygr0yUEQNgLgQAkCpeWRIIXCXLuDK/5RB34VeoUQbAo3HVApg74ZN
tqOYDGKpe+u4YPZ9EsJFKYcJYA7nYyPLdHlqKFvkudWtDxYNazmMsXKTGNh5
zIRj7jdLZQEm0MaMjprSvVXyMkqgbWjEhwaEJFPPOJzzz/no9m7iUGJiwIOE
DzXjFT6G/YaGa51aa8txWBO6+2R3G4C6FeUdkXaXFMyNeZCJcf1O2k3F0L7e
gfKFycUccgltg3BdHuuX+2VfN/lnlZEdnY4BAPrxPc+AR/ifHYrYUUTeqlbX
z3UPR8nCfaoV93aNIHkxoZIO2eGNmBzf0AyVmVCrGzGT54+K2RuH+YEH/UAm
/yM/ZG2sf9KXvfi02BWTUcewtkEYAyEQzLRn7LRmbRYfZzdcf3B709w8RdjI
IAvO6gqzTetTMQ2JpNyhTTHiqOw0Rm2ecZmqJYK4UtVPvDPmuedhAIHkqB1g
rTyM7G3+uosHgB4FnJyNQ5hdP2cmHTVCAsxR/LkYcHCNtJ5H83t8ek8HkqbC
QMCLYgpSTAek4gVHD1DaPZFJewVXOZ/XGySTq800/FgegB8106iYu2A1u5Wg
mo3LgN26DuS2i7ZSIadbiridCO4lRduPCuO6ZFvXQvuFssxBWSMqs0TyNlNM
mkHLC5BZwuquVeNwVx83ir6yI90X08X6MY/b7OzuaZ10uNLQxhhUqN5gZw9/
2tMVTO51YMgsgT8eLLYsKD0/oNPbIGgusZU08OyZpnOS0w/QrY6B8kShKyVb
4PvCfgDI5uAmaRYCMXRXsr3cfefHwtZNslycW9zxhlxf/PIZ5rWaAOTeNSGt
vv4EYoa6/v/RgTgEtHA1htoosy8+rnwAo/FZEfoeNgxOob3lQ+wOASVT2U6r
TM8yyigvjX04vdOyQIXxDvFCc+SIhXFPa5YBDPYezJOqSYzo5sAfKu/+5Rj4
hRY4DnwW5PEhUSOAfpMz3HHiP5Ps6ulFlnNr+mlEaKm/QyyDzvt51ZeWsRM6
PQPzRdAiTtoaZkll5OXnBOWd6pI6bTj6jQ2zWMqMtqsb47sP63A9px5I92C6
1b0ZYit9tWP7Iq/lTM2QE0ozqTEzxLe9SJGeuoU2GJnVdpa6uPopWc2TYrlS
kbFOrYsGk/381cQv0dT6WBPtQkkPACCg6u38qN4PoT6LXQL2enC8hLDbizXW
4LNg2ANXjKyzdbBO0d6flnDTdlrbPSi0PVfRdIk5g+DRCW/JVfS3NveK+ZaV
HG2iQI9mvFHEWPoFB071pp0UYgo6dp+CxW+HCwX3hieQURy4e/eJ1U0hj3Um
KswzdCeohWKExFNZbBn71nDycU8T5809RKwH6Zt+7L60oju1WLf4aYv0a7UA
VOkOZcm3lTeBUfqiBOMigR9l3TtPI1aPrpOPnPubGT4KmMoYUMrflh4jBh8+
/WpgR4X2vS/fl7IMIplNL2JNOpfhxRctLhszg4Z9CQ83UTIMQ4R+hVVPzEO5
b1jWq+cO+UTc3tME4y10hJXG8d1dcC8muuYNImUKQu0X9p+0D9MFcsi9LXad
sSIc2nsR49yE5EERxrxLx5Kr1L+RN7jSEYFeoAsHV9nS5y63NDAUviFYL6Ua
jjrjGO6VL+RJJGyyx+D7qTbBP08K1IYCI843PZcZdz2cBqQJiF3RBglYwr0T
sdq1pko79hZsP3J65q915StVKP3Aao5KwDuIVeUjT8f+hHbYg0YAPr4Iqqml
Zl2cJorquwSGu/EYLGZ26BFjqB7N+CQswNBqgAOEFeltB7+ZfjN1A8c9Ad2v
RZ8wi7xJs06j1nRVB2zhKoBF5m4POL/h5NWr0dPAayEA8tkjf9Tl5wNb2zZU
jXu/WLnCJJfdGf7vvB9sH3kplvnzdrwLV6hZcFyLIZSH1Ip8xus6I0ESkh8B
rBlrUlLmLRjQkOPUQbjY7grT5TQY2ZcKmphFH67DJz76Uo1mfcJ4EGx1bmlH
dbqlANcvbLzSIQ4i116fgUPOkRxdlppx0Yuzcb0n9mST1MiQVJJ3JIjqMRjk
ew0VR57OoC8bZdCvxCpk6DahMdvJ+/5OWQonrcYGeYRPTuSOCqPxnCG6IL7Z
bOlUZ+X0b1WkXzFFmPHKlDMuhFr/o8iu+NTpfbvp3Nkgzkti1vZcB4WfFrDe
T5V0y6xb0e2pnkeSCQrDN2bNbZD8bchoTonhLtkPMCsS7CHLEyYQsV7jTrgl
/KqQKXaXBj4GMltkjas5EhbFsk87HbHTAHgmVBW2EWhvg4YeMTmebme+MKr8
E3qxxNwV2/8MZMh94kOre/yUfnNIFXmMyJsMqm+tlLXRLEWwbqf5os9B11MW
mWh5T9aA+q6R45pYFpZybPw7D6hHSwjhtHs5Y56EladB/ZX1bo22fPmaio0e
ZrUZY7u/JovfHELvW+J6T9ZzPNkMle1PufjV5h71Z5M96R5F0i0zghCRhqrR
JuHIFM8qnzH76fiDS+EGWhC1t5+AJdWUDPNRzrU/J+phk7fIXr0qb6NF670V
vPP8HZ/cMlrYbPVoTAV4HHV+K3yBSoeaN6qhdL8+TROwn7uMzGUIf5ExXBf4
KDX1kOWLONs8j6iEReqdOSTRCcFak80inAgtYQ/45kJlWZU5K8p5MuKnw6Yy
OcrJQItRLH/0bdoHi71NA/0bXRjFZWpbWKa9ZoKRhLkXEXxhCMHGG5XVQ+yg
U+EZAcqLC6wrFQP9KEOSDUBl1YnUzBYoMdCHD0AAwaYiOS3sXjtNZFCQSMQ6
c3OAeWgNLdjuI9ucmxqo94+QrGLL9OvCNQCrHwMhx8JAakNkIcw+A28JMImY
zf0ici+njQFjMM9tIG0kW1zokPPflgHaSO14H0c+3xm8K7cYOCMKXD5PXXYB
UJGHXp0C7Re0xWeF6MTDIWPn34QRY9ySOsTMGcMMiD101rbZ+Lfg2n816YU2
KHeSeDQH9UrzSmykX1gk071paKaY6R57JzfrgTbH0F/hYltN1IR+AU16w0HJ
Bbi6HqLEDWGtuMx337BrUrQmr9mAh52rzyXA+9BaTUKMSjNKpItbFqvR48S/
kauYpQ73k73bMNnVdYtODtfrK6WEZyfayYra7/Ami60WaYIR4Uq6sirYpfiJ
jx3ajN7vY1y7Hs3I1Q6MeUSeX4CTGL8+sTOYDF/E5PMGJtpZLRyNXV9+IwJ9
wfdLP4dWDxAh79nSU9dAwI+RnH0gFU1i/vkcFxfgZ2RlB5sT1zrl9Z4Ldr1O
4fDb0tpMLK6A77j5WnpzA3nCJ0GgcqjaHwZI3vIznHBJxeDD4AxovE6Num1x
wmTgz1L0/GKbb9IOgn7b0IF3hFzEcja4V0bwl27rVcHnN785WIqmbK1N9Uv1
kPVHIpNe4ZxKX1ANm0syQ82bhf/ohdtCpwn1VDPEwOtFYZlIbqooSD1Bw+xK
7pNQizXixr19+QOTNnGEkTrhJjja+7us9IR3Arc599s63K3Cy0GHg56MT0WD
iB2O31L6/RaTpuJS5IxAoCv5aUJ6fgJjBk3n9OIEEbeldYc+z1ISBGlaS9Q6
eR9Fcpzr7jXDzUo3gQycP4+9PFJrIfx/2QowpyhNk8GH1Ny1yCEXG1j0TTBd
x/LjcnDqLECXqbQcG+5O1Bw0ielqRsne+QZr5G/dsOxPDwZPTqOV71EhUGAb
JYgt+A5NiVJbU0A7af4F7M92IZUTAGUAc9N5vRX2s52rgcxIKmw42mRxXOMT
8bw0Cu8K1gYqdnfNaD+18W7iI16r2o12OfOrrRx79MFTT2HIcuG2BUTwd2RT
5wZdQGBCtta8LFGaDEEVE+UzSwTPkzpvIi6xNz/N123FTMmm4spG+foorQMo
1lfEJnXpKTig7P2nINRkn0ZIA6uwHG6aGOVRVBOuDFO1B65y45WGRC83Zf1m
6gtdhS74MCEuW/elHAUGrL8VLnMXkAJOocitK1iQphmyB9rZeaKV/9DgtNdB
2JKLa3U+pVbyvTEm9u3/xbfo9WAq+vdud02COL1QmNyqItL0zvm6DmFSIIKk
qJqLwiHw4AslGH1cOrpRrtgp+kPb+M4mTaqFQ5Q9p5MPSCPcP0zAgWkpkMUC
3DEMb2cyPQ3hGYYlgunQt1m5GE7WExq+OvkoyUf2JdHlWMDDEclwWokftffX
EofVkiBCaT8E13u54dYhP1xFzCeQgTkk84NPBGVLmSAlhk6AKXdqQSISssPC
9sJy0wP22iVJqPWloNwJOdWPuFaQlU9A+txYf47zx3kisAPeD103PT5Vs+yt
5QXI3Xbygl3WCov/CBSKiIbYY/0qToP0+Cctl4KG4ItHKTxZoxZhdo4wxpYH
uaGw4YB/dvxiudeKvV8C/Fj5R+01Fdgie3mYy7wu/X5N7uvDmi1C3cSg4UWI
nkIsLz6e+JAcbsWJOuKLW3levQgf5BKDPPTi+3OJUF53xLQDZ32h6kLCo32h
PzoHFQrrB3lp4PS+SF7DJV5FaKQoj86ViYBc27cWq1Hj8Z0WS8BkmBz5slam
PsZSjE4XXqnf+wHYDD+jnurH1Ndgxf7nBttwoWOkmteC4GT3qE+Msq1nbaf+
ueO9/T24oZlU6kFzv10PyVkALPdXpUIXM8056sNcOMOxRtsJYk77HS4rmVj9
+Hhsfr/Mnpj6Kv7ZMGB5IZlyoFIkd4dQp+cLG9eTayBwHUbjB2mwMIfIFHDD
+ZjOahM7TtvziWRBxF8jYrpcO909DUp6OaBGIH77s7iliVIRLsV/GegsoPC2
ItQMNBMVRw3AammB/eZamW74xnZT003Tvb7PoJgUNjoyUirvcKzEYYdMzyrO
rzvPzgraHH9KjzsZMrlpLiICDxchHgFf+/BA8MMYygc7YHMU3+FYSHMSObDP
EpskCLf0EJeh86g2YL38vsYHJrn6YPjOKb1byUeUOZ9Ex81BiHFoO1vFWmX6
MNaORIcuSz5LTnk7v4GRyB0qXw2U4o9vzhNTLEvQyttOcIKcP5MtEY0vK8Bi
zAjAVrlIYBcFkGL4TNdH9BczNoMf7XfAdfQAYYHbAIA3YKSi/i0s0ovv/gTe
WPx8yhFRZVYwyOXoN5ejsy1SPAerimJyb4CQQM5aeYO7X4trq7vAUZehKbcQ
T041ge64XZ19KCk9CBmcXVK/jFUv6ohYfs2Subvmyk/ub4BX0afhyF3FG2zZ
4wpl0rZZoJPb5is3U70i5Ox0L5vcxgtpiyNpvGA594zP8cbiOYFHEXWMgb9o
xCB9PjWuRcXLravuRHldZNZjdSJ4Cdz/BMMHga3LpZhEme7aU4bTa4ZLmcnu
PcWjrlyBwe4cftqHuZh7J7DbV+fAFYNf4rjRFdYgbJBiAorl0QNELdy6AJcd
uFI3qH0sgRsRq0m6ms5MC2l1SY/sJ8LadVmfx/dK3nxA6zE4tVPsHJa2V//P
40osey+Frqv/PSa6xIztihUjWsSDBC+VEv2stAOFP5mc5V8T7fJx2qLTb6IT
B5Je/KeKrrGqfUxrNH4McCdvJ6zUi21B9J+HfRiP5oOpkLLF1DdF3ve/ZlSX
KXxuxZx198B+G9zNcrp3g0+JOFJic/GHMBP81ynoMqwbcuZt1hbDVJrwSCDi
xmnYiMblmYmv3DtIVmPvQpQxw0Oz+qkJvTZtNfWllzlUXJH3UKylp1Xb/1qR
URpevGh+rJda88zmow/OeDoE/aSi+PDBKZAGtDei/re8R/2Yml4IvwCij1KE
2YB5hUemxStz949gcbsTr60PS++24yYqmuq4caFTeuhnHo2zCo8tEDuRgtwC
H6mjVbHQb6xXAGppDK2oXEY7UutZv801CevQ+CG6sd5CRMR5l7CXDV8HQ/Df
k8cJLK/3QvqHhpE5lt5/GZQ1G39nHtTodaRc3N04mMMD7srBjvlIiZdvwyl6
BmksecZbKRTjT9xihfa4KJrmKuC9kuwLrg8HWI9EP0URd3VnB3ngbjv0izoq
3se1173vbivxpxvY2nMX122caIcJZV10EWo+Ec+SambBRIVTOLjEeI9Bub0y
7rWaWiaNW0DN6VwrEG5eljmoaGyBavzK//FvcWgaDvcx+iJM47Pj0U4IRY96
YevBD9IYyWS/9JGlFhecuCBx5d8RY4LWb3+eWIBHm40rwnDKvaBanu9dKHNL
0ozj9WprVmNvMn+r0omZScuCSL7UjOzI+HsfyIAgqm6t64iH1quIVzRHDpRq
4RW2bl/MvHnMAv0qi/2KbFa8KoyjM2fPWHvxg6gl3IeE9whpeR+9d64Mkinh
Hrf+k2B4PAy11c0GsPb7bPWWCoZ9/F4suyrcqFdGKYbC3S94faodgrtdGi/d
POr0t7zzhpUc2SJw4jADZZ3N6cJoKOFEmFsnkOhTBZLVqH30Kfiq2PmmCJi0
oY7RO9s4HmbyHN++p2Tl3KhxLjSMHxQRcN0O/vRVzyioj3iMdkaiGfsElyyj
akE6sur9Xt+PP7x0EF2Zus2PqtIidXfFWHwgVl26e7dZCylOFh+qohoaiZ08
wcf9e6G94QGi0B82mHb9M8q1O8r/19CySBsOUN2FhjWQT+XB0ELKLI7u1leK
UELmFQ+lgax66dPH4h4wz6GsvZaI1jpW9+xyXLV/FintHB+NjK9L4yeb6/w8
Y/rGn1tppzxcsxp0Lh02ZeO2N2I2ftHbG4fnDlSy36hHY+c++ICN3WOK1KrH
3mK9szzUER/ZKFjlyZlsjtcbow8axpym0L+ZmQzlgauHObAOCfV/GEnXGGEA
cA8kMW4fCBt4b5DFSMDrhzTFZEUR05imKcEUA/zYvYNgD2O5ZzBqmNZFH+WD
3HOC3Fj5GQ80TmZjvc4dEI3xMM0mXBqi3by7+gIF/nQ0xj5h+sQDf7mVdBVn
6HzfE4Aucy3FRl8Cc8vI34TdTsyqvIQn5veIeQ5IdIudJDH4/ya0AZ+f2bw3
/Iz4e7VS6HQtoj9ruyPGzwLmk6nqY6qEsIYsLkhYukWt2vslF0WZvus91K9F
V/x1bwCto2iQo5/o5FiDsVFVEdc90RxX6wEEti/OL5cMxMIjcWrKG9O/6J4/
4KUqcRFuUt3WpWvv5QP9mLMvgRoBP7J0XsbxyypTfZnHuY5rCZx6mdDuPBRd
zWQhboyRtcrHqd8LgxVQVsSWrZ9MFEXeFgVVdVKTPhTu4cLc72N7uhyPijrr
0mpU92Ze1FnQ/aCCjDxsDcHpgk+q0kanscP5p9UPguQV8hI0S6QYuyHEFImm
rJxyPpUdWRk2Afdtlte5Y8oimszhdJaCHWsDdJZ4TNxlgidmE0HxwfevxCJM
yzaDlbo0nQMn1hyNnalja6TG1fdE67KAQFXtQxLyxkD+QR1T1wr5M1Ipa1sz
lm7bG6/ANtT3Ap8sBGq0tcasiU6nQbymvYY9RUXgBIouPi3oJeN4QY00+la9
SU28ostr6DYj6q41G/+7gy+vR7uU4rwfVtW9TU91rp0kub0qUfqrc7gVa6S+
tVE0SbdStGzKDUvhbgzbGmHfPTsBfN+xbp5XWLUsjqgfy0XR+6biiHI/AJVs
pkkyaOp20HWn1P3y7Rbxsr7rAEBHTfJG7WOVQx1Be2TbZWEkpsCmXq1Bt332
++zB0y4WIi04Lg6Zw0Dh/uywXA8+ftw2nBkvuh7qmjaVc07D9cEafFN54aet
TIOOndJDp/GXTanS3DPDJgD0VcdWxCgIWcoujOTg6ILNwynLC0FGaSBEarLL
R/cIjqTUm3oXbtLQwzqnLCih2jEDhlUFkgd5UL9mdoKHLz468YLgBQUE+zgv
XZOk+07IL1udhbOpEWO35LpY0mfa0t4UWIi/3Il25Z4wpvDLPzLmxj10sxb3
DWlb1/xj6q8+tTRz0+fjTGC5EcAXrzYXuhS0gaF9WT38txMcCJ8pxq6alPOE
vnvyru/zVnoKvIW2vYGDBYe94p7qE0xLb+FtnwQJcSscEcW6WyQfDTdE5Wig
mueQDKlzijnnqW94JUmB+aKgitXPnAQNE8znr4afLQ2UotkMP5g6rRQXnSY6
L+er86+bdmoHIaGbMO6ZfRfWZf4eZKjGBHeVVENUL7hKxcLA8NReyzb0hhEe
wTFGskbRh5H7Oq2sYDFumZ+KgtkQlQKv6Wb5ZxlRLHlwbwCxy71oG0DFxf2D
x8yAATxApKqWaMmA6NlqlRTo6XiBCOFlK1e7sLH3PWyd/yCxzuN2silVbrHC
j94LJUzvU8udgMld66fxcBdkFpXaFxHTe5eSQSyaIMqud61qHVT0f2K2VnOx
eK6DH87ufhla8jogVERKMM2MBTkfL392ouIqCiF6ofSo6ybraM09aFx3uxqA
swUwSp/uGpHE+/FIqzPdWN8pGzc1Ad+leF8jcc5kXaqrTztJ1plMkHHaBYNu
Meja1JfDuA/WbRRtXRCs/egKk9QbBOiLPbHsQJwKH7we3iZpbduTa8xSEGRv
6Any7hWuoCcTpg4QJd6E8Uyq5eFEfIDZ+ZWrPwBy0LhqnM7K3EeavnnaEfxP
B9zGFo6a4g5My/Ky1ECHrCAjnsBBMayQWSwFzWdujsFqPjBNZhCkDeRndbfh
ZGYXt+5BV8Ij4ZBcvwragc/yedB+tCU057QDZrOfpCig2wXkTdfvHc3mcMyY
XWwyO/FPY/qHwDZzSbhhC7xVKe6Z95sOFQ10W7JrWuGe1wiNAJdSpTO8i6tx
qGqjn+pidD5xI4RR5n5SEOxmuXcEnjudp+Xk+UrCmW2ZWRnJNtGUBUWayuBK
5/F1cz5btw9eNvNcQ4lA2cHNEGLa5wikcKSOQZMgx0bfO4pkAj7EEKAObyED
97Bifo1KAx6yEcJag0tMjkMQQ4LasBd7F2b3hNKCO+K1pKjCA8nxYvHLACEY
lummg0SkM+fLpwfLOizIw18aAYSIjZ98ZuldO/CvhEq5rEio+wUFjzZf9b6E
Fc1ZIis25px/XHOMEg+5yaDwPQWUh8+U9eaPKaoOw4Ob5aZ53i5/tGFwbKO/
FKp4G98QvZwsv6FpR+8By/ypKsSPsoz80UfZP/ns2MY9JuaHxB8/AnGsSDHq
4i/RUlXKJP5H5u1xKVHsbJ78FHmSIs2EpG0hkGRvsifeC3os1L/1viq9Xoo/
FzjMQBYtvjDgMMhjUG+u6Qi1sVWRRWYNQPpXsuRkZYuF+jawrnXCavdqDk1a
Ggm2lo75cn1EaJ5hx681PdRbHut7ikfbP19OnNcIKpMUb7RDYw8xITMGRE/T
HfaznJpDGuCcjygJb2EMaf0xjVvmNNGFF3gaywEgEZ85LydBUivOYvZVAFbV
wWufPTix/4ppKFOgySHD1RlVRh4Izd+mG9//UxQBsuAy93GgdXeg04z1Zlur
GC4WpN7cXgsOnMZ4y0kAArn4WmUmjxf7YT6u3ARBLBrkLd/bKStO7OQYK3PW
XBIDh6ATaxWQUjMxWepChz666D/rFpUWXMiD8EmmM5l8GHtsQM17zyxkkNrB
bjOrnuwObryqij1RmtQ8zFrDn9T7jy25sTeCzN8JFYwX0E50RYD2kJZmxr9B
+WlqufQR+V9QShjKKbvByx8U4i5Cr7EoTZNeGCQsbcVdAYTXLxjOMAfgnI+C
qgy1F8ZxfDNqnNZkw9VMWbZYwaO8Od1C7ZqL7g/ZYAo9y4MgRmywHeV+apmb
Z1Vv8cH0qL0U71z4pRIebJdCbQkT2nRfztUaVURCiIPKvs6dVbiT3BT6KAI5
QByczFhlJoVDAEnR1K4LjVqsvrdNznmgZOPrsa0D+K427u0RFNOb8yrz70J4
2sxk3XHoL5ZHnSgZUPzPQ83Rt/F9JieYNMCgP5xMXLkg6jG3T0A7VvJ3jI3v
x6J7+L8DYtfnd7QE/TEqIgJ7G9OTO11swr5vX8b5G+bXgW1C3gQuyng1h/K5
TGRdzFp4dsdmRsZJoDdrOLOCKcu6Xswmd3tCpKgnMQWAqqGDkRNOP4B1MaBJ
BvSPmRBnwsnSd6H/cPKTmx0fT9NIuazaz410iN2dmp3xBV+5fZ8mLzCbHmac
4TMcbJictXs16626YgcbQOdLYfStcnZvczcX51sBxg7N3l/JzyS/ObwprA3C
ei1340vJjjoqMjaXqdNIVBZUcRLrX88XyoxUmRNY4aJZYVrox/WlPOWqc97i
px21soCH4JT50qpUkQtNuPbHcjuecfNM4PCXou2wddv+vgFTaL9/Qd+FL+IG
DZi+yn7fyErz2s67MwGY3ryNF1SB26e3a5RoQyIZXvkmJqyly2xpzDrlGh1T
fPgHkJeyKPsxU8YQZD1UiHyapC10i3n2tKvJUoR3yIOYMTh9uSZmkubaXz+g
12/W2BDfXw9KQTRnjsWhN4VL4KzeCbNkkiIcfh9ooObDj8RWkmJz6CwNxsLJ
eerwWVDx8SBh6VcnmKI3IDkVIvJBU0l/BrnDJizlh8hGd7cUL1o8b8lQlIn3
WLiAF8vv9/uqXNx+SJ+cgUxktCzwOItPwcrj5Srx50NZGq9+BkUG05sNwfUO
DmvPzVcKFDMXLetkPIsWVsMg7cC3gxHUvTydC7nXHtbtW6E6l1yhGPhzePpw
tOPUtUp7+SBwp24qUua/5ebFZR38DzAJSLzb+C6aPdYTC8jrO7Rg1peSfTDj
TMzLwguTu8ATPP07Mvd6r/hrRDDFc0ZrO0wP3Te1ThWOlxQMedxqkBPXDc7o
ZX7YaozijHKS0v/PSpewnnpwUr4z08QQYPv6sWdhWA/pS/x+Xem+Q4f5ktXx
I3h74hw2QAspCsZdEjd51fJpWAeHkpOHpXqvLqq2+jNFtJiM6x/4dfdRv5n5
Mj5VVhnplCtDyzM3MvTfeKsFSSDdKHjc0hHCmw/JfLLy/S/gNUQxQfoGTTru
G02L6/OJJYFXBKbBKqmGz2IL9rj1Oktqasr3DUeOh0U8FZ2OO4Ybfx768Ck2
4Eh/4b3sH63mNVsGxtfG5DcZxi798uD3Nno43z8uJmbQec20mWpgWy43AkZz
NBD/QsosjC0fgViwSTFMvN3YqXKYmBqWXXFvxGBBCoDKazB3FERvQQwaNW79
SoVAmRt9Rler8avMEMPBrT3eGWbd1JsXsQfhCtwY77HK7IXjYgO3P/UvMU/d
B0IV52nqd3hB7BYtTAwGUbuEd4T9DbTooRsq8ILUCnS+suM8qQXUoKeJe+Si
fea5GmVMoog8X5F7TyBrFft8Mj+3BBjb6hxxIK2ZEN+d9sx87vX9iQo15uXC
pwu1sNX2Ik4svtM2T5pJVyAJGIzJeNsjZIvRQqTqpX272uOZpmJf+kzEnkIR
7ndNS3HxmtTPmM/ULP+UuOqQASJ9WcJbs1gqLcx84tqwmDxWXI8M960bl4hC
blBcNWGvSduIMbic7OPQesODciUB0JjWNrC1DQrqWXWUaEaVgyGHfOccxMuN
1pqijWvl7QfiqmTQacf42rjSXXzQIPeWMM/wkjonjNYNsts0cw1X2ZDWvinQ
AFGdcl4S0meyE445TloIwub2+pazEVpqHyA+Vvtt5NtcKJYqrI0r/4q+zcCA
gRVfIfVJj+qUoJSq2ey9UkzCPv5xYshHJPDr/P8Emcdj6ynwbQ2TdARVvF9n
Q+JmPz+foCll9k420I8IaSiii6WMM9rZ1EqyMIaUppOOHtm+KQ9TCWLW9ZG4
DXRCEfTZhyFZDnjTpyu9OLxoZWrFhBrvs6jWkVfICAtVf9ilBkJQ7t7zJOmq
NRWnf2enpLfUTpdjRbP04Ig7DpLy++zNl745G8hw/CQAJ1iWCzKcrpAhrDG8
pFf6DxxrUrrApGTGncSucfOZpVfb9vGOw7cKpvL1ZFcCWl8sk1ItCIzY0Nb0
lR0oHtldNTLgowtEUdD2O41BzAsoCfuqqd9XQGqu+xOknqvEU+7ZyF1gDgZL
FIv5RYgv2bMzk3Cj8dQqHL+qKMMGLMzQiiuWp8YY3nJc40XepsVTsAgBM7vH
HU1IilPABhIm4MtwhXK6fZ+l3BO6IE24UxaSyKwkq4tB8r7i431o4FEGVsEe
H4t6DOP0brssP+wWkDQ6Ean8hGcR3eHweI1jsWsNYqHStIjJSHjq34akrc9k
uiqycoAHQ/hndyEPM33NgD6esoQZ4jXPM7N+66uiXdcYQkLrERhaQNrf0I2D
3F/RpQ/1zGc1lgaaPDROtbT1a+FMCEb6uNnni5y1OJCOYqUwVMsZayYDL/hC
pZFsj5YlG2G5/BhjZWe1AMfsdcocRd1RVBxv1OcUkC0MVHNapI5t4ZWgFCSk
lEt8c1M5gOHLZCafMbknZs1IDTDEafKNmspsy9RSPl6q5I83uLuBdmOI3vL5
GXPDKrn+2JEqCmyf/UpT51DVoFFsjEGeA8zGtGOMwZlTfLGzAhcO9G4eSa4S
Gx64UvHs16arYypyubxmK7W7Ig03o/gTFAf7mERkcHTnv8xCnlb94p6byzu6
K3CqDB0bysXe8H5JYD46DWrSKBvr+zWLNG/B+m3WXaD76CtuPv/kOElTw2v7
W4XN+UW05kzn24KfQI1UTg3BECW5cHKu3tuLjgnEZp8wJRwqRaGTKR6jde7g
KZqBo/4xlK1jSnPpF8XjOAHeS4OZWllZS5+rY58bDL1mAEOvVuYcrRbNqV9/
ESfk5M0ZURzDxEmErsrxtW4SMaCvawIKh3+G8VexLozK8fJzohvY8Fv20dgW
72oFGD9JsO9Xrxocuc5F1XLknTGAg/Tm5jZ+nI5c1E0wXTvvgJ6B0Co9sTZ1
eH+XCl6d4xCOqYwXW+zwkJbOOSQTd79ouZwGTOF01bBbEIs1ZX3rJVR6kKzf
gmPxkAhHJ2a3+rkdGOkfBfvFjV66iqJaYIk58aQokNRu1tFXtGne2qXdGbgc
6iRp24AT6puf6S6eFfjGj3Pes6lojAvacJjjBtO83+QCHG311ZAPGur0SNij
FQhdwmsln9yuwlPza7ZDHwQWTe+/K7L47ZaWkyJ2hQBbW/HLPVImAVCbG/Ud
mcbGb7/lNxHxlovOIudaU/oTUA3FCcHMF/vrQaR+yYA+MGLkHll3oMJVSkFR
bZUWgMA8NetPGPGHKeNzpSXsna3WcdV6FnuKZfj43DD/De5/jim1aLimy+Y2
v+wn3Nyvo6xLbEMOf7p6k5qs0jPYfw+XexkI0a26IPph6Avi1KVYVe1w7K/G
vqlxNLSG9neVbLUdw3K6Twpe7hU0Ug+wPL+5g7IRIuiyx5W7zl+Sm/58Aj/Z
5gMCZqq0AfBAzbOBckBIaw8pCfwYIZYcRbnHEo8CMCQbkdSwz32IjlsxD5X6
O7BgMBspGomoE1tQhDQiW2jMeyGkZQipv8iAXQv5a4OkLCjN0Te4E5jLiST9
nmy49ZQ9wPIcLkPRcK5YJharN7UYwCGRtTziGb7+cpOTD8EtH/ZQMYTnvKWb
G3AoGiNG6Zr0eWxcy98IiaNHhkaGkL9vb1jx3HUyozUsXLuu4UdhyVYth9lX
XKgYKJDRcqAzbsZ6nQkWtpHT1QPhWSPKfeHUHESgWXcF+XjhCzipEcgqgoae
RtAsUPn/0cZFxbRXoM/Per/U9w6Gty4+DbjaCAV4699QEOO8iVZrL5R9MIYb
9zy0kuFy6k1LHh7QY7TuEoVFDQfUTg8M39NWXoSb/nn12UjGzB0USlpJO+hM
ap7GX0BliM1kq2HEPL/dnECnmSwrQfswlYjpzBq34gHTe9Ubp0rhVO9E8f1u
CnFrgfVxYAPmeMXXJM0iJbVKM0d+cyQ7ubFJgUZ0uO25wP9XeLHY6u+slxN/
DSDAvrotJcsp9IRHdPSmSlDUPhwVJl9jIe2lYag0kvQYWB6ZHj5tzfdmGJxh
ZFPyl0I2zEnqoNbut5fBX/Cx+EzUOWRm8/opA1ApDiMnQ0vKKzc7S+1sCXWd
6ZHjLBJhjJn0OLhDW3OG6CrDBlHGx0w/HICs8dlcXRA/niHC/8Jakzi1f1SL
KFna/kfdanwCBUvx1VjFsQkRJt3P/lrqol7hmADCLBA54W3vzvxdv4mrLxwX
TYfEIZMpdcw0sqOlczZ8uhxac/+4XHbmYr4WAS6WLTUqSL0tsSqfVOFnFLdq
mOzQsXLzg2lMmiWzy2Ai+rcgT/ag4jd8M5lzRX9/rBeVkBqjEPuMRIzqBEuP
nSPRUA7xH5ABqn/8d7nPmoeEsV0W/gzVP9ZDZTtIL+xwi95BmrA84ynCo2hz
2LOfZP5QHdwvFdkLwNbWMgAViKB17ApcybyY2X17OKeRDDcLud3QE/nxJdWa
mOY472FgE4wdyPPxV1k+BqUKkv3f2YHBJyzm3NDY6DvwHpjXBM529AFlzKx0
qgpEuLqU3wSuZGjct5V5zFADEIGX90t/AB2RqbLvFRB6+vcXl29icw0Xvme1
gfbW5TtziGUR1cjKrF/i+FcFFHS7b38tcTe8a/driYh+/B5463IDXozXPjS9
nu0ljUm9OSH+eBNLG6YDoP2fNud+rSf7OPHt6uxop9lFJXC77PaRUkVc0W/0
36BTxUSJaDajUnc9FEVtMpybK8bYJaVblKZmEuv+JeDj3+Ws07eW4DB+tQnv
eeRV9RGw0HyeJqSgHmqjX53Ki61AxJe9CE/mI2VNgeD5JRYRz0H7FOmmYz8u
+J0GiJMeNFcnwSfKBFZJi1BsBxBf3yY5DkV0KrV810gLcz0kCBLttr8yTAdx
tR5dg23dFy7Xe7MKXw9i4uOT8hP4YFrqsnr/QHEpl3bAU7xbGDDPp30HvIpa
NSkHZm5dB7PmzSXomDTPnU9MNMmmI+q18YDLZ7m3nTm9PvsR96IQ/i404P7P
Yhy3EuE1b6mrRwfJrnrW8uGY3S16vmvgUBIZRbef8Mt6Tp+GLjTd9y5WiS7g
K/akPVG3JdTfYgyigJHsmsLQO0OJjL9r/l5fR9e7O0YnRDIDSxLMbkA3bYVU
/jJWTHjrlrPnoHKqeWru1wzhYHFz0ennEJfG2XK1spsOmJ/iGPyCSu62ps4U
60lAB4z5XcRUtUprilLK3sk21WFBMXTEHALI4hEXK0q+YfLQyp8ntmpOOSj5
B/DiTN/+bwWSRmJ/NJQIZ56B4gvYnEEkQwIeBuhOIV5EWrDylGrVuqAkAkA1
h2mKocaQ2oW+Z4QFZAjc2m35rbev8TTRYuKAgtNq13R2Hi3pSSDRh1fxD0VP
guHL8KHj82RBFPaTUER+17T6DfQ78n15IoErogA0qRfxduzxNPKp2WpFTOZ4
4C5HzjBiJ7BIhxRS9IduTaQbFKqt9VIKvmOOXO+hnp/FEi5lgWhiWp7Gg6Le
ux+m8B7nZkpkNzesxOeMm9DiJBQ6j4Nr/H2zdjc/xxW7CQjxK5rdCy5i/HJv
YKJrguH4dKUNhc8TDhhz+I4Wxdl3kwdsDUUoGc22CxMjzdcly4wgvBkCFPCV
2f9+Jbq9UnRQGU4y1tf7+K5deF4DavmFyLVTcD48dVVWmY9SVbnAvvLz86jY
+Jh7BlASqO1U1RTI3Cb8EUPJKdcbFmDG+ttIptNWQDHt+BYEwSg+iWyUd2mq
QS4pR6utOXX/DPcMUDOMCgilLaVzFZCyjZSarGMdpcS3A9GP5MyeM53/YQ5K
1GuCbGwLpLUKKHNRwji/hMR5qPNKXEFdLmG6pKE9TB1xvrDeZz87oGBnHGyG
nEfRvFu9toXCDMlxR2NmWGiRpnHodyaeboxM3C2o2pv/ez1D0Lblpo42qna2
BVWl/pGytZdBGJlV4Vdh8E0fYF/KTyorxX9JkbbY+mCrM5FpX9qptxwNXU+H
NoIC6i8LvcxE+TyRWx9jEdpRJ/jdWA8X/bgR4ZOhYVwElRwMjZb7BOOugCK9
HVkgURoXLnDCWd4MUQYWdbR94ldR64hVItyRwjtwiTUWFSgNkh1HnGf8BKjU
7SolgS0eZFOmoVPIZtFnaKd8tk+NiArCtb2N/sR77w+NpKp9Fbddi51V6grF
0Yhhg8D0FBP6WtWmOnGTJTJ2yU6k2c02RIx9ECJkh57cnlng918Go9bChSWl
10atcaaGugdWOKFjmkOU4j81kCWl+ew5cYH+ALpqyPkJQAZgFVBHKTpJTkHP
DcCXPdHmu1ZWNhNvdesRHcOTyJ7lv46Zr7jVnyGPkfqyxHniAlr1aMGAqf1y
OipKewW7NQXCO5cA0O9rFASkcpFoC0pKBNgZeiD/TPyHTFTSpDc1DHMY+c1L
NiHWbUFw3S6gjVV0znquwKLEcUT0gFvv+EdoKm3pAPxF15LcqRYoVGjk2amM
wAc+I0l01hUw+ifdch8WsHEmTt5cGZ3gCnGd/9uK6pkVfwDHTbbVRQQJk1KR
KvxeC7+1u+86qI1TUYKoPBMaZjRwDC1bmRoeTEWSl8BosTIGalI57eoLoJ4O
yUx2EaDd3GfjDlvGs3NR19qvo6HiScAS91IUTu9YQwr9uxv6qjZkidmK4Jgh
uDXE7fLyUCk4EtPsgDD0H4/9wumMZmo22ZM9elgR+j3JUiyr1CVTSIZ3fWlq
r1NPuUirwviR4cRr5H40TtpIu+wnAxWFoxhWbT9zVdlNic+/oi4MJPk66mFv
VKQW45/up0BOTm4RR1ngc8dNQdD+wNr5lWgp4lmikb2dOKr/SyPH+rOO+aZG
qtyBVUi+evwhV4cU+Li+WwUKCiF3+0mCJzqoqndWiP4kB5Kk/gAsAeZMyw/s
P2+uLadUi7OGlw+5xq2QfLKwsfhUBKuYRd+cSN6kHGHk4CAcKWDRCrvj0Xss
tMnlNgvwyMVHiOFOGYjIH3DWhZEjCfvFRmGuKD5LT4k0OlK9K66Caql9EFMd
o3P1HNiB9qy2Jx1rwUB70KgmhVlvSqxRjRncVRNSbpivyKxhlk3tCkpGdFMS
hrHKrBja829qWU1Of84GzP+7fd7UDw7arKA3rLMX9rNbKlpA0AokTzGWRouh
ejGlex/R9VEMl24UXFxbhJbNigQBYABVfpnUSucTzPFLjMfptnRW/9PYopUQ
ImO71GolgcbX6lxK4lQ3jTIitErr1rQNLmN6VOsRB/MIGSmRMKk7U2rCk/vN
kJTDEuVAbR32opW9dDQ+nAgvRO8kfmfdyPOMQ8BbheqLyprfPMNtVM8uT4U+
o7bBYOSpdXVayOAnnvqfaO4qcVumoQPrI4fhAfoPePFlmeWoZYr/0PloRvW0
d1XUgSqHw3KviLnStacvUHrFNrdbvarBdJk5zGNSwMfxcHcuC0PdKnX+I2QS
vmOKZch4r4Np/7nYr7m99FjLDMaGRS9bFowScRDZdqnz7u7OuMSTAgGsouTN
Q9jkFPx4fzKS4Jut9jIytyYdbil9M2g5S5BlMTouUdlDizDcDcuSDCiS3aIq
u4SmDc2J2G9PVG6FrU1LxaDCv9pnK2Z1VMMPbXbM7QORFuKAHqnOWadpL3Sf
OztD6BI3lf7IeUxI/W2Ik6euTnKwtX6ndIfBENyLR3yFRn8iauHjz0LRp5mq
rpf4yezDVOBBL8dVPFUWJnILoEUvzoQTm/S015sQTq123rQ+1KXk56s0tg8H
TDFNpBy47yM/UWTvsikxQrNhEG+PT+S0nvkJGEPqX6Ns+LkUVEgJPiPqLgzq
Hfa7dQMGd2fNS4mAEYbnG07isuu00SplBkzzYDzt/CwYi/bI0o+k3IpRjrs/
ZzHuh7A9BGsMu1ia2OfFbUjY8zOxNvRvAefvD3kTXxYap631dTQnUMvyNrJ5
xJ2vCkK5EtJU/h4bFy2AWCjX13w5/QsosRaBACyS+VHNW4NB4s0ZRNHtjKvu
w2/bC9FYCziDCeMuRCIcQ5yYplSL57JhPVleomx+W/QSCrKVD/fCVxAjzHLC
HvJOvrXDPRIqeVEYc7vXtaOeDxXjR616x8/Q0DYpR6GVtZV7TVHeEZY3CiCI
aA6tKse3t6KqmnLDyAd205pA7b/gPlNWS4N3QizAx53ujqRAUDMOpwa0B4zj
RHeEBodGR+kXQu+jyZKEepzuFieSjzedQyWeAjT/2mpeGsGaMsPNnWvy0Urj
2OKyAv6sKrIbAEc/UfrVZkMtakc/XX/Jx4KsM/N8xwiUb8ipybcNjAopjWPx
YDulw6k0kSF3yzNzsa/P4tzCS971Sx0fVkmF6HkA9iBK7wpLtNNfbQR72OTu
mgDDQvbhl22VAhozCcYuPQkiJzfd0FIsmyOWOI5XjH1PSsc6w5VABhuiy1DP
iSUNCZy+fJwCqIo9Uq1G71x0NbJULKK9qCROtcFL01r75RlrIplWMrHQSRNe
lSKZ7O7IrQVQkQc5slCsWpstFMRmbFuWuz5fRifdu8jY2aZM8gDcSTpynoDJ
uRKsUiVzq3OZqpUTtK6IoTyYtQixl4/X4SERMZ6CjHdBjGD7xEpSQ0kNFTRz
jOs7XwaLmD6dBfjYy7xbsGAmq2S+DVYdbJMrJNk00Y69BM/85uCnjlo5HrVB
pn2j7ywvqJUYlXnuVVkVUxaljreYjAi1U1GZwBx686LKCW/rRNCS525ysUnY
TFSPd4klLRXpMBJ9h/6L83cGDXVaJlclfJfFuphiRqoOyZxZ/WN4+yqhSPo1
q3XQhCvUlJaPu09jhbD/RTBJan3GnBg/s1kw1xpdMYLgViOGg0fTpB/4X9XR
SWRaiB2hHgM8/es0ycDZl5agKE5D/xGuHzbMahNv14nYOOhIpks2i1tU7Rvp
TNpuq1+HXtQY2MFjPcoSfq91+gpnZzCTOR0koZm5EKqcNHJzfYqT3o+BMZ1S
tblUXFdv/HtjH8aNiatgDbjTYqKxKtVw2OAaskqW/tEYdgaIhQdVAHCl/E03
Qn6kk370+E5LdAK4H/gsY/BOaaW6dgLvHzugJMUgECbTIVIynw1EBYJcZZRW
Y2bC8rLD77Ee9+rRWyfHOIwHRafgTlDTh0TVCz6f4BT3Po7yQ+Lz4fsgUceo
9SE9uR3zWd090Da7j0l0NprGgBGmUcPHLpwGDRKrUr7sWBTg80btvWZNp/0D
2BcWc6v6VUtJSXjOs9OAbbjxtj9yYqQVJ+HWWaSIEB90Xat20xCE5LWcMJO5
o2O9c/phxTy4yfD7Ld/Wp3jID3yJIOQjUSRZRyKCqQh7sqQCpX5d9sSnLrax
eOKxgoajnPbCJ9n8ss+/aoBLpA609UqBF9RP+oQFedEFoOi5/SbpyuYgW6RA
LlXfEb8cFcdsMT5Z8Bn6IAOFCM9PWW3tLvKlYTg8cf9IHKNJ7Am/WnslBJAS
pjGwnjvffbKL46rgJQ2l1WeaqwHSQJ0fCo8BhqGQCXT08LRVcurcCcarRtrD
7UXl8TiCAkXtPyS5oz8XOIM9Ts2qkFJEe59VaLxcxc8cMQS+kYG0Db10yOU/
4pdGmcGGpOPi2ZDg81vEiPGUcMgopcvKZ0gTV0bKsuMcsJwRNxg7+WfdjuXz
RRsF/u9+PqSNDqO46FH7SkMK8O/QazIbGaL+jKtzQA+p01HukRYdXBX8Zi76
5/CnRKSxykkLYycMuz65lHQWsfygmdM60SOmssM400YFAsHJySYLghwhVgMB
JHpY6QiIr+ZWndjSMx3p0Y6PDpnDilMpb7T8SphAJx43CRoAdVKht9rBy2rt
JjviQrbCKI7Z0Yx2GWWTvjuE6sEFRjhUl3+SSd68tPV4LsvfYs0fdsdCC+u4
NgnNAS98qJSLidCdnoKKm/JUTBb/OQKW6AOzAnoGqMAtwj2W2yZbRFaoUTMt
8zRSgPM7PNAsm4W8yVaz8Uc99CZfNE63uQUx9fxmpZxj5k+FIuGDsRwWaUhE
AgjDCwlGwDe40sGl+xu6rvpumstYVWF5k4V6jAg43wAIcFxzSmeHUUcZ16jb
/6RO3PNNLsqUZsMV+/olJeBc8PtrCY+pLErlYXvKzRWf98kqHrYHB26hOjkj
Hhxm6O38xmSpiD03QLbi0ruL25d5DngrQKFbuFpEncetZIfA6/7QRfGxXFsV
H6xAJecLviIVlV7NC6Qk7ikL4RcsslfDAa11oEC+7MFWnxff4XqrgtZTabxT
XLBwbJYxn7qAcL/zYV8tUGIQWTU48JOJCcDsLePUEjPVpO9NWjtGTFuzeYaQ
QYS7zgqVd68U8ZTxdwybSweCY2hN+ArMZ3PLitY0JVLnp+XXBYNpBJDI5MTy
7v7FG99Cuv4GPPRZveJudNylOm4plez/jTugISVeyRXfjAgZDt0YVMABdaeH
SkZSeleLLAXTnJlN+zejlkIuEsBNdZhrZbZa72QSbGFjK7RkreXUui88IsTk
L7bpXhiTuQVu8JwEZAYswxoPmsT3tXcaTXWQELJwMPjb2H4FSueVVuLcej82
m5ESMlYlyYNW28Y8oL68fDFlMUAYF6rrPcEI9fhLMDKEFH+ON0x3WbWshdC+
b/EKeej8U4GPquW0eMfRuwOdtA9bf61x8ejznVOJWlpR5IltlWnDmTrluT5Y
W9jna9u0QPLoPiMcTTT18Q/VP7R4OD+x2zjPeisCi4t9GblPzxbxJllQEJbm
BnYElvsfF7QVLbc2kVB8DLh9WZzsNIOd7daWXxwP2RRxsHNEuD9p1urhRWph
TxOt1slu5FUIwlsbdjvCuY3mvOdGnwoORxT96paBO6TmhG8PCftCsq8qE9MA
px6WFHuUf444TZFzMv7YA6hrMdu/Q92FRIdNfbtk+9q24FaPFnpasKUNLaOo
fnKOlGEQMyyTL2lruqTeE/ZFkKzWvTTkYYLMnQGwCAUceY6CgH4GRILvL36+
8lmUiy3l/WEBg3rIIlLVRo7B+JRDPXu/JuWTZpIp3QWlpjFVaK476xT3oORR
HWlAG6+68uRHsB8qsq+J/rT3m4U2a0sZIB/xYHus3oxSeepA6aaw/KyiFr0d
f4TTfqWA1ytbIoVpMC7tMgwUzzIN5KTj0U0Ym08/iOXZFVDi70z3pmLMAsJK
FQk0pidTR18pXI0SF83ZhmOT2NGfne/ChRs1oV1MwvfhhQ5+Av7hdlXYKZvn
C+5xWCSnAZKJ40ExKgEgE+oq2a58Ir6t//hO7gHnVBnR9CclPt+wC5bDLjrD
WL1mWbVt4HTq8nYrIpc6NilG+Pxgr3BKHf+1JP/WCFtFG7vmHk5z/Vq4L5yw
Sh35SiI42MOqZViDVHPOgW0P+ZmLGD/hM2HN0kFVDipYlOzlQod38ClYrjJV
mXQQs6/5g7kxfw80BaGksxZjXloS65gZBxrgS+iHR41Ky16E0NZtfSx6cI/d
Sv+MIVmeWGSJUWbDxbENYLYylZ9GArZ7GI6f3VcJw5lKEc/bLkIsiLDfrbX4
AyVRjwEiiprRb9wCgGtXB89dINepbbLB6qLj+ZHs0KnxrJzljKcBEHBBzXHi
w9zUX5ht+fiq39VY6ngdwgeNJ0HOm/ddt2eaRiQQlkbfwLivL3UVQXL2mJLD
aIVEAbjwQ+qGo7yOMTD56vBtuzLqdnPKpbG9sbcaZ73Y6g512IgxUrQxDPNX
5VIjYHe44A07dZ4q3x3GNffyGhTet4YrsHsX9CS94m9VwfkvRsCU5eipn0EV
Z8lfvdXhQSQQtsxTrpRAOmIiPBQUL87+1DPD49dFu2+XToO7Ovdyn3v7h3mQ
6wYg+X7NEux7yrD9WfdxpJ4LUxtVLL4Fgt91mQyLCHglZy8/RzC4WedADV1/
M/JUS/iINhwsu23nZhJn6NgoLjgKN8eDkbZJeM6TkjzZUJNlwzovf0W01M8T
qCMYJk0PgTCChXe4yzw91MzI8YEvWAFw4coGdDZT+1QpA2iiXlyJFNbXds48
f3oInIuj1V5WK23QTP7Ua1QZ4i5UnTRUHGPrDXH9UJ3HuomKFLYSlJ/rkQze
sj8x4ULcF10bH8RoOo5imP6b1YJoI1rBiXkz+HIuzeifXYR4QiRxhuZgKQc4
VvbNbEZ/02vKnDe8DsBThKECTa0WT+Qdii4Okp+Kqot8XANwM1BQzRZnyXq+
cryJ9yPJy6Z/ZE8/UmfB4hTXg9VOXaDvOQ3Mx6plEInrAIyztVFt/JDcY4xa
WRhF5LLDvt/FRZdVRZ9hiPgUqIf3Y9t0SiN5C1dBJiYc6iWi+/KoOrT/SOpV
Wyn7OI7+DSdVqeOooLItB2+7JOvNxr+rX11NS/o91QOrAv38jUbDmWAOXn/R
iBgm+s5I/ivDf8iPRbvBJe0VMl1GkhUrPDPsIQUmU3HybKbocEs0ze0Jm2t8
VCrHLU2Nmy3jeACdW8s2ehjHY1oxf0xKPnOY8BUD3rvC3Hetgy0BQtRgbE9h
gEa1CDN09L1OR3Ni1ecDZZcgNi4cw5lfmTfvRwKB/SuLEV2UGcmSk20s6d3d
W5BsUfiQC0Ju3JDyGMj5mzj5bRoQWlDgYle/KrmJ1cZehzZ9JZCK5ouni0uN
BSymWayUfEnJV3nkjwD6BoWZCDWYI3cGSzRbLrzNkIo8By7DCZSrga3RLSXJ
rvt41q8r5CRwa0ksWzOb2U3kbFclZgkAJ6SJlzjxlveTZ+XozjxIVp/PKceq
HcpG2plGYnTV4kARqbQZsXC7V4Xq7YA5/VsUYuZrbaIOCkwbUPWFLBgyH0hG
6AJrRSOv4NKquuLhNQzhWsDDwInRQ9exQM5DTgD12ejeWDuwakKECcM+agwx
MEwG/uF65iI1yDChINv4dxDUEHu+as3jFLhQRnZjtHqVOfrGAAF6hTIjNakN
8W0q70z5wKEWipA/7Edgwc+ISu7kxh/cSfCGHuTByhS0etqXOSZM4e/Y9G1Z
X57DFWYvpdx72jv54oJxo6mmzZgVaZ/ondTiVYRe2DfIGgSfWzvlYXWQRmUO
+qctIMnIFruFBnZEGWZVtlchE0C1PLaxZT1vHYWxxY1a0G5o252+Xoz9BMWw
L+12Mt1BdgnOj4t9iUOKGTEc2dZ2nN8bjj6Ky1LD/NUJvpAN1hYWDhKMGp2Z
2avNhnllDanGt/h4gviIVgkKn55G/XhL/I5WxS/ByOROemvEz874Ly9OEuLe
R7aCuzDUdV7jVwQpYE4S1ESSJkUIwYXZkpuf3i9xFackF2Ijhp5h0NeZAU+5
pdfnE6oUSThOt6XQZD3DNSm411SCNGvLiAwsM8wWDs8UtQ33BcAUi9fLxdQH
QUl93OuC0yNak3qUSpABJkf8muE/NJPl5rr5UivnBuO78hZ3oQ785A/+evZz
uNpPulwP6SNFe4HCrPHmYTyHlyBBR1sw6Zl3FCm9Qv74xNseF1Rfz9O13nEz
865A6Jv4jwVliVqU8zXgAqWgr2N2ujxjzkXX5YhxJ/eTti60nunbr72fNEzq
rgLo5/fiirDuFZOydgNE0RjUNi8XtL8sEdngKGvm66WBQVusQPPaj5W1kq95
VhkQNfsWGuZvxVYl08UDbzbCZ2ZHb/PmZoEhkPYFOiLiiBaLCjQAPvRuPwLS
FJCnmtHhvSllqp5nguUlF7KP77B3YarJE1F5saX5QUSkeQriLYKJWNaW1S02
iylfqJ1wdhW1EZz3feSr0id9y7g7aMcwH3zMoS3GZN25tT7LwKeucSuL8snV
LDMDAN5fkUFQthf615yPg1Hlk1YNFlo7b45nhGSHV6oAFvTnCFjLAhBvjh4A
TDSb3XiJFoCK3xMfSWAf8OXLi9Cjba2EHEwYYUpe9EGBev1NJ9VcU+5LRnoi
wn/VnYVLotIBfbnl6u1W6pWuVBxOz4ZMCgQzoOVg7kKLWltHAk8LnvjeuePl
fD9DBxdienFIAe325qy7QkiC82163WWKa2e68nNoiGJwjznRZAmS/zaWzbjE
iEwd93SBkafQSpur5v8W/f4X2wQhynfICeh2m/4FfoQ3H1fC0us/3rjWazOY
9j9iMO7fSRBuc3Oe2HG8Hq/rgsX2QmO9f//xhAlf8ZpMz4FPMxMSPAM4s7aw
maS1me/ey7WWDGO4whP6Jv6q25f3zupXM1JtgRXJ6CHpRXSd2LPk9W1hwJOa
CMxbGZiTLYFYwFRgi//sEQa6Iw2uAj6PFV5VwcglrMGWm9smMrZoJvDv4XDS
URpD7bgNeM+uQKM6DIDfhDTOC1ztMVcxvS4OEv1KlGZRLl6ZNIUKg7IyIaBU
kJhA5DL+i4nKsA13+Qek5BPOxxU1BmEvtAIi4Tw2ujxVm+HmWWfCADOXh4We
OBTX2Z2qRQW9wiMI407mxR6p7Bb7wJt7z1T3weexdNvBdUg/91BcIiPF8L8k
nOe7RwGwN7rFuKZmE1TT06LkhHUEH9NtQrA9ioiIGT7h+C/izgyCD0DGdkda
whCGIMW19HAorp3fX0c97bsEkNFcww7nw3gXi9no6tjWWI+L30XYD2guuvid
nXxcvsLaGyfFlqKevtnYpbzSBP6LV29wlrCm7saDZRDKU6onBVvA7WhIUvaf
9qqWbGT0Mk1udSaP7rFUFc1bCmZvFRXFzNOp/GljiJZewbMjYBZ0d5ZIoTmX
IKzfTfrUvjPR9s/7P18XaVataOP0qeLbdl0Zv/LbPJXZMxRX2uzcvstLQSgL
/e5p4lCvTeaxc0Bgff0H4IiAOX89DAVGqmUTgbgqME5ZLyHc/7++n9zL8Biz
7lCMLef04p2YzM+/MpYXoERh51f6pC2NhUg6pJD1kLVxfB/PqnVcR9y3jtN9
mT5j314oaz2F0jz25MBnCDOgPRi4JYfX3sjpMfADNuIKbws7SiUsQ2d3oZnh
FjdhArvX8ah7bimftTPPI164l4NauntkjFQnI+dSQ4XTQe+CI/BsSeef8ijG
Qt2oIDzFpn1F5XDYaK0LDEwrTxjG0cXTZHWSmW+9SnmIub8YDWG2W8SPL+7G
mMJLtOfNY7TY+e0c6OwEIAfsAV/zXRXYNPjXWu+wXvx6mElW5XUvKbu1pm0O
btSH1zhvp08ITCoPt2/RQy0dcTaXu5RnaqUJEx+DGQ3Zo2wGb9YlXTwX2+Na
mv9ZR1qhtjUASntopGpj5kuN1dK+11MhnhvtiiR33LQLEKwWwmLK6JW6fjdn
BLWPIZ2xwdhIYE0w2L12pcpW8ZwdSc/8Vj2ssSHAM3hoGrVIy9oYfbfI/0FR
6p8aD2lZHPAdMPvHx2sr/L6MaCAntdl8L13O2g1wmewnmziUbdMesOuJOlhZ
+vrqeaF6aIvQsX4+UUIu3xcXhH2KThi3H/iV//dUZGJBuROvoGJw1EmunSZQ
ed6LIMi+eF+YinUq1ncpXAFrwrevlF+1IhU4b6Z8xEAGgGZ22X+ezfgkcTI6
fWN/qDdGC/PQX74dgirXOT0C7qgvXX+D5gCjw/uXZFYkvU5JfHuEMaoAwjCM
u3jXWj0b6EJ3so1oD7UGZVwpWoeEYfxqcikZPpe35qqMGk/5NNuOxesPT/ze
kxB4PRHg0iZ16cm0hNLiJZnH6ZjBOamszPe+O5fooVGojXiqkTWbscaRWQtm
296d18Rylb0CWPL+K1h4PTBQcQHden3bwmEEMsBihTahTZkzxFCnJp3/ORfh
s13OKEb9VFA4IZ3FVpY9XhRUB0k60xrdsLwVm3l8SXBE8b16ieRbCifsRnsB
4QArYYLfhP80FSsE7qXl4ToInM1cSUbWnnqYE/iRtCsYzCJEeGFGsmWMxB2u
I6JNq0iQNSCBa+yzThBzZedKJbNRvGiSFQMQIrsxRtUDiV4cXs4XJxvfnZnJ
iYxxi8AqMHnw3pGITIvLnwXgiZxEwTSE/xhMHxU6Xc89EAT1PA0ZosmmAkJd
dk4koVjQ/q//vx9rQLVeNJ4IOqv0qpoOkbKpKsxjqvVnkTnPTP9JRqow98+o
Yz24LXb1TzK3O9736UAT6xb4OHawUSRaIChXuunatnNpYbJ6iWkCbzBrpX/P
2d2HMQF66jfS3S9X4cGMPo9E1tbY1d2087nIPa8UWCTnT6F4B+O+tpcgNsqv
Udwf0Py22G0SwDwhAU+6UY29/lVJj5rO12O7slkkVHtS0Qkd4S+dpPJ75v4E
xrDgGowv2dtZg+N5E9lolZqhrzVgPUMi1xNd6Qz8Q4Kh5tuVLhwqlH2zIh5s
3FLH1Bm5H5m5WkgPE8wo1LVt68pPHSVZFcmdeD0XswcxFr69EHuANBvh2Pyy
pwGF/pp+s92YnaHffBt7w17qJ5r1/t5m09YcQ8sr/J7VBlY8Wh4UeSReJiKv
lH6/hU6m61RoGyGnMOi5iHBiaRxkQlDYFvouSTOqOLi/dRqhkyg/3pHwtB0f
4MidwfxztAu6Y5xsrP6M5lEPk6sVZu+gP2rUfxaaE4FubOFyi0RPCm7j5Rrz
ZLyi+2tzf/0qiXbyi12Rmb1XhpTj1v+XjRCzG6rr9pRzas7d3M9I/Q5Od2wO
1caX4j9zYfYvCU8Ud+hfqfB5uB2IZQzkxclt1yPmUbQxk0gObknZVox48ga2
LQFZIrVaePVTPxyw/PaZz3m4DgxIFOEE6xvlgzlQUqK977i6Lc+mIYcPHZ18
y72D4IWEgLWe5CIvQlMXJd2vMTAVPG95j5NU2rOYP+wuPLWFW++tzpNwvv+c
UWX2yenbleOgHKFxFFYwMKbtYbK3fUwRqozWJnB3zC2W5DNQNrehKzi2lutA
vpZXlis6F3sO35X0hH5vzfsmMDgfuGBLZH+uDIUHWPfOmP1chIF+HmpWCqSv
Y2j1vpj8LuEUxT1va2giRIcGfyS8OoyBHLGK/jaZtIFAUVuMeyixWl1JL1FM
S+iaLdrNWnE2bFF8P0wDW75CfbGppye/brRp5u7TRI8jfcvK+ackEM5rPI18
oNt6C0EkzQRYHTs2y83vBK5sPDHjEvvnB8Ld6upQj/rUn6mOtkSsS8k8tKyf
hlsifsPgXsQwBu6b9FlogqVKUYyl9bcQ6w5bQaOnEhmlkDfXCdBYxLFtZmZK
uH1tRc4egKoiX/P0yyiAxWXtbJ7KYpe0bWwd+xJjsjURfsHXrXLwFCg3B8Uu
kNI0AkkprjEA9Um9ljGaWbHvlKI9slj24icD4uyYHGFuwWndaq3GjllcktD4
ajV5BAqP6AoTWVa249Qcp87sLqasc5h10IC+EfbD5Pgpfkhw3meYFJKWCrJx
N/4vKqKUPLHFajbs/Y3SG9TLLz9FCHrvKWXQk+rV6JYGWsCWoBLfyoVCMIHC
rEJvfXJF2lUa6EYxAlvvi5racekSX9vzl1AvOnnTYWWh5zPtR3MWx9gtoRvY
5P2XWo9cdx6ECE4YDAOcyQmKfJEqT0y61s4nrYr0CSctTOqUTBi7qqe9RmvM
p4/nI33TBqW1tCU/Q4vp3pSq9s6CttIPrIJ+V5eRUe2M3XBn4xFm54Z4hD3l
H1p2qqSWe6ULM7/GuRkLE2h9ZNRIr/zrv8QjZpqDq0NXJObT66U24YMvAFmj
zihtduVdpUcJROrP7+VaWktRou7+zGUNl0njIpZ2KWQ71pnP8D+dGT8skXZJ
nTq+o/Exf0B6kllhBcWuR9fZdTS3McDxNUVFXt74ws1C2wWDmdDcdiSk9at7
MQeYYSg6ccf1PcaVGFAGb2HDAWHEbFln5lZ0JGOVryicTckMjjEpltNUpa8F
l8MW7oIoe+wA9vYxXxScGyayDXO6RUo5b6E631t2AhoUV4iVrZi/moiPiKVg
GWjYj0wV7hl4CfsoA/fbSwjwh4Ob6riUBq4KYPBxs/KW+t7/wF5uOZgb8fZf
Modyzq78dTY+sTt4u3KoOo4Yc91HreldnM11ODnirrTjdVo2jg1QkdZDy9CZ
OqkgwLVbmzgVISz5dYP07xC+uqfPfzyKi8Mr0rAT9Ri8EWyPq+H61MNV+LUp
vi5ppkkoBkyAggiYZXmE82dABCUPWN7FU8aBqvdyxjVAKYfYaP9JLPKKvgQl
Zzh6Objko1rqcbychFhEXM4kfxnN5B+cRg0Gd4Oxd4Er0vbOOq7rY58oS3LN
txDyGNk/zfYqKtNsPRQV4/e36LtuDELrN9rglc5Bvm3JYKOizY6uLo2uD7A9
dml6LocA5K7m/+YT8Aq1Vx/uT7oZSNSFfF3NaCiRQ1zcH3OGnDXsluc+RdZb
RRUzswUF7HvVMrhi1Kw4ERuKY7oURvd02VjiNLS76GyDPT/R+3uI/egucJNW
RNqjrbaSxB0lRuKwZt4ZHvnIKceOg6i5dLCHQt/JGYXbSD4K0kfa57qkqqEJ
0WtcWb2JTQP7aOhIs1MVxMyBEKxZ02Ry/rzSRq2RWRMJ9G3M+Y1C0zMj/bao
nR9iLtRJqUeb+3UjYHAG7nSyRg7tanSsUoaEPI8PvD6Wz5wQTz7KG8Z+/nM5
nQADBC25Sno/5TK1PiJ3gpqQR1/5PBsrNyss/plijkOFAa+Cr8wDPPpoN8ih
K3dl3qm9oOiKyUxtUWThhvl0SPTGwiICtI0Rs4brpwDw6fizOakCh6hfn3nW
fk/2bnU9rlVCDVxkw++SSMxdSLjVU5EyjbQ8Y+Pq1enrgGUlRblvg8pM34l9
2s9m3x7kUdfbucnqeF6bEeVjA5CmIr7U83g4eCb7Kqu3n4p9tQjnyhpzfeJw
o8SnUvnee02t/YxW8CT3TQb/WHGig7Ptpf1vuglH4CkFcMaDS0+XrDJf/czQ
BXlgb70x29a4t0bSqipCr9vNGZZ1u0GDyHbGzQiv6M2uI9TZN0+Nb2wgKBlu
E+7PQ5kgFLEMuM+g60P3q9ZWH5DYQ8v2AgHtGtXn0hrgMLQVzBW3NEne9tmp
+ZqWHsHrHZfY0IIxANT1lq3Uf+E8PLmn8IMvI2ImkDHkkZx6Ej7mfy4Wc8sZ
uvIWGBiOGfAcGswuTSZMJEn8f1iGapFBFgo9hUrFeqAtJoIbC3Z2wP4dSRam
3mLVu8VU56RkTSJkpcfQGVVSGe6ZjFtNOviBtpKQ8JGELyidjo7qEKjdgXJ9
+4wxSdy4IaYeBoCHa8JzLzBw7SprvmmCzFoCElOc/IcBnKJV3btuVXS/8JAl
NuemtToKGTf4EAlSZwokU2OmTCmmwYGeB23ifChSNtQLrrsf9+Wm2N0pIlGV
f38ZIfrUhwVRZmiCRmATbbeF4OSpVGzea641cZTgphUUVzJUWDBPY2eGxZfG
p+m/+IoJwmSW9lFAL5Y1C19Tf/aRunmNL5z/9oO8913N4nCIA1G4ow43WX/M
jqWptmeHFHD1Ee1HfDt9xh3nyZPwhjGwhu2FVoZj4twJCXvRHC/C1UtnZGR7
I+L/x1CCQkXXEiofHwvE6NKqnQMb4FNht4U7AoLeyh8AeJZmo47VNKnr4RBo
7yZCc6Wlv0kmNtVmD0nSUfS2fTVlZeM0cCN5zHKAzjrK2/DcJ0MuVSFWl0O5
gy6v/nwMRLBuwHdD3xwWxVbCrcJgHpIy8bllGksUP/TSp0sAEXFXnldq0K4X
FSmDCcdgR1+MgWdwNb1kxxURGXVGNxZEkktSJo6NNt+bADPQZPVpgnMtwdX9
yu3X8hPqkcVFaohNmT5pCOZMZ3aCVX2xN0tM9xvUvdPg0CLk3dhPc04LW27U
xgexG5VteE/JJQaqSvkzsGLNni5zWCQp7cBSvg691ooZQm9/yeai9SB/U66B
MtJJbhWPW4AB8/yDFo450HXCDfcHjGNWzYt9yy43KbmGs17A7x2mlW71OVdn
LRjxbHpYMc+bc70NSu0DbCicvEFTM0eWugwF+EWvU+kULdGMjpRV9dqw+/S1
Af9Bk0mLCk12Y//yhmWJnaEV8igwNc+4Hcmn7ktJ1uLVMbGrfE40ScIC/Z3z
vt8i//Mu61n8etojlJWB5xW92fHN/+Xyoe9mg7/9qW1575iUw7XL3u0WocYt
ewGjgWz5g5vxMbSA+23e9vnYFM5ANCf/49R9szTSwkr6A90z9a+9RkGDsPfK
+wZlrImE4rdH2eXcQeUAS6Xs/LqxIBR+p9dLeXEnRzIMYRLncFQ2IBx5tJ8v
WETPcwUH7WyhwIJ3AnwyU1x277jHXcAA4r/EoIgUxGYND95nvgOXSUsER7/H
UiCWdRmWtpgOjpQvFY1z6GUkRYwKS/jBmkHDQRLpJXdd/7iSKqeyChIR0DeX
kUWMkWZXJXUX8by6WewXCcD/67k64X4zyAqQdordF0n3jOqyAo03uyiCEmUM
atSu9795ckm0G5LwyghwFJTfJZX/ODIHepxi8DE+kkujyDVJPVhe69lKsl/C
PTz/YYekvDKPIG9cRGlaQPLE6owbfUc0vZRXQcFXEceJhv8o8hIRvEyFd2SU
uk3W8f1fDH9p5rWs4d5W81oHj9x1GbKEguqcUlP/26O+eXrXXBRQc2GOHXtc
h3Qrv+6cIaQAdMzIwZznzmocHVqZtPXCS2l/PVYTBZEiWgLHemeR4BRQplVw
IbUo1g+ffSJ4LS7UyuHbGtbIEa7QLyeatRu/n3TgsWobM1gp/wnSZba1H9KB
46n1iOrqYj1fVk2B4+FdPix6Z6uBSSY5iQ74iy7Z240zTifLkw20V70f8xbW
+UbMFrVN5wyoIPw8VqB3Q8dgLmE2pxkr2pz/Q/uMX6x7IGVtym6PLqUAs4lH
7Q4ZXzhR71zmrvtyCxZi06yh4yNtLoceQCAoCQvcOLZrKPR2PN/CsJp3+c43
MPkk0j2WHjZbZnE82H82+VoGQtVZ8gbFVopoPG6gIJ8bd9KlZZ9vVbdOK69f
kScVM6fLP3p9gDW4Ws8uDs/FvRqAtANz++GEPUM7wSRfkZn4l627ZYGyDyh9
NEboHTkVpy9cUFhOdceVr/DcfPi1oLPWnmFVbimH2ttB1NU+WdTToGQSDasP
g/+xTu/NnIfF6hgfSkaPEqcPpO1P+9o7PHqh21oTOYwQG2ZnfAtLSfUXpmF8
2SbI4G/2l8A/RsHoA4qTwvtIxWGknRxrjjTSatM9yczAlY/039Jk/BFtJsO7
ccXhDuc/+TB3+CUU+j4y6ex/X8Mr04JlA9bN7JlLn1qKJGOYW02TpnYRAq6B
fTKmNoIj6eqpWTJetCjl5ULuokRTes7OuiKUYykyGVWsFLG8zeAnTCb7ygPq
Bc3HVtDHQhs3ZueZZiEUsKKhqGBmM/3LMic65fixfbSDNkLdz2HXCdKwHC2y
lpgSiOqkoIxyeOCgw5cBoeZbjiVcp0fUgHnUJOsQUEdo3EH2anxymXH8FCmZ
T4furMJBrVrRxaN0GqXa6uewb3ePkBF+oop7SkaPZ6A4YQLmnEL4JAzRc+Yq
da8xfiekcCJN7xNdJz5ThPH2b1o0/aL/IW8oI9AFcxru8TdnS1Ncu5UDs7MY
MFmMT7A6uQPDu4+E8Gltf+ocOjh+sroib0rXJjdpiU1zyo03UwIVqMvvmTjV
GvbmJ4Iu+evVKD9y2sTBDYYXMcCfdrFEf3IPz7ggmQj9x8Suk9EAWcxm4kXx
pDNbnjvTxL9pIGXY0Z0XmNW+T1S8py/QeetWUuAckjHqUl2AFYdMnMOdJfM4
3drK2zQXWOS7uGTn9WlGXHgeCrCYlU6twZAamVijNBEoFE+XDVWLcIDBmF+H
StF1ckfqKix9wOkaTCAuW7OMSnX+9P6RqqkFRmQUvw4RaPGXvVhLcX9Xjnhg
15xHlC/N269FgjiuiXov9JCk0wBRZamC9Ip4Lint+cnCIClJ9p0nMtUvGeWv
TwIiFSTkCF0CzyCPkwFhW7mGCsy5XeJmhHXWXptFQSDvWpZz2YKi4SIQvqQz
F9t1MVe0eiC8VvHahm4Jaz+m6uSvI1lZSo8DW9QDcFfU3q8EAu7yPsWu0ZPN
PsmgsiE6N88V7AFZCT6CaIXXrA1ZGEkeOyPcXOTayXu+VowCimZ9joWv3yM9
FYdssNOeZ6QxmnSy6oFk9pc+TTXIZsdh7vI/1eJau2XQCJf3lDTx1Hg5UU5h
RH5YTu2fC5EkUI18XT4BL6R0bIrvzz8I6fLDbghVl7skZBckazWRjAPKvwIa
RcgM9y2t1j0tdCKxynl72gYvzQ0arPl75Uzzy6cjTwKpuU9m2C30SrDc/pl+
Dn3j6bEfl20Z+69rcsMs2cql8CWFwRjikGjYvC2tFgiUITPmUVuDxscPkuK1
6e7oFNh/YP3yBjBYo7EJQmr3UPx74UAAKQ/z/DcwujZtUk/AhUqIadW/6lPG
Jl6UPxVkyCZ2tCO+fUowt+tlP12zZehAT69x3fou1Ra68IVqWAvm8Upo1tGA
QE6ZXbKvDtxOIHlkdWyKg8Luti1eVew4baDwmDJS6AswFfC5jYfVO84hqkJY
rfSUU54DHZeJFs/Y2PgibbQBjXHs26w6brQjt51kDOn7JlXEIRDyYBzDFdc3
4Spw51X+BfuN7C66EyOzBOPUn9+98CAYQLU4hUt2cHwNdtctB4qoKWzjSmcZ
y6j3FON7ubXykRjuc+ENyVAie1Wr0zHkssOfCJEiNxoRlwLcVz4ngyIMh6Yc
Jvx9M2XOoBM5zUXwGwdQ1rn4wueQI55izp6Qn1Pg/ywj8QpAHfGBIzlEUkKP
uKfIf2eto24nM2JSBK2T2qDe+cByNsNog1ElfvciTcIvPz7lTdduejeLOdtt
lCWFE/83qwhzrMkK7wz8l6pUNcRwD/RKngePffGNgBEGG58Q0JukEDAhWR0n
QIIhVXXkPtavWr64ppMs7izPxyJ61ajxqaZTcyJlFLuZdI9+9ul1SNdNX1dF
GaEoIJdhXXUpERRkKDiEtmNnl1+olh/NsxxtACtsVc+0hmjmusORYangsDgP
xypAHMCZSATsLgubqK76tpPAy9qXXowN+m41icsFNmrbNIL95hWn9Co2wJF3
Phqa5AHpuEYHsGV88nFd7olufruK1OJygOOogQfWZMZ/Uld77OJPhGp5SKFX
dCpOzJ2wYAHpBdyeSwF0E1pWC5nuCrITUXOUJ84eMX7HNijH4fAA0FA5ujQy
gYaCGPugGgqxzYoJKMlut/9Uxv1V5QuNKbLaVws+7RmjvdviKbCCu0rYYpDz
MwRrFGSONMX1Vms3L4oAqvzPqTtTvw9nFp+nANszNsFt88QkptA6+1BaYQd+
KdgC7LkyH50UXZ9E8Jpn0/dPDCHQ4YsQgdYqYAX/E2J4mrW66ZhAEZQhFj06
XuVXKfuRlRienB23VLGWEV8hGf77bLqNwL9Oi+AfxHZMu0p3jKXjoHH6GjVp
9iZQ4WkfEIvNjS4RXSfYlrk7Ps53yVG7TZFVfvF27dL+97AIH7+kQfjjvFRV
5jxl9FSTWyocT3hX3f6V5FEtCrim9dIjc2m0b0p2RkdQK+Jsw+aXDxvZO5r7
0ePFEbm7gYXhSNmSauoMvmt5cZFCGbY2thZ8LVsy5wM96LJN2oCO1iopXuWB
bIUi0exve1H17NEViBSiSdAM0bxbwmMkboCIfdMDZDBjbpZlW7+mKiojxovK
+ryqGHxliqdENHvYyDKSb+yxlS41sYswJdNz2h71FXDZxi6w0NVuKVIg82Kg
+8ZHYuvSqisLt6Z85K3Th4CAsPWXFVOqVUiuYyQIgzqM0nynT8630Wnw6rzx
IlsJKcAmKa2FgBPhkOLtlOuiuCEhOyVzksCVdvrVFUBLkQK7n2YLmY2l89nj
AU8Q0JTXKXPKM6mVAageXjTMp9rW/Eu4yVKDlGgmg0cNYT+gilxwuZxkHsQJ
1yZO3iB7Tk1uPyejuEI1GOWp2Pj4DgzXZCbylWyY+krooQnkDeIR90qAF+lD
pIsLti8WuRlOAvpOiKxMevyo4IrvaZT4BMXMIWynC1KOBHt9Q25lWlvGrTje
ZYkD46eszyiQ6U9jKTH0Bks/rhKK4JW90Rb4XNnBs0+JiL+u9SwR5A/6221p
fEXMINaplJYHD+p4nXRQi170iCfmtS8zGyjI3WksXFfH1IHT8Btt7hqzvoj3
b6V8X2bFUUexeVX+YjVlRs8D0hz/11Ot5aDfL4y9H2I3nDJekgWFL20PAjNj
UUyMpcC+6wSEcqRpm7Her6WWGlQnRVFay5u8JgNltboAFQP7THKLuqm+V/By
uyVuNLOdFAwzEH1vjcpe6ygOe+LznFIzyd6VTyfkDNNOg6hdtLoVmu6XNXPm
J4o/weswIgFWqKYnw8+wNJXY2QZ8GSt0x1SS6au+cdhrIUyTpvmlqBL+oCOY
GdLK6i5cnUnhfJVeEchii5DYAbs46hPfqAa6BOeMwi0JixVUaQJDnVh6OlKb
l2M3pgDHDmvbs5l9+6IGzlVhQozHHPaTo6a7eb2UxeoZBy2lPA8uEFm69LT2
V7CbgevzVOjmDOOugeVVpGjRQPbnbyZtVMHBM7x0cCnPzIuMmFNGEml7Hy8o
Q+J9nQGeOmjvyP5/gIRAHIXwrznytq44tn10JQt4ZpQxmx/KvI0kODkcO74n
n/QyvBojhGAfHIjWODFwRWRXohDuuMKOd59EArbYt+/X5eOoDfEhp43lxxH+
tQae5peirswgVg1PgpoLkISwaSBO36sJ1qk2rTKHFqj1VBwqnGbooxlxEwWg
0QrXfu1m2CwDy8X3tf5sL6jrOMqGwuMvjU0oCLgR1aT3mrrQ+iIgmmsnIPyo
3CR7gA6t+OuyoprDu52vCRb+S/ofZMOZmHvU0aoiGAqcyPqthvKxlFGzx50+
GufI1m9/xB1/y9ZN7Cd0bH1PZQBQyIneJqeH8/Wy3C5MWGrq1VfqmgmGXEH3
UxYdZ941tzUKed4VDd7HVsFZ20qjGDkC6WDxsLHGUhuSj6CWa9IkDxftkbko
UpG5zVLHYEPqGNUhdcJJxntqumNZ28VGrQ6/16X/KlwdmWgLrzg8182IKqSn
pArfTcVVc7QCXwB9a9EJVR9UbIxAmZD4BNHEuL009TBD1EcSw3dy5+6DU1pR
PjQWC4P8w8pM6Tre2PrMfIEGCFqk09vVia9PqJQxpv0cBaD/WJs8YGSuevvo
OAd6YD8iy5traTxB+ymCJfTIlZqU8F4i2k7BU4pne5hWLSGWxtuqIfWZZmNx
zsQmVFcFHKBGYUBMNXcQHVrL1jaTijByzKYnlxzaVWhjX2Zhx0VrehtnMsTl
tT+ESCJzP/8YHU1q0tQFjUbF2LHHcNqCHutUSMC9ef3mWv3hnAg1mnKMsnzZ
RkbFukzRnM/RYBccszjuC3QnSan8jE1P6Z8VhG7SOu5grlRBnAE6HN70Kvjt
Q4F709Mhn5eSrv96+ivvwzMx5GiHM1AqkmjycXUQ1h1JzjZzVjBpgmIM3T4w
KcOqQs1BFfkbCSQckMswLJ/pthT7RJbNkGGlBSqZDAafnJ/+BKN21iQXmaQC
Bcpslv+xoMrXCRHraFpfZREtiZRne23V4TvT2iRtUjQzeodewyh07KVaJxTR
8iQj41N2umDhiuGgA7CmIq15RtVoKXbu4kApWYdXXzme2DCpC8tRamvbeEJc
YY08SDKh2fe3zP/L+eyWgN4mSbZYUwrARpSSeC3X6n7STbSm4ppzb1anMxma
Rqcdl6uEq6LYLmrPG6dwDyc7ZvdrzXEHpv+sDvhcMNjlWfZWUU1vL4utqnmv
vlNLmSUmqn1gtNvA8EPvq60dtfGW+Smu2Zy2QSMOiYTtYYA8LJPnj1P4RqFi
LONfum+dtUcDZzy+5uWIozZkBC4rgppVOdUJIfjpN2JloxzuC1QJt0ug7XJs
EVP3N5NlBEH5FGFgDJu1ykJZkqyWsbTMIb8ISvsXTgPqsRsL3yOQiVJaFljN
6e68uUS38TtRYZmCwt8BMqP3VSWrz97XIB8fkkfOQY9mS4IJShD7L35oS+g7
qKMLWzPcDOeI+M5DAx6DJQkl9l+LVzjyp5QJX0LNIJKSbIrikovKb6YLocdH
zDjkY8u8/+unqck8PFSsLa88v9AnOFrzIBHw6NV3xKnZGOmSF6d2Qz24gVyg
FOdcb/WZF1P5FQhT3fTE5PHKA1chfXVotUiSUfuA7i3gVS6ARRiFV8u2jmlr
apFTyA5G9G6V4IXp0ljbFOVreFbOe+du/OVMpfvtfULiAsJzVdDQqJvoT2Lo
DryW2SSToAdHQ1YjOQs/ApLUlYPxvBwQpCtR41BvtGzLNmbXeOcZN+0Uv0VC
kDXRyEZ7BGz6cUj6afgkyG5PTH/n+NiZ8pq+og/DpaFfi99CJ2xKB0uVoFmV
bEw/2Vx/CZpO2XbY/7USbllxHHDtNAEr6fAYcG3ZZ2GkVzEsU8VJugmQPnAY
mUuhRZONMC99kQecMxmordyU7eZx6fDnzgMxkzp3L52QEd7cAmhtTmBGq3e/
03ZQJcAugc1uv3F47NT9N9xr70HQVrrv8VUk4L1m8BmLbMKUUkEm+IpsMNVM
nSezXqNAlMz5lnFUodFgIpgn3SjXBFFCWliQXiU0Cy3+Cij+3Gdq2BcUueS2
c7qHlEIU2o+dh7tkiqVx3tHaWCf4Wb6pEeNrl6GgdrrCYqCI/LS/ZfM7KRck
P7mK4W9j886WLB0rYgSk2Fz9z6UQbK4xaKLsIqY6twzBz6FHW4/3X+uQP6W+
7akB7jQUE3D+MZcyeTmle2selUmMU7CD6xtmCDWY5Uk/6vuZJU6PHc9c40fN
8vyCJI01K3dF0+lgFM7R2Tei8K6bB/kqvtArfpSkWWGyeKHm3ShQm7UF2fod
0OJWYedCdnGkVqMWGYabBoHHe9pXnqG8TW4Nz8bR1ENmOhbAln4R4s52E3Zs
Q27B3aDXmK4FDf2v8VRUGSPCyZCIgwC9hqrt8AbY8gztssNC0LpAhTEsiYQb
9j2K2Ln340IeOpJ+9BovXM1nu6yPUWUd8PwKEwFHsxRfLU7BiQm/WseUi6Vv
5cdxG0Y6Z6jCHbto8rg0rBdmYQxvIrg5vV7gEBr/gO5VEXa46IABf/yfOZiL
Q2rlW3/lsX1ovzbBIgxxtfBflcvGFtyfMdOkCuM2r2ozo4vqQf+XfoPvZCJ8
pb466ww7CN0UCQDR+Ndr8p7gMFcbMahdmkmREjfAYPpXYvjroDjQ/8Lkmko+
aNLubY83Skc9g0AhsEXGY6m0w3MyWr8vWhyVKLJzQGM7PoDQi0eWNjHAgJIs
vFc8i4P3iqm+d70XeBoPWZrLhYPA4eLCTkK8KBJGO2rpoLzoaMsPtuhU20a4
8/fobChMLQK3V9BlKL9vg6z6Qag+EkQeowFToIN9xsaA64U3yoNwujM94NTK
cbOWuaTQBFn39dTZd4gpM6NzjcIicI4AoeS5aWJjICo3xaHiLzgwv1VQ63/y
a1ZOcJmYj54E2Pwroo4/x3Y/yym2NNeO3Q9mNpd5bR9msp6k2AgyuQJMhxaE
J0n3oLoUgB6HKaOiGWMTkN451Zz7zBt3ydB4WhYXCQMy9Dcl2Ikg8UxC0kGX
45JTjM/gwOOUUdX17p+p98L3WLHPN+z7tdXTX7ViU8kmY8wiKMRzQFp76tA4
eO5/BZLDV/6oz+Fn2DYa3agvjPvJdvEhQJVur++ZbFLYmxCLVG2quTalAA0t
6PQOYbHfq2nRB2cedkqim7i+pl1M//uMUXS7iOIpSdjsbI5ZBayVhqQlkhgO
WX2W+8/j/kktqO/gylShTgcoNlKa33vANAzxgMSk4uKk0VJgZGJ4zt5P+6ZS
H8nSdpGwISuXdVgnKdC4+CO2JGGUpFcSI/8Gd1d6l+mm3Ye/m5yrdGnGF8+5
FusJinY2NMUkzKKxgT0P475Jabyxap3VkIoN9/5UmK14F4N6Tzo/c90HzvOL
kFgexTTuFc47cUaekMZx3I5DhI3peiRc73Ok4urJxwaJeBtPEkOSn+/CA31j
1T7Fidz32v9Rj5Jx+bFOv8HXCwzCyhqKpfboTnWxkVRVacfn0+r3bNVhAOu7
dPphVtk5knIFqchzbwgJfQotrpE8welt7Ucq70IqLXof/e5HrihfsVBvo5y0
UmsK+ExuOOaU2a8H/06lSZazJ6R2dr3Cai+RQ7QdnrecurrkKn6USH/XsRvd
XHCKzzbUfhdwoYweDYXmiYTRoCf98HeA2ZKjB+rOlI9dPA2cKJl/+wfV71b0
KHJ0aoaAANh3jgGpmV4CssmbapXF1vNOY5YdWSUthv8SGjuu3Z0cUzynEv+L
SJzovED6D8AezNpEO5gAjOzmQ75PFndjqv01nP9d6LOwu6MjO94ro2eHDRHH
/xsowzoYmmBalrP3ucUfhjfuURCKULN4vsNO9cxro04j8qwilQdlVeH1OCmj
SPwDU7F6mX1GxMBMxjS/aTqz8g3sHn8Iz2BAeQqhBB8Tk580BNj5TPycIyGc
podebkQvLfIAhgP7LgVVI5WClHhAxQ7K+NqKx1ycrtqbwnvXCVu4/kpcT1EP
2fjkkD7z7ZugcdCQ2DFpKFyAgmWpE2dMQPDQ3c+vliZuUh/rmPeyB3U5/HWC
KcVmDrL2ZvpUWKVVBLUIqiVS1jt+/oOJc4/uwzH5vb1ssmTOyMXJ/DrJBHRY
y144pwc/3MDjRS5ZeJ325eam/UVoH+j4J8kpjgReI+g9vIJWZG/2TNhA3w7h
qTojS2YrhClxybh6qag1NyK4sDRyWscos0TCeRdxoluu2/tRKYWZwV+yhcpv
8gncxy2GtPx4RuSstX5DweYX90WjY0WFlIrPKMxj+9C/SMxNyYwMHNk8TUG5
Jp8+r6dtq9ejMcxNmTnJVA7dgzJ1289cIqqQWCXAUxAszov32SLwlXnO1hoO
Od4TP8r7193tA98HGGfGIFr7ocXeypYnIehkgSnsw7pY9YX8R5gVuuPQOiTH
8J0sbgtMZKK0oPq2RYJJZjMMNM6BcKrbYgrLYNIoZBktSE1/CTQjtZ+BOLU6
25kih00qMwEsctfka9p7rZbrXnwe5XrD01WxNLKKYnsq4KNealw96U8tX39f
nZ37/HZzgRI81mksgeaSJ7dos5mu95KDnquTY+Az5wiaLVdzeePC22r+cUJO
7E2UyBaShuCvz2QPw2kAWNK4uHscNYIQ/73PHiXpWGHZtCZfInlW+usDuaRs
25Yn0kNRxA2cGVQnHYcGJkmMd2vAsPrJCjlTe4sM/7biGIMYoOPnlAHhqW6K
DvxrFNx91RNmFPn3Rq7qmEwcI7Zriz7ukLGrEaRysni7Rhg0DhmBG7ZzUrlm
JjbVNFV54FK+b5ijUlOs3IbYYHodWkKtGnRswhQ41S/zcHV9ZKkgdiOYehAa
RYr1xWn3wtoCnR5ShsWc/ir7Y0voGYJyagoJJ9SyHBh4IOcpFngV6ucz85pJ
UO3oNuvluYOm+Y9wWAKPA3Y8M7VlE/DkOpDXdPqEige3a+TPwpRXGyvjddgy
B+FgaZQw6pBr0Vx+l8bB5+Jjub7ZATc2yUwm4ArtnauZpyPI2RdHqWTbEsfP
+9HBwSj8s260B1C8C1ttKHf19jyhYvnkwM7LQ70JqVulyM0eVtr5OvQzd3zM
oBWHGk2FCsuOB3/wZnhUuOfjF78iKAaMaaxB7MtA5yvLivIr9XStokEwqmef
2ZK5bQnSJe1BLb1/Z+CQNVS/8YwPNQO+LcHyHkXOcqOzi6IgI+1HGEywl8WO
Bm2zQfrF80ejdDzSeeaFlfpuWsGHiOVfWXFSFFrgRKUi3hLmOVy6UujONkPS
ROLd8QC6t3LvEYYvoUrAwK2ipeNO7NDiiiQbBjU+U8H8JII7AEzvim45ol9D
u69VS80NioObLyA0jrad1ZvTkoNnVnnAJiWwY41CXmIAAdRfb5CLgTeBOiPr
QzPNk9QjrX+UgBr5REN93UFk74GAIT3GgmVkXR8kYo+OaWpST6j2jUBsxAoR
WD38KMNfw4dqagtOLMZjBWygRi25cEaiEA7WDTIxbQenrTFiouxp9ti6wgeW
ZmsmGzX0lBCMGzSH32FDGcF6R4WjDgALrHiRn0yXOBvg7j7ywhGfKqbEHBTn
TBK0gOvsG0Dc9Ru/K5Z45rtBb8a4QOu/+jE79NNSYSg5IMY0K8X8+2iRasFR
PgYFQW+rvPDXRd+KaTgn5jAN+DJU/1yHsi2naJ12ZrAvtRjjwPb0VvAiDOVh
2dY8d3zL9YGZSpkd2wlnhYIIpH+sirwTL68rBXjzX3xBQ5AXCGA9k3BkbkHb
WqoY2OfsMhIqbPWia2WM2Rgq+My9y8DP+bBS4wLVwnH6CUEdqSzkTkLXoxZI
JUFOpHKSfMYXdOXB9lwxO/VgBItq61JsymUcG/gLcCn84Za8hTQKfA2x+uEb
eiZdFa8KBTnQmKL4Yn/PZ1WF0o6ciPy2M/hSD3wuAFUiS+qqcTziQWMp3ZcF
bXwWQNPK0PQVa4Rc15Nr+DCuKZydyt+cGgNv4gyqehk9zpovw+EUuQc9kgAM
cYR16a4uI8lhRPCFKbZajOoddFSb9RWeCoPTi4r0nuqQGO2BNvHjS8bv5DR+
3nMgUKhyo3sFE4MPsjw7RVx6RmN6iceVkGZIfabYlt51VWU1I5BXp9pYAwZV
OAyDJpuo/R0qaXNdqNW5Oqe7ph0yNsdcavoFrLWah0yV7NF4X3fCXvdu9/Ot
XUxgUwcl7KGYsqinBLXSrtbusWE3kSHXbjvbTkB/bBPAMNHTM3nGaLw8htuq
aRP8skKiBJqPlNHt53+RK44wXq5uyavGLhlYLX2O1rytO5DtWSLbFjjyATiZ
yDJhnWxSlrbpC0oVslRzVQYuKuAQeA4rYYCCkOu7Og0OqwVm8+16oy/ot1W5
vgX3p4d/2sCYdigdJd5LGo9yuU3u7p5/AqebHFFgjRX/p04d2neJ6EISsud2
sC21rPJOHi0LwIK3yg6db7rKl9uwcsz+wKYuM1vkVpMkIUFbvM0l1DajPLlP
YumnDojO2PDodpzgZmsn8tyOCfeJ/ceZnYC852IlMHy/+H9HeH2iKSMxZk9r
leV3WZItB1SdaP1UNB96/rqixH1cq7OP0k26C38mtk2ce1+kEjnUuOpScvNj
mzyBZe/y3XuZcZUZmCLLiu06lejryMMbQdWxir1UFLHiz7xe+DQI/9ALs4kY
5N0atCUzXcsMOZIxk/puVdPOQKZq1t6djXOjTN/y+aawTwV+c6DViHvm9a9n
9wqy30lgX1ffMM4qbG+UO/YmGdD4mplYDsXhWxYJyH2W6SXFyXyiyWDQXBfj
dFTOCeFgOCG5HsgTzPuMIvPT8rwelNZDXR8hXUCtWPx3vm8wXZdMPMGuspKw
Daz1W7KVaMvAaaAVQ9arIZmO0FkAYZUU9wgXnU59qH3YAU3EgEMPOhCDb2UL
+itV18BgQcBWcyc8EPz9NoyUcMQFQSDpG6oB8+3WIz63w6IBsNd+AdPOlBOz
54Cz0Ou3CpXTsn3DYlhJP3ze4Z5sWHk2DMd/o2XLZ2vvATZdOO9aoXmCDc/n
lJ5ClEp0qdcLrPjrz+ka4HxhL2gHCH5WLvYSLEAyB6E8HQ//P3VCxWvcLtBx
iUd1bQGOipqmOO9IdGh1KIYxC5dZLH43TZWUk7euvqF8FxBXWjwB6m6mXr5J
t54I2HVU4JkWMVRzituTF9FUxFG2AbWA8q7HkDy6RfKkdHAKnJh7YyH3LBlS
d6MpUgXbZbtwcxP6diFWGJGWxGPLtCs2Ip6yIetrB2xZnyQ+FY9LqImjWcD6
b64syEAlJtadukly2SRlLuA9NHVyw/kmCaoQH1uSHXf2Zc6VBjTLWl9CrBsp
EDdYDQ0DBhj87qHH8telEEXNRjJxVoKcuKGBSiQrKlQZDt8w/s27tLV5BM0/
mnzV14qSrOHDV3C4QjmrOMFHR7TctwsmR9glFgQMtR+ImrxUOlMlbwm9WafG
abT/YnzOV+YLJZljJ+cgy+m/cVrY626fvIE8zd391LxXuDvwe6LG3e55Ps+m
rAHk3GDZ/D7IuOY/EFifJBVLFPnt0sOwPzwzJnCx8/s17N7abYphrsJM7qiF
DZ77QRbupNwtp7XAeyTWc7MsmZXv9yhH9hwBm2ImWuJTj3bcXkzBRoNNPFKe
dYzLNKC8AuS0723hMutELvZ4WrxgB/VoRZbj8AUKVdNeaZFOosW9OOm+J2Rc
eWbTW6aarw5MxSHElnS3iEI0YoYpcgjv/PuSJ/VtWzP+U1yHb8KR1B2Rmkpp
7+e2uv2Zqth7LgkPilY/6B3Sqq85I6PrOI7YPx7DYqFMXqIB+lqOa/CCGjoC
nkx2PwKmq46QgoaRimo59C7m+CpJF+HM4pNhCduxyFGOh4LJFN3IU0nBK9D7
oIoIho8LIce3ED344/Iwm451I0NW9BzyQW6COPdfLnxIhuz5g9IB5gDJFoAx
jw7Inp4j9gOhajmGpYb3Pl8LRmDKkV/b9VBRVPvlActEFEr+4tSHFgDQx4nX
QU2x5RU5yoGxN5auofBl6yeH90jxoL+eDEpCRz91efdj4OxnN1SVSPClhB6E
tiRCHSV//JoZnR9g+6PgGoWMz51DAZ+cQJppCLdBKwA8RF5NXMqTtP29nNv0
+vLmtKmmNtVyuf8Y72k9Wc6sf+LrOBwxhO24oBSUgFv1q4hybAU7sKSE5Vfu
zrddlUcPPhQZH7BiIavSGvzGb7RSzHB6/H50KenHd4nJzJaX/r+ffKMcFbww
FbtB6bvbrEYNmX1AgQhDhC9g2ufP1MRjc7PGbWmYtr11np+BQoDqPLSofB3X
iKlvdRuPsrJ24y11RDAL62zjuZJ3FtMv1tQ7CRVdOmHE3Nr7wemnoZ+8xi6Y
aXYRhLDTvowcZ9DhpM26KIm7FGqsCVhBp+FP9/wJNxcm1zrLH8rFOQ8hEXI8
FkkpXBgk4fwEwchiL5a4oX685MRzK1Iir6TpNtd3NQMbJrLhpxMalEoPFCmp
GnBszv0KpqZcCYCSzkcbfzL/0k9Be7bAlm5iiZH9Do2qjinOFbdgD78tG7+L
hUaPinTUsUV9PhNr+Mr2akxdEikNd5A0Ihk8oiqbEMRUKlaXf/u9Z8q/mPS6
FFgk/8O9dJfDmrXvh3FeYVCp6fZG5733hSet/nkv6trFXNrtJ08eyreyQHin
XFqzLtnwXL6DIs6DpMnU2iwpSmtmcrZ3R1h2EA8SYQKixG7IaY3zydrIkK0c
5uZlpWd0pJ4EJF3si8fLX0MsokbELsJA0nK3uBHZ2sVLOB1TLwB9zyYIIi/7
atd1ttgcX7ALoSxH4GNsvsSUBHD54pB59tc5+QerPfihk+baPfFRd4/1u6dJ
AZsYLqEaDLeP9LZmhBvgwhGiYP3tywlabSa9BQeICAC79XjZKh4PBi5mWjzR
nqi63Rxy6EmRiThHn+zm0YJew4r7prVqWscqFlMEkZBRn98bgaU7UGm9Pogj
TIL5+r97b9qgVArsUTp6mQYXoe8TsUMNDtS1m2i/ZQ4AjNmSHwEmy8irOczo
kgaohvUMxhjT58tHQyKluCHA808enidbbHQZE8ttilVZ+hJLQFUqB3/NRW+X
X4JKbq1YblmREO9LHnPVLOqbVIuUM2faKCDMZ3GbmZRJLH74dvq4wbs2lSlA
z2ROG7pk2lCetp7Q4a/MAchFF4D0kBP4oHZ2O1bWS42H/qsJbpxsFJGKIRec
Ah1JoS3MYz5kQVcLVKvNBfjwN4CENiUrr2vg6SStZbM90lQShm20a8iSjwcP
KQV0GEW8xDxqyWYOEVp7YCqqjh8MJtbFp4afn8DW/wTOdj6uYtHQ6PnwO+xz
I8/KPfAj/AzMaKR++P2p4MARFFMCQOtpWBD/3iI/sZWN7zybWQyu/OUHFOp8
d94IKJhVNuDQBbVig3TRYo3wFXZZ9+fnQh06vx1ckO2EYKXa97oKh1EshLxf
FYBcTrSoMM8qQrgyOKHH+cuYGfiF8/bAZM0EMl/PwfzHo/+v83W9O/fvXkNj
WOBZT4Ca3+nrnVXoTiS6IgqZ6j3jt434huvB8/vuLHqQKdyRuAFTa7oOv0ed
AfU5ba2YGFlg9rPrk4qvWGDs+XQE4AWtqi7oK7a26v3fy4SFt/RAH+vUKm/e
UJtQN0c8ib4aR8QFl8sfOfW54gaNa4TilUodZoSEQOvX0DmjGW3ByLE9Cgp/
fdUrpU40TlZmwk4l6D66GW5JJeEQ5ZLaFMw3vFB0+KYYpdO15q5K9GaG+rGN
db8Fcx7uO3ePhF5eOEZTc6k5vGY18dWYu459+DlrpL7ZFZi30tPoHNtkWPOa
bB9cUDyEm1PzLTh4j+idCsLu/BF9ySuwaL/7FmUW0XijtqaZ8fzqwJSsDTwE
s5IFJWQ+Wahh29UqWogwoiRZJa6VOL5sO0jzmaUZbgPWXI1ItaDtOoyO1QSO
RZ3GzOZBvTaV2gaUXVNWyJEgj91xRMukdlWbHjn34eMfTrBSNm/ZYOd2WAos
u+Eeb1sQo4RNM/t6A2xGi/ZV1sU6Fb3Tbl/zi1agyT2M+SoOYaYZ1fFFYEU/
UC+rlU43IwpVvx9ya69HPZkoYXkenL9ardpddiZYZYevFGZpEmnRmEB4lQ7O
AtwoSqnv9ap97wNPbLn9Rgjrb3c5mg2ePzfQ60h/rrpIUmVwlh+aojhUIcZu
tzKmX/zMOZoaCmvt9diFL+1uggv3+io4mkxTsc9mOk679KUG1vOWcxH4s62q
Al/UP2hLxEDh8dZnb8mYS2dssCQzjCAtJOqd/gB+Bp4LChzzv43z6n8YDB5R
bXq2MMGHIRCWbFfgZoogt6268C1kRaeIHu+f7roHX7PhdDBQ1+hN3+G5Q8ot
unCkmBvR7Aq4to7HmlZpAuChZ0YkdpJui9JQxDvHCMpWONQjHrn+X2C1TIKJ
xVLEsc598giph7CwBvZ/2xjLykmewZnlpXLoL8Tts3UJhlnd2Jy8Cu2cU53l
TncNwH3Yk3fXl4re6WVlKUm0AQqKjVcu/MXRtQeU0STq7zrvgkhXa8cLB+ME
ImufvssegDC7TeSgIQJPLt69oV0P4n7SXXEkOHWzgGx86bGZBOx7ZzjcmtzT
lVgKQSHH6X/Yg2RU8rSO5D3GXjT7MOahAGAjaZLeccsu5IzOLUmjAAzobg8O
bbE5rbzvlJJI73s9tq3Twt5PJzRFJGwPqrIFqK/qlE0uaC5ykzRDSEghPytD
n0GqTTL5ek/5dzaBiC6gLR5mimeWHAMz3aGG2uRVYNp3CQip7w68kO1B3Lzg
y+xS2AMW8gQ6eOGMbnecosG/yjr0mwlUq8uGDdLQOnYYmjUMY3uXk69SDzzq
9pL0jSszRDPJH9GmB6RaMAfEfBe1llwDt5zBZG+M3j5/FHWo+d3qa8pJuUOD
CgZje/emtoiZuYaan4xRGaSCpxxtaZJxKOq+ZSF4J71YTJCWYvkYo+aIRLWi
HW477wGgqwO2KWhUVTh2EP1lP4WEzT7ORMOPsChBesxEZ589YyXf0xt/3chm
2SsCDl0ougQs60uWQ80XxLvgw7LRtbhvcd6PjfZgJI2NuZ9f55eB/CxyCp7P
ivP62PLSD+k5m0UyzfIg4pjK6iazrLnQPppcwae8ZZKlmrrOddR+Zu9vjwUC
neDl9AZD0dCop5rcIoEAZm1Ef0VOa1oinLc3wrF+kTihg4P59QdTR6paZTK1
7NR1LQzgrFQknba20sY+QO/ohHEamqnh6GOMvEbtSyX15YYIQfr4FAPdXGZF
hkJMFKpKELduNClEu9Fav5Qfwz6Mln7yj5+mlnE032AiNcdQnpDe8nsoK93M
5xebnEQjCH0lBoAUoCZdqJkhdrXZtHSUKDh2rsi1wd0NkUKSHL8Am8yWEjJc
9O9CO2WPHlGkn+yA0rZU4Og/hjFr7TsfqOHqL526mMkUVlJ8KHL5Y9VVfn4V
duTBaylb/pI4HST5MeI6pf+anOb1+eIdjp6RnDC4aCR9lGIBY+/NpUM7bYvj
NZHEHD8dcMWqd8M8FCTGnBsVGlWtlsk3UsPdE2w9SqWw+vFjidKmreJSZb43
zzS3IJ5Xl9UU3qb70c4rcd5Ie1shW+fHEIU5i9K73giTDOZtIaxx/hY2is1E
TJvJyj6i2/RVFjNcpuulAhPkJKw+ihTGNn+OrfXIPzhI/Sb9iroIgs9uxrfX
cwXuWWuQPwgszPN8B7KW4EylVf+aAWU6LUKqkGcM3kdn1WsCLMUoVizIgfFF
vcZGSGP9QD33pEj7X3OwQ5hukXjqU9rAUe6W4FPaA4o0rj7Zbq9dOIc6Zls+
jpwZIBtuY/YU+5FTOy/dUOixS9tdu21VfDJ1aefr7egv9OU41pyWrixSobnD
XYbsmD0ISVTFZ8OB6/u/n9qWyPB5igLPj9OZ+JR7GCYRO9+qa9tYkMWwXrSa
TdNu01jmkY8a3ff5f5BVwAUCmckl1KLVhNogPCbkhNn4EyQsQ7MOvaSzpIEn
IkXagoQsQzlwKbHZcNT33RNQIXlUEn7IJOm80dK9oTgOOQlx3qRUfSF2CA4d
MEhk99DzE/itN4ve+QNmP4qxaKD4WdU2wqZUbLtOerYTAfpAzyrSP8ZNuvUl
JuLQ1KaM8uh2wpR1pkKPeq7MbDJ5Sae2xnpY0m0csFe8NEBFITGbJdrrq0qh
SrWZMkt5uykew/WZ8637EYUkDZFuDflGgvyfMMM0yBhEXx98/WwzTdecA9/M
GRZYi0xYPCVn/2vU8AsYyFBd2A4849nJzXKfBYqfJWvT7YLjGOLAIP+UaeUS
JxhCVUDtaYOpacXIPdifGD0QLVRFoweiPoMgmhZcZtBR2PisICce8sG3TOHD
yucuzYe5pIlRyPPZpijrmolxJ5T8VQSPdpKcaVzs6RDHGJcx1PkyCM359b3m
6egkgWaxh5AWX/AMhCbxHkbQliq5FmBhRLIarCCioSQs6o3EVi6p/930yH3H
gkcDMbNjW/HnixuLghH50bPTcRya5ZqglzmogD3QjiGH+5rav9ChaGNXf63x
CFMuOh1OPwyLvPQtVNweY32mkjmQtDLEjqKqi1eYoN8ArIv6AjqW6Rp1uZSN
CKa0XiPzfv4RRD5LsUvVQdQnjXaSu/6ovolPPevamuJBrSpALVrVo2k55byU
fNcLA3lPqhTqlmFKpFpYRNM3pFkiaCUSASsCLOsL3YKrhJ2/Nu8S2N+6jGz3
i40twYTPgDX+I3hf78GdEJv0J0/ksGVW7vyYXCBIY1SLByuOIjeikF5d/tPK
nZAN/ZUOxR9erfwPgXzG3H5I968J+VV+JYcSD9SUn6gojTARkPFP1R9+Exw/
bT4w7BCiE1xXTqHFcduo4oBBhJZPRXWOuw1AmWzNoppCib2WrJMLRwr5NW4h
rnJWd62IvCmvYKrm9RW2lDBwaqUShJscVwyf3ID8mKgCfXjnq2JKsc3W/p5Y
I5U6EEYNWtjfhEsWFs3ildD/UwOvjyAgPaL2w0NmpX3CZtYhYOAjYBw70w6b
FNjBhcgkzxIubHOAPankrK9niSLyU9FS0R/mI04JaGtJ6f2LQ0kDWGxl7bhO
ry7xK2jZDswXzk0nQMhOAWkRSGlyt4Y2YJy74LgY3hIhPOH0XYwy8Rgu8dKy
a/nPsqtQfURD8ORv/V6RLwObQA74LNIvGkOTnoryLDKWoJTL4En8zI9LPbc5
yodl0ha89yYjQyYxkaPm22U3kX8NP6QnDc/1lBYX7IovKxNgGC6Wk1cE8HdR
FbA5B0g7SQglQoAcYCXFAOjep54y8JVaNuF5Zjky/2ilGsWbU70Hl244vaUG
vRHgrFL9gQrRGM382WgZBq/zBknXhjMl9+PggGRNbcO03RjGTNu8AmP1uv3Y
BsQp1yC8KOvPEqoVXQukNKq7P+a/0YVFZmtFY5X/3NvLcmIEQiQ47uqoMQ8V
5c6vI6nQeyDcygogbvP5iCKfFwF+BfUxag0uGFvy1fn5UbS+fwPNexVdURZK
pM2wjpAAO1hEAgQ62pThKSg5e1eHNc+PFEarzPK9xxraUAqEuvgVIfqU7DBY
ARbJfxbM6iJUgM5cofCQR3+hi9ZwDFjct6F/Yd8NK1jHw418m2GZxQOYWpHR
i668wFdgZARN9+J0Zhu/7Wbg2+VWgnP10zsEx1y+vW2tzRdgJU4ddWQLyIjt
e6pp2kmAuVClD+Co4cXddAdgo5d/vq1sZtDqnn2qODqsYfcavBIf8H3Z2y+7
G1V8CkEBiL2Dl8qRJOS6h/zmkv78G62A9corxFAxfo2O7m5fzdkwkSSRscBC
MWu17mDdsCkPEyVaVrr6ePClzHhOakoOan0obo2xCEHUOb+sGTDcqrHWQdBR
ibkjoK+2VT7UJeRgFXe4iu+uSSK5Wc5aaQX6hwjy2Yg7xwMo0LPVG80h3/Z2
1eypO2mod2y24sslW7s2H9GhOl4JmvhQJq3/XdR6J2ERk1YkOxgFz6O7gvrI
C0Nqd+Bmbd1gRX9jtYgSM+WduEcrkeB+YUK/K0tFWfhEzGpDUq8WWGL3qhWM
oGhOH6BSEK8z98tltaiu8P+/jG2PXpwckbJJRSDJbsJqnfZDjWlwqp3TEr+f
1fizCZX1gS4bIiahu74KlpYYjG5DoIc4EtWFVBz2iwpkbLzpeDFb66zmzZ9Y
YYdoGgBRp9hIInamFOMIF1mOGCj/ywTWNFBoXkaQlu2rzZqc9R+XbYT4XRoj
wXtyW2vTHhTJtm3uKotKD2+QRsYQp4XvTfptwaHclBLrz+mKguKAzf5FlcV/
5qOdADaajYefwOR3gHd7Yt6FlRX/3NWTwhGxckS8RooNiZoqcjh6rCZz4Muh
ZtKOdpCmeAlP9JgOvTVHjqOJB1hHb+pPDwjOuFFodTOhZvK0N4bMN7Lt7cOT
ne+Q2Txxy81G0PkzJXZAWi4SxdwxifhjdENdRrrIRTSj9J5zb9aznmDhrJRb
BC0ztlWOwieMlPLWBk2Br5VDRBDB4mQJmZn/WaVP2nkOc9U5W8TEZ2Ij/VmR
VxjLPTGw/Wxp6x0vNBzVuRk6oAUQqIOXn9AsgAWCYo2mP0cH3tqO5m5DGu6w
DJyJiiye0btjzGSLuIoHrj4v/Rhx8HgdYMKW/IcgAqanoeDy9jnL3SafR11/
I46PpljDadTkb9ZT25YOoQHqmO/lgGwkTJIpgE2x5K8CM41O1mYYuJlXxJeN
L2/uBJUH7OcRKD8fAURN2TgkMm9ZXsjYO+P4mGj8NA4NASm/wOP6rYuEz5ix
WGIe6nENo2PBpCZ25ytFKdlShvAbSthfIx/D2OtJi8sQX5VDfCIFau08lAlr
rmKkp+rw5aaKFo3Q+cFyCryBuA5Bik8pDb8qYiW+Llys/lF63BMHQU859CgL
u6/c41y1vC+H0hxBX18cwG4xEGrdZ6YWZ2+gl6Gt3/5ip4GF1V0VLzaUNPwp
zAU1hfi1oZXackBZYztr4lEw5dsB1cYg8hkWz2igzc8RGdTjWSHusL4yrJa4
3buIcGVGSla/yPatCoTcMx8PejEhcqbHJwx6Ly3ABUG7BD3S1g2A2QsNpWV9
xtHbnePuPI95hIRU0VIijp9Eapml/8QEv2VYzm6xzkoi3tnWt4t/Nxzf8Ak/
LA/+JSe/W3ccvsKP0W0twQd4KNu+dE+YJPFyeG+2KwddLsuQhRvGyeoOFCIv
Cfcbr26/nA14dsgDfpsRCz2muPy3+Vf7xNVnlln67o7CzwD/yp8BrnYfiYAV
e/j/EitfYCyPf0G0yxVDLTaeXwLIbCRFXcTlflV03Tf/znJjEJp4wFQXEnSu
1YogXnu2sH6ZjGaR5ju/SgM6RX9OWqAM1+ftL2c7Wsh+9f+e//FzcKUJSpza
Sv49B5vKK47rHxaMe2Hm8yaEexsfhEj1FfP5Z5PrczWn7OhBUKUCXytWcpEk
XuBpeJrO1VThth81sqbk49bKVg2rUcAHZXybrg6uDzp8fmv4zl6087G/8Qnh
FlYytuk9zKRQWOMxyqqWgzm76TKpC2Qsdn+FBTBdw6ZTxOR/JGE9Wh7fyNgm
PivYdsWIfFIYO9D16mWIBQ2rdjwvqQbvpaOTFwvDDWPfJrOK/dDQrTZBzAHV
jFZv2D9LUtSEgkSduwl/lbXG7LxgAUOfHTJVe+idTC0Z3m14vR+FYJuDzqIW
V1UvPzY9wF1E54PZ8psqK9BWLiGrd6+Tx07g/K1K64Fy3w05RGxducO4GnhV
qnt95tfSDDLJF31/NYaCFLzhAspDFMYpVS7I96o4jpE6feCN2kV6S7XEQO+3
3zSo9SB8E5OZyX28xGiMmU6HTtD/xfHuHw0tvvaaLKxlt/wZxcsEV/HRaUbd
B/XHD0Yxze18stEFUOMPe6ZObqmjuCCW2CyWEqc/VRiftARNLVRY4Y0Am5WJ
ORmamZHsDwwYHUUKjB5RuUaRDSZJ4g9v6+JehvyJ9nrCFgA/BkCz9YdUwb8I
gp1rWQnNEB3xe5niVYaf3vEEKK9za1AbLUJI+aholmVPGyV6HZVaMBf5+soh
QxNbQJXl9iCnhsklYZZZsUpQOgLKiPMllBELAdhWYYD5BPFXkqw0RaAdacYJ
uwjXTIduCwSCgOQ5o1A8fnj7mgs4Gdw93BF4se4AqqBZ5LRbc4K46UVu8NaJ
ztdWBkpOYWhDfz3MLrv+Z0bFQG3i1oC0ra324CRkhY1foR/fxkqdTfE5qVC3
5ZxWTKaz4napXemBwebTwUz390x/Y/5qhoXsvcG/5RW6O98P8iAgk/yXTDqj
AvDdehTos3GG/+AJ+KbNexIzOGe/PPJPw6Tc+OHRdXIiFe1vAZHfGQb7hILX
dmP3oCoL2S12/qkmCYf+5ZZQkBzM4qkl6YywvxRRQfh735bpCpmPDjEbVYTB
irp4VHG4qA5OmPIf4bZHb1TwjMSn/opD/p2+s2MVdpEZlUH2KxNqx+a1x1uR
HInqsjZQuevRorgYFi1u8ypN8RNbpc68n8IznRVpeKmIjm5oEEPSx/79xcYy
NYMPdmRbw5Lb6nNflrXNeFa3uD6WeCKrbpiIZBo7ENJXedTLqEcYkd4lx3/4
PV2IDQgrroXHEtyXamqUSeK2AOm7wAoU8KDLOIPWRfmIf+VXD+ZPRl+cRpSN
fJwDWx3ddPpxnvHZK0IEOInOl45h59hSXbSa7bDMzhHYWUbgvb62yfRCNsgc
MF25bRlnxhbswEg1sqLwvB+spEUoiPZ/NK01Py20k28CV3/1l9GCvsdzuUZf
w9MaPiN5khD5lnyShYNw85yp9yoOS1GaPH+NRFC2w8nPMHlUZ2Eh8FymB2Hd
acJhdEgIwsCITJsPTRxd1XnnA4d2zQjMBPavRsKoWRLcl4KdvGcXhWbxkOC9
5dkbiipgRAZux+wgRRRp2qI9hR9mzB95bY+UtcB/u4afWej85ga6aeH2ThJh
AfijzSdYTfN1BCvY/ugIyqlF17DmdAM0pXAbmlQBpHceG+9Ki5JMB+EP213t
Oza+K/dvLvg2TUeOdhKJTmL9FKNJmZwUJjkDUCt4sKrkVMWF0F9Fa6Q64V/I
x4rSRpDBXiEHJnhzHzQZey0rAko0Y8nKgbUwSlQfg8CyA3SWHbCKQo5gxuGy
s834C08LJXtsbKYckokkdp4xY/R1JNczTcI4mH0AtBspgvXvdtJc0Nje2H8H
BsmRfKQ5+hMXR5x1poDjNZBMOZOhzkVCBodHBbqVJZF/YZmalrWumVDOa+ao
hsRz0Of7Z0RJJmJHA8+xS/FbeGU4k5IvR4TXJ93tMbF4VmnUr51q9DhGQaJn
7ePVKcEUOLUV5Zgp8iUU1Yce4COJrI+04IKNbhYuJ7XHWMs4//Vi5XZpz4Q8
RLJh5hqVeVWhtxVOZndxtoDMg63hRQf/5vbwzRqH9tYt6iRCejNjOauaqZRW
XtnytuIqDZBdXScvydsrEWG6bDPhYpqUTYrs2G4BpERBxx8ovF95rw0zYtVd
e4/q38nWTh0siThRKQ48Lgt6XJEFHl26VAhBHYtoq4fK9PrZ9pZZtNS0MECE
BVU+I2F41DNL7MRZ7zXWCPDq7eBC6rwiUt81pnShNzfplqy/Qik62f8UlLiJ
eJ8RPeFSkQeILYptv7NbmqCXULd5fiq4hEH2beZS9I2tJdGRC5+4aZQIZY68
ttqVJx8rRW1UTK4M0RMCnYLXXmgxq/0uTLYM6MPna8ssjLtBrombubJd3GJ9
bSzovCEBXcHa1rnSNonQ0ZUp52cn77HZ0l/zEUNvJy0FxBnHNV/7y9Cx3ces
1NlzQ/8w0nA0OfsUlkBOdRo8rU+uF80Kam/qOHpr9bZrthn/uxgwq2yN7AG9
5qTfLhzmcqZ0BUoSzi3TJIj6v4ZT5Ubfr+76/FM4QUE2QrTXYnkE7C3dd7Y1
kJliHSO+iAC10YFiD/SefwcuqXTjb1Fp47A2MuZqfAiuxSAVThuBf68lfoAM
Pz2lxD4GYN4pdQ3zUNpHyVBl4puM1uSR1JnI64IXrfs6gUuS/7hYTUmzqupf
DB5hvsfk9mYZ0GfbiELyMEpM1j0PjDUFij65vIKOlipwm3uBVW8hpGRw5rTs
H1IHJ7IwyF5bi/m8TCa/t1m78MnvfFvqTKaLbcsQv6KnVFiLQmLndYblM3Ms
XEaq4rGQLgtJmhjuLGzOVs/Ue/poua4cr3dUoXCqEzR+h5efW5ou7Fq2xfOp
dMpN2WmKLaVA2vorBX/7EpjzQyQgTjA7afyC+rms0ZcK8MqtubztAIeaSswJ
T/M+lgp4qMgWMagHyiIMhoL6pUHB8wHZmwYxIJHL4q3v0aYVWt8gixuetMxk
dkzDwgJP+Yw0TbJerQwIKBh6vDVIn3LWxzPEueb0dKxg3n2wFnZVzem5mv/U
YbhleBLdAOg3Q7rLiOTtuYjU0VrtmwP0fYlebJi8S5pQOVHefVTuVsWyVTze
LGjbOTEf6esTLaR+t0vIdhL1QKAwWM6Ft1vphwgG0uOXsiWfsMId1DA7B4yG
3w4mQHP8a8rRdwgYS/vpEb803r9KJ0VIRWaEgUfY6HaqPY6+mDvVcMH6tWUw
oF3zrB7Uvbf7EgYhvyzG4cYVOToZEgrXbV+J80AHlzJzTjWkMq9N/j8myZgm
pLJabbof+Rny7ykt3yHgS3zputjg7fUCqkXikp6RGYBTYdeRLc+D/kGuzPJX
nst1azjMRbsq8fmz+ofxrbXttfdoFMwybUOoZuj3Kh2CEmo/f1OhlC4Pexkw
lwsMjGP7icobVYPKjDQd37ujxtUjf8NCsVuK4TqVRer8T2qrWEfRHLOedKKc
O5KoQIbqhLtEKHbb9SJ4EzFmpJa84i0AnzyrHs+DGPsi+vW9yOKjsDNr6o1Z
rTsO+mTN7xe0TBKKTEAgg9dajGysu5xENXZYikyLERtu5bcq7FFT9Xw57KpA
vBunz4da7Xzb/Fbv8ETNazLIGSsaJRNZIQtF9/2yKD2v7S+wNt9YcayQMOsk
c4Tl21u8Rr4pGW2wPPNDKcPephbB8Ys8ByGaYGcRWgbxxWBAznwowPIG7CAU
fhQB4q1ZySnuZsnsdKCvj5BEEq30bsTGGG86G8ES3GlINGV860JwJBFWT5bv
4m55Gmh0dIJwN3TltOFTe/rtEUVjVI6ZKuuFgdU09embHe4781dpYnvKp4Ru
h/bYaqUxYCGCogIqNSx+iCWgfu6T1nNV/PGzid9oXRNVSUj9eMqJptrUault
iDYNdYGxxZHt9NRfXMSSXAtgjUEkCJ0aODivvy6izqJBBpZFxPzudNpZHEiA
3A2l2X24xnq+0tpmGQfTiYGGT8rCdK+GlW97SYrvq6XQVgYzai3cCAXho+d1
IVgkx1M4+rKK4dxZmn+EBX3hevMwa91+DOeyS1AAZ6TRwApaog6AK1G9SVHP
DnnXgYtiaY5Y8hKM4Iwj/sIOQEPsI56ecP4V2BspieOtIaefn9KVKBfI9Xp/
xUPlgWyeWhpdjxNpMsyXAq+i/4VMWEBHpZus9srvXcT4qa9VxP1K8MEiFuBr
yddlhcl2Pk+SU2au/d3bGig0sD8XuEuuCHJQuvBIPB9pKpHuM+dDG4Vtt/Db
nkfe+C0o/SdAOhVmb7AWE+Wp12sOu9V/UnfJbByr4Yyb4I+r25UeZL2G85gy
9W1/MUAuMVgfBbK71YP4d7roifLBEe/x3HK1G/IOXSjGSBwzyaDVlpwrNpW3
jokkanY285NbX+tjEmb0BiyF7pjBpSCdcURPSF8fWiDOmv5Cs3W1CyEcLRyT
8PNW7McFaj/ZDuZWOZiM0vltIDbIiwpOnj+3flhpO7ImoE/na+zOb6t6cq4X
Uef9KJM1z6uOX0mxvqSDxsQ9ljX5l1oBOU9WZfY87FP7VZyFJ4ebU04CAIQ1
2MQMFMjafu8uHdHExunG+eNuM2cDVurVJbGpB9Fotr8Fdfdf6M+H3VwwMkUW
Y5nAVcNjGVAwLMkkGBsOXfNpy8JfQ1kZcoZ3HQb6KFRDKxisiKkriEhMZmoJ
AofPTBfA08fB2JH9ivF25+vFHDF4xrmO/mHmKTi92udC/DvN/crJbg5qhmu9
S0gdsPzHn5mZDQE575k1xsPVXQ8cFuk3jDBbOv5wC+7an8F6Apav98Sl15YX
nnRgri8ACc1hdkz7rJUksp9vWYV23vM6tyJ1bYLOjpZ4UoAi3+YgJvwotJK+
oeRnxJY+FID4QswWgP+qeuWQyJrUYa3SZWPtxbvdIzFYItd3i3lblmsOgr9d
2zMD6i6mlWe95Ccn5HrOFr2iabW7HeDhP2OAV8q07c1CO9qni7PVYzv46Bl+
f9NEBKIunZCGbYsRdzJ/HS6NmQp+5KlGMg8q4xX0cfpxMIoOzyZTPBF4vRUq
VlUVJWAME6rePtIIjwUY2RvQNOPocpugKNzdLHP308pKT88jXfWtKd+rmRa2
lZTeYKONu61DOWBtQqY4JNOl1GPwHlo7IU7oRj7Bz1jozJf8pyOlSkvM5Qbh
SmegYMWmIiZNp4SJc/WpniZu8C3gxMZXapq8CfPehjyKaN++3VkkIBacECTg
ckypQaqLMe8myyiGIatpkU6yNmPpUrf0fnDx+GFLyDOuJUZgXEv7WG7mwu9R
uxvn40++vJFHloOw5sht/HzF10ztWBpbzWW3lIDJWlFNFhnjCR4+HAB6TVaa
l1NTNmJytYFnOy05QwgmTrYzzpoYHpftqj01VAhtIhLlu/ia6ZZiiI8wLHMD
b/+cn1QNRj0TqTFhhjE/0RKAkGPRFTrJKdHmCe2t8KefKZBvM8UujS6kql27
KYe+zQuDe3sGqFJKk+wKu508B2WS0cKahmNBn9QUG5DNAFmepXQWHF8gdwzg
v3O4mhI+v1dURHjTuBZyqGwXlk7aDdvhQB/oT3PbVUFWYY2TqG+vnmK4OyjK
6szEVlXNZ0RBxvRCXCakGP54VVIjaqRyLgfHb5TV2CuJ0k5TFQSEaK/KZD7t
B93uiRqAs5x2l4ovF8cgxl6w6nAwmKlFJW7aYrZNIMBWrJ07bh6L4mwLExJe
Xcq97gVHgy418q2LBShK+tP770fY8wvDAzpPQ2XyceqLUTPlAdTMvuTb4WAf
Cwb+PsnCZ5w9mCmoTKwrnyeE7d5buVMt8vAKisjzdbpYI0KkLgdlsVPRRN3z
eAMFdoSHnb+zmluL/OPBkSTn4V1r3nNwpVN0wYnkpBSncqgiltKkUslSOD/3
uWmlFIr/DwPN6mWdASN/9WptnvHgVjXrY8zZeyAqfYv7WgeZ9+Njl6YWmGmv
9wKOJUMvMYdh6mJQkvwIL0Q4T4VnAlifBK8IboX4xsuHEHnJ8WDj+kZ09CIA
Gb4HGi5Y8xZpcsB4A+UzAez5FMbJq8R20Axo9WOEb0NQZByJs+knjbqda271
Sdu3vuu5NUh+Tl2anvoeNIxSubOW6mey9kjNHojhF8skmr/Lgnd+zL91AshO
duDvoEFW4hGCD/fRMe2XhDENkM3EPiOGUzBWqlmneLUpMg/UeKMX0n52j8Ws
+DknkAJPrcCz3BJFnosdoPgqpyATtx7YlW5qrH5LBcpZl+NBqdm0Bvn42ZPV
Ndywpt2QHO694NIx98r7e13W+PRf4QziDWw/3H5RlbEG131vH+EBHQLLIpwU
D55XFWXa+lj8ItI4eT9TijJcyXUJBkovrU3z4kwaBH9Wk6Td3L3jx/HX/6+D
c8MZGlguWg+phQUJ0zs5FnEVpIRrRAjMw5tlVcdK7fBJNqJVNixvCCyQ1qPS
ohU2ZtLRT730SrqmxKk/DfoIt+Szrlnu/zadgf9Haqg1BeKLF2XqzZv1gEIf
aar00R2cbB+Z2Cik4wzyZ+92meyE7I+iI94rCePwjG9PCSULRsirAnaQ2L6L
W0RAocRtSjQJlIUfgmhZe/ECbQWDBSSjyNBe4HdEaghoQPEZuxzOTFL0sLX3
RP0qhtOGWIL3Klxn23RGLCcl9qbVKd0z5Wa4KieZOXIFZpe6bph2QgOXNSy0
sTOQKTlk750GmguAc4A5kgCbDSFESedqRU5IOMnFcXmukLBWgPSuXnkrBg68
DpTLAHiAz5y2mxYPUxVGadM0VpM6P/fwoxEFllKUnkaWZVD+h0PvEKjGGWuL
c+xxo4PQ8hmcxj4RcWgEK3Wy9NxGF9dArEQhkbGilhQQPLSnIrOpiOPZxm+G
ndgm9jN4vL6Jdi+Fz9q6Yu1TeEFSmRzoQk29WoE/KdR2FKysykCXKvO5JKJ5
OvlvqjK4JHjn3mHM7d/sZ0ouXv4wfbuJTAgNbsriWmbArCOAfp+XAo8JnBEM
If7UreS1Vb1YzzmBNbSlvImasvpZ9l9Ig1hjMRqdLOZLGEFYCDxYYjbqkB7b
vdSSFTdQ5Ez1Z3pvzvbNTlCyMbmFVd/9IvpXXsUvEU8N3jz3DujzBefh8tyw
yNLLw2y3iKEQFuF+iL4v23297fVHFhZ60Ds4b2wY/qUUecl6585GHdmubxA8
v1Rb5ptBaPDSyfxgI0AcXEi+kbN1oie7XRbyLlFbYci5GkdBuhpA2e3yWmcB
Z0ER8pGU9EOA5K/o8mm4xJ2CDNj66BceBA8I70V5kCjv1ldRyQFOZfLx4x/r
ZqKc0t4o5DRX4Aa98ZpcHtPAi21eutZ2EGJWW1PPVEFzXTMxDv3Q3Akt5kBV
lv6Mf3JztmyaPTsaz5mVcSD7Bg0JW+ZtVdLubOd8SsGs1sStLg68a1jJTbn/
RVPxQruDE3dUaGUHktbAz562elvYBEcwFrz9QpAU0X1u0NmGZlIL42rutC9B
kc0NeTF/UueuyEjIgQI8HFRVcifeauIQOc8JrG8ifXuzmn6/dbZINynGxDgT
ZBHqQcdW2QU7XbKoOwNXz3CDSPjfA4drkpMgewb8GGSrfZZgE9HWwQzKoi4a
2dtYFaHREcG+L15EQCdLD1vgbokszce0J8sVpJ0K63tjJ59MP5P9XLItqvKY
9RKaPAoAPus9yS/z0ERwP/YHLcFykebUL8vlxio2DZKErA5QucD3H7F5Mh0u
foXQYnoYW0ca57FRzMhRi4vwDmXSykPKMDchaVJf7Z8OpljFOEcnqbYM0pFE
GoUaoljEpL8CZSFjajgSVsrYy0nKUPg3Dbp9w6MpOqxWAr7BTaWK0qKYkyjB
JmDm87CcIkt3Hf9kToYzh+oYvykxpx4oyRDnjcsWvWSXVflvYpILB+8VDOa1
xoHO3WF/2e/CYByqgRzNYJw7EyVZUsdBvc/bLlqvCZzGr0V3jc5evrBEWt4u
XiaSWYkBJTYywBiDVuwav3GQ9bAXbkjppqRzPe1sdWCmTpc+/K+J1KhJo09g
ea6LBkmGMfq4jRUGeuuqI30wfc8hO+hlXTEftlumqeO8ETqakuaxkAMsBgsI
khOhEtgJxa5dT9oygZcJblOpVKVHAcwvFdg125bBCD8R1w/EOzIs62sn++NH
Ru2Ay4Byu+R1PKcnBfP85GOBOydK1nI7w6vaK+OTKfl3hdgbKhBGlAGqMUrf
rsa4OIVg4clEl1gIKuympGcbAUDd4JHCgkbfz1Qy53IVREXuuWS1+zUcYeOR
KLwuxwt390iJ1kkiybd7FD9VkV5q+LxX+rOhUlgV0DMpiQEXyKCXpo2A3No8
TkG1YeW2tfXF+5UE+aMv2+WuGUYt2B8ip75L7imiyBoSxd6wBOnH5fipux4O
R5S2NqbNXPMp41dxhS7e7ksOpMBxhBQ30Fy+SzwQ6SC05b68ElJm685HANyD
AJRTq92DVR6yHs+JgH+l+nPuvLInZq0dwoM//kI9PaHjvyy6+rAiuxDi7lLF
1QVMYALwo7y4eFALJuPPaLqv9pZB2uznMCBnc3ORjVE6UAcW2AYXMhWr3POt
+HZgLEUZKSzqE2suMRouORw5Ow0AP6lsEsxeyqjFDpS0hQzVER/SzOOTjNz4
PG18HA0+8pPlWfpKZsYODrASNl32UYokQY/T0XcqJTCnUpuxwT8hMx/MiAzf
LRxZoriMf39alz3B6sfZWa3a+f3p0ar2PpOv/oFTtJSN8iKY8QMawp5YY3Vj
e4aneC5ru06w4gmZl4gkL05P73+ZafUoxBB6D1S8GRmf2QvzsH+3ZfmBaDz2
6JPP5qKcXpNNwfN9/kXr4kip6EYVTXviDOC7o6fVyGYNBvUHDBD3wxD3NnPW
fAJa92gFtrCm6cufUfXESJl3O7prqK/bO3g085oZqp+kXlJuExRM2PorMrt7
fPMipWlRiixwUnSMrsvn8FZvq2n2umFoIJOGxIXMACfDtPQ/TBMWikKdyRcX
8QOL0RHDRXhi/QAnKXFABI3N09sKjI7QV8zepV97R+zQtkWS4MGhc0YCLm+z
YeQMzsXLmjh9Y3RWv0VldTnSnduo6CpZGLdHQFhQzC5r6rmWF6wCRn4DeNSw
/OYaVLc7dqKqsjL2Yo14gQ/OnI1DTPe8fr8Zc0GmY5dZ1Zo3Eq2pQr2MyLak
kJ6SRomIx/EB2eyRqo+u3gnMaAJm6WM0A2QpfumO3rD2EfJYb0ASXVV6i2ZX
+L3CHP2fxUOlq65u6G+OSjhuCijCivRMNoui8+iuQMOiWI8e1rK3bNCMrzPw
svWwRUPSUY/pIDm/OT1enmMe6ZrIXKVEBtMNWutlYAGxUw2/SEImlJy/3xfS
BC74nmly04mqrtSuSNrV/XyvacGw5nOs0kuhGG6hcY/4TVtW7RaQRv4mwCUX
OsLQDZcgUL51xJDnsUQjPNWPA9yZcneb3bTTneQsUNfJcPI+2Y8xASTKFLKr
UdboKjJVKhyq7S1ERFfbb9/6LAxeKdobPtdl4+sbTJlabiChkfuoGPr+M/Mf
iWePw54O9FwZvlAweqNiBgdvnhtjItxcREu/BsZAXFBxaD5wpam03sPMm8Ye
raXk6bXqg+iZwSEIyEi/qWr1l+IFv7XE5BtQuSYF+rrKLQxyrqqhiuqv/Anq
UNgO2bNfyadSeFAaIku7vpWy7NdEDISBWCS880Nx3/ZmZCnT6rfx3o4V8oAp
VIY5zKv7uG6wkV5XRZ8ip+E5fV3/D6259NfrWQvLXXHuxqm93xBqodKWU/Ai
tJKGqllc+H18Ek1J9xvFcSugNcIjFqZPipjLseuCTSha9ZKQJzW6k0/Yyylo
QkB0s+01FXIm5ZwBoUtxjbrV540B2oAYuqi5urHnhmFnbgDU7ag2zgy2Gnoj
rRWo/sfifYNVctJ5uDGZGMAP7HVxc1efKXU2vN7YSR9fsj2QQqfo1gn9FWMF
k0O/29NwgWbqrCzdTqZzQsZOi84IXpJWjbBhdflzWaVA33taDwywQFbH1W4C
5I39A9GDG4oM1ixoH1i8TCEMZQO+8e8r//mooX7qJFjHUslmOZAFA++SPkpL
7Wf6qqvQtTdFxQm4acy15ks6yAGYy7Moglfvc41NEs9fzKf31qXSnGXTTYu+
kWtP6fd4loJVMpmPoHhbZfBdB1m2WYIjJaEQTG6a1A+7OJx/tmqFV1loOo4H
wcETEVJp+yE8s8kAwLMEynEz16BzI5m31OeK5oGgU6Obd20LdC7iDSflMlNe
Bjc+poIZoSedUglLKRHAPHtCefoSZjqlXXflg0B37H72v80bNhfCtogCaln9
d7Bm+UDhYJZ55Wt7Fq5fuq6SGJ4Qvz4fjSBoro8dNoQyWOouVmpR3rW2lEt+
qrK9i1CiJk/y7xBH8gujFa+efeTMFNTYyLT2jeulYHmoLdDUj8gdRzNl+hed
zba1xdGax7uzOVqCknA1wfaG6rsepDyDLPT0FkRLvPKbaDh94k8odmyVITkA
gf0WCnh7Dx6uZf8xRhrnMA925CjbhqBaq+RVROKVIbKqwiEl8IgfWcNT/LKm
FzE+UZaXEwbQNPzbm2VLRiEEy4kLl//4nQ5oKpByu5eqglrHBtMkO+MNBNIZ
pSSC07KD65TWYRuhMvYvI2fQUP7RK6yOnz8z5GgiTK3pLdthLy0Pw+jFUfW2
eMRO6VQF7JHmYsSWCFuvncXtVjcqP2igmZ8zfjYaFXJUl8SABXi5isoMx6Ih
L7eNorA82fs9oBYtnoBxNFdFvY/Ewy5iOH4z1DYJmtH19F2VDSK9KkrMZqaq
N15W6nOlVttkMDAsddu6hyg7Q31HYj9krFq93f1GmwwWAuAcPdcVUBHJKIR2
3LlTI1NcCLckJtUKDZ5CPDrQtTCPgiME6qU+eVejcHk3yrgHCDm4kwp2RG8F
Yvei1RQO01EMI4JJ3IK2Tw1BfEczttG6rYDc8sZE95ZQR6hK+dKI4xXR/+bE
7lhAzP6qAGRW9dZUMvSSeZFYdoIcZqkQK4GpzhH35ZeI63QG+45mCrYTl1Dy
s5/dJeN25j5dKiUWYXcLKc3Z9D3IvXhx4qootv4j2abdnKEZUHh+yqnpwt+A
HM/AJY/8GNy7bDC2cj+a6UYjNRqpq/2TgOQcbfkJUg/APLDwMXoc5PkgZxfO
6mPWEuXSZ2qYZx1TM0NJwxDjycdHLscboMqcUdlyexleq05vuU0wBE54yrop
Kfkft4ZBAF/tqKp6rVvGfJ1yYlsh4w6Tsydr7qLS5M7ybhHYOKZMCW4OXC61
Lz7YwUCljcT3kFzNCQPtsnAwO2SSRfk38UfH8i3HNsK/KG+GyyEZW6Cp+3BT
5I9WEJOJ0bVhoXG2vrKZ10Xw30fzzMyjwW7wV3QqaylDxMOGmODvbL4SuKpJ
uCjHQqQWumGTKxoNjkWbbEsoJcbz19mw9iEKzOElpJvrZ+uSX3hgCrI7Bmhi
y/72+Mj05QruY4BoGzRW1GpHtVfi0qsHrJtU6iIfb+8lZc5/zhS9H5oGPakR
fPR9gJQnkpO1lMsBrcdalT5DG5AasXYsQl+cdDAjTprEAQ2Pm3Wz1D41W5pn
mNwEoLyQ6GEkfI+uOsJQgie5my2ZHIDF3lcsx6skje70IE6PEO4sEBNXJEvu
x7Y3Y1tKL2aLqiirEtdQoyC3qs+2WwIO4WZFYyWFzAfM7Akhw6blKXt1N7tr
WXvGbw/lqpSAwclHAW0126lHTVW7PzAUSgWPTc5i4G3rMKB1UJo8BpwGyT0Y
exsb+NMVz9oJWg76nG+hfuWwUlEWq0wnkiVqnRXljc+/bNKbXGCgJjqxiX5I
5lguEmZAHZpbSmL9eq092dx1SOuqw4Rv68UMWlbIR3962X4fEwSFBK74bsCT
W+89T8jbj/ZamUtco9nblXbQoiRaflM6BJbgOMyll+m/2MjX9f98usjqr4Il
OZ1mgD2ls+0ypaQPuEevb7PEfsBUVPeHHm9wNDWPtnPamIwAkNarS/9ncCOw
98o/SrLVMlYJ/uTvr1M5x6FbuWfVwUQoo2x/JTLksGNfacLeClE61uafn/b0
iLYqH4Qf8ALIlhRqM6uKoRSlSIO+/TrjASCdhKinP0lPxi4uY9WLUqqduVtk
moO/GhfyStc7gvVq7WHfa+5XYrkGxZAX7wCuHuVmi2zxZ5IHVPH1ugs0KZKa
x7R9rsJiiizMASwOGM8pWvAtiAU5n4FU9ny/YE818wmsJ9CsPsr37EaZ5u98
CR7oj8Qak8n+jHCx/VOKoBOA3xHlTfdMg2sLqpzXl2b04G8sDxYhLg3lVr3H
xBA3Djt9XFly0H8r5xUJj9W1kbJ9s+PYPeb6ngdat6jVyQ+VjDtoa/yW252h
zP1Cm6mDcQuRBsIbHf6JDjIRaLeWpAAXdBEqysGlA5mc3dC3O5wjTvCQLQPr
EZJ5iBg5mADIjhFOnWNOCLKF3KyQXFEHRrLsd/dT09MNPqt8iOjubOQgAz8O
h2Vmxc4eiW/9Dtb7i2lecv8+1TAkiEFY8AXGyDfobJ+fGne1wPHq3GtlCWgj
bksU7H43ePE5WUNF1KNcpyR2aM+bonjPYQiHnZ3CMVCFtnZCexsTozZ9VPOW
qswuJzr1cn3V+K3w8Kevi11beqLai1F6aS8I5prf6K/g7e89iB48y6PcP2UP
hUTgGDZbRHLjv5zHQHqXyvn6JWQMkEAAz5eHHWflHo36ITEfznZrbwuNwH/4
AUzCsEo/ADdHkK8L2xqo3EfeyjAJ5Eau5empVIKKPBBUi3hQoJnFz/72I9ar
FV/3BMj1hvERTr7dFOsoAgybMZNtc8t3RM7Lo2JqDK+0j4n9Kqv8I+UApEEU
Xg9dzcIZxmpBZCZZWqmlwdALV8nE1qArOZHruc3g2zhH1xXHxPM2Iw7/UPtl
CTP8HeP5ZngymcIcCaBI+aTnBXBUyEXu/9Nl1f8uhsoQ3lJNWFawGsA1cUCD
kQF0PwnFFStGsYQtd1iz5GzKwnWiPoOtzTqGWPpqbstECHM0C8g0qNGrTK5P
416C5zKQLXJaSW2uCqDrVvWYAOKVyeNZEpcQtzCifl2YcSbJT7owIMwooCn0
ChZM1Jb6wy1ZBYp4U20hajxRdCPuIBAUrOV85x9oVU1ydDFs1zR6WLKbme95
wpEUY4RKNfdzSrZ7sdGPKrpPZ4eIPyZccZ7FW5gsDdH6duFl+M+tWHi9zXJ3
V6sXCCHRcD8XQH/7bfio2bOxhPO/wugdXRXWoVOkZJ1FJaPJrmP9SbXvkDwI
DjDkl0uvzyzv8bTLbABvP+1AHcZ98x5ep8PsjUDdGXhBo3NzC/PE0L/In+v9
PQVz82wlHM7yjd7ubtBPvgmu4LYH7pk8KTPPi755pGEvoFv6jDUk2lCI9rmY
5aOqgIi4+d+JkVpl0/KRFyb1bd6NvXfNLfPyVFcKsaHQtUzAGcwkkNUuVkjF
1FydKK9y1/HcL+xfcp3nlabnnnGDggn3WQVOJ7oMrRcLmd+g6HI3RFO/UcNV
yVk/a7f7bRowjU/XoS4QKKWwGT9cIOzBaGFYnzUn5C2wVTskCGO2fy5qZk3w
Xo8xF+jQVvfdKUSbco+Gn6s5WAz/j5s2mEVeAIyRAPPqtp62AIFvI+KILGb5
MsqAjQQp5nX2qq/0M/DfBYjq8LKtVbcuAucHzTdEIh5BKhF4JHEs7xy9APEB
+EOZ46Xyw53wSvyT3UQWC0mBBVTkvkItP6aRapa8IAGVB8Jxh2OrEJ2Ssb4g
B3UMeAZmbJG1lBRlXplMsr4EL1/mbXCTTC07ISKrJk89GmiFYIcueGQj1RKw
TStOTGmvHL6RYhQmZEPJ9zy7mJIZIcRiXZyrC8HU6VkikHG5d1E6/5WMpCLP
pAFEDGDY0ypBcnZjD1RBwh2drnEAQ+SSXEuzXbKa1EaiojuJlD4rxXDbLTKv
m/UqFXBX6gDykxO1ajiWbQFk7i5eY2lnQ95Js30ytS+pZ5oSn70ZfrUmWih8
PQc2XaGIIp7lEXU+3/P1A1fGQRs8QhrkcUtK55k8yPEk/rGrvwk7UbsOT3o6
ZotEhIxLnODkpSff945iXhjPavtjCzyW8GtUusN/0p5/e/oE/KdwcIYe7CtM
kZE/1cHhrDEXHRaDkLz12k4lWBd2kEVUzGWtOx7eZpy6TCEgfibzYdCACEq1
RaFucp9akyKINiFNWWdxpgPOcShy4NstzN9gixXJ4mj0JuJnHBrKXxnST234
uyWFbXbx85fR6SC9W8BlhVUpoU1JSSzCaqgdghmTVxxU09KbBtuTGqqUg2Ra
OgrDf33kYBAW0Bo7DTc+UkiTnPEIecotPebZipY/xwMpo3oZ6vDnNGd09oAn
SZNmoWTfZkUVa7Vr5ZCgYW83pwpfPH6/53CkiYjPdgqORFMfC3n2z8+MSCGf
gs25BJ1XIstb3jlIrj9BxkOcPVfPcrSpqqY0Eo70bsv3mCVziiErAiSUOOqX
E4+ZBxdJIHKNM3GM+Pel6/SR6WnWT8Wx0qUSSjunFQNwuCBNbMnE8j4evWBu
95KS+wp27ToZbSofkQE7x36MVbHZusxPIiaoWErSCWTXaNI+/Vr2s2UAOQ+I
CGYvx5SgmC/NuSkUNCeXd8wzYWU+JOdNNWthB5G6iZiZOgzWM2QrHlHa1FMo
1ApBp1t7RH94cpapFVrlS+tkwcnJq6jdh24vUlKsinPJpjGHIBdKhi6rpobZ
pSbR5t9js9t0McEGB7+Mz8Kfc6TqHuHpqEp+b8a5/C0LIy6X0m5EdyOPSUmk
ixBSOltrsKnrIQeRuBX5SgFiwo/5i/vf95wiWWtdcv8W1o6TAJQ+tYXQ/BMz
IJ4KAffLk5RpTnTNk5fc3jsC/ucgCzHg6dPS85QKRU4kbi5XpJlyvUprUtBU
xQFxKt3//ar2/uKZjqyHXlJkufaevCtEZ6BumE9XXKInhh1e7VyUezzR88Me
7uefIEDuTo6TPM+lgY5/cb1Bt0eUay4TUtNIdW+hhhgc+DGNHofOY3Nks+7o
lgWkX28eTYetZNjHdW6xIXvkkkkM78S33UCnp5rU1DORm4uelPRa/c3cICM7
k/GH52qjCwIWSnwkjShe3lJo/1Ok7IsbSjAeoLofsk4k6uhDd52ygwio4bXT
2qm3ksIF+JNNZ9AR9TF/SUe6aixQqgbQKBxxwsXV9/biEqQIDld93oeoAMbX
35PJv1Rf3fSjt+fjKHmR/c8DbWD0wXDOOGzIJVKt+a/fsJlHSymJgMy6ze8/
TwWahWl5NbEmJrmD10SC6zo8RbyS9Ru12Mcmevl6kKAkzY8cUEZkDsQ0QsWi
kBR+UpvTQ6ERqqlLcJeVjzIMvv0NEwTWEKTuWoGksCFeEuVPWP4ROjb2khWS
lTqPPqBRzINfPnV+o5IpfktXPhKZTM3JPdo3iqUawONdXFvFYd7RXZjU4i/x
eKcpIQ3g+pczaZ9YZzu8hVgwd2E6BRwZl6LSqMRHMWhFvoAhaT5TEK9uoqLz
CNTd4Lvn8abBi1I8Zj1UUgmgH+9XQ6EzNSQUvc9JpTkYQoS3ltdx80jJZ2lP
kvHvfqWTHkIniCJcNQG8Ceo7qUspWVE3TAJMUAr/Op165y3CDqQO5EL2XS6m
7okPIaVLcoSkvwa8qPe4tjsDeGRP/kxxxpJtuH1FYcd0jbfKl0sGR491Xxn3
fSBnQeHmv+qYpknoyefgSNlCPW1/bZXGi+Pph2bVHK+TLY2NtzQs+YmHuRtm
2+ZYn7ihQ9TxqssJp0OKmdhTG0cBDINmJdZUyaouyI0neUfQRxWWEFYJf/q4
xFRVaXBGW1Km0W9c48MNmUeWYNMjTHeBB5mTvaUC1UrbiRHnTIFhDiX22Rre
gGB6XXFhOaDPGfQg8hQ39W7PIyBXiAJI2GDJ4csoyBlAAtM0kHBOEWDe1KpI
oB6YzQ8Z8kFKDnOWztiNAzy1tVZN0oKQfe2RtG4uMIZZrWDC7t7b8XB+QbHY
FdLsbULH8gS3qu4Bf4Gi6T1RyfMg/w8bturkodQz9qDsWqpXk3sz/nJ3F2Zn
Mfe8GDIv10pgIMpLL3LnBb6GQZZOSTDAv2sdS0Q0jBmnZI1Ybn/eMoAaloVt
UF/xT/xyNOdmiSv45mg9Sv1xl21mP0IjCb228CjUg8gETdnTm2LH5v8Lpr6F
NRwG/K3/BRq5rQ+BBApZnc8CTn/onysOpm6Y27GJoir83imaCThAre2X8Aoo
3dN6qOl9lqmbvcXdZPC/YKMTYjKK83v5bD9Ib2cLDy70XjxJrI4giEOz1CN7
ohcalX0cNKt7reqpTSAp9T4nYmbU7xadsKH+XBP5rVrrODqjFLI6KhQMxZU7
FsFk3vKTev/hySnexXIuZ9MkW96v6UINLVP1oZaBhRjrnxIolNsVfUArIvYv
cIQhxc1ujmwHNYGQNLGcUSDI41Se1n8OJ/luV0JOwwyWxdqCkivKqSOXHXJY
/JbRdP0QdyG3gwU0LC6MHlVnEChAGwm1Of0j8aj6h/mWTnhR5pitPY2mtn5f
ustRD/RLJTXRdWHHZN/HxbWyjFpV4kv/K2e8mAfB3oD1KmzCEPL1VNgYrDOJ
RpVu3fKLESGiT+S69QVNq1c4MsCqd+xbZJm8xdt9T6eQ+IgmLgJS0L2Yeor9
V1B42ND27m4iZTLot2GFdVHPD3u90TirCbS0JSJTztWkLmhm8K+CnRXFaPij
BoGWqqim0T6dduOaAzqtcMiJRXRlq8zZA2O9BGDjU1T++jC5JBDtuR1NEm6L
WI4FXthXz+YGaxWwTrBDIIpqmJ7+zkRqfng9E7sm2gCerHRj0U9D2Q1A8vr4
9YAslmLBgEDuUuVrX7WynDXfIwyrPIufmhzKBKd+tipAKr6jVCvkWn1WchLZ
xpwRNq5t9TdSvpNfnLEDpH68dU6Dv86oNstbHlZBcAxXKj5+rtDudrQ3G8iV
EHO5YB+1y5BRn7P0w967Kfw7IugOeyk6j+lHxHnm/YbZETadtiZCcmkpDZ2m
WhPeUP8WRa8FLHQ+gYhWp0DSI3ottrSdVtrF6+79qyvAj5LcDKu9OXoR8jRa
Gth7DR1sPk5gXs/+X5pDeXFHJOF6ZYERa8//Xqj91nlDDqyHpmB/V0YJKf8x
M2nJmZ6+FADX5yT5sA5C7+cJkvbK35vYbkwfjXn99m722UBcdil084UNL/UJ
JXxHRFCEA5X0PR9FCnSYvslUkVA7YFDQk4G9x/xJxUbAquajhUstqW8OwMh6
cEdlMLTsOcexbgGXd9Ia1qBI6aKOmMdfCJc2s4ZqWYkCdNZkGnyX2/pP4Zcq
9SjCXgqHmgwcQvNBfuM7BO6xeKT3q7Zo8T8wtEkypzsQINEk5T+8r+w/ikZX
4klw/YX3FYaKY5TCrNNMw/27IVU3SN4GOk7lmXwl6LMao9tIpLWJ21MiavwF
W7kC5PqY1rHfhgI5cbNG+sGwoFG0e4emIK8vSn8piwhwLl8P2vxLYzvqFYa9
Fmq1S19f67iK3+S24qFPn9+Egtm/BCOiZtwMjUS29jtBiyjKy3gNqj0zC++B
eWfCfWuprla4nS0kZUd8DgRl/vicJLWwY9luAJEYrJwWRJNMlPthxCp+JE0V
sQ/vnll7VaYf0NrOBBwFCmMmR4Ng3/IWzckDbH+X7SC76Aq/xNjwaLXCVXlC
RL0JPWzjzTuIf3s1IXpkavsad60yf34gD8Q/yEVUwAukOfJNlOiwWgK0iQSI
oZ8Grom6s/Qfy/0SOV+osrCnHGLgDu5C1Jkt9PQxs/aB/bCyDCydUeQnO5vl
6SvulMNZgDgdcSZ80yes4qEEvwPBtKdcjFp3GT2ETUbmwnvaxmR0OWlz0fzP
H+FBxOYZpJh/6kk7/NrU3st+iyezP7IHOqGTIP5E3bKLb+STyW2bK94wOmgE
FOouQZMsAOreGw075lv2eYnX2IWJi2OOtkQth1g4stwv/bBR2lQGg0ykC2qT
B2jWZrgHTChZaVKJZJSh9POFNBVD7kaSmsorttli/DhlvEEriZdTIjQ0Q57y
Qj2YjkRr4sVIvA1AAwy9/5eh6q+yas9IIEDK7En4Z2As8hMwrWSJN/+xd5KN
cbk/140FRxl/Mv9dX//6ysEet6dKMILC8oMMeHplgL/Z3V9tY507d6Fuygc3
f9fNGxDTBn7GYEdCrUu0FxJRxsoUxcIYfJp1J0+2MlrYPsrJ7KZjlZJd3HOF
UeLn0Fluo5dfb8pHklDtJ635sckbDR7cb9Ityv4zKjbOQmRQ5s24HOhWJrQ8
C68ZOVXaWWf90uTCHNyccT9DI8mNoT8t/vXn0KndCX/2F0ETsbagc1g2b7rP
hToubXs2mcgbwENTJcu/8c40MiXQQfWv9b+LiojADSmk6CS77o1d4cvn14if
gvNWihQ0XXqCd/UkmY9zwRT4Ac5HG1cjwXqjMKkF6CFAGjIM41ZeZkIQjVE9
voxDN17DEkzssUP7pUi1xxQk3TtB+hZnMV2XiVM7wZGsnW9lYOUb+3g+gd7r
bzSFBxVfVp75wqKwpUJXeZUPtBNGGwSdvfCsh7gsZ6XyprYrbXlvLNtRdiSu
jdPpU7pY1GhaFME22FVx1vBe3SFWmm+sF9fewDu25NnSDsqFCJAzOvlcQUpk
fKQxS5Jx0cBT8/fVY2y5S40BgKNjjckuFlzXCOSoKTKdGC2sBYlFHm9hAn3q
zuNC5J8BmhFj7RO2EvRLsV5W0kN1U9uI0RblcxrlNitNeRrQV9JXErjxkxQu
48H26ZsBfI9Z5yhk0Ve7Fg2oj37s0Xiqg00VwyWbMIDUDEw/jb6P5Bma+wJq
AKUoyPU+HwvJMjibNbmgtPp33R6mgpUcldNLdb5IGwzJZOJGLJcASvY5Oqm1
gi245UTarhfNVCto3eyYdXYs2afsCvbCaFewcC2A8Fat/SBk5eXNZOATu4WZ
RmBILDylKxGd6UU/TS7wOxtdQwpf1fnHFa9wWNhzzXEzN6kfiTVtumbnT+iN
aFuypchl0x3wJt0sMp9uXJchefYiAz+vNExjskaiLyfrpeVBsOZjO1mk3ua7
k9QJ9G27XqY6evtbxrKoJAYSn/Fx7SDp8TsC/ggn4C8EKgEnKwXSLdb2eLfD
mv7WKLN9MpHaH0/SqzqOK1FAldll3BxmF+niEh/e0vOARIe4EcYv/LkFD5CF
lSoTU5sOmJ1H1xvvR5hF5wmkXnXkeBNXdIlFLTsUv7FDm0Njsg099eRrUC6B
kUo7bZQRAXkMXznR8oVp8Z89bsDNsOkR1TjvGj/cbRbYd/kDgEj6Wz5vkZpG
T4KuUdX1Vx7JyaSxQW9XoxZQsg4gtub4VD4lKklg/ukj58UJn8+IZvTLS78Y
ONpxIYDjyOHPHcc6qa57wKsiNF0jvecFzHtnEJ5E/71CIzZr7Mj+3aF2shsb
CN8nZABlpBOzrpOJoIYRptIO3106KmgT2eqyGQwAhwVyU83sEzshINiGGsfx
tO3iF6Egpw/N1mbwbNBbBNdPJCshFiuvFeKnHUxFb/k9rOsJV9HBJHRaRh0v
ilGoBkODXpYkTkezPyNCCwDdSjHQ7PwBQ8S3eBLBGCufunsqL/3vrozwT5qJ
7ymA8WS5otPtqSp1oV45fMpa9g2/S+DX4HG0GvfdJZzqWHMcJiPpH74nNyEl
nKqgkHp997AojbZL8urGb/fcLAscD1DPNuvMuzCwymLjrpWOOfSjXv+/vwbw
Xvm2L6PrdkYy9QgH++eXJi7L5D1LtgQH95cZIcEnkkcKxr2kWq2o24Ktw3Hd
siaxV0pfqh/ZzbKsI/SSnkevlAV34y4nrr/4e5xAKzcd5YnGUEmTMYgq93pw
f0L/b+Myj3a86pll8VIDSgTIh/DbWoVtGQTpTFn/NI2BYOesyzL6fBuByAsa
I21HiSjYn1zJiOw2q0EQxRkZLCs/47xKccnhYk0ZE5oOBCZf3eDcl2bj+9YC
tdp8CMmEtRKWJKK5NZAmhe04g7vu3E4Qp8tG2v/PHKnbc5zRqX5qtJ78I8l0
t7E4dWZueo290xoVDK87RGnsSnn6qAuw2MhM/BxWHzI8lQrcc6B7i8z1Q77M
mzoAT+PtMfiLi9oAsfPX3EGFdjMxwWG5tAJvLC2efVO+NB8GsbU7WcWinB79
VweIUWZB7QcROyHUCmIfsDSQ8Nfspa0nf8fXEzwuJuTLi/Ts6HH34DaJn7Ts
mAWxtSmvlIl9u/4htBUlA8zWnnzlkUJmie7wY50VFHLi4isrLzrO8ewGSYiy
Uje2syEuWhBIIMkDTMTF/hP0iVd3VyDqeg/Xodnkhf2Uj7gB+hzSC7uAPkOj
+uf2i3tijrEj8+2Ybt//A18dwM/2XgisIjNbxvtpNOoHbostxN6OPQbf/5Mf
MPYEUjoQ9/KlMC/7TxBUTlI+0lOq7MZVb1LrL1lXAiDYV659LaMXY6H4nhLJ
/oIpQWOqEEK+D0aNTYA7IWOypqMSxKQh//BU81JawKRs593ULsxonvRIAVOg
wAv1X84qi2jWmLXulmp/fdIO3bGWiatzwUHJlj5OML6Beo3DEVvcE+3g9l6e
bKWTF4+P7Yna0lWRcnrmuN5yMbYXQXVF5/EH8kT+QfDeyb41DvEam9+DOHR3
8E8JvSXtZkvdQRdhBhepOUiqCpo69MG59MDXooNtNXWgB9fQd6FciZyE7BMa
9G9FYEdqutPCSRguwJTVT3l2EZKX7I7cVc7Uu0mRTvgPY/i1Xcek/oBC8reN
kpteRhyvtDdG/uYkKiBnWkDxtZO9BAZRzu/6CIDk0GFBuVbUbtekSIVOgGAP
5znUaX4f+akagmffWsTd4wG5yHLm5tcATeOODWAQ5rgsiiZQ7ioQtxsnbJqD
+U5UyBZpuanQac4fdGE0UmMHcXNejDoMbRlS5ki8blONSbFDwUYsxInv5mZf
4szJcn7B03nBnG0ywlgsz/6KEwElWPH0LJXs6nTMbUYPq0nMrYAJAsKRKnCs
cOk006JnVFrWiR8J815RWdt9kaIlJ4xo5fgeMUy55bV16RUPuyHdl61IADPQ
628KDUbS5QwYapVAJ8SNmo4/xWzybMIPO5tFpoIrkEocfHgKYNYEMCve67Vw
AxvZJnA01n4jir7bUB1nXzvcKadXigubxfNxr4nojuAXqQ1XSn2IQ8Qk8wY8
WAxGcTCSx+tzDhpFRF3YFU+2zNdxZ5/X8ubN7F4I8RdFv/RT2/IxQQvGc4Rp
z4B88T+ESgnpg0+XjqM/1IZoeXlIrvNlDwdS3l0KlOd0ScARBci0MfcIOxp/
+gClR3f3szirmFYB6qUkYc+266qpfkaDRmquPZN2ju+a6nMYaXu+2dKm6ort
fPO/3FRApMlBiJXNVE2wP8BWOZkumpAP9rvqp7twieJExznGV5d+sUyzi8FZ
Jog/m3DE6adN2odtGufH9KEYpH7AltPm0LkrCw89ewjDWWPLMgldaSbcPo5v
F79agzvOWPozG5iEcNH1ynjn33wcCON/g3p2a0cxqvD5WoAUjq7VTUn6+oHP
1f7Bb+ktzQNAVmZXcUQZvyN6/SPxKACaH0Bm4v2TNyIm1EFhGFy32EwQO4SJ
rmLfYpsXEhg9LR1EE2IpT5/oO1KqYt22O+fW2UAAsdnHdtZA2B8I9Qr6oUbV
nB3+58B5I/OJVMfLDKjiN5ulcvrguFOyISN9tIq5S0HNTC8kPLPFpbqUxWXA
lt8JBIK27bScdHQNOPWnHz00XA5olghhmhp52cXBkTgtFcNba3udLsRMZtNe
TkhuEjtygJDVsBNiyrj73OzQ2tqF9J45LxgEdeL0VqZbTcc5PU7BldVig0rJ
LKJatimsd3pmk7saryX6H1EU1iaok05Ef2foUXRJHxIBTj0LD4rNm2keOVoT
qC3yzWLuyn3uDRcf8d8V17125GpKAui9TDnN/TVAEiD9lvLP6IchONUFIkMq
4L+VQvJRlB8X1RfcxOXiZNXy3EUUPu70jYVvpuA6j7w5QJ59sxdkY/8SCOC7
fUr/Ct6Gbdl5Buh5mF8LuKC6+9Jr6yYd2m0TZmNHr/1bnEVbpvATdIz18TBy
KT192kKK8HCy7As1FgrqyakjNLIzP6QB7ApYnW9b4bRtiRWcAArBz3CqoSnv
AsfpxiWjmoV/Zi+FRzbrdgQM2kXCk9sb5kz9BV7r8vwjvrKiAx6Aw9FWawsn
PJm6GBoFCKzOsLK+0oimuvJRZANVDtrLj80WfgMoP0HxGEpk2u9imL8qM934
WBJOSirdE5k6i+x+rOFPMS+slVS069k+YM6MHeMz8Bqzyb/EX2yzQ5uUOSuo
TKmdXPkBD8DoTgiceqJplr4OWmNlH4ED8ifst5Hu8zwwsxI0r3Db4T2Uj3I8
7+xaVOAcXYOvcBGRbsTBJwxikd+QLsqFNrdVDLEl6RZY4kolkvmazR6vXvGE
KNCrLTT5HDcKIF8ntPab+IzarcVpkpRjKK6fupRGR9TK47vjQ66obi2m6K8Q
Jdo4L6DnG3RjcIsGzyI2Om81fA2IhkHGbTFeZ3drCWm+8Q3mjRYnAQQw2uDF
o8HCqV343MAJOCWv1mu7PJPv8JXpQiRqzUL5at1IgYKAVHalrHuq1jVC0xeM
kUB33f5iuTFGss6jftsxP31QLFK4o178l2lnF6R1PZE1Ib+QGPa/q513Tqzt
SxDvBSAjvLKLt30f7rF8hEepgIptoxcMmRlzPLrr6MTAW+BDmchWPiia+YXd
WwY7ZxCo7epUexEPMMX/zzwd/gwofJiIb+oPFWBIKvJagzwOenvoM+jRjKqM
q6BJoDkZzwEJKV1wEfbISYvwr/ChtwZsMsHMf6MkreI0HpvDMMmeTpJIeiIY
AVM54Qtmgyl7sbemgzHLy41maJLTn2gD/JbNqSRQfpJFS5qmWFVcz62dcL8D
z3S+rFS91QBw4VHQlChPQ5+IiRvlckUQeuZes+MgvjI+EMPHNljRCb4gvJBI
e0y0kLwciqKCB5d3oOSylVNREmFg0A+iZJ+1bqAFKZHwgmEtJrlmnUPcPGp6
8+1MVEf9eiPBULRhY1Oovt4GKQ9om7xo84e2GLdMdfcjZYoIZI+YmtidVCS2
Nb0HZIxuLa4RB+MgmSGbP8KodXaDQKZifQgww7BH15S1buHPAkdsWKt8A72N
hvpI37FR9uJa83pg2YiLgWaQzLjMe8BYbo+zjOQJEFccYNlda+p0YWnI3/UA
zFZQNjLHb7m5H4kCbcUtWqsuq3uDdNVYcoRLSY1v2UpHsMgdlzQU/E/L5kJu
9Gh8nNdObxDsWnH2nrHdcanifHRONdNoAy+7PYv90CGBn75q0L/aBGyaZGkM
NZTbY8HoMq0H0FR0JIZymOLSXqOmOznyX8Ce++1ubhY06Pjkue5AzDWILGQe
GCm/iw73k7xiWsOlVXZe9Olc2bMnNRchUQHpWi1Te2XyFIPwUjHZlKBHuNBb
se/MahhuEZqi46XzUigO9TuB5GENRTeT3nkvfGyhWQ+heka5st4COQifr0U7
vuUQd1Quq+xMfclcjUuTOfATnwTWy41xgnC6SSY2iOBrfYwCrSAj8vxHZvVf
tm+KC1ZTSnn+2a7s2Kmq+fpGngjabOidhvJjv2MoPcfr4auk3QnzRr+rK0hn
qR9Al5Xo4Ela7DAe0wG66pLYL4spTC0hpWeUFQlPAjkRkVzdlYAWOWBisnmk
8brrqnFZ/y9ph++g8XJVJy2E9gihUKXy+DtfvdpyvDiccPBmlHq2GscHrPGI
WTo6eElXQRLkRCjTsnVEV+zNvSSvSsOVEzczqR3V3x9IDU71uqtf7A79IH5V
SWw+yoY0UJUqlOMpaUEeIw8fmMePHoT0CPeKTW+vpPUvuUtsxonurk7hrp1L
+GMezffIfGm6TD7p6PKzkZiTyYgxWR+XzYfjlbSlqnpcLQg13wDLMtV2beuQ
ZL0umnuhJetHbtiPyQeYOG4cgsGL/JTXTfHqa9tyMjDJ4EmHJnBXH3umt64R
g7VbHWA0nwudHH+ocYO6DYn6jp2GaOf3QNDCQAL84vpjRBPNYoanP4gWRGek
k/sg9wzwNTIa9N+VDsvXhclj6bbga23GQIWhH0wQRa92u39Mm0Br1LXeUxa+
Jq1wkHwoTsoIZ5pVlvFUa5Mj/EbMbOaiyL6a/1IseWdugP3GAsqHRzzGRcFu
geZjZYAptNqFRHcHrLXiPHErOOSuNV24GEifIhYkNevWpP/I1bU9zsoYomTr
58dxeyI40aDdfg0GphqCkXaGjtan9DDSUr7DsKPEEqOgHKODtS+WXeOvtzOa
deq2bJauoRoDCVRMy0uFHudnZ0lRGRfWosBqwAg/up3wkJW2HJHPmt7+sGn8
T/36Q6K6nMUXLf/pbQvVPALxZLt2xYCx5tV16YUutv7s6YqaHP/tmeFtuXB8
jd3ltfzv5UBtdtG+Ydk847W3x8nNoY2YmklJv1OgPmOiReBMJ3e2Q+DZT/C3
ddxrQShPXlk2Ch0UiIB3k/2eviRCOvW08Ec6qeioHCGDCMpNcAobpN/6zVJs
DxrZQJmJKZEuuGqxapz4NjGdgG+0z/4ZxQ4iS4TLeRYhAWJqDmR8DJ6WX7Mf
kvCv735N+EihWib4MyH9oxp5vTHPrz2d3ryTAhj2Dz5irMKL4QfKtuS59hnZ
jqyJuXJqxqbXd2Z3fXVLPRRgATHy2HHZDoUNva3UWQTscWdxO1vXbLgp4+DN
K9T4u22EqPJ1j+Xg9+uxaHuUaJci5Xx8PYZ/2J9T7Wz1y+9EX9Df5lsWXRaO
UUZacz2wN653OuzxlrnS/mE4QZJ7pU/ErlNguLhT5LdSq3atw8sa6HNlNlF4
4VzRn6MnuLQOzt6Sz/6DAgSxL/DKycUsJOq0KWoxnC/oG1tOLkB2Vv+gWbtA
1oFyaRO9vtZSE1/ZJXLDvSm572q0wQ1GafTIB39nx06tdv+bmAf5uxCie5H7
beItLADP7XUVkM1KchsHPEPMjOno3LsbaJJ6kAczF244stq93l6UTmUfkpCx
Dtyb8jenfTOu4EJkGuzAoIC75qguynI/xnL2yMe2FY3YnRHeKM+3ZPSqnhn2
nhfblUFtNXgO8LlxabIUYILTq/X3zbFvpjAUOqo3ssNUcF3HF5hySuv4QBY0
hWgRS1rwoTzNypyd7VesXHTw+FRVHRL6TP/kagnpAbasslG46lm5KNs3hc6v
SUaUbnniwfh/y1ZYbTuJQgqypP2WwvJypgIQH+Yjek5GFYwyzF9vf7t4CdYE
Yej8+I0XqKXQhy0JfB7vSr3QVHT/Dcr3Novm6rTV6faXpsebFy2PiDxgn8Ci
EJK5Qc8CnBB6CfmrQhsdMEhill8mq5zemOInDaxRaO1e/nCpnECGOi76r+6O
ukCELGpChvj8AwHLJTCZs+udxxO26ccpHqaWm4CZ7pRk/hLOUtAdzzWRnJM9
0f3Pt6aIP2dYW/KHxOaRfj18b5TpoBGfLd8FTUbiWboxmcdacRkwU1/CTuOi
O6j1HdIpBbxuHBuuD3UJ0q993qwdxo5RRQ5lgbBJt+56+FyfqKTM9YAPky4m
wXIFzpioM96pg0ZEChYlJujuAs8HTjgYVuYW4czFsBliTo9LrKIhEWQpFEv+
UM36j5cIRzYbTwAwJWqYYrvAhshlKUWIqQqtRafI598IOx9YRZTx51JO0ZZY
zuujVpuYTspg/zAVoCkb3kMm5/5FiA/cjYhWu6eJPYqAsvjQ2k4+rd6kuwPL
4wUiF3x677tOJgRFSBP4l6tIVP+4XDYOxosPOrQislYIWUtDbnL6B8xEDIuE
nb+gjkLXw2kIox845m36A5HDz8NcoW18l0BXKzinE1+O5ron3dRtp9e1dGWI
YwTIyN8ONUCwMgrSCHKbcUuXENM0gmsZcBGR2R/9zprHiZ87vyIvxo1FXSpt
pA/NDRIlTgCnGUo37j0vasSWYLHfqwIGuNVZWwCBCAOnX5SYw1SV7FfgGJwc
M1ZHXCHwR08bY6te4/cSpjYQsE41KM83IcORxCR2ypbZcmtZqYi3gE6V6GfH
f1W3TGOklaHsEjqE4FmhOwiswkrdNKrkqsi9NICFxidTdzS/mZi+99h8MZms
T4A8IrxAW+/0rTWiAI+SeMWpJPf3cA+p7ltx9+io6w15rvdgCtugHMVa8BxH
E7+E2BOCg4JUgHraSn79Hbz/NsMcCAkUhLaWS7ol3nghbidq6zxRN1Pdxpjr
ZKow4CyOlaZgwIH8ImeRo5g7Pgtt0LtdHYcIKGaOHEznBBVLfkVj2cDLToBo
C0OVHZYl3cxpmsk1yh6tP+SE8eDRFiJ9lMeKMejYjHczCEBAeUE19RtqUm7v
ZoU+Q1Tio/JcDqXaKGQVahzpYTXxI8+AfhHNmiVgCjDMnWMMjKcPq+EfbN0Z
IHzwRp6WUseKDer0XtLRT2AhPOLiUuw9Zksfy08LjFbOl/ZXMC4CUbNvstKL
dx5cSKk4cOxdxh1UPn4Du2t2UORDJjuwfIJy41Cx5aUPuI6aiyjX1y5/qpV8
+unM79iS/il9OiXe3tfQMGT39Tpb8+3kEeexK3rNlLE6RTY2b+fDqRlL8L3E
23nZHILlrcU1A5jp3fth76GrjXXM+T10DX0LFDcT+dpx8FIWn4r6ehs/f7Xy
qrT/uA/kFN5fzUjDv2gooMJdftj3CfaRYiyM6+L+nZY3LHoR3i86F5oGp1tq
eSttGXq4NBdsjbue2FVChhXKb8XvnK15LG4i3KdCIKDULA2B8UkexqUSesya
dH4kJlWm5s5QGJiNe9VTI5HAIpL59hKBJCI7dInFKyaos/gm8+gmubnfdHLI
PE8Q/Ve0YVJICS9mhSMDpmVLRvgwDfMe6pT2GhR9jrRUQS0yaEQg2xUmPqHR
TdPh8w+sVbC0tZlc6RpmSMEOQS5OXqOTPR2XlrdiP3zc/cS0V/0YC3aWSNGz
N33KODbSgEZSSLYHXVM1tIzjGGOgAy5s5ZOUvP3s0lXLMkv7F3CRUNld6C7U
/jbbV+7ckb/svCWBAwxJ7ZYdTIXcbsb/ZXUCD9vkrIuGqHjByN+G54PGJzo8
lmOhsMEdmAs9yHuPJccwKr8YqiPAldZT4LSgKu7+3mqsanceipWbW6xDXTeM
iBTSmrCfajBn8JeGR7C/5a93vQgaatpTYxfiuqwEvDWPoTiSgWhVggWP7ZGW
U5AOPM6Xe1++cn0ZtbnNvh/TrpH9mDUTB2yz4q3nU0NWRxKoCZy+bobkFM3r
Fx1ajxJrlhjA0ebhvWhleSi4FfecKAH3WVAhCMyv3sg9gBn8fRSboML2y2rj
aWKw76PH7GPGlFraiQDAp5l8k/+SmX6KFs+6a79hPqk1AcULvXOgDZvDVIf7
08EMTU/RBRVawe9BhCteys4QSRDX5KJipRCorrW/mQAi13bE2/Ky1F1k2kTv
GxKxmltLHMt/JLwmAKGQyJL+w1qH1Zb+VR3XrQ029aKQMtQ4jLc5Ci/37kTG
O5Gi/RBJwk5p85pjt6naKPKLtX8sVH0qTLIpNNMtgCdfVzujmvEvL+X6vAQ/
Ri4uuQaKq8l94k6v/n96KaqwyYWQTgBsJybfBOByLYDo5G4O4eT5uepNBA6K
fp5mPXcdb6D5cHWyDewTE3w6I2UljA7itm9lFqTNH+1tg8erNbv2SSNd2Ier
xNiTzn6WCs5ttHBYvK4ZXbN8dumqYaiwkydhkApHNWtkrYKD08y3kfGGojcJ
ydKpouiW0RiSnpnXYt029xRkDloILjXfR4cOv/886gXOpCcksilMX8BRcjSS
MiYedDkz8gHzftSDUgeu4R7uZolYqcSH2TWj2diJqI8Cz8PhRyQvmcncbY7a
oJMxRf8yT4ciA+hFyhnmT1OaxbW+2q+lg3T/4LV83W6dH8Ywu69o0krT5CD/
OuAIseJCgmKTHnxDeFPGDXr9ZbhrIi04qTX0akj/4w9sbYrPHuWFwg4VLAC0
pvwREQtwgC2RZ4WlO3KKrgG0MRiH6lj+1hJZslnjNb6cXdsDDwa/poC9tRjS
3q/lify80JNdwBUKrG9tho3Yy7g1ODADn3pZUV4xqo5ZAsftJiTVNjideMPH
V4BtT9KBqe4pgiQ3kYNmTK7Kifk89BR20R1pea12T8TBZ+4vRFMzAiANpx17
pVP0ozag9H35NhrPj/z+8RW0JOlKEjQTubC/DxDGzKb5L5fzSMSI0ZbDeOcd
QakjgjEWgt5RqR9PdmXz2kO6dCT6PayB7HTaiJjLIp6FgbbDagKnQGRuqH54
IDXM3pf512TLCQP+0QA3CPcjPitjkQiRbbAXunsC7/z4HM37MbosTsicNYGM
xyfOVJ/TkwIopZLB80o19dL1K8OhtiFF/WzNLN3BH3wMDZSDBM0pq0luYT9t
G4E2FvHvQd34mTtPzlkfEihaVhfrAWC1+y4KCedqkV872HOG+FdC3WP2xjDn
Azoxx5ZMl3eoWW22ljQG2hbcJhsfcijVi2XvgSiQ8ZcbUCu+stqgw+2FA2xo
uv712i73QN/tFCctIs9HiK+ubU0O84/mMETd7QkWjdJYW/J7RNnS6kaD8MQB
dDeA9PhGNAimukkeSYH7lZv0SIZ8AADavvUDaDwgwpNXw/IPefhfCLqQ2CjG
e6W31jR34dYLHOPDJIkDiFoLcTkO3H/YF4l79WM+JUaMP+0SlfXKvLoR1Vva
32n7C1BEAQ3+DUTPYvi9oWuY5pCNB9i8+oczI/mAdVVkm0OWtDl1iS2QWC9j
r49KfpU4KagG3iX2NrkKJl0YU5LiXgoLx+3EJiKr26Vbsx3T533qvJn5TsM1
FcSfycZf2N3nq/Wrd4mcvpDhGmpn0QcL/dPqd6ngXsdUtO0KV7U2hzTebCZg
oMiG9rUqoey7eHyITDY1VgaPBEYIsiAJMT4ldcC+ANkcoifWlx9EQJQp2h8R
kf9LyPZbkv10QRPtO4xqSnR9kBFJp6htmmN/ybwB1cVV3mvTHJFpxHCkFLrX
gb97k4f1K2KX9ZDmofwS9OhAwfy1QInk0+E9cw3WcNx9cvI3Hlo9AzT4LrrN
6TNYxWGGUB11AkS8qV3dy2pWN1xFhtMgY/dciIrlV+yrC+eNg9W1OTirEccM
f8ejfmGtF+uiTW+3UD7HLEY1tgk8/k4rKt8G/GQhRX1T0FBT5EEvo+21+FbS
0DO+SDgjjaFGtEjG4tk9AIidSh1hPBxi8qG+ycQomwTOmuuSQuFFbVjeQs2y
xiKFdC2zZTd01iTU8jfpA+cracyoemOdIW6qYOBix/VYwK4yhv7N0jL4kabu
ih2wlmbD1Z81DjKK7OBcW3dGQ6hNZ8rp3Db+fXZSGcKMQxQBXaPeEqJAlIdu
bgwPSA/mQqmZD+HcXsLyonJG1e5jaSvZYve7gklXzP9rkoKDZPtjQI+6wZDD
ofkKxGBatpXliVKkdxvoCIygs1T2/2FMrR+hvvHZwMUR+OVInlb/pySrVqr8
EjMrwHh85oIKZeaDNlJBJJKB5N11V85Tmhr0R5uN0Zfrmt/xYTJqKlU6rtrl
OgIdFCkNfpl3a4qXru5py2X1lWjT+42MjSQhRLHuOGLFHNWEMr4DVYdMW+5P
1bzRLZJwfdO2aoqGKlED4DKy8DV3s2qjZC2mypGb3WjrcuTFCCq/cReCXEDL
mJtEAMju99e2lPqFH3NYthg//Ykv6fAFBzgejuHP7aGhv73UdshGpri1IkDp
KAnFRd+rjzAFMNIGWRViZly3p3wfbaEWc/WhYRmD7zRQl8q+qUt2NAmjoAhO
RIbB8fqLSN2vkxuNHVw/5+bVeGWhmV94ziVC8ZdUFSsRF7EdlDxRVABqo471
uM/fQqj1sUQ6vZ3BuLG6IXjrJ+NkvPZprzJRKAywevV+shK3sAA1L99G2Vcw
/aBjo/Ml2FPIDyDzcXirED3c/tX/5EQV0Z6tKUiWzXyEaU6mbMtG7yerEQgY
Ip3XUe2OiJAa99383FD+bgfJ3mY8qp8riZUwStptvrYw33lrDOGl0NU/BHer
zC7q14aNGHDsXaA8MkqOT5cHudey3S7+0+l/W+9+bJedhbN/wsxRjd4wUEGC
J7HvvUqQTbKqQULqODF7lFZES+WjPHCSWE+ejHeNrTVnbwcYi8PhDRwjWZZ6
WnQ7gRcHtelfo0cNCshOXUlpFZLchnGJPmmu/TPC0sslV/52hDjkjV/tL4D2
o2mjiyCwEoQHdbM9Fxziqus6a4Qtk6IBs9FoF+v1VkyCTg0bepqgm1rG8ggx
/J3gY62PNbnf4J9D+nfYDtAmfL4ubSk07nEQbAkZQsEeM6tSU099VW/7ZLDi
DDD8h2Kg8Cdc2qdESwTHeP1QMhGi7s1cR4PwwxvVVG+uDyKmZLBuJxmk6pKW
1axhQ/klbTlu3IrdzizHaK86Fo6p1wpat8ePe3tTDTcsK5soJC5bObC2gaRg
Cog3s1NW7nC9NBUp9fJPS+Q+P/Nre4PhTgXbApEMptGHtsT9gbmsF2BRqH+K
tMgyQvrL5I06liTij7xoBBxeHMUdsyI+avNRIE+v1IGFNH1en0neg7YyW00s
t0xPYQuRar9UqORSUHXpJ1+NiPkeV5J1di55GAJRLR6QjQtnAw0I5R7L+G+O
IJi3mngPD82dxfBjHfzWYNJXEj1YgeWoWDdfzpyVT4Ph58WuHiLG1yokV25Q
jGmBoJrmznqC263fE5WmR9w21KLi3d+NRh7cPXPSDUyWPRLWyInxKMZyaxmn
RdKu0xcOoTLJR5AnX6jUM6k4J+Da9MovHlm2KCI7wLUxprqdf9ahGHMoNlRc
Zf9PXVqM/L8rW1gJUaOCBcvvrVIc+TyKc/8LsM0sdxGybIUIg1L7rYin1J+V
tq/UtMaL8lPqzeCseH1DXrGrMOCySAqrl5xi2CWKuX9MGaih6TWIU6e64DTs
REr9zs8fakgdr8faiQOkd8eo/qMG8lwfW4Bp9BMZ/nshsBIppsGvZoPX5+O0
f1vcLPuvlN8nX4R7GGHldHYoMTXL7ndUQGVbrOeRio0vnoOCT83qfr/M1APC
Jhv4K2Ry7CvUjxkYJfGD3taOFELpXh9PZevD7BqagisijqRiTfvm79snJR//
C1GNQek1Cy3FZBDRARSr9bks9EPMpLZCxw4oFSeO84ZVCTOqQ14gXrulcV6y
sgfdn9hVEIOKP7f1B3c9ltmqDNDubRICLhvLIBH+Cz4FZI7x1XwnyOGfn0vC
wRtq7Kn2CuA5SXG+q5XMaJ+rxopkjoMhrCQ6XUKmJhQxU58+lOP6bHG2LGRe
SY+A8mVKMxD//6EGY4gGyLN7fS0oYANkO4u+1XkMG3drYgQn9RqUACYGjk/+
wAnnagMtG4d9byCRimcZUvP3Dzd/+gZlhWvDMftAKhyWGBceMMWmVazW32AG
yNvjhNnkPGZ49VmjG3g22C/SWkvbTCysnaX32QDLTADMIEWkDMQK0UvK8SSa
su034jVbegqYUaaCHqZVbFokvR+4X9xPETdh1wVRq17mQX/ScWyY46flr7nx
ulrSPBkNPXxstr88Wlv7IHmfiht3POneD7rZFsT63w6fr3hBymkE7ppdToCV
WtqjHe8YSVqF8TVoMHfhG8UhPFER/WD+Fs+RUNYEdRX6j1ohB6HLb83K9yaY
rE3BxJUoQwT5V/Xo4Xvi6l1o5Ia3dm92nV2RSR7EE2laT+p09qkODXbS1CxS
Axq/6H/m9LR4MJn2R1DDBlsSXbWJhobzedild0cRU3WEg5F0HJidayYoM3jR
FgN/gYzY1sF2hbOlaNaK2dgglB8GngnZOAi5UImFBW5zYphA/N5JrE6NbRbF
x7MVKqiZgmPXwBcFlihd1+UJVaaQy11KAtZpVs/Gf3pHru97FyNq8TrGd6tb
9VGkB2odV+N52JdVzx3xjYY++oLP6rULq113vi134s4+A0M2cVzajboiLRkn
TwBih58B6JGYrqMhviIohrmFRJWsgR3pVgEpBqP9wFo7NeT2J832llhfyWpe
0ScRt43R9XIzVKkcbUPmngc9pjBr5ar4UFZaxDRgQg31tXQARmnJ7iSMtavg
YVkGZGgzG164oMnsODTPBlSk459LC9VOJ7Zd+igZoDfXQdCQlzktpzpW1oDx
Bo/bGMCX6Le9oXFlRYQtACs1j4ZsFtstPIahSLMznjay2y9Dk+coHHI3M1t1
W3SR8S5NLGlUJ6S+cPpDDCJ3VyrHS3nfkXsopMrT2QWl5P9ugKcJkldsGOL5
e1Ckz4gERfA9AZwCgzGwlxLLfks0Twoql1du5u0dV2jEQj5qT4E/GgdM2Hud
w/lVA2bpIX9VhUrCBag/V5N6sWBpG+c8pj1mBOS3Z+7ayNKfviycRU5yNnIJ
r75cdcMZxsWOMSQD6Jhr1W2XrLfELPJdaBaQuJXrUgvSm5/IcT6n14RDqfuR
syOYUgeg/20MOT1cke1GSvdcVjm02cSTHOMvzqVosVcOpkg/2ut0Jc6AV6Sw
wOUnI/eKJwy4Czn+rW3fYG/Z0myh977nhqMQ1eW2Z8ZpMJCRIZ8diT8qFzqn
EAoQsldafnUDsuwVuLnCczDTGlweLnWrw3S+zQOGdC9s5zYMjHdgqoGkfkt4
pKG1KLA5EAOAJzPg03HTh2Z+6XpCsEGWbnBkIdi42RxjX69vaOmTMEhoqMhQ
8BNVZZeAHfFZT7tjESUc/UH7/v5Q8aW9pIvtCK2QxR4Moy3XE0xCVi6btL4+
QNs6j2cM+Munv6S/s27JichgrPhciePIqCxIBdL5zpY4boU2KSMREe92AlKf
DKd+bvmQAeNfjzlCvouknWFVFovhuDE7C/Oli6k3aeR7WO8DYonMNEG1FBeY
vs52835ZhLkP9P0iMibiZos5dgX9hntT/KUPQscQnFjFsuLNpVvE1zI11d4r
E2A7fDS8sFCSJrwjMnRKqi7YsMzTITTxldjyh1ONa+ZQzOBmU8j3pkm6FM0q
SQFnfR39uc67bWMcx4xcWc71SY08+e659KACA141sM2DlJPWOPAkcXWwi7Da
st4IVTc3ymtpiRgwWzHba8atKfs7Mx1cXcc9u+WV66+uaNq46LCMKKESkOCs
jdB60ydGW0fd855FiAgb/vcMc7GS7LrvdIJg0bXhoU3FxUfXpoladcSnn5Ji
ROPAuu+kmKpHbf6ksNkrGeyP6/qgEWKjXE6T0KHqAiLyy9Ul3BJxJzsYl8Lf
ulrxVcl2m1UX6ZCUWTeTSoH94fQK9PpobaH8eFMwMiTyztO3VS3f31b/7wqi
/qbKeV7x7Q0Z5m7o6Zzxp670XXt29h1G+d2P/ZKEObYqPYWFkKb+bDgAHJLI
x958iQIlURZ+DAja1WFNDAW4KuQ3HKHTX7lpm/xGT/2D5sOqOL7YQth1/X8e
xPczqEs970fLoVo5/KCtrJW9rgxXS5IyDVtOv+y30eIojFu6B1NPBgz7j5/O
w3DX5UJDFJDLiBjslmxOY6T39RWJNORXTW1REyh6wiRdXSqvUiozR+300Hnd
eQfbK5AWOktdTgcezg6IwIb+y5pTWkLUeHXPBxoDG2hbX1CcW8UPsK6YoXi7
n+L0Cw/WZ8fW72ojhhnxwMSgOwqRCEIhoQblVKnhFb5xK0x8JroB+0EQ8R6A
x1HwyUdQweSFivLcmcDbXg+49hCsyZhGa3H9sLk+NhuyzoJcz21cuNBPAEW5
Vhr02NQUQpEoPnI6uczt0gPDgWLTnFgoLWfaVlstn6xRz5F2qHZxfV5YgCnf
IJnx0QtGBAZmGEGFSGeLQ80KrjrRFSsdn2hrSls6OGuPr6BKhsdQ13yeGFK0
ggUsUGy8ulq1JwC4FCBJjZHF07JhqyQKTXilHZPjkRAsyozERKCZkoXjJtDM
JTMLVB33YK0gDik/4l8TF7WNCLaALMzuWVZaPRISyjlQ59UPkiau4TXLzJQi
gihLqLSs19ixgE1Fxd7O9zTFgRaAIPo3zF7uCqzKp3MGalQo2vTpxOBzvhf6
m372iuE4kkIpKgppWJYvA+yF1pm5mmIEN4dbNFv/odrbDOSdJ0xRbgLlr+Kf
DCr8Zb2ofCPV++Uyfong9vgQf42kmGKXmaegg8ETDy+/eOEpaFTUoav5NPs4
rBKoxrZ8MlO2HVCEDx+E8ergVqsDYeyD19Z7cV9Xl329yNAvwn1YHFNFJNuZ
vPJAmA11RNGmv0SE8sWueqdrHKRrtC+x/MGFX+Lm3sjg9MMcZO4KDtcOldqA
AX3b3kuR8Fc98PB20NozOJQOLH5DwrJqmIJrKFJyrgzAvX9G8fJkdpVBrIcs
Y+BByTeBVI0LRCHe7VpEYyQiHJ8dps97b4pLUrS/+cDCSDDnw4ckYgonHtjB
SyMK1QTMCd522Sema7wQYIPxdbSNonXcez5H90QODsCZZQPI5HD7WjrmqZj4
E7ywftqJxyhYv3OtmHKUweYTrMJNiqu6imfNcVvQDQ0BDJGmafFA54j5obBk
Lovis6D15FGP6MUROrx5+GjDA/UQVXdy6QxyygsSR3w2n+Tfsnui0bFH8B1Z
9wRyGdIvfIHCYLFgTlUuDxJjeNCM43VDnCp9bv9cwgAL3qpzb9UvnYoMDeec
aP5MhKZPvKS8cm+EIYwztA7Z2zwJ7aoyCujgs9W3PJImSPpO0rUZLzHv4jkh
/7cSPTtUl8mUevA4EyF3Smk4Re5e0QsMgHFb1HMf3HxEWc1UIqfUtldO6bWh
JNjVEwHP3wGXNz3VHy9Mc5dV7TBDg4Pq1BiyZEjuVZOym1WwyJ27hITFxCCG
u7cd7IzjzYCwyqGambvhmphLX35GQ8NrMUZ5Bvr4iK98pAg6ok84wZbS0Y9Y
5nxqyjG/Gaz6iLR+PLPLbQjMA6Vp8IEI/ieAVdvNYrpW5SxlUvRrLlIDag9h
65mU1LeDmIarTvlGlhchtYl07Am4xkrAa0o/BYn1yHBScR/eJcoWXGmXxdu9
dtZUVtPSMftUcGeoVwvG4S2nWLHGROEfUyoLMpvMgkkAGyPY8btBlFbApcrr
2MVb2HEfvwBaWom7bGy4XRl8Pz5E03Xa2CaDdMdjDehcVHSgJOfxRqGTWMJz
rDn7lON84FFT2X5H4b41scy7MRkpQ/hjNzZ/ZgWadrVHRATu7/t9deinjGua
PhAuF8MZ0HpsUACoBoSQU1KuPBi6T5BDjniEgQEVJP6e86523sf7xfBYTdIq
gqmslh8yteuLBpegoMIIwTfMGxWgKRhx5maURnoC3g5jDl8jjhHiojOOFl41
ij/AXwcZhGwVTDbr8VawcPfvN+cxrFHbkbVf/XO40hWYDwzQo/QWMHVDnbAD
94CQ/bd/OZHxLxelzgpiaTc46Cvb58iz6/sB4iHOiQiC6DR1ygu8bDrDwqGp
2q+rMLV+3I9PsSaPmjFnaIrRz7iEowkY2Ms/JCSV9wTtXgtyrwQiLdBkA/Vh
6J6buq+OGH9HCNBfG/+ivoyD0sjTrA8CQrlz2vFr0nC7zTE5uyCdzPJGhS4g
7jmz4W5PlI5DBIsTG9bEkbZmvlAvIhu7yG85FXbFW2a1tuvJYVC+1pHpZEiK
im+HovAYesazlMh/lsQpKJES8utZAx+LbFP4fJ77TyicObm86/4G9CBFNEMj
lU39kk1zDv16WeyERa9IzB6iNPQqEtXbsxvQc3MfH5hdT0I/rGoorRtTy0EC
2bjIxSwX5ubpwSLGkVKL8WlwbAer3ETcXOTNsoDUQdoKouQ8KFJhdg/vUugw
ZW951CvVOxZTHFlsqWO5m4wc7gDulUNbcEEGVgN5jLqND/yn413lMO+aUPNx
VpPkXFPmAHNy4WgLmeNKkL6K8Bi0Xak7CEw4koUiAtAiw5JngG1VbicbGV0R
n4E4jW20NeUqmjQnhQXvWcVoIMWAQsWBc5lXx0qTXLt4xF9VKZqJ7YY92uBY
LGO5r5lAgQpGM10m2LAtmqcANXyflPOgmd56j1nctBri7wgVYgOEVJ93Xk8A
VvHoqzz28b3RVINPVbf6XjczTRDCq99BMmrrhQGQbiNeqb/tKpY4JzVFzo3d
NxBJHRgbfPeP8sB2rpVPUvnMGaa77Fk+EFxNPqjgHBh+aXirsG6psZ5xZ8q8
N/nI4bFTg+fsddbLElkatvseHwUxCUOJ/8OaX/ULyzYYWH1tpFTH6oXkxIH7
j6rZG9uwg7PaVsR594rm/EzgZJH5kVzZHtmmCRP7E9XgwL51mlIMsctcYhsG
NfktOq9pIhKdL+fj6imxk8/GazJR250Sj3EbK6RnnyXfQROXKCmcfTkBcQmK
FPkT5a6kfhbdcod6eYFxMn8FSEaGTBZjpv8iu+LEcZWnB9k6SwMlpKNcfn7x
1S6N47ItDSIjPkHmbW399gKJg+vcS7nMiA4hhwMXgecmARSbjnzfQh7TUGoe
OxVJmvq6hinFoUQLShkEPAacEMzulgr6NL+6yAR/TNf3gzscs5Wf4G/4gCSS
biM+nzH0DqCx+prGiPyIhJr9AccxF0SploJVXqoiN5nk53azsVvWS3zim9B/
Odx8ovYLEd2AvQt4MIpxzj6PZGkXfPZm2I/sQguZho0LpeOsHwb7xB4DgUtB
RLA0/ZPUJf1rmj0ZtMeoa/xqwQlT49de3zkBBltG6OhqXVWWKfC+GPfLkZN1
wsTpIjfUbHC/msC4YZI2cZtaetK0WDgf1pLsDEhsvC3xUblOLihkYVfbTUSD
IWzDInxws4K/2TR1/6lkQdXTp9qEj7I+Bffclru5nIddzd/3ZreBjHt9kGo9
zZCbZGPgTPpiqb5HN+l5tBORuPszVNjKeG+xOicSQ7t/mN0+OOc6DGBAPD5Z
g/skSB2D2CASvZimGJc0LUAhX575k/fIZeqMVlxa6elsOHkT3fmaJ3yXk1uH
jjUJplECOJG+HL+K9+4EvP3nJljwpZkXk7WK7ljKZz14CQtjv2S2nFHpnF9S
T3MQ8AvfohvOPnFF5K7gmyIDymaxncJOjgw0On1TMJvXsZmIeiRFecID9ymf
tGh/BLkkcRYRgh3R3FpTz8Efwn/VMi2EFMP8vN0+chXJ9aoiMnIn9O1DIRPq
/hoiTAvmF0xJ+OYzRyd9i5LUppnwtuue/RNhD2VGXic8ovXiVEWYjZL9Xhx1
50Bgq0nZ7ek1QDE0QMXvbwIzJiXRVKAwjC4uj+rRe9r8YHRmoQY2YEZq14UP
wtn6EarTNfaKm7f2YZUiMcXiXPTj1pQM4acsLk71F+Jgljy/vZSkzeF6WSLe
A6W2a1rjtUVuu5KpgI5jGR+IDsLxa1TygFzzw927o4i69x8xa+w93Z6pxJrC
3aowMS51sAFz0rgoZ6russ8WbM6LSQRz7i6Y4ARQo9jr6mu/WGzgtxmTO6GK
PEK4OfIirJBoW6IiZJgAkvtHfu+GmJU4pejc2i+ZOYmrwf0L5MU8/w/6TS7P
T/qU9ELpl0qFy+kmhwMFdusc0uTMliR1aKtxXyNnck813SFgsqwaaOhBMIQ0
8aLHm8A78IKWdSFtiKH8o1GnTSa+dWkslgz6B/8w0c+4/fKsuxgca49Zc+dS
hAzUBglirBrbngG2rTnT4HPy0jOZQ4olNCYCqd/E3n+HNdESyAUT1Bzuut0Q
GjJjS4k6cz2KnttVBCOULtKl9KljFOAXYOU/7Fdh2EsUNUHKXXHW7k/bK/Vk
P0O9JFFKF8v/k0isDY28t1SmbvsT1y/nVzcH0BPPlBWgohAfRLhohZ+n2j/q
lXAKQXwy503MHyldEU4OVDFZ1mJa3IZfCvzSoUa5R9ap5VBeOLUkPRFe111y
kH/iL7POC5JxmLf9ZqTS+EkVfl1wqYua2YmLLJBcISnR08WhcTfo79X4Q/W4
kv8mVT12mXob4JArOuBuolEmMbmgidWgL4Z4g9YVJwVlyH1oUkyZFhnmDcW4
OAYclw5HuqWy2XYYXLVyiR/WajAE3Bqf5eqmEVrQDEe7AixUvt8B0pIqD3Ij
wRUFp63iG24ijs5ETW1vW/UxNnIhKmvBMvnLnYUEtk5I0EgOOR20aGzq5BS2
FZvr6DOw0zx5H1jm9KK0WsnvLL0bfSxJqPxWwWg3ZqoUGF1EOIKvIe7oeHbk
Z6Fb2iDwUU8BxfzxnGfX41/yVKHaGyZCj+4KRl3EAP3oURXx4mZatSGPlf1O
S48oe9sK7qNoMbfi8gyyI1LN2FP6Wk86ZN83wouTTwvYqJaFKpevNCQwvShl
cmJLSFt/i/o8ndTqqT+ocjyXXpV9OVs7KEBjn4Cop9ojiMcs4Ud02CRsvX1h
dhIip0YKx+nNvMY2jsOVEYoFFWvdaH7gfmDM3SvB46yCIk8Iayz/ecKNc7Ho
sjPg96umN5nKMndNUdG5RSNljkx+Cq+FfT/nj4rGgyVxsyASL07fh4Ugpe3R
K8ktWbGLGkqamk6sTGuW2g5ouv68fl9N1OrQtJFcXz7RQvSA+cPVSfY9raOQ
dg1ACjvlXtErfDYMtLaD8WhjnXiP2b1Cd5aUbhIKkwgvCn5NWMO8jMBRQq6R
ObeoOyWcrXsbGge/1OIHGNk1zN76XUqgsTADzpdiD1k2HxxXhoMKrYFgwZUw
IitcB/HiCRG00f5EV+Eu0xn8g8wN0+PjA2ANpKY0+xrXXwGe+YEANZdLeGE2
bZqPqay8i2cmixZc5Zm0A2WX/mY1k5ReJ5bySAsChBZtldrujwvhEeSELRsx
FC5hxOYYhWt6VjP0rJSOcFW4XlLv3IyCPaPoPjStXvr1aIz7bu6JrOJaxXU8
NHKzwR0F+Vb3fE7T1fvWZma/+V4FS+w7Z6ZQMsR1wTHqiiKM1n4JkLGM2FLY
PXGb4lj7QnChHzy4sbGJuVdR1zfaXhwEojwvuir7PYji9AX6rUTxexu608C6
mabUEqEG1YdAQdnKrlLyblNZtawyKo7wKlR4l6kIO9TgFLUDTQo1R2o+RmIp
SwiEgc3m1NtLDo7Z/0EpBEDsOvsAGnIc+BzmPvP0EMtdCe9NcleqRHmbiFch
+BnJR713+WOflOXGcee4YEykp7ZM0jTZv31qGb+G3cJqLk6qmYv96tPYBPSE
X0d6PP2V+KYvNW1JU5aa0K6RzYVaivwq7vUsnpHdumlTvy3x8N8PWR3VzfIW
1Bh9AVMtQA5kTDG4fEyAOoXAQdNB/puedImTHWmJBrYfcN3RKXIwVG0N7Vo6
IGAe+KrKdRZV5eUmRnERPr9I4k8f34O85f6pO5fGYZD4PMm+799wI9mfIoNa
u/SDFRDMfcKdpvZvpW0zGbKTUhILvrlrixKMph4KW5eD2u4iUsR/4vYDniQo
t8Gzz4CO95/gEBUuOIad4CN+lqyC3Wug4OYATt+7Z/jIDGmdjl2RUPYK1f1q
K6BsJLq/lqGknUc6Q9A62Itpim/tGXCI+kUNsAApG4PxOvlogCjXqs+nxpnv
KIAwqvWKArdW0Fjanm9yNXYErLLDYKzcMPd6Euzveu9hirN2E+Qvu0h9CNvy
LzvtEVxKIilxHHA29gI/+3OMsuhRtiYF9zUsj8WqZeacAcN2kCbTMSEUnJH5
PgVbfwkrtFF8SiguwP1pnDbp2fa6V6ejQcMo81MzYoZ5jKC9XeiK9wL/7FS5
jdeYtWJ7xCC5ciL7gcHGt0KN7Ok55ANygzrilOo/iCdPeZntULCtJpmKkA5M
hCrszq/HFFyJO5zdRy5qiO8O2m/qvYCErfPbRgDY21ccgtkSF6fBCx5g4mz3
if/P+mdnbfjtcPfhUtImm1Fbav+gA2gSWK0gXzqcYyw+zuXu1DeQYCJ+h4hp
YmMAmuxgPQTucXeMhwH3MyOVkKgJeER6Mg1y27UeGmY5qh4WYUTguxYjg7uJ
AwKzTKYBKV5Ketojd+kSDvvjqCGISgq7DoO+17sSy4sUInFcoRtL4RNqtmnY
MszX3QyZljXm1lIrTEyFpGrYYoT7DDhCtxv2u2mDhpZHGH///QeDfvsLtwkD
G+J+g1Z6KozBGZbW4MJ/S4p8ublxOJtQmiO7gEcZ9HdTN5fkBe5XLsrfmrWC
Te5bpXkb9GdKvG3rrqU21AiChW38YdkgKHN5qVO9846mPG6psns5NQR6Mu+o
TXSKW+zR7rk3fxoaO8qu0eOuRuYp6ya3MzmDQxiBsZ2R/iLf4HNDijjLtLsO
yZk0my2LjBSkKjXUhweSbS/tKtw7a8rECJ8pl1lwHNErMnYCFTluzkOc3j2m
E2roqDTK5Yv00v6ZUdhA7CBSzJLcezeGUJGCrDK6W99GsjTaO6eZIyI0mtN2
hEF7tgLxTJfClYHVyIKYiKKjl3dNJ3Lv29qiAREFixMEnECMusfgzQM2tmhV
JkuYhoXmUF6t/fdOoH5OV+P04B4EMc+ecnAApIPaPpcl4ISLZhF8teRNeU9h
67Y6qAn9TCHL0Ov3kEHf/FkQQ/IvGP2+S2TT4fo2HghK0xtcDZjZCI3tvMDl
6cwEDQ2pCk0PTg+4hSrLcZnjMTOsFwD+a/xV6GumRq1VrXL7o+X6HQec+z1P
O43TJaMG5XSbsq/rlmBIRvJ/kWEAURRG6J3v2/53jiilaGGgv81FeJPCrFJ9
6p+LB8GbZEgMPs2uiIJv8ffT2V/163HCISHFIYDAcKv2/ifefbqGsQUZUrrk
8Ju8MeSxZA40nz/4D+91hQNyv9N3EwJpDeyjmLtX5Qarp5jZjKbbcOzAygSs
0k81RFhVkfUyNHZOiWu/FABoLnm0qjtGJGcxJwLE0yfSDPaiO8G9ewn8iLq2
nDslCT9fZvIyf2fUHqsgvjVstxCAW8JlMtIPbaRej/lXb3jjWxgI4sz4rbU6
w1iW1mX7owq9MDkZ1Qmo6XkENaUSZlFprsE/UzCYzw5GWR4e0mINWxUVStlq
4RyFKKhuFPtk2J1CBto5paDnf9akA+gUN5QccPonxKTuZOD+BfqdJYA+44Kg
+GisyS2nwV+8h/cMPCpNxEYYVk2huNuWnSPakUtJK/shSGLFsCMb7J0dqbpQ
8QED22ty206/2gv2rTLtHKD3pMD/jw0/ePT0RhwBhYZNApj73WXwIxNbu3up
B0JqCpPnTpClGMAn7m2762RqVoWLBlIm7RWMwYnIc8/aLwYSTfSQ3MO/6I2Q
lW17xV5uWxpcQbFNU/nd8FHDjCaTnC55WzQs5wJ5s8Z5ep9cgNozA9mqw/vn
MBeyEzIY0kMqBeefsjaA5wiUbfTV55KcwB2mpjH1KH1LysT3MI53bJqGJVlI
4TpMtCRZ5kSe5pKWl65iUJ5aINZ68Ynj0kPZSR4gEyji6Oi2PpTWpgLytjTO
P+dGVwrjXL79HjquuHAXE6lQuJxGA1EMSIRRzuXo4/RHCPNUljlH7MXhEYoZ
H5Kkc+6IJdPSy1YMvHZL0z1s5+vBf6Lh1wuUH80J+AJGWBCf/kMgvaMZMmUp
DDSzUBHRjBu8Mscbjlo23bFjCciHAJDMMgqwuJhYRQ16Cyfmd5odzdLmdVwP
Dv92hS0R+pGPtDprYf4zJ1JdgA4rA66kd3frnD//3XtOLdt9P85+G2pYRou9
gBLC+j08eKKMptQBKX4NyRDri7XjdmY7M3pXHtROAjzkZptt244TgXLaim16
Uy0BqV3o5jt+42PynuaC1oJ/H1O8vuJYHxntZjJbxCpDlIOHJiMArDP1p5FX
/cIcPaE81gQRBv36M73p2qCI7PmvGn/OKQwiWZ1HSkqtUcyZOT73RE4u5gaV
FCDR2DKZM3QxQPC5zQXEU+MkZFbR4NY6gbEINfXMPRPvokgtM6lei28b8Zt5
omxFF4+Vepyl7P761AFds0bzpONi5RwzPPpfimj6k6fnt00gGrUWzxfe3Mfv
lNuKy44AmuW3mj3ItGh4ouXpTA5PfykvPsdRyiw/IsKT/Jo/rv7fcFi4J5vx
yS+WAViNXOV4IC09P2w/a7dyE9SnzXfmTlCyw5T0fKJFvgTORFUFV98iGtD+
AqSJ3bPqDWaL1jDkhR6j6KegZuGE8IJrAuVcGpPmPC9n9NA7KeYUjntrRSig
57xa+k8L6AfmHo1auISHmcJ7myhe5SL8g3756s+0Ys5EWI2F9wnkfXt80af0
QA4V9qhQ5AMpGP1NbnhVacreHdP7uDAglS1KqOHW6gJalXanKUxQOmG+gt1w
/fGlvagylcys/L8dLVmKJAgbHkp6HQbdjt/mi6q5NBNRtogeefD25m1ZfscI
85Mha8HemdCkBaZ7tV38RtGD4sRgJkWfh+06b/paLxhGmu4lYA7sgGDLjR/r
6jiCnAteLV0/uYhQidCD5atM6yTSaa2JOO+C2fJvd5zhfs08BydxYwpsgJmN
v8UdRWqIgkXvxSojpZMRKkadmEIg1LqQfqIKXCxwyS1DvDUCZPTunwhQcs1Q
GUm/i5rnslRWSM8JyWhs6jMjrdLcM0MJVmSmOyT05VyhmZWglxLPGKtLkCTt
UanRYMy2FaCcFokKMGDUvhushEP0blud4oNG/T8Q1IqTY6WPPe6eClwT4bEU
IT4pI27QRYCD+39pp4PsJ7bxlNK8Hv6ScGe+CdnYwObNuhFJrMwfcN3cOc9q
a8e3uVT0n+dqXvQ8lCTaM6dFK5+ZvryQRpqMbTTT22YYFlSb12Db3GT1ASVy
pG+7uHWO1+Hp7moHGx0LvdQSSfNur8MFR20IagKiWugxOPktcbx4RFuuYrUT
XdnJ5bElpdMMQkaRSIb9PMLKOMMubUqNmBaHozYXO+J8TL5pSJURHyyo1+vT
WqPGkfkQ3vT0A7wyx6+mCXltK6CjC74n6aXxcRWdbdjGIJ1jb3utYxkSuZwC
pBX7WLM/jJiSESSHcLuvFKu+2qi4wxhO0OY7KD93TEZHElMVxVC5nmJe9YUo
fB3MVKJBTmbwWhzUlbiKQpOSlCIgSqbySn9drT907TpfS2ftpLUdLOxPOXDa
qpYDeaY5I23IWkkfpjCA4vPx8QEBTISiyIL6hJZdnqP0otxYfQpFFPhx5CDs
PYLTAs0JNGzTFGGBL8g1pBkdEIGKnhSetyy609IGez/lrHkv7yofJKPoYnd/
RT2KNsz+Stk2zSBGU86g/4P0xsJ2p2LlxHc6ZV+G5NAowgI5Jlj3er6sSlgm
BO+OhJTa6g0quzX3LH5zOdfVEbuuNuFCHQnNkEK9cndH+ZKTFsi5m5HDAukA
dpflAyeLBGKszHOz/zVS/TMKlG7f51w2n/GLUSWuLFEWb6KrmFRI81RUI1Ph
emEqKhBxNW0dFDLCTA1/229knkit0rgEPGhoOMdq4f1kdH8JIVKXtjljg6aZ
7YXddVPLW1VUvGHCtW9jpNAZqsJ7DjXiuk1ka3FX5x5iPcTMLoNhHdnBRnuF
AcoEfmXb5jWvCd48dhCz4C2eW1Nrr3WLPEJ8B8w3vbXadTR3aNNkXJwz1YC/
bkLAH4eSA2UqEJfYED8Y30kxaQts+8FgUJpt7/pAI8wKwMaclEEO/4MewFsK
rD2GhNvCh1YnA2hj2UNc5/NOBFjtlaiBN4XYWdWYqwM1A7vt74tThBuYiG3q
XAWTQU9WwjHc+cVYaMDze7Qda4+alHM8Dys1lzdP4w2jRekGs816wuzA9Tyn
yoVjI+77Nk3t6hIsSjj0CNx6HHissxCxue9IZuAUk2fFggtxwCJwP+gtKkMj
9PBMDQQGpzxq41f7Pk9lc8bj69lsnQbxM87BgQOUDawVowrYkjM2O409oDNz
ExppHOlwpiNDTz78wAhZsPulhDpeib30H1wa3YRPeTiMpgDo+3bJ8KURVBGW
7+byF2xgfNWCazSWNpPUUfssK81/sFOqwETRB8vtLMZ8m9GIx2j//eEkA38g
jCsF+K7t/RPVWSHrEaCGvEBl/YEDmZSrfcUR5m0mkw5nRAPwOTk3Izva8S19
DCyMV7SmFft/MYhKy0/V1GK6tDUKf8AREqzEucXM6TZjHd5l3xxhVOlHVIAF
5cowfKgWSIaEp5tbTM90CaFK6EYefreiLAcVKSU7ye4q6NxcUAwquzLxL/Sj
nKir+uQhGoXbQOwKzEGQj847vJuCUQXRZNaMK0OwrtcJdJFlljILdLzqNWs+
2jHLyZDMJzBQYnyNBkEVNRyqLf/J+BSdeiFeFvcLdBI5GnK9ZCHcHwotM6iD
QhTfO1IDnviuQn5IAju99eDLGG2HrFBGor+H7Ud1sWrVaOF5ZahEkQOWaY6H
/LPdyhJrgh+XZXDz/DTfGkJ+FN0Kl1upULQxOKjy8XwRCxjxVpdRoCiarmfP
PertHlLi6nlFTzib0bRVCjc02khdGSn379XGQ7cthEI/sXIOnfnJiXcjZ0/b
4CaDS0JebWgX0XBZpHESWQDFADaCzp97fTXoAgcJ5dWpYwIrQ/ioVIYvF072
UXWZ3pd+C/MO+OkMmiBwsdP5nOSH64eMb6q9sIRA4FUzGc5i3RjZJOw87GpQ
qu8BkGfzAufWhUqMEMMyrDmVt82hl7JW5/EyhG6Yty/EcrfjXMfW/Ulc9CPJ
BS4xZyW55cVn7XqX787QcKUnYPwsobY2CkRj6F5zKpfYJX/zXivAa9S5Qfj9
P7VoxfaFdb4vDSwRvBUFJVKREig8ZsS7O+TSIACsmKIGZ3EXrHQexZ2OMxsu
n4OYtYfKjgwtDQba6Wh/q3+rNgWmQKmHD6nSzbRc36DMGqu8Z0Qpgo9t51Vm
gz0YnsjoTLohWCynP64WfCSeEnfZtZg0rHzRrqVSEX5o3LrcKf+948sKEQAF
muGO0+Er0KjrWrnZO744uFEX0bMyXNn0DBTRg+i/7vKtrcI9mRBqOX4bitVb
CzghPfiXATfo8aL6fH+ai0LUccT2jxxKku+M3lEm7AkZ/BvrHyPJInVMVMri
WAifszMGUaw4QuKiLBvWmCf2WoxLW3GLBDlUcVhUkKKBraHj69JWCkHYQBn/
mtjE2jMtXorVZZDMyAIxzMPOnqdNl/IDH2uHK4fUTmHDeLKbHpk4+ftS4OXX
gJE9Os/xCLcKC6FmQR11mdNHCJsalqL9gXhOMhLzoaPPcik6svbwX+kyP1ds
Tv5hjURiS+bVBGksKbTAbWaTnbOSSh4yHs99jVgZgDgANsAGxd5n8Y73Cw0v
tU9hI6ptX6iF3YgOYT3xir7NCwlW1ZNcYnxFbOJFOG5in0Em9t1xJVTmWT4N
32k8ZerMwydIHgkTy3rqkfZMvfLYKifftYeGzdI8NQUrwSYPd2XBJQ9O3gNy
VlBeeDGENonYHFd9WiLvO7bJOwjKAu6O7sfKgdgJpMoa3mmrWZL/Tn/o60/Q
JEV38CYxR8Zs1EmQsT5wpbeXIhAF4zX2YJ7vjH313zShuA7ThlOluv9EA4+z
c4/qmm+f8lPlda+XLtPqqWAWiT2hkIXYtKdEfk6Neti7h0MJNQTc2maOguB9
aX9knQqnEiO1nJk1jSgODJ6L+1PH647BRzouGzQYlDU2Ep5oSdzhmg63/HCG
zQhttoe4iBEuz3C3cdJ/AM0XaoLhpoAmrOkkqztbzMeJdQ5+Derblxdp4H9J
byobmXWC1SRCIpnc9yQf1TVIL3ZeIaNAKWPzI/Qwt2nmJF7jpxVHPBlSuPrN
eFFy6qECAoSEITvVr77jqSzmKMkJrU1kK4mfOK1kVBHzQ3kEbRg434Dx1Mcb
MK/5zkzfYSlsc6/VYmUVJsXoMPAG9/roJ5C+IuuU6D4eqlj6l+m7r2hBNRdk
vPFo2lbxwInTfq2S5LUNvdp50UmoFFSbAjn26eN0rFYHqx0SFdLZUBE0qTRH
Y3ZPRKRjnGf9MgZX75EzjMmKkcqUhOSK6jTapxfQBF6xulTB8yrVnFUnBIG0
Mc1x7+5oX5n6uo9xLCxRxRCgGqM9pjxJNYr71vaAxyOEzR5phWmTLeuXIVzU
/B9hZuWyoCpUTCqkgNcQEbnFIChgMpwDPamdrgxe8/I1InA7AcDzGmnq/GJV
GeeN1HIKcCaWbjoAC1hfIMRvZRwI1XamIng71/O4CXcRD1QmkKNEJc93tkhW
fqkJEDXAbGLcD4mdMb+/BUUMlCCwrCPfD9DCF5Fn2IKViJqFkWloHx20hLLW
97OSfxU9kne/28SQxfUkhECMe4L6LrUj/r0oxueVuwOI1HR2P4yN5mLvGxPR
5QIBHvqygI76nVSxDqpH5lU/3TncdkpbnA+w37PZCW9zvYRsyG27uyDK92aR
X0hCp5dU25ssyUVHv0e+XR61YFOzBnmO3LWJ6QjjCSpFODN0RMCyc4y9vFnP
Awgl39OIiEX/7bQvSqHTd8z+fOmFnBQPowOH/GVVx5ndhlllOgYbzjdVD+Xu
rdHwe83pQf5ggCmh1xHWaSuOSfRfYsjthOv7FHffmfxannwk25xNbSCEdIMm
Svgva6xpDhtuiZSjsFNywgKqzLC/BFDMWuG2QfrRSzVgzT/YkavroTcIK+WS
f8M6D9WgX2j6oucrw7pQ1k9FxrCwRsCGsWRLBMPFbzYcMJ2doltB3iawpbLd
gL+wZO12VGDXtcNAHyi/tyau63xa7BmlZyzY54vWWOxGBtOYWCnMAEphMFsr
dGMqMCDNZK1qQB2abEDzaRPOfYqBHkFtU1PMwjC51MvhXxTvGY7gi3m6m/ri
hgtovPfPZbmZBmRD9A9ITMQFS7x2GCA/MDitMEpO+oZdYtJ1aROhggbf5TOQ
3LaqvcmM6lA4N3wNkTGu5/p/naqJxTtBH1MSamio2+K6krVg5WZbt7UkhEIp
hh4vLlfw9fou+iL94AYoi2Uqspved+bsBvnRM1l192qTrm429jCdtlQ4JSEC
QpX7CDYiksJxX+v887yxzfXd77Z1j1Bc2vnSJgl6AEfo9AZbaq9PqgOMOPd+
FG+JfEjgkjncDcSvMIv7O/1+HB7f02suShW70bAOWibYqAFFBQ//jY0/3R+3
eFZsW+wuRQ9kJevka3uGeMILC7R6XLgZ5FZK4QAn9zwztYM0+vtm/xfqwzP2
Rpbe55OLIeqB8mGdjW5A37J/ztebioTNd8ESfmbZrPmnQ2gYQwuV1S8c9OCR
111P4Tc5Pd+5xECzRzBNv0blLMV7Ix+SI7t+cC/EcVkyZiiwcRITM9QRIRbt
ORX5rZDI4dr/ykvY3Rd8VJGzPJZGSww6cenrdjMDa2qg64Nd2bzjQT3rNxOU
Kti1QsIxlP8b4dTpvrN0Cmr/+ymwhhEUG7GCA6CzTOyO4VQ7A9H3JAOAacSI
G0rBd/OGnGGRkbIsrUqo8zvUakNslgRdnZDNOMjWFVG3ScPfqoVcZi5UBdPA
UUz+BOrLwIwqcTJTFeNOhCvD9X4+nEqUASlF9m4qrUpHxFN14W11ROMdUsV3
ea5fwn7DYIPHdtiTYhZL8soDg+1VYHrnN7otJjr4f4UUfxP9kzUK8nCzQKA7
0tHw4Ie3pFo4ycR8VUWHb3YnbgVrxVnKZ2ctikB1C4ErLr6y0dPSjjivsZuU
WnfJafPf8u7H36Udv8j8AtwPLOJ/KcnPArYzCiR1CUPW5urn0pI3Rt7zQssF
rRLTBo10FLk1ybxPjxcoE7+yXzakMrG3ADHZwJNAkrcmjCSQghq/sJsMoakE
kLiGzoFTvNBQdbsSS6xRL9Wp7BxZ0kZGe5rLDEmoH16IDHknpPqQikwAHkax
RbZH0yR21+xQd6TYcNgn2N74AiGC+i5c9J82cvfymhjrXvcQQXmOr4CM53fy
lQNcfmWX6BjPO8chAaVAAoaTRpBq3T6JJSmw4vrxj2OhmfuYLq4j+XXQxEle
xvr+TrDJmZ6Cx3VwbUCyRmb2ZZv5PMcIoMHuQL1pcaAUuOH7JPn7UPJwAR7j
1AbMqxUTPcU0CFZH9rSjh8KwFTxJ0Rox9OPsTeZtr/7tepuevYOanixZYYxf
j7l7Ov2HhZF99WaeLeQ/zjDFdgRQc1+s59dlnL3H0md/oAw4RI3GEiartBQ5
e+tmzeLGytTWOvVG6kodn/8Wga4c+e7DSaAxdofPUglC2J0u/B3lquoUbvzZ
LV+H1WGmBOObVN0Q2MD3fEe8JxfCFD4K8FMw1UlPiXjzjQb43GJDuWPSOykz
NxnobDl1mqtfK987WljXYu99KcXn45UIthmNGfTW4Tpw+UeQXsp7cmzMrVw3
wHbnVJZ/qGt32LAuTzcQQLoqxGj7PEhcKL/vNDrTKNcLkXcBpM5CxUEgxfs0
CKGdWLQVv6RwsOUDVA3J61VoxMtjGjV1ZNFdp+/FBRRXK1t9P/bYYy0FHcIK
achOOyUvOk5U3jHkppcLYIXxnfO5ZwKVNJKHWfAL0O8BdBk7HgXGTRfxiKMJ
ApS1dlgmACud0S9mn5viG9n1DcisZGdNrGvGgMB44NpPXWYgsbauOhy9PiwV
J0K1Ws8Wx0xztfiPVKxC4uBk/5qAfkfOkm7MoPnEdC6QuzwQTT4nMQ6xW7zF
j4/MLTVUdirCA22nXdtnK36cKmVgJDlzEfHf8t55Y1iqZq8zaOFcaWnI5EbD
C4BkXGE59XS0s8Ikpz+7zbQQPJfnutZMVtkakudLRu8Gi87YdAhzkqXvRWUG
Gl4B+OqUKl5NGloD4sL+6efUpFX8sQ4DCK0eRD5w7f2ROMTSRPQkEFrpw35L
O9l9Fft65xi0cWsdgqoY/mlx3K2K8Tg9aoCqTlFYQzFOobNccjFPZvdGtNOq
FxQ75CGzZviuBVXcTQt+sqz5EPrk+/9kFLTt/FCr7RW/OxP8Jg72LUC8ukVz
N+ZgOOKvKipEmdcJyp2ko0GXnDed3Lp2qX+hj/qshGgaIzv+Sh2UveodvOAh
43ojhswNY2ZrQ19tQLYYpARkZVx6m1fWpjPL0LCoUIr0X44TuHenvob+PDL3
WbAIo6GPP10ggDGBlYYSYnPyoW1DapRC8Y6MkQga6hA6yPK9UNIbxO9jEpc+
sprP4ADNUMf7aR/tKdhuw/yxCuuBzJcc+8dyQwkV5I7XstSe6FUwL836EVxP
ZA9mB2Zpox33spYhSAdqefbaYyOG43uVU9QRqwp6W1xGEJWBK4ZOOq0xvB45
VaWqVaN5ZBzneN/BZl24OOazwDQdHtqlWBluZJt/QMm8OFAJ756gfeJVeu2k
TStKc0Nj8quF4CqM5aw2CdRl7DU/aUf2rTSMtUyz4vq+0feJ4mgzFElCP7+f
VtuKr6xLJtu+ngUULhdD9/WcUpOcC7kH3mPYNV6ymU39+DZU0I5w7hRzQ717
rILWQLAXVQwfoolROjc3TUhMBgLEIGDPgI04Pkp+HMNrSSS0FjMEa1SOcTS7
iSVcJg9e6YE4NQ6p+NFngYZJD2iH/bEPm6RKWZyC68I5gFAs7g0OgcbX/bs9
GM76g8wrNtKo+zNPs6CTgCOeYlMp1bm0TEE3srCLJWKGhl017tiHMtZt4m/7
2bVisB9fBnqsCIYLdC2SkptKUkpOk9AQFwzcU79cWdpfu94YDWpIqwwoyOwN
5suRrc4oyBT+MFBunVBMjO/WLEe6MqjiJscUkuN0mqYZHY/SBSoEZtNfxWd+
Z+XbnloqYwyUhYepQL3aWZBmVL4Psn52AWa1dKmhFxsUxzqiizW/doDDPsK5
G1ciPsVCPpzStGqhYH0QvankcPm+8jEzXDV6mWwlqVpQjDHAZXCRifkgnFlL
t24OvFx81stJ47Wm0jc91OSNWv4n8aysRNDTPUdIR7brxGPkXx5GzwIzO56G
kEY7f0zLhQDFNNvALQJZO6bz1Tud7EMJr0lLrnPjQft/M1T6gcg5fxj7H4SZ
tfX00RH3KhC/QGi58q1z37utxrLVkW42noo64W6i/f7SWOaKI93Y3pw6lkhz
ArOSbWsiPVFWNPAOCPKF8CeIwj+QCWnVDQWiJA3pLTL1Rq3w78eRDXGkIBaP
oBqaKjsHjtkgPuX1zb9qdwq+CVCKT8nkHjZYyVLPV1D44nfnSEtzqhc5bKqw
0ibzQDym0hkgesogKtMt6QX7Vi/R+YOlkDDeka5TUv+6iDVTVDzbNL+/5/As
JUlq67eutPJU0tfPNmqsS8xi8iffAHWxpHlE86mvo6yiealxOIx3fj3GGLle
zSlOCLjPQKT2BpD8MqWyRo1hjfpCetIQOEuLLx7Ms14q4UvngxWsTtYWZleE
Fvoaeh38CQQWYEQ9R0cPKUbz1VV9eZWkNZmcdztR0ZoqiCJuKG/gMNdG/Dis
iussH+B99ajzkpkHirizHTjAE4i5kDlmVy59eGoAgL+3zC7xk7q6F0njp4ed
JD2Uq+TvKipm6rRf/nLtGkCUmLfrQQOFB/rqAL1kcMgcCmw11mJJCu94ng+1
iyL0/pAgql03mCzwLmGEqhDzyb4lQbMXGMz89QhUKWBaKXX6Cha6gqUiXXqn
M8bhRo5SqujH1s8UHsYXRicnccN8YnYPJK9HIi/B3VJjHTh7hRHzRURt47OM
pcRPci39TjqV2Vj3RE342qIDAymsos2joHRbXVqoSx4xlu/HQc+XYyyiLAC+
0LuE8A1D0RdxP6iLkXC33waOT9iyZEfpRq0Z+I5gz6Bc7A44GusMVVzRBemP
zsRamx2Z3RcYhZ9gWN0ls9ZnBNDGVvgrJHaFpGDkR9Cux6r4nA8zt5Zz4k2n
2V2hIlRIl5xCw4g96LnEES7HY8x9WAX0pU26qjN+izGTlye/vj1WdNPLD2Uf
2i38zFK0Tc0vvrqT85vMmF87kGApdvqVs6BXLWyya5/gYA7+ja4ilBpIkFsH
HqsPCQnTuXHJHmuwP5tLhXVSg4iwHFpq/KOMdt6xnDPN+QFDkuC/24BJqiUq
fBug2TwP7ce8DJgJ1untUmIF4+nFNzZQY/VffnFrkHbbpklz+4jiLYtrgyaW
W+CtV3FOu7yKIy5DpLlX4M7eOG70zOhUuu/gz3iC99oAyRKPrCxSXY8vE/6l
wtk2ys6hw97KRpKiJ6DOaNczW00uLOMdjeoxZmoUaMOCmeRzqdPOJKmo3E9w
7XV2qDxd8irzZepe07s7k0bXUsILZGeeFmsXxWOikuIoNiyIqtuKVrwvUm/z
EaH1TlricDuzTecO5yqcBE1jFeLBpfhKGd+OgTDq9xH1XsbGwQwfC6Plz2+G
K95mHSPxeFw+hYDNN0xAY9PpfxeD3WUfxxechjePVmnXEKB5kyxN4F+RSXPd
0sEbbRvDmXQkTKWgMiGo3mypbtcKhA4hhltUeblLts6m3rsHk+9ZRWxFLJBT
GzNrXg1WUcO6f13Il9Nat1fwlevzKvggjMj3raqWfwZVx2yU70hJSswHBgK+
oNscp5Dyl3cO0tP9ge8sfQUr8Ui6U6UUABJQBlv65zNG4LlC3Bw0fxcEJd6L
kKK6aFzQzbE9kNqO33NJSUYMKYte+KnEHJ7JWp+zkA8OxhY7TLpoT0hKLh79
3jyw14dXiM09baBROPp2Y6LvDc3eh8mZjqLr3VE8AcyEW110au3ImPlOfaPX
GWCVghQT2G8+0ZTZdN2RrRgB1oVDUfp9EEBm5SyPnc6USTmf7lp++ScEKQkc
I5KkMg216UAu/yAGYw8gcEhhdT+YoZhsxCWgF6Jithor0Z9jX28ngpeiOshy
lRxLilscNwqNau2GMrGDRrLP42Uk8SV6MIVNxigoMkaV+gT6qoOdTIpLnQw+
u3l2YRcbpc7wCJXBrxQwy0hFPLq9U+vFy0BFxOlE8wOT/kJp/HwhtV2R5ko7
cILNM5d6gnMNAJd21kwX80VNTyeCmhnYJ2MV3N5wjitqjMp8aRhJjCqhJoZS
6xx5vEZG99PlRfdkthyt9OuJNVM00+NjtUuP0eHFnAQ9WIKXs49xTdEgoSvE
oKMRT3oGJgXShLvcCNnBtYv4UTQ+EXprcKTMKcWG8tpDyUapSAhce40uvsrV
yhSz/S7EsVsfoPzfp3bWgVAzYRIx+9btcPqRPsxSBu8fmYz19jD1mrCFsHnQ
mPEIfdlmJADv7CdYVTE3TBP7gQNXDP7qA19xFjEyVowGyQWqE5AboFFEdNIw
PBya5N4VZbNuyRQhqwPGojTKBpNTUOBcAM9Hk9TfQCQu6X/fOfB0CLkbZH+c
VFVRSf/X0aLM98Rr2Y1sKrGOiYTVmJBkdMQcLsIHjnZtwMNVxDDv2wAkhncx
aabsnHBqI8YjbXhWkf5X6cYSS9Kpd6rOg8LuIyGF1M2BmPKQRIxIPqSU4EKV
hrTEWXrQl2iGDKf26Jt4zNGrdrcz9LVD0GTSHpfs6xSoRLtLY7uZqonlHPsu
bzHua7qYG7i3AmsfWXkDU3OeeaSbRBjl1YKwkX6YVKTvEjARv73kMhIMZPHi
S5pI25QAmoWz1Z/k/wM3t752aNfriH4ufwtb/MwXSzDYVJE2q8+SROtTVNgs
ejmokTBAmdRrXRNPwGp/SR1Kzh9ycx01J1dWZUw5fZdH19KWlJoCwo9YRDTC
zkToaS17VpVMcx9huAUNXqiW2xwtVrlf3GQr1DvaFCGY1feaJ/UjT3p3HKeR
jPx8uENsYI4ZlLMiAqte9TnXY8VhoAbwV4HJC+Mxqa+kyRdVqZ15LOdwfg6V
vOix5NNPmZ9myQzTjnRrXF8vhozBTdRbfdvVHjICjO1SGp8dM62Anvq+IRY1
1xLNZEQ8Nm+bTR7Il83dITaL+udl8TtRbUQkyBPlOp4AKitwQ7B8Nte8/L+9
qcd85OcQSqoWEISJmTw5a4oyj9olYFPwqDJBXDCZvcdglBlI+y0A6g9/JKk9
ifimavMlV1OU46gBnvdDKVXXajyjNDl+rNaASZFieb5RYYM39LBCV5zCQEE+
uLvxnmzdfk5k1ouCg4WPsh8A06lyTzeR5zZ2WL9hX8VVMPAjR0WPvWFrj5Ht
xdaKp1ezfP+w2RMRR6tg1iZIAwPCWJgu2KCzazObvBi6ghZONXkOXIiJF6bp
cvyfEw+uq4f7pIAsN4Iod4NBemFLlFQuJl+GDZhpz8obot8GHKTdqVIrXFA2
sgJB3wI1EPO5DIEW4rwOG9Xfz/sZggFB2h2J3FySgXzaC17EHUdM47zUdjJL
MoW/sytQUbvLPJP6FJm9AOJvX2QWE3Vj/Hg90YAn94Ms/pJjBdNOIVvvdmds
IW1fvbLWDnUmN70LnhN4SfA9wEW1BHOYXJ3Kpf6pzzGeIgi8Fnuz+Awm8IaU
vpFTYEcjzsicEHKh3h9dD7zhENqXtuT8r+u2+udjN/epV9zLvTfRIgNPwOVA
BLMk9HKfa+6YN1X4lnwh3ETuvjHjH2pBImb//bGpsdv3PV6sPkECkUiyx4/m
pcDE5Z6f6G4zeYMqoK65VBJTo+qoDK1f4Mzoom9biRCdNbdoB0FxwDgpxfrP
YShck7RFkw1rlDvN5SfQEUCmwurxfTR1Ty6cw+jxibbaJg+yGSRLciX1T66o
E6Oewyi8uz5NXsSRPX3pqMETnPWxMkhjk4jRgiPWhBnnRPhgaoNQZdg6PWYp
pbFRs/2bcSwFz4pnxjKDGVgkEJ3P5vLu3wx8l0vpTt6+lpVvB2zG+b8/eFAB
8qHgHmtfGVaFItGFb6O7Fn9ltvv+BS5WQKstig/lOvD0iO2hYKP2NXuGZugC
d8XYTRJ9DFDGyd4H270HyfIx73e1MEZ6huLzbiasQmLE81T3UTCTBIT51ewW
qUi2O/s/UPndsfO3/0HtPwULNgBdCLw5zQUv5WnWoEBiB6v2FtjjMjiFWqvR
/iFpqR5LuEGzj1KmsdsSaZmfI/4E8MKGPVIanK0nQfkxQUH2/eRf1uyJi3ck
sl2l+HKul9cHpW0985qyPKgCm9yKsK8+21vPwXguVP7UpWp89DFPjKfw3QCQ
MpdO3wxu+jH/B6GAtG2kq3qgmb80pN3pxCBHKQRR3KQ6BPFmICoPqeZt6bru
2bvzVOu/X5+aBFvq7dHkXUumRVX+Q7xpZTh2MuWYuxszMtSnny2vq97aG9DH
7HeCy0Zm4Zz2f+5VUYu5EL5/urT35JGOZl6DP9MP3CS2RmOmBXLjye9ysKRr
Jvov0hXAnXovF++4gvVSZefO/d4DBUOTVg3HbHywsvwjKoFhDVDOVIGe4pCM
9XYN44X8xwUc/5vwz9+1HvexrHktjhHNIw4YMvUOz76+KI2SQGzT6SLB/WWd
CvTcIEQaXJLb4oIslnXGG52jp6E3w3+eU9dcv9lEbI4r7TwkJ0AHne76z71J
p6NK+YJUfr5XjG9iNY2tQl6CYKmP85xXf7OKF1YXlR+AsXv48EAJl2UCbNxA
e2/8b/pBF0U6HrSgwYuI33zic5oaRfXBHPeS5WTHQwaSzXGEKeP7ggJvcBSi
aQxOSt2fZ8evJK3geKqHNuiJXEQYrGVRnUh6ENACSwSzODjF1ioYijUltZev
T4WwUPkMWacleu6uhVYBkrmUwff5j42cVUAdtxFHOlOhTOXq5h1Hri9KdDmf
OCPfQyzYJo92fDd+OlxcUPkAOh6/LU0i+efkCokcKvM22b/3ix6aYSf7PzUt
taPAuL3KF1icwShJOhu3aTfE2JN9tQmV9HXilB65I2/inIEQPrHXFVvnPwPj
nbrPBOgVmFTirsqOp1kQjNwLtf/d/CRZ1ItdobIu/Awx3aYzE45jBNcU358t
kvJOtequs7UP66MLA1R337OknMyWOsc7WH5OeIfLG4QOL8kgZICeew9/IBY2
htAVL1+CUukQj73zTnuM1V/W3ZfHgi7WTXOdbALUPiDUrS//ecGfVWFjNrmN
4xJyEpjMkiXgL6kJrzyNumPYL9KR5tQSC3TZ7GtpA/GpsEB0A43VlyQYaLN5
xoBkvH2uvzwP89gQQ4OgOHXeJwuES2cwBc8Rjk23UG19EiXOA02GWXhdEcsm
/dgU2pM2fqlBYy3v+V7PDeCPbFzNJYlvFbuR34erpudZkd0ux/VC3GVM4Y0v
qW6+C4wU0L7daKX5l3oxURk4Gr1+Z3LixzbvdyEHVSDwSOauvyrqhJQ9R7f/
ohZO6Y/aXdhzKfJjEm+wp4k3KEes0YKju8IBn1SMKIAY+/Tpg7hWnAPklG4H
0mYeAABQnG6p35D8Il7SokxfwREnQvoE+9u6MJE/ZDcJ6KukVNPn0NDeNpyE
sPznSGGZ36Zz+yotRcxLcwiwOOJRy4aolVKxDUc4mTSGHgsV3SApCU98FhV5
Jn7YYrkudYzfMDUJZn0GyyK8zvKS7fj33rZqVmJriUnRMGwp7JWpaUq8o1yz
rNIk8XPMH0sAWrf7qg0hRNx/OvoH4dPjZYcMJohv9JDFeIWpijgNHMoHSPpJ
HGcATpde1gc5C29dousXr1WTX6gvK3nnSj7bGvmwu8u3WYZE2vcGfgPjVAuF
SJijMqlwnyZo1z926BFHT9kNroKZDr6K7YVpgYT60GUMs8rWSTEm8zwSCwqZ
YzqAqqT8/ReLrUuS+LTf73Ixsiujik0iAX/PRirEMQyBnViUrjo+voRSMQoP
Nu8gbx39QqbzV3sH/7+7KhkbCLmkLbmrCOFxqDzxoWEzuvKGrULmVtl6kV5L
ai+JdDcvhKs+NmahrbbU7uev8jMgERKxTrThiPG64gH3vNFaXUwX6B3d6xom
st32kJPfWm9Q+0fe6vX7j6OcVGW5uMypE5gv0VUDzURHLEwdSHbYeAey7OMK
VD0yVkJyoZxwmJoaWMrXu1tgLdLajZ47JhyuxYVF5Q5VyeuvM5N9IS84RzHk
FUXlZpZYpeejgZskeK++XhKgkq1qOQP5c9obSlZUrIBtpnjR+V9GYIl0iEsv
UPuWILCi8dt2AIhYX3flGG2LJzQoUpS9FQx36wEDrb/ERY1+JOkL6t7dM4SW
OINvXLzQs4nct9PkFYp2IbBN57MefXLNjV5XSql/rb2SdpMp8cYPxNEafQm5
yRYmAqGDYj5L1iUKIiAuM22I7eavKaDw80YzvIL/EtFEu6KbLt05IL5xDFyF
jKIeAZCTblBD7Qtl6JHLTXFX0wPDDgXvUTDq0s07qE10pOnw2RIt6VBh+XRW
iH6fjOguHzGBsjlhI1ixCHXZx5oDZB8xzBcVfnkXvRU3ebJYyoTtwc3AtC+g
pBAtCU1HJucdbSU/DDYPNou4Q9RMlL4yr3nWlhyJmzeDhqJbwJA3qUJdNDqG
lR8JB3u0FsjZCOwiHoGhxqVddurKv+LhWerWMxFuQ90GsH0D0VaEVbt/uR8j
21XcT7zINHrvmamDe18WsRMAFGFBxtlnOl92LdrB3USjm2wTetKWAGqs6B/+
LyreJ5XXhtB3C1a+oGWeQ8sJ/ih51P0UIBACVVOksuyV3Dy9pwz5vO2m08iN
SrBXN3pu110qOkmWqN0SJUg9LX+3AI4vAXcWFZgv1GtFeIYkmAe7oq4iFc4O
KGftdKEK9TxnnMUNdYd0B/WuV2kh9j3gJ6gb3MAWRbwcEOXVu6T+7cFGpqtX
E3+ATkZnGCRUisheM/4EachKNveX7S77supTgWPbbD5I2uVLwhDCO5d6267d
eFQfr4GaxVKrg1eX6rBnSYxHU7TcMN5/JCbxrfQ8Tmm69mwhmO2wx9LDdajj
6cIucabbY9VXcOawXt/jBn3vCJ2CEfJmSlUj1NCw0qTr0zm7OCl0y9MQJ7wZ
xRIJWxM6OHY/zZMsFx4y9qBa2UI12soXkVq7hl3RhVA9s3jJ0f2POtWEowrb
Bbhp53NzIHEKhPGbKAZU7SpG25Y4v46J9jc+ZXHSUxGo+6PDWY/b7CYAFkJ7
r3poMG666FTo0k8kmIxI0bANGvWiA60A2oNHYHiqq4UeHB92gXajuKw17TG8
P6OMDnHPFUGkeKvNAvYI093Bei8VDamcocoXz8Hs7hoskc8t4TpYGvdFPi9h
wTz/UjaxNPyyPVKXkAoLBVYDdzJ1v/1w8GQC99kuvgShBuTHGc9OdXrluDxL
iUwGCcXD68XEXl0C4nO1rBm9nDitQlZibcWgRZyyV+A3h/Nf5kJrFV7ybcXG
Aj2siKP9XDdA+E4stvFOqn3w/AscFNuKdy9/+wAB5w/AyPHeWyflUFlkCEOs
0zc7WbCmeigmDoa/Bset7pX6AwVpFMbR8n7gHxQdD2ozCuk6bslB9YbTzD85
liYiIvtEBwiBP+M88PoWJO5r0fvaoaPkwiT767T6/jqHDaJ5K51koz9OsSBb
0G4ixmbOEzGwosG3FWICH4l2wTrMnIN+AGNg0re+j+jkugtzf0/5QN2vcpYj
NqzNmDDhc0xC6B67D53J9m5VLmKXb+NPHM5vMSx3lRNDaFfYHyWK4GrsHNpj
AoDXRtq9w3WMR/IVxKzP11Kqts2yY5e7HB5hfXfjHOmXv0mFiHRV1v1JD9AU
j0f6UkpzAQs9Pa+DmEkEHdNPzvvqs9CkvdGqsZYoD9v73QPWtIoAPm3E3J/Y
Yak4XpayJ4HioJ+wAdGGh/wVbkTQYY4eLhkukbpB+ouzzlAY1Awlvm/UZT/x
+Mx3xh8bOn/12HmDY6m3bpn8jM/qlUwbTYbVTczUMFYH2TzALbh4yLQJvqoU
H8T8VtnBJe2v1NsLXn2Ty485cAuiV34jpqwCQ2naXfJoNVPdFUQa0Xqo/v+V
IaJpZEmW48+su55fomIqD5eJ0Ib98nOsBUlsYKwKhT+lAh6E4otLJs2h/9UF
i7IbK/F91pkAXl9JggzBBCtG3dCSxLPQw9kcMKRfs+kDtsPhg5QyO1J6AEqw
LCOfX4mc0C3yRc0+mIzCaacg/8tiyWWtOVYFesrrTiWmGvJSXeTNvKKOe9H0
J4np0ZMnolTUdraOJEXRGKjDEvgRRTJqFE8LxfAofZphvW8iOAyQULXVlxNP
wty9nMe87x5YB1pl5KVEhCPALGyK11nn7+KRgdowEk6UshSLk45Th62TBSFo
fUENA7l88VeQFsDPDH+42nwfr7e0wL5hIYdzOaoCqXJsR4nEtnKV0UqtYy+/
Q2w3MQ0hy44RJ0B29GJ8L/DAALf7P/HVV8FriTwSpt/8Ed6Xy3NifiYJ7pmP
mynVJAh4fmNxTzIz4hdY2Suouz8YhnZF+5tK6i72Tcn8gmlnkb21Y9aHPABf
H7plgXJxFyazZHxeaqbiVdXs80sVZv+DquNTkk42GbGsnE2Gc5CJP9zDQq+p
cI08KlX4FntH2Je9mZAkapyF+BKGiwpUrV16qaIeaBqaoyO3LFtVWqujpAb2
KNWRmiYxRdRmJ22SPqEQgHCZ3cXidwgQs1PFnVUbF3qFTw0I6ZaICA6nwAZR
GN89nRihMErRBlgv2CUXF89imtcQpB92ojR54FwUvw/ICyNDfZgU0fYBtkuF
Lc5Lh+JZgCZ8z6pV3pofROg/lYEIFIp5kCrSVNTBnRKbmZ60JG7cKFGoSa/D
fXyyOZVgUmTjG0syd5upBsEG15WyAqSYSln/3ae6N3WmUI8fui8KwBlfiMmx
9Q/54UCQrAAmyiMKwVHeNOPh5HtixAGTNcZ4nyzxv5JKjEKdjpKs1kOBUZ4J
tcwHDaaGXxImHsaTN2EMZr+lbgjrHbu7rv8aX5ARZH2Y5pMPOjU6qDZk9d8x
Mun31hhefoOy47vdI0mRUy5g2lUqYZo9dex8vHJGvAWn5pMrri383T8PKB1X
t6LKgUlGok5M5xAmBQzJpydqHAlAnaQTnVfhNnK2sF123uzV3hxkoi6Zaf1O
M1bYzflbVidEhT4bKNEmuqiXvFPW521Hm8+87E5XcGj9IxE6rrKYH2jC7MFt
MAkJNCHNgGLibIapOuFSHTcaOF3S1opE7DBimKFyJFvKIKYQR+zfjdLSkU9P
3wJbTM4esUwoUfrfdAccZ8nOCRYpjRFuNbIXhRBw+iBlH3FKy9hCwQro8MS4
6IVolSHAI/a5w+H2V4xSBHp08AXVHQahfCk05kOP0nqCurAx1N3Oj0vfRgh5
KMEvBrAxwyepNvAi4wfHzbze42Xq8/IGA+s/1WJOqNkOCnMQtvqZAQJgQsKq
zvCRY5/p0iMtrJPY1AhHTSnBB/LMFQnFTYnUa34E2lWcFLuUH08Kkz7GsvvJ
23vd9UzlDfVEx+6ggGUklnTB8g6zz7v5w6IFZSuGicRd8PLWEhKezOhb93U7
mb3aZR95nxvYu8c2BBydNyrrjnu6koRWdPb7JDUcUB319jcq161ZWwJ+rt1b
twF5L5Gzr+HAqS+ga0TUa4sBy9WuZgGgW2Pchg1KnRUloUMaM477Txd7TVNb
HhK5/kEB/ji1x9fZOrFRGGg8bFgAVolcN1iywB2VKCRm1deJQZr6EpgTBvaC
jBkmSvy5p6mX/cV6H7NhAwdURORMz5cWeeJEsVX/EMF5IkKzBogQrgPk6NFR
BFLSdQKC/awKzl8H7Rp0lv5L7+Fkscq7YqHoUb8YThFEpuEBySs0ckGr1R6W
da/pPmYrLUsIX+mfwVEZRqbih9RX705iuTO2/D74gZ39t15epFHxN/YSy56c
CiGb3WbMembIcbpa7HbgzrNdeBJXqNe3KK/HY81SDhv5med2h4UYZZ5faSXI
ICSL41DPab19lvyz4DfUyqcAUUhwoeDfhrpqnhPRoqZn6O6brw3omj0a7usM
ElU6huUv2ii4YqVYLgwl23bocGpZG/+nEWbhin5Z1pWYLZzsXvW3G91oA+/t
aU6G83Vns/29/zH2OvTecBdc0kGf9U0S4sYZrdySL3zOSJgx8hso8uAKm7UA
bfl2ptC4pWEMy3qycHiumSeYw77xk7YBnN+quJrTTZcM0yV7V9eKXXYQ/cQ/
KnfGr2U43Pa2qmouO8lfksveT8AScgcWOKWZ295vtvlnxPs+KP4MqLL5jKYf
zO2Q4Rv0fZxuxqJNdF+B4dkhNLvS19nT6LyCQ/VEJKLbdJZH0AmOy2MbkmYZ
1Se+zVQ1kZamti6MDMjl1QR+zzWegHZZ2TW9/Koj7s8tlyt6i/5hFbUE5+v4
eU9jGl5tKB5qmgfZm/531FtvC/OfDYRckQ3t+KuaVu3d7crkddgMGcBqaqqP
gmM3rl8G40llRRDYuk2mDFLscgZC5Me6ewRNK9t0XrDxg5RDD6JyJw4trevf
DYIsie+5daHTxceTYnI9z+TNb/OI6FhXD7IQHEEJQSg1+ho3bZLBOUoLYg66
G5IYXT0GyhNeZtwghsl3R4/cEUfRzmONOv2K9cemgLOg8BkHs51xXpbY9VFz
1swPVOKso09d/Bl++y1fllVS2fccge6TN53VTnBwhhj2FJ6EEj3NTMLwI/Ln
jyg1sAi6rf8ELW68gL2Qoa0td9J+TfjPB3Odx7tsxAlu7eLHlKwZGrqz81VM
Tf0qn6+P9TEyy8kFcVZWTictZk/NINtoXiOax+vysyMOCJUIlcB7roeNdtai
3pxWJl5h7D3gp1I/r3hT0b28/lgPmlqbVZeI8NDzewCAUTUDDYi+RGwIrn+5
2OfXVv0Xui9GjQm3nfU+11qFvpOncofFYfdImXReUFafgqC705ZlQsSDHmxy
SY5bPRJH/pP6EIXgy1BZ3DAZh7lAGtx/0nfj/roTDtlIMKEIZ1LSqsMGYZO9
SFuRTMQNrY44qmG1szLTc25rX9B3/F+y77WL++XiBZ2UizkWnzNZ1Q4QKh31
3vIdrk33YO3KXSNnGq10/QZBYii1o2flr8/xa/EwwmCX0sa0b5y8SozTkxne
PEivP8a6kgWGL2uyMGj1gpDBbOkV7piE0ARnziZmYLsgFVQ3TpUyxPqHCsqb
SFkm4dtHl9MMkswS8g34VQaJzrqNE2o/+HkcxS8sJJxUeu/BZWu1friUNZY7
cEq0nOhI0qUMJdSywiZq0DfvNMHLUKDjJ/gNO/COmZ+LvdpjyXwJZVP8xPlA
jXKksEg3eOtDGtYrsQw9jiwZ337TjjvWv8D5quDSMsVfZpXecH7OyvrGMXx4
Qt4Uz/oDD6XT5qpFPdnjoWoHH/MxChMrrkYQtg+VQwohs/jjQ4ixyHW5or+P
mNeO2NzT+vvJrlJT2WN9hlOuTkMMNm6e5AmrlyE+qtO+ZjxHX21zrFobo0XA
yjDNKDtkli4dLqsUAE9kADHjG0CiyI00so2kooaajP0Qi+EkPIm7ytjaCZwW
SqVUhXZ3puBH+YYJVfoH2GEi4hb86CMJlRGo5jXN856/LuwvoeKpzm5NdKZY
zANWutDEapTbNzgiLsPgruhNCZCSfsV7lkug2RWv9TmkCcqPEKZKoXjLDwZl
67Kq/SOfhUsnKsivLntqRToEDKuZqTaldioY1tYjBwvDMELyFB8xKrkkSeyU
NEOfJNXkKMaXCDIpWIoojIfwT8tzzKfo1fa/+jF7WzxZVUK52cC8PZuiNKRt
d0Ak0l+HaV5ECaMNGqIuBu3fMR1Si5XE/v8z9HRRSzs2VastzUkaAWrNAR0x
T5WixTtWKxI7fSVPvAlXHo8YGUJs5CKKrftAD79l8XK83l/4WnSxUJlu3Db7
cNv7eY4E6bL3cB20iWeKgtZF7s02Rdp6v1CdtnYlRk5zqW0cKXn2l4qzwKYh
2If5cnxgP93o8q82X036AmO0rOSzxDIQ3/IqUBSPTBUwYN7nKeSM9ee7GiAF
0CIdd8y0VolwOJP7x61v0wput4+Gr3J+4GyuoqaNxFMVcZuXhf6bMqkayKcD
h4aeLZ1gIfDsMGYhGt34QUKbVfc53zAu6r6fDCGSPW01BvR0AHYu8orOq9eG
1IVIN9NDkIOr73KCdsPXqwdbG6CIiGr+pieeNIgNm+k2v4tKZYPKH7TNRhwg
bSc+/uCUkd4pRP0tvuKyaRroLyuB7b/PtGdIfqOmL86KN2T/Dn2ZDGN1LGGE
W+I4/83fNFmZvyDuVDYlVI40JSgXUwzGYczuKwoyTKUlbUlxOAO0mpv/WScf
wh3fea6UGiysMU2wC/H+yckVf+CE3uz4k8aKDApSnveUAlL++J17i8Q1K0dQ
j0gsMlXzEAabie4lylmPnh/6Dxm9RMMx/ZJLXnzNsSoVeG06TocvyTSgq2D+
ZxWPligyyMFWCGTt4400FvLARBsJJ10aOn361MpDZZrf/4zkGFMtbFIrPYV/
b2tfgkkWCfUvKdT5m2BZhNO7ElJdNGheTk12DXsg9LW7L2xKaFZy/uSSnE7v
vB7/vkNmBerGHuU4Dz0KFYIrYmtQhdPf4reB3nFBXlUrKKgz7lLllY338OX7
w/a6/aaPmUk5o6iA06t7zE3kenLxk9mzuFRR6ZAOQ48lawQtTJO9dM1Dr8uy
ntFNbf+w0mER/PfSMuyCKF0Pc3A1/+MBLdZHU3jsmrUP6ChBZawDXxYBhysB
8QqZq9TwiYdHbLF1X51kkh5OOJAzwYHjRUmGtOt6PPNXytl9OrX4oZv520OL
wm7QhCCKrmipPOP8ZlrMNymMyBpM/ZE8b9w63LTdBto+MEnh3Ke8qEFLnybg
i95GpDB7/Z8UkYZjqMjd7stEtHzFoCTnA7GS0tWvG+wavaVJNTwLNzHcwpkn
jo8Rz3xMCB4gdE4uPtX9UD/YwFJ2u6y1blcTu8fXA/puFJhrZAHwKtMQy8Rn
HQtFqgTEh9iWoo8P/Er56jN3sVYjed0y2xUx8mxVpTMtZm9bxN913Eym2syL
I5wtIA46U2LITwM3Lzn1127ftBwWU+znI275MHPi8AFTQwKtfCLvLglXJHpj
aOez9EY6zhBvCIJG2SgoP19hPoj9pm3PmYOVhP0VnlzWC58i2d8KMBi8nFjF
u9uDD46ve/oVtjKyI4updWGDe7D3q0qNryJlZbELRNDypr7rVUcbGDh2NLIS
5QRI8PEuB4Zft/YBG+NmFX9yEg7vv06H1ybAVuZOh/q5VdMMfN9Ag67Pn+SG
IIDFCHPyV16pLMXf8joneYFS8eFeO4m7XtYKljg9hCA/6vgehY+7FdLS5r/D
t6g5RBaaoTIi4NBP1A4Yc/uJf9qBH+VN321TcY4eOnYHuHnhDvVjvgJVys+6
ISBuDh7sfOxRehgmms6zQWRwTDo2x1TgoV8pvzEjdvLvxLWDGvz3yxvZG/dN
OzCoX6sLSW4euae0rOM4XQFuQUlDp5yHD5xV3/Sy3VEnQcU9MW6eMzFLuUwW
a2i/9wA+hWfJPW0IR7yQP8N/EP+AFWJJC2Utql35QGtawQSaXC2mlPhG+fu+
VPwbrrc0u5Dl/0cNrir870FHu2l0/P8CJ3mFsgipCigwRNcLqe0enXkIoo4b
5CGoKWO98+4+ILr4Xl4MUjNXQ4ty0W2Q8NCkZn2Ajkz6u73RAuS1O5ulBgtl
VAgBg/DYPEvZQV/KC8X7YH4oDl4L958fukjp5IeEwdivsaU1ju5ErCGp4pH7
sKQS/xl4ZKRGg3KduE8O6MZ0E3WZg5k1eY1uk+cVCLxHjTfDbIMQZWdQ44hU
SQFAnRFWF1cy5APQbdtB4vKRYCCRlxCB8anRKMwrrSGJY9UdT8zblZjZl1/y
/rzlI12KAtyfP8WnR3xTSFQUL8JsTB24HpCe3ggtYNY2GPGpUu6imQH1LalF
UoMaRgmAOlJFDasTfRNdm0nyo/cRDTPQHUT+/pKSCKXV6uC7izibQSThd0we
FceS3/Pujs7hIukypkcQHrRHyauomJDDnPR40lnus1QGLA3zjec6CRn2pyaf
tQaJTlgIefXNRix/shwX4kyzGtwqdtoUKDldyDTJo7JeCNKLx5j4o6x31iMr
E14ltDRptLHa6GHjkz6H7zWM/6CqpSDIKUEOt7jUIrLrxzhJsrhBWj5qdEsv
YadI5oT2Ya7RnMcCMgxJGSawxdBA7i33wVmIndGDlEAyjkZNGomXhXgZK/t6
nvjBoqDnDHWkq+P0wr6SJAYUCzHHi9pt96L2kbKj4CrqnwD6sHYt2Dof7lFc
nqQxSp6aZA5BCDZxUuK50X4C+L5k2e9N933xu4UaJlIQkWMxABkdYZflO4hk
ecdpIwhIULwNqbp41ryB/qoXdoxR+BRzI2q73+2KKrMJIbADxsYmeaASZRJT
nZhdF4ji1NNmtgHHrr8A+0H94yCpwH52tmSiKLVnEu4vFTHSiGXnJpPURe6g
/8xnqYFCkE/MNr1t5keog7VS5WUzFAQFgLo6t7NFRoVmJZsWmQ0Yuidvhi48
YwHZzMpkrAuTAQnbPYbvAJ+lixEg81YldlyQcaE3dnjTIK22fkLhN6GKLDk/
OySJWoWdrycGpS6Cu+tqI53xzXiV6xCblqMIARIaAc7q9y5aVFEw9T4OsEW4
w4dRTPH+Sr0x5mHW6PyXK+gDTF/+JmDj1S6+6QeYq7eOdyB8QbndmKSPETei
YjwmpYv70pFXCV34g4cBsCVJx/2FgNmIRPqHEF2u+i5TSJytm8doToR0xNNi
4FmhQ5x6Y58F9uj1vGhnHPv+CPfaMOvLtzC4Y5HCH+sl35j4g5l9OfglUdU/
61N/S22YZvpnKKMv9MZWhcUAYmsRGS91GUz9xPP/in9dxkd58xqDRGLgZAGk
oKhLyeyNmQ076dHSa9ijlQ0AJiyGQIgZnzjhg1Ony6UA8lTEzmaffZwUXD8p
IDqVMBcWFOI6wiJrJUsZRV05ha9D7ftsDk2pTLqPB/EZgDqM2oK0n2U8v3kd
qWJ0hcLN7hULUQXZdwPk2Nd/6b896lWJcy4+HksBucZK2ntQ0hgIePDsRUW9
RQ+KpG3QlTSgWRd1BQikCVwcfdNkM3/rfHSRJggz7DCT/bdNuDWt+mvF2aUN
FUuqdGBl+L1qhex1CuxN0GHwiqRRtpVd9kjw3/OMK5hgOVSxWojNPuhOiFAv
hlhjC3vNAN5lEB95pQqAUmjXLY+PZIeq672206OCfNi2uwAkVuDBMTTB3xGE
6GvHJ339vYdgjkB7PCC/6PQXHKc1M/diqhMB8+eRjPCkObsrCHiTeAlVVvay
ya7bMO6EjfRtYK+xmaPd2B8YnkLiKUbAfoyWGWZg0UzCuksmJnUC+eK+WQUu
I5w5Vhr0yNR9fJVvxSqu+1OQRuK2dJPrW0H1TRzKMeJ9uB0FYeCd2ZufiB8p
CTJCOnIRodZjukFoZ/mXwsxBvPhPJ/YdM743FEi8TL8qlXCcAbgUraA49xY6
4KDg8RdvF+KDuOuAX4RNxJrC5tEr+jH/2BB1FOcCCmMzZeIN/zY9xTY6ISFP
Ct23ieqg7MzQRvenKViIPO7I2aK7zbRqqXCjPMd3EKa9IkJ5YmgKLA93jZku
vnx96ZliYdC2y5tGIl19Lx3TX8ImEW1JyqWTp3f6dM4GjIhTGJTlRR3ZV3R+
LIA0A++FWF7QcEg/ahTR36BJpmUN8g0Kf11IV1vYZhsCDKRuAoCU0Z1Yec1N
KFHMZgWlo0T/KPl/PKc/cdYgtzszyHTinDrt5HHs9Pb03WMwtAy3y3qEtfiL
90J2kzatGi9IIK/ie8ehTIdTqSs8jEUcXiL+FWv0phdE+2Dntai01DeyqMU7
UsK8BlHZS9omXT9kJSin4yF+WcaBxItsGc20wK5/wo9GROKHivfW87Wq9Ihr
RBSEhpPbTy8NUQmcerPzisi2b3Lrjl8jFXOy68KLduRdHsQw3eD3IQD70dM3
26Dhpg+5xDlt32ro+1Xze4h0jCB5hFj4p0Gln+VHRLirWPVbx7Dkqoc0p0V3
42EB8AlwJbK/PXqLpV3QJ74v43bnsFFx8152SYm4X8uqZz4LUpPXRiWGuJdb
TiUHxnlkwYvsRQaGdPQJeNmvA9IUQ324T8apRuIzN8bkgOFP9MREwqJCIuwv
T1PV/MBLIXmbBbRvHontp8LZD8pSVZmzBgmYj+CEz5VST+3nFd/0Mf4gdDFU
bS1M5qWnOrdop9JsBXZOleoQxdE+Hzhym+T1yQUrnz4aY0mS2D5gZQg24+cT
cFetw0rAnqkNyvoTXbpW84pSfKd5IaElbhVLb5Zb1PWIfDSEK87sV3CTVq38
lLL5HOwqz967J+qrwD7e7MoLv0IGGIDeqIaKAIw2e3Te8fvA3d+b7dpTRRPQ
etHziBnr7y54IF6MQJdBLYPjXhgn3ySY29kRcgmsd76z5bm3sm29tDi869+O
ibEnltmB9F5eXAkrBVp4b4u56W7KJtxalaphx3X2Z53Wn2dqQVD5HQJc3yCH
xC/joTFmKV4E657L/OIrQkUsearnN++hgPUjgY0pewBWBCkfVdjvXgGbeUpn
gdg4AmnN6KIFSIJLR6T6uDy2qq5AMHsOb/bjbVQutDoUfBqHDcS5TvecBk/e
7lXEmTqffPsvrwQsaF20A2VACPuLLC9eRxW/yLUR/zG7DEkGUGG4e8/54v02
0dXBMm99dVdjU0PnpVtJ4+GguwIr2Yo45BEvh1hJUneXVBcejcmFpQadR4Kr
6XG0d+2m+IZPIi0hMK6TK3mhUyW00oj8jVzOQpZMT9IwUVv94yx+cFEpxFk2
C7pVu0YEu/EXElnt5KXOmj/2vDF9HTlIhDuONYkdreNogHxwGfnJSqAAxh4l
ojMns0E5WjbsCaLTtO7dnpgVLel8P4/78wyfqN0ENvczWojlNFM0eH0VioAY
F9OcgI7mNLx38LIsU3JpTxcgDOcC63iKNRFnN1RJmCfm4i+aKlfwYlRJUUCs
gT1BQFkGCc9ozzZ9dcSjCDEZkrBkOtfPmA2eP4FVVdUAxOmJdF+DD4Q6xhNs
ORmOafmVHEbUktORqj8iLVTSXCSOxXvgn7wRWFfEU9dACKm/J7dehCd196Pl
hUeFq5XExnO7RW/qIwkJz18jc6PmKNbWGJ4n+u3dEmxdA0jyqWZO1CPNWR7p
8gtJVMuLeix1p3jdjP8IkDR5ppuVECV6uRicmvwbCdFYn8SNNHthnoqqVWoU
wiWx3Dpbv1labg+5I4KhF/W33m1vOT/fQirMi/D0n7kKdRUSubNwEh1g9LJK
9rs0C/DzB99bDLNv8sd80fSQ+Lj1Jh5Lh8qt5M8uwpiVv7Lo1zG9MJbzd81V
pfeFqb2V54tK/V+VMgL+kT/LaxPiBZruab7bnNnO8Fj62SL7bPHRn/ql69KD
2oX74DqQ8CF5m9eIre0dLCQcDJAL4jEfixAP2TMd/Q+rmbzMgNyGgRoKmURE
UzVykTJ4CKly3yHyTT1fneu1Ui5/F/TMv/5dNaM9BkEpwGG07X0a/GdKCdWK
JRJDiMjs3ioK078JcQOtCKlBZ70uAdE1FQVdJ2/U8jb3m5JB65hPMy8b5Ujg
oQtFTTZgET2bpuUTC4I891OzO6TOx2+a9svMvfoqeVSEJxFhXy8YVwD6PIxN
V6W1s/BelfQh0Meq0+Ax6D/CHEqSMEo4l3qOMTFi0pfQppMqzfNQReZgBYE3
FA0sT562W3jXZio41KPN+ZlqbVAP8GKcasQ+laYN6qaBhdjxTQ+LF1n8p36s
PkWQNwSWUtW4pRLlYd84Yk8yIR0vCdaGyko4vxZOrfidJdbqWv20ud9SXbu/
lG6Ocq//vMudgLnjCGXhBrRwv2qgC0tLTdsyDm4e5klvzuIkFTdFJJFNCNJO
l5umkbWr9fYhkFduaCLaU/uiKgj6suJu4LcyoXZnEkJgAoef5lUrhVLguZ49
sFPbGhqNjC0790CHn2Gz6DYhn6MUSMulC+TREJUSAvFlHGhViGDSUOVPrPF0
qCKOgiWvM3VVmYecBzm3WKnKPU5p76vAzRMA7NGF1Qh8SCITUbPChOcJxE1y
T4V645OHuylpp6x1zTTA9lLBv5sm26Uk8CND6KLIvq5NGYzJMI4tcvFbXix7
TfhhVQkP/hgpdXSfUmeOgvLMyYI5fyA/BUGbUkbYA0fzfx0wwsHpfynxbj6i
MTwxxGgpJslr8GKyPQiocbSEkvGIUUWVihtavotSva0m/93Z/EPtNHUPtT5G
S1XUGehe2Gm7tP82hukuchAWbHRw1W9dVqfikITFbGfyLU+p9GiFiTPTU5Dz
uVK5e1NERWYAYJYVOnP7t2pPHKa7dTT9YlWhTYfMgYJPaHVQpuXgepHYb0ub
cGLjP8YSKq2BRnn1Rg/R5Za0PW9pkFWkhgBAjnf9B5CeUwvrF9aXNSQR8SHF
CU9OWYOpZN9vbLiRCsUmlv4vXYwQxhiD/yO3mSI5miKt3X1wdPOnFbKeJ9oo
0yMueVYz0Ixldd4sKaCT7X1UGvTG8Jv2WvoxZplopopRP08EVB2hMAfJjpKH
780/4oowy84Zm/1lOkUlAf4Rccmc6ks4gKCCGZ5K1dgl9Vmqs/twg4SZUb59
wC/T+OS39UNFaL6DMNbsIjMffY//mVXS9gx1b7nqWtGvOswDAsgjDt7IcOfn
/JucsLO8YgAMw7svE8Bdw7LZkOB5zT2TK82CGb5vV5JVplf4bxlbWaSGgPOO
ZHYt3yDe6iyci3CVookbzL6RlfyWoSk7kdOzX0+Jh5Z+YgbEDsFtB6Atsjmg
NmQiEbz3O9DJmAT0PBuAyEWJepJerCPMMk1/kYjOG16hvTvo20snKnlmfAgK
sC+zFkUwJAjn9A1j5uIKfwLSgsCZDZjWVwZCLoQDxpmbT9FsRuZRUCe+tVIG
/P6mS8jrcNRyUyxT6mewnzfokDOFAzsRDcIgKXrCjU5jmkbXypQkWQzUp6CP
LQ0KGkGty5sFM/Gwwses83/9HjNTI4WeTPfS3+1tIeHW8CLr4NGLyItKMht0
x6kxzRL36o0tQZc83DLV3kqxIF5ie9ZL4gAL966WBH7txj1SkEpqTt6wUskq
TyVtNxpOUsQSvJRmr/vWqHlj+P88+iDY1E/5BawryEXxTDEHeZlOwnaQ+KLI
84QqJh9OBtsH7roudmHOnb6fZK/rrZrOZ09SHEEfmiSsYthd+qgPDCNQy6Px
kPH/OycxeqmDgLEKp1V16BijfGT2z3XKcc3EBZgkGrlc/IaXYNCHWlGQs63C
Hi221zyp+gTrZED1ztKquHTnIj5GOpTvVuihoFHnPhVGYPH3zvBQAtlAach7
9/euJ8R0pI6CLaTj8cM4xyH7sZ8B1x/erXcesLXROkFvYaNv7CFUby8zXrVE
7QnnZ9WLOKRZGwBNr+Kq0yvKP7f5yr424QvsePR7yqXUwBEu7rKxw2mqBbVT
7QzQNlzwTyOgQ48GRRyoJ7duCgJmbfkvuTkiCGoNQY9iobsLc0NO4lfoxU0m
SEX/GPN8GNlSnIX7tj9azSQ590/8XtPnInOrmzYzGnSVFZIZTHObmKe0NrRC
XlsygskevQ78ZdOVZupJMHRdNJdrY7Q34AzXN9X2ivor7XCVYIZX+Ad6Ovpa
tMtXcSfK1d9kYpARq6AIUcG+Zcz4Cw9rBxGjwOHFdKzjjOAWaq8+wfKrv3cL
y0TAoSftRT3iYgs7nc7iigV6R8e9SxUGsvxKwll0y3ENULlDyOUQgVJ5vRH7
6cVOJlsQyXGUxChHKKouucx5xTt+UMyE5Zivu0QypRjxQMxKTLtcnygvkXSx
AE1hqEpFoGjNTFpsa6wyqyDxsjQp73it4Do9NCdTz8T2W4KMwYCvK5r1RlbZ
DVGF+SEiEzWoj5llU781tD74aGjMDoCmaPsrb7dblb5j/jUbKiu5U1PIy8uR
y01AQc5PZTZZnQ8YMhpxU9CJ59GUls4ix3rz4uN/eXnXS4k1kbzBiTtHXbJ8
GVArCXeJZZS9RzfSfpAv5Iq5vGAOLKzbJ8ItKhdczJbfNeg2hL9HeHl7e24r
fhKA95hK+ImoFakfFoEDv5wa2x3Enx0UjIPP17CX3KZ7O0vmRq0V3GZzj4EZ
kM9ucTQb5yjh5jVRHan92Clt3aLHBpZtwvxX4IsMsXiIh0MhB+L30iYF9EcM
xXOkYPPpBz6GapFDLdUmH9DpOzm7rBNPdd21Poq38TG0EyBXhx6A10pAviyo
px+dKd93IwxjN1ILCtDCCQuCGacYCmAPnQz+vYo5v36khNWwMducHerzyoh3
wKGstJFFPJRMnDDtleDYSwCS3bfTrrqIHyoLmdqbBLWx9iBOrXbbzySZA4D1
aNobxZVHa5hyDCYX+Iy7BTqpSxjijg0RhOufJCmuylB3ggsfNTWEBrpu1jYo
uvB4Gjl+5fULNUkv6rw6OcbbJ9w9FCR31L1lbOySJBXxOqbRN7N4JbtKT+Ps
vb1keNK5KYM4V5CD8sxe+te8yMaYe2BmrJEq7DtpNQt4cfvDx0SDLv3pk0og
UzDR+JxTircmird9NbNLcR2QE+WsWW2XjurWbx+WCFp54Arwm+UY1UDoYXxE
dPtM9cixkBODed7FiXaqZkIKcYG+3CvQlMBZ+DAleIHuAUUwtbZBqakumXtD
TXjBhoSKvobf5ofzmo3TKYTwL/gHUEZ9Oub4xGcvnf8qJlS2NrQh8QydvALJ
s6IFnKUcqkjpqpQtjVCtIZSPuA2VezM0tq8yq7VyjCLEHtrYPTdbK5B+OBAN
iwPOTeReSdxmYf8YsvaMUJFW2uiJAyoxvBk5qqhVzC++ZJIsBVBiILoKvUG1
1JzRt5ZUHdO0cmrGyoRMc6TZFHsOXAln+UIvmujN4aTBuJJyy6hFzDEa4B+l
MFLwXFnoorMYOUcKf7gWxyCguO2Zes3CoM+JzJWnvhbwHDJT4ukr1MyZSuFb
60STa6SesIhwjU843X05U9H6zRoqp6hDRcW6Oag4Aw0SujI2UbsZrDunkVHw
0Dg0+kBBErC4i/jEMYXLMOhCYAJEF5VV86eu2TngAcw+IezRNzvLJx4FZ3Qo
e4UQdt6BCTjTm1CsyQFTmoaWfB3qWlb9sMHFcG0p6z5WX5uRlc9wZAtCjWO4
rtbgmh0twmg+JsPtNAoy/N6kmXg42L3xDSfbOdSoqYvnT10ojXely3gWOL5w
Q6p3Sg0fe/vDBNXNtFVAWeFCJwUuN/+dqXRbyYwyKMjMNCu2FR0Y48gtu7ik
wlA/PFNtxx6kX4P3ZMQ0jb2PeUr0on3pWt0DTKL3BObgRH+uWOw/b/HmbEks
0lG0yyBWhd5vQu2CrKMUCv0B/Q3sDzJvtCU59BMq9EpUx1dQ69LFtVLLBoX5
Seyz+Og5msBNKmADiBJ8t1A0PaCQvu0A2O4O3qnEQK8Krhq1qhaCzrDFwS2+
Oy5M2ZcS+lB7PnaRFC3625xcaSefIBz6MufdIqna1BNzkGN1zFA4NAKJbi6G
GTYQiKQKOPS3KTtRtNEej9GbgZahco2O3rhOp6TWr9H7doLj+s3yx6cLX7Qm
rmr5SjGtlz3t0p40cZeDs4imexc9+204/bPj60zxF3K1cav0fPI8Ur+rAlaC
sU3T9TpqtS74UV0++8YVO593k1LrLqkZIbb3qKJJYQJi6lZMLvLH3GpjkNut
UD9WLUNxt2BhwmjjvzJCafMmi1p4a17lJuh840Uo1owhOSytRwuESSrdfW6l
oesu5dZxoXabBwtF9H3lfzzW/0VGw/v7yVTA28JaVHvjPfehUlZmwNlKWA3y
6iZJnFm5T1dY50vUIvKyIbiv0AZCRYj1Azq/8sdFTfvbVtdY4fHqjPPp4EYO
NNSb0iyoIN5BVYQ3wiB5ZdeNimq8UZZuXuFERyWv/DwQ9PBaVyheby94ij/d
kRIsJBQ9Fb19o3J7vaOIN+Rf+46bByWbRAktEQADDHonkpSCJX9m+neMOLo+
6S2dieTky2BmVkmm/caXtmEM4pYpZo37kYh/LO+gm5AeF6UO83n8+mRMMrIr
4iSB0CT0srbD9A6NGvlj2XaAjx1YkbdrzoqW9UdVyZcCGZHhXHE2G3i5s/Fl
vChFaUy5X2/pmVQb96G7YduahpgpiCUgECtedbfIx2pOpUWakP0o3GYtbYk4
fxVOi2SoahiHzOkyAwXM5LRM1gYulYf8BKkXGLvrJfhU0jXCJZrq+OUqCFsb
0WblCjHiB64euefP96VzdrFX+70EsIR5LCrhJ+fFRPyz8u58YDVEt8eNDoVe
1uAchifjAT4lWg4URbK9iQG95xVjVxTB9PwFhnzLWbFTn6+d+582QUsuMdUr
GU5yxnWR+pQZPku4INpEBidSQn4WzvlybIr0pf8ENOfVZGGLFDc5mG5OwrlE
mDRRGitVVywpF9EP8imANALnGOJSL8ktuYHbewxIdXRJq5bbwlBcDDisdfHc
7vT2Cbnne3nrFXftHxWiWOCLfLQrvQDhgLSWg/Jabo5xgsR5QAuUkHdI26Ff
Sg4zlV4ypJ8PN8s80R/xoygRdUJXLn/uXdK42Y3GPVXTz5mENp3wqkJZ5DwY
5hp33TkjhsHgbGPNKyyYcBfvE7Eg82hqNcQvcCsJiIKBBwQSRL7FSKmdwUdM
qb1aGk5uKRhuQpITo4bZavagi2GAklxx0aKDVOS/zlI0jpj4/bDAZCT+r7Bl
OBIwm31dLe+Mm9qLvOj6gejyd3DwRY0LZ4Mkh3NXXAd1PJpiUk8P8wL/pNKk
CzwqPVhgS6wiIfOVuu/xBxEW4UQEOJqhDqhgDQ8+BhjpLWD4KLtq3muYmUv+
VV7+ue2uL8zTqXhVU7aBBT0qwiRyHagV5QLD670tqy+Dx10JBQjS/2czChof
E9+56Dfh3uW0zTdE5mypxaE8IonuCADzvUjC6tg1jzhoSdrq0QXz0AIxGe+H
4PZoHMn1KYWMG/CUd0oGmn8OtMym38sku1vIsEihniYWMONbNpbSyBX1qtLb
mTVIp3qYwRPkzELfWGS6qa6yKxomnAhXb/puWNUAMWmD5CqqQpFzn4VAFRVs
VGvipwBOyYERs0E5WORjCy9/J/r3G6udcuyG+02rB8+tWLZxooc5IfkiUYmx
JU/n5WfjOq1xu13lNMeEDVqa7tvSi43+Gh3Hnimg+9bD4dr/SlJCvZcm6x7h
e+vUsBUnUPuWPQizymRepXF/FV3Np3TPaLNuNBhK9x3Wr+IjpBVd8q9uPm6r
ZLFEAE4t0rGPgLWAqXbwVpDEANOEyWKbgqkVBPJ4lHAu46sUUFJgpiLzZcLO
p+D1Il2zP2pfY/fE+lQVR8fe9cuVLJAZZnVywKo9LFRVsnW5NzjmD3wuHScZ
yyMGS2sS/OaVYrAjH71gMOtMNFAqiun6BGuVQE6kVWJFlqMGUiqhxPqdSsSH
TCjWDPCb2I4tjdbHszY/SgSXGZA2Q/YopFMgRU6dfOYBblQ4StJIsG4PdeVz
lvkTGERxwJie71b/rvXuDXqEHdRScBmK/2SCxwIsmKM18oXJLRVSiFSzY0yV
xf3wCessQgSrHX0ZKq3lVxaUKyn15JZF/vY56luSCpRuhsWxI1LoUPW2Cg0W
butCvnIkBr3toa/qNjkU3gppaS/htdvNDHQ6UaMMiQkkPV/x1Mhvk3BzA7xe
uoDSO6HVD903rOmzECEYHkOzxB0Mp/QnPBWvTl0cojq9N/10P1ngQRZm3ZTi
epga6o1A5/ZEspdqURZjQ+YFbotu222h20Qlc9hToMg/c558TENGttycpxm+
+MPlC8ujzsWBHoJEmnXrllPkjSn/bVBMk8fQ5xCW4cFKWjsqBJnQHh/LvFEY
wTFjw1Hg3xIufQi3NtaPzgw/jup/NU5vllrwQw+GkDSfjOwNDthJH0j6zEWx
5CaNAy3of8QH1q595jp8j9y19JbrenQhoq0iaVjNpNrXbhjWUnTqDUiS2C96
zeqG1QcHB4fQnQ7B/MgrylLRNz7Tv7saUCXnPrS3o/xRvBhqz86c5ZYOJNYi
PhbLmI1tZJmoslROyl/yiowbhyZxFe59YEOKSMNREm/pt6ccTuFHCAGvdnOW
stfaPjT68HxhRucaQ6KXdk1N6meBQvnHp5kvwUbU/gxHyw5HSFZRl/0eUIdd
mjGB+u3EGBBWiEcer5hNndMBPdRsjWkxIPIUdGsfxbAppGDNLR50WGSZ0tSI
6fXTvOSnB8pGHOeE80WnOMBSnLgiRDSGOMdC8JDvz2W6VqGp/dbftApX30Fp
YDfvTDblC3mADmSikjYzs/3FZ3Nf0DvlvQUJG2nyc9uhmx8mY7nMRDozyRnz
YEfklAub8JQp6l/mOKR/YcIEY9we4DVWw0635RPk73fI5EV7TpqkBB5akbZi
8qplycC8heTX0lVerX4Ki4rTNeQhSlwVm4wbQ664gH5PIUqG+MKgTfJB0Ui0
9XKJlbLciPxxB78kzhXibrdnK8CrOBUApUVzsWgEsqjNrjJRNGo/wv4bSdmY
Jkhcf+mX/yLFHFeI4a0SBD5ns1mPbyrWW21vEOBlQWHnVJQalJVlY2azk988
i3nJECtg+kPZdkBzT7YPfCNdmJ5kVm4Oil7G15S3tjvdogby+CYYLh3WCIsh
+mG7kz+SMhFNLjI3/SV8rV0b9GQxHFgQznXmDSf3wbXjTMdIpMhcNT4OOQCA
wVfiBAwESOvm8rR68DgVwLoNo6QL9Z6eYtr31JcZ/UUyW7fBZwVLFcxdOAdV
n8c7r8+2LE5DJsiCIWrfkgqeUBgLcXadlJvID+CMUlU+DhTks6ertW8yiP+b
X/JewzySjh7P5eDUtCHSGxbeEUKIl4tYl7zhamOw3xjX/W6XYYpErdRMZkrv
vL9nmmKGuUdqzPQcSoDJNGsn44s6AqKarEKau6r6ZT3+BQTCbE3+jr+L1RWk
ql7u1Zg0WrvHbQrgVIQdiSAo7mkK/yCzQ6jWKANaM0kOohSLWPsYaukbAMLx
wUVJUcP2Ihh1wWcTD/UsigBLsdgVN0vCOkoRYplQHA8tKDKX8pKAn58gTGT/
NKDxmNhaJBexpxU33SMp3jxtf9eZO+4vUt+yeaWS3N9y6XZl9ztPaDwR4wdy
rmRuU7zLCwCf9XOoDsqc+n6xSUK0UpA0pXNROidj/J4UaYmhG5yWvm/5aruw
Ur/AWRqxL+foe0Tw+o+zvLleqHRtkQawcS0lKjrU/wV8ZK9X8knhObImYFsp
4w9maxwxqT+stzpAzW8Q79rvI9AS744zPA/mFlFEIX8Fa9FQEEFp1/6v8FTv
IigYr3XlZPZM8Mx6HXHhOIxIPUM9aHwzl0KFQDypClRaKpTwMd70JXLjDQpo
X/eb3yxzOZjkhFWepjbcQou5U3GLpvTw9dtKrNglFGP8xJ9MB75HKhOFWw22
jHN49aT7Shf4OF/7dtyv2Yqb8H2/LSQJdEaOza6Z79P2BeRPqZ2ZbT5qx2rE
UkVOzMm61yb8KIUFhpdhSAStRQi69N3YA5nVKbdBa/XCf1vleVBs8EIRvfcl
7np35oVbprbgbPKREGXoXy2ir+XFQqKK9zYLCM8Sd3var3CHGYhfHPOQ/suD
4TugoZz4lPw89tsXHnxaoR1dinM18Ph+iA1GOntC+9b3TsWyoE2Z18l24F7D
YD74G9J9EuBOPWQZQg+zd/5XTzt7e3yXFgd8kuBTpyRMx+9HsvnkNxoo2n70
MB+89KrMwevHcKEjTDF8+ytOYw0KXRuB7UsfSZ0I/1wgHjSvijWgWzNjkMFs
FvqP9IvSXU+9DamBix0pryZBTF0iXcg/tF0vjZ1s+1RXW6TTIM/H2qVgo3s/
eqa+Xht+ECrSLxNrjXwx4xUCE+fNd9Z5d1x+URJJPOQr/+YULl+svXSqroH8
s5OFVMbrsctrTkxOSlWPuhxyxHTdTcObqFcwmuQoFs7JtFct7g+bJEi35PDV
AVI8zEfTd7KUpQqEElEttoSXviEAZVu3A7zUjHEJoZp+eEVec21Bb0X2BWDG
mEM78YlRxaJZuSjWcqM79JTLqTYKHgM5XeyD0ovys0G6/Qdhinu3PNJ5uWdI
c8SDiGS4x/ghudGQko3/N0bBUNMHDOm7ouAiaqqEWxvloiPDshBbeBA+uQWw
pZZk/tq4xdSk+lQj2w7r8wN3EOi/QBDcKSxrsXRY1wQwel+9qgUchO2dUkIg
6TL7Nq2/Jz6Yt31sKg9JBftx4HitUhjKBksMmlsYs/x3B0QXk0gOoJjT29mt
Vtd5CQoRGpwCAkDRZq6lbeiqfJzBr9ASXhl7Vrc6OX3B8vSIln+SeXZ6LB9K
5T08ah5UA3gTYp126GoHG9iDKh8FHKi3MrEyj5/XQu+DbU3DGBGPNFHdo6wV
U2xR8d9h99Es5XLxE1L7hWca32axLkVJBQg1GT8ccw+mrOx3q/cndOa/jmO7
BbZb+5n9wx++XcUQlOZxOTpYMvZHOY6ou1dz5MWjD7LRxwgIw/m9lvfWZ4sv
+EZy8i+2QcUzLHNRj5gYV5nx3lsW1wWpg9/sn7tk1UESpeWQv01ZFeBYglse
Z71KaTvQ7uxcdWKDSb7s3GV00zXwGk0phQWYrQos2KzQOqy8jE1QdpXi8pc8
Mvzq0FQYtBPTVUZcIvnGCAZ5ZWqQruyJ7TJKp55F1pX8+5NKRQxoh01tMVPh
mFIO7ucaOGgYzcmJ2/sRp+6jzs5+yx8H9lBID34bBa/steQIYg9Q9nDlMS4t
IyK8gyigrNLS29+UMc4YTuxjFn5g54eRwigKldSFwknZRqYV0LxJ354HB+W/
fZb5ugD9S9t6f6rW5V+jLnZK+PgvW/ThHi35f2r0aqzcGsGVmGBxDbPSh9U0
VJg6ES71cikA1QZ9YAUtdswmtGmQvizQi9mXSSCwePPhDeLG1B4pbx6RBGx9
3gRuZuhoGAOanNYCLMrtZl5vjWhd2lymQjeIZ/k2r37RzFjG4Yf2HL/diY9l
VUWDQNs9Cqnxb46DZVRYN/hc2F0eq/zD9/BWdtMaTsY7sXGtDki7cvD7QI+U
FoogvZKEnDKeQXqU5Ii/FsdauJMdtUHr9VUszo3ijWp2XazAZq6xKmippS4m
D/rpgSFn7khbOlkW0xobFo5UODl32dvTnKPk0eVPFD+cZS11KgM72j1Utk6I
Lg2qJr7QW7pTjgQHCnUVzThxJD0xJ9+g3n97VMrc3YGlz3R3Ld5lBk7deSWm
sLYsLaMRTykodLZ1xmhCbmc/Suo2Uj8qfugOB/UVs4HUjuZ6zA8ktWdtg4C5
N/dSmc6q/YqiC/3hqYo9hioU5yaS+66bqOVvwGqGRI/ZzVLeARMEOAcGrMM/
7b0iMppbh5nKgCPZ58zGcLd9F6XgL1TECxH4DsD2MODkYud3pd7uZ3oTAgNP
mAjze0NVI3CVxC1VgMgYPA/rgWkexmbaRQS/nNN0HdZIYnk80gLSqD8fT2D0
KqSH2P30ck23ZRtS74cxKFJHFIbSxoNEvDqrt/OuuuadzGMKFweeGbKRI+hF
ksr39HSezGQZQXbVknhdWXQwVTmMQKR+vH3EoOmdEmg/UneZv1QhAhuJxVvp
5RDHl8MmIX32v4ei73TUfeeaTklhzQwSam5dDvIOfn4FNDPrvjl8ueaNzUnJ
KfZDzEEJ8Yzh+cGzcv+H/naxoQNYqkmocG07vAoEGaaajOQ8RjuuSszSA5zH
thLfjNP3jotRF/RJa222d0m33KapEsmUG0zN/KxBmDhW75uAQk7Y82NC8nqW
rP3DzNy+3Vi9QfAbYzj63MW6DsGFG9PTWlyEboSzW92sPouoiAyE/BOyxFJE
Ec5nbXZRzdADvfOAe4hFF9uM/0Dqyv2Z7UhvBZWL2YJPIynjDvKqvhmqmNtb
N9FNKyMP2MrGv9HKlRi9S0fzqGunyggYX9yTGQX8OY4MJJtACUdLmNv+BzJ5
TeTNPnLvFiAae7OJqin+ab+NC1xXeUZCPVMCZzjZwpc6tNUYa2Ac5kjel1Ys
Z3XaOUPitbQd6DvhXjtlPLuvaRBiEzJdF3cSkVFFKRsV48z+tfFV5QyKF2xl
AmDK7pC2YKnP91RF+cUVU0cJbVW5gxiBVVQbhixbDNL+Iir79VbTe2o9AmMU
EzJrdgpPjXBcg0LrEwLdHQp+wxE0ZCZyq/wL7eXLpzDwRVW0Iaw48L6W/w49
8LeBz+gbVatF653DBo+ZVaraeexXQnHV7p004nhDFGJHemKrFTRY1rcMoKQF
jPn6Zdvf2XkQ1SSBvKV2Q672bCECMg/6A+2b3axAlGnce3bQZbQa/D5vW+Wo
i1j8SqQyie7pFwnvvyltDNfnnbtluGoN0cMjF9W0RhVF7AsZFIQaHdhl7agK
t5ghaYsbMkLYrRc48OfCRmLtnnKrO7ichHSjILczkwTCd4SloH0sfOHpAgzO
PpVZVvueb0xCiraz+G22bLh6cfzXWkeOatgh0TrJNfortsHxB2ovSCVuFIVR
wn5pti11UtJ2jcA1jeQDEZzvj/SfYjChtLDvuNwc8fYjN4l/tBkQPFeIFQG2
CbCuACKy0CI38rmY1su1ThVLO8Neix0WrrOvaJR/SRTp+Kg3J36KWXDly6NO
56uD4yhXAr1q7NvlMTimOxxBp5M+t1BBs8/yBnFLClLDhCATK2OdHmW/EuRK
lq2enZUoAJSjomUakid6m7TAbblowzouwJt4uREqZY34GMtJ9Mk7MJDoOOaC
XJAk/BbtXC/E3Ln4a4MfwcSk8xRjX4xZC9vgWTPJ5b7Np9Bfd7M2SmEElRUF
/0+qAdsDi8uVw5UllAGHDVetdjUbWkr1hz89VhUq75tTM1C7THDCjOMkJVHu
/vmusgFnjezEFRaXUyxEGLw+H/pWNd0MIO8Z1n4Er6pJNIvr6ZOYdTBFVyIi
3VMnVXGS04J1wVhRkUY9y+iR3ofizPSMNkd/Wcbn4dkvkrqab4I/I13/r3tY
tvMuTFgIAmWxW4f+XJbmN8aRNqW61RwjgPI7f+PvjPZfZ0xnQcmumzLlwpRo
OBvt9Um8i+PzNHK/wJahHh3iMNOxs8OujoiFxQ6gx9++fTSzjfLVkL0uUUIE
bx4wO7ErATVVjtq4QXX/KZSsg+bdG3Qn0tvfJTlLmJfwLwW/yiVbGtr3HiSb
Y+ceb8QMSkSXNLghR1ltvU0tUEWKH2qrEIANFwX2g9sGfaa86bFrQADeCZHL
5Yrq1+EJdUIrd3U+yIfwlPgct7qyVQkvTe0C9SUGb7Ahclk/Mz9JIjgIfKAZ
vG8WsxxFc+JnFUJdqDYjmG5LA6Bxoi9Cay4+1UfHOCbR5qSUbNWcRhilQ4C7
uTeMEAmPp8/B1DytTFKkOt4RtAcZskaA81FR5EgKMJo6zvy4tvu2/Pfpz34m
NkSoXzXBjPlgoAQfE+K3+wgWPD+jwRG1gv0uECxNLAIJXNghki6ernuIngrN
2js87YVg/ZpXcgi23AwV6wZJ66xbGCgAjHnFmeIR1AuJGrt/WXKXEQTyEcBz
CCpWLeKVen1NAxWsxZcCeoAmwKemclppJb8mr3CUODjZv0+RjRoyRJE+XV04
xe3ssQmgiqR+85sIIGUWlbzzmaI3PmKNryI8vP9CyMvchM+fOJUOfTHk9kxE
MWzRCKnfsWqpYtGrITmIWL8sMYJ8SB4ligGPf682bU7OHkg6uZdt+eLlY3Uf
ikZ4M/mas7yjs0lWw4IdqFjqYU0AAKn4objxshd16PyvhZjKPKNbu75IQKia
u2tnWlVnUN9PEz+uWK8xni5KENNW+szyZZ9GbvB2dx1FktH+9BX7v4TR8LfD
OreNVPP2vc3zroJkDxqzRQWcLPzaJ7HHVvpFsJMrKy/th8jsTYVKMOZkhcFu
4ymirlu1A447XnyvjFiwXa+sjNQkyMQj2cmhJ0k3RnBICFmsGRgg6MKvOmFe
nvxRkOs/6GD8hU2w6otWP1/JRdwjRqAIZhNjs7PVfZ5M5XKwKsw/t95d/u+b
o/vvkgkW48fkhX2HHtZ7mf0loC31cEVjjpaN03WiF9oUDiuf+A3rsx3OaKf9
0DRJ8/CbG91yRpuiisOP0c2Xy95IM3B+U5h/wEA48ln59Z5ZitoHdafze9Mo
4ZmcqkeM7qmOnI4ODtMyh8VTLYrfaf4LMEqSTud23CBrgvKv5uc0JxeHpJfw
7ULa14f5GPDJGR6EzTJkgLm4msaw1li7SbzleQCE2UCkfMj+fOOU2nLLvguT
yyBY511b/0bhumb/ktIVkCfpSAbx2ClGdbeVDIZkHoy8x8gIxnkqoiAxNlWC
9EDv9h0eehOuNbTQUjJAcq8s4q2mXMQSxwQtjj7gGGPtNhx5bleeukUjZYcn
U4dLKdDnuoOmIECm0Vm7ZZm1MxLysX+lalcpxm7R0nNYw63kiuuJUrfxWuwH
VLD3T9kwH3/HoSThWSDTwyNxof7vDhipOUFNfDMEYrEvcRwVrDDc+DRWbdAM
otGY9//FhtLdN2PEdJB5zYNa/6oP5SLUW/zJlBpSfORAcpitmN8D+nOLWly6
j39Hilichk7P+bstzmtwyeJIzOXczSgyKA1eNf/+gRuv+e6MqTXmjKHSY2U1
lNP72nbGq3gzrjL1HtPIoga9ghPRZRDGoL7F0jEjK0vQ8+aLpVX/AHbyFgZp
unUtdZlxbxGLWIMmTTkeQc39MCOwwIQIjVbs+1Yu/jCGmAJEiM1I91YkZScG
ywQNEFX3JPWzcP1rD3EgJmXQYq77VGeKz2zyw+9EBf3O89knTsQ42BE3QH6E
h9w5WmT9ALowLK0PfevPn7Lg0xOJb5H6NPNMbDdIQ9PIRllFzRsJ+o4Kgm/1
DE8hVwX1PT+zYkGRR6IIwq6FHdIGAOelvRJbf/LfFZSgxgDfBUGN+QNVfwuU
QkLkC7uJj5t301FR5ZMXxuCiGKnuxeDOUFQytK/mb909od8lO0Quvnt4u3vX
yw5d/yfEff2fXrlqhL6bTvH+G+zdcgbdvP/KiauTrdet/zvZLfYApA8suiol
7LG4525j7OA33QWAjh9SrI7MUg+YRPgZdOg/DwbPK5AbhREZDL9HYy06Muyv
4sXC90bKfYdPhN3LBrZEbWLYry7lJZOLUmqC05T13wlYxOp8VdFJAWZczxu7
tghu14tF9Ota0ekrYfWcLlDovDFDr/dl2rpCuQ34KkCGKW5bkk8Z9YIYe372
JuCHJyNvbnRVUh1pKkLtm2bPXxxGb612tG8CSahYO7xo92zsAYlmlaAF+RSw
QucsNGU4/SA2hEtivNrMHpzUoHi/dij3CAUDUJjw2QKaWuJcVQcVyvPEya5o
ObZn8quN5kKGeoVIdzcHj66+4N3VdtoNvw/duC+5Y0DPsq17Dhc0mpcjsUeS
3tehTUeXn0kjQ57Lx2TmzQmIjnnrV1CNcHq7ACPGVGCIFWKIFicOjJ9Hipdm
OrcpCoUfv5xrFNUeaXkHSmQfabmMBt+4rMOXRFHsEHw4+sgjtOaNaSm9lmRl
JU4SekefR1F6WM4Dc/GxanPJrjSwwTyZ1nwLtUlg6J9+aOzhLdv9Kwm7TVfH
GzLQGQzhqr0v9ywzmRlFpinP45SldGLcC3Bnw/3kDNE7WSL6ZqzAO+ppNcBo
lbdxez2s7J3w6JkOWT//+QMdo5O21z93fghT2xnCG2/KJi2qy2jfiXqC5C7o
SsBtxVoEydUgblGFOBwxZkcRgBlODmrr2AFXUv2CJ8PFZik3UJ6nPdqbnFBS
f4rcYIUYTV/QYEA9CcwUaht4S42fuKSKfIbdquATKTTR+08+mAFmhQ8JwG0v
LJDOwpzZEmWnZHR4CrHbj4RwEQfJWN9/Lbe0DpqU2geXdjcS4K2oNEcwYIJ6
KDNhdZwjWw4t+gEf92jvwu1bzYAm4htc7pVI5ALP1hwCkpNj7xpeHd2F64dl
Pt8DEEX7rd01N+EC8FB7J9OGT4OAdLZQ4j5Hrvvr8Moc7wB0nLxMqX9lcMRR
31A6KMiufr3YmjZ9KKtBqurSB33zy7I+9OJrhhyEsVXEB5WJLKhzn4k7UQgV
fVVK5snXKACUzatj5eptur5HuVzRa7UsjFiHH+4x2xoffT77BK6CNDEPMU9f
N0fbdrXNxg6thQb6y5SXjJRPpHmXu5axUFid4/PQ2FTTBbUzaCr+0fSsGuqy
MdUGV3JywjbveV58g4AnNSfGbsHJjBxBqzJQQarOmyICmGypM2ark+3L9f54
TX1ns49rxskeVAOv6nCTuPL/WRAtpHK3bUa8GKbBF1c6Z7K6DjKpIzGJ36qc
J8CbHxhl0agWmI81T9sMsQoMHUzx0TIkfu9sr1HecL4ImnttAMpbMmLKcshY
BBNGJxCOHz2vRZpMSaZ2X3t/rG0cOyyZ3rV4cZgY/dmmEb7V9P9LyU1EfY7a
zwkWY+ZsQtGnaKMhW+q+Ef9kXfEdYt5wqdMrcSKVIuxKTKHO9m6PQAel82sJ
4slFsY9Zngzppf3QdauN3hc/cPrLQ7OW/veOooVDxWdJVpai6D5eCmc+dOay
g6Qfjbpw/0txNqSSo5ySxFrx0mCfKVQedMMqsYs6zVXKG5v3jYnWtbqLUj2Y
y6ByllcL81AkfoQFFgSuh1dMu+QYsN7EcG97PJPs/zkE/kfZw6SMnfvV8qHf
kJGbrwrCFo6fjmBRh1LIuLqBkUmHlzG0NwFfo6XFkBsEjvoxW1o/X6WqpZA/
5n/rJSwT8tUyLev+Zf6w4bf/JQYbBvuVQuOufHwRHnADommIGRCIPWoehsWC
kKOYdKHbuFoGvydVEukDkGmIHUfJLZ0qYzxfGXrFzFaqbWR0LLOFnjrJqV7t
cgkdWdz1WZg9Xc0hX8u8BjkGY3+iiQzClbFkGRo5LOOf/x+r5xaGkF2m3Dh+
1d3GbTlu+3lSzZgsJ1v3++mWw3h6+PpP8hcqXfoZPbmU33yTlrFJa2g2UsrG
U/HA2CHqAnVIo77akclcPIbmxDuUEfq6BsQxj93fKzT8jFmS/X8gSbWO7N1Z
a9tB5WQpmeJut9qIXSMSTPqjSuI6Sskk92XS6i7/Mgmb9SH9kQXd8CNLDOi6
m6UP6NkrZ1OQngixao4bndv+6Ahv5pAMiBE0Ndy3839nMcrX75RyiE/n8S3x
b7jsUBgobM+sZCBGhhJt8nvErWPV1SRCKObGDxqPJ7+WUyONwDeLLj28vqZE
2j3UsIv7NSiQU3T57Wc4nA7LNww5jdGP05TcYHcYfhfI2zk5VT1DXRCu5JfY
cQsrPdD/4QSAooiz2OnORQ8IWcrBl/VKtJacr8FAcLaoHZtYo9CVpn0mr+SA
qOOWNuWIGw6tnqBFCaMsn2UtH6cAP/R4ZqVxBGDtDj0YX/JDVrqVR5Ruhlv0
z/p7dIi77pU+YOe/N9HQ5fM0jN2EdO5cV31WcEA4sxU8/jpVUVyjCvPpbn/F
QMRhSLBaLo+9YZFignJtUsIRCot44ND7M+zDzB91oBn0t4ZV31FpdmkXBJkX
BLOSHhxm8xKLOxCTTKaUgTL5geXZ1hGWsMaclnrig8vUTsZ/IkH4nI/OvJt2
L5WrNFwGeBG5nhw4kzZKgoY1jiY7xCk6tDnQmZFZmsUzkilJ9BrZ7GT+5gAd
Ki/ZVzq4J8yKfZO+84gO/+J+UKjpxGq46nNSUIM/NTIBlinpCVq2iZ6tgxFH
ddLPP2rilxDF3+Xlmvd7Beuf5ShktTvWxjMOS11fa8j6gboVgOTxbIh7sU3T
7fw9SMQ4ErmPLnHluhIqz8M63WZCs5R1t0k/DXOdLoN5jEgdxxsRZ7uIPtch
Wxqivuky0zo+b27/kwRhp2G8+a/0oDkSAU3gz2ZJodslaKhJot7YByAbZS/L
PMxFObVcMJkgoyjSdu/GkYS5TG4+LTQv8cExNgU4yCcX/a9KmTz7eHmBK+xX
x0WUOUwCrAuq45EJhdMdGG1l+GYznBdF5eaaS72aFk2ZXGJn7gms5KK5cT5Z
5DNvLRq5TbPevxFufwlW5phU0Rx2k+VIQUV3AcPPqZ8gs/P0Oi9KY/rN6iDw
YLe/dVhJAi6UmI0VdL972TaAKm6WLBtJTjAXVBb/ZapWJG83YmJN92UEfN11
2RNejGrULsTX88ehm7AWuPmdzLCEdI/fw6Azp2EyD8nkzuvCeKIYVYi8wlRw
TGBnVZmlqbgOXvdcjFoO1amfCsYvNBJB5AMfKJpYTyKf0svMKgv3FVTHfy9f
APXR2C9xNYRU6+1B2L0deIXgghz9MOdflXk3b6Y2YNfo2zuv1viFAylK2tI0
hbHOL8Cz7/KPZGrwn9bZmIZsZQudGovCXKaJLlRGnU/emC6zYCYsDQqbZIEz
/cGEBvG3mRMz6VfRJHrmqECqdYx8TojDGnQCJolq7zwMPkBVscGgsAhvc3J9
qeQi2IR6wNs+GnqQ/s3hFzSrSyr2AScI4AuB34Kl9C2fpz5n6eb4dxSkRYGT
TzPpKFPnkMpZe15hjulhpo7TGvMlL2F4NhtPFkYNa3YnaCMZ89JbpeNUK6si
rCJk34X3RMY+CNk/VEHa78ijf1FUzwbdCXpH9RUnEWc/ajF7GQNHhzyiXuHz
WOCoqp4UiGuRytyIY4qwUwWjazHTBKqEGTwtik/r5ZS3lkV4WxVjquMtwmqW
hn6Yx1lmxx266XiWO9wqRf/zmkae+VcqMa2i6UlCLiEVgD8bNj+OwdtmIVqR
FHysltBnPYSUu5s5Ai7ei8NzDo7Bwv4P65sB1ChEOqxdELjjAqQZlCO8jkXM
xBH8SHgmLwZQhgE0LkpqP4Ih98CRwiOLlylaclRELLCJ3P8oWZ1eEwklL1fG
WDqmpvDXoFO8NCK+YQMlNyQXMLayOzLJRTmXFQlZbNlhRYqrCQKtMe1Ar2xy
12QPyqTGXErvPPMuQVgBwYUCbnLUh+aAE5MlolrxoiDBcdWb6liMUr80W0ea
Mx9FpWh/V5q4t0ZhY2xcJDqWj54laQuqabWYCCteGmFidhiyjCa6avm659iK
UvNVzOMG97xsTnjT6GG4lhfsyBi3CPADHsyaax9dxVTnGJ3KKi4lE8jhvhXk
7PyG955diRlAUBNyekHCM7+B9nkezoe9Jum46SeCZY7NP4/eAmzKKXOp51QF
qT5n6IsIcSgIJlwSaIR0LHX0dRoUdkd2V0YUoqbNABLHmip27AMzI5jPCU1Q
lSC6esPgkzQvIHYXCpTfXIXsexG8N4LNn/BwI1YEeFutCvaxxC0oy7sZyodU
8oV/4Y78lvgzgJsQyvMFON8GoLe56ILcV2eAGq2YFjPxg15jSJE0hsgqn/lE
7O6cbossLpgiIbYrq6lAmMxu8NyXggn0KVFhNSBq3zX+kZZDa8I4BOrDlBl4
8KOz3yL5oZSYR6QeqSw56fHFkM7K3Lf2C584JzVQ2IkdV82TdKP8G4Ols6cW
FSonmfgYRID8CBCtvD7fkm2u3CxBfQtuWZoSZs8e1O/QXeN6oxpwDpD44p2z
9kGvWnyVtlpUns7mT0863jPav2Ls7lq0Nhtj3AawS1ehielsgncA84gHjVHX
ETY+mnLXpMwxngDjEdfp4brjCmQPylKoTN6W0q1ygpZnMChA/EVcvLiVLQZC
Vj9Rt5zYBAa+jbbBtvUk2/g7ODra3SjSDuBPqch9dgRTnBtkvUjYT+Y/2HaA
rKhtVc5geMHoajt6lOkKEWrFr9ihntlFd2ani3vPVhbPbHRYJ9vSTnPhSRBE
RKO20aLqHF4qTJkdWDBVDX//p1VESmkcswBDHn/9F4rjfoRiWACamqunuQAL
pXAr6egkkk1ZGhbrHC9v2iC9EQ5qsBi1ghR9orbXfL5wsH7RryDedCoetUhk
rM6tr3rVjac/an9ud8ATWa63CxotC5ZC17NUyZvdgbfxi93ApH290RDhHbpk
F1qiD2p08IV/esrjHTy+QSjSezWFkYOhFjfeSZt7wDnboJ6EvnBWVs/c+t9z
/faiiyWJf1vWlxTOhndDYjdtzvpbHSjKNVkuSs28145M5Rh94K6tPRWt0ZYu
GoVhHkfk6ryphP6sHZXIOMhyIRs4jD3WYy7w+w2rXa5V/4N4OxXXsJNV8keJ
117ACAXJ3pT8Rs8XifRH0wvEYysduK+EVbRhz5K7NBSO2lIoA2/JCL60/tD2
M3wKEWlXSgPhqAQonQhn8gZ9mka1hBM/rxF2KdA77D6WBqzRAhcOla1obAkJ
CpaEgljGWqau+vA8hR/iR5lR7qU/RtyldgrSfn8nXhuXg1cD4cFJrMfJ11ET
YDouN+xfb1NAUZk59IS3z2xFYPfcTSftWpa8CBs7lee7q7z3lR1cj4lbGgEB
vzqal3wBOAkmttPFoP3m5KKxcFKUdKenQTsWgzSuFrwS4vkeA184RNM/6g4k
l9auNneFl8bmFTFe79GnabS0MY25raiW7f+S1TqfPCVCMF5l99GC8VYiTgyB
cwowujhqJhMqX1Zgw005Oo/vGQ1XGWMY6uRdfrUeCAYtEa6BzXbW2X8cCIbU
SCObCHJs/m+Nv9M49QAkOqKL/PIVKkFXA2n8u614m9RP8XPALma6tEd/mvCk
rghSnimiIpWIA1RIlz1hQk9Tlnz51A9efcKca89TyIAxXEMryIHKrh0ERhE7
8vll3SM9yXHKsn7IE9VQQ/yXWuEvM0fKhVz+j0WdigW9oV5AJjAPgAAzepN8
XslNz1fsq+xnC80Fk0CfIfrp2Qi2LIGsbnySPeKHHsQ7upbjJ+tgYwWb8n5t
xc4Y+OHmq1d4LRtBUVL26cqN7nL6fZ+iS8zwPZrHYBQwDtxfJs9TQqX5YM8f
UtmgIKcW2P1+wObrtSFGPqj7jAvyUsq7rumCeL+sVielwcGjP5w+uN2KW28I
gjlTVIDFEyZwxkkPT6oyJG9nRUdGSBo7+QiKy/dVVcpxoY4UnNghc3kBMyrC
z4trnT20hhObMWP1QgjRef9qW3MA+YwWLM51jQD9/axVGDRAY1BtVb+CQ0g9
/36dYAblBeXh4pSQ5CGK6ISA3vVtmZ5oPr59B8U5T3spqhF90jxZqaI/HkRP
fRPeUXcGaLPuL5xOf/fl+dPMu14GpsdP8nAfJIcebXVaqIE4lfaEQlyvzuMc
01drBxvZ3NPcoBNhn+XxKkja76RYnTt2MsxMawwTT/fKJ9onZAwOR7SaVQ3G
+Ek/LvTFniUDes9fQS9pF5kHllO3M/sG5iH6aQpgDjUDMbVMIWO6yQEvj5uc
0QSxjuDUjN6lZ73Y4dwT9A+gDKyd/ygWl553xlRbR55f6B2O9ZkUV6JmIrTC
g6BDNomZnD4GqX36B8p/WVsN1vXOLWKauY9Cpu1hxCMlp3cpB54e3V6+hGTV
c1iw+hNHnlO3EcKcmjUKalN78vUONwX+dQ0sGi7Z9dawlAdAITaCDyzx5ge6
iRaPv8MZKTTciZdhLvLSYGKM3AjrpUNOPkoBkyP2HZ1OvhwruOcBR+xjO3Bd
zJpmFjnsGrvCkG0gx+/DtxYPdVnEJDS8gMp4hb22sakht/jCFiqxNEjPc8JD
E7l19aY14kXETyZvwVczQSlD4vjh0pCV58OiRNWM+1dMuvdfKdPngfbjOTg4
HPPalpqero/fuzvjiWTWsvChOhkdJE2EqCyH5klooq0tDcaVQJaGuaok6NVU
9RBV5i11gOjXi6kB/0kgYhVLj48iF4W9ujQbSQthqnByPfnCYrRBh3wxFC9/
tPDtadsn6CptMdbzFcLxyPvYDAlOBIvrJoFrTsxW6kD+85zJJxYl0Zg+xZbR
W8qZPnQJNiZEysQav5F6630cD8QbMQbiXXHd1veOrrF6PrsruTPdka0NGtYD
rqPpuo9sSXd9+ROcF52jbds1yjCtdBsVRNrApss+DkDUiv7IXWc+15Npx0Dl
V5kzORxNRFfyIlZfuoDZ4gq0LSwIsEmoILCMzbzma37BPsV7d4Y1Be4rMMKz
zutsMmKMp6mZOjEjV12qqHD0JLnoK715Gb3oirDqoymQ9PG8E7CJNvXJ6nnw
rfTrZcxx/RHRXwQiFMF12VoSmB3yv3fkwDnHTZ93s6sPrA1dmJZz4dE6cWns
OB4uXT7cAYD+xhOe5geXKjmxdfFcacJcnuxN2JJakzgy1Ic4VHEOe3cmbw5V
0a/zvw3qqB8KCYKnOCjOz8UCRWnXy/rdE66vLxassly9GwUwkzr0rH4UxRVv
oz2abVfcgrtETpt7ImvZ9y6EVl4o/gZPAV5N548K956UmKkt0QA26SS+5qBG
nvXjLDV/6c5om/QlNK/vUstAAOF7+HEDfmkNaCeXZcFae/sCjPxMcXcL/mmN
TNkV0air5l8YAtZHZMPj7OZe3hZyjl2t2bGTbNa5TPWVpeDbrCdxSFsXPfV9
D+unbqf6jjJwUUFOxCsBO5VVJdcz6fnGxlvxnDEofOBeZoOTqjvOtJ7eKC+Q
Bz8CsyL7CA1SIrJPNuyr4y5zD8FFy3CalSua7eyUrJf8uAGLXWbmf75DTp8a
RCgtCWiFjTbN0jifbEMS8SjumRRXhChNY9IfdsNDVjcCxzXzBQakam2eb5Ov
hMLEnORL6KXlqaz3DthTfocgdg1BS3b0tnf9ZmwXFrAWLthWPhPvZViyoCfE
8x1SuTkCPa8ez1DPF6ChEgo/u3ub4zlS6nFZHee9pnO57h3WNMJC8jNZd9H5
vl+pUY2Xcw6h723AJ5PBznYrkli4RV+ZKfczHv6xfOBK39TPwz/FHU1qL8vS
Ugw7brmE/pi95fQkxb5GxrEY3Xc/uDMGWEDTHcZJBxuWQ3ft1JgvD1Owf+8Q
CuqELKw31L1793iEn8KS788ZpLBSvjSy/guuYIgPn3q1Kll8Mvmf9QkVvpga
BJzD7SK5+p+7KFiXwpQfUWkJHaVBGHfZ7GwStt/jMzMTkJUMCCJgdIvuLyqq
XaWrXdj0RSbK9q+9EIP7Wrx4Se0va31jgpmHEo7b9hj6ikwjsSNUYPwp2dve
3L/ClGFMdWGtqupI/d4nRX3b+2H5iEYF/5nEpOrffZWFErLeAz2pZV+T3PcR
t1gMCYn06B+5E8hvbpOLZi63MeCzR3Q/mRkQgQZS3Rm2VJFcZy05m2zWWy3B
5j/2H/PycvRaZ47RX4hvH2F/G267AqCNUs3+nDXeadhZD4HoxUA6z7RLI5UM
XOFLBANP29pnfSEJ05euOq+lwBmdFyG39PVZ5KwJO4IUEc3t7seLG1ckQdHu
M6XFJLNcybg3kCDCIy9deJryAyw/8cEkyCAHyvdgsgapVaNPtgRV/WjBd5yR
vBwsB64zfc4nmtYbAWUD5jaBGkUFyX11br6H0YUXhvLbjMeomyouSqI5Z4KY
anJ3KNHb7ijst1Fc8Eglt4XY7u+r1E9EGBeV+9RG9f2jkxy/CCuL6mGmXM7V
sB6fqF2kitZ1c6lZsDkpn0UhdJapQUXwwSDmigY4WX1HRsvhSG78iuwAYxCi
w5df6oq5E02atwvMwR6HL+J/iMUPzyD0Emy4SCkSs5mD6pgarg7fatE2P23Q
Asq3HP1Oqy8+tN87X05FDy3d5pgZ7Q1vcbKbZ5j8pM8Fmpm6cdEECKPf/ayR
zp2k4zQ35wmCqL3um9yIh+VWzN3XoQs7WGsjcUbQx2rwjiMDJiFcG5OK8sEQ
3ivObGPhPRaE54RwgJfPiQ0Zez8kNNOE9rZMgBcTCNHCvUfCHRLY3kl+Hy8H
SFOSfm9dS7sh69p6fEMnjyp4w2XEHsdzEdLd2v57qD2/wviylRHVEA7/u84X
qmBHJbmFpoKZlcVYhtPo6ubiqmV26g4gEfysUY0TF6H7oRRszTi084QWciCN
5EgdyZFfVqAQkQUJPUbDRruR6lrMeEbCdB9PIghX0P6JV0W0Zd17xVwc0Nyk
g+hRJ2nh704ZsCgttWsxQ02sF+QIe76JplZwkt2pGCg8g2B5uajOb4F7/mrl
9ZVf8qCM9PyGL+PziezFi7SC/g0hUkS+i0CNSMRniBTx0HoWAjP1dW4+utSI
GxPXr+SX4W1TKn0rL5oMds2e2TGyj867mAdwPwghEwVzcvhy84Wpte5qUnlE
usb0lxLurOrlGvLSRxrxhyEq+NC2R6Zdli+JqiOccWBS71GRX72dPJY28yDJ
usezLNwsAnJDN02q50bhslSgAf/p24F/1vUTcw39RHo/Rbz2mjN99v9i7wUN
X7LLJ4fg6VidGVRVsSVuRgFtotXImITXw+fTLJX2DgavTs9B8IBsERs24VAP
9RbIHeLV0NmQ2U9kFNaPmL9iqsrbw5izgdgvomEQJVC4GHiCodOmq/wtdy67
0bSDlsu1ohdK1viE6XC4QvVFb9LLesbsGS6sz3iPrHexHhiC3o4qB1U0vXcR
J4oVtBF3k+kvSR8LCz1+qLQ+cHBs9dXt/PTqioDKIK2dBhkwsEKkyyLsKzQx
vVBCjVjcOYibHEYtOYvQ2tBEh0akA+Gjidxn900SoPy8EdiYN9+3KpFD+9vb
qzm//CPa9mdueAJnXX1BDEl4jURYPpcRRjydb+NXo4laV89tkyhxQh/sBScM
ODegBJbW4jLs7CMCS5b5TJR+FjA1u+7VbGGwiLSPCB5UVnDc0fbiTXywuhUc
61hp81BWwmOpmzUlXSc9KLzcvKaP9OgoNcNgMNC3rtohjFC92Pf3hxfSy3Eh
P7YFwWfopSF9FZUV4m0yWV88ESrzJu3ei5VR1l5dspHRK8ByRfNF4xv6XZNY
UJuJXrZVrh5kFhRGjC/GGShmoe/NY1mxGGemSfH20rcAsVGRPu//Xh3nYvek
1ECAI99SIvhXyVgXucmgL+CWjQ8O29397vXLK3V9Vv3ryEmmCOAkamXJEEaD
Ckycg1e5HmxTIfOEgWF5TzmwqIwZxJZ6kvsmJnnlMExXAqxCjFk0Qf2Yz6S2
4to8Rg+iAmnIsp+SJX8+lUIbVDCf3BSYjO3FRIqIrwv/Xtb8Zq7DS8cI3bpp
GlmAI1m6oBcjRCuDAvTR0nNkUbHSyX4Ax88zhWH2gg+pu8cmqXw+FlT1dxhF
PJLEKTiekTeIoGz7hXGyqdds7Zbkr+6k8fXTqq0uLxE9Pa2Kb42paH4B8SCO
1oi6oheht5aKJYnbzGFe3Fxz6YaRf/zXHA4NnbBDOxfFJZpqjhjXGFzsldwc
l5DUzXA8VDLG1KncLo7PTuP2PkEJzfrUOpDIyWGWLJOSwBWmnu4/diuEMmEe
5CRaL9JQrfBlYsJZ1YiYwWRiawqNQnrfPxPEF88YR0RdRyOvGQZbugiy95rB
/9yumQL/bFwa5qcdOj/NtK81eW82wHdLHfjrpoNIAD+DAD/wJNzA7q/1vv7F
GPt8Cl6Xqlaa78moBrslowdHqHxr/6s5zBBTgTDFhd1R4wQ9xXIhUSZtsLR2
plWKOYzG4mmAPBLKSul6JQ3LtMkoOcDboyoOy3n2Mh+HBGRe75EsjEgdNWdf
Gn8nJCm79q8Ht7N4fnP8rFGAMU3LlTGar7sx5mBV8+kq+ZvIKEeWbwSH6nrd
pP1TDeHRhHLx7ExhqvLvElvH3zWZh2+7qGanZoyX8ojzGwVO3ZoZEpPUogw4
VuNxwJMn4M1d/kC9oKyCSwHJ+9WO3MifgC0vcO/PoIT2D4CMjaSRaiF3XSvq
986Mjvh1tZS4lcCfflq8WBH2/eXvzGNS7Us8ogKCxe8Gx9gsYadaW3vYTtW3
1Phstiefc5NKJYfCsCa+nsI4sbEO+yM3MMR6Fvm1WE7aILwi8iCZmuO+p6aC
uPO11MlWq55MnVgSBw70be8v28Qh/dZbi7IxxNAdptNxyn5b9/XvDWw1Os5c
Abh9ByyzuuzLNg22hsebmmRejHKc3YbBqs3RcJrCNCdO0KV+St8OpVwQ6kmD
6sBULuBey8n5wvaHl9unhZcun/kn0PGVpMj5P/K4380d9xhUtJfhnm5cS/iW
Bs8iuh3r6nIE6J3Ma/VO6vpoG5nJzLN94WB5SKdJkJzJXf3GPGMFMkehn0Dm
xfEcmzH2yxAo/hWfKFabu7DMwPsII+Wq3AZliob4Kv6JiXLdu7Ts5U8jDvqI
xkw30CdorwbKXSig1cJe8VDoLMyma2DUab6WHu84gwXKcijf4zR+W79m6UJV
QEY+LxlOF2YcOM06b2oYj1NPR2tNjmmas3RtygUzDJGDFoT8t72SvPDiePR0
kovmrvTAfkTGgEM01JwIR6U56AhHHajciISRrX7ZrDGJqKmrhG5Z6igElTAZ
h/BEdILA3zYr//sUDqkj6o1TPqqEcbrVSg1btxkgXj5sk3WlvWRkhoi7oXJu
p1RyKBFxrFxdZ4t5FSYRofKa21Su/FvgiiaIm//4rjVFyecijK4g4RP9sSLP
28iyDH9lwemFc5qV7PnejFXojnkUmuR+y1LkKmQJId+vb4bNSOGT7JFcfQhr
91VOCiW3ARSm0UNX10zJWLltfzyXbKFglb+hF7pW788UbiMH9y9NdHxHFK6/
ZlL6Ga5FubCGPkNIIvaO47XlFZftPUXA9sw3DEF7uWE/NHtupSF7+DxOxFiq
Jb31JYNU0wEYvGppEd7gJQCpFfnJXapYlK6pCK7RrNTyaDvAGSPsnUqmVij/
6xUwK2lhhIQi1EGlYSvsTiOZ8XtL4H1v4FtM4RF3pb9sWIpM2nR8y4iYjoi9
42IufOsvg5udyDNwj7eReH0NykHAGXSR8ez9WckmNmzIVNdN1ey8bvEnSBj5
ujMcp91rI+1DWW/LbmlqHeQoCQDdRh8ywzN5slvquLapFVNmqC80xCVciD9b
6tNSNY+pTyu5eyS4ZJ1NFY39zskBDCWVlitVN/oaMJ7zwcrCnQ0pR5EDhwsA
CaDH0DLkR5AP4zO4tSAaFEFf9EsFWWwv1886K8dViifLObE9INCoCW2iu40F
dpglpyxWMGP1alhhDeaeOJgI2co5EqV1RqDUeyVIbjqPpoeiUlcW/P0wZDay
DlwabteWCsEIFNZwpCkGjbq3mzvVybAL5VKAik8O3HccuLD4/ecB9d5ok4F4
K0B3Q/0K8CsImKVPs7D/EbRvVbO1C5kvshv+6kSy09d/HTTe3KRBwuV62vv7
e26iuQ1Q3fjvvuJGui6D56ykwVDyi+q8q+o78HToVn6Hy+tp1v79tXtAAYIG
pF1xBVMCn4x/aDDIdM8m0bOw5KG0jbrj1y4WhDTo8JeMl8vefrNCWdz5e/x1
2kXBz4od/j5PxLYsVgm+hjGuj6yuokbkaY+epxBQGekS/UK/zxm3YdnWrrH7
CuxL159BUpZVNWlwpQJipWHlR14dbUzM+mjentfNppUNCk93C0CeYeNL8GLd
bg0EEljKc9la/xbxmkRlK4Je36h94TjSEdtz3eWJ2E35D/fHrySOvsGTAxzP
pvFKQebne+K0uJphmKSXzMSUfOgAu2QWMntpbRHOZBLQOQ+UuxT8PLND7zWj
w9be8rmPMbXc1Dhz20HFz03EdDsihijsnSz2R8lE1qGEnV/Yv2RmZh1iYbqv
fCD2SePT+rA85u2kVkMddaifdYK10u8h3sQaJgcIEfmcrbaItTS5phL8ZbzQ
ptvIIFbDFmaeLnd8ZRnLe+aZg8ximcopSjlOMyfkK4sCp72W/cd3346ik9RW
TkBqLHnPdW8k9a3aOhHGEcgTB8pW6T///u3ZqlyxBs9Y1PIbIkpKGRuYXlI3
cBUXzNJimaWELuks1I01LSzFfamu5XgE/y4g6520dqWhbt/BmSfnbusTMvXY
VMjcafUuEzfA84tlL4mjWfd2zbPGss60csTgc/9pjSBY70NWxryoQZUQLdn0
6tyCkTQrAVquXnKYg//amtwxSS0F/I7DXFU4TwNVB4HUPd4r/IWEbbILB3Wd
oIU/bsT8GUIqDW2iGLUGopeULo88qvcpl/dV6Q2+NFKZiV+er4K8dVzz91el
GA01PmT3DHXpVPLUrY8y1RlXtE7vqpFLvT5oUYrf+ziN9gngx1t69T4H2pPg
eyYb1oggcieMLSXNLgAwRgK3fBs/EB1P2mKry1MB8XYrOBb+bkeNEVfhpBEg
8qken3EE3PI7/0LyIbYY7GqeJdRRJSfcnOBHP3TBgXfe62dF4Xmv8wIh5bz3
bfdtJZYI0UQkmdY5u2mDs8bpjrdb3k4hv5wL62fj6P1uX0uKJsMFDVb21G9y
/qnHZlHpXryQTBhEo3tVxpvTTQPvZPsJOvXvI6CDfeA/HZ6IB4/xGKkPy45+
RNI2njjkkWhYu3NTTBe1t/1qnaRSHCamG2lTpMGIZgF96MaCPVoTSROSm+Vf
+VwdJ8x0j00epq0lTnhYPx1mF9Yyf+VK96W6h3s90qr5tFGihR4y8E3Rl5V+
XatKe9bDECfrjEoG+PsHQ2jPkV7sdrSwrETgmztHKm7vuBsl6/V8dFUki53a
43SBSte8AwXPcpaFZMeWfnZ3qK8m9nwF31sCqvq7TIzkOOVT6eh2bKVJpH86
dPv09fV4KkpQSORnIWXsVNebZY0qgENsir75lFyzvYfFln7Er3NM2U7pioBE
1+lS13byfD+7fIJ0j/mfxPFh3duWE0HnVOiwJh8kVNi2+BZHvywfMD98oB6R
NhyyXs9Jfn5gHKj/CK1W9faWG6IOdH4nrX579/K3K0DxyVqqrvbFyCFlcGk5
GinIaIplcIy2VJ2h7xmU2yi98aNQf3m8px52on9s9SL5mCF6g78XhM0CYE4L
FZ7+K0gTqobhnvnO31mhnjhHDDL9WyFN+a3p54sHZUbmEXQagNtGdDbodrfj
CLdjKuieOYApx+N8flA+3cgLp1UjvFehYQdcRUJ12yYjY5SRFd0mVYAt0xJg
TRU5bi2bsoIytdo42KL5LBnVdK0SeRMtuES28khKd/B5lGCA5ShTZ9uGyUBp
PQ2lr9ex8YlSwvp4qTfRRa6T/DrhebFvl6W6egmpYTQKhs9vNfRtqDcGKAFp
v5fi/LCc0zN6XYT/kI+qOTDALnXNSiB6p0j5YfuJecILjHYQoU9rKuU96SV5
XGgsLJzOwg/6QZZ+TQND+eZ5FrlN5qPPiE1CvQaVZeOJF0C8/sgyLAWsky5W
gZxUoeP6yZr98X5ygYt3FuKobH6k5+lw/xOJp8Ixtrkp0jXSWlVPMOCkqIzq
OUTZ6RDlyNZGK6rvZk34BkOzaowTggXKKMWZ38b9bSlC5E2KPMsGbewnBBAm
Z4wyVgtZvnfPIZEqqK0yyjmHKmnLpi8wk+vHScLcNwJ9BFXe+oVqZfeOm6gf
LkFEOy36mE17CZcwed/YyyoSXkzLKrobpivHHTOdKmFvE2ai544a4Y03Ti/5
ogdYSbEVJePNVNBHNKfH964/R7v0ImoEcuY7HpMdWSmu708e0G+aMlEHF3i9
JoaFppMNvegPFs48R65MuPLt3/VEIIatkKhfxM2UO6yY8QG3DOcsGVE7hVPZ
+PRhKs/pdBnkSuFuw6eVAVILoN8rAJ7p2gOqj0jQX3ali+lOHl6jxiMRn0nm
/+ygTQAX9Mz7tHVXMqznUaHpkqUWar1BlAEVSG3AbkNhHru173vh5F5wy6EF
TQR+9ehsH8eXl74X/FlTwQ9vgigB/cnNqav9xSzP3oYUm4wH1MkwdUj82vJC
g6d1kAGegvrcQ7qtqdveJBLEjEbNLCcrbxe8Ke8oRLRKimvnMH/atU41pT3L
Jjxip/ds6+U4Aikhnz44JwJvITtYBIvOArb2O47Kq86CSJ54k8NW2h9OMBNJ
xU4AIcgDBsy63ngyChL7fU0on3tZSIsTuHFiHkWJw0iYAqfl3e1Y0b0Y6c6l
ZY20tnE86Dg96M1mXy86KEZlRPXKsSUICCXmtZY9Jh3+dRgNqhIVnurhRGss
2NKxPygUDKpsAmdElb8M9B92EztSRHoM2dRuVSbX0c7qU7dPqB1ske1G+dl4
NQp6co/zMKpMO/Xt9o0B9pVhP2CT6YzvBQb7L0x0CDNcAx+a1D4L4arOMHEp
oirmrXuQvmzguAPOMcCECnfpGNTevQu7VIVVjDTNg/7mVLgK/JxLpdfwvf6X
pKQLoLiBrBz1XLShwsn9cEcdcRzQ7ZQAIRmCp078O770++Tnt+jlNItUkI3I
t2EZdh/SlMpF4m+UwYnbvdQGISzn9AX1cMKPpOpU45Kz5AJoupD93NetK/UE
esLBLQ+vmyBmY66WEGmsSHi4Zad2hG/di7XR0mPmDzTPKdyOtMgnS829FCYu
LpHbXqMtyA21UVs/pIi8ChzK2bDQJm5dSGpjU7zsv3m7gjcXHqDQtgkVPpYY
L8zwJdjnyvdyHrkP90HT6LAAJ087GjqK3RoPiraCYKsAC0ayEobj/ueZvaAE
LwnQnnxGeg37lyEhAyDVcku23c6lzC6wKiN5xAfVIwdb6SoeOWcjDT0VfJvX
HAAOFot1XSkjtsIgmaECwVJ1DojVmLEuidaornyAFe7WBe+bcV8VhWNzFu7Q
NzyE36KZLpCmvsPLN+M8pMoW3y8LLVz2QhWoPZ3sBf3TJrF4O0RCywuiEpdy
AufpFOZHFhRg0FRP70t+O1Qa68eYmJIliByWtL6Mk5UCes5MDOeT+MWPUxSO
taebJmdMcvnD+I8umbyws+WhCgXkCsb7mO3mLszHOZmRHrQf0O06ztH3Lqld
jBRI5IarBIo/Qu8Gxpm15XiBk/K2ry52Lzw1xIPCWopond2bi3FO+MupYfGN
S7H0y3c60GmWM8SUgDLqcHFnvKmt0w633O4pz47eluuoIrCygjdPPRCvBw1L
A5FIvThmtWaPAh+ZbrDQ1QX1QQ1XgNQTgJC5eRBODF/BBxiS+l5/0t/kZ3st
zUy3qSRayPZ0D9pBvrdbV9Ruliy0b4fnBHNXI84+7hakDgwhsmtqaXeW337/
+H5B2t3ESjHmvdVuEWM4BjvAU/5nQcqqUvNpLLBxL+BL5LCNMZ6yHcpJBplN
QXkegm1dzFBZLr0l5MtTbxF/KLr1BXLLEgA6AgRcEgfISs6kGCddUtXeLMjB
OVD86cMxr8HZYvksJtE0wJbFWCR5tEJYFrWSl22YyTI2fCHIbVyOXO/H/Ote
RxlL+Niu4fDBLY2hQwnYu+zyOPv+1BW9WdlDCGnI7G+dJ789OOE6Hjs32eqa
UTIScQhsspkzDDTWTHJmm3JbACDeZEhL4b6dvvBKCgx/ruSNoHBnTnuSxMnE
W9YzVt7h4SEDr2RNUWCjVoQ+jMX1GNuI3QihVok0Q2khpvfeDFZMgOmi1u8n
IWFFmd/vTpE3V41d8AlXZQ22yYndqp2iDx+Vz31r/8/zDodX/kpoe96ltvB9
JzNt2nK1reRh1xYux+IhxQ2LU11/1Je75eDj5Prv5B753jDPIrO39zirx0DY
3dFM2RIfjrsMzv7gEsSS9Y4LfiY3D09175MxGtvbWZCc5JWNu10kqhpN5fLp
oyWDxeIfKJlg0tgMqo2krgAHwNOAZvXRyFNMQnkBxpfIS1v43S06wwzpugvd
GoGawEqWdvnnoApe78Yc4trat4VfTEZWSNK70zaH1m4TObRjR21FT8W34K7Z
UVz+AE2nadKEDtqPZQ5vIeRloIPhUXK8qqi8hBp+x+Dydv8Y4awU/dPUN8uB
V/WxmRjYbXXBDeUrV0eGU6+jJca3QbNyC2UikuOx0MFMWTWkMxR8rRe2tetl
FKPbpvSH+W3W9XVMoB4eWpxk77nEWpgy/XA7denID4RkvCQUUCelhNlcmdMe
Vzw28i9ah/l2behkCAI99SPoH20K1omu84bOcVLec2fedXeKsZJMQUxzQCl1
HjgFBFCgPVeJTfEksDQ9HTYiH9FUS0x6qRs1eMaPFSkTp3taaqEBSjI68+ss
vikdHJBrN6aPMH/R6IO0XnvdOYpyz4D141+rPUptKNPPfm0L1f9jBZ+ECJu2
ObHsIchUesw6/ruVI7UPmYRDW3N36Lfg5guNapedsLRpX6d+ySfZG2MNRWrE
s/c4XnV/FEY36+kxdAWeGQ9i/qF3RN8x3cV7LdsnQ2Hek82Kl40ZpvK1Wlbe
75LuSCrbiKsl7lzHLQvXOTDUnoaidvf+VgdsbH9HihREiZiBC8qGaQrLBE0M
Ss8n/XRfjMiQ+T5rpBTr/cZdDZ69xp6dAzzcTov1YC3mOkAqQjYHzNcDzGsW
2lwhIuBil5bPWeNx2ksXat5R7GPE7CveglbN8TaGU7A9yZbrz3F6Vbl88lu6
xyoO5Xv7YE12CgqtC8e1zgPccYhCDhDF36yQkl8iOppuBpN7OMBQKFom5I/J
uR+93R63Te8oxC73YgQcHEBFFPWEI2omcecV6/hpacE7jFFpBv/89RMYNWeW
f56z9bKl/7q8yBczVnjO03qzpFVshK/9RNfoQHUULyNIWp3GzUaoB65n2WBZ
PypYNzdvtpxYraZXA9kS+7f77n0MTONeqJgGK6uJNflufJDqPwkYZELWFynq
hpup9b+MhNyvufXng64rBAeiZl0gCrmIF7RPxga/0tmjTDdNCNiGOJ/HkiQ0
t7xJbg6Wu/Aa8aJ24KZrjaKCWyEuhe4mUW657WuIQKnkBmOe5Jjiunn8MySX
rZZkRwC0Y1RnGDyBbYTXOY3rKFEo7UI3AaLTLmhwcEgRCEKasks+Xqsp9X5A
7V0wv7UqfsT+37Li7mU3d+gAFRUmaKkN7cRjAzbUGUX6vHQTZo+sMJoDUFv1
1nYII7Tw96TxqonTOSGDBoGVT0A14UeTvUwBiogRYux2ajV9Jzl7e35veTqb
ufU+4aVG99H8vIySrwSD6QV1rIhlPdjdBhDXOI/ZzX2qTMOrZiYU5g2buENI
qEANJCFJCOdTQlI33oKfz/UNsHSzpmoFtg5u3V+gVOA7QtIceNlVdyGKR6lJ
E+POy2sPk4YcNykUGylpa6jJNI/gt0jO8JwLABGxwgDFPq46MKWm23JplwLi
mcay/eTC7zIINW7Zem7mUmBTixXrRGgxHwr4+a6MqsHP4zeL+g6NEPB6lgc9
DjU2QvQo9dgbtDcEPGnAJ8c7DK0PTRE6wbdX3hFrx5oJ40H5ENOgqtYaNMPD
f/INp8JVpHTKf91eFD6I13l56wmy3PTwa0kzi0h4kamHyYOd+FK78nXXbg/O
vdKYgZMxqaSDyN5wMK2GLIP+qSmgZhXYqivLEIwkEQN0FybeDubIiD/DTfz7
N6OuFWqzw4N9a1wemcGqMlk1DaTO0hmsxlNau8rfG46fpuCi2VqjhdtJAUOj
aPqz7hBI07YwVwGFC66vDaJH30AVJcSW7Q3zAeczC+FXWgIjZkOFTwaLx5F6
sb6vAJo82ULoblvuHJengDyy5+AoSrkBDdDIBOZEkMG1OAY9pFlfEqdMVXqG
BX80bG57QjGV+nH/URe2DzmmfNy4Qm6m+8BA69ONltuuuFe2J2rpSR59njWB
QMTLo37VQr4/W4ethjoq1nqQK0aRs+goKJ9eTC+W/4Dxmkw4Zjq1XnUJ/xEj
/TT1kgkVyHn7HD67AAsDrlf7XBf/csjpJBy45eXwRRwR9RBeLFM/xprtF/aG
sPkWNrX1wISB5Pd151npASJ7LSeEVAloPC9yyDHo9OUajj2V22htssXsOJ21
IT1J7GL7G9F51ahN+5aoCHuaoXKBd+ntlZ3lLi+CnVQZT7j90VnOW6nuKHrr
E1eDgwtE/WI2IPkXZxfXmIGalfuCpw7EavGrg3qFxdwYc8LW+U0gLT9JZ0zQ
1OQ4Ojmc25rad+pW7hBhkcUDsa+bD3DnZDj6qHsONOWHbVxNDU/qHFVsIqdi
iPjBCag8d56unpj4jxJ5WvxlQ3XbA6qlytFnHomYwC3vMwCRaF/199RYJKcA
fnTyDcvTeMlIRVgIIEbj9yhusOzVyULnmwOvnxQQNEdbWbtGM5cDuuXybBtJ
vdl/wha+BLzLA7U2g0rvCa2cE3Tr7PJ39GtF9ZrH0SwPxL5e+qRVLtgfkej4
FUYEu2OvVc28akEzhRAExQkMluGrUbqnlHwL0dkfsa0tXYDf1rpHSawDPt4C
9BGpSX5sg/awymwYUQ26d2SPGE7ZchYXpPyMCXB3EpRISfjz5WamxhQfZ3BS
AtnkcDr6m0Y42SieA7rRFaFr8iVtFN9+whsavssgF7BfWtQTm75qwHKRJq59
aQJR2FvCMQDUEEHG99Fywxk5v3x7lsDztPnTw7dWpSbDKbzMfSJ/wJOcVY2d
KQGRoFezUXoBYauaFvh8BzDnCFc4SDM3ArHgAlS8AGV9HALio3r0VLz+m0vs
gDy5XBvKdJA8uyGL1ySLqBQN9PNWozUbrFy7JV/L0BuJ4rNxRzc48b8J/ZpX
uHOG9qal4FS4PQ5Vwl8l8P2+WN1uPIXbLqQj00+VHWRSJbe9+SVTdS02iqxo
zH1fdjKKZuH39pRzmBM7uHqvV2s4jDvGdvh6AyzwCLdt/v3T96Iec5np8F5s
IV4ECjbLg9OWkQ0TYf6zgduQ96RlcpvrY2O+Pzww6iN7b5RPyVN8H2UpxRe6
IbGWi33vhIgA9dt0TOo2Gz1vvLNya7W25bilZrsXp0lDnSNKKvCgfJmhfMGN
V3TNd7RCx/MO+f8lIJJxGSj8T441639tONHvnJf6Bwo0pCMGV9eKOGqVupev
7iT3/ehTymYfkb97t1rUOaSAp+sR8k87B71c/B7jHtr/GeOxhCDLUdyAcHBs
jAiKQ4u4j1uTX9CefiJnfyOo024+L13IsN+85noUQ2DzjgItAhHYtjhVghsB
ztt4/FE9x2MJuUUv0UR1R3AGj06ZzWuElvDk2Ju6wiS2LTaphm+yej0U0E6K
+sJoKPjYtDaoKXOZ5JsFE8Ds1LSbUH+1QyRfMQFYpjKV5U1cUhfMc2pPYWQA
C3b3Bz8JZV0sKiqo0/0x4+KrFCW7sg/ImIET2NLyYGQiHII54BPNCrLULFEq
2rtHYMUHPhr2EpvAf7x2/vaiALbA91WXwUYDPjwmEtNcCTOXpBgs+W0Bx7QK
xykZ+FoFmqheTo2A4q9Y50zAIzKlMam1U1+kuMYYkKOu/el5d1DOjEBUqAFH
I5xxk0y2VsGNbVtu0mFNXXF6o48HIWhj/OANeGHDN9aSWn5KtU2uPxbKIShq
bXduKICJXZ+olbEjDSWaAVdH6ZHYBUO2nI75lQK7n7fuNeUnJOor1G+M3Fsa
NwzA7QTM3cdg6URl+12vSzFWa4auvVtTgiwFXhew8d74W0yhIZpOv9NlrQCD
vrwr1Dsd9DxCVbxyOT6kcsC2cn3N56TBloQVHDM8ZBPq+ZwhftIfI2aj1QvZ
SSjnrKsMnho3TheSOfwxri/O6DJT6VIqHbF5sYv5FEDI1PKjeUh50dORCyby
XABTJMLsWxVEqa51vQ+b+eoblHUeRKqkpZvQdxhwcj3A8fLTYZ9ly1vMqtqi
xvfHJiHKYusDFURcoBevhU2vfQtFgPTQ1Yj1DnJKMcGTma/r3B5EmRXlCoQB
crjMggkHeFdAfXUeT1sAE5p2RdXQ1cBRX8co0mLDDtdT/oR7VgwyhmCN38ee
ZyWMTnqafRJwXNQZly5sIRIHwku47FQlPOD+noTUqV2lKbIZ7vVDZy+PuqkM
LXhYfVqLW9AapuW7ILCcM2/zvcepijEfLIc4uOZYNGA2UfQHcGHFWAhQyd8b
jts4LkRowTNIRi0FZU0Zck24SI58d8S6swqhrBx02YfdDB2u/CgmT5bA5iKh
PiPz0v0vdqPjfb13/vnpy2sPU0nEX1wwhUvCRjY2q7fzCMHWki4XshL478pA
J0ZC5oJTSfnNYc+WBLJwvhsf6CFmW5BsTwLsiVeW41Cwxty1g71L9p/uiSsq
2d6ciWsDF0DduyHPYkBSLuxy3m6YBSsDmatdUxKElG+Jz5bs5qSaNinfSoDd
HYDDmTuxamKhYyknkyu1KMXBcmueewnRePlHk5HvNqyYbtvZ6HYKxeCeYLzr
fj2UB3ZvHa2XT3CVvjrpresP8HXDbPB/C+eNNuaCymBwL1lu0BwTvN7VPKIk
3ms72suVOF3NMgRdu1Nq3dGW0KmhLTyaZzTuTZkJ2MYwSOuYR8Lw/V/mTVJk
3XLVqO1nYpip6hQytbAOAPT3gZ5iFBDdN3zTd0Og0Mzda8QZJsW0eb12Olx9
OOI0rfv2UglCzu9VMMR4+EUzsOkTkSFUS1IfFxgGRRjKcr6xfLBNp7gqAZmy
jGSSQyGwOY7PWwkwyxaenc1/7ai7r2FVN/mTtCw5Oky6dBwGkp05s1dTfWzW
QL+QqszLJOECGN56i8Xnx6iohP41uEwDDlgI6stAywR0TxanJsQXrLZxS3zb
w3RuhfNXVReHpX5bcEkREM2U3B6SRGx30f7dM9J24Obn4HuNO8IsMx1i1GhK
ahDWoEKJoyjaxu6RjduGhuLtHBytSy/QTnXH9BwrzeFnYBIqqTkt/Ih2pXOI
7Xf7tSkG+dUEaJJVWmtXUIMY9q+Stj9Pcti5940gWCEaToOga4zyxcz8IMvz
I+s8AEbTPdsD8gUWOzJx5PTYNNPfqx9e2RUj5+adAr5xyNJ4UXpQue1lmXwG
olCPd/393mWHy+VTPY7b2LQatc/keTJXOwR6lCyViDkw3XmpK7E7++bwjpfY
rXNbJbkRe7J+zs+eI+FLLGvJFLANQ61m9NRrOf1qZBe9I6sMGBu6GNWXQZFu
rruF7d+kQ4DI7aBFLpftSsmUc/DJpXKoR/cKe5960QoaOZGrEiAWiKpCZFLT
yp5G81Tc76nd4PWsVUw3/I4I5GEUgliPMlIbZZ/t4gXJi3fv6AM5RONIxzed
nF+tUAOjAuTjbEquiOZSYgboqndMsAil3dKDZFV93SHZeXuRqoJCSO0/awkM
8jmFwHehGr2O+emS0xi7uTTP7Y0CaAyglj3+wBUh66Ts/FzxRaF4zUrYll4e
1XKdve6ynrBNaTTImqjoFZPz+FfsdkwgUuRha4yKdihs30QObN46aRLJ3NJz
Yn6kuFmOHTeBO7iV1D47y5hZRCOGmvtFpC3fG76JZoMWlqL7BYe8F8Be872D
WaWfvo+0LqrSQ5QzHDnIj8pnlK3lnr3JbsIzG7fF7jlws9UJoWAK+PXurt+v
G2z57wmm0Bqv/KLdD81GCmv8tgbN08ADi+4i02FJ7RLz+TK1Zj9KEbnL9G3I
ZvUQTepaaza8u48H0KNfWUYCRvwk/hFMGi80mhaD8Oj+VsVzgUh1h/2WT8uP
So/oR86wFLYrYIzYlZXmsdblJT9pffXZeY0ped4++sOOrabyMnvzFhq2q5uW
QKhhmsaEkleyHuLMIiNeV2FeiFW7ZWSjzhS9AwimMRHefXDwh6RrMRw2hjCI
LxC083LcL2bA4XteIANPlssThltDBcy0PDwEScTGdYJyTyJtHzEzT34Jctro
J8iQp7Zqhjq5aQi+HRktdIAyFBGU/dem5TZlDUM38K1HFrUkJ6KAgnVdxkKa
P0HYheqRrQWJai3v+pr04bAVLZnOgIKJnwCaLple2t7hsbQ4EBts02SHtehE
SHOs0HJvn5c/E0//QCbJHxdqbcA8VnLLOZCXsY7ZMqDGfC5q2YHhWNVMZ4NL
TD4vUfFzi2jGxAjyj/EQDFjTb9zP5NcGWWFmee4rMqCDqmgaKiFl2xb6O29m
Gb2H3Q69+eh9G9kqyDMn5xE2SKlSlwveqpwY2/WobipCLA+6yFL/SLlPhOKg
K6H3WikOHbCnRdlHY9vhcYjFxgSZ4mXLcU980OOnjgYrT2Gc+d2oYW8XE60p
hbT1tO4KTBW8sdSHkkUL6WFtiX5Ihlr2rVuVq+EfCUW4JjpLIWxCcrwHe54a
Vgc0fYfSv4wkOGSnrgS176MIJm+J1KX8UajSQAnFL4f+SkGYW6eRpWJVHZAI
3xLY1VSuSHmOqzoqtBeMWZXm89L8u9biWxoP/4olv0dg0h9Z1liPBQXiLOPb
tnBnagJ1ZmsgPwMwVUzyTa4Vj2Hn/fO9HCXxdgLohGq4HGaH21wG37dXZ2km
oJ3+FMVNZOwFINaw8LwgShtyHLK1ZDSEXfNse2dwFssGrCByKNHhFLTcmozO
Z1vL41nrtTT5d3CeRjrVW8gLY8U8P/d4O/dwUDGP5jQj6ckjMa/CrUSQRS91
JtFS3BqFW5yfaRAKfQZMwqpJCoWzP4ffeWnENe9nuXx/mnr4HshJOU3Yk6l9
VV3Gt/nucKBucu7icPxn/nbIftGNiEUAfny1AAZE6SnVRv47aR2Lf1ZTcAxu
MXkl5UyjJPWRvlxjDsIhHJM/DPKgmT60FKnrotTou4t/nmKPnXVNRPX+nYbJ
ht9TgRemLVkvYYwl7pGVGM6n4GWvYsaRb91PPMWTtA3GQduLbyoK0i/1IeQs
LQJutOk/7P/y2CSfI9YkWPs6V9Fgl7VZQoQz2OEk3QlEh70OPV8Jm8xjV4a8
7ai7GZBNGITMJUGzIf4yMGFBRWi5eSU73S5G+8ZTaV1UtHh4ZHwC7cKcFzHY
pdTy6ISWpxVZdhKmhToy3n7O4/U1bXCefQ0FVxl/bJnZiw0hW9mWzUwMlZ58
XEElvKHjQszphE72J8apKquDIQk4CrRDmGk3rf3dO9a6BcapKNFuXQtu7pR4
7ml8df7m4kqeVV79dhQxYbP4F/xLN6MrnQa7YQ0AwNTgYkFe4kom9moYFlNu
YGBBprDba8GiDK276G2VgUQgGFxJWRZma48difof/lDbebWgWns+mTBCqT0R
QLLg9ST63HcwfzvgTfZeadvA6hjhBx2jaUM3CC3ITe0zYAdzt+3banmwMsvt
j6ZNrmUBf75z9ESJq0hYIV5zpliLwXznRj6Ew2HvL18ngZNqgWwq0RhPLJ4J
33EH+5nLUPPTzX7t3dHVg6vChv2EVIgAjkJrC/d4T4V1PiwdvYtWa7fZCl6E
qIbB8Y33MBc/hvP+QmkbGPqPhW431q2yJbDDxim/jz1ayr5C7xrE4wUyKCp5
RngQb9mdXRdWZbnSJyLkLac1UROaMqqgQ4uPUJ2H8h7k/dZi/qk/53S3MrXJ
FgTlZQranLRMheYA5nFezFgtiEciI1oVZ+pGnZZmwxeMBvw/4JZ0W/fFFY9B
RAqaXmbXu0xFG1Jmou8yAIwR58Q9bnkWLdNlSRgNS84B+E5RZKOe6Rqouk8o
Ni4z+pD7KFnzyzfwtMFEvznnrmiiq8clzti/ad/EoljYK6943Rxg2giWL5vU
N8d3Q9o3adIU+TauF4DivL+xB2crk8Lf1l2xn05pF7K0OC6yuDn1aZJde5V0
js4FbuFd2qW1Ca0JichA3nX9Nw8tA7tvPOyuL8lbfoNQKiI5Cp5A6iLt4y7K
4wqfu6yyVwVtVmUAFjRT7LvlIjwqvDdquc5Za9tb8FKCm9n/NZ+rki0BdLns
TnsyWOjCrvZTyoSQYulzMFPsrFyptiYA3K2AXtvdG33zgpfZcNno7W2M/pY8
TQhbJtPFbg+nrfeuxkom8qB3rg1GPW+EDWihs27vT3bW89fkOD//5l4PIDN8
RJQwZJeW+XHwhxQ/gggwdT8amMPsGBASVOHekL5xTARNiHtWsD0yBiBKviSU
HS36o4aIO0J9PcBk8bjM/thPS3PfKL0Fzr8wGdSXo1BzIXP+afHETzBQqh6m
y9AqGYbJX7ctGnCZyuRqJRCGdWfO4WfUVrdrTd0QU804hCeh8uOOJizcFu3L
wuHpqs2yQA0uxYySeDSmSLAgBtfAAgWzgeoTdZWHKM1YI0iZoYuKJUaPX/az
WxS8mKJJ9ZF6uAua3jGgKLqXdkqTWs/Cr9GMjaIMvO4sFVdax0YSGmHucZvR
7eOdnXTnoX/vgDiJCgkB0gOPl4pLK4gSLxYZwY6saPjT4h9PjkL03PjuvH4h
cmo2BBMSydVTqGsm5I2Y93s1vHRKxcQ7zdUbas2/lIx7Su2EKqbQAeZ8cFva
qj8hJosFJPgtvc1mJt0BQPV8QEbgWP4esdEPdCPP7lbD33pXtbXOCo9z7l7M
mrgyecxZmJ9vRkDC9F0vQdiIZ6DO/FOy3TcGJkC5+2knztDe/FRMAG+Fgwec
qk92NbZ4BlcW6DhQLgNq/MT8m9USbeFpBzKg4RN8oNH9ATqLE/C16SU+oREr
SNNC9AY1y3YJ19/C39QNCEeb+iavFIeLenbUWe1k1CqHuyWPl2w2q5XofufU
heCsEElf8Ju4MGDEoYOBVqe0u/IVjWvwBasvL+ZFmhd83bxtJRNjRpp5pGKC
QoTq2wZ0fJJwhIcsWVMD90h58o9U1Nbzicm6i2lIhJPRFqmjDYm03Y5jQGgJ
j+2LhNLvIL4hkcdPS/iHQ5cqHchv1GUhi2XXSUIEJ0akDciyiZ59aL86caXF
oc6cQHRDpwbRyoYsKL+eXpdw/nvpH0F9Qj+AYk99NrSCd7rU8eou+AjJef9C
e57sXDp37N3CwrY9o0gQGzJwhcQg/q4MFd5XDi5e4JCuSPYieyDFBXb13ku/
wfYM4x4ZMoDYbYkU48iO25R5AFAH7b84nR8x+knPtz/wSztWSjpIF7G67njg
e+g1kEAqYW8wRgeKvYvg3iuNfQwH4w3fVTpCc/O8pCi0l/icPqXLGtz+/WFF
reLcXgmMPrjRjZ7z5W449fgd1403SGeJjYMAp5V2X/w1u/t5Wg6+/3Kh+mD7
Drhj2ZCDMdkBjgk9mvEQrRpofw0EtzeHHK+zej7fac2Fna/fzDnIrUretCMX
x/ADl3IiYoYTPwfdt/k4upQzaJ3BJfpPRlZ5453bP0mR3k84iZzi7fAxYQ50
Wi4WJ3pBpuZqw6/mZ1FCh6tbdhf4F7PVpSj9GZ/WDMcZkJObGFZMoBMStHV/
4xEyRtoGe+1ScPVElbCYRIQrd8Ix651ZcJLsKHmzMo/QRp4Eq7dgWKEnFHLg
aUXaBltyrvNKFFs1OxntR77EYXJCbQ69kvjvUvK32CyNqUubSUg5eHwmwU7h
Q5bA7a7wv1p3VXacNFE9nbohcMszsPn3fwehD/RgHFuFku+PFmjk5E9UiQxW
zG5zWcSDCQ/re4/D6wMYTTkPolHa7S74SkzZRQbCEklRO3yOx8msepkHXM6A
9KR5oRoz+LgQ99IkMm3sBHLTjrz1xTucSjM1V9vRdMUBGcNbu1nMXqfA7NWU
QAGX3P7Gr8Q9deoazS9rkJnJKOoFylgiDsWG7VS8xOai0auca1DYC3fgCf5y
QigUAsJRxGZ24s1BAx8pf51HCG30rpejxtxedwgxe1WcIzxGpQivllVE0DXM
KcExT10e51MIjyhLeOfvP1cVug1hPONWcw9IL4hcA3c2Si/Q2WeR2dglAkEC
Xzi73ryVGB7CpUN/oWEwilPMMhtXJluA1km40oMtPqGjFwumMivFYgTEBhGC
9UY203znTXFgjfdyraNgzSMEHvY1XxXn11iLmaEd8h7WuDGWb+vhMKf53TwQ
cqUfMYPfJ6iFcWryhvytKXv6YfSkK81Lla3Pnu7LJ8l7a1YtKvk9NJu/cr3+
SbnkNWMXxfnfh1EXk+NdWyYkVz8NSgHOHn7xFntZhs48VxKYXioZdGYuwncw
u1mn5YXhL6uRRUqU11xbvMOyVgdtMlrqqq33k3YSlkoaT3E0ORXYSEzqHyyd
GAkTm0OzSbbw64UxSX0emdCE7dAl2rm+IiTPhQkxGvtgEVq5OuzbdTAtee+b
3r2QQ9QxXSY1F/w9+5OeCrR8JYwuw05v97PRqCuc66G4eF5gFqdBUhcNi85q
rOWWY3kmDh9NDATnA8+sCU4ifixXZZv2N2HkMnDSFx9f7oZH8Ran9WznCiJA
1HxEpEXPcw+V8RuwVesuISx9G4STdw4/VsTesGCWxL2HzCYIxSbl9lxG6lGO
GvGFFqCRZTRC2eGYyQ6sxWBSBvx1emhJBo9NjChb1AIO62kHP+VgwilVr29T
Pr1T6GzuK9iDuGdCe7xhfQThL5xppdECmiTemNDvUOnEVG5My19NZlD+vyEq
0KLcXax5cSn7sz5zXZMdykgP2BJM4zKMp+JyEn0NjE9lwl2MpA1fGxB/UT2a
GDG5WQNdXz7u0isMTCjh2iffqjQ8CNQWsb2LE1dMRJHt39xMxF91lkjLWIud
hNhDVlxF2jD1a2TMvjrRr4cuFy1jj5CUIgQhl5wI0eAJpKjgRpv9kRkZp3SN
jBN17PBl2YSfBH0N+4PIO0xT6YhfdUenV4WJtWtOdTt6xETE4qWzagpT+KMp
eoTmX+2Pkct7JXAky02PbFjatUqztvkVgHdSPqp1XST+orMfXndEdTeWmeYX
fWLqwWTUZmqMz7+FJmCWZ+fvnwYbRmBsBnT3C4RrODJ0sZoSKC3PpQ3ZAxK3
3Pdf/s4xJx3Gkkc6/I5ZaYzvMBZkTBpnXIq/MFxzpVCc11osHF/WBd6pp0DE
XgFQM4wZdlT/O2FYkDOH5ktH3N0FiTe/M0J4X3TgyJZvFkIWHAe0x4Cgyzrc
xdym0oDbcH88RC/IV8SYEQr1FC9AMByWqlWpXcn5hDmuULTpL484cqMuM6Y7
xJO0kPReLPpsvKQbuJuIgNv3segpok3wrzH05UfWabV/eBOk1xJPnOIP+/9z
NWJb0k6bWIsetUKH8enjyubsKslOw1A7KlCwarTyWuoCBP+OYtNfMsLoGKBp
tx4Em0fRVOteT3K91Za62YqOKxOTr+ZeMUNuM6FjEXofWcZZ1151A5r95RHc
A22nQ9TL39kMfwoYZxZ9PPY+jha8jlnSS/9QMY0YOFy1Mmvh+z+kGCtCjlGy
KINSNN/dmHSpul4IJbrHfr6tXujeTAJsOq9MdbyY1EBS1lc+pfWoSbyfdHKq
Olr2btHK7MFuKwMcXAa6FT78N57vAQiI3AjidMT0a/GTJtzld9w8WDa9mge1
t/MUa2NIPw7yIUtEWWdjSmIjMISTDgj+Pk3AjTwNvXVGDrLbheBE7Omndjfy
An/bkUqvuWYl8/Y4BAQ1uApHHp9KjMh3g7HehAnuqO2qZWoASr6Hwtuu4/KN
CxCKcLoVRYok6IAgsZws3ph5x33Om37o4BhEbeIM37lWLne6hT33w5T8ZfH+
3n2BNyfkaOv1lbdRkIIO+Gb6NVS+0h0p38CfpRZFZaS1oz+cP+E87QkbAD2V
cfpTKhJpBKh01gFGC3NkrZ4QHBp1Cfv7pgxf/w+REZm4maN0giZdEWpOdru+
ACYJpgrPf7RWEgQNZFy/Ve5cP7It0xcvgASQl6Vt53Sm9fK6hsJmgCoMI1ab
/BfkqDRsxopw8jKmEurP6mF68PAQtqNXdHkeKLipAiF8+yVKc46sIGs+M8W6
gVfHJ4bwl3GWV5wZoh8BQ2NXSJJfaA+3E5iitzEuX7yxnI5uwxuVTVJydbru
Nm6k0hYo62eAogcgi/SyKBPOOwH0xTQaFcK761TVue2GMiGIMan1W7Lsikze
eETv1eVdUkq99CUzAGJlpPrNttHN0LI6G29inKI52vTu+pm0sEJI8ukx+Aw6
ujCV4L4sgyayl5hoASj8Lzsyqpymz3Uog7IrSFdgrsd6/K71QmgwYIW7p/2g
S8LzUDSGcNDF2q8Q7b0r3kgU9v9lQz7UVxl2jpY41iysJ8nkx3aKM/oS6FyK
P7WuglJN7EuS+wlNbHJ5EBXMxoh2igu7bXRGjAlubw0yr2xL62rnr/UmQMZs
tEynUy7kJvEohnMubrCQhwm72o0+TGgCXDK/6hf4eyFUF1eSdDz431hVOa2o
RibknlJu0535+99ljPywOIXnPfp3QghbeZWU5Mcatb5cD8wxpZQgrZMBpzmq
bqRJ6ip7IMHbtOajG+fmaAduV8nY3DPZw6xwYAmhPpG2hjKTUExKHsCBVtop
z9vzQo8kZBA256ph7zYeLld6W06Ut3ACMNlSuFK597nPwc9u49scUYIc5tGv
9MDa12PfQjQtemDLPF3PXguVs6txUrtm/m2A/v9p/DZKfg8AECFOD96nogbg
E5Ptk7zr0z8/cmV/1mvhDj+XqfYDxUFB63gUVRU7YhXVXy8kWFGLHX3t+q/i
M1+3a/Mvt0sQ97LZZzE7HVygdR0zpKWLq306hn8mkPOD50k62Co1KZZzA9s4
aj5nqIYFhmqHByOf/IUldWAoFdXv1nMmLSslLrCnOtyT+yz3oEMt4ufE95ni
yek0AiGYRB06YC1sMkRNIdTCjtDvFlNjbf3FCwg/UnIkOpGEXNtWRmUHhAjq
vIupToDiWEMStuODWA0ifU1MxUDjnolDnOICZmbEPWpxzNE8AdqsSYwNSIsz
/DMzH94SVMZoNFnQQaSI4muU7qTmjg0aK2yVczgPQWuv1hQKD+ilJh5jGAvi
u7xFzi/0sQjesbcPtpfYyCiehXTyPo7WYjHSu2P9qFjAn42mEM6IKCk7h0ak
GCFAThR72b4ARVQH2l8mJ0A87n9/HdWpmFbbOljA/Lph5Yrbwy8cpKzSiB+0
Z9gXxxCDeNM1lq55V4vSzoNP/tBwVXFVXo2WAuRSIGOlKeT5S4kEiz7bvASq
9boyra9ctz6kFe7VtqI3SbTM2DuWUV7+tVUVGR+7TxxU1Eq5Wnw8HVmKugZ9
0bIJCAVb1mSSspsW/4vHv3zwYn3cCCP/mVQG3vvBi37UTm4gCj7BMa6Rf9Se
TjAkwrBggCZaT2V8h4pXPW8NPzDb5/Uf4bjTBMmSEzLvxwzKss2THcG33TQR
Cij46aNwssg/pC58NCTfdLzWJVHkXomKre0fd16UWJ4ADFwdGdF38zedrQjO
IOaiUZyVzhU4cAvFPYEyyF/ygKt4Ije64fMQM+YGx/gxyw4vRY37cl7u8P4z
U9Zfc6nhlD8olVkUKN+YjCcr05WQcC37HNw2jmkaARW2iARnREl+1ZZ1dvqt
AWtM9wQk9n3a2fANVaw2hBUz2QS3wmi2Ssv33+IkLMv4fDtAwRzOMzEA3QQ7
/eNIHEiEOy3rOOhn4dh50/+r+lnYOlxsLmlxhFZ5jOHCuQY9MqKH6MT3mc8G
ieTnVKaLDyXOocNd6CxEPHE8vo9Bl6XNIuhWI4qGBJ6xvrESzban+Xl6H6i9
HmI5Zg9Nj0qJ4VNQpWdRjTReBrpjhYMYMNuyzDs/DNb8n8XFg16GZVCuOY4w
vwdrG8TzoB2t4cpUs6NM5q35MKREAMOQD3ml/0lwwc9XlW9r5AGa23axSR5E
Ne/p2sE0hHGZsNGZH6E9UNVFbZCfTtAv/mr8NXRBasl/Pzq5UVKAq9ojnc1n
oGVQcFBag6N0dhih9ojqgvUOO7pZNKpjoa4WKdt+KUNIh1BhH8oTmzh8cT7U
l8X8UUeKYRWTq/kAmg7tiDa+OJ0CKb1Vmo7NL8r3DKYD3Q98Y8zU0clNOhLx
7B32urmPwYWfd8PFkJB2A9FBGWdZsLD62ifa0/NYDd6UbQksXM+kvwHhtCvw
W9CJq/RO+WOSLhF8RM2RGlo9ZHD4goDfKEr3bDi53a1asxsxKbouZHw+waYB
/WBXIdKkEMKFAVpNIrF5CBgEHi+not70KA2Od/8mvSHnIjrD5dUKF8Wrpjfq
nywT04mm2e0HZqBA/HTLe/VL6WmJspDFZGHOvhhvv/s4IL1LjQpX7uDGvxsH
tOmLRBfVkNTt8Jkv09iPrvWAUf9jvrB5mcdpuL9GcVkrN1pK3xHhStY4eIVv
C5rdQx3f7LIV8SOs+6er6pmgwatJlwPvxzFW+JRxJ6/2HlEeHyxupDAJqaIG
5EB9OMlHiJJaUZWZNikk+58bA2bhrnxWjcrQSrAw9DBTbduWfQZFQKgofFWC
7N3u/8EdhFzIKGaXMlk4XSN3crI+CD4TooqHhBMB4rA3R1U/rUCYCJ550zP1
aMEZ5i1kDnrUXlfyQ6x8UPyOlUstc4HvYfY+6M2x6g4OGHNLRAn6OzXfn3n/
6eEYwcGPA0GnkRgzg0kZ7YLcPnbN2XIEZRpRIAc20Tskt+O1MZWiPq4uom1V
h/JjXxJrm9Xr5ba6sOZePqqmeO6IlXsWICGqZh8OSB/8higB369VO+rfsc7C
QnSvL3oRnsd0tzWpumdokRSrhx1+PopVWj/4u/ECid3gGmWxY0iSRJ+khA6E
ZK7EuXGC7khmacYX4Cp7/UBfB3Ezecp2i6nRUDNN03EOG8C+cp1WyA09Co7u
r4Wytd/c8yo6EuVEKxaAOAkDdkypyQWPZ8BwaPRQ63RxLL/oIp9pW1gaMbfF
FHWo6iBP/D+mcTt6a7pIb4jQ9SvWhmRWHlcxdDgNDPrPKYIOevK5jYPOpf7v
Myso/Lio6xuJIzZaXaU72nNmaDX35BLON3uehcLtvsmZ7S5nbS56RWIjZ55q
o8D+UaVM/Nj0AvugzoThvHpbZkVeoo3NxRxaVNg7SAQUr2OyKwWfEyJaIQ6G
XmJzaxGJ5zGWZH8Z6hW2hhmiR5oTmr1lNAloG1Ig+Tp9UU4a094WnISrMvi1
cPvq5zvgXsMPAXVRCSDfn3Z+O6nPZgfLjqSz8jaHOb7w7pFDvlX9RHZqEilC
7usBt+VWq9Tmb1cSLC2r90yd67LsKaPHgwV3q1flzQzeaRInFOTEPzLsBp+N
2O0mRX9ECW/5LrpDcEpKTGGmA0fYdhuVXpgR+g96cpflgtOn4u8n25DSYNmD
MeqOxJ/v4FonMju22/xvJCAER/jZyI/7ZP5fA0Au1pFocDss/ZfFaUvDuhYY
aJHAJvB+3K3awXnAmusKLRg79WXqO5H+vYTqp6eLUs+Ov8lEj2qjzqScRJFR
Qv3sfispeByiBGksFeqFaWwtSgXLhkBOWUG5XjA1qL5jAOASQ4pg2Co4AcEf
p+DuLrkWsQzUtOvWsONdsXDhMnxkP2qUtJjTT2SmcYXTGPaRtFc2VfSaNWFU
sA2MoYqJAJi0S6lPZqAGv8ssDy2NImAwGwmyvut0frtBf8TDK+3TWGq9bhYW
vNeUQ0vL+elmOvUh1h1/n+4jb5FuFP5YvkJxEa456enlIBtr1a2v1F1Q8SgW
aotpvjESerGJWdmD4VT0SVbx+MpwhrZ6S6wqBme73QjkP6HViIqXwE9QZD2d
nJddz2MSTGriq9yXfVXweRNR9NL9fRBzQSlDA8z7/U1erG/Hp1gji/ce5lES
B+GuqjmYRbCgPIxyYiI8QQSiluNcwrK8PT6w9A9Dh7h1Jxk3Pfe/DQKlg12V
ZtjAy2gY96CAL3DXCP1nZyVANW4dQqI56T6+SiGHgybAADyOJMWhXa8yHA+t
YBRM4skzq8PBzc8dC6JdvWh+fjs1O9AXp7kbjEod5bkKfg3dV2tfxwsVTyJT
8nkBIvjgFLNyRF+AD+OsTR5KQ2y5WD5pwNhYmOVE5FREP0T5brNo55BSiW/M
+dQ0TluAihSbt4ufWiDDkh6ToluvEl9oI4RdMf4ZcQSHsyXTugh+0T0Lqt8r
J7mmfgNfRxkhBdc7hsdLoNXFLHJdLNQCOybnvmY7SizMVB5KrgENUNbHGUF/
XUYIMmU3XCHS4tsGs/UHBMoZ/Yh9g73XPtc7rpG80zbxeclq+fVOv8e5R07h
7iaG9aNG9bk5GvCYlJKsSZlNfIFzq9PglOHY3vqwoJQ8iewwHzTgh9hwkDiY
rHy2RlOa6qGWQAIlrUilSvSlaQi6WeI4hmA+OGV4tFtowQtl1THm6O7vTqr0
ufkwBL3wFl7T+5wuabCJhJiafYLpo1coKL6L0ebb1VVuuhvN6e8YqNPlxr83
3/ERUz4axbdOPIykhCkz4BIOp3xsi9DqX3hie8k9vg52IY58i1KMneBhvyhN
jAfsLYYYtM9e6lFAzYbbxIeQkQhd+SuqyjwGU/BtBI8y0sOiuGWoDPxP+XGI
hG8p6/9Mw5XZyz5MTVE6ceGPrrlTY9JMG5IDCLjNyoDZaF8Xqic+L8Dhjxqe
sMO/eGZWNN48kMlqLdyO7pFDDHW/2MqioQWS6Xq+12QCIjq4NFfUlULoOwzT
SWm/vlOilWVkGAqmcetlxhOG5v2Oks9bmZ2pImlHcw34V8jD+8j9bb5N7wZ9
JIPxISvqFEsMK0LshwvIVH+byEpgaW1Nthf/d0jquhdSGbSNGLToKYsHf7QE
J7hvEp9g/CG7vqLBVufX/64bs2i3ckHJopo5ptkjDq+I+iwZ0PZUCS75LEqM
5I8NRNzNDoGtoPiUvyhJ6IanelZyZgnk+EkNAjZggWtzyePttd6kalHjRZd3
tcTQE/1/NK9CgX39YBotU8L2hVs5hZwUCiTwVODhFk1n4sVH0EJdqljs0i6b
s3y3DgiBewi+D8+FPW9crbNBE0ozIjQH6Q9ODTJg7q86yxEeKlLsxPOWAyi5
M+SWE5hdQjWixXLhqf3GGSr80MUhRkmnPehw1mpjlXsGSkPt97r6ERJYiafU
4QSm4oNxYYSe1TWJMAaErSACtJPUfLci9aYdxzX/lrwqoR48dJZuVONkVgD8
Q0SOY629KEj5XZz43TVpOQP9QhTK3AVW5tnAUCkAE7h6Kaz/Q0YLfTq+7TgK
A99N8QDA9D7CRIAfcCfW0VXUgKqX1YdOTYg6U1OjtogLhdG8eFd8mstWveAf
RNyxaNpqai8MPydM0jIkKtTaXoZ7RzqIsqSKBiZorRB4xMV50uQvt9pCGeca
Uv6xHo3CQuCE2a34X/L18v3py47m/Fy21QoonKVW4dtQzYryTBdYD1RjVjDy
4LaP2G4aRjk4FEN86l+YHaSCU+I0dYwvvpcbINxPvlKDsJJ8+U3FQD0rnadT
R4nkuLKVm0u8vKQ6IfB6p8ZCWoBgUEJJHqRPid709dQ+jqF10RKRikJtTf9X
NHUsqvpfaaGw7EPlbhi1I+Lzbj7w69zorKOEHJoisuhxMnV9f/1OvRABJIlh
bxckjaYuBJkUJw1Hguxtd2wlExeTdmjJJouLzyV10aXVg5np2HHyW6ltIPXd
TrVH+MBsYRd/Doufzg9dytcdZIDty6LI6X+sIqGz+h8nz+BFQbYVLAdcOc5/
l2fYQb68OH5EEM1q2k0jFXIxpQGZBh4XPYOubzXDXz3cclyBHpZ65UmAVHcP
YTGxUeKC8pO8uaTL/9uhZkVKphp90GIkWR3PA0PvuG8QgofE40C2v9hR1DM7
nNRqwDTfKikxtXzg72zgKiotljWMWqDtFd8WjrXk9zFT+Mm4rnk0TwkqrBEG
0SRl2aSBDcJunOFUK3sec39vkRB1rVc9s8EB6hV2twY/Pvqs1dr1gfGoy1lw
/kP5RKVixk7NpMFdKppTVcQZgSGv0lZ3l/yRyE994kXhR1EjXEtBW+HcoFsB
+zUBujYkbcL9P1Dy4Y9CAyg2CJMMyXk6VQgD2y2mjcMDQxqWcP2P3gc+9sEZ
yev9fa0eqRzfzUtt0AjccvgqHkbQRmERT4+TNdDM0L2YjoKFxeOBnKGgTjzl
wnG/ePV2giGXPbDJCU8l4KiXvwpQBp9VkLt3W46IER0+ADdm+27HGrQunf7w
3Bq/y9y9D/JVzx8zRHVMluCIkwHscRCB55xQ2QIm5+iJxuYskvE0MZcqd7XH
ZUKyuiUqrNpwi8IMzQxvOrhoVYuCYqJ97MkhYY2Gq8N1oZkdDA1JAJshYRl8
wZaDt6aU9DrdkCyDh6vAqbUQ2gCIuMceWeBFRrnyt8knmQanb6M2vy1t+uoe
9X6Nh6ZqU2lv5fGl+bM+9r807+iDF6My89IRxi2mKsU+fpa0Tebyz2Mx0qYZ
4Est/tRx6uVAM3NBo0XYMaZy2k2QMMuWp7tQ97eBCgwvDTdmhXIJvgfpY0IA
Bu07cjmwV9pGE7TMms8X8Ds8r0ljM0lYSsg07l/J6tOyzlsJgDMoZUywSjE5
Btl2dk/iXwlgBiyy19jNmMuReKcyfn0k3Nw6dsqP3rkrgeNN+dY62ty5y6f4
+WlqaFhn3hasoaHC/qAp6XPwRfrSoKlLRhhP9atOTN0XgYOqIbFmo3KviSk3
UPywV1/1jH7yFnetY87+dspeW3f+r+CFyyXAwbPs3KxGQqt760ioT4cGd87P
44HFyTqbSoZJbOv3xXr1voSI0e8wnPnGqjjJVAHB81/gEYtfkAkLxc3IKcUb
hguHwArJpzYi8hOkPp49BP1kjPewwPJJC6LIeo44tB/On2ZjenhzvFd6Bysd
BkhygDEIofkfsljaWZZnResaS4rdOrq+Hcx5VhK27zNoJOD/a19hRhigApin
+hO3hGmXtLx1ov1cfK55PM8wFkrACvG0+0U4mgC1wEjNVlK7ybumnQFqZfQS
KjMdkMcP64ykacu2bhFPIswD/uxNKOwGVAJ1gEhY+7vhlL4DOjrOQJUZxwgW
J4XqF7hPMGLr6MVCmL/Qi1mT6XMA+rRrd+/sQWw2rftigG7HKWdaGdT5gpeh
OgpTMBOqbba4vZrkFua0jSqtxgpY1y219+s3LvsWkHFsWu4BVmsC6xFcLrKg
S2g/tihRnak4ldH/CIvBKHVRpkwpdCYVbLhhjJAehRwtYehgUsqLcOqP5Du9
UQg7XQMhGm0ZWqC2oCAUTprfWV7KVA1OLBJYGfiEpvfiAFu+GXNNV8XJyRvo
iPcZaz7A44a5bNxVYucddWpfrXBuTQhE/1TDKzJaKCpSUBokD8DCz3EynWET
jCjddfhqMsyRFTYZPlHElWM/b/cmlilQqQIvmT+KoEoeBDsPwpkcsCVb3J3m
Jd0h3diP3D3aU334jP2hJWI1DcXXlxr9L4uNgFUod79+8JwQt0j/6Sw2lzDS
1fnVOqsqTJUrLcEUnUjmsrd28sAges1ZiuOrAMfBfr9Ik43w+3SctPkx8mvM
JWs7/cJ7GBSWfWBssDDf7DMQ0M0Zo4DV2uUbtuTRMD9fDRUZFW4MXjKNQYAE
9YgBKmfB1ItOJA8Wo0xFiiNwrtIts2XuT2imC3w+ORpAFRzHJKCjv8Ey/chd
TL8bx2bP2UjknKaRl3f4N+OUJXF1VLOAJjlLzh2o/STeRAk9m7dSS8c3KQDx
CWGhy2Fk5N2Dlv0cgUuzvItRxaSj1s5qA+fe0AnqSHK6DuG8i4L4NTuUQFYM
qqYlROCN59f3sqthBAGDSBpJc8PEMG6KRAoFpl+a1Kr0JkLYHAeM0VADCKJ1
8ceIuPGnbm/Qw0e6sLWzAivH7tLYFfUyqBw3iHfxckh9D/+txywK4YnozlBF
lIL/k/ISg5s6bWccN8gqWmCjKRGN/uK05VfCcYP4hXGyq0Li/2aHInY82lCX
O8CUyvu3+gywtW+ECT+M4ClNDs3IV3SNQBB8tp1VTg/Wmm32fppv+m3M8UL/
XHX6IWeKjWE2h0zVMR8uSpeVGxJubb1IetZTNYYnHhxSF+IU/CvXnwhi5gHB
mx5FPIxqrrnv1kln0jffoCZwNgBeCNgm7leRApa81MuM7mpSw+scqGrUoMEs
lPy6f+ZtwiBwuggrgdxEKg755q9jvzaraWdS50YsMBdMCN/h4Pjn4kv0olgp
TIzCUDruX7jPYCvYwjKqaCNC400Lh79jO2g6njEVns+9Eva4UTw1tF7xll9X
yQLlzOP6Bk0yjNVGWdXdTsxsF8FfyfhcxFDlgK73rV4Qx803XUOae+45bvRc
fuRqHO4A/DJFcKp41/+sUte6ItIacnD0t5LGZho9hIGrvcc6hGb+rLozN/mz
0qOikMYjVfVPL55r5NPruUpYYexEcPTnvNzudXPDVzSgyV21nHFDGFMQM5ts
WuJEzPbK4qUvS7FksEFQuSJNM4bs/6z3F5yYLn0BB1QxdMM5aESuZDt5/8RP
alKglwRMDEvJYj8jQ3vlgjDpE/JVlW8jctalyPOB5SZ/semIi3f0eEwF/+lN
PRwBjgrJRiw7M9DecurBS7cIlkqsyDWE6vn639T6K/Kk1L4Jvw6DPZxqfuoc
q3A/O5cqA9JpByjFakK26uGfGiC7nNMAQaD3hn+5lav9fFDNEwA42HYf0oWA
VqvTjLrYdLfoyg584GSjJ/iBKCNBe3cXZzFhmHTctlOna7unnRYd/5lo0w0s
DfpNoNDr3JDZGOnbSUv6cn4B2MT+6TxSf3mniAIvbL8Lb/vrERkyWpmsR/8o
wnR1kAJReIb1Zn4Am3qPsJIuDaCyUfdLwgR+K243Z5Q5oUIDXlj4V1vUnG7Q
MB9pna09EglzA5VINS2sXdcsgZuiV098r+H5dJT+HHJmSIkqRApXd/KaRN2l
1gRM1sxxnITLZkz/qz2QhcUUGPevhdZmRtjRqNHZSiYBneRIgpNqoerSmuNa
V49QDngDT2TM1+lUaMrk9VqXU7BHUDbu+LfDpsS7zKLzx6OrPehoxLc5TpyR
wY3weotEo1pzohpWv+J1bUhLZnxz4qfXYLmF42nxAY6eAYGEyKpNDxBPGTv0
/Hsis/9Q//poCC+W65BifHmSddXRUOaM7a3X9iOKVQzL+xEC3HjZ1Gy/vK9g
pfBOO9LHhJxxXbgKlKOBCzLG89aLM66if2fBAb5/mqntTdbGKZQQJ8kKHl3P
W15ci+r+hJMuukN/mPNEtcs4CiG06Ji6hUvZZICuwSba9LEMzUITjRmCCl2a
WNtRMCV96o8AcHSZEpot+vh5abg1CWJ8QKlZ9TzEW0FVLlFiS4fia7Eoq4Ki
ne99+yY3weQgHRUJ6eUMpP1zRL1TbVigKhHjPKYmNyc82pzyi4mPJlRnx4vM
oTQ3dmwSsHcDmZ3oCaKaIU7nNbOOIi4P8k0U494GX0L1/W9a14ArVGPllJvL
t6GoxZn68CjMYFuzCv4ndxB6POYZ9RfYsyM+HKQVblkSJhPeAGo7E5adAWJ1
5/gI5R4Pv0EuHQvn3crbtBu5aClJDKk6BC5SFb/KkrMt781aXPBllUiwUKVP
5VJ6sRRQulMoJwdUT2YXPsDOiEkm0vdfFOW86Aaf+2cMIppykjPig6oXn17i
vuwf8Ms2Z180pHC55gXZjJ20nODkd0wFoNuK0DXYP1cS0zNCQGmxzrr0mYpn
e1EM2Ry6nov1tEpPPtOYjFU59iaXhasir8FC4869ABR05b/YYfs2KSk+hKDw
HJfyhSohQoR0LY1BEX6WJBXL2iCITsVThb7o0FAwsK0hyVRmA2hsvibiiezK
GnYWsnqKSQPLuM8htwUuYgVALnkXbIHTD+MvFLmXtGc9jDIm3Gp/9Lon9QSK
xsArB8qp/6vJWnFRdhHvK7++nGSFYADS5E9pvfF2HjDyGuCioBTaBzUlOAw2
M1o/O/Il8vokDwqIOGk9xWsBsubFw7Mkq8jCHVJ/06whb2zWC8mt75lF+jDR
9D9YoDUK9NZaQj1ZehplrSBWe/7P2e5VY/asX0GgslDsY0dvEJvBRvQ8wqdo
YpOuy19M8RHPr/qUAZkVkhMyrn/enRkisIpa5QBEBb8itXOWYIM0pBSejsm+
uF5kg+T+uktgY5ib8KTdUEF5Q4AEuiQhX3qGhyYL/CDQWtTlZJvsrF5FItOT
k2AmoElSa2rRjytFOrd62ngK+LF1hzruUzM5VtAZMIednZEx73Ny54BBEGPk
nLqik2nNf36x2+qdeMpfpuJosakD5SO5XrC8RtoYFujV0qd2+FqP40d8ODbL
G6fNTr8JebU4MAk/99ObiQWEZ6WjI/YZGIFJThMPj2FfmL+64hj/dhZyvBps
glpqf23iH7Uc0pR0hYYAf/YfKn/pc7rI7zHQCsN3ncjT4BFYvHmErr6lfzao
RekFz0OZHV7+vFiPPRx0LnjvpeHKG4ZPNZFRT8QkS5Xtfn9wisocjkPtrWl5
jUy2IpIdSSPANx7WL4Li0FXpPLme2H8tkKgAl/xbA8zcLBmahW1gOzWT6Bg0
Ls5PG4uO7M2E/MSY+GLIhAz0Qy9JzRSCJ3z6enlcE5wEx8wxp/O9P+9ACnhI
o4ZXLsd6QTM/lKTpoXs8lJntHIDo7ZQwU/0HM9A/Z4mBbJUzFd8LWGb6QPd0
r52PiK06yvtZaOjNtWa5vTwykTOg9GDBwAh8ybQ1tneQShrnKIGzLui/Nbfy
+m/EN5+F+qLmM6flPQM6o5KfGpa+I/CuIjPTbLaQahirLe6BrOVLOpj+4sh+
DfnKyfUk3S/3ek8WHDRLeQxRJD9RYX6YXkZylGT5zRkDfSu4oNR7Jyq9J9Id
/lc6swmLGjT4UBX+gqhfP6rmESd7xl8tWZy5qA3/uMGzyQIZEwW68sE31GlP
OAu0kcITIxYI02lFH0ve2ypOmkFzBJ9WhIOTuCZluuHBjoXo7Vjy3WofvxOS
4lzifz3fZrgMZRIxv4US7/+BLem4WUXRv79Z2zD/KrOW5mWGJue07k815sWd
/E6OvmYdWcGCcMNCRuw4CAtlcfxas2kv4shrTWX+UtZj2u3AhGXDhZVR2q8Y
XTaWkg75UeMW/rfQqr8H3w2eo4jZHfDptcUk85CFvK/kMMlGkFNsugCUmTxG
RWXf6dMPnbw9UJRn4Qx+fPjD9XfOcsxOrczfO0xOpkKIoS3pDVBR/5oa+22m
vbwtnmNUqbQjIPWmOq+UvU3X95Wulk5kBciRj9WGnns0MB1C3EDuodNx+Di1
WvNVW3tPkGcQm4x7JcAvFhriUnsM7V3pg9wcEUTdMhADXSI6xpsV5hZGN8x5
4d6p0D20SqYRqq1U7YYO5lK/+t8slZEW7V+6SHa/Gv/ZpOkcqKM7Nx3T38/q
nmrUfSWbxDkDtTfs6bu5bhLjBnv5LLFpvjviMyUdUOO5ayIm2v3z61kYwRew
8+mg2zaWYfEMWTw4KovwuZB6c14v6ageHOWzSEJnX1ycrkH1OTX9/vcJh9sU
TvLCqIVltP7veTneTAIooE/hMFx9kEJRHjvJSIUlRp5FOPXBbKnPigq9tCDU
3l/ghd6/eJZm4rAvSnJ4DQ+J0d9hPbOPeWNniHZOiO7YjYg+xECr/HIbnsJW
U1pXBN6gHO2+nxtVUlSWgQNrq+1uoDyEVldWN62L2TuLIpSVsK37cAd6VqdE
lG4KqFmAzjJsav0Diy1cd+MxHMe7ZEu+D76zOJ3FSK/d0HM3tgO2kua/Td4H
/f+X/Lb2bbz1q42qO0Bk1U+An/NHvm5IExwVu5ybGdgYWlPj1w80LhnJOn/G
f0vXbAKooxi6YWbrv4rn7bR+lGUwnKYFPdGmLPZkJF7b5FesoeOzyxDOQ4Sb
kriUyb15M3e3n2UWPhr5jDeXMCJ4JmQ1TEii98Dq6UuF+3MXnhzw1zc5a1hn
5cEiQoqMgcTL/df/7BuqGrhu51CUEKSeStJW5SKCmoGU2R4sRCZ8X+mBo7T5
XcKj5SdvCUbqA7FPzFmLQRVyFV89uLtfrQUHQI+3o6/TzLxXE+RVtyu6vWMv
CD4Pm4FXcgCb2T8rc3wfT+i4zSCOlP6fKe3yhnTctjbRLwwdHJXGiWAy82AK
sMxxhBhYNwfgNz1t2RDkteG2/dpPc4GRed1JzL6Nq9lEtUEF5FD4g11lF7xA
bRpvUpbI4wbY4mZ/IVkmC9MzrO5WDCkA04v4TaliSvOY1dzgfufkt8HKZQfy
gcpVjD6EH+fRXm3jChEcSYnUFKo+Eiv9L4xN+yk83qsRapOKn+ieOG3Xv40H
/li/cfv1Bjx8eyHxqxKwsIkH64X+Ekx2pNgBsSG88lpP1b6h68uE/qcYTyIf
drR8kWNO6lBbxxHQ2Saie0o+wJfULe81B74TByc4qeu4WJS/mKKZfwetr5c/
DeY0YFSqESB4lXyr151sguuP/f6FHDqKNZwrsOokHZzF7Pde5U7QWCIQnM6N
uFs0F2nm7zw8FbOx0xMjDvdxBsOpSeohz0ZX8LzsLpnWkpVvLp5leFIESZGZ
Bj7Xi0hWWs/lEw5pIGlpkXeqyXKOINvBH5OsL1jXOnoSR1ZoYLmbR+TZBWJG
ObyFSiNjU0RnpoNru6D1gBRbTZZEcX2BixK86QN+N3swt0J2nq7dAz6uQsEU
6S9rCrNAMKBwPa2fh4NjBJ9uj+Mo0X5aGVbZY0l+T+/vmZFktl6SAh78DXm+
xOgHImITwSY/wM4vDXsp8g3Pr3vAI9xa7O1HZFjQziqYyjQjMdLEijL42kW4
BUWzFBGutu45XjrjeTDi/jBF9K26CkwUWwcNl6NfZm6BmxZuKuPYHUFH5KlH
2D3JpSnJoNtFLLG/Ay0PquJvOF3z5q2AM7APqdiZiMkiFx0AYsAQwBqciIQu
QEuIOYrvk+f7Q19dagwWwGQxlyQfbelXBqiP/1W4DLPs2mA1DkxXr/siDMas
5X/SWcA1pDCyrCPcrXmeasxA7f0C76g1eB70H7us8DE+4rCK3AMVkA3iC54n
WBp/VognXE3njq2o7WBgB/DD8PFZHOze9JPaXMjwYLN+tAABxoUYKh7s8/KQ
jCGBFqxiV5fZUH0EYB0rXBM/ws4PnU6mBnAf4DxkncLWGp7GlrguorFbk7VP
w83sseqYa9H1JMi1U75G3tWWN3G5KzFDAqKNP3KMYksq4y4zEz36HY3b7bv3
GDUzD0z6Jnv1N09XjqIadsH8QueFcFfl7/xZ7Zs3pelIijUVn9JPvD9Nkqe2
NxLypLB2D13GPJozoVczSKZzMqcJm46e+oLDOq96ULoxCA9/WA9hBp33p/M4
NUoJ7EyMIOy6R9Dba/sde95zk2dguDACEGaJO8Ie9cWh2XKOR7ewIvldyf7K
sS6UfgSAyz/PdIdB9SgxeE0LgfLPoaXCSx+iwZrs+Mjg5weP116l4PLZpZo6
nTTuR3ExjNXBc53IkFUlVTU+xItrEFduAgMlv44HUeRkCVBvPh8gOH6WBeM5
MLsm1ctNVkTJkns11jf09avYAciYMoqBhMqlVYVBBHAJGM+B+EMY76rBhicd
iYxMIu74QoYZTg8POw0dI6yIikdomtVdMu4fcDalF+5wrqVf08o4Q63WejZv
hpmxAjioElNxdbT1VRY0rTQg+DIft5ERIEJmiT45o0I/qdmpjXfg1G38+FN8
/4a80Tq+5Os1ZSYmAdMbD5IPMSiG9iALvk3pszPr3OA7uNqSEa9uEOfucnga
a98rsa4XLp7vDWyJZF8zPTH1O/eH7bAGyo9oN0v2AHhXq9vly2jJmRLCc+nH
UgZIEr5BQsH0ybaqbk5CcA59EwQDvWpOtE2iXq0+LzD24TgYt3bpDkwA5DUO
P82GfBuGVKo1Y4+BZw1IKVoS3Jszt2ZEKLHOyOmWjwIXDrNcid5fws4wSZ8r
rQSj34JTMfaI3h+Tb4bMG+3Z2t9EY6Dqi+OOmMq4cyy0cfadUyACiSdCKwg8
7rr98P5wJNsTYtR0GgN0QV2Nk76rfjBg9f6uDC1A6sqVGB1AhT0z9s4AY7Ko
xUBch4Q2adFM2Dce00qwrlFCrVlhvQOWrlJ6/ZewQA81ukZ0T0KlSLbViBa7
jnZ+lwLGjorcW4P2zxRFPun0xHzguieBU51x5K4CnIjKJCk7+fzTGRSyt1kz
v/i/qLdzq+atuQbju68n3f54VsqK5S5QjtepR23eiOQdAgQfnJzwQLGVgfab
sf+mYeqF1BtxVCAv7UpXgl3LEoqAC8AYRDqUx00mPauT1xDfcvhiENF9vBDV
y2fZ9pWJv6JKM2of58QW/eiqlTlyio3bjo1mvFCmm4I44xFe4G4158Cd51yy
aJrJNznFdb6kzoX0hJoEcFtmEFnO9HaavNc+oT/0HHjXjXtpjTE4SQIHbdxr
GaH7IPKC0qYGfu/RNzdsO1q4iHi6Jv6sZe20+8BorPz1dzAocNQwKN6c57dB
rXaYP/yiDcwtO/RvhQy1CDRDN5JlvyzB6PFDHqv7NxM2Dyna1yzR8NLoiYk5
6sRCEeU6dO4cUPBp0cHjkEeZA6fqMIcFdB/1ZsvhzmzcMfUzaWBmnTrBn7Jh
GuSYlVUNLwfLmlhZAUJeOb3xydg17GxY3n+ORWCBCxTASa5Z3eIEVASHsk4R
7jPW0DrirRXLyec6iKH9c9KQCbxQ+s176/Fizh3oeY8h2c19ec+p5Fwt3UZO
lCE3GVE4qjt5SdKPiDEoeT75S530OHm0AT/Pr63Lx8GQR+58jkoJh7AO7DdD
PSErgM8tkTbL4gwykhPx1NLZON17o0avQ9tInqb2Brm0+Jd98N5WU969Gizb
CVfbiwZfbOuQAIkxojWU2nNrny3NVOKWjf+QSEaHvoWLTFsmfxivxOpc8XRf
TJxfqKTU2PD8dKwxOr3OimdcAcsBjRU+vN6bNuy64hfp70Q2SNUTmDKmn+Jl
9LSOsPq4mODL6rmOlaojpuqk8sGkM2zE5aFLaUMFx2Ni2Fa6jPW2sskkpdmQ
oimSSFYWGkQzg9vHsbLYmTRXe9VcmFzqP0YZMTw+7AWe8bLvJWdH1gWTCS7o
UGGWahTGzYX+Zaa2fUMX8+1wZhCZl0rr5bsdBXgNlqS3QEzqAh1tf/Cdb0am
hzxFv76A/aXgrQs5NscVjAVaBaXVBS/JnsntC74tuCOGBckrnJcOS0GgpLDz
fyIKSlZVKju0Oc8cvOYPgadNWTl35+gpy8Hji48LosRJhVKxlGfhiVahitSX
SI6HjQbRVu00/YfOkbkZ+yE1wVJT2W4gkIyr9oJh9clpedTlbPJM33d2/BjZ
sWtTY032yF4k0OjpFs1/qjPlTYfws3cBS7vGOus3gmPuf4S1EKi7LNUk0WPm
FP7z+h+dECs/k5qIuNHZFJ7Hk/4+rotXoZP6M8kUN2+cg+gGCcoTs3rbYweq
FwuSg5Anp6EmBXn6EfKbhZ8NbKlmfaJQgAaDP5x8PI5j8oGTQ8irUOgQU33d
pFtegCSth2avjkxAHGi5dZ4NA1OfrVRsrAPfMZFqbW2eFoE8o6HdWR2KMG4N
OiydYq2Mu5/j8kav73aTRWY/SY443oIXwZERznWTvDYpLbV3+7SLaE1S1Zan
KH0YF8oNwEl/wKF7GHvbMLkmDEpDkXAmk2Kl/NP0Z7mdUg9U9GtJNGkiiyKb
eucvpgqlToXaNQbxuE95QTAlrKJ3ii8aScUV36FDaX6ltroVKpX2VSnwNLkp
yWzOjLDaRFlpABgcPiCCH0OOKXm6FpwvSOXVWEpQ4289kmcnblAhksvLTPcv
g9WuJHnnPM205Bj/LuA8kVNR+trDMEr5T4WzVjfB0Pxo94P48/PCacpBRy4f
2VV6ehkwrjIilpTIUkYELMdqNFMVzDG085Z6q94WUuNbfGNoSvKblPvafopS
50yRvuis+JjZT0al/C+sDfpNcbLWo/CI5GZELnwWtF8UVX5dn//RSGZbikrX
tcV298fqMQ/Vg1fIf6GG9dYhr3lLubIisaBDB8yLqCQzcBEYsXkhzDxxEQwX
nwOQoCSsvKRgjX3ZsOK0C34OZtGKBIxWssZiD8GcDDzcm5/tYiyO80wOl3as
7IJD5wN0LyGnq6DgwGFQzg+UfSHeMlQSGAxzEfzi1n3FWT3dccg2aXI7A2Dt
WDMj2KWiRFIn7LBQ3VMZoI5k6/A/ai4O8UQzP32PvfWUZiXSrP+JrIgwQ1cK
FnviKjMP8WYw3bnCJCz64N2/7IBNydo/5xHUALFi4SJWwt0ZyTT7t6qNTt6I
xsUIGX0G7XTMIBIOOY0evmvct89SJhRJYiQEolBggnPTJgjHU+7sGFLnVF5c
kVMyrNMiASDd4LajPDU4LLa9uaR4BsCXBA77d5RIg52SNNQIQw71Qno5qZEg
OSqh3GQw6FVEQny/wKEI7NpKf13LPKWXCZSgAVw+y6asjJEtvpamIy1KDEDY
/OkggzcdSdHy6Zz/Ue3Qi+zf/vLDHW54lbcGDMkGhNJ35EUhksXPKwUjHR0g
sIH7flq5Fpsc5QJ4xgo6YsK4BOXKHyivB5sYC7bBT7OuewB5olaN8T/jIGR3
xBi2yWPdi8Cfbr0tXRrMQnq2H1viOSnDO7NvhN9kn5AqAMP4ga9syhzawzKD
DPR0Ou1UGcDMXIgRIsOSKiSSSo83tuvm7vJgsy+QZ+hPf+lopGB6NB9J8CHt
Zyma6KyOjmGs/wYz3qOGQQKsCKVRqkhtqmFlp6qnUpoVwuwoJt7/rpx3pjjX
2JVF5LUVHbBgyQahn/SWHZSDSoJVZ+3w1296Xi0+xscGRy/AklS8JOaCbPpt
jPsmnfnkWbHIDVBcnYWrIts9N9vr05BTohAHIOHZkxchsDDui4ZmfjLDKSEX
RCysz2Vt2XASjLd3ueDwfxDPk3oARatJZTUzhtPBzhUysb7o2k3vxhMPaL06
hzSfXJooRvSkVWgKsdJ2CVlVMgwtF7KoK8u80k056MeE64YMAvChhiTSBtum
Qkibll6W/B603UXs6MtNhIvSs2UTXkvfWs6v7wm4wIVYbqXM7Xt/JTPmprmK
G4+vx0hO+zFenstJkAUSxtTvWBso+dDQG8xjSYRlgxpOxM6cVOQ647UKnStM
5GnMO0cdQjrud0uxHmmZ/MdMTIFohF8jvDP882YjsfJ1hla7kccluLXj91Ia
RE87ujqTGXYx1BfpDeyJMqIvvhLCDi8BMcdG9KLWd0xiNlBBenOm0+uA4ZrB
jzuq01xsI0VO8xK3fDZpM+8x8f5Dc/E2ZZnALVwT03efLAUt/WOoTG/Q5yNg
6n791BWAw3l1Tbo/it1MTgu2PSvqg9hsZ41ALQzj0MCN7V83vBVISaGE/0Ie
ZgrgSdZcW70KfTl+O5L8jZa36BIGKaynkk/Je/PQDMaEdJaRdWXLpgaRqT5O
j7ZBETutANBV+eLngQ3k1HK2KlIRjLhBdGW5mnxf/0h4Orzx5jgueAUIkVuE
Qymuo1tWzcWxjCMW8xw2CvXmkSrHn0eQ0NnJRt7Y2BXAErGDiIgXmdxdfAV4
d7IhIxSyfUfy7kGu6OFHGAMrbjlGZ4sNBkUZSf063GN4QvHye3lCd1FqYLdv
VSht6XbXewdSkgC7Zmi2Hld3zDUEApvCPtnGfJMcQpXp/UzuJdlMxfkgJtTV
FUcGNGUlJ7I1FMzsgI4A1a9L4270W56k33DINoGdi5AcgwLwEqjdp4+hIp0w
2sAAyq0YaA+U6caD2dfyehwNje1XPul5gtZahp9U/o+j5rEeh+oIIZib/GVc
f6xoPRRmDK7b99gfLC5kBdOjbiVTtjKpi6pD0hxqIunHcwC0iuhIsf/PdkO4
+SMUKL2avjOCnWG90vjfYacMuSzOMZw8+/eMiqXN64Lga3PhHwx+Y27dzSos
UHDQ52wmw4bRYoqHpurcP2+gCNGJ0/cERZsA01oh6BBM7fZLh6K5gj1IY/xR
mpRklNhcPpX/16dGaxbH2+hO5H/2Od+SyFOieHJpucPHT/yzGOj2EGQVkOxZ
QTLS6GfsW/wlANbq11IGO5PPbD09G6PlqGQM/Xk+JqC5nfhNC5v22Uuy5YQq
ttT/0k9VfSPf1vY9EcJ6Lb6yOed8UVkYyR5xJTWANDwYuvEPpi8l2cxMdVux
HysLpGL0Bj02yFuVEE8YtMj+uYWrSNC2k5fBvt3LhEeDFpk6WI+OjAiT34xS
05CHvNPsa9uMllZjvwjArWua5fEbOkV+g9zOdh9tpGWyoUAv821/xLKTZQFZ
61XkJYQWSc+Nddu8tDTg+dEwZsh1XmFH212Mk+NHe8JPy65uq9xVxTb6x4Sm
BV2lV2FHSwMuE9OHqIc7LoZh/FQN/jHwHQ7TdBmzActHpvbe0AMzMYkLlfew
9MzKE10pB5Fsot2+38aiS/rny8nK5wMf5e0qqmTR5v4UONGTMjTbWyugd9/O
JMzAFu0IU04jL/askNRKyCYHTHY4yeHqRSvCGz/003SdosOigDL2Ixn6MN5q
7LIFDw363pK/lI1PbJurDq1xRn37zi1TpDG0O0iidzC5tR03yXqNNHPKxrBC
sQZ5wyPuuHohvATwWBf4CKBq3BXWv31WLFyTU4kO4GkmTp0e+OgnxWS3BwAH
KF/a4HO1NnYephTRsXzoV1LsGnGioE3iQ85QcrZv2FszS7J3+CY9hBEoWdow
gcwfGzdGzYEctVeivOghQsZYTvwUKClR/W3IfdLmYr88gd3aFLwn4Tpt3ZZs
lAEXcnijBKzjrNhRDdPbn902REJtRhR6TqZwqVbl3nfZhPSm7yDHPMizZtvi
5rcc2IjuLxWobrFLSiCHEawxALzjXUeQ9TbjpabWAnuZQO1Ot/VvX6cH22HN
zJpL9F8WQVwKSVQ2hNRTlUOUOE8dzj1/Y4sIcrabb3RHXCiDqwI/Z9T1f/UN
D5jDp8Nr4Le8gcWP2wb+wJbK+Db9WrCayIVJz+9lgUSNSe4MdSTx9bdGkx/i
Jk9cAA24//TCqRqZEz+MsXEk3FBkHgxU8XgHKR+eiOffJRov/TVWPViM+hgR
TNm9C/UwfdU79c/6ZET+w4U6Lz90/DUh5Hg1M40woIIIKb+tvACyqU+x000f
vjl+OzHMLpiwNH3ZrN1UDQW8qd45xE+v4XTCYNjjT7D/2XnAwvGhqa53BH2J
Pyg5Qsz9dE2I1xfT3vZoV9DesrkHDm17bkbCF2RTqxKb1DjxMsMGaHuwNxEN
a2j9FaTn3CY59O5p+9V4+v4XNHjDTnNzsGdHAuXWHLttMfj+/DOkCi+A9s1k
2RIGzfBg/2Nw2W6bzG5TqrZV8hD5vAumgeQERmGUuIbe5Tau4kqceUY+mqzN
NNvpxemz2XaFSYSAITDZniAAnm+UIq8ptFu1VfHp3tEGvE3gfGsVeYKSYYF8
Me0m1urVNiNGNKWG+MMlb+0VqLqioitM4JBdbM1eyYq9rMfbydlfA25tRpi2
dgNKnvCAQiDDKOG7nIE0iGdIAlFfBV7YSADcAAhpneOMTkoedC0lXHdjvH8Q
vQ7+8Pfn0sw7XXIMoTt9mLnuSVnycqOL8xbo6OdGp42LmdNIeRj4wxi+ajXt
HT3B+4AAtokCcakvPDFC0gpeCoY1u2+YX/b5+efkA4Aa7BxTO1FBYCmPT5Rg
9M/pRu285hoWbZygs8YSAyv1HBa6hm4eHuEdChn8X6uXR98o3gihi7fIm5b6
nrl7xc0fVvFXLx+3lymZcRaf9QOM3ULndts3pRPunydsJNYgZXGoXiRATqMv
j6Zw6F7kp/ghwdSwWXMrvHyFfua7Bir37q8AOf03oCr1uo7HFqsO6V6M/eKf
6Hiifo2g01NgeuNRYy5wD2nYT802V4JvgP0DGGnNLoZ9APM9qxER6pIzvsVO
e61/mnACXdeeFirws7EYkxgOaxqYzIaBNNNtHutHhmEBYgNdRsA5jPe45UoW
1PW5UsK1yrdObvZLlmKXlGSQGwCC6b2t+KaE51u8YaZWNbXO5B2ZdDtj4dMD
BQl/byBpN8fx6go+bZty9ie1YgXRjbRwC5ETbGW98UodL1LBRfp6w7G7jbdU
JY3WGSSCowPNaXdou0luP+trYX5DdGgtkRcfdbucUvwCd9cgu/bgHK7mT8TG
49MpwL9fQSxtAkZC7aXZohbYUVFyqGKWfHMlbvCA7K0ZxPhmIdWcCF6rG+fi
eSUlHpA0rXZsDjaBybReKGxXm4XXRqZhHKa0i15xNrGp8uVLLOaJEECcXHPL
YNyV7rub+dH2FZBQXaPsJB0BE13ldUQP8nozCHA+N84Jnw/R9xHcSH/gT8a4
62rZzzdadth2rM6q1Li41YcTb2faaFcCwSOxymsWvx+MaNjZYx1vDcboKaIV
xz7g4TivnDyqXavtmY19DFxpEEY8VuFPPkNO53qZ2zf4gC/hyGwpC0GTzcn2
mvSlCUdlr08Pn65pe/9xpGylckcLty/2yL3DWnHUy49bkdPCx78kQyZr1fIW
RBQLnOKR3rbWTpj+yw9NpULFy3o9Vp77ZhW/O33WX1LYgnBrwtWn0VVY+lpb
HI9r4YUOs808Ax29mIECBw4upRhqFQHzEiCeRYBwzPcZTQyN4o8jeh4PSXA7
Tez3F4KQ/p+FGIO754qm6Bamhg92+XVzAV1i7PhdaRJ7YJhLh+kc1snp8A7J
yoV3By9j6nD0gZeFdAKcbdGZm1otTMxfsOKX/FRVi1Ep3gZTtcKFc8MWjB6q
DPvJmjC4KuqRCAO0bKMVwP8u/syqkL+Z2m67UGAMEEsr1CGvKkkSV+kiyRrn
WpcxYV8oCeGw3Jd5wv9u4/MDzCHsgjelO5d+xM5TDqDaj5Joy9XquDGKeGh4
rfdsxQ+QarBl/GqOS0a7+V52CY+y3dcpLk9JkCzI7WiUs3AnvNboMtz3vfAX
p/REAVHVYlYgfaHbPXWugO7a5hhR1Zc3hRm3OOeU7Fr/0pUBV+Pp0F9h+9xP
IjmSuVkEVO6Js/2CquyI67NQEMtt0HuDMKz4VNfZJOE8bWVe9yAVT/NyXvA5
eUMwgUzYBaLTflK0eP2W4qQpfjEZuFMqQWwYAJKYG4dyGlx0AA6RZkGbxheR
Ql+3puMfVnxjT6tlcfdHFcvIsuovjcnSWiD4AFSjPxPwtipYqCu1ygOmY6p+
4acrg3zbT9P2UfRVZbeHqsjCsbOYJSscuHkT09swiGrQSzlNKghtphttxxxs
m3K3Hp4CeuK34KLGtyy9vx0AIzMKQ1YTL+jaG13PRWusFvwk3PNzlxU5l7an
ug1uKiIm0xG1o+FOe9wyXGxY28Zb9Z5jY1UkS9HnXfWX/d6okyTVr+hzpooG
We7e65/LSBDyqPx4GkY7MyZqpdIKT6yC8fXOG0ScESqJ+4S+NBqf3kQ1Zjfb
ydZkpgozUNSQs0l5ocgcayCJkne2QQIaX7dc7BrEq8rqt6IJ0Q9NSViZFoyK
NPdzviPGTKxkBKh/+avxnMSTHEEmVtH68kY6LGNoKz2Tt12WfNv4L9L9GbUs
SZcXD3tn2PmqLizAXrqJwoAoBBn6ItdEyDSHt0D89+NIgfPr5rb1fXqdxFSp
pF3j7ENsJLEymucRCfZauOOewhdQjyGt0U9ug7waP0uoL7suyGEN5bhd1HcD
mwOlMXt+s5i1WogVxwexJhFFx6vbYOadgN9zXwxdIu152VUyQr28TvyD7MjJ
U6jGgX5wN4MTXYQJ4TeFWRHcULX0wiBbZ9qceRrqGwfVl7PC2beXOcjy5kKT
dqd+iA+OSSpqFxSA2ziVavu5DE4LYe+BsT9OaFWnEZdu/h+nKVHz9dYxw5nk
wa0/BI1pb1U1isaST086/ubWZniqtfmbth3lLggizzIBv7pw1ERtihoURkYX
Y1Zr1NeHIQaa7F6SqwGhrl5NFfIFWLFzm1aokV5cNlL1ce0JjYg+j3q2YvTI
71R0GgblO3YZR/C/dMnABSLMGBtLcX6sIZ8iQuBX2hYkTA4BlKWmdIE9+r29
35JKO0jpevYuqKz/GDrBirDJsoDGlc/gymFN0iy3OF78qUBrTmyA53crR6Zn
E9EpH6hR+DqM1zuPeKSYyixxvfbURT32XWzkahNn7cXi6hdVbqXFKvmSymjs
ErJrfLYnfMMPUA0OuHvoos0I/0b7TcTo0ptSs6+Gz7opzaAPKrkJPrl7k3QC
RwGKCuoli8EqDqGe8+/vZ7hssUI/RqHX4khh8sbntVGM9ooELW1BLHw5ntzS
HINmxU8cENQ376rLSn991b7jmJqFh4BkHO2/unS0b2Y0pByDGSIKczqB9h1Q
88WMQVBPToYh8wjrpeBXh4sqY4MicHL8GAB/czLmUbSPPjvT4TIbPb1k5dix
QoYsNJy89BwD4vIzCo513URjuLpQrQE1Nx0WmlW1N/iNuej5CBqNzUGqlgUI
FEZAHRPsAJHZd+oiFPYeyI2SUkonTAETW9MVfttAj4F/YaHoHYb4Zat0jw5R
rcuVVMTpI76pfcDcxSitsyV8CnM6oYYvOcdSs93cWJzi+yXqKHrTH06iPOjD
YuZ8y5QF5OUkfaf7os61uhy68Jb/4UugU5B7u25iuoelRp0YuTjz/F4CbunO
ll7PGy8z6I79Mbzp1K6jRhaK3isFMD6IrbnSHJk2pbnPF4oJpc2kIj9abBav
i8a5dorZ2oEAWGxBafEHN8IF5wsD561J+J2i3uKz4iN0uPHXglPzLtXjoFYY
Q8sRtXvKVOWTqL0JRaWMkqzhnE6hilVYvM2awXw1nmZqCYDXmI22aP8b5OB8
R9q9M91m/UJA7guk8Ui//8MD2mg5WWXYsb2NDhXKcy30oW/ekY1pRXNvEAX5
84E0KPZKPNM+DGPgXjp/NcgW3SwVDRMIuj7B7SFBCA5r5rgXWtONZl8gs/+P
6x3NEoax2zFdEfrLz064mFHv7UjYGdp+vVC16H0Stxa669mp/SdsSP0+pOJa
mlpcCWl8zHr+zno5Wmd6mgLyiX+Xp9cJiORb1k2+6dM9v4pEyDnCizHaMOxB
9rh38v+Duu+Nj+CbzPM8Q74XA9KlQryJAowlOTHcBDg/WipN+7im+OMbT9dC
jLjmIWvXWFEVA/7CCbHgTIfD+Hbi0bbpBhk4qyeeJhprfVmBGXUcKrOTI7vw
GkhVbZiRLkMvDtpVRQ2DXHRoDNo8V3EQepVjNS1lS4S+NvuAz5syPvTA1OMk
9b1VQDtCOU8AU6yVNGfmyhslgj14+zYFwkyslJXkkSiSCWMehEgBy91DarYR
6Uv46v5mZBYKNBjlMHDGg8hnResb4VxiTXXflRQkaaUL3AKWDtCo4P2f+K6l
UtGvnPHx+RtjARecBRsM7ha7d/Y6b2PknEB3ArCpx5bToXH7YGrbpBCObx3N
R2kkeDK1UJKsYe6v7lD25RuMUqGlzsA6DB/1NukP5Rp9K7varcUPLKjZJSWh
DgYO9gXzL7S+3gzdyMvnuJvjLbzGkoF08LGmF7rXKybNvzX0i5T5Jm02iN5G
lS34D1Yp4WVjX2fayh2TpQuCeAltq+IfB1LpWJP6qIqcmv6zJ9ZTeTEHN5ZR
sMNJW0jJgi4ZoB68WuPhQpE/n9k2LJyyrpooWSbH9bvYjjXjQzQ2yJfNfqpm
4RZvG/Yiv9S3dy//nnJDlSclMWzq2ynnYucZwRSxAVY+aSEGbAJb2eiwP5sW
GOwTBETEKLphygdSrkuttKTxQi1MrKgkPKuGYlZZaMa9Ff8N/oUixxuNBNDU
0DzCXInnkVd9ybPDn8iLG/yIXLaWSryQs6iqeNZDgQMIam2L4oq4VVDYKRy+
q0QAcnmrSzxDPODUI1wVj1+SKDk2qN35ZYaltuIx8splbCMiBIXiUxizsOWp
FWdpBE+sMdsSR5TTmRvqRI4HlMKeuHvbgPcJG/Vyok1S6HKKBnREWuPSOeP/
hDelTCXIcngY/GzT0aIyxkuKmbgzv8kJOhe/C8F2NeaXAF1+/4ZNNW8OQe5k
mCBVcSl6G79GpJF7Y2rzcU/yYKGR19wZLvg5o5teaT/rOBrpV5R45naSfOEJ
nAyvCWMr/AWRcoi4WMP4zhPWWGXO3uwIVZhAJUsFiTGUfiAaRMSoJClQniDJ
Sj4dWVGrhEOxCZ8SIX3ZLON2BviN09TGYqvf466LLmND4+aHXkYr3WMBDO0O
0RLqilUW/czazEn/V0YyYwl9UW69lEEDZUG8eTNyazXXfOZ1UVY4S0qrTuRc
zdIdUC36PGASdO8kkq6g20f4AVsBnSI1AxevjgcPzntoULdrAwGABFrhuUCJ
eZ0Icns6faITHKZD8vUJgInEj02DRNTsUq9Vtq2RVN4/PMo05iEyrrlXJPZO
uQtJZ3Wq/wbbXM7Vie1UZmXc0VMbz4GebSFZJ9FlDntCdE33CCcxzZ8dtnjG
dUwzRkmp/YCerQIbg6XZSBabob46eVnA5oJK+QiWMBlD6kWliYNFrHFcKBG/
/WVYuUFEjvtXyXmUknbBpIZc3e29wxU4Y6G2Dqlnb5AZp3S179dy4/tFC1Di
vcQAWDalbq5ZhgdcUMIqK6eCvpqTN6QVXLkxiHFGbmK1ukAkmlrCpaqmnwQX
w+26Y6rbqoBVrrT5E4eC03cDQ/dkI2v8ypbaWZW+MLf7NfjteQ9GGOQT9j4a
L/sZt30n+vloCtE5JRTdt8asorEu4NoCU7nIPSFxoyLELWwJK/1jHupbfWBd
bG0TPViGaVVTk4WYWk8DTyddSbtKRjSIREXO6JjL3RK5y5+q8jML0eWO75kH
CtESO8Chc1yhLMq5zy53mDxwyq/Y/Jaf2UFJyEEW5sNYeMPJ63b2jc8R4qF+
7VdmYAgX6M/pAarxUz29vGTmE7l9Ez6ZSukXeuC1y2gL57QiZq0mOyjfzmQD
4goPZD5GMtyxQFlsfTy/aqFiI167gVQpbieh27ao5Gz42x3q63TAkqnt3Wjl
Sc7/P1YzwM9JF7qtnDWBcRx4HOqCgnZ9jSxfob42bfzlpcEJWLXhRM5CTIWI
/KjoJHR4s+UGaxd3px0KQxVp4dxlwj28l1OEuiIWd2E5AOzghdsbBFtHshxp
8qOJlopsQN7C+ppoMGPD+bpW4OIWQYRaUMj36PhzgWAUkYJG3g3SoOyrp7+g
5CJYwYDap4NHU0VTjUIiRHCR/gtiM2p5vEGd7YXnBAbGooQM+GiT56/HBzr1
DKNDzVZ0nJ5Xx80LL5F1MbMlD+hQ55QTtJB4xhAR3NQIDfXibOXzryesNV/4
YZT+9opbpIGknek12WKWdE+KkRcPkBnZF0sCFYMP9+EQ7G0ZUoaTR/bLLREQ
MhqQ//BAaHEwW4XYFZHvTmP243NPdpsDjRX6Kv3AoJ69rd8d9C8lc3LFHbv9
Vf0JVrxntelPjdlsRWFl+HsI2xGlt1YJizScna8Gox9IjgbMNjzapxMUT50r
thwIYJ+GKgV9YucKRJI60/RZvpR5fROjXmCEuSXp6gIuRN85kmtg4M1NOj/l
fASQl64VTLEpArIyt5LA/KMp5YFk4fgKqLhzQZbUa9YhQIFmodD5au7X+8iY
e41+36DmVSqZUTtViLvBN0PRZFRCajJ48708LpKHbokCbTC2MeRq08BKJdyH
dNDWbpa4QedXvJhlphy01hS/GqVAJ2lQuoEKYVFV2lr7bXmR98ddM+HN5nkQ
9J52lS+Wjp6V+6jriZzBqqY7XKuCg+zbZoZAqCIfNSUVk5Pns4Uak+C7fgiB
aCxfYUNVkH2SgyIa2iZt0Cnf2upw6J8TQpRUJP9KLGl9QtR1CG2Wk1Kr943Q
m7HzmXihzgiHVVPdMHRIPfTFvKHYNjQKX1TWEARZANDX58M/iRX0RGifyT6y
XaZXjbwo0HqWR1pQ6DthfmsuK7tZ3hjJmMOfgUx8aquI1JqUxzfqFA7WTaAY
nX36PQMSfE2T9YWpYAbpDiyFu30Ln1MnJA3fTuUP6OEfmjb17mVopwmVgbM3
a3lZ5OBc+/4Y4A77Kr4QMivtHIxrcFnR80e8z5rLLY43lMU5jHNFOUp41vVJ
L7g5Ij6+S+17V8/qDoQRu9fMbfs0cZUtHJ15FPFusFjg//gmW6jvyeFjCdrH
pGX6oPo6dDpWyjYgitm0p5LS10CRYazwwe1wjuSQvEAZQph6T9L/dDl9U6Gl
NDV5QyBYJJOTu1+jIUT3vtHGhaa/MDpRkXi9/DM0CACHKPBwiSvADm5BUrx6
58NP5FMq3QwrmMUBek0yhkAcSRa7DPJQ7xuzJDPTefIkhfxJd0LCPdWCmLVk
lLQ1TErMNKOdrZjUJ0zl+jwMJwKUKXsUWwAzgXnEAYL80iyjxv1Scf24XlhU
evciLtsgXIgOCGrI0wkZmnvV0rcZC2Y8Qmj38CH8om9ELtyXbZd9ihiYSb2L
3LbHOrRaAbKgBwdPhKuD782KFV/9f45zqafvGg6KmRi4k8ZjzhJTLgPer2oL
fmybNdff2BOCvKEIC9q+lZHRnTcNplDcoBcKzS9sesdC8EQ258RtBfVsImnL
83gQC5ibGpx7D8jduj4b7OW8Hb6Tc73jZof1IpezKIws6B8jO2fIjvgOY0VC
M3nw9ZpxLR1iQlT52A54KqyUX7jTjFF/MAngPuTQX0B1sOHUpL8f23oPoEf7
ejO0wwvsmTh8Oh+kdzDXfhukqN5T7WpouAbBkMOf+XMTsaWwRCZ60Yh4+EPB
dihPYhg1Jz7s/rkxYVwvyhO6ATaClxsRVAzrW1WpQrIHVa+BnISQxyEfcaKX
tKY6nOsFvuu3myELNZiUXGJPKF24H9AqqfU4QgvYuWJyXoyQZEomZ5qINyG4
3iapw6uzR31QAtYNHs/p3LxnYQW7Eufz7jmCiYzwniCC09S6ZRtLb/f0S6od
QRwkz8S0zz3Xin3vdO9jldf63sKEPwTsLXqGenQ8XLO88topwLIWUUF5DfzO
lsH2yupqYq5FISemkeqA0yMzho3uaZuiuDy2BIfnUCE8LfxTgkzhhDQp9eWd
fequYHKpoDIiM4HRr9C0pAdjUxj+82tp45q6k6QBStlPpystainKOUo4zOQJ
ikc2gSyNQWunkWuNqPXYHPkFX51gFaq3gaAyGiDLNWL3DBm8giEmJ6OPXLyY
rtqUAOBcklmADMOWic7i94YZcRtQbwQpJvB3TOnC7tVqqcBYBlgkse/oLaEB
YrWhRc61G4RJ/PKuIYwN3Nx84MRT7nOArByhvd/J2xoqT4WKYpWb8kmTMTNX
wDjOymg/3McB681KgWQ+t/hpg2kC1Mbhm8J8RaIrBNQWyVs1jw7jIqRKpNDP
4fBXOlFUNg8/ve8cHCjLT9g4Vsvga737s/g/dxTh/2fQ3y4CJLQF0OIqCj2V
radEPNN24DrcIeFwtdNeDwfpBTIR8/QoXADSPxKOS7bVNiDwZ5QKybfKfYrk
PEH1cTCysJcqJWQVWKhFEY7hYrB9r8NC7dTmj734iIG90naZwnMCRMCMnrzj
jxE9jbN7yLmAMXU9rCJGK7pId3SSbNKmG4PSPzDAJN0ojaxU+uTJyWyBGOBR
IXETG9EwDoVQmA3N4C2cARLkK8GGgG7jcgx/scXk3W3+xFm7vrgO9zOOgvDM
KLOz8nDujBU8eRJpMDcr3R6UU/tqs+57oUdw+FnDNZjOyYf2LFT099W507wl
ZCYIv2GkG+sdAOghWKEhDLGAUidE2le/wY9oOstPsUS+sCeCAKZYO2+qhYwd
RubnQqo4J8gTbPLIk4wbaocveK5X6KQ6pVm7nH6ChjRfC6SpmJpRgDJgE91P
cUhoXSEUqd9edB/afOOVys20B1840LT5wYfwtaBD/METC9eJ874NTnARk/FX
OSE4ayWFxrUM0dstPq+wGtaIeFRnybHXAY4XeEpSyFl+h/+M09GaLAdvpmgr
VHoFus+xlE6y6E2/sgw05ICnrZDk4NCKey6yGXC1XQNpFeNu0RCkLkG9P5I4
8XuhTOeE0/R8+vGUYMBT+VCY71HFF+7fXWnlDdqAb2UyqAbYzFz74sCTyfZG
EgC8GprJSoSxM+v2qARK91MopMAvczREt4jY/JUkT5j5YXtHohj3hElSLCHQ
EKPuMuyHthx3g2VCtYh2nIq9URKwntnLw/mVxACGsmB6S6UT8olvTinqDo+i
o+06ahxONVBOnNbLtm6SkK3dk7KgBDedNzL+8gbdeKPPUCye5YTUrkrEgb5I
IwixR1eHT6Xe4+z7QtLzQViWfHXd5x/us0jK3SCOMwC46COyZ0SZWkORV1HR
lgac/fPFJldWdyCgpFzVCAH7+ed/WZKKLyCI6NBgrO02aUhwJhSZN6TR1VTS
oBZg6lH3N6XAts291qWXxd0ey+Rpbcdhy/LhOsLn6V4H5EEh/sDi1W+j4yXF
UNk7LZ1VvdNZVB4yxlg+xOe4i03XKUc6zA9R7h3+pM5XcwH4+MHEyd9Prpmt
FBxM3JYUJfLxR+ijRlbkmBeGSt5x8EZuF4NsacldKvAsmFReOZbO6w9pk+n3
SBiFoxpbMLwL02lU2QMOFQh6J9xTHVE3qZV0ayDOT/Gr1F0GC6gtHQKgAeDO
9d7rtVCemj+Y74qt51sgmXaAZWsY/xHLsDSYR8f6+XcqQUkImssxZxrdbQ/r
0WuGqgUY8cd4nrXyON9+EGjsQSvtw+G3a9ZTAZenLkRuKz9/upuVLvOzl2tc
YWa+GMSzl7Bl3DGNlErjMbYTkX6PM97yNAjUuBVp9PJCRh4n6GNxW0YNQd2d
jxtFLRC1IrkwS0P/wFR76hDKcPxqdPLoKLOZ5ccYO7S4PQXT2p9rNFQnikZI
5Lfx5jSXhu2XZzz+TldO6pa63vOClzIpnMk6jX9Kr6JtJ8qljEY9g4UMhzIM
KHS39vq4knHxHGkGUvDOeptyKBVRbXzk18JvkBaMD8rOGYi7+jaNhkE0QJtD
S5dvKTc4713Ejko0SRstGHcEZ/acxwmOD1Ca7HlLhxcbwxbe1bDhWyBkgDXp
GmEpFPuI1T1Ec5Fj1C6vWAwmm7+24b6+UzAm+Wu+JhgIfPmqjy0f/3oWDfq8
ZlFMZxFEtDsTTESUh1f41NhFsNJspEY8IrnuGS6N7ad39Fp8Ur9X5LZlX/PK
5j/1ny6lFMiQj6AL3Hcr2btOkkeV6ZmiehTZjIHwNa7xH9Bx6OIJgnRBZy3n
3JJdxhlGW5VGH5T/oa3mAfeFxAC99POWASOtcji4McUVoTXKD1Sg7l1+5hVB
weRrTUij9dGynx+jbnAuK+OI7jKxb8pEKmyN43HjfdeDk7yVZDW4DRZ4kk8/
gUDFbdUhogPvGZJ6vgYzZZQ/C/Gdd9pyIp1NawpImPV041zHiBNwuC3o61Cc
ZSBml/ei1baqmFTGsr/3jxJ7HJhXzBWCX7/LQqggL7UC1LF4HD6kGR7O8Vbt
fk9XTCTPn82CW92RdQgra5paE/Z2/X2jj3KwQu0uFo+RqLlK/xxCOkUSuGG7
y7xK1htLCa46EnqVWXowtIUAV43yYIMgI1FCznIm6dCayedTuauSYuKdhZXX
gThnIx56qBMx/Z+ElIa9sC2biQpTT3VRmP7NLrhW+DCiUs97cQ/9f1qtO9fE
IIOYTYZe1F88O66kyLl7YcekWVCUtXnGGfsImAujjA39f5lYsMft6NgPUhLt
QpfFTAh3qk3bKvvBQ/kDUUMl4O+GEmL1z5++idehhoMggvB4HB+v8AGPK1cQ
nktnaowpA6RUJso2Q2KBE2D68jdzm3mLKugmRpDDyWAPr5w6hqJn6RXCYCn4
Muio94rkJvYiC+dH4956PRJWTyNCX7v4hE3nCk/g0NnKVLSyKmaBp3u8Bkso
yM0CHww/5pUBDOw4wMqPJp/eufaiY7v0fZx58rSkCunDxjqxBOps0xx7yJrw
uflPKKqcVIu3nzLJJqrsU+tTNbf47TiYtpzpPskGOzJxsdpAz6w4imh6QzeL
345TOEAi1ywjGW395GvQCifOZeRzYJqT8A+ByMlpJnJi+b79+VT18NWXQCSs
Vo7WCKIE+CJ66dQ/kot1AXtFu6z7AHLib3ESKrZf2IlWZuUlXOyiY6tzjFxt
xLKt2EDAnN/iNMX7gOePMM4c+jVTEKFKi8F1KH1fcyvO3Q/gRPdo+5u+CbEi
P55NrENmTP/VZWgar5EZxORmKEf45TUDfxvkH5wv33GnV8fLIg5dDxbXbK1C
qFg1iAgol35Jq5nVixc/PLEh3r7jUGL6x18MqJjGuimTfO3xuAQIqbnhKGpY
c5XzZ76n4jxyyL590D5+GVq4sj6f42rPg4YSB6X0TWegwxaiB984joIxtFtE
MdtBtQTmItH5ZULmxihzBO5vFovaz841yvnbOmbb9ojPlbGCBgc0PbuSHlIc
1KqVrO+lDWS2cw83c7NWvkYLu0+vvahBshO2vFox7z1n9ZRaqlVxKIG91T6j
bnfcq7hwZQGHUviTIyw+lZ2GXz3TvFx0iz3QCeYXXRhNha3/oAqmBncSzd5n
9sV0sEkmnFAgUnxwfPz0ba511Y96TEDOPz4A6769p2MDvyvYAe844lcuUTMb
ZYXqSKR3dDe0V8Z37TBWuC5YBph36/Zsc4wv5zVyNuxHyn0bmU4vgrmrSm4o
Gu+XM6m6owpVBYwqD7UtceQCQ07GoZhAAXI3l193cOMC9B1SgNmO1dQ8SJyI
P9+Ni/CZDg7uS0B7gSTFhrCjuWxTkTWKbni543iOHdDlXl75QIdm9FkFge04
yUp9m00PDtuOylvzvanEsk7+0oHJDGW1o9friy4E64b8s1n2CaOCXz9iq/za
wz+W9IwiOIsvUhfnUo6TUMJuhULe8jAbU1nzXN0lCMTYjg/g0AQz8kRMDJwq
/0FrNQFFiOAQkWkPbqe1naxLigUf8w5BsHYJ74Gapo0rD72+7MIz/zNUIdlR
Ze7ze7c/G+4SANja40orWuqUfLGmivDt8iZP3EYTLjWYKhuDiYl/pzZf4Fq6
YQa8kZPD7tvDqzW6pi3N0EwkdsHS/wmGk3NABtRPV4u/uMvWzhZTg3GvJF0M
dS0seArS+d0MeQEiKRAJEjCDQ2BfqQ9vTyUw0FXAc4MSvxc01j9jAgz1p3Aq
AlpdRc7ngv9d+2apTYJEbNNGUfKV8ULUDTwuRCpo2GxJ/8fsh3MmZ6EF/tN0
YTrfx+N2gMCLnrthyQ5B3CFPwRVhCVAe79AbKqbUecGXMHwIyJ233v7g56eO
1du52x04ZEw5+uQ+FDK5HB1s/qlpYsfuNvytiV7cDPeUSsDJqYMPlbYtKH5Q
xHr8/MQNQGvCP6Vc0mICNK1RdZK/EtMZ61lgqaxrOig86wENoY9PHsXOTabM
C1BTVSoloDcajn4DTj9Y/GrGNLFnhiihMvrqpUjA0ZwM6anvqlfI30HYPFzx
aSHouNyZ8ylqRtdStMdbodidG3StuBEdmcbCZeKgTv54kVSKTfCOHB1vUelw
P83ZsCYnHm52hC6WcLdULpawGxUnazRzgVqVq+Me+YRFfpt/ORKQw/c7DaA+
X6mrczb/PmuHmT/xEDm4gnuqPgIc+XkzFeTUlX5ewGJijwJM9+9eu0t0mDL2
58M+7PlunyBDeBM8WKt/Er826UVZ7fs6BILYypqY7th0V/NNNk1ck8lpRCG5
TbCqdjzD1HRBnA64HJzmQnXYuvQTpxTP2Js4n6Z4j2Ro6Ph8KLFioAL85Hmj
OV3RZqiMGm4XZu648TiSD6Q1Lt6UlJxyz685Kl9Mt5V88aVbRvF3kGuQdoHX
A62fAgK8aakjfrAQUARvHHgbKTqQp0jRsFmn50sIn5cRUqs2FUOOWzZnaPtZ
zq0957gxAPGp1OseTEWY5oBpG/+0gmFpopgn1q/TcrPCfcMowZZDrljeSe4z
+Mg90NFqvU06a7VPGQspWcs2CfXWT/BAPeQkd5U2ePvFTHKahi9O+oZJ+Wyd
f8hMzBsB3FOHQWFkI8BsD2zWi1tuaaXhM7nKH0T2junkmrMSqkwoZI0Pk4Cy
h16byVmJm6E4cyLrFR1tnyn9i7iVt8Sbx0W9u/m93rngZriN6TzKdsQvVx/b
X0uP99eupI6yTICYWXUIhBbg2m53/ElhhzgDtKrHNycH/ebaqd8bNzAV9KTu
qj77VJQDrXMVku0SZ3vSMuzsQLZArphqfeUS5EP4HZbm4nHqL+oZCjPeg/te
EzlN9PHZERJxq+j97JZFIqoT3dNaJU7qpOAxWE40QufE7qRUKPCcUNqkzrkH
WrUmd9m/l0Pm+QuVoVlW/JPwEfX8ze48D2y0FOW1sE45Y2nlBc+lNEvsEn4L
4UqzSOwNIXGLl9CSdhqlE7Nm6CeN3B4Ku9B0kdA+BHBIcnHToC+wrCh0Sbcz
xLW62DM36wLdrPhni6mFSjFe9s8TA2Y33OQUdyz7ulg7neY9biVFp+IO2s+K
QHaZiA/T+BulHTPMAwLuOBXR4STEsfqdw6y8UOPkvMoM2so5cS1wz/TFMAMJ
hGqVbOGfkYBPddgQBL+DVXE4jFSHTQ0kcnmz3HVGpa+qByIM4sDlKY3ERjEC
/v/I5O95fzvM1tGA+oxGtjnlpcROrAvkJKxtu1y/DHTgGNjCWXdQjq+4kBJx
IFjOZL1XuWOgwFz56gnaDKzqIgNyhF152XmrKniHCJq57NEEim7OvmnZxl/q
hDrhJ7VgMzy3WkZA0IE5mJHh5G4JjMee3u8wgsXXv2fVyTbG0FtiRGeQClZu
kejFnwuoEjyAb3Bf2j18mjmbNAU3LgX+qZ4uLCA93bTWdVDEUPn0eNvftKuy
5qe7335xlY9Azb8jgZrJ565WoN5F3/PXziaZvAm95qqlDGqQ+WN2GkWbe6Wa
TiwsuutGKAsCvqCIJtFLqSzIs8jQcolDrs4VIhP0+LDkO1yOSj9M2RuCUfQm
gDSc8kpGj6B9oNXKtdX65Gf474fcV9br+af71C65+W14f5vCjt1Tq6h7d9Mf
tn0eqZYAzEEzzFaS1NaLG0TOdEioPc8N9P//WEVxWS+ClK7iN/H8fcyRYjVl
BFqq5UOSrGdSN7VxnrvINye13wfEppkqx5t7qzxTJOc/gQd5uoH9BYy3aIef
L0kf9GDiPemBcVIUmqv1FmwtlA3tYF1JpzDvz5PliGGYnk0nad4ePuiUBDEF
i1FvwGB7OJ/mJ2HEGujflFFhGg+9rixkpvvz/BRuePPDkdCiGFz3hMI9w/g2
gVHfS5/riMAHsiihc4gDqGK4NyCe6mVbZkNJij1m8u+F9Yp/TDzlH6n1vNQM
EPMctOapoCy0amCtrYoDbtm7LMKsReZ/PH61Z6rhpfmCsXgJ6OAzu1MFQjk3
Rj5oEbMHUkpCiQqW1K/uGs+TOK+S+IsOWiTTmaz4CYe8GW+6FrrGYWLqZGcu
HpKARHVP31XdlnV6ZDHVDx4c8fswm3odM7xsPeEZ8jNHVwa/AbjKXiysy5of
NI3HRblWhRb0jnUDmxOxGvykHdkD1heThOjdl9Jj0L+f8H6TWUU3M5S4JiIA
cW08AU06xINDLThgXOUi3LNN/BOGyK4ozvoINu4i4ZeUo7DulJVNoCL+yAyG
No7lEFCE7IAso6vEcYIcMuAkkY2YAjUpD12XodzA4PfRR/ZDHBjygYnqERZc
CYH1YGHu7PZ/2S6E1ByNZMUiVm5K7xdgmWoIspxgrFK2VVMag28ZR3/AUXRa
E7xuZPy5bs0FiR08+XyAKaV430CxT59VhiIobqbH9GCOC4VxleTHJUg+IZOR
T1fA5wNEj5DdwWVso7wlRoXgPl1i+kRSM2AoZWCkEbLGY6el9I0EyTOq6I8G
16oLmGp4LAkBsZJG4t7PrQDSs9df16QgCBgkXjzum0YfuuzGiDp0IZFSbUNv
xwss1BvYUS0pvrGBhOSmP0whRccwUGBCytRE1YHpY3yOt/0Hqi7oBzoAqkI6
W7r1FJPhL6Y7+/seDfSIBQ2Ri6Z9N9DAJBVb8uJH3gHW9Fi2Tp3N2TPDkz00
2mfeTNmhK06AtPGt8EkCqBJpzp/X7mJ5ewYrgdLzGnD8i4DaHWHeULA6B19h
f8ERt+KJUgp6R5Gfsgq0WyAbRfemwFwF9HtPjFINKp4RRyVpZ0jASjQusxCx
xUYFRUuUrBJxaS8H1iEuUV0lK9LUEzx5tn+WGD6U9FL5EKRNE/c0UJM8lD54
fXX2jMI3DdNSodS6umm1oqP4c8GAv+W5Kl907QguiuDSr4imp0C/2rhspkRu
fqayA5jxZZ6ecLPnAEqOkfaDa7hwJSVYoIgiV90OrclmOSfeoUIkgcHTMW4s
at2zYqKgProW4fgF8LkKwC5hZxoAjf/RaAEYR1EtHriWxzd2fQ38RmgdZFlM
TMXd+KN3MzTgVbEhwONxWNWjEJxIoXkgV0gL5czTIahnnzy530MlC2UB7D7z
JPtNpS7kiew+Gz65w7bodOXWLG1yL1qVmg+50Gbzd+biIr2GZPV92DNDauJZ
VCXHisMlVhMDx1Zqsn4ginQwMioJggt+awsLdG1pCJMwW1KbPh/YF6ZHa/V5
dQ7n9RougH37DNiJXe2o08yvRgfRYNIMs6oaZaY+kPg1OmF4VO6wLCxS4KSk
ylNpLadCyGjC8ZKIKBfVrBRLX6aFat5oHo/+Rc2CDejuiPXHTFpRgteUCN38
olkM/aEikNuaFLxmRChmqZXjPqgWLRLF5WRUNUP+Zaj2DsSXxKuV2XY7wBYF
4lMWlWdbRvcVEPNN7SvtqwEp9CGll1YtuPWwo96GPVXAxRX0ntyeF7XHdxAo
MVzWoxvuDuDU3sJl6DXiOC+Jo9iLBCqLRWVhYvoPu03VteKGYOkaPxhcs1hH
uAsJyogGfQo7URR0QRvx/HM91vZ0Rx7iNyC9hp83d9oOx4PYHHOpnbuqIK0w
vQ4bFlyjA4vVh+3CB3D6hduk1pYekImg+xxBiFwUl4BLtMHZ6uAcDTZ6IH2l
NhxgR8qUD7RAW5zCCmTD/5fyHPaGufE1pMepOz6uNHIRIjSY/Wo0b69Eh/jF
VYdL0cw+298BJ7rle7H2mb2tWwZfvwthgvclmd9q4nXmRf8sq1SqV9PcSEP+
anATtyPRolIeq6VJhTBhdZTuPpRwLiRz/YlQyW4o7z+E5cpVv+F4uIt2weLk
RDW+GAfkF8nJoK+AQYM6oBRrMxykgghCJrhEf6BTWGV2ANIij6VcMIxA7/s0
r604h59i0FO3i+bvhp6VJXXN/k5bWt0BSpD2jnGDpOKu9vxTlDZ331EfX2lk
zgr04/sfvTKZ7Eyx1OAeMjRqMZOZL/+jzTgVJOqE5Ck84TEApFR1b7lJb16N
cJf2NVsbCpBtdhAUEJxfswBG6lwK84RL2j2ZKPeRe0eyTzEad49BDwFPuJZi
/eSr66wODTPYI7mHUyEdfdTx6Rk/sLdzGktfZlEIc/OThmfEEB+F4cvI2zbK
r87OR8IQ8a0DMeZNfHw6ihkCH6PgOFdM17FAWC3adspmzzpXokZhQiNWk2BP
r1QlORZrvq41hN+WMP/QEI0dVK91twHFTNEL8v8P/AbluVLzhtNzXaFDce49
bd8YH9BxOU4OugoneTPvyfEPnXYG+Xokvj1ZTwdfPxuR3fRPmu15lHWYfe5D
fdc+6D3+TJQaUuZEXZ1SvzpnN0oMuEhrQ4hM996viXy4OnuO+9zHbgS6jX/g
3fIPlekz/tBJkBcWPd6ryigmrnsotvQapmBOjGq2HDQaGaCHnRK8nOiXwF2L
arArJzyFTcCVIhvAoSqH44zxM24aSll+9jfRMrzJtij2c+56XD4q3vpUI9fG
KSBCUaV2kGThLhAoOAedNk69VB2sg0QxPe6MEKjjZWsOmHYzCda1Ktov7LhA
0jJ1A3U/BxNthDSHBoBAFuIkZwH3UTLP3GWNDEiEyzI3vZQl3me1HiGyfxG0
tV78yA07JrXCSpY3nisxltIIQQaC4esyq0mR3XrFQ2X9qLgQHSvSh3o2JJop
JXRwrJ+UitX8vzqmIVR9soXvJBLiKlAbF7Lttp/Fen/simvy0Xq0ONgUDeTZ
8rd/fIT1SA44ZgXoyOechkOd7aiLUyiY1IZoJnovChAGrd26EQopoABJo1I9
naPwyFbS0BSNfzMeezmR77BCO0Aos6MAPxqBgy4iiYnUBVNXgKJNQ1H7GJjo
fxMvNTNubmJr5vukoE05sWPFmQuDHzNW4a9UNr/Qix1w1k8Cou2BT3wYOVqn
+Tud1tWrdY4EsaYm8e3s+gN7Ox/PfxOISsX//AosKomM/J+8RvjSnWBFq9Px
KuWf0KNBNMNDD6b5nJNDEIqkGg6Sgf5i3lq4Tp0n9mfHNTLjkOsEso9Ry5An
5PKUVejt0NpYnftNip/OruCQMqk0HDsR5XLRqgY+H+EkVr0AuzVWC5bn21JA
f0hJB4eApQg123mXcaGl6QfavzWiO4wvQXEuedF+3Q47b6yGrwJ/OJ+oOsHl
BeZuQJdeagnVrFw3AZefCYplS4EEKVQbe9zh4yEfZcW99RPxGr0ny89RNdY4
4aKXR19r0YnLfecuJ7binOZjKREhRx6YAOXBKoSfz98s/IzQlKxubmegp8fP
fQLUz+v6CaHfQhTdD99GmvrcReCkG5Ur0TMQEsW6z0yYyybYnefjSCMEjWXm
c0WZ8Ozlp53E0HsO0Og3n+cFTtT3cQw1B04c0Bi9fdlDYz2Gnf1iib+qUJUr
zOm/YtxTtmIS/Z9RV8xiHMClPyA2HF77UN0BhjElEI74IXbsCSaM0FL30ZpK
18bTTjKK0i09mtaye1k2zorx2eTaBvIgdPW/syUK3T32K0bisP4TIPTFgHjJ
QwbXGNQDgFVOYKcD028rH9UgNK7Wq+i3IL21HlRNcmb8ETj4WH0ByYxErRoH
qLwD99Y88AOwx54arAHBRUYrbTI0anYvZ001EEoOII4DGkajS2qryI+zCAXt
5h8u44/vjUIUx2uoZ/d1XEBBzDU1743+hyCK0E9PDeaqr9FpOkQDoJWJetaM
d0Hm/JV6T81e62KPEhO4DxlFnvzkNkWBokCG/uCR/9k6sn/oz38wTLh0bGf7
QxTTrWmMwqvCNAbPZAKj7ebuAL67QPL5pxiGI5SYfSvT6+tLnoikuLHo4Uta
Wjmp+LPi53qRVvpI9ptX7qKlUyRgcZeLv2x2qSN6xLHmW4erqvO23ZMwfiGJ
h6ND5ke6Wmk2ZjOKKob+yWp6G1YVawliX063a1kIVZdzh8PEx/ShkeaxNTvA
G9E3E/xtVR1gW+/wbBNID7BTfQF5hxJwLBzZrcfVF3F/sdnSmYgNhJQNCkJV
NXgPD4L+GvHBHrwoHzYfJmnMjqvD8lAWmbZq1o/1/Bx7wP7xh/LKjloPxSYD
Kjw5Uwg7Tdy+0c36CrtGbnczKvmfb2X8KAkN1WsVIXMPYvd+7TZLdczJpCpL
ljQ6bNam4Z93o6f5zP6NrwNPDVnm87mBH+jer1xtgOxF/CuhTo71/c4sos5R
RvOUDB9ZxvlbfGWN1Xo+Ivms+E4xS18ykGrAvDEr9NO92WFx8rKPFsYS4FaT
KnXuIpOFJU7ye50lNlCUhQju+or55wKI0M3mlkPqJCgHuFTqvMcRpj+saMUn
363WGyRs9IhEK0VSn2frO+o8DVFOmt3F3Ha1f8mBXZ7LY/rHCWyV01pszPmt
9ZC3xpI62OVIqfR7KvKGV+MtJPvo/vUXk/SBQi19w+nlMOVyWGQEfquZAQA6
Xbn54oFNlcfYw2JECiM/YexuNUnn0gXjjgp/ERZessa5TfXrGKp2vdAKFlM8
3pfnt1cwS5q59mfOrqIoAuavevN9ynf7IHeMN6rRDuEFz6bbpxtThfpF+gff
GtXreZ3QymelN2Wy89T80xGLftOOMJbo9HhGdt8ykgvqHC3C8yzHrGHeqdy0
wyffjS2QuE+9JYo/f/0Bo37nfyKzMYz0Zge/HbVSVl0O70fkabBYmZzdzMOD
e+g0kif32kNbFl6rDyiOBkgWhpvv9AQcs0YCiRk6bAi7u2FwUWtTsmU9Tz8x
paf7dqrsL5ohG24Sd7/DFiunMnjFhbHDLM1odkAt1IoMBdFBhctuuwBc1GX8
//2O5xQBE2eCJDXTJV5GVfTuYKHR1X1D/FQL/7WfjP8U552Z4qOAJJ8S9zoL
KNIRTzD0BQsDLejQYIvJjsJ1noTp3Ex6KmVrLVr6PhM7dK5NsrlAekMun08Y
s4f0usjivXFgUxxaYNSaaFzAbaFPKkfta6L31GYWz+bEOG9PkmPjPA60eyHv
Tq9nAX0Y1ZqtAgbGlOHxitQVZVvFR9ff+bTVustojejnonSTRxO+fnGY+GiQ
zCJDdOrlCdpv1lqclbwAFTVtIvwJ12izsX0mjD/ivVQNijPJxQ5bNq8AyJYY
ERF3aPbF9y58p2omHMEOw7IQP9XsYlr8O7/bw0hAk+uGTnjr3acKE1qgsvbF
z6pFA3Gg34X6dL1luN7MAU4nv6zaxE1EUgB5riPK2/3eahslDXbdsTfB35iq
eppgWcvooWhDGNAgNkSSmegSrCcy/H+8sGaiyq/5sle5f4sya51UmO6ShJQK
6yvYkxOt6/IGe9PYPnZvrNJhEqxeQXKtX8bMVrO64P5e3Ak/FH+9XDUsr/t3
fjPGRvjzwCsCD6NXMgG6S3SlUZxCeuG1iCDZILMTPQ13QitoTuhhgDx8c3c2
59eMXa5XspWhk0pzC+uuKVYx91S2A5AxqxUWVVZyc+MEYczYC1Hn+UUbvS6g
h+s04jSpwxC8XOZ3Q1tFhK+vRKA0dVWFsHsLPWFKFQyxD70W4RgDDdc+VK1k
de4XnKLMUAPQRK4l5KESxNtd5s8+6I3XOEBAIytBPjU6wJU1UkLE+lTUBdh3
mqeQQ67mwiLKLyyaQduKjFe5K6Vs5BlnxY4orplck4gtPg9Z2F5nA81Dk2J7
RMiLDJDfPfC6u6h6V8L/cpkmZCUs2KSzeZjVWApyeE0ryXPw40F5kBEk7sbn
EJi5bPc7LQJp0lukEv5JW3yg6lJz1N89tKf7IceSGEt9LWkl3YU/2Dpk7Pej
6cQEDOu8pG+MPExvViNpEL77Q5RRqrrywmd9+2MNXeXBQlXdC8GCS2w9rjS9
tuqEKOg1Tpw5yXUExNaZmuG5/BH2EEjxLyLsS8/KhhwnV01a9iDjTW28O1Wn
lR2GXNTw4Hq2Jv3U8kKc76HNKE3ds/c3u8+Exw9Eh+Mbm3kEyHZoiceTOBzX
ASPBxQeUW/mFrHLlZOni5/fGiXdNmpM+7CPCDA2kOIjEJJdXPUU/WaNAD7L4
BdY/sRVXKZIH+L3naJIf95SXi2XkadYrlak9qgDfGfS1qEy9RMak+FolJfYl
M7jz4o3ZebHIeCI0QXTJ8NkGbVGsCByWBC5A2Y5fZQdGRDgod/jE7sG3B5eQ
cRlzup4j4789RCSqEgzkbYm/iVpVTqNBwq3a5tkAbwcrCx0fqsJ1KS+GzpBw
ewGAppNOU4mAh70Ix310yh3vDwvutWKulNWyYpF6KT56EoleXaGu2MyuHZJJ
EcoUk47FB6nmADaFAnp6LFgCvDtYOmpL4tIK0eC9Bh8SQmgvLAqXOEE4h4oV
mqr5QL0y5JAKqNAMYtztZxORKX1ptr0GiBjKqW/lhWgCWIiVtBrtILeAJHkd
Ez2ZlGrXtmbRaaihaOjUZygMEAhT18vPebEwRA/vH9+K/y+rHWxl3GMxr3Va
FokjLtYgGSlFjXuP2AEsmIzSsaPCuiPGOPgVjC6UBZUoHQFy9M/cTNDIHvlv
TZU/oY14tVPIfEs9hd7Cd4q8NB1/Aunc6SskxlgaNgLiGV0oh29WTi+o1XzY
EkdbG9yNbUlXnDx2gYj3JVMpxBvXToHLCJni1YkLgUnLzYy0+39aaGbhmV7j
Kuzj872m7qeel8N/HvUlvMNSloDe5W9/H7dztdkRD8HFha4frc0wq11QOrKU
KjnZiCgfsgFyap1MsCUeSJxuDAI6/dj2WqYPczBvVACSES1++rGCWPc80NYu
Y4RBZoIoeSSXLA4Zu7KTPqe6J5FVsbzYSq3zo8LGkIcIgbE19SHYX6X4PX/p
EN28hrrUdAEdJTn1siSL0dgIh172sYr65AbZyUK4POfGf8L1Ph5tdebqKWiC
zEoK5Vjvl4dAvwcE+3RmEKcd1Ad/TNgU+700SVLD+O0rHTXp2nCJbHAlFGNS
vjouXYFmALoXnG1SyQOpJQrD6a+CZlLX51lmXAca8y80hm7MFoS4GIEq/xgQ
i3v9weU5Qj4+XQ5LpDnXNlqPI1fjPWS9XTrChiunSYujisxcjdF8QSNCc5US
W5VJJrVfHAZbaS2o3kB+be1mpvre8uijtCmNVKeKdnSIG32o8XAGYwFeyNpa
CrH+3HYBld+OptlEJpA97UJPagsq1m3Auv+wzdyuHRpyCh8KyScrWEaJErvn
GjX/26+nqIVFLP0GAZu99j3pzmTy7qhGCYdkB7fjXM/cNzT0XF5CTkNddBtd
GaQk5cSRq2rELDMHR8G84EC2gS/RcYRuc4W/IMFtb/IkVZFhfVNUbiUgu913
bMtgWlNvMA+W4Ym+Ovzom9ckLLmwuOVpZ6f1jCo5UmAnES6p/LlDUf20PSTa
6H6QZ/fA8u7kc763JoMj7IBofRTWQhx1BLvZBdy63mRek+u821b2EXlkVrFG
6MLGN68imQpVYCJ6jWyMJwo+7LndYMWq8ffVPfWG4dFQ0BHmbObbKtnGdvTZ
U6GNyFkeLm3+NwYjn9StzaLBNAZZ500yvqWMjFrM12hS5HBs4evJ8OvwqLmi
9TEgDmwgfcMCJrotcEmslxlsN4tLvOJKU5hq35I7zIR7L3tHrggsgsv5E2AV
DjrfFUXtV82IeHR3nSUsnjInL0Kp1NnbaV66LfkQSGJQJlryE1aqDV0bbjyI
99bacu948Bhrt/9et0tBDKV5nk4Wslr5O9xraGyi1U8ykss5gvB8mTB/7N+s
kjROKlqUvX1oe2kKbk62TzaEY2x+k9xMY4Z71vzXwmgvLnNUrsfXrlu3He44
befVnk8mhnmhrQpofvffhpiJkDD0LT/IMUS0Q79w2NWDwTRj48kPBqt0fwvl
5WhEjM0VOdSo9Mct58GCe0DTx2b9jrlvCoew0Q3sOXrcIqduxl25CpDQd6WQ
/Fmd7Yc9ZcSFwdiKIYU8NxgvObWQBFjNNOekl6XFqIkLXlJ57a27yamzyMCm
JL+dRjy8ErufT7wXyWzd7RljwhuZgxHFWdlvWkY5LPVWfXqCcFiIrpy4HI9t
PpY1U8IZ+YjHaIL/aa4Qxf8ASQ1VfdPgwRp2LvgLOOoXgOoZrOo1A0sHxB9I
+YhHjM8yrXCbeIPBpSDKVq/g6Lwl4ihM2jpk9+ZoLE6Pyca6xcL3UvZAxlty
typaCTVlVFw+GUqYKeWC+L8OQZbcUxXB6PcZxKeSUhysJUFCBJbJic8X3Pl2
RyeYrXdYjDIS5FemACVlTMAKrXog3Q2nI5NZwgCto2D6LC2QGASvbvyX5jNv
ATS2zTxDXy8VPukaZ9kSPlKKLvKKelnaQRiEeowe58Dmywd/PzpugnV8GCaN
HuOA2YcioxbuHViciIOv0NzAL7VI9pIJ4+lSZPCzuJus+nr/Niw9DeD7Hd8p
82AuVwwngks3eh5TjXHHK2HPn17cR0ICyVtwPI7PIM10JxdR9mBlAbwSYDSD
FOdSCXPFi1tvVBpOK24wHo1WYiHHaA/w8YFLWtZavcRWOYX5Sf+OTok+QX/U
lwQpyzW9VJn8/t0sQ4+mds+Ewm3ob6vIQwXcQwq8YHl7+w8ahYNc1AaE8BkI
AsH38qrv0brudvT897vlR8gm4XUQVFWNbdZGYCGUF9AQ5Sc2zPvT4YCn0vh4
Q5ZcmO7TKmY0Os9LUi9fvBnShC2Y7C5NGYFCKvJc/0HU8tUphDqdnQSSbq0X
OEULdhwBY8hZA3T3rfD+YiMCU14zq6DALvKrncIz9wRp9U9+3zbAEl9kgBhn
3xFFo7aUw71jwqn7cBdAgRuMwOlW1EZCktRc2dlxk8wqlEk8SU4DJHxI5KGI
yMLkyWkx8BdihlKCQZAdStXKEa5D7aJWgV/ZOf9gC/UuOUJuiyOefa/gpGtV
qPvhl1/1+CS/0f3AQ5ctfhD2WZnvGa+jjl2lODF+oxkqq6RKRwIH4GSBRjUW
UDyuVTDCF6TezPnpS9+o7MiT16pD3Jh1kz6WtxOrmQBJPEv3WBSd1HPmWLHC
tpAkBG/k5pwcwgpyw7tjUkb+2SKcQU8XeFDvedFWE/apnr/6avg+kXOjnN06
wTNff2ClPkWlum6evY3SEhRnh696IjvJsAeL6oL9fM6XbazMIn2EWwjYLpp6
NURpONkJmhy0hMbIwObpAHFEqGV6OVHlypkdGYNGY0K7Q4MPeVH4Fd9UK/48
GqV7eWBmXulJcmMwnHcOTF81j0TqCGuBPJX06NmEG9WbWp+XNYUzykFntSG4
DoKToGkDPV93Hc/FgTYPeEm0MGuuLYDwsoJLBolv6hGrfvyNBfbC+EzOWGoB
d96+LM0ll4MLPFUx+u1tpR3Fp3ZS80QI54aRJAEsQ3zP8U+m1lx4bKm/jRWX
Sp5CO7pNc78riecMFOHP93GcdIv+v7dH4801JMcmSn68xl6gaqZg+XjSOBTM
ZUTRxyP4VlzpNilgecDnhUb1PfMw9ZINzdv/Gboh+cSMRuK//ZFW7nZG0oiH
0UHDfLuI9qr/syN/QGr8YcBd1hKJHg35LTvUUD2/XNyx3u04wW7UsTazNVAY
2ymN446z/7v6gop81H5NgJbX55f3FnfWmP4J+StWuKyHJpd2GSobdVpp29lC
JDU6SHHWt/AlvAk9x/rv/1MixEdaxiW+7CMUQTeeZvc50y6RHg0R+98bXf8x
CY2gFUAI/KCBzSEohxat9plNE98+55nOAdJlb1R6XyczgHr8zmjzKZTNIdRw
+FUFj8xpOUQ/8jgMlRvp57QlLplDVMX1EKA/d6gitkuC7sbq6JEV3KD0hsbF
IlWDZIvhtvyRbUgNTcV+NRu/5KNr0GW8vLdFRbzKvi4hNjnT0BCTp+wIZo2X
nlNe7ByfiZCFsXXa2ZCivcWB7GTP3rsZjXOq7VcLmfO0JDlqLbuXEO7OVNXa
9cUtnohszC/zh4nGoA+o9OyhZwSHTT4jN5YupiCwGMJqMFqIUplvvyd+bE7I
gtMZLD4JR9mcMd2OuxgAHHUYxBKHJ6lkHO8BGiwza/un0TRRZ/T6EjHohCQb
99X5d7lawEQzG8pkhV9B1wcB4LKiXlvlg+aRfp6/mEQmgGpAJLxDLWDbUTUq
dyWBlHOtonb8wg1cAuu64XkTmJjJc+ekKYQIsfpYLzSz8pYnCr528cZoGuB0
GZSL8AwEf6RDXzCAX4cdgeoNEcEvy04Or5cwnUyuD/1V/FdkBSdK2N+4d3KG
DCEa4ohonLKkHMdqwXFWlG59NJh3bkUUHNiVn5eg4q2F8ow6pAnHYKEdX+YQ
edNB2etlqubjLCZlpXspcJzrWGfuJGfX6uIscsiqJtUyvJuefimBtv8+mTiO
oDOK3I5CbiRiNP3Cyo6hnGNJecJHcuQAa6bV1CkaNhTYcJGhBNXMVRdYaptd
Rv1nhxM4AlGJzxnRpccSbEAWXqsc2a8L/dw8dMxjRdp6JYSJ3xZG4363Hp5z
MEKkP6HujUsaprG4ZeJIGFytASed23rxp1ISMOrEvFQYRpPkpiRtk2oTpob7
DTm7hvDFWWPOWJeMd07FAl+mvqm5Wh0dpm5cb1p+l/TJRmygEITS631kgCgZ
VKJU8x0QgmB38uko5uCMotR1M5+4sriA4nU11aGA3fA/ltr4NBW+paIgJM+P
IJVwffbvvHUkQxlAo8W6J5uhsIykhnsqYzrBJl1UgBnAx7hQ5kyFtM7mRxPU
ExJ0O37zhaas6yjbzdg9/ncWuEQ7u9W4Wi+lQrK7l3uguBYpCsbXiafHB1tM
f6wXsq5pRylBu/Ihs78SrxGzsb1BDNbNJa/qw00euKwsIYoMEQH2siJW7oA0
TN5KTkoUk9QZj3mupNLQGwJDNISW6iYxL5BHxBEBSwtz9ATeVyv3WM9Q4H69
WDQTQLIqvPkbx5CmVPHzwZE6C7qVXkKqcWa73/wGajHMLlVnz433tiZE54zW
u3Dpmuz6u3Yb9ePJtse08Od2uIWVEewfzrmQyc1+O4DXeFqnCiLimww5Etzs
aG+xoujtvIhGGw11cwcp2y80qcSp4LQgTpggVXzzGtr9xJAp/a1VmuKzr4RV
p/DxcILnVuEq0K/bdpjFNbsLVyME7lbXnc99yaLeUxzWByHvZ46wYHbU+zQ0
HTmFMdzWnRHrPr4d5FEPyLWpCKsbv5iM5rDpNVzDP6RkkJNzQc3GK3c54wUm
/vueokxhWGWkFqkE0oibtHWEuTlbSTDFjRChXb6B2nj7qkNGLhqN6OiMloqt
H6ZpGG/5WNJpdTz7NlxcUp8KHqiA0Km8ZSWSH+WWEWE2Q+my6sZU127aFfjg
/K/mLZvsKlAjJWwz6bARbgwByc55UPZrMVJf/Wc8wJ4RHNWrE43AyHKLFhHo
owRSAjkVNo1KA+UxAsV4C2Cwa0gEhe7WuMxvuEfjYit+/7KFaInI4oI1KwPf
NLqAFIwwWeOEcHUsksbqgQ1+MN2Y28Ki5c39rx+OnreibTaESi+vwyZwhOoO
14ialoUKA5U29bytv9KgOVYzsYSc+mN5XgjwMZZMSW4+qpnwjJYSELHBa5Ti
/he3nw+MwzAoWgQ1a5lGWakbm0hFpKzOL2RzFiNl29T3BzFGYEuLGkN8yhuh
RArcPur6YpxvRhaTtpS3h17VNoFVx3/5iCFXXWB8njoeLnrDczZpbwqi5EGj
WOAdDmeBbkXhvxdGoAAFiy4TIKqafEsX1Xft4VA7k5UZfpdiEoCsyJJ9GNtR
b93mPg5qXHW5rFtf0Ih8n6D5Ftu+t4Hbwhl77/qtvBmWKivnUd2Bj7KSC81T
VNyukZqyp4Id/ZPvY/y7nUpkZhpdg87dgkaKTN2142nr3SKWxyf2sA0IB9fK
UGzRyxPHkrMarZtccnkAbD68WFltQwCL8wOY4yZJ9FglKwzWmSYMHx3o98xl
MTUCZklDnYXdO4tKBjAtaeb4848p8dlVhBaICO6WTj2UA+h2BGCd2vwFcYRK
qHpGpa9H877DsFx+jGMe0doCExGuWwdDgDJ7nRFy4JGwuSrybhTmPkGS3zvv
n5fvB7JVMlHUNFpXqqVYKkwl7S2NEZROs4xMiVadNtdE6WkHUsqWGzR8tOeF
KzRbb1G/oWFfcwfXs1DupXEeYaKcszVFj4/Ty+orCwJYCeMDI6GXBkYSvZMn
Y/CLbSXnxICNAwogTB6UJLhUc3yGN2ywgwrm1yUq1EiV1a9DH1+5Va6a1sbE
CAwhJO4kNPp8PgcEuQL011y1UEr9RXagAfbTZBmJyqiIPT6QMl9PY3bnxXYt
XAjjYxMGMMH9esLGuwo+Om+uJ1C+k6c6aZ5DWqSHuKiBjoq50IfiE+3zC3Ti
LrlAUv9EuDivo0LWl1LIpCKLnkdK1iV0ntQ9lXfq7gwxzxCI3S5sFGVD6LGs
D9iID1piCWGkrac4aS4OhBWjeWumEr+IdTXDk2fKsykOepT+w5Qvo+YuYs0x
pfbzmkT11BW9S9EDrk944uCH330nqXqYMZolSjjZu01XUO2C4G/FWEh/7X7l
bphrbSyGM8qCFagYUklxCGJDLxEZBQ+SWF3hdrzMmubgCzb2U/e7gkf1IVko
3I+9USKMNe4z7V4CYarvU+SctUCP+4QDejS4KEr8xzuYf0XiTzFMVzvcXqiO
0PbcNqJQOOEcSpuGBJ9ktpL35mkxzeAoRaspIP5HW+/HwqE68KNoYEfY9Vf7
M4AKl7UpPHVVLcjYjcWNJci1ydjufptbmA4xlSPnOSz5eCfemTF0rGrXHn0Z
Wt/WwUS94wElCLdsKecp58LQcpV/qo5B9J3KDeAkOkW/J67vQUCeF11AxJsN
f6RCDPXvN/nhta5Xo2jjs3vAfP6UnVP4HJWNH3mKgNSYK4q+XXuIxuJCe6D7
EDGZ167+cAIzv+UdNvMEH5wjVR0+0FqBceyBTvpTr4VAsVbiOU/3lcfKS/EB
g0PctQgIhk68ChQ7ST22YUS+atXsNHZZMzQjT16ttaBj4bdwmxiW6EaYhwHj
x5H4WSrPtiXTuyU6lr+/4FWgzxdzCB42bCL5rrVlpMVUvcjhxsSMc0HSffGP
vxywtuNkxrD25/n9tSulbW5Fxt4Ffx6R9njPRWnsuQrqRWD5wsM/Chcc45Dq
hn6AB0kgtv4hqLdof2KMxzuPK9M4EmJg/YFN1PE/9jgNJPCStUkTIyAzXsYz
q6b82ASKEm0We4NUgg8DhH7izeb448t0QJYnTv0g/N5+t66RdvYEDi/d7QFP
2tjUm7k88M43CBM8BMQTpRYPgwBXfW5OYN87FKBJGm+TUsfn68ky5nmIO4Ru
vvKCtx7ZZb7Est28WTJboGofT116wXgZGZvW/sVxxmTpgViB9+mziX/BjGng
O+ditNC5qTd1xT/d/Bulv3jIbsCn0intPTKGE/6NHHq+z5MvsGfpGhK1uv+a
SvBwxu64xk7joi2NovUqL3wxDx55H50EHylBt8wGmwqXY/HhQbBWoBi7MBDS
xhHS/fQdUt/Oj5kyeiHBaZ6+/p4yakvfxWjO/aUVxJuWIYq5OBubvIxB1BeA
yMERfGS/U5d0JAue/CILNY421ESZI6zfrzUrfhxoZq6dyPhUS8/bCoqsape4
aWJJiuH7fS7zfXSyzor7soq+p2PlVWrutqhSdS3/oIDXptfRj5c9TzesUlvR
s0qOe7Ny84BnbcwK2Y3iO2pmXm2c2GtMd5F11wXYH3qxm4vyRdKIPSuFF7gE
rvr0WtDJ37P6uMbfqejcI17MUevYXh8N7u5+fuQhfP1PKZIjMlzp2o8QqUED
iQewaOkX8cMC5GeeV3ihNaZoaMEUdA3uAr+HYgW+y5MnynVvIVSu+COVWAQ9
tJ4xSwEtX+0byUL5M5+qQqCuPQbiZrS7l7Ou3E2bBX0n/IYILNDNMqbW4ktW
1KnLguppGoB9/1xbdXda55dGlvTbZrYz1j4kkXsTHXFA4PUj4z2ecvmnq/rH
QOUD7kY3GCWITttFons10EdFQICmLg5Qr9LG6BhFgJDqbsD44ZtjfdDHMp8l
H6pEfrDoYLSIt07DAgfnJghFvNNlNa1O7yYbyt22iwJtX/TyXhPZNa12h51v
dOzT+wX/aQ43fplQ0Z0/5gxoYyZNkmvYT4YLiiIpT9fkluSQA78w3rtjSWUv
34os3UWutlMKlv655ssZ9aIyFwXaslT4jfb1J1hkJ05NdLee5Y/XwPcX5gRo
xexQ7SmJeLJw55Ok8SJtFjlXFtu6AS1nw+gJLZTUTezCeLpVKkO96RUNJi7d
nFPCcmSzu1FD+Beh/mnu1rmrdyTntCajmPVpIs98K53EK9i+uXGv9OotF5u4
EJcIiKnc/SsczGzhGHEP3SJ1ZWRbY1ey1y8C112c/idvw5UyDwYYWET1688T
v4JALoJjcSGYOZMQ9qHFee940iP/af04/PgFAzj6nbYzScne3FNEToEhyP9r
mrzl6bS22WFTSIKNgxOyxiDxEvV5n4zfGAyCH23inKTRVlx6eL2JR/Weju+I
DAzteM/dbbI4CZrunjwqa8uEBI/9OqW5SBYfOO7nulCAPwsgY0K1YPSZRCGc
+0yC6ZKyjeTEY97OB0vbcXTXTufcDRdlHf/M140xHjjFzzRf8HuUykeW7g62
6TYdoC9+S32zDTI9+Mp2j9is+FK085S71IiL2OfEwKIFP1gU/HY56Vmiozhz
ybdbkosCZjcSTKXaBDgqkfhyIuFx9puhau9+5VKHxnoOW9r2mg+K9XvnKbzt
Tp/b5/W6jS3KvOXaLXIsSXa9Ec3Qf2Owc2yOnsbKODuK6aKKcxxmVgUxV1yl
xOuEA09s0LlOPdpVXwCWik4VPwcNY0OqS25qRGpVT42rfPJYEq5bfSFQPRP5
I23NW7tHYPmW5spMA2NNZnybhFilQw2cUgNrzCZmGGVEqI6SmM+sTYtP78KA
DyoD4sTHCqYo2VlnY45HXwJnQulQoC8rGhk0KcwSsYIOn41sXLAAQhtEdDtb
eTA54NxHZbk0g1b5mbR1kYkJPw0Yhc/WbRPUCYIo3/+Ned0/CejhlNgxqDQo
4YxlBu94jDboKbQCnIEwZpeyqC4s13l8B5E9fwHeSUTKNO07HxGaNEj1YWu/
WL0ZPhc7KHgwdboyRebxh7DovuZCCM7tU51kD4sjYBrRM7AhA5AjGmSkQmwd
qEckFUw+ujVu1rainCjudHdcK48vIvYpHnTPTv3DBA0pQpAE37OymRfBFjGD
vKAA6p6X//b1elAPB3O7pFHl9mALBp10n6xW9CEL8nqEOUwEd4vdPqFX+SdS
JMxxCdsGzgWmAnq0GOuJxu5ULJz/YX+IIgkVwItoM5MCklp5xEIIwU+SN4Og
SVPKOF1bnXfHtr3DIhqXOEXZTP6MnWpml06oB5+Xtm/nWtEinCbYeAreicYm
xJZXjne72OWxAsf/7exlRAFQlfZDDB99ulTRmTXoj0mSsCq+BmhObAW8YPv2
ZSjYTeT5n/4wl/wdGdPmieruN+JDMNEt4YQ9WjeWzJyyeZUcqAn6VyzmqgIC
keIfu+tTcqmH4QfWGUaWjTUmB3lw0b6MxXw4kTGnBoffjqNxL0zYXpGvYmof
TDFybMy31V+41TM+1GKO5UteHT4DFNa9J0zDtbgx4P72xQOCSIgk0dEsY1XI
2yegIU0NIRBIoDJOQP+cH2HKiSpqBWBYeS9swlQCZEn5Yw0KjBnyY7Vsgn2Y
vURoLYfntJKwV+BWeWMOu0NDbc+TBqJ1oFc8E1dFbIOErO9dqieX9CsHfJHA
nNyXNyA2P6H6N832cXASM91T6ESn5Zm+5iWXndcpsrSsXIVi4sGFzi40BDnR
NqaDwfk16gjnxlZEEec7M/PfOaWctEqoZv8gm4xTsRvMsX5sK/e7I0c9v6xf
6BhHOLJ/pdIHy/JXPeXCaMMhwO8jVgrF7XbnEuzBUSjSHUR2ltwP10+H99bX
K2NflgmuaGDLSQS9f3FKDfOn1wYvP9YfK7OkU+vu9XtiuDJ6RlKoHT4WduFG
qfw4rsDVMploW6F5+iKf8kR3QdkszKRrkU0BZ1lKvQL2bQW/SJRFhkEyXQXf
Z1rcftDQPvdQiFPpOmdATxFgzrAonA79J32I7m8Zi2+CKMusXczMR9WET1wa
YSWtuCBr/KHyRIZlV87hpVnvPfkPxKkt7nqQmX0qdidJ7n3CqlmQ066XDI1U
TaqRNdZb/NciMMez8jwSc5XIvBCp3tQE+XRy1bHWUD79ca7AYLGge9PAVo1z
Uu0WyDvvzru/0QSs++OEiD5R/vpfGE7CnZfrvLr1tJKUb8nyw1mwLFhMeK/5
PUv6SDlke7Xi6Kj812oyY8rdDNxV3vbUZQ7tBDwM9STrUSYhaM1FPnYu7PyN
pppSMMk3ngkAQ62GBF9mdpXBs2KkREUOxjOV+0LUTFDA+RO1Dj1Xk+PKuXQ5
VpZe90IhxBkbvELwiiDCwverjXwuDOB2g188CE7hFA5lGDQ0dKF2uNbdQc7c
wAY2y8J7WtrY6kpXO01OmWBh+Natu3HkE9kkFP13U1Kq57fVIC9Mfju92Olp
uWjpZQhyN+TnbSzSiBiRvZpP5vgZImU2QvfXvMVNGZ0eZI2futjGpzMlXNNV
AzJ/Kr+WdgCKRULJdwwkAi0N8SGwU4uNEQ+z0RmPYYswPNaW16iOtLrsc6Cw
bT/RGCogOo0tCmaoE5RH2xilqUEkxcI0Pjiz7AC1o89skb/PyBFamoxKNuR0
5jdjAuN0f9Tx0hFMzabZWCjF3EGIOClGGrHhQbyvSkjGfWH5lQYFQ2tWonll
Sn1L6PjoehtGcMiRnBS0DgiyI75hb48HeIP0n+DusrLvtSSytT0NSZKYN4Bo
dmtc+hFlOuv7eChYqJRt6i3/bFtTplit3GMIEn7NuBlWrCNlZG6vmW/7Bozh
L1RwUmY7mwxD3TS6PwdNwmzhkAGtmEedfoq8vzwErN+wbdOiqepo77dB1NSe
nwr+p9kADfOPNGUvZyynEdgEtXNBviW7Y5giPJyTkSSgVGeaAB3QYfZdPihF
v2oud4K8igyuQd8ZvUCr3/gheiHdrmlGiN/WYgoVDgdfGhWgEev8i1GS0v3W
Yo1To/69fk+mLX4RM+tmZyJPapREOECZodiPFVyt4VtYm1+SwFybWzc9AJgt
LaITc9MPud8JmHyZLtzyDGtcaXl6PPdtObsJaVmH+AogZNMCAjCbpIGvPSke
C/y/DSl9G2GIwzb9s3/YUbCBIWXnEIQgQJCVlVQs2By3Xlke7dJIWAXh58Bc
rX8pUjjHvXkwjW2T9tZmmRHL5BZ+KgZyVHnNZBGR1oXcuaxIIZWTGe9owWSI
iYe4mWLm9EVWJcgke9iLvrXGMo4D7t7JYK5Y/2n4QPMfPSjV1wwmvO2xO3xO
Y/YlOvA3C5HTPwtVvvXLryPiS7ERk7gfSLQC57ChuzVaBVq8Lz0Wa/Uy5JkY
HNQORBNjBZ9N4UDCGb9UbeqCpWKaGmG87Lew23zBOaIsVtmU8/Xn0YkK6XRc
ZhnWddLV//LLS6qlo7C7MgWey0lV5B3Jm5eNdYi3wTu5OdtpMJMbRwyt73mc
hN8eELG/+CXoZVI7AukIfWUWv9lHVNSxz3y24W9eEIFU+i1aqXXwAFd+LiG5
bjxDVI7zzbS3HejAFi5zu1S3XBhhvPcxZ1jsOetBs+IPQwpKz8uUItot5fTr
/AhUrw7qWzfFb7ejtfpNB2804wnAm36reJXKxTabYIKxW2gqEfgoMFO5krY4
am6Ivb0odU7Z1O0QU8EVhnXDjVgNW+2OaQWYjJuIugNGI7uMrqVlpYZfZmdr
TSjbJ1i7tr8Pm72t/s6QmV6HhTe/dMOqwgnlAoRpNW3SiLLb48xC4WcDKD59
sBUWapF0p6hC34i7zkeG4gcwJGynZf6Xl0ALnGRWR8lTgFy4a9stxBE9OCOq
oVeXYTU1tGwCj5clRLe7u4mMev1tofdctH4BBdA4wWyHSN84REOA+Z39kg81
mjWjO9lLeia+RgqGriY3UHjku6vuDTp7T+bSN54e04lV5T2S4DT+Xki3+8iB
gl/AFqFKvZpVUhrqOfyi/lFPdS8v+fvZjVk/nvRZ/UcFZOSTIaEv30D5F8ZP
BkxcykXRxQv9SV+MTX1uKetM3UPoqvC935N36d4hOfj0AdMb2o+2Leygfyo1
J9AboutOyBOm9zwJ3AFcsnBUyCgJfP0mbDSnWVIw5v0O6Ya+X2kK2l3C8u3v
KeVLe5KFK+VzDnXhsnVw80DGivnxM1vx8i8vYJKc5cPncUnTtvgXA0jlMxYo
5SlUpayazwczbx5oXr72Cqxn8Up4awX9VKZJtSRJvzu4FXssuOJ+z7W+M8vG
ZTWpfLFPSzSu1/i1r7x2ZtFHAj9DZcHSatUJXq/fCoRY/F2Tq1cv8ankddJY
WuoDeZvKCPu887ylHFtDnqjLSpnlABcWSTRixGDtfycJzQPOsRGQ9G+kfJPo
r0QWl1iDM315vhYOS7dU7kt8Zh4IwOzkoQIFeoLMgH/WlTZ/NMyKJCtvvnst
bWNIo27J4gxBNbQ8ov5JX8XRBnmPj5W6QTrv0eMJxASvdQneJZxRNMxaK52y
7Q5zKpfgfaj4XlJOT74cW2R1UOAA6R2bI+Kvg7uSeREtVQvJ+QMQdTIFodMU
BpxWlUqb8AxgTi7dnXjDLZSztHdIWz91TapNIBWv0M7TyNF7Z8KtMSOagr6n
7bwR95FNwhmz/c9jiREoSBPN/e5Qk1ZwBOvT2B9JCVRaO0pNhJGvLIQAcq2H
7gk6Pn0HdTodi0WhCwijSqjDZBgJI7r11x2GZeMStG1SKjvA289f3tDOs7xh
wn2doTXbSRs5krSLFLkmaIx7iwRoop1GCpcNm0W10ksJ0tSygC+SXbIsgNi2
kq76vjfpEZ2RKFpKZ77FBCGfPF8fo6H0dSeBLcptE6wfvne92yoME+YdUB3v
V/1cprHkY7xNSWw/P3X3Wfm/n5nnBJjRA0z0ef8IvYZPO0Ru6wKBe87/hMsm
PEXgFt9dpxGuOZaTQM/QBa3UDhULBgAJCWTDo4ro1uA9Z35uj0IeBXVgQOPU
LonaTAIY8Es3gGhpk3F6lf+8k5ixHtGDyBWHkQN+zTsbn37i/WppGRSv1sAC
4lBZsR0drqUjtnY0UNUEEx3cp7UP0KDQ85Eu1vs8ceeZAoHjRB6ynhpolaIj
ipSAAkmBZiCQqWS3cAlilCZ7rCW5gJNfVmO9/2agNpqeS8AuAe88GV+PMdHJ
ZxQcEQmvlFX7OgcXnnnF8vrkJfVs7SQTuPGgWoiBsuNduD8N1estCawy2Ntn
i4/wEU1b6p5M11hKUEIhso401w8WZWexSU1A5R3Ngqyt38KlmVhlDV1Wmdxj
XSq4f81X7KloD1S5wU3PS5xeNwYTMks3oQ5y5JI+LnkROtefXemA6lvT6HkH
KSpQAR3wXEQm4/dLPmPLNuvJruqUhaqee3J7WsKwChlDRPhDkKnxKfPIjsPX
rb190/3MTpbGo8A0S8g6RKZGXIgNu3u0lhqZxQXBxdIUyqBa0rpG0NmlCjex
k0v9fToIyXM87wVGA1cvQ/vWGbP6UP5Yos4zGy136B7jIiosH76PCTT1YAyy
QNgX2Qqv7ik2vuVd+izpPXgxedZTsPWKTMFSX9OpMowzBAKfVDCJl2S3zNVI
PTe7/I9BOvXQ5bRWz0ZF7amoh6lBYcr55sR9vTiEp2K61lIPXcxX6tsYGSNw
ydMJLF1sp7pESNbKLpG16XaJSL9+IhWpqA/s05PmqFtM47W3zDSEvo1n3hYR
9IihkBPDXcOfVhZl8QCu9Sr8dK62ql4ZTvCwJhZTT7Ny8XmLO50xuoU2SowR
Tf9uSrJ1IEHd3p7W4GsHpB2FJ51O9QHURIU4PtT20EBL/ZJ876Gly3PfuBF6
AGQlqp82W2fuwpo3PpcPFHPQ1N9WhwbVTsCpADXF2EEkugc8a5GJJwKpPgY8
vxfWIJEAJrNNTnjF6BNgGElzsu8EOHZcNtuIJwZui78F7wG28fgpys//qCpz
ziJ6lpaRa/80Q+IUXXWm7voP4GwsXRugTbkS9iQ00RKKXfq6VBpvAtrTnKkw
mBhPwczRG6uVSAhlMX+HUWctk+G5jz1Wi43tDFKM9VFVrt+KRxgBRhTVcmrr
TSUj1ebrsxsw3nvmj4JconrYBxIToYvz25IKuL6Fu2iCnlgxjt7XXxb3y1Xt
gq5Z7tE2IZaKOxpSadLPsJLwB0sPwJZKTFwBKZW4Aa9p4Htkq7X8oZlSz7QZ
FI2XUrXTo5En0/N6nq4tdPAY5Y0gLaRbfWHE4awC/TNJKOHscSv7sjnJweX3
lrjGyVLitt4/F0fWAhIPY54d+bAWkhp0nX8Npyjy+Qt5SdiF16K4yrWZRTBS
Rlrv0Wuup6sheJKfY4333QDl2EduHR2pepLAGXx5g6fmJdNhSOCzKpX8harK
4P2n6gBz9p2XUgkD1wwKhtCqbl0nOd5+hbfbeIFF1zv542BsSEUT7DBYalTx
g1+tVAEOZrddGuxgJcLhgmQ3MQr47WoIWsp5zeNcJFJn0d66JLo3yFcZXXEB
3PkemnnaYJmMf62Jyo1ExKxjlK92+Ecgxh/UvwOFJM7W9AvYH4DzEjnQxx/U
kMj/JBbHA6hEZkBmWDRT1j8kGE6UFO+AKvlNIKPx9illNCBD89zfbj1POkv3
skMoQmeMaV9FxemyILmp3AMMyGo+NYccGrOeka7Ca1kJtujtACDeHj6QIbGd
V880EXbYTYS5xjdFUA/SR2ipyqavVLl30FxsMupt2hbsPKTpCsSXqguXbCKc
K6C56FralmrocC5Zxzy+FDadvJhZIOMzDUtHHeffGPTh09ZAG8LR9Q29eYrY
q5KC/USzulglyQfnOb7J5d1kvs9Oiu0+vKvSiif7eZ3cvEjEErFJKRKKmrcA
lEa8yLiqo0qfdP5fRhcFPnETtQzVvao+lk/WMq5EMXfqSNAScrFci5enMv3k
2/txiZWrrY2/4LaIBAD7jq9MjXyYD7JoWPg/AJ+vdRg0UaRbRgAHFeOj/YuB
gqtculf4g4afpL8RXyTsPxfOcUiywjvbMhlDx+EWNWDv43q8UpbH0Y+yzX3d
XMTiKqbT4bCEzkFT1sar/yXxtnZhIghVnV82wU56hciARi7AbpC7FgOJsZMA
fwXcmCEh1E0Wu6pH4j6ubw13U21gzLQlK7/u4KbXTecQY34ogR36p2KuuNXo
rKiWOT0XZOVRPoylZys1bvp5umdKEB+tx6p5gmUK9k4DdDbpG2vJV2fRf9Ou
oPZ1nhA9AkJkft/oJ8OxCWKQ1OzNVA3NQkV9xFEtoj6CXIXNDqIm8CTsUNYV
DGODT83NrPaHlAx+A1BWvoD/d5GtT7RxNNIGdZAbSkf1NiGRylEooQhZ7ini
T2xxHRGW5ID7/nAVcw7pKsTkImJfTYRiLfkxX5SaGAgBK7L3Vx+Bl4ZA4FGR
TcrDdqbcHhnhqncLigAn2U4WwsLIHtuAgxd2+mKS+AwzhEHN6U9ig5fuD3/2
ubLD1iW3gHKbO2Qx4i8YBLHo0qh4wWhgZ49xjKENKqjEONe/oq9ITBqFUOth
3fVpDr8y+oG3+N9yDSK4MvIMxDg2lTe26MeuG7dEyPZ/3zbpGYkbQM0JstMx
t4EIFPJZJDQdv17MfYG5OBaWMNaOY43qeQHHxzBz/b6wQsfbgPMCsOx4LNy2
dgh67JGNU2/y95veVVuGCOOH95wQktguFcAwZVq3qga1LaHOB25/zF05juk0
BK7OYdmb7v+IFsVqKvxuqol+Y20xdGWCd0xbVnRen9aZFe1VX2JxKmltwE21
j92BpHstOAFiYi9LZov/C/YygpdxhBNap+OFaEZNMraOZWt6W2OR7CQS/NZY
N3QnMBh2RcLqK7cAg5wSnH+PeQ7zDXvazuemfP8OGKWT1agWlwW5cdPy0Esh
DJapPFsD/V/DI7SCwTrIfenmY1c+r3KXviP/5H8GpwUSmUBdYfPE9+9Xysfi
fQ0gXuykp9Ci6yb0u+q6ZeIUXh3QxWajS84X9AiC/BDmqjzGyS68lZFs8G/b
NlSWgst0TjPME9iW5urAZGSzKmF3yNBr230VsT2XMtltjgFyaI8gnFcmVIo1
s0zakZExktZwmhCNDrcV5CM38ywAVc88pb9DMmFOyhpgnotHVlsdxhQ1H316
7iIJRmrkTQK4LkS7Jil6ZIF3Tl/R7Um7K2LRDw3ZX70KjiKjgj5DbeA7reVu
O67lVbIHMVPG1fjfhMNkgvylvZP2oQ/ovqSYi0RDFU7eyJS0YOqxf5fr+jDE
7XTXvFHxadoPGwZIVBKOjACbGetwfGvjJzRWTmM40OU4oV9mMRnGYP4+Ogni
fZNn2cttpYB23o7hEB/lMMVOMemVbatyjIVm4Kel1k1E6PiLkhW53Cxs4xA0
u3RB0EkdusBQRyNrIGOJBAV//7+VDFdjWKtDIKU1ABAHnvNOZkuVh8l1ZoR/
bW1dIy3DsGADiGD5OmCfTatYyAx/WyU1yLMEyZD3e+QB/HGGlVDgkuHP3GVz
bTvcFJhUhgqUZtrr+ioMxI3LssXfgHeRokFSuBHgDDW/7EMrK4DFuBEhaUpx
xMdT5mKfSasR7r+Uyr+/INJy61fRHOGKrkRbO3P/3kEvmIxDfr0kH2GQMcvW
kNmAQY5AQgh/S76WJJpqhdONcG8ks8KRqgQQYWiM4FxdDC3eneYfZlYtZZ8R
NnuvNwHm6CSoFCf/Nnu9Fwgx+LhkXEpKm9fGBe9YqGZyjUEk5QmsYm0aV2NI
O3xX0xwnGr8gCkELSm6Xn7nujIx97ic8DGscJbEf3pVOMfUWKIXqZNcIfG1W
7rG38aHpA9qiH+DWfrFiumN4MkWtuZhMuamdKWCqrqHvgutxYfoUYVtVsbOY
p/seDm7Fn3aHnrzT/WT2GE19Gw45dMtWYl5n5CVWsD+J9u71Xpwqw9RFJnwa
WJDmVUMwOg33NgISL3++2YL5QOzQ76rxWEvJwQfYs3vCuNIC2UhWhpZ30B6N
Ph9DPpmpCfb3bCHoVCxKLX4ZhBZPFmD/4SWNc0mCQuT9vpLUPOrj854px1Zr
SZKqhbsAKV4cm6751dzER1Wu14khOBq140XxrOj8Eov68/MxMWNKQoP3sBaS
ZDmqlovC0+XhAH2rv8NL/+nmhpcC/pJjCVG8Lp95OBpkdUsbiMIDO13Tmd3o
7/C2Qg4MG8MWlE6AUZubmGe4OcfscHbMmsQW99osD21Vy67A/MEnr5N9+n4u
pz6tOXfTrBBnYthogCEnKunNO5k/SFw9tljeoZJvEl1ADcG4TIOrl7MBkjWc
UpearMt6yzJRMlRE1iwsL9UrryJsNfFflv3rWhhrtsdejsFoAntZ5pKwVlF2
lGkHaWGvDoktnrvUzeHDQrU8yCjTEcRkpBH2z4JQwxYoYrOYq9j1kuoEf4TQ
adj+BecH23BmLrFU+GjGlX/tWGDY3fCD2j072oKe4lf6RN6QsT9dg7/UMRHp
+7AtPRz5WraNwdA9+0arCmhB+VOaCeKmEpB0oK5bdGRVNqswydMy+1KkQMzF
e0TZOpK4dwltdCYX54wzabuVJyNmVSyjhy0bwxkRlIJCLCxmsTt/xcUttj+7
WFhgAgLDFuNGa4t9xMIDOlEG6dB1Hc6W5rPGmWQE7NTz8OGQizWn2a+PZmj5
R7VFDRaT+3Ahmh6r7Q1ZuaTJnP/U4VrtizUnhHACb+qk1OjzyRg5uAd7xqoT
d/vVkcDjvRLVejm9Bzh2Aaa3AAm6noi+9IEWdrXaVKE6N37IS0KLKpi8S/ZT
thWKJRKCCyEeXeJuvrywCAJDbCN8UbSSmHblbhR8s5nYT2deaad6LTXHVlks
OeavAX4tioyOTGfNpWevZ2iAVjFQB4G3yXUSRvCDYtMpuXXi+KlDqfe9Iwy0
znzi+2MdYN1O+xhn/Jb9ff58f3Fh/1rQfnl0DckpKRm+Tf0+T+DVP8NlFRNw
aQVp3k/UDv2+y3ZL+fol7j27cS4/8COdvMIozE4Ykj0R39P/4uVA4wz3A9wr
XMFyBPFC5qmwvdWu/+hc+lcXwnNJJgGBV1MV6x1g2rCMAKdJHHvGD1FgrIi4
sqNcvtBnqxrFVnWTL9EWK1WqnFaXoOlXLFg9z63HeO66Ppn0hLGMxh4/B7Bm
0QE44l23866eB2SwkfKlDcNOw9wOMnRBaMfugthLsxwIkDMYsA5BRL7fmCoV
ZVW5fG65WzcrraFnxWntu4jSIrjTW77w/v7EsyZTMWvV6/bSuJomtdW9HRbR
QH7Y/ppcSghUW9B8+7a7vTY8nKxECV8+NVGnse08s++c8nauN2AfQDoU7mUQ
z0ENuq6rvmkuBZ4tENRnQtRTiphjlI4kl8kMBkEznF6WVEVAOCexAPjchLeC
LN9/5JRmHD+niZfm4EGGqJXgMSQHb9Ua06x0qJGJaiSpetxD5kyg1mg74upz
Vp5cuY7e4GAqPjaVlecHzDOy4JEVR9jkGbl0AK+1FNigxfsNe4/2A+URQ6im
aEWfZ/TDmi+4+aXVM89npcW3+VsbeXvR6N7e9B4M1YpcOKHg3bgYBUaNEDdw
OMrmMiCzNC6ik2kC3grh5bfe9pkPh+yVuoeQiLvDQzljbZ0pQxmILVAC/U9r
gvSynrF268AoTVjRkvU4sxOs0zj+8JzDBr5aG9qwUyojA01mpkARWW6XOUNX
DAzNE8BJhZxtoNEQ4kHOLFjOovGU1rPQuwGMargRfnEirR4S1I1+++hDLY1h
3D2gAJExko/7aOTWV950pffYzv2oRcNiJJXtZTTGYr7GqHlH5IUqBms6uAH1
Df0K92WcJIlfFqdXGIhz4Oyu+HwAMnA0MIamZoVbdhbBsdmodyRDmd53IL+M
mijv3NQTkhX44vF//CEPZaFzx4HdFeluLbF3gY6xXFOSKvg3wkR0H1xHu5pY
zT1WXKCruNSgjYaxTVgthMm0j5W42FFACSHTzAueaMrueG8jtxb1euTGLicK
K67nk/8kFqdRUOkjJai/9sp3IRa2Jylz1x4Rq1RONpnUUcjdymOTEOMnCIJA
xSpXTSAjXRoGuIOdFDPPxnSZNDBzgBjeLfU2/1gPoFtGx7k7V+Fv9uDE1W87
NtS/9Mwn9NvbJPGDpH70emw44WkRLLF8Rux9cRHfuvePtwYF8R0lT2WGoLTH
wA3vATHG2Agh85bzkw/nWCaghRVdJUMt37MXEvCdlLgKB7mr5aIjsItfg0LN
JGA97Yd992/v39MzCNiHmq13wBehvI2fJNcItYlfiXqOj6UBoxRuRaiDsV9r
wUSoUJY2Q6gm7FfsBkYK2PdhH1MD5Wq8+FCrBwbTp8P9uShULnN0zopwcWMk
sq0PBg/9bFGCbi1FT/OSj09ycWBfCOstom4IRLcMK4gnMcqmDgh2iIkewGzJ
QAkol/OZ2DXJORmfci3FYn/dcVIdT0gl+0m95/pbSZr4t+fhS94qQXxh0Y3Q
pURlCI4dZyQuamw8AohI8HsFjamElSIL1lfzwpKxM8FxXuIuJoPyd5311QoF
+C+PUqivBUi0A5W1NFanTQCrlv1rgQUIJukP0x1oP013zRRbt56riiux2nSt
RAr2bjFVWyAzGrg2mFKubrujeoZfUnq3FaXSALUK52S3oBNbG4s9xBaKS720
b7JAKP5d7haK6dXMHgpUTZ2MZHj6gyfyPlEG+DZC2WPC9hiMnqIc84KgUqBS
jMTbX/Xp3Yj+3QNXXuPM+lv/Tkz4Q5SNP4ctPKqUbIwmIZj7B3zVfjM6s9oN
4yis0bh4Dm/bzdyHzBslvhCXcX2wD6EsNxWBK29RVFhbdxFIDY/jdvnTUFF3
RVK6FYR5doBOJmsCTFygUmbAEK02lt9S1WFeX8PJUlh9Uxkmg/9c9Q8qe1wy
ADPfl8QcNccHVrLtMNlkQXSUf2yw9/1dLXQSOvyu/MYClIghyJzakDTYScdb
GE4A9tOGTiBWCcxbOrDhwKbu5tSYrr+1qwVgfxbYbsxfiWY/hKmg6RT7v2FC
PSy05NuTzZrTZkNWodudLzhaEBGurk9Zced4IyhSRarAlbrXi6Yuc4F1Bd4L
XXMyRnMezRNdbNEGviLzZm5ghcslbHUcQ2+x76FJsRDwVlYkDGSjGxxcZ2cb
DWHA73hP4hC2oOAJcWiqypmmFm9Oh7selACyuNVGQQW71cg2ouzDyt06hKn2
XemmUH4IBbJ3Zj9ZdSRjgaUH5oJFiNGkn6yxrNGZTJ9BlQevWwLE1CO2YjWS
K6TyFLzynEHLe9FeX+CLyCPGe5NzlFRsqt+65gAACz/zln5b+Q6Fec0gcHoK
W3Byb7V66fhjWkDpRzkGwoQEnQc2ufIuEw2Ip4YY1TcrtDAyWWaoVYBf5THV
FijDfs4S8b/jxeMb26pqvKE6xwNuDmoSmpaxyydqOuhOz9Xxvplb01nPveIy
O4J71KzMPUPror+/A1vpxJjiIxHxr6Poz8DgaO/d87kR2d63UtEfkdyJP+p9
ENSmddQbwEMmT9Uj7Y/ujcAg5yGdwJDwMNfkC7r1kmtSmDQb/BI8nrtAeGoa
dK0gFlOvzlIx//lQgWX4HXru+VWsChZOiiQ8lqQskdmuOKOE9slVX4FbVzGN
4mFKsvDvmu+RR2GEYcRZfr9ikKoSXuiNO1jKSD05HBeBw2x8I3XnmDRhLISu
L7Wo2GnzaLXPlKjCiZzwJKDXrIdzZT5ApSt1PaAbuCE+3gSaILx0HuF867i3
KM65+X74GD/bSUdjgvtNaj5NLwziu2ZQq5ypG7fdZ0aV2t9RC0W8WM5/Q50B
1G921PWIWoqJ7HK+Fty0S++NWOYeXohz6624B0j/4szQQ+W1coJjG9UpDkOI
/90ERwBR2Ci2LdwxObutW1nNDwBRaW1ZeNADWjN1FR9Xh4x0q02wyFjvMZKI
vstTH8j/vxz59EbPibij/tXFCexy6CrfX22uxrYBuD+wDKpYN2kzgYhf0pkc
wa+35Z+3bzZNy9gtr5K7zFV5aUZwcCtRB5+sO5jDAPn59L9ZdygyM2IhPtlg
P91/maL3TVCdujUjHlHTd7rrQzz2bKltVJ7fLvDrSY4zMeqQS8i+X4NnDCbs
nAIP3x8rKxkWLEv2ZcQpqgG9d1tEYXv35aJMbaPf73UuLVteRqTMEpF69Ssh
cOlr09OF+TvOPy9bc5HcFK1iF8T5/kGvQa/INsdsMLKPG6RhV5kqJ3ivVg5a
v+SZ4X1OPNhEhliPXRC5G3oQBc6RFjfJhbJMw4TfUFGYyGnmA63+pBzdeqDT
k1ekNhYTHddAsYkzVe2F40NUfN7YIVxv+LGHIiZeoxqxnT0OlMicRn4GHd5Z
ucdCDtyT+r64qbDblIJq8JOQ/p7y6ZQhU01gIorVUSfyly83dlmeiOws6OMo
UrFQoUpd8EgChODTfgh1mEFFqPuoFh5MAVqFkQdKNpgyBX6CsZ1mI9W+6itA
NXcgaltdzzbTexhBSuHKbs+SYGXDiUvbJ3/Ols982/tuNsNJP1/F4cxXsUHk
Im0ZpUKTvf4Db5Pf6jJ5NDTxvdvaDumGsiqi3Kzne5KbVT2aSxTsAJA63IVD
9RFwwHwuybfVmxxs1B8cJ59HhzOH3lrZCadbYvyvoE6GPS4/F8HhTphEGkKn
92Rsq3wdr0lS6S0TKe6Agine3mFVsgBr0LVDln9F7JPDHbF6+F9FXyKBJxoS
/RnbX5JzjOR4qsXsKInfk/sdHggjj1XNZw9NqJ+UT96E5D697QB7gOMBvVa8
YasK8n3mAcnY6G2+JwBBOTpXqNIkRDSKeWXyLqgV2YYbpbdffW/tXIVlxxW9
+eYTtxg5UtWE2SyLjaXHbKJqb+uyohpMWPQmhWJP9W7+a2IzoIupdhRPJegT
YD5UdNB/g+AuosN0EGw5c3zQm8Z7Eg/RnfzoZIKVNLYmJ3o9gRg6EVuMj6Dp
t/ydVSs3yFEjc/Iw/XIhlq56CyUZdVXOIlkm43N04rlQ/2tBwDpHFlO1JaKr
UYBmxu/32LIuysv32gGJlN+/lTCuPrygHKJNSKqAdcUvCct0awJZNvcgnHjz
l/Dcs+b4fQA9XnNhLycaTm3JtYlNDUn8boMPeOkSOVZWju7zLgLzrKOD5ZpL
n946LzvgaW5+L6D4f3idVnMSlHSsu5yP/nuLdjmzMNVojSupTDeqEHiEGgv4
XFqKGmkEVbWXUlOK3Cqp1uiY3oAuXMckNwtKk9VQsiZsdIfgOqK4gqVbnbd+
bV/UixE435Z10Cbe0YdZcJrhypVKDJFjUtmDe8xh2nIPo/ebfoXkwPQm2zTb
XPbie0Cq7I0t9LiI1meuWNehR4fz9yyBI7/L3J2/7/nITH/gKLQBUUXbQ3x4
PIlMHewPojeUmbnQlNKXikSTpYmNAsUn3ajT2NeCGzNFY93aeGsda7oBU2E9
EvDpFEoiw8a8eD0rhZFyzQP6OZXIPajJl/7ATP1YeBhPlLuPlSYGPZF7QyKY
aFCIxV3ipbo+YChb4PGYj08PWkjunkMahiiHSkSmzyfj1Jn1cXCOls/lmcoA
NzzMZXZ9LY2WdLQ3Og4RSPPSaNEWiMW2Vl1+TiNpFm0qy7ohOaANzGqOT8kN
A/ROhaH4BRAiTF27pQjhbZVMoagm7a/0EDI1MHIEFnuZ4TYtzBaBk14kID7/
5ENz5MyH2LB0bZpsc1jZ+PgZ0f4pna4jrgnX89xrjsEGGUUV8N8pY/Lr2IEp
4YVIcCbK9y9g/HEOrrI7GdqQC3WgTeo7H9mhow5eh0rmGSBczc693uTTq4br
/K9rJDAErVNsPhuHmSX63R5Ih6Lbhuqz0Hk8sq0D5pQw5U7t4WtRVCCuePUh
OSJOH1V96JLApXth3on3RTZuHjcKJfbCGR1I53327TgxautpBKezZZ1fF6uu
PqSX1IgjjcKluO8WLE3TT1hGwVfLq9sohtLUFBtxX8r7CTs+PpFpt/arLTBq
W68Y9o0WfcxF7itR7SuRUuhbFfexFHkVxC/KR9BAK4NiLo2459KsIyaFWCTD
jQCUcL/1eRMDEtl1dx7CY4nxtJv9+7IA8drh1YafnNTerwcNOUKAz0N3w0YO
J2/u65d7miRZus28fYAHMCmxKWr6Wpl96S0LwB7nnVlRgC84OUIDTkMktRbX
Ii8aXlNGDYRRiPchQHfFH6WYt/O3V7Rzuv52X1CqyY9bHipxGH+5QbbLThku
2g2zGThYP1lmv4gzenyODf8CEvgq6SLPjQLmq5jWRWmjVuqDGkAUrHlLaEkH
EjEOF4/TRr1A8hBF5DMzaKhmfoLgBHFpwGNeiU5Sphfy2EdFNRCQcCR+Vx3O
T66iZy1kesfpcQzGi8wXlQVIZhFeEzw/hCBUC6C2M0EI1SSI/3KJLRU74zzr
sPbRLBGfmRh0b7ibigMfoNKfngpmkcG1A8nQad5vR9UbSggsETkzOnUtVtla
9WUXIRP8SaX49WnEy6pI0E56owk7gyQEiiwhvJtVw940pdYnYY7zQCTOgRfu
9ayDBbk+oihdDPJYc/apcfLb2AS4+5Yoznq8PjJmsnm0U5qDuecGCSpjRuSq
Jgb9xCW/RJzYvqc3RtrQ6aCvs9ObDXLrTRvrWGMhucPpYR2LUqyfEDJ4/OXD
rN2s4cIHUEaTA4GvrJVs3tUG4Z/qNU6y2NE1qXKU4SpVSkhTxFEbAdfapvhb
S8Qi9vuUcxMSScWgYJk0aRUnN367Mpdc0RIz6cg68nWoB4oYlhbhIwf59cab
LQB9/MjPc6mdx6gHvLNHS+jwAe2uKN1jiBzrA25SRBt+TerI/OouYiK5XMuI
9QOCjt64/eLwZcvPmMk/cUh2ab3UOIrHBKGpi31YvtaN/DRkFXuJupFCI5k1
J/uTQbhy0eDw7/WG0mfKXSe08dYNHeBB7EbtJxg3Nu8PMYTPh31u0akzQObt
dnKPQmaVLgZHYtqdAEVldyzZG4l2k7hTkd3CrAhbvh4glAge6erHH7XGEmX6
sOOJZJcrzQaAZiEgITDwN8APbVm5t/pi8iPBamp9js1+9rLHQZ5GCmtqYN1S
3g2l6mM/RJKtpVPMoM7O65WRwkyxc+KAkhe4hKYoZ3SZQIebjE9gNOCOYLmU
+j1llmRWEAQQt2s1KGKFYmiILKhvgZi3A3aLWQFFbHRjpm7sWPgdLo6Jl2Sd
FZTxipqMavD5HDnUhbCjDiy62dQE/92vhR+KEkMitT0eXvTyxr4DMVR30qPa
j5eE5J74bp1eI65Fp65Gyn7nUI7ZBWYzz23p1RVLtfjzh35e/w7jumHsxn2T
IjTry3Kj+00dTe6e47CMu0CRA745NKAYdOwzlW+oVqkmWv1Xo2rhwuSTjpgp
FPKVWhyHFzbGyZzJ9nAuD9SHhEBOVSaZYq43w8SWx/u8d+eyNFZHC0gR6w4E
h6r84ifT6FqQL5Js5plK56ZU4NUR7MzMJO/7Zy00L12FJ4AfqcckO2VqHz1E
L7J2fUHtxPYWuE7bs+SlHXPacNQDdVBJHNB//7KvCOoQTTYLXh1OUMp2c++y
EZlDpMR9dpTh/m3An2kdqLXDAjJjvHxFHo1J5riW9dRqKXUTvc0TwlHxhoRs
8mzBJCMQKjNJP67dF5eV16+NTIkcq1OI+acr2akj3AUJC78KHVuZLrVJ6kkg
dUutjdTCLgfQDvLAXn5SvJKMRjzOIlZfD8mZzdP6zDXm8x+3Lv4gIxq5BXy6
32gJtElVyQ9UDeWmeX0wtVpBl9/hVxlqwbxTf3e+AramNnPu15UiHe/aM8t4
Zx0N2A/NsOTaeqbxVdmRGR9mltaW7FM+07c1I1GlFcX3GE9gx84+uZ0Y2yix
UIyJfx1k96IpRCID3zOhCMcioOYEI7y3UTOqSl8fBA6CyfcBb7vOkwGmqMSa
+76jKG2QesOawSayzWvu1W7nhgpIqqpdG5LDFykZBDBplq4VVqvcxfEZqoo5
Cei8zhKE3fme5Kc0rCNZYVKROOJ0PCfqyp0KNytiVQTI1PS2jgr/CDudc8Lv
lRs0jvdK/kGLNlxQWESwaZNu5Je4ZZXGxIA/8jEn+zvopSiIXIPGdPY1+y48
rkAnXV63zTw8WyRh7nPS5eOA3uj+MlOdw+l5+7TVlZh0+pTVLxpCzUDCg1In
4LxHbPf/gqZZ/dTzQibWR8QEl7sDwa615pNuQ2BCQW4WSd6a0yW/12s2+S5Y
jAEwRl7O2uxA/wOHq0l7qVxAtXzhzjlb9ydt25DEMxD+g/P3xLcQpxRIHaDp
2xdlwTFDGW2CLSYIuVPN/Kqf79iPz8vO3hp4hCOYDXVWBAbw1DgM3UyINo0c
SmS1k/fQtH1U6HCEwxPWM25Nm4Nl72dYtNgypCGIuwaxoQoyT0GXynQhqVFM
2e8AnI5hSoc5MCJH12vwkWsjv4JRlvkFm53hMRDo9nwc+pSBckCMAthPUnGG
zm2gS0XYgb+sYPQbOo+ApIWNXvwhHwIT8T37qIxu+Dkr+Z3Hdg0936DE45NJ
OAz110obJfxcnASv7IlQbuROk4oVGPzq1MC15jmj1u4adF4YlYRnacz5gtMw
RjleCaxXxAA0UCLVG/8jposxBYIac+pGf9lCykzbFZSw6h85BML0aZ7DWOW2
pXTXlvaBhRKjvNkrI2lBCwekWoN6vd6R7qeB+buHnrdD/+t3IKyfxHPFFA7i
ys4m0dpXqM1udfytgL3ulr0PtNwIEw/llFXdw787ET2JT4nz1GHbID7pILr7
7WcerkVxEV9nIEAovThg2z0B467Mx0eH+QxkEbp8rgY7QodBl6tlb7+/ITxT
VDrkabXC7UU4kpocJ9JUxdhkv8k/ZkH4FRXaKffm9ou93ufCKzkF0j8EF1f2
yYl97kIYJlhFIt1lgHL4UGZKOQTUdzu3yw/F8aw/B0qDal+bqde99NPHyb3I
uRP+L89C2ui5BbpMVdZyHFThcBjt610OSiWTvhyY3R0DZ2p0OYp+QIoBM34S
Zrzcj0AuvoGKavi9kBw8NpFU/el6bLHWNqvy/ih3tkqwvwABXvYqEUxp3ZBC
mutHRBp0YmpiO/OOUN/qBFkJy1GpKtcOCnSawfr4VJ8/t6GmqJS0qmP5sMSr
aLAK5RJoA5Nr/IbWJ4i/Il0YSsCZa5mI58p8CZVtce5R4KJHd5B9geB4ffKQ
+5zDhunXLlFfXiGff8a/spASL1nHho0WHwAO7Zxo+omxXX6azA8BvtXNm5FF
b3E7wbBLGzCUW8m+DmsS25518jRIWuwSxJbNH8Kn1Ceo3baC10xWB/bT5p/Y
srMFiFEZ5ROXiLV3cPQi3QL7QPx4QIaWkRtVvT7Pu27C0GZAUDjtifHqwRBT
0iF1O6iCf5CLgkyp+S2KZIJuY2etAcjpA9V91kpYfoqkidGyIp4GrrFDwITI
jeZZ9EvljhaRpWHaq40A//ynnbGjCZR3ANRW9qFFfAqa/JpCjmNlDVvjLZlP
W56K7nzPb9ljMCXubpDagGue64yvF78hX0vDL/bwlUQ5KwUv/vsq1kGQpkaR
FZ+0vUQiClqx9XdurJfi71EB5wxwKCUKx6vizZ1VlqS881bygfunyTlWb7jw
aRtKlxg0BmXqzoRkuWX4cHwOcnjFaOeMgo6i2jXlVFEbi5Dx9WkYFJz36L5E
xOFTCy064WaRvHcyV7kXd+50P2aEKpQnRSL1P3vWg1Re8rmo+MLEAcW0N/k2
RmyxTCPasJe89rIkC3mW2bKfk24rlLqFO5miJsv3jISE/NZ2jrC4SOD2M5Zv
i+bMRnkWwqXYDh3qPa8kZ/k7GDhFL2NCYKQBJBKVUM74BdaCQy4ia6WCW/SQ
bXS2DjfEnzaSdBob/lbjybYFntnpak9Y0aoieBJfX7KZnb0nyuR3KVXB2E6V
3x7hHav7xIXc3HcVHr+2FvFNodjpUs8W0ktxt6WKPHoSOUUh8ZGZNMjFDAsB
hXSiANdUQNZzKY6Mx7HbAHZcbaHnnWROqSsaFRMuV1C9LsNMEBPe+kqQYQOG
+ohkqmmHRULulKWQPK+oB4Am23jXkAx52Ei5WJW6MvAE46ns/0OR6WjaMB1a
pty7O0styaSB87bP+LHfPG855bI8QKXPRNMZDtQ1ORoqWeyaqL80POoZXBdj
qohyFuwsI0uJFxbdAGfwGarLuaTiTHHGMEIGIOzjRVawMkdSng7Q5Ca0E0/J
RXFrWHKvgLpNUfRWfk0sfRFMviNiTs0LILdxtxEY05o5s0eYWEDc71L5yXle
xwocitirmVEtYskrOt2xb14MZRYf3bnd/wNCXvHgoMHOl8BlFB9o+uu5515C
86n/MwoiaRswiDsa87ll36y6exIR7vPm/HVBLZKqg5F96Pjpbfg8hxrRiAK3
o9vxyGcBt7yWdyBuiO6RFzdo+PINnLaBcOm2iH0myV1zpClCaN29v0IAPLXP
FUoTkzeb6dHbkxkqTVayE8AT18n66yfRUd63uI0Qv8kz+Q9pXtDZFnmXbif7
4e441mHuxgRl5pES8qIrfvZA5OZEaD+wkPJzuDBAre1T9zqveRZudSIAH1AE
XM0UD+TxH1nUKJaZc//73MUbLoIVzhbvBLq+EFIPCxMFMU3sCv9cjWLMdYzd
pRENPxD/kB1Sm0xMMcwfJxfVjLdrE/nx/NIQp9m+tSMotXRWldtqvO1gxAqN
OggSIXRUemcNtOW/HW7p/eK/PwEwUgGw9EV9lqh8TEXRg4JtHu4/r6BzoToP
GVfcNHtJQDlmwg2Lr25fLlExZtpbK9ERRgnPvvR5Kot5GsgKgek60ptxDHJK
R3BQBjwuOwp/uL6/j1TzPFQRHfJKFu01X5x1wTd1qL201pP/Eq6lxO3qHvwg
k1rZxpKP4jYJ8TUgpXwS956wzBygr+3Rmwt8Tzpey12WSfxAdRCvDEElvr7F
5EH7QfQUIjNWkIy1ziyufIIuPWk3Nx64QGvhSMZFXJH+X1FlABuI6HVSQ9Ee
ltnvmQt0GVcixfxc4BUni86Z2hMo1ZtIy0XJCTFoC91NYFq65KYOvOG9IgOI
Ab7S9SUngwmgJUlMLvehRvKnSof0FlI7Q6Nn+AHnx5JMnlsWtjZPMqvgYCmo
Beg2VqO+AUqluuI9C2wy5HMV0VHAMZ8zc8ClRJpJJ8dF2h75c8aJ+nK62OsM
w2bMhrMIHniBKgHCCNQblSKtA54sQ2RKqLYerTvv0nXU3Xhrn+mddFRfK8W1
NkAoOw393V+FaixwDFYCKXSEgybYtuDq5mNUXMoZmhGd9Cd7KjvCbEGEi9Tl
L88cwhKji6OdUiHwprm0hHW2NJmuDsRpI7KTW+US8rzaLu2EIETvNPJno3Up
J4bauB/kR+6Vg/MmzGC+coJHGDHIZUwyDg8QZPl2TxIDh7M84JET5Z/QtOpP
x/4wpBayHvSrk/6gDeEUwuWb2uaof4FZ0wpQxQLhHCgrq6oPRJv8qUWehhA5
42NO+R19ULaNvNF/fxLQuVNHl4o5lskpy/S16vs+24Gdue/hK+HrM6jNnCWD
x19/jk/cEmJIg7L7Qc2qq+0d7U9z3DetQuxdy/gfG84CiACZiFaA7+6OxBRN
5fS6tHTdSjp7Wv0jB5qs50AJ76GCPcg+wQwE7mOUr/41/CwhY9PYRyJPLAl5
tLxD6hjL5dyXnWbHUaTmT7YX5rRp/GKLymnzo60H1L8LyL5YXc595BFLVm+a
RCDq3J4gCItNZRZVL6jkHEqiU7odBhyaWi4MPA9CexnZkznBTAeDgskxX28j
tGfbCc5CtmX+b3Ul0YgaVxjj3mR+6va7CvHTUldRU0KJzcZ4Co08s5NCQaKD
DlSFuEURs4PYPxPlMZAjeYAt9jRt9qdxbrltmBZOmoPTLZae08eqTYuBLxCg
r1nNAvM2tLWMROpBVgqZIgheB7hprMBtvO+sp7KSEMa4BknkkMGUSFrRR9YL
Sj5RgqtfY4vzt4JzIG6CBvYh/CX1Y9cJUeYypzn4YUYJUkcbHS5O+4+K8WHs
vbUm5jRVWZH/Gpa9bB93zsm9MIRfo8ouVzWRe4+rQPfgnXY9SEq+THy8temt
3PYVBgMG106rhA/H4Bj+jHdQ0nB9/UZE51yQnP7jQ8DDeclEKDTDHwsaDtkd
RzYELGMH82Nl3aGji9sqHBxqa1qCa80AR4jk5dfF5F4gfHrXkrvYZDUS4y+S
pm0ubgaOIVuSMQTNFdaFJM1ZS911DAA5s35eww7mGunwr2IyAWwkedUKduc3
hp77jZ17PbRObJu7Bc9ghyxICr6u7H0FWcHBFeBqYgZJ0vBnjSalvfBZT42U
/mZvIe4UBJgXYCqstKhNUVHiUwgSqb9l7F0GzbVUqXwTLtTmz7eixCspzLa2
AaOlIIZofKDdTeMvw7lVEpMf5TW50dqJ2fDiHhAOBw1VpNkfW4pYrUYXE9S7
p4AEJo9m9F8F45qOeUVAGgxiCg8wCHMwdbKT6lAQiH0nwirQ4wP+ya+/85UV
UszchX+nFtE9ON5CdylCV45ZOnFsQ6e7vPLk9z00A5rnTK4PFXWyMSu4CzvX
UALOCjXi+8TQWCg1mXiV9mz2EjFM3Typr5HoswtgeuHe8u/sw5gCEb/UezrE
mZ7yMJtyXpFtrcU969pyTdGSk39ayA9Nmbuo2WTTCsAMFlH/nQE3i6rFrKHn
ttsazsosxZZrcUerizLGeBwkNUCE11G02vS6/UISEk4Kyb65YfwPOcN/qu/X
vPW7B4Q8vKFXxQRvod0n+DxWheFW78bLSED2PlQNSJVOz1h4k2XHwolpECv7
nB+NFa+/YCEXZT1aKnu/so5uXhHZ8cePSeGyIYTo8aPpiDafEAPNfARe8+aP
mhDnTVNztBmw4x2GPSZfHe/ac0crKjQ/bGLFif/4Sbd3i88bgN9yQz075ifn
dYoAlQOr+R0CMz2XKATEOG9RU9WfmsRYejo47l18BmczJ7Dbq0HLG1X12L77
MvNa07fRKlMihl/irsucgcky+2QLhzx0Scl11ZpoS6qkK2ZpSgc04uiGvJa1
wGPZZUOPj3HLENZ7MFkSc7DCVQqe7P5POJIX53FjB32teSjTp37fGbtTMKFm
KqjfXGMqqb34opkqThA+ugZmFBnEEBiJVE4+2dBIc+URmz5XzvfW65jOadp+
YQ4Prnk9vXV/0ijgUBgyDVtjXj8oKFWYcMtvgvZ8ORGR/6k+sSW1oS6Tcf1T
t7XnMTDNRxKO1l3m8XzLsJFuWvXiCOzbJPpDZn48EX1ludqU7TKYKyBJTFb3
7U8pdyDn8hEXjEfGwCk/3eo4w+uK1Kf/wm8CoZuIvIDdQyFce5VzC6WyZ5d4
99Pp9u9OiZuIzueiQxxLIDmJXp9Q7TjHPDCB+c3Ya96Dg9tfGEtmshkoq2SS
/w0h09uBnY8xLI1eyFzU3HRf+5RmyAyMfhEwYTaQv4tV3+rIEisfgO9Gmjo8
AQOGNxfJ3R4Y5MHZuHStX+AxsWsWNzzsOfaiB7lKkqESpCjlPo2xcJbKTotj
VSiWtVefcUjaZw67DpsN/045slR0IV31xtTuug/Bzkb2f7PKytDaJYa8OTbG
uWnO8n3wtyeamFoqLbKdAcWMl60MCatnTeE5lt7PKZG/2D1tZh7xYF1+ovNr
3wFSYhcvGx0ZNIEyy2eIZm8V1bvxKXLPEFgAfXJwe6XcU7qBl/Jm/KQc7uJg
PSejsFmG/6G7r7yLmQPGckVfavulYENS9Ya0agx5tKvHBBU1rEg91rdAfDy1
Y7i11xk/+33FFGkLwAf56ii4N9r/lZdmg53vJTf8nJIfXXj1Waz70IgyCnEk
exo9CG080f9x1fm1w6LShnsWPFBzwsKBx+Pcyh1aPDnoE0UCf//Und8hNbDC
20mnmXEZOa21GpylESdI0jbgLKMwmDyr3xs+i/Or3OsZ54X9LXiW43oDnMTs
nQzGz3vKnnR8GxnmoMbKbIdIC6sQwsP1L/SohwwlR7ASD3Xc4QLssCN14tvH
F3GC0u+ncXtaPoqawWmuhtQTTcGFYBH3YbWRkBJS4LLI7RGRT9kp+EW0ebqL
cwgMmyvKwWSvyapgVF6b5D0G9N6YuL9gmZVO54kIGtR+jJ8UXf7pFVIq0dmE
M3bk8hAobEn0N9N481c/sU3xT6wivqOoiUbxFvOz/LMVF27TNKRUTmgr935t
UwYzKtk5SNYGoSxNRysUEwBcnQ+URZ/azYYA5bRtGOYgIOlBMfvsUDpUXeEs
fVy31BjQqP/q2oOe6N8sO7dqm5XYS0p8Irx+AVoYV07/9CkBG0XrONGq8dbE
p1EPDejheZU/VcXWBSXSAABBf6qNhdom+8AT0mw+mTElz3bartAebR4Rdjts
MbAENqXtRpnOjCPSPmQcOTOw+IygYFvOSYjxpHsBAMIXcDC5gDZIiRcz15tZ
WopA+YT8FKrZueeF3M//JHlmZEvAGemNj7M8+EbmJFAP4MzjwxAsgBWI0vsW
1iumbqd9c1SzseVWxzJLZ+qHH1KiyQYw9lssC6Pupe4dimIsPtxP5NixfRfi
stEpPzRg2eOo9tUrmM5qHk5to5S9ZjQjE4yg6abEfcL6FNooawK9NHDFQGmL
kFWz2c1Z7natko8ZlDna8agHXbVfX2Sb07WRPHCPzE1UASqZSxhx6Wl555En
i0Mb8iVOmEPss3yReFy0LJX+1AF29PHbKTQqcH/bksf2yX/Jdc6xpOszqkg9
GcWsJ9eYCFsmGLSb/rVZ5ckuRL8/GLNoAhHz3FtjVmF6ywZqwnB0apvqYd8L
zR8zbAIm5jC7qCN6b0hUXOxLUp4Fc73IJ987SP/0J5+tq+hzFid0RivjJxGm
S5ryS/f8F3PvqFbA0QwpdItD9J7DkpHoMgcHHEz/CYRZKy10SWhc/fNzowbd
16UatPNWHbc7xpf5C+IEEzL1Fea7XjdjB4dE4SFU6S2g5BAH1nFv9Zjs1LpW
nALqvZ9Q4CUSXoW3DtBiJoK+emNx8iD+erpTOHikKSxnhAdEKsVtIhyFIsSK
YNECNNxdcFKxz2r/xSEn9oRTjbKZf21bZtzjZIrucfS/rcxNfUoOTMeox/3r
QNXTXlPqZ3O9VtZPK9C1A/QQq37M9Uz1Z7JeyXF0rckFC6ReVcZkhYC9dHYB
cLfp0JC7zHDoBKDlTzQuTNaKS8MB+3j4H0F9LINLi5PTnqhlOm4sP0se4ORe
mNBXp5FqzGBR/8KXNz7DetNsOBhXontUJULVgq/BX9vAgThk4D26RrYza0wB
R/0tU4lvelbxOcPPw/9Ft/8yJF6t/WVxaI7FOSPTJpgyTXpu/LF/86cR5DNs
hShPHR9edjBTlAcizjCKRQOBAaLtYvZ+v175tXmfC0DvI2W0uKo9t+fYu8od
bEL/UW7gDBWCpNCGEEWeigA3+n//LHB87RjIGqAGTHJtyid5vme+Sdze8CTf
fdaWzkblRFA+htDsdwvms9egA3lV8RqnREXGGE4WIYyS8FBCCHBQ4fykd1Ia
WHWPA9QnT3BnVuTo6mMMsgumRAxaw4TVDrestFZ5H73Pk8Upc7BK9D4SjRhP
TQDFFkgqa/Igofc0KePKcvtuXMJW1oo7Csw6UzHWmnTgh09GsuWHjnl3Gi8L
OZHmt1G8Ea+iTjOoexKpsnsubTTqL/AS9YClG6Ck8hhs1c0C0xJbB76Yywh4
vG/9RTsfVDwxQNhNxi56piieD+axNr4xmIbgUocg6rt6SWKGAOklclwT/Pw7
2BIbuU514h1P4reEG572c57ZnI5vOkXoOWR03RoWk4UEsQeNh199huCI/o9P
EVrUdM1CiTez4DBL8xLIFKFof2gecSNPS2hH8oVqqGEE/zqxnLeiqcaws543
e1SQoejUXXXg++ingcJVZRWhAVtqxz/JzHtW5VmL/aKXSUii3OBOMUmI4mGI
joeFr9CoKwEzZCWrs9QL0XAD8s+vi+1FCkvFBPLX1YwIdmH2PgKkdtTLSoJy
CLxLlYCLxFlkv2tgiWrQYe+FPJ2g8JrMmNwM0AOg3FCMTR1JVRy3IpgfzmIq
O1Uf4jjyKRW0X9w2KlH8foSnO77PvQ2zBODmlWVCDlLbCC1bfou+VwQR96Hy
tLcVDgTWOwdH1iDTAUaYooRh5KNR/7Ex8J3afD9QGaoAYRTTg0IPPn6PFM4D
47PRNZpC9A+GtOaPSkssbQnGYdS/F8N/qYTGwRIKPOzMLRvRL2W2HkIQXFLj
dQ9l5g1Nku7Px6uRWfYXq2PrIG7mPeFWkRqrUJzNRmwilg1nofKqXCyrhLq2
awBzm5vYm9x4TmIgHKKZ2fx0BAKKqWMqEKbhMrqFY9e5b73iRqOlaS3Wn7UY
YdA7OgYceIlujg/lgLHevHLigVIf2YZRKYGFhnjszemjCQUwQMy6gZIuWPc/
ZfguZk7QoG1pJ1rJo+vhXxBf5P7P/zTXiIX/qJQX6U48VaD1q4IyDm27RG+x
orbtwzCX3/LkIu3treREznojwg3U88/YT/wV0j00NY53V/xNkvnp9zrwqFlS
Lpul6h8beDrebJQRRTPnJwPu56aF9fv2yD/Xc8nljORbVnyo+bnzUFQvonNt
wQFdFebInS6K+ILfWzqG/MrH521AFsqt1dkIQ7UGd8uKdiSA+MhRgfp7+DOa
7l4Irz/MMF5M+I5hHRd3vkxzmTeIHwQB27NV2fiX7HYAeEQ8i9ujy51WAECb
KJ5KisvXDZASZP4CA5ZpZUjq+xb4LAQO5icWc3hLIQnoNgzee+hgictbuIX2
SArAvh1B9OEIHGmYktxqJDvN68UoF2ZBNyHq/VAVJXzk4NxYDzLPu90/3+BI
pwgUbtUY3YbwNo1Bv9/NbDrG1NIIjxmy6DTmzZnxCsr80IaIt+phLjCtuMyg
VSKhdJVABzaADd+mCmeGuoXMnus2MRFsHxpt3yYMiTA1ww3AgHGPnfbdUT3P
2X2wRcBvaHDw0lQhnWocr9x7WL25tTEeR5vTyHU1PtUjFIwPgxwG37pjbSeK
lSt/vGpsMI+y0t5ARIVFwELiqLoRi7nHPnJDn9pvFvHs3fpoxRnO7NClT2gQ
2pomHfOl/I/kBXj1gPBJyLfJBRhzuNYGJOB+/6dWsnuvaX2e20dz4Xhov0NV
5MNPAiMsj+6yHnN9vjLLs8NgrwOep+WzUlp7af9nYmc/kNidJ0mjQIQ1xD28
bcvr6lXIXcbjQMor+63gMbRoJntQx9xbkcP9ORs0NXnKJb32IuXBYzZt7y1i
aT+WgcyiGmnF1pGX9xkF/AjlRErTFyOjCrNzFXMmRjk1TSXTN9/DPxrLDM3W
kA+qFoSaZfIuKJtlYDGoKHcqoKPFG90zLXxdhuu7sq+/T83xtNdLSXXWhjZ5
kob1eMCzeiVVxVgXtSga45br97JUPfMxhTXcAE9OdIyOb9sIaB9vuL3sLy4E
ZU2LMupEslCPnP7NQ0yV7N2nEA4VRVAJmSm3OTLp32Jq0B4df4HA/z7hB2RV
XS+LwmC0Xh+lsXXJbGFNAjN/f6GqJlrMAtu5zJuNcJRomFLWF0C0/HlIvBFD
QT2ruVWQDNuEaA0gOuZ7D6k/OOKk6PEUr5vP/XdcOSdZmY+l46y3tZMa6WEv
nxP9UD51dCKIptD9FztzD31JOMjswF9hY0+wl4oZBingszKlAL9YTOpUaeoJ
sqGN6ZKST/icAKidurC3+F6V9h1M+xJlBvwAnMgtZ8YxHhK9E2Sb6MAaTktb
UaMAQAAZIbNQOEJmBNXGU1Mfv3455WsbljS9XrvCvuGW07KAM9/fG5vgKVrt
AAAlZGecyWSbdu+Hq5A7eHnPubkl1nxboA/YC5ScUcA4MGVGsLCl2zcoc84M
zWMCN2Hcm9vVY7tXyoRHHKHbPvEembFHOOoQ3U2T4NvfDGW+TMw3GnOSjN80
vY9x2DWeglIzdoWSGUgmZULSqnIsqoRmRQ8NiiDF7nT/1f3R0lryCqL+e/sI
XAD32wV1KkE3td9HOr+/YvW4NplIbwY5tM1/c661M17sqgdSEPg1cF8mYpGs
1XJpwACNUsMBYvvCV/bXpbwLLSYGtr6DnNJaIIwiYsinCTvwVA7ZbOk0lmVd
9wmBOVpeOgBNBjZXJsgUC+RDVgtcjbPg8862Q8yf0s7uoHjvpiKPMhBazlnA
bfoMNW1+9BW8B3TL3R/dnsBDPO+MwLo+9mcyRszv6slFM4SHWDe9MIbIAB5Y
u5J2RlSNQ+EiQBhG1KCzzxDIH0Ps8zrdCg6svWm+D0OYGHJBJwVjhnWzgykA
5VO3gbQIOHT6iO5PIZDJSyx4YWjuXwosENN0xiQmDmT6ICyUUwB0x90pRrYj
NHpLZPMZzme+YNh/ngGDku1iVSvGcL66YZUsXVjxWD+Rh6lsCHYJpsmj4j6G
A5n9iGsYIvKgOn7J5SEbPj1YSDLsA5PuVONEyON/kKNlPJE7ftbEt3SbnZdx
91unX3m4ASsnGlQv7J3uMecKOsJegdB+U+4eHkftKdrLPceXQbxuZQwV9q6q
TksmgawqW8YydPXn6UItwPU9VTdphRN916oNQVVBZ0LJI3ZINDway6PBK8E/
sI4HEe1psNUSUw6C7n8Ac2PgSHEVT6RrPrb8OpigBJiCKgLPZGk5LRLNLka9
k/APHJeDJRDjwtJ6d+gYSZSYFlnh6TIxUziLIsbLBFw5VQqgOQuzQxFTObs0
3mdvpTxDo69MxlAFf+1U5P1x1X3biBtnSpGLk6ojzpGRmoukxdH74j4XZ6zo
USQH9wp8PHQHBVkYA7zczNjDivy7EAnKqCWYks2E0xrXRaFvCFH7bc91I2Ob
zjTr/xWJk3aRLeheWE9uxbwzckdrijYaxhW/kdtCxFkotMDFERJ1qOTeWz03
DVCNZAbeFqy7SpJUpGCatOhx/JEmf3uNMUV56/Y5xzyF6r4YhY7hJDQnUtfZ
S3hryF5nRlBMd71pBxDez4ugP5FuuiyHcZwfuh1LGgHRLp2KRYDjrzSpZTwp
8Yu2F6vYJ9UZO40qscOwbz1ScLxyDU2rRg6kYH3BV3RjiuAL6hfZ66U8U5lp
nKLdMRWRtJ5nlZa9nPgkX5u9IcIlQevYGqzQNeKBfNergCbrJzF3aZ/D6Qn6
GOF1vVhib4LDS4Wd+aaMEr1hDUaFTnrgMZdX/Y+34M1uyjgksyPxpDrstorT
O858W9/May2NGds4kqRctRmfIWecr2iJRz8iYYh+urQBlSSmfELqonrr1Gig
3dEGrHuZHGyySdfjgF9tJxGCmO1pjxlzkD1QZqWswmFKEzYkdo8HvjNS9o7i
UuiRs9GW7Mpk+oGYxMX9IburVetuRal/Xnxg6hjt8wfVcHs9mb7AgXDBZ6tW
vUozHXwQdy1F3XLtmOjLjQmv8uk4+KLVhn2Rpu6uebcL1xu4XcURY2QTGyF5
pR/olg37LmtYS/ON4QHhi6Mt/oN6gZ/1DoJFPJGIh0fdHrWcyt8nJmcANTm9
E+JuwwV3V2vWqTrEb2noewBsOrc67lkD9U0flOw0sv/U0umfEjWBSNvE2XVI
BtDLA2YT+IrGh7mg0ddt3vOXe1oNc7mAVz2qBsL2dHAI4YomSjgg70REMNvB
x/FHbDzLjxWU/QL9LPabATkw1UxpfnjLHDugdaLajQ8ekXV27BB4o7wN8OqC
MMkZ5ID16O2KS6nrIdPF4RESZZKNRVfjJAI0Pvniplzmr3lkNDoyztqFpOPm
fy/nSs2gLUbQ+T0t3nu3WvdBvUYVNXaJrNIs3oKXqC7jS+aSlO6dsKWJmslw
YoMiB4Es5QWn9msaJ2VWZqD7Wg3ZpwvoEJKJvv/5FOdeGW3TdNHWWGwp57Kc
kKQFei4kONL3SiEYG7oQXlFMiMC8EcUTLEr2n2Ar8wJC7PYPXhWXN5GrD7z/
S/76bvrJ91gy+8nCTBz28w4/9criAhS251gf3JlI0wtN4/aQM+N/Hgil/Ix/
MhvEn7dlpuABO9hFkhU/YSvw3ahVCcd3FFZlBKiEHJCklLdbTuk/gFvB+27d
slDfAYkZUb/TyHWdwryOzZWC6h3A4dwLLZ022CIFn9vB/b+nVJjqbSppJmDZ
XLu0z5uC7L9frprfPGPRr+mnF6bX1PvFGXyOi5hNvZXt0t9pQjTNerQhRm7z
9TE4y6cSXkl4y9k+KjCABAsUTSEUlP489yGjgm40CeRKqJab9dnM3QhfEkyg
fSmpJOZvd9wfnwzizfVzthyTOFY9t+GoBnJ9epdOb3X9NDlivC6Zlge9b14e
rd16bfQIg8emdkTm01nZEH9JDSGvuk3P18p5ORpFIEiKOCAuRxozg+ARaH1y
E2IP6Q+AW75YBcO+DwTfkIyxUKzTL0cdicjwJR0hTnY/9PqoZ+lpiM63by/H
+TrBzk8haWbvgI+kR3kDLlERjULo1LsegEoG02CiBU+JxHi/LI6Wfwjkut+P
JWKzgQjwZJ4/RmKKRYRrQa+mYac6BucGyhiIPqIHvQX//EA9IzirIDqYKpPC
DuE0Kl4kX5d0ujC4ZFcJBCcLrCLHxDkW4mcVYvrM+bBIviWnRuZJ61rTmh/z
PbPrje+UFV5gLfqiF94Pnrfen+Y7XKKTPE784/LDDTJ1Oy+VKSKmMyJSsn+a
pj9ccp+dA3KuO02XPVqVjEmL3YZXdfk+HFsj6Q8e5+eNGpaFTGngvtJ2xj51
VSxKAmK13VM5XFw4XnyaJkV2UTmTSRsqNABMV8Zvv3ttsVZCTZuzG6JqxBuE
O+RKKSR/3OlZi1FWf9GDZ72U0k0bJoZtpensRQpA3Tc0+fPsCZbSwkdC58Rb
CHf/OFn/kxj5YNPdxlKYfy3iPjLB8Qn2My/3fMmmUK/kBt/FV+7UwgpoI28b
/rlpnrksscH+CJvp1no3/M7P3+K/MOERLN6jAD5A809yIMhR1VIZg2sc3bFh
9tSuzdmizltcK7vCYUj/m0rfGbljrcK3xSfjL3odepfsxIGiJN1vjmPF5gXs
zHbnaYWfmFkna5YOBPxiNoJu4xGc/Rjd7CfCgbLufmcVHAJbFf5jMMMVSPyn
LxOnePYaKkwyLFcZiczHgLuXYqtFwDSl9UW5ZJRmPT6jcYb9ILuMFG6XDbb1
vrd/OF8ATzQmMAaMgTGSgdoxmlNFUjpBnQ1/KthPFsLF4s6AqBRHd+H3LwcX
4izqq5V5CYMAi5TJ3cSzzqgM6U8Xd470W807UJB+ypkyuD4G3gb3MTufx70n
4+u7uLuZK6TXukc4pGUrL4eQVPocHxTHoRzKS+DZX+4ejQITiaYrJIYQivL4
YpLv2kkGA6PJIROL7DB64VtCIryfzXrVqnZFsSsO/YUgJm2spG4Az/2V9Y2c
2g+nkIRDQkTglDBcs5WYbLMkwEgxJ+0nwQ0ES0asdGBsPedt/PpSdzhkc8Dl
f28rI8F+px5arlBpnWq8f2k8pVL4h+Hv3jfWx4reRK5CS7AW/t9KIY+BQqOw
ihaYsE/eVkSttvNrXjiG7juu5xf4CckQOs/QeMRXQvMIm5iakG+ZB/pIUtKn
S7Lep7aQ3LC7TkQtCpo4FWbAkQpnGHG0IKr5+mnhdr5r4n6TNf5lqfNCNBrn
cjJvO2y/XF73cH2UPm/r5QL81EflFtllDXr639MwVq701NyQYHh0xKAR+A0M
i8vAhEqaWpfaZjNC17cMLVmrTU/SgvWR4lSG0RN4Xkxr80SKLbHUug57Sx3O
UgULuc3W+Ly0yVmDGcMMQNif7WbEVOCQyzh/dsr0dU8PyO0pVMQcAh9NMuzr
IA4Bj7wSCzO/KwJvftTzsIdx3rm29InH9rTW/iS+7GQhNF8YBln377jVud4R
CznUSvCW30kZj0t8D3WmMTG8fClGrLsJIp2a7lJW6vKKNylW4f+UjBS8rB7D
JR5rTlPfgnC+tIyIbkBKH7xnDGnq4rLXJ5FcLB6ud4ShxVWdw6qGSpTKOkwp
MgAe5zDjvdc4DrNvQLgIJAgFpJ1om8IMmH/xkOhzVm5LrVz68G7wYoxUA7rs
u+dAoc2XodX3pYjnZYdlJIaR5GSKoxJk9YiM7Do0U5Q02QB9GCzo+irQuhPC
ePbGmM6wBeqHcD/J8Ec+r21RPKhCo+nBsDzO2rIDVCis1y35pO3dJ930WW33
/d6vcsmZCuHU8fcK3uW1EG8D9lUjmfbcES4+uTEDa/71/VZkxZyctFs+qvp4
XuzTfqgil10mXlW96uu/mXJpPiy4DKoFrmUeh/Wzt2s3Qz1axjNTezqhKzY7
rdqT9cSgjF7CYImn3vXtpuFai6H+EOWYAhJ5lO35tdOVYdN0kQuR+Vp+4D49
5iZoLc7R4K0xdO5NcsP46O806SV94GN8bRzIc9kaUGLJwHBMThhtlFVuUNLq
ry3DEfvv/rPPtrNpEtCAP8M048BTw6DoWJl6n++DfZ6cl9Vo0u4zUIoNIjPz
Om47f95lFKm3pRZ1226P85AnxEXGewxBjcasK6B6JAFRxM2Ns78f6K3yc26N
drguLgOSpqwi/jfY2sfBP6FPBOarDlxbT3cg/S2kxLuCroWiJYefoc3/b76d
kBH2yc5g3MgClFhI6Giw9JKUHU43hhfsrKJdsf3noReAeYY00MGQ/PTrePHD
hyaPRg26iK3cDlDx+MIQBFKb68tzPxPtL6k586d0WoXOOdXy/z0QnB2lTow+
o2NW6R6wDrDl1MG4ZRj3uAxJE6l1VVBE/tNdHa5sWz2dlOPTdbDHWQzkUVSN
qHT/g9KOcdoPC+m0z5rXhdrOoaY0jK4fJYKTvgHpoGt1vNr1R4hYJULZMZVC
HMcPIvIJHul/czoG4flEaNfSGo1atawMcLcVNGUpR18494Le8zaSriXfp0+s
B0mahn7AJblj0jivF+QuNtSwjqxX5Y8n2Sywf2/pU4aHMOhbbogHHitXMeJp
2hvt7FzgwKqKt97tq1ff5lA8a53Y7SGfqU9gCpapqUP585Mer6/GZ355FTO0
9fZx91biHbBkJ55gg06s34eFP1SHbn14G1PeorNsAoa+1QAA8ZgxXjkW4hv2
/itxvckktutvtFqAfk9j/HVo37Lf8m1InnBBB48TVtTCTxzfRGT9EREud77i
SFHCtifrTSAdhmBY5SFNIzQYlKXUKOsYdAn1lg815z+NkBNlGPYCG4jUBwwP
EbEjD2WYftxckTTaLVKs1V3D1iHItqEgdsmzj3GF2hl9QtJ7RGbkUD7qA8Rh
d/hoTiisXV1tQLYDBzRWH1BQkuSIIOTGgYz+BLFNHnkTLkDhYip0L+//dyn6
lyFGBNeuc8W8WL0SKXh3OiW7xRUDMXbiMh3b8kDX6eur5mvnq63j/6j8kvse
06byzn3h+DeBOPgdyFxL38XDJPPMHLVHvqoY84v1ggLZbyk0Y3jtiQFFmy52
S8g9FsIuju0I/wltMuIbvvftFVexx5dI0JOGxygerawdDbcsp5LKkqDZVlpP
kcgWFtLc2v3sEaK3wihmhK8G0YkZ7GBqwFyQTAPa/+8hmvDI7tXzlREuh8Te
5+Jw79dBMaDLZc+anpFL8EWyVi3ET6ga7/XY9Zfx1AnY2lGsssnnoOR7fxOw
mHmjNiZFZMgp4lUX9N5uEIAuKlvPZVIArDh6dWy4rBZLb7/1bVRkOtpMomUI
ZYNzyGKZ4BLJoriLY7Ywpij5Auo/ObtXMFhOteeqgrMftUHt11VIe9CFOZLG
ckHky9whlHdSvfhT2cjALH5yw4FGOnRzs/O/BYLbWASwNI/IjxpomKtgBzES
ON2fHlTorNZxys9USommDZLuxDmdkK9jByECI8Ueh1oHmwTp+wC4HMA/XqT9
aE0eWe4PigVu3Xnu7w7m1399sT0bHer/4e8emqsdXa6lrGsAGG+PjOAy/6aV
VLrGVmZf0zArcBdVYnhWhfgQDOq230o4/XJJRKv1UATikeEmeg4m95ar3iPs
lzTfxxwrVFdb+UNYqMcNtbYajnnNcz7AkfXWLM7CJblzdputIUEHv+9AkrWd
6s7FfP1rD89E3HKP8Pfh9cQPlLVjpL+2hXv+3zrp5KV4AtOwQdnJFU8HLGNP
CBnFeaeq2FA6+Z0+ywXxNboBhmwgVezLindfPI4t2E7S+8KnM1LWy7YlZp10
ZQJCq0TWmCoCAnuaBcXlEOEOIMGze9F7O69fj2MClfFf7cnDKehJNZXm4eKQ
JxKZA2oNIRkcHnE00Ti6xbwDcW4tl2mP1LyChz9ktxrihFrWo9u46O73o+/h
2aQNz49K5D3W6m6J3O/mgJkIQy7JCnf/xjpzszydYftMgGb368cUiwmx/Uof
Th+5yj+xpIVGbUO6gtoCS0NXh/WKtKggDnp1ZEjxDUZjsgskEGDutjfSHEJ6
Rk/B+2N89Ej4SGepEz87EZdolIbBIcQHRJblpgQDsCb4zIMeFP7HPygB5BRr
2kVDXbc80ezz0QR1uBNLErv/WnxUaF1yeWq+rVX13wE49WBmbWEBz3qz1L6f
T9TBkrOxxwnI232gqeGPovdmksJXYMsgxYfbjt8nFN1dFEY/9w1jF+Wah4KV
cSNmHmKi6uqsNIChXTnrM7A1mwHheAfQXctozwRmswnUznC71Uybia90xVoY
ZckNTzhcb+Ua4NUFBPRMwQFzPiqNWYBulwYOrTi46pln5i26pdCAbFszQ64g
pFZP45yukgGrzg44c+pu9JZA4waS8rcuDOeQVRFs1xrZkMWuVern+CA1NnD9
0xX1pV9YHL0RjPe14AmBRh3igmx/FeV6WKdDt86rGfWp+INzR8Hm53Q/FCcK
GClqPVS8kWe86PVi6+MYNa+XxmXWfsIakHWgC3cNj5LY2HjlKGDZMs1ap3B9
PddkCGZ72hQimTHpxhEYS/qo4L+QBMYlFAIwPmsfgrKUh19VNShwJVaBcVBU
F4AdnKDBk/uMzWQyX8woSKKEr1eURDJhqtFy9Tosb1hZn/wcUJSL+oqQKkiq
lRMUfEiBfTJtigvBIkZkX7jF1y1k48KQ2GXPqzKaowJ8Eu45yms8F8rjTre/
ntIP0MBdmo89he7ZBg57WfAfO/UN/g0NRr9JyR8WNwlVdIAMQ1qvRNgSAnh8
7NtydfxM07AWCYcg3pRPJvsGhBBLM7bhogr2lr3GhT7Xc2fy4CFR+X4zV/s2
LTKPIRZaVUMaILu2TYOKq187ZM5UM1rxuVuZ4xOpEC2ahZBgFPyK0ba8XdUv
9WNL1HU/xydUOZjtxjA3TxRKYgJnFoK9upyZj6JVYLOn7PTUadZCwzfZUYwx
hw4tjSYjJFsg92SANDvdD5UZboHU3Li8sbFpL3+MUSwbExbkMgdbrV86w3N9
+0zdOl7tbpSsm8BCRrP+mloCsQ1Cl/ndOGjqJztIt0ZumNzb9WXJ/1mTZ03f
XW38ybAIkV1uruxmL3x1CRrDRhlscXQB43K7P/Gi3GxlCzSKYGPEkxnRAnjK
hQmCkl/cw24SNMwDlBfUt5/XITwxMgZh9aq0ci0sUExEj5jcEZLUccSWG5Mo
nTJLZ1IqAhSGl4hT+HMprrrOTJV3B6q2ID12R/lC8OIzxJOibLZQv4/NRXU4
tnb9BO/NAw+iGgp6So3gsr/ACAdnRxQNnhMF65WofpBqCnxtTOojjp6LSgM4
3TtDP9UYP7P3tmvWa/hNUf2na3dc0zDKS4buwXyx1L6icICipGAijN26Uv9e
9LjgPkqUhTm11mjE154pFFUczQkdugEQy4VZV0Qxma0UJhe4vlqGQjtM+nnX
3g3IUt1d3sda368gyKwc6CN5oZbHSEQ6iHfOK1JdhVSJOkXnK2mQ2uyzLvz3
hBvhVXEt8LeQNVhdMZt5IpkfOLXGHB8HgpOmBY+MsqdKWEn+sztK6SWsF7dP
cLr9j5MWZHGXSsZxY2ushaTAGeU9mn4AK+Dg9M4KX93kYvMwhCeL8qpMY6IH
mayaBbuimtcYNw6jEMZ+PBrDvF3WRFYwQ5xyZ2qvWX51TJxN2N9VoVp+3SZo
jvG60Ki5eoMGMGr8OX44fGfP4lDWZWXPdIsXh+t7XDZUmf78U6UBCmsAgfEP
ArpZPrXvGKF9IFGtHYSdgLYuOw93iSwSkdji5DLcDsdqAx7Wx8Zh9KyeYsWD
xDONHyfZ6JwXWmufXfNtI/3KX2VrTmaMrLM+vH6HeHJcBuy/jJWLihAeloBo
Kh3aZq3Rc4wv4YLYaBjYt3R4jsg85PAoPTdiKIkcvkxcd4/Al/9VKIVaSJry
qrI6BauScT14cRQE7EOh7wcJXSIqQoZqL/X5QuOIfCR06YMBTR7LwS5LOaa3
jqpXsSzbg8UY9jfXzezSl+cBlyxljR2Vq/334d48AC3ArsXQei9ZL6OTeo7N
AqantsC6SDSwfbPw5bbGEed76V5u2A1vREc2IHt60pT2jN5KRn4LqWmA/AzG
L/w39nQRCmJdRawc+3xQFfm4b/L7dbUjq8ySDkRN8VPtzALLGL8vNQpNhLqG
OsINU4L0gCLk5be1B3Q0zaYgd24bPorVg2rxZnj3rs+qi/4IlCghtVwqLuPJ
ok4ReN3O4TP0Rep0s7blsh0KAKBqb20TtvwbySOj6a0MuJaw5s6cLIxV/DbY
7+nI4ABzkpYHFukuz3v+FJl9yswHGm+pmb2ohfES992Ile48xOcgtyDuLcPS
VUJxx1fzd7l8/kQqlQBvZWlonhBwfMlDtWd9mekO+ufpkrjpkBfrvC21goLz
8wb0UJuy7W8o2jf+1+2jUBMtNBzcoE6s570efcbPfzTDtaGV/JYDYHh9M4mx
a9FxbUGkMA03GGkYx4K2tqr6QzH3XNmWAipUe17F5irvpNayLixinS8SX9EN
5QCbgSIWko57c73II5A8aMBZtmIXCFUnlo8+9UksopWp+P9hRM+eRmaE3OfO
NCR9hobWf1fxt/SQEoDMZPO2gPAreaqdVhEozMAfyeyVhm3FhUPfYfHuAjr8
V/dPmXdSP7Sf4KGhp7bc9ucK+gLuerdtw9DaAFRoLfSQay8VZT/bAzs0iRpZ
i3s6t1nCFs3jccERrwmyxf/McT381HCnqgJvMqQW9cZBePC4vs0AmvQwHR8R
4Oe7Bg8HLt+VS0GP6onOv0FXGBO/vhfKhWtahtmsabwK5Kjji1wP8tHIvxpx
fn1HX7pAR+ohde/8NW/UYS6pBmZjAhstx0bAVylrLA2I8UdIGGOKrIJG9EPZ
owEL+OITs8w39CqLf46E9LCQN8488FD8BMwUyfBX4Qi3FGK4u1EgtBDzd/EU
Nk7qMulrJQHUqZgUDImZeHax7duyhEDHq3fRvrFGgsjqwCfn01g6f7FuUW3d
UswD8/nPAWFH80y1NGSR/ZMXED+tzl1D9yeicEwUdwhNmnxJ6kkDZ5b+WHGi
xZx6DAxZQz3KfoM5Yz5LQhHzMHNjdgxNIY0FD4NuF6lKYPrdYjLylSMopnGF
S6BKR4+UB91m/eT6vuruo72ZjJ/fM00D7hxvJ0712gepsqNwlCPFf7pQTRJ+
CIDLfJn6bnVIMlsQfwESa+PMx3E1fM1tue1C1lhT/KBPSMmKj/ow9TmMM0ZN
lrscpnNZu/jzv8AykNOvW7p+EkkE/8Z13VusG2hsrD2qqaVhKoPIwYV79hOO
gExf12XL2kTGIRGEfGi0wT+K4hNSgmw2yPzMaAVICEyjE5Vrs6pPQoBmaaLI
C0P0CztQ0kV/Zw5CTLVkC5dJNCXsLV9h+703jGGlVLbOwIHyuARmy9Shcb8F
npRjmtoplGBW5mXcyXlXQzZF4NdH09IXClesmAyKi/2DwApv9RnLS4ZcETSR
BX9vatMQcGoSBDUbHz8gsoyK8WyaG91KbkZY3FDkLF9mhOvtjmtf+wmV0SzX
IStqXx55JkKvXJEViXq4qfbyp0aw7YG/RSyCpfUVi8k/VKn9jv1dmQwUmNyu
Z0Qz4FyV85GM53Bl0XgXMAj7tar+xSmGHExPFRGBaLWXvSK74fxdRhWX8ZU0
XNObNr7dzAuBJoHetyHJdO81VHbGhVw24FQfOZ1Ktv0ZLEXJJs/ZRx+zq+Ar
YAAbFh9BOE4WqYmoQ8otu4vVXkWbfqjmsA2U8nMHuOoEnTBm+7OjYWuGRn2P
ZPb7DmJtALyuAqD2xqRPX/fbLAuuxHf1cu7Vm2duTCtE7vteenLKIuFNn5ME
hK5A+mZG8vP6CW9oeOxJuCK74Kgfm8kWhtaDZIjSozjxfSFE2v0j7B2hBRQL
F5LbXA05YyIVGuFkx6FCzKewJXthGBU5CkIq6b62iBZnwCiYmn1MoDpuuYhn
T2JZy8Tnl6pSUxDK/oe3yJsykzqYQYqNyTVW7RCBRGfW6eEkCHexoN7rm/Zg
ihMm6ZRn2AbvTnCk738YLWuJoo/o7t6UKNjknES5BoJUDmEz9tc1ubGYEE8/
loCNljLas+ACNw62SurDV9IY1n/pIkXB69Ao5MEbBupZQQotjp3l/lVmgj8M
773syumZe5BRkAhtXAWlwGRy/5hXzToZoVf+H66fieOmctDLhTfI6czVS67F
9OaiIv8tdTz3Nm44VoWKBTh02H+8Mp8vJtkUxY7hL/V5idVuyvwq7ltYPIgb
LDhNXXOqmaeQWL+smZt3IJwkiLbKR/4rZ5ywydUz81kESDOl2mfKuh0Llw6n
2HspBYG2np9NbzWaLCsDiIJM/IAlnRAmYjAuxNj1Nb7tqi1iJ8QbEd2PrYQM
gN2QRPC+951rLLCxwsrPeO8aVZW6nd05actN/YPew+/0WgVRWtPdRsdoK/Z4
JGHzgsSsdRlm4hjZt5uOw3ZghaeaETOMVSNB4iE6LleFCNIZNpTZSk5tUPaD
MYlY0S4bTNu657TZOdKYxUEll1PNPyZ9p/sxV7Li9lS+Nwyt6g7ob+E7CWfN
PokvTfm5SJa6UknFQoRaE9MpQXm27I8aHxkzfE4KG7jUy3HVXbUajmR3MADv
fMvfYIjZQy1kYkqug7s0NIepfQS7N2lvAztmvdNTjt3GqcHI1lnzwrvAz6xb
sL9F8rmkipLCWtoZn1Y0esbhsWUs8z3j+MXp5UEyDvga/WrTJWAeORRWljea
CrVS49FwXXGHedFY5tQ6oqZ5ZolMdgEIMRgwcs+6zofTu0YRTIkAUbLz6/kT
uKFTcDbywvRBZJ2+W3s9H9y0zthZ76QrWEF2YqGbpCt0Cb3cLznZ9mz4R45v
3LNA4w+trRpRyo1wm4GscPfCntZZLG5s/5OAUBgdJMwjXdi1OoqUHLTjcoXv
tJ+sk5HglHeU+VOSrZnl+mFZ9wPjQk0oqhfubjBS5UzLgVn4MfVRQfwO+3uJ
EKSWdh/r0Mi+jUbZy3l1gT0SMuOSld6hEoKwMt0OsIgaOc+naDjQagvluPSs
Pq25J7QjL9am8rpUQPO34crB5F6N/miRque2GaBpNZPmFfdV9lO5RCpCJkN+
CypXT+PAabjuempK8c9KOnzjGJrlfYXPnDkYOzU0Mw4DdmqX0xvyMP9l0iho
v4eMxv+45ZLl3i5AVn6Qxt2DziC/eTNP7zeUOUEXfg44on2M1bkycTGr7kvb
sKJO0Ye0IP+3uNSNAxAEnaCQBpCLDHnPJ+sL9cA8vI3HZedidTFnXJuLSxzR
nRgqn5PwymnC25BTZqbbi7JeXgzYkyN4FjBXfKgCrkr0TO2g/eHzQuy5Tit3
tE139RifcJeExLLNlY98mXA6Z/dOFD8/tZZi9omzhMgIUENDkX/m5hU1NhiV
Rflcc+0T4oktOSC+kJWiRmm2vywliVRc8jiBOu8G4OCc+tva/Rvzh2c833/P
C0UVL2Z1Lxu3LT0jFJbTo2nClawOqcmhBEjXok3NffN0Brs/95O728DnOgk1
fKpt0SdLNhMQxCtle4+dBjXxYy0/Qx97g2CuSoS0hZiV0okp0QmhMleWwjlN
MDT+ZMBY1zHfMy/PWL5UR9VBnrkt3dxbMBtIynOsFEfd7ezXh/2HcunxSxiT
aRn5TOwcmJ8UceXCDOGbnZDmg6XmHyEizKHh3TRHSOik57ZPuh1JNFGBYc35
VY4GrrEDtPawXrtkt/LSko29IB+OA82qbmj2ONpR42lFBLvhTZAwLmaMGT/E
ZcvZfTP1BvPmFYXLNxNA1wyRmbslMI0j6PhcsZHVRekouxXwi3K0jaa5lU6Z
Ftr/dxgTcAvVT/6iyREo7SoVrR+kiyicNgcNO7VaZmgLbxL70tfdKw2ej0eR
z2eDqBS9lu9zLAExIdalZkT0xQg2EHiTkE5Bq0azdPT1KRXrst4atC+NsgyW
egK7Nbe/XLuPvEnRkaRYWHt7RrwUdLl68UxSykUjadl0OzI4MpMf/LONocjX
6ImjSexGFUbH7TmOL4LrBA/mAohInjYbRvgyIlW3a5Z5d3xORHm+UzOCHDyg
YFKIfkAAOep95d3v4GQSYY43uIp0DNYxbcz1j/Y5pmBSsk1+IdbEsgCXVCqR
016r75kyUQElre171rVEFwwkswl/pmyL9RkmljdeFg9DRGWZIE8pngdUYI/d
Dod6i7NDRlqLfMLKBqa7E+KrioboeBjFIl04/c0zdbXz9ecfhrXsgMDrUNIv
xxWqHnggIpEemKajWNJ/slXQjVqtY5YUD4eELYhk69o0V0M9MIAQPvPl2cd7
4lTfKwr3YxpjqEOzp2UOU3wY91yHf5aumkiafBXTwE63ctFAuhlvSSjSjxmV
RvvKsNo3eV0KQuk2aavMWJLt46xPgBXcLyYF5aMcvjQrlfFGtJ0lUgGvf9c2
o4vaneuJyFqaab9KkS9y9Nl5ZUeQ3CnLukBek+MvO8/R1gdVN9kJYlXy4urF
uKcAPEL/pLeCpJ5dOCHd4PrDNiYb5EABLXOD7vKZu3c57jKM2ql16HIqPgVm
ZSHwD+TtAJ98603S5Lr3oyPUPQ3wmKxv1akXMWIuf/K8zPV+EmVsA8JD4giv
da8wx28Bw35pk1LlJccHel8Bb3DgeqWjcbTFo1xhk7iIA1ImgLtK3nppdxNw
zFX5IZfGZ5cTenLAZGyjthe/inIi++WNGCxL5OezBsbytUDIQQ+WFybZ97mI
8zVE4F6VOaBh/Boz0e5ldIAmXRieDOdT4XtKerg5KwzKoIe11yltE3iKlwsn
kgP8GIw4c0SEEn+qktIps7DjIBWS+2FcTz7s2TjuYCHFNxHVNDShkck4XkI4
GUeIhAUE/4pXa4PTamJq47AWpILYaCx0/N6lVk2/ewMhG+3+jrY3snU6Pqsv
GWkynPd4GB9culAuQGk/BFPdQeA7cHhwC4leWKyFOpuuBbfhWlJELyXqGJR7
HO0XZyrHfOuSDh0sZZ/MU7KsAp+f7mlWia6H5jMnjGzcQhKvrgWOe1XLaEvI
UeqGjDLvWB3QeogZpDyLSPK4KfupqGVvOyqUJX3YyjeB+CC2EbWhtxvrQ7fU
pzIR74nrzMuxuON8MdI/lrdqweEwEGBislwfmklmPk39zgP9AWBDOAAAxuZH
dIUV2topf2+1TAcMtIUR7t+Hkg2T7fWe4PSj3+QoBmeHJZFgLFf72mtQwKzs
0gQFMkSgAIB3eMYymeZJC1mw4yMN9YqWOsWpQeR+buCLtz4ZDPo7hcOf9LQD
lQtz8nITR+i4Q6NJzTY4zqzIT9nhNeF7IsWelf3pcafW9U0wDoYk6VAn8l0j
G4HStCVRX1fv8LQPYFtup0jnx5XJHMoPAvKk6wC5eSLsoZ3Ox01Ne8cy8YgM
lVqbsOy74biO668oxPc++KfaO20LKS0AxO6C7s9JITCHBEBbbepdIKDwYH+y
W8qj1JHkRAD/hoBY2f3CCV63bsMBQkh1kvzImsp4Wy9IySGjAk4q65VlRqmo
XMloVaCoH3YLsWw79Xz8NgibFrbd6dQFYYw/gApduTlGhC7dkEC5N5FzBGnd
nOPQO3a6gDnVkza/wX8QUFHKv362bubZJgE5jEqz1as9ZIMsvmjFyzRO/gd7
qcNl+I/WEOemTmJdDk5nsqeUenyYe17Xe71SmY8MYR7UBoBBFtnub59VAQBh
sEXVmtf4/lXQNqiO5k/Q7I666shxVr+ZaATFoFonuYhNKNrNw0zH7srOY4JT
5RIwXzGctCvjdc/5K0sGSlj1ZlsyuDPaW2U0aMNHTubXV8lY0yaQcFGNQTPK
Z/QAp+vJWcU/xaqbTE1X2D46MNPUmaea4O6StTBYBiQWQA6Dp3eB8cMIDuyU
iXshxRmJwUf4QN8kYlJTYfdrH8Yus40Fci7Ylskgh/oGF7GrTnMdVvBSBISy
RbZrCtBxgANj41CCPHH9zmTgQ8GjLqVN4XjMcmHBNK/e7bbM2lhg+UNW3K+G
ZbzCQxI52yVyPXN06ScVeTNSBCukI9040eBHYDQlrUMaSMcrb15bsnl+kO3e
J/fPVuQjX7hQUNSFkjpi0CVRqu7ETVNM5Ocf7ZOKEjHr2acjfOOY5vx6EHvC
VwVvL/j+RfIia5tmsbxoFeoY/bVmujNWd8vEncDCg7y9pZ+9rqiYelM/KRn2
no9xklNpre1cy6xhuPSt0HOzygIrHpnvjPm3gRAxbVHKNlrlPkJCUqmi60pX
FmDT9gq3ZjLHjJs9u7Y7Svdbw1tRQ0u9geHtR+CX6fod7puh2UY/WVh5eXW5
Ubv9hKnFHUbGMOv/YboH3cMY1R0g7fEWoZJeGIj+6hhTiuL8dZiJULlbdh8h
TfILogj/wd+TW4KaqmIfsdo86XgrezRqpRZISXje7Fs0I98v1bESBL84JbVl
1fKXQ2/YJoapMdawfbHHVc5QOVdmS+Jrzn+UYgcS43NSwaeZqI+I2FQcfCh5
xnJPO5GNXWWX0mKpNGfFYBif9epaASaQzTo3H5lzqLJ1TsdJ+zWLtTyqcMoy
mv+z+Oy50O+nMujU4dW3eFBsrCyahhnt90OuJFELvz6uCImnaI4lZmxug/Bm
0dvHHViZrswKUEnIIpBWKVw3u1PZRxGbksy67Ly0+0Tpr9HjzIdXVbqHXY94
D1AylPofn7HKkVAXMNIEjGcwTPfBa4Pfuc1UdZdmpyi5+5p5ALk1p03SbqTu
2hyK8AfIJao1GiqqVNBOBG500ykaF3ynUKpT4dHhr9HADuSktz1sHAYVcewe
dJqYYeclgqzM2JGbxBnfFVjniG8jeOXJe86kqVNcDb6JpiNWkauMbF/dRmU+
bDrYS6W9TIXgkNPmkBY7i5ks4EZr+S7gRJ1MHnJTgKrGYWYdlFVj7//mHURV
IYRkH/KIIM6770NoyYx06zE6qHeJpEmtGxmDrR/1ZLKcSYIOkhDU4z+U28Uo
y4uPkA==

`pragma protect end_protected
