// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HoWqUxy+1ACPDMRVexvIwt3MClxsGLNOlB9xHyEQUEf19Y0j6XGSW7vnsdR9
OK+EBCg4rCZKAzkt6Fw9gzXENQjh6LK1XwH0/KQ1IGrVXSVt7+rb0QAZtrJb
tTbUm7f/BscFQpFLrLyryTZGIhI3Px7EhoJhr57P39wxLolFXgf4I3Pdiieg
651GoUpOgqW8BUzE8ZyctE03QYNHDmCWQPJUhY3D7cK8o88JFHjYrNP5EUO0
I+azzAeLkPNVGosSgk1RJ+tWIyrMRSPFmeZiwi5FIRq21Z3Sj9oKA1+TXN9F
T/PjiqcykJzIDC9INthTcAU7ljKicdY2hcKMz7v3Tw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W3vgqbeNZ7kzyWeEyW7srqxVykSH+C+GDHCb7ntOR9Pjp+WrIz3U+UkxjTbB
NXk7h6ASh5eDNcWMQy1t9S3k7xBpvlvL/Ia7plFwlXeGelUXfnsDi03/zABG
TFiAWps/H7kCsfa99855eYnEs+hOnMEhS2avhgvx4fFmN7M/oxBWXCYCU7T5
Z7sWgG7dDcsSCCNNETrlprEt/GLzI+Zc/iacHELshyMVDxSY+B2E9uwYeb3k
7qnR8w9Y8ljN6KTGU1JB9g1oYMjlzidtpqZAXjGjaSyFTr5wjxvRko7BNrJH
LYWUYEYw5OQKqL7wDP071cTeDHBzOW1Di1fq6IT9ag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IOzxF1D0kG0dTl2d5vRuKvNQ6640w7sQ2/isV/kUV/JGtisZe9AaGEn8RyHm
MX4yaeXz87xI/iHYHGZe8HkyNbbJibhpY4xCj/hXXxrJtDlddg72BxHOYQX4
0T8040BdtfsgBaIaonhQ7nYk6CL2tsa4uiY4j/QyfxXR/t/V3sViV7+O0vFH
ypORUhKbIZrvT70lGcfJGfQhBNTz2WwBqCvEqMzd6KQRrH6HPahGcNRc0Wrx
v+9xbolskILnZ3Tx+teX0iEq8EFoalF+DgDFIIcl69bVi/bruamUGFct9R6D
DoDiLPlezjBqQzLUYIKCN+S/KpkxCEXopuPLv22ThA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pTK4ASMfceyg39/6WtGdJruAKfz2xsXIaeBte5uIKMpmB7n3DRN+0TRCG4yt
OQCTkgXpmIOJ4OSqQF7Oiemgh4R9yzxrald7LWMmsh+/gyPdYBoP1Csjk7Sy
OPObER7HrV1Yxg5/Txs2rJo5v40Y6RjVY8j0zVmHBDinmXzF/KQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TEaYZWeIaFFp0vT4mutvWTY0MpBrB7PCyJcLDHCEnQ7OrK8kq9SMobyIv0Yk
L97kf6/38Jp+s2XOVKT+7J/ebALFkQZ0Gs6hQZWb7RBy+pkQCT2yIE8nIE3x
wlYzDTcvF4lOZS+g+C/uGM839YpzUP4VmQI94lpr2V1iU4Ac6QfagY+FPHNp
AKbSiMUJLi8vt+fIkX4F6V0EuqWViXZKabjbf2Wo93hQuYJJ65QpVJiqZ8Lo
J6USQ4LmOAnJ74ghwqd+0XNv8DnF+Iqkq8JCj6lJmpAc5TyFBb8pRiy0YhsJ
j5cO5CYxRM/7TkHdlbmKwmFQA/Q+52/PFEWbarXp1afYUksKIrOBkkekj1Xp
wJgcVKypNqhfYCk4J9ZUWIsEM3tNk9VDRJ6jJJf+xB2gTaLug6Q+Mbm0aRfO
Oy7ISJ1eyxT2DVA3MTT9CGHj3yqKu7BKVLumN1z3WEqZtcQQHPg8Az6pxMUQ
Y9h/hcNSiRqWuXAmPU3Itnos+lBB343A


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
StD8pEWloWKnyEB+7otbugo5ixYkS5g/TMV4wd8r/MxrSBiMF+TLNlCDzCNa
fv1pFTDv/04yvT2yiAmAY7dWKiq4V9sGOaXc3MFOofuVCFAcvJ0L0KnKicLc
LLp11Xqs26301nrYwPfMnkc7mkQk3e9oDXDGmPivuQ0gwlrR0Ts=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
USEQS07zMc0/T1OwoE1iTwztSBdpVSxTlstCgtxWH6MwxhzznKyrBylWsdTm
N0URktVEONgYbbhJrIWSCzK5qdzaCHRSlJk64IsocIimTf1nUFafTioDvw06
fwxw5fTzkcCVP6SzJ0Gno7YmZJSxUBJQQC/vfIvU2EINsxABdV8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
Q2Kp8zqpIDiiIFrUtPYUFtdayAADdJrALDjwRV/WdW1+sdBPOm0uZSeEXc86
11NsOXQD4D4bJsZ3BhK4Z6Q+1bomJ3elYOzK0PNeoXMv6pWO9IdCYg7Q//sH
9Pofo2SLrjLVqIT7k/CshYwmj+dIh0CjuBR1/B6Arl+HPL+qG7ou9J04edWq
LR7Vva0LngJO6tsO8FF62nEq3cbfCoUZnT5eBntr7KXSWMdprfhUKshfuHjy
QRYC7Byh+MGuhUz+X9FantWOOVl9tpioY8o6TovpoWrrpk96nes+Wn1AEc8y
oQZBA/T2/QAWijtSqK/3l85MV0Bci2JpIJUBYka09opTk5JuFxUtV+MkdVg0
SbXrxiFStUuudZBLtyac3CpzCNaHzU0kAx06N/UJVez3t+Yucs/alkI/jvjk
yD0CFZPX+L2tF1ApvE3AXEc6S0ZB7LotH60y5xpC1D4mphB1wtNBG+J2zLxw
enqsoGHW3Hl+gXOmKYXwtLFhgvwF/OXxicGcXiHXMzZCoxypzDwXakYf4jeu
35J+nsz58zso6syglek9EGIFRnacO9NGlJC2kA0Y9Sh8diJCkSxytG7RaFL1
Jnh9gOyJerTqkLwBcyVCbWACH28wzL2XdlgKlUBxtL/2wczzryD7TpXov4kO
zrMKRj9DviPN0vRrhd7XUzOUcNYRtvm0P46WkgnojeUvlq6Ppis1TRMwUfg0
bsdmtN03nvCRalnd+M2GnkzLq1h5ql5vzo8CyZht9KKwo6PUqdScyFPHpRt3
igseEz5XWi16P5N/XzgwCjgbExpN7D6WB9HSr1Ce4hh/sGQz4/8LKGv+vafV
XmEYkks5lgndyY6AWY9r2NkvjD6z8YOi6PSMCT0FZ44nQggPXtijGdOawqZA
AFDtmnuuSUx9uug+EbNiPyVh295gfbKzbSlPb8htTuxib6iVdylAjWib2qxF
Du6rs36v8wNv42i49fpQeTgtzUZBqd/FP7ZNcvnCjGpj1mHiP+EQZLzDjrFI
mhKMPaY691qg704prNcLFMpWHV2rdsMQOidRL2ypV8TABazzNtVe1wk7S1y2
8nzkyn3rRCIEU++gBVxvvTJNjOcL6eUfwiAV/xXV210t+smwwDlAnMkxIl0h
AYod6ZZ0QsyjAMenTMc/Xd+t5Ck4C7VaO+na3s1gTrwidCh3COv2ZnS/4ePE
8zuW0AH+uaUJJumhxkQxCYsI3xgHXqAj4e++H37FbQtgO+wQqX7+IuNjVuS+
GZwBL2usDSBEgctJ2ytneA06zT6bISBk/K2mQmNXgHhr5gftQZni0nZjRMBQ
WvnSoABR5eWVQWmMa+fHxKXXFpsai8xOvo4C/FStwBkf2tB6Uwb9EH9Atkyb
ZCGlbKSDD7ZHHnBz+rEwrcNmnPT3gDXvS6Wg/3Gq/rmUbdUw0XPmm0O95ZSL
YUMi1FBfPQJQNWS4vAojwaaOgUZVpjaxQggN/GzKCZ2/64cQyTkNC4AduOYG
edP083LlQEsoBSPKVp7eYSHsgJcXx61XQlH3ba3yoyacK6P9JgTvaoMMlljq
UFupablqvSgNH/sBqCnr7kMtfjCdaA2ZCMu9vGuAk6m/pmcvju0My48/TLR5
Q5rHufYptd3PXc0X9qgblmVfuVA0IPebGKet2Hk6CDCDIzz8HZRRg0cWPdHg
RufDS+S6/uOu59Il7/eoQvoAbw3iLEqb4SG8sOH6L/fCssktHUjBiU7u5jnd
Q/SPSpuyEbc76bKWN/6pGHlmIZYlAeJ2XLpUrnyo2/iAwxvW8e+WCZTsbuqI
0VZTqU6H75bwKnXaS91apaFsl7JyPG5w9gE=

`pragma protect end_protected
