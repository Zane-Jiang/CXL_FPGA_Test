// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
4eXeF1lVSXssS0OV4TcYlDEx0xIPJJepW+jUiT4RohLTmcR7AXwwYQz41lpPqn3w
4u5Q3EpsuVSO9F/RVD52GXmW8jdxQXAeYxbmk4za/1gwLEYjNj1J+aBGuzSxpFVQ
SWjjq8KtgM8meZ0JiB5bNMesXIEk9RZdLvzr18vzLfZQwL98q91fQg==
//pragma protect end_key_block
//pragma protect digest_block
LSAO/wRBobnPY7ZV5oalAB428FA=
//pragma protect end_digest_block
//pragma protect data_block
/YVVDE9pqplyEKANzpsfL3Uc+NpB++kZIlEZJVW7mjNGCe0mDPqhCh7davVb3Ogl
1ALPQDpYM1UX/XiQIAZIXIE1fF2njtVUumdj7OTi5nBNPmfbWq1wDE8FB04L6nE7
JEmZelKLJv8pTJX0MNqCHcqHggSJ2z/7rCrqDQE1Bv4ID5GPgdboVg5S7ZNZTyXg
47FKpbLeIThZJbvnVyTwYrYoFvAmZ/HIebc/RAF+PTBRPcEY2mm0I8nUF32Zl9uP
hVKdnPG826D3fOwI/YyenHfIR+wXM5/Xd8VQR1cqLaixUKHRd1UeCOJgdpPtFFM7
5guh8aPnXDUExH+LFtN2mNCvixtR64C/FfICBsPfcVbKheTXoXKfRy97JbGbWwbP
V10a+FcAx9Qct2wD3T5ynl6UCyzngSC0NMkpzDWLCVqRpjNP08kE3RjlWrIgqR0S
vpxT87wAgNTUPX03As0bIHzhK/b95i9/ORyzpfuBwdeP7hwHJw/HuYfRHb49ae/T
f2x+LT56cedEkLE9OXtz9/Iixo78+GgKKh0WtF09VN+EPByUI1tp8W8h7/5l7DME
a00XPn29yU2e8QLRuiFS+AqKL7xhjxZUm6R4ky5TiJLtsmkE7AgQcWBGI76SVotO
QQhXvKT4BQMJvyDO3Ab1Hu7x4ykFCU9WuE80ZppmrefodSjxjm+12HYfzs6Eeu3Z
62Kvw6HaCsgDnVPY8QTBGn4eImNhEECeWTf7YG6KmIRxIlANxUUeqpURlvLBfUDc
bHZtt5lk628TI6RgAlnaLRGdegVc0INiKRpnQ4jTzH4pP1zXKKGmwkweBlGijyyx
9+vgg0ZLYw7PIWd00T7wijXwahlgmsAtNgIIrf4MESxsMLn0VPjp5L8D4fLGGSwB
rvyMVnHKe0YVtMyXJHJatYpUbCgt2lcSp17bB5tBMNmrimaKSwWBwDdC80Ci1iuS
nv1aIsGjHsUU7o0T9J5RapgEW2TwkX4hPReBo5QvR1zmWxfqQqtPmfSDjGY/dH4B
LPs4ND7mFraETDzIFZeAsi24XX/3IbnIbowkVlO3x3Reu6TOM7MvthhbnMrd6Vfx
H1TEK/bsdauqYBNg/7/qU2EkKixYcc4B7LLoSxQr/AAsF8Bk3nZgMkw6IF9ELaFj
nQK+ppyPGHyIMY79JEHtVTiak/OQ7kD1NgVJdBZXM10VBkBPwuGC4An3u/hcC9NG
0i2s2b9+YHH7oYGtVi+RQ3VtJGdrbKlyPaT+HtKZDT2DTK/8Hbr5D165giUHUHeW
+Imd6EfkwTiD7emTPmWN0RntvYpIoOpEMZ9m6wndVRTmpYZK4YO7Sfc/WbaMTdaj
XA5FUZsE6N+iWPD3/6mU36UvTKnq8eUsfdZdbhMAZWOeGPdks7NhHd6RJiieb0S3
2BsN4qb6qhuQKYUNP91XKounobjOn5ztWUMXPEFVcPfWVkBp6NiqjjKSX3T+725C
K28jPDNfM4uoJKxi6OJ3htbrC+kMiv5ZXEg6MC7kIKhxm+SRbFTksOoqHccdWwQW
/NSgVUAcjVIjGxm1L1vDeal17PJAZB/P9WcpLcO48NudSjW+BF4axXCB9twDrkFx
oJgsbhxgj0AqzkP334JVzrOaJcY1q7wonYng1vKvSe2PTYwUG6JqJOpGLV34jJ9B
5KMzgr4yL8GkVQy0CudOu74c8qgQXuvdfB0J4elWhpyAw1NiNNSIUXfwL2E27w6d
pfq+I/qg1H0J9SlS/rQb48ZBlsX9HytiNsk+ZIblfgwSAsAZUKHAQdmO/rE3ZaPo
eJjOD9n33OBcbmpJp4WWESP54dYOAwZfyYLjC/FbY3zaN6CukBi2TvU3d2NIJ1Am
fre1usNsmMsymD5t5wLM3jqbShbVmeciHIT1UH+D093qiTvh1IbpdxS2ltdqzDSW
4YvKsUxH/bL5mLIotksEf3IkUzCUsDXtWN4Q4FOYwek+LTdCwwWGiGwzwB9oDYtd
wUb/CZ0HZOJGfenAtbkAs4FgUG15z6dapRX/QzjeLFmGyl3EarE+oeybx8u5e7vo
DtBtFQu+7yIGU0zbRofxPRo9s+UJ9ytIb+IgDvOP3BH9nJAs8JqgagPr4dnnQcRW
LyMi6kBy+uTmqkRjqQSVwOUvSISmbM/j4I8kqnePOafpV7BzHeNDNUhJ69suGZ3f
1PyDNA6AuGKptKuM4tfIcKmV9devXQmnzBtU+pz8CieZ+QWOtEU4qVnNOKcgo8D1
7tRJWhus3B0BzRYT/QJaZvMcdG145Cct5gaJZCuBLFeldd4pgbc3cQhQKBjcBkyZ
2bhptc4r5ej0KBzzDdcNTs2Ra4pu9clLROQeUJsgogSjOw5QlRzMIPCfVJiTvx8q
jYotCcrvcABnt/k1AMX3m5mqVRKj+wOwwTnVwBfh5AaqIJysCe64Pvtn+pkZVu/v
u4wShfIYhcwIwwG78YJamg+g+ueweh4SWdpxLXfN7LWBaKZE+6uD2E9+8FQsAa89
/uKc1tIiAq9r/4u2cUXlAEG8WcEX1TKzRu+ZZiHioyEREv60OCan+bTlAln6iC3r
AQJ/W1xE21vsTAZhnpr+5v9cN5KtLlXji7dKAwI7M2JlbSq6fDe11AO5+Hy0mg8m
RssElUzwh8azmg94YBx9LSDJTz7BFOFhUDKejk4PFXopBCSkLo3E2Fvg9frvAqB8
TcEZmhwpSocyWz8XF1/Bx23+dALlrYg3sFlb0m1zv0LUbLooX9TziIy0rSaF5el3
TRwGQTrRaSdMRZX2IHF+VwCDd+SAT1plhXMr7ZjquQvUElQHsT7Nx/7a50sioxp2
/8AcPCo/cXWRL6Z2MLmIiiKnYI4Zu2aj3fLIl+d7+QgCjFY9tnTPB23i5J3eP2+V
yFLPlR9NHELoOaq7lKYml/A9qfD5T+JfyAPG/NzbbS1VT7yUpyJ3ebsIDtd1si5V
OsdA/XVILQoTs1I2lX0GhWSlJDm75u8Ghs7PC1J+sgSjc+XaVahu3gQQedOWEjiS
aMD9m4lXgho2g6HZUtdswI9DFVx6UH9G4EKlmW9roEFn9sRONSAGpL7xsouXkHuA
xUU2dxHv2EDbQobP1CjEgVVZl23iyD9NoWjJo/C/cJ3OE1dn0QuFGWs63hRUCNxk
ZzYyBj5yFVB61tG7AE7TCmdGMfMCS45DxFce5JMN9p9P3VOmvsrLuXpXU7u82d+u
st3fAxc3585HAoekqBAmD+sarQGig7gXJEbJh6arHQj6VflL2WpUaoD1Vu6hhTQJ
e9HkxwPnFXWWdqDUu0AB2G0lRJOQjo4BvNOjpo/Cbu1NjDbb0tkFyG6BhHBk6F/Q
CJXymu37EN4B/pnNQ/pzN+vmkQiwyNKMHNzlcvG4LBQyMw+A+6+SuKQAt3oSRPce
Tnlc7dpDrYvqvr2EBMTMrwrsWNDKK2Qhy1a0zJ6K3BRp6vn1FZOYuTevGIXUK8q/
f3I6sGaFB3uh0v/e1NAJCfwaxQXQPMghQxaA6TqbfxHYU6G6mRAQich9/97MfYDP
8t9tpZ9p7movtMSShzb5t/m8qOFuqP97+0nZh5N2yJKPkNF2c8Km3AGMDurgXMta
xtv0mZDJ/WLwngxl7j+XolHRXX1qh8/ISx114mVRN5efVBHuUYcqEDjJ5fK7wLNl
rpBos+qGsDUnSh9rr+vEQYPNsHL778ly82c+lNDjHwi3Ee/+MzKqBWFrpKjhwQoq
AQkn4YGfvtZoGLB58co+Kjd1v6pS4bSjQXMZaYV/AaiX9HuAvj098N4C/w2fcS8e
2JTgDQvVY4Pto4spsybkjUnLwjwu+mX0XYOx6Em6Y5wCJg1NI57q/vCLB0zBVdwA
N+sKpqkhZZ0nOJUhtHvdCmxa8lxnQJdqBI8SEF08iL4WrFP8tO06WGouMHEHowTq
fin+aypk4e4KfdndiS7eLJ5dQiT0J5nhn9RmV2Q50klzYrqk5xMWE32j9e2rAF05
IHXzVyIwc7btKxiYziLXtVcvfM2B7WPdtrL4mNi7Ry5IRDsvvy7sDHsbvozpcQG6
KashYb0Y+/WY1RCbYfD0yDl7Ee5nCZrchadLd59oNkpa9Z5OlMdVGfsph5rRgeKh
+4qopoFw7sM9tAb4jELeTOGpI3eKBauOltwqlN7R8Q6qHLw/HgYSVnQmRxgAl2t4
fiWjYRLIn4EU2zZ9oWA6qSZ1gNnRrekDeokS26aAPy/XVahASOczSbDAQy3eeV+Q
bx79Sjpc9aqqx4uuHX4sOGjQrxY9oVTOKp/l/mgPoR+bTnBeNW96VaPd0GRU6AWy
vUQE9uu22escDRI0HesSzJbJ1KJr8wMskrb+oRQULMGujy3OPgIkoQLIKWhFTYq2
D2+Y53BHcqW8qPpoPhqXFC2D9ve+3pivoJEIDV3Bcl8pn/o++k5iZViOt3oSVszZ
kqZ3OIbVp3oAgWmGEBosUpAhJ0i4jxroZZkFbMZcgqiYi0YtGYgcltEyTw1rDPjw
5wj3de4t3Wi+S6mSzdQ5s4Kme+/mHJVQCcTUpvpGwxkvPcMfUlB8FRnyv+fa8hIc
6Z4bpOd+SY4iHnv/TfFKZ3RLp1YYGqR6ZKdcwsIGY6z3WZWG2MMhhmZB61xYxFVT
avdEdjuQr0E+am6v2BhClVsQsCaqKNg8aXa3w/pWCD0x7IrmVlWqKb/b2VYFqQGm
LNWYtZ4KXNVu58vctdF8+O6GW2EXII2i2/MAZwYD4hTqwt173AM30RENj1zVTYJJ
0xnFaMRkbH6iGAgIIzlr2Ronp5kEdPO5AZfDPpSw8hzNwAmk6AzZJybl0XdiJw3d
4kYnztu6/9n/pv+uqksn06/SL6wdL9rkRqtNbVjXt9/Q6ctGW7BDRZymC2eUa2UF
sTD8DLnZJ8IUTOmnnCBmCDe2JxLhGwWjJembQlmHXCyZVImzsw6Vy7xEoppxWh3+
n54b835/c3NlHbEGbOh8Au4owYPNoN5tRtvk2sSPtNQasH1UJbhsHv1Y/TRJQ13i
jIIOfHAnpLxtC8fcLEadhhFxZDBzcUv3Lh3kxkj9y8w7c0SvUYDxIvdLWHwA/c2m
M/9xszSkLQHGpqibikcC1DkpbChx/X1cFBUmmlSpbZeskQCgnvubIT0WbLjOqI96
FF10MmTacPH/dWAv8zOclx7xI9Or1VAtujZoiYYV8UCgftLJ7vioVC8inslgUon0
ADLm8tY9OAkZhP5akqpRsXb3GGoeEJI0Edvk9T08w5SCrA7qRJT6xmxMS891KHzy
yyegtGeIhtu2OnRm2yt9acDGnPGWBhPpbeVVTXOZH4q4+FOds6gK2erx6oEvN7C4
gWeK/tlDRRVnNdI9+vncxJewt02kLDgJeXdfvaARVg5xXEkHOZqWj+OYFD+imcDf
870kbFqUZ9dxK1u9UyqD7omz1WHpln6h/S6EGDSAhtep0Uil8EAJUaQYWo3qB8Hq
tYFZM9mVIpgTXAwsNNFBGIg7bsMrsEIZXX3Xp3vzCjYA4N7rTIjWBvrc3b5o3LT5
Rw+2UhgyYnA4kW+sZhiGr9vaoCgIaTbiriJy8e2QE6JPe5wxn4aABBL74rFwnjlP
ri6MRBY4wKe/YV2GBxOsH0pkzh67Q621UEoVDtvbV1Gn4t1/HMX9Zj6XMz2WTzAM
uNCbaHDXnIkdTOa+79HpG044X+FjQARAPQmMh3Lbts4bibD86joAc2yq6fS9SXFB
4IFRHTBb7tsWD8srDjrVxnZnVqAF8xuP/8LK8uixhwObIwnEMSv3Xf6f1WlNFpab
CHBiat3XuBVKvE3b5VoYNCiJa2rIx14sDZZv7MfrDRbVfHvHsbK1QKt4Jn9C7q9X
WXKIcxEKhQEEwb3FCA1dhugAnDXxbN30ozy3prpxueFKB9xXUWNjQKpvFiK8J9LR
kPFosdhAXDkQ/Rj97IG4yjN+USFEv0+ESPAzsCvOoedGjrfe4TGTRW5eEQpBxVtL
ynlYd4vDXBAtz5TmNdwFAJPQyiUMBbLTH6fDv9sE5JZ0UpYH1jAScuS6Yc3IY4Ti
5mrXV6Qn/LBMh03EbphYLcZ2YnIfXRoIC+tyFiKPdj+uTUVIW2ZXpFrb1edySPfi
+5qa9gigkC5Q/+2TVqDrzE91UH0EJm2nRKZNDSzltfMkKgjQvJdSd0DR38WkC80i
jjB+xcXshmEOVt2NOm+ua1KP7wUiBnPSLCaokasWfKB7ZNIUxJB1AAswf9Dl6l0M
4TgsNp82bbkML+gZ4ZD3QuwIGc8SDuNc4UkOQumYbeoGKuzhHHULocY4XFcpKkBk
l4SU2HCLUnmdhjHfAeGrJPvlPUgSSLeh+GXRUMbNCD2qKFalctjv2Q6R5VH7VBZL
KXnb1spVeKvEUHEdJGier4RnSWPCpuKaJMRhnELEfIYmrpcUwUTll6HBQiL1zDLw
krSouRnWdnoAscGOJqU/dDKAmJv5qXbyn9dhOvbLkilPkc7jmWVdWiqbo/wRfjvB
p5gEBpQVRxvgZ20qCMQKZNA6yltwUlkhBL/RvO/z/eQgqQUZz7KXQ07QRaSiK+TA
FIqlzf95QcFHgshrJ4Bq430ldYowasBEa49RZ++Oqvm2YgYccTsEx6ulTwAXAues
QK6J3UXEsaoUP3JGI9D41seU32B/adToDptEV5iet+EfbajW6V+bMq0cT2vvAQ3z
Z8Tp/Hs6CMCH0Ds7CqcSsiLk8hA0FLtq3ACeqqle1w8ns+7UiZy/vy6Xpv+x7wjh
hT4ao1XNSenGRGPS+tBC7VPoqp3Qp0AOqw+WbJg6UlxgTDVUNWciPe8Gq4IGzFoh
vhQfoVloN5fopiMXxJFCamSDQm1+le036ofdBfEmlDeAXu/F1mT2zQafwsuUA79U
9UWAdoTfqHtygf4dcb0vCJCcEVF8aHl+42WZZ/kJD39mVfexyNqSfing9MdUXAPg
8hOSo60AhJb6i5e0Zvyafd4aC/FvSVPkdwEnL/x0IMYEx9EgBdZs4fQf+NvLWAGi
gnJ1xhowciXZolwl03AObmvtgOEpQs8ilWe/dmLCWCkq9Pguqj2aJaj4GXNRveR0
gX7IrREB9hBZJhOfqUikD3Y35oere866pSS4Xn0+7t+KPGsbZx61SkMdHoxqhVCw
/EXUeMdha2eAzzZeFf+GSmLIDio6iah9oR7e23N0uLQrKZ/JxzFMQOQ7rc7Tv4nW
2MiXwMWeXorP4G8/J0GYSwVlJNfYwncjIFaaNRAonOoJMWPSJz0DKr7E6GC8oUFZ
FeT9g3ZhAD9unGOu8EYBuGXD8Se4tBoT3DdK6ZGgk7Rzk6hUXQXzLdOGtgUVzyJj
LYWoiVlyVJZJFaNwTJsugDX0Ajuudt+8Hrc2HFYbMc7J/Hfxzx1wF1c5QpvqLf72
bJgeEYUQMttt7p0/8Qhx+xhboDIvox45aIVS00zAe/Qoh9wcE3IkO75hAdhmvZGD
YAOblY/ONlrS8Bq3NTcx1faYYwJn7wQ+IfLej8RRT+KPKTsj9ijWwmrxqGz8yw7y
czHISIi/6ogMJed+GzECXpeXVzZ4d2LVc/4yYz44Ln7X+Y1sIbmDyj2zii0cjf58
t4cEspEzTeypSkHuZ5T20Ii3njqpKkf476T9pJsATgxhJyKPIalI2W0GTqdnjAIW
LO4X2w1HbXxmB2ZGKaHu6evAWYpgO7wDCEdMkWG2fqABA9r30Bk1194pHhL/pC6c
wueXJ0vb7GC9rnACJ4lSf7UJScnMmpViLJWL/LsD30lbdcQrt6RxWWUO67LvCTbN
gfFnwa4BYYA+33g2dcZ5h05mxHywU/3hEKTvm3XpRutf4zztlZRCk6f581CiwH75
lAsE2Sy80Hl/kR7YP5FRyC+orL4gzT0DRARJH+iJEUjYqI/ECW6gX+aZF4soak/S
j2A/DyC3L/vodcuO3lDfVaO0ek3JisDPTntprR25OUvpbZZX04pb+P3XOoD70usH
dMTH3oVbSzj/nz2WyDvjQOYGeqnuO+fty6Q52GjIKaVydjkKnppvw2LB0AVYhbc8
ctQf4sJUMATBHoBkh89izlcdjR7crDnTy99N8d1z03qL1rFVUe39jBaPaC+ThOza
lndfCtlSuEKi9+EBEJKLQwb5VP9LkBma8/8eMbphn3rDRJwAduyomDhYf9xebsj+
71rXDXyXHGwwQ31QCAIRAGIcU3uPPfQ6bjYmCaBPcnO1F9XItj8Yu1dW4/WW5MKB
SZNSAxjBQJbwNNfMHTGGd41kFobiy2Vk6bzF9Ize60TUTeMKaok3DCb2B9D1JKn1
zovoF5N4hQJBK/CqhBR9sWYfrJkbkU4Ekfm+rdFDQ2B/EDXb+nu9PinX7TWVGpVr
bL0dnOKu/yOfdJNg4Ddwh612bC5EVcLjJXd6BEL4yNnMVk34ZuokcQnIu4e9YaYa
871OSEgGRdQUtuiUPlruALA12Hpx4mFFm3+1pTosn7+myHIRZpOFZnocbN2a7PkI
d7HNShF/4PH0EUP4gmUgLd6u/wlyXYR2C7ZQWM558/wF0ZmIzZoX1iDI8FL6lDTW
lR1mriJ5aHQIkr5kD6v63AE2dQVaMgdeayGx83TxBCZ0REnHh8+KE7bEh7SMfDCw
8chFW17hwm6xHjGkfMsvCRceloymXOpq2WQzf/NMSkNTj+tXvCZIs7wUJa9hvHY4
+PPLCw8vK1Rd3lsoMnOKA/cEI84Y1kBXT1o7jksJCipOZ9jRnW1noBB1Vs7w/3Ot
Qo6hSE+ZvHpwv1fbeq0d0Phh6w4zzd4UTWa2MIxmNKNVYdH1mDpKAyn2b0+r5e3p
KtwQq+HVYeu8Z95tZdqgbCviDmZz+v35I4/MRxMajqP12uZFDmdMR6SL4PIgQ9Hb
thCuzyENngkiotqd8vzvoOQkGoF/+QToA5bR/9MtBuHtGG60KNCux7XetzrIVEiC
npUGuwEygeBVql9OCFb+wpmIOLZdFZmdfjz5tnjaH1yRzZ5HhXM9kFT6Nk2PA70D
fM8Igp1MYm8Ukk36yzxpPP41IGiUvP0ry2t1IOkkJY7Lq69Vkcyl69RAeNneYB81
JM+0lQABtv1eR99BBGuhfsJ3Rcb22aRg0+EeiqjxvxCkdyXZm1XjhR54EoxuPgC6
apS4QAvvVKbSalVaNm4089ZQxkvUcQKeTrhEANQOGd2AmVAbDlSr7nv2bPjoU/HZ
jmVR8Q9BJqCM5GoV7vfuv+hTn/qO+pkDTPIe/LHYbae5xQxhWV5vDchF/pd02BmK
cAIzdSs9tNbjRBA/x2wP7WqEvTJVSmLwGuvb8wesklFqsKrleifLZ9GTh5JwNQx6
VTSqtYTgTF3q6jt092fhCtii4XAzrQJcEFgZo6JdSmBLYetW9wy2atjIAfLORvjS
ECu1GxyVg8YmafBZQXY3A+146pXd/fi6UZm3BrN9/Z+dfzTKLVA8dNtI/Yh6x00y
MEo+erFKrFY0arDKQk8s1xqUDwZ4La37MqV/LxnbCx9oYBhzcYgHzWocf0smiuge
tnDZWKspLwIZIpLGvvtBaWi9B8j2696WiMEEerrHEJ7hj5jEfoD9unihZJYMWFE/
U7UN2GeTL2WN4XtIr6ipGxKAOeYre6h07jx9VCCoVDj0m0+O0WC/FhuSSfIjxUQo
mkJXfHJLUqbOhjGuFyrGmNaX9GvCijNOQH4mtNHmQ0NEd+LzlP9+iqvGBUHfScLO
DRN5YNsuzIbs3lpxqTHcD7lHJTJx0DXekJiR/SIlApa23gbML490xZbOqpo+ccoa
l+PhoU/laL6+JuiEhTyPplJgSG3i7zGEH4G60fBq8CLJ2eua2rDf3BjqhpmV3Xbb
s3ayX7Sy1FdCfbbW+JMv3fyuLWIaJMxXeQG4xdywizBwu7NpXrHh/DPLI0BbCGXO
kFM+z3N5y8yaKg7THiX5D5gdc8iwa70VW59nVMRZncUfGJ+YTwRYLIbJn4Kxb7m8
TtlSnz5JLnJXSjcZmjH93RCVvYc7OQsIpRMNbkWsao6PC6YFVR0B2kECPxO7GRAu
4SNjygz8k+Gcesbb6AsmUHOMm9URSf17vrVjxh6FDeBDdNNPMjdARkxQmhQWOwmZ
9qNdJt8UI7SsUZXUrd5WEE7nuuEUUBjvpviAOgHulR4BWZyqxs/PrMHwFwalFTgz
uQhFg5wpMIEZMYt5F0U8ifMO2RJzXmTMKcvuL4yTK66snOktRhISP9lSkI9szBEv
s08vrJEl+S6hzQawzZLFHs+fYMOoAjZ9QVsK4wUfnea0NPfBQhOEo5hC8NCf1nIa
gEoJ+EWUSsh2yNJvzn29lgtOYi5hTbPCRYdYkguxGJa/4ssFWcGJR3hm4zWAP/0H
W3Y3FjfbJQvv3998V5cMxDD9jxbNIl0ayuM/aytaTrztU+0zl/rkddpekZAqOrgy
MJoMRIhtMMLRxq3hTOjnl8Zk6n5mtK9ZXxpCmcV22gx1fxq5hElquVRlwpYNlg3O
wJ0C32M/BMVSLP0eO4xYECGGf0HngRSbglW7rtEtk6K8RBA/eHG0zkh43kxk1Vov
Sn7DTMkvxw1WFWe6r8PXSFn+aaP/GDwyw8Hhxyputi6XzcdDhjpUuRnAzOsxQyJv
lt4qrJ4hUvIaAwSB/sA9oeoTBiZQl8Yf0+WRgufpmP1AYiqfOUp9JjMsth/rI8BF
vyj4+hlrGbHfHkd3st5EyCY+H1+2c+1zq0SErnBAawbF4L1rCgkhZ9KyxulI9wBq
AnMC3hsPhRuCMn06yPjhoLW9oH8LkeTFqLNXhAER2ssz+2WqxB2EY5q8MX33ZWj1
nL5X3zcrhGHkrosozLda3mZ+A2w5MQXTQl/DwTOBiBTUOmkff2Ju4EsN5KVnrVRr
moiZrTP95i44KGb9MBwGH8ulz1eGtSqyEOpqxzGpXdN5aq7Ky/h/hYqLT61Mhodk
Q/B/rakiOQNGLvucQVKMlhZYPe9b2C0PMbBpzwMBMqHSHRnaGkXcG7PXxTSaoPZe
U8XfgvlIvqtRqi8D5wqVPF1SLvw5qVFwkxUrSqpaK8pKnUSVSpDeIRUvMc1lCZA2
Qu392N7530oP3TAxsh9nzOaV2jz/MfcB/SaARSeyQH4bcy01+KO5fw80MKD/MX4g
a7s7C+LT6Po44+q5RVBPcEZ2S1KyC0J/ZgJOfG0CYXEVHUPw5uap9W5xKdhEcoL+
tWyLGNiMw+cTdB6yjYwuW5zU1JMQBNmVNxTuNLkfVOTXBom4+2DHasTlJ82+zxsp
WjQtZFjIdOeKySSn5GceeliNfB/QyVF6GmT4dyAHsuyZvMKDqujfjGRd36xCzyOU
IaG1x6Tm9mXqy6+fQDEjmqParrz2Umplj9r3N00V6dL9ZodVSnfhwrSBqJ1LUTWD
h2tOqfzHHCmKGv1yEgwB+BJthX/+4U9gVpmh9T2EnYFwzMToxlVsxaeZVpBb9jGi
EPTOg+88bv/ewO9UAPhdaSOlb58zQKcDmBV4n6D7E1VYY2rvibZc/PuLIi8PpwSr
7oLlhXK0VGECF+kycA0XqC0k8566Y3b+znpD7MBGFjpK887xJaqmEkFAOMlyMsho
pjPwT7jFCcX9/diUK0Z4cuYdahTFlmODQdua/uNd34IOX2BGSQVb2pRNqGNrbnLD
Qn28BUOqBiY7agc2RvnVv/IwgquB6zoE2DlFvsyrsmYRfq3hoKljzYjdruN27j1z
ZaKuIueS8U/x3cxZgFT3PU8CzinTA3TY/emvL4Xuqz90UTdUMKad/HS2Nk4sJqCq
IHmgYmgbS9TRMU/fX8CJPh0D1ZZKU50O5CSqN0cQKhpC9INWXlMGvO8lUfM6DX5+
/tRIU6hqYb+Z8p9x6DG1gKSZG8LQ7AqYHvziw3AzeVpcIre0eSV4UzI68NyCHGsJ
tBGz6knymiqKQPa6n/mnAzWqpNpT5VDxXgAJ5ZF41qjDnFq5FBrinU8JJgJHKJRd
9yGPqx7IYBL80NQEy9Ph3trV4AvRWMY0xDMRCJct9Vr7Y07a8y3lKMc7IZuwluBD
mbwuLFEuNbVMdIGl5wnExc53cQkzsLYDVP1RiUcAtpa1wl8BibDbXJz5A2kLaC7P
W1e4Uw74vMOkwp94md3zWSaCeBU/oFAvRdMXbw5TiSXag+1hRbacmqfENosbfu2i
1i2jV4hiRxth5f+UUbFNyIhH9q2HxMWu7qHEC/k74703X19Icd81CQNXXT7Rvwk8
KA/adoMqGBiqtinVDxscSxpwCEdK91rwGbeCh/obFNMq6dyutsQMPr6loGMaiHQX
fbKvjWIsVWiYqfRxn0fmRJ9hx6meBqYYl8BeNAZRhn5dxEDbNTYc6TxKbXoeQGiy
CR6xgqlJr8idJjO4ZCADw8bzMXAZJ1F3VTKcStAAiP4zc5ph5ugGJTknMOSupDeL
sQ/eX2XK5uIa+GsYmBSvOFh0KA3o5I69cOBb3FRMFZEymgsvCkLJLPkg+FPfSK9e
+WQQtQoBar0ioCokVsuyrejlegY4pUwakvPpV1UpFOU0wyLCyb7euHiVH7SOVIH3
G7w3LH427psmAiXamOzmiFJmTv7Fw8JdSFjovD7h/fHxj5cjIjCQTQoarle4dmeO
2xDE6G2grVwygWakHwTrl6F55ZJ8imWF16ZwDjTas6RLiTQG8Zb4yq6TG5C0jdcY
wGMebWJMg8Czpy9Rq2UBw20i0yXUh+MDsr5pdvr/4Fx99awpCvpv1xY87ZnJ4dbo
vu/pP8OQ6sPyIWW0yh6alRqZxEMp+QuYtJZNwE4Yn4WrzZFXF6jXk13DHDvfCWho
mDGR8OgDiGoE7wFs/mm5gGrv2b/iyNzGn8JRWFlugZNhgOck6qmfnH3PLEyLRXGY
LDD5N3vLjjU8m1e3YUqFT9mlvRKf2oMpnrZJMiDR1wZkRPFucyNnq764yBef099s
K1Ihevm4rYUCFlPZqqgMb21hs8bShWdoF7zKW10BfIeFD0bYvhZtQsiLvfGboVxD
t2wNHBW8+MUQ4xBsygEMDirztebQXm8LfALzdKhtH3vS6urkuBI2yhB+HLn4sIzg
o3CLwagk7nHuBNhD3W0IUtjxa2bqF92mbfhA+0CetHu/FvfpV+jL2TzX8/ce8uOm
dSay6V9bbreMUN30o0FRkeu/rv8ZkBSBU7vbvHjJ0v9f9zlDalcFrclA5pu1uasg
4B03VOabarmDsMc9bTuMz6dXvfx93Cw5ZdEVUUcuDDRWjMJpRP5xCUaua8FJ5tv9
WK1o7ZRhQQ5sz7yWogPl2M3rRWOYwxZOhGR0vHV1JjXTQYn2n4/hLrk6hY9NL70x
5TVZrjL4Gi+sprmNyh//o2mDwroQz+Q2cocODxx7KFR9Y8Js/JP4P5Hv1vknhjUm
WpKZ4BIvbZcaxUaBTDp5a4TYLb1zABc0vPROFh0hRh21QEVgeFBLWziAl//auhm4
O/4VDekRizi5m5FFdBwTo0fBkEjHHNJXJ2/RlBUHzIYYvk08MDGaJCl5EsVJKUoz
4JwR4MHJm5h9xVfFJcB3YZGmX15dmMNi8Y0HYO4J3YJYcTkEtqD57yjNPn4EQqs+
EiNJyK4bfKWpicJIZ+/4R3t6vRybCJQfQCCdEvvBz9bp+TjxRsmeN7UeYH3Sw/a8
5cPc4ydauqO8aAfPtjHnC0xakaumc5/aDuCBCRVsz4w8wUMaVi0/kfdcBrGp1ofc
Kl7UkjHA2flVfCo1Ye1vdkypFJAeQt+shn1DRvBk2yZfo23jCJa7OpHtQxw/BCuI
Cs7g3NlEEPckpPNRgf3W3OTFGfqD7SZxNWjOorOGkjHMZZv10lEm4lBWZfPKgVKZ
/LrJeHqbR+BrOFUJq6sBdCeiD42rUiL7ppRQtOj7VzXjNUC9LshjKD0+MUYgDtTt
wHztqM63mTE1+G9jVlRL3/vtGd8QmpWq4dajFhF9jgAAWAHdb2dwc9qbsNAamGtB
5Sy2/mYkSUxyjb3Gatd3ZkaLOJ1ICdRQt37NDDuGo2dz8EXkgM/uTaS3cl5brObF
3h+QUqvi6cZdYUjDdCx75UQ03UESelds4q/hy/FtVZUWDqYyTfYnFfcVIRSq9rG9
Uik6WBrxfUhQbZ/qykiAW87tsRhZmWAyPObzMQVgVQhbNcOK5tjdfj6ulpPM6CyA
d8EWQsQfZosucoPPTvNF5eOS/bjBQJJatceycToOS8+G+s03iOXQkpmLKfeYhL7i
fqFsv+ON20ail/ZmZ4hVFF7CK1QLGD324zgQlHq/LHT6bN2SVagVi9KXgs4JS1Fy
Mu7m0TZSi5BbQklh8ZKXWhfJ4EvfoZ8xU8Q/faQC+xZyQSvupN9Dw/VxBbGP+ghP
WAhZ92fPs2336MycT3+HZtkYf7B94DWXQPuDz0yNmC0w5GkYbZC9PGHqqRsuB4H6
vXfEqv+nZFgb0p9p1VxJ6CnNP5M2LfWhthxFD1bxpZDp+vapfqH5/M1hfYWPQenx
/ircioZBVoCnvnnkLtDq6qTtcchhlFRCrVxgUXCkOk4vcnZiat8gmGpAeJcV49eX
Ycharp+wa21HlYlmfoRDRWn2pPz81/IC7+X+JyQak91KyTgNikKELPw7cV78AQED
3u4b6b2f6pwaIXpifNLgqUv+A3Ct0ENu0c8Z+FErS5Sh9B0tJ2j/W87mvT0k1FBB
WS17HNpzkpMPQWuOXPOsWZsNOeUPGLXgAJzfhkBBmk+XYTCs4mpjpcPt3Ywz79Bb
1GhWfFHrT6UUSPrEn2ZGBGipbK+iu0oTztb/8+J2uNnGtfQUMv+Lbn5uteztxKwl
b70jdqRvX+l0apP2rIS0ehPlmZNtf7rfEBYPdQpBWrSTSkmPyD9pfNUSojNqpHqt
JMwjeRm2Pqry5bOfeZf2XqprVCnOAernZHzBAgphJ/ZJtR5P5CtlqxgTj8lMqVcR
+pwPM8ErN9N3FqjllQk2vyhQpqfbt4Bo3MyPBKDSPc3zI3emkkyM/HVOSZNPhJrJ
HXCaIFjTU0CvvHuRZEkS98/h+cT8pmwOFT8rpSWkvFt4/HNWd7ovbm14hqMHE9Af
OBNW7Nsf8hqRCw+rlOoaEnh4nYf/7aLzcN25fCPqmhA+0UcIPa3euCEQxRmew1Go
68cKi0p5YKepLj7zX0KoHr1cnxNodl6rvOOw0nfNpRAqmX80BWPABdAFqRc1oZm1
5hzfYI350ljm9FP9VnuTodD+0H1YEvL9QQ8tNTHpjFBoaBzUZWDMYegwg8KxDjk+
1sVN7JsLrgR4MQtvtiDUou0PI/rFQY0oV/5iWRaNu2MLV4sBEwaNGERw1wp+aXAv
yMGdtP6rD6XIRLoFsI97naCrDsEU/sLnihgX2Gvx1XxERXXbQVhOZmjd8CwfA1Ii
wIM1eGCQ+iILbl1qW6qWdNfPo5Eku6aAt0+C8lGiA7dqB2ZcbFlJsLqB3ZdN+9iO
8E7cQCuym1LkUS4taQW/uduPzew/D3ekqtRX2kAujQTQPELaNpz4stiLF733+I2b
sBgXflV58ma4fv6s8NkWsMBCbIWjYpHkfmGbj9ZoP6dpC2z0ofST0Z2wU9OStWpJ
Pt9jG8Y4lgCMrBaCQV2c+qvg7Gk4ly+8UhDRH8oiV0NKof7YGd58v9M9OJwjBeTQ
j1hhWIPrttgqjyBezjSKW/MH5//u+1F7IaArWGNBbHyMA+krSJk1Rn9tGuJXelJi
CA879aWRCeF27xfcNo8Fr9z7Z0wDlQBXQUVEMHKuNBeidNpgoZxLt92CzW4MrGwj
RlEqYbQqEVMlceS/SiWMgzYNSl4IlVp29FiCUchoFN3qRw2/vGK6kria91HiD7k7
c3V7IDviUWsO3dJ9i/kwEjWz1NDtyHD9VaGhgnT5P9cWoWtuB8o0fpIF+Rs+NkT3
A0hrphssjF1OZwMHW8Wlv7nXCjP9SbTpPLWukyyWgcC4GoUy56nnMuMbFh0CQeEm
v+cFJX02ifKpMigf1sY0Ngo0odelaWhhKurmbL8kWR/n1HqCJS4d4RCVC8rV3t3m
IfNxnruGeW4R3TqRSq9xP77J+GSJHcOY0U60Iud22P2HmK/hKBLd8Y5IChk2IZkA
v5TVbQSotPGrM1yOXPd21rwBIUM48Y3FCAW74Q/l2i/3iPBYZgDtZ/jQlRC89CgD
4Vq8rT7QhEDCnVg5gq86jc6w7Rlu1heFB1GFAAmSX6TZq3EqxYq4UOiU0l5SIdXJ
WrP4o1lrPl7iQpQxrbUNTPaZf9ACbat8RciNHbMwtNorI8eTFvFvms9EQ+9mmDYZ
mHeP1d9slUoLEKuv5fFGGnpoqimPdjt1ApZHo0tJiHGEalzDhWjb8q1fn0+QEg9R
dmtXbmVRpdAWJka7/EQmh0VFnXd8HDW3/g6ozfrsjCMZtQdSFTlcHeUtSX4bNMiC
ga1W7sm0aJ6PYzIxD1XR1feY2maYnGdMmdcVZv68HHIVtr9kScf1eVh6HteXiCzI
f8gfyq5/I9D700xQST4zZ78P+xEChIDSlOzjvycNcSL1qX+Ijcf/xi9al9vn+AQw
n6SJjQV6HlZLgXCNKOwBcBPP7lQfNrchifRlZjdNZ5OQySAK9II0wF27may0oUGj
dEoEvDh3G5FKObAbeQWkWiZOavT5eZ+XpQVFLyHliM1slclPevu8yiVAwFccCng4
Qii2vI9Wp0U3/OVr/I3VMf4bAdDm2VcVSj6U2QrNHHsMJ0syqqomwxjKFiBBWUD9
5rN/0XKuUhre7lcB1fKjJjbnP5bAxT1y2lw8gqtO2kIdt9hXBKojV7zV/m8g7ccX
fLHvllH0KT+VEYer2nl6GMO78ynp+PtguePaAsv/TQdUk1RjnYrk537qkfkx7e2J
0ch4ZEdTNHWE23XkPMClFe+nvFQNtIEImiLl3C5fte/OIkAeQ/qIqgICJlpKUkWl
6FoqXLqJ6Lqib32hnSCH71o1oqmTN2Y8JwP4/QL4iTXDbzajS0wqb5wmSM2hToRn
aoeecazkza3Kcf3cCCzUK56ZosklDS5HHsGsgiZydRrfOCYFg+cD4nYWXPoNfa4a
+2X49c+FsvZ4C7oHtVr4RfrY9HWeHRujbJONzp4CJ+AL1Lm9DJaJ50493dAsVXlw
d4HoHwjKbDT34zC8NY6pwo+8E7st2TChrev2fNpFJTVm/MyTBZcHCeBm6SNFcR/R
DAwVjb8Lw83V3114l+jP/+RQqgNQPfpg500G6BuWkuRMI0AEKBTmf0qfRMTe52Ur
gVJDCOPZ3fwJZAYJRBXOMtJxsLTz0KjhF5szbuXW3GVazVmGsvIoSfSoibNODJHr
o1yPJH1HK1X3WpZU16jRL6dcmhytQy0XTZhY963/TqLdkkK43LUFYcd8QyZ0WRpA
8QApnxw8Sia9gCjbJcczstvbSjHTZhJW6rPZOE5fWRBMUAuPBbvNx+UVyniRWpYx
72e/6dTNHMa/y5iZtFd6E2SC1pdF03YeBm4OqFeq41fqLOA0sG6zwA6vzr5WA7J9
NiSRXoQuFH9z1Fc4CQdS/pFnQ1ViJizk6tX/D6eD6P7ipuNAS8adqgE4422mOt1i
NkspIA/W21VDq3K5NMBsv9mqvGhpdMmaOY2fm07faE2z6xLdKwDmhuaQQwlLXcqM
dPzXTwkK3wk58uBe/D+ck80IMRRsDHAFfG2jLw4YkMPDXEGXq0+wkzqsHMEswkf0
AE0FwQQMD5oJSon5zaQyNmUJ8V9hDpI9jOHuVibZw2fTfjtX9Sy9gFysPNf6AXaj
eWjY8vEIjVMlqDJWZuHmiTIYNyxTD55f9t45SM/a5ZUpOSeXb2F3JmlpuxeeH6th
Zdx6lu84DMp79mLmXZl1Wn44+o7jRQkH+HfYfvxo5DDMU+u4T4YzUv1U6Qv8oP0P
xCCtGh/vWE+0SkJlYnHGeoctyXj4QElIWf2HkJUY4ZYv55qiDC49doCbko+4hheu
W7/wXJvb0jH+fJhTpw6G+aZgxA3eMop8jHyIWg4RVJgWkJBSRCJByh0ncB8hiI/e
Ylti/pG2R2F4D7H1j8Ar2EhMTPsCT4dTZOVwlXmEliizUqxjmL2almJQcXNBivUL
/qvFN633iAP8TMDbeB246dC/V1IA6aZxYOZj9BQplL/Leqc+yHuhedVUQTMNV09I
dqr66bZsCe5I+6qUXMvgyGt6hkVNA9I+2Mv15raDSTD431w6Uncqu0fZI8SIV5no
1jYE2aPPhg7WeSrQkcx3AHApV9tOpzy1xScf/5DCezBLk4vm/BsNn8m2c6uxjKnX
wTHOeAj/Y+QB08NfCt6ZeFnKTGs7q7Hq53Gysg3L7G08kXMmgzwAjE04owxZdNjg
3CpUAadNTZueqXTJAj2XQimjnhtuvjnXXzsPexZ9XHRgXT/WJ3nQk1mRAiPEPTSZ
5OMxDgndLhCzfzn3ns6BlBvgxRYyMy4kQ59lAYONIB22A8IKCagj96Rc/OwgayFE
0wMDOATiWG5X2Hqnd1EIil9KqWdnHdZmvW2te4+Cuw7Yiacj8HPi3DMD//8hEStL
njkqSwAPXnG8Iwbf3ffmlsieWy05WpJSqw9iyEzsWiiWdMVdfmsyLWVNFVXxqx8p
pQpKdU3Dh6FIHzUSBv2xAa7PoGEcJOhrxk3MFA+SLo/gGl40Kr/yQn9UvPKQ51Jl
HqpeYziaVxbbvx8Y3MCoP3b27CN7ZLGxP4lQJtJeZ3tBCcamRlSWCEDgMAY+uO5E
cw4vNbrZDVtXP1ylf4qmhFCMWHq6KEyZFygBUx8cDZ9eNGgKD+Dm+FWAty7e3LKL
SNYSv4PDQm6+o2zlr6tmOjvCb4NqLS9i+Gg9kjis2kNDod8Aue8lf9TDnu9Q+UqU
a0ExocV+VLSen9B28o6CLoS2Ii7doNW7c6HSTKdn6aTArgks6Ocq3U5xzbYcNh/w
Nic0JgQWoNbQsXDkCVfcXIWjK5J6nD83yimIp+M4ea0hnKdSDicfpi3HkW6OSLl0
VtlY35VyUcdUMYgautXrk7F8pl4tf/X5eFfUyjn6DtM8TABnB2tn5vt7wz4nIw0+
MPKMAppsFTNShx7eft3smAAHL6nxbZodI1Qktm3psDKEI2a0kh+jXnKRIOQJ8n/j
wn5LP6IOHdkMB3JCEWCAoMQTO/ZFSs3Ovia2nG+GD8kTtNWiwYtJdjwdbr13aKbR
RU1+sO6pqU0kwV0P9JmYmvKIFEhkIVtMr1yTtGIr1nDMJhERiVjw0qwl0NRUTNdF
6IH5KFn8RBxNeX71v7SfZcvXDWuGL9ZWi42HSJ2cgMsPUR5YcX6KqwnTG6fSW/eC
90m6v4PAFqwxPFCFGZuJD0FGSp7OZAHjYrS2z1iKYlqJClLVEulcZmDQm5BEse5h
XPcLk/gps4dq2J98gV0s2doB6/vhoLBh8aMZZnPS9URIbSRFBuULASUA0kL9/SzZ
ojhhCnbcYFfJrmpzxrnSC+tCOB2oA7nL9dw0lMeyDxKXtWE2tUPp/kGP0qPsUTzI
bSDV3kmndUg6ELHxIgIagy1Q+Pp+dW68jbCQxc6ea5vkeg2vqgMLjfua+c7Anxnz
QOWavQ37aRvtKmnRulpzBeNPEiUf57Nu1Yb37RlFicxXbVOFoH/HEfyN+/PRCsZY
3AqztLr1UfC72g95gKutf/c6bB0BNS8PF/VhX+UfJ4HK0yc+EzgnAOKsm1ZQdlrn
CUNjyibKGFoo+eoXrzTk6Opfsk9l/6a1CWLOnGbSloQ1WOnHHiaSApkHbxh6Uhul
1s9MIrcwmSB0Whg/HbmAJHgZUf3QJnH2tnBDTuLVdYlAFChMkiem+NPL2HGQqAEF
NEmB7rJVqkBbMiLztwrzp7X3dJtBqA4GO+TIv/IzR/eKj65c0f5Wu426comLHDOa
DZ6Xtnx294NItfF1dY7Dvvf7gwN0QnGjfkxY187qCOYwIYBMIZsP7sCo1kn1E6Tl
13b4hlB/hId+T+g+GMOnHpkuoclB/T85WMiqYbw6s8ofd6u7i7WoXDl3F+L+1PdC
m2BX5h9N3iF0lYC4f1JuAeZmhHD3/IcvYXvB/itcTgf1K/hbY74iq5cJYL4FyWNj
lp6csdosEHYEb+bmRSctbWgWd1EtS3La4Qn62h5IUsxdV5bjZj72pCQ8lC9Kq/mb
f8+BfLlhABCYd2/oeb1v7kYcKBeUxihHQnC9Tko2+Q8T+e+MK+Ndu8UQpbzZj34Z
TRSy5Ic4py70Y/UeAHS1xbNd83VtNq3lzxk2oeYgxnfQWjzZvX8xz4qV60PgLqr/
0YhLRFxHd9vP9h7T6ihN2b1YrpYJrdPSYNfSY+RQcuOo1ORLU8vW3hSosa4Bp38T
ueW+tebVVK29ci/1M4lx/AED/o1BAISiB4JKWwdBK7pUdnJCyOfsug53DWw8sYz4
QLMnUcf5Koszf7hbrnpphpEzvrFTXBaeiI9y3OQiWyyLnxXb1Beb7G2xiriOb/aJ
OzcrUhbwATJgItn4k3gE2VJd2ehaeWxP7pKP8Ex4IZL9eVpcn+szhOknYWNf1lbz
MmhtcYDxpGxzU45d935f9dYKrZGr5CQ+xVbBAQiBd5eCIjIMlXQE5WRnxXm3hKi/
bTrOD2HaIljJvG3KJBkVPurwTt/ysJtDa0/+UjY3+Anxx1kvHR/mC7zyLVtG3azX
gsQ3RLySWDAPzXhcRbKm+VQOnHBK4Q4dK0Yo7vkp/yJYOLLIypG/S1ULjUy65nWQ
HoVrse2VID3tEhvGRVs4uuPLtZlJH3WJqF5NPcAZjJ/qNlmonJPzVdXO0ZSgREtf
Jdyqv84t5oHLsjhdpLKkir3zP6/epV+189VBXSC1G2EDlhEeL72uegTHvOozuL8+
E03vn95hfHLXmrBFPIWwnmX8BPeLA648DBZi/oN9zujnkc7AOjIYJV1t9TYJoxdy
ryIMCgXGnxXnayNLxxnuDt0/uOtFzZ3OcmQHtnQkcjPD9+WLPfPt6onrXv2fnaRy
i9NPFdonR6eexp/e7SUToq/+w7r7+5VOCrDv7pu7XB7oogC33Srt1K9EWMZx022D
CqvC9GMuA598YKXaekHvyy9NGNJnWzSExwMYQ/WkA5INmp0qIN3hg8Zk66wrqBIf
BN8ZuOaLGFMG3anC4eCiPI5E6mCnYGctSHjNCUu1BJTobNcfbskCObiEajUwvKRv
J069s2Y0+cUJN9iVQPFeoWqgtB77nKGZKaAvHinL++5q1XrFr7x/LYERoKqXQn77
bVYNl4H/8cLAnveS+Ja4uF2ReKgzCZRhAFhbLaDdt3VaNsauKJ2QC4X2YtpDyPAq
RoZyTVLpdJrqnKTUePWBZvW8fI14RL/eRGOxZMYdzSTkcPtClZYU283J5jJZnRLu
v3r0mgIlF3HB5pdhFZ4Q8W4LqDcSGS7wkUTItBIR/g9uhrk4PN94Vj+mFXGfyPJv
8QTL1t1o/LO76nkB9BGLBXGNKHh/Ha4O5PsEl7w/legEaJgmxVplZlwpm/E0wp4z
oWLWuF9+GMDGqVzov7RUIbFy2LB+NGL1s356hHOK2bRIOO9WLJB6CVVj6UyyC4eY
O5+h6k0jdE7SqzAEHkzB07SFkD2yNRSbi1XmYO2BvLMzHyQnFGF0sALOPpQn88TU
TzzZAPzt9W+IGSojYy5mnyExvUevPUA9sF+fpJEV/J/JeydkJdKOsaiPLtu35Owm
Ti0QsqChvBAOhKZvKuX8bdFu/qcD8oWOo6Jrs0Rtj3f8KZV1r8y0iXnomA0+Ipzi
eX4V+UnSBr4FI9uu/vHrTmGYyI7w88dtJrGm8zqDKLx2EiFxz0LgG2rZy6a8P1p9
ldiqnEtLMsIE1OjoH7qDXIXPDrU5R2yLeE3jbJ6tEtTfZ9nDZKA8S6sQCd8BMZza
qkhPUkE/2KBXBEVcj4kpGGIvHG2TPeVS/neEUX/KAcEnzRxKn4P6qmRmdG6MJk87
TDXYEgUfKHaXjVsIaUFA8V1rn1CFgZXG1yDggMCZsX+COUIp8Tu3QJvY+YVUkGiJ
hopJqygK7TvTSA3GtBv0dezfXq4um2X6MbW2rXZ8g8fBN+3TBKHBHkIYoc3Zctuo
arX4BwsaUgehK7zosdO0DXzIxfE4gAZ/+QBUH2EEYYBjgLRrVBjWOKuaJXdTtGSW
5TetpP8pkCsz/x9a0pM9GvKxS1jzrfhuuRV/jVJZxY8IhbZgMImcTlYsCeoHdqiO
iuV72t+9FoTM6eIHktwiWUKE02iM1kanLJ6kxX0Huiot36A8SFMwB2F3x/KUDH3A
tlgcXBfhDdG4UtmA7Xbg4H5OHLdgQ/U1zjuomvAM5/7pPJszW4eDFo2Kmql8AQRO
6mez/+Raj7uRt3rP8dWJBW1R9QQgU17Rkg6gq5Qqn7vQjTk/EwfsufFdTG7iC1Ok
TYgeIyIuClPx4L6iozT/LPGvfhVkM9eamZ7Vf6SqOyPo9pO+w7y2ksNgCr2amnA0
+j4HOMrK+ATDFB4sPha6u5md/cy6VrdHKX5Nfg/xZC6E+w4UV6hjwJcP+bQUnS6s
Anple8CKLaBzfVOHpBm9ZgW73P905KJYnljVEv7uzUCg+Gv6SHszJK3xYl7Pl5hv
PU3F54FIVViaPnTZTycmibdPfdAK1QLWzHfijbSqQ34/PLYqfYjugVM5D1xJhTJ0
d4V8z1x49ZaZ2XkfNOhtSjxkw51gbzaD4LYTo9qnxX4XHNJItYkn+5xYZkMJn0O0
qUKOeyPCh4pFvFxCer5sJMXjxoJjzMddGn5w29IkhMxghdj+E2YnZtZxE4k9bYub
3Rcz5hyeLEVFLrlOtgTRssP4M/I9vNfKY4BClh+tBkhM1MpvS5nQcGrqHv+i+/dC
Oq9ODIpV3AC89o/5hBJ7bazu1Xdw2ZkYv1q8l9iYKfXn57qoO+17nDwS/fOd7E/r
az8JIV+BwxGXAsR7xIVRCHLhqExCLa+nUiC6ZT7m7jc2r7IGPOm+uIregMofIYUo
5B635QamkkxjCFh/AidhXTxKbSKnqDMBIoCyCDBVMHWOonGuzHv6EHLDA+AKIJXS
LcCIS5tUgQyYzH7CFMNiKtXjCPOyEsjV/xA4/s+e8eX8DPgMjG9zuP8PqMRO4wA/
X+0HU8O7in8M7obZQS6sarJciBvjq5W5XyfekwIfFG/v+ykBv7ozCCDHtPxzjA8/
rP1QibLvsnYJuqXSIqlhAOILIcCZEkNkKvXs1SZmISXGayYnV8DrySWImICIQZhs
hNOKat+hguks0L+XlhtiuoIKgK3Xj2cCXUB42WpVEbrlTZ6LJNVNc0LIRv1qi5Jc
r0mMjVps33tKLf3rbkl/u24YGI2zMs7/PpZ9MPfWRiEWGV357n3MWm3Y+lS7+Zpa
q6Xlo3VfnmK7P7tfbZCe8vGmAufdnHz/9azh/iB7KfVZKUtokee0Jwpl3XgX7LxG
Z1geoI0w/M7akjwU13wkoL6eH1KlADwxxFL8R8fNKF4iw/sBdlSmUS/AZRm2swje
77VS1NodRGzd9E860Im9IvbUCRU5Ht2DPsJU50qxaLHxmDsm5beeOf0xBxtQ1rsz
XXqinqnf6PoN3gIykRoL2C5i0q2V5fIdaa2bV5yCXKnGGnyldApX9uBqNVETvG9+
7kJE5ZuCCaV5Xsp5uIlQFuhcZXssFmMFtxsjcMysUIYZnP0cHsZ/4De10F3Nn+w1
XO6fzeY+2Zht2PwXqMp7VLTOvZ0SbnN5+eYVwVfvperWqkNeQrKBR6RrL99VfzTh
aFCHsMJVxo3yJu/JB/30EFpskbjd5ajW2USEiGQO53FZIAeMuvYniF7otpoIUjw/
CxmMptbj6UcaMmtP/YGOocZ2d3787WHVTdEj6EpVPdMAwUYf8zcedxcS4o3CbTc8
/muC5x1Wc9pJB456l2L1O44jetOow4xRbrVLva3WaXVa+Nl24UHVPfVLzZLiixcW
g4IA7qvOGmGZTkY4cm+CQ1BEVRfT/sQn1yoj4AJhyFZ8qRHX+6f5ocLKumnLQ10g
h/qgZj0XLSpUm4WhrdVhFq6YI32brpeCfLYfEFKxxIZa4IIAfMpK24YWBJwsqx7y
OG5gNkZrTiLYy0xVo3kRGWmF4hCU2dqcqevWP8bPwe+TNSq+znJEDRQuinBrKY74
7qG9Z57kZYkVPELQGqyaFjrWmS8MpaRsg71k0RhKX/j1NMsbtsEv82tnc3LXTMZT
U7X/uYVKtZH0W493NBzJXdhyffMnwRdkMYRLBlQkHgTXZthJh7/HcWKhUJeXcfMa
X65YUsvVdLJ+fD7v1ciYJrQJzQil/ksJljZhbo5sQ20Ymx8AkMQqydhqy06i6SyH
/uU8xTmRqrOG7hgTmH6q9KP/a/aC9bxBp7wYpCLj9h/0wl1cV0sJYotJH9Ut7E2y
Q8GGNLpguSiKatKlPrQY9uEVVMRi0ExfRcwx6XSm3zI8Lkldj4/J+tAcw/cbsevo
Mcpdoe6VMSHEgvFC58nWV//k5tHmlZwSnDdWvDEh3g3qEPQVYDhPYMX1hykYkDgN
MTSVoYSbwA+jdz2yu06MJS9W14GhyJWqHE9/jQL7x5uic1WLXnh0yOzLmv1kF2fc
MZ9fw2FVSbECA/57UnR3FtgYaH6OSUqWeWEQj39ZfboNpxsY+X1n6rg/SNASm/a2
Z30n5mjr0Q5mN1Fv3nLvSn/SnfE9cDYfYktnGSzxjyX0hP6i7Py1xDmgAGk+T7wu
RDILQsWtq2SrQyhw+d1+3J9hlXoUTtkbtIIrKbrmlje4QgcRzYe1eGEkYVgJHE52
UGGN4Mzy8+3WmkTlE+5SUbtZbuTTN6gdhK3ii+psAxjsbV+YGsZe0bQJ5kOuKfpc
15e3OvBV2SeveA7/RPdg0VP6fnug8UVP/roEyWaO8GXRYcJcRHnJz1ZsqLSZIV99
9luA6PZL1GNs25mFNZ8OJRDJIVS16j4Cs8Hu04ilAwTZvfGqgANHWCV6msseB7e2
xBTPnv4EU+Zmr9r9GR0TJh8JK0O119LQvZ0J50PmSvGlaCuWssG2aaMUjf3Ddirx
kufW+NCI17f+wUDJl1Bw1vn0nGePxKorKcsk4nWZ28CSuvBWvWTJ3lcntK7ul2rz
u+dl0aiQxsd6xdCj/264oMxF1VYd0TPXoXOfrGvwtcUfQ7sJ+s/2uI2ROvvh3qwL
XzK4H3ZRSKHObbL9WIHXuxtn0CpwkTFubqCe/DjfjwS6rAi5u4aqr5fbBrLI3qLt
KxuNwJbNc1mFy4pCk6WAO91kinHUbwiwNp7Asq3D4ha9rjWjQLAaRTLiRl+s2Ere
liq9KjZPK4/oE+w9YAUMwLGKkgAyTHt/sp5JdHUcN2+Jh+5bsXJJE/pethVAWuza
Fe9CKtxh5HhLggzcUk9MfZucI5bRpP+VZGoGIF/jTf+2UG494Hr+vGaDNsBjcXZE
LQF3jHz3OV0a90lz32gUrqurM8WpYz2ZMRj1XMTu6KBvIQwyBDsfElHPQiWjlwIL
45tis6B9XCcfl39yHW5KI1Pl70lZoz+Y1Zk9/RD5q5T9jFL9PlndXWsMOhz2Sfy1
nZmlKFByEekaAeEAIww6278pI/FEDNQ+xZ8iIlL+g2uAWe7mCVuviFczn7lU22xj
Oku/ZjHqIhie3HouGZba/DNtoYoeZqX8ReZx/oaKyLLlpOhb7WYVD2Hife8ekqZT
cKFiqD93a1p/uEbyTTvQkrLqGgCIxBZBolAUUBmAK7TRHOTEI1eIl2Z3cIKbTsHm
T9CQMlTcm2PZUuTSJT6PrC461i+w5nzcXvJ0ABmijz2nzLKEaG98ExODbC389wIQ
OvKLgKAmmDWWkZcP0k7UvQDREZwlauiE4YAegbRaQePOD7EvZ8UZK1MqhtPseXFM
WGKZIeVPn2qLI20OK2/VpWTLJCLpvx2CtwwCsMfxTVXGx4H4p4RdHfN7v8r1gCPi
kBAdRV8SLH5pWygjcs6A7Kt61zRGrerjCPd2Ek3JeDLcvPys7CQyGJjGlyv38loo
EQpX1x/sTns0ivJDbVnixuoqJFVl9FjNWeuY1RX0/VecFo4pY6awFgt9vk0GAMYh
gsGADHY6IKjKQKRolD5C4Cfn1Gqb77892USjD1Us9gmWK8KMD7bOyG8ExMzAOG52
oD0Snf63sHee+z+5/Aqk1NcB3/oAG1z/Rt15H2HyxVuoaTER7KKVXvbiSfUQ2zjo
tEzH9Dk6rokymH0NW01MZp66f8AzjeVRfhocd5vmC+xbQP1PiGIQLqwYUV5QLQxs
w1mD2YzhlG9i3dMBwhmc7aDCLesoGRWheSCYFU639vdU/KMr1mBJWgxDMOftcoMu
I54PQO1UnT9D8YBC8rm8DTQU+8S03IN3Fotb4Rmrykz5IycALUzgHAy6NllEMwLa
7n+e43V07SEuxImMd1BxyRiMX+BLkWyn6RFvM4guW8idWXVtydVmTZvwsv08VYh6
nJMHSiopBAcVC7zmHkKTiJr4oQFOAEXxpPF69Oxvu5gBmCx8GInETe/Mq1B45D1U
HCplFyVTYNAZ7WDn/DPvn7NNv42q6cvxtW0Yj9i/S9D0kmYjEMJG31RlbUYahm2s
CjeA34gVE6joqT+dcvom/odTsB/Zltkx5QOSwYbJrGDb8IsIuxU2qt2sObvSuZ9e
tDw7s0yDghoIsXpsgRqClzp3YZX95Iaft8R1eNFBFTdICMXEbEYTPO4i1jXn5rm2
jl21KefoX9LwplYJCgY/HheoQN144dQv8cHdV1Bmu5OjJp8PHdOLeqWYW7zeTMaD
gx/U4DtbMVUcqqYnulRvtUeZBYhuhJHgx4pxdpIFRHEI7h4cwVS+lnTxSi2ORFnU
6VTTkqhOS9KaoAVt2m3H/UEgY0fNMAWGD8g86XMO1WmW2ZIxi/7FmPBuiBfRkGqX
LPscNraAELSAgbeMgJXvZQCtXgah1ZL3SCSqTDJ9rhPLefL40B+7gH34KJRd1BhZ
yKh1Orkr8lcd51DCKc2FHQuAU2W9aotXv1cq9J+ZErwcdnGyVn/aXWoW4KQAw3YB
mJpgW/gL5X7KiCgXDpWPkponnbowexI8QBI4f9t5Q8JCT+TyG6F70bkASl4jBSF5
JLKXmL7/yz3HYA0JMI0MNG81/W2wyUGnEfKW9UMB7buyVN77U2u4fCy03rEQoGPJ
gAGDOrNIVQswpyYacaXdMFJlmTNzHnBUkltwh85qYZKBsnMt47NFVCVu9CiSd15m
Ib0sTm4ytXiS+SWNH7SBCxZCh9zKgkV6fkIaYM6iqHHpu2q6IrICNEFyEFUiRxJU
ILMVes1fMcBha9uiz30MITeOjKJdAg5GK0o+tHdNzioRDiBy6cAK83dxeKYNyisp
y6MR+3V/qcd5HyXfM1K9G6Twf7yPE/6j1wyxxFQEpRKSimlUJTKNGdpCjUnXdTkA
/xvVW5Qi0h89TAZ2o1uMJl6vT5f2qY+vjPJAGP/w2Oz5f5jCwkAOPt1l2K4kAUkk
0x3GVkzwIpRT8EjXVTahNE/DnHTL/qceM+QYBVw8hs20Fl4/CUkHkJekzkZZd95s
6vx29Xdnt7lIrmifxOdQfsdrVn4Qlk2eKpPB+xKSnruRKINsOpfBhZ2cO56uk00H
HgrRD7XVnRYRNf32Gq7DwPPLOkZg2nhmD9VeEg8iqjg72wwZEA1l/zZm5kKhtB+6
bX4VZyOqk+0DphF3cHJg9owVvkhmkMRJ5Gg+fl2ksaWp5I+7e1aOk5KLIhayJ8Nq
2Eq5cSOMg5xFeEwwpQSJokZAnnLr1ukLVoJRHDIYQqMJpMLPeSIE7nQZbQZSe6JF
5FWnlcoN/fMqSEf3IwACI/lNUL9MtJ15Q1WdYlj6tmffGf/zKloNGbOyD+a1btqd
fZTMf/EGJNGFL1ThCFDygo7hXIBJMg/9EBhx+sLoHeneRVOak//fGGX/ucMjzYiA
fC9+KZ/WwsUow3hXBxLz0b9lZM6uimVPSZepPk0g8dexwY0LjP2uJVZ7MEREChyI
H/fdxoyc77WqLHn678SPMoHs5cMlcVMgEdSN/o8A/YiXnMTNoqLYO9FvqZoTlxNP
ZIRHyA2CYavyA+7ksFAiQO1qyK4fC+Aqi02y+JyYBI685jilr81oVUx6pDpioq5l
bkzbUILeP6Us37lAYbxft0TOtLymaZfEYDZgbsB6LJBzFRUdP2IAl0gRHP0rSbZF
3JZxLZrkhBNFTe5dyyqJdmfTJZaYM7KYthgT8J9hAfMhLr3dLEGql6m9Y2Oa+bAY
6W7zWClms1Z9HSxw7v2IJiq5EwL6w0ldK4FkE5RY0vZu+oZ97ZSHPaKfv/9jGs9K
W90t/TkIuJkGZb0MLyGNqF1CmT8sJoHLBH5fW7JeoeqrNfI8KklHSEdoZdyWZtOm
iiQ7mmoXPhdZOzpI5gF6sheMOIInTHvjJUvB4QH8htStUkMuzH2IrtLMYjbhC3fJ
HFIB651IpyiFEnFs+6vhMPGHgx/H9FD5k2zd5HqObw2tF5hmu3Kg7vR0Oow0QQMx
GrwevR3rxrhlO/JHeVXwZ1NS1abR/QKxDn6RAakO/Dv2Kr4cs5EUZm/9sDaGtiqH
Bv2K2LTViiNLqhKSUxC+t6ObIyuhQ4fF6pN6z+yaLZeoedVxrCfvm+UqEDzc5mcg
s3DLLkH6FR1dfqdR/+9r2mgN5lnIU0O1f5srN5W47dR01yBSRQwNnb8x8PtLXgTR
YG+H79q9DgqUiz6EmsYGpWkx6XKJS8Siuxw23qJg+DkMcmuDbWCMeEnM3ZQTCeMr
PC47ljTpOrlpVf95t3zxeStIKpBsVm0Yw6jgiKM8Gs1/oIk4nOR6PnH6Jtaradd3
SZpum0JTmPf+6Nq6EpXD+VfhYH6fEH4Z511zK/2FypIMfEDw2h/zAM47NrofG8Tf
Na80fsYBJEpWF7W7on/N/K7AtmpjdrC/2i9QJcmj4K6sanjzGwdQsyQXwhCGEmyd
/5UPJeYH49R55UqtY6NOTHGJ1Xqy2dY131e3po1dROmNm+SZ+E0fjHhabzd1gg+0
28c1+099ECbcTBbPEZd9Oeaxus1HTnoUahwLiurriP678MjVTwVZHDeNvC/+qeuw
/CAqRmlneTa4cYD9ra8ixbXVrMYJ9PdMw7kbLr3flEwef6YN1XVi/xRaFISxXxxW
hrevarzhYTSy9QICgwfLef2FYav0R2XNjgVt8qXZ5C5vMIjberdlwXrply/jaEiy
NxqnF8DFY+GfZX8Gj44dBEmnGkqlJLRiy1lWidu58Ux5BziN+TcQ18uhWvXW6AiB
0N39DKdzxxINh8vGObvWhl6MxsNnEoi099Xv5CQRo4kxORd7rphGpjpwrf59tXQ9
UE9oL6FcJvkpu0YcFBmtaJ2awmpKEpUh8agR+HJR2eYIxHMdQA0FgE124VwL+V9m
XXVl6vWOOaOrrrBVg2V87Y1iKk3ENe5/ej2k6JEt//bvjLPYHrGGLTAj1D65BhAy
k8JkMuXHKc9DvjEqRw8tH3fJ7ui2Z38D/ZV/wRcBrn2r+zJTedvuv39dvlTf3NkH
rnpbQIkVSr2iLRBy494RbgsIncHH38hk5KLFnFj2vNwlepiEVkdCmYo4hwxhuxGb
AgryHDbjqapa09vNlYbcFGj/4o6pjZRUVbqd18UWVLVvPvqYntK7wKZx/TFnc1g5
HirwFm/SrnMUrt+jSXr3wIFLaqueXs6n92jUwjLwvSU3f7v+7A0IVpiMmhd0T+ce
LsHMYRz6E/8+4lEO60XuDMUjvczvsCWQx6f+0HzXSroSJvtom4VIVfm28kI2WRiF
e15pAsB5zv7AeDpsTQDuwQ6adLmanwj2UuLLLBBeUaYlzYiPE8nuu8fz/qCkqbwg
mxYJGdcu+VOWWmRQT54S+4POocsCAR85fNmlHYdtHrIDaO6ysvP/icXJ1i4Z2QLA
2+lyuM+qoig5sAWvt9reCj6HyMXu2kzPoKS8ZSV+lIVsdvtgZTFKBoLko1c0qOdA
me02e4LW/dkS/v5+CTMLgqnfwisE8zHxusqCtFIQXOQGA5SOTvwF0WeroU5UBVX3
2XBef6+PrUYt3i8DilISFNG9ZiIiIOzu/wILiwEzBl3fqQtVWQAFpvkfE4M0uStX
1OgqsPCUG11Alm6SkAdZcktwXWVjBukgJg3bPtRsIQ2gGenfyuJUEjaCCUDr8FrJ
ZflzYIz+LJ0AsXIZWR0obQNTgkHcK1IMlKvZmAcOeYAeLRTZT4X/x9mOyMNPAMAG
d2xX+YtOoFe2htOo0nMozxuyWEnfEfi+ef3i5BfzTOvwMzEcP4Mv8q+Hn3JAO/oX
z9C9YXbKIaq1zhqsqWro/nLoEESrvDGx5IRIMeyCoylikQsGxTdVUJfOUC3vOUo5
8qQiaLjOzH4Q+V/HMuu89gWQWEehVEKgKDbPWiR1RqnybriKTzuJP+N+OYsqFDw9
/cDwKRjWv+TT6by+jLGGVpeFquaRogZPwP1Hhu4KsbCmnke909+ztvz72176fL3o
+/TVb6FfcCQHy4GuUHqBJyKFiBx7p89E8YSJiHCBFxVSy/Hq1qLiH9ITR5qLVx9X
miXKW4RycY7QZdvaImsLXI9+aBExLW5wqiSeRir2LHxjbwUiDCcbwdlsKMftPM3n
J7V6LaZVmTdu+egJtg43gWSk1xXGdSIFtEfK2pvBSX3l0zznyewzf2RhMjHS7kWV
12Ek76B4/TC27i+Srt9SIVVsGnyVZYObU8WoK97yW4HvZWTMivQKY1VcGNZZooTP
ITG9fXrPPhkNjPqKpGoO6lkBst0lIPFcFfa/h1qTrUyP0ICA94yo4Nk/hf7nxNzx
igvbY7ftcJJB8dcTuQeDMFJaQqk/vUlIgZPZ/kaWcCJsSTineioXL8K2tldJxU+1
wCD36IWiSQBQCgS7WUqCIX/6bRLrDtcdjGxGxTeS355AcSrIA4gClgDwcCe0JJWP
4LtKVJ3F+vtuSxLTM8CZ4kXNHnDru3uzUCxsDXLHgar1eXtOmUCK7Loj5A2EGBN1
mIh8ov6Rpq4gH5qFmmfYJht37qK0sEcn7N9aP3WZqtPCenotfYqz+oAwmOitKBO1
73B9aHqY1fDs9T576yjoP/d14ofk7wVhSKSHi5YSVKh7T+dzvS2yXbcoM/I2ndEE
3QNfx3nW+lZET6zT9cCUkjRF4ZBsSJ3MhjrY1VUGFXZqC4ea9i3KqDiiN3IrXjpF
Paaa5xO3yk9xcoGh1Z3hRilEnG40t7u5X4wuxUTV+AYLIq3CKSkZgYZppI16srf9
nM/fwnryROjgfpu9JnSH83Ur2wKAGKkjXhXx0KahtMLzkd89twiBSB9TjW+1Z6WU
Lb/xaU5UARnn8zsx66zefpZ4593wFw3/XoGwzevP5BpYjPEGrZss8AL5wB3q3WwN
rqfFpaXP/ru6ryoY1p7yLPEhuBLJsaxPzlUASCUjZA+XTO43nJBDnQ9BOFD+2i+h
QrPlObOJx9s6arBrrsEW3vuqxcdzPpteBKTaZh8x0c7g/7O6J6cgVIop8exnQBGI
w6zE6du6eLxtUT7gY+y8p+5r8k+a5mLgx1BLa2uTnQIk5zGnTOLQI58QwZOu7uwd
pLJWhfZj7Rv+e64eCLHPUP04h9OP1TcweJmeoQjKVzcbq26VFsqJRmAxRyLy0nRR
rIMjsQJ+qu6kNKAuvERqHpdWs8usQNVLhakfbeDAzigTX++0QnaBqm70mXTQQk+m
5SFyporCHy3KeoR4oNKPEO5wlvS65dRJTbjQkQwHnrHiiDeNEFRwAaC6pFjrLIKK
1/ozxIS3+1BaQn7IFrTuttmTBHrkDT+POO93LgdEz+Z8AEkVMMbRjrTR6EvwJRmk
iH7qCv2MaOUpmyYB2alU1s1KPqA51hKu3UKV5OoxLMxm9Tavu9TUX0BjsomPlTF6
UYIthm6LTuz3uHxFmI+cn/qk6uZrFkriTFjAY0q1Epz1rzB/MRMRLECckuSV3bEs
XZvkvEAiMljQTiSoefcPshtewbIu5kUcUQ7OqEeO4ynvKx0EYu/5BViXAWNIPR+Q
+TP3UGa+sniRsA2wMTong4Ud4bKD8wliuodglpqRUKv4XU4ZSU2fa+usnfSBIX3S
Bg44OUZ0GCHeIIur3bP3rny0OFb4VP+xPLoVUC31DOnyjV0Ytjj8gV0IYYBhYs8f
0VZz5E5ochWQvLgNIzgEt02a6A5Cp3nbfRBXVn65gLWaT10i5ZP+55Xfnu9fYIpr
mDFwP3T4jCNp3k7RW2OLERWHOSI0aq9vTUuXbxCNUSKXc6GLQS6UDLoyBCWDRc3v
U+vZZzJJh6M8SNw5/rLrpC3qdcbf78roLH0GimGIXt64+icqpur8tP/usopz2cho
z7hZHYGTmojFolqR/kJVhu2YEqpD6itAOOC4YAKiKZENoXUpzUdYR310xQYb5Qf2
v8CIgHwnwzFuQUf2JxGivUFEIcYmkYf2RFE1ZdkMPu2V2hX98iaKiyfhWHwgaedc
OwrRol+THNU/b2z0HVPu1+5p50puTWnHcjWrM9H8//h68FyKi9aLIWj8F2l/1xic
V0tkdYGsqaULOtmPAEzq/PmQ1ptIihrZplm4ChTZFEsnfT9pmKHP1+dZs/hqa+HR
vlOiRbLxYDaaHkKac4hKq7D4LANtapaDge8XP6TL4+Xbmj/2E8zZpG65AYMRPmYw
YrSUJEAwHQ0VrgHb5eydeDB2gE+rwtKRaCIJXWkmjjbL3KePthOIZWcDkATtkseV
qgi589Qmk9YsEMyaPBgTSafy9hgCTrcdk0tEfw9PkcQg4WkySJrE6v6rKxtdd0HW
gs+rAddO3mxXInypCqkOYO2E/gt1xesSU1gFMhevYHEu+lMjCBbz5Rsq+BQ890xc
RQx/IuEF5mTpznwLV1XJjoLaWEjYs/IBSU9NM3R1grIanoFfI2FsSFJccfDOude9
ArquEqv2BOTje8l8LcX0A55krXbcWPSmVJpeCWA8PWguqFByxQlNPvqFTHFMPY9z
uWZM77wm6vy4UIeNhSSnaEWeH+8fXIhd1wpL3oj+4+A2di4i7SeQPMyZsNMym9s5
CRK+U7qO1lEcAe+ldnHBW2/s9puLWGCSKw9HrXZlc+p9YrUk5XaUOBhOHNNs9CE3
7VYq6Kv9/hK3moD+lz0GK5TY/nkS3dpmlTNv6K4BGWEfwWbtXwI1e7WUT19Bzdch
8SZ0Ya8PC1l6W3CM8xH4K0w7RE0rK3TgiyZxGLpQGNYyBU6EBj4sDLIDzR2029t8
bZCV007i4mmZl9g8VAQN5b7R6mmruCvvu5DWH2IVWTDj+28jHEJ+ZHvVGdTF3ADi
XqvaWjpzRdM+iFV+jCLKx5QEBxpqB07wuOh2aMhilS/pB5v3LcmIo3ww0rqVwK6b
nq3zExBdmNEvrGI/E5LJ0IwA5qcCsj42b3CZyVeXCZOy0UHq/3jty+y+cSGMMlor
IZEf7AYrV5fK2JMLHBMg1OQrp9CsGEteARlsgc+zf9oiyPX5R7QiQ+9/JiXOVibq
WB1JqC/2u+exULQuH+zkPhGUq6c1PnfxXVt4PCpgUIBz5TviX/kfEzH0ckbWOTQ9
BHdulvCn6GYz0KMjcwMdTBX+GCMLi9q8uUyzyK4mvlYpy+IKDKhZ/CodFOjIkcBu
bqtDuxugw3lNz0VdEOsk9ZDYE1z9aw33qaPXBnsHgk7JOQML3y2MYJwlDCdgFgJ0
QpoHPy9/ndzzTRM3IkNz6jqvhYRXvwdv+imNbRiuUq9gQPXi/jgXxeamMr7uEHRv
FiYT6Z25ubZ7oAkXI13lOZKb86h8C6yOkaJz1gEc+HRP0I+OwwagDAqn92EIeb9a
uAAdQ+E9BsNTPF+e6Uu0yvY5MiDFzPa41fo4gTIXLc0VTC0wtjDanOGHUHcPmv0h
HjXkxdbQTO1gF9cPV/fNA9LM8Q7ejeJAtnudOWbm/lXLjb2RAPQ1gcaKIvjeZRQh
mlMnuiLMP9ZdDky//PIox1R9cECEUK4fydQodI+AuRUZjzM0lMpEi6dxUO/G60ys
MVymQHmxPKZzGlasLxHznf1AsBAPCLliO9AZHAiAJ6jXrXFoqguofgd38y4BEIhp
Hmfl4jRvlabVQ3KapTloYtS2bV82uJJYpxaNlg8oXjMwMwejrN2a6FtcooDGwGlF
iJEgWlfoPAMzfl0zfcLgf4VQ3D45tVYuyQv3u/0+XMR9CezezsbXHiyT3Ls9ikKY
vOGkSugYCUMgmEzuulRoddLBPZ6gJg7xZqGaWdURJCtrA+gv10HyyHpHzAjGnf2w
rfISH8XKSehiYzDUMYOb/oMJFBgh8xTPEuEuFLaZtkLknUVwaThYGFiAOyO6Xwhy
s+HS0Djcj6lNhB8kMQawzfi/RRo7n3zF336SntHlxL8xugD8aaYGyPBqwAkBVYLI
0MhgY51S/RzZB1GvTCvyutsJJdIH58+TBdWqlQEKZmgJjT+enDRA9F9iHmJ39mtS
GSXg9JAkXu6y02BRK5GgNyH32LGW6Jr4RAufIbgLoAa9tHJYARZ331c9rkubJYC6
U0gSsAVqnagqahUHqwrS8I0ZYQnUZ/kcam7xgu5x9YnVmui6DgL4EOilkVBDUAhl
tMe6ym4Z65nDgUAv+0HmCbjAgtIpMwk9JxIm12UmU7H0MNbmMOgq2/lt7KDsCaLh
rqt25LkI3zG+VRB+wHtY9TnmVO+hmBjqQoDXHztNIRw9p3qr2qrVXhNJ4NzKbSgi
RFPXqjN/5ZyauDJWPA28zcS75OPIEjdhazLtGgUnvKKkniNygXutwQX/KhWjic9x
fjshw35Tb+8kd44e0K8qf7Rz3FlqcYPTALi6/q4yhj1HVOZoQZfoju2bhvQQU859
GmcVHlfYlTbRSOiLYpF0AkAWKXl5aKsC3e553Vz3ILwHOLAebDSwm+tEjxI4K6gp
6cgjbZTuGgo1Jl/+aEzXZYkjG2azm8u3s8j8iRujXGMBync6fGr6daLVe2teGNzG
cxFgUGttf6O6Z0w+gTuSkFXefNL3qQHacnzN0usdpthffgN7OXsvvbfu/J9lgcBl
7dG5eJWOuJSEZune2ai5xb8DvMgNym/9PUoXXu+tJI7oSYsdIYmD2l0uemFCqmbi
nY4dQreY7CBDUHuA1saZAXTSR4xBslCZ6q0hPlyHN7K1FSweUmcAFmqIc+a2yEMd
yUu3ULSW1sKjllGCgHmD+q+S20+7PWjN1sf+gAIvMyI6POLDZ7HRV6mumNqQUXDI
mvlJKGOt6x/s4yuTJxwc1FxuvLbQVFefcZDtkdR/5uGHQYthjoX6xbsmx3OBZLCj
mMOZWEB1daRTyMJvWPh6woVkdkPCej96lNJkDAk6ovzQoKxkEkiaNweKIjq9MfRF
EBjKFVCv+FbQosLwFhiqSBBJISnzVPgMvlpiUnuJwkRaiKHp8FNo1dbZOw7rB/sW
as7mabiDFTZReyxGXnAhnUDq/0zm3ofXcCbLnEqT9M1g2f5re9juj7UtDyM4+pJw
gy1WMC2borReHdhIjbcU6a1SwxSB+UaIsBuvBBRNRanm+Lkpb7+iN0zHgAAGpY9n
ivQvNUwPsr5KczPrf8tqKCkMibFi4Mtk5e21ZrWPjJz2Zr6/Ck6Vl2/4E1U2q4j3
pNzR3rLdhnQgZjC3gRbLAft7XfHaDVW4WG8abtjgujfabq3oyj4azQXlZyLXnts1
yhg1rA9ZFTI8F9qI4qPQCRtPIoYD0k2sznfyuAhoP0XJG3tNf1RRimkYCX0qTO4n
om/qgvlSVT8Ijz5afkRcdE+wCcVTuo0G7QkOLqiU9jWMarr69Njsycat8SzKkWEV
m+zgSZeazSqr+dvtAUjM62anrTFdRVG+BzLhkdi0KM5LW4wiQJpUbp5Zkq7I0BJZ
XBpnZ/o39cbzX9yrHtQC8EcoF1Rwr5vU6VXMkLz8Qmr2N4JbDRPk9309aZ7MmAGm
sbTtvglYu98LyeJUmBrRSiGtJEfPR4ZZoJTHwiJTyesX1sVJBMSNTaiw6NGBFMz8
uCs9NJjARhhVAd3u3kciMVrRnIamo8xvkY66APSr+aN+f0zpz6hB170acnNhZsVC
+Z7TiwPAy/fPq2pBAgVb1hbdEyOJhpRF82qZ7NTfA+2kYngK5a9qOkTsiljLPMdW
hIb8o3lBS7/WWsSy5B7f9+MTnMf66ftJiQdxJPzQHMdQbiV0WLpcJD+AqPONo9Yz
2ZSJVg7dpgVpxfQRt0tq1AF2con7bNhg5ogsBpeNMmhbmS8flnGtUcSMm+g/xYgv
BlcyEg/DeOaJtDIyYyCWh9H+aZVpxJkDF7tWHfwTlEny5YVUkM4orhffcAuqatXY
1sPqbXOTMYVQF6RGHBGUI78/I3h/aL2SNKcAiG0Op5D97If26EC7ywrm4RoMe2r1
aAlhm8CfGf4VKY0S6sgdQHHjC9JmvQqjzMU7Qguboh8U5dCMHT8TSrBKlmfmw5nx
1lGsfHU7A3guIgWEIjQomyhdFXWH/jZ6vEA68W9/a0G1yY4yfPHsbxMbfHMyDOl2
AhDEkhkZaAqqxdhJw3tkUZIYj6RrESL6eEq9fwYPQd+oc0Du/Ei+XNCOWgzlfqME
VIfFrXI6PhEZUF0j2usiC2xlw6U3r1VF+a8Lm0T68elQBL4LUfySnLXqdX8P1mKM
y6h41Fs802jMDfa673TazOALiC1HpLGRUE2bD7mjB53enDLvzFhu0nfKwyWdmYSH
ZOQPMZIXecUnkaqYiE63RBwq8Z83KUZimExjf0uOk0rDQfcs5V5qufwtJeE/6m56
+5WjpwOwJnyyxwRPVsS0pgNfAs6CrBeg6IDCEEenQsMfNwpEf4/3f6P5tPjrXnUf
7rFoefi6qjX5w5mVGR/S+PxuBcJFr+gMrD9SFE2NlnOd7NrUvShBeYhct6R2HF0t
0ZjsW+vNhSH6FkAtinJu5QDEZsRGOFMg48n+T+QxJ6KmpZ7OKqDCkqbjX0M0pzNn
XNMRxi2cacR74ctMr8L25BMfrHPR5EjRlxqUlmCuKSxJpbainpHfjokscAy/B2Vk
L/3Y6wz1BQRXu205zxjFI66pz7/XHcpPmgXTMIsNMYsHnrGiyoqE3GeLTCablcb4
ZkWQKzsctPbGlZTE3LEMeonrpcmFU6J/xzEtucpvjQkkHERFPWO237KyIEIBEXsY
DbcAPR/nKbcM83+t174LRbx1VeYUEoZIesAQHyHYofjCO6nnIQlg+TKSXLwzNxNU
Dr1kNhTacRP4qbAnPQM2tYUkG0wRKtUxrlcCM8PbJE+aEx+fQeMz3ggw9y0uXs3h
cKoTe7MzZ0+ByGdfv5K5aXYNXDBkzkLHeEH1zt+BzA9T4yrMI4x9kzfTNdeZ6ekJ
SXIj6MtmWFvXGJwLk2efBcKjFJFSJaAQK2s+eWXvDqu9uBEW/fNsQC5QNhXhLcEZ
kFnHZWrMputci9b43fSuZIGrO2OHB4BzhXA1GCb+dmS7GN6a7Xd9iD0MFe9GYMiZ
xr9cQUmRCJQA7swkctwgt6oqlRgGuGNAcjUJn64yzZnUru6n4+SFKiHhvnXr9Ggr
HQUEEaq7knw5sOAwN9yqPJ+Egi7/ScaCKmXOdn2cG7jptE+zSRuQvZ1Mjk9w0DZt
YGTmBExMcfIXcS3qADXHpDBVf4Doo80BKHyD7K3u+HVQJfgGQ+Zb1iX3k5fxtR8d
RyUJH6YhIQxDySXR3KhR0073U8LS3V6FHZDXWAxv+OOlALihE5fSiR3UmCP2tHWS
YM/7YO6Yx7HpyDHkCYW33CfOzXvJKeVz5yMAitT4sX4avwTIs7W7g/sGHQUZ1xxG
r4gNkzR2HZnHWWa3saiN33Q0Ks3GRx8QYz5hqxtf4pQt8woVE0rgns0ZzLta6LBx
MeYj0wPm8pV+Bq+hH82TRFyaiXtm78892VaO25IQ8fVBsTmhlq7WzvCZV3jqSqht
6i5tGW9Ygt2jD5UyrbbUsDYCKLTQQ3tpO2mZNthG5i1zvepaATGuK8KI0Vi9xIPp
kpbkwkhkZKFx81igMo2K3yZ5yolLFAvdW3l5A4FtTrKvhFcm7q+yVB4WsrapE7Ft
liyeWEbiSNQ9lHV7SDDOb9ThYC6kecxgH0ukOIQ1Kc0apVHjNwcabjJECg501oI7
MD1mbH1+Sof/9Tjm2cjqfx0gR6xoLURBTO9+dhNGgE2r9TzxubFRzPbqmn2qqbAS
IfUwcl1tABBGed7XTHWorJsBopRQFtEsVS7DQ0VcEiOlGKIi1/OZue3oBY12X9+s
OF3sQFYrp+wNUcj6RqoNwa67UCRQwfBSTfnsT17MK/x5FwPNjyTJWx/fQkUB3Uw4
7iHiTiM6vE9lJOaJ3vr9V74Pekbk5VA4CC5+QAvdANqIAVD+jbbSf5zS+w9sksOl
mL8ByID4jnIIkFbOdq6IDTTaxDjRjlh75rqVXGTvj0ba0UcBC/1QqNI7+w8AteS3
x5bP6oRBS3bq+UQHLF5XM8ySVEOl5KNhUdJ3dOXwmB48F4aCnEyv5z8865o4TphF
/Nly/IUJpiyC4tvj0cb3QG5VUP1Rta5R4c5ZNoW1jRseGpXGDy/x5qWwB1hrBuUJ
eZf9gzSJmlQV3H4eI580QXYenaXMjE63TBIKnYdw4oLxnsj/k5sdz/b79GGf6pEp
puDQneDYhz1ulGx3d+mFjZmPHBFPrY4h99Ogcd7RGy1Imax7TZKX6If17CROYoD+
MuScqNav02n0SnMsmK6SGNDCmrkOason+4SxbtL2EakMhiMYGfEH8l3F2DjabijQ
OwrHAhMo3e6MK4YC6wWJIjzmurdiOEYihM5YVWXKWsYh+4iFUW0cW1o8p/zh04N1
xD7I3I99FuDZ08xdmy95Asm6wiI5tFb843lOpjZkelIA8D2vmGOmZ45muznoMKNv
CR2LhzXHSnFUR/X1aGP9CYlrXOv4zhiKbBBM+fcc3vyS5OcBQviWd2F1wtUB0Ow9
lw0HB5OjFYgEqAXLQds/5gMuHcl78vFF7cKPC/8/YSI4idsysZ6+kgDL6qL4Eys2
JxZjKFvHXYW7nbOaCtuhWh8fwfXbFEsV8EDQqaAQzW7dsSgUYqFoX35uBP4XRGiJ
h37CwwXGohSYxV2RSzyPSSNhrzlCUlNXVYnDWVLId7/4/SgSQSukJxWX8CEMfEnc
UGJqhOHRskLC0aA5QYMBmv+vSe3qPVcKFJrGDuz4WqdkrxUhnRMFEgMheBhe0aCO
i/2oJ6nNfu1thJoAna4ojR02bQ9F9o9n1QqLcmZ/i/LxjmS5jJoyovdu+KYSynbY
3e2dXD7505IIqsI/2/v8g3J7Vg2BLYN+91qMwFupvA+NjGxir/qfRG97SQ1gmiIW
i20t53PM+1X8W3G+Rt0TsLYmuzHPluwwWx7BTo45043ou7IE95oI1oeLO5QrkmXl
k/t5gb8Seh8dZHr7I51AAv2senU2mBvdc0IrcqixpI8BKv5KbUH4AqBYtKb8iBH0
0h9m5X4R1IIV30dMP61Y86sYl1SxwEtNjghOZslKy/zr1mo8PtY3oA6oB7CbstBD
VYBELVaaTQVvlAfzlB2FpY05F/El0JYyKIvr/DdIQKJwJS8OOAfGA+T12Rr3bw6w
mtrhK9KWZd8s1dKJfNmzOXL3sje3hG3TQDCJm4hSdxJNLVW9/Wgct0WB510uKK+F
0OS0fuL0zzUBAl0ujwWXXTbjmpoVDBdzGqGXal4JK1dQ0yEJO4g7fl9lYFzDR2wu
GEeSEMkA7p5KlwLijTddZG6d3jEDuXt2fjPJFvaWruxc4TIujiMo6ri1/58OsjbW
iJ7OCl18EsLAsmAQmOGMP3fOegGfLJG7IpPCSUo0Hte4tdAYq02Z8e2FGgdNkeI4
WmDlUIBPtHw6wiqpmaQwxVM+JYb24I6wsWC8QVE6HB63R4u3VGll9IfhQU20429l
LzBhulrww8tSqch3RP9LxsU5FIUFUHxp7G6QXZG0Vke7IPl6HbCUbqCW6RxuTmDS
nBYh5/u6npbSk1HHCjsdr0SsehDJRhyA0IE4gdpq17/ii4S6GMy0j/OWnOVfWvia
I2KXdjRBQkdE6stLjo5cZZPPvOAk5QfVZ0bWhUavnjADpw8F6UjUxakM4HEE5leU
5mTei8hgocIL6NDEyGvmCBY12hzzfytzeBbf0iXWdMStKHYsIsIyTzu2JL1tvQbF
PNfrXN0LrOmfbF7jVNaarSNoGFIdicETrbf7E50TrP335k4gEm21+l75ye68zTp7
q0jQ1+nTEXt9RaPpnH5SfkOfJplf9YrIAESNdp7NzY/r/n8e5ANE971prWa9pnS9
IFF+0GfnzsYhdPgBxTFork3mlyf+G4NGiWp+4fN5bHBC/4Tql4bBTRKMLPd3I6zB
zl0UBCHLyAV9vu5V3Ns1BnFP3L+FBlC9LURgKcp3xEpuX5n5Kr992fMt7DbGTg4Q
Brh31PoDqKUPL8E9rZBnBkJbGhyvdcbz0vlr3Mh5G1hzoV5Rb1dVXmVxQuJqKUKw
N6xg7tO41DQzFpwCpiXhBKgOfyDkQ0DeJBiFaKScCpREjOYTcQhzp+MqTCZtyCfN
IgBwjJ5hPDll5iYXEWu5RNfTbf7Jgxv0qzP714d8IlpZxE2Kuze0q+YH1I+tGfhK
mk+zykEopA91VAgnXyhDqPZDQvRPu0wqrctiCXwibR04ifSDl3/L0Y+AhXj7ZV/T
As9yzFxH0FaQnElIaidaDJk8pkKWiCbY1aDJr+JQQiXmBdjT4OW7+30GdvVCB0pm
eWrd8roPXnB0Z/F+ChZNo9pH3TEveK5CP5EUWnDUC/BPufIRUfsXfvNdZEB+5m2H
cpoBl5WbDtTTkYA6QDFRMPregSGlTm6+aci99fvdIUHfO1IkNfQkaN6M38NTp0x8
w5pM4JVr5O9lmmRc/iysJ/9qJN+Z7eOWx8eBv2yA6aArFnTZgIMeLK9DmE1IRkzm
HLKFXqXbkAxYvD/7yRWwZxw2g0WoX2qMDEziVEuIXK9ouGVoTD7md82rl+5mPhOt
OMTDaldyleNJYAwq6LO3V+hR0dRAj4X2gM3MHqzzZVJSxOj8msaSUsK7dfg/YxOj
A28YwEUFGRRXlzueBvXkxbFIY2pGbUBo89iH7/aT54X+YxY8UyCeX3WkoziDHxXX
7PpK3Bd6M0LXW3YxrSGGdkxOkUzLPdN5rZbnrJznt8z9UglJW/Jf4O1am50GoCER
EvHpA6hJ/jLMN4bjc2edlUD3KtTpvIYrwc1GPJFEE89KZ+CdFrj8ErAFvtVvUrvs
YebajJUudnZdch537vS8Kv39tADKRJbSN1mF0N8Gq7cY2jBh9lTMpzQDxhaUsA7m
8z9+Ytz6UY2KUaO6IdjPzjHo6UPZSpZE+H8QW/U9F8jQZ/KTUa68nq7J/6WwmFE8
0qYEgkbFNQ69jscyRTMfdGJrpWGo5SfbkgoZlDg0PXkorhRbu9PQu0iCJfbzxva5
2OCJnEyTvkbjA56LvTXqKr3glvDo2+9foV2cWuyZFBQlqC+7ZyNopfZogQb6J8pX
VPOnxOXIQ6JAblyoPo2yI5aCP4jaS0rxi0e9ulBAgzYGJej9q8cT1LPGuIVV//pI
7N59RrajpC9hg2Okd4LbpKnWar7hMFZPCIrEyGT7jKE7OfjzEVHoGNhq0dawMOcX
SBVF5nfiSfnw0paGxuVIiPqJbbD3kdWY3I/bLMqS7yKqS2GsuN6yUUCHCQLJpyfs
5z9DdtRe1YFcqRs3iBjl3MLlMDWFj32gjAZWvGEfCu0=
//pragma protect end_data_block
//pragma protect digest_block
W5JOgHSnHwPgdtKhrujswFeJIsI=
//pragma protect end_digest_block
//pragma protect end_protected
