// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KMeM00vCZcTdcelMnsgH+inLX8RiUNPZhjkvVr4UeXG889lA70XXV0uaOQ22+zw2JsSfmzhuIjRI
A/2P+a2pEvhCyy2lfwD5AJMA8y56LM2pbJwuUi+c5/1gGB39ukqNQKyTQeqY3WXHloeQHGqO6l1w
XlkSbr6Ji7HtgVTlBUryX+Hym6Yj7Efn1xOKGQtjoIuBUo1PvSi1bGTyQDJTWglIqzKLVQbrR98X
NQdpbdhj9lgTjSfgzUFwXUtGbqy9s1j/mHMM5wNWsbTwYRSjV6kLKyCc2eKXTLdWF/MW2JZzWntK
7qw9loIGqvVUAMN+cdgW6eLKY0NmdgppvSOIyg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
OtXgAKD21PWCazuc7yK3gkwxBgjRGjx2Eiks811K1gq3T6jPmCl0XDs5KZQaLRLSopdLvFcIU0tE
PSuOD7FgiZPgN3FtOhJ9Qr+yXr9JUcCemwnLmBC4SmAPiqmt1JpBVtokkzRpfmxf2/11uQT1rZdU
rc+o/YqrXABUe+A3/ZBNXfR8KbpQhHYDEi0775Q6tnwY1A/cLt2eUH6y1sN4H/k8H7IDF25sk2eN
xeKFWmuYycP7pr6T8sStUQ3CQ/AGv9vysNAyhkBz0Y5HbjQdwVxvYQy5uoPPfdBYziSwXZjBLF+4
YSOipGyhlyb37pZ2U83uSSUwk0RuoNQoctGaM40dEMGA+9CQ7vhZSHPR/Vuu6Q4PKM4eB+ihw99a
VPNHhOaK4LVxrIo5R9JHNn7gEw410kACfl32vNyYUb8avjM90MZuf/+miZXHoZGyLfgBHCexCJ2W
AIL09ZQkI+sMgB1fGexql7yUyJwyIpmKyk1OXe5eDURYMNRPbTXnbnCQ2cYg1yJBIsJ931g4juFt
Ep1yBwCu6ArImW7wx/tV4KcAoEHtQtNQHOhfFBkgrV9duqeZkxK8Slz73BZ/WQwrYGvPY5dncATY
DOV6MKf5D0GP3SoC5Z4upLnm9tnsZRR4mAAj1JDIrvIOZ6RrN/HAmGI0Z1IlG2a3mt4++56q7mFC
R1CjrrvTiQtvrW8kKuShoUWHReeaGQ4mE5zjRPIzRsK9ABJGkZy6eQgB8qaAq5QbkmIb+dEehblY
JRIUF51unVeJxWHrzk5NJ+fMtT1EjxH6Tt/0Kr417WKZm4ABhgHXtabShgqRLQf4eoJbr9RkNNZz
EuQX38D9YexDniQG7vIX3oXd1WHG21J5KMq+G4umdI6/vZi1PrCNq5HPuJVLJ51COA2vnnWC/Io1
iAnc8sVJJDDcgVtBGV58PIcGR1CIKaCwAuxjdyvO+MT1+pCsxW9ylgZesoH1Yqg+nSIPsErNqSpQ
ZCPqLXslnfo04DzL4Eze7Y1sTLg0UX5KYCcwF5RCVCZAQkQX30E5dNMXnY7rGU90S3ISg9aEj2uh
8+M5HhuOAqDwtMZJ/b2pbwNuvEkSozh+B3L0LpJ+7HPmXK8JpYY+SxG9c4juWW11TZZE7k5Fq0WA
FEhK4L+CE+1+lg+GkAY1uqp4y0gv5L6YanKpsYesd8u1q14G6yTmlq+YPwtQlDmb0OECvUIqPa6S
4kO51E0s9yfsDB/wKmBMNvX1MtTBYFdbMutt+a9ffDA22+rM6SjqeXmI6FROq7TcJv/Sg9tvdYHA
rXjp84uHkxGHz+BdOeFUISpcsqmdXaB4UQSu6/PTHujETL+60VdZzSPq66JeC7tC/xWudeWaENf/
EqXqa+Cw7RSSl+YFpqJhMnY2wV7/uRhoFO1Moe42eNuhpe4yESAAomhTzOqLP2snR/fpHVpQuMuR
Xv9huJEVkZcK4XyYjuxtKwNZ0gZnnJUWFANhWz2cfBSZqahJ54PHoT/wwEbt2BG2QRTVFvCBc5u4
Hp3u7FU+EAIp33Ob80LCBB2euOE9qPH3EVuhFYQITHMy//HIRHiKHfFi9ttosUtNRvWeSuqpPldj
Iqpl9LABQmqyXU5zihKUg0JUWcREZYy/p3lhHfgUCVTMAQSotQSMyp+kU5fu8wSMfhO8eMVIu6HS
CEtllBLfFWwfMZ0j5hDyGQPHEEHEIglTOxOQ6rUKteidZj/pAHoLj4HnXhGbLBor+kFlIeRr+WfQ
pSSNGCs8ZVIuEjaZz4cVzlUyv3SHrcH/YErt58GW1l36KB0r+ZBCiLrJ7JNFtlXJiYevIMH+N/Sn
pLiCVxKqQDeELOCzOE+jDvDL1SalUhdBrCsrvmkQqDIOMhPbE3MtFJyKIV2+l93O/rcStDDeKlal
BYl4cj2g7S9hrUMnZlT5imsw42TJ7dKB674JvfRikbVXG6rgRr8myt2L5JaNUK+PsDuZpz62wX56
IlPRFFG31DBRIZeyTvdJqiUnH2TtmenRfCjElbRvb9IIYaS8Re2MXcXTqFsXegcONchU2085Zzlc
Tw4oTqB84P5l2rM2sOstRpZen3GY9bUeZw/TZSMnBTOslOUNx5PQ7U0TdNJX/RSGk9paMNkotHEY
6oAkm8+tbjVbf1/z4AzV5v/lusKtBx4DlZlit9v1kfxp9HnABBccvKLiq4GFe1ruf7CXuSW3ojoU
iPO5mnGcoK8VLhxg21QF+NXysc4VlDiz/a/5ElkmJukdGi0FEQX/40o02HPX2tAVOnOv9XBQg6zm
xLPn/4iTry4tCqmhgTslpLY69NA5K19kxqTPBw0nmT+GcAgTlW1glrwlQizRIhCObBz2SQdtmQo9
EPdAP0jJb5fccwa6tfYo+wjoDC9vlxKrctRyhJW/Tu5eAu5VIpZp+xHehwPK0b9HIa7STB9tdFxz
wluea12rO2ideRjyBO16oh8wBc3H5Mf4k1QDcgiRhEAkKlPv2v5f+6c69OenBuP9EXeNy7cVkkIN
UCbs8GbC9igPX6pUIBZ3cTOldB+f7/rlKsYIL9jBvaogx6VfQhAopPfFuUfKz74MOTnHj0nmMpFm
JXDcbVrj+xYiKxH+HXs+K09yJBcNKZXvRGU5TTWxsiNlx11ENbhfK+bcqFdhp6KB2Om+ABcWLVs/
2CE4urs0Q0rzd2MEAAt4PhTRZdWOo4I+XejmoawwHXUGPgS9cAzNKv/yz70WbQe+z6uvqbV3d9tu
ViakXddMfKrtJfXSOqpZR0dxReKSO346/JL35lqVaw5m8dLSnQKRaTM8m2F5VncJzWX7X1MBjgTw
frRVUjkYuChfEA2curxlF/hKOtXmIXwrOr8Xey0SrifEVg3dggEMCzR58F5+9DN9+WfbfYi7EwTV
yX2FQLho3S6jgX562TBo8nrL+FeLPlLduhauIE8fD8cApPVYidB9iYOvptG5FF3hbHtH7XuX1qaB
nnkiU1zQ6ksX8ad4Teqlzl9n/49b0Q4SZQxgKMO0sVE8y8L8vMceBaL2dRzu75zL+lDFdrh5DVSs
Jd2tGVjvHOsYZVzFGLoqrDvqgH4zqOr/bb53N1jshjYoPhtvNlDbWB8T36ipNHB7h8GoawKza5nB
O6LTlXvhYDnjktkXYBw8W2t04q7n6VlgpxwD4uXMkMqVY60HKsMLRikJ90CjbULVq4KlrpSlit/t
CzfbcxHddM+w8N5HzAKJ71U6E0MjVUOg0tovv/ScBzEoF7dGnu6rIxp9nUsViQWOiBgNuJGBbaUO
Y58hJhTZx6xHVlbnNvonQwFpRi6RRB4heNfeLShoZQVladSczCTem/ysvPxZ12bJ/cdwwPGhLNny
0dce1PuukUbVzjIvw8kv9Xqg3agw2+hIFXUGlNrJVBoe1kHSLLwc7zeXajeD5sP4ug7kGc9Dr78H
E0uqVI66yxa7d4cROeTZ6HICY9sZCxcXvjTflvi5URYlVJCHGo5+3gCUhWtk46sGI1ZbRc+kiZ8q
VF3Oq3NFIuL8EDPg6awuLFx8pjPmYn3RUKtmWfkQgP67P/N782AjG9xFmHq5kD9BEsbzvrAdCTjX
RDNUOuyLHMmGXIXm9eYxyNoSyXVTejbw8hKOzxgjq7BGJIqPtG/6kgZFIRvXYAM4aTwRr+ZQ0Sfq
DBFL9pwvFCfdWU+2vjH3kvOkT9Is0vIiVkOP2A0WitBM1Ri7Sp5nCgQ+2Ra4ZngQj25L6JYGI8AL
nlAceUw7nUv2O0G0IJe5LyKlGID1JADhwTxcHphVJfD1ihxe61TpCQb71IXSTtfLMRVV0UsfQe1I
1sCPGkatU6hg4lr42ZKboC8NWkg/Z2NUVwGdQ+IDbgAtx4Jjrkw1KA5QKtoqKoHRGW/vQrvRBvMh
vE8xjwQ/9yGh2hq2r0o6NgUAzhr/DTN7AF9r6rX+t6Tuyh9g/q+oEKXowC/V4hd/M1HbE/QO2F/T
NzAXgB6cqnFQzqiJ+4h2v0DEfQkVr1HydxY0fbH4Qp/2JNVCNwQG3iOLo3q1lR1IBL+wusEvahQl
j16V1D/uQZTOgod+/iDoAV5dSWOAPwC0SLWk2U2ZeJnZWVygisbTBZ1EPhmTelLAtZB42tZvjVN0
3zRdE53hxNLAe5Ah015V9sdxUCSxu182x6w/fIMrS7nvhTTp/835HfwYBIbJI0Zs6YObOI5mUlix
KeUD0CpvlyBopjRuVd5wcVuY4K/pt3IXhIrmpPnhTxoS0GlgeIrkIlUBrixCXW4RvqPShQYQ2Q80
Ioyk1zzZ++R/ucgfwqcNoc8CHmz8NKBm4DfF8oHgbbt8fwF5A7t7ulyzwIGAYjOvx4q9pGOtnR63
KcR3ACT9idMRQLz0WAdWwCBcuk5QuIoVqTsEFTbzLUsGN9L/0HXAdvHRAf1ASKzmZEiphlyWYHks
qzmdYB+DE9+SyzS+L861JuYGvOELxFKUMrXb97MTUj1caAU54NLNd9WTuGlo42DPeE+7lsF+lXbO
bkzK6+buTgb0dBZyqWmu6L50JK6+cxkC9QIfHLhaMkaBWjEfNFQNTWEh9A4XvPm2pscR0aDR8VSD
RS75OI4eNdUogbs5FCcuAxBAfhpsPsgKlngoeV+jUAyz6BsCvBlb5Srru2/B4ujFvcCrh3eU9nUN
DQj5fJEhLqTX1rqwBsZ43Z1yifd0sfh15TG718yabt5obNOgSIKs/DZQPEf63ZlU5AISxvD4+WwN
HO/rb3ZYey+mJFanS0xctXKXRn871COPyr8lun0+ftZGB+llxdI2hQEPogoRAubYU0oQ/hg8WDy4
EmBkudG7cjKR68YC8iZv5zUHGx/ybYiYHFqFbIbia2wzf/CrdpAEoX+62PY3glInLIhglxFmR/Fv
m6tK2scPPPHNpmZKv+2njWmBFIftTCd6+GZHmBN+nuUD2YdmxqoFdACY5RR8zh3LPzdBNLmy78s3
BnxI6wtqtRq4KDCGnZSaNnywLRMAxWQcdB3TO4MllFKP2B+G4dO/JcxFq1vAGNdGJdAvn1c6OYOE
g1mmxg6zWS3Z2RWabqqmHeE+3QEvM5FCuvRFcsA46Z25XMl/iPM4dCvwR62BQmwf7HDdWecB5pR6
qU23aRuJxXpbY0Aeeu1aHcc2/RYxIobFhez0a9ZlbjUIpYPKBAMds1e5+fcIxMnoZkZ/6Z3uDYtI
+vm6IfGzfZ3qm0J1oSAB1OS993e947aOL6XuVzwtoIwfZ/cCcA38Agd0gW8Bf+blMuouUe1CcT7n
HsXU/rfTdxFVm9FRd+64GWF2m4b7VluFVSybopyJvxJ7paCyUMbZxrc2TKciLfKqGkql/TdEH6Xi
l+wa29e4SJ9RMVvhYV4sTHEVYC+VK5H5t0+x6yIE3hxG7DcvswH0KSErwQiUt0BWIbBG7MV6Pt+J
jZd5EtOUtMlDScjSKCgvcr7o0opiZE4pUinzbH/5EUVHnusruTkCWC2M7p2Pug37RqcEcntTAeSl
1fN0WkDBQPWwGFCo08Ie4i1d+4T4Ne4P8XbW0cTkcbpFXxG2+g9hG4chYC7Hnb7ybYy7IyyIA6G4
O/v1quQ1ojrECkjCYZ0GPo/Cpri/dM9R1XAII4QRsGqz2dftX1ymFr5Fs5FhzeppcsSkUu4Z0g+R
psbwvvNRGYzROybiYVEydLXI6BH90DtUNh1WjNIHYNPsoWUb5hl0tgnFVKZEXN8rhSMXx90+g2G3
nqz7EdYIFZhoprm1DsGbqK4o72GqAJf8hCCkBfm+UIhFpC8K8mPkVqSOPoheq+FrdUwIlfesnkxk
/HxofHI42myULJXvD11/ITVttRJiCGh77UE/5n1vHYTkp6V4WpwLcUa79mloVoWmcZDML4MmYbQP
geVtuenHn2ThA+naWFYviE/AswaMhEc1A+WcaGvSi8OndVSTMDWtIwBnenffap6ZHpgKJnd9SNKR
mju1LNYvKO4HqDtrZIlVSo50DARQqCoNZFVtJIx1sQPnYn6BlBusWXY+r7Jq7FOldYmS8VhIojJp
8pPWU24khzpEEq9iKpmRZ451KsafWQPu2Xw/QyZc38I5K18uDpeHqW3EBHkGHNz1bS/ijPZ381gX
di97yn52TTn8r4KsJa6P7zoQ2DQPLOxA5yiHAnicQ+6ytEzqcAVLiGm9z8vjKrSuEgIa4VXr/rOE
S9+4RUd1qEVIebAuzZEdQX5AmpXgzYJmfSofwrOfNyZZlOcFZUwtQPt0u/e2J8WGl7ZYK49cD2GW
03YCqSOg6xjYTI3KlGvbtinVitG/TYNd98Ny7pYbuDMjtzS78dgCbyt2LwAS9plAcUyyB4g4CGIC
OLIgonIKV2vHbrgcFBRMDSgDvJOdVH32fkEp50r+yYslc9pImLEKbvMSRFoTpj63QNyXa5bJe5wS
iN0HIR7LBmbTxs6PCYlSOKgWwwtgrjL9KCD5iTlVLFArFo2vupLmpqgVR/RfBNuFdGjazlcvheSq
yEf+BokjIuXnbKF2abfpauQoNjl/MNPMT1cNCsgGsxz4F91tG1UFyAFr2bAaUjyYVLrEgvPosYVG
REtWKfHEZdjwZRHdysItSy5v2HufW9+kqpqnAqY9y3L4R0gzkxeY75egHzNHONPb+rDc3u/Yq3mb
iSbx+xrNAHvQRTEq/ACuvWgasifXgydMSjy6TQs4p6Ju92w0O8/9ZDzS7OuxrBlELvRbwFJXvky4
EX35kf9NrCClTfLsaxEZfdmV6X0xShGDObtUU9FagpZXASMx9QDVLLuqduY2tlJruwiM99JdBHiC
PI9MbBZNjC3Y4jWOlcVk0X+oWJcXV9Afjv7lLOE1+xoahgjeEQ/8zB/B07fVT/crNRWI7n+23hk8
knqfo9INwEP4Fw3SarzFwO/yI9bd2GKoALX70y5HPBn2yYyyzy3sXmNgR6KkzKFJr08ql4zuTCV5
jOMwXPSNDjfPw3CPMUgc6KyBiO+t1EQRsfQpn/irlzs2GCfv/ELDzVWogVbTRc5GxhzQgyYX68uv
xa4t4QnTL9Ymtg/V1UuGAThoMMGaRuxUR2mqqvOjsDi2iTaW0wIBxcPEPzMsYvLrtchCZm/SEcBS
YZ+7F/CnkE6gohVwl4P+3hY4IRQqgGDL8rUn63VOmE97QsP43/jPuF2htfT0S3pBrAfhA4kxqAd2
KME3IswvPzg7dt05BVgQ4x+h2FvbUbQioQez+L92j1cltnV3V6cYawT9u/FKMTVfDJZiFPmm3pDo
Zj06VAhp1xBpX4brE/yUuJESRsV5XhZH9Vyk15MaQ1W+99IXHifvy38X3iKRAU0lyXdOllFzTeRS
CNc/BqK7kEBteMXTjN4L93n0eZsjaP7tu6wlDrYGOAjR5xYlERihCWhbS0GgDtXnV5vba5BdieTC
8E6DCnspn0xQFozkrLHi8QJK+IUO99yiwDAV29iIZA5d8niJYl7FsE+k0mg30MnRGiNO52D6zWrt
ozRMHt4Rhki2IH2jSJIM0qr6pf6Yrxz88qJiYdyCS7xxGC7PCjA/WO3Q8OXcKOjha8bOK8O3ofUA
afY5iRk2VW7NQR4weFHqXo/yaoyAQQIvhU4EEwPNqgA/cACoPBgk7YgzVMzFR3vDFR8957E4VNgE
s7BzoXq4tMTAB3M5anksoDZK5DKGswU1rnsQrza1/baIZAsZ5aqjwaGq4eYvsXAlvOC57DRAC9g5
jFcMnfpH4JVc5qq3Uo8iHXrqtW0ilryU6Wjd2BR1/xPUeNN2BiGnb+b8FwsPzrWC0FIox/vwNJGs
+6wXGErkyc2AX4csHHVkrA+4aMHx9Su2SPtdL+k8xQsisSMhsXxv2NYz233Nlg+cMtACSzT8gbu7
7IYtAy5YJeLz35WZaDShi/1zR/k/vIAIJ+xt0D7eWSmx89XfLCdNRbM6B2oavVpA0xSaCWp3vvAW
oF5SP/r362VfC8vD2ZJ9NmA05UNRcQJZhHeDBiwnH2h3CQvlORhnkYaHqIM7BJhhhMrKVlBDMJyr
5xmXbboR+FWwf9/ErveWvk+Uxx8K/lKag+yvIrvLyt2fpz2i1PtR5ihAl7wXXhQPpHJfsGRHE4t6
yRCWQkgAicPFDGXGfeIxg6+pIqqVs2a3DtZl1BAU0Kw32ovJODpfXNIk/foDrKOVVb6oU6GX90ya
4Brp1c8WOG/qgsVb0Q3vhYgCmQU92PvB/5Kv0fHYPzoEX4iAgrnIq2J9SfJgbAXGnm2dmxfix84i
lEU8b3yuLimfqoiD/ut+RfUrZGKUwfGkgOYE43NiB1bpW1yFiiiuiF2Sknp2uQphiT0jIOzlgKPn
D2oc+anB2mFcjaOaWPurO7gtdGfePAjvri39T0PPiactD5jsVDJkiBia/0l36vz9DmYbCYQSV651
SoZI2C5xANGpV7tZyZZRW4mdFF/t90EzY/gvRaa2/K/u45/BvdP6BUE4i6i2Ezk/mIsej7zMCGvk
m6HA1bjts6QjJyovBPkxJRIiYB9ijCrwtpgOk8Qq7YGne1Day9bRW4KUm22E7GTlS4q7N0XaAKQZ
QCuh0flgB/pocWhWu7ybaLVJ5r08t6seyslU04/t32cEy10iHNTQcRE/fZonLiVhhTwgfGAbO7rd
LDe91kO1VAk2dsSAWPKcHBh92o5MoOvWBzH6cycjApqNqPfuU1HHOx+v7LoeF42Ko9NivRcCmTeO
aOdgj5t3sp9grCqm5n15pw8e1I5OQXVPn4AVFHaCppK9I9eTDRBjB+Dba8nvCgtGF6P44OVayjxD
1kiQsWzeFYUP/FQgttbbaITEsXNGUJG0yYbGuQwciD5kYWYG+ZD4K2PTAsFuQVSGyKQHgL8akzPT
8anToZV5iZisOBfVf/+pGLnkna+5bv6QCg4Z7yVH9Kd9TOH/lyMQMpd977OgELSdLn2EnyMd6uIi
Ed1GhlHnyFOJ1+9V3sc33o8zKEVBtBts+4ug/2yQ+rNd6dvSV1FWZWVEsYfBSXNYE54LGLmbilCb
oGO0tIy8b5AZMLLLz5N2iZj7vaNt4jcuRbdrCI6wKDnOsJqU8Da0aZM/96CvY2dPZ7uuC5Snp0KT
bG1rXANEhWrbOAab6mJTPg4IomczxPrOoKBwbYmi/jRQ3P+WmyvbjMn5cQcas/0fsnlnlUjAg17i
KIdexssCI+iALRlVQC1PBvmXsWcc9Tyfsf7SfkI0gcF4pyUC9Z0kD0zK8u7SxzFlad+1jQezcVAy
OewaavuXx1auV3JdaO3HqlyNBocXyXjMItHo0Tqs82pWoO8q3yvQWUwyD/j3Gk206pwlY5YVajIo
D1m4GNYBWibDUIGQ7G/wz9bEPCVf0N0m/9bP/Ky4D2SjkPa7PWjY1S0oZM0S+zwSmZ3O57KHsKeI
3E4nE9wT8iFOwXL4l9IXwKsiIXHFz8LRkLxWME/pQZfj30ZqnUBa4JWrzr1LMe8Jb2y2ogC/2sWL
CbXu8CPOTeFLZLjo1t9HGJgEgtUxzb65T720TGxLT4ESGdAAgKiRNF6jfdipplWrR+CTNL/vCR+F
lxNTjy/0itK0OuAGu/4JO87EIF23IHxd+AG4+Pk89URmeY/kfBgoGlaakPjK0TR5gKCbTK7s0Z6v
CnomyPyjfyhM/dYl+pLH7Fu03loy1k3snlSgUQALM2+p16TH0AuuAl1hKBoPIHpcg2J37/3/lgZM
5y/NoSQwpmJsHagchU4sk9WZBz7A68B8oCZOMNyrUIT4Mw7LlxE4A4zVK3v1Opq7xPbjvwsqwrAG
aNRLkSh2wEmqVwxEZDKmgn3ZhONaR48FZspqrWvu7QwSV4SfjAep3v+Tly1FYyS+Mws01QXVEnMs
Zc4lfPv5USEnJA5dVATR7ntHvaNuGLpTYC05X72ub59mSx7jggL+09wg+CsVX37T5qITveDuLtLe
mF6GOsMwn1mmKC8ZHBtHRmt9vmjJqCzv9taeTuq4SyHnZo4MVRl9T1RwWDOj0v/dQUZHq3QTIJiS
ZiCZsqzkgg7LiA56W2H+qO7Jppdte+mwTVZSWXXIQhAV/ETIWOyBSPdjHsvNbFRzJRrTeNOes/fs
XsBo5Lk7uHLiH5BJYt9o9czS/5mcnANgQKFhFkElplhqgIbewIQD4SeN5KCyGq0F9KPCuAEpqXZD
yhrOYKRbyWYSMQh/EXIySMPHmuaZl1b+6OKS6snfuSwn6d/werlOadLYgsxDGueDjg6UFdbMS0Al
OfAZCFRcnQAqB7eAjqe0edX8wmQFL42wER7xdf1hjXhHga5mq2lTyb39kHyAJ7/YIPlCphScjlT4
GvqMuiH83McIkYthxN+ihHdLzobD8/8Chjb5vE6QZo7Ak4DjhzD8vhF5M17ohUpZTtg0MiLPPkcg
DVbYD2mE5TYpTqnE7+xrnLxQGLOA23SGj74tbAnxSOZcHWr+ziMgkHLfW4kmfj3A/FpK4mC19MET
HOuHSjhqWmGXtaVoT2N/XCPmzOwRQUEHvmB9JrL5RK6D5T3H0T0dZfQ2a1iaHJ0vkgENu4i7w8Bp
lWg1z6zGEHQsG378zR0QvNoFT+uHP1q+swN9FpuTms1msWfCUHhLWB+T7wyfGqzrI+Z4TIF0CePe
tZF3Wr84urKAIAE+vK9dV/0UUwSunnpUhZKR7bQa8V+doCJwmzT7dx2zpuRSM8TnJi3WxRQyCclc
bEK6nytWDkPyBTvbqtq33L4Cs+Z9AHc1GvldOxwW/1nuhBCRAOm754SjBI+bbgBDY/mU/BQ7QwGs
EVRlLxTa55vF9h9vAa1AJ6b281lmgv+V4EuLCH9wRBbVvAP7gijxewwlIJrNvomcj2STyoRzVQZG
OpBF6bPUpGMRergfIACseiURQ47t87sHAGWcbotoJ94AAyVNipSb14a/VwQZIvHyZJZUXgOpWooo
UQbbEO306knsvgRs34PVZcWlMBY4UyFKi+XXY9OrSd/wklDv7Y8Mu2cQbvFRRRFw+cuVG7WcupIM
3NIrpS05oSR32CVW8StQpclf1614AEBpQpm0p2P4CFq/XIiG0IpIcpRomIYuh5WElWlrbR4quZcO
m5qhqXRB/i+9gtL1HkEEiA8q6+h/yI3hYA5+0ziCUMXQ8w3OtOiJxRXLfgICXyDWTWYJoXSvA3FY
JBeka587x+YvgWmY1K0swKqIKqFg/TM/DSqCpTYK6GRsjyd5X+qsfHES+RxGn0HBm0oUAAnu4PtE
ki9tbr8uMrwHJ/LDQ3GBZSqg67DNxcx9OQRLV+rlX1otQngOSpTS7vKcHNw5UWXLh1+9I0aqxihB
TRuu87CppzAfX2P8/i4mA7iCPPMrNHeTF0iJFJAy5/a+UaJZbaA7iRIjkLVVvamrKAjsPoVU9+z1
R5Y0
`pragma protect end_protected
