`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Dq7DF+QQMUmoH0YzVqTI2uSZ/nXDmpw8Ft2rQVtrpNQEd6n9mUgje3D/q0Hs8u4N
Db8sESkcCiRePiE6o55su22kgm17R844WZvRgLnEiumwNxEu/eXAEO4ZUe8gabcd
gvRDFtbU1T2jUG1Tj9vwx9dVeRa9046wAneZjuZ4AVk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 22816), data_block
BRuBTjmszcHQyMCJiEPVOIeuz6Pk/rwSZu4J0a35xMsS3KUOLPgXBL155fWtuz2y
LRp8HNAl6n0nw3hn9pB7CC8LLybj9ZI8ih9DYCweQn4ZYruSPMh2QN/+lNXRRr+p
TRR6SQkHJq0pohb5LSoY3XgAso5wl0msy+oezIp3npY3aWa5STQkBTE95zWrdVZd
f1TGUbvNCgdPMEAMO9XeLhy4X0MMdJQmkqNFR0oI2fnunWuMPLSz1M0eJpawFi07
FRZMT4XJFPmIBM64jWwjuxBaQwd+dtyWIUjZ1cAIqRresgc4lbTjLOVSwuahqDR1
8J7S18Yn59wGYMXfwq+wBz9DZR84k/UetF4Ff0X6dIUZpTBu+rldjmUYoSs+h1Tx
k0ZuH+QLBriWtRXa4+sIqHh2XRekuj0L0NFe1wFK/l8usyVDXSi2754e7fa1nIM/
2bCXBdkcrmxF6S+86NoUDuxahC2yptWpnBJSeUg95N8M80F/1G2bKgpu58y1vH8M
rUfI0sunucusZ9i3YEzXZMuNgd22D3Tl5+NqSCU/xGdz2l+Q8pPdmgm8O+mILAon
5dlshy9S87l8ErtHCbcoXKE9185Dcc/MnwfEBAYA0rD7VcnxXabzSNbn60kOwcaJ
gUan5WvoupvhNeW6vu6zUT6GStQxyECRye48e6l+qkHT416Ho/OktqDiBCJ+GKhm
uBZMBrfJzzbuUpbAhyKVAqLwDa1m2JidQr1mlkhymYv1v1QGHIrmLlf5+TPQ7GGZ
obXcmH9Ai1uanUd47qGO/dYGJuswS6i/4nDWjvFQD6xGYqmCQ6/zFcZ22DmqQ7Lw
NmgqccqSNNMYjBjBwoNjUK94HDNiHKSXgFS6pOXFGYwqGtOMph70McgSYBSfIDEX
3cmFQRehqfHNF6yoUbA9QwjRhXEXACXLQGLr+c/H6IHWW64A6pdn+3n8y2PdaTh6
VDr/Oe5SecbDblDaKXTNu0aY6O74lSG0EjjBufqbyjCe9BDXkCNIPoXtawSOPf9H
I5UnHzy13YOMI1DCKB+UbNF1zniq4tQt3tLbGX5BOGhJmvB+Wy6ll1752zB2nB0R
qKZ+aLoWRsgZ38qOsbp4d1brHO4L57kjjO9ZGq1SWXTW1kGHeUN2SUKxu7tm29on
+MqI7dFKO4l459dXM/WjmOOntpMzu/wFlk1c9vpwG3AJIYGxoxEBqBsRyPH0yOr3
w0oafOTcboJU4cGDC4tTwvPH9+KHotTpzlI8nzihOWG0YdLNurZLlyVez6suKb/1
Ak4GsmLm9WBOYmnSqqiUPRF/0t1/AcLdRL46ucynouwBkaYVvzZPBGLEkB0grsb3
vixxL1owZX7vgpIeRoL7KoPcxvRXAiQVMY0HHFDwP+/7gHlmpBB8rvfe79+Qm/6N
SlZM0qulBL1DxO/HKldYBVuERFgcvH6FSkJgWudhRBs34Cj0Sf+el/QiNHrXCZqf
ta7lY/Ddrf075JKjP9Ex88PHE20D8Rf2Y6vuLqQceFHR2Hj0BZGQsh6NJ8TkfpD6
9tu6Ftg4E83CVBNeVGnscgvFMxET+En/r44K31a0HbionG+OJUs9K6mN7GQ+xz6r
zhFH9dwdTlbaSCDplB/IEw7nWc5SOPdheAjf735dXstT9H5exxs6RnlB/V4aVK0N
vyUACJf0zpzn5Znyb2tbfjKRVQ2V243/ak4cmdnzSr8NQhDduziQvy3IzABPxvyE
dkocCV7Zs+ZTU+1Rpgm9JQ8YS5sM+FV3TJ1XCZI67mzipB/Isj9hbjz8BYoOjMXw
yPx3RdvIGbisLGWl9XGQK1/gSv/wROaAamhu2YWf6FkI0/fem1jWdYx+2g8Pt6dC
6Mv0EStzEXiZKr94HmJqy5xvBnslQWvG9kDnOUn5N5sgXcmrMRNJREJSm6bJFCxc
mpLV0YxdFHpeZOsS7+rNGvkBaeO6VIqrdh30ptdxCv6wcFGgYSXs50LXjuPWUebA
WI8R1091eGk6GEzJNDCTH2wu95i7sImC6LGn7VJ53Z29zEm1anP5XwzpDsSx3Hve
fEfziK1Bru8X/m3tSD5ilCIgeWH9Xv3ix6jQehoTAhuiLPfZ8nfzkb29XIDqaqRd
0vSAGCGPZt7PiXCseLdJE2bH6QLmFkveluCbE+6kGxsniOzO1/0NBYO/v58XQCSp
DJPHCVfaNTzG92rLbNk0fIl0wC2PfyVA93YxIdHvNFcl1yxAjt2d98kFufi4uyp6
adVwNVyCirwG1KNh3aFRrRjOJrxZQtBS7yQX/vv4kDurqZsmi8YSytb8RvnfIe2K
kSTQbb/UQgQE+44goFRzw9h5wKeSXf/FW+W3YsbsCM/z5oQOl96/9HBtkJkftDCV
rPlbY7hgbHcUccUb+LWVgKZYbJtdu0CGCfEdITJ8anWRvT0hPYKBNcnnlsEXqfgE
TgkWvyZI6ty46m2Lrtb5CHXU+9nTFxes6aU5J3fl2/CrJcmka2h9QIPDKAKrgTbU
ef8goQ9gj07axxS04LhCwgiqKVG4/WYy/h9MD5wnV3dN4Bv0+uh6fUWV7XqNhWFR
RKqc1WPbBXjL5gjUeoOb8gdZQ9B3YoYZmvnKvhpWqAjsr3+1bUnJOZI6WLD7R+Wc
IKQKdPy3nwlioACpkN/MAVcSw8YbThuXmTq+C+zfyp95ymBrxCBDFz5bRHYYt8Xd
zheNRw6OpIOZhM0GTvH/AAcjf6sWs8P775ANyRlcSkpHMtDmyGemnit847fhuWzj
hNhWiV56hR+bqT+1jq6emb/KEAQrZ1Oek5smxdM+Av5fuYrG0jXHvjcpw+/kZpFX
8OS159XfBcUksRkr1wMweEmyQ/vn3NNI/roqYwD22Jl9O/USJ+jIgWB99eba9lqc
a7Ry6FZ+OxOf+ah0sG59MEjX93nE8DN0gMYI7zYiLNCDCQuzhQ3sibNi1SS5cEcf
Y+uDdAHr2YEuxF7WE2QMr/xtwkyl5eqbsmrGWZgumb1lAmDWoAwqXrn+Utv5xNm7
7OeJiffVDqsbxxgAoPfY7blc6xtghOKLLgMxILX2UMhOaLLL7YKnlCrx2vp7ya38
NOhO8EgO5URzjeBS+3aiBINukLlFc/0V2KPz1HlVcU1bK3Mot7ZO0+UTl10evQd5
ugEXBRMyRhBGgkTtZek4/98Gobs5eqxT+JLrNK3nj/5k0x0h+/gD9wceNmGiB5kv
D1CokC66nPBgLRRZ0s9jIq1k8P5R/JS2mq7heAM1oNVoXy+/esXSfrb+T3iiHg2+
LFpKepsEpnzCCuInIj8wpAcoi4R5SemR72LjH1TUjGbk8rT1ZLroERkx9DiAhAKA
drXjtcGD2fUdRcuG6WkWOB9FJenK60gv+pSqBcRGfSyo3WMv5QFXCAOTtA8XVnno
fPb7WhOgfOHlhfItAduwzEp7xfMxFXSpAGWY0xe5LYnwoy0sFjeGJbnsZR2RGUiP
3LXfKtbtuQ5m8TwcD7EHSzK9R0bVQYkRt7GApj9JWBaCQfKGXWq/d/rXtrdHdjjJ
sXC+8I2N4vSweSmM2QGO9woN8NCMkSs7/oBXNCq2Rz2iyZ6Va7feVFR292spxHh7
SBjOliCK8zV/Vlj/4nNYgRJVeBAdS4WboP4a9sm5FehoXO8dft7kGvfIL+ewqgEh
CSekJJMjSjCDIXo95S5WxhwFiDmqrc36+sAq+oG1EDDZAhngOcUBB+xnxOvmgM3B
CIjYZOepv0KYk/5fRdd3D+Jk0G5kFIaJoJJP5crMtFBn5R9HQxbXaZSM4sJfFWHy
A967/oMohAel2YEhyWaKLC7JAdzl52CExi3oJNinkephilB7hOjiHIaQoGuNeNww
W1M/HOMFpBZLrp65G91+nV5taz2jxpbpcEhAirxEgUgQx6uzfy5Rl9qStl732rBM
iSldsQuG7JYX0doHPjJJTwJF4YlGmvnHyIv+i2q+NYTRdHljTDvqUF7/4/q5VH1o
EoPAsGL7ClimV+Ue9V8BaD53kDZuiK2JkLM+rwvMIFytADG0FxeyNei/htDzuyVT
r56EdrRqLYhqeQzg3qazNKvIDz1qbvEsI6dHONLKJQuZz7aqC5QdYS3kyja6OK+I
wDhXmVTdrp8zVdKIb6AvbsfzXJpsb1XANTVhazk0JVQtRp7tpB6rxNC30So45t3O
sdH9z724p5sP0Ik66ADDA6HXpwLMKvwEe8Ox3QkuC7+R4DTXUj0NNpGBLkTjPVp1
NfTYE6iwFnQ+MfJX8UEiqyHVUAjC9bjIFHWntuvKrwoon1rKE0bEflTstqz8+ier
lLJCWe1VgsQkLyV7aijxSKwVHaXTXBKAs+7DPmBWmCpukXtYeGPac/jrHiZM8TeH
zi72gFK3sd6iqQ1jYmfu3JYh6j9VMW/g5j5WrkRkvBTt8fA6j/gJ899OWDFPpjMN
vpJ78MerOw1xGRQXbRAkIW7P+KANClVGjpa/dLt8OMd+FJ4zsf48ZKpPmyhTHmC8
STdRykysXhAVg80+aSJFGhYleaY49FDaIlJw6Uqj/gwQiPqBNcd1Twv2E0QkBBcz
XirrHcVpc9zp3WbBewe9cpT6qJ77NDf/+zKAq3a3D7OMYGC9egR8ESYQ4FfkwEbg
wXcPwonzu7+P+227TFbtA2hHemvZwDxeoYTZbjBW+gAABXB63Et07njsMNpArSfm
Wzxa+HQ0XaK9bHFumnsqXMP+6uQLdJaNoXyGFY0k0dqIfHj+lzOQ5CmlkBwcMh9B
o0RJSa9LE/29uyY66u2qBnzGmqHg+rSqweqP3G0JHjIFk+h6c5vlcFTEkrgQdL+u
NJoWDPKC/aLnhqhX8p6ZLVMiZgGDoc4tUGw9Gr8BiEkTsXb1kar0vbkBpKtIXWHg
jnSElVYDIEsHUmeHWaA5Kr2YJ88148kH71poLoWYRNHeR0y3slZGrvCWNLQRACLk
4XwIqpPO5rqLoSH2CnbJZ2q4+itkZm6zNvNZIviI4N0MhqMOZn0p37CWgh4FAsWe
1vTkCm2XFGKIlID5EDhuRaIuDhgA7pELW3+cvyPGcNJ0TMGRuBJs+N2XVsErMyGW
8/2S0GeZWNiJcA+H4JaVncCApvOxqPJAk+TJske3UKBMCFhZESTmk/qyay5z/KK+
sdJd3TiZ/Bb4cnHc1C8JXBMSvNsXA93zNoEj8pxswLISDHGyAapXv/p/LTEqU3cF
wmXZbibG1z82Fh8+S6N9ZZHy8pD65AfVsGrMjZCpEv3ghgG76SKNUqRgFgRoZ13L
xHgCdEevac+K8iJA/56Zu+6jT7You1oZgMCUByP+ApZJfgd9rAdJGdOvLBZvW8Nk
Ghc5LiP0IN5cT+aSlxLPLn+xTxF3zq66aCvV2wyfhsez5moKlhvXVI7aKQPWLOHC
m/qCBNtXHtGO7uXpnjsnUTnguIw591DKr+FP/+hJvkMlDzvzztylQIdOTM7hk5dZ
3oPa3PcVW5Ovyt3ZKqBRYiAie97rO6A+io6CmfbVbS2BDFSOalZwegmAYMHONvZv
iOVYu1J1oloWXMcu10ng03ekhd6PYrM8jr/69n6U99Em6SpmmnxfLkbzMSlyZaBK
vgi4nHhSJzTjBbJrztoYdNFlKXA6sT77sWujU84Tuz3+Yd+Bi59wLlUyEM1rqX+Q
3uyhNLq3nyGFAjw83XZ+d3XzgLoYKDXjJL9UkAUQzrYgOxhvfFOjNfhuxw1S3HKx
jLvydEeW6bsPI5YcksIbF9rVySF33McXZZdTtXj/oRGWWQ+nDTyrjXyfqOg2boHe
oC4QbnsX7AkPxK0QwI4gB1SqV4yvQHAHJtiRVdNCWu/e0+RiTK673PmomEW6hO9n
uJT1PZdU45tNvb7Z9eTwoX8qAHbzwPxXi7gSdT1oJUFVhfv8r2cR9ADCa6WFyqxB
vhVdDHtRqpq+sx8z5NGVFUIg2tQQUxOUISy6qpBd9pW/qBTers7FaB1EjSsFlZdJ
gfNmT9MqZlYrwI17KVBnG6HR6kh7yGUy8/eufrAM1VuU6ZTFk111kFsVgOzEZv2J
j3CpNzl5zflijJ5XXCw1fgg5PNXo7R9tK9HMUtcLxvt1KKSVziThPUP6Fy/U9gFa
TkP852x7RuSBf6zvq4HgFlsM5RwxA6CuRj/kVLv1oaTuUMCNhmV1tZE7Um3iG+2H
Sak8SaKvAIaHMuWxgeyNujJyx28HdIzTpTmRr6we5u2Nzmp1c3LvNHQYq8MQsae6
j6xIXMfnAtdrpzPZgbjt0pqAvHT/ZHEDzOmuhu6+T9qtdMthoue3/VDGQxyifK0p
TPzfLABalv6+QiNnM7KCwmdlULWlxdORQ7dm0X6tkgrO+YiGm/4I3HRcyAH4G51x
FIGzTndp0bo90yoKo8+PU4kqDnb4X+Y/hTIf7JAp53yRnH1IYJD5+VPtmSoIczFO
ta/FvjEmkUd0fFbPQpAS7BG8R4ztIl9HWcBG0DexZC5t58LszoKWEib2RBw+HeJm
QmDwOSko1U5jouWmQdOKa7aQ7CKWrb3LEtLDLabAyyNudbO/x9J+rk+p19pZkY5y
Vy/t2xqXJGNoZRA/1wBZxMusKSTMrcoIA9PzZ1D/MbSPQQW9l4WjfsI6xEonkPnR
VP27oDaNv01xTs33OkQMR0eSF+L1eY2BH0yrgGFdZIqkhFC7jB7zCpBad0lz6cdY
1CMcncwHCkgM8ZJUXPiJgFqOPoFOFonRaEZizOz9dagEdbtvy20t02X1D253auel
MK/BXzekGWxaTt/yuhjc1jAOmH4UB9HVcwNM3+Q3QGbJPG7kKPMvSdPknqzc4Q/V
fS/YHW4U9pQI9Qon1uO/U/bGA3np/VCihq1YhblwkBpJe40HpYapYuWHZ4A7t1A0
xFbVEDSFz4c4o0Eovc/fFA0hQa5O3kamd79s8ZzyqeHdIY5GFcgslTw++0D46x8D
wCDGEquUnSu9yAb0qveXs6uu4xOKn1+xobpDDjirZPGfNXY/KI1KQz8kz3ePZq6j
2aW/JHv+e4wuzpWaAllx6HgphJxnVaeM0l74zWOCKKKukPTetzpCXFpNIp4ruQ7S
xmbvef2OI7zMWlT5yhsKMOVhh1hjq1/r8LuDJUQ5BW27w8+r2jGhv821BPlM7+dv
W2Zy/JC0dQxsRB9xiU04u8y4hAr7cVzcc7LrgAbiNiEAvBo/njz9S2T3oprsBX5D
MSb2j2jOd8wOYAjWVYvuaBfVOvuujQS1h2m3UAV5/q7Vrcf7FnhU2ME/ZtstJuMK
YxHfjLM2RgETzi6/re6X+9+725DmwwUkNzre1doAu9LxTeQaiOHmOBqyKgx68OyO
Q/cp1+qOmOT+FXt3KYFbD8FOK5M+ga/BfrMq7JwtfFuljoW2+fUGiamckeo+YmCY
VUUlS75g8PvJEpLgEIQmUHLUUffVR7HHOspW4BtMC1BhZUNHniDD6ADGYjLXMVWX
BRYJNPRflnJevSnQn1MjxViqVmM0DBLHAXHVHxUnTcE/McOowXOhOBiPPMDvjfej
2Z5f06UJOU9oAyrgwmOrQl4PpPlkGg3BEaLdU4gAvBygdnng07MeH5Mu4UFDpA7a
Z+DEZqlxAv3Om3PdXk2SI5Trm6iQJJaicIQSNH8wOocq6X3IvN/p1IfnGhno1azG
mjfv/jkIF8CyGiaT9duhH42cbVapuYTdxsoEptYG55aU/Q6d3gORcWxawFBYYFNp
WG24uac+oGuk/DIKEyoEf+gT+LBRr6Rfy6DLHtjfcZDUa5dE1/cVRLIDZTsgF5Mi
bMQWG7aiSp+sVsxh9bJs9Tv1DO4t3jhCK27H8YBoAKBnNVy8w29eK9ShqPgkj0eK
TM1tBASzEPWWi+c37rnh+sjO3Sut9wg4FzrF7b9UwXHICQeY6UUN6j6imVl/wtMx
CLwxhTdTaahwFLSD0l6VYHwXvjfVR2lRM9CXbls1WgngSU2nM1jorHOwgx7GT/gl
4GyS03j/02PvgntHi3NpmbdtM3KRwDVR/vdjnwysi4kSNellIeVX5ov7jhNihZNF
I2FC1rhXg1qG5OUVyMrg91NoQ0V0k6CoWI96V7j3Gi4XW4ikfmkWLUYJfi0LFjlF
uwXooAQ9/jLqEqjCkuiZ432ebSEq73FfbQ0KjLzEHaSLe9DEh1Kkqei21n6PwPPK
Fnxw0D80TX8wZfZ7S3lc87+NrGU7WZo6+RRViTHP3c6T0b5BsLD1c7Lj4pz1BLfE
pyCbOpDFKhRj/eUFYnNHGMQGGT35C+6zyi59sdSytu0EPKeeaCGQ8ZNFZrAn5KBe
VCUfzowGCc8Mg3I3yizyR3/uvbqXP3eARyNJOLlJofZW3YivucY9O0CwmL1EIX+Y
M0GzCG3yDCC5B87xVS69/CFalEQ0+fhXAr+9Jy5N62RfNmtuzUmnabatB+h5JiTK
jCrggDe+Z+piWfCOsr9RWt4vDIwt0fgWpfhRTyRqqYc6OKTLrNlQZ0gINN0IrIF0
88hBucqkgEhTx+rSRfXzAmVfRpIsEa387YPDG3Vpexja9HikOfgYMhoBwiTy8hCI
9w6LGI/JPN/h9AA/GrVKm7RLUKntkxQWoiHZM4uB9EtWzMsdJerQSfpIenU1tBJc
EmMj1VaET8Io8UMqhMWwzvPCIt3b0ZliTQBrJECA+qzoLyCmnthwNEPRx2q6hJIn
QKl+/pokR2smekSD6fR//EAct0bHV23QlwEWF7535gf+avzylIqI/1L4opZgnR9Y
87PzaAtgXHzOKk8dl9lmKjDcTMuYsF7yJQoy8Ox7EPc0dz5wbOXzDAmhwXdPcxeF
Z3Wwwt0B7wE7DM01ExvkEdZHnukIISyQVyNsKaqWhoYgJ584JgHfEYGKAOnsStS8
pD4fedHiRV2QgBWbOTyjbA4vJeWDQqwx8h2QOMP+D9NRnaMNkGrDC3A5VUVdDFTB
q981/WdBkz9QkliRbur1DF7lnB+lk8+raeWf85+JlBKAQmKZCqwU2UBCxszNFHl0
s8xoZNS9mkF3yEQH0q711xhlALGXi0gItWaulKjOutDPLBuhd4DtvCqRU1avbZ8b
K2lpK+paYrTV/RgDOHaCzrtNdkkws/8xuo911EFiJJiv6v1tgqKbPA/J94m2ED6R
Dp+7hZfrZb1KSXgn6rhIXTCam+oqlmofvvJG2+RKHhu7yKiaXnK5P13gl/tXqX6j
xYD/F5FXG7/1Zy2dEhrwZHwVY7Ar0lpG/XLee8HQEP8PZcXie7yEcI2bflSGNReP
kEiXgMfy+ymdHHmYQWIY7o9Hw1/P8brokLnpigUGxGRVHwld64EB2nROoidCa4Yw
A2HNjoYtFxe73R1VrdGUjSBDRuhX+q0lGoM+J3PmXQ/zs/lzjyeT35g7I6CnF93/
33vqXUD191bGqWXnmsdq4Lh45N67fhGC+oZdpvbdhfRuH2opqrGNQcgkRVCr7KFm
6oh7/dErGM+lgUbUrmdmM5EytHUwxL2gLX7bgKnn9phjsur1YGF28+pyWqDrg23n
fn/KIVZ06QK4e18+s2KYphuv1bOmXuxiTXWp3t3oBcxDpr2ETvGVtJWbYL4jLH1W
OhvJj2BENjEzkF6eQ9/tGe2d+wmo9Yp4Y48VpvMLYALxJMsy5uF93uwjLNSyqAAP
dvM7n8m5zxu3z71BT3jWM/pPBAtas4rDD2afQ/ZuxPdWIFLzTp+CeC41A44dlGkD
YwEoT7Ign8vkp6UbwLrDtRsroGWxH1v7mF2GlPEo6R1KZJrH6GV+OvEAjHNQdd4U
innZIjLbK0iW9GAs8zMKtpez9yA+bzLN346ojTV015/KvlrvCjGn5h0ktul4+ycS
JP+nvxdJjbfeu0PhsoiyQsIdTgH3kRG+RqfwZ0EzvKLydu+gs3EoSJUytQSYl6oy
WgpoJ1Bbrq5vu34Ee3x1voyVNZOZxGoR4woPybIafpYkVuuxEnBX1dDi63Vo7kp6
gwsDDnfm0v9yKo27m0ud4Tfq3tLjgTcg//1/ovydJt9rAb58UDkmU5R1rMtXZKOx
sQ2Z6AV0n23Ju9gzz00mnvBDX3vRYuKykI+6i759JX+3mcum74czIt3f7seOfMdl
Cs3CLCeM40wC1S9yjXOoZmHNZAB6vu3vBjdt0Fze7f1z+e6Tf+AgJOpXp0WvMS/l
Mi7gYqsl9c3yiR9xJMmc0uEighkkw/boiFA9AiklOTGAADSAS/jgWgoiu5aAcRiH
AZFUw4gvesITmBLJolYVUFi+Ld5KGzmX7mBbsw+W483t9AaPi/cgHXifJZ5ancnS
etnhEYbfXQ4bCMZpokQy4wDtRopOh/GNFCZ3dESbKX47qycKh3yGnIqq4md3/u4k
LanuZ0acdu4Pl+CZMWqxwf2ho/b7o4bTtkSPC8MZFChL+WihXcpEX46F6UPPxjSz
u57EiaooRpBvt+gsz7KFD5eUDM17ErZ84zL1d+wMbDqveFoHUFX97KW7y5TCRtIm
B8rF8GyzDMLKdsD34lNlaqHwYH+MeUhmthlZpHslMOmZa2VNuSHt0J8veARystty
aiJ7RANNPHRq4yyj1CMQT85/DY/fj/hyS5qd6bHCFYsjIvsekOgvZdF9/JBjvWYW
SmoW3W3IEUGnDE5uKG0ctOVgRk5njnURSzxlSwiQrz+4O/v6z6m9KMXRvxoCGbRq
5e/4j+ZllO5tpz8KEewU55vNVNN6+k3k0USkylKaBTB9p+SKWasctpPuOpT208A2
k8HnCCaDaIkRPQ3Q6puQ7mnkkRYI9n01Uk6HYSQ7Tv6ST5NhiZsMYzqoZ1IETH81
ZBROMSyaM0tgLJCF3N+jYQ71Z6Q+jMKjadnHROW2L1gEuj/uH8HMv0xawo4mwO5/
BPuVSuOu4esUP6abZtVcwUE28U0783HX1SAbnAz1BZXA+aQqS/lJvvZycRVrLVHr
pmwyisvq97Qe8SVgnNB3x7rotVTX/XQFtRCaqLmjjCcLrxBewqHrYT8DVvrGjYVc
H1A0JqSCY9o8wgmRf6td8m54A2wap4IvR0taHKHjRWW/Ad1u+MgOrE/ISfn202OJ
z4tQCcQXt5PCiWSmc2xmGaa6Flw72u24TQy0S7qmfIPkQBiC9mCkwnUhKbnCU13e
B/YsqUqYVWXiuWkhmL/8q9IAJeq22HF44MTn4SevYBciVuQJNOtjjzVhKl26Qll9
w7z+9I2jAerkazaG+JaXaly8gk3yOdfIZMk4PhtEW1qgTvl0EmVPE4L9bJteBFOh
zT4OkVjUq7LrMISM+R+EawEm9f4tRTPcqqXNcYBuSU2V/37s/3TT85PQc4Jxigv6
2aLOUxBgjCzuczkx68+WfOU5xygvGtIXEtPNL8/wbdOswuejslIr+Ku7fNLmjfE+
N3GjH8lpqt+aNrmlcJ7XDLgC5MxoFQz25/8r4IGwaxjXqjs7eCO4nhSjCtUqvvRF
w1FCHNr9qDkyMyZxUvUhAQ3g5e+uy6yDv4EyC3VEP6+Pw5Cj5vkLhJ6GW/Jd0YZq
8tKn84DPaO1OY2aOJAud5F7Tj8Ap7lkBx/moO9bBHTe0GdZllP17W0iR4O06dFI/
m1d2LUIkhmWb14xZ2a7EL3+rK9KS2keTkWHbF/JOTq/SFzh23xJ26k9x3pqpcv7T
4Zay1AUCD51MA282TaNA1ZFIFFOKtfC/+FUcyyfgflS5bOksP17GTiUxxAxmjLth
sWfGKlpPbrbFmSkD0oisVfAv7h19Xfk7b7JbuPEeLSnPqSK0objDoGkeeCNCHpC9
k13amYbwlz75wQcrQaPwfu/hmOntNU1oHrPaZoqRLmMModVGH50QAnb7GXvybOBx
c78ytbHHCdQ3xUyFe42Y1cDDCd/X8sFVzIqrLpmhOkOUqT2C2PfEJkLOLEFW5y1a
tF/GDjseRAwLcmB0tvvDK2tkc9vLp1DrpzOR5/Skffee/RjvZujJZ73fpJNl8bMD
975cnDVmKgIBUwfL0bmQRG+VMUEVQCGcFqadlwCekJggsEknKkbf2JZIwTn2kWa8
LbUKeNE7qafHcUM3h8pm+qKRKZkNNbVYr09Xhki5cUgqmT/oUdyAaeFK0HveNnDW
ISLFBZHelONynkpuUGEiSx6XwCUSGIRziPxLbh+ETSjmgc2oh3dhZLDNAUuyWsPf
s2XVikVYLt/3Ri7R38O5wme5BmsbhiDfpIBYEGuI8s9xEhpWUBoTiJWAWBJMePCo
QH18z2n0qYpMaO5wUPWncyyAn7X6g4QZJp5p2ywvGsUjPWuYcLeED0Jf2XOqhcLM
262l5q9EWKXwbsHpVLu22+zVCHiYjKpO+B0itoJJy16bWX08acOnNrsrf2rBLiU2
BlJwME4N29sqR5FYoSNxG5GVhwHUtGyHqFvi7w8OqRSm2+jc+FmhzDPTOolyl+wD
o62S54dJwy+yFk3p8ohN1CQYL47hLkYU7oVcY9Ie3CfQKHGyPbk53PgObCzvU5U4
fh0hkm9aFM40UZWmmeYzCXMW8LMCdRnsvw6tSHA0RlVcHgjnE7loKGdwPEcTWi+0
tr6/aIChp172b6sbemJLyXnLsnTlFgkGZH9NWYuNNgWPklzlHoUDNgHa3okUSypW
FYnJQrjpwEZL4+KLP+4PvECOn+VPfYvUfprCN9QcfmKrLxDDkMssZiZwOZARKcln
cKyQHMQ1juiRBikYq2IqlzhGORdj/NFxPqlz5fVxadtntVYjcXKs7TuOXEztg41L
P37n3N8IP7YPF7YG7CDcVBRcKiRHmG81EQiauC5VZWK9uP03PEH4+1OM8KsPKKpG
WXLlbW2mX1JW9K2gvUxx9s2/MKRosiS+6BV3YlxtovF0ft/ALrjK9iecBoqJpkBK
RUs/y8bPjAb621agSkeWf9wqGBx0jBzp2/Ux1aBF11JKDwQy53BljSTPh2k4l3UT
5eKG/FRzSuJoyQ8XAzgnT3FRKnufcWP6h5l9HlDk3sDAlVnwCtqC9NxBaduQGrcv
N+0trWPx9tgP7C25ITqNEXIJp/9IonbeHk3ATTT2zUcNTqeODBHWLc52rQle1HA9
MZTjN2UhM1UVrDAv47YfP+uAW1XsAd6yaNeEED5Gx18poGVBVNESRB9VCz9HJzBc
QRLgBo5MM3cZjIzuXkXluOpg6K2b/oM296Dh3siAhhRTw3+k+ec2hpJXNpriLT2j
jdL+CoQ1ioRcxmsoWuQ72y22qCt2mbT7hoyKbK4Hi930jX+MP9aiSDtj7/EDSxYG
/K2Rt2n2M7UZpJBQUkJWlAL9Ujbkdp81E1wfN5TWiGRLxrXu6bY/Qt2knm/Jk9dm
4V3JfOeC3rr033XDP+Mhe9qpkbTcc4HqyHmqsMYjXUnZsel02FdYaJx/G2/b9oQ9
HbEKgzKygPlWmiNPs7sO1B7Hh7t/MNmTF4gmkkLk5tY3M8525ZF5fM20znwnw3/z
FZFaS69+tRlWX8X1gOOqt3xH9XQ0Rgv4rVEwhPo8QEMTiyAgpK7eJjXe7yo3h4vN
20jBQj23kF5iOHkKMVMcwFYX7WJ2LuxzqOqF4BHOcpEvndNKOjX7bxgfvYUeyfAI
Ih9b5UgOHDDUtGYFytrnAMD/qmPZc1b951ytV+uiRkoRw6YgAnv2ssc3YZ5gce5y
8xwPCHfFJLesk75pmAZfP86zd0UZOGZsr8dMm5cxgh+mFas5ESDtwJhfnuHd9n2a
AV+cp+IYk9rqSiqWTa6pNVhNo+xIVR/4uLDbAVQIAzJfSq3uxfq8a6zRsPdo4NKW
R7P37DKWhpBdftBJ0Vt4cjfNGhk98PfnQZZR6X4lpYrc/PHVxUZAb44zCt+ZoXUn
ayLhoNaUpj71ZqGx+uffOuMUzquo/n0mNvCyPpjzMVvXGe0gA5HdkRbrfZfqpilr
jLBC9i7iTQXnsAJW9XwbnGWF0iASN4/1rZgCJ2KZzvYyFlCz0fuHKKh6yXCUUJiy
mYFV3fcLNehHSbjsRaQGzuDskS+W0RSyXrt8SVbtyugbNEYpBuYIP2Phqe4COgiY
iS9vI9rjxBG31WqzY7fGTVFBhn6hFyP3DuAElp4WmIw7+b3OU4OtR4rmsmCoWlkj
c0DKwbh2AJsVSFJzyY3DwOrUObtbUaiTUmUN3JP5Is1QxNe6jjrNiRNoTGFvphop
QNX1zrRaUq293jvw7P+nv7oLi2xQ7/LQ6tqtBkRBC6bGf4KyDyUBt81fFZ4Pr6nf
Psjp8nBTRS7skfxU157CLPenM0sAsPaSROU1t7OA9PkYQbnkXFuWyosYrTmKSLNH
nRxxYDqljiFODoYHfKztmfMWWzOPfmn8hW2GkvwUUke/WYclRDkMHFynCWPN+Ymm
v59gdlwIy0L2QUDR3FRWAHHI7UDAXPnmSH4a9WUwzALYwvQcwKwQb9qBoL/ybTug
gFsOr42XBwYGFah7hAKstJcZBJrYDWAKfWS70ZwX4mlvp4vwQEYYdZpcWP25g0wi
ewQ4eVPG9VSMduzInc476o5IbIJ3PT9b5T/FmOCQEVnd9q2g1f+VTUxazNEG/dxh
W/67Nxovc4Dva1EkbG3M9bIDWEL4mWtxjswNFpZnK26TXV3NQDyqaSnsd09isYLo
P15/8JbHAlI8i3vW+5bodEUvaYuklWO1Yk3X276KoDPq4jddBhHetr+ZzPM1zywM
1zRaVpfqLWhac1T0miT2I7TBbQveWsWWRYwuHWIb6PrbVSOTFH918FoDuv4+aYUW
+KZ2lcI4YV0sIDMeqxSFW8VYKMmoLV/g9AFIAhu/m5yeQKKwwOvF5dvy1EKc+bnn
3zSwx7BRljp+nanyPqbirGi++Sm2lwUWA4UyMmjy9bBCjdCYKtM6tAA4Py3gjwJc
I4H4o8UX8v4Ooxxlm3Ze97XfxVR19ngWxVzKnjQ1JT6x42Mo5nx6D1mlbsksNgqB
tHVG66txuaXhcx752qUAqvdqCBxF5oMinEKAMOaKofBPr2BJEsqQRjE0mwTTaR+U
QED39AV5KMZkxqQEQp13e76sUpMY72L74Fb0J0mtgC5QfJXLrt3/4Vtuy6Kz1bcI
w7ydHSy2PeXIkD0EEhf+fZxpMQNFnRyxbZux73X6BzktMyx4XEW96L+qn1sgJ9sd
XGO7XNJO7b1SZCibCJrMmAU/9pGVdwN+671ckd9IBRyd99gYcyM3wqmsabEaLL5O
6cnIObSsz21kpmzqRic2eWUecgQUoiVfIpZjWGHSLPb1xsvMVvye8OgT+H6on2E0
vZWP9X5M4zfLXRecJ+u24qr9AbyDRw0nEXaA4nG2CNjnRpYyFO8Xe2wCo3Vp3H/Z
s6YArbHFFCHMn1TtyeNrxbZsM7kLfiQp9DlMTlzS/qgvZ2+W303TCJZcr1m3PA4M
O62ZjEHgQ9Ah0IQE3kQ1Aoqn6TURWIJ0n0EP5t0frYK0J48wvorYj/L/rjI8MYYx
DCwFe+Bk3mL/dlRiMM+vv1YH/K+2d6koIRyoAaxxwGjEncCV+eIk7TrFGxyalaJN
zFJDee9ya7Rt/XBEqHQhpAbnOMFwEfYzwUTuNg7jJe8H8bcx5/zJUYyURBa6hMsn
Dnc26o8+FRabgmYjdrT78av/6HsPA+OL9CbclRj4YBAk3+aJXfXgC4rJlRuQZ8X3
3fWASlJGsqA4oic+7HJQYm+VvFSkAJRwSli/1l1QXepclnXgptj/RDfIN13mZmck
Hdg3K4ah8aqxhO3dMu1HHI/iGTu7/l8F6MN1ik03ImUWjgUVLaOyfpOlUU3V41g7
SxwxSj4K3aYwepvxH8JcXWEVAjNCgvQzXhC1yagVftXSrf2v0dDxb90/SAzIybNo
tJI0BXKJ/EPbv19SGx8+RL85rKdw0ouryCSX05JRrZYqhLUT12pUijlL20ch1X/a
EgPQhsIO46NliUsKQSOTxGZkYYAQVXbsNwbxC8Oz3n5z1cta9AlpHj8tOi4IAd1l
KoAjjuQBExVSEyPz+fr1BzTY+BNBlS2ljJk4Srp9DG+bNOMxdauYrT6xic23T8P1
7OdNP/AS7XffzBc6rie53Ma8UTzB385CPVsKyhsNs+ACQHPcduhBo1hAQkBVaVoe
1ANXDJZKznMKhIaDfkcHcbc/rpL4ZpvFOiSjvZbjvSXhKZjugMkKNUdI/0/jVzG0
bme5cK028+7jBgdbOhla/uIl7GrAxepT7NfINWuXfVH2lsVQTCxLSWjpfvBwYt9H
wSo2chfwknkvUfd+dpSTtAddcjyor8+Wg07nrWmP14MWl4Qtkmr4YXjVjfMoMeox
oN/S8Q92UYwOh7HOlGVM3rxt02cN7UXpcIP1jToE0uvqSnmw2cRC/jh3vuLl4+Nd
rb6wdJ22U1UftKd0XbSK4Z5DE5sG61iWqONNSRlDyQKSJcEgF5VPKZcHbCP3hqcj
wwE1db052TAN8s7/E1rk1F+08yGK8rMFFVMMAIY13ioHFGBFvgwrz38495jajZcO
JnJ9Pe9+H3mt3dYhAIDGOntLJGuXZ1kE3ymfjy0q5tJ7U8PVVIPOpbsLATN7TueU
0UfWNGwpP/Z0FMK0XJ1+TDe/RTeifcv25ghDmyzBjKZRByhIEcRfJNiOzb/G1d4x
ji9InP4rxSAyL//ACLeyGBMV3STMatgccMlCAnc0jWckh/oNqzCH8/8jYXEHAmyM
DBqRz2hHSzup7KgBmpZrAdptvQwgPXUdZiubLQHY+0x3XuKrQlTQVH/1igpHUZ+s
h5EzQcjzhie0wYfIcvUg2lz8mvOsF3dzzRgqel7pAAFkWqsIzcba3BphuhuZft0N
1WPvT9rYyEqVN2iUNMivchYXxuRcKlvygnwEHuYU2606rrhoClvvKq2UNlunB0rk
fnPdjfPJQgcbwhZaMzN8Tl/lJzTc/FN4BRAiHZrvHzZjRDl9RZuGFrY/gKdGHsXd
sLjafwi7dT+fFztxOw5wOP9uQIB9YE0zFRdfkTi5V3AyUw7USFxwxYoz4VOz1mFL
pBMAcofBZ0X/0SetOTMh1/GBoAIoXxy0U4SS/vLnlrJdyt1WCs5MRcW4jX3h67v2
BB+8mR6hHMo657R3+jUwra+Pk7GMx5IKSOpUpz8P3A7TyqgRcDoAQCdJR2CP6yqq
l1uijEO0cW5FyQbZ1GK52sCEhCq+yxhvgnEPJfij3Mcg8B70dC9pGdb19UVJH8f6
bMkmAZrh7/4DN3M7aS9lW7VLG3sINrrdKsVSDDkKx5Wz1FkmmfEN04TDpoV06sSv
qxu3ErJXq55MTjk9bXXZR8vWtX8GJt/FZW7Gk32NV/Es7eFnP0y+p8b01XU3fPfc
a7AjWNLO+uVoMkr4vSi7ZlTBEvDgTrf+Whp2WnWlADOaXP0xXDKnYPv8QM+jYtdU
vbb7Wuhzma7Z/KyvlOqTl+drB7Glqwf/mhonmwYe+YPmHLt+To0qYieQ6a9x9kb4
Iil5amzyjAzaq8FUkiFrsk5Iber2ssW2lkys5ljl7OzXUoOB0/BmUroIiKmoIZrc
jZtWd3nMUzhbASmSd/aAkVgQksGPbN7XLasEnEqG4NZu9BX58tvG+WOCNLUotJCb
Jk+X/Ks+ye9xcIro3QFTH2BPahYZIzgLzr9HCx/y3ZrBuZzjNdEMGppPvs4TV+xU
9XjNk4/zYMRA3infhbWrhkpNR5RBQ5peOw/tQZZgRWpeAdXLsagsyp7CrLcLZBTl
QtOhAtdLQSDco/3t9tb2z6pUKAKXZPrfecOnmaC0sL59Pw9TfRkjj55bFo26MNdp
5Rq2B6f3qHB4ZID+u/KnC5q3Grm/GbSgl3bG44xucDUor7VbD9LxaLBYZUljWtH0
MbHJlfUJhaDVADqfqnhWX1wVQ/+8awPIeCO8pXJEmlv+uyZhiLcGXSzP+jsMKChp
IpWBafdS1K+M1og9T7IMzi5ZDYF0xPnMcqx/Co6SQxo4bVyAYlQNVRl+E3XUcKrA
UsXZ6AbUkaziI2U4vv+EMBc+8+19a+fjZosy06t2K5Xa/R9PHw1DYdyaIs90tymG
QTcFplcAC+Zb8lO3Fkz1W6BjwT2dmVMK4G7v97xNXRbveaWN5HAQMi86BRFPQwb1
Md0aU9JGiuJU2MH2+Ekj+CXvX9LPxlKTGX6gcAgy5GWYVt2mxDfX2a1Gdz13Xdqg
8ZhoBMvLLXI4jxRsu01oK3W/lM0nBaCml4R0GCedeo4yh2BzPLarX21woVhyx4Fa
1Sk2PYV5z8SbxzQgjKY3mnSuwm+valDx0jvQBHU4ZDUKb/cXvvadFedinkPXG/dT
49p6vUiebxgWtGlMoOU6hHb77Lq0NU7u+CJ14qsJQGUPcW2MvppobXQoh2SIyItE
owZpGbIT2uLbT3OtRdGgFBZWuk7oIqcQMZ2wSkP95Gp6do+ctmF7K6ZlQrMZBab4
9oevn4qdS0qITy8xwIQwG63/k36ZwRRxEcgQG6Mx3XFnpQAnP/0RUKTFEMqYmuCG
7RsGJc+4nGHGz57hXYOJepjybiQ5V9J4eZZwGK/gliNLucKANwQwMgUUEAPcUED/
lpNVmvU3XvpjPKCg4YFFjK2vvl3ze2nmE1vkR3LYCjtDfLVeHHuIg99myVouo8L7
dfXtlS/1Q2wSQhUVydcTsmgGfPQOHH56PhxozAMopPJQAqrdujDN1dK8WcdWqVko
9DMAjYNWkbUkwYT3ALXMtL4Yfy2BlG8rdk9CRuG0RxT2XRaql0Ci1r2wn9gntF7Q
3bpvHcGt9s2TAlQNRUKKfpWiCiCWOoj8YCB7n4jYIXdq4SlRMVQZjjoeqTSuYV/h
vH7GLygR3RkH8dPlSOztCRozx8zcnBKwzh7QzUzLS6RCTrHdJ83xWOtoM7kOuuSz
G5auo5rDMZsupJx+4L1dWwQaPHjn5KnsArMqfdL2CpoH3LpE7I1pO8sLCUMAn/k7
uBrGF9KaayRg0JPQptFCWfJawX8lIOr2HrL7Ey2THtlz1SvQ2TKmZrWRTCa/TeKq
MTpGOkkxvedaRYkgth0epzzwaVpxEn3CH+lOY+lMjRVVRMAnOtlT5PK3TMeZXjwe
nrkzfg7d3RUYJ10SFSU1u62Dg4Z4zFq+Y4A30FR9Son122JmO61uZWHNJ+qaGVWQ
IaCP/j5yVx4Wg8+GtCE54LtrXuWKjE+/3FGKxP3Co6cA1OZFPjpkW/8L1cX//HkA
lFhqjru6zAakSJL40lQhphdiQEVRLTIa0VE9xz4VnudVGxJx1tiNxqtVMOBLzggj
2HX6ZnPbNKXZCrCRX3kwm6k0qgqt6Ra5BFwXEMRCF6Ur/ITjg6wpsztqU3m3GSpi
HAj3gPA94L0NPcSU9TJOskhdAi1+M4a2gvlYbPAlA3GnYXFFD+QHpbJQ0N6FhKNs
N8YF1CoY8NsuDPk3AuIYmwQp/DMEcf0XuAADZB7p+nQ2yUUR2//GlA8eZqIyp89p
FaqC8e74vRxRx7LqrjCzoMOyGIW4z102oIDqB/BepHmWNOaUg1Q8wBTlQ/qSZ69T
0EkVjf3Q14JIBFgEnD2poLs6j1OYCCr2im4rSGKOC2lBIF71jDpi7qS//BkhPcV7
Y8cGZI5VI4cA9PcrF6g603vVpoE993AUPtYSVNStvheZPfcuETvNf7xeDCl6I+Gk
zPDurDY+kkofWq5LNcEFH0+5GmU1N9YNtzvBVvKJcRmxGwbz5SsrcS+7tBJ7o5R0
jgbs6e32xZXPxb5jiILpZOfX6ooaKdH15Fdg5xuHNeJ3F1pESl4IJinIExt63G3a
n2pMw1vMPPdcrKPznes9Gp4eDEXPNv6n40leP5gxTyALn2srmxnNqkFg0RKoJDF6
2VsgZHfIekyc9rZbuDd+Ah15mTJ9m7O2lMVYXGBfMhOz2vJY8NmnBaL/SYSpPuJa
Jjab5yIL3Oo7sshQUFlBYK0HRhR4CtnzhKT6UAtIJIchSoet1uBUdATSDV9ztNss
JIVc06DD0PGpuqxrcCSXR0ef4nQWg4MaEVTtxNV6aKh5G26TwBtVCJWO7rJpdTQd
K0Tqd95/8jMwAGT5qRcqu2eDhPQf5AkXMwDsRswQdBkOsb2jUIpvSg+tiLxvcodQ
3btQ7wDp5bOF+/SB89VI2YWCK03rfYoFPq75RxTLKsMbvDJU9EOYfnmxHMkOtufJ
2AFtRLP8HsfHr2HG9BgG0mlW8KTRoTt8P/t1BiXVwB2swyId0c8vyxIOdAg/uk6N
kSpNzedE3yBfa02winaZsYN1uuZ5KZabag6qLvsxfx+TOpfXCEnptajjAoGBCb2P
KlLEUK+ELStRLMC0Aw7sHn3CiwoWZzMo2IQT5cdNsx2xiIRhs6fiiyj9OQOUAenS
9CLQvRxm/D+Cf4TSOdPWXf1vdf0kPiX/+0AzUp8RgqVHr6Sq2FBZt3jgI8gfjisd
S0Xbw84yY1PoRe0SmiXBMakBLWC3mGQCQvc0zvmSS2MqBKo8aZ8VUAPmJdsiqtnz
KSXZzwpBkairQDg9uYasDs51XjbxOqaVm4+P37vGUYaowRjLKDyM1clAYTnlLfaB
bFj392hlAosvSTm4YYR/LEzJU/0HhUIkrFkfIJ/uhqa6gDGnkB+vVfAsgE1XVHsQ
cUv58fAZ7k8PriO0Hey4nuiaCYjcKUrmTRdwutjEaQmmMXwJMRXBQUoGuyZ3kx90
vtP4ot6nJthD1Vu7ytYRmcnwaJ2tA+3YNP49MfpRZy/Etv2gzPKzbIGl9TMKugOW
20hX9zAdEHu55EVgD3FOZweIDayzv/Dy1Zz919f17OEla8QsfIuWJfSudx82AFeK
jKQJvRCuI8xkC2ppNTJd7ohPWtB9KKmz7lEXdh/xmXdL8bczwQaoX+WxqsA6vRBM
gqqE36L3knDgu2n13yMlgvOjtA6/TSLy4dgto/LUVe+lcUQEEitdqfV74O37MtC/
YTNDdCmsUw0ZefYsPedRQO66aLyGS/Z65DtlHN3NIQrY0uvRrBc9m4O/2DhVAGfB
18RZGuoFYiRDQdb1l88z0jvxe7/Gd9INaWlAie6Xym1Kj4v1nosLZxS2lgnkZLsE
llYdeH2UFuTaweKmJRs1+CDNVj1x2MYfQ3Kh10kjy7wEn7HmqzRSxdb67dbVCJUd
RcDVanj6TXTld2u8TIXvvXHHeKhKJJcS78cIXFxdDwneHGO7Ypp8iUjB8kl8pVbK
wASvYYlQo61ryKQLZIUglhXbtCwZKcFoazFvWIYfunRR5P++3N7oNsqoiz+ocg+8
bFGEvaIig0VHdB6MuxqzYSpZ6mBpRZnNKS5bayA0rQrEJNYxGEevkke8vPwOXVPh
iXdn7yESDuIfwamx3ni7WTzemUy2fHiPziEFYCtzwDv7Eon4hcxxyhFn3oixAR7Q
qIsgPSkjxH5XqKw0aanpZ/n3h5Gd4A8MVFVo+xL4WMngUVZsPUtO7hTh5v0N00mt
RDnQ9FeMLhPBRTQfpIoqnZsQoUJZQcvvQKNUS5cAg7JxOpU4ETm5Z15/X48JOd/L
lw6AXm61Hxft0BLTBsJmeI+tAm/Ii5F9dMHenfAv+kKjGHAxy57MHQd0Q7qg1pkV
D6lSQcS8M3YKmj7Cd28lTVEXfH/FH4ksfG2eNK+1hMu6r2np4KV2ys+krb+I9jf5
erwrOkRaWTon6c4YhZMx9v+PPTJHWXBXwrKnjAW4Fr8HZtjTEXxIhqjOcxXqJzuk
YhcmWtOPIZ7VH+k9TYNF6mk05d+5tlurjhS7HKxbM8wEO/7mtkKQCt4K45ypaMd9
27pcgQzUOtRVjX5i2EwZAw+gOVJuOA5gSfjTO8liEp3g3UegqCZORUBP+2R7mA/O
CchCQyhB2iPgOJ1VgX1mjsYl0WtfJivk6pD1wNgcG6y3afQAgojKqys6fCWAN8ew
0RKT96VFVQF76StQkdoiF7g59cCHmz5LTJ8il8Y4wpU7ytpg0ACHC2c5Y/zfWaVN
KbM2V/+XdnP3rXWprkyUTe2Pl9pzLrsktC4Igk4NObR0TtQWOffCMKpOdh9cXmtG
DCyxdbyTsZikngiC4icyxol+Hp/WkzxtQd1iaK247Q62n2sY7e6W29q0iqAIr3Th
V1Aue1nFj1shCfaVVMRmqYqBIUjk8sR6NY5Rbk076Q1M6Ih/Xnn5yXxM7hVe3xhi
MQTF2z6yZOR3wna6D6IcXjefglhfpfepicxXVhu9xNJI3I51QcXCKzkY6EbvXqKj
REuP11zoYJcU+fAiV5vE+bPeTl/XY8MTYlmZUJ5nBzoA8CBVihgg27x2dGkcRJ1A
5s+K3AUDm59lUMC4nADrfyuyHL/OKrJsbL89DznFfCRGdM+jogRquMIQCfufWMAj
VUb4X+DHwKtc4MPsRJxwo16iUpmnmCNXUVXT8ZsndczxYvZ2OqgGyUR9pRIQBwrL
fLoRSVdDGnQmXtUw2z0cAi+1HbtLyQCV/3tr6CpgDw3xIcu7b/wSFvcV7vc4rMCj
bG53vODF/jl6dU90bIa0/i/fEiR0BlG4AfY34aYFXJ9uEy1haUZx6pQXV/fxQ5C7
vffgcIPuot8qxcwkSS0pGoqk74N0dbcRFFmwtP9VSUSirLELBibk3mZKwkiFdxOO
8qJcWZAOMM7KaVTDWvwGpGiiJ6I62LMrUdae+B5IXIUerIVjTT0vaQM/gunrMw8t
85hTmqZetbYjzYMvZQvl1AcCDnn1YXrcdDsA4theEpgtOZ3nyiStO5FJdcDsYSA9
giqSSvPaAMvfQ47kKwLIoOcApl2KBcB5x3Zi6GZ+X6RaZKHNF2XvIQu8TohXSx6P
yGjCwXkC+0gwOxMOnl7rqnYZayOu+c/vqAwSM7cHU6vCbs8XpmJQBRRx5+AKn9Wx
lFaPjIVXzO6lWwFt9xQpX8brnpKZPPMwrQ/SzRPqhwQyX1OaJ3YW0H261HTg0J7Y
YcDsT0hjbkJDgwd2BC/+klN+53FvdyGeYzAD4qJJ7QwxBwgXFf6fGDXFiTiQFWNW
hLB4m8dNOcNvCvE5x+o1//5hp9aeL/EP7YIovvOYa1hF0/lL1eYsn+s3LuSxmY6L
NulTGWVjo+tS8B0bUWs7oHIAdUa5sPF2hUIuSCi7mRpl+6L89fQAvDmEbrAX4gWI
w/zGZLtqERkX07YfbqzKo8vvR+ta7cU39PECOsOw5m6Kmg8KQt8akfqoljfLQMHH
G+gYE9H2zqm9L2CCIkPZLQa2kiPUIWFf10FzDNcBGsVzhAGNOBc8LgqSYUMwWXSA
KPCZ1Qc6ekSZb8Z13aPd8F3t0AAr0RPXzPt0kgSiQh14aFX+Sguir1IF4aonrlf+
KjheoB2ZQhAhCDqyDu0YKs4/aT0P2FHmKv91Rdp1gbitMRzbHrDgb4sX4fKjHsHT
+hXSPpsCb12Yagiq2TpuusIW07YUyN7MK/oPYZCyeDakfq7Px4KKLh0egiwk8ql2
zyRH5mF11Z8vwuRUY+E+lCBaeyN1sPQy/zBmjy6wBAQ6YJvDciHi2PejuOSri0Fg
rFUHYEz5i5qnmPXOD3q43u/fsLZQzbou7VY9OZpU+yVQowqA6smjP4T5DCTrKLI4
F2f7WhrDq8qhLknpEGhERnjklaIYrGG6h1xWZd5hCSCW8P7IAT8YLRbCS8AITgn7
JhnwmazHR+4tiF+u5co0p6+rPskIVkOCQkYfHJhjAjURsOZtj5rVFMyxjHbj9bui
T/G4IDjKQ/ccZK9Gb7+4yve6+51aztQitLI+WWMQY3vixN8THVOIDquAG2q0wQRc
ki9TdurebYOrW3TBnUR+mzmsBHJsDgliKrAfXPwWLcZE/IHGdL0h9DzNJ9b7AaXN
5hZ/vpS/GNTQb8mowfe1sVn04FSUu6VZzKYzZoVyBKxEsUl14L1MM/WX9Febku8n
nnwboAmclSimi+6eYpMR5jygavD4KoUgVZ3kMrGjXqEHFNvIw/55id41ICyan/pV
mMfqI9egMoC+OXi9RsPc9jquaEdnwr7GAIt2VHr5BgCK9PIV60PS+AiRvLPqlwdl
jeCq4QuudnhOTnr/ZXjx+Af03QHRjPkKS0OLTFrmHpUWks38TOdQFeFJoc6TT+PW
7r49xpOjYm84ON8dIqGpG9UprKj0c4vFBnPAMMJkuxaDqmmD6SB2G4toa5r2qnMD
eKLn7kD49b33tzssrzsKP47PZgR3qZMDzw9dMSEepiX1RKiDxPBJZl57zS+cIpHg
EXGSmvJPEl5bfOnNApThz1JNwcFvun/8XEBYd5HGdlSOGtsiIIVr4wLkCjoymsCJ
U34nOrStEf1yXNEmjN+HnNnUoCjIBxzqVmaoPv1u/+6drxgU9wmd7wMAS2RqlljA
qbIENXf66hk1CJXtjPcprBdRnhDpkJL7vWwlDTKbST+Kd0JFl5zWwTSLswYX8sNE
RNEwISDHCp7xNPuE50sub9/z4Z7ozWpc+mKqfkIS6bhBFTyoObXA12jfjPpAOh/l
8FgxnHDUzocdGEN51D8J50ozxgvvH7wF72h3ewPULx8eqS3LG+ESa9n3dUI++9Tr
RHCXZOujHTUGI0Cf1QD2dbsgAW0O8aEWRmSUDptSI6oqkXhrV9YlDOgh872vyZx7
J8ujKLWBnl86+9qV6TtBVt6utr32PFAv2wWvuqfXuLDt2xCBk1maZxnC5qZ5T6Zi
Ol8tZPq5RQQPpkprz6rW1MLemNZm48WU8SEq5neMyYAS5AIn6v8Nm5yAP7aiVT+H
VUox1gnysTcFgFHSXkq6PRYjjtxsXDBkTaBSoFXG96nI1sCo3lGjZMSWXCqkcYv/
xxOzwvZGBvZI7guJ08vosFhffoeTZXY2myazpCDxFh+rsi+SwVmd9IPVygB1e8qn
7Q0bzI8Vm0bQpD3uPpRyC7/OBZrMRJ0cYOkKEGWKK87t0gIit5UaUW4OZu2nM8nx
1ufkhwJtbAgprK/xYBuqlJSaAs4AVChzVl471YAoC4morC4OFaAxfbV7xwN2WPhp
9Y8Xem2Ke9SE1OPvtl/ncXP4PyJDNs2qNCiPGGIovNoYLB8IwjqdvjgYq46QY2I+
Fs4hjli1qS8GG14/mekhUY9BePNa8sj512HPHzQ4UhCBBkNsZR/ZFFAof+5P/A4c
n39Td0900f/p4/3Dk9Dtzb3vWvPFc39dhPa2PFukhFm1mKdbx32vTO3m9Sh6N+V0
jP9TZiwoyLeGyr1hkmBDc0GGbuAnusw2Hdw2/125PN4qUJyG9nklY9mbximWutKs
ADjsvrurRP+I7gde2P9jt8MYVd3AySICs/6VxAFvu5pl88SGo0BGm3VZi9Y/3549
WAe4cNnjx/sLLbp3thr932/LJBTpFn41PRu2P7mEyho5mFIuu57dKtyLNI+OrJNz
A5zBmWVdqySAbTm4EKguCPnUbjhJNrV6rlr9FQusGYZ6Qcftl44IzrYVUhdV1p8l
1nai/bCGDTnwlIfnBG6HAPrCn4sPRY5raVhhhdM+QxvOBVanSCnsfji8YeaxQOPv
ctWiyCa7HjfnCNLqAOUHZ8lOsJii3Kridkr8irZ+Q4qTU0ZX0flUJQFl2Q2c70pv
aWAlET1ofXJuzPFy4z1X+ZNC3zncdHF5gGDemi2QvsK/8xJS9u8vCijBt3jO2HWf
rzsQDYq2L9y31wfAlpVSySKTX+voqysNbbm1xoU8i9g276oK2+9ucBah3KHbTCk3
IlSV7xRy04uiTLN7I42MUUhf4sERonlqF+ppoXAvAO4kxHNvAaMqqSCX+L+ocXqv
+1YFRvf/TxhnrVUzO5TkV3sWuogDfRc0eXPV+X1azBg/L0StHDWGNrWrk5oXApPz
XwqSujXg1F8QIw5dD6h+UOzUXWoDOUahuJCmHtBdHSOjUMyCFkYGXVAhH/0ZDWXm
f0CXdoYYZm461WbSNxEVHxIRyVnvE3kX5MzUcGJaEGg6/32Q4piVnJb77ZchigWL
5+CJakS/2/N7s3PvjNAOFCEI7us3uDDHe27qe1CCRQRMXyFxjkC8mQ+CaJ+71p7X
DovBGzbHA7SWeaRurpBhRj836hUQwAJCVNWtNxwtqhBNj4EJ48HACz8ksE4SEqBK
4TKzLMpgSyoJgiSwPU+bMSNh7S0Y23ynCSFxwuo4e0cO6X1JOK+Z84M9p9k4Kr3r
gBiq4YKGXf2JV1s1xJU9FVZt2thIekgY0hNoCrPl3F84DIeTGtqdSm7gdV1868zF
N3e2j0VAl77NKn4nme3rjwItJ0Eg2VPB/U41svZ21ClJ/0XS0ur3OK+ii5Bn+ZSN
ctRd/qEwpkA6J8Nt0TNvl4szS+d6ljbUygKZFu1Qiu+g8TRsjRL4/bS52+tAsBDr
vedqch4WTungGI3WEoKZq3kpv+tSA2f2f6a8pn76AUZS+/Rz7Cbn5GHUauGbfiKl
A0jTjA5xrpv15RqU3vN1C99vL6JBTWfipalEDBrjwc8lzy9lmKfxpEM2QbWmVIjx
mHRZ9uHe5nx27rBGWqysVbwroeu9SUJH0Uvqy5kSQ9Q62ZKYI8G/vvTDg/PhfZbg
S/jNwn9eG2auD3rNgGu0nBbHKzCSQD5Qx6poC0yYvRFNjNLBjVxMEFxMvXBvKO7u
5JFNRTSphozW5vukAxfVqslg6dmW/gNB698DSdoTMw95dVZF8dlzYXCsKLzpovfx
dTheCUT+it41iYoWM/Vt4sTrdcXlrBzjUidmT3uZNaxMC0/KagxlqYpyh1azXPoM
TNEFmdY1Cz6nODTUH11u4/E+36WwPrWgCb9cEt37cYQIhd+XOrSJn5zPxlgrIbPM
XvLGMgtEOlIX6qc0yCWyFpAtS4RjvoXlIU3jWjF55WnMj0LcVqqGt6H5O1rhRTm/
6q4QmB6jK+W3xcha0g+6L7Nw61Wu0oBPdUfp5X+3CYAq5wm/XdKDQjV+nSrQcHmm
iTev863OSnvjnjtlvVREAIvLaiUDcnaD15plvXCjb9EEkiLbPF/FZg9yQFosgRUJ
yK+OHC69MJwzlEus+hEPYWoGGw3T0ozPtyE0ki4hVTmavCeqbZDNBFWcFkVG2ySd
jG6xQdC6pwnNKIHKYmbrWKI9peeH2dH6A88D3v4Sm+yo+bM9eZ6Sh3VPnVX4VklY
3TEK8kwdh4/U7HFd7ne1+XriNDY1ma4tiFfWAJK5whKnON0Kqc48dNSGaZuf3J+k
hLncrUrcvnRVEvE1pZhSIWWRSkK+ci/QpoTj3LYR4FStTAI7hoBtMkrYmtlyFlL6
Yq/qw6c612oS7kXG/BIuhaXsZgbxaJssjBy2N6z2QE6BxuvE/DKakqSFlxvWiVKn
NIe/5/oE4EgIN4NfqIeuNZwWNUCpIa/Rnfy1VcQzzW7pxU54n0n6v6uL3PDmIkjL
aBta+MAtlYjGdF5dPYp/QFQLWAfmy99/NQIbcRVkw9eNQj+xW41YfzYyPefQZ/w4
iJOwa13gY4eipYOuuCCmO7j8mU3lY33IwblALHT9QIPnxk4Rmkj2wBvPSwj30pg2
/iXrw46bg8PdftyXFfhBKSc8A0jyjt9+X3gqH5KgxAZb0qRkhPHPwIw801Pk74LO
KJuV7WZlmGI4vS8Z2doZwzGU76QUQ7w8W/FaueYc9OVIPG4HDcEUEZlJTS++Vnmx
0qH0vp3Ekav0hjlf4EJicXihbTX0vMTp7yOyesuWqccr4bnWSWq/v05Dh/FvGg9A
CZ76cNhPH2+g30O0sZzGNsWKzaDnKzxrHb+cDof5ao6EVswBMSW90OKMyefK7MB0
3JTYzBgXGnizPvq2+NxxVTK4aKpRtzy4CF60GAvsJmUYNpw5M2S9P/RoMrdFhs9e
0JA7AzVf42Wy3revNdndC8atVgk/CVsRTMi1dExJg2HhIFLQ0HTOSWB/t6VOL7Qn
7zeUstWyoimitrKwUtr7y8Kjxlb1fgmaIdPra0vyDOyyqRjUPVisQyoL2qoCfbb3
inK7hUxDfAWfSOMmGb35ag6txPBq7nUH32nzV3yoxeY/bWFaNqQSDZ79KqJxqQpz
HKUD8rr8yqbBbFtPityKfM3yEtQjaRBrDNfn02TQqTB/7WZ7c78fdGsXlFbJsmEF
t+T4OfySvvwcy38eLXwok5PB7vw53QosbxBC2SFJo+cWw737SPQrgqIrEaOWHBUi
rFJKyNx8Ktm/WLv62TcfuL4kpRclSA0ot+kpTTy75XFbjbHXG0V2ZBQFjjV0r4wz
q+0OokuI8bfwNyw/OQHu/tzbpBLMEQ3qGrHFRL27Vknbv4963SVdOkFuoRpzuvqm
Xk0A7hBhmHe2ZYIBh7oWrh62iG+OWS+RGZDOtoD9MnsGvML/cYQZwGokDo4IGca3
7uJsSFY0wl3/1ttFNfmbleYx4AhDrk5loEmR/CkE27nDOvEFDuiOvH6GOlxqsYnJ
NeTYmGH14VZsCzJYmYcrJMKLFCcSsLyV1gJuD2jrzSFW5XirIhu+G04FFGXZffVP
HE5E4Ye4H5pkg4H8+6MHrHMZrTrR86FgGqOCqZAafw+8GXoBGepcB0Dj+fVjKq8y
uq8umTsKrhziTsOP+VE67QV2DiedV3VtCTe/WBKjX3WkJI9g2jv/DyouBmmWdnDa
XdGH6W/AUT4TmQgm0m6ZuM0oJi+tNhLdHzRd+JdivqD3EjGuWpLHZ42iHb/e6gM8
zchCHvtLTQzqrjMevneIauAeL9H+utg2BY+ALQQw1udozVtYSmGLmm2Odxbb1VzK
GftpyT0BprYNxySZUckEN7HDe+QAUAfWrex+aYpggg4j8J78ztoiilHPht40sWt3
KAYh/3uFTWxN0zwXYNmig239oNRVyA3O5k//+gtxcCsvML4Dn+BASj3K2MxAidTS
3RKd3Vrl3cZ8VLAsFUDppyVA0mmIKjEAAWgo2C/00XA9QJhoPDGi4gpI8g92n+n1
mCqlrGRtRNut3ut9kZrDimMvxNTbLuEOuXxf+nhkpmPpkxuXDxXYcU1eWWK7LNfZ
g/YErihDLkwW3XMkX17cGKhOTqXcaozUFxyFODp6fYtk+LVtQrkbdm1ilKbdGxeQ
anw5UU3TVsAYkG6zGESk27cl57htZmyFPbKf2DLbcf4JSYIzzzGgXwISEJbPDlw7
DUxu0+ZmGMYZ16yzIvNnVJS/TQQPztW7Yfaxrb1oxG5m1DBiJIOB1k+GaKXNrSxl
Qo2DYkzWTrxTEmkbegEWfIJtNHvDW6kCPQKI/052yHN/lU2gbkqxujLUURgidhYw
J1TfRBLsIQM+vi3qQ7XvlmlsWv1dFauOXKYeaoHKEPoFAsT1LXAvyxqEIIeDCvzQ
bg6oY3vaOjCM/JQIYcKkpZG+D5hM84twwb3Bx8WLYasMeIr529MBNzMwBTNbXvZs
RMAGyR6WT9zyimkIHtgR260bMW82S4e4hlFCnSlaC55tkzYBmkpYlJ88/ZdRXBYw
uQKvTySYek5chXsyke8febqnW5avLrptkX+5Cz+kxlG4ShGmgqBhOPLWvHNOYNEx
0whk+YwgNx/34m+rViRXF2vz8hRVXvAGpiGGvGHUMvRc5aRj7Fn7ERRSaNMsUzir
ZCfyddewCsubdqRtqaRbfVZibexcBPPmBozbOK8EUzFIcS2fldnWyYO6/72purFe
mb83eOF5atVKwXVs6NsKc/l55zz3/DM3rd9FzXguCfKjiobKl621WPh/L0FnRQu9
koA4cY4+dAlrcAvas1Kol0viosJVofMwEIAZWWaeGEOuD9AOvlA2ubv4PYR3Gidb
I8gv7Qb56n2bYMycows71ACxl0gTeaacnddYtfJ2J9TTlL2YFeNR6rgnbZDCpN+W
1JpQqNRCJiTram6R8KAHzt9BJ9SYvlHGffA4esjW+CgCBujuEdT0QZL15bGYO7IC
yHC/kPSCepZ/g9A4pQL5Q84bgBmT09Mqe0BGikZgObTm9FWTWVDmIyXqiQwyAmb1
xhPGF5+o81X7DceCWhDJftLtbuG/KgmB46kDAmd5YUoWnGfptiYmCVp/AUBdyaxK
3MK2+ulKC+OQ/I9SnGF9GW7S5423dZsvR/Jnu1oQKXyNrjLo58wSXBp0+ouJSpDq
xQVFzP6w8JHW3znofSpy6YF/T6MxXDnaediRGzjg8KvgIonDsl9MJ5Tb3e1+aTNz
VbWqXyZPDPH5wOWixk8IxfNIdN/OjRK9yOl62TDluV0XL+LafVi2YglJ8o2ZJxHW
aVRcV+8E2bUwEbvzmVgKPJ8ghIBZH4BHkEHk18ogLhANq0h3kRgx+is1LQ95nDwK
L7ahUOS5lCAcjU/uzxCQ7ksTFCJcySzvXDsxrq2AmDd/ozSuuwYcPZjB9JzA2Fh2
obBYOrFNleBxazDKVWN1nhNiyDI5rjLc0+X0Xp+RkxQnpN1p1W5pHX1H7ZBI5jED
Yn/DpLRZjGg3f8+o02W9bVbIfFhv4AZPqz/egYNDAvlQpMVjm4PsGVBdhIDLtcV9
GuHYn9dKKVEbBU8IJCRNc+fKEgDl0fv4zzoCfo+ySWai2KUC74RTc5pnBLNK4m8z
T49l61ymYGq/A9L5ajAjIUttyAgcEsEsiD9UdUPfhz7JT8fi3Kxl9YFiCPs1e8nS
WamczOZjR8dDiYrfXPfEeA==
`pragma protect end_protected
