// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ly+b9B6ZKX7A8fsES//+6lLNJKN+yIQbeREatKQke6E+P+sMOJA9QK/jo/1Jjwn65l9Da69o7EsK
PMJ30NTpD3il4d9ArSsrISP4M9AzFg1GvJAzekZW6vRHOWqsC/XmTIfhfro0KCDuGHu/Z6ZoTOwZ
lfjvzosUEzDC/5/tZMSg3QdHEKb2ugaRY274xxkWhKjt0/Hhdj4AB/RZJuZHf2XIoamz81URhnqp
rklUjohtA5OUilNAVNVWBia+A6T0XneeUYXjdbnVX1UsdlBTFQA5NEyBmDFM2Ma4kBCRobzZ599N
xt2QACnRJdXhCshmyxpXUf6FYaKOG46gwzTEHw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5920)
xh1eGf5R5g7FKPgbYk1/c8BpdCI9rLbbT4ELKltUMmFCgNjU74hZjxaohlmcwdZ3C8AZ8X1bcmzh
lEJfrhFJhohv2+8oPOi5ojYNzdOJzzVMAC3j0xBje+b87r8I0IeBVstP6nevYGVuFnMJ86mDoii0
+eb8eEqVOPMkmomXBkpfPGewwJ+oQDp/VxB7WrZR2HudrZTReCGAECQ948IwF6cQrv09xOs6KxmA
VqayrpNrZXxCOqJtPznlqlrDE01ydR0opE74nwat9hPbNJwFTxfIaZwhWjdkJe74H2FaCkcJDm+K
CcR+RVaTHxth5mogTMCbzqaUZ9Nemnd268JgvtO0f7dQ3yKm4+NwdvY2HxmyJpSPHK2gwqX5pvPt
VQ4rZ0rs9PTW3fUOOVg2AgBvVOHh/sR5RIdi3NBhk08yyUzm2FkDkT7Oo2x2pEdelawVgUWq+Cte
CklhmtwMPuhzhSwIwQVSQEoUDqPro2grX3x22vr7rqOZNisMxAPZr7piYc6pnIY7sxEI3QlAboZs
uHjiGDmfZms2TGiqeGQQlUPF23psx+QN7dmAxfn/bVoev4feRNMK037aSLH0Cr0MVE19tylq5hhZ
a28gBVjpftv+cZDQpj54BiQQr2qkVMz7f4A0WY9NrXHba6G3zieyk0kxxt2FpFdtAhhsHlyleLH3
YQaUXcpRihIxPg/N6OxU9yqSa+qWAZfNIsm0S0G73UaWLpPEBcndb3BuMf/UDnQIfr73sx6lAG7k
v4ECV1Umre4gS8cZW+rPQ0nVowcsVCp4bZS8mTtilPEIuRFF3QdtXeEnUYInRqUh2RdlH2newbto
uuiJ3E9YF1m5ghF1HnocE6MIKHaszqRC9+8xzmz90PvJfpFgHkIGT0EBYh/War2En72kziyST2ry
E4gGg+OLfIAng29TF44AP9P3nsFZOChBA2LPr67/KCcErYMtx8jbvUqR0Ky/GDVktegya7MSFfFM
IkzNv5YZsT+Ujt48kWXPk/xkDz7Lz5MGhubFcuyPttZ2Vth8M0+0uA+ObER81UWMr+oWzgxswadB
yNrgYRJNnNtU6jxUPE1eHUKq/ERnaXUgtPdxgX6PAFH8Wr9Oh0xQQaAhAObGFKwpc13ZafuecON+
N8HNWEsZ9NjJziVldjtOEoa73dLjLzZXLLoE1LDn+oTTCc/RApNKYXpzmhNV9NmENR4MFg1SW1/W
qs6kgF1NR1vTTrAFWOdL2sGamw3IBoN2lUyoE6lKXsC4SsZFVQ5IL4LRI6lj5ayXHnjGgNgERo/K
gaCW4MzKNWGTJB4bLHtRz8z/zxMYuRVdwHCLiBpT7ELGgg3OeowRJ39t1nOqVn8oMjVqpo8lrqdI
WgRSLTrqOde6sj0zwk4Se4Dm3KUI6tjK3+xkwG6xFiyMMT6F/K/OaJ0o/xB+Cfrs1RlEambqpMUr
Dtx0ZZZqlIO5EvP40roJYCVHNNt6R++cdEiC5hGdRno1LoUy6Tt76DI6/wr/NGRM420tQAcdIV70
iT3umm0qK0CLh/K3ix0p9nsqxjLhMDVMDhnN90b6qHCKJV5n0NIZBDZU1nZ0jP959DkJbgGncDqa
RtXkFUyQB+yBy2yA8facnnk/aQ36zoZnPLJXSakD6fsRg6ptEDTnTO8ZjrAmB7BpT0xT87+Xn2j6
Xhwc9RtUQbrB7YfQzB6PeTLLDiX1xZ1DRRHfZEuYZxgp2a6bTwSiNiZxKINsgamRyTRDQY8IWXEX
xqrZ89BquttwkXkfk4P6FONtevihyorjHiXMUz/cD2tu3H8XnwRFAsrjeWWe9TyRTr4YIrJWvqmJ
PbWrFM/2NfVs5v6vIe1kai0nzXXAjTBimY+w2AEUuayIK1Ko6Hfv/ZPLwtlaCXR5CoA6JKIeokXT
hkwLWiN4itKkRpPQZC4CVgtKgLkcmGIfoo+KUjYU/6Ge4F9bomRd6DhMOhAI37pJ1xdZzBx0920R
x0KwEOgZJSF+RU1jKd7ITiRr2uGAIh5S8muSGpgHqHDjdHNQVLZxLVgTFL/+ixkfYYluPr+QIIwc
HUs2yiLp1HWaXzuTYZ02HUDtl9foO3kcT9rfyKcQ4nO2zVdOCjp2TNsTu+v/+o2FkogML1+7oInM
xhoTQIgDbsSweit+09jBSCxhaGZx4eo8+gct7Kn3/yuRBwjCfO4CgFUwqmQ48O1/iQPz+T11E2B/
rVl/FsEb1BAZvelOEgJZse5ZlFlaBB243RcuY02ThgKYCcigC4l5TYXbOiN+ZCWSMLH1cjugmBjH
xSf5ieGyMcL5xRp3igD9GQYApq112Lt3UHkg93wt/44xIoZiIUz/cYQlAQq9p2hTh/ORo6+yuDhK
LMGyGeqkQWLLkg4S4VgOgzOp7hDJXUdU1XKsfrgVwjQzav59hOtr+RX/TfFjmX5U2s5UaWFUGTpL
en9OLN0Yq0GixOAJwP9JBn4n8rqln50Pi/IG4HZrXq+7Uf13mLfjEt85zXLOJCAMst6Pt+cNE8Yr
22KBvOEILrv7FBa2qlAu0ojVopv+n+KjKVL5cESlOoviaYuPrEzTaBflRtCXTiswqxNUA4aC9gu6
jajIEN2CY2R7mamTESVvMmrf6Ch+p8fiv+3FUuTuqbFQ18H4jSjjZXu3LjS0Astdi8RqPquFqE8F
oOq5M3S9CJbrEw4zDqHRl01gxrdFjnqiaCnmKqdZ2Hirb43ygz+RlHP65SeX/z5nXOk8oKYMnS46
JLNNDqkeryu7l1XQJHGaPLxwJOIwMsQGAy7Z+6gzRB96ik2ySv8BpUeaqXOHE0JdMsdpV97BDYXk
AJ/7YTYKCqrSGfY1L6jO7zq4UGIniI9+vIZf95dZvXWPA9+HsOJXB/QPnYCSPgNRc+nUr2bNl2XM
LRIYUKR13rQz73E4l7xpjZj7RN6b49OPINOOHz7viSCVL+Yu534FidcKaiujsP0glzqYZv52xt7I
7nzdJ2FkDSTkgVwmLjeKQJTXv/2WU0W+H7nsimuM/PpUnYb+C6i1dmZWHjOjIOW1Zt4u9uaRhPHh
h0WJh8+onH+ggC+dqlBrOMg6KMwMOFM5Hz6zflM7I6vdoaxYl4Dwq+FetbzS9URpsRFzGw9lH+xu
bYjthPyuSVM8PWF/Un4fkF5TUu//TSHTCVlRUI1EBcX67NtBZgQ5804Z6SsU5IBMGDERi6wiH6Yb
M34mPfPISXpGIByXiIbfvBihSJgau9QovPZ5WIdkpKDzGayddLlODpyBrbu1P0NsxyDmlzCObTJt
uy3iNp6/BVJEcMcceA1I9u0IGf+vdzswP88t6Lj3cAZTZg3oouGF+Vtv9GSa/yvWWsFNg4qhpdId
3/FINhQC9MY5dOrQeJ1zdMF/WuMV5oQNEpmbIMLUd8v4jsxFQDmhfhswKfwFTbS+Cm/Nkten91mL
dgMeprbFLopVFdvyOqqFgxJR5pI2E5axNOXXRmnolLOu6y38elBqyYvop9kJEm136vuwkvu9mYq5
IoifZ4bJy6pFKGM/Um2tljQiaRPVRRKiKnb85dGseJLUL7bdXwEhuBWlJTtZ6JmBzIO2tXUNH4+S
rfxZ5XaSGl25mxJgBMVF6XmLQulpxJZwK4mxPGXGxFAWjwt4f++J2ZEublRe0Qh9o1GNQOzJUqeM
1gIRy0hL0z5BrEoWJpo3xyDiypnTdj6y/4sT4ga7VZbNLpF/II6+tHWrkaE13N8NEW/Q67/98nCr
EHdkqY8UeNsuSLk7SPMWNLS3EoEr5mAICx+V5+7AVfC94gsIq7uXil8RRm7t+8aMJzxKnvL8f3Vs
lXBIogotEedIHSH5NxW89Sh3uKZtMaopAK7ta/JaUPpsdXadqD372Fgrirn68Kb7MiIF1yPBEwC/
NKAXmV/XdSknHonc4rhQEg6VvgkJSkAuTxJGvysrpJvONbIO8DaTIgYPq007ETZL8cZGZ2V+G3lJ
jPD3qziQrrCzXB+XvHahfV6eQPmUu0jCUbyvPJUlfdwm7chG1ZPYn9nGBEnXNCr/r3VvqU3JdVOy
TCSzrfb9HPltYFr8Gs9wpHznY8lmUq2vgzu5+uNRDvUJF4lK0F9fDCEjVR0NXqO8YVk7huAAbMyt
udrCP3URFnp5EVBYM8OKlE5t9CkBiDsWcdRsGtXLH/LbgVQ7YQvhV0lRDr2PIjtRgry76Y26C2wX
wW51gpMHrah8VG34wYEW4UeJjdw6GHkUWH58jBQhKlZyMjgF4jsan/sMuYbxh4Q5pmcF0fkfNe6D
FZXERr9CLyJJnk0TVEv13T9ueUW9RQELJrnYhe/KzTfmGwe+1JW+kssZUUQtrzrIOpz44v1VFIbu
R53kReRA2ocad5QpM0VOphoyKr32K07vcRabMQp5Nilur778YGooB/KAUUvpsABIz4DxisTRArMg
v7BqL2lBOAKWn9HKUGAFIBnsYGRuf8/VxsL888EYK0O8DLwyv/eMlrTYrFkPH59MbR1ggkD9AnGS
oUZfWtvW0WEW164Rtst6yu66vfbDzt51mL/cZXigi2ZzN/ND91jAJU+JJTGBhKl/zJvwltVIS7j3
NoqhI/rgOR1XleZ6dvJ8UwfNQpPyWUm1xIal/7B4TbO97tVhzRYF2RBClyF3TNlLfRaqRsj529KT
6i6sldehVfNOezDn5Z2zGMYdg6xRPwkk7DXyI+Bww6yGHqxADLoKOdxli2fA1w7dQKlUw8b8bid7
eHbCAkzUnTWZChrQLuPSjK/3dI7Uh0vpKm7vleeSdg2YNt7zsVFEANwYkEJqzkFLNGpdvh0DoOCz
naDi22uER7uKHzZOPbUINIOk928iULAX1zVKb2vJv/NHn/wKjyTt1ZueBkJNyt9T1EPyWjL5c2fI
IgnyHk9Xp9wSnwSwT/i2T5Ljw9/wkjdTz59JdOAkOG9T7pw1uwgcP0GN4/n5LRHRgixzV/LGEMgH
y7yvJg7NluPewYI1MeXQr9M19oejnWSf8zmPzSQ78kONJPrq4PVZR28xbP/D8UE8dG8fZQ7yCNTk
SiZnSXERxJOcRoY7E/qpNxN27jJEAQkajbQgAIj1P5D+sT8C44gZmx4V61oesXhpOvlDa8ripQHo
GaGrU1ohLP8h5CHVyOcLbyRxX4JKzAcg4JaNVgNpRaGjCl3g+TeMkokJ+VpSc/IuEJ3W4Fu9+tJo
mn8PZlP+iZfKrswfHMZIAh98ee2Mw35OJ3ZcrOY/RTWe6o+5UHrIas33T0SY3LWcSAY+s6jJPTE2
Rm2Cwc4QyDJY4Ba+u1U0M+pXT5ZqiOTeVnCzhiE144J65fcTe5Jh6FlSHOs/G78t9H2mck/541so
jE6KmKsLxw57Ygqkx1vaKEBltway74zTeXTVYUkZTMGXrGaOYHhCDlJpikarvtPyskFoHD4AER05
180MLPuInLlWTsHMkklfLeX2ipEZZAOarT4OGCrXx5qquH/zMXTTkacY2IguY1+vthBNLSxIU+OD
5FF3LhncUlniX95WRYdc9TEEzymKYqwe08XgCUgwXFtLL/hyFuIRQ5lfBWnx8aJo70Hmt6DhCmoF
JWSJjiSqEVJsgYZYGxWSgAzehCiVjCwX1ekhw58PofzDQibvJE+O1T5KIEFT2PbG8jq9+kvNCuQX
XSxkcnYodfARE9+19lqxYnH1S9TKHEbBEjeE6NKosxXwrjTE4eIfFFFSnyl+mvFYUE+CPVRrRwsr
LWjzFw/jfSTCr9jLfbvc1XCAvPCPmR7fSAVNyThQPbfD9DBvVJzbmrI63y31rqtW8lxymvvAMEXz
LcUh1uCk/yDX3N4lDmbmIrPtyUWGklL/l/0vyg58BVtTj8fcTHcD1Yf5rONcEuhYWMbDb1s7opFz
a8mEqAQQ5NSQDklV2/BEThPc9HQMH7eqBNwVGiOqjih5IroB8zaO5aaO/LTI1nzsVEsQGmju65fk
rq7CGLVemdDIzL/kdbLRQoWtcvPWjmQShzWi9B54FFXyMWfvg6jeMM81+7XSG4xMrjQBxDOHWSee
11xMHP1I1itsMtQXmG5BePKgWQIxwMcnhzLIJK4DM+7RNyp38YGEOXVeeh38re42u6C5MIryAIYx
dCmj4Ji28ESIrXaL87vqCLjWOwUpSLO/EzLnVWX1B82I2lnrQ0t4fsKzmk8/XNOKSwx/1hZBuEqx
Gzaj9GHDNauGrTzHDDL2izp0U3WwHzRDeb1ws00R5CMlxREOgsF4MIiJ/r4wo+lMueSsTkgO3w9m
ho570EqYKDzQX6hdtue4WS+ksuBQrgGkIc6dZIpwdrXiNSYk3fIwWPk65JTDsYjfsCWZ+JH1ZDX3
VsHSVmPyKMqAEgco1nx72q2rW4DHZE7hIsao7MaLLKSwi6iT3sB2VBOVuemYFmztRUu+KOvPZkLn
uplJWNR08nSAcKBPV0TeyDx8912A+OrbifHm15C0X+YuyNAYLk5U/7yabVjNiK9UiD9Cml1VpDB2
KzkRgaeLxRQu16TiXzLFiITkGNodSS+1rOLBUNtZZXXuh1bmUpNrm4SA19AbVyParOg3XJDq4XsE
i3YJRpSAembn+pQuO1FaFraa2bKOCp3XA2XNSomo+IIYWyNXtmSgVUbuMOYF1TYyPTPGssLX6R3t
v9MQRG9l3xkqsj25LTTMzo0KZjx4MDYvTIbn3azrB8hILj5cXB2PqGjbTt9kXlnfl9hO6QleTsSs
8j9YuZ9s7VIWOO8teGYu5O1o+leyc0h1v7BThFfZr3Ud8kXseh06w0aE3McdhRS5uVDkIQlU1yOR
QoijK75lYrugmw3f75QRjVXQhj6FPQ+EtOAViIOrIDUQ8ToBMkF38tD8PHULcHQs2Ck7RUicW8Q1
SwXk2GCJUC3mu3xhBiCDUNA+ktlh3q1NYm4qi57WJ7nkUc7wRrH1rsDB+vhQPDJoIc1YQCSEYac9
BP0HsyvGa7RWc20tGnTzctcCw7LgtLIaEFynFsQP2DmYvgJ2SfOGTYLDbe1NernZgQfmp7QihDhC
zK9ITibtXqPqgW+pCJDuHyBHIboyw1gNI02zhl1eK+ueNXmaoxGW7nl0NpFsrhef0E1u3pNqci3C
Q8V1N5l3gBiKQ/aFvzDlLgWxRKIwgEvlXkfgUsBTp5B43sehMKAGUDJF9PldeBman4+6bDQ4ZgsR
6SjDRBV/yO0BLvu7xGRzKu9WvX/uox4+pCm6doVlfNH8PId7eot6O/1XYEGIcOXjIdjGsayJcCBV
k/OVxWcTojBwM/b3T6WeJaPTZFFFqs/4jvHxMccQ82D5Zuwl3TpyUjgwwFnJHvjZ1RfhlrlMeOQX
2i1jJ2Im1zj//2jGj8EjCogtxSGyGsMd1sEvrvsoeFEXGDomL/dF3VtLRuIKGmGSb7KrdIbDW+gh
ThEUmnHzGfFS6YyumzBWqzmLxhNUPK0+P62wmz3oWe5E3qpHFMm0V/yssMrmfAAso1/YpenYfilt
ZBE9HPiu5A25Ym/Tu4JnXZj5fSmD/dpEVfoDVkpMpTsXXKRfCTy4ZXydiixU5DF7MtpMXZcip9cp
z/zDEnfsgWT4uZXUWo8HBn2WeeI2isWf+Lo8M+s94ulZ1PHi0lDf6uwrVrNIUvWNxr4cX+SF4FBb
4Wmbm0cyK4at0/oIbyv7vfie4VpQOE006o9aFMdOxR9rPfq8wcU0UVpJIujHmrwy8lDEk8C58d6X
qKdPt4GT+pfYA6qxrpSU6o+SpHgge9QlFnJ6dW4Oo8eOFTNbfxfIT6EvGa1eUx2ogOn5GKkGMNvK
5i4nN8Qw0MfaJ7GoxDjPsgVZu2v/f3iwfT8dRsJiL/fqqSKCKGpFsjTaL1dV9TVjkgyqd0i8ZlQe
zwRou/s63WmiXxXj4TRjt+giHsKuzudWL5TzF+RZZsl4p7cpUB09mGtD2xfVl2QgtQ==
`pragma protect end_protected
