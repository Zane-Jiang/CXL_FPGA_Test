// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
IPkLViaX3dRFrVudL4Jl6DKOPn+/Nv0/oMlVUtCxR3EwVr2NqCbBZYqjZ8rjGQTM
aW5NhN9x/y8nF+94enywFofE/gmgdW38bckml+SKI115bJSOcmIxMGWbXZDraKI1
aiTDKjBiYMj/SQ+UcnDAeSBgpqfQHk4bnDEegjLmn4U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10512 )
`pragma protect data_block
xye+aSmLM15g/agrq1Vj4G48eHsvVT41X4wc8bDQHywfcF9b/7nM6NKbnvVDgGoc
Uig6WeDyvUM69y7HPVVF5zjnZcPqgpM6DmPWN4XIL++EQ7A6qPLlWwAheHa42l8v
LGc5AeIndo/hGrp/5wQpArTe9Y2xRB3WTgutpqP/d1fiR73Vhr1hcIy0SRIOoA6w
rGeWNFDYeMCOK+zHC9+S0fArSRlGrGdE40ioxMRGkBwAkohQJEzrcuCDfUnUJGM9
r3XhyijJ7a40dfG50a8VjO37RLvSveMINmFa9Zqmu8viJqhPozC1XtOjCwMaoa1h
Dgk6ny2IHtaEJ77+WEZ6kSSSPRpWWKWIt8aQiD+CT/VXPjqryuu7Tm+zwFXATM0d
VPOyCiBWz/9ZfAG2SZNTHBIiTadhUXY/idMY/6N6WzEwq2l+5aEo3YppC/F3NnDf
y2a0J3rsuygQsDwXzAl5dZT/xAGjZngwmZB9KB9GKr1kaQoCQ8Sj5rd6zjldxITi
aG80KSLjcH+ASEJhWvv/xOpARKqvT/7Buf+DOPKEQEn14sObeZv6DI/ZMgYHqsYO
surSYc2KWznmxTPw101FRycboQARxiWUiINNFnC/1pHXsWLwupQQ0a852DjzM9sY
BEzmmoZquYu2uTnS4+Lej+mvB8EEB2z9aGkyMPNq0eiZde3bofbi3MWLpRDAJ5QU
OGfCgMrMnS+fq/UyCQGUQXOnntBEelda0NrUBI3IfDGu8KyD90zJpS9LfrPweAC+
m0xwh+Omv/gBJDXX/ja4W0/J5wqps0ll0+D6sZuQVjUnYdXmb+jmaro2qgcGGbTT
TJ6ZAEMPQaYJcM3UA4ufgxaS6UAuvSVCgYAcXDjAL1biZqpYl635DTn0WBUSqldV
X7oBkkfmlj2yTF+MWNitXJ/8S0/gZw0ZOHJU9mA8ShSuFmbdMl4wK7Wwd3EQ9kt4
URgsSdFC2CpT+rSSf7lKihEQFV66J8B5P1DRgiOivhicYCTeRPfC1cFA8Dm4I2ZJ
QYSgBHCbm3whtnbr2j7l/i69iAAu3povl2Iv3QGnl7n9PaeOJEQTp83e2KZlMCiG
utTTjvExurtr4dPrTX240R8CozNh+ypPHasen75E4E1PIklRJc6gWqnFLgXhuTQ1
J3HpWfeNMzWgIGAA1+KxaU48PVt/6QQ9xcjcrNCpiiMyiTiJnWtbjLKHlzumvMG+
Fc4mAO7D8DHZMC96lQfXO65m3RJXOv1sNT11zMjfO4dvaheIR288/ZyOT6suPoF1
RE3JOyKXx/FG6CdYNDt8Ifi8LPoNF700ZfA8TrY/E2nkCg/cqtWXyEUwi7hmeEvo
RitBrpOTok9THHYK3GSC0vA5xBIxUa4HXiczTrxTrBv/QIl7pr7KN9/ImqEEvYQ5
or0rfWClJSIlb4lyXdBh2FMwLIGeNPml82zN7q4PV+PByPJBeGj6t7unjfDnWnyu
ekQ+O2EeBnNYJ6MzPjhmeTXnUK9mV8baSariAkLAuxg4skX1SUmkzzbut2jRfjHK
yxJoS8SR/v8RP0uKBMcZfllqQ76xIGKIzQW4tQlx4pWJBjLeDbC/PGgWfkmmDATg
RWb24THTXHKrffHNSMJL4L8HwB529N4AhwU46Q+OwIZV1HE9wWLY8BRGRsRUM2/O
VYpawO/bLAIFRag7TKTzGW5eE9JczjjbutQA4b8IQy2SZ7nIzWyyK96+rlRnr6uP
gAX12t4LtH0pdAazY+XnhBePM8nrDCg4dRr5u2Uby3AzIAw+GJgds6Bu73QtwV21
Ogh/83gKK4nW9XiWeVPvpSKn2eevRbN9p8mE4qvMke26Dw2bwgNZyrxZN6uzZ6p5
O9o33FNmt1WZTw3Fzi90J8Mewb6/8gIKEMW033JVDaPTzHHPonwSJcoT/x0n7xqa
B64+i6qrqusOFEYpJaUomzbRHeQCJZa09TaukekI9fqbDW3i5UqPyoCeIadTlM5l
YhVUJSOiDbeklL7r7K0W5u/X+5q4Z1dHeS8SHGMY55cqOnnrbnK6ZiD/qax5CPZ8
PyMfcu4miscABIechiGquYRzh4PzJMXZQ9uuXLXe3DYwkwQfOaNwubDTHVYr7NH4
o0LqsEFvYAqzpHLYp9PIb6zWUOelkUTBobgQIS4H1lK6LQl0IAyvbsIcbtZQL/ce
xjJNZS3KvspP6j4GkaQwojP0Xe4N8gWdLC5dtTDWAfqcpwuXngN+2veJPXstMu+v
/Yu19dB102gyN0H0Gb6JGVs5MP82L1pH7cFDoMgKkbi6eQvac0Ee5T4g3fYpzblA
x8zSBf4mSu37G5eQmeTJCly3HXqd0lvMv/UJmdbH8ipPO1iknqjuqBispY9dAn6K
fY5D/syqwJ4TZdvZgxrYUAJuVFl2l6Ahq0mAs7n29pYrozNNsCu7DvsXdvJ0cwau
dD50D27m5nJpC79UAv0pRN/iXaJTk/XKCztk/ITxdPcWoBVMfMZtS1LVEEjIJx3i
i9UWHLl0USaZbKjcjOYD3EDJ9qvOjCYihNPAhPAiV7igqQiFd36jiyNmgXvZAnzD
MPNKZvn3zpTdOeJrE5UXRyenGrARz2fWLVyz4C0Ge6nJj0VCXCyK9axrVjLR29+K
WNQKOPUxCyAI+uVOaOfmEOOJv3yPfbLgmV8n+1dfecGOeTLjZu5NEeg11lyFblZr
aOtvBrhv2C6IGoZWyCpS0fMlCw6JRKHZeub3NgtfbPU0KNuMbfK1Q7s5KeCGao6g
erEowit1gRApRihYjPB3oNfftt7zFQuh6fYnUlXWh7W4Tc05+Ki2NYcM4lfWEKoh
FWxFQsuTiJALfObU9pw6NQqDAq01NPYNgvX5xR0TXWeLEWXgccVMF59j+xW3AUaG
n9FSQO7jj4p52YTEVkQKb6qqVLQTFkhap9ND2dchUyg6ZgYS11svx3DSq+zhuRAd
NjQFZuvKJXwHXv5I6dnANRyShVKphF2pL3m7ZB6fwQph+vh8zXtGNQe98eDLpIwh
OyTUwvMwVc6QVoY9q3NNVPcxGM2vgt/N13pDZkxPvnjdpwNoRvmMdMJQTbQLtle1
AExCS0RIkUqMhL8Wdd0BWicKkpmTP8/htxf5Ask5LVpTPC94B47/ApJqJxz5Kv6m
0w8SG3fMwxYVJaUONjRTLR7fIoAde4kRotB/Y6gzgrhdjA5D2Bj1cw/BHBZnTN7w
czu788uC2zNNffa1Q8mxDt7rSdmljt2xqeSeQdb0DspWKGvKJ1gNjVyEJynlHi8q
Ua1RXtHTIcW00qk6b1Ol2um4Hvghw4gn8v4cE7oRfSzyteA4isLBLHQwKGn0vV4h
rqiTZ7p2UrC8831WUdg107FlhRhnW2wMFtR/gDAHEW1wiIJIlTrEHj5+eKcEKd8H
XOvWTb14IPJq87FlRi/+vfwLeWFdD0/ELuPKBztvQDY4QipMHqsfv26HjDD/WBMZ
/QdaWen0mqX71jaYlDULRCp3U/aG5nm6edOfhmB33j2sFlsmZeboLIj/RmxkyCWP
QUajLy/Stx3auPKkx0NS+f0efDY5Uk/JubBC8FPt0+OKwsH6OQ/6NsmLohFg8SGx
LzF8whmUyazVRbs2P0+BKJFAsjgMiFGgUj0VuQ8W36391TRtk5J3CUtlh25oALwj
eBMKMlSNibxDRwMKc4POXc9eAezVZw7dqD3OG3n/Qp33re1sCpmfJGo0DGFdHLNf
bgTUiBxeLVwuijzWIclg+fPv/To4iBLaki0tS4WB5b6f3kwnLW7S3g0rqha092ws
o5bC2ALJRsHep3smKOZNY6RiwZFQbW6mTvN7LfR5EmoP/YFxfzq4igOUF9jUWlGs
Xggh5X8CaB3NvWxzbOgyd/su37RKH1jshPPcCNsuM5JnthkhbD39pOWeIE7njrLU
+3adsdj8iCmzXVetJ+hEPeaxhshSrgadZIleq+J8vzX70HoQG6ifMMKrIsKl34iI
d9Osoy5o82DD0fLdeQm/TYjTriNTRXLM/EN6VyrWp5vOYi8aUANW/Cw+/eXpp6Sc
M5+XpicqUcliVVpy5bLdkhIF5P1pRQTBxNJubV5S0LhXn5LtOHDwmqb1OcpWroX2
Is1nH06+P11FAl2/N1gp+AO2s/gv8daRAIsHWwUcI4WqqkBAs+1S2j1aNxEzXV/s
6p50/6V2h7KciC6s48IgI9QJHNqfBYwYuUzSbj+aAmvcYvemzHsGXLrhFEW1nHNL
dnjRemz6u0iN7DtBuiA/gjLQsuwROtpDWhpgTk31XfatD2oxlVmGsKQC5heSRvom
rWRK6TBc+vNifChWNYRroTQRKA+KQRMz9082ZJ3XN3x103ZuPGyTEnItD680O78/
69i54DEaTdrnt0uxeMjM2ERUZr6/Z3Pv+8w9L+2Y5TIWivdbkkMmp+ndFxm+YaLT
G7RLMClmu6nXU//dRLCtMw6nonZfRZS8qtazkroN3LJMl80qTH/fxjHjunx20D4+
wy2w53hHoSJZaz1tqJphu1OrOIpv4W7VGAcoTYYt8CO2lK7eQRvVsY6aeHDUBVSR
6+gdYF7cfAUAfidI4vCIIqUyjfSrlxnmBtDyymL9shv2utc62AUGJTQsM10NIu7M
WjMbZc382NiAqiBj8WCByB0t1rwbF0kCSUN/3VsouT6pjIuSOMecDSTPnZHqNvbK
AXFuoXZjKcKsnUJb7UfXMN3X3yG9/qCsWvgWmYLr5CsqI6jboC99OXL/lv9aoSEl
NK4aX2wSIzlHL32z7F+J95MJjqKJj4j8io/7CQrJFWzwfPka+q1xTnKzRQ5o1bRx
/3Ecj1I2BXu0b3683LGqrc/mox4zDdzGX2M38ChgeEqQcPPDx3eNZb3Ok8OUkriV
Nmse7e+m4QZSWHjtD8NPyV2l4RQqYx4igiFpnPKqbxK+ScUevL16IPkh28hIm2Zd
/UmpIVPGyUREXZPau7rOuFOBFByMGd6hNfwyHvJt2ZRuIg+g1VlCg1NTIChrY/Rc
QWW+VcWEAeBRne1IrfYby45c9SwDxhMh1UNQwZ3kCq6z9Sdhf2MiDe16MEbhxhME
IN5We7iFT5b4pshvpevqgQll7YxNRt3xyApayNgGoh7cjAvmAQ2BbaDAW/2OUiv5
HKqJzOwkDD+HZ3jDaezTHeZqbJa0MagMPxse+9qGU/TiaUHe7Salc1YkaLrzimBC
jUpLnwrqgPqnKHZVLjGO4udFDNuE/vcG9Ku9HVY+/0G66zzR4vRJMA1bfY2J0Efy
j3aIY+HMgoBdPWcuo4gJcCd2W12aDnPyoCCWU1pEEv3j7y2jO4Be3fl9TUvN62Yd
DRBLaXlBC30Mtx1m4ozT12cTPejRUv5MQ9d+0L863UVPSFGfty47I2rWbhETrIR1
h+QIkriMB/pk3rQBczHRpgwA9attptyoDk0sJ+BJ2DYM7F5O15IPLuEfxiGWzmK7
pyeQTaiVsfJxKJd+EGSM9EjV0u7sjKuyzb/mZ2V6QTtHiisvbpmRUx0dfWfCQY+j
oWaBQbPrF/+p8qYI36SgI1MPWP8vLbY1QW+4ysLC/c6ybELIPb9KxBDpJgc7y9Xe
2UMWoN9USQHQivp6DSCzYyQ5pMMBTCaFXjoVU4NBk4KJT0+JuzJgP0YNxkrFbJ00
zf64wYA3NpIFkfoHgG2DgjTv1ib9s3RYVttbW9/rVRA7tvUOVoxR8YegCB67oq1T
QG7Dv5rjqTwZmaxJz/VA7pAgE9VSgD0PZjxyUHTI07W3AvZ8VDdGaqICv2xklvQA
ZEnyEzgGThtPRKM5pjB1IgKE16ne3R5BFWbcy/otLGTpwNNqZA2cBbCuLZc5QFzt
jG2jrmQnwlSwsnKwSEcOFucZjOsJiGCD5Kmy6sJ0x9Bll7jSbX0wvybr1PZ6WXi8
gx8tUuTVqdODXAekrGPtOTAX9cAhYSMEF/i9M9HcLyQAtGFd7cYttJfisivDLkpE
fx475Yll/yHAud407UBrWcc36VzvWaOUGKd6bzuksFq9g8NxfSTj1GvkJmEVKNZD
twrL9IEUTiCQAUVGI7T9lnkS7bT3OOs0yCqqck9WfxDbHPVIX2EN/kqK0NqX+w5A
PmyJ18CDDlc52XB+0QPdQrAmjEmk+aDl6BlXbK/MBEQam2RAYT4gDF04g7HynStZ
egoND456DWqGoSu+PoXHRljPhNgCuFVUQHvmNMmQZcRNuynrkJRxxrKao01BALFk
SiQIH4chcGgiexl60z7038ZZcd+cLg1y7hd4SsN4MO5a/9iryxn3FUrY74HHmQSL
zD05+TqNlg66n2TCx5xa9d29QjJ5t6bpEdEiZo+ZsDBPdtkoJvzh4zqlBGaDrLyZ
MM0TkYFVhG8VJPj+C+j8iOL/d7JoZWj8GZJswppAva0gxU7of5CvtqxKQh4J7ocO
KNKFmDeZvsLP+srTtEPberNn/nIiHbuDgTSBRbr7tYRQkAnum29n0b2YfHvVXCsM
4CS6Gh0bliYsg9QXOSd5txBtbtnMpE9gkDKkW6aabda0v+BRWuvuurxBBpYCR/8Z
KR9obWwj1XdaLdcaegkyP1i2zykgheD3V+q1SZQfcd1S08hXhBmxudTCRAWzYTQZ
WJKj2TOyVqyhgtfTPbsnCVITGTC20QBCHtTjMY0ttcNZ24th8JB57rnMtANrg4Iu
cL70Jsvv3ZmuH5ab6/hkEHf5ZHRRzNagpLmoy+tjfavlLjApHwT1ZYPBOexL4J8G
nnxh5Gg50il+S5O1P6w6TfqbX/mySljberKC1cKDAKX1g0u//ecw04cpvHXEOPkt
64LkKgYMi72MVOgrKyCwy9ASJ+JvLk4/UJ/iqXWK0g+Bk66BdVKxtjhcYaDqgYHR
9dfhE+Jm7CJCqvgw/08rT2QP7xTM+51EpEPpiFFjaknFb1WpYUT1Bjks72hn6vDK
TaMqm9q3P3difFCVGSzW3PMSbk+08UiTjfeS+77u7hG8ZScKTQ0OTo3JmAAHNZvD
7riUcu3yJRpRybbANGKCWKWR2Zq0UxUmIUz84uzuY/mAXQ0v1aU6G/se9eJeClAq
chcUAjbynBhgGvRLeR/Q3TOnpJxXk7nD7+NMfExatqpl5tCVgXxZmkvlK3ZYwT2N
jkjOdkAbH2I307QY7qkK6sGbEFgMal9L62nncMl9r2UTEIAmqqhMb74+02Um1J4Z
NwLyv9HrRtMNT4laQHkYoWejebh8W9fn1wHkEfbJPnp6dvqaygsQ0T8LbP4TRdke
y0VdJY2+n30+5I/nq5SJcJ+U6695G1Dp0bc764jpW2tOQtLQUohLRVK6zCFn5pZA
eAucAaUTDXXLWXqIyUrJk2wYWzLwPvjN5ZVK4KWGVTrE0DZodWLk9x+ms1rANXzY
MN1hLaQMmQKzwPGxx53tK3oGajZmyTdIntez8H3M+SSUoAgw/fdExxhB2nVkAK1n
lPe86TuoL57mB/pFzoMrrp4Z03QEaNdD4+0JiYMxOJb5DNKEBekSgHqKoRujSsG+
HpE2z2N35JdwoGgK1Mf+m5WqYTLvxRp/qBP59ekkealAYVY3vNRy/AY3hXcSTHBg
XzPjoe5DlnmHyGSF7SQ+8jt7oYA4bfVuYYHoxcWwzpp5L2o/dwQCXpU4XQXuJpJ+
sUq8PGh48FvKM81MNoi5ySaiwaC7c0RFwAYIDRbwz2+Dx6PL5+564LQRnSsjatZF
8x2d6zkmyQYQ0yNU8xmShm/LIacJrjJ7SxNqvxYPVpKwE5Jz4OtQDOWjxoZmeDKK
ol0P58A99p7OOBZPEW5JGMxqEP/LQ5vdq22bWnK9NDHiZkDa+zcGW1bxdxa0o/aF
FN2EdshnY5mJRKRYCbH5Uw8nCgAefZv7/AnouJqB54yAPsGJT43hF32FUMdI3O29
HjuqGxXeDouwlSOdwA5zTcuDRSf73BooBaGe2uJiqDjqkFCx0crl2Nfnal2Fm4HH
EmiIxp5FSfW3fFZnQ06jHUUkexrZTtFUQjOUt6FDapYaeScZMI+5H4bB534HMh0A
KkAVd/nCxIfYq9PuDo4ZZWVzy8Klvi7Fnsaq7Bt4fb8T9dQd2cRakvISrq3RjIW2
FgFHtIUuq47quxAVobEJW9TG6KGfAfrti0cK2oCTwqtxTtFsM9vyzI3i8yZ/5tDa
V+z999izdQZKv/jqvxALfc+D87KkL0e9+7GM2WsjS+bDTPyYCPLNRPe+v0Btw1Uj
SG5RN29xGcQ2/za+sQNbZ9iOr21gsu7pQfier505PYkHvHtxrvgSNSsaaGA37VSX
Gyl1jIeafgb/4pt/up6l7Z3uB0E8NjWjTbjB/jKz/kdhEGo4zU6oCGP+SKCCtc8S
ox9x3KJxAxItrHH6Zs2YasgwFzjy0M0hwOH8M3a4yKTc0cW7Z4qgF535uhPiY+Y/
7H2pSWU2dRS1MGFv8ZGAoBNU8PNt2SuAoLBtAvU/s6tl8MaxcQkYMxUHijJ0Tbhi
Drai3TT77iKO4Fjnvn5GVLPt+Q7aW+NBIqcFtO2XM7nCQbH11vO5eQH2HSupbsOc
uidbB5C9w4OIG5+Bzu4JK7aHESBBEFGizK2X0SgzNNzDwMvpb1BOjPy6NqCTNl+Z
gr6S2tRA7VFuinABON0gpYaWzBs3F5Qp+SSgXU9pQMtpO1gpHc/JcWLYMYhL4Tpf
5XVe0dx4sRnwb+ZtajVSLWi8XZbsdqA8ToB7sJ3OXI7OAwOELt/ernjoZSq3I71m
46VysI/NNdxqDWLsRwXUj1sEiaC6f+YZ0CSpv4Mue+q6tzI2CwPSpi7DRte/X9LF
dEBvqTgfLjTavNwzTYD39Qq2dPd6BRwU8sZLt6XtpBgWF7VL0MhzArHFeY8KhC0K
IgwKdouhLx7DwZVwOo4DuJT1LBjpnB0yniIE612mSz575SgcDPhTqx8ZqFadvuve
nK9zb2vlpqqdGYM7UP7hkZj2ZpVXj10unttMpQp8l52ykm96mmwqC2bXXiEAz9P8
CBfw+wTwirJWmtxwwqQ371v4uGpR0bbpulhcH2yY/olrAekjUdREWRWiW0WM9npn
f8a/MJmhGLHRo4C9ssQy82L8W9Glg8bNJP32vTNQojRYMN3fQCrBsTxwOn5QnOxu
AkRv9KgKa6g4r2aF0Egy3a5nj6qZRWGHpB2nznte7wKqdw8f3i808JrztoX23jLn
j5FdTQJorNSlXwCmWv6/0lX03RYWlJVeugxQbxA5KX2DE/IqNlAd+56FNiDB5my/
0oJ5/gRP4hx3xoi79+TpufRCeE/O9CiMXpGbuVmc7tUs6CJr8OfKaycpabImM9UW
lSmQ62Cs4bhb1kfDYfpJv2BlVD4VGxD0hVydBY2zZN0dYHJaKUIdw/bLe+PZkZHc
RXS153CVN1YdiwQGJ1PoPX6A9UaZy8igarZuD4VaAhsRArOl31LOc/38jVLhuxYF
iBOYluANMRyaQkdBBfbbHmwnqrnfbXtfwyx/OdK1ALJxqL1m8g4V1WpnmAvW55jY
OdPyw7iLQ0sJnJvA9q12va21edneR2hC5EnXe/qBVwfWIkGc2r9s1YlER2YNniSO
UEXuQpiyfpdWv6J9+8WAzjaWk8TnycLNg2C41/JaaE4u1dDmfO5DU4xX2bGs/PLS
ECPWSmjHQ6L/tJeEB2xSXNROlOO3lfMmNNeC5bubSzq4q9AjrxWdY89oUUZ/WGYa
W2lMo9b3ntGtLQkj+zg2ut0t8BjmXspHzAFH5hUqrCBR6S3PZzdxrwxN37LAVQ3W
QHQ70iFI8MiZIHDAtR3zP8qVoUF8otphyDrHzGUYD43IdtHiSMqZvwOm1cTcm/Ha
hVLSrbGoAin3/tKfrhPhO7n65NL0hBBpUE98nfeaBnPYxg6Tm6k+d7JrlBA064mR
Mx1VIEsYtjFE1qD37B+gyUfd1pbidD80h6enAIEvRK1l0lZfVKKX/f8+FZ7cXyWU
fbLeQj7KbjNZH4N1VkCWhwiw3/WZ5MEaWBEkd8gsZVTLw3QtQc2vlm3faFESzGkc
AzU6n+kGYceUqmDmcn+0q5fEPhxBl8CPo5xwQMrujRS0fsJ7AoN3e68WDzJqKxnh
awrozgVS9QkZtsUkPWbddYW7M5weZonsVsaHKNDvZp8hSCImWW6nfbWtnIjmaCDm
DnOhcHhobHG6CfQp2ph54Ghs+/J/mF27LXtvTKtLzZgjotTg0VIQ9lAMPju6TLJc
KJDhjALhsfHzn4LYG6yzy/wUrrYrgjj+My4OQpCj45WVrxYmti8fb6nrcpTkng5/
O8uA5SzD9KjfujL1NHEnjUIdIydp3YoSQQW3oPXUDplL0K7aNFrpnKnJYxVNBtof
b1wSyXtBXX9XC5UnQMu78m4cNsI7mt1pjFAlA9vC9y1WSlGzrgpAfsjOJ6RGUoZj
trg9OXArRh76QN5F+1J/BuXdQYpQL9ZE5TNoBgYd80ziLfgps24hOtKzv4Qit3ij
ubks6TivL2jablTXIX1rybHZpof2zPD65jN0GuIypVqWni81zKNwENOSliWxa9n8
8z8cAJseypdLZ4ViYe32o9IlMK+1GRB203QTA34rj7e10p2VZCrx6oJkbxydFJuu
fuOdSHPzE12es/G7l5Ows76ywkQy5BcR0zM0SeH7VDjqgfCKK0WjcVvXxbktiE6N
9XVhCa9yjcTiLUrozXyrlAvMDRWWiXwgG3Ufyq/iP5XMT7fDBTUIues8SpmBMWL1
InrJcfqea8lWut3adI8cN9FfnAk1iCrhySajBdvYpPHEuZVb6qcx6+E8FJKFl3Bl
k1TLDJBKzP0tzL5nV0r7806QL7Y5mC0J1LcekRJni06hkcjwEK1SXPRcznQ/MMnL
a6dc3A0/26QYMZ4gIYzYDVbXG4mXpC9igrVC88CmQif+B6esdAjj9KTCcMGl9Dq8
FFKTXSaQulmqW4WFr/Z8hUTnp1/7zPPOrYDrWtZ5c7SgS2uMOeDMXjGzFxzdsLp0
cKHyfY3h63hxMtZAcJ5UvOKvlmoNRIgCWJIlh8zfIozDmMN6bKAG3OIcAyi/olPe
zkbQf2DERjzkMPUbOB5LWlBy6uM1RD9NZGLqfpYgOPwE8iwxk1lchzSJvm950Adb
YucACoXtqOHYsaMMFPjR9qXHk7Dl9+G59+zE8Pc/PT0sk+kDcCiYEDfcwM4kqiOt
LqbgT+mS3+HtBrDTjE/S9SaBAWTzQ02PoPtjWcQ8W6gs4QIu7JAiNgKfAY+Y7j9e
Fkcw0rQo+FuGyRSLIhTFgF7LqnIN9HIa/8+Um5J8RMYCBIxTJrObjK+06lIx2Wjd
0Ia/rP/UAzDuT2LYh8+dxNAWxeBj7jZk00yNUQoc7aG3Md+NwgAd06nv13ix5BrW
26svWUynVDgG1IBZYjk555lPMlENzqlvI0IyCid0xnO+ckSMiORCMSCgO5VRgXh0
LJ0Hp5x0sV4HZvqlBOfF3+8ZiFeOyDLZ7KK1xgRWS4e1ZPxTD1uDC4bGJO2DNV/G
uUN3sk6HQQ2eSmyXQE3LjNsiBmvyrf8/BTLVClq2bXIAZMCiOn+Ze4pJZUcJ/Mly
Xjki/7LDiX3gz4+os7QRcj1fZToIvSAaEp7M0LtAs6XYjc4UBr7/TTrvc53f/LOy
1bAqm6U8sTWo4E2zA8TyXI76zyPnf58FbhUaecreMoYPlrtv5i4SLiku0susmJsa
tQdqphDCtAGKhqELRWNuncXsJjHJql9rLlQ2Xo1sD1xxMzJhJQTrNIABaZjtQJxN
85ys73dSLBe42KmKamtTviX9JGXGSrY9tV3FpAY1yCl2VlhfH6r0YJt85zE7MriT
X5ei9bd1pAEDnRbyxWUZF4DHXoEOOMO77PFrpWO71pDlS09LRyj8q/UHg/UPKCNf
34/9lIiwfLROM00hGieqigCmJIwq90KOCV9SDjrWytNzwvbXBmK0y8Gq5Z/0j8po
4078dHcOxnv+VH1PiU4e5dQ5XmwHlSBpVTyugovJDpE1xrEqjm5mjjiMGgXuAsXv
RRSsAA/rAc68KJB67kxE+LBqapU7p6R4OuNXu7bezjFj/ZWwzjxAKJGE+uItxohB
yxz/9FHIDSGYt9TiIw6pIoiss9FXBiu1PB5MP8N7QMGmT76pE3OPJWMFOoe+67BG
zTUn4Lcdz1t1LgutnogvPn0QwMmMxM11tKVzG2Zfq3gN8xg5G146TOcW7aN3BiNK
tnOqwlQ0NmeeuU5DEmctVDdkno+bNJ+BlFHcYhwnBM84sFDm8ShtAyHxrX58H2Nv
lkjZm6uJRnIY6fUj+6uBNxhYP8mg2f4aJ8qAn+82D+6759wmJqYhVbeF2ImufdxO
H3HrMQDqgNYw80/cJVORQmY0wSM7J8hMWqknLTEk7hLu5vPwqDZnoiNIZOlV/Bh8
EI6ZBtNX/kMiNhYumWbiMANQexX/WwRO8pEsxc0HNdJCuHLkP4J5oQbyHwdRhp7H
XAR29z8qK25wcQJU4mB4Kp/+hFbTNwmncPl1C7MIZ1ijTfU9TsqHLLUxAz6Y5cwa
VjD07xBHU3AbRwgRpVdgx/Vi3fzf5wq17FZTQvBhqddwtemcJMoDxiBv7sXAomDI
rXAqrfH0yw9rLdfwvyV1KhopHYQ/7/iQ6hjnTeI4FjeeHEoPpVmy6154+l3AWNS3
7Huq8XhjR+mwQ6em5Wm3SxMHpiVCj1wiVB5JaLsHS5ZWOS4SyvoGC0q2hxd+xC2c
YgcK6WJ3D1QxHO39LXE5XRVm2cERpNVcyw45OxjEr0AX76pTH1ze+faYpO9JvtTE
rfrPnUJnvWW53CSgsxcGvThjNhh2QVNdbapdGd8d0YgJkZXh7u56Wh+DVKXRiZdv
h+e4u0WJ4fbKqljtGr4/swQOFMy+z3K9PmpuNrk2bje0ctwKtt0QZCnGaSJShoS0
NIIGiuMia+ShqccwuI1wU0i7mAq6W3v1X3p0mqd1Zr+rFQNcTqV6/BMcuSxYkT/D
+uxDLvQ4zl0v9Tf9UfjPUY/xjSPUl47nZ84uyAMspH6EimF94uDWDGaae+4UzKxf
/3jmPL4IbhTsGMIM3H7+iTz/fGZZ/JTD9KsHmZWkkxHyHJyRSRjmkjnlBdKAsR13
6v//M7sPRLwx8NlYCPUaBu0m6znWyECKU2vhvMReahaJOou1nw4qkpwApBLw00+E
2U4w2FzULKA3iD0m4o07RG3UL0IskQf0QJLv3WsZo3c+49tlvc5YBjEY77hYqqBz
Gr64fVxfIDKhMsIsS+s66UNdJbnR2c1q/XFLLB/bl8CpUVuSc8gxpz9BX8of3WfY
9/oK6to5yt+hQl0Q7/kVmwqoZwxxnpe+pMXUey6SNuBsch3io67VLq/Xqp/BXjWM
JxEaA62yIUta8u72IuFvzBRYxWG4FLi07MB7hudLSaB+9BfyQ3AlZ9RZgiTIPX5I
00e9P+4KPP+hs4hvWF1FmexzeRJLWusBsaeCMEzROURGtjTPFfBjdofFDIPOjUh1
vWKWdAv5JYJr4XmT8DaaIGfAGnprCIxSVKvH2mkYjvs8Nqx4TwU06kF9sU3iaClV
881+V9UWet6DaiF5tg8EfPTx1RSKf2gdi7bzwERK/6Yp+5SjbGl78lYLjwyvUmVY
N9ilEFAKA/bKz/m3mWFPXW6oNRnbACv+DjUbkSfddlfmib7r6gd6M+K+qww4rPZj
qhTfG4mhL7U/ArN/DZT6CMBqWXwISmg6d9r1vGn6SaqZks5Kcsfx4vpMQNav8rCU
DChCVaLcgvC+r68boBNydrwoMBxOYiWbm1BjPv+2vhi11Mq0XsKSY5bC6GczPpHH
vHBAsuWMHbboj0Id0XWTOGRYAn8CjcsdHvA9CYz/hbjh0c5c0V4RhF793sy7Sh8Z
unDzMxsyhm/7AEt4ZfzZ+taFoujvXb0HHHW/0Knx6Z2OV4Ge+Nq+EdtCpnU2UajO
0nMNbhdK0tbQ+35zlsl3Ydm9kQ95BxFa778tg9G9wyNtiyTLGBW4uP7lBdYEp2x3
iR1hzw9LQuIs0soG2dFUHcYB2hbHIBaX87x1UEtUzS2Bwhdv7HG5zXq22oulp65C

`pragma protect end_protected
