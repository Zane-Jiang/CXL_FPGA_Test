// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LyS5R2aMjO4GE8DYouZTOc2U9BPsugJT5dTdifY8igFaPnMZPeDLnhT262Hq1m2H
a6aolUa7318U/i8uHdqpM4fxnPb+otD5jsYYQChczVS0quXbxTATaZJpd91FFlc3
tmbIbnDPxT0AriqW25rNJfLCjHT3ciRfPn83WZggPdI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 93024 )
`pragma protect data_block
uL6tLV6K7eELJXCX0bSHKk24Ezn6YG2GKPKWZmD8uxgy4xXyDrnAkHm5OqhmHSiA
OFDEag0zK7dbFmty+QKUAMhYVm80xS+a93NfXYqQLkE8WBat019dXvmgh5xcELEo
Of41I7bTB3Av4x5rUqYNx5XGeFvNjjrCPHVF/RVMFTGu8mglddO9UB6/IDvW18mb
S/tfvylLCjqd+FZPmvz9DRhJdbJHmAbliVOeHI6UMK9yRu+xW8FEz78iloxsXDJ4
/EYwHH80CgTz34/gQsspsDbX0KPUv69GWrOcBVHP1mHxauR80QlTyqe6hnd3ZZWS
MxvxIVa5lPtDllvTdgy4I3Vq6y7xC02rSVvwHoy5EyIc+oJRP5jvSPl6GQspKMIX
utEPWCKaZZcwRpLVPYkYVeZ4N3My9zgjBSzwFNjRKFlWFLINLWKRPKcOvknv5vyG
7gK39Y4bTe1eLHLp3qBDnwzMTqlmi1OflivUSOKYt4YaTvHPauNbcvj+aC52jY93
o1rBfhi7mLn48EPLMIGStFcxVXfqlsMAPfIkfnqhPxNY4No5wY8QNKglqxqu9OvQ
NTp33eAAXd0oT7uHVNoAsQNqmqlZjE5AyYP1v7bJGYLlC4NnDrBcQXojwEQ2gieg
yR7OhW7tw+zIo72FZp+OacxumwOcSfUwDmscU57ejI/MJsAhzLbafEnnZfFZGzZP
0WSq8MQng69ZQPbvqAaYV//MWBmObf0XrFYiULMlJmyXe46sEar2QppDohQahPdn
3pcjcC8VjYtEi7nBZGYwbBFTtt6W19FG61vURwjrZk7rmDXK8yiFfuziTFdhq46q
N+k4sUcq3oD27pTsntFQhV1GcxkKJzVDPwZSDBUqqAxJcWE48INvENpc3I6fdEZZ
x/H2XWhHlXxxggddn1yjnLAOZ81gqkXDw3Ms8hQfbENFMTh0AjJRiT8lJdTHvKVn
MWxeBgHPGyp36GQCqfQp6RRAEMwfqNxs+tN3mXM4LBjXKjx86RjirIsjnNsDr5q/
lD8kyQabfBRLWhX+wNNOJbyPtASL1d0SozIAIIhplI75aGo+HVUrzU55xIS6M4TO
cVhBpJwvF3dL7mRpAc5paUhBtTWhbnsl8bGixIzEl3FhybqxPuIEyVINJmUqwDCF
m/NyqQIQI91jeWJ8qRVWg9KZVHmMpnnNi0Jt6hyxLqUVhoSWuGGiWRx4ewwRUxDL
vNoWfiy2P/fBP+egYh2/LUfqICxWH0dyYYeht5UHyJFcwmGYHCs5+oAhytSRUU/1
U4Jd5LQU5DPI+maAyoBAbbARCCa5E/mwsYcgq95nk6ciP2S+nvCktphGm/TQHy3c
cisM6rjVi/SDRhtgwytNX+c81cPt2Sfo3nX9Y7TfyjKfi6ewgNxklXaFzlX0yd+e
Xl/cUtOzsQ9e4bZufYX0/k7eNfw+YbaBBDYWp945BJ44P4it1hFROythGWNrk9jV
F62Ybn4Rhenfp4W6l9WkeStU8K3j41vP1vDXdkNY/WuJaU0HUMRERxTZyQO3Swa4
RI4+jyZ7LE763VtSQ78oM8ejoSctKGcQuU52gRO0Ik1hcxZN3pWoFd3IfsZSIsC8
lIaPqzGFhcwYk2SUpfIZRfI2t5t4pLCuyBlXivYIBdGqekW7/rdqO6nSUiQsu+CW
4Um0RtCn6XyHuSl84pgW2Gi930Yc9Ygvujp/bIMN5f9Xih4OqAfn/+e+HLm8Pch1
20qmwD3gvwtHD82XI74snQ8txW3TxmZq0fCYbvJmCKZNHKfNcDD8faY20TGGcJWt
6q18Nai3IcZ8X4F67MWQKzh31cdpzuPxjk/2pMVYjF/zncpC8+Pk+Xs8J1Kxsazj
w7H1u3k1bvGNPB9uDTGBkzL0YXfm/cC908+c8JQT++JWwFsqCoIkEGdKDsilVmLL
f/intpAAtMpffzSnpIqQDax33wO2wElPy9QBj4GbFNm5Gh2jYSlfFQMMxyW1X48U
zonchKBnNZJIeESWq6B39E+jqJ7/h1tDHi5dwoyjneSGlE0TcE20JqOU9TaB/rUq
LlS0gZdyc00hlZsf55z06zS3Gzg9InOe/OnLZ73msA7e27vGAJFGZn/sDvtOhpAv
KmkuDRyOZfXdcWj2mtkTipeVAmm67JdRk1ent50z6SXjMBJyZ2JC/KTR0SyubzjG
rRPVXmwqu44l3pVyfxwFEPcDJGBBchMsP8+khVqY8YLoliLu7x6OKqzXLXugheIt
AmKrhmsrBR0zT2YvDm3v9onf275bzTLVHHThl+/5gKYi1iw0YYhIYeY8+YUmaaq2
cwy43LuT0HgN7AL7K9V3u+FUE6rc0aNpnQm9ZqGPzDrTp3IlhnDogNH4+F4ugFNV
YYv/DB6RawnDO/P7a1x9c2hWr1gKsDUtI4bp2KL/ZcM1mjz0RDRUdE0vSm8vEVAD
f/v2tU/h5UFkhtIuoVedWjBaprs5R596ICleWeG8LiJddIPg1awyAqb5ltye9u4n
YZehraL3+aChLpMiqHWlD6VlnNj4+sSKkrCrVS7xw2fYi6X3QiJCMdJYskON1yjD
HDyhUDAN1DodkxhZPP0w9ChlAjJF5n+wiOvVjox+2qUmkOAAwt0PcXnZKuuQrWph
acfNZfd3Flk7W/jl9X0kdIy5zx8c+XjNblxJp8z0vRJKRYVb4W+NFpqySCtoYlEA
1Me3Rqm1MigQbRkOhHjZuKDmLbd6bGSp7vQTBwQEQL5PVlg8FKY33Qk11iEuR2x5
a6DlmeUPAq2IJoK5asLQrqhFz5oRc2dIZxsWQjity05Q+9aVSJNLesyjF37HePXw
cbhtnr6OCqNBTHOzyBIGpdDmNgM348JVAUQUhnyutr9G+GXkw/L218v7JdSLteAS
SKhWA6Dsv1qZpHu/VDRdVH8aE9LSz5zYfFCLvcN3vXsnQzCH5H15EDDAB7kpvGt1
gcX6i7a5RntCFAYOrfNTZZiwhEmPbqQo+FqtT/AvOmurt+e0VIILbWfx8GlZfuV+
/xJKqzadcW2JBWzSUUCaq/aO3bFHLNb8oqx+z3Ka0YDhSImwxbyRoPtPFK9nNAzI
+9bc3QXlXKLYKJ0iN7vhmPAYVhQujY8oyiXN3Mi3KtA2DFG0OHdxs+46+lKBZMWY
Fl92HgG2z62F/itFtO5T3HdKXlPdGikvyKl9Rl4snVvjGxLEsjVICJsFnA0Jgh/P
oWD5CPB3/xm7meOBOSjUdk4FGA+2QS0hkiUkOm7vIPGDG1fTzV3XjjPo2b7MZttV
SgdeQzrppSP0QskMInTR3i2lzJW6nHph13ZsTipXVNdLpY+RTjb9ez0P4ND/4l43
qpt296CZqM+lhOqwkArkQ/eQzvW9lr8kM+N9qo3XcEifa0AmBY5vTrWvQEWSk0n6
vqLgDA67ds28LW7XWHZvRS+yLOtghqYcBNQSxL2QVTgVPblbYwTOhPXG2Dnt1fl+
kItW+zccSqEVrNIVzlHJQpB8Bzu/CagDksRwExFJciFcD69eXvcN5/6NMeicgyLY
+fxHQayz2vGZvZ+40t+l/H2gM4mxQs4Ikz+Ozq+skWHxLWRo2jFopEj/0YwUhx/f
n741FTtIeU422jPYEYSVx6ivWByDqrnSk9wY5W3gMzTFGcybghThDiEMzuJtHNeB
JkhKbumtyXC0G1GXseDNuPO0MnzvA5eTzisU4xz3snmUW7ax04Y5QMZfUOUAT+Gw
raJBnftb62rR5rbFVutvwktPQLpFNIVVihRtVMGCbX3At5YSuZu62f/cILLaLmJu
TFqTxKGn/ZuTwySpgASPL1p5LDoOqTD1skbAzcccbMNuu0d0AvCWdUOZE7+4zP5Y
3rgSF5I2MKPBXUQMql68aiZcV/vliX+uqBq/MgAfAlvPY4AX/hP3rhwyXRJ/SsY6
gqeJ+lnIPSObdk7pp3kCkKL6+bi8dsm1+HO0MxoxHA4edsQjZTJqso07CT5he5+Z
fGIVL9zgQR76r1Y7OMFOpunwvUGLdK7+hWBNJEJUPjvRTZDtSv/7Lz6ZW364pJwQ
5JJXmcD0C1BYsFpEk7DWeor6OKOT+gQ9FNr04M1xLc+qXel/sljIvp3mkS2WCzxc
NOirjxRQcWQ7lOyNmJEsbtXkb5P3UA91PD8g9ohLVPiLsEpVXwj+u/BM2pHvCEJZ
+GwOemNWnkVVCb0gJMZK520TH2plrNgcwYCZWvxF7h3qYegTTzXQg/Itu6qf3iei
mh+hTa1c6p5nExVuPK0P2h9p0VCN9b80HXlkQWQYQzvBxqAmIRp0k75DJSxD6HDw
XKqqqApUFH6o6Zio+8vmSaRKFUUz89DbNONYK1bchD+ZKGd1C3bPnj9al/z6ejkT
XdzVEbgvI6FLoDqmdgLXqDNfc7n689AT6GchgDZ+pw/VtF5YlXDfWq8Idbo4KQjD
RYr8/VMl1kdJgdIWpR43rtcoW5B8ctkuEG/Zs8W8ApQMu2eUOCcQS/ODnnaeZfcn
jpvq+GaPe5muRdDapoT9gtZmpn5C6y3n6272OdPTOf5vCosDlXglXsrWTmwRmLzc
Te42RX6mGzN6doEhBp5g3HHBuOMmpMIBAtTSW4nhzqQVPG5uzFJyuxC3Ekb2tbE2
bSbUDaj8D8xTTFD2Jr0UdXjHip4CxzignjXQv+XGBxYNdAoBYd+bQf4WIiE32EIb
V3EI1Cux+bG/qBxiqDnTOLkIGKYrn1CHKgi74eyjgVXzohh7iRicGETh4gerUOJ6
RKfQ8ZcWmm+5GDx/yELm4/OtCTxa8m0NlD2PYcCTz/lXPLDOJHDLofUCW/JpLuor
/wW/iJVO8qGBPIq6JnnUoiu/iuK8s6c6HU9iEmfyuob/ROMePWXvjXVKlu3dpXLu
RPMd8UD0UJQcmP+SbOLY2KodTa8Mf1vcgUdvZ0arpNlvcZcgu2DtmbTxtrMWNQyu
FqeRt3ppOLPIsWIrCtPw8SIsBY4s9/b1kTdBDKClVG8o24Q7rNEoKWAgqIPFem8Y
jNUFSSK0kQYY+p83tlrt33veg2Cjtpz22XN+t+6ifsfieWOeviegStwLus84ulc1
7jH+X3O7ykL8H9nxkALw6bwGWDGrgq3kb2iyAJ1/IROdJRreHeWwl3ZdzOe3etk+
pDc5cifA8lSoy+04r4j2LRPUFOIyo8B26TDV7HwF9NpoPQPMmvRNhuVWbb1DjuGQ
BvzOI4IEggFlqlWNaPRn7Y0jiqg0Gbmjcc8KS+wvPBWnpq9uQrJsIGQbFElV1yp7
cAUdULdeEeb7zUpRdi8NnDfrArbC3wUAxZFsBq4E0O+bfzrm5lifQlzB4FrIfoeN
xqNgagpO6YHZ3JwbaYRt/ocM5Qirhf7Jw7fOBgqNnKyXU7iT/MrODZvuaauFpxnA
Wowt44VywRzFMNYbaNh44eSNWYjxGY0Gf74EZVbUKa+bUvEcxDy4l4Gr6MCjfhJG
k9qyyp0jHN8xlUeGyaHUlm01hr7I8BUtRnBP+RCyr3/FI8LtB5cHmSFlF6z539OC
0jBwVNvlpOxwT6wjGIeYbLf7rCnfMGc6dZLmKjbWixXkO+mNAU1Eo2tiCZWPE8O3
YJ/LfbX0xN98ehOYJ3i8B5j/xecSthLE+PBZBvsZGYqMivGIHL8xqAjNRihNJuqO
I69n2EBp4wMCb9VCA2he2oEAvPeJc3OARtpyg2QJgNmmY4JCnTFs0MQfybQleB65
Ga4kR8I2C9tZCqd4RiR4muA10Z19jHb4znXy3kXHEazwo96WtieQWEfPm71ZPt0I
cLj9GNx5rMCwIFeHHfo6xBlGcAkt7BWPc6bE3ibVbOP8vp7lxfRddYsiDa+IRJbr
UczNuYIAMa6aaqX1lWw9maUVVAj4Kna6BCrzIbNRDe5hhOiUCI/028fC7z+gA9yC
pUahHp2e0noAbwtr6evOJW6RonGbs9flS8ngrdFWxgd/gSCDTIW8MjqiV8025wPY
Ryel+PltLTu3FkphmCeeEmyvHcQqAtMMvsaRZ2MSei2Z8QOUWtEQLJwhxH+Oj9uf
uCesaKVZaNMvJAANCofq0mOWSir1D1gkROX2LV4wedgoQ/jgS4q1r+XdbxwBAJib
i2UdM8NcOwhzfXC8FHjvaGCC1v6wRtgDA+FZ+Xdkq+03cvkP2dMBnVuqTKwSYE7/
IF2alJm+E/mOQOyS4GEFaBG3B+FfRR3AOj4gDCpKtpBwztb4zmNF8QZlAR2HS7Un
VyKDOq7n65To+5KeHOPHd/ojZIBv4B/KVWtnHclywFlJRMQnqAnoZc8pA0EKlW7q
SbkJDGqUGLbW/NZdqU53+ZEXyeAG2XGotSMlDA+b2Gw3D+flDwXJQMfpbRI038Df
nC8D11yGquqQk/pfDgZX/9tkn9b5Z9Ys3pcJE5RtgxEhmamv5L7xHzAvuSaM6aHi
ZlpNeYqaLyz66nACn5fbv0tQuH24wgtkC56o2o6aP/qPRtfZPNUdfHcvttqxIu2X
VaQirbqGlhF/xblipr2xUvffabG44kKm75N1C0SQbtncOSHuNQr7RTyoEe8xrhBy
ptjJrKwd5llvcua2eZ4bO3MQhx8ixFhjr1lCBWKp00hxeJjLxKQbgjpyR1uksq8n
k9sqokEagBsU2/BF1f79j9bSdQIw9g8gZ92w0hmSsNl+c2+jQv9v5xvK07Nc4hg8
091r824dB5yltsZtYGmjS8Pywx4C3PQJFSVphCPjlfeHekESJGUp0vZGX5y4f330
O8CGhaOzeWL/t26IQxvhVhbg3KPM3xG2i+uxg6gns3XyyOVLsOkrZlbH+Xi+KpLu
vMp57mV3LktdHN8uNiuZuGKuQ/MSTLxtePk9ZTKfC4H26XeLxUw4Boh7QDAlf/bR
sPoxWSdS+2+IIL64r+8A4FBBzGZRgg/Sj2UhP2VgODsXY6hyA6uSHYFxVxUYk0nt
2n7/8ZcdnV09Q1utogQoZPyVegleeiErXOzho81OhjSZ4rP7NTxsIYcL3rWy7b82
vcL67mgCwwyIrRd/dm9V9JqwhfSiCl0beKYCZXzGiG1U5/g6S/OoBqcNEOQBGc40
tBegfu5+AmUyKvPYOz/HT8C2VJB13uA6Z79RSccCBP/jZ7iZY4i+99isXQCC+dCu
4RsDrsTCGZ3jWIf+TDD0uPkQDQN8qRdTlk2fWdh7oovW1TVKVdfkMibXKUNrqT2r
RWF4XQ3fR9yfZlx2wZnwfwpTeeH7UVhgRHxG2rxEekdYaF1vU+KdeaU1ZC5VKedU
oNw9/aAj2xtTwN+gNUj/jdcJD1IiFJDT2IdTYX95dH4DiuzemoGmFf38SqSspYis
MimAmAolrOYkN+RBxofdpAJ1sa4YSlvuPDKuRFrwZTjqcrcbQtTePsRU08NQvati
g8YZFno8ulrYlki/eeH23CfTGEvzr1Ij7Ov4iMF+TFVUJu+12bDxqGIN/WiC3Hks
UWO8SvEcbyoXAs5YlVEE8D3027IVGurp9fxFkJI0yVbcIJ84fHyTBzmMTTkQng5V
/omTxexlxm/2+eOn09Su5cvGDcygfg1ToWPk+cAXEXyFFrgMcExYowTr8xTYPLQF
aLUasyy5C7r/oNNnGOpRpFgVU6IY25opGygBzwVRoDjALRjrTkh2Yuk+f+VzAWzT
8NElQTozHS6sjoTZI6TZjcyejrFIIT11yzKcYBOGvBiZNO6sV5/RbSwlf9V+AS9p
i67UtXPeRUuVy5Ot4uhv25tphs80BpugpS+g5Z7SvvYxPlwb1xGja6Sum6dym5ZD
5KznqrkL3DiIAmzLEsJkWMhFOWMqj4/twZMyhL4mDkAH2iSAmj7hKuijgIs7G7MZ
FrUzMQAJHTD5yc7JDp1eBSUgISQSQ4owkXFOyM1inYY+FCDi5NczerR4UUIqNxOW
zDi6Mxrs+ZVj5R0cNZYAzcbR/Rbg5Y5+2LZ8leG+nYWBE/Sc8IImpiV96jS3s0Cj
ysJxFOxJtgzhixfCbJjwvlknSVQpI94CJ+5pAGmLa/W7MWDq4TN4OdcQD5a5qWr0
kHW6JsSrOO5tGEgPk6kEvOy0w7CS6Q8OgU7I5Lc2vSepArGReI28HmozjiE6S/QM
1QY07YQB1V2vWOusLcirM7pjJ3WNovS92I59Evzs+053ievwBnf5UbY6Q5tRSdvT
B8aQ7cS2u1nv232Dyhu1nHKhLWFljQTP4KgRa2pC/lrXtn75DotbLOcSDi3WRhZR
VOkBwVVtFJc2WWmFc81OcPGn47L9sxunpi2lh5jwaOQhm9SqPQKSb8U1CZyYNSf2
BacewkM+9jABompB++SHD9zY3i6wMWEB0S8UCT2vpLQGCjJVHYKgCq6BXV706o/9
kWIMs2XtjZ9gVA7tQ/0N8fkKAELLOktbO85H5TmAwcfntz4nBHC8GCwQ4yB7w+lZ
dZX2CreLmmLpcpwtkJX1ZvrJz7AGy0ERIkW7c4082G3NADNrQROavT8zoZw1ohJV
M0EdPzYoC1If8b9csNVyvoA/MjdRxLuZtrfibDdtNu0kdVoe59OPqupmomIWmnCb
OdC1ggtYyhemtVNw6eoIh9T5h1tmnS//Q76eLzCKjqPZSPhG9naRgRJoswZ8p9rt
lJxlER4jTBELR9zr6DRTrIScAehrdvVQssxzXHK0xmg36w3bb8OZjDgyx4UV3SY9
n+7hIs8KgUAkpY3+PtKKJdl/01Zvrti7soVZ7z/7Yfp9Vt9BVJBVR8mnFCfB/266
kDbPLZ4VI+JndZ/9yGxjOgZhQJgOZ+l32bsEoLDuqTxmb6HZGeIjkYTIJ29uM2z3
sH05WO762pbRAIj5TZXqULAJ4l4yfhjQYl9Yjw33kNxHxLyqTJpWNzAj3IY+ykF4
yPsIITvDgQimrjUauZOU5+4ze/rW6WbcYKKJC27xipNv4zsH8kMcRSqIL866omsf
CtjVsza4qT8uiJFoOD/csrBuUUKbiH5BfqMIfpqRwim6gHvI9SlRR/oa+e3kqdXv
b8RRUjJqwpxhbAn/4+P5/1dIaJpG8OIrjXwJZhoXeFaa7Ns419aSIe1v+OiZaNVa
t9gZNhS5dHv8+sxkVJe1KjkCr59JtkiBuLZbZXV8XCdegRC/VfbIk8njviGwtJYo
b9t8GQDAnIf2ngmXFZzuOmpeAgfT8ssT7a0RDX0KXQaPXciow2WC0qhK67/xvsTr
ArGBrqH6D3pOA4wJWWsFGKBMIuTiuyZA6ZVcvh8LfcTnlF3svM2JjiYXY0xTacCm
EbgK5xz8+2TpAZ2ek3YMkb4RMvfGHckZUtiWauXewvKQy/rQKtcKhT4d2yKXTv4k
oDWbl0qfxL73GDlWr9MIEe6jbSQjUDxw7r1FT1+gFwbge4kir3SYFKXWDmlWq741
9KSWGu1FuNAqe61Gcxc50HkeRoiKQjrgpjsbFnhGNqPlasVR8dFhBEdsQF88SQWB
s3bdjuXGneOv19xMK2GsjJVTLZKkawJNzrwaQPdX2Eqb4HrD7dbJ+UGLmz6bKFDq
qRzOaOQdqN6DGfWvbpYYFPGxv8Lj7LYOd1noMY9cFdZsJg1SY5a/bV6tg5HRwl6R
B9n69yRauQQUwpN6yV/5wFjJZljCWliQhE2qI1zFXO8Ql0Whoef4J0fusf7qBO9+
+5ncKsAdM3z5VJnnQa6HjkhlbmM/NPAdwz6H/pqZWC8M08YwjzEpUxg7I/jA8iDB
iFaOg3P6x8OWzQCPadj4vi5yKKHlHB5kPquml6IVGrAXkjmbaWUtYif9WtVTgi0n
4w0Ggeaeuk/51isaJFXbAtRQUKadzXHKHxV+HbQhEab+mK6vB/YBWBkUPtINWkI0
9Lv7awjdmIN2ZIcpsBfvNErJPuGUhe/8e9uzFt30TZcv7KARpXjZMzy0X6l3PPSx
WQiQcJAxUQ7hP1hQKgmzyP6gVepAKFNFq7AxHPnyq466nLjVaAnhr6Wb3b7Bsqdb
6hUTTXhq/+hIwbBDOvisHcRpVcnDqStXuwbBsdFLQmYTg97CWrF45RyzLfeekpVv
O9bjGkY7BNwjJS+JLyzEyLqHM7oWXk+2vaowzfTHtJ/liGK2NxVL+nE18zaKCV6M
TYbNURuo5aS5grM9TRArfLnvdshfFU1/ESSc/oDspvr+DfgeCiTJhBC7Ezm+uJKp
4DqGMjUbfQAOk6ArgRpukkOHLyu5NfyATy6CkDksDI2mGeW3mwIzYQg3NPtzUOVh
gct7zlVvmPQ1PN27Wcpm6oQpyxVBhAMh/t48cBK3OwSWNm3EJOxEqVVZIpdHfbF3
GZiiuRYGdbtTtpYgDAoeyELSpe5nQ+W1o9ScrvC3EUz1Miqvb7DzqRGg5BoMvnjF
p2ElbmneGP4xhkvXWE3w7WaO5h0uKdFmnL839/aEqWBv4Sa+kc1chQqMeFf9v0J0
8YMdhepc0QTXG1MKTm8Q/B5aQeqjTpIfAk9X7gFGKTbgSc1GARvwP1trdwJVMmE1
UWCTxDGNdsUvnxLDS1KBDYGGpdYAGRJZBv9qQpVoe14ggPNjvyCdisq2C/fesZBf
+5jYsG7Hnr0FLwyhOsxtPnQBxNLeQLNpkyWhuJusai/5Teafnt9d5nojRKG2Qwyp
lb0ti8e7a7oF0XOrrxBil76gTbJQfaQZ6r9R5DmerWiYmm9J1wmZpX5/NH8oGnsF
gV+8mVa1oI56htPX7N78NP3m6RHxs0MZ4jwo+aY9KgQPhAjWw/Yp0DyXGRRhWnzC
WI1CT3DCDYJtD0of2eKfYjUyp6cQIZCxpGFaSoCBHH0gI3cD9bnqkyuXQJlxargU
pDdJ2gIMepeGy3hhYUiAlV92mg8b70wLED4f2pmALh9LRKgTnqCq1FhCoXsGvrcR
CtFKBzcT3ki6s34V15oQEtN9RkIsIKs4vjdugaKTt8dRXlqJ1u7fUEbIpM/iUBXw
txBZQEiPHArFRajPpLo55D7BZVdb0N1aaNN/V9qaIGJEJL7h97TXtBNSFOb6i7T2
HIxHyuwQLvBoTgi7IEslrqnAT/Ckau0ZYrIje0GKPdlzeyjOaIYGqzjlT8G9njzg
BgTfyI0Ox63ymrqigQOyrSuJ4lZi5VqBiGOqoXBJ8imwDj5J0sP8sqhDazL4atEt
xdEghiobaQSiiqhExRl8aDTzAvliDstjFYI0O1TchNDSAlNP4M/97xpaQO9Tj+OS
OfUdv+ywIYSlfFCPLtpTczrUSXgD/5MUFYB3Qoe6aeHMmpNDR2jAa5OXPXegY7U7
vHV5Zq6c5VAWS8NfnbY040YGZ+ziE5gCJ4TOtpWpjveGkSo9x/AfiU94O/1rA05g
sG2t49SPxY837gIRInoAKmaEUc1jrmyb0eQlBhf81o7A8KN8r9TvMFvIiAFgCUSy
CvAnJJWdWpOg5V/DF269O9jclJHdzy2Iypg96m7qBqXa5HOqU2AgcdthKeA9/KOF
nJJbUd0T0AbdpVNkJOmTgc4MdJd/Lpqn0BiK944zGZCNT1YpVYlaZu+POGW8zCYq
O8Rad3zEY8EkeoM2O3npfF1ewy4/+G6ArFbD8OBwsirTcLVWsB6HvONzTnsP7oxY
IGXeb/NUnQqkCZr6OQW8/Zw1yLNTCET/WhBFUN9g97nmifUIGalgg3G/lFytZRXX
m8i/3m0Ztml4j7q5q88h8u3VxQupjKFjiwKaW2nZCmZ30Yof5wEkReqD3t5OYWQE
bB6mj9ngyhPbcmQ4dkfXo/nlrrxFWcukgrbWFoAyDViw5/0Lijt+7bMJc0TvALjH
4OCcb0XDQc0YWzzlSUjRcAh831cItDAc/eaov9M3jXMYN+Nrsg6TDWJ0o15OoC00
LMFmXAHtmJWbBwrcBbNXiRpMz5rxz1/AYCkMv6A0azIU4ngUxz9qYICB5aYOSyXj
lUlHUZvNG8VDnRjsb7CrVccM9nR80t+OTWGIs413BvSjGakZCbEId7eC7+gYrN2r
OfzcPu2aLkWToWNlsWlgjWQEnHH5HJeAaHr6ULEwXTehcumMzRbSxhIcKzE1hmMf
ndGujCowDcRy4V+/ndQjF/1Nj0Pwa1Ss1Csy3HKPUf4M1FL9IssVcuTircPVUTC/
EetF5imxnzqeUuYPv+pjlX7lcNyQPUCQVmWqgSJ7ttAwdinb+ObP7a08DT1jOqXP
5FLOzmWbwb6rICzDrgaFdqY/ZVCvL8U/0VWeYN2ZqGK3LHUVE4bmgRQZXjeo77L9
jumSwoVhNeMUMncpdRmaNF0SvXVd5Tq7SMAHXQHNQPhSt8tuW6jKATQ51qffCNwe
eAlYxiqZgsbM9d8tHDEGF4TkR1E3FkYGX5Q/3waxAn75svVJsvLGqqiiEPvEojLB
40w68Jp14QvU+emrRgxWEv8v4c41B4RyCJT7k5Jy/xvIYGNoJ3jKEvng88iFCD/o
9GaOepaJr5rtmIf30dRE3sei/E1dbE90rZ+ivKSicrJ5imtCbZcRgeUsKMiAACOr
eXHqIg5gW8cZVYLTLxmnMWozlWZ/UKiWXmUwKQhG7aOawdMrU7dnNgFVlGaPW0c7
bFpdvv0vJ6R5o3CERySyfQO8CTaOe7SkyncivvUi8mZBUmt2tqjHmzfOwZnltlAo
rgGQGy2VA87f34Y7dKXZ84myB64ujH1G4K3+arfPpYYNk6gWQB6VVdw4Q/KIDMIW
/CGdXEkTBytJupPp1jDgYKlnRXgJaMrKGnQu++AQ4fZIjZJrUoPA333czk1yPTPN
F53WVff7D+jH2D9nTNYP7f6CoqgL78TmsFoSY390PKGMvvVoL/YUgQPOCe/0tjwE
x6Txo5bmv91k9FTj//C0XtBfHQ00vSzM1vhn17R2YY3hfHCAFpbNgFXepkQnsIGH
bSIZ+mT+ElPPtPDG4pCzCLyaXACIoH0bA1SmqMi+GYDNmVnwNv/m9m21Z+GJd3a/
yWEQ4pQWsBj7xmUE3xCTNmFGu7frlPI9DE9sdvXGyh4kKNLUfUAb643O2yqna7Fr
CQAjcBHgwJx88jZ2h2YjUWbdMQOYV5SnrS3EVZhb9bypatHwmdf89Zz0imnmF14z
+0LxEyVArZik/E1HD/qPITdELqpWQqoYMkbEOeGHvuk/2PUhTBA1ISCEkAcfUKsC
7AG1J853oG5Tqgiy1wm8QlfKlkFTkNOk94A27gboBg7szpSywPXItzW6N922PXmc
i/uXD8SXeSlHAzcseG+deCIfJ3LOAO67vZzylNEN386+V7Ctc9IipQgLTH2dTHJF
UtjT05CM1lIwl2gkKh6Kw8rtsYhd46VlD/fhedhL+i5IG1YBULzYqCtnZ2x3NdYU
xAMLHn7Nnc9h6DSHDF3m7z7jkBZaty5SyP3JIc/mw+1OfudXuOtGO923vqmiwjAc
Pc7kkEs0FEWDIqv19bVtt0PWx7ogNVfdzrJbBJWkC6505Fb/EuLDFY3obwex3Mz9
NgDwEO4Fq4Cv5/O5L8QjCaFgcpgPa+spt/pA6w55lUbicWxMoA5ER0PaKaF9k8di
tQGkrJf+TKUp9nv2KI5Ljkyc8DZR0N62Ac4jsrnR4A2vuoj3Jg2/xYBYfc/Q4zJT
gmRUvQsmKRV809VoImZDvzkJ9hh9PbZu6jRHWkVNb54Vf+05Q2zsd4O6dZ2QlgWd
L0HMRIfV+mahzH6eLbrhg28gIZ7LdoysBNUSHxyqP4ViRmW2Hhc5wePJcwjXBnEm
XFgTkvBLmmbZBfRlhChxvxAPM6jrO3zXgFm9A+X+x4aIBwQXaZEOyWGvxesLaGSU
q4ppjPZtBjqHo4LYjArBXY0CMhr46lDe3WMIOkleQuQakE0vPcHY/NuqbCmjAUZF
VMCAPdRu0kJ/bCuNtvbngoOOM9fPDVB5UisdvwhvInYeNMwJOq3U5Xd/qL9vVAQu
iC8sCkZDC3gSOmWOgl6dgmsrPpOcOsvn9Cfo6I/MM5Zel3PvN+CQF1/jAhQ6AXq1
inV7Epb+ZI58nHCw4oeUzTOex/Vo6dWjGn+0F6FMieCU7yUhWLOp5x7l2HbQEBJn
oczXFEOHwBlvU59ZnOawSkvJpDFnCL4Mr1M5wezMPJb/GWyJXMqK+CD11OzMLfR8
iSl42mgD3ZSvUojhDxkKiPY8K5xTrxESxTc+sdNe6OA5aD8iNOy+WpjClExBur6w
H2GjEXV1W/K0D/ikWxbiamy9yLO2EzSLlh33+Gj1MHI8m+M+TAnH3ToiOXf1KEoQ
Ys2d9XDJ39X4oLC4YHeK2zb2gUxoj6WIalXR+FcUtKS9ch/pFOX5OAOAJro++rwn
BMfBmfjRJqkv0417j7dpCOoxGWZRf0qn+FxYO80GtGg+aPiRwhWg5F3SSvLOzAIf
TPlMU/WT03uGzWyLqNQoRFAub/dLWexJgvnzhdjgtEyBsW9lDaDWzvG2Krsns6rX
QvdfOHf2wyFdn3hQVU9u+KLGyuRrGKgRY2M1ID0C8/zjvKUj9/et4Px0sJQQ4hkh
uot0/IQX8Adv6JTPdz7XX0LNdFpnfwB/Y9p8JwQS8uZAlet1kkRtyZURXVUptKte
KNzP5I7nIj+GizIflA9jLpugBYMDo2JX0XUv3UTgXekd68SWg56RDPuX6udw5ctw
t5rIlQBGSXiXjWfyBk6F21tlGA0yauNNUwgns0qy41k2JmsdxsUCrnPi/FKDkyHu
tMJEkH/hAjm2S1OFJEU5oZGvM7XiUR3+15cnGfKoURYc1rIdRl36MontoyRJosS9
JCOyLW+uraEizoZTVHaFgUvw5JR6+yOXu0eOXaTZ546EeHVyBiHTHsXpeMb+p68W
QZSB0gzKelieNvR4bSwlp4T1oGmT1oclnWmBMyhj+rkhr2l+hWAgnm9fp1sn56Dh
p8jkh1ji4bdQ7W1z4embApMLA/IT3f1OfOuGiSQN/sn09ZHzDURV6O/xM39oQGyZ
QQi+ocgqz+vb0RceVQg4YQHQJrIu2RluMAstX58Oq23vrzIn55MTHuCerAOlpBIB
0FVS8kNbnPge4ph87Kr5V4iON7L5Ka4m6ua3/LYQNtGwLQp2v+aq+vfWLNf0gKbS
d4n+tWc/ReQjeA6Aej82Mgv/FlQWAkK20R0ylkaY4mPx94JUIldawgi3nD18ybfJ
avLT03TdAqPCEhChkQbQZTqZDQtSVzHpRHFlOwRSgthh5wijdxfEfM7gjrLJ8JyX
3uNqkzq/jRm1JAoh6wFAL8CeJ6t1gTVFjvrRNk0Mknhv0yBz3ZQ3RVeZR69Ywk3I
N1wr15vNQrIDfrifIfNoKcGNbr0Pyihu4QVSVkl+erwIPFfSE9QbUdOKBLJqb5+1
f9L5W4cO6DEwFbbywPTsKbpm0wr4JVNBKgflc5v5vAXsP0rdsxCDglV+GHZyjuh/
GLUVmjGeDXUJylk27QFXNkx4p53xisoz6Cyz0hPP1LaRrh3ZRAVw92rAK+V5kj35
/EgJPHrsxIlX4q7+gBdtgvlQ1Oz9Vj7qbX2srdig13TjVJN7wv2dy6c844/AyLGU
zsgzfPwmWGegFL27X9cR1Fi2cw7UpK/vkVOT3eXgOIjFSSaujgBIM/J35aEmBw7M
qexWNSHfFmkeX5IJ6IWoinJ5/Dt/KZIk7NDNniE8ukD4p+JOn7f59Q2m7w3iQg47
ghCB8QWY9g3uvQu1KfVhuKlNVN3ywbkIPBp0Co5yNURgtxSejDyTeI6d2JcAxaBS
VhCOSo0TwbKQmMtqLZTKuTco523Hpe6RGhza60cVGgrZTUpQwzqywUyeA9ehF4Vy
dyCFa3w1UO8YFmCBsG+0l5+mXmJnZVTKixXvOQ+Cs3eKy0wbaXZctf5Nx7TDBDJ1
847bArOaHT4dqNfAJsEwCAD7oHX+2QLXv/eDolaVJnC6sKasKWhoPCCPk82iJbwN
mIzkEjg72404U6j402dVSqRjKo+u8N2ElTr5Ak0J/JCEyUM8irs20Ux+1lG4qt+J
TE1y8FbvDWveEbQ0hmFbCPNxzlkFjNxNyvX7jJfS0gdMXBzOz2ARhONBoKt1dcTD
8ypkxnY1qmC/EuPhKNNyG2dZlRF/JxDGOWbuxiO23SbtcvmiRTZ645HMINPovAls
NWLvADFGj9UoDa1GIKz1ZcShz34RNIz+jcI6MBGA6dmeT9Utd5RhLEF4xyzq+NYO
FUYy+yojWF685LEEbXTxN34VjspwiINE+SUo4l+000b7OIJnfG/JLQ67LL7MuCAl
q6V/bsWoisn5CfsnOR4GGhhnkG9MdmbUUoMB1Ga6rHmUyvcbFH0SqeaGtop/5TE2
z/qWXIe07skq1EcaVQOmVmKctrqPqavC/G47VnN4faUzcVIS14qbgcgiO21X3Po1
SWPos09zS/+EaWSdqGpA+3pPDqOL5W963TnbIyxAaRbUNrstKyZ1UIYgdhwSJb9o
eiOYUPNgvHSkKPxNOGtHR5Ru0/u8Je81fWUvvgMssztFD6xLWf2pKU/VQXfMdb+G
ean+JLctO+eX180qKksJlGDoXHy38g896cZdjfrnLUZ/rWc06E6+AuvreydfTVUF
C+MkcirPufjede79sA0Yz6HG2UujV3XhbcA3P0+2+sRE3JI8lQEYDBV6tn8v5VBf
QgqZFKfyJdketlEfOsswYXuWrQYUz1Sytzl5lUpwDbKfUgU8KFA/jFkO6GEcdhzC
2tnIlM2mNC7VLLhx5aCO0ZIzkr/ZNWbUkWAngyaxdj7Cmjk0YkRnsBJHDaCRbAgP
vFQn6ylXsBLgPBtEQ60omHbAgm4LOXNoNg7WcsPqi2xu9RqH36Eo3qUO9lwDNw+1
auksUMwsrBYhvMseH0SDgdbWrJWRoLEgQYrtoM1okQEkcWdwa+sa2Dzau5aF9es4
IypaRivU3iqSbC5/dS1hbS0qZST2YfACjqQsVAjWhbUc8Hefnf/Qnvo+6MRS/bUT
Kkzhaa/zET07cUa/BZrGLaW/dzUQVH4ABwTJZJoQaCncKhbo0N6tNMXtbSOvW2uh
sBQNrV9PPt6DgJEXfJnoNhlKt5SLEsOS8nDRRhzCK3at19xG7/al0pOcrQ6KnAUf
mgV2Fv5gZAp9xorpwojShV7xqD6ErZPTWOxEVtIY2KF56PRK8yC4WF6/9PeRP/P3
K0VDhWvQXni9fdvewbtWvxh6pEaruqMKe7YOKu31Q6wXW3NUbbfN7kpouiEwCwvQ
tfHPJmbdI7PkEAfZ657b7FMWtgSj6eHh+3CCQFdaT+G646mbdPUxr3iRC+sSkda8
cIDz08RqOtXjTHW7YiIuyU4WLx3jcpvN9120QR1iD0O2wTOnjYa1RAaoWmryws/r
Qjt5Gnzwy7+Xhd/P+8d+hzfz6zmZbqweyjRlL9mqWxMg1dWvwhzFhQUPgO/lzx43
teLHVV11zSU+vdCirtyorAz+C7ej4+z54omH7XByHR+NwrCvbh4zZ/rg+mn4lOjx
gRKm85Wk1JXelrmlKyzkU/aZth8bazqgH4XfYYCwwrz0uwV/nxKe3IHnVx/5dXZA
rkvh/eRMh8o++50UuCIBxq6lS8l+F1CXLr/G3Nt/jenJ4aw9/xYph6o9rk7hPJF7
9PNlYcO+F7zp8TV8mPDC9nyCfLd19BYzunjr6vo2TuKnPejE9Lk/OfYw7XkatFzV
TALm7M7EGW0bF3eJdJeuYOwr9/RsF4q9tg/71lL/EsHGok/pEo9bQhSVqCZ48HGy
jO0EfQj12wk7RE29Ct/10fsPpuL1bC2Ry27T7ZnmVtL9IP9/aGLORsav30ZXvIDX
sEyjwxvw3i09FTeG+VcfKmi/9LdP9X/euAEQ/lkUxJ6ITQxo9JoWTJN+ooOV+ddt
PoT7I7CjA3jIvhX0gdy+fDUx4QWZugUsiB9+e3cEu2rTy8Vt3Kl48V65YB3+PUBP
t3Ame99I5JzTe50uetOYIve3GjDs0KJApJtMn0MHVOX+g5l7xwGhZ9vny2ReZpGY
IgfWIksBeVW3ovRSqEf46BQPRvIve6h7mxoBjdPhcBVEpsicYGEA1ykRMF0acaI3
bc56HRZOyTL/T/dgMOJFt2kjfKjSj5SayUhEesCcLLJzJnFunOje2ueMhTYdhy4B
N2aXmL5OjRucPMON+2lzLnIHYGB3b1YAWWpr+s5X8Ynkioq0JNYkQ/TYPYvui+U9
+ksm1Y4mkN2SAxBcD1AiJyNlizk2mWGCM13oTisb4B+9ra53m+wmRNENuCSdmR4C
D2U4bLRCY3XJATtg+KsQ4vvittV/yNjusbe1wmmy6sXQViDnMVcNQYuboo20mxxJ
/IUtY3iEcOAP86YGTsc9FKZUcNpOH2XhvDYfd2CLmx8TMbdvCqms0qx3T6NHv3B2
NtPfDw1rRlC2H1eZLLH9Ft6/mEC9G6GJvpbzhZHhTvom4KQPe48wYUC7xNMAgGFe
z8R61fyAy/KJbm2QAQh8Qu+HYhZNSrWiMgwr/VK3ua7MIJISyevsimviTlJGUQqX
m/xeo4J47hB5KWhJh/DldAXlmTXNmapBFihbqj69+GkNvz8Tm967qpDeSjoouEko
QjDV1XQmAGXyGVXicjzbGtyWdlnyV9/tz6JImYp5O1tmcFpmq6OrjLcwbPfYcYu/
KNnfziPg0SMzVRaj5gSZo57hg4L8p/lgbA8BieveDE+9t03o9AfUaf5QCVKCG6aI
15xKEE84eHwR8fUNjsGg0QronNEkSuze8msdgGr14hy+fBQDYVJbMB4KJHWSKXhe
0FX6W2Vh/MAdSjqpDGipVlQogmjCG/ZPIhlbNhnsW7PQltm/B8fbSO9mogg+m6f2
GwE2TxjxK3CDADdDxc+bULMOoiK/AbKVESptj/OgRFtmcR5U31MxI3IuqN5WGOpl
yiiXWR/cOYzz9BtHDm5pY2+AzPxWvPr6LZXm+faMyOxzZdokOgLMTDrWCJClKX7P
sweDs2fTRaYqofFx+cTvJD2yzMaNRqfptmRs3dgzT9ajVN0v0UZFkI2jxA9e3UvX
MUJ7Ui9Wrn+vBMCu0V6Gg+k4ISTrtAOtHLUH2sGAWeh1ndSY9L3rIeL2tRyZFBJc
a7uyWZ5A7GDUBGxpixdDvRTtrI/hHArG3zict/WNUaZbQr8Nm6MZclbzCtbfFOuY
UM1RH9Isq7ledczdOzR/CTNm3tZMDO+LpfFx4vT5iVZozinAco8TqZu8bsjIzeGO
nRcb5NtjGK2qXSBMqLHTFnCbeZwleYSBiBlCAWAB1GMUXXEOnemRCThIOM2mroRv
VIf34rDFcECx6HrxLOVypByzaH1SPwvk8pFuU66hjUXHYTzwRH5zbC8OqSFPA5p5
9AqAB+S1/QMDqG/XlEttbIFOkaNNLXIaC7+rHtFVbiUEgKanpnRNNbAW0acVxxql
BLr8CfFZ3WsBfdvPE3dBKSzvOQjSux1PAlHsn7W4S/mnTf3ygpSbXuwZ8A4Q4i2i
uooGulW+XRmw16AmXzjr++StqYSdpHB4ZbT5HNdCuEv/ISHngsAFdoYqdmRdP1Pq
ah7jjagaKYscwr45Brzk7WXwfTrXYoi2zEDTPSfyeYg6e7fZRq8s+7bD4RpntYPU
Z7n7O/7c78/o2qU9JoLav/cF/c78QE+rQAi2MC2FNHJEFVXOnh03CbVgCVExUE7J
um0uQ3J2MtPIhHuP9d5xykYkZsHm6rQ5KEW/PzC2RQK9RgBvC3nxP0AUz/tddNrx
CH2k9c7GWlySUVCryBZhuEE03Qqr2WGlXImLr/rJ0QqUMP4/PLiEktEoLMHYif1H
FIkbaCMJ+ZxdflHC6xtrPEZLMuhQlg5nAmXgpSLVNwSa3uH98nIZmMbJgy0jo2UO
9DFwYMIjx2kJr3oEJqtzG2MUrQD/G7/yozEcRR+Zz3ruY97LV3T0tWbN8hVTx4vn
8qO/p8UzfVlQh5W6LwwbklgsWNm1Yo3X4BcAPvGMzCIwPqCddlSlGHOHkiKAHPbG
2Eqv3cF3vZLJQ9fafh2iLup8yS6eTQl5fKrU/eOqO6Iv38oYu6Y8bxX5viG37/AJ
5nX49cxMyGW5SNrtwel0a6h1LDCBs/wramW9PLs5t37g+AGvpHdUh/OsKwKecsfP
HN9rB+/ssq9TVKm+3CYKss9/mE62k5nIDJlgEuBL2rS8bCK1uWziQn+Vgzcwo0lj
bk22xICWDL0j56ox3h4RaSsCdz0/hyRcUO0LufcXsHe9Qs79dJqmhXoDtsM3OKX1
zwWcqC+k+BVMCG3xrmY+dncgHGowUa/opLJoaFAC9XbkUOvdNwsWHIcJJsmbz1tQ
JSorhpQun4AjA7J/IObcRzRPGB1oFiIwKNIrnRt5z2a3F/1z1O9btpS0azczVA1c
jBog29dVIjMcFL7AdOz6UiAvNcOI5BMmnwIX9IJ0Pj5yNz0mKXnLjqB1Hj3SETd8
ruGuCizqUx5lAAc9HgGt7nkaZ7x0aUJPliH2KM2KVSt9obqCUcqrRcoySj/vIF3y
GBa2Ws1TMVTQqAZEOCEcycah3m38Q3tJa//WHexl4uUvEymOEJW8r91q9hLKcaWG
uECQmNsCzNnisljtPxlB3Gm1+EsbC001nov7Ul08zIlCysu33LgWYW9sFPAQFEPi
HNDE/qZFDfBFY4K+Aaw1Z9WbCR10s3bkLme0IEHlVwwE6RVHQ0S+oq1+Rc/uKvCd
4BpioGL04zfmH/S2/LdLQxRl+x8ZV8R4LdiOKA+ieaxDkVHrkUcRSYAF4SX1gWo8
CgQqZeF+GWv2lBHfTSG0AB0yktK+Pd/VFsgSnDuODKGSg+9fuUgeO4dVwvuAlbOg
bVE0qEfQCcDJpJXieNvt2dOpedC5A4+cP09/II4OyHGspQ4f1pihW8QYKbI8t61R
DT8OXdd0kmpXne1Uz8EwtnGLgC9oucnniVMzVMFo5PuWNb68uw2pOprwnZ14Wule
x/G/wqkRQd9s+lw3h1REY+WuNsJzgk/OYdbprPRqNOZcm7f5Fbfqw4GtRNaqloPE
zJm10wznqmCT8tW/PHhPrTdfqPvEjXbGQ1nHJ86vokLe7WYQ7icpNaakwipP+ZIk
yuHrYTliQzZXJeHssoslcmIN2os4u1NfgT6kzfl9+RqiZZxvskutzx7Iqta9OAlc
iiq/Li3msm/Be6bG9tWbOXz04vMaZmXQ/q8YkRdgw0qemKA11EvNCuxPMgBW3JJo
tTxpMaNfup92QGIxPT0bEVfhy2pDHQF+a+2PXdMsUd/xqi/UJkXVMzA0TiPc4JwY
UbN/oRzVICh9pQnJkly4XswU+NgoRFxbrKQAabqAm+fEaPDABBEF2C/AezrRYw9n
XVmO9D7QU1VLRDvwip8ujVtWJMUllyTq1R48ISFq+Yw3hhRJb0ZorMen6pAkWIHx
txtMACWZWT6QtBX0eRaXPDrzaboA4IZYn7s65/eEqcMqE0qHt86ps3a/7nihA/JA
Z57zmjH1oAYiiMj7NxjlOYuakSGBksLpTaCHuWTsvSNkdiDfzQ6769YHZR+MB/U/
hNligMkKFub3wYOzxTQz6n2UD64Ttq5yxF0ir9WV9+z/MFg7V1q3RzZkSlNMhlN7
ycNu174OS4CyjXOY+06JRIxuV1pDiUBKc0Vdcm5aiDPMpcADHHaU348i32O3O0eo
qm3+rfRDKYnaRmzNZZwwyLiKbjZNXGLsflTfQZozt9yIe8WoV9TwBS85WH73qxEs
x1pGYn722nqZY5uHkGbrUP1mWytHGNryxdXlalvWLqs9i0oNPbA6XG5TEaTnY1nC
yXJrW7+fUa7TzEl+7G6MeXcHSNARLKEEqt6mAO5tOi/oNGw20BQvRg8q6zeuy1ob
moEIJuidXGJzdpKDix2vmzTWRKF1MwnW7lYHKPNWo0/efHphQqnqgHqpJx1NQIAi
qhn7BrHv6XvtPcGI2rjw5WVVitVpRPLCgNNJtpNkhCgL6d1ZoKGFTpm85teQT8pr
2z3tEOH0IZhmzLqCvXzXNf523/KXFlQ0oABIZZe+T3PV4SsLYqiskeA5NCflSvj+
3TzA/2x4U63H02uOflpBuSp0DlQVkS+/Dr/ALeaH77IvLIrjQa69H6m43AOTBIht
1HDPvH0kdsrVuZwokoHB1o/PiZoFezDJd6tZNhmItbHKzE4nLa5twjUAKW8zw1ff
NpO6hItZ3+Smc+O77KNqbC4WZs5jGCHcsahvHP0blEDFvfbLRBPgCGssHICE9f0r
KzKeDYthS1/q1C/WhGL2S7vZVojChI46wIpeQ0p0xqlbpcuNvw79qpn31fYGTl6H
hPNWmhqtiQbSevh7mlaYVLlE+WSbZc5lEh6wq6LeyVuG24WrxYbsFPBka8kcHGxL
4r8fqnVjj3Rm7fSbf+mc9xH7b2xMXdSyMLJ+SlGfEtReCfAff1ExIoPxZ72XL2Pe
JgaU+Pn+w99Ml5284dpLOk5MXCOxayi9zZQJkwlj8NX7zSGwvpY3OPCweBUDHeYV
WsGjW09Y7VUjO+YOBJJcxzzvRYD0ZEVhLV0fZx5TrXN33SXGbwohnwf77uIwlHkr
F065+cNWzWKzx3I+4RM0ysB4TScJWQrocrQfRmLECNBTRfecEx36xIdvwE4Z5qZN
CkrefdjuUC0ZxX0XlqDOSfVvD1YovSHVMlNjyo0wVjkHPwgt12lb0QYG+HNOng/X
p6VLZq0HTLZ7U+F8cw3bNGB4EmatLhQaDrL/OhQhYTdkbDb7fQucBUk4VLLrUncZ
+Pv0cBiEwYEoXjqHKJp6r0yW8L8OzKXhzczYoSc+wvPBa8KjOdYChb/PcmHHYNFN
XJhkig0JH2Gjz44lSuB2MFDEWNhOAE0KTiXlXS9o+cQEdIpxFSKKnFcl58gbsCcm
I4JtOlCpRykIUiHB01NSWgX0C7vHpS8RRmYBwS7napC/gOkeji8ZgoVFr8sZxnar
ipMFAY6UTa1yhklBrTq/RCiLuNPS2RuL2024XaLM1koUTiFQjowRlBqEnDtdUI59
mg4JUgy30o6ebL7NRK3h61ZurQ1BslM0PbeK7oCbEwrFwjg4a56P+duSAarIuod6
itneOM5IUnd5GTeMHrj9nGsMe+upP1pmyvwBqjnhKzYI5HkYz4OcbzIPVhTPWtgP
LNxZuTThopi1kFRt8nbY8Fm/t+aQK2gGV3KUrNx9sabQu6LL0B1ozsFLKw/Hlmt4
IHDKIY0yiODo/+ZXXrPmwF3OF0F9w3nhohbVUfCjIXQxjjPTWn1o2hQO49vya7GY
31g95rqx9VHj84fzL+HVYGWURiR0RRXGVXHDHPqogKhgUMrdqBL/h6Gk1n0pAnvf
c00wV6/myzew19VyEaYzq0dJGmmRzSL2fRiAKAKF7eyFvB4ruaImebqD4ctFvlW5
HWCuGEBAo/Rphkkq+S1whqzGbiGVimdANGGGBStObJLghXbgEACPFcNyy7m3zTrV
ijIuoBycw38bEOxoIZopNev++ZtRBVfbqh4ZsVn0L0p5ce/lf1epQuzdTkaHzJa7
uiKJ5ad9PCSMbmDLzZkOX9uD4j8dx+rGRKDaPUUS9gdfbQsPb28rP98lW75NBCFe
IoM84caRTZW2sMBCCIgf29kIhEk0Jb4nP/CNQ427A5TCn88NsX5PHBG4/FmLYspj
PNSGZ9VF1Ksw9pA8ev+noTWgH6G3abZ+/adqt7Oat4b/0N/pBdrMaWQriaBP6UjX
g/c24MndGzppFtel6rHTri4GDJK1Fn8O/14CtjKVea9whdhSZR9CBaG2eumBInlD
s99XpvvqBwj4jeh/pH5Jh8Avsp9q47irt6DG9pAqoWIp3sMHcv3njGjf/lTzzBC2
lcvo/fbGXAzDJV/LaZMc1BjQpZU3iTlPwdrsK5HRscWXGlPg/a6k1d0xPQarxZVb
F/3g0Hns+1CsrW8dGBFpxDFhr3UUGMsWJzPqosvvvf264cWgcWPEPyGdkEam4yCD
Res6fHN4KQI8+ug/z8lH3RZvkLyprm63q93TmACZs6G7cA7vLXhoxSCJKtQIcQ86
72ksDwMXlYLeZMppdiXN3X2SQfTEcKD5JQ5OwtEXXWMnp857w2i7ISXP2Lece0bg
GYQfODzaqcOsP9lL/iYmzjObMeQdgVf6R4MslwZG49rh0zG+Z/HLtL0U0TKB59hY
HgCZz/123hH9Sqex7PBNXrurRJ3vd7lfrqVi+5DUZ9csQKEhN2Tke3TjjlJIuBiY
nQ5A+eXyk+VfmGmN3Q54fn6b6NSP19LDIlRpjHLDwe6kLKXq1gVe6a9X999s30iJ
7+taS1YfZBADeLlZ5cFntNbb6wUOGynjpRA9YocwARr8+TsiaH5y9Va3xr4Y+j/1
JgpSGbQpyrF0XoiijQNsT1obqToZ6S9IqVXUQYRAQqU8zt2CYBUh7t6fdUSSnq+e
M2zA2Mti1/NnJtYKvgGz7a/CPlfPP/tQZKwNyNlzUgefgC39U3fNoUWey1kYlHZ1
f+W+nWz4xcwROgvtPXamFxUclvac5TeOibepTizUknXA6iHdnUASY+oYpmZsQV+I
ojMXh9JUW3cywdQZo/BNmnh58vPbKZeadttf2VQStxEB/IQOrGOIhvcymwNDcGXH
m+kYUt+COxp8X2K/sU0lS3tyH3CZPCmvuU/0svaW1KSuNvc/eAdp8zr8S3lWb81Y
r/aViDynLwO2U0fByhrtPaX0VOQQU3CSrCAzpUnjOb/QShLSskw8qUWm9N+8SMhA
4vVW2UZ6EYpK5t/vCvu3o/hd2bLDgQsjl42LPK8fgnq0Pi/SViRxFL4rYTH4Gl81
oE1li8zOBD0tx0wFXZNbWzYstYVxhlTAt9pqJi93kwCbLbjNQRT558JJJF7eBuIS
hAoUpPLBBgzxpB9fvpaMKq56oY4K41rVkn9+NPay3X4KJH9I7YRrjMpQpznsWAl6
O4ZYK84RjTcueuN/4zJ4Zdp+vT0+kTV9b0ytgjk5iheCkUssCuUgjznrasuEBkBB
hSc+8xAkf2BHf0M9KDSaDd84UjNTXascYtzMB2M1A8k3u9Gb71FtZ1ubC9zCkxOa
OJ7ICOEewyC5tuwrvgf/d4An3iBny9T4zXKjbFtkDgiXOhenLHI+MC3O6uPprfUy
E5/uF5suCWQTYj6ooNxzhA3H1Kj6RP2dsrvZ2VYBTcRMDefYZ7v+FSghvbbG38c6
tnqhZzGyU52r03WROMosI3IOf5eK7FpGFhh9EyWh76/jwHSFSOsmguzx/P9iLk6m
DjXZLdEUeX/M6QiD6scr6GVS7J5zHcnmQwNlfMgcBs2yfto9j80UGmqcIDHVhSw/
Z4r5Z+YHRB/EIywrnF3YCdPjKmm4QGZ8p5Lj/HDzQ7gw+h9VDsDDLvaFaJvFzGoB
Jv50hd/ux/Re6IlBlKc/8C1U2snDSvNQyqXkoLSvXzwg1B5NwA/iuqEDWZTTEAgc
Hr7uglDOfqM/chpXlvZKBUwGenrdRX+wNL9Iq4gBikCBtj8WynWB0Va+G3XfYUng
wiUgFfD8eTjQf8afm5rABrjlIVVaaA7ljVkQjDxC9Vo487jEJTAmqFI3idiSzQSL
QgZeFy4/GzwcWwZxNqmUoobRSC0B5h3rmffSfC1m2RnuRLGEd45Xq3/KL32GVTf/
tCyyjiv0/GKJ8RWFNwI/nXDoPDH8MV0U0/3W64kog4NoqKjdseh7nWNBx1QXk6JD
/1zvDIJSPQCtZpm7L7mfS5YiFnnRNtyzqUCZI/N1ikGJVCciRh3feRqEiBdvjVKO
pOcqDotOTklXfu8thRZHoSV5mCctf//GKqtCy9F5Jtm7feZhuFf+4UuvyCcxPMyI
AG6+4QPfDzaTkI2WZmQ2rEhtmC/yZAfH4CgHsNSJQtnsy3mOgQr/hrvscGK4gIH8
zJPMCQ2g57N+DIgk5GAWEXtO2282+uJnkGdASZXn0eWlZms5BIhtfaO3shfYcbDH
SjkfYTH/urZZC+dXWndVlLeK1KaI8i7/rRIVD+X7xch9dEUTc5h6x7hN/kDwm9Bi
/1WBSChajPYGOHIDVNoF7MPF9T3O0mHS4XyJUgoyxq/JeNrvkZQQePVGGoJideoC
GY4kuijLVt7yu2VpjqUo2kNiuNyG1xkLFDHxlWEFgF6EolzdUnQKJoIjDVOkd6tk
G8OA+Y8IwxIbIxBri1DbBnVDzbp1lODpddC+61fGw3Gbntu96oaNL6DPrSubw4LC
W3tYJG/ROM5GrconggsAL4o9gshNtzrTzcXWMKOXHRRjhkP3MYjH+zdT2E0F83nq
iryut0ONBqUUm/m4rj1yD8DQgr2hSIFDsdhxfx3lqjIIhaBnMSiL1ocxWWSznYOw
oXlRSaKzq3tmzsv1zdxR4pMGkF/zgNzEAW4s4x+kkHHeQr8WKjksNlGvt2Zn8kI+
WgxTQSOE3mrXBvQzsVSh1BCdN/JK0x8ZEEbiC/r0do0yY6Iew2WFjIOKXSCCFeiU
LOI/bQSH1vx4t4HMmdSyh+YUbl+PHgDJFmKyg71nfhIUC5BVLgbWYQf2fkIedSd3
pBVdVCXeqntsHGk8wa2g9588lpjlmQwboxlt4zOhthCUK4F9q8zuvCT7ApSVXGt3
kQDyhAbMPG0bys8AAvW0UrAeC7JN5QFHN5JVGeq3+9iJX4c9/hUZTHUEbpSH8vEe
Rcz+pavnpmoVDIZo5tj1khTOSFxjDeienKCVSjFobtzewq5qtFVi0+6OuGkq9GGE
3QohDtOG3bC/eSPfvN/ePZ53zSGyiVmavxmBilPiAEn98BakiU4C6KOwnaM5dD9l
kh/NTH16+IOVpLYnFBy5nySu5/9EjFgLMLfxbnhOt4MoWmYsak3nntRYmpbMjAqI
wIRgD9qVexlajUGyMDIZ9WD2m275acXq3dEFa1c804fLfQAt4Qn1v4i/a1lyPqtw
Z3hZepB75hBJgfktgMM5rrtMs02es2RhKUhaZ+sWQsZbrGSFOKNyV3oE4BR3gu56
pi8hQilmWjS1qkqA23f3N5XmGiAnepMZmcyJWsmywH47E8GLo9UIrJrjiw2SYLb+
bw2CZ7JHGY1WlCGBSv9+OBdcK4wjFpWjhQrJz6+5InrQs2O5OPMewYWmCbppetk2
fl3E/rlS6ZJ6Y9Dh7LJzrsQWnVDYwE+X8aCxf01Ax3TNbR7y8VMmh0jN7ZWHRWsg
XqOr9ggdl6bxL7gCUhhZf3JFdg23M83L45tSfHZ6i7lfEU1zaOnu/wRRdkU0GUAw
7LZ0d68Dhrda6K6o1arokM6xson/TNAeMaYHyUgWo+l7JbA9t5/qTwbfOmx64v3A
6xylWJyz6YZUxmQgGOwtVzK7Oo6UTzi+PrOAuIIjG+y4uHSF4KdxkZzn99A3nvUe
0wn+ryY/5S4aVHAacGViK7mbh36+2pva6sx4mlXhfFQGejRthS9JGM+UqU7SgHv4
qbPNlkwi6X9pHn7O/YczVP+6G7b5rUjtBW0Tzi6ANEPL2f5p9dFjURSSfb5n9nRg
7CrBcLwn+vHGjpi/8Axg26FRwTPRtCxSedRw8vX1FCYeFLcTMFAthQVHbNwiDUYC
lUS2ZZqOM0Q/q12ra9oBIWV0/pgyfWtww9icwjTOnxf7dDXHsQN5pAMDnPYys5n6
QzduPwWJOrNyQbNgGczxhE5H7LpDtnC6rp8AbxRyP/oD7wpNSIDFdajwU31kV5WX
BnI0LLtKQ7FNShL9MZYPvMyKeAi33T6H4yA/DprYPt5Mr+Tzst+2PCXJu5Do5DWR
aj1zp0FyK6OJOBDSK6lLpoeeknIEmMCd0e0B4IsaIzEoX0EQNR7bfO+doQhHLS3W
fN+1KSlCCTgkj7yG0GNc9v7RvIWb7IDxZpwrazsxamHq4qYPBgBiYrl3yvQ7sktF
2CEfgx4nm2XNw6t5RKXXX3Dm15d+4jIMFNWKUn+OGnZ6anuTR0/S+h001Y5eVp1d
7AXNxFwER+A1Yx/7aE8fTRI7Cxhr/Re4svB59Q8bOmuJAdNCsYj2qOwUvJk5N/cr
6sKoC3PA7xpU+rd65Zs3dvPLw01gUFDRPk9wZx6siT3tnBphXeBaR87MVgJ8iEcp
AkKeK2re+aJvaiOcTL/gnL6BqvqWc8ckgy1UCCpnsxGlj/09JZXs1kYhBESYjc6t
b7zKT/Ia8dFpn6hAssXGV5MucZdyCeFHHvjMIeRhka7lhJRHyGNl4fhB0B6ptb4T
Sq5RxC4dWQK4xTm+zQPbpGEXtkXneFeE2AS4mOL2CARpfNwDC45PjJVJvmsBefNf
0TcPwkm8jzFaBvedruWcQw/p95y1GO2t1mdrVQji91VfNDUbUfjcVcNlGwZr85f4
IYApMM5Ex3Bi1VD1fLTHksKsApo4Ju5Jiqxlz1/xu9OtRxcpNAhKZQXEj5H4vBUi
1/Roww91iEEkI8/aLrBE08uTFOT/rYIVk3EtEX8/9cq8w9Ea+xcwwgpz48XzqLwi
Fnq09A1Sx/npGS6pClNYWsdxnNVv9SPGvAnx1cCwJ3MWgnsKs8ROfskY84qcwPfl
02i9+bX+YAuoCpTLKIFOvMUe3XLGGhhMqtoHcgYrtIU0KL3vykgRqaBUAJG01eHp
rUsl0QJjPpkolxGL10fkNpmS0zfjPpuvmki/cvKoRQiramel7fnoUHcp8DhPGH2A
jGn8LvGJ+AGW9/5jAA/Q4zCL/oYkUohOsaxz3RfvOv0tilqn6w2Q7wsgLNI75mH6
Fc2UgeQNxQ2R2ks4ea1+DgMn1rnf0uYrwhuoocq5QKuHaCHlQnz4xDhP0v0f8UuX
AvE3xCdTIJAq6fKToV3Tx8TRvg12CGQpw1lbJXVzo8NLwwyzEhr+oAuCHqf1jhZd
12eB6F1BPLchIpV5MOW87PaHKAeNKRiYAf35PG1sf6IjMJ4bGZzby5n7rh+/JCmT
rPOhBwQp2jAkwJO1Dw5ZlVIhhRBKTz72ka5VMelm6o/5Bqht0lLHj711gbXDrgz9
qzhklPfJ/5DDE+kvpV7TOPuLJhemsZICn2Ior/7tqgJtG8tE9aeg76o9jySamVAv
p1+jG3OEl4hksQPHxcQ6IrF/e8v7auYNmlmK5oHsb7VhMlYl5MmxKQN0WYpNzFZt
BsaZOWtKyAW3vv6DzZ0ahla8GWgqtJzEjz7ygyBHIE84G7wJcsQh6TBAzI0Z/T6A
6NtBUcPUB+IXU05ntg5JhnfR7P4yETproKm9CHuShnoeumjG+X03A/kvYouU9PHA
M3EPmYwT4FDBsl11m19RCGZU48TIKzBK/BcluD0UW4H97YRbnV4TOQTPH3UTj15G
Naq+8KIHtZf+0+QlKoajq/jtUAaPtMiVczxjQB1CrRFUClNARkozDzMTCnjtNt7Y
21UB1Y/4XmD94g1XOziLuiHcvYChHPdo6Hz1OYzeFLxUR2io+M3yG3SGU6BnhDur
Vqb7wAyZh3v/q7BqUAJ4JIYYRMCMiBFqh+rjAjbOC9MjHK5R7NoOeTJ065XkATj0
oCsHkLG7gAljBrsQ8//fyqQTCp+T4axf+mDumguM+NPpSgAoNmJZMwIReO5x0Maj
jlNQHf5aXYmhsGLE26GCnJ/dJcDFc75x4W+9uR7ke99or67/Ov5PFBk6hLzXKW26
PSLoc9w846XH+7HrD7O3AWg0BHqAZfT5bZY7jRKr/rfgsZZp5KRiGWz2r8w4HEQH
lOZRdBB0SeEmVmX5TgIAXE2hRCX3gCgBfVukinOXtCWndkkvmWbH95Ldal+fqSCA
m9VLMeRuyUC+WwUOO1dXeZAxGyB1OlF5Wb07Gj+nhdrR08K0UrDrtnCuIu0LxnZ2
KcCS1z3gKKUN6GYm/nZrXz5+DQKuKY03ley0r9Q2RT6GyWmsS7Z+JeNoaTnZQF7l
Lyjv51duiGyoeNzNHyKpNje3ziMG/m+pod+yf5X2fNNE2Txkj0Y93/ulFd6vj2BV
pKL/g/rlbI5NiueYsoHlSbbk7uIoW6Se0RXkJAIZsm27cakjURjGF+obYmbmkmjk
RlWOVxAC0Yq6aeajj6XRyJld9HfCKSJck+kw6Vc4PVIAjg4kGhD5yAaFIoXyMHBZ
tORW9JcD2oe4UQhsszOQLNe0B6ksteQgVpxILOomhnWQPG6TQWzzH6cnELqv9Jvz
Q2FPmSXLnFWllQye+H5n+CmmzsVKfxcsioTUV26xHcIubCav7CwsRBEvSkLYz9Kj
acEllnD9vo4HJh6FxmJoMCcnql1wgCCTL4hr1dsKF7c9N2r1CGBusomQpDJLc2WO
1I2u89O30L/n52tCByho0elLRmztgN9wSxrdErLmKwN1gOLyOz0WVK44tuMgiCSC
R0cso1/i+91cI0iiJZxVK8aK6Ff12lYVU0L0CHO7kO3/f/t7bUhgZ1eUcr8G2S/A
DXj088l4RMXLIFdwY99ueqLl4uA2bOO3D9d4VqUSkp1Q4MJnveEI+Ab5I4ojzFNH
NV5aZPi7tai2Jo4Urq1qPqaqADok50JKWuiyRh79wfY16b2Yj8zpmw1StX+bHTsY
akLpUmRfSLizYLbDh3cA2nwRHcUWOzVQG229S7yDdxX85T+Z5hxiUULaKL46M7P3
O/0LzvgF55LRoiCHLIiD/5zA23AIgq3BM3VY92Ul5W7fZe3PyBk+jYuCx28mxXgu
Te07WKCnQo+gjmYBVnDpKKspzaijVAiVXVkMWV4FFYakSTaZ2+ZpzyxvXc1RSFC+
AzId8ifekcewS5HWxfgrUCK+i51eSaDiTGihIjihRzgdnA4RpEX88LCraRo8LZF9
YH9rYf31Q4q20lq/wumQ3t/4AIewePYaYE2/Js5pwPcwcvkyaB8dND38r1AqZKv0
+88JwU3TfeOElyF/XQbuj/D8VrJzNy8UVLsXTgt2n3qtIJsCJ4OOxXLe731ovR0u
zsB6uErImpTTVeCEgYApdEUybw0kn+2xb6OXhI83Dhtwjf4Cf9XeYN3bjiXNwR6n
Q16I92MKx8ozzH2/yNZxcouvVbh+5QgwmUaPYFU11H3fB9g/Z7fJUEL8+dPhvwkb
O/oOiCPl+0s8wQCbvDqa/L1UnqsxKW4n8Au75U/OLMGAoNotg9GG2Lt+LAqmQ0FM
34WicysFyvZQ5TFEMC0jAMstk833RHsdKa9vuxvTxOsSQk0Fn3ISBPGGzD1VTSgd
DRdn/5BELDJHeJdR8pbEmExM1HIynEerKVjqdVo8fVVp/8QxLyKJCpawu11/m31m
QhuvuRzd/9nFYXU0NmDVPaAuyk3pyfbwSi1xnEedA5KK4tkTzVBhXni2GqtVXgms
EFBR1dv+vg2nBDNLG1iVsvl+qhLLCcxKq7N23BKSbHtl8n4V9UJijAZHFeNFIYiT
g3EQhTreUeW0GYI0ycZSJjVGl6DG5wyF16O56BS9CLRvuCU8FZ6ktViEEZl9eaHS
+S1HHQt5+psH4koZd0R4/vWnnlGQkFoCbt1s5yT1kDShGN78VV1aKnAr+rDHPe3Z
jQLptak0buWreA5ILkqh0wXeHVCwWL/yuimfPJ/ega3Bu9DHIMpekF6iWZaLON+a
XIjADrroC5RbeFZxFCUHIuiXNELcAfQNTMPX/oDEhsArUzFkmJaM1mOkbHpehmIn
ioeArILu03soc83N9ShgCvRX4h0e9kzPNuXkOoblshXjqznhq8bN8MJPQ1LURM3T
8Bdl44PVuThiWz1fgvd5DpFlP7lmFifVdjCswoxah3OASSuFfv3LlhhEYV/2TMFY
medRdo4XLzc4b9yhSc3ju9XVfXVA5Z1TFpAHOcgeasnZZjw7OpV+mMr5IF26y6pC
5TlAXwkh51l87ZbrVtavMhAbyk8VUuVFHDr0Iiws8PZNkAGrTW0DC0i7lINntCAt
QTdxy1099BAv/ZBJSOvD9S6UbZe4FRvIEc2EHUT+LuRRnKRDpGOMOH7UIgKlewz4
ihyHKSenoZ/0Nfh7+0fRwv5TqDpwcHzg1PXB/axEuLFcqrFQbabXBJVyHn58FMZc
iWA58wav3zO+uqzaet3SYLqKCLVzRnAqjEqP7ZH1okcIOc9LxBN1Puc12hjUtOaL
EJ226zy/j/is5IVDXGocJ8Z18z40p8jcV1Sljj5fLAx80jf6aCj44eY9HPXo3dPW
xXyV/NC8SHcTlN45aJTxDSLzBtTPyK7Y+RTk7XX4jgQL1tSRicknET8qJcejPvpp
X2L3lgouz5lxgeIUZirR6CQtjEb/HmihKnWczLTARVqSPaYOHULsoXdtlcI4aaJz
kBN3DY67jwX7vOaFcMTreRDE2QKqY5lv5dxgeSHkhsDfoSIg5dFrYIjFSSkVOtk8
YRR4LRHOW93kTOGSkCWCiIN0oaKAGaDstq9PgPB8nwtwUiTjcjnW/Pd/wEgc/jHJ
xk2Y4K32N53xkGLdAVxByMBIUZj7XGqlpUydxGB2dilUGOMmAUI7iGZhsZGDOvjJ
Mm6hPoO4q/ueJ8CI3R0wWdnmUOHRjR1iqEkv8OFWbOLkptsdWkf4M+NBt6F58/LT
Kj4SB+kF4SChzkB781FiUpFDn93mY9KJ1cl+q5RcGfo00TaX8acLCqLLZmQnJt9i
pJuzYLacnxG05JVUkIBjscB9XDfWtBEyU8GiPM8qFy/DOV6KvsYyCd5KQGTBEHeQ
k6GjL9VgOoz3R0hOQtLVY6IGO48KadHP6Y+Uxfcq/l0LTNTXXLGGiQhA+XLe+NsF
ymgQ540peGp7QvgCzUgcakIP4KIZXuuvcLKDR1Bc2JEi2tAD3wB7VML+/uBhX0mr
6wgVId9+8iAW1Yj2RijofZqcZbfQtRg7JdimmQYH8zGB+H+biF3r3LrR2vPUd8A5
vJpUqIVbEv1bUuGi2YIhqaYhDDVwNirIHJKZyEXRq0JUsTjqOBKFbI/MCQMSjvQo
sErWbju++/cHZRa9TagO5QbKGfSWdWmDyLIr/8OO7o7ZIqVqrDO1AFs7AMyeTkWC
BkNqetU+v/TW8v0TRLoQQXuWzyutTVZejchUGsRyjZUaphRF4RcQWaqCgkc5tLAB
0ZKc9d1PVqS8mfMqyIZnige+lL38hn/40BnaI5JjdabUVvHtAizupOWI/uKMprza
HCje86aSggOTEoV7ea24iu9GE3YUp/YAY5NQX9bQDjaPFv4Jp+SFb5+7d2ms4RRw
jREr2ET/Unb8xuXdDbaHKRtDwwKCT0FNnvNwYZNbPjs1fGsP9ErOH3gChfjzrBa8
WKLF/raHEFjoDfnGHMVWX+3rMzNUmm4IjEUEq1cK1FD5Lod0uMV7VJQnpHAN3szo
cL8nmz8pBYyJseVZ1oQEpY/sq4tngTPALf0LibaZbxD4P/q6I32Ly7/3peQtMRjH
dusjRrR6B1s6Q7TrtSUmO6XZVBeYEGaNU/+SwuqMAVmNWqhb19rJu51ryw3BS28b
NENh14Qc3ghOopP3Tcwazw9Cdcvh1k/aASwiz44/EQ44dUXa0Vh91tDiFKV3iMRO
oIiiRSbI/c3UElqlxgiGM7VeLHDQ82+d6AnF4rKqk6UUWlYIv8DCSvHV1u8ObPfS
3p7xizQ7FfThNtm5sAV13gcaTzO8fet0rqhl6b9uSlxmm+kZnCKoXWcLq2otIPuA
zw4LNAEJmwL2r3LbiqYGpuXZbjPFOTLyKuIZfB3v55nWOBWdNZhpMcPOoRudvKAc
qffgAdwuAwGOV0j4wLR0X5fDyxRI5q4dZW8aFs7rPF8kw+fOi0UkAvNi3H1MZwh5
O5jMihrYHEeLXAaWRS5nQtJpg6SI8Y0RhnflgSvLHWBED2/wgVycMwJkmu0EFeBB
1s8CdKRAWGmD1XFrllwFDquLKG6QnKVaNS/+YUtgqnLPHo/tdq7nf8m6NyHgMf9u
bfY6wucN2nCEI66VJvIea857RtEsbLCe+GcT9SMDgnlL/b86OC5l5SIhZpqu75an
jjh58to1iphnASCIi+0kk+MG1jqGpJx9SBIXhDW5BoStmA1tg3eSkBYR1BliM2CQ
D6LK2o2DJuO3YAQkUnoF5IiInwvQ3LaZ1bAvYTb8o3JzvOCmxSZo8uxXUxSSqvEv
l27F20fxIHNGJ5q2F2bS3bpMS6mAchrQiXdOrRMN0FNjZOJs5lJrsPFl3uOoGu3E
FL+qfjwzaEXz8tN4vq63/SRwgQgLjbFNLgFUS5uv8CUc+pMFMaa9oEeXpookX261
k1IjZ8DqFZps21qP5/qXWARDnPfyW3tkQfivTvzuKXnky56d3ad15WZ0RYolQ5zh
KG+j8ehOhwsomZW4lM80VcS+G/xJhHRjOiy1BA8+javX8WcJrO730RKeHvZSVYIA
pSvSE1b7yBoX58DEEZvRX4lWHgPrNMEqjfYA0MF+2RTKlSyRwlYaB7yEyfG1fGiL
Zq/M+5/lgw9RLdOLV+snYC+edO/4ayXrMXHf/0XO7y2biHidGch6XaNFMzlKW8QB
9V52FFICY+vktVZxPNROZeX5yDTngEaGNyNUXyzvx4Y7bbbg3OJTx/25f6YF5V0W
Cy6B2pfspzaRvMYup9dHg50ttbTTq7GhfyjcVgWlls/dG1dHEiSf63NSmN+4oouy
nRHy1/uFlpiNRJVUF71si396255CQDWIBujV02bZ5ueHXoO/elFoO5hFYvlcxl/5
Ha70TySWM0fOlSkOL/5jNbhPVC+hrkval/r6T3ZA6HJIXmV355JSDo3mMhMulUOT
0ki+pi09ZP0bGSbFNUTD3RKv1fKQOE1yBdIWXF+YzHDN3E3+DvWfaujmBimW3on8
9F4q2O0wfwEb0ROmWoML7pJUkuJKOOAtcMIYIeXV313M28W5iA54bktKcnNvwf0x
5UBEeazWSE9p7lWC2VV09VXtqZiJIfvd9sYzDRqtN606DJLmEIJqPqI9bxXch2LJ
1TyJvz3hQvICodHWfXW4oIRdeWXyq7HrASnj2AS2jeqhWZLEsPp54b+pUgsC/lqT
TnEQxdY3i3GMHdLL/KZdGztSl/uiaKqpqCC+1I89OalBWB9uUEkCGRsE+iIwPlFS
M3nojtnnbhQrc8/B5SnqmMSV7wDTL482HB2UoIIb1keWzJrGwsi5JAKcM+luomDz
CJ3wa4mQLHwuCdmXnaHRxy5VNtnov97y0nfYjTO+YEZ+yjP9MhscN0AMXIwPsDYT
XPASSOTx/hp0ZGdfKQOWpAHE3kb/mLusluqmPwgI9weGyuYPHCJDDhaTkevhBARu
8I3wmpO442OkCLDqiVJUZxs2MPY0uOM2cRlc5FU2WQ/IzKWi1T7H223sdabF7qWB
6Gjt7tyAeH0BxXX6ojZmd+zZ+eEI4PvHn2+eiHfd/q8aBIROg8941nBGb0lTaeVw
U8OUNfR4LM3usPXTNBV6il9T+ZITlQxpsCxyYfPbIey27BInNZ0UFUx+/d4OG/XG
vYzAjYJ3Ho+GOpuZ8m+hW/xo3ahkeOp5sCkyiHPSVkzXWhff16v2FBxpL38PYcsi
xp/3vZZ1my1LQsJKK2s5yzdT+MLjACpbTDauIZijNPJ/xMS0v0Q9rfRBvzA6Lel3
QL//LP5THZWXLd75yE4PdSwPfmyS5ZnUNDqKut5SxBQIqMZYt3BYrN/TrqaHrm82
WzrvXbPU/bD4uT02p1qxLNCg+3/B6iw2z4SK+hi2kzyW5Gb+8UQ36H/cCOPDkwzw
shBrTz41AXsL54CjmCn4LaziZ8cvAUjmnAapC2Z/NlHcvQjZrpO5XMJ0QbiTHYW2
2qp6jeLHICM/4OapE+IPGFbrUPDd8CqkYTgYUhKHeyujPhKB6FdQWM/SigTLFQBm
mgkdLqSR7rPJqMejw3rUbqBVr8JFGIkX0VtDCfvuWqHAGABDGZrXHxm0AVVAsNmL
jRZuw4nf78VFS4J18Xd3Uo0J/KMCMUQxZECd5TbvxMACApAgsO4gh6+EHQubq9ar
KaEJxdPW6p+MMsghWpvp5nQ60d8vlGZEJT7AN9A8NRWL0LbJKFcva6p0mjGe3NUL
9QwJSaI84YiWmGNoI6bImpkJ0rldeuy5Gr6MRW9HLWmcXmGjgXQ0Oqq0wvvXu5GX
zPi1xivmyGFNeepdK7uMWRYawxKIfLiH1E7YDqxv1aLrfj0ACIwVdR5brWFYKvSI
uRZ1+8hA2zGuSA8SFfb8qzZghZo2d0pVcvO6b2ISGJg7vfop49TzGB4mTR1pSMAa
OO2YH5CXhxJAnGj29GrTaG6q+xv9lUeoNzIXdicWBf05LHthdI9gWtg4NeSBWJu1
LymOV/cJMXPf77zto+AcG3aK8C04CYCI8BxATig2W9h1r0O5nKjyas+ZTPWO21++
oXFj4qAtNyRqCw7Y5Zzd7ftm4Ml8qJwgIusdxBqochh4GK1nhyYEYSH/wLe4IudV
Bi3Sncob3b1W4wYxQQx0kycJc53kbEKUXWzcba7kpq1TjhCF3UCuBUZt81Lpej1u
1Q7wVo2CF0h4R9n69vkryF9ZyhLjMze9qFStOcy9MeVR/hZV4UYBrbwif6+7wf7U
Bstf3pfTegozxJEe1KJrjqYiZu4b7eZe4zm458OfTWfUY4L+SD1WKFIqRqJcUTfp
sLEo9y/ATKiUA8wH9wQfPFJ4FR7N/NINnUdS9vVJSVq4KgKflCetKYuai7l8Me+U
Abk2tJmdzbuTSdYyHeLfw1tAeEmZZcwmovQwujl1apkMeoqXfsaFcKU4y49aW0I8
6rUOOLQAThZNk5gSPV9fJLwcNX3Hd9kF2bTxFZMoYFLdP1IBOhd/hZnLOqbN8okK
KK1pqRjSYF4OjzbqQgkqXcEnwhrn+kXdnm5hcj6f/pMOvYYMVY41QANzpJwjpVDm
j0vfzCuxxooLyrLFwzcLdCYxOuFFy5dgxUl+1psckDWSV8MR4vc6Fa9bhBpWavSf
4NnNeLKWZ4B1Ei5fOy5xkjFYFUOeFalj/wsmHiy13b9z7nZIap0VVzqHPgwipVgX
GJp6y1mMrYEIZZ3ToDXVlfJFxOJEfupu8LIzbyDBdw15HEAU/FIqmRlRIrB/Aajl
Dhq9R8Bh+TrR9z6nIclgGJeOrxzh3IWMssyNkfACZhTFt8psEWiJHV8UPwcNeFzn
1FdY9cTWor/9Wv5vzc20MDXzMgPBk5r3CG+h1Rk+k+0fRuO+eFkaExOU2OS7WJpI
3C+RGpHetI7IM2eC50UPP80BDpRV0PzwGNxrp+wMzqiqceySi4/zQKS7OtIp68Ln
MnzQcrOky6XRQ4mkj5f4lOi28krfUceQOXAs6bgEC0dlD4VmkmMHpuOOJ+dekZah
ogfG1zoM/YBCSefy4sqJgushJQvm+iCNna+8aiWhZkio/D93/EOwu/AYNB6DaqmQ
mfRtE1wgzpZ2e3xqWLUrP82qZAihtflYwLcJ4+Kt/NhVeLdPoJYX7QZd+azZUI5l
P+iVzWa1vFkSh8rpmX0jjijg3fkMkDu8UDBzSeuumkAxWj10iEMMIWaAaLVX5unG
dwh3PY6XZ2fMlO+bFvSddzFNYWnjtR2mvBmGFuTl+phywvKSCu9xSJeuZnzYLUgV
FR6a+HQQElpGxLTSgC/l2Mh0sk5EZwUbdIqbWtATF0oDYeFB2MsJt2Ju3/TN5/S2
xtUoOdD6G1qzUNkJ9WIOl7CkampgbB5HP8TgFxFRB1JspLPd0JLhyl02K4I6iO29
1bEP5aR/IOo1/OXSmbH4Ff/RzJu6UO+dIqSjP1ghmetL/BpApinp/kdoCIz2OXJK
jPePHf4vzl5w4qD0ZD/FAi43/Ixur5ju6EObCb7D38csdxYTdEMzmLEDT3A+ZT7B
is+TmnokVIig2htpOAwE8kGFQDRtHdJGliYaedfuWWQmdi0EbomcS62CU9szxjDk
ghgQj+iTjfLv3G4Bp68uB0K1afaQ1gVO11UYuPYDtSEMaHS/uyDiNat5SkDopqIN
mwzecPtv6Gdz49zrCPRYt+DsxBlc+NOk8abJq8d0a3ukNzRHzT7VLP17SJ8wvHNu
Tbunl8WY18oJXt8T1oE0GuZCf4xHpkwDzh4sH6+qC1biqXhar30qCX9CbmFvdEVS
jmsSMhuCo3+TrKaa2acigUthwTOugWhLEzJ21+cAfrCts9nsXDVpGd5CN+ugfcGc
5KlcodeSCRRtE+ocOfoFb0i0/uU3utvCa5C6zmSIFvAqnHAj1rBmZ3rcgImCOPUo
jxKRRGxpsKzcKUaDs7tQELyGevb3yPe5PmmCemihOUwSoisf3kB6xRu/RklbWmr/
Q2F/1+mtRHkI+P+7+YHLVgFrMNkw5sHLuzMCnTZRVLViQUCJTrKyMqJZTGGl3LGd
cvybhpwmgSVne57Td+/D+xn9Q2rPc+XtYaiUHi9kQe8oEajSm9Tv9gEQYrHWsjHG
fgLVo3qFojNDOaUBlonhm71E/N50FjkB2wOtIw1HzKcAEOelYnbxEYD+/gLEHWTi
Mnm9rKC3i7/+APz4Mf3yky2Ha01RVNAs8egXirceQyLKyAuhoG9iwe4WfA8qSf5L
2LH/7LHEHQ7Mf7UHLmzNIet8r5hPvSO0dKnkk/e7ojv8n2Uspd2CdibkG9EtIt6T
arjU/rU3b5TdSidscjjLB1see1Ag5ZcEzaDHiXscLr0xzKSRbN6IG9y6b1wcg3Ys
e+QDc3vCAf7mwYAezXHkdLHgWZ6BbwFihHaBY6i9tl+q+1NQwNhRJ+Uydbd6UZJo
dEpDQQKyz5RxSBi1h/UJ69ToIas67kJcW/mRtxh+sSbehX+OmC6viZBBE8x1QvvA
JNShGJpGhZYIjRp2Gr32JMm4HzugxZF5GGY5XYz9UlVqeBuamFf/b3pBdOFAg1Rp
BrdFDUcwRemD5hwckH+rA9hmwC3fr2lpPzMsgClE8RfCkiImKZUD/66aMFk39mLG
SOWitTGn/1Ckh8rItlvFhU/wLkI8G0eEGz4+O64hBPZHYHpqKermwUj8+f/aRon6
Rh5FdGNIAtC2S8EyeLZzvZzufZByZT2RT6Xs3S+GceRA1puIoiTL+eTThOevLtTT
1ZcNe/PWUd86qdwnPaM8aDGApOyD5SmI+QcMF1rZdpyLh3AWv/LwLyK2hjV7U5rw
xill+odRuGb92FdI93xOtRTNuSt1RW6mdIJwUlJr3jhF5Z6Pa6aS9eWWyNVs7g7F
XaGKmBxePA9iI66FkCcDJIiFITCMi8Q9JdAlb5GHyb0Qi2DY1oW/k/MwbIjDfjJ7
yRpXZDggTWT4cNl2K40Pcj1coFd7SD2D46rlAHROW+LnH+BdJ1HOGtaIvEQVjqq3
ad4qvWpXICpCv3NavWWh3vAlH+Uhwbim8XeMGH+Bn+VhPvmrubl/E/IibEhtjF+7
jcdwTchNAZbpG+wShBPPR5uSulq+j9Aj+wXLh++KxVyGljLbDjhlaX5u/8OQ57G4
gh5J6DGp5xaZh/F36CB7ZWhB9JAsz/BmMhxbWHTPIhr7kRmkzyMwQHsPF0jvjE0V
LZnuh2xFXyY8mcZUecfN6mHdZ0eOD3XgR2iDpOTpfEoWMY0cviCJ36QZ5fLXroNr
/gUOHK2PxXjxRwcYxwgvI/wRZiV2tIoZ7lEZAjxyBDTK4hHr6YD/hiD0sEXQpVFA
AkA/x2V8WEeG2iJ+ucJGKqcUSg6RtogIcOilMaBZLBtXLd0S8r2pUoYTifuq4xAX
hSGzn1ifl5qr5JCQ3CkEaXoi3Z1Ir9ovg+y6NPX0MgMwMDyl51NZkUkwlCNFUPP7
nOiu94BCHj3E1PMfY92qY2nn8t7djkMxqqWqq1iXleGIWbWzrx/I3mX0F6SvszPP
Fb5FSgaMchuP23jtMqkSL82Xsoebq532pbwt1RpvmKE10Ye5PQYsFji4n2OL9B4Z
7cgbufg95UzXXObsldku7vdRx61zjcfyoWi5PUx5k5J/ieYAQnGuRFru8kgkB3HW
uQIZ/oPZKEgVDegYNy8pAE93P1/esJPtkzrklWCOrZrm8ZGLemeCFiHDR+LVEnds
4rWJeneu9pYTwijMZsM+oo1RXCz7zb5h2s0H3TwueJUoagD1ZE5pTFeRqNbCUNhA
u/W4hMQNa2k1KDYHMxVsn78BQqoRr34Npam+xEa4ccqJuXKRCXAjNn2aVS9EWce3
ShnUFOw+3URA98KfP6LOpAUyrjo/G0laBAV6RrYtdMFRSfXNJKfvY1usgqg5cZCv
IGr0zoyBbohVyE34OZHII9oIPYavF7AdsqncfKREUW+2Kkd3jurjrE/TKqNToEJv
4+FWdKJEnsabobxgpMWQlf+Di8bRKGputUTwNphLRnNdX3z9gihoGXbZkEKJpwbg
tV7e1A+8W7DL+wdK747u7Ry+E2t+2HU8BMr2wylNxzrWc9VQAseWzgEol8vGjLqc
sjt/LbrBRAyD8Q1rTLMj4ZfJulm2+wcXmvq1Qd61jCQAkw0OYiL+I14pIN+Ym8RM
kkWhjPWpFg84cIWIFc/IHRoD3nH71I+7lEnUHoLvFhaSbHjP89NNuLhZKR3gnhsn
mcvd6ZBqd/Vb0nxEezX6RicTXowLYZ8qbNTBhXlMKidL9OOBfJuvLtsokO2vWg6L
hxxckFjlas32bzrc69w/eFxOyUuKlzpZvG+7+TI/sXDq1gkARovLPrTYLidr9e8W
LJxG3l88rTuWr+9gwYsoiiac8BuZ0O/qkS6QYPz/gf6MsKbt/mqnwzRssIqu4iti
/eu/jRzzwsxFOQdVt5vwcfM7KM2L2H2+7dWbJ920Pf5AxJ1E6jucgmBZs+PzjD4d
YYI5vuyaxLGRMexlBvyeA9ZiRTmb9D691tpYFM1TtcrlJzjXwB51Q0FWr164+Eg3
Ubhgwby7a3AU1nFPEuxstoqFctrQUX6BycKPGZrnBX/dvpsdxqwCRmJpZrHmU0T+
7lHR/Wv69rqBGUSxT5hK5EYxw/T9YqsPen3C1w5i3CsdOX+1fURH1kOyUoll41kh
rJ7v2s06nch7IeGXuXhhXb/UtBqwu9mW9Kpk/bw3b4wGBUHxjtyeKNY+B/wGsyjh
y15gBB264iIr8FOdbr93M4clc5hH9HrroVI6nWofEArzZPZOoSR2dg2Ry/cVrQ0R
zxgunMQOWauKGkwqUCKWC2IjeGv9mahH4Jb7Qn4rLkX/3oD8QVrOf5ZorHB6D7W5
ec79bljlCVmLAUbk+6Gl0dq2MR/FxzXptC2dMrfmH46NOfLfR+DpxTG4AtJ0F9nF
FbUGAFMEq0FGy5FZJ9oHvSUwssOdtWwjL5/t4wGDLyvcSOtcSu5PUWqS2IGHJRcj
fjFmtpo+0F/fHJNwxTSTrpBWHlmycqSodcgr4aceDAVGrbAiI9hd7GeuyUPF68X2
zERdKvL+DjWSaEGz5FeOag8+Cgs6Bi/m31CwUNBUruXATAh3WKZBTpD5zQ9WKLyI
Ec21fLzMxCdTcRxF9EGTED78giBTd+Hdgu3WB6JVP9iGoLz3mbFl7Vm7jtcdeP59
1IRQF+5lHun1YB6ora8PPRtA0FJfy6Uk+cz9o1Jk+dSwpdN5WongQjgAHLeYQX39
HF31jUi7t7BrMEanT37jM9UIUXGQ0oQ/0z2dlbxwpeBlNU86cMIpeZsx/mjQNlEB
z5U5pWVV2bE+HLaLmAG2JDtNBPekpe//18S7ptsKSkWC8MW2hKK0L+OsgQOYQQsd
9nln2P+bofz632Xr8zmFiF9Le71NgX1GInoCsykcYvrmhOxvmPaEic/3Q49LzMhI
TyDtEkrvKtFBwdh4PsjS+aA8yRsFRfNRlUz4U2aXGdGML2Z5jMCUIY3/Ic8V8Qzm
2VpupPuafCbmFjJeX706a+UTzYoS5WwN8qmvFOJhitRV9cLWpiJ0orWJy9VObCcI
4kFrcMMugxN3gPHP2mPZC+J8ByA9p9GOSbPJZdnqawzg0oA9qEIRGuzACAYLw0v3
EXXlM4j4xKVCoHBkb+1Vb6qPtHanUj+V34wW3MTn6ENldGKKqDY/+1IRmPmTRqef
2l6/DGFuUon8n+77w03SSMNU8cthKp2+FoA+15Fh4LqR7jcJzWazk7yjyiCaNVlI
nQ+JR4nY0MHDdX5Kl47VnJoyTUSlY2OX6qxrIrIVsqd4ecAH1QAHgN7VAK12jY7M
CtqM3mww7G7vKeWbb3rXQAtsFHEs1JaMQc6VCHRcWEiIfUIjG//UqPoUVr5Hdv0X
RD6/hw5JQPzjPEr9wOMGIG2oZDoSzRerWf1uVIFAjO7YE9kS+oQ8fn0R+z6pyRWg
xBDkK3u7t3wXVQlYYTn1xjuQcm+dByqL8FzMVshg9WQetksgi0SOOra+aqMYhVzf
wnJ5CMCDa1zs7myJKn8pXOQIb1vGzjgmYAtwzPWQN7yD3yf1otBoJmoO/nNCj2uB
O/iGr8447T/p7zwNIPeMd07ejEz0Qmu2Tr1HR0BituabBu38GD0b0EBUCV3JZH60
gM/Qz5iyVExswCuZZcVyOp7zNIeCh6zfv4fsKeSss0LfqxLsCHVjOHXKcR6QcTsY
CbkqoVkR9lLsFAEDYN0RWZB6cbbFz8IKML+mrKwWdieO4AcHQ/MFvBss5ULto9/U
scHqam+FhYgz5CA8jXGUZP0rZVZDAa+Krla9YZMDGef/tTIpLrMxz6oUhdtRs/VF
YWRHmvsdqxbQ/43N0BQESwP3iaLJEbvY5XyJlXAyzUVZP6iogjIyy9eX9qYS0oeR
XBoqWDtvlsta9pNGnNCG5kdJGheVKWC58VfK8e4EVM6jfA9S6RS5N6s6By5CEp6+
+Q1p4/skReppoJhadHpd/5ZtLOcCUz80Hy54Ma3ilxTuEOtaKeTO1We24dy5awQE
jLQ3w1L2+3CPOhp/sytilpXQxBzVvnfVw57oT9vX/f7CGY6mtHZLJnWrKrK3mM29
1wGSfYwORCBDriA1RKUujB7pmOUI2AX/L7kirYaHEVxGOx6IL+bLoAKa7dD0g7dd
PpZufBKoh6xM1rj3lGSXnwzZ3HGWDLgKtUnioNDAmdrYn6WsIS5vMI2wy/uAYTSf
e4VvKISCgXkiFAQPX3F9kHkD+7ifi4DHrE5rxIXKGJC2zpQ9qeYG6i/ohOaLEObK
V9gqBTrQP1bCCatka5KQLj/x4fbftVU0am96RkMPLizMVFIMDBNyEqXgfBzeD2Jf
1emrk040vZv7Z+Ig8F6RSQ8jnOLf5jCYQgEM8vuAwTsZAU4l4K8jpM1h2B7Fe6EO
yynBIr6jVGzyqdqbjj3t7M4+G/g7iOZdVyGxsvq/S0ph6W2jsYeWFFyW5vhdP4YL
x/cJvpr7PhkwQVUeiBi3XH9EWuvT88PtiJO3sRKMTD43LPa3kGEcTHBFh97igUup
ISzJPheUlosqGryG9JQ4lLrlaIHU2tGFNiK6Kh3bONVpC8PU+WpJktLyI3DmRzMi
EenXJDJSue6f+WIAtsleBJavHOdPVoNLelXQwGvPrrfIKvAqF55OUGa8Itx/2DFH
BjRu55D3KVg3dJJdtICCCDcQOWePQErTMckaAA1bNLSrf0rUm1AIvMG2Twwi7P7A
b/JG6ttJFmpMfnF3P9EiNzTQK+waPb4K1E4H6xsEoBbbxW+A8iRc39wgJJqWpLok
kBOlSENQgnXMc8OAg9sLslvWd9dVA2i36DZDZyTc6tWTQMCEL86y/3dApwOMUkwa
Tx0G1CMblDxH51eDrKTWUq2vUuPPR2mIdX6mMO9PFmlS6OnjBzau0+Pdcgnf5QGF
8SJ+sGFXMblMN9NUaLugXLif4bNq1eWtuqfcP+ed6QZjiJVQDHqeri34Nl3sMNlU
rW3LU93fu0BXnjQXtr+ZJWAs0i/QQhNQLtHECGKbDRzwH5j4BVqusqcYFZaflJSk
p1fl9mg071AwJK7pD55wVW+lrXOVDe3oDcBHZmNifdk0jVf+Bj4eYWQxIvUeNhi2
9TJDEeG1Sdmb3DLI+2rxVMqvrc1HmSjpfG0EtRHQYFclb2umIzGSBrGzBbbKGt4Z
99mF7800ImLLXZCiR6KZ2de4qWb4pSseRrKqOmV8F/T3Chltv6URPhnB0Ed8LEA1
RJilvVNkxvSIk+laQRvhqU768E+3VYrYr7hCTSq6ZQqYlFHJwe4E5BWbbfilNs0A
vwHIb/4VfscKRXvLk09qpV+P6qs2Me2akGj6ArifMvp/tELObQThGwQkD5jO49DS
RuqLJtpfjyZWu5G7U2faQQ/Vd2s9QBSelNAqQ6VUaQT8QYarwyH46ZN6NNLvrVSn
WKaYtoOIvx9ZtyIxgSoTbiCMgJOZ3AEdDFS8yU5qY5uCG1Ldpytr/E0PiBjUcLkN
Ga9NO17Z4vknchV3OTMacKdUSldmvd9lNWk8M3mljF7DWSBrCA50zLtVRQ/8n2i1
SU/bsGzkcU92go0+xRZ9d+JZMDBEyA+HRKmWLqSoiJuScpTf2lW5GScRVzvt3R9c
I9kjRkkcHE12MIX2jhPhzj4FWtO+CusE0+xYOZ8tkGIUKInGkvagDy0y6rV5WUGh
865HLTYRmGFk/1GiHeB2XKwcNahjLQSSVRhbwY3cqNHXh4Ocpe0irpMlLZGTvBBi
o5Sdl5wEj12YePAoGwDtTvEb1zbQPo2IirO2CPbCvjZhn8HambBvj1+XiLD7EtFv
BFfCPX1gg5wT/Sx5PHdWFDrnsgFopo7ZIyKFrzY7T5y0TTS2cYpyYrVnq2MzQSYe
aiBUF8c7g8gDf7kO1RGlyH1dVYA1pQH8byJ+C0/bbug3bLdsgtCYdrSr8MR6c+qL
8OWLuo73RBlBKgumODioGm7m3+DoHwIw1ryMOdbnGrzZoEKC61n3HAxNaGjhIRJq
kIWb8U68XTxp8dnisXKCqw1PsJHgvusqMfrQcVSYcJB06qTRl9Yjrb5WWfxe2EGo
9XOR0p7TX4ilR2saX4o6czEY7IMgadA9iAT3XIxPqwrA3KdQXg3ENs7+eE8Rmg0G
fTxYiHv1xOvaFRHI87mQXxFqMsiIEQtIsvexLBun8gxQsqT9393BEEClvjAol1wg
+/8sB5FMMwizTRXqFeJhK2qXEn0tEMGSpJYWNOHfIYWYBAOASMMGBgIo82dlJRs5
DA05zwk079Us6DcmuonY2hqVoaPLMbFz54BFUQWwTuKih77WiPK2TMiUZdm12rCa
ncpAilqNCA3BoK9IZIDEgfyAUEarMaASr9CaLO1x4RQiqCtLwc0wo0rr00xPbGf8
zbvyDvECEiiVPC2sHTrbMJ+IIgq8LzMlc6zOE5fW+afTDHCoxiF3UCyet/zPHroC
qIgbdncLXbbGqlEQouCFTR9scIKj0l9qq/VjixQAmyXB+SffWahamJoP7SNXmyMj
LWiqQ+MT8J3I2+7BZer05ZQqEhjQu0ableZ5UxIRvZfx6VzXAejp5+RaDynPSbOl
e4WYu8lkFSkAen933qE7shmnZKyYOmmW8PPMDSHg8Ufot6O3SghMFAY1boBHmRYJ
j96HWBc5w6/vknsNFZZAv7C08jPZRR0jlfmJ0LGO1a0oMZkhqYiZUpxmd2jIk4lW
Dg5hBgojnuWUKmzPLtvYCWpwqAC4NvBpMSGc7Io1UQOVMloELvIlYoqcu+IbXUZp
roqygr2+pxfrhoGkSsLcYhl0OBwpIDU9wVB5P5ya6/NVqDAbM0SpYdmHn3gMa97E
A3A83rwfowgSgfJYtzBwv2eZuHnF1DQtaRhmHzc8mf44Uht4R3j3mNt936Pzqs+/
wecroV3NloC+9PMJY5BtE1P2V3T1T7EwvvS0l1LUPbog3iP8JgsRMY5JKqxRdKRL
4aHMtrdqYoFjf/ThVdjHuLz3pUZe7dp5rmy9rt9k6X0vMFIgKbcTS90fkqT/Yx11
UZ2D/h41nd28u368XXQJcwfk7C5C2RUXoZPbeat9cNqQqlzCF+gOR7+1ac5c3FVm
zzNIcCgzQUxRaDAD+FBZS4ugOhIgIZKGu7K+MsjR31TcbabKWHWNr4D6qxbPlp7r
FlJc+OM4JOUo3BqCjYuRcqKGN9UWrdRnbTeAM5UeVR//pxwyOQHI4KWFym18HGg7
5OCYInPMt9TmTV9wQ4zTDAt5xfj+R/0dsEKHlJgZa/P3l1AP9WyFSraIFO/yzj3m
JclY/b6JJ748o8Wjgn8UdEhp5BcDtiBQAH8CEYvmO7zWhzpxb0m6LnveHMAWGqQO
Va6GOWi2p146iAkN/6TjfUCXKsXwtK9PzXW1/ZbiOrmXqKP2Xi80c05ZMjkuvTrz
CPW1BRbIKkPROAt3KTTQs+oUSkgat3EpNJUYbIJREuSovYGEKXJCm1Y3vQDUFDvd
2PR+a/Yyg9BAtssz0ZT7ttTB5GzaHg0YrDf7gpr2n1nBtFaeK+UN9mcmgBHseF41
YDeng73R8boD4evTghNMcLBEMyOpeUuK6S+qFw6hFY4pKrHvat5nunfGb+55en8c
QH8pcpOXasTGEnaO3eRVS4Elkjy/Sd1xoRblcmA+c2DvTuDFMeUcj5Bn/A6qKrC4
R6TFMA5uT3l+toV9bWN9UvecDcUFEaFIxRXA96PH9kOsLMWEdrk6eGiEv8uZO1FI
Lt/bLmVS25iX/xYX7fSquybbdkUOyOtty+blV688mdjJPRz23iasI3hFNcqotft2
o9TqDSgp4XsKjKPacgTYc0lXnH1rNkkyD5rd3iJPmngRo+1feoXXydtEGWf2sOYU
ZWflySGBfvZSTdCGPnK1A4O1M3Gvi3RnbcsS7cEoPCHz5XYjmELYcJMgsWqELxao
OEenw55Pf+ZSazOLeVEJ8gJ0GAzomG28TSu8M5W7IDB8aaUZ01xOFWSdXuulD77v
ETfC4wVo6QQhEHMrZlcSIRHlz3fuAjvsWFj3geHG6N4LFveTODqCY2kI/GhxqtR2
8xKWRDAUYGqtWEEyVURg2rsI9QDZt6fYgDOoY2EQNxSlD7hHIPG/5rjSvXBBq6hn
VyevLnwhSzmCdZ1wBbr219pLlWmRuo7OkgelR+jcm/cFaofKMRpOS+4MGkmIZTzK
/jI5fcmKHtTVQvK13REdwPoFEZVruYvdhLBSRTFPtqpWKRIJBSGvmVhuUZ1X/zxj
Jg+Oll3o1lrhzoDcQEX7M+mHUb/HgbbXLOtu9hV8hNK7lIQoANLEoODVKAGUC0Te
WamPwI3v01yV8WyQ+zmUQ6lwEKrXiVMMetEEQpTf3vvtonFO0Yn7xyn9Bq6HJAhj
sVdYGeTnS5yz/cKA6dVuiMQusLGckbdTOC607Sx6capILWPhhBjcfSNqfY0Q3MFK
0PalK2f1l7GA8BJlw8q+CobAyABbX2QdCDOwwHLw45Y3x4WasfTdAB6bCiZIJ1fM
ljSqvaLTedzSQBIgOcQficrmikFPgSvr9M0dj2g4x57ETjdInOV7txF3MNwG531U
r/BCzfX5Kt6W7tmKTajZlrrv+NStk5Nhbk8gQqRCRLT0Au4fszGMuWbWHRL1NJuq
93ej+fhewr9EU7I7srcOBhtShZ8OZp+wo045OYDIKGwAnKwUfYscZ/hBshCZtquw
+SLNGewAYGICabduA8R1V/hCQMcC9Pcrb37WScGIs2UMqKPfCFRYga79anyMGEWn
9a/2N1PdeRIywT6bn0SCmRikb1MzPMs9edV36zaF8bBj8lhuhVc+eUoQQ41dAYNL
BD7Bxsg+rhe5VaqAeSoHNqLjfitWBQi6FGuSzsy7ngv4Fz0poT9mrZud30lfNr0I
7WAoZxG3y7nnpPHaTXDSQ50PQm2rCkOmSv2WUaV/b+zLjgvNkcl6v7PaqCWGeXRw
3mDQN6GVnpU+wmATYKDGuE16RVGlCgmXR2AU3Cg5vVqYcWNN+W9g16DWYQc/h8GY
QwbwkuN0EyQwMGtY4SY39MiNC2vZPQXzZlXRVdtZ4GJcQIbfBpJLANQSaKEPxiOn
z7Qx5RZ4u397AARlhL3LYFoh92ISBatMzm+M8ShrxPgvugVnu/0wvZM8hxV+OksU
vTjsbbqtQ/frHrJstqQSJCXLN9F7+SA9sT0fTRfKClqv/50zSpTOxmdiYg79Ofob
5LJBO0PU8UFJiJXI1oMT/GRvj8/atvjCc5JzY1NntuCXfOd190HE0YsPjDVjFD86
Z0slhCHXzMft4RYvPEibsLXjsGpRczCNySr6LPJGJM6uQB7PrUYMQlNGgLTMgZ5P
QZO/8qRVpxTZMhH9tF00pBcaMD62nR4K0XzFNJAItKsf69VELwjFHIKVhj7axJ3L
JDY8DVL5lkYx3Im5EqRG5ufWrFkCObCSuYeqSAwwnlJdaoCd0mojqDtfZw7fmO+O
8dIDcCxeh3uFGb9IAGieDlT1lxKK6e0IyKP2njC8K21cOqy3HBIqcXHJdSTnblla
oRQIBusM8rXV9o0rq9FeAkKdOQwYbLjcGXz3TmHoPdfjzM1BubqJ892y/R3+cNgH
iTJ3qwywYMYTBJ/+SCYFUk059W8c+i9+hYZr5bYdtL/ORon949s9AcQ0T85AUkxg
iEKYDbR8j+n4AtGiSqpoEi/W3SEYToR+OINUeTc1D81EKAAsHSw/f4UFmPzxJw8l
WYo+hUQyjErmse/9MotflsTYZYfAjjmpjoGphtTYcaEC7cBupij29Fi42cEN3siF
1xWK8EKSl6TAe4DUuQ/qyoEyC2PIimlXL1GJgftoFPn/fk1UvU9R9LIs8pj/x0Nj
LkswtEvkoOseOeFrAzi3hzdvkZKV9WcG0LZ8+hhBEiU1KbYUO9x5OCB41yXM7/+1
5qFflsbNw+9wia06B4BEs+zzLI/oPGq8J9OM7SX2wXj8P0RSNaZ8bDvVI+Q/kIUF
IYVYT7+H9DMDOP36CrEr/ubm+4laZ271iXZNcoi0h6HKuL7VIH0gPO4HbOTG3jUU
x+gjlze5XaiQKzfiYl62UbEepYk3gKrR/l8miY4GnU745GvKUrRHBobOfbTLLMqq
KVUpy6sf+N8HhICVZ8cmVbbyl7Lq/5KfnuAG01tjNaiTEQLFUVnNE0CpTXFnA5BJ
XmBe1pCyVVwHKYhXiarjx8LqtUT2u5EXnsXrAuI0AvHcHC+hr7W0gX2Hoyam8PGl
SiJVKBw9KR6rVgBoPElYyVQTe6jn7zHySmCqsN1mIZJYubjzU9jD4RPIkCwlliIx
tO03kFVYDJX6XZh4sa/lQCHyyTGJb2BojFRNrBraxW38NpZjdmloU4oPn4ebx1Ll
u9IL0CXlITwwpSH1IJ+//zR8GtraKIPejiYd/HRXeM4EcvVmIC3EggHASqzbTfwe
O1pWFgn4APzW58ov2hkWHIfcsso2m2wGEy96tGSeiS9hzIB1W1TDgiPRu/8SR45x
xZIRy+znTaGUpuF7ZN38skpNkuxi3R9qy7AETsEI7QrTuj/eLa8mlmysaXM4AUmC
8TKEkbEjv8Ps/9XurAFfesrJooIqPEgYmXBItJVPKcfmxSj3PvtDFR9o1DXhY6b0
CsoPhYgg8EHW5qrD4B7/lVqAXQZM0fKjhjn6Nyij7WZHGMxwHzA2YPVHDjSMRLUS
VNd8GnRMp8e9JX6dbzBiLCU8byhN7kBoLhTvZca/q1P6SuRceks2ndyWSATGqMdN
k+67OBuNvv2GfVfieyc+KTyBqkt2QCfWJUGCLvU+LTUIDg2ECCvA4fgzprstqrUa
idUeyPl4raCVIozXOxChxe/LwFLhBMHWPlpAToEscGrdp4PQp66jHmspzvQHyXri
/iMPFTKfCm+tH1MUdE+YUKykar/atIkU46oogwC7IP8Lw9emFY75fK4sm1iUsmKb
1ERBTL6cQNgdEZgbwEiQjS0ljpDJ+J5fyxqIgJtKPDKSvnzbWUk+1xe3TzJEj8TE
cAyvstJEPeDKAj8TkcyWuYhMwt1pIKAnFM60mcbhnuSIRWLSdldQRM6dVtKxFaBm
RD1eVeRWHea8isDUIsPbGS+e9zDelq/fqiAMpAuAdR/RqC4wvakxs/FCrKkJ3nSW
tzeMYHa075r3zleyX5wKet2Izl5nkSUpbIZj69wHR0OtUCNUR7HIEWe9tgt9rhQG
XLUNqXCjqkHvnS1b3ZB315nW5Pq+YiQ8KwyxyHIBaLY4QmkFytwO574fPPNO7/lV
fMX1Il1mJ9CdinPgA+gTTtj6M+iEKU9PaARmqJNH1Hp98ci6Ki6/UDzq//KmadBa
rHm3nbYiClQ6swyiLzdkBv/fhFLLM3gdustuecjXid4P2nGGm1wzPzjJMsWrnvfz
WEqOaabu8qMzky1uC37q+j20/hy6+qdBctIcZ9lLfDG0e8cb9oQpiyTYmAaTjZts
ITzpuWbE83M9bwmVhPv04SUNMnRtc7ExD9c+UDNEA7RcT9ztaqYdiFZO2H/dCo9w
ABUCtCkkKnlz1lNQbipNsyXZxlq44S/nrBKrEZiPDHNPxBkhR8d5rHWxMXCbyBjx
EeEg2eNqV9X7HgW0S8LgG4mJnVoEMDuEf/08jekQCy2FHbnqkqNOcAo2t5KqE2VJ
9Z9B0o4OAoSVpWKhkHSLWOOJdaCdFiWNbphucHnJmgXDE1zXRPpbdc/2xHzC9Eet
13E1/+eeTpGzzhqXFBL78er3Ur7WnEf5TldglE0b8aaZknoqTFRBmvVooboVSGkz
Q9dZ67OjKBSptdEepxJ1lrDCi/3obDIxvrPos0/BpSquXuLYTl3y7Dm3TA17btn0
ww/VHTB1g9R/bkglfH9tv8WIYLnwEUboz2vXrcIJZDxZzpZZjNmC/6BA3LoVLUry
9dHjlYvkE7kAIuoKfXM6P6vONTVFtN521F/1Zgr0IKOlh8eukHZ0w2My0FDrFreH
mhoqcLd/vKmer/GXRd4V41KUso13u6d6x1xNtAwzKw+2i/+/W2Bh1U7kOIgcIsdp
CC2m+g6w0PcLBC60ujcTZyOMFs59StbqmIIez6r8vraq6vltXI1F07jVDYz43pv+
W4QlNVOe1hEIrkLj/pKC2wdwKzylrtipal49MdofQ+Yxg/kwr2fSuMLrAvFPdPKL
teRy62PvkCiYG8GawW9YleQxehM6DqyF1AkTrao6EsQ4JZCMIyns3XGtqbawPXp7
3KTShPNCepXiEQ7IhO3jhUf7Nj/hgXfTrJhA4PKnvp+5ukImB/VpvvmCC7WEwNc3
/bS6l/ALXEDAoOUVmwqmDe8kQeMZ8PhwN0T7X6XSKqVFJ7Ulnxz+RxcQ34IcnqQN
ceziokE3q5dySqWvJUWS2pwBjSs9pUIs7qH+WwC3PkBGvNavOuroYUur3nZqsLKu
pOf8ttB8f7HL390WX+PrZVkUmmb3XHp9qixYwaDxc/5TujehsaxdUwunnKGQfH9C
xn2uO5XC+mm5ZZiaAE34/xfoduLXH2mPBJ25rCWZchlA3cb5MtYOL1uloklpGvEt
o9Kaziz19vYw/M5gKZ2OwSCkulxNjhemV4R2H9TJpcUwgr+mBwFKu4UdSK7IJI5P
DCTdQoBN81QkO5ZwWmtsQX5qoiX2ROPPXAwSKTNJmA6WgbvCVXqVrNukgHIGzYJy
GWRQZLKjg9n2uViU6vpn+bf8Rr56AKjF4sNVoi3wHIBC+wpvX9wb5p+TNCvUB1ui
LoOtOkHrXpBajLqooQRczHwKNybPfGo04vaV89qDh/8XWZ9BFZbwEwR2ursKFKcT
mu3KR8eydjgJRpn9A9O7K7SN4wCfCH7L07KS5u3xkZVLpKmu7jmHUZR5sPp8AL6Q
Uew6kq/ICqOw69tpE7/iSix/fbWmzuNQewqMoqHsFkVEgCfGQSFWsb7VvFPmaGB9
l7HQg3nX9wuLskzNYILQSVeo5MGVpLIfast0zA2oMyIUNT3psHOFXZg2vMqe4Aj1
OoUJ/E2hMHuzhgMZG35ZwY6ZUqT12d4p5Nba8S8h+J/eyzADRBXbHth/CTEz04jR
J1mLRCbl748qL5P2CrcMPomHQzrfReiVNX4G/cduWbbra8HATsjOJ3dwaXTFrKHK
Gg4O9Gh1Tjf8sLhuMqeV6YFr5J0PYTGLgrHuU5IrW9f0HKOpo9wCieAF0Sne76pH
pXrifKMF2Qt/gYMflM1LEzgI6PptAnrS3p/BJs9Rk4qTAxuKexIA9PcbmIwOT2w+
jNRNxPIPanmhv+3mClA3qlAzax9IvylBZ2QGoLYx/yThibt5mNH0Bet7lNejEwZT
OCWz+11oJy1yKuXub+UEyMIRPRrhW4q09f30y5JqWzX7Fly5t7TlWoC+e+aGd+YG
RvBHcDdFSoHLKllajRAQM4oW5rS61D7O0On7AuExjSuhcAZapEA/wPH0xuGOaHNx
416ZCgqS07NILysl6ADDaA60PV5FtY+Z1J7HzsPMDrjVRH1CmAmTBZDtD6mo/RlQ
yqIvveqmb6xKoaTf7ZUmEwSiqJ1f4V7o0293GvEZ1yhOfS+pjMA3mLVVyowgnwNg
pQrxhlzyamQjyPS9hhAP0n/w5Fp6aPqPI/se1RJa1TjgielDAI2le0GvMoWWxP3b
ENbPLlgYDFzACblYbiRjP97cCJ56HtNBj1mwPL0UV1RpD3dN1Qs1tYQ0Nfj1Y0Fv
J32BYdF2p1G/F/vY3fw8a1hAiIx9FwJuinoyzuV7XHcElrAASkIrvM0SgMaczege
vd1GdUk5JlvNcClaEkOz8QcHwHqyW6kWevsfXp3APtHFMPhfeSF+Ye6OAxcpqUft
uPoe8GfEShVu/Wpcfp7oYY0vjR5y6VYHdqSGGUXbdFxY56+ooKekRlhSoj+iTGpm
gRbVv8ATdzJ6dBxhn4lThL0OHxGvWAYRyb2PmEQ8vnCt+rd+Ot3jccCIEfcDFIZg
KWv5h7emnAhPXvojggjKv1xIXHRZhSMnZfqD0iCJkET62jgq9qB/PJkFPVIavpeD
6TiUZDSsRfb+aFWFfedb3yRNn0csTJ7HyhxIQGYiYsrJzQH0kYkDcdyUZAcN2Bd3
hAwlSqKwCTIKOO5NHFY6vDHTabmt6aagBF0JfI7JfNn8dFKBokR3ouvykUFTwWeW
6FnbMPuBRV1douX9b2kUXvCH5hOK7EegYBLXELyaHlAn3D3qQL43I7h1kkRpUzd9
O+DNkelxXeW5BvXCAKzt6YIAskTeo7+dY4XeAavK5dkWDP1yDYMh9h3PIRx1C49p
i0+4vjYjUlhTNJmVxTMtKv8GQ5tlr6LpM1rd4h1Jrrq+pSK7dfcxa58OjtsH3IvP
YrB5pU0epwp7Zxl4WzPZZikt+wjZShYoQKX/lT+br4be/5sQbbQ1xccej6CsY2z3
sQMV7l5nqCzvxOv3aaRePJv4VhRC0cX8QVQ6Ppzh2O4IuV86FqfNG/ejdp2LP2H7
Z0NyCuQ/HR1kjcGDCb4136wYOQHXRLeZf8LAn6Q38x9TzpY2xP9y+99WCldvk+ng
IvSgXj5rO1VCBn8xr8cDkqxGLzWobuXj5c+CdJDtbWApAuaKRMnM91Vl5kzhNwxI
trDbEXnshfWBB5K+RQXcjGa15Kpi9OhibAonlpYybtVZDg2rGAWxYI99CnRyM6Gt
zUWx6knOtO56PKqoVyXq1VlA9v+Jn3g0iYKhJ68GWFBw5nKW1zKf/i8Ddvh/ydD6
wyPOqwLQnmRW56uYzae5ZbOe2t8nynz9JNxUkFE2elGbeHQYAs+rsrAPT2QN6G+v
Yc4gG5No0H5v/fMEoK8yXqahCC2VIRIlGWKC53OECoNEVydWnGwtRSa7yuPVO5Tv
ox98P8vbCBe1iEKIODjgYD1nWZMX6//w1VZxyQZA2wy2HogpICg7EHBCDwdjjQRz
DtKPe3KOmwTTLTxVkpoAB+EbGoewqxoLZEmlGgOzxqVFXc5en20nL+mipDjMgVQD
GxVf7tCCx7atCqfKM4/TwrwkCxRKpxG4GVm/YPyE1veyU3/eBA1orjESI9FM3wnT
1uC8Dr0X0yu60SN2SAHXNXJgG8pGNYyUtYM8DOCFF9fcOg8yWgSRHxF6bt1rpndv
RWWSdiHVbDHPMEESjXKiPcZOptr8DlQzssWTdd3DnHrb2uBrvooOFt8EG0QavL4z
hD26v9IcErmNxOsOCaVuXXqx/vuG+fXn2+DqjrU45T0j487VNqle5E+ggFdL8g3p
4o7orB3X+hqbyDiUbTbL35ALM8BtQEOWJkhp2MWQL7odIE1W2RSN67VRSF+ax59n
doQiSGJ/CjhoWvpQh9uVKbUASfIXWRIO4GuMdLxCJeUwqwfY2I0bkG0bdYQ3zERh
AsIUHt0gqEGxfcCAXlm6fSEuJ8XXoxp6L7yqPX03jgjkAdNmSm4XXg9QRkobP2OQ
/6t27tnUVi7kN6OMS3iLRt69ftlgLvea3FFEV9/g8n8MbZ/2SpSeXu+qql0HBIl0
rZcbTQQjYOJ32ej501TdQXmuLlvRe18rqRFjjMzmSXGkQFVgkiT2FZd/v4YOHPm2
jF4KOQVp/y1Kt9JKq78k6l7mDMhM6+q/yKlJF62xdv5pgLGhEC7YeLZ4Ho97i4OY
uv+aCAqZnE7yM2tSy1hZzGJibvCRd90zTgFOHHz3vgdoiDSSUPc89quvUIP6qFXA
6XNRMoWl3Uqrgo2KiNSuE5xpyvW4wh6vtvzcwsp4uN9J/WWqPMDWx1onv+0+eKbv
kisPy48HS3Jsh2+h0GzLEy8PvZTllwyNmUs3LEPgYoWnd6QAYzl30RuXNSPhBDtP
yfN9ku1zlYCudh6BY43NzJIZeGQszTXgMopm7OsTPZXjc6qjjzRadcc6i8ob4Eha
MDz0+UoAvH55VjM6UrpqRyq7m7QAozQMLiuk6n6Optdu5tTXoK9JHXZxJ50aPgfJ
8s2/wjSyxpKb+I6vL5sDh5xEifjNV9dZOJwBr6hOACgBMaErs3Gj/SosuieAg93T
aXSDvfD+fF7iukM61IoxtaOw69KiRk6XgMRAeDNoE1bzafQMwjiz0PKkd2jjQEjv
+q4z68G06lV6b3Ikm0YItdfnNakngJ/ibUlAqKfWcTtEQRRkxBK4P9F/CMdQyQVv
DeUsy/PzHlwypLk+NvsXx6e5WnCmhtmnFHoMwCXp/ECVdn+1+JdGNIBVxpHwrkdA
d6QorfkcQkvFC1d2LxiohITLRUZTOr2Z+s+sR7NyBTZeIA5rRazadC1yqYz/BLfo
90m8XQ4tA5Stl/Al4uS3lA5p0TcWZLXis9R6tOy8zJsrxmEuG4MoaTEKWFcwRLst
gBG8FaUv5RNtTqLsZEj0tj+IalHHz8mxj2Kbzj32OUugMhdumdsvx3KW5uQ/IFrJ
ZB1ICRLOBYp2A6/Iw/I5di8HKi9DSz5qydE1jxgwNaQuD+8LRdTHQJVbkM7RqdRC
GI81e1dB66rVlLaqxsUbF2XAs/sOnUQcWEKCmH5GfmtmHBgPDrTgnxwdDWDSEO9e
Ne+MRn1BXiCINcLfSTmEhliBLw54qncrB5QZ3Rxd7zynn7zrYamDcgGMWG7upN3j
C3A0BlLdQre5gtDMlUZWiudvV58Uos3TAWxUMjo9GtsdShsP2KSRbCuUzDIyxfwQ
eeTz+NSnwfiaURuQnchdrjGWcjuPHDjLW4Y19Fq8XmzRm9yGD3/VE6Inyvp7kelf
ur4ujFKJzMXYF6BztfJPiJZ1+9kye1dAVdFW3y1pMkBzlhCmWyi42Z9PEEpdH23h
0pwAKy2h6op1M0XSgtWf4zwlbRkRjmWbxMPW/JcUgR8xQ4l8/zAsncuZHvxuXZ6Y
py7ix941qA6dH9Nf9CxXmLqj/mrkRTcOUK3yN/GpLn4Lp9kkIV0DBcZVdv6heD75
n73hjfvz7ZCWUR4+1RP8hN23R95Ibxx8fM7W8jEJ8vEBr7KS5MeTH4wvP1U3ITYT
mlUaz5AsTxkzc0j4fwqhERxc2o9TqCc9c8WYVA6TNHEf8QSjOP7suK2eo8WIwCWU
IDRSo/J+nP/qd2Sgwe47OVIKzeySQbJ13Vptqp5Tw8h6YXm+/3iumwdFSF0dU/v4
tJIOKOnGBTWmWqutS4JzgXytf4ef6aIY/L4SDUcnJutbi67Lr4sWC7AVUUyy+5fS
Lt3v7NgJ6fhVIs5nHf6tsi1iB1lOOvK9bNWiBVzZx9hdzS84dSMSlRgYrmCWFEDN
lF0ADlmmi5L4dF04FsVTcEoATPRsZraLA5oZ8kU/ndDTRRHBnVMoGHWRoXKxnksa
9sSM6RWc5s4HMXmiiL3vszu/bh26+yxMMiu12r3Q7XWFQ5T+NIOkesMuGEBHi+kx
kkSGivSzlDki1n5caeTPwuJPfwcJVOcZJ/j1khTl/5YakoohpIwcDpcyzmICEoH7
+fjMwc7xA9GFd0984tK8FmPs4+NdQuhKUS90uqNeC9ficFsZBXMsGaV52aCgp4Uq
2odynGUO+9Ey/UcwVPYw5njNFr53jCmL8CR8C8EK+x9yFQKBKTZWsccG7iMmN6VU
6FIywxqRehWjcQW18tcx9BEJmJC88OyUTCmrg7dVsmWM7n4kx6r2M3feISIWgSyT
8ws/LUkRbXS3kZz8gfRxKjXqtLVCKOWIEE+gAhmywGr7j2MsExT8gc/8O7P4XVpK
7vwFIMO5WE1J+s39k5azdcUKtbHkvWgDEuwUu31pYMNdG48KcOQaikDBaZBdcOEJ
CVN8gsTwWuNx90Cwtp7w+r9cXhCf8X5AqpuTYA9j+nLoNkobgvuZqnP+VEhlv5Yk
fm+zLWwquLmd3kZ3VVc8Wo6iK8oWNQW/57wOE1nthetht0gX/YC1FOqdv+iliNCP
VoV7TKKizPalNV5PKI77WrNwBUdPDnAuW1C1TjmZ/XE6+RuHbf/AF74T2bj4fZP/
SwKtnY70DrCaZxKjaUj3AmWBkWWF3AUMP0dgxUJ4/0/nWZT7tRe/GQiDxpD5+Bxj
wXgb8y46FXGhmTMr4ndWhxw9To416gbGB7FXhvGpkDHVLU+bTHp+66JQ44eyP7Gk
0IR+fdcSrM8v9K+uk3DThQum1NSeKwNJeHpHjmaYNQZFafHpBag9py47X3QFRSoh
fyjkpE+9rbnBA9/WkHXry1sh4vTYztDaaZx7A5tTp6N8iOozNoFmlwsSR+bb211M
ohWv5QLkE7GyCQF4o8t0mYQ5xbNX2hhJpwGLqLq0AMT/BxLmQ9dHa17YNKeEOOGj
0euCvVGperkTxo4MFuCREv8vJjAznJAr0zxN3x2H2A2zjp9EBcLqS6E7K2pdAkzT
qbxQVx/CEuGAeAZYG4UUq1A0wrqa/u1eCs2sm2aUTdKJainjM4ADjcdqxRmsrTbf
2iet2Z8HcxE2ZK/9m1k88fHDYvgqMcaLrA7++lCg02MFnsMXPhTVgIb7D3pHmc0K
Aj7tTpMa1sfPYT0BUfCtqj0FcoMtB9LbmryqeCXnyWsjVfDBKBk/lNwlAIF+wMP5
Ne7PemyT+BYN5/lXqLVXB2pcOk5E0r3S+KejEZALWKriWbDebmRO26nC2qYvgI+9
JslOhHZ92iDxTT0NOrCVutSJE3CNZibazvz0g0tN5TbdZwJo7sEPOaKH2dgh6L8c
RfELuSQaE/oHh4ksV2D7lYPqo/4vqJ3NVXug7h5J+aJJPZ6IhyFAFfd62vS+hkqx
mg+I6oQzQSF3bZNiT6XP7GCZtWVEY73vT0HZmfq4PwS57630I9+SRdu5UzFpp2/d
u2poEfEM1ozv1Xf4Qi4iJGOcuGim38cWf3siyqf3QCZeU14sUfQukPMxo5Jwp9w1
zqQUKI2t+h6BG99Uc7L4NNeI5aGkzP3IWHrbtheqqahOix3irA221DTyHHdkuRQf
eDAPR0NnYApDWOHeqvfQSHPX58MnDWOrULKx7+NOwafzspt7OZlVvs1Sw7CQ6wX2
kEnjZHC+81Avwa3eV6olgOkhg6gB4QnRgC2lNqRxe5L1v4JWF/Uvfi/QHM44uKKx
yN0NQ/LesrAPZxMyD/zb/pGXeHaQ5/IRgwp2QfsWGZiwHq89Eij59mEtLG4KiGhH
53SvjzkdqsNHiIRxDg/g7mptKt44KAX6dX6gc4Ba6ohllW49R8OmcXWaTlCU1Hxj
Z5xlSq4ihzCioD1x0nqGCzaWR65Dzcn7PKltlRFEOgVvmAFX5I4ecS+snkljTxhY
AKezTG15+1dfnJPO0wxg7aJh9DDA6/3Wjgy4T4BXHv4q1hJQQv+7yM4UaVwB6QP4
l8Brc1IWs/lgkNKStcoVcB4J3dfkGiOjoEQF69WZ5Ii+FmGHC5WE4fJKWBG+CS5M
QMQfIRhY5vRBwU35s4ngzKtTEWm/qZ50dksb6KjuDP/Yg6TTuzBbEQ1jM11zG6K3
4BEWLu72BYfrz1W9XzYPjw0h+FvoxxHmpPTA1LwiQkb2I7D68ztDy5LqMioIKvE+
uI6Ct7JWgRDBRN2Ct6v/lgC1WeWI2oO6hYyMewTsU36fDXxsqcJHJURWHuYJK/vl
yxzHCejFfXjp+TZo8TIqsmu5zrKfjZUCfyXvAhSYiOcuUDHhg5ny1Hc2MjUdaMx3
SB0FQ6wYafC8yqLDsCCV/1tLIZLA5ecGzvHD2FvwGr/e8LMWRi0y+RJaEGqxMMls
n/KrBf29SQpYzVcKSjrlVG49DkQm4vPUmj2PAzDL6t1KsCRFeZvRFUz1d8wZZ8SF
OGrNLKRj44tc+lhps4lHtU25SV6YaFdhiADD4DH9MVfiXaaC6ZHfDNvr0J8KZbiz
KGKi2sfnyp5M0qkH4UtkjM/8DixRYcQMuHZ3Dmd2UOSGNcoH1mrm8ZH0ovLH9E36
CNUG1iBMN4EcbfaDLNk/lf/WJ4/TMuDVtmvxuuMkRkRdtc587PvIeYDsiU3C1Bt3
wMaobNE2ND1S+RBLD/10OxqbdMU88kQ3QVyXJasqFKRXQ/IFanlW1kQlf1lW4gc6
jEo9phMGQjZ8aHxHG5hDZdPitESDQf8JPHKc5PeO3pZMZdY19T3VK2jhOsfVqk4S
Sy/cDvlDNx0+1p5V3ciZwlrxXMM5jyPCeLQEeoQ5+tdimp1pTZWhufK/LGiEUxK5
K+nZl1uP1V6hJ6XGpA8Co+Xz52LIr42PkkuUYFaJTn2c/kzYsmglYczHpDnZAqLl
9dC1wzvCYgfgUFS9sm3JJhDRXeEkq8Qn1tXnS9c2wMqS1HFmtfsfxRjObQD0gc+D
57ochSdbiS/vYVckfJO72mK1ddByMoYyYaqC4BC0p9YgaxVD5TZr8o5qKMUbAxF2
wEAb1VqxhtjVzci+daAmRqiKGHi7CjNtSzvA/uRfPDRkh1HNr4O78U1umndS+JkE
ql5jI3MogmMdL9eC4rN/v4f0niZgoR/lOOStfGCWxy339bMKohC9uS7cP/Iast5P
eboWOhgWqReDHabXQJ89VQp6tJyvdWyBoxaQ4KtL+YIgyjnzZpk0c3Q3B/R8dmE6
9tpxkgJeJi2vFKBfI8nMgSD/Sv8FddIiWFygaCPmIdDpl6x+ku8uPWQvf6Xq6bK5
0UW53+oKXXbwJ5tzN2gYdkJLfXFfZWuvdpgkDcvyXuRl2Tq9yOTUSoyG5lcfqf/e
+lWtSuIROdqJ0FBOa2hyw0Z8xCVs3wqC4OS1AyiWkvrDw4KwWi+bDwfNOHleDeWb
gxQa2oFOyztveSZfUeBps2PLyKPwRlQJytAxIGuoCsMagQk3zVNBCsnoPCTs0ZNz
TywcBnRiriXKdhz/ABVHCBnWsZyv3xp0HPKuVChM8oDAQJVH592xbo3zmE40IxWy
ECr/Yb/cW65rgsPwyfxB9WW8ms4Jo4ofbeOQ1PqdWe3/3HnHxg96WzO4PmzzRjmL
NuWyFk/wmQ6YXv/X3S/9huQyD6S+Cm0E1Y1L3zgWxE1Pp1veUMT3nNzdLrhRu/ih
qqzCxQ153w5552qCQcnYNdtX/vel8xzqldU3PgohJVa30msgN048BwbJifhO/ZJk
YLtxPZr6+P3Ra3GKp8adm52oIwehJooHU5G4y/QAgRIl+Z6psRoZrU+pG8Myot5c
4p+UTMfZyRptJZy9H0QmGKGUq939oJDBWe1Wimu3uT9LnVoHjjzk9jZBHtLfYnOD
433KOZ4hj0uvuadHLbU1xZol9sd2yS/RVMWyB0L30Ryp1G8g/V5QiijgcnYWWa9T
vB6dHiJxOwiWE2eo/HGZ8cN67YkNqBdIaPenFG77EKlxN/M61hengO5KjZVkP1s4
GOVOd1i+Xcoz9QeE5OhgJurY7zeLxHJSbKCSRYDW0X8hsXyQFDrhe8dlq7/ZnDwu
N+r0Yb2C8uH2gqxX1pNxs/EtgJecB8V81z/L5kLtbWBN/3f+NMZim+wJckzW1em2
lifJiFwHmmgc+GLf33tAH0c5Tza/A4Ro9Z4KHnx59jz37rFpy4ke7A+H6yom3ntA
4tVvCl2Z7iftnLyieZJTS6iQWNEdr4DR+kpTLqsqQrYqX6cARFbJzKqpuRF5Q1JK
G0V19a6DxL4jXNlbnGeSl1FMV1tA4DGUmLCxytvaw9hedTIdU1zzOtR6fcITDf3G
uO9MHRSW89U8NFNNlr0BHiiCV9YvA4fnmPII4ftbDXA048eY0ylR60LPW8eb3WHb
jLIQGGPN4yxANP/KynFeqwdkK0+T2VyGxgzuOag/ALJlmCZTxkPmTlHO1ckmV6uJ
qNSbL57o65xNABwNTwOca9c3HvxmRyc9YRrooYGx8uUyyCE7eW9g+GjoUgz40tlr
yHFZFztPorFfH6k6GHL1qsIk9sk192k1EJrZLL3A6up+GoZo1pyls4SaEyDKPj4/
kDhrJogCRXjIDTN31kitvtzzWjiv6euEBEuB0NQ1Ij4c+0k7io3rrb/LMh0351hV
wNf4lkZTCLrvrGmdy9j8+3GqZY4ZzMg931YVMZQv9NR9t2togWvGUqudIWGn2WtK
HOWR+S+A+3dcHopohgzlJSsZe1r/r7KtCskt0GRI0Kk/1CY43nEEHX7v7dj73u1/
Yn+DLo/8RqsSkagC1RxehHMVpcjf3eqUCHFUDDfOU1OeKxLILiysdGHhomNNMzfT
YmM7y6iEB/HU303qzjyDVnuTqn22oIBoXw5rIcKdw/m/2IPiH94iLke0WN0wzl/h
gaZN1wDqIY7oLHz9RN5r4EromLKmF3bNSTyGDZpQn/Qh0psvN88NucvT2pk+lvia
ie0bDrYuhVm6TGBFL+0ljOFGs0+0/ZOx0eCLPK0jj+MqDZv0binvwt5p+SNMCeEd
sO//6Le/c6caKW331NOoLaMNaiBfulzZYCai3FLGABcCEPNJXw7hQhPfmEOhYncM
T5LMdsEOV59XAS7J3KRhXpjp8tGItYdj3WoFIz4E7p9hdqQt2RZV7ULq5Szh5QFv
jS8vmKY9/n1qSks6v7TJT26sOC9RbeyrvmVSEzHxQwi6jMs8T/HRUrAgy5GXMuB5
ORoEK77WifKaRDrZt9BdlRojKNHbdSBtUv2LPVyFZ5MhbPd/g3G7K/K2z4jbKDd2
8+ZICnTmBVeJBa/hgBlRFxUrE8b0nigx2WajTdeqesPzo0WIKLRPCPJoLMI79zcC
G6nBryh0j0fyz0vGjSlYKyraE2Kjupu93JzoAIBjmoTAC91Uyosgdiv0S/JAd9ez
EQl50T+UmSj0V1t91zIS7vRuEIruKZ/BOYZGtwAHpX8kSGZzqdDgduIooBUThi+B
60Um7zDE+ZO8BXl7BBYrcoRZbYFbz5FS6n5Hwd3u0e1smv7e+neNo+FDFR/YD8Ho
VPXmGEneRRLU8jqJaI0cRif5vSgmGwz/FiIbbQRhRx+QpdieogbLBeSjue4i5Lj5
FUDO6HI/zAZTftHiZIUZvw6WPSuc9Lr4qo8rwwKuNuEFhcuzCm85JLaHl5CN2WZe
4ibJwHqNsSa+63GOuOG5xoIACNH5nenw3lhiObg+ItdCxt2VEbKoTZqAOO6QFHuD
IRsD/Al7xWXS6N1Rx1yV4nOX7kc5dxV5EsncgHNSa1xK1bheq6Q4lcURwSm3IKEt
KLplijYe+A//GpfckcUC1KAdedUpVfAp+4U2QTN+Cj8ZVT1xyVJGcPqibD0A91kA
jfiaH+xfxkUbIxL36HYWqjoccgFER7xrnkUds5kZyofU3aGFFogF4HvYZdJZ1LGR
fDwbLZWWEctb2X8heoKbOKTY/wPjwkK5fi7o/3ixGSyrMc3iGTsinbFlHRXomLT5
HnzU1KKq4Jy1e0jNfNZyqFCpUPAHZdVm5slN7dT9FFIJnyoc7zmApoGxK48McvSd
foa2ToObbygnVMZbduIEoJp6QK9NXE+Q28AWWACoEqbW1qApyTW/tSFz6yrv34IQ
IXJ2CboSjCzWjzOQtV6VUMCniMpUSIsjd0l1Hew8FYWTu2+X6gY6vDsRnmsafavq
FlYdf25/v6VWg4U+dKDQTXB1A9kElEoF9+TW5BvGudtqkxBj40OSv/MBAIfw0Sts
mMY+/JiXl61rSGfjIvPSphdN96t07fgXoaEv9ud8WHBwbeg6nV+zZSCmuJ1XaGK6
+M8z9rPbqe4L3tc74GLSIQthKvrGFhnIEMoII77OeLNFLtG4BhMfrgzdsCwgiM5c
4Y29e2vs2D/Nxi6DhM7eNd3r24oNZs2wSimsyFAj+qUSq86g2ZYH6GWPN6wcVEZk
Xm/DySUxhLtYVg2iw6MOM9r/IYxa06cvQNlEz+dLDbHN6Ohdd1xd96ZlWJATHl5U
abJcnypeQBLPpXtxPpkjhGmBAJBvCpQAYA8BW4FYLah+rtlbCH+E5K/NXrexv91L
iKq7eKh6YBjHK+GnOfNefgYqSIm9IHGZn85AR6gpO+O2GQk+nH8GtiZSIM+DYTJQ
ln00L9SK6LUgcqVnwzexzMCvgESemLyMrjeKoZ/cObgjnrtp8tEri5NfeKaJi/92
vnts/1YBTpSMWJN46Fzc1tVfkc+Ndz94IG29ffTZwuUZI+UPqAZ//6tzKyNnWkjN
GSIlw3XFLcX4qm6pJ+nEe9AXMWaEYsno3RP92h4Qdmn7OKyVZx3NCSUQyihxHbAj
O6v7g3Fi0VLqCftjb4GJFmeXb26vPncMFP1sIBxmfXzTpw6ZXvWmVuIZjkIKieDB
TDkf6zeGaTAKFW0uajfHORMtzM/3/UH3yORAhUH1QiRiTMBptjSh8YQVaXqjAfpB
A64d+Yu8KzIS30jakJI2i9uzFCG8pFYBvjMPIwKPjqDIA5sGpFlvhJ/Jq3qZa9Hs
6WjKbAgpJWxtwZGbEFvlQ3P5tjTRrAOINU4I5UhE1Cz6EwHhQLQquQT5v8bkdIgk
C2qCjqRzhZADMp/jzG+TymPsbFiPuapzjHrCvpfppzjSGkbOxCz20X2FFUYPkiXQ
vUAq5ktm3QJfQ9P4UnLxIgIyodPB+O2kdU4IBSsjlpjzY32sK9XKRsiwEhZDZYUX
/AbDNNIJZGkpjKSwBJHwNH/peV490LPPV/ohoOclN6xGLsnvVfTfheaovbKabBU3
krphEMc+sjnwdjFJ1KLHUAF15F8XPMtYFbO/XHxXNfuO3jDRCJdLgq185V+UQln0
fIgomRtfiGWUuTZnJgZYYL9Vx0sAVtLwVnSe8tcBC5dNkA9FxU8ofuDq7Q4klniO
DfB8bE6EZChbW4zrKf9nuXd/tGELuSF0gBdjrF1hYgWET7LXI1YNQP/O5DmViWEd
rookp372/NygiU8G54dd9rtQPKOy0TrSK5jUawSasjQMe8NsEDraM70A8mNNQIIC
iqOvv4UWCBtjoz4IZILQ46N4Ooxmd7uMt4PlYFXe/DEcjeY9JmgjEV5amAsMifcQ
TyboMhq64+docM6WyIkAmuaYdhw0RZtowV6OZg9pAnWRX5vT1TryK8HWfIX0U2zy
n+/TAd2Z6fRYcDOJyEmMM8Dx2JP5v0I1dWn1xCtXm1j+lKFFyirIqKbfK4V7H4hQ
pq6QxJubR/sHEBwIfkNq9c5xT47hfaVrTXhRjaANRzQ2wy4bAQYmbXQl0QU/97TU
HliGhvFBx4Rwog3Y3pmQQDMNoCFqqOrgD4i5BI6iwXry+TAFaJGcX68LhSTg0WGs
aL48N2oN4vqVopR1hE0QEmDb/89IYV9Hg/sQ7sCO5PyZFuaXOVyBohwII9v4C6fm
RQmF3xQD9Znc9ZYZjNJtrVUdKGrJP4Gl9ar7Wt2QDzVOUOgDra7Ds3Po8uxwLr7f
S1YWODF+Z3DmeTg060uiihg80SPFfTH2EguYh0YuEPs/QnmGuYqw+esHxJFA1eS5
5msozjgUwOj3ElR3CQJOvp/4BlIm921k1lfgbks1+06I0MELWg/DauLbhc8yroyz
LxW24eFv8/alSlnn8bwZBre+eAzTd5sWeWYcSlDX0PxCjfbrZFfY/Xwt536BIRGL
22gkDg7FkE5DwhZ7hcXjyi5dSKQ7yYPp3nZGQxqfpC09B3pS3C7F6CclkyaCbYBs
gZiyQ12TebZNF6O7+waUmYmJPQeeQmmXmVuJpxnoRBnAdwf9BWlTgbPRCkp9qz3s
jM79S/KHz4gxJB/t6n4QkIRwKjZ4vEBQPI0Q6DuagBnvLUFA7HUHMkSa5olVVAIk
S2Irbojai1kBUuTeLHh0Ehr9zOjVgcaBUcZneIlxUcR6524aUD9qKLdSFAL5lsps
TllUw1CBfDLABHk+i07LEOpwrqEfp+xn1AkJLuuUKbvmnlv2y9p92N2yUkb0OXDQ
ihWUbw4DoXFue52JTSosXM07lzIfc6qIo8d24FwBWrAjX1X/f63f9j+ckD2db9Hy
0vyM6PJFfLKXc4UANLqTeOEIam8YcHUI0ARuB7NN9aqM3t3+gvaKjVZg374dMMn8
E46jNMZ2L6A3od7P52QA/E1S0w2XbN/Jo8QeCQT+tKTus8qvKQKo3imAvGYxNLeU
+JXgrShZN5Vemagy3NPMMZt9cTC09Y9OLhOAicDR9qnu5yM49pwTmKTJODV4eZGc
YBdCTJo5OWXVegBrHR+uwslzWMuspsC1Y81gHfuiQIbkbNaAOiO4+kTV2aI1hKoW
LWfX1dBcTkesgzvP/+NjhZ9PjJQYQBHp2UJ1RRSKGTU9F6vk2QAQ2dg4oOPmqr+L
AEtXLqay+EPYhmHjKKzlTZl9RgmQ38flc52IEEnMqWrG36qJ9FIUBEY1y2kAnDYW
EBHgQ53yuNdhFnnaxT90CPFvD19JNnhL90KnQrLpVff8ZXxvNt9EAwgrtpMYD+oT
nMEtetaNrBO4wIzcWXeIaOsCjmmzp6iG9nUAKhsTzChMRNZHCn8oaM+bBBwtjamc
0UMksoCpuoxWRrBCypR2095K3UO9zg9UjbtMP/vQGBr7qY5XkLOk9FaepFrnv5vn
8NFk9qdlZV0GxKU96Kr7zN3tznEbyUsWbLW95e1DrOfiOI1Tx4Z0oa39jO1EHQIW
UKk+7XrT0U2szINtJ3DpVjPxO3FiA8xn+XUtne5yhDgT4b+1XBRsMZqOm+bZvQli
aensMzwqC5M7bRkJdErOe9Cdzes5EdpMsdBLyo0ysZB6rAocp5F6GrrKwqSWrVxG
vQjKPor/79kI27d4PMn1llbjlF+1ntNRFKNMhsYGjVtD4vbsToVqjxw+c5gCQEyB
RtI2v098B2iNDto0pOhywUL4rNHwlXfh7aRwfY0hlQ4AKBou5GBlAxAtSPN1u4GC
xfghhCaDrO2mNqggnVRTYfsD89OHw12cSIZ/CDEysPrvuUs27gGBf+W4gQxrwGOP
7D2cP8Y9g4zH7fpu7YanAcaffe61YIsxbNFKzZmGFuG5Qi1uqZ2H4z3GU5jG8l0k
qyh1gNqOVPmoXNInrXT0KhF2taLYqZQWc3aWMcBM60NKQag1Iwi2C/jdETz0hcOm
9UA8gSL9QTgEUNNCK7dJa9M2CwDWT27+gBMB8932xfjOMAtSF0ZxkO/CNcRsX5eG
NoN3Y4v3bNSNAeEZHqPjosnU+52RwyHJdmGYx+3eFU5gTXe8/ethJrKPw9LQq6et
7JHsMMVovthOz+/dg6O/fJtFjIErndpft0idOkv6iO8SsGthqX7gZg2EHWl207Q0
irUZK8qDhbmFbaDd9sn5xmVg0Z2tOT9Frd7ZwQUBNd9Pagr31OKA6ZfiQRuVgtRq
i+vSxq24jCqS9mIlPyw4MRzPhzchZuPBySvj9yUhVUTrM+CqL/+KdGYaFhfXH/EP
Oy+BmEVHQgQv34NuJzCKKCtRIE0Bc/nVKzBbRTFhvigsZV1ASzyQBWraBWjSQWM5
C0FgHFGNNSIpp7YZ6ddkXr2eqoMtHpYp4IjADtc/lnjMSTYWT+oTW5/t7jUoHSTq
OJUXTErYB2zM7M/IlH+rb/LMgY7lnDIs0E0SbCAEb0/Qmy9Pk7FfYCWCdPFwtJRa
Raf0e5uPJWjfkcDEnNBdV6ceQgQ1bCqPd389JohngWcfVYeEIHvi55Rk8XnIyStU
QYC35ysueH7hSyCJETYlEh3/GsnNsJ99ao7kdVvRL3m/kSVghiGEv1Hi/m3lQlI8
ZRog11XUWSVecwNPScsEq6rEtIi81KcdgaZKLOvV0M09pLGlCAaqZ4Fs8sPKdRXZ
te+SGgn7Xpe7q7umOk54NikokGgiDr0FxqixLYa8vI3RbJesrU3mjE7PP4YZaWES
93iAfPRgiF0f7OdXFk51u+A7nyol5JdA1mUd/hT4bQqrjDaSHVqmhnB/BfU/VcrE
vROHJIt1hqcrRiVrYXM2/CbHCFleb3B1vd5Xl+VVgQG6NYpknfJR8tD7f7BkTTL3
t8CzuM78RyB5jKhL32IyxOGRNDeey5T3lOya9JPwjaZ00VaxwGBZPgvM85TMHptf
+6fyNHNsTwtAHKHw/rvhjjoVUBDpwr27D2oz4RNOe3WNskjKip6Nn+tmOaZ7O9En
4i+STZyrWBYZR8Nj8eBxcRoLcpzLaX70QHcL7g4kPiThUft9qEigkedQ4y7CD1GE
rj7t/UB0FSCnLko2vG4RiA3yh2vKuNzrI/ZxG8S6ZQfVEa5m0qPQKBXn60GJb0GA
aGo56vJbzEDrZRU5++J53s63rH0o86MoTlNJAHD8MRpgKCwxoY2G1jI23UdtNvuk
KWnQ4u0BMmDRhUi4EJkhIzL8eSGjZRUJr4XFj5hs4KstMwVtkdYLTq8gi3YHOfCd
FBlRy/4id1oeo0N7CS5YWQ6j6/8ymamERAX0nz1aS8bWmQZgvGaOKzx7+UH0co3v
1QI7mHzXccbA0j5gvzH0W+VYG8VSmPJphHjZHmM7TmEoiOCd55HOE3t1eGl9omXY
Vxbk4nx5Fxi1sZAD34Xdf0k4toq2DZif9TMkhu4hvxPmzDg9CG74PmLCT8da32eT
cvNchUeo5Y1stglS6Mybg4XQb1UyCttkR7IUpRULjtBIrPFk3nWK2VfkAz5XCFhu
yzjdYPD3fl7hp/9N52JOjMrsTKrp3Ms20RWmZpsMef9PrT7JMv7WwjBTaZhKbKMo
5pLHHb0sUCS3on+HF18GoV4I8gwCJ+wPcJOisAR757srZRNAoO45t4PcU0YNX4F6
T1bjWUlZgy2npYKdSIr+J17hDomw2EXYL/Ggbw7l1wbRJe51OSYyZ+P+cvK1oNiP
No4JdmZj42VeTAYjJe2kwhVRjOZlqhtXeg5VlZoOZfpgCrNXiqZULgQNOu1a+E2V
Kt+uqaI3Oy4lI1cTV3DMSxF9adJGzUEjec3TFPBTbKt4tl6tCOJK+CuXRtPLqkYg
NMVcyVQicaHC35kGRFlDiiXkM/HhznvrKaTqx5gRkUnkmgX/hbTxr5F3x0AxJih6
Ybjf2zOJ9G9VwiJ4fJqvV+XbHdCjYodt8L0V+9VC3du/6MjUEmn/LqxgydF+4vMG
HrR+P5FVTFWh/weEYboCCE1Y2u/a3snq2X564z4J5vlRGqx944xK8dojHVg+VQZB
XgsBWYORAiNDJshMpGFBnjd7KYQlEogIcOjIzS2U2NpZ5Pp0ZcVsVd2aizAzg2m0
0Nz/pcxDg6ayM5tEW05WEb2mI3TLKd7nPhW4oJZdssVrdGaqN2B6jdlDjJQoE56Z
XxPQdy1XhUzC4xZeqMyphs33LnCf809mPcvP1aORrAgb9/a6/dofrdQlI/iRolCx
0S9KnEf2fY9LRlBCedx+vv7pZmftmD7igR7cVvLdUpyJt5ckJR5BLGcs7ihFlvGJ
ZC8lvjW8Ti0FLYkSpAG+Ek/5pKNiV9USrgWhyAvm7E4PvWOd6GQ91jipz+8IjVoL
a/pm1L8DsNir/exoV7YGWqiAlouKVZ62+ZlXS2mR+cevaGxQLNVUZUr8rXi0LbQs
AZmqhx6agnR7P0KUaXdLHdDpnRvSgL52NGl5gfXrAEaWQcpPskPc+/tlnEN4z9LP
qFftQ3rTzFXtcQrNP3Pufe6995Xx7ye8tnU1DeWne7IlrleFrGw3mIbsxsreW7uT
sHMp8amiMJMEIkDdN0H9JQVLSKzUyNi2El/tHTRhcm3/0V50ZTuagp6yfQfbfnXT
ZLvaotxDzmADixnQ7LsEggbb+F6PKH9tpDENYkzEHHq8VIbARb37VYb497SrnQwB
4c4xc4SYFhxbTrpfLFgndFmCP3bn2LJ7SuIQFsv+Sku9RNP9M4KBaZ0mYF5Sqkdl
LxgMaAVZ+gPrMJGwJkPJ/o4gNFgcDwkLrY4WzPuJR3y2c2hnoSJ5LnFszNXI6AHi
g3KEe2a/GgweVWFnAEl2/aDjEMoK/6/aBBT5VYsXsz1AXmiouuMYvSbOY2e4GjU9
k6UnJLJtQ9sbFXtqKzW52g2qVDV99xfmyB4VYFc9pavRJ2viwj+0JMEtq35I8OM0
cqyC84ZvupzsTxIdMmLSpLr4oNwJ809dgJ05LnwsmffSDgOMG3q2m3fRBY48WBYm
ZmOCvDwvsW6QAbKENCirf/LwELh/bZaNgtcSlQ4UYgr0O/hvTd/iXhKJs0iMTL5x
r33kNhScO3Na7rJ+YiXHr0RTcVOfUakjL95+lb9GUcqkDl9rtizWWiOcpi3MfIyT
FsvEVDKv1TXNnmC62bBSapcMfsF6LLQ8Wh/lJ4ZqLce95pE8ZE2pqBiuVKTkmJw2
WfSz19tkCqXhqCTEDGh0Dz1MIzajPvxkgZeWJQTD9hvIGBU2Su754wJA7VzQWuSB
fy4RPUxnfAcNCBVsZGP/8AVsZuoOrZ8tebpLK4WYk0kKp7kTsdoO3vYhAiBMuawK
4riCKCMVOkR9n81tztmVtM5OGe8RoiWlMax4A3hPY8IsSYE+vq0UK+Q2ZDSO54No
lE64F/rxDoiqbTtMbZjGaiHIn0pAPCJcQxO8x2WDLT9ddt0SxQoT5qlDQQmRnHiH
Yz2QA5nMRpg4vPDHJo0Hq3UeczWsUz7wYsPqlQqhy89hPGeFc8Av5koXpWtEwMvd
oW4jhlNvrEQN5KDGTSqn4UIQEqFzcjwZ1uCf40Stcv+I1AXxzUkFtD4wqg7iosy8
vxub6IEv9KQcHCpa5hvUEx6j2Xf67zo462twoqSxZl3Z5D9ZWhFIigwWtgJAS9kM
ftpAcBVfa2SIvKJEN6Hd1jj3fn9Cii7n5MEA+tn4kxflP8KskTadFUFKFxQoimc0
+yoNAoh2LXD62yqIKFhPMwvHlcD/e7YGAxZy3bCgHZPWj7I6OOijz0Wpt9iEDKBE
i93tgoRkNWRRNOblY4vBbG7T8cXbrwZzfX2Fk4C7cImbb/535+Jrl6CGUpKiZEsJ
XjdTfuw6hV5yoa/IwNe1TKYxEG5r1Mxf03sSHz4GZnDIxxQufHTF6pgXRFZYsN3m
5gldLcCiwcisP9dDa/rWJPHk75nbYz48wXRmU9TUQ1wrtf6AWLC7cR7Pq8P0ubgU
H/C/p0PuOT6H0/xPqxliAoxVospyLNhw40oRgZDWIBCAxObQXAmqYHJcSfeaPf9y
W6b6pjzS0bkb+ATwMUabSjuNkkPyCZV4MBdO42GLGYGhp6xnRQxTUG3YPKX+Jzt2
3vlOeFghM3Ga5Nm7371nMIPnI7Xecc8vei8XDx3Y0ImVaC3xX4EdUFf12qPYx0uC
Edw95Lff0vpYbPuBUowJjJUmNGlcpMWsAhLf3h9YqJmRfnVRfJuojLofujvUgK7c
11GcAHnMmyi33oU5hVmBOfx1CUoq9ncjvDTzAlHlMIXrB+fVmtEDtKch89o7vV6B
XyTptd4svrZj4qlHecRs0+ypVbgNfz3X90X3cX8vfhP071VTz+DbFpEKb2dM/zor
JTlnoBoTGffR9FzRz5GUaKDd4giiAWA+oT5JM/9p/HlHxtDab+QYR00uBVq4ApwB
kZ27miIb6i54SRLoXeK1hP9WyP2k+4YFJCcGCu0Nlzt+5zjZq5UebfvT3iu7NAmP
5XZ9hxYqa/mwKeHlaN27hKsxuxGUNRNbL7dhfcR90MGnps3TFerChyVeUVCJb61N
UqLkPigMiNJ2c2ovY8WkqOR0C3lnR/3rwqwk+b71I6tXJkMtPp8Gm45C+iGuYy7s
u4HWF5Dkpq1F2segNkZt1InWpKUZv8WDY6dPnfsaXVm9cFC1wYRcWsx129L/l+HK
Wsn6ZGbSAP4657buXj42dWbNdVuOdA2/XBXV795kXVW6iPkhWhEvschBIcFlCSSP
4yVP0UmSjXmTj32PHL0kyqPYvC2L+MghdPK3xKJrxjFQE3RBFhf/ZfQ5OmN5w9em
dOujUix9slGR67t9bLzKvxm8fPDnWCS6cXrtowsxNOA+ARGmQ88bXPwbKDG6BdyE
ZsddMzYAPR7+RAeRQaAphatye/UvBHVaEbPtq4dJ2lcCHSRPCYHsbs7mbBUXKQbX
Rz4Kk7LBnAUATvCMPg/I81s17vTQFh1TP4TroU6n061snnoZELh1xLCTcIVBEqdC
59/ojQcSykx7UV7DXtzAFfWNaiN2sqBZH2B2gJKs3pbWn5d5XkUhIMYV36CyvqyG
Hy8irQx90+YYurZT5q0COeEAXRjGeX90a0xCYsQMDe5xSC4ge/4t2jaNTy6N5RwD
eUpc+gyILw8Wf0wNX6cX1dqyWVYpDwF6HsL1DazWdseTX3LRJ3PJIQN9SZsB9VZ1
UGZ/PihR0WHEl1rGpfyEvzlFggtlkxxxAtEnqOcRkvLQ3CNlKYYveoKvPIqEC38r
w91BVDP4CimisiSoobvTlPBgiGJOGYCwc74DZ39a3YY//JgZfmbqMY6MaIMmACq4
la4loRKVSEv59T+LWqchzqFKUaTpa+7ZINoKC0/rifBTVmM7TScAs6lt1mVWqE6W
z9ZKq5MQzNT7zH/ySaaK+Ahec+C9YvT9SXu6qnRAs3m0hVKamF9iFHajMAQrljxO
RwRASia42vPIrrYml+HC/xdWX3iJlurp0zPW8ftfx3Ko0q6fQNYtDzWS333hkNfv
LjIKhVk38wk5zfOoCIpB+zIHs/mdmwa6l/qnfMcxOcyAfPvhvAKKrmZrCgzxyyjg
wxhPgEkoJCq1oDjfwl0GGnDzmV1Pe7gbMaBOptr/ezZRZp5xJUlQuoCk+lXVFmaP
G0mtoHIMaMRIHucqDFswfygYEyqzo1vs5d8ZglQzS4wntsR+FolbtKxk3XJdNNRQ
r1b4i5JgvKNSA0wiubo0OQapHYNfTFwSc8KcFYP/dbTUKJaBxXP0QpfpbvnBMAi9
7FSq/8+7/EDqBmvFNK8Lymdlg1163dys8ckeft91cD5g2yFdR+H2c197pNbrWMK9
jzZ/NcyB+g9AwqSgPCpCsXxhnLgi2Cax4j2o9MG/oNsHmHZIiNmeX7m/Ykj0o+te
kDEXUlZiDDd91XI5C2aRDH69LHuN3SzMvCPfvFN7b0eGmfr3l3H098C7iVCZjMsu
YIecFl5qT5lQU1wNnVjHlwvyBfVaA82OSJJrIe8WWJTE79lgbV15PVJzZ9ZWxvl1
8CLKn04ZNuQSgQMVLa2KQJH2W8+/KTqktnnjHH2pufgE+3iRvWAfdSO+z+RmffY+
bnqWdVC7QDeOiEJtGo6iUKNRh9TU/pWWBfDjPQ8cQ27glEye3SGhGbPdVxNFT8bm
TdIF+CP5Z+Sfo4o7uY7QTMJpua4trEqVXeZrtXcCJrjJMjHvLAD2ZBPwWf9qdRIa
FUTU+8BU/tlAdrsEjUoP8TOxVIY0wGeXZGOCxrFP5POWNPlNsI4IX2ZorQ9mD1UL
A/QAhz+BkWZ+uq8Cgl+dmoXcv38ZNhQ7EYIcEtrWvOf0MaXgxgpN1CBhO1iLw4EG
FQEb7gE9iEXVQhcelN1UMSkzutHUF60RyT5vSANA9E31563UqWJCN4DLpze1z2Aj
1ZvZzodJeNt2zI/zdi6uEGmkBZq46e4OtLBfuL6fYS+q20YadYvjwgS37ZcpZ0vF
vUmXem9dqbM2Y0iCYGGkFgr9Ck/w4Ud6HCxDvhOzrbQe6oVhXYWPtRQgTGvWLj1i
nYFq/O1v2o879UK0TRcL4hqA2z7eqtlEMCBlKSve/g7aEpO/SMLzmwk8fVAVjAIf
TwkCFrleZOb9pEWabAErzmNgOtc/Sb7M0oA3CAJ88xWUApTYWytv8RDPP07pgfjm
lpGMv8cDie15Loz7GLhJbIYleaqSU83pMcNeBvPBvvyyfuNKsNTT44D5p4HezPZr
G4SgSyEXYo8sJTNXypItM23fIagG2o7Yoh4hDhBfRQrHyM3s3pBGbmds7cAnNWxQ
MjKArkQN8rQIxyOjm4m6ov+ZOqSx02ZKwQGvIpx7k45mqBujfXvaCnkdWJtAvlOW
1Gaf1Vd/XxHqFgV+fEIfqlpVnyzWQCMGPLyIjMx3N7fPXbwyvpspMDYSEsUb6jfn
EkEZXgp0nLgk56Zf5N7IHomKoNnCF4mnM2M9mFOBwSvlkvhbzHXAegNQXU8bdaLu
dEXIL9mZmdwpED4zxChp3YNCZq/nyZwnRB9KpsaOteBnwWo5pCTzKl7HbSAFGfe3
wvlyLKoRnHj6KpZKgOHGWbCaKmqv1GB/cTftM4LRLuZRomQoipLNy6g2/9BXfJtn
SIIp/uy25OBWBo33kY28Rx7nlfn7iHxW5GD20hQSa0DSagltd7CeSZCMxw3YK3XR
4W4V/IrU0G4I71W4p83/9JaZ5qdSLMUNNCEvAyOaaGV6C/9tC0G22Txg1xNYTv+r
VL1Tt3tdS5PkIcsx+B0G/qwniVjIc+5InUiWV/DYQUbIUyXcgr75qjpxrTe26W40
fJq4jqC5E3SHb2gMvCSbNPDkCWwQr+PAILSX9VMuvlUOovkWcozPJP6QTVM8qAnM
DHZmJBrYCD+V2/zYBFeoWrcFqS3Nuht9d2UXBKbKzA8WsuXwYqhom1xSGid72sS+
3xGfA9KTAj+62sofF2AG+7m/gheyB/5PG5Mr0GKumLEarrZYo6VEcb7U2CnofCSs
Ox93kYb2A186UG4tAOq2fVDZ9M02qAEbDUFy09AlrGuHMA/hKYU/scvLG3jpnrK/
C7sKL0SAlqBMojR4acX4bYdOzuR+fLCw7CiIbA4cWPG9QdkvXfyqL/eCPGU/0gbx
MXAWwh1kKer13HOI1qqHuiBDqZndSPKKwy/AMeANgIymBJ9h0njTZUszwr8Q5iMy
AbbrDht+lsG9tWEhToXegnzSDbVYO2Hf7gN5+hc2el1UA99IzCTOtkgagXmIj7QZ
SFjv3UU7ESRnsn5Y/DsZ7rVpx2sYVPV64+BmICQDmP9O2aEmXRR6cBA/g4p3gFVR
MoEtywg/pdWpBPhLcL9c1Yge8v0B6UKo8Oz3ujnaCF+oygnTKp2sKOWru/gyprYC
GmIzzWzFvvh/6sUqbvJ+AtQjhPtYQkK143vzuscO5DesiZ6Ah/2wkATdafqiTv1K
l9BAPWHJdfscMkZ3esVuTDRCuGcOf9TN4Yb5lJY70u8fyylzAG9dqrw9ewiYrJMI
8YCfRpRm4n37/ujJTWX9RNH65FUXLKaQWdnlSPedv1x5ZiTKY9jmM0NVyKuJrwcY
KTcHOIMrdrV638gD2VITKfGUaGe03TUN/OiPS+g35To3dLdRY6rw+oPmRZoVex/9
v2x1QaC/mKu/YbtDHHEUYtbTYagAvN04AzkhP2VNGpZz/SmNXc5qgVIdNhSgl4oJ
0G0LShxFbaL4Gwf4nL6Srne9mxfHafeYgqG1OkmvMEPYWc8jANCmKljvC5w9OJru
MMwUbbH+YdvWkZkf4eksARRGD6eE3pgga1Qh6weXSJXX/DOFiSLRJEWSxl9Juyh0
KQKwED9Xs80Wjy27lrY10rTknD3SQkdv/4jdTpWhB8cgCWjgtTOl5AiTSg9is12L
3LfIAR6P5Mh7iBANso/mdZlGv0PxDg7YDhfPkli6RhGnN6gflgjxBSiub+I5t/Ul
znuQjpH2/Ofi1jtZzusgGahHTin66uIlqTkKMgXSmm/No8Qwp/CjW47qOnNW6U/G
bidgq27oMPxXKp2hmPbX3YdWTirNUJu/2bqLCgpcSBhm5Cu5D8S5NVKWzQT+0oli
ovzOE77wvI45JkegXIvSOQ3kVpIhtp9wiY8KdunZnWRfPJNai/fy1nRD6Xoz8L2Z
di7b1WTKQ50ejvWtj8fT4MMCqzY4j50Kq2aTlr1hnOdaLXs2o9Ayq0ulKOB0Wy+n
l8KQL7AucBxqLUgqrdntjmxyNI6OW8yg13ajOeFgSsVNY3i14AbeIxs4omaNjYwL
GRZmfeAMlRp7QABBR8csvbJr3Q/8zpYsT0U18M4SjXZDkV+ooheuB1lTthjSx4N7
XQ4B37BO3TU+PfqhnLJUsk+be8uKl+D0pCDYxbKmgFQzI2tq0KhWCtlORuhfKxs3
fIF6/GIZknnlqZ7a+HS7CksamfjjrawhOnukb4zAZO2qaMekuUSjibHXOgtJxrrO
Z85ut5kWoyTDYOeWPdZKKctiql+YuyP2beC4PtU23NQKdiZWXgYoxm0twFQYcIge
r7SYIJ1OWJcrtJl6j/0TdzW+R0Z6qseJEbjQ/FklBDVaquYwNMpvZAqrgDnl5lJW
KYNjouREH6qJbuz5cTTcg8BsL1TcExQ1IsGOVlF6kdIr/KD/VuUlkjHDZjNi89wO
+Mq3Z+VXaCPgIS/hylgqTRxkkSvbvkNt5ir/ohaBKKg3AEtD3zMPMQcHooqtFYdD
UDQ3fFzozXmhnKyk/FTHPXYj4V3tRUw+FIyq4JJUF/39pysWRXG9jINFpNLMlJKb
3RZP01r5+3Qk2/Jk+hRbRejMXlhPI/GoOkzl5WUQFsrQqU1APpiSSJSAz+ya0j2y
kYVNFNANW25pgHMi3uqO2nZmHywyIWRo+hAww50N5pcXyt6M0agtz7mcwSBk0njz
oIWS6IUVslGP/CsT+cdvT6kaj5ZOIeOxm/Y2oMLBSfNidbnkGTeyJRoUFHzeiIJU
XRCsSA8sZ3MUqEIaW2H+Aqi+xnTqq27NslzpSSUe+KUG0zx9C0BA3GbMy3v58gaG
J2v/PVqoHYRYdSn4d0H8tWDP4IR2UDDgBLvzuBYoEEO4nej1lnV7q/ia8U30zKQl
JYjEQ/FBOdnaHAOwuGMgIDhtZo5zvqK+YVQq5+kKNXSSQdgO+lldkwC1q++9wq8h
AEL011PQOi+22/7ArtVf3gVy6XJPIsfs4DiAx/mrbSja8PDGjXYyHEmS1+gQupGd
Ihn/EZFVD4F+pse/Rofazxj/v7Pob//Xz+or8lHa2LXrh8nFzGbYfGXpUEbReCxn
xBj24xUoC6O1pO4pzqUTTOfD/T6qd8F54yO9Fvrx4F5d0llyfPLGpE4dj3p4sasf
Sv8BB2sHKmXSiqJa+K/Dco83dyYj48RWdB9M4eguLZWVTbyyUJ2FGQm9EM4p3AwC
DKu+trRmpGyr0+cF9lRwx74gICxGc8I4tUdJBgbUKq1kbCmN6UVhiuSC2tFcJG9W
Cv/Wdr2rgGtMMP59OF3iPj9aL5FdtHhCTVUND5wKB7wqdh19A248n9+nSckZ/ite
16iYHaZu3HLl8EmwJDdS7V7jXRl2t64q4MvrWqd46aTvCZLiMmdR+DL6IodTY9jr
RTAlj/cMvRJ7ImQPtgiTlgEvwhHMZnt6jHYXW8XJNQnGjO3eN0bBDsoxdeAXiWjW
HH0vYpX/1mIHi/KQMa9dIVJo2tyTWmV3UItCww0Xfb+XgzS+qikvbEzJvf2Wd8Rb
vlz7Gd9tieQGfmfVu2Xu047SWEyCOJ0yCOngFEb7dGJgONI43sEHNu3ExZaS0Tyv
bCl5YEt+yhBjuxnpMeE+dMVznmOqDrgW3bPWNYZX+uao2OvAxgecu7WYUFtvwY4x
cs2Y+PBJtlpfjUjIEOvnlflszRDS12LSE5z+INzRFFGoPNFUbMw12FbJD9sC6fs9
5zvCgEkyCN8KJY36SRZ49kCdmaDWqAExsTXC9rXe0h96iPlNnY5Ld9vJ+ydS5kTl
zu6+Lc3RWjSB/Foo0kaX9eoUSrHs1wuGWdWIe1astoxh/exen2TqAawCSp1Ccpyg
ktd+FK6PxqaoSJV/tOC1JyEYlUVUKbtOQakC6ES8LxaU/ZVQepcOddRrSJdWqLMK
xXvEHWW8uRGQQZ9499DDxSX4ubAF8DI22/WFEdyDwqcQlsaSc6A1zRGMFH2Bfp+P
XQuELZGr1rrCGg9VY+SO11ZQTabpSL+fj2ZGfCzxFwYmYoZAkzFu8HnX0OPpn+cN
aWBS6fbHoj7Yb6K0iSYX1YnbvED+qV+OdyuVxZOmn5lQSe+Z42Xf122yT0iWULRZ
nAE0ee57qEtv8AIYvFSvfksU8epUZX2dQEHRzybeGZoInK0+HuLXs8p7Ss39tZBc
iJ6u7DyyZeqvY/w8bilwYA9NPnhYeIgrDVePlxoBpjTlvzsKaCg9FAcXspJbhitm
8rSc03d2xzc6/Zkxy8mlvHxw1PmVP293tesfcOEmSIdqmT+Ag7nKR3DNC2PHBYAj
2ZYJsK3ZkTklvIm+k4wOmaIza3GPNuQewxJDZMvHcJHoD7VkE+Go3IEjVGKo8AV8
L/nn7TWxvDV6OTgJ01d8oPU+C5nV5lWGTrTcPcoJoX4dD55qFMdd9GQ1OTzgJg9M
rT9j1gP7wbWaf+faJdWGLJS3njkFJtm57dLfoyyIr3j8M6Munnu4NFDMX0nKvBSc
5uVy+se/MOeK+gfW9zjepceVexUR9K12fD4HgYF6pGBFFwnZh6gFWe4eW8FZjnpj
4UFV3J6RtoXEDLy+jF6/YACIlO4foIz2C5Tfkv7SmOtcEthS8Q15ZDhziyX2yrBL
i7UdebT9JL2AK2IuVnsxekpgkUlwp2FXy1m7nkmvTHvhmLa1khO5bodT1kLnkGYT
k+krXIuSlD4m7NgxA0T8A+bhCInEDAtbUvuz+0Apl7HXeTOk71f2Ufn2cV0NrxbW
M2fT2tjygiVpZ9cQnpjhqnsyGdJxg6K5SvR+TusFcSBn3sbdlR1cJaa2Fs3zsjpb
LwSqgYqjWpvNGI+lZbsR5tddUYEYIPFLR4gc3XpmFIltmXZFmM3X0iH6biT5jqCJ
aYFGFMadD1nICxGuhCfMiDhTtOUXXRZxuT0ET/es9oCwXGqrhPVrqVN27zSV6H4E
nQlD2qfVNo7tWZGtghzMXeP6TXogomSxiMJf86U68nDN2YIsKJG8HcBDvtOHIPvT
2rAfFypuJU9iviECHY8/9U/6hA45Yl5euZzf4NoN00EkQhY3gDPATzxGhX2LorJX
nvmJvZK3K9/XcQbQfCrPbu6p85h3T9ogMD3Bd2RImtEO1DvC2nQkuvGyBLKgxMnh
s1NyaWGoeGz6HcDATiW0quKEvLV5/7UqFGMSudxvHlobYyiozck8IxxJe6TCFYr9
qqHNP9dfh7BzNeXcCkj1Z/az9bM3snoZ9RJrNDDB1L5WAUyLxbgzC/MVcaQRhUmD
71H3fg0pABHANNXoN3XXixPyutwqBr0+xIMvFfmWzuUwR7Wm87G16LaOwNdqxLgY
WzPqp9Oat8uNcvaPIJYbOPvpS21B1Z/KFe/rQ8kNbdKdMibLJlCZrPk7bAVkWhsU
Sa2KTpbDzsLTlgRzoOIpQXRIKwfA8ytqvwBLRv+dGxU6tWlF8BIfJIo2i8LMDqiF
vhXukV5TcEgvJ2K0H3XodXP8bXQl/f8JjeJkwSDeNfNgeR6ovQS0ZGpcZstNGypo
5NDCIuBDln9/hHD7PGJMTYbihy9akMZRmgk5pFzwj0SJ72IYYo2V6bU7uz6/XIHo
fp6XHcosPdwgxXtySaRUP+bPmx92H2rthrRiDiRSSTzH1yy5iXPj+XJSWvwZxkTy
opTJ1m3XRgtINgdvLzLf34t7s+tjksAoKVUgg/Q2UG5wWU0RIYKgrqnqcxe9WjTM
stHXx/JwxsSaUm4qRmRmJOaM182c66l5zm3KfPja72V6Wgs9sbN2EBmXA8OTGd49
Jh6lgU1hm+/PqCNuPeAdC8zHK0T3sCZ3qLJnkN1le9mGdWmib3O0kuEUy2t1e3nD
UImmKWnSDCXNfRd38mJAPF3RfYRGx66Z8oxq8FQo4wrly0MDtJjPtYIp/5y9LS+B
KmfRCKhZS4hCqODd/fv+rk5f+HiclSMaroO3ouQGoKDaEQSvedjxOX19gp3hnl9q
nmq5y8sIeztZGVbAAgws1h+yh3vO8R3qVSaHGSvAg7KD4cmTM2KgiGk2s52W2MRv
gn9IbeH0ExaihBAbAjDxwI6kenSOOvk+lUasn9qCvfMzh8EYfADSJNv1N0psjXRF
UsMhXY55CmRyRzpeC/kK5tAnMB5RrOUmEEZQecqM/CWZnzHomIWr3RO/vyHNhSBJ
rjch+TMx/aKTucOAsq9IDIlMkryhelI3OFcClTWu15ZkEYDBldDj8LgkEhg16Rqa
j3W68FFnj7yImHX1ikZJ21GLuTHW8cXLXsuAY7vfZPIpMVjDz5DTzqq1WvAfvcBG
Kwj0py+CKg3GHkLqo7dISbAzKqJfkTTGp7GM0+bpGejZw0FYRoP+E4vCCNsMoLSx
OgxZCzPYiukhtggBNvV8hXDBj81ZFO9bEcycEAcmIJu/JwZXKu2m3Of0w1E67kX1
BFTrorhNeoV+fOgEVrKt9tEtELuiIncRhjUP3OicWubf6r9tfdhLxJ3FfGTz5q3l
nbQv4jKAhxr9EC3kyz/5iyjtIFeKYCm4pa2iT2mPTjuaBQg8deo5TVlK3y/zQXyh
s4oxpbEaYu+gcIxOvIUVsWbi+2tLDYinMJOogY7+h6Pbx68oJCozdtac1Nlval60
63D0vqLlLjijbUzt3Qwew6pSSOM4mjwsfxgr3QZikaLHN9iuv0TkU+JO83+Wwake
IMt3iOgAFpQu2hEV+NNdmxwN+EW4ndMJWHZQDKVHCfX7Fmn1potAJp0F2W3zQvPS
bvx28VRQ0fH53xth/ZjB498INBxOtfpCYBrmMWjBHo67Z9a26Mk9muBLo88cfZFM
/cu6diEfWVsm9+aoDeA8s6D5hNgXa/MqcHWN043uzSGAbnriB8WmJ6EZmm/yB5Io
TJ0kkR8B55yQIW8z/yairAdnvn2DY8ZyOIgKgtEjLBqBFxmXmVEGhk+qYLsWsFrf
ukZkgXQFzJc69KrXSNljMlcueo2qSR+MWAkK/0qtkj3io2ORNdbIPydAmyCoLYgS
n1e7bwRDHVZK9aYPTKILPot9gjxQmXE5A1Gi/BN5reYVdqxwl+m5vdlVhsWmnWa5
zCqvNtaD+3nzP1SV+XhmmUT/YjGEiL+rm20V2qs3Ck68WVe0a6GDmeQrNAE0HJ0y
iyo2DlNiw+ZxHlyvQu9V+rpp5pwqS0Cp7e0Z/ZWYwO5iah0IHuQREQuD6hokXHDs
tD4pgSjVQ18TdK3jNVV0NM9heWJHnqCRyNHyzmL65I7uqLxbW2LNy1wvQYulVlDa
UTlEfC4QFLy6K+0HFn4+tPbotGw1Mi4rSADzrHExfRQ//QfUZAkm28s/C9N7RCTw
Aq4G3dUXJkJhs1R7yiorz8MRTucVwKGFDwXZlN5AQReHQ7M2TI9/Yz+xmzhO1xYh
ybcqT2Xw5O1n45rMkiXZorAdGVCk3TX0TDxlisd7ryJwpyx51RDkXt6tKih4TVwa
rwh2M9ljD76mAaPdGbm1h52lgVifdWZKoLX+qr42zsIw3FofMiYlFDM7uv+YMp2J
4Oro6YSMab12D/RdrrbCvzPXOhVHupQM/KYP3RZdpk+3FC9EGP+PYfmHN6agkYEy
dsAUFDgd9EsRzqgubmRzvdGHGT0iIpiekDk0TD+gcMTh2R5ADWAPS+W6CLS5P5OX
sGdIg4o/1qCugSDo7DaDXkczJkZTY7oi+/ZlEhIpjlPthMp/3ude+e+1Sej3rnn5
K10nWcYZDtH+hPGOEzn1LyaIYUKXPfzvrP0Q3LaR5/qm9wvF+m2/GaJUoqabjx1z
+WvAOuPSHhlRsio5hLPKN4IfqiIU5A/c1JUs5V1LV0vR9+x0Ra8Rto4+0KWc3XZJ
L6j34ZKgxfy2Hsn1n2ekBIdY3hmVZ1cA1z34HTgPacmZAx6J2BzMzdUDGj1Qg/DQ
rjLWrGXzDZsolzKeFRSUjd9SIbXEvwsAGC4UNz91i9l/b8A1vC8OsuOc5TeHZkP4
2iUkqrLo8CjkzCfk5hhc6+k8EEoUYFwN+44979e9sagDYSi58staLiMmPThelQhY
n1OpYWZuAvncCnOuRNHtLIt949Du5Bdh2aGHrsiETRhkKW7pA0W38Qvy3+7B3Pxs
VM8Cy8w3o630WtdcIhsCdXIjQJwEktViloj7cLM49lPRuxr2LBe7u0pu6mSe2gCr
rINLj1bvkBvi7thlx/By/pgJEhHUcS/G8Br/WXkqUIQJT68vuIullG76bG4y8sbc
z0MrjEwC8oq1OvL9M1guz3eeY3JFCjfrnt/KZ7IY+Yytc3/4gFCyyZJBGZWFuglv
bLPKwAjNPIIsjyzbCF9od4kroylMCY3sj1VI2ZGKblcP8d3Csiv/VReaNjzWwm/k
VQKArgOZZv5i9xj9DA7sOtrzWa/DhF4Jk/tXs6GkJNVChBM1pmU+HOS4k/dkHyxH
R+JsfPJlS7rTit92gDCug1992FDSbJrivmuju/JFme0d7DJxi/udDuhq3RljUpx1
ZHMq5BcKR7f8Nzt/74/jfZmOg2+0NGGlZpQAl7uUEt/vyywjjZnLOCvcO3z7pnpx
6bI1BfrnPJGQBONKkf89AujsbDfjacRYOoT7TvR6Hg41ItjbS1wfQGyEOp6lhFbL
+9UzmjPX3bEbMlF1lp0LK+l3ojJ7FZ9B3ZumLU0Pz28MY2UnBPkASypfmgosLC6D
BvdhA7RPk1OZDeMNV3RULq7nsVFvWZbO1kmkHsvKYHhN1UyNt59mH+Dv1fi+KNzd
d95B+zEyQxUiQKR3QwMv1/Xnw83RXfPwOPKJ7i9g7O5pK1+MoX+W9CgLCXo6CnGe
BxbBqbyNakWKoqvnMHUAnhWCLb1f7a9uARfOgmnmJoJJfpBApA+k+iFUdo5NsroE
FAzrI2Arr5uvrvovVGiOW/5K8oNP7/M70EhqKwKTtnRtPfqaYtiVXZ1IQjwrroO8
nV6QSeJ3rEvzLosX4AHj7loxLEqe0pSBtSNDShoHYqQHFnctEvO28m/hSE78rTud
4fmsD/d/lgGpHI3uqEsFUM4/BA6KMKpe88/KDKWDald7j4E+xWE60ftNfBWsCy1N
n83H9Zxa9F/F4JAp+tMdlh72F8KpqVvNWzRn4REH7VfATZpJkwjGO7QYaR/0PrsL
PGWW0zIGBwZKa7ctVa40r/2UZV1KXWs42Da2J+RJt+cpYhIfBrYQHeKFVcCJwuNo
s+Lnkp2RwzeFHiu1nYFr3ZYDEZ3s+Am9wCBNXYfkD+ddKCm2EVVp+JK7K8XLB11I
8a77M2+AZyFSZFrqeIErlmYABLYqgo/tNg4hAoWAo7Sw0O4UQEQzGWb7kS6uC9iu
PU5akXDd5mV8/dg88Ja6noyQEfTQE96O6WhNwXkZkt60tvOui1ipxSNxBpY+C3No
jxN0Pl4P92oA7S8VB2xJkzSUk4j5+Bhr+gYQSNNvhbNnlNbRC5RHSeyS/djB89t2
+zpOub5yA3Kejek7ne4a3BpMMe8z+i8vTJ+0cK5iOvhzmEZEtUnM7LHee+nn9NqP
DZy3LZdIu/SbQECInWuDZvBXdMhXW5Oefs2e4SMiBJ92gzOP+moDm1DzrHOC9foU
CFxZOT9AhLyeklMgkuelt7yuwucGedD1AHnfNp6sGwQgIcBU/8dUF8NXoZeWG8Zq
bN/gABHc+3YKp1JUML2a9EzWy5lDKuJZFRZpdinuNtuKvYMZH43kSULULXRVLjnx
6AX8rJVRgaVQj6S1OEYuC0YQcCVIzWYj97mc24/JelGNBn25TketRhbhkA5cTbpy
mjYkLF86EuvWSyOY+HZhA9TVMP8RKQs8W562Z8dIaTa+uMCcmllmupLsPQejLEpg
3qVgL/VHoUjyDZfwxU4W029u48/fqU95YSOtx2pTwzeZ/DYl60eRzCq0fdHHy+JW
X71mE1pMRjie2xPPy8kFObQeeOViCTdqLXKzthH7Ob6mcWhccpZpfriakx8CAXge
ySYmkk0+IjgByzDtRdDWQvKkOVkyT38W6qW/7YxVh9d397fKKC0YyDbyPu8CECyF
WbmivfaKiSjXFSIv1RqVo0JiU5X/YpH7ZIt/Ii8wCy36/XIT3OOc/HCs6RVDkoNT
rsTbDCyJca1vHOoePEX9mbbVjyvEfIxOXBx5xAs6nXNTIw+JW73vLf1A5TjTiXv7
LHgLDe4BlzKUCjZCaKvkorxy2XozPGSKeoTuul5vEgD+gZiusjvI2xCE8LZjrQ5n
YJDibg97F4UNZrULEzVeE8Gp2xhEXrlWcG5pqsMRuAQHYmixzgO+HbWm1cX0UD5H
XPjGKO7k57nbt82/4UXgokMeevi/iWLb1xhcneJAagh4IMkbbjxxF0kwJCL23Etg
k6uooVQQaFzYgt9LIqKjRuWbOQ3Kmzp6DRI1Vg4FTOEfKU42S0V+28wiJOlWOgTX
8NHuOvOVFfm3UfVWigkTSTT2QdaRM2T2hYxwX1bB+QtH+RVqUEZzVUFUWvPZK4Fa
LRvEL+m/IQatbVsujUx4ERaPtSSWUgdm1OueZI4hxpI/X+4J/S7tgIh7/LfNin1X
6U4Ff3EtXM66phS2zrl7ohHmjkp6AKV+a0EQzWtYj/zr+jPvM+LvWoUdCvMBkPkR
pTfv4DHRm0NzjMgb0U2XS1Cke7k4jFpxXqeyXOi4jTlYNmPQoVMw1FCDmCAMXkzD
5hPWcKLmogULnfx7L3e9JPEXf/MpMSvMnZLbH8kirXjD4pjSbjuRXxQ6nogh6+LP
e8DDBaUqElUaugmDheTNbTDR67aF+9uEmiklNiFHW0CAHnxaXWEB2KZ9gw7j1P2u
COP3XNJS3nclfKN9V0ztavIMSfWcqqfX6lwo0tyrbLKVOlxVIg6RbggT5T/wbW3R
aPMjk/YGJcq8VZoPDAse3LNYMt2FvYNHzLpkpjBqE0XGJSJ1r6EWkfZMv5IsgyoQ
NJJ856OEIz+eRgP1MFFJ+Nms0glrCfPUZcvDd1ZQP7VroAeugdMheVXHRSj9cSHw
oAe07kp3r63oHc2jVcO0RHPJviAxvl0xUMk81rX6CqATRAcnOPnkM5BU5OTOy29a
o1a1Mqk9+BAa5H+J7PJggWR4d+burxthvgs4oH3zZB7z5XO6iVaqZ94xLBCIvF9h
w7hQ8YHaoQnxnGcG4jHrYujD5aEIbk8WrWqq9q7ivwNkyz9h2ofrrV94FJbmT22d
KH/nAm9+3eyvO8s+afjuG87o4gVz9OtVb9k8s8QN7aj6pafBo3yAaZUqHfkIvm8C
Vku6pet/WfXZ+OaZsqeXI1X6IdKvGpUZbU21swjVOgFZuu1aQNGNyoq6/dxnxXUD
2Wh8o+s3RLyn3ZJWOVzIFM+X3wu3e8t8xasjIiJN/ZW18WaKPq8VeypB72ly4Rts
Sg5E6pnpJD9aB9Ak7mauxflSKeubmMlrNVnDwUQmS/fMHG2vg+k60aYM8k+0MuMt
OQ+g3MUkpEEbKYIzgPeOSsNKy0HoqiUhIVy34UtT8q79d9v1NE9OePsFiFQ8qv+f
h7374jA7v5TPS6w0nlfNjF4pKP7psdUG62lGnz+p/bno0NJz9nOPprLvdmmv1B4z
4xIUHlLEMBh3atmvfQnEpjHD7KpPs8EsVU9aRtOeDRhv1YntjEAJIKDdx795UBCP
xTtJKikCg3bT/j/uqyBkEiNr6wHroOxfLtsaHDCQDak+34aAlkpYzqzp5sJIn2cd
o+F4fyUQeQtmgpQ28mtdq0YVC3+fl6kIVPWRcLVQkiDOdj5LLDNVSeAkj3kUP7s5
n76gEV/J56YY2ZEUkCls7sovuKXKbkOWsJVU0m4RUNlgzpIH1BS8uNQ2GmB0m093
f++B6XGAvobut/cG1ZGsapLk30Vk1OSlgt6hMIuXj8q8+80w0TIpJVvTvD8q3FLh
011hCdc7mUFCuAysU0FleDm1kTVT65uPxDSFfLl+Gyx2PwJutFJkf0pTFi0qrW3k
ESz2KEAeu+1fQqHGkB9j++SGdJhojCvC4V5h04u4d8ikrwEHBTM7QXUBnLuN/ts7
mcwWXWoANkuI23HZc2cIGrTGoxMxukOPRcWtoblVUMS6CDtGDTusSuZm2fUC1Unf
/L85p3UrjGUodmiPasA8/7z4WdexL5XwcGOgcDg5Cc/abJugzzHmICZ9zlW5p+VI
7FG4fYnFgu9/ybYg7ndBdXby2MMpBKOQJJL9skluulvZqTH2bnoRWNh7OKknP9/q
E/Z+kf2aRoUV6IZTFsNl/kgZt6C69wFsfQ+WMjbSouYda8uMsGS3iiz9NI2WhhBS
WxtJJDQRvlJ0BXIWkiYd9KaFlGt/pao12myNVOQJgHf1qWBPqPF6oCSIx1OYp1Fe
Jvgp7sPHuik8prMxPh56eTkphclHmNadw2cEGd9DVsmsVsNKtU2ca3hVL3KvHk1/
u6+nTElOMmtvZHKaQ+D9OVDBvj4DkauWxAOdb6A6mgWb/78U7FwCOGB+81mlR57y
ENpFEF2sWfPgpmWeHdHKLoekDWzonEFAJK3vnhKXAg6h8GDyM+U7yLoI8ATT5hmE
gvtQxx0CvnVwmbbpinUva1OeUdXLJxWiAKzF+NVjZWnOB5BXYpGdHDmdDAdhSEWg
ZGQPPmHlYxce2dxsf72bFVK9hR9NtSTTWZlp9xlKRG4tjqk5QXjhUJY5v5IM++7N
kpydofKTVax/Fpi5w+VC1q519H0KU+at/vwssT/ft04AmkqfSaD75QoNhFiwuSgX
FfoBZFBGY80hF6/p+uoYpm4YLKXSiFXGROstCYcjs07G8m2+mBe2QwOS4qrTkUJA
O0TbLrSAKUd2M+Yfkj6KCWf4cMTZpye/Ps+Tl2u5NxPxt4gsyRKdVQWzfR1lrG9m
MrDI3a1R5OTgCYn+VDzSKLqvg6enZG3KdBQLAqHX+Zn9J6WfCYBlCNQ224vTf3iV
RYDVJzLr340gBLSU2827m8USP/YCLPOhvNssisuESpU7oxFNoDd4LIqm9SbxzWVg
tqgwt/uZwtfPTW4xrx1BLf0O6ebqldwC+J/DODPI15Az0svmS1Nz70E8L8O2yz+O
fKS4EZldoYlI07Mt6/zVkXtw2Z8/7AEhxTB9HjxgCkvPudqhDIRnZXrmTExU8xPa
bGVUtK3ciIbWKy3EGuCOdmC9vIkGrAipsg4hXQNl7Hsg5Kc106ln913ih/fFONxO
YkUELkMycWgEj5DAsf8wAvKd7rVRYsZCrzBdT+mZOMywMdUJiGdkXbib9eh7hOSV
nTp82bOKut7HqcgnIzKXmOk5UGHQEohTgzMI9VYyBRccGcHK8Tln4ymjMRQTi8+r
YJatsXqUZw/zJHDlfCawuhcmx/5r5gUew6YP8xPbddbal0JBlqztrILI1muNlO4F
EH3U/SCKk09r7FUl1k2vRNrW2vIOHfZUp3Gtkat8ZV1JdtlPDcOx3LIzaGYOX83X
lzNwB8w+y9y8V/VyFQwSf+7IYovu2UGZbtSQl66/fiZMeZD9hWRJWzRTlmxRctlQ
kCb3M7vQh7vbw8BEwM+AcK+GZ824eVpJCMSAQWmvMbP1bkiEA+2gAV2yQI5h2zEI
4TN7+qWkKqiqTSEo1al+PKbt5pEFexmgxIYf8B/P7WArr2oEWCiXJWt5VFkKTaI2
+bNSgt0tkt9uI9iUUenpVCJJxzs/07G93ECgpPvcxCav2PVzV8UCfxsQOG4c/zs/
c6EAfyC2nUGFIzqz8LpeWvDChBfsDFLerviZ29cizIDmwlptQrsndV0Fj1bjtBdw
hXRCW5wzYqJMLRiEOzOgqW07q/VueJ9AJoJVFByrJKrTXT6PTlmlllAIxQTjbRPx
9kYmvPUrkNbYe8208fm+0mH7PXKsLEgH7cx3oA8rxAXeqoAeUWWm3Qugh7bSgM+6
6szEgygoMnm5xIi2EtgH9D/RhKUjOpElITSwMSGLeszkBmsFY8wz5I/qtsq/t3u5
Ufr+H8qfgGJSFZkGQHktCay8JAFRP0iG0/3cLwZuTgPJ/zNf4NCtc2OHcXUdT9GI
EbjlMDHxYvC974cuHdQrDsO7Z3/YGWZegpOgP75W6OCFbC/xY1tAxAYGKyCm1hz4
PejEmunh17NXuZydSNheCimvED/n2ESruvF55YCDSLzhk7tlTgH/EN0LxT4QdkFe
X6r3/yvuVGzIuGL6Qx6YUQ5j9SzkfQdhdXZ5qnnrMfCgr1joTu2OuS9MPDnFi+Ll
m6ZoTS6f1Kn0CJb48xxDdaZq8HuE+GRPqB7RJrho4kP73sFI70f/V3tIPu6Rh+Bq
Y3fvUTzVjYFAk7bixGM//IVLW4bUlhNrLI5BG3fLINWTlVbE5liz7Y//Mq7MYosr
0mMp8p7EiEaoYFwEzc3zoLblzF0CWTbuds/eCKuKN/PQpGzO3kbHUwoaKySVMTNF
3Tt+qZpY5GrEKQFMxECy3Y9TOvEJwhcByQZbPV2WYeGYJcjXbw0A6rQ5763DkLhU
zZCyORRtxjcAXUtd5FEJRJONS16L53Iu0K+DOpeEyaYeorzADsPrwPU0KCA/fN59
F0rj/lAHUw8fJlYI1hR4LR34InrVYMWFniDufy7k/9Ut6sp2vhDgcyXIZR+YxOe4
RnmJr9CtOMz7JXCFH7zoKOLLk/xJUIfIs/oXKBBD2HNK9S9PgwwS+u6+ltrgeWwV
GMcQKS5hsXeI0TqNXTkSzlM2c3fqnj7amRtBzrldrhaXttcV5qvttSnh9r9Xb8qF
Wxz2PQUiQHe9F1xwdcaBAyeBRMfkPwNuQqMQAaus3Po0skPtDeSp+jiSjjkhi5Dc
5Nom+04TBy7NtlMLhlFDeRE/YoLt0d4H7QAvdGeZ+8NSFOUIZsSZMk8lJN2LgUJY
N/32gnsLdyN/ghPKJukKbRiUVkWJUwFaTvOkVBRkx9QxlBX1ej1B5VmvkcPhRhij
2OLBvGtmvW1Zm5B60Ol47va69rP3Fn//RDX4fDlW2g9W8FWiWt2PDAvqU/7JJiYe
ZnO8BoX2kwA5gipe4AR40Y+zWhBuaTOQ3SQkAXEafjRXccd2odLG/IXLTuW3AEB9
hG3ce/YJV6r7Grb98S9LmOxfU04CPC3AwUW4/s67L078zqootCSQ2hHsF4ApgWOW
VSL5N79Z2anJFXPA+2MOvF1OPlahLbCIdlsgIEXGvWcblMHQaeFh8EaPx0hKBF5F
Y1e5ivpV5wpJf51/ZL7GjWZ8yGgNfQhg/l/d63MoG++8sAcekJ10uyvIAhnuttYW
zYLNAwa6zYHHrPt5czn4bwf8gUyIM+SaeXL7SYlVOX6i9RPSIpEhC5uFU7jpBftV
OLYUp70XgFD1CaIvv4xKqEHnbM9Zy5DAzDkv1lV8MKVNQEBWYLKE/VZFM3jh3GrZ
JRJaDGOFbmDIzzbYVeS39+taWNJMfMZ1BQ1LVpTrfQaI8KAQHzebKlr2wegFmy74
+ab+Epf0dIMn1CPlbD75bxBME3fJ/Qwmptm1LIO2E+vQZS0E/COsmrRzEoadfvoU
r0mpr61GMmgYdUZbY93V9Gn31hrKAsd3Sd1cwQmitj30sqv2TaQjRnElkt9xrYMF
AUVtlJ4P1NmVpbPjDA0ErNZaNOLuVe0aGre6scmKlxEnJE/u/SS3M2iWw2pVUjMF
tnM+8TZZsdDm9b4kczD9nIjM/3o06JB8hGCaeM0h8qxhgJJM5NrWtH6rw+xHFTJR
c0lf/X3W3vFerSiNqDUM95rgGFcxz2dfwRUGpqxR8HaKXt4rOyup9y+YiYPpRZjR
eIEq4A74Oo/6dKZ8dPOwlsGUDsQjgr/baTGKXwTVsOiAfWFkXmzoCMxJZbzgqs0U
gPHMMm02C++D9GpYzp95tWXy80vaiZHhct38q3g7L9crpvNcVAO/FdXh5vaS8i9R
eR7KZp+isz29ztGFDqWncWk+rfB90d1CjnwRWsJznrw3vzKlSGOqCHNJ9UsUlf7C
MKLwWiR0nKatqDPB72X2dmgzwNzWO4nTh+0zqBC+1WTKchgqyQGZBN8x4XIMLBBy
f/0aTwWMfjnYo49FdlRIuLXh0u/MmMYglF1qRZnhEHCGNN1q8FUqnWpE3XgaXmuG
FOwc77DS8K9khlucZHXK27kcRiR18ztAIZ79W77TYzM4+oXdRil/tSK/AHzLm9d+
o339oCQmzQrKUqvNKHnBGm+iBFP+NVB+bOwlldhxsFCk5dVm2uAE3KeHsDD5wtju
KblbtfzV27P2Oahs+nzxo1XUb7YiUWGBD+uzX75iJKFpxmyYH9pDogK8bn3j9HWs
m3aZ4uvuCIgG4QrH0JlTnSPviJ4MHXENN214z2Pg+Bn+69jjVoQUVEmsDSrFg84L
j/LDesgeYwdfWl7te9DWerTMzaZxAQUL3QRt2djVt3TmTYiw0MGkOrL8nRVYblO1
VtB/sAVrphikXxbW027MVSLT7DRX0/fs5I09VNItcTwZdStEznp6FG8usKQnUtA4
qGIHn9pQmtaSt2ywGBoC+frdjDhpKlmTAQH3gEzoji2na3nRyU+j8+eJRhsHUckI
XjirR86UR7T+8bdzwSNAyINcXVqzwIKJVfvkXX5uUoRZZHRsRvh8BG/0QJWTQVHR
noN/7nQI+CRHc9udpXJdlAz9SSMQNXpQmlD4yg3ySs2NO4VgU6Q+n6bO1TrwsVpC
MzkzNCW/M9CGb45sqP3EJZgD5UUos9gV1mvmMuVMEXBPHIoqRKmZTiOQYTImkLWI
tOt3rSDbcJDo3dF/VH+QK5QXhZa4nmXw3jjYDx1SFVwvIjn+K7rHEZqeQvN7Eqki
q9Ffy7f8O8KzKeNxiIutJKkZ14YYoflygvFPFjfx+iljMgeYwsXgSK+6qkRzdX7S
UKEbC7k8ht2JDoKrstXfw58wJpFFvJIpt8etKiZ4neiCSWqEl25OB6RBr2gXYLPH
J2bxzTvaU/OvfpgK2lwYLhu7NZ+fD9sQqA4xUss6aSJQJriBqkgQZh0N7QuA9l+N
ih37QXLFLFlUtgfsVjnasoPuUSPoy/Egm+VzlFBfjjPAiYJYX2ytlrmq91z7iL/N
BQ+DP3yhyZRA3pp1Zq1EdFKMEv/5NMT/dovxQINYY3JQ0JdTSedJDGrFu9Cx9IBD
dpGtQ/WdQ5xiX7zzbj4Nz7aCeRbO405ql6zx5zVUq+avvGLHyHASzGO0JHwcJEYT
E//tDD8u4oV7nFM4GMtgZ1USSA9TIbK3O7cjlN++xEnVFoWa5JYf4FFt19jQUsqM
yexHxYU5yJYpMkkPM/1V9CyQOBHZUud7R5kJp/UA1773wxqejgJhwVAQj6Edt3TQ
7kAoMMYgFs36iIGfYyJSksz0MtYt8sDLbC3vKwYhv12T/cGvyaOewLX3XrZGVs2Z
0EUCnxSurwgehxaTALcbBrnMA6/Ty/EqOEzfbMLP6BJWBVxco9Ug6kChaUotwyS4
vyxfZX5HF0Udi3C/LMFbPv/3OuGr25YFUjosjblPtc2ETpmlI76EtP6Bn/M9MzPT
5PjxpkK1mYTLs3qGM/aePWRstrZLvmt+HApUBvvoUlEmE8uEsbzGhzEjqSY9v/IV
MDF3/PbtajCOCtrRWg6DYVrL9qLsYlOwSoioI1+IHwhrpT7U2fPcmUtkukf9oBQr
I/rlj9lnYgM5HpPTBp163LG8L1lgPuDqs7FYaYrWIiZZkia8PjPRhdbZZNuBwMSP
pHMHINX4C01oYNFXLORXZ4gvhabMhgbAqgDTNM0k/iipa3IIRv59w5QskSlZQ/o1
BzSOwfsUof+31JBXmKcMaH6twbs7z+1HfBYMd8TydWl7OPQSigRVYa7gVvVkACEn
EyRnBF814g/NsZ2vv+K2FraTqxKzTZm+HJFugl23te0rv6HCxSxwzJ7xYlxTE0ow
kS8WU5jgi4voqLKI2P7JXsNirH63LtebZ1C+lu1pIkt3PD3COyyfjzne+hRIkq6U
wB/jRPHjqVgAvlYtArSBJx1IHpOskgA8RhnaljMgybDAVvTfLmn++0T0tgApzLU0
qYXumYlfPeruEcEWoF+2CXmRx15oDIdeEUWob7K/yEv1EP0SW8jbfErZtKOT0+H8
9IhQKU1Mj5E8fCAqoYnCqRMQkj85/hmP1igV+t448SUbz7qqkDWjnq7311LHnFzl
/ShlXlur7kx4NsSK+/ucspbJH6M207ViaNOI6PgkEOrozwG75FI0bSVrl1q0qGo3
n1UMnigS5NhrnVcLuHKX19L9i4OUf4A1HgbCTduZbupjN2G8NHfLGTyloJnkOUHa
Ltk6iIYSaoFhKcQlgAvsnJ7Ok15O/NyteWp59W6dSpXwzYZuAF+00Sge5EX3+uU8
kuDx3C4LJwt9FVkyu5k+RZBvDJjlEZGbTBe8kDDuzqqv49yc+hA8vWndpft00yEg
MiRKEoWGZjfHtMEhRRckO6T92kdJTC0klHMsDRQS6O6rHTcKvmwT3PS0gdk/p0S3
Dhk1CrIPmo3gxEwW6xdttQFGfWLyAn8Nogos7EIkYt0uG8T7ODmrxpUZAdvHWatK
5Ilbpa/HSbTmoWoTIzN9vjKZjwOTyaLFf6qvUezVM36jO3G2a9g7aJEihemLKM6o
KNeQWhPxlxuQ+v09VOzsDpWhYseCp7ZYVXOf1ceMJWP9YJYEqm1kN29ml7qJsi85
xRCmsy2B0nJPmTxWVwg8Q4VNo+y9Ezo7bmCYRHjntcLUV4qwCbomsfm17TGmtx1h
QtjF0mhvTfMP5ZsadBpMvdEyhAKMjbHV0QodjmKSF577bw3W5uS0Hz96rt0jNfJz
3eZmtbhjR3fzQTvyL/s7tvK+bjtTORimqz2l6f5NintUMC+JNTKNOSXspHonYR4v
sdd4VwcG5RusvsggcaQVe7irEleHI8rcl4yxAbwx8Q/+he7u2Bz0JHIDcB7wQi/R
6m1jqKvNRhjy4yYIL/IoRSKfA8SMmxQ0YLUx2UjuhNrU14xfsLBP+Yu+5Ks2ABz2
n/Wu39h5w/WE1d6U+mm8gWUVkh7aTEPZbcIjyqPhOeXVdcH018p2ACauvqC5B1vG
XhIpokO2AzlvaIYe8hx1dPQLC2Xacd2vkzVOLrJI+dG8sZSCg1FV8U4RqU3UoIAr
azqwwhfNQaEQjye78ghosbWd4fJO17vqy5q5iykZVf4tXQIVBLWkjsJC6lFr9nyC
+AJ8UWU2SNUBLsa3Af7y3QokcZIH0oewmN6fBmA1KQfmhbaQYgaakUSMNlFmOlSR
JLev11dx+lN4d2ya/fjNMwV0EXPHmPBVw0JEya85NWTtHqh2fBBEtziIDbfjCEtd
ssyotvT8qxdJ5rrPmsBzo3+snnRcTuMdTzFsThW0B26c+RernRIf4D4lfJ43ee/Z
lGX0DCVrMAqFsbPhzj8lM0jryYX3KC4iDOl2CiGxkMbU32NfazV82cnNHhKQgwMG
NGGpL0xq02/jrEuBhowhEe2FT6gh2QjHPiaOedis6ZtU0LOiQaVm9tLfSrd8Twia
rTFEGbKQWWEsATfMy3R2IM2A1mQYlAM7ggiukKuZaIVkUcx/uAGB7PhmPyv1p9mI
v08QbJNlqnJ2gXrTIC/R5dyXZOHK569G960AAoO+e7eSimlnPSUXh/dE9XQzIYZq
XegEbDAJobRxVBn28ptIwaPuahfNc7rwiaC03e3+KaiD1ix/fzVaQEk97QYN8n2X
NH3uI81TAMZCzGCeH5aostDL2fCY1UwcjQVpGhPJiZtqh8/uDCNKkLEH43+USjIL
wMYYE4yK8kf0IeoJmbw/6BiFKOvjE5a/XuA01KiEY/LDiJqc1NpRTTsEUqrUORIS
dBjRTwHlIjJVDmUVqu4jPpt93nl+JtJzGiNWYdkYXgs0M6b8wAqc1fzrfnFYFfwy
YICU9DBkoFTtjIMcoa69FST2lt3/vVx+NVtp7t4HIscWmi4sEQWxN3XgsIWUDcRB
8edoO5H+h4Ogk3AIUrfh7qX1Y+NR9xayCfuEB+gzVOHfh9jNIcYYgTnaI+pRQElH
rsWMXNM2xV1yN7pWSsCOyiH9T8TXNkKbtFuJiCh3II9SUFw7+pUP4H78f0pcaBM+
LnlCO96RJ5+I8CDqKc6/UErJRDf+wiun93k0nZ8/q4MdCaMOuAVqS7bUlSuPayBl
b3BOIrdCGHG4DG2zQ74pINESwSnlduYBFgUaLpL1ym1q3iTU3i9Z5zECkmRjwdU8
y+4iQuK6We9ldNQJtQ2tGU5oDthtTbk3cGFZsP6y/FHzDmqT3zuIN/xFhkq0FrZM
McmSIM6I+/UOgfXKqrlmbCSpntyynuumoroZmy8dqTR2f+HbiX2AmevrEteMVZgz
7POKcLFfhPYDfBTHnjNsz5l0WVFF+ZvJgbZTo9YKjCg2YIBuOUVhKHk6UPKtCgZT
axPloZoipXWn9guJUTTcIZuHHvPqWUSx3zQ3VkdVXk7XI7u53XcaFmvlO7ttpoH4
h2NsjKwUYr07kI6nqY5wptre2uUWljBiJWwksyPhv45ZEkLe06DiOT+xQdQ8Hb5S
D43hw+tK5Z/qIinnydAAxU0TDaaNY9SaLhAq7x0SEXifnWCY/jG/WiBjleXlOf3n
MMXRnBRtiPFKI/ePDRJs0TPipmYVRteyl4xW+rOOqm54lhku+Aa721P8ob6xBSGL
EprTldh57aTXQPXPwKboeNswa3HODgVu5JNkFywiNRunywU9a+K6AbvKOu8Vmb4i
OU1ytqkrcnl9jxpwV/bEKVD7ZxERzTmc3d2m0RPwn7uzAq8SImCxW1rBSeEoIE6F
MFQdUGlY4IPAN3MVkKfQVZVs87tlp6wNrD9kjwkpfBmm/hxzDBX2CfuO3DW9Bbtm
bhOSDfOTXCzVVEEy456gRxpSn0Bv+KSYDYko7T0JYWkeLYe1FQeg6+fsfVKg0SQX
yXvz3tjTfCkNn4uwdfzOaofV8+wVu5wcQPyIpG5gO/UpJG2oyXQ8MMl3vNqaOu/3
2CDlUUHs4GytBg5lnIv/wJ+U4syDcmYeMC1xbjoUBlERA/Wgw5yRbrBbqHtq6mpW
y6bThgIyCPbOxDHIVAP5FDJMMBXZ2B1KRXNpSaZqLDtT2tbDNY2Rc1QZyrc/3iQz
kSahlGHcxbjuryjyrSi9KoWpURT/qi0EJ3GkWysbLCj8Z5Cw7x7R9T/+IB1zgMv1
InESinslcGYxLvkyPGu5+ioLOlsYMSwzqaxwRBO4s0R4osU4WgOKP7VbE766Sbdd
EN+iCYe4wqXVeLAgHxBbRceMzbNSP+0gYDqsL8fbVk5qaefbcpWdF/OXTapSbpMp
FOMI/Fd8qpKMyAthb5zRE+uI8Ljrr51DmdtfvwpiGHptF3OGQHJeCOYNN2N/zo7n
XjBAN84JiI4WIbv8hRNmx460ULUbjqNlqpVVgllXkDnILuu9byPslnNssriycbOO
lt2J9Ps3S3DlV5niaFXMECyp2VRwEi8H0TZVTjoP1yNfHCcSwZA9eBU/kkzLFXri
uAVZp3e2t8osk9fLiXVNKdf0KPihoC821eJqsAMcfJCMIMKZtOGwEDAy9sDeW2vd
VZuKUfPziWy9eeRCZsziOkO2hpRRlUQO+XCJrTQD/jpqRvan6tD/1fZses8ioORY
QXLesAAHMJY2W8MJ8WW2tGg7Geg+D14eWN9KjPDetXipTYQ0Hn57XfxlLDs+642A
E/iao5ATIjXzw9mpB3F0bGWjYe8BeRJRopEmuwSpsWHgo60weAZ/mJHT1VugGXPt
+SWHUAo4ThO9inBZOrNqtPJKJn8PtBoxLfQE0OwZJNHUrHPJdz4BWdXu8dNz1jUq
+9hqsWdMrWp4LlmwvbqQN59hkyb4Buvh6x/FyrexLVyeLgTC9MnwhC1SpUinh9rr
DjO71TgGpRE+iL2a6krqeJOr8Mha8MHumHjoX4Aaw/JnIq1NwhNNL5k4B7faKwEH
ee0KkeXH7luwZ85E8HIeaQfkH+6DDnHp74jP2FU/sOwJb8eqLrALUqkNeU4wSYgg
DTA/DmCSdt4DWdJWXrsEnd3se2C8hBJ9yIA82Jewd2mFEHbJ0P2DnTGc5+c6fJt1
qo7RBfU20iKpAwB+acVvE2UabBKAFNCOE7C5UVWXu+g3knF8ow9KvZRlJdnfdesj
U159Nb9Wl/5GhwDUXnEC4iBTXgZSOGR7j66qh2hTv8ZDloCLtbPoJWPMYgSfNNDB
i0vbcOY2uCJKiMUVuVxVnHSWAa8zGRR46QmlxKgwtfcA832hpQUUKGkhldR8dFan
MSRBD54JXUy/qSEcKEZ9vELhU8aJsUK8HiquWDU3git39Qz2leUQjMYvWeMSYcJG
Iy1oU9feg6IkHEa2Oe2BNGpAVfR1wd5I0ExjjWu++46Fl7yPpD0JZJ3dLY/2YxDz
bbNCs6z+ihn0qBZBmLMcioiPx2l/nrIEeH1u9jwaCw5ZBOWpXJRg2UdarCxw5P5W
vpG6/QbniMjZfsoQmHkgbDoqnpaDfLq2ggk6EGyZmszpR/Za5tR6Ec5oW7YW/6ks
mkTAvXnKhSGdhpUXdVzKwV8vFIjJwQKWBN17M7iOTpT0y6cmn1wpAr98+tvn4yLn
h9IoPS5slsr8mtLBI4GzUE7waEQo1HxavKV2G3wTBH+CSfK49Zno2MNqnjjPDzKM
S/gBjU9D4QVxBWEDex50trgYF2zlBbNUpBfrq+zlV0cP/7xUXxdoYxvrvrSuO/+L
I4Vntcy7HagEk4clUBcRFHrt6AFztW+a1IrdQ806OmyZ0sYZLPAbcNXnsLc47S4D
6dxq2Ez9M1PtxDvfmb+WqByW/iG5dhT8VNyu46ta9ziHoM1bg+ZtFV51XswFw75L
RlX5K62u3/aRgaHMMq/ukyQCYmDg5q5tAHiy/ZLeM/daMx91oKNt+TMXQxv0rCsL
Sp6EK1z2S7tHq6shoMTbPNQsfupHmbDzL/izHiz4AzrDzuwXLKqBDdhmqi3c4lgl
qP6vvVLNwhifBqdTS/OcGZzOwMrNPlZWon2+nCP2Et6Nqnt+QSMUPBJI51lQ1XBT
PnKtNpv3iQkiatnzsVgXKXkUH5Mdf/yOZ/rVXOw2Ez22/oH1v2c5mALyeUHJP7cw
d0N/i0hvT93NjYIou+ueRUlyf7MLAFueRbInggtEb2XLYxtoL9ilWa433dCAlhUG
7IH64JucpWGcOi5T6H6aF9lrRvUF6BZuvds2Nka1Yd70ek/7SVAPvRWwjQ9UkePq
WFoqIrc3ebnZZZoek1M0SxvW0QyXIFCsr247lHOtrRBACrLUE/LqOoUC8ABOs/ns
KOrCIN5MKzRHI2qCInueCNOupNQ/9ueIZ9TRyzcvL78C77kZzDm4f9KLQmMU/pL1
c6GD5PDcJ0WGYJMi371KmbCsUlohdewBSdE/trfsVQn5PI2cucOyZP9RbL5aI2Sc
gqtZNKLDcgYplf9zaEm2dIOGQX/hloi/0/oVS1OmAc9dzBIYluQRSrTN5HfFtGD9
h9bcb+mP0JBZQFicF0W4bdjq6oFFyjyrb5r0qMvcwd5n4coXxUhIXo03D3ONjJkH
SMRYJWwrfDEJT3m5rSf5VhZ9jv9hGRIS2ouGlVgoxNFKhXzZcGRnNv+2zt2KeJr0
X83d8x3XOD5KseJ/YtKAG6ix28s/DOLHOvKQIXJyzsRV5h4JytQ2Eq1O6L3G3kH6
7HjVjT95DdZs2139zmrpvp2HzqL4qFmpDGb2/44OEM/gDYFIkB0XgctQ0u/ItKp+
HAaAgXrSyg5+w/9ZxOoFqkIGEI4s3x5G6MZptKiNYJKxOIxg+bO+sVahoy9TlkXf
vMxvlh6Ce5tUF2c0VaXonRgMMgUJMR6SiwtbFTMqByRL50Fj4fcp0oB7QgZQKHQG
/Zcztf3xPcLzo5sunlhda/Q1teJ9cNe+BqXy4LZuEfSLd8JxEeCiopzNM/IBwcvU
XBzFrtJyg7ssrEuVuBkSyrSVwT4uGD3rOY0bJeotk6LaR66Gwvs2at4dX6butxeH
5XO/txOS3g0We9tenyb3snvg6pEN0d5Iq367ofTdqwfldKlyf2lBvbSTD55PeuOQ
YYKPKx4yHKIgEaIRPn+kzjEeuAldcivya0fR6IgJL7FI3SCOz8c3bKmqsbcljzUm
/TwWAYMiyngrcaQFVZfWGyEmsPMANnCSWYvAsSqS1sPjU2J9kDwcllLP5EA21tOf
Ns/NqHtPckxP5/nXKar166Z1RiVYvT+etqke6gOXVpbHnr6HYuOGF+SFgYS3KFdJ
NMXNL5qN8rQjaVeQOkf18ZpoCRY3suxiz0G8cx2tqouTVtQCygxHXqJop9iPbo1f
1uN+LPbHI8e7YrvKPaKkstNBUu4cN5u41+ilyuDqRAIY2n8b7svDqm+gXuMUSuvz
vq5MGMwTZs/EktX1DuuDNLRdUE2NhYIOBL41wyIny+G1l+45CYIRvX9nB4SH/29Y
1+nFrAhYGAQ+Y4sPw/edRPcSmW0O2m9JgEHk957+F4M7NEEzLUOd5CYY/5NFjHU3
p7ThKGkc/nHcVjD2jhc3UKl9bNtghUe70RyUWdTajYGzK44Zhe7u+gq7b8LhqL7Q
3MTVCUiLorcaE2v8/NZ6t/zZSCCKynDDk6n+iehCq5E4HI/E/7tlecq3cge609Wj
3j2ysZmLHxH0hxwV7lEl8qxg/XAOayx7VIKJ+TwMhXJB9SopkkDalBI8bJxup1FY
3aXMn/FG0SHMRCbuCUsueLcUr4QqaO2Z/hPmGKIeq/h+5YzpTX5Sy9hJlWIk1iwj
CUoodj7D6son3cCNIHF+y5edBC0H4sa7xR2MTb7hiqo5yYpbJ6R5KuKocQRsyyYg
ARp3n+IJUmDVbBGeOoYPxHhg2sMjnUqr0s0R1RHAkXAtLIW2A+glikUyJAF0MGaO
f5OPkCKZnKgBXKudSNv97n6tf2nSJ6Y2cZbH7nhitn7ZfKBF7K9RaTSTIrYwXdwv
SRD2ogQRXFyTgF4kSZBWCQKrfgX+DzAq2aPOjCRtHOus+iNs3XbGEipV4A45EHwb
NL+SSr+sL1oTmqRVZps1C6/iRPBF2Wplp00HGXje7CtwkMHe6zC6SkLtGlJvGHuT
fdok+lfmj9Qbeb4swoOw2TtZOg2SMnM0dRu+vGK4MBylLz7oxbtQTvozLQ0ie010
+KMYk8QibArpuV7VSmdjj1hjBAohc9CRBQUSHRvY/vM7y6n0KYeWb646QPCvnjTd
fR9g3z3ddpdJoAEHt+kvNel4qx4Zmn5evj1gpHpsrPOdwPPXIuJadEQRCGnGIJYV
ssnxh2Ocl3ECD4qboMtIRJJZ7BsagKdHaIdq7fBSN567yo/Lbf9Hg03rEq/r6rp8
V+syle+NqLSb+Bwpe/uPgm5qW3S6PxbA2xuzLu3wLwb6qFxJcriD/FPvsk4ZoVLI
2kso2gWu8HBgL3xlb6Q47Uu9gg0Q8E7hTRjkghXj3UiayoXe1bQDiOKWyH3Wsfo8
eg/1+1rrduaL/Ctj0ysstq9OylBptD5CQXQ4T2mZ3uUjEdTWASCBciiclQgV1xjO
MjClfUvXiDnyQUf7OoWvZE1qLEt3xMMYGtqjQa6c4/10WtLrp8+ipv8yGJj6vH1f
yowCjVJv5miQAk4/4VUiCRdnRRRYNsaelPb8MCUN7/Zr1StR2hCMXuiFxLM5gmeb
Rn7D1d1qChFFeL58aPDqa+PK60ufi6eydLAB5YQXyqaLiFEA7T1AkRIpdfG2LAMJ
fREhchg6ZdC45qF2xEGjtJo6SEsJ+3/JKIWSyfguCmo/vkO1fFzH+LcOtiK3uCU7
PPEPLqLt1KEsmVqn++biLKu9FjHvYPIAJfJy//Mb5JWY7TYIYbIExDvIIm83EBw1
6W6cqrCDNVE/KHc9Kt1khjfHIU3Hh6VSU5IeZ7sQqXfIuVLoJI1NCviDBKXnxlxJ
sW31F1ZvbuieFXE2uUmeJ8GpGefSRcOmKl22EpmGTS8J61OVgu5NX4CNnAevgAhP
zi4Fz37fnsh7geZe9iBGzOSWN518xbLVrrqF6//N1lluh59cQEyaCZ+b30Wcs4Ea
Qps9XYE4uC72/Ojs24jBgtlfquHe8tXzVCu2D6ujDOPq6+i80svDvn2LkSMbcJq5
cyabiGA3uhrW9XksvmhR2dOcCCpC3pgDIh2wGbEZqfM5cP/byZVCfls1nvl2YuJy
xndEOXV6J80vaujsRtyCqLj4vSoSajGk3EYGvzGy/qsofGWocPA3LuNYMWfgCRTO
y9IWilDnHMXSOwqAztZE6E0ZovfZeJWX6QsayH1tw+Y6b+kOxYQUZpGWisr3X5Rr
ZSvpV9zTwrT5eGGfSpDslWcRWvU5TL0rgSRgHfpgXLMFgGUKfD+YoHa/leTKVkmQ
593UvOIuqpiFLd2jjtSlYN5KJN1ux0RwuEyoBvqTH+12eJysDY5KN81Otg/GhwfD
ZTnF1+DFKnnMhcZN9NHFSlonxQb45+OFsC28L1p8A0N3beSj8R9jfsUs3qDDkxFR
LRltanBWPDBBm+0v905eRV2JoWYVD52r8mSCd9LhN8YDUmTdqcOO6KmC1koxeFuc
Sj3Yq+5TFEvCMO0CfcajMQ1dLrv10LgtoODF/Dtwdk0xS7ILPKdYlxpn7aucNLBQ
0amdW/fA6p+ceDIEOzxB1tUK79qtwUPHNSkeZt338+p+I3ZYCmwoWRWyTaWGRA7m
rEw4UyHSriN4mcfzxP0Flr7U1KnbMS0ET4AYb8qMxOJeiX/WKJCYjVMqIVP+qysO
8qr3vkV6AWUSXbvOomMYBTg5UhWOXBFtUBncz44iebrm4impKnhZYixE1iPH+Zq+
8O4dksJhp6Cmd53KuOCQ0iXeXB+6+idkFX+JR6qLzTuqoMmqNdFGi1ePovFOkRv+
vsjZOWl4NI3PbRK+4L3e4dtbaS/Z2ZgaYKXBgUTvlkK9kqJSogo9HEVDpwN0F2nX
11nZhWafNuceRy8xAHLDbiyOJ8qw533wi41Nime0+xctaLgax13tsnCVb3cqMxHn
/+QYsHomOR/AJ3/uAjzi4FJIFkDXG6720bhicdl3VsTbUp+E9B+mT8Am5yqE7DAM
cewmQn0iIXdlGlKTlGb9OLchK3iceSFoup0m7O8BButy0YtYti785BSHLwyQIiWM
PjJupQ0fR+4EV9XCRh8eWmo/Mey3JnYYXnDyU4VGsji7zfPspWarpgUElQGNAypw
xD9Mn+2IkEszAZSTr4tmoqFk8EJSwgu8HgnHJmFlHACdw+uRPg2NG2EF08BiJztv
oYqaRspfjlxbceF0AjoA4Y8UevgQiFf3sbB1oGQ1uOgP9H1QIOIWYuRkoqiSs49z
wR1HmJASNf0cpBAuOtPH8BFHyUU4FL18tUN6Ysk9Hfyeikcqdqmy3Hm9SvNx1qcO
7AqghA1gO86tG5BxUn48M3Dhm6SIzLj5IYtoy2pgEO+dXrKjSMdJ+NhkzW/5q+ML
CtiEbUxxhTKjybAFAIxekaOKfwfVS/b0K9CWBXH1DA3cP1Wcp0cmwL0xcell/GO/
RHGq2c+Kv8GxG+RuC7Myetj1onwuTeA3swdO10mWGowmTgYFVbBeM6CDaU2kVjZ4
JJl9CuAvRtfKD5wz5VPRrM0dxKRyxd0863sh5TFyPavisuKcXW+pEo/2PufmNgNq
y1X5pi2TPogSTqJz3SR9gbEmWX/addzP39MzTGoSz5hR7kFlxrm63okd1F7x7FkH
jSPq7w6lAGP2Olnlexsg3wPHISvYgx/GEj9lWIQaSySxzM3ffEbnCOQ/U4HPakWl
SdzJIHR8YmHgOpEBPeWB+o0lZ42OoNGb3/Z+M1CXYmFophAce/mtxlTPoiSBVxim
WAMwAOKN/JTGfkQF3d/WYAyy133LfPQYIMxmvlukZ63OcqatlDQ9/OHKQho7j2PC
+l5rUCglCQgXl/7gbP8H1cexV6hZ7hbgacFbqZRJ9io3qzwHG1LQY+VKE/u7JxDz
ASnvKrWOalsGelGXVTvYWD37s3+SAnbOngPpsPqFcLpw1vs0PO4C/8DKKjOLp7SI
SGTp3/YQBzU68rJLxeXnOVOONXYBMzEeSgPlYM/hyQ//39wQbk/ZKbE8bhQW9q8W
o6qLOcvuEbbBYhMceiWSKw86Wgn24VvvaNcZXy+Io9Lu0gevRp8Xu3GCCkALApPx
LYmofMw9ZLvzllgAf+4/tc/TG/Y8zYQu+tZEe+X1gpAchChSlwpAteskAR0C9i/5
MPuk7dwjYwWYp+y+dfSWAlszu6r+jY+xDKyLGMvPwfJalERtaIdoi3T0xNJZ13AG
4AG+BwrxbKTzWwJRyIHEKffQaSPSFcezGjnu7lTV87mjldDGzc8JbNPPESfmPAE5
bc9BjrvwqnTl4dKP3OVh8TiNbRjOVGOzxI3B0cuKkSCdnAvUTzFgcMBem+xz7Pl3
PmtDZXXzF533Hwiy58FxzBTmmEYIfV5LaasIBrPfAPoD5VNQ535Cmm5hIFvOI0Eb
OQ4iVcns43KXJmDhD8tJZjJl6k4oyxEhw4Z2SfLF1I3PkqlTV9nIwkRG1HTIxsEN
pMhoH6jZW0ewJI/N2JAGf+z/rM6H4C+FFJSu/FzQ/AD8e9cvKciWIvmRLogapuSS
HPc8Zu3eIq5OVEfAqDskNRseHd5ewMPhnz00hQigszVFqynFajU+iSNp9yzi/Y4n
XB5EuWR0V3DjurFW+saCajHHtm4AAxRJBkOf8LK+YmwBRPeYQ4jwm76vycWdibvC
PDXsE3DzlcImQtTyx9nm//RqC0+SgLbSi6h1D/jYwX2knwE69G+VpQEVNQFVofqS
dHmTAchGFE1aNPAPi1JW0d1jqDpOT9pqRijLG4kTSeVQDpOFpheyVUU5QqwdG78M
X/rZk51AQgjraBzHZBCtlubWnCTDtux8BJ/ZArzqC+5Ui2nLfO4RSsuaINYzkYQA
Mbw4JZWKhfATEh49kYEMFYfvaCs2IfMMNzBR9LV8kwCd3v+tV7GGc1xE5hNTDYoo
vwKQaFji4vu1Hx3L1SiPp4cHiiR291NWHZOGSBQlVczWHL0DgY1udjGzlbHrl48d
Lx3UiMU1hJT8+gGkesfkXs5wzAD1ggIyVoqiKy9KcGivmAUoRDaZh6XdWV0LBGsP
KWeBcTzgBdYQ6WZgPl8KufkhUff3eJFjyaL9araDaVcM9jMYUFoPeKtPuNp71kSy
SFrJ5IIHB94Es8N2bSdYsgYTaqMED4IFwgR0oO/oFtq7a4rKi6AxxmI6k6U5mi/R
s42J55fhb9fBd6WMJHoRmSjVJfp2aYIJLIynPI0TA3Yi+s6dS/lpybLS01YN7dZx
wyq8Whc2uSPjvO2NM98VBQmHdIoF8UKM6A33GwJVxtzv4xrpwci7yuc2LCAFvvE8
mjjW5r+oB7FAzeIGsj9+DI0YgsmIFh1D6c17kiHHLs3a8ATLetFlHt03lD8AXAyr
Db4ADyrfg3zA42ao3sYwu0CKMxsKT+fBqNytyVTU8gcQJPjZmXlKuy9l9YA1jP2p
SOFafivErDTimxUwvh3mcS0bnNOE53ruL7gP2TP5dl6EGGlZ3dM+YisgC7nA3MlW
10pf2lkfBsLyENwiGwMYRVrSods5Td7l7avxwgOFmA2T10gBm/U//79uAgDwzV7J
Uw+ZUyDxZmjiSQIHlAhrBgGrwxJV1tMK6kaFLF5AOjmr8aLYkfHfmIcuqbWDubL0
lKQwIjHvPzGD+uFXvtNeibe7ywf+9PvKh5GM8wTZjCOgI0NDzkvChAzjTYyfqeFH
54ualV/qJoa6/Uqvr+TEXpnajVymgW7qPQwjqt2Ns6GfLRB+wxQNOxipiBI1TOBj
wZ63MSpzOnM8nI3LrvXkQ6ym3NLwieMDQHOceBkzJnav7BGodI9e5N0pjHUz4vzr
16OCp7HewIo2fSumXBIHPgzCPB/T6lr5AblJFlSQZNNJccUvMUqkuW+f7JmHqgbG
VfkTM7xTbf412xjYnet6Vwrk+fhh1P2m8O/Bdw+s3T6/vuyVu11+hwM6cK8WiBlW
ZFgSMepbmiLyil2lDU4Li2DDeX1ISVGNpkU7o7UVaoemij1Gf9QC5FACfRWcO+SY
jw4koZOIZoY76zP0sSVJtZnnwzwP0dc4oK9dRme/oOv9Tk+C5LngCTVrzd3g6XPo
SVKUY3rNrmjXaEYy3Yv/ks7pZPgdg2oTxgf5YeLD+QrYmhXt4L37pZOEixs7ZNzx
eXzp+RUIqvhXaooO+SDKH7su4U1hjIkF5Ew4XchwYw97D+kHMa6U9M85k5n4TvlK
tFd4vRO8dZT6TqphM06v9as1aOQVADMdHMoVfKfd8sP7h8Kb5xu0p6oviJTbgjGd
SK1OQJAV5mr2n46sDUAwk3IVSihi+DRlblpxSBmSZIMVA4gZjp5Q1qHzFtQYtV/A
dk1Mh90am53115oZpNEbahemg2ZcM+p9Qe67FSvMiIDGw771Wyf+TcsNxwmqsBgJ
jNO9uvSJjSi3W3V1n+lkMKkcJZ7qUZVz4EfobygR95+Ff6SYuXa3FTXBaqgKg2Ry
Q7qzMtH/s/zOgKacxoqSgFisRgRPoWeT92ihu5WcubuaqB1MEnCUwLzTSJylUfak
5CZvE02VuJl1A9Wwi+9gWzWZ0i8eNLfPRbjGfxvx36ha2HWeHD0yR146fWLwS8hm
xXooEaUgkGjxxpnyIt8gVQLFB3u9qKvOdm8Oxm4DBrTH3ZWAbpBqCjSr/ONf5OD1
pg0mEtmee/ZaRFEiZHArYqIGbZIHN5oV50FALDj7jkNKf+oH/PXl19pJgzndfoSz
FT84AgjJC0Lnus3eyrksBCoZFBMo7g7Cui3/1LAhJvWfZSEGZa5/IPgH66eW5qsn
597e7Lw9Q2LPDN1/Dzn4+dtGh2IWjuoUo7E/s1pxurvNm/9HTCmMesMuWpPMAyhe
CviXDLmwhz+viyDB9J5yyT3W1PL9D3hisXX+A0Js8R1Q3ia7wNz8dI8JLx93PAfF
cg5rlZhDoUzl4FMGIUn4mGvz5cAEeBM6nsJY2YRFZ7YV20kZvUhGTBuwm7FVY+Gz
jZpP5ho2GrCYDmr9bn7cWA5rOG8cDfmmFGEKcktnaHYEieI5dTvYXJwUCAU4169e
ECLED+6PPtL1VZTwfJY9rvno1NqeXFFprZ1ZfqxhT2cXH/tMEcBHfX4rMg127tGi
+hKL6KYGLBf/Xww7qaBiXoXRjRYGx856S1uNHqT3oFeFUxpBHEwg4LG+sjkWv3rK
016szmFq9MuMac+xl/lB/y/tFE8/oRir8AgV0zXF2OZrWC81eLvA2UMBevce1jQ0
9UlsuAb9v0IQoKOQxR4gpc+5lEalTZcOk2liuVebwGzP2T6rJLCegtJEaF3vABI0
SnL/NiDl4ink+8l1QBPUT8Xb6/wjXtm+KCni8PEKR47MXP2X6E1nIhART8SWnslf
5KNLZ+W6xuKlv/fhgoLKu7djA9d/cxKImZ6jKONF3p/pX+qHRZ4TgKU+yhLD5oEi
ow8R+Pr32xBqUCaXAuCuHQs6by8f5JHKkxBV+xYpJGrLyIIapOjDABKqSbzHjxrR
ts6Zd2ZB9uZ6AAOHd8QQIOUAznZ+94sSda6C4/QUF/pxjPKMUvDFwPAdn0LjVtNH
WeL7GqHDrFWnZUQKR2St4dRMoUT9s3rmrLneJ4TqCbPRbbLW7M3OjZRFy9tSQLI0
JLr+wgb5I8e2He7aTU2uT9P7por4moX6bHVeJX6jtoIEQanWWcOtoNLqA6px0TnC
Gd37exnuqWvuz/Xk1EPxnoZVUdddYWk1NbQzWHJjse5ggvbdfE4KfHbTrVHD4AT8
rGOuL9nAy+sYE/DNW28cWm8HO7eonT5JUD8cRmYEGVdXB/tfugwAWBFsJmkJTPPS
BWcR9T9EdxsEqzrBP98zorGfd89wz98PWuyTxAzajO6YV3n6wykbUWdcbChmDgNj
4iPZNxZC3iKmvnZZ/iULFyQkTShnZcRYjLtGyg2YfEpB0vrt9/obCoSeO8rD6ZCC
DaS2TjZ+yg/K4qPH76/2PE7AJuIpRdnNtEnCeq24bDBIz94bBHGY4fYA3DjtE/uM
HWdpAY/XcbnM0kPFcvnmryY6xWlIbAUauBZDvWwdHM2FoOh29ke25Y+lc+GEWwWY
Ow8bj/jg2Z8s1sNePh8QEln/yhaV6uod8h3KbeJv6PkZyZv+tVc2K+kv1pfSEkL1
LnQaAU6imlgnG1KGzYqd1BD6rEGi3AZypOTMoCcN3eZyaWhh92CgTJXJCkAIAXoC
Ok6FR2ewUQwK82g6wuOrrysXrA1Ac8e5HBU/i/13br7L7w6Mc7d/efoDwV83+bSM
0eQtVhjPMe1Yb+GoAyJKE6cU077Em+L+vyyVj+rqLpB5LZfJGyIHmYc7OFBwKXiE
8wPQYnZToZtEYWEo7iM/Zm1PK1ehzTY8rqg6fDsqFbJ3XEv4XLNHG/x6aGStuX8q
+Hit49mGXpKf9ZFldxxhb8AH2iwMV3FgPsVKMGwUn/citFzfnIYsY7JtIebGio7Q
HAy0tuScLv3mbZmm9zGaNl2z1ces263451my62amVe3+jv1lDPRy169xNBs7277z
uZUGUgbw9hLvEke37a+G3NllmRNl1dGXQ7BfVHfDTSBlUoDEeDdAzhUu6Ch0GErL
YNBdS/H0u8shw3/z7X4cNG2+HH/oYKU1qt6f8Tqcl4jekWzAyALLPhyVtHh54us1
yzqUhTV2oT+/dHdG3Fx2WDVLVGVJsFoiRDaz0+m0mHgX/3OpsE7/AYjwjd+P/8XX
7LdiKyizAl7I33ZFRbGkzdm9JnwwhltjGu/JLztZI7hQfGQ4AMR7N5kLCATJYPcy
XIb9OWByJ2hquTXp3InZ2AWO5a1ElCnnV1pWDxNmH/BCpSwSv9jSOK/9PE/OpEp3
/voaG7Ta0G72LCok2gXWdJI9vwNtMykKHjT+yDutV8eX0SDpIR5PEDhNAVHyc8lv
lAKgaL7EWK3wfpJQ+qNSZu5Yluqar6LK3qJWUpfe2eoITQ1i97nX8E/hVZUrsSue
UimQToxARBcWZaNcynAGEBXM+lyVjnrHD3Gpw/oJXQpO29UyteU9UVDRcaUjY+1K
lgxaOScPaOEnjJk9882CbeNFZBCWUkXiwR59f1gj74p+CH0C++4eunapkmDFW3Vg
yoeSSA6cN3EDlHppXClA+aTpEYG8xMDsMqb/3cTIGiAhLesXMUK3SbzLCc8gNk68
6aTchZRIjiaRBq5fSFvEwqzEdnBjujvvpb11emLzcZCUv3kCxBct8RSmG1wReYXF
unq2EqO5dk+TPMrbLyHq3QdQkwFqRGcxWcuJuPqYymvzIF3tHKvSOURpgwF0Dttn
ByRn/QGdE2IaTh2KMj2LoBGG34XKcDN38j3b19G7dZKZqWuv/VQ/j5C0F+6LFy5F
ylcjYi0TBy9NRu5o89eDo2UO6NqKaDWWe7lqQgEoFjIstCQeQq4Hf/50PNhM/ika
zDmB/YzRhbf3xYoRnn7jxg0IoG83jvv3cLBLt6CE+/9eGFJzEAJLQwtU9Gr4k9SW
n0AmD2zGN6PQBzSor/H3sSMI7fYmlXpre2OLNZiUhnwYA4sblRvJQvkMG+59lxi8
AJSLtKHdKg6zFgIwFMMfnmykc0F+UOjwkzoJYFHduh/9tOkpUw96j9m9GIHR6TRr
Ob+ATbLgXhG6Uh/YzM9yPnZ7FF4iTy2b9e2VtEpvt5PhiSFNSu7d6u9JSgBV90Yx
3G71s6YgwmcdnwStH+I6vPWtStf421IyRVfKedwPa1E5YAvj81u2b31N0pgRANxK
o+HkIVtenEcXTTxf2sjuUcgzNGuGWUXvAYY3x8X79Y+uFgmGAnhjWWvOeTSj4bBX
DXPuRQQiNpWLm9DS6Cr00Cog/UOlrFXDEVPxlBfz5NEQCcUZTdqvQBJrVk4RJ90F
r+ZoE6VDLRb3muPn+G+JoXMti0YELYhqwDHUyXekJw8MAlLZDGd8SuuNyvYIt+oQ
eKS0J+Un7dZDJENa4kEpqYcs8sBNYnZp3XasDMKwiMLdCqvb81qpsUwG8Cfs2Z4m
1MGqBu3dtTxY8qdLwzwVCwHOwvGbjRtF52aRPsyiB2tuzxUZAhToojU3DOIv9Voo
jF6q6O53L29ZumfCG0zCBZk3QnjXZeikmPuD2kypwlV9adlbZk3I2iCR2Rx0SkgZ
PuyjnyitDUamNDtxXuBb15M6Pv5iglFff8hjjHh6ObiQrylMiimyKwMlRHhTImg2
F5iq9OBkDofeOS3k3h6gWRXsyOxkmyHewbNTCrE/ykXHh5uZ2/PIJoyvDr+Bix8z
kfx19AphEUSVDrzGjODbCJbUo543PtBs4869vk55b61rH9rEpwLVhCpgoK/wNQDO
2cw0JIO+fzCWLOG3nFFgyOIjogeDSEXlIRmxpamQEy+qyyzgTvyBmGi2aW16PmmK
3q0TK0OYYeEDQnT70m0U51c7Y6FYjQVAcX/1mryN9cWDouPh9Di12eE0mxrtPKbC
zX67bMzjBsHVLgA3xT2iBJrc5JunKoYqHZHST/UAhWON/EAbcySZaJoc0m6A6fYI
d4moqgfuCSzOsRYikRgfYaGwphq+gtYxeMJ2EVsYyLTV1AUEVWqbSSH/C8ya059h
APxRXY+gFOwgWwgzwggS9VNcWN8efl22DMd5jVUwFYM2DTyebLs1V2gMiOmHxKQO
rE0w8yFTw3Oh4iQt/z5ArWoLXnm7tlrownQZsEPeYYqpqCnzmhffK1RmRuOZmYOe
GgZtMyFLU3yT5VFKrRiRa20XqkyWaiSVb20dzBF8F4+oO1TR/8s1Uk4airBMYQNj
4rI1GCG5EBHAyOalb5hLwjg0Xx5gW0IsN+3FoHSgp7cSzxSy3nUGb1ecfamFYShw
kQqO+f/wXDXOXJ+lwwuovjiMlxqkxvsW0Zq0Iu70em0ZXW2BO3+MpkLwnGw9NdYf
LMosEnfUHducXyR+yE7oV8iQ5gFY91L3K4nN/xXW4av7gd/rwodt7sg18ksMWQhN
YrITAgYk0QOBWSo0djHun4GnbBZqOKCJ6OdFOJIuN4EJdgCNWUMqXpQG37Ua6P6U
HJrs8uyDxDVGHInGRLnO9mEDkRzz8x7bclL7ujdyzjYlm3QOPj1vw7LxQzbQl54G
EdBDb9EQCV34Qmsgvaya+tFVT/gZWwh3kuC3AEmQPV2SH4/DfNg47x9GZe7B3dDv
/Eb8guWySI4L+b9XxrehWqCAR43diI4BozZAL7DTOoJjpkX+c+TXcRgLhdAVihu0
OLznA7KSFl88f3nd2jlZyr8v20NE7xQ9NlLHRszw+aDsbQEWyMMGOz0tufSCmdJO
IjNsQY68V951EFoawyWveCt6QLmsitdUom/gCcUjKdRYqLyMfRV2amWyXO/f45o0
q0F8Y8PzpzCpfrKdwUAjAxU9SXJ8djra1bbOSIM1BJfrxcDwpXYQ+O5fMo0lqJeC
ezIRfkOzUcIXPOaqRYYw9P2xBeYFkTedR5wn/faMSOQ7qB/vAuFhhXRp5c3KInPj
/hGOgkcPi8P1PdBXQz8M7HB92rD9huQqbLBH+6gp6DHqRGTBwxOumDnUEgNDzxmv
I5EkZwu78gRglnGGnD1m/BnTtBKJ0xIOOcMnv34ChRoy2vmx6iBZQado5+WU3P+v
0xY/YAl6nyXKHdKvxmFXqgsI7UZJhd8UCNgj06ZBSU6+XlgEs2VXHDUKMSPOGkC+
eEOVqRjYliRP7sf2489x6fKex8FrGbWTvJkRNPauwUfRYqQbcJlL2aFeGnZlX+1a
SV7if6eWrdUyTtgEvjsUvtOTd1dzjNePA1lEHhOm+bwohkshqt8dHqGyAgZMfexx
hUakVk8Dj7A1mDK+xs9KBpQR5yBuyZlGdr5JbcoGXCoz0VEBJUFPM4nkPxT8mbeI
0g2V4AwE8ieq6mABF5kqknlf3qC1NQ/Yu0UgOEc1R8b7N7lDsyxqrOxaNRjzY3Ln
PbmYheCm4XriP965aD7jFiBt2IrCb6FBcEl6D60/+kABxM53ze/SbxQWzzsd/a3/
45HbKTg9JYyrG5oD5oMcXHQ/41O+o+3gNrpWkZbXTuayqBIv2L+PG7yxh4VcamKJ
AGbw3qiqIlkYYCvQ9NqfZL4Kx9h2YTJB11eUlaQZWRvHjRYtmJEnTsW/PMZdqWG6
M3rr4OFZ790MHlOC1WxvXuYJtxLunr5GmgD99y/h8XWcc3diYRXGspZi4wONEsdC
IdpB4atmgkVFPeOUB17Wfo0S36Vcf+c/jFDbu0UNiM0+agA7lcwOGAYhtj9OjGD0
SD9y4inULHA0mJr8LobbVuw1O5E6uB8zNnMVIilIpnGSt4/7OptZSd1QFy7IDNlZ
5X8g5dvqYLhOL1CrTTT5nr61u0jwJqe86dJ7grufCp8s5wE6lBLopwLaPqUplTpE
2T9VqPoDfeESm7oT3sWevINJOsTTo5vuTk/AnsjArznBrsW2Ywy45H4+FL68P6DU
gj1w6tQhW2gaKZehfQOYtk9ottDQKaBTRUaTr7H3FwREpPio7WvnN3HcGwL4EoOq
BS8NFWugFr82zd19sOeQz4Vz2jY9+N7iNsFZZLNczB++MvCblBY5WoSfQXKvuNx9
ulXAb1z5b3tYu5ICdH9O+BLLENM0uYKICRmEQ321NlSnvfRQixGxkQ1UTAcH88gz
d1y4/HAjqMcFcMNnvoagrcABblryaIbQ/1EcY5lcGawMIyXICOE+3VbXiwigD9YF
1OgT7VPr+Z5epXo2EpQSyAilSdAZklbV1Ev4bSZ4vEj2mEhfgEelepoEJgQyb+R1
H8l8W4Tr+OBuFi5iw/NmaFPboygVlysXtcY1pCsnQg7HsAIrrhT4MSi9OYcZxnnE
+l2mkolcSkZ4OnaveKD2VvJt00VOhSExM4RxrgFtcFYXEZF1uxi3O709CPbqIXZs
5BdugokRbmHpmh/YUMppnZbEzOFSkvwWCaw3C/5INmHtSJBr8L7Q3XgCAa8gw6gi
SbGTSFnIWbgQrVikO1PvhiOXvelrIwxsA0X7KxEib1Bovv5ReeYbg3G3u2y2yVFp
2vLHNOmSc1RsKsV2n2LafrvPtHaMv6pgQ+z6OztptJ8U0h9pIkT6ICChZ7iYSNT7
uw5sus3Ynhi1nAxJ3lo5UmzO+hQGtOjRUlZHT1IBkidD1IohPKvWGAJzmi2z4yiu
R8pgwNE58bHk9rGoE6gurGJa0XAE76OEdUUlvtvOL6MuVsX9BWILchTAQplhfgWA
lgM0jg7L2D8iqAbUsiaZLDe3xizKVMHO05kMwwXd3ZlrcDB/BxiKk5ZjOVft29zg
OY2W4VcCY/Ah2ETP9BbBZIt9sTk/e0Q8YKKd/KGocMQ9LDScipIHfiiAn9SzEQtA
vx6HE4Pa0VjyUDVkEcJ/JvzvjbZm/0SGEM8Yx3y6hUFWxuTcS7kx+4s9uPBPtNvB
9KGLqi6XHONFO59cRVvIMRD4fHPgFS+I67ffQ15PONzZ4sWwMQ/dsqhNU5Kb1iOq
H8mNgN6E1vK44aP9cdBs2nIYddZPnMVIJELapPIMAnctS7aTcICEiLcDKEKrWAUF
2N3FcCuF02wOZQXowbX7rT51yJOLgRM+UJ3McTJSz7EEwDUHv0O3mltMvYcdVFKs
WmCsCYiguxdCUTG9B1WpIbdCkIJ5PSxdukgrpdKBDLB6M8VXk6uGZZ1ckv0mksmk
oOOvlg1b1pFjkKSWu4vxe+ZCGHOhiYmw34lFvNd69rjwgr1lr9MkRjStrDl8XtY9
omx8J2OfIKHbVp5WD+JrfPaDCN0BKysoJxB1Pc5+CY/8v7B2ASmXtbAPQLqHkqkY
vb7G8TaJ0Qf0gWRq+5AfiU2vlH5UlNzQzrDY1Ti2yUdCuwNE0KtVV+e/saWp0TFA
xS7RPMZovzBMOReJp/9A+HbHGu8SsQKhbS7pPfgDD9fpK24tAYOPXGyjFzrSoFOw
LP2uAG8VQAlgKSgVhQ9NMWy0lOgg1toIb0kocBOYEz5Il6dIBFf+wMtksAUbot/2
Rdr/Vu0AY/O7v/ReSy7KpDenUsPlK3HIGRvU7eHSmLNQYrpWsbnwm/AMtMvyLGvh
IGYRwwAA+ylGtALCo00EpuhnNAhXw/1kmAY/a/omlzuCZzbPYAFdvz2SF6uwRrVo
oGUdBel+27weIYp40CdDSspUjw8rAN5wwWxiloXfNBaW0mA2q9cSDwarnDdnWu/u
SwEsTqX9noi2u2O1zFysRca//Tc+7HvkRxueQsOAWCjxmypnO71HvfkQqGo7rolY
CUpVYSGhQREOw8VSwbZhFHqX0oMSE6ypWe5QqXhJaHLfKHYymdnjBEbjH8qqeAYz
l3gjlJ2qVYK2vgjqieHrEZjmn6DDZ1ws1fLJhP8AXUpcnKfmxTam2Rmn6VrtCO2F
krREDyiAoc3GS0Q/DMWpAv2PDs6v7/ThEt9lmXBaY4j54mg35P9Ti2qkmKhyQSTq
XvDMc/atVuLmS5dBlibukpfMf/aWIx7hkxkL6tJf0j6ol5ySXa9w4TRYuxeHT4Qy
NIUgeLk0vt2vEPog4e0MdbCCkZ8lNxIR96tkgIQKkCGugREuQdqkRN4vTcKTinKX
QFYUfzP3ZDNYswbESLQ3BPVhdCbjOURXkF4xhJA/TkxV4lrJr2Bg1KcmVkndLY0A
CBlNKM66uQoKJT9M65HzTO5xZBPhCphHHMYIfuAyFZ/pBbCm7cfobYE++O4tulIU
VwdhpL36x0am90HTHwnZYQM1y/IAyYkPuV+MCoCLdlhJvkeBCzTUszfYvgChN8a9
3p5koODQbAvgjUkTGJq4xhI7R6QWBInMFKs4JoDKzKoXjBvYLLjI4Lmwx7jvhWrY
SVEEllfD3Kvl7t7nFxWevVTWXZOdKQ34HpxlTng3FPNozboyK1mrYpYSoVEllMeZ
/Rqh0B80eKWQVGh6oC8DQWfBWQ3eaDGvNUZcOjy5SKIdg7n4XBTDZWnaWIlqc8th
U17UCufqpbt+28QQzW8pCygKYqPlqIbksJPysPsSIHo9XFDcw3l/YDPMYg/TGwdC
rbBZLz24XSvQaLOTdp/YHLY8uHMiKgJXsymM5MdtiApo4kLuENk6IN2ciAsyvhXl
vLzuzuTCGA+m1kKQMp9yk/tPo/RrnZKVe/E5wjPLKZ/fnmgsDOm8djOT5aAseBOr
pRq8UGce4yjPw18UPfu5gk0vKn2USUFXwWsqZ7522e4tQvh4pCUYBIRGpIEYtEjq
oo8LSZRLygaI8k8c/5sqFWMo8AiXSmu2dsJGdUrRJwNjF1VnqUhGq805cMOPCToT
UGHhY9Yyp+jt7bUPHx6IqM35rcgkFcwuBz3WDH4gVeU1XsUbYMOMFvWrzVIrBIsK
0T6/3wxDxUgebKRkybi5pEhUk1cE/JyMI3O+McjW1f5VLStmfSwxiF6WdF5iPQK7
qHDqS+olofQiCQ0a2KZh6AjegzXDJm0sEs9BO9ovD42DCo7B5sy5nAclGh6N0byn
hWEYAeEWo9d5BnjEDv6g8IQRphZMxKmTxjXXk1tS1D3Msmlk/XCHoPKSGAo6HFEl
ZRxdDJy27lb1a8ZRJSQTWVLTLPmUN6e+5vYTtOlJN7O1C0iIYMyYZ1TW5E5yDRXn
iUyuTIHoBguwRzsYD4R5+xKS0yu8DQZ+9DMGZGVolfHLd/biEHC5pug8/gzD4VYE
9zoM4H58rkaY4MidTbkjP6SBqQkc/K3k2fF/67n+EClM5x5idoPaMd2+GRkxo960
5MCgq5Mgsu5kwsKecyMtFjR5OY574uluyeUevkOahdix6y3WiRJTeCSgEKa4QOB5
ACP4eQDNppH2wABoJJ9Ffqa64GUgwWLtgTXPcGHVzTGQNqgzAkfcZjF6Z3IkBiqz
LT5yvmqFeqwFjn0SnmwsEohrTp9TOYtYgUal6/DKpczivkpGjZg+z+qT57xJudEf
9it8yaRIKTWJ/rjGkFchr1jw0iKCD+9eOMZWOcqgXHROUFDfFqw56HddiQY/NT4r
v0mTpnpIAQ2hah5objvb1FhrLnoJUkBQ9bFrFQgXR4ONNc1okSe+beI3nw18OfeP
hPZQUIZ8AJhpEWYEnaFWcwMOSphZeqIYPA7b+kcewSrsa4ytXXt5YM+k7bPRvCEn
Ua5ph0gPlwyjMHRZexHodiIv7DhfpMfe0M8Lbi05P1zUmkUFvlzzRa8Ygn0qVrJq
Wim8UVMHPO/g0YViHTGAAYlpzldnvow/cOfFLUsFlDUR6GbkX9hRBZ6jFi+GlrGg
T0PPghx0jTXz8RNuE4zNTW33tu0l93Z2P8caLuav9IDFPmidUDI3jzismLduUilV
x71armmETdntzGfF9BdPqwbKZ+bLL7rAJHRQCj8xFITD0AS50UsUz2ZlBVqKIjmQ
ekBeOCCkQzLfSgEyjbHQXEclMIoCEvfM7T8Li+dF81lZXSaJqgxPzN6bfcF9hzVB
Sc5YnM3ChkEBzRYpvOXL/Cl0EQIW4YfL8H4QZJw5FFcw8SLniweIkKzKittabnOJ
Kngc0JoX1kgOjHbl3MDqYwuPx/XtoSAT9c4q3e5TgOWt/Iw0LmDiKik0WuIRpt6j
iCYT0ShVRf7rygJZhszR+0ddumwwkoTZCMhSS93LxFJQL9GbDwAw+XYhCjMRQloe
AfCJy7vtarkrXJ6sBz67y57rY4gFpIR80H/w2vgdzBPj9lpLHSXHQgZBxXZePoVk
KY6GQP3KIVAvog8JPtZYJtXNlgW/fzV/a3J0J2iU0SntuCYsYBshOazWodpF8hzM
L/3P/xwkIzKYVYDG7N/240iNS+ypp60R9j6pJaUF7iXER6r9rBK9JnmyUWdtg1h0
6yIC9CDpNSY/oIxSzgVakys+gK6xfb0gdWHkp//KrDt72Sl8kxldK1H0mMCLE44r
uejAyiELb17zSsSWtvdbkP0uHwmOI5o3i0oFWeJXJ3gXNHBbHXZvfQilI5di1icS
R7apatrC/erucc+tGlo7PrrJUoWmsmD5pLo7CzcudO5mySdny7AohwZyYw517wkE
lElO06Tm+fyedb8Kx6VElK5qUF1iyKv8LnWyQF+JIOZclNtXJnzS+CCUXERm6G/M
ikawdSOLAF+ss5EnElY2E8lWe44aYXa5IPbo7sjFZbbGFOIJZlLqKfVrgbT7ePfY
sNCTPCFInBCyMb8UyzrwbPtGxNzQYSPQNt2HIkyMsKJpNsUEcRMR2ksXbiBvYr+Z
KyTuCSP5GDATzDPrh1xNcDtfJtDYoZE2qzgJ0pP88UrXd1+HYdGGsYZLlYCaA1GI
kkmfrHKNCASCOEe4io30TzxatVidW3Bfmi23p3imwB9UUYfxtvldjeOUGZCYbF3w
LmcPDnpXRTfUZBuylAi/VSZqFBm1FbULIpekDH4//ru05O/cJPhx7YAFB5C0qoEf
KorKwx37sEt+BC0jialhnX8mdBpw5kpoZscXudm6dG1+iBlNhoVRl4+WSxXMowLq
vQNe5vVMiH7zzPfZQ1QWy4YYI7oZSXngvjzEXfG9Jj9yz0uG05INdobG+UXt2Myg
g6MOeZiXz5QEuVkCKEfWwkDOObd9Fa46yrOS2L3GBJ5d8sswmRoFFGjXc9K9LfUJ
EGTUqNCXjTsLGWiXqqRHtpC+lrkcCl67088aYl8TzEg4hw06s5l+yeq4ExHXRJoE
IrDE+raqlhiOcaK7ls6VMSsnUQCyrxxNfpHJmLofxKYVgc6npK25iJHju++K+kTG
QeM/76b3zbd30R+26jpKjX7Q496S2Tk1Ix+huaetWVx+X/btImVlXeBPx4snug5+
jrRDI+PWJoZF6ByobY27WL6GKTblZOZaT40paip5JrqLYdP29pJiLrAy6QMD260R
Io9ydyRm5hI3jRAY0j2eF1tFck0ptEcxEO2aXZkBrJ/4ysNPJ0Dhd1PpE6u981oF
NmKnusgq9uIu+DhHoO47B1wgoH1ACHN7BO2j9grqBitlXiuF2YzhPiFdcw4jtJb+
8H07rBNgi9Z2er4e0VNSHpbf4PAaj19eX/UyAzR+prLnUdiquq03WrpS3BqGHATv
bfN3T+B1Tnw2lbx1xqEif+zRqMm/8FmM6AU5NKboOok6MUv/FH7EfZswr8JZlsgd
qyMYjF4JbCqgRiqzmvap6aBaCLg7s8/FghP/CPUexERqp123Ks7ylolotX8Og+6f
8vp1XBOW8C8CkRByUxZHcSXb15tsfeIfS/Hpya6FS9KcjhMBajT8yk7ey7Gtfew8
cMadBXcJHOTaQVLESapOc1LNEMCryEm4tmhZvUN9SMXuHAdw44kQ+t04XkGUGK7D
UJkeA7CVk/WA+KroPsZhR1NSJ3ffnKjT+H50ujvSOL+n5NXUA+79GaiT5V0RNCck
H6Sh9Ynsbdr4x22rZ8BUAy52XR2zYgzlxos8/bJtVXs2pnef+Af2sw1APBx8EiDO
Oa0Qy6iGiELaBcr/fsVenbAoNSji8ha08lVDp3Xqxrw4eWV+5GFrzXmNZ+tF9MKq
lA8r8uVUf96IgZzq9UYOfmuNqXFX28XCh/JU2lnnRzDgxUVV9iCHsiSTGUas5K3F
QosLNHTffjSGyOz2lg/sIfkrhiRe/vxc87jmzyTgVHitDBfRaJ2Y559mklejJwQv
7xVUGEWani2Q7YuC8ydruwNennDspsAjTYb0DrkAUXe65NXllf0lCD10FUSw9oio
Uydoaq11RZ2FdHW7JtWVEOVlM7eBM/vV/NsJE7GW0ktgHF5XmmgWxIlZlRpUobSn
FjRRWs72LlGEz8/cvVVKB6qtt6YURd+MeoeyAq/bLFSddIaQ7TTHCaiP4WfPzwyw
xrNUAur4PGL/sbeed+fH/cqGGbnRY9k5aboGjHr6qkVJ1pqIP14Ka3dYIPZMoA+S
kPoDY+/VtAMpj2ms7raiTAQObMMRRLx0cqR8cGMCnxwlhvoTBp1GYuoDq5XBm5Kv
v51gkA+3Qo6NIhtv8fCt9z8qkMk2En5NCyt4sXAxYFuqXt5jQkz2S9DmWaPICJnR
SZP5Mf9XTTFG70PqKGcl85a0y3JGeitBDMgGiGbhdViAIi1bumNTO/PHu6nMelT6
PghEvch46dX/vwGPxCS+D6DuPVT4f8A13dVC4dIb3GiK06AH63zEjFrYoGrO77KC
2QF1gzLdTdTUImSS2UTgdTZsKRwFDhPCsyzQaXWYyqCTEXIG9uI5C1utVc39SWXU
KSA1Dvf5hJ1IomBbqMMZD2oVZvU2BxVMtiQccWrptt7ftWnF0myY5CCJ2YXHoV06
0VDUezO4JZnXUwzvLrcCC/fh8g4yL7rrUYupAlh2nA4eWdwJrzHVZfdAaR4ap8Gj
6pe5PT/aLFSAwMNnP29E2xRD2HvA9Qm3TcgIeOaQwvuET+WMcKwThtGhS+3qCFU3
TmlwemzvRwH6EtZuWXm+5DydvgLgxnMMvFIBcAQdktZq2EbEnlYw8Sp2n2dRSjDU
DSDHuw6hw32kNsDzJlxQv3hIrG/bgNBmwIQo5ntXIo1Iyydd0Miu2lAN/BrvA8W4
CViv3Nvx5f86lJg9/XVxC9QPnJ9aq+0I8vZOvKWHGRfCyyDbmqHb/NzhfPrgHroh
snqcddW/5g2kc5oRNJ5lSEqdl970BhFj+I074pufeBUY32C8Wi0vS8BkvxF7H/09
iO1t7ral5i8tsv+0ngdDKUe8yaJrqu8ylpItgYmIrklTzpDytLTOw1pWOLztHyw3
8Z4oisdeyhWWygDQn4eY3wqZod9nh6QNSMBK9kXILZgqtELWrgUgC/3J9hmmdhb8
CpNdyOVX+nk9FOey4iu1i0sgbRSqk9gsbIboouaGJyEdd3h+DYDGBMo6gairSkG6
OTq1XVw+4tAWj1hnpCcA2hfoUcp6eVkIiTBcaoMObDlkRf0pWMlSvjrpqOaz6cFs
GRz0tzk5k01cwGQaJFfITcu/v5dIY3kncJ10Glz7egyObRmFiTV1zowmRJriEIYg
+RE4eOq6yhi4koL9liPopLXR6KbNFpuAguQAdNrRbq+D7Y0KpKhULPT0WBpyvKq+
jEvT9thRrB16E48KySfjJlm65AIHgtZ6zxZh2Zb1dzcKxXNHS6mSbwVp74+CSVar
Uzd3yCPOpbFTLCFtc9lSZK0kAJ8z4YXQy2WNXX1CebqfKcgNmL8UyEoD1XJ/1nTR
hkUxWRCMYRbcjB75UrnMrP6JagA/V/QId0zM9fWEqb6YOFB/dkz29k+LiEpWB+Ys
gYReiTI/whfR78xSbqn0zFGCwdVgBFw03JKlP1xb/BOFZJxm1QL886tChVjuqM84
nKQNbI4IqXSaPR/7B7RXz+FD3GliBq05ZdPq7kX6yXcYE7zUeMQVT71Pf0sYhBdg
AY3T2TgdgjX9F3JVSBe2r4uqHBHmovsweypRAdYMUKABX7kSzz0JTQCv3Bsa4Pdg
roDIx/Yd3aV+cIvxS2BznhHEgypIF2K/wp0j6G9xtu1t7nvRDPj1vYuY07jB9Gjv
ftCQLQwLR7a/wcjKTEE/NUJ5gHMlFImRRb82BnrrDEcxqmxvHrix2Fo6VRMfE6bQ
zS2ICW4dwJiCtE5Undlg4DZ/FFGoHTBx60hQmWNjZyRv7xgP9ABL5tf6AY6nPwIo
xIYmyUmTxMWRJfKtfBhbCyJ1XEEfSw1nBdS8J3Xb9dWncEsEtUje93zH/b5awI3w
pis8GI08AeJwcET7ht/0115X2w2+TDjWsRNkPX+DGFbnnbZD+EHVzL234Jk/gZSx
vDmnL6/w5cnDN0vW/hk6pgJ66AqRGkWKpDm4rdSmWEQcVg4taG/grlyLdhSd8oU1
qDWO1MpCFHjEjDiu7J7PYxDnSwYdkj/U/HekzvK4pxF9xuG6kRR7ocL+FXZMoOXi
2DQ7NOEa5NIvpK6sPsayJPlt7KTDql6raV4yXsD/N4zl6OpKwiHYUKLNDj151vCz
HIPmH9rpYHmpfXzgmOWNzOC85a5dzC3r/xICV0KTzMqOQ4g/oSM6QGvTD+a6oT6+
0Lo/AYrz8PUauw35K2Dvk1TvK+n6r9lV+1i1CgAGl4qy7t5syaoswn9BsZgwkQw2
Ozje0YtkBPkXL3y0WW8x/lq15CpWMqEopYPlnvS/sC6LUH5+TUdo/nrUi1KKS+s6
uhAjfI1f4332byKi3TiMqc5NGKlZSIhRoSY1ib7V0bi7LgpcPan485qz5AbWTQhH
7PF1OqS5Zlaukxgpe5x81Kj8q+muU48iok2p6SVpC5PQTLNwllfPx4KpbqJVJihM
+fKR7NK6xiFIq5+dSbKlHqm+5XqzSzH5Y+9cr8f/dd00qydNNDsKCpKvbvrLBnZ7
dLA8Sgc3Bjhsc+3Irr5bIEbhTDpvuDULhtEQcxGIr9hN4U1/R7k4D0I2Ysa63gQ3
sXFtERuvvvLEf3fXcSXrEGgPw9bIsiF8rAUyum/aJzhI7VddAVL/HIFpboZX15Fz
FM7G8mCu2CHe7YXWQLY/w+WY0L/O+tm/N4mwp7oXA5fQ5IpkWfTG8CabXcqOrjpN
V0UOwBFTbQktjmOY/mcUrXVS29Zj5vdhFRvqIoWMmOmn1Qygmo5UEOLljXQ5BIWf
RCHen5a/Bd5X47BkkmmMuRcIxq0Lk0wIG095WNMEuRAxQFgICQE0yJZbz6xQPM+n
RoEq2xD6zsgC4eMOs4AmnrGtLkf/6DJrTxiYao7RVsK910BMdixRCpKKMIfbELyv
60sxI5jQF+E/LfvxNfq85sezLl4qqvFlVOmPtWU5ksWnh0zrHs4dpOt8lAmPo/WF
tW3kIfEewEM+omQ5Q8Zvo2QfqhSA0XFImMvNUYHCWIJikoJM168VRkAjYo0DUS16
BKPkcCDZx5CnM9xrURNQloYLCbdpMgdKRQlQRHALaqN9IabKcRFXu4FMX9xAlkBw
28QHBImQljoGUKKZcIcy305MVHNYca41COKMpGu5mpQvnXRM4m/rIq6CIpwtisAn
vLtJz1X5X3280eP5DoItscvCRelrQfRuOvk8jWNnSWPcdV02Z5ZllNncEL8sbBCZ
1gmpAoPGfU8UfdO8BQVRdh1vh2QQDHbuaEm1YijyIklfgMhl9MvvGmSd1XRs/FPf
N8ZggH3mky/J8QDlh2OcrS/Z25EdSsrAX3LhCvm/g83g56O3/EUlYPafR6LdLQlX
tWG6qECN0oJA/EZG/KO00/cL59uvKaktqoKORLVLZN7X+KMe++QlKWO2IHm01bQR
Latoy8APrdWAmVvpE+TSAm4q8MT1tXkON8YvX3t3sUG/FaesrVRZDWP3dCpN4T90
Y4aUkXIoXrwbcAarge8A6FmoU9kTamrRtdJhLolDoEmb8h9UTzU2oTQtFACaYXRE
tGh5EdK8F87Xxqn8VyA/+atY5yBbKcli7pgV6U33tTq1wE++2CbvO5MIWkLiaOo9
YEmHa5h42SDDBZtfPKacoPr33/Qkocz7ZljSbOh+yZpS1vUvyPizJ4TToOtSIHiR
6XqadAleGA4dQ4iDEJZfDLip2PbIdrcu5oA4U6KsWGM3qC2gY16UqfrAEHQHN9Gr
ODQQ0Ay7yYA3Z6Iy73EDmLemycocI+z60iBLxbjOcfj7VcjKcOlr558ca0n1ZJyY
ETgp1dSnoPd6BU3nmiW06VhcgRIhsS1EBRh1kTPG60BQHwxkV5aJxFlRwhUDFL7W
SION6yro/dHxshhtyIsyCcrV+ot5u1OoAfXbUUg3M7vMpyds5Vgmy/KhPaHhESK1
Eaqg8IKdiF5+tdvADKgBKMjG5Ml9N6VE9iPmylinLjsjcYH2YbuUKkKCfKNQqh5h
uC/Jnks2kcMRtysa2yyVi4qQIJaamC8hHEooCnL1NFfULkLx4WpdVfKyRorENmTh
ndpIZOblcvAmAiwLg+pmSYA9P7jBAUIS+x6etfcF39X3HyXRr3XCokbkqWWgRVsO
IsbRQ6pcadnp4XGFBOT/qiCGaANj+kipw7pELi2m9nfpr29VAPoKz0KGVDrStE6O
6J4WQ4IvSyebsq6zuauYXhl0IXPQT5WMlhOfDqolR7fHMdKkydCLaE4XR2iODLdX
fxHQNmlw5I9gksLQTX7aDdpeO7YXYl8YbrwP/Acwaz2n8DrZ8LquQ1GZE5u4p3FU
gOo6wiQ707/zEYiAuCPhVGMftkLhNlNs5Vr7Iz6nJEbd5ov0Nwg/WyZVHHRpLC4a
tv+JN6XJCKWWzAwPRsxjXxnJIHUNIiluxGLfdM4Vn8J1ARX/o7QACiqi4mzvIAri
SmI2Zh2wxpNfV5l6DU70eRyn8EcJPYbAGJjbTu62/QlXwvAmBRyjajNhxtkdD2uS
q5jerLevZRgCFCrKjspx4Ah1yVREdgsGp3x+z0HWqQWmddLWYicKzplwmDYzDfNv
h9+By0e2lCYswXMCgRHQ98RCcxjnNWNt4e1OObRs2luZs3tfS6yK2gfJrYpp/SQ3
J9V3enkdP++zb6LZLFROL/pouGhYn4cL9oPM9X4MmNhCS7dxDp0t/NkfbS2MarwU
GBjp1aGp/9KJJlC6XvOlNA3gWsglpLGgEOZ3FV1XWpfykrqqvMPS1vCROsLUEhKP
OKwtxFdSTDuVUKWPtCw9sNIRFD/WVGPcbTs+zQpp+XOSfvXFCD+xGxEWTgyiHMCZ
SIi8Sy+ar1gCLgsXNjyNWwpdhMnYdy4h88MIHQbxdkbSSJUaEGEIuK/4PRecTdB3
sGPRvIx6ewEeVPkUxe7TyAaEEpU6ARvCULglGNnOz9h1Elt2xOJ+QtHR60m8eMmT
K/BkNqb7KzjWQfGDH89cWne9RPdqasvslNVrKtwgNO4uvHXLH+2LxvD7LTwWOlP0
XxNPGuJgunSoBlGL1ngjgvXnXMgMZ2wJBxssW1OA9WLnuNDcKEbVFkzzSejS6lbp
o3Ztwy5j529PSRTq58Nl7UZbFBmqthgdW0il0q8HE1RFoC58+Gry1ck6E+RTZBTg
EdD2s9jQRy9LlGxJRxd+P7WAVgIlxSx9jtA7K35EkK3Q4HLT6Ir2/PlxehQcesYm
WK7FDXIovH46yMsAEE642w7J3G1cgqlcsCP90/JG3F2T/5EL38fEZtPuVJOoeV/O
EntReTALHx7NuR1eJwQExPDLshFTBNjk9rhJkxnPgY/+69beH8WYOqf81FOtoAiU
dUo0J72VjbQvtMEioXIl4pSTR5IEiCSWDltbb+j7cmJHFX4V51spg46zhLviioN/
5tRPVI3zFYMWK6HpvsToZJutSLY9l3b+XKbfhIeBeSewfPGUHV58Qk64txW1zbCD
WDOUqCozdtc/NQVZNzbYgHsFDQHRlM2ir9fip/LTt80QodFCk/iBVpnh12tXR+pG
I8sYaEMzKxQqHfFgkQWCCJL1en6pcXvSsMJkq2oRl0O3BZvm99GhjG/atzgF/+BS
8Kij4gnaPDJqZPOVieLtrcFPqwmoV+YtvmEML1Gswu4ghS27UG2H9CHwQc43zMZ0
GU5Cq02irGfHpZ6f36ZnmD13B4+toOGHoRZ3hfcRoD9LB19UB3Q6oNtZhmVWo093
QnnBEQv8kGJqc6JgeV1XJFqtM6s6a31ojomKP/4NxH6SCv582fsL4FpzidwX7M2t
EWTuzrV0yKDeApdOboJGQFK9/oCWhGwY6k75ainqeO7g6055zOF2U4VuopYMJuWF
UzDHXH+Y4rQxzKNEya9hIb1MAEDCG+44FGDt08DaB6OOzTq2YFlBYdsaoPsOO8pg
zd6mH2l7hAFaetqi1zBd5OVVnkLvl4+UzN4kDPQBHyaMX4vO+Dij5wrL5AKOWEG5
PR898+ToouAAtcCyMW+eEEAV1MThd1uUlzXXAR7PUc2Mg5bADucjWNi6xH4DGg5r
QjBYGuOAAgZTbSV7+0PAV1lM3DjCQ0FeKifhz5l8XsqZC0KjkrNlLZXjJxYzMdYi
wnIlzRMLwCrhC1j3AxgG2bFGxxja0AGDK4gjFMFwvcu9AN7EeWW8Nf3XXlwMxMph
5OIee3TXkBRt1oTscPbyqRTBZBy1Z4aiHsYW05OTm4CckQ3KizHSaGkTVsRBZts1
N2hc8MVgA5ktE5aTkw1x44eUY2qlhsLf/IeMMwaW+0JxZv59lav467xPpxy0mRdf
M9Ld9/hpEVd7jN8hMabVgSk2/KhHCU7ViQwy6OFwu2m7iNLhbVtcWF2ICRhp7qDk
uxTpPAQK5RJiY+oAucW6paWzVv0oy1CJP+BbFbmX/m9VYAz4mmcguLqvMQ87cDpt
3O7lYoTk8X0QwAkcLW1u6CUC3ASodw1zPGLFw97EWVgIFi/+tqUWmjLI9+29D+Qm
lfIOlzYUrMpaPieabXUEPNQPgdtoMiPcZ07qkm9zRHj4w3+PP+OWbaITYSvRFmlW
zWJtPzm9NyZYcgiLG2qplib5AxSEkNrQ3DjxUD88nfec0mwq5nBVkT5qovQ/gSFm
l+U3GD27DefCJTOifIp4vyCdvdBDzZQbJhNAIt9TLoLDwu3xFX1ora2W3ywtttyV
p+enePia0ArkzSNFoI0L5LIWqJxOQmou1KJkWVBMAzZd2EX7uwn4Ix0i6ktO9Ir1
hMtjPPlsE0qqizD8dltv0VqwyY7NpYcSmShi//6um3dHU3aV2sIj7YeVi99FDMKA
d9LYbWgshGC3pHn2CXdkITUh9VGbK5jLgIZB3IPB8xmeGNBLFagbW0DYXn131ROh
QCHnGdHT9epSBCLhCyiFEjtXmv7WlBl/InQac0vJpvNWuc7uRixYHxo5Fkj4Qx0M
+DktaAKdPrkqLQCX6vIWl3E+TVcSZnjzttvC9U0rqc3OqAXUtgYTkcP1SnL4ZsOm
CQoCcs8tlHDpQ7Ydu4EqeIG4I3i0ujWDeNF6kqL0ny2Z4MB8ORCP94xhJ8xcMvCq
sE4c8/qSXoPhs8XrWJHyPx28rxAEboy0n/YDRGkpVyW3WGfh0U51uY1ynQunG6S3
vsdNtiboGDNWZbsmFIOPhtizydzavmbRKDwrmlhyNGMb+lGoDR+/r0LIJbjfc+nz
1YvtrVqcRL5pwSeKwLSWshiGzcCMtvOKQ+YeyXNeOjR4Ygu1xmSzAGmaiQSAbSlm
83NTMRsSyNY/+Zmdv4N11Bad6JvfFkWhjO4LLe7T8SCy4IPLcn0wZucXXBbmdXX8
TDfGBC3ZPoKvxnzreyiixNNNbD+Kt9xfTvAEchkTHctS87E56qGm00CaDgv6pTkh
JF4+9IBkGhy9Sy2wz5t5QFz4NtskSmcX8W0QRXTL1qN9VzVdn5AR07hOPG/VWoev
0V0yBKEcs8qiXQe1NFxfSWEl7rvtW0Hh5kv/XuRG5/jgmTIDebJ2j2zdgkqhl3XU
WVU+ib45BVj08oYiMU7i1Wd+ac/4LCTIfRM2nK3B7CnCpt/HEfkjUBK4pWwV60DS
x8IDq3zHSDdGFjGXor38rJdWUCoP4TZXiOX9zbCctlIUKGiWq6T25bedg9DuqEIu
L5T/m49jBzY8JLXsaE+DHDVTjDWjiSWSRVdfbhNghhIFRFCz1++PxIfy6F85HAvB
jiRZqPmVXO/blJ7z/5/14FBlYmhq1KfZ5i7Mg9Jma66pv6gsMNP0XfptKFDZ6bNF
Y/VzaVCWlXcLrfjWvUThslKRDF1IUM/C5fmFKkX3nHwnox03EEWucLRsg/mKJ7pG
eDpfurJ+tPE5wNJNK9pPaYxbc3aVJPErp7WxqhpQY3YxWPkhVP8tDnXl5BmCooxg
gcTBJy1Xzmvj028IHbPBedJShXxgm3jcbqsx0BtcRbq/5vpZsM3ymIiHc0J3G037
RgUEjqBhcOPLE2/tuFgX3MB3WrH7jIZ2Hp7fG2AfjQmDhn4MpAGREbiA2mn8opei
FEMM8Y6enYnuRcoekcHhCIrC3RfjEsEW4yqQt2RiUAjrXWB9OC86qe9MuvczZjkJ
QZ09wsHQjzj45nTNRFFywVOwNTFNOqWezKtVwe0hwA4aoMaZPpxzrQpbJsQddYh0
TlHyEkgaCDAmMk3zZo/oNp9CkzJHAx+LM4Qm9pSYguHgCo5y58KVIV42j/qcUOTr
6r8kahnRwSDx9wgK80XuG7/2AgkyzJkNxYsca1+zM+fwx386XiOHg/hk92G5Z2oV
Q3fFh0XZr4svQ8+y/xCMJc0QOlYcbtZKpaM4X7PPdcqZ4tKDyc5iegABwd3pQ/O3
9rj0piJgqajibITLdFkDzhsxjbTane9m/i8Gk76ehBzzWgO6V8TAuqqCSseMG62w
WPJ2QIep+fRrhMosvavYnER4pFOqrGdXgGz78oDhl2Tz6QzlnFxK3y6rQ6EH2Ftz
rXBpbdBkcVwbdyWtlorFClB0mZzmF8r8llx1RU266LP1eWK2TzvFecn6lmAA0dZC
9m5rehsUDzEakYDNjPfoQvB4vO+ooJ+Bg5VgqKNgGfJDTKyPD0jrroWUzZA4edEi
OmxOPXnM5ntDXGmVEK6ihFhLTw3egRBz72Frm4yO163l+7ET7ccgNUUVmdGmpegq
elbwGo3Oy9P69mvif+MIlq1xGcrUMWxIaTFyUYUOOCanKHIB/kbNcpjaMpciHTQc
xcmr7hzcAdjcqJnG1Sq//Tc6YpDx4Nh9xlwkm2NUtmU4EWoaeF3MBVw0uJfiMK/Y
FBpB7Ljb+nwCbinx2aoXTSfr7p1eICM/MH2uHHz8plG4j+CU3RzlQq1eng2FlI2i
8Cwc2tjTizWFW+7s+jO+e90VhuWGMvm5xSMoa/lfoBfMbYn2RPIEnDxr9/a05KTM
1056WLp8RPUDlgfEtaQGBMCFUOpdqo6yoQoER0ejL/8NwfO7pWcNhcsUH73bMxJc
XkCbrfaCWIckBAgYsy7AB2LTNzlM96XanuBVP/EyLMFOWujZ3e00Ve5mEgOoy/b6
UytqH6v82BHdmByr6Pt6jqtTrG+v/a6c0cu5pOyGMiys46DRThdMe2/5YCQo5gfe
4aMW3J0Crrjf6zn6M1bDkIKMwhTkKvupglnZgBWiClb/vzLU+XoQ1FGp5rNcoCtE
NwN8v/IMzWyWd60uSD2ueYBEgVoCwGuhdRdKEPUA9mMnebYUC3DBz/wYPkJx1ZDC

`pragma protect end_protected
