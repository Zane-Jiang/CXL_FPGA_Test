// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yAmSKJYuUCmx736OX2RNMI4OCp54D1Aj+V9vyU+Rw4oNDqbj2/SGoXVESsLi
fH5aCW6pa+TL0UId5cGve7gy61P4LGC2eerbSyQn2UkC6UfPDiwV+CfmCizt
03VXw6DhvacFF+zbc1537U3vAo4XeuShA3ya0ss3wMUolwYgbZZ3uLlQzTP2
mrWz0CYjDYysuccQ+gQNnYKVYAi35SlloaosqeGCNhYOA71ExmGIjyzdmT4S
MNMHUcw06usLAAUml03ywlA00MdImKHZKa1uwEsbbObS47Fvkcyu22WqKnV/
4svomSrESGbpgmfwArh0p4JJFQu2bB2q4ddtGq7QZg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p3f8UK/tnWjNenAGTUVl/rXxLLNtJsIroc7DmI29XAYfZOGLmEcNF56CTdAS
VOpUVCE+twu0P0DwqYK8BFEv5KxkV2jIWLaH9/h/Xkb3S/TyqVYylMNytPF6
7/O/LiQRd/AsrS80OeBNhZ1bxeEAM+g2OYFgQSFqb+OQ28HzoDDgc/I98Nnv
VtM4Vf6HradKwLcTlnCGz1R/3x74U75vWU4ZPxeF9wmUFebyK55mOrk52f0c
8lmaFeEtqcB7omghZn8dcprQ3z8v1iONY+UPH07pRrKvORq8/TdPvn4qCyEf
0cFLpN+o2s3S9VpxzvIGfG2SovtoDwRME78xwYnAUA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WKVwXzUZ3Y1jOFXHeULiw/GMBqJ0weFmCV4t29MCG3XvNP+T9kU3bZ/MwYnY
wfmEx7LGHzXBDkwaooKsi1ppSOia7PDpcMAif0pBwzsvytAe2HukjpHYBt6D
+EeB1LNaqWXZBrWCJ/yyL7pv7bzH+cCSvfzUczm9itSApLnSM54dO0YWuMtD
EcYsVGZrUgK28T2J8bO6dy4JEBvP/5hL1XU1AuqPCjjSc8SSRRNjFx3WRCrB
jxD94cklsRxEKB1FZKRpmYNz85thUO97VCRNLvefQXeYwffSw8WmHoG2AtTz
1oG0iTrTjfiJYEDcaQHawnA++Y8YXClWG17m/H6arA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BKt6zlvhPaB9r5PpnV0I+lkLxncQwparNijBAkpsCD/w61g1JxbM6O8Jk0EG
XETziZmDZ5KV5x1l/LFlpbTtZihNsNPf9PqOILlWXqCuo9gNE1xNa5w11sed
pN5UQwyIqYjmUuyMDPyYpve4TJYaW/LP8GuQU1baB2w2q//43kk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ayzmqFyHmj0ST9wib8//2sRZnyK9Fn8GzxRxx7SpqrpS+NyAVcTEbazMbRKG
YR7EQF3wHhzah3ZfNfS22ghtudbizBwPDCxCfoG9PaboDYPnpiRlJjmhxgdB
/bNxARUqMe9vnd9fMNjnO1u0RD9YFlwn2zdqBgVtOreixgfRjqXxSjJpJSNm
eVRWnUInPcJzoROs7PJDJzQzD1tb5qJoKd/Z1BP/KFwv/RbF0K562O6zigIo
cNkeE3Bun4xTRUkF++iJXj5SrLilqrTW130mi6lu8TUdBPLtdVVBY05iChEz
4LYGqcWV1IZAunjmeVWnQ+GH6RtGrlBgLOjC9emXZVbZMhjOP9cewOb0SfgO
q0Q0ZsZZdJZLqq4p1CHwB3jALxhFxeE7WKCZUMAomPoCaNNCniJj3aV8P+hk
hrE3y3yhNqpjYzTd95NvDcfSNx9tS9xcbjraNKukEB6/e7577SnebM9ft1Lj
6IbYATv6UZggO+f19istZOEwT9xVBc7y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aMp9iIJgT4WI1SC4UVRkcLle+b2RtBkNImkaEvmEP+pzAtv+I0ZmuU0fBeOk
yr1n7AFQuPA5BFxPz+n0lRk/9Ej6UuTmkV3bMRMRM/C8wRvf4BcBXKRr9Jsk
S1IyYC8L6pyN/XA04SSNvourb4qzF4EiL5bw4RPGfe7F6dBbAYI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QaSajnqfHtcAeTvW8PyG1yPM4slaYAwP6ern861UrVRXcdnQOK1pK6WJJQQp
W5kHGZGQ89V+xJWbHBCcFrEkfB1/AizmtO+wo1aDCde/d55hPX+R2nonDOyI
WYrW1wAEykg79aO9PolNvlSelsOJ84KXBv8YpQtshZcOzVHQD1g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1392)
`pragma protect data_block
gAk7dsjaaqWBStrmv5J6xFI70Wi5L6V930Q8lHO2FN/zaUJ2MnOwxAA1tcEr
qO0RQ4wnWp3lGxYmXoHTrMBxVe83NcRLEjRB01mJIsEzRSZ7Puc8p+SaHu39
p9qUs+wXoZJXJvtP92icfB3qs14UpECbRB+tWtva+SXrNh5ATmvNpK5cEQVR
oAt62QuldR1rbgr9MA3+skpKd26u4vJLbFqHQfUMs9SbBrEcUE4xT8Xk8EIa
Hb8QqaUUPfGRgD85UgzzZDzZQtTbvknFbB1TXlxI2uCgrEbV+r+BTyVhcFri
HtLpDrykvVmU/hoJFRncY4V2lHXf2WvFWEPP6OH4AvlTAE/5LVxPVgFwriry
ftJWV9Vj+/eBV8zf8pfx8azvCvBoo3gqlDWzyBWNAUji5jgU5bTUz8a2t6Qg
d+ils14XOCYwBWPcX0Y6/7oTk78+z3FVYBSEFPWUS3iEsgj4QO8WHhAPjtsD
b73OfhQJqgCBE1MrCrrub6HEWkdSwAqqVqirEoTp36mvkZYzVhVWpEX7U0os
81bxKjXdW0zUveV15Cwp3F72alvMXDy8gp32nEBxjG1Ha7yhqp++mrnT82BI
CBtfbxqzVu16nNX4d+bGeuLaQ5Yvqs5XCzCY0b6QlBTUEphJm4FHWXXu2YJQ
QYKCZhMFlKGOBzsrhmouQbZPD6mcKR6r/NcBEwmK8Syfl2TzfGw6Rr3jGuY+
c54kwQ9Qbn1TIegArWlczmtch4c5lQh5qEC5WKVJr/pMsiDhOOL+kZ7jGQIA
r3aR+5QMj6o/+uJdd3pT9bL4EvkpuxPYjNKd5MkP96GVpv0TCoia3PzNNTDm
Y1wwvszJYwYDFm5T/bUwAR9rjcEvlMzjfzxGsXxkPQcxU3Ep7ZrHjmViofWu
8ckoyq9PZ3z9AqMWhm4yRkaNHIyecuqEururj7wS9yJ022evSb8D3Y/NvNgb
1YFNR+708I5jpdv8epTxI14GtVNDBu0/pVLjGmr0Yl0pMZK1Nvt1BgjlaSCu
yRi/ltXg1l8cYUGCkt1Y/4zKngwUaHmHbfGqwTJM0rCpVK3TW+TbnCPDddx7
nmpd4x4IyDs4hKQKD9/uFvoOmzdXIWf4aSGSIwZ0d/ihZJVyAhdFjMD5NojG
OtKMbtMaI+v+4ixhGTA5iwQCtyjx8fGaEJnnY3gIjKP3I+7oQXp83rfSIpXP
NsNdQsm7N2WtBneghbCe46G1Vao+mjmsm2IRFXLt69fGyD+qKY/lCCQgclHW
h3RKqlGj1+ajr07+xVueSR/JWatwUL4m45a+fyeG6pmPPbQ+YY+TGeixTO60
PEKiX0FolA90noGpv3L3gBPc75jv6kQptYhPBRp3qToOKbTICSSDHVypoXJI
ybtBIYBR+SO5JzYEnTK35qOFCw8Vvt8SQpBNHyUIyD/MXuQ/hrmU5rsebXQI
tHWb8B+y0IrbClQ2bktljRCA2JBdTqJ+E3KosKHyMh1EHfKBvWDygu05+Yiu
zgOiiT+2CR7vX2m46iuQJpxyak6+/YZ7t9BkI0MGTqTZMHMUw6659igjJfj1
SGzaaTRu0X1MsNJntpLOt6RZ5P3fQWZLakBNLuf2tj5twMnlFWxU3P9VCAvr
3xQNObIdAO/E/iQELF2EcX2hZDy1esENPqHDdSn5w/IDq3R/D9ZKr3bpSMBK
gDm+rewJu/h5QKhQDVHQjq3Ce5p3MToi3TgbQByYN1ylcuNIV+N5Xktlqfsr
vbBwIitNk9w8AxhN+Gfc4zeepPZS+WMlNNE6DkOkKGa8nm47meM2WNv6BPH0
GIc+51RPrqtnyCSt6ENXIf8nQokyBLwzZDmAs7yD+6/wjV2OA2s1wm+d

`pragma protect end_protected
