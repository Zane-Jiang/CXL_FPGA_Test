// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
7oWFLJCfvwHEigLWieW1izlJZtPS+CK0Hnj2lm56hBhpe44oUAQP6WCtuWkSXF0Z
WaAJNdysRZALojxK+KzCxSM1ptSdRS5xQeUhXDVdnZYu8KWNJyWNdBQ0IKaeor68
Sqv7pyqECTepnVawEziazmYmX1pnlCaop9z9q9qeKnlgOwGdFe676Q==
//pragma protect end_key_block
//pragma protect digest_block
X6zFXxNoUm+tvg39uzRaMI/scSY=
//pragma protect end_digest_block
//pragma protect data_block
B9+TJpBQsm4PKBX3e/v9YIySUlQqbVa/R/JoHnz9zBj+VF5BLtTtLiM5bEPdQVwg
pg0iFc6xcT5TX3QB0jQy1qFTXPJMSfo4xtGbEOe8x6z9p64hxRcfqWSEL8vIWfCh
mWybCKX9UYHojo/g1CouqBnFXoimWuaojF38B+SFLtJ2HvKWyd7GeLnITtVnqIp8
IEbxrCYT5zIlFCjLSOg4WSVx+v2hcyKsHoZlkOoElafvE9kWxcV+altMvYsMPr5a
HUlsETq2pRpMu7BaC+to43eOKtfzzgxjOsVUJoaBZmWuP52RT8UaJSJVn+1jGtqC
gQ4ayEewzvE+9AV2FAJrL/lAC9QyKqKgpz8MS6jBxKttvLHm1eeV6lsfgCJlDwvI
iD1hLheZM/WAyoDYacbFavoKQAyouZX5E8FaWlx1k0Dhx7hWB1b6Rzdp2TVKrHM+
kPGGxpZOpO+tFE7t83MWoaP+UsKP33kFU6p1HoDEyt0ieD8j8ejlreT+fhrqrxQX
eJiqZHAPsQhN7Kf0YSh1GBBA42eBM5s1ZRfU8mVI27JPRQJxUOTtL25wuRAbnl/Z
uStdAayeW1e3HDLKjmQcsIj80cxSl14L7GFuRuvysAx6c39X0BVy4VahxCpVD4de
evI4YR+Om8VU9NnzI/BEEw1h3Nj44utTH+GH0gkWkvjx7MPoOeCL6hhdUqtmAepv
/3Buv6la0hxecI4vy2c+zIaUzXgpUjnDl1J06wBLWtmwkfrr+IY4Xd+ucZWGwley
43NtXoGhv/kCDzKnKtQqPMN31QVDhxhTlfkvOH88DkR4V9KTweJ8s5Z+lYiQAZIt
LI2WRJuLQ0r1aBLJHBuTn97x6c1uneISVDMidmcMIw9grpUpwXPThl9KKl4tZHzK
QPVbwaEOfj9MSEgLloASnuB34ymmGQLIacbpMmQUA0UsE596WbMvyNLd4JZKEgLV
t3a5X185bOzxBSSuIXLRnktHezK0pmtk5WdtLy8xfhyGeOjOH+oMEoVIaR03x80/
fXCqvDI+v+nW9jALuKZbQn7mhr0Oahv+N3YmTRDhZ2Z6Y/x+WC4EA2cG9gIC4yUl
+b0/gmN9+7buLHAYzpemMgxI3VTbWCU0M3wBZdyA6t4uUQJEkGrTqdJ8lu+0nDK9
6P5CAoBD+74rdyj7wg70l1DZg7yP4dI8FaCIUJMlqfHNpFh9+rXthEDu6tEo98+M
tKGI0h/YnkHroWYe0z67Yf3f1/1NBrDkj1qILxLDkn29jWrRIjL5cc/qyv9lbVbP
I//Ob5OtYb6mCTonU1Le/dHgl+oPra7xfVwhxB5MqJfC231tkueLQPAtvdcf1cWU
MYU/6Q+19u/qf57eqAzUuPs15Y+ucjfCGq/7kdgDwMJpEbfh0OnONAu2PHn83wYZ
uEchAEDWM7nQOag4tkKdheM0cbB3IVtqqbdDgnFwK3pR6r8GzTTZ7JTMOFeSyRtG
0pbmq5I48GQBcRd2Lezlu7JeB8JWvX//s3ccPNnfhlcY++nkt5tCTuxOgZ0uFqr+
u+MNeMKhvG5laYObbYq+ILc1tT0eWLii+pZjNZgmuEAUsiup1j/8MJoQyzrV7Tzw
Q3O9sqEbbx9JtRxsSyYqFopkaLsdIKLHQCmvdtnCsmgexFgKeyajV64kEyH3OLHR
2tevuMlrRLUZKJ0Di5djWq2BoeILRlt8Dnw/KR4LlmYP5/wuByZXm8EQlt4kARZN
8PmiUdCuv2XuTInIfnDFBn2hVxv4rCd71kLfCHlW8BwHvIamzDFmBeFkKWAyg+Bp
BkNajtsc6ugVmyXZkLrGW9t24XcVJCPPcqVSX1Up2ryEyCyLtea1nv6nKoUXGh1v

//pragma protect end_data_block
//pragma protect digest_block
mnT9T2H7KxGqG7abwvpnpXuSsmk=
//pragma protect end_digest_block
//pragma protect end_protected
