// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
nvBLqr6fT5mmFitHxeEUqoSdxUMzGEKlY+WIzaVHupsIOX58S7Hs76cFZotfYmFa
4B6Ie3c+rzJFsEmwyVcRd01uNTd3anPUR2A57bwrfphvQjDeJ26S67TZwvisC4cA
9vEh9yHJhCkw+q1zYhD5QlUuBaYsNc5Suhw/gL4mb95OVlQl8dtfOw==
//pragma protect end_key_block
//pragma protect digest_block
dYwXvxN8lEGWh/kLGWmtpimRkZY=
//pragma protect end_digest_block
//pragma protect data_block
Z8hGG3JY3tBJToYQ3befIBrOkjwDw0uFexhR92jt34jXIiofJqHiYAV7wWCMY5eH
dVB2bu7fH7cA3ViFERrjqE4PIR1S1rC4Ifsb+RWZle5m8dEFizajwNxD3HIKyTG1
LR+rHvEzAz5mzuH80IMUkbaIbOMROwCermPONCspTzCYDwsfxt/3Rv3ExgwOOfD1
2NVOTTntr1YDek3rOwYqoo2KdzIGOy9JZjiegm6fJOipdphJmmd4FRdfmhEItV5l
EZTsMTX/ehBdmnmG0HfE/6uGVd9hP6TZXVXUmhiPevzT1lXFgApMlRcQ7oJltDLo
xw4u0RIoH+HLIM/zod+JxJROWdyWrYD0nFbFLhclQ8Yrjf54qQCJqgBBBy8EgxDM
zhr702a2NOJM+14f9hwh62jyz8upjzFOL/lYsSTzkAi6jfiPx+j9koJPuoulFOxz
y8XdtaDpsa4NYWPggbhizozzZKw343szawFPaup/zMEzzEkodnN7vS/R0/DHD0Y/
HPqVyLZ2Sl6xE+d5k8WG0nRFQMYgYBGvKXP6BbWqqCSDlwhnPnzf5c/0cX0YTPMh
g5wSUQCpITJsQcCsukkPzpb9uIUjjBGQVyUagDQNDr5GIfHbQbYdfWmktD1NQEXi
7KByfc7TX7xqVj2JRwwXVslilKA4x+NBOkOvjypb3wP6oPPSBkILaKdNr+cO+ThL
rFwMrqrQF87M7QGtr32OwPD3pHz3QMOZZSM4S+sliLc4u+HlxKU6jomagw0XcJTA
wvYmjTJeDouAeEuCZ8T92l8pQGTD2Pwg0+jv7E2GE1GcsKSwwGFEova30VZXDyhL
itGe5d75QqgJVKug82kSEpm3YCyhDKMyjwtfPmpxNJq96KOrPQioxPWshiNZ9g0X
X4K1ZMhSa2D6NSf+Fz+/1o/7XFf0ImICVlOoQ3DMKrc/qbzxqOtWomGE7GQJwJJ+
ii5YeLCUc45hIJyJV0aCyGPUFWcXqneVE+qpHYnmpxJAtGAddEsRAjpqS3eiOzqK
XksFHYX1gBqa6Y4t5BOKhwqJlcMmvItSEZSfR6KQthzkK54sxXaXbEE+c1LDBHwE
N8Nf5T97/WPnRLnCxrcBtldriZ9WuKi9F+Jq8FMVLuL9mGdMcttdWzNyATA9zR2N
l3IWGyr6Dd33j547aZReKj6ciVXXdggswhBzTQAgCxw8R+dK+UVcH+DP1RkSaHHc
q7aONnTBH9N1jvohGqZAgNZs0lmbROexE26gJXm/l69kY+pNtDA7dMJ8BxpE7kVR
jQ/mjBnQeFSRoeJmakZGYsVoKaA3f2rEkPuHE9DqcTsuPAdqPRKxGJA7yiGGJ1IK
Aiz76msWxizNdjnxh+XpK8SOYfftJbXC8Bp4Xb4/zJ4gOanNSi1K8fw0xOOSVCup
Yy4iKmcUN4pIDZy1mRjWMqtN8kQbRun42DTkeq8qd9Ypl7aL/+EjaoMO3pIFZgZV
2+j884/JQ6gAZPxbfF5zOLhXWWGI/wShYYKLSK/UvK2D/VzdtqANCDZUyZFoAklG
wr48EaP7/WoFEbZMZt1DpEeKrnszEFcK21pyHbSuGwruGlqiMQ3RjRNwdvMgMezV
g6wYpobG+7gCG0J/+nj/qn4LfYRGE2uE1y6HWtKJfY6mneULMCq7Mr6qmDZ4sGLi
ZMEQS+CB/vccBfcHgbjX8p3L9Bw8bcoX/kW+xFCB7m4fh338+YMus5tCVSE8A0Ej
F87H9yDPk6f1yBGgzq4zS4gj3/O9CmyjQLX/67E6xTtGowD6Vz0wpH83L6TJaJ9g
yWZ9P7TEdkutxY6EaFCTVvHvYgpMwDCfUz+6tnxna9y92aHBJy2uzU0ZKQso0qW5
pRnurD4vOmxM1+uMOrVB02Q37Nwof5z0xT9E0xtec4cjvsMXH4Jst9SQ12WFIBPk
0REFLBbib3DsjuB4Zv5/DZ0QpySRSB8zPra5rue9qCY+p2x42sV7r1sXcluD/J+a
WSFhQQgcyInr2Fbc+ndvOD5cE9ljTdec77d2OBKhQasCFIGNTBTl44d4Zmmj9wLH
XGHTjSsepGgejD1BPdd7CZAtDLvH+BhiLkun/Th8Xlaw4Y7cnnHTEmLlb5MViW2u
dw/E2ekI4ZdCkv1depYTxMvqanuF/BLwsrziMnDl3xMmqTAfdJfykUQ6EraHGmDe
K7v4yUCSAFQI7cf/GVnQXQ0E8TVW8kg23kFv2SD+GzNYbyaUbr/E8T57VevkTpIj
OSZDnA7IF/hWworlU+RleZSrJs9Aajml8s9SRYQmarNjit9grceeDVuLozqW66le
3NcSQsKxkC95adMYrexMCOhmWRpYl/64TK9NTgnRzqJzsrYECtO8KvHzUHloR+K9
F6kbYelVQfs0PRuwhx8m3a/kk+HsBE28q5umf1rgNd/MReHsnuRaPlq2tbmNrQ4r
cO6ZmiXdGtzYT/opUUU1zNIVLvqmaseIrCTbWa9RFpuIjWJsRrKZq95FIAH2Wgsv
iHs2EnxqGU1TSuJ+wbIU7Y+ZhM0QFbC+sDSPvp8tUPUO8oVBgNhA763wUzFhmwyx
6esWugCi8AOJFg14PXuYbXLmqqcQ4XHM6bLNQpTEJf6/QF5d0Hpn1ozuZ9H3Ho4t
cthLSQPPBJGsCaBrf41y/LzIZPxZ3WVVuIkjaqjponskGVbszlkLoHKVU4/L7mTn
HRHpff/NupeFAcSAwKcrdQj4wPOrvuu4V1ebaKq55NvLg+hWXJBo4Vbk7yEp+6lY
uLKwPoyXZ30FMczygPSbZNhvC3cy0l15kBN6aVwS5VYZ0MGM/+S22nRCP4qvR10f
sQqkkJ3qOZyUfbRJ+UPPxBrc7BfdgDWdUt4NVJE2VOsZyaTL4tpx4S2h7bp3hPYS
tQjEuXKuCKMBRaaRisFtncSEGtH2K5wV83JIJX8CPcUZ/zLnWdQSQ5AQuWf1fY8r
lNiHPTaYs5EU5wPWLu3Qf/OTM+/iIgCuvBrOhlTlmC5O/nJJf/J9MW/ncU47hjwR
XVuMOgU8lzezBqtbN+NfnfhjqnF7gEtKw/tBgAuraQDMquDvTT09kHMGEFsIteLi
bRDulkuyxb+L9uS09uf5QIs/cN85nxjD4a4cYWwrViFbTA36MhApNm0ND+Ey2/9D
yZkbaTJ5sWuOSomjSNG/FAJQyh+FvI5V4YgQa8y2XkIkzB2aZ4HRmTNy/C9BnqnP
IEE8QJlXNDDDhtrwva5qzgIIkEgVIZEzlsE1fagDsPM0UCt1Bc3gaSJ09/gxpUWg
nhI8UN239OilsDH42HMkt/sW5SdLen6FvuhPlY6Wj3CBI2iSiKGh2w9qVX1JCTY0
qYm13DXSbjJqN0Pgz9zjtGYZpkj7HYT0Hd3NQIkeM6oMsA2MWouy8NcAw7GqH4GX
TEY6udJg6RY0P+t8YMJdI+FxFPhFBRxGw3APHnOVaFY77yKW2yZ3KFyjotGW/Poh
IjwHtOLq2DroA/ufKmfStiR8d752wDaBWVWsiYuEDypugbU+O1I9U2tFKk8WzplO
GGW7MI6nP+zGqe/8ZwrXcFoW5aXcVi+PrqPpufDTkMY47G0/pzvIQMoF4NmY5zxw
N1aHA+eB0tUoo+AMUd7iw335QeWX3fqIZkNph4lez8ifi26gTMAFgar0ZJmQJx3u
/GI+vUkIBcONDvOF3HZcnuRyICxDbdErw85dgHLH5kv5xO6gvu0FR+uE1XHHbNM4
QMeoe0ASwtHLuoy2MndV6JofcW9qBPfiY88wQCpU/5Y+iFMJzyhSebIAm6a5CRuV
+/gWZSPZP3x2B5G0YSviLqflXYRhNcuqaETgmv642YmAOzKZxTPGqSztIGuMVJ25
bFXwZ4Pz35ReQUdFlAkFoQJK9JmgeiHrhMV7JQrDBhX9F7jy85uQoxGJoEOIPW/G
XHn7R97GlWUUnPKUx/BLf626VHHkntFuz9lJYDHhu9AoxNW08HnP03Csbyoqhtf3
J6v3Ale9z4XsMBLsSm4zme1wmhq33QkkJ/YY6XFSCa337cMAjI3sgd6JV9k9PRvh
eWV0V9tlWb2gh2XY02TINtp1JVpIV5d64AV3LeL5iOm3KaWlOkmHQX9RL7G10um2
UIb8HEADtEGX9wmua1Y5NCh+tX+ESJmi4uOZuldgqPUeOdCr/w37nCbyrH5QxZCv
qyqKDmyZR0YmDpRh66osHca99q/p4k45X7oPdIOaJfVbsPX8rMNHKbXeDcsipCQl
bHQWjxmzoVSl7oqBsN603wi/4r6Wr+CRl5Uo/kBOQXzUHSysyet05uuksc3WcEfq
BTZGuLdZQN9BQFBfTMMvQUSzOklNOgMuP+8fuEdJsmXwEx2nhkVT1u9N3fqRWc9q
KqiuEspp1l8L2Q5SS5zKSfVGvhZ5bfv+jE3xfwcHUlr53GwUi1w60KZZTuDBcxvP
3b7r3B3HlkL7QbzolHR1wPkuyt63TbOVfrLawj+htv79GV3/B3zuD4FG6gzV38yS
rAJHvK0aAtggRqgQkZZPL/loyc30gxsZjreLzerdwggDe3PpU6qPS73kJVNd/QE4
w+quT06WvYGzHy7d7y+s6KjHHKDHpR7dpWJz8HAa1w9sQjDvb5uSj/CG0+rz/Ewj
o/SLu317KmwmzAa+9/kkek2uTOwnDZ1dun/NxKGd2njP9rVpQXk0+0dwTtBBsMD2
chNZIJt7i2b0gOyZsO3FNperKtZD6xearmzmwgMW4iuyyqyFBR/XEPHAASO28hEW
5XyVdm9aTUThAGktbbJ7CuVVugOqgyr6NsCI+Q0zphOYBbWZN7BXRCF0GSLFRKIX
0lb1XBBaIRc1MMBRMCpuGZM5t5RZqvDytD7OAhqNqE/FVhTca9fFSrXl7fwlR5kw
vd2DZxHYKxfJdMuGKhc6Lk5ZKmf/Aso1y3S8R2Kyf4DOIRX2BJOIoAgXVc4WdV+v
5W6F+WrAUnlDAuexpYcgd9Dau3eyy82ptcL5tBnbMFOHIVh6qZcNjzCmJO0c37Cw
OxksNL8KHBpgJHywB6mv8ZoyYFOy7pwGrgHVJP407G73Aw3u+CCDH51KF26kzvot
s8cFQwQBAvZI9dY7YtjCaU88AMe0Ew2N0hTGu5EXWF4ID+67Adfe9cB3fg6tN8XH
tkfDGeJmwHmqf9hdKAwUYOIcx+vxp50VVMNOhW8HrrEBD9BMwGkSsIj/wmGZg6Oh
NJ6Yp6DUFSg0gryJr1OkQzoMaWqHuK0Z/99TgqIoSxnh6Cv/WDlsnPnj/AWbm4fW
or+lwnEBZG77XucTRqjEkoGqYG8/dcgwujTvnS6Z8LZ0h7XAp84eWdAQxIPvbsSj
LNO7X7gWbZKvLbeRsfIRC5K9Lkcp48SPX+JWIlyxnLrOzpQ0tstpZVd1urcZRiT6
69J7mCsLtlpX0O/Cr2l7mzHwrQj4Nw4SiAjSHCy/Fn0oQlL9J138/bUqU0jac5oQ
F7Mr9RbtPCp154Jsz5gMuNw6jZSNNs/dsgcxiBM4xYNgJbGSvYv5Eiry4KqF/dZJ
9UZgLAdKZ7mxf3sdDDp/weRh1LW9RUuVBqfGAJfLqueNE8bYKEBMupMs/m45fw3T
2wItlybruv+7s1CJJmSZuzhtpIYiYN46kWIo7vond1lfWau+wFkdhS7jBu/xoIVk
eF4f6E+Q6vCwXkkhuqtoZbv2N5XMlTnRbSfxqvzYoLtsOW1pBEgCqydupcm3tw1f
URoRQmDzQRJWDOCvIy6+cNDsO9NtPoSLk6edePVYvPQxh4sEvUQLdTNoL8BzJjQw
3SvzY/8UJXw2SDLnKPrUgE0I2eC+9vvkKAmrifg9xZhVy7S9iLKw/IMumpKVMXRl
XI8IgZb1Lsbp5yYlaN7lMJZAQCNJkfI+iUUq9wWjbSnew8EMQwc9ONLixhDf2+/+
4VglKhIWJen1+NMW2QvKFFiBtwP3Vo4ot+Pz/8+2JajS+Fjze263mKrgKP3nEZgg
ehGPNQSO5vTw4ymXz6TWj7f0ouIcqhMbu86mQ2PsGGkqoDfnjTyfKERsVdiaYd2r
MWIftU0urzUu1m41r0peikwbq9uc5UZn7K24sN5nRWOoUUFeOGqeYKNV7SPIi9xh
3t2uYeN7RaPwfXAhVXLcC5km9l6uH9t1jsDZW/E8l8eptSDPDuvEW8J8tpnGMXpE
drImW6WI4FN5ieoEx9NFHmwt41hRE1N6ocA6YuxMYJ7YUGg+fgPM9iCYMmO/i/7Y
qVLBiZ6WamePY5TlCWO3KUd7X/Y87rm5VVi0iFHacT9xWdgIuYqnYUmxsWO+68z9
2ycBZ/qMNDq+BAaCwPjTU4lz5xEGKoZLfPytO9xa2WtXerNsSaB7nZOt1vhN51IB
PdP9cmUksJHuJ5M0TDEEVqECoNmzsiTggrEzAct979eMw+oASFjIUqA4nh+NIkF6
acp771WjCRx0dPCG+Pq3bSHiybpSu7dHwDGiRRljwcF3eUlgVvS6jIUOwrV59r8I
d0/EN/k8IIfWFsR6FjfJBpIYl6jX7XxkWrkaz9G5HSHqZaRElorPUp82MrXgwWxg
pQQnaZoNYPGWVKKCtB3CmLr0hMuqC8Oci7s/gS+HuSov/n4r4wfS9bJoxgm/5o91
4VCAwOFWXXn2vedklcpZGUDdZiR+OQdEhkTSnf2nn2v1fyhk8G80aPyjrRLYgS2g
9+fNCwNQEeXuCI+03n+GgSFwXM+M1pYepUJ5sVMqMnmCfcPT5QeRt16ezDFZ+HbK
0gqacUr+9DdJ+0Ng7Nrlc7ENkGwefE1DADg4gVFeRAk03Wv4XveGh9vXdgj0rUZH
nOH5UlaW/t3jj0ilvoHa72CzfKaiJAu71gDPoB9xmCdqhH6TC5ihUAjz0XqzE+zm
LaJbiZ93of6g9OFjHVtOi+9jQxlRGVzQfWcD5pisQo6vBxvkEv1yQJS21qTgq+zR
HNhILG0zLUAylAQ2Bom9Jo6j5yU1U4Im3u3tn3D3nQ0bDiQyamZ/NqilNVYdURt3
GjiSldOulAjOCXWyptw4PDyuxMPJ3oSWNqwbZ9oVuDyPaPu1GljqM+P+xO4XM+T3
O3S7UksGZ8a4bfNg/PhJxJXjRwPtcmrkUyUXVQZ93lIYaTDDeJjZYjkcE+cIyd49
hcd5vms5uaV1N79W+BvqMScKqxFsVzojoUGFz2T72mEBntuqnfQBzuIe41FGzy4o
LBUEk3rv7dcEni7G+ziK4A8mQwBR6lqEcSL0hvpZyrykdCkESETLVR/n9iw3Luux
q5fierwMQy5cK+0iHOP6fAwoyQHiCBThZRK37p96BkDJX1hEE8B6Pv4eP+DPkKUM
KiD1WH5ztuysS36DbtPFdVrmqEAdNRB+ssRJMNqX5FDdFmeVq/632qvXFhlO2t2s
vtHpa9fkitxMMnbE3tYcLS5QAXIaIAnwxAFokB1A0h1V1aRquZf6NlzzExGIv+Mu
lwq+BbfiXauqKbhXUCb23Flb7CG2kjKAr1xuZkjGGWV5qVyNUNuMXOuus76R5y/l
co1b3bQHcwHYC3gIc6tnyPo4+KAPU0PzqRzyxcrOEXcrdZsir6D90Tr3mkXuZGzI
evAQzyK0aTNrIcAXZkNU5FdwI+vPd3XaT7jQj3fjXZWd/BcQLfHscMKaqYcaZ8kS
d78wQ/yPl3I6vhebvfBOiMH15GjXeSuMk73bSgeXUYZeHz776XFF3IztVh/ZqN9b
GW20E8tkv0MqKL9of/DMndIKxWjXWegN8l7ldc8ytt3bKj5977SXinXCqJYUd0cx
BolWxnP2QUObtg7e7PinDFawJiC9NFIN9TvqwctNKEROPJAMfcqlPb31KOCreclb
P11VbA3sMXrxuF6RX+C8y2p/PSKdirEiO2O/lxevF+iH/FZIA1zMzBMFUgG0sq4A
twZlYasoC0KUd2xLjC/EMkXRkV6iVVXOzFueY8gsDOVSB0mRLmABj8ZektXTZX/3
lw9VKqUBy3mh+j0M6cNUeCiyk747gzLjOJJ0pwgsvpa6jp4UcxLtlyEpCIhHFjmZ
emQJes1yvR/27kZkrT65ICXI1IYjw1fSWQO3JV56q79gx+TfQ/u2pqm4+CjK9Q/0
YFzK7E4uVTEEXDy5kk8ScKvi25G9WRMT3Pa71k3Or7TlZUEyZ5AgNFBzD3LqL10/
2gIeEMhBJHcc18jR64qZUiSaxLdXez2ofXTezbzH4PH7yvkpWsn/nGxbUHi66Jr7
y/4MXDqHex3e8M+uUBWech62kanc172rwMnIjOgKy+xtibaVmjpVmRRLV9fld4id
N4N4m4qm7X9NOJxfQIOzTbBB5zoCjLADj9rYWAS5pQCEu+t0NAvGYDZ3pCD3PbLz
QgCaa41aKr6dQPswf17HV8WckEUcQm+6RWcu20OfGsBYDbTSPOO4oxT5+XGJvTgA
fIuO+KGBPP8OKm4le0Gkt9hc9sfLDdpjK7hiiiYReETvuhr5wQJmx2dgEi+1a4Tw
mo982FjD+VqA+wwF9qPbysKynd/Z21RZaquom/aKncGvL7iE1/mDaNP/MszkDhrC
kZocq/3E5jQ1zO9j/A1tNHudsAJqgweGB5bXdKfEi1K9IcrO/L7D30nxr9I+/Wjn
j1lySCt4VHPsH1gG5OcToz9YsIjf8G4FRf/s1pF6neXijI1za/WGu2R0s4gbD8CN
PNGTWLGr3TxXY/vLijwxAVpEPtN3mWcWYPfEMv2PVlmbeh3YFPH3wXwiMV1iEBLT
J4FBnVpfEPlZI2IlRDwe3BoRrL8BUScQvhVtOc6dV2c8vi/q0FrynqobfgpUmq4P
waIvmyW/Q6RidYFOLV+QY+HwH/QDIpoGb8VHl0erwGYt5uigzZt1gXTvwEZ3vQ+4
TXBiqBkNuOmlrv1WOpkFM9HVcq7BI3oaYyzL9lOgjblqwblMObBxejQKqEtI2Ztg
S/pHPLfrBRXjy5s0j6es7yRux5Lr02wp6mE73mdH0txdLDie1lt6ZLgAMsyBISiI
jD3Zg+HebHMpbTB2Iy3mT4Yoz2A9Gc7PDJsDJOgXGO+0E0VX2GjxO5D9ohpT+MAD
kKue5L5oENx95D7c+jU4jjelKD+cYy1WigcOnFUB0exQTJzzMJ3R7e66Vt5KFrh4
LgsKA9uLr1F2jOCFbKmduXKrYqhPfH3TdnbVYLjhcSFiwj0ragfQj7Rlt8FNZyBb
qH65fKdmxlbMassNzMxL3bmKNB1yurI3JjhVm1314Ij3byRVHMB/RjvQkapYoaLF
9SePpY1mtWV7JBn1aIPYJuR8xb+/3fuELkyT7mEFlFEP0c138CwSuFydR2YckvEH
Q/9+MrRNeo/Xj4QEvC/aT1vfv0LCm0X9MXUI0qgRRvoepqc0SMMGCS7Yl+a5Q/1f
g7OfOG1O2n/KECSEqKwexTcZ+Y9RxvAqyjZus0HoU+iCUVCinpQa7zERrc0lKka/
nO8w1CkGFxwv/5S/XqA227XXOzG7Bo6JrzkeYq5QkGpRwGPah6bU+DRf39e6Ees1
yr02i1xI4LZyW5C/SllXs9bAUfztW9EprhXv60+d76qyYW2ATQl5gA5iagzPZKZk
dUBnEs5v/Y/cdEi1HfC/8/JVJsHOhiwAoUwB6qceJe7KBhAk+X24npgFnFQzHO5j
2jIztPMvvQE9zNVPiToPXtSy2QIhc6jgzBMQufYpig//H3Dd7sc+bz3aTdIJVKzM
NRmBqhc5/gioXYw3SPNkf2QwjiE09dPAfQ/BEK1x4DfrGiav4+RtbfGvNCtB4qes
8NXbTppzM6Pexwmv2bvIczRoySNprKnM1szLyyPFZXDs26o32PC2h1Yi8H1dF0P5
j2ruFQw8fA39rIKKUwogug3l13pzafMxSEnr4fHcnc9s8cus0M6xq0WokgRGq14F
JKLORqzFTrNoYnJpBO2Bo7lHC8Sqn8kawPAB39LTQjowntRV4V7rKU+xqraBl4Nk
vxxEbF7g/IeeBNhX+S6eeq7gw7qrHU7vhif4GPlhjiBUdce9WpFCB+UWhRnBYgaZ
9k+vvdypRJZr9y/hkMvpDO0of3m2pkeRL348T7Oi9CEKmjQrTm4sChKjRM4drIis
oXa+DQey7okIr6QbOM04Dgw0WbpMt5PE7Qa63EtTjEWxg9O2PLGiUVt0GoIV5PVv
qNQF4MrZlb5pkBd1ozGl7gYJlC0wGPMbRVK14APFM2lqGIb6vDDRUCEZ1FT/6yZa
VTcq+1hfyhYZgwrHqYsrxQg7qIWL0ouoIG+AM3JeOX+XKvb5OzzbdsK5OQJozkjW
47w+ImCrZvTGyTwKlLXWgzfMib3Drrq9yT7RCxSCpkX/DC9Z2TxUgg7Ml92rd4SG
Pm/BZTxocEy0B0ROO8/34EX6vkMKVbtEaIdqoqjbr5kxlCCkvII1I6CC7brVkNiv
brpF3KJr07nisc5ZSYxqXDRqBjsNRKn5GpZhq0vlK6vV+s8vtOFCscLAunBS4Y/u
t5baMiZzSTL1K9o73Q7olPWmNYsjXvoVecidkfE1Ilp+ffToJ2hZ+jYTpf/scqlK
wkOylGJhhpCuZpUXU7Om6D8L1Vsj8C2uQ8BeiLrwaJ2U34JFKubj9g6EWCFYXSel
j9PtKqkwv1UDcle+ZetFMmF53F80tnhi7WyldPorWYjYpMcrU+weqFY6abWHpAcz
pVe2AegBh4XfevyvxUAWGfhTx6hZ3kw1ER+uqORi0Q6wEwtf9oxg8oke0TCmu0ov
n1Kc+N/ts2nE5hwKT4j5dU4JcmrljUWZUFnWh0XERy+3pVXqoAUN5Tpx7duHoMUK
mJ8+WxAuq43NTs1is2fGQkQA3DfXSEdChyTV5efX1bk1Sg/Vec+aPIQJk41sCMoc
6aZnxx3j2IIPZ9lSVW9MotDjf9tpE04bnLdo9k7sqNUpsj5t4qFC/xfQrF7P5yl9
tFiCf9zq7RKbO+KSEnEGwpcjhvG+VWX8hhOJwblLAFZX8JJwbXpZO/s/szPRRxbH
XbJ9XU2YIvpreRHjMZhHgpKdUEF3kCJrwV4Lg+IbtebVc5ntRvg5YN9DfaDMf5eN
0/HsEqCkNC5f4lTAXS8bCvFxJuAnuLq7AfxsQ3LWXkFdAN/60Z3WSv15f9VIwEGe
P1zP3YIa4sXmHwOlOFabJ/Nu6fBxf/OXqYbFDV5E1Vej0xKYXaaw09fsmLY0H6rH
D22V6/nUX+U+zusFlJ6aw+QM4zdLBS4eeLUA8egajvuvyRBo1Zt464NMRxCxX4Oy
cC0IdOTKZit02wBWmn0PbSvcWcIQN+hPnm55VI9qiT99WIURgGowmksu83BfPEGC
6iVZf/qJZf8JZkLWNBBfAZB4ATKXFgRkvEOhYqV2gWmDJDiSEC6c/kaYIZqCn/kP
ObBvmP/D98EZdpv6kIuW4X81i8YYqq6q8VXroLsQ1DDkzqvhE/JCO4zNd4GVX4QT
BuG73ul8P5uFVQNCjBSTBCAiWZ41HMFud8iYXCP6ZUnhizRpdwm5gCfMLOmS+2G6
z4Yej8axZ6s+oACNPePEIQH9Nfv8Aqmvn+0ZkBe/641qqXI5p86E7rDLphY1DMgX
srzC9CjeqLlGVLOk4+DI29vNn9G9zaHiEq5vGkUveV26iSR95V2Sp8W71F6Tumar
MmCIOtnuPisybzEI6NTOXr0njULzfrRRfOp7AxU8osIRipoM74Ydq9uFvBUo5lfK
Qz62FpJ9EGmMdLA965hcoJn4TbkWt0+ed11/psjkwlKUI/hWxjWnpN7Mz+jN0ebs
SjqvbK5LCSLbXcyn/ovW42zK/AULiYPDIrew8bERrhydAT3QeZ5ih8omIhAZEOUQ
KZSLRU7RX+HNQZ0huTGJ4UnFGc4alCYs41vkXCfC1kIZcehIHrJsf3TbxOek1GVK
HO2+ZwV28TjwR0ssaYtw4e2LGeW8EjIcEQ6TusBNVVtwO0pNFU0gZeZP/4phcIx4
EqpAEuNIAMwNYWhGM1Ayc3GB07A1cNzrYNCPOAm0Nl4vcWQ0DR9vLTfYBgNQ5s8N
Zj+aoHOO+ocwbNODdbumn8/Sr3yas96b2G24CmDEK8Lp7lytHguGT86eLTM5daSo
dFi77QPdhyGQfj0VRM6gZusqBsSb1FaYGPJl8InYZY0rac0Guv0Uu8Sp3LbWSvom
fVKa90pryc7kG9HsN053+0i06TR+U9Q2ygE/EDPaMaEQp7dJ1k4tpEbiSKNP9LLa
v3JmdSQQ2V/s9DBBg4Sgm1P3usawYhRs0vqLaMreZGVLnxEue1/UjlFauj6vAcPn
QzKR0BlLemKL6fqsHY65u0IX8zNe1hyjd42WG0k+vYSEkJyiz0IUdNLQmVd+59Cu
LNEJKQaUu5Gpk8ggtAKGj050blXjf8et9VmKRfYkolCqgBCH5NhPbpF878eWUQj/
niR6eshwcUZNF3H0BXGeUyDCoydQWFVHet9wAbZDZOPpqyLjW4Wq55pCo9Ihx+iz
PbYYJmdsKUanHbWDb4uU4yJFlXU1s+bEYqfgTKVlpe7e5H5CcAm3YldSmKTXAiJV
/hH5Z1eOBMzw01WthO/F2coqfBFGim0H7D1ujXmbf6fGUqK3i+UEUejxR+L+4mG8
PMgVRACQS5V8usCxsjosC3zL4Zdds6ZAZcBCHL6599mp5d6HXKUygkG6KYharb1B
edRJxiyjUot9MWZIGWxKrgrjaNjr2TQDzyAxe1NCRD90T30N0EGj8b5wVg8qeEdU
nMaDT+GsmiM5ph5y0napg/6no2WeG9qdW+EoOWQCw5pUNehOIfw8J1e9lg39N/Ig
ztL06Hmdufcu90JZjzLoXqrEu4kMmrr2riHejdwNg5H8dE92iJmrS0mG56bYeQoj
nGxuQWqYpzDwaF8X8nJ4DJv4LrLvbtbTDOiyEv4sMCeJ5Lqn7yu063gTXTSzTblP
JEwyQKUzXy9L+CJqrQ6VizdCNDdRGYOu3JLrkCzglFJcPkfjjpsfllHPTuwtV8Mw
YGpdm/SwDwwlBdtAThkhX7Ce8SGTt2IOPnsFXoW48YX8DV6zvj1Lr+pWnAsBsayu
9Bvs7Zg/GfgNrj5G+qOEkifKk3HQkRpLkLwREw6OYRFwGYLwbbR37zarLffMJyCS
IiMd+sVUKCzwkpaSKudvNtHls/ijEzlIyG9uqjJnbNOhMfSQYG1rponZH0hvbgLt
h5I5eg9fEshT4PiRwVXKDndjvyarDHyuKyYTZbJotVAGelCEeNwQHP8103gTTmV1
4ZP4RFacVlY2Fguu6Z81Sclhzck5DJHqdrigfstOy+b385BpEj2lZP9TIaOstJJQ
VyF5bfmXNPDnKxHbdzp1PE4WhO6W8h5O+YcQcrJ5uTfVJs62E2rMoCXRRu/UfYds
VPfiHjUAplz3A4pP1ueINWhOuh6KOGrlQPT0h1PqSlyDNqDTgYWhR/E7s8qIQnOk
YKg7KsVYYnBPf0x2K5+crP//ZRhUz8AmJTyAYWyDls5H6l+o0rEoFywNYh8ESAgw
sF8uBpT/kAUwSFrA9uQgJdfh9Il/M0WYcpiKkR+2UrX0Xg8s6o99B1Dj9ObIXWgc
JPb8eKMor+sJRgcxOBkPUpR+pS65qyysUZjNm0Qjuxyp2kR6AJE0oeLCen/768Ds
8xE5Fmhh6tdrMu/h2fbtR4hOnYy8sdfOu7Q6uJHsqhgCjDWdni4eYZyaQ8CCEhea

//pragma protect end_data_block
//pragma protect digest_block
bZyXSYtrDu2iCKTUIskkmf1f7s8=
//pragma protect end_digest_block
//pragma protect end_protected
