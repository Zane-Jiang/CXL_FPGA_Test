// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
37JhZvYpm4N8gpNsx9wy9zFgGKzRpQALv0RtW6psLU0DbBrSOHtZ9xueT1AD5VcV
eCgFm15Gx7PxRxtJsJnxD7rXzGm1XRPLDmVhvVWq9tigZCNhktZPa34tMTAUSbDq
NolQObUs4Qj8ETwEyMyll3joBuN5Pwmah1LuZ7OgTKD/AGA4haEEnQ==
//pragma protect end_key_block
//pragma protect digest_block
Y3YB32WyyhVUfqaoj1ufvQmgYBs=
//pragma protect end_digest_block
//pragma protect data_block
VQPbRmo2NV7STXUjlVYRJpeJwumA8quoc47ZMT9gr/q2HJ20mAXgf74xXaIULLyD
t/v41YJORGh5ftBJqwvZce8w55N6BRVxSZPF0L75DVSj1FUq9KmMkOduefDu9sgZ
6PJKBHRAa3bobUOlz2WBKrK4PqJ+bXTF6AtJFMCRBQv5vTPOd8LUalr540UqfiCu
cnCkM9UvwPZu8UwEbtehLMbIMMJjYLBRgLj0C6K/VcM3t7YEaLCrdFGalRzC0O/b
oXnGk57B6yLy2gBCqZtj37rSpZXianCSWgj8VCW4+eM8i3dwdGEMrOoouvQAfHMr
mqkdmO7brRqbr1x+qdLFQ73V5nPh4Bks/0HLrOKJZDRbWXn6GqRZLWHamJ/nBlxP
hU+pw1Wq96prvWafbcgyfAfWwwhSkfyNLn+ZUDQNLc1gsxn0gBUkMIdsKe1oOnfr
pEz0T1Be/1RcG6E1coAGHmkPAUaVLZLLDHe10ZBgtJkri2bHrIovQL/GkEOz+myv
spMNwTShHOfQAdesqOREPdpxEPZMGuxVM4YfwmMxs62lNyZbiarL+/QQN+7VO04M
IRomSsHFxqKa9WShfN+o/OvTNC+CyIS0vZ+FoIGEOCaDM79pJOoLSRItTDRlGBHI
IDXLLi0mY9QrEZXAf6Y2hQrFmv3bZLugOinmX07sZPSblufnu6KYcd1gQ7Y2LZn9
lRdiYTRDoxoiDrhgBNVHBNdniYqMkdX82BxqJ/NmZ6L4uG+BzZC1rToQ8Giyi3QF
2aKsBATUmc8iY14dzKyfSnykpy8zeCmbLS0XPiYQiVtQCGc2vgfnEhpck1XiiXhb
XGLs+xlWruBjOpeMyj1KduobB+CUqratDwClZiKQOPwGu9JcnYKLbsgM8Hei0fsy
utxX0N3G6DURYNWu73EHiqOO8BXysZI+5/eCp4l7HL4D3x47SvM1xzcbjT501kM+
7ioHhM7NRY+1SqrpnecZiu/9z2QSIi7SFNb+uDzT1QFDQXab4OkkFBwklOaeQJ+1
xjq4JqhanMiWWmzhwyNeqBI9N4tvgLVOr9u1VUcY/+8gmJHSbarOqcr3Qr4WBEzq
KYzpssOsuwz02ZHjsNSXZPNTaGEnuVxlFBFUClZpiO2qsBRk/4TbV7v16vBst0Vh
Cvjqjc4tnP0aDbAb+pL2iyklUT66x33gwLRv8Z3ZwyNO94Pn47kVn6nGI+r/AfpM
A8lZadiZM0F2x0HGXU7NFLkgPm9GaDsEKSzAB7FduN3FPYHiqfcFymkmVPxXvIjN
hAQ3vIHCvFZIGhNpUWZTVBF0a3ipZuEOXMH6q776xu+RmhYHMfZxSPOpEgbXiZok
8znRogdLv4BTUGFXuxw/SD8ymu6CTrwQUNkvqBiTkjyPsNx7nr5sXzYBr71F/3Kd
yQMjFm0q/WKUANm99CVsjajuKP1ppswyglwTp9kmZVEVBbhNVVgya9pHggfPfqb+
+4iNVUtcTGC1AmqaGo1PE0bH403ni55nxkE7SkdVe7IbwxLa4B16edSGc8phk9+c
rIACkXjf3IXX2l+O0qmsvsbtHUUP9MmsXTqCbyfAAwKaEr1ljveMx5fdHFHVIFpv
p2iC+SvYpp82ajPjpZEZowK3uwc0cRBBkl64mrSRMKxiPWQikxb3cn00t+MMUVMN
rr40PCRhUor3f3NMaoSeQhaubxPiPQvVAhCxGL3pTzvJD18OWONSkgGLq1PhlSis
vrJuqmDD1gziL4n7l03kB1R8Dd6aBv6Iqh1DTjR/DE4KshstU+MwifAhRaPPI+ez
6H5CY2D2HozZHl3/sKOUPadVar7xoeHlVUN6wexhbMu1J+YpMU/3YwFo51ZKHyRo
GOAVkz+P8fRecUUq8bcFc0ZiMQSsd+RamRVyQV+4p/ncUhYJlCKpyILv8tvlrqyw
R0LN8+njMeQ8CwfUm6ZJeogO4lOXmuWRtRaUwDIynP1xq+WhUYjO6AqSTd4MkBFA
JcMr7Y+JoihBrSIiDKh6jLHHiAI8M1pkS3MWVhc2MHWl2va1gbHnYgIXfedMLIG5
a6XBKVpyacq+s2BjyNBD616iWnLv3HkZpctVx9okLCogFmo/NB+YFSuHzhOYqLqH
ySrMKT/z66yYIZV1rDvhTbZNOT5etDIxYvMtKy62TGNpHVkJPSWQqd/sFhIGk2XD
wGflEwD/78D/N3BlgXm9h8CnABqlzdE3hHtM9Achj3db1COF4xf9Nm5Y2TdgSjR6
lemHizneSqUgRpXdKjOKr9+aT7rnqvwAJvE9UB8ShoQVg1dc4MxHyKKDGrwZpDVX
k/DRS7M/h0PHxaVcLpksqUzrSffcySpBZb7JrJEPjG95jBRFSAj8B4ZTzdW9EZEp
uKMzj/2jAwGO0yGbAOBssP3GNxhZF10ajcd4tx4HcF69ohrvAn05b+RHjgNGZjOX
reRT2eUdbhvnWE0UqWzuZlcUZFJVSwew3ALB5aiyqszc5Zz8/rpgegKtWX3T4Dty
IpPwyg+NEt96KsvSnKu+xGHwSF3xbum2tWEChH3siOAWDTphzVRF3uplRLqZO4Do
naVz9fijnls28qZ91TAlUtdxrIkID/LCDuDGKkHpzmP0R2h1kNalSIPGWDHm+tCo
/o7KuU/Sn/EeLg6Gbyuci3zvzydNXAtrhkiiUPMyN5Z+3+JfDEMj7t48M97RduCt
YJ8bGx2u22b1Hqv9bjYLKd/exEh8xyHTMTBYtxBEjo2pcoPb38/SMvMaAH6X2/XT
TE+7QG8u1IDT2G9CAz5zj8To1+LI8uHKF9sNCSvbxdW33y3pj0nG0TLKC9AiEZLc
b0FOOkmh1D8uoUsRPfA4HfuVrUjYR6NHbltjIb7GtCLRAt4bIOJ4fPSN77D36xNj
P8mFq8WbfAWc/IzkVSXK2OPVo+mHxzEL8gqiuNuCEsO84VnomxgVXXHnwbYsNtTd
44wl6HPvtX9YhTp9YcgFZYFfwuzbSV7FYcoIXcDmawK+m15smF5uOrP8Z4ssT7RF
6DC5cY+j+CPzt1DvUVGbD2whC3V1QkMb3CwMZ9c57lT6FhXRfTmkix6ixOhhgTVd
2KRAJ8QDN8jBiCP2bYaR98ZETd9gh71QAOSoZcYDCkuBVgKNeQSLVBQHLuC/xk83
L92wEOJHkGDOWa/6nPkDHwE+X0TXqcDDQuVYJDEGI9zJ9th7UTp8Kb+yUNffZvJt
WAhtIFR1qYM44YEr2pFTwoeUkhyysptYmALWn0dg0RFPXiI69T2VfcK6n7TnLRhO
CmPV6173tKkX5mvARrVf8FLdW1U+h7YqG3M3/+r8BppGwmCqCeJxIO0gtw98XJQz
LS3ISp/m2+D/Rfe5Fw6jBkJvVqtmkIuQ4KjJGg3afmKoQEyZg9eJJ5lVGGp+tQ7e
L0TZyP7Vvp8oyqAa3mVf4I0RHUXTgkpQLnNFndlVtMxM0+SrPNEGj3tcUnKX1s9y
/o0nr/W7S5ghquQmzkEuux/uIJzhMgjrB68NG/aSvR1QxmQqoC1SZXh9OoFQnSJm
PS4/qo7c0JV26wMiwzs2HJ9fJ6GxDdiqKenCHco25QYN7TpHoTfmuxB/n8lCMEzM
C4/euSmPZMdWyL9Da5pC3H6oViywH6CWGeaSPtrsH+9kld22eMTdqCL17N9e2iNc
r3fkHVEh4zvGu7a/J+8gdSVIXsnvaUTnR8TVbRQVD3F8ziamME2SRwMchvkM+jhi
vvmL72rLHEacJFdBkZeWKysLIFCptfKtsqxkfQbjbZmBwDfZSBDeMs0p7jz+er79
Dw0Ua92kO5X3X0g/oL0hxaiHR3DtjE8pv9yXR1X29oEo0d9LIMqiudbA8UKKSV6+
OMiSYkwV9uVxWDAH/XyAHoizEbjl1Y50vH1imYdSqYoY6kmM/lhlDxkpk6WJZavc
GqddSDzGUHS+biqWgPmKQU/EJfd34EnU7pMUixSeoyh03A9jUBBYjjRTkuVB1l4Z
y3k2gUl9aOfHIquVhe6/AELCfLIR9LAQ23PEvPn2+nYhXI21qBUHIcUtPX//bYZZ
PYQZFT6nhwwvIBQoESviS4+Db8xh2pgk/ueFqaQ+97NZGhK+o+ShYMKTk99gDblW
q0d1lDeyMPvYij1FkxiUDejV7mklBqzS5rwSg2+fpx1kL1HSQJDWCGuCpUQWhczs
8xaqtPP9NxIEmvs23JhdNJ5EDOL/Y54+vy9KLeT+GW8QywVR/e+u9RNwCgTrP8oK
9ol/VlLcuq/TYHkuj88eBu7yIRj5OJ+1QfEdo/aHQmzODFuKkumb/EP+fNDUaQ9O
fVAnghHc5TRU9OWkQeCvGXDhCDCIEB/tQKBRFLiv54dyxrFjamnJTSo6d2FvMzgQ
sFWdrOtXQ4FRce5tJJQuBZtl+Wx6WMS5ah9sZ8ctFGC0oNIhuueDljAZmegUilH+
ew8b1/E0fc2tpghHI+Gkt3rzUUXz7FuDhysAHmB6qvsSGkRDd6cQjHDDOHOJL8r+
H9zmW+CH+0v/ONnSSoyEvclBybthy+gaHaNP+Wpt7EnaXsUQjmMxrB0OBBjs0gcm
fsbkdhhHyWAHu9EjasTQENV9z34nji2+NN9vayCem4l2mamkytjxV/AaNm238PQs
m1PlJ1VsKOQNAn5TP2wNORIrGlWiF+DhvTB+j/mJW9TxH/xn6v1BD3FqZnCkfEjj
qQ73KoKgbYvF+/0ogWOsdvFwm7BIb6dXol1krKOKIRg96CbCVg24/5pr0lAXUaTm
4PWnIsQvmjRv/rJCItgIP8GXgVRLHwTwcO6rXLSeLZvYNnP7TYwytUGxy/CIhljv
mrTKq1A9EW157B/q7KCjHslsq0c2wHZ7ijhCHtNPis+zVnadXckP0MKmy4fz90a2
PdqmXNdSILehn9Z5cr4mGQLD3dXu0D0gVREo0NSqV8vAAJD1gEoSvvGu2ehzRjbH
PQFKgRkm7p/gjpbfZ/hHSUoSaXweZ+QS2a+IhrbXVuYOTTLh6M+R7wirWYbSsMbH
bCI7y9Khu1NqJ0z3M6q0AKrCwbQGGHyv2rjG8WdNl37/AptKWTBqzATR1P9rMRyZ
FkTBcI/hH6mPjvYFcsRKMXFn99xe0l3Mx+pq6HbxozIkN2g+Ht2U6NluNThkznkC
Ea4PRGgQwci2RwdmfUgr/yelS5Gvoysja5yKABsE/zU8kiCXdZxBHye+M46359Mg
C7NzxNIPSCpxIM1suR9G0I4ht83axgIOlQ5W+IqFef/FCL/x2b2/KFwaURhS8fWk
JWK7pBTKQWNPJhN2FxS1vUBeRgOE0j72L3URYme49KTQBdlFwa+QTdBMsr3b6HtH
Vmzs14NhmLWspbieF6CPCYmzuNShOT5i3CO8hehGAFIkR94YLpjp/zaFcMXULuOx
uh8mI4+tARULO6vY8GIBnw2Din/yBnq5x880IbARgT4Y1u0GHBqj4EW8TrhSm3mk
YbNzVQ6ZylSFQEmnPuQFyosPnL+nVXVuW0N5OV7ETxSOoS0BsEjfRGthSNrQ7JEZ
1+O5AbatqJ25mgZmXtyI2SwBcCv1jYK9bVG0F+Quyj/i/VZ6moKfDStBFZuy9OhE
zQ6lw1zsGGiy3QS5snNZpspjCBYWuGgGqYvVWlSSfpo5NzL/Gxs8hlVMTX4opgLL
RHjJ8uX/T1S9GAmaJ3K8+RShkPwgKZrnA9tg/DJJk1krGX2donPrWDPi2AONHi73
zoM16oA80IQQA3xEca3ULt24H1PDtdvc7KbqBmyNICbg8KWb4OlBNv6oOna00tF0
EqYO4VGq31ErjkoH8KGYjz4YJh/BZOs1B2YPHrgZOIsRUSn5Ari4kzrR1SoMjdxv
2rqbJvqCpIfUBWPHeh57LB1QjhVD4PkbyrBzq6xvAbWBP/PZ4Gq3Nm5IZffo8O1l
lfx1IXtWDm3hzrSnnZUKcDKdqqgk8NaQ1uiNbaQWCp8OHBfaL5QlyHLa0Rx+aomL
nzlWF7Ib9zdDmi0YgGLrHBvZCoRxDEBQ1GD0zN2lQOrEBxHZtrCLiFaCDxR3916b
k5J/uv5/ww24JlBMO3KKBMJAVHG4SXxXiLXqJC0InBxM7xKVJUgGmiwBy2PrZty6
MJzZpRIPcSoFwcdxdfvV/lsZOgvfpivWw44uDwpdbUWmPSKAiPmNVyYXV1eRscr2
1giRofH1CmWppg3WqC/AjpEBnAsemnRm02gnUAV4TdVSGpF2lTxGo8F2+7quaRCk
2HbpG1VYtGSR7wCEBzmDnomcFwQ8nUVUwV8r2jd/Z2yunHxvmbBG5OJ7+jpRA03T
uKYA5HlwLdB1pDraVWFJV4LKRYL4xs9t+Q/GhUP+q/XjIf2UVNfkiMsJrYUfWH5W
HZfYAQx4VaG36KkXHEbwTWNXcUaqE9NdyovwyehNrjMasVmRmmk0uAOYXbUS9NrU
zf+DciskzDKQ0DHTfYRBWWGra5KzOiKbFyUKWEIPvo5sCTJaGjydBVPmKtbIeOhW
K5gfXWdw2bDMMYKwFv7LYiJDJmC7x6FbSJ1/NWb5SKNPYecji4semUH7ajBoBTCE
Qw5Cklc21IvMDzE4cGZYqQYVbEzregSjXtkhmD6CtYDTe5kc31opgHUXZQmiulL0
eJp3rWkqNgFUt+/0eBbWt2nE/Bff1o0MD1w9VKVen7BG9M9bxjNDrdbJjxYNcgLQ
HZoVfDt2OQaPNSy31SgtGf+YI3pkwW8pSkjRhax2Q5qvXeNb9WjIzqn5pdUndUBo
6S1Y+Tkhr1JDxMFyPfqwl+dQAZrkQESzaUQSaES7D7jg0QTOtnbYSCu6eyS1N2Qy
WVHeuYLiBZAGpMpa/69oRy4p8PrfKnVHv6wVlEjyKZ9XuetPRyvnJq/rqzQShtK8
igwpHH9Fj64OrBLtnzZ2vUOkVkM0Flvj6f6XWVdHW1w4iPmXpvewM4Z93pnec7GN
YhEzfdoaczZxkwmSbrEAlD2ulP+yvHFqbxXzr18RCkVt2Y9vY6kKBHmF1QEOFYMk
uxsPSY6K2OQkArcLBUvOeEkvdI/RGIruFalUKNznKgn6KAKrb9RDCbuHN08P1UoY
ndFZ7lIHjC8F3nEbC9wnAc7Y0hnb1PgRZ9DsQWzN+GNNs1+9jmaM1aekrJXKTPV/
i4nhRtJQ9ZpnlbMUEmrfFsR87hM7GesXj8Y+VDGZiyiTpMS3ODZ2RL3yADAJ4/kT
eUVjDkO+SJ+BtUL+v9b97Gqfg5PKRGMhO6WMTkYa4g5CPC67RTekP4bu56aVLbLH
xvmRi+1j3Esx1kf/vdtRiu3M1pG+YJqm77DMPXj7VEWnmNXqDkxJfDJjMBghgNxx
d4F56KtubUAEl/+y+8YVMgXOKczwZlloz4gW9w4eQrYrC0oRBWF7dyjXC2uKzb7o
L7A25dzvXHMRvCJcUSnfjqrl0JYdwlcHMc5SQ5gb2d+tYlULJUesuGyzWTkss8Qv
SMUZZEqZjJXC4RvyPod5ISzwRAo3saB6MuSAi3WQ2+pg4DXXilQVngYm3kVasuLa
txkrYZ5EIUfzocl0kf1GcJdYKkJlzwZOKiigFY30ksSvYuZJ+fqpAvy5gdwWkwU2
5IP6B75FQLgcxgFFqP6SI7SOX5/GXXctm9TkqE7DX2pK2YzCuWbEH7iSk2BjH582
peXm8ntHi8i9a7ODrK66oC+/vsvUvEt/x/XBprkPdfSCvu7+6OklurTS+J7WGkae
4sQmPbCeDoTsmHmi99Krqh6KXnMGRYAzh3uzF+NWlm+K3GSEs5YM4zMkHFYF3kv8
rKXHlREb0VJ9kKFUv0dP3DMYKS/gihwJGSTofUAtJ0ALXzfDciw6tkIcBQIjCMHv
goRO5Y8tdt+SbsAf2O6i/LJwUg+QgZmevm1a69j+o2C5dsECUaeRzATsAw04e7vO
rYohrlyn3sGI2wE58I8cqNq7rBV4rt22MFOSrwEcIapqnRJ4SwLeuKL1DPU9voFX
uYTurDHhiux7ZAORWk0eG34zEw3aAj/sdTxmW/oLvQNcIO9AknGpdGFoYhxUISki
WOHB95r9ALuPmn/i5f9QtyoIef/D6ds/Ac+g6tL3Ru0gyCFgyYK9XsUxR6glSvwZ
FWlrIeH3901EtXVlzxMNHgbfv3rdThhWLtytqFggVfEj/IP70crdpHyZa09venLs
+Ezj0IqTaKM3z0TdgktwuNli8DYftZEGRkmKXd65S4xD9ImmkvXKd2zaDIpAS8aB
Fg5mEtk3huWDLYTdy9Kbz647TXmB7+D0fkapD4KxFXJslmWTy/5oIrORSPIc6jiI
enxHsLw60Jh9GN+oWlydq/HqGJsXuIJd1IpkHHerohnuqnXctUUFeMWkJ1NBm6dH
tLvJ5RuJYfplv5/DQH3sePxVSP5lsFi8XMSoW+0hPe7UaxHHfsPD4Ip3/JHvBsWz
vMORo+TufB4DtbNa6jx0psk9EfambXdsH6r5SJKP2PE1PTQlXD6bIyfuz/pnp1B7
9ApxH8z1RJ2kAeGiFXWkKGGiWVDIEdadRQ106It38dBAgHQP5ynyVzq/5MFk28gj
HJJlC6fRERlCSi4V1h5lIZ0ETaRbbNh9lmfCTtcCn5cTZfr/Dpjh4EE/lLOjeZej
j3os23oUbcqY4guHexjKbw9nVhNMLjp7krqv5upyJ6b234v8aNwEam0zSX7M03Ir
A/EhDkksV2sktsPCxsaayCCM/RjMCcAxfC6tb5mEvBbre7mkcz6ikqvEoOOy+cy7
WehfycLl3rgI0Yxas53wi8gYZ/73rxRNg5Wr1hSGFwnCBme6h5jAgBubaeWW16TE
njuxgZPcPnD87v62GnkomLtu6SMvS4QzpOSTsdzTaYFAGRCaH4nFy1HuwYWO//1b
49+SsXm5GR1G+bt6dlLWbzBDRepFEJil4XaqQHG04DtZh5rJk3f1xrOZ90tVWUif
6UAQwH+8xTlkMO/vexfPxP/dPK1OzSTBstN+s8sFh5RII55MBT6xs8Ueyc4mmXNE
Mah8/dZYkuxIbuo/Ndga+FUcGgygqIeUIR53lB8J12qQb2c8w5Rs2na4n/QS1DqG
EWR6MS4mzq0TsjE2BcSu0e9b6tAUxhUHYQ5Be+ZwGCimt8bhRKi6+APT5DjNdT2W
JImLR6LQskn2MuBG6WWunVuAEGvSBfPoLChpYlIjfz5ExhFrHghCJGp5yhEnTvQb
zAiA8dj4I+KUKkY7DPZkBhAh6JKYgX1EkXrFvI+tQMW3ivOntr8hhzLczITGUFOS
YrfMxjHA2RExKHuYRO/g+XpxSsoHg3klL8QiQIvdUQJ4P1mK5gw3XSELF1HSv4T/
loj1LX9dr4VGfe9gqbjcFiOK2isSp9VU2QsUiFYInrjpDQ0Sblp7JguFANwbcv1P
21J+MpVwrNQC6MwROcN3BZw4N26dru4q5nKa2xKL4sth8TzRF1CiTat43L7T5pA7
URuxrd/xcDU595L4uU0xaKi8Of7x4/lQgqqb3HKFFtQyjx4IQLouOQczEg+T67i9
coxfI+Kd1WU/xL85kswz+v/jRd/1HrYaI+xMx5sUrBCy/YdFpV0dPop9x/Jr6Caq
+lswa74hPWTc/bHv+EjUVbZkgJ3BWVeUZPzEmqZFW7WquojAfsUjbX2olDWwq220
oxWqRRArUB9hlre26h66vnZGuTeTvypVr9LUkAbiSkvd6UDQW0iXz3I3puBiXmib
HAq9wGkkVfgkp+QaxLwJ+tuGJaXI+IRLAWTx5virZx3uD/bhQSVwE/CyCHotNHcN
ieFx7iV9wp4xjGSK3e9bXIAgUB41TfyWkGurNuJyXlAXK0w7cHrdi1uoCKiScubs
IpmxCzzDv0PmpITJGVH/WC0CUPnc6B/yirQsjjiqVUJznjfAUmvrAHe6NOpjIjkK
+6XfwBnxNbrydaE/Fb9v7ghiIx9cK6uMuJ767d1jXP8ZivaC8so3r7N5T9mBV/Vb
ZA1xZ3W4pN35GR0wmnFtbOplUnJZ7gOYS71Yxa9gZtCP/SnrC7CSYvqOVf6lmEnl
cOb2yDSJO2CBN0vED4rJkDfgGg/9gfycACAZu1dJWEFuSe8MdYMb2fJmSENmIT7V
AKnkjnAfUlkH1IeHWqGk0Dsd8uecDPewLPxAMmO7aEngvyDGwNaI58Fn9NwRujYo
oddlMlvz90MZsqZDt7vIzo9B7UE1X1hxXjjNMqQrQbwd/sKvrmxnkuWuvCqJN1hl
ggIAugbc1iChbSnsSwwYPgg5nmzesATFcjPmSxO1ncq53zz7IDIoJaZzIaicW0pI
iG9KJoPPXEN7QWJIxT/otB026nWbjO1L1oQ0z6kzbCN2ECk7d5EcxmHmrwI6F+zz
poZGuKrvCxH6ciCM6elO6zBbzSiXENMlGOSw9/ylvaYpAERDl1A2llOJCnEpfeAX
uR4Xl5YuX/iiadudDxlN3X/i2rc85GQr4TOlH3i+FNQFbZMPv9ZVIgDcIwt70PSt
IZigfkWymFb69Ts86b/2la5TM9pfZwGHcmkwP5TpGdan/9CHDRrU35+WtsCk83sy
aGE6mskF5nvzw5GgbVqPOe/pPKhU42D+jZCfEkXTqV8C9nnGnrT7n1KXZeSwr7Hw
n88EwebFg4KzCpEpFS8QBapp4XctJ8Ck+M5Qeu7H86nbIfgCt6NVVm/h+PQN6Wfp
fBeu8PnKT6n38ONqefATXdfGLxYFhRIJRjTATCT9oOG8M3JoZP8o7m3n+Fhvo2lf
EXHRqXhlGPrFvwoTpKsjtVmudXfA59yGOxMrBXxBLjSXpcY272JGeo1pJSLlhFN1
L/jNg31i2q4GAtylvuLOG5wETiPQO7iOsyiifUG4Gd7ltBhQiNYtd2BxymJzsyOJ
o4wT2nlUcCNlD9ZFxzFGL6LtniSY2tX1WeYgHqLFc3Vjza+i4cm8fd2+63LP5twj
4LOuR656ID3ep2e8g38CDGy+0fYumlAjkP1l/nRAjl4jX7zfdRMRDFPqUnytsLD+
NJLaGozseXWdyhYQApLYyUAPOlPF/pY54e37C+IygAEk2zqHEpv0bJ31n/w99Tuf
xaNJSTWGReESX1VCDh9JjtrLfH1f+Ek4adPrnWBiAzP9d3Opb2iValqWLrmWGA8t
bOB0Wjm4VrD89Rwari8l7hUdeufm2BJgDFg+UV8qa1omElFs9EMdRylDK7Sr119R
4wqnZ9vCkFqJ33Eguf4iW0i2J+fK6D1XqF5IPnFmbIX6efYZlx4mwR/iXwTTtZvm
AXPTo2AvkgMfV56OmD7+Faqpidgy3SchlDJEEf4SciCE3EPXPfnpt4V5e9orVcgf
eaYlCFSK26f8yDG/x9yEEW3GgAQrcOI+zykhrmJLSSaS9Vq3JhtQ0N9W9+ZeV50o
cfH/r+i62LafmnrULDqVUrPAiD8bcA46kVo9MoohQG5wBhGXqkW/9/k3ZeVyQ4OH
PFGYr1+L5+y3mh3BuCj9DyswzHJsjJxQojh4ChYXqe9S4t2QF8pKvyXV4FQjFRfE
LUxcDudF/MjWiJLx5x/wOhW7spvJHS8Y5Ys0EOSKKSbbVbv+aBthS+y1SLz7O73n
o1fPJHFKD8/tlivt6J7Nxea4Fgio3kK9PYFuvSHHS5Jj/wUGV3zJ0OiWtH0dk/UM
oc8tbuHKbBTRPFTcwqXQvYUwjKwOXMLZKz+VZLHLXaXr+HCO09VMemYcMSwuVeJT
PnBT7q9HpfhscDKXCgFNaKTOZB9bsSBS/jwXE+ny2mSaEl5G64w+MjUjl9baaqX1
7bAZ6GInuIRWAfve7MvKMVNxJ8CVZD7AsWAMvMa7aQChhZXE2aI3UKs0dBPC6tgD
bQ7KOi98Bpw7BuN/A2Lcvg3MTo15cy6bE47zgwBu9ucOFVrGfDNVtn04wJcXeHXr
+k+K5FpFqldUBKWaZk5LUy2QMONMk/QfpqEHAHziz7M4d7aWU4mt3cWE2wARxZnf
BMDla38YbdjzDOzkLZ4oKnl6s7wULbjVD7wSXal+Y1VYqWlZRqC2GU2fvLPflpDd
75G10t/H8rMJMSoXrdbhxk7GJjIh+XTJI31YpfidAU+uhM3fc+1OExlhu0D8qI7I
MIR17KmKlUxYuS0QbjDBwiWNOJpXgU7h9QW4sSnUUjhuDwGWgab8povbzWnYpyqF
khhgrbhEXx6hX3RAXHswM/YP1wD1NaS+SyMs/vCaRyNBAJpeBDjQQZfpmjfYa1Pv
M4CzW5mfwb6Ms3ceNRO/sfqU+vsPQG/VTwyaD6HnHWK+Z9MjrJDAv/rqwtwofaqx
wLTbJfU3jgadczrho7O3qf2bHcCM81e7uK011AF5DSTn/0I81lzxtlK/SBU4eymz
3sQ7FmHRcqy3KFoMt2drMRpuVpX/+2rC3m9FxTrUKolBQugsTzwBuexbbTyIzNTR
VlqkFPnGWNYtR9tFGkZwvzpdhWrJHv5jsGgpahP58SEdcF42TAZWgiDuyrJyvBen
/RvfcDeRULbuBOxlsnRM8uN4TWYMxzxUEDnKvYQWq/vcvVfwBENqaJke2QTvvjOF
Qyqy4Bb+D3DHihgqErv5cthRyquzhSBDnP3I+7s6RdivElrPdH98qm9WAs2P52jQ
0NhXxrVPZwIiSaoBNR5BeGo9j6BGAUfPSKMS0gWO74I5AJleUw2ye3y6EVMsTkmf
/fpt5Oj6k8/rk1w6Mi1pDCN29rhgroEgof+V/C42ADfmqSybnAqVgGWpjBbpbwBx
nhM9y3/F1y12VECyBLWKDgF1O65hbZ3IkBFRqyek8g+YrTYqPN2AO+j2hNld3gWv
Vvj0pwwdDvgLzBmduL227KLegy4EOmr5cDYraaCHRaUc/5N71B2CWXYnKw5gyrrE
LGrmNW5dnKHV+FSNXqIoNR/82TCJW2m2GL2C7LIAPuQn+NTvombbMODnzRMvpbK5
yuRhA5A/L+gidX5+HUIUUP3foA+c6gMJgySy2YByKvE16M/eFpmPpfiGmCCVQxSJ
ziT1xzde7ubaCGET43ebpraCFL51BcWs0l0hbdZQasu19LVYUGoVp7wGmFm+7o0K
7DzOkIPNZcTNwzWGgqXeca/sN5M0j7hC7vmFvKX7AsftQnMZGr7B8tWRUgVPTIZi
05lNuCTYzwPHKRMxgp7m8SfJSJENJgy3cVX0pDXxB2txzPi/Spp808nvcO0+9h0U
4jXI5EIxO3k8JPFauen3IZskWhivMkMG+EifnBydHH/0AmT3HtIBm1iNQcpaL+5C
4iaJxpec1EpDPnNS4ybUDZaJa7jHPQ0clbJ169DwoLV+iCaeRx6GeqNjV7Kdti70
1QAUGsnXeGVrCjFCPV9PazXXf0Z/wDDJ4JkMuwlndLZGaaEZ1aaq+moCPFLeF3PG
VejiBFMYpSQjGK8c8MIjkr1V76vY4NbtrRxpnEBoJ6QB1R0jEjCqEuujmW89E9ZS
aw0kHUv2fV3i329sydxLLc4gfXvEgcHoqXyfV3tjJuRUx7h5ur/TKizX5X+jnYsV
lPI8fkJq2RFFreoWuLOJLITT1QlJrSWvfLTn2yHJJRBvYDEhPMdQ7Lb2CriopyXS
laCHhaxb92Nvm6RCenwGX+neyzHQEYy9yyAvl38bmdZuhThdOqLEMz6DyD7lrinz
EuYwNsr96FuxaWmboUwhu9vu+2yIE6rO2ADzkYemr8j6HiUeKu4GwKUYLu6frqLo
Zgb4iavqf/JIJLPKLv5LtsV3qa+/7FuV0AIMg65TrYgCM7udgcnLILVZUU+Am7aP
3q0Ym8VpoFeKqssN+V4dIotFgMfr3MsmdtDFr6sEg0r4vDBRKSK+yCG6dcpmeEb2
hY/iOrNhKAig5E3Kvhr6ioWrUYnkRwGBuGM2ojX1h3ZEm15BkevckUECAX6Ln7Ef
4gU7IbBmAY9AOJS/+pXs8dmQK0LcTdSnKfcMTp2YJY1g3Do9ktzoOMELI/nOLQtU
9IrlxITIwQGjCZMCFUykqgfiVK1GQVbXrFd5CXGkx7yWyk3NIt6agKYPJAzN/a+U
huu5EpcEQrGiCJXI+1ABDhnp1z/e30tumT0aIlZJXbgcLCpZ4f3o26dg6LghjFxJ
l/BjnWxguYtN6H9tAftKkdOjEJTeiD0PCI5IP6RGoVPZ8/8VitWM/65176EnJ3mW
k6J+Ps7oBJFPcFXjadoZtGBZbGhOlGPSnmDbafv4qbWUvaPvIluaur6JUPY6i5Ib
OiLI/EVkJSC4c/3vnREMU+NpF/Nsfn2KXYK+aFxZkwJX01+bYVBewzWvRi+5bpik
6bR+4J+Wjwjthk8NBRVycOJl9ql3MPQb3ITTje1cvYwleU9QPJBbsr9T4uYfVAQt
aqdlSdI0gXGLQiWX4swQkn6274LMyxKlPvSDjcnNalE=
//pragma protect end_data_block
//pragma protect digest_block
8rmWfpBmo4Dj/4eRrIFDswXN1K8=
//pragma protect end_digest_block
//pragma protect end_protected
