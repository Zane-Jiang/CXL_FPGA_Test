`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
eDFGOG4xFzv5oWwYaHaoe8OrNeet0HYkYnWK9IFcxkvxXSPpg2e/1vwgiw1Vrra3
R3RlLrZvpqqF16j/t0s1jFNF6vsij//9EhJnXTdhL34TZ1LtTESUc6YJa5VXCo1t
iuZmDQ6b/IkylpoEPV7A5JMTAYC1n9VXZqYO6HBo8fU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 91168), data_block
MRPnOhEHLZMKxLaOBviNVvi5vBXuwqOdu8o3x43cTcEPs65lNRCSjrJGKE85Uei6
6ACAUGt3u+lsaOaHA5OF+dhkFzdWPzsede3bfGlrvAm2fDBW7NLH+MZB8IxKXxVH
vZJ/h0rrdlg90OT/ArejC+bzLuLQXzgi8gcfq+NIDPGyjqip5b8VGBf9w+0oQs8c
0PM9DB7D5SPfX1/lZGUAOA+iBX7D8CiUBU5iezMPN6nZAW7oSpMBk9P8XZnSVm1y
mH5FXdvYCYbiUVdoK35dWd3WrwNQmJt0ldmhWDojx6XmFFSrdmHtUaVP/y3x8vpX
zlBqLNr8pSIEFZHeYxFdlCOB7eoDThNB/AoV9wmyZog4ETHi55woAgASJmeXOCQb
l95QqnMgM2gL/QRVo8uSSjpePBWf6uj28hRojmP8tfgaHhn/zvZvPM9P2s9QqDrA
cFN/HBSPpMDbaXVo80HYaQ81cm/bsNl03qMwQ1LA08gyq07wGHLupZYEA41IgOAN
TiepPBz8klw9pObjbfMarTGYkeRZzO2SIJ978XD0rjhAX5j3Z3nYhlzH2CgOKlCT
LnvZQ6Ka8oVOpXeJnPY2zBerKQE/TRlxYilh71ZN5uVDlPZC2x0UD7Ee8P8Ey5qw
WmapcKndUb59meOFmCJUNp3wv7W731/EFJ9o8an9I60vCRgl8HfJTYcVjte+K5KD
YX2fOhfPkgYjjipiCZaVqeRkgTlxo8BVh8Ckk5WNEYs7ca3kEG097HQBgK2OtBwC
NBaJt3NjY27zLh+L3mu3MwUT9t4iYaIMztb9WYpwYXLUe0E5oxAka1loEdHWOiLa
b2pIbBjwTaVIbEikodZOoA21oAa4UoV2U3jh2fQqxY0ekvZxKYGFy5YIUAxmBw5b
zLPcmRAvklh6AEXVqRmbO3sAkCAXL6q1tLpag8wpNzGEqRB8fCU9qcHRm7QS6Wvd
+gKO6Rvyds8GU1AoIpzK2/qHETPLEt0Nq8eAJTrW7kUlJlINUyQHfCtvbuOE9lq8
kyZ4Yi4ES0aIa9ViSVIhENQtqayGnS3PjBQc5ti7NK4ddaOyj1ZV4sUAkyXuTPx4
4ET+6gWnSEvnjMu6BdS8c1OX6vLVn4EHMaIiQj6b0kiVVra53nsyez2II6ZsPept
Q9MqMZU9P3Jo2X5qHdeH1nrUH+ajMYHsk3gmmpjzeec2g9i+atCDRH2/3om7hkFy
AFL3VG5mdrhKDX5aQpIONkX4dJ1XgP+5ia8KMTGxuxkedVbkToTKQDrcYjov8auG
JPwEMCLeIKnLv9VMY2An9S9hkcefPv2RaX2NUzvKgcdLgOTC30m55/W4GL7Z29hX
AeRkQzt33fQaMgm9n3OsO5NgZIrz3fqj4A6kPLQUdXoD0EYGKiJ1+HgI9O0ORbhE
xwPErc+brqgLpTFAsumJvPBZcx4/Be+bYx/Iv7sX9rowXewqIhyftr4OXMgy1mTp
QcHp6CzcJ9TntEf7T9uCB6vrhu7U3e4t3ZxOyw0YtTZzCmqP6kbeTora7sLP9fBs
sOdDbH6os9PslGSWEiUPwoakhM2ScSdRxixKc6YdxiRduK8nUt5S8JPujrQydSCI
tApXcnadiQNQ6YlZzZAjEaTSZwQC6Klg5ZEgyY4eQCDv4LN1MJmri22iVtpYj7CT
4Av5bUFKcj3o3/LB2jzGjYu5V/tfklY3Rquti/Re5Kk4Rv+RPLQhGiwL+owTxaPv
nfooJusahviegSy6LWRFzQQnGyfpAOyT0fpUW0Q1eGCN+4KRi97QAslDE5D4PxJs
G+1fMlNpmrqXI62juFD6oFQjHjQnpfmYkiXRwWwOGFJMdtN/AbTXejFix+5X69Eg
5DK/QK2QdGFrj2SF6BWEI/JAWBbADQUCRYMeRnsq7qLCDoiOfj4XuB+qR26zG7nY
pXcqzRFLkN0FvYtD+GFwdKpgANYnraA9A7iK/AuxMjRFLLRwb+eKU+xsYthdRtzZ
0a3BKQqH8ej7kw1IK8TneMycQ5RQCVbZHOasMszylHeTurKkcvHfPHEJ52bEeR4m
slqS+KJV6HfFTYeXSqKFtACTqnVPkj3LRakZWyn+44l6vZv0FuSbCfBL+TPGr+BY
cxOX8qae1zyBntQjPRwEFSjeHzIvar93iLTxIEtyBv9Ic+LHHxUhamxKTVf4UOVX
UxFbfEXbY5LmHkngPtLOJ/iszRW7ZI0TXbpISLovCKHLzv4/oeaYsLMfM/vmHEuf
LJnHz7NOApSgpwciMlTB9KNZ9dL8wzisr2wIFh86U4KGtGhwqAKeF0SfHmJmyu/3
bGdg4XqWSUo9sc5HIltiRD+1gmrpW9Vfghk9rjPmMrjNZ30FJoxGTemeMOnpCcqs
MXRKlUeIjZpfOIrq+73pSiHSs1VpVQ1jE9dq5j29rwZQFNU+j+c2iuaA+j2fB3x2
7O4qhgB128dA5hisWjpQGgXcBs+0G13Qc8dXh08sIdQZZJ71UaUIMCP9DtpFhLvi
ofqoa+y0/4FIHkxE/3yyEUE3YEM/oH3UEdPA8JO9x9ucq1T26yH7TOzyw3lqPMBS
RD197t3gj2X9LQMEMCUsF2RLhoM5sjPGZjbV/SeVyYFryPBVwpOvYaIJTOBcngnk
dKnaUJuLmLrqwOAQgFGWkE48Vx6ytDmkvXmsvxv1CVWjp2JeLDeGEWUjVSaZv6zY
03QbygpPpql282Batg3nxAErOuAu9SOdSRBIfLJMKKRE0exBDD/v8NipO3Ek6hwz
g1dKZ4Fl7ikRtvxLvX9SVIptPSJ4hQkSDrc56xMSI/FBN+6e0X9LYpIHv8O3tSI3
VZ6r2AOY2aW5+0/vxm0qG5rdTcuDmuISXdmLbwxIHC+pbWAZFSTMnEoy9/t6I2Pq
upbsxRtR+kxsna7EsCrX3/tBaCmCM8Vg31CZsCcD7cuOj1lPcVjm/zBJyavY6Wh5
Rq6ZjTR+Tg9fW0W2wurWRCjeDTdgatzJ+Xs8vV/ivn4fu9ASFuKSyA934kLCEwDM
d4heWTtKkVyH6FNiZQzhg04qrIjk8xu/rlSokrhTJnLn8Ztpi68q6HujWbEtk5v/
V6Tt082GJaLhyBNFFto+aleWUVJwcxWhs2eP32pwGOa6AoIPpOeJY7JIrh+Qph5h
bRtvEqa9PTMLw2w6qC/SaQNVbfteoNWjk69wrCTa0jxuhwl2faMYebIbvqMlaXCg
PpR38uh71DY+jIw1MXt6nGE13CKohX1I1L4IN3C0tUpV4spIplg/ASMRuO1bKlKy
3qgZB2SUyEiDP4xsJ0GlriXYm/jQGryRspEPEfmYzoL6Bllng/kmWSHApC54tC6r
D09/d3ZzfhmmUIJOKaj+N+Tl5GSkdvKYXa/UsLYlPlcScor2DpcX9xOa+bEIhhbo
F9PDHO8hzrbETfJD871/LSrQWBHE5Ulg55ksGQ0e5iwDWckiNPXDuEHSyn1i7yBq
lVD6v58U52rHGTClsYckq0SnpLZaxXPFHfObDO6GnjvE44aZvLfSyEuTosPwoTzW
HhWpUy0bYX3yQkRcnQxtrpfj2YzhuMvMTrv08ayDi+JskFoqfUaHH7/ojwGqRki6
J6sz8ocluDu86h/77fw+3U53NM2C5EiyfMd1cv2mDEId/VEWpEYy8kBTN+zzWBQI
pypvCQYqeVcLAgkuYne/VmlLBiidYX3E5GUodhvlavuadlTPd49ZyObchNjzdXJ/
6OclGMG3jfKAcgcFsJvehyLVVirrMqds4w12CAl6+OxzvuHT6L0xEnHFGzOOaShr
zvjok1MWQv1JAJLG+P0FBwWCQW2CNi8tNSLhGmnjruap99MeLPXko19SKGmD+pb4
CAeHAom7Pe9IvfmCU0DqFNUHjocK8uRv4gZpjmWAklg1HxMLC1Q+ol2HW6jfCDqH
LWEULAYtFcXDevGbYrXfqpq5wkToaSWgCgzBFt9CH7H7Jh1mVQpZDz3jy3sqV59q
J/QHTVeOcgnZ4s3YSgTMbg6kToPecxDdCUtqbqexCxlMMbBou0SIyC2COomNJcSM
CqEnvPMlywlu95pPXbMPNn3Ij+R3LIfKnEgfvAVb8cwkfyAFfUM8TTaL7Q7pdcUJ
ltWGh5xdpsEFUvjoxGtn/G98YrNxmEA2VH9hwYpbkf5iZBn2jEJDGgqed2T7BEH3
ap3CB3KuZVDbRq7WTFAIPlvxGzChqMF+oejICovhuDv5oQ4+vnRR1YYTA37ZX5hZ
fQL2I0Y739HfoupkNZrc+K9mmXQyqzoaCtt+NrmM1FtnRsAQgirVMiK7rOeOOqei
VyWkgRwDUL3zWrMnkmhw1HmqARov//5C8fe3JSD+7RArY9/KEXC69fk0jG1AKQjW
/RYOixfh0qcVTkOrC0Fvhx5W1uAM0SIgZqvDMe5g5kxDhczjryOkjT6X7OI7MvDc
rU5rWyimjNp2rfehc0KRihn31oWdyLcfoIjk1HEANrJ9rxxx4GalDFtisCgy+RV2
keB+8RDGTdtkrUblLRxKRWAYIECrUKIguE9O4Und+8A2FUBU8OC2xne+csMDzKIi
p30wlinshKBAW0+lMQz7cbcMj2awHLi2SfD8rBH++jP8b48FscdWPzsoW/ueFw+Y
NTlQa/N+S1dSdR/uj2ltRLF6+zUeck561ZCyJuxWohRFeMxV43nF8lsPNOoWMpRk
eHHHJVtntoBN3HN5KKeUEerWunjnCE5VJyxauOnWUJrOr4aS47J/DgEUL76DIlLd
peZJE88Y7otRaB/EK/+a3f3sRLpKftIFFqF13STguWMsI6BLUZWuk+vINeIRFQZC
2yNYuM8m6QYVSIu5Ref8z2hOfTiOqP4prBsEFJhcJAZe1YTMVQo80ei1XAqYGyax
wobELqOGM9XaoWmFmfs9jmtDCwCm4WxHu+COLtaWrwm/GGj3PD4ezRlMKMvnd62d
3Hgy4xj8llzIsSm6KoC8O7x0QuZJoSE53QdB1wI1zbZ/5tYOtFLsapCAjNON770r
enJbqvwRLwjU+u2zNHa+siJGxDu+++BbXZHtQ6Y+VrDLK3mi9nq5jWtxQG+TA4ac
A9Yjt2/winTYig+ddiT+L+RYocR9ckb4rrANDn4ooQZ9tBN3hewG+l0EFBFvyDEH
lf2DHnoaVV4En4JR2lHflHjRrqeBj3sakg8HKYFGYQjF0w/4/1+utIeRKoBMIjLO
gIq4zNppWwxjD/YPFWdn7xBDVb5JH7PIxRiCuZvb+aHh0if0MvKlKzD6VB/llg1h
mZJdwMb300Saf9vEPobNIgSEF2iOJD7hgXCBZb/GmkZ/LEQZeTQVpd4AeQZKlwcr
lM0cbY6k+fAze/JdP6+k+Wp3Dy9efx2Espyjk/NhCV9mI2JrhWFFZj2jmtsJqkiw
87TRKgkokI3KNPRfNHAjNogP+Z1ypQygRg3m0R9jEi/RoYQHVzriGjOooEYSgWYD
M5CCJ/7dqp7oZsVaqq7BxBFHzhat5weN9oNjWjpwSwhwCuUpPzQ4KIfa9lFliq3x
sLdhflaNCUv4z1urV5pfIv08KZiD7PtlTewSqkyY5TJ4sdpMePsht31VHG5Pth1w
fkxe3HwVIZmgi1fWobTnDTVEcuALpojXj5amB1IktpgySUSQStIpQqvWguskMXH/
kz6pUczNv8y6B4CZqUg61HxAjTUaTq6XjnpwVs5fwLbwK5KYKjZwRhNy19aUsZ6f
kto+VB37nAiL4Fn6c04ZCVLJIK0K6yJ6X5+ijIJKumb1mHXKezIndqTHz2OTOle2
+4qkD7Vn+uQg57V+vE5mmyCjLb1vT9v+FtaetJoPNQdA6M4eqI9TrHyIh3qsUUhA
TtxhTQHB24KWE69Tj8wTvR2StPGW4Qt6o/+FzO+0WFpY21I2mzA5IHNpU6zMHrTW
v6umuAIGDqGuWcqznhOFBqgCRMKxexNDIw0IsebUwVed1DCILjTWlgVraSol7NIP
f5eTHO0d5ZkK3lmU35fd++u7+lxo2Hfa9w5N++YsgMc1g0IzBVZqhlHKkxkawT1e
0FephHTr6LKb3JJJDvJKlDb2YH3kriWtGHOZSro3y4ty1QBbN5rhUw6E1JokXN37
uSMA02ggNx/ild/dt3YQOUFQW2Osf4VatT7NUDVTD7MPfJ6FNfjt9Ewp0vryeaGU
pm5+VA0Ra6/hNXp6kdVLB89UakXt6Mx2w/y7QviA55owo66+vxCk6p4hIm2HBLJE
BUolamQ90IOFTCald4Mw667NHQ59KKzrBChiJPbs0nVk0uN1xCDZCy3CWz40Ru69
Zf74bolDtdkVYPpNN1Rrb5qOdim3rr/4fzDcIRDvG1EmxedRSC/4wXaCPkJ3Kgnd
5UkwBiZ1qC+yTMVAWjgkITr9lQPRny6uM2bpJoBG/E1WAP8U0S9BF0Hnkm60NN09
cu7V/MgzqcI1dDhWgJiEsAj4+aimOHIR5+8pxQfaUVI2SX1Tc4+0CyAr3jTxgvpe
ePLDOFXAd8o64BWfmcJ0PEVRvo+MXBm/T25m+5B3+zXpOp1aAh9ZbzCZ0+WtqaXM
3sCo/JdN8ootKAXj41vKnrwYesMfJVdanvBMRpMKJMV1WpnbA5S7qW+uq+4j7lKA
/MpgCMoQv53uedlq/OKg014+RZVtOfj56O0jQhw/25NY/gsTBW60naqfF1/70Z5B
Pd+YXZ8J5B1UAKZn/4E2SOCCmLXOrB7oP6iF7htZ/fGAVcfNVOEXTH4YeUpVhBTH
QXQyunrVfzTBVbUl3I6QE0GQQ8KMiz49kAO5r6gNERQyki/ctct037rM9wZzSOmp
Xb77q5DfR/6lvfzFt2N6pCI96NiPNrA0/lvUDdu50l55/N8mUrnlZY4Gpa69/IZE
1H9d4SVBST5rsKkCWiKirBafkadCQIZhCXap+m89ydDMfX9U+3UtE2JKgwSI2PwI
wjBRKtMZ2P1CoSANuHnd3pnbU0H8vWFJI4MO2sVlnsdAhK5FjJWQ9Y1KJ5bGB9TH
txzc+40yW0Di8xhsVD3UZXk96joVjgX7JGxd+hgeCaCOrSFjLOt5mJDN8EkK8OZJ
EOb6imJgPhUX1yrfgo2C6LbRlwcl9uLMdiTerqpPKpmV7Bmz1TbdZHrU+6/DOzHZ
Zjp8DiIHTq6IHPuge1PXov6qE3veZQgbbxLTgFss8BUKjtK/AVxPWgxLd/7+tLjY
VWpRyEAHjG1HKO13/Ie/1X+X2IZJhOOZG4tC0VX93VEU72xgx1wyuHppTgiAc3T+
LkKPjioWkBAb9RgNTaJ/0TSb0A3PXtYxExBh14jVxS9CUanAgxD2F9RD/l7IkIqq
r/fcZHfXMV6hZLTjvqUFtwYHY0/m78pCj0U1uX+pCpGZ0njHgSuqHYihSC3iZ35P
JgGOPBEoZir32oPqzOUF+krkRgmrO6b+t2ENUbjEtHl53yKdHGKjPHabqPn7EzgY
UWVWlWeKacrzMd0X7Tg7i+QTDg3dT6TFMgerFVQRso26my0g632Iva3SHUP9P5ae
aCTEH7Ga+TYmbJ3J6MRkHxjRJuaeVIf3j/Q+2Dppy0gK6uNt63MbwljjVjGYmwiJ
0VDIVgpZqcZWVU1lk/mbjurNTG/XEVu3TQb/TS9YRTw8Dzpp23s3QDVZ9yyxP5aW
jRjFF6laQoRAU+NoaYujsqjPlmbbRTgLSSvKLa5XIjHgyaLoG9BRnTtBNR+bVDjq
FQNSgEAwDOj6+xXTd0hcphujJ53qflkjIj41FtX0SEzuxs3O41pfLlLjgaSC0Fkz
JGcOlaSUTXe/qfJAqXZRTdCQttVf7enbMl1chag9Ie+S3Pv9kPGBahH5cpRHGIWy
7CfahT+fne/g4KuoatGU2fymBI+perFYWe6HY8Jdl1r6rQvvOfmIHksVZ7C0B1oW
kdjBQGZG+QSjqbstJG4hnkxQGYYtxy8dbf65kDjZg20Txvd7XCBhTdG6xzRTJyKU
yLLaSGvgHalVJ7tDBSjxNDRcFOv3rTSvvNDmlcXTpzR/PxwBdQ9XLJCQYSM7bmVW
liwSmc/GQNZvhAsEJU+AY7rnkxRp5zsgGxr4X6pZPtDym4od5kaeJ0EQCa1hGUqj
8e2cp/W/F/Pz0dXwfBCaB6YzCQgc3ls4USpujw3QhzYXpklfJIUnjPs2D0qglSl9
ZmEHV7vR5FJsYi9m8US3Vy+c9+YJuR5RUvRJHeyFi2n4OOsTtJEzAUa0B6WN4qSX
QfR+6urC4KOH6s/qxpJ8XmtfJD7wLZUusIgqtUKKyYaNrWi3J1LzlJDmy+5WRfyB
Iyhhuj8qCS1wGSw8ko2xtqde0SPHMbcsf7+G11G8g/TS8lHKwNYeNJYGpLpc5raa
3tDBTmfK/EI7hxIXDOo/hruvvIP0y2p1r8xTOvl6DyPlzzJUDQzupHzWZfgsmp2P
X9Qz3rV16OvFCOb0FX4I9Y8hgrOyxpZwYJGMFHpeldzCKtqKZEIN6EUDzp3jZUt5
vSgwwM1qywUVHfL2BM+kS/mblUAEoImVmhSt476YlfoxIhDse5Zrf38/hT8erB3N
a6H/JI70xI2Z+02j1/Mp09xe8u5S119o95oiOJIogTj3da/CmbZW0BunfcAa26SF
9l/ZwN46zmUdVy6qPWlWBIkm1CjASopziZvpNoJqB2OAHJv+XxO6Qws893mtFwZN
nCsNmeOUTn3ta9MDuSkwHaNeEecahylzFT3AkwvoVbzd26Ql4dQElQx1zQzDbK7T
nKLbATrPpL9sOF1gtT82tWmOJYsXh/kAXEKmaicgzX0sgVrZE5PtvK7GmfsX1hXh
FuU3sldwKyCtbJJvPBiwO5cVO/pZ0Vt6NZyHbVzoSsBTme4rQPsTyEnTFX3odNJh
xnP1glU/+rqX0Qe4tMPZuEea4C+82MR16lfU128i7JNc3Yc195/wwOBo2IeYilSH
gy7WOmMiduKBobjqfgHGSVoOybIH5P5UrJ/dGtACWKfPr8fLLqEAyE6t9ysYE2p5
rl9bw+yL+Vz1OQl5Fj6fyxInXNM94o4uywaWLPjumEVrmKmepOH6j1r51VdkU4q1
lUDiDhk5ir+gqJA3Sq8cSZoY52Q2JOosi6xJmbOkC/vNhsnS83+ywZ0L2hrsXV1D
9Ofk8NjfBFfUG4tU5J3hqJktxz5xLHoQxz5fwD8L4BvHeZhdB8xsn9PGX0CGFJyq
ducNHoFBrYnbBgSSKUdLyWKv1DerpmU2i4CQEt0xi+0PP1i81omjKzDILjZn3GeP
BEPQjVJgb7Qll9hnHwKvaPQuntaSc5U79u4NXbwSLVkO+HU7X8nNRgHWs9V3fNNe
7PtGfrt+i39jDVX2qi+atOxdBaZZJrJLGLQ6HcaBshFFYK0c4JwgDCsR+0cHTEu1
OUYyAOSoT20OSsukUBZgr9mB+9QTlL7+sxwEnr7ITpCV3mP4KhhBcNchWuVZYFbc
V6GMWcqwidP3z4iHIKFmJYLyvSPMXJJqujFQyZbvpW2vovpTl9LViL7Dd+JqgBlI
R1sVvDkOre2rt5ljp6WOKAEru67Fuen15VDGyPljg3uZQxh8qN1Rx6UeilogggSV
Gs68DciPCat1JeIOGWXNeC+Z+0Dp+PGVjAUoijAYp7nip9xSi6tkyQ5SMCWYq6j4
7Y6hR83Ojrx19UAVRAcsivBlhIKUT3fju+DN7oUpsQsvVnRxJ3INyTEqzPjH8Qqe
cVuAzVd1amEhfo2BY8SbJ8EF6eRkm150pXAUWSMMEeFOMbtxdT61Dsb9X75vIdwO
1hcaUyGWPaFqe70XLKjYEhkd6O9Ipm3XmSprh9Y2sIPDdo3FWKTBk7jG7f3kNL6+
oF0QGx4xESGSC4Kz/d3E30CZv+HbxL4e9SL9xgoppuuLjCL70uOVWZJm1jPCXHa1
G5Xaxq5rVE5kVLT8ccRwiaLGm5J2MkZ3rK3DT9DaLES8Cd/utZ3o9JpaKlEHAMFW
0EypHamJmk1lEjbDK196yq2ZNUcN686+2qo38LzaF6F18nGKwhYfeMG0rf+P3aaU
GLAsvqrNnxLujjzyvz6yjCGjT2tD8m1TughOWtoKJ/tFgtWImCodR1MPYnajQF19
Ex3DRRJQbVA9HpwvGhZGlfy5BTLAlNCHvQfgsh1dRpr7Ttu0k9tl4XCHAta2Ryat
DON5yEJjFYCP6MTw+91MRE2PqKcyXP1vsJUV7Mk/a66RWEK0xcVGnPOT/Ric6QaS
WLagcCWVkXiASCyqSe/Jf84qn8IOK7viVyFxuOZ1Cs9gA8JqMiWgurRueM4Fk9jN
crNSXds9oonAHUD8b8XFCv/BI/akXoGNKLrV1rGeUGH/kMDF0RFjmKGfBStwYkd1
/sBtC1zsJFOWE3qVngde92hbniX2lMuZpbj7HsNuJTlC9oJj9MRCngNbRwJJje6x
180hrDKC1sY3qT+v5MrsfcK3XTFGMwi2hnOvwV+6Gswd4z7ba5xtVaKPMsHuRl/G
4tFJKxGGXwmpzalFlsd6OO9WI6IrlM7qPY0PRMsyILedXEH3sMt5UqFw4xNm94Q/
otv76h0KeIiLNUkldYjBLngP1bBIxPYl2bHRZUY3zimw+oN/iEIwzHvG1RLATcJW
Vl98OBHNUo2B5VIiU/URl3nWaoCdLF0lfgkUPNvHs9fdXrX4yeBRBW5aSX0/wDqz
DvJ3p6ggvK7wyks0UvqRYLaYKLJrWnHXcIJE47ri/ZqT8kQF+S+VGxx+ajG7BZ5P
bxSy3EGT6b+XPqbVwy1fppqTJ8hj9qg6z1oCyWvYKdt2+R9QJbP0mMJKSUgow2p/
uij1GxSC683xKuMMV0ts2RB3xWT98aVs8NsCshz4r8AdDNz4QCuE6x4D11EB8P8p
jc8TNrWfjZ5ldHg4Uh3lDSs3CpH8A/6i8wV7vEKwZDzE5bOl+uSN7p+L5Z/E1TWa
hOXE84wFT9la4xBZCow+upmTFIs5hfoXaMLAMj5ArrolEIxKccu2/GyHEIM7VPVt
vKaDtLrUYR07BVshBJGZ0fcOz8jZ+yWWRNnNBB+okGYXW38ADCQbCHAupGSbm9iB
SA8YMHsMkoPszba/dcummrpRyNgfQzKUGIUN7fPUI/FEbFDmTBuO8vnOgyltbgo2
nE11rwEbyS+m+yrxqpOA9PXCvcUmMXYhCfqh4jiuh1PD1t48Bm5kj60YDnvq51lV
9QTUAnCtqWIN6i1SdF92lpOmScDy1SNBf4x9zk+IAAHw3NfrKsKE7NIyN2J2XPS9
aisTRuDjzqQbryFl9KMFjSUPRWka7rScPyHWB5X4jh5UzeHjzphJqDuGUqzvzIGG
5ZD4kA0vCzoll06Qxqg7z3sBT9OaBowi/mQl+HaCNby2TQhhRrGWpg65aLGRkjwi
7vE9ZKtQHqgLE0aGNy/u4l4EwWEnxC1a6oQMTmO8hH4IONNms4+rsKSUnDCLHy2n
um7YFZD8DM2b6nwtarPrV4e+AQ2vM821CTm8NcKGdBnUUIfeCvqA7mcxsP40KTXA
Jai2Gh7uzw80osIYuNcYx2eo+lo/a3f8O5WtvGycbrl9AhIbdf0vf9tvjelz9zrE
fBrI8Mb6nqgSIiLb+wRvwJgjdSmZXRWWcPCeQ2+j4rqByyowx9dTm9qRdReV22v+
N4zfvYVgILAMX100w+JR3fy4in7N+/94gmbegEOtRBO86lkNrYF5aZhLjxgl/hrA
0cr+OjjdBmUFvoIPH/SHRS2i9AAEcCujzqpQJJQN7LOjES026uv1R4fkDJs+I3rX
vKiZ+Fx0LY2kmhhz5JeDyqXfTRJu+r8JM5w1Sy8tygGYx9pgkDSnz2VSRnBI6RJr
HXXV3kibU6Rgbn4TuPuwtFYI6iEOzUTAtTP+Ug7/b/RGQy9Ybo+GWpiZQytDmOsk
qIeOkCE3NPdKw55FcrWk6pM3Dgl9wUH+9nqsRASm41oI2pWoSJgMdq8cOLJujfSB
goaSUsAZQha8zOrutB7R2mwML/wjVtFuTYRC862lUE6DUQkQCd/Ukd31s//H7aib
Zg4MZuKugWa7R0VR1LTCCB9Dfwh1372ksZjczvq2HMZCjl/y67237c4kCH8lJiVa
f+ZVP3NJX5EoQHtxtXGmMRmcG/A8z0KtVQ6LRDMVeaH53x74fDNWAAdAQgXS3TG6
IGJZxKH9c4s6BJL5uFT96QdtHcsXux34MSkwkFWrr+C3uEAbpOOQwByS9lvkwi81
2HbVKbPIbALErhKULHXuFZgybxs2B2jSslOLYhNGMHZSEjlfvekfaARtPJ/OhjE0
HsDAb90t5n/IFeXUiPnvxAGrI2MnTMmHMpXsNhR1BWKmkueaWpjuIHUPeJ70rEh1
H5FAGUkraZj3nf2RsOmItClv2U+duQr3ps47Rgg0DJb+cNQsrJh4yi3a+jHYVrk1
MRpevILu9qY7MhsKKrwr8EeoGsy+O+bSLQdaV7yxtkCgLc4R2lSM+ynMpILKiIyS
sbe21DKzGDcV+ikDYdALljP2IfkkL2HaPp/n4/n13uxvlxdPtWj5OmUR5P9DojOh
Y+GsDZMi2GyWfz1HPH4ARC2a85T3AqFChj8pu9i0nr2nO692bW9KTW8BUXwhLhuP
RCAlNrewm0dMtBTEc6OWcC6uybN/+AHoaOSS+2qszpQplpt2MGtHdixd2ahGsJzI
MRs1bQsSTIl0o8FkUQc8pGdEKCOCvYZAfmexYMoTVMT+qbfcj0M2BUk/K/D5Owy3
0LFLBykEoO60OOD4vyJxTQGlne/v5hcetQJoQN16cYDVvRnGJmXeUvOcXB+9Pws7
O4TLFEfBAJFvvJHJQVLQ8d+NqeaFz4lzJsCVC+irdA0cf0ZfVUXEmNCQ3zAuskiY
tUuVFczVvBfzVFTZevNn9UnSE25sJdj6Grj3VgnJ82E7tVRjc2xCBLkZxE8A2vZk
JjzyxyIESUc599yuafkLOn5HWpQOCYQnX+cATFaOkri5rq5be/65Lucoomy9PBIA
sk5iZfKFtojlCt0PirE2+13K9BwaJbWvHrN4woG9LohVZpPMKPlkpos2mFLWK/so
PaMfep55oC8XsDeaJZm9AewoH04DbvXUPpGCbIrxCRh0/h+EEq2P1hkQ0fd461Nh
Z8HMAz8Ws/GYq4EeziRjSDBRrBL3x7lp66F73fttblJPgGqJKfIgXaK99mlRCkpZ
YeJU7iRryBY4G6jYL/rt+FSaJ5h807Q8A4pR7YyAYA1n+MQLiE+Efs6UrFM3qEJo
s9Kbu4Yqa/kOuTWXI2/HCRcn/vArewaHXpy3/wJriofIwJo0YKkV1f4UvSIfLZdN
qYdZl/FU0kJaaj5U8KUBHzBfX7jcbDdJP6LFY0IWhI5RKiRYUL43Ajzor0g/ci9R
3o1TuNRqjvIgWcerNJpfu2PLuFatylkUjYNaxGYIsF0DT1QTt06UanG5q6gVzHpM
V6p1+/7w3rGr5tcZ98aiBSYNOOaDBW7LIASLiUL7ydaIvkFCBGPUm8ykyJigwkq7
1kIGYW9SR5sBjrPirUyKssVx90TjwIJwwGcECwDEoTjTiNXhRPp/EemEEhHYq6x3
lnehufznT9Pul6WbH0h4HijGpdYHTMEK6sqRoKqv10eZ1ZXC0nilAVvlTdyjONjl
aAdLTfn7AZseDBS+lA74llQ5ZPYHxB7JcvBIzuBCaMPEhPiWPphpAASvvx1LgAHO
LL1rD6s5WLVAI/AKAInUIBuZQJYJUs1Z1eAcPIApmN7k8HtaINqs3BFuSkQNxpIV
6/0VxTtbYNocwe3VlnVFTaEwQDjY6Ug2ZTydEXIPayq/0P0JxwxOSkVdpkryy0ga
7227u1Mc4WxcPYRlNtF7a2cSzF+Sy7ny96S1YlVSwVPJviUqCZH9xgMUkpZmHlt/
pELQws0lJ/cxuDijFOaAyjr6fanMgaZt1Nhwnc1DhmWJsMfGa1v7uF7etuTUWUiS
b+sr6mIMZkQzygsT03OE9xg+2ZnpbYc4Vgw/lvpaZpytiohfadvm20XTT527LAcm
HKSoOj/wH/PNY2p56je4UUmr3++SLVChjXN0CYj/gCVTTotIhfSogyoOJOCWho3b
kseUYE10PquXlfDSDpDc/6gynJaRKxy5NT5KFgYL4/FqjCW6YOnEKOqa9g20OltX
oajQeD+Ut3yUr3FaVGfwG6UUsU+OvKW0BNQbEMG/9mvDUzeFWfl6VsQ0v5LT11fx
iV5bCcAIyvljjC1KV0swphHP7IQPJxuPuNwmGAsQo73nLdiP4andkLbynp29/4Ks
VXprtyoNv8VM87whHYbOfFtTxy2vurAEZj70EDQLeRl1PpzJTiGI0K8cbvCaDAeC
u/pWJ6Zg+MLGurC4DuepUh/W7Cll8VrzC3bPs41oQe+hix5Ibqm43LTi5KA5PmuH
TW8Py7BcBHFJx1ho8OrAa9goTW8zav83nqgiZxyzA/tJvHR41GHNp4szN+HLobzy
D7N+L0SVF4wX5DH9ELyiBD8kymqAI57rnYRMVjBaoFKE+8lsfsw+xu91Mto9rAmW
Gjz1KC3fDynh6GgAKYClU974t39yk6XZN+69T2ryQ5kvSQ2BJT+y2emyDAcl/hN7
MGfKMCuqgFTwlXXk+h8Kd35QjpegTcPiFtUt7NrXSggMv8MaCBWa3VrWiqDUi5US
584A2euJsJmT6a+s6Hg/iGIJQ7EwpfWOH0XTUHgyXCVGoGPGniclFu7mfc5iPWXU
i0+Lyf1g6FiqzzXnVyMEhk9IhNaMwCggafeKb1GII2hCSbjkEM9lyZRpbi+BjeRT
4uxfMQoY8VQdicPopnyU8W0+kWFjcvyeYFAi5mpsmZSEdXvBW2qeqOMnAtUCdCPl
iNAuRaxZ0TJTvLlF9BcLf66Xu/m11PQ8dpcQBAJWWK47yrUiiUZiFcg9feFSGtlx
95/c5kctjx86qrcB/g1qLWraTLpOQCdbrEeu4MddgwyEfuqG4xw/Hk/myCFBaWM/
GLJ/u+dBOnu7N/bLjvSNzfGE3L7W956satb9xHx+5FL7hslEVIvN451RGBltgEMh
7MqcgWfoGeif+cBP6qsDr7ZxehugK/WAO5L01BlmAy/lp0mjMibA/prMrsE3hexf
FOkQWWr+Ds0ZpRx54hT9UuaqOGQKvPPhb2IKgpjsxkOW7LoTJz6dEUyxKG0/02nb
LJL8Bj+ogq0ZrRIAaqQkOwsvmANA7N8jdVY/hIrpkq3ZrlZ7yF1joqq+RcXyWCgl
vQ3y5iXkWXvEZgpZd/gxbeedO5OK1Rhq3fmtP2+6NZjYMtzUJ0KUPKhmmRSMt4rr
ex4SmT/WLqST3Rlt/JShoVVq2HOGYvvbywdukEDIeawKB2v6XqBvBIoTvnOeg8tM
AgoL6nxC3bGwVI2oID1qW7MNk9FBkGjWXJSyeVz5nTk4x0FfihJvormgf2o7r8/B
zz/cyLiK1P78ShXNCl5MRMVdtryFT425ZIzhj7h+sk40nsiDbWFd9tucAl9ZzxX/
416RabICWrv48iL2ycbmYSr7FJjeDFTnz60cEFckkuICUOnDrhPWliDlPUWxiycf
YV4C0/EpfXzuzAU9aS++Hc+O0y2Mud5aQVyunwrpVnKJMtQNC9VDSgiUSds9wRVN
ZhQaUzkaXRDRhTbYjnDYoevSIqKnCq6n4gu3hngqL7efkbjkn2XgjTlW6vYiS19T
JAhhQ08G6yi+G1XE40Mg9DdLAEYIX6aRHvo1yFsOxeOhf4ivmkTeJ1yhCBVv+R9G
b0xh2hDt3Lw5KgGD6psQgd4AfAGOf9qyv8tZavzcvWFAurforlEULzkQoFSKBMGr
CynB3w3PCPfQ+4wZwjshDslN8/Oeetz8uKPi2Crn6SBHVbQG4zxpTSH6Q6Q8T7yc
MtgQqvSs9iy1Z2sHQfNpzpIL4WRIwcn8kDiLxAVLrqAKtq+LfVADTTGNJtDxeJfZ
e3B666+1p9Wyu6X7MDBG+m3dyeep1gvUQMrx7ETzFUN9PJGO6GuGNdIfMyPIFzZH
Z6Xs80xH2ZEDHzu4hMcORXMDJ2AEqOxeirrrIj3+z/fzr+EjbJLdwV282dE/0SnT
QiZhAl2+jlFmaTLa5YzFmCEXNtXAE2/EaEyEETvJwEdxhi3pM6f/bThlPv4zZd2x
Wgzeh8rUl94Mwcrm8OI+6RS6E+xXu1qsAmKrhPCeymsHQHnhCJR8peiTuIbhzqCh
teUUrsKXeBv6Nwz6xDUlPWCX9P/z6ArtxyoKxNigLOkqAi3/geICVv8QUwofZ/3H
QyC70sDfBwTmejsgee5IRhjpCZzbRvIkGtQpeLjgDgagdbFYrXdAVtmi0lBhXEyT
yrN8Fbu1i4s265YEv4lloff5B571IK2KJr2SMzLTzffV+owMCpVpPbYSCfObHcp1
KRUOOJOQI5yMvgd1znV0Txt5HYFJenfRTSblddFSNJUDavfqfWx5jjAt/6E+XxgD
TB4gdaKxaCU+sfN9p7A9nwVfx2JxvSwpwHOOFKJw+DQ7MAL0NSOlN1pGzFJBhYqU
Akgm2nQW3PBm+aFMxtuDzpuCH0rqL/3UT3vE0PWb4SyaPOzmxcIfkUnu9dX7yDni
6vdf2fKVaSv7Gvwg9KW9dVl7mFNtejYzKFlW+lKeVRLuQilqFzXn7LrtE+KoCUd1
fFtGn0s2ZQYf/tOBRoNHa3xUBbNp2uioPiFCswT6Afe/CXKhGc+VIf1Uutgy3+bE
AeHA960Nr7FGVmpX+J+ng6iMo6iQpoc6RmBaKcB2L8zSNWt4Zj1KkKvKXDX8Z/2X
g2FvK1t7BB+okF+/cz/3xkykxwQ64RwArTZslzxa/Ebt4PtB8svB/jludmwvzniC
O25jm3ACr/ShxtkpHtWs5+IYoKeEWmw+FWDorAbdUA4aHfXhssJzr7Ml23CrwZMb
RsQZZPq8J6br3gPmmfqcMxTmpA8g/CJ11JB4S3v8kN4IX+j+dtnrqADhBgeh8QGa
eeSmx9FGlruTnK5Pnc/luvyJC27ySsrfVJYcL3boT6WgK4pw5Fe30TGMJGFa6vIF
zz0JCgNRhN7/E2t/4tTPiC0OEVXZFUbds5mVTf/pV1n9tASP2P4afZpnGKPGK2ZI
p+pA/h5UerxJxJitnOJEKPSO2FvlA8rxQpWKwVdsnCtFqfNCsDX/Uc+5xy9T7CPc
bXf9ZFLLZlWhey5aqKmvOVlQNhz/Qn9yQq3oG/s+k5gIObNO0FGFdKN+JuXu0Jk3
IGQRocmbIf+CxeLmt0rlyHM4/PosH7sRxf5QmSxzrcuPbQ3JCc6SlQOrsvaceULG
v4wjILSSfohrcLkWkYa3yEnOFs29Fc9A2E/GjBoAgUuDnckcelgZUbVAVaNTHdMP
FeW5fxkJg/3tMcWI26iH1jRvdCsw09Ss224a7KF/mzlWdyx3fnEea+4EtV4ZrcDu
xKKlRMzESaiYZ9MmkEChzgAIF9xda2NfniPvULd1oMAJaeS7lQn9OMIvMoJEVOrN
bzVytHjKnwpHuKJlDCF483rqCCssrMnjvkzGWWipG3C6Bo7yEn1F0x0EZJm2Qc4q
iUpIPU/m/sErzbsUdlauLoQvpVA92P2L26nNsTEugjh1KRsKVWxFEJlpzcSgGorC
Ckrmy8Mw2h8yxb2LjJgbbdoUlnvSyZ8pLEiczOpKzW/a0hXRUI9l/4vF6+y+n14m
QPN5ulyK8xFS7tDuruV7e5P8pHIFrJreY6JWpwVy853Pi52nopjcCQPiv72bdxjJ
gQ/a9MvcnaRddF/k5pYFtZj+6arKY2qrfTDKdnDFu14XJ/DHTqaffjhLLXCAmbfz
nNpRMWM1OSNI5Q2VWupEZe5mVJpu1wqXI8EuOso6nms69w2uP+QMWMkjZRYfykh4
BLmNs8YqI20LtDvDYd6H12SgHJtnLft+w2iiUfMdfk1UUnJRiD9OT8l9Mpz7iWwd
MECHZCLpKpvfmyIOAnE4CaZb/5PNz8SUObRHq1VbDgWJXJ3Xmuq/Inj1B86vc3Vp
A7sNXxf2DR4kXxr1IhYhmXnLlDXM77sGn92zUNoOCob+Q+0WEqblpfRetgHzY17a
NgvXaBT+vUz8fDwx2VYstuBGGzzfjO2fO/l2N+p6ze8Mxl3d3Sp/lXuf365iCf9d
CzL+zBLpUpYYNd0sTJZ7EKJzJhGSkMb+lMwQazz/IRLVdLc8Xm8nl3tKg3Em7BM4
sUTEC6UP7FRNPo2sJMxRNgFr0V0i9RgstFnptXbbo1h2XYMCfZQk/bRxURh3rYWi
R/4tR6I8dI+P4SVN73KRLnWxzosfIDYP0iJH1BnrCMyhGRei2RTjpzoMCy9xjz0S
0WzW4GTiayaT48drRzzPwRl+Qpeva1NUREAEBuawZi/2/5SOKo+mryBXBeTgd47G
uA5I2hIMLstu29KB1asjOas6vsie6Z82bhvKAgmmXrOohSqqeCkn5nV6p5HdZ35N
bu3X90sIiTgUMsAMQXL/oynj2teVXGpklx2MSNtRWjyyzmEWME8I6M7vqpyYOueB
DtM8Ee/HoKA5LJTRGET4mg5Xm4IqQA/FjGwzS9+Ij6guJW2o+qIb7k/RqnUdeolT
j+GQTojNxTnkOJ+2NoQtCLH6StNZaqpxMmzlSK8t6oIqJ5T7/X8JC//j9Z9+ZzVx
W1LovATgifRkseIpHDvH/qIsH5h8kQVpLMA9Xz//HvKCLUAMmJ2R3d+8/0OyYUsM
wB0rdUVj2SosHqtKR4UbqreiTyX2JfZ1h/iCEYOda9JlbGmSOG+remI4PGCMB/9f
jBxtgArBQkFZ6/S0/Nr2FO3ZIYFM8EQyo5ZkNi0fFEfBC6of+E1ElNt7VVLLUFcu
7CvUCldFVw+kdm1lQ1O2SW/haTMVma3Y0AFv5uLSjVqVOMLAp76xOXo7OGtBnYur
gbF3x1X11NosPcJxGhE6Vgk98WZLJ1whfbHxppyfa9DFz8VAJ8PFP87zGNM4QSAK
4/THBuYUfWdHkuIu2yWsklVJ4S5hAAB3+0YiW6+zNUaROSsSwQEWb2ODK72PQ2rL
pihKu6kw9NBbSnXD1hiLpBHini1IGyV48LyArW75b9sQM8MYTfw7dWoNt2NtYRvB
meKXEY9Ji5c19xs3yXLl5dr8J4Q+D4Ds/+xvRVwqQ0e7HFr+dsokyWfpJXgE25T9
fCKGye4QxEPeWE4ipX69cfSeAfkyTzWidOo4OXmZZqc1UR6wP8ytjSmgebpQT0cD
oB6ASfcROEP/JXzn3z+DkKGYSXLzjPjXg1vkMv9JuGy1OmSorF2JgunmLLttpwkQ
8lJNTtADfQigQ3wjqMlZKbqCRe+AVlpxjMwdOgmQOVK5sxrPnCtKdFsmZcaPrrK6
n0P+iw/etWH3xLeYzfyvv0EbsBQV5Q685mKb5Qz6ghxhj/9sLwb6ED03RbT06/h2
ReCYQ/emBDXUITRKvt00AiZlG4A3up/XsYDRLqL/KP/lq8lFwANi2pMpYyxlOiRe
TBglzVISaVqkWU4/+Fcdqn8mDHM5SeEHm7pJ7E9AcJLK+gRScRHdnQfEau/VkGO2
KVqov4g24O1eMNcLS9Ad0wVN3cpEYoRQWH+LQMU3HvH3D+G6MjUFT9J7rUEd5rnF
iZWvzcOrK4mXEHyYKyS/J64Q/t3qk9ZBTvHLi8o0WNVW4cHxHDNhK3SUsiN5QTHc
Q9eq9KCcPGQcR/dGOSpJZO2mQRNk/WBmkyTa5dm9Wp1+rsQgwsv67Ifrazll7FwO
+zOGbkB69VdDYJl2mTUUkLJTxvIyzVkMPkgN1icwDVDqQhOKXHu2FZpWU79ftMNL
X7iGs6vF0SnwCJbkhuT05bsvpRBxWxFJAsbAEKUAuRvqxv8LeJ7hZrOidTvIwGyp
vYIvy+VcgCntaYRdErXP3giklaPcDcQOjXLi6lETWDjPz1fAP5c1Xz6ZDNn+UCrL
EKTRY3/xKzVl4F0kbJcOaU5ioXegoB5usidcdkBbyT9JHRPKOcT0g2YA0ts9tbN1
RuO+zUm1Mr/md3mu7g+0gRUlIiREz6hte+3Ib44GTmqX56fKb1CQGBdPTlm5PnRr
fjgxS6CHsTpO6fxJRm16lYcjjuOw7QSihhzDpqDKel4j5l6NMslC2xl87ogTpGak
ydA8gViztkrZTOGz28q/ysKJMxPqWvvahAAQVV3E3iXxOLpCC7aZjwZ46Z8zUiwU
rN1czLiFBX9LCRbTMngTQGYA/wh62WIMVAALU1p/BYiWkrpEZpSKxV6Axr7wPzej
sa+15VR32Qst89qtpceWIbzCPBriulxcheaOPSGfc/TePXPBoq0lUUO5+5rSpEyN
GWkFxbbaMO0QPCWkPgH4sSaebf6EspK7U2nFo/sFJjaGBlVyS/KmUpflXgYqW9w+
lJR9AYE8nNzx35DSvg2GbCNSMBhvl3wDTl2tDjH59IohzteGKcRd8F8Fvq1lKLCv
8QZAF9q6QKbrT10IehmAbt2jY6nsuimM6p987qRm4P+2YJlmcHADrSlvaVRcnvzl
vAMY4UlmzEIeWyoDMXcbeM9PpZASh6Ye/r/L5KO6wpp+BZPlD4/zNTpW7FJLqo41
f7cARO6J6ESkWEVaZoIsAtX1rp2Apl7ZMoxJ1mvEFK5frrvH1b/gkZckkmcDZpG7
T6yo9zvANRe33L+1KB7+hIZvzHZMP2WuvfDw4J7sjNQHymStiGxezDfcqjcbAvpa
sasAid7Eq6GD/WroGSlfz8IIYGBbaL7WlhOEcQmkTUXO6hO5krO5mUqPetwW+/II
UwT6BPpWYKWqo3llnTjItpcCl82Nys1GcUqaE9Qcd/TwS2XinKv5Ho2uJpIDsRiN
TXiqgTXvO80Lvc0Vd1h1QMNLB5+WisBWGimiTvGtZfGu8E50lzp8XByooTrRVY6d
jt5xBYgYNWT9rI21cd/aSIIaPbxG3d63j8BAjYHIlauc8Zr1n+YPZMMGzBiozDea
p/+u+LFZPpqK5gbmNhPmbacaXVtGYWT/8uHRcogJ3J8D70AG5X3NyFyboK6Lu729
sAapBqeS2roSuyZ5fikSDSIZ38ZzT7MgdasAIwRJQr4Ld3Y/S2Dvxh/0X8iCtSf1
XcMEKungH1PUJIEFQkOuTUccA2lMQ1YPdEemphTNorN5I1CH97R9DPcylPEh4T/G
cvkiokkH5EEtjhvSw321MjAqytWsi1ZwVfWVoJ7BJaIk5MZgEBQcDQIA66CSQTuP
fWLmQhtCcDGg2Qe/lZAwBgyuIvsVNJTI461QOdyC5sh+yoHIbhoGcowrNx5uyq29
56Tj3Lf0RxOtLCBOlOPI2tho0TwsrfTdOaPqnvRsLf6f6b+CGHc0PDRRAfqkeBn/
rpB7SV29wYpVeYwTOKbJ/+5D5BIX9qLmBZeRtx6q8Ao7unH6Jya3yDxTOVelq+AX
SC3/O/j5FCW1DzPmH5QrQG8EGleq93r6I0GqksTbeBzXYhNCSM0W2hN1VSWVPVXq
Ikt+2eG3IO0nJjNXElRHqmvfSlIBq57LmLxgc5htdCzwpukRKAEKWFEUdc0b5q0T
JnWIlBGNBGd5aoW21LlTI5Ez7pbGlHRLTaF1qkq2aLkHf7Yw/BoeHwyg93rn2ouB
iYu2dJZUkcUILjfRxGrymo1ZeF7SmXqqaJ/F0gxqsqQlSiP0CICYRI7IhkJ3lLw6
167KgzoU7jkqUZtuA7RkWVc5DYQC5ovAVuK1VocOSLsn3eQGNM8SYxhrMSP4xoHr
HKgLCc2obXu57rLjC2I2uZSYbls3Bz13bHQj4PwftvZiyTNhdIeoou7yRy+LfMD3
AWEvoZEagXH75Nbbe6rg1CiLKHfvudbRZYRgJAt1ChVdzali1LYX20wU2my9sC8C
1GRcbYBbLYpp0+bugPZyI0LkMJLThRM2XU/r0/KivWg1YRG+E7TK8XGWicTo2VOP
1VMYuidOkAfepi8GeMBdy5mj0KP0ZzYti0MG87+kAqAFQdYOKgwClumZujZr5Qor
kyIoCYLgXXsT2Ulhw7B2afym/WOwD5s9MQiXIpU40rfFzEhrWsJOdhrF1u5Ai04z
8vuF090h7h3Zt8CYX34M9K4XiG0FFX9tnd1zI/TYG1JEgxcgM5c7NPMgRqzZZENE
aCoVaGcrckaup/d6mpYyI+NnFHUVqemFDfAWriH7RMU6v198SRpeCgYjHtOKx6sf
XHy/Y0RtIGnWAdgAMGQW/HqCDKxJiyjeFdLh+2rCnO2chDJDmjEXbQsBZoMjjfYc
iHny8i5x8EIxG95KsLL50bogN/0nz1gEkJpBehJAXkoxpjsC3W7OcuALrNBxCv0m
MZPQRyxeT5lDM0JDBw1eQooyxkspWLcGKCp2dpTGXH9b8bwlMPtKNt5WYn/M0OdD
lYsAcNFFdiRzYAvMs1Zb7OTwZen3kA7YL7YyN+emXUg7jQ6NSyam8+6mxq/7IFUL
LIspyl2Un6maPIHoavtV/kYY9RYG++ICoPuR5lpqWXyJ5VlLMyd84Cuf3xb5pZpf
E/oG6BbfWX3zyGAunFQavURYu4OmKsdb1kWf2CChRThPRlu9LRa2U+JxKOTv5E3k
hL13hwAI29vxmFV8pDzpaK/9WxkjxVo+a8Fzw1TNu4sbvX2nRXEpuIjhnDcZfQq9
s5ljvazrxqtSdi8xMIPu6+u08siEosBG7K6ta7LKqP5fXm2bSRGroPQeYK6INiVJ
ny1n2nrGZjSg/jpSmLjaJUMoEuL8o9/H9DKBUgQmKvTes7+IknGyngRUuE2J/gr1
CVuqZKP2CAr/W+NS4UXu5rzqFYDF4iycwQzfpzfWKesjvuOAVUggL4wOvumPHnEW
5N6NoLChacuw3eTk+HVs9s0Rw/rRnlu3lyK00iFam8A7yN4zZeh/dztrLWis3/+d
Svi+EQfS/9NRRnL9eXjMncArAIJozP3zcmhyBXTfyNBJiGsxNWsucmQ7EYzJ2y/7
b0bv1Sjau3xBeyN+2rubidUFl2EqjzU5g9+g6jqqpOzg2dAVR+vAwlN0P6Vkqg/G
CggYfOmyxgMtB9+gjNbzvpSsZ/R0lCfZfV7yajC+4KHjpTsk6TEUpa1pO8QRQZCA
coLm1vGKInYK063I+7adnk32UZU5aYwJtn5t5XyBnXTY68H+zl5yW+g2+7i7Cftg
t8SmSQWIbP5k6kXA1NBUxZJJL5f+FUxpWuMRGiHnfgEBi/fZtIaJLpreIefwlsfb
fN4ivW4rgAj+SxCOXakvn4sw1Nhl4qLGC3ENA6eyNyOtqQgAPlqV2emcn9hJDnfk
JjkQYqrc+ipaqj9dhn2XB7yeqcU5ZrzHdhBut/ezRhWRVyTZXg6CH8fnQUK2pD2d
+tzPT821C1IkVSJn1pC5HRZCV0uyAq9T/3tLjsI0YhljGDx9ZTtB8u5cgADjOcaV
2Q9s4NoMbX7D4JOhqcAqcJf9CydDy9qVAqT3EHJvG1aTgJNhSMp/gHS5RY2/IQpv
QfkAWf3/cK3o84azSibfU9hHsmP3WfRet15b0VhFR1O8cOARxCu+wN4IsJjFZalu
VOnuyhs5Uap9jSiVNcuxqfqTUI/C55s85me691GtR6cSvmed9T+7LI1Ai2d4URab
v1lpz/NlNrk/FdEgOuN/HkiM8j3NEMXtuUu/kfizH02lN9sErz+/UoUj2ZsfXc2M
VnKvAfRTS9xneyxGihE2oXGEvk4i+srv6uBWJxA13dYtWW601oLXUR8evBnZjt7R
0YK45TXd0t9ckThuJ9cRVWPkaM3uP9BFOWuqrJfzyttNT1brbOY4pVFrYeVH4GuZ
b3XVgjDodt3mpGPF4YYQ+kf8k/tuqLKrm7kmlEKUN26QLy6Ca58qqCbos1fwYr0G
JzheVh3MwpsKTzQ2ZVlXtNl2IvmelgkuekMZpSMfwV/j3luW2maCA1BqCkfvSq4N
jiXCcoPYWGsW/gWUqLQyDEyrPhHjIQeFhlHDu5BagIDtuRPBQTJdTHgIpFllNgTY
jwxahe2GYYunX/IUlP0tL9QLqjrmX26XD2hLVzJJCfYhJKjkQIYOglLF2MSOOQET
OD/HdYJTRlrxaxUR+o2fxr95aAkRUt0sAjX4qeamDpNhG/90yQeHt1fjdB4tljl4
4WqTRRANO2dSPqXj/dg9jig5A6ZPJztnQJIJnBaKzI0AaLIShtGZ+m+Wl+3RWoXT
GDvuU+yWBI0zlr9pU5/wHp7OEpU0xCbZ4qw98rPjEg7yLzOV4CWeGkeUsenv1Wqs
MX2IlDhaBiH0khHypSrRhG79Yyle7SJLSWapbTrxGvL8CI3r8/mlj0bb5rSTGmf7
oTBSKKA5qnU+d18yCt3TJU6iovMEK4KykmWes674sW3t9Je8qz+pCkIXASyX3AIs
oYMrml1akVul2Kf9oxv2PbTA9PMYT+rUJe8XVeQHbYxhCB84ml6m/1xh4IgAG5Ly
5Az40fD59wZhR9r0sQ/5xPW+G+RAJlkSGlFhk1BP8MWVPT6bh0ZfeWkPrsfjHbWA
zw/klhgqMLbbObDVskRscVDAPM2ohKL+NxuLPNLsUoTD/DnDCBPy2rUm/TcpTtS+
XRS8lXSTdU8ZLAMyd+2Ht0WzgESdUzToUf4Uk4rbWnbP1G7mOjKj1GdK8Y42/M47
oNYpTHccnf/8ozGrNB6Lka+3fvvtC6AaVL7y1JhfgeTa+aiIjHCN5+adErPfoj13
ehgduiUgoiL2hQmq/hQ/WLA/Z4nk+SwoaaE3pzXeWVenOGUxndqF0/4sn3A+J7fx
+jRr2RkIxy6d0psfPtaJZ4Z1FY2jdERkWQEEvYNB2/qCczYl5uR8OVmLzmGRMtsp
CWb0qB3Iukj0Uuj4HMWoA4VYLR4glMAoE4u1qRDjLjxGXW6vl+8AOgLUd2NHLhvq
0FvcwF3NMyDkj+ULCupVlowutzvlHf1JrqfhCvWCZn7OzqZhmZVcQqiH4cVQoiq5
++c7Ebx7CGR99pvl2TE1Q1izy2fz9dM9VYpWanCCyntYWMSPVdaVSC89+sSWCtCw
wn2Pw/h/TSASUma2z77xsSurMg+ajc0zGN2qgQsGRRZOOTO18M5Q7/f/ijQSa2FK
TWrM9Vvu+QgTOsHHFJl0pOMvcxpHTsoXcxbApWb+fFTUcMkerLpyyT7OlC7Qt66C
Irm+RJp+3i8+cKJPiFSk0RtRYah5XMy1hL3EdAfnv5IYXgfuPkBFNkGnenyA7AB/
rp5bIDku8CNypAgJD/PiqRBjiRudG+pBzNLFUUJoobzc3KvQU/iSXFywxqII6WZf
tFHzs2Kvxaq9GzQfVQo3FbJKXD8tjCO2lO/TBKHK0My+RPBY1aNb0Pd1Aj2GuMS9
rLgby0d6EfNec9xqI16v9ssRuIBffeyxAlLzjSkgJj+Q+CenfGlq6xQR75xKCywd
qqFp5mwIS9EGRtDgRA6uFs+scY8kTuxz8+ezYhTPuAQWq/leTuakucbmIMAfoAXS
MqqmnOFek+e3qYuMvdLwm3yMYSDt5GlHUnwbgedyvOY+HlJ1Rq6NWYHJdnfNsZyy
lzaZinR+HzrkcHVitL3rAoN/doK597ooi7OOnf6r7LzW9iPObc3IEkD8Vi4944nk
0nLfGikmopdjQRC1QK/6v0LkDB3fVRZSTuGl11LEUptVD8u3By/55L4dIaiuUDtt
rb3pcl8MGBp4EWLLYnqHyMFwvBLTboN4ip2J9a9DEg9zH05ay8fAt2JofjYOEFHV
cJTKDiGxNSUXHiIXuLmlFp/RuqwWy773asMt2osLk9hEGlWLMf4V6r/jBhX8temT
N52cSaAD2a+U+r18mVpfTaPi2hIgHrh2qmiJ5vuInP7zmJwLtdu8aRZ9JrRXToBL
rjFlZU7FwZ/zY9dlptNajOAertIFrpn51YGdEMe5B7KdUASC7o4c6ZAISUSapkcQ
NsSw7j98xPtJxIg9HPA3RHVrEV6i676G7fK7vb9clxH9ebSQkl+zfyLptspNGzb6
YVSdVHD1knCaSZTxSrqbhrVdXxbpIwNgsqjv+Y8uBBZFg+gcwg8MO5eeyuXAGNqM
3wFNz+0Q0Y4UGq0qvl7tbCOpQfF2OSfAozV9U98kuc++SAopKk95DA3et/PuhYeO
lDP3mk6GLoqeInnCHwcBbs9WMjUgkl1oHA5fKRpGZA9p/Y6KFtpfvoUjEBcFhF3r
RfprytWGOEnZLsQ6e7XctBNYwPq/o158wdqXXsZ1kSAkyvqa95n045BqVbOiGU1Y
kActoF1k4ExHSRXLCWBoS0T5JNN3tYpfdQ1VSEzq8OYDKj74rBYIbpHDU9rH9iYD
f0OpGWD4xfVNVIM4eZzXDMeP/yZwNk8UNmijJGw4dJVyq4hKm3bpOvmxG+OOEOMY
a2YsyITfQY34jz9S+YAt2W+WOhb4nc1FpdaGPb5MWuZlr7J1iNFJmQvDW35Tt1p2
9VbjsxWRJP2ZvnVHH4pJQuKLO/DCFRLQnH5trrFHYJnO0DEBh8+Ifrx30NM6ps/6
cfOdTPTcgLxq55imubaTSljF/DWAfkOHhpSfffg8VnwMGImy488eajj8WwHJ4uwN
0oDCJCXuQwQUAN8K3UCii+7NhEnE2L2EnI/8/K20OHJKmQPZYpzYle0rSFzctKY8
tNWWXWsNu8wSbHfZ3i1ong7N09X+Lfh/udlBmpfhSXAKJWEOauWwsSYD8LIQ4dIV
MY3zIazzjXf+q6cfQ3cLXEUas2S6PLsS44tZgDx3raEzv6BcH49rOLOOwmR2ypIx
gPtfUD4508rktotwBP3Pvd5LeNrXNIB/8mqqEq8KBB3OAqX7jp7GoCIcHr+Xq1Hv
GSoRvHz74zRBfgmL19xnerUIAvvVAZtN7llI8Vy+dW6uLdP3QmhAtAGcmti+Sv6i
LYhB/l9+RHAeUXpqWehEUrogXRMiribn+l6VpNwqFmWWrC46L5Jand7FEDQx2CRB
tDzLorqQwJ2rJPzEOkbjlUMro+SeVk4xqtU7xJpOkhkC3vSEgP36YhK0pvN6HFJ9
WZA7kXr9XLUEPRmaGEYvNGNVx5sZpkVK9wIrPDlIHOhye/Avkpt/Xr03Id3FqVyn
RzkFv9vCmFlgB+l7YK8bCqXn4Xx/Y1prU+TKPMuw7+kfrs/DsueXbIs7PUk5FOn5
jKhZ/pYogeJe5GJlh+lNYuZulZ1a5DSHMfI9BUPys9gtjG1Sjg7U/BBy5EPOhlAh
1StttTRItyT1TxqBgTLMjCIcCvBu0D5dlit3qR97N60GY8s+PJ2vCJpJvjpGkD48
bTqIa3Wzb016byeylzvcsYVoD5YpLwyBYUgGqU17eRVTb42r5tzrns+XWj8Tiv4v
5JOa/te+3q7CWs0Mo4VB8yWvsxsH9/HwlJlWrn6aj3WIFA4+ezK3nE/vXiTuxFNf
dle4GmutQy80lv6RG48MmfNYHbwKCZEydM1vDQQr29kPntwwujl2ucGnI5sYVhXJ
zTXV0ByT350QU1A2udrCRYHHVMJ5BSBm5ymEF6TKsg6qwRff81g+rSpuErFdxt6e
nEYmqEu3s3oGrwr1dLULdnkzzhU3NwMLRv4qBpKKVwY/oWLxVQsJKDctxlO3pChA
VSL411F3QmOWlMKDpcvbsxPFRycCK6y9QOmwPBKB4oWSzuPDTCS0l+xR9od55adu
ibBO48ZvWGy710DgSheWBc5MotkiGF8r1e6emVwjmAKJOH2pGowa36sUp8LvgY66
1++0VZcblXxDLsDt0FTBLCEotg8kkICowCUfnzx3+OIBD8QfBOONRXfbq2Ur40I/
TK6fgKJogJmXnmgD1juC7j5BAREyWYHSlepFbMQDd1bMBYOHaP9vgSUgtRozVx99
YZ/MflnDw8oRuDeYBvwbpjJ9m4rUHMA2rpIlqDlMTtBBkwQfE5nve5xpTgcTA2zP
zjyFiV7n+vOygFn9EqboMz9UU84lUDAhl4HUDIXNbVsnfhxqY12RlFl71s8HdgdU
EXqu8YY/4tBHVVoobF6TIShKtfKbd7DxgjdyeqRQl2FrJ6MSVkpFEeRkPBZnk0mL
pMIsI4WoUUmcnyTZnyooHIvkecyO4eKb0No0OcNydp84D45/USB0ShOWIlXpAMcN
h0LiVnjDfQRjfKrbMzQx9vLw/gFhNitk01llPc+Zb33VMYO6VUCDAwhn6jlX38g+
+Bz3nwftg5IKDaiaEXRtGODLQeTQN42OA9KRWfZbH7trsYiUAapp/6IocLbbWlTy
ZNCihlkJQ9hoOQw0IwCBkE/E21or36q9y/DgIoUUtln5C8xOA6hr8tgAtZKWXuJ3
xn2xeeYqxkvVIYXqOifKSO5zthZdyEduBUUK9pYr7g6Rz1ZBrczO+vO1iTHglCcv
f8XFs+JTEe876ARvk8aJ+oLIOY8RgQhoCms7zp/nCoGtne+VpMaxPewxWG0PIDz/
cDPIU53WQmPX7va8Hb8v1QVctUBMB/zZg3g3HzKXkSEDioyV/UbfnvTxAx1sqA4f
qk85wjUAx4ivlIs3T2G4KxleQDfsLgxoc5wnwowIzfR5Xi20g8HXwEkJj9quyTsK
LNqodR5hsCS4ya5XnpKWrOf7vtg3aX9aICtVELxf3m0PbZn9K+0xoHgYvpuGblEU
BtB+XGZh021xcSudxkQbPO8UdJfdb081CPurFeS1uvBw3irp2b+1nE/+N+mWp7xW
Kx2faexIYmXf0IzlVivyWPEe9R6rzH8IqVVrYw9GR16B8jw8rv7X46h7kibbJQlK
YUlbw1ZAuVNFxGyK1nMvPzgImJ17VDa8Z1RsLlDeBwoyJGI8PYJ7pTSrrDAUEi8h
tb34I8dmnZpb0LjfZ48tFYmdqM3WHBm5AWi95MB/q1B6V1BjolW3wJJyE3C+DK2Q
V6Cb+yVXGo1/L0HMcAwIzEfWJ+wP0CyhjP5f2BfNdOt18Ew7SsSxXP87bf3M+wi+
zO+LKBnaQkZB1ILAz8h45JW1O0cB3ivwMwHcy3VtipCDfqLOBNemXIzmq0MIAewP
VgVhzddwB5NGkVVEx664kUIsW29iurVdUDpPB33ULmzcg3rfO5zpvxTjrCUiwuxv
XBnTy6XdIdtvRDrsCnBK634NIm6Bc1IBCqGATbYI+DBC2nmML4B3YU2DD98VAsDh
DfwtaZi9GG/6UgVaKeHIHZhbVaXgsibscHfPq9JbKhb28acDZ+PZNEwPZ3ER/Bu2
SoPF0e4ZqN7ssxEUchyiUkLul47tJ6FIXBaeLaPf9ljhMDnr61AnLJiFxPLxnata
I3UcfSTQvlLhnlrH3hxNUrTQLcy4gPk+/i50cpdApltkcv62gtVCZEJ/uG2uXWMf
X5PYJyVVl8W1qFWOrHcv/0VEyatlZV5Er/8ZgMaWcr6CgtEo6i81+81uv9Eypmpu
O30AKP4jk6ojbfRWbYBpBuVd65fgWN9IpVVGmHvKiSabflIRuZEbuGAyZNuk7nJy
SSSRbVIx0QUv2Jt/2NEeruoojeGrPncSVrhanzXcnY/ivOBoIGGWkaxyz9ld+8mp
sOioCel2wkcLRvrRaxvRt8d1p4c7kXb6ZSPHQjmhyCxsnqnm2VG6Xr/PktRuccc6
QRv6mHuN7nJJfC/VWE/xo7WyZBMSWjv8C7EuQcZ2FeJ5LqxHBddjmPL0PXLu12ci
090CO2BT8HogI2H8OaawZ6mxYS35eePRTvE6GkPurLrxePQAnPAtjduxLpKDsm3p
DgOq5V8ysxhAuf7jvXYxmnpFHWleZ92gyo0oY098s8DoVoej/a40RYzoiGLXDS2a
vAnp2ljHltTiVhsJc8V2E1n/tpbRckne2qwBzQbwvDEk+ZSvnAKyHI1e6nLlHuK8
WI8HXzEBrm9ixK4H9L7tS+t74xXz03pFcjKJKkVp8Re3z6cPrfFpxvkB6NXSdvGX
W2Ch7v/E8FxemSCzDLFDKKGpx1EFVjGllYuixA13VKtvrDJnXTFiK6Ir1Nrkr2bi
HZbA0Dp0odU/whAkBYnqc+O/lgbLqsiHop4kuIS9SPsUxI5YpZprjlfS4f5408pn
yKyRVjxSkgbNrqshvAPxSEic+MQXwnendM22swlbUnU2RHIXPQAYxIZenbNpvq13
kUba2a6nltS0R2x3zYYmPIRjKyMGxR0WTUrXKfWHApLvRA5ouYeYZ4Phu3yKnpa3
en0zG9bQWQ9/d+PoPIm2UCMXnyp0I9b1CtH5vdU3eoFNjLYSE1hpwg+YA5c/05lh
aHIVLCy8lWuns7iubo/EqIJaKuJb8oDYUy3J9V0T35c1ykx6T60nT9vwWJ7d1Cty
Cyu9B3zf+J+g4tnxW05uMm231OqdyYbCgqDhCQfMsg2IY6iufGc1VY0mkVtWHAUa
yePvXRkukxMVRjf8SKHfjlpU/j7W1LMEqZo6VKyLWW+Xe37uL3ofeuHvjlz5Ui6w
TQUlJJ+/gRQufi5sKUvZ0a1F6d8LfVSEEtSufs0EEuVjYiyRtGQABOEsraLekNc6
Fql9KVDb6HgloH5xGmMBrYHZZuOpjnWVqMmr4wzZU7I3Ot6qBqir8SioVGlfND6c
yh5ZCtL7Zz7/2jp9jVsRCkL21CYE10QXrIRaO86z/evOsWLdqtn2HQHVfm97fY9a
GQhJ4uR9zY0l/xPEruXIWTaipAs//kJaqFXqvv18hV5bUur5EzYesNecB2IMpTT+
O5cR8o06xVIwpdIXjFkol5Af0dXQBOiJRi4hHhPuMczZm3Z3X6pdwdx9O3895MKq
nr4C/aTG3PT0DA9KYahQaNvh7m01aEAcqecL0C5rQjx5cTKcol69ctMab8omOK63
4a/CqxdGmwVwPdqK9EJJgpRS5UAiuWFd+edcHpOe/KKymp0QCwZfTgCZLdw11lwv
leyb25pVrrhJ0c/h6R8HI/3jGD2XCq2+PHJ6BgOIQdjhKJrphqZyRO2JxnwK8o+B
r4vI99NEFDSz8KsN0i1i9yi7BaRf6PFmHeegql47XS4FTMokmqGldvFHMlYV4JML
2kmiROenLo9cS3QYD6Sgsdy2y4uclBvDfdeY20nEFamUrQWrbMKhfXgjc2mkUt8Q
evyrc9m9X6Ce/L3O6W4xJpp8CbVk2Afcljwmjjt5ZPmyoobdp+HVUAb1MiYl0tz1
/Pdv1SzeYICPvAMBD/yR0xj5hICV8MLVzS0rQ5L7fUBK/z3mSPXj7IS1SZWGED3C
zevVAqfzl63f/SardtTvv0+tpWLfBahQWorzLyQHr5ia7UxOrtEKFz5Uwo3JME+S
J1pY1OzndQhBRfEBH9aFPw/jNW2T9pt2nXCpfDOh9v+f5YmT6YcWgj24JAWlt/jx
e3OitgTv0/ZQ3bWtQtI3wGhqOfaWNBgYx63gCeMrR2ugGoDvm8d0HDwbgwVfT8pz
edHwm06eC6+owk89DiV0AQAtGCHc/YU95hBFS8H9Hqi8nLuCqh++wQdhr9Ltx9L9
89ghmr7gMoHqp8grTSjqVSojADcHWT7POuRwFcT7Sfnrdf4Y/qzbvjCKFEfV/kC9
oiVz+sKqPevJo8Q/AdeYFnb/m4Urfsvc0n/GuEPnuu5QyFZQjVbVlsMsQ59Cn+Co
K30eUStPrYgLGzGHg3YSkUcdf9U2TXMjZgAAVcXIXu0MEMv8sOOvU8W99zu0p68E
3Jk8e6YL4j8zJVR4HW60gu8Sw3E7MzcIsWwU3TOlEDtffZSgL9biRWQ5xkGgOYOJ
iVEUMTeQ/K0VQ1tKPBH77+uZ8lF8w1IXq/k1fFFb/a6bj/TANLjC2g4jHE6BPfuE
MigM1YnB+Andgwi9tYdfLJ1lrD+0b6O8H0fB6aUoL5hMxpAF3PURKMVrn9LVx5rt
bSlv9+9p2zsoYZYB8U9ZJBmQkLWiq1mO3N3isdU6YbUoD5AX6nGv7LzqeZB0Z1vb
t71tVFcAqCW9qKiZ1q32HQMExbJacvZaRe4kwTzYsYG3UgRrH2PWKlT+Yry4C+US
3f0doP5DI4TdBhy8KaEPut8olvD6Ib1gytY3bgL8S0xWALMs4G9DWzbulG2I8+ka
LexxQpxhf1/pFvbA/dmJPLstNB5V+vNN5OQPARI651x66CuVL0+rxGkralO40ocn
RbYwAPyBFzHDpOtTBchoA4cS3o53MgjP0LBqEpESrQdCaOqVq/xfcLRyqTWL7KlI
yY8hyIKXkyl9Ys0g1dYk4WM3DmZub8fTbFmnnTIXRFtDIF/H27Pvw8EU1DBCBUiy
C9oJYhV1Qj/5UhnaQrGB/znP9bN1e2N0v0POY/qTR4Vb026qZ/pzNmB67pbBNDp+
ZCBU+olNPm8EFt0kdZd3ajMSkItKsqafFURfKw9qrH/tGng1E7mNZyn/cvd1/fb1
yl9bIx4f0rms5TOQmmUz2REdQPpm8UzP+y3pcPIzo7/vzAYzUC71D0lGKSpk4yER
/YmS187vaw694EtGHCLk4Qdp2nI/lyOARKtt/fo67NWTpKVvmFq8mS2NR0hmgZoZ
yo5+gWyOSd29oNnSShFgZyIFQkVq22rbdyQdte3CZl5watnIK7kpXC8N5bDNYlTd
pOs243Ju5I8MdJjVrXA6/jSAq4YdY/aD6CZ+VPA+u7jfMIvvwj+j8Wem3jsnSeeF
wAkwI4uGJaX7LeTwYJs42TnFXUfgKHE/NJeAs6h7J2ZCjqU7K6m2vTjmCpGrHG4a
DV6fX8acdDg7h2x06dCG4nHgC1O1OPN+k4UvQ9/Q4qIoEvT+JKAI/byjbH8vmwHH
Mz0dftk1FeO34RIwpMe1H/ArvFVWdVnFrMj8hyQX7DzpIAbWwKY+HavKkLSO1RwI
Bbdbk08KA3BOaMCh5JAN462JiK7stcD6XLxmmsCvZLBVgNaohh/A/d+0Rg0mT75L
deTlny/bF6L7a9a6Dex49a0volV5IjVfL7E82zl/zb/4ib8xNBiVekKmy+J3a0PE
yKPHXcp0RbP4fzJlluTcovWlprzxIJ+lQcQp/jjAVi0sptzIZWUENoq9paiL0F1r
u5vcUVzEydJkKOwNSISwSZFNiCL+haJizMB1MjPetWnJx7kRZycCvbfs5ABkE6L5
F9X3c1WrNnPThdo4NSrvde4cO5i8CEWeeavWrCl8RuMwHVkHVUJEzz8ZBtj2Vm0A
dxqIiVL1v3mBkX2ZLeFLAH7BOEoDgQDqqthbd4NjAlZ4u9C0V60A5i1MzL7itzYT
dxg+4trLSBmfZUAzXLGX6mimwmw0JNSB3L4fra3fDW2Kuli1Lrkoh1ZJZgABofwO
5EexB5w0nJSHu2vjQsiGUU55F4tUTtQOFYnUbRGAvrZzoI022n1jNw+5zUkHtBgw
FMwj6noB6AYw6NUXufqy+O3BRw+nIoaYsHvvt01PxnIpsEJ6B0BuN9sKm6mmvOGn
vQpoCVLNVBVCciORST1u0AgxPNSriaUD36pQn72VL8RJztaGSUsssdOfqGLIcytR
/Ze3NwjoQzUPoD1vdOIi3cf64zB4BreRP0NI7DNCg7X7jzCJYZKNKazpu05vEvRu
yt64g34JjmuMnamHRMNp5A+ts1/D+cynqW/Lm4LIcZfkZHmDMYo5LZeKVPO57tjV
E3lSKY/gT+1EvCvg5WTYNtUHWDwkzwvZbIN4eLP/Lcu+HL1Dk7pg6kq0IoM4nnJX
XPfUiluRcVXVTBjlpQ6Tlo7smYY4UdE4P5ges/8b40wRPK5SG9CVo6glcywuJwnQ
HmG0B1X22lLv7iXAun72jxAOqkPybQMuoU0QAulxKZB+yPja202MIKUeKLP6APyo
R2OYsMJj7x/TNDnyKOCRkEW+76EtgLTQU+OMLJgB4hdErh9z8JbxfkZ71Ua8W2bV
orHhd3v8jkr1pPmUBc/59jzEkb6H9lUNO2ru7F3clY4E1MpXIQ8lxOrp+zgt7Elo
lGAzc42lLVawYGM79YaZvhh7FsCx8vWX05ppOgvZJBKmnD8LPUYO4JxHVVZsN9e0
UWwpbQl50L7fF1PLke2gnl2OaWtBD5k92a1Tdtuto5jIHoo1Pj5RRpLiHQox38o+
aigG2sG6VlKBoljmF+sNg2Je5MVU0dJ4oFtI5ZhkSCQgJfUoo23LErD5hWTTvEfP
DoZOi33ZRKI1bUfEA0JSUQCGSgRbTKyjdQF++NDjkHc2cb4NGjeqRIbKRblWwQGy
PwBO0XPYVkgr5VLtlyOr2i08/CHRhzCreauX3up7lQw9nh8Fv5jzYro6ixk5YpH/
PlCobT5YG8MuTBy0etKO/r+XxTwXUfdXSRsLZnjVfK6exaMRPaIzYd7m4dCdUmB7
Ua7Mf6n3zAoN65eLWBba5TEI/TlN2xZvILOGXZPWgTExmdY1lZjcZUiiF+StF1tc
1cCOuemHGdBpBfT6W+6p4iiQlAuj0MH0FDdTqwOQDYKMZQAQFJFvW+qaBzBGxxUF
CCOBOppbHtYpVSYBxcylgrJ8QLzDb6MVzbTFEVZ1Zet9ydh6uJGpjVC606RVU26J
waDJase/Z9tekgihcoNcuADJYsX5fiZ0JMAw6u+DyBDsJU7TXdesq7eEvd79QB9n
1AYFfZIbtDtbuZK7eatSr0KtfeGtZRcRozS9KMndH8Bmr0GuJJF2oruwmfmJ98b/
rUdOS9uIPdN5X2vDQ411DllipHgUFQgcHNgxfo2idfvV4NaenfC+GuGWVAAjY6MS
F3pitTzMa36fDJ1P1R5g+r6TvZ2ViPVgMEmnYHK5GnGBFJe91bKwQrAR7zOlkAj5
m1DD2bor5vV67qJvXPIZHMQ6GUJTngd69RG5v6sTIBctoSRGWq2xrrA/OugQKUPK
w3Q4VUEzDVoGLaoy713eOU62W/uM2k/AnTvQ5XzU8en9yInLh+HyCPC7nI6Gc505
2y0b0VJLTFKMyXIfQFSzCTrXbkrv0lQHqITGDkyQZngxfWgpY3s3oUPPe44fVqzK
bxU8LrWvUd9ssBSicPmy86GJNYSspGV5tf4DnMIGwq0lNsSNoJpbhyDnZ74bSxXH
Wn3HCCY0L2MqJ9fvZvub9BDupfOjyHErq6tuwwGbovbDGxQWo6Jn0dgqhsxa+N7P
EDChsi3xt2SflP6/XFnDskJpyGYoZo9Ao96VhojNqkclC0hql0krmZi9O0ljVrsC
BONzv/sOccHiCmiVfYdyYm7+0JHn2QjkmDWLI5mZaqWcmFS5DYjpERDEhu7R1Tic
qcY0Xc1natKE2Tu3HGcpmFbbeOAgIrI0+cDdEQAGObe9da+vilHD4KE8gIt3xauf
41Blr78gvlJjUegBfTSJzP58qcdvbNQVzLRqpNp9i0eyAvGyn9oVTO0JuTJy/sLk
GgyDCK066bFE0f1eP4iXYkmYvGat5VwsJ3jsdpw3DvV5x4RS0AfTWrcPfLXgq0/o
41bmRn6vnIKXkat47SsHzJYSeu02/qyJIob/A6iQxnULDRlFOplp3ie7txelXChO
fd2qPuQGOanpwc8hfjZMktDpkQyAdLo8Q3UxLuVdYyjAe+zqvrQsJ7ghNWutrnne
PsIEXAe7PL/qQE/BxmwOirImOQgEIoixnZysLL3JqttGXTfznttcYi2vuBqpQIIy
vUYhS4JeICZwtYgWlIsPtMuZJMMnIGibBhwezuVk0x2TU9DcIPG1xhdQEuRXXggL
JNi8Mh98e2rAFUwe4qM3lm9ih+OI64V9iFlhn4ahFpthI7UI8/MVWSJMXvEV1lv7
n/kgQqbRb2hIC0MSGLoc2PI7aQ+anW32yKAMQNrBznl8sK4+nWFG/cfbN1svSwZk
ag3FGksK1SDD8Me6PulqzptvJn9pLiy2r7OYLp6xPOUAzv+sTB+jf9OdlRMhJzsl
kuzRHQdItBqV9+qbd15TMYHRltqbBmbQtpnMR6Jp2gN3MC+duhq2YkxrxXJNthym
jm8z2UCf03QL0wGnhdJgmeJEuMO5tEQbrmOxnfTPHm4M/6TTjlehV5RHdmOCYhf2
DkWMLjCSs7D5Das6KzcfyFIV8kSm3CTrjYXV57F6JDECUH56KStaM4loCBuPT3YA
sVIY5UEDN0aHQBK8gVXbmhr3rTjRoZy1UKCKhAPdNnVvEf0Kt43pPHD8wH8xn6oc
90MTSVU+GU63ySy+KIu10RsiMq3I/RDggCHFF9XVjNyOxF03+x/7jWVngfSF4i19
hyTRQuAu6R9BDSONe4SoJSD+TO6fzSPgIzpJupuTKaVvgAW/cOKJBtoA9vfzRk00
YdnF+Z3ISlICr1odahhYvpR8y6jLiR2ojBmdFrMZ/OJEedLLLsfttoPPkunqqxY3
vXhS0vN2s7kSE+43LwEEhOdFbMFqzeYWRYX1F0iTtAC+K5FyROvDTdyufjqv9VKb
14EXe57C10gI5MHkAhjw8oRTIYUy+UteU5GSv3eHbts8L7bookqTw+n5rShbUzcF
fHFrTbR6TEBTkzgF/dF0QQzC+/bPIezIDsyCi0OXgrrxyH2uABB92IwbQagFOpFD
xemeM+jAB2u/CjdGw4YiW47n4cDfwyk/f8iwcyAyon3t3gW6biNZsQW1js80KVNX
d9KDumv0CC+XZRsqnOEJnaKRSi6HLv0gCYq7GIQZw1EHysxamqGhBh5fVT/bn7M4
KvDshCfxlw5pnMjzG4yvDC7MkXmvOKme7nCBvwthYSamKoYdt304sRAxBQJrAmuj
SdgfaBnTmsFBwmooCESKwhUPaFrrqAe5zCMzBoB3Vxy3PHyWX/SBGRtAVZuk2QBK
kr/ekIVL9gPOtoprSV1yIwX8Ge+0bxT2zaCjoxob1bPRzuwkmxrzmRt4ZYoDyJ2B
IEuZMdmmnxOjShTHmWw9VOAnvev0LvlXMipB/Lbdr1PjM8BCltC287O07By8YeZD
euSKzJlab9oxiYYmJmkUFQkkiWk3HS0okWN4fTMgnxzmwyQuXBt74TtMQBVvfUlZ
xqv9iP+VMDPsCVk5jMMPWjT3naJThI6Km/4x2+NbuGmTQKS9Qznqg8XF26DvI2/F
vMVoOrdiLbNw0hIuDxiNF0hd1BX3qvh25A+lGIfUZ3c7jqlfO+Sou+phcpysRs/U
2kGG66LfLYChP9zs0Ht98MdtLo3/wC2bQClyqVVkTuBcBYRzOM4RK2gsDG7Vi9zp
nNjwYxMhyt5CNbZxiqnfKjgch54s1Luzl3f3g7vpTW48C26tnK/0Vguqc0zFHmf6
6tga8uPRZNea6E+uYZkGNl5PFz0aEVLjUfrBVWbO4GzsbGQqvQgbBbHfx7t8PwkW
i1OpTOtn+EVtRAzBKzITWaIMGgluVbaKULnQZbMEbXREYUU+4lyDPY1vKIJmHBvf
r+r3LCWXEJfql99dq9MNLq7LPm8HQHrj+YX5QBobkV6diXdpg0Xa4c+xnFkCFTuC
oTg1F7K6PlwfwZ5t/K7WCemBFYnZvJ2A5+zeL5MOisPWkDdPQZROW2+BEakLmHGM
g3RZy/roZ2iau3AgcqRQ+cbZzydZZw/VKcndZW58drhKsrRXB7YgOUkcK9GRXStb
lbEQYa1m/13lmh7gj7syzG1UI/BcFGAmognvW1zf9VSu6IXJdMjpNBmOfDdPqsrT
JaZ4qxqcc/KaPUaRiYi/VaDmum7gJtrW9/JCeYEKBWIi+wRow1SpOj8ARVLE7Gbg
5q+8GX73bvvJmYxyFWAAsSS1f+h0xXT9oaYzB9QoOJ5fgicBdJlYDsnrlDou+PUH
aHFtcoxl1/V8t7xJhBimkuXCwKGH1XmErYyW1aP/azOEiOxB/YVV0CUz5PhxqQd9
sznNaCMS7ZTR/pbN5sM1Y54mDFt8MHYUzyB953SX7xQmibz7RnATJPK5Xn79AllK
u32jykMlOtsk6uQCEs1ATZ+u8D7jpn00Of6OGqcHp3l47M4daWURWNNH94rGf2ss
ilORArmunClBdKNYTppEoWctPZyGKrVETW+GB7XmEcSOSZL2vweOs+DGCkqqL2Og
vi5yEUtEt3ub4j5zQpdwyQ5qIxwfdj+m0pMeI8/c6WAlj+GxHCIhgBs/ikp7OIIz
kysYEcYog1vlKzwi8gLR6IpRj5LVbccNzraYu1uNNbz9HUvFbyMpy2shC1EF43gv
6cQ1eyAF/Kf1BWhTZpGIJWGjtoZGtXdwH4xugHwd6rb46TsaHEYkdHP6wlGto8oM
L7Sc3l0F+amsMqni8yKRoJjGTLj655UtynsTxEhd072Wem9ja9TXw8HEVilDX59a
hMN1RLFiEfsfV4ixFeprrqRowVRMO641rfY52g5Q3AMdfAx8DNSDk1BXNa9KWvY2
+25kqfQk8bcRI0+8EeFQLwCxoRp00XklxAee+Hkqu67whm8upV93hLXm5RIe1wta
Nk1ZfqVhepQFNHIQrmPWWyAg/zcFIlvMFKtuFo0iZkIYq5TOyuJzDtLwOkQ+OdzY
nA/53XNuzR6cN4II+FqJmCz0Qarr/TrWThExn8F0R/EolO1+HRNNuDHfMZ26JZJr
jKFxzHqujdS7FjTiL/nApqn18vgG9yq8AReacnGUdL+ZrEo8oL2ZPrk0MWujuJEA
R8z8CrPP9OPIqSxsbD+GtZhkeIj0JyBlc/dFfVARLwpdTUYIq+VdLtw6KFZL+C6G
2k9XS1cnIaCNrKZMnCY179X9KhnJDd/YedVI8t4uN/zjyXCRP4DpqYLklRPvCFzx
8DhuoSPkSWxv3P9vhObjh8CZZsxmhfvus7S0gjiMPdmE/+p0NUrUkuY6x/MhrkEc
crrpborNnprtDn8X5zYIX15K6QX+gZEyfzKwiyt2hL2RtnufrneaUXbffRYeLxMs
s6CW9I8YnbMkT8LCb65OYeMfg2SU7dfpEwNac2Jr6XEXnxKS0MeXTdvr8pUEJIe5
ly49TBmS/dC8FKbob+P9mmxbS2KskHZxX++myfNPLZZUngeWAW8pT5FiNmKzg5xb
xDTnqka0yNazCWlGDxleRoryuDFV5QwTxgMsQfMspUGTx43mxLDw+z0MmTaAyG5y
lWFzrdDzJ84rzU06JJJfQxqzdhT9LKGqRM+Jk31fx0sJTVrnhJ+ayZJvczLVTb6W
wP3HlLFX4Zy6+fIq0FbDT2N50hDLeeLkZBBTxmvI6Q4NUpgS4FvBy/P/xdDpaWZS
w0Wb7Qc57W9Lk56RyQxAT1zwGiYV2HbUnFntGVkjcoxhrd1Z/CxeFR1jRaj7SqGa
jYR/T5mpuCc0YJGIPERrodw7IAZ5bdfObBcwYPANdgAErzBraTBDMfYT6M3JuuXt
Oe/ukfzb+/cdazGPNV5HzuOH4osBA1LnAos4anh4O3GPSm3dPOSal46CS8QzLa19
+5YNkxRS+UliPX9r00FpSkmrp0qYIw5fih6LFwjFLerDD8298igEQ+zWhnI0wDm8
lkuMua+iZ9KnBvws6FDHwLhfmhw3DVNja4fBhQQvp/UvOtYDJmuPVoLL/dVK6R2L
fSoEk0t9LQvWWvhC+cTARSg4xId/Tr5btPO7aN7zbHTQ4FqOBMJ0VyMSSRo721fJ
fFjg9HVV6viDJV1w1HqcEhDNcydEs24OUtPzw8yR2O3OHmkNwqP/+rPOz6W1rr1/
f2QJkIOBbgZAoJCCfWEFd7R/S2WuB5TBtzx/qwRD71ofvHiL8nio+Sc1Q23MGaW+
Ws94U1OvDrBtKe5QGVk15NRVrdjN+Qs7RTRa3WzF6qrFtzPFIi5AXJEjVKKzHZLp
vGIapEXt/1eB6jQIkyugS04RMLAIV0zw3ExhvE/AdFWyfwx0hX+JyfHu0kVdXBkN
oYtAB9FKezoxvGLO8toBdPieGA5NPPer4OyxMg3zBtb2t3VaYzLsWDXBMRUUis+R
qiPKR2DUxJXZNETVoAXAXADNhS7KHcCaBMNh4ppuwK3u6y5cGxJ1PrZ8Ou9geEZj
Zkumr6DFa24CptREv44nR+O9CZIJbOpnfz4PQvdBmXZrTk5mymiofXw1bS5KFyxd
kYT3BPcDVid3LesGrC5yxncKGlLp4lquzM+FaH+OpexaRHm3vCbXNGui7/nBLEpX
f6FLc1SZvE9+Au0JwwV1KPaKMgtdr5l42NJnc9qqeZRZoR9UR5hQ+cXY0Yovtp1C
nF/kkeyWWZ9pfclDcs1IOYBe1HClcJLCp8fZfvW2MJGoXwS43cHMU/zxe5VfNiPf
HL/2E4WJ3D93UDp1uWwAptTKZ8N7b9SMF4fH5+30JIp6T8pyP1ldsQeoYPG16EF+
lmlV6Y+ZLNodD4WUb9x2pQQI/3g+2UTPT4pg0C6HfwZvnaQks26OilStVl7ug3P5
dECWIAcwBcSTlpWo8835lY5/1GAlxhu8TtaXyXtw4nrIBkItl3GUsLKuy0Yc2RHo
4KogxOyxR5e0DJxk85FGXr6RgiHoc7wy84AJUYn841K6byF7PuqPAZe9+HQmbvFu
YpRY1O6thRqmhSDZcbDykL9REP+E+InPLP5lFWPHl72XNbfJSFoWnOnmdmRdw+h2
LytOi5ijBZEC8Pid4usU2qzOrAEqvbGqBDW9wCA4AOPVI2PvzXAuSUflXuvn6rJN
6keTIYO6GaN8jAKXfwz0X4lVzz/vS7rm9/pSfZwKdWgyWrZj3bsX+din1MeH32qR
2IcZKZJ3ya85rFNX8SwB1zeRKKa9DJOyeWFHpU9CC+Mmx5PGDjCSIusPUS8bfB5Y
I8nLCQjf4dw0w1y42YH5UHPswKwj82zL0JggOAC7F9YE/YVS7HUwprtf7bs3ojWT
F3tkHmGyPb4/xDYPFn3ibYGxd9UhXJqv4TTvbVtdoKbuJihETo8Pr1wZGL+M6qeg
10paBtn+CeSVROiGh5+CtsLNG7pSJw9On/rncKPfRZnsjmY1ouqM3BUfYws7iKHq
pyWkvVcoLdXFYu1T4KfqpEO98KIefChgO/eZD/FPCRBKehSRNiJjtFZQ+ax+yzbl
Zpy8eVVSjaG4f/SMrObN17tH7Wi3tsCBhdmaNvtbGzViWJSjfngO5ntH+CwqhD0t
eKUBCmUr9IBnBgGeMcWz8TOgh3n62wmkoxgTAM3zXkQesaccsythrWhZDkpclbeq
pp4RudnAAJQ+t/shyK+/AlgM/PATT/5OcUvE2XreeyPZkdAD5cs5e4bBHEvq5jeB
eQjB7OSFrUDXeCEsAdPFQn7n3qaI7Tfcw4xHnonZBNcUHzrIA7lStzEKwXhrcxpa
R9R4ZaUGC+gizyxk+Av3kGPHuR78nq/He+kyNTO4i4nDYiuY4yuI9pV/3/Z6nmJh
7vB2ByHc/c2Bxkc1yhIX6n+7tRpnqydSF1bUOp8sc2P++pIViHjZN6oppltUoU8L
i3FmfzwcyENxFwwpQ0AW5GDnNzeDEquDgZtabVJzwHEhbOchvV2RjGf5APUhrWsn
B+NIG1dD1T1P2mMHC9AFp6TvZbMcuF4fl/TlJ3fzjUipMhCVNLTcoX2zUY1j0va/
9ftEd3ZPjhLelnr1BYFP5+aw5QnDTeXTTAKf7hU910VHDpMuZuzKMEpNpL+133It
r0b+weBxFrsyi23E03GcXSHNim0erYPFTBeVGcDFsAqZ8dGvRmEw5FJ2p+D8saJ+
Emqz7a7DH9VvhB1qdEYDBppGDwkGcnWLEnkwPE1n8l/ppt+fr1sXdQoFnVJuKLcg
hb3ehqUB0mqZzoFd0V9C4JKRWrCDOEgiagNovmE30M70llfmfcbxOl0BT0lk+MJm
sfLeYJM2RzNLFesICYhxR3fvA44UZU3JFP+DlSTXAKuD8j5/bddiVXRLh1vN81zs
QNzEC8i5RYoBO/UAMkMezywv4ew2pV1p4Ss8CB2z2v3iZ+h1SsUge4jZb4oL2PdX
ivBPmvYjXXXuJA3odbiERnYuQQnm9woViUqUDMtn2iR9VwjD2eIymQy9/bnJctwC
sQItChinYRs0xXtr+6aIjtIfTJjHqGqnWFWI+5T1hLYFi3hvwADLKfbYxFV+zEb6
5+50e4IglO9mQePdCgUznSV8B/1xK6qzXcQqXoDn6PwTCW7ZaGb4MktwtVGcdiPm
+l6IHfnJtT2D4Jx6dkNHZBuZbEEH4CUkkFMXtdAwIa4eNB1WtAdSLX019ld0Y/G6
bR0ecxzVlm0MbxhRaN4v87JLiXLOTF9owdmK2asJBnKiKrjVc8UhpaEu5g+pD7tp
+nEGdN3FIWQpmAPJTj8TGcP/+adGIsDCvaZNuAKn4jXNjao1HyL54rVArYi+RaPN
UJ7ZMFi4SUuZLF5mJ4zgUqWM5sV54wwKJLXLES0owY7qo0nfYO1gRX/Dj/cbzr0g
cyagK1/L3xOpcdIpXslnR5epjkXLBzMiefpnyAlm4QcsDqAurldtwafhK9mvl7hp
zn2jjaoSJc12IdE9kQWkjT2E3OuL9vKWCTRO7CTyQPDBg3t/7vxn4n26eBJioh8u
7Xa1aZEOxNQ3cLxxtCOUCMGVvwGqNjd3iNHQTmFuysUDrK08d7whqrF6yXY2C1d9
InFX3cyUf7pFWiWKm9G3NpPIaFjt5Z6kCofc7ia4BAzWHcBwrxjKWewsLT39/cUG
tqPIGhx/WOPnSfk+Nlpkbu8L8eDfFzqda+CJvhpfxMufmkym9HOaOnGPoncN3+7Z
yF6j2FdzEemnCtjNcZ9TJBWEXRA1u84lxzWf414MjKURqep9T7kVhnsiBrWYnYAO
EUJjN9OWu/+eHq1z495l/0MPgJN12xvl26Q642juY3O7XsN7XNjRxr2C1iorhQKC
CAPcVrIsRaH2vGERiTqjLpRuvX4iSsxndTksjp4cjdwqH8cLq9iN4/so868smXTy
6G2ttxjAmTgbE0WhGEQ1zbZFM1R4KxFPahP0SgAmNAFfKFx2U8Seaa7WKQagxo/9
Sx7473AGasygNP5sSNpJJgfKuGRdZtANODOvpM1pEqlGPmscLGksuwf3ceon9fGC
2wmiGY7KkuOHq5t/3mZ46KFTlhneycXJfnolQW6UBuo2t2DuCA6SNU4DfqSdeAIx
HUfFiGhuqDFj3bFgGogrUqDilQZyGQho/e8KDrPO6zeM9HVgCvfYUGIs9N79hGda
kT4kZO+VdaRNfTcivDWU/dazm+J8lXX1pMI9dU7ohES1yFn9qBcNA+qpjsc3gQlS
NgBLW+kumLpjc55fxSD9QBOU4AOMMmKGzckNEJvrjeYEjJJOmpiMZNV+rNpdPN0w
/oh1a0CxveY7In45d9JLK6TVa0PjGjUQhNsBvrjreMZBV6itSODX0Ybul1KgxZem
duZgVhK1jt5s1zoXaO9nggy61WJCBEzxLZD3fm8l+fZz5FBwdzrBENOsWSn/k/Ak
/Qer/d8FhbV4d/zLlBGkXtK/yGUzwpBpUWOfDpdFzVL8p5WcyEWMqrIs3BF+l7m1
vEv4kbCXFNUU+QM9AqADFuBUMeN7OaDZnivh0C9+sbnlLkYIR1M2yd4Zru6JFRU1
Jv1znJLAI+aULr7or5kgrOr09xxcmclMkHDT9tr1trGo81YkaOBqoK9b55NW78LO
EE6O51djS8sg4L6u63DRYoVOVJgUAEvuJTum+PRI5V1P/cPIdctnfsWBP3vCPbej
kb9r8454hoqzONj4LolwD+4haDuER+YyVJjV1ZRSvcqq3oINv1Te0d4yfOR98TAD
43LyC8g6FnijZYH23kdeLwHWBPsDqY/voOM4poZo4EbPdvoEZy3yC63+j5EiITjc
xu09zy1r5kl+S4Du1dLo3I20sqyL0+m9qQyvH637t5+Cghl9PLfQ3nJZ5J1/qdRY
zKM+3IIrDkJzN5xj15J3oiCUZTA4R6CY7swLBEVkNyAu+Ks+T48QLEfkRE6MMPHq
N8wpaP8KKe/7drjhzPGJ3O7/2hOqH+8ByjeAtO4VW2vGJ7IzzCyK1Uv9PLIE28OB
XVasykY2aWFbgFnt7hDQjAOY9t4Ai29llAqYGjlr0TiMaYRvywZiNo+/GmT+agoN
O/bOPH3EMrcZBrU2weVeqCBkRMEKL6vlHpPFfpHe1SWSuPLLmQHY1xpYRSVx2MGt
uttS/E9QbiovAQoUjPriYFzx2bwk9RY4UKLFTk+HyrNYPfO98P6QN/uh+S3U8em+
GbjsYyG+ARJralE0Vy42ZC2gs7gL9iuipt40WotM+BjV91wi0qzFm6gz+p17lLFg
4F/0zAX/VwhXDE0eRauBHzz+rFyMvldyDovJXGMCsHX/tkuVeNsgC1+QVmVLrB/x
8nYxMt8CMC+MZYP5GDEen1sVqJltlbQ8GLvFuUlNWPsQWWu/gWXIzBNuMJI8zayc
pige/Ca37h/wTmuQKfBNzE8rYpNwuIwhgePBhGarMToxE46038FedG/0DyUsVoh0
vYbZn2EqSNEY6lvMbVxP84nMXo0nBgHuXfB8cBRiypKcteUKibrVXEnQHQcItkQ5
iMy/flZITakgupH16FQJOCO3o3H3LzP4lm1nhSuc1UzC4HU8S4UQOGzF92Fl8GOZ
XhoRyjAa5Y6QOSV5ChSnJY1Tu4pXdD4nrH985cqK9UwwBMJyuwvGo4+krozRGhZd
sX/5HVO8K7vEw+IvmKaORJ9K2/gg5kF1YOXe6VRpMrUnonSmlnuZLpfPqqFKUg09
qGL4sbxOGT04JG7MVCvMRbnWZX8ydMPFBJyag469BA4lAejR+/ZiOMUXMG50/PUg
vuYLNCEowj9nXhlljCjahB1jJApMFZF1pD04SqShH1HYP/pzdXKoIKGrduCW1FwB
tKiilN3WX48wPpKZa32Qak9AeCk4DTC7XDz5ANiLCF7N8Rz3ZtNvF/1qWYrj1My4
UiTw+DINdck5NervYCTN98hWlQDfmPaMQq4CTaBkpnM1m2K8YLigJ3BgicvylD6x
9GDJRyhWdqqptZohqXyZHbN9UjI3K/x1LlGpIbMN/GfE2iclE0puPz2RofmiUYGZ
1Wh6RrBSTJB6nzv5OplZf//rB46ywHpnwvNaWInGvjD/wsk8R2yqJJlLYe2UCiPQ
upYe4UWvGvhDPBqZ8N1mnTlPCg1FWTyowTOuNz4JELE0JwhfalhHLZsPL1HzpCz2
cagDP5tCwzh1qwAgyITpKFqpJGGgtgld6+biXQP/KntHKhkCKc+NjGcKCFOrhq/z
KdKOFAvelwT1kQYHP3S+jDa6FzS+VL6xhBNbWMtDy8yHEVb728UhT0RSv7o0mfib
NDKR5JTFRPTsi+15P51q4ya8Uz/IBKaaZMQQ0JEDRRDqw58uZTi4ZR7yW5w89K/V
oIkhufRjSwDoAXxn4EMA1k5z+6FgA88vloyUZDfG/xEYQDnHH6KoeNlBjLzP8t9q
Is7+DBGoCEi+qCdcGEoAR9F71RJKjCfzifqRAsMzwLNRHek4yQKbZm3nrg/qZTdT
DjMcv5EuKOdbAe+TGMVNdIjj6llB6PX26abXTv/0dhs/p2MqETn06mUW0h4uURld
22r/6GtMIKFjaNlhpw+flS7g3WUL8QkcLKjALLEBOnwlSgPcY7eS/NWN8O+qE+/D
FKeq6kUINaQPkBSz4J4Cjle5AqfEjjJqr8jMjyWicdXdvP1K7fjoMe6gXyOsSf4P
NU6ZaU/Etb8+dr4eh4BdjOFcBE1T4KXuJNvMrAqjUP9BYtX0+a5oHu/p+riQg/VL
WmrkVmDw4e0Go+QPJ2v5psVVRnDuObNnkI8277dBh6AESFNo0rWDRN+MHf1ZDjEf
uy5wlXLJgt29Kcmn4ZLKAK5t8N8/gQpDmGoKPnsivxuwSNYu1DYvMgYXgSTMpP5J
WiXxkEOb55oiaJLOEJfi0yKBfmHwEpw3+YZWwWqB2eZYJnYNJuRs24u+3eoIJrmq
MCQTljGdVasuIiyfj5zjxUwY6yTcP6w9NfTIoFYhe1TJ7xwZedeX9v1RgZWS96bc
cJ31AGzChpDzU6wjLpuMV5rINxcYRwSnrkF0XDT/3qJSqdfJRuYJqnl//iZUTzuN
Ea/FU9tz8ddUpco/JpkyPwRfPJCwXx+rbLCN84clBhtpt0ikuNIyxvNPSKkkqTPN
Uxu7ecclnPZsYTRUjeirR0KOHqdZ+YD7aFnQiXde7y3dg0/YhKuKMlT4GVOuRdGO
D3IO0I4JB3DpRBLmONyDUwthJemk9iqyiB7BpdMY8D7KFdfDDuUG6P+QXANb+yGY
ArjIMP8kIcsi2BN2ZgMlXKfxRVOcLMGohmarnBF1L6/8Ft9szSTjf1E4GSiEPqIm
Jb5/fVACdjDy8UHujlP5R2C7M9ML+ORNT34jYUZXY3h0kRUdrIlpCcdnZX0b9FNI
KrfQtxgiIzZQPu7h08rNYRRwasf6jNx08z58KhEr39O8cBWmq7bMgPATXCX3CuuF
CHWS0Ohne+utjQxYhcBuYqVmJOsN86jmoor/zhO2LIR30hRmHoGhXAGObVioft1z
nM6sRd6asqXxLlk6KTakg49TKaKJUCR/ZqWKgN56UokjWB7ZmRZyXwlCAETvFtKB
MXhEKW4xkXaIKGuV3OG0cdpg2SCjr2FMW4dAR3JnZxb67ndPxlczRQQHSHgKmOMJ
zJUO6zi/lNEKVDk/uXVFQELXf6r149Y6hX3XGrxfpYH1XnsOQ+HGPrTQ5J5hfFZv
BXxaWMLooD7HguV8wfctt+EiGnV3YOt4Bswb5hoq2Bm0/4OKtA/3Tnd1jBnZMBkg
bN5dWJImfSqYdbrZr2sFAcSGpnTLVSaxR5SS0Mfq5IuXwStmyIdiy/s+uwisA3BG
5XwbjcALrBV/NgDAKLKasgNob+e6q+MZiW3jtfoyeHwE22RDIiTlImnIoCjD1MMz
uGNfmtL925eaN5kYPJHv0Z8m/1iT0Wu8/5wwHVP4mnKkSLY+zk2EanF5Eh4J8SpN
40fGRWNJf82hhm5MztPUjxRKMx3BGAIt+JdG1JSEguW4hnWHYZ3qZMXUsKr8fpuu
zYcZw3ZPq9iYHcagqOLLbKswZxV9cJEDI1oFKSh+DiiBsO/pun6qZzDfGxrmRJHE
GP/r8+lVz9Psk6w00zgMK3TFdu+OemadSr8/5NzOJ+13QkoKzShSiK0+cJnXTgKA
oiq7fCqEpsAEjVOFrAfOhaX7zPyF8bdYMl0CneIwHAH0+fcUjSsUX9ty2n+M4d28
c81KZ9rQEcNBZAuSFSq+kjW4PLdTMGF6MBEqau49wscaDVJK1MG6xU/Ge4OSgDQO
Jhz3+Gd7WVeWfAsO3O8/ZzJhRGfsKRmCMf/rYxR8uczq1hDHVwQ2Xs2t67U1G6lb
RDzGJGIMm9+tBGv+E5zeuGdstvMh9NwIQbZX/0UoesM5S1I6/G45X916SnvCnU/g
u2lj7m2mfw5Xhtfhuw4XL1WF1YHm7+DMGr0NnY+sbLMwqSzYhRS4jkHk6GwoCpVc
sMKbfyUmAKDPsnuhyASaVcAVaa67QaRZQjOjEkBFBRW6sgdkcDe7g6fqJ206anE8
fhi5b5H/DNf6RUCGVj9LJMg1HbaxQn6G6IfcAG4EgYI55jwa/0dm2umGnzPMNvzH
T9Ze9LRIVBYlLYFldFam2IMwIltr6/hS+g93e1q2d+xWplrGD8Tw4t7Jv49Y5oWq
qmqpevjsxAxV6D854Xx9bXed9cVrNcJMIC89uD0THas4EV5/M2a6wCvxnyEw66n+
GBcu1XIIJRxdXd/cvb4+adoeI+Ot2i0hCjxHGQuKFSa/ftja511J6HYyayshWRIp
gZzPxEQf70wWQXrkJETA0ChySyjb3/Ev9u8pnguyWgQ6/fWYAa0UQ604d6Wx4G7i
GdvBsWqZaenelcyArLece2WMdV0YoKj+VRjwIEmApz8DlPEvlyYzt6YUaxWXqfCe
VRsRH+266n7kTqr8rFthEskvYSARmmqj/HnOlLCI7qIfzBNmb5EZLmSiKYnAgYJd
TX5wG0CBFGaEQFh+tnYMKu36HOqOkn9N61Vm38X44X7OXU8QfeS3ld2ct9YG2fLL
Q4WsPgxIDXmDhu6V2mcsKvn9ubJ1ji7prlYvioa/PJ1a9GOfbKhZuUjoROaJpoaq
SyQoG0hFRm2Y7DapuN5Az0qryHvBkow2nmg1YjbDeUib5+Kzq7z0IEcSwF9wx2sA
5+osXQZMAzKxRQ8YghmR6yDfoDQgN80qSiDfPO23rlBoEwOEJFUn0sh0srs8vnMl
NSLV1+x7z0uAfhr8bXt9ZmEMK2CMpuSrB9Q2Gxho9Utqku3N0kUUMOcm0ZOYD9GI
r7S+zI1gQs+HbTOqU/cBAdQ8idMeej9qWF8ZFGQqmA4qU5qkmDpSYldZvrlzqE91
bjnz0bf7Y6Gm0ObzuxvA436SbrTGaEFD8opBskNwjz3bBdQbbHODLsRTFiq/LDg0
O7DWiVcN0prqlYt8UQzu9u5fJZXulCOPQ7HlLR9E0o9ZSdoP5MV10V/L4Mv2Q8Zk
gfciDwjZHkxcIQ6cInnFMsOtcdHMVs/mGV3rV7Of4WnecS4fC/kBhh5m62QMkXsq
CJS2LgwWEYqF/aPhz6OmLb5zbXIrCpELs+WL1SQ21vr6sVUhdIUnKRWp2TPkU8Xo
LGTXo/blwaV9IO6YANAwC8qfSVY96CSa2X1oQrXbSSwzxepXJebh1hq/vMbymA7/
WuEQMWy63nZDKNx4Wfe+eQt+b9M101Dabn3I9fEAOSdJj+eZxadyPv9NVn9K5A2a
tcNMYg9qyjK58p2wfEk3rRy+M88YW4xJATjSy3ECvKnry6PxFMSyPmnsbGJCUKx/
1/0RQY98jtZ72oLg8z1EZbYsAgqg7ycO7tyXGbTsxHqncl+IDDjCTsO90e4erc3U
P2PZJ/Bcek58VFm2qZWvTBmm9EdBxv+t+l4oCw5FVUvZ90wplVVG12KR9eHm0hhX
MH+qHcoon76xLL7jyTZx7R1Jx/LJOeMbjVNDg6VyP2rq76yISa96lPgLNpWfEAxS
h+jHjUAdzesb1DRn7lidvx4GVGaRMmVlyX4D9bJXjjNtc1XhQEbLsESFpRVRjqF4
VVs6zS0M5mp7nCBrSLBf+uSixdG6oXv+AxJOxTGk2+FbQLjQ2HafT4kLvbz+Zktn
RnEnaf5OvONgHgUyA5oDNvHThLj/Hmk7AChiGnJzhqJagl9ue7BchA7BPcU/qHQ/
G1TmhRY/LrhPgeS9PIjqF5aUHRHgXpQwmXl+DfVEpsrlvOy62i5zu4n9mJhipXks
min5wV2AjAPf/N1Qo4NLYBSWZBbYD3vnBoJQUpepp5epK0rHxtMuyqhlY+t4Iowc
UpMqLVWMtaVJaoR4mAhKEb4QSRJnXmr/iieZqxcv0aS0G4Ray/wbxB6UljgIWw29
yWIAMga5x6z1mvRA6YGCeYrxue52IWFFgPrF7whu1fVl/mjMBrPo1kbU7OvrDpuB
WgfronTiM3mjolRlibjoDgb3zy43ovEvfj2M8kyBSp1BwlsL1g9WZwpr/lc42t3E
IzFvDzv0+Z4oaJoJu4UX1PqDPoTtH++0rYZwkeABSD6plS0o8WGbfmn0E6YfRXOt
IojXHdBbZtSDA2e1d236QI0BRe6i036YJDOxKw6SqGLvX+Uc/SCPccq3Ukljcp0l
96Bt139HoxzyqgvR8WnoR/87LxL44W+l11/2OXrbQ09ylZOsfIEMsrHcLssrm5/g
C2HA4nzADfrTtu6e6LFH2XLi7vud1ev/B0HWDpkIttMtApCAsmF3GG64eMR6pdhf
GFuEwswH8EyEU5anfd5FbFDSsfpwekfoLn1rzYaAkyNdjFqcNKu6z7V3ok0Hr3Vp
fcFhQ5sb2vycfnVkO+FGOLMZW4+7S0+7cLk7Ib1XGJLg9xdNdZ7Iv4CRYW1ws8mz
jTCXu2xxnR407ZU2YLaYTl3P1yDp6xu4S+xHLq7LAOe17YPz0/7zuM5zYZRZFTcV
QQR6Ob+sDTS6FJgk/JnawkZdbDC7pv+gYDlmNDxhMJOKMTvKiZwKSKAcADkFbHY0
EN6Dh1GlIVI/2QbF2L/l42RJ74iIg7TUWRO9FquKAJjH6cHYAr9hqP5vcxSOq0C/
A/AX6ll+dMHp5SjdXZLMLL8G5wo+6/SpOqwUTDxZdkSUb9G7yR0gCz3nOAg9DgAF
JBED6OGyU3nMA1JljHqn4KMh2hL3fJeOrPIY1tjYyoTFzSoxFNbzupDAisk4dL8t
kcn0/yyH2VhJo/ZCdjs2104U9Vj0ffcjLtC/RQNRWMXV4ExTecqIiPHH+pI/hEL6
gd+tlj1jG6y/sv/RijsHQoyt82PlkoZXSb9npNObT1TkYs70L4K83WXxkXogpFxD
UYjAUVlbqVTBg7NAh7fh9c3Iq10npjmQySBFnYURlqpsc0A/2gnUzju45qXT2eLK
Go0ZfZx7ZFtCxw4sk8YLt4xIDvvNcLuV0vp3gAozxNrl1SvdnbS9Z0WUO4T3dYCf
Dd3MOdue+4xyqQvcyHyoVYmrrZ1aPeE9sFpwowXEbay3UfUrmd2covjW7TticnOj
pZrHKeOP6ez24FUcc/helwprnTioWV/UAUm2rd1yZtlF9H1LeD4yBqEwRwO5LLMf
3g6rBqoRNZY4VvmYglSZQO1GSLAeb/tsKXe1PkebDJreFfygukQGbf4UPU6Ur8nm
KR8lj3Qsin6yyyolcf+TUPewXAOH7yHHWPPHCw/YbjlG2AxTpN2sT9rvYJXgNAGL
4jlqz5i27JLWzpqNII6buLPu02Hv10Fc+ZAI4CSNhjOlpleVWSEuCS5s1DEO6CMJ
ybxykFMQStOlBboXapx0ysKCOO5Ep6WCwWFruGtNlpnThUVECpms095BKiq7YoEB
dz5b8OfqPYe4VsNc+5+1ytx2b47/RA4SCTCfFWYRZyQP6arMxxWyLf0qI2zwax57
t1sDK8Au6mXxT9OJMXMmEx8Hrz8syWa1TnOkKWZ2NfIFHBD5HiKXPoVaJELyOc+6
LPwvideSyhBn+CU397NxHPSYWJTw/j7jZji89314QlkfXLvW/Gs+ttweMztRp5om
WnttO9/alRWYH9A/zWYHT+OEran5HcVxCQORiAp6yWFln9WUuICBOm00C4MmLSFt
nWFhnhipzvkMD4bf5adk1g7UTsi4P4f6FP12edRHZqkKSNlEes5HSpobNpIjz5zQ
q6pQ8/PUuT4RENFhAjwlQQXm4os4GfZVBSSXWZak6xZw8UJgb2VNaXXwMCkZxJU0
3bCkCZOPv76cmdSITjOovqnZ8k7GljN/itQBFsUtYphSuBg0E1rRdDK7ViZ+hTcI
TUWd6V5IxazUHEeNc+Z2Zvz8zRwomrH37n8MKlzPiJtO9pavsyckvvivzsq9y4ie
TLKT5kJqNv4ZfW+fSYjkm95JWvS2ZEDFz5VjOa7WgISyDaLvg8FQctZxF80r4Ixj
qBfu9EWBrj1zlt+UoDGGcBHnHvPDfDoa2LBefkKmkZNupCnC/wvUHLYhciElLJa4
f0lKd+mPSOR7YbehQ61UMeHza4LzcuvC5BCdGe3LpiVQD5Boug+gGsCbALqij9nq
+5cOGqWsCMVaYmSyW9YSKWnYt6y53Qdi772vA+WN2rI6yW3Jtx8ntCTHH5TSVFgp
9yC7y7evw0EF2PnKrkV7/YA1vS2zhRzFyUVO6OnBEiEXdIrWW34G01QrcdI94l5A
uR5vIwh8Xg9O0hXfVtvaasIjO20wOxpfmp5AlhZRnIlvS/7LRnzzk2nVASJJMQJh
ddFIoc8BL0npOnVVE1J7vRxmubnC29RH94ZOcoorM5+wuVlNz1lsYP1qvgEVYIwe
tC/nWRIaYFFkGFfyNxlpu440NNdwlD0cKTPhYyd/5EVMlvJ6SdzepzG3GjuSoxTv
Y4rDTy0IkpCckNDCc5JUTX2kQqVG1WO/unC4sk5J5GUAKN4XSDbTFjnW6wEZgXiz
FkVJS+Bod68yJVLRa/xPU6CzS/4lrLGa6C/iIB4kVlcXqZapYKthtiQ4Mo7/FtJx
4bAURCvmUv5EIhlfRMcJJbXUeMwUu5IWIyxJCoGSfoS/5DvzQ3ot4/Ej3pwnShY+
jjfEbl6yBUzo7Xx1LtJKM0wfAsbBuIt19OJi2KqEvuSa/xtg+jwEFJYjIuj6cQ5u
xlWfd2rLk7vkDZEk06qgror8F2XF4lq9Ksf2ScinMMYyY+Dyq+IgrcCCdKW9+4Cq
4rcvQ7XUnCxFfnudUSXAyUsY78wKAFqUmpgcFEVwly9dJ9ft/w/iVPC+f48PYrIa
2QKtsHLys9hBkB87EB2ZBKGVdSSgwKB+xFHzXD4UntIVYDj7cRIZsUxLpxVw6Sez
Gzc7gmqrnv+nY4YTdfmqETJBiALqSyTroD/9LhSv702xlLBjymdMnQsG0zMO2SIC
48CmleDsEwQh0Xx2YNCnyoLOOr1n0rmVn8SuAJR2AP0F8ZosHSDCUfiDRY4tvNMS
u3o+00KZtAefdRk55LgBQKpnSaB1tNCeb6dYfgI+L2DrzOdyLVWzYR6eyOvG/Pbh
XsY1V7kWW+9oG0EJIh1EXQ9PaZrVH/qGpTAM+rXZCi30GzgJA+f0J2sOqLbfzHqb
mDJxAsQjWgobrASLYU4BwMqMV4xAmFJ9l8Ok8ebKaHP8GusOaYOxLIJv3I5d5MUt
mREUYbcJlbV8180XeV9ezfx1SFJ3a55jT4bNquUrnoCRfEd8fkuUBuJ/m8w25mWB
Ys5H1QoGw8WxBe6MapRMs1hj2Ng8ulnQUMI4fYTfnzmrMvKxFbEArqATVAUojQrF
zlM8ckHG7eGEeOvFWJMXafdOe7PA7isZX5Pxf77yRRntlA6yjzHgBVnf3vTS0fko
hOwfsQlx9omozYStIrc18qtYGFGl++7WMOL2QxTr7eDwQ8yO6o3punifZ1doJlwU
sTUSRd/gg0me/hnQA6jDOAuhyRKc1P4/XqoN9qBTYj3jMiKKnPqkpswRIodaPa0t
yIhe7qvBjYrvW5PbFCAJ3GF/9bUcdJpc9xk+aWunQvknfVxKWjx995GhUC43+wG1
nVyNq/sePcKi4bhQ2I/nxP0hkJ1Rnc/09MT/9N5zam5ylYGlBncnco84huWdGxNl
zrbunSmsYF+eBNyARmfM0rfs2Ic94YVgLv+Ukl21ut2fsC+H2rSwh6aRgb0ucg9/
tTYUimi0g0k6oJHCt43e7qO+wljYwnnEg7m1G3Us+JcKSt6vWAvzjMSzM1O4jsbr
6HOINfzO0HBsZ8fVjuIPB3faFtKo8SXQlZfdODe52Df9HOhhBT8gQMQgQ4KUqzBo
XFe+UKVFlvDLxXM1rDMQSB/1YHiwt6zI8J82KQMVuglRrHOBN2cwnJPX8A2CS6s1
Ryz9TIvppErnSM7u+oyypQna3Gcglg1dv869U0z10/30fkkhzxenVLdKNUn3QvVW
3vNvi35bLGHUyxBi6u7DXgeCohReq4gETMnrlX17ELBbiiWa3piDVXL92t3HO2ze
ZCjXOwvZhNoGrcxQx9Dj9pgUzhjvkZAzlBgSVFlEnkWFEdDpAhwESO8fvajqeFTm
/4i3DRljEMCoy9v8oH/YYmxh6J/wdvV3MNmGuZ5Q8TNpPNbiJkGlYBixb9RpOV7H
l+ez6jV5SvtY9m2w1lop5hK2zV8CQ/ho1r5FsQhisimmpWJ/Sem0eVQo+o1oT8xx
5GtNerw4gx57MPT2J141pd5Rx9YGuKa3vDxr7OAhswRZFM69o2Rvccn0Qo2YKArs
yfQnBvJGbXOkn+r8/36Zyctw72o75HnNnTJRucxdremu3pAzd8WNeYGlTo+74CkT
yYpCtLRs/iKP330VMNQhJefRdWB80qe0SnTkmf04vqBvQvQRjcBTXFfpN0zM380n
hc2u9ObcpK9an1FlPwm35m9aXk3e2uRD9B3oGNGBh3aaWiE6LEpB9sXA69xmaIC4
BhJ1J5XacLce6uitmbJ14LrnxCUYBbP+8ATiBvmAzupzvuPW/QL8IbndsZVHV5p/
czwai7ggSrEQLIInxV/EcSLIyWY0kA+Wy6KE5+bCb4XOmfbRji2Caqvj/xf7CtkI
lGduTOff1tXcvzzgggzz1FwltXFPascLVa+/lVpYn0ErQH72EEBAIoobRMpORe19
3l0PT7hQL1qEg+0WPbh9HV0Pr/zUqatU6mf6FZPewZbMkA17xV379WqCW92kgHOw
lDfydEmDncJSJ3BlxiHuZ/Be1GdWd24AMxHtBeKejL1MptHsEONkvXObiTapZPbe
wjNPvoPKQ2fnha6K6jyUs2AGkhO9cuCCVXYnawF1undhZjISuIriEpka6M5huq+T
e8/qWjCqIq/r9Va5JL05EtiXUmCg5jReqWfaaEBoIdmoWBF8/nkKcoe9x+M8/I1I
IZdWQFS56SbRWLYajRXyNXxrqT+CBDjsUIdhakNZFb3JKCkb4kbsP2FjpwaHWvqL
gEouQCW/ADFzf3AT7ILEHitnZQpKkol/101OGSApDJnzXZbatVV7rnHnXabhIfT0
B8L2uHajc/2ZrmscArmriNlVTU6LTdAHpf22KI+mQUgDlT3MM+qOBKTee49Fl8/m
lmGQ3lUMzsKR6r96NToY6QmZTt/DoUwtwKKASs1Km4fFjCuwyDIMxzK7vvdYIa94
o4+04qCbny65oTzAFJKKBy2jMAItBa4/QpZymCqR51uoyJcFhDyPap2x2IDKd0MH
abvI2BpOAyhTKecILMyK4ZdVBH0gWKUL6vTOJz29m5Hm6sLda9n4LnBbaji7fivQ
BtZMbxNSTvtr7BVGeWqYUdYzqYMTh4dDq517bIeWBjiGcxZKsWI6Ke+sketnx6RF
0oLDDKuhNasip0rkk/bWQ1mtMFsJFBSDtaCOPQhxdwMPxQXfOvgHzBnN3BeNG0WD
thPqwDw+9TlBSCJGeCdD9knkHZQ62pO/HKbkKdrDVC+xN4eA2mc8ir6s7Dc3W5AL
zWjMGflPnopf+nPUl+CeX8Q8Bt88PAdlMB7+MPM3mTNNK55bVuHK8jvFdpYjg3U1
5bOrXusu2u3lHHqdLqbThoVmfnpvqpoe+S7f8Vd6udZeMzfeHnQbXOLaCFAJMO1Y
Gcc3ttWuiEMEM2CHyve3BTLpfSqkt1DYntalVdTXmTFMAfw1ntaVehwhIGqbOHr1
UngsKcWzImfRmmqifHsNOpUdTRo5R5DzW1//ttW+qetw3pZ1+biZTneV/Hx5aeL2
OG9UXa+871f3sqZsJk1smuFgZj5UxiFyOAbp/daWNZF+ze3uEazfT2/OH9H/bI1t
gsAeg2E8C9Xb5MeD3zlDfUcEgxexmiI0UIuZocQY99WBceKChxb8uVJ6ejIsfAHg
XeaefT8PdHfBkak7Red5QXBDNcMbh99xyRErsNmsSct7glJ9xwkR/HJCyogJtFk6
DwUPmBiAvkwnweja5O9PZek3AHPZwQELrmRyjh3QBDb1OzUgNEoo29gY80izBcbC
tB2YSaYwkq1rhzyfCmUUMhMKKd3RUkwYt+6mylTSOUf00U8KxeKUMAITxTz5y9Rr
mfSbmUTSH+JjParnrQctwHhMPeNibYCJ4f7KvipDZKjROnjpJdnJ77N/WYe50nTh
cNce6gYKzMQVeBrVJztONFwb4+2dCOE5ssQuBLUPQe965W3+rrkYCGnoJxbYgsY2
l1xVSvsNmEesC2KNPQBHeIgh/Qir3qeDyx09cHoSjUmVjLUbf9yoah55xopas1tD
Owq3RZal3UXYNbIAqklaeck4Ku78YQjw/kvZ4auASn9GMPjEK6wefzViPGmIeKQH
gn6k9gVUxg0F+fhxb1EvTQbiVDgtIxMmkWxWBgP9d6gyxDhGn8IUJKoLYNxfNiTP
seKbFN+U1ElKiAUS3/DRrzzYLcvmD2lgEEM0SlyhWDTqE0yZSAN25JqH/37t+4ou
TQrdG1a4qtPCySx4Ra7NIa/PtjIXL7q5mqPVL+Cj8KakeU5P1O7gKR7ZGb7kKySE
P7R5dCs3fODJUb2mA13mtd9Z49o02i24Z2Y/AZSIdIH7dIs0n+ZEwDeTLys1u+CP
qwr9QiVtAzSB2O7aJSG3agXJ6XWirnYhPOYI08cAWN4yizbQwNYit6TOGQNtu9A+
GfaKZifOKjQrkhQmUlz/KEMGmpaxlsH4TADZBeNSRcYUFV6xOZSihtip8XxX5b1p
kGVt1ZGm/naMHokzT1p03M7jeEPnNZJGczAjVeqIo8WVem5LPSLUBy09oLdFk6vt
HwqcsrabAEhgO4oU2ZfPFV59U6hrl/dWCJE150MpmcX6OJ9ZBthOB0+hRvhDYl2b
emv9dODVxq55E4lueiin80cJidg49t1oZy/2KcAKwYO7oX0Ks/iAJNdAQ+EYDfCf
tlEQCqFxsCNFM0zfFmLIMdveXW0TDvKB5euQq5J4BcfIfqNfdnURWvHCoLFQusw1
01MDKb/edeQ8TMQh9iRot8UCxakaxqvYPS2Qk8Cb1WJxPRhycD4NfuGyIfnw7OHQ
FwYwaP5CfhlB7VVaANGWrx7jsCrykd89KOXpnvd4NC20oLu2gqEbEp9P0tWRnSXh
WjuMd9LgMgYp1+vg6dJQ4UlwBKT/+NBmCEGClFZd/rIsmUdTtkCsNK1112ra0bhs
O7vZAjX7cKsVBlsztnYzSzoEgZnJvcTe7walGdpbkweGl4cmLXR6AAg8Iu8o7fBr
raLJ2D2wQTwydBy9ymcC9d4m4xqBF3db4IZevMvFcatuWQBr//FUPuaiuc6d0JQA
SlmgjqfNJjl8NmRlpXksPNYYoZGP5AnsRDAUR7QMEuP98t5RE3js5qv4H+Z3OW0P
P/wK+b0nYOsBn8Z/PXdUiT1leqVY85+/ehq/k0px3XUaKXgEDQ3YpMJfvwnk+SyH
SQFjRVm7RcRYwIFG824oRMTv5U2YwOky3DGNn0luthdg7qXZe+9+R0e4cvnOc0qr
fxl+/aNpqFWqSYxHph3DLEsSBYnK4jOtbfe29j022xyHGY32Cxnap0TmqNRIiZBi
UEQNgaWs50TH1EWyRAwiWD7TSQsiSUmNpvlQNhsIe5U3kGWrI3LTV0Rdu6ETWSBE
K5u9g5B4Nz/2CpXxmyYQskewiZVNL1QMYPQdjo6McbBO6ZFjyPvhjqaEG2OW0xcd
eRGoiZ5mRPp5yu6OhBoLY+zDMI9QztprlrFT7X6rdd48uSJ1+WeEEWwHSSrRMdOm
AvnxUKlic5t41tRa5/Gk6ElEo7YR5/hE/3kCNzg+/Av0LHMxo7sr2SedxdbtgkTB
QB8O88PsuDlAgLPxiJxT4mOEZ3aGntnCxcBWimqAzBQiu0zwetVLFBlWhlpKAus8
GeE04pt26tZTJwHA/bv4KOPLf3kYr8mw5ga03m5IlizYNR710rXigTCBPDh9gY9r
f7eBnYLLxBv4suPvuDnZow6IXO6jxnCYaJg7Zw+S7UIn5uhRvhO/wynIimbSR2mv
QPOAL1wWj/Ca85cKHkjdfsrnMDp5cFUD3AHKxHdbiJyCSmibTmdz6VoNRrkk8bTj
84YMk8b049V1qzk8OTB+1gKgiZjbIRX8hQxUVIAt1jeCK73bjsNdzCUt7xLmTJeK
WB8cy9vTNBc9rFBRGCjfVud9QNazouRv92qqpmkr6O5xP9iN9+CaAAgwAI/D2VSu
+uIGHTSEOyOSZGrQ0Cyx1FD+UQO1xrA600R/Hn4uWkwNQ+mydkWuiuEi1BMfhlvd
uy632d9Ac3GtcRs1IepS1g4h7NRvp3vBC4TPKojhNmA4i3u0tCbMFpBSTkjczl/+
cp9AtNy/LMtKdvHdLtOI02JejTPdMmfS/J2u8W8FjuEJKbuZ6oNzA03yTMTYvVsB
5IRb9CUpAhlWWlRLuJH+osbLV/loqhOAQ7MtWA5R1N3m4Q+GZOQ2hbw+x495AUfU
d0zLkntgG7eTkdJ6rV1lFrkyPONd/Up+6q1VzhTusedOOXoL12C2D+Dmd2Z4dl3H
RiK7On5EX08IJ0QGTzU569FdgE5v49jZD33uKYY/WKcddcH+5U/snSLui06KPJN7
4UrGefiip85cDNCedEJxGk8zKwsidtYtwEMxZYxqBwJxB/cSw5mSZcmcFtjxfblv
S7/N7Dc8vVyDIdP1cQDk3Re41N2+lPLxZZZjpyJCbXYWi+bpd4OzBb/X+2IodH3l
8xydG3xMb6hYovCpdQH6jM1hMxj7XOgNzMEHIkBGs5DFXd5kUjEbnboVeU4sjbFk
6lFvpgCDzPzTZwUx9joqvogI74njgiBgv7RNfNOOXmAwTwrsd7dQ/9zb0vWjrmVA
9QopDYiI0qD3Afd+40X+gsjOc+3LeLdDoUpjTPJPMJn/pgCqEsnr1hBhfuK9bsJo
D+TsFwynOv1GdqJsBgOri81NrAMk29msAMSMyD0Ny7ERwqAGPOSsMqNKC+ZLwyVO
pj/d1I5akW6b5/MAUF1BB8/oCRZyX7P+O4Bt+kcqyxZxqz4qdtu5fmC6kCAqM4oR
yt/S0Lmza23HcG1LHZDOot8/7D7gNxjWp9Bft3hzlEoWfDv9DM877UfIOuwZ37Cc
k09IWRoeRl+PRd9QxquWXioRbuSVm2Qg3u5+ui83NF8kGqNoUYtDFJ+op8XHDM5i
7RgD9P2VPi3ZBDgPsYS/lBS+FY8vZq6aN7lP7PeECUpQRTsHVee0z3jqxvX1tDud
gr7xd2bw4kt4xJQUDnuP+339kkfW/Fisu4XxWY/P+5kRhdZ3L7Kf6hSi8TVd5CdE
/OEQGDL4XLx6F8zIUxPUNr4y7hUeBuxv1HPVR1otnqpOCh2CjA8pkYCNLwbFNw3j
LpXdCNSFllY6KsFGWFZHuL1LY/TjvvKJby6KE+NJZgyqiGXy4+mA87OVDQ1LAIxY
vTzIpiyFmJwsganN61eJKaLjK1gDsG/SXMOpliQOtrRQG6RXhQrwRfH67S4w6rs4
IoKzs6sfFbtJlGLcsK2svIE2ypoBV9UiS6w56AJkeUNK/MUqRBoZqimdDa1X/n9V
RzK6mAhvCMQKqC3Q7wos5xde4t0ScHkYCvotHcNSC9BNmcZ3He7lvwtiMVlN+8YC
Zr2Fwhj+0LvjrC7vTCPShhi4ZYDZDTYaHhII/fam2lCBwmqjOXQomLSjwt9TKHik
xadPlmJro4O3y16OEFj22wxyQjKfm0RzC643rPy4t2jfbPir6/T/q1LorNlCm8s8
nzxS8FewvOCqLLwHlDNasYDz4I5mdxEmlnk7Dsi9WR0nWYk9q7lyvV3jETWBHIy4
IaFQdTXbJtGfDQL5rBsBrq+oiFSKoYGw+uEICoFY3wmS39e7Aq8AKq6o088UIwyq
CRlyw1VYGtLbaE3KLbwd0uBmIZulJkbya/23FEuw4uRF/WiifLzHUcxgPQ6wLhgG
HRaCTjE+ZXnlOBXLSDQcroNHO3ro2bUuLXid0x1f3AMwnqLTcVWdtXeiOXnewg4m
9/X0ezftNo5g4poVPujJ0mvwFNTNOsKCVh3ztxpQsaoMK3z1MlOe7mNfyT+fUj9c
R8Orvd3c3z7UNqEogqGwp+tKdK2sVSadiEd9W4h+xvGLVw7qcOabsIb71X0IeG6j
kkRVqcd/FyFyrUWa5t/VOEqenRyLP3WyoIoHSibhazFjGVh7GjULoKZLiYlOASad
hKGPicVJxVYnkmbSruhZ0im6cHqhHZEwq9kO4Ollzfcd78S3vsY9uGU/h77cwKW3
/nTq7LmT3nNGx1dsQlsjnIKRtqK6dORJlzaguRXovWQtpCt7aF5lUNOXDdsdQD6y
oAUa+9I2w15b7SL0pDO+9UuU4UBX3ebIPrVfoGGK0LxwuFYO3Sv6n/+zraOWhPIw
PJt5n7Nd0xftp9zSItPJgBSkhLlMBfIVFGSJoMkko9YeNG6qT/slz0Js0IxzIRiI
k3hT+d+QapZWuDx/o2Lh/hs5q2hch7Hy5ObYF/OXVEXj8bAs9Cetv81vq/QDQBAE
D7XjstYb99TS8v90DSR5ngvhx+BlH1c9ywhamu9MnKG0NTyyeLRxC2dZSO4VrBly
KlTEsJb/FyINGgPhMjKvEHZe3V7sHmQ55uDdTmqIMFiLD+Zbevci/86bgc2JSacF
Jwdu3mb4Yr2bZ7lgKLURfhZwwzdhmWcgu0G2vQ9ANUF09NDaR+0JpY9mVZ3R1Lce
9lHFvouMh9XvmEOqvT4hzXFIfUlrAoOH5Jn0zDYuEeYIDgVZENKdm3uJHIfD3wKQ
5W8emPWrxHzy0uXIMBubpIVGz6zmjzUWUye14w9WXHzHka+9UrKO6G8BqdCLwChC
f6CrzjlbJjfF1eF7Niu3Lm4UqpxDazfs/HeilJ57+Fa33rXCe/UcJirZwQO2jZjd
pShBAxboIqewYgpufIigKy3sqmA1/smGg14MXKeMR+HP1HV5Y3S+BOH659nOwkKc
DDIY+c1HYa7DNoHBB7IDCq19gGvl+kfpNUdvT00hfKmR9Bxd4SOYClhSNUziPEep
2lxgZgWIzWi5T0krSter65k+G1TMvrybQJcIe2Acn6PcpsHSNXbtY0BKMmZAbqKv
bJTzl02oIsXvs3yz1U4xTlv2wSep3BLxUNHO/ltBBEuCKbmhwYI6EvS3DR1izwAq
BU8FpTXB6mmjMKYbGrd7u2iUjzw2B86SkgzJ3tvCSAucx4omY1EAWFHeRg5ct+k4
g0TyH0XUE3LShnCe/fE46MpcD/pTFGaVtQ8nMxRFO/QjTrlplerHcwSw5ktp1fM3
0sDA0UVH6UcqV7FF9Ax7+TdUqbmmZiE3D3af4392/j0eyoGDI0cNMMQdOX2Vr7MX
JRLEdYSkEFqBns7Fx6iyO1A+quH2k72d9odTFXrw9qDOpduO4qQpw4KTd5gSr7O4
CU8gLAAF33gLn63LPU/z7bwcGcCrYBWjUpExM0GDm+zG+GTLWZ3fTVcZDPqsp9R0
fUG/I6+vmOdf0scmpnO5e/1n+XIKusmUNg15pk33yXVYUAEKwQxYkzlZ1PGravS6
KjN377xThRb2YfxmcbxQ6PBIF10USL0NsJq1EiCHEUpT+inxQ1HQbS+QnNLpBrWA
JUTzZcw9oE4/smsn1BZ0juXCNqL7Zj9Hi+nywW81fmbpEzim9NlgI7FNTu9hl//D
TdP82akm/kge2mlimim/wPSV3fHrshfTeSB8slIrQt2bSdc9zRdwlpGkIwZUl5K9
To5r1N6Q+eIobrlDys8YmeNLaX2MT1xiy8THwJ5SVBwWwvdm/hFHCfby5dy+gMi1
zc+XGdxeZVH+JCmMmayOKyHmK3+Ghuzu5XJaW+cuwjMBWrUIF9mYZhHIkZmUpuUK
JHyk7JxYohr7wzP2Ft3RFVAUkxSVkuAhvPZ3d3bOrSA43nNoHk+ns0D7hlaX5IuD
+apE3Nk1GipJjBNJCFzVzBvD5dVIFoQFUyq0bg/iOd6js2N1uIXW1SSgw9bzAiiM
Xl9t+Ks/eEv0hAGIASWTEbGpYBTz5W//mnmY8MNPpLurqkspMvEJN/SG9jqJQKHw
Eui9VO8x3W2NEu2v8+IDB+z8lYC7pbw52agiHguZwmm50Nns8+CBhlKgxhWGWOD/
dqFIqlSNFLXPowtjn2n9kZqOEoOIkj67oFWr/9YtYB6l970TTyIMw9UuOplAWGqF
mDrSxGbcuGD5SKKQmrwkl+dKXqREH+MhjnpIwXas3Rf6NWR5gcj1liKfK3W6+zdk
JPdJiNNeu48PMgzeIL7aVoRgQ+r/mZouP+O0iCboL6GXpVF2o+oJtrKSJolWOk6t
kOuAyz/yu3BNOWENiPraY5krICd75htlSbxKaul6BE7+kwdGdAd5RcglSWxT0wGO
wX/eaKmy4aSyVz86rFphpBSjV77KzdjmaNg2cPaZXcVluSYsIXFhMVicIkd2DpHd
jIo5uHAow0TLQWpWA+X5E42QiXdHraTZaZ+onN21gURJRwo5CYqh7bt2ye1UBEwc
+NaYRrH/A8NN466JtuTAxIqdTIhzp/MJwMxljSByn11f2QAvg7ValqPJMqe/IQTz
97UDV+lN3jQenpP3lmjdohKw/Z/NfcwsTuC5v2FjwgZfqRWYL8lL97fakioMsmkF
N8dcfZL025X5kIAuWOFyjjSfhtfDsA/+Ipkx/6ka341SHHuva0L3sFlQJCCAy6wO
ZQaOefSIXHpcjcl5vFV/QOnABPqV1tYFjqQHr1bl3F318PL+7O29FAIIRfeKnlgJ
XYVxfbOLWDW5ELJtVB4+zui1WfoeX3FBLC+yA1CQxwvOamBepziYgr6/TeKBjn8Z
E8zT3jAnvDbomNRoyaBwxDmy1SZEQjxk7j1hxYR9XwZNDMnJ9ka6nzDLD5gdM/fr
NkXtl72pSoDQK4gJanrOvywVlJk2J5l+EA5o3UlMWWAAeVAbpgwD5LZs9cd8bzjQ
IZqccU79CU98B35mwSvR0JuGVNPIlA8pl4PKly4NcmJQPUhk7qaza7cWwK/yt8rx
NELP4ZDg32wHpNt5vnm5Zf1XBoaoG4YLHbmMTVlDAVgJHhX6Vc2FuSRqI1wHXpFc
g0s/sz863ugbUItGmUWYN6IrA2vYnRTv54sHKwK8bRQffqMyz6dg5bpozz6JxHAA
7QQw84WKUZTaKR4IqBZIWKdt8HYXiU5UG2JnedMHK8M+iTBn3am6uc7xe2R08aO5
UURBj+dhS3/1/SjnXJH7xIvZSV7pbshYz0rcWS2FJnjbZCyzI2FjY5RXbM8SbSf+
QQ7WYuLnU0vlU5rN0cuemRDgazawlIS3k39xoOdugxQYFrgkbtjN1L9oItNvoP7w
Npz0VjzFgcVi8JABZmy0EDAd9ibkaAASQp8u82MKFj+nNZtY8pI9/dRL501lHiZn
OSas1AhzS88IPvv5SXbkzOErtDp4RPNojj7hXruHlBmz59p4XD38PVS83yUtm6d2
Ivtve4vw4+gRiD1nBMD8B7DR315z+YWub+NFc3Qg24H+UqlrJC1w/S9weOtDshHz
l8O/ztFrd0mz1M+QSlf7WmHTpBFJkMag6OEtWQpck8HjKtJ0VT9sPvj5zfKvMwA8
akdOSULG/to1pV8I6AV3fiWyYnfTAii/EhXspps1vSp1G2vEknmlqVqfGykCRko7
fWlXu6blFfajm8WR12Nhb5YgOMJm+oBxE437dDMHvcjaxJQSs645oXSN2EQy18u4
wpoWupAeJY3BXPEo+ViSqntltgIHrBcOTzVVFH/gh4plhoAI5j93WPMGuGpMOm8n
q9VDmUxVa6g9E9gNdAaGEYPWeZtx+0HYhc5rO1Rc4Tpfdu2ppLOUKHbSU6DadHhE
iiSm2jNCA98iBro36L7m/CJrd3wFeR2u1k8aThoMQyUcOWsGW/0vJdl7kY1NUyFG
nFgDOShTrbCqr5OzqdeweYsYJbc21RJ1tP8txC/rV2gYFPDzy7wy23F8MTJUy1I6
I0hQ8jQLcP29N4M+jETUoWJTT1fDwrcedpwOtNNImhYPiGyeyDPrV1uuHS4t20od
W8G4onOSdiNTdizx4S8mZqhGjygfnd6YabwDTK2GUKZ9CvkLX47EsnspntWoT+J/
QKh6oHjwOxV85uzNZeN0GqG9Z0fjIS3qmP6Guy/zx8s5rAF9uTd+KjqgzzSEQ1vQ
L1yrAx1wG+wa9iceLoBN1HHZzTIMTn3TLo0BrtLZpfHIOU2xf+B62LP+N6zBOiLQ
9Jd7bOxRbmYPAC4RemVbVpGfgIuK5rrnpszEumEqRS4slmEaL3PecdSncH1LAbRZ
j5oT5cyna5Ew2kQd+qtMxoZvhthArLDqHKTqNKwvLBUkmFtXH190frWO5S08mTPG
jKuGwRA20/Okar05H54EalYwzqA0GIGG+KiAxE8QAQaZ1IHuh8BDgX3wdkf4ygZa
erFcnK20B7E5iRPlLMFgKOpq4e0aAT0ztmt5ob0AXK1tswZPxQnL85nwM++xrmxI
lbLW7LvMhH0r4coPXAhR/rrIliysPj8//8kqjJ3qsKsm7mkipcaDFkvc1o11kCpW
P9oty9pPumpgpsaAgMahte5tplTNT5JCAnE3Z+CVm0za3Avfe3T30y5l2D6wWIXC
FTMkZMqIUhQww0A/miYTCo2mp9eBaofnlu5goUPl/c5dB87yNmIXbPm5u56Bmjhk
5ZHzhEfs2/z2BqaQXHVZU+cPjjpx98TBGbbWmMpiRBLQorNLvQvT0h5iT+Mt6aBv
ff2pFlxwTJSAM/7Wt/r8j1ctYOdGaBENLx8N+4D4nDsTs0Jf6lx3B5Wddeof18p4
K2fpX0EkGow8cHn4CyfVIfhfAvMYkWcqRtVH74UZi629eL5RCoO/DxGMP+8vxrzV
eKIBfApizzuL1GIDc7abRHtjIcnBhoJIKmXZi0Ucdnn8M8wXm7MT1FzbDq7eBVhB
z5uVbR3ICUkdcoICjcl/wbeLOPtytCWPMYSnOea+KdD1SIsXSYniMoIK5sMIellp
y55VXRR/3uUm5SWCpMXx/F2mRhUhinxu3fpR2eBxmJTDPw5nmJlAI06GTeMqJyYK
vw4lOVN4Fxa5kQnqSMvBxQrCxLQhVq6iokUmfzbF7fLosd1E0X57IG3ABIMy1z05
mymV5DURi0FQ1HyOTT8yqsdAd1dBS+G1L5PT/X0k7nr60uLZ5PPfrixvSPY2jSQk
Xw8K2/0gqBGAmvO0WGGb6H+Vp/0uzVarlih8+0FLxQyeyA1clyv/v6mhObjLnVBS
w6Ff3q/syGiSg4AQltcNLIkppfpC8Q5XIdNfo6Roqk7zwvaYUxs9aCI5+dC02tgJ
mgvksh0E1p2rSTtmcAB/HP8FKhyzK163L3SGUDlT0CFA7Ltc+dJqjskTukx/zqGI
GVOW/6z/ZS62N8sMF5eFIERau6F1Q6egUcvSrku9QnjvzXM/fbkPjY1hQdp3JGf1
PrZjSArq5eXezO1xwc2b2EW4l6uPvonPRYuByGHabAmOXac9SqiFBclBw9yJUJFR
IK3LfCIK++DdXvb02bN9PWuUC79NqSK9njr6Dr9qStCIbwNfD6zA6Be9K8XsM2Z5
Ng8dPQFSesIp7fCOHjLL7nyoegN9do8yJ55/XiBmjNMlbE8pa+LG570zIqxEupmO
ZvC7ESiAj9845vuPwBbB2p+acYlRyMGwbkZb5oSf95LL/lQ19CZjxaTCbIbkdGja
s89NEDYUIIA+VyNxeyGyMS1Yokjz1dCAt2hNpRZ5WbN4/vtyQPeU4BQiIvpuncrh
N1hh3U5Hy/RaKGN07r509CIvA6Ys4sRipXi5CGAR/+y3isNFQskAmWNiygAvivfG
UQvdTLmmnk0kADtpI1sNzikGJlJMSfb3efhdutj4R+cRq0DuFYQCKjppLJDn+osX
Wqbq1UjwgxLVv+8Yf26VrmOFlhklm6Pk4sh6cARPi17MzManCOxjD/8Hanparvn1
lyLofAJFgfCnne0BfIBNH4m4HdX1bVgACrGxs+7bpOVKbZswA6cDRkKsMxZNiGTx
5tAV5HuDItaxR4JARN/z4pK07doSExprV8TK9BePU7qMmgvpRegr3Xk7WFLSYbSe
J5b7bcuVtvZeFGLe7meSsevxTdcSu4dHcuX9B2q/PwrUkGUuQDO4nw6kkWA8tXhq
6hMGq4N0uNIvYNo3h7hWYQA3LlefV9H4z/0vxDanHvhH9zs4WDzMtLki/CVf5VRc
xlivFrU5iYwqNDPTnKp07lPcT0CZXLfd7/taluhZZfYgcjUExDZmgVLiFPD17kpC
WSJHR8sAuyAHLwLtsGUV849cgIuwQgD7e6ufu2MKFM1lYKMoFEdk+ORBbBCP7Xat
cVeZS6p6KPD8AvdLl7F5nAwWHjl4tU8miKaVBMONPYgYmrWFHTKOzl1o6lYozaVm
n6425ODaizouqLmkESo+2iFcqRf57UOLY6vyn2dmgZYBKVroST/B/0R5F/MMV4T7
13ql86DgmFlU8k1YPwWNhMMVMHrqzWWUNKN55da/9kV75K/oGKsu74DVZZBgDhs1
9swhFcrNB9NV2Jj0T7nKyxEnnQdVzlpXkzJaNMYX25/uYP+gMTXUR0asUBfS7P2Q
/ExgrzaSOU41QFo1o4mR9xJqYtu6Q6gusoif8dSauaCIpHjNiRprWM2wkOv613Fc
31/no3XnMzMOs0jtBTYFUZoq5utG0cwsTkodSPm/jKDoj/W+W0wVnGcbdFhjgHM8
mw5Amy8NTy6iX35ciBRw7RcemqI+PUAGH2/8Sz0hCyCm2C3eV6n4nVeMj/iniioR
YTf04/37FBoN2N6fHJ1SvocAUqWhtV+K20d5bIec9PcaA4w/8vqgiS/r+X1cypgg
0XneCrcVFP1xVzI8KlDLgoYmn4YhqWQbjiFbjD99hYBWHIML1R0Bk6o9IkBKP4Nh
cBJQhtBwRNbVUHYsgjN9OEe2GwFOgzNCfrip0x748aIABEJwsj2Edbta8CgTnGhm
JX0tE4L+TMbhSFxBZZuqdAjn8NVKtgmBWAkzOcHIfN99NtHlrZB4eMFyrHFw2Erb
8aZPph1MCHEV5FIZqqCvppNhe1LSlHf8Osq4f1Y+0qvEXPSP69a1dXhz3eV/kVva
PFIZqz/bPyvII3Evl6YRfmWGACzqs+U+CEneqhT0W5HH7vDWlZorn0vZ8hWA3LbG
jhLSs90eH/bi5xI0j7X3kRZfbEsNFTm7RrEQ6WBLFOVgw4HpRva1DxK5FhuWEUA+
jH5sDGvkXcrbxrsCoRVa7GX78ieXfSfT9vpubfDFnlmTpNJa4FTZUDKoj0Mvh8Mu
niUnzTwOqtOyRlQP4pQLvoiaKaS39UDZTYuhf1iJh/lhjLjlP1/rWhv+w7ObyEAe
LFd32WnEt9nrauPKoF5O3LN0TzimJ/mPZRKPcPIkU9pC61wB7CNuDLN6uSpPPykZ
NirhXdHFH+I+cZyRrFafCPhtbiL+Gpn0zcUEyotJ1TVGWbNsXW9YoTvmVLMCpnDm
Mk1jCk27YQG8F6Q4OCVfG3h8mC4OOs/mec4MhpjpkV0e9hPNfz/0A3ULBND0Xeka
5RMWTfAVP6I4gYjQWIPs0uOwpnieXQZPZiogtCJ1Y8viA4I4BPGKkSWoasSwOiOo
3NroGccPY6WHOV1k+XgUj1Ov4tU8wFpXueINBALrmorth9CAKHWHjecPE7PVDhl0
oYUNbno39EyiEKKsTELAIW6NBKjcw9RaU6esF7qixr0Tp0f32WCUwkLLY/Svdmj+
kie4eDi6zbAHFacULEYPzIZjWWrmiOurfH1NgKFvpcSwEJadEuQVZOUinX7aVrWj
bgEp9F7t007FWjesYyvG1VFOXjUo5hSr17QJam6jF+CP0KFfB0LJoNaKic6T79La
4Mz4HAN3R6BXvRAaT+imNDnaMX2QXXJzGPkvTD5DjXSyOoGo6wW5cny7gHSKRefG
D6UIR0+uCiGYyEMtaLC05Q/IwHq/YUZtGloWnkVYslcfHZ+y1ef1vg1XQ6tBxyz0
PwRZVuR4lc+6YOWRMN00S+Rwj6s8wQ+7So/0YhLfy2xrUUrIIOto0tR59ZUI/fKU
CgBA4+a/eIEz3GEt3S9zWgJWi38GuhYdBW0vT3xdXOnVdP87E8TaPnOiJIBEeGoK
e3P+LfE3rOWwspnoz1YNED4WqaTWP2ZmNDSqdYiFPqUn1b8Fibz4XV7DdwOsYyDM
KPmCYXo/IR72DuBe8r76jMDvzbfhaUqTemzupTlF3sQ6njbdmpGIjTxpbPXE1Ga4
/Nk8OW7j5ArTdBAha9i2bge8b5CAaSXs4a40rzO8Olm3YJZR+kWzsVH6YuKe+J3f
jEMdVjDBjrwGtQsldcHy4oiUzL+KvelH1sGe7CGn8jB4j0AR9RFgBfRQN/4zJg05
IL9KHHuUrOCXW7RdsBSMFmIqoZtsFDc9+dS1FhCy4P7i3gbvdA5DfCapumd+pSaw
+iOWVGs8WIBF0n/J6DhUzYFncI1ISxlWE+AzU62fnVma56Aj4MfLyfwBCYFUfZAJ
vcWBn5yB0ZTNKwFFWpo2cg+7RDQ6E5Ithw+Enm7ME7W47qOv7Bn/oXtTYvv+VilK
J3JYjXEVIblX8U8KTuEOcRS57M26tSNvLzEl+T78ppqxuwuB3TBSZhwcdO/dOmHu
Y447h75UR9vH9JDJFQRpsvhrQCZ+RrgJaGjoPbYTkymIx/jEA1zk44i1fJ/EdYtc
6JeMipskdd9yJymd72wkEm7mPjMRUEbNzVWMvi3EaUa/GevTNFhEj4zncp7bmmt4
px1S69qEU47ZetrMaDmjlD+tM8v2GRiTrqjtJTXpAJjy+JME6/UhZ0KhTpYxZUY/
KpDUNwBTYmGic2GZyUmStXZ6vqdkrcfrIUi7VyvKPX+KM4/6P9DysqQbHfwr1bFS
7K7NYh+vVBNIM3tYScXkkLWObSq/LFIeM4YmDC2uTB+tdqYjQdyRZdjwPRNx0f7I
Xe3GpK5cciS2U2yF04yIPxQvZb+b5hVmuOzXRJG0/GrPGaeO5t+VX1eMN4c+IrkC
FU8itdvpmYKMp18rjSM26p4c2he42yn6+t32uRfDrSCFe7mp8/dxmt62szQxbmVi
iLsN642PD/X4BbIEhsTyrvypcaPu1qxTBeusWcmtZd9G/9TWYVVNh9ThVwqM+Get
nIW1NhCGMOTjVpJ1fHnnoJhGs6o4erVUnw7dz20RZeBTeaPi+EygQczhHkGhxYt+
wSrOGC/7yfikMKDkqmC90H33Md8RK5VfnP7QNJSL+5ldR+ICNbhUsJbCNcuVo6rX
wAf4+sOnGqSZ4J9Qzaub+BBxdRZRWmbGSidqxu3iDKxruoSn6oee4Wf7ZmUThIGd
wrWh4lGiFtITvVB2ghnKy2MlsHD2dcY6zJbHcjm0SuFnrp29O/t8KkncbH42lIAy
oDtHaalz0DWTJLLWYgl2yOGHAz9pEwvCP0nVnO/nKKNZ/mkkGpmj0l+0cm2Saz3S
mcL/niDeYHmbV1rEo3KxOSn9shB1rwiU7vMrRe6qo+sKE7gvCBfvZcy92DDBep4K
PcaDQEN7WFYn+gWzLtfFhdyw9I9Zl3Px8FE5O5FShwMNcFCwevbubpUPOOl+Dh/f
kl6BeFXvnFoWpvveTj7MnZf0AbZMueIoyOCAKntR6avkYfYxpDORr3hYdPmT94NA
O0v9F0NjS77W3xJmBMBqycqiE3yPe7AChmcLd0B6AQND5Bmr9i2jhtyZHTcc2514
8Sb2yLH7hmH2YbmekhbxCiJySub3NEXcMzrVxp1cg8GwzAakE+pGWB1UFlHTB8r5
keTWnwpW7+/9QPGZvFm9t2RoSzZy0mj3aROpBgi3/Qhp5Z/7u7wL4lR1Bvds93l6
iMFvQr/8z7+TRLjfrSdc+wOooRVwbqtHKBJ/ZzBdWWPzhlC8YbZS3as8JfBZHT5k
ynHeu8DWCckX1OpH1Qe49niz5ecNkzQc7JwgjQBc+zsJm2hDhDHHvmbHYCilMhEJ
U8VWxKuMPtrCpik6BK8FaW27f82a4bHYVcMSn6llSYEsO0MYtddcrBBSgZ/LlYkn
B+vjXXAYBYRuDR2VS3sRltHxy0VNy4/KtX286g3CVdOW8cw+0fSC0DYtBVw55avY
bypkVxa2b/vbeipK3pRwHydCWf6q0plWeutf+8cETBdqcOYJIEhRKhGPaM2zo68D
LGCyrBe72pFyzi5k/jgfW76Sx6/POI7S+seXnKXkbBQlc3ZUvfr+XehZh2FuqUOe
miPlnOy1wlo5k8T78ywplbIM4p/w1nv/lXcWC2BoGz0ErnBSlyX2RHyA2cXFNUkC
nfGHElBUOeBSwm9+6pCzh8GGj1tWz3wuXMr05dqXBTZQoVGWjv4VubTA61HayXpp
88S9lmZfYRKQPGXlpIQ4SztuMr1vdZdTHB6ffXkaEUas5EcMeZWWlAJ2/XKvyF1q
1tzLErzONlVT+DbuNsp7dBEqQAT/8njw7PxkW/rEPdcq11IGWs3tlFu3gl1bGjeS
YRnIOzCDaI3uTv/Pf88LrDKk84M/cLCNMyPX1nqht0CHBChbIYxO8+awLTCqaT7T
2unuSdAr6vCqC4mSF8DFrHDVLM+2y88UhYnpmValqtOM7thMPpdUvAAIslsBeUS/
0SIgFhLC/ryMLOPBmOs860XQLSvbg+4Ac0aTAABLmI3Vh6cyOkwWKxE6WYJUWkh0
NrLo3H/x3N2At1DanrPxJfZauSScdH61sp6N7ywUFD5Ncc6FGVeedRIFHvxYVMTr
bR490bE2ZgdwFv66iXfgKCKjuIg+fun0Rpwu1/ce/0qmDodlZOjGyYNaMXpyvKE5
Mg/RHpuR8h0t54qPKNg8FXg3bWchL98JsnW/Tv+7xzQeAE3WKvxIH8dqfIhNqiEF
Nws6QZHekj/shxi28jKZ2dLwMsenA1VtxxKCslJztCFGTtJgTznAHRNlffZ44keh
sRoLaZxjMY/k1ZYuhmUtG1bMZiIM+W0nkyTNIqqbSdSjCNTxWyRVF6owKQ7Siubv
71NlV+va5PKD3MQRxINGLp/EM5IzTXlWpKuZotvuycAm67szKLD01zF0b+MgpKeN
f+vjQxzMOmsUqE62RoAhk0+7UuqPQ/9mXIdKTejciv7RnBKpOkEA2XVG5DcV2rzq
s2Jm8H7DNL8Ej7UVEvY8vOolom7/RBvgSTdufM8ewBS9QNe/wEkX49yz/Pq+FqK+
mFNi6tQqvi1bN553WbaINiIMDOXT+SOP0VRimDchVN4KCW/xe3KuK0f/8GJBZd6s
I+cSEAtEtioUWfAqsFVFykcesVbL4O4hbmqpnyg6vd3F/DKWP84vslWqG7gF2xhC
tyqig9L7IvLBqMnpIxS8PfjYCG2h2RR5JCVIcdTZn+Ju1HOkH8WAiYYU6dbgeY5A
r/F/I2GKtjcaAXMeju5pKeT4TaeSg9BR9sRxoGRkbNRWD0cBSh53eFsWz4Z/CqZV
N3qnRU/VfaBCTM+3HedeCjn+eP3d+zYw57F78d1LiNlPN2PciaUCmSg2hJ5TddWw
v0TbAHhQAnu+caSKy+I6elVjA/66RfFibF+VjwUhaX9KliGCNuGcyaoWtHeqUY4S
DS/u2CWAcJBBlNmTIRyASBa6r8NqfobOwVScveUdX43GCWdk8oOdK/OUN54X4DvZ
PioI6RI18LzoeC1E+Hh7koaHJFygI1DU32LzyLVPbHlWYuMBet+1iURbuzuNESwz
PRy4FayMwg9sakoYTLYadJccmp8PQa7shn0oxB2otHyqfyoUhUvH1pZl6iW5ISYS
UUSfVh3WsUJ/GB+OfCD9Ckd2NJiC4lG9JU25v+IRS53fcGsjkOIDqaAV71KuSZtO
S4EPgkZ7DP78KoqoztPw/VDG006oruFpzK6lZZ2NLkI8lGjvpr6Yq9AjQPU3L34x
OG+xbi3EghWdzVRYe84cueqCkHj1/iMaxvYvAlp48QmprYU+ndTitD2cav7gE0Rn
uF/wm66YtTh9jx3Q4bXJjq/waiX/Y4y1nk1isrWBAfXoxJd93RStga1BwQbiO0CH
6G5dw3IXUtaLLgDwOB+zKHMtXLBn6egWCIDCClC+Ksx0+7K/nj1oNKu7DTlSJ97U
02YpLOPxNgLryZB5PSCRF3ocbtWIlduKNozA7FhJN5crykFSxsKLFdZ5KyH88+48
hRq4zegQMrZxVpmhSmriHdmzKiTqyUhGohRSZUJ6Qu1Eu2DsXMzRGw/UVtM2LWmu
QZea71Y4Y09uh36xDM8o66QutUwVSBw36hJlhGyJ9F1MltwNEZe55XkoKjgCU15D
lFImgyGq5eejnXRpKohJyzIMyEvBS66zyNx0KOvMXpy66EvQ9E0KjIOKu0XyiFJu
9OsptEjJPmA7quoOonrpWJ5SosgOqptJ8z0WaSDNHONy1K1iruca9CSr5xcfedOV
vPH3NPXJKdQX9DrRWjkJyju+JdJJDh/K9BX9WU92Dc/GfGZcl38b2PT7RdXPFjb8
sNJIXfhHAZAWkMSEDkB/vQ1qFwI99m6papIEDCDK2ZgPGNI7o9p4dxCysOJW6+18
OZkUBaTtRka3ksYhMwS3QnX2H5h3z3aX8KFWUHXNLAGnUEi80XFLGA4knZYRTzCU
nhOImuP1azl3Vh3uWEf1fw1Cx1+FMndnWmXBerXPOTQiPRBLAFYNyyBreDq66/tO
C9HSTFcAkfL1jMhpbITM6aqWX1HcKcqw6R8F17o1f3sEtg2ebsv9XgytWenFGL98
aAWbBYK/XzXeU9r8u7znTxm40CMeoggFldJ2+cdrrLhfQjmw5DYd5WrnLx3MpIoN
iMV6RYOn9X4z/k6bbPKZzdOAl6NZzXBGs4W3lsbwMU/6V20gyifSl1dbr6Fg9V/j
Jx+gI87F74dRUw0ipgwYQQbwmT95ma7lzBT7b8Cm1M1Ze0bYF+d1DsMqVk85iiKL
La0oMOSYTanF7O3E0q5BmXIR6os1/srGFfiphhEMgOb4Lg8HuzjCybawYA7R+3QL
Hvy6cLjGuPfGGydT9PlIO7kGXNCX9zBpzpDJ1JvUAvjLZgYGOUq+rrzX0kWTn/lJ
RnJ8bkviQwRJcI0u3SdU4Ht8j1owZy2xEBelDdApqnxgLKX2dsEPI8HodC9Bh6AD
yMhKPRa0GymDXIa0CXcZajTk5yNqwpCaWJmqOF8naPweG+3FEHV7rp0CPx0bzNI2
iFVGB/B0YlKOacSJNLEonyP1TVEvDxLFnifgCVdYy68WO6vNqNItJoNyLUqv82RZ
8e3eanO4GM8T7zLEItyy6lQIA2R2ZI1qeZELWUh6aNkO43AvdWvSjqcWQZANFufg
b9OU3MdQPFlukO5++y7CP2O3oXFETsHgdyfv4YYnpqIyDkJLPxiWM7cVBiAo/aKZ
LczVjlxPjO5HPk9iHQFvaT9mHxl8QJ2iLxgNFNGq6pd8pj64D2eXPnr/dUfpXfUq
cnbulB7o1Bp2HQ8HIJydOaEE4E1naAWhAyiiHiucH1MD+yQIZk7gOEv6YM2+2Vn+
EiG1tsBzGL3Znmxn40bcpbF3HxkQ6oEqFilSbL3y6SUST3tBy3NroMf/zs5/S6V/
EeUrvKaVlptoGUEbI8FQyBywGEAnBjT7yAjp2mD/dyPN1aXBRXUFq01PNNQATk5M
ApiU1lVJ4fJaJwQvKvwwzNJ5sXrKiHfkECD3YNVvMmXOjiGPoYr6k0KE44gnc1RW
cgQKQbr9qWrMIGekkGcve4iDVJ6gfKR1zME0nEn5EyxCZe/OTEFFxAKV6QLvLcRU
ubZS2on9WrEbHNjSY33bKINdlrq12aaZD9e/efok/m+mrmEhMyPeBEFjm1V/Xhkw
PJuxIXvb3I4MDjH3tH22z7vUAwYttx2kg8GRJ47lEX+kX96h/QPwZDlxWkeSixvS
opIhiNhPHJoZZ/vANqG0yKmAAD8gc7OAlJcyQCSPytoz0N6mni9qYZ1X4PLySpg5
c86+OomovGu595MwKHS1VIwhNN+zxZlBAuJSmFtMy/IedNXZLFSz9/BXiJT3pZWC
Eglff8GeguWp0rGbcFv1XqhBqFkFMmJiRGvsITMo609Fk7dpTF5kZZ1CS34Tx2oC
MxLoaSno9/58bSbzkacf5AJdcQDYrE5Q4t3jQrB8b1pkVwVI9BlSw3W+XNRCBOB2
e/pKtV2Pqpi2jFNgEZydhwn5U1kcLZwgVzxWTxFZj0zvsnBr0HYv5HVpnr3E8ATE
TOWhhCQHZhbfIahwXC3yanoKdtsKM9hezGb9Jaum1tcFh6WOLVg1SLBzMfpaR0CB
wY1qI/Drxw76r60fTfsOttwZ4x5bUGghGqYiMD5SAQ5NVdgugjU+YQZty3Tvq/Ql
jKzfuCK0JYe6L2dPRVzuW+hwcF1CB07ekxBAAH9cTUcfyJLugGh6Z1TVv62FvECi
3Y5jjjAkW2esdWtMixbmWDOD5CaOZWaBgg4WnHJ7gP8YmU7dHVQ91Jtl4/EFCEmH
uWqiKErX5mBt7JAVV5jsjvXbHRi+Ks2Tw6IvlljmMB63iHQmjjd1yvqfv8ILRX7p
18fsw5hqCI7ezII9xAn5cvNBiGNTqDVPt/OKRK0thn0MfgdI2EjKzs9NEv7i/k5T
58X8gSJddTE+zff/xE1fh4Z0d+6CeFwwbTjLRpK7bSmNtoyo6S0mUiCZj3+RNhQC
gaizAQ7FtaeBf+u043uqwrSP/RLK4WrDaAf+Q0xGzlLWcLFH8i7bMuKxqYS0uQVl
9+Md6ZPUW/trAJyH2xeyTp3cuUdW3/NrzQtLgCm2P8s4V/6MABgO25/Px+xam0pA
BEj3xNipP9nCm30VVfCIGtn4xsyOs7KE5CGHZ0arkxiE3NXNt51fZkcyqC1Uixq+
xWe6TVAP0tAvuCxgSm9il7b8fdVhfTDzagS8vxsPi66iK1uxDRiXT85G/Ufm0yIn
1XduopywjkvpokTpiN6I6+qkSK6WNqva8ZXnqUtbVoxW0fveA8WzG3ruTfz5vvPT
aZC/SmGuUAlGqRvqx6znFCTfC9SE4RPnx/ll04quXVw9i8m/ChDoQhHy+qrwzk0Q
meBP2G5HuocP7hlt/pNr9xE5jtU/ONSInQ8dw3xwyCEJVsi0I1Y1brmiWPW3ATWZ
waNF4iC/C4S+T1j2yxhCXaV68R1THyrzlqB9DfLjxwFPdY/hYuiKnC6MFqDfZwyf
h+3JT8YousQiUt+s0qryJRCLweoEZsvFOexw4LeFsLYZ7H4Cqyz+N9uiHqeKt8M3
BvdhlYLH7uiRdDB147wKE5CtqN50WsVg7IyiQ6040QtSpYHCp45zKmeBCgyfvYob
6NjwyWgm1Zfusy5/azY7CuZd9XvoWipcl6dpzO4iMFgIFw16kfiW9nFdUG3cAII3
lkbDm6BPzogGeN9xky4Tqcb0h2ecLq2ZWfaLAaAj2HPYK396H6nrqzTDHhKnAPAu
MhwrcMxeyDv+n3yorxvfCmxpiaExWF/k+Ph3mfiOyiIkEV46pOMGhMRNbJIvus01
ubBrTYbrfnanA1qXEMNVnVNxbSjzK5R7oayhUadjiuvALI6AOz4GFdsbiJ/3lVuY
3blS7MLtoWDcPvm/dDdfSEJ1wzyRLovIGn987mEgVwKDw562Tnk5e5l94bgqH/Hw
rrWddB/3+QEiQdwu2saaUlPrj9Esr9rCRam/Q8sKiPOlC0q8L8nUb64FEG5PooYd
g20PZaKeteZj6ODBtkGSZ07DyNBb88Aw1wxg9Tkwhm3OfHq71Mt/m0GlBfRXLEtB
ppkCV++WecH+/LBjnt/shUL52Bw6gp8MVeVPuy/VVLCQHITtcgDHoG5oFE9TXeHY
nQKWq2h0vLE7d6ue8zsEIYOEeonkRLncp9Muv1ArQkqdGzgWJa29q3wVOFBtXOYy
xTv5KpQ+7hRjlXRuqK3z2FPQzVKe0/Dpqs8RjWLDa3jtFmz2dcYc1Yk27Kt7bToG
qpHCnQGOYEtD7oU8JGtbRYrPcBJpxJz9CfhBBrj8MCLPy1xTM31LTCDx5RmwPOiN
8p0bf3aPnEkC5PCy39EzHfbHJIFqDPKUbD6J3y5eL3goFdfei2olmp3SU5Bo9Qnl
RHOHf/FnmuJ08AOy7PQjRFyNmJ9i7vDG/Xma13SytFDqb5yli4PxqOcjanjAIE3U
CVz3m4JvqOyJd0zGuweHDxXI41zZnPd5PmVVKLSvowAuzqPy4Pb+Z2pgmCCOs0e9
vdDezCzyfMiMbuIZLCs5bVZXKyXN0PWfVlLygNMRBa/TdIFu35oRegM4ol+0Yrvo
oGxcAwPs8OGX+vDm3hthUHIj+xPKhHXZeUVHaeI9y5b4mWY+MX4FpMMqbiSXTPOn
wz78sD86oYnuTpChyHZ59kQMTtsRrK5yMjo2OFLRoAwcdmB6fZZTdqE6f8PmAbpK
zFs7weO9Qa0t9F8CvHs/DE5hVgX4t3DEtiCeXQ/w65AbIrZbbSNrRUdoZtY3/ePm
FLClB/W/Lleco+eoDvS/rsl6JTVI+3ATaxuKdmYizLroKKUU4bAY+GTFDiKd97A1
A1JF6DNND3QZtp6vxO0NLJs26BrPjjN+5K9HcxlfgS+KBRLP1emoUcFTlC0MhXED
93s89EfoZuihoVlZKVxUKcvc/9OMCgBgrNusg12NaV4/87NO78D6M7JVS/Oiftdk
h/BvnTfZaJEisMIryb1xM78GeFyWVk0Gckd60NYd0Oh9lMpaahp16qFS36NqbHLQ
iVpe7HR3pcd0FNAWxJ8U4Bmmled69rctoDzx42kqprmLUeQkl0nsxyvyQvt496RN
8R0AsKATbLOzFQg/f79dZge77eyZr4O4b0dkV6JE2Kvb4x2sj20q0LX4aWiri/wW
3kLNaq/4I7vkmoeiyWvVUb18HfiugQlgf9cKmaYAFO7Vvfy2ZujGSakOGg00/VJK
qIuVB9uHmSogTygbtUyQDJCAagaZmdfH0A21FX1wy+U03r6/6hRUW/SQfbRLSZCU
49HyqvORcY6mfe3Ee8dAooN6UK5P2cqWFlHCy2cX073rSW9jcZ1DXBqpTYK6UuTn
vjFH9wY6zH7hRc7xLu1oazTrWE3OyrfokvQRBuijxaEm/jbpNWJwnlr+34Y2DYVI
J98eUdsdd6GIY99Au3YvVV46WRNGUeJ2UhbffQKYU8ajWMWIl/VXr2fJwrC0Ozo4
ctUIQ4BBkKkyWLn5DseMRQvZjSc2qA0OFdircvP4p55ZnrVm/C5s7oG4bDI1upxH
kw50tpKPuqkDTweNBM0I3q1fz6kKongT21hk8fJ9Btn0Jno4wanvCk48TruQTR5W
ubRopbwBKam5T9FIJFapL1NXqNUwaN/f1wRACalTYk+MDhlPFxjOyJjAOKtyljoo
Lim14pepo8Sp+GdBhRqS0IkZAf2No5qXd2MpwRGxPNQzAt1K1JYc/6o/67A7oj99
hIcieOjk5x+jk1nRRhDXTkNGakxqoI9mtNpmzkw5uociyx47ZiAcAXN6IwFB1qtK
mQOtUBmcYflctodUqfXX6wynfGepImeIENzsVG+pvdpydnbjKntwqMx+E0xuIgsI
49zBAHPIn+V8KgbZ4WcK/LkKDFo1slWOXD4nf34OY9MDTliD/zdvQwMp/vXKi1tu
Vdx0qJUU4BR15VceikT1j1fDbTo93CmxNkitLTAWSmKTrYDRwJ+CliNet6/QTJc4
7qaYYUTgcmY+P14jIBjv1wcbueeVCkc0Se3Nlr2G6D/lJvymzZokLWwxLxdcoBkm
zoK4sW8pPBUq4s8QbGtEh5I56bIYQcFgAk6ev4UpeSvAak6TwGUl8233PGPr2zwB
ltu+zI7zOiHrJGpsStemNzlj34ETLht4rl2TTk7yWA8e4pOcNnNIsBHpV2W0zslz
4l3yXgm9gXE/fMjhAKCZ3Wkfr8MKYcYnAKvpxqhLRlymnZx4PEbNTuJZLG/tDRrs
06oGyiRBJgqzlyhXt3RgRw2V7y8MK8sfFh1hRt/DWuRvBcHp9Q19mk5cgUmuac9u
x3Dqt0wyL0Sx1MGLHb3xKTWBINCMj8MkuOL6hzhliDPoXDLTXy+kFhhR3S/ZaS2Z
ZqGd5oPdkUjkrd55qRwgC5xc2QDsKXEJS500OxUN6aVOL52AUMGRD6WOizyLBCvI
i0KTDoEE5syKE70jXu1t1U8JBjctVIzU4AJMO/4lJEbwT30PxIxGIlSy4d9dM2bG
pcf7lbDzQ5r1zMwA4jRAcJgvpIKXEd24AGYzrdR+Aoe3aac1BRlMLKvV8qYGC1Ut
lY/27I2rhYZHBLXSwUZXfqviaArhMB/TosKys7ImPDKe31XSjb1bWhWa223gtIC8
Df7D6KJyq02wdfMEXdTswqS1S9A6KIWrlHttBK6L6VbtUwi7Ia+ooitUsmquq2B2
uIc06Ou1YlsRNUpOY5l+PPJWTGqxNx6786CD6Gnx2993HZuoCxEF2wnPwGYbgCt0
msm+gzOPe/GahgdTXOyALfuynRw0T3ECUexZLLA20881FjkGq8bRp3r9dw6VRKXz
qjQy9gO+jgx6srPFp9NiiVovvXyJyEAZ1PRJmBdmGCts8fqaUsK4oqAFfug1eKV9
B0wOZr5uilNqY3PmL7ynxmD813MtRqlx4/e9yqL4u6sfMzaDuL3BuJwY/srRWSBA
1ROVugwMc37gIRk5UHwTX4IbRaYVH5CNgGg+lV3ZRY3Vd/RPkyOe+dYIEN36ykI6
kkRRMQ7OmDQzKqeJrTHUUCBei8MPbRqR8XNMipVc58U7xf85kHwEaz3TqiIWHQmI
sQojmBRRodDiAw1dxPPC/ndbxuwNOIpXDLq9SYqY+E4Va6GYQRTmeT6+e/zkJLpD
UEclqONSz4Y6Hnt3CHDXj6KWBH2obz2UES/cfKi53fYHjXTM3KunBvvOQ0qUWezE
KEiE0+ooUBw1O3+doYU4+AAlVdtsXvXQvl310ZltY41x7XmLJJmuKX4b9aZVnhHZ
Fw/1W9Oe/nXmAf7wkvN2FlSsUOmQxzLwoNOKipqSED+VCRCF8ohrbclQgeP79+Jg
tAUHWI+zN3pgxv78fNLBlX8y4kZcL0EFct4J+1k01Aq0PR7Mzyj2ZDvtwrUb1Nho
xRvk/ut3eNeFmOKfltYxftFpA73/WDF0NTBLQ6bjDjsqbpTsKCk/Ixn9vUQzwfLs
KiX5d2EeCvr1HAJ0irS6ZThHCYaq6jbV9d0VDrIaLWRT6CSIycpmzaZBjD+gP9aM
PLhNJ50sf1JQPkgxmQd+5ro+4F5GMnRSi8xi6VMWgkzhnk9X2O8SrMwfiOMVlvyb
IFFF8c0IstI8Y3//aYsfOcD1m7dMCKpBFdEGieshud3SDZ19S8p9v/MBNaT74O+8
00EJVrJMLkvXevVXVpRg+7HEoQdkYFb3qWtW6HU3SZ8+pCsgdFfA1Wx6/JvJbsyA
JpGDevr4oyV7k7d7j1wcCcO/ffNwtCXNVXC69T0PPgUw0oUt1Lxeh+kctLrmfk8D
6b2dhfPxNAA8r4hzx32rzW/UfSWPTq5599IfG51kBs8qgqVRzr63dgnHx05m/flM
zcs2FjkvZMauJNCyJTCuy9hBHM55/My7x0mPNmyFkuue799nfFGvlq83uSOjzjPk
RX+pMrD6Ohhs0d+g+pYNFgGEjaF1jmQjzdntsZQQp77Q46UqNAiySroaiBH6XATU
3dRTJvBh/mksRF3hynBwL2Sj3C7QnyBcJAOM3w63SXGYe0xXlKCe4IyUVVpYwqCh
BcaAoU2tDzNFNPcrT4qQUZAe7kFM2Mzfe5f0wC2BjDhDC+MPxm7N7WMNOG1ZhIrJ
qoKcdFCskHM2JKWtRDIgTwETmxdI3QWV6h+oLIuHNslB787M/EN13ZHLoXt4wGII
SHGs23P5OHM6QEO2xWH32ATDsFe95ANDlafJhcOgrm22dYdiEKPMasTI3X1gaKFo
zTsFfed8ggHxr4fm4wqyNy6mXGvc7CUWnCDXZIJbpES+6oeN5Vhgs1GJkbuRU/IR
5xILXldmsF+o1mBh/pRqT9Hw7NaJJXWRRtpELP48OUBHLh3vu8lM0Gk1gLVdJXus
Tv6QYhDBeIXvH4eQehZCXkfIw8tEQPz9+C9f6j51lSr1HoS9Nu0nxsc+wxZqJnjK
GmKGqbFojI5OMEj3B3+HhShehMRLoZNdVwup55/9/xgGLhqms2DdY8bHllAifUAq
RIPFQaqlNAu6SVyD30DKo6j+ciqk2JghiYQnCc+O5iYOnJLkxk6qnqW1fyH7PMBv
0T4qDbfJ2HsC6oWcOifVevUB6xo7m8mCHz5fxgVYAfvuqDO2WLlFUY2hqh0DxiL2
t0hORxEuxHCrIwIJZ3WKlINWVPikgQrJChOWoQMpWQSr2/vNC6PH0EYnyZeMZ9ty
kVpEx2XJ6cxGqpA8NIfEK/CVcOA9p1By0RmGEYmVh1SF9rtwdjs+5mReIhe1et5U
mdS3ZBL5TxMu8fe5qqYuAk+tDbACdhCtoUMjjfaw7v1JqSDva9U2ozBPFAEJ9TR/
ojcH++2LgQy86tm3oorxOsbAs2bioVJYjoRxEnrR5ZTHlDNaNa6jetRXtWlg5knI
7paEjTibN3cYvfRm5exUQTjAVDilKw1qgXX6+wuwv00Zwf3tlSrhhwgv7vv8Moty
tnkA4uF4XvIGsM3XinyewEsggog3QavdCHnLx1+XjG53UCaqllm9bqQRynG+1Yz1
+gkhrI/Lz6FRQAzKKNZJV+UON2e58QK03UQFRE6c78C8b2UJso3p91zLIdIU2sP8
Uv2V8qWjHgZcFwIix/6m0bb5Nrk+e8uYMfI9pgarBQP/AB3xuA0muechYiNTIQo+
y60JUtKocXWQkrvWsX3wlSCpZsnUCnhUnTrtT1RayMwdrEVcpb84pU7UxqlDNKb4
lEQnLpWlUL7DzKXMW1sc+y2Xeo9OIbEchi3yTwvdNiRL42FHIWUXhToOBpHjLVhW
M529gZa7aw+Ku2a15OTJJrIMdPCfkodh3MUkjKpT/OhM71Oyc/C7lAAnOQZzJ5cJ
MB/6A+jqaqxdC3Mcv4Cw4vC5AHevpGJL38jV6eIO7LiZKXzvNX5SfxrPhpmlJV5H
v3U4ES6n66iKzey0Y9FFGJek07Tm2wq+mCAJgiKzbWCcV0S8aPyHVQxWfhsHeNRY
E9OmZClseGYEOKrlpQSClF8Q4D6f43fbB4G7r85jDmZ3fHMHla5lJ3ERpplKkTiz
sZ64Blu74bmHqozPQyfa+MoqDctCNN7IXov9M1PgT50ghdDV8Fb6QwY+BYLrGNAk
fgmEdz6vp3d+yWf1Twgev+U+CGF+3eQrcnalP8Rggyj6r/UNuU6YZj9nYVtWw5KY
a1nOZa/5qVSf0J03yPUzvT9VCQe0ZmHGXXKIQP1ForkSopVRwpQSgpWTlmjgUP4y
45Yt68ohg3D5/mZmenobFjx3nDmcgxAUIy5DpQrngNsGYYWpqhBGxzkm+Fdv5CHl
iybF05gO9OMS7rUVrfRaKn/P/bRmDRa6obYdAO3zQ+TAvNYeitq9fokLqQO+a+bC
nEhDn1wBQk1RWjMBP8VZFRviud9iS/S8C7SsQ8UkHdB4WARPdGvo1aWLUO9EdFmZ
Cko5ATKuoL5vYZfW1CNYdFEinQDmEwZJrpJSTead9f+SUNFvkOlgXnRsgtPcDYCa
Yt3Yi41inBYJbhvRZMQ1j8YYnZmvScmQiAXUWZVIjpcbUcJAR8UONI/8/b1Uprst
/DFqJtlkQEAh7HRDp7KUakgBWz5kpYLB/t7h5chEDKxdUsmNrF5j/sQ8XwjQsmq/
OvoZd1bDQT5lbSIwkbpyCwR8I7DZC5DDnbpiApv2SITt412zEXhNf2ekSuXX1TeG
Z/Y8Ta9YqdDnqiCg49C/ilZ0PORDevdjTBqHnVqHx5NPrJD/WsV4OrwjAcy0v3zB
p64UpNK9gPWwcm0nwL32B4uQgfW79MmpPsuzMHFeB6UW9TWjk+iJ8hbqzUhfeyVB
PaR8LNHENP7cN2b84KjibkugQKdxzSQLmLt13iiWHSE5nSOLJ4voxraZruGibgdn
RRigaVTuGSK88XpMMDUkEET2dAnfSEUNqx15IWUxoIFbwk8GS4uupxByClXdB68U
CgHt6zDBM9mETFflSITZVU9mwK7pj+QCQpeIRWYcIMQozM5o3YUHQMruG2EztnlQ
KxHvryPiJMJTX9RWwUvXoYO2mHVXxlL+fF/AVBVxkVmd0J5/lJq2VK6rs6ylqZh/
YSvxPONfGSBjURP30qFMw71bdinOX4XFHsiGSWfHVrbtBpzsgS6cf+zWTckCe3Rz
GMHRd3+y5Qi4l25Hbn+NaRF8YkEeCQFktcE+YG3c92JsiyHawoZlktliDNYO9SlY
rPnjwhhQfrKSfRLYkD1LdjwNs5dKFf+bD0Fkxpnyqp+o7w5E2C+rDcvpQgGo7Esk
Jn77xdKQ7l+4IShMNUtjIQTPPQhXD8yh8GlM0yG9LYJqMHuCCWciNeNOVdnlh3+j
jNYZEI65c62T8ofwHMJuZSUqCsi6ghnHXVT4m06dPLdZB6lh+t+2WevvTcQ5pfpp
1yQlyivdH3v9YV3GdVtaWzYahhtUbvwJCUcQ8UTwQ0irw1hLzTTAFVnnH5ppLv7q
1QD4jJR+wnjBBr7MA9rgLTMT49jzYYWCfQShausm3RsPpAIldUhJEYvJTBL8yZpb
HCMDAPxdNRLer/XN5/kVSPeGI91Kf+21vj1On6FhRrk687dXrBk6vo8Y1JOTa9pK
Yd3DmN1MKiynC29TZ+EIKGHipcA+dzhBJZzpobORjkFHKxukl1gkEARKg61QHrN5
8Rgl78Orei5IxqPH6sIcdtHzVfkdahJvkHb94x3SCLZ4JC2LsnR9v9Pa5fp1yV4m
Rmgz0Xd8BNZVlS/F1wRk0ixMkn9JW/F7XTffnLvzZxde6vmrQTSqMvIf2H9HTD4/
kv/tHydt3qvSG/tBpNHOW5pl0SWfzPiCEr6XvejtalaxbglCtfdxWWD5W4q8S4ju
y2lAdWkFBH63Y4l2aqgKBnm+A83cpxobeKCnLGPRVN5PJ7ojR/NPyP2sKwb7iJpM
XCQIkx0/2Qe8bv/ZmkuVjnenqnNhwvDwUy/VroTqXJJChBBCST9WYHqjkqv1qM5f
pVQnPkjTqrp7VWXtTr8QC86JhYvwJ/LWbnwUc1AYgpt60CGDdxzBckkpQqMxfNiY
IfXiXXwj5Xh8ih7PMkmJQd3x5XV2YFZDQPhZC+XHy/3/fITebrhGbtRmMNE4yEg2
Z375NA8KLo3wkbsQ6BLk1qsclPV3VkksFhYqAPVAdvBYZrlZKJvW87Uql/fQUYUE
ANEAKShrzNugMOlLcPL5Ag1KZ5lGfreM9qTpzzh7KwYYT9/8phILrknWsuSxq9at
uXdgLVjV/vpV7RH8mzlu4jKJzhLEP5U9+SVS/ChBY0Y84FZ2iKdZWglXF/AfATPD
LRiS3w/ieTYEj5A2id815i5fAh4TLX7nP2H4gnI0ilxUPlWuv/b4DxAE4FJ9/yvU
incOMGPQlf+lv9yfNu2UoL8mcFK4X1AFfqYLvlbWEeLyuiT2kzNMjWMxyUht88Pa
azbiv5pjm4C3cgjIrIOgGIpN50GyjKXfPTuG3wzFLxT0ZW7clRCgJAaC855pw5VY
dp35GpSsFvRGzHckyUOVdEY3vD0AsQtRN6Uq7vuKwxgug1FBZnOk3C6VWszvg8HK
3WTwk28zTaWNP6VDO6sprXdy/r43e989MR0ukZp/unYgHKxICW5vxk8yeMYYSVd7
CendayuVOx3SwmBt+A62tBsJUnpRsr9TNkpxD7MAUA1fXFiKmzSSnOn7JfA52ydg
7soEG0zs0MTeRarD7IZq7wc+N8yvUMxF1yQ6duo3+Wx7zSuoaeW+lvTa3dEK3vFo
AeNPgSVeOrzdEBZjK5ggNAZnC6H3r9om+OEsDtit7rRa8RVdWApmyK6ym1DkLLSJ
j+TBAjeeQbE1z9OTthq2LVyFj2TPCjOkSLnRChTpSaF1Urz0vb762E0+TJKNXbi3
dp6YiJ5WxGwEGFbFWPBbjSMwgeqZNOwjEZ6sTXIxU+5Tx6hRehnM9BMrS2EKgbcH
deCkDdJLvS2EhYmxQAR+PQ5cLFiBIUUorC2CShquIcnzAKLjabJ/E/J1hHCG9Lk1
iG8asHxjKzx+XFZky5nSTBZS7uzc3OFc6PUoyw8GpsoUuPCTIpVHYGD2HR1emrzR
rb18S0M2AMUtgIEUlkpB6nBMxrhIv7DrNM5sWueFz6xoKdootpD3O41YkbFlUxZV
KcII+hUchHZBd2+J1sTUgvGL6DELWlKZJ/n/5TTfyJQLO6U+7qnRaey2o4reeUBH
u8oMYxpqCtMaSoDKjXG5JTKvjydUEacWq0ECBiI6Qc7wxDlBhmuMbkqi3nyNS9jK
FS21quoUnocxIOsqWrVNKsgS7nWuUCiVlcDz+2gYv4Oz/Vrb3dLUDiTd7t/ksmsx
DEYyziFjN/kKCGGDp1kpyPm4sd/kB3wCxZR+sORlcaSBNPU3hx1ngATpH1WVhZly
VlVXMEY6jl6SOIul18/IdUoVxV15UeKdDWa99gEhe3vv7xbcACxPp6zzm+Q+Vm3c
IHs7qDXZEjE7g49kVc33EvUkrcTOCk8d5O0JEGUmWsqBgdGBOaPwGZYhG0qm2LU1
qtsgTiip9JvCYpoYBxEe+6k+scQqvasJnAvvHtZevXid1Ozr+yCaLnMNAnAA3MRT
2kG0Mzgy8SzXiGQDd89yFiNgXi1IBzUNG9wxjZYh1uQjr89U+UewU27Iw1hDVqH7
J5ncFc3QXcJau1sJ4CYSKVNR46oaqStvXYE7QM8ioX6V10nsBkaJdtev3PbDdWFM
TADxlPuUKWlhWuaW3ZQsvbhbu3czO6xYF/hnWUYM1Lk8RP6CKroXRv9sxdhitiM5
F/GBXEOt5S+nAzI3Ewz5yjJB9fb/pVCx6nu0FauXQEFsekF6OD/qMeG3X+COrpIj
PvUsKjkSQIV/iSzCd+D8vLrk9Yno+m9HM4l7S/6KOjhyNjdWgKH1iimPpdStsB5O
txBuBQz+FJdOBlqsoPp9NRB6K0XXO1TolIZ6vCSpK+Pv2DJBj4iOEh3MqGVQusjv
JjwSI53XgKTXv2lq65KP+dMxWSIcJ6MKHEIlXwYvNF4Tj3bXkj+7JWZqDRHC7u7r
VDdfvaKMlTto6p/CyYlujXQr6uqoJuZlm3zD/dpei3COlGLivuqwBBJ+DiJ0I8D+
OqgaV87GX7Pt7yjR19K9N5eYkceqRIB8wXvA3xIgXzg7iT36ymK+PcA2qq4DRRB0
m0zjZFM6+yDJjhOliCg/cFXv0yIVWKnQ6pVHsheo09hwGLIJ0CVdm7daPXzTiqCT
hS6TCCppYbWqilMlQwMCT22OLLQ6z6+kOZiUkqxIbWKwNkNUAi3rlyle1iGEIMM3
/TJ80xaimdzuUk7ySa5KmhVgkPN5sOs7fIZaGfZkEzGM9wUj6f1OJiyZJYFcd1QQ
m6RV5xPiIo5kvc/M1cW1FqLJ7F2T3jO0+Zz+LB/QNYAcqGQ4HxpMdxGaulaHdopM
JVXOITlSo9ojUgW9C90+4n0oEcPep8vknJN0OpBoKstALMWnL9gzjipiXeWJXp9V
Rgezik9xT28H13R4xolMsksYSd3FCvm5aWNwQpI3hvYCy31RbVm7hkeMw+rFr/s7
CMRR0quFa+heXOfeIlSHYNOcmkYhKStdbZRVV6suhkIc0pIicYBVe/gZbxNzc0S7
s7H0uis6zD+NbUcxsrYB+LZZZhRkOGG/MUzipSXrysV99TYarhfUfeySa+mxdVAl
MPLCoSL86aYq+5Dv0iy2XFAXUQEuSMcC59wwSccCaz0X9DFqKfe1ZF3rSoIaIsSX
YJ+F5044FLMyzl/igh1QZ8IpKKSoaBtjdByvG+EPN17OsYCXzxiZk+yio31kDjYw
q6mOwNBd0wFs7cPQQ3QZPC0zIQiChFA1sFlO/lDuPkUrezpAddmPmEETG9SxB+0V
QQMEbKgpqQHn0RaQobIcJXjdDDf5tG5rxh2Aommt3mW+NRO18SUvqGkVR4Z6aqRX
J8WRe27BtQwO9jDgM3LSILgPO+0965xptPteCI83PKm/QHRuBbeE7D1ctyxA6myW
FGt78zqzuVSLYoV/TMRF6ZRRzPsD3yvDMrqVQEOoRTV6zA3fonFkC6xUYTmsmFtD
C4ifj4xrOZTAst0uzgxWxBnqViKlftMJ25DJppICWGkXJltymbJ0DTKPkeLpk1oX
PR6kLtj43c59b+8gf2YcZX3G1RoHKa5/90jXEPNkRcK7t80FCa3odRVzgwha+6UC
jzIMkuiEpOHXGFDOa+NGNiBQ7ohEd6S3/KKJrhkO2RPvClnP7g/eKSQYMt6up37j
Modzj1LHdOMj3qr+tHi2KWJgOBvw6yKSjqcgANCx9gNwncfiAInEi1k3gm0M4uFw
VwRmvvB03XPDEWAkSYUmjMxjObsoMNobelmXxVuBH4gTZ6+uW13S9MVhTU2CeUXo
k+7Xzj7tbAEn2qnEMVwx9kqP1iP1Zx/9YLhlxszTpjsG5n8LNwZnReFm8tK0rRvS
XY8+ZiTkwkvCUbqtwiXIUIiExSAZ9B4TJ0NKn+xG1eKAUp90GFjrFU3JfvneJv3h
hpWYc8O8D2mYrOtqvBeE6+NH8yPG9DbCqNNtF9wi+Osj6Msn9/scqzn+scAndddT
C9x5ZIK+4ZM9rW7tAYMln5WeNAlNUFB67bkTvag2DZiJHAJZbDStUG0Alz5dqpz1
hEqS4EmqEqkZWPyJSaRkqvvc5nIYOc8pkllVY6Oy3BXwqwQfcN55BziZrWmPyTcj
xfJWLxdyn5gnllTXvjUZIYRt21wVKroleAx6l3GyhUHaVq3ZTJCOSzBh2uQZa7Gk
bg82RlJI9KQFe3Kvv58WUqhTh7lg2yCTUWtmDC7DBmZ+E8ZkrCweXygHHO802TsK
xGtUE5JpS6/8dYztZWv57JmlQT+XODAJA3cHN1l3QPyaoIo8jnijhpWDnmFdF0Bj
zHJ519pb/9N3R1u+xmOtT/YJpPLMBGtHKdpGr3kVKxeQffU4I3WgShazVIZzIvWK
nB6ptjoYwljWGah+6iRSP2QT1IoqY1CRIG/UZ3teKPqL5YTmtiL/qy3lT8dXjrO4
pZiP7hj1eyXRkTUC4E5Wi8GFXj6VtWZ49xK7z8kuZmjdqxLudnUqXNNqN9gmqShn
0mbQO+5qJioTRvALWxC7dEfeUFtzembTrmu7trKTC59DQHTJC/+6DZblaSeAd9M6
evh4sDKQHjzGlK7nyHNFMFs8PuoBnjSe04jMh7uJA96gqrcARHVQvcIZY4w+kAw5
w9GgEA2ImlyblrR13lBI8sIxp2fctuibEKn2FYbA+yk0OPc8nE6TQQ+RW7f1AsfT
Co9RLmNALxuBDpL0oDUCEcI8SAzLLEMCibNVYuFtIBXaxJA+k1ALMDYODlK2hOvj
poW+lRrFpu09iyUszC3qnprGX9Yqbbm0/NiVR8TutEkZKONw8MS4I5GPmcrpIVHN
MDVhKwVH62OhtQOL6flbjzoL5dFVWqw6XKfBm2RcYf7w5HzUsi2IeTXGZ1L9XP10
h3ADfyhd5b3WDVInVIlQetvAy3617fElVYSH0ffcLVb3YcdipXYSBc4HMbMkqeVw
TRblPivMq6mU74OgjPmbmi+s3wqIXdFg0TFOZneEfNdCiVHFBgw5AO/cyn2zEYtS
JfomF+TznuHWkj70AuybFw19MGIvDuXV9LesHVPcQUr3qGd7z+GSnXmW5euyKBYu
60m/mt7c5Ryw0TgtqNVdRXtO0kjNt5Yt8C1awnQKzkAYw82/rv/LMgsJu3lu820d
RFY66HszMksPd1BA97P3nuSyP9KQRwqUnowWyzp2PFw5fGwr9IVQJJEt0oxyMLvl
d/zNyUnNNYjS/m7dbaks9peM5tZ/7knG+vPw3aYvqy7zqcaNoom0ohx/StpH/QHP
tqGplh9aHXx/kKD7F28wyTV2Y3Lywmb4nzdpYELDAy67pzEw/jwQwEGlbF2QDHcJ
HuhA5IVOUXtTnVhBbChTIKPIPu9OAnXYzkLV7SuofyFBOquTaeAE152TdgsO7WtJ
la9uiu8szcap7jDXtmg1WuFfhHTpPVQLPcfx2MantAY2e2X5VWKqbvQdlBxDIuS9
qTxGFsxzJaizypKR0/vaY3BM6V9vOTr2tVUeYczVy0ZQf/ZecjiWOF8jXauOjpOX
Psot+L0xrcDDctJM1b2HgLjXL7jn3KgXcOF1CqpF7NWjmDtrEf9y8tWiK3ijnZim
1B84lEUxKsvjb0JIzlFs3jQOhls1nScDQ0gwrUOEdY2KeI26fivRovj5bSM7TTl2
5h34ut1GWoaxFLWlq5c/acfLtQN6z5+LkCM+ngQCpMKqvIwdrMvHDJBVTPrETqVi
bJmQzQDouBqu92F9ItXGv5oMSWL7BPyf256wSFLHtmZOq2Tsjw2MMX94NknEH/4v
uaoCrDAMJPaDHsLrV0PB9XEfx0GSBDVod/dl6ew0k3QeibpBGsBrqR9WqgEM0qqy
ebgfcK3/czmtXLP7pJyw8d8VG/y+ywGLNC8KjV66AyRsN2fSEue3Dk5LrnRjPhIC
a3NKuYo+x6yfWiskpFZ4YLyXgz6pMuD8UZaCu7Hn08JWk0L9ivxR0Mn4TWozAqU/
sOprL4NESB1hmEsweUZQJcb7157PGqZNYZ1NTlMRFW/WLUn/Ao4Htrh/K6jZ7oGP
vUTwmZuSKxWNcTxvt2u4w9DPTGlmKs9fSJ8GKJR9WhjmdoDalobH4b5j+k4bdywZ
y6GXsgmeBIOiHEh/tCLTSE0yJeYQcO1Vy3kSbA3YWupUsa6P4xX4zqUL8TXc5MGa
A9l70CcgcTZwrbBEBck/8A4/zTG8fUKX//bq6QzFDGjb/8XJgdkewrTSXXs+uGIs
ag7drIJwNg8yZhgWF2Q/SFEAp33nLb+IorI397CtPBlmcBlDCHEVKpJmey0l/nsh
Z/rZS/ZAFVhXmY1odtsrXPk2+abVWXYVMvGk7XxxOzgTHuRbHlOnT29aS/M6tUK5
/cLj5sfpgoZfFk+HVtzPlAoB0VfLp1t1hdcH1NoEJYiDiveIuN22TRdSBjAgq3jU
CGUMh+ndKHaxd/Ie/e3b8SbfPJyy1cQS8VqAumJp53a7ucBO4LvSMg8PuuIYqJaw
J5h+3yN4OeuA8UBrfzd4fc4X8e2jMStVFi25ELcOf4xSpIM6cGORYXoh8ekPbRxk
UR8SAccfZsED8VhFgFC3zIOUjomX4BuASaVg3TIiFgGM8tpqoDDA/Avb3OuyxO2V
V0bMwOdqQ+0oCLP4ZLWLeCFrzxbVf595A4SZH12iJo4bT1C6XwpJppL6MpQ8pFjR
+zN3izbL8DfOQB/SsByHLUoWD1PRNJVnz3wA9ETzaZEjYIET2vl+cGqjqsn7F2nj
552W9opx+4eQnlX0EqSqEXEJGAXPI15YufS5R8F72gF9I+eozHylK9wlQFeFO89e
RmLMasoluho6BWC8t7+WKaD6PSgGmUCwe4Qko8HAUNloJ1BtS6aavzagWxoIJr8v
SnTD3ofzB7U6aSUTt/S5aQwKfD5kZLb7qJR5QIr2knr9h+cJ8mOECDBnS8wE+Jg5
fME6C68uZjmwWFHoL+k3cRtZv72sjMWhLUTcDxogOdp55mvOKjBs9oGFmrVrzHAH
356YOv0mUyiITykmQNuBQMlYzKXLjLYA8+mcxh2ojShaPZbrwRNQn9IFjK3GjdJ+
IcGucwAf25EBzabXx8gNSO27bRYOFQL6w5qOj9MHucJ8dotq/+XBkVV/AuWTdIif
staji+Qos4Q7CjAkqbm+il2Li9EXQFhJROtapeA4ksdE9Q529bxnHkiDg9PU5HYn
aSWnIUcBUQxTo6nYLQ+ZfbqCTLfXXPcslwKpLZPFqavA7ua+OdNfGbwCfjt9p2UR
8ZC0edt+l9AD2PFhyv5SLeNx/6THcRnpdMYG5of1mJiNx96jWZ/QG/mCLzzL8OFL
8zeOEjg/gvvFTtLobfBqv4hfDC5jP73JbMku1MST0AH9zUArV5SUH0zs1O0pxBEK
nS31hR+5RXqkIvf4Vq2UEyd0ahR3uHksxHHxcuAp0dCIAVxKgH/PRSbs3C/O5pQK
QBhItvicn1jRdBeqfSkL9t2FUVU768c1Un0pwQqgacgATHWfg64H1fs1vxJ2yYgF
VZpvFhMSkio3bh7CCZqjlOMwcZKzYJTbpISfLqws2wjplvnUmqJYZFz2gg9bsXJz
GLg51SvmajsUJCWvyqVR8tFKDEmkUrkonBy2d2TKVMSY5jRAoCyy19DpKFBVnkNv
AHNyDzKmtTE6+XMa9Sy235iK7eNkDLBVOJa93o5q8k7AvgAc1hDxydKrXsha/OJ0
VaKmerooMxRGLuD8ZmLn3igDm/leeWWobaOaoN0rkFIG42yLFOVnPjLklUU9vqwr
k+K0YwBchb3Up8nG/AaIDzwexFfKwGRhGxzobiJNE6NCBl6mEC5VGMvyHOwi1jBj
d83QSJjgErHRtIBsBnJI+NYfGWnl/ZEo9/GMY48KQocfOU2/iPsy0EAAG+W0aEiw
GrZDk5BO2CVfX+c3EpELPgYb5EfJw60N9tXvepNe/IoihGP4xldFDEiQrInaIp5N
aj2CjyE4alOV4iEIItR3CytXSGA7YEZ46L2IZB6jsyK23qSu8XlewxWyMdtdS/ZE
Y0XCCOVsC6YV8EWU1aNknXCT6ZwuP+JUeIa1LI6oES8j8Xwd71d6As8aqKCYwkp4
qLL5Em8nf2oZL66DUCP9spTvk3iueH3wty3S56SSIFzbTt573St3OD4oeKa3NEYq
1tEuIcs8aX/o7zhe2tSFnHxyoWh6UQcqIGp/UhyJnTQD2WvGeGoKOcL33fMTKM9n
oNUd44evEUzTG248RPd8dMNi+wdDZkwjwaiLDASbbP5fwSBqnnvTrdQcxVW91f/f
9xdbfTf/64MvSsnkISQNB50TS0wTHkAgRd/X5qrGTcfnh5FBkx8L9nIvNlJCt+KH
brMXq+Lej6P8gm+KkxHGd5Yr50jT1FWKUKfAHyHwsC4TDpenXgkMRnLphwWUdBly
U6asp3huwfoP/HYEiQy4C6pDbcMN8g7jwT9Z6vNffcJ3fLOmuFG/d3rFj4MS5xP/
IGinSfPpSCrP9X5Co9MQagyvXTidqmpfchb0EVHy4eiE1TAPnu2bFbhT5ccS/OT7
LqAMNpxKhVmFQwNDAuw+ztjNoLZ5l4gz87fXkMO3CmOGusq+d2Ih5PLxiDBuxsl5
9zhRvLB37EX+4MC3SedxleeaCi8U+1DdeDYrOhRUzF/5VXdN+Nk9Pj7HCdS5ga1I
vHv+2RCzS8CiHVv/iKZaeK9Kx1yZ6Z/EUkr+ZqjK4io7YiiramVlDaB2hAP8PIcb
/Wo9ORGtcjsoYxIA+NsaKNGaijGx897tWOgAIJ1oABwYRjvTX74Liap4sSAQVNjo
sPIyDIPx30PawH5MR/mS70HQJ1K/qSJqSBJUow8nEpnr4WWNvaNlacxFmYYsCLq2
uxbuqRioNNm/wQVWjQPaUxp5fydRcFAe6ExlpnzzJtbPzMOdT3AUJL9GVozXAtIH
hSff8RVZKhz+LO8BbgPdK6YbwcNxuUNRheg0H2m5VSRj032Ur3qzzhHQp3FsbL4k
oi5Ri4vMCQNd+NfoAW/VEP+5wLnzaS70FyT7x/wIoU4Y39vzdajz8AcZxgAx+Ff2
l2O1xbxJXb1zViuSznkmLAZixw102RbxP9gfNq849kVe+oG3BIVbIBiFMvev91cx
79QPQAv65+zdM3S1nLuXg1s19ti+j+tt41iSWVFn5MYwUK4mACp3YdTZPDAntDW/
pOsaEiVjKbsr6C2J2o6SgRGtIxz0mO0ABZmW74LuSacFmdL71yLOvTWnY4J56NCY
MLbhuJzbfo94DsPMRkZSNkmWnCfxHHo/xmOlZmKdLE4NBha+6S+zTEwNAXV769yG
hQ/KxLEsXyBANZzky02zlzntUCdAfmxgxJcXfIVswh4OL6XOrQesvB+Ob7KXWg/U
8+l40Pjqrbk3imD1KuyWJkxCeW389hMDdnA0niZYMbrWh5fZzzsfJNGJHiZu/THy
I4L5tsvM7bWxBqjVHmHMlQDunervZeblJAsjPBCcWhbIDf7gRi6xcG3q7LowFrh7
D6tHFjCOMxsoYNN1KXWRJXh7kJVdVhVF11LHtnalPKRCzRi/rTDGtT4Ue+fB1Pr3
kIgkol/vXpKWJGCZej4yon3+C8F04RX0BuvaLma/l+I5f08ozo3c6TrAnG8HfZwE
NpLEdqKVzaShm42oOnI4DQicS6tXcHSSxvMVO4xjpfMaNu4D7DxTaD8Yuib4E/0G
RIyn3u3jf5A1Lx6qTtHtaMl8T9kSofabe7Ffd/D6i0aHct5i+Lc0SQkc4jX2CZGU
KRTemQB5ckowSL4h9uLJWohkwqkn1kbnieDNdxPFSORFhSlIMsWQEJLvjrXdX3Fc
w5y2FTfWv2gbHQ24pUc4nYUpxKiNUoZvSLlUrNenY0MkvJFFzfSgmZS89EWzCkFY
chuhNyV4u7J/HAXiRH9wFwx1xHK1pJNXfSh1HeCz1HLrCVsW7WA2kAFUEUmxErs5
PUsPLHVDadj0/pWchqtjKRCynr28O+BeWrh/2bFqMUPKbdgx9Z4ZYjudrELOKu/Y
HGYHbpy1D1uk2cIsu/wmqeMuQJZCkWkZ8uoJKecqfFaVmxEEow6wiYSPMPuOiRuu
7+QDPBwkrZwpDyC1+Edtfokcp9ale+WsPzTUZlA7AhvB92clDCEHCTYF7uZ+ySTm
etBe+frEE2UG61vLqWens4/iFLvfo2u7JN5TBh6vWViOBfz/geP/2VRhGc6nZ5Nd
0rYzhGstY77j6Nhj4hNkU5RNvX84eERbpOulrCFUyqGRI+b7OaWXFSL7wkE2Fr3S
C6qjgAkHiSxwKhsCK8EEWWKozuuhB4nuJaoA1eFzDytkdsdbCiM3NLzknpw6kyLI
RNUs3WkIdl5AdDkCBGUZdgUv6MkBEEaMAGBmWmtlZ2az18Wi63A/XsiJDwdSozmk
prpJe5Ov3BdmO8HvTEn4uGDR3qQnr0P1Z4xY0LOGr47Su09SmGCgjV5kHjpKC9l/
XMRnHKbtdHmPFZySQFapGJEQ2roTy1hlSXBCeRYR9rx1O+tteChdqqLDJeB4fRUT
16Tv+X4layep8oYWgsIDGBQOG7jlNsCIE7ro6ByuJ9zxPglPLAK4+rtjMrAWcU7V
59z+0O/uT5OHGd1FuAQdyruxQhZOyGLlH80OYqdlw6wRyeKXb6eWUiiu9kaJhNw6
dSDYLVXcKHP2dmGszmryIJ8/8Ht03H4oedkkTGLW7K2a2zUUcyOddkaOoMerNX8F
jGw5A3hoeSRWmBVxFApR5f/97qlj+neQ4n4o8qO39rBXJsX9EB8uJ+fEh8k8IhPu
B9BCqhQTMlbKiMN1+5aXY30z9atoEJQWu0JcL3unhRBpMPkSaTXw8oHoxF04vpRo
5s62H2iYtDiwIF2IWscoBmmhhwfp6XSaPeo4b8YItzGUYnKj82/ZReJQ4P/L/pdR
9SPucaqJ34ItGxwnld43+Rcfuj8kjidiM0Ep3OnyvjyDwVSip/NXAWWvAMxkYTfs
/Y85XvysfjdhoTaIbe96PIl6YocUiZFWDwtQ59NpijZVV4qvN9O+cdMLIMzQcz5W
ZImywFVEvfmsUjFvwPz7QMTlLOJp1HFCvnVH8bU1XePd2K8vvbpadfBocJA55rdE
26PKjzqLPX+Z3n01btoLtDxNKb4tUX7etZbutv0q0ryImUxIGYDwCrV2tqmhV9pK
OckAzv8vdJr2oH4xExFLuJ+wOo1EW8A3PGso8sHOej/Y0uLaCGRLCGjYgs3gmE1J
4n5CbK3vA7heatJ4TSHBZnSbZ2Z5m/vn1FIWbLqKQ7CIJ7Eoj0iU7zX0f9pzr2xg
hJxATqd9BWbJEoLJS3XeMG02FaB/1Hs3Ar3sz+a6O2G8U4VqY3uwyrMnUHWirhm3
k/u3rAumnNYW8R+tZ7N4yaMeO9z+jHZTBpSvVHaSJK+ny1g8Aarv09LVWrwzq59X
chWNHaAqEnd6MgOJ9zFB2jirGNoW5sJdgsBmNqDH/i8BuOJJ1KSQDgWktQ3PgtG3
PtS8NikzvSUOau1i54UvxwPrZ45wvov1g7yg2fxflhLc87qCIGwCmTH3lUm31tuq
7trXtqnlv1vpfRcTcTHt8534A3Hp2da53BLgzPgFSbpk8oXEAIwLIyKqLftxS6xl
fAJDw95thY0Nk6W7N5tL2XODVFd0b6W3QlCX102Lhnbuv358LMGTdf4/xslzfk7F
B6ToZmRbU7a4/z3AdS+H86sFrmTRuLoF8wszdlybbQ2wNL+ZL0NWJ8negfN41v9e
FJcT/YXqK2Q80n4aVMisfUqzDsgMMj9ircbBvwMlyJ3flZL+xtciMaQlDYgYhj74
0JzCzs7vERSXHKIbFFDOsWigVxFpbK97BIJH0X5pe+xaHIAI214dOvy+LY/gefwf
IXKQBKO9UPDFrTgkxWOiQZdwH1BotXqE3hS83LCajT3+OORfAzhxeF4Qx2w3OUCx
M3sXBpMRbQvK2pScrf5HPIL4j5RIyLdI9trsWZYN9i6AnQEnR4TEUbdS4rkZjqqi
85COIzKEhvHyiH03/U3PJG7yABRpzF9Ea+6hxYthWuUxvcbFAV8MmduM1t6n/gWr
o6l6ZzhfpeoRnRCmKfYrUhRw41AHSQbDLzr8WpktqeCBk3R788Y9zQ/UP7HP4onp
oMmXZDO4+uaVHoiJgx+loMPR1vk9KtpKBzZyq4+DPN4Zb1umrX5c3IapNp2HXgY5
4PnBYVtfuuz7ErRlRsGJ4yPAOTY0tRsLmwBA8iwDZN7Q1tuNlg2G78tAK+J34VrD
q5w7Lt0gO8SCpg7GLw3y7Q0NYe02NC6q5l9vMdxb/ULqbbxtRGfd+RX9Y9EKWgUZ
7SFLOusdCN5KZ2Da5nSg7YDXNn6LY+pXeeeZyaQNCTGSGVD84aepbtungatIaBkg
chuU9KEmhtKm++qrIuf2PVWkuIZMUYuLxTBYFxKbxNZ9blcKc8n2oV2gREnA5xz7
KMWDKfwqNIJJB6R6U6DACeLxltoMRQnYiDMaaF0P87GHZw+PZi4BY6eWGlrsh5B2
W2voiaukbSxtSQk9y0SGB9qejel/IbbZH8D9AUVa2qqfdx0hw7qLrdWXzSGT/eeI
Un3S6FHQl/Yhfi0AUQAZB937Qh4G5OcVW+dUxTUojDjv9GBQLf0ONSJAZYAE9elD
9gGQZrW+rlXxmGaByG2TIWP5P3Kqmhl4GNcT/Ux3lf6XYGCtdPyO740/UbxcBu+H
WzsNgGz9OxySLvXOLpF2twQPKsqOa7qU3EIZiEfeX2a1wtg4JALI6RE1OdoS/RJ7
Vjkv9AGMB/0Uc8itOX5aMWjIiUJC27hk8Lai9+cW4esWu2+t40E6K668QrT4YOYE
awRNUeR0ZYcVrpE3nb7leexsqNeWpC9TPugRZcPmst2E8hb9DoZTko6xVgZPviS2
+Bg0+v260PGUoSuKKf5AJLHUM4aVPEui79iCY3qiph9gM8pta5lWJU/LIXUF9Qdt
NJNDysa0oBOx2u+J2h7SQVgzCoB6WZ2JVQQJfCvn/Jz/M2spOJ/GFDV9rojgT7nc
0b63UQBhbyjrHl8WALTMOx9qnYfQ8N1v+iOpV1r5NfRNZXUTEiuEGZ0y2D3xDzG2
R/V6wE/Nu+x/IHkbcngSocYg908+V6r2X1yb+xDNCMu41N6XCP0kOLUKVs4Wc+RF
nctZuO8WWLJ+dFvwwwaQfsihZe71RUFYcdCDirSycHeUJIN1aB5djlaOe544+shF
KIgYPfEYPpoq0ymI7j9xn0YpGshhB/ovoHPyO3zYHhEMaOxz+MmXejKMhWo7p1F3
eoQ4cYcfqwyZptuE0nw8NK1HWlPIGJSuBZmyZNpfK1f0B68Nx/a/PfxEL+ZdkJKQ
sNxa7Diol0jTp3/lG4GleOwBHbRCEQAwv34Rx3Y/1B1R3blHR/VfPL7uVg/IXNAp
lTe5CCuift5TzBqarPBq9ItsaYq4GsGpyz5786DOmnF5uAbmXFi6UrE21RgiyxrZ
Fc5uPXpEJMCmRwBTa4ostE8e2tYI9nEKYsGkOL+7SyParvsNKnI8PJXNQemfUWre
oYdUV085+IoN7GnQUYma52z3kpahsW2xytzD4omjP3iXdXvdfYPcD5C1BYzi2o9E
WNJLMO2wE6OWk915DXAAbaFAMSy7x3dISRvmK69E7WjpOgNAth/4QFZsYrNEVyFY
/QzBXncTUBaNJ3IYQvvYw1mg/HemlXkKPZm8HEZ7gK6kc4B1KPf2ed2qljN79gH2
li80gySe6OiwMarMAtK2mfNGWn0bu0vRxNmG3GmOz05IDylSvk0x8yBFJ8qah80z
VrkDZ2/zWfNamvtw3foN+KMdUpWRp42mWhxlx33WFrxImNl4plS1w+H0DebgsMIy
aK6e2ZNYjAuhsGA0TPdX8cIWFpO83/bh6vN/OYjSYMFzlHYWteHp60YL1FnuuHNp
3fOLuzkIdmKP7KhSDm6afeAh24fb6PKcjBL9Yc72eaCl2E7bpx6ne2AsBgdi+7Tl
zB/OgimKuMLNhb2XozEKPNJsY8+Cf7+GNnPqcIY03h6IL8hxkPtDWWPt9Wb6AcZF
qX2SV5/61EL4TXNeoebB3qZxJcVB27r9OTQ2EMe/I0ZZ5al1AarynpsL/FeUR0T5
SG5l6Pb749+kguHZitJ56J+QyKCSgTUso++sqJrr6c4vgi/8RJUMkWmGleus3D2C
fWdNrTb4DBLnF9L3JRmkG2C0WdZDLiuXQQi05cbqj5Wn2Q/zkNFJxPdzF3kzRMCK
EmiTT5p7RzWycDMNmgv2pClQ+byYAYcIBKXp2vo9Ga8kSs6fBhShXH8kyUHf2UhZ
xD31ZRfYols1rOsOt1jezTQC3FPOLpStBuSCMnOCRocrf5F59ko9a/76BmaPEMk/
jbG+PXYmxnJroXO+R8+ml316pQ0+cgqy3zgN9UvqKeBSoCaka8CFZsYrinCPKzJs
8Nh5mdoVLYcSo2KEnnT5W+sjNukoCC6x+BxKt7UeJcYWYk7M6IjfyiyHzfVRZzOx
cZCCpt3py+OREBYQL8uTFXaicaKivNhBHY3zwljIQ/CttA/gyrORKM4wLE+kJK+G
9BvFO1Xv5mS/Avh5OCi1jf73LobqdJULV3k389Hx19jWaXtBkCy8V7iigtiC/qKL
8BKKzC+RJk5ql/3+S3s4DYy+Fu+Bf5OmnLTs6GST0AAPxG69hQev3sSP6CJWn1h/
i0f1fzfl8O1q+cDiAO7hrO/bmiurKuNUWFQoTAewiDjX+O00ti3Q7HXilD39yvE8
lwzOESuNYyFhjGVk2TvkHBJded8Q5Kjw+an6c9nB2IWKMlnCDm978qdeXiJrHLks
vksiv9qdRIGy1Kkew3H7F+pSx1lvaiI15/c12YAeDYZKe/TU+8YdpAomszjIIESO
l9GSefjCOSbD+DieJz/ARCqgCWbsmqhsStOLo1Qup22sCL2dvOy3IdFcxD4D27IC
xVYeqjtqcFd3Dh+phT1ByHBlHKkh76PJzfnTsx7jpRWqczD27yroAu4TIHKqMSc3
7d4dEe7bsMBlcuccGRnxplsCIrJ3kkdXuqywPLfJSTGB+TlqX6cTNvs95/Yb7K1p
RRgdAGat20N4Vnj8buCjQJaOdscifTV2pV3o56Qgjjk8AVpi2TdUyPltkuOaRVRv
bf5d0GJC57/TTlGOnkWdaXk8oIJo3dbZf6hSCPsHAslxKSn7P+yVLHV2bBN7WG+7
NtIpfCWxSn+CIblWefDtzoDhe12rJJEMnYGxiFQgYzbF0JATWH3Xo1loFNcBvgie
h5ACjkiIpmS9MMyS9ex57PEF45KW/mmbovvWoZfGofYQUcqy9eVAfaZDw245Wfxd
LKXh29KXZutQ2Xx47rl4c6HGb62neb/fiQ13OGY9XO9OSCtmw5kmpO+s9vNUKaIu
t6Yn9BwFWyU9WouJ702t5tDCXUcaU5eQL4i3/5p6kjhNkKNLgCfbfGJpmZWJnEfP
v9X98WKveo2kCCwSRZmpQm7bimG9zMr+cKNNzqTadUyEqIoQFg7KjJQcqXQeGFNr
UknywHfI1nf5hunkEYJ3Z3adGPMRJtRJn4yJzGCSgkakbFT8CfdaHv0elELxhSPA
hUnBggfnFugw/rXA+VbvJc/YC6LbKm30GvBzOcNa9oGuk38h+6fZhmoVaKZH1OWS
QtO8EMj3SSPRHjSNevphBfknzPjvUnRfpbdi96jFcf3hW3FeBwqbNCcW2ufLt3GC
g13lV66ovHQahKE/KxJ6Pl18KHQk6Q+15ymxWuUYDmTCCFSxqc8rN1gOyK1KzIQT
O7nL8iQcmANFeF31uQsRYRdgsx1uDH2haTmYe4phqTBVpCXq3btRq7ax8Ov9BGDC
7/JSt9wewbGDHUDkP4KtmxH425YJn8x/3AejqZYjz+ZsuqJGRCGUqwEgR0mA6dXY
o/6aVRgOQdKtfXKYkKjDzq6Qyen5Nl0Q4G8JLI16CxAFpnHOM6foWUZ7boj797lE
ozdVzdUaq9/PTuNwp8FiTZAqdRemmMud+QF9PKlFmM8ivNPmhg9DUmWP/q6OJ7c7
ezhaxe4amdkVhw+8f6gwKG/EktjJVbpl5OoFJrternEdwtEhzpx98L/LuEhVtO3V
BgCJiGhU4n8wBO5CJYyXp+1hCWUT0qEm0b2UeVqhggOQcUmMHse8Ek4KjXW+ztW6
1AMyt6upLr5fWYuMAphdZuN5yLbj8/6M4xQhmvbwaqJzBC87WPwlbrTikm0N/NHW
L7bOlhZuEOHqSWcSV2KCw8wGhWFSAgXrngU/wsLji6mqby9zrpYd8PjAjc3j5mIk
75IrGqj3WxoAIaAgVjZ7hlG5sj0ndT0uIk/vWnAKp7vZz6XofmwcoCvjVBWMQY6T
rzS8bQR91MQXqTYDKMHMT4cjM+aKtrtNjlp8ewt4LowpV5fEal1V3iyoQwTIUhMo
qXX3wQt3fEUa0LoUrhxX0JMG7TFlDt4JrAwCen2yndEm9zQ/6mSV3MRysamSHpLh
sjcAlNZNFngIVQra5wN7BAJFk6A9rE6RJsHhDfF4dN/fPCdn2Tw61RfdMRuES9sO
utv76WyU5uQmfgy+xSoWsksgxEMm9NcVubTUJ0OeZ5VcSm4abcx7E1vgefWhQpY5
GuhF4ZOdUZDEf+cdE93zBBbRxHBVsgjSdhs1utcoEeUgOmLHLFHkuRqxYVseAkfD
gpJXpoRBUY/o05dyajeNLbBgn847on6U2xXqaUQw+Br8fdOeKDpao2BG+MmWhwOW
mkvoJcXETGBOTLbT5xMZ47nArv0sju5feWhq5YzgU7UK91JdcRPnbZ47w02Ppy9F
lwDYRtFJbsG1T8hlWh0HPee54RU46E2j7CBoUjmb06zk+PuaDaq4osQAGaWzwHRT
IALxtAfKtBVi58q2jaZYMK4SMgyfZ3/GEOP7LylA/U8i8tOKdcjSPYYlNRvXUFHr
QuwdWLfpVwWniYJPwsdGRuJvdKYDzaV5U6kwH404+OnLJbtSasXVRfAKjeOOVu6f
88M9cF/N7pSxr0yR7dUw9COkZIyQXC0YiI6I0Nn0YUcqRaDHFf6pPA4VSmKymKwW
3mYQvrR/B/9+fozswgOaRTvaD5qLkXpdsWXO3DNOyr7VHNNvpc6UKyieAsmJb65X
wJNEgMT8z7VO2RZftdLmHnUsUVqFDH/jnzCrFX2jMvPy+/4fNQphBuflwsPyaAT/
+znUUD54MfdFwJcQNmQcxfZUsUPcUn2tthmDL9VQxL4eteEcAzdwhRXLRmia7Nmk
j/VRUd5FYILEjPnM8l7X3sKm/rgRTfPErIKPqdFFQtNDewHX5H1SGpsbJHZKtF01
x8QttFZfGly4vDOey927RGM66YYg7RofZ5R3+XDeypCA3p/ykWTsdoKE52XUE1sH
PnZxx/GlB7bZbHJbql9fugFA1szI5dOroFbCRL62W1YMVfsjTytxnqX74YpieTZ5
bXo6V/L+1L1HoZ32hDOed4fhBXh8EcZOMPV2H0jQuEKIJQ2y3hrvMeOBFXxK5YyH
vRXAeXofD4iadJl8Y7nsGCQCK2tlFsifqBma+Jpdey113zp1cLgkL3TSO6LXdsGm
JSFlLO8v+kHJCx65A9obO7gN4HzVC0UGkgB8lrJ2bIPwtACWADhJLZ9noaLUi86W
/iYemumjp7UMB56huLzWyk7ofQM794CTxs5NoEyYWujQLPy0QWLoyprWzxbxhbYN
tuMu5sx1kTgalHnOyxCfPr8tn3Z5JyBdACDWq6fYkG3Fy7AcPvU/5Svn40+hbtJ8
3Om3TWGm8BCrSkmjj5KMhIac1b7foLZd5aP+DQ1Qd3JdznbsYlWRgVmdu4SBFfkj
WDj4w678cOJFOr7IsrKzMsv6uQ0c+qBge4Q35T1HdqL5P9I4/oh2G1G9JosrFssT
UnnL1kyeth/qgbAZLaEOLJCyv8MT4smyGc141787SC1hixB9yecGdIf1RXFNQ8Ln
4GbmhcrlSqxQcx/dU9n1oJnM1uJcletkkU6frQPc9b5HGCuLzDuOPicn6z6P0DRF
I01dPi1VGVZuLIJEtU9i4djx+RsIyyFO9lOCv88ZY2Ssrt2H0kWFPlJvg50ipNTU
OJPB1iUCvuwIhJ0xvyTXgC5bZHr50eF7gum8bqDL+hIaqsVkvg/tceev+iaO4pnR
9bqlm3IrL0IVF8UIjoynU0Ynd0+WKPU1VUMwXWZOOt7ZS64k4NGm4Bnm0tqbx81L
zpJYEBb7yVrDQD9MGcKpg21zzsUQtAlN/skgUPcGd3szA2ywBi1i0rfbkmDE3M8e
AvwOhEAIICIRgATF4p1HQ4DvrEO8UXWVbWEEXpddENXiRhCQYi5dafR8vkAaPCIJ
tGnd45XzvF+xMM5amF7TIWMEe8dbMbNrbfz0eGXkG9dlYvHSo2T4lpa/zvAi7a3f
chKHqsr4QZXKdZmovn8APXhHYd5s+yps7FWd1idJFkmHpCEmNjIoSWsVwjPIe7dp
jO9ps0Tv+wuzZxcK0p5GMLRCzeCADHl5IcBg5DXC+mDSEMIVTviYh083xNJnql+v
/ZWQBFYHwTgYBhYuzrrn3dxbz1xFTX1qjQGge9lqevCwNbYVLYLw4Mo49yXDjG8M
54hLsdAMHDaCaDz6Zn8Opcfr+DceiDHVmhUkjH3dBmENV7ljTxIw56Cd52w70KUc
Uj9bHsfJ2PwhsVCl3suTc48kCgTj5MN2ISR1caxND7Z/8PXKJxoSVs/2ryYklNvF
wEMsxI/Q/Gxn3ZTCBw1ThjtYLle8MsQ7kpq3lsdFARJaPs61tEpgS5v5yvC17s5V
hXuV3XosExuEogudNMloLgR96haGVQmhMj+c72QIKMY8yLFIkpRgK0xx3OWaT1XO
hHTmZUojGPF+5BAZkjptkza3Q7fXpXomJDF2d0HUb1gaWkAWvqcD3rjipkFi9ctJ
lnk8C5TT7/KeDnfpyavoOK//7B7tjkUvmrpZFQLX5RODu+YZk7HS+PP58erIpuDQ
m+p6pr2AXcj9pRT1PGqqGtFUbrlLpGS8IP4NCcWbT8yM/3xioAEs+AQtqk4/wEot
0dl4cibgfPZ+R0t5/Tqx7GIndUtA2gP0OKh9hHyjtdDDp5mcaY5t6dlkkwZ+GEcT
jjsXQhoeqrnaKCghVImWsLG46UbJAJow0Z8Rv2zG+9hqIv99pqt2AHrNW00Y+2Pk
KiPs+jf505kotPeEFWSaqCBp5GzydcndS++0zaBqLk587F9cGPeJLy7lfoLZ6ZS9
2dAB/xGYItTYyCZPQJZCo4M3ypcnLraWWFN9U7zpgyXYj9pq0EPQVPmBgoJYDxUS
/na5CeNXeZgXhaYpvW0hH/zB1VEqO49b07fA6zEBtNpN7a7lGzcuuhdkEgqcj1La
j9zDfBSyhDGla53h9KTKN4TMvTO+TSPDdtOnTsuGWVEyiKSnXeAtN0yEvCwvH8f3
xSXZDTb5XzyLxZm0QGIbKI3U8Vj62quVSp3iURGZDAW0OCjGzYTRRMQH9ITf+f7O
FcNHJyfrGxq4fjdZs4zSstdi5oNUaDbTzzGD0RFG00ROlXJnzRvwnOwUASt37qV+
hMZxYFGKZb02LSCU2dChEsUbBSh1m4HmpbazGMHCIcqqwpqwZECsrVKi7UkMf4hj
Rbyim4ZbdmeEyv5UKurvr1S9FeMO3UVYOmyWzjLvpkxG6BgnbJgdaDXfygUUe/lI
hm28zxqUpxAGxICEwJhfvfDkHUItwcmzQTGekuNHAazMHHjtpnH5XIKdRsDBESGw
ieX8HV9yJ0yxFPB5GVnpsFqL1pEE0HuXnBdn3NVHKtQlx3VQg5ljLFsnT7jkr6Mf
sjFmjr0dNfh9VD+UX1VFsEGzl4B1XQXxPeRVNY+gnWIdydQL69LzOwG2YkTh0IJh
8Cs8MKdgQ3cXo/ATs5nI/xiSOKeSwUuwE3NAyNk//e/RQjl3dlOH3RT62IyYibYI
LTswA966uwErh/HsekcgRazSxAvD/ylcjP2LXOJIlTpOjBsOVcsnedkzeXQTdXaT
02jKlR8cIYppBvdrVQv4FkjoPZ+4L/jHk3U0F6PW+tnwozROj/yBOMjXdFMPQlVO
xflG0TjJIgSfZDGrMS4eCEHdlT2ysJDAWB8R3UBs4ZaLdt052+YJxD2dBmCkP+++
Pr02Lwl4mPP8K6GnJqqdacdlYkyR/OW9mNY8X6VSirYV6mOyR6qHAhQoUX/g5v6B
HJVvKH4RRG5sOlneb6O7HxeUnNZqtTy24atCLRFVNL9Ka9xi/2wSyP1aR/Qh8PlP
ioyaU00w2xYJCDHU5dZcwXeo4f5PkR4HNlwIYoNHgNmYTJZpPe3iwzrO7Pr9VXTa
pfKqy8xajGZYoUJn1s4zwABcd6UkLXGLmilJUyCIQe96tYWX3G8r7sLkfilSdVKH
s8fm2asBLCOCl0SvZSV9+2fTytPjEe/XNg2fh5fIWbX1hwNCKmTePZr2KyIXTj6i
aKQgbteh6iEtdnm2NIu4y4bMWe0Q5pehsDRkVjgceGfVL1fF9UbC4KAUd16j2YEN
dS19QxCzDC+rhWjx0L5vOf9JUpv2jZuIEzLNmaAE7qSSfwiIq9pqxfQf7zEpp8uL
Bf6i65dFgaWDjP1ml6EL1697ziYQK9YEEV10bUUw3SZ1NzW1Byzv+ekR5f8zwKpN
GH/FAlar1oowOshaTi5VZF/4NnJh3D+QMIOhfb2p2CyTbAws7FgeUKNvFkDFqVgF
IQ673Po6JBt90z7sWxwLpzIfwTrK08+K9cM1QOiMbAZfftqcqqUvieAKaQLacRyh
XTIy1trqQQTcDkSo/B3h0QMLfaF6n3g7yw3hKjnuRblQMrx3gnuW7sgRJyyS32lu
+fAQ8e4DthzHFF6+zFTzs5/tfQNhCkUrYFAn63ZxKxFLvNHir3WMpO6ZiL2yf7Xz
uSJPD2Arfi0F5QBWco44omOQE1erqQ3ORb3X//kFvd7aqJgwI7h79Zn1JJiC28N+
ma2px/R3LKmlMqGrWdomR20EaNwpCju/EfN6Iov91uwZ4VqGmvED9sr6OhPX+eVy
JNGUNsTmEpDIQiicS7ksDHY+M79rv0I095f1uQSq+Y1KD0qKUFsjBCLEfPLusNUo
l3jMr7hYxjFQseAPBs6X2MhWX7eq+MrYRnchWj2jkDY6KQLFarEeLvrRN+1ikQhp
awv9+LeJr3YjJW6UZzB+OqGzXHjki86mFZnyXl/SvSt28+k1RflXNp42hgzWmwcN
aUq3KcnF5/cPzEBRQU1Khk7JKLry8xUTmjsXjQt/P/wm4WqaZR1A1NlyHnuv5IY8
9uUcHlSolOUIzemeWGYj74kZhS8tSK6FBQCrSKXqjJ4rtvalLNqs4cra0yH4ljoS
Sluj0Zq2OfjG3IeOBFYGUKjjBJJPHrc6+kRlI3bwa8qQOdu3VrkEQdhg9YFWBo05
7O0TVwC1BS/ZVUT0vn5vGynFYq7DpTz2zVO7LWeScGfKolvmvu0vJr1+ki8k2hVB
eRMrt1ke1UjBfBoLjpNi+6tYshEFWI+z5PxzOjUQ/0Al+J8buWksl+DlEIP4U+0I
NXk0z4070ZGUb4D5pw4AgytTkcf4AeXow6/t59d6lRqRLb07wmV8a+HGbSB5mv/S
xkXjUEnwchudDn6Ljp3JTicrOJBHUKsfh+uEoifAF/wfGri8mJb37djrrHHyZ42f
kVU2nABoTaEq9HHFhOy9HNd6QbAv5jl8YYOoMUddMAH9Paf3TiUExqZLnpAfYYRe
E6po7vhi7hB8Xvdl/GYTuRVc7zbUNOlTwu0a2aV91VtV2qTb+R4E2616ZdsjSWrA
zatki5ifKi7JXvuEHVUqVsr0Wxql5y+LuzRx2dR5ss1NFngOlU/fOBnhB60AtpO2
/MTZidDymMZPxq9ZnuF/pB/O5chFbecEXLW/iG2z0zRze1acnaap6L1kSymQSzvX
Z+5nlUyauyVdfjPB8TEZyhlBr1F101EvCstmsh11JIDXoMDgnO0xhEPzCK/Z1DoC
OJXy05k3YY0GbtzPjeAEXm6M2jeY/30Mmyd8q4tze5eaudCAK0XT1/+ObAHmAcv1
sN9/0X1kTl2j10zjmpRmR2E2Ogh2OXgHT7zYmMAUu3ZBClKTy2iv4u12pQE5NF3k
6p4KTNH4/QQUhOhCkfuW1VfpXHKbiXWK8X+HWwrSL1XvpGoRquGf9c6VWL8TeTwn
vqu8fyfJX8zuixx4E+P4cyQ07FCIhGWcUBrMJNhMzTl0+ikevsqDQWp+CPOvaPPT
wYCM8+R2PKkRT9DSsIYL4SfHM8wy9+ZDMJKJ3G0PJ+KPbuDVz3BVp5O7MBfxy7t4
pEQr53L88aeAmmnWsPnOSIK8kaKQE5F3X/u1GYOq+tmmwU1+CiUlGiYiJwVLzF+p
zCCMRNcTCnuJAlLigLH9d1Yyr/YZvXs5u8hcACEYFgGIo+mV4SLjF2jo91Hdpcoz
3imW4K1LnWYFA9YzfcdwoeuCJJ0zEjvrtSX4T4EelOZtbmA1zhLodv8B3rmT1W0h
VkQmEKrbE1+dWqqtPD6OANC8ZBhNAwuhY6X9lr4iVhK3qN5i4hDm6u3sicQ3dEri
mYkaQksAku4NjLFRVj5e73fEHWbkwZ8rVymYv9Cg71iUwAePWhTwJKDPDTUnsDko
WHrZIiFmcQVRsRu0Vv7VSwQNldPQfVSTr+0YYAiXOpLEAojEFGYUYlWzQgkOc82Q
VKuA3BwlLzRt60pETG0QM6h5tDrq5OgUxstTi4+KlQ0VBsC7+J+a0Y3HqwZTohnL
Yr/tuXKLGFtTLTyxhZDzQUpeEGeOjAI9RL0n8Q1YY3wGkfl8UD3B7OnB8XzNXSfi
ebUFtoQDFf7CsCNY0Xr1OK8z1MLRtDhoMjU68mhxJ/lH8+eAT41qs8YR/FhJI5/c
zHh3kfElx6XUs3Oo89iIkjpDv7BBO5FKWe+TKC+yxiY8HHhJHt4FvF61653DuNBi
0AH4TTq2rEVaeSVqUhjujZOmJyWrjaNj/FH3mk9pMOQUVF9w0pB7sW7RicJxtf+7
dSbV0LvDZEkxZWcA1sXPtqb98SRimuHsiFrJBOHLJp10byfn6pGuNqokv8MUL45M
6HK26DMM4x8DLBHXM8g/Ii1HywYSJeY+6ZNlAkjQL+4TyMKx68B3bPhbjKBeyyiq
j+OQ0dqOraJmFvRKBSkydSXF1jn6hfZvJj4fKCrG9vuz4FyXJ2wiwJN7SNccBkiZ
MLWdXh2j+YKW6PJnEMJ3eHZkrJ9ekn40UVWXeMiuWeINOABT5APn6slMrBO0jAVM
7PBU7jqlWZfBVwDs8Lo3/M9krh5JNjQ02T58PTc2C9lD05HYr2b6PZJBrLFjh6Ow
Xu0Nc4Hi6x6AaVqQz9NjesW6+UmikJk/5MXMBdylvMaF4tIbad5b8obBybWU2Yo6
d49dqcP8L7fEY5oW/ESNFgP+6IWWXEA9bE/MAuo9x302Pk6VHPpfuc6OvPbmfIAE
PA8PTkveAUGZFHkhVM7z/33+WdngU2759E772hsEBsfdjT2a0G+EC3VnAGi7SWY0
iItxyGsgJksCMFymK7IjSqB1/Hq1gYpOYHM9PLpFkpasxfWPTTxdl1hM2IcX3b7v
Uk63t1GdY5P4173aPIN+UJUb8Jygdhig/jVWOlRQznEq4OS7ufRSCaRIB2FtZoBY
fbrvT4RW83m3YoNQ5eRLjrjFXiR9NGW9UDEN8MNBHki6kOU/7hfBtb7citXDV5e5
ST9HTY8R0PGUHvxhPin4aqABEqcEawCv3U9YPjMCT70HBIWEdIlSHV0iig8HWhnB
XVA+IXxps5Kg2E/y5J0QUhaLyG9Cl+4+5rp519DZEuP4oZObIqCsTDA/+H3Jj4T/
UdxTV1tgLkbbH8L0UEviznursOVE+V2FoqJ++wtsNJJG7JOykvCsTg/CMnH37FA3
oFSZXIp3kF/Wvf1qfTpqM+4FXbqG9k/IEc+VSyFXhqY95sVW6034TRMo40nBlPiG
Mb1hZOICFLfAlJLNPkJDu48SRylxbfInuNdNK4ndfIUhs09ewOeN0VRsh0VnMT80
jVBBpx4R1dowRxqD/0P8Y6BDYcPLf0nMme6A5H69HoesmwmRqQ8SajfbW5tBII2b
lg7VlEkDgqVJztUkwvSa9v5J2BzO1GvniZmZnHNUaaUxN8mDxG3q3IzWu3KukqXx
E0u9JHCvBiXyy2tOk3TdigYmEqKqV1rVPdnpNp4zV2USDztH1+1Q5cUYnhWLxInH
Eq7+29q3Ep5mRxVV24yXSEINK8mcCJEsdojZB0MUx8P8pkumpsQDpJoXd/7iqOSj
e5FpgJ+tyxh+Cu/Qgml36lziPQLvj5XkYRjYuGR2hdgjSLocYpDHt/t5dyZYU7oM
IfTEI+cIvLb1XTL7L0eI+Cz+kEV7reD6SvF7yt7XAMyJ2+wIBkG0xwBuieJtKlGu
HkrL73IlUEuJGKjYmBHwBEtjSo8LDYdezNS16KlM1J2HdRGQESgPvLDlFFjG7OMi
WVEUaUOkx2m4izAAiG5kJB3EQV0IAuFNuSlyusCaG+b5nfNRRrn/ujt6nmkU04nR
QhGJ3byIVE6A0l3KcncP5NJEt3Q2/MAjQpnMrsxtgBS48PoE+1Eh39/n4Z4pHOJB
eoNnldHaLn8q1TBYSYE3MQrDiYCC5UBjwcW9v6WjOY+dnJll9i/YH1evF0PfaCX5
1jbJ+abnqmRnwqP1nPSWu5G8QAQ5zWbRMW3CoYkfFrLs0xTJLXvQ60q002hOUror
FmKyp9jjmGx/CGWYBtFyncu4shxmOcYd0n/ojJ3ez3RkeDC9LSiybHCWzJwRbvjm
9gL96vb0zkfn+zmJ3fdi+phWJSpvZDotttZVaXRQm7Ktud2CmxXqSp2IDzGiueQj
HCf/hCYsgFKTN08duQ0Ro/9pS12vmGz7KYTFAcRCN0YJrXGC/C9kI+y+uiN009nb
z662O0w++Uy5iPzM8kqSExbhv6aOojk1vfMQlz3hPvcfjNOEJb73/ZnFDAPvxwFV
7tXPU+biBfSuub9/8AK7xE+OmVf5XBCpiDfO0bP0Ti9jXhzVr1x/HGTisTT4gMiy
bl37Yr7t/2OdKWlZIkZ/+o4eORcIZVU7NuVWUIHR+Hac3pQKQjUFqwLbbJoV1xNf
8GNmeNiQXDlVM51lsvQldlr0gSZp/Mx+05nJ6JTBsIDqfbriMm00NA+yBZH+G34W
EVKQk++Dk8Z0Y69omN6njjHOBbkOLfjIn6Q1eWT5CF2+GNlU6b7YSZHJKg+sukEi
DtvuUlN2pPOD2rGWIUzrOeuV4+ExpsEL2JuxOllorptSGFcnD12F9hII2nb44KR6
gsmA0Ldr2UWCb5lnUZvp3O1i9FsDt/QNiFO4kdMhj3UbnIPUUDfYrJqr4TeVhHGh
aCOl0JuvMVen5TRc4kE4o6CffYJYIPihSkXsZ5etGmz7CYLIpInW1ZuFwHHGAO7r
Aggs196zXxEA1GGdNIlpEbdlsT0O2dSipPEutFqkZcEgLJ3Dh9f55yKxr/9fgdUP
YB4U7UF8N6mPfvee2gce3g0n5GEgrKS2a1AcH1E6vZTbgia2w4ou580+oCvJGnXF
xcRXMtcT0/jougGYN4D5CDBO6DnS8A92euTwSNTCbiY8VB/Akbf2MW2x1MqzXFFw
UA0wjmAk7W41bU74Dq2XbQlS8aD0P0qrjJFxCTqTO69+j+Pa/y1lFCfzmCA/qir6
3wTDaGJH4/jD1yB1ye++dxysKGGbukN/YBzWCuOVauB2hEyl8vpIJfJyYiiPTjxx
GlKd4Bn+BJAFT6FWe4If/XfJVSmIR1ad4/Rd1Vm0YXiC0lD6pNrM2bN1rA6Pob/m
oLje0o5Fx9O6Gy32vp4AQ/oryfYc40nARAEo0OGSdqaAJ7UkJztKubUvK0iyotKH
THWig3mgHT6WGCWZdtkzbGCfQy+m9Ex7L0mYD2i3/5ft2O3tZ47vycRhg8N32WO4
V0V2QxbXtL/VnbaIg/7d44bJa83ezJgwhF6EMmRRkJs36ISTBZiLONskNz6glL2k
iXw3g2KK4F0/jX8Vvaesep6mJqD0Ki2fdMZtE0LsuhOnuFLzWfutwO1gIZlxpVI0
YhtVzNZyyiBUxfKqIriPYlxoZLzZwTa9VwoonyJbefJfD2Ki6XdhUWMkAKpQhkOx
o55NWKfdwSDIDPxf+UyNZyCCa6rnDONvcaO3QvR2RlH1DobS4nYKA49Nx/YHXvqB
AVOcwZ9jolxgBQrJ6qSOF48tW5Cvq0DzCLwuC525W7gb6+vaYCu9++b7CGMxSVfO
U688nI2YuP8kT3i0mDhi4VheSFzky0Qy9tDmVIWpiVdtcDxF0QI6siQnvgueygcP
tP1dqeBy5DOq3QtUULCN0PaxnzuQVXz5eHskFEbX1+i8pU+DQWc3GOKy4OhDtCsj
BDltw8TyGHvr0kX/u81JJU2yrHGA4yLKSr2pno4CCssNQqAWVwI/S5oJG1Un2m4f
I4fGt+fT4oC7BgTajZWE/3LY7SHbECYlNUAF2Yc4hPrkxBxL7u/qPhJcf1Ppx1lg
JqzeYLO4JbQ1LU7VAHUf0dQH6ijkym2kC6vqBJqt97/AkH0foagyj43zrcSy1QGQ
5Fczy14lp1mqx2cpYSVusY+uiWajAx/a5ROBkmEEociYUk/lOWncUzfWWjtH7vGv
rtW/Pc+wpBprLR3xFsEPnfH6gfK+MaR+/4pCEYBvsZvMrxQ+3ZYxUV4D/0Uz485c
ndcOtICFL0odA4XJqJP9mGQHW8tIAMgCFr5ADO7eiRR18U6TD4y3x6RKbGmYvPfU
v76t9nAOOjO+Z9f28DxpSnnmU8H7wBf7642I+FX5yJgoQX0A+Xvm51iqkRKOtUhf
vx+uUnKR0YmwxNcJ6NWQ799vqGLsmPiKdGeQ9/sYUSz/ipkkSJMMdgFsH9Wp0ytn
jZscWxeAJM6+vlhuMLvMV9bilytvSTPIX3nYipMl/xJDr9mTgaVuYPuxHj7Xfvgn
VhIDBxLzk2ADbBr/1fGg/HEz/CxISuZPlOyhuRHD2RyJEil58M5zeNL4yk7jTkKa
72eiUMsL+7DtqhVLX7Ty7mG3mMw3Q9pbH2AgSdQ9/5bDtygYaxHkL2ZS65QWSNNq
/m4yNw44iv5G4aE5Mi9J1kNsYNTzNuSnTe8iNb0jyHpCNn5xqVFfVmy1q/q289aL
g9dUCcvtsqYg9oPpRUPpiUystakHhzni47a/K5A1Y5VZMgIaII8CYN3iyPyEczkm
UBKs/vXJpYxB29CAUUgb2RNTnDDw7OyNNF/0QYjmBXnPiDFRESRfV+a5pDphD669
zrhNGob9Pm4OFS0VkMse7ZhvBfiUreyZrO/LzbgXHD4klLP9xRXJUagpeOyPPcDV
LL7zszNt47xmaImqyeVzNCDAsdplp2un7BdNsLggnJCEwiHUVYzKiYK/n6Etl+h4
LUss3N010gMgiS1GGTFhmru+0mAjzzfp8nJvOuvM19C0l4woU6NO6fPl27uMOGQ/
IarX8JJvaK4SJXMaGM6vqQNtTZo5v9WYDJkPeitjHF50vikXlpIfmGJKnrj86DUP
+TpEOkUdCs3ItfCekCnaqDpS8jwWz95PeVpETOtubBUukO8YjO88BDCpXZig29GI
iqnmtHGOcPScJTxUyCS6kQ7PZ5TIuYGB1ASwD0pvv1lbcMveBTOT+Ef2oLio5HD7
IMVT8YiXPWZYHQx5Enwp+XnqQgadHVBEFsp0/htHcRkDG2cmA89LCvMwq+QVL4nk
+hFYkxOhiOU/8romO1tmuQ9k5IhIqVM0rPP5o7GAtjEC1PXOFjxEKiSNoUnAEWar
WzW2inkPlCSd3d7zMTcKalE6t6p4a7eX5Jomu8LS/Bi0Ar0tDVAd2QIV2GErR5Ki
9H2Mag3SvkUy9QBsM7awk4w/jbWCGv4KdIByHYf2IxcBehSR6J4zR0K5puGN52he
fGh3he7/LeA5MAsaPwXbhYYwT2HFBnFzDAGCCRMfb1vhof4TSPDURPtMQATAq5nu
aRSpIjA+3X3F4HPf2wgYM1WwGTN6wj0C3vcAG2j+jfnlj6zBKy/LGfzxFbjdvoKj
1OHcyQgEd2Vqjqlzp/3MJnquAuZHpOcPjeHOoAniIthk/SxnprcMy/2YYIrApBqB
ILx2vPO9srMoWtjm5uN2YIUAikvv2fa8KxPMtBcGJCB9Xynt8xaV6l7+ILxvnQpo
7ZBTjC19izHAjq0V7hm7mophMF4fdQj5C/FYbzmuXNAqsCQ7daBTF47WYaAxmL3D
/Tc8C4zmNSwC4CpdGIrfAuWd6wMGzNlP0gkqAjaILUVg5LSYYfe4TudYUnjzZZRb
JirMtCEaNUI51STAP8rQjcPLzr/xvVt61AqvrFncbxlvvxQUWLAhgo4Ijz/ns/WP
YEQalm40tj6YcJto/Zet6ROlxdQRbkkjqoWosGKWTKMJFk2tX7NbpUrybwdIMr0T
6Ovg6ZB+YkhBG1u9ozjW1JcdmtBZUISZ4amb5CbxY+gYCElOZG1thZNRftw+D5OO
YipWZk3E0Csom8HGKX8tOqw3L6MkNz5H+lIL9NoV3Ojl84Kr64+A0MyvtsSTy8o5
HfDx7XbRfxCBSj7Qrsk4G5Da3xwrkjKwIadqZ1RqjrbGPmsIzlDB4KuIkHhtjHCf
Y/jq4zkKcQseuEPaO8p2/WUpmKUIm7GgkbQI6YLlnG0OwLb8FI/QMQbjIWEkMyRP
d1ESY4lXG6BPcjo+QswbZRDXc7EBDcHQaIg1RB7id7AHX+UeeZ5XvmMmTeo9aWQk
6O7q7xt2ROPaaDP7OjVIQ/sIX0S2w3QaftAWkKz6yQkzh3C2114pCnxvTcmJgnUf
lUqt+m9/Ooi4q1iA7MdUqgIMfv6X5gr+4oQLY5/bd9kQeFFUiVPoHv51USOIS1Tk
Qo/19VMMXI855tj8QRvrnNEpFQTnYNuS5o8HxyPK3s2JQlRZgjcQk5Ud6fBtADeF
X9u4YDSgnEKW1OnHmxk/Xq/6x0sSz3CH5kmK+ph/8RaNxMsJaMh4e25VHpTUTQpS
lA2WsdOwWkTVMAnwkEQusCSGN6bzprttezfQn+sZVK0fni81oreY67iEizRIhtKJ
7heOB1IwUKPDwmUIL6msUtiCrhBYltnFy8+1qQVMfXtjVmFLEzk2ClddPOtb/jH7
3cfc/rrDi++eQEuXr+9MYrqG5+r/6V0ERLLWrFxVGdRXl/mydPX2WHGPb7Z2MXeV
dlmThuLRUicAbqeHguAHXRPlvt29Y2FUPE6En7Jdk4GnbAPOFzXslmZhXjBgXPpK
C3XwntSKVDpn/+CgO/ShPRfDDDZinCxlIXH6co0dXfb2KDaWTi8wLCB/49or9AP+
qypy/TnNNt3Be89Vv1M6yIS10CKzS3LATsZSNigdlvRszzB/bvULzG9gAsa778MY
t+MKeSuOIuFRVxBRE/nl8JV1QLRcaduHUk63RBGIkRZTyCIY6VR8AV7Nf7uftsv5
tlTg39xrz7l0N6tOxg+j1M/sOdcf+XOA11XLvXDyCRaRDgYKywReefNSJv1Xe8hL
1q6vEl+9/tWKZrO1hz3geQiRJqthF9vuc1By8uqNHntfD5lqMKf7jUUHUoChC3Rg
h+QWvtgsrwCWpMy3Z24wmOxP+RWr4SmcCbY9WZYZA4fLPHiRCvPM0yydF8lLlA3E
waimZCPGuc7Otm+BqG0pUCE2vScMGlIuEw67qUEg6AJpQWuDPDLbHszdv3Nzhos2
kUIW+2v8Dpd4AmIzg6sypGRD12PbvH3UVXq3oCS/84bIBUecL0X8lQcwoKFAlKLC
1qt4OTm6VbZWpebdc7Ckp5NTr8fGF2cqldbiqyy5MSmZC38iVcV7f8eUGi9ciW7w
WtOAlJsDctuJ/SAo9pyQD7gsiKF4eKliX1g4saFmyYvGR2zif6QlP0bHlPdF9Y+w
/XbPhsP0qH/t0QI3ONXkVIBVbnN4XdVeMuNb5y7uvtjbR0vWcV7eqXMvDpeyxoSX
UQWw3zCNYAqhdoDQn0dwXrpYntSWkS7LLY4eDv/IXyBiCOnrnheD0JbxKNyrVRoA
LdkY2AetomzSkMD401nqtM5GNXDdE7yovGz5kw1+BFfZOwst/R1k4UG3PCShHnrb
G3hDWtz1nyt2ZC1Ldo41Kh1UNJaTjBGKarSepKT1MhqtgFD8wd9srGeE2GuIzNzO
sQbLBzu17yqo9U0hr0lx7KjLY+cy4Iq4El973noGkxQOEve/aTGAUgK1ANAlM3At
QNEu5FyEIaMKl2OjzoqflznJbw+qzCRXP1XB1Hq0WdLnL3vLv7wtniptHaBodZfi
/ny5kTMYWxVJYudIDuJvl/Ca6hUZNqMYGr8kITdubP9U3ZC3xUFh9VLiefbF4yue
pgF6GMOC8ll6A+5K5av+sEb/CffcccFcinbp08hb/EKVFXD0W7aGCsx8BJCkIXsg
ikT+X0lyqmsueL00+sZTh2q5R57QODFDIJsoK9J6WSx7waDpQ5sE5XsTjJxZ5LiV
vfwv9HKUKRx9acgfXmDN05jn2Y9RXqHe9QdwpeGnx/oWAKCQHZWj6XB4p+vbxzjy
cr+d7LZrgghuTm5QbeoLfZLoAbsh2dGC2MZyFdSGXPnz0T3OiS9A6REVjpDfElE/
WdG9K81OnEcHmRpow/djApY7zYShu4k1kN7lxGDlnHokor5zNfCkbPLjOL1tM4qW
X40jEWRJwziFmPDNyZ6IYRJVCS95C/1ZyxBEZdSkUIAPp7MUtlSXN/ukWJlaxzwe
UJbfPIA8OYKJ+jversLWVHrKvEnEfIpl3mcAAPSfBOsbJwz967mxuAvOPznug19r
phm7TvLHVq/5uylSqbuEqlkl4Tk+5yuIljddkVzcutrlmnFqtS1r+ubV/tepECx5
NkEyLnYJBGXwwTmnLFIvUtVtYKLtABK3tNk2uQ+c30n4aO+7AQleLnctBAMPhoif
SR6G/ehk0lrayVdFGExPVnz627vHidK/9u7Fb7DA+CGBJIaoflVk7tMW5e2rN0AF
l/q1xfAbnWakLj9i4i8FXAT1ob8p+Va7EOUKvkarMLuhxk0MsLPQMYUw8GhGqyO6
QwHYSetNfYGO3Gbo3RrRRSdqlLf+TatGpyirMzL385GUV9SaIwv7JZ354j27p2Oe
GzWKQDbD9wYhUCMRfN43VDDKo0s43E73gOSJw/IOE+szGp9HUQKj7fqY7VeNSAkI
ivhXsWn0mGUg5IB4bUWzA/+Clkj9ga6T3TRigfhX4qSwB95CBP3Xs3STDR9zkbhD
YBLQCpoteBQLJJE024z3n7DVsnOnOvoIrtuykMQiC7IIbkhBeVEZGaMzQ9N34OUc
4r8MPbIU6FXYrmU/cJM2Imhe6ysI/trYe1OM6pCAjQD4xpH/YIGFb0W07tq/IDQ4
zCq0tZxErpG109RykA86xlACKCvMLxmc7nXylGtvE/6mDAqNLfjJFHp9U2Rc2f7Q
eMwSdAL4zVPu7vELkYg5OEEPy/PVB84F/WP1SPX8PtvhAkq0I23xHCzGGoUWbo6z
j937Lo7RCL8Z13q9of9vtf4AKcnNw8qP6escXe8xayfnnfYqZyYJ4YtY805XF4aS
nWfUhM5FdmQvJlcEhayHOSrsyfzt4nRgmmDdtmJ6l+VGFz0c7eZBH+YjLg6Pf01H
cnc7Y2Gm1dr75CdkNHVJqxpbp9oWK494YV5SM44j6lfkU2mKK6IRsECySG1nzZ5N
UYh7w+D2OuGV2fRvPsyVjCMhj2kNvI1aKST4bjJ2FQ4N6yj1CTvVtvF6TOV7souC
V6YOiZ3bmx+w1N4qLZvCjX0gANsxt48B33Y0PT2l3XDCcaKnIuDRcbTQfCavrLiK
ia15MdeGOalvzo1myN+peMHHwTUlRj0MMFJsbblfRcDUPQs0Uvpf01hDfTopLIyV
jj99sAiM7N0l+i8J08uMIvL+WmV5xy8lH5j2oTTmc1ncyTnKnTxzX+lYGr3H3TSP
JmKbVZXFhlt3RuscaQ6vD3AZ/pzTk4jey6TVmwEN6NTbOHmagrummHwL0xWnnhvL
57m6TdkqqAhMoS4cWAFYOx2aQ8Y29Fwlvg9bpaU5RhW31Pxia0Sy9ormkDh7dCRE
O6Wffna/hk4t39SgjLx8wbPnkETHKL60kOCdMCKsO/t2iUgixO3KeJIOYwnDGn8V
h4Jt7MTout5f/sZE/XD3+6hRSSfhItOnlaia6mcJrpwYUT0AFbt8DW11VacZiZYQ
giUAfNCJUn7Bsf0lpyyubRvI18G9WwJGlkYQl0AmB7Yp+4FIwUZNl/cSpnwbRJQs
y4ysmXfeD7jo/5/yj8jL2TafmYyidtfwRtBb+lwLmnHfpzHOIYtRW2d32js2eaiC
iKVhyHTM7zOSDhvqjJpUuFLBjUP4UsZtV4wFfzAarGik9g2F6vzC6UJEUY4vTVkA
/SXYRLVdNNIx6dbIr0CVtWzR7wca/n0AXU+iXECmshR6w2eI228sZVPfpOfx+rns
8zZwHrYATAvrbkd2qGwI3vu6C2GylKE56YKBtzD8og/wJeHG2RGZ5t5IgpGri4JB
3bqGCT/p8J1ATUxE+WvFib1mJQ49DQ9ilbp2u7Lf77UzwHdNYHGKJEy5yjpHHE6S
civ85OGPqhu8juYzNlCVi5auHLGbm2CuCveLKh0I7vm6GSWcdFfLZrJiNzDV7svz
JGVnk8qj+TUyT7Ds94SdnKp6z2AryR0WJlRgM9VmM5GCFqTZQqU9N+PhSDpdr4cJ
dw97Rj7679RAepWgaoCHp6GokI6Q2h4h4mRmpLvDn1jVVtN/CpQar4iHkxxl4VTZ
JjtvFwCdWoy61P+RaLF9M+FVFXr/9vdwecT3D6cclpvvJ1RTrp5/Ask3ZjBbTnv2
O4Y+PZr+cc0ls7HoMDNtSeSoVZnuyQ6llnpVKT+UrNyzqKmVUjT1zats1sU60csy
GLjTxHekqMXhQIuUBYyjNYuF1OmCbb7mEPO7VSC7CyrP9Xw7lqLl+kVm7kqIW0w2
kUZSRPo1+dMBcwx4b/Ud+VO3FlsXytXN2tXyPR2MPBGVb0RvRSu4wXIQe/w19Nan
GQRDb5pQlfQM0+py0ppZsrsUc785CQWfmZno6+n44/Iph3ngew/nqCpiF1DXimGE
VNEpNl1BIq1Jgge7yuDqw9Ow1J9sOwqDD/KBBna48IgsT5Gr4u4gdrBvse+kz091
k0kbzaHRRF10xzSUYwwOjm3imJRr6cbhte/lJsa+xNTHpFT5ICItEASD1/9Cpv15
cCTbXFAia0VLQrKNOQgDz0eGlB4qEtIR7TFwMnpOPfrYm7PJQuAOTWRlPlJDY/6y
bWqNtvdEV4ld6D6UDkMOJZkFCxiJZ/Mxq5OPhhVgMiFa/3ll0/DjE2ukqhJwofR1
Sq4XsFgvXDGGHtOSD0XFm/yfb+0VRaBy1gvOL5oPxlt0I6p6rJNCGv518hIfhlF+
PsLbtiPsLZeDmhvEEvASKOsJlQ/Sdc0HDFoWZgIw16MT9f68AceTIgrkp7QK/aKH
RA3kgPTy9PKodeTmwg1RK+IBt0c+hNWnTuWYubfgsfPOfBvaVX0ABUiFdqNJpQFT
VFsPpNpS/HcnnzzJH2q2mQe7vlCddiqDnfoUaLtlgQynEFPLBnnki5MNWqk+EiEd
VHEqmv/dsUW6vnNcmjiVZGdMXXoz5OHPlT/88/vXCA3cYR8VbzwC3z06mhI98FlJ
ubJ44DEsH4wwHjUI/nrmD96tQPxsgVLQiycAONdmE5sQ8TIgUzD3Mx8S+u3Ewe/Y
Rq4H8IlS3Q1L5vRGcl1340thkx9dn9KujWYUjzgnyOK9n8CRMhv4E18VHHhxbucX
2WYB0pzyKRJHxN9rydYNV6L1ed5X8th8A0iVUJ5VUPnjQ7YYruSYnqr95iQh57Yz
UdCIiemzGcluM8QuTSvrM3lDv0PrALFZb4C2IdrUV1yVBKbbvV2GQfXqHV9XtWT3
E4fvbJYL7ALD+/mS5JtSDHS/cqY55V8GjSzv/86XTMHtmEk/ZCmicLedG5F1PsAI
rmy7M+WOnbbv8CXnfttMNdu98Ip48ybOL62KlKFFAV7D4DdyRsWS65tbBvF5F6/d
Qca9z/qickmD0fpEF2SfZ+g8mgEeD/QgiNWtdlINQRQFZ1UpD6R6vLQTMjb1l4BH
/ssdaCymMTx4hs61ud/uDP3x9NNeFCfsBlV+14qZB/F5ut39ZtJ8entHcj/+pHA9
YXdEj43z7aoPUQCr7HxQAhCNm31RdhbI/r7sMufmJldnlvf04tkDiuPGEqa3rm+J
17oVV4td70PmyNCblnMoXKWxLL1xm3/MXpbHUWCFYG64i7NQLcPbmDrRysXCd870
o3xvzILGwIueEltkd5W974jraP/41fQ3CRnONHYy0AnTrwo3ZdZdC/2rw4wVptPh
ocm9Ur0W26IsoCWTIqV4IraodLlyKyYm+W/deGVRPScrAeDEzew8JebXubfYNrcO
cBeMZV7Iyb0Npkt0UFnJsUy5aTWxaAtsEO2JLr6M3Vc2+tkQl8EceMhiKjLZZPKn
YwdC4p1Cc2/UpQSLzDJMQQTXS2IkpXu1PklCnA1VtBX1xVVOcMnejIbZvwFjlQTx
CD/vjPRN4zvkx4hqzvJ3QILc0PtGPZWN5cfgNo3rJe63wqibt/2DwXKlgSSVS7s4
PGBkQumr/nHgQtZ4sPYqfLA40Dn+euG/JsFFoI23W4s/tPVAeiBe+HOafW5VcJn/
AaDhsoo8cxRRVtBpyMJD7m5K2p8irpO/eomyAgSZdKYzQFr20+ZriFoQH2GyNcsU
uKVMCxHLLcSLbWd6NieWUng2aBCmFXccjL7/5SlGCZvS2ZIVfSkJ/2lGJVMqcIkh
Fuyts+E8meUgfrKxbdqZuVf89+ROXVHiCX56sIQvBMG7SymieuwP1ny2e44WXyDl
58GVC5KWP82hn/3Q+yvVIR9pAuWZKTiX16DsdUX4sJc46FNCBulDM8LcfGgqAf7F
vbhnAAOIiOzuQiB6mXcJ64GT1YX1NY7ZF79hbrxRuDamb0avHzYmhMulXPeYLHoc
/GqZm6c611nIs4L1/PgC0JikxwENIRi+WyjoAP0vgu4PKSTtuXG/8yZdc52LCBYU
DUx0V8RK0sOXfBDye/orXuDoJSQYSbge91mDOItE1pqXuzSfajEaAk0qNJxFUL15
LxOqu7f5uveafmiZVeWgNIB1lU6cb+u4pcrtfX9fokzHG4fanpCprjjnBPbeUKbX
2qYKnJ/G7DS/BEvDjezwnRygvpQkONW/3cQx699Zb2A353an9Mxn6atP94Jkkd6G
BT6wWG4iaN0z2y6RJG3uXk2QoosQ6w4UqhRHxYRRR4tuWss/Nng4Ho17Dz6kqNPj
oNwB3gTPo9aE+VQDE/wSQrtTXNFHssP6/bfvr/nE3hU1WDVCKmtJeiHMUYFAPRAZ
fDOzEQ7wieyl4yWgB++zvRsDG7x5ocI0aaPBg7ZyCEo/7ExRfyzxSHt2+6h6nuaq
sOkhseimvA6dyiZ3DwSRJAfyCyf+jehwn8U7tgoQtOmyapzTKqh5eBMvfPqyy4Ws
9M89wWFuuM6spIHwutwuWmAj9K2oDzLkQO8zOhbZmVeoL+AIzM0m9oaYAXr0pyH+
udw1yt/jxjwUr69tvreB1LFUWr9TN+RhbhvtgT6Rb9kVHew2F4B65HRgamGjvK3q
C/swK88IoLBteKmiF7EiHTJUtgY8Y7qvHYfwA2aEtEMJMqlHC8WRYUuoM+B8bHf+
1Hb5P1UTUGPcqFiijMW+wA7HNHs+hsNxfU2XJStB9aqn1wqYldQKrtjltNIWB2UC
QTmEVirdu0u3hK/Wjr8WHFiQCEdo+sw/A8nx7QyUIHVsXDwOJ1ojOq+vU4HCwvHg
nHEar52XGYwgqrizZwucKNe+m3hvTr7pCXAayB8TtJ/zefW1j0vsxz63wzI7wUcK
rZxSzS99TbzjnImSc+4s2GFEiLUQEAidARb9X7L5Ld3GoLfSoft2LgXxV1F5OcJr
WapSO17c7A3vj2uA0fgUQ3PuF//4AgSRuzOrWIkxeJWgRHnmz96vcaMZ7BjGUsC0
/y9a4fRMLEW0ygMlbducLvtr9hSX14A9Q9PHQe0YUQjSqS9/etXCFTe/5wu0K1Ks
ub6fWOkSf+V7bbgWehS3vk/lrmZHrPwjwfzoZYeL1VyFpqSKwspuvUYq/rrHrhrI
PEeluJ3ccj7czQRRW+hPPCPobz9VQxabhTsL3l+R/HNJdML4xKcptihm7R9IiJxo
7xTAhj2ZzBLG9R/tYetg96/HLVN44HoPp/m8ajp3YCrNtSU6wYfNHbK59lKGesud
ZFeze0QyYsp15OhVybvpzNCP4Akh5+/kHbeUYQWwBZVl5sugF/Cm10t0FNWJhut/
QFlCLSKqXOGwldF4u49hWcOAHaiwO3/8uZqQUkAGkTN8C847WbAwXHyXIAANFuHH
NAcCYUCMR3Q6V8Sb/pIutLZAKOaRzqJHwnBoSpe7HAhVfDfmN1EvmTwHTotW9FCf
8Rhq8ZKxa66S2Sdlhc18CU1u3Pe25dAs18c0DF4gsLEoLvYdXlgX9Gi0Ug7Jhm1H
SaIvUeLX5qLmQRo5zHxDeFmK/QEKD7tPmiir+gKCFDNxhHW61xJqhOp3vOlpydTC
WBwATEwpJ+p4qos+zyQlYH6Q572+oAzXPglCcalQeNnyEifMgOV4wgTWigqmq8od
fbJf5DaJ/n38osf3cOi/IYSD/bXJIR7EFgIml93Kp9YPaVN0QeDqNbKIx/5lcMof
6z8GmZPeTlPiD4db5h1PpDvx+Rkdy8YHIY7ZYEt6/CQX3WPU+BCWU4KA1gtdvgmf
GxL+Y3ZqaolhOeE3SWnGtlMfyjuYC6nx0uJPs+kET7LVKyAxbuPMyleU4mdqSc/y
07/N4jd8hfrYRUU21fMvt9BwxMySUbrTQ5jBZ98jBfqvZoyaGXzgo5N+bLbo/bqX
c2xr3r5AnWDn4KS7Uxs9Fv9HhcObNay7HQxeflNTtzTVhlfofiwJyg/pkGwMUCe3
rqwsxhmTEXWszkDqPnEy0KwmYj1j4t8kFrAw+vhMwGP7ujD67pPImfUqpCUpzDvi
FQd2aoFPCT6dho8qflhY9hHQjw1Gw8YYQl4PBDRb78ZB1cBwip9GEqbbzE/4rML0
DxVY3BewJ68Gmjb+ct22FRvWmlkd5s0Bij/BKTVmlkRUc6fAw6oY+adIIRLLvfBu
CLaHgK54ku3/b0H01R4Dceoq4AA1GiLDPKxuVGcbkkV7ruFOBdE1pZ6MFQrixKC7
csPDw6oTIpNhYK6HDA/KdHUvthB1PGgtVkf1i1PZTiKhqdfoXo2Ls5bJI4SznUGC
WzYq1mnDgE/p38uL30/80fyGtWl2PYIkZjTCwO0L4DxsQVaXzm4ggav6GcxdgGu4
2VSPaWn4rN/+y7caQVvVvJXis1+XblY3RqjSPluQ3uUSOafX2j3c1IY5NIFLfxiv
3rAfpGA21tDByXbYkvrCG3h0UVOvX34d6gMHpV4BpA8jJNr1rKF+V3FNaRwIdTZu
oltYEejicQiuB5eIS88t+7mtXi6DZHB8DElxQPBYv5Lnl1meoId9uJGjC3tfdELe
nQ32kxThSNeaeeUEaeug9bM/ZlsY7nY/5Kn2DZk+OV3O2QYPtc1bt4hGh1A0Ogkn
+lHV8Ol/AxxYGixf76a+kzpPXF8wWABAbd4kXzXJffRkfNnIYI9QHqqwrtuDKz8a
/XASJlDQuuKCCa18b3+c9KegGfuj6qe0gyhZeBcRC/6YwI970DC6aDmvgyYgv4dN
ujHM117B2RfyvSadIbNuLDwkrBA4gzIbUNSoTVO+fEkN3QzpdvQJjC6HW8ysgmqx
svwS4T631uE9hmubSghDNK14oN7rU/Xi6W7Br3cidfB4AAW3AlfYl6a4yl+/kqM3
FQFNutZ1VUEldfKp+hfH/p6b+TpfXDb0wQOlJDB1EbukOwxfgKFEAG7yUzl0SYoD
v8R05FsRe5j8vZU2TaxLSPP+J61UglLUc2kro2EQKpCgdXyMmnfZmdP8XYoxQ3g5
jlexWa99zHOFuDtr/sYaHDZc+r2p4Xjf7qVNBAvKQuVKGMZX3emjqSxyVwGT4CjP
VsqUCc2ZHk39FYpuUxaWl+ioqebfGlgGIAZU1h+lplxUQVV1oqLIUMNCr54r5ZpR
nMJUB0KRz+xcqZBw8TmLAxhiAJM1j9eAphoOOPy/38c0SyLPNSwaepN89DfZO8qt
2RIX8i1N3fL5NNIZTxbKWoxxMS1U+k+USQQMmScV6k5mdAnIlvzi5ZZ9xryZrdqX
roCaOlf3jARLxvSkdnfm2gGCmio/W0yAb+/BTyf/uWcbKwZoJQcbHB2gn/7qjqoS
qptU9bW27wLWC7uOdVWtSIQbU3mioSHCfHCYUAzz/utASuqRcgj4cppCHrZSXqHO
4M2J1qy0AWvrObIi0MmY/g+zkGKuNfEhxV4a0r1yzj522lc//PZuDPk5O4aqQL6d
wJebiHf8X1hOg3oCGGfHhFXy64TJ93lLmmjD03CeAhygJOI3yeqBfQJwDUaptSlA
dx2SemywQtT481ic78GUklUtXKOjLky2xBtum0sNEYa04E92d7aJxhk8VZQXkcMN
ZIxLRjsal1jYM+zWQSb5vbmUy0ZWrqxx6P5pT8oXbYZjgONRN1a0ZMgAuq7d+vUw
0VyEFeBvBXkBYfHNLZyHmoyp7URxjX3carO+fwmNiKCKnVR7gvAUh5OwzWmDRp/c
bJVTI8HBgKd24yO4MEZAd+4AG5Kze6MCAAMMMOJ2lhWiKIFYn1B1a/kTQaYQ4X6c
FhKkUsIfjgHMvaVeulo5x+SCEDX5GLmOHX5aXM8TpGCMbU2C3bp5TKjN/lQBvQc4
zaW0ELrHc8+TvktDKwCBKll2sz/qKrBakjx8KwchoWH1XuHMMwkBz/DwmySNR6SM
rhSOCglfDWgLDXJ1e8sANIoakxyW8DLHBwf6t4KhD2fu1Y5cOMCkQxguGfD3fowR
thyXdDOlHU5ic3FMsA0KbT1Pd7iaL+XMV1BpiYz6YY1hbJN9VWFHiKz5tIac1QCV
LD0cLpCISJ788r9fMYeC+zd9Zky33OSYF9qnF8970meHEEkZBkiLMSDwM89F3ttR
SByL03ff1WwDFCGIRfAp9wWGW2UoeTWgrrDr2gW7fxioTvQv+EZ4REpZrxzSm5EW
xNicEoIZudiry5nZ32l0WyxIJWufZ/I/qhIytegshf9IfLwQGv40iTp4AcB+Jrg0
euKviulXvatb3Zf8w7GGOCf3GY9CRMfOeQopJIsqrDL3OHAO/R3gX3TrocCSAodE
HRLo5fdmk1qKQsNLtTF5qYXdT9LjoFn4mG5xy1tof/2fDpCM+mg4bh24TV4M9i77
vcR5WN8k/9mDSHl688nJXqd/QQQWv+CdazYBpYbq7KZRwTVla84ia6Q4QsVVRU4E
OgngOaXB1po0adDNkR5g/y0dhStJWOoOYgWFaKm0PqiT9ZWoZQLq/86arQErNz6T
fe5qUDujQae7n9ieXwMcnSLrxAGsJb3snVnC3USwRUsJfvBXHvbSmXfGA/2OCTam
FPwKGfZWk70/zet+HO536YgT37g7Yb1WRhrOBLG976aMxY3gTifHfKgkCKlq2HY0
t0Ggi4DLHCMVX8s6H4fKlY7TKGQmXv4LkaU06NSFSTSfL0M1CqkqZdaAw1TgeXyF
gUidPKv4+/afoHAMso473+Rjmwj9X6wGfPfX6VULFnd8oSH5Py88pzlcwEiSzAlg
Src8uHESykjkcZcyNgKNqg==
`pragma protect end_protected
