// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W22DEXLIDdOiU07ABuqzx/kj8uu5da6AWmWE0aA9CPbEOf82n/UFBGsUsDmX
n7uEXEZwdAxcFeD06ieoeKoi1q809HS7WRJvM4Us9SnqQnUcCdF8DJTeSFhc
b5fFZbZfIIct1GPdW0zAWc2ACCJRK+p8GgVP/JfUuDrmNkzlOV6beJBUdpIO
6d6IScZzjd11C8SlLW+AhvrHLXeyC/d6KJvmYlZ22+5sXo6YGLv957OxQ1Bu
2kLdACPCzXQE7Qa/2C2hi0dkioJpoSgr8gNd6CqiKCR3X25oumt6fLrxiN33
Ukx/uLVgLjOPYO37lAf0/ff2dJYyp31dEGJpbR4Sdg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GAWCz7Rf/OgVGFSqPj8unZHy49Kc/vy8e7TN1WIIZrJui7gvUtRwZ+iQT97d
okl5I7kGe40w1NG1cdKkA/gIsNt7OmjhjoNw8hiKunn2oezrTBjy5o25VtZE
vCRk/+QZnHGEPTe3eXA3hg6S9JnZiYy9Zsn0P69VNQvvxqezZJcLeScRPMUr
828YX2Ks4EYdkodKBZeP+cseP/mhy45Kxts728cyTypHRsKXWUtli4AcqQXz
+koebkHNmMReo1I5hC37IyyE54L7xxIDfkSfjTvPn1UKprNjR8OITVi7uzOF
4OJbMZwOVmcFsmphMMzwukbYeNOMkboa7ThVUEM0uw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XfxegmN+lQfquXkUgQYfG7hFKP40tK4ygYHUehmgixQDccyv9LqDXoOpnfro
9SVXGz5fCJrYz3Xi+6Xyv4SxhRkaXFUjyB5hGtpwgHZR3QRseNEyL3l8rzTI
PgtElO9/4iVLVkHGD1qz2Z3Aamvarldf4UzOOZTqXJaUKvHcIvQxHyp4JAfK
mDNEMAttcrBeR3R36zgrW0pz6T0XniUxmLybtGJHIi6BwttrimeOqAbVtahM
XVGvEBtEmL54+/NgqaRg4B/EU7ra+33kfeUSXN1cXJ/3k/8D7mHuYdH4X6BE
eFe3eTddmZGOWXQbunqM+ZZGhjjRc2PXkWF1wFF9Pw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cyXpgWDDNiY/b9qhpE/r7lpbzaWGho/lMXZ/mBuqJiNA8D/EcIRZahUBBt/T
EN0Z8szXqhXVqWUNs/8v2nrlaWucPaTQcqZE0Md0ySa9OpIvch2i0813p23b
04j1rUQ/mdWYTxlZVP7CaG36gpS0Ot918IeJ/kzM6tFSGUyR9hI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
H1zTBw4CMe0hZcwBlLLlgTsyzh3fGBWKvZ0WgtKuOarqhMjqFtQH8ACodhE1
KlquH8qcyJ7VBk9mWQpbcqEU1o01cPqFW8Vytk6AB5p7RVxg+rUXs7L0hLxr
wgmOydIgH82Z+0DHMAkX1z7fyyJtd1xMp8pdU0pRDsQAbX755gv95dJC7juR
xErPAoXFw6zjiw1k3iFZvShgbU0isPpYQVs6Pzed6R2+3rLPCX+lh4X49fde
jQvWVwZ5sARK4r9ziDCIKkm2oqd7HkYEZWmwtXgupelIaNJMwV0jIiBH9bIt
DayienG0UP/rK5YKhAdFBZi8pSoQUo2ix6A9vUJj/i62lkSW6FMdb5tbA4mm
lxY677Ub0bvfzJufHo9B0ZuqddDLsqbYb5f4kna9qpSMV3qPJeBWoiFDW2ZX
0a2pnGWNDYBI+JT5p/lyJeePim4BTwmDKYrkZVLUqprhh2Sn56QsWzxKH1iF
lG49qSCB3y2ssLVkTVGn3AABEQwfxF4y


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
saOHJTlMitmM2W5qI8miDs1eK6WoAgaI8sb1jQ3pD7Gedw/ZsL9NDzPScvZK
robs4rB0b5OiaE2x+xrNiYooAXTrhsra/GimZYopQOWfwyLnNJX0pKpTUnnB
mzp1A9SGYmmmO0Gvn9um8gebELB0TtVL9CKbnZr33IpV+W4ccF8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oCk0FJsE2oOJ5lFgSdQa9i7ZYM2uigg1cFebmiyvxZnNZ6N7ptJ0qrsnQxnW
tI/7hwwct5qX1cpkYkA3byuqyELWoKT1eSSag42xEUQlT884zJPWA0BhGGmJ
7FNQ3ZUjk/BLs0qs17ATMCHxOdK4yNEeZcZLrIWfuWYPUm+7sPo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1248)
`pragma protect data_block
/eDWaIC/4lNkTgXbRct6TTKeo5TlQHlTP4S5FqE9I4cb7bdDAP13isLoG0SG
EwLllRuMZNXaeBIcNQcEJgxPqd5Vtmek6HBWhzYTm6q4KzBWcSPFIvJvHkMt
dOf/dErZpPK7XzBACyJ7Cmeh4JNsDaY9ReM1FIGsufEp2HQ+rerefDlCjWuL
/HFUpGgBpKHeu7/jLubx0/hSiyXRHz5z0y2ziWXIk1TEwHKq5eHOJ0r+bm4Z
m8JWq+b4lvO/hagJ3uMyrcK8HSXqF3XyXL5gYnI/obeN2ehcnUPQgq7bnaSa
T7Tba5kKVw+pE49rg7QyrwhBpHEUTh09srPZ4M0jCwLNa/Pplay9fCgz0o78
MSQGeYtULPHxa8X229bv4NbsmQEFb0/ScM6MD0BKU5QKN3w7nf3p6v19xBzb
hLQxf5TDavmJ9ipZg6QmhfE7LBAek71Mtm+InPm1w3lLBT5E83Un0rLuCt6P
TQulx+dP5qLVYrBqd8bc8e70KSjTAhU9nAUBnggVYvuZT7U9u0t5u/Sq7Lu3
jgmuWsCIpreCKnW2xzEmTzV6V4opg8ZXueZLogRx0NS2hsyDOzEslY7SvMFB
hAsGDhLmnJ2Gu2UjnCm4x1PU1sSSd/RMr3DW/qwNI+Pa9Siz1J3bRa0/nNoO
yZYLzX8x+vNfd2Ced41y1sDzwxBrZQJt/Nn3zna5v057dn8bK8OlHzgck/NJ
t9VQLD6rD7shz7EjZxzLiALvvWWMD6ziWZUfX7q2xORGy5qCVnDGwZNo4ffY
bnb5RhghFCT4QT4imI5a597fio68h+shYvbDbTwsgOyRB1PhQ8wOBJJFfwx6
7ElmEPTENZzAdmxj9k1DxgJS5zfr5t+S8DjN/uOvY3vtp40EA396vLCVzpwt
4cqkfvDRpUVwzq4ZEhDXGveAHJxJ5ggh8oPdLWELFs/DBGhnLOCOypxDsuK5
2DZVTdyothlSE/xs6kWJLhKEpvXl78i2Ucm4GIb0KNvPnyhdq+5qCHEhNUmf
AmGkMD08gscj4pRlFpBBnHnxHh3zIs2dsd0Gf9q9F2j8bgw2JeJTneCd78X3
dS3u3mKdFeeHDGJDbVxwlhuj6MELo54H4P12TyCyMVgxzUD6F9561pyojI8q
MJsIQWkJ23UhI2Pao9GKwOLvf67IthDBO2g/4E4yJTt/lc+4pv6j5VV90+lO
DvP+vJh5XCej24Y3QD8KvLTtpaASroAwv8nimcyhiOSiY0IrQy5f+eCeleHN
EnFyt17iAZYSJX6zh7vb29U5i8FCBndU3nosZMSDD4yEG26IMklFEgO0zP9y
9Xw4eiAvnOx3JBMaoOGtVdxsWCNQ3EyByaxmEW32uPiar2H1L9aSPibMFdMu
8hseqmyAbacOEpLZUhdiab9tsA+rMan7R0V081geRhZw6zmY1CWd9JJk6F4r
EikP4oJwtOxfHeyvPGYIZZyMnzHpO+MxiGbWxE4SWPx/18sCa6WxoqDdhnX0
95XUWU/MR4z5CIBSUgQDqMuPAVflHG9ipkaMty7ZrH44/oXNluaPTK7fNe4a
nga9PsRTDV9/Nh/g9X2QeXFYP7ihXHTJxJwPak8gp1V7fd1/1hGbnQ3pP9LS
3DNuMNBVyc1/bst92pDZB5k37PxXV3fOcB5M3tzItkSU

`pragma protect end_protected
