`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
SzEgHuGeOkXsB+MWb4WnNQwyKsp+im9S5c4iN3pU+MrloQ02x7LglW0SNdi84PbB
4DqpgkurUuGIzvnTwnM/EoSH7xs0zE0itEWAi05KTwVrKpkdeqE/m5LFU8tXbPH8
wZU6aXQZREQaGrMCVObZUh0wVVUkEwsuIxGCZPcRUbI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3552), data_block
xEd5umAYVwAdiHdn5UyQhC8mcW1FjSZjh/K62W2NpH2LO2Il1HZHBBV+YAEgckPn
9NtUR27FrKMspIH3eBX5VQ83bg2QgMIrCD76gObr5z7ZywIMw5K0OLMQwoKD+Lc4
ph3B2qRYabMlta3A/aTXQTXLmkXqmoWQsBfi6tg2CuBOTrUXZrZrVPGnAhIKhvWy
DwzcIaMFvjRH819bmsnVYx3p8qZMRczP+JV1le35pwLNZXUnAXm1FK9pLVg9NcE/
R/B6DORsoQahbQXC5yFl56zpkvK40+VEbFguwVih6ZLPqAZmFRQlqOJsRTRr/oh1
ENfssgqkmxyvjWMdRsFd5TCYLE7YMj7SRbSyAX45BTCJ88+WAEf0BzWjjeA2MO4G
VHZirnXtLwRWHBAaXjJML4TnCmAroDOnLxE8fOzvaosPzrb8RiRHZRmUBU9R0Vku
l8GZdgtRMqojH18+aEggF/lhAFcc+yYg8rKnmjPG32JuG9O30NCyNC8VxCOavlH3
c9eM5jhZN5RpkCAYUVRoyUkNXOoJtVwoi4jccIVhz261NlZFkB4ILFprjNwytSF1
gxrq2TcO7aeAcm7xozhMNxVinsiDOTlctpMrN+8Z1k0ftFDQICkSQutJ10iTWbnv
Lba65lI6vrlHaGApeOCmQFqYd6004axgrxJrZK4uvA88nke9TOOiD08Rp5KLPITQ
QP1GI0wkhww55C+bGQWlnk9fMYNwVO09Tvx+XzFH2vBYiFTXyjtARgoA+srUWe4f
WVW75PvfswZ7IjFLEBaJdo+qaaQv8h4m9w4+JkYEtPqQgzK1md6oneQG4yHwXF5m
UgogI/MRetcprkGNW+BgazIc0SmK7ecJav8baVyIu9snfL6lXcnkReR7bpW8FVvU
YZ0SypTV1tN392yD3P2mAknvI1rahusw2Z8cmreNj8aiSrOFIwLggcCIcTYnuk2g
8Z4wIEOYKwVo7N4+qeQQjSQK4g8ds58apBtyCKMkglR1X61suvF+rB9OqAqoeERK
x/VTFXyEJtPIX1XM4XzqlO7/qW72NvKxZ/UVmuXZl4SZI3fp312o5Yur7lvjHgTy
oXg3N6TBVOYGtDuWCPDX6HFYbB3EpX796cOBjJuvhnhf1sTT9PYrNXYPJDIfVd2V
McD9TSfwGozTcBsc0ZZJKZA+82eQ+S7qwtHkS5cwng2+eevaezLZXcltrGYl7WLC
UllEsnDkaHjKQpTkUMp4ZughDu6wqvw29y5p5/I6wz95lgqvm/NYU1uLJg8bwm2N
ukiZbpCcymDp9hMb0Mu5I5Lche5bIlVc3I5F9fgVZjMMuMrrXPX471Nh/Fk4tt1m
dozh71Wy98wNGI+sAJXRpP/Dfje7AGMQ+5a5SPPVKbkcCD6U0nKxNBG0TqURMhDz
e7nQvqEo0HzoZYPnhMWMpTk6cQP4Y7I+UPK9lp1Q3fNYDqd3byyw5JtldKFTun4n
xKwlLB4aStIP2qCjmEc4FSHboWU6vpK7e1AawXKBaQJEXN1utt1F1qbAq0XDF4fU
Hqamu10A9L92T48Jwyyq6mTmwH65BHUwNbof2TOlM2Y+XmQnV02w9YalKf05byFC
KFAtrUTh9DEzeVk5W9MCA+YPZdsm7ig9agR8990lMowP/QbaOobIvqyf/MD32G0j
31vf5V+xlscLLH5EjGk48onlG81wWngJzlOHw4H2esIy9wR8NcmJlbDMRa6+4z/R
NvZvKUkyE9JTvArSCl9k3LDFmK4Xqg6shNdbKsg5Q5v8M3mEU7rp48ntmROjWLEk
FccA5PkW97SmstvijLSedxPHVKZso5XWxnV76MBwlGCmoXi1lhApJxCduiKZiVXi
IsuPNSSYo4oo4O4f+CTeAlASXv3ygAJnZPj5nwLAnEwKnMZfHLpBsZdgETDmU7LY
wykuHg3zPVYHwB17e1K05iit0asxER/hwHhNn41dWghuFWuiUE2l7O5IrxlDffEr
6xkiC0BGEHeTmRrAWINZ/HMRuUFFbfx88Fo0pkFPlAzCaCAL0UZWJrtGAOGrPLUS
TAJvzzwd1df4HPLVKiBOLen7e0JpPruWPvWnFCvV5ZaOVeqA71AvdBdUaJS7IeQ6
i1UoephYrVnwGNUUmfYk+rTHgqht2gLcTNplTyWODSrhspbUXhuobWjyKInSNs/l
g94XC7ZiMJrJ2EittB5Sn+20VPLTIvupuABssj9fP8T4Yd+RcsEtIvUKG5Apx2nw
VOZQ1iz3Bw+wMsO4jvtae1FUtd19sJhnLf6u+qAcAA4Lb2a4tk92WCZ+UzauMhM+
lJNNYuk0XPfYbvZeozkGi23inX5Sr4lHy0tv9HmvHaA+owD+iGN/FL/I6NbhO3q9
xQ3eJ3a5/kGa4lNu190e0Swg6HfyIoZ8RuVtVnK+8xaJISl3p2We/dqu4+6a7LJo
QUnweHSmAEUZQSa18kYUkpa6Wdo0peXo3UXL7XVY2ZUQuiqBmUPME82Pu+t6emvF
w70rpH3q2WJHtWagK75TEfymoAdWoc6zODv87VqnN9KgkCXIwmRIYV+srzwViJh8
WpPT3dBBbbmMzA9WzFJxp1HkjRwMdUrPk+G5DxjtEYmkMJ0zfgo9gMM43UgywBsc
AQVzv6WyyS3oAgD6+JbW5wVQb0RPhFOX26wGx8Mys9qqzRDVTskz3JeuP7+DaN2H
3JKZtvPQ7yYXLRGGt1tl83oplFAcR2e9bx1jX27LyOfCwB30E0bBV/shSjbUHELB
K2+joHjBq17kJjjenpG7Mxjt3UwSG9mzqU9QJlbqYfoj7o9sITAzPlteWjYmy+bU
lxzFXQuZFQjoV7fTmiGqVVhkvB2th/nLbP1WKdqxchLZa4MM/1MLUuOnECGo1rih
54ix4qxQLBhfposzH5oNYIr0BDl5JrZwi57Y7dK3nc0G+xp4uHY/DCKEVSCfbpHC
LMQEiJuxExcbVL0mkDS7pPSuWxA/iW0sPuTUUcCq6++apn9cDvHOq3VbwP2Y5O5P
6dT0lGfVP+WgcoYDV21blwgNp1fYEsAaA964BeHAEa+5prR/zNY6n0H3JU0YFnXQ
09XAjoxGQYouqD29JC2/UIEG65q9vitW0taKF0hazahZT3XEOcqT3/MictRQyFEd
E5vLikFUaG+aJLmOcCEGLL0bjQdqHtmJuEs2YB75l9inO1if9jUzqUe1sriajPe4
F2ad3vLpOjSoDv7YSVCQA4Wr4HtBp+2m7zJkx5R/t5p/bgABpxXQWmcJzfeIhAaF
wIEdQK28Y4sScg8CcbYt9zD1kwxtYdquigJVUZNDnJejXJ8lfro2M+yCLMhRXNFm
GR0eOa1nFoG6zAQ/EoZTtvuiumgLFlYO3e9+yAP/F7PX3YfhwsF3GGTu5nP7ir1g
MXENm93pOhKVf3VRnr0ho+9aasj+m+lPXG7wUa7G7cWOZ3t64jTj0HYLYyXhTvDb
wlAOu8bKrBazhXn/VOknyvACoj8IarRWgFxhiUui+THTZ4MAHB3EKWkrJD0sSiY9
OVjZF8f7dsa4Kc6E8VuyzuWzfgQfTHQxiE2yzn7Y5bpgwMIKPERbNLGpPwERaist
EyO5gmX2viHlhxCLQYNRcKdYXjc/RovkoZ4OQSnm1TYIQaUL15ASNnni1JwpSfxj
MSHKzJBeP6njZaA+aZ850/+YDY6a9f0NNZiThCtvFpZYL+FDIxmUxYTT6dHYENRl
7iIMwRo/Z6lUcKmM3SBDQIvqfZwyOpaZeDXA9RH7rUZrhj2ma6FYV6WmMBwkG+Io
b2yrxqCKXHOifUt9WNQRahooZctjrQmtrw3vG9+gBNoDmzCfNlmShApB/mXN2x2Y
j6uRLovgTDgJSoT0fWL6bCtB4/piJYJS6SWeWNgeAbjahGZDo1fNy2nKBTYVGThv
fkUTW0rAfBu1n6u7waDf5oZALnkw20ZwISXicxIaVB9bjhgwPh1Fa+ZaiyuOAcR8
Eoe71An95ylHQno76R3mSoQ6WZ9YevlrUO/mQxoxyk1W+yLioc7w6+JOuX2nxI3o
dFbyhmjAuQ2eOQS2WNxx0t6bS1fOHxtwiaeyBrp3w52iAgpm1JbKFdCbnhV9ur1F
fg1e4rmuqXRnUX+cQs6JFq44kR4ln/FH2mJLLkTYctaNon3xLXgiBag0fMbEBn/Q
SFjRzavXKHbVuPufjYZiFPMYxPLWdqvbfF0nJUFPtBmiu5UxPWLQJ+yCzEDxYGLz
k2776TI2wujXHsBUygAu4b4ReRnpRiWqv99+RvVTmpVFbUGaBtskv382ofUV41gr
6pKmDo3tZGXM7TyqiH0uWKQQS6AdOQN14UbZyW5XocEg/obKbyEBMwMstIwbL0Yq
3mdfiF1McUIfcH+2f6EVyhghN0WGZFUlzUWEFvGTSqFJnKF1i484A0BdSItqNDxh
82EWSr2uDIytGSf+Vx5xlwKb8gGBq2BLAFyIpOCQsdqWOfyacbivdzNoszI1hNTz
vxVoKnSh31jkN7brtJcQtv9LaBW2gXcRb6SOBlSkckP8iBhDYKkusiP9+dCHiolT
dqCm9PG9wqpK/PH6OUYvUDv0xqBmSyisZUmGi0Slsux+PrBtBsuxg5Q/hLDYlSsI
x8EU1ECS8jZYs/7+ujjNfaJUgPSrjMOamt7516k47x3TYxTEO2Cr7N1D9LHcQeqT
IVR4JJG4o7u9ulNnah93yNwjmMib58LLo25n/wJISLXh0zLAnMxjuo0aUfxzSq0L
`pragma protect end_protected
