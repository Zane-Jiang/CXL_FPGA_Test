// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J8z4tOds2we+/rcUUywKNfJPwg6vLPzjUeD4BzEgQn8Mh/8lJybxO2PDfGpQ
eJ8WLNiLUjFaNlAm94VTMB5wgFSO+VqVGn0Pc7JDQJ3A7fhkPiUSpsEZF0xC
feuRAHalKPFZco6cs3wb1HKYcFKn9OVLGjdVKUQ+sG15Lbjehk2Py0SMMqPz
qw/B7N5OXA/v/gl4Xq0LQmtEz++utDI2YcLtGU3DSMki2Mhl1apJwwi9DwWn
VTBBEuLffhjCP4rNJvFOFjMQG3Szj5bOrU/UmgRb6hu/E5lI1Zp0cniRtwOV
xgiXVrgdDWLmgNl1V7EvK4CUv/hOzhpQbcQdgWEYPw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Uh55zDiVLGV1ysmyQb9Q9pfshhoDLx2hMQ1FvynKtvZVa+HsBrnpHTqIYQ74
lxUw8B3dlZR9+kwSRL6NyNebuo2rd251uI48/Vmjoa2I8D6PQE2Y4kfbRK3L
t3DwUZOzsnFggMbS4kv7rI97nx3iuw7v7tOp7JLC1j5HDaSpQqpQzN2hKICQ
OBXHQpO197/9epiFqlOhLOrA+9MQ+WJKumoLqWL9qv+Vc6bRxdnXnWald732
HJ8ZbeRb9/9Wpk6pUutnCgjaveGCPN71SyBosEVvSYMdf14bouiI/hF+ApTE
agUgZdDcExDoMwa8b5TAChK1l12bsi5JQtknijVwUg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Zi9FTdWWUGk8tBBIBJoXKWLO8c3w2vwXw35oqO1H31E7Y+k+EdP3gcuIUf99
ODHPdhY7kGypDENzeQAdEllCj3odI3g2loiC/8In4KgW5kM3/x5xCjVwTFWM
0gAbm11TD9lhOk9Xxuk0JtoSf/nWD3FxQ1bhp3Tbi9h/7F/p5BXLQpll7x0Z
W9Rr3FYxaD9Mmma9n+4uASGlyGcoybCSqE0dirNUMZsh28mubFEBFeivlMxA
KCup1Qi50vhDes7ku6Oqagul2bpuVmYxzbxn2fBhpK5k/+DGfYZU+QSCcHzA
NQh/3hZbTxCEef6vfJFwSJ/yE2tHna0CfBKvAYSY9A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mtbf6i5/9gmrkIAv3yLDAmKWA4LNpPBXM0gwQZlv7sXgpjHtkK6maWwLuZVW
FrmCnEBuJTacReJ6x3zAsPCCB0XmSWPqMxfP8xndOwhQwKECEYWjhz0W1S/M
ps6mZCeiN3sGeobkKfug9952S7OJ/vM9BJ7x2vVam9OQPLBXki4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mpXdX7yXPxL8GI2Q2XkS2nvMaSU6oKtoIwWhrvz1R9aJIiOpYj3z6yOYeTyj
WX9otOX5bts8zOd/vOes7IArkgwP4x5aq3OaYnDNlKgbrZn58Bh7A4mbhzCF
KLT7Iu5c3LLGD2i4vfAuPOT2oQJL+e5P/pkbmK9NyGJhu7s0YzawvLjkEy1E
TaC8Pd2holqwiqi6X+F5JCJohip75KhVzHTB6f7IhyjYw1IJlld218RhbQ2A
bdbczVuAt+4zvH+QphK05vvycySuPGDwiKJo7fPgADyrHZ0UU3iyxOLIew4X
6q2sg8n0xB+dqpC+lGQiVhssxlCv4wz7mVKvnsvLCeJPtLS2a+6k668TGa+R
LGXNDf5L7LUJtGKJWq5cA1bcztt6YF298WpwEdLwyyJFSWRFJGh1v4YiQjK3
s40cDrUVPuJA7rfp1IwNf6yJO/R47ceLnrdpmCG5yML29sYB3jkFzguzW8VH
4quQAM8toNg8+3cdXC0IFSx1dS7uMSlx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
inBDkmJVj6VoPCnu7goxZ7y5uf4+EyashJDsCWfPxSyhPwcJQ9p6u9FTfHJF
CoiCFuD17X3ZRNho2FKjgFcAx6JGOJdz5m1LLA5MtbuDtHbxRZ96YtZ8qO8R
jUy+2sFkU+ii2+Va1H0sMryghI3/REaIzNCf5Tcf1C+WntM8GHE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pfucXzeKa2uoAAVrV7yUg8crEXZ5Y2i9S3iK9vRcIP903LZIx0+BVgXZx98x
BXiK7wJrTfM+wM8Dtmnil/WtEA/oOnuYi/hpOMw7Q2pLEWE4MBZLeRJ+i4DS
qtef1rq4iQWc7hpTYe1q5hF5KCJawz9FIAw9FpAC/9y6Zu4mF00=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
Lkh8muu31CSU4ux89KvYzbXsUNIVzROx4C6IVKefEdlzlLXRDP7eZdTdyusG
fzq53fhHoY0IA9MgoHLhj2uyf3K8Mk2OIDKHlG7MxYl8A5mbJoc+AMq8G/s2
HBpCdX7KV/pRJhQ5eug3otlKd/MIBisFd0R6cbM7g0TkjNWM5e7iaZkE1k6p
G0hJO6J+iIsyCHP0mruAMN6ayR4dAxe8yVaOlZBsc1YxJxJzeYrKah2nY9PM
a18dvehVXEy3fhaG260TlMpSY7t8+Pzl2HteTOlTDSSdpBrEJvE81DnIJkNc
xAh4E9pylt9UHknSBums94+L+w9tb0gK2gRX+7ELNA2L4ku1mXcdh1hIrBun
bzNnMTr05oqOpNk41N14PogSzj0DDVaeD+q7/h2cmT+s8wXFIyqGMrrfEJaE
OuxNJx35oWIslvmNJ5Ev/R1z91YLdp7DEHv1tfCIIV8/StkrniBjOrFpHWZF
IQjsik8aQbaA0qWiU4L03iU01GlvXLoeuLHZZa+xtx816r79DznrSVo/xgVL
WIBN7EAjtBGiuGbakSTqfslZSrF7RjMgrHZZZNM4aZ/0X6p+0Qb4xpeYLIqY
rsKrUsk0YGvkQC9lgMGwPa2X2YtPoOCzWlj1A1XpkyZihhAUSX+JQlwo1C9c
67c8aKbad3sLKmUexuRaXjFBdY3yADHVrLnno7WFih6G14jPlrH9yI/ZBOXl
CTHZu353RFMHXrcz/odqw4KcFcga61GNjKrWhKQezxz6Vn11acZr/XtZQW1D
dAWeh3N6+VTuWmqHZhYBerPv3OEOTHMCzqMsA9nZh9OFpHITnkwwAWwoqF4a
lqI93nQrnQyfr5zkMMk0ocPR8TxNaAf0gutjVam3YOrhjdjCCBfPRghU2qm5
6YHSDkUtYkRjojTQbQqN+1fGWRKnlbOFYIO5FYMiGk7MochFiDXekA3mjz56
KNL4jsHIOOnOzPSY5v6WKfpnnAbsaVNlMdOaIUS15Vp+I0I0jETrSFV/Gpp+
C5/5+m9zgDGGPWBkh1rpujRamNZnhs49QLGTqWWOBC5KnNLNNGYw4WD9KmRP
C3uAlge8t1+fSto9MlaSXBn82/T5LxvKmoisDAZp9dxXiAmkOSY/MfiAeRqi
L8p932cZJqHAIKw+zRjd17hrIzl1LO21VdbKIXn7kP5eTP6fXW1rTumQHkI0
FpSo4/CEYEEcueeOgtNWDKAoZTVGuen1vzo3Lltm8t0Cw2WIjLMs6jzQA1vr
MuWAFAlXKhiLbt01V4Cr3cHo9Tl95Hxr58R7pp+YejGRzXciReW90Sjhrw1v
IZcdIBvyLidfjaLKTvWV+YU5Z6qa63avLEcQVWMPLtwoDFdFdTmpQ9FLB+3v
u0lazzHU4xNTGwl1e32OOmZV6QhcLVlNGxZTJVsmHyUJ5lRu0BiuryT+DUU+
BEwuLR7jigsV008x9uyO3+rhMRtuYhVGcMziN5fHssz17crd1ocnVpFSGAel
ymaTWS8KokCBMisKiJcroDvlKoGfYX04yye8yAUMYDAf8RQP8CrL/1quKqSA
oVHZa3Nt0Rw6LvKFtmzLbn4uWrfiFGPNm+CPt7kNua0fpMzprMnznCjh70Pj
vs0yBKsvGdXMUWMc+0L/tsslaNkaAPqhLDpuVIyPljrA/+r0NQIuLExGgzGu
T+ffi5HRz9ggrgwj+YlRcEYfsTRtkggdeSbM2jsK54p9ZpN1eVQEiugNgB26
saKq6GfB9fKqRVHby5ASBRaCw0hlQxVKtpp8cV1XIPvOkpbCNQpH+9oRodK7
R0HjHDMliXd0/Ln4/jwOO6D7V+fg8z5dNyY=

`pragma protect end_protected
