`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
in0S/wxJLoFEf5lC1Y9idv7LW9kRXSLELN8LCHU96tr5JSgML62aThrC1nec+iU2
CHzeErT+1kpMPb0r8c35k6yfxJxDdG4FWTffe68bBJ+6B6y/bCZCtLrJTrW9VEcK
iTlvoDIjWNxKJ17QesLkf5JyLo6mQKICnDpevH4VGcI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 28736), data_block
UKwERBqlQhSeikoteSfDFhsxRqTV1AYUPAl5qkDi4HxmHQOzA2oloVyu0u5dTycT
5JApQvLeYZbA1AfWL6ctCy79pwDmTUKYs0cCSD3xdSbNMrUZlKwCSxQY5WJBgA8d
cuGiH32cnZuvxxfRvPx7VOHqXyjyea2OlPW5j0cJNd5ZZnYNMxU8e9beGXxvVExI
XG3ur8CpTZGuDsOr5k/ummUW+EKJIV/u4sjF/1nvw/Yf0LLtyNAa7IF6jcHJ7HXI
cEONdYHANKOpE5/LCaPWIwugxRPpDheSPxO+g/6jdOwop44okLNYsNTDJBPW73UU
vIoPIZYVq20sz5TMY5HZTrCt/pBYFbnMErmqHHqqaiIcLFqW4clIO/vRuxW5vD97
tt60+sioDpTlS278CVCYL+ZGXs+y7P+fXR5foLJm4+t9afzu2ssKUpDDVQa220IW
NnXMWw4dt3XPCJzhqeWEX+/DknMAwhPyty/PVitts6Cnb6HpZvsGrJIaPnVz+3Up
NEAE1pc3LDNk5qrJB6z2UplULAAlwMmDfWrEO0/KmCw1UkHB3HhWPU++wlgyPwVx
sdZfItAKM8kFy8aWg7MjSeej58qNo0M/GDGhhzsSUMGzvtQXq6en8jNZmOJBesaK
b1Amt0rDo9do/VFSVxAL2YxxtJAdP4oZlJFRHXEyp1zrkGrMZS4NtF10ST5ktR4q
2bAeMs/CxLejhBljB8mO0o+ZDxFHNEtK1kY6HBwBLimQpDAwNAX+EsX0PNgtucDo
4i8rxiOFPFu09bjPTZOzFrI4ibL7hpOYQCjdMbeZ2QvzMyisBvIiihGZQtwqVXJM
HB0n5Dy/Pmq/llYdDJEPQZYi8+YhMGUmhKH07IPR1nP7bfp+TqW3SZOcke9KntXR
I1+Cg+U2ncA2rk0UZCZGl52YCvezu/h/UIUx85Q3uDguQPCczpiAN86Syk5m4pGJ
i2s9Z73EQLodBL9cLE9k5izmwQt6BkZ/YjKcSvqUKaZsE7lLu92LdGa3DP51SDHN
lmx22+WiMxyGZt8czEPYhqKQJes5Mqxj/xIXTYDbg2Tj4BB3tibweTUNIMaVkVm0
xI56hoHi7XajO/laQH6qE25h7W0Qce1eAIn3Y/atN07qqiZY96rMyerQUfm8oQvj
RdxdbxOAegMdSH6kmwqvct8uMljLL1Z788v+vn8jVLRZPg39AVxSodXyaeHmAnIj
LxzcmbBAoiKkMzZ7gPbapUGfwLZKhu+KLF0i6ASaqckN5vcoAQ4EtDc8NmOnynfD
cxhxJIgG4ZnXl9uh3zrMPZP/sGmbQu70LeZ8Lwddn6TMk8A5HIyOIgFfeKSjCkYB
BdHjGOmZgo5xN+U65J7vScTEdHzy1PY2ko7CT7l3TVuT+X8H0MEcduoPQL2T0JUr
enzvRZN94lp1c+1aZmXZi6CgI38aHJVdF5m4j0/7iK+s+2xayT/z+3yrhXlmHm2t
ukliAlD/7/qoVbyrqF9KJyVCcrngicKz4YNcoXSBKkx953kzLLAW1QNbhEOcY+aL
2vztyXhYTiuMkQIv6AoxpnddFNEvnvexBQm3mZDSO6i6vj5FZ68dFCUF6dFh+/Pn
XPSHpOA/sGyNh2hWQvxpEFAhpv2U+Wh8Lj6y8xYW4OKg40ZIBxFkjYhy+kseiHu+
MDBFF3JAJll5S3cBXnVSSyb3dG0oQyC5pfrZTlqThqWSWUnnZtohrlbqUT1m4I2P
XtuzFTfEbgPd2PRTAWTGP/ZFyp5YvKwjBMlw5hS4uGfEi9f7o9l85BtqZndvXXjl
gdD2el6R/pdTdSKL//e4KT9X5dClRWNhTvaVWRbAv7WZHn3fU7JQDR4hYyaB64Qg
Jx4JyDCNyz6x7jtJiW6gGxQMYPwuaPYipisktUkSjXUffXKe6VTdsS8Pd5/w/5Zf
FjlOUmtdQDWxDLrUVK1k+LVJUgkebgiq8GkmiHWzOGTK7bZ3aTbAiaD5ZhD9TXJ+
xnC0WQ7y0jw1mUJtZaoEMdPvZQbK70wkulfDh0SSajlsTiscC23ReODUcHl9qY45
qPMrdGT/67Sp8JutbD0ujJSAhKUt0h21bu4HrEJWt6kdreQYMn4t+28xqjO0meAI
yyRNPl+iCMGJ+CIXLi7wryRLcd9f6QY2tV1Wk5WOgq7DEajo5jAFRBOuCETPKoCL
WmKCoK9EQYStNXyn2niBz4BIu2pz6bQJdNRbEJd8pYzowftylDWW/lS3SXU1UOv+
Naklhq8/4b17TgKRUnNAbTFn2t3LXDInqidRAmdFjkVsCKoBBwx2HQBGNBmTLKGd
JijO/jWH4l2N5jKqbxFGCnzyjHv9MqEdtJy5O9ie2JITvZbgKdARKwCjGIzYfs6z
0l42HkClIC2xCDbBvW0UpoxSeoODXJSw8KyAVm0sJ5mwR+1yPJ9y7JmyqsP9SUhL
JsS+xbzw+sv+MCKuPke2/f4hWBuav6mMXJpYPX40vd9t0OISbg/c9d7iaDvGKRyN
prXG6nAvQV1kQhqQNwJtsKHE9/SEGDrdVl//8p9XhrH5UggUtlOwYrxS5GCcgEx+
haBl1y9X7W1F3FkpnYzRImkAqQORMxqVelRwLUQdLUcM1+SL9FVEDI3MTtwLM4X2
XqxPipGKbP+85MXttOtb4k9gagMQ+9u/zqxn5yoAawyBOiktczKlq3MY6bhU1Mwq
Cyjs/zM7ddlHQxOIsmnrsm8vuChsm9lQB4X+phrU9jEry25vSrcg7BQP7eiq7qCn
TMmtjJZuvOooGXpz9tPRMM663jZ4N58iUj+4tlRKYZUpvfYqmFUwtVtCrjeggi6C
ttdws3vo39zecf/tYmTwuKM6IFWrckkEIPnJQWJBHREwoMHlLMyyGO234SmDBnAX
+a8IQBCJ0gDj+r4uuq9/z0vGhc8cv6ugKx+ctlyDs6ErqQPiABxF1cxjJLiAXiII
46vUCogUJaLVIRR/mAVWiOb2cNIoOUti8iAH0XsOhBGAhJHZRnC4MZ/OEoxBTVzI
G8skdmf5XLiiG0BRHwAng1gNyc8jjrmsJyjqjNkPqA+QJXcqaeFQPSwlq6S6+8KI
f/QMwofa+6liZkdsU6p9oPj3beqVB2dI3vV1csqWWBwGC2Aqo2YM3/3iu62R2p2+
MNMbenm+D5FMPjBVrtO9RAPrF11TlK1SzpH5yeVHr7voPQN+dFlAc6kXko+xII14
K4WTC6Z0VBsq5LqrCBNqfo7VA01qdg9xM76f93R0+I/FvayVVyljnwcy/QER5lOL
iTYnpaL+H4ohqngLXtAT3fC/hBxYsRzK4tr3ic4Jbi0sXj9ZzC9Lgk44DqLsXHH1
ii+0Jowiz11VOM9UPhXzNzGYnCoQSgdfk4upGcnJTOla5DPLppWX02LFjvGjbcTF
NAO+h0YXYXg2p5ziOZztC2zbpqTqf4+P9+dNNqLZB7oRcJOVbjRzqRYCFRxpIwe9
VvM8oLCoj0bvHknopC15jIDVoiGK2+FI+c8fhfpb2Ks4E+gyIZUwbsxtyhdXskMs
txI2v8Ifrd4K4jjIs+O5nzZKX6TtfseLywi5BN7VnE0x/QasynqfWVGmZt2WDwDY
JXNW+I4I/vPBt+FbQto4Fz2V5xUy/3on4oOLV8szC8g7J3Uh8rzI36HZL28lQCng
I/bqbxoMPoSyGvTX9DQH3r/WN6k/at1hm7ddO5Z7u2Eqjra6qEbmaxMNvaY81bz5
uLcfcUPZMt5ucTtyJNvNqpaG/0+H4BqeyHlMR1vpw9a3DP9NzEapHaJbm93pllLP
MwPrTOGNLFjHlYdGSgSIX0kilBeK8UVpgdlzFci4u577oCU8Wdidl2PmUPDsAHBO
RVkN6g8rMBWpIYeMkxneaHxs/n0baLSEkNsusapU5ZKe3JRkt7QexZWGMXaHHsJ8
EhQ+GX6eQHTZy3eE/FgPKXa88DJIg8VSf0x0ZOmUdZ01Q0ICSgPl8+3lGugQtohr
A1AoZcmkTfIwA31h8GHseEGaYDNy8Ccw4X7jL0MoC/xIE9abpnR/8T1jPOKqrhcz
aqgBUJk1n4KpxK4UgDwpPRZ1zQX7rNJEXWrQlN+MhfxqGB9Q1wmSPG8wHhhbXH/+
nmFUlUozBiI1aejC8gizOUfNpzhMbqbieA8Oj4c/J5hvqRCZmLqF3hmVf8JqihDu
HswzNFU6tgMAgxPADMyaBvVcG6Q5QjTU6VbX/ocfepuqLc4mj0P42OFCvUHKXo/5
5JTvFG1l6SC9yIQTyHa0EvTsoMoMODX5+JrVZQzuT2yZpamZqYDnkEf5dOPx7FQ/
63UPR/M+Jl7oIiRifK4Ho90Qh67YPf1VzIr6XmATgBQ/T3hgTw3tI8TMG8mQwtjX
6M3/9pYPvErT1psg32hlLf155WcFP5A+3CmKFBettdS8XA8kqiEsNcVzzeDdl/R2
uYkKKCAMUvj5gibMTRW1sW6eHHGW7NdwXytwUrH2NFmxHrd/XuGjimflXFEuPodH
bqM3rFnX/ssJxjHl9I6xeIYAu29q5M9Lo8RltL+q5lxlAoew3ISlIXhbaJzUhURe
mcXm5UnS2v5ZdU5oWkAzbEcJ/YhwJzeqije4F3SWVrMCGI3FFEuvpJmeeoBYLo1O
KcyoU38CTdDMtrEC4f0IKLnJKS8ULhO7vd20VLHVlHCKEEXdvLL2Sf8K6XTschHj
EuuEOqDx0V5tgUFrETC8OjRsXLI7QmiORtkxHpsYb2RyacGKF1/h5VIDYrdwZQoW
UIjj1voPry8JKNjA7VIH1CS5ckRmrWu8ri2qrDVrcf7toZ0lQYHSsXlbwtKDEKIY
ZQkdMensF6JrP+Gyb8twHNX1T7h14UPB0G+oMfDsekmFvGiAlM2y9o5CUmz15qhD
L+NP6J0Jstr8kMLrg7DVNCvbRQSfEDzEgUw28rn7IYZ0nxdQbB7c5L8Za1qe5tlo
MPb9+Nt1fp5HykUxLd2ZHUMgNkpClKxO453WeLUJBMlg0G1ZUlGvNvq+TFy8YjsN
CmN8fhQ4tGB/dHmdMKSuuUvYVnFYU18gzhmgRGmpbS+6+l4Wu4l/VH80PIXt67//
VftSpkwkyWluAHgb49pvxUjw3wjOYKldtABr6mXUjlwqW8qsIwp8e1W9WBKyOz0U
z6G7bJ2JpbZ1OiUDQsPqVv0H4i//uKOlnolAyR2+gnyhMCWcY80LK4BdVczDfqCW
wCkHjD7ppKo/KYBVghjxwttU6UmrIXvzL4dBzrz4fW0i+ZdlhiFnzc8E46schWoY
JadNLpeOebYe2/o48HUjs5Sp1qxAAoXxF8L2XhXvtXPxDkjl57UYnD9fS8zQDYjZ
lOhOYCYXMqGWwvV+44VrFGwxxqOCHkWf/r/Cb0vPnyZZ+xz9eXScxYmvOFwWr32s
VmXviWQHXrqYI6FA9UCTY9bkAYwMVu7LRB7B2ImzBzYJGZliL7hB6nqlwomaIsxp
iJ0VY8AAzGKbAKMJZq79OXIbvkjz3j1IueZye60bjrWy+EGBKW4qJHucVWFrXdQ/
QqDk0dnGMlMfY5xlY2W0X5HIfXjfDqgifv83derYXGeHW7pCRW07CqAUwTjxEsPZ
PqF5aGp8uAqeCu5iLSq9KkMmVuHczOLLUp8chUsmgEOH7Lhkf69ycqDMfRpgh7Rk
rYdZSJUVhguhgJEZc4meVq/bXLCl6Hr0SZS9xk6dQf6zxBpaiyiAQ7f6vGGZ2+aE
pw4uSm+Ohbi7N3dE3DXf1Qnwy7BQtSDjx4mxtTKKBij1Ni1nGyV3SC64MwIJ1/uZ
r3ZGitGeVRODusYuWR378G3TyrSlqdgTE8u4aUyzTdkRt6WUrfhgLAe/7MlDUapE
rJ88VcrvduKUHBVXv9GLcsJaXvgIewxERrnwJMv7mEz/D1VwKxs3OE/68bqmHcf6
qHcWDUN5XI0iTt3SDxfrJJNaGXAIdJXxlxnxFAqSETivtxJH4Eo6HrDLv3qXgKHz
0mTjnZHAlE6q6LgwO43WQFSJo6Fvs9nV/wkmSwY/DPywX41IEjKoDWJGPvCtuMdL
pCRa9bL2vcznZvhS8jJlC0RCQfwRKLkGlOtG3A0EYzSccDYe8if71hXwyhePzY56
y23CxP2P0t0nheVywqVFDBdjPzFZVZatb7fYJDefdDtXRDwlg/sGbcLlYuXoc7Tt
j2G2SsEZxX7HW4vHLK8PlKJ3grQam64AcRsjXWIPSAZMziLD42AJfyV40eZ6Jbis
2T+LCIWEepbuRyXdEvlMbxvCP0Qqi4QSlcEadmCpGMipoqbj6czRv+S3DWe3Eisw
HpoarIq+2ZfuDyI2Zm+bNfU+/WGlTIxGuSqDyplpCSiYZLgd5BCtmy0n15qWOwd5
okd2KlV7/BodPmQbn5cUG5Xv4lWyUESU+P/skwpHDFDy9JPnVjUuWHXCwwrIL6dX
lMK4tQceIHtar5h8gazgBqhksgOB+xEKse/x0HYJcZTUIVfBw7TywryAfMmRj+9Q
niWwdOAJYFk3wpYBG5xK+7OwmOa+W7PmZbItpU2PdeNLHslU7YwtdyRMT2lYPHBb
d6w/uWhU1AJwkgbWbdKT+IqLPwwZKI/8IhJSv9WffuovcGkw9+f/1RkUavKuSdDD
8L6dZh7DFrAzGDnUbuN1iYzjTUNZWq0/QJLgNGBzlCDUlmq7ZgAuQZ0DdAaN6PRG
Z/IWdL258zHAo2gH8/zeucFlDmYvK7r5Yp75lOl/xT2CO34pQEUYXmLhr++kMqwR
w1G8c+Jk+kJj8K3A+tpNaEK6cBamTlpYVMHwF7O6gJTgJ+oav4D1HQx83DA5B0Jr
oRypZbFUctDDJeqjYhDQWfrj68da3vM/zOUtM6rLA23VE2XxdOU9gXhgmZcTr1r6
k3A9+vhjWWI+meMfQ0xtWIjDFSr6ofqgZcrVBc9OKpKoHqAceiaHMfX+LQA6cH92
M+eXG/DbxbEhtIcCCZbAWwZgVRHHm+afFveTofeALkSLaXNbj0+6r+9oPv/ZYJlz
Cdm4FXzKDCmzNLEW00iAc+WU9uD4yZCxlM3ECk3OpMoM++dMqumUPQH2uazoWihT
XliW0R+WsOuNmOn/7vG1v7ymw2e73jJ4x2cUZNE8gteGH0Vqnw/SCNiJV8S/kv8u
nhboCnbbUw6DzpHrfi5YH5OLus8q7wDLhh+hjuY2l+C70Qnws0yQAV2yEQLeIaeP
Agx3wTCC9HxM/UgJIwwyhpNXOTE2g+nz9L35+7nu9k+4Sk/zRx+jFojovFxCfk0f
Mec2+yYZNvLkDxdOiFMBjYD1zQkSQrRkrG78dyfGSE5mlFJ+UhjL6XqYSwZEQbiv
H+by9XTDFF77X9bMi5tGI97/WerOOcEZQYbl/ULQlwsGQkzBdJiN8TGWNZAYjltr
R33SCMc21OR/EYsx7mjVL5wOokElIDBOc1ADgQHpiLwrWWIbDRAS/0HkdZYPy5FD
UIod7PcIUAkj6pUsmDFX3Nauguz0VtjIQSERd4kFhMcnoKUPA6/XVGLsUCfyP7B7
DHJJCo1UVDfkrrVZ1Uf5n0VNpdqrBVO207NWegXOYp7IvxOjVHleZ9mdLry68832
CqPkgeocHbhjWKQiWERQpMdq605DcAlqL1PrGbnfJwjuTmu6DKVdIhdQ9HFfZevz
VaHShxqSTKYiryimHgS6+bHDhieGv3L5jZKsL7qb7pihB34ojnbZUiUWMpARKe/q
Lgmq4Ki/Ct7MwbXhD3N9WCdwZXGUoJDNPY41zn4/MizmraWy5sJLvNdOg5lRNfS2
Z9FUj4JmnG0im08CR7PfoSLnJkZk/7iyU9cOqmGgG7y7OwJLJZ2L0A0ff9k83tpX
ZrA9gUAhTc6O9TwXZ4sR/WYD5NZNjv9+J4/lSJPWJXaMOG2duwRvCFJfH4aaKsfI
EY5kBGy365gq+Df0wxziam5x1+WJ0q0XOf4cLJAC5ukoj+IAd+Fm/OA0gbN4PWIy
4R25pAjaDXBc3HOhw5L25xUNx6TlZOLz1MeAuKxROo4JvUmzuXgwq4dQ7Rma1iYZ
Dv7ye2jsuHOsSZQ+B5uo1DuEAhi2yaq3sgrbtEvZ2rJ47WbM69zX9Psa1DxIxy+n
yrtU5S8Z7z/gc/HOdyqxR+g9dCA7JdNf1I0+G54ESkatVyGuwHzWRHq7UL4/cWqg
4wA9YpfHHgjMHOI9q99XYxGv1ypStB3BAnVXBrZl40Ff3ftZFRdQb7HqoFuTaRh9
I7BiT2s2T0e4+3daB25fcKIS+lDPDv2lUdSJqPg4XxhdURTVfwHkkUfTpAWUcv71
BpYYmdp0ynccn8efls1AhkqVzSgLyJc6fpIF0H4N68qvwLiwkkCWfNs8sng+5DGM
GKSSxmnSAC5wigAkHNJczcytCf+VYApd1mJsedeviWdc7m86nA7eOaPnqXOoHJ1l
rVs5iTCl/2STfLiSC+Sh/bT6Ynd562jq2taHiv66gWWNtTfIjTUaFvrRRU3uSeAN
YKbAAWohRBCJwLcImadzTIWl6ur+0JRPGxVbvBFaFxpTzP/ptMdpLp92s5xSgGsd
+HzHg6/ec31dejXNYvZIFkqrffBJu//NPr2UYfvpJ5/KCj8CosfxTbVYNAxOoVup
J+BIhac+TQLFWm5d+vywJzncIlCZgJap5aBE3vZLftyt4jQKXDnbw9SmxVYoQa73
SNvWzRmF2Y0QkvD5bKrdGpoMbJ+xnfZSm/Njp928yONObLpnF8AkgHbcSAqdOIbS
VUDpr0isUEAG69sur0PyMM+eaBUlAh97h4m7yRSuuUEPjptVW86jg2WuPhjH7UnF
3ZRU/tJP8ROCG48dsF7ScKO4zEfqcRXaLebFoUXAZ95aPvVxSjEHLyurFTqbRWbK
FxbknGJxJy5tnJKNUJa8BjzQsRfRFKHwzL9KEkXPCWQ6u8C424/gy5PR0ZZgC62X
2xyNwhfdKHNcD6bV+kIZ8VCNzJUehC/Wr/tMGQuU95ESiZLZt1ZGkXzoTK2ZAzZe
bu143vzCqP05DmLQqlgsYRpQh5Bn1LAeh6eb1UwyWb3F25OCzIdsipQkVmq4DuH9
1ieulnNwhgaY47oj4wVjJH11UKskR7NOpCS6Ld+cOqyYudvnxXkNVF6A7qdmRwHd
0QE3QDX1m5ilxhtOujGGIkztpA/U0FpzZUb9vNAtCydJAEH5f8d3qsLOAzJW1WZ0
eD0muRezltq5DUAkRjWBLdnv3WsjnJXI7IrfLSWAPYwjEpVIGfh2+q0GniRqcQwS
E9aIV08sOSZI1c/0ldcd7f+MWkHyd/TyzyV46Vz2n+8a9MCC4Kn1SAV/NHjIGr/C
HkuC0gEwQBJ60oJ+kCyJgFBButNkRQZLZVJk6H3FTOMdRvPQlp3E8HPftsVkjc3Q
t5SYfJtBIBhLAnpKN5+vYD7xi16OVwMcyq0BPHYtXZRtYRg9y752gkk5vlqwnfGm
1JPjxYkLTIUzL2y/N6ZXaY9gAV5pnqIbUJglgWOnA7TZR6qbruJD8CntJ8p/qRSj
LxN08CKGRwdkO/ECOjoUIKkMYwloj36Jnbj5irE+/wja+bHBgq1o3rO9QT6kEsrg
raRRi37Wgs64+CiofApG4i1EVNPC0ynQFvJaTYnU45oGNJk1lFyJFFfqd3Ybeamd
ysrTK/AHUxtVu16ydJwe9zCmN4Tf2h+VpYb7l9eM4YSVZ6kMZ1AIl3D0ohwg6IXH
uMLTmMk2PWCdJhS6/1DIdWaJ5HrxBhSOT0vW2idmsUrcYCHZJMGRRAsMyPq3+UJe
RoS/bZPIBJn7NlED+Br5XxOVSF3sET1LF58EdVZzQlM2+ivheHIETegPtbavMvda
etvlyc8qpZPzAteb6O4X00taOBqc7uusszGaNhcygAJEy0NsFZ4W8Sly8AVYRAjO
NjLovvbO9Ze3deyaDf6GgZEsWHbpQvWa5JJXuSEaIg4+cc0pnxZGF/H8J88g4nQy
62xGGUjamVkgIBsQvMJPDHEnh2JZrtVjjGcRqa4afacSxmGryYAIFyCtRkQOLe3S
MtiuE4WnhLgGO24ZYO6Pp1rImE0XLT+QxPxLoxdEBwjJxd8h/ZxUXPIbLNXOyaav
UyoLZ0SeBUFacNIInkpKzn+lTJ8TuIvqkwQw1V19c2MLv3fwNBIyHBiyCIHY4wqE
63GY6EjZrdydIjMIq8ARyWH1uonO6AEiship9e/fJcjkSsBCwwyH5xXq6V0zE8p8
zW7NECi5EEt6vfBgPi3R5oARotE2FNY5HUVwAGR43LZJ/n7XBmch9UEt0wE0g8yt
AB8C2qPrSlYKbjaTUNGopFXoFgWMRVCxIcaCDb7C58HJ58/E/qlclt9+cvAtftH7
SI92MRMyPP2Dldg28IelK4SVhAaz58T+q858D8Sb9ziCBRzMuZj2dDwtMTBuZeHR
lbFYW97iLETHHBGGF9uy+1Ya33IWgrEyH6wBbCdmh3aMcbFFRk7nJ1EGMNVcuymq
2QsKd9YlTEFNEcUDVj8HPO3Eu6+/9Jqa9hmiq8nByXXtRpWWG3/Dg0K4OCuNJQVo
r8MldurXi5nY8yVO7KDx0jSzvUsS8zjH6GYAEJPnq6lPCZE6xqGsjrWOI+b1UFMZ
L+pNRTF/2B7cvg0fYFPUJBHZvKwXZOL9NAK+n1sg1ieC/rSpmXihiJngZBOjxtp6
NcIz6kIGeGizC72jOt2g6IGZUo+Jqz5JQkVUDrtIrdE8wM2ln2axBPd+LDZGkgjS
bsvrc+lBuczIjfQJLWyv7ShsVgCWi8UK8/eSXv9AEwNDiKZHlLauMAQl3aUABRXt
lxhF3XcfudpX98JBqS31u7tpVqOk56qnG60WMp1L7Rq2mfOCGmVL90mdGxw0bb1g
EdRuNM7Y/xJ8igmaa4fUlVuPEo2srYY4qIM713estyYsiQn4SgletiO4KCSWeccG
vJyLCpHXxZW1pvneIu1jqT2bpvBT2f1U30JXdKwkas9k4MezfK8vRLQaAPq8K+i2
9g8SfXvqr+LNrpvT3Do1zMQrNouzS584uq4odFVvMZJiczD+ZQqH/R6XRYWwiNx4
pDWYPFAbf1lyThI1m5+8pbgtftAZcNhyndjdanR9AVa5Qs8gfCzkiDjvkl0IWNZM
zxATBj90qGRPJFlUhqyTrbLWVi2+Iuj7/wHfVcKOFRZbP74YOMBtZKXUYVo3KqkL
vXlNnn1dzxRxxVXvhWEKhxAz3a4lP814R3Lolcz45PF/A7aynvjBmBoZiExGQhiS
FwjOtKph81ENwJRaFhRO+kPcu+QcRqAOeqvwpvNaFQeJ7jDtoKhnDeE0H5QtGPHz
swkaRXF9JCENyPcijqZEj5tKZctHvjAE8J+nXinalMW4BtzcTpXsC4kspvnNkzFK
/sEeDQRV+VJJBbJ7F4VyzqWeVOI5ESJy5NkUNYxnL2uWpD15vqR9bCdb2W9bsoh7
M8hI5mPYHCLoRRW6ZzNz6DECmnBdDCiiHuiWSE6R3hluHhRcRgwErkislowHXCXk
gMfGj9aDmXCz3Jc6FSmnJi4gp2Icioz1WpBfuk1LeUxXArgRwYDBsa1PLtcSyYYV
M4gYgZrBo5ITRz6KFYHv+WtcvaLkP3ll7/RffytzDi9RkXBmccJp3GXEKfY0SVhh
uwObsVQVbvl653xrC/5PA2yDaEmeXfn+zHi/NQwPmNDlhK4gK+s3qit9apOA3O/H
whxzn2FWlUryt/2Nr4GQKbS4k0N1k7vDgnuRoeTAsfuCsvJ26HWXwT2rJJhWjWNK
cnP6YgxQM74QXz5NXCLRrcw7PmWnewv3kAo77IRPymO9gmyDHfk79PTCaoFeFdVI
IH9pF9z33XhD3MowkrhizxCrwwa4MMmaQzQ1S8pEnqdyYh3IivbCtUmNr/Qb1zDa
TJVkYjId89VHKGTQn678trE6RZQVWx1HGOU2oOl4Gl+qJ0HbURXBXeWntPc6U4W8
v8Op/r6BiICpBWz7xBpMvjfnEcXFlUWXlVK4MjZi496a9c4SqxYDIGAEaIFcvgDA
r40Y420stM+TLS5cXG1wF4W6L01mKypcYpGLTIrXqXKQPpSmlcJ+s0ygmatsqCCA
VESh82Nb35MCVCl6F6hMMQ8bXTsGL82t3lsotzi0Gn+xTPscqH4oybQmMv+oI1DK
SWE1QkTalPL06ecZ7ZGXY0tzecToc3YIWP56epdzMBdawNYGQzCiog2TNlkjEU/s
Zpd/7S51QCflaPeqH/b+nzNmCxY/bsvdLQuusbLBClsqS3KUcn6a3xzAIcvYMvzL
kdzFlsH5aujGNE8iwA028fkiwfqGfH0RvOUHq0jCJkRYqMRhO/0IjSSi0pR6Yp1J
0VqMcVoF0tU0JroQGLiXqoN+S+FAoQx1LM9jB+9IduSp9hdMk+by+hMZSeKtZe9C
XZTSXUyqXWzV/tNXBv5fXbAsT1/ZT0wox+HSlWaaO7C7UIKP1o5wYODchzqwetJa
XTp54/vBEKXI5NtCgGWyhFYE6XfqtOBnJv2cpMHkHeMFgCFLPc4po2ZgtepdWYFI
sfNBsJCO4bboPNpCR83PuSeEQJLP/Aok9rwpZUPj4ujnqzzsSosj7mmK2w7F9ldf
u69mUmQo4iGkHJ6of8UHmwp4PlzBVGybT0gfDF8M6k9Jam+QsVGjZzsDEvOh1o+g
W1TgEjrkuDq8GsvBvKVIHQChDzukvhESErrZ0BvRdBC2hr/IJqhWvV6bEPchJ1qz
rdhp9gb1y7zR8rMt25Rh4VTxaO6Nm0D6hhK6MARNh1To917v75PTFQ9nfwmQCxyP
tbiv2iomNigUfvhoXOOaGbRZq3W3nyiWIPpE0R9lXqUaH9cYkrmO8Gp7Xs8+QDya
iWbZgKWq8cT+7dRM3MXs0v4gNaGVTVpMn/cfbxEwzYGxEIVLGCjjtNvUFysw27ZA
EnC5oj12Do2WR4cvHj8B6qABSWxiBqnVPkC/S9NCMzMMi6YM5w38RCqYwX86Pf28
DQGkrxiYnTz181s5w4d5zpRd43uq86UIM3lsjwvHDtpWSb1DfIoJ3NYQeHbVS6Bu
xQUgLLJjVVanfuJz91hrsOiJAhOtoKyKYvy+4/k49ZaxRxlOgvlrpf2gqfFm/Tfq
Fv5DTf3s5xGnpVtMwMj8MrXce+5dt6Elr5LDdpGl2oQl6aT+uSH/sriecdE+mw+7
e7qsi3guaEkbdkKVs47lfqfGxQNbWoz1BkSBirIuP+TYjbTdY/l8GFoHkjjY5HR9
DFYXOtX7KmhEKlvroi15l01IKzM1rpdqAgYO29lj0vTtZPoWhHzOLRgvh1dATtUI
GpF2GjEnuO/rYsJ7wr5eTvvgGNaMppr4mhvb1c6TSB+dBlAOnC4us3lQr8+w0H7A
/KZ/1NWEOR6tRqoKfpz9uyTUulpA/odF7vMEaxPM+HWV8YGNk5DzZW4FxDn6fjFE
J0/3LOz6Z4nHN0+pXtxs2Swd/5ZhmWOa1W1FiahuuqZAv7pdnl71I79MvACAV7L/
BuDieiO4jquCgbxYOgnH7TjAdoVf28/Vrv87KzTK9yK1wfn+mMp8G8znZ5SENuHc
TcxXm57lkmCqNYczSuCv791pa3eFkU8bjRzbpzmDA5ISz9m5EuGLLfJm8N4G318U
sVHw9twPod4qzoVHevW484pU6KoQI0cAAsL7hwyfmOEeBQ++4AovTNRCvYrxOQvO
DaqvaYoOxjdcRopAbGF72btUaZIn3983wH39FRweufq1MZZLiNlvl6+kNfNH60aS
PkjxqGhZ+oeUJnmO3aBfEP4G7aA9aNSeMg/5tDO0ZV12v1ROVKcqeLOnSwjeRMM7
w3T/6Twu0HY7zW4ZdpfbvRT6zifzHy/12UcIRotscMDjO3FlEZRFA6wod4mcWmeJ
A/IBL0qAheSKKkgTm0BtaQEe2waHcNI7vpp86BTfAifk6QUucCCgqcsGc6EvgY2i
7g3O3VuDJDZcFE+bYPG2chYdXCMYDvTgzz/BZWDlvTiPPAbbhT/x77Zz0HBk4Svw
JPBX8wqt1EwM4XHLa2/h3lMu3ALtEwcRRyKtIfs1sgrS+jWcKY+PCYXX0sfX17qk
MLbxGM5qR9nBjjcs0jDKfS7E/1AXncuQw2Lhf4TtibdBKyR0Dnbd7c4iBtEPSuDZ
1zl3nKhp9MwN+urtJnrk6Z4Cjs+Dwuiv6Bju2lxWm0HV0XMnmOANveU+UmbpMsPP
vMj1n2e3UiORVlhI8GwY/MU028JkD4NTGnlKRA5rKWzSu+ADQtV18zpMWx9+2c4Z
acI1WARtVFzUx9ViwqAXMNwCwwtGF349O0G/Ag3COtcMUGPZNXWweCxuH2+GUSzx
xuGE1g45TkHPQVuJoDj542CXflPkeXaoqDoLSrslZS8iznlFOjke5S69G6zINSo1
py3TwfitXVv2kTSVMIu2CA1EDAg5FVlnMaMb08HSnb2m2MdAyG+l5f7iOdOOoAB4
6GNPbrOuFRyt1EjsyEfL3yOkFV58Bz5aKR4pa3nQ0oZM9V4oDYaKu9dAgDE0WtAV
ty2X4gIfEKPCdPfBL7cL7U6HMYn3QQ6ktZPcxE+xn1F7yF1wP0GAP1rw8SUkuww/
/g+A2TfeKCE41BGmOx+5f8LVKVCkxvV1ppYfP6EicK/sUsu4PbD2kGh+oNzzSuIr
s65xw6l/VsL7GebBRBIx/Mh3CIThPmtpByrS5UDns0VmJXnouGdsY7ASoZqM3epG
fRIllW5KkjTurj+BNtM1wXVR+n+UqzNnjux7oUZMIriwDcMvtj2lrl+zgOL5V5h7
vzQFnxrja3M7GX7/NGoABxq3ayal8+xSnGIsxQtAuUektFN5VaH0S+eS6NUpulxB
shwqbZmFrreXdPIt5ISVYE9xAXxEy+eERlfglFD6r6dF7z2vaKC6K+WKeUGOI4re
YSFfQgucLeI6mamrb0SA5gAcmdUKsGSBTLpaWuTlLPQumLsvQfiMFt1MCOUtspaN
0C5RLsVOkg0v1eHwwyCZGjBw7SzfkJ6UlBtVw53yOjKHJe/4Gc1+nzpjOM50/nW5
f5LR0e+I0sB6WpEIcZrie8qsC725L6Cn6bT7GQKUCufuQABo2bsbe0aqR8Q+A/Xw
VQEeDD/NXU/fdHBnm48bljEMaIV2dVqM/VXyHdAc9Rkbh1BtEOplBs9k1xjDBgK9
exynZHJE8LBqXF2mBOy3T8iAXSVsevbSrVVkSNtWR9oiJozUmIeUKVJSuShthwG6
ge2LYzEBjOZ803NJHH63DxwQRdnY2p7+Imgs3NHXPGFnd1/GE9A9u43LKYwAv64X
7zbzC04YJMquwCwS0Zfrk92V25+zg1F3+cjamAy9NEvG+p6tgJ+9ZFbFwlGhNMhU
1vbE8oWouIkba3/gtoJns6SPRuvRsH9swBi58xJ9+dZos6Ex2dQ8NsEVTUHetH3o
10V5cXr49LtoQ3mAfWpOfIbAOmM9n4gVAQzw8OXb9C0SgMI3b418CEYWIhJniw+U
z5Mp5IC+O9MiPpKxCDg/+lONTNgChFukI6mZD6hY+Ah6JRDJDqe8pnmhC2dupQqN
VUM1d5aFdaK2bGhmk0DhduQubmijeOiy02/gL8J0UJShTdyy3QUrJECUKDYwTzdF
skieyi5iFPqtOOOlQm0ZZPP2fG47LJ/WQWZNJ9kobc/QM/TWsYZTaYhN6q6F3Sxi
KorfkN22gqZaiYuT7EKyY4Yohg/Qr4Mot5bSaF0VqdDpgCXWTBoyLCb4du8NjiTA
sKqBgC+DOSNENuzyVy6BVkT+HKwMJJnnPwR1FedgL+5ob6YlApTGLTzrrfFskdQT
QVNwYeYvTzAwUEj5rE65mDhzjQUfPJZYbenN9BIOFCPgPKECp/nlyiVKoGtAbeU7
UTdu8BkTHx4SSccLqCM7T71+4z8APZvfPNQcDatuK6K+9KimSGpXh4eY/IMjNQ5Q
o5UttkqTnDvsuC6AEd9cW2V8Fvj4M92T3/p0FEc5JNmHgPzqdhV4d7aF7NDUjYn/
00ZAVdRrKh7Ml6tThp/cFdFqY5Hw1tUZwxzzLS0HEVv9/tsK8hIMlJEKK9/IByuH
h5CL15ZrtJM4EURavVbfGMdI25ZJ7nd44YwZZu6r9S/ewmcenlCJH6A3mvKqUBsG
+JJFfPv3Iqz8bwWkIC8kpr/MGOqZxkqfr4V5M38r4VxRuEl50PdBcI7d1ZUDJpZT
EiS7Nh7HfqzEBe/uZ22NrkRBLiK45trT+UKcIXsM1kr1pSNYFZB3nvVz8JcST+JA
rTarKQTcJpi1ymCRmssvC/0faK3ziW155GtV/qMN9LrvQeZu88+bDQ4tkNgi0fQg
GG40Ilv36qMyEBvelUr4JZvHRRknwCsLY0j3qq+tej3c25TfyztrIIdNsnjCE0fw
8mJztVyrkJKTmEKhGD9pB/14Daz8lxwZfpsVPN62/NecP4NCnwn4VXPHA1nXHaMJ
sZ97wv90lAX74rlF76fmL5sUDssVMs/DzoszBJRXD0+3EOevhK1KRfbrsCqLctOp
J9kLRiSbZS7Bw9SdGEYlzzyUENpjQK2fd7P/Hsl2v0vxMgp9Rjzq+2vd77jAhpF/
I/dtg8vhR1Q3O5edKZv6tGogbrSmJxRNHkvQmXrfu90/vnkPA+TOuhP3S29zHSND
wdYPQBKJbYxPIEFUfQ3Nua7IGRpytaJ0tSS2M5YGBabThF2kOontbq0uS1q7DqNo
VWOolzEe/P7JF/yQWnkoNB8kirtKyd2IUGFp5C31Nu6maQytcRZTcl0ELmnJIIAd
n9rfYL2lnsWbGEeN9i7OMkRKhUbaThTMPSZPZuQIj61Mu9UQcHTfgitXsUoheEDU
8aYVYlfFJmhCCs6O5fjDcqwLJm42v+riykoLr7UCI+frgK25T5UCn8yZ6DmIKjl5
wXwTaGOUkBVB/81t9IXp+elu4/tDMH+edWpky0xD5El6RUG9jD1eJf1Djnq+Uujw
YWniM77vxYA4TlBJWaXgaYVBxNlxf0qLy5SFIuojJgHUsSneuhOugIrEx5nzSuq6
wc9QKdxzPy62L1qSEL289VnuqGWTFABQqPBjTy74GeyLAVKK2AFnHmczxKVPGpmQ
UdLzCZs1b8/R7Rdkb5Aw9HISOQFnT1/SPdDBFogMTkjHwY6fEI0wDQfpB2DVjann
3mA3py6rH8smeM3fWlHUFFY8geZFBbkneCjVmYRIhPvipqI9gJ8ml8YiPIdwvQVt
DMcioTNCSqm9/O8e3ypIEaQ43+PnDvMf26twiLNpsTL2Aomc/EXoCzL5LIO3Kcg0
gDQQLR3sw5SY/ErAJhqqqtd+SjH3183IvE5vRKAx8+hF6Z740YnZ1lT7zwgH8vTu
lsuT1OES15ZUg2kTRhylWh1KdrlpW6dza5BkGOfCje1U+jtVvpSMJN3va9pjYyRA
M6VJyK+W94Y2OaRm1Q2jCYUVUKtThw5JV273uTbMYbFZRefamwU2aaahZHGrxcXD
ite/GnAxJgHF2TeGYqKF0O9Q4gN24f4iwciXu4ElNVpor+dA065sfvm7xXnszCu/
zMeWHUUx9XuuROYcrrvmKpzWuTKEN5dTPtngpc3YkUfF/BN8mtxR0FR8PysoW3x6
Au5T+y76HUToUeTwi0yivbaZpqirWlBoMikoY2E99GCCUBaW6sY+K70MrkTSebpG
XqPZtWL1Mk3C8k2UGifL5YZ//NvVFVhdcYHwEPanAD84+pIn3Yf6KmujVF+B6u21
Tx4f4PGs6dwkJig6o6GPzFcAO/TvVj36rXbfj5PqUgign5tqscWCwkEUs0MArLjH
JmWvc5b7PYitZdr6QOIwIMuxxusCo2ucyOtkmyiHzF9UrmQBLsoiudRLkYdZEmf5
XMvRqV1JcSdoDYQJjM6K9lXm3bU1dink15kgqH5/9Vm2/WI9Q4e5xwfdTJNZATWG
ADF5EXRYPiAvm9Y3iJJmn6f/9gCjrzI2Jc/rCY4+dDecgW2adaY0egQX/+6wpVWw
RjUcnMUuGBXcvPGWNzgHP4n7NyH27BybkRN2WEurO4UjTN0Z0rNrin7bdDdXsk6+
mn5LWn0RyovtC9rIen+GHuPRlOl5PjAtKzipHqXLgskVtgAAwSzcmGhvCmgfgMFm
GmgF8X/saBrx1r6cXlDZBIXAzaKjVxPe09Sbz3GmTQtC7hEqdPpf7ghO6W4k+6nR
bjUhL/1kG1trlv3WJXVmgv5bwDucSMUU1pVe579DRvTjGDnwijqIeDHncscL/hsZ
NLL8HEz8NRX8F5T76Sl9O7Xo+/Ikploxqpr09f1MBikkeYCjqsYlPI79szTjPtoJ
eRAeLBg51iGJTX6OzRY0X0AzG1I+iN8/1LvyJwY+Szq9PujD61lvZOg4IHLjVCoK
6QohFHTsmjNSJWSqTy1GaVNwyNYTdl3bsKSEPT2WjGpnIPmlPcVRpNMv2CL07ysa
EqFqsicuGM/zxEtr12rKZnEn7sBMZESk76vFQ+pPdX92F/EQ9CmN86IyIh5Msz30
gIJ/zk6OSro2kiTH3mJu5+c1MiyT5OFTb2XSwqzHB/zKqIoqnpBfW9fLSdohXZKu
Q9Z7874VzXQWRF2sVob4yYNab3ueWFJ5O+0Z/67Kcz2PE4dJeml33TmyUoZoNy/W
OlMUxAoBIlEfJhLvFmjfB1KcVVct6lCuMZK0Diep70P6iekikun+IOGC0jfczMbD
NQ8KWwSa3TpThX2TOjyJYeQ6C7Q6nQTUVFv6taXeB9eXjbpN3KkUsjztaDZuSOZF
1MoN5u6wV1OX6mEoxR6S99iOgLkbDa+ouqRLLgUAzBkVU/uAI76m5OeDyq4WUCTy
uXYIiqpFFOuBoVtm8wFoXAT5oL5ej3i4IiF1UGuBkk7aeJ2RrqXKf6hJ0KnhvKmR
+RwAcbw28M+ogk++amPpX9gsIMSF1tcOjH6hdnwO3WnVaMZXrC2wumcrj96dpZ/C
KrqnN2DAQxuyduhKEaz0g+5nuzGONX4dFxGgFQvILI5sgrY04NQC5cENcSigmJRZ
4kpictkDmxDFfSvNjpANTH2fkTDCIe7ehwMZRGH5IvRJogQ8oKBnXGRjWbC+LSXw
R/s1sDx3AXEN1wKbg1ifggq2WcYH8SNrNJKkodaLW1Wfc/XRArma88TmtDid/Z5X
qRhN6W4J8X6Zncsnp1akwwImC9thhCUlxziDVbJFgRdIYDfjOn7SzfHf5MYLHwx6
RXMnrfi3inV+XTmcLbFbFWJXAVqI1BRyWMN/aqhu68EyzcF768x+IOSq8xCPw1bV
VAaPb2Ay/mmsTsmPG8+gWvN/I36bmUZAjlPMakqhkrPhWORO0rxs2KPPJQJSDn1V
qerHriv9DKFip4tI1oqy8RYcvGuGCnuSzSb1WO5KgBYIbuk8btbe9l5HcJVveMNZ
TdrjjR1bOxF6aSGAUWlXWW1Gm8auKIwpilNL9GTv4CeslUP4EhHUorUQMeryoIa5
gtlO2W9PSsG6vR2twPHAFlVl5o3ypodgQYsmu4I/kRlig/NsO6Y1CyW50xKdqqcL
7tq4snTHJzJ5g5hr0Iiqo4EosTls2LcCMSqSjsLF7OrsWslDNbJLJ+G75SSB8qsm
iPd4yAHsxNhqkkb5KSwODkMZpUuzvgnUAxq+rwDYgMf4eb4dXai9sfPaPEIT2fY0
eBnb7sGlJK+rWkli2+0JcM8fVPjntWsEfelKGsjd+XeyLKIKPsFDrQPFsRMpz+7e
MS7pO2TE6FdPmdZJCi8XhWToquIZLp1Jv1mT33GLM+BEZi6hgj+IeKs/Re3qC14b
hpHhfR0Est52H5pMok97Otg9ea4c8etXUSZJEaVWQYrn++R6dJtwof0h5dspGX33
aFnKpBOZZkUhEJXRwVXxemYtIl1ICXPozRGP6ESMoyEkgtLitJPVGQJuw8k1hZhr
qJRG2s8LHooWI6Dts9A7++N5LnQySR5M3AZKFbPvWhNqJLsMH4SbsGYEyhXg1WaL
3n38NaCslPMMhIO8w4grKVpW1uy6V3pGjTr403hHpXD1z3TG9Nc+rwiRvKG9mOFL
bTtLrGFRcO7d6Xnyb4hNP7GPmLHzgEwAsY2WL07sfLPTEKTOopVeUF4s/TxZLtcc
4dtwQJWPtVT6KqweDaeHrUN26TxEuvuGEcgb9YMYz1ZKKJ9xMYdzZXxwn8u7++bP
VfWFOHbXIC16iw0v61ZmcmWXjWYxGkKbM85BcN1hOJt5o95G7Aj//mf2OW34QYGa
NzIRDV4KmNAM7vtEBVb8LfKqvQh8nh9cWvnipmUkYVJMz059+SpwTHjiVjt1FXv4
0hgz4DfgOGdOMYt6CE7V2X7zo+4K6XxS7FUbZJe1YO39snHekG4oPJEhwBDTAGqd
VjQ3htj2pUapPL5YGyfoXd4GzAGaHUWf4ei38x8P5Uq4g/rPt0EWyN3QHwY8lHbJ
9K8+drG+vjG/WZybUnbDdArgt4FIBRuUnrMy91JIUtO7pBoBwamYrSBET0awq8ZF
Mhha+wCWFKJpfa+7QC6GyBSuTDfDItrdyIQ92lyUBuqGKblFGW6wxJQWjHdTMmIM
6PedhkSD692AJuPOJMtkobAnxiRoNXFPxcO5xZCA41RacZTxrW497cbSMjQiaU3g
VjhERW6A2K7iJledpzuet5qlhBj6KjrPOUFvXQhVsb3skc2BhNcSRbZQUqfGQzvS
RJsaC6RmjXVOF91RQ2/x1QkyWMwQBTWiLIS2Av9+Fv/GMXYCFTZsoOFfxDgc01gT
vL6WV0bSu+vQq2JUdRL30+H5EsB/G+PaxMmLYGRp7/0wN9+7YQ8YDoGn/cAFYCbn
KtjKr6pBT+1c6UT4giULMf4tW05XACzFnMHnYKoRXIMNJ41mbxgtnkBUJUmj3Y0f
CGSq0epTQQMkUeLaN48KOQShodLKG5HpwyOIDA1hlbi25Nw4xSo+QxmjH5JPP5bs
3TEmqwokHLf+iLx3E79BrVStVnL90QSLYnEyXpaHYhB9hnOw4Wz4bQvbTbtHBrv4
EF4Z94Y+6YjHLWai2eh1GWos+fVaajPh5NgPTL6kbpXQdGSYk1RKK8xCAxMuodP7
HGi/szDjzwPbP+Ln4BaBDR/ryd4cx9lWj4ZMQL0EM8IRE7ncehiL7x5XDfwS/fFh
WPNnO1iKKG5BsvNh3ZNMfXQZyexiVczDa3qsSDPHpZHdDLlVG6YKEOSpTghUtT6N
GlO0K3p5qYb4/SPpW5slHQS8m+0sUYcgsXZWUNigAFyUAM2RC4Acj1sbSesGFqwV
e9BJg6uwCQUxZEAcd3wTJG+OTspl6M1qRqHLtOuhAazeOH9xR9fyMs9AhhzURmwI
j/CRqiHuoQN5rPVHfC/YqcTdxcc41yZZ2U7Xwo8LNW6aMQpOYsrUxy/9V9S+7HM0
p3gEBWtIxgmJ9cR3LrPV8ltKxnXf/Hp+SJR+NvEAYD+v4JV2KCySrB7laiHd/Lg0
LZCbHF7iqAm9d1iSUL0pATKoTfh7NqQW9vFy+FtEeQSvh5mNvZhdf3a+5seGRCli
gJvb6oOsj/Nh69XkfIckeZx1lmPp9DqYe7FRDCzjXI0FTNw86cTh6gRQtIQvl1F4
8cIH+cWTrVp8r6TyXTuWdMae3JMQicPJph/RLgSJ5JQ48x2vd/nK0BRJ5dXZ/OLd
GsZFP9MQV4y92Q3Rak+qAsJamBBCVU42nWu72RB/+rmNSxKoK4JHh18RaIdAHSQt
zVpwB1mYNMmKy8GrHaNeZcG6Mch0bJQkBcDLotODTxtKKY8lR+XjnqSpvOCFfw7i
Dbs6/f4u/dcNYBoccsPYMgnsY+aiqKDWl2ctfWYhfLRWhlkR7YLupPRWLwD8ayLk
ir7y9QDbDOQyNhcuBTEFjRGbtueKf2ScgzonYeYLO1LLWn7SdTrO1WFLxF11xGpR
1C3HPAH04E1jcJ1R8n7+kz9ikReDF7ElKXRMGXl+5F6a796LVKMaLJeYU4sSQT4f
OCLxPjJ/MyUF93+PzWWOSoWkDsIFoDosrpYV9xidG15f2CEpmSr+MaWhyFrEbLbc
RXZdI7wZInkqMr5H3sYf1zlbMTufYxQJLKGR+6FBQVhUyQhQM+Fxjtgk4XSEA9FG
tabHvXbywQF/AcJ2djkE9bfavK5KQJHse9EHSVkRV98j5OEFHxTJ/KPcHuvhWEcN
ajn/mwIReHEcZq+eUADFEPUd+aU60umQjKdsUb1gZQ47NhgsPPgpad0WnfBT+Ue4
VA3/RNjGPS7QqPFL/VQPZCbPlZZXjCI3F+KhJMYrm9fr+f3KK+1rEJO1MwD5ydNU
NwRyOBP8PeVE8ZF0u9gXiP6+hRDfPNzjqFXD0gpJxXogYR4/ySEtQdy9nV7/htGM
NYjbPCksXUAnVZVDVEJMPltq2uPgmdqMexDQA7W/PtGK6QuKf4JB0+M/5qy5jR/+
X5pRJtj7tI58r246jlfyWpC12QMe5O4357y2YI4h7LuTOmH0h8VIYFxirWXv55w0
Dr9hhq/jLSOG8F31X+kEXjELO7fAZYMCw8AjiGVg0MfguZ/q1//YwevUNiAmS9Gb
EwUA0qmNRvhFhrX4M0LuGPNUIuxeuiXxmAhibPCDZVuEDYZVhQzrCq8TFtkETRhZ
3a4KGyAvzSiKRordhtu8ocrZRT0DCgGdxfqCqAEo4dUA1SAsXYyzTmEzwWRBlPqH
98UCUWPSvuzf28lpLt5Tp5EQXKuw6+5qtBT2im3AWao4Oapn1BAPQHlrIkcK7Hc4
PwCBOPE/BHnZO3SA7FHw99Ue+l23fjNeN4wmayqJtinbJYRWZ5kEmurW4NxbjSM6
nZcRVe8qHZ85yKjqgnotYy92vurTTh2up0T1G8mOVaI43L09yvmk0jLcbz8x6W5z
WoSEzPAEM78nd9K7A+f0pHwyY6QMuJG8wyUPPDomG3uyJFEmSow7jdCQPLhlS5RH
a/6Mm2QKKpyGhHYhTxCDdWv0FS9KWUNzD31T65VUO5oOHXJev+trqWM6hOQVBAWL
KulSrbYqm1Vr06RcEVGAtwZmj84oFx9YV20rswWUv/nmMzpMfr1EgZOk5KwrwCL5
ebe5vx8HyjQb0oHBdrzfEsVPYUEfAKWCPQg/rPvfBJ8JOdx9DZxIk6xnLrevhXd/
7J8vvD/AkrW9FYr62jWZm66Sw38fqKLs3EOPlFu2qnrXig0AK7e/R4kh/mj7dZvG
9m4pXEBYAAf27LDdjzKbK6pgt7QKYK/VVZVRDGzanP70GR4v6UQVqmWAsCdRJ9rm
PKA8o9FKVyo5Xt8bK9WLYwTHmq84bmI/60D4FHZbG5fP9RyRC0gBkDCuO8ThQhqA
e0W8o3MDPW79ymvOLNYkFIT8etBAzhwkE3+ukUBqCZa8O7q36hiXJtVeXQJqoZPg
GY6abshuubUwKYl5VH3/ScIu3HrutNUOP0UY6TRme5NDEbwqz69ACUvQe9d2t+zO
kNyR9sL6xKgiZy3L3zQcMoSfznu7jGG9+7af7W+JOhHR7zt/yhA9cBr54oA9qfyw
P+3xZ7bPuH7+1S2+H7cRIX4x9n5oXjM+i3oSe/fVg/7zKblVslqtSsXxxCZ5XY06
y8hOU2Y0p7LxZ8zBKiGBjoC8Lht6PTWurz76k+1tlUNKx5nJU9f0/Tjx/I22b/R8
s7SfdaO0GTEsY5F5+quXTg0cI6W4f2bmyxPU8HbIYn864u2/BvA2Oey2QZWv6GcP
EwmGAzopHKxTzb4cnu7dReGplawh2bS7yYAib9rbDlBjzL5NxdQ7GL368SGfN8Hb
DPraFVXbDUnIqJp4PYzZVIqYZDqNQJbXdf0vCAMo1YohZ5q+r3bLxXRCRat9dy/U
wlur6fjLsZIsMDAZKy3UC/istw3YUN46GDPm3XTyEc45GWS8hgaVLujzgKcXXz2k
fa9Ek+zTRnydGQnzVQdxrWCImWhi1aTwE7L4Pm5seACSiQhaOW/7/9cVCVJwcHyA
n07uttP1KMROrVm+L75YfDlVg98jQ3IimbGpu7uiLItx+LkHPt8wf+Ib9ruSH2aG
1+Lmo/Bc37MIaNBSXAMMsNjg6pFHQnc6rCH5cTLCZRNtqzjremP5CTjK8R0Fhi7g
5ywPr0V43D34fXtdeLCkk7knLYxzg8aQ46C7RHkcb6bF/GJIb5jS7wbeDXF+BBPe
3GSrUmNkMpbPPdw314xaBxq7kEBKVY5CnfpVWyE2NlOKQLa/Wn1zOZTXGjTYin9x
PDdb5JPIwnDMvXyE0f+rzSo4y/oVI+g6GseVeG2OzmLMTA0G+DMau1b/g3KdFGmY
2GDL+Y3a+RrfeWo1oqJpptTC32RK/omyWuVsyeoYMDx+I8YX0uZg3NKm9arFG2vs
NxCb2YveV1tKtk8JeKorIqzUGcfy2ljb4ggwN77siZzGgXsmF0jIdJbLpbdAZqOh
Pp02+20p9j5zFSac5JwchIcNueNOb1+bGQhw+n2MAa19Tr1FIxLsdHqn4tSlEQV0
IZ5ER+eI3Etr/rgAPQhHhrzOKlmZDSr4mDoNyY3OlJQ+x/SC522tRXYPT2uqY/HW
1+zmqT6x+dtHSXjnfuVKJM+VRvSuERAv6Tt+IJ6detQz2pdS3KiC9nUgIGcwCSKL
5Twr97xKKv6cMeY92Hz9ijyLBcNKBmQiaf8FJnlRVSlgL/5RfCatCa94YP+GXOgT
GOh2vMK1vbDlZZoa/qejW6cYGliI0brHVUSR8ZGo5umS2wcgTY8MAMnGtfAkm3WS
pBFeS3S5A/YlcWqvWKWj7uA4HzMHgzbeOaYo0iktDKKGjVRMcyQz3WliVSbB5x60
o9+S4YlTlHY5IN+8/k6oh+UZUwhxpGz3/PxU/OpNglR+9PE22p1I6C5qJKn5fr+h
eCp0y2ld0jtE1xby+M+esdzowzXlO73OxOafUZGD7ZdoibywdxRsZyk9mWpuuy6i
5v2m18G0klq8hln5P8BS+iKdv2JULUOVvB8klaOTpzhgDXZn18DSDVCfttDEzhzd
I2j+ieqXo3rEN32UtZAoLOzZmxAi0Kr6oKNTYm84EEcvPqQzY1hNtSJLrVAr5oLt
wcPDVEyMByv9HJydYNS/cvxTbyRvoLEvMfMt544PLTgGFrP0Nm9kdv2naAO3GRK1
iqhJ+aJlB5guyx94vx2FCgH76SptYpVZk4rfIitneUF/wK1wxcWz6EzW+Bx7HlAk
TTGP1CIfhD4ixNX2LAJolstolwmhItiTDMExiahuAXcnxkBhRbU84gOrvXWj1wzJ
PxNFGYzmDxsWQzx8c/QiJOfhlK5yV12OCpmaTd/OmNyGQwsxRF+TFmVT4a/z1Hhi
LNRHHrk6UwZ66yBkrb1oRarPtlyykVCLVlHYYZaLiYCgPH9HBgFs5uGH5CnlhfhB
SbYFP38rY/3p47VAIf1e+ChHgPhTQBruiEH8t+RDGHoCML3IWpX8x7MJW8Myio+c
0Hb2uk2cxWqD/2AFpRnMtBQ5NQ7x2P22gVnbiH0/umdJgpVLp7+eH7/oeXPb6bjw
W8KR9l10C+AdFuGDoRMXPiadERYLrkL3mw/pWi+97CIbxMH4n/ZQtzcPvuEAFa9m
zOUY8ZTkQEuoHPpgLNbkgp2NL0O8k9GiPiMmMWhPiYVVpT7zkhbLvvhvaS7pUews
Qg5pZ5kW/3GVLI1zByPd+Ixl3Gpjhj2um8lA4bZUrNAP2jvGNXS1wbqp6zvLC6X/
gLZOqqSxmdkXZ6nsVS4nMkxhDI8EdGXXf5uBvbe99jbZplsGwD0h36uTOao+nqtL
C3nyK/zHac9KdBEbIarD6ZYMyFgXBG9fYliLndJhva8xDxQz5NCpFqRZiSyfxqvP
1YWiD0ehzcG9Lp3oLmisCDn7y5a2TVuNA0P67JIvCz6fP91Akz/0to0iF66UXlIW
jxhkq6e2kdPqbW8D6Hue6ORcOmwJ8R0FRrW6fEa6Tc3Smxytx1N/g7OtVn43WClr
g5b7vFkXs/LeKzv/60C8g+PxQyHWX7ezPrc9t5qyGZdJuDCDZS58/44DTudEjkBH
GDuzvKwgammyQLd5gbLSbn4xueR9gMudtlZFsk7tEqL1YZn/gXSBTHUU4ai2X+0m
DQWOwlFap9bmefgZcLAxvCXwAnaPPe2YOufuQ7goy1td72RFvo7FiJF9m1qQb9y6
ywsod24rknqoihsKNX4tJQZHWQDtz/gZDN2yG3Ig0DGQgYg89JHwsdlrHYvPvIDh
SZUOJZV1GSbWnPXLttQtpa6pMg+gWz0t4ottC2kTipYnnxQG/HdLR3Y3uupAmzy3
rgpfFQap4ftGFFHRvVj64HXIamfpB+9u+eeDUQFKeLmvt+gNGLMshV1EneCntS94
idLvX602zq/cwT6FmjZJqZM1HjXpeB4VXV/nbuFa05Nc3FyHYcO0jrrFqtIzswyn
1rTaCzvkL3nBPKyoU+PQaF0RI9dFdM7qETZBaJtcofjVgohjbDvswqvt1SVc7fJ1
CbntGi7mGQGmFzFfLrMO4GaErmPFsKj6yp9HphIQjomaCF/7Up0TwI5PsaHCgSFT
dGdX40Gct9JBqDESUUzmehJMHqSns1ZHnBPOhlj4QS23oOKrxbxc0dDDVCc1YHIj
51eWshzyblmKTtpeTbewqKkwYfd9PIUkTG3T8YdPlZHoEz1eKr1lgOmVAz6kUlbF
Mnlnw4SodcHyxcnv0R0uBWJIJ1aVaxJn5BbdbWCm8Q58IhXESFsKTp/zvqp9/1fS
QinH+FgRYRZK/zkTVMmHGhvK4VFUyNHPGCQnnrELF5R6EmiOsjvRwylsMdawgP4W
SHJf5XBRbsnHnafBxCAqBWJa1cEWhJsiRw5qrxpq/g9xyfRZwFHFmVBZwzLG71aF
HxNAbL2A6X/kVuyyPWPGmbuKDY8HGdH2vN+BeWDi91S2kC/NwLsD7Qi5t7j/hqqb
JXkW9aP4NLda7R5rxlRQa9LAimEHJhfdgew1WD9ZieDFdk8aXtqz/ISj1qeYFXjM
wlpakVNVc2V7LxQfUM2TtYz8LB9lbs5E+0rubqscVSKnubLJLxsm0zZpcTJw868p
P3c3RGCBZ7DrlqTzn2HvUI0osDkYKsVaF0DFqklieAzs9vOZyLQZ+u7NW4ADngtE
6HRAA40Btr5W14SyuD1JkjcBNfONjPb8RSrzvoqABBYiV+uLIQqZq+EjYLL16mGQ
mRNumsicxswgFoYcSqedUfBmUW5MU+GEFBm5Bu0hKXMZ0jHAprHbp87ErzGVcVB4
//TNOz09DXweIDnv5EAj81XmNoPZWVdy6X1AS0KBI41ApmIxAzHuTlL9OkIFeuLp
mtl4jDKdTPzLDHQ7fiAJ6DYIG9CbVwwzeuy6elvE51rpLTcg9zfrr0eboiweu3bC
4sN76HNe0TiA2GGm3lhGIpagDCsLi8dkW4X5W1BGVi1THhyKwDH/VT/A/qG+GP3v
/fJdNaVYuls53ha/tqPKUVAwIKHE/9O22j64a3XEaSCt28EhIiPtCG+nncaEw8Am
SwyVzzIRj8IzvSBk/dsCKS8iFeSQD9Zy7YUrpVLdODk8j1qp4bdtJslAWJzh0I9Q
1jKnpuFwDUXxfRGgmxvWQxLiOiFpextI/y5UiE1DcK3XSxFPeP5OaMPBT2yi1Evo
MFAzj7dicVCLBBKBhSbsgOhTuddBeMkKdeUxN2gI8CqfvC00TNUR3yDosM+DxhXh
PeGXU6wfYRJxPPUWphvTYkc1dtdei98uimLwNQgqGWyywIN98NN7H1zghJteOX2p
gpRC4z50BtCGxcpPLMj0kT1Itx0jvbWXDYbYKPEJIYXzU9hRyODk/vGqMqXsCu9/
DCTmE+JcP3BgtdOf5Y9u6JrbQ9mULukt3uub0Z/y1FTdT9aSOLDn7tz54Kkhc3MD
1NewHMY5y7rDB2kztv2gP0ylnD7zBJ4iZ0nWGL1Ni713mHg2yjUYtiMUmZ83fbBO
XIJga+XjXEQ1pF/C3xeHxf92a7p/c7hOt4FTMSZIQecylGhQBcs035SLdite/TP0
9iYiwXAEZOwVrqpHsLmF6bYYhVL6Wh6AYPRuk/MMzGEndvfneQjjFCqro+JOzxyG
pfyTMJK/X7JbYU5V8NMAITsscWxSt/kHItJfUlNnbTC1lE8pI7ZqVL6dCjJShuAc
6yB9ybGcZ8hCnqxU2Qgdc7euLg8cznT38+TqOW/7NYLMw5ZyXUOApgWBZqpRiV3C
W2tokX1W0uUv/P0ZnUbeVPp2VfD6TOazcY6ICC+RaIOvld1qlW7k7Muj3ojT8MQv
dOU/ajxlPCwBmtCsYu+j/SwtfwFUS7kkU5vhDsA35HJYg/vmdpiBa3kDHaiJz555
I/Qaz6G5FXKvw1o59dV2DwNaGoudCsU/Vp97Yo6Ij8+9o322ORLccw8ROJz435Rn
IhtId4WBYLc4ASl4g3tK4e+cKklOqeDRU8fnvyZQSL7YX1eWnT8/23MA+kRPrp6j
LT7et3jGNsEfLmlylammVHSELyLsQK3GVmyXnfIntT3mQEuikcmCaTtwCUbWwSu8
IC7mwSQVOvk8U82IfF3jDW9TVVeByvBc69GtMUMaQ8UM5VVLWL3CjFfrnZw6KkMS
FnACOk5Ux4A+vHe9J4bS4r4gfHiKKG4AWrY3P6ZYT7y+KCzq2y2W+Rs97LxC2vY2
AVcPI08jIU/iaf/Ozc4eD5hlgRUBPIDEwD2DDuNnU8Q+mSPAy6MQxkydljzMVhgY
cqqvdTpHeAvI0gA2AifO/k370hVlMnOlweTa+n1XXnoJyeRXQN4msaNOGxUI18VN
/gWzq4bywHu+5KJeFdOMCQ6vVzUyWlYaTuzk8gpRBqjXlqwVLP9lNIzXE2fMaRmI
4D7HBy7ZtgMtquze2o4dA2lLSfzQCBWVFWlJ7nTuFZWrfUoWm5iENJRmv9Y5KyzD
HHih981ui/49RzQbFHmG8rNUytz+SNADkaNruKE5S0DdPi2N3N4wFX1oyBggxYiG
J+no7YSbxGa4932cbRzWuQHszaJCJfkXqXog142zuKigYmsX6H6pyuPidrYQZ2Gf
2r0sg7Rug7jX/Yyag4592Cp4KwLiNYinMgV9Rgp9aTU1j8l77nR+G9WwvWTYH7sv
4IYtPn2wjRCXED/R7O4DL3OpT7IT8AOcd2t36nUJ/N5vsSH9/Qo9X2RdV4y9hmQz
7xCOjuYAcVKipfDdMKyrpXnr3uZ8oYt4+HQpgKpWgPteVZVZx5YZd55InVl5bcPc
VUezRo1nYKweBgFgf/kLhwor7IkT19MrSQJxVJR4QDXKp7vEfEbLqwgYuuKA0gfJ
1ws5LkqMyP/aVpQqKcEGk0tAanti8xEHdphSyc/xhigv1GpqwNiuBfRFNxqbz12F
lA/XYrvRQ7Rn3Z1Q+uhuoFJctoWKjDd5b/W8SjGNRRq7Jxcrlc7Wg3UFgnP5CgCm
SuI0v9OrsCOewoHfid9FnADZlzHfpi0Uo2xUU3KsKeFgVFCoZ960xtnn/AjumnB6
WnpHnp4tBj9unmXR8wSSrcQP5YGsWzcpvKymu4DY+OLpOcVOre1XIzmdniPdpBnf
36G5Gk9+Lo3Dtx/zVlgq+eum3FIJbhwiENwN7/8UpkcvzzFzgKvVsLEt1J/82hjO
waa2NNbtbUdjFWFnwM/2V64NfUtw26Yts5q8jksipaaYdS76Qb8cUyGtJwPX6KTo
Sq6SByI5iPlr0ur2th286BfWbQrU+cDtbV5tWzRNCW6lQQBMr5wgsitDPbTAl2WL
YtdhK9dMWmpdtXFcu/PjyOULBfw/giiopkPTx4piYVni7hSuwEbWy7ahwrPJym+j
J4WyvX0ZCvURq2a7hUjgnChC22L0IJe6Yz5w9sRN21uxaNJJkDhjnGCeL1H54vpQ
YDQc+l8gMRb6dCeIoABjPCnkF/eZ/ukjssbh4yAvs8UYhmKCLe3Ga9bd4zyTBQq8
frX0J0vg7e/YfGDvSIKEuddSpyjkgVAYVpNPHnlCJhv3P710FASfw1nHNpJWp5G8
pEgBcdPov2i1BZ4INe0yYAGdGE05ar46IKoHr5Me5BFu7TLD5sFKTzxUT1WtPplJ
9HJ/8b2hAWaYyXefxHspozTh8hFRTEZudPNZUTSl0U2uFsnOiL+vD2SMVlJ80Xaj
fCGHaoGUtocCU4uU4//ObAnbb4MzGLi2fQg29rFrRxgC3J90qsnn4mpujT3WRlPu
hlKuOK8Pm9siRdvFvcwc9dJh09BROyYiDalHD2eFu4wqlOqD/OUYVIJEJGPOvsGU
R4PY/x5I6U9WhKn86Y0WTvhSvIc3YKi4PD1LzwA1ZhQa6PZerrRqlIIAFHcVRtGo
lWemFni5ezxkqhfu3MPlgqM1DBNn3SeaM7u4Qh6CPasK8fAETrAxbwPF6P8y8KRh
2xAafwkvRX/b4s6SRFLq+kqFoItNlsvJdJLDOOJ/8a7dVkLXxcNNX5I++wwX0xEA
BBXsGW1WYE4Ai2e/HGu84Wq1Apl6x3CsTqTcvmtND04l7Oxlj8fc9IVv+5i4m26p
tmYM/TWRUXxYhSKPiGC2giLJyXmpAaBqm30vvUEOw+zOFA0PbmmTiK1yTK43zKgI
4YASAjFOXNrv8o2Lzs4EockSrK+4ZdnOf2zugGkFWwuUOJxL4B+iOruhrddP4LW4
BpGmkVfM0zPKf596MV/rFc32IbwF1dHP+RIW5gYIuCseC6ZNppKuonwZ/XVIJy0V
WTBXy/l1p2MkWNtzR8NHJ/p2I4UUEailSFQ6mQ4zNTPX+e2MkfBC/S35yF7e2z6l
1INqlOLZ1m6jg1MSj6ZZWj14VxioAikALSnfFXMQSHwwGkWYej23vq74UuJTMNYM
I9hOPBk+S4RESnBEaQ0qWKTsRtt0v0M8N3eJKE8TdLzPLt71CqDTZHVi14AMao0l
/Kk07szA2m90AEqB3/X+DpUbu0ue0obQ+zinKtv9mF5M6T6NbsrPtpI56kqzHIKQ
YuObb+EDFh7ruAkh0WfdjBf9T+Tixyn1qYJvpOkTrgeD/x1eXBoIX8H+3JRgBht1
79lKPPXVXaQapvNeW9Sbj9l/XVBHHR5+z0QtQPxrWbuwO4Z3vWBORSYNmSURD476
sjVqMzZMJQLO7ljm0kO0wBbivX4VlLKOH4jdvFK+647ZrdkkcmJg9k8CHkf92agP
fDPq6bhYSoCOfZUMZy9wc8+5Aeo0vqsIGJRv2OkhZa49BQP3Us6PxUx2cPzeaCO9
/fBs4uH00bCHKn9WXn5ifpMwTMvcaU020Vd7bkdzruhT5XgbPhIAvGU7MtSZoFpW
WAR//ePj3/sSYots7lczukOy02DvnIf4U4MH/pHljPmhkAoCqFSjIZXOZIoGQsQg
W90wy34xePoihx9Oq7V7eJpIb00mGBmhDQ1TciHL+NQwpxqUaVcrAiibfQie8kzN
VPhVbbJbF6qC0zvet4zGYzOJWKJxA1JYiLItoDZQgEEbrM6TrktWtC3JbCxWyonK
JtkQbY4/+OFArEw/GpRVn/Fnj8VVxYErrg3TbdCLhs78uHDz1erVq+uCgEXD5lqT
qaudkV99GMPdpkfgXjoyKE+9J/FdBlUfcV4u1XNc2GTo0qhVnaItKmsKStSiyG70
YpT0UqeFW7+q9CYH+O0SKHtCp16/eL6mPP8/xBk5u4u7VaccIKJtRXaR6eu3kXzm
4HM0D4SWRJujzKJ1Qisl6px97XhzHEtjzo8tKkg4KJRoHAZm5yV19Fa5XvS3zVpZ
o29DkBbihml8PT3NDPgaV04edcpuhfAKTS8ogU2Z4in724oGUpd/XOAV40bVNfJH
1kZbH5xeegu7vWsi/hEWoMD9i44HrbNac7Kp3N674qPioe37yp9987XqHVNFZl56
WCelj1xwGVY9wuYvKdml/9b869aWBZpM6zf5LsdkgDPNbClt3zoj7jQDTgfD32Hk
8vconZ25A2df5AtLAlXHhs/qjS/fAgoLFL5pE9loNh5Sh0eCeLx2sDvlSGETlZqS
B81o8J5/e92vedXsV/PSIbr+2sb9XjNPb5N4IgXKWs25TjkAEv/vDdr428o6HWyO
uU3LdNUYmY0UQ3Weps8zlZXCJS6UyqlqqogdF33hWujJE4AII3clRmJhIYfabY2k
va7nAN2IHD0X7nvTt1eIbNNqXQfVq3IAm9rzTslqBlSM4wE6b+QL615A5PBEZ6ZR
vwDReKmRWQ4Z1UhZ91cYkb27SwNQ1JeMWaZsWvnLl/enrgmIt1tnFfd25R9RmK/+
oLfLTjFdraAuKAzMCehO1e2YpJZXl+y94x208opUJmSmgkkMbtHlKJYl8HLLYy+C
zqt7dXI2+sgpCVd6r42n6dUYKpkXAzunJavw0DKjHGi51z+YihigLw2AdSwS9X4/
ld5f/76pmNnju2Xm/HteXxSyJx4l1vF04ohQ/iDToxIbyiDB7iUWYdrw+ishDjHT
yGxnz36mBmbnAMwAbOTJOfptw3hV4jRYMzHYSdf7hq/0lNmyzWt7YsMSEZrnKEOS
k+ZrPgkZjcqdpJTVkiGyMXnAGSqUjYfmI8tbs/ADXRbYIr84u8HioVfWNgk6B0+r
opKRVwfOSLNCtvkFEbQ2yOL8vobLoRC3paZ90STis+URepu11SNTevxqqigBVrvr
FnSu7n1tCsj030WL9N4xo/wIlr7/8IA5mTdjBB0eN8saOkSlRzrIwgagi5cOdmh1
HuMs4L7xrc0apbDG841rk+M4+nF3WtICyT7hy3T2jxSl5b1PKODvG0b1ZXhNS/kr
E9ifC1Rs008vm6QvvIN54lb6iL3IhZj++YsrS34qftM+oSUYE8/oetRbr9o9LlcJ
8V/yPpJTWQnHiDOWzz1ZDnGFh9IFin/9bx/kTUaIATprCz4DHbVNCipkSZsMaWiL
fLovXRWt7jhAcAL6B2Dw7zRWGo+ySGn+zTk971vIEGRpVQZgFJYUAygb1lhon50g
SqVbKc2kNkyrgSbvRrxM38jLzXE3AVZqOZEj4a3jmpRvlJeZpyYabwyjZoRje8Tz
nRTYXooR1MNZndPukUznTUZGeEiubrZbh4EfQ/xQ04SZNNYIJNtvyqkmvCc2vdYF
UT7CzliO7L10+NYxJLyjnVgTG95NRkKKTDhNcRNetdD6vOO6PbkOveGeev9jnYDs
GvlhQM43WM66lAaB2w3ywQ6Omb1OSMA9e7dAkktCX93fjNqXdAVLdKTyxvINEZor
SDx4XUS36rRuDl1Du5AV7vEAi23fChyeaXzTxNRV0cGOZrHkfeksXk5Cx8yuObd1
WwnYc26kxoYVn1YdThAVALk79+UbSubLpG3u4t7nRlWsTkN17x7Que3KCaIth09h
RSu1HpRcp6Q180dAgkbuBW4hvgPrN3lmox8NI8SvBEpueWnDyZQBXEXRhrnJd/M8
6c6OR184WqG0n1hBIzMWpiy2n0f3su+u2antzORLmWVrW77PZk5AdufXFBlWFEtk
CAJXCE4H+Ci7rqzPbF+DWcnD9pNDYHjFi4QqJz9+/XHWbbSVWnv/WIu/VQtwUzkA
/9H/JBBSZK8Ob+AyLcv3VC5D7UpbZGoBUVwrmWNMdIg1BxfMab+JqpDLGRFwQL09
UZkiqwsyvJLpBQWdgS9r5loOrJcTkh3qiHMkOERrE2qsLVtH/yiKZ8KoXaRyUvlX
yjYFbxuKm7Ik3Nenf5qkXH1UDy7YHWBNig1p0wkXZjG0IrUrGhajP0gr/pq+WAO1
KPpp2a7TLkaVu4IFcgGtdoTFYpjpMQ2xxhkeQEXoFlG2DxLC+izNUmS1knXG+75C
uXkRGy+mjAYVes/L3non3OVrwUf9TVGohQLjL7kx+2iYj6ade4p20COiMkLMQ4UM
vRR70Fucb3DSU8a4VIHkPBJAv+SFTMMuwZDUYSO2QzflhgeEz0WlfavnGn2YFApU
WbENT2b+4kcSNRrYUEgWwHpuHhSXxl78uqce5+gtlcERsnvdZ0pOqh4habaU+w/h
SisOQXfJeqxdufG3iCC41F1MXuoAeejR3MH5ZvA64+Vj3GJND6ITqAbAR9bmodJh
vbfz7l6UzHpjXWyBxlqOaqSC+RtClp6iJ3ekfpoFEmu3b4v+GmNGzppM9cDUijBa
Lx6FCSfCAyNOcq9C688kaie0hwd1Ylt72bkoKaRDJ7V6Y1JS1SUfYQzfWEe2h8aj
RdlEteiGv5hNGgoYjKecQq9aAizaGKFwQuTB4s1lHhcimbPsCotlmeC86/2unfeQ
3Luebgnd14K+TiaCdT26HkDNyhxO9BRO61KGGlxUjXrMfO4nlYIy65J/qMHI3CVM
Tr033ty4Pwry01baMev9OzPzvdjr2sLV3PCoYKnRfdzS5Uw5n+D2d0f/mnDVeFp8
t1Xx6jO1KNBX/qRysOOyBgxWda+CU8a0DWm/WYxrBgIOtXXMNHbp0lyLL/ONUZPc
V3tih5dOOPSknsQyFFjhruqqxwq4c5MTNf05cG72891cU4tk7WvLDU6bCkJOnDd0
LQCxZWReGalr6+3dIs4ZkZS1gPMMfhCLDioEFXiZTmXyNc7P6+fZ/oFtuokEorLd
6jvMQHpGr19Esd5O9N6dFR4B/Mu8XuxjmbII5kM8qxcnHSA5LxlMhIeCvWFiwekD
SduyeZtaC5wk88eQ0nKzsLyz2AhEPvH40gd5scrHU9G0+rgM9i1QSbSe1MSiFGrR
n8xwQwxxKOOg+5TSyiqkEQ88oCr/vVKC8VF7ydJFtO2yzTNAbNwaSOn7/7YpGBln
u/0ELx1NWi2lsNvcayldoB3ojGR/17yXpiWI0ItnJoI8mv64enamvN1Wb9cHaKVD
0LerGFfm7QeHo+dVXfavEcRo1XoFuQ/LknDqawKI81X4iPQuSjGj/pYLsoEWjdL1
0bOW1qkKS9zR6RCzVp2AJ/fuNHkI0Eus2rK4G/LNwOeWzkxWla8/6lvotrRQBzT7
MHdqrkedD46urpLokaxHpZb+//plg/4T8MWboOQCA1u18hEPuguwAikF8wJ1yVkP
bl7XygPFnC3nXiZNiuUWx1VqKLzsB0u0LMyL7jGYz3eoighAAH2DhQcqhtK8nmb+
EQ5xyOMAOpz+rj2JYLTrrMD0VD5+rdxlSpo3k95iBXdO28MI5+mfY3NRJ2/6d1pw
ZyYJ/674y6cpP8PlRo9lHqjsxexdN7Q8t3AXl6Dp0fHpPnfQm5wYw6s6pEQHIh49
RhNgAea4mFK+/T+SSIqbcS8+jLwo52b4nZbKBMyb4v8sZMWsgUaSp9bwchRNqiMQ
Yeng0+bO4toT1Qw++i7H6aNeh+AF8r9XxLFO+5QfrRMHsYEaS80ez7zkwk1J+Qbj
cfwrDzlECpXX8ixDwKNeUQ+rUhTXmkshzofxnNde9KbRYU/qJBSalpep0B4eBRBK
0Ucts4PCZC+cT3niPCnpWNeZ+d28j0CJMoAC2OlYFG5F0j9C6QnzDMkPr3s+hpYp
6n9QEElJSL08aNq6S2vyDGWJia5fhwb0J3I4l0ukzYeFMumAzQhuNett00Bq2ybD
3N0yO4fpgetKXN5SimLe6Zhtp3c+Py364FNnvKtdiY1SKVFXVHEvuEBRr9VQEhrV
/hl0r21CYs21Tquvby+EbNkP5wkaRdAHZ/bEVZFFxipuTbl7RpMsfdkXRRGEy9we
uabCvuDao/Bidx6W0BYVcV7aiFSSuZ+6sDlur3CRPa9p/3StnMxS8e3ilMFaMgqk
lRiBR8AVv30zI2kmxpaQt3MGbzklCXQoZVWvgp8cFd8jPxgqzcObX9mgvDjnsDxP
AtKdYeBltX2vhqjsYmN9hHX5ksmC34CQIXtkbA6FcP82UJh6U2q/OP/A7vL8LdrM
UXDyzgpiz8S5vdndeJLv+mMTwb51D5fk5UTqxVqi1lcwJkPAIQoVSt3NujhtkTsj
EGmpsoNQ/taYd34THvNEXQn47NCwNIJmBlzW4uKGkRDVPt3zz7MJUs5Dk3BTYgEt
c5E1vs3JhoBgcItzF1k3kpIEgO2UvcR8GNGFNNIXnYwrKTw1w30sm0hTEpYNvCWv
Y2pVW55zdgXnSmwZ0dJ6QRJ8BQo3S9MJOi6UUCvRS44z4X1Mdaqnq3JDX2W8Sln0
SxEshYh2CDGA+tEG8mzyw3mPyn4zKo2r3uO3aVTXwJA6/b5VdRXffL7bUyiJNv0b
EN1yKHGKY94XEoYwmsriv7bIz0zae2GaguwIKw53J/B7TMVLz4TB/o9wIJ8n8ufZ
W1OX0qPNoKDIsc+p5w/AJPob1VlfzE9oJ5yXS9VaL4WNvTTM1lb/LbyzOuT7MWpv
bIszpDEKiwNY6KbOGZ9AwlrisG6ezp48Q+8zhxFzuGnlcnCy9JXURfCgv4n/Ww/A
oeJpQoswoPjLeJFJa82OY4nMR69AjbWoqeLlT51RUJzkus2Pf3F7F2G2hHxF1Zj/
pvCD8+kW+zgHMtezzIv8HjZahwE6/v6wxkNhcZpHjzE3ooZNlM3DoOLqf6ACHkFd
alybvuOiLWn/TlBrkIHieAuY7P66jG5Apo5PmX7tsC5OPqykZpUaxWvisNQU7zKO
1Y1QH1/43LIiepSUeyE1KjjmDnSGPWE+atY9Tpmvjen6/gn/Bg0fc6UCzyCrm/0E
sm32+/44aG/SV7iAV4Yx6qnVuXD50wcu4kizeX0a3YYVSxcrpLB5VBE4bETv0O3y
SYx65c/3cwMg50vrFhiZ2x9mgtiPXs4I3Rx0it2puEeDan4uVwXmCWlPIZtyhDS9
oibtZ1f2ZTAlRukxePz9F8irOlyjHYyu7FCohbOITeKeeTftvOI14jgfgTh4XOdv
HAlj1mZcoeTNpngIAE8nudYo4W+bmRgCANumrE2sygAs2aiySuYZlPzMhpmrE1HK
X3L/5ioYqqv0Gse5exPLWs8kIufhB8OS82QUk7s5GT4QiOrobeo+cTdntDH+gZWh
tCNlf4v4pANTHgYbNHfpZNyyXb8mjgu6+ExbyW7XmEdU3klT4zPAhD7yK8VBsXWC
i5s9BAuPgvX+DRg3AVC11E6SVNqJD50pJ8wPyS6HlzlcWFGxXHw5R1Hpxqi1Gi8J
gRiqTBtXRI/jnO622U3OUxLCpMN5X30W8ChKmhJ6vRLZDj/ZIe1z62rSgR37TiRu
zXznxSjMNQ48TfILZxBxOUf42wJXptDBt76uaSkVT9K2bEO6IcEkCu2wPHSAWoWy
L4tswvEq9mbjO9tFfeV7xloHDRC819FZKwa3avNv+YKjBkiRxSXZWYXlyVQRsc2s
+lYmS4SyN2cW+EOVwalJz5rW6foW4vg3i7+sOekvUX0k0sKtoA1wgJo9MEJ+TEGH
LUiTKxdxIxgTFMyRa758emuQj12EdfFIpl/J6sc5+3RUZuv+bfMRugUw1QLe8Fcg
GCWrRI4t7h6SbZ60RnlJ8IbLzbcUFbXiXLd5dIuJ1QHcGGclyTOzLYdpmYuxjHJZ
V27UN4sCb12KDQ8KF1+QDnOsL4fTSDCpldsOH/TajknRglmOe74ch5yPXiCL5y/9
H6vzCNUPgQCWIklEddHUllCSc1OrYrZPdjjoXpTlmv+CS8NK9vpX4g5uK1kCcqn/
+6qD2lDlGfoXFDEEY7hp3dQClNrzhkyZaZCDZ1/53+LeYN8jIVeKqRzyz65ysi57
5SBfcFYLy7ozoAUo9gD5ozK5L/Q1UsVytj+RlYGqbBaVGvsRXOMFbTbKDXK8l0Te
/9ZZl9NgyeDiXxff9FHl2bQPyOrLhdcnGwfQJHFEJV04uy4XAxLr8gdNTxmfn42H
53rZgU2b6igNp+t27Sy/jXzrMwpTe7WoPHrPv3qcflpc/53Z8t0wQJdlrTsM3zWg
kcFaLTIkfwQnyAr4/St2k6xZli6f/9oIgB5rkLjvBgpqT+6PWFvW5bK7W6aiXeRn
4CY6ZHSg48FOJIZwd7JdepAJh7n8+vNnIFbCRl25YJxuercLECRUCusHzm7wxAf0
YynwKdenuH8xGKdy8MMjp6YyJUNzdNl+JCMM/fOq3YJwW4xOSoPvKnCHK5pOE1Kr
i8NJqfNvTqbyyySmNoOTrxQowAP0Pn/qlaJAi7jycvDnmmGas9nieajyIljscf+3
smtSOQplm2RloxOJamEWSRmzYWYD8/tcAJGdSjFBNyd/KKthfpiyvS0P9TOn3OQp
Z00Jd8NzpMrEvozoZqju+M5Hl9IpZPZEMeb2gATzl1L5+wDg3gqDEirEVoT4zToN
5NkASNgO8gqyx7DrPA+GtAvk8bFpimpR/P5B7CczeXPYQ4g52qVVpghY5aPpXjQg
2jhfjyq++ygY9Ij3F/XjU+zEwfsmi3icMuxQ8X3rvrREN9mrnWoH12EizvoqHKnP
R58BgBlqzt57Nqvg9PHApa0N2kY7mZum1p/ZqVUXCkGN49pA4VnG1WcRNwhX/+7a
iqbmJit6k6Q7D8UCfQGCeCq+osVeEaGgeCcPJMjH4CA=
`pragma protect end_protected
