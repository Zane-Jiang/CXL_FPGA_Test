// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iQS8E3a6ataJcDIScbqQ7dLaqBKoDHi63gUXsJrkF6aN/1d+m9tZ1HfkJRUB
K+eXQNFcJRIVdXYx49ly/9OwG2tLK9bE7kCbaIZHxPz5J2Gw3oRcNZjCl1ms
f8ak63/lxWbdwEMDSlwJQTpsPmW6HwSUQf10YNUACxnSpLPtfyQb+B1LrEbK
6E5UvDkluJUlJ1OK/dfyiovYpeh42dywxTnI6WqwpxE0WvozuqFMO7VCGsRc
wh3tHsXlQQ8i1wrfqsYXjBsPxx3d1lSSeQ350n9Zw86mC4xjFqI+mq8tt/3d
6ZZLUMHTBzCMqGDCeRYGTOL1xpzVZNnVOW/LQSb7Bg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
osGN2IKpsXeFlv4+r0XWE1jk1MsYYkexmxjII727KAGQnMvqO6E/HxiD0La1
aRezPPPCfazUXVrTEJ9l1DmJmphEff68cV6lsgEqSZZAA56xnd8LLTxWw2Ml
29rpAOnbhGL1L66LUkEhgn0R/mN+tqYxuvRnfJ53VkYRAvoYfskiIj8OklNk
/XIbW0f0OiamqB8TKYtTZCrH6SyR508P5yISFtQLorsmAZMM87wnVyYCKDfC
Rjv6wJTfjHjceuIdR8RDedj99L40NR+ANAvrmXKyoNA+P5I0jvVtbOovxbS5
TaJba0Aof4JbxuPKyJbiAxeqBaQMuulcfYKrPstF1g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Tsswj9C+thPOVAgQHgJ4PrBNDf+rHDkgNXRpufP9A/dbL4QDh75ICcoIY9LE
IkS6lYXhn3ZNXb6cneHN89m74j1O1WKNRCJ/AfZqanATSvJ7P8l+E1xeMbFf
JwgN8AL9isBnE9MglZzxZujuNKnJ8Z96H2B6QGhK5Bqgsk1qY6AFVBb8p9tw
hidNpDayVKEtZxiC5tzFkO4KhWyNJ7i60U3ML/bwT8icCQc+UsmM0Tjz28NH
TzWoqrCIyZ66oWDJdQSG3tqbYpW0ebNQl2ZwgLCtsY7lxOvLgkFqjpUfSZvs
Rq0r34UXcYEknUXOmNvwEC96KQmc2AxNKSAWqsqw+Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RfNsPIGqGzS56nyg+HcwYcE9CoHxSXTt0Dmpxhqiuni579+G6TCtegDF5bpq
9Ryicw3qlCWEZgOOx/Ns3n0QdMBWpzVGjTSOvRh+L5dMmr4MtWw0Y/MhfhII
os0+khcy3SO4CN8+j0Qta6lv+UIZFKJjGYhdxAmhcbOZ62aCCHE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FFVOsNTjjw+79XuVEFrHhBU+13qw1IROTWyAqM75BeZu9E1qkCJVu2269yw4
HP4xvtwA3KiNOHNYvDyuDeQuxEQYHQJ1fuMYZwsABrv9J8jpegqaPUvYeBkI
O1njnhuj3VJNnJg661ODHfBxR4b7dfv+b5iSa+m1SMZenhfKdtZWnfYSzjUa
TuCl5XctJuNffqwcp2t/t2lulkX2Nq8GIGkymGy2ySZBesxiFcVY+/2U36hU
1b6nHDUBVnny7WI0RNcQomvuqBIQuQg+B/emsG2mPf1K560j6Wj+oCuuNG9y
V1hguBmBl2RhclSIZMf/j4QyTk7pxVKB6/MHjFKI2K7fGOqzUyGzWDuDO0wi
XggPDfQOJPY5b5shIlZT6QnXbKG+YkPWlqvPI1TifPiAyL7LCh417CvnlHx1
OJ/AJvobB0x7Mx5XvtvEYasHEp3nyEoaZLow1DGH14gfxVPMXXgq8jXgmJrY
5wn8pRMHNfPdxK9eMxSQzzpCnixnBdgd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IP7y5XrQA5wVGgcE5lzrqGUsZFaw7z5XK7BDfThrHyGwMRdROZrNAjTICinl
mO/ZBVWYtclVCRrbbIVupt6hemUUfLW0g/fUsE7A6En7KSSIUV/KaVaLKOnD
M2OYtPmYp79JwhkReAxy1cL4WKPd6Yg9O1D8K2NBnGg7nkmxzaU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ByIcKT0/SWz19Wwcr/ddbQICx3yIDKVyp1OLvstqFPDU6Gl5IFLMTRNVDQWE
CTuKzqyL1M5i6q9MGtw5+jdB1LN37y75GkRMG42oPt45fjyW2h1vHwXbz7t2
HOTM+wVdt6fAbxuiObJ6Z9y9E8CEGiPMU65tcCUiu3gE9rpRN38=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1040)
`pragma protect data_block
yxPav+ow9JZ8F/mVtY7yzbImHou2LajobljTSZPA8aUsNde4Ir00VB31GWDJ
9XMS7ACLPC2Nz3Gzi2OXp8cTKL/v+AOkOokp3PjT4kGA6jOAEoV48W8LEakv
bk/9oGFfaeDX++4HiAUDrboAR2MwStwnNNZxMm/4qOkfbyoAZjwyFCcrz7mJ
ERKHzVTaYyU//d9r8q77gveXdSKQ64EjFbQTPB/DmjXCl8THGJEs9+nHN7+r
0nXjhgZKbM9g/UP6ja35elG8/OIwKg4M6YjuPGTKZKYk4eiZsP9JnY1bskQA
v1Y32ac00nqyNiHU9rYcDjCS6DOq27WtlUNXU8zlQOFi9bBRgWoaJvYEfdAA
o/HIQZwT3UJG4EJuBtRRnklCtEE9rW0or6Q2Mgc4+JlJkonfUM+7QiNRztcz
iQ4AFOrRlAmIaGiUI31BU7PcAfXMxD0gVEIIcVkMY/v8FnbdfGQqd8OFN0eA
SH12R/JhKB6g/J75pT83875eSXE3itx9J4vwkxidadIIaDs0Gk1spVF+vVK9
Jta8fIyT+ZWZFy86N0a3cqSnQpI7c7Ipcvf8Yf/kEqkrOXFjOpNbHV1MOmsF
3u6VzAE9lwxeoAYBy/NPQy6WVpz7XgioYHEiGRDbVQFVJZX7dfPI3Ao/q7Xl
OX+dZ/OSdhIsI2UV2gRaVHa316JZEQx/TFNgg2LTgmO66BDs0riEdqUfoXfa
Axfqj38nc1h6RK3nJEm4XEqIHJ0Sly7yhyjdeyslRCxYzzxbgxWYC5bAlF6G
6Y2V4XO3z0wuTi2Bw2oPXRkSbiB9y6CgSkauQNiKFx74FQH8KW5UnxOB8F6x
DHhzyMUGpbCfSORkpnOazHI3hDS/+WxeXIb9mVpdKMFw9sETcwR+f4wPe8pn
3k1iqYvz7kvlIBw312vct/fs29zh1X47BZptW3znT5qm0ikOKENC60Oqndnr
9O9aA7AVMkWYFilHhDDB2ZQ06ahMC5kE59s+ZWxuzLYYj+1zf0dVFD+GVXYP
eUNALHea1pk+odCrukhq7FGlVvx+/9Zq6okE14q2pk8A59J63sZHHSwdKQys
XUBxdYHkAreZogRAQPvaHWB9uCusGBYN+n6/Ap9TxCzd+t3Woq5VmjFGfGBr
z4iaUVjkymhZPF22lMcKD5qQLlGL7m8rhbUIkdo7YHRVZZnGcX5TB75faYPU
rJjNeZyFeaYSOv3oKkUfD7tq9pgHQb3bFPjxbfUqdE1Yau+YQTk23I5GrjVd
rDGo7gmGwl6uQfMJivmz1PMiKDNa5A9U3QmU/LXYdydXWv1zdpgIBx2PcWDZ
pj8m8YWK3AyzsLKQ8gTQX6rWQGElHpziFu1tJzziVzfShiVq7tDsd7P+Oxx9
DJNM/u4=

`pragma protect end_protected
