// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ncDNaR0DN50Vnqn96cLyEk770Y1mV01Y6LC+FaIGmE5ij16TodqzcM1kmOiMoZwT
wYnv4741Yn0Wikdz+cYh9GE1B4xgQtGHr3d/Xxzkx04JffOkIqDPpb79alN2vbuH
R3t/77IrE6qy7Oc2jDrT1ciIsupQwsFK5i68AHdDnCazsxaHbHAK7A==
//pragma protect end_key_block
//pragma protect digest_block
Aog/r9WckL8nXYri23kswGPXi4U=
//pragma protect end_digest_block
//pragma protect data_block
7cz0UoOkIDwD92X71OlSrsZexq2TbJs/PAsmcPqxolpP7H/1fld/CQPc7eJBkcam
a8ez2Fj3Xjt/sdyfAQumx7tRmafVTdYphvBi1c9Umx4AD7HJ+/XXJyoZkz3sUZ21
mlHfqUUY5gElzRc6Dts113DA5YsMAe9QfUSu829S5xGNJxZ/mCjETdsy+M0YZP+A
vo5a7EBlqoowIoXXuHQHP9gnAOAgmfZSRcrtv61yzHKDnzZAmeGu4Vld5Y66NKXC
Mctm5rtBrMDBt054XOapTStDHzPtEk/dHP3mJ4H5BL+zCB6if13J8a7cjcfUY5Cm
StPm1bf7eHm846bVX0s81ntqPxyvCOsW1mqVWoX249o5x3S4L8QkHaoH+Rb/ADNo
IITGS5w+kHkTd1gGBzutxyJ3dXA2suFQnGLeaK6tVGDNEI4CC6U907kSgDXYi5C/
jU5Nfbxaa60KQijgddv+VEBFRpvCVzEXeq0jMw+XVdNTvIzIl/1MK00kuK1JtGAe
tqBEVzxT0mxP1BB3TD5/LxlfnIc6JSbsCnXG4xvpLrn1Km/lQf6lpOv+5L3BwSrV
KImp50Wg//k+nmW/NsbYEdninBlfQGOr1jj4Clj7SNzD2l5Cwcms6cSf0MLHE0iS
A7VvvyzdibT6lKKg93orgHzKa1DmStqttkD69hsx8fboCZXe9cKASs0lgJT2yz44
3J4jDHjYWfRIDlSC1SO2kKiYyHSpD0KQWrXHX+UqQJSWTwyPBMvXu2dRhSzllTAt
dDzpwArO5D0sojqbxNVLgPMWl+uka0YlxUFPUfckCdWFpYvGII3/W5yvxKogWDgX
nV4t+R8UZEO7Bhqc3EH452hcR4DkfCFC1hGb+tZRs3HWoKk6Gp8iICI5+LXaQVpN
87n3Ri96GXC1qIg/7eF2K7bwBNGQqbGikr30VAcbY/r7SjjP4eubKn55ZeGCX6zD
l45Lkv8UqUAeuCpObq/jq8lucyA7Wzk/zG6JYxi9uifa6d87BSEvNDj5VUfMwuzh
/ivAw/5R+S0HGbyIoiz2ZjGbaTznybCKVX0ecriaH7Oe73079/isFiYqED3QeCm1
atBaDrhQLEUuz3hF/eez7ATc/gO84qcVUXrOspHTzt/iDZraKDRp1nNxi4i0Ct6s
TcaIQDAGnECX/ctjf0Cu1BIt/lMObFFXU2W5SKSr0kaQp5aOgS+8R7+M3+o+h+hE
ak4U6M3YGj5X2kUxkozlBDz66gyCWmwXp9DnAP3ewt21hDi7QsDmMbIrU6LEOi7A
Mxuu9WujHj+laTHJ+PW/PM5gh34PCq6BLrQy2dThPxYBbBcNp9ZSJYJwrrQtiuG3
lnpW/P7Q9wgw2MahXbCS01VXhbghoUhv2N0r/j3iyZUq1oZlwgdHwA4WOnpenFon
NlVn5Rs2L935KaGUACz0CDr0pphp+QVKvfA3IZaArrkojjHSsCE8DQA7fIkDvms8
4cyPdikznppG8iUAFTL4DdKCGQL1jQCrTKA80aamiXqYsDVGJySx59s0gwQvkbiy
HmdUnDgPgQ9oG3eo4UlW4UvsKKhLthTymjVhxIQrkgOFD8v7R2UetF1CIoJbDizh
vHb0p4+npg6cms75IVy0bixJz/MNQufbsYBx5o5Xh+7i3u0nlXqWhsBM/kU1i8FJ
yLzLDNpOZKpt7woItINbgnZeQZmz2bx974XoyLV2X6avKob3+z3F1Xw4GqNT5MQo
l/hq08CRKWvLw4w64/j3feDezIiN8P+aAy8j7Qu5/jDDG0MmtEsAZfYSskL3S0Co
vDJ9BPKJDLnC+tgmDHMx0Yb6XO2SUxmbJgUbuYNg+riY96k9KMOROcEYMJpgXqzg
Hl5LqrPzL2vZc0OS547zYbxJ/CYMEBR7ffkQ0UpGA3Fo6idsxIvS3b5NRQtn4tSI
4ACt4O4YNQnLKFEBC1MrjAUg4QKWjZWILyYcXZs5z43LHc2Xof4sUhomrWQLRbuc
hrQjOOHUOCIXyTT1Lu3DIPe41vWWHf90XPYZLDskCBUhV9f9qUWaOoQYKd+2ZaMa
+RfUal3xTP1dMXXbDez4uElGWqRd3Of0hdIqK7BoM4ZIp1Ix9jTt8FbPFagCI2Pe
YVKyNYMY/wLGdnPTfe8l8tppOk9OKTdBlVQSS1QapCrXY7tOtRLgAGrYPHl4Qm/j
udSoh/MWPzohl9ytpDiSBkhdazjaDRuxmiLp7s6am2BEz1NXds1gYGJYaYrVyjB2
yDd2Mj88LZFaU0XcAqZnVMR+A2KH4gS4VEsGeQO/qkpX6Io65D/IwlHIWzIPSDiD
kc3RaAaasfQOdsQ2UoV4qYVVz3UHWPcOBbVVIAK9HaV1rL9MNZQPQjSC/lPBkTjH
24Dc1xV4cx7fUHJ50C5Y/rsL/5RpB9QcHHdUgY5TMzqqONGjUoegEf4+BnHHjJRr
lr3AdX/cDn7RyapnRThD7RWYekPzIwhz9B+rnwr2tLqP338b3GqOPOC0F1s8jtJo
38Ze71WjE+3qHEHyr1iQjdfiOGsJfmO6T19x239vm0WEllzP5YOx7qA7Iu58h5wm
HW7iKfr7NcpFJhJMMkeNesxbKTXa2jFuOSgMpAiAsLnv495tAho1asLt8NJTX6AK
oNCR2gjxhMz8mHD6OTHUX3t1Ua8imVbZghBq47oxTwMW/KhTQWBEf+qrnODfymCY
OzZpNoY9guF45gk+i3FbJNgQg7P7DMPGZ1tcpt3h04zlZcJpcnTGVRHpvLLs1iFp
Iy98Tq8RheFWPN7XG1WcmijiEVTGxe6JVfToR7q4WV0Jo3CtM6p4ilQeOlrWBWbb
SO7KnIsBC6dT38ODiaP9yd7PPfOZ9TVoEpDuwBVWfQkmpH6b/7PGOP1IiRmCL16N
8Ml6EgjSTolU6VpcSOj/xDzf8eIFvOOxOUgjA64lsmGuHwfeWmWICrORTDL654Cz
dWesSBiHjAV1IGK0NhcvVg7Jm5bTwnk7seNyWvQFNY3kxj+K5TdGpXMa1rLL/NEz
rXfmb5vjp3bm/2Fl8/5/uCzEfbKBCyO7M8UE8ewQyz9C2qgkJfs2j2UmJT81KGOK
xnHUi7YqaYkBoGT8/H0o841v29NWeHE9v1Xnuk9BUqSEityzudXrCIUbi83y+6YK
OyU38N38B4egzAs9yzFoaZ1UKN/hagb7w3ag6XOk5JMsL5pGY5wQ16sJI3cfo+xA
i8yRwhVt/91WOTm4tj0UFqHmPzg5VoRrtyMh/e5gATSBrlQi2kPz1GL6iKRBiewL
qQjd8OTnmk9Nnx1gqTHlDlh6MHeN9LeAQDhT1aIfzrJnXYZ+EAMdR056UPNk6OU5
e0GAIVdoBzwKbB/+xUJSkVHe4s59QeqCkOU23gKL+7u2totF9tLQfjo8Neahk9hk
Uqp+MZ3tdYsMWJIiyyjBYzVYXkkcB/PbCfSokNLsaOjxMrew5ZmeMMCnaI53FFYn
gdRGKxIUSVOMCFSmZTcM+gy8dgpczXJNrheMBJcdwiOKNeoC3ReNSxagIUfGp06C
nTi6ElZP2+14HK5n5Gx0U1ZOjX/DyA9pVfVVfWojukxf79S3vm+TN897yS1tN8VC
d+buJOiEN1chDa6pBD6S4b9Us6RrZHQUAUW4kPqi6x711eqw2CCPpXSEDHAZUt+q
t9vlyat7j0OSoEOG2zuA4cZgERaOh3+fixK9+R3/DdKv4e5V88y1ziiLnKVswA7O
ZqWMaTMWO2M4QMBXOX1CObLJ70g/zAaWuJYvviu7TfxeY4PShv6B4Gzxjxxf17CV
u7tSX9fSI4DudkwJkWs1kJZBQDQxeGW8bKPhTw970ElnvDSTWXvKw9KyQmCILdBh
E609u5thtHkAy/EiV95oT7tKu4LhChVcXu1sTZPuKogEcD7kIdbBKWiEU0Ckb4kk
mYx9JrHfMU3XAEdnskJZw5bv8uMLxbyTjahG741l2wGLDpcmwh4JJwDoMdDztrtv
KK3ZwWk0ks3nrqu8o80E2UexjZ1l5OjKom0JveAHBE5rZ9mEdE3bdhRJdlSxWGkT
jwB0SSPmgmCTibvLyrwUV//OFXiLkLf5NJ8RTqTyiB9rGAIRyWLOZG2edGyFlYNq
BgQr+jxCEnQaI0jaRIkuXyGaFLUD/pYOZAu1pFgxs7vhgd9Ny0i908Mgr6yiduLf
Sjs9zhyUbfBkvbS54YoXBoWbGVv/rCsZ7mAwIA6lY7n2mi+IqtAQ5DTLPYxSczVv
yglHA+K0jmi4rGI9rOFkxQ63cPIZCdkPsRvM/ScPf9dem3Fi6T//KToYQpplTNhn
VUTxidokA41Ih4us+eIVTmspEQqKLlXBwaSM5IUxXQsaUqGEOfOiuoW7ahe1qB3q
EFDcRuEJgOoPg39GMSzupP0wzdvV2kQgo37jhLcy0dwUnC//hIEQPCF+klPB4Fvt
/12nXiacFYXOGqkY1YTx4OI3Q7lcpeI8WP+//pr4z+LFGZp8hmbWBLPlP026CurO
ZfvpYz805k4KJTpk1/fTYcrKd3Mx7V/PTzRPPPT2N309G5EJPKWGlbc5nhHckOVA
w6gopy3cQQNdpaX4mKVVfFYJBsn7ft2AJ3r4iaxZUXtwtJb+dmBIuECLbCeql+8X
511A7cMCST3ymFczE/U2cdiWTNa5Yfx/FKxNOlLbjYiDvKNM+vvCUz0J0xc2PwtP
ebe8NS5et7ErSVd3iOrVfJbwkK7cex5m+rXgXX75u5/YLAn8G6S1CLXvXi6/Rnp9
yT1BLwqEeXDq1PDRgWMa2ZaIdXpb2fWr1P0OaeXjGLYQ9XLVN+KTVhtPNmmNIjqr
Yw0mYnQXJMh2p/qWDg4hgeHMZpMZG8dGxYKOyM0/xuAHXPs3zgFv+xjQ5wmSDc9v
iKvHhVzbf8vwOMutnHzh0ayhxp6YHx6wF8IrGYzf1VX2Mak6HCEzP6hI/54P0o9M
FORIUELBYGUjjcteEZHfpSmOuwh0RDygJ9r6V8H5bn0/Czfw1H4qZTSDiQ2F0nD6
mONZPeLmJzY1tSqfCKmD1us9zgepjW/pQsEePjwYP/YMtgfTucrwX3bHtn+MxU1N
9YujCFcNOS4Bj6lHXhoPX6THodA9LVhBhtL4cCf2ZbyRupIol2EYMGNbdzSfbKyo
CxlSfVgsOlKTS1WLTHadYudFep4mlIN51s6oUKEavYwWW0q+uNYNPsjb2Rf6UY7K
0bCCFZstvX9lX2o5xDpE6ky524aAi3oYtMmfeLw5ov3f6t7DFGYxo1tEl1zmkzim
1ND0NaDvQOWYgWS1F58lOQ5sP76J/CD3ldCKAp5aC2UmUBFKodVQ30sEgVHwkv8P
v8s25hD9tEfCX+P6sCyEENcXG37bWKRM5t0U+gNJqDurKhpisq7KV5G1I5YWo3re
57FD5gkD5IYcVkpYujYd9zstHCnKTCDFHBKWATIwOklM3mpfaDx25UM2/2+synOn
dCyC65TUPWZUt9nEOIbBg0ISjwqOTc5ljFvg0yJnk6h9a/KAyZ9KzYHephkMyh0P
yiiCGs9Wnkl5ioWZWACQ/tWtO37wppzdCpS35XdZ+ukeNDjujgNu5K6clsxW2W+X
qLQEkIIOxPQCf81EXEjHAIEqSMPoGcbOVDn0FFTxXtd6cwN17ARGDThj2qw4iAYW
vkIChHFHajWDMrKA+IMPg0nUL9JxpBpoon09NfF4FtpwRCoUJxoll+hSZ2dmj4Pt
ifeafFiMk0tIOJ1DNCOOztW/xuWV7OR3AwK9bJ5D4u/kNDpKIIcYZNlGhx2zwJ5X
8bDretcKg7lidDzO4oBr9Ri2C0k9+idO4alxggYZxCBc1jZTpV6ixOeFkUHtI4Zt
gEvoR+/I95kPIquezRt2kaNAruGjqA4agh64hZbvZ924enc2cbUzh8rvehdu6xAk
Wlc3G2NxcyCSQI45O7j8Vc4/pFNoafRSHDmtceqUyShWMMd3/HWUKMJQWEb81myF
yCHhtMnB3gQjoMHtRqYdtUyP+ti+Z6M+jHAJvxrrfS2FW5ZKLEAccKZE9w62mTw3
TWTFP8anPZZE+u4JmtEqX5ebdG9rWCqXi+idP3qxQxiie9famatQYYblgFjjz0wf
FTfwRk8/3Rbk8LC1BH8DAxiBoOIKgTi3vtG/MiobDjNLFdVHKxJGEbpeYytxSKdU
Ed8fAtDmpbvkfyGPEDg/iO9cig7wTNv0rdDxGXkn2tS5EILcior6iiMIj48+CwUV
mSkuMg3QDMEZduiTXJq5Kw/Q7SYqAeNfiE3iAUQQQIawGrsG0yGI/re7iE8LGQAz
fmZqO+KyZTsmzafx4qBS7hIhRB8azvB8iZVJmc4wVWvGbWGTuMzRW27uKViEnVAg
DVgAgtHwf0fAmQCkHeYuuL1daEF6NG6BsS3ycaHZjX0WEyrhCkrG+sMnzht4etf3
eNA0S3C/IhRELQzKRP37kV7tTTWqD0QAZW8HHfkZxns+g/Il1/4DdSTDFuxORlIo
tDty2dmxZMk8ZmFA7mEX/wATJlZtV+nzrr0DOXhQ51zOPM9mXEAo+z5nfLHeCGbw
kjVs0pEe7iQqTbTg68tzwXzEDC1a+zBqGC0UGRWXVdkCiXfh4fK2NIvvzqzk2GmF
HPR0sn+iqxUt/Hw9Wp+oGeNusPhUWynWqn6hUkV6/LExH6lfv19Xv3NCNbaAlzIS
OJwNrbxugp1AtEB+VyEsU+G0NOMq1uM2VmaJKgpHKjlAgKN+AcH4csnKciaAPx/X
RwN/4cM6HAMnxBEgoYlZCwQrpSlNtcdh01mXphln59c7Ybf7hO5RLw5zmTUx3qU6
Sfg3BUdhwGZRQXyoh9lWPbnVGM07XizwP/sxZiaOPeFgkfU7KXOJDNMNdcpwGEIi
JrqRCV0u4tMQKyi0DUyTMpFuyP78HK0uuzUp2KGvFFwyXRTlh5vVXbpJ6H0pq66A
VpU1sbgl4tqGunBeOZTRvnVjPxGFLu2HhFkI29gMjLegU1e/wn3UbYHjHnCpHrAy
xiHhnhX/bDxfgF3zrErwTV/K5hktlU2EcNuYu/1nYIuNGaKftHtW1w46krbY2Uom
bmW9kZyr/w6pIAMNnKeFlNLVy7MvXCBqf5UBRBpMk6DNi0224lKZPH7PxidEVjmP
EsKh05SUCvFq7TYmWFH0UwZeD3D2MOgkzYntNpVFXFV5TgapqOl8Md96pcsZLwZo
yLesoX+ue8u59hRu7qPL/LOh3OFbeN9kLGM/jw3U74TIQhdjP1IRtGIAq+tJke52
1Rjz+Z7OQ2M5Rn9etAsA33V9TS9pPMWJS6K5gDhkSdOSEuzOPpA+nE72g8T8REzh
ObwsHnoPG4jgiLr4N8577PxsRoRk+IXavpQI/nEJgWd4TcikqXfn2HALPw3rpT8g
AqGU5U4Ze5NZGc5tVLEAM+nlCgKZAmULo4SIXwGr3RCQbL+gGkOuNT65CkldPY7C
H9S17bLGsr2UAYvuMin54oEsU4WR3Naj6iRxHFPoI2RgWtpWRIjRpugPd5AdUGZE
SmInw9LdbrAkK9r4/0XhGtQnp8SwCOEdhfKEpFjPAb+XC5cYUH5T0Scoyx61hZmX
7dukF5VcBzhQmA1aO6QG8mI4LBdoVyiozMhA4OI456wPt2h4mB6mOgzC+GDeb2Q1
Najtdhham1oVYrbj5RdBMa8FItkiKmND1BaWf0n33Ovs5yN47WMZ543AgR0lRIQe
GCZ7Ol84IxBip5/N8mgFZ9k+e2v1wsbKtc1x3eeVRAMke/32Vo1wgh5lcuCzUnvl
2XTwoe+vdianOrsPuNgb6ovOrmiwzLOYeNAJX9I+0MSrGMeeTW4YqQ4UwD9A149D
aJqOdLKhHQWuCVvWJa1I1h1ADDpo6AzZ9fUMnuD/gjWKeWchoES7UMViQdFhuNb2
v27vw8I46ATl+eDpVaVd+cGoGhji/orLfUcDhTvGf1HSwhIBfZ+e+5vY5/Cp5wOD
Y0ESRdBl6QRWSr3X0/5EFbXhi1pGzu2apCFUs0ZtXpkW4y2Ny8KTfXELu1UTTaEH
W1b4F+SAYpn7zpBHvxJWcNxBZYJ/eK0p3G2au9BCytTIGSC9XXePQ9xBFDQSpRNe
8GgEmBmixtacbUEdyxVciDqJaixQvJzDYF3oVnQWYGI/pciO5+Cx+bOibAnSryGK
4mNMB+v379Ooewl7FnhtnhK6Sy8I1p8n55filYn0OlDpHToRlgMLbTai/bWmV2ql
+0+LA3nKA0vi9yfDGQBoZfXhKm0c7hpTow3C56bUAiIKd/vKs+goEWdOokQXH/fQ
EuWhnws8diNeAw2Pj6q88G3K7dlxP9h8Gq0Qpxm9n7fBVpOXqghNoyD0BocrNAPP
uPIHrreBw4vy5c1DJZWNyX+VO9mIs5uA/5IOdFBLq96/xV3lsXUeEj1tDWjr7oIp
6ZWA3fcJlXvt8CUGkVNAZeOicvBexqavSRcIyoc//om2/uqQPTN7SeY5P669Pex7
/NNPkBVtF8LRUeDr/4lhphBvfkn6hR40sEZZv4dShA42Q2iZYgA9J3CXocuEGoQ8
dovT9qz725WHmEMWPYBvc8Rae8vfbqAx1GOSHVfNA/No9+buOj+V7Ohh7tT+DaB1
LfgR08DMD4NlCDjBE82j5mRENmhBg4ZwFpoQfQH8P1hWlFozBGxqE0vwgqR7+5sa
sO6m0lqrghuI6oAR8UVp2Qrg031HTVOD7XToPXE6rAzKfZ+fMbQm3yOC5txCF4eH
Mv0r8/l9p7u9vm3At7N56Z37CiP1h/uP10cMfpyKGTnR0GaEJ1kCCG6GwzL0evWr
TNmFDGQRz1Krpl2UXisLcPGGyk9KsQQK+nEAPRRMBxTfhXsJaLPcLIPND2h3OH5d
SQcp+QCq0nKeXqA9AT6KRq//vIfrEGqTU5od/9T2+h7pgyrEbktFzDZ34zo3LJuu
cVwWcz98u40jq64S5ewK039sN3mHVPBZMZD+qMTgjj4Wx9/UAnYyHKuzjW5ieidC
F/sjQO4fXXCnubHrmis0gYd/AhiJd/JgF1oDWBw2ctlrylVKpC3k6WCD32pSmpcu
Ckr5wNLE73siKqc2sAZjzTVT7MLTKLHQqOQV5Ze4HRZwyi0RESPyIROhqGYuWRbd
zvvvqO1e31Ys8q5rWtTM3g+EpP86ZvaS2Q/2md+C8+1Fk6np7Ls40++wnLwdqFCq
uHreIyY7bjK64PnayhgpB3NNq2E38xJpxwXGTUfnOE6z45aLbzPlOltFfiomgVYa
1uzoejkyocQ+7LI2ypVLzlqmLYuLTtPVksXZUyMeni8QukwhYhoZK32d01jjfzaI
7OEoi3puyCZXRyRZPnGrCA2twtVHdzaoCjCd3TMBwPZeaaZclzwMvC7mg7yUgC0S
6TeUzQfePHhdQLobE3DY8cN59V6ksoF5Ufg67TS78F5DXnmJHMyK2hygiWLmHg9O
Snlj5LPjmbRqA39az1N8AEMyFNv0nk2Emx4w8/u0r1Ho8lYacObMUZC056eWaFVK
onPF/JQ9t7CcXCmTo0htjaLTtrHUsoXYeP82ikkdy2XFclVks4rU1nHJqOxFGp6p
cUJ25s3PxF9NwZdXe6M+voKZCIl/39DMQiZL3xVHz0xIqK692RgAM1jlw/UBxpF5
yk5d+aiXcq4NDx1BqqIPNqJKz1TjrPY7km0oPbmUd4AeL0dlF/Kj5cIp/TuNs0KB
53rlr3dND8gcwlft2mojh01DN0xThxrIBf0jZRLip3nBTLDfVIIuEkGaMcWrFfvs
HhuIyWoLBBFMCZ9LYqmTzDnRcEiyj6ru9GgbrH8ZYLK3aILCy8yqH4mS0pKvnPZ7
rw6X835hEbO2gx+3Bn15tnv3O+InRflettZrudCdPnVsXAGGAPrTkjMGEdpvUseu
6TLrf4pTC7THTjyycm9otOngegwn+fh8mSB806F46n3AtL/fUWse+yUo1TvN8ayu
7yNnNzBqXQC6QbPpPWrMMuP59frBbOdw4zadnwMgWfgwF/kpE8VpYCFWg4KK2LHd
dHUkTewvcjYqW7A4d22bnB6aRnPFMH78sLZ8Eu9tzezOUoqKEQZL4kT6kYSWOG0G
BUb8i5rzEyHnDid9V201FxPNRzOd6C4l7yG3waHw4g85fpo4Um9pzAGL2oS+ALWZ
KEyBnKA22P14Ysbxz6N9jqZ9QmxqRSRBKLGrnbfVjMLmbYm0LJutuyYWV+3q8gwK
Nf/h6Uv+bDDHq9MivrlJlbG+zAbI9/rOYgk05VxklBCt1HP1f2IORKl0NRllvwq2
KioScfg8rT8xtI6KCR89+6zckGYfgFuSf6b306+vuzb2flsz0nCtSrYVqIU8YBiD
P2LIoPjpTsZY1pCfEP+T7dRvf4GQ+qfsAv+EZsN5aXqh97cZLvLpW1FJhsA5RmJd
zUXAIVqS6RodD8yfdr5dxrNGzSRxICBaBnzY+bswCYCCyBnLbgnjStAYhCnWZ3ZI
CvWI1qeJlOky4HKV9wEvRm5sMkbMitRTroSJce/xigS4GTZspR1F+5zCqu16DwBt
rpNCwZeGLUW6fwRJp4PST7VRCg6JzF/OM+H8rCLmtD25THbLLw0pavwtmaRCdjDA
Bm5FcmkduGSuzW+Yvl3bY+aMOd9rWRgP9WhIJGAnMjSJyipk/GFZWB8NvmvQXZsV
tcKNwy3hORnqiChZ8sViy3BAPVmmAyDry4rZDBRM0ZsJwtNfO3qQs8BvvAD1SMIf
IdhFJpDoQjhAS6MmXb/m8HIprDU5lqjtO3zyGlzTS0ZfUAGNlaepJBQK/HsNpjMm
ULIdfIXBgwEWYJgEXFFUF0jLGJyl7lc/3dgIL+SdvI9cvQLA5Ooo81AtMJhJVmJN
1r4Fe7dgWM0o39xZCZVRk5j13KL+ShFbHLy/zX6efYMgtjyEKNNrRms+kSDLS6ho
ihApFyOwClZmgIXloyCfr0HDmUSOnC5eU7FMtARiCKvLTVIMnBhW40m7DPNTGqhn
4d5Wqj/XtLTK2wpy+fGMNznlwj6b9vtHsc8PCBq3GxU6rhEMwKa1IrzaYR9Qf3m3
FzPYzE7v6Xtkt7G8dGHr4rSSUKANXEWRJZUilVnhIFLKzr7cAbQB7N4hvvYL32d1
H0boETCgdwxxUKqH/RvOQZ2PaaVz4X21FuniFVdlVJ//iXlKxyAQ57Tob4HCEtAA
m8CZBK6zBMnRym6zR+JT+d1LumurjmiKNhL5U2X8DJkkpxQx9eCLwZ4VlQoGAENN
Blecx2BTUTrF4burJEO+/fQn1KXSKRoKXNx+vmXgYRFLZ6Wn2p6l4zdKDCqaiDfK
X8D9DHN5SlILp0hUNbSrUHx+Q+3PRFNT0ZkXv8Z0AV+5Tw+DYMPYyV1dQ7eJNRFi
BN8Sh8jvtOt+cxGCU7V6JFKjT4FysmBmzsndxJaRvD4Wa0EC0itHchG6Rie7L63O
pi8/YCfv/5mZdLFSMEZ3c23D50bOLfoeg1pnFXoTL8nm/El9QdPJren8Rv5uD4ka
N7xo7isqKumKvd9RvN54R+cv6NHmU9k+sfttu4DgX9+UmHWoUG1ZcGurgdIMU3QH
vjNlgF5ci80ZD37wn9E5gZyVyRdkbeDA3QnabmjDLthtR0/q7j867SUyD7aNNblk
0GbkX+Dhx1PMg9mo+SlMKxGu4QMQK36Sp6sc08RWcdn/df+GLuXQ3F4R61Dq4ZoK
Bof/yKDWcJzgwi11k2blmWGoq2XfRKf1YNjbOeyAfRQpcUpohi8Ac098H8YhRcIY
ZMucgfh13wIBBxs4zZn/00CDom4Q/UXiPykWDb65P/SPDahYkx9mCc30KL2qBNcG
CbBmMCRc5jJNd2vGnhKMX99DkOMexCMfXjRlxAtYPVMWStZbmOH7QuE0d1dtT6XQ
qMh0tVxJHvBgsDuRLLHZ2wtwuwlIKGoFSG0AGBp/8+x/AqkMz4YEDoFQFNshu2+2
psAIMZp6BJtbWblViE970ySl8Lv9lfd229j+t7rZEPAoNO1Hli1cOA3/MxjZ0yrS
yDltPxeQVALQT1F8uVZ+sLHAxOvfBhQJiLBihAVsOrYGLYGA80FjarpRCLtlZHSZ
eyVXF6CEcjSNtqom1VepkL0D+cuBY4EnO6zrccUYW0XS26HapcX39l2FBauDLCZG
CHyhCmYCBI/uiCgBcmUR+Nb4+b/+p0ARsXGjzNjQYSD1CO67sQedhJBW0/S6x8lV
wOeP8xFwLg99/NBLxLQ48PiZAxCStjWSBI4YGzP7mHPi1crwJjOGCYxs7Mvm2FVj
v51VQmXO1w/yj0A6chBoocIjzM2V88pcqBSUdsjI0y3+kTd1Q4cJWfNNjND8Ui9E
I0hLlqtxA3/f2k4K86pc4lPi8seXNUAbKFa3Ig7OnVVFdhrUtkg6tSXktUPQWrU+
ZDJAQ8FvyiHMcVrBTzY6os3Kjyzav7go8xLT4vXZYgqqa0Fb1hMFdntnlVv8VM3/
SFMpUVrfnTkjrCGpjECHeTbAuD/q53UPLT0Xj0SXVC0gkjaFLskFeGvt0Jtk8LFT
51mmIqr4md7SLOn6ILUcpwiVgzeSLlhS2wAlXFdHPKbKUyTAdRYm95wasxzSfZpc
+v8kRrlYxn9ghrmgn3I8hZNOJ1SrSiozVY4RXnbJRIALb28QtJuhuuUsTSzUd13y
/uxhVrebi2AxRIMQ/iU/NLkrAEhx+D9iVCSoWJ+dfLGIwARax/R7l128+U7IjVi3
YI/EViTqcGAIKyRrzMUx4gby/odtqSEaq+2tHfanXPvhIthblUBsoFnYdYzKyDeu
volFHrc/PTLrcHgmvBR0VGUyLEMVIGAT33cJDyQMKmDIeiXt20uV7uuQsXS8bQmp
P3Kz47Q2xl/+gejbRdB/qB83j9QwQeToI6kIcyV3LrKEi2/Js/DKEur9Vb+nkQIG
zfQfqSSfjxU+qJloDtsZPfvDj0SFazjHZy8V3CbhjhEjwuEhaurpPP5pixwYY4N/
mhNAii5EjLocTFewkYfCc01DyIL5ZEdxy+KKlqQ9ssRKhFUVxlsuRtHjVtUbFRlA
L9QJ8VBMSlo8gPIQoaDxeSLDURHfN1jD2MQNL7fdTjEquFwpEX0EknlSq2Brn7hJ
ZtHkvb2o38L7E0EWuqvP2TaPKR4/PzpHNHlRUJNg59/keUBEYrlEwa17V9m3ceh6
GZWa/V7iXJqhBh8hplsrKWsSbFT8yvL+91pZ46wTz3gnTZG99mBiq5uwYE2NwLGO
oIsotPF1WdWnEw56r+qgxUWj+5eXvMNvsZliAQo+akn7KKnglKbYWDhO5hIiyOrz
+ICeloGxdOvlDXah18ugrygy3sYTE6w4SzFyXjFUKiNjemVQxTPopHddNhXvFJkh
qcolov88CwJWt/fsB5nMvEs/GiM03NdxBm+s3rmtd7y381RSs8H6mewXQ6OFxTqC
nEMET2l850CX1iZAOHMID206qK5MPreOklsbE5QCc2FldUYMKWB9+Pij+kMwtf7+
fPNkp4YRFNPQQGiWVDAStZ659v7plgtJ4mwHs1ircqh+A9zXmDPSSjWGx6mtvBSn
IyvsZmdeqpBC7n32+ol0sC1AM3shcU3H+xA5I1Lq93sRyUa0RTWZjMv5pmaTQkaG
541XgEiEPzvviKYgzxmPOUGb7tmeqxwXj6NztXDD5DTy+B7cTRmrc11yG3CSg3Hh
VPQYHHmpnZIl4vgELVmFngSSuw3wgTXtmmsRkTSyxiT/rpNvpLmX8UV0gmeqUzwW
WicJ7hIzzLw0fSZrvtHSq6TLF7VIHcbTcrdm0Af4mV6pBhdBmIKRvW4FaKBc3hgS
i3BwBn3ZoQ0Qchy+xwi6D4wgOhJ6P6ckE6oMOX+Z86MZNu5w+wQCZQDNoPq60PSq
OdJmw6OSlLtEGgDcyHz28EZUSu0UvTH6ES+nlLTa0paoE2KyDdn/pNDlmXltF8zn
6S1YGo+ED4bJPYyw1iLg8nYkhl4er5c//8w2BpVnIAIGOmwiJ9wo3c278Ltj2hfe
hPKNI6CbjlDVqbNthjpDFGU6Zeu/P1A8H2o03d7DFYtRO+ynvNdONfriqJGrA5ds
U9H15/6PFxYKAIXEsL8/oJaMfMkCeRuWqpK8ph2fJA5yTk+05g3/Kvbph1aJXaYn
x35CTXdy3WzDbT2HD6oPE/+viA02yhpSbmJs2dSG3ExSXPV8reMu3Tg0Z3/yM5Fv
jT96PEuioaB9QAOyns5dId8N3Yjej60VFAbBcZrMjy7k7lYQeTZj8Nx/PyIbLA4t
eSJgalBK8j9mI7HKDl8UaXWp1rpr0R7FCqm6Ef1u0XziDis+osFnTOzkLJODoeZA
oldY3fjBPg92eHn+6HWUwE9KiaFEV3NSyA7SAVjMjO2EDMfGuWGbWfecvxcQ/smF
ZWPOWpaPCa5I/EIZusi8FewPZvvCpv2MXXkTOOkLAw0L6HLoeKit80gn3wDjQRN6
TH3OjCfQjRurKIUjZyGXTbI4GL9fHGoIDzYXZWZ+LKlFEAKTF2PEB2fv95YmIxSy
SkaEfeA53A2HGu+ohViIR0jXTKBnQejnB1gu4iuP8paNgn8XhojRIm4SQ57Z0CI3
KkE8F2Am5uDSxCAVDcT0rsST0e4iobTQtPKpnbf+MZhbolcUtsSNMtO6tlelv86b
jmZAxptpGP2ZLA4jJ1tv2OSgpWSvUhGdqGobee6zobnJKckCi5lrTGFMBArF0VlW
UzY8MFReexXbyJcOElU/AXwIgcQJHTVczwdYTKWjXGF7ZpoL+O0gHf7HxOcdgrzn
9HuHcSbWmSFZBnfww6OOaq+qAbriMeR7j9EMXnMI0HHf8Lzb45RxR8Fy6Bnkr2er
t2llgv2SRGOdJuKdBXGQPj03HcdO6l6TAf5AlKB8AtFwcIGuBiEQTJ6dxcsMouqL
IGTBDDHP0Ulb0SN0NtCLZbcUBZfvGvD3M+0roHgPTQ7RIAAgj6FC+VobgRhmk0b4
aFTIbvn5oZMATog5RmJR7EMIFNR3z4Vctyvhn8FEYQxJShBZpzQ6NmuiYIwJWB44
3rgRm7Liw33SODelFjQxWLzu9+dv80LdpnKEVsHC1zE3rExElJCaC6Zgxo3kUvqo
r5sTArwFMFSdkoqGIEqtujmP1ME9a+LD8RqxgvnppxLNyyRZcHWZOACPdPYdU0sW
z4mH8Tfz9PBlbMjV5EgAPWnIANXjHWH0X4W9llj2ShqeL+4cYmt/zscNfBK9ZrVq
9VDGdrlDnzUKNoVyH9CvszIFRGXTppPIrLAH6y48gPubzR7r7D2qMBGXJLlFGrQz
aW1IsFL7/Z+RxIk8QvgKMo0ZZ+mvEXEPIZSjh6xnC0lbaSogaLxOUbxtUGFnlK8U
GCVvq2ejRs1u7+/MzB/WpAHjMjgB1oE1AKKwPCfX1Q5WYqKcTFkXXoVIUBkZB5Sl
n5vfDE5EDQBu6EyNmiNWNQJc1rbGB76kSO1GoNDhmnIgrCB5LPcOnZ81EDJQkade
1k8LjeLcgGA86Kdk2FCJF+BfZBWR1+9gbpWffQ+nq0gboacJbo5vVKyHu38PntKL
E7nT7lGSw9SE6KfmVxq5pLpXq6UdLSN109TbtN1jVqvIp9j89hhZqn+sUMwArGKu
UtzI8fOvlmcK9sIwkBkfKpMBcPw0y9AJuKmAmevnRd4AyId+xXZG2yp1YgGBB1Tu
z18ldnggiNYAFHMbGwLvC8UR9x8PRVRB+qXhbTVsh/CP7H3CGoL7TiXNM5wjIFnE
wpe8imUtgjyJutvCXG3KG5ryX0KCdeLi97yoON8uGXSwzHFySYP1FSdAoiBspy7e
U4mEGCZCZ9ZlAjUoOrlK1F2UZ/OQSHzCjeuGj8E3UPd9/sncs0pbPOymAbGGZGGR
vIgfYIdYG2fTZYaiD3F2ER63iJru6e6n1NiFelXD3NTkT3o4eqGp4WSI/nE1WpNY
vc3oFjm4vxyFXI7H8E6FeurNPuL14TWCR3ix4NrJyvFrUBLzg0s/xEXAu1dQznRt
28gDZDWw9bjaam6oAKuCos5R2yXYt8z7jf4YZ7yN0z4M3bMeHtDgWDLAK5W4qAdX
o92t1SscgFJReL/slLKePCwzZbtbRvysx0saxcUL33l23Rn25r0wmQjmAQW6Snzz
SEBb7Hw1TiAiRkvSAlmhlLnpLz04LIBpJ/Joz1gy5FH+XRArisiZ1+wA3Aly8329
Um+BgosDC8uUzV5RBpbY75NenGtm0adwihQELLp00sddM8CKJEFcVnAbdXWYAfMZ
uJdgqKpJMQZSYFr67IyPQ6MjyHpVyCdLuI7tbSAkj9GuLW8iQfJ5auIAsubdTdK0
qgPDDdZt/yJClXl/TeZMMc92rsHaH2elxQwVS6yWSvPnctE8b3l4grCJSB62iVkD
tcL22R8BZfxBum3/csCa4YbR46Dx4lKiDjqlZBtuCh9A+61RTRGZzAVueibsbVqn
fYiM0qCLZaZzN4bMkzGLhAlFjeVsV1H0CZD8bXcX2d7ruckUm2udQeApZ6f8UnYF
KQig0Opg0N+9Bb/yGJzT7I1AS3XCgM5LaAUhtV0uJJC8NkkE1L60OJ7r3xBFJfyh
DQ8EXENcUlYNH+wOoAuGP+/JkgYwjJZaARaLI/nEhwT5D2c3ORwW1MeD5NiVrwKC
9SHTJbUMU+HpaNp6j9Sw6G0FwaJbSoIyEN2FWUYVEYlms86rjH12cHY8/oaz21lO
MoXqu013BRPWroWjhUtXW0er6sIhDr1PX1W8CVdd2wuDxK6M0IFxLBJy6f6WJtfg
AdAq1CiekOmMkHBo+Q8sq2J8gqliv9NavdVmt0ua2atM0d+rxJKOiIT9jMHQKvpz
9P84/xtV5DdNJepWqBRymils5zfBNWL//vexYWEwVThA9uJ3an3L3xVARyTiGwjH
MhGa7L4mboNzQMOkXKBCyNSrwk4i7ROiQDMSjd8PLyZlsfoXkZe81QyiXKfEpoJx
m76biXM/NfV3+pGLr7ROSzgl7Iv/WZg6tYUccthwhMJ9E6wvPqqxwb5E3xYBOByZ
pV0rHQzqmK2hLgAneI4tvlIp8ROrI6N7yQUcgA+rA4rd/555esIqfbohXypwME3D
cSS4fdJ1OybF/JDE73uYImB7ycfGIoCbN4DxpQ5NSW5UrWkXiqd8zB80Hw9mIofD
TfeZTTIcqG/P4DrJInyx89oQ66l+AC7TfdZX3h98o2rmur6oKnz+lQAIM8RB8H0v
EaZr8l+eX5zqUtUFsKHOPxIa2+czLE5vyq2Ue3Voth62IrXOG/DwtAGphYge+Pq1
hNWhAzp+e/WdknkSGCI2hCTnXhWi9jxVZt/VuRW0Q2B6vVt9B2uCl4aQ2lEvSuuK
97htx9lQ2PGuEqfK5P3sfnzPbWL8wxAEzTq+6Y70ePIYQMuCISYpE7JvrCYlpXQH
ISqaVROMVslTQtjf1KABAVXA6GrS4FrU8SgF7r7pMp4i/+QFyubB2HmjlYMY9lvD
pG/Q0Oo2j9ds98yQxmHcJbsQis/1xvQZooQ3y1IE5K2ZkbVX6SO1Ja0sdaYvGUmB
A0vA1pOLBGGwX4JzhTNgOorlvPkenB05VqviKGSFjo9easJUDzBv4n7OZkWEZ/lO
44dL3RNYoC4TLvRt48uVxWv6XeypIKN1KDnVrK7CHp4LdtOEx6HSDqdUU9b5xa78
PJXX9IK5hQg7wI/gjY+/FrfyOBsEDrEA95vmPNsuNbcouDJ44mEraLbQQUdqPVJz
/pBVEsbjgJANZ2wnO4mlfLzgyjsUvoXNhjm/YP1BSspTMhe0mnC9wBgPOT23DTvP
Ut5iBGa3HaPmVWQhZWlW1nfub0tNeYZdfz19gXqZ6Hh9IdIlx7ttcVSwpvubk/p2
m5PeKjM6KSGPbqQfO1+GaHNm1hdxLrP8sQ08ySRQvKSgDH55CuJXBaB8dxUpJfQv
QAQZmhSo34I0LlrmDVB/wuBHeePfLafy2lRvEraHsmjgOxDfEr27Q4mD3BoVZxf6
9SC6w/g8DTbsY+BZ4fCbDkDo02qTqKFEw7ee/LSkPBcQh1x16WF5s5yA2LQaF5B3
dX30fFX97i6xNzJijklq33wCnyLOq0s2M5MMrU+5D0i7Vcwk/0d/Fs9wY6lYUeTg
eJ7fF+kli2InZK2lqZUW8pNKsM6G9kS9l+c5TImTX7YviZa3fUKQU7G6IjNYOXNq
4ArJBG65J3I9LdoD3SBkEH/7+U2EFamswsYQzBa5y4QBpKeCYMpJNwy7AuhVqRpE
4og92cj4CmZxe2raRSasdRG8ibIsfQUTAdZbB8wjHh3iM4hz9/3LnBGsv89y5JhK
B5jQigFKmZWffUWahzFdyOlS25tBf+RnfqcG+/6mBiJliylK3iPp0+MyleRQmMkh
NWDuSbat7frDQxLw5f0Rnuhp8eqw1rXxClpIPxJPHhErufH11gqIHXj3Wg4r2QiO
0F/dMcC4eRW3nQ0uiTI41i4akqo/KpBABmFtWb+uMg0CMWCUMYo5Xid4sFyNNudT
aL5Gr2QdFVVb2cabFTzOmkIbOdTHVQ6SEE3PS/0UtDQYHto3bHy7cpl+i/pvoGBQ
lJQBzs6+IFC/ZMLXifNdl8QGLC2ODcoy32rb3Y+27JkzL6dUbaI+Xh7B9pQaUnpt
aSqRXkGhimUsrUYlx3Twl5HMYZkJBOWRjLK3lNXa5L67A9Ps/GVKBE1Ubls2ddc8
WGC3HZib39aG0KDnxn5xuEpV6pe0TP9YvinjDR+/7Fp5yl1+pejPntLMj/YzJtxA
gGdUbqWFnx+JKbLamYQ7rXauwF0BVgyCzk5h3jL4k5nUoG4NqHzrMEFhiPfxhGFT
mtxWzwmcQA+cqocP1peDMNkWR5PV3cn5vqbmUGnGT2KMo+hIrarrwPbZAmzUtiA8
sXEoNWrtDAFumVDYk+W5dKgEt1Dvno6Z51/+GZXbYhJfdS3YeVVrJ9sI1jFYNuKj
pllz9SAhJT+YRh/l2H09Cfi+4zBJRwzaCrOTc213a2BJlx/qyGdHiScs8lPZbuj2
QKxKdR2ND9YmLucIdIHm9BL7F3YD9Wq4h6fQpqyJjqdsw2RyTbGpg6AXR0BGwyFJ
Kg14+DIJpv/CMkC2dFj3g1qcCBpg8D4VHfXAs+dq6lKpCs0PMuVZC4EkRd8gs2ka
7iEr+SvntjxK1ZXY8id57tygt4usegAqkieJzd6Hm/yRhCh4WdkALsGroCqsZuE1
IXd+LHj/mkMejWLxG8/BaGzxLbM86vHZouOFze+gVh7YC9EdpOSgw+ZeP3zyOTSV
MAvZKNtSqkQWi07UFH2VWhjxYfEOvlZe1J6IB9/OAzFIuebryg1ND+ROpzOS4b9W
vk2+ybWE0L5/Y3f7zmnYBAXrR2zEGCu0vmFaOUVixcHRPY8hSCmJtoAaX/in+vdW
PcGaDqTOjXmg5vbtlprLIsQqnnNs1+HcDv47zjTeRgDmHijkFqScc85VBYWTwq3c
NlTMKMOZiMS9CBRmk8klas3a9DEAsVsI82XRLA6omhB7qcx5EfjKQFMkdBP/BNgh
g0t6F2KxxAcUX7UZLXpm148c7Cv1nhlU890WnCrId0F/F4AYxcJKGdDcwpV8V9am
VEE8tqdzjSHyqXjRIx3JdkG8MIZECzCsUYCRxk8m1rTvIFQ4yDubcIdyb/fjKFs2
hQvp1j22k59xoaMFj/MNvQ28eJGGj7mBmPXcWORsH/T5iyk0AitPYZ+9vt/y56eE
vtqGWzk4Ou2USJhXYj0DZeT2F3CFZ4BM7gowEPumrpqck8AVeITEAHnmX8OSMK+E
d4q+7rBQiXNGD4HBnc1EEyYoJOS+BhVibT+9pl1OJ0OuxkliLAxp7rhGXQ+QDMSY
YVPjmvWVCbDLcBLDCBgIKaYbCHkY/DzFq+JHYcW7JpzOcPr4vtkPI1lkRa1h4zmx
aAD9VJSESS8rGRjhpAQa773FoDn58+UOcEM3dOz+cMevLuy7ywCDPWRqqczX08ch
HLes580kYqgUT3qm4qNPgTShuiCA5tlmRYDambejCq4MkQjIwxfnO2TzueOqnSdj
OnuBSwBjhUT70uwLPoAEzCUKDyRgRi9p+wK1LXLa68J14X6ZVkxN4x05DGrNY4C0
g8klaShb+fnUcknu9o/6YFhHOxK1+XavSsQAc2Vgc/2/MxHu+OLXIsiiw1ngLcjC
hq4nTxNMVjAe1+t30upFK8+G9mo0vdJPviCu/HtOU7jpeFpSUHGrvRfx+7jfeTdN
qDybjpdVgLf+0dtbkibuH1OjJdS8ci2JnDlIyzHYIYPJwkd66NiDq06WCGG7tUvr
DAR4j28eQUCrZC7Cpg4SX8t5fSMpAFk5b5X3buKbij/DPxUMCqv0KQNY4QzGQv7T
AeFo6ibbpvakfdNwkgUa9xhceoQE18pOjkPznq+q2uIxjK7xt1LzI0QD6AoWZEst
6DFG8HwQWcW6AstS7zUD+iXR1rRwpF/8qkxR65G+sRRiIMnHa1PkG5OYofUwMCZP
h3l6fwIuqCWshfhRiAt4ri/u6xQJrPMW8s+akbdhi0jXUp/PetlMcFwcsmdKsqBu
ZTrrv6tVTuKEnELWPlvvTE6lda7a57KmJHXL5OACRBpeEmTmvKhrgjjEoLHyu0Lh
+Yto8jXvhJrMDLSZiLsxflE6plyahn1Z3XawUlqD8WwXzwxhbs5SHXQtHPD9lgpL
JZfMoBiUZqqiFm/SBGhjv/hpgo8aejN/fFNbA0nK/VL8iIFo5B1fFhVQfF2NSMyv
wh6s8gWZ3ghF2sUH72jjeSw+yKVSSySRDug2r8gbRB5c00QVuOs8o7YLvH422HQe
ieWDjEs/kNc/7LpfjzagiC9WNpYRlHGQRlYl0GcMs2zpn1nNjYQmNsi3Bvun2fGj
Yc1q2ZuYR6C5ldCcSGSaIjdFWHI2rPXDkpWRh0SfL6HdQExQ6zrNPm4xna9S9AlE
1LZEoFaY6hCjoe+2YBG3QgdjJGqEdGYpkXWpto5FKLtryvu8taNYU2tqYHGT60fC
EgFQVvLKg6tADcbmBgxkyhfMdmNF1/tdXh68CVGsV8XZsohBwt3/U1tQxcgc947P
mu3LjYqdqlONQli5gq6eJDELTVmCLRO5sfN+ytjf+nGAhr0BbwphmNKXBJjgyFxF
HWS0BVvJXUeqtX4HS6eLibbEGKeaOpIm9WuYE7XkRcjv/1Evf0d8kXVRzJQgY9+b
u+b146MSMPN08UCpTvntHT2WPnEfjruWoOEdC0//FmJydut62/6rcjbil6eb+LhB
Ri5DPxkIMcK8Ctu2YoYNRapLgncUP6yOkv2cYUW5baNdwal6+JoOS1iKgKMVUPCt
EtR6793Kmd1GdQ7i51CUbiT3RxJshuipKzrLklh8ODmhgVxzrbvLhG7ZNA8lYLyZ
GOrpKXpgdu8sQxIk29rDQZMFpXWTyPMFDL90tYMBA2p6QEaMUIHGszSKVrGmXlzz
pn7vHe76eP6lOz4Yt76O9nRHJkl639/U2e9CEWg0jVldHqbTfz4NjCJPGzl3YInS
KF8oTLSarcNWdtol7caTfywQcZlGXPLhucGxaj3LVS62ZZVOG8qJkf/JGATrck7k
OKj+G0vxPsg3D7kMb2rMlRQLKYpDwGTnhjxO2HcDYQpfUnohWeZOqdE7A90vpDct
vNGl5wQe4ySv+6R4d/bRPYtnEiuQNqA0hBQVhiWHJW1ItoF9657CbSUKPr6CE75e
GZlNc+3Ubmoal7UFTAPGEbdYdVOhAcPimlvgX7Yt+O1020+XyxOMpwG6qnL71Aa/
DB9M+E1ca/6ZKoLffvAcY9i9KHZ4JC0BQibyVvbnuHWPQIxiko10mKYecIDJr3NJ
ZiRtvQQMgwQzz44XguGHUoqC17dEU5qIMgcZ5jBG5lG9SL4tWyVW+6zyds+Szdza
rMTp21ZeF4ygO+MGg2JD0kD4kSx3JoH3CWCGRIEbbnGcjUAyJalUKBp1SHA1pa6i
UCJAKLXQaPBYJq27nPBbiZTlRmSyFPzEjJYwXlfeDDyt4rT6bQRFNRQZ5qcJjiKq
NI6p3s8DOQgnBhr9D9elOVUW4lBEEqdPxc2WOyTsjJJimEMjET9PiQtpXx+L/RDO
Vv43B6e0Jn+pExSAxwkrHuujnZ494YcNZldT62nj5VaaF0MAfsWY0XY7r0rTF/HD
/NZesNiCBEHV6MXfr8kXtAFYR/pM912Cw4S7t1ygLUTcZmstVjw8uQac/w/6gUgp
UU60wUNk6CGv7aA+5KojThaheqgM3VYHwR562EeaI7uKvCCRsJzVPMV7Q6Ro/IFU
62+nHMUux5U784gKHNd1wKCDQ0TljhxqT/m9z+tW59VY51BT9yyHkQ6YQYpZjdCm
VvxGrNR9USo9R9wzLOESsoprj7EPwI9Lf13oo9HWfAGkzMFnl4YBzJSwi6Vk3nUE
b3ezsVLWz18kzER1u9X/giZ/J3+TPM061CsYnMC541jf/9N1ocgGUYUn1J9IMogL
ARAAg+ojRO0F4SAgCOaD1eqPzPDJq/itPtpKMr8n86PkIQYH+l0Jg1TnGJ3il8H6
rAfub0hJBNA6E2zyeAhcuTf4x16qmsCeHN5RKpJUYRXpSKb0L+fI7RJTt/80eNSA
TTvN1dKuKtEOUj+74eGQSigx1b3UHBqppmbpLmbA/TOVXm7eli5b1lw+LNo0gzP9
Ly+QEuRNmPhZWRQlTI8EkWjIGyqdYW08wSl9PtZbMoD225YJbXdWAUQtldj286Jf
zSYoRU1mMlmKkd0l/nSNmTwna7mHcd8rnhBjjejqxhY0yn35tMXQ4zDA4NIu7VCV
Yx3dsXR7ivLZoGUvWG+Ot+zx3As49zKDFoo0tumqMJe6v/2MwrA9JiNhCD1TG7+J
+APOvzpzCuOzE7gPEZPHu4chQZ3KXOsrObqTkzVmPhcEgcVlmDV2uHCl4CrkVBkT
/yaK9BZ8AL+ulvQZvlCOXx5jYcIuLTr0jjgQFLGmZohM+S4tU1WDW9M18lnQuJ4m
M2L+BcMDGkknEjiuCEDKOKqeie5lb/8PWx38mlmkSaGU+JsUwTvWXYaqHCiTYAIC
5ll9u1hpOXjZrN+Dxk5UxtaqwG/OD7cEVQ1e7Ic8oEwYTBd55kGeoen+Bj+6bLQZ
q1hmxMvPg/qFA3pi6RQp+6AWVSBXA10P5YX7c8z+Fc65O12WwL2ZnauYw98bnRyN
1biqPWyD0MBGArGq02Es/g0ERDOtixE5jU0ieCJTvz/6APPa5Pyt1EYgkPNsxLCV
QlJUbECVglYNci6MPYpx3qg/OkQ221qiEioT6Whu1OC10WCsQqurNHq8K4fBRCB0
hvL+r6fudWKEWQbMlkP0DL1FsEge38bKeB1ldEzsTegfEgFfY61wYL22lyXJsWoy
1qGaCeCINrpu081ApZd2sDTNs1etLa+4W2cfGX0GlqZgkJIKyG9912Cfrd9H/Vbc
+4RxgTgk6C7exci3WjFeEx5vEusdK7XxAq4hA4sMtWwvRm05kxnw/3JgM1qINokx
g1uNBcziR3N5qyJ83TEvZydVuM1J3/IDbF4/gyXk+GUwNTUNR8AFrvRziTV4zT88
ugZML9/WPa3HnBB4IbCX2gGF97jzG7EX4d/SX/1Uav432tLfgOjx7bkomW/oj86I
kETYRz3gNa7nS1miuTr1UDF24m45Mn4RxmTfTaSn4QSqfzlZJ+DyS62K8cEZX87V
iTWpuIRZ6rDbE6lu4NL3wEAkIWla9VTrgQHJev5joUUEH8F561RPFzXr7kkxXRcy
cMx4UFC5oSGCCucRQNpu3bwqVLcR5UXSjaex5OjhAvxJL8/IH4E3pjBJlbi81Skv
G0vFpB3k5tWqALDNq57pPoenZFsxqG0ufIHGhIrJ1R+/8uruCtLiKbXN2G6SAmTh
DvxlKlPH9gjtuSoBV2T/OudJ466rMKvh17p+VDJUsbqtGYfCgCxOns5QU5XdwHkF
IYJz/21cVuCZV/qDtKGUzrojzlDN2qn4UkvGbOcIoyek+J5tYu0KEArMmh/7zDI4
gJHwH/2fRlEC5HXB8if9ZOoo2OREmXcWvqyxvwj0Eo/SqnCee3UZvJkZV4CkVaIN
5QeoeK2rFn0f8p8lqJCe2ED/1PwfPFOniRVNjWQM2K9riczuEK9aRgbXoctyLtAy
8XRSNocksM41lDTLPNjkqxtJfdrone2qaNDXgoy3tlUUD5xARe49vNw91HcEdERp
cDLFyzyAC/WtRhIWILRiBEUVX8BaKD9lx4/8xNm7tr7gO5VlaytZscvdOAObg01I
7bGY9qkfyopsHLxx5H0cOCTX0ht/iCGMO3S3oVBNzjnDO/kcMbpAKnqo2i1NjACe
S1t1oxYMve6J8VSbwHBEgLkf+kT1AR0wNQnsgxUgi99Qmr2ChKtOwJqzt3E1gDJG
KORFyDBXnAkhljVNt1z3GX4exnW+zk1C+/xV5UELuKTsi1VSKZ2yIy6bQiMDPwrT
8cuHc1OXK5PFDJjKW8sY8hSlb9n9IGCt3fpO7qU3z+7/b4ZFUe/cgRcoZVFe1LQL
UguFumwD0ZfXqEikmQupudJwnX1zflgmZtfTHYq6bHeXAo9UWXrw904OtC0h6yHL
pIs8Z7+dY24MD5mFrpQIZ30Gz/xh6ObyWOf+q/LP+l8AeuKPL2e0nVCpb2adv6Rk
4FhizU2V/eTsa5CsLrlPEZEg3oKgKpXxLBG2T9Osx/fwUvgn8WrmVvaJnEyVhNih
97RXBqd5vGB4CusiOY1tnnYgj79W3ETo4tFlFVGuadWHi8hgukuS9hFqFjgsL8mB
2LsnDTesnPqkwgok2NokBB0CyI8xFILcEgAgqkaoDHDqIBKtS9kmsAE6yRvP6Wup
bUoUtsLpCvZ/naHWBx3KDMxNXUo8OWtb/3Dw/7OiIE/s9tI0mMsy50Zi9u5uXjP9
kz7jPrNiQlP9M40nRKObL4wNpaSNaO8k9HXM8FYlzXOtcJxJ9zPd0qQ8Iz65whiv
IplGZJB2KR4NTKQk+nt7Rgrx+RCVsW8KK9ItOKkOa6jjCoxQHnh9pLTThEI2Jpk+
R0bcN3sAvqPhJnGiUWHWesC+SyD0JCb6fcm1F8ult4+PWtHS6wH1H2zbtLKtpzvW
+T36vD0LUfKE2vAO9mjX8ZXt6F8fvfhTjHB+Rzb9KzjSbJLsOFYnIORsm0PaI9xU
lYiPa/BG6whdFIbY7ndE3ZnXVhzzZQJcFjFN2HF+RnHgAa771u45B/eIQaxvTp1s
F5I4V0Cj/87PkST5PRNOMR8YrUaNkV7zONKxExab0wOWCs2OMvp3ts5Zc79cBWjp
VFMbqr8JanG6gtAtXCfnB8OElYWSjBvFI1w9xDAA/5U7snTSC5VXlGxV7CN9xSqR
euj5j4/t3wGhoSLKa/fAQPAosVQMwiM0b6CgwaPERfxVdJo8q+KPOiBp0GfHFQx2
7Ez6T8L4LBYNuI6SoD6D/uyICPQ9n57ljvmJCBo4/1wyMOH2elFm2s4T820g8R2x
MOmDfyAC6DgDUcS1SMgKBYHJQbbCgq8xXq6q09BhdZ3CbbCk4kI9+GZCUkLj1g6J
sr4ks4hRBSp+KVjHSxU4ECOI4kvkBHYRS+JvDVSYxaYA+XMqFgKkeOeNVXPVDlWR
CrDXDlXC/iIPMMu+FA+DGSbg7y7AfQ0vIAb8laP6KXb5J9Zl2zfBfqM0ckl3qG7Y
Cm9dsGudH0PFNo2mCgFrBEDSL221BWRWPip4gM2GPbYQfFJ41ot8hYZkf5CCXALT
d8j2TJtJ49Ne63qFcSd+ZC0sFNz3g9KKkeyPm0uwblnz54Vo/rf+Ser9m5snyJQv
kwNnAGkNy9MmYK5wYHrU5DDtotlXeHJDARRBMp9+iYJMyqcV3ckYMHMsOIm31wNY
wugAGNCr+QxHpwym3TXSOWBxTAip2731EV5UAeLPKzx6d8peds6w2wa5JqxzDtwh
T/KeJInoaXlKboUHIei5+L/l+oTUfRNVrVGGKuD5Sb9Y6nywbZtFcTaakuObVZK2
uEgk3tWSsR4e6MBLLjsIdxhX6liFQn84/acxky83GJO2L8M3pqc8BxgCWlrgGKql
e8581n2oKfyC4LNZpp53OgYPuq4yQUp6HQ3OjCK5kJ5YLr4Ed+Q/pDw/phtsI7Gr
APJ87GhkzP9e8GfMjKCLuTby1yOi33oXKoWt+IcioXZqe8XRKjMSQfkytPlZP5VS
+K3Axigl1v3qllp8T5DfxzK0qy/tRzRDcWuEQkl1aDA+TqH1yQg/ddgSu3sX5tT0
YRk+0G9jSsWyJTbFRXiFcuSyjeooKcgGP6qFy9CDmg+g1UfqGQG39MRaoOORJaFl
FZLE76ZZCeg9Lhg5T/txq9RREWXVdcdJ5zHfT8PjZA/JSNIwaYLF7eL+Erl3cie4
G8q4AAqY+cJmDCUNQQEKwB0FcqFJ2qHYlg+6bdsbB/SwU2XzVdekb6kNrFebzjsE
VvVpqp5QyHoOw8Kynuy5pZI3SufU0SDAOEG7evtjQeZAiUeywuITJlSDOtQo1uv0
YvI/OImRmud7Cr9gUwR306FlncSJxn+jpmNdAqbQXljD5Innc0nIhIwTLuuqH8DC
/cU2T/a7b97nAT7Ztq/fmz511FOGvpee+N5IjIvZRJvu4lx7D9le+ua4ViT/bpgk
J7/2SNXcvRh9JsF82baWvBUkm+MWQwlnvRc9zMqAKZXwa/yISITGUC/ximgylL4m
dSL23FZIGgGQ0oNcwNE5zVa2DoPfK8sWoXlTTpZhG2qMXyPN2NLsp/tir+iD6aYW
L98g/ehdVh7JIsmSC1Z/UsAK2FU8pPV0B9teuyvu88xlV2FYfFs+dh8JUH8UUZvf
y3CO0fWHzPO4IOqZ3Y4vViFctd9maysHC6/2U7Lz8eaSQRh3ihbiQ1xHbciSMNE0
iG6uQKATjkdsd+vYCQQpda2O0+vV1gpDNthG685E4s0EIvPQImegSdn2qsleVzrU
Kdp35RjfTReWXaKAHJHMTDj1Iy3C3SuDj3vA/cUoqXpWX8QFl+/MQXFWSeAkRXNi
sSO/34sM7xfsehmXi43ixEJhChMXSbsB6sHw/QMndTM8d1e4spHdMP+Xxphi4hDN
DaH11caVaM7G986tn8Yp6VckCRLfVaGzQeEeD5QLLry6chD5H7siijeqGyXar8qu
+DOohR5kEKsVBprBQoT5tl0vjObwjn+Coabg/9fpFcRjE3QMw27+tUuAv3rzONvD
WcB1s1xa7Zqdn392Vt/Mqlowm/NWi8tAH3qFAzNPDkslFiHFu1O5X3KMezoztjlt
mu9T7bTw9Ee+4Cm3KDIcBVWZ+cQypZuO4CcS8aYgULVDnOQCQJoE5QUUsCX6nnci
5+YxzWRWiijgMu7t/E9mPatbmhodc31pz0zlebI8lGEKat2iq9h0cNhwcv2lSHTR
9TmlUM3waBH600gKC+BqL8jbeb/74yNIeRrET1v6NsLMKR2B5CyC+1frnlLJGJng
XH8TPB/aIf95h5nUm5YaQEFriPUNqEMLQoutdlQ3CJNEczan+iIUH/KxcWTOlhXV
eU8WJ7UYm8IcBmppw+I6QqYt/cl+GKsQOFFaLYruxfLioBNAQePaEk0ml/2xx99O
7oMqGhaBqP5vXm+t0AhTVcGX4rDCZEmVBEuez4bnDDn9XS2PwTx/LNREWjqKAm0v
dM5TczQkKdDwkiJ58Z8a+3kJVmAiiR3cPfojYf6J/00NYXV8WW6KOlhMCPbaKbG7
TN4UNBAVP7XMLHOzfim1/qMClM5fvPcUYJ/+AnQmA+UlsEPSyIoDvaMIECYiAWAg
7Z86X9O7fRMYJcRMsVlaO6XwIXKpen5Phxuu6KcqqORovph4l+giDVy2WaTGWukz
5GwdFSwexqj04iZY2Dxww4iwZUUxHXZBVOZ77Gy5kT28HwvE/UGHnBEQWGVs5v65
RkPxSusQNVa+Vbf6QTTdLDgat5eAfJY7IgEvwXWoVi/NiHlYckMEWkkHENRKs02S
z406u6QUksSMSpGxXYSD5a5szWi1je9qeqOq/oJ0VyoLa212NPmKmGBihquYWZhO
bWbaFFEwebVgKIc4/FQB606SC4CMDNU+JFF6aDNd1ETny0Eywf7cErz8EprTT66D
xMAymRm3uJlRbuT2O+1gx1vnEnhEHPqd6lmaUKYEvINvN3UqCNAd0wSlmMuClo39
pN/kSmgSh64waKwSj4zXK3S/Y1wPWpsMzAWo9B9HtPAeqf8XGEFYRHgOkmXDhF5Y
Pifg58TplKYImFga3WehpqKNKP+UeSjZsEvmys3+fS0kN7cgEH/C8p61BGiwGSKb
9ePATxyprJZBpOIFyaHpJ8GXsox72qmxI1XXQwiOmCga5VdMD8wboNl1jAc/ugy+
Qtk5UliuTai0kRtxKvy4xdlo4anj/cKPag8piurEl1knEniY7NpIbNrWYZmq0Z5l
ppdWF4OaGcv+8tWWkuDOvPqVpLdULOs2/hrTbvoPEsjvgzYtkllQxLcpI93PMbej
luO5ER9EhMfpn5Nq6ECjXtqGznqNXvjYwgZg+nLkWvq5ihkt2DUIxYdvt4SqA1ON
Se4siZr1DMdKdNqFaHv+cofnrDx9yxiaqlW4vc2j4v252ZNISarkOTEZhNhrjhyq
dAti67pi7Wj5lLwz1I4571jQGksWuKxn6wraHMBgOoBO2Jx91HBtQxM/II8NahwE
UhwnKy1M/O09E04yD/AMy4G5fI/VLKf5iEZuuhK8Vxw4MfJ1zUryE4BJzjIJtejR
nFDM6tiE0IbJsmN1ohICFBjPiCus/LBsJJHFuocdkfhzzj7oGEbfLHzTqoMgAkIR
QDCC89OdBBjmYK/fGiWxxtYdhu+MjC7LCRF+D93oendEpizDBLMTcQhShjUX8gVf
4TRT8ildVbuXXPN14U6hGEEOL7EXou6SpTlEp6RhiIywpSTRr1QPQvthR9FL5pMi
8G9zP/Bhj3RWHl8q2w0ZmnUOh68nVoqSZrtaWKi98pBM25Au/JEuSz6OPCARRi+V
1GkK4mrBVsqhvoprkVX7PYER6UWlreJ42Mx8olkDZrh6al4l+IzWropd+UdO80H5
fadPpWmL3ogkhPWPwKgCQsl7krdxUX4UmoBa3J+vNyc59xnLbzdg2ODJKSGp2Mkk
H4eIy2EdjNN/af0lJxIENZ6c5fj3KHC6mtEtdzIMDyTLGdCMDI3jLiLWZc4rdxTs
hgio4VrUQFWnTbFtimdLuUe5Vcw3i0LrqFHMNwUOSmp5DxJPCUWAk1n3tT5dp5oh
Myu0KfBrq2bE623C1fBS0jBJ5XFvP0juD14/T3A8kz+dKNk9aDfnzcR0pBwORM7D
ous+YZzi3/3eVoiYTELqA9lPFkz+cFcymLLj0UsMJaLZlHiOX29gzXVP9SxDlZm9
UuHPRYRA6j/Dtxo1MR6kQUjfWO6g+uBnXjGAHKZQed1yrKmGvfUs1zuqaRNLT72i
gcOUSbsl2EA8R8lXMyqiLAA83z1bddq/an53On6rN2DfDxZp3LGOm9YQBXdvg8g0
oEiMxPmqhxJmORzSggCAHC6fW7WmUTMXMzdS3US+iL2fB7aPVO5+MNJvJ2GBNN9q
whyr1eMyE82wXuY24nRPEuLMxUiROAwg+3OOX6J/ktVbFcAwXOSzkjGv9qt9QXuu
N4yKt5ystRqbUznaY+0NVtY/c4p9NsGh+MwuS9ELGgCID8/qHy1iDrCfB2FARSuT
lgknWWc+I7vDk0Sh1y5RKYQn3bX9B+EMoTn/4QEE30GnbuPXh+8c7EmjoKmhs0tZ
nxBHVxm5oxksMzqOfz2C+hZhMuKUcrS2rOO2GnpKFkFz/onrDfwrCXhkduq/3yiM
dgYlHUwvFC6gw3MYjkFJSp5q8HA/8nJl0h+RsgVtEyzjaaL8JjYfMUHNAGJVOiGl
BJgrmgex8iYC8VkOj713NF58VHK7uBz64RQrK0f0sqpvqT6ALtVOrV+th/E42Ypn
zW+6jPwfscBPDiXbk6Kx8cwX1dBq6f7Am+zGdtDNREHOoffP2u2mDzHFNkzoCvjU
AUlaJxMRGmdUo0CpBW6dIGW4qgIAbCaqqwELJOtup+LM+iAo8Oc8j4c+rSjKKPiu
MesEfZkYAMizRGr0DsYnpioTpLQzsZAccVkBJerdP8SA7C2Ldi6i2uuXIjU2oNtC
Vo4kgkXISREY94+0E0PtT7xHez7bclCeun+pl7gT1a1UZtDR5AYOvLJaRV5qe6m8
WoZDRka3HtLZGSkD580TccsjQYXQ18b2fCts92X+nLN+sbl4MG5eiJO8gr/WlBeV
RVA0++AnxrOgQYqTji621/7sO8fhJb6htdDOwEfB5inh7rw2XOAtGFvM754L4HwH
MLLuD8P9Pal9rLMA+YmmKPnTUIvkqmHcRxckCrkFxYjIcbYcGFShUpKplk1SzXH/
do+7cLaBeAFbubZW8NB5CfSbQI5vKzMICWcUH30ahJlqeJzu217naV2+hVBSoiU2
L9IFaAOCPK4l3FLL/XXq4Qb64mf1NL491QYKknYHgotiYur5TMxmid5DPs51tD7Q
EdtXzC1d1h33wKbL/q3ggfhbdlcsyQTDQCsDU70YoQ4l4GvyNarUyrVYqgy1/QWz
q43v9HxqoWKjnsjJrmadGjIRGNsfrE1iskQyZ4uTvKAtHTHJfvbw++2g+Xu63/lp
tsw8weBinn90WUdyYy19RrnieDcodtcEYj5K6NbewwtHNX8dJ8EYnsya8GQJerf3
tKHjzqVLd6PhOV6kLsINYbrRE+PYmErZO6WfLjqHGSfCETePxP9RceO1dgGKG8dr
IZ7ePn8etw8xrJobRFUyZlXnAn7ruAmS4vuFUBau2hHayj8rC8HSCWa9TsicLlUR
cwtyA4qophiyWuRp/MfPMPuPPV6wlbYjTzmnoh4oVlRWBDEDIxDkB/5G0GnHPL/G
0zkj04q1kFzwAcE2JzKWq8RPaCtb88OXkO/tw9YEljnpgLpmYsUg4CZYc4XZ9xKG
wF2jPn8vBqXHqTADBpO3MyvplCWtTS0Z7rDvVyTGi62KP5lQf3Mt30cE8YHv/0w9
5DqELUeZ5cw0k+qDVpnAsdH1Hqi9VDANeWx+/A79UxuqpnC2Hk+76YC0edFvCSmd
8NhNg7VA74bvx2tE0T4HVPlhVKvJqpDYvRhYLc6FBuriH0ka3TBvp3HnT46eZVtp
KyNnn4MetXuQI18A9CX9RoLMACK+kVyuWbWJ6CRI9Oghu4n9O2RMpnQmdqRgmFT/
w+wHa7yDTRoGr+ab+dKIEA/7N9znshnhUYDgPykOCPJjlUqJWcQYVnLxUIdPPCeT
9DvA8vhZWhNUJr5FisL3vJuj9Z5No3mDxLZR38mprBY/KPZ42wTZYo0U+tuespuK
8S+ofLbzwAKDc/J+pEx9k59LiM7UfJnbXfKV186jUphliqclz0NngDW8pb/k6P0E
z0DeB/mLj8PNwksN2fZZjhBWxEe65DhQt6Wp1sJIu6hnprqiXWnOzwf9NSChgK8s
mVg4SH45JvI1bgmjWb5OyUQZ0mDK+kGUgImMwSAd8uAj5ty7ohecXr0qo0QGpqm8
JJ/ZqMtorp2XXLFTXnUh4gOGOBOrWFyRZD9598/YH+Hq3d5m+YTRkbJPI+8p9uxo
qhjNtVSXLL+pEDCchWR9/AzWYGFo9xkXOchS9yoqCpYjL+H1QjqEE1WTrYT51Oov
oeBulQ+NrsqlF1/tT0MkQYWE+DVxaybwwjeQAW7uRYofKobsfRYOxKj2jE9Lk97s
p5q1PI5twY7amohemFAG5M9vyTgnJdqggSYe0P0DrW6rrtx0v764fyjOVQFrryfd
ichSRN3hKocV9PS9AXQN4a+OqCKcPh5DZqyh9QpK9NDfKXlJnxftn3p0gBzE5XCo
HNKEE//ZXHy2Hi1anJKH0shlX8pjKjEGUU1v6SBscNG6pBSNWPArA0PSrsa0c7eN
VjP+ujG8uLg5RzQvgD5+QmqeELrX41OtwUJ0GPxbYwfqn8rGimcJ3W+576htWvtD
59+9ARzJSi+k4AuLP+TeTLQqAn1ZP0fiB81L+Bgx3PkPQpcDlvdNzym76Ymi4JDV
ICINwItpjt37z7Ne1okmp/rukPamSEQ/COKlJ01IRSMPu9uIng7xsgnse8NFpZY8
bgLEz5TgdrXsxEWJmOAdno6P0/OjqXPD7p/3c6fTyPY6h4Jxw5DEcTkjRO1k5sBt
YUO4GYzsrYHMOdUTw4MZTEXwzVJwIOdJKsoSHeP+SC22YiJON5B+XlPW4TOLOn4m
VTOmCvP0HI7bXh3cmr7d74trqwvCQjpX41z3a14AOUYAbAkQ5CxKdXwqoTZMp3Bt
ClfssBMlAxbMTQ+dbQsMI1W14oQweUj1IUBqVivyzKcY1c4WhfLyBOrtYILcLkeh
AtjSW00vVxmsHE+88AH3LvYB+9WZXlG5g62V2QktyhqC0NpiYifWxtu1HCoVcQLk
a4grKnyU6d5ZsiQAU7fj6eL2VMP9VP1p6sbopCf5z9yPrl+WZOUBqXJb3BSErBEB
AqlwpEovk1ghH5Z0CbNd6Ja7a2hM4s4z7HvLgXTsllQJ+W3odPEOtVCQeeKuvJRi
Cr+d9DwstavzZBXaTACuZnKOhFIbJpKRIPTdfwabnpm3zSzPMsPcAFIAZ1wSWij+
ysHXx1cmOMFhb505PH5kfgQ0eDTWii060+25NTjnFmgI07nBSRb6wcNwgxCdtIi9
i1cGVzUpsLj7K68RgGQvCbER0ejwmqG8EaE94dxWhd5Gj5BBTeOh7jsd/N3Wg67c
9q1HT7kHq3kf2T7MXCTRgFwPEAPefvGNPwgsSHlkUdB2Db2gw5cUAXtyDtUWzXxz
QIJz29yDOEnF1REIYNmfDn+60D2mFoc9BL8bCdMIhyA/YdM+csQiodsVpOhNfcOE
i8+Hi6UgYXJkRNEQE7Ith5QPhFS9QPRwElQHZJZSWJ2KL4Y5J88pcqakndyNyUsx
soYo5mPdyQnJd1knyy22frcpumsp6XMgjKqXsE5f139YLgbs0xQOLYArVJFQfVp9
2/9nJSdkEUr1MN1Aq4Ux/eCWDawLEnsEvLSF3hHx2vBZwKf1xMb9kgn5W9r4Q0zf
0g7ygpHpNUAmuOPJwyuuCHHCIQ0FK0yRr/dIenj9vFMX176vt6TdGNo6UIV6lLJS
F7IRYJyub7m6aygI0998pScNeNwCkFVN1QdhEK20UV5xwAHk51A4dtHFCr8uSmxU
tpEKVo2TaqbH08+uX7cundSt42rSXOcvMCJr/OHuPYMEB8+hoZWDtQRWj5rJNtZb
2L6+rf6MgmW0D83tJwwNlkAUsRiPDja1QekWTx7stMk0ri1JIxl09ow+n7tmfvHD
l0LrFEi+IEvqNLFM55XQhtRSugkb9KZ3SP1cfWnqs0i9cH2HeGdcar+bM+Ue00RF
lu7pHde+3FlTJ6Ng+qG1hdaY87cMbn9mUkBwMEouCr5cn+qYVM5NFcXdYlgfnZWi
/RAZjUOtwLUQPqqeftLmCGfed1V9zOCfyH0SkLXfdOu8iBsIEx9MQSuAoAse7XXY
QJt26FjFAiyg6ZiySda4sQOBYFp/v5ahOX9WDH4b2tOHp/Y+dZSThYx28pyw7mjH
EEhTFuBI5sOEjzBRHFkFHEod3WqTSNvYTknnyhwm8tA+DmcDXdGzzCgDmsoVR7kv
A4rcarzNgG/dCP7Z42F87bKFmvBnBdC4puYIw5BLzVAwX/lqZ0om+YulxngKJJNE
FHNq+e3AQ1XqzmqVyEpGn+eTZBe+1DwJsnlZ4ArIyrR3SZvTLEYiLDI3UohVNtt6
bDgzru2AqI6F3dFOgxvQLugWAl2bS/C7h/zdNtTBC1ULieMY7Bay4zQ1T9Y1Z9cj
1xxsglrkFhnb+PK9P2/1Ck8JqQ4izywsGu2C2P1JnUjj8cSh2DFU56rd5yia7R8P
+ssxfnRmcneeS21VXMdmRFX+R+q/M47+Aa3M7Lv+XTJZG2zXIRBx82hYEmoxDZu5
k6PURxiGE0HJhEMs72aEd5z+GDSgXyCbPfcxL3bFaKEfbRQYBdLBts4zUG67PlXx
6K9U+1U3BSDvQfCW6jE6PSyPs8PDDlW61+eK+UJq+u9F5iQk4xgNmvujwbzi7Jg2
5Ude4pzD3+erf4gFKHtKnb/O3seYQgO7R68VstdG0GDooscE3aZYzbowqnZXRfS0
2VXRoo87/OabhKqisUSOODgd9gGHowq5XGnkP1XPVeYU6uHJeHb4u745caYjy/Kl
jE7/b/Rgm9JqFGZSsh66zQnpcGCMQB2dhJTW9qdoIGjxPLdFwe+iC09thaRYA8Nm
LAEod6Z2lD18GfLch9C0kzBnMRh7wKJCIbQVUAi+gaQCpkxf5gFJDYurZ7rHjL7g
vtmRx8L31ykj5PcWZ72K5azsbzW5EXH9YJodzzUK0DSjHBNdg22Lli05Xe7j8tBA
CnHQcNsEtTA1JC0HA0Tz18vGTqqc11PNb0FNEVCCTaKh6SCBYLxSLNbebGZWNvq3
UG5AX+KT6v8UBtPLD5TiKRcv39w1PbaEfv+LxiTPcgbC9KOWxCv4JXufMlIy2QB4
WSWeyz0GlEXVT0v63XpsYf3U2HjusRqmL++pt1ZtCcvclqG9NVT33MEHtGhRVP72
v9QVwbwT+JhxkxhVud11HwL0Sw9XdiJPmGux9vmyJ/t0i0zpOiW5Ht+JAMzS86Jg
rHIVK0Q5V6rwLV1lK4NrylbUBILHDbvbMMxPdmAA6kk6QY/dgepDjQPolKrXdEI+
C1MbdqvK/Op7Xq16dYQpjBJwZzs/HdGQwabLGIhQl+624AfPvrEJNwFO6fG1k+gP
gn9nZaqWgp6Kv0OHHxKlha6+VlxG2mkXiOYO/ef3GrwkcB0uhnLQmiCghCFYqbh2
ZU5+UzcGzDndXQZO5GfM3G42tgF2lSlZzd0YFkkXizp40Tfy39yYCVPzCRy2jqhe
04PXNMBUafsqSSUy6k4VzovJ3PrOwdRXB4YP8UIUbP+sjOQKjvn4lUAhfwzXOTGu
LnwT4Rh37EVDsgDe1tYjNbMsh6X9JTYQkH6OHRQUxZ7gyva6gkgeY2MuZaZCdD97
lRm3lJzfSORRB0MK1kfkF1tbLFqbAGeSfkzgXQb5bO1eqkYnyzF+G+sFto9PQOnZ
XJ6NXkrHVZRcLE2p3QkqycKUBuzG1poCAyTZ8S9kMe1eu7UEeZLcEsNsYnIc6wyn
0w53UaVm/mOhU44hBg3M07pDH6YSmQIPtdDLnmDSh1ARjOA7a1P2hQvpKiLK5MGj
mCtInirFZ/oejsoOEbcCPMggg27i8s4zYbv3zyHqx9YgHoapV3AlaXTCiT8XDLrS
unQdNrA55FLX/6VE3tqR8Vub+6DlTafg7iltZicH762FJ1b/sxptElwvCM5AGbR1
4HXse2b/pgOa5Gxw6Z3kVoGLMoEpaMaeLNoYM/qUuDO1/MmLLA4HdukUTkqSjB56
h7XcZTui0wL7t0igTtQJNT3xNcN5zXzs8aYRSKjtnxr5UjQCzBiYWC6kLPaGSqpr
YJL2HaPTzkXMGHOYoziUKf8FrA2ZBqlYrIQ/qiuBRGx9UyESkN56jbH+34cF36Bg
ZzIkyg2KUQvQ1gAgcOJ4wRvwH47bdiDGjz03l0F1W77bU85V5kVi+WuAWkH0zdew
cbbcuW9zP9Iw6AFd4sMijS12O+PlEWrxJP4kglZ/QZ6/PUnRCCcSCzi/3Z7egkaU
kVFNXoKS8wILy/wL5FPeFjVU/RbBxf7qNQJNCfqIMm2e6n96exN9wYz+j8nHVaZ+
aZu6NXwvQJNJPbJyZo3cYGtr7pGHBgAjYkLy4SbRUq5rullRZy44hd72Sn0YcmtC
lZzOBcC7dv5Qr9tpP9fJ1DRreqac/F0F6aJ8GVwz07EtDjtInVB325ksFN7arcYZ
tvaiBgW35tv/OHYlDW8tNoRuhSXMKzDtnwIzcXt+uJvbs9jpqOF1K+Hsh2FpraM6
L7GactKvxsIFBWrh/F5hTC6AeSVbmEu80BfVIZojdJW/TcjG/snPR5J0FXJZ4jOh
5LYJJIAQ4cBzR1lDWf9jsJIIqKhLZ57gsrjgybs0jzWWIk3TfCSjKUT/hgf0cvEl
wLBM0JQNBAqhGNc1ZK6xtZgn5+TJ+sZcoHcUKo/K9H/z7rPuxgAHEEZp4lBIz55R
v/ZdHkFsbOBz1upvbRVfjIbpICgiZjpBoT9CN4RFjqrkpKc5k2/t15yEOsdBlJue
bXw+vWtPQVfpRmqo37p6+ff99EGYAnA/3yUf3PDWrP34Y0M0TR3A9K2JkDA12hiU
QhD+c9Vgnkudge/c55ZWS2c6lGFp96TXHQ5i1M9Z2kkKlYflu5dQ5b548KeF8e+C
Nq/0y/0kjwkNrD+/fyIa2mYazLvU740qgLeQmhhh6jQ2qhhS/wmZ2gufWzixC15l
3i+oS6/pGdOxMF+cVZShbcPM5qyMQVgmy7QSyW4AlEthTL7+UjtwYwzbvy626+ce
cEImxFeDVszCF7wI9re9mGS3/I/PiRYuBPZN+4NRlS9JFLuvjd9tL/7HKHCnhIvL
GmcQMAbUz3XBz6jkzsAxiIII2wgwgR0UrSlqtj7VyVQ9XR4WFe1aeZsQ0Zro0R2V
nWxsyF3MVd2Nw285Xv61coJigodT34ykRQ1WJ0+1J2B6rOi9ebL0OdERKnKsm2P2
pAA1mvQwdIWBVId3NWyHI9u9NBvGKEE9G0hqhN4k/uMq0WpMSr0BRAljVLCKX8pF
d5/aXvdpE12I5HTITzrg1QTAuyH8ESjEdOOMovMvKwv56Cb3iFDMx0ECNcOWnDvr
yOQIBRNWSZxIzCWSXOmi+pu7VheeKhM/RROh9GXzKWPECECWZACZ2u2rablpixaU
/Aq6jUAINKw1CTtmXmy872rB0dxYZL25T35J6rWwhfCwh5XZr2GXBRMBv6J9Ydy6
W+SSZUirsy+Vupt1ncU0v15JJLqfKmC6v7ddcFOgV+rcCzIn0ubQ9/CGcC7AVCg+
dtazO23CNFofAWHUh8gEot26rW5gsntRZ6LTe8Mj14er8EDdVnnI24Nbib8osgkZ
QAR6179MVnxilmLaJQXO+1iqIxERKFR/0IGcIJTDhe1H4wCM+BUcEcG1QTMmtSqI
RnzwZCH1PVOdmrnUzqcxvK32G0RBX945So9ZWbcclzRmke8U3vBeM2rIRIaTPRxW
YHVTVxJzuY/e1QVN68zXmJqtdE63706H67cF4qMq8h3eTp3dUrJhD1qYtFxDJcLy
G2MklWF6ZG/pmMa0bJcD2qinZhn8LIwtF8OhU2NG88rcXumP1Z19YHWbQ2VD4fgg
NsAvl8z5drvL/0yDJd6w7WNViIXFbvy5ctVVX01Nq4paC1KWa35OUCI5soDIqgVf
WXGDNEkt/vbeTqMYJoouXur4Ox+DfCxcCVrgCcubzMDGiLdthVkQzhI2E0P1w2ph
7sXYqkiFztpRMY1J5uYQNu9fnYbDGFodAsO3YfgmaWBgn7ZR98yTmmBOYzkbONBM
yQ19N0tGmTPGA4AiQUv6LaGjySRmp+wz1GZ+ClmPiNDDcJduqPiGBdWDX9jU3Nih
s8MWXqyrhAcqyJ3ovIOoWYQeWiY2WZvMci3R/qyhDBOe/o1dhMryzIm7vByr4yAe
7XM+eEk6+aLGKgxYkpl0BCZlDNKwVbYzVyawvwoqXJW38mcIPaE5xz6w12hWqZir
6GOJd+gkCT8UtRMtIHZJcPv0zw1ecowyJEKuSC7d//3PQO1YONyFIM7bCVOID1HP
x376IYh58rPf36bsA+hSsGOtxvHJ/nUWQGEYFTp9lt9Smr/doBPtZ8wgJXPgFEZs
vcyusmwapCQGb7/ZejcZZ+/F+17k9SgQQnwr2JgnWc5hw/bsQDBdfGJRtl2fUX4T
yeebi30TBYc5CjW6RpPfXKAcuXr8/lranqw4EsYYBrju30e1Pq6qCQLCX2UVSjmV
vZP6LefkJpa7t36CaEecvn9kGGMitSHYr1Xm3Go4hwbGJ6g/z+za4bgUj29FNV3L
Rd8PFk2Sp29152+zSIPYvB2BEtx+VFOjBt2luxWUSnH0sIY68xsdH+LD9zUVDwoj
AKEALJeeN3KDCkgJ/WzC3IrmMPFN5u7ZvP1GvIj3SxTke7DqBZtKAR7qvN3xBa8X
DAv7+6r6PJEcoZRAAI1mMD0QqrAlGIv6k1dvexOoqqfLLnWhz9bFEQM7C8lRtFlR
2MnwkkH17gmDc7EzU5WujgfOxVjKB52pnb5Ou0mlRCQkelAzIN3s6LiMveLuVLXj
BZa4g8lGtNjncnhChBGaxZRQM+3tnqdEqTUfqUKj/5mZeM88dROkt12Si20fAsPj
mxx9s76O+irvkUFGvBLf+6yv/tS50smSQk6OFsmZgD3ljy2xhKrP/3rJrr1rCeax
sDf75fQWI+j0Svu+OZnqt6tqoKvUFgERp7sfQIUO6/D3ZtKCjBkY663O7rRtGMHH
zz6cHjocm255qsvWucWsnIfMfoFj3+XGMjZLhQxazZ+ywD2GFqOlg+dFWLhEL2TF
Iz/F9KabtHjMdWTQcv8jRNP4NXuSX2dYV/DOspJW9O7ij+6JWV/LdieLwxF59ioI
H6S3BSvj0CGe+Y5bKIvZ6QfM2jorY69Rc9RcgOflyWhXrX9f47tEkZt3sxL0UAvN
zkCb34UVlA2gvNNtkpcg/BM8OarybKNUSlwyrZ04IuYBXlamtIUPp86NkKn97et2
fOPJqiPbJIRkh7TMpzN/zifFIAzFCLlyNHE/Y3pBw3ia7r4gvRrz5J3EiiHQDxKx
qWIQ9ZUZ+ybXskD09JChX8ub9JmYGYjiGno4W7BlZzGOjmkDeBYbPUIUfVgJViA3
Kcr80XPKX14CcSAsmTs/tcADx1owx4bi9ANDPsBJsEX2v8iszd7mZGh5xjP8LU3z
7WCBy1apCpBu0tKaSzBxmlcZ9OF0cpbFKlCNo+4za+1tQgW7o3+7zNqeh6+Cj9FM
c1TXWCEr27LLxNOcYr8TX6lmG1Dsg3CJEGRV0Y2KFekZHr9rFUCAqpG6S1SYO14s
iX5q9HrN2bk2PV4a+Hbrfs+Idg+1uZMDwUT4qmYg7L0kbADG8nlrVr8OWIq/UkVI
c2zrqOC9K9xDrCkzmKpxFy7XuqxEPgt4mNxP8Xt1Ykgt5dkoDVEd6ksxOQVawhx4
MKu7hEBZ50ys1gYvr2JbWGc8/GiYMqtpQJ5/o22UEXx11vznZx3A1MxcL68Dorum
t4OOFeVbV4EfCUJeRRPfSJg8l5uBeN7N9EkflxQxXIRhDXbp/ecampJ7ACU8IroC
SirdMESfmoEiwqEe2t0pnQqP5PcmlSqUib7COuWilzQaDl6y8ZJe6HBYz+V1QEeE
rojh06yflKeB6JjdquLrcjHr1upc35YSaWgR6Dk4kiDtPfYYehP8BlnzPNXbRFDl
/OzHbmRvfjf2Ohws7I89XyImqF4v2mINPykcfUb1eTYVXNiXBJ6EDR/dPjgw1hnD
dlooqa2wDODyuAI+WbXMpKyCFWnGQyOOu2dM3d4/J+yGGnP5i+uh1qg6GAh0al69
9qiwMWq5YW/KgSurUiAK6zY68HgsAdL5qTrTkdc8L+0oU2kJ3PxghjD4O+5jR34k
m68qsAPsnY/H+amdUwgo56qFe04W78iX7MWgQGSx0eRXN+1QrcjIXiY0AkpRe22d
xZ/snHMH46p7bN6/n9FZ4PCuBzxWbhKH/TbVZRndojaTMC94G/i8FLuyCYLV4vRb
t8zQsoFzIPbw+9wRxqNIvp/nuP9GUi4TILLRH0Cz1sNr5f0wH3k622NaGmjlT87I
MigIORSbDpb0AZwOtTMXxHThpjTLnkZtZSc//5ZP0uf4pwsvLDzWstV6ezISaNhI
kNKn40WCBQleJE3sd6nGI2nq736z7QUAMKqiDhPJGaKmp6QH+1sjMjLU9KOxEZfN
sLEDvGI6CIxEkV67FDcum0EKIhYobfW7exUwReMj6KA4Q8UZS/JngO5Plub/jgMB
Y/Bz8V3cwgyRJTxTDEb0AeuK82sR+6jpv3tPdVUXhc9gmVCpScAnQDgFWYrArduz
apZylAgMDzMpMnjipfFmLWTQ9FOKFe2qhocdRjQvijKjjko9sn4wf4I4wwHnpHXy
Zxy50k9LrME1Wq7k+m/b5lkfITTPwj5tsWvcRTf7A+1jI+fxUpmUDAYkQJuG7p3W
U2MIZFxhDTfFu8K4Ru0oM0eN1PF7YJeK7Y55KoTOBfPqDlGjPn2XqFkVGcUEbgs3
SQSq8Xr7lrhib9ZThXAJs5e91y2yWV2k2xjr2m756K7fVYw61Nd+843HXqUgzOpl
66vhBPg5x67qpP3mdOKvsbApo9JKhryh1oxwbgkP1s9HTfjYc2/9pGV+C59UHfDu
VpAIE4NaVdPm8S+fpuhx+Z7hf8PpvjTCPTuwbmwRAmH9Sy7g3uU99w2g3RraRYNQ
2U0dx2hrGygBQJFLsfjejuOLcJJmjIrK+EU7mvykaH3KntM6EajAEEwUpadcGB6a
hv3tdewA+JO7cUSc/kxMbKQbXhCg2mQZkPZJbwbJoETrdfOsGlI2NSQHnQAr+mmb
KKE46SO2IEJNdYok+c/lbBn8xDuVG/Vfe8RKe+HdELfPDahXgYqiqt4JeOf+SCke
KK9FDHi3upjloYU2zoMFxFHu/9mgaZr67SQZa9laXhgQ95aXUDL+mkG5xX6RGunx
YJb7tZ/Pc8n9T20a4M2/Hg/kd39T3rmpnnranAi2hBpY3SinUtHjuR/70Ub8Kfmx
bYNNZEwZpxQO0CSroiDPBhwrckRLzGmGoFtKYO5yELfm7plfStrBNIM8FYYFhp0Z
HZ48JEqIEuK3qftVRpQex+AEkRwyI5AtniaL/382kKBHjwJlo+EiFA8eTOExSHog
8BF0OfzhqpYvyAG4ukDqIDxcguDvbTlzqR1uw8t8/3yD2FBecTgmBkJ7i8SGgFRS
I8HfINkoAWrrheUVxNcLimqY2SdBU/XqtfgeB5TYyWnhObPr+Nfi90BXGMR2MI1Y
LZGircbTgocSTjrbTscA5cTv75vDW0JYQa7HS8Dkv09Msjp6179x1KOKPhx4Udho
O0B9iCin1nnGRxa/nYQRLlXKzM0WEw9muK6Ecf1scAsrK8kv/G7fRZayFeRT2Blu
GH+EDibY4Ni5tgoBvhyAohPlfjD4ZgtZ93unnUQOT2A3ng/RrKzOPHcECkYORMlI
goF5vH+/EqTCWnuY2vzJ1RLw9ea6H/c1DzleUxV4mtgcoU4GMnwajKMZr6rUt+cV
FHyIGU+lp52pa/eNa8cMSSjf2J+xjYRp5PrHWQIpJRHXzAEOpAg7RVamMbOhuUcz
oOnzitSvub99A13r2MqY5ptf0p778i+JMWQ8qXz0bBUh2YnCgLJkVGj3+TH7/a5G
GIzoSOCv+pbjjehyzMscuMd3Cg2rOdAWd9yaPQje14GJF7RvPqIAOWqbkQ0vAck0
UPT6tp5OayqDGOdZuKQVMx38aT2KgDXTkZZeV3TK0tkaT6klsrDEEnyHRytu5T5P
Ft+GGHTJb4Br14h54OuhA+sLOxpdAzLynmdk63Roq1gr/CvxA16iwEX9lv2gKoyc
Ju14J2vtLh07JX+H/7TtUY4dkkjjy6tLvlkl5cUr6F7fmmI0fDo/rb39jxJ0xxkl
1vl9crh/b7XJTaXfjwIgxPXWh7QJzk5BaFsUSWtv2s8R8URHZzS9ekAbkeo+1E2r
OEZziyRJhVIDkRU1GOqahfWK+CwMjoLZyzq7E3wrG6RWvvE7nNOZ9TljpYP6+8pk
FhdnnW1kfvYXuOsIEzKPRJctiII44ktAw366TB85bJs7Mdzy+FSUBKKxJUU/tkU1
+PeQ4famQQhZXYJ00mMTHnVsddWx68QpzS7pn47yx0t/pstFfhvzpXLdddueWyrK
84H7AGbA7y2IItvBNNBAHIv33Pt82vDVx0UPFc7lByGZGvsum4jfdO/kh/dBArcx
0S0NmJ9DTF8+rwww8Ei4QcAY2x7engiELDObrdCcYq0bja2k9IwmIHJL7Y6wPFtp
cG30Sux4u1bDpEle0ewc3TzdXKdtsJwNolTZN4jdmC7YaUA9pWVCQx6ZAEf45byM
X5XOZnl147HnQT5R6/KSWIpgaMav5AcANPrls57p631gdYeakcQsq1x7ldljNBLI
6w9ocby8m36fTmFxlIvqsLmxhaPRjXrwsZaJtU0ogA1WgPkMnJsYaXhNaeZtDYpq

//pragma protect end_data_block
//pragma protect digest_block
GoBgTsu/X4xDFP/Iv/lALxofvRw=
//pragma protect end_digest_block
//pragma protect end_protected
