// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PFeMAKw3JqD95NtCr/kFbCcEa/hu5BbWa0oqZIOFa7n0oKuOFDT2am4vWirszy1nyCzbRRHlDSQa
KH+2ZK5tVMHSZ7XUvD4q+pFxGMuFbszVCyegUF3Wd2kHRbHVCGL7OkwKRGbXZ9W+Jg8BNxp8Z/Y0
rtzy8j70/VwB39TWE3UIz66obhn4svwZzHRusvUvoXzD95GW0h35F1V/4YJ0RLzGtUOdXuOjM58f
pQowAWpP+gsKf4ceHFhxfqImgfXFFVHwULauOx2JE8U0CodLSYfQ5FLapgK6dDEo8LlSv9TLvCA0
nHLMcdpqsVMJzJ/2AhrmJ4hJzaWFqFb39bFUeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7408)
PwJUcDtmLIhTvH0zFCzUPg71f0sSdampLT3aHiYw8mtuBYemhQudorMk5W3Tj1+15NeSu8R+QcQ6
VYcBaItrAbes+lqDAP8wHtfYdc2PiaS9oLG2ObXrmoKPpkuLXMgPqEXs4q66Hmb+Or2UUq3257yj
8CyidMjbtoibjRycgDTLxyOrufDVpSwPW3NTMLF+H1gVyq46JVRcS8hr1twMzzhZhBbxLnDxM+Ye
WFml6voxeH4WIQV6QG4DHyJOgyFt+E+YqnNf3njkxlJVEKhZ8JanzYhm8GvYgWYziz/ppUH7kFNj
/f9gtVIUL8AUcVDj4qj+ONrW7ZDKs6DZkZe78talFoSbLUYdJ9CkIlMy349nEOLFkM7BLY5oVw/E
sld5BQkgA44Bs8zIzdoaeWZuxuDePIcJWxxPVidJVmD4yxifPv/Vuvjy0zpzDIu4nff/smcwz4Vj
Up9kzYDb1c8StzUeZ5oWCccV2DHLC5ITMmvWBnieXngUHCgjEI0/tjebAOAaoLRUr3Fn8AxXiwHb
iLprGKarEDuXzSYmT8AQeaAYxXmBqFGLBj9nh4Uvcbj2rGOkC4u/Zg+j8lSfFcwTrG7RmImd8oLQ
w62GpQ/XU/bxfIn5yOeTmAVVgnVGdfhE+hA/AQEMhIzpmv9khqegWP6QxtR9qiSQReJYY7BYyvyz
xoWAFS5w2qAAE3wQa27/Wx4PHjIaq+X8IOmojWy7BvIfp6HAYxktv3fwRRbkx78s1WeSi53vABTF
FVEqp9p1YLeCkekG/iEqDVlAj78cfK7l66oSzCBKMyeAId8661dbCWylUE2X56sLG2++TfcVa+Zp
zM2OcpraIjo1P0nb3Q9hSGdo5/LqURRmJFQ/pIXMPmMOxMBZ3QnYqXFrlL62M8+SXUP1KaIhmD9k
XtIzjxr+F2WIDqbsS8nonSIxTMpaZ+1Y1fklYaU7fLUvCez5PYSo4cZIrIXmvMXfWe48UVyo6YAb
CMqWOV++bWoWSHYWCRldysY95DZQb2s/XBOu/bzo+asV31/fgacgh98rihK/ZBi34aUX7Ve+Z5VM
Ok91n5UHgrksWc54yI9QY1BSTWyVEPAXb9yym2lV29/i+4qklXUoXFfrwPYTXwlJgEEJG7/EIXns
hc+CGo550YuRNYYYzsOjq+wFNbmQwh63aLDCMRvt9Vz+uvjC8Fw1+xUKSZY8AwC3Ttq+gilM/0Bf
4mJyVOc9xuk4xSFcPNgSyF3egHSRSG80TRQn9ectKAotSXDNLrmEgfQoiodHS12cqYZXqBKHUmzL
cVsCf2l5na96bISA39aXQt0TH/jF+dmn/sOUtwpveld06TRppRg0OAsiqF7x29F/hVHuTwEOD49x
4LJLUXlZhsgjzojffSz3LzkgYwMFMWmQs1cv0ZyX9K1wi3apzjgl/4Es/9dh+nUj+B039azTF5P0
nkQnbb43vvWlNROLjnh0pL4DZ67znZuqg3tYP3M8xIUo49XAo/6nVGAYNlLtr0ICCIbobvvLifCQ
t9IbmFSneYVu/6BxGm9WvBQKwTuwTonu9WUm17gmtQOtWa4jD4o+/YVIg/953dbYM0F4Rcns2RZH
J6irjhyKFWrrOTOaL/wgtatk3nhBLCtOva1W8xkwi2NNdejH76ZhmEBfbgoonHEJ9w2jrkYtjECa
gBcsBVvcrrk0r6OcSwVlDaHxog3uslIJXvoARTwLajuhThlBR91b9kHJtZpQUIsZWh+UHinc5evx
dbaPuL9GMSLiYohEk8jkilmrMfbDrU7wnvKHRMN2ixRiV1sGqg6LcOgGwFts09IlF+psbH6gyQah
MEVTAKPWINPkwpKK0VpLN1n3x1uGXHXaTK11AiW+k4AdirLseFTx8Y5ELMw25gOrQZoBD9gFoBKS
umF5jbbDm4CjF4dVlXUTtPS2meWGO49fz5GOMKYyxet13Hcpq8VTRuSSf23VvqKvFQD7oxAFxc9a
eZdRXjSN4k6i2XuFfS8w713Tf5/r9av29LbqLt8HrxxD1sjTBHnxwYoiP7hFUV8SJOM7LWG7Be7a
clLXOqEm/ws3WNjtllBbSW7mQk4iVQlgH2ROMY0L2UzVN49s6LkGPFjBl9B3O/EYyel5Q7otLaEQ
PoSo4oZAIlaczEJZ3/DvbrrsHSa5nsIFedlNqriSdsIiSm/ixSU3s+yoUT5DxVN72ApyCcjTJOE1
uqimS+MbdXBKzb/UPJp64fGtoTxlS9/4tSZcjELPkk6OeyjlofSLnpWy83Htd+aso0v/KqICL0gh
CRRsR2koKMREgc1v/Udza31JgvjSPBduTzNjuO/BdbX9JV4REhHAL49ubzWkW5N2dzYEsHAKQQ9n
cslspK0PZYPdWBJBQ1pOThi0FqlEsrA4YUkIpzfu0nFekHddcYU20c5WikWOelXKELfSwtNB8yVP
WeTy/z73jRlytN2aFil8031vnlW66JUXT2NODHth9gMTa4meM7na3RS5uEfY1IxNWbuEaI2oHfJf
FX7ZLrG7XwqUwDKcRK4V8ojilPztGOPPjPwuWOuOKgSXFUDG39zFp8pyABCtDD6eMAbMWjyvPqyP
s7QyzlKulAiWOvXJp2YclbxtYKtLhvnIyOxJ6cRBcY/TcVK0VDLnRraN5qa9euvH9eHngzCSskVU
O9yV1joJZrz+i9xKOsmQIuEyZcJUJz+vVTJYB7UFqG2KYzPHrlNM3DgvnJyADQ7uejDQAVF6SLJN
CcQ4/8L9mKRZmiR5O+szQuH1169S1tfGWbU0+duE7woizftKPkrjQ43hk2GzUzzVfrggQYUVzw/0
OSUX64GckhD8l5udCERUxlBHrOLPNSP9RqO0VVuaxYXgAbN6tqSOCBIk2QLERnqVqKlHVIOa3E4y
6o3oFhWdWqyumhcPCG2FiSU3pk+OXxwulkgQ+VDwVuejymt2FbIe0MnHgJ5HU8wj2NAmP3QsGhll
c9Itq+1eeTuWtmfFobDL8cwKgPy5FDIihZZfgBT716CVvsm5dvRbI6DcUnr9hU4/ELNlaYRQOS/U
+2BPBwmfgIdwIhhmuRKtN2HxangnByL6rbZFPrDo8ezMh5Er9vn4MrI6F/tgc44dZF8eh4XEFL9C
JSzSA9eFgYNuRmzHmEXYUXHD7LYXR6m+jqVqOkVhhf+7oTogMixj8lCBlti4FeSPHUScjnqXEGmE
wFNBrbxK7A/CrU73Uz6u2W6oFqgPc3H7nLLYFJMCpdvT65JwfNpnyOMFIjcr9lB2ATD2QNKBBsYU
X778QYS2U1jejPERaHNzhFrSgi9Ww+/Xs1+Fwzh6ldnhzYKAHMna7X6rZLPh8FOs50rmKe8BVBJo
kTyiwM70cHe14XT4CaojDm78INSCFQLTr2NK4FZIfR8GBK/7SoAsB/+MI3oRqCN9nn2wUb15Yo7r
pxOXdtXb9RGrkfl+IzH6JyGTTCj6Cyz3CNDojxZGyHFJo54VK3sVajvdPvNdl3G+xVGqJoFM4B9/
qUZZYcoKxr/FY+noQ1vJ3Y+NKq4TFucuTjYofu/WdVMpTWpTIgzl7r3Fr0rhc/bbhZfQ+yzltp46
iTDx2/AKa4L+qo8H1cG4QWWluEnqEp/TKTJ6ZPX85PUIet70+iOnI2NmD2A8SjhX+jwRMVK5hMGL
d18YeYi6NtUt08C2FzQRm3zv+djbaFR5eRET+/SUsRhS7j5tE1zN1aSgxT1TRzPaQw1inn/93416
akiTRiRcTcrgpcctbOCcGKxKr/n26sNyE7m+jziBDROX2CPNcJaW5s7RGqZy84V71rI3Whthl1B8
qxR3j4StaRSM3o8nfbIs6rmcUdfQ4D8CQkMMG+6TS6V+v24iZh/Sw1pd+kMY+8rh76nrrMtFisJc
ucQNk6+AYLYJ8DtGxrwH7+Nl6H3o1FDyKuVCi4tuHDl+e5YRkdxLi0bSCYo6emR/ay/VNDXlQJY2
BDNBt5ToTYmBdnrU2e7gCNZKy/gGnFUWb4aXbtVREoCoaU1B/FzzqtLxoUZlM5NJpRhfhb9WCJ/f
LZobuRTgmUkrqA+14/MlX9GVok/qIrqA2ID0DlWZzf5n8SBfulH6suiDONJFK8mjP3Kf21HJcnvC
QEjiiuih3R+H1tsA0lLYxset3XWCptWKJBBBLK+Kt4ZsDPIzDPVVwMrsF5LGfu80T2RxVv4Z/614
OI20JHof1I+5gkcfMmXMiqZ9JeCuUuFnRsmnswtPG/r9QwzGc7+qToo4TVK75LgThbOK1VKX/92P
S+PEiEkds/jg8Ncj0CZz8L6K8z1T3hhYJPee4W6YHOILtKnzjHEAxD/hewwVhKYC263SnHqn3tfE
GhQt11iVIfMId0NUmL9j3hJruOk3x5ePOvSnJNkpyBp+KjHejdMpFI2xpCi6XlLyYKhnEAhheQR7
SUdtTOgb1CdntoaFKkeQJUpll3bzOO2m+EqL7j3pNh1aHckQqWFXs4pEHptX4lJtp9+aB8eQy+TA
FCZ9LHJzyAkkpZkRMC4/X8fx+rmmusbTMHdzNLfHDldv9KgUJOG0h4PxQ6watFHf/EG7WSIjIDlz
jr6cPfE/fnClJwXf+vR4xtEdvqNlVYfHYK8TDLGRAyfHsJX9sy746HJC0p9/Z6/rhylcnA0o6MMP
d7HgEO0wWeEuBUqLn5kVeyZQrBa+CihRak6XA5suVqOZ8XHKKeCJ1SC3hOmBTu0s08TtPTqp0hci
ParBnVOs5BJQOkJA/T0FZEYmoDhOezi4Q23x98mL18yfkN4nmLcv8Cs3z2BOt5n6NxOtV0JdG7vC
MaP0u7pwnuDtAdP7FL2svb6Oocklo7uzGTeodIW0mHgBR03aCiMj8iDInAHXTST8K+Au6H7oDajG
GjGHNGysLNQqqyyifoALIjG6lqmIFGYIXNP+OCp5rRQXw1UAhrkf9sqi+Jc0TQbKgK76ZjFIlJ9l
/drh3HH4FDxLj6O37PYGMEdFjhJFZKmE7t+5/zNVHTbTqq08ClX/398nLp2mGd0yM1GYr0O6lJFw
4WWRzJRlIvqxfM4YJHY2E1yPUtEoBXgM84gMZ1UtatNMvctR5ocQj9s9I2XiNybwhpn9Xp8fp1fD
l6vYtaOYbo98iWwBhs4Brl0d+wFZkkX/dpahon9BnXxFKIFH9vgy/UaB0ydfVD9j7C/YdkYjq137
gp3XvfOobJD20c0t7aC0v3mIP4AO4AMeggiRYFs313yRL3S93/6crdczC9/c9ZJJCs46tTAIhcaK
Wg476WjUNx8PqDo7oSTv9fr55paEQBduHxoPzdklesDPyZBuQdEIMMLEfLs+kLHm0iOUi5FXZ86U
7GfxF24GAZZFYGsh3HjfeSPS9Z1JOULk//uADoZJJAHo/4Rex5UKr95vfjOaSaVps7vCdvJXcefb
wdOe6r3wMRhE24Hl90L+yohfQuSQdoC37YB+trFX03ZYeqyEIsPOHQyBMCcHorGQ/+RZ37wytt8F
hYO9AKWBktBgZV2+Krm3TcANP5KngHfUvvdWOCew/HDxZYuxKdpORLrSELp3SFeA9WKTwg6DJtDu
YwQc4boFmk/JB5hLVYa3h9o2KsyTNQS0sAvUKwdhDYjzq05CK3daLiBvz/IX8yNIGd0WtpcRVXhT
9XW5lgkXYfsxE/fxWH5pVM9PkHMQjtCzb4WH3PNFk5Lc+dwIxg+AtvkrllXnAE0bWYS0Q4W4ghRv
sazKs5wKqbBmn2KRFaNKJ28J90RzGi7tAmlBCGI+k6mVero75zeP8g8vCVkmgrLh4k3Z9diKQC/B
trPIPt5Lxa4zDW+c/kPumobrc1+Y2nWeVAfjmhlAaPmcW8hO1iU6Hlb3CDTYyUMj13vp9DKfQ9mr
ZYoJI2CYcbMGxIkWR/w4aIIZdMIuC1QgnnzBdXOcgSMGuuXqkQuxgMpOzGV3eMckTZsn6U9yXHA1
/YX7Xedcv6FfaFAJbjjAUkIudM9UD+KvAyMzHB/3r17HulhWJJkJeIusJ+lv+6yHKmFjQOzRyRav
43N3vOoXxKwMP0R8Yf7yn/4MBcBPkCqattoJTDS3AvwWskyunmfsoEadb8UhYd3SjI9U58Zql1Qp
QJbuD5cgziqUsaAZeH0QU5odZcUsbVnzVbIeUpiIu01JPl7JoE5lR5c/vxJ6bZS2vnXehMkkMJ2b
aBg1YRSoy7W+vh70dA0SBbp+rH6xvWiXgr4Q3+3yc0b9gIt2Nod4OEds6mbQtN9t/ZOQQKFBIC40
3gStHzzeV9HHUMUQPwmSdmp/ft6IyIKRxX+NJ4ajLFIT+j9dxKzBf4PJ7viKk3AIzvBPOwGdYGpw
ZBOa5UBdlS1VJ3cVsTlCRSG1I8d6PiWVgbZcXXDGOP0IQFgUcgZkvyOYpg8bhIfecqI/mVa+tw3m
oG6kpC2er6eTafbpqJGdQlJ7bBFUNoEHD1jfIia+JimeyKyNAlvy+iyF+4UoDz3ItjP+HPSbN4Av
CSYhNwPck1dJTDxt5iiTE2GuQViKaod0qPsB7OvIPFpJCWCqynXHSGs48CbhCYt4VUtZdRGvBdlG
95OeaZEzOVoatxh7C/MVyN4DUQn+v5PLz8RPi5vDmDMnZOThwQciB0m8Ju3jxeMyPx+3IMmcYEtN
dt3K4s0YyfB/yDZi8XukTQ1SS8qorCnKhscrbNF1OYK2xMLupOEJMBrq3kzPnlFQecEKBfgr/9Wv
PbLcZfcqfnuViaRhoiChUlDa5fGRt8YE5h3q+qoKWPPAxL0ysIdCFx5QugGk9UBz7ZMpJW/NpBM5
4dgVcgpEykfAsHAbd9z/hZaekCa4vYf/M+I0Q2VS2BZ9FixPoTU8KvRL1h9Fh64CaHepFSxZR7SO
FYInKBPUrvv8rog3V3SgHqH085AGJaDj6CCxMbIq3w6fL+0tfsOdvIEOGWGRYStzP5/MF6AhzEPB
i1llSXfdj1r8VcZzw3OrxUhBOC6a8gfx6zi08K/NQ3Hxcws2tDdshvqn50LhnxzBwriJClr4tla5
SiaA+0BW6QS7zwYhnMtmBivI2GBM/VGq4nJVRiCRUG4jPu2C2Odv+/IjkQahpS77R3ESd0qyQmM/
8Ng2PT6PHfNnQDTsTsQ8+G7TOV2Eg7ygPyR+x+E6C7f6DCH/pKSYeSyfDprhWFZ4QpAWMS/KtV2G
VF91o2RFAuTicBGim2SY77RRyd6RCkGl3uT2caimKBalJfGgqVvcnRoepwb5U9mEHrY114vztAKE
BshtDtex/gzGjGhWYdIqN9vPQK2hlQkvr8sNbMJ7py/nT3/olV/vgt4V/Eau24B10YTyzkSqqlWN
ko+UJdLoHsbrRrqoFQRiz97xelVGLhmZLZeanuNz0lh3lhbzfJEy0S2UMGkmYU4TC9a25S4iB8bb
+1Sv68mmuUtvPsb396x5JfU4TTBGhqMputCMsYnTKuAebh3o5P3X560FqlDFG6Z1sLe6+0L8Q7xU
O4wHo8CbZuXzNSnAxTdanlK/KgjP/9FekZ4pRNk00uTHzvMqs/qUbg7B6eWlt34J/o8E9ON3XH0X
NYhwmlWvk8Kah2JICxn3zGy/LffM4cHL9KTAqNfv1KmXshjuqyBv8rNdgIXRXapujomse7zdKla6
cfzr862IkKapX8KjYcY/coPA07BUU3zWt+IkCBLj85n8B+ZJcdDDM7cT6N+bc7wSDK7QuExPapgw
FTIt5oiwklEVtt0SRdOuHLXZ2mN2KnCMx2sChk3XuIW7jzgRCglpH/weTbgdmgmXTozyK28Rr/RZ
PFJUWzXfNdbzQ8FY56NLrhckrdTMD6IBBwRxNFz3uRudug1izPm++psMDO+KppK1kfEuZKG5TvGo
R9O+4lmTSbmNTFkBvwWzlmZEWoZVTH8CCJc339zfwNBa0RTId27Nd06PCiKHFKfsLTi2/WcJw9m9
ggSgwe36ISdilI0sv5tLeHMdLAG2nT92VlZjsgp59Rr5TjMEBOsxQY4K7x317b208vRAHcJUEPS+
gJ7vDZwcVroXzPMyGxsMUi3zbsSeObKp2q3DQOFNsOWRsDeszUHMymlOQK5u3GhDDx8YtySZRXZ6
NtueQ87OhwJuZsowR7S61pRNT5nkVXokLouvdwfoJw4X1oHrBilVlQBmZ2zFzbpt84cwX7RXFY/I
Qygm2HPz3HW08fMssP/IljVDOzdy2zyvbYCO7KEZys1SPYwJHxwo/49gjC2o/Xt58CiphBbErdfk
wEF5gkiThfb0kO5TtnMUjbLAbC094GEeUrjpRves2qSwzouUWBcxp2hwlthVqM0ffGDm6vFQD0JS
PRrMCdeFoY7tSWOu8n7w+D/iU0jRxkZ9JPW7Irn5+BGGk0tXodxuqxnF6p0E4Y+UZXpSvxUAVVhF
y/GSV/NDFM2plOjZsfY51OKXIo2nRnrcXIm4QZQI8jzcAu7woY+jopLUjaHl1VYOzo/FrU9V246q
GyJr6q7v/b3RF5hsN27vdASGYp3V+IgP390dV4tdi1kBb/b3chNdmnc0ov3UOKvV2j2smfn0UCyn
UwOvRqifEWUFAg8SRuKTJRFWTsv9D8u51AX5OpomGU249RAPjG9fDtw4xCW/IDCuj2WBqJeJ8E9f
RJrTNMivVCMboZ9nf4BXA3rgECMnVZbnoOfxCPV7fw2z6POjETtT8qhk+Mr6OMYN5Sf4GVswyvtk
pke3ksIAfPNvItCMnoIsiFZcdrI+/psds8wqyhgiTEdFuflH19fjG/ZYBTgLXLbMJlYP/46sx0JK
XvoVv9+sIh4ShYl4tWNql8WoiIu6VU0vPlcTxTOEkLMXLH+1csfxIWr+sjbr1xJ2sYLZ9EnJkmBW
k4xvCvz7jveVTNmhKtzxuuNeHtkUewnSkkJQWKPoirvsbIUmo2kUisdM8q/gyXC3INbO8wDhzVqJ
TH8CbCFgaDh//RtOWLxQJq65fK5fh7Uam1JLf3ocSIfFahI8lWh2IcutWfya9nCW9PMBoDwIIylt
R/mGGYeGXN7hg2G4/Yrr0ZgppsTFdvckDei473QeJyFRqVV3g26yJJ9+be6JxLrXNEied1LruY4X
s4Ag/dgFyv1hZMbFDJ6xESo11yn/S3c5Yr4pVyJxVp68OzjRJQKlRKr6I77cwYYyENysuPniIk0d
v5GayMND9KuU6VTyjgWxRPT/3ZEJMc8EEl8MQg25nwVoDjhBjjz3qnLCz7cjgPshfyUamKHYThI5
RL8HidvmnlM7asuKZeclEhMiVhHhC15iP0PUBAgq/wJqA5hFIoI/iCNzjpJYho0eSjdc630d3kVW
IR6amf/nM45bq6dOo7EIibA5aXdlZmK4HRfaO+KyohQvbMxurRApM1PEGRijXF6ki/hzR/aSaNu3
wjkXyYj137q2x2+tUOXvLlUzCBfH3ObvB2wXcLXaCwd+B7n4oo01jvEKdi4coKAgjRABtYREc9lU
RFecXN5gwV5VoQHOtPVUxBY2Mr1MAt3LX2VgE7PV6PQkLiMm+IeJ3kAu8eXe0Wv4igrx8EUaon6V
BAa50/I7OHRDysOyIygYmU95R9idVgIVKJaKEhtxOBPsU4MdX9IsBfiBvjGZgfwvTUEG3RQ1hUQq
thXdSV9vAEa8+mVr82H7jNKoJ53G+Ck628NtVtnZ1aQLgauxJd0YMAvnV0Qw7G3ohEjMwzg12rZE
dHKpADlt6wIaLw1SPz7yWXIm0P9dD/ILbdyxlNbn7vV9Lo/XKJUfyWjYO3MSq3aLW0R0hW3UcWSa
6gJclIARjJKkFTiWSkHcI70Oy2+3oeyOZgaJNIgWF6DYwRkjpNsjhtnSBZ+7LqHqehvA1IJ3hBZo
OWY37ZY6OPJB3P8RuckjZO9GtrKmb+SefqI4Y8uu7QN772HwM+pXwsTZ7h6XiWkipGGudxwPsw==
`pragma protect end_protected
