// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
PeGkhBRBa/vQ+vnOwPw3Vb0UcVUBoSCTYNNdhdfHRyn4kpRjUlBaGmk2LNWFvpSE
9NZCeVoCR+I2upyPIzFJjFMYC0WS3wv92zaOeMekN836nwTR8Sm6jLxG/oqJod+2
7oIphqRQ0JaCDv3kNAv3a+c0x0+5tKAlA5BTpVuOqhk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26496 )
`pragma protect data_block
8d+V1ZuN8IXKVecio5vZj65IOwZhgMjhAjSGeThfGI7V7E1+zSMCcqgAlGd6iOTd
l/Q0xWt1v0KwG8bAW5c66IB9A4iuy90+20hyPV3iBPNEcqKgaMPAQ+B6tUdKX0dY
UZYM+c6U+0XW7e5cLLZMOSjJzuGjT5Ot7P7IRfTR3+rHQUMq1l2ysz+c+VoWXmcW
OuSzlYUcYW0FG4Ou2mJ87pkDpUqHDpsMG1s/Z2U7o/haOOZD8KcPv6RftUIsa+En
GN4QB5U4tmfreDENK+DVjIEPhJ6azFG+VSGWbslrbD8y1keffdpeexFHth3VldkM
hhmryD2yMEF3Xaet/y/CKEgMBPM5OMa3q0OrIefDmIr/sx6F8l4jfrLds7f5bH3f
6gEhUosLdhu2ip+Mf4fS5LUKqfVQ7fCrlMY97t7tRjCzXDbiG1R6ENNPYSNyow8W
T+D1+EcKOlhikb1XTsdyTap3fBDCn4IMC7t92u2s+Jjfm3hMg5Ld4flW46r21hdr
F97bESbKOdpoYn4vQKdXplL3iC/CMdJbF9U5kmj0FkzYGZRqe0MAHUtVPqHR4t6V
kvPAxbqXx6gy1qKMwyXSl8NFDsL+D+vDJoBCvuB/h8+rUpZJBx63OMy0llDzwV0q
CnwcVynIoB1OblmRwKd0Af3JHiCsHc/h3KvSYkMpCnFHL/4yKN8iiTPbNr32UUAA
zkBGehfxhGe+1X4EK4vDXM+2iApYrJSQ0AXmWc2ASl55yHjxGhvmxe4Tq5Mg3xvI
f2ZaDdDs9aFRGrirN5S3AFjSeEbOl/M+T5uyOG8ExzFEjR+TXPPJQbnd8mBpqSHy
a5v+6kRcOLshH8sRBqpPVCA+0/bXKSg7xZsq4IWu87Qmu3/fNbZafjE2vwlkQA6N
Jp5/byqJLJIHRSEGevYleRnMprmgGUt87B2c6BEc16UyTSyyn926H9dPO/Ni2o+j
EtPCVOrjNZngJ2B04th4FFYH3H/lmFU/UCpE3QB0/556Qbq4ClSdZiTl579/uyfT
Wp0Q433+btx9GS9clHowZpTSXVsa0EVqE189BN4ee06oreKXz7q3/tw6w6Y/i0O7
gQS4uS6cSuR0evtv7wH7O/lXZJrGcOzsVdZxgOPk7ISuhF8EBQKuMQFv74MQtg9Y
kg+74aPwXVtqyqhI+v3aDKQd2B115ATNgrsVT+yP9l4Cg88lKCSr0TCuoGSYiE0t
ZNhWJd/94X3D55GeY5qVtFfcos67YdZXq330r8aYIWO5o29eW9Xy0K94p4gYzx2F
9b68n/uR5covZFS5/ySclZqUqFSnJDV+g9Z3bld8CsGnw8gLUSM50AdbiBwoqgsR
u36lqa2uIt4ZCxkxLvQiPAM0md57IxCthDlWtPv040S4BrK9IjNyby89Ajq4uZSk
ElfRGfHMQlpQ6yZPDGLtl3UyKn4hZ4kVsxdaHfcOKfLPkLmF+tbHwmUxpekIfs4j
xvsgTCrZmt8BrXzLA/lGo0brcP/gq4j+aycxgaY66gYzD+8FpcEmhW+IVUaJpFpp
hLYQPo6VnljAXyIa5BMDJFc09o/glHmPq8GJO9XJN9pUsX0R4sUmzMSmypqLMZql
aM5jXBDKfpiOSn9VzVYdgHnKmKjpsNTB0M9/okK4ZO3C2fyvnoDHJFYjC/DTKEdD
xyRvJTNpOI4K7xxoyg4dJUcpn4Pcdo/y4z4wLWeLXG1WsCmu1I6lobNnosDc7aHR
qBgSkefayS6/7+luFyY7Fpk7PLCBCPo9hmH0M50T7hGsKEG5MOZ4wS/3u3go4SCB
AQsaz01ZMSBiTpeL1Hqm4H03KsEsHFDAAYvndRbsiXc9FovKuZ2Eseof0wwXwS07
TOdaMZCGt6uZNAUQxifKd/txrXaMCMEFhutUFTLPROnILkbehxqNG8sWIz+KQ3e4
99tSMNhRFf8QogjB7Bd/WxwtX5uCqnHm1HblUwjoG57oBBl41YGmtPnKl4m47Y83
Oz3YFT/ympJVF7ZH/Ezlyo0Y6PlfdggwRRlyjzB3bd/1wSIY3Yp9GEu1CYnMy9vu
OnE3wCAQGYoUpcCmhfr0rnZoZ718ZaCO5kDsBKv8UP//vh1J/NZixDY1XOWTnUM6
uA/vOYtcEGYCKGVa+FcCro7Xrj+3bU4Jj0NyzF2VoMWZFUR9+MthSINqW3/KT/uU
KWtlQUei/ixJTopYwZ1ejTKXpp1kNyo8O2YRsX3hhGfW1EsKXJNul5Y14Y0h2M9e
4/mAb23dHYBmePsR23toJUPXrvLjUQQyfBNUnVF3jMXv0Gx61FbtjrNHeKy+5037
Jc+kDxTiXRjBjZqUn2D+4MWQgV/A6jvfYM+S1gqn6GOKQRsomRCr9uEZq/wNYcph
WlGJ3SsN1BlFbS1nS17yP1YuWojOLjKUXviFnSF9uw13uH1AZ13z4hCWfF3yuGAM
exDp/s5gU8Y4gOhPUqAnJH+6O+Jx2NRLiiVPIxgmqGuvp+FEwS5YelexqWQ6hGWk
EaqbtBPMf5TxTogRpq3T3hhvnY+qOuwFAdf1opP/AK83624tkxus1Qi3+MZixaLw
i4bN7u4n1L3fEw5TXD0S4FjEUSbzNjZ9apiwjJ9qJwUKsqi/BuOcSvBUizmfND7T
7SjnP/9cSp3aFWZseYvVP7a6xpZaQNRPde7SG80bo2rFR2Jiu4itoqCWLM+UgbWc
e6bLpEprKVTM2sM05jrN6pJ3KAbgkNqVIOk4eAoslOVOr4A8E2ve/sOfbBJXuSb1
oH7TqzKgTKuamMHc5VdVnsuPSXB+SypU/X4ovuifonkBDeOubuV4TfpB4Ll/Tt1m
I8fPPz+MVwjkbYoqsETsw7JIEhN0szOwMqg5XyyWrM/r8iO1JH0SeEx4Y+Dx2jjl
41q57xdNum82O8jCfg963pqwWhMXyR5Xvke/thK6e7hrJ2c+noxkl1D2X5DCdoSu
3t7wQc184CuPKQPOMti/7Qeq75WNmFpdyCd9utItwsU3schioGJz5gy7zKRP4jsa
EWQ8mAfEyFib1O2Ac6W43/U+iRzfeZRwo1L/pvQPX1W2EGuApXe/JUQrpTPNsM+j
RpiFmT6IECv4hcDcjYQOr5C6X8njLXoIt0HoEUtdegrr8zaciWxXJTQzta6hyXXm
ENMo35PrgzS+vPkU75Ng0V1f5V/BuoUKDzj5noH0FQMiwWoSh7r0n8YV2PfLsMYO
8j+EK2uHf4ar/HvQrXY9UkTMWFcH5yi9wBv1BNIlN/76DGSlTaPOXVbfO7CDXXDi
FY325c0LLLfSAyrW6+qTUksLv9nqIBs5RWRYMyiailQHsrTON+UuNUOA7ac1epUG
bGWLd+hEAMG7zo5utEFrLh/hRwc+ESRAOm1+3AdfuDVkbiAMuZlQcSMUZhg/Ahwx
eXJW+fUm+QErvNUj0ZYe/2UA62E8Odwo5LtZcHOeTPNQuXI5lEUZApk6htwpRo3o
bTIcR6FUscqWqFGIDAt+a7TJ062bfZkGKl5N5I/RM8Xnv88MlkqUBmeOl2/MvVM9
O77/FdnQ/lcR9DlUxa+f6UtCVm2Om3fKO2KrfzsP5gNrsog5E6FHrL17nj+qXXt7
LMqBI4vlIFZc7WEu4th3AVv/WwNPuJEsOrYxEuMQq2W/pEqPZzye39OYKMZxsSYY
GXaU3sG8eaeRv58860bPuAER59SRHn0N3V0Igk06R+qce5K/qjWw7EyYm6pAo2+D
u3teafM7onSt5yxHW8X9Qoy0cn6Pj+MYYHNEuMGKFkXxFHV56xTlk7qW1wcMy9UR
3cNz6y1XB/9vZZXoiZhj2JjQCNJgW906UHQ1UQJiUdApDGDXwSr1/19c47uHyuHg
GSrcNX6PkyDvCgbRcmTOxmLHbbkr1IK5/rh0976sOJDzyi5PFJYKo1d8UWxN1UDb
E5NATJgbLSqVKD0QowT8U3qNT/V3F26rFyOOpS8gJ9Zz4pp9Ld07079Zzb+jIaV0
KiT6W+rHqYodOzlQ7hhbGW23sRKwrPAcGeMd3T2aTX0dacNyshUc8LMSbHr28iNL
JOw4nT1eNnVdCT7nAA60j2+SvAhlGDGUi4WQ7+HdzzEvTnV/krkEAyHiinXml+Cw
+rk3RHpJWvxmEak6I2iNhUev8qIfpp37a3IQPwonkCpr44ktZLmtgz6yI5qkb5tU
AnLm3ostlGcbvbohp+81Ta5y3NHA46Mn/ugqUONbfTsOSiPliAZnxEqN/cgetknW
U3n2FKGmWGlM+OsIJR+BClWoIxedm3bLj5lNK7YMNFPJ6Jr5kXPGbJHRiekhNKJa
b66XDAEVlzqISoG2kT2CRe9dnpVNuXa+kPP2rlj19jH4rpcIi8hMn9W/ZYd3PuVa
qYjnPxO/MUYbiSq5D09yCNMl3WH8jztZMv8HYcdy8aEzNmFI7zISSatgIl5J08we
JWLIVm17eWTn6BMuworq58XLnhN5KN5UuEOJC51WCCPg2OWfGgnbhAiWWEFt09av
pxfluL7hTZhQJzt+8vs1FrNjiBAK5V0gUux4Xfs8fH9ILtCi0Qgm1R2DK+hzMCKN
mO7fm5rZyOg/LPkioej32p3suzwcTGlx82DA98SUPGt5GZDL9PMKJB3WnoNuYpFD
bCKRsMszoQIGqEBeNRwpS05Gz1e4K69RURA6WhHXnjOh7eNmeC08UkukoH8dYegI
NdSnojI9Gr4waNNznI+4jTnY1Qa/Gs5X468ZwyLT9Epr8Kf+5dMIo8ddaA13uBMJ
a06aBmHSdCwEAoCZUD9yWVvHD5yD99b4CjyUD0hIH7PyFvF6Fh11NLsJEyOI9PFJ
2OWQN065kK6LTr4rGQTT4IF92qzlOsRd4aU1dMt6tNhYPcM+m/viBimMpZi5Ur2o
iT0+BC5WFSBM2/h2KUuXAfWcKXOk0N1SbHrUAJJ5dAGJUsHM+zr0JyP1iifqSWZM
i0RyCsbrErV1AIW/YKTYBvTDoLG/zjJGfdTcl+vvPIptmJ0UHh9glxhK+DWg9Sid
aTcF8KZoFtKofILqRPJYLq73TRqFgBDiAguvIlv4JyDQVv8F1yPWuO4oo/Nkrxt+
yCRjkJN/om41xm8gjSz4yfqb5uYhr2DNG+vyxL2uYisp2DPyk8eYYhc2HbWPMfle
yEsgqPMOyskFuUdY7lKZrj7LxcLLzH5ff7vaAT0eVg8ZiJMZf+T4WcfMtTZnNEd+
g/bH3qU1g0YchWmEIPusWGXe0PlK+bR7MtOnRH/RsTyPESkSlfN+F4OivAfbOhqn
HQLJkby+NXvblhq0KCBdvtlsGYaRG+0Yd1eQEPC0qgDqOw2tPIc/oOj+vO90bfbA
BavRDSYMFk4KPaKGgQwX+MH0QC2kUt542krbn4wKHH7l40mDa37E8+USG587cOWB
PG03TQY1Rl/CH1/yKxeid3n61lggoJMLItM5ALBs/9llOGhVNXl4tvzi1+8hU5UJ
ocVD4f91WNZq1ps3cBNaRjF7CtO+NsUmQ0NCJ2rCTUwnfxeHpeY/HpeBvWVA182B
XxNAI7TufpPzdkHairwo2r8fYtbI9VlII/7T5208NlYYQR9W6SS3pcnijQeXaqgz
Lpq2VSrmBAPpuXO2jPfc3JLwL5M2jy87IPJW8hnAnYq2EbTteYGPXKtgSLs5oNSi
FVd5yHPYpsozC0CUaXKPXlNwGPb26Mh/YO64w7Ogy4ouBp0Z8QPGNViWP9jrw+55
uPrOgi1gAFYN0Fct1GNx/WYEgDsFdMngGuIexM+I09QA4BBVq3DmT9v4B6xG+Rnz
AInSjJDLF8vD7t9cX9UCLAAm5V0fff2Z1JFn3XL5Osgbsu43M1CyzkumfQi4eqip
EHDG4nDsYgPdavHHLQg1MaF8AY8Tl6Uezd4HdFFfuUpKG8HxIFFfd/FAElmMnx0G
ujwiX2ljdIX8qmR55JgmMyay/zsXKpIZwHW6SktiIuyULebuKg385/pBcpBtJfSH
n3NfwL8Lsl9sS3/AeZshNvMNxccY3/1cbaRD+y1i8+ooyHfiiOGJ+cPB64HaVdV2
BZkkQglNk2So5RKQJb2tTFd3FyjsOOTtX0a6G9xVtUBzQlXoGJ3clH9jYPgdkDMU
0G7eVXS08e8V1TBnhlJEeviNAMzXW9W4HX6lBLV0P7soWRg4kirLrbpcEK45VZvh
JdrZyMHNtsgm6YNuyLgf8CI570ax8p+fv70Ynq1JjoprQFG9u+YZYEnKsazLabT2
3AVGuE4YdiSG7A5fj8H9OTGmDQZo7ywxQad+yJx+QUQqi/HbjNKRMUmxvUfJX6de
QQwsswU5I0+++5oqbIlX1H/NoSse5bOwtr9nCnYaU4Dq95pMxMA7QVeHGiVpU9aQ
L6fR5n26DM/ilGw/IwE203uOFoya44SkD6CLYB6NEbrQXW+q7ZKWX3VjtHs6TWyJ
HFkAYUu42IL4ho5z3AJJCkQsi4mE9MLZNilH/AX18bHnpQSJuE+/3lzAv4iWTArn
nDlvpdv43MmrR1b3jrn9Nc8d0cDI+KyZJT7rXMuNcBtszRCtDyfMkYchcLFTt2mv
RiApuUnNAJ+rufM87qpeQ1aAACrDtA51YU81UaudfGpkvoN40qyqUcDAMcnh9DBR
CfN797PhFe2J6yyubSF0gJm6gNIUpRClFlD40K+wOJTyILlKRCN0UI8zV73LWyXK
NOzM6nsCDNGdNZVMIWuHvgWcn8uYrGX35Cxqx5UjBphBxPMtmjBoubwseOMmKg4Y
WSV0cKGkMlij2AKq1zXvAbrdXaWG57D3jfDjJEHejbPHWfuQeifuXe6E+WRbwdpK
eY4MTfTX5hx0ucBoflBY78te0ZLUciyjaBCdJW76ajastGTcxBwyQ4yA23u3UZMa
9XtyFk5fd+8sm9Q7+JYZNW1Z6NtjiCzu0X6T9kGS6XodmxvrBz6vXwXdufFTyu/q
eujxH/ULqhQmb6URqUY9yfxASFYf5NxZ/l76l5oYE0B8aOupGRUD3fHPvXOrcw2V
y2JhL59fIBXuXH0ucM2PQglUWmlifv4+wEBXGBhFXgU2SfTbz+0RQKmy/tE2gL66
u3GWB41P90k7NAjbHc/YskdGIW3RjLy++z8tDsWLh2SKoWwSSVEH8sEmIg5rj3id
ICx0yN6mUYEMfZ7Zn6y9Qkln4u8k7y+UuC8wesYmXXzubYSQ4lmRI+7WFTaDycwb
RA1CJ3tcMAYktH3LWX8Lf0oZ3vSFVVUXz1mLfA2hjtuReOy6K/yhb+PELK7c229v
3z+gPG2sZzROSxbamd0Jdgcx5YIt8B4pyPZgouKoOOXdkNVoX7X8c7yj72AcQC8v
K2/ooosOYS3khlQ3L2hPd2ripmKCqrWIwaMwulfE3Mz4LklnCqSotCCkQoH3AIKz
bpRkjJPOZVzAWQaayAndyryjJ2NxLc0rRbaohj8q0RPG/zW3WuRwbD30nL1qz8RC
BPkkEj0igFnQN3naeuRlM2mVuEG/w1hQSiOi+w3SD+dZIA4tbem4SuiDGDBcUVl+
kjLmIyIWf8TyCXCuGvI2Qt9uNcVslNNgE1vB6EdxGDdyZl/PY/jrvpfjS52w82QH
y3qq/3VvFXO82zVi+idkGc2ESjcmgTvDZQCD80KKo/+5ZgdzUcgbwRHmpgrII+o+
avXipCA702k9V5NJpbmemnIKrSBWuLeKmmixVmu8Qtfr2qFY8TwsO+Pw2zUZYJZa
K/fC48SUWt8ONFqBJnTnQTZSF2rh9w2EgzR3pxSEOoRSOHbJMUj1S/y0Ud1YOjZT
8grrmRuc4aLHQD/VYIhOO53CaRveTZENzIFsGL1PGptEIA1/oR2KklEZihTZXqbW
URpR/n3iGKkocFFdCuUpStHMxT8iq4LHSKBjWpszMPimRv8LzoUPf+SUbRAEW11H
OUnkbn5AnOhoJFh5+KrYoA6KmNxbQZbG1RBPiBzX7CwzF6oLbeew+nzDT5HEpfeP
vudjWimVrJhFKkxouKpUaZPPeuA3Gk5og0g3zz+jn1I6BZuchmHAMs7NdTh1JtP7
1//KkBqHml2SuquUXQJlTTYt3OrJsswQ5l5eWNzHFen5us9/K0DyU2DLDIi4nf5N
PLHQcaOk3DTi48yksPAhdNck75RTAUCPZBiZ0JE/CcLBauF7WAChv3cCW7871NJf
2hvbx41gG3fNjTBPfYrYxVdeKMDnX3E9eCdzCjuaQTX35Ymhv/VCdjjMRoFxdvsM
NPB1xB91q/hx/gblX/nDG6WwgqQ7hDhUBhpDXXIUxMZjfj2oyNQftaLW+ylMTqaN
+M11gAPSz1/rb65ZR05txNnyJX3uttnwAr4kTz7HV34YdsVjBFMvf/guiAet6eRm
VYzUhdrn4XNB3y+0oVMUJ/pm34vaSZiF8oCrDEw0ikF/rHne6X4rW958HVMm4rfj
rZWUGAqRXG075Sp7bEqG7GEXUFiWxYtBzIYlteFMjx2/f7UUxUXaIGkv+MgcY0SG
fQSFkEpF9pfcJVh8eNuvxbTrxY+ePzJCxGWxhoCr3JAjVBqCZagz7+0IvnBhrzQX
T/LhTLMKX1HJLa0CFcEAWDPlVJENJu0OOXCRDavxMQlBKp4IcRHM6AKYC5PGmnK2
yewbn4i2B0hHfFK6tCx9LhB3bjo0kxtUsBva8VlV/9RNAZ3EWucRr2120A/5l5Ef
O0ycEqwOisjqnIzKvr3zK/XGXOmT4aUiWWu29JL7YkYLVK59/9l8FoMvjl/gS8nw
4VsH2XWNwTpGcc/U/6AcSnDFYfnbtA4Wa1Dlr+VcfZCqOFhnLbyZ4pW9Rt97+xcy
jv/zDJqq0GEZRlYiUOxBRFe/rWfR1dFVUrQItWFCufjIg3jqMHo4npNI8CJD4Vvx
yDn7wvN/X+dzwe6lV7Rg3vww+ymdMBgbkM9isbGZhvOn913Sc/BOuhig6m0/4wAL
z+SNpKCQxlh6IzwGy8xIVFRAB6ZPrG6XSP85BJhhKtE4gKW9FQkHsaMSFoG0MGg9
CDauvou9xV2Hm9ALzoIQyJ+1gVotTOxJzpGEH0z9HzJV7y7X7ze4urk6pM1aJtTP
bN5+9NuQAExS//G+wYKeJHGCkL1xIxZVctNJBWqeHUmZA2CnCOvCTcTbq5mELs+e
weaIBFEyocaYrfBjWXHZNx6CDyqO5FNJHu/VufpXe2xY5p9l5g2PwaJoLIjD9b82
oQXv2Va9QkVV5Xwkku4Pa4WV0d5b7fkR1vBp7lXzK3PYkDm3GdZK/kTMpjM4X5o5
woYTnQoFZP7vpuM870dfa/nZIgeyS9ijCsddj+BsxQZ31YO79IDcwfPhdUSAELY9
n451+YILbDHbHMKozdVd2CGhR4O6uKNke11mfAHT3Lu5HbV7q5QdcDO1KYOX+kPz
+Fw3EekgCnMnVy/WZirWhvv/4S2WjhwANQI22sbBihEYYbdH4FCG4CNXuWKVMIA6
xQzKtdGKIHQyE36Q2WtnLHpKA+4xOwzPuGhWKNqCPOFlMfrLDL0YD6h6CDp8BVC7
tohVDIkZqaAhory2PlAc7MRo/VGc4UUmKh8+tEby/BzaknvpQjAfcR8Ye0XnB3iU
Snb4pni8PFsEnwgeBe9TfjKw0oYXtvJILJ+Tf0P6fmdMxiUYtGjzAJ8digpUZ+7B
+QxMLNALY9a2feP3IbMoQ+rMazK65UFgMobk/rVBwH0rMgawHQvjkSrYFuq0/0sB
1tDg5WvUf61vo2QmWxs8SluRDOWhKoCHKu0tBQNUnACNJJ6RutwCJB53PkawDtV7
8oV4woBBfVyEenS2ssp6Hez3KoM3qqbePbv4UCrRVHcSEYNhw7oDUkXQcshadrnR
CB6m0Rhx08ScnOtkXlfJrR4NzjrfSQfyWID+6jEHzZD33wyqUodPqYIVZCYBA/H8
DbYqLKecYHmC6mEE5fPPhOoaKs6x51og7018DqHWx3XJ8JQk6I5JZuE3wqYef5j1
5sHpIogGKdZaCPKoxZVCpcBQhaOQqZpINEddAdJEWzhSXT3703a2ry+3OzLMD9jP
i0UfqHIX7WZWTiKhMphsXqVkHNzniuPDRjIaW3xcW65zCH+iSgHVNf7ybhtX97Jn
KyEvEDUS8bcFV1jiuEcE4Da8/Myinb5ueXg/u5Gyw9uE9wOA0l8kuBTmd+pQodmN
IaakCPBqGIDRPf6Pj6OR7wxfflnQ2ewYeVrbVm6/bZzq9lNQidDmutqkRNMrF5Ft
+Ob4fKFa6vVYIPyZKdwEFjyhgVwQtLocYCFDdZ3qyDSx7XWSCnr2KaWvLW50valM
sW8dISZJzQC8hvDLDkZf9lfDYRfgNhzdZwyC8J/NaUt4AyLvGH6XuGKBt+cn7zZ7
+wigfKMOx4TJsdxdyRilFXHH769xYKvSijQD8gs9y+zWohblrAHYhhLXag1byhzj
LSnhiIZ3H3n/VXZ5j5msR8pYFW1ho25uIUrMBZIVIcH+BNCr0KvLDbO/AwikG9P6
mlwat4RfEDicenpLQSp43IdqneBs1yg19FnHbKiSmeEDcKHp3DHQYjLaNxw4Bvhq
meImSX2TsizOvWp45TRFhacQL3ERWJfa/+VovwUgj12gHuk5sG8sOVX9XDHz253S
pjRarntGXKlv5mUrzS9JWh4QdaXH8ERqC3WFi9YKAbM9zvkOLb/kesYY3Nr1+O2C
fVjRqYNVhnR88ED3aMdZD7Y18gJ7NtK+DVY9xG7vrWovM3XpBbXoIr3BMw1TXV4v
wMjLOQMxuPbJgWwW/wSgqzxYe3X1goYCv2rd3u3IyGIqCxmxTx6zzAEnuALjoCsz
abZ0dq4MSXP9XlCB2jIkxBYPgE2YbfkfT80lGZER7Q9SsCt8pefWplmj4B0rAulZ
lzITV7bvTlQE1ur4TM9BqUYQdY/4oSToTRjLqURqwedxWjKMutg97K/YUAYGLrg3
sFlsb6AizO7d7O5DUXHK1EkjlcQR1PiZxfNC+UHbqL/7hjP+OSDlfI52Xdf1LjnM
LQlR18FRUy9HVFfsktXGKR0Yi5Zl8JqXgVyPTyKjr+RDOQXRHAgU+C1ZitwuKlWh
NSqqz08K5ierSLc75tB2tcYVmITvB6cOf7VF8JMu1C9nzwavV9TguUbGHl6AuSyD
3/ZTy2TroPL69ekytUfU0J+qPxNwTRLbHbNocUy8hN5p32ggKBSID+BXgWqQLmDw
dChdtfakiejUiX22KI0DICC1xazJ8LVKS4lO5eGRlBaDJbN4zH/CmVPZnt2qODEj
Ya6yxbqJFagDfB/AhogyEOdjBTcu972UFhttuygNcj9LmBHqLO72MDzfcxgUQWHm
cxLWrBkY1j7QtVNoAFNwfaUwfYb8yZhON8jRCpjqbXV65LEepMCHaRwOJ3UFfk8n
F01uGCfeYXL8MUa6rTHvU/4KCRvX6yor/OI6GZh5CqXe4di+tFSuu8cILA1bhDr/
jyQRGRjW+Nc4C0DJyU6g1mwwE/I3jajDpj3BBNN1nrZKdlLy9bcQjdDKIPoaHfj3
7i9594uXzwenBzeXxkonvIMw51LQ15UhdtkOXddEl8OG9V/CuGmNbqvTaoVMya4E
UiaW16iVboKsmvZLlbuHV9ziOe56SLYQmmEh9bu2ss1VAH0bBicSSyQbEwOz7M8k
UMkavPzPUPdIoLaIPgO/Cm8fkb5veVqQfYFzNwPkovncarKk9d/pyc2k0gtXrmQt
HKlzjRr4g6N34xn57BtCNfv7GzlLPlNZpYFCp2jAV8UZAB4hLYy5QxZJ06WJT47I
T/I9AV+LAmIz9l0DxSNfz+jj4wVXTuXEhrSERyp7KXQZiGS33kC9gNoteM0uw2TH
uivDewNrA9jmnOjSLnb1seEFn7J0L4uv/WqtCnRdtjGPnNxsZWkdNfRv0y/+Wdao
ocdNEOFKkMhM7s/jSIs/sXsyDE9XeH9LjE48/i9b3Lrd7+7vsRROyq4BSKVn5UaN
J71iEpdLRmMokT2Rn+jUlRazTn7Wb6UgHYLlrwXlpmOA47zB3wi9dO5xmvY9Hu4N
/xAdsG3TlkDDzz3LP283/Yq4Tv+J3G32FL8qJKqhqoObFvEL62EvjNzNZRbNh3sX
GltaoNhfCK8DyZIkrJ499lcsvtx0o0BLExddR0FtLBKV1ITuLn2ByHTrY/rhWPYD
6bkVkpLTA9pdivDhYtG+w1e0oC8dEiMGpcUIaeEu7GHMnjfR794etz6+IWKE2tJr
2Fl/6iMef+IelpBgBchf8FiPt615II82EKEEsz028fr8+diWnSVZVXq0lNzjgPEU
uFURI2n5+La/cVmLL3dwutBZWaWc5Qnl5cfSWSOFoRMARreIB1pJfQxrEgQqSp9b
5186JtPgalKkF0/p/mudbubjOUEzWZGnWm6VAh8LelBlOD2Pi0YWwyXj+rLNBN5i
a7eFD5m/JMptn/nCfCsZxPYD2PmGfmHLH1kTZVg0LaZ4U3EVnZlB4NocTCkxO9Dd
XCvb3wA1nywMEd5okVQ6XEqppuWkVsalRuCrKYiaF7i0PEsbFHqmNi2gGI8Y9n0e
FQi+wLI/b7fC3cHfMGgOFVDvCouBdNJlDrIQBlyLuJn/VFmNFgse0HAZMxMxjKm2
rOW0yoe4XjDwhAOwFZlg8QDsHE/HFX6MN291kLsFQT+39DvTYQd0WKXis1SHp/fD
lRCUnnOS+kcgf5bZ43Uw5Oh2c70cISw8DjWa+3XFTQZDv2/gHAC4DeH373i3cJsr
JccatAuiESHc0NITZ7bIPvHB7g40h3yG0LnY4nwRvQIvrcmlv0b20OPJrsrrIPVF
XFGF40e5noEf5rPMpTv8C8LPph2CrmeaD/5NcaLO/EobuwSw2fll0xFUKYTn4a2s
JN0PtBWlB18GlZ1ZxoBQAriimGXeRUyqm5b04sdWAwUDtr/r+U723RVGCvol+pIY
rXlnRackPSK2/9agItIyAJGMgzdGD15/1TrAi8nky4HONbrXIDKCTB4fkQf8uvWa
3ptspumz20vvZSOEyipTspZd0S1LEAAVLoT4EBTIqfuWPAr6rJiTWKZKNOf4NFmG
lOr0V2uHgmi0Gk0G7mJvTD/kTZ4Dq/CLYYW5vTh3PV9H/it/2wIGRejYmC/Ng/zQ
wo+o7WxSEmAlyw5fqtEGM26E7btczJz3bC+VogpjKc+XXnU8nR+9bc+tgawOlE7Z
Bkh0X56A6XMXEr8yivLqOhXrdcjnOQO7tPaj4L9ToD1LT5yGWniRXbDKsLTTE64r
4x6rezIvHOjt9oSX15C7Kk+/jXZawojCRjSMlVVptmJmocYYK/sU8JhEilOoTnVg
gtuJiDg/ToEz+kXOD7r1xsB6G0ELIO7KGohvE7rRJBszmKYSrfrO6L+6bUbWjAG2
rBdt6PTSjAbu70uv1PnZMHwqJfyePthd6kf1WkmHPPDvSyNcgYcVHwKpPjTJvsj9
/s6pIS78CMH0Lm5m/Q6NUJbFbst11z3vxb9hqBDNQoJOtIIgcux/fcciLvG0/54n
3szylSm5ZQHTBFF8j0L9ul3ujwfUmYLBEDTuY9GYfuTZbFObNoywYgt1FJFXvnD3
nqI0C8vpRz32HALKOKgolxG4ihdnyUQFKkHCsLCCK9kWj8DKbxwvhqzMCHq3qa5z
d7DQYGkCEkAIpfVJF0VW2p9Dx7tGzzOodwdMcx3MniNqIrtQeUi50MN66fd3NN6P
BZ3FkpcJ3Cfm6ZWktGB+y+MG5Qc/Rk/b1Lypo47B+zMUYDWklhtfC4wSDlRxyxEI
RiFHm0h3uqngH+On1K9YtiBjze7UpWcppkssUUOr+z2yPGG/PMF4WMMfGXE3iFM5
uq/7Xb2inX/IBgg8UZG1mA+Qe7vi7v6FGxR1nPfm2Yjg+9NBcUntDwEcfRtnzoWN
LXplfLh+GnJCjzSdF+a/iQxtlf2WYaUobaT9WW6Sj5h8uONYXEqEsodUIUZbq5U5
RgqC/iCgT4nuQ9v5At32p3pgg4LDGYIxo21M2umJSBHPkmHD6/6cR0iWVaXvr4yV
xuyEp5SlkPhGoRFdZ1GgFh72sWJKcYXtHlG4k+qM/r+/rChyY5tOUtSNgB29BCv9
/RSOXTv8GY1mXO4P9Bzgtzhpuzuq656NrGnlNSqCOwZ7uab2MbYYIbQLS+GwnFo+
89zWDosMZ8mwx2ulDWC2X8abD+iRyLyIxcShEoeC5tvC++uXAjEWowTrpBZurY4O
phgctNyDm8I5eXM+Mx4D5uej+ere1j9Uy++DUn2WTpK7V+j/M3g0gjxZwyz5RC7g
GdJKpw0DFKcKyVzv0NlZ14wL6JnimuoVxWcXxuYdyuFyJ0+uoeommbexlpqZ/rev
tYoE2CH+JKr4Bvl62itTgoFnCG8qanQYtXnTP+PL/9CccMBYg+EtbamkWslSTWjt
27BiH9aNeJqvmYXA7zPG5bpyXDP9t/d4BEmUxH67/XoAY5AZS2oQrXov66dPLsHP
0h5EbctsR4SYVBKtS4Ctuzx6TJBbIxh9y9nq18DSbi+BXfkywFWb/KYeL5dIK9tp
DuS5+qLCGWy0t7Zu5hgcPZuYolZVcWzWbm2NxDY3cBZhHo5X3ZBXgTczibxpM4sT
vDkI1svxGMbZcz2pTzX7Zv/4n9NAdSLXQkNOMl0QoLwip+Ww0myW5xO+KMcgunvx
gQ9gnLnOw28F3YQA43/DNqUFwHw3ppRwVkEf8klFgV+uqkYlHaf/VdYgs82qvi53
bP3rObgLgANCQWSHQ5CHkD2PsXOc8Kn5YRYft98zru1F+Mrt8ZajWBDUtbLaC+Xy
9ksfK5RWr7eepX3QhMUi6532J9MxDo4t9NnMxItUG+j8UO+uYgyUA29agWtsAK3P
6U0LB8ntf8+3Tit/NF2PLxMfI4ayMEJwTXEBbcOJViusSS4ZxfLx5gudM7GX/loz
8Yd2KRWNcPPZYGJkSu2jhb1J1uv5/BjZ5L6psnp7JksfnXaug3/vFnq4b0t4ggNK
KlBt2Pmm5idaLj6blB3yqhnyC7uIq6NPdXvK9QNTOygWAk4JNGYCGo8EHHSfXLpu
tIeiKdsyUh8+k1m96yfOO/dY9L3rpwGyrbBYZASq/xwjln3y33SF/62ZICeQ/BVQ
mT6utIwO2394DSowRjGCuxtzgXvcN0epP6P6FLYVjK8GoFr7FSsey31lVzD6Nc8N
+sk/Zq6BCKtPP7lY86655C8+TrOVI1w+mf5+XGynarxXRzk3Nq2jlrCks/w50kPx
L8xJKMikK5Ux7BC3c88o0Fier0CbvVukGcefSGwUd3jgtazJZ6PWAsOZaqxrgDPr
OwmnRxcHiUUlmZZt2A9PYiJeUKMpCv2iqGVEK2d3XDbnQR+VqbS2tLFOj+Aowwri
xTg4dRKjOYDsyucYuH4ytPUR2RfdhJCH3E3Gkwc4YTWCWYx44uDBS7EksdEW8kAZ
qahKbqgqAVRlc+0GAq59ah5HjYVCWyKhyAF4P0o7C3gEnwbgStD0Y5dC5Wstuqo1
ahXYoaDzNXJT3jeSnGeesLHDPCj4lGT1LNxnqi2VPI92qvFUU8rBYLLmjjn33K7b
jfeDHqyYhTmIJ3ViEVkIFNXr7pMwPqOkZRvjfKItjVeIkyYuHaYlUf01M5+eLTqv
PpyPKkmXGqVUmj2d9ALTMYOvT6OJLsTLRz04MVFZDq2pi1h7Y2n1bY47sUxEdVcf
eH/F0odCkowKTmA/qLrdW+e6vLNzIG7ehLqNdIDBbldkJK+iwgohy2OgdEmqdh4E
vnoy7nh1c5ErBrAHn4ZCIDHyJ73blg34jd5BFhPAzBDW0X/xRdhT5BDjwZcEqBb5
SsDNQtULFTs/c0sMtcN+zPbucWSd4wHxiwhSCGpBJaFpuTxk73Gl2p20pDiDIvSL
trSpSC8yC6canJMxVHiNWxFXv1qFzVPTPsxQakhYET41+nd3hDBwFWozzy9cv1CQ
LvlLm/RgR1EiNRnuw+5uWJQ4o+TgTP6gG3RBGRz05HnklNj564Bus8In0lBBkA3K
UO0Lt2iu7yCHlwrl5wGMvhZ8VKQbWQC8dBBp8+fn9wpRXRMTXCckZtMto22ZLXaV
c/x5WRjgaEVU/zdAIZyobHcNR82C3axy4fM/Fd26TXyU/MyykvgoUugp9ZRXlT81
ux9SObfcEY5zgccLw7pJTZkqoUpraHKPuLMfY2QbveSEdFL+5UgNV+xALAtZbngU
Q363tvFRP0rZIGJCBHKGEPTkfWWAVoNUjWgcRZIha+z19D3YD27hUvRkl6aOausP
Phn0PDoA2QG9yjchRkjyXN9ELhlDpYFeVC9UAu0sKtVYjhsfcLvCp75dlgy3y+yG
/ScbxtONWO5mS/5SWG4TlL7hO1vHnoyHNqS5LvIV30eF+dT4+Q/BgVa0TSlnDlza
9zC0ENTXy6QlK32rsd3zJouIntaN27VYaztcxWkxIpzpMysGxaxU5DP07muzwfbl
WPGE6WyVKCmKUldXTWWVmb64wDpbIIdSlgZ0h1QjRouIyXLz8/ATGeOhgHWUYt15
526kMew5epUtnY4iDrFIj2SBMU2GX4ft7LwS4TM2JUAKoIptmDDR4iOXU1L4HS3q
qwnk+t1Ssel8IYHiZunj+raDgOZvAlV1+yEQmEUFjeK7jeCJ8e5nGZjzVwrHnQN1
ppyQLajwH1UnesG5c/3e6FTE5NRCVd0o1h9Mt7VtcDflciI7zha1wDRCZKU3zGmA
lV1zYSDE472ooSNqYXkd/FZ27HqqbWGFRQhPB0N+zYJiJL+T83sVVAZ6i+q3JfGB
ZMJX38TR5YGi1lvWMB2sfh3aS6DvkHDtgi4VwaAagujK5zblh/OwGuQw+XU2Jw+r
jUCurgVhrSGfAvUNfwp7yHZAzPxEjYLsxXUYZ6jfFWAS3e7sxuqZdxXR5dt0Cn5z
g3DA2NiaMcvPefccBBVuJd/PVyRNDlsslvH0Xicp+IykP5U0/gqOuF3WokCjF/RQ
7lye5MwFotQHO68ck1/bcuAKqxSJ+kjPW+hLqpVbV2mF+eFTa6PkAUW7Kh0x2zOJ
DzHc8EyiTlVYiaMjc5wKGdoYnbxbsypuMn2lv1u8Bnd8whA387lt/M42tQTPNV3k
lLRHW5maYj7QtAGSqW0a3IF0U57ODl2D30VFDbJaOabn7VgS4PLqQuasL/ROAatD
pCgT1s2KtXTg6ocd4/QWZbBDoirJvUOXQsNOz8dOSNzfvqkeGkBVP7VE2bT2rmBb
toJK0QLrgPtN+OAkulwv08Spspcz8kHBVMnyfPQXFwIE9SW+Io4OlvJCEuh+2wo7
HKwBSl7wNp/LO2Ay2qnfK7K95hBDMXzAFjHWTbs3HjdEqDZUoMLerXjaRHI53T2G
c1N460naupPUf8a37t5+kLynM7u3Lo00gWdy+NDOZxJ07ON/XPkLCznbhNTLic/q
DTKSdePPV1niZ1o2+QGGQY8ZUWG9HN1VzjdWRbsyyeFDjyKdef9Vcbw1YJxzcnwY
223vkN7IGJckcdmS/b12K25CQ/EN6tPYyj3+pmr4qAz3wpdKIeUJ/1nWA3Zmer2C
K+3Pqc+TxdqboLfgPJwZNU6rn8YJ1gwyoTqmV5D4H8gGflRiBBEMC11CTiqNIZF7
R+tve8rFhI6N7TrrKbyLs7AbIJfS33QV7uuLCrQBPBkdC+iFQG5qvLiK0BMTuFDI
rjLnuTXDdypLfkYncC9KegqQ1OEnzW+u0duqwKwAvwa+OtPbEW6sFngJWZAp17pc
G6EHlGk7SD0BmMn9zpWl2KS+51S2iNBustjJTU3o7ffZw+wbHOAbgG3dMaHcyS9K
8hM9z6+GImw+bX5U8P1yqNKHyF7bOf9mex+Lydn6qRBjC9HV64lkCMsGW6esuGAc
e0JEKVbvppAdKW69iwnNee2W4599ZQPG9cjwDv8YwWY3do2GyicSMTjeRRWIXJNm
3ay9bQEL6MKITkdQLJ+98jGdfioN6a9A13lL2BJzXXvEhYrfxebPJwQsMIrXOu//
F94sl1Tw/1ccyk5kldjfaozBFgoK9Xouq0zuKvG39f637YgLIMc8y2I6TbuZ1OHz
jPcQ5RMXgnm2CAvUDM4arxJ+5MDlQRcs0mt1xufoxFkQeoxm3+56L5uZP0IPoMW1
olmoqGo3m+Q1PpA6xGKM54qFXJEZWCsZOLgl2khY3mIvH7w0xOuB9gIgT2q6ZV6d
JIbOb5Ng41c2vS+/dLTFbYdVHL1N8QVKUK/LlfA/IYRRch4oHtFm1VKThFJl6H5a
b3wVbO6oQRtzzW1nOHVEW9nGPkpXRT3zJnu3dqgVaIi+mDf5rcrt1Rax7tYjvmU6
sbCsQ7YKHhBu7xCRqM/ZAJ6yYLQ2KJNOOuMbK/euV0qHpRHaLv/yd4zzpzKU6bnT
hd2aZ1reFlYCNJS8R56pW2rLdtEn7k49X9ebFsp6J8jaIsGZpxDIqNuIq6Fhe+I6
klakZCWrFDBoSu0Q9WsFwHzFDWG95FvNPxEN7ZPemvliMKypHLBcsH1B2ceM0/Uk
BzBql9SxKJ8SbQeVvkAmXVuppoSrj7Mn5ha+RdHjmhIDsROz7kELAHLmTOM1TUD3
XVCrtv0kjFHCVzEOBV6XTNjRQn0KUz+VgkvNRk4abgiXF5I8S/NUZkPSmKZiLlQ0
K6lqpHcNctW14Lai6m7ecI6pHzbnBya6fOSgfRRDw6fU2l2TuCzAYbMYit9pHDpj
3UloXEpwzeG1Kc9c1j0+9PFI2rsLZzK7nz6vF8AJJdaHaMEdMfDf5YcfVGB2xK1L
9r6YSbKUGhF9B1TJo4AZEPY5Yt7mw1kl7nOfCD9E45rUI6IwjF050JWfEgBNHiOU
sNLhODwdpu9EciJJRg0zkQ4viFTMXxL7misN1V4jG70p/jbLF710i4C6EFa5pRoW
4OUHRAIoQ2fxKZ1ZgFmPVCH/N64LRkSDvTlGyM1WzXrUx69vH1NZ2P19980DO63r
0uwBxr00zeNqxe8ugxO7JvNBWx6h3zpYn0WSQnR5+SQC1zHiN5NKa33Y9EDiJPCk
bI4ipu/SsYxXKWJLiMANw8w7ySItjK90PKta+4f3keOnto1Q7fk+ianEr/B6XNWI
zI36lY6Y8skntbCCw2g8kNZk3nlaRYIK1jGjHFINX/JnYzv3m8OGXLALUAzGekSB
0X+X1TSyf/O+9hiTEE25bwZQSEwJsG3bhHLJqjFGHDzDg0WuwfK3S9JQBuPW5nt/
NAvWqZ1hgyObF3SvU8/491u/XyXrX8N2ysVihChUqcHYiSqclux2NiNr9Dstdg+0
1BBPId9dV4Mh9jA4VCuGrJn8tqiMp7iEXIsFLEEjO2eF8oA7lrM8XkwlKq9IaIms
EEhANHHmOeVFVz/HyCEUM4WqE3tdn72C14Yclzifh/DgruSmYAr2LF/l6N37sFBI
6hPtZBO70OnK0T0IgZ98mjgg0EVtCqja9RCfCtbnpCe4sQRpHMaufNgwoBRUMTmI
O26Gg7mJakCleMa8AJxKsAIcPXmd9cjyB/0Rut2PUPxeip3C5XujkTbYfJCHd+Wh
SUp43rtRppkwjTGiC5I/juLLes0a5E8+Nl82cGHGYw9dsBG+nx7AKga/EFpi2opr
NAVevofpP85vWhkqM4815uQWYfHLvYKviVymiJK3sQCvcF3IHlwbxgD3dnyO+rok
siv581KnlAAM2qsKJ3vx6Zkw60aggt87ROnhLKlGGQu7PgFVTiBKC1swm9OASNhS
bwEcsMGUVkNvj8L9o/Y2BfOQeoCwcZyWIwIYvsLqdAdMsDDgwP1qPeuSL/gzL6aC
056074Nxz1/sYzBuoQRZ6UtiLS/s4RTRkqZdKDH3/vYU7JtyHpIZddl8GjNBRsp3
KAOKAOzizeq947GUP5bxvGzWnTv/h455tfpJYIKBPzVxP+DCvD0KTb70qyFDQYrB
clRn81BxO+azk6paJtrnGbWRzcxP4y5veTY3/JBfSh8rr6G1073kcKWBNaqT+H/r
ADjv9e2H0v4ZuHPIvQVDcsfeRk6JT2iDX+DbOorTYTCIfwvnaXiJ1dRCrPO+IQr3
JCgnLyO5/xDWPHRRKqpoJtTbnFSFkbHPmfHMXME/Alc59VEnO9+C7WmjgwL4dmR3
a4TSkkAuR7KiPO3OuHkZKdBjIwcb6X8dO/mToxlE3K7XwJlLi613uohKPIUk22m5
IIA7fa6ZZL5+vDt6YlsO5JjP3QLGSX0zn7sFCv1X8zgD4AKBQkt2vibmOE+frRfD
bMTBTd0rcLApQF7FcQo033StI8NPNIQp+BV2+cD1fHsHYTbt185UaFj4zthhLZzn
JSD6VmGwU5jzju2f5FnJJnSL7nvJHbAIQ/IVUYk5nbphC4WoMEuzkoUBXsQjvPPT
mlNU3VNZ6Awes0sFsUXZ76/Z2PndyEUqreVJEWIiFV7ejuqZ/jBCGM3EtLYOskWm
yKmy8VmaerSvvIMz4a5A6deuPPzlIx4omxSygDl/hSFEvt1e/qv6VAt/ojwcNdtb
Npg+BT3zTrd73HSbhDGDj3MbRL229pHo74vFXFYGtDyzHj48ixXh8j3BvOm1uv3e
wPzbMmPKhhAscx7AbSP4kzrbD7FmsYa0VnRYVMbGUcEIKoxFsbBNVETbjBArg6nt
W5N97ZCM1vmZvRX/UEsm54fC0xc3Hk+e8PfTbMczPNlNkfxtM7oVluhWvyDAC0z9
vl+Hnnspj3gRTYmP9QIk2LclSF2fsIWBR/NNuDS6CJTOfn8W1YjtP/7SZEXFMJ2B
isg5zuf1X8rmGiVFh2ZQW9NirfRgZHs0FUpisKQ5ABvU67W9ZWcNpy+3aSGalBSP
Xn7uBlp2Bf0H3WhnXF8xLIecZo8imObO53WCpf3Jqj/mg1I1tbBKPKu0fHWQW5Sr
xjQszhdAROOVsnJl+MpGdymoxBrddlsXTAtxeCPyPs3n3U/iWu7HmkH9k5/NW/Qm
Msadf6is0xhQttLBBRBzqOwAAXhyyXSFC/35fymjGx82M171aXhW8iQqPRT0h1Ds
X+swHVRqoVt7f4pxq/fRGY3rYmtuvT3IybhneeBpYNhGdWNKRBpNXdQo6Phq2hGc
0B29XDHxACXwnqSvsPgDsuQnLS2WjXicbEXaZTlCN+wV9BO8yRQduT/K/GAxvs91
eMOhSVVCBWNQJb4gCScslW8A1j3WwDAUuz5ojcklk5YNG5aq1IzlHqpo2upwAtVq
wIsO+UslzMvkhUYnjj+1SKW5xuXzgtcLhfjrG7souDEkbULXInZtLQhG6yJe/nls
84EXqlseXSR0QHbjqNQc2drGRukXWy+E3qY3gcQ1eJJqlB7R4pF8lG2uOvZewCQr
huLOVIO1/eb9Cc9Qi+8oB10CvW8iKX837RS8X2jigQXoOfgxXtQRge1AeKOQ8MPB
GJP1c7gIrWIyBGrG5Z8OADXP5/871rCe+5qkl14KhoGmjOV9P8B56JO1iiUC4Dob
IvHtotAehpndqjATJMKSK+3DhbcWL8XJUeAS38pmcAtnpkm57zYs4MLInjaqioLR
3vHDal/VWX2MZcctZQr9GWiCfByoXOuwzu2tfUIG5px8oikn/fmzfqEhPFwCjt8/
afnNZv1xp5k6Hu+dnz3K0cOQNvPNwjGdRl6gT/YvyBe5yx8796R7Pn/qyBcsNhB4
+hltjJ2H+4I2GicmvBEOCwmgCvjC06nHcvIwwnsQzWdjYNYDdacFmLKWtbT9bpYH
M8CXITGg3gIMlJqa/7yudU1B/D80aVebq5obICVRDawGXck6PFsJmz6lcNOLu4kh
c+ukDOoA/mDdM/gRuFA+pY6bQlPcrfjGK6NWJnoGB9hUN0JY2Sf2NG3sfkhU3oGZ
xdev9l2b7d84tA2TUdcuI7VTUfhc3ymtIVAkArDhMItMFPCCOMO+WbogRKmGE9gw
acxIee18ar60LQpJ5gWrJohNzubS2ajTopD/GagPCxbzKRhvdR9G4ZUEPuypohTg
dlchAb+YEgRb++mmdm1Wx2gj8BdZ8nqRk2dddtEam2/k0dcRHAXu47dg35v+Sbqt
AZU6L+HF5TvBZX/8m1ptyX27IirE0BkXJcaR65guZ2JwqvbBjo1ZQsi6eFoeary4
DBghjFBJ8tN4SMc6T0FgCOKll0NZo3/9YXnkZCzn7PAqR/j6FeRLjL6qHEHbSVXK
UrYKPgl9VtxisEUEj8lLZnFgrjo2x2xawSjW4eHEOl5QHEw8ua3Ud/M4HwgTTqLM
fGpuZiXIPdGM2LD6ToGFBnWZZ6wznQmOhECF5bUhZRPG9lgG03CrC8rnmD6NKYTG
IzfsSoAZlzdYEI9cnA4zwoJHrkNWFOCAfQ/oTqvVBKJVoDGKyEeBK/R+1i9lhvJ/
IgUTxZqhZ1PZU0igcaWCYmgbYNtiaMgwn7Ut5xEG9pod9JPIdHEy6HcwgvJOD/0o
ZGuQbq2JDhTx6ysoNRBQSULXtfmsX8Tq2jTIj4JRJ914jJUo/rtun5By8Eztf7OP
SO13tb79SnRxfu+OS3ZArKduw/6H7wkpuLK6PAw3JoLWf3bm62Hk8FBdWLNlwAuN
8qDCKCLYukH+ZLazh+JVSdPxfQMsP39kVG0bC1e1hjJ3GdJvsEBoQmMtCdqPo5If
Fmyf/tWlVRzkjr7ZgCa7Ta1f0x9qHUbYgYfSjv/0VQwPDBDY1aa/tdngl03tW+6M
sf/bVDsPGWeqHPYwIhqE5Rl1RarKMNYpkl+yjZP8NMHTLyseCwAiga3Aphi9rwSl
RgLjCvmaM+udhgfANrv3s3XNXvpovQeGdyrSsjl7IBFyez3DHQ20ftR8g4WRpjuD
eTFCqCRYYH5Pk7Tx3eczox162xZy0JLgmN7UX0JuvrmwoQDVzwetgt8M1zswhx9g
zngLAM9H21+2a35B1D5PEu8CGo6y5dj8uDqlHsBQpaMeT+8Z/8P8HwjVlxA5Jze6
BrCNfzK+/Ze2tjSrI/bGmxstUvckDssreZ5kWYhCU1D3FVwWxbHyhjXRVyV7Tsio
BeDsTOHIwQ30abaYrjx2RiV3ZtzV2xX6tLpp2jlynu14qCqFUMvrPFm8ndUQA6I1
XDMqSc/I7fwKqMI+s1PitT5H3Dy+aYtzQ7bglwa/Q5RmiFG7eRPdWUWtzkvuiE6B
hMKSQj5yDKPxngk55f4t/SH8qfEljXCjpBCqPvAVtyPfKvUwsfx5Ad08JDVh5rCF
hRbbBwbGtQazscAHHeMg99zADi9Sb1ZbLcHItDN2N+QDfMlDTboQMqax913kDCDb
A8AjkVxX7T2+b/XFMXHfKsSC7JZ9t0aDbczDtsPBf4O+gOYSkM2LG5VTUne6QyQa
r8/x2YLMFFwKVUdlTLdPi0+b8iHy9C2AZORxXvdQ5PpSURtd9lCE32/dcb+/dqBH
EizKBbdcdUNT9VDcsjjFAa8nYBtMyFd3oOgfNfO0o08y3UfrF0fvC4oyGx/vfvN2
sNXO0FrQd/G9P4bWVISj+6pvgG2hvVwQjv8d1IE4Dpb+hUzcMu+8x66aYsQz27qT
eKEuFIrrUsXZGjKDwEnVEDenLNkLJgbgQ7TnG9+X2tBaF0isrRflzdozc7U1OdT2
mSgWcFmYam4Q5RbzutKhy6eKWs7V8diCtaI6VSyZhL5r+2Iyt+7iidzRkCg/ZR2d
eCKqhPNToCI5rrSYnKhu1jsQK0218/zRxELxc1UTJdVi70Vu44hQ1aF5PpjAvVNE
Y8FY/QFpm4k1bJNO4AnxES8Pe/Rawt+ivbPstjyQfhkJDZ8UmQUQTQ0wzluKq8VM
S/p57YawCWKPUVvudBgP8+XDX0UKMKmPI3/SBvz3/sAgW04RQJfzPtcWfXLS+lEJ
nxNAoS62gYRbWbikxeBqFCwjR7ir4p23JrHXvNGzwfB4Go/BcGNIsKd8AJmsiSvi
fNecTawymKjVV/pVBhMz6ViuW6Q0DClHicVO/6JsFgXgX1YEyZZh6U97R/tpCC8q
wEf2LqFXTXCWD37eUa9018zwAlg6RNAtqnYfUqHvFStcIT1r2amTDRIpmx99C7Lh
9ip+Ls/civaMxGEvr66O1pVfnAUsRxtQtoCiv7IWiqZ5hOB2DptTI7jOc7wJnfrn
nMCQTZBiGQCW0rFdlcE/pNrNJcX5mdHtjfiNvU/rvSPnEfX8Dt8kcS6Jz9BHjZ74
U3z2wA59tOaFlhc5gsGOAk7lHi32tX3IuPgfyEgs+fSFoa0/hKwgRC62KXHJpl10
6HW82CpOCd0/H9TKPuJB1P2Z3zn9b4uREe8oImD8Hq5dSdT1NFwczGGLPfCaDH1Z
VjgmrvinRj6KkOFalxPEqToU1QmBTEApSXXksanMxPb81bOfpbXw/BNx/gbhfNSW
AAxM9UFK7XSh8w7atCR6YrjSOC8kyx0+gZgmi12fJEmM7KGQ1vXSK4uqCTPBz/uk
DCKQdZW75nbno53O+Odd/dZJOdNNyENRLf1j6tynlVZ/NvG5Bo8ulpDAKtLlhhxS
CTCnzD11bd3Y6CacWYsSm1kUX7flivuaDzUKza//EibGm9GGBxLzh+YB++FGgOaf
B41pUTj0xbQv+Wn6HzaqKDRpqJbok8xHX3BOAiwgobQqZb19n4FAr4viE2JrD0Bd
VJxRxulk8BuZtW85a4kJGvTuq4sMJF/tAowGF/SLIqTsXiiC3mmNTBkGsUQbO5sc
sMxYACwghPZqaT93cKYSe4SoIOrzv5BtTMsFhlVtd0YlRgQgzHtoRmHiZyDkJMrn
u4lGTNq0b98fv7cYeN4J4NPR/ch5dIsDZc0HWz6IgxCpGounWVi7hUqs1wHijr7c
utrTGZd17EbZVyXeyQFQm2YGB9eyY67RlJGR3DVd3jumhiygyvoIKXRuVkGFAseb
1aILIoZEWGSSAY4gKJiHVYZfUwowmMdWluJyOTJTO4Rki51US/4HsfjvEDWId5VP
++kyW4Xs+IMhjq5QD2J4xPtylCxVAJZHgw4rMljHJJJx31m0e9oQYYp1al4CAZaA
dURutXh58sMc8zB7KbIkuzqvd7NMJx/i5oG6wX/Inlh4PEN+4F09AJ7lyt/MkEMy
pL8rZvBrHcuXkA2ZL9kU15xxrRmu5Kl4B/Nl3hXIhusW51Se1T7GeQsFf8SCgevT
swm1HqJgL+0Ory+88kh06T5Pb1pGHJfF3S6P1nUDmboJGAfP7ac2i7PRSewp3hpk
pu3hTZxyPAlYNXDgF4GO0x+RiaYdk8umwbgCVtgT9mYrBeNbgVaSSYAPFZ/K2Odm
s5sTMGY+HtuFrwHpZa2oW7BUwpf57/G6KKCoXXvo2DHwoaL5SbCrsoGlYn9ZxvA1
QfRqDNWpTDb5GOrULF914vQg68cOuTp1qX40Z244BpeAZHiRTqM3o6MPegiraJHS
ZGz5Ed54BAmjwV4yb0YbfhGYruGlxJwa9T4RkEULqYh7LceNWYRGL4xi+lKiUKlr
Nwmb3RRf39LhsUdZ2YHaJgTWhdbFiddL4PBFXSz2WS4R4ji5VWTQyW8YyBhxamiJ
Ii2hriYImSa466J7E/SA3o+1WsdBJHdH760sL1kI2UxlydizW+KY4mkqXFTWlh1N
MIZLlm/QDhDVlShx1X3xQmjkqwt7JqfGLDS5mIJVG2GrVK+aR8PHXr9GEjwfAxDi
JBi6RQOCas0A9c7Y9J4mUDq0rkIfD2c24g2o/yLVfJKj2a9TIdcMD7PNPZjyeCf1
0WZhO6ArxngCH+EqFjTGqFmpfls08VvyNYIQDusPIHEvnzDYkYp1YES083Wx0F7I
uU9dKfpp+YowRi+yC+g0v1WYg3v3TRIvfe5J75LFJ02g8LItF+ps8euxFy3nhKKa
z+wkUohCvMf4IkvvZVNLXaJskucog+ppey0dYoNUBbAmNLED7pxAUwoVvTLaa3Oa
WDm17rNBhLPpuHHDs79yFofOwbCNCSoveYMFJ7qYlQKFM7epYYwENFfQ0qUsawyQ
qnjhHcuOnkQH3p4FGgIqKAiTIyeEu2Tt9DvmpkPdBbM0HF27VyHrrKmrlwoWVTEI
9HzIG161Sp26CEXYpFemBmHsTlRB1kkXx4WGIKE79V4cfMwHmVfVJca0TaJBA6+F
NFarOvLvCKFyJnxTMoDp6skMYwXHHK1xincaeBMSG+ZGCyewYIhAM/5VdWxKG26J
dPia3w+JUJOshl9vDvJLEsDhMAO6VOwIanOugKwBnVaGbrJjaHSLsd/r04WU73a6
UmDebAI7MnzGVPj3E41GgRywRPtBtSCGV32X0xLwD8jcoBMh84l73NRdVUMgOvg/
h4Z854lDhrW1WYK4faaWpqrDrgGqzSQ81rGTQjv3RIkpO2dpJUhyr29PBg5htDu/
SvMp733RQAj0+g9W3yByLTHbISV2n0cXnHtQN+kt5FSpRi93lK5zHmt4z2psgsYj
XhxXRqC0A6hUFVqQkI9RfoAUjhkstMVQ2U+YZOFTUijZsZB5qZ4SPUOjRKqyF7Bs
OfAmkvrNe3iep75Ujne+dNCSqCEF1rM3Z/0VU4b99BUZKmb+SdQ5mPXDQFAOiqH8
BogGaBaNkPzbO2pkU/wZO602HknWC5nhdK4mMgH8UFFqdqSX89Ziam5yCJ0i77Gk
9nKCF+eIN5nNtc0p2U0ncLshfvZ1iD9CJpyfQi+SLEERxIAv9icphlvL1hunKyUN
2MeVsDfIE6BSq0M/nepGsz+mm0wMkOejIFBzc9bao6SUPP2GWuu1k5Qoi2/4GX38
neifXTMnicUQT5dkOA3Pw5jyyYLE6GXQ2BP1JuyxQYcYIssSWU9joBRwb+r4GGRp
NYJns0zH1ocu5zO+zGNOys1ZU13lde3W4f1bEqzBComaQRg9k+fZlnsN5GZ/HoBn
yRSzYe/2+suMI+fBOudON9GDHBFWgTaG59nAoym4UaJ97PFdR7n325ENkA2AHt4V
eL8gFvhtdBeL8Y7wlUu1r8NJo1Z1i+Shi+OJyA9zzCkcPoQt8hc9nuVk70fwn5no
nvKcs5RI9VvI5/Mv1YmulP5B3JsuZWyWbGoZCSQZpIlZyGJ2ZmSlnAjMy9OQS3Ww
g5rGG3/gtCOh/p69GlE1bcJhYXMB277WoL+47gMnHlBfrOVjiH3RSF6kHDoNbAUw
u5p++QY5pj69T6vklHzQEBP1t8JMxijGoeD+I4z19/FN0ksubHIIccFLQgvW/rdp
nqVKIx5fvfboqrRoDVqWniNDERd9Ydd12XyBsX6KGbblYZdxSPW3Jgg7puklqY5M
dFnXIwgJGs7l8r/uhXH697w2c9VTR419YKOvJJnan7duE3w4MgkC54bYOjgxC7EI
DugyWayuAx5LT8b4iCEhPhCkCJDel0QOEIjcH/x1h/Shr8rUtMsGq/dwbBTf8fe/
K18rg+wY6Wfhte5JEeE7VGG0WRf2ndoD8kGThf4Eixd/UD3nrRQ9Ns6LMDi6cSwA
Kn9JTAm0i8Mf3nB0xdHclLP1nQqx2+7UE6iZMgRTsSxyjugmAEbIF0bN75w1yQVD
tCnhfdYqmlkQ9krdgqXyXZhj4anO3IObkztrtOhWOEAUw1oyO4xVjVuxB4gOkeeV
4oNEpt1mGMYktSi820VaIjCwnSwAxj8OXP7Px50o2k3C9yXuDhCxvhPrA22eA0VC
zg6nfubRN4GiMTX+w7dtAIhmBmHa72yi6t/fktQ2L0U0/UMmv00aJexPfCe0Lip4
MMuvlh/WjIeObzur18Lq1olMJwuc7pkV+eL1BD+TcNIIyQacpV5GBXYgSdqOmePw
egPdHmukzqv/KaaOrM4kvabps64vz/vT+HcDTLV8NLUT5dBNBcT/xT2VWEidKUuP
rUxVS7s206VUCCLttWUmWAYehd1opVHccnVp4uysUccQlAQvVylZZck2spcsNQln
I9wbbVqO34C14omc4R6VrculwxP+8dTD2un5ktRJspzDKYxoZYGHixnytzug+WVe
84bHY8zS5MGSFHg+JyLQrHAeI8JZX762a7RGNpgL8fmqf5NJOCS+oJB8IlDWOypk
H1zP4IhP7Jg7RTYyADeirq01fPOUe1v6Weak4Bl8JN6aFHl6jW9NLBuHwXuor6ec
sClUU/W58Bf3uD4mf8BUrmt38nU9BlyxsB7v+sr3OmDzC8h1QGIeP6jvG5OBMGUw
EK3UwFhbn5A4+lHEP51IAamINj+vDXNAgmMNqvyhvzMbHZ/4ybSkJIKV4OH1vte4
205TYSrmE+RMVicF1WmmgywSA8pe8YEMwIDousmUrthKnAtspst3Gp+JQiadfUVq
DjPLYVCz6nWqFVjYu1KZurNc/s1nRTWIds/3pT1qeJ2PijM6fHpFMiz5klekTrAQ
00UBDefl/852oxZclnmLJMY7uuqc15RLXpthaN/ks+Ehv/V+HY8Qx9R5g0ikhNHH
4URCTx6WqRhj0P5pjuOGZghszKOdnytCpP6r0rMTzRt5+LKcjRva/FblGupJQMUc
NMy74Rp9+Sl/yXgEE+asjDI/FafzbM5j6zZsD4KshQI76ZaRvo+in1TniUvQMMAx
rBnFpkNJPhIBGzunYinKqVq3f6/ejGbdWy1vdmQ6Jm5gkTdCs0RPmlGaTjL78+N6
ZN0x2ZmUKt4xEzT3q/JguL46625bwDTkYJq2R5kEVgYfVKhmOVaYQkfCU+Y2oHnf
rgYWpbjrhEViuwywnpscwS4tibn0Q0KIz7o0APRz3Zjou505SZe/OvLoU44N4yzR
bYesBZWZZ44E8J6+yvkKKK9q71CmmMGE3nh9bh8XwDCieiKBjREfHxVnDQgtLceI
bvzQ2TO0nX8QWz5sbg0uU8BASBoa5+qGNNSALslj4stLgrbXnce/hFXaYg7olOdY
6Lxa92WySFpNF7L5pQZIZo16uyXA9y6nJqBGzlorw7OYu21dESk6h7w4YeuUJ8Tc
YTIkTnfit1mahKLnsm2EJySK7B2GTluyttIsQ0WJbZXk0AWqxzhHbFf/KKWOlJeF
cc+WFzWsoPxPFcm3lmn9ltGL19pPAlDFjAy9fobtMpUoPTYpgmbVfC5J8y56HnIr
6MaNw6sPuUPw/DHo6mM4oIhCygtCI/u++Myma66R6jY5hnfU/1YoyF2m+J4l6SW3
2vZP/d3J1Ja116GadxjMbnPLZunCvDSyBWLIPHYt6Uwc7JzV73GBNPbxJCyF7y+E
MsKuilxE8V3PBLn1KoOrGgHEsEm56Yl2ocWHU5vUKKf/Nyhbry+dpT5HrBzrS5Gw
8UKQllHrYtSmJ2H8WAd6BHkbNM9I5tt0SZ7x++MY/AAnLMu5LOJtswir4kgTaLxg
0X6QzgbGQhFuWCVzFcuLSPjmptDmu8LwCjJXwkMV3Lp7gfaqVNjeR+iRCT7lAGgm
WmNOlBR7EQyBHx57aWpUBOm4KdxcHHi1e091nx0dYRzsnp1l34Fq00mVpvVl7zsR
CvBGLlmhz5yApQxsvZkF/Lz/PVYJxD/KenrsuiD4oWqturXOggptN0PJtKfQZ82Y
1VrElK0TN2+Lw1FstsKxAKvgmpAj7qU0SHLTWjOegCTOuUjupQ1wiK19apwdh2FZ
VhAOkQdwSOoMzP1Tyj3ZofArfUOI9E7qBPKbal9lTYXJ/lkGtyTJLy3BWHUsfSe0
Rh5x8HnsT1iR8FzxN0bhab4Nomw+JCRiljxrwQyCW9Xr6KJc50bCwQ/T5a0mQ8th
IL8TZUTUaICYGlpmvnDrhhCuIIp4GypErjiXvnQkNv4IhXXEdTVxGZEVlXEiVgwo
S3xUzLNAl4Y0Ba2nwiGy/ceK8MsF5jCwt5mvhCiyG+F1WydFqjySkiVaKk/vDv6N
OwBiIGLRr90IKW96i5mF5rexofo3UFifQRognN5ACYVBjhRJysWzxVLx2l44SZO8
yKiDg4ZSC6/+y4FeUtfjxG7e4ATY2KwlY/oDWC8ggd+PCQV5VKIaz5O8YcxvbUx4
z5wyOhqlOvn/PZz1juKBkHYIAa5co/MsJamhKCB3g7V8hUIikB4jZaz98ePVpS+1
q/hQjZiz20uZlqugHGSyUpOCAESz/CDLpDpZgEXtyVEqi7KHLr5ye4JXOfvAlCa1
jsPDy4XHksbwsIRmcP80kw/4sHj4C2OCxofEzgk4russQ+FL9Tgp7XXbFuRMT3+x
8zBRmx19kshkrYJfWhR+MrW+EQ+hfXf7adVkpj0SAcvRBVcaDziO15SFT5WWsufn
1Ejf6UG+5rOar5jEqs/rrtlYv8GjKfYJxpRW3m5mvDdxk1gSi8wIdINb6tmkNzSz
stYRCc4QGdub61d/jNuGJ1J3sYPoeg1TrJHmhfeS6qdvLJwzqe+oUlCUmcQGZeRg
6EjlK3arVE1ZiwfBbtbGmp0AXImnEhDk9jezjyrTJ/NPknOEjpGt/3Lk+47RLl2d
FzZCwSPdFt7iDB+7IEucUHRxDSbqgawLPZ3aLi0r7eOaK2FWPb7rVimjr9AgsK0l
10gHyrh8H2rg0hQI4RJpXwyjJD/sGsqCQ0w2z2qRxvydcYLQvHyexWSNhoebEjBn
NkJrG25ie/Djs+F8Fl/Up6CsNhHUGpfgYaveTdCUkJ1MisN/Aaq9mkwxn7wCxzIo
bD+mJxRctDX/OvkxorW0CffW/uhrpPLKsO2GpW8aDo6amugCTY0u8QeGVFIuh+VO
yGtXKXGN4ELMvhhhVxEWw+DtoxoiWUhRYfokErPsrThQQR7doV7I9Y2nkygzCVAP
afucSLoxugU9gCIN3prvVT+lRenmBCVqNc+mUqHUmTwh0vQfgSc0ngpQZe0hl1Gk
TYo918zcNcOrLi9nsAbwYPdBvaMZ+nRKSH+2ZxA48ORh51J1IykD3P9ed8iDtYal
DFKTqZikKODG7JkFrxf1Iwaq6zSLFZjy0I3lVSJ7u0mVtdiiP0k1kQLTnxo3auSU
6ekogE71OXo1ew+5yC8HhV9DU7Cl4Wj1K+U7xZJ8jxRH6XMRirt9mBB763VXTkK3
3EmLlU5QE5CJPz9NR5NdYnEaBm7vMlDfnBCDVT0mssmk0RPSDftFBlQxkwBz0GsR
xznY8dgi5LN0s5vqrDZ/odtafKjz6C22oP2hHdH/dWVL2LaYUIIQ/kRJ1U8roxQA
sSC66v+iWbxsdmZkT54HxFAoUz0Ep1keVQoiF50XWKXNk3qDmiG+Uxxa0Y+gsxh0
Ftkvo8sHxEzVHO/BVbS3e+FyYsByh/V8d3PvOGdsrXBAUa/EEfQO4+mcy7Ez/67o
qFWSX7BEmBCIUSXxZKRd0zl14qo3z7snAZ4YzjVaujod2i6jBLkw71dqBJjgtK12
clGpqKe6Yrza7SNVqXr6DXwmx6NijPBuRFHYre8LkXB/nXrlsix6WEFusOuKcBcZ
LirYfZbtbVrf75j+IiWNbdmkh5zDOBRdpUrxOlWm+YaHlfkOxCLXSRSEpj/yyHwk
T5rMEP79vjbwF/5Ee2QusMBz84teov+NyZcyBQPcei6h16zWrg7a6uPsMc3OeEU6
VlQe/iwUwn9pnm9xT7jWSkRz6cg17bhXKHAQbJIwH9AN5A+a8ACLB4Su0FwK2G7d
s6wBLxuZ6v30f6+TkcVaLgyrgaodGDjeIY1dRg/evqBKgm913b37BDVS/Mi8dZ86
l47nYr1cuutenNroETCNyzP6Hr4h2cmT71PN+fx8NrtUQb+6Oj7ucpc86C2TFPEG
SkOzdN+iaX0VR0S0+rqlPzaUMHIiWT7gxfQyrmSyrZ/vYsFGP7NJr/hK7xreA3IX
KILyWRaoP+aZFnVPvLXclWPR1k2zLuu2MniBDdVaG+sgL2vopvJbOBO5/blFnwVo
SM1/vzgaqsvZVRdMOQhY0GPSftPuHJXhuX8+fzHXAsGNwTLfDz9ToLKmOaZfEBh9
P/zePwNeCcAqu1AvDJgKWFY+tji1EiuOzLdcsmT1mlIPY2YB1vEQYSvW0EzJHCGT
ucYpTESj8Njj0nufzKuz473cX4eaNCu9yocwijQhI64UPSKBhRGt37ZmtMqklS1i
7+xHpP794ofMcrY1X5p4r3digiTb9yRtzkSMBnYyuUcim770z15oljcgmzW6On+Q
7vCeli0AfHwC7eet2aHdB3hPFAb9maMh6jAEBx5njTDO4TdMDYRpZZF+H7ZFK+V/
PYH7KK6Dn0Ig6tsso1pwIaUvVd3lFwI0DnDD0Xu+z1cZEPoZ4cdvrY14j53mhZCg
vLn4UUdRZ2offl6WahHEuhPPv0H94WRXU5EgQYdMYPGPK0rWvv2BGScc5e5TyZ58
I8KQgy+cLdwCyH4yFMLUeyvkSkScVIA/QCnbPyRVRbBlb9K1QNIcn3bC/X55P6sG
8ohmU+B3WlX98kHe7ujqBxtrt3TqFRGOb1VlvdtjjTG4Eh8HYbCE0s93hAEqLHMV
5xHt5QN5OrSJdKeemtKcWWQb1Ym+bZ6hH88/ZkcP/EWot/qvMhr7qf0HqWqOp8to
xJRTWAb/gnU5lb++ZAkflVwkTWaugCRHgLUrqZ0P2b4qyiFwYQ9aw7moAXuMmOuS
LKbokhfMyJrVw/P1EOiUSMfuPQIrpWJPadI37DcYfCnJPXGFXz2nLZx0OlgHkZZw
jNlUdw4ZsrUrEz+7+xmYHqmCK6Fj1RQgsXPwO6V5X2c45VxldWZUEZQ1i5aQTQjb
Cq94ntBYSHGWPZdljUBn2BJB00pTO+akqN3Hf4DAA9/RKqUZYL246yieQYgIhHXN
9ZmdBD+4a6Vm3Dcj7K1o1aR/ftWOjk5jwyy6Un+miXaT8O6mzBTL0x77qQ3Pmv1M
0VZ4VOCxdklArxoelqhJ3W8Pa892hjZrlCVptxNZrNsHgUYDa+o0O5vJkBPVbqfi
7rf5d//U4C6W8VqfJDOUARRWNie9eudjzt7LKMWPVcy33Yp/VCc0guL7Oc592wld
PXRtXZKWtTKiZ87Ac3l3C4NmwYzm5xQquu+iC6bKI4d/ARgxiXjUCIgFlUY0lmaH
cSCTzIQfbMV56BcKx15e+o1JwjSEZusNFDCOTc3PVt7nefyNPxYnnL7OqkB5yNFa
ZOwsM2ahNGI+3kqMo+Q6Fi56/v4w8LoItRlmealxUEJ+MA3RUu3zfgthuYj/8T/1
nrM9fyVok8wqs1lZbBq7jjSg9BEsPH68ASugF3fS5DnxtUCIO+n/IbBaaByVBYdl
/vkIswYtgoIq8QzYyL0r8gsOpMRevqcj/L+UiAXXHuQ9OEraUQCAyGAc5KSjbLCr
nzqLiT9ih7/iIBpGhpbWL1oBirKkWjwZR8X9nUvhr/7QHRwEbZzzaRVERoNueYsn
PFfX/QlVcvuXTqPcHLpCDNacpeGgZ1tzx3Df8+rxXFdUQM5NkRqgxo70bFXWG39O
DJD8TtPgVlczne3ABAg0JivxvTEy5X2GAaCgCMCiWIan2hL1DJ5+8vvVYbVn6pJC
UZwYSkRLyum+XJnFfRxWKQmZ1bF6PE+m1RScOxZFrS1wSYLXteGarBSfwemmJ+C7
rd3NcUubQ74M3Ol2NzfZNfEZE+vU8i8IkPMmVR+SPRp8goInT/x0jSMtbruYr3rT
XuqSV9G89/oSey9IwAk+jymFXnOmhBXO2GoPafFSFUTYB8J6DGv+LLheW2/dPorF
SogIE7FbHyi2YU3RfxdRbqM2Z19z/OF3RaXXycU4enfudGx1GTkUxzMXsjhKjDsS
PNL5/GsJAbr2p+r202yHqtq7/DC6x1Oy/Ykzxe8Kn1ZFydaT3cpYZn6Ct1eikzyl
MYQ4BeG2ab7Za45Nr3f44A517I+F9hcKGE406W6cbGN0UWqp/GkGBsrfjkWluS2O
PIRzdFZd1m0v8GtlEurpohwJqrSnITRgZXhBpkVhlQBvx/vNs4jdzfEVLVPzMCQr
KG5pw9Vr6108kp5eT/Jf64yr8/AyS+epaaV8FbvTJR9EKejGVKFHtUO7WvJEKljY
ZNy4XK0l6gED2rZaI/uL+7z4OlR5wwQTfqjjM1hCMfDxCpKEbYlvTkVX6ktIH0bX
3W00uYYNEVh46yqCObqqNdSGXcnQbcpTyY+YSXUzDcxAkm4nfRSOqCcbKwsk3bf5
KSpAHFw7rA0YnME4GpkeD3JeLswbHHUEECmRB0kEWYsrg9PmyrDGB8/o8NuR494h
EuySlNUvCBUxWUnm5kXKSS5xC8BFdtbuf5REnVgOVyH7v+bqqayd7swd2IOE4KEb
qO3aY1Y+kN5V9Q0kS6t21SQ1AKlVwYKe0MiFzu7ojjf5sacl9EC2kqJJJLWL3hIq
M2H4cgl32nDtqEbzIHSpLAn9f8u2Dbi+iqEeZtXB1vn6ObH30nuARuHZLDNihyML
X45RrRgnZ9qRG3XbyTM3B6kavQZOqNrBVmsZpw67vPjz6T1E/paPMe6bmdEdyu8A
1QntMNbIil4MNF0upRW+J/wzyt3/cvzJIntUhMgspAl4k7hlbIC664MGXFt6ClHb
GZvcxdb9TEDWT0D7uipHTffnNkAsQJ9gCbH+66vhrt00DBg6QEp9RXaeDfQ62CJe
DzaZc8vYjchfOoYiarwH4uFVYiotVwzyXHbRrN3tR3K8fN8kajjLqArfMKNX5S+e
QsLSIeIiVeRcePunt6sN7SEI9AM0sjN4K9zNvg9Arfk8KpnyefiKD9dIScVJWZkz
cScfwXL/H0lkyvYRPbCqwGWGcn6OnMB7hOWJiYJlno+K0IXOVOdEmYnnERtLwRlA
YtxhFzMXIUCNMQXK9ZbClU7mvMuKN0szBIHYElhSP1FEzHeO8Ej6AzYqjy3L2nSP
T5Sx24vktrQyKQpER7XhvzHvjgLeRGGod161v3A8QljKAifeazpsTgTP5yS1srjn
bzFJofnBMD0EUtsz+T8a8bgWekfzPNeIFVImEdlZYhOIWs2BQCzcyVZjwbrxGMqi
F3i1Z4Dcv1hnmbU/mnCSUfHUhx0rRQIjHGyy71OvkO5sagaMF4LX0+7KLKZHU+qV
f1Efldv1LFV8lbrJ6rWoWTXYPaHDEIuj0dqiYxMErzTkKYgoUjzWywe23flXpDs2
Wk8Qm53M5w11TjswGpo8RsyQyOhGEUeNyA86nRcdKJaMG5HiOqzU6p4eTs+4Mt9g
YGH766NKT1xFlNNMlhnKeYhqOpl9uQ56m7vp5UQNqyeGznKX0C8s1D0e65Rcgm/g
NgETIaaLU8d5jYnDIsdz7meIjJruJyIvHWYpZK//ylJpNxh0ruoztiXGkQ/MLqXY
44gG721V+mMAHzyc60tBIWveDj7YQwI1G8aylcuSmAsLGEuJGyK1nIwb5iYcEDSD
1T4vLf/epor7J+ScRHuIgFKRYwEzgCHd3wNSv2BqH+p44dVPwVJP3X4jA7dYk+pD
Aq5zOl8KxQw+ot6BUNlcOcjn4dezlDf/OFO91FCN87INOfrDoy7m+SqoTV/66e56
Qr4oK5YP6lL2PNI77hi/FZ+nPcFxN4gpyGqMG99/G4Xy7d3r/FAQ42RJte8HDuLr

`pragma protect end_protected
