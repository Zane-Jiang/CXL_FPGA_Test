// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
qzXc0WmJB6OjAj3rw9I8dgd/ur+EwaKyniSOtsrRM9AC7o/lipSPVFVuYramaNvX
lJ/B7LGQSIdYX8TCplMMfHW1ROpjWk6b9hqAZAH4WfsRziUBTtyWIDID7A6CyvZ6
GdFmo3l41U6GLwpspJ5HFdRoRtuYsZPzmdK5SPTpdqA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 67280 )
`pragma protect data_block
Lp+Hup0cpGFXpT7l6JL7apPGFI8MmPtU3jEvZA1wquxGJuQcff8GJHgWBLkKsQIS
C7aGL7EGvbbLeTQf9kLW4j1lun2qmr0DYxJR+h/etiSE/0tY3VWsLIxFhW49osim
4ij/cb/qjrah99m2YL3GZBjMAV54zvyHxUhd7Z0R5bsx0qC3bEu2XN+AuCBOFttZ
Dya9qUgSghXchq5PNhNwROwQYHHBJ8U16l1nr4wSjfNmXvn8Tzp+0nSTTd/g9rig
hnBhdBrlbMAWK/Ieoq72rqWUiwOZZpZx8G8GCrzxxxoQ2tgAUqzhBeX5o2Y+BUuU
oD0W9ILdDLpS1YcdX81g6EvPwgL655JdsGVKw6b393WslzHmvtnIyQ8sTO9I+0Kd
lngJxd9McmnaYEOq3HjkKu4JZSqtqHQGC79FI1eEjydpqpRkT+YZTJ0W+26WfZcJ
m+c2ofIQcLktbEMKbb/pNJMbVxhnjrGuIj9m36GW7MfAjPdV0fpkOYQtraJZ6skY
ss8IX/RlbLA7OdePDaWsFfumFAKZRXp1/vstyAfVh05EZnnHwLUcqzhnzqPe2Ymv
Te0p9+IvFHK+eONa2c4O6nvc4p5Fp+lvNdA3bPoo6o2sF2rhIrw/XxHhIW3E7tUP
6YuqBGUZptrtf1ZDUfE5reczpvUQ/vDiiFm2z3wQl+PWnQYvzhKjl9dCdC55B5bn
0vfJ63WCZy3LrSlzUP+a0FqNQd+AAXVXUqdRTv7ScFj62j+GMPaVnX4r09aFELmL
URDbcILqAu9rrcsCiqLg1Gk7D6x0yBKR9z+Od44rBgtaHANwZYfvVVRHfbBavH1W
GmA4qImOH+72I9DsFqG+rHY236NPL/yvuNQH9OrXJ4PSbdghGbraSmqzJjG5ejQl
g+QuM7UM3tqGDdUkHp5AOWhBJdNl3EfKIRvEoQZQjE083EB+x+vdnGMCqRb7V1Lr
7XWeoF7E+xq7TD3V31ys9axvhoRzrB1dLr9SFcixgrBgabGk1XfY2tsqcL5TxPsR
vvNWcb/9nkczzTlC6DoLl6oArMsD+kawxXQKgjsM0cr/cMyc3ZyGwlPosQzCExha
8LjU34vXYBGfnSoX9+6PKPFby6Y/P+KG3j1bpPIQo9c3YAI9DGOOYUnzu864cTRI
SN9rsOeL2cemsSuVeWJrx2yF242xll6oTMSyR57N7F5fCHVofpKTabHyMT7NBXf2
ana8Oe/QzCy7+AHoVdtJ6SzPBGsGhBR9yZ2ThBhSLHKKPYPSP1SNyskti+kg11Jt
dxF/8f8dJmsfJa0zT99ar7QNJ9JFP5QBTHJ9sCb3+5EwaCsV9AGs7E8VE2i4akcq
Qnn5hffz4CoZMMfFXpj0Q/tH3Y0nRNMRkl9ZeLnw++8VqLpPhDEPwuxCJa7VSVyL
33xg9ZGvaNET9qnDIOEPKmtuLrHCUu0FRnPlB6dXgv21JulPSaZtFzmYx9mpmRjT
y8hWEcbYmkulLY/Vd6JRqYbsQcRJW5Lht2LamNgyHnk+j0VBOTmIDK+9zNBgHkab
P6pnpwG/Om2CF2DMUZnXoktxcVtPyO2h92T2WVve6hIWVw6aXwNHEdrZGa4pkPr6
CZbty8vqdCaTkF2WdZox/wai4v5vENBgcfdtjw8+Hrs0JkP6ZE2vpKRwV1fpBLog
UwyVBipqnXa853ZSY8uQXA9Y39snhYEqYnFxHn8KZKCpN0zh+riozH5x3rv+z+WR
5SolJwVAQr241RqU8eOwzJNvpNSONF5Lrz8uUoWV8lFoqLhTEA3GalGCwWTDWfx9
3IF9M8/+SpmVn72fy6P316VID540n0aho3MyjyPaUMid28gimMwyjxNIyMZ4SE37
tBvVXYLvdJrfJb5ZxDArybxqE0w+iGyn3SNoABOGIsMwP2d07Au4PJZn8+jx6kLW
WTnsWDP6sovUfMVOcRtuzAlqiFh10I6mxQ+/TPbRCgS2aLJk+X6q7dnUT/s7yJp4
Z7zGoYBUk5euQAjPtCqqL2/4wPnjSVMNypZ1PfWydr8hJZlTD/E46H0EMH5kyEKG
CSWrmvloMt+dYNZKyzxlZ3pdvmlYHrP45RicxBlBHBbQLu3SH875ITHX16KrR5gJ
RJJwTF2tF36rGpMyImft7A8COfuQxbSWQgf+O46iW5gQqVAqJ/AX2N1GOjczh8It
/OkDLDj3peBXBQTi97yMJIJdS/FKb92+OstwK4VVBfnuE1dy7LrUJwc52CbSRwPX
nwakLcMkrvz7kSsMhC0J9/lC+9ldpBnNDm59NUcjlJBetm9mPP0urNS07Fk47WF6
4Fh+yjPmtGqzZ8UeMyljOuqo/WEBwYpCHNEtFP9H41wqx44LFc9cVb7CDjDDplpQ
J0/YijGc/Kcnf0GVgwLvcGdmWL4ZV1aYxicAlHGFumhpSR49h5nb9g+XUgM9srOX
UsMEGWj2MZgjy6dvxhl9zHhRtXROUPJ+L76rugnnWFgBB1k3oVA6mxB89Zs45SlZ
fImz/K9gMHhY+69T1dWOyCxULZccWat4vtvFYIP6D4ShBa3X30aLfrk1qCRW3PYj
0wl/XuQoMqtU92FTFAmQ6ghM6rOIAg36u9ABsORP/qVDupOha/Xs74Qwne+r2XLA
+Cb42F7S3GPGbQvwt+f7I9sv8F6hbSsMPMPKJRcUZsvU5FqmJ6lkPzauCqk9QZvt
HfLXh4bGONh9Yr+F3Dgq1KLmssDMXgVUzJjOU24fqIUajtsz1rI5PPRrzrFb7PPO
fUdM/IMcfdQ7RbF9/EWA47yLC/NljK2yNukYpvAjlRZ9Y3IfUzJl4pGujuUXDz4H
7AGixaEOtXNrrvvA/bzYAlEuPrUwUzuSk7exlaAChqDX+GbgahYYDLjb30vGVQ0N
UxeGmThpHZf0i+Cp+yi3jlBSDjlHHEg1B+LGV6rpdPini4T0lGGKkKzRhKkggA4z
QynCeX8MrrxvMvfnTDPagZ/ElK3Eo2ij4roFQCGZxTMCvjk8FA3xxecz2UDCKQ1i
YlD6Rf9AwX0m2t20PwxYf2iaoRpLNSw/7IOvuf86KI2eXWJsoeeZFUkbS2zqGRxu
omgklY0ex+0eBIIqXiwOrr3KDoBhryCmGWfDdDWUZsAws6XUHx0zcT3dhvw9RSUh
yK2WFXq1fgFEjTa6fuetCbgRn3IjOaSiiuZwruApE8okBBM4u7sm8RS/D+UDcA7a
hlaHb/DcghBb2UAsE8rjN9YvTF+hYzg070lhcinFheopzjN3RKZEtcMXlPcuQtzO
OvdqNbF44tkFLvZlx2gLLxyb0J0BZjkgyJB1O4hb2QUNv0wsNd6RWJZpK1Apqky5
8wG9hdHAArnebsIAw/z07Stbl4lXFxMnDAYYgg0lGLccgB42c/FfQCPj5UX7AqXv
va5sbw8wgnBUWEd9KR0PP0sBu2OIcYOwkMo235ldfKWdRRV2wPzoiuLwyjbUH0OO
VF3p43bGas/F1tVliW1FIj1N+y94juZ5lBYwnRNgMd+LRgxtb1PyJWyjy2tOK+mW
nDfbFx2OQEcPnOfIJks+fxVebDGVbz7RGss3FliVPoWM66kWjKnPHEBNvj+/3BiO
niR21HdXocjPY9zPd4az5LgWvKvGW6vJPexJbQm+BlAnwSWL+IOXZeY/6SV+TWdn
eMxAG4AbmvavXC1XKp84dQeVy7tDy/dfoMm7k2D/8zWCAgOeyWaxqnuOuPKkKQaZ
k1raavpk+lctAL209bS8tOxgwY6A7jq6d+NMj5YnvfEXuyd4LooQhBzz7thWR7dw
idE+b3jyJgSbxfphPwA/p2cflNmYV03IpKhRjBxWPNKSHunPESzChd+0o/O/1RGt
tpDWjuAQ/sf8RJCNfa+3ruYy300hHrqxwcVkvnJT4pzHh3XR92Rproqd/SOVM9ol
DdPCFmI091/teyqev0gVfE1w8tkJWgnyzU7hyJ1tjMmU6D8Q+aF9ZrT1+TsW9UuG
I14IMYoAFg+zhfLnGDBM/GXofZy0YwkNdptfwZwXCiNlZM8yD154G1ODXqBXWAd3
vMaVQTzooP2Pb86skuCmCuKN2Dx/s74wJTveSDBFcopIWTXtzdKJBf5/Sx+7GdF2
CYyaFqzj8ooRPTP2LftghN3AMuQCjTFgJuVd5aq9mNRuSFcWDbwE3sEhln9OlLSx
ktqCj1NhZozyEFgQT0PG7jYp80Q/dljYGXprqlGJqivgxy0ETNm93dBfmkNpnrEB
NanuTfwgaagEngRfwDsSlIttCJEpxB/c8tUh45RlWNN0yS1VGou6FVyaer9oHhQJ
o/yjszYgwdaGxr6y5iHXqwnE52J0GCfTFB3JWYOaSna4TjqIYSvAnZ3c9jCoZfeG
vh9exOT1hjYkKlH56Mr9QYL9Nb9zuifeDmc1lBNbxVLOUdekDTwFPy3GQWK8INiZ
DdM9LU5PfS6eRFpDFjDVEp1GozCo1JnpHpzC6O+R9oG6TidVoTYIg/MWah5T8SII
Bs14nSA25oboYBh45mrZwz+F7jLnUT2hoxZ2ggFqmKeCngGyauatZC6dGjnAqbER
tpWO4Ddbw/s6fq6PSuaQJ+PKObxTA5ddi2OvquLXMgTxzqKr09AVWiflaTLgg5X+
XgaC8d9UVTC8a99hn6iF+/qJkI7HdSe3WGvFYa90CKDlsxBzBFyQdCcaDHNOX8Sk
N1bNiILDzMGfTRAFjQZ3GF54E8/Y3EVo7RtDOEBiRUFom8nHOyvL9tX96yfVJLZ+
5QwbRM+zjTokLel2UEiT4dd58oo3klN9kf4AkQRq8YnPtD1Sc5CDYtAm7Hhkt8TR
tDypHSqbwK9QcQYvvDYBpi+9F+lQ1OiygYLlg9yTH+qKH/635i8GS6XOtLqcFT8L
BDbgG31r6xJWXGJL+8J+V9imeSgfJY/9RUOSpFWZ9JMDAdFKB7fLiQprOQR5FEc1
vDzYBvxHMgt6lMEwNIgu/KM97LpY+xZOKPSUW7zS4rmvxzWyXlAbhYRgan5LBs8Y
DOVj5szjRQ92yQ5OgkflddrBCJA9JKbpWGiNa70e4Ww5QXDSvpqdIZM1cuRi/0os
kCyMpnktSXvVseEoCKrZBVKncHtCqNU7uVdoLpmjxFqFROVqurdwQP/aZ5PAIoqs
D0V6HupTshdU65bUgY0Mv1d2WZIAm8nR5e698K+NFJsgXPMdKibFQseoCywnST22
KzNbEDIIV+zj/JKYxOuKvejD85/8T3aDgo2XVp0MgpXuozWehPk+TsqD7e47xrUe
d9G1wPsM30Y6Gm4N5AXkdXMDorvRxNVzTBx9VrMJ58MjEDz4XEa8GpRmyJZTsALU
g8YnmLzynzw/YncT/hO9QlgWmxtI76Zf99FElCia2a/SEJLXXJplN0cKIweZYcIt
Ux4gtN4MZZRXRE6OwSjcikrQaGoDuS2qHR/jJmVYj8/ZlR7ijIllk40C08JEiNEQ
GQvxcsQJG16jdwzG9kmHIfccbfZETRG1idIVhz2FdgZUQcF+QyfUBSqu7UEIKAN8
Ug6N1G9pv8PyaUAvzvCmZnvf4dUodeE9FXAGhWQnRGSc0ipdgaBujKHKYRQ3hvA1
J9gvHf5/wto/OJmDEr9wrjbtrrCjtQnc05Tag6J26r79vzp93jk4paIC2HXcSbXm
hqamE2+miXENI4R4NpCyitFYCzuGEKrLZel0GB7P0pRntxOofT4Cwn753Gk8QNnm
3YsxqCdzzUXJc1XJSvWbNCTS8iHF35EnVNbCOq0y8uStJgqIRsnZkF+TEz+Q++Q6
e4HDjc+OXBTtvUwCEr/jXD5f5yyv9mfOmwjCjhui3VsKJ9kExHRmOBAcPmMTNyfG
7yj7uQ8xFrM6eLan3igtEZRL9leuvge2azjPp7fyu29JelwlvhukjPkkk9yZWCp1
ipddeWTRO2YgrqIc6YH+T7ZinYbMDzLYf9R8FfY0+jsqv3kVg9LYT6+VYxA97y21
JG25f0kFTm2PSAf4G4qmE9f5wFVDVYDt/iMqdKCfWESaUGApdqC89YYLwmU3bex3
KKkxSC2zEoattZbrhRFt9ssi0ym4CmwGnA8sgpEQJJBTkK67XMtDh0SMSWbYbtnL
jO4zIzHtyUUXyk0cDadbErKtx4teLVQhwwxMpnrbG5hmvveqvtM0fuX+Tph5uZhx
JfETqZjZiji04C3FE3ggqtB0VtYBsIju42XAFWrbCK3lboGN2Zi5dBsE57neMs5L
sh2tJ88+dqiLiG3rr2udlV+jaMFLWkqUDv/aLDUbEUC/vriOqAd+9hOTXNvfT6E2
LrRwSJez9DS5wLDtUZWdvUjHbwK2wMnXbjgAFL0JmmnZM8gjKSGgx9WWruPZVdlY
w315cZV4Fkg2nhomQ4PPA9VPiSTHfu/g2jZ3qEoTtgYgH1mm9Vs8+miCn897bDHT
2ZoJwPm/MaDUJLTUew6pzpV0njoZub9xv2wM42atLZVQ0KqASSbywaIiDu6+TtRy
GIcoRXObxJ5GWlaN7xfkNVRu3ZEH93jmPgJG3DKzQjH//HMiFxCJwrX+xeuvM+Uf
xpFphjPMMIohHqk+ILhTF7b4KW8zknELQ8gTjtEvSLuGKgPVsYE4gYjf4T0eTheP
Q1NqWFORl1AZt02+Dc+0hnEgbKt2052V59JKOHL0NVLQLfMVQxkAlvGV4I2GhwdC
hqYg9d9qaLDJ+2WLnpQOddyuVcCKvkPr8wpPpugRACshpi4YNQu9tpuq8HhxEi7c
Ugc+26dafOTSqjYBZkKZ8y60X93mEIeNzsdlJIFsJtiLyqZWADzSkkNEale94p2K
U8LT6zYTTc4U1jsflwi2vJX/plcK7Rq1Zv8pFdgavZzzmR00D+EZl0+ybCgpJmAc
0/qADUJDMUhM7I745TUX5PGToZDjAvl+KH0yIpDqQlwyOm05OEImNXAWbkvbhNJ+
p3qvHh2ibPzo25S3D++Ys29EeIwIxISiZFnDGGB4o13AHG1eVYPoyk1OhEQn3tfU
YxLek0ERmKY7NtfD55yIUZhuXQJYFlq5ko4fJuChsldBUf/A9kLDEx3JZcUfNEGI
KQc5rAKaFmXP5KGg+zuciQFf9+8V+TknVaowjqExoqt8pmknAnuMu0zdIYeG2ORR
GiBUOuTR889eAyAyyr4kgQKSEKeGY7qx6Mayx3yBmV2MlyTtAwGdv8QSPb6UM792
JLzusIP2hlK5N1yDp5wMdTrmis+B1+K8xMBSOVW15GHftSB5rXDPl6AzkVoMVJn3
i5TzbGxIl3dVMib0FcUCJMNPcj13eoLgl3JhYP2oGyZIjvw35EluzcSn32+2Oxbs
qdXFpmGBpHVKeKA7tbUWAN0rnhyAXQrW/zPEjj8RzdvLcsA9pypu15fOGhi8SIzs
tQy0aMw+ot35gc8Ll/O+xkDLpYzc1T4U1T4CcjxQKeziNNdtZLP6KlUjKdXcUQLE
gajH4v5SicGF/tLT5zVLuAPo5PPhdsZQv52G9CV8Qrgcq1Y+CZ9iPoJtIVgY8iGy
Jg4NLasZkgb0AIs3gk+8Clo9l7ZZY4dsaXoXOgyxEkE1tPdF3VexM4i5jOX2+Rdc
IBZWQZSZT1FscOyWv9sD1CRPxWCAUz7tq00uZXJ/XrblkMa4MyO0p/Gp0Aoguq1Q
30rkObOAyKa5t5auSujnK4wxXrsoDyNAVLtz4zqxF01KT+fv+inbz0Rzls0+BBrL
l+LJhuH3WQukVM7pRTBm7nGMx46NM6iMmB5tuPb40JZHrvxTLJbabT2h16BvyMF+
pKWfas7whbmLJwmEKblkrU8NqBp/c/kkUJRRXU0zQyWQ45veRyJHFwVk4dUyry2W
5+H+qP1RUBeJzEI3NVCWLOGJFsvR8dwk0MkBk1mEiVMsX18SiJedtbshBlT/2QdY
1YPCLCamXSVnmE6xYSru7bCGCpJpttitB0sVPrKMC2EefMI1wvRhy3VO+YYCpsXv
gUed5CYaGJke2iJZ13p2iis+dYnVyE/w+BoA0UecYKSCWdVtLWkn1jT2p2TDOcZx
HGo9xzJVAIifC9NkXShumas+7cxaKX+BjP3RqZB0T4OympYBgIZ1E7xdPb3qoDrb
2F1htO+cNQ1/Ltm7Rv2IyGjxGyjGtjt2t13bRQiyttntOfNOxI02q7YGthmy3SEX
bZI0wcXq5Xi3WNpCygJRQ084DY2LL7Qnv+g1j8b2CUkQPxWrJ0KbsfxP88GtfFnH
Ocqd9l9xa5OXitcjkkXCDpjo2ZtL6RFEwuu5F7wbXdG3g41C5FkRUSsRK63tfq05
vmiqcMlfjDwzBZ9HtjEk1poVCdKbcCLWDWoNaCe5GNK5JBzIcf95E16FL4C+fJzs
mJBAHc0WD//pCoZmWMzrBwZ07KeS4M81ZiZmKBmTqt8M0y/1uR/CbNamjEl76m1X
WKJILGU/XMIVe/Z9mWD23yia9alGtyBK0NmBn/eAJ9SWKAbifyrYz5C8A+Hg6xVd
ptalS+bMAQfl4xggHUGV4lHIiGLmBlz4e3I+SuJ6Ao6Zd73q+1fMQBL+qyke3QKY
gjDlau9/mNQy2wWdLECnwcpXRgDugZ3FNjmkWIrzKz6Amf1fCa526Zn6JICB/zyv
KOYDK3zd/pnAMoHQH6R6gCxLSGMOv6LQYJGKCV99ZvURxq/9uFx2slbNuY95n67f
bnjvhbQCW0LALTZGYFw+mp8jkGyK0S/2U5z7N7UN1GYT8z9K2B5Um3F7pvJdFq3u
PdiUdJNSxyPkcYdi0LqyV6r1QmXYX7xezUNJmC5koCgf4pH2VngRNzgbEKnicRmK
h4A2Svsf6bocyQvN2nU6fpXIOUjBLiLqsav4zprDMrkYIQB0iERsqrSgP74vRrWH
DYPUeYY6dEVnYZ2SROBCdxWH64aKAGcy6Wjy8ZypJTMp+/EY/EpSe7n/xm+f4USQ
/zZP6k/5+qpk3TPk1imUjI/JJ+dt1c9BzRTMu2r3SE7Ef0sp0Y7N4IWdE2xJ0kv5
sOsx3n2awLePUbv9Rrrdi0nZk7kshX0+FN4TOlR+QOGIf9LBrVnL6tot8QL3qPsw
W91xy+DPVL8IJAeZ+1N+hRlLNRvWrRHsT1vtv4q8BtV+7GMXdjykQKKQzg7tVcQj
V6x5VdWsu6rHXzRrrIOyb1OUKmuLb1LecXfjwMIfyzVR3hYlfqoGutUYVSHOoWcI
RurK8ReZgghsSUBpTdWAn6bad8lG5U0gZ3spLy3ld36Uq2QNFuwF68gPVFrYPfqE
Rgkd1gL/Llt+HVb249Q3uKMP0CbR4NZVbQx0l+/0CbUZvOhRfeOAEKIPvBoWkclq
D32ndTwOEaXKR/JZ5M3YMqKVp0c4nqY6DIfeI3tNTIUfi+172BX0Yprg5yAAG0n+
GJS4Pebm+RXC5DHuZPC0MHS0dUjIkqzSkTTTqvg3zqPjFtYnvx1tDgaLNDV7mzDr
wovvZJec0APtTFnOr+2z3DS0NBqFmcTuJrEbws6jKIwgiramaKymTv0Ds4MXYkPd
fBbL6uZbRIX+fdqxDem7swdXxdynyq/PfRRebkUu4TgNeQOzuNidjrs6ovGE26rz
UmG/FrVrFrV+G0+yBQQ4dkYmrcVneFONXBk8PMGfXptGW2R8+uNAod3VNYUBD3Tv
wcB4QyOiogGQ1sHz1VCGEBCUbZujjW3SX3jfswiFPMtmE0lTF3S009W+vrkAAsJ9
vsggNd/HDjtz4f3sNs0zj/qfqvj/cyXJo0tH17mZ52PW9/nrz1ZARIDAGlhFVxwg
wpgQHJ9s07TGqOBQNYtn5mn9/6UuGiY6l5z0Hnuxt9WzlWsjHpDSpUjmddwXXmzc
/GI87B8CMiTkUASXVZOqqhv1s1sWBxOGwGLH7mOV5zqJrW1TT7vk59N+X2ffTmj/
FTzmpvok0Ya96y/r2djZ6bNKQ8BA73ut8K/5jM6cmGALxHvXyVi9HA9ssKPY5CA3
djPt+Cn7Pfg94H34Jqflhy/Ne81n+3wiWPMK40NxwWlgO7ML768nCyYZr0jQANXR
6vc8CEhHoo3LXXNlIeurvsVFGMjlaMOKFo47TV2MWD/Vrf9N6/69XCPvVPebwbhH
WTa+Yfe3C7bhpb1ayYFL7oDjDSi3o/uKFLhE/gmXFjPSHGuwrIrl+nMqPdvHtj4u
1ERlIm7KO/t+k3oGISkNisQyU3zVOcTEPgctrkORE6jJCr5RatQCuc0/hYJAKOqm
zKJNOcIL9Z8lJPFKkA1XswvpOfaX+WSMchADGufi2NfSNnkxrj+1tQazW+vm7Q2I
7GJQnFmlohb/RDcTanP0+Ze/Hs9bPQxXmEB76Dbc97kKrBueFFl+Js8npq3wBjJP
r9hjBNNsRW0nNbzJObZNzuD16ihDd3JkHx1vSGRsewxOobyVX1AXrm/4K02KxORN
3yZkou8H8oGJhc0Y0HuO/OBvqXCd82fKFnAfOm0gPlzjRtSFWPM+ZVIBZyFB/D/c
5Af19QTpAwOEPD37dG20buvF0VCclZOEonlEq2MIZ/OyLYzMzYP9OXNJW+kRpe8D
74Cp4trHPCQby9ac0gZ3i+aS/5uNkBER5W50LKeuNssV9/mK5s3bmvu9uGXEw6EM
dBdgzYQK4MWcX4nxvOecSZ59LJ6zyLiSa2GdPT6x7hh6GFW/+fNtGJyLJ1Xs5dux
By2liLVJXre8dOIe4Yz/RKieB/o5QT0wuoeLwliRmkOqSHv1VRlJb5wUWcQ02+EW
DvDzDFIaEat0H/jCypEkGtkK+ZQT7xErk96UHTHWqUuYqlO+73bANnRGnGp8fQ5o
8V4yiskHnxh7CcSBIdILT2nLWhv/4xgUO4sq3/XvOu3y3gRP8/4n6KDsaBu/bXO7
TwvPImngJJ3HFyVxiUQCwqVeeSXsUPUd1yUDTk4zKKuXjiEIaovi2vWoWe5xZA4H
UTKbUh2yIebPvej0LsroEmjb7S6B+MTbLyNTNfBzdvGS2h4xkufb0FUvxI6miU7s
fq5yNZBSYqF7QAsU1lBjPIZLMcDjnYuLRcenH3zPFoqwVlhaeuWKs5/D5OmhfEBO
gyrX8UW9NFvdCkspvOdeRdn5eT3bPfneZKCaQGnNh+oSMDuFGd/bCaCNCkOLEe5F
M0LVEDpLfp7EFqVc/b5xsXHcDJwUOEgDFok3m5zYjM0552c1Uomc5x1vzQ/sp71U
wU8tadck1v30kpOF0T2JH4Y9AYrJC1zTc434AxUHjUEPDzY7jOPQCBqyN7OmpXkn
tUPAhwHeKtNQNfmBHnzFodbKofYcHTqrf5N7LZoyJORzzVrcbIsyNMy/EgjTZBbe
M0HkS0mPq36BtoP+VocjKukQBrfbIFkWSslt7Od4rvRxz9RcOJupnt58Sx4I1/n0
5IzK6uJ+pc/etVCCtbJ8C5f+C9KjdiMVjrY+xzAzbfpeRGjjMTlJ8CTHsQSYFp6F
ifjwAT+GrSn05kSmiiRk8Hktipbob7Bjd6ZgaHwkk1wcIgwc7iAFzUVt5kOxa4sg
CdsRwdqmOkgJdPil+3AwXzIHTo7QFFlH/uwf0Ap+Ibnje9XfPyXj/r6TjgXhA9s7
FMy/gG/QCazof8i6NTT3xVoMt/awnfPsO0MT7ENrPiaygUgtJy2O9+vOs4hpr45+
ZpgG098E2nwOi665Xsq16gjG9y/JKJ3MMb4vYppOUq4UerbAbwJZgyUMImNwq1ai
LgGsTPxU+cpCx4j0IAhPwx9hHqM0F1t4iS79vU1hzFeCQ/MSoRfVlN2l1Vuj8WYY
uPO2/VUFQrd22yY2WdOcUGpCcr+S+PfF+uiR5IGiQwhYIZlS7mzEsJc1ITIR5dnF
JEr/BEIu3j7Xw1As2q7vq3UIwR/FL3Jntfr/rbIXPRWdDbXPtSCX3+IrzlBiMCPC
t2Pt8XS/AMtW0e97scQ5VhRuADpvCM7lff7C/LY0Nc206FqTnbtrd4ClK3GJHKTC
9lmt2LipYO289YHCWGpadcQE/0DxEtlB0KA1YrRS+kWPNoJHhCNGzUTUotSIcvHD
+QrEtva1MPEkz3zfH26MS9otV1TfZBo6ncE5D8az/RMPmkQMsmUvRuFze5KJdpAL
0LLfEkdTWBuEiObplCBkUqinSAAEC0enadLnQ16jZ4/1PFteOjK5fXtNTlhkbTGP
SXu/7SQ69QyPiHjpqiSvAYyE3CxPgCnNmDJc4S2zOmWeXufnUur0/x7Ebc8tOk7W
ZHmuPITMP9mgoFC0PK9W7NhKcptp5NumXKHZyJQdsHnDfu/jqXOcWhQ3ZrH6G2LS
Lifztzze3ra32O+avK+ObNHiLfYuGQ6fuW7fhETevBeLMmTwA2TUQ+XRckN8cmU+
Vbcufkqi3ipreBQ6Ff27o9tVgEJuKi+83FVX1SXlxyFiwZyb85ePQXyH7TlcGa1v
2oIIF9mDm+fWZtqnaB0YQHn7OvWFAFOddbV2RkluFWMFyyC9TWeCMSUntcheOvo2
nR1y1V5DL8Xwwe227r6ZfoD2E9NaKYlDbrQaMGDInw8zvSg1u2JDrAhCg26++ScV
+nFs3oW9e3QA9YCx5CiCiqNzpGBj5Rf70lZcKKjDD+X+2DZBl7fomSycAxYMTZ3z
y+LNEZ4mGcrN4CfEaEnIPtoqBomPkCVJ3fhsg2GPr8rRzjSerjkdeuCUkAcqzkRV
sJLpDrgxMBqTkQcvlVMoE5d8C36IKUZRZWuEKzw9U87SN0h3za+ENm3xLRPjIrfE
8JaA1Ej762FcYbYbDfHTkYwaUXBj6g0VKsCWnPtYNVQaoLEA4DrTrRCSS4V0nn0+
tvxrsuTwGV05prNIIqFLeBmJoNWCsi6tamwbfRf44v05PaTjxEMuq5fKHalP+Xxh
h2iimAXPIOM+ZmnadhPJVvgM+jIdmbnK8rUoEsPq//tfM+rgnaxOVnDp9Sj4S2EJ
imAFfB3VcIRvDMXlaEywIMSLL6OQobFqkEWq/3+MP4N8jInEAvdH8oPd+jY/qppc
F12MiICguAW9CNEYz0D4VleBMS/zWatjlUp7m4YJxmdXeYB1gohHgYqaWgYKdd8K
JD8UXdABknHIubdUw/ARVrFlxilJdGV/9C3fcsaAIemLZtTWdni0Do5HBxdO9caf
j33zt4LNwrMdF9SNXwlYiP60dW1pRApCKuOceHCgizHji/t1QwjAIt38t9TvzTWm
iNQ+6Lv6vvWHBngHztfsiUO7sBONCRoiJus3VVn70Z/fCDgi1fjLmKV1othODDY7
78jP6EnFG6ADGBHHaHkChVqUQoZcdSUxNXs32DJH7OA0v9k1UOVs4JVPxWXI79aX
PvVrrkxMDdxiyIHl3nb3/sEoa0hf3LN3DIKgst6S9kLOjud13EPOmFgaARE8we38
IVp7BfcmM+OIn/aiALLGXFWh3w17MW/5S1uVrEfqxViUB+M+P00DpkAfL06SG8oH
fONiOe3m9vrOxSnJCwfeZyQ00QAir6/njuSWNZjgyeimLg3YTCkpnhhZX3e4LCGw
8eIXpDVle+eDeC+OXdSD1SMN5TWfZI7/mlAI+/pO7EzGevRkho/BjJHNFmJPCj97
ZPwe/dBlBw2z4thzKlexrln25Eh7fPeJRd4qOZwXfGjgTrhtMJWDxDqeaigmwT5i
DsT8RIE6BReSHa+u8JfLj89IqwfY7abWr98/9Jvn0tzZ+YssONu3CylhIyGketzH
3Dykz0iihvnOB4Hfgi8XMYxbAoKry9YxTZVsSFPGb4L8oJZ5EixZkby1aYvp7cIT
QLOLei9s1U4ZNyJBxCo8CcY+zXQhTN2vB370p5cQyhJpvAlR3S9joy9Z9qTzVAC7
OkcVzUua9kifaiXD59+fiGFg8fLjtDUjIqrQ4Zf9QWAVdpPcGR/X5/EOrZ06mUEk
WRw2a2dBvgaTU8wVGj4MVo3mThlZHM16xFKi6xisPW8GNgvMSeNwsGSncwgnoOSd
JF0RrygWLMtnnz6+v1uG3NUXlx/CgHzg7uDvafz/33a8JQ+7zGH0mWizVWolWbWV
tYVqmB5YMr1BGDmr4Wws/9dCaNLYUAmboVw3VaRsDwo6q/TvF8NgHIgf802G0gVx
z/vzIVIqzF3t3oUfxmQoS5BwoZR5HWvC/T00c2cXrIbMeDAdWz9a7FB8hUcsm6G5
p1Rs7/zvx/eZS35g5Z3re4PLjxuDepFqGxyzj12QuWRKh78inAJOrN48RSHlsApr
BNBvoxe81Lkum6Z25p4Ll8xjq4tdbL2BnbWrMIyeXofSje16xHxqV8xtU9wOpMHA
WOElQu0wVzvMZpFbV+OipPfJlVbzIpn3QcayMfcw9Dq0nVlxzlzEtSSXh9s3RDie
5k/BhNHdKuAn62D0JpNFqorbn350jyHd7DflndpCXwL9ej//eoYJT3v/CWyf1D4q
T0LqEOod8joDfiuupjp7UugZfQFUVWZ9hGKV+QwUnXK1lLXNkqa629dRWbugVU2M
Z4gG0muXe3V+iAEnGFHkn85lld2+a5fUvdmvXotOd4OwcZqlM0l6Ccl0p1X1bf+k
h0QUFaD9Y/nNGYENGcMyvFb+/UQG2/MPuzPMxx0EbOBah5bTXXpWFNcEM3Ysp9w2
56MHBc/ODlEsuxF5i0p4ZRLq8HiMRX5J8m06L9cElLup2PYoFpXzXpHtsAZXkrKT
BOC740cQXVCuBnERjUJ9LEiyJLUsW/N/8o4iz2caaSq5cnGvwqiLCDBQBjXtTIar
xnLgY39Rkuh9Ss8vW5wvgL41NbU3jpfB6ooILRWpf7joRwjzKzrE/wl3BObOCe1N
0jjdv6LInCw/HAmdmoGbBZWUHwHguId63cgHUkWdqxTp7koS4Duex5WHfq9+g9uE
BaPYtjlvGB/eqTE5bGvTfvu4yrRtfirwpY51M8Dfcd3KrxzB9kDzllb3B5XT4S1L
wt2Z//AesIMVb/z3fEU/2Yf7WAUrAGtvnQtHA99A6+u3bAFyr86eVRwfHpriKiZW
EHlS7mfDWVIzNO9rqS9ru647om6Zb/7SMaxnuLnQTvhBKN7DyK265FQK3xmRk48h
TEwp87Ly3m8Hn77gepqAf/tAH98U3gYzWy07Z1Y34vlhaKCGcs9Dxo4EM7we1dgN
VPxGm4Oww4Vsy/ODQzpQjbvl3sC4L092CcheNrK3UNodmWkmOjK6aCn10yT1H0Qu
RmOC01oTyWXEWVf09XpyOi54RbqfwCfS/5NSiz2mbzHUGS/z1l+G/2FJL57J2COQ
ArjyNGnEUVlHzDRATcUfYKMNwPlco3O5TXnMLT42D+sCdoFhx02otQW/KgQCHD3C
L3tsjy0QMx0vibw1isaZwWBB5el7gaInkvn6io9IVniP8BYpSBncBhfFnTL1wpwO
JMKN53QaOKY318bvSgAEjMeCa00Itkk91el2aeBi9ARSvfexvRrpb2Z5y0xW8Okg
2a4m0yQ67MkhjjCPFrHYTxtvCRuXQCgCBxdhDcu2P+42F1fJyfwvhIz4itfVhf4a
P1WLQXFQIafbz4CpyEbQqIdL/EvwqqE1b8Mt71A4B2Gwd1xVk/Ai37+jgeRcIlxi
13qRBReGfWu8tns63rH+npUxr53fMFCrZWLhxz0EM983Kc6VerbNlqsYqrBlGroS
3tihNHY8PP18lpLSn3j5T8HG78if0SVTBT7HjFkO87q0d0rUZDve48yx2JZhR8n5
UbfcajztCQllixs72q/n7LuwfYT3BnL5qSXBxSuGT9tsqROlLVuFOdDe2xnWtlrK
Cs7sDPUhcdQ/T6p+z/evJ88y8vGCdoI8Eqqjd/tOQkiKZnDhk1RnVRVi5P/QoOWd
RRHghYWcwbxwzZAbT7Yv7H6M1pRIUqYhF78D6tTKIMu2B10VXODHBYqu/Dc1kzgI
4t8U5VqtpsOyRnVOeJW9ZpjfPLe1fROdxMX/CbFvIoD5C2nGXNt2D/Olz2SGKKny
nmxdGYFtc+i/vC6mkBI+ADJHehtBO9p5tTnueJqTU/wUoflyjFB6pXAg4SiJ3SxM
UGO+7bIyMkwoIFnca1wbOii0neBjpFD1tgTmSF97g2wZfe6e/uDSaRHfpreWEl8l
298EedacwvDh4ggADkR5eVsSBeC5bH7xOHxD+S1KvouA/hhrKxuXG2gkH5Gz0qPh
zZ2ireJAqGUnFcgBj7CSCVkVzYOS1Y2otTv6t56bAG0oOWCIyPYkjol60FDhmNPH
9vBwokFWxaHRgLTWq8H4X8lZ1CS4rtjaIj+J2JrmrWcJMi2QFsf52z3Nbz0EIZNW
rIXwRi76tJsjfhTNTLmyFS+aDcigSOO15J5w0j3F8J+gb8OBeg/KVg/yB7vCpYPv
9HkBtnciqPC5Djvxzv/jxyBY7xTpt6mvWwcJ+74KT6Go1nwgILFZIFxwiRitr0B5
mrb2kQtCUDD5sBTdGavuX3JIhQESxgOc/RLlpIuk4/JGr6LxmkF1bv5wrBn9bVm5
UMJejkmtqwR0AoSB5aRlQFI0RDDpVChvwbXiKJDgzZaNTrb7khLZqexruGbyIP/5
GPkjkYroi2mSFaZcgLrf4oW9Xc3dXtPIxh4Dy6pr8KqU/jsXjL7vD+lD/6Xlm4DQ
cMK1i1Jz1cuOpmK783XDBgEOVKX49DTrz9bPl/o14UwxMUy4aY5Vz4B+nvVYcINT
XyjqPjxqfsveb4unt+WZDw89jpycaL6ro8WKzwEpKIET6Z+Z8gVmeW3ND1FyYHpy
efLR5NFbqVL4T+zQXxuuOrpRX1pjxuNi95CJjEb5yhWKBzBFJwJq/HTTm/QdYe6m
n3/ujNcHS4tbYtMMWI00rzm9XszxmP2Ubowm/A53xh0eGrE8Za3BBtlzouD8wDhI
4QZZr7QxtwBNuZ7KXjmM/tbF5S+E8dV33xEw/EXO/c1H+NFkB+jAz4Ke8/OmTOqO
Jf0xGF7m65jRFiAlUFOWUqn7wPziALY2W2rl5OLQc1MsvjLeTEi4ggWeWO9XwpPN
593txeL+Ols0yhilhq1/M2G85wDtCq3Y6GQWumpuNgsQl66ciYNZ4PF3DCUTQSme
gLdRLHx0vC99iwszIhBT0jz1rf5Rp+OH7vRAkjsqA74ABPNxQOpZFcR1sSKHJP7Z
vyLIeMebeg6ZwcmhCGZ3anT8d5V5Q+3jv/D8j/qnKnZ1JErG+IRvT7gL54REsmUE
ksQTdSzzGzR+9aGLY0WXb/FPdr2Sv9leSb0ivSXinPSQAB4jeyH/U9D+Fnk8XVUJ
i9mYG20k6dhKUzWeX6J14LOO8J5O2OzLJgmPbLcJ3SRoEV7na/rDrnYNRm1Qs5LB
LzrR104jB504pw4hf3LGhd0mK16UVjvgRz0ItucTmFIsMXgPU5mDMzhb+F7OQHUX
yERtQe03l2MBnWAs3x65KK4K6PZ79CtVnk9HPavRf8ULaEd7erkcw71AlXvPTctJ
eVNLIdRdqvjjsJPye6dA1+KgLdLJyZr1k6PANOifYvRbyz5VVbZpZudDHOB4O/2Y
SCzO7i1pHWKcomqp5bCzyXDIBOBAlYZkFqReOme+hwGCPWmzkrdYe93Emyu7nKbC
EZRHPqCV3lRUw+LTuIjAiGwQaUDj5oFdc3n/725ozEOrw4YzFovuJYNU310W4dSx
Eqnz8VozAjKjepyqbRkJea/hGdyykVhXJPFlyQA+4mm9qp0+ZqNqnz2VG2IFVTTd
jY00NyGs6bP0DIKJ575z3F7XXJBjSS4AlNxi2/F/Jz/C7J6ZAhpmlgbsYnZoWba1
SRoYEM0/l3Ln2L7Cpi3/h4aYVynz/4bip+gO8C4UJswePvuVXERrgSfCA+y369kg
ScHr7x9ymmHZdWwT/QNmON8/gu9gKMtHEpIXREXpUEJznBN21wPngwwFOYMgsyEq
Cis8ZuxbUD5LioPQsS9KaZA0/gffO4sB6H+St0qPTYJl6PCc8zWTo4huwWtVaUFW
4W6Ak2/a7OFFcgM/6Q/pn3Igf0/qO2mOljc8FeoezTeHKydY0tOzXYr9nf42hv7b
etxjAkkq11VIAcB1XBiSIeN9JEcImKtsKiee4PcAOMoUnTbiTrFJ6/IxCmaObPZT
9fsGh+bm2x4wIvOvUipyTzUkXB9eE8Xhmg97S1/QZUouhy/vTPB17gzcT3QYNBqs
9j4ow6fr9hH+OMpXf0Ts8qQgzhTTpUGLCh9C3LcZCYUGt/InkRKkHnTDEafFHEwK
Pqlp6nCKzl06FzuLckMWxdAL20BsSWkKEo6Lw0iAJCoDl0Ru9jnS2B8b6yD3Gk06
0vspSq5hyZualJzTvBAMWcV5wMReXKpjxiWQsW+DtHkqF+mVeDvoWRXWidtCdB8S
p8euOY0pGymAEsZQBf/1eR7tlJxo8nwzdr+ut4OHOMF4ZR9zSOw5Tf5Fi7k2KAuq
7+Crtva9/z8hXXPjyfuvFF0kv6nLMLu+dGhiwtdM0Rv8g+MGdnpQZ6vBKXWobNGU
RKfKf1KrbAgibDxboF5gPEuCt06zEynTVXtQWzbWHsRXg8ibAB49aRBkR0y185qa
hTi5pa6OnWMroxkVzhPZCJJch+xo4L9vTrEUc39dkrFAJYqhtVRI9kdTmanUmV/g
vjg5WVxim2mTFnkz/PQi+gPRZQncwA4Gv/SP/UxV2OkCaKa6qfIMbnKAZNcdhE3M
o4dsngE4rmJ13oXDpdhbPwlaPjR2YS0pb7TrbbhDAQimmw4D29jZqGYIV3BeCFKL
1sjqQSuPBcq6qa1HdzZTQXfMuVnqFfAvZ57Wg3mJChJUAiju82HJVRcrvxHs1+TX
Q7llqwA9gxmq2kYS9ipejv2TYcFX0YN8vZ928NqDJJCWIu/andBTjPQXyaZzTmY9
YPgS3D+r97LP3SFD/vQbHiAyR4m9MUhOb4LEz+yVFjnFBKZFZdi4pzYlpRD5iwjN
OD02lDE9comXhSam5j54hWlgrlBqHuQnQoU83JJB7RgRuxQrPF7LP+uRkH5Nb9zE
B9ts+4ik6a6Ekq0Qmn0pGiVFQTNOLBoYNRzSC4nRPY7Ecbs/1lTgWwpAGzTQ1RWL
/tMNIaFHsrUVPwd3vQf8H3daouaVBQeCMbawd0E3WRZXUdalFn5o4U2RnOgvj26M
IVaQc8lb0Lt1GSE4K+OJ++MQ/ltIEz/EWPlompp934pqQODy/NoHe3AFBdEN0qfS
aV18JGIKIY1OckD2U+1xXYesRPZmDX6LLvp2A1wNBAym46E+BjE9aOAnl7HyrCGg
tE5lwd7MJ5B+eSnh9NvaN2THrHyAFrn4xqGEAp13GuzAfLVtn6jOZPOJW0wOgdN4
KtGrwiuXP6KqD1itJ+iCGH+p8XRe4EnfuBI+o90kdX9JbO7Eecl0eOrmHW/6HkjM
u4ngemt4ns4vCXwMxQPPgHOuPjw6rSK3aAbT8dHEzPnuK0xEI6Uz7En8lZtehN1Z
gteJ3tABtK6vvgVUT1UDw0Ht1zoZiSV4xsXVfhdA6ZwQLCF5Yw0VCVl75fIhIoT9
Rn8E93n31AK9apCWIb0VU7hxlMwepvzbtCV7ixBJQD2QrzQWUF08dG3zeSTWm1hq
rEmWTtUgk7FA4qNRC7VatFm8DyLvJsI9cNN5+IdlONULVbSGof7H6ZL8nZJx9BId
9X6AkewYQbB4+LNTu1iesuEqHz+8nbcoJ1dEmqo6jvStf3GR1IrT00iOGrJw2VH3
dT6tiB+VQLyoo0PP2UlhOWROcJeZgZE7bYgQZUQF+26WKWsi/eC5AAuATqFtljxY
MnBA88KOFXq7BmhWA6wfwTIjpcqC5reaamcIAmOZdWdZxg6wbxekHUzggStdvtFB
Q01cOfBFc/QqK89ND60hgEPG5B8H95W9OFyzxF2uSRkzfzUjzuAhjT2GJKcdYsN5
NbMmxzmx/D/4NPEm0u8K2VQwfzYVcSUBhXfR1YfE0qR0O7r2b2PMl0pO3P7k7se2
eySEmlyFrM1rBfkYZ/G9oBsxugwYvxvtFOgUqa+SzM0LF8/6y7dqKXIUFaiPjd8i
V47ph5qnh06ChBwWKjVcAQHgH1xfvInhSYEGhPRjmnejw0IyF7e6/3CqgTXfMORV
CGMoc+14KgmVa/0nmmVvPHd1o7sP46xkri3kqGBu7Mn5vcnw6TcAhbRtTIVC4DDl
k1+Ty1s1c23FHGCQbPmS4/BxzYjd/UUHerXZr0PUIYXJIeG5+PV0gMVJGeTwU+z/
2+wnBJcC3f7D91hj14OjJybDB3sL8SCDeBauaPPTtsnYtYTW9fYDzpouJnXrZU7n
14ISxRGW+mq2hmLYkj1y7LzkoAcz5PuyVusvDjaGJc5leNH8IJqMt7I+p6IJXs74
wtFZaDzAGATvzW+cvRxZeX8v72u6XyB6sgpVM35tIGOaTHFWQshutVdm7+miqBPd
RmdHzmF6xG3XZOCJcG0TcBGZaO+Hj2q6/L7bBBHd+RYPokrHYXFU+0M5zlZ4KeMD
0V2wLSa+GrZ3HN75ye++riaczYDXIStzGBh/ui9bVeEftoB0U37xbj+8qc72ZmWG
AF3hQ0EjfwBnZsmop7VkAJxbEIBnzu9AZtVEDwoZKuoX00xSJfrOkURuK7R5VmLp
uDxvSCjImbCUBDocKHnAJYFLdqsvd2gFC08VDctKbyuZ0iUY+fmKNXfdmGyMQFUG
LNyqXhZUq+B5vJ0cgOX7n4v+gVPi7s9GfmWdd1AYD9jthEdLhZNfplaOlyfEqp3y
z9f54rUhO1Nr3mHpNk58mj10b5h67afKFzjC5PIRMH4RQsECPQOZCvczba90bk9k
pi2bqrrLOfT5q6Hla204UE9Gp4/nRParBwop/KFTbM4JllqFYuRuKH2dFJDWOciF
C8SEUDzVK1tcKxmxMD8vrfnmOuvy02FSVuLQZtxSD7cDIvl7y7Qr3YB1zPQoaNVs
oxZmkh3cdj6zxc3soR27L+fKkMFxRR/ZSqFbg1kLiVz/wGMc2vDQFfO+zpLWov81
XGmm0xJw5RNX9CNGG+phYxqFs8YgRGdOGcrZTwMhcX8ntqYauLMCOJsLm4SIx7Bv
d2MX5YPfqO1f9hNPM1BCkC9qMU+tJ6u8zTmNecAr4pMuSRrmWRxY3Eu/JzG5o9yM
4860KYJA3qj2+CVo1W6Zo15rFbAyxK2pPwEXnsGMfUHQM6/h4oMDKoCShO431bBB
wBrxtmiSgfSgejIX/HN2hV/SilG5kBYUE9AaIcEz+gMt9R7avAZgTvC8XcKvG0jg
2TIHlg7SzMBdWfUl88CMV35rWjpqI+/wT3ssmc0viq5L0yg9pHEsThPqm7oTNT1J
t5kcBpFVg5Gqqk5dF9cPJC23XEMibZomqoli6YuEPJWfj3ZSBoQqJ6bIqGjxEe+y
tlK8C9kr2IGy6hysSK8RGHJPw+AgwWzxq/Mm+KBJYa7E3ZcRMuVd8cO9dV4u+QSh
gBaJtRuDmUyUIg2ccaHT3BnDNWBU97gWQXyvfY5aP+hrNFWkdDPppnH58GrSBPUX
nH3Vhkrkvm1G0PjSlhbtczCR8XonQTT8ezDr90JlqTiQY/mkhEQ0k/P53Mx4XZWA
KscilbtQ4Nz32ippfRg4rSra7DwqQijH6xXTEi0VviMuJDI4cbnqodm0VH37iWDe
5f3+MaZWr9Da9hIt10h037t8dR67UT/t/GAVMP+eC3l/eHIIVzeZHUxl0GFs5/J9
jKlDffIctFdLyrubEHvyXspCYP4c88FQuN+aSRMi+qu3l2tnMpUqusYWcbbxwh1l
f+5QAfOorkSNetyjcgrsyFiy0tta7Rs0UnpfjivhAB8saY+FeHz36+FH1NAjzYx8
ZoDFTGJfDIA9Iyt/FGONYpnb/DGmlDSzsvokN1fBd/Pns1qvXHEA7kpqxy4PzMqG
99dldQp20goMbp3DGxTsF9zcrn1doq/F8qqvdDWaMF9pQju2IGKNtor50qepx0g4
ejfsvgJcYp5K5JXqLhD8bcKVaSr0vSy0cFyimMxeqffhARe/A5KWiEAOU5E17Hkj
eQgIRxebRaOxZuTN3SSGDYJZIrjhGbqoniPTI+v0cRqKJ20576/+oNV3oiGv5nUv
AqZphXkDPAzrMV0R+cEdwxTt0324Y9siI+QQV7w2+q96Xz/mWUSIKxTaEkdI42xp
xtoVcAoc1l87gw5I8fhoT4jcn5OZeNE+9fvuBTsw308wpK4cGzeGpe6QrogOYyAW
5qaiX4RXRhAgeuHZQP1Q+AEKyZKBfiwAWJN0dnF1BShXR604z9D1YG4O6caheU4V
g49YYXAsTUyGbVvyRRwX30l/B1Ksz7R/w8tGehYrrs4PMknQyXqvb7B/tCxpSmvZ
QmbBPSM+eZcY4h+3bx1WgOFS9wr7fJCK7lyG8pl+Y2iwtyMIhszHqV1rqh9C2K5m
697j1BYtNYT2Uc3fbfVTMl6Oak+8oqxXLMXzSOQ4VXuUD081i2D4VVacTQqUjuOy
Zqcisb8SAtgJK/0ovt1RRWJR6Btf4FlLOw54sYdHbK6GfctjXqfggVpmTmzNBUA1
jAfuVDKQ4CPmwRh9+/Y9M6v4b933SBWbWjtOxxf3Jkt7GDJjbkWQrLYuST7diXcA
Fm6zElixRyPheiOgLqHm+zCvs0DCBIwT3iy44UTMyXpjnqtkfwj0fHgSQ2O28aMH
Xa0pW5QCT2mQwhxrnu8Q6rhTzXmaJRMY4dHa0kcLXeSXreXXQDLZCchwb/37IYq9
xYAHXzxgLr74JUk8qPbHUvVeY3BRgcas9nns10XtM4ydeAcH1V89HM0f8SzUTQu8
ajbNaJyYeujBPYCxFDuMETIVh0SL/zfj5EvkmpkEoFCnWkTSfGNAgtX68yLsknH2
c9CTcb9KMy8p+Hkr4ka6TIMLTqDnsqJJwW9k3/cCnlsyzop6Hs5DQ+veLh4OJ4cC
BMAqiU8eI/uCn44BUpwqB20IIDNuxSVoID8YsaD7iv2a5A2e3sjcBOEqVJrp0cGq
qWA6n1eb/z3gEHURLhzcSXAKnhqehz0BUAeIjBG2Bzch4eKrHo/SQwyDFQ3F8EaQ
LrjE7+JE5CwKBRU6v22jv9X8AKJeymljm7QzfOZRuA5RiATSfXQcfxM8wLLkHgRT
JhIZrPZJwtmcR07jsRlk5xraSDW8LnfdQkld1Feva4HGuQTtZbjYgDngwIKpE4NW
8XO6VxwuM5657h5R5WGZswBxvNHWcneHTVcijoZJPAceUsMH/Vbh/IP06D1n5VAL
aJKhewaoHkFhph8IeJ7teKkU6G9J7EeQ30GhoCCfE3/4v1/WchS/BVKOZX8ub/Ka
kszfGTvjDeU3Ki4WgcKh7E7jA+QmI5LUUIZ+d27rrSk8O3BCgQDzNy/dG9TfKtvB
SoXTxO++gUmeJ5FlFSh7m0a23okANd1bmwr6oDRKbAiCgGkkGVv/X/dxCkHAoH9g
k8HL9qWYCG4uu/MxJyuynReTIxgIbUmeZzFS0ynUtTQ8YkFz6aLcC8sDIzn1KS3u
wy7ByxtmHPi/MZNsP6DiAYFRRVqV9ziq5Z74OyFgtqa2DR0r5kYmcRNaMkdzVPdK
jZJioR3SUsWjrEiKaGoPklK0rr7e4hVbYSiIn/Gm4MpEV97mag6kdzDpjSPybeiO
Bl6NDe+dkYsNCnvtyNUZi0oQGfAbvhweIwfyd4aNRm281c4Ysoa1P1Xtpi8q61gP
TnZ3xWMlV/RI9T8ZiejxCtsUrODqo75X9nmoJ1Ynkzw2dEnn+yAACYDDn+2s8y/u
zywjAKIYESw++Z4Szqhu8KMTndWcn7O2tEaBsrx2K5NQst2MTdkPJ21bvmrWtzHJ
gUj3LBXl6/968OEZ5X1howCs8YS8MVmDeIsAcLEaPn3dydpDYhd68mkaHZOlVq3V
Onh1yZhHMo8efemtSloj+v0tDpilNiaKNCKDqFGumUG8c1lg9K/WsIF1jN1MoLOS
4byq6u45iUBWQeHBmCtc0tNAldA0pFDiQM54hq0sxV87kJSJ5oYXbFpo4GtNwAj3
wgecnsJjyuWhibsYdVWfvwkmbqliL8mWIvEuNW09nN9s3jhX1PdPZxX6+bHderjK
C7WvS5hmxld6/CVL9x/PgePgREGW3pouFYNjQ20UNbxW+j0hbPKy8Tf4zSWT8oF8
LBTZaaNSkRv8lZP5M82qSjwTN8BWtjekFc0bjQsyWvk6oJ6abIQpFkAxuRY2ZP/w
l2VIEGpOM1ox6KqDekJSdybszcQKxJPwFBX5O9ekjA4dGdQYNfbhVAyBUXV5oPQP
+cn5+eyOQTiluMuqg6puGq1/Tm32hg9bLc4Abx36aAt5gArSO20TP1H8GOjKcTPj
BiVX0g8rrid5vxPafmhPsZRLWin6IHHzGC1KKUKqIdWgYxU9luo0BKcsXKo+iTwP
HyObiMoEYdLOTG5g+qat0K0N/1F25IJ7+2FDZN0XFPhJ5LEXAjMeW9LuJl8qsKNH
h+3BPvjiAGZhdW8zVOy3dmwenr9KRpQe8eqpQJRyAS/Lene4PK36ZbFiS80AC0EW
dpMuE/JF3jpO6rjDqkP3fC82cVvBRzrSKyVFPzNjhnjlA2rgzCpKY9TJ4OzIc4x4
ESXG0rbu4n3uWNc1AZfU3nXhA6Neifyzq/j5FeKh7i7zpYJ42PId7O0xcWlDLNw/
rqI0cFW+q6OkjUFPmTLICNBYwKDPiZbrjpnOAg06eibYeS7fVlTb70HRUBW3eJ3M
xXW2D6SnXLTFDo1o9PN7pNpQN57RjowYLGnh3l0lc6QWfejHQDO2QKlCeNXXH34q
/524czG6QIrFpNYZORkeKrPWSGwTy4ZoAHQGc0Po+0afTBEFM3qCWZD7wQq1LGnd
+KnkRv99SdsKq+/8iOGu8+XZ05YaOhXqEt6a5niUT938bMTnKDmO1zsNvHBm+ETz
SU1auJfVw6vwZUB8ISVivFS5aV0RMkI0GuSVgd5cr0wVRJIrAzZxn9g2WgZlfnEI
WFZ/l8MRCV+ulan6RYm5NRrsAY+abwwcHtpSa8jly8WYHCipQqp6l6cEu/yLuNBY
fRdplZP/vmZaGcSXGq8cGPjziQkCN8+Af02C/zXAO0vSecqtb3AEmM2nppEtqyWT
FxYGenU21rA1eyhBoJeSHpmBzaVpsmLKyxuK2R+HvjKTBtUKOC13hp/+PMbWIeQO
RGqv2Qrux1q6G711EV6L9HlHt1dbkSA7BDSY5nkxqRqoVtfNXbfO/9uEklzhqQXb
r4VMUL7ApfmMsDlsVLmFGKKgsjKuLaFYesWyRFgTqRBbFiqSJvgt0iD4uQ5Jhu3F
Za0NNhJA2uJkoxxg3VnJY6F6hGJnaQVKe74ipa0tOdYpVvr7SABGMeD0X0LsRovX
l1p0ynxR9rfo4cO8F9GkHzG35EFpPA0ejqchqiSsDEI8WKUZaohgg0+bIHGws/IQ
0hGl2SSN/oDRgoFsrtO1f8LUAB2PLr5flxnK9oyqoFLF0yTq42sXpvy+E450H7/+
bnIFqNeELupe9D4o7pVhuYT07Qu83IrnhTTBf/JScZBizhFlhaQnNfJqnHmchf/p
BFD8m/4/DbtFKsBw0bd3viwo1J5y0FOqNywyNrMNGjRH6xAWWoRYYfrc2UIAglMu
42dmMsxLyegbEZmhhsS/BV4JfjpWMhUYQbNSQYqkYtwWOXOmu5l/n585Fn2iuSX1
578IIBM/HzU1+jkzTuH+oK9jYAhgmtGFCe/Z61+BEQHI5iBWIsfGHK7U34XZ85F0
rabxsPC3oyu+yeFWcCMmT8vH05p+P743Rl/m03HFdmjpePGxmFdSQ9gyx2zo0DV5
uo3SCknX1uXDrUO/KtYrq0lNfzWR644rn/w5RLcga+ro2P6f59KvU8KgJ2RBwVns
ot/6XIToxKSahTbouXSoGRvewtUlPZDkfZM7QrAm+gl9Y0omzO72hE/lQwsMpWM5
0nAFXc5UgDy87dR2zO/qpqJbhFzooAimI9VciU32CQwze3/XR8wmhhR+9810Ix5D
TYUXYIX1P9dVPhUjWvu2FR9MKtJ04V+k2FQKXyTjHMgPM2xCJpETkJYgPv6p/OCS
wVH7PR8W+z/eu8/8i9eL8G8fHGjYrcM9u2gcgGkHzLKp/y1aHrs1inAa/ZLYbbiv
p/vCeoT9O5WVLueSPzQHCh5jEaJj9p4YumqOHOMvM882Yy+7BmZnl2920UMtipyv
1RY+KOqKVp0vhO8ED4sbrZVhutC6yzHePbZpPBfDdAIHXRBB1q8tmNh8d+LWVpAb
GVZeg9vzmUHPxlTGlzsc66Yh3yfjhv1lwTg3ThE3T5mG0eoc97AMsv3r8Ah00RAY
ZYEc+4zYavFRIRfTLQZPi+5DLTaFLjsQWeaPuuoOjcE4yIw0kf4QN2cuFts++SGO
oHWe9q6EZ46d9W56tLMqHz83wGhLXuOPlqnKvWoZaAs4YRBAmfsGd35qh9zGfHQP
diklIyo5ClCwTjndj9PsoCkCmLEleTSideCbJ8y5B80CNEQqsB9zkEaVsm2ojcxV
I6oyg/9i+VkaTCxfRGKJyids9aaE5uV0UrP43csg2UcG3MuZxCeiA1rALgWG92fe
U9ZgPY6SLwKmdF7SmDbueYf7chmASsLJWTACS7tf2kooqenJtxL1G4bhjEniDV2B
wMCedCh9LvzDtt8GY60z1hdVrpc5SPH0med2dgNRHTWyPxoN5c6tm9vghdZ99bJI
sIVfPzmYxLw622F4vMDof/2bDU/f/9qZ+slLx8kRtMT+SDAqK7A/F452YIv5vOqe
pUUauOAUhkXxIx55efwxSQg1Md1i0/pdyOqynz6zmlSAFId7b+DpzX+0yquuNFGi
d1T3RCU2lNN0alFnjV8uYgfXtZXuFoMDMCQrLeJ4r2kXSTYfOh9ox2sfc9jdx4Ia
9K+9Lv88aAjMMLOAy10KVxKBfYfUI3kBn18r5dJgh/tVgc88z36gKxtADnUuRk4U
3hTLbtCLj0brYqFBGypdbmAAbnb4+TH6N+40JAhnniVmH51Vlv64g0M/mT8p7iXN
0s8nDvG+PF335DxyXXDFfpdXZffiglhSMmHIHsfW+LcR5neMnYlysD/H1whW//yb
xK7jm34D9pfHP5cICcF8kRd3G55RDSHYz8JsqBhGD5JX20sQo7BscRHBbL5sVoW6
u/jdt+VM9ZEtP7v5aSoXUombZROZob7w07rCGv+l94wIp8cE74hgTumQaxrMkpCI
/KmY/dSFrDG4jKnbIr3KHBy2wT/fwf54CNZr5jJN8vEBC2Pigy9A8MLNe6w8lTEM
U1SOfErxze5OkWgMranztjOnOeOQeE9NRTErWjsCiYhjMKn8xLFFrY0JHB7xKiZf
bmrYOwRGJnoaJwwaxp5iFsaYVdAaSsAMbOey3Nt85Ng/d/WFGn54qvLZMxe4YXUx
aXnGnE92ttCfnCxF+IJfFjEwzurZuzjwhVDiIzAT9f4/rK136YZg0cRi+UZoiQwj
n2aMArRNB8uDOnPA3FdumflmovQBn7fuu1mscAivuel3jaKC3hcJahIUtK+nu5e5
rnQtOfYmvDiv4oPpF7XROKYpqGLTk5p0y/5p24QvDl0IiIKU+AMS/I8JDlyC8p8/
bMJu7NhhChIZJ8JAkrXZ3wsoCyAXIxJPixP26jZRvfi9777I/bnOW1Fd2BestgfN
ky+WOU6MGEZuRmkZDXujCLuVkrsnO0YY+InnIyK9WcjFHccLvEXyyyQlEL1O7zXl
Z1nTsVBjnVe10PlJdo2KEu2UEEQ4P6f7DxL6qsJtZaiiVM3h4zUSXPq64KU+Xicb
WQHZHojwaQ847HuHgBxstbjSAbG9kDNU+ToHlUtRib3UcymlMz9GbfXbNTabXjC7
uU3TJZNMsg3mgMTBY52W/VPnsjqtxK6fZJ55263KBVWtVIsdDib7kiRYL/ofjmYY
dVJFugXj70Be4GkjY8LZ0xGVsKtxiDnegGQliDCIcaO/s7IL+FB5K9QZXYDjTHPt
BIvzjcFEGZbK9em02pSdtdplz/61/mDF48abTiLIXnA7DUy2wmzHDuXnI/+MzlKe
p2JlFU/tWgiu+DtpVlzrTIBYC8JMU6T6RIbUME5p0n/a2c4tEg5ZkhqGCFxeWrEq
DPQXw+LxaoJSspNYzUKIRC1tx6mdeeKF/NFRlTNDnPUAFABlZlCoj1Jo5LMi1IB8
hGr7PG9DPPIiYc1RJ2wSBpQb24R3Yyu5EZJOS45i4fGUziIpoth+zrdwhcIT3DPY
csKc/pu09yzu3f7FWKRy52sYi3uCYo0I1KIoaI4+ARORkmloZexFrbpsn6G/Nixv
/I8brDkyzsCJ6qN5iwQPqgXxAv5tXXu+IdUb/3b3QNxK2CwxaR2LjUFLMfhSi+qU
xmII1FwYYPzwtV1VXpxjJceth2dR+i/hHBUcnT241WvqlPU7FmJ2l+Er2n6j9/Dy
h1vWsPINFlE5xrEoPpE17X4ZkcgtJdfBlHTp0uHRl37qm+R/ZAWBS1K59ACZo8/9
zVAvSEJIHgupqGdKT7QAjPDh/gBlKKouguDvuGd/EweM4dQhDisR6Hklu8l8RrDU
QhsDATRRb2K5Vrjo+AQ3kdtYe7dIt6wTg8ParyWxXdnArT72ngZFv6R3JSsbaRP3
up4HbRSy6ZcTIOJRdwsFlWBahcM6BR4IaDqlvAkqYws+uqMVaD0uQyuN2bLnaAWB
GDvZIDjbyQnZsyojQ8jvqeTJ1huvVHLMS886FtH7HTZRXMFfBbceoWVPP+mlZovN
MtMxUxKxBzusFKYc+tz1GCxMXYLk4vCepQ+rgvNYdYhPnsMbEBHeNn4bZpieZIX1
D5W7rc+smj/2E8sO094eQVAuxXz9xPDR/kGVGAOGwnYi3AKWBE6FVBThzzqUvhc8
mpnJB0gcaj8C3hF1RP3uW5G0T1SgbOhXuNrmMRb2SmiKs8z7ZUpwI6Q8MPvy2Qcb
7X0mVIg1t8mCsC/urFZ49up4d6aQeAAWEKOfWnkAOOuUmmqdIdlmCVKKfzu2b8lA
Ci+J4fOo9nZzUcoC5dJ+9RALbepbkyM/qWDqak8YOdqviwYFOIrtVxBZVyAMTuqx
ZH1tf4VoTna8tTmrJxRXcTTlkSbvR4pH+6ovb0khxkG8nF+7Xd5PCVtVvCO168Y0
Z2ykvV7YI1Ne+9odolxiNomoDdsEYzzrPkPzt7A6WuV5IUuLMgKcULQF8fmaWEET
io8gCf8R8aXFwxYfF3PC4nPsb+vqlFLu1VvoJAca1mRvQ1UWVEWQdnlXBHICLCK2
aGtoxE69z5/O64Hq0z3V0N7t97WqseGqSdJJjiW/rs5etVjO7TgOhOXIf207diTI
lpxJtyJ64w4qa/zGTFtBHJtG/V7g8syXmDjPn9rxGvCh7AXK1IUIPk0QYptpSoqB
iwVA/Z7VRxSpLmVSVy7H2M6l1oBOR3lZHarvdYjSIgD5Z6orFIbx/uqoCbRO2DMm
6YbebOm6JKiJTiGsHQ7WJBLSA6O4LcbzbIl6CBdiKMT1Y0IMfa9Ilvyioj1ZcChn
zmJ6TX3fnPulCLWq7LngBk49i2081gGXPrKZFMIGM4DDKdR4+XG4yB5+Tme9f5EO
dYE3G6W6GwKNjrkNV8fXHIgaQE9e0Val+A4ttEBx3i/19sjRO2jdMde0SGCIC1p2
+2tHh7CpoGMU8Mb7pSa13U4BZUOCTIRjA8nTSpt3y8bO35/5AqOPW4llouOFBLmB
0CzU4XTE9KxySXugKW2kuFSj2IehZBcL+fkhlAY2BrOVUl/rT8CAx7P+Ciw5thtB
+n99RKGQy210Lc66Fp8hSJSc44/kXyfjSplDaVEBuzaTFpcFF1els2VamL+oXcnJ
Kf9rJg51L0lDTfbUJ6W8bWAlstMyMiFi1J+nDnpyAu/tLs4/YgAwOu3Sp22Oai0K
K+84rabyyrLbD10JAl/IgO85Z6tKf/ZhQA/mIiqtALWNSEBZ1QSK/UmEip1ZqOsp
odqolsFHCJJtqcg/52M5hL0Ji/alX7U7u9TqpqkYsRTSiSw/jy75903fal1eH7kr
tJJ/w7w5sfT7vR+kUFGEMERkutYKgJgRmTnYcfMxuRS4g/ymfO+zWRVji5wicZdH
E4wXqvkc25x9+o2UXwXBPYwK14fXs7BeqrGpTjEmogX+Ut88G+q1+TAoYrgK3HD8
j9s/zXSfJXtXjuM/xsLfsp5nenbeNayQRCkA+rGl917yJu3+URpiKjqNNugylB7M
9TgFbzk+fH1Tt31kE+Mqvu8BAJlbOHVsHAw621kOhqni61+Hc/UVQFmIgbo//qJi
NnVhT5ukTjSR7TsyLGh3yNt8+oNf2PnpJOt0utuVIdCdX7Zz4EOLarjqwqJBxq8C
z4F/dGEmVe7uR+PMHyar2SEX4ZWOPik+O880StbBAPj9wW/+LKa1IDfF/G5eRMcq
xrsvunOKPNmqOv4ERVFGvf7q2Wwn1yvM/El0wk00yZFxHMeRPsqxATPB8XjIELHy
f/dpF6RMYlJNWjaDKgDAHukYlLnGa9mZhFbswc9Lduk9hMtG900c+Uf2+tBztmyQ
fpO2C2IAc2kSkq+7ej9dH74xll1kacArnSd9fsBrFqBeF8O4FY0d9Sr/cCbaZs2b
r4AjkNT23xYy2TvZyX0koOR/ZNgnh12YwZDO4zSIfRNwA355QewAxw6rzyFABX/J
VAFqmBqcYDA8nFxav83HO2xyqNaXUO5JKMs/YwhXuF5A5r8ndosBDXhCFgimnkCa
0SKCmtRznIL3X5/DhGpY2fDjR6Onq6exIWxBFQhn+g37M1KJ5Knz28kiaXoCUS+I
rhKWa9BBBEFbBvb8Oq5Ymy2bjGRX0jWfp4ovF0wGTwTOan13lS5AuJdvlLvdHdL7
gjXbFG949s1aScXwUg7Eebw4iHajiBtjqEEkTBbSRkZLOcoHXVfY38G0iZmNfKdB
tvyroeB2GMkmxDLr6n/RAt3GKP+EYtzxPWdhDLt2C7CgOdCHj6B21W+1nUy4ixED
YLrpsTZBOC9OxkUjr3mKiTKY6N/UOirtbCU7ICcVQdhd4uSrOCOcBwiKEaHrH3ap
lAb0JR+z+yJxAhVH5cbiIffnO29UXW+WqIEmRwkQzSisPox9lyJDjgozgFGyD5uF
1rM40knHScWk6eaGTApVitLRRlHvjATo4UorcxyHDgY5l5wXpCmqM3mf2SA8RGmZ
UTgKgUNSkz5epcGXZk1G5+0MOp78rzy5ZjfDgBVrLCQK05yWn/8iJysl0447+jk0
e30Obg25GuhXHHuxn4z+eV0tQE+jW8yfYLWoV4tVFbGuyo1a5zgSdzjge9gNLMir
VwuZI7qF+qoykSt0i1RfRupSoihxOyuMz+EblSwNDjWKzmtbUl/YSceMOAXa88Z2
kPUbD5THFxXg6AAGB6hoPbPxnqS44Ld5OiT4CgtAKi5GZDVFrzY/bar0bUO+Psrb
L0KBkGIPlysBlD9jcKrasduggW0UjvfxC01AKj8n3pAaVTeI2s+3xoPiwHE4mlFc
c1rqKDJBhhf0xfIFnu2suTTnWJSUXiC753IeGM7iulNb9VQVlAIvhBXPQ45veGTG
mL7NqaZJoMakjS1Plh2DQAIEHGrU9/i2yuXsAbnUho8npWwtSJifPC64hyxef5V3
kz7LW1ALJICg3rV9P+Dab16zMF5qTKt2Vc1/0fMflI53JpmHXy4sdGX/9VRHyd6E
QeERkQXzoImWp34S3ymx6QrNl+sblgmOG8tgzLiyrdWO/65KEdcxRXDAKbrrZePf
CpIRzT/WpvhFZrtya84WlXeImb0r3Cio20C4HiYwD7gkCQisRA9V3UOF79VlVU26
+ZkFVYdscG2byLNDJcEmtF0ge80aLFcAv3XJN2B6hHp/2NnYY5NmgLXTvzntLxfG
IWzMgV14+l/Vror3UC1cK77Z3bFdunbKhM3O8oKFqdR9106/sWBlmm2USbi8zFvx
ruDOOzLsyOYO6jzKUuzX8WT5F33RuyrogL0+JGzboX1Gy97MAK/vsmmykfvektKb
ic2a/hyrOw1n9fPcjtH5G+iJiOdYVOCwZqRCpyRoKjJTZJItCiyr4Ck06SwwvVN5
kwJ8VCtccCDIbIhQfPPh37pgn6lyKGT+9v78bS+kK6qq0l53ka87gJ/45Fpt8A4H
IYxD92q7bGeZxsxUOPRPFc+8STagmmMIGB9/907UdyQ3l2J5ZPMqmTWyGy9LpD7r
jJqLHRQiXFZotIdT4ea5umbj2dDqkaVnbVmCMmltpGQAMObfieUxxLmsb7swOOvU
aFmdIj4gCFdYw/t3icypq+ce6pKjdaP3j7rcx6WMHE4PbcsdUQbv6M/rzMr9Z4r5
IoGpUWvFTGy1cBZXtQ2Q7CzYg8OgEPYsIcU92jcNUvKRED8pK7qjH2vPAjsBSGuN
+3K+nHsjFzfKIa7eAKXizx8gMCS2WVrPq82yuZWSqXtEDIx2WQF0FK4uZ2hEHmst
dzi7raRgFGIJpg9NXOqILEo9MH9RPLn0lQfG7AauXQUb2A//mZWQW7aFeDWbIs2Z
xxEwkONsjCP9T5a7F4LlSRJuHx2ZuqwUshN4neK6O940Yd+rMmqG0YU91MjUB4Yh
V6o2kO9BPN8psMBLLUfaTm/ZbisGIGhv9XFWOW/5CfA/tHYx6C1SeEEZsPuh/JOB
gVFOM37tMQcmKu2Qpf8J7gP019z3odMjbPHgYDuS6b6XfOfUv7qMu58c2xj2rPPD
KqwkZEtpJaIZXLCBHYB/6SuyEpXujqUpEpkKAjEueNl0opnCM83212GYEIViWrYZ
kGbLln2TLLi1OyL1a5EUpoxkB6FRs92P331hPb9P6Tq4AXZUDEpSOaOQYNJvGRo2
2EPxLFWfNSRiLsz4gGlm7G0sq8xVzRNaL1bkn47SvDm/fI6LTS1MHzZg9leX+vzs
Qcg3Zc0qX2Hew/6eI+KVdlYUTf8uF8nzCnqgjlfcGqqAsTx2633iCScg9xv0gCD8
9Jj4NQJRyEBE0Moe7cScUX8w4mQtZl2v40tAQURmyfppTRnXKPJ/IWGiS3e/vVkz
Cp2TdpnYorN9KJmE43I6RFWX/4o7yOV5OhK/4/FW7thNYpUTG4ipehVzxble6AOT
gwokPTEDPcIN8YOlUJV3Xcx+7WKiC8rFqT/Vmt+k4NcWuDvzT0KHYG4OF7lLRqCw
lVVtv1lIVGuTQAttA1xS0V0hbNhdKitoghZzMBAk5fsifHB9wZDY7ngmosOplDqf
Hhq6VQnKQryQNEKnjQh7WZFnJD2h91fhEe1DMYgyP+48oW/3IFYVFXWPcc+Ljsa9
XQAf9+A7LnVeMwNnveMaOVSknO63igFRTfn5qaOi0a1d5WNwQwW2IZ9+3kmbrD5K
ufpGXc9eGzVPAR2PuU6rSEzdfyTKHkRe0Rqfo97/WQRVs4zSCfaaY2OO8BkN97HB
7qhXWYhksw//xaZnXRNoA+TZ5CzH9sJ7qK471hV+ZHDk9jpZFK9JEoXRbDfosgIK
G76wzhW4/1YggAE8rx7W2OzEoGlHEVoLLz9pu14aiIvTNzweNl/0rU33yj9b2l2r
ZMsHYN31FTBXq4TX89gD83eM9/MtEln9q4Exz+hydyk/IdEytwdv7J8qkhNCvJbl
eP/FXXsp7KC7b5nWVghLViCmmniKhmdbfJEZlXn2xZmDbqoeuky8xAYL0TzCLKKF
Rk+PrQIX5JscNQ1dePwdxQZC0bRef4X5F/MhZX4/KABXG9h/TI7C33YaHgnxvGFE
uWXHl2JX+5ry3in3+3Nh1lDtaD8mykbkOitrbuBh9UiFfEp8Bzq1A7YRHjFup9VT
71wQeUTz2EcP5O7byOBOnai6j8IcGbBo5kjM7WVeldluU4PdZAKoQIskqykCc2lw
epkSSKSPFR+YyFlQxMFQ/IWF14jTxtgks8oRvRaueQLE7rpjF69e0Lgv1JkNbuIg
nLjLuIU2TdRAicpGJNI7CfDMEyKX2u0bQ1e9NI8Y6g+bEA9wRpu3kiuIPmzC2shm
OpecF2qReDyjfUZE2KiAiuhUqBetAoHMRkEgO4ovUJwQGDWT5RXpx0EkW4xQlIGh
1VPOYS0cvFyz3WoZqHWEuCLPowKpLJhOfNsOQ3O6saov6nZfEf9xYifMW/YTBI7F
3qzGCBPcQ532wMgo1MyBLAx/q6AgTuVbem6Qg6lNeef8yHVUn1h4bckO1o9MEZqi
L0s7JDDXQzIVfnJme2jQ5AmaLeA9VasNwhFqwaxVPNMWNOHIyHGHm1RpVm7eEfaB
qM+G0psRzosRm2lgVKoW3WJ1Z4SzByaM/Z9165e3t6sahiRJDMrDVrKE5naHculE
OQUKEhN5yoq/YkF9oPbnuCSkInUgJXHRMdbFHGKyEbIiHfLHmoBn0JIWGFGUGf9g
y8DFg0gRWkvJo9akqCpZiri2L8V2Mcwuyy2719A50DCJwO38uyZRuuX+CS/AVGWU
ld08VgTJcKKC10Re/ptItwBNz66obQv8comOn5LAsYgCcs2ot2BCAr69CqMT8iVv
sWXuQVAGkCFSytfgIZWR1cHSQBN36N9lf0iauiWr3d7/7CLZeqREHyIu9QiVxWx5
2t0G0uM+pL0OJaUeDZ2UKmQ5tlw3K0qGNdcYSu+18elU+Vy7yGfIXOvOnyvXKCbY
VcViUvFTmAKIdaSf05/LLM1X4j2b3bV57uR8PGjUsYn5kpSRfT5pnwQrCN1pXuPf
PQ8tBa8E0645zIf//G7FVn5Dx53YHhYOPyvNFPIJxGTAKg5eLENoyl02ea/jI81W
L4Z66JqyrehicAERqd2Zt5zDDsThuui9Vlysxqj/leAQk7lOggtfoxAaWcvejlQl
yhACJ2LpsFJU55ScAwC6UWtC3ZzKz4+HpSFAl/X/EOnA7qZjTXZNe3gy+1lUYai/
VoNLty8R4cEjBeLOb63KZ0iNLJhAWYYr8CYOdKj8O/kl0eP/BpaUaNMFGow3qlkI
MH+B7KOe5DROUvHkNHdyBF/Hh0q6fn05SDdce2GV/xC7tLLE4O8Mx0FKMPu2vh9+
oFsnmWHdZOF3Dzzwidk4LtVN490KkAF6p790JoFvgI3gF9aHaWEKgziSk6qwYIom
78cSybP4GmNesPZAe+/8DpF/0YMW8i3+5INX3sWRZc1QVhPEGGWgMJwNwSDBTwRB
xsjf2hOqGke7+5iM0gjaQuJxAB4hiuAZNtzRZJMKDDv9dNTlahCvmxz26ybxD4dZ
pm46QL/s3l/pBDLm3bc30ndAgUTAp2giFzEyBbgXK5iWUVbARSSMF6wB2Yc+nPn8
n2F4oL4z3kuU2PstMyTmxQ6GKkDmbh0l9l8D6r44aLk/cmgCREoTOaVwUM+O6sZJ
zpwjLNSmZnjb8MURpEUdSOsrgmbDxOpj8q4/s0aolZGkTBJzEspoYAGxcaiq6sJ7
/cVPT+zviI5pWEqc3bblDf0s1oZCb1R9vl8y93I0yYajQYBrCkqb9xI5drsfFWHF
FfAWg6TyJ+hIoA6VYL4zpAKg1VX20/afoyi+s8WAZhNxOIqZk9v1zBLPefTfdVaL
tXWQ1UZNTBhPQdirKGucQsJHrNbPtLQVkh61o2LI0MkjDiL64epGmPOlqdQoJTr7
EzqSIJKhmoO5F0+ZvY67ASzm9/8YIGTw7SHqHqP7JEBgEjkaqSVoQB5nOqBHW4bl
56Z0UTz4AvvpC3lI/BlKdwdBjDNBcpvZ/GEw6Gl9tBoLlJ/WRyzgI/r083vfn8Fe
nFk9mXaEw5xM+VOEMV8CpsaeC6RX5Rnqv3aoYTVXD1GB1aq+ldiRGke8fzSVfGYE
uSa5ohmd4F2MPFeL3F6VjIeHi20ynrzhMy0bApuNBu336b42hWRlHVr/nqPfWQ+X
Jf8C1MYU/+xsXY6Imp/C9xypErDKF8uwdMGdYeqZwjkjivBNuWfss4l8WLAo4Xvv
3pVoDoTg1Bds04D5wArUXYFIBrgtI/Fc7fLu6P8zSwwvMThW0h7nLoDGSLAlMZVJ
776J3T6ttiZjHtW23PuuGrBYj0pL+Q3+M44yTJXTgXgKh4NTbXzCz8mJ76Hp77Ub
uVcWZV0A+BlldefNIMxUCHt0lkrhFWQuXm7aKzFG8IyHouRVQmBW2bU0B8F0L7RX
8bb/7QJDkuq+RuLu0wFHeQoHL8rbWnWgil6cQvNo0Y67zscwvua0ywc0tX+p23KL
e9fxEnaK5swFVwrRBTzrVQnZ+ye/rnB82ewgdqjpRxAPT2ZanO9/LrFT1ZYblm8N
VjtO6lWA+Jy6K/5YeN47BtU2aORKAaKtbZcCNPSUOJ5PiFgbbv+OTQ0IixFQRjwJ
uc8Y6Us8eazIJnjCEGCX8VlZ4TtuiDXr2bHt9tlpO/v7sKDzMSmioqsUTO39mTCe
XGgVUd7qcBFnKi9xTavn2h5VujeIB0EXdUMRus8WwqBVNJROrQB6jGPGWEAvu53z
axQxCAXuXnpkV2MiIsL/y5fTBgC+hOLHid0wMtBIXZGVQ0wAI/aU3yU9u7KnNqxt
k8aGToSTbNrTxz42uizVVQvKbI0LLY2L+zaLuiJXaZBgKgiZTdtTYk5TDdLcygcv
vo851Cmqis2myRU8dRp7704k9FYQbuwFOniYx9vxh8ZpM2DaUSkCL7Fys7GGHeu5
1uAuiWIiZnGKtLibtaGGyFLHiZgh8jloP/MyCeRArkd23wWeS46mHzUqXwr3IUZX
HJIFmD+Tjj1B4+ywA9eUWKMAk5xCO8W6XON+bER4XXPTiMKRSqnm4mKJrXP7zeeG
OE2CJb5DGR2439WUe6+CXXGMFG1t5Oi9bwE/ZTXwJsjtkrrlAGFRDm/tH8zWTCTU
oyE/e7+Wtvaxi7R87aytpzk+G6ITYpHgj6RT3IGtO3g0y9fgoTnPyDe84KlMBRXB
gLV5jPUt/w2ZMJhF7C3JDpRX9n9njDBPvcMqLHwLKrySANCw5r2IWADhvyKE5W9L
zfiLCRouepIVJtc2LsCEfhNQQq8a2BxZdKXu9rbeqi0o5KrV8uSRm87TW1b5ZGab
coofXyDuB1V6SQzRePxMEXIDrGMBmaRQi5jCeVM0GGlHyVSTH+X1SGONf8XqlpGF
tg4kIJsHq/2SNeVBts6vrYV72whaQNn2b2j77qdqHZaXXnRru5mVY5ddy44RrMya
ZZtHZpg6ETE4K9c8Bn9v3HhXXI7cbH9m1LlGUQ29y3a0H4C25ubUbj04TTBQMUrI
dpOdDZDlTr6LY/S874cO4S8EcrLilmacJxhN+j4yR7xrHgkFV3FCOYH3l3DW2B9G
oUJrZwtXUz3A5sJiBzxDX+0hNVwUImsY3RvLN6S6spiToZKmiJnVOmdScJpp7D3m
pCiKcSqZqgL4CJw9G0yysdQd0wSJBMrnGaz6Z96Z4ZvRYaMY2H9K8elU2Nkc175J
g+FpgnWydlcGqOoR/q8l/aSBR7Wy/5oL40IS77qEHZLBw/MxaRkeZ4Z67I4pA2VQ
q8lsU6uCD0/i4wmBOjUUYRaZz+uu8MN4I/neiZ8m/Mb8chS4ZvMRps9AbFZ2+wot
rAx81DtL0zfmZI339k5bytt1e3Kzw4yuDw14Qpyus91ePQhIn2zWDeDL6Ukyoigg
40WjiFPT9h9PabSRRtn/LLkANMVArvmolikdO24ODyfW+4euNE/lVkEu7Wil2BYA
QWVBZYNvkCPr/AqqG4OqLzL39Vr40nJXIMYgMzPhxe7B1sPQ73EBYZh52r/aMI0P
xM9V56eR6hBWRWMTGzuleRCVMdw5MzuwnZKag7Px37xMkIHeajRukwCwGGXe0jis
inYn9/kx3n27ofkacJrio5UN3lhTqfQWo96xzyNRgR0OAxtv1Udeg0mrKFXx/NRn
4dnNdZI7YueWJNW4VgAh8QPadWlbh7xulhAws8MKV1+vfAKeCStSzFmXD6dCOzPn
dojof2AoBm1aLYgJJuCymqYLPpxLpU/+yD1K4eSxUfCqCTRervEdvNEMfaSRUN8v
OwfRa0nTEMr4KWRzDqB5cjAPBY6xojVgucljzdvhoj1ws2gBUpkZvpikpjLrWAmk
9SQ/b35NpjOhO+tZB7iitxbAyjg8T+eAWYpC1JQEcRMqsxoxCTO0BEn47cygRZWe
KVc5v8iUyM5ywxspgtObXj6WUR6VdHM7G1Y6dMtOgipirBZq15vPV5jHKRg0IJql
Ci1lNN1GcJeP6PPtVrblDLpB5EeNTBGGsXrEcr2TwHzHEoAQH2v5fEJ55W1GK4dS
/cKkk1xzus9Hxi7VbegXPv39PZuzMA3EvkyGWrD//HvLD+LXU5WI4nDOqwBv7Ih/
c+CxPPAk8Lak18XFz6Tdkw1KOxSZKuSUmGIJfOZRTnMpNcTAOL0RfGKh5XkPRLdI
K9ki5kgWFWVM3GV2A5/3TrHL1bEKwTPUW0BBmKaCAcVro5kO31s6rX1KBD+M1i/a
i/XGYRdWwG3vZvG5YclR/9nApIhgpXxPnCLt+JwLtvpX+uQI310ejqtdgG2Uq5Uk
CGG28wzV6gENlOcrMBN/soxC1f5gX1A2BjECz3tEkPn8UsHAT/gFbHHU/jjX5V64
ayWypT+WknCJjtN1uiFf12jbHw7mMfxyBAoZtKstmA2e9+anOfIYCEkSLCEC1o62
wVRc8Q128xIVlSmsD8YGRhPGNc0q1ALLus7OU/Quf938IqpRmbbQyaGwcJupNdGt
P36BGZUBMmxlcr7N40Lid2r3JIanWkpLA3uc1EDDYjruzeiQXRLvSqPqF/+ZqBFZ
sDNcjEMWnaMez7SEA7xH0/3PQY0T6rk4UUv/cXrtAqFeosfuWo39z3lO4G4oFPYT
Kh2gMaagTtnTN19M2tRpJWCe9Yl89cLcq+kRvcndTKAJE8UcqrBscc1oTjL/8igi
30o43GZMpyJxJGNAXRafk+KMI1vjlQfxmQIEdZVbgIp+9hRNI+K5wxq4W4Pa0YhO
GJGtltH0b9gaSa3vcLZ3SMwsdmvEOYi0crpkQwq6og0jYkpGNt8NjdQiVpmoWjU0
GvQkRgHcd6BrdRDsgOEombUuUUXnRkNR7c7IornMwFuiSpuJFNp0DZjvbgSkHxCt
9p02WP2sMdiasS+kxE1Ef+praNLIKpB3l+A9MvvKHe/ALSjpJtJ18fOSHYYNl1gw
qEte75mxzrn+vbUVkSA9AO1IkU7/IHsVGpMWuna0vgPbGhGP2QW2HhSXZBpgSSha
qybri/W2XTnUjJJQnOAn0i6aCBTFjCmdODyrx+YFz4FY1G9TZcLfKYQCWPy5Qj6/
8gEw5X5z7hBKe+/iKrziEIleyraeFN7TJ85p1YLmSmxi3v0HWGjAMfL2hrf5Gn0Q
Hdp06W6LbSujnTjFuLY4OYblpZ8Y5h3c3sbwyunRqENrFjXsTcEVfSTAdeeBVYZ0
bBw79FUU1c+MZT2EpLu6wAIh10iouf/AXMcuODtdR3bgDjueNo7oG+sBBWc07c3d
57QHRuIatwMRLVIzhNh6ONjAIRw9QnaAGfTUNIPS8HsXGpzwbD92EN7Q3ifLUjdc
gqFk5fDl1yHZTEd9VbzZCDWLeDv//7gyWCgaynZNYRjVt4GXBz+u/9N8R7z4KW6/
3UiVqF2q4S+rtDpepvPQP+Ta1z3AKSBFJJ0PGtBp3J6+FUemuMftNlw65WynbHQk
/cvejJh7yt9V+CLsHZWYJOULMEBjuZTqw4jdZJIx4DrdhF5N5J2a/TAdnhpeYhTe
wQXe313rTGs4mEC0RKpzr2vC3qfetuAOXcQyi7PYKlajvpJJLG5zYslbTeCZtrWa
IdQdEARPy3Md8K2XA0gOjefuIWpvsNH5UHcsovVtFccodm2D5pJX8OvHJsg7joaC
JeVpUK6WqA9Je1bv0Gbllq18vPRORPGRkRpSFKgS42Td/MZUwqRHWRtrFyAFlNwa
F0SsQaMa45I1+qaafRVBjcMUdvXnBaiHxsWR71qDzOL+Y2yKtNShQbE4PErsQLBF
VDuLHMRZYz7M7ldsqTzidMhca0+Df5BMC0GvQmu/f1CfPPPAGuCxmp6Rc9fOKAzw
OR7SDuAp5d1uaNtNeGeUwyPVfZe+Xr6IarXwsuChfzgh8pBlkC3hxxGh6dvlicHn
pY3KR+/DSKzYp0NHgpAeed7Tv4Rgxm2rUN/2CuZLsAr5muNstpmlOkFtod8rVg7f
KjARPRozfmsUYfudXfYXiYN6W7H5aAcIAgjtzBfD3GrW1YNfy+x67vZuYCLPFI1I
QWMwkutTFB+WVv6l4nEUqIxvw8aq0ByFPw/xsDQjT0/Dp4K/XSu40ZGWR3JwFbhj
fZNluILBZpm+3BVFgTxBJxN+HVWxee9i20c08SWIFUIjGUSw+R+MYhU3xzK/7sbX
s2Q57UvP1d+JbuddsZdwLp7EsgLJVRCYhYe7Vp5nvNefylYSTavT4PoVid/AAVja
O07JEtTmEQHeWc5TfEL7GavNEDD6luQQWDYcz8vV5D6mt3Xxd+I9jT8iQJZ6h2NN
fdpNfKayWvtg7z9w0HENnRvDvJNS1f/s54a9Ps71CN2t08JpI5y1HNGZsomiHzAy
oc97aNDXPXH/7sSNBW2hoXAx/WKN6TjKJmJR60gqdfHZHSfb3NDTDM9IwdFFWinP
PZsueGoaEvGMi5LxQyZFXQld2VWcoO9QJs0myd/WFv3OreIDqLUm6WoILOp+ZZwr
9eG24XDHDI0ns7j7OtGwP1kXso2VaYgQSX0Y4KG2ajiJVtoc0oegXKGyKtkvg58r
MfzP0dJZakYoHCstrSxc0GxOjPwt4NwTfea0rg4+sc9aAQyjqbMWwT9uTTygs1Oi
ey9LpnBm85qGrd3QlqJz35yxy5kiBIbmD5u2BhDrFIl6Jl37SdYWvYGCUTeKM+rq
fHdcFB3iIr8fUHWcGlBTELMbnTEz9SvGEt7XTZNS+Cm1zDQ7Q/jw2GbURQNQJ+Wh
qs5Q8QbJeLVxaYoqAe1emOMCg3FupSFYA7xPQvkP91zrFsbptEBer8bVyVbAXhMF
S5Ji6suP8E9FTnNpEzO4BfxFlm3JPs4fQKXifzDg4mARtbpQKHEYD10krtK6QBMk
MlrEA8gxQB32FqJR5oskrJUTZP+H8sP/bKpaTKwln5xeHy+zNC79uTzc/hQshBF8
h87ZPVnxIaL+XCAiE5/k/to8ku1bwjSf0/W1VY5TpaMDnMAICwHL9ojLroEPX/Ie
yZETWiOu8df5LAMbwtg8h7xO40Ep+eL3qkcafo+qHy0ZESANyJVa4QNyFp2cpIRh
snSmmY6x97yuXkyrNVF02y4VDDoWMYqfxz2NaVCDOAIC+NwtkqZDnOdknS13wgNv
53WxIvbMs5S069WeKS+lU4bTWFI0+8F+UzngC8iHfsAN7BfAnPybMbmMT3VZSQZx
nPxnJwAlNzoHwU01OeSrcrVqtw+OinhJ8T/0uhTcu0sw3w63/TUnoxLCPTfTdLiI
GkYEHhT1EW+j2DvZCGFBNctnq0NHJlERCIcncsWEB6vv9kDsUTBDrLhJo8G9YMF7
42TrPP7FfGI3zWX93+fzxHf8HwIYnunzyxiPcUe6YcFX6MEe/G2sPJ/znbYsjuQ8
1n25oe3UnFY+nLyuBXe/8q4FJzg8MSZp41cnt6hZqsiPNJIYT73arHhazaTbcduw
Nh/nHvPi0Ju9FVNwMTuGSa/D41LT6GmBFwdfWJ8AhdVf/voyaTbZIB1+NuZ63jEM
yR61wwsa3+QFEsfpORZCt3xKw5r0WZLp6sgYyfoDRKb3zbVJji2GnoAUPIte1oCQ
dEtw8g5qnn1BeIaq61xNpDt4HNSM4KM53y/WSDyL43xh2078Nd2DOMX1cWV2KijG
m/X44TPsOxYjXvi4SPvp5czXxbCbaQwc8i7Ycy6aBiNQEMEm8LDklAn4R7UuhiRR
84kq2XpxP5leE3VpYQROBa/zOSC8nPNT4Sg2tbbVgLad9tcnkS4D0HNn7IGPhhQG
DnzjROv5rRiTxujFZxp/DMCNG++bp/hIir6N+GoQ8y9d0XH7FbOR2IZk1g917B+V
VsXNAkc1qD/5HJzeJU9/OxT89LaQcAE3HOAr4nyzLJEFNF0Qhr54NMPQhLB14TxO
aOt2qY3s3ZM0UphFYSTc9GbtlS9OLoirA6WfDDtzaR1G1Y0cukqn1iio8K5HL3UN
TVWi2gzjMmQJQ5nt3WYZ/Tk3duHDOGo6Hb4zY9zM8x71i/OwaGZ0csakDrDxCUoa
16iLEVl7OwdGECCJBMRAJXuaRRqckxjGotoOCW2v5rfwJeSJH8I3eOZ6ErY9gX0t
4LO3ZDML6L60yJm7cPgexqppFhbnonyRmUGCLePc+Q+JkIpho21ds0m0fNNRVfu5
SXZy5LRFoTajUQnIgim/ksuKNn8NpVSB8W+3HjVAihCIdagrkLtEstdeG5xOFnA1
RcL9I8htLHWg4enm/PsqqC0tBXFxfWwoDvsGJUA+XvSMdM6ndmB1iT6EzKGfUmrE
Ak4lEELFNf84w3k7vSa4YqbyD0lSrvKXPMumbqlYUPSTGeaTchMHz/X432Hnmdi0
ytpYg74Xx9mXvT9OWDJcLcw7oJ39QNawjJcs/RAPeGZVptor+h60iv8KmNCpnAUi
2FBJuvXJPdQLRqpH7Y9tGRQFfHKNr1JQJvEi1jmdLuzkVMYjcZ/TKYtJlksnnISX
yyv5EY4Vx9y7P7iu7Yeswh2q8mL6rztFfX7tjcybrVTFycE1e5MT9kOwqztW788s
bmKudx4DzH8Dr9ZMdAX0lL/ps+lRBg+tnQqlywO160sW6JoMRG0QMlFd8JLreDUG
Mz/YHf7jw8173ocmklU8tWVkkCJdFG5pIth7fNf2qe21HPEeL2C70q+aM54ieaIb
vUfKyxKnpSr5OMVDaM6vpFLQKXNwxd1CWxiV2brI3ybXLg8z15S3E39W7ZWZVGRT
2K+qX59HNN++rR4vPqip0RZ8sV5EWMk+qIEA84qHzKExpJIFk3hsBfed8XzrKR/Y
78KiZ8OGBD996RJkXtduxVY0D2gk33U0+i1lNVcgBWKrsS2fMxyOn+mwSfvEGiNo
Vs/OlZ+QB4o2ojNRhXdjohfJfAgcM0Cbv8jSGL1Sy+F3K5Ouw6hCKXBkvKvejaZi
E/lMoBHkj/yfti+Wh+7+sSkMjd9nXXpOc7Ur9Q1I8nzLliWnPR/DfhfSrSnyx9VL
ZW/Szq+sGi05BUIgkvU9v2Jctzjotg/DQ+Ut0E726OzS3E/RHJ8w98RX7YkC4oHy
4rsePBn15eiJMZixriDd3PUyUZ6e4tgvKMCr8st4TLmSTTT1AclbqncvDkyF44cd
LUjVIVDNRY4BlxQ0mujgmFQBvH9AaIjKcQtmIBQxKAaqb6ZLm9LFqcXWWLNlrLLY
oMbVOxDE1b2je3KVSq2Qzjprgb5o54aJK3ptp/wuouQP3ces1gbmPqnW+0LPP7zU
gVplxRPD/vSSos8TNKY4IoTTNAF35FeHpxyL4fbcM/pFbrnysHtRceJ8gX9a6fD5
9qj9x3jLIsSCUdz5X33IeIlXkkf8Tdo0NZkKjYpzWYDAAv5lMPaj0FGDjqhwSNgl
LhI9uuUyPDoz6U/ynTLH6KQXOo/gPP54Ddc0CQErcfjqfC+JMkDjhe+rHF31b4io
gFJyMRUpJCuGO15pTnzwm4dW3l+2owDjxRT/E6mFDuv/QkqwDQtz6HFJgULejMYl
Pv71fANeNPTsgWcIe8cJsRYy6Sc8G4T+SNjb6GnmdvD7K3QHjy4ZVNHtdKGXUZDS
ahjkMHebz6NqwcoZoim1j+h/zHbtX27uurDRZdO2bKgxsnCDhoB6GhwRUrOq/E8k
WeC7pziLDjfDCfjkM9jLwNiqVSdGQmfUn2ZKeEFX/d2WCPT6go8Nh/3eyoPt5pKz
d657vcExjspCJ89jzg7jGSjSkO2tnGcCFnNgpR2YPwKOHk/t7ZMnqRrF++GZLe+x
l0vNatFEJ1r2mjIWbxdUzFbZgImSFNvuJiBhpq2Hw6aoZLIl+r3webOIfwTyH1CP
EdBWihTNj1j0iiK+vkHhKPBPJJrrg0xBISOzI5Vh+SQH4SfYFbqQ5+78dvZD3F7h
wJQi7R0Mq8nhpACtaTtobmvDUeFqMhXDOP5wjWNBJzFdRQ15hGHAoP76YPTNqGlc
cznqFF1iYFEIbE4EaQUtSTKuWwIjhQHx77SuhRgK6fh002eh7FN+5MoZu/fleEFc
NcscBF9TzI/YsClcMesCGWck9xO/uOOnG1E7FSARZ1EGfYgm5SPBYF6pNQP7wToU
crSK8wPsAADkz9wOwb0TeVAco8dzBl/WIMlnMog1OxpTXH8WETWyCCkm4G0iL2dR
QWUbaPyISnyyK6wYlfU3Aj0ApjrMskps/o85QliuAB9W3lqbnghBb02zBDRuu+Tu
+vodLjPwQYaLGThyX2Qzvi8qfiyRqcobtAJU4xRjZWbKdkyLWx/rWtluC3psbPHZ
o8VWEsm8hKFhzZ4DBsTbdpq2+LRBk++slIRlEBmn5b/bB0W0WA6/kG1geFXTlHQl
g+eIRYPpavOKUvuXtl31wcxr55eTZomJV0SiZpmBQ4eDPS86JyaJBYon4oQ2svBu
0wYtIgL5ToLVag8q7dmNBSy6bOPZJdYEp1+PRVJ+bBcgy/JHPoiVB6hbUat2mzTB
XlTMjbcd374Z7hvpgu054fNFvfJk6ZVCyM9cYa1KwxggPmMrGLzOHWzj4U3QkN4/
Wez9UhTjswu6yt0MWzfTSNFummENm2oSgzueCV58Dfku1//QE8Qs3QpzdNohPi2U
XAnXhbmrtpr63crhAlIPYf9aOEXZ3OfXoxi46KhC42pA6/X1MXo5SbnUjUuOxBSd
Y4v7LyehoV8TiNRSy1Q0fvuSonYF5BafNfPErvAdTRgjGvbbnBwU1ADqZrmXk5T9
1SbN/snO0ndXe2dXTUjZ0Mny29xvnNnTxJWgO8gaMPETO9jNojURTnH7GWvF/cxr
A85394MhOZMnrFo2gCo5x/IvgiqIDZ4tsXg2C0Oc02EMCCFHfe1Va7okchgcaikL
SDJru6AgF7xx7DtOXF3rSRk9zr8OrEyC5nDe/vzIjZi91TtgOh/Bm1BUo+gtB113
nLBJDg2fDnNPVniippre7Vy2LumD0Y0GTOAIe1HalyEuYSYWEQMT30CyfUWiUyoF
cWzReB1w7y+6p8ZV2NdvBkoN48aLnPnrMuYH4vwLlxYIXEt29u+rCBnRZm9D2mEn
a3WTmrUkUkUCjg29SzTwpR7BChO/ZGCIxYkRyK2wZnRfWxjaAYaumf5a1JgepOPI
bsQIWK7Qf7bxf2/DjUhoe1tUHuqIUXL9I9jMNqOtG90t7JPC7WJWc3MWCbgrGoog
lOnPn3xOD1r5UI139iwb/D5D6o3LryQqXPTLEc1a48kRmfV+Propi/KHLBGn39j8
brn3QcqpW8lQhxYby+ki4QAnZTWTBy2NkWe74EF1VyZfP8C0o2jBSkif5xE/RhL/
ACOyUDYJdiD4dhW0rygOVRmsc4y1h/8D63MlhcvcICHwOSLVibL3g2be0/qdTpBs
JfgV10ql54QJsn6ynmsbak2IXiJqsoPFwEfY4DWjtm+euD8dcQa57TyRQbFVVqi6
ciVr6gVPrgDMY23zOrWIZsiWClgcwN8M194L6ZTXsvEp2QXCLENtz3RTcp1g+s8j
/7FNyvFBwiEca56ROmIDpNC4Kf91IJ9eZr8uE5OxMkVaAbAosjkoVp7mOqAMrpOL
236jMILBZFTegudCRrIrpLSCFT3s+OHilB6505uRPsqtGhCV9Dqz+Yj2t+aXJe7/
1ky3rGmj7VxRF0U+uko37zgkcU161VjD+9j/3JcRqajsfAKVTYzpwV1yZ3piDzqJ
VOJogrXp2NO8SS30H5Y4oFaLuR9QieiznuBA73eQBWlaYJHGDUpnBcGM4yK0tZ9s
SXpgMFfnQ0gT814X9ojqAZ3T3uTOCJxuHiVTIc2mpUhJ3CwCwRyiggeGfJv0eYWc
KW8jl17GlC5nWmzo4ySqHhIESUhCAsBHMZhWygCLfGXifX7Xw4AYzjiY+vXrlu8Y
ilL4GTt1aDrPiMlMmsEqAaN770qkVfVwElJZ7OYSMrmy1o6pux5R2vFeUypc05AX
TT/YFZVNVT57YQieRaJp7Mc9sPELi+uOIvot5CpEOm6uDc09B1nX9ohDA+GQfCtj
vcFW7BRJAltzp07RPX3ciVDcdBckT2OJlBAViRq45bjG1eTgDRrYAOlvhchZW5vw
H0avbRy2pVpdsTAwBa16dWZ5wi4yKdvx3BcXM9CyklEYVz9stArl1HWT282S906W
lfbv4ohPzvcfQ3GyZVDjLYP++yEhRrvmpA6XrWIWHZ+osL0LRXw8jYoAd5djgkDg
Jn8GOH3jZxUeOqIspqkStsd9FETE0xYB1nTzj9xk99kMWlxAeqE6KVzzwxKqHx+B
AKHPBxg7wfBJg/ntLyYbUJuvxRxwbvLsUkL223YCNSlp7iBpxmoYYNiy5DRuo+sl
nDLCze3lPKgE9lptc7SW9EegEuzbyWsjpP21jmrunqITuNdLeXLWTjLVreIaXQly
OLoca/81xhqucaDPZK5Z2I5SHOWSyhYFlWVgedmRheIAllMFhQ3jjHkWsDjw0EDV
uRSOScQrQ8JGkQcNvNfDSoK1zCK8lah+vZ8wjJzMUSb+vnuxyU82zdhpL3A1yHsh
D2GAps0FXwchVjH6Iq32nHhnjDeDOlnJafOGyX+jCg3QDnnQq2IDYfBhYb3mEs0d
lloz8t2pKui6F+AIf4IUND7drFxsjwdTUMTeznaVmjjHv6dD+RW7UP+73ZHcsZDL
JDIkEouay6aC+sPkaOpI4hmK/oRXon44yfxFpwASJ4KmjmHPAqMzAPfwpLmIrN9N
RgEWSZYO9pY32+YRiZUgHN/3qNnz/3gcO5huThVn5YY4HwhQJ5A/EBBjoW2a2rtb
aHRngNAdcoXQEs10tyAgGK9rY3H6dj73MWdvsQJ7txmIGHn5PKd6FETfG2dRj8nF
kIdjrBZI8d1R7WYImjO/zx3f8mNhAuwFIzzq/OoVTg8va9NCIWn1hNTmajECmpj9
a/ZIgb3GjceGoq9tA5Ig3ihGRxXaZzbRgh3NXb6bsND5Aa+idDTzW1+FgQTQ38tH
OtStthE6TdUKZRXoCUH5qHHPv5bO+0YutCCKPlRUxp0K6Lu2BtjzB4SG/fDig/js
W72P75miq9S9Gv2wX8T4b2ApRmgSLp05SPSQDVT+vSk70Q+T2n/10XiEKNiTPg8W
2PwbdLfp8wfUa9HVn+e/2NinF3sEvpVZURG6iLt53iAPI2fms0xuDeT4daMtd2RW
8OD5nRwjeFdCCnLdZEeq3v8Gcp5z7+hwrjtub60In4mUZppAr+J9JrLWpXUb975y
n/TTSOr7/eZfbsbk7J00P/k1Q9LxBW8hZSBwHy7IcjlsxXr+UWalLzsagMLJFzRi
7IGI5Fc3mIKjsHtiQlpWOFnDF/b/RH1K48LtornAgwpVI/cGDQbfpzYsrFC2SOc5
R7LBhR6th5gThrEWgNaIFu57evjfZH/hMY8JEay7R/zMctc7gUHN9RxwHRZkFChF
DnlR3XX+RsMjTohiZ5+bxFOoP+/aRdvG40oySQvbltso/DJ+g6IFu21k5OE9XvrH
mrnxYpp2fGVR1+kuEj/3qzD1FOiCG+b3DqENpIUtJBcN3o8b5qgObZWPv0ghRaAi
V1cGIaItgm8QR9DyPdNpkn8T3cr4f5+RmZFfoEJAW7P7DOvvSBe9AJmXGpvUVCUJ
8+5zquZAwFbjvqAa1BnMHKfh6Gkoxj0xHVB3zZ6a2n7XaD7WChKzRLLQxOSg9mNo
0hb2GFPhP9smWjfxLdhLnn353h14UCxTc7dKl8iQKyImb2vhDkBv+OkbXVsJi3gQ
E3PygI3ctqbFMSnNBTBqlJacbwMxRsphBSwMSPokIYtAPziWXOKdZJuqhGqdmwJC
98l4kDeqAFAsLI+LQzwIkO8O/KjN9E4ZiJkumMQ5LmfcXTv2II76/tRTotgaW1H1
HQt2MmHQoFmwli4+JUHFmT7842Ke/yFo03YgtMSZHzld1vnWZj8VAwoyjHDov7pj
ZmhVzVSgRcJmZt7XbapLpst4Yp05pbA8y9VjzjmkM5JduVZ8RDn7IimnVczLe4V9
caZY1vOwQomiNleFKa6cW/6FaPFs/JlPy2RvsGz5+YkEMP1cWOS5O6Y9O7G3+Xif
ltvNRLZBvPkgrYtAbzM1V7mlrTSinKtucGbjgaPqJ8a1VV+fjc9LO5KQiwE9rGO/
uJWsHFk2Audn9+Yb2/FDoHtIafRyyV4N4hvK1YUpJVCMZ8RXEsBejRhOx9hOj26o
skOUIyjrJunVE6zR5BtypHaHRkRPrWMBJOnKq+KEO5HNFHK93g+mtJQw6dDsdSGQ
SDsPbEhPPFRGx7t9iaTlmf2T0BguALFV/hUf3Hfl+RGWq2N+DHyX3xypKTA6cMkF
syDI16ABDpoNTxNiOlECS8y7t2cK0hNZn7NX+kSwp3SVYBF5cy6ZutX/8w8tU3T1
GhYsidmwIUcqUIc6RwInamwX3ftyRfyDiaKqIIU8pen5YJjHQnzkM0udMkst4R2H
pFy2WYrAmkgLWrJwhoE05OYfg47XlaknmUPYlacOT2x4vnbuoOgy5Hx36PG937qc
hyn+XPrrlAfyj7dQ2tuqThi2M/RcK5yOf0UvsIH2Hm0ZI2y4TKQw4Wm7Y7yMIM45
qoz+35vPFEuB9U3yoLO0rC6LFgbvokAa4lgftLh5n/QPvdynATp4nLWbX/jbKoTw
1G47QQ/VVG1WBBSjziDBExt486+Pwa3i6SAgr/q3rpBugAoTJxzdNfmjr6hn5sPC
Y6oETOw5h/bR23tzAurFlVilkOF3taHfpIToUDSEZiGxQ+4abpSpoZ+H9/6b0Fbd
QdmepxrjheVyeLMO2jSHpMPynYNzuYrvuCklFFa0+J0QPJ2/Vo/QGQkLol0EkQi0
c8QYBMwLxv3dczCPn6Ec57hA8DAgngCm60tgcJDuDECiwWskpgotkjgd7nfjRiS5
DuS4oICuhzRfYBLYtosVpyGlJ/UJuM15RVcIl4Pk+22ZGB9fJr1cLamDgvK1H9Tt
OC0JPYG8kFU66ZOapjDuQBC401kyMJXTCsiy2c3AS0tEzcSDCenDj6FNKQNi2g62
q1GwbmNu7ee+QlIz1TJHHii5fRZZxGkWBMC/Rc/A+BONhS4tAbIqDo1WW+/YsZiE
aDKc5eAZxrEX6ewOyM/hwoC+oWXetAM+g+BNw5T+xGBzgOOymiVUY4jotoiw0bsq
RkFUipah9pBMIOfP2rUm3Iy2s6MzJiQaDNQWI71GG9njrNVs+th0VWFm3za0eG77
xMrwR6kh2nj1uL4O5xNgNy0LbbDP0op52qURPyOBzk+0ViR8mpEa1Up1PhzyxL9l
TtbElEhuQJad3j1d+A7YTRFMNA7HFyGo5ggKcYFrF4NSQTNqYrlT9Jol+CwfMxa5
pvzAxRt2zUSN9XTnOrcJdj62ahskpsAfL/PlXjCcfwrrcxJuevbJ+GAOQUCQ3Lm8
ciguTRPqhzvkiNxSepcqzlGDxikMx8Ka0HN/054b5T9J/hRwJiIq+pzAlEZQISEh
o5hCNuZsaZ6HS6ZoGHKoD+LVG1lGP71oaBZDyA47lWV4zKp+ekr229/xC1SFEPfR
fr4qi9aWhEV26yZPnaarsvY5ziUVqPJ4J7AIOAQwyWXYROzkLTp0EpXFee8Gxqhm
tOsgt2sIrgXlVxSlDnXXYI0MHyI+ddr5bPicBgPMlEzQw5F3NJtkUBrP+BdrkkUe
QkUa7vRlrN93ArQImBzZxGZoqPYIdyeY14IrjNo1i4zeSOvrM/Y92SJWswg58hBF
XjaCaqEqD2nicf1TwhXzzDMh90ivw/IpBfMNlDr2Kg9Z7HqBg1JNFyWaD7Taa7GF
0lai0pjIXiu9m8V5em+9G7ZlcoLR5TQRkzUY9s9imib7VHWr1flvLjw1i0Lkplhp
vkluwvqb0orj9UdBwaKRpqsyodmnWwdPDvOne63FNSuehkjLroIDfJj/HbP3V+eE
jhoeRG3kZNTXHwR4ZXeFvjxprVoPuYihdV3iTdjgCwoorltgqIWdAUK35jOTTVVH
Sez8bdiG3Ua0BmyoTjvdxb3XvCiyKYtpbNn9cuES7O5M68BHHIhxvwd/qZEHMV2b
UBT3OUTChgowDjBBC5NuxIzAYyQJzZjwmn14/rs59tFYukHeXxDCYSug+KberoaU
Or9O2FGlnnsPIKYbhEghML9juZda1wI2CEjTnDOSaStpB8m9fQMhNTcO+JdwZjb7
OwTM1OQoT3cHTtZl4qAtUoatryapOXMtIsE/Wo1XpdhSOy0EiONKSwxHi3p3Vekd
Pn6L8VuYdsyJsketL1XyE32hFSDHX0w1IU1sI4EowXZc6U87p8DKbKzCBlx2HgP/
smHDm10yAbfuzlMm+oKRp/i2VZkYhAxq15rfoN/Q7aydrH42Z5E/pj8IVSDfSBxP
PIHwaGYrhsnr7JTCRfnBvHHgAo9ukcT6wGRhi2AJZ3dR3Ms4UOkiG62wg1+pKnX7
g/sn7xj6asZ45Hb81lNdKKQP2/7jc5ZxkfEnuv9C4oMVK7LYogVgb+bbOQ5wILXy
pz593iYz+A9Ykz2uhEVOm8AtJiTXnLt3XS2B4rsWF5N3ww0eb7BFMSECh1hsrOJX
9HunR1pQj4FJkTIvXz/A3AdKcZZqEZB6bgJNK4W5fMbcCUsEtd5naHJsoGWBFbeU
RXioShSvbfXIqEC5I4+oPsNLJXwJUvMhLoaIrRCVMrA6EZkXt8BM0oyrstet2Aw9
4mXuZaR/PhWQSK2j+JeYjRR31LGbZK7Tj5DTs5oh4ONMZ1dZ3oyWXzOAXQCINiJ5
rX5+PmtkffHYUHXPZfBEWfA0C/+RHGRcHpZyBBiiAq51ilyezsQk5lmJeZAzPcu4
FMcDRh47L+hvgTrRPUh/sXN+yiZ/I/QyiqmWPAU5DPOMRUR1jcgZlqs3BEgsXtYj
zP5slKf7Y7FNsc+MHUuIozW9sBwwJWTCN7WD5qrCPi3y7+3oJHlK3zl/dIzhuJRU
GhwwG1mLT3ruLNNViAbhT9szNPvc7V355SKmxYZA3jQRFbStWvfXB05ydgZacCJB
WcbGDMTTOlBj0zEuNgg/vxOfZVD9dhZ7s2J4h6lq90HboeWK+h7EMieaZXhW6fc7
FjNnlp9qzJCWZvL1fskZ0Vj8l1LkIylv8mtuJLSLQ3HZmUKi8eJHkTVQ1S07/5qu
3ZhqlOydrEUsQJ6EA9TTqxopFrxxqkb5rdWf8rOkJNh+b6z26v67ojwTuBFeiMO7
ussPU8JqiQAb2afrLi6Op8jilvC2U2frbZ7VwtBNSpVHq2sJBlwn3ZfC3+9AP1CC
jsfX27gGaDz3Mc16PcKVTcnz3rQJeLRWZNAdghXzDjNW8Jbz52prXZv3K50AcL4N
advO9gWprAtJDt47uAMTXb2ZMJEqwA/XduG4y0TvJ8apy4DuuQ5qaQD3CyKfqfBd
j2OMpH6D/DjxD+y45InOOiEplHFvCziB/jrwbAXPwylUIJ7F+0bkaNn+RbLqXDLg
Xi596CJiaeLa8REpdP6WzoFFiH0BpyNNzJ6Ded0N0JKNnMa7H3qAXQ8d/WYhVn78
19wTR57Qohag98F70Ly7WtbRbsigDfdItIzJS+lgngFs8q3Um3AYDenONKXmgwLG
1SEDzR1rQxKfeUkj4sdKxsfkJ3PI3ZQjmROB+vidNktz6EpEQCdxgmlZxfzUd7HE
JNOLbcD6eB9jaYYn9f1qnqsfHuX+y1w+O6fOyH8nhM5hDzSFN70tDZgai6rIMofs
vyo33G1IwhpgVPlgubWWMQ2NRa0YZuewR14L+NdC3slGBNTcBMlQOdaOI0gG8hT9
Sbpum7zNXkUZFUaAJO1EoyZViqsaQo9Z9xBsvQ2nCpgTPC1jYitLgptUjbNgLvNN
cLTDLamRi5fT1O8YEcqxaBZuBsjR+J0Ld5FeVk+DHrURtEaqVDSjEyV/7DglCzTQ
E5NObAIXydnAH/+UV368UQ5HPM2KFqVWQwiATzF2+mG5SqDK3vq+LlqSMxVV6I/+
wv0ck0QOqRNeT2KN+JsTZroTWfufkdqnM8aZJ8goQml5ZpbzGxddH63J6cTzSfN+
+qRdGL2kPrv6sTwMttoxW6kQr/t4zYgUjTWlHBKeDL76QHVcHwrMsG4bhCN3V/GV
h7oZg6s3pjUrKTOQ75lh4HEkWYr/mHN3c2Mom2F6SEy6foVJZhuu3s+3eIQ3xtab
AQzQHZMthIw9It/sYiRfFxLBLq0CyACtHrVvYkh1Cb3RCmpvToh8Dxj+Jw2KllEl
Ih+hvOpkymetLEDVgwVJ1+Z/EWxDW7qEFTgfoBBhXt9Gm9E6y/4joCElBfLr8/6T
BKpe69iu2W0B5iIRgrctldN9lnSimXl6SxRFt/3RqSceB+bu1I8gT5Cuso3h5L+S
kL1gpDe5e5FR/kuMDBGCn7nmuO50BQstIPpDjB7xrcvCHttlYWcRbeE/zJIpakZP
fu5FnwBPegRnWi89wy6OalSZtdhecXtL/YrqW+3zewLkRWjE402SCNUR6Jl/V28j
1+1r1FGukkTkrq9SLj5h2BLN1a3Yj9xlMU60AyDNFYwmQJcqOzw8yJ8vkNrcQGSU
oTMGvTI1IbjNkFESspQkalB02iE6MUC1My27OfN4KWuYEfjJa86U9GpCg9vvAk+G
v3DpIWcm4jyOVlKVRzBke/5xfD+FFi4kpk2+msz68rFtuXG/9dGsmhg8uDX2PdmT
kl18AEiRWMcI/2/vRhxEYGcLeShToazc5ObG/EpIMWqHYssC4zLMyYaI5ds0HW+3
K5Vzvc+bLaqSasm5bC1z1BvkmjyH7XLQZi9EnEx3pJYXeEVxXUhYH9GW5LTbg/Yy
yUdKL+krSsd/0RSxEhYnOczrBw1yImcOlMZLlZpPqVlqG/qXxiEmxFOQUMW987Nj
VET6sWPao+qirysIZH0Bu4+5LAv+n/xREBmgjFo28mXhvIf0eR8mYPvDQrTq4DLW
QhLImw1+g/QIM/aeCzgnDWbshaFX/wr7WhLuVxhp17exx2TIr05hfYVoY9X0UApV
mstIhUi9I1Qf8H/ERKCwvJIFhB2vCzHEQHRjABvvS0LG+PoJA0RQ7mhEWQU050L7
KqodEilZmNTWgG/cwpF9O7QWVG0wGhLVb3yJ3TUmf6s5CVD3TUEDq2ZY7HqC8R7O
Xg7EJ7WVoWWWxMMCvjOnkmGAK6rnozybOpiI9hxRBbbsk7LYiplYKETY5vLoY/tp
Q1lW0uAKkHzCle2Z6jT0t7wr/Ep7OH06rYnjeb8LHdEK+RG2k2DmP9TfCSHK3sXa
Jm//pGfEA4wtnTsLp5n0FjgYSyK0w33AW0FCA5P43OYrxZV1BKJ+CGNupIWvKwFY
pAzzGOYNT4qV+kCbQsxNvLzt1TTZzoh/oBIN2hcSpPkXHKboJRhfQXvU1GRA6aKB
kTSybPPAMuVlpVPj8yFEqeljkHvoU20Xi/aRmoVMOcafnd+fK0RkpT/5AUWQQ8I5
BCoxnfTP0g0HA5NM/MA27/J57A6Kn5nXy0B2+YyoPIK63CkFpHs117bOdxh1+s+2
VwJ6NcAcsYFvFwKPnSNLJouPo9tYIdD07kdm5dwhYcn0JYEI3Q1/8U1ZcBoH+p59
f/B3ssUhsUk00cnpqiX3XQvI7+fnh9oaI8YN0FxxjPXMQ5UWGlq681bobZFnRMel
uWL3Pg2Lk7tAbbyW8g5fXaOZ9t9Cua9vcVb0YEF7Q6VcJLgKU8LzVbB5YBHnWdfp
Mdoqrt4KMFfuWynrsCdBc3hz5dZbMqxMmGpK/YYu06lTFSXMGMQ6Jj3plU08HwQA
HkzhV0mNw3BqcSnObZkE5bFb1g+jhK9C/ykKJ/sgLpqdWvhb1E90KrN0VMJUCmdl
PSJJ3Ml+F97gPE7y4l2Eq3XXX9b6CZjtabsyWZ8JGZyS3CcZxZlcJc+kEVRYS+rS
7mNxwTSi/Hbv01wsGvoVFGaIBaEJSpoCfMQVqBvNcMZ5/jK4mSaijg7zknaTYvbN
q9YVHL42JCgqN7XMpgILPxT5kN+uuO78eIE44lgD0D/sVX+RhCot6VNRhnBme08e
Wywqsi7+nHvXHnFqlxkX6ViWk8d0QRZorceeYaTzE2kFM2TqaDxqMgIE4h5/PbKH
x7Pnspdc9OE2ISJlUY1AFPSWiI4FHX/MQINCY1+fwqRGTaIeY1BN1hVAEeavPQgB
zFypAKfwe1ZR4i8cKfqkzky37+PH/3emVFW9h68/4of1XqfXO22DQYWcWJZ1TxhG
YTcqErhN9rsR07aWk7k2qBFgFCiSv/Uu4v4GZRxlqKJu1+y2OezX+LQAoeUowLMH
DIY36mADWjnK5/n6uvcZ8RmUxkpdFdFRIY+FGjBA+tDHvTbZ9fF5NgzUoMCrX4Q8
kzHTW6lLCh7Lf7Z6VZdEbRU1Xcbd49Dxxj3w0DdCaasrJvfLnkTR93GzQ40Ktk1F
UwPldwQGhR73oZQezK4d3wXxE+TVqkFK88ABPvbZzzSTdQ0mh+r6dnvSVdC1txb7
8yKZ1/955xmth5KlvK+QfApeZfw1ixvBxIf5B1u2d1T9i5rhA/D98RJq9OehIMpr
l3ux9rCGJKVfvipd5d+EO9W8/ltXCFBC43uaJJvDpIZpspmwkGY5K/KsNyaa3eBp
p5p2QZumyND03Xen2jl4j+7/3+ZAOiyNKpvL5WPLhV2o0QJKVrd4gB0vArHs0WH1
Xv6siDVRKTia2X5/x9Gsxa4n9wZ07aBpBgU3xdP0oQrzvr+YZc7TG5S9xkxWbXz+
sL8JMay25U2tfre5s/s/mniArdsrTHKd9p9FLoJ7AafJtZP/75biTiiK9SDhp2f6
mHJ1j8L+apSx0dYhqcOoCkXss8AK3Fr35Z60rvmx2SK0rutKhi+P/MKIqxSnS1Yj
pfcnDG0LitfKx4WdiDCO+MNlrDfmcI4lLdq8I1WuE4QmGQi6rSfyTdz79l1Q48Ff
JDLO5+N/Dae5uO0yubjcQ2zKF6/i1p5U7OE+QCHuDqT4Y5hy+RALSy33rjpJGIKc
Ou1I63CF3OEdcMJyl4WBeugiyS24pVdWH5VkwmP1ro0qkknymh7izZaK/ZYVbvZz
+BuE677KKwwKqOGTZGeBVGYwmwDwsFEPPmHESVR6wcoQsCp7WbJVVkKZOOZ3AG6m
uYz/lIXi/pkh3StVzC1ri4HseYGPo9yEXHGXoP8GVqyCTby5gQW4/9PUrp/XLTek
G+RAD+oO389u4Ko4dob1AihETUwT5rNhUtpVCHp5kNtj2uRHfi0gXMYJq98gcC5S
fFPhBE1o8Mvciqrg9XLVTNMhueWRFxWK1n607h/qyMb7yRQR2aIrk8BsnzR3Iv//
kfW4JcCL/nVB11zuGDFoG7EX3fq3JJPjkTWzNxvvCiJ7fVIK0Y5kXCFJlAqym11c
7+Y4vih4Rvw4M1wMlDebnKofNioFi9Ynfv7ktmfLtQIuf8zKOXoYIuMZXqiP9EHM
SpYnGutrz6k+7pjSNIwDTCmG57xly7iay0q+MRUXNLCeArd0S87stu2PkFL/psPm
EQ96L7QmS9q7jaYHn0g0SjKg0mqnc0Nvdqyf0b1O2D0qjDIi9gmdzRkGMFKtFR/Y
ywIN8X6XrMGBzcDC4O/RSnaOUdce9GV7KCTjLq5RGQERaB9nzZACtL1+pNmE+1rl
lq6Wetryq+jVAzSndjoCF/tURVcaKBbLyqd/VkzvFpk1FkCB0DwwKXT7eX4Ad69N
I9KhQP75TUteWuzvuKa+WNZb67XCJr2I/3GRO0RHIMdEsrxpqRTd9Qzh7S92LfKT
+aU+EuAA6YfV7e5x51ua7z578HLlHPUYN/l96wqW18DC059JMjPGHg+T6RPTWk9r
+6xrfnlZNpjOMu2/q6R/8zdbp9VetxnNmY/mOKuq0KCTqh4aks3Cxk+WrUpllVYE
cmmbOxhjrKGma0MNldofWznCZFhCKYMDfzaShvElm7bG0KTTG3g4lpiLgr1rJxwR
TVdOoa5+nWm1mfFHa9VV7PVmzn/H4Lh+giElgsXZJfcnMxRWKACAXjNNlfgl8vXr
DwU8cXM1V/vo/ROnlPei8Nxi+dTYXGiGPP+ZEL+Be3SV7P/vvdROnvp3LzgGAbq8
6Ma+rMFx8LcKdaGAijkSdGXs1gXM7N407LV9BvN4y/wrFp3dgsnLGyijypZfOONG
t94SxFazr6Fdij6u6278nKAEzcdzW0fdSt4k0fmYxDVLRZFozHhH/Kc460769St5
tuhBh74xGU6x+fGB5MKiHv8xXpo590Tw8U3cuf/qUn/GpMmZ99soZSvx26VSmYCq
gosM7K3SvL6CmihTUA76KdJNg9FLkN/Ui0svGm2webyZlHb75tLwKCSmZR0maM4+
HLipMBFMqPARp9hLk+VMz6q0v2sGoMxF8uK+RJtyKPQEaq56KtoD9Op6+Q94TZCP
6AnUHAfhLkou1NX1VTTD4VJtQYh92BVRoADBs3E0jkKl3uRpiSq3u4bXDgq1OgoW
w+FTzNWPTPQoQxXV+8wTipawBga6NOuJVzTWbnHW0FEjEij1KYg9+DdxlqTaRwg+
sncJh6g/FdGKst+pmNACWyiHTA2MJV+4CCpJ96xVyAzi83JECLeWu0XxyXfQH9Af
W8Bqr0nGNKdhmxRXHmsp8p2Gpp5hXJlEydL928cLDElUxE+YpS/St/p0T/UjZyw+
RPOHorbJ5QaFv6+fG8NAChLCJRDL83jQqWj3yWNFJ5I3h1huq2WJun/pysg+FOQe
KRkWNmg6CvMBmA8XmANvy8P3nEWgdXOXN+0mvUB59JdSGPl7yjYWupOF9fxo3PRD
R8rrzNgmOU7QlIfgLwJsLm1Is6nPcnEwIQ+mdvjpiAWM74otyhehg6LvsW/n6S2/
hAIBNQOmHetDneIBVp8cpg5ls3zHNCWluPngqJ/PXQktuYw4sE3qCXg8ii2DSS+D
yCzWJ0V9OSXqjAG9zPbXgLbjsA97AKwwTFM7G0JcMBWxfSiDsv8/wm5/AlwUFlgB
LUs5LPZmz70nUdq5DQdMAtoEKsW9FMyHAjrxWibiQRWzrrIBQecU1tax+ltc/5cs
hIoAt83t2qKGq89uBSultnjq7+S1RrhAX7/udRKTCQlVE14D4ADb8wo15pgOA2C2
JkHlrwGq0EUrfrPEkh5L8ramRKNNKbw/pJxzKh5x5GPkFrtkoFkytWfegAHhclhn
cmoBZGxb8TbbUbuIR/ZcahddFOBH5imvDUGuHu46BzCNNjdbP6tZ9hQgBKGwM3yR
quS1mFJotx1gT8sv70C87BGO4IbqTHeOf0Hgf0h0KiLpzU3Yv1KYMMzljuxgFkx5
U2cV/OS+0m78JUMukH6ZORnigPozLm0p859W/yfCBEFUTERdG0Quu11lTglnXVYy
6vq8BuT4FZdhpz2kBpgeXDd1Tydcy/0wv3IiaK98R/xwN6Gzr7GKe48mWSYQwjxS
ae5yeIMd3DJFvjqu6gGfaXLpg1se4Kos3V5sIqcvAG6iw5xbazhAuVmPF9aockUY
RvUiliQTy3iXOq7FSwv4Egy+0Cey/rgQiJou7VOq8v2C8VUAiBLfc77+WEL0kyCs
z33ZvFs4AIFcrGgeeeHn9d4CxEQZ1geJ07LAwL9HvmB53S2wl27yie1vPLU+WvbV
bfpGPF1iza6tMcGJGgTuFyr9PTZmIjZH8wYKlucQcnf1P9jQ0NZN5n0+tGIWFmE/
L33+X+2RPUsRFK1y9pI1fCxND4si7JhldlTxjkkgP67OPZYFuCNmy9svntPazBvI
Ss+2khokTT8151/BraHXHxHEYWupGfrS+lw60n4ASfXpQgnirz1lbHcYva5Swuoz
VrN9D/NZgg62jJorNu+H00RwJyP+SYcI/5pISSeYUx7wYEMtloYaijPlcRtPprQe
iTfneirENgHO0ji/7ifVEmUh+MjzohNW4MrngCBvOsMwxNj5zD9cjFj8C/jrMDNz
Got8+GnGM0uwfuOwMpWFDMSjrdaovxRFXeLZKZyxcPTl3XaGhsvHxllXY/i2QlCJ
B7LupRfxwv+oWUsMCAGD5OJHtLRucmTg6c6VnPCEdQ0UCnaNtF/kFv+hkfJA25eR
s4mV5BSkik7j7ZXCova2DSHof7D+bzt6FO48ofiWBm3DafkEo4pK8F3xEYNoZSma
t5Dmqji80IYeMuN56GBews/S0FBcGKQnvHj3u8fkUeJNtp8fJcjmzEyB5+rNY0Eb
xqyMxY1Bj4/hlwKj++otobj/H0rNmpUGG/ds78vFCYhoICQsCnl8Re0PdeIyOVAy
mspR4Rz2qVmxl4nsiFY7I8r5y95v3whWDtcYs2rIoMBDswJDOwXci9Lsc0XNYPCu
s+OKOods2C2Sad5aj1PQllqmtmhv93RBt6RumLsx6eRYVU5/9h42qqZ++l3ttp2j
qSIVYU0sCFoYdbI4Y+uG+riWY9Gx6lhs2MYG4Hk9Pg3ihnaInTqzB6FXLLUt8WTc
cveh3r5WOnFsD112bSjnEYYvGkOqBE1rWKloRyn7+zJKaRTcbvC49IFl79/teYLr
Rg3zl+6CX9lQOpoykoTceRDPtaIO58GpIQfx53+GJBPTz+rjSiB/wOWkT8oGOuIq
cQz+I0mFHrVV23uqSndsqsYrHR6+WJ0/8ISe/jNgPddmN5nZkLpXBAQxWBqnU5tv
lSfyBzhg9Ozk2K/b6Pz3zx/w4WtC1+Mp5SvoZSs6Z5nOEXQTCOFvQGX1t5AaoyEK
nWTtox0MwwzqqKR1g0cO4g0LTggMtW+yWR+i762wKStB40rLNLAAie1o9MZeUwur
cQz3euzmuwd8z7cebR6tk1LiSfcQ2G5qJnb4wzXcfJoeXRf9QPvq/9ROjQYIcIsW
fv4lyW0VwWQYoMYoe8fme2TeNWW+hBROe1m8ALTRm4xznGZmMud/FiK8X5AqzMTs
iLMbmAZ9YYnj75j8Vt50bqqRbk3aRaWM/u70AEjpZn7O8CgvPLlz8WZuJCpLwfWr
5pA3dS++KkkgrKm+ZKxUJZN1x9OdQEq3yoHXDeD5QJVLcvIJ98NPgo0p209g5uww
mhU0zNKXbA8BePoikmsK2Ft7y/s8zArwYymgjbz2vYSuY1+wjO2zvg72MY4ybzjN
LaEeK6+s/aO3OhPqjvk0KYLWEVijGq6WKC+xWe/mQigsindOfAEVfXdUy8Yfvebz
wHRzLTgObVaMk6xxQL2+4MbGX9+JC2Ru49hzhsONGewtFqjplqRYpEr74lMwBVEb
J0KynJqkJKkrD063nJ3GceRBeylJdxNNoPHuAUv9BoZpQhcBlIi657FiFWX1USOM
UOssG7Oq0/B1rA+4CojVSrL9nMggXyvoYUQQwqqIUXDEWR/qllrJiOauiwjJkMwM
zUIHHmX7L93h7x/HoDnlEdrLdSc1kNfH8rJ4k8qJsFrmuykkSBzJjTs/iuBOA0kK
nKrVUlMX7MXWW3Z1L4oBFtu8Whq/Dai6yE7Nm1ZVlHlcnUE4xBffqyc9u3eruYe6
26mCHjWDrQXTAvMeY6KYq30Bh+f1eyKd4Y+ZkfThTUDDyFL6FMCJWWGkmgPpE6HE
QJpKxG/51efTURg6IqgPJDdnNq8nk4FvYRNe9IuJc/gzmicTbjOEaVmG5UAF8+be
tHylo1SrPzMxYaZcgqP+oHKFmsupbcyB8CS15/jblW3Z6SZhPubQNi6jJGJE48wv
CT0OsM3P76/MVL05aAJyuKcqD80FzjTfCuZixVbkg5izUly4FhXVqEobtOWpmnr0
CYEia1JQhzyExHF9bZtjT5Q9MWvlrxXCS19iV6n6T6ykooPCSaRTzeKe4AKWzGBy
voFAE1/Rtid5bGL/Q62mJVqvmN7acaxnrQ3l9ZfrE+oY+qHHf+eqcOw2UYRPt44r
T97RdWWQJuxRk4LMDp69C6vSGo9FS48MzoRykZNRHKIxil86vr5Ns6lphG73q6hD
Y5K2fqQ9d1hmgC91Xaly6a2BMxjwQIRfhtdqa7m5Dc4mqvNYCeb+/8AQPP4TiWhC
prj+mzAwneLx4k3sE+r2T/tlOlvlJmLaNOSP+jwpVpQ0w0y8/nRhrsZVsC2whQsx
x3oYOapUPXD2UnGBjFPL/fCgzeTBnGkIQ9Bc5AgL+cA26NZ/EmyZMcZbeSTvz/kT
d4GF2ajS94CIceQlyVfuj9qli0sg18cblde5EqxN5riVz9ZPC/bkC+A41k+QjMdS
SMVIpxBjAZ0+v4uMiMEgBPaSlUvRr9ECwPrcVURBj+moNsZoaQkp+sVnVTWLiAJy
zeDpewpxmMlwTw4DofvcgzmI+c0MpHBPKPSjQciKPXEA1vscGK4JMnOdGHUzcwqQ
oN+kt1b9B/x6H0Fu+tYnGKSiPgGU9jY2lw6nvzwxGl/SkxDuqzuT5jeBfRTSNgTC
U81kpTFCN2ZCLJAJY63dBRcRgN1G5tovIkxxe0DH47leGZDeXrg3aPb6PHbmLSs3
3f30wzmNsfFKOdOwNMnGgqo+k97tAaepk9qQ/eEyuk7DC7Is6ntadzx7AnOaKn/a
IE2paXlQrnnabN5vIN7Vm3bQazLAfBAwVfx1PQQPpxZ0WpzJg2vDiLmFjndPeWwO
RRHkCI3gb3Vu/yiG60LY0JCaD4mNuiQ2VEo2BhdhfbbWXulvWXYPY1oXPUf73Sw3
PmWn2Jj7ae5jNWc9ABEPzUaidBXAV3bMglOhDNqA2xaNB0ztK7mmMMRyyOsQKNkz
jAsD3F73BnL0pDQCZZpgn3vNWlmARGa4pKi4boMIGi0xS0GQB4ZNiTseI4fgAQyK
CyQ5OPHxi54HG/91Em1dG1dh8uHiwZiYPxnTYGuWFVQ17OMSjeJ81FAYRBrb5C48
bzx4lQPkwR+rYW1MD4lx06VQhuUCWreZTE/wU7mUiA6stgBO9IrTmewId3omyGoS
3MROtAWeW5ngQKLrg1E32gRMte2O/fT3IgQI14/4b97zisYvUd7yZmOl73cFSwjp
agcTO1MeoTrYr/kP4bn1ScjWpE5zj4ZDIcuDBwV1VR/5l/sNzoWUURLGNZv20Z6b
u1iGDt5qDSUL06n1ep+npyJY4gVBzexrQQXSUL/EXV1h7S7kutBO1jNmZpIu0EZh
UxeXc/zNu/xJwtwsVitsK3vQRFsEv9P2PD8c8jPXtNdGHwZoDlfzFNRLRB6Q2FPY
VB5Om99Eg4+MhnaqVbsyE/U+RSzkCxrEX3fI74b3tp53515mMJs0lZr9WmMw7zq4
bwtLIb1lDXqj/PJlPHuUtFxkObrgFMC5fh9sgUR72YikfSbeWKRFrWq8+1lCFBSw
NiWTLLe7Nrto/4f5xNZ0mky1BTFjVpvBiEUtfNC1DJEjufJTvGRZldNHssVAG04h
f0yeVZJsMf/jwt8hsC/Jv1/qGH92Fne90nwXPFpuBP6/IWn4e+zLyhbiF1wbCThz
W5ZMcI/SDIChVZDRouW0qWgd2m0WDXpzBoz9oyoC+zeu2pRzDHWCYb9gvaSHTX+X
PjJvyetdGaNrYqKXhdFzygYev+ycsgrQ33UD2ZpOC/MFg733frPfaFz270QzPK95
cSsKoRA1fsrSfr4tDO0c0UVljAcXYCZl8RoO29txuYAF5Zo38hcgg+LktF9Ehkrw
9ZReLPY4SL8pGxZfxKS9sykdwvmCFhYh3kMoYREtbmx3CwU/YGDTfeeyboO8secw
126O0nxgYFlzQlsZR+QF5a7fLWw+XYzIX2pP39eusm43LcoFOEcNl+KOXeOgmGg4
QGPqnaO3Dkb9QJpylddMv5Ati8vzZfiXWAdD1y1/5s58fU+/UAEudbUfqtOkoHqx
YlUdZcCrRuBq7V5+3MGiHwoQyru+TDi3wfb4JZ5OPrvpY/PUo04XbDXGOMTvs4iY
EBiwnxmV0800LpPCutajQ2uT1ZBqQl47aUuMPF27c138lPK74A3Rv8HWqygk7k9c
3F92jhveSmAR5UQrZm3zzLARZU0l3zT7TTpFCqL0P1zUVTn6dHccLVFM8OX6PLSz
fc99cL9n5qkJjT8u4o2UK56v7v7dr4+kAjkZOPSlFmdd+5YnS4il5/yHaCKwy7Z6
8orhURVJmOTwxM/8IA7PAVF+OhoVHZUNpwjXhFoPy1KbR7DwkcNETfb14IMe0fgI
WezDDgAsun0dNw6a6NJ96NqOb0gtUfIIcly0hd15rTUDdCRD0MRGRuDE9AQTXTbs
oM5CxT7KvDLZts7YHVdLZIGyELVmJ744UwguakvwyYHGEP79FI8qwN6eeVwzGiyA
7Tm488+fZaYnNNHthvNl3nRZLud0ooWvyv61KIlBQB8O/Z7+BWcerSCsNsyPI5MH
dLj/W79DRqhegfwjCANMelMpjxUXlSP3zHVNQUmmDd8+MhA2WwjaoFVcMc8PO9Jq
G9LYqsb4ONRHN92wKnWw6Tms1T82toaE0nlSn1LU2EH/+DrJeWTiTiJcdvSj8gBS
8xarNyu24VA51hs1ZygawubZeacUT+bOXRaOULyChiV5i9ydNv706m0xjRrrezS/
i1/raVSgpnIYZtiwToz5SGAt8wQEON/H4ijRUQL1xuBYOr8TvBRqJY7s4stkJh2Z
tvIYLXTVDGdJRNdv4YjnT113rlMsCXndjBDQ9+5x3WEtKTh2z4Gvvbpemy6A/Mdz
dwyv4aueaXh94AqpopjC4CtKDr8rAM40jkn//EkDeNmdLJFnlwCEnnC0TynHH6ut
lVmM+vByatWG6mcX1xhPtarVKE8wOrV7Fs+P69SR417IqnXpsKDPkdp5gKMw+kYN
/XA4pECeTBeWjNzn12JVGfQ2APDbInZzkqFGDQslLZfTgOLbB3y0kkC6deFp9zv5
gP1b9poOyPR9nHQctZ9tRd4zBaKVFITMsh5viD53T0muNSsyeAMAqt6DwJbJio5Q
mV7AjtC/kbILXMbS25kRcIsA4/iBPEynhQ2RAUZxBf+s0LlRyWZsDI57FJIk+t9h
rrMP/oDztsUuJ9vs0dPWRJQ5mr1iv1SQ5MiuU2HqAXUWQ8HLeyQ8q7uQ3LMnJMwJ
GQFsiQoYTexseUrF/t7V8hpYWYlsMCyDtGKcTO7773oiE11gjS740iBPuIAW1GlE
yz4JVN7lGlBVYkISXi5AUYc/eEm6BDHoOOYyTP73uo8n75SiCy4lf6pnX0HPlQFW
5Lsijm91O7QBxWkFbdDK4ynUrUsw3jr1gdCpcZ0ZhC9flbDoWSjvyDmkyLHsN63c
cI2DcY/AhgujyC+LMvut4YBXdmjk5G3wfIb9EDCvJmL/31ge4TSM7UTPyF+WcyhX
9N7ca2H0SgZP7WQWsn7IRc5Mv6Mzz3jPbSFuAnnDMk5bWbMVDtS3rI1EwlC4MLm9
QR3GlMu66aHn4nU4xWvXDsqcdkQlxRahF7KeiacpS/CeFYcvVUBhfvM1mEVod83J
K1l1IWj2gdfQfKwA3B3o8+nZlEMhBmPGl63hFoQoJxvXiJP4ZxmARLaq1fkECfAJ
2wfPsMkYP9thWMyvIxIZaEWZQrYAuMfcJyk5brfab62EDff8bJVbkDyR/3AUurR5
Pyahe+khBSEA1i+W5P2O2Y61MbiYc8fFNgNTXKqT1XuloaLqfnjE0IUAzVEjcODL
oJwfIwtRngHmdpQYZbn6sR8CbFZWpdrp4hTLJdUWL4Mukv1NyxGPOtb8FdChNu6L
IeTBzvVwKuOHdf0spvNg59SkceOUu8lk483r45IZsibF5PeE8eoj/6WN9rjliLO1
UT+LOQV2Twks5N5MAuf5XvK3vfxzAQK6+zWtXBQO/vnX6zn3MoREbUbxRwAg3j4Q
OklrRirCG5LbVBpRqriTY9egiKkaDi7b2kFiSfFQ0//RLUuUU9qguuP8Ocltx13B
kqpIETA4l8ul7luE1O5t/Zfh6886m4doxkSC5h3QjYRrxiZYlSz+MxpoYLevXWNC
pxHCnuoEBSHang6X1UIEmZb415u+yfHz9VQEjuMes51JZujJaEpA66YAue2bRXAH
jghryrvcv1gV7VQSa5K8Z5+gqKiltto0Yb6iCr/clZYyXYXb6K9Yvw6rW7TvBoI4
YmL3xylW2iPXgJjdR8c+1MW7wvsyH3eoh29rAJ6qboasLX6qrwiOTB7U25x69icH
Peh76O9pgjYT/JI6YEQhaKXBDX0gqxVEiieqyXoVrN3eLAjaEHDuhxKiu8rt5NnY
c04vjMKvvhoSEloEpKfuyJ4fy8V+MYmv/lTAPLOLsgN5Pp0cWKpk/sH3PyntmaMR
JkX7EvvcYTmUbDmLEWbPRstzfs1/lu5Ht6CK3WWRqxS/4Xbkac8pwPa/HxGqzY8A
v8ucCfh6+hzDSQuLdun7UTyVkBvVNptRzgCOrrhShuetgHC/tdz6oyLCH3uynmkB
x6oS8sP3gXJX/co/Vwt2EkLangLgt06LkPq8QtqEgY8JnLu6iFEAUjqWlfPpw2NC
GITKpBSvG5YHf8VsauwuDnw8myWFEplpippXcXLNUelXjew+tT4CbM6F8hB/n2ki
e1m69ZyTd261BMy78Y00wIkRPH+f75vZH++S5CFxwczHk3p0HVH/49yohq72CV8m
2Hx/CJA6Bp7IkBTLneGFFRFDOr4hftbEJJclwHYychNdw7YYQKDuiDl3mb4ilL4v
SXmHgJf0g6kSiHCNdUjktacsBaDOdNO5eZJjO3nosNTDG5oWORf2QSuaKF7UgLqM
htuZPCXNzQPWBRVfxvKmXEcXapFxwE+fHdd93cHpg0r1XfwAVmESuKX0BEoq1ZML
Y1/DRBej8lgEotii+TixqCAC3EVb5iLcpcwbFiokuFkVL1eirFE2B7gnnJGKn7wU
2zvWTXtUT8jK9Gsxpp5MyCDHmMDywXELIdXYOmh84v0FLXoQY/VJo5g5SJogD5LF
BDtaurzxIhBTwj0kgnSNSeIwvaMICf43vDdDhF1KDTd0EYyR87C53IVkDbEVcStH
n3VTSN4mCV68JNTJuO1UubaeRmPUH6B/oVWv//4aMOgGU0Ow6c9Xlrjqr60/5r7Q
thobxlCqYvGppnSxblUPJ7uVzLUhPbXS0qxxcAlFPeBotK+D95hhvQHGROjnIqiP
sQF1h/FSoGsV5/Wk9yBmMCUzWF81zO9v2EuHbm4qh7DQdTIjcXDz49VsizAJXxRJ
Ov7uqKoBVN2VRXpj4YJW6ivDEvMMg5kpNc4C2FC2Xr80ABMNqDCcFxZjhgl1LrRs
ho+1kC+gcYR/jynIEcaIFj84fmueQUl8J1k5WC+kSkGReD2N5E1GnjaCUVs1GLpx
Tu8M/dC305sBPdR4fJkEOHIpXhmrALYYaJT0mWbCdNolicjlrItYg2VlP0QpiCZU
5rduCvpTpBzB5ULYJKRc6iwtt9wnnwQmutlS7dsd7AOPkb8xDS3umvFq6/eMIaAw
LcKpeXAon21c/otGNlrM4zcpEEbSm9lY0yZoSnMkUMMueMS9DCUEkyv5Vym9G5j1
0TSWkMA+Zw+uRqghopMyIAqx3lhCW/FJRdaFyoV+h/XAwEEtuzqLe3CUdSM6hQqH
tCDJlx2GWIEQe9ksPr6ZYtQc1G9OG2shmqsLToDd/IGtGtsmiD4wg/P2AjOYiM40
yT+m8G4/nvNTC6Y+FIy8yrsWw2p7ueNy/8jGVc7k44ySS3f8UwWlEpkqg9xV3aeN
Wv5dgzPIbKc/Lzrb694EEuzmIJaBvgnUcC+FdZjf3pV2jKhGpZ7qstW/Pg/j6oe8
bUcFCuMlBnoDh3vQOajtl4ict63m/5WilfdJejjQlwLaXw9zvBUtmZ4W9acF92ln
RakymJQj0duYCM86kSDM67ExaqK0j0Dy1KUpjLXxX6WBBSGwAbhstJVhR9hn1CSm
Nzv3jjyV6T+HfJ5js9O/7rkw+cTVtR9ErSS9F1VQbU2KUd28C/Yf9fZu8gUHpMEY
8uyEFvqVtW3Hhsyq+pb6OBxZGXoEWnVbEsrfJGxwdyXVGm6CuN5l4HVvGNtGrH0q
8OlXqUcMHL/IqDJAXBXflzv6VnFWQd8l7rZO0GQZWcadcPEDg6TVqa4AEQ89ouMy
ptE1SVwFn3Pyk0uDZEZXwhLizWX+KfozL0845gxx7PDnfdtaCRbqr5lkIO0GFcFQ
GtHx4YM5q6g8E2fXT+8PIvF5VAmgVOUXGli1FTqBV8rlxl5sO3aKWSPzVuPAg14Z
bKuBqfL3R1nr0V1KDv3CTTl+/6PKKwqXcdWPXc55zFvlhkI80vm0UlbSod/rxLoc
+qkv7uSh0o00mG1aoZeoLAbNYcxlaH5NbFGcJdwGgTAH0vbquzE6kCFHmg+RZwt/
pQIpxWowshlyQKMNRp1fH5xuzxEDLLVxSJE3RE99DAdYq1WTtX5P1UqwtyNU/BGG
3WOPsAvg0Dz3TPZU1JyWa7Abg2KvRifgO3XstRCEaFQDepcVtrCVjQhQr09yqmZd
kx9BpnhnVZTHabKW6hxbcqH1Ek5n94BCVf/aljepZGeFvhJ8+A6+r+vWRRfIZHAh
odoDCI3TIbrKYz27nuSOVIGeY0kWvZniV1z68XhGmhRBtbtRR41notLOq/wEOgDj
DApSB7dkqPn0C1f+1UAovhy5CngPBAbW9jnJ3JbX1AxneENsIunjuqZS2lG/kpoO
OC2hUS+3wzF7+WT5mp17o+NswJfRsmAdY7mFWQ0VWgPwHKh1uiSkZzVmZSeqbBpu
T456Jq/y0T5Qi6hZLmFdbTzkdyqkHJeGmmwrsDP8587o+AxLkJNHBiFKRvTptv6J
YLQ3Geic5DKdCc3rIrJU0g+VHkDMH34RDNOdWeWpkWvF14iYQFYohqnukwgDVhqk
F1pRVWXomHSyhBWZEDMxvsO3WEyOhPPyViBJKbQ0COKOSHFByaIHBOqmt5qFS244
/rUKowLo8lFpIV49wVpsi39urj0DmwiJ+mJIx94+6xo2qbhPD5bSbBEenRQW3So1
Wv7bMepkJ7Ga8jdg9p89dAWZgNTbCMmlDDx1bt0qpvMKoZ1ENht2b3nSfxc0bAgi
O/e88y7poBfwi1eYXvmt9s6sgdSaKGbe7FP5VNvQVpm1x3CTwv71H3iiMRF7dCRY
q6oFjTRxD3Qf+c8VCe33B3a4/9AapFp+RCwhQ1zoRhngGe3Qpscz55pkB63Fwm/U
wkndyosskP9zLUFNOCqJYgwJUpwe3gfhSnYbJbERrJUwElBKRIXwAmJBuDpxCS+L
z8YkAPgUFnAg1MgxmppbKuUWY9bn9eWD1d2f+sir9NnlqrONWyCH9KmR7pOARTMi
5M20yAc80MwuMcIjE68iVcum0f6E9nOzpXYWlPzC8wVXYxsD0I6fOZ3RpRARgV56
t5hg0HcSobR3vam1eWU94wcfH+cSrja0MQokZoJwsb67qjE5mIWWdemPfPcNbDlV
XkU8hHUGgbkxUeEu5Op2da4xw+wlKBfyr1BDxibS4xBFzFGunuUG+JUkyHrbaf3t
nCRp9Tz1jixT29TopAxkrDw6DaaMiJDOYZVzuWopJtZykmgNdva8C8aWpYwxOGp2
HHmR6eNXrfz3v854eMcFW3fjfwWoepRPfg9DYvleenIvVCXa3scL/s/cQwlfAk/C
sPqMEiQVCsVqlRtsUa8yLu66GPieLHkctIbLDzPBIOFtYOdKQtL9fr36jB8kZ0Sp
PMPLdee2z4DwcMFPv3cpxGJ2GW5CwGSBSBNdIL5ooh7w3maBHHdrg4LRf1Pjo3Z7
FpvvezTjPE8wEbzafSSO+ue0egSIRf7OZEIGV2esH68ceI4gUUOizetFiZZGYeIy
uhfIUtDMJu1YNttuVUhZbODVG0w13imQa/XMpDx6yMfEybWbSEzCyRbHL7MW8FSa
XfxMcQ7UOyMX7NmfE1+FCSkwHwIQkAivx6NEgmA8LpApdnxIlnL6/8A+pTUatsrD
zfH1zV4UGuBH8GfI90HfX5ka0GNzkuC9ixqAeCrNvXTDtJA99JeJceDh4B9KXr9D
bfh4HclJQmC2HzJKMccvbJF9joEXMUhyntvdngaU2e58KffAGQ3J2AFwy4kdEU3H
dMpI1FIhHJhM/ql/HVwjhiCwzAaQ6J5CibX7o0RbhpG3B/F3647jqvUhL3lS3fqG
wYSmHhuMDmD1uooU1lpgw3zKIkc/uGaAJWfGzYMdI7SxW5xjfeMw9KcH8OqnD2LA
dPd1S4XZ4+1LDXSOCqUFSIJ4vy7sZ2wIfeQECprsV6sFRbZ/znHW3tnI0W5eHCf+
fS9Tvuzxi6hTrQD9LMWaVIm5TR+AG+pU/J9Rz/HfGOvIRawferqkEfjV4aKN6wzm
GaIfOsXJpeRCqOc1/C/Gmz6YN4/Y/naUsf0216yoje4bQvsP2cX+3c7POA0Nt0cv
Fpaj6QuZslkrO4vaMwctme3+p5lDQlb5arG2F6PcsJ+So9i/gAuQE6O/LQs/9HmQ
W7pkqP2vWHEntxkjUnEPXnS8QwJTzPNaTfO5nb4oO8Faz4AWZ3lTw8PcI5tt7Z0K
CzeYN2lIkNl/rGfkqCKtdR3d4s4LTgxxSNb8NkmjtQenAkwLRKC6/AL3f+a3ASZU
xbWhv1SYv3mhMJeor3o7yOeIxT+zqoPHyG0lhwZuqINRL5Dr+PKfs24D9EWTE/Gc
ruubKr0CBVgM8EHHUpnVhnPc+Dmu6sEqGaKT6BXbP+vPhNMUuEvlTg9TtlGdGzHa
3ryG7ARz22xm6uKVrqjuEqoT3ZwkfzxFBSH9D5zBVbOWbUJMub+94ntICY3QqC4W
i0efuxECf97bzbJWba10afpWOTlXG3gc+UGfdY7r0l7dHP1Gb04nLo/WPOpiZH71
jw8vXkvUkUos5LDgUXcfJ2nIn+DEnXHJZoKeKX1ZSL5RYPZVDhmzKCPlzQOPKtNU
8VqLJQgpC23HoqrZTBtkhGjuL0DO8KUsPch2pn7rl01CrOtw07XZuwo/qE0CPPTj
DP1Ae4NHEFTnX6EXbI/rmu3pd9SRWvQbDl1myVmqKoe/QKA3yGoFO7k/V7M6unsa
BTl1GmuoEh946r03pIwp6NI4gvMkjY2nwu9yAdIRrxcDe5PaSqwzTjBHL3SmGpm/
yyJ4Fgw47xbKMzEo2pWNHGN9IQIOzfjlRyGDwTJZJW1/sgVmWntNPfrRwXMb9dZp
+PkZSLRtWLJ0RNsS5fm8bKc7Hq9NPHstN1Uw6CMCbAB98Keh2Fmnx4G+Vf1n0Feo
7VIcZ6K3jdjf4EV2AXnf7zhINYZ2OYzOUOPNEP0SmloJT/UtIQ+psMj8sJVzRvBl
bp4ZDHxVi5AxpAr28hJtM6AmY22prplsaM/rqBanaThJF62iZMRXhmHONq+QKDi3
i5AqwtgJoKFtq9e/9GRsrh3kTkzGi53Muh/wHvvRTL+swTrlHVeP/sUJS+Ek7qO6
kKd3ykqW7Hv9Bhxb1V4nD8b24O7yxILha0BJ0B41aVKJ4hrT19VkFLpMwCCzDWsg
wqOpbGHp56yW4yduFlDSUQJ2qGND77qS+HEkuj3l9JLE1AKF3WDJCY2DqZOeO6It
DeJEEuM0JnjG15hJfmdSQqNQp8Auuxx9l08C48/DkX3lfdBIgJ25f4J8wNJw9twU
BGb5pENDJtwy7sTmoP7cB56qCMRPOAMsXXtbKzLiM7sSu88lmS1IN+Y/MdqkwJW9
65mwpqu4GSj34zOturFKUOAXh6V29SJGEY+nUiA4mNSrGEV7hltOKV3KL2yeY23h
rOqz3PkIuwT9+vwml4mJXLZRofFWRnARdnGeNxGdHD/mQr2eI7jkRFmKnvwCaF7i
f9AsATXSBqrjvcM4tLBro6BzjatBkHkcONZBIkttfBgUDRR4BWQKf3UPq9fGHmi/
DD3HvnYoSeCGRWaybTvur61bAs8OJVJB3qT2/4oNk3xqd06f6iZQnsHGyNQnfY9k
PGccqR7FO+WXR0CPxmwnGr+wsZSdP92m4i4l8Va7Qarlrrhbl5UPQmDZTRnhxCKn
rLosKos6xMDPcgpPjnY4z3A1FmUyxPDh14doxMjeUNzbPcNfYx0FX8l7SlrqbDgZ
0Cl9+8puoXjvuzd9HAK1GRUlGaz0f9AcaptM3oJ8wHUa+MIKNJgo1OiX/Gwrs8zE
hvz35BLhFxtqDJY43rB+muB9651qlzZW3STxkZsetlrESN0/cIykZt25SgL6E/wz
N7FBj9XyiNQ/4i5S3fUQ7VbmxnvRTmViWnhlI3Pofy6QXOB/y1gq6uS3ylVbAIR6
o7/GWOUeD9zL34/mYmzg6wAl5/vQEcEUAkE2/8E4ILpQzhtUBY9ssZlNLojSbQe7
fQjHbeWeQq/LRyCM4oylOpwtTDne7DP7KO3OXlAML6M8JLPUayvLtFRpooRNxlL/
KmCoT0KQMGqLXWxiNYldLumL6vRgrlb14CoJ7wh6ceMBbiL1rs+DAMOR2MhCiYnM
k+e324sdkuOpgimFUIgkCD7jwxkqdQBK5WuOiYx8x7yXr01WK7gaUtoItMbcqVFS
CTIDewf0dk6lMESSycuGq1hL36HBrbmDB/ZOyGPC5XtpDUYL40Lrr/W3WcbFpzTY
aSEu6e9/q80yFvLo4bLproy4fgn10Rndh+aHEEgiW3X64FIxyhxBIJhEkWaOWndI
l+JUj9RXb6BrdrvLfjbrutch9NtrB0/HCTD2jiQGPha4OAHbyg7CFx2vdCJeh832
VvOTgqLaXvu4k/sPQjD/RdpmyeEI/UVwOHTqzPOTLV1EDeZBbxKm07ltS0jnuWSe
ySPwqqHytjl9ksK4Zj3/vOtUHm8Aw7wqpOsjIGWntqgeIHgtr7sokWkRlTmb1XA4
ODKWT3202wjzFVmmF4sQ0ZsdOq1zfUfmJCDd8emxoO1u1Rlo0ReWTX4l3I4vBuPN
qaGDd2HpQiGW8WxtmoElcsfJE9KNRDYPGzi+CV5pOQ1FMFObFvWkFp80jt92OmUk
JJqR3tQ2cbFMOf5tMDxf5W8U0rZ2a5kmnDMKQZyC//dCz9a1MMdKgpIb38zREEm7
xEiMqZpGODP61yTkwg0qL7rumKnTTIemwNVBB06yqGuSTP3hRzTWdINoOB07QNim
13JcJO7+kRqnVuSfhUYH8gNdWZ88XgUcHhNBJqp5Lm428Lsz9+iVkAoRz12d0wO5
o5JJbRqQ1afj+e0JNlWWNONRD1eHnexwdcI9Z7IJRBF4MW3HdQ5T19sp1735VGT2
CSVta+zOCIcL9p83IWubvqkziRfMFRES3weYWX5BV1oyPdIydfPA39Q10DSIrsyg
QRrzfgupHvISg2NGNBdYx3TYhjwPnmNJd+gf+Mg1P69Wjdt8Capxu+yRR2GRz78h
zb7ump4mPl+UbJwhaMiufi5iHA6Mq0jQ8Oq5mveI2wGw/0vkANKU6NCctcOBVEQl
OTRW2/PmBrn0i5tS2d9h8xfsDO7rKt/yCNf6NcZAtnNuHDLg6UKIjVMtrxe3GZpX
boZZFD/uMvN6FbRew00eKJzF+NK2Km5T8eIbUB3jE4Fd/1vzs/b9CRZWLcj4njgo
Urtu60ElS+c0p0auSwo2Rg72f4Sn6ekSEvs5FBzHZYenrqzg3OzIM/HtrGINMXip
rHUs5kO+HszdhKHCJTVeWc/w6wlg2iasHnGeC29uDHcUYJSuYXPzG9zNuV5DJhAx
McbwfRpcWt3NHv47uvsf2TM3vp/Ouk9LhmZGO0BZAZfGQcC0yLjf1YVp0lmFqJO7
l43nAeOhZITZmAUfFaYR4kG2uvFOE7Zw8yYeSp42LirIT8gPStEIdrlP0H5tHAvE
Oc45fenXaU92jNrh1R4Bq+9TJdUi4nMLj4wUC75MQqdx8Hxbju8pl5CzM8djuYkC
ZIhiivEk2vWm8FRY8dFNyXcACon1RxYRSp4TaaWLJSdDWxcq4tUx5Xu0AVktWun2
vEgwPUupV6XSDt2FitMOcz7YcczCGUYtGb1289gPFZN5uI4pyKIdn5ZLio5CCSka
aVyarKUgHLHge6rXoteAWgkdTfvYsAEypqBeVu2bPPr8VDFEFZ/l2EzQl0XfVwTw
RwyOA9aOKggSLfKE1WbvU+V0syVqjFgC8OfyGtJ4GSSC5MPyCNDAWBq4sv4MP5if
vnPKk4jZd89+zj/xyqIDKAhDuESudg4iI4kNlx6HPyHeVV4e0fZIkLZyQREdRQ7O
vni4tVYNc3kAlR0yZ/ROabwpqFd6Wa39eTHqtbCPIWT5x9nYq+YfR+tNBeruj+Oz
0ZlioP8zoIBs6Vt/7DFDUX6mDSU9h2meVxz4mR+fx3L+lU7XcX79RfduJ3fqmShp
vklxRc5KOIX06OXDLiGpJbKuFo5yqgL/ajJWYKYKwuybeV4v0S7A+rTuKR+7ITfd
j9hzBtIifyCrxkEhrXa3z/TTSFCrkYY/cDp2K70TuAh7i0QSSizNNm5LOEo/Fhcf
ouy2MJOMspHBblr4Xr86KcZp6EEQ8FE9owNb7Shx8otHNYkR1vQCPhcd08mRCp4+
yNQpwh6dWr01jrEfWHVIFCkfnwtKBbdDzdxJWZXopxClXmmjG60XU24tIZnO8Pw6
21NYD3lvYVToAZtIAnq+6IJzMvNjcZgrU1Og1JpE343ErFnx2UqxxEADu6kBO3PY
g//8wJSCKfQ2qXWmHKR1mdmMe9vvBJZ235WiNthCNbUs5txJ1pQKyNiLYNgQg2Rp
5COwk2gtKMpZbEZrKzZsAQqeWpFw+fzgHNoVfdrVk4wt7TYVRF3FsCHn05yFfY41
mW1ET/P8H/NRtS3zRJD7zaq/y8d0WB8b5zTs56A6PNrDUBQujFd3mWbGbPAMdD9U
Zh4VYcsMB0QExWNEiYtePmteYlBSE/kf86S2O2upeMM3h1nku9o411W3KNpgiAki
gKGoJGrw2R40FtAMcT9zhMLXZxSuL1Hel6NxgovADBo7fTwUHfbRU2yIMeGIYcoc
6mV455B70RTi8j7lQ0NozvB1SdkIimUzhYwkI5J7WtXfF7mYw7cItXsoYTrfy445
0LD4e69oZ6q9rEjesA+VCgGzO4qoTB/gTUBXY8HZ8spel6BgRJaWwtVWcPFakj0P
8RO6oLPzv9DOaWbkLbdpCSVbKmLvifr4VK2PNpnXA01xhH9sp/z//Xu5jlH19Eh+
BdO+0ztQ7ECtCl/dvoEFrRWsBn5ptgIxcqn8oVyhq2waiZlThvn5mjKz1/lLIkNr
ITZH6bx6F0SCSueRyE/rhFbV9+I4dybfbrl4CrbVBFt031PWcOruxiFjh4KLc44C
cvzZQ8fRFcnmnyp0f3FeGHLHUafiqGvL6HERs8ZS6icAX/xbl4OR4eRbBNEEg0r3
+WCkBIE17NOhwQNWSulLUb2LpkV/r5tRR8TxI8uGLV5cfRu+AdLHyO+I2YQQFZYS
qjAXW/8vY/qOWWVZHUrXYcjfNSHZot4+zUdXaQ3BXaetetHQvQ18rFyf/QwV+g7P
zi2gxVeWuXCh4rD6IpEpsCu7R6lw+ukGsJmTtwKOoFz64uKFkMg7qlTWbjHd9bM0
yC+RwcvicLYJy9P1vP7RZmZnwAnLixqMa2Cuxn1+wY3hVgF58+lH718p6AN2cnFH
Gb4E9Kg1m5An8V9khl2653TgNHd+7jqX5v343v1VA3r2WqUWiOCljT7/4IaoFvvg
bqH3ddvMax8Mk+LRcgVrRlYvbEgzVJf8kLzo1KKzRSNlZqZulKIQodUfPHqBQiUw
/Fy4/7TBwjU7LJx2rsBbKvZfMTgveQ6q5672BPvuvSUsCN1xbdnd109n+SABfYO/
LNWe57N0nXe8eXz3ltwg9Q0FRRBtCW0lzDE604iYf8R99tPDUBCeTfrYL7qfNTua
h9MDUPr7b7ZnXCQ6ljD9T1kmnlyEHalI5Wx7jsBz493i65xfLZyTPQB04wSVl1l8
n8Or/sY5r/HsoG0bAtLYsRpsJtXGA+mjtRloCQEzRS7X/GxPXjtoNIuwDxLoJMJg
EnqbJPi5ktlzr6Z/RGPEioUoiDHUCMPXo318aETLS7vRrVzvlU5/GSq1BBMLBbJp
IQ6i/9u6cHV/qxJC7/iJgwXUNFHvQHPAyBmijc+gQVlJSc7wNoGIkU05MappoxTp
tLnriRQ3//ZfxGHKHN3wH88QHLmDoLHgBkWMiC5c5g+6j/xissH/YYgtmv3F5SmE
FiUaphlimCzHN0Hz3iwezK0Mv8BJFbVUGK0bEVqXCY8+38BepPqGRbK7cGjZIjeB
9o+BjvHZyk7rnnVp5TCq1VimH3PwtWh13FQHc/yRaUrWawvMU65dBi+Lc/SdEYGa
81e8mv69z3OGyJ2ZA7jLSVkbsrLXNMVBmuT7kZmMpmIeXxqJCwU/A50E78TThsct
LlZXvZBtBDuWeE0Uhl9VhNhBaBRCD6cwAoPkJuroHCEDZP/h8nRJk1ZV/njTJr+f
kIHtOcR6PkD4funeFKa8WDGQ8myEiKFD/AhgssW9bmDFAI6flLdA1/d+0/0NiAOg
Et5NE3UbfNchjawfX7m4g6PTaBO9ibm5mW0dqifRtMa3APp5z5OYtFVYarcN0AnV
RgkYKaYDmXgX4CDQCNYqEpKJZtPSPGJzTsD4wzD8T0+UD8kbKTCGmkw8e62rfJlL
jANAl0KMaDLou80tkyUpyxr95RwMQPcxrjeL0spuOJvZIlOkcOdIA/Sjp1AgCaAA
Mdcm+5Cl6MvKXy79bBoE4XJmXi+2Vpx7/yFCzTdsJCha/w36qpkKRuha3HO6EkwF
rddllUd7nSvZjF3VOSnKB9q//xQtMomWbqCmROmySd0+D/gReWAmqKWGEJJJjX3B
p9o4uM4BR3Hdnr7Ugawqh19ndOSR13tWNUe7C0kCa6viJMH4z9QjG5ToNY2x21mD
jDH57MtiDyCNaPOGJxcNuEPWCWTpIJ/DsVwg8UFP4h/b44d0X+qNoUsQtkbnpALd
wNDmLK5OFEsPKu05PJ35nt0SESVZEi/Yj4u8u1FPQ8DmCzlCf2LgcN5ZHGxY7mOb
MMhI42JcCbaUaImGBVY5gylhLu+JqrclWEGMJNMVaX+OFQfJpcuP6y79exULDq21
7kaY/DyZsXkB15cs9MPfxsJooYZw11arm8TmKjvTpYxsXxqNa7amTVApfXGB8mRT
ihRyhKajp2HWTldUZqqvvFSO4zYe1nwgscIoA677w/n9JFJwJtAZyHOHhQ7LtJDU
TkA+kVnSVuyxc094M7UykllwXObTBbufnYrmKebD12rSSXiB9/waHeJf1hyBkEqq
mNAgh25l5g2zF2DFBNQT89EUSRIhLqcRivOWNr28jXywymL1LAeQgoWzFrcEHF9o
EYnsUJvsg7W64o7wMEgaS2CNZNUphUktroBz5AazipryuIZGmMh1SkeyCh7pVG2/
Su0JqyJ25m7QCsopeuTFPpaok9izmtcwSGeepKGCrGO3IQPwEgWn2rDm/XMD4M9+
xGgF0x5uaHrlSN8KTgpcdh1UTIGx4E/EAOPOw4wsFKIhWRWy0s8XrlcOOJYh5QY+
Lt1VJ4EQulcSIwAQ/+9CbDjRfXONJSXoXE2IAzhKGQuJGxeRn5tyjUEBZXsKfYnV
Dlm02+teNnAugy2qpGlFCZtTXIQA0dcNWLutLhhR3G+cT0QRuLn+eZD9qbo18vkz
+UB8j7kkvCtilBEMcsVKZySU2fdU2+0XA41bEs8xBVC8rvIbWRY4jbJmPJ/6OqRE
42Kx2vf6xE3nzQgNvh1a7yqmt54uHQqiPTeVsNApvEKSMQnZs4vpaQaV18WfEmyn
l7mUXHEIuBkZhNFqWYVF5cW+xLmknv1aqRhkjlET5bleU4Z/EKXP7ZI10u8Mqkqi
Ryn0CfRccfpPc5uMYn6OD5BEzUqbcIS170UEcnJm5SFrikklWqJv5hXId3Y5iExt
xA+kRocklpXS2ZfZLp6y4dK8KInKxUMqwJutkJXEfjAIOxfFhOfK2NImpj4PjpdK
gx0xbZo8nWMpNFxb1SBx57Zpk1XCJfvFqyDnHQ/kgf/kzfMvub+rfS3mf8mlLMEy
8TebpNlam2Odg6fPpB+ecIkvJVi299OQajpzO4fqNYmg2KAs5ezY0h6Lc+a7tOG9
lRLo6Cc4iimNX4zptA+CZjpR7vgmmrMmIpjhGsEaktvzr8ydsBR7AbknZ/TdNefc
Ebt/gEsryMoWEkrQN6d2KgkkbpGxKyHlPXMpNkyT7OqRDi37NWGRurpOZe/oKs+H
kH2t58kCk9BxmGJ0Rb8hZabnEJtX0nIy6KqH9USyhpimzOMiHGJ94bOCV80b3t3X
WIxF28Amts6F4+RFfoDD/yipMCiINONznCpiXSncAkjxHskww1vbZn9YecnX0ZzV
s+Iq4txvkuFBHEfcPpl9Lis/WDw1XMqwjqnZgKFDCf+3B7Q59W8GYQqh+jJym0fe
UAMXQQCbxGtU9vXJUEKsYYc2WYNpmEIIySECuaCewxac6rSUf7/O73cxpfUAGZBw
lK+epRhapX4Lig98bqfCoB4rX4D85cN4j7NKdhJQgPVrjuel5S8VrCn0BzgexAeb
XE6jTaMz0SCwy190Y7/hUGBUFlFuRqnoXZV85AfLIdCrsl2w3SlEBEB3U10kVtAl
c7OYFPPH9AExQ+EwOG02NPNW57I6eE6EVnZrkcA8Gr4ygbHEZOSrWL2mXn3Ky2bz
xGjHBnd4Ri5r2jkaEYrdKpQlTlv6B4YNQgTHH1n8BMvdF8s+3xePSV0eOj2ZJuyr
gKRPI4ArrGe7gc/hxFgxE+dbeyuLny6L3L4LqkAMpcNK8XkZygXo11cLJhXMxkj0
wNljSq9CYQ91KiDCozs4VeW5YETsi1SwnSMVLjcC5XqYScvZPkQUgM3IM45MSQJj
TaInxmB7W9b+alj292C8uMOR310ex9j00fEn2CTeUcltA8fGPArtgZZ7SV5HMMse
OKEe8XPpTDM6/6EDe6+eIcnE5Du2ZvkTF8FnLvSRy95NAARxa77OXbpLR/4rrkA5
q0dZlG25SGRSbOpyQ/FwJhDy0nmK3aZqD+ZKrxORtsa5PxMJQ7LobSHSyehSVwh9
x3LBVQgPlHB8eYBGQZZ8dyniDFm43h2dRGW2BtbibENat/QpkXKmFYxyI0IlfNx+
T7ByDAH9iL2qlObJTWSmzEOexu2pO8uPJ47IfjNmnkv70Ue9WFjsCgF23jY0qqaE
l9Xe3Uxljyy709SMOLnOLofOND1fsv6aAAtkmUPXa2u4FooLI4nwSyTRF5BaHel4
wDtSEyZ+oQcjowFBRtGLQmPvHmqVbaNDjxNUkFmTnQDtqZ2xpnnWoVvXzPT6fZhJ
ixduNuI1V6TqoC4XG5rLcSDpPsxUKmEqPNAvs5nIzm2hMRmBX7STSZ3rRljf67lw
TlQzwOvVC7Be9bszT/aGgyYEsNM5s1n7N8LstP9LXWFs/X7wYyQhg3HUA2jgbpSz
bJGMHC/qEQ/T+AFLXg4ZvbSWDh9GN8w7XWKiKFmRmX4qFOqxkdY0rbxApIoQaqJ8
DNICOlONgeKgeL79PbgJE4uUgV9X38CaLlD/R2I3cd5jVKpR9V2iBRB5V0ByIuEL
4+WKC3fIypztgkDIm1T/su0cyS3vdPKoYwMIagyDgamrnlSoy+jMD4QP4p6TpNlP
AhrlGvKsptlDhPiS8XriMvNjanLDoWfjDM7nK2oDGsx2lqIcfFK+kelSoXGqwZS1
eIVVH4Y7PcrecDpx/FjD531fEYZEgPcd85DgK3or0WlOQW1+QU3uuyx8cZrDeYJm
Upcce2l/q+Pb23CY5aw0OBrVzDzXoB58fa6wl9fUeC24yk04zcxi/x4gqLG/eqPT
/yw5EsdBSD7txWHsSGwwt4pN+9sHha8gxbBvxtbDhXbbvgD3aLKBdmSA6jSC26+K
nc3rrz69rnkhX526b0JI5p0rtd0iry30fP5vCEheIgKXB3YoxTzo62zfK4R2BskK
l6C3QTkYNtU2OH1LE+lY3O8qq/Gi2SkZTT2fNPzVm3wHRRnpihkx0iSJa+Q1Bkph
ia4gO18Kc7EKldMSTmYkYwRO1HYrXbidAK6umXQFEOWatsqklIapm/HCWK1fvnsx
WASAPpspd1wRYEwth2O7G0V7ENRreYwg7syBxbOgSOW/i6RdR1HeSVK7gVGmoh/e
f7hft6Eb0TU2NoHdrY8/J9wQ5cuS3tvmjz/B+hOO4x/6/8PVFcWf+5qbX0p/JjaE
jon0J1q9aRdBAoQEBXEzXEfYWNzUR7yHyeIyqXvpIgrd6FrCe/HqU/9fmm6BIJYd
irKiTq/YYq9ty3N+7qvwmK7u883oEhKVmTiqs/gdR7GVTlmm/a8bNwoA5xb+Yvwm
tG9DFwf5NFn2N4/jnw6cjBPyhmIXtW2Ih/rMWnwUZs+LhCRAFZS6Z52yfMYrBeAp
ap0AYq/jERtE1Z4eS2JfyFGdpyUgPqw0m09y6V8lNUUyZjdYcCN6ZzsUC7qTF1sj
PBLr+gqfMUVorqm0Rjx3VP5mf2eNeX2ccXLbLYWFbPFzDLwjHGe4k9/dxrJ5o/0+
vxZL0VTn8G0GkXtB0mNCfH+uVVSwdHKI8/wqGUZfhneMofBtWx1boyc7a2myLAED
2fhwHMDZA77AquW7g3CeiXyxSFkebIqFEQS4XGR1QjLMLWyo+qDmBpgG0hljyo6J
hSIfWb2wRqN2NprMNsAxtxlqGuzl2U7g0s2Lgtfh+8zS1F5T6Wgb2QV8t169Eo7s
YOU0QaIM1TuAhF6iCUPW4HisSNd2YsaGjevhzDTu3/H0KI/tE0wmQAyFGCIHfMHm
IGSYAeamaYFCziV/FRw8G2yOU0XUOgw5B3sopSpROfQFEu7oPa6Qhy2xsguiRer/
ObGDiORZ98FzTPtS3O5BsohxjIP4QqRanjXrAyGZyza6SZ+A4bev1cFHkzsKNArm
TJ9ZT7SmvgjrKIpxmMhOEFU2jv29egp3S51QYtnIfCmi+RJQoWk0AvJDMHt9oWCW
j2lfq+sMrt6Naw9fGMlyAQrZVPdaIu8QwBO/b1r03cNo4/YvMUtvmG8QJDBcC6e7
n4MQAfNGtv7Pc5NIVAHrYeGIrXWjFyNPZb2Ef8jr/fJsULgp7ypMxQJubdkqEezD
biwFuZePR9d0E2v0GmOCpFeIP/nq79jZOpZhBCss0IEWHP4k+9/n4Bw2T9b7vVxp
KegL2PngC7wqMObtqPH45XRizmhTG8NSkByUqWL9YzfiRj6gvvDd0yV6Fl4zJsKI
N9UmYHF0AwfoA7ICPR9DYaQFm2RD7aB28X3J9nVE5KYaoTFUro0VstnpB/qO0mOu
i3rATn3G41PlhNMj9z6WGlYuCOAcgVg7+Hk96bTTcMzD2BE5d3vFH1Yj+vuVH6pc
7V/9ZTYLaDGszJr49D9mx9ScZy5/ZPYy0XNldLQNu65LOALEpIpfkrtw6qRSDzvV
7Xx4TTt+m4ge0JxzQNF6+/2XOtOZ9CisknmWMZwFgoGKmLE1eT0W/IA+MR1DF0/D
sDDIoqvjlwXHDnXpp2eG9wpsXm5zmHlGcsGBjdTKbWACyqNQHOKEPYFXWYeEKUOF
9psr6/Wzhatwkdxqyb7VimE83e2WFn42Fq1+JBvDH4KXmpRD6s+6NE10PiiIKLkz
2lKRvR9gbsTaLhBbV4qrS2laHmIjDWl1bxBbkz5RP6+tWiQJJo2+smIJcCFXEjAu
97L27s37cfOjX9/ZMsgPBYUhzNly+cGDKiPckdgrN+kz/djnMExpg45Jgu8hel+E
Ey2rYJeE6OkBsoGNKmPZfLPBZzPlPVNtKK6yZvQRZE+MW/ygcH20GXPfjQEazrhL
+7jiLj/bnIvw1Ynw1mZAd29ai1R3vQBM/vYVnV4b/qytdxnZTBjRjKxM6tDxIERt
Hppw/6EE7F5H32knIBrD8o7t/SaGMbo1o/UizLorqcDSlUJb7l/+JhoeyIAo/MfB
bGudobrKWBteAb5r7Taf/U4M/TweruFhNzaBGuGAzrF/4aPZrYz/ZbjcZ30Z2H16
btrNu+3zdHdwGp1BvcXKRC6s72ard+a89HGYGfzVSozkhAdPQtTZIY6A3OFao4ux
hootiKDe2qtJp7lSxTx+ySG3f93BWgYffgn6310sUzDUSo+vqLg5tHzLTZxRyiGy
07LDLReqEFEzRqGD0JqYoXmNWsn3oPunQ/Ets4EEH1ys6ZdTP50+tOaV+lLddpNZ
Ofok6Txf4TG5k7mH2o7bA8Vow3HBGSOQobynXmPsRjiTFC94W9rP3eqFZTchVH6P
wm2Ww4e4Qt6Dd4EJFL+KKx0AJaX2MWrZIXkjZTSx2q+D51r35OR5xaBIjjGfqzyR
W3dW/V5k/oZMv8Balf1c9lEPzUnc63zMyP0TVHha7rttZQvzOUOR4M5sj2DSmIaS
55pnzMbwgOTFpOYPGdA9+jR7ggOLu0XFCYKhuofaXRTv3GVMlNwP9cGNs1vN4jS0
L3YS8MHJzcw8TDq4H81GH0tv1GwO1dGGcFV5Nh5bd8QSRwh+kweMf50vxdIm0N5S
MKEYrkBTyTASXLUXOFbbHUCQydqgl77D+05gvgAAaY1TqX7lO8vN/nkpG0xV2NvX
rr6VnNnBcMvA6+/C2dirr+ddMh8Ee8qbRiAb0dJfk9jGwdMWdr78agB/cOKbv9+C
naO1xBoLyay6jte1p/XiMtxcVR5foUXmRzROCY3vZwL/8ty1pDZIu3NoRuOvypdb
vvThr3jFv6/9n1kVlBQUOaaUZKDZ23EhhnIzbAa1n4njaLU+Ac4iHPuSjpaK1/Bj
e9wjN9H7R/Pu2tqvzXCtt7X5dFwtRCKQ40+rJIT9ek7OFzqtw8gBvVPT9qZkKY3N
gBHfWONggORn8dOGmj91VKKne+W69HtqnBvb80NixpcTHodfk36OJSNfGjas19oh
iJq/atjdhrcRkkalqJKqsR+KPAXoXIy6czvMxfLQ3aCxb8gBL210rO3GnOEW8z3F
RGSJenr2hnNeFKAeEs8OhkGvp/CccqtJkjChXs9AjgRgiuJzwQp4ssinsVTTe2xH
DxodkddmcOmxh+wrvstwy2tt+nFaxaEn5dAJiVUbokjVfGMbbqyG/qim9tq24Ajf
KqseFx7rYvwytbd7e//mwHGY/hToR6LOWq0Tr7mdqS7ww0VY53sV1HFzs1P6B1pb
5td1KeFlKKl3ebXATIbvoZBxjXG+CZbuJHJdmgbx1aHJ5zLm4ZH+kTmxNx0/XUXu
0txgq/X6aORQ+iK4XZFU3JOEC6DSOw1lQgoEK9M/Wvd9oLzgwW2zzFpMA+lELJVT
exbdjub+QCWFVNiPnHriYmkAs2HrUVOnhemLpakaMdWXZajLOVD00TzAL5AbVxrf
Vy+tFMg5kNEfVLgWw3obTvNmvTqC0Zr/6zRSZi2aLSTSIv0Gb58CiByJbkt0gjZ0
dKIt8Q/R4mytX8ItrL2xrHkplAGz6zg9hWaGAfL02wO3RgJCXUuSAiuPNCdmL5N1
q1MU8ROElTgpCyGJl8PAVcUJtVIHkdXlxaz4fIzhU+N3jTjn2l8TnO1I0fvaMLOa
4C/YkAw9+RNmuIdBWlhN6E9qHDCR0BhVKIx5MhKdL9hmkyWTD3aggGkBPKX7ccwG
oO07E+Xghtx7YxwCKuQrtDa1B0Kw+UWqP3yOB9yLDEEmnBvIKTIbhaSXMtzr/igW
oYcw77ndx1k61v0kzpGlWB3Cr+bs97IfQyr7Wd3YSWBCfpXWT/cVPqHbCCp9GY0C
X2Tj9b86JZ6aa1K8iKsDzFrCJBs7LhmfvpuwCbeJACMyp/7FjIQDxANXIwMrca3f
3P+sxvbbMXs/fYqCz7u3QhVVR45DmHVNrnY1W6ytiCEj3OxXjluyxJ4IOZn82n3X
MvvFCB3yBWpwB/OIqnYKYdQKRukormt0N5OYWdqHY2ft4so5ZXJuWGznkyXvaxTx
1cTIE7jKWs+ZMDzeI/yip02bLEs3Rgn986AS2gqxFRFD9cvugG5uY26h8GR8TL5l
A+DhzZvaP/jafv2QIl3gnbhkLBVxuFr/CrP1tJmA/+p1gNoHNgCb2a9+rVZPgtKr
Aha+fOUJF/MiDDFbqb/91kKjnu54AtCP+tHKcsxfD+7FTTcY3uAekTaVBJIzOAOR
tfzA8HoPu7yhYCFoRT5ubTUz6qjy/kyurylHjYcwLL4BVJricbtzv+Px/yhPP9BX
JyAFidS/bncce0/TcuV2FUTyo9mjY17rvijq1+00qbjbzrYl3aq7E3Eunr1RHEfS
0pPwVk8h6bY8CRP5pgwmaxQyvrXqQZJ9e1HZLw+NwfojcFfnTmSQMrE5E9Hcd6u5
Vq+8gx6YEnz9mbUAD+2mdxAy6ypznYqDKOd6PT3bPgb3cAnMhTO5WuQY4yXzCoo+
Fsq4LCe26X38tFEEO/yK3lRQDxFiCoDACBnOB9MoOpSOlHZHnVQspNGOaa2pzRjJ
lMe6sYcMuDFMRWkxfkl1+hhCwumYqxmdbT9I517tlwoPvFLAZak6YihUSROC2ist
ORW8AnpJhtlivZX1H8hFoo574wmOGuwXQo1ear8L9s+224p7b5rNpbHu5Pr097Jm
PG5PWAISUIrz7uetzWNI4LYBQomD2uK6ReD4AEnJdEF/5FFzhm4PcsH/jR5QBfS+
uTU8vqlmHEHBYI+Em3HceiRlzbPrNur22lXEwJ3jSicjGWNUcn/zCW2aBzXNvXOn
qNpD9/ZjuoiF2Ll8oNyPTFWqSAt+9LVrkz6YS7zFk2ZZSrToP59CWuq4gtRpuQda
89AwfYeh3+TV82SRq34yYHxXVJIDk8e6YDxVPOwbWWmffArBGgsYqkJfhLmcxjxf
EJNvY1YoqrQ37GblGKoWLcm6rMkT9/G2JTApY4B55XvvRCUiwfkD29ZPbn9aNnb6
aehv0YYOOfsF8WDF9uBnsPiodW5/FcamYSLjQFNH7SrpMursFB4XTQQeeZiujwL7
LuVM+jBZ5VIEfS3w/CqYrz/mM0RDEL41CNPEoRXODDTPO6yBu9xI8ZiOF0xYG3yL
dlpRBW6812oiovhQ6Ff0luEnOAgmO37B6bGh0SpbfFntQ1QoZvTyDea+7UUwH5VS
PVqQpxvlE3aflebOuWLwG+alXk0vtafHrHYJBtNHkl3BFhCTV2iItFxus0JZ/Vn6
7J8pNMV1L4lLl0j5guUlDFF+j9/uJ3w33Na5Nwzo6ZvXFJ195kngwbAqIJnfdgpm
nTReQUjW7OiOkBvpWgX5OxU2U5PAk/LoGeq0eKO0HJTR+nHLsIQj6OOM8CP2bCWD
+R5AeCb2XOT3N04uGJ6SXPjKGZYPB6MkonHvY39QwYX1JZPlZNlHQ4Cr8ckBxZKI
6oxATnKjmZjLUXD57+9geWex1+iUQM4thtVHj9RTPgH+VxSfP8iqXIxeNFTkhpnt
NEDyX8RQRFUMWcAANgAASUWBBN/GvlctM+zEn4hVLSTZ+VM+o7QHYEPniUFISCip
1Akh2oDrfm+hB1TrrjWQwmIVjqPA/EMQkZSZlJ5Vs2j/ZhjkWQUDQlD4+UxZ6FRS
M/ypC3E0pBF+R/yMVarnn54xz4joFQCZLrZdhmne95QHsBI11OK2KsyuZ9gwbCPC
sjivlYtqu9TJm/p0LXibtV/FNcIIN3Z33R3BZ4i0W9UKCYJUnVp4km1B/IPyWrIM
ajLTkCkIxZZ22U2bVT1+xQPT7doO9YFRKEnvn/WTICL6GbEnQZBGMCZOdMbKNknn
gXq33oj0IaXaU9FcXUI5fVyftsCRFvywZyU6tqfTNY4tXiqyMUMCHXQoXwcU3K80
WXwtsVl+TlP5N2diNMcLYhky7K0f29rfMWrESzds4qM8mugBU5WFsxIoFmobDZmr
YEj3rnAYl+EC79LrA+3RviAYeyDxbxbnkCsM0iGmP85w1FgGXpOOTndZK8+jzEhz
TccczjaFktcIaud+MHZBNGb6Q2kEf6hiHVfPVQ3cAKqMBK4nlrUyuAO9h5XdlLzz
AFYYRpFZpr9rzOSR/inQNd3he6SfIwbkIYpJIgtyROY8l+8F7PdFvwI/kzDq18IN
XW8SHXPu9YlkPN1pi0mvOGU5JsuqGQMf1HEWeHxQAJZe/vRb3H5d5HD/Q4VGWTb2
XPwCJyhFp8VDRji8CBNAsPK8ZuKymzAvpdrc4wG+YzmPQSQxGp4njc8O6EFUZnzX
H5AHgq4ICsRA87y19ViQX6jpkZ15qgAuhGqcohmyEEhZsUYliIz+bA55Z7mbdEzg
V3tO9ERtPqPjxI/p6eY8/Wp0c7X0pr/3zXH4U2urjpNUS7KdH8syBOH/7pfOXMrq
DUMbythrzCfagAO9ac9NbAV1BRI93cvV0h7bNfzqoRWDlkHiUiGCeV0UwaeBDaEO
XhiqT+GynWcK7bdCs2vXpIZGbb2jkjX1KZpKcYWkhRsUpDI3UY69HtIR9rJxHM3x
28R5Q3TIjLnggML+RQBfi5KJr45W+cDod4c+l8nCm4Cciod247iv3uDdJe81ImyI
ehPbmsP55CGjM8uGijmB8MIWmkxnaSFpjoYwkZQGjbvgTsewljXS/7+EriOXQ4Yo
A2Zsh8W3cmQBm2aMIw6IabtctE1i7W85tgF41aA35omgYcHENEzO2QXIZszryZhh
uA2o5ybX9G0krAxsgakW1WAu6zng0bcar8IhHarx/bIas2TVXCTT4ice2jkmKGM/
1IH69qQh/ivgnPRrW/YU0zFBuU/EpPOm13akjGSIBcFJqHgcetMbidqC/L+0U01V
H63+93xeClFCBKSD2bBg5lSdDAguw3bXU6B1HO3YQLNMDSVxKsSYinYLb/Sc8XDO
+1bUebTna2y9N+DBhLp4Ruf3Mqk0/pod5QPMMuQFngPPgoTd806b6NEDTdEobAto
H22+4n+HoYuNCQ61e9PlHUMzdT1kTNpv4Ay/rJ5tfxonUuSBNfjYZuAWtR0WVrLK
wT8LorShYk5uW4kqTxqCwr9V2rw+GyqutHj501degP+zzkYir55wCRv0QxFPdE0B
Oye1Xs6F23KdtH0UVXqm/f+O+imnbtQTEzpAa8ioUlkalrRQfjWeFu6ueRPy/+of
4DKBphFxfOmpOreTN/W+fOiUJB67uLP13EwOlEEk1gd06GqmMT6/dXQ9Vveo3gMJ
7JpNz0Y+9+/lT2M4wNzNRCR9umwDK/bRgv8V0hk9/3SoAkOICLTMmOtDSGktjXca
4vwDyyLXadZgFQgUcgKKqeH5jz57El5XXsSb3eGv42KHPxgtjU495Jq/PT5Cw7b0
AwyJhqqL+JIMZ4eEhvtHKaUhHHd6izB6V6xxUIwYqVsC5wM4pnwzRuzCBHEAPnvB
RPhcG5jvmMJYuCoWl3Fua+DG/RiUdnPF4FID8/4rI+ZWODEhiAx/VdFFWpwM0Kku
F8/Eopsbjxt4miEvt1Ooe8u15a9ooSvvhp71ASKo/iSwWF2j6a1o0UeiJv6S+buZ
3fuDlpmA1sjBx6vn8Q9VuHb6HGE/shqLSZGLaTQx3qSWV8J+FjO/dG9SSjSgJp62
65kId9In4Zvtbs/nuwU6Z/2KBBhYNKPKa86jifhFsGw4oEDBDt0YrCYl3kQ2rTGq
DpI/yYIc3eT87coZQyi+aWsszbArtH7IKnfQWUyn5vvn/0E2ehuvFYCebfVZGTLe
9tVmajj8G+lVjlucbueWNJKj7qxr7V5HSHSLjoO0WUHeWqHu4f4usOzwYiN7ikAu
xZoLDxl9D4vhefpd7zjUV1SHd7CISO7+6pOZ6Fwho/IpoiStGiqfmypcCHT4sMgu
vWJRKquZ+zpO374VXS5kOfe0ZyiBz6yBcOen57uYpEKdDTQR44VetwAtDP4PUyUr
FAMCU9osw1Ql4x+75ZS6+9S4xz38jBCtYWdXi8vNiQjZO5ZIk11QAO+Qef56p8XT
Pop5J0yB8sp+6CkeirPTXlt5k2oHE399++kNW/3O6WxLZIHKctcxe+qnO8cym+xI
dRHGuO54bHEiWdkMf27lgWQomaRQrd6GN8KylNhbBTfg14oMvVhxrsFZo+8pgqgv
c1T8oE+jwwSWOts+JceIQo3lZRZtbk7F1l4xZA03mn2Ur/iUkkLFXdbpVnjnqdgK
1WCsLBqMERLWNnDvSVaZ3wLtwZPckm277rOYrkouhQNSG8gbqs/LInOC21Ud92MA
AA1RdsiN7XR7IW+7e8okwqmhFnsoUZUEm+uQlX6Zf6okTwv8A9Wje7foFw8M3Jok
Xp2bg+vEyHWRuO4r6C0VGDvChVpGYiepRqHtsS6lJl2bC9cbMqEHLWEa1wgUs6Z1
7P0M9E71d70BHEPXemA/RaNGwYgXv3Wq+lNe4ALQ1SMH9QK/t+qGZcjAdUvr6Tap
m9ykVWY/MBBr3dbOIHgu6tCILOByc8051R9LI32bhHY4RUpLnN8A5EYl/1AKVfGg
fsbt4mZtl70mHzz97qfsw9bsYcMkGKP8E7bgkCKgdFK+b0I3W4LxBCbBoEvAbCbT
qBPNmeFnRmDGyRuwFN4X2Z+9u5eJGeAFFBr7hcCYxKPy6Mu0lABIQDSWg/fsT99t
NoKd5KlNd4LL1S/oLt9Cr73RFnl30i6auU2yN07U8CLR7/WMP0PhZAH1vitmHLZw
qfeYoe7HhAs3S3Z/fks1jCgGUUFCEEqi/ZrfkuQ8qTzl0AYqYtBPM/pSeQXe59GG
NUQHiCfEPq7n1cFgiKlfTcCeUTJN8koKAOwognjg3c3acnIC918AsvUgi478Kpu+
qra93Qt+ep0AJeno3BZCNelqwWmJTa1r0XKSLbUo5U3SwbxyzcndduhFH5I9fLTS
Bi7lgMZMx3i3tGo7dC2PobE3lAaB6MDFIJgpcnUOrgagFrHKuGy6begPzjBPpiE9
6qCNNoBC229J6vpuRwfauykN8upwq4qQxaxKJa10I8nKtig14FXW1dL26XUJEezm
oWlSB+R9e8Fv+mlG/4U2WI+e0VNx8Fie9cw73Pq8FN75mTDiP1zcjZIsszSsUbEM
AZsuXNCHr35jTrT8cgA5mY1N9UnlmQvzAT2fyzH7w+OEIV0BzDtrZeZPwj+la+1Z
E/9snn5XDayRvyrXgL9/Iw5nr9aRYeJmReS0IqHHGWu0xtMxmZ9OgKaHG4LbGghH
1Amv1yJGbvUZ2zcrJqbtPUoFI5z0Z2+KAGB6MU0N+J+Fc4mxSk0fuSo2IiHeS8rb
wS3pL8FctatrZcDhIZt+q2K79pPU7pIYtkWbaK0h0ohL9id7S5NgjE6xC4UBwqHh
dAkYyDuNnpR3jp3CcslK9DjQore54WUzslVb5TJL024BR+p7x0pZ5gEXSZU1WOAF
lDnkX5nchhkUSLuEVsJaVo6NdlzkPHOoshK+0S1JN+XBUTY+byMybRBUmJp8O61l
UznXEWcfTjG0d1iOGElAQaIl6OZGeUfrWXKXPRWbX4YGJe85VVTt5XYWx9D3x74L
O0f68mR1vMv5v+r2/pqVgjvzjTgaej1XU8OGafMP5OPN/fUyIWr0hUTfABCpgrzj
dWSpOtxvZ6zNwdr6t+9qV0fxXbqotpJi2Z/MAbnbR12aJxchvQYAubtKcs2gVXJf
3VslZDn/VWvdmr6BRECh4rU6YmasnFvRUojxM90dKPbo8fcSLqK1iR0tsuSJsfrz
JbvsN5KGiInamAb1+MBqMc9xswmiyH7jr5BpppBwPBV/bjfpwunR99BhcnShh1eB
5NLeAepbP7tmhHrV3rrr1zHe7idawJx3ylaZl6bBiU/yY9MwpzUVXuIDzCHchaUZ
Qna9EpNNfXL8CbwHiNoDCocbqegn9Qgi/Y+GO7EyGGqDxqfhqiob6ut4D9Fxv+TE
105c6J1qzxnAHU7LunGn2tUBMkL/JCARVnKRBV18YqQu7fWui1aZ5lQQCA2P/ljk
EitgyspEkhoC6p0j9/eMhh7roU/eU6rDJYLMgdgsVbZKZAX1bNV2Ks7BhFfDV6s5
hxv3s3Ica1igGFU7GJDtU7Kr+G1qnjJCdPstoeoGgMkZcBaxlxN4OzrnugOeF50Q
ce0MadHUkwCI43tbrHTdGSpoV7OVfLwTuF/JXWoMoG4Lswedbx69aPr8Jr9+nT4e
ZgCnF/EogFlxtGKCuJKd1/YP8mfp3LIU0BfVwrTI9F6mj+cjFgbUq2Y1cRmfRbC/
yBsMF3gqiJgoyFf3Ib8yRKdS/nSQVsmQI2NM5s1B3zF2qa2mNxowFCgfV3hQuA2h
EaGuJZeTcQefXwLfUQBoewaIr+dBodJxss1Qwq8220GHFJXx0QH1lcg8uCIdPIzu
1P5rWt3dvx3KL8mMoLK305ueP73uNW7JpFCcazLcvPwGze4VanWOZaDIjuaiyzvc
EkYo4nOV1OFfd8iH41JbLCXi+gIB2/MawcoGO/pnlYXSV7e1CqJgNnv7qRewPkV9
vZl3jloGZE2l/AK/h3FfgmzK7diOwwp6+UeMnsfvxqXTJgf4+SVB6zO9SVaL00If
kGdoHPOccck7t190h9D1IFETVDyIwhLpBmgFsdQQUiDr6VgAAY6lnSGgSwc2/gQe
ekg5LF+dKAZrtkPpHMHHV6xNN7GGxR3WKMeWw/ms48LaMjUR1RLcMghE83SgbX7a
TUBN1Qf2c5ra3/slS/5cq3dvr2jo/p82jRl6ZqZsX0KOS2d+TpJ1Mp/25WeDDLBy
TCv2sBHNK/zaa9l0cQH/wQuQjaSegEz7J+aJOSIp5+di7ciU+Hu8KXnqD8vAQdR7
JFcJZqRL+LCOgiozJuYHipcz6NiPiM1+2wprnd/qMBqqv+BZbGd2KWuTrwB6iIIm
/fDIWDg9KvPSO5GMdRy9ipyFHBWB8wWCC4isvID1n0IG4Pm7rs2Ak2db4d5kdIYS
r/f2xISvF3epvbQCR06UBo5+wmEkzHR7eMCve455gLznIRqq53aIYq9ghssNaGSN
DhxTyoMIt+q5tQYvnE8R2CYeEOu5BWPu4ipFszQ9gB4cSGixzMfd+bMVSLX1p27i
2A0BdrEDATW58ukfGFZ+xP63Awy0S8kv+RFL2FUQexKeZ0nVg97H7tr+bEmGxiwL
9Jvk3ewpEmgp/jSOyTtpm6iKKzbg7V+bQTmoIZuDGDEVIJOy9XmFMkHinCLbKMAx
0IN8HrVsRcvLSCVCMJr9v+vUg0QnZ6ORWzky77vUGBWULSzQKCelFluuj3LcGHH4
4cviSb80jWoQcS53LNwmNKuTKlUGqQ1ct7nPpmhZFKYUbNSNZXY82K1hKkDg+crt
vcmE7jLKrXxl+UcOmRHPSFMsI7XpT1y5nPdpdqTyH+U2NvAfglCXNM3LwRVGswA+
ScJJo5EXZ5Nin9YAnaRdf1Br2F9NgTsZx08pxhIDQMU6wBYNHr8sXIowuDBmf2Ca
9Bc4P9PTfl38pylCkQIagtKH0HgFNJF8c1kmWD4+Uo0NnSciDaw3YlsaO3tJkp9l
kJuXaDhYPV0bWivzja22V9PbhO8ZMl5KlqDA/miLBFRJBTcDymyAT2H567uuINod
CIS1xhqPNbe0ajv9oHaJsqU7Nk9xb6zkuxw8lZ6WOow4WzIVjDURH02EYmOfBoBo
rdYrT73mJb443+v/6YtNqSpZ9vWYC+fcWTbNaMgPv5zL4Rx5jxI4wSfk6Zg28Uv1
Qr9rlH6Ei0QBZt+maX/W24KwYjC//mA4o9II/JiOr9ZPHJRcd3Aed9B7EH7J3wmS
bQBKM7xuUh0i1+Q1vBC3h0xVZp0o7pftM2syQnlwXqEPmWKdlAe0AN1YVhdFy5ZB
fRvdXYmHFPkfqnoF+cAl+oYpp3xkyvlJr4CaGmiBni7zJgRJFdCX92Nf/BceyeYY
6mIkYAWyryvxkcQ2OFmYip74AaIX0hMuCDEWgHfAh4Q=

`pragma protect end_protected
