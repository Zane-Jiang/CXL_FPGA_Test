// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wCXJaZF8GMpli9HGhH4/58NoEuVvSK+mPiY51jyE5/xdWofvrEtlz8VD519O
5RIqCmZMrdqQnCbVv7aVUheQxI+mslPIc6tJcmDZGxgEKUxoM3jIn7iUSNTK
fJzOCYjqqATUV7CDWVBnOM99JJsDKB/M31aeAbg1nC1mo1hpkC5H9D0CIDli
EoD8683eB8Vac1OoF+dpaUJjofL+vWbv+pMZ0rRCkaOKK6GMUEppPGM0VdaQ
0haiQcWnAFpbBng54T24/42UctF9Ii74Acc7lCeMmz4RAp5WInxiBlp7syhP
pFky3CQolL3UP/bpQuLOM7PVH5hCvYw5N3itScfi2A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RGfiXmqx1GpRBkrJXj3vZyh15KQiD72UqckPr4BaYkROz1KVumR5pogh15ZR
PiNvgmhJ9UDWBOmlCDKlCnT0IHEYvhkVpSTxjo/7zhy0uSZ5Whg2z4AjGRJM
+4Tyd6iENfV1C0AF2ldPQsGXGbH5rPmTxWSvFRTeKiv9tSq/zbyYboQLCokx
Dud7hoIcbIy6WW+Dyq2DGbHK2z3iEjAK1Ywh+FTyz5GtBHEKGBoBDtCswmtd
Tx8NDToREz3sffjzDRfOeXEjwwbGeCaKbjsKOqBvea8qfMTJv/dumOoGqY8G
hb/Pb4nBBYae2HE4+uRc9NUNp58Ux/4rfppSSzxuRg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZMXGuFLdy9vhPeIamW9vZ1NFyN1ghfZq/mwRVFd9IETkljIlRYoktrx5S/3i
Kg8o0Cv69tZLeF7FTvzrFVX4sYSoSZHfH8//QfpqGBca3AEQ/F14J806Gew4
/WXpF8FIA2nyC7uOmrZCiryKfhN8quxHUckftajUChm0/120PavhEYBy/d9T
+UE6Qq4YSh5aHpj+aqdiokievt5ndr09Msuc7LVdY2x5qSv13EJYmvBIRyOh
0zovfkXMZKZvYmuXVCFOZPPdi8SvAmz3WEcLIKTIFiJR4Fme3WuvRawbotr+
V2oK9QUQ+SOD6Z/7eAVTmuLrwjKcv/1h2xOqopQk3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IJJvvBdlbjZbpidWlen/oMCENxi+ddIwzbiC8UwAYXyKfzKTAtJyqhHl2792
38q7/0E4BMa97qo3yS/J4/vgBMu3OTyqfpgJM4JWKrNJTf5etxr9bLuHoK3r
P/9V7ssUqghmrg7hXZX8mYPf1o4W8bnRfkPYx+QVRB7yjeQSf/g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B0V2ZF7vQZY7ibuiqIhbPNu5gvYaXJrDSZ34hycUSbMxFF8pPZ0ItujOLsjE
rOy6oyciW1nuduyRPqFu8Fmn+NPlaUOr65WGA863IqDDlsfncM9Bl0vTEP2u
Sj6Y/7ntnMwQpqS0YLKRtEgloI0mVnYHgIGS0nm2JL/+gKJW3HHBVFaOpybG
8DW8XuJd4AeBYoVz4KpZJ0byV7FgRX4Hl75L0mZuSBGyjgOBk1c857Rf0Vv5
PgTsb4YYa3OhgYd5IO1z7y5imTKnWEzlLUkXrjpeEaNIVNcKRms7KC6e6h4D
vmU9Wm5ie0xrIIYW7KfZ7OPmjAswNsgZpkWu92+qLsJjOcC5tUXAQgo081eT
MD5QSyHBxymhiHasVA0xRhWsL4uvHGbBCrr2/uCctx54Z/9/gLu9+grrlQej
LkZ50rUKYgaT2UBwhom0Lf886GTyzfPBijVY18Y/O8gVvc2E6G7AWD7DPy5/
uZZVulnV/jdsKxrHecYbJlFu1K1iTSU8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JzZNe2M68aZrC2dJbI0hrPMzKQfeiizD0xe1t7rCxhQEf2fjYzyBLbCrvn3r
gpnVqe8BSSs1eJb6Oi6QErC6afvfii64MIeXQpHj/e/JhlJlnMcc49t7W1ke
Jp0bnFcu+m3ETXfPnXDn3yHoMmlq3MxtOZ0orqMHdXw2sPfBlL0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OgYKzhZBZsCE4H5S2dtbZXRpXJuAZgHgIREIf1uFIdguEcvSL/P7hPcNow/N
sgrm2qJ01KxF7o0Dd+7Brwu7MXxC6LAIFd22ElFgNtsIjWqanENeu9/kRp5/
IfASNHdUHWnOmitRM+BxUeIGn2A1MbxIi1kaCRH6jMjlRSCq80s=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
4buAxu7RhuwbKyvS+rJREjrB4H/VTJzPlzK1Wb7Kw3Ivy6faabKPuc+su5QY
OxZi88c+BeZOXm+BZqqrU6AzCFiNjI9AUhCj+gligemD9EYUZ3+mwxPZCnN3
Kju8dQ5Nef7b8sZLNUU187i60rrnULXjic5Jn17stBhylHZYJkw5CL4Mp3ba
FdovjeG1DEWuo2kB/sqT28iGrmZvXJeM0oZlIqKQBxPhrIlSh09F2/4R9jJi
M8eQs8IFoYBD1J3piArbAzIyfmw8LeT5/fCUQfKBOjcwWX5HBuTz93wkcr5f
dLVldEtUm06O8Wf1KZ66BFomVm0mh14CqOCWKJeci9nji0pGGOrQuYU8pSmQ
9Vx3QKQtyk3ibFv5e8iBaSDui39zZQq7oS+s8nZQwb0e9l1zzv/w5DVOPnXF
bgYkPjlylaEwpU1Tn23ogMAYRJld9m4jy1u+ck+xKxd/NWRr8ldtvkcCBUx5
pMJC2ZaLoHWZeq6j2xFEzy7I48lShNGXI8OOCO19pAno4kCCzpwNABfT6SMe
61yReJDJnMpTenuOnHuxeL/efTwShzj2SKkZyVjGBrOR7woKJruilbYICvZx
9PfKSA4Ip4OdFoxGaNGU16IJu7vQYejRP7d/TDj5gRdu9qlyX9sH7NypSzou
Cdjys3ix9P696RYvUrxaSHLWLrIanUOTCdPahL80uXfjVgoTb0WeUGio7TSK
0KQLviYab432n1ApzUwaauaJBZbxLfGJ9XumNTubU2MKVsaw2Jm3ciWJ5/RF
ROxQfQgMF4nc0cy6AD/eC6MPwgqutgPj1p2AE5WTyjImHmYuH2SP9zt5QYti
OkLylNwycS7XQ/CEWGJGqsHYmDjdyEBOZvWPEM6pVEttXbwvXlYaO2p8CIdV
yCgFngc7P0VXYKY1uUNh6ddHTmzxr7284ueWwOfbCRXSfVndQ7mNdgHKri/z
+FhIFDF09EkHXt7KZjqVj4WTxtcNP8d2f3zrmJs/ifOaShlTPnsCnyQjaSWH
PatygTTifh79Qt6wq8Rih2V+5iH9NkJciV25yMcmmHaujLYazcLC+kSP0a+S
j8v+wh+qBBlYBJTeBS1E2f+a0VFNrFebbSn99iRtxYxXLgxM6KeDGtrzgbdo
KhQWY51jX9fvp31CC/E8dp//D0H1JWWVjouIjF23Mr+c/zE6v5wkj4DMgXwR
HugsEBbMZK9cXfifuaZknNupFH86lXDV4J7NnNQkex6iss9KloiPgM/BI70m
wqIgJttpjkxd/NWCWaMPlkydyMXwmViKPFmU8n90sRxWFbz2AxPuyxkIwIU0
BVUkxdE/lnE62L+dF4c6dPfVBGSGzj9TVCsIkR3tvLFoJZVYdu+KqQ2zgcrs
ueDR2pv19tSV/KPl5xxVrOo1HAQYboLc2+ekG4VNjsb3e3M+E8G3/zjEU/YP
lrF8tcAebAjKoPQN04qxuZKC3QW27pqxMALHGus4ppuRYq/laHHFgOPngQux
m6s+Ggq+oSbOZ/ZgE1lH6lHnS67a1K85aveivtj4bLANhgYLrAgp5y1rVlvg
525lR6sfOku4ViuJY79kP6Ra+nbeb/BseRVOUR1h24febaeY+1ngkQ6KuxTy
fWu9ZTJ2PhlUq/CsoIO6OKxROUR9uF+FdyTiLwy6AK9KDPQ07T0FBlft4AQH
xFwG9cusCHdHuxMJUYMDWGMljwg=

`pragma protect end_protected
