`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
FpyiqOmoLwkZoye+ibRIylM6SGDHmlrHaT61+jTpkh4eqJuuYe3VfGZIfEkqBvwG
gFjFPRhPZUhhkxuAMjZ13GAwIKGtthH0aguTHR203BEAIpPh5IwtDmWKb61i5+Yk
9E0DbXr+m/LbUPGIszehcv9hxKbqnTX7zAs9dUzie1Y=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 46432), data_block
v9gch0xV2awTwArpaaaTj+R9uqumeO6egsLrwsoknTpYwmcjaUtfaXQr4sCKMtXv
TskbV0Ewsuu3ZF+BY16hurjUjbLt1pgNhW6P9MnXkT89NJk9XYiOdBsQEn9vMJ8v
DITQrT7+Evcm/8duNXqLy3PsuIRCMRvUXlWoDP1OnBmII9iBj50I0aAJ03/Zyldd
r6jkth+z7xzHiJOyItNGl94iLWuWi3G2xWRvUE+PmmTpWPUVO1bVZgXwtarejCY5
dA0FtRiHcBnOONrMIchYcWXwiAAIYXoUm8bMuAAwXkLh+MGqSFwflDuhKHSP0EQj
EF2MkdwKlpOee+y3zo2EsZbgXcmz24WMwBQxL/VJ0ygsovH3LLFEqgNaZSAFScqX
UG6tlnSUihQnwN2KwN1Zeg4YQT8eRcExVoZL4HtmBowfowqNJs53CtFe+aPsnGJ2
hM4c9zBQFiItHHbCnWIYwTjCNFXCBjltUCZbYFtlnF/17ucpHkyhwSqb70OQpZzj
b7ssDn+AcXHczL3g+U/Io/fdvu9m6QEhrpqiwCzZnlCDeuZ+dmVt+J9cR4TcyiU+
WBBNreAUD5Wbe25x2pU2zBgBpAKL3cvBtxhebw65iBHOMG0nl79w1rF54NifT47n
NMOwawO4Vrl8znbvJwauzfZlFuGq9LC0MYU9HGmW+oWbxvdvEn73J02fbWoJdQfA
pRdz4c2K5bgI7gDw/rhVk3+x80s1UV9KpcZ5zGgU3r5e/EVFiE92Em90qC9JZU+t
hQ/BxqtuPIx5yUf/zwDj3PeQ72SKtX/O/LIsaJrvYoVbWq4mQq4rKRqWQ+CfEgpJ
pPv8lMB2B3Hf2yrOU4BagJqEwINZgTLcl3C+bZVoVG3DKIqVSxd1bvMxKVSZxO3b
XcsOrNdfh8SXb33k9KGijOWTEkNMSG8/crqeBxBDRVOMIBEk7OR4xD2x8OKny2xc
fWXxgdUDyZHgMU6D5KbAx4/ZwTDJ/jD9/0Th4N1BZURJrGPlqM9jKT0QImr6+4LM
Esk/JxyW3XRWTZvpM4Y7UmFqNoKt2BkqeSCW/p+/N/icyOqSkuW7jNBat/sQ2FXe
sA6ZmTeGqLQr+JnbbMeYkFoxxBSaG8EwTVca8C6m847WUwdsEcoOL0JY/fzBBMoW
fhc0yKOqYRBqVix3WCnHqXS3D98lR4wJqVhRwTSasoNPo0mpYcn/skngtoX9X0Cx
QSkK0BxPc/r+4WgJwfi7gL1e5yfhdx6zhTRVEwUDdwVEzOBuPel8vkNQhOgLv6WX
0jhKsS53YlXAXY6hVGVy0cBCN77FfpidhqgHD3fKKWjb0IwqQ5HoG74g0wufltT3
yF5QI0fwQYOFt/xEuvqWYMaQtMb+E/opPnax6sfTgip6T4z5p3+GuQYsXEjvzRFi
A/bDI6gZagwy3Hbqk66qqv723l9kjdl613f22MpARxFI2Y6bbjk1Uh/RThI9x2q+
QyKtSrYLth+0RYg7i4jDeHp9+gERbkCF4nsVdzd90F4PkVqqmTicw0l0Y1p+N3RU
ynBY77BJlrij9BWP/C8mNZd5hHHZkcAgba7kbZR/Ef5eOhNQaUrhSRJcTp8fkgFr
4hB19vp9fX5aRLgmdvdXPDc+h/iuCHXgoexMc6p80SqB3XhPZ4pe39Ca5Ly+OrA2
5vOUQ0SFScbbiuqkPXuHceKI4UhNhusHO3f5MQHUNkxOElK8vwQ6foJ7BKtfGKzV
hCvX04DlUcDSqyv6PU4/IhGzGgGLOFD+9qd0lvMNJ9qn/KpO78hQRwnp3O2cNgqp
jW4ag0n7cjhUcTypFP9sTvzNKGb/6BpwxH4FrGlcKP+Wzw/bqOZ1wkaDqW49lHyu
mwnXGNi+3qtkc5DW/PKrVi0NLlSnP1RmbeYQMtDXumeVwyFt8oaMMVGB5LS+xBtN
3GlLwzG61Qs9OwndokJZYyXxvK+a07f53zCVYHVdZ2LmuO5e2rVeMJbvgt+cFv0z
0sv1isdY9Y1PNTN6PQFuKXVkzyQfECO7J+yukcoKf7HjMArvOi4g1j56rYpD71kO
WeqC9s4DtbPzJ4AslDo8YIsR4UE3tCwiNTdcd6jJ+KYqESOegOJeDlR/fVrAwIO8
Sjzo1MYiN72jxxlhAsq0UTep7jT3QoXrrXxk/en4lzp8CTHzsSprVLAzxk8uFJuF
M8yOXmgRbf24S1/XYpuZ3lw8pQgz3sSfpvM/23oZzYCJ2xg0UT35nGxRhs9KOfnr
2ppALX0iqdn9OKM3Dj9cYRc+eNxGmny8m+r4HH9Qw5uxuXMHbZd5pvY/bMz3htfQ
ITRkkGGaOI9/+disAFZaosqn7IskzZgM78nwG0Rjv8+2zMVBaApkfUZCj+d+QmZF
R4CAv0aaUV/BPDOeDLqm3uMx+y9edwsIZo/ITYBYGwXRgBoXPgk2FWq4yeB8GyUF
iOeHFJWyxvPLaXL3AyGgxK2oXOclt8t717G2ubCCmHH9dgv6z0nftJauONx+dibn
nCwyHemxNUy2+WFQsPtppGhe3se251F9AcdVi5/Jplv3VUbGKQqvQxpu7CVznBTb
GzYl+U+lvp+kxGFrhaE/unrVT1PNVjKJI8HuzOWw4sA8BtRpNHdvDABvZljOBzov
BfdYogcF8HmcqyaKKx55SbF71mXa9jOrS/hbJqg09p5Sss0/5mfcz3jtiA+qLuIZ
GIpRcit1ASuy4Z9K6f+hRb7aNqEBY0dIBd8uae3xNHrq8f6Fn5HKyOI3UFFi4w6y
CSXluOqVy9u2mVvRl5pq1G8dKDKFoWBLwPuWwEUy+lVDXxeoIrIeUcTRLV8OABTH
+fnmmadEbRhsPHCksLsjEADdbCAESaiUP5K2PGq8ViIIddTxyAGrdmj3kE3buS4d
XC+/WrQ5FZ3gvN9quzzQjLW7oARI9l2ilokBUIDZNxyUjDE8CjweEZ9itoeQjHdm
FhHtvDrrDfjcoedu5XFqe3TS1wA1+Xswvo6yDA5XF5TVc1LZXArxx6tc+NvhsY+b
JZOFdr+JYB/R8H5JGkB873adk+G7pxweuQBYBDpcJ27bkw27sAWG4FNKkSqUrh5Q
6xM1u9NyepDFhaKsGGixIAu43+jms+PhToYC17rVnhyDqE1RKC/tDQAGujk289CW
usPsDcu9Lddcd7LeDaOjrz6S07vd4JfMFx93+s2OIaUWhTS+pvGf/Vi36KmWjnxO
jvY2PE1RxqwmQKWt3+TztlLAM1bFMD74GX4gqd6n+fbeGz2Xj+MoYpVGPjk26gNm
j3T5FV3NQOdvCKx2p65ci/TSfoRiDkSpuojeZr5ZiEsI5pZt6G4q0mum32MMy4Pp
mN1eD3qp5iDDqAa4SyPyEYVQJk9Fg5Zvozmi2VhE3Wl0Ac0ybEDQvb3uWm0ZPnl9
tWrRNpIoHs0tUupHkwl5uISF2t+5RGQoGjR6aogdd/gG8Z1xk3kCYLM85KzSTYPC
BFi9Ue/D/H/sF4fx4xAJ8dCj8gLk9480aw+qqZo7gDzPyUIF68lRuYckhP1oH5Tp
uDB1kVP8/cPDrHrE6qdUqdU53ZJTwkSsLsSohC0a+cFovH4QvQesQi2QMsHmwnDB
j3VswFeJZY+42amnstma5+cKU1+Zr/XC1NlOpEBSCZPUXieqHcogjFStCdu7xYYe
eVH3RiIO3BxktiLm6wWkdasha1YUvOFrm1vlVMXpjVuMJqg1F8lGlzawr6AuNEzM
TfPk9iRYi6eewlo3Immv61GpsT1q29F5wE9BSh3PdEBwnby9BQ5gcyfexZ7FJK48
s8MAPF2DxFwvo/ZQiPUsBWAr8Kh1cvnerNC5p8ROeQXPbiRjbzI4m59gF+kdmucL
yG/ctelvhigcjWbY6wgqQ7YJepLnjn6v9Ji4AvT4f2UmG2bEDtT7eqvUns3J4Jo0
8jAs8eqIXhICcm+ikv0Kbm0Y59aVfWbclZbjdxfn1FXhnp/d3c14tzC9e9bloInk
47OoSecMuxNwe4nIkoZ6Vaz718mDFthOwaTVzelzDc56az08lr6XbicHl4r/ZvH2
c7yemqUUGfZs2DLHDDRCBR95QrUr5ifCILncSzRoLDPyhTp+YrCY9a3ACLJkm35D
iMSrMrT+ecImzrsInQuD52mjNRxHYCzMkylu7tLkiWd7ffUUtHgCl5QVhF4yoLjZ
seZiqhjFy1xRf3smU2m7qj2Pnl8Ziom0PWS/8KjPQ3xw4P/9Hh606kmPheCzJygr
J6PRngaqlXCEeVPgM9h4Y3jUTvPwchBawOjhP34WsifZ8IdtS0XOlyLDLxJB+4in
5sQ6gziYq9/gUvmWRcaKWx1CiAQmpTY02lEO3X5MtMWM+gjxKPkqRfLr617JLHJI
v8oJ1QdLBLccHtd64Fgaox6L2wNOY2n7JZPj2ZrQIaEc0Lfd3/VMwyJQTQM9+iRH
KhjLVzjCwtx3/XyDHv2ynQa8HayNDV/Nn//xhTWV0yr3lOWFlwsCN0xQ+MUfdD5K
a8GMiiWasUhRXSoGRS5SAEsUJa3mRw8AjEkLfI7CPrOg4OAyBXPqX01jCrTOuX74
WvF+JFvWEMISEb4h57rrlBZAz77w+bPaDZsqldx+m/+b+qVcoNORzkF2niOWIVGn
JlWAAdgFfGqeexzfY9mjdPHW/Zbg/YNzmrVca8UcG1ILbOh/Ss5MRPkNe3BATnZ6
px//pZjJdu8itsm4Tn/jOv1bywZLSvdvumpzu7D2zc/ec7Yr8cYzLxMTvhE4ES15
PwvZEPouK3DlhlgA/S7nekkBaSoQhUAowrY8cciD38IkqKJdmjEivkYmJS1wcKFS
DWFHHPPwFv+jksSbi7MX3aNouqb15tI+pF0q7SU1foYrwWgjAF1L1w/kMJyifjKa
APQblH85LYsHUyNmTrYNMAMmVYKxnQClIlIhhg4dJfkOqsSNrpDyW8Ke+SwOj74m
TLttkltEwyrlbc4tJ4DHUDKwwq7vBHI+kCXDk5cQcQkarnyv594iOlQwiqFCPZ2m
lado+PBbqwxUlIEaBaEV09tHPEtK6cQo/Ad57Qt/FvHtNrQRypVti0DSAtZmf1U8
/qO10hoAgCR8VELxKV/JKXBxudJYUrcR6tV5v+w0F1amq1CN1Yi5LVgeWQ41kCC1
OCBFRQEXSLsy8MA6temiRGeC1Icah5NlW82emBhMeF5D2mhFt1+TClGPVocDzGq7
vv7kHh0004GhB4kddfpu10pMR6f8uQbz1dj3LtLnOBxD0StQEo3QMC1Zqz4DKTjv
cmFibGvAGxrW2Gf00fKn2qrgj8GS7sUpAsvCUa0M7pE6OQtASOGI2CqPlZHUiiIW
hfz9RYyQ3gF2lu/CWM1dFkXdSnh2r9674XAWNgvzdLfKWT9hkPY7UFE9RedUAVTu
qiLX+DIeISwOFhF/GeIkP8lBqiNGAhnsQC0/JtMdp3dXDXzIhRg00Gz5f6vcPnXK
4+wBTjvV2vrV6V+R3FHSsL1OkRAX4YvdVqKRK7fDoP5qgyGshkYSyb0XU1DndmrM
4fbkmZXTQHqJFXs6EIlIC1z2piJgMeEO1xdQpkhIdA/hV1wqPk7Udl2eM/ARth0Z
d6FPgEpcglFjY0RAkbGc8dVaz94P2KUQUZt/0tl4zjpAUDvJUc7A9CuVi1IdwR7s
9/M7WldziG4gEeJx3XV4h+Hlhkf+cfTK3NiCcjgvdDWkmzQ/kQOhsSfT5ARIjkvq
Lj/87qMcOFceob/4S2U0fAtLPknm041Y0JtwdD2lwEDhBeSqDur1jq8Urms2v9r7
x+Ly/87U6eWck0KEBSRJEagYxaEsBNh8KcaUbMedgMtgk6bEfQHtpscHOGrt7cP1
PTNoDVfO/ypIqgSXCtg/zgGQjp3caRzAP8MI/QAfhP/YmDH6H0BkHKtGqhBZ09H9
65KYOVshUoITGWGBPHag/skWn+E6S8yyNlvQQdRXgF2X63Bd/a24zDUwEarM+R6J
gEHF097bWNrlKWoO8CGC28LD5PFrrIMrRDjxJXJUY2cD9x3M+fF8N/hxJ/Tk7Yum
Ofcv7KZYIOllTxDH6T7RrGHk80OMZruiDF/JgJ5AR+0YjGggp2boOC/IvXkCrroA
im0mcScP2XYgH4HSvHaemCVNOj9lloQsRJ5Kuur8whcxVNDXym93Pk8rm9uGCAk8
aifh2GgBuQuu8/aCw2q/nqnBFu4TvHXBd7l8SfN6AlpwFB8sDZJ4B2nJYGljnl6K
y5qTidugbdTVOwphroX5hmHCo4SMC03Y28/oVja4ejnI3KUxDtm+PrLdyoW1Pyir
QmVbxnJk35sC3O0Cmn5Dp0iUhIX9cgGpGmEDToagzc08DfwgDK5s/BHZTSJRFQXp
crtbvV41KLyI8VkSHJSiXW+NhBxCl74k6zAwDnHPrzEWpd1XGjxRmFdSfPetG2/V
0pF5T5UdYZxV8wu/e80dqptLg/bq+nSEB7tIXuXsWOeAhWnqBwWpCum6oQrGRcqo
56B+3uc2l/Lff8Hn5M2ZJ1geiFFHcFltOGXeNG5e7T8uVyJHNXXJCSr3cbCh+NGu
Ggxut1LmdpCLHd72ZVcDajdOpTtFP+ezSg8WIspDLj82q1h4cRek0oehzoGJhV91
VpLpaLtT+8r15YqFHgu1msH+0ymGOA32qWpAPttzRwuCa5iweSMBzfbe3mGy7vTG
InhshDDyVpalGCM/20v/hvTS6j/oAR5Rp920aTSnoMA5M45wPXsGurFHxiwfoq4u
xwsqY56az2qI1XuL5H9uSGP8q4gmOD8vWMC1xjXXDTSQTS2z89W/kNBbI9cGqDSG
aFL+OlbXf484eLxxEjLnHF40Z4/YMWlluuQgNSQN4sW0SDQPAwXfV48QSOI+XcK9
D5Cs4dNXHIzsvh1TedBfWRvadWlYGmz/M8rnHDyM7iKNgRaUy/7UElgeR+k40Glm
GUN+M48QhImbjxFbqviPhVTTAK/RmD5RpBp0kpT29QfXtXGT87Rhppy6yWeSkFEJ
aeYd9hR8zS3eQCvCky3jpntTrbjEZGTPNqn8cFRTYNID1BMAs1u2aw0hkMateFiG
XI+SHNfMaURrHHhfDU3bfVQVChy0IJdQEBFzLJVLBK8xfYjJ0OE8Zfi03xztivLv
WYvU1Fz+Y4BQCJBwghg5NjLDSSsNF0zAwN+8JjlSJm0pxaHXPDWXLZgbe3gCeAfL
UpunG3+wF995Lj6uRlwH8IuR1yTxtZ8bae3y1gTynE3yX4xmB+aV1dkiodiQNMdl
ptbFpzPddUy/wzubyEzE12/y12bn+jDtNAEbmm9eCLm/BIkTPkJVbux+qDXtOK8T
Rmj1CZKEK0X+fCQuj41lEi/DUr+JugcRMbHWSlf8Q9gOdnUYqTHXGf5JO6gbfHQd
3Eub/bEtiM6xermXmM3HeaHfV9fWXO6pBgSe3qE8aRc86O/RHOG+vBN6N3db/fjY
0Ce8jMckRdJgFddILCOVMMdBg0HF4po6LgbEbiG5VvuwGPVK1FtBDZevPD1VRjsm
2wFIi/cf3gS3U/mIUDq3zohnfH62DLT9ybbLvd6eXRlWYSygHoSueTVkIaqLHRpM
9Th71LWXvZlBVf6xdVisFQFZl9B8u7Pn6Z/Tpt5lmZGd2GuCzJBGMtlo+YPipUwZ
ygwh/c0sajlF4/ZBNo+BLApmc1sVHBa0a/1WQ7K0s/Mid40KfEFxNa2F0ylLCF0u
ZupwlTLJz0GkophuR+Ur5NheBPearyJHKqFUzeSTx3h/rPXhhPpYJVOjB02pyIkv
ej65HuXgFB7fDAuH6zFXs8+nwJS75gvZH4GSE8qhCp1akzZVRtCucjSbYtMFVWGI
pn2gc+xN6sMp+9VOdllcFtnn2MgyXBBln1Eu4WsxSjpcRlm6JFIYFAa8fQZAaZmZ
EO02MWQurRb5VLpu2iIBRMRspq5KlxlhsziQ6GcJEjIm039OZRC9kixwibdlvQ3R
4Ho7z3P7Ah6+V/p/8zPV6M6cFPY4ojufGT90Xx/X6TmnWhXolZ1XtgJLrpOx0ltp
SaFuQ1QtRBc8aG7bu8o7z1sauz7toqSgqAEXR8GXSHIYprpaPoXm0cppY5tL75/c
Iov8cVaXLJOZOSzwEOIlMWK6ecLZrUWYcQlzu7DHPB4x3s/Q8/6yh+5zkvOlAXeI
kCqpo2Zj6y2mcJvZh3GnYUwuvp6/y1FJuJzuAylR4WDc2KPNaSQSit+9Bw24lGXP
23N7ynEmC0x3qqLWfTE4neVOdWlr2gk0DmEFquDYBw9uTpTCSZs0u5Shs/mMiKCB
bFcukLfzvmLYjbnqZ3ZdFd6k0Qb9XsEIwewh9QB+Z2AXOP85GAEeUjsUore1+pyH
JLMH5G9YKgf+zwaQxuM80bzL+ruXc47KMhiIGLP1JHMJlsvF6/pjAVQgVxJxTWg8
ZZgGtUT4MkzvrdelrQJSqdN+vvp1WHH8kLT++QBSpL5anA51VKGwgzRG/ozh/N+U
CpMOR/U5AWZo9sKhNxC+dUhD1Ms1kwYJo90ryZJDT057EIjciBcnWNay8PsDNUWm
SbgIXRbZ8U9FjeKbEYI6a4hraV7aopnxmJN7aoj1HqU11viTX8mtD5kInqWXHuG4
N0YE0SPl5LemqiXWX2VAVrcLAkqAbI34VshxWRTE43w6+XwYprgtnT1/BJ8UhgjJ
huWTAoiP/1wwneLpfVSzikL75bsLTcZILe8ZwsVunW19J/TfH+n+nEcAN74PNZr3
D31BTkHq01qmSu9iVNCWTNrjDILJiBOryT2i9wL8bImFkZHBC2XGXpn/0YsLgrq3
xW71bVyyzJSj+3TmqbxpWV2+lSqZbkasBSvZgX+xP5HmVlBzRSdjfPDPmZdzMPxo
Y9+MuCzrftRVy3HahCgp1DmVKppctUNKR5fRm1RA8tSOqByFtgEfEx0m/6+2VBgd
xNEpk5tvEGJti+On9VCP8Ee9IhU944G+9jcPfl9hBSdUXEGv9ExajEpBXk6Y+IxX
maxg9oxViuHxYreYNbei6Lu/mWtaCxTSUhQP0I4P3gGqHa8Cj2ymwLTGcq7wwmFo
lDrKQZ0udfdaPgSuABqXFs6JrHW5skOdQ4PV3DOnSsM6LFz72SSNFuSSVF3IJ7O3
/mJya+Exqr4Ja5razf8vAtpy0WoFfFNvc/KDs9XnRPoiaL1PD22Pfg9rUzzog7bx
yw4QbGEtRTcHX5kdccm4hcEXM0Fa6dfefteVpAryqwfc7nO1CkfjfQYr1+CFtVON
ddPcaoj1RAlLY1Gybdw7o9TxpONtQYXXv/9nP9DMGYzDQ9B8slKoFDiuEv3qRY8o
CWNbFyXYejADP3TA7zrEs6n/N7FevlRMxosum3xsc/L+dtCWLLFtaKYHWo9c2srV
XY5P06X4LbnWdi/7TvJ3jWYkD2OeTHxfkE3SZ8A/0w7aF6vQCB23hy3pakfDY+Mp
/j3HqDGuXI8+H5V3nD6TSlYJ81ZxO47xxJrJ51qO7ZsYAo+5/gZTQbc6bnlNVX2a
k/k/R7TWDAHrZTnHEi6OaBd4QGIT3h/d6rqYX5L3VJ2hG4ztAI9KtaR6lPFq/E/z
0HMun9idvGPGKQ2d+bgnem20ZSG2ggOpVtEeIzcI2dx42YqniJMmPs35kxarCbT0
sDev0Epta0XZ0cK/TlNlqXou9dewy0XMWDpHCuSiXYyMJbVTL/7tHEXrL7BCbKJM
zXD7B6nldP6C+GdxZiglGJXzuR3Jt71n2yb6dhjkQyDJXNc730A+zdLARZga4FrQ
nloEl7rUxTOKYQey5QSXYAZj2BaeCwmzqCTpPJn7R1fP2v4Iz5QowE67PfWtp+s5
Fg7SkIOmqh5AdNADfAa/5CCu5N9xkgw5BjuFdqyK55cHgwPK1AWTmYwTBr/6XnJ6
vHOXEwUdB2XANUz4KMz1bE0Wq3LGlpb89bilgCVufAnEL0Mcv8ZRAwj+b7sRcjxP
+3/r9mz2ZcRQMq1mbAXSSgEOh3pQ9iI8Rg1y1nH/tO2j9z2ZeB4t5a1Xpca5OzSG
XClRj54UsAT8Rdm7g6WhsOXNEGP8JNQFe+jOXtXsJi4CFYGMlXBbS430mNANMM1F
m5xyeHur7wKKwyNYwnlWASNY9uWzVrLqvyvaXuscUjPnVRM/zwWWrS4jOFx5rllQ
se2qLp3p9NR3QdKbEc/z95EqoqArQCuOky0meOLT7d+UdMY4jAPn68sDJpHuPn9N
pHo8nnOqLFTbV3Xt58ptpNK11d2IUXrsTUcx3QigeOFTvVq6JgmOEqmzkIOFvEFQ
cjTgozqKkMw4EIlyOpUncthsIipam1j2IWQomxZSMA7K2e2OlbjQYb3kUfmIdJLY
doiSWgkgVBGM4MawVYa6STRe/4MZkDvydsp7CFKJlX6ssi/LiLr2+STmHZ6cMZfY
XRrAoZ3bI/xf46bGzlpKImJAr2TDUftKlO0y6NQ2No25P2xfYJUx9IUTi+KKEQRu
Tr9uMBamlDljtGIaW9tIEOloyF157Jpmp36/KwahkuOQwj5JVudoxLrRQjW/0mJP
+HT33JdgNHcTnaYObDgFDiDR0DuF0EjZjsy4U3ksyopdTx75H2hPVZxpIWY3sfTO
vDf19td0HeULsxlqytsQwu9pnRV4NsBX1OsKzRaMcgaXMb32VdMvhHoyup4QlfCh
rB8e/RtbwXFYPQvwqnVWtMONnjduXjuWI78qzqkN9OX2Cpj9h6OFFjmHX7VGn1uI
hgKoViVts5ge6O0z+eF9zh2o+jNgkK+JLBDnwydJ0oQ9swV1HooDDht+IkAtr3kG
uVp4l2/TpoboLP2zZ/4mW7e5mmagr67Ukh8UUR/eb3ZrN10BmRXNImHrF/sp+KDS
zAmo+iENAyrDBHHBXir6pNcwHhP3f6GS8Y9o7RFFxsIiT5v1Zb9xxQxN8MrAv1Rz
y7ipeUnBnOS1/SOjB72JKfRwjdm4xXPw9P/6DH9RkQ7/bgkf8+RIwdTnRguZWacK
KXqrtCXZWDbBH0R47MGzuF+GjAI87mdXmhtQrbMcg9BfRsxUaZd5u2hBO4xHKljS
CXLQCdgyl7AIrfP3acZn8SXenjtHupVJHp+HD+cidTppl4lgxjX3sALjxirUC7Np
fzbIvFRrMEpQRUODLrMPy5OHtdvcwanS9O6YNmyLRa5BUc0pRQxFY5RYMXLHrn9t
ZvrQVL0kZLfBvNCXdgKsG1mXRbGmOG1/lBU/oJcBGFFxHq0LOEkDR+xM4aZArLP0
9em02DseENXbCQ1MaEUX9xFiPz9o+TrbzbQpZ+fXK9HJ3KHkMywq+wbcyGluRVqm
yQdlCX8WdqQWFpotHaZoSSfen6Qk3y5iGASroJEoP6QQTvJwbKL8XJfgkOgVbWNz
eWBzX3rWAYgukHXUjNxZ/LyXffwjlOL3nKJZukWG3wUzF1Dcg04IShT3B+gC+kVN
6KJld+kKf/hc3DpUL+p5mmUUkd8c8lJU+8cZcx0Y7umIWr2jwt2MyW83Gw9mG8Py
0Vibo74FvRLC9N3arXk0hNlnDdqjc4sik2+I+DT5pBEMruybGmmeE1af9A79/raf
9rARDOw7gGZsQI5S00DvsJlimUMHr+eUX3Q0LXHAIdQ1zwBxBAXnTQkpLrng4Npl
pyaRK++58Wm0yyJ0c5vvljBV4EsUVMI37cn2+PiIYaRY6fyTytKCZ+dNODbogD6v
EwALTFZheMbsC+rnAIFK8o80MFUCcjJukanT6Eszlg6uHrl8Jq4P0qHoAEHeLpKD
dndRMUgTWNmzOELWrGrGyYSPwmX6cJEiGve6N9Bk4AeaHW6MLAJlxTDYFast8TFP
Wz7sv27Xre8dJbcsHWvYd4lXvbYjTnloa50DRP1DpObC/9NZMGuBkSqZ5k1ZQ1js
IzW8qTTnLuM7h7h6yFu4zi3Xf+BW3YfwTxakoRTUrTtfIRG4fp6iB1gJm7TFFHz0
hruKJG1TP6ehBK93eVVggJPauIh7QcWxWu/5MnqLeE84cvvHhHp/LKrlNdjsweIq
FtQfddAcMpBPhcFwSPExLw3Xs+bzl68+rNW/lQr6qWjOZyzfXUoqBYZShw7XESWW
MvNtlJm5wAxboXvUBiJ9exHdBNvTIgWRqgWOg3FZ1+/2+ga0g5fPQu4VTKALdRMU
0TaMMq/TyfXyKS0MWGWuFRSEr+4zTV6PFfzFMjX7F3kMYAWRIog2NXT9pn5jiXNs
DnTwyZFzgMeE2Dwm0/WHE18r6UXAYbrYblfd9ammYEAa54Ar8l02fQUTFVLSYcXo
4QSf24KWXYgKsAuFuveupjqpEWmsN6e8b7cRpJAo8SGnyuTwpwfHKuedCwThtsc8
q/BXQz1non3VfTpF/6OSR2ORCfmjl4ES7P9LPXcewyg7UvTwL5Ot+u8wVBPIeQ7d
PaLYF/BoeD1Kj7+gLR4oREJmqS+zRQ1r7YDxLBxGC+cx53sEjldmL4hsBY0KXgrL
w6GO14vog8V/7kN+lPqHPIGmQISHSmTbiSpIGmkZJaN+vA6xLM7DqdU2uYBVv2KV
X7sfX1OWrymOU1JkNrOgJCrlFUIckDqMBkD1ldPAYhnw1ezxwSQbhqqtq87ggKO+
7Df9nbe7iqFN8fiYmViltEvynHp62Y1ekgU0ocGIoJ3AJ/SxPnnPB0a9xKu61gI0
BAPYfnloQ3vOJj1ygj0ZFoRIbNuU2+9qCPEa3GKp4unX8LIHCsG3UVnAglfbXS5m
2Vmd9B0+yU2xjXaCfhj+X4CuFaaRcCirxbh0/hoqE1IMXy4CkMgs5/GU3QNeYNlU
GeOT1Dbj0QvP3E3ZWH8EDXgxaF8jq5lmf7Z2HlnrntqUXA1TKRQqNSdieh0M8V/P
9cAMWUjx53xAG01LQgIz5RoryrAKCcnE958qdtU/RLN2hqihpXUgR1NFv34lE7hA
CkUcS7l4S485vWRdomHCELDtn1TGkEexMWz2C3UeRO8jTHcF/Lxbm6jlaZnEL3yw
rizmLNpnAMXPUL8ybg4g2BXe5lzHsIEbxSdRx44yClUcQrtz6FY9DFwKC+wToZJc
CEfA+pJTrncO7OtCpAbOzi4bIS4n9BA015SSP9DvUw7764mHT13PVZ8fAs+4yTKt
x52Uy80AoFb7p/EGd+s74h3D3GVehQ4nrvTRVTdTnqedLBnV6wro0NldXyv9a3s0
TRo+w34Xye0nVPh/RAGmoFfPU/brO5xk/1hwixkn+Mqh8NjxrOTqGf8Ghs1gDXfy
+gBK6wYjqpG0dMSQzqddmn3jR/nW9NQ2ewHYb4mnptNp1AmR/4rXMUQQcXBiRCTE
0BcwBXFEQxVZMTqJqdZaKTwYb9PrEhDRIfsXUfGZfvDMlR3S/Qca0o+QaEYxt8xs
Wy5iyRcg+Eo9tAMrVoHgN3pGASCzah/L11WtNRozfvW3+ZRtfW6+3LgrnUL1I1ZN
wV0BJvb7uCphrSUvkwiisgzc7zm385wipuHB0qnhtvgfCTH8Ksd7wG4FbHt7RNFW
v+l4OHSBPSQWiQUSBV5wTyLlz7sqq7X8x9HSK0AI4Yvz12U8+b3SwTx3JkpV+BcM
OHZIZ86koRKncwFhpxMVjY6bd7LyVD5ALaLZH63V9Oed0KLMrGW9K8C9vzfxHlK6
D8pjwUBnE3R3lsUwEHfxYPTqqMxR1f52i7bjgR6AvZf0PkFju7lhKur1RXAH2DVq
uQa5vYZcZByBUoHeZGTJYESZ5J6lPsJimWudwBMFx7k/9Y5+SPfjCTJTqqhAU/dG
jCAUaCbZsZwQMyJIFDsDdTOR5trvUxRZuCV8WbWC63prbcjh3JUu02r5FLUtaAvQ
I3IVauT3Xz/1z5hNXjFA9hOybh4g/ToOcFrbD6i7QFX72ZdCF7yT23pKAFnNHzg7
9RIVUygNsdyOw00VZy5hXpbmzJMSi8mpA7nuUIb+vaalTVwbC5PXNUG+7qP0Z/XV
j2KVce5xMS+Efly9rzUwkMQc2mdsMq77jQpHVPbF8MscquxzG3UnmF7jnI+bBE7x
0F8IrUavWhHXhi13Ny5uM9/4nQ2nsxgwQSacTtIeyWodp+qbrJuV+AeXYOynltdb
mYcI3hRX+ZcQZ/rTXigm36sGeplWORpQyxtS2P2VUGDvB2ZnLoXY928t24dNvjpz
ujwqJUvZEHDY61ilnR2YDfF1Qwm/1udctmjXw+VGSzyPLHqfA03Erk82xLvAZ5hV
GT3uV+jm5hEhjYbNH1k7lDvj+dam3nRbzT5eDVqSFGxBKLigu4P9qCh2fMFcx2W8
rUvH8O1lth3BNUrcCc2+YUEesmBzEQ3tIsvF7T677k1HpGQtWryn59VDS0pPR1pE
BSJk7Jj/DTlycqGoSE3kaxMqBK0e6L/nerMpkGHfUHk6sb0t4bjXqQJspm1z11jF
t5SuF1bI6zhnErA4P4Cz7g9JID9rR4g0DCWea3VXPSVakBR1wk3S99cwOv+Q4lh0
nKJgSZfrRzgKV0rWMK0tRHfdNWuIxY7t7YZfiE3wYuVDeW4soeSXfjNYqNijL4s3
F/5ALZU36Be11sUVPV+YP/Z64JRN3MHdM1LDlMcna7pdpjfb18LU7JEqmcRek/OW
p4JyvvUxj5PnS4o0Jn/4fZcG808lRTwLXL9T+4FsFMOs+FN5W75feIFdqjzCy5tw
yVSsughDPQTAFUnzhFBHyTB6Uy9d65ejXuSVNj2C9PlUBfSpdGjKPuG3tXMpbRfr
EbU43d9mIbMe3tXxiJX0RU2NDCayeBOiDmY+/ZPNvbQLpL0tGMAyVNxGYZr1Two6
4kLmoLara07dlmuPmV84PITJ5OwAt+UUjwZ4blHDIDZiSTOlYh1aehayLD7v3yJM
w0Oq+dCaifRg5UEvpo5rITmGck7ausrPiFu+oqPmj9O25HnJ/k73S0cxumcW/qR/
ZwG3Wyzc/5oNDXiCERBKbvTC26yQgppoEi8kfA94UaG6ImLNrd0UDJCKTquzF3Vp
F2pfMCoZMh4yBwtGsz+nJQRV2uVxMBXv3eVeMC107KzYXf9pbFjdXzu1vjM1EMwZ
V8DrZt+9+1rYc+1A+xhqZPmvndThc7w9NhnQjWTY1444vDPDlyxcoU2D0fqdD8MV
BB7B9rpUN7bQZc6oqC1UmQzDxg0PGURUn4VW/G7zfDbhYkrC+REGa9UKpk3O34fk
DkA6YcuMMcr+8/wF7mVSNa21RClKqigns+gSmZxecg2aFktFXLZSzWBRXeAjgnyt
pbEGCItIg0euoYCzDChJrvYgTE1zc8CdQ55KcwYunwa56lNd/UviMoyd43ALyeKF
H6y2vROmmnxPtm5liwRWAvMdDpncrCaTZ/dHfh2YKufcopJWEst5FTXtR7k2hxWT
IhXab2AgvDXAA88CrDLGPHqvLvyjPDaDzPZMxRm1AM9THLSt708vs/JYYGFrigC/
FcCQi5kn6PFXAYcjhMLZyNGNNNuSie62tvIvafmYADAkDTWZe/49Es4g+h2D3TSe
R8NSuMfoLtqnUJsmqrgnYELANry3O+i/caJpBxcXxuRIsJnm52Jbjwfsy7ORVxiC
cG6oZG7RxQlZu3FppC1YSlcuNoncOrnoLzp52gneRKacUX1Q9mFrJWVidZWSvwAJ
HIE+3EHRuUbBrpVJjfdtfETRHo4NUy2i8KqWOod9C67UVJkTmEpC1wXns8A7CI6X
yxWXvTTYjf3WDmT/0BBOtOnUChjKuTjYXE0HGl/BgigRg6vUN6AJiTKbNCCrUWS/
X96PonYvLCL1bH5RDG5N/qnBcY+IB4Ka9kfGAQgfKHg2vkeBpACKmi7BG5XQoTpX
Hpd0NoC/5x2R2ic+HhIHX3fRNKqvzhRxyLltDJKTU2/KfIsg4yXp0MzIGQIUFiRO
8MB/M4pap0x+rg/alNzpTtfG2vvelppSKPblEy8Qsj6UEUur8T9gU7x1M5A4ontX
k7uqUZ9xHW7iws6s10nsIuiSy0IVXai5yupjApOlfsfB4L6vZDQ4AoFoUY3Rtgm2
r6laCjKVlTxM9SE/tcKnjqhXry6nh7bTB242IrzzhylCJVWyghM/H5gMvWJOgxMC
p9QVRF0F90J45SVc2iV0AGGRNb2JAW95nfT4HCaDM2ZK5RxqPBmcEbV2XDEC2zzc
63CJ2v/pmlXT1nPUvs/zsESWzGRDbXDOYefpXjhniTnJL3vVCy+czz/C+Vcf6sPu
iGX4iOZduv/+EIuaIboPWMvy3gQtDImBiJIf9ykSMcr6kuG0Dx8xUL3pyi6T0Sdx
cdPqPlOJvNdrM9vjn2k1ck8cP0Rcw/oOsS9onlyFZk3KFpgrWypUKJy12Oxer5lX
C4q3UvQ7/iIM6d9BTPFIvNcHjVWIXhYY6kctPPckW99rkqXpA0awtvvZL+Qr9Aky
4GeQJ7Uk5zMwDKoNhujtFtD98W6OwV0N62k6JRKzWhq8tn39q2vgvp7he0RJXt+h
HlRmf3Qw+r1I3Q/0he3ZdyQhRpWL+lRTYJLB3G2/aH8wfgyhxA4AF8UH07NAsMet
O49ipFoI5b7p58+8X3465yMUTdXqEZhn1VOC7uZxkvPoWlp1R3h6mbgQ13jFu9pc
0bxAismA03jFlRZKpu5iNjVBs+Q3vpdbk9HFhJ9h83jxS+5nAO0xN5lscjByx6Ii
jIammSpqCNXdLdmj8gF9Wbfj8fD7UK33lgaUmyITc09QqYiyCjsybHgvJEWB82tg
D77iaF55HgJ01BRHJtqDDugcYH95A/dy5JJHJgY3Gvlji0nrU4E4e3+45kBft7Ho
fw83GcQa0ZWLJae7O/dTXV8bHrw33R1a+6qoF/8cOqT73PmtiwZz8a4HegoO5Mas
CB2byP1KjAYBaP/0/pBuCnZ/wbM2FyvpfhQwemTQk0+20JZYufGkxiDODc1f+v9c
1t68hwO26klcTTMIlL4gmQRG3+Q0y+kWWz0AZFjq0CndItx37/y47WL0iuIYf3tu
it2DAMxGL3QMWIBtNDAK1h+RZp/xfnLq0Kc4xWCvA8JJl27u84JPYik17pB3/4iQ
ESqQXc6EHK9SMgCQ/11sf7ytpUiVt8QTXdyrbXy6TRjgf6HLvPrHylmx87r8IILG
4h0k8pzUOma4F02s1Lzdz96Pk6mS/XoQcwji5VhQVkn3pAyl+6uBo7gCVOqmwuJL
9cfBOBFor9qwYraM4F2HcK6wrC3BHzho6ieQnzrKxI8tLDtdtsK2suWCB9WhNPr8
cxRM7Kk/Og2EXSCWFm4OK17YTv7dutBCvtAO0hnM3OKLPzQaXvgvEOcmtWOJWUb/
/GgyIK9tzddPO1mE5lnuuV3gDEXNtKvoUe+M5H+Vm6w+ABATz/rSTd2b1kl2EE5F
M0LYj1Od7a32HZRh6RETO0IBpCDNIYP3JTQ8q1jxnjCr7S0BoZslnSa+6TP23FXS
9ximziVB1P6VM0SjwPohO0LpRCRvXvmxAb8vcx1MRMBBEhfpJHyrONDLubmyzIcH
J6jjf/ukmoNLAoAVFFqoKKZrjyO8RWkUi5c9AAhbt3BWiMeEXFdUmEtEVW0fY1zv
I+qYowiw3p50cDQCIY5bUD2FZjIOXIkT4uZDtqaTY/CNc+N421UL6XuMx1uUGgUP
lRzmfNG9bY/eEs7uaM5LgIfTJIwYUtkm/1SsluXVHD3t0AjKV5+sKNRImtuKyo/v
o9Q4JVuPNQicxsHzICuccr9f5ES1/4uQFD91zBpCAFmsOMAvjSjonWB2ZtwkD5wK
xH2KsZp4kBuaDPIeFPZ+dV8ODSSka2fnfd/yk7tvI8I5TWcazUwBLCnvqUoSbx/u
n1geOJG1fjJ9wN7qX25OCYcb5zMUi0aMVb/VT+mjSH9xPHuSNawLeGuu1J3uuE4W
KtC/R+zkeKps+szXoIayPWy9OUGKF05vXZAd0DhI5csvfYx/vZ8aoBaGAod4wZ+Z
1I9OvS6WAFTfm5fPOJG8YuRdlSbR17SQGBqtUvSy8NjazZfDUkhdEQCUoNBMyNZA
YXlPz6piyIJnMWGHel4sFYbbnwOBoRFB0r7OL90oJhRUrrYXwQTcGbwi1Dzx6g5J
6Ifye7Z2ZskDxE7bUJGNqlCoPnlE7+outtlXkqwDsDaoDEsL7iNmgtW/AoGTgPFp
bYA+JdxHXFRbLDiD2TMjj3v2pWJ0Rf7Eb2ImFHPcTpjxP8V8nOPUWZXDvbmK5Koy
MSjAFOyugDpKibCjq1WoNdTq0ngJbOE4hCj/lJxuwVz9bEV/FZKjZnX+Y2s5QuJS
ZedJjyTdvSVsrpwTfbejeFl2VTkbAHXJ6RdhsYd8K8+v4y8HH/DK79JSt2MFCc12
3U8WX241GcrxN5adaq6kEas7Zk8T5F1nTqJBCXy0UKDHF505SvqyXrssPhvXI1GQ
kyo19NqydzrFg3MDH72bVa7fuWjpnaWz7aV/o2TJyNlvunky/rg1pG08yIr3LenX
+DrksFaO6XC0uhFrVwKBLYjzikzzoG0GyIVl9GDhFpv35+5kcE75Lv+ODOTrw1M4
gam/UGGbrePqFiqvdYkbkXhIzv+NolGvcVWhQdVRnIWkBzODfJwBrK/H9hY8IPfO
f+bdxDx+W+4Yt5E1M99GmMagSm4lMBGwunP6F9zhjojfLBIpWE8m1Mz2e8MxiYmS
hAb4jXiIZ2i4fh1tl+A86oxaAYvl3DPAl7dWMz/II4Gst6qE9tNlnHoigOzL39lQ
OHFphJ30ATrNlFYandrZwXExT2JwV6T+GikJRJrhaPX0TT1bXjUi8LN5qHTyLp3S
/x2MlZoFQHbt6LHcVqHiMBpEKHF6Kfp0vAu+ySGZKcL62V9F0G2yma9natEGUWpQ
tu4V3p4DL7rKr0o8IFKiiJukfVj7zdO1uqDrnDWlhr/fc05qpXJ8fHGZRhT5ntgJ
yzuYKcMoO26pJKu4yk+D98V+DoxJvQd31yLxzxDjiNE8c6dqJHSA+pzj96G3RCAU
kruoHaMGw6LLdq2HQUrKjlavXgQxjVpt7LcCGuSiNjipMeIyEAxdJwuqKDiswTdk
0VTjYU+niLl8UTi9gWh4YmeMlvwwMzeTHXB+c2B2pItyulDvflRwawjTRbhbkPEC
8IbuDxW/DgzGl4V7XXp7FLqt7jT7cvnH4Pl2rfemOaczqKjgWomrN+6Bo1aI8woR
v+aK7nyr935RkUMNRN8QJvJuCDTFbZSEE144txszRb8SBWo5K9qO+0QExbotgbs2
q1ld/T7wXn0vnHb+WS1D57KEpUHbXptCPgTHfaKpki80H7hu9Q/Y8CtguoTlKAIb
zycPwH6gBq+kcYq+I31PO5H4CSPHPLVFIm8MV8uBYj9XvVwcsnFLz/thV1QIjACI
lrmEUJF6qMZrm6qRiD8fNYCqO+in0L6twhm6k8kv76JXfLYUyl4C1jhFLcC3c9ZG
SanZonQogebgLkraNaYIGk4+o6rhBSegf8cROOB39hpY7qDtjuxZ+yuPwTpmM+QY
yi+Y/qXPs7YnJBaOuzaIfibhgIvK2tmlu0Rxlw9PSwml3GSOkuDh4cGKTahu46Dh
WMuJdv6+EgKs2BY71KFSG5kOw/dG15dfuNCz1R3CcNQLoiyFDLx8Gk1dE9vmvEYX
9reX1E0lS90ucnl6EkWvquCwrrbVQEl3efxYdD0Qi/Q0q++A6ybcKxK60BPOx4xO
EblS4GgIiFyjuI/ARvy7KcatYH6RAYBurM7JoslFGxYjjQG7t5T9K+BZcjcNJVb/
MH2dnhboeTio3hHo3/UQZq0FudrAQmx62KuU6Pw3di3n8sH9UBMRsLtRjxZl7bCL
Y00JKk59CU4g8xEvfQbWxNiM4bhVgZpw9ALaaKVbfZT5FXDtooghS6qmVLSRhQW6
uiWM9iqbgT9Z8J68ws25Mpj+W0kCQoSxGowlXuyI8si92+E8xE6j7/n2/G1RDvNK
RayHomqSsNlFJLpZ0m3YDkmnkt6c6lPwhySVtSdIVeCfRJX3Hk0XenYog7uKVtvS
GWMRcnw6rUd7wPSwU09BoSFxhjgrKRNa2/i2kagGaVEpaJJqqbFT+YOw6IHh/g+s
Y5G/6vl70qbvK14rjgLj2GHJMJipwpJLQefT4ctEJyMuSM4nZS3vBLsCfR1jVqkD
pI8rwiFfxVz+yxh70xobczK7iRkQXIfFgCXgJvWDr2EcKZuF9i1FYLcJtdT6oGRp
66fqiVtD0RNk1vLtRSCAXpcI8wp++TUhI5o3fpUllxsEy6mQjIKxA9Myno3thnR6
j+IuZ5+j++hmDj7SCJCvhXFiXOMOzi/9G0T3YViljc10wSIh9dW9Z2uTcrpivHVA
4c3V9igADvn9m41rDmbK6jkE28KCvXeOkxZN6GImYqd/juqDCMlZXJzHQ/0LUKKN
+guQA9RtvieXS6Z4flkuqOSEmiFJmUGEA4XIPkjvbtiJMdosq6eUdEtXpV3cFwiG
GgvhwWJ49XbqXsAHX6cVmYt5ZVQfEZmKQ1qZAHrAyhHJyTW6V/HTX+ASD/ZQLEWE
dSbLpZZvS8u9XsyDzoyPdC4pKFaV52aSN9bQzpTbguJmeY2Jol/NtbWgx9YFX1LV
xj3aqzvf4DHEbrLqvMqqQCucVZK554jTnO2VwvtMTesY3EwirxG6Bx4GzGvailPv
wB0uwxIoqhVEJ3RxPQeVrDPScfCfIKa4XQE9/oTHa746/+yK6YQsDgEY4qSuQ+vV
QHU6KFcEV/sR8ucHvs2q0u/l7IwgYy1L+7/7DGagIthtkgcIlUHEipyTOSbzPeAe
kT02YEO9Sd7BmonAWr7swRwLk4zs54aMjcW0oC9nfQR6eBHbfiiu2f4CBkpbxvod
ssFl9rfKN42oyfXsT6ESchf0SSItN6hOrAR9X0eU07MFNPI3YbIbNuTVjkNKIEvT
kPd3VW5RNrUcQoNS+zbBgqpnVe+mtqGeD4rejc2Do0gYS3JrzMRUZwIsXlhbZyu6
f33McgLoz+MPEh0VRLOJ39hf3CGMEBcA6t92Ol/w4jF5ZrSwg3QQFKkIVW5XtqL7
EXaBsYgaTB1we12hJzwQ1R1m49QIpQ7NHpxtme+bNriBvB4g3lGwy7WxtA0bH0UH
jr+JPBacDWuYP4ijkauxxZIE120O95KHaiRbndpJhQzwcIjGDVMopUJd2hkafXCA
lt2esiWho+M9rkg/NjLospBLubtIxeZ/rePznYq/MVC6ZMfMIhxupZY9YUcf5fum
aJkpk4cYhAbk7Q3HJtpD0cZUBp9OqEqzI4b8GfYU9a5ofr4nZeuvv80Fc+zl5mk2
BJt53wZJvNKFdsP0eqGV9ZwDPnAXug40Re+/x+UR2H9Pv5DHCl+8emydx5Gc++mu
ZdGSBXmNO1UYZYDUAmMkbzeV16slCUMOccQZy90MrdngC2GS8/31Pj8Npy/LR/Uq
l0Tqw6O+RGYX8Aw8ZR0XxM/r7o8uVkuuetzgmI0hMyE8sPuAp17+iSNhJOZ1hD/q
7s37odew9jpF8QHXm5+vaq09xe8LMf5dVhq7OmpQbkbHu9oXiRcsciU3ToYkEA9j
R9xe2wB5fR1yAS6XxsB9WSu8GYrYPXofJoAav/0g34SooKnf2A3IsC2BhTGhdQ5t
+sg31nsoF/QYvzGrX/FwCFosPdr1vAXguCNdSHKHiA0bZtrb5lrKpgxi9hGWnKtY
hul6RmyJnrIOV914GEai/umAFbYEGaLdcCor03iRQ1x0o0JGJgb33z0RgXxDpZQd
iKznqesWnNs4BmHg4ZHJ6jjLYPLx6IPnumqrQUzaiBiFUrmXZ8BOUN7NTPmLpFWI
dFtwjpEvKsatML/HyOmlcpcOzlYTVIuFjAqER1UWDE270cSvADg+ahjtIoQQV32n
X0K1CFW6Oq+01p5v1gDfsIOlb9mcdga3Y/Mk64bZR9roTcduME1/xEFs+f03omRu
JIOTOu2K9oY9kLZcWAOvF7YRJArng4Pai1pM29mCeMzqMpfDlz4QB0qRLShUuLph
g8rzNAT1Rp18RDOhj4PYjxFaLh7iZtoVbooXYZOq96gfpf/my1N/sRNDax1ur1Zm
38UsA2qQBYWy3xtMOHbbhQuP7PJC25wZimOvDoYkqZQdoiBZrmj5ayNcabtVZj+i
/P4dv5/MHOPPy2U1jUYZL45O3TCaWA1XPlPF6XVBw6aszuWTPCsXWNFh4GQyAdrI
CCEB37tiNQFmkINV62ucMO5wpsgEJn0AbfF3qdGFm7lQDVJPvjCtHgeyP1i+Njkz
H/YRZ26XT5Xn61rdmTpP0aI6LzszROfHz+/v4c8oUqI+GaDaoTnwpDjUMQtfw/PG
d8RRlcS/xKJTGXOwUjCRrmjiUhMTFSpmQjR/X/oRtl6/DBNeGgPheQRwQeVD/5N8
SUuvNVjo0SbHKe77QfkXRFUwSPKqwgMgVB3jlvRXGpiHmIB5MeA0uGlSMbmrcABV
ak5mFrBxjK7KGhmjJgCxXhOyCaR+shX5sTdsiO0IMUpIv/B6yiTf+Ju/pI4+gZys
mJeTQCANBLuFFH1yfMUwwK4UXKL7BwrjRgkPBjtUPx2XmEmMxXquCA6g8XoslLV/
4YfacBRMzP3aKgsXmljuuiYsrkGG8sJSmQMjCMBKAMISSKNiy5EDFxnQ1yg7aD3Y
QePwIqVO8lfUoNLzcI2zjZdH/oD6G5+q4n5olHFIvOzCchmD8dYhhQD78H0luQnP
N+r8E3EnyBn5f5nswpLhpfX7QGa13deuRbhmUHQsYP+ge+/604+PbbcQvHlhPMBj
zASeTAof7zjsFpQWUC4ZUffbFGJpUNP5tTXNzxNXJMylp3yLnXSODLMm/DSDYmxD
ipnbxmdYif7ipQRCIa3n2BuSBBG/vUUCHnDmkkTazDdl9fgmExNw4tRIHeyq0Fy0
oppfe0z/r7pUOVK5R1Xi80WwGJSHBdWuVgnCgqPS5zE2twhqBtZEcVvPNZi7rSbQ
8DXmzW4RJevFS3gvOcGnFjfVfEwjPW02D/XcPObfX2hFDA/LGp/VBIFfnpyzsByx
KQ1M2vu0W5AF9o3sCwhObPNjzYteDcoAcghMGt089LmSTS2hxQDypliJUJMkkgrG
VTyWBdLSdI5dHP+sl0HWQidU6LmyTel8JJnrlg5wrmBo4LD2FXAJ3c6qS50RYxG2
wfsk1B1Y9dX4ZvBaUahfJoUK2A6+nb/Fg6ezhv3bwTsQA81Yt6qzTyaqdjzQHhrF
gHNLRroPLdAi7ExN5K7d+rpY8GKpZAyunnfNfq8fXvk/R8jUSIRI6nari7fobWCU
OmjVOVErRc6cU40E51gvke0SwyvV2gTAAtQ7zWJNS0L8Uve4EoAZQ2zigahPPomY
x6AW2pueDmwUpQxAJVnLLzTC2bkvI17DEvLcZfglZLqtdtchGOd+9Hpo3Q+5B0Ui
qGggJ8I9q4MPCaFEM6KS0JARLyRGzbdRlb7lxNXArR3/2IdAL1CZasOUnPjlAH51
hu9dcFe+71ZPzb7YHKnUnsH6bkPcS8ep+4Kpuq/EFJj+p/1Fk8lK9Qxmb3lue/KL
4HKWkwGgyngknGjJ5HoO55a7RHFxWDTCP9ZsMuM/RvMXW+ODifRip5cPPwkgB1uC
hoWtDyNalpK7ui4Xge2ZoidUKi6aRehgNfP89cEpHqLxi6pr1zlmakGLebWc7tWk
sL/RZitGd/RbOeyZmys6p5IYZOo8IyKyJ4tzAIP/jkN6mMDC+a3vuiHDX+a5oXQe
sV6jSv2qslNgBm6CMEg1PfRZU90ZJhPMYVGA73zoomtU4Q2/snjlg1Uq++KRUMKu
rxraixhGq9gUPX+feE+WP6fVTC092dlZK+aFbBQnZhFqivewxVghMZDYMyec97jK
KAlFqaxwApJiqSMowKwJdFCxxrt04lNheoYZe0OBRIA9B1jYKl6k3OcX8kWb9ddl
WiyI1knfqOcEg+yF+tfcxl8sYtzBHQfCG4+tU3ARgbAOCatjlFCZkRyCsAdvr4nz
dtce36UX7he7wC6V2Aj+X0mgOo5W5haEXo7ZtxrSnzobDMiDhtbe5wLmGYTe9C12
B0ztIgE3gvrPPV+Psrh4CNJqjV7GYs+dP/g9YGchP1XUchy6igugB0DDu4oYPNCj
QCEq/Dz/qHVnknfr7o6xddR38F8i9vCcAs3FHJtdf3+OMmcFUQjJNJ1hKfG0WdUY
FNAYbqMZ107x4CBViHe05ffX72C3AHaG/XVrxFtc494My+JdQDKW0nrvSF7uJ2/m
jURWt9q8eurLRGxfcKxSGp59UyTo0HJ/q0hukYmmzTEPuspWq7fRyblJLft4S+8k
ZulaTOQuCeoJPelwRK31PSqeNomvyHmyVB/pNEZtMAClxYnvAmlp55xYPunvidDj
3s5bpbvlp1AI1oT4OBjV4b6TNvvDeMAONjPGkrnEgbxqICs8ZDXN7NAKNMJaD7N2
OZ9eWkY/dIeN6kk7j6/hySclbEqLuyvqMWgfCcCskBmId9m++Vl9yiR0H7AxK4lP
L8G5CdcvEN8XlKg7Uq747BmIIL8UBb2YZ+kHMUaCZqHKG4xWWkC8WgHFfOz23tvC
RplgMnnYybGdpd0fyawH/A7/EYTRSTGk6t/YOqk6hmr50TZuXMS2DH8tNHDzi4ns
NjE4X+LyCD2G5feOeM365SSWpsuyQb2OKqsazzNykyTIlUhT4byWIzJBkN9LSnRa
pKHDPjf6W0ubAuaSb8/m5RkRXWfSO4urL9QDQlgCyeYizkZGm8FCZaxO+3+ZimsO
RHwKB8RB2IVXsP36U/KGAlnEwoDm4CQJcf85qZX0/VZH5I7wqIxg+DA6XOAjBJgC
atFqYIa0rgVBVQ7qnKjShA9jcjlaJMY77Hxku8eVi8GXoTTqYqPjscajTyMAWMUk
19qH3T9Dud0r4m0DZaxaef2RuWyGXnO+06M4e3ZkPEf/RqIPwYuDtkbFhW/cD8aY
RYOSA3G+95xxhkWQvwH+/rZi+HOsOWIo3ecRhcmk8WuoPrhvR5DKZV43sxGpIMHd
q/XApUQzZN5ULgVk+Qza8hnfvZfpMmw+1SHEzzGMKz1ezXTerO1VXzDLV9ChmCOB
wU0oINH5NkxJ9XYmUTePEawbf2upA6EtplDB5NTLveRU+5GLOGueHmSLVCyNeNjt
PntTPCf/80WHzSb08qQr9BbOYyKGjFStBGzcb/WAJVJcfBbCEFbwxZApymlHYXeh
MzAPaWq3ZCMZ11UIzhN0mnBzmp89exjCESGY0jbzbbtDKGdSMn8e/4tO/59Eav56
yWB2xdVdVVP9TQFTCkFAapTplE0YSX9U9uqjMuhPEiMBMGoqpCQ3tfpn1Z/EpuXe
Jzv4uhV3rGZddRhXL30KougUB+/YzM9qcdowUNJ5X5acrCacKsnAEMa0xq1VDbAw
LYAFJr5qmQU1RwuCUITn70vWj8wK4Mj85F9/CNZFrIl9pZFg+yrushazockQBrTN
gLMdMJS+tbeLFbixMVwkTywWWgJxsbO+3SW1JJLDDs+IDTODhpznAVu8PnlUBPnK
B2iucY2LnJ5fzZ4DNkme73BTm6aKp0BDXqlTOVJJIYF2qNdMbE8BgaO1cvIxbUGU
vQweR8u+yJSLxcGGtOejYYKL1cGNYm6fA7D6AO3bEgN9OXqVYfAYtgTS8MZwccNq
6Xmk34yA5F1a40ErGvh96aF9BIUeiV18U65JJLCwbvgr+/BeVuDcmtpBAstW4Zrb
a5M5L3viqoGkqp2o5F1EVEUpOO0hSrTn/xot95rEu+ICcegFpsQ/XnhYN4jvhaYB
LGIm0vy2qIAq+KmsdisSF8Pd3dXE9ACwOrz0L2FqMTAI4KqFwK2V0iFeLDshR2fV
tFpm/c+Jv4UaPReFyi2AA/cWp7exzjbjMTQohUS4jOwE+NlPAa8SBRhcUODlHlT5
5wJ3Uduh/4x3EzGdvvNM811su7Qb7L9b/wA52uNgtbHyPJrm7+pytJfTyl+Sq0mf
8zFSPtf2Zr06KiddtyM9jbmDD1McCeSt99Z+d0pkCmYXfBHg7F8QETSYkmZOc9qs
aKyPCmuOvGuy3fE1IuazYRRceV5wDpQmkgxhep8qXrvwHqCJe98Tj8h6CLrIa/xt
1v4XDL45063I4JBBrmzOildrc9fVcTPfD36yWczhSkH1bGPGEyv7PzCvkI3joIFe
ipHSwF+gR+2Q0bfiaMxWYr0GnTmWz6map+cvwvqkfaDsNsx7HMUb3zJDD2xqN8wg
K8K9tKwKNsuBx76800Jz0ozNXbSMYIDwoWouGRilhURZsIrkTg09/9Apse/sLTqx
mhhBQeaEAkEDKo5WE4T97Ltojso7hg35FJJkzeya/V7K3oS8+ps7GtBqR6OTbZPA
D5B7Cuq4M826PjtDhTPaGqcHs1S8WRYjcB/GmVZ9VBiBKU5Vhm2a7f/fznWzsAkS
0/I9+JBt1uIJMeU4qXZqQChAb105KE4vd/H4J2IPL8ueO7O84j/kf/t0vpDRPZun
vsXFTt5H9EuUyakavpXs0SRDu1bC5dzSuT56Ky5TUKnp+xf5fv4Pct5hpu+Zn4Ba
M+urOLym7kTcJ5i/QJ7rQgBOf3Znu8Dc6WYBOCm8dQgAregqzO8VGZTFDEr4xCaS
fSsRCo91nNYqyA8dcuwYsaGp7VGlDD14WeJWJtpfjLZWUTxIyVqZ1nsTGXN22qng
PguzswRm75DlSsvJ/+MN4wLLOEpCMp+8o/ZonKLIEjpzQGvhRnJPOXJpXH3PIJCM
HRqFWElqcRP7CK5k1Zq1KucvkBt5s6XQCy7gk1lZWNy/izQ2WHr/fMY4tL+3TV67
0p9oydJpVttqjE9PD2732w7aV6t1AyuZ3nCU5iBK2JILbSOXbHibvWAhOm9xO1KL
jxcLdCLp/5Eh4IboR1SQtqfpOWc+lgJL7u9BtQM59JKYdaVGvWKWtQIVGpyz7+6i
4eIZGBndLArnXeeww07BhoE00XfU4vWpoQng5WxnkwpkyWXJtS+jBCNV+V1Lso9S
jx5rysoX+OmTj+NDXtVW+o+m4x8DZ0o5WWMZUaJ2Ya/4Um339HxaLD/8HdBYkUdN
t1rfoFhdSkpszRoQ7eavMFyVT/q2Hh0ZRDtFnQk1korA7gMd2u9GqhqcGaxuN/Qs
ZZ8WOatObTD8ejMAKmPlVv2uW2OFpCw8lXEV0d1fuVWKUWupsI9MUVn+mswyUY8i
E6QXf+CrPTTcYD4lNpQsjtUHHfneafn4ChuMMRQC1dxuTFXw811TYPU4s2RrvfGH
82yYReUTG8zQegrFAO3PTSsXc9kKkoxyIToS/J26oRtf9FoML0I7r6aOP4Tt8FP3
Z0t9ri2MwCXSQgNS38a2mQevqt/6qBQiZ81YRX/FYr/55+zCHBEy3g0daxge1VAL
dORSNmKA/Wnwty1dy5uEnC3gjUFkKo2L296ELERseT6fwGknOMOo0i9ZosxeaoeE
YJmjWAPP/vZ51AOhv2kkZ+im57dWE+KgGe0DXD96db7/o5vi8lXhVJQS8l+CLM/G
JNLvfWNHKmq83cd3HsKXn59VaA7wE21nAbWta6Xc8Tz35iq2ntE0h7G6htbvHCM3
b/Guy7DtGWvsLxgdty0OqUyId/a52zxMtgukSsLMS6AtB8qE9IX8yeSW3UOqNFli
1yZPKBjS8KVA7Fyc/m/Mbzj6s6a52xUwM99oVDenGLhzoIKgltBavmsCU72o5yyr
FyOTS93AgFJFepY5MAFEPduU3gs4Bt50HUx5TFiZq3K+eY+mZIP9petyidi2fkp9
heKsFeWTFkxGqXO0CrRrQfN3sV5+TWH1nWL31fYB4oBhq89W2vrNL7glGSevjfr0
yWVyd7+UeJ79VGGDPCtnSBN6eb6uaEMWuKzBFhT+zub9gp5Uodg9j6bM+L6QxrfZ
yysC+abfttIEFBUfGThkIaahhCmczIQMeUrV6yw50HKn+0DcD1f3T0aOTvryRT01
u3PLrXyQwkYiB9MTH+i3mBf7WDrEpJ2QYjIOltV7cJnS8af6SmBR1Z3cXg1FTAqk
HfRaz4Oqc7D9/YDH1mHZ1D1n3q8dClM15W1vewLvuPQn3SOfQjH13RGIU9VdMUnY
Ni7ObyOgATowcZpfRWMN6BNbqACU7ffpO9psd2zPOKWmiVEdLR2rtnL56yq/iajK
jCbh9vOafXyKxn0ED/rFg08pXAakdymt5i88pu4w7wF9okAQfQbM64IM+hLzl2mK
oGgdx7MzOLXtXitbDcR/gv4LoBm91x8o5ne14N1rrfGt7lKm8M8cMu1D7vSWkK1I
fOWWelLX5ZD4LhAQBMc8l2x+BP1epzrmrlflIAy25zJHhSYaYwNO4rHjdf0Q08bp
hDpSQdPxQkwWTAJyK7Vty0McaAkGArDxKStQjpkteZhS4GFQzP2wZvgnJ6slupZz
yYKJOJt1p1iemBRcReWSd5/CjeT7oz61ZfTXmCWegG/DOeNqoZB7K7mmmMinevVf
/uCXFPE4Dt/iZGMuLP6lb/M68bW/ElHleJtW/PQ4Pl35Ms+Zra2RNUXDHohFzDRa
1lVbm9cgN5ICN/71ZB8ZXNf5sZGyUrHoarAqO/dklEFHLvhlMXZs9x8O0Vad+yBZ
7OiPkbnoLR/HRnLQ9MLyO4JwEL7TpH1RYga4G70SbYDHeZHk9Avpjkz1iy+7rjM9
Tx5vOAqMg6euiJWlig/oa4kQRJRnMls4qh+zj7pJaVICz6RK8dput/jWE15v0E69
Li02KHD0K1LNVa45TTI41/sG66TAJ/8dVJf63dZ1JPDpMbOcdjXj1paSHytHlooG
qZIs1RowD6x2AteIWAeb5PjUCDigCMDX8RUkE8AXysd6PMMdHSte+dIkPDHzsLp0
qVMfymI1w7QEhq87zYafVOTr27M7y1DNroMaLZs4rR5sgJgPvnY96dtGvj5ld/nc
FaivXll/pyVUH6JYWoOp+gyIqwYnTTCIxyARtfhN2VxRjQ3EK6sPyLz3gpyyEH+p
9ZSc5HxyQ8IobDD6VuBz2EAwC1FLtTJ3N/SQMMET3qIOJ43RMfXEY9zpan7wvljW
43qLkp5cc4OzZJESQGj672yQMN0/xZtp7DoLRop6B1dAhq/m++IQgS+aWMvsBHtC
Nvo1pO8FgQvBBtHyichjLzygGQpQ5anCwFgqSoXyUYQbhhEOQzfiPjKPJTXJKg4T
e1rLpuzxiwoOMrCopz2XQLJ7CjtpJYa84kcSgHdcwQDczNtJS/FgWPh48BHiuhta
LOArhZcxR+yiDgNh+x6GR5mJGL6UJR3x5vVkPG2+3/lcJIcQ5fokz3qWdRYNb1A6
e0hHnh8ycsk3zkoXmOZF4h1MtTqcIL7BLPU9gLbNkmHcVCV0V1v9Atb0S/TEX7Qx
5BZbvMKGBN4//2PK+vVzNyQPuhqfZiu0i8jny7VSKMLQCT6fbjXPdw8JFR3PWUWw
j6saQbdqdoiIFk4hn+yLcVrfppKtsmuDnFiun+AxVUpimhHzQFjhSwjPPxptCG1F
rAFc3rnyUt944otJJ1FHqNOpg+EPJDc1dEnSCOEjao4Fpajr05gJOHR6f3ccNKVa
4HxQMrFGovL6+/hElQK+2wMQprTLlNqAM1aY9MACqMUKBgz9mZeHHU5aOwssgeIu
Xvfj7SWv/yGMzWpHtAfRw3aQghxdv+dr89bEz+WIIgRFpOdrJo1bfNoC9HntKgoS
L6/j9cYRq8ZCC+VGol14LNqUP2XsZuD7JxdxftK73YXbktE2OrwFnUIwvOr9Y/sS
yDC+kdf7yM3YZ+Uymjp9r53TpfD8E1qdsHr6/wLw+TK02DglGP1/d5suHD4eDw9S
SPVFnsqyPEw+BdYDQXWz2yJkCwwnBXMJqQ1tnUa+wvmaFH5M3Y8f2tERZxJKEtli
r5Zn+/u/TjAmr4hzyydGMJgrclSgC4BWb2/xmKaYQ5nrpA5LcnZcaHYHh+UkaM29
e30pXXGqvkHzuS/+iM86QrjeMp9eY0VnyDmuSihhl9LmZHMw15NqhlKVxutWCZ6P
a/GHoLAtRp/UVBOmv96bfDj1Akc/l5pADd3dueWdKqWdrokxQyf3skfD3InEyDSL
ezN+81PT9XEhE/kT58XqQrKQ9WsTap4FkCBHFOJIusTS+mhQ2D0tdJWG6/YiI7Xv
23XcuzwOmeSR3AbXisK29xQbI4Rx37p+j6LV+IBoI6Px74JvK0DReNEKWl5P+m29
IQrjOesnquSOcJOmljQtzGSRFbLoKYcv31eYUUOcvdM+MaUJYIArwohH1v40ziyC
fKEaGWAg8ICctEKQLKol3ZUp6P/iQB9qsEyJrNTY+f4mWYWHTs3GUj1jhqopLuwn
OMP2sb50OSsXGdWLyKrYwWGgaWDcV4qx8sbluZvL1HR2dONxUZI6LW/rYXehupeq
GrFKNzdCM3IbxOfU3tiOgf9Yoy6g0AwkCuwbfeCMRrN7/ncEuyxrK7vwW0h99p/X
m33RpV7OJNLiAI3mmR5KGDx0ayXs+dBVNBQF0gOtuYH/jAIfBI/macCobGNdidHE
NepaRnqmRS9eeXnAjwnZYTHHsH18iXOj+Z3XELr4miLbMRrsSwrzgSyRRvVnWLtv
T3x5gOYOcknSD0h2fE4sEQVtbC0eBALTuEQK4rKGtnUueL8qo6wur22z4489AqBI
2cQyLLwfwW6vipSI189o+Nc2JId45VhixQpRCv3UJicvDRNgZE6xGjiKuS9ewFrE
PANuGFhnz3BPlF/ONOIBQIaHJq+9Ikqk5RlLo2R+6qLxdyysDCR+6SsRlPO+NFEx
chgX4BzY3Jgl4CwTATMnIOdPpPsJXCtcKLyD3VDT42b15PJ/YPUS1ltogq1fx+Rw
hB2Q04VGmJ2OGDujFFdd9gITHQYr5J96n3UyE+qXgwVtpI7jeg7TBNt/tP2qHIYm
z7exIPmL51k0CraYoqlm5s0mDLbmjHU+QUW2sKSEcg0zQYe2AEU+VVCoE5EzDzJE
NiL54qCCvnRPO6lbE+sC60BTMHmJnvwHoofGwgc5B7iJ28pIkK/uOj9ElV5QKfoU
5XH9n6rqe8haTHAiElQ/A68/Yi72NTkJkny0KCXI6jBlOjqcNs2ouUV9R/rM4GL/
GtqxQDGJQalb4TzZz9oZiKfHsgrm3HR7ruOYyyoNWNt3m3ZR90mXn40lfXcXbTUq
EKksGVgyY0mjyLEb6E4NTN5Xt58Stic0/ZkkavHgkbO8+A88V8Dxuj31+/i73xR3
D9JCE21QnMJMBWd5gZVuy0WBMu4neP1arGmZ6lqrm+Qd1Ag6eCJIjePYDyOdPiO1
joRnfXUx0b/mm7voP5TCoDcuXMAI2ah2z3bQFSVdI1rC4RpNbZqYZYwq0yILKKI5
HLkToN8lN6CfYnzVwhC6iQPleSBYwBtLfyaGK3qlCDOijreDO/LlVvlKxFRe8SsS
9O5di2eIIg9/BwU8DJMf3gpxB3IdzBRvE+Z+7CsEA1LnX3pRMaU6giiFHtUUOaYM
P+Y/hZFqts+Spxwz/t5nNvSnUg7DTdjQulLFv2vgk7IvQZHszC+5p2Gnx2XdyhY7
nYfTCru1ya/cZzwEt7eLvjUuU1Q0DGIt8GyhOs7HWQKE3o6BOh3Ns3OYzLqzGWbH
lfPhegrQjsIuplNhCX6+AEEV94qClR+6i1NqtTaJZprEcviSvRTE8SMZZKrHzRSv
S7eQxTo8hWVO2/O+Btyhx5k/oOqjdx+5QZpU6Cv+QiGBPcPVXDKA+0hGqTvGlfRr
peoj4akSlmQhCoGEo2G3Nw3skucDoPPOLDzwxPJPpxXVIkwilAvw/qJS9k1rrmWl
mn9YgTIYwJAejMj9rFtoqAG2HeZXOkVrXI85BnYSnJIlYjnoVySgStSBCAY7Q25o
sQKjmljGkmUDZ5r6TPmTW3D70nutUUOuFnWJTrQFB5/No4uhrAcPKISozME0+VbT
GKPHeoywkSS6pRw5vn+o6S7uc5Jp0Sm3QtwULlBxr3ACJ9ed9iqodp3MiF7rF49U
7e96rpSELJFcnPw6R0VJXCj6sSa9SWpy9Nf8Kp31olYB2YEglCsjzoE2/MKC8+MV
N5KkiZuBJGUGzJfi0ksj9WtPArtmn8T2rwySVxcjzR5Bxyf+dhHwAYumuwkuZ7iH
7UnVsTrCc1/3mZWAAiai6XeSh3q/HvM19BJKrjdS4B7GGKosBFhUFhAV6GtKUQlj
NVF1Lgr8VWsmMVWhGtjRbUi2osElL6adjz+vFwT624xGon5s8TxNY8613tI8uB3u
OIvoo/L/TUaw+LcqqGCng28plgz/HSeuk88AGVpBmIOluhVPVRdXIJrKtFGmlyNz
pqKGv0YRldf03jRu4g/KeybkFO07OoIaDDNmBmMub1VZTLQlul1ebJRRLf7anTp8
bwitO3r4GhHCmcSBbX5qZb//Rchu79rS19LOjXzk8PfhoBGG+HdZgv13DZgZxV6h
V6LzQcW33FK4xMncnrVK69yUMQ4bsJjSNOdHT6b4rzsXYJhw9K62LzVWjxJG39Fm
pRKVDHFw711ixDlbmoE7CmLq9ny3+I0ZXtI6F7TgKTXd11sVs8Pwu9j82jIkpMqL
BVvFdkhEFvPS7+n1e1khY8JfA/MF3NYgFlLFdaDruz1Q9Q5Ry0p6BlMlBLUS/VcE
9xJUzudNYM1pIH4fqxiENGEcFmu+yRWKxWGk7OSD1mdTsi+++emjsrgcIH6Yzpfx
X8hTo4PrOfWUpC7hjjoDvOjTSvZ+vsC5K9s9/TnuciiKh1EbR/rx/QpSoeO1Kp5b
8yNSV08rvZLnDYbi5ZRVeGmcn0Kyc0O5VWJLAM4Sp97pI+Tr6FK/0ctZYGb66cgK
kIGH2Kqq8yu1c7AQkqi+AY2ZRatuIzTrOwGG6ZVK3NsATuasYJVHoUP/fYmykIP3
neluzxBqZzUo+DpyVTOGth89Ycvp+6iP7WSjRoP7uB4yAH7jroKinb86Z0J9ghiu
PXfaC7XH3GceQuTmlGFW6YOa8kv2sTGa3SN82sCFZ9cuP/zSoneLHcFCSMpPj+5q
AUj81D7+Tt82QoNFVi4pDXRcRmviP+Njzat3S3qoMID2j0DIs/nn8y1JSNaRFKwd
sG1vzbq+hmCytPph3s1Cy4+3tA/d/A/ncVwvptomZuv4h9hk0zBKeT23DVusFUzt
lYyPl2GMwYiZNI0DGbFufeSHamaBj2JyOm2Dh4o7pi9iMDozrM8hDsFqXGbvhI3r
Ole7+GdG8WV7VkhkPOJb8SGNuv8XM8T8Z2yAI3SazoxgRojKywNqeQUCjotduL03
s5FV8xwrQWTZ44E3FtOHsZpGqxEB/R/GCxAEN2Lj1iyqzrtmbCTJUPZzrirX5UrY
0/i73WcoJACL3X5cjjCgAB0Il7tyCIb9Q/XwTNtgLOrrYyOhEv3Bg75K3HZ+GbIv
DILnXsLe0lUVO8AoKtVR/4z4FyryEy2a1PT3YpEdArRwYMNEs4jMLec70Q3Vv+rJ
Y3EBBJsWahUX0+rUxSqjj/lQ1rb+/TaQIl2VMNT1cT2StIn/mpP7Bqa+vvEdy8Oq
GUaNGXeIrpbJrv0nuax6vwpyWfr8cEkREu/3QrzjAqUoRXzkzfe1klvM8vaXLP+0
Ba2dBM/ERjnDxXJyizGOD7ptJRG9YVyW2JQrX+0D+Z7AUR5hgy7R4sgbqXJXmwZO
KpbC8i0eh/TvY5WDBvYmLAy2bFsCNOOKY9Tb3l60iZ3pdVVZ4yTH6CyJ0XA2VHGT
FfTRcR/DaIbuiRZdw8s2+OyOQa5SZmf2rZZPuh2LPHEqAvF8oM1dA3z1ROQ3F1Wo
ZpdrlC35kHX4uTtKmU51tE84HY6DAWvELp+kP2uCXv6uGqD0aXvFJTPtVXibHXyP
Acpv7d5P8BjmE51q8VT04FqW8Z0gr5tMULlcuIBfk4bae9oWrENxCzetmdw4nCdA
n2etFo4orvApnZ1buIQPEBibV5GYsxFm37GBq5sSYJlDEDTdJN6CJ6TY68AY/ZSM
BUYGLeoPlZ8Lo1OsxQOYw8LealquyzGYZtku90eKYHMNCNLoENifpZguzg83DXf8
9TqFSIkiSoMYHKPUtw3+9YCjPW4gaXoaLPxE/bfSG/QBCNW7i6lwEwLxChBEq4Vl
4ixBXQ/Jqh0mzjkGki/1AX+qsLJezu8Lu83wbhodpfSItcfeFQWlv7BnSbSQkbMp
FvkZaSJpFA1LRhG/wDKxtvgbbDd4Sxv8H/KvH9V6RiTUE+d4A9v/EHTV/mltwN1Y
TUgDr7ZYW88OaIyYciCcH+3N0lSXFJ6WDPtdlza1KKPxr6/wdbXbzoxAkV8fnRdA
2j+PhpdhaKAQDu5zfV0QLCfpTMXYgFTshHCszqyDFDKSE6Z9pADg8kyx+g8H5by5
vRGVFZSvoV18Pt+8kW1zMk14kXpvNblsX7aWWt0UOchGXd4FueVSlOGs/+TgEqRo
PaeqttIt2FSLcolPAYK8qHMk+KCktAiMwutqGh45B+qAC/SiasTX7r+kHAM4kgdx
mHnyvkLO0S9uldEU40mPVrkOzAlfk7VBffdjPFOF5bgZGSr5uSEQxPoRDrSm5C0b
TWQ+md+wC2LTvs5tTfHJCNzm56RMyQ4gWYdZ1GETW3CSOQRMJ+wHvjAJBXU9+29U
jQnvP6dNxZOyKsdEZlEu/9vc9ct4s5TMoxk7dV/1FAH+wBjUd48xQgveBL0+VCT0
8iTdricmpp3AG71tdXd9DRiVG3JcDGrjWiI9YN3wG2+6AephJTmyzuMfZBAN8dRo
QY2Xf88s00udBhK1cdNyjCC2i8skVsbErHaIxf13EWDzq+y+QxyjhYcVWp+xyuPK
+mincyzQZuLIosWCdR4XO9kn8OiT2C6WfZq6c+qGabXGpzbtoMPdeBIGVF8wPmOP
3fo50Bsz+o7pEPMLiILhnLasHm3Rf/xOKULAJ/4ESM9+qruAbsrh9J+clxt1f2UL
uH2mugz5v/V1Bq3sh/fK22JV440eijiy4dDFCDpyRwkRMMVAS0NQf5QIe7YEPpKF
3NUBsHGl9IHUwvx1MkiSZj1dfByVHor6wqhH/f0E1ziDtjtJN6PwEDcJBd41ss+/
PdF56qsKQc6tROJCPCacxYnEGiueJuGoCzR/puiJbipGXcOTT9uZfGFYIuZY4Sfb
oSH8YRG2MFfZ4TQWgVkWScIimHCbfXIewvf0iuLwN5aXlTlQjKlPYCF8nlZmWkZd
4zK6GTEdcZ26rXERfKdRuH0j42n86oDHr3rFlhBiFX2w3n/ksMsq6takp0B2DJrp
cmPkOqQ7HXQ/Lg8AqFtLRolHXmYurko/FJUbIRRGztNdrkUSspXq8GGrnBplSUWI
ujycABmY3Jb9TvMpXDyvaxLIP2CiyfPb9Z4mat+nAB0brhtVoj7fzn7H4uUBF0se
gzo4Zu3DQrGVziIbHLtivemoYgEAmGORjH4bN9wYo+cdMS2aPj4IkidnbgL1oOJW
g8ILhJ0pqbOkP1x20ikPKA44ZdDUT2Y6ek5L2tYBR3hDloSpXaj79f5UY/QnJzof
lH59+NcyqbrVVqW7fYX7WDfxdhpwzZvdICvm6b2OTKeSIZhUrzuxrUEt78rMLDxW
dvxMoV3ioaBD8vKLYVpqChBGWM4DcJK53hTMJOjTC1t8UKhZp2/gqJXfqehvnk7E
d7toi4kiIj97XdraSSH7YZBg9HXSdgTTQVCqNkbZ9YzOh1K59HcNq+1RJLFmHx6u
V/bIL3OU4SOjSGsx7GRrl60fxCV8weQLpGaPEAgRQ+2+lbxS7wphjAbe4sfyKCfS
H9XwokXudkqhwljdZ+dWh6icrI/lp7G4uU5Zdrr2MyQVFZBa3hLeYWuHqWoP7vcS
amXxtUSDi4a4xBxbNL+5pwfQUQYybxVqvdPABjXZmAYmyEGzXuf6HR3YBA6YiKxk
LkK+f+Duye2H//JB+LnjBujYE8xGgpdvI+aeEWTLJxOe6MbBDazSjJttoDAMmgpg
okzP+POq98Ej+cFwZowmG0sHwJy9ARIHeTsPXABDMgAPfjzv79sGTMi4mxmZe661
Mgmr2E+INuvT4bPJ6XYGs+oAuAaDbVJXLfft13v51ii3emfRY6qwJyp1hlGEnBV3
ki4aV9vTsJbcAb/E9XgImpbUrNiRfRipDmQiTM1zYgGse1VoYyBt12N+QrNfKk+2
390LxjXy603Sp4yl+legWs4Xn/puRaIex/B66MktbyHSS/I0WWYKg2fNw83/XPjd
UZ7eGVJoxsiGWNlXaAVf+EYFv4Q2uL7wrOwIuebI7Svd8O/WYHXepXE51g5/3x/S
WtKL3Si/d8I6cwKQYPKbMD5j6QCpgEw23qg3Oquf+6XgGxe5QLywTWMVVEHXqhxZ
PQkYEGxakJctoc+33Oqi0bvX8ck+ggN5JtaPxrEH4q0OaTdGdMJWjSTqvWVrZ+Ns
h9hx9zMAcXeo24pQRJi8x62A0h/1ggQWZaMBx9Fwb243bPQ0zE4Sd6Wmu1dZwAjp
L0QOa0Zw8zjm09Q2sfIuoGCUiI8734Ems3sLbejdJd6oHmN+8hrOmZJ98kYLL3YV
BcUWEcWb42jBPOQQlyLh6eEeu18f/WF9z+Tt5vw9miW1FyZ2nm6Su0UJnO+mCD1f
tBd1DYLRRXgPDHIsOMI4eb7F81h9br2mvIqPagzRDFM8CEgvABbwq0HFFtJ3aA/q
UfIv+Y1SgvK5Dwr2w6pZT2OnQOEod5OV1cVYtWWT3z9c1Yo4iqfClR4P6J82rU9V
cBx2ulYYxv5GYJL71IU5b9vVus6dwIvy+hcKz8tDzaLR40bA2uSq+xvRnkviXTCd
3+LZA1k3O58N75tZ/9h1zLwKhoKmqEdKqhfdaxlCpExmn7WqtmQjoJRUIQdOyIPm
UD7UQ/ff9fMqSIxetpnxWu2mIULC09WSS45tQu0wXbAMEyy3hvrkvmdatrXFcAp4
B4leATn9VAMFtzx5iwiKRdYWUrFl4E7aKcfIXYy83BTuMEyKTuYlwig/8rj9btMO
QJhZVgczCIKOu/oAF96pnNiQLFvB3M4MjzaRwyugvTAtPrpx+z0j9TivYXbj3ZTJ
/K3rBet38gmyCMD7dYNfbPQazKpiNFY8ZpyJcr29GmUSAiqPOLrXjiNJvEPP4G6M
2ANHZzV7p7ReXCBbuibKsDYP/4Cs/RKmungXAihI+PAfkaxIPS9xLAq8c1VCmsQr
9ieVz1XjKU5nOjLcSfXQWMuFK1PO1R+6ze0uIPjGhTeIL84zTN5bHoVVdfwjql05
WDb0t8UMHq+z72v8E5QfWXzYVOF4o+BAwgsS3PHBRS/7617domX3/GUcwB6BT+Et
ntkB4vVsSxA7wMHFyTLKdPQrzkPZMv7AQ/oOD8pO4G/eO2xQmU12BTJIojZUAKbm
2/RGIdA8oERigJziCvVMEACMg8Eo0G8xP3Xr6t2aq8VraJb30C7vGNF7hjWSe58j
aLLRpoH3fEzji7++8gL2Xu6VvAVWkWsuFh+CZMIZuSIq//dTOC02Nc8lF0Wk2GpB
d4RqdyGo9Jo+PczWFehrZl8OupUgMMXknT5wC211F4i9P/On+DT5416ZxL/wWyeA
hXhUtOc9UrWNnrGNOsBforH1CA2m2+Fncq45aZPlOOfBcDwoUwhfCu7TAC7k5l37
+s+LAopp6261SRRVPh7X3m8n9TZDRPS5vxNx4MrL9X2IUM/JH+3N4CFKnc7R9uoK
bXswRmXaFj3LkNBn7wYANxg6p4Q3eq/yLvIv2ShlOkwQ9Hrtuks6NoA8Me+o+43p
rxPwTmneG0NsjFadvo9fJhUVPq1AdRCTJd/LkuxXBdk3Vk5laOCVtkjaFI4MBQqe
6GeKeYCUsHw1kdgx6MhNDLhNEyoCEMpm2RcfD+R7e+KwG6grgxtmgqNS06tWrNvC
Na0MZ9ETrAzVjiwDRN/iWOHd1eawZWM0ofF75DtEFn8xsT4S5vRDiwOGVYCl7w0T
ziz5FHGlzRxxGJIfABo6S4fA0XhFqRHfwF6USLtbXm+6iF4JIRGFlHfT60fspmyQ
Dtn6rn+q9saDndUMT/vh75oPpL6gb4jnr4LNOcbfCK/O7lsEfP75RUejYEygLxeC
jiRSN90FC+4uo3RVRrLNJ/7bQCQSpBxzxSQWVcEK7PX8TZQKWLyMfqQIX/UPxiBS
/0i93jxW5O/urZ0woJxmfBkCAkix5hEa/m7cFX0f1Mqz3F4b9xnU9/dA9m9bRBQ8
0LuBa6qH3yj31l47Y/Tbf3ZM3EtxYYb/a1Ywj49/SH3llvjTYhgnqflh0PqwzmW2
NV6vlmxhGP+R2a5er4DRy/z+edIUd3FwNwgUV0zRl5aIfgBP9AHnsCvIXmlHb2HZ
42Emf0q2KTYhshVNt9+5sp4FW+78qQ0w5BWnlB/kB9mm7rZlCnL2Ey2eS1y+IzWQ
mp+MhCUxj4NeVFaVOav/Oxn9PfyOUi61yeaiw1T93xR1w6H0nfPdUFl0YgMfmeEY
ted0Q2hFFjXE/GDqHhIX/R7K5iOlEXy6xaC69WRkvA2HM1YYtRHPfQtRdt7iBcz8
PVFGBPYE2jyCXiNddJTDRuMALJ38zllttMJ/Ulvei+lBJGgxWfbaRR51SOi4nrq1
jb8JlxDZKexCIIzdwtU62oHlX8F/B1G2ciSucMWZFpdpr8Qsax26AtzyM/moYier
xttX+G+u2SwlUZDqnZKkGsJ4qcGlSwt5IObivPF9/U4kBCWiVjp/yXiDkmygYmXH
j61aciIp24WEMl7xZHHHKtfEWblHEaiAKUkea5gerYxkZiKOf/YHO8GMoJkXUOvc
/rxKt5KzgHGEDDCaYp24W2NC+URC8wBqSA/yHCu2MQlerunmcyjfQtbHuIndhyfE
PpUuIFlLMiFDPDI3IGkQIstcaaITzxzdmvjnzg4qF6Cw60xUjmnPmbtt+fcgZU/8
rvpn9zgwBifcauzjuhDOUN8XKA2xxQAW1iCC3UQZUIMbtuCqC5iiZ1LJpOJpbTtT
Dkow0xmooyB41nP7NSgJHnKl5B7t4+ss7p+3O79CekNKwGewPKUi+v3D8sAq9ryH
uraSqgCJyDjf9+kQbqEY6jETlONbdhIWVH/YNW9N/5xghjsozzse2Gt45vv6I1sx
k0sVwBwWa+Tc33twXeBvjUNYlPjfMZkty9+3YnEVWcgUULL2+Hc8AWXwF3UDYkDf
PonpHlrgi1krEnyEYg+5afoJ8g1Kl3wwB3oZvNR76v1g8zsL6JqVMd4218EQpU5O
KIvQFC1FNJrv5xT5hDsLzSzMdSKJ63SlOd9FNErhfPRYm/DokUBL49YGTQYy4iyg
F4NqWIBqQiQodoX/njJW6YwEvZWHCdG4Jw+lSDUyOrxy+as199MEa8y9TFBuCx3m
XPOEnJxNvzT5eMjaFh6hbVsFS1MPIRfzjzDb2JyixM06s191B4KjVn4XHiKU8dC0
Auju6xJjT05+D+ymnXp7oaBolZyafBr+7PmeE+eTwg7fH5sRavJKwDp03d0hwhhO
0pS5K5lhlMTMRmh5HcC2xGersxlfV0CzYQ7hnH3chcg8nO4M8K9I8p6NsQtV+rtN
uW8FWciR3Q2OpR+YHfOpDZLIrPCGoBrOQOb/6QfrNLwZO2siBM2TVXTd7McPm9de
LrqcYUbdzagV+P026uVEsF6SA91ZrwiNz77BEK/4rM0+zD8zLoFtcCQOhId4H7if
0y5KtPdM1rG8xLlYBQAHRGXJFUIvX2JHlI/zHBzmERA12/E8SVhPL/ejorqsyLtn
9pIeunJ7YaNIAshAfUimgfmumBB5NDQT0S+6cnnRcx01cen2hjiPmT8CG/jFpo8F
GPTBqAAIaoqlzIB8E30DAxN4vYq7+cMmxBP1+k487CIml/Jwapy+E9b+OJIOhqD+
A0/DAxVM+ieYb+GeZKfG+dfK5Yxzkrlwbar0rlvz0RrCvjajg6kMPIKgk2XU2xKp
LHh5UhH1+D+de9iane9NXCOxh7hxsD9tLErGn+gOdPi3Na2GJTct6ytCcXGYpXeN
fYsmZnTORta5dPscXtXtCR2NAZ0zC0vaX64qUi5qNLzlDMQInT5pgpqPt2KHPk96
kBnpuw1KtBFzf1kffX7QssyQDRFCjw0PeIUC1e/KZ3/AtdPeyB/0pLDmTg9WOvPS
SPTBc8xIkDKI/xxgU7vLRY0uMFb+be3FaCZmqtoMR+ZrCnaXo9/HdaLyiFxPxyrj
YCSFCthiffNEgJPh6l24qVMqWVGP8lGkLAMN/Z3QsCDRZyZwsudqFOkStEXtYA79
ivIWYdFJn60r9V4F7xsmRX/YPipiTCXnbhcUqVSgtn3eZuYZ19kAESKkjlSrrRRw
xaNo8qKkIcf+SOoT+Nu/1W8x/sXG7Z+1pcqsh8DE4k8U5SJhWgNUONcLzswPub03
0JGas9n5WCKssRdkrzz6NXRM6fRckVcdonhePsIpldFTmeZgzPm6cC0hWXobZJ5C
hK8oCcHXTSbzzRZDF7nX3JKOSxvS89/g7sZSXf1wL/n9nKFi65VCyzOyEhTNUUOw
N7Ngv/0jiNi0Y3nNMegLEG7SXAyW2QpK0SIqw9N7XQjzNrHiILwrkEVKYosa8Psy
v+NotFtl3NKxys5wnEhrjy4msTFewLBSpKT60BDZC9YTG1NxbIQbaqKKWpqHijSl
uVCuF0OHfDMaLtnt62hnca3dN52QebQFlzzflc4GIqA4WzY9QMvnczPE6ve2KZ2I
p+yISeCO9+8ZS//Q++/iB9/Z2EZscLhjR01kafiOz60mLjhZYFj2nAcdHzwW8b/G
k3qXdXtAH9WtgEdWqLT18N5TlLFVN68CcuzDTRhI1V7mREcjxNMi9OZrjVgLQnAU
ol1qqbpMVcx1aPiCRvXoOKylQccA9OF+qWfq88F9SO9W43Ud/OoSoxq88bXogt8y
eMw96pXjyN8/l8YVWHEK6ROKSxs9B1P7aqChuw3Yf7+nNcADvwlibDM7PghJZr+W
w9n9Uc0ZzFXZZXtfi8RH2agIyQL6+F29hr7YizDrJL2ETJhR/TqhbF0HboWX+edV
T8cuNFlJuQcSPWAyMZfGeQD+S03gGQU5ISqzD21J0TUN4sj5peIA9oEhXALTX5GI
TxmFdXUMT9WPSmp+vUSKC/KqF7c1DIY9oZtDuNa46vg2Db2ThmcYvxPVw10ZtpMB
79F+qBLYx1C8lBpdoZejEExW9rJLM26CVPQM8epWzofpAOqh1xjF0vWzUXIEmQTC
94qQZBo5pTuC+NWzW+NL9BJ6VIffOy759c/iawsCO212DHMTg+ELu4bWEvRCtXNQ
9shHDXczRi4H3DqGuyb0eDCqlpWN2xmYKTqPAVr58GXYYjRpl9EMZQomXCtnUVoP
AdqhL8apWOA/Zziufm0Bkc6bi493acR3aj1DJ64Mef6VrVvOxaTx8euhVHzA7ytr
Dtn2ZxtNdB7I/dUs1KkTQ5uodotM7yt18kfCEIEEo1ZHIUdrqHZwBam+ABjC+EMz
dpySEEsMSfkjSWzyz/3jBYWhd4cQtp4jOkxrpN91BKhpUW5GHtOr4b56OP0AEH4E
YmZIam882LpHTWpl22omv38Gp2+3YV/JhW97LtIe0MgUvx3NR2/wqkUGmVhIvIKG
4198NSjjGb6exuST/IbKYejk3cBAEAo2D6fdOp8qfgAeMRY0QZbkp6actP33uY2h
QvtZOclofYzBkuFzDdrHm2Pe+w7MqOEJTjEF5iZItoygt3F3rmNJlRBPUmf3ZrPR
NFEyerlOhFldZT7VsLe6wfFoIrbk2P2rf3PzAEDz5qDTsOVHHc91kqetr4ubH4JL
xbbXoukvVfcWmO1rkCBffQgvuhe69av7Ff3A7Kjo6wbK9pRRpSjmOjSKEMrUwhkp
9GRfyxGaqnikfLRPmr0+1Xiq5+/aC0o20DCbq/4DE2b5i2GsWyNqS16S2FB8iWKv
2DSHQ1g2UMeUjca4pBf7tjJcAoZOtVfdn05exQjZAi3rvX0hXdDdPX0e2aAtTpVq
KKKup4sjRjl2f3s10XVzY+zqmTJuvD/cm7OlaXXmVX+hmt3bFMdlMGzlO4BdLl4m
+tfbMCWfazput/KWUwcaHEmqRcsjkVbuveMqDDXZMBIceLwptrMTFs85P19X45OP
p4fqsTmANk74pWSkocmIzs8LHwWfj5o2GxVJm3MZ+KplvDrIa3x3pvtCqno+Ya5o
K6K4856YwG3EikbG8qjuWvdx6HhswlQQc/e3qHlWaO4Mk9e6Cje2kMxcxavLa+w0
WbDi0dmMAde3rmgOUDe6sNdOnwASI6+m5xoJwVxuLKCtMAXKPMet69ze4vSSb0B3
mwHghCGUpKmXLEUwDSDqZ5nK34rifCVXcv2herMVLc4pnrqGowS9C2XGbCSR2VKE
SrHBTiT/yQ1g+dcqq9ZmXKIE377s63eIol4bXhHhFKfcDtRBBbbtYu/jZr9SAZL2
5t5HISksE9h5Jkdf1LTKJ7oEk6XLDuIvLrFf0vrSHFXfVAVmpDuiPBGICiNXoZIW
iGSy79EcZA78DPaBQ48VIgRQa5i4WKM62jzQSBpQCw6ujBOX1mcAB4PHcq4W6JR6
OzB8Kh6WYlYdd42yeXikFRDSrGhhgQg+I6A6KM/1fNKlY2KCbi8DeVGSdTR/+Kt0
9C1uom+mpOxXYSg3ez1jWsGbIUZOKQ0KOH+fuVvghxkn4RlsyEVd4+85Tfo/KJmb
z2AL9dtVfc69NOwmQoFI6hdqSW5CP/X/PkJVTBvx8i9FIZbh6bl4K/HjBVWEuIRP
WVo4iA29qy58zSechb8kGam2e4uQyQi/c23uOE7HVgWgz0m7J6xxE7Ec2BF9NKS8
6smND59IcIoOApR/kcvbHjIgqRN/XsmX1U0EQw/enuHSI/SUusaadBq9OcWJqTFL
T7tU1qPFu1x+rBv4EOgh0AUVfYAljB4VusWm6n+PqZN5kV9rvVsGqRp3VS5ul5zI
cal/J21JX9ZcHgDsozy1TGjKleAMe8xR0dBFHou2/O4JSzr/6KzgklWORGSADpeD
9+y+5lTt/Y9F42B260Jvo+7pzKhtxM2r7ZEklVOuhZeyyvYLKlC6DhjRiLbuEecU
qz1bVjPXuUi2KStLyHOgVNGoKiMluTLgvAoJ1wdoj2yyaFYa2QYykzqJ/nRUmOAr
arGuN4FMAOEoitFa9aysyz7wQxhlhSV4cpy0WWOB22dVHdVba3aOXAmOt2SVXEh8
932Rc/xrHUq8Mx2tquPIhytxt8Q6BxYPFbIofGPxnCScpWfLJahzDasB9BkkhoY1
aR0jskB5mZjmHk4+RQcYW2AsqoCFaOkaIWHi+Wl6WeNU7s03Inwug/CdlEcJqyV2
qYhI+y4BUnJkjaItxS7YSMVrOaerZdWgBqXbKmO+2wkvcVJflufrGNdsP09H5COq
PQpf4Pif6JD+PNAAWADOHUX/5I+wFAXXD+juyqr5xe1PcATpkcpefV3ZqRCQoFrY
uitqkC7q0IdA6JJP9LvMSnzJ7EDwiNqI4YftYPIU2rtJALzVNbmOIYVckP9SuiUb
uK6mwgp2ODLSagWYc/uOo9xuIClxrQArRgee2lkVw6kfpUuKQ16YMLvUmeb/heKc
WtX2d4VtPVfXCp9aqtKF/1/uvXz+mCqlMDVR74wKLS5XwgsNti9tvjGiv0jIAkJ4
PP03RqF4pDxmZRhktR/3umhD2I1PJ5qTb4DWmidy4eoSEY8Wmg2NisMgCexiTyuk
6dQO2gFi0RBtne8/UyM87UDhNdL83KHCcoJGVe1Xr1cq6yRjjADqbpg0C4bVdZi7
wK5zATnuhigzPGgzGE6gtqNA6ustJ/EDcY7Y47Zi4NSNI769qLeSMzSEq657Tiib
f+99aGKgpUG/h1KPOVXSlFb2805+jXuc8q213gCuMYU3Wih2slfIVFcT5HrbBU4W
fJT/Agbq7FyeT4AE+b2+j0tHSNo6C1k1joPyh9pim5IQVr2kKdgnm1hs8eCV5tRO
d9jKX6/rGWOg3n/ljE6NTpQFcyRQ5qMosron1YWhhrbBx7a8n4oxfpTi18Z2RQfC
rA36pUFnPR69KGeNsD3i+ugpD8jfcryxCxK3f5qWIitYLY3R+6vhDfzWy3KkO7jk
6sMtLQAksgsB1JEapGz/4qfNcXI2CSNDSVPQpSm3ReNStvEjRdUFpm7DgtEa3kiR
PeNoXCDz+8ZxA2c0qGBa5u16IckNHYMhA+2g0xLv47STy7g/Y6hb6oO+R7m4P4MR
ypmrkPWnAGGomQWxgzv2iDjI/rqA7JUqxq/W2cX19QdMkX/rfszeCoYfyTn6FZOi
6agxKEztdcHMmoEPeUTOrww+hGA37WNNwAcMJ0m7sdaeDbQECfg2hp4qss7kf6Ia
Rn/0/u2FGZxOL3whIF3Lop4kh6hjrW0JyteQEkuTKXrAtq0ZHXrccd9QmC94jks8
pfBnz4tSj2ktbrfymZMviR6kL0N4+lmdnBsde399WopMTGzHfqDUGnTlU7T/pVbF
cUts3ivS2uW2uDGHyzOy9FrrsXBlrBW1VuBpLETDU3yHRpmSi9GnxtOMw0PzKWnj
1vYXI0G0OYWNApdy8U5VMoEfMKy+firDgs3j0t7EQoSU4sMWRsQsoemGFGM6y8t7
0warTPAFtyiPWqPrBapE3vKVk1uxtVkOh1o5VfHCdPD+uOZL/y1eHy2f/VyVAFPs
UetDQRdGnsCWbBQx+dLL3T+xB6mzlMkBxx8LeuLP3HPEvw1poJmWbKrI+0/QuruJ
HUdfVa4UDmKt7tOjrPtWwaEWSbiqPQUTG1RpwLZS9NLPsIAqTp63OtFpNT3pUUo9
fzUQ6YVgBhBQqucRtJot5zNAD+/50ry4JU4nZjEY0AX2sYZbwxuz6BDhm/IFjI61
elUKB/54tepLF/mIofMHlcZlhDsxkRalSbR9t5m7+XohEXB7mxfvr4EnLN5vMmGl
KToUWs9PfN6XAjWnG5Y7sulR8/v+VUCGCDYghVu9x1O2+Q+kQKSWAfyyuSvZehRo
BLE++m08Oa2YGdKBH3iEMcJWfHFydmITOkixpCHhPu4pXzLY9nTXH/80frOwJaxU
L54I/Y3dcN0F77zmMihA4W4SdceiO2rwq9n6aNN1cnIUEb0ywxZ41mBUPD4FZA/d
x3reEp2wdwmWV8C7aBVyZcaKnldVDHtsOApwGxN0xqqxswqtMjNU6DCUpavPHXDu
xmTMVnVsePLlwDQrq1L6h39AQBJUMScGXRC/xouc5RlhFhab+cmA3KQYd457Ys8o
0es2ze6HOt/drmyXyBC9AvUSpZriYaf5wBpDW+QOK2Km6HaJte5lXa9DQUQ9j3WS
rRarB6NdOCe7GY5Z88+bbLpJ7hgFfZW0E6oQmJAfO0CEVRqIs+i7chtaZZ35WDim
+i4QNhs38T//Tc2sOLUoU1O3h3r/H/bwhxUnKS7hmTaFTAPI4fTC/5VhN/RwSHrv
WE9rubyQUwtLVCKhslJOiYPXulmAee+ppFyd0lVsX7WJ4gnOCKwzVQBxzdtR58bY
RwRXb0s26nWKzzimk96YDC9i18ufgMoeP/fmRmJ3IaOTTRH/ndaWwMxme0Gs0EHX
jHCg6kxmSe42xDFTvoBoWdHSYH/U4qD4WD8Q/G/feaRN7iQQU+/Cwsu7ZXIK1v86
y/NDZWy55/vy0h+X/5J6uM9TDIiwZcclkTwUWLD3iJR/FMiBWIBspaL2q4PdH0du
fYaiUzzmlgtWuUXFa4Y47rC7Me21iNOreBXIwr2UvnzDcs00zqyTmVOLYceOB4wd
11FEfPTp92cF3GrkxLXTyIjNCeW5TOFyeziMy5IQCm+qb8KPRaSWLxU8fPRy2O5p
dvlPFf9edBl5SMrYzAbHTfOyDjIobFapeGT8sm5D/vlTkhuXluoYPLVoImWdsF5Q
2+tL+PfMfA3M8PsG4d6Elc5aizBeUmulCHMf3jra6zNQ5QIR4H5yy/dY4FpY9vsB
0iV76so0++P6YaIdWCx4J3Eh6rCENy4dmIHGz3lthWiAhnolYGNG2O+FKzPTvGzY
WPRRWT6l8S11AEznNoYBgk2aOYFVgXxTZJVTkrWrZj2mogP94fAC8c8NSOZjM3+t
m0ZI0CCWKsjf0qenfaWd1VT3rBm3rSuAsfep/LvC0tox0HCxQzash8it/TAwg9xV
+I5vdKy4DlK9m0Rri6Ah1e1FUZ5ABVvjA0k4M9ZBi8PSI/C5CmSg5IScVium19HV
KVrZxK+SOJRZDh9J7drm415S1LSrkRNd/4kFNfx6KwVl7aZy0+vG42iGOiQVC7Ng
QGC1b+XKmaNLxuiowzhUDJt2qk/eYTbDC2m5oQbpYX4MIGPMMSPg1v3anRTo3RbG
qo4u5XwqFkVCeqL9LaQbJx9r/snYJgvvvwNwM9ZYXbt/VGYmBWGSzV8mLVQ7YVDx
pexpfkUL8/CrqZrLVzNXNIXQz9EiLJPZuuMj/Di+o/T/VxYj3i4y+3IYd9TimIsz
gxQufDd1DLaoKaAUDfkyHKMIpREjnFONqMKbJAoGw5/4tlfetjk1XsK4qjoJknfH
avc3P+sVPeUMLdTWmdQFW4yduuqVg3JCInu6CK+SQH4ppmBPH3P4EUsPbnQSoHZF
RUJz9vcLLi4ogomUCKzKP6xqvQMRDbKWrTwwBdFsc38lNWFmLTewrp2H9vi1Txxn
STszahlzIfhgC9kDpuReyix1KtFzrBNKEbyC0VLQaJkY8/SbRQ4nBk1IlPVEOakX
wybtTNgb8lx5weGfYRWwK+/XkgxVD4RXS4o+VGRW9gs2lEXZ/TZjp2MmScIWRJMD
5zZ/OYqdUlYahhmyRjNLPekFMDxK5zJU5vWI+JQZvEinJLmIoxEAyYtijBLwjzAe
LaRowx4d0QfWyezZNw1XGejnpsvzpM38d1UkCnHxuuunJFCYMffiN1J9O/Z+/RJZ
TWQvtiuxCchi194RmvS+Atll4QtkhNncRq53e6fwrdndnK7KmK88KxQ3X3V204FR
n2jm67ZusIGw5CIh1Sr2OPtX1VDcjg7FLuVeYbT/0OYZeI/sj0nr2UZ9O9DozJ6a
m45DvUW88AnPTteYAfXwSie2/IP4kgI14oEd/rqr3RTYQGMXWPhhTqF3Wh3c2DS8
RWUyRtWI+8k8dk4AWIKzImP9Qoyc2Em7lFxR7lu7NoVMXR2ZU99trRn+wDX2BPOa
Jpylox9/xLj/ShFhQmk7nbtm0SMCnSh6JT0TRBsnW3GkznYH1RkMhqjKqTxsuubs
XOkSsxy5xhfbQHyPNywH5kh1KG/7yMvmSyAL1Zkj4ce48MOVglXfmyYxfQ++eSlq
eHoovmDCypzekqLoVWIX9C8uCaC85qZa2/76Xrgo1ahPrbNh6jFuxkQhX8G3OIDl
TlMpng3WEq/7sAdGib3BgQh+9fBQ3knv9YMTQCwMfTiflRkP41tTBBkcVEsjj9Jj
n0lrLsTUsz0fHm/aKFdKq/jdc1KYcazrRYUlumHxEysVsIKegTdIQR2qY8fJs1cp
vXAbvRuf5+yVcI2uXRDtNx3B1Oc/TnYqJQzCuKayRg5HMqbV8xQWewayiEWAnnbg
PLgvRC8uLMd6BNl4OfilJ1FAFVEscihfUkk5lAU8rMdktwQcVI0TWybxveZ8pspN
epvAbYcnWEcc8S41MTNzn5R3A1K4FI0GMwK7NGiEshkJISXtamJMLZbtSjw03EjN
oFUis/cM4zfgqZ/pwMx4g8vKr/xs32G5GzTAtf6O2X3auQ0v61fBzUjzjGgqrnTW
s9T2o3ebQlkOVpD2nrwslxg6TTmgCKhwt8pPjvUrLCtAWPb/6XKjU5xuqRVR4v8R
lpdJHeOwqIrBYdB4x116DOjxfaDQ7q2mV6SP5JuAWhxrKDBuN1Sw3ArJpxEGseuh
8p3K4SQ9Z2ykwM1xWmYLuJCu2n8aTu9f3uCetkWfeMej5rLZXxNdgn5EdXqHCz/X
3SHNxNUiVQMDGCoCTj1CW/PD5mhxnbVmxJNLQgxb3h39ZgTNWCQjmcqOlVob+Ate
xRJugI9s8LgfDo+WFpAI9ADlTGlOTI1f0Z5FL2Ai336u98uvqPDMg8yhw0UNmPsc
LbLGTfaF/nMzl9aY0xKZYi/tD86eDNrXHIkYQACHkhUHXtSYljq7rD1SbJczaKLm
1eEWFvXgGI089nzT99SXKfK/2rFOByHwPHs7dBGOkNiHFbzkozCiB2yj4yL/F83x
K3XbQz5JO4ofq+YgKOVmMkkIe2zX5y9RBTGY0esniu9rN8vEoQgel1GhrbmpaOkZ
3A4o7yLhQydQth/psIgroAbyGRi/Y+GDxTbJ+mIWdHp3X88ry7meM8N3XMCNUamG
P7Aqc5cD8dyJnuwHpE75c8c0xLRD1S2DIIGa5V9F5fj+GQYF1McdnlBUBRZsofnl
HZOQaUCUy9FN+O7ghj6ZWUa5d6YJq/CCYXF120hDXuQ7h64UwM1RFKAfIdweH7kK
d+PHAewTnYtDPQt9ihaMpBuvlwVxS46gMO1pMz6gpv/0PilFf6wqVu5RttqcKwYB
hSbOqsHkCAMRhPJNgWl6phn4S8B2Z4sfNDiFzrcAvHCOfXqzb6mbliYkAfvh1/rf
0FwP/5j7yZkJNLMesOGZKl5mbUPpbkTEACjYsnd2q6zjBraRG6y2dLavLmomSZbH
vbabo3u0GEK+qExsIFdFqKF+n79G/Au4x+t8dRqc/uRSPpXbpXUEP8Gef7IG2Uj+
bHPgoTQJpWB1asM+Cb7sulwVxaWYJyguDd/RZ2/1N8A2blnvRtmeTm/2tg2rTHmC
SPa0K1sPU1Kq3A6oq+YWe2Sh6zhhuLGMHYSSS8ibOxeTxllntGgEKbVzxV/aD32/
t+wG/Uq8pHeu+o+DPGZApH7lSr0j6pRGanXMdaz2s4BoyogUS26ahU8HmsUVkr+k
j/7wqWOgMl0cQ81pbvvPwvSxYV8h6pz3gxQuPvW8I80sWztewDKb/SRGab5QrRFb
8XtRyuDXxpaMvqw7FVykWoLeRWVouQTYPWEfTsy/9U32pMgc/9/1rAS/Y/yuKiZY
LvebXN5JNfyCsG4PQAJ59r32/1FJphvkS2wf4jejpM6y971MQ7SgjbJzjE00VIxj
QbMC2Yru9p80ZIf1xJnQi1jQRf532/3fDSijLH7x4ld2KzMb3fDcu0dIoZWor8f+
GNkvgNUMZlL6Ufj3fRokCUl7ik1XaJCJyjneW/kyXewkLVkUQJqDWjTVSEDmOUQC
06djge7ROMvnjI95sD6LzR7uBikJzqyYpifYrfhys9KYK/fggDNzQPQWP8cJ7c+C
5lA7yV74PliiXd31WkFKJl960LXHOUNk/fXu6PhRwZvxch3vPEkX7pIMMsX/sumM
fdQQ+T4AkQ6KpTSZwhU9St2MA2MOQ6v8PI3tZnVwrJlq+qA+Ak26tVGILV++cig/
pckUECxFcuWrR7R+qlqum+QkP6/9HJm0OHHx4j041jvT3CxrzdLDhI46CNmHZCHB
Xt8HEtr56ZBkjXx0UI2m4c6/ZwFSs/TPsILlZJWO74/gRnPlJP4BOGrcw56wGYpS
HiUiUqFfYZ3lCWt81Zg4bkZL8iocmkUtrgWYmAZz5GnoXfPfE+sXx53P14FMw4J6
g4g/F/ghudjLvnOofgLMi5cxB/izLbLzoIoK2J7i4ssr6qP1cBQS4whIzC8LpfdO
e40m2EPJavJyQjfFFKrCI6gFud10/RrShzUhMAxmNHTVvoANKPGPUsk/agRJxndP
YcbJXXruX+AVrp1znXJe79L4a0dIdAiQ2fIwZH2hEjfJoamOkPJg9sRL7ArnPqH4
Hz/vaof/Z9kZveOasbBj2tEgUhnrRDlxYK92X5vwmODRidlM84Edh7huCSmyDCCk
MIDtpe+S94cUKuaWTc8F3NKI1h0O6DjkfRuAeXGffFDDlzBCj7hQjjez+WlAK9RB
034q2hceEgC+4FFVNI4kW2PMdrKh8Tb8jwW6NyTjDuRizu557e8rjH2cu1PMuI+L
tUe3jZywWAWBif4sBcwcZLQ8Yr4kQUdw6pdhkO3qYOxmJAcz+iOLPqjMxpaNc0o9
+1ZO/NNxrpV0bG1Yb/40294gpciJ3PUL99WdUggfD3zPKaDokE7AEwnErLc20FI4
NYUVh3AGWSTRggetL02VymcHZXwb8p7ezGmCs8/MbA3JPzsEklXeW0fMkAmBFMsa
IIfiCyM+THROPi1ZRFq4tbIcrlNzatC2TzTotUZXD1RMTDS/ujuDZwXUqk5LfNhO
hrwNi2XvIUmR+IHJaWkPVG/cQn7uCUEDU0PAFsvWjPZcjJBmlzjAt6lnvhCjoA8f
HekKg+44917kBLiYgHs7oqSvQyRJqRNNdMi7YGVXkqAfNFdbJwkr3fNGeSC4Pg8c
LbVAMtp8aAUtYpslrEH3RIaTj5gVyoopfZ8kQPm0NFH7CJ6W6VHFIryF2takAPJj
8HaylUqu48hmWL0QYUO4Sy3Vcl7vNSzFa/M2MNamMCFQjnzC6zEeHhO+H68U1fil
X++/5g0Qp6cbOkkeBjwCPKfuq1T6JPjFRWOvKJ3UQEtCqs21Q/1zFJFGcVau4/kX
lOy1EBiAWO/m4T3BNYzCV08GfP8C7yI+QNkII1yzPW2/UqlHviziQM6cHGjlU0rL
DsbwJUelQBIIUVKVdK/2lzbOPTuQsGe0WQBG6LjDQ27VZ343KJTyPFD/1zPnrJQ1
A78Irk+7oWv6S/EsRnjzoAThO4ktItkCqF3GT8sQLKpa6xLAenP3tz+kNF4xCzAt
sJMkDBjvbx55IwC1ooEcv+mJDM4sfy5W/LibLW63a9m3dOML4UDJm8J3aTQHd9wj
q6f60mx8Mvg8/SiUj8O5Ets6YDOH/+NjAANY+xPVHc0tYXFxu5c0XVcocKT6DkFg
1J30rV0PwaMiWEZV4E8vx25REc+rRqOkmtRTjNSD1vuoEwVelsW5fdvLHG3e1Wq9
PJ+uhbVxljcVy3zM97MWznTtQXlWXUUXi/Xc9Uc5gx9MT8AjA+4MZoAyH4514NSE
nnPgbc75fA2rhSjKmlCb+5HhtSE7K4mmXVhE5QttPu6N6vlOGNFMyS412SVjLSqd
NzXxnD2IpUfRvhyK7WO3lqNHj/cexVthuk5h7kpT6koCKnK4m49IKQEpPU3OSHwZ
qtafy8c0VcCNL8SEHS39aUvB4+WJOwthDArvl3mLiZ3U2YiJ8KEGhDu8z8Ds6Xfr
TsXT/BEqafEWZh7zFJh5p76UPgrlIibHvbsu8ZzdIAPDABbmci40fL/ccNjc8JbP
L/Ndf2+ioX6ai0UswG5WjTfRIWnIXEQa/A+adWI7XbX2CGm75YcEftP7gYFfnuAN
a94sjx+UVagSl3BDwd3JHqcB88Q/IDzIsXeGQKSSD/k+Y3vY/yXnaxqQScXGT1iN
Aw3l8ggfA10lDfdeEuN7v095H2YJjJSF5Ar0RYV1VEirWFJ+zp5lJ8w6PmIMNlsD
gEVzPP+sEzExInGTBJtn+7v/ffgBYEXu5OGjHJqn3j/Y9Clf9/YHGiq4QfFv2eya
tssEsclagQxANnmziljtBwUNCGFA5waxJfpV4DHItT1Ff23NM3N5Zqv0O2QUM4Bb
p3tzRCEFSxRPNr6kNnbMQmpl3WQ7zrUZ1PConBlsc48i+i4qaTVDz482/apZjYyr
IRSkoCri1oZLsLCiBbTFr1IE/uJuIAbyGAlULfhlqnZ6l4HQJcFo8WUnaqElBc3j
v3UAyDBds5yFHyv3UOEliQLDkw+8h9QEDRcGalUEANY9Y9bEpzi1bfHpP5ZVwmUl
TpE1e5mhkcjIdQaHgwby1wxJAJbHYnmGAtbBkVXueIq9DIiYhO6C3dEU+i/MuZl0
OrzN1NfC5Mm8zPwXexAMaWM9HtIZ/Wzbcn/ilqbJYuaSGetmMSiDexU4R0z0O3+u
stHOo8Xzu+YozglYqRlyLkaLmmbD2G6SY+aUzcMNPaC5DSzFJakdewfkGNJ/YnA2
MGzmno0+LfxSUAs6d2T3DhOVoZhG1m2/iUNP2h9LCPFUr9QoJue83nRI+505Vcb1
fh1F/Z8UDrJQ3J/UhEt34zmqMOOfrDapNr37/v0OyRXgqHePan24AJ8cXkqQ4Nce
bETIOgZCbn40gdL6mONa7jClEGgLRMtNccn6IlsIk9l4c+Mgtl+JuYAt7NpkthIg
VQ7wlxY5d4stHdSgnY1UAnhb+gEj2U/oJLPrFjNzujcljGYClOjU2aKNoLoJEHzr
b2elZS6nxPM+sdFpIiqT98EFtJqgxx5bu7UipFJ7oqM84Z2yQxVDEtM9hxW+YEko
YRYKhH5thXyqR43x0D05uCsjAM0Y+Ub19qh0ykgz0Th/pXnEnXH4XN9FJHUjaZdR
qFm0vciOtEmAMHTfvA/TTi2stBjQIjWXEmfwJEb0JkdtLCJozkHbWt1lPJaZy4iP
0/SUVhARnxl1IB8vAPyP2n1MIw/Rqc1Ac1/9RN5B8nJmQVwrHF0zKvXhy4spRvJ1
xaIngKMO5IRpxheZr77cM4pnpsreBp76nmGgWsXgGZKcU4uCM8ciDxSCAanGVXZy
pUI7h1/IvoWic2Vs+BrdXS0EtqSQiLcfAUIal8VLN4FqfzHi1r87FwRM5lbTyvpy
GAGyE9ngZuwW2xyilviFUBDWgRWWTv9jgtf/XtnukEPDAElM6TEHA512X5C5YmjQ
mrRUPafwx9K1kLht/SINXMxzI+l1R1PGfbzOYIVv3dccGQzI4rkQWkf2/N/I70fm
KUFQ7V1jLo+M7MOQU1bzVlMFh5xn45Zed4080by84NQciGQhlswC2HtbyD1DiXzK
msZCDJMVH77k7ko+O8+ZrOES/akBVEy7l50nfu7T6yj1AxVa7XwgLk+em4XjILRW
dFNXDJ3MnWMyZpSa3yGEYgjEROLXgUQGukJS4Rb4eiFeZzTSIPRfg57yeZZip2W+
Fmrv3zXQz5zk9M3eMnnV3JPPUwL7D6cRL/LSO+he1vONUVWTny3e/gpPGQVYFVr0
vs+f9q6hxdOOsy4XoeTqamF94b5CVkILL8Gq2ejAwQqGWmnX729obPbkE6R7t9G2
DCjVZOn2la8kIszuJgJ0AQFs8jD6v6HVXNsQmP/N3TLvWfpPootTudexdjHpRfHm
SaRMwjCWODWS2O2GS3ihh0tKA02k4Ovfd0lshkakp68wuBVcF9ZeX72NG6UiFmA9
bdtlmE/8gdmyZRm97JGu+Tdr96k74Qf/YxK8w11TuYMMNUCxfBxjE6WGfn+xKUN5
vOdbJCANnMdlMArz47cZFx3igu5NwcIwatfPfQeKfprx7ebtnKxf9aArU94YfXMt
ZAr/MP0EfMKQ7+onY44h3RKdJ6xkOMs/xbJGwYJ9oCLksd7Gr3DALSP5ZMqeXkQf
JyCtQHesHLrr7UonG7o+pR+vgjbNJYhmng6FbdTj6A0YXPl5hjn3B9SH0CCWxLRE
iQ/bbl3KH6b8+aufNFY47dfHL0vZMEq4fx74msDmCfvGo5cL9DzJvsTfBIDFGE3H
cnVXZApFkTSgI+KvBtaxDcxOtZ6X8LRmoVeMOJCN29J/XUeZChYtZsasYbRhw3hk
CRyiQOwP0SPrwWBrC3QSYtOp0kExz93SpxM3O1fVEfFIwA9qdFmOuJ0zP3Bt+iYE
lq3JbpzhYBIYagb7GyW1D+6xnaUxTd/7nW13UdXVZ9b4iOy/hMOY+klc6YwNhsFy
e2L0gip1bCxxXlo7B8Vn3TLRQ9zP8EtHL6bNR8qB/42PjEgvwkppvs97dbULjROb
2RRScXRTSAvS3/dtTPYBylaFTgV3Quz7N4+EWI35cHSHUaaAIog6wAd8pq7khgp7
oIHGYiaiUd4glRarGT/G2DTCh3zsz2veZw8YNcKNjqFk49eqdc33u8eJhDX+hugy
dyr4mamheUca3NCvRncX93BSvkM3LZ8TQki2JccQGt41Y25VnIVrQGOYHW993YbV
+/e9L98zd+0LjXnUi9jTD93+aqLZt22cTVsN5LsHZ4VWAE0dTzIWj5mfAIiivNuk
ZcbzcrjKD610pfMACf9Y3DB7mrTe86shiAS64jjXvYeXmNzkUC6qoCagUacga8Uu
v0WlFcPOsYhtHKz03eC9JODmax0SJHo2zNYxipsIQaloFXl2JR6HfIl8VEjTCwdI
q9upBMTD/z6AE1T/90OC2U33ODQuhlQrpJf8eUGRuPzSGvlTnKLNdY36WXRBprrM
wwOfJgH4IV3KLUewSmlEfP5wZ7gmGh4sXI59B01b/v/26uUUdVZ37+QGmpvWK7qy
IDGv4aPWgP4m3mBfYtn8Td4tjnNrNlCxzO5bzhdK8tbdSLQ92YGmxSKu9D5t0xB8
Ff5LVpywLLwiXrd6Jy1exY+mQvWJ2bC+TmYsMeiQz+unWizZqsB2jULLzeSmQJfL
dvKoQvBRfJUvHyH7075hAq5RprL2SPd/kUu/WzEPTv/4x+wqU2M260o0s8QZ9F4a
7VCcAoOBIbI31Rcq3VyKMwX2hsbgLneT400gq+ITKWKnU5I7vU8QtBgXVTx5IZhn
UsaU+voGwd5sGsCA+0CktUhKgruYFrlbl/7At4B+OjBZTlv0/lFiXdSFASvgNYwv
SNh6T0ixksBlZLyGu5qqMNBD3FkKo2RIqsYsSCp7YV4+PgJMKbY7KsP+NI8OnWZ7
RNhWRXGYK/wtG+ug/+bzcpeYO1dqwf7cjQl+JsUMZ3uvN7mA/KBt/mQuB0+Q4L6n
QhPAEJGYXU/L4PmbB4n1Vrihqun8sNoW+S/T50L+wlE23ObPvreq6fIEhjKiKCja
1hYxD7Z1KEnkj3/pZ8Y3tBUfiuNCXIu5VFDtdDxAuoqzj1WTBmzw/PntR345cLmq
Jn/zzZ3Ogy0nSwyU7s+tqDyrnLtIkZXJpmrzSapADId7iPMvqmHc2OmzUxMtrfEz
7DMEkJQAArUJ17p93G0oV2Qvp8mjQvUbzPGn9Chr8eZsHBM5Kfs2m3vH49IR4B5t
Jdn5obDR1VM3j39gh9IscDH2ywwFBEluxF8V7/FcGBNbEojsqUV3goZCJ2e3p7PV
S7eNkvmwWl60OAhFWOm7vrY3sWjL2aj39cVaJH1v2VIjj3v0ou8YuBD91lG6Nwlb
rd6CgJYGCQTrThuoZc8p6Q7Jl+W60ZDlZnbCvwykA7yttYznURCXH2+wiAU17XiO
6lc/2hDnhl2F0Ep1kosLeHL+PhExE+jNCkqMO884CYc1y9LhPmPw6a3m8yOxmlRH
xZ9Rqc4Ob3XR0CtD/ZNmk4IAuE0w9RESKE5f22srvdQAbqGCmMdledIaQqEdFiZE
TCSWUmh4xNburGPfsI1+dNP8VM1UBN0mCWoW+fGrj9VCP3SQCHycVGKbe0aPXILc
nmGjrVMh56W2wN1GGzsOIKeyUpGyPMcaruE66k/ODnMEIh3bO+TQOsJy9zdqyc4Z
CqgwfX5mcIAm+JkTyiIFLdRTX8kiDro/vwI2MONMQqlKpX05z3U8cbtEyrnt0gTk
H+qJhodjPhKzKWmOIh00c553Tf06Wy4T6GvHeL63RG+CRKd6QwBTAHD2bKh90TBf
4HtxWLWpnUiSPOf7nLajh3485IV8xCKT5KWcQPEj66Rl41q87xu1U3QVRj3iTcSz
f8SgLiThYPzQAPtuaIkx3kGdOfxBKeS7AyAjKks8faBKzqzLUSQ18HJ4DPy/QTxZ
SV8Mkkvm41MzS2XsQsnVO6o/OEF1fouL/GeHu/imlCaz4fenCjKDg35Kjl8M9sso
sEfpcieVHy6nVhQRyKOtbIKecORHp5SI4HR+PC9K1M8itlfuf+SA95yLaJxvk+DU
2ly1AdEO+wLhF3Dpvw+GPpfR9H26BvEBK2MJqBp1p7evvwIrrw8S61MvBm5fRcyg
yS0KKWV+jn1kg5YkRulnXGbE907HuPBGiSx1q8AuBcx3j5wroI72/etTM2ejCM3X
XHaGBCJekXoIi5GogYzvq3FyygejEbRc55F3aE4JeVzlJOqKnk52d6l1p34x3qBG
V5iGYbwYIDsfsQVikM50Vbrhp80fRmkVpcTEVRaIScwV2lhofWcETVFZsnZyKgq2
PhMMSZJl8MTIpLMeEazvxjya8UQvnF2y0Lx7/u0ocVV8Hh4q/YcH6OpWZ8wuWsUE
eu8RVOHvpm42j65m91nmzHx7elef+033+n1y7GOlTD1vw2pqv6l6gEwG4qyWf0bN
NsJldRYcDXJQDqZ3lR8e5Wp6Im28WaIK78n6PxJd8ww157F9yvMRaMbSRKsOKFIp
BJjUZXd2HAKqbgS5Y4c4MtYVdBwGLVcRsVoa2RM7ft3b0CVjYeZJmpk44zUmkrJB
g9nNWluhSX4r+uPJEB3KhFbOvdY9x/G0VMg/zWRhYqqtk/W+A3Crb5wEYbqDSLsj
isNXss80nmbzWrFXkvMP/ywr5LMk+2BTJrNyu3sXpciOSX0u2M0gD0dkyg22JOCw
9SGEAlWrGtAhX1uJdpM0enAkh0zi+Wkg4o56bgJ7Tl8qE39H2H+5pdkASpJAOVRz
h/s3H7bjgFCpqwvNpYi3bPIUqhPSl9yM8zUBgpU7sCqoQKznsUafvQbrRzmoeMqw
b/O6F46fnm94YsolnVIxCiq3Zna8TktYOj/kXt4pXY2QeHAWKVj5LKOIgv/RMJKj
Nauj0Vu75c8b7DL7dGG93xue84LmZtTcDM0CqYD2CpJQVb9EyWnkYxguTp6V/2Bl
BLkzGMlLjV6OcNDmMxLSpe6h+qVYjFBD5CxsY56c0FYmzfL/B6k+SZuNUh1e9ah7
kNOANn55h/VJNDvoHSaTG+UtbkwTuVMcZVzf3szVU/bqi3Jb0DNVEViCO/Pv7Cvq
ov/EQn/xE6W3BVf4vXeDeuBpAz9w6LaUhFZwkcFPgt1v2sqlLh+gdIlqJjaNmdvi
bjZRwU8upAvygaGM80pB6sQgmU01mkSml/GjsduULy1402FDtbcLEg4nQPiME6iy
M9JjyW1D2/QTSYHOr1pVhwXOzXrr79sDLHpQBaV7xA9fAxNhgU6PoCOsWV1ee+ki
q6yz0w6inqsuBM2KswZ/Hrw2LYLKsfkVwCbZoBYYYlexVYnctt0pCeNLu5/a8L6j
l/750CEU5zkMwuWFPFyLl+WX9NbpoKxDSKg9KUfyGrYpBmqyWaogyKNLuCL620hD
HIxIktGc5X3jGQC3fgm0fHwB7i3zh9JWoucy6GyRHW98/Wc+FOXaVkO8W+AEdS0Q
8eZKktFsqQENHOJ08YR/+oUtZhPDYRtkKhPZEQZr3VcVQbaCgiqQx9I4Y80J5yfr
LOFMTS8BPD7vs/wHSythVfFGLr1H4co4DfLd888C80wS2ZvmAFyzX2wIK/sTr8/R
FwAMk9W3KpYSULsrn4MCN3a/zekiXPRTCj9d9T3ZvBV2E1mVKcfg3YXX6owtNxpG
dsvLeWMdWFzjkn1xaQE51XIi/ARkiprZxLveWnE9sVXPVdoJTvFPHFApu/osXtce
PAyVfzhoihj+E1+ENALsBD0y6BdFDfDUGyCSgJh72X7Z7zaJ7vg2VOkV9RLmQ1pw
Fk8kK7PDz/1m+PBi4HXcHPF4j5rFbDrqdzz/iFJkpecRwtJmySPDw36H0rb2JRhc
kq/IvZ2FzP5zMbE3XSd76zbNXpYPr8uiBHvoQB+EshnNFit1/NGY/G44zXf64q4e
TglDcd08vCLZDWYo9swIOC3ytljUQvuUiyIzLdXeaSteE372H52UVe2p8JmRwPWP
gk3uHqbNhNWNZtduDuUG//UGHMIvNUKNll7CDBqB1S2PJX+ZT5Kq+AW7fpC2GBPr
Az6o9Rxaka5hfzv/iv3k0JDKnS/hxBasmzRcl1T9KvbwrheDbx3+EmUkR3td5vus
Vl26KRsy7aY/+7kTA+ZLAdIcgYIOCjxlQBJcqFbSi1tVe+A1yoTZBsEa9axEYkU/
srnCTCsVTfOGCD/M9e8krNK3SBjEUsvfAp3j4Q+SvQK/KkI9I4bSIl/dv+u/pSU/
EoVgBZFEo8taicKFYdHLdsFvi9sfY9XscEOW7jrQPFDhHTjdlJddAQqNmxHiOG9/
MdygtmjnfKSA7p8DbYpXSeQqe7pqEcJDT5zp68AmaNvkV6pCnAFU+ANebU+Tge2+
b4d+5FnuokkC4bG73wvRYJlulZOc/8/spZvSaryxV1XazZY7NDdP9w4tGW0Q1Wm4
HH+P0ovc87bQxyRFV9mlJ/CDZrjJ0EgAaY2Yv4JjZoX1oOrJ6nqli1AGvXkHuCf6
7g3QglE7BpiHMOxC9LFhXTx+LFXReJuav9xORJjAMyDAOMbRXoo38dRmRPw5LZ3A
WUesnn9xOAObMvmNI1ckJMLPLqpTp0D9Hal/Kmd2hrBt3GwjifnD0QWVcKmUgJ9O
hagdJxvPWIT/wP1XeJpXibBv74WYsCtoqqs/nek3j6nMHlNt84sqTmBcT4ZXkVxl
bYNDlfdCjfVph3zx2bzrXcY4RrX/IMreKQSSkIEiC/wsVem0ClUtRQVmypvkAZf2
30Zo/lYXemnL7Ay0VFmRxO9Cx/qjDhVVEiWAyrDaDygILaW+lNWqIzZSiJbcXlLM
ECGuFXLGGoCHYiimWW6godfjoyNbQPtaO0NwIgW/FNQ1+GODTg6R1m5U2319wlzL
Cn0cmWx5P0BxVbaCLYTobjLT4K6vCGN+3Lvt4C9EDEvi12yIIZ988vl9Ucu4B9qw
zhXbJxZTgRm9PT54KnH1CJsox+/IIkH0UBcYDHNHS0vYBNGqrxnXZHEoYsD1JnaD
Arbyz2EP4QO5bo1BA6TLU0xjWQlw2w/y7WcieablO0gn2vvuOZ3dUHF7aN7TEA4O
L7zviON+Ala6MljxdS6XLejFXOY6zGCC3nHjMEsLcpwlsY7p768qN7KQB7ZgufeS
g1z9dkzY90ecYCDxbBOaQs8bFPFYV2fxikkVU+39Z8jgHC5JzmE7WTpsfFbCLDGu
evXVP8cvamsvdNzL+asSbL1kpJpUFooIFumnS2rdCV4OH9OijVKXIR5qz04H1AAh
uLZcMFnq6wh5v0n5j3D83XRufUT3hpfuMgKSUNagO5n9UW7YOpQbDEkZMNFpft1g
7+orkuzAiKsZVAFqIcRhwMvvgjOrRboIdiV/hI14bROTcPDvSewPIcOyrRZSlCkn
JietgLh4qQKGuNdgoM6x6PBvEceoCIKhVwMxQ1ERyd226yESOa5+Np4QcMW2j2DK
MFSyNAtz8F+q1mEiCjcomKsTYtlO/FfJoVZewb3/qPP9sjBmLljcW4iZKH60bPGf
11yqud3hAxdzIGwsQ8Fsw+ZXSmvxQ5l8aqLu1SjbQDUsP6q6wImExBGHXhojBsuM
IDzTb+Gr0lO6cHPhTpt01HM4pBxDzaSnQhy1wqCQIwe8I0EVSVkvfHF8/mmTc4tD
MG0ENJftTy+lP4Tp92lFgRPYLgLzXW9W3tOf2sg0L5ZNbb07QKHyJMmFRU0iUvfI
6MiW1r8lJe/dAwG4CPSXk50YLz/w1vX94KhaeISSza5Eidk0RNEODQhgh7jGV7Kv
E6ocLaqdEREXer73owahUO6mwVrBwJUQXmig6Jauxh25ojvPtijnkbsp+Wt6LAVu
x3srpp8FqVnMJe+1pySYrSlyTryl/LWOWbaFcFCLOLPnzPwA64Cep/UUcFpxQHe1
WlvU9u9Czq54hlp7x331e7WCkW5P9Z1T+PtKoaLlqqRPgh+u7CzJMXAFmWLM5dxG
FZxzbSq773mPWN/LSOvPPT/6L2cancoOSH/7QZsIbqOZfO/7pVcRAGmMfaU1XxFo
33sgsdv7fh+L6bnsae0seH4HAwfYlpTOdQNPW0QGznqkIFOa4pjQppRUX0cAudje
9hi1dP34ryzVf8ykjUNG7auHg6nhigJ/fSxH8xD1Om7ZQwlUuErgTp8T60tDe+wi
92JFDg+WPtPraeM/8S70rS/tcu5ZgpeH8+bqjc8XfRt+PasS6P+YKmOG0yRflW+w
9b+4FbULwDsee+0wtFYt7+irvffrn4QfWHrZ3m6e1d1rz34Y6JNSfWKFiVJgBq1C
NFE5QqC54nEsu9isXvO+ebq5bEsshn38dHwPKrm7RmfUSU32IBSB4YyHcIvExqrS
y8/d1ZyCSGtPhWJQj5gz6Aiy/QBNLx4NuBcZ23fufRldemhoGT6CZCmETFcPaPur
xsjCJaPluCW0FEHOvkgt2PJ4dMBUb0F34w8E0Gi54CRgx8VTsLjwvEx0Oi7Tdqjh
XpMOSMdO5serHNtoPivZHe5DCqaAzOUv3qN8MIltyEm6UqhiXKkfFpufLLUfeVSQ
6mv5pN8FNZHDrJVixcw+fgGs2TDNcRD2FLye88GHtdzpKGC3bzFuYNr5qP8qZLCS
YvA/NO132tXEopqnJ1+yc4B7wgnI6/owIoxcsoPR+hQ/ARZGxAeo4mUb7UwnxTbF
Ao6zLfk1y5jcxtoXMixz8OK69PrJ1xpynstYFRVi1exZ9Ziov/1l93Hr/SdS1HWq
lZpKVseDBjl2oOi7DqxRuQ+5wj/HeXBdHGY9yi0ayglhN+OJtIHVzOyYOJVjErX5
pWKzX16CTYK5z93s9Mb9tMEJXX32e9sNq3HpwgPMcz2Vn9puqt0mBWmmwkglzk3l
HON8lXZ1FTR39tB4wy2fG8SPSbeinPMaKpiKtgb/m8NK3K+L4gzypyLsDel2AM0f
QQYteTacX+KA/BZF4mNeKXRuY3VFPX8NLIoKGfpj60Sg/rkPHspIQPZSS8+QrRnS
j4TUZ2BOWQT13zJAQBYLzoFZV+qMEFThuyDlBz0CloT1OWMlc6QlCv5y0iwN//e6
7mbB1AbhrpkkDfP2ughDXlzabpTxRwyDj0GtR8lGzA1MwEl8oBmCOGJwz/qgfa0P
N6v1Xk5OPMVwXbsXXBBlNYrvatKKH3T8BU+lxr0M6MlH40RuEmM+0UzYQU4T2Oc2
hUotKSS7dCsocyx5R1/v3ouOOIIo3LUW6BH+ZKfDOhhOvl6+jHqCBLT1/p5uaZ6I
/vSpHp5QtzZ035/0+HiMMY7zepnv9NpIM34cJujzV7vtrxABxDc7n1h3r7D82FVL
5KLMbf7wLeGH+r7MzlNO6+bYHAqyCYmMnMbehPbictqiqE/BNckgWSQ5bRNPKU9J
GsqAG5AQPnKkaqYNo5YQFs0FVppSOWfWCCYMdp0mGqp9ikq/Ki3ksK96oP/i+sKn
DQV5FFga8VcJ1VGfFhH1v/tHGzH7wFCcHEwWCpsyuTxLi71LiR3rcFCjAqQpcPZs
dfPE+Hg/yYbzqoIh+jwrQgnjr5iBTxoUf42fhzor6X8Zj8S3VZ0QS60M6BPkJ8iY
GnYjm37L+05bG1X2GR4sm5bkSCwl0U2DoY3ZBNl8+egNrMsstoGVTbRnqdVAUUqI
JyK+GPbItGzRND9QDLg8KkWkar6xlG96Co3qRJuLVuPGWz4MXTPg2mAiBT4Jt2av
IekRt1iaidn8lanY1/8pcJAYDj4icrBG+wXkFgHAiVSAO2cUlxCGa41+TBSZqfRV
9aDljrRf3T+o/5Mfqe6iAnOwFNRM8w8V/JIJkpAA84PV4PwhNNYHJvmW3oNczOKc
VyromjIgUDG1TKdN1aFOCzdjFgRSUnFnNEbI2Wa0uCpJYJadV1BmfQDmUwqmRf+G
/1vOSvUIreY2c2WHhEWhSTqZUvnZEc0rAXf79kMu+ZFJaq1xGg9vuj/WNxpVweQm
LBKLr2DBtmvEUkM1OWUtJVZ1O6VtonN/TLLEFKf3H8A136NW9wj0elVSrLBWBkzZ
YmmV9QBglRJwmE24U6tfpS3CoXWnUtsyisYLsVmRYU2NxFYzUeXu0Wr3Bl5QTcUq
vPe9/SxvmTw1R3zgDQ6JQ4nRJKRcxAO4F2/DDx83A+CSMGky0HTYAVCmb4clJBPl
pBLM05ySEakS3ARwlj9MTtw0uUqh0Bua3XnTMlw7BjZ3HkKLs4DY1/SZxUTPvxrA
pFIqLzZro+UjKYTday1s+ImZxAcQqqYYOEkKvwnlK0E3S4LtRNhgVWwBSQB/oqm1
AoLVgvoveCL/GbgEqmYHXQ==
`pragma protect end_protected
