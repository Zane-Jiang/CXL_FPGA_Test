// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
03uiIcHWYO+18cHhXu5Erdbzyo8q2GCmpUSVQBCkV1PgsDhdwR761EYxBRjK6zkO
05KS03rmy6A2ETM7JrpZcp6++IwwuaHlYo5L3Wn3n1UFGWQWiPfmeLKJ5MPGeIda
/tOTdJkI91AdPn0MDp5cBtznM5kNr6f2f4kUlw8nKobjPmIgjBYJ+Q==
//pragma protect end_key_block
//pragma protect digest_block
GNWY0LYjOr54KHT7oT7rTecQmNQ=
//pragma protect end_digest_block
//pragma protect data_block
UHcQXjmkgR2FEtQvT/QF16HkLVGdg8fi3qyICaPTzz83fBtkfF2wtSiJvvITY/Sx
DDo4v7iksToZfJGjXAHnVXy0QeaqDVtRT6uNGOmhpGXwdqDP7f7/PsgrMukz3wBK
sXLTXpoL0WjQVmTAiNGPeaTa2r9r+h7N+PaCVIqflqXXAZKb14yAoRR5/Aizqufp
C61ynas6Jt7Xp9edAxSA108HSHDjsJDczRfoCzQCvMGAFz5h/zfNoG8jR5zMPDXH
7Pz98319qanPeu7GL8VCP9bBYhegiNmgRAD4u9cJlNIS4NaxRMI1wMRHH+HEBNYy
/wMuYw9ii8CeMMWmqQW43RPZ2lT5o9yHECtwldIUbXu17raI51OJX/eUdV6legvd
jAcAp4J81DNBz7T949yS4yM4Dp/SJfxZTH09jrRn088P8Ax72L6jD56DVOAmtppb
dYClmPnfduOJlW81VwZuu/fvDPbzFBqc+vRmMVLLnq0o4CYYcb6l31Upd/+YWZoD
G/4n5DMHkA9Cfwskeg+MVsoTR0ZsIW2wCoB/74S2Qb+vGg0fapDFyrocmx1LyAxe
aalui37gL4Qf0NG48AAwIkLexdH5RsGqrA4tGdudBz044mWjH2eJDeJ9gzuexqb7
+CQySQ5HKejBfO5y4Zik1U8eGK9npxHLiM1UBsAmbXrrRGTP8oM3CH6Bd+GIvaA2
cl3XXuXwTXCRDQZelrgvqcERF8V126xYPYQNtT4l5dxtcw5jPMdOICOuBrTgn+fD
poeL7sl8g+AA4dBWFyPgj4vllmvCAXYL6link/wNN/W9YQjdM2n5fnN1nSnsWrlD
Xb1y2UFcKGqrQEsCUxxnJJYoBANUkE6v59JEHeTWxkycBw8ZIWqFDcj8lgpsdF1v
T8Z7+rLm3nPce3B0zDrA6jxp+qUVSH8XuXEmx0ElvldV2Gl/OS87uujlnMSwMnZy
2ds2sOF5IC/seMjnSgPSfEIGVcrr3zOoodEVE3g225sI3UxBtmDmDNcJ2P63B2lX
lxmN4FkOb6yyemOcDEfh7b9mxDc9Yqwp9HIvpPHUPLwPZ/HMj/fSxhp5vH/zpYij
nGRh7kFG/JkJykClReTh9tKpQeG/beszr0wDS3NNId9hL3BF9ZiG5kBIS7zuUEZN
hOfcESWSmsqdxibUY/B1Gi1PsjHluk/43B/qFAKD2iiqg1eYsmgmtP6nhd/yPNTw
/sWJ7V94ms0juCZRp2Tr5x6Nkv/hUNu0wX280Si88KjWNHtOhf7UtWuBthFGLLLH
GalJ9KVdmCmT25Pt9uvNJuXFVzO3ld58NddHlq24bNhK1BA1dUgBjSfCz1p40z54
NfOpvSHbl+tVKinHDjIK1yQesZ+hpTChEX6yMnm4vi+tBWNnZ8PX4gWqKlBVFSau
4H9yyIo9CVH9nnab8z3pfHIY8f76LEEzRMh8cmoXxxKmYlAELtoDPy/7GWd8geEp
SOruw2mDEKlJoywd2m4XFPL5se8alFLaQN4t75vd++Lk5gSjFkHQE9oq2aGHNyQW
7sy/r79cEb4pnpwdPc89iZ2zscpig0+e3ARiamG12atllm75b6HCKWr8GzT46sqY
rMF7/uSk0yWbmN1VBNm+kQR4ONcTHFFcXVKRPjNh0OpCyiJu2iHlzMjcm2TM6/LS
6wDc1EN9pyBz2ONVtHq4rVlzKzXKX89tUrPPIBiQhHx/V/S/if/mo+l904nWu6J4
vh9f5h9ddJW8wb7IhG3sMHQR+xU7JJfLyYMrsoasPrQ/qWoMZQnc0lWROA+2fGpA
itnuJq5UizN77fEVksnWqZocooJW5WHR/seEg28FD3K8GrwvSj5r1k7/HzJmCM/q
76acPy2HxB5OX9xProaLASOyL8tp6xk1CjmzlfuglPTC0elgf8t0tdXddb4LWwyH
ZPKKGPSOtH8HyAIF04M5TmVoLePNDGaeTjrLzsOnW2vQRThjftd8qEBr7aznDovl
atdNY36NwoChV2VWbEEqr8M/4w4uAUI9nyCrr7MD1JMmJ8xnRryoxCl0Z2Kekl4f
frTBb9ZqqQNf3/Ln+Wbmy0V7TDDq0VXPVG9MRpm08xZ09FZpFSeo/h5x/SLEb823
8wqIE54tvrt9YTzaUn0NL9xonM6McY4C+/zxufPSGHW+Ww1uos/qFxbh5RYWUzUn
ceFFLFWkvkvRGhl+qMBG3vpFSq043h0fhwGEaENNLLcHgWh2ZFbcDUoRM+sZCnOj
4zTY7iKHWNHFEjd6CzwxC3cRKZ9cte4TAG9o2E95RLHJ70OQyuTBDqJgXtpOWc6J
mTTwYFzqp5UU2rIWIKftjVyS5y08h/t/tvVEZ4A5RHZVOc7IItlgAgqptW7l9WMM
Z5XdqjaO8KVV5Nt3vWoRU+2mcP2/4tnkswvdi73rWBZjKkoadICbxvFLLvJ70yAI
6cgsXO8QArEwFa2FoFuIDNxqATxReA2SzJN0T6r9QLCADLkEr6/jI6m/Xo7GUr4x
b5btRVqOi82w7S7lwdZUjWBQrFVFkdRn2xiflA59pOen2xBQ7J1Ys+HiGPzNqE3B
rojR7jK89fWqHyATrd75yF9aPrQ2AIuw5XE/+sUORH40E2HhafrTn0xG/Lz38/WO
qicgN9xVyVvmX1U1iFvnSjn6gg+jQh/gAtyTQPfGH11g1iarmHtPaPkRQJgUACOa
dcNRUVOfFLNKBD6cEB4ezAcwfnkm/7abDDKesKnBLaXSWMMlBj0ooNBKtIeXqA12
39QZLXhN/RdFpyA0jecGevL9AeZSNgGE18llRwyiJrqzL5JyHKkytvT3KPeIRrC/
4EsM18nsmG8qGHP9i6dvrCq3rCrk9k/KVin9ADdfp4/OchX1peNTHXSNi6RpTRW+
n93iNC4OxZoqmrf97mvBa6Pu6kLgnLouYJj4hExveKO5z4BitgbdNNQsOmQV1aQ6
wQUfPqYd0X4zD1+B2EyKXbhXdaw5ZjmRqFLk311VadcrW/ddyoeZyRD86Mg42D+i
0x8GdFk1rj9F6/pKAxZWUDuO6dvRfmfe8tOAZEOPasgyIDIGzsu1bZiwj+LOn5fY
j54vNlnbXhZNuQusF7PnoZsogQm/Mb+Oraq44LsgwUv88opbNSGPgt7IsxamlHkw
9gWUyBHyCs3Im4vgHx8pde6gAvM+TLk8gvKOKTjsPX1OXwa9l/cwxvUgxcMuaXjS
rWj6/sm1ZSxcEmRr5RjO2i714gkF8ae8wPgjx3zYXcvEmXHPA4cNBssIVCxuLqfT
vtM/MsUVc0PM7YAtoV/J5Yw5yEBARHcWlAZ7dXEasf+dHz7uZIGjLxFJ5DaKXJBo
mZ+ClLHh3J8NcOwfpzLNyJ6iEb/DDdvBMOB+nmiIoTdyx8xOAohVZbbp7+CQr2tJ
0MmhGZSy7gcwoQjVM/m20H+zjmWr6iIID2AHkVEjQVewLt8uRumFxlKfRldA5wsV
4OF/1DtcKXqCfHDGN6ShWoMN8+DSQey74yr2bvd612unwY+pcrbznqoc5+P+az5D
y4KOTSKaoshTgHScBw040vRnDC4Bl+h2AU9OHvJmh4eBc4b+K5RbdsYh3iq+mxIt
2F3grjj3AplhRsR/JAUV5MlIWXWk4D13X6v+8Vc1AhrjFSV8v8+KKEdRxzj1tvZc
XSSF/jyXv2oHWsIEx/iPKWDHZAbAj5ZtyF0cykfrEHYeqd35v+vaVw4YIcPmlrGq
nt/pVtIA+irA3j+8rrtiJ770ijArM5/oXNl2z0JVaDvgrVKZQyamx/XbPIW8dnpo
GT218wppsCr/CHF1jjKFhac0S0gsgEIlICPBosLTHXB55MvLqXSFm4Y4wIPi3GG3
Wc2jickBaOwSNhjXPVqWK9txjctV9G5OOa9kB8IYXFOKi0y57MLxrnzZp3QUN2eV
xpKwqhd2Dv8ojiEg1wYWCwvht0UNKyLx1ep0UZ9OSYmxCGvdukkn6sN1evIipnEr
WC4yZEHLWI5J7kC3IULujQ/V2s5MIIEv/+vo94LomBEnxxK4R0T9dTqr5iB/35gM
xeRH9WzCmJCHlQwak62WUNlfO4QK4JCPqHVy4vySophxGTRRmjw9egGQpqED2IHc
GyfVM6aq4UVQorw6e225KlZbldpgwnE+Krm838OK+UVvWekr/EtWU9HBmbE+Y5Rt
5kJe63Psx0BXc6ya0kTPX8JrcSC5HoU/eXosNwAzXpd5KRvFizTurENqPMMIq+OA
Vy2ahyvf81W/BdnpZGBqHWYP98bueXPPnqLF/pclrzZ97bKuI75YlVEP6n+LN2Xw
nOoJRRSs0iR8V3UBBGJW1zy4eBO7LKtFFvZ3LAWB3D5jie/EBoaFClaRmIPg8Fjs
grbU6yOh2LOHRZ3lbhkHWFH0JBTy1ZMKy0iCKecdNzNQHMWkvOfA6q9JCOD3KUUd
rWfMPZIrYvZguxeBio/Wc+az3VGsgv/FJhAKKoW+fcOevuNiNu4TeKcZFaJHiMSk
wXfrtdLGGz1PFzMnYIw5QwfNufYLXpVHEhPWHjG3mS3YE+WftGPmejxxYNzPQKYO
Y38VVw+nOOr06LvqWemu/85gYj7UKBIPpttHiDdrsT265LYj8IlZqNcU6tXtDeZX
TdmctQzFGlqtj8MgPluePxNBy8vQmRMFDUCQQ3KJK9vr+jpsT+k/o8DEvOzIKSwD
4+7V+JWJIgVrF709cBwcjXi4CDyRKnuIzl+2b+W/uT9tDNMz5LJpV/eCyLrYJJJX
fvqFOvwY4m2vnE9h5ujSafiaF5PZscNFVYsxOhQPY7KeW7XNkH+7awvMyZhuMToD
TOeKraMLs8I/8soKpzl5PeUpQif6/oCxrV+SYfUHbXOLShmboPptXSXHfuzahlV5
mHcQDtNJxW2W0fWlQSeZFfHEGOYDWTnHOzgj24r+0uo7LwXZ4UAIxQd7E3VKJfev
8b6vtVgseXHou8OfKEpRBvALwSAwD3QiIcgfva2w7SJav4l3dZfEs+Qb6ooQdQb2
KfvruS2GH3uqQPE6v+6ohquvdEoK2lWtA0Ji5B8MBzF5QWcHt+bTmXJ5V2WcPgeF
e28UHYlV4rgtrHF2apSx9uvGypqQyjSXR1mMwAHDHPPJHC5SH65r5gNgwq+dSoYU
RJNoPK6e0CXWD1b8YCDQD0LKilfnTFByjMtkTApWm2Xck9Zr8u+E/Zdm+LiUXXFJ
LbvUQakfEQ5j16jf94ziH57pmehARuWum7q0McBAN3EwRvlFBczAT+R6scVAidLm
BGhPss+OlUo5yY6Sqwc2gj6Zv9PvndpeZrl8bBVEatG2tMNp1J/eqbXQrK0cvDiC
2wZTuaPmZG8O6DfoYQgEcrlN2nrKuK4ig2crytZ6ez04NmU8J85tMA/eImr0b3r6
UBxYgY1Ay6ZS7DtuPiTJ0B7leGC2h/SFKPuPdnSSO6p0IIYlFNwEWjQt0g81dgI5
fs3BfqpzAGLT/I9YEA/04HBnn/UIsdGtaNNETvH7Eh4oQABqnnKyk2NfULgYf3ev
31p0ZP5rknvIkoanAS8SiKVy8uVOQ9T+q+WH/IWCqd6r3WvjvV2jtc3wr6YmXbvC
4p8aFPUxW3ojCjuZcd1JF0GvVXhrBGtPImEOnnjINg0sZjcRrBHU2bTAp+QDNZ/n
7Gc+HiLluBlBpEnHTJ/4tqRoG00k6GUbU3Y48ap/qtHWGMD68NY7lR/ZVc5qW6hy
roCYV8vkindP7Pg9iEdV8CDobWOFhfIHUE+eENksPGliuAOK6KgEh1+fdNF53OeA
Pcv6FZz4uKuEkenmBSim0S3mGrvGXxlv4fjbP6QQvkCrnbST9XocxYupH1cLhYb8
nsvonVTLIHY8wAz0Kh/xHBQQzFA1vlMm8rQBmY6WSSqE4QfzzuFOfsi9PIjjGCvS
d+7tw/F6gkHqk1wNzlvJ/Xc99Iyh1iZdRauJYElqDhgp8/xJnoReOqk8ipwJ8Qqv
aUCXNyEWvZm8OORiVNDvAUZHFpxYki6Roe+QpM9yIzPecrPI+v/uqEsn5NFzcjW+
vYp3H65G/VR/IaG9WJfYOVf3yoGhl9/OqyM0QYT00CJ+azHcSTa26bTtO+dXzddn
GeOo5QjSvyfSLjZDPFedmMV6qTR/m8jU49HbjYBe6FIObAHvFi3Z00Maeiciz7Fg
tSTAuTqQkPCLLFG+u7T4coXQmr5bel3FDPrINGal5A3Hs66wuNlQFvw2lBCxIISa
jIy6TwzhZJCa6FtvPwTdq+SVkUbWgEC4nngnyVnLfjp8haiSeEw+0It4Blu8AkaC
Guz8F4daxxiTnKngVEJyZOb2tATb7cfdQppKNCQxh6fbQUw/MjbpOFqPis/YNWBS
le/rTjFPusVgyDS/2uV88inmNcE0h5ubqmBQvZdW3NPjD0mQ/ca3ZacGufCTdRq1
CDbH+rOp1J4CjXWgv4EZCR7oJzvZQMuFC+qR/DfUQRKVWSLJlBl5L0wnZiaCB03W
j0UXu0QdMaRuVNIBbR1phHYd16t+aMevzxI8K+TkbFMbtXoE6+JBE6Ql6FxFLBks
vFsmJd1YdKQFa76JEHw/xjA2+ybaeeFPayfLAwhxoi7se4E+99Ef8uxghC16lI/L
mRneUkECCs3SqRa0oDnPXyGv2//oBNYFzgLKXmWg0am5i9PImvJoYlWw7qnAnnO8
fxrVlqdWG6dS8ZN1kfj+HWapOP22mP5pQANRclsPeEVWHOZ8fpA2QK2oxaQyRn6d
PVJHJ3mIjEWXI1lynncNFlQ+RGzxftwqP56AHIQdHdsBhswb3NmWdE3Od73KqdYf
ai0QHM13QX3sn4TXrFnNJv0rPJ2x2R21L/zd1xxMCzB6MyzzEgOlNlCirynZ010L
YoA+XrPn/pmB3vxDUxaWRfa4wGgwqYtag5JflAEP7vPlW3Sh9u8h3vGDMoqVRvzX
7keonbtCpaNaUiBxArMfwuhG+ANvuJYao5KOYr98EbGVk27MN18cVyB/WD2TYAgd
d02pIQd0WQHY1ZsgDY/y6r5ICsP0yusEzLy2pPgYDX4lT0qELKmlDJbywKyY+/gY
i9/vaXTMnUVHi9zqZDoOqfrZZsv6FgOgClLMo7XVGUGbvWDfiWBK11ausCEnDTW2
uCCZv6hPn/ZvS3fWe5gbBW20jDsP5oFewB7LrFhGruTjGg31JiybMecJbk1Sd/h9
JNDlKkbuCB7lzB1SP+Q9ef+kRr5Eb0+sVq/RrWfWkReY5aR9LdS9j9D4PkRrjyNF
NHsW49YP6+9YUS1fxR9VkuIKDIfI4FI/I1Bv9ILaZblrsrE+a6ruus/tWBGg+AV4
Hvw5rH7/kuK5KkTbw+MCVFMxhJLUROhqhzbWlr4ml5RYCOamZhVewaPRILxsJ10n
VDLG73QtZ2d3CvSrR+gzM1InWbeWRDebmMzM29PuSph0G79pNGRt04abYgcwPk84
qcsPqJwOzHS3H6VdcYoT6HurSw91EtVwjoZ2MugVLQSJySzdAyTgA685UCi+JYrz
lcBOtxKlviy4IZiIsHcCw3iCNHZHEJIvftk+Q+SI+YdO65qXOAXDXayNj7pw5uKP
uyprZu83fI/2HEXcSpRNnKEN5kA/woZmDLPCp2Llvtz/bQQxSO4CMFrytIIjYmib
K99R3aL+7Fd8fo1/h3AIRhzsxBu7Tt3nlSk+09Q+qOJi/Wb2bfvQxMFTUWy0SXBU
3xHmxmQq5T4Z6CY8t7dc+RhCqS9pAOCohwv5h6MML9dB6g++OC8P1BTPYn7j+gbQ
XyKlUvdAp1u5VrBaVfxCEInRDV+xj0nlWVBQCUHIVo6SUXpAi8RiZX7IIKAU+pfQ
99ObCWFlp4VMC8MDiJsjlnJNbmXiXaMQg+0DS0KxLz2U/b3TvDm5KX73/ZwNFkMo
lGjJUlHhVBcmeefHRRf3KqCg+3s4eQKlNSnsAS+xYGc11mOcEFrwOZ09nlgfzsRs
Dg7APO41pkGhlSSj2q6MBSI883pJbVzeoqbvL4ydBbm0f99+TDXWCOYn3iLH7kOB
icBxpYumw3+zMnK7jljD8Ryp7ag0+3782za5HtpUTPc4hbBmpY7MmAQHQfiYlqzv
7oGieDXSokglqwobBo363wnIneQa6Ur8cKNX72M+dTVfZpi50+/u7ZatiZeFBjZG
862HXFFHm+YAfotfnIQ7ntCP1Dc/r4SRCPOJWK6gpmN2A9z6o1nMBITlX9sF9tz5
Jind8b/sqqv+PwlIrd08yR8yQTpdwL54zSI8j35O6xxC+8Cwt+DM0w/60HJ7Md8V
nKtdVehQ93kmFFj1iVzbDRhQQNbUVY/Jzcbl1bOmNIEWC0TtGUPAa0U9zADRnvmn
7nVcJmnSUqpAEIPakwOh1AgJlX9P5Unc2SfMa55sC8z3TL73O47PxrQi6OsVfip2
HMzpro3DIFgabmQVljXwD1uHadmSP3invsW+NnRgZIrO4p5mYAvOSMcAs4xOjDsr
CNhNpsHdeeJ0Phnnk5HnPgVaKooyh0ZDkP3aedkjo0NNnxFseOacyid6qfZk85KC
nufkuU8HiDkgukhGfotgsY3bwdnOEDWX1zg/GmCnnjmoH0UWDS5nM+xVI5Il8BgP
h5sbOjBLn06bct3p24RBp877Sdi0rR51CSptVLkNwfk+KnfdqdRJwbIEMQTLvJYh
gyMaoUmm1mWRiMQ2FIiXpbI23TgQz/QBLjPiHRME4L0AM4bP225aWP4CH7QAMLx2
6ASxOLCwYlO2XZDzmkKf1HBR/isJGCt4bvcFTzdJBOB4PC2DgHJm463vp5HOCHEX
u3joWXkS6eCICScR+1Vj9eOBymrmHSfLMwTfBMiPJ4DVgb/xMXFyXXmtYHR/TcNP
m+Bq0LpqK0IIjtLg/rk51s027MFXbia/U8VtP1gP/aG13sXaNPzj9fxdWc8pf2eJ
vwjh+IwLuRpWHHNKrnYkKKidVvOIAoH522+/3LzpnA3uADpCdb9atkoPbqVam8FA
DJcEYFSe5YpHRhX+eZnjem+JxWE1JL1G94lIhREPeNBrRl9BUoEmHf2b0S5n8jD/
5rrmO7uaA/VugnbiHMDwNoRY6cEyycTBKWrMaVwV7aLr3FoVs4wtyjUwSwo6OiUX
Pd7A4NEqcBP9JR95qPG0ZCMLQXg+GrJlco/LSNP3eajeOckM+N0avXYFjWKT4YR+
d+lJs5O4ho9mG+ZaBmUAFqnI8o0oyjZHIDNzhkLLJsFBra1ixWNala/ZqDfvO78i

//pragma protect end_data_block
//pragma protect digest_block
0NawkPvt/oSom+OAnXLGQOV+4VY=
//pragma protect end_digest_block
//pragma protect end_protected
