// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mM1NTWuWoY3tGjo9QnkhxkN4MB7r1ASAOpXhmImfCuvwa32+vmK8xN9WDP+ahQNiuIrIruR+2pSm
YDzYS8AGX4NuVpnXK0eSB1es2swKNNdbEpujVMmLoKfm1EwqxHMGAM0uJcReOrrwuGq8O6kZf2xL
u2+2CTgfxWyldUYV/yf/dwrxPfOMlQn9Fq3bzkrVeHHmNNE5PZNTHHM69mjIboftI4c0m+6vCvqi
ukwJLQYacgGzakbcMNo3UqkrpdMa+zFDUY+g6YJWIr+5MPt8BN/B+DGgh5n/KxoITvjIZeLNkQrf
8/wUaUK/2y+o9qkYvWVZIKn5JcSQZbhO/6HM3w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 20000)
uu762PKowuMhbofOh0uS5/IkGFx/To0vJL2+XZA6cCy0P2aARURJlp/U6bv7vnIzlYWrWL2sjyW0
OXRsuA+Lx3r9ee18MbpqKn7o5WggP6WoYz9K+cfzPRjcftFu1Rts5xX0O4Aq4Xaav5Qb2YwT/S7n
ooXoLcZR0DGQbwBgP1ayw8jsjVArr68VECNrHD0HUkhf77fyBgBBCv62MKudlHe5qejEshQ4rD6N
6lVls5kWOi5DVY1N95J7w/qupgFKnIlRi2WDeaJc5J91GSKhJyV2sIfuOn3GQW3Lp1BV5hFCO7VB
5XsXYiqzhY0oQ4/rl5eIVSI7+1jTXdZliC39TrXvrWK5SSTXwRNnkVZbYWsj/XzDAfORh1fgH4nq
TrMpxGIt5kXBsKnlLuEXucdKHsURMGRovPt2Jp1nNnmO+k8kHTG0ajoD/VByPgt6nkUCFqDQPmtK
IMBDTp4ZRk4B1PXwaAhogSLV2YsJzI06IPfMfEl/VcjIXnjyVo5rdMLV0HqCblxTkoStYmQxVObM
2+vy27yjimJtNfhE5SOGn9QwIrgzb8g0x35/C47g8k0Ic5uxNHgOU0hqaIkIHizQSb+6bK/oSs10
9VhS0ryyvVp4Muhkt9vt8A/mkNB9rPJovpfvLotXStx1G0FVYXO/FTnyV1fLyn8zwGlrZG2qwJJs
/odA8kRsdaPHvhI8Rl1nzTRxYQyH49nTQbKWUmEkHgqItJOjsN3kfw0iO8TKTJJoo/fTcbqcjYkT
MjSFDJXZAtReTH1uaLs7KWghcMU//JihQrZN50A9MgCf3/uBSoAeey1jGsQCETnw3tkT3CqNMixP
TD6YgVqqpg9U1uNo0ZfieOFQbGlb6k2V0jTJA+TU5m1AfUo/DWT3GIRHPhkH/jBUOpAAr6Yetkck
iM1n++baBm6Xl/RT5DmyaHcc2SxlC8XddEkj/vdxUS5SP6flJeLS6diNShnL6xkqLwNbZNgXlARD
/IiEaiI9K34JJSsvZWI25U/Lmib5drMZJdlVUbO5hNrgRJfPMj0JdVJsOMHHCXgjG8c2mTBz9DWo
OXd6YaI3jbCFnLHbAcT75YPeYsVBqTJhBf2N/ikvBpBDPzf1Reb8EyeZoUIwirsHKWRZHGmB5t0E
5ebui+dm/MXfXbh/dIs29yKNgDgU7IKHeWxoPS9BuMvyILBN9Lq1c6r+UN6p07yTQ2yBlgVhxtUU
VD7Z+ldLD1ugmWcpD++mOd3GhzOygPbB+lZIs9rxNvY4E20iYidpqY8xUVxlTT1b42mr++lVHYz4
xC+b3slAq0CFzpawbID01jfI9AM3myvrlP2+O+rCi8KLJ+HV1aCyrCLaiWMB0/8MHc0VoJmUApkw
nCK3Zo+B0wTrqrPwhi/CThvwadz2EViTtX/9BW5+GSIGdqopBb9J4zFpXVSmNAfSGq4oQqDO/LSE
L+RGOz9L6YcwpzZC1yRESGW/pZznyGT6YlgL+AU+kJPK8ieOlJeMedD/6vFbFswxY6DwIxAyikKs
xo1m0XnCFmj1MpyxHBsyQXTOL+M8C1L+xiwtB7biFpkHUChXf5tpM1Wo7fbOcWU1pU62ZtzGWR/5
jKbPpqdBlsAN85pzrMW2R1yYX9IzNzIMf9KXosLaiGqg/6wFN1yPi9992Zim9I0AAUbDt/M3nUhg
MATjicniPySzcksGAVWa4fC5nTVW2tjd59NZyh4eCPUX5NeKa2xBKStjYZ+X01b6mT30jf4MWtyF
C5nfl+CkoPw2EQfKDoa3yG7T1fwZUaHE2Hils563taRnVvKpXmea3jqB0t9L5c4FLJ4Dz77jpc6j
yIYCHSF9GTA5Y6yb8FHk17NDQin3DeMhIxLCQ0xmHnxpog3n8RcVVKrdBo4CGe1A+RYuf2/0AvGJ
+fx2u2E9IPQxMOCaIauK+eKBYimKwRZZF3VSEH21mPlqO6jZV+pxuDm27ffFdqnU/y/1A83jUsYr
7KGNZGksMlzdff+H8/QpeAGtYj8Hu2Lkjb7P18tQ5UWDJ/cjni1+UXTvyjY+j0B8FUHL4XNnN6ME
rPQlXFQaQhTHQBAYsC3ILp/nrEbP6lReXWUlqgOhRG6/UrTZTfYNWz7AJeWtEXyjmHPoObKulyYl
ghUGD8b7UJPGnUU8TDf+rXAAf/zUqxm4RawN099B5VWubhtS/6WTm3sNZwi7UFcAYZh/ZObcqQNj
+TxN73l71BSMBCcq07uQIXT18IqlcHDFWNuwB/GsxThM7iKJmPOTDZy5ikohPR8ONy+8cifqDVfG
9MwROMRmK7D/jYGcEyKP91vKfJzEZljXiriC4Q7d29+fWQb1gGjxg57+v9DKxyuJ0PDGjGtPX5MY
WECjKAa/LVQXJd5BgvFLfDZrsn7qvUuOkIng8LSZcBruQ/+je4FSEHRyspTa8eZi7owy2doJg2+t
Lri2cxUKsfdy7bl22YtH1EDbT9geRn2urGDSEG3HqzsHMUp6IqQ4SU7M6JsaKSt0F/hKG630nkVP
cnF4Yh6iZzPR2DsVt1r5VylPZTtur5YUMT0JqyNPDFucaGogmnK4gfRHUliOGj1FhzRORgUvqik3
+vK/S6FlrFcrf6rYXVVQ8ZJz+XzvcnnCG0NKa7oN44oei2CkuxpgO/RsCbEJK8vLiZ9LMqiWRr9g
SvyDwZxD7MD6OZWDrD4N6GR5KtCELGQX4E7m0kvPkvGsoT3DvWXhqq6uI6Ll/ksqQ8lrr22xVeIz
PEskIK0qW/E18OQYyVZ+6Lc2qdTSiiWX7I9cZki5SQDSM7bs8HyE/Oc5LwCYzY0HRiOuVAIhk96D
kGsMd47kUYG03TH0kf+wwDBeUqINosZdIeH1ULqbmLokZDsqgkx3lhaRanG7JK7HBLzsr4kHP3YJ
hI8/GZ7P0WgE9ykuavxCaNdrdL+P0Vz9fL8UMRpi1NEotAdyDbfvXU6Yqd3c+mzJlBxVnLdqaTiv
LrTeE9pCmk3vBLGDq75/mG5puHKJP6WY+BZ4E1aYGUYBkq7dksK8uRvJ++DoIaWN32z8NZUtZfhS
GkiLDO5CVeRFxEwBKDwy9rZK569N/FEb33zaty8i4wHemm+kqPGaiqlupk6S0xvG+PhZuj6YCcoN
BHvwKDzDfch1mRphvDXWH/cSKP0nAmMTcNOhmNPqoMSp+MVnvEbk4EJUo8ld3Y8rycxUlIc2Sa23
fxR3QIlA+Z0u1b6hnRnmTjPEYCNSWW5i2NIDWMFyqMq2x3B+oLy7WI86VFRfPW5KbCqnImdnPrNq
ZlGLuTu9hIu6fEkusqOOCefpKKCiIqYkdxHqSbH6wjJ/N12tSO5KQW8HS5ZrtjEkCNHNLFCZLfof
Y6cf/XPcz8zyNHLT3ZZOmlQd2nWh60h2gmC8UajglnBuSZpvkfKm/Ok3yA0yKCsTD33p6d5I3CtP
Ca+VjNjxgrIO3JaEBJILKgBKs30KHjCISkFQ7wfdE2VxzsyMs/X9R3o3i51XfnAOnblfTMP6Of6n
vQAoZ2mnLXMGi9DUL+01YPq0FklPQ+H4qghByd3F8Il79+T55zH+dbveKw5U+WgsDV9WbXvrJUKY
FratgcF/EmRfbkD4aMgrTYAZIhOvVdL2tNHm+ARcZBoa1vl45i6W20K07G+3r7NqMhLVkw9uNOvT
9uWqzDh7JwlyDBAmFLyzVTmpcZg1ejoruaEI79/cUlP34q3bAvJm5ZaZSzSgr00Nq8CzUN6fNnPe
xmlPlh33GptO0udBvAkbkjWFPisXY4TYzpQ0lloYjxwH41kQlH19BGxGPF6nL3bxbND3WTgAR7Xx
9LdzdCY/CRTcnLINpcKW8NNwu47Z33LAI3osOLUpn9BDEs8spFd4UTW71bpOuNvF8xofS8GhNXr7
fdyNqYixYOgFDexOxxn63iTTzqRWhATq+mKSJq1Y7WSFi3ShmnHCyNF3zEov89ipQbEF5JjjRLSo
snKYfxNpblqFwXbKyWvH03FB5wXQwx9vj/m1/BpDRWaZVx34oS4sff3e4nDmrBpA2fKKdOmyJCSM
6gI2nlDZJXK9+BHicB5DpliGD0Y9LGPVI7eH8ITVouz9TuoW5T8E2+C2cTe36RdwvQOTXJ2Ucsxs
kpzX5Xwf+Leb8OImNxc10mO7udd9eZrdJyqnAZZofG3nOeGyUg33Uw/oqqYPmtDX7d+UhtKO1Bvw
1+GyblggOacW9+Up2kIQlOXw0cqjas/4dOVizMbTUYtxssx4oKGA64xn8zw95M/Q926sojTjlcr3
3rfjIwucp7nfXzm3MRwyLl7THrslLiWN1jTFWj8dHtXLZJP9MOiGp5fTzdTn4zHf4WvXqfDHcNjP
PfuCR0g0zexN7ERaBEl8nyOBx5nJLXtssTgosten5zVbUnUz7eywRENp1ZqMfz+/Pe9msZECu4d9
wNB+shcvet1P8DbLs2bSGX38Ri/e9XgMtMB7atMtxw4G5T/SwOQ7dq0nOkZntCaGhtwEOsu8MYQw
B/b2hLnSVOS73tOwyaNNeHr2tlneOc7cj5GP8V1/JD6s4XiFHYoEhYRvYwztqICXRn9igGlm54Ft
RhRwZJyN3Ye8aedfXQAclvFkyAtUnN9czg5O2FyFK+upDbV6D5RUAQqEicKmrTIJVwPtm9rV9jiD
snx8ibHRnlEiLVx7Ozti4ytLNHESkTYAq6sQASnFZicFI2QKgCIiBMxm64WHgQ53aiERs6AFo2cY
MFjG+A8c+nVIrZcdDvMyUjtYac/jz85f8KWXQH8/fusYxq8Qgq1XalzeGDH1Ur0dkmpn8M38mNwp
SFUXDb2BkEmOuxHsgXwuEaaiaukYgOQzCtWv0Z0MkT5vG+cqu5+U5/EkYYItgfdQX2Mu85zotv14
3qDpZ+LrisCb2hCfUeReZpkMxTiDJQS64IeN2Ip3YdzEKmymr2KR/k5BpZ0jb0NrK5AAxaMmLJti
F38y8XWJsztdQ+ZnXtBiENzufzZxh9q7YC3dd+G0F01kVASIOXWgylfhFAfDt+I3TuSoUKKj5TQm
/2RtxeA4RQysdCQZ+eQx5rHre2c09csLXSlFce6UsDi2Toj1GYE8X09jUL+0KUAC5OMpyXbn3wsW
j43lKFvCfXlWiz58G+9S67p9D+OBOhQCv9v83nmfca7O4sXBPjrbtUKWUaXBtmF2O9r2okb6yR5r
7nHGFipDYh7TT2mZB8ZzFi1dfUYgideBxnEilJxQ2/A7DT9jflu/IQdDOJ6XQnglt2LL4jkd7S0c
tC5pZHRxmuvOmJOCbhy/ttEXGlhWkLIcQgIkUfWBfHVcZVkLG6/cY/EGTPIkTYj0goZo+CrN9fDx
5xDLv2Rr+NHpt66ZUmtZC6ubKmmCtJDCMYR1fWAQHFPKWDlcxNYyy0QaqlLpADL+NIJ7yDYjH5Gf
jCsOYHlyg/IjWUcTNT1diPsBzKigNW9m4nGwVJhYcLT+9wO9kQiEIiOqTD93tob1xqrlKaXhaVR5
+sOGc5lJmFK5A6liEVkDfmixXIu8O/IEOjg3lA1E3L0JcS0wI6k1aedMkWyBjyUmf8sxFWeaamtA
9/ZHXCZtLubfUj3cTREZQEaRKJMLMqkBYd6zfBCQpZuFLOyklmIqya45A3vCmCDEQ3ZsiqrqwecU
OATzvoMutww+/zLi9hBdJ//kF1RVx919zD/8eaumas3Eji4xQsjD9iZ5j6izr9yHc0Wmq9hdcu04
NaU0nQzmyeajJ7TJMlTiFq0zZrN7j1DfPnZci2F5jBs6r6YANmU9CP8lPHOZAa5mJeBviRBd28TL
tQOyj/2YG3yfo+oUM22vBCXLEwfkw96t8D8zK67Dg7loduvbi1BBu2RglGSChX4F3TYWrbrG7M5v
3czUinCb81A7fP0aSi1M9wmZLKAeYQH9jnWZBek9MwyOqHZDZR20p3V7JutovHznv0PiwuTKPnbw
5Lx4WFoK56QwARiU68CtLe1IMq/MYBpS82At1/ydkkFgcDlY0QSzU1nk2O4mU5kBc1zkERvNCVo+
aW4qM1CQXocvEoYsrZf1yTOHXKKSnP8afrnsMDYhUMSSLZUtezz7XyD4hyVDg8TPHuh1B1LJpirU
3ltsyXrNbB4UUZVC2rGQ0+TmFBEhOE/dEt9o5fsme+YY1ugmJGvWLUXW/d5jt3uSU0U+G2X+kxIZ
RQcqEJeB9tYGglHXh8n0eWx+UTDI0pyO83M7r654wkg1yJ+uOWik9SP1fIa5V1lpfQHSZHVqUcMP
Z8V2eyGT++xcfUKZgTh8HLsNzettDUfdChde4H5ojHvgzqkfxDQPDrNp13P2eiHZNB56jx1aUsrT
gEpi9MbPXXwE5wdvJ1UKK8ZxGZZSsBbN6SgS3XVFG36A4mLtLjqqvZOc0MirGaJLLmytovhZvUuI
Bx9Fxj08W+EdVqu0BYfTQN47BK2NwzyifcyU8aaRDioHP+VMF0eMqgpLreuqj3zMYs8e64ZYx10x
CIg5nyq2r5WnmUlerSPXDuLYYayeQXnrnlnf0sednROl1SLKlP49tKIadFH1VWEDruxgxWcantsY
gQWNCAxEsE7mr5fQ5ug6lMYjrRXFHZ4GaOulfp1PNhS/ldAZIir6QkZ40f9iijDkXDPmxHhtkggK
mau/epca95c5HQMCIHhAtrV8aonX0ohTMYR1uFVuuw4YkWYftlJBpS/rcyIYFi7H5LdsrwSA8hK9
yUfaxzPa3iylidLjg8orKfPz/HFYMliCGb4muiVE7ck+mPgssHiOL0Xm8WCKqmaw01jFccEW5Bhc
O8wTyEjYYTdcr2ZN2Rn3opht4W3auNj0bioavtyEwIBuB7L2lb6LsfFUol2DHqOKTG8R7FzrcfKM
jsuL1Vmzkcc7sZ0MNH1UNwSMbjwTwArQgimeOPUfANOeU6qEyseTAw/dr57dJAoNFfsf5e+KPZvZ
GX7pvF2EJTX5p3ZGpK5cevIfbcj6e+Zxwdtlw3o+7o5bU0gFaLzsgXgohbkXYqd6Mc/qbzceR22J
IGhi07zjLWvynnLNRVyyaXogoh8zoHUmU/ADPw9Xnmdkh4JpxvIff3DsEU7NNVGpJi2h+ffb4TWm
4eXXLU4sfqBS4NZFe3l5iB3c0xscKcT0zTsVI8KvPxv9ELRAMsAq+gxda+VTUJU8GMfjjs8XNhtD
xgGlL2h9Q7+A6YwnDlOqGmmRbBQi1vxD8+7Zk3v20+jDzmgeaf+V6JUJCFR4ADXF3qlFANpdk+X8
XloK82l1i1ZfBUmLASKk0o/by0mIzzWVnL6F8z7PE11CABGTP6mJ8uex3BrQ6QDR/XPikFBMSMLf
Kk8WXWWxD4ZgOx/Fza/dFrCvSTeV1ge88RoCen5xLw0zOiXkW3rEJt+YEwUomSLyC1EXeU2wqWpz
K7zw0Eyrv2Bv8hAGvNHWTbztaBk2hnPUbDwZVDDX6Z64JQtjzk+/rbomZ6pnCkKG8mVipo52oGGe
u4Wpg0KMw1u3FCOpvNWS5KT5yZoqOkhKxjEz9xwmnbQ2xQfEM270R77LXQv8g2CiMmxeqxqw/mRG
eKdbRLWzKGEjv++k2TBB10wbTQw5nIZWW16EkkHL/Yc7h6DCsjabtOzCrMjNH2pImReZ1Sn3CfRc
RXB/x65OqKFy9BBSrRDX6YbwkMA8/tAx6KOxr//VXtBCa7f41Goj+xoHvvHtpu2kBisK6WUVV1r5
FG8klhr5B3MLz/8RbIwnNmWN6nkO/3fyO5qCObneGFaZhoNhNwRVPDJdJ7p4sUiU8ehawr3ymDIl
VnZElC4B8kBbQHmRyNSCGQwl0ohkgEmJoDfgwOsu6nLEvFUb9xl5jx5PPZRckHtU5kVxY273b0zo
Cg+a2G/DKG/aiUYd/GjRtaquZNq27fI+9CwgRnA4/q7DiDdHOWy9CrxNZtIaWhaWCgHCPqGrFc8C
E2Y112L61ReDgqUv0mcX/ttwpeoGhh1eiJ8JQrYJaNUizsZlqYBzLEU/2/73rpunZnnHguPBdSw0
5taEUiaxT01UrFqfMTlJMiIWxRcVM43RsZfjfkcc15NpayHev59RlC4KmMnYvDiU2SacoVhES7e8
ol3Rg4aNp4ceEWl4J33sltRNTi0FpPLdrZm3A2dBs2mbFT5N3w65BxY2B6F9It6ag+5X5NU16m33
qFVb1zzfdk5HYRswL7PL8DjAvcJsIG9aMSjdMXP7kC7qiS46U426wVjxo0B8h70YlwguE2XYeNZ5
DltN41ExBtmOoNIsredf1JztZq5ZXaOKKGOYD7GVxo24m7588qVICLTVY9Zrn4a2QhS3fTheWmXO
YaxHsEb5xcH5xVidTtD9yjJIVEPLlKb16VoGBP7NIAuXj3nAI4EtCLEJc+7fOYHB9BfB2yUR9u1x
8itK/BotWgcX1xknhDBRkca4DBaUUFDPKCwHE0nA5U4qct5nm5p9Y7jgnrH4++13SZCFj4NvLfN8
7b04ECd0WIgALTAbN47MsVrLyVhtaW5ueIVh6Y5UjZd2e20T5Mi6G1TtDsyM5id0Lgb+u7vaIwft
lxSrCYUZmlMWy5vZvnCoLkrWTssF2po93Z3GX2sQ8cKWKfHeH/aFNLqyL785hhJVZGTv6cXUtnO+
i6QCU0BQUFY4o2mnh76DlF/LLEeZ0qJz+8a8NJ4fc2Ev/S61tDb+SMAHRGeoWhDyn3Sm6dFZG7Dq
6g2FjjTbuVGINYrjD9q7Q/9PXivbxRc6fWnvMJavC1qrM1pUcTwlfV3mAkLVwGl/qgPCUTpsbuNU
Oy3iF84/qPXG+gniq4OH8SzLRMj0/Vt8nucr/TMJ7Zb9p8wbj6K79XE4f/6W2WcqbElezXtrFs7C
M+aEpPwtghEGxH+4vcl3xS+ArXaj6fJcbyuvBnpAHCMtHh2XXh8x2Mpr5NC0EoQ1Y8K9dSW3JXZY
bGP3IohVG5ws+jU4QXtdqicEF9Agh88OVVZ0x+bbdT4Yl8i2U8qBXcH727D6aXiED1NlcB8EEo6+
mfosmlYv4rRveJpLt+NKovX/SnuFzf2VXMOfxik4flM3pdA58/jjH7iwSKekL1ohaExCTjc1I+ba
+dsDESiiO1eQpKAq91fiTb/2lTTgo1+r9lSB1MxA80lg/V6P6a6Z+BKvSsHo4vk0WLcQM+8BghEb
iYKfudFx1/QcoHBT1g4fJFh7RIqkCv8HgOAEDOw53Cdd7obsNSZZ3JFqMVmpT4Qyqc9UNWInuoUS
35x9kKA9qlyv5KkGOvvWtyMSIBOlOueEGyZ0mmASW7FSbaIfD9wQ/wq+wJ9M4Y6LW1E8EkEI7LrY
1VKKPv9jwn5PdVnXtgI1jLuKoAd83+VKw2TuFyjr2VXpNfAPkQpSCCnM6Ozdu+5uhl3FtW0GR+BO
Ut71x0mDeSoRj+nvtDuiOSxZpa7z2XXM+4pmpdhDsVlctLYBIJKUnXCtRa3GkNfghv02Vpevt8Br
jgeb4ck6k4gBEVfZaSJN3qnGoz+0m5WAARYSjEadKMgD1ZAfrSaSBCkc7kOw20Kb/lTGZisk3wlU
94QXDK8+IYvfGnDoYWK/djHlGs1MmN607LvV24KFi7IeZk84+X2u5X16uukRwYdRxRUqnAj1Y6jq
RmrtEaR4Yq7eMOXSLYkBE/8RgHnh9lNpmwZri40C37MJFfzmTIK590IqQ++4ybcMYcD/Q+52m0iM
5y/XU8MUjMl1URWyjWYAt5o7mnqw9sdpFzmQacQjUU8i1j5G1oxez+AQVeW74MKaT//NI3lmrnOi
ijTQUdg21aFZehgFX3iJkibm2UUU8pnAlr9yDjYMtbEFpfzi4QLz1KI+ZFs6ScZ3JupW42v8+KQL
fdmJWLCVKT58aZjmE3E5RtRFtJ46CTgmar5knz0xe6MN/8u+cmNFi+AU5BMtZ8mmoeS0n49KvYW1
74v2c0crHEYulwj39wcS160hKhAfiZrLe5l1V5y9t8emDcbg+IITJTr3P/oHY0/gu6UgHUAUzzSv
1PFt7ORgDyhnAAlved45DofYLRP2F/7lHCYcr2cm8FwsdVns+qB2hNQRZAwFRXc8F8hIoVdaynSj
L34Aq/fwHImQG51w87UOCsZgjI2xXHM8SKPFzP2kQQZtb7KzOsT4/FFKmVI/gPUo1+/I9DeKIEb3
huz9n7V3Gu9jHF4WZUqdJKE+u0lM8T3unrfGx2ToKnK4V2Lt2BUCtjQ4DfpOXKihg8Kl3NH/AfMA
tYoE04DpEiyr1U5y3aVhHTOWYzxwHmvOnH7xt4TcWv9eFx5zIp6q3mNLPL7PPb63sNnXOklbYawi
o2alEfJ+yv+u0r5rcTfp7NOk4AZyuzGow9SImrKb+hUkTx7NJ9lVZe8Z7ntXUfvge8K4FmFIFRSi
o8uGnO4sVJ3UW5leNlgxJd8JCW7XP6n9DwiPKaxQsHLjiZIQ/Yd8ZJ63yma4eWhkl5sG3L5p/54w
5/mTwtrKftcvBVma0fSAvHFE97/DXTzQ4BOU/5gsajhF8JYtrCsGM0+DQYcd452MGolkB6zHn0PB
wy/VSgF7R3Y7jImJbsQ7M7q6LXPf/eDk1FzbhY/r7crkP+lxHpTNWBn7veqcz35LKJSWzC81AEoS
ByeuwEnu/tFBOKtRXmtAZCSrc/PQUSo2GJ8k1mku5QwZh+Iam7E1Jp5CAK0yKoXLnErr8P2z77W8
bdWlBevhpmt8+Q0U+R8Z1RhF0vXwUeLLj4xUVfeSJ/XzsaGgz1jf0OWCm5wRx2U7ezsZ+yV61YSD
lLThWjosBK6RRdXbn3zslusud7lzEsBOYkrfEWwpphHvy+tFvlfRc30KXTUjg1GI2qA8bW9Phvz5
LaJ7RCiic6PaZ5BsQ5YjVslJ3PQh1Hu81aQpXJTL56nlGQeeyVhH29Yh8bLOdQ+iuuHSLkhYtely
q0Vr4nNKQ38fT4yS9qgACjlEXC/hGc+VraQiYA50bfDydzsf1C9qJZoase+z9umBopCubA5VCkT+
sYFoFlq3jxEDjo50Ysk4oXVUVxtnthSYkxLXuWL1N+JTAny9tjqY9/YTUOi0I4bMLoiRARXAhDmY
79+NX/mzU3gd8hzFQRNcsWuyAnY8F8qSCBlRBlC0QMvfPWFgbDXpqGAPJHQ7kLDeoFilQsiTy5rZ
ayLlWN+3MLz9IJL29WU/2VsslsisXtggB+g46d5TtRq/D5umAepXEI2E4edbRyQXfSbVBtour8yZ
JIxgJMI2A1PECoRrmIQP/NH/ZEbNqlA1HdBuvfSRHw1PDcUslqh3AgCsSJH6S4+I/fLwxSBduiA/
WZdJQ875uIfFlB8LukSGe/Zlu4/uedjUfzYocUdSKGCxid/wXLxrlXWvpOiwA6wPyFMk/dO0zsmE
whe26cWvlhLZxo2qlhXSQiYNndtA7sU1yt+UdpJCJh9SQLbjig6CK2K4N7r8QOJR1CN9PTIQcbwu
NLSecutjuEFJddSpDBKoJm/ulI6AGdD81XQ/YvqexbBeyWiTDwOS2agGFIhlKt0VDcJZFxf0CNhy
e35vf1vlKtwCFHZHhex3CADPX3FROJboEY0NQHCbyhFZ277Vd87n6D7D5zb5Z1wLjDmGfa9a20Bf
0VGI4Kj0EQLQjnPhb7Xhr9K2D8NRYzCJ5XRj/J56Dm2BkgLGVtZ5MC/zUU8d232MlJwxjVuZrDDx
fSrB5+01zSzZMeT+rZFxRgt2TqNjDqexvW8QFXDzcY+EsA3pypnhawzrxaZYtPOYKBQbeIsT77mt
wpFGMTObzEd+RDh6RKcHdsqfUoVLHFZxLS6ns9/UKVo5z/MDRDOy9eF24Xu0BBTiEffLv+VAoLkX
VCuj55kFNU7+l6TySf5GvAbYrOy0B0AqwsqcmP9MLEGMJ2efEVjyU4/oSW/AfRmuV94M1uHnbu5V
VA17ebnhuzBNu4UR4eIzsOuzDbqANtPKxMUrVTouMAcTSWPHxFmrRZQR08Dtzx/JQd2gQis45lG+
bUifTVm9CaS+2gFUcVD545O3osXlHtrvRYGZ7GGoGZfkCXboYEtT8UrJQUP0vcHdmRx0pG7Xq7Pl
DFVfi3wi3+tCDw7TSMOS3MZ3s7ynRCZItBP/EGFuAznWdh0TRhIRbnvj5Dzpt9lIAWolBWmoipri
hhgXaCZdRpIWkt4mxkX7gbJ7sJAcA9mP0s9S3ID8p8euDlB/O/Bc32xEk+mbjT1/uueng50k62Qp
GgYYkYKhv0l6M/iWg0KngZfr6jokn1lg3+Y62Z4WsYT+vIuoIRSpqfbBmMQGg9T/4TdMzhawIVwE
LeUkGE0QnulMsT8gponYl1urDc3DMAfqGZxogu935YjiJvp7ezcHq+FEh242qSrRbm0xv5G9Ms8C
M7Ju03D5G4BKZ8NZBBuQWlJJBQZrXw5hcRnQ4IcavravXKWGdmM1ACEVtKFU3RG/M0jry+NN4R2U
0MC8wszwUg9Q418M0OGxU8o32eZahz4NbPBQOfJdlU5CZKdmWtp9jexFvG/BZwSkepST+Z87Ye3A
9dehL3tnZOJn8oCTbVbqZ12QrDek+Jpge6CTFQuLNpAoW9oNboPkor0xSEhYyqdshDFzzE67f8X1
uC9KQDDHhH40b5FtsS9dxoZAyfmypvX+KNTGH7xslWrLgJhRWyKY7m4TMUIA4P1cC7rNI1TeQXiH
HUFAqbFS4ymiGS7ov568LbIbMjBY8cfvbjKE5dsmHmxoyYejb1t+8wwAKABKrcQBFR6ou4XZVjZo
250HBqXmF1xOG+H9bil30WZevCf3hk9e6AGbZWR/ewsPh9GVLI9/H46oLYuslpWTDgf7m3Z23/8V
UlJqOS9E5h8j/+X5jp65H6BX0ngQr140MfrnfRlFj4+i63fVf/1vMQHhQoyco/6B+FoR5AdnLaEI
2RmzYJJtmgJfvd3MuWSbsqWPl4jjlDsp+aE3YcWjbvjQ32l1SySCNXkhvp/meLdUSMSmGIwoA73L
VZwXT8qKz/3TKdSJ5rzaoeroFt4wYSYEkxy6bBXu2hY536PIBXDefA0zDy9wJHwJbRacDvXXnyeo
LO5N4haEF2hWd+tfM2WtTawFwXCM1QddYa22xEvdK0SNV+VOAEDFlS6GNajDMlNUQhoc4Qldj5nW
ewGa1wgWAR8khwx83UqnjyxVSdPd+ZjYqc9yrfTp2DXS8fjta7VN7R4flroJyjQ9/vu+oNtDFcm3
vcDD1Us2TdYcS3r+8tqN28+uTQtecuVU9p/PTUpf43ENkL4+plz4fqDQ3typPBSeeCQ9jC6a0/8F
O2/FB0fLG1nMBWAkmkVqcbhqMOK+YqOGXVwwLOPLEXdT49pFDE00KueOmp3GGmfPfxA8ssYnzk6f
NKhH7dOW900naNI14SGXxqvPDMoPXM7RCi4VyeC6zOeh9eIc9S0EzF6MitWJ/9xzPuBJJxGivcgs
iLuTDIyGl/vQctXyoiAD14IHVWqaQZzmdFHhoxqcVUdxaigau2DtMPuApSDpurXf+VGj7GtRZxp3
5ZiPB13DaroBg4rI4b7nlK9k0REkOW57wy6/2JxsZZ+yp8bK7b4PjgBn7Hjw9gkXCmndfXTn5VuO
m8w3s1GyFSLbseDNohk4OFID3xfFNsMGhbTiT2ZGLJ2nPF5uFU0ha6lQMpZRF7cbJxXZil8dcyAh
X4vEJm6yMZ+qLyGxsMm5yzZtXnfgvvyVx3UWB5zRRoxN5JovEINKdsZXRL/+C62OURQk7aUNnEaN
HJx+mgyXwH6E7EPyg6KHITHngapkLTqmW7X/6fugwMkwhIjeyCGXkyUoIAxoK8XhIE/2WwKV7sLV
4gn0zg9i+QPA06LA3tI2txUzMK+pZYca+S60J9ThvAkIZt6LgYJeu2pDQ3oP67mI9mSH1autKdQ6
ABGINfDx7gOhQ8B+d5+rrz09dyGP1fs4OGR16cNaaLit3WHa5WvuJoMz/QbE6iWT5cwRVkleMtQq
gJGLMcEh72T+BO8uShBufeaKckmqy4wH6nbAsMNqg9QfpRuJRBGq3t9/DVJo+vd8T4HHiYSgafAk
aZB4nIybdDE6i1tYVH+3DzTvZLyX2igRfV9pVRY2D2kKVSrT2wMje5VIGUhcis5mXaPnb3hUp+D8
nN4xNxj/Nem6WZmKBTFliUf8WS/MHNg6niCititcCcCM0afGft7X6mSmeyWA3WuXQNz6MFbUqKaE
F3TyvUR/H7hV1KFTooT3stPKlnxS3YQlh5zv4mGNl3N5abBC3ET0LpNXHOnPogyNY8BKNbNYfPBq
TpOwLZjn2BalT+zRcYMwB7yKJ3U/Hy99uyHYLz2VY9iih2iNVMslrI7vD7c5mqx28/slTJPFjtay
o0Ppsprc0ZSbZmlTqDbkboN5aiAn5SJAicrVivJ/qPVqAvxSszyyo73nIxM0ogLZVj+wF8eJb2gZ
NeA9u2b4erm7URSPRGVC7I9nJeed/Qw69fz+mtJ5gwAru5t3jQ9yPadEMBryZ1Yhd/ZA5HlLY5g0
4hLp0jy8iV0ZY3PCPZrEwYLTvxV3Vb5yDG59bps48aGQy8rG5tXhJKuWwzOIM/lZdlV/6Q3KeH9+
iONi5RugqV6R+e7fkjXQad6zpWSS2zWOMBaWKNtK92Ixtmt0fG+4LOwm8hawmP+79R+eTEcVrvcw
Jh/Qn+OunrGeOKxVYhsXw8GkL7+vO/UydJ2lUtY5x/QOizTrwaudL2WCB6/spAVDF/mA9hWy9y4z
9vbj1WJwa+SXCZhB82qc3H5dt+Bd13ODUFTYHEeYMb8qg6CPZ/UqmkBJaMehlMcAets5/rQGIE+e
kyWOMp3EOwm6A/3Og41ssbzwn+XN3jFqjyx/tb0vX59s7ldXAKbwCYC5vChfsDfahO841m/nxBJd
J0Tz2HAdDehhFzSbEh5mF3K6oVbK8SsRRCUDfuIP81dbRUf65uxbygMd0nXRG825HyL83kVXYyIp
H3ZUNM04WgWNm8bHsmvjEBHI4DUbpA44a5wFRS9xjgXqFBm82yeO+m1yLq1NSChCF7Hg5YavDS7R
E58l9+geaqg/PjvUGRHU0ats69N+00sZ9vYylmHcxvviOwB4bu5/6VoOvBIRTBoeXAkyuXQu7lZs
WhgtAzCRYSaU6N4rylLhehJ7ARiaSQIFZaYkf9IIhoBso64ouUek8jG8u5R/y2bAvXWcVEIQaJF+
aPnLcwV2HmcT9yYhvj8NIj+R7cE+qAOLamsC4m+RaR+F4m1jjXHV5dX7DkmAi/xz79OMTeHNBMrg
diYOPgTqGgty5eaqjlbM3WqY7VfE+Twmd4pLNQ8RNHxz01oUUaMzNLl7IgxeIpkztQzcEW68mWpH
vljkuw+DxpWezKszfJw8P06ndjHot/r0tlHM6xhuy6RrXzBEpausJrIZVzZf8+KCBz+B2gQr6jVW
LnbRpOJEy6kvw5b87Yf+swwp9ulCCQXnBHM/wtNHcTa6HPaGae5fvS2mtQJgFCdVGChNceBEsO5p
Kw/wKWbFYAQ0qQtDufC0+lPGAvPFMCzHVXKg7bkWYPhVkhL9/PrrOU12OuiJL/9S0UuDfjJaj4Bd
qbNmsZYGFkOelxJuvonqv29RxrZLcq1ofHxepNAIgS/Ixa/4hRkpewu4W1YavhPE8qw1mDOKy4nY
VVIm9/tbHfViqFCE6aWUEal5plKrs+UvcbWAHaICf7R17+EsKZ7Bj+IzeENvc/78kF3Q1nxzk07d
hEVI3CETyKrPGwbbtaYePQml5hTk1yphwyM4DzeWtFS6gCsbpscrRDEKwTJJ41T1Lo3nkY4NuCE1
Knlo0I153gTuFlBS9644Ri3xY3Cd4c6/Z46GwtWcChZbG7Lkif0UO1pMYlybPkzgkDBUPjoC9ICt
NTV6iTaltOgvFq0I4vxkAU8F3npkhNo2NBBI+ijb31UZ902yO9Y2L1WwAdOVN4KIawUdyr56+yuO
uK3G+bK/slkApBxDN0VIbAvN+QmoNmYo1txvcjswSOVrYwYbgTOko+j1fiifA/DByjpSfggwdGiF
n8AiH/Z46y0eZ4kYapPS/Elpu3SBgoMqD69APBsPoqAo36meHWREMnIZfGShLSmtYKD5YlPq8dd7
/Mr3OVrnN2w/Y40gFubtYjdRf/8pMDmJnabKn4cWByftaSRb04Y4wBz/6npa1hmVDSoDJ9gVKvZy
JEY3JI0mli/bSXxGg5nq8Kpc7e9Yh0dB4N0GEZnBFfxnKEeE+VnxG6fOjfm7JP92JLHqBIvKZDEY
3Z0TAIwY5yBcTEJBKWd715dMzsYaqtQjE7OnHPg3M04Y88EJDOy0YNoYYmciXW7wr/Sfvt63Utyn
YviX5NtsrbaYEItGVPNB2cmI8tYf2M8nf5gFzY1yGezY1LvWxHQg5NUPpBQzAeh1C4yqONf6F2eV
tORhrhO523WmnDeSkCaCWzI/sRUL17T0zBw6tpIC1fAsl3wWdCp74IKm8psimYb4NSr4qqTuEbzq
HFFz2XRvfZZeHW8OnSCUbEKZkveqn4FnFaAfy3Px6A7psTfJ5wV9oAt1ITnrbO6C0V27WOdknKD2
D6ihr5A8lcUsH46w9mNzwtNBAveV9bTRHLJbqVXsM0bzR5hIGKI2eKYyE8RJJnlHtcO2OG51GNQP
Kb9LvmHftTbQdQw7W7a4OqKOAmGQyrTwZxGXcWPnbSDjF1lobemi1IOjGYKIET+LtViTmS7CA2uN
b7Qm2roX5gyfBuEViypxibAvKcyhvNHOsr8LbDVnw08Hfh9ca9IHErO09ko+bJTnHPaZjNO2RblY
PdQNeoZwoo87dTwG8MfkGCpPQN1vhrN/wvgcS88STe9cQrua64+uU3mVvN0NRqT1JCckl1NT4bD5
vgSPfabRXu+MgcgaS9CxpqxsWFfzKg4J6RrffsqRtq3Pwn1yhnkNJLwu/jwP8VJmahKQTNcLNFgT
N34noWSBzrmoQK6vY77utXzk9n6ON73BoaZpqnjU0Zu+go2F5KnQrgbgSVpD0eeGYKyWwJr9gGb0
cUaEAeiJAgjh0L+EfKS7LVinx1cBvvqQ8augufVCELpWMDnOdg5LI7oPxC/EsS/bg2X+fqR7g9II
92ZCqlH5Al1T2nafRjcDExww3qYWtSGv6IziOwV7J5SGtSHM23rDRZmy4xCvXsXCX2KEFSmyYxr6
ZjVh8AQcdXPWHOJcdlHq0GPdO7Ja0lb27K0bikOA9FEQK4f6EelK1u1Va+p0m2Wy1pY52DU20tmn
/C0Evcnvk8Qp1kmbADRq4uSYgzCz/26aYP3icXg73GdfZknEGceJaMmi5sXTHhKNhJ0yKlBaFo/+
1b6LXCvdEbHsGfeWzUdUhyudAqp4NZ846Hg3QxqpCbJT0aSHqkcOLiennciXzvswDOve1ixcR7Rk
pmwEo3RUy4byyXizrDNKA0ISdL1gTuQdfLfCJJ2bHvIj3d5wrD0kZJGbpbaajB/DdyTx1tUeU0zA
34RE+bAM4ZkUST60VXzPdHQW1hZ68zcpbs/XH3MpJVabiIWpeHRRHIIgtyaXyKdp1CGCHBs+PCP0
h24c353sfNgCxawq+JT2+nYSxS+QSoqsecorj+870SXreV5m1VYU6r7m//5ERMiOURfbfXjuxxzf
/SY10kyRw8nP1rihhFbafVHR68phGCtMJuAEbGtRT/Na+4KwTEGOpyOzzHnE+QIovo2oS1XsMMP4
QLAiPa5zIQY5GH/nvRwLYB1QN0tBxpZgem+WiJ7ZRHTtocX7heA5ERKdFmnrYHNfTL7T3EQ0RR68
SFWp0oObBDCZLXFV0Ru2kK6dyS5uhW8Yb9V1C7SHrG4/c9z3SPHnWN2DZsF5nUeI4xr3JhbBwI2Q
+gFiZgn+/0SkCBHeKCzCaWtjVYoN7tiL8UEosgZKpxYG7pg0byJazeLxDclUtfwTyqLiw3VjKHuK
jw9EQl7ELoaFJJ+0jtrR5c7OSRZ3HKeVzheR5ffs15c1Ni8IEHmYXG3+8vdK3UGLpfn6/Uy4Gpgs
bqogPw8nnDk1tkTCO09f346VX+POnC63TGfrttXnrWaukyiGwhjcgCnQllfVLU5PzsrGkAPJPl+N
oe+A0z7m4q1mbLQ5F5/eSF6ZqXxfjmHkgD+FDUKVcTRRn+Rbck/1CXNQXDubacExOu/5YpCiYH5a
oEVbmnsncyA5haoDv8+TCWOqBKnSkBaK0bU5X1kG3WoofQPgj8f9Pe416p2mMmOLNZ1V4ZO+f3Kq
eGiijrpKP21difXRu1fEO3mVBXY7llIe7Q/mCUQwBdHYXYHQfm3A2tC3SVryT3vcEZXNKIoUpsB2
udJ3VaZxiYCOXMf72b24yB7T9bTsMd87uTZNEF/Nv9xxhgQ7f8xK55fJfKp3OMMQj8/74EIulkec
QRG1+N4hjO11YgVeleG0oSeuyfKPOk5Dl8Zs9UrOdH9Sr9UFfv4iGi83Fh6a75cNoa/cQ/i6I5lv
hw1cmcClOyBnsFOHvR8od5Cde6/dzSorM+9PGv7pnQP7fn5Zcj117AWcqozKUPyTQepjfTk2fIW+
z9gI3qbbxjkTuXmxYARpxdTiOGWFYQLQvm7NwI+XYmmqJ1yVjnp2LawaTat0vKwy4F24nbpsYqdT
ZIKi6LKA9frKzYL+LJrKDKoIzZMSCDCgQujL3t6B9LUmdAtc8NszFW/MIqwDshDXWDqDr5Ku+sR6
f6sYNB9WpCuXUMyFYMEmNKe3i1c46M3hW4UvpWaEAYQ3V2ma+w5RYHWeWwEMpJ9wpaMQth0KrHIm
Ymnfoo9ITBgVRud5c1zgTr8ogwblSj7ABXtY1jW0APj3diGwiOg9Zxr2Vo1m/n/wXgq8vjs2Gckb
qZAuJz4VMIWv3B5BFM/Gi66HLtmISgnFF9IBGAmeEsyF04pzf3lRqszbr0tRAsv8ikbQ/fHBAdeQ
lBrzLVXUaNm5xWpoe96cdpMrCrLmBb/hSV7A8qpthWHihxsajmGFw6F/s7ebkrYn45Y2GPG8z8hg
LWWOb/j8idbx0x0/zRkBy/C2VFeJ+l91JkuHvujpgG9EwYhWGr97Hf3/BuooWTe57tYcUo1p2BH9
AKwOYnbbvwvLF651MMW4soZWjg+dMUmrLBgV4bszzX+ILmb/IcFUZzd68QmfN9tNnOzfzE/N3fFS
uDUtm35eE0pXrKHPhviO1qR8jM/I54+PIBGQqoOtWTxRyWmXkolxB2gSqPxyJySAb12D7vgPVtiw
F7S5mYZ5Pnn9rxLiwlc+iv2oNxGI7E0n0UsiIpw8n/zeBtY/70D6ydYFd82ZDxbSNGHqvMG7umTZ
8MceC0XoxLE7aVqjp9zUkAT8KVuQXS37qT4YYkSChIqjNkPSf9d5p8l75ElqB0w0sCmhoMD6Zr3c
84V7nURW+RCT4nYOckcUF2neDp91w8eJ5aJ4lcJeZ7pbfE8FjavzJrq+bh0J1f1dw320n/KK+4jS
9AaNyLqZREMedRAt4ILl1Tl+p0Vq4y+FmTOaOs2sSG4yzXcaPUUltyM45xMspyL52pYsqD8F/JPL
iy3VQXfpn05q8NO71syErCQncbE59zBGK9l/7NuKIaCCYbFCFMXacmwivuouLNchXZnnhOsfaJcd
pWUpL6rEONg0H9NarW5COso5Ts8PzXYeS2tI+m/id3+3e9IIEgTkGjOQlVfgkxyRGVR5AV1sAMwi
spCeLX+27v6yDimuKqUYqDe/PEqmwKoVJCKwDgQmRPHQwgu6py/d7Ayw5xirWr33sle18I7UtdVX
nx4MJbwm9YlBZEWixhUHkMowZodFaKxCzcsRIa51xcj//ajQFGTM5UyVnH6gfKf7sIZS35lzzgCj
xCzRZUsRIs3g/cdVfPtlb4TsAEGrbffVEbk/0Y2RFc56GFq9AjY59NUaGcLI1Ljrab3nTNugY+Yn
nrWB8hBhsyE1oIYZxBCi7CAmmsSjsF7fduM8tRSRn3G6WX91bmV/kbnrt5ONh/ld2gQg11JpPVqO
rP+RrvqNIzz5hebiTUXhRRGavA+GCIbw+ULj9zi3cirgg8DqCuhiV4sdFTaorFkAcRvZjl0Apg/a
+Zmvypg3ADntEAIuk8lJ9L+NLFUpcA6j1ObiEqIfLahJLxAUAzFdtp81W6m1ODgB0kiV0ucBnJ/i
d9QMeWLCjyhifmvr56PjsEjxTDP7Zdb5Q0Uq0GkCt1Z48oK7Urlg6l7vrpVsMBudlldd8fnPDUqe
UuvYqD+CMyXtCrH90t38TL8rH2us32Km2wHJ8sfPaCAZE4PUkUidTuBAdemLzFCHAlgCevn0pkvO
2P/PiIq+YuYRPsI9BneN5f9WYa2WF3BtZTGhUnIPsMBVZjbvSHugTwz/QlB5y76mKmf6UaxLbT3j
HakWjYbyLsZMq3eQ5zaO7dh2afrAMnw3HmZ/m3NnnmJ0DQ0lvqVMiMtttj36ldBdAQ4K2sglzq4z
7V18CHonXFfzumsE7GI8FoMPoJ/b5jsBrdYHJScLF6Srk837xlnUrIz3ib7/Cybk/Rkb9kg4U9w1
sAWRPM3BnKYOSxcsgZumCbYf8RibmmbHtstf7AqbSmtG3LD7InyvAAXB6TWC8NP1XKIqYjq2h3Wh
qFx7CoTCa84eoTHF+22e+lb/aA1hQIYpbrimqUg3XyKY620itWDZcj1p+LGPCXl0NXMXJi9H4SSq
IW7z/rfyqljS6K3XEj+la5PzuLv1ggR4zt3KFLrbnKJcvX9RFdf7iwmj2+qTs+6b6+sTGklDO2XK
0/3EhZaikkwrWoIS/IQ2dEfdtg2H29s1XieATJ05xOZgVdnib32uXh9Dea6QYUUxciks9K+1Jpd4
c7/t65jt8pY4RZzB+avWxUon+37NhPLvW1gYVkC5tD+EtLQHl/K9qiKLwf4sZhWSBFq10nCtr0QD
t260nRbnpyWITk8M32ukrxda7Eg1Z42hwoOnEDiUKzYtffWs7nH/T9eSVDF8kmGtNoGQd4G4Llg3
1SUA1WXRCM/BHE17/Rmjlo6evmUVkylHguqE+AbVWHSlNnUs18ot/INEGOf26droyXGgwWmIqFa/
Cp4ZfFK7yGcmi5rn9PAk8HpUD+/DN82fOG8x5Lxk+3xseQJkbidTbRTu2FmOgkPQVKAvcW4b7E+f
JGPxKJ1id6jLOtw12IK6+65GINWXyPgH1FfbrqNcj24lavQMmjoAD7i9deU8tgPd/EZo64yB1B2w
+xQWvvfXbowUkv4onMWTGa2vVne5DWzc9tzUqm3CFxMje1suQWhL6oGP5gBaOL4zgGmV+ODizRwe
TfmmqoZRVUEifcwJgOs3SyLONTcPY6OE+l6dRVegjYgCK4HGZcpftQ5OTRUs0bx899vfce9ndJRn
yqkV6HsLo+VgLGjBNrAEQSV3vtMsJsct9anj94IDHHI5hx+6heEOpQ3Lw4SyGfITAy5IKnWZTmRq
ivOM01HmKoUAsb6FIzoeV361ef++InFqKSR/Hf5pvLux1IRJg3hg1c0S/Mwu1Smogm0++vWEC95H
VDjzKM77bfwmWqJZp9Zz8QAAJOUh4wAuZcxvpxPZ8qu6MAUD+6vtXsb8oypXVQR6IFDUXNFP/URq
Af/NTFHenjeEaUcm/uUfo552E4UFw+qgoMSpT+KsCj9BjkWO0cn1+A4+zJ3ZbCl0vgTXzznkC0Zk
XCPYSdXGqClrvcRmiOKZ8Su/D7598PE5XE58MPO0qbT1KJaI33/DlxMjK2fHq86HLDoBC4GqU/am
V5NO93I16JfN7Z6ZxVzygscopRgy78PXnOiqfWV0+PjqwTgCWp5trGmz9C79nyf5clkCLdanG63z
bjk+MI6stiMTAaTdGrfPfcvB0wFfDLaDA7/BYggROtjdTzstV8pCkKwKdjD0qCyI7qETz8BB5QgO
kue4OBvZ/c1WMKx81D2jWzzfNgrOt/tvNzeWVaNgHybg0eUjmLnnQCxlNUYbhkQXKHKVyMavXxqb
kQWKNYTDOHycI6hUk/U6D1nGtw2dM9qsbw+pVWVn53RYFd/u11KPfq9ccP+ZIdtTKqi7TZabzS0t
034mXUL4pfyBIFRJ5XhjVo4g87dMi/1TGaehmemtO3nwPliRZr7LO2Saq9L86aZTqF3QhBBOkJy0
QwH6a5u/WAdeedF+4gwkOduWvS7zrdlw2QLph7WV+5TARRZzaIGwwjXDheyrXrsxz9NZYmF7hVnP
sF4Ay6xCgE1e8ocqHHSuM6M3F9CwI7WsXb7ZPlmVT1siadmPuHdxXHgxlcI1GEiHhyj7TTUXVcF5
rcnkMMG2zEn0/jFHak6TDH24t5ylIBg2qIf6l/UkspUWbjRiEKGDhaBDjyc+zNTk/kx5cbqPsgUB
Ir5YzzzSr+zmLaQOd+ogjz/lE11oLsO9yWjF6Et88pKLDlgXiP//T/eNvhhoMN3uUXfeYN3+nypl
XgVDxtQcZEt4LKdLvwWcsK06lKALey++UlqUr/rbPz44Beoatr1Ub24dDtgl0aJbiE1zENj9EZfN
1RBY/QQZdMYk6LfpD1SiZlrG3bavviayyeiDu13yTUdi2qPZtm8Qp70rAgOLQq6fF84DsqT78dsT
LvKwHMrf8LGvrgiCpwE01K1pRXd/azWBDJGqWY3RdEOuaF0zlfvH6pgPgPpiIhmgyXWovUHUa2wS
L2xJ1EuAq1KjeGwYvKXStJnfxsHH0P+RrFMgsS5l0K2uo6uLrh5FNPUxMTFn9NRgXQ2rJ1P2591y
2l7s8o+lOwsIc6BJHhgMaUM+Jl4R34y5xAxJf6gEw6Qx+P3Vr7SXYPx92FI0aGbgTBPwoiTwmlSW
s8SPGQ1tSuL52hE40lBReevYVfDfj7CiXlBDWeg3o5zEnWMRBOsQsRtQc0tcsd0MujRusUSYuNDO
ofQWZQHuV2fjF48Eg7mZiQHqqgiQCrirV5DKmayBqukmKJ9NwM63zXzl0t6GNOabmJKGJQPCC9bV
2cS06h9Qe6N+g0lKgCxoCOaGBNQjihyMVKWxoKQ6XG8EN94qgtqiYA9gW3/7R8dPE/d23zm55UWk
/0gcOZhiU3rfpagw4AwBb5AS1Nz27k8HD+5ytMJ4UncTs06QEHlqSnv8GK0MSFUlM14RT6Dyic8p
R/jy7W6U6YR+QZ7hVKQQ3qj/yQsaop4Mx/qzqFAEH+imVDok9+mNYrKzFCy8ROR9VLD1CZm7N1Qp
qa9aJF4HAKK6i31fzG76IAksbmuZp/cAt4BkV0kcDelIHmxH8AF0++AFIeb8RbA5qR2Y4sRHYbVV
vCdH45e9dHBKgGLeJ93YFam5GN4ZjhNFg11wQWYySc74kVvwDE+qmDVHaLd3GtJ5NXlv2V+8ARUl
B7GXDTR5bqd6KEyo5RaIKVgPAOGoyfOVWGfFMYMjLuoXGr8wy4N1DWhc4BNSa5zsLxsdU38nCzdc
3V4dcbEPUYmdZTO96mx73NUDnlPEDFpi85lj3YCLZ7oPX5v0aSS0Vg4okffNxgNmlXqvAte/6fTm
bdlH3XzwDfaTssfcNsC3Y7WNn6ExrBVCccNXEaX8/4ARpFSszM3ySUUn1Y2kSp9ior48oIOZ/PXG
Kix2vlj48ak70LIiVyhjDbVQFj15YmrywiIDku7XHd+IqPBMvPWK1460LvfiKKjSv25g9EIF1GQI
EhF+tFTQUjzqG+XUv0HWDZlMp6IQiDT+KcrDHW1N4fAoT8NJpMroTSp+aJ6YP1ZUoeRZsqWwOPZh
aDqiNcLy6/M8Bm+uqG4uCQaywvF7TuCbO3DWYGG/WwsRWMyf3msTi4vD+a1ojT//rOQp4XBAfNBk
0WeMFKYaXNrMzrE0BZgyvzsHZKeUwHHWfiw/5YmPpdp5IEvFFjlQPWsCP223aPO1tr7ZZ/pRInWc
VBVdLGp7XxHP5SVG3FoPvS57k/GCtS9Abvjg1bmI8pxMkDPdBJQxGVzsxZcgKEYSGufYfDasbBKO
6J7UNWluR3kCDal8rOLk59lWNvW8nsc2FSEW5javNX5okLwk/Y5SJllPSRQ9vgAFyu/mQw4uMQ9i
3m54roL7O51/n3DQW6UaGsU+szC4QXGs8mH6sm/EGzkSei5BlHSjhP0y3C8nSnXD3jKvzpLkjVEY
yumgti+M1Bs30T9UFSlEJwgm1m88Cq2SATv5fURTxMiyds+B6rdMVSXyLFTDEPeIA5JPjZjUGU6P
YD6k8HA/T7qjFf1fK7fpSi/EQL2FCn2aybxVdmy5j82VXnIGUfG7GWy7T1tLosy1AuBzQ8eGfLWy
lyg73Q9gol2mazyoZRZgtaP1we0mlDQ/IRpfC06Q18KtVNRXBQVGhVJTLeWr7FI0uZ2T0tn+ZEXa
RXM4XPfpOGD7LIruITNcR9YJLafh/lbfWL3/et05+MknVw2gjsxGckIEIO0YWegLE1jSww/oDDle
9wMLCPqGbRe8zDiQd/OIvSWEiEWjTRUEE7NXBWpyLfKjTEusIGGuqUlKWZ+1fovk/IVupkZICVPu
XMzNqbL11Phqy8gOupmG3v5H/P+KUA/SZOVWGLM/V9EdUTKQRFMdURnMsRh5ONgCK1LGi4KZN8tz
/wh1qQR7NIukILBY/abAIODtEFd2nB5KGCwwtqQphyZ5SHXqYOWu3qvWyUWgJ+/7pvmR2EtA83rP
Yb5VLPQhWB9biYF33c0RY5ytz9D+bztGsrGS4/wmXjZRZz398WxK3rx9Q8262Vz/1U6R4tF4K+2u
Eu4WcQgDirinYDdgMS1h5B7v4NV0mRWr4tJn8accmGBxZNZNxTNHa73wPj/p2mL2wI5FVI5xSyGb
s+nFej4vTPwNifteLKjpfEqJysH4XgAye/WzmhSazqRaeUgLoEqbY3TUghQenLoHmsvxvll/2W9S
DHcI+GzoFJGHJrQcZHVAiuoSCKN/DpYP852nIevb6fbw7oYHAwfQ5AeRfy/n1fOeAkLip+X7l7fS
GHtkMNaaFsPPXH9GUagu6rQgP2kH5f+eSBpRYShFtvmSc0dGXGKBtC+O4zZteBpte4YTZMJllD+8
ncJyzYn+uVdt4Gs3WQFt003mm/sdjARVlLUqttcUUSXOzQ+m/A3uLzKUSUq+z+ObuVx2SQZsGlWb
DFIKpI/xe5hZSqGeWjpUaSxphiOU3TMpsElMLXt6NStyCuVqJZS7zXaEz1NCasdl7OYPbMiC2P7Z
PEwfaQUU/Hz5rUlfvFdOyhrk7rHi2yE49D6P7o4q6iMW/A1RE6qsrpFzYQbdkl3JAJbu0EdosXVI
25JsWzd/aIF3rQpuzsx4H2Q9sJt7EWsROHWgcvA9nyneNRT5vI3xk40xcCxfzKzhY2ndfK6B1tU4
Hbc8jpS2D8LaVD1pl9v5ja/xQjl5x+lGRPP23D4/bi0vTLVsCcLYcAxFmit3bXtDve2F3HUV6P8F
7RI3JvRnkqbBFjGziUDUqyuSQwGtCTGZRl1uzes41ZkD/HkPMwLyqu0JmxawgmAzrWbyhAIpXLFB
Clgt5UxGvLdCnwwAg0L9TQ1iag476DkcAKomkOoWJ4scCxQ+1SSoijPMHAfdcZcyhvb4u8euV2UY
in855bbQSVcyu9my4A5EktlLnXJzWsi/s6G9Ds8jRLOTE6h9eRwBB2aR7wU9FLNWRWHP9Zj5Rs3P
m+WwAQL01zPT2NwGGjC204/JtV02ku93tetmoUWwHFmniquDH3U9/2m7XYGSQfKdRazCNHeKW5nB
t88h/AmOCMuwIEN13KoFiC2bZ+kylpW/3O109kigcyxr7KomHCQEcSpN+WQYMbM1DJ9jgTnNDhQ4
BjXA9rqWfZUBIfZGkNoIT0YmGG+9jCYb8zNEF5X/ZhWZHrCdFAfLKD9vz5Wgs79HQcMftFWXVMYU
u+0bS4vN50x06x+W0L5F40lzltwamcXP1aqSMQmfvIkWNHgocrF+DCLdKfvUbjcNcJDO1PNzP/qB
b1VGg2J/bHUQ/iD/ToKL1JaECX+EyovIoEAMYWglheAd6C2sz9DSg2iE6izig+yiMNMR7EIncekr
fejm2I8LikugZQnJdLuEq+/1chula8fuPplfIMVAqigTX+KwmhzrvO/JbsZKrrpaRobiwMPXzZu9
kwEzewtqluUXIGzbLxy0vGYv3IdRYQR26eYWrtmYkqDCSfS6RAIiuOjOh2pjBwdOd2omDDhz/mII
q35T9Jjhxoeg5z1OKW6ozdOSYH4cm0oQrPDnmMmpdQgb/frV50Ml6PsHKHq8TXSO6h0r7StDpSPT
D5e33OC3ct9EaJgvBqwX86WA9N+zdZLtaR90XqIsh7AqVqr/Kx/Hmk5XlKHvI3XG46Fl1AzvxGRF
wDOhTB0/A5zomFQ51Tfh35bIaKAkWmox4YQU1qkyMMDzw32u5m5YDylXw2laO8456U2FcN0xyv3B
DFKF0bhYGm9ViXF7NLbGaDL9dd0NIgCZIIs0DpA1kcr1A9mO9U4dEvjzzoYj8eZVk7BFycmo3hO6
OuVC5pXZlourhh0zAlpcs4cENxQRDoOJ5JEswjBZ3GbUe48g/cCgjWY2nR2/Ro/19yDj16EEJUlr
bmCxrwMtfEPKqEFAQEYq5zq8/7S49sFs5HykBH2aDfBSjx4Z+0Zi8XRMiaocBf6eYke+Awlj5YPE
a1m4J4Nnd/+tr2B9I9U0wGvnkq0BY/IKcHqIULEzWh6QNnoHmDQILlW19uRUjfyblP2w3rh7SAGA
8Rq0BKoRiFUzzEzpow6nTdJAbbkjnz6NjHNOKa3NpMc/xdG1s6o6VogkwDkitShWUZg=
`pragma protect end_protected
