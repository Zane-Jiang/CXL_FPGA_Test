// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HMEwygN+5YJm4UvauhMlE/4Reo1xxVIzl4eEzjGEgzRzbY4uNQfm8lAfeWap
ZKuFuo1aHGRB57Xhud7oxc3g2SyA8srKoRFbrS1XuWrRAv1zRRJnziTSXy8w
u3cJxoYcTW0ydLjZKNZ2R2rkzHO9ZhNLpSISiUE+imISeTL3IDD5aPRU76nZ
oqoVTFbjnMnOLB1RRKTNjh7/glfE1IfC7KHwbItP5y4cBm+7bsLVtElKBX5k
yg0q30baVspv5H1WK9TesxcXHfhMS+k0ZXjW77ZRxjX3g2168GifmUIoGuUe
C1xQ+KrN9SjBwj/ICSZS4UxSmq2sPY+K5bbB4Rxk6w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TFbc6gQ8npP6Rp35h7nRTco5Y6XJq7gEnleC99W/DthHuzskwP79ljb61wm7
Vh4V6DjPS5JJcx8Qlwgb+LFw6g9436ABS3ebgovl6oF0T81bN72/gvyPpBSL
ADFssetREEo3QGpGjUtS2fn1uOM+/0sn/0bKtIFWboZF9Y1pg4CwEatoIiNg
yEXoq9gj/cCzfdRwM5gnjvxHZhqQ98oisyQhYXsO/J6UhLwLg+j+5bRB5VrT
OfPwdn5bRz658iRgDjyJEbV8eHgU1U8qXrFAJUIqwfs4eCe+7lrcszByuEgC
QpQfHAh7Of01hrg42Bse6nwY9pAmTFvj3fhmFImzAA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LuX1uXpbnMUDOCr3ieq59XRy+OpXJPJCFdsHWzMyyqB8XP3eTvVcqro9kUAG
McHFS+ODhiCw4lgprQoIjeHxzrj3QKUrYIuV/+7+bDhK13lpyGaqcQC+OUq6
+aRZdxD3HfiFN2MA6pYRSzIVqgsXKKDTcleSP7iHNZlIYFbs5HOwM97i6x3K
f/ch2r4YqRmVy1RZHB1QgGHghI3eBIGr2d6zEL0g5gKg7Vpz4k7IFb+lCw0t
IXEtHFxnlIut22+RwXD/ikovzRhnpgNqAMTX1uBB59d45pMfoy+AfEtv8i1P
bc6JWtgG9GX/WPjWKQc2nlu2IPJu4Mk+ZeqtPZp9ew==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GVaX/xCX8uBUnnPTQgItREy9MmzW0diI3WxQomgoZr0+YjUAnVgSIplDKWsl
a4tTyEDswFylqC67toRoFFIoiSDplSNxmo9hpvQqfg8dQtE7GHnG+xEjEtSp
G+n7DhIkAiJl3wL70WtFxgdBxUkR//EAn5xe0McL9Lw+tHGyEw8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qosfW9c1h1xZ5ieYAJXm1HbAnyfPVUB0tYW1T8fP2LOmNQVaeiTrFZw2Lv1P
0f4cgUGRJOIBe3InBYESGzNB2T2E3iC9RGA/Zzkw3+KLzajJF8C3D4XLb0ou
IzU9P4oir5K9WO13KOiDjoIJQ8BWzYcqJfMQjQDAWEmZwXmfNzBBRGgheulM
9yInL9gGzRw8d7o5a0vQxvJUjTdVQrL2hYyMp2vPtB2aHT4x9Y++F95BO2ks
0nkImgTOUxYh/U/R++nWfXoQcdlXpm0o5at3veZVAd39cMfkyUB09B74poVi
A6HxD67jS9XQ6ou6J2Yjdt/OtLJccsxX9zeHFP09IB9os9z3gIqFTtPUwO+j
x7RrN4ioRJyfpKjYL8Tw+1o0z7CLcceXQLuBMwk1tQ/1S2FDV3+t8krN2HlT
jK/9pBvFKYh23kPMiZAGM4alzUh2m4hfsUiGHkMOpX18jNz4qdNPog77zD3z
Wq7FxNnIwOi01DZ1UKmhxtqy5PQn5f34


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oab4Wzg4CguSCIqi4nma16TySmQ+G71t8S0fi5+PtdbfBpSGJ83DoThZNsPY
gxuM6WPByIWCQsz/vwVD1HSwXK+Zsya4Z/J+0M64CNsm2d7nBn+Xbr1uJyZX
SuRmIj86GVGvfKDC2GOLNuTMHMV7tEDNMZelKms3s0e3boyi8DA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ktXTH11PK+ydKviJhhYZoxoDrgJMZwIM8X2TN3wFUtmfTYAVcuHxBff4RL/K
L5KQnGdcROkBUuCkZEH9YZxmKHAzdr5XEFfPbNk7zRAGz7bB5aI5onMnw7Hg
qK44LgKPedjs8Ii1oYDOaJbEhfhs553f0u1YAHoBhskMvTaRt5M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1232)
`pragma protect data_block
OsY5q88L5TuJFHsPsvhOGCCS4Azawb7Cn9JzenTvLBCyqUai6uKfU7SVIwrJ
fFqlVRpV1gfId6bzvrGEnbb8npnFOHYrfmDuk3l+Vkvo7zffuNG985EbOqHk
ZDm8x8/4G3RDGCPgtAZ+f+umWL4DKUQkGDTeKumyWCVgn3X618egomosE3oy
sFAOMxrnjhf+4Im4Xzz/oKOWxuwf4M4Y9FFWvkBb2POdzkON/hGORoJV+cLN
VsNbjI7ubmtZaMcaapnJ3QJVzFPLbPCAe4rf3grFy868ReNwjHvqXn/gUFDr
T+EKT5T+zywok6MoRacBbtiy0yAIu2qmlWi1Vm+0cYEunPb/LfEjF4JXzTqD
gqlQ0y+MvxV2ll0NBH5NR7D6Hj3KTbw4SlsBQdYgedCYwaTXiAnvw+tg6Guf
wsx+scd92bQNIssV0KdXEdMvZKlriMqxdnhYsVeOynxEuzvB7+dI+nE76oVJ
a16uZ6xed2lE4m+esZN1aTRe13+WNPEp/aLKTrISDLvCvqEq9zaZRklMN2a9
hkxKRi5r0le68xtBYyj1r/G1Rgh24SFc8eZIW2EnJaeOyUwMO63mlAGCqWgE
qCThA0fhQ6q+qDCEk3UHVS7MviFhl1ZCwyCpkllIiramufnJNj02zpZYAY1G
2J/OCDCpv8lo3vR2LIn5/j+aij5JNBra/zz1xrmws0D9BOeqaTodc1YdGamT
bQ+uifAEte1zVqfSIvf0hO+z5Ipw9FQIvII5qKQ6MnA+Q2g2EBccxOVA9FmE
B6Egfs6HF+y23ByhEVWKO8Zg9mKHmm+AqS+fgQdAfNUfdHuMaUVA5dNizIdS
eMLkMy4g6DfJchL2hvXPHFzQneyNex61S+li/slGREyN8bVoeyFjCbe/p3Jd
9wjicLpP97Fgctu4Iin8FxHO9XnJfDUDU693OFVr4NJAqOB58gGf2mHkE/eK
33kBlhxlBfAfYezHrcT+a9LUYTZ/buzD1tc66wiZ4wPGzf8H18WVRcKtLkfy
Bnqrctjhhti6a5hYJ2nKWGSb6Lo9BqqeGfVFyRIlbPJyfmy6M/4qPbmuNHrs
orjB4iRLP/+iHhc3NRHPNshwYf9Qde/unPkSq5rr4zEWYjlcJRofcULJ+zay
NpdpxG6laKuKo3TtTxeQmP83etOP8uSJpa43gCELkVXGCTbcFcwByHh9e5DS
gXS5/0JM2WMKw/Fy6xBVIrf8vvGU2ZqlqhlfprC4j40zXj0r4NCxsgeeg3go
f5j1o8y1XNmt5tgWJklUwHZCNB9OIP/C7YvV9PT474vAQp4vme3nb524NMUK
/xplaT5SumetDF5MaQnjC6zmZApqo0jmu8hAOQn0kyiFDzjMtDmZFkLdt7gb
vErNPMkb0aVUbs8kWqns/Cp3Ovg3t8Xx47mVYvU54x7FHZqbWrdJEOHe8GRb
uxgPLpV5uFfRA7B+R+yf1E8WGJigemNUhrpdNgkHJ6qtsoUpcMf20vaJIsGo
MA7ZFjLK3uE+LOt/+ndrIlyEWL+mgbfiwufdC3LZqUkvQGfej/ghbWeB6TMi
VVootdQ90W7ngZHz1L2gXYwqKHy2dJc0r/5ZajQW1eZajeq2XK121MFdfjJ6
FdpOPmsrLu+Siu0wR68VTzY=

`pragma protect end_protected
