// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nKntRqY8Q+Ox7vNaj6ZYalotTLv40uHIf2kJ1FB4oqV2Wjne1MbLQPzi29+c
0rQVSm9pa39UUv7fMiRdQRcmiE+YP/JozFuWG2qc28quGAERTwwq3FgYEeKY
5DryML0gn4Op4x9URmQGKRZMlTUaG6A/ex8QkpCxazAKhDAxBg327AEsuLih
5Qe/ZZnHFIC8c77vbk5XFFOrppfwN+L5dB8XeMsoilqgYwoI03SloHaq6mdL
1lAUToxz0eIaBLaYTpNQIe1Mt70bjyus8LMDkZhsJkfijxgCMWO45M5WMklk
Ify4RovHMFS404p5BohHTG5xZVAH6Uj8CHINKB0NPg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jCTkFpJ9KVJMP4CpVCXMTBkwsSkqgzjHHD0ltZ8ouIU8J9I1DKpK/Wu+QCbT
voRFKZvnGRVp4DUlI7zX+5jLup+oyJUYc33jNUE5jAgnxE+a8SsR66sA3IS3
K0W1iz1Ef1Ijmd7XtD7MDV17CZAuO9cCcdhC+y13H+G0Jlc+chXBaEzjwghL
ym1WVWs8Yl25kPNxuhYY/r7Vt+nti+zA1jyCxkPpQC9wkrT0vvDkHaHEhJo4
RIHTmhNkJsrkTI1wDBaz8DSk0VEMbY9oLeTTV092Necag0wH5hvIamYhsXhW
OByXiClI2JsPYGd1myO4jYvitdoT8XCVt+gwuKd03A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gaglNNiGj+HvHXvwzntxdGbR82D0D6NUmbn2fCyZcX7u+IBh/hqWUgTLP5tt
ToFTrzaT0zQEYFdJ4u4dPbi/QHDewazGHzDnAmieERqlQrXvempBuVQF0JR7
SdGkuo/4E8nD1BV7eQAp9s7sLeu5FZBVmb6Qo6leCsc9YR/tmA1Nw97s0tii
knI+Qs1f1zj+Hf6V9nmpFPUgdBshsGPOE2G7eX5NJY+18xP5Hk8AUoXgxVex
65teXDD9h4U11SFXl61a64S9A8b8k+2nEHaIUFK56eM+BC8otugk/lopTujn
M7AuYUp5jig3pRXw5oPKl5usJWfMVFssc+OWJ9arxA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pV/IvW2XGUuybFdrt1hYMZ39rU2qHwB6VM5t4AsR1c2j2cR1CPpwM4k4bV6V
dUIX1Bs6RhocOUWLa5C/pwNKRBeW1atD8U+NmMdmvxowIkjHwNXZfNkE+Es4
zCRX/eBgOzWkovTwTfxXUE2LWDZQDNfdeugFvAYrjMrUv/SWMJs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DjSLKZn9JhgRUIH5FWwBrAbkR6UlqYrCEhVZYqHBmj2udHmmsA1L5etWIU2W
eJaWeeT0Wjo6t0OgEvwn9nnlBSNjZ4J/k65MDyORIjblsh+E/F7OMbG05HLZ
jbJHZP1SPBk/gk95xQuu1W7qJlAyTZMxVoS7zvnVN+lTJZIDQJOTynE7w3Kq
ElBID1NSX4udOmhVjQKFf26BCDc8iNzk0kluQl63tK7m/XHP5il1lYSHQpvs
MM4tOKuOnebKCpwfgErkHrP2VMM5PAAztUUQWkWtrFY2oZ0q4zPq1SBFnyf2
PLXASg5ZT+dz7N8BvsvjSyjrKr+eYF0xoLDY7YvPfo20Py5tLw70M8tqtzAp
87TkW0XpubbfKmZDBqiThTRXKqv5TqtUVpAxbzK959W/lrW5CUZfxx1dyQar
+K8d3ai+rcxpK7RfKkcE90W1X90fPXgx4S6qLFbnpHKHPpNiXafkXKE3/qjU
r2Xivl/lH0vM7fI8SaveerIYG/8d9ixI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cplckjHBySm754AisG+B/zMaNPabpCq5o+ZYOLkwewstWPkj4uaTIHLpCFC1
0pB1QefzgyATxEsMtNocb5dCA2OptrOiuVcF8BeLtlXwYYfjwVNXr2Eq1hjN
taZQOVRswpJR4qrZHd6gQhwJQ8e8iPSl16x9NsXQWKmK9H5V52w=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P5z1arRG2zoFN9TI6ZTHsyIxOIOuywwkopV494Rrt467GxcaAwrfl6NMeRCs
RZfbwaBFVTaDIrFYQiezA7SFNflfrr002b4wI5re6AahiWLpOiSUbZu2jfQg
63s4IQvoi5uDEQF8VVFEI+R/oJ60mkOXcX7uxe1F2FKuJmvDBZg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49392)
`pragma protect data_block
+ANme/td1Az6oFPeBDEKqpWnuvW6KGojjBQCCy+8bsK3zcL8cPQ7usMJ5u+0
c9jj5pqzSc4xM1AHtkkI4h2RkksoM++aGa42oxMn0O3Iw9gKxm7wceicGMls
9PimbA4W3YoGpUiLYlBE5TGamIZDDKgsKGUoychjoS+0czvBwFdA6+2MlVFy
xl9f/MCEC5XPUZTGIq65HuLsmEcon2SAJQVNiF4dy7Uh21ej7VapQhXqEaHH
KBnIwWt4T3Upq1N7DRJNKkgYKzXbKZ1dW8QaPasULe/aXLOd7zoZzqIENpma
8SQkY1vCeW463HKnbAOQfR5YTiSWP0W10BTGc+fyxDoZtLa1BuYfGp9n4zCl
hNxnVFjCAqtVOcscdi3+eGs4mcKiakA8kqXLtYp5Y0swBL3cqjMCd9NyDEGn
QScdiqZKoPHiZQRoDRTJZHqBy2KQktSJdAtn7xsjUjRPFtphF31uyzxBb4YY
p7CG5gQTosfmJl2oTiKpPKiBTiLizYGijSoaVI7AaWOCQakUh9jPKQ90j0C9
rYI0kfXPTuMmokNgpeNHGbGqA5kr7b/h0OeKBvtOTFomRN+lP+p8uuamuevO
wmTjLP8DejA33xFyPSP+oX/OeqD1wgVfI4fzg92z/U2GqFNNDCAKrWkxaZw5
RTSfE7CNJujrJ5gqkmK3dZHLAmUWRmaKDkkuXneUY8qYOjIl2VjZWMYpimqn
GVvh79U3ulW2vXqw6NYdaT0PR1BasYUMxiT5+YjNBgZPR6COd+BvERAPgP/r
mFFL046Ro9qO/3yb77owSKNMzhCUVdPkSAwIHFNgjaFxLn662zd0uJNgQG5a
cIhtpbNhEfsU+V8o703vjFlnX0ETDUOJUXsQP2bBUcfWha8JPMVvBSch+L5I
Ly/moSpPjbGbcmNtxi6Gs6iuVavSioCQ5Qr/bKeMnjSmQS/91iFum/leZ+4M
DZNiOkfGBZcHOd/OfJAynRhaIpZydNOGxnKNGZphQN78U8OzZaOcHzEZ38nn
JgFmGVq7qcwnJPl7heIddDfJCdJLQD4RrGxnrM8Q+dp62CaIPIa663WQdQOk
Pl5y0p4eU5G1XdlijyMH0YiUxvhifALo5K9QEf1kujo5mTMfeC+g4GQDUiU8
IM34T1iPps63JJVjm3JBhOIlpUbiyYYYO1P4NxtBR2Bm90kE4qgeEfMHhlvW
ofMfFwPONVQNrnXRRI4POestL0jz2f5Q/LoU3RQpiGuHJl+/PyruTWKkX1gR
zVbarF9vAXD3pAQQ+K9n/a5zNUpHx1Z/eixlHo7wOJcFud3B53Yiqq3bpVmU
GHWn2RtOlIan9iWyLEiCvqMajqtzNzJ4YqgSvmkRsiRb2nXPnrm7vnXy/PiS
EDoRAdczjCy1xFdo1NkaYZjmPSkHbwq97rFQX1B+Tn5p3Rdch/0OCBuL5fuK
cUChZb68m24UsKbUlUA4Bpjmg6EQ8ZNRP/GpAVFxOBlwPxcTKjrfNUSLBnG/
yg8/cx277VbcrXEUCcuHMChU1yEQkMkT2b/AFYhRnxM9kLon9CroWRKtOsf/
rEfIAtbFuHl4xtHsDAMaCHOh6mXizMwvCDFW21srr5ldhLTa8UhqpjnFLElz
wIeFTQrClirIrp7O472HoRjryVngDxXmCUPbnGWo0idNlYsp2TJlAJ4XAZhM
Cja+vOWEU6DmbOAtXLUJfzAWapoTjq+C2QjX2GR7EkfMSouA7LY9O2zOgzHF
jXhIBJLPs1ha6NayxNP+WlOcdfY4FeULuF9ttuU5vTYxeBYzmZEkU9VkIKEI
3u0NlU1P3b5MpOLTP+8mXFhZvn+H/QCu++rM4DbRMhfLFEmv0//IMaqmNXks
dy+k8sbyrNE2VcT57QuoQq5G2MldDiaY/De6KKVaJwCyGimef695MRX8clcC
WsYZ29U+2inOF74q92Zb2qeJEqP04MBsmzvS01EyDGvzqxO97u4ZgDONR/WC
ws3FRlXB+gSF1uAO6XAKZjUANLLd31i8nKuBP5lVFvsLo01w2LLk0NP+JUvi
SyKnbHPeXc+XjMFg3ANiLdEiWxQyhgY2slG8FpzTHnlIw7Nxq2hqIgcW9Xfg
qnVyTao12+dwpitYAL0VuR3YETIS1w5dQOxXiGiGP348fqEev+9tgRpKZp0G
0X4qtTfdwakLF7lkZjeuzOSnncrdLdQUILbIhBqc6XB3tBXL/T0UZx3PNJEO
mYpRPi1Mrulv0CwUuLk0e/MG3uL0nqcEbQTYkfHXYAizmB4MoaV7cbENqQLM
aixcilATgrvnhnlDd50dyx40Gqd66AhXbf1+YYF6CxIin6oesCKmhJGpqjUk
nck4KmMk5WR9lMcOXl0A830Ljx8hLDPdABkRQYnSpOIUFsnosAKmayj6Q4jx
0pvblY4rhoMfz/H7bpzXt9HFh0c2MePR0YEcqwSguKPZeb4Z1ypG3gBHLN/j
KHeAgFYNwwNX4Bf0AKhXu1NXNBoT+Bt/OfWywMvU8KV9tElT8FNes0jizK/v
z1tAAe9kzIER2U5lPcfYWnA/8vxuHJ/U7HieQll778cQcV27iNLg+whSs/cz
Jt+aqfO1OQYmBSF11WHZ4klGz7x5AbKWuCXVSmQMqHlLLOYzNQ/2msvSZsyr
Fuw3OOSKDoQToohpKeT7ytTctmhSEwlQn2bcTbA1KQRw8DBi0n81whUTvFCw
k4E0tf22gv6NjeBcEWQr/qXhcLDVML4Od+rH238zntOcpUBr+5I9u8SuBv0z
P03kdKAJd8kJfJQ0c+/0GQFp0tfjrLkBo8UuhxvrOB2IHAp7Qb4C969s8/Ne
F2q8TeOxt1MyJAm7wJEIRrhP9BAwZi3mAdzm0tQjanknVFy8MlBZbb8D9TEi
o5gM+44qT1V15jrfW4hJqHI31U3f4CSOSevDBbR1EKNoRSqDlyHBcCqjdhwL
XDMjbLwLhl67+MPTOCFMacj+i3MhMCJD3cT/3Ihns+3vZ1VINXcldOMaT+m0
Nf1fwrQDdJkKMKT/M/U7uPi7BLXKyKGJJI9R2n30T8mSx3+wlmiZc9uo6KXD
eb92f9w/40Syi5/KHdxHc5R6pk1ydy6VccfJywKFe5I2O8o8+kp7bNb8KCH7
PwxlRdqq3487syThaOSO0Yrihmd4UG9szoqP/QJrEKShW0PDR7dndIPA/joj
Dec5QhCWku5rInybcA/k6Ag5DzjHs/PHaScpAxgvY0olCRQf+o9waRAFvq8q
tB/h2Sx8CrwHvRxFSEhEbGHfIWka2oNVG2R0FwG3+YeBsZVEG/zX9Og5SeIU
kKAd48JxegU0g+kypIyhPe3622IhHkiR8mk4vxFHdwmqKyv1RDc008ZkWaw1
Ct87dJeIn8s9TjSXMz65gNLmH3RsX7LtHgBkbbFwVX74J1IYv1j8b3WPwVmY
4dpMPIqmMpwOeITLCd0GWzJLIjXVzLZim9E4mwwiQ7hHv25hIPsrrLIwmjm2
xOv2mTzXxPVMGWh1/vGWEdpwt5R87LLelRW1CYvaZ4edl39xpr9JbJmWX2r1
Wk8r5T/GNbfegtr0l2URHxoX/VSvn122bCiyVqwPZfUO3gGgBHu0QGONpL8p
0eNbEEV9qxjJHvvZXGYxfouAKPgJ9x27lU/3+S+w18DWdoSRN+Urf9SrvI4+
SD9DpMHDexoPuMjRyf1++wCEUrn2DhVOztwrkrUzZUM+7Boq9ceyB8KdK/vB
9eNAXsfHYfe0hvXMnF1fRG1F5B59r1GcuDAseCgtIiB/VeG1yMwV1kTlM4GD
D0cWkbbfJQsSGDYJWniegZZP8YTz/5T+MtfEkQrnhIsR/EmDCV4m/866WVxc
zwaPV1ephmMHk72Xardn/Uu3hQN5UpsFutX+YDEhkSZ10WJz58kDkoIgWfrP
7E6cd/fbxzc5H+CCdWytwp65MY6dHXcBAAddpz3W+iLv4gnAjmbTOXhsYqFd
fC3J+UfAm2CkOigTBHzg+VPYOGogAs62pXx4YTYDBDN1Jfmd0tIgymNLi6qU
OCmmoHLhkCJwoebdJP4PlBimS+GZx01uvbInhrnUkVqjwOTa1YhR0Gr4hj1u
zp2P358vgGsIISHg49e7Y2gbeMuA+9PyINlndKhi4I8o3lgveZCGFxQRfn0p
ExMtEfXLhe1Q5MoYp+nWqu3rewexuBeENW5qjOMmZT7+j3CfESkrVLWzb+af
Qhrf3sTI1YOmI164YWyY8Mr087tzvOS000axbBWQ951xUR1C0X5krl2GDL+7
4mUo0rD7IrZOgbXDp4t5+cNcrf6/3PGlP2Qlal7aom094vl/RNZp6p8dG71C
N3i334eQA2L+TpkwYz2O6U1ao1nbq5UUYsSeCI45k6Y2r5EbcWQren2JlIrV
vTGL4F2cUKAp/wWb2NnbNc3GJKkqj6anT6xbwtNHF+zJwEfSTVu6IEuOisqj
EaAGJSi/k5eS3J9qv1+Q8IGf8pntQMxxObBBNUJ9mfOgDeE/Uqtf5DJof4BG
e8Mc8I6kiYVN2qWVIOywsfLXRyNHzevy1b0ooPE6+agivBX8aB14hwX3u2rm
y7ojFnD6/OGGLDTwA+KloRuVQFy0QWbd0aKJzoPIfF0vRbPKqvVSgF3KKsBG
jZJIHmiKMo7VA5OHEPhiAskxipU7UfWc5QVaREeeRGik17yaMdlm/6bl+I3P
rtt5aLOyZDgB0okOaFffxKRHJTv7B1f3zH7DEZEIEsJ1/4OsPG7cOCKHFihd
9ZIYALGOHdxMio/+SwpoxHJoZ3KhNQh87AGKt69ttj4gJ6eLTQOcL4YhE6CR
rSAyX4q8FvfftuzLUYAg7rk8LwiSDZLmGE0TrfMeQfwVRdawdDG62oD7ZA3p
BfIOuS0qQeYw8ETKoSuJJMHMDeCouygf6UF4hyZ+iW6dbMMa9OX+h7EIBtLc
XYSg1Oq6bsUfSUwTtXrxRYveE6L8OJiQu0VTL6CrtM3LvNoTGwFyB6H3tbaA
w72zRt1b291f84mLiyHfrYSk/AM+H7Cra4dxjf+8oIILJLH4wBKZhEQrre3r
jkLniifwNgup1hxsqkVKBMBWSlBJUtOJGRjC3QqGCMmZteQqe9zl+gw5T8aN
tk2zVqvXNIiPk+Eb6mccprL6Jf2Z/teSolG71X5pCcVCINoGLIFpJ/oED5ko
LKws4m+xEVnSin1xg2PQTr338ujcWadKtBfO/5PW3MMJLjwX/TNot7cG7gub
Mc4i4q88Icmc8kTO6fccZDuy70117lKtqVxnbuwhG+3b6jYS7yD+7ieUsa7s
IV9Y+yGAie/8XInUrJR0v2KdIoVYiF4y15xwUJJOvxRDBlyJq1qsNJxFzaOs
iSKN/b9WvkzFZVJb1/QxkDxkC/xV3VOllL80s9yYmEORIpfdOHCKFtpnPgs2
UWXirDkVDsnGfS/ScHeMfVndQad0aEx6LjfUr9n+aMHuEiYbCmjcFXCFLZ5e
z7aUrIYLPILOik7MxPcyltH8txLrI+jexIvJSx5CwmXPeD2/zV3a7QSLlrcS
J1vbA7aFh9q/XLokDNE0sOtDW4a00+l1zTttFpD25+lmod/MUx7GwjMBWuJj
K3yoy6jVSnLdWJo7QhFEAlsG1r25HUJ2t9KWOXTnx0o9fApwzAjN+eX0SZ/d
0gSOJt5lPgl5ExZgZEHiS0sqEWGrf/QJFzyL014GilV2igj1ipfxXngc6olt
aI08iN9+JRZYMqepcRuuLLENffJcu0uy7cOWsEljOa7IdrTr8DI7HuQad89v
e3XK/eh1gUaWtToiIQ9wO5+hkJx2AY+4yoqhRpwRh7LUFA5GCbOB5MNN+/i8
jWl8WG7jNC8tCU5lvYnSpvNZrtUi11+Et6j6BfH66IezircpGtq1Co/nSLUy
T9QfNcjhMAJXexnV84pgm/LNiZfByAOVerD5DpfJrLLS/kKYehVHcIuM4xd3
C5Qv/QbkQ3VVd6qbiIjcIQddt/tzHQQV3/fiVC0O9QVFEZPHJeqltUIzILA6
V4lxv4SqvYrQGvfqe/X1aBOQW9YAYEafcCoIV6ynFzMB/txRuZc8tvBz9Pqb
mW7o9Mt9IfWUsi6rFLKzgFCVA6/MZO2RnBNiSim684XunEEuyKlSG1rFMHkW
aqKFC/2Sdm3Zwj5jWOQeBQza51bjYohrbc34Ro3eeZMfU3V6BkKAyVxM3OKR
D+Eagc5bWJBZxi2xG8ndASVHkQbfYkd4OOpymYAPoblipqRb5DjvGJXyrj6j
rx8Hw08G6ltYGIv7ntRbPfJ1VRrBLnuhgA/3D8/y/ez9fld+QKfZvINWVRjm
iYNxgrUbh+M3didZkD+MSVtQBZiZR3KdayDJ0Pzr1UlrMP2hBGzuTN9kWNU5
MAuMJI8knu3CtuOTeVmoN54RWW4TRpE8SvF71x9bocrp7kszVe8D7p09FiXU
rxK64z9RkY9ZZEckThlUx30egBimcLqa4c9aBopU2IK3c88lsDsdugdFG2hW
8ydjyDl16Kb7FBabwwb61qbW86pB6x5uWx4E+KDZ2FVeLMPPWZIRw/DUe9wl
xSDAbbb5c5gHde4XPoqKnN47Iz0QhYSZh6eYf0Dkv1XUsgu0fvuxEha6w8db
Sxs3u6nR/g9pyHRCHuzwq5rFcroy4Byk+0srb4mrvHaZ0gA52xGHqoNAUz78
BDj+qWXG6mZgPDmZv6tPvk93c2fv6l4/5nHuXTVa2z7eoDRbg6aDql/Baic5
p/bKbFx4A0hchQPBGJkgnxaFhNtQKkhAbZ/sbB9fgvlig2N/lJ5eH/AkDac/
t6P3n60FafYL1+yiJHPwqQYyTVOOFljYPT+7sT7IRCYjtDcY9j3DfcWl2NKk
HmX9OhmuBgUIAiRYbieE4pWxghid/nhk3g8MTN4pq+MdBKOqYW/oyd47CABu
OI5ZFRqv2/LZ6y5fRrUxzTN0BJAhTCH3/DMm7xA+Z6XK4dhnERe2aSJ1orjN
xWkscauceDRM43/70wKQ+OwH21SuDZlRHYK9uxnLUToSPIKinVKLbe3CQVno
ApW/piQrCCmuSgyqsUeOUbQv2+iAwopi3RdVdd2CkpWBufErGLUX75e/1NHV
luxt8AGxdK9qb1MAwDN7NkU7ElyiuBZoO9oiIzAzIIAXYbBYl6L8BCQ6gTE1
rx5jZs0cmLu3RgUDNqhktBiq/6HG94P1QckTlNC+y00hHGJD7akXcgAHAm7B
hQp6C17ZSMmGcBFUFQT0nTomFz/qc3H/V1Kkzlhj4RFN79DnU/7ymwnLRLbF
I6pQM5k2zIAuZi/Jd3I8GaTSIsKmDweAPCxzoruoiWs9mXzjkPU9inv3/lKx
GMW8PA04VRRQJKtXUf86esJRGjwCyY//giDAQkEjVC0SJ5CzG+DZ8l+/uTGc
XnBZ7horoRzpQNcMUlbRnPo5FwVJrkoZAsrBWhVxHP1kbAlQYKwh9wX+hGVh
4jTRgyiceo2DPikYvTAirye6CQFJo9UU/DhUsJIRcYi1Zbcu740N78UbIS2g
ek28VCfjWR3vbhGuWTzHzWVWH4vntuspSyZhPg852Qi8fnfksTsgC4sRxo3A
8ykvCYBhpJzQF7BYewmv31xXxVhQklCXwa4fPjE1Q226x0WLfYW61/i+OcWe
LTpwMgWn8ylULBxowkjzTrkdwaO/gZTsSO3y5e1+NI7/oC3sBfhJH54YXKLj
xpgSXVSg+quIpzL4DsZ4m4HClZhN3/CE5XPrT7vEAJnlBB62jrDaANG9DZc+
EVRGAK0Uoka3qY5DEas68U8c8nfZoMQ38lzvhKQbuD893x7Ip2CEvNcX+MND
a66e2Nf5T+fK6gsIaNZTWRN/yCzj3NMqMV3sMTFDJuPBhdUOIGuuiw+0j79S
R35FJXni2FTb+Lun6YH7wTB/HL8xDJ3adEcieZ1wUafs59EE+UZchRbd/8pt
wK/nz1StYJ9cDfnv9+BjLkDPs3/0qDkJaMIAQ+5UzpBNE+t/gGMRNFm1Cdur
vk5JzbzhWtAuORcmBxWf54y8O01dIG/jqRB2JoLeMWLUf+Hc8QLaWBopwiYL
03jy4VwOi63/lH2DP2yN1Ef/oZzlvBtjJ3x0H+i+FHG3n4mKQyVtAbDoe3Tv
vBxKa5RIzx07yFWMJTJQJqB1igB8Dj5xDoZD3ZGZukQoH2LrTAIxJ8+Bq/19
xFM9bbtDvCB7C7whJZ3EaaIHDr+G1H+dN34ItKp69ozVxL4JAwC43eFpXlWH
21X9dP7SBwcj/LdwVMDViDxvGj4gLfZFOjxQKYtCe3YLYW3Ijt/Fw3eDCl17
hWNjyIC/fyu7S5Ur7hi2UNKBsRCeSb/yr3PI4dMBlcdH9dTWQzwROHjKMAqH
/9EZo3lFutjGQXt8BKE02yO/OTIbWSYTF61PGUqw6NO5hvDJvVRLYdMthXvn
+0W1h7EtTwN0aTGoV5tKEnrvoyZzpkPyCHnIrz4Ls8loUH13pI41K1+tiEpU
cHta4B5jz4X4CHwLNaombAvKygDH5Czaqnrl1wr63xSVnH0e+Skwbulr+uUz
UsorsFbJp2Q/AEUUgUr19nT+5HfdiV8aENYYHqvPfIah80Dnp1sDrQ7DnMw4
aPMSNdB2ryGPLaVQfnIKmLl2R+g7AmPQ2vMdy6hQcZy2TtsULp/c/wOTzaFF
QFgfOxiSCnBXGAmMnFvZCUsNG3qCk0V3kPePWI2I2M+CVijGIw7NJFXqM7jj
JVM3LbuaFcNy5k0Z8EG8ng8ob5iYHOt+BNmlm+BeePYYMaGxQkY1DPNb+7NQ
E1qzBGqa+Xxw+1m3KlqYWQNjY3xFuQuo2iYOVinfoJP0EFeAOeYDuSxLXJ69
nv+LMT/myDGBwfBPlF+q5pQ+ZISTtorS4iuQghn2BmylCvTY+Gm9HfSUMeEk
MZe5S791/e13VJr65qzudyA6UKWWdhkwp0V/7ojkafDKkM+4qQEDfP2rw2wk
ub5vXoE4S491F9hTTVwDIEzVGbhtTejyBs8FpdHHBUkHtmZ4in5f4Nw6ZBnZ
UBc9ny3NUateTmL0TE670DI0m9sLoqKy0cOwx+EtLIaBBUCxUt6OPeRvhZrJ
mbdGzg9uanpdTzGEKJCuXX9JOD7qrzW5HsaYmdPLt0SD37FVMv67QTaA+8Hn
t1nUQrDkBo/zDcQwF5qvcgzHtwMK8rUz6bwdJsi+VNZZQXIS/Kipqm+fubKP
5WOT6AxoSTrLieDmCz/l1xvDapNvvJo1jjrIxuVoCpxhrYJgYtvtPWje+/jp
PEzX2pNQG53v4mWzfj1Fjhm6Tp7fiBMGoeorWm167toOJESuUlB1aTWpPxp5
b2HuhuN6TD6ZqaywMkEENsf7qhuTzfdu9JlguMynK1MF9Pe+usUAU2NfvSNu
jhmqpYCr/dNbi4gHorggnX2CuJBDxzsFngR40wv5XpfwHUAZfBLFyJv58K77
zQ4OmHs4BBJXIVZMvWnX+Jnuc+7EB/bcYqZGbv+liso4jVpnSduuslpAgSNP
at1Tahj8arE6dHBzOgpZXVucu0MSFHxHiK0qMWt1D9PisgE1dHfjxjD6EIAL
yG2HdIXyLNehH569Mf8in9oq8YqJTN85lsxePsEsuzLCZyzYbr3Dh7vPEiIB
KkAlNer6ozIkhyR67iAuBqn4r/CFVnqPjHT83JjqHuD7Y98cZBmSriWG77zG
siCTKGGCliZNetMlIH5ybsVcIh0zke+C/TzTU3CltvEYhk7qBAl/TU6yD3Cc
CFVJyAooo7TK8WoWNYuFQhnBWd7CUjKv+wzcPbVM4t7ub0R2I3fm+6hnJ2vS
06QlBxxjgZRtG+XpMnyU2mT658Nd8aSOQ6j1vLznsuKALiaWVy8fCFtbMPRy
LKh/hFluDXijzs9zWCBPUtYp2wg2RD4QBpyF2pq+C28gKCl4L5UjyC5Kxoz9
uZ3KOmameu0T4aI4KbERyQ8VuxebfMk9sTzd3/zYi/npUu8lt7ZM7+79dxau
hpGPuRcL6wHRLsAA1vSJdMkyDC8UC68A3TEH8IkBohERZ1q0wm4uF9zUIJi1
tuQXdJsbRrsgS1Gi0CE1wPg+y/fkQyoT5DNvah9PWo5QsNUFU+bI5EBWuKKf
mLzzY8npHe7PiWlybVZneDCbxnoyQr/dnZu2mzd8WUsmmqsInJWJHliGItE3
ivvelTGVIZFpUworSzeieZYmssOL7MzxBcHb9QDFFcNjtvCBTfYmi5Eudx1g
szWWojRrtTo90Fa+ZIsM+j9VZEYjFZNh264TOFPZj+X9iab7a3HrZvs7/+2m
Ml3WW+qnMTR4TYI6lNBdY5hoCs27poTde9/HFlRBjp4niF1GPi6S0Uesf2tW
w2wIELcv2KWK94iPYbouUaE4FOMvVVW6hyg/ZfBcmvh7/KNFZ8HpKQndb3/R
aeYknux8DJGbI5RhpVgTsqm9prQh4o9wsm/UWHfEtuU6INTgFq38QRu1izxj
xRhrmz4ACbW+K4FF25q3/DnYqdBB1h6hqmM3Gx8VXEFruHvmuKFNGIs81seU
BG+BFxe6v0W103/lL5PTeH04SRYZz+pIDKfPTDz80dI4hEi66KpMhq24Mi7T
kXTAhXAqHJntSfbQkmxQZpQco8GNF8+myhhzhFan263uSx0uhc5u64yDmTpf
pf088JnR5hjzkYtv8OGFIoy0a5mx3dw+xe+PC8DiLQKP1QK/u3n+ayE0ZAIC
yLUjesYkm8Mef64h4pWRskbN62GWKNObx/T2qtXLZoRoI5kTXOLOLcCE4OA0
yG7HwDKgd3aC0dsN6diEYR+GwSaaN6J4E/565a3pW7i1P8oaZC8q8UI81uS+
zIImvOA9YpIjCNmexdoQAETjeprkLgjM+sEKdi2qKSiUFbWL5A+rT2RjKpbi
aAGkSKu+eqARnmn7kPNY5u8KZ5nzHMMivwR0UpCQvSgpPh8VLc00fjLT0Ml4
DGCLTy6XBJwR8QhVmUVeyaHFuCsRaW/avQI8GKvFbTJndTSQRqF/2GfiRuzS
dwkj/GBKGko7Nwbnz+tNfW2IcaEwlHYWEvUjx7z07y2utqyCzX9t1n4Svbsi
sAT5JqvfP8sMHJKPGliyu22ynZLpQHDJOP2+QVSyxcZq8BS5qVEgSGi0BLU7
/9/mfZm0/kGJayhB6NuhLj7eVauUH3P/qHv6CY+DxDpDr6NdCB2k7EHGpY9O
RES/Mn2daRIznOE6Qocd4Pi/yICSMIeQg7n2gZfsYQzgcTmIQyO6CPkbT44C
RuoEo3f/tDyC/1AiT2aw/YLaApnW19J8LrWmkwG7d3Qzo9HXuu7l3vo+RVk3
zZOFFmiXyeaRpSL4XlKsQFvs227qS3nYDkc78eD65hUY6Y3yqnNwLYCU9evn
D0co4SOCNBWuA4qzDH8CjeFWMjWzXL0ZGKmb25pTLAR7iRHQt4JRrQb1Jen8
keaxIckfrzCnCMqks+8r5pAtWE7gSUiMeYJxe/ra1vv8YbChTJmNRnbM9PgF
iVs9extLp4BrBcl7ie9iDEbqZe03iP//LXOrdfqU6Hb4u6BWJqiMDugFl2MN
3YrJCSxt6z9jz4JDkQlg+wVpW4HNnHMw3+Ee/r5hDgQHa4KW7KB1mWuotRDm
N9g1seTMX+IAgb4YhoV+XgjODbpx1R734wZM8dE8oAHEQCyGuCyifXX5rMu/
aKgauql3IQqxFAOViFIqyLjiP0ZWs9T8jqYEX51gVcdIwKHsijZpUAkwEXv+
6hvxhXsN0rb8nX9m2BHLhB2whKQhUFVCr/YRmR6t9gcgD4pPP31pt0PwrXJY
zMrSzttW/Qfxbay1hVSQD6A+3EuAVE9FYqTqRbgyfRPEK9X4H8fOic7sDRyP
RLFIR16OuMTT8+x+krr7OowHbe8bp6nWp4Af2vUS9hpJUP+X4kc1rVLc1WtM
SyRizqKhe1+6b2lhm+BTuyJvWhd5+QU3yJ21oUrWBOriZNW0uiISP9lHcEwC
27J7sYe9VdBBatyomvCF0k6pU9pIlH6/lvB/qxWJt302FnsjF+QX0EvJC78v
SlLYbOp5QJtKGQf91FBno/3zNkSo0X7TH0DQA1P2MX8We+wl/z9EAmHlU+aF
FYn8krLIspjbfF7+TgRo6MRjQe3BG66osBxcZbcDYtd670V75bzdD8lmKY4C
myR8RMmEVtNIF2OMEaklwcwdySKMU4jS5fxIPGk7NHX3GcR53sNvfXf2Ggic
ydMeZOdEdp2dhuKcK8TgXqwaO2l8fsUNXBVeZEEzeaOB8FgOIDfBVwV9brKc
tTwYztXM/Epr8aF1VcFydi83aC0FJs0AiwNUEWDNrvIBKnQcWuKuonVE6Agk
avpBvf4MFH+bdTDYeZV2PHk/aQZqx7UtGOaADT2YLhhBlgJCXm6hNSQEA85O
MwcYX7rz9+NQgsYPc6fRnxsY3GAd5OdMg+7kiRJZNH8vOcshJlEY/8mEg9Sk
mHU7LVje5XZVB3TtGKgP0nES3daH7IIkKy5Fa9fiiTcbh+9O4gALCqVp7tqQ
oCPQ7LV96z0qXvM7VqCdSTCd25QXuoITIEftywGSbC3g2vZHpE/EjMhfxLeu
sY21XMnS8h6qB2N3knKDWXn3vaKB5l/3fvDIlPZhq32koKMJujuPSy2yMwZq
3TdYaIRxXEw/nadx+AqxRUDNmBVLMN0OppWFmhQj4gg/B3ysXT7qJs7rmhTO
5GcrBeV0WILXaKgU5VSzkcZSpiIWU9+WdJjhleEORDIQ5WmMIBvnhq5IA2QC
ZbDCtLGgEqGeXP1dt2Qc1b7ZpFP6N7W8b3bP7RzcIqDBJ6diOFqs046qDQIm
CfFEkVzdLjm4azjMnfIpsYZCx3jXoENsLP4KAufW3Ds050WYGWixduji4yMA
Wx+1wn3TsVvsO1CUm8b3m73n0CjY6cPGtz8M5kKuvEkWKhcGtCmb8Z771VBx
Os35jGVuI+p9DiwyJjIszFcjkVke5RPCBKrTvyNKJN9qpO1tJYjptSRdx1wG
mWbs+iXRGVQrwlRarI1qQSkbHjmyO6ZToykdf9FUFmZ3osIgLopejWy7OYNu
KWtG2DxdVnTpFRASpLsa9JlVFN9+jVzAPpVxm2qddsS8TCBoeVFBgGHXV3SE
SXA7QEhcvLvMfK+eGoqSDfb2yulxx4G1A83XwxrCpTb3cSOC1mtXLe12HU/y
IlzJGfo3dMb69DK/v7zsWSWBNcVsuwkhSiEiU3apG65uxNlWgb76V+BBvsS8
HuOXKbIlS+JzjsbCq1fpLnsSmnmzJnJ+UM7RFi25WPMvVsXxL9TcEmZ+UJNQ
Qr7rtIiEFh7G4d9bS0LeMWFeudPX23vgJBfqPSqiwTe+2T/wPIYHJ2g+gRnX
CpTVnp1N28lOpixUeL7A3CATbrRqunD4gjMPrJOEAPcJR6JR6lEeMS9nCL4n
P39ietgPr1mSPwICy85av5kT1Bd8sz3tExKrDIn5y+C+DS5oC0sG+ckdwUVF
cuc3HXK7TYrdsbmXCz1b3PjkT2wwYd4suaJ287CyBiONLd9k6h2+7mGaWY8k
LbSSvbCST91NGnQB7+sQZbYfzd2F9KTzjrhR1cpr0AU2yNQEgLp0bGwe/eCD
cLDCKQSerP8xgMVegst1AVGGQaB3PAq333Cl45QNlKnrd93vKb1HP4aJL461
8z6Lwns6j5n5xhhtZXIiExoDYId18NnarvxzzJQPY+nHEzJyt/HFhPfzgBlA
NdO8S+BDNW+4AUlPWwZvJt0bwN0CPKZ2wyNQxmD6brEUzZshKTgMJD4iKWu5
aIdE7yRfMaD7D2zNpHNXpiD9wSxV7Yf9JnlYPBLF6SkztCut/CTa1WQtCtY8
4gd3pu9wEv51WnzIZAtIXCQTSBrcIKJjNRqb3RhhBTe3VGUp5tWSEzuqhiDz
EGJAusSIuk8RJq+Q54WXUUFVfjo77TUKgyClchG84/YlNJU7WlAQEuN72Het
qKHNgOH9MfOpbdntYObvkfdqRQhzxOl5q4IyfUhttJh5eTbTO+b8yC2oVJ4H
GNuLFD/XbUsgw8GqBeArgZr4nxVp0gSRhaWM9IssoeU7EwJaCk7xpfDgWgIf
keFy0+EL8u+ZNerD3nxREQ+kAsu+bVo2FH+YFoLnOMD+UY+jc36uVlwCN1xy
NGcvHy+6Z9Vn8zPa2vRKN/Wcd06P0xRQerKIOBek3cMgwZHrJ3kNnvAD4Y0P
Oq2PHUKWxw5I7ztPTQB7geMcO2bY2ZBYjBYK6ED9mVqZxwRmbBvgVZZDcMXF
UD3LNrizpS/xhqwiflvCSIIjUh8zSCZHA+91mOI67us43q4dDrlg5+D0NB6O
uhqnwDXEdcd6lGYYp27jmTVouX4F6B+o7qG2OpdYoILZtiOyMCGi19jrU9dH
3pG8A/zVqIE19SoXuGpWY02U5k9oAk7ituCRr9PMZSnyeFB18mj5lITNaSfq
zevaiPNt8/dDElfm5Q6BhswAf4BHMsDEmy8ewH4Btg5oOxu0ELVcAtJvSL1/
p3lXJTzRjNP4FxN+CyyLEDljHuJhhA40fMT78t5PuPnlSDCHwpgBQOBtRAlY
BowWGzHIPNOYs37Mj2fql64rLkHKGRVxNiE7bZaIDOb69oRsEE9ybQS3d/Bz
mbgtScJRXfvSSZAkjX0TCUZXuTCWFK3EFqDNK3t4BOIHureMgb4Vx8/2Hpyd
VLnVc23l2LThhqr2L6KZs2A25MpZ5Of5sLoFhPFua52esQJ5UzwyFSlfvopL
mlq/fC6KW7FeNTWl1Qm5n3yXsFn3WMEHLlHvJpK2BvvVgMrW/VIQTqXj17sX
vbTLpTvaN2alaQG5kIkeOKZ1kfnt34IiL1z878zuxUzw3/04TL1qBJ/feXCu
yZdTpm91BFQy+4m3A8ijZXuwHSTSftH4OzEFzOVBwmVAiAn0jkknYok/3h0m
DxR+8VWi7CsAFyo6f3u4wMGjQ6NUN1wK3TA60Wsdm9OvnEjcKk2+jQRAHEJn
Hmca/MWQEh4Xz5JgDmIebT4noccvxbcTuc5CfJs2qiDP9dvoQxj0fIm9r6M5
ja5IWKKcW0TX/XlttbNpIQXP660VBhvQGm/Pif+2g7DCaIzQM1UEc9cD8HoH
O9nBM4CHqJLve+05eQep0Rl2WMDbe631jOZ2VRYFAdiTkqvGfNxpexquoiKa
INos9a/lAiZXLtVY7fyGgKw0gRBMNfmJluOSovuSvL2483U1CpafocIPSKUh
5bYI2ImTga3ha3BGblfvFL7/Ul72gE5kjVEzbMDRVqT41JxrKCQD1DiWjyPo
HaQ7HKsKJAMyfNC9dfZkV09i3vQX1HqkbtiM9MCgZhqf8KbQ5QQty0KVcNjp
158+frcnFj7lanwxsyRPcRVpc5i0vN6lGfk751UaD4+MauYMG/ZipIxoIDg8
rTcB3Eg4xYfuLEfCkPFqSNW4m/CD22FELBCH2uhzii3WvZT5D3OMD1lbzBTc
L778XKVU7GS7Q8WqhffL4HpExnPOefZNPRldHrQtrHA7F2CyquI4IM4qC7xR
pVkBNsv5FoDAjfFu46G0E9DNfWOWpH9kXoI9/k5eFimHWJ+65mAxXXifc070
TWeSZZwqpVVoQZfS8y/1fxBMMoGf0WU5G0acXddo3IQuf2leLcIDN+g6XdMH
j0YYHbsfSUfnpU6bGDrdWATYHP6/Q+3ca0x/PKPm5v5WTub+zw1e27VL6HHw
0hrHgjou8115mnfj+oQ7WTfa0jaOhaUBXSRk9L0Gpu737ZVTdzpkvC9FFICX
uU4TKfMB9kRVahlsZaa2dbMjkY73pJQoZbKDhrMdYoChK8IRUlcqaJ99hj58
vus+1wGM7rdulDB7b6TQyvLIllC+kdfqmWWVDcmHNiK+82Sp9gnTHo1t246U
Tuw+35sM7jSOdYkv3i+s+fAaq4J/WZOT0ERgyvBA6jwliThMkWlMVLPFPdSr
sfLNZfjmg8GjEvhYLwqSOqqhwmknvGr25VRvSQOKG5BDN1iclkTjO7N5b9LD
WmAD5oTSUq8W/2yqLSuzK1nv9qbMC3vS/tcUvlMJ5AtEmurGZBtHU5wqxiGw
jyhiPJURNtJQUGNKn+PiFzzcO4V2Qan3e3IunjP8VFAZDnlxeRBome4iwxUv
0IhfhEVY/3x30nvtDKQZoxmciyDikkqrU/F9bgmIdCZHpmcHAOCAFs4nIPaU
TTq0yU/SOpWALgrOlEOpSLxrl2sctF3iZdy5Q41UC5+ltDOVV6LRYY9BfjDI
1c5XLDU2GI3SZ6bBNA0XZQ+0qqUk3ZECVoGBai2kJN6L7JkeBVvdf/8Lghkq
Scb9HlklSQKhq93zPfBx/6q6B62aa6/mgIWmMjhnx4xsR+jXIqFrkPfd6aOm
kxxEaY6adqMkIOt0+hcr4ghPBO4bOuea53RjKuK/DSisDLkMAky8O5lhRHHL
+mYqRZpBQUPSvloTCmI2Il727PAOI0z+fVUB67CPcoR7IDpDyVP+yckkpW4d
PHfup5Oxibf7TBRuvQNglQEMmG4kRO5AOoJYYeAwd+HMSnk8IqjfGskaY/aH
YGB6L7SC+8PpBgFCI4443NY/BYc7PTZnv3ddoVTygwYJpsU4py3btrggyP1N
oE86kSkFEqio5SiY7sRyEoA4y8UMnvEe6EDp2lb/4xQaZSRVLZpDaromw/51
qFqvS2VTNzA+xeAjncRByO0L228x9xNl7ZR28uXsQPF56ECXNPauF9xO7tex
mh/76A1xV8VWDqhJcNmkDj/Pb3u3lm5NCDoTryeAoJ8EiIJ0M4FW8zBzU65R
aLU13ehldUZcnhXMc/kB+7cSS7i4qJNsm8aRcv4/qzkZiLeypJpqrnAe57p+
YNOdrH27/KGFaKx9L7d4pymVUca18kBQXYW4J/ojifXDpQ06E6hnrewf9dB6
EGvxbEipca9WNZL4n87yK9ULxTdbrFX9cu/EzbMB3eWg2wi7BvknhMpQeatO
HkWE018076K9tOhLIVwztkpOcTgqbX9nzr/7DBQEV5psAc6EaFc2kKHUACyb
Ncgy1y+YMZUj4vpnGrJCS1VPpG8OrftWsdfXnnzRif60v396UgKlQ97Nr99d
0VFVKaobrpzGXn/zxJvJXtl1TKx2CaRAlhXaCZL8RplpTAqayfGEf9JhzGRv
PegumYC4i4GNUzJuIDEDGRIQ6cu2QxUUfZYuGg12f2lWxU9x/cQNecieudZW
N6bTfO05E8tStnZIuBi9z8nvSPwy7LKqirb5U/oi08hskUflSculFyTBsBSq
s91PU+O5mIR9hK8UQrryecr3Tvl8QOon0nxrk6d3SE00YeiNm5RfwBRAKQq3
V/yUypCEOaTwr5FQYbfdO9GxOH+sClu0W0IwjbHaQ+48w3DmP3JuBQZ/2WER
w/1Mcw+dcRd5RodyUHiwVfyk64T8n4SXdKsAmaMcVe+85een/SXhbUFoGUMc
hY2JpjsfLv0i1MleE1B2ivVK5E/fkiYlfq7Ei8yNs/YdWzpqRpZGOoNJRBgm
S+P/feBC6EDOVJrBSWwsYTKrdnBwQKpDlHQtu7mdA5L7m3r1+f041aKNwaKR
pOElgkadcYKkrTpg3a6fG08LXldiEvWCTvvWSOzNw2Xf1qlosuQgc5xrg7HG
MAGLpAyTVEThZATE7a0KlWi5LaV1Xt1oL5O15KTZr5NDkTN38IcmeAYuyYM1
+v0UnMB9nX5NXe7N7rlWbg71LfNrlDBLJRG0dKNYymuXuGqFCUsEgCWVa0tX
ijQTukonKbp5ijS9PpQPa9Fs/ky0SeOIUiRvLUS32egRN+MbhE5cT5mer0TP
c1UgnbkyIZa83vbODiXaMn6Mem6lKuyMwZSxgZHvckfiYI95Bn7g4Z/Mbbss
rz6zUQ4ie44dg8KXZNlxkz4JavWOnNFJTw9xmzhyLuNXPIcSSEz5WFBngBXO
MyhPTPVTdwN4KN6L5bwfA6ItqPJ/T2rjXattLXCOyfyOUsi8Pd2AWWlcyrqC
i+73ntuvuVYRImuZ6FQVMEXL0l4druEfMCVMN0GDwOe81wV7LdMFSDkEjU3V
Ydy+tPYanzPeOoYr3MSuRivkMdJFUce3nrNXehf9E9X2MXotLc+b+8UxpaZs
FzUcM4IRkNil3mwSCIfQTjROoxDMKDzzFdNNCCEFyk9NPsoYbbiRqKU6xsrU
yHflhBRY/VtkRkkAoMciowJY+M/y+ITVEjlhi6Ff6qHzc6j4hT5+LisGfAIq
rvWm0s6d+rJIb+XYysDyfc5pH3KBDtiPXJgMbrzHtJZfD05JsVZYthNUagGw
okLrJaBdU02rNk/JrbYmb145ywvvTTFoUzfVNbycoEHZ/1pa9iMEWODJpT55
WPXEKyR11x9RokR3hkPYjVHEvd8/1rl/UBd96dP16oABxkENPlMKPzKBJ55c
j3/KNNw4trqAeqmGlTVCaW8I4a949K5wGK6h54wSQHtQ71lHB8/oAJaTBn7u
8PuJUJ3RjzeQM1bWEgErbstQNqQkkFUDSmFx89aul6Fu+hulF9B3vLI8tf2X
KMKK19/n8Vzp+s4V5RRanmE6YefT6mPiNJb6jV+Bd6ThJEY4DHegjlG8J78F
7f+zaMZAtLINJg/JV7HVli/sRHVr4WJVWAL44kBjYmo6rLiXTiYMATMTgCRJ
jmak4fJUl5RSxzg5/AgsgvMeLs4ORr9kBueZfR/00evT8wsAq7y0p4Ar3T5N
sZX/jUeaHJLE//himo/h8VdivGh2iCLt8AeILeuv9SgHYY+os83x1wQBVSRK
wVB+CH6ZQokprLOiRXsCDQC0we8qlY3IuDzHUZ0upJw40MKv8QsLRxSCWVpT
Tbz3rjtsxfqeJRXnpgMlDbF+Szy5XNar+bQkykVe9ypSxDXi6s0erfTZqzNC
gLHsl42GVymepwdUfEWFZi9mQ74RzijXAf/fyyquLZKTHz3dYuG0EZGyy/dn
kFwrn1FEiJ4awgspm0nRUJ9D5nW1LpwqY7fzzJJExqPSbjmXudBf4ZVA5yG8
2LCt3n4fsCxWmt2TrUlbmBkr7tSVnSZPSAEMGyWv8HOPDw+gnvQY7Dppt6L0
XbaZYMr+qZNhbioufwAjK6zvbK+N5vuiYo5TsXo6pkskBbhN00PCQCr5EZYo
8Sw5hGsQ1smAuDlIeaaEZg3FfgoGfBLrKjKhorajPl98s6bW0A5bqYwXp4CW
IVVSj4jXV3m60Mk4WzgVhs1ZG/PFsXRxskjoY5fJCmt2PO3vxJuARCfub9eo
e41OPXdffummudxXoEhm7NhutkpHUkZ0v+LLUaqKuUsSKdM8+8rhNhbkU4Zd
5YrBDERjnwdNxRxjeNLfJX4i5iMdgJnG5uCk85NFD9qDZ/0vXS3WjNgru2S3
wqQ+FYyFd7Xsx0iKIY5aUMiYf68WTz+nrgwJ56AEwM1in3cWVnYeccBqrM51
zSfc/1qT5NnFfAp79Yf7LSI2a3U7YbcUqpuvzYhnQ99B8lEOf4ThK4dzZ4EM
eCFFIEdmO1v8s4phHZn+OzyR1rVU7C2QW5GbA4NOVTgVk4Dx2S8DrQohYXO3
KgIz/HRK5yd9AVeo3uUocUiAvw+sm+uoTIrvHUcJcAzmT0bqHzrb61ZH3g0f
IltL5jwnjog9C1OQwi1nWMmStk5yPCo296YfaOoCqDrtGPzExQoUoBff+m0w
Hyx48XhTtG7IvaasdQ04bDEl8X+vbF01nWsdy/UeHB/LRoqqMtkWgdFIE2xB
15lrhmMYDfey1lbRDWapkhudsNZTRbMmGH3eRfD921fXsvZ+SqEtU/3TVN4c
NCiG520KJPuLrd9WW0bam0/rXfR/o46QU/Rb7nWvRYY/IKtaTIx6FwpMtayF
a3qyzgJnwsiQuPmPYM8NRHAQxXjUlnzM02jOnxR9wgU2RRgJpC259eL2Xsds
AkMc2337ZGNYRtA3Y7BpANEC2Vwa8/XVRIP+VR+BLZe3bmEtkNSSsQZf6zPl
kdMKZb5OFKvLI6LQ3yPBDKFlF3Bv1B+NFhdaRDHMtSFm8AoZJOvas6DJRP79
fDVxw4gUnd7J+NQX1IIdABItGSLbV/0f3igVh94QgEF/tfbg2Cfai3sd4RKX
GryBarugTEKAjnbCt+mDcQlYiGAjTCm713IbQt7DJRkMiHp1Fj+3wdjZW/66
+de2SANHAflCz/RW/GeUXQV4l8Pr+A1iwCB+WSr/3FZlhln9cTTRg//8Gf8Y
nqcsZH5ZmkOSGQ5BmREWPo1eoq+b78u+uX6WfteZLlJ8F8+80IexMTD3nM2g
eXqnhjp597jbPkw1+WS3KScKQHD0CM764z7REoC1juFvPOV2dknKLkoFWjmV
t0tHE/y+V8/u/63B4xH2PijJaUkjX+iWLYT1a/J3Fjg+YsUxIbDog/yVfaGm
K0OobZ5Fkvjbm//7gvVI/Mlm2r3PkhPZ1nD4cuTMvO+F+0L9L4L+vo8hZ8Ic
zoVh664VsRGghgGi1z+7ZAY5D57mybsnSIxWuWO8NTkYlyA7qKGGw5us1a9K
r+yrZo7Hp0W26p3beNtiWzdumh02NHvtSVdAXgSvr6/ca0O62CJinYcw0muX
QJ2EZ25meTH8pc8UFygdZlbiE1pcS6vFffNsOtU8eGYjqMas07hhhRDN7JgO
qeZqhVWJEeleNMzcspgnehsRf0sXqBipE+ngwMQxTJlkF1xFeAFV6tRjzZsA
B+iT9+tWlfR7BRSDrDmTpTPRUWJQCptac186CxENqiz0PQmb0ZXQT0SBP7TH
B5h8yHErGfZZtb0wJ3a+gue82AgEhQ3yB+JTFVUAOzQyFXn01j6le6hfRjb7
vA0ipUuy8tdxiqjtijHpsPgzc1zn7U55K9SPkjMp6WbMrfbHjtax/QqAc0y9
B7hU86n+u+gHqGm+dUdsRzeHOHJ2pKyF4eiUHi4aOHlQVNjDD7HtkJA8JYuh
QeEHFfqdnwq4C+/UZEvpBKmlYHS2EOt6tOVdo6HJ9udnL9yOAffH8xtYjBcw
eNMpubKCV9q9+ZiUQyBI9uktEtJa7lm88M/4hULoRI5QybmrXmjkZlQAkdnq
umAWAAV5iAYwkTMitD2+qZ8OcqaKWu2M7rCV1VRbFPUioPnXIBVbOqZFdK5a
RlkYXte3CodxnLrI+spDYwo0hC5ffGZJD7Lo2Is3PJ1JDHg4WKYsrbZCytJs
U3V1euJAzT/RmBuN1FBeqt8EaBj/DiIuFI/jjcsaRIQ6cCDw2HcYZq9mHlH9
1d/3UrL7Uiw1oGucJERFJ+iN9UdWUe7P1YOPtGa17uwx/QfqH72+hmJTlKFi
60x3N1yXiQmqVUnxVUcC6Fqc+Sft/2iYRfTSyDv++CamlnUleFrNOKc5Qwhg
Q/sygUzlgtdCLoNuBkmX8pLf2lz14trAVDgbTQ7p1tfHMhXDJX023Q/RGOZ5
PY7vr+nbUPgSM3ODezrP0vIwcXe7CDpIzh47oGEftIG/ZLovsRCivfVp+tqp
Xj5GiC5jtDLyY4uuNTiwNC/K10DGeGO+RE3iCmJaQgtMzZ44bGgQWPLEmwgi
o9VH5jiVwF/6YIgHizgvJcvvlJepsoewDfwGJxSd9+BVQcoxv6wtcPZIIBhR
ZFHgSGYHYJmvOMbGp5WfjZllryjbrDh414gVBkz+LsXFqhpiE2em3bL11KkZ
oEP3iOmgvlIII/T+NkhYIkCHDLkASE8btrTcLRViqlkbKH9Z24cf/eN7z62V
2foJ7LbysV8KIfYbDSQa/ejhfciZOM/jQ46PXwg2mIAEeum3ROMzslQnoJTz
6EmFui3KhqtyT5mC2Q5zA7TAR3kHANLwvwdy5JAg0H0XZQiT1NK6hP+qFkeE
DPHmUWNcqtPz2vQO9hXip5BH5aD4Im37IkFgj4VXgYPTRK1fa7xcuEbMe6Mg
yG6C1AEKEM1CcVmxLj6mhOroAS0fiMYzJ8uzUyIwr9eDI4IiahqMPzAGarm7
0QI0n/P+td2di95znd3UZqLzK6GvNjUf3nIW13J23Ms5nvJUu4guQ/rWg1na
5H4qZ1HpSGOhEAGj8qgLGSrJqKz6cNXazPw4oy6mmfpe52SSapuoB+kOCeKS
9NUrSQFn+kleqAHfnPvSJHySENTwbPOk1/gjWzEFZ5Cxzm3pR0ieU6uQu05a
eSvyFKblpUTrMbwvCItBFDBa345zx7aEMKTSE+jjv04pghNcck2ZSLUQQR3/
+yhhPC0gfcV59sywO0y9dsVUBUuu4Jy7rjZcomqpcpTl68QuyS+U75haQcHt
YaouIu4gDQfqEEHsnl7nzdgvwrxgjaTqrYEAHZC8sxHr9QKkGeCqoaqLEMbk
NqsZXM+okRdwNUh0OVkVZxJWhPkvcAXgt2Qh1aGGpVhExS65UE/tLBPkLzim
80rAmyDYnE67Krff6lMloxpnpSdTvSSA7C6rRSh9Bq1OgVF974KXSA7uqJ4i
AM2wl8RLpI9Avm0aD6mLGgla/2dnHeLL59i+ihIdS2hyaW/z57vrYalbvboM
IHLr3wAvOsAasZCi1x0mAdbA8AIkhrlqhRT3VAp52zyZqkXigq3IJGez1OQc
lYAvrq4SwLvUoPowsv00oqbsy7y9yf0O/sNFZnkOdz3lzTB2HtmtcT5XrqEj
8ZosSbRZ/jZBbgAJcEsikv9slZ6eJV/+ykbsnPYhLQ5KhjXju99iBlJ2Hmxy
B72siPkeOMvAsOor8UfefI3dyVgTJB0RZtboZdeSV1MgTWhotqTRGVI5WkBq
lZpoh8mWlAcC9ecQnNamucnxvU7N37j+KmAwiJH7m0ExsG/o3CaG+L6ckZz2
gvmoUVI4MAi2OzdoIQNFARXXDWFvTwU4e9jAOqbTkAXu/pWcupIwH/JPp3Jn
Jw05SfcJ6Jpt2/nHZpG3Kw/MB3OKKnWsJUGX+F+zABAsJrxquIl7iO2W1VwU
TDas0DiPOhmDGqsCaRPjGJG93IDL30rcblNYVoVYpKtSlCct62E8ek1xdf7J
0vVcwUrCw6A/s8uXt1vBuDc6lvMKSCjttmCJu2dzlMEuL0KOmw3s3yNrwDpQ
4dlvd9iJ95ZzCOSLk3RXKezy0BaVjpVjzsca1iz2Owg4OTGffeLGbDpEejUk
0aqr2k8udS7ma5mpiMpqErAschWu9qYFKWB6v/k0Sor/wx32qivG5u0RENTt
wacXC7JXepAu3+6gnQQjBOjmEO2N9sdMJxa7BQhgjEjKSYL/Xhjme6w/c1Ff
0NX/crrUYffi7rtItRbakq1XtRWAijWnBolo5EcSkdRXJXLBKqwm6D2eXTTP
6510LfAN9GdVYw+V8zopYGELdahm6LiZkGJKJFXf2lSt4RZCUs1hZq86gmja
CzFyNADUMrS4zc7/Yz59nKMvoVGW1XrJqQJNINxRt7DicKxBozd6kYPhdhdP
GlhntPl9pEE2NibCPeFJDhfLz/fsHAXjhYYD7NVm1we/5RnV60vY8TIncCx9
5RS9Dvac4F7gEDxUOPdM7NNBnqqTfSkYPiqCzoi3rBC+Ui9bQDNwxbZ47+h2
1lejDI0KY2tkqLbI6CYLcvdqHUTunjhm2J7gK2rRyCwEzISjJvpdAulPlABW
0HVsmjiGTfnZgBe7dE9mB6OkNOwXHWnQpTpsX23titjOZDh+Yi2l3Ms9ul1c
PRZ3fpQV3CylpIrvf377C/COhkTK7GDVKnsNN/sjVVkqfDfu54NK9pw3U9hL
FUOIRlgrsPq44tSEmh9kZCWyyAT9dZZSocYDgumJG9m8hHRZwGOT94+DRVIR
JNf+8NE2SpaE2VM1tXJ3y+r3gqL04Kd6XWZ2wFoQg9cX+5I3khi70KgWfrtd
/OvhZ5INypvesvSMDY2kTx8+m3SGGqRcyocsG5RMoEs3bSVuEbAsgVSCOlwI
0CKAl2FRpNdKgcWpW9pnTU3N8P2drIqHfkVnqNO+Do5YNDUelNl/5KjO+iMj
rE/dFHJ0fgUbjB+w0lZs0FRFO73DWFEelH4WQlkklomTG8ZSf94QTfUVcZZa
kclwovZPOlKzHRI6fC8ZDceYbKT8N8wzBNjpWH4xhzV+H8D5Z2iaijd5x0iD
+NKlc9jyUXqOgs055PgbLzJaGlcW2DIAxH/jXwzevEQ1uL3HUQ3kIvNZMyZs
Yqlm7qFp2OpmtPaCyZYsHkSmUnJoyT5FDVF2LCJgspTf06PWiSAPtx2uhE/z
KUN8iBV9HhmHftNu93mGUE8kSA/VVTJs7HgfUt6AR02O0FxV8KwgbqnNAdqv
xn85xVOU9c/bITJ21h/7vViA7LSQCjOYbvqiQwIpb2X//0Tuk5UyeZCFt5Ff
Hrw5OeT04XNgbxHzdXJBnFddfWTP7y1SFlud7udEkETzPv+6e5a0ajiJnHWn
yc4kJepBbHOwcN12khhp9ZctL6pn/nP7WJt+FzMQOrpGHDb4gjy4WSexLVjg
anNw6eE1thkrJgLG3M701PmOBbGKCPwQ+qbTd5RikaflAdUa8cqzrzlkd2TM
UNXRZO1JnwLg3JudPwDvFzhMPKHTpobUzDuQs7o2rcFXMcSmSF0orZ1wNZLn
N6d+eqjapCP5oajA/hr5dv3Xz6XWcMHKoW/LWlQ7XACNICcC2Q0AEQm0c9N9
rBQl6gDtBWJ3YhnhrD/0ne3OszcX0nfV3EqS2Fxi3BiZeA5kxH2n+ULf0d5m
HMZUA6iZHLjJ8qlcfCxzop41OY4lwKZAv2EcEMDqHDC9kS9GPj8WgDVV8JkU
AAJLLAZqTPwDE2Gyl/+G+/e9URN3gECu9oMvGr7Xliq4wrg3y6nFsKEKNrs7
OPlBKVeldVRfWP+KtGwykhOuon4mgGv6lRKHdp6ld/dNS8maTl5docQn0cGy
P1tZZkKzl+VGjHQjB85cbn4ajbaV8aDnXZZKOs5i+d0kT+nIhiMdYNJ99K0g
uPwqRMqLDV0id+RtfygXiZ3CZQONj2vdbsEiAdNsvKd+SYk/p1ns6JTxOlFP
9GtqkPheCRmVwoZ4iiF3cc7RI/GKz6+2CH7KYdtprWyqofof4hGTFxwFqv+s
Wi4jHminULN6mzLxLQRlKDeJUnLvmWhh893uXQrwPN8tGKa4hcdzkNPjWeye
0rzmWDzBez2Ea6eVY6ZKs/qovVRm5Rch63W3nBrWOF5t455bywjyWfl57hXJ
1b8tZdXe1k1kx9SOqDlADOLFk4FwuFh4lEl9WYPf3usRM2WInLSBKIRrLZG4
RmfbBaF4slk8LPQ8qSM/rWzOeEZRb61QkzsrdMyHDxJV0EwjZBffE5erwBIv
XKEd0vrWgrSlvVqLRQSf0lAVjW9mVc34fbIbVkxHn9qqxQ8uj4K6AINufwGh
QJmPqeK3bV7L0NmZhkWRJnaOBW6ddKOcCUncPHnhOQWULKKpDIPXYUKgy3EO
ywbtL2CbZes3izzO8AHZU27P+L9K9tPr4C26FwhId0ZW+8IzIX6vk5Cfgeey
l/wcJGsXVvMjY9niJL9kJoMMPShZVFSVU6sfKD7QAgOlGaV0xVhrHAgrxP14
0yeq2D2lyrQa3+hxtEtoovSQbF3cvjcY4p8/0gPJAylMjjiD/yp7NRgYEni2
QV2+gC9qQOrXh4PqqhyjXmL4jE7rv2XLTy1AHwqfqVjh/cI44jG7Kx0/1EUi
hPQBfyeYsqFe5BdcN1IvnolGJ2COMnUY7c9oQwmE4wI8Gvi2gwPMcpeJR4V2
Tb+wHk9myxbnP80Ko7pwA7379mCqw+WQtcrdQOe/Ms/WQ7Uw1vtX5X5xT1Mm
QV50mds3rfOQSJ2tZ6YsIQWSSXSUsKlzBtLZg7+/vJtDKWFvcYSn1Jo8AZL6
PIIgigMkKorQC765QtUgy8mS81RRJerMqzx5Qjzix4lVCdy3wNTyUY4mNUSu
5v8coYdOH2xLKafN+hBPIz4NPxhWzotaBqmmZW0HAFtJMoNwz00v4ioElQbr
11cH9bPZGOsimzBfs98wXT7W0uxLf6NVQLtScS7XJQbZwR1Tmtk//oANGvC1
q7ypZOYm0h7yXnuoYMcWRZfyLRDOrk8zTVAtCaUUrR+D0ldEaoxv+62jn4Dn
IVXvGde07y5iiIl9oOlRWw1zhbbEwwoUm2XAzHnqYaCOc0flwNQcj9DvJjSQ
AmlMRE7RJLbdEVLL02Qt03p44uywUnZTCphCVC/xgvV1o3lBnj08nV4qDagx
L/YMdedZ1iASzVd/EZK48+CCxwHpa8LnvArOxXw5jVjBfX6kenpRS2Mi0JYE
QpUhzVchBKTKaizN++FzPFZw9uHFJnmcTSs2gr5NW+LqNFKaMHLx6UiGJZDG
P+/iHqA6Ao2N2YsUCmJEg2woOITpbyGwgOVCS+Q9T+K2oIjxgeLhWGiBdHjR
rvEH8jz2q0WolTEdw/orkRnn2atbVRlfwAso6ca+xzX8nbRRLkCmNOwKTuYb
HI9GbaXIGo/HTaqpO5qIHZkrtpu2u9WglbOBiyBZ2x5/eikJSluG7ikTCJgq
9WTA755c6P+732/u1RoOCO6/iJCdufX1rcqxYSuXsV7gCcKkdaxyntg1u8sP
uKQWaHsp9CqGEJXd/a67sAHFR+SI7GN3qkTiWDIv2ql1mgAJg5Mo5ZQYx6EF
TP49Es46euNIK01bzl68P7NiIoPl70qgo5uaYkaNb1Ajsea87efPHuWMsUIN
kfCFWb4yzjEbtYGnCUUaEPKaDh/9ReZCdnJMKs5RXK8Nd0s2BFBC0E3JJkn9
BL/bMc7VzjAQi4XXY4Oferi9hRrzKbs7oFIfH2x2uq0LT9zxOy1ybmyeMM/i
EJ3JWDnQP6r8wXtjyR213Sn/i7p5fdKvNFTaWuBfrjSU77mH+8NkHP9eZjyc
CJVb9CPNeQ2gZjIFQRVjDseL5TJfT+9Yml/R2LjguQIAzKS5ReLq8YEBZYY6
wuXkAkSCcFZnUbyYSqzxo7YgkuoKzZO5zoOtC7cR3qYkencXz1oUZ3p/OJWw
fYDDZOM5BvxN4NlbnDSFebnnmVJe0X1q0j28rDDk2xhoO0CTYVEEHxynDbZJ
b/Cm9lE2kcqoMAFSeiYVr33O3JShGd2TTMGYNSwFKtWznCk11CR+RPhWCzpY
qA9DTSIZMjDgWE7qpVnwb5WUNDRV4as70WwUbk/3Ddwz4CPPXqnv++1BWgya
k1G2yh5ZivYe6cS4Ez2pbwVHvViAGpbSr/r+IJj3g3RWWM2MypQ9aEMwam3L
EOapOfNUxPssjZSy54vGjel8zs799ViAiJ4qqVu8ntNXIbWMhnLIj/xSgQ5c
pukWTPglVWTAPWj1a7Xxze79x1UnWJCScZ3Pla/MsSjiImekRQu2CPQ+7j7c
MvaMvOeM8UffUR0Xp1nQUL6ibrmIoHxD/Zpjio3/hxtQsHePo/FQyaLk+DnT
jikF+AceMCdDVeDUrzgd3+9ulnhGQIg0aI7UOLORX5jy1zhetJJvwbuLVhag
mltgigM/tqrPBQXWMT7e6LcQF7AmUs5O4kuaR1PIs7lOKAV7DI8+1dNdlcxa
93DvrWHxsomUduf29FcEaFxKuTVkyCWWo4coYaS8mLl0WiOyk1sg0G4hrmpn
2PtnP6dak1lSiwC2Q12SOW5hIqY5kBsFT9CTuQ3yg9E9c/NVSyscYWSOekMq
CzEmmgrLihKOWBrOnPo2+G+hX/MNx8q4LXlVV6LBG2wOH0Ug0OLEsMWKwuTz
pxLXtDtZJ4nnIJaO3ox1/n0LnVyZu1o5mKAT4JFpEcLuGM+icyYLxqq9tLoL
fG63FghsGxZvfopQ+UyUFooejmry6WEE5/iMEY44RmTLXh5Sb+vPsdEP49K4
dX6xK2esKRFN97onWQzDHm0rJfFUUbzylNDEaDKBdhmbdkm277Isvw4roJ1M
7HzgQeOPU15SCGKANerJewgZkqXHI+rTNdp1s/KQrLjsPNqxnAMrdYTTZJ4Q
EDOG4YwFdOynLLma4Z2AoChpc0+wzw5SP4nmtXoiJhn3akJt9wWp8ecM7e+7
vt2gAuwfH/t+KHwJmRDWuzAW+jxHMwRaEvd5R3X4FzwySfRpYmNy8F786P4Z
2mwQvc0TcWaZT8goeLD0cRQLRYYng4DwzTqIGaBJgaKanyzSDByD0fHD9o7c
gwoJXJs2bSbJ075YSNZpjhc+UzSBFMkw4pI1lnXeS35ZS1ie85AF57t2LJfs
3zBC7uRRwObT3Asm92JeenXaS6nnTDA/wjBMuomerdMRCzVAARemkZJJvdoD
0pYzVX9J6317HsnVMhQ8ilYKvOxWWxMHYfOV+0sV+D4xT6F1VuEdfTHECzyX
M23k0WLlWjWBQqeyTjnjLAOK+5INOH5qA6AWShSSBVKlpdOBwYaFF5nMeOOH
Pb7TUyAM/EIEODExOIof1u4+1n8KSAhWZe13XvxPg39Qbnfr850KkxlGSLMr
fnzxOV33VzPpMNNt0dI2ZrwevevSSo0DmBWdKUm4poM6whYFtTQgXLIr6cOc
n66hafOA/w+Sovh/ST19L5iMJm9d7YXNgWAyAOyv84u5OEYpuFHfv6yFgjxq
k6YHrnesOT+gmAJOgzcWhZ1+hCe2VLyRVPdStZ8fJNCL855zuL6qDE3Z8mo2
m1zbtNdpFX96W8bT0bcKaVaUibOlr1FP3leAOQB+cbPdOJKHoogvm7vmDzUq
6kG83uMi1muirB0X3qDHYdqyXDa4MmAW1Dgva3VQrm7NB6hPRdl8AoVvk5uo
rW89KKllOjV7AjLhW45h9oQfKZiQCC9XCsVwgs4kmJ7qxma7g7dZtmy1RyO4
MCMJ52IBvm1/1zdIwU9PqOFX9sv3pXL9UGGY98fvcH2EL3sBNOWsN0itl6qF
wN1eZIHd62K/j4J///eiVxnEMwoZFoFmIUQ2Vqhh61kXmNk3ZagornqNvZTC
2GcKedmuaph+55m76zkGn8r/zNKpDAnkUqH5LJYTfoABQFBkf/TWtQRZyyj/
WcshIfjhl+ip2cKNsHTHfWm7evQjxzbVb+M4/daIMDZl+d6V4nxf0RQmdSpn
ICFmfaB6qbSVj6jDNOUeLAodQ4CJcYK5O5EkKSnMLZlbhRU8fpQcpzGTU1Y0
wuNLNvVCqA2lHgertPJLQJ0W8GRq75YyZM3ZibhLsrB4C5qgatvs8b8nxvOL
8w8Mjc64IT8UAE/P5Yel/KKY90aiveLKqQdZDXxBBvn38Ihr0gbVdAgwQH0b
/1kzw4adMWhOqIlUv58QLtKvz1J7Fydkw9YygllhA3v5NTPNfkBEVz2/S13u
qW8mVzvBRxQpqGXLMIn3Xlry44aP/NAo51bB8c7q/cboIpMBNiNDDE2YhtQ9
EW7WjYt3BaVto6l4L67Dt8nZlCGrokuEkZlie1d1eg75+rnWotGhz6773kql
MGB4HlaZ2+5d/BJxCQg0EJOHq+jJuxraeRjiQZDWgO60iP2q+0s8K12ORUYw
Qvw50H7shcIcwQwgBwuzcqQLKPaSncc9KWFKOHmSs72h86z4IZRviXLWFm6G
CAj9yTs9tXJ9Cdwid2KOonvEIIqmZRja/qp6UG0VsniKw5782xLFRWpEwX0Y
W5FMshCnVzjnbF3odZBC+EkCXwoSko8wp07tpsJxxHRmWI/exXZYyOGA4vJg
0UHusZ0NPrbnFTCjMxQkcXQJh+HAQQwdThuv6qXjiIDdebZqGiAQNhLnn0Ok
xvp+OHeuo2rX3td/Vnvd90Kl8NdqQgPUOw+8xm3eyPWnHBou7t/nDW3Y2Hnu
OZK2uzmjq3708TZmqi4edlo5wCQFxl6ZPQg+IvJFAsbVnIZeSDRtOC9wgiZ1
QJyCnfy5X0PwQvL8brieS62c77Y3ujU6SW0VfmAdMIEbQHo+Aykt8AaPFpaO
+XwoV4ISfFF84DwDfkQ8OymSXxKAcMcaU2Zg1Wzz0683LLJ8opgIKsBC63Nw
eCR0JDd56hVyhsU2MrX8M2a1+Ey4cgbEb8m9Geufh/Kz+ZFcZu08J7zBjE3v
yiubJPIMwBG/UogFnUfsJE/tn6XYG/38WZcz93VrcjHYLPZLBFnT+hLIACvG
NzxLnehYeSZ1qcUBSmsuO94RvzC+C7nLcEqlYvsHQQBsUXv8S/Kug1S24gpL
bNVau+a/BLdncKhCH2WzCDRb6RtoKrBNtm0hJx5poeZf6YF94OaRHIAB6u1G
DGx5s35UCCsCdkubhhF1OuIBaaaxja4clp+OUO74vJIlzkvY6rd4BkU05OZd
UkwPzuFqHrna/0Uf/8ZMvCS+g5/EPr9mRrCmR6bK0rn9Dnn2BPE0cUaZzVlh
KUe7BbAfIDvO3xSkYU8HMA6ipELf5Y3wB/HN6fzahDy8x+0gzqMbwKhLMwVv
S5w46ekj9CAuKVvz/6n9x5trUIBzN/HEILA0UY2fFXQOyvEChVFCAXzBI8r7
zL3MTIpMK/CFRY6A+PvQja3b7BsfP6CAskgBXSTrCPwhFPfy4oNeoK0Ltlgq
pL+J/n5Xeq+65lUAi7nkvTN5VgNEfscH4b0SNl0R/8yi3ic5BjZm6311d+jW
FfsDt6QfNnUVc62/S4FlrB1TIKcX+yL07g0/VSxc82+gzKjs6xIxrNs9HxLK
kpyRChIJ5Q4I8WzvdWkBNzKL6I8iR3aYreBdcswUN/jC6ueBy44k1CZwszWq
SVMYrxTpUyAv94eGnbl2LgGy/0juEaaVEZq+tu0KgmWKDrDVMVkaHyNag4Pq
iOJJSz1RRFQ2XlOLhx/FPfvA7J2EMiECPKIJiT0MV9Xu4n+al5n+rpey5Vz+
U/EQ4wu1N5QcQUl/+PPHWVRbb3trYEJoGv3gWVOuBooJLMRJNqOQ3nXqKWFC
kGhvpn6Brla9Thyp5jafSAthf6I8qmEA/oEUcJQkKBqDGJ3wjFEDxJuP3b/c
fIgANEVf/zihsNb1+eSplts2vcoa4AKBNQETM1jAJ3J7OntLldFcrpG1nF5+
krAMJokVf0iqM7uIsFkPbo6YcHqb6fWmCKXgSXJpnjEu7wjNZsaziw31a6uT
TbdRbDpPTdANlMpoj28HBm/qk65/olRS/r8JDS0YRHESn+lyiClYwj5oseMS
ZJwRj10ZeUanvtfj/yD/le7idgRrYDd8ItjEheOrYYT4trMt2sE2aCuXx30b
zqU6zXHkWGKc2vXJXJVGRAfXFJvhbXI2BmrccT8tEAyg32Yog/KW9+owctYx
E2blWeOgoN8TX/Ha3elnInJQk/7VBFGwFB5K8B7Kc4xSV6CKRwITW2FtKDeH
hBBwlroHP29kiOX73n5xj0c0nNFHhs7jsJQ1odEChw2QbcuEjkiyH7xyK9k0
Cmi4koaOmZVdcXkJHG8qsniFAh2uQRTwhWEhFaiWRKYr5BIFPY7Js/HsWGZP
TjfcylAd6atGGxd1EGf36+fZWJyxoeCo5GRad+UqbrV+GTJ62XwbT7cCYwvC
21wdoSsPJMBBqSgvs7K68ptZEFKbxeH6+w26KXVS0hEwaDjV2S9z7m/qiZQn
uijUC2QG4iUFRKriWE7TizbvZPCa3WISw0qhVsH8mdrC5Sk1RYOl+Usv5Odm
W58nyapGVzwMgm6M1pAIxMuwkJBSKywOK6qjVTdUfkKNrBprerX9bbpz4aIt
LTgG6HQ0vaEfPAUanTgpGv4GpyGCk4W9SsjQVo+ktTuGsUsDPEamWMdvtaB1
n/MXSsUO69T/9Rbrqu81rqEcqFuhvfL+PS2EC6/A2hl7TQ3L4iFAkvZ/8rUo
TCdAbfL17pFO+OkUUBonGaFDR/rSpLOXlTYMwaFYD93txlONEbRWiwOQz9mg
M0ZqEmOkICFquG/wlYXPYw7Ix06YWs/OuU34/oaEd6F/sQ4xNitiM57GNsXX
3NKxT1EjNZNYgsxYJUnvKeenm4n7ItsGYDyAB/a9gOWnanwBss/lCKM3jbt3
6n8VFrol/V0Fiw+rFUiv51YNTNayK9zmIe5o29jvYGiUErZh+2z5zHyIqoVR
v16rw+XkoOZumWll/+wFEBVA9BX1FL0NIL8VwCKWOSIyAXjL/+xk5CkYsxyj
0vS8VMMQJPqyiPcNROX6/hvSzxmGR0PrW3LFxI/oYrosqF1csVfS6uRwop2v
Dwl+eFPW1eDQh9FJpTFWlSm8xB5X0jlMrO/wDbh6WcUf6LRzDz8jW8FlyGdi
Hu9sLJqqgyUTlpKqMKBqvZ5BE34QM93ROqsZDivefIMOhqyYKlKz/4nKZ35K
GsimVdbXDYDovYbT9xhofmxauuCujm4zHpkpOHI7OEXI4fp2u30qiMSfV8Oj
q2L6riSGP3fqGLAUD6p1vD5TP/QDew9IWzpy2VfOXEr8qqXFsPUvGEfRsGVB
ElKn1RiFwwdhEODrI2e3BA87+rCAPITFXXJQKU1HfxvOAZTq0fHpqNhNiYoq
2nUAG/JzDFzAeax83ZecyIqPQeay4ms1zTv5B77lThwedgjPKpX4IQwkoKMQ
xTiLiEbu36IN1+uNLspUGaWirI4VtdHf0DlRatOVRROvggtixO9/9zHMD3s+
z/ufn9gaBSkg4oircz1mxOau6iq1U5R/Eg40WRlAw2xgaI35vNI3ZgkigIfg
CHLaifufcVefK1/Nc6uQDfdHw7fLzP0Kxm416LNwxrkUsNY+xi9nnPZmfgCE
Hl67h7zRcmwvaRvJsF1xKFvUs8lXfdW2UuKSzkt2AHmJh1YiPz/Qy5euSDE/
KjrI4XUTwBBXGXujGUWsVXg4+rYpB51URcQJYdRbL2mbRXxzqpti5c9miFRp
xEsHoUu514BQUmfcZO9KPPfpqN/85QJGysOocEIpbCB2B746cT+cy7QBZRoI
iNF5beFSbqtHPQ7mqGZVf85+lGoTpMyXG1+FqGXIQ1UTCAGwGldKclnHpWv5
16digfRS8POZosbg4iHrAYsk4QwI4LB9Na69k7hfxO5jIuSUj1B6s2fwUWVy
HlRT5fYM8FDezWgB0Kl2YeGEnnMHkPMx8j0aW8Iw+8r8UQDXLrb45+CnJSgN
qmdQ4bL4DLgfs+R+7BLVSf5qz8j/NJfdR+jyx3VlAa05Rkp/hX06ZGTbLcCi
5gu59khbPjRh6roj+B+5NxntqghdsonmOHooB8mNTdcNxrUEaLzprglC/j4F
bCOYDhg6n3G4eh5wYKn7mxWa6YKw8C1qahWCuJkVywxIgPd3SsZ8wWTbFhaT
6YYaOVudoVyVapSvf5i1zQZAOP6PtvsDsPp6c+7eKg3SoSI5C3qEqVHchb8L
Pi+AuOU/s7emcr3OJpLvJ13okSWOwa9JbcKrNSm2XDvh9jSMsKc4/+OVYXQD
/vhMFPYSTiQ7BpqZIL3TanZwichQNakUB6I96DvXJ7CdlFmQ8eX9KC5NmD6d
W9lFl0xa/1CFjz5TaFdef23oerduYYR9X+3BCu7D9+4gSPDIMqHp40d2/0Xk
xQ0DkDQU2iZf4GVphWaEukgo0wFmA2FrghpRS5lPWZFZU5D6nJd3XKheEB8o
3yOTAx41a82Pu+IHrq6tUu8yfGSmODwDHdVgZxbHdBr3Mo2Hz2x875243Kql
XoM8chRXQ71f2ZpJM/pW23rFWkB3kf7GEADPOVKlZCVJZdQwZ6wwX/m50RA9
G0rAw1ItDk0r+PocV7thHNwb7mUCQYF01+/JFL813GPXL+X2MvRhmVHrjCXI
X497toWRpiBIhDV92j1t3ZPDOUHh1g8gQo+3V6eh6W8t5+kXm/uuvtbdu5Yf
cxBEj4Omk6TxH3dItC+whhw0DPaTU2nlkeaZyuGg7ydThMnRTILF0ZaP1e2v
DCgo4sJpZeP1Um5CjTQ/Rzevlk7XuX3O0MeZ907av8vjfUwfKqXvWgsF05aC
46tfb7ktH04PKs6Zxh5mme0qMD3CFusGPCptCptZl8zx8N17DM2U33TZA8fz
1Pf/wvPispFCF0izzo8IgIoQxYyzR8caHMCovAUyfR+wDux5/Fzan1aHy8bQ
cjMtktYRhnWErLGQ+vi39AmZK5YE0xcgTVStgsi09pFFUkHx9PzTfgmDEyYS
2WYOa77AfjkxL/7MZNYxMMLvfR1D8tTnHisJU5EQbhUP6A1E0REIoq3aZ9Rl
vK366G64lhTDasNgS1H1yR3VXGVufHbTNHg4Gd0eSQX3vAUkPDxuvI9hiyul
vgLaRI60ci6t76c+ep4lwmoQPtN1p8QQBQfz390DckZfqKfVBHH1XtjvkmIj
tODLHesPWdjbqtOAgpkqd+qjzwOu44oHB7nQJJYlEj114miblMwlwOJ9+MLA
DCw1BKSGeGbvorUrx1+JGRf3vZu8e1FYBjIJCvg0LNuG0f7fXSnwbPgr5WRG
LyBT4OHA46Y3hfLWGBztjbv0WQ438zeINrNAsdyVOs/Z0dsJF/NtWMdV4em0
KjM/G6nj3yRbHfdB/1Sgt0AQNSFd7h9vaqDdvkkCNeyXicmnHjsikXdcvKjs
4kqjqL7WaB/IsvA97MODwEpuJcnGjik1dB+7vdrCpE/alkX0VGg5F9BjbNv0
xZBvHtVBCNhWjZwaMzRznnb/esdQ2ePpifIek1rJi3AhiellmrtJCXD2Jdws
SGTU0otmCQjG5uwLN61Ho/9Y5flfGpzvpKUQLSTeZ6qORbbLUfnjl5FTcTAy
zpFxxg3fDpIlQ8EHPv+0ZXesks84NGqUwiWEo8cd3S3Xi2lXcdV5A+ITvWIZ
2qiDTS0YZGhu3qTpTjnGmFVj1H0IDhuuuJG9/GXTSlCZOnymTXpxDXbXm0Mu
dI0XWWzBCMcvn5ni5eksd5r+vgYzhZdWfVc062YPi8c1sBlrIyEYzd86RS+B
xToXMka8Kw6sBiimx7qUmPrXZuTXoxLVHHBtQQmuGzhH5+v7BOvQCmAEiWN7
SK7WrQiFzOPk6lNdZURCLWJh0/Ew8Ntpj0fxD1XD6vR8Faupo3zntIzkqmmh
BVW60bjlYgdy+qsdjONbTIRBfg85JwpqM92gi9sjzKFrk0Bx/hG9QsOGqjmQ
JA1bIppK4utXcDVUg589uU6FSfWe6OkN9jYQAII/2Ul350TOOs9CamBR2QgX
mwj7FCPLd8hMzfr6/LJs2Rp/omdUGCL+u28cYxDMwNwqZehap3Gq5z87NzLw
1axjrVZ4KY5NoORDziGZiE7RE/NMh8m/O71wB69gupsNYThqKKOcJGi9CiDT
QDt+P844U4ozupass5BpEf+mHa4aWnJxVX/6Tx5ydIHmIINkkrWlzTUUE/BL
OgsFpgp1KyQZjoWdnkcBhrSanOQ9eu2EQZ3RolknpNZlSewmFH9Fm2HZaOE2
Nzh32yLnPGzXWYGAwdT9N+OYuZYtNtfawTrJOV03zAXlkBG97ljdjEmUoXIk
m3bQPMhLmms7KN60+5qJGwcQObkgoNLXLyJaL1a4jisTcjtyVGGa9jt2cDV2
9J0PAsCp9S2PtUyou/oHjbuA4948A2i504oWmCuiyamKUqfCPbfSYIQnOGFN
gbCPnwlhy9bEe8fVyfICh3j296SrvUNGT7CIyqnTMNhHz+Ffi9Sth3LFqyn/
yMdm4Dxe86qTwEV7jSZtEicDGeLVQHDhJE8h66FXH38ddSnRIqtbaau0kEDU
2uTPZrTlaQeW1btg81xA5sUiqASm+GP29jXCJ8Ypw1zY/YpdANkZWv6aGqxq
ith2nb5C+q0p54TnYyskgWXv7TpMLDn+pvLFF7ipzCtUClPIt0ST7cJNSKKw
SP+thwWMJBzZ6+FpXbGptFfEvToTkMNjFgYBgzbBtNkPegZC1ZTGKYJu/Djt
MVO5mJK1IMb9A0FdvO7L0OjxR4pKTwx5pXRXv0bfv979CffVceCnIkM7ZAzo
IijQxz5Z6HUjrhGnHvJ7ve5/v+I0E0yWJD3I+KQqr3GBRGk9eAm/CvvoGBWQ
515L3m4DIx1M2EhA9OGXB4FEsUlTHbVgHcXLj5EumOw7td2y6OT848aFz6Hx
3qX1z/T8Ordm+T6XicZi7AJzhhcVBGrEXRDWLIARm5w5ABYoe/yAOhgsLQiX
aA38Kmf93IpgPAMwTMXNheJ66HHOTEeEy5FjFVukrPaTV9Ol+ABugTKHYRGX
vJnBezvcwGkGDCta2jNBkVa8ltS8mQRWHGAmrJ2FN8E4Syfx0NQTinUeGeKV
gUFGiqol0GMcbUa0SSrG78Xd7JelaIUjFWYz8pX0K/E+DpZnfvaypt0qbv6M
Sg7AE1yoCW8GDlic1R2Z1zd1it2LQI74ukmQqtigU2ex1RURwlPaLrU9Rrfi
7nZQ6VNq8kOtIT0bcA/tzf4XjH9rNQ4ZTvVg3TOzRN2ZBlJe9+iuYrv2pGT6
NrirEIcrhrdF51hm6jxUJoGDob9O9zuDy8r2dTpcD2WNEYNHg9aU15VDM36v
PKAYnX1WqGawMC0E9BComM8yeK+crbodaDVxGU9XfQGGTSQmLHa0aFkMkSjK
wbk9qc5NpuVy5EANm3qz923S32/eqX9mQJaNNVvEMqPu1ftxg6uild0Q2PvW
3g/uRvELigqYPe1Sa/YgWPrXDVj3umtpMl1LdbzuylqggGwtBsMZDg9vn1+y
SwS8JaqUCr1Ub1w3KJtuFWXidDPNNRepehBYcbPoQuAtYbhqvbmfoffmPrQD
lymZ18atvYdzJyCFWzzotSHnbVk6Hm2gk4s2DORuyC8fbc4omBxQMO93h1vg
aTMeZq3v4ACKpLj1CgxFCkyUuX4Cn/eQA3eLelwn1/lrPl1fl8omfnvlNzVg
aqytt1z0K8009bSpnCkFkxVABk6nSy+nmaZUXQWbqHkefHPda+C659VYfFla
0Pq3gc/BOQ/pR9DoNv6/sgdmj3IUuxUjKnjVQmBXUSEFasuPmrFD14EuYf//
izE4iVbj+/iiZN6OGIiF5PndjuZhJ67VBYqrfmNRBXOtUvRkIeQ04XoU3Fc/
ALikuB0RlkQYKcoqpQ4NNUnPunBQrPhMvKcmA06xkKLIITdoJ3PjVkYxI9V5
iQoxA/d7iz4Ltacvs08LkIRrTCpDYpCDXGW9LcR4syxE8XzAn3MfN/0K9Jvd
PrLtPOhEUSjwk5YRPwmCu6xlxG6s9MSlBU7YzYg42lSUzVSGEoDDjkzy29u4
uaZ5xSrEeInPqk/7jiiLDrMskLbn8s0PzdARnS9Zd+5oOL+RSRq1E0sYQeZ6
KuCtrdwX70vMiDTyypgXpeHnltkiN6H4Vc+xBUpCDFY7DPEpDCi0sVQ1wN+n
t0oGpiZk39F/eqKH5sswZnyP90vlRUCPH2Hckbx2hQrgg513o877Jc3KEnTD
LsO/AMo+bVvM53qcupWrLXbeqR9OcA8UAmgppTZKpBCY+iVc1Udm7ZUQwdeM
3m7BgTAZHIPw4Xg7AzVabHKdl35KSYeJFiPgByYy/7i4bgW1Xp6/kJZFtl4C
WZL2/eklyb1SWUXkGHdk49WZKLIiRd6kdBkZ+Plv9KaE62uE5dl8giJIOq2n
cpvh8PPa8OytTpwR81FMv+l2F6UZDiTi0H95oQ075GDS9KjFLOqBvq47ajC6
bcvDp1WCJX8drRY+12/Rhyn9tNzMm79UXHHrlFQO4b/W+264vuFZ7dFIpun0
L2maYmSZEuEK85idL2rFPKmQYorpCapmAf4XG+07esGyXfj2HqtZgV7eObzO
YQZp9Ip93+DUXoGC4tK+DUy2LiDS2Lzbzqri4V0/CCtM7dcIhJZnqG5CjLuB
bQX8omEtYNJWsFPtSukboToIaIDTM3RlrWY9eD6sIi2Ezc1Y82zmTLa/P4kM
MLgWjx7xewymutdR8wnSyyNq1de0qZgs6A/v9dT+AHtXp21T/Ub0U8wJYhwU
hjoMnfoxAl1GziNd/KJAfbmb8BZFes1Veu3WTw7PbUd878dwvXRuO1Lf7RG6
9/7fA80nI6k8qeQoZHhZE6CYbz0DoSkUv+NFezx6hISX2gBxX379TB0QEBuF
1vG85hmpYaNmTYKMYCOKjdRmVwT2IeveMbo2NAtnBr+8UnGBMQcIxWqsCxsE
hwGbTQQKZ9b610vw763ac9sSHjfzoKZ8CZlZGM2JkXM1YHmJCG4N5RRIelXW
GSRSQE5b7qZtEhsZrTFf4c5a9yJP/QjsBJzmhxh1iS07YJrTd8xZCQmpmxUY
7aKrY4iU9U1hOnKJw0nS2Ag/6ewGAyULmO9CATDgJIaewl67xx4aocA8IPda
hvYe9uEgcEwRhTqOJp3gmwxNGjdZRCv1EIAHdrHCtLLLqDs+OEaLj5B0NjpD
zr2KajyTV6L6PB3K8+Ac/LNwZUvV+7ifpuf/6SIMh1ZSk5nRBOND5b9yN25f
cJiOpzLe7kAkpa4ZFQF06yjJYXUuoUSNESPMTKkD4lgYZSBI8cr2agST0ksy
iRzfOOEcGBaZzA9+3CfJOR79h1hCecrv2pg3rnefCKRAkOG3R8FXnnk/Cgrp
qZgI/0h+FEDs58UK/QTl9qIB/9TfAcMKFwjmFuFsCoPKWkya9ktDY8g6Gxq2
eIBsANChAcIg7pPph+5MA9QpxFG5/TcfZGFYQG2bnuxi4gEmsfuUZqUSAgTW
h2soizntoiqPVvQI4QkjFKDbJRVVY20SatYr6UFDDAsjBRl4qCwDoyKFEQCq
w88HW6g+1qwackdOv4gufUTEsZUaqBbfxu+CVNaJY3mhfq7MvKa1AXSesaWX
1gi/zENq11WiDOouaGTRLZFz2EQrqWL1kTv5GXm2M5OlY9nQJjCtUMjHiYcB
oFJLVYYoH3Y0zy1Q4M+OKszufk8A3cp/MY3so2F+pPSi6MK6jPn7U9jkz76b
NYKdzZ2GqCaEpaFDAT/mubnrTwsmqSHaPPkEAJ3OUi1nyb5zcloG0gPmCST2
dAqeMU9coxSfGFtD+D7t9hBYe27+ol8w/P3vkJeIL7JsuzqOD//OWfIVgjPC
rszefzF17xUhsKSR/z3/XDlsFBQRYB3bZYTyGim9NxKh0nC1Unv62UvaU+ke
6uosN6ar2viEohJ0YBXn+ITHETeV46WYdZELDgPMcLeyDQ6h3S/IUlLWME+s
28yzLWNY6ohNXPgsuhb2QmR93EzIhf+pN46a5auSiNDM3C2xjFuJrLR+17x3
dD4ETAUY3BI8wuNsPPO05E3zucRfFc9zKkITgRO7NI6Uy9d9egKhV2XHROJl
ofYNGn5THrtTzgIlPmDVaNE1LExozpd5VZbzFLJs4lvmsDMYB9tEvFft7qYT
yTdNkkWVo0a83n6POn3xNwsJmgo5OwQ/KNOgiN7WPg1ah6zwPh3Qpz3xZPG9
ZrWV6IWYYCyDzhvNljDSu3dx8NaswwzXnZShmSEzKOJnizvWMZg/jFKEZoni
WWdZFdnFdQcQkfwgw8/YhPknQEvttspUYFV/7yB+qe3Jkc0t+oDO1wxp0GUY
ewkkpdjsfKm1LjglBRuIUJuUCcZR4jhGIWOTqsDoSYdsXreucM9NSs3dkYww
m8wDxcQ8eUQykmPxZjQHIrYZjJW/lX4+QwW2iKqNvhxEZkc3hEXL0G2SU0+i
3NAR0O1aGcO0FQcBRbUvz/1PKelYdkFXe8snXyRo9FCtdwzy3NFhj33lFU2O
g+8hMDQnuxoT8qftyzQ8tq+Q3qp1ZXkM217nY7zSPDbB4wFq2iblWU+qVVz2
T5PYKLLcTxZNhKE86FAR7kbjlh6AXgvg0PH63WeZ5CzukR68/Y3odic8i/oW
o2gu27wv0aj3wEEgC1MUgz97oMdq3tk2whciJogsPn7YzmOKpSqzpbF7AT1+
8WTPoCyqf24lsh5T2tmZNZzio6dFduadrP6WSKk+O1pulA60xF4BN7z0yTH3
awACZX6m7mWDStys2AAmbbk77OjNKohrxmURLP31iLqL88piFqsUjPSBYZ9U
eI+3VTZ3PAfW5SHARpTfOPVKFH4lF1hw07e5C2fYGR/napy9+j8SvBDYdd/y
jIF98JTQTJk1Ymq2LlWfpMxaPSCvNF5IjV4JkM1WvWDDJf+4N5jys95IXXNS
fPAMswDADNLmK0+Fb7sBYxidnGE7VoiqaxX/0mWOfYWb0cb3oOxYy5ehT4lZ
vw/AFdFX+fPb5J5rUaLqlQqVUJH1mdyD9Nr9upJEHMYkVL296jgRGNg0rIVF
Tt3TgD2JxwhQ96Rih4P4ctKne36WK8KX7D+t63BY1cXM1sDjgGwBjuhI0scw
zMpDphR8c+p2/ZvNS/OAtf5eU2w5yw+QtPPAy5c5eP4zYy8IQIknYPhwok8W
QP2KV/+AMSXIvxMPmD2c/N6u2hsU1is83/aTVBERwIefOskVVRd0Ax6m8N+e
cs4Z0QaYC9Qtbn09w7nFaC4Ca4UwTcgh7j9I98azUPgqdMgwGPMJWIeKC0ps
TOGDrEpxyLaTxkk4yJAq0kSP6m/FDZoTzVXDOMdBGcUygEHeIjfOEzk/mFsY
CPa4Zqvrhg4Ewk0YEM85AqWnNrsA9A7C2EA2AvHD2lyAj7lJtmGH4hjOV+Wh
fX+Gc6wPDiLs+cokVLPAH9OhWn2wkEHPepP6PgTAu5T4X5ZG0xbtfyJcjljS
eivMOwYEjDl3SlAv8nuEuTd8IULbQdm7+JY9Vr2L9APEFi+LzucaXxFsied4
AfjIo6QshlUkj0jcrf6/j8aKsd4+WU0OSDBKV4cf6vrZgDM/WFzFm80t0GRi
ddye6LT3HVxmXi79fwMFKNssKO0k5Kl4sZn3W4gPylbY7SrY3jDrhcU2jA1Y
TR03ZJYGjmzsNOm07sg450lKi+shCsl8Dh5AfzKgBZE4il8TTr8hRUwuIaDe
paV+U7/E2lAS7bwS4dK93pk5IMiIWIp1qUi5CMiK+vi6fkMBxERzWvbIeAYo
Bot+Hk6FK/nfs/uIDoOJGOfcFJdJh0WknH1SAlhMaAhEfJ6ekdfeXyv43l9f
yzzJC3eOtZSDOSVmDDj+yFndwJOshcTp0/jl7uPI1UOJRAWpMFTpAH/gz4uw
eELHH/IqU/h8RsQrwliJA6ytIpD0rOZ9t9MvZda0zEoNVEPfsi+aZnBo7O7u
teZ5tJPqhilhBAH0tzRjKBqZlPMn+Y4FxHZPBFrcMvzUPIfSL49Vv4r5RGy4
YN9Srvmq9qaIsXss2Qzcn9aCO4QO0k/8m6l1RgImZWjX8BtjefwhrUmI6XOR
40+TYHFUxdRzfLwZIxUOgb+22ajfBG9nMb4AgrinjDPPq66ymgWhFXw4+yNF
+Dav5YJm78MesPgz1ge9qzWrr218/V7cUiQ31SybQVeozEgpcmilIhl1yTS1
WlvLcLOQoY79D/0WgL0osK92cnmFoW96KYe8i2ZYhtuYtOKhmFkVkBlxn0sh
QbbplQL2XZ1pegZgSyKKo2+ipOUZE9+Tf30EJATnR+g7xRxhNEADjib9Iys2
YsTCuiu0aiFrAOG4YGp2t7yHHI8a8EGNvuWwZijOtH+9nOn0Wj/BKpne3T4u
UPahtkNktba/yYJheJOcrH0EUpRV6WK9wCBIq9+3QWIxY8+N6j74tKtT/ufM
f+Tnj7UKkykHkbjO3K6DcKXDG2Nd7MXxeL/vIz6cZRXbhF1he7xLInTpAF4d
985mivl05/ADWg1W40kywI+6dThwMDc7KiL09uktP7xgRYQEgxyMQJP43/F2
2uhy0aXggEoMYzcj5oYScTKZnxbLS0H74EPbZUVReFsds3x0JJ9QH1+cpPri
PcKj9eFY+jURJnKM/hPUdTi5tW1HVyXJpolErAVLfV7LiPgm+ZnPL36uuMCW
8l2TS2aI582VaIXH5sSsSigz1qcF/x5TKLZlBVyK+OCfRd0RHTj0UhakevlY
2nYqKraZfvoY55Wt36z+K/OSGX3iBGnwvcXZCeyScJra5a+HiDByi5foI9Hn
EbPWSKU5/LEEsbslhFFfH5e0qdIOrpAsiNx9ly6ztjo63/+DSIEvgP9nVKDU
UZFAUtEE/N5mg+C8FTFK/DmYpG0Xf3a3m1TeysieWqqA0nKfRJrAr2GsKEjB
2ZwKQWS+7Sesb9pXwpNEithv4C455HfZbSbC0psMZNcCKxgTZe07AuRr6HpT
8Bkx+o0yQHoFbPFu5JZOEcgNSojloGxVbasYDGz71lhjdT+Fs28zuNICSgep
deecSgzRrNcZqMj9NcfYXOIa0PgqzdAdOQTZKOxJYRKBIegUGQV+9bn7a8As
aW1NvPiVNTckoXBYQ71UH2HbGBi9sikgRtIgohlHE9HWghyRkjKKk2Zlnpc2
SKCaJgqQWYg72OXfw/SCfUiGRFr77Wh7XZgGx5inUav6FkEsiw7eCnP6TKJX
xcIsGjM6rm04lI7FbXhdVDl75TgHYAUMqrR/Vsb4blBp0bJFWM+YXAYg4oHQ
2VlGYS+O6Je/E9HQmRPM9tP7DpaEQyNEhXvGXpmxJf9krzL1k9rfOxa9os6D
WPRcF47hr+iJEclk0WjSQlXmabgt8sUIQbLbAwQJEojbcXJ0T8gK9AQG60Py
7Q7jckOTGByAIShGIqjxz6NFjPDCvwLg0prGgfV4UQ6Q385xYUCOgZ75zds9
XQYTpUi0MVvXbTMCJne8pVGZKCMx9+qfxz5ibv0S3U3lmDwNNTLONmCSSPHh
LNN1shJ5i9k2zoUygHDBPIndQj6RW+b4my9Um8RPyIMnRHNlX13hhzjqQS89
RdjWR061YfMyWqPNHgUlOXPkPj5qeRaGtYVI6PQn+Fd4LA9dGMsM3AoMjpVP
tFOsDTZAVyjmjEwiUIOpDdUNejSUZmVpdqF53F9j3AMQySR3w/dalHPj8puZ
NWfMWSnwXBusNuvybX06+5VyZyCzNh6tvp16gMyChpDAYBPsByNvX9jBFWFm
STjhsFRrpu/ML4aS5NaMULBEPsiQwKHceckxveZHQCMSvvQDtVN8nfBJv1o4
0gJR6fIwsIGXqGiMKWImKg97sVpi6nQofdfqQwT2fdWBJ+2ffI0Jg6eo9Vu7
OH0uQyZEHsi+HOYj7LStqS+gSh0GrEZzy1UMrxIFooN2aL3+J3r4k1nnXV35
UP0iUNJb0hWYKKwz+vILvziO4eP8rvWGu9Yh6Cb5kCb8g+nOeyI3zBs5V0EY
vLAco0Z/U7Feew/x3OdspG740hPkpz7B6eGiWIGuZxYQvTLYYCMfC1qk6in0
H+0Gy897+gVrVinVN1kRebWHfr4WK+XK1mOa/jXm3amhOo/m6KrIFECGAM36
G8uBRbNMLTchFkOIOjZAM0LfugcTfUbQZhgudN44Bm10eIudYKgoM3Ln4+Rf
GHp3rHD3HzZFCNLacvxjNTDJ96DcpL8hYgV3vVKOPIjW7z9sefoG3iN7ZxlO
EzwcaJT2TuHrfu/LqeJ2q6rdiWOdMxiIfLnx2D03aH/8z/LhOcLYWy0mK9gv
vtNDESIg6Jw3Fh2gCLp1LGJAGh95CqKloi4Xa7dot967rMfloha+AbXUQNYq
87GuNb00N11xYnzxjhDCxJN/XHLhe4KZHSBfDP0+WEFZH3wCVTeGGpRScVew
l5JGUPssy7kIUKSPMEkrq9mH06c/w+bCfLHCSrkKOslmvHARDeYMQPTgVQ8w
Dfq9d5Qpz9BZKkSSFD5Rp19+Qd1GsBfYu6BSlQxih5S8WesFKBG0ZSYL77UD
p4IzmROLn+Cm86gNOUcR1eIqD8NY8KJFrKv7kd3vVL8XM556vOVGnhWGkBWv
IgwYgNZBcnmE9VulthqUuIfvUlUlyKMtDsSsLz6Z5JOvAWaKcxQQX2QIIU30
0VADTcd0wdF1O8eY0Z4r5C02+UtJxY+mpfcJ/PtDmb9YKZL6pp44kERkX0Ji
4W3nfFJA7HJNpfkaHOgE8cEUM1MRuawmaTnbLVGUd5/RjCvn/V3rPKVEB7uS
QveKEu2yiMlPFx/vyPA/Fbi7N5O9bUa8a6tJlXWNS9rgvrbaVxyRlguQaQvq
iSBq3AW14OSoeTZ/6ghR9Z53VWtWtmhsy2Sw4/3eOuWt9R4PjkAmQItPWnzG
MkhIbFa+ky+wsdYV4ntNGQ/1AqFMh8vUKIWaT6e+S9c7cFCR+5m7bmIbZKsb
hwBP+ZnsacJ4TUKY88wI9pN2Z9xTYC8t8fVYjC7O0WOTYe+6rrGk+QBMQFtd
94ZtEEg/5hC5ZMuZp02o8xPdwngTqQfct1rVpp6YAN8zGew48CNpiL8+z2gH
5QrJzDBPiLIiAYeQrYREYv+/0vVK83vgg11b4RfL6zSvMFdetTuqRbLCra7Y
sgRY5BGzV5jb3VilKFiyBZFHeEPXPomPEC5TgmxbVVK4/cZHJ/ASxwpLPmvZ
o3t24sz75NycZSFwn6VilAfDpzYPQjJc2FQeayqWUjl1xG/RFY0G3478H+Xx
aRrAxObFucGmxAlXt1lrm0ODph0BoDT5EwpCWigmBp2frFs7KaWWuigpCWdY
6xVecYzZLkLFXZ8o0wh8B3YObrfcMBalXsgOqbMbXwcy41YXYKRrFIvc9VlX
k6YpccrDakvMHR4pRykb+ciUI+uBcQRVzcfJurLDpP5JU8vYsflqlYFXihPq
lKLmp83DoenCs4fhSDmyD3+zAtYlYo2bimKg1Rj7uJb5jdsCwUMZtklBx44R
O+6YIc7rK6RpRmPxa/mMozYH4EN6qVr1iR6CD1DG5yqqcdsANv47TgaBajds
qFqEEQZTbUWUF/dWLR4PE/4MdWcioF6b0521v/iASz5oaTnqNJfBJNmPeAPb
loitt3jTo3QLOFgymMxQqi+NjYGKq83vp1KanFsPUIR/St3kYkvplIlvS/Ff
4YIuYSVcbnDp+cPzDiGQAxHh+DawY9GBMNYi6MHtxZUYliM/iC5Rn1WqmEPw
gF9mZ9JSjoLhyb2SN5JMYu+YDwwCRP2we0fDLNjl5mMOujkI1f9unKUnZ5KJ
+v81kSfhpogvL6qCG3Jmp7CVGbQ2Q5SyCjJ9efohhAiO59v62sswgcqzqx0f
ASIUI32XXmB9W3Qid1xdBhbRmSxA1z2HBOn/womov410ttSKYC/C93iP2WBO
OnCoV4SnifDvU9bX6jndM7u4Xfy+XSmEF8MUYGU5/dHJPwUOkqQbS02L9w/u
ACBgLk7CyWXMIjVI6Skrei/r2SFSDYgIu2wJ/9clBYE64Tc4C5mvJg7Uc0yN
8CoU6MoXPyNaR1X4hJogPgHEKyecVWy9NL3j4SLdEK5pk36jfF+RrMrAr1/d
+D6zQuz7Z0uNocUqOpmrZeJgBqjqalyxilCl1hgAcnRnPkBzDFza1D2uQdD0
CGcxZCqpHdAUf+Ksf/9FSEY+H6rc8g9hs2wPEOVw93ud1Ii6gS5S2yhWBW19
ryCdizBHryrFN453sJdWPEE2/aPvkk34Ao0RiNOFK1QGY7aaTOTtMc+gcs4N
Lvj19sRUfQ0qJsPhb++5eeyf4VGNRcAamqwHGFfiuW3vwbiTmxF99wQEf/zB
RXDLTJXiLp45kzTnBBmTFeHXRMjCKOE2QaGwoztARAZi3nMDRPsD6TTPD2/T
Io6fvG+N7VgxNt8o3jhvIbC786XcChk74snLZRXFG7BBI22fX2xnqPA7XzIr
nb/lssxevz7JYkcLld7t5xw0lZfqHHP8uQfXpsZIfqTR7KkpzW9vDguvP0Fo
omFBEplT6udRmJqmjTkxmfl+roAokZelAal6wPv5vFKTmmmcM61pPd8LeNYc
c5+eOnmtmiKzcGlkmJFa404FI45yPRAdicuiaXvPzDpfFFjcq4bJn0WNOikK
j0hGif7fdN0F6VV2LUJFQ2Rov/AHHe4Wl+n642dWwrpJimSQNOALSVZCuE9D
Mtw6P0d3yrwGGDM22jv2Spe9raCwtFgMRusWJEQA449enHbqpgglydqFxguS
3dNAuovCuRcEH+qo93LmYy+QYbiGMJud8CkoNGHVduKgOfVWKFrlILUGDXmf
vr8c81Lh+Orfey9pWixL0w/PDgfEUfAgnWEFKSiDUHySmjnppKcaQojbSD/H
9J/JPgfznhGS+CMr87Ue5xTqODPZear8yT6oqkjiuHUI6XBhvI/EVDRJx+Sw
UGnU8CMVoMvqsMLm5WrA5x82S60zF4eVKZBcOWuuPjNFWCRlGpbcX/JG5Z0h
TbvPaJcTlhzGGvzZ8n+htP5rRo2FtfaVjCD8BMxw5/EBsVs/ets95KUCVXwt
2wbI8M8LIgJ0EJICmBAKP8ju+nQgms16cTpu7PmF2atvP01UpdTy1xwVgFYs
sB29LvmGcUU27v3T7Y7RiIbpJz57HNSnEu4p88Jxz2zy//2DzGF8NkQOyd9e
dJq4zjsRvgqvwTxr0i8whScG9LbgFU+R4ROQ76rMUGB0uOrStXZN+c543W4n
q+TzOoLqkLxz8DpcIgcjDimHb6QlruUmCw5B0O6gi8uv+S/1+TxlYry9mK8g
go1sUl44QazkK35fWC9UJRjD60eFmPdgSatSaSC7NZokhvMRh1Hnv9mzzseB
lS94DIqk3usB8Z+Usz2lxd9+DY7Sn4CB2N76hQWLWITJ6cl2wtiQkkNGiYT4
IgKG4CaLvWsR3H67pOyos9Z6Po9/t+MBTcNhnOKrbOxcdqeZSlfvP9K72Ytn
X1E/zJcW/K76C1628ksG81iW8j+bhbRYilavlAqrUi2rVKLFkzGBQPu9kDxn
wA3hs4giZ9Qe2Wmr53jSowVcRTQ6dXLLtEI1zcmWTTNOv3Z5FGa88mj2oYYL
+LDOZeCPG9gabLFRcZiZaReHHzy6+csafdQqdkJhuM1hC+PGkLnpGJ72/U7F
1zdspNy1o/jFOmF0qouGdjeACCpdRRiiGl3O0U4axZvattzsWs1OSZkuGq7e
/qSg/MK+MU+gY1IWec7txJkwf/ysSyq4v7QL94okqX7geze1zzdx9rlDv1G1
QNDrz4Fp3O2hpaz4LI1/iDLcIEo7d/1mYFeW4mntMUFs83LjxCssbDsGFUT1
Yt56T5m9wYb+fO45NKAQoRuYo3rq/9mmOdaHjrOfLpAXU0oXT5GhMXb6sTXi
4OKrrUagqCRoSSQZK/dEF87OwtQzKVLVkL+xONf+wqmPilt67lK4+Q4CVq9P
iRLHaXDFpDgYJDBy66VfxqLG4hpjJ3kYkownVMUHJpsNFMBOy9HMJGxj+sho
YD4NxzYGWLqMkuW1Kr0Twcr4esJDbDwooQsvi5UyfLpV5q3dyOj/GHw82znh
U0FlNxNmkOPpItUaXURHy5bE5wlvmljBGLi+tPtlBDZXUtcLa032A/p7XD6d
t7kIox9tVowy68jYhmsGvxP4saslvjG2dcDqbk7fg/nckhXZRR9gaKUiaKAm
vLHRaXJ6xwkRyb2nVelJhT0G6KSL+G89Sle2AXI/IJZNKoV1RRrXQr22nf5W
PWwjdAA/knsAbVIPFLGPFTktaC3HZP4QCVq5XF+1JmrMTC7PNpaKydAVKG6n
aM3ccQSuzzKdvtJDxnBS0DtKMnaDz9Y2/2AfWhETapulHo71tZHJOjf98HZg
0bAN/Iy53jLwhQmfhtX9/56U8wwcQ93Zpx8ztnDpFzINlqXaH/J1y9w/zir5
tXa2yZCuqNXXTQ6x7Wz+EV0Nwgpm36DXYnsMM7wQGOCg/wXSysmS1wCy0HOX
bjcQ9J+R5ZJ28VNB+Pb+Gr7G4SWV3AU6h0BVrz1k5tdSHhCYWTxFtMerROhJ
lSlJRIjxmD0FxwLWyMJ2POwuUynibWVjQOoldEjkvNr3Sj5/Zq5kxGdpurGX
z/tsTAjBA7Ey2gmf+c8qau/ap3vbYqC9tHohAkcDIvVG4RaZUWJ/8UWuXIxX
d+tj9u2GwbX86ylxsaBlOi1zQONI38Gn6YsRkpX7uW6+/DXK4PVzUVr4jzRJ
ADp4+M5fw8o/IJ2uNlF2CQA2tjuQR6TeGG9wzJ+KP9TAQmtG6ozn7QKbxGZT
AZY0DjYUKM7c/yWRstcGiAIwW+YOkS6nmjaJxyk5h4a6tYZX9w+Np23eV6+L
cqdsiLJJEkfxwpWotK8+Unvfmg1/iG02WfhOJkgg9NfIreuOa4Y0b0+pZhoE
Qplb7EwMBqt81hXsspsULG2z498JfBmQoRsrdbruADq5mt1yIcHFuZ7LwFbh
44VsjcU4M0ainI6Ekd+DNo/rruu8vujSGEu15WJduYp6LPWjO6xPwxhrWdo5
Wji5lvmoROifVCGKqoyDMBU+n0KTdP61o1HScVU5sfTALyPYefQHKl7b17JY
l7e/zUG8HDqrl1TwPrSUa2G1pL2zCZoTeSgEWILFnRufj49ZFT54AAiJHdga
pzuzqrNCJvIofrHWy+18RLKlvkod2rX4b0FjTDuzIRvJ5/wvMocfb3vT7kxq
TA+JuXzUDiGUuzAiY2HVJP3+giWkc5OYilXIcNoGKUVnIzdlb7VOn92sGuCM
2lS9hAzkUvD79JgBlZrAHB4L1VK2zXglGBk8PJXH/jjl4GTFbRU8ZjlfjQti
Iem63LIKQVOqtASB19cVVqm/1QsA/7pRSKCMx5FlU7LzOcL1kydN/p2WebO7
sIpoW0IeUoWKJ5H+/xOPCB4P5hXPI2tRTcoKTsKHUfAIWNoGV/NL3VxMiuo/
eipuWosv7Slmwjpd2tODyp8chCdd7N4jPsdjUKUB395DQEvHckXdJow+X5Zh
vq59TnKFbd+vPy1IeQkAxy2zHL/CFzxswYRAheImJcU6Rej8DheMfEFZGhL7
zsTTIDG0uYqj0cCWpxBDluKajjm8GM23AsVTDt5nH97EymgfjH7IR2vuwWse
WGdBKF2ca18LOhLlpm1Qu/YMb5VpPIgPHsjkIgPy0PUijuUy00YpmiWFPZvB
xm8qqyKTTI7ZdpmSCcIy7MnXGHm0khN55sQTV5eMNrsLzMFbhCwmfrT1pNCO
bT0EwUMJaUwz+R7Nuv/y0N9YsSw5fy1Kr4DDuJP+1P6Jxi9Jx3DpHeM8afir
5x0lLVg60GqAP7pREdgrKb3fm+ZvNF1dfxo4kF1kLqIh1FsyTUw7sbPtSqRi
ltfsbbox536lpJupam0gXFyPoO+VBM6LiEaQQhIFsll/4tshrzEKxK6eCieW
wjT9gafBEVP3f2Kw/y9yUBruVk5d+bwiz4HMT2AIpeuXstTLCBmi+XxFcj34
SRs9TlcyzEKC/qeKdyqxNtIz7Ky+odYBjGgmMltF7/mSiyujtwOK5mFJedPH
BV06DTI0dzMFuIQPNi5/soa03zIYaoDpBnm20LAaWqd640+Fnt3m6AsufRC3
/3UO5A1JpL38ijuIRBRbseH6EZvcDrM8Dw/pT/EtZC9yF7DhvP5m07NicBLX
weXVSnEjjB6mYgMTJs/DnVqkQbkB66x7aVl01zHXoyz/QiLxgeQ7UxmbluMp
45LcA0hRh2hEUcdrr3GIdHPU8iEctHFrclm1HXZmy4xtlxMlNUOutKV1sSRC
FsrnhYu7gpoGSAAPEaWfkTUeLi/Pua+TwqHIHkw8VwLHA+aZHELAvlrpyyPj
Hv7k7T9CytVev533ok/T5KMZMSwo+8fgyd+mRcVun4ySi05yHerOsCpTYIn/
qUAzTl69I/L4b2lAj1SUhDt1h56qkMeXLhCOJF3/Od+uTaPlNtj47WfbsIe8
7dNrvOfkYZG9GTSUdYhvrC2qIu2xceVNbe7nJxbYqKYqqFpMrwrlMv743mDJ
AsAWOePcl2FSz6xvBoWESIacdh+7iOFOWlGcmT9Yan6Otoikk4+Iq8e2+t3g
QfTmrsffad++VAa/LfGnC3lv+gCTB9ZyYDtAr2ulvQzgMpxQ+hLcDWhGcP4S
9xFvNxYtrNntD9ktpXPzZM8W1OBD2/EtZqCSrZLDGwdNIjyMbyLclPczavRJ
ffYvTeAHkBsGAR/UDyDBGX5s8hQPkj3VqZLAv19MgiSY7Vly1NK0SHcUpfkQ
PixD7M3ObbpgLhb3apTBAQIAqozf1UX1WVs68zvN78bpnrQdqVGiosm1LDAR
IqRS1lxjRGTwpB2tUe70Mm0CMPlXnRRnplZbTyJekh/aabKcJ8aKTrd8tsjQ
Jcrcm5FvSmVYYoexksvpS4Aqfgsix3ip2V2VapbofoRddl2acLRH3ipUcwi4
VBvbEoCzJhNmKufUxIK/sGTic/Q8D/zvcYtBz0f7Ln5R7XoA2Nth38SxaQIa
MVNGmNa9qa7ZGLqlDOfUTLl2MWzl+SIGEvIIc0aWuVP0yppD1ERujsR0L/e+
Y1VW7RdUPUCeDatiZ6LqQGAV6IyRqFJzOFihunktLqvvFhmcFxWPxda1eG1y
y7f8ZUOcCQkumIH7piQQ/ohK+SYB4ffcvnuYWcD6WluRLB0eVibf16hktQif
Sjd13fHSAM6KRvSvw+BzA+BD8FsOicoDBImk819PIpH9N2ugzzd7vv9bChJ2
R9d0E6ndDAi+uXNtVY3hWFIk1Wpmq0Wgsb4jX3442MHN25gm4rL8MUqmyonh
/5Mb6klnWqa+O7UnUsMKWTEwWL6BySdF/WPIxG6l/Hm+CMIB67gPdXwKY43P
1O/bIT0idKFQD6dzd9IGJjksNUyVzNlV5XYW//gOQknnjgpkA+V0o4wUrzJq
VOr2ATh2Ugr0X0kQgxHyT4nVlsf6+6/ELCtUe5ukt8E4RjBpyfcP4+Isokf6
l19jmg53GsF50lqc19gqNp45quUPGS+TbKcIkKwK3aH/u6H2kMV5eDFlaB2T
+eLbFntKNJS8U8mZOnIN+Le8VYCeMkfSi399OILprdDGkwol5chcsRivHpyG
bVpQ/iVVLjEo2Gr0AXdj+SmKw1WVBQJfJukAPb37zdYxN5i4Fu87ru2cbINu
6EY8MMdfxSd5yag3wWWrOmPzcWxS195q4YI+8HgRmoHzwFKJZwfmkX5gE2vY
s+YVSlFgImQkuJo1j98h7J5Cs9Jgr8Qlb/LDlCffatCE7Jwlz8uN0WNXX2uz
7XP/gsARNnidaC34MsDrrTUeTdQbf/Z6GcoLawZeECR7Py52stfUVHz6sGlK
zVks6QUCAkGdYP+m4b6zRx0RH9uLEGKX7uIPkbgfZrVFUbV570c8KkgG4Mj1
jIz+Pmg7rzvwQIH76sDYIun+Mgyj7GSeCZiPqtYMBgJxfPZQj1W9hExgTBWB
SG9kGLwXtZ1SlYyPOwnBL+JVysDVpJQlzjVoHn0ma6VCbXuSw3Y8PzoO6vMp
aT7OnsdnXvohC21zoEV1SOssqFFBvcGY+t/E2xPjAJf8pNFT5ViiS5GG7sOQ
l+L/h3ZV4dfQgwtRLHiZKGVyOy4ozcVjkWB2Bk+8EW8vismXmo9g+b29AlM+
wL+4rXWHTfEnLugvqVgaBPVVkvkMRIHgJcTx9xgYyKWLwmVVaKDcaYk2DATS
bBh5RdKRgZPQvNFVb+KWGJKhzs0/a7I5z6HKq5la83jNLdxCDC6JSoNzZxYq
4LO7iNK+B9/Bumso+bUhcqIBBv+oUv7UbFaJGtGm5SBXn+EEDlgaRdEERNuZ
Tb03Zblh7ayAWg+1nT8qtYXSzJpbFx6LW6LgkjQOSyXxI8OPDh11f58w1mZ+
cBaWOirXYxdRUTqqqziPfX50e0Zkmi+9kw55xGvaSaVXLgcQsEBPsumMwTsN
yY6qUMHh5P5nDRaAypImaCrDvfmfLozf3dqwyJldwQOPwxpstk+AeEX5AHWd
JXhLi8hYL83BKdZFUOGdYjkNMc/kXZFEgGJc0gddowgs7gQlu81q/jf0WV/q
js2QpoPwet7dSxWDcWcPJIM/mCcLMVE/CL0+MaCdly8SXSacTAETxKaQflyx
Npnh7h2ADTKrJSrgTYW4OOtEAyELPWPcGTuzY38zGElAoCxxTvlHonraogUn
gLw/VvgdijzLz/h8uYiCdJRMev/+5+1NAQDwMsDy4XQBzeNYCABEeSd+3ZQ8
hgX6TWvC7BO+YZDCMNevWRF/8+s1S6LtY9rDTI1Mw2rhA8Tlbbppobxv/l1J
K0qJ4sd/nYq2v2LMLXWWTILUjk1/wkboG8TrApbxCuO80XQx6xTE+rJGJyro
iyJ0kZB7s+DQCNq1w5Y5oehiuo7NP9DD6M5zkLKmyjiMGOMYTCe6G/1tbnRB
sGSxMZ2fkVFZAubyT4yth/oulb8ueBBBk3qH6T7pvwuBq44Wwe2uGAZlgeMJ
xcbwfsWhGcRERReHn7Gn67+dk1iikKSxLJOElvhloP2+oOj8OfZZlaSowbAp
r8RatYVH0Z2mpakRg3LFKx2NhJoPikP0JFQXlHNnSHGkJ7pX2N/uBoZvrO7A
hOL9xNv140PJeiuSIDPscynMo6Mpz6Ag+XkxS0seN14QXq5BXBgDRcHwYRF9
RaJ3s70ZRN3lNql08mUph+SzHPcodQKTeAkQ/7kOfnLKwWFMJT1I3JkNeabP
mPZJiwHM5/+vNntDFt/97I6Qpo9msMOTnO3VslD80m9TYxtOs/izLkHsgpLw
n8A8QATNYzy0yMyNq84+NqMH2gs2hNRafg9L/PNVRPzvInrll3itsfs0kZnm
XZ3kcyxiFxiC+QE8cU8hWNV+kiAva5QCFXnOFz3W9/dcrGfq06knj0JXkO4N
ytJ4M6PovodI8y9M4D+grOua+E7kCKyMnIksoUnGHM8rH+wuDILPZKxP5cbN
QtGO7xEszf3JuprZE/zPnziXYgjcH+zcTXZoumiRCo6/iPMAS1Kz0ufqyaz9
gICLckURLvwtPyoQNQeHggt28DRb6mlX3VuN513MqPdn4K467/ZQekvGO9/F
R4+LWzBZVNuTA2F5xNpwBc2QnDCI9UXd585TWrz44U6t6Jv1CzSOU9K1GLi4
WK7AjljU2AS/i1IV/EKAytsPKUJl9pGQgWB3k4QMfKL+GqtJ5m+bTqdJ10Dx
pu/zxeAU+U+UxK3oPgRgOQPMyRWW69wM7Eg7qpX8VF6ZzyXc3MYK0ja/RPp6
tYc1cxmJyld/afiQPS4yz1TFdzPu4jLotj5DpZSofffa2NMq7ns+6aF3d0s6
uWlJMQZ2KzISjqRce37CZvGuTg3S6s0bg1NFIwXA/RB2wDpwaYTmRA9xzOyY
dKfU+uqYYA1dEHTbo8XuxwsRk7966Bko8W/YV+hWuFs1eg4V769woNdtFB9s
Q0a8Ypbs1AgGELBUyYxMr7sORAK/lUkf7OcnjHmxkOa4OaE+BTYkAi5QyaUI
3q8Wv38d3AneWhXNAwvt+pKCvUuZnFhXR+ph5RI+yJPAvB4xw9DusNmuRQ+5
708o+sGj7wadMR0Ae1Uh/1xCVQb6sVd2MY+zcNRA3QUlGsVeCW+wfbZuHUDo
vJgmu/1CY5n0rXQkeUoK1p8UZUy32M5nuacrG51wrxInsuD9COzT78l+AhAt
l1xSKe36Hbz4dEN1eBecHKvz+agUxG2rrFfYH3nXTimH8VUuVw5PnCyXBWBa
Lkuo7/hTxTb4o+gRYc60Y5gO1/SDSQyUGTB1edRZ+512pfOq1Z9xR7dYgMrp
BSVmQEWCuWoF2iuPZiZ46Nss6J4zamCQ3swBE8CeeBXbb2rMNq9J96DxTU8j
e97NgiFOfOo8DsGK3G+AH9SFnn+071kajPE70Va5H/kGBE4JEC8iIB3NsEz3
iGOVON1AxHEc2yM1GHK73J7ml7poWd7l2PcBLBSDd+Velbx7SUlRnw39AZ7i
a6CfkRMxjPbpnSoLv93p03a5Cg2uZiD0Crqb+k7l3s/zu+GQE/r7EnfsN1DN
D+kWYJTWMK2gazlf2WEwKN8TDlh0qg9vWj0DY+NvIzYaPbqGpi23qRtnTeij
jXnJnKWiFScQ+Ty1NpVpV0P7udHm85NU23jM239Zng8Bo21XVj86SUdkXG7C
yTokyp+RHSYQMc58jziTWXmezwzU4ujcgzgJhlWR78xQoSGoYGW2/lexcGcm
2xU9yTNKGmAGM6f6cB+hGq4WATTm/17nDpjIuWazjP0nrNLrdHhWQoYT4G4H
mUzK2TZ0qX5lATWgNZ+9hCXA8xnYTilUv2bn+B4qTL3ULIjHzqm43WLWmbb5
A1/eQai6z50HKxj6yLfL2Pib2Kc+alNRXeLuGH2f/JB6VHWGsimkZ7zEJzws
+vMxfDt5F/atjTtEt2V1M9S5xrdZZ2kUUyoS2VkvIkRcpDBJ5bR5HkJ0aqPb
SQdXG+htZ2CNUxA2/99ML/uHA+1p/r0ZOIolLZcN65aBlSqFUWsV7XuXjqcL
T6sDX1/NpIYx3YGlhljzg4F/lqEApS7MnLcZLCIS15sjKmgNU60DJn24Vkdq
mb1+ZJvG4wVCH4af/jyNqVQ/35itn+8opImnUIXLYaY0C9YPcsAmbZdIdXCU
5AC05yWAFzYMWNImhbT9jDPXTE8WO6WdmJRZ5+g3qBVoYinu8Y8FnHjkC/bw
GY5ZAN8MTgZ7EXaxrZLq5X6CwKX5bH6DgyRRx88zR2N7P6JDp9SeIIBvsGRW
MVXFcnsqCwMTWtPek1HArRrJdyN270PMJdEdTPI6zXaJVYr9lsVa46rOnz4N
q1vl6IQCEA7f8PpJaTO70aQEfg2syN75HFfkl2JJTqq3DZIBH+1WU3n/QYq9
mLfTCdW/2WFv7VBSePhy5NMgpn7DkBTVDq1vXVlG/1zV07TqcpbwGKVk7VNo
08iaZMJybbsi2fcgXHqv2sbu+HHq0v9Du5DWgrCZo+YArfWSBrW4MlkI2Dn9
KsIMWL3KQoBcrzmMbC91qqpocU2uij7jAPDC8jQKHr9s5MP86icd9Wm3ylRb
2hHfhgBPnEVh3G8bJuEJLWj1mRNM++uRF10FtJXqyIqtuccGJmdQ17O5dPn5
OHVtcHHbRQZN1Cn5rzi69vCrt76zg/Yvb2HQaB9nZZUfT5Tg2g1HMlXIq3KW
42cpMugaMQJqZtsXbKYN1nbHUZCJKbUJbrio70/yeiQUWK6FMXs5X1/g04FI
n97NEp3oxW900CiZpw18aYs5Txb5SJxR2cWjNHYNK1UNyidhTlkrPtGze4oy
WgCd0t/boxdWVHvanLd8xKgAtNFJT3oMiVD0Awv6tOBBV2+8oPhtR+xQF5D1
TsWCbrgEOEe6NSq1xF7fsIYPyqob4IVtuAGL1AOPyGFt3/mKMTwmoDXlBc9J
6oS31vcqmtYn8AhveVrZeqyqNpUJ/Fl1VDbW6cY0bp29AeEGqwEFbtyyfMnE
OxYaN0hrV68K/LsJiaiMV4CfukyiiQQwvbf/RQfrmzRm/Ghe2q9KE4rXfXTL
LqfLU1mqR/4p9mFtnGnNhoPArJZSCPT+jBpPs4mVPoqvzML7g75hdwNOwAGh
2q41uo9jIatN1pVkIwRFEZu/hGD0YyRhJ/X/Df0NpZOXBJIZNhiXA97ozPw2
jcitJ7Brxh9dFZaURWbti99rYoKYP22uFhqBrMz6A/mAsAyvBygtx/tnhEPe
X0xLyvEb9smLaq+bWoSaapHzNVzPuin5HKP3G68HmsDPh4avn9wMLUnIyxCz
njWlvhgxqZys1wDlU0Vp3mtbH4e2xEOtq99ZIZIkvLyyHB+VpkxVSkvEJKxb
A55Y1Vc9D1rBoWNuw1AixokKZUbsWY/JFkwcOCng2HXJSwGUJugQdjj7rWHG
2KGbNKNWqGNPsQG0ncmIvpqsQxB8S1QpUAxVEdHMk+xYP20pEc6upFHxKjQo
jsLoI0eAiO4clBy8kBF38X6bs3F+t7XIh1yHxxDDvkmwFppWbT1w5rjcldIc
pr488zwxYGvz24kfnBh0zKplNmfyxBa8C4577QnOyihUEslLXdnXEFUL7O4c
OTvOV9DOUyAG9trXkJCO8xGsLn26KMgRvnJnF/nBF1aSE4K0l7NbrEUVIKdX
KgoPl66rT9qmNCLoWiuj3Bj9ZDe+L/NrRFHJA6hGyELD0FQoY7t91++E+Uon
2Xeb4H3HtzUXq+FJq/BDN8myWiWKP6uuJTO0Lar88KRNUIPD6jPcFkdUSPhB
xkPST7j+XX7ujPBHpDhMu9c68R8tX9T5tjTPIsRCDyH9N3F9fz2MpR/urlt0
DJCUwvnv477OldlJASajX3MIjNvhdi6n5dGxYYYPuZHleqIc/+6VsPY5OclA
ug+Hk7dbpoGeczwubmKQ1vGRm7rQeZlnMw6E8jmHiPWNV5nPfdhc6T03SUC9
Yu2DoSBKypWiDpGKIO897tv/7fmpbp84Wz9rsRhEeBC7KCjDKzW0H6FI2rh5
1YNBDmoFjpYhQP/pzAw+tLZ2XS9U7gZsNT1btWGuVYTjuolIuc7f/NhbtjaP
/MhZpyPZS3aYeFGtT+8Q87aoCOPqZf3onTaEEs16+pJwaMVvVQOR2JSo5rYN
OOgg9bAbm9pYOBpNRuIuqaYJBO25xWCWyXAzpKBdFHFT6WC4a3vfYBPOgmIs
1x8Qb9DSCYQ8lcrOqh4OuVohlIWf93LdIxXJwiZ2MILG5e3qFnIIki6A7T9h
+1ZQBAlu+rbMngD1fH8Xuom2psMNYrmQJ7HQQB4URA/mXME3i9NhAQRx+bb8
nvk0uBeszp4v8dZH0PvYJ672ajBXRpZa3C/3fXn3o2J0TW46ElqZFFojkPSA
h9jQveEF57k0+PtkUQLxwLVl0UOh9FRNAlX4GxoTL283/3bWfIijtNRjyHNP
5L2WY4hBvZcqicOVA2RG9xPZpgprnNhw0rqpTm7+iPGXw5c4olb+kBjbnKmO
wdgbOAS3Yud5P/uEemrteVmC2K+JbYoP9l7P5TXCmPOYATiWxoRF0aYrKa6b
G5fOPtAdqjAaHYKY0zlAgnhuqL5avUVP/DClxj0s04OioNz2ty1zqkhd1Qxm
5s7/NDHDpedeN8LuB4Vn6WWkxLil7TrBXd4V1BLSPsQEvZaujT7OAExOFcUd
D0UFkMnoPOx/LeUN1Q5aurHE4PvlY7USo5eD1+F9BhFsG6R64MF7hkiOL13Y
NICqUOiV1P6kc7Ypwft5WU+1v/tuQN7/hbec2fpvL73PzdBIA+EZZ5kZjUrM
JozwV2mfwBDpeJEDl3D6+WgPjhD5vlg8sK/XuGH9lwb0LdR9RPLkw1FYzdMG
gmokmu/xKjGddW444phu/Py1Gwsor7iLBJQphHifjKJfIe6/q5xTZ2e4I2h3
vIIQwICFBPhIh/+28pP+TTDBRE/30mFpq8dZ0vLZ9A7Sz9cCaeP/jPTMeclL
WHQxj4vp2rQx1BxZt5HxwdIcDxpQSz66wAJ1XGZaYi/hC5MbwVQ2Rl1BiJZs
vV+8Qy06OTRQ4yfVKlxy/auxspuYMyTp9LV8v5Vv1tMzt7ilbVT9O2n/U6b4
8+6zPKHwmEJ/I7VuEvv0eDVYOX/rz0/n7A3JVqEndJpiX1j2fIZYOeQfZBlX
CH67mtB7HqSB06gzd0pnMUMuESolW9f5Ch5B4o0dIxbbaoWEI7kaf04jCP2o
Hg8hyuf5nnb4JnSzBM1lkz+Ep1KfM9fsU6D9y4lpZnIdNURkhDfF4M1sBWfC
iParH7oifMeIqUoH0LGxnyDCo3aUybbJwoOMbsWU3SuOowj2C2fSWEvF1/UJ
v/VDer1fMC0Ak/yuqE72fWdqRAqUouGq5vapwrSJvx0aSmY/epdvoNjXjtll
cmFyC0qxkcp69tNTgNKH9cxmCRPrCq+0Ia1mfZJxOCnwtnY7mckaiyRyFGGh
SOMYtjzrPkQK11EVk0fv/GYJsC8vyo8cHPQbGXa0ubBSdM0wBXa42+NmNlgG
L1x68bnhAs+TwtWC0vdlxoInowDlpBxZJyVGUH6LCdZvhnPEtn5mJ0ecg+bP
QIqn4D57QpUOlS16YdckfNCkyZ1cVJRVtH8tHS//yTC2ghlgoY/pkQq6unzH
t453O6odGwxRHoOHSciYI2YuFiGw529W0TYw0D4KKdfuTTUYY7u+/vtb3RYG
L018rf+z0rJTTuT/bB3s+HE64zeIPa5fZRUe6jL6RmrwHocq62zVqDfiQkv1
FxB/hHnbMeFuxrDhZzJLyMoqQA8S7Vo1J/IltLZSJG/QnDoMzoHh4La11oPh
nBfVNDsR4W0a2a9zOdDdpMp/t/jPjBJdRg7xRGo0F50iVA9xDQFIIFqj/8Ls
be1jsH5QXkuqu5FMSzV0HXG7dwwuPQBb6xNStekVLnM0/988O7g2NigzgKjy
c5uCkbA2kwjGINZDI+4bbkTjqpVmp0jMqmzO/GPFlu2QZUilXRbzIbpNHmTg
3uVomjigXiCW6hJ3rQIdyh2x3fvpORMhJsUmUQAZP5Jp/Ew1aqY5iTJDeWzr
na7q+SCbic7PoU3/9HGAwS9f1/qnhJiOy89O+PgI+4O2eUaBnHbi/1f/AV5T
pFO7Q4jrhqaNhhRNEvubz3b+e+vip34VXJtzPV5Rzq1CVjrmw6NuBHcXsZdc
R9grmXmKkGpqDrXLTV0GqmpP4DsjJxaxt3o2PtfJqaurVmN1dP0DUUcvTHm3
+Dup4PRUpsWm9E2s8+k3Epnb+Jk1DDFTT2ATBmm96kTFadniBWkakSEf9dFm
D1hZ+THCCc7SNMjTjF2K7aMEkaYLRiOlK1iDlshh5V/ROL8HDS/pUwaJ7kio
dYr+/rVRoeNKGt6jpl+yJTLzyU3RoLXHM/6BcMsGbpstbd/PAaCV6eMHmYE8
oCysvuqReShvzsf3yJRYwXzqglPCRWCwylq6/922sJ+FeJ+uQQ+iQQnFN0RE
+6z7cts1YH37NHOOj7kSILSjgnRHASIQafTzTp+8a0zs7DN7xAknKSjCwtkb
tkr2cPn9OE6UUrFDESXIbSpOO9K7QNy0ATtAEcOkP8IIALKSz20WqfkG4S8f
EDLRKJjTWhhpYk83pPMo9baaHUejyLrd+NzmWXqKZK8PFo6wOdLRXMx2QRBZ
udc0LIZ4/FfrEkAg+fTBwQOzxTATwfmor6NKQXK6VDG2RTL70/oP81/TRPnL
2DPyNynHlAP9UDfn/qAX2Tne2osegbPYZK1grouvoXvweyHMteWVEO5GKtQR
iPK814V3f9z2Ews3V2Tn7jvfC1ljiwM9yyvCj19Bcuxa4x/mvG4bYBh9f+B4
HPzpKrYvO7qFHM8VwWjLb4IqYr+2ZCC7Ch/7RFszQQtLZwo7+7TbXd88oC3B
G605a8allPsl07vsszb+lVzstDxZxr5HNkO+Jm74b6/AF+sPV2E+cjtcmIL6
6Jiw1LJ7Yy1cqSnludnoEZ1AqxjXH2K2aR/zOY70NHzvEhaLIqCbMuDvDRWv
v6z9eAN7CTC9BNqmaIR9BF7nC9mJ+by6qyRd7x4F5ISUGx2d7kUFu2KxcQQ4
87AMGELtBO7Nx3oP1mCg9z8aFIlg5ZS6rgCrcqqKOKU4s6DLjiKBtv000P1D
xA0A4VExGpmMhXMPHZDa8T9mHB5J494jqO2cNVfWPsyJHSofJ/RLUCiPmqC/
2Ai9yBUGfGNzkwbnHJ93kPlyVHsBR1TWAnLfbWVLUsfPhDZUbV+mVbuN730n
hEj7cfZ9WGAl28+egQK0xM0PG56HAdxUuZyETVgBKMppgxArXJ8HscZ5o1QI
ez2mrsCayHz8c9eTxsX4Y/cegCR9Q6vI0IcspK7UMtAGXklX7QWiuap8sAlj
z/o27HNM+bRrH4GvfeQouI11iPxf58ZubiV3xDs2MJwGojf6Lf63OjAfSrdH
tx7epuDi3WPWLwEj9A833fWlCqdbXaQp6Xk7cEkVLQkm4Km+H4cpPDkPflJA
ylxJpP5O542IelhZsKdlqI0mdK9ojcqqyMDKI8zZxk4dREiqbvK/9YsdTYWW
0evqU3AZJ1On2kyCH67xXDZeZNiugGZoljImxlKAYs8Q5DO2V7L2476n/no9
dWc1qAhInQcVXiWNiWZnrJKmmsnuVEIqpj1CMUmvzJgbDFkuHaxtuZM5UOAl
5q2m9OoLF6IitAzReFsSpdxqMGBFbBKQ2kgIXshx1MTcSyHc3zEJHu108InW
4qnGAixPMynMd3+FDB/PvWDF9rfe465pC275K2fx08ZPtzNPhZ0fT7xQli89
Tg+2hFV0IbSwyNGF4gB23B0PdUmLWDHSclxnlvbw56f2CyOEAwmCGvdFCSLD
OarCBaAaXYV4RT01CEPAT61pK1wB5YuveGiuzLaaz/ZijhL2+SDU5+qpn4X6
KQjatiIIoC/uKmtu29ONogRLxOSPLmsgJvuItj9dH1Lt/MIrL+B+RW61Ofx2
7QM5w+2xxNVxjijBlyYd91dqxUrTA8TSWyV53rX574iXyB1zC8CQ/OvEC9DV
cK4uNsaOg31H0VzDo4GuekYr0QWPSj8m6KrwfZ5i9y9CV4uLjvXo4NcsZu3F
FCJHMQTHHYH448haRpVWZlJV6qrf7H/ozORU6aXHnRFWAyXuI4hSc8/B8r5L
DwkYMLQy0mj/C7P5RtN9hw4deT9ZjaNpTJsdfBdhjhcmNMcEcGmh6pXpedm4
ckjSSsX4wDGHZVKjvsg2BNoYWpRPLqomak1RE8KPeh1pc6aieH1ACUmq1AaO
0U7Xpvh2LOID1f5BfamQKi7L7Z9/8/C/GaCfdZngX/1AT4Rym4PtstgSpdGy
XSpKW64Ti5EQPg9+LYny4VYMjGrgi7cqA087b8SjZ7aqrkew4GEdNpEJ/Zrq
viUYIRopW7iuTPj/NgqWUxDg6Q0Up7A0r1pOBXwNKPuvSKqKzHNMJ3SuzmqD
wssX//RKmRDqsk7itHAJtHrK0IbAqMDsqOZnUxBYu8PRaGx1TJNUcClG1HSv
l+hMXP24WCwTJDWuiNQVOrXt6DpkZqgYQWFI3HhrNoQv3L4xDIE2G0Ldv+fq
raeO5QMZUbwegw0tF5z+C/XwdemR9jSTcTppbLFD0D+LrFMrqKv4fchXCu1/
3zYK4z59XxLp0Mug+YVG/3yU15dO4aTtKDz7YIDOiByZyYb6C1F/m0r9vunr
uamTkwUHfFC0pL2Hv8Bmdlm+6TEE52OEtHDE0z5hmw8BFPYvcxheu/2+8P2p
cy83eYnfe0k/vT22qkxmoMnZiO+M6XN6zmEDiowJ0dOZ1UKuTD3p7PQ/tvuN
z1t9mxOEtsHwavbJ2VOQ1sqIz7ce1XGW+FuwiUnSUIJr9e6WsIi3L2UzoJ/G
SQCmsxYOxIYTGfx3zlDk3O2rz9Wdg9Q4MxT6JXY25syCsOWeDk9M/4Bbumvm
BJnbR5D+uCoOaJhLeunTaWmGiWUP7SMVYgM9796r/bf9zhvfAxgMUkFIqgin
b35DkLQCWRyEFMnKXzrKTawsX0XRqq5q+betVmJPzUAZDHaGiHu8XjJbbzER
jchRMbYFLlIkOgBJP9KuEInx/b2/ZV096nP97y3ZEVyeBv/ZwzDF4IJU/5wU
qSu9PZdRYHxL89QH/TXDI7IQNYj+EArxWeplB+w2ol0XY45n2KePBnrdVC/N
k6TBbRoCQWWZWz/CusLQARBsAk/yqg5dHGfUU2tLhL2tpCWPyifENHWIWwFH
yQSXAMuOH74fY42uNmTt456fh15OcLm6dAtFBZOXXDJAWLLbEerN1SW1K7Gl
M1yF49KbpaY/fSVgHfCC/TGtm2uD11DXD0s0E9PUQEQBgH6ODfF+L+/JOpBJ
nCX7NjDlDSOHRwKOslrDq7dSxt6l+i6iVP00C/Gli9Liodbiy+qIIOc36Ons
lNV9l0ifiJvUNoRi3KDaEVctrWLGwianAY0rt9Ie1Y+zJA7+ugvOyewTYLq+
9UF/6Sg0WlkAIWu928iyBcAT90klDwPGE7rcnv3CeYdjtE+p4W45PJn8Ofcm
IFx/85RrTjRIDXOPxX/Vi2CNPxwP/Gpisln+fJo9mFmx48AVQEnb4LoWSoht
dzzAACTj/Xn8tHaTffZ6PPR68k/15CIrsmrymGKm4KIW9XWemyHVRZ08CeUY
ptjGsk6aEWdDq4UhRkl4wfOgLScA5UXNFElQA1iO8X3eWH0xh1ywvM8+bvbh
O989YRjbJEzR0r7fY9tyFtvh5HpV79BKUzWIAy6Ex0Dnokbc4XY3+zgrjBQd
UsckLonceH5lnO3teiiJPJko1Dpa10rlW/0PNlJSCiIa5lR5irGH/jfoPPv1
5PklhHDv/zuolff1nVpjf+CMta0s0TUELRiXFJxw/npDkSzHhcPKwfSAQiRo
mUWmKVhKubmQOWzuWH9Ma9oUhDzp/DgohHWXSggBFJzr5t937Yrj3a92OwCW
UZrrjv/pDP4p3LF7/UO2t1GFEyyjmjsD4sfwsostTfCcl3bFKp/UF8Qbji2s
JB0xK4X4zb+6gEvaNxuVsykGh8zkojB5H2SDCecjwI7ct5RS03trEFhWZcMj
n+zskHso5VZADGQ9gBBJmttCyTuBgy0pcB4WpsnQS8kZRyXFCGiq7KAQHuvt
z6psPLFHNCPK1B5ib1RGC/mli+w7FEtpV19M/zPhn/skUAGIhT9yLCb1iKD2
mVK6+3b23tAsWpQuzlL5gORSxb0M+JfDI+1rf9++fVGn8own/FYFnpD9wmFT
mvI3uVXzZFt36pr+LmAiprUTkJy4h8d21HYHPS+POCVjise4lHP7HgrqUy/p
pPnX0QJU+ogUhGQTGJWkHJluLqYtT2GIcDCm0fwPWMHXxdgGnwsGTISib/Gv
xJkPCRujMHrxho8LyqPdIXw35X2tC44rFn9dYLsO3KCOCj6Y9AjzyrOrueo8
VHKEDlsvTj5en0cxbFzt3/KbNtsvU1ZWkswzg99bSeLz+Nnd6qBYJxTtIzB2
0CwEoQrRMlk+ssODqcg4kPu+0NMEb6qMsqYkbwjl5o24gSrUqLLeZPEB8V29
7MxtA/xSNdbYSlQjTjRO3LMJ9LUWmOLFrCMp7aHqUpqfhIkNY5HwS+kHt0VZ
DSo5wt+e351hZKDTsY/e9kGAd3RYt0TpGrVNNtJsa/52bRWEgKypf1vagUhq
ny9coGAcmbDG79SLSGAWjFx/GCArRt7GxRnhMGiG2LOatHq1qxkO64kKKhQ1
bgccmhO3FEOPP+yBzPwRjbH2OKA1MrjYnEJi2URD52ocyml7Kt/BmNJLOzSM
ZP76SWvXj/anvaT4oDFnlmtPP20fBzOPd8DdEw+W/z7zzl566m+hcm9cQJWi
omysETkSRxtGjKNss0lAtktlDy0wwWER90DaJuR06Zj4cp+SFTJGPTXmsc8k
lZ2l68abhHoQNiwjEIIgkME6xM0fgNK1GnpFwGL1zd+t4h6CfAqIpLAzofhC
TGGWWf0/+CS+iNDEB89kmsKN3hLocFeiXtRVD762fnCsptkPNZnh+akJiAK3
aWDeSs4cgCo4b08aHYRMz9Fi3yro8fPcy/ySaW4iRrJ6Ku5o+D/RoDkxxcTN
/2iL88ofUowV0WIRyE2QXGMFH0x6bgUJmZNZwCjmnESwDvLvslTsm27M16Uw
eIVo+ULfXK7jj5hiw8MWyyyqL3N+uEhJ34hdr0U84oSGdR4JWr49S4/foViX
hS8vTtTjoFNaETjoll+SJjruWTphb7zT8y0yR9b60AdspoeaST65tu5BO0oG
pnuWyNGaSY5EEQ+SzZnB6PX9f0jbsw/FFl7yMVzNgvzpUoId0mt26HuziX2X
dlHEoAh3AC3NJXXtrIld07bChnBxZOiUBWJ1SynaLF3ASsyacY+WRdCfVJlG
GkDtOZGwsRJvfqWrzSVl0OiXaofits9UxICqWLpet38Jqi2Rq70j46Z5QCoZ
vIE9AAH6yKg4Nps8brEDny/iC04x0n5oeaUMVhJ3ReD6Z+kQTk9wujaNKEk1
6+ePtrbVkga2ftmGxoU2M0xD76Am69gEYe1MXUqLCMtIgTUGUaakd2uyoErX
k6B+Q79DZpVeRyAfrvW6aKySnIFhBbKLQXoE3DMZjeoNPWpBx8wODtDzcACv
p7QkUk+Gy8okw0BLn+TzoOqwfbSLX44AVVzZXznG/Lp2DTc3aAgIxZFQTEig
AFcAs++p7UDi4bMrtTpDAec+Y5TXBRg9tYvM/C1fU73fHJTFZFrSPaAOP9+Q
9KJw3ATqekZT4ElZGPm81MaZKRqWQeqZmj1KVujdWDfSUQEexoip/R5lty9E
tqy/zzVyoT314CbtZqjWyf7yaxpgHAsf0Iwd8muG8QzyviaAHb1Rtr7nSQyJ
LKfFtAZTERwET76No/2csuavX8XTuYa9kKI/NIQerCQiNCg2qorbdAynX3lg
qmYbGhnTyi+buD+SjysO1uSE5Z2UXyzKBGgPCLgi7RnDJM+O41MhuCNuLAfH
waR/dHEJuS/9/pVhEKGYtFZRaF3BSLCl8cto22F5G/cRwMXf26QLZ/dvZ5Ug
wDdxpEQfGNu/dikegOlj3EWCA+HGADq6hBuTD9nmU8/vd62TE4jQ26q8YZxW
/5oTdLRMMwcKsLSexqwheHrpv7EfjLiaeTyOneM8tTN4X538cJhwV0oKuyBA
bvOkcgOBxHbeyEwppjox3WvXYTYbwaRGzQNnmCHXpm0xGzseSSkG/pUlxZyO
9CO7CZ6B+XrNj6QidL2tA61XKKPA9p5Bj6hN0lmUt3iKRGNRWeRuogCwZO1m
H6CEEB4B3xCs3Q7P+fIAGOgkHxyJZR9U6pmDcXb5paOIy/jT5+miVzmQC1Mg
pf/wZLaOpStzDMINLrjzRP5coot9tcyKVT+z9F6j++7On5tWnMEHNuHQfJKL
TQqsGZrAVLdHfCN8kvCtSpsPxfsv0gbFQLZB/ERrQRfdZ7ia7IynAL15Joz8
EW/4Z0O4eDi5eDEjK87cbKciq+Psv+Q6LMXpK9oW3vGNW3w6APBx+6ytTSKQ
DX0P8/bhTjsHgIk+oT7kPsz/CCnw0dwJMbRI9ax+TJR84nx+Qv0Fx21aj2Qo
2QtGRMkyPg1KHObxx1KukQWF52c/gjijvSB8JZ7o5fCqt9Ps0KJ5bR+OneTH
DUhp9ebhAk88LO61BKK7flcmPz9rCyzpQQZwvNzhikCONJveVP9LI9bQHPcB
THf3KLjujtIrlxlSkRlT8z7UOypW16i/WMRqvnSvyk6lQB5i43LmyZBL5ECy
z8x6UPpZY4fm0cM3mKhYqFn0ayAyAlZ5DJ3cy94fW5nuzEBVDm99F8JLvzVU
WaonrCykuaPJQ1aedd4ChJiA3DoNoDQNEmBpApA8oYibOpSlMtlgM0Cjy4/a
9CBREYprys8yEKn5nZCQCz36z7TwUYp9dFD9PCJfEPTE12ooNnY7P50gywiW
QvV8bAfbfctVH2pfyrBeIFprDi1pVjoW8phokTJ0jditu1vSs5fnXFdJFLUc
HT2LyNIjNpRS33ae5OoQom0+G/UbDeNiCGPbIQLoevk1Tb5tqTIJI2j5gRy2
goYwgi+YjmoaCrTGytEacHK15ANAc6xeWa67GEA6OxDE2StviBwfPMd/jHum
5p6529VdGgp2yPXBeSKxcOet3ogAy0VNTCrZl3YA7Rz2aWh44CJg5UavQYjN
UMaPodUfmKImZOtFr3GeQYu3Fdjxw1baMJjZWUkeaGWNv0gV34NbfZP5Mv7p
FZ8lCHKXks1XrBxugZ3fdrwQOhydoYFBuqO3gLR6iMKlEicmDEDMTZhsLoJ/
/gS5a+Otipo3DUF95kgc+a1UarLIZpzGBwP4qX04ylmHrg4QMFIz3XzAl6Pq
1oOjyMnj9LQ9lPXOYdA2zJDpxc8bksB5P6K/tduaPZCtQ8WEMdd/tQ3WTWqW
hsEc5n8cKl0K5SREmekWvj9m3+nLeQ5evBWd2KuuWc+tWgVGQcwS1UmL6CtH
JK9NCtIZT4ASgjKsre1FSiiu41M7x9S9mhlLJKYVnLJUYokfKS4cBqWbFHAB
UhIslmQ1CHwiaC6BzrU8o6tXKq4YFeAKWcFIINd1NSmbH1TrISPf8rVcD0BR
UXdA1XCOAqQSCas27aux6Fh843+oDdi+J/gjidSBNc3sbKNvvf9fOsq9AYVp
AbBmDuSZG78UbEPS7ji448C+28MrtkR8uhzdj63rDEfQhLJcm82ueKmQL5P1
nU5xa3fmmft0o5hqUp5OdtmfJsGOV7+nFFWxysoi+V3BYP074U9weI9ms522
x+C0cvAyd1pcalCm/Jy+RR6Hjp6e2HmccCuOIZ+k/LO/vBfHFeEGNguaczA0
/UpbhVp2TQ+kMbGNQQM4UAR/1vwQoqyb7jm2If7kxZG4SdIlASqarrChj9sa
/cDAzC/p9oA/nGa1VGLx1vsHE545ZXgVZgln

`pragma protect end_protected
