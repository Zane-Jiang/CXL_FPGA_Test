// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rmfUwWuyfYd1Pat8VZcqAmSh2yLt4xDXnAlCh/MjU0MnAWt10PWhvX6YOyfd
XVmpGTYJH7Ep7lPadhhC88v/oazV+tHEbG8J2Szfd1A0/cD6jd4OAKMiZeAS
elQ0VB/ZAD5Js0xIz+bDBjTuofpqbMO9r4L3/PThH+3OnCnrwssb9u47671J
xSVu913w44xkxdJT/vhlBns/zS0cp/q7CulfCMpNw1O9tXv9jzNJFAGlzW0M
x0w0b3W55HH7bOa6vB84747TQI6gU1ODphVkeQCmtyxSKATE4qasFQnkwF1f
/wOWmmIPrVx1JkuVO220gKdqeP4pow+a4wEN5kyvHw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qsR3GNkPg0Bgdur87H6XYdUAxuTCQQBLQd1DhxciPL7SIJO71FvMaMhHczkC
Y7nbQ5NOJd+/0nicHGgzEIWzwrDeGBNrhT+fTimzOStYiBzZugdnNrzWg6wc
ypFlEcTfG1miiUdwVU86FB8JzBQ2Di3WsvgEwuZ+Vyhq+H5H7MMU0OeOaRpk
kq98+j2eyT83lzQ3pbgpoqOJzMeiM3SZq/0MzxN1zwrncCMoeXiJ6tNijTKf
9TsveQAhMEf8H44HRPhcfuOyDweBByJOtRq3HmM1iuE/apeh+XfZ0zeFGtCw
Vb7wpOVuoDTwa0hP453KfJnPUiAFWe4d/AYbzKLBQw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Aw/Y4PxhzaCwTSiJS9pn/ocX6jeOkLtk2+FQ/s8i8yQm3YMnlWo5q4RJQoLK
XgeIwf5ssxPh6oKqAr4MDaB0eHyQXNtuNZpdZySUuHWq4sDZfRqqDsi/szZJ
0lvQr/LFZVcJdmRUruCU1kqPu0GdmqW5Akc0pywTOwe/BiPK7I8THXvQwdFr
+cEcRTYlelYQjgk9b4bZtOWDEh+GZVvSLIhjX88DzjcYTCZjoNR+4Nkjpnq+
ZT80WzuuAuNEPqKizRFMBbqvrJDsS9/RrG8nOcR08gwvRGLcbBlR9DEJ+kaz
4FoLEeJnEsZpA/q1Hq3ZX6yUkP3Npmm1XLW9cZUCOQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Enn2O9DWOytNKDrkGLNjITy5PJGtagsreTOGn+tQ22H/x2dtys6ztHf/925c
dkJM/P33Qs2vnIZn5k4kvbwj2wkl1az3/4U5geftRC9JDifl2FvxXk7rSC4+
S5dSQZhQOjrLYMMHMkVg/sMjKNKHjJXwG4X+JFlbXBmXX6H75b4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hC1HVhjuNhYtYRrFg0LChMxmeiYaW7PghE6HJCKEaYmQSyN024VNnxjCJyUP
Am8Y7HgNLkDXZq+nS+YWCKWsYqFMfElPiNTxYl4o/OdVdDB4Hit9QYnvCA1d
kMPE8ZJ+XcirQhQh5VCyF4BF3C71wlztoveQzBqzX9N9G1jFiF0ckD+dLO5Q
yi+vKo+XhUXipriKEgLRZ4sGPgz85ukjGrQ6lNA2NHIOh6wR5u4tu9xgPKhY
K0fQ8qTcqrjZE0Zww98PXx3d/aqMTfI21YB9Y+q+UpcGQFzRTEoXHoXq/iWf
yW2ZX+Gn/QWV60CZ8AuaItfBYfUQV3kU18sm7vKOQ6EYL2WqQ/bpn1fd9SQv
GObv2lnsihofY+1skNB8EQB4a/084JgQvPDePFOQRMiU6i0Bw+oPU40PFuyz
ZgdgD+JGyVTwDIZCFArjraF7XkxMEmPUoeQ4Cby1BcL6Pun+WwtZrs5KkFGI
ksV3dLt40d8zKEygXXv7iRjTW+F+TzuI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Htfu4Vseqm1wZW/d+xbwKCc+0F87qxOgFPUB8nyfGZXSxssCLzAYmLUnaQT1
WTks2HbbD0WOXuiJ4JVrcO3JLU5m+plA/chOLAhGjuZO0WjDO5WsLUJ8yJeL
EodraxLbO08Je1fiYIw5gXoEA/ZHsuFHp2SApdu1PERZ3iX9aYU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hp9gk877whY+G3PjwULxMGBN9oWV3lLTYgiVfFMXKaMfGV+yk/+2SfzU+dlz
mrciNsjQLIOPPeF7OsKD3kPs00kEWfJk4BmrFLKcXIhf1XFqxDffeuGaWZrk
4ypgglabaVHkkMnRYwDIGLMaTsN/uXQqAn0soRL1SgJ7uGzzcYc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14704)
`pragma protect data_block
CrKtPMcj45Nh8kYoZoOn/M67HHjZ8mpoBTraU90n7YLGWm5MmhDSQF1w7Qcp
7PRHEiXl5RqTrJJoSkLUtpNAD3teugepwKdmxqhrO1EU+7U2S5GFnxwdoBrT
h9I/m3tfAs8FNU7pejzDlsjdeO1SrNOHOSSZSvO4lrzYC+urrUXKZ3HBN34v
zkpPDfrsvmJivSB4Z/luKbWOuFVH6jFjn2whAcAdsTVFUjD1617FGLANxj/l
KB4gs6AFE6MXqjp0G8mZE1QfxNextkVUMnHIxUCOuo2p2d4AsnxFofh0t+yc
/8yqbR3kcbLaRi2QpvViRH8vDdvPhZdJrYmfNQ5OlMwjc8eznqImBGZ5QeoS
zhCMEA/PcFsqxfNXPfzX8cotKC2csGSMuqbiyo/uKeFRBHwsnY110Dt/vCqC
mWc2SsgUrvgylYTQ5mPGxuIiCS0nV3e3tDu8AtcS45dQzvtPw27q2nRUcA2N
i5E3ZGnxgaBwcmfkcJfpBl3sCVG6dJZ6TLmcdspsvlX/u/vuyN4aJuY67kLX
owTORJ8PDqS7CDciWXDAbShWJz504tez/6vqMnywbYxpc7eVlPFI40AFQ3V0
7byB14q/Xeg7KWDrS1XZp0ymf4ydBs1SUW+MbyGs27phwZm9KmH6gRVktvbg
k36Ax5ZWQo/ozNI467/W+/NlHGlxPcnOhYooOTbsU+PgV/Xps/ct9DaI7x2A
6iez+bplC9X+xpIDANbyTfsvxJB7X74VaYccn+N48WRDNjWnotYQklFDFh3+
T22CoVj6Lgjg0AIcw6Q+8m5cf/OecJEVc1h37b5xE7HuyKoXsk2AmRAAksor
lHZDr/B8FC8Z9ZTeAC9y8FHoYJcwcta2bJpGy7vN/F8XlQIgOhk0vhEuQEJv
7OIBxL9RzBuKEYdHBjaFQ7NP+N3loktf2hNTIlGrnCF3jc0tYuieBE/X9yHQ
mRaca3NwzrweSTljdYi9HUqhZIsBNGixO4T0C1reTqwd17AJaCsF22Jaxqqp
KzBhZrZ7DJ0SxK+Kd+kUuEQbu/vJDfwxzA1hV0Nuzdw/N+EVsJ7cLz8N19gv
Hvyz4ZlK9dGJ+djVIGu5caS+Uk17bp2Eyq/4julYcUcCZcP8nfDdC42CM7e8
5EgQCoOLcC0gK2q4XGIySXkw5QRw+JAcRKHj2eWGITTEhZNcsNtIsEHZ1jSU
4z3v9M1MRoB9QqqW5JIHlSgACvPfbQgXs5sH89HsBnZJPITUq6sP0c0WDmKQ
HNBE4hWtyZC+4TQ0vHXkzv4x3PFgEvlZaM+PyLu+4Kui1mukUqwjIm/3s02t
ged9CMyWpfr+u3Vf9Tyiu9hIAbPtOyxlJVeuFIfunwrVTua9F+4jfxvFK4nQ
bFWshP2Do8URnnTyIQ8VrGqQHJ0x76mS/7ScJWRdoydBUyrp48AS8a+dz1+q
Px+aSUwBTVMDP1mkQroVVCrhqIpv5ruY2eRjmASeGHsRk6ffSfABHFZ1Uyik
3TZdgDT75RsghW+wOGyerwx+Q9NBB/nmq6wJYPPg55dt32IcnyXx113kBCPh
ka+u2Hgb/L0dLNuJ2nHYxHnWwSFQidH3qoodjFCa8Vdmp9mvk9Gzg+JXn1yz
b+0jCJrwku0W73MK35+xOIpba2ZKsIbvq8esM0gJBuxv164BoHzoHarstxbV
ViIb2PO3NzwuORSuEfD0Rk1GgzDMbpGYvUxWynom6E8PeaIy1k0rqJhO4kHd
r/1jgcnr2pXo2j/wbPOuLWSTajhIKgaKxc10RXPljvX+6n3LVRu5MdZu0Aky
UjZOQhdVfMdNKJrZe+eize+YV+KGJy9tgJEK9c+Tg1IRwvUZmRpeOKYsOrHu
2bVmvmELf9aXPsFqycMHYijN0tyXduaXNJxDzbnBckxYM0c+2NBR42SRJf6f
j7onWx3h2sV59fyd/G0HIYLBFAXVxVToUPUpNWy9nFCuHt0T7rAJ9b5sPAzf
UY/QbwzXh6x8OgH58mhiIad3GhOih8ysDojQYNPFX+6v+m5H4lWkxuDulBYV
Y8O6s507zDs9VWBWZ5O+bL3kxBF/wiKaSMuk9U7q06ndOPZHXl7JCIrNUzSS
Jx2XLO7J2wlvc2C4herjLa9nJE4VT1qI72epvo5UGG3gZnX91ymoNEmlBvs5
TsB31r+9ktq1IVB7oPlE9TZ3Q/aknIMHEbdzAOof9xkhWEdSdy0WpRu1Ytnb
3y+wENAJ0vO/rR+/yIW+hzeCtFcl/7877D51RviPp1O9i6wUtb6APPMXSC5B
dgDMMMy9Mtylso3fZ76PVEFnUbA94eZg/DSZKofPmiqFgT90lNJ+gQmgZ4/U
LgdPPmBaZALBjvLO/iD2DbKgjDNwCIwFj57vCN9Qu5odZQmSOAbLv8QUlX1T
VYGnea0zEiVN0YoLiKVMUPVNKbm4+MycEgIR8pQ7MuBzbpCYiiMXzzfStaB4
I2kC7TR8qflsHeVsRWqGB7UKzWZbCxzhcDVQMfMJqXroFTTbkKYx+NP7lBDv
kpTIbpWvudCKVmYYbgHsNdBP1F9jf/pXI9Kn0q+vc0OwORZ+Am3VLWvW442i
9AsX6qMDg5xrz3Rp8M9qMs2tUzbMa+yt1wHM5xbj/eUyyi0pidlR0f2eIkmn
3ifI/m7oNol1tLUr86P3+x1TQSzIzEse60w/N3BHr7uzmc5LVDkzxAWLwEPw
lAoHd01bE42ui7Ywxe/axsEB4r3pCRGwA0nSOG1adI8V5pRHK7zHERPPi+A6
2AkR1i6YUZ7ie/+YSdEPxtH+ijWeZKzDYj97OM28zytdQ/cM+CdHJu0bG2L+
NR5vK6751NlVa0rHHPtv8TW1/cpD47cjedQ3ZlALX7wti2A63Xmud9/IBobH
1Rfs1L3HyQGBTD1raKCMizhPUci03tBAU4/WKiTTbkN7+8W0ZhICwvvq2UmB
xxM5Nq8gYUn3fc+1hK1uPRDjPNOPOPcbKp/Djg8lzmp5z0hdQEujxJa3V74w
J0Fsum/X4AEtmuwVgd7h+JawRNeR4aNi/dv0LkXdExdUkYF+GWf6iTiPe4V9
Yop7SfJ81QYqKAMXyz4huCrGbcZ2WDeCjJC8txctZVMnOp9LkbJPLZeLpEfT
hn/OgZPZoNr4Mg5ZipeRzWglXr/7CNLYWnIVJdw08qYs160+8Xj83ACOftJT
3D7nJsrDpu1WLEbE1L2+1YeG74FcNAZi2CEV5mB3GE3fOgQPWx0mV134YcPM
5qJfsLL6JB1XOnXEt/J7oSGdaYmzVQhUdsiiJK7OXuOjQ8tw/zhoa2sb8AAa
1L51i0q+3tclw5+9HBnN6lPEhTd9vpZ/Nf5vUQllodPBmwWQW8JtvLofpbqQ
BHezSKOKDRgI5zOemNLEpIzW4GBbc8cHNTFvMzPs3Z6YiTJT/+zxJuOgu01R
kqi9b0ib87b4IfkaJwSkf0Okkqse+3/dmEttRY0O9rsD/HfxRZR8BSHP6zPq
kZG1jMZlgS5uKNbKudq6ptNydPCZ8wz4q8miX8H66UbE9GsjFbTz6LWLp0zD
gtjrl0LmrZqbSsVr70Q/s3dyBTJ0vGYYil2xGiTB0HMwMCDpPGksyeR7TLZ0
+7mJXWh2eWtHhan6fRLIx9qojiMq874rbBbN8wV5GM3a1k/srfgkCV30DdNl
TymRB+RDn03aVa64mC00QY7TCirAlIZLY1XX0LPrn2Nm5E65p+sSq7mdWiIS
+a4a2Mu0QTR/OmXnYchPk0n+WZTK0Hhf2z1wJq9YtVHTv15orA5r0a4UTD+1
8U9n5MHmCLU1hvNEisZU7jXxtlkNtjvB4VcedFXRFlhu+RAjFj3Uw5FVcKdb
nCmkHUI2oFLaiB3MCnPNs4J6IGpMtn6b31p35KNBLvdccYjCGTlHb8Yx/XME
4mQ2qHGNse/FmeQNhz57DR2ZWmOFzUWhGyVMPFctqVJh2RNjRYPUu2bCvl18
h3tK9y1or59ShRujuVNci5G2ub5xVDD+eWEcYJNEDsiLvYjSF/nFzBH2/rbv
zsC0IeIJ3qTLnFL06gj5aCnb5g44x5BRXdC1yIo8GC9flzWw1OrNWXzIyk4R
3aYe5eQzxFFadkZAgrrW1T7vhXfIha6Z6VH08Pr9TU0ATLH+AFrA2i4q4rFw
t6eNfN3jjbbr3/dx03VNZUYCtrCX40RV7kK9pdabmexJsT4GNtZhHf/6ujZ5
3CBiSz6TEDr2CFJESleNkhMD+VvdHJQyKuL7gUCJk3Gd3ynAbEXyO9SQ62ON
Qn46/rDsIh/TshKCVn8RmHJEPXby8fqEGEXaqHwd0T+yB+L1zn+qd5Wo8uJL
UgTc4DuM2+OvWzXDvj6D8+qOdoMOQtm0Sjqq7ZJU+hBJLIUHjtkvsedUbfnI
l9aVfM/9JyExJVyOd0ftikC+jGSKB3PIQlfRggnB1F9SggaCwNJzQ7TRWxBF
Goy7oQKw4SbAkehvGLZjjxcp5wOauWng6fhBvAXCGr1vFLZtocMW2W6AOGxL
1RU8b/ln+Y/SrEr2Jeu0tYA8cLPLndrmgPuvdlLxSlxIkce9LCMeK9C88Ewo
659T7H1G+7DQcQHIxNBnrpTWz69OeQbnsCuB5As6hWk6nLksAQYKUUxOTtBs
vKJLIQEgtCIPUzHAu2Se0pFo9ld7n18b5sveWNfkhW72rOnakgAkS0Tew0Th
W60Sxqc9eZQiLU4hTwXr8m25pC5ccF7KFIx/YPGKsjFMtWYpeya18KnT4vmV
sq1pORQ7CWrnrKWNXKKAEluyARSMg/D0Ytm1yeA4+h8gn8YD5Kklahfdqm5C
IX3yVQWSJsk2Qe0RRkoS2F5O3yRJ/Rb8k8iRK56VZyr6k0W/bcH0UghhvQWR
8BH/3pm+9gwH6JrkgHSKHBS2gAyzZxEyIsJLkRTxmPYx/AUdnqEfUGfKmyf2
vTl3VMSII66A3WMzRJtXH+2QldF3CXhwJvUoqW6FpJW4GFCtcuhGwWKgfhJe
j9zMkvoVTHLqzfNHsZPcArfsbOwmSPHlN3LWDZicqaBsy1N1XZuDm4p6bGrn
PpkDvbhy2uVRVkWQKJBQWkv102CYDjP3RUg4LFyuMFm8SG5bIJjNQDxa0K/2
PDKJ0I3pXseFo6WooJn7XnsVxhyKp3WlcPiqexW9AKQ/vZ+LX1JlJ//5bg7g
d5y0uviqQZZTUsZVidY7C7nvTYXIBMIYJipt9ol4dqJyUnSh4K1UCCUxkrms
sYfqsWpc6cAWtJGNRdjou9WgygHshwyY3r+HP1+mkTplfRqsWWnWuGAVJt9U
B1ajnhvKdinwfXYELZMWXkPK28Ffl+sdSZTAhKFcj3Ab+MmBHpkU5cQtk77T
o9k0+f1l7QOLdyXQDOT3S+v79E7e9niNj0vsFrfYZeR6oNy/jDanIwmg9XDN
hIZIO4mx+bpRobjGMneMrQzSX5w6+TOETTTJ9Whu3zQrGomAI6KLXlWT1QAQ
wZXFHnVzSBStdqzjiAlsgWaT5vdIm8xwg8xj9GIkWwE9kNgD1h1GbsTzuJ/r
rdL365xAL64bG/KotHafRNIGKLqgbg9pJtTZgv2CrHuVPaethOOgidgn6YgC
L4e/YPFeq0oFsdV0VFSltB/YAIMqV2QAk820Fq8l+K/OwDhTMSqxWeCrTnpK
cPe4mmjNLHnc4F/DlATfmPKK+ApaoPnO8OWsjLgnSHrqmbO07bkTRX/mW6/V
Up728GjcEYWUZYlOl0E0MIypbIG7PZNJiFKBn2c/GAkJcjLKZ9VY3n9Hg6TX
DkNhlAVHN9ihDVZytBAW7c99Ij1AKWLyja976xC7GXuRgQxMisNRKh6ZReAR
/F37GlGp/Sp4IjOxsRqTFtfLAS31exbg88d+Anh9RFSOGU8SlhIs6efU+q7x
wi1Fug0nmZMOOFEYxg5PgSZedgPYqaAbgii4z9Pc64UoLa9BD1uclKD+uJBC
tQ7pSHWAkZvhhfFZMbXdBbGLcwjeUtXYI2lActyHCuPrQP6v3cugzmrJygS8
T2arbh7Yh0aGzgpkKL98tPyldKA/dsBbM12AEyVZVpRc7Uxo3VvnnasloRDO
6fgYU6bWOTAHMNyngI6XkS23enihkof9eVR3PEsQospUQL0l23MMU9JwJ7qD
6hYQiu3/GUzHn9tjaqir3XwOA/rKVEU4V5RDed8uQ76UOGns61+aCGLkzKli
3qx8vcV7ZXp8ql4JFZqweeUPVOzvBZy4WlkT1cd/2NbtufftXIUr9Y8y58zX
ImhBiQ3qGgLhpih0tfchOxycRg40bhuyKkiUNhJDY5xkdGjY9fj3ytttiQgv
OLrV8Bkoevm23stPZOPzjw1x3dQ45OOuTzFB59dOuxwkQffJqTRExYUzSC8y
lHosckIT5BL43sLa1gyJfYrpogsaG8XTXUR0a5kZl6VZg49Jn7J0YwcQVpor
GW+j44YkQBf3w2FpjPl/ydE2lgRVVaJWTrRSYBic93KmhrH4eO95L8NVP5cB
J6WAaKQRd7ml1ACOExArqe4A5hZuZ9f13/MBT7YaAzjd6o+xskIWm7j2xIWf
fil2vTMvfH1FqfrHgOMHtojlWo/nwoYGc3tAydZ2HwZwIiMd4lHiKU8IXIgX
YXKFfM9KY9kuwpxpKdU16cNqrJM9dIBZRBS6Wz2L+uw87ZSYJCt+qf6mDZ9I
NpieM+y6HX2O50pLwMEgNiny3tSW94wVPJYAphxmpe1DfSmZdp+t1EoSZbr2
y9lE6kdpeGa80bTtqT/Y7I7CjhuyhiwJUsyTcNoPqNzoPvWZz2L4wW1RXMrJ
pmcXnZLoSTCoLa/e9KegGq5/vIPiKJKNzCaJ1ptOp7af90kXhg4b6O+D4XP/
tVX8qnP1yIBu6ZiNB9zZTjh2F+7lpWcqGH1avBTBhS0rQsIophQGC6tv+rlC
eNTR/rUPfRGJZPN6Zzs9AWn432N4s3SQIRYHYZTx0UJx+KJ4mGrM6z1aMOWc
lhxIVTuwnpnTTjoIfEJVHpG7UwV4rJ3dTPFi3Vj+z2sH9nd+v5Ufmie3eClZ
gDdOBQmAeVSay4EwaiPWNmg9AonqVFctRI7CRrP+D/3Ga2vHIXlxXKmDxZQJ
L9+ztZkMhO3Nmkk0+0nWt8jI70oI2GB+zMhXHwPNDpY0ZtH3FagLB3z4WFmf
YD1wDaub2Xyxo8nnIjmF0HZ7FMLXcbSDFlGkcMnaWG8aQV23Sx4XHIdRUQzC
fawoUvgSzB1RCrjTfTSsxaonxH4/67HOnHlVDEuSVecbb8XmOxQ26HSI47YH
7+YqOsm8IdUPxco7LLPUCNV173p31yAUQACu2mx2eHIMRM689+x5c7PyCa11
XneH7X49xSOhvYyOpGHrsdVD2S/a4X6LDPSXTebWIsWN8Krq+sm6FMdWiu1r
N/xzaMgBLUz7a4Fdhbh79MLFyBuvXxR/Nma16nDgjqbvayN69H6T4fWVtxSF
//hzENq43LunPbUEx00V4EvQqpvvUdovRhT/NF9Gq5TjXRTGok8lvfBV/dtl
mjqWUounz7jVBEYYZGntNHGGA1W54gMgFahpBD5Y10yN6ZTHIdavNPBQV2P9
Jkp2m2+zPd9k1QI9cmRK7nxhBvMP+E5cf5SMLr6QsSlJcBQ+WTnhRW34X8Jr
YR2MjiVzAzN6E5RbqCFD9IkCKUIQ1VA8YZvo2FfT23bmDFIfY5X5CD8ODtvv
19PBebAIVpEwWvSww96VfPp2K67jiL0hcLBfRQcY0nT6M1bzKZmFLe6gDX2A
1bdRjIRGPf4wse2PqiV0RwruXy5G/+VLG9co4SZQw3KmzNxhuxjCuYuSZr2q
qjHQyHayFb8+8RmW2d5i4+1qOijrG1LTEfu+ENQ+sRy//3FQ5IhNhh7pd9jB
FyFNi9tk513zkRZ1ztVebFHa/+3V/Eq7QA3L1KP2V5/a4n7W1cacZ4G3fXaG
FupS4eJLNPtTdVBhOcKHtMXDQXIpszU1BuAgUP//EhHLS1PiODwAlJot7TEf
iMg26NrIxXiIGOk0k40A4yXfM2oAfpIgnXuvWcxTsp6PphrOw+wP9fj572xM
CUo+q1Lc3Y5W3u4RplLBfJ566gzSJkv+/yycjcv18+mLY4kkFvcDQE3x+WO5
XEaXTjGV32BBiY43MJfOpKm+JED/BVz3hcgbllN0UkOemefdMZAbhERCDArO
rHlI531dGC/5LdOa1C8eEsPe5xi2wezEOG5KTlPwN657ipmVCSxGdPQZoHnV
T8Mt4bXjIQkU/kPOSQwZAZE/0rMS5xwdm07x1ix1df8qEURuN50/cgOGEIBw
kld7uVU72KNRMafXmOj15aPgNGnVDYUwmYyBo6GwocnUZk0BXjtJ96qdAdMw
atvprd0HO9qkT0xvxChT/jAS+4WLWebTdISwHg5EByv+Y/UPLvc4eCh3s/UC
9Uc7l5gk69eXgVbB8Wp7OW77wqYWgn1M8e3LBhON2lK4UptaNlxWiuLu0zNv
Ec8IGcMSmpO0rWDiOA/nyTW509Newm7067tsp00ETjLrMvRhr5aVEHq1ODfZ
hi0Lzl/khp73mkDYsQVC90BvkAPoTz6vuaa4fDsnAmhXzaAaMSc/uWFn1LYa
IFTwKFr9a214NUBWyZ58RXpYnp5KfO6jqANUuytBx0+66s/0bS/QDlp3lYEF
INBn/Gm6+DZRLlnXlShVty6WFa9eXkXpnFfpBOVr6aq9sbjw605n3NYTT9yr
Bxw2p1ArPAAcl3zRzrT6n+BF4wGm7xbr7i2lGWtiMuJC2uRUS4EiJSKDPzh6
GpYnR+JEcxnAgbFzB+cuMKqBiK5afm1fQmDa7CMZ2vqoIVNo1qA+NDu0db9D
qRLYQxK+5rmJIUtPK1L3YCiaaCbCwDYXU1MRuj+vOldd5yt/ztNKbheu/Oy7
7If/7mJtBSZZmtHLg9gHZtwzZrgDacWOb4n3nca9q1koXFEyMAIBF6gjfcLd
Glt7zb20FGaVZgyKB5Eb+6Fc3KVE04IKr/rRiJtBvq7USrP2GPmsma9VDL9A
HHD4pxj5WsK+FE4sRbVtsmnrvLeH9/pvqPGben9HN7vhlmTkjaOL7xxqSkTh
7V13YEIjgCCo9unQ+nZiGJIds2xQAJKRJCQhrBWCzhkNpANS3Nk8QvAeOvnn
OSvyZCQw9rB+rcY5+0xIxQxuMJgHetlYMgjs1gtgIKWxX24f1fvYqNAZWSTR
l6H3DkslChgE2NTskl0ao7Qtui9VdJP/7uOIRNaMV/FX6xAYPP67Lp7/Auny
irV2n8spFEBnASK8m6OvBv8mOwsCs+64SYEkB/zOAyhvFGfnDEGQWZKezjB8
/jfSMKbCPuDjMwPAHOVGhgy1lODmewLegJzAes060srBlwAZAy86UKFpnjlI
kNgAWDoDnOue5zHGvRnuMI6JVNy8mXCc8kOMWeiJntTfpe53bqDiPpCILsWI
/0LlzgHmOcGeHfJb0hTG4BtwoyBiAnqbtbLEascERkJNitrkkWqKXQkd3iyk
J4Hc5Se+/HFZd4ESsVCiD830EdayIxXGZt82vAAYHeo4xBi7AmeqDQh685rZ
oNGYk5QNNQDOCG25j2xPsMP6V3d6etnZLypWjHFakcJTVFK4IVWRAyAfTb+5
Fhuljin8TWtuqwDeuIEcGMK1TEcS8odwsnt88srhuxXmB/SuKF3XFIX9xztE
eMG+kj/fw5ALRhbjGdC6VVVX37l9idFVCGJDXR05Xw9ZeSizoS9/L+NCyByJ
XGIV6/ZXZ+BTV0lTvpVawS7yFS2e93B9T4X/aVfDXi7kbiuvhOXm+Y6KcevC
cHsLP2riwU8PtKb+T/xEyrHpZLjYM3P7YF9JiL3f8K+1XWKnVjhvqsYJ+Cnz
GtxE43WoXEbxL67nEh6C9dga8NgUGGuOY+vQM+Y8uqQlxyVHqs3RCDHQrcWk
vvp5cPCeUdUTJn/+e132wd5U3gbeZeeTpW8VjR9o2ECIqRIGntTy9niymoH3
i3kZymycgVzuoyOkZLRCjbZbXcCN1NMa0RA/i8tU5n8DgvI7ElBWSV6s9wAg
QzBsj2roe0TQ0nkJ9cX0wBn7uho5zaphMqHP8syDRMgmphykc4XXSBar4lCh
SZxBGrmsbLFljMy/jr59bM6tpHrWNmTsa4p8baqhO6crfeXAqOOyCecz9te9
mD2uwdF1m7mtx9MJBkUNE/hr0yhm+7+MkLqSUkGf0gdoqduRG57bQQU6qxPh
IY9SFLC7xAKvvug/pbpaQAUGdehCjwHyGzFULJdsQUqMZWHZKmt0CrrlnDfX
psQtautWaaWymRcGH8h+5PKuL/sYj73tzWS/Fm49hX5MWoqERSRefQ0dxB6G
cMBlF2+kRkP7+Bv1mKqnkGYiecSI0aIbsf+3DCrt4KnbfEXO8yWi+rC8XW9i
qblcFSGwJfDrbSzw1stm0FJCTnmfJlOp3GF6aTHPQIR1Fdv+FYAy9g9ZleRV
AMdAaRQPrEwzdSzdH3qXxMU84SMwAOoHVZTsQtm9SVKUOo1piUmRex/ygymG
Y0K+jahuJMJrKE+mm1GPezVuJHGll7ZI2wr3K9us8lp5qgeB2oH1RJsTK+Sl
he6gtOB1OMFdYvw2RLhPyJmXoAqsU1TGJitHPwInQbaHeYrCJoRSOe4Phzlu
XiIsJ9E4tFcNux3BC9BVzM4/SRcQfDVyVqvnqZlOxMvhxVnA2XUoNuQKggGe
t6NxxrFC+TmRqCYcm5ElmhP/DXmqmO87WjTriAq90fS4YhulQMH5Qxbms/fN
ctxZR720P4o106U8iH0GWgTTuB12ZAK8wVhMDRaN8w2Hk4N9CNdvZ1QPZj6a
FBpiOdziwVVdYSArtoWwaSlLJIWdXjzxgz06fVzp55i+5m837TFYeDZqwukZ
qiF4BzGWsg4nPwFSfo+IxYSAOUeakO7BfSZoSPFQf0fLtOq7Q6OpX2fA5W9L
t6jIMz471WD6BSHjmk9827Lne1+dehG0gNfgv3uFeZg4ViUIVjUrk93Vw+T3
lsoyxAELZu7HTeneAaMqNndVfHjRGIkwsfl8elAM4To7EWtZg4FvQSaFemkq
0H/uTKycIZaOwJe/e1/L/qorfdoyn664RSn6X6Txnrq/2W3hhtmWVZn4cUgY
9YaqzMtRBr3eqwq+HqyiXhew3sgI7bT605soGuv37qk/7gHwlXQIblr7Xf0e
TwJKnmOHCaVeI6eGOQCbKoTnt8DxInpXEIrAHQ2p3qhO4qdk7Wrs7aMVr/Db
iUz1UqmXQ/Uw/JPb4B4TZrOD51gGVbJj4mXUCTha7X4ncg497mfLEBJi2SoS
L3jmwJJhH8stVtikd6Y8RrA8r0T9FaG6sVELW7UoRY6+M4u7r4N5QeKnyyqw
LJW2m1lYabDFCOOz/A2+NVgNtal9L8qMPYTXeOB7/nGUkNqZtP4gOP+7hKPQ
S4b20S6wquoO4GU7TdSlN+Gi5ZlMOblPsRyPy7+tLrpLo1onS+fkiKm81Hin
qNjPSwB3u/Tm4n8pwNPYofXWtJ9juUvxJ9RkdDhnCK90IjvyyR2TuffQWqde
F47Cok8uX7p/GT+SrgkTLATWYD148lT5pWQcdSXpP4220j7ONGlgfTnUgXYd
o8ZjEI/w0emVgLalBZnER5I/XcR7lLbNw6RALReWG+2ZLkzhWm48/wg+RKPG
nrAEykQD9ZAeNuJD5sm/BJ8nkDk4ABM4c3U8jFVI35fdz122eSToeio0ToH5
KsgP3lYAs52jDd3MwD7I1XWAYIQj8a1GNmdMBQMTxERHA6xtv5j57ovqHXnC
33xm5GeLZ28U9Wzbe+bBbO2LmO3DVAp0vuCr3r4R1W4DnCUA5VTs4uDJI3/m
CoEvZT1G0HRV1EWaI6XdnmHkVSrl/dWG2bf4nhFqinp08I0gisMBNHec0Ee3
3pMw0FP87Zd0osbxFGFvSeVis7nA1wjF0+yR0Cmc3dwqrutXnxJL74Cm3x41
hREnRnbeBHlMwPE6pBydFnb4oxL6Bxu+/LNiWX4fja7aJ1brR/UErUf/w9Ed
+lAcmJBhAqk1y7nXKw7SYKa9WRdbLD0vqPaumydni9WlD/liTMKFmBLhRlii
K/z5Rvw+uv5IfjAKaKBFY4UPgIw0V3OJPvjMKMRSBxsS1NEDVCYP/GhopMvw
6d+XM8sLdf+PUEvPosA1Q4xsNYEHMInXhMoDb4VTqxRgomJl9FAmipdutI9C
43q03Xsr2VXVP2txzvEkI1744AXHwyzkYtwTjKmGH2THIyaKeGvdNOMezgfA
8e9AkifNnewpWaT4oh7WHq6Zyz9+jugVkECG6e2rijQO11gyJrui/L/JTxaw
ab/7F9F6r6JtXg3HNgrhOz0occo7aNcY1KrXYF18fneO0QbpGz3Fa+dAW/k6
6o49Sr81eI4T9BSna7uNL7oSUEIY8qhFdOhd06I5EKrkDXhQjtSEhkrP4O5r
emF80G2olSuul6WrN8ARGbKaraQjL/Km3dtRxN6Oxkf5rOFfjvz/JNqkuMYC
2IRY3i41bv3iyuTeErha4ZSdnyY+hcMFEm0Dna5sqB/4lmbyV0koBWugJsuQ
nuPYQN/W9D7s/oyBfT4dE9cuu0WiFyDijEeDTC6rmLy20IMI/leRMxabFU6a
CUoZAMibjW4NbSWaEoma6JnkuOOWwN1yqCA+oc+tzfy3PmUBdKrOTQ4fDunH
P7WY6QcDb4aApgwvS007s/zADJQSfdhcUCfEuZrpWRaqK3GfRaJfXs6ZcxZA
eX9hIrzH3+59rzaxVM1NH1FtvNIAIxj/DXVjJr+L1bSus3Zxf1yiun4LnBvA
ukBHx4cm1ltHY+hV9gj89WrhHOEUR0nlpvXwZGKvbbXzjHiQ9F6UYsP5hHLZ
aWdioljK2sElV+XqmKR+dkwbfoTf3OYSuEtvx1BDHkbzZZ/4IUv9MRQ0naFY
r94yrSuO+nQJ1mm81obCr2THkjxoq4X6zYDBknv082L+Ynvp/2rTNuOGpPwR
TQHzxZ4fQZ8N30z2r38PBe1yXTyiB6yHukT0+86L1Dm6HTlFafJm2/VuVywh
/EHmb69YEftokb6ceJNAcCGI3y1C30AZ7HdFCxk4YCMmAad8kQpF4Dap/ss3
7zohntrQIL977vMXhFld+tVfSbg3tmOF4uvF8sv+p/xFRKXjJYvWnUIMCUEe
wRKqMvn9bxVpRp3GEjQOdJW3Wt862k6X4yD/7u4zFLg0wI4Z5g295cjIGnW4
mO89SmYnrwZbviQnZk84+9upi7hDwEAubCY8djdC3dvN5/zwS1Exy47Fkrsh
NDxY9rCxdEN06i9X855Pl72znoE0M0+5e6wwFylnL01TjASKA9s1uIpk83pv
H3kJXKrgJ2jBJRwZXxPcxKFTtP+pfpoe6XRUWURt6nAyR3HuiK1PWMg5gx+y
BMS71cX81MB/zbxt+qDfoFDrcLOLlySlr//+MMCx0MsLZqASS6uGsxM5W971
/EmpZeonLQNiAeVGcJpSR0s4btKj70x7+orjHWnnexrb10FsE+j6SNAQDUn0
eW1yTw/eLr9TOKTbPQ9rEM+nuHhU+2tWM0kcdmcRKKvJH/0A6XPjkCjTi4w3
PJtP6xmb8TalGBLpiebPZiYmk8UgiLDehWxmVusIUmJovi7xsMj5ZIV9pQCe
LAh1nYr1H+z4y19l9hn98ETstqBn2AsZFUS6KgzRFropun/WHsLBeALueOBF
+WB1s3SRimJ7FOY9kYWYH7fZJ4y5jIePTl/wgTPctpy52pOydyiFaNaoGXsc
Uvnp6efSA2Fmlsb5YoQo3bYKLYmLy3BkSy9YtK5nrAf8E14L1PQsH/7syANR
7FB8yUoOZIHwbPCwKq7CkpkmRxofUzlXs7JVJGOoSa5FC4dbzQ1yJY1xeXBg
+pIM0nMfUClMNb30ia8FV0mwdscHpE0XKA9E5K/eItm+MOf3MSVhysh3EqGY
k5OlHLhxsGau5olHuU3zqkvTpZVncTKfbC8VGq5sYS12nW0dqIsoQvslP9zf
Tm4aEXh0DV90l45RuqHW9HWg6ZMgccuI9rqk915HhCAjpujjtk23RTad6IUZ
5sMbHGrjol3+onBj8JFGD9pjrZ1VUywMvONzNoVNJWbcdtOFY3eowgYRoyLv
VZHCkVzk6z48QtvrCahBwA+ysQ4KTZcVwQGAaC8lbwGM0T//vQX0UOo01cw8
23AzxcMqkNnoRA0rpMdbSPE2iYagV1Egc3J1yWYj12S0VeKVSNBs4vcOlk/D
0gwS9dRTNypjESByJo/77NDYm8xmX5fMSnhW8GEMf0Ct9EDZtnBOQ0R4SDl/
l108LYXkz9eSIo+fGzVUrpcCkkIWy74YvhXFUAO9TjAk9urD6hSxAinknw8B
oUmuMVLVCwAKIbTYmXBz4KnjmWYx6CP3VPNQ0J/CgRaG1436BD7+5+OIVP96
NJ2YPcxlO32XryNWebG4LgESby0W9PYBH0m+r/oTqu/uMR6alXLHdiu2j/4b
mIYhzxmd609I4XgMW5OZomC9dYO4Xh85z1D4MSdWmA/j8D6FQnuS284EJZvC
UFCctXWtAQucaRUVd+KkhpJhIgwYz46nvmBAdz+cHk9SmoIkhjkjM9ANKmTO
t2fYdRiyrx5eVSAF6KPGZnDMofs1NOVjjx4XKMu59ykw5Eb9MDUPBF9C2YU4
/bXViJIa83t6wm4c3RCb6jIQqgazWIc9GesDVMRt4qhtLtlxgntrGAv5virM
mISLER16VYkn4Nl+4DATWI/K7w04thR/gHGASmc2O6UHSOTp0wSGVjFoRtZ8
INbdBLZvoNWYd9QMkHZ3FMnD7+Cu9+5PTbIQs58eSz7urg7iVPUlwYNghlgH
QZq74NahsKIKk0NfVDaIEmQ6fwoup9nLozNVXiFHAfW35iME7roBaN5bkAkG
uyaXIGiFXzRk6yIlG6HVMeMYgvJhw2rFsHJ5deQ6Zlg2dOiECS118k7HiT4k
x4j7fgYiZk5n7HyFOux4GPxP56HXU+YqBIhtwBL2jvOaSqa5xjcns41E19G2
rI+wQq2NG9IdJtKn2JgpB6AoHZo/vmkwefPcdvhGmv2LMptbCVzO6z0Zg1vm
nUZ7JPJaDr1RJVUQleWU7Q69E6k+B4Vz5aHK+GuyvGBckxh2T8ElrbQqKFAt
vopmVuJ7jqTe/2J6vEtyeCOTkShVtQ0MR4AC5HMUd0hs8IPEE/ZSfQvuIT9v
GunEzirZ9rpI9jfmFJXGGIeU3QkHHBa8bwLTiu7mQbElsz2xrbOEFy4KhLlc
u4m1tnwmxpURf4WBvPig0njObZVnv9pQhUehAbf5Cmz7SoaeV9AxXxPSLnNj
BdoFa07Mg+TvQFjb7QJnFnFR98Jdr5jt+FlYSO8xBL/3BtzeV8xsO2m4f0jC
rehZgM//6XCeGPON8nj9R7o+lzORcRctlNY8C9+8zlhWDo+1ZmfOMaxVvAh0
K4pJc37/7PK02Rru3aEf+4ZwassxUpcT+JobEo31VB0c8T8iqyhYzBzXyoi9
qYhRE5Whk6VWKWfrEo4nFNjZbaqJd0eDi7gHIfEaPk7cJx7V5GFeuDWAb96L
B+bLQjUb1fVYFiXiaUahmARFfFMg9IOIln+g1xnvvyAJXVHQ35yRM7qvt3qk
36z5C9AFrTEXaH1uJB6xfeCn73QXIxhggOcuYb5x4HaTE9d/8aZtQTi9mAIb
sBT7Luk9GeHeiuNSy7lwQ91ZephHCQ8eFslPKtKwGcoSXdR6ToaOjImtqciO
5/trEBmJiH41AkT817fLWUiD685Z2SzkjJ4BR+t5HsYX9ObRXaAHALomp0pH
Obk59dkEip+BALYhPU2sjffpofBsGvyGbmbSdYeqp510Yx3zzljLlIYEePgT
7D35fIGIrlETzoXh3i3Ddv3Spkd9928M275m2ImnmCYpYiamBgZcV47V9XTF
pKxTdSdIlIXM40a6+duMp8tBCOEEKNdHVsH9PVcejVGwZwBfcRJo7Y0MpQqE
K/XaUe/6/pWKSYpIurGRqdVxzG6nJ2OTsGavaFslNtKV3wcJNIi0sEvkm3JW
QATwdev19NOq8DYpSuPcaWpXTjiaFZC6TAXuWldygMMgYfE5iY8/soLPWOBT
sZyKQ2lEdsBQqYqlefnoXoDV8Vjr0ONFoRLxyhXlAjb/VWmpC6pVkT0Z6QgO
GKX6ENyJjmpxnzFR0IeT6HDPsV1WgHRgHnqhCv6SqDhZo7ynGSabaNy0vi0a
0rWYo+F0H4an0PvLKTWc2GgeiFXiBlyGyVzZ0aCrRiB8juke2jcy4AEYVDHN
/dXDBzg5kGPmwR8Yg3uQfZxNL20di9AnnfjVeN+9aHLV92+557rJIMo/minM
II+JPFKG9Dz9dmbBiOKgGNqNT4Pu0FeY52hy3JKwnIOJewc7UrEh1ix2olOS
OWdg4OIxEbmjNgRNdtGCW8UR5spf4w25+LWC/7KdMLD9Msag4BUVU+gWhioI
tNU+sbEasoNqrlSxbwmjKfWxSYKbVGqv+/6zCAwUeZmE2Ww4EKJQJRE8hzpM
XB91hz9zOkidfGmRw0yLbVDHhIGvJmcV66Ls6igBIYkpJcDVoc8xBpy6Q5Sd
PYJB+Z3zeizyHUeejJOcT3+NVkFO3TdByUmbP4urxd2UuLv8JdJrmMRUWz4B
reZlYU5N3Q15NFH7oRpyG9Vv1Ruc57Sv8Y6qs46EbX7TynWSU6lSFusJ0BXV
kL0Unm+oyGOSco4iyMNF2qukOSN5RCAPysOtpCQHWlGw6ZfOjxbCX8C0goId
fwr7kO2PrN1e4/A5U9AMvnvZgU7irgqVdF0LX/OB/2mKdJ/bGXFwP4p2ZHg9
9bYLoklWQIyh/VIzHusTX2lorMTWRhzpkauK4tYE0kW+I0q3VSICBgm5Bpqt
iN6MhQKZMPL8pdYX5KkjpxJ3h0wwWDVhkXPuAVw/K88TSyhcVsp3L1PCzjXn
4xvIVVNeLQ/oAxZZwAfkVrDRL/eIiFEBkDUCARHQh9nZFt62EY3i/M+QSKEc
s61s+kuX5/25/ICPzZVE9RsSWpHHQsXkcmzeQzfMXgEg1fktQA6t4+E27LLo
1hdIoFd9qT9CY7v4qVx69YZoniVOVUO+kMsDPUBjuKML1Y0/ndrco/lU0b72
xy+zGqIFW3txBlImBkvL6wDsA9+0o9LMHo/B6oK2E+AEBZEE8LIgmxxHGAbR
K4GusaT2WQulGZ1Jmat6udxJv1tQePwQnGNfJrP1Ve6psdwir8X8dYK7WeVU
3/xXd6qol7bNmU4MkeCE5mNJT2kTd7EPK8K0Vx1ySMC1DOBlK2tOLF3TnM9B
kJUwqMgndkpSmWkzMOMkbehRmF3oq1FTDYSFVj1lznb47tUGu/JWpSWmAAPH
fPR4LR+U4dDQp3Rdqdyq4xTXEV3ezHwev4ObdifompPuBJR7eoBm4wEDhU/t
nxDXh/XfqRocGWkPu1fGOLOuzN70wAlw5AEaEpX9q5QENX4/ck5zt+N1EPaW
fB1Efsy3Ue7JY4RPQRCqcvYAiSAnVkERczJJwS6IFe1HI0Pi6EkEkKmkst4A
8ySgVvU8JrNSn8taxHWYtzdUYIkzzcIOO7RQ10FxSS8/uA80SnuM5AuzoiHh
ie1wNm9FENoMKREz7ZmrjRykL8HzDKu6J09MZ8wXVJKhuwoxAOCmlLRGSbNo
d26x4iEU8hPiVuUTEHtWyXwZ/a9On8/itbOz9z7ziRnRPyDeq8QEoaTDpnhW
1gwUroECCwfw7qnoljxLcxRbzfrDgSnGBWpoNUlIyF7zgqAbrhcPtoEi55mx
EY3DcGN+L7bJD8SxAddnqP3okrvrddtRzN5QHi7ODjpQfWscujQahIHCHatm
Qgt8HUZb9z8t3hObWQlnGThZsdlOyorULPsD+3Y00/Jz7U5Urb2YfiGdyY1u
GsznGtpRGlcvZpxkrvcwvMVt25kCLZjYXnL3w1bwq2Qa3+8n8cdrd7U9yxNM
UQcL5nJTFNDkgZ0x6B2N5tjpT/0d/E1/dJgPji31tExT+XeSmiVz7yWCpJdE
NYvIyNXY7C7wTxtO5tUDbzYLvtTaAFfFcMHN0Xvejwg/VRgFGszYFWmaEgB2
UO0QzIwoxeEPhaqPbRu1cwu/PHgXN9GF5AyV4X8xQoo25Fsdo4r2o+fx60iP
rY0qoXPPBXDJLKfTWvu04JBcOiLqZsOYIu5N6ylpgKzC97VZM/4RB0G5ySvx
CV7yLm/gxE0MvLviOYIxnq83sgvTpgRik2pmL7x6Gc3um9IbK5oJYrrCWPxq
z3bBoMIhEIFgBkZLcl84T4+76FiwAXHb5hSZNpUUb6AUjNzeTOsFJXaPz5uT
1/Evjt81gIsZtN9d6FvrhVV06p6IVajjwf3goo3W+3F/KqK6uf4N2qRGrW5B
6ITKn0HgfL5cAKgA0DGDaIrrXXkkvQFJmngZpyLPex2SDr6tKvgSkG1kwb4R
bNRobtgXa7H8DJxkl5l4rh8ONVFaydjFVf16dKLqfHklgFykcexGJaqvsrci
pScVRNss3SjVboBegYhtjRXgg8on3rRVPbtN9mRiztZlj8fGw9JQqX9IQae2
A/QzOVNLAk/ao/A6N2cJg1ILctofZ8RsrjKBCBS0UZ0eQxXSu6Z3Cr94KwuU
ptQdngX97hK5BiCJ9Izc/xHM7JiMYS4K5x1s2F05PDmxxotzb+PgASaaJkIH
1BTFmPiRf+7YW+QE1fOiWXWNTnpMBGoxEvsvBY5yaoNiiYw3VxQ0tePvmUbE
KF7AhDdVQxrNnBJ1LFMYDXUVE+VXgFWeMsA7fkNdee1icULf7NN+F6OQKOn9
TMrGrsUmRlylbDYV1kdDUSBTORMs7ChUQOt5RCt2oJvNZMR2cSAC3ALPUx9D
qI9oQdeah+EY/UOOTcJgDqhfSAC2OY5BGKbp/7zHiUU/n0RiA15KLzVNjAlm
k1YFEgFl1ggs4qIt9rMYE0Izn9kHaTmpW/CeRHem2pogbjUWe2sjeDgwMsPT
iGKNDpvwZxc1zYvWIb90ZYdJoBVleXDUGfYSlZJah1tsSKn+wItYbDNHQRAV
TxHmJ4pL1j3IBSLWVyO61q7qjnfh1Yiguvaug89oSpL0Re8CY+/6jd1RpPQL
q3XkQ45Gs39dQgi1FwoEQFpkBb6Q+//fn3M8wtosEhxTG6uQAu7c0wENaEWk
S+8fgpAL/n17FJmyvrPm5rTrFlMiuoQCnj+7iginap/NVHB+qFuwJHz0OWWF
un67czdOAE8EYMJnWP2lzmTDtHmjcDpF2O1U527oNvMZYbp+lV8zNdd4TtHe
O2LgVhcieNn3aCCF4SGo5TE/CFwR5ux2eZ+qq1iKMLe7ykjDP2MThFK+gfZs
cX0BbSSROqkxxATNAUK6R4GguzM/DgWcWgdAwv5XWzHL4YXKF7cOw8ReRLfW
nlAOyGuWSkGJcthJZ8PpX6EoKgKffz52LvkEeDscXkq0du1X0nafW3v+hVZJ
O1RmCmEK3FFx1SZCCC21VDhkLGGdHtHf278iW4e3KAVtpll6Fb9OPxyceDQI
j4lUctz5e1tTCTtWWwvarxulvaLuYowkjHwo1Fbhk0IUIGSxxFxlGNjRE12m
XvSiH9SE+UdrDW/olgBZtxNrp9OAXRJSIC8KhQ6M1p3OAA==

`pragma protect end_protected
