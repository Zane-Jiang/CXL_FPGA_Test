`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
i+q2qNhbS0u+2n935h+/f8TZ2EIwf6WyoQ/jURwTpqAoCzcS8MxKHx4cgjkfz695
GxSXM99RHuqh9PbkHtNUYz7zpf4PDAQvanXlHDfOdhugNJAmjdiTSXhCe3gmhiZh
itX7uOv2z0TpBOQ4+EtfdD4GBnCJaHaAURghAJ6uvVo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 11216), data_block
ST8u5zWfT1j6Rp/hlt3G+it9hjbekO448zivbsPUp+ZEAuqqwkGuiFKhTU05a8ZL
3+2FTq+7EJdqC105f0D2lF41BHDXHn3w+W3yR4qDuXtCmJ+oENKI3ikiyEqPw2pB
uz4ajFLeaeyT46mbvJVDKDeiqutDf3M8PunwiSu65kx1iabSzqd6dX8JJ+XO06Xw
kEuzIRGLdUg/tks2eI0qBiupdkQIo0gKbGE+kCMw4/HpwNZR4jNPfB8H+pmWcpOv
IE20rKUKmUGqX/Y6q16CiEYEd9cvJbbgTjh7sLV7p4SHc8wdiDKwww7UWRn4EWkW
djLxhfjUP7VQV63pVzANRtZu+agnNU1h6nBQ4L+a5qYEnPc/sz7KOfOJiwbEkqXR
bLlW/u8fomtj1f8DqRQKNitUVeLAHTs7PS7qi2aWDpQ0LfPQmtr6eMbH1vfzgRG6
JerePtB19GlYcpb74Bkm6sXm+l30LR9FPKI6LcPZigG/Ec8FB7PTtMQXTrQxcjGv
fCrO9/Jw6G8UP0IL5iUoo5wHumXM+Mos7TJLBXbOI1hGzCqV/rpYH7ITeiNjGYc3
aNZJFysXd3Qv3cXx9Ewd2rPyFryxG7QxednkfDd7I+jpIu/pZIFfyCHQdbdbP+Jf
JWWO0A48/ILQLm1YymttrmmBhXPI8AcMLBzGIDDOtYumPnzgdTHidKaEjwGI+FWp
qp5ClSAOqDMM3kyPK4cNVxu/6dFLqEd+mJqaoG4GsiYd/ShTbY1kwr+aQ72NEYi6
lbRwW7l0qOZ3/3eI9ap1nLQ/rA/4Max6b5F6upCgOc6T97MoiGRUT7jB5sAC9uLm
iQRRhvnuaVzaovnCZPtXMj/UGgdnUc28mAKRe2FQzbWycslcRyLOgAO1fzmAyABE
An2fmXaDNlU3dUsc/RY3eUYtqBLFDV3h1lKj/QXHfGraQmh0qchC7IgIslLoHYHE
36nTBsjds/uEfAnQjne95BuwfvUUghzXuaZ3CtAn5yJ83UbX1CLgCbjvCD70lUro
VeOR6a1arvD4IKXciWhetGFqiGjVPQGeCRra+hzULHTlIY5/jHA6glax77HGIhDl
kiwEO/uF+RRzRp3uQEuw1CblU+aqAZhvSVk22nnLk3iPgV5iq5qMrrHn2FWHAjtK
VajgCO375fQQX2H0pQW2eb6a5NpwolcBcrMhxvnn8w/NZx5dSA0ONbS0C0DDE2zo
Lv0XZsqs0oW0Xvz9wGQTIw4J/DvoMLYEd6nJh70Fsc3z2s9pD64iPj36pHWNj/j7
QcYxXzg81lOVJiea4Gk19ggO1n1fUHPgbgSDa1Xag/NFUdSUjwvkAjmVehrUwekp
k3gu31M//MYqf9Tk/qsUU0i1j2vEsOUpwG3Iftknrvk/vrjF41nu+OZyzai5m4xZ
MMkQQJLU//2LeDCu5lqcVLfdX0O2yUUw3a4Ku4GU8DN15+USoIBWDIq4QDJtjCqz
uodKKSj7PkQPq7K9yd+IJzhbFVvQyjXgPXcoTBcpemtWUwOfJJM7lhIQm+C9Ocwk
kQM+loRCRGL8uZKpGwnsPdBCkVRmBLLsSUIR9z1GHO6QZqejB8xKtxq7r8bb8AAO
l4r/EZ5vNTKnjtd+7myzafdbyC/dNgoXQaJJ3BkwyfhS1buA6M2nrm6PiICmXuc6
DOQRlitkP44yLV59vkUwTjbHhXSdKx++cqi0SiWmy2O+1B4ygxOCbPnsSOecsd2h
8CyaWZi+nUluQTkWiI+9rPtZqxSPwPdDbBnWXFL74eYN2NeXXWucNZKQdFm5oIOv
cFQ5VybCPYHttR+K4MOOFs5TU5QtLGJNNdvqUUXuaAKvduk5byafvRf3g43+n36p
85+NhdZjHhibdObUrryAL1Wk1BZHrIDDzNmPUOhWwjYOzMefLqfKgUVPrq4jPRU6
qAUyvHZkob2mvmUZieMIZrPn1pIbbun3aUZ6K0vhYM2Nir2nelhJvSdUx9nLh5Wu
aX280Z1uGrf7aWBDDuzsUQ9TRFYCbhj7r7EIpc7cKDqWamXsqrg+cD/puuEKV4IA
dGRf+cHi8KRGDyyY6LpVIiw7FRV4U6F4sYCcllEJSc9XOgl4JuGFafOdkKn/3Lwf
zhnwdp8YvVm5MdeIDjIw5EXYDVo9Hxg1QcCyOVZ149JdYTIioEUpvsqlyDvraFjd
euqKElodrNILj5g1pYJAfglGnp+GOWRtA3CzZxORaikj2lMjFCxhcsTBzsfnai3G
NxzZ63bfHXRvpggcF162/2Px11wFZqWiknTE9jO0cEHIVMpqbmef4NXgpZOnPD3w
j/6c4NCv90zZbEE1MNdyoEwG4jYsUk1gIgNJs7+g54XfoQmlJ8sZTq1Cv0kJ1VVm
esnQ16yCsGCVQ33WAutOj+1Yo8FP3djG1QOeCQJwzOqcruuMVDSsd+lAv2Wy107E
W4Eq1w2S6DeXgQ4H4dkDzyIEzAo2uabYNdVfoWcR/iD5zkhJQD4kfT8kjCVKdAh/
RiY5R92qfeWwri5eJCSw0DEsowBA4UYgsO8Nk3LnWhv90ZOu7p1kHAoFPTh1Hg1t
8IcXPdEorz5oQG545JfxBDSOPXAiyd/I7mafBWZo59jidZQoqDOSHTl+A85uyWYa
iBi5M3p2qYPXmiOJbAEIHiDzotkJzhDqgW24cDYMQ8tZiGFrXo++pin+0JR1hV7f
8KcVYtEaoBeBuG17gktGZ4QwhlCADRLQaKfo9BH468PGCJoP2bpktJRl0Tloha2v
qkRGeBA0PjnrUhf1/47/uSePqwNRhXDrSKRGaFEGBuWx8ABfJx+QsQNB3y8jbmN5
ElGnmz30/bP6t/A2PpjILB6ijAzOPONAGcqmAXG28LNAIt8K2ys+IUUUmF5I+pN+
k62XZTFQdgbZjCSkbKkXj6PAvIp9WQJL07xJZ8X90uGerYuRnHcptFt8vE1Aza8T
oP7R1hYC+k8CoN/9NbLzJkp9hs95Yk3oDxPl+P1ehOL8ZBVMIW6cmNNRnHKIilEj
G777vyypP+ClD6fsaKiCwg7rGn/GZtCxB/6YsKhkLZcn9YLjVZ0vmpfoQiU4eq8f
sLLnv9pV+HUkRPm4vIu5YpMSzAkOV6bqvd5okX8T//3PXEWKlS62qXxkWWQaV1Og
wuXsOUfdhsF5kRr239qPwAXIGCbmVBopfx6UDnBC0YkhppRz854+pmm0xAsIJYkB
p6AWy07i1f7qmNL0j0XVYWcICxHDHGsa+XbSrey8WA8Fbhz2X2b6kOY4O8JwdUbZ
Kr8xdyP3czpOeaIEUQWkK1sHhRLH8DcGHBRuImqseKQJFvLki6YDTJvsQKgaRD9/
9Kjr9KT6Sh+TJO/kD7U/zF9scS6UYAKHzhI4uhi9UNqShi2xgClF6UsYw1ibUD94
bLEC56luQZG5eavZ3FziMV/gXwczaufvAYwlug0TjcPAGDUO7OHjQAfYQI+PwQVB
b1HZARTHiOvkqII7MwHUdLFQoEMT/fQXHo38B8mTineSvvXFJlwyPiLjDl05aGuE
pwQe4NWQp47hmHSxjOuLi1ibGKxzBsp2NpGakvp+1/Aox+9CbAeiPqZiAYGD5cWV
8Sbn+Tro+thUEq3CsQ+M1nyhBbKOYSV/r/sa8B/2PKyGjwDU+3N07yClVC3BK5iv
WbI2RkkU9+K9SaWfF257XNcogttz/UUb8LNzpG59ClB3NLMrVbR1xwFpMQ83hCVj
PW4T4spfRB+bDdUJ3Gig3qM7ES9U2ZAGsz4d2Tq0vPrjZRIvKx9H3OqfXeXeawT8
Ix51TNJVKISP7RkeB3RNaqcgOheLN4cpp5AC4WmjuhwOH7vl1KI6KX5ZboDyt3SE
ExPqBki0dn6YbR03JGi94cePt5ReQqCC47ZR79te3GKzenX4M/MkI0sCnJLnM51E
2n/V1oD8ioIqcrldo/oj6DyusGEQIAesozBZqq9b6DGSP4vHKWVBpH5sbHs69Py1
9slqc9uej1drSXg45LFP7C7Pj/xlUdDNpcwRGWSSgYzRzi2+vT4zLfzzz1WP8ITw
UwufS6R3mdJL9+npE5cziNeT67iA8swguwNYpWOfPJczqyyGjBBRHo1uzKKjzjbf
idrUmdimHGZuBrfAULv60LaUh8EeXveuKUdWKecv9O3eanp10oa/oFJXVT1EHOyO
Md6/Ice4grafYa7LIEz3Z5uBUZERB3WWdWr76WF2a/FSVzT3uO/Mqq401tDzZYJg
1BCH39soSVgvvSg98EGuWqK91TdDf+hZ5b85iYp8l5iYteniriypvTgRQf25OU58
I70QD5shFwc6mDf+2I9DO4E+Nj9M+xc6uad2JisK0M2GgFd4rPPpm3sHQJkGV/Av
rI8OcoDR6p9MG+u9qRz9foVMVQIVanFZSo9y1EZ3qNICmkoizMXKrZGwKkUO2ImP
+70lQJBHI2V0LCROMMAtKA+0MOps+4Sd0atPsL35t2ykkedelrzn+t6BNQqM2sFL
F00EfX91Wn0ACEbvvi59t0dwhFVpMkPmi41SCKrsmNpXFPnJqXYa0Y3P+Gwsmz+S
ewKB9AvCZMUF9hshpqmxEZI0rmgbyum/veT75as5qQjbgZoeXrbM1a7wKidb9/ch
53oNQx1fC34UjBIwKI8fNXsd6wIk5CcRQpQqQy2YXyX7DjXkMX2PDGOpWVjm33fv
LCatWQJGLKSHZ+Gs9obBGEXJOd40FWzo/BdgUUNMF0+a6B/j9rvWFw96fiZ9Dirh
PS+9VvdOimwoL701I/wn7VU/YC6oIpv/lxVeywBbjY2d0lH5fHLTAuHEmDW27Tp9
bxHONYiviqKzHx1OuROsgp5QVa9glZGEPUQqxd6InFMryCptNqdeJDM7jN57vHVY
4wL5IKde+zvdUE4wsu9s8kqA2GywfLm1Z1us2WUgKheFyG6hoTR3XEJ9D7XBr4Uz
ruWQu4WTeqlkNmv89Vql8S4jWgMx/wksG4vSXnmfmmOn85YmpjcfJ4qvsD5/ZD8N
wZSQ3N7FO5SghBbPN3Etz7ZM10CTUSlSSgPSV3q28JNZtz1ozebd4QYt8MMj3OuD
nFzljob+VqulU2epaO7HfjarAKd2t+dJDoteuaMIm7EcUi5pFfWJyRlzFRxadf76
cJD1Xqfc3lotpFEE5kE5TdrcJsY9FuSHB6CHZDGQkkMzshxbA/YCUxdVNlTdyF+u
Tphhgjl6awi3lCswgXJ816oj+wPjszg2vFUqpFzWjjjiUeBT73++SIn8NzqvBpB/
QQpAOq+x2uh/AXLW5zLoCafGYZB6GJddTsRb5mDp6NdkMB2V9x/rcVOjOV3klQMT
f75oQHmtKNbCyOX9Djx3LDpTqjK5+4RxgGjG0AJjHxVJAXBIhFNogVLJu3b5w3SE
AxlHYOzsiSP7hBIBtTlriqZIvwrfoGBCM/y/Gsej3mKXj2cNGc/LAaQReTJuDZdn
IDmkjKYqrmxM+5ckETXHaRzu5MtQ6RAa8K7QjIwzBEnpVu4eu6ZKbKTXZkmQhjOi
E5wZlf1taxyppALZD5Bx4Z8+XQvbky6erg3rArULMIPuRMszvY9pKhzdbm4kxrNM
9FDrMUvFfKoOMq7UYhzER1rHFGEvOKGjfklKM15/Hbba8YUJSpDgNT0MkPsyrbLu
p66IV65AGaazBs+huxtw9HbvlFKiYWRkBVDDuPzEKgSp0IGAFZkY6GjB+kC0fHJV
c6f2VVdsovwEs6UjK4Q9MT3iOu80TPGuCf4y5g792IBZmV+pDQSbOmGM5Hu9Z8BS
1YOzSuFsZ+QmhOXiAfL6LF9EVRMFFnyao3JjuOGi22OTCQb1rK1EaL/2B9RLPKa9
MaQJ9veEsJHh4v42qFZVkaSxSl18+ga0bhgq+l//HnE76k9asZCXxolGn3WEAK8I
eBkij9fpIdmfoXecmP9poqiZfwgJvZUxvyUjD4SeKxy/qtFB6GTonJNYi57oPqB1
ee/R/MTva0PWt1I/Pa/7+2I/YO/UNfwmRPMZGO3fwAco5nhUYUnE4gLV2zL6QGFj
vXBsn8NViW1flsmp7QYSxle4qCdEpY+kXiWKKecqbeiX00pNdNTRxW7ee8YDvte5
pCN4sHNmhWilkdbm08ZxbNE4ngtKrETQT4/bNwnqC8yFkcyU7l7tfJvVwM2u/s3P
FcBYi8q+4YoscCuc6D4zGw4DF+diHziN9iOlMcIlt1AMCtaDkfchq8OWRSfyhrCS
YoDJ7li3eeepv+L7OO4SWRWyf8FFdIrSX+Ay1ajFRx0eRhgdYbRWJpqsLrGYtaH2
0Ew3kP31ZaMnfU3BtNzV6DUURw7tw2TlXQaLrco2iyeOfBthfMibPpd2Vm9pV/m7
qnX9RWrK4tk+R8I+LusWNnVJj7E1bkw4qQLXnKfe56YMo0Ue+u8SX/arMf/BbEbg
4fXvTKA0XIGKK3miSYVmgKoDlFNE1KO6NGYdgDtl2BWTIuiIFSt9xaRf+hL1kM6g
ihXt+kcSoNjzAs86SLlVwowl6a0oWgE8Cg3BJv5LScEUptFOlbHscgBwgwhW3uSA
HMg321iQ2c/2raWXvp59CgDDHupjgIQfRJAYjufd3Fgyq4ZZYsL/p1cih3vPN2kV
XrCqLXtNvsse9Uqd5lIEfTsmHKfHSxufZBRTQxLiZUA8+3SQkB5gH+feZaBGxVi6
Bu1zXdEdQBrw0y/aA2p3u8S4keoTd0AdXEMmRaZRjP7L7I//iKU4ms5/2fDkc44k
kiGwO/zHdO+6gy9y5uHXCMWd2Kj2e+sGwMPq9LqtVzeOolXQeJw0gngtbqfgtn9g
GThdJ3jkx5/DaXBMks7NGg8pa33/877W5cqDpVkOo+f1nBrs0q9x3GhvAPwFtvd7
b4TPZkFx63Wv1ssuulTUV8M7YTtDPqQd88RVP5L1LZLRDfCTzSU/GI8yGGnGDSmr
PTl3LaV6qdPUXcddaHVc84koIckEuXVrAOI1ex73bLYU7oTUmrdTKl60Nvu2MXTr
nEKP9D09VRyu57OAV74mP2LYan/tLQVRDckGJdsTRkmk6gvaUPDivYRqsD585ZAO
27OjGbIIEvG8qWT7dPMRIlG6l7d35j7EQ2xHN2fwcplJTw/5pUA3kQ/bJzeBqnw3
JzW6+YVOVrfe3fYR18VSOIIgEHBPPCBYABqq9O20WmiRbnTGUcCXKEVRRKz98k66
mPaS99brRBJPYdX4WupVQqMDKtJEM6u/Y2UudK2j7BwD7WWp3v4eC3T1Nq/Eynv4
MAibrTNNFypAvum/fOW3XU2EPmp5Or3WTNomXbhAxTILro1UdikcPeofJR7QQLop
60/rERlrGyshkpHNM0AFhAfHjblrTrMOYIA3XyqaM/efnMVz7Tw4Ev86Vgu5HJHF
HGM5w/ZGtK4RlSgDi52BEijtuPnYqMc+Ekku+eAYf/0s9tRGLxMBUm6IVzngbxh/
1Phn/KzzpQ3JlLjRFeR5d8F23MkNIc8AilSiDqg7xadeWYgNjWdc0jC+v37FcK9G
/kaKhp0AdVkgFRoxtxU4V5D75x/NYcNrpK5Vr9R3voponitoUq37XJxOLaAYC2tS
yv7lMcZ375ckHRNMsn4W8mEL4UkWES5dDtnLEvvt8nYKNZnlSoSFhr4FkIjfLSEU
n3RclyuwNnvZObG7o50j6hVFQp7ImnPrTTBo2Y9O0xCvy1X+sld5x67oTuVamSs+
PRfCe4gvI4RJ0WMFTbKZMJXzzP7sogl4Xg/0q+NHzCk5w4IUkO3xcoPxH0KJumt1
dAA0uuPdaYbBs+jFatniU6SabxBa16uP74Gk+cJSb8JuQ9linoz9mNtJf+bgj1z8
ayadijc8k1in9ShbUgZ0V1wsUnBX0T0mVDtlgY31yl9nZ5vru21zUZX6BMhpBvcs
D/VSYfO1qGYqy6lSoewW7uURAjP3eQfA6bTibBk88T8FwW9wPUOaDi60PrQyeCgy
b3Jl1zX4AZ3vdsYl/DirB194n7//3I/8AqvBC2iiYRJoyUM9xt2HMR/ZHTrLxEQ7
ZsghSljVvwPetq5bCd+xhFMOM/OVdIgceb47t89sDjmTZwHqa/xyPtxAbNDPgWZO
tl4RkzCweIPNjSgTXoe3lAfGhW9wSAGUUZ9GlARi/VgT3lHoV35qlxQRQr840lGJ
rqpOVWmGcChE5rbMc47WhEMR0fKuos5kGy3N6yS+8idnFpOLP2wRU+R1VDUQGEfN
QWcpfonn2vR11/yVnkPijQYulXhdN37DBhYTV3aAOC4/qBqqoQjO+j++FLK4qI4X
91g0izf1TbrvQJq2Ru7CFnYpujS/JcCnYPcQhkM3AhwrVkFE/VgkHb5ZphXBEHCG
3N62nvReqw9U5Cbb5U0XOFKQn9UNY7GzStIxfeXB/a0qWjg/tX6tAl8GFXMFEMNQ
O/3L2Nte4stUF9dpX+s7E3Kw5LIYQ6Fosudfxf6vcLdNzqb3BonG+wLlsnENZ3Ao
2nCMVyToPLSvmGreHg6oVVXr72EvWdRtTYmhgDBdblgOsq/8kaEQ7bCjbHv3cWic
KkKbbu8QIMiHOdra459yvtj9XA21uwDdwZoFxF+3P4n1ZrvpXMOpcttNamFXGd8z
zYiZ9hDLzQgHXdb72thY1kzdee+ZtiOkEW4/alFCObZqPLOPPUJeIgfSLREt+7mA
qlQxmUPh4lXwJ+PWcb7joEqG+jF02z5xZpFmQiL4rBZj7XiJ+wNgT2TYyzjWoX8t
kCgWyu56UX71/nvEmPdxwpNlLGlgTWllTQ7snBtoiclRBsIrnJHnp8bpOJSVV+X8
N4HMdhWViSjjRHNC6+FT7nVjU5S+4GXXdJYuZkp79khNtJZ9nSw0BH3zWR28wbdK
io2C1w2ioh+AvPs1/xUCi3R6QSCVfYU8JtGRWgvbNpz7hwJK1W5UqBa3bpmb2pBm
2yhGlmnfE1bD3kbMCakScHYyLfhvvtWR74WMF1PrhAgftMdGexDkSkydReWC/eQT
Fgqh4upXUDIMIa7gScZOFjdiMj5TwOpVDvHxFGbHSKNlY1joPyHEX6PraYDyFB0w
DRWAoC/5seg9M0qfXRQ1Emwh6Dfs9huYlcNOZpoeWZDffmJrSKpYRS333cAZ9g7w
XhzrFIndjm0sU96Py4mB+fDfekZQUypKdjg3dkcC1ha6iXNUKblEgUN7kDweJ5/y
/iUR9+E+tojivc/rG6FkJfNjkLtpymTrwZVvdF/HdYFznXgfoWq7pMOKhZmi+h/3
PZYcYFicvHA5gf+75NU83a2soSgz39dR9g3DZeLz6pu5uEwvuVW/d5yOtFnnWSZQ
WLf6DSUDA4LUkLOZxjwIFZD6286dUPMcVWiBlmOHO5HN3LUZg/9Ht2jbs3TuoJGH
eBgjnAgvutni8mDgIr0NcRR4IixMxSSz/j044AOZTNgeHcHtorlTHo1JSp6xPsyW
b7fTOHHdbF4iiMOf+ddWjv/Sp7yX3WAsy+YFKaKHim4W4Fm7wjSw37ijoLm4+lkd
bVyy1it3P7mPJ5WB5s/tHLzsSx7ZJFLb9KvLyHYLdp5q9TFTAW2uGOVH/xroMPFN
XZC0EOtILTSq2r8x8lnXJFcYPwjj/im87kNJJvO7auu4AsQ/bz5oaPESBJulNQXx
+MjHdG515dBrV/7ybBnlY3OLh5NPsaPjZN745CjlFNQmf2zt4A3tF+chGXyRm3A/
JToS05NUU7i9E38dXpPVZkW941Ozt4Y3NhrupNpnu07NlVGf3q1f11ZVhV+9W73T
hRGzb2amgZ3a5Q5i15nR5uKrHO0fKSstAi2MfZH6xpjGmzDsIwzXMZr1zTlt8FbW
INIoFF9/Lf5a6o7T0Q7N6t6DuwiO0cCbRCw1lHvnG659Eqlxr7zuxzfQIi8HyjhL
qLgB9wLdJd9oIxdTRHwh70VRKzWXVcBxrzbBK9DHcyyJy0VzqrK6CozB8xKz8Xna
Pbo/Xqw+eGoBlq2UOp041SufCG+pqrpIN5we23UrCYoWM5u9iwb/xR9WkMxkox+L
WYNnCFW+TTao0fQDhKoKjc620oLXp0u7nYccVgj96wjXc7PMNNYFd46NchF3MBFk
nvm7RKAyqLLh10rgDCUZTpVOAesgbcI/d3cyQX6VEaCqIybibvxSM5UujWf6ybU2
aEEUbfZ2MWG5miUK16B3yGGbOLVtEJzL5kzfsYZ17Y8nh2i/NiCMoDgADMs7xPhx
y6Bfa+F3As4V5yvmMz0w1O+wU3xkghPu+FyuqWe/8z8gKTR7aQHbRzknYOZ5Mm9e
EyPZ3033X/MhOdc5aS3f3dwJwglBV7JusTC00YhQvUAHq49JQJ6Th25AstIQEO+T
/99CEnGqHOM7Sp+AHDg8Ryygru/wEVlAZnhiD2BeGOASdri3HW0kvNSrKXcRV1s6
Ltxt5MPTUyshoBSMo2y9mfmJI8cj3HahezjnfppRXM8J6G4wsfO8E/F/QQ6iuwpP
jqf7jcQaRqbBPKwx905iYPwPEPEV8mQgFFwrn9u85iyz2VPArTht4qRVoveZrRSi
jBMV965hpY1s59PkTSkTN6Fbpp/fmuRUvUUVctXVeG5fgARSFTQgzfuDCcdE1WRE
tYQFVZFSfhoKD5bIwvas1RNKPBIP6Le8d/iF2znubNN7yIVrmL7bgnuocUnjYZzY
7UpU7yQYt1I0yWViaPiEPR85RD0kufa8tyqDjOVx3ZoI9v55SluyejCLA7quuVsk
sqNtm90FZq5+YMZCNnR5h3s+uxyKxZS92t7agiZYgbibCKBX/D1hxsAgR5njvXLQ
sH5jnZ844i6CxknE5NAaBOu7SxJargTvpXWQYHy11JRMQuySIx0KI+2Dtfl1a8Cr
6weYGR9WsHVnUB9LhoLmfSiALrNK+qiu4OouqsATaPG17YiCujKrnOF4s/8vpWv7
nOXkTli7BHFaBqhb7Gz8nvyo5lDC+BQRgW883cXCZ2H0YV2S6jf98BekyaYuMNLf
Qm/ku/jCbLgPDm17Ft5D0i15vpO46P0o0E1K7FtV1G5ZuHAvyKiSrRx0ClIUgiNH
iFyQ5hR5VRZuITS5H7oQ0puyE/EtKQZypMUiGeKUUoYAI9owMgHT5bWJ+QxMtBUm
c00X55MO3kWs0B7jTGqrCR1SAWJwBXKNIxnNqm8S1Gt6958C7jvXEiKzaW4ZxQbN
mSxdc7VpT+IHe6C8Z2FNT6g17AQl3iQUtm4+L9R+dQZzLCKATU32si6Gd01ZR9Of
OZ6vNfQKhhGKyrmQcNzduEODMw2DDq8u7NWdvo/1ULq5EnvIuG54k87NcUXarqeO
ZtwB2avDHb0Wf/GS+ZrQiZLV+kFgBc6Jn2cKAJIR+WTeZoxtokmBJ2zRPRCu7Jyh
v/m+IjfT6QFPHy8C6cbis5p7HF4h63Q9fA2sgATuxCNn8RolSuKVyaZtK58Ut1Qp
a4XkWXRyoTmNelOlr0QJ153GIn7ZjSZuVYwoXvL+rvZ889Rt6T7j/izCOxrnwcFz
sZNvl5DTk+/D5UjEkerXhZqD2M1BFzBTiWhFFvrtbqSw9wu7yStktc4fenmG/4rT
dbQnM1IFj6qb5chqNtFRt+3R96K5vlMCQFPr8CBMhExtPXfOLl1drrLDHigfH2bh
H8ztSko3ZwZ5I94NgCOYSItXKhXjmvlQ1ojPnThOJCxZozVVcJSjQvyKS4wpAEOQ
nTDL2EwKAdOie5OyTGhzJr6EeNQCaenLYs4tIXin76HnX9YoQmF3nz7tJTgGKcrV
Y5JgC0O1onXPgFr1rA7f2hJkQhYzeK+b3tzSYhKhhxCm4tCCfu1g5KG0Mlofrezs
3TUJ6MGQov2DagVqkfGJmIJ1Q/nvdX6i8j4r0ZOlHH/18vmZNWNcRsQptXffKcF+
G+qIcRdci8B892a+8NClWX9UrDOJrycOFRyqyCtBcuZoTKfpYmQ9pV0NEzy+6ASW
UuxUCo+BAJOlf9eep+VWl/dbbUskrVseLkDsw7gtitYHqBfMoQYn522Jrvzr5dUo
5Q1/+4N2R61GT5DlySJaCRnB4cVg70sYs/8AXxDDcf3nQ8bY6/brSQExaiFiKv8D
9cYScaPkPMww9TEQpNzChgR0GuFS4t5O7d1+Junh6zjdm9O1ncSEhukumw2Xbkwx
cu3gdct4l7mJ/Uqtbk4EmlECSZhLgOseLHcpeEooxtB52RkKuzra7b9+idLyW76s
tEf9bKM8png9YYzHPN9/ESXwofBDo+0YgXrbdBa48qCprgBqi7858iuGvcehZTWr
QTWdBUm/pSRslx/4CZk4upV5sA5wcGG5fgy09SjqcC73ltYDFhtpf2UNQc5Oo1cn
C9da1B4fqVgNExk+klz6MprpxeCtmAPHRrQE9fZdrnYgrzMxjUV+2LWrsu3vGByw
F6XMWhRaXwmxvWunL1m8WLGttC/L78PaVyxIPkSr7mNz0yRedvy3dBJY+f4ZRKRk
kVTX+/eziuuRHK4uEqW9YOqOKdr6pFbM5UeTe+3wqrAVD6WOF2U2MTa1Ral2qdf5
yK2Wj+xxgX7GaK5BPD3e8ogrCeSelzbVeM+lTnyeBllrwCIPppt6cheCWwQ+W9Oc
1vZ9rjyG31Z0tomhjnDjyE+c5PpJyIO1j6MCrPvjEl2CbsLOBSYa6g/NQjBl3k0+
x10bfnLxVFbZu7GycnOXMa8ja7cETcnGQ5IF4DffkgOT2lIooNqDi2H0EOlJLvEt
tQITOvTUIkBYwHxrwtnuNNd4Nb14gjPtzF2utYaL6gjHl86dCcRo+K3WkWj0T+Ba
vozfsBIZviT3FKlUC2MuuA6tcFlicwQeQJ089sPmDOrDBr1buRrgEWm1j8AM/5Xg
PUKH9O4/J+RQAnebvwTcz57wIJut1XR2pa/o0TvaP7HzqTdV0X9KXn0q7vGqRnaL
vjVPa6pbLzVuFhec35F3VYQgYak/23Bd9hn8lqmGbU90+KpQChd59CERuUwlXrvU
AwLW8rx8Fo+HViiwnIYrim7RZ8yZh/imOoWOWaktjY6Gh2OjIhi7NPx4h+ZKwFs9
74jtS+RrwNcKeOsFvYukcB5U2u2ombGlGSD1hSnPcsqe8AECsY2F1Q1mugK1VPw4
GU3ivwNsmkQp3W+Ofebcw8UusjXVP9OdtZS4pyIf/xzyiGhRAh4HZ92s8zXY03Bw
Vtohq/SCtUNXwwwrkKv1yqypWpXDWZlMkTqJGAoXHj7NcwXlSKA6PlBcnaMhF8VU
uONgt1Bu6cMIr3NdJVsBwp8X54XxP4Tp4FYxLTWZ5SRuWtRVCzuOnlKT46DO8NEb
kkP7ECDUTIUKMIbR/+JsWx7G3y3d33lgxzgzdqdEN3aYwSGVA3j+m3r+EnWZRXJ2
78gkDiuojus50VdZ512agkpyBo6tlgCXfo0REo3uhD41w9s0K20BhPnl8HKBPLCS
hXpuFsMS01JAb4FcqNG6nQ9UBDfznh3EiC8Qgul8WmNiiBW0fyGtyZdJ2q+94Ncw
OJOp4SLa9G+WOkEY3ICYxmirmnUMMXBwvrh+5RGP0WpKPnvpqvOjzViGwcCPGe36
7rIOoxlJBtO4fosu+Vgm6nBamL/Fm1bQhBxQ+WE+2s0tQtcsXXdvRb1tm48V1xBO
fk6NdLw5d1oByDku3EzvyE0rKElHP1NLknfDX2qAXqsFO5+sZQ7A9RJnbohw4OHo
r1pTy5u7zUo3G/K/of7P6kvxxjSoB8w+SGsuMIMJjFfCNNPK7nWfzeQz9+bZX0JQ
HbkIf12cmdLSZDG/C8kIEETixBaT4DKyUz5yDul6ruO9aFlcFfklpdOx1R2RCF8o
bmqEM4tak2H5lPphrlDQEmM78gI8ilAdrWj70cQu7LmCybly9BtqFpps5j7DutQZ
7uvG4zbRI5c87UG2dEr+EC2Is5e/KDmkYHT10FzgLrWvagPw3cGD+yxrQOU8U9JQ
k4hR7ITkfHHW/6Zh+xZAvZL5B2RLkgrJXVnBKVTS8KAW3PbFjWL5Int+dlRvaseu
adwrE/oVScQa893HdihrtTccnmAJqQ5YtW0OSOROMo8w8Q0tgUuwtYn5pZKyn79B
c4fdj5xDRbPZIblvV7Gle16+bC1JWcb+VKMeW75qZn1mvxdWQA1bUZQqJB7Nu33o
6v7kNVQ5mekvjZL0tqpJnxBqesX8ewTniIIzUuxgPJIgcREx1YLuzzKBx12osm3I
OTYvXxiuqd6fLOZglhZy3VbLn0dpUCyF1XxS54ctYk2K6nBwX0yAwUB2YkrHIS4k
mdRkWD0LxOV8EGpaL4YyZisGDanNMfrFXm14aZzObEw/z3zZlny9yixu/pGnTiV7
kLwK44psxNpBSJoW8u0I6e+k55u7njrDPY90aDofCmD2WoSdELFoZl+0XGNXrOcJ
nzk2mqxSFBOgEMjuHP5u2MQvvF9+xmXa6V3IQOfTCKQy1N6C8u+2yhx0zcbLNtvd
Gd4lOT9l87JNQANbNX4ehqU1kyfXjHUv7LpvMmFl1/z0fxi6DTKbBSJpJXlEM5SZ
XX5gYNO4m4dk4RyQkoGNr/O03CkTwSaBgeMJOyr6ptr84BnpO1kiYF4yOs7kOJo0
vFIFmBiL6dp2/KTJLZXGknwiNihXR6icUv6sH0lIFw2iUez983bHH5uoS0+cjxH1
JLmIktDJzTkeeWx4H/A1YYPhD/MHQsnpXKLSJJ0yYW6B3j/0rJslEz+xMQW7Ovy3
cWQeCyKszF6262MXq7T8LDW3cGT4g+xGf83mclslEzeCr1aHsXhE/uP9B/Fmc0tj
UISXT3yvvE6oBIgKGlx1t6FGkRLLc+7IteKF3i71/wWsHyyln458OxdK9a5UOsr0
dVL+UKmw8NaLmYcVzG9Iyb2nAUbEdgE+n42HlgdCbewatM7+nUAxUNVbOK0kcoZe
pRVmGfxi0oDAjetkva8Tn1HKkfAxXcP2mLsGvwcw4dV3es2935EiSgjr4rFon5vQ
wcAJMMBzWWAod5Mx9lSCLPme6rW8yeHRPVwRtADmWXA=
`pragma protect end_protected
