`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
InyJwiLLWdXaVVCUWbzo5wbkwX71/2+0fgsDzuQN6VQ9v4oNpLuPCqCi3C/Zgr2I
3oTu8SW1cNMAFel8WvAL/VdNQpulozxToBxKtR5d4eP0MZV9tI3TsWcNnSA3ve+B
OswMCAgapzmdw9cRS3qPNFmAhT5C7DnstnRgiTiZ4R8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10640), data_block
eq4v+NCcG1rJVlxBLIkzrsm2ycCTJuuy3e4tgAQU5/0CV0HhFdKfjc7dO8+Pk6LU
lv7/0I+2L8jGZVS6OQk6Uz3Pn7VJFFVaBqL5uKWO9JTcWLrKRBfGJ/MaPbhL7PkW
3qFQLTU/LUCkQVgDlQD0nYQrRwamwN3UCabvHZZd9C+uKTdryNDJJLV0u1JvcgnY
/dqjf5sJmTK8/zh82poVuJ4hEPmLg5R0mJEJekaR+TRExzwQG+z4HnSBEHVwGDbi
N5FC9yp4VI+RVmO7wQPofqpGsUWkFcfFuroDQoR0saA+TA8RotQO3ofBaL/1Rzpw
Jm80QA3ghQw2apzhtb0SZJMFAs1oXDq6H3cZ67fEVdW4gR26q5GqcyqESI8KDnXN
G3xUBHMrZCJXkpfCJDTkwzrHSoK/mZFQz2BHIa8g24EKRk07BmDWzgEAL0eRysps
XVwlK4q0ZVe4hdtaSKFFVNMJOnHzjevdn5bKTs1zujiCe0na3Fm8vDze7tMCsVWL
z2srm7mFS9k/k+3U3D/9/ypto2IHKUdnwhmcczkbaTV7CkxrA02rdS3t9/6NvF7i
oU0+xa8P+NbjLnM+FyGVSegsG5zGjC5mwaw168inK2gRGuVwqE++ZRGkuvQ92SHS
CPdEK24QeCivNC8im3amHEo4+QSsgc5Rs7Yw7ugiftTAKl322mNkxWyYxnRwMMX4
hbdP79q7npeg4YHEGYvx/Aei+2evLZxoXTMB2+fpAMoxPAIWP0OaYioC21yiS/x4
4Pd+nlVR8SbDG3D5DIgNDsD833r17TVEMJHbBVvyJYcopzbKS/Lm/fKrI29MIBnA
mG8EhIC872sLtCf7Vt9u/cKq+a1JB5l2eSYn3KBTaxk8IBoQIaJJ2jy/SMjsvTWH
iUDaEOqpnLJeMaSmhyQNymlBaKDuIc61UTAiRKySiXgRQ0n2kfPw2I8edxISzykH
LDBsCAFAqS88Szsp0esi3vihW/dbjtrXeEUFRYqRfQgLaZ24dyX0vwcat+UP8DVZ
8MRWwCHonwelxdIydNI/Pq7G2k5rXQ4siSgXMtrLokeG1foh4pE5FQ2lWE1Ew920
JhHbF+KE33JgYUWtMmBDFyw0vMotm+WqiIDZI7/b2RdpL4PR9JJlcVw3vjHkFlg+
vEPebgubyogftfrWwdH3OL/YNWXq0oalhi6IwD+hgtFd6lSxPKWr3QHns0VJ/Nky
Gw6L+CK6Mf6INnYWM7RvhBvM0SHv8R26itvOmjqYFRLO6iPNRX5629P7qYxi8Cbi
BpuLFBNbPzLHLclyaoKsosn9eJxaom39/3MxkDbi39Vo0Y1VF9npxDkIlbepvWX2
h0YR94TuR1HumX0pAq9IV8CbYxcpdzHKcXEhyz6b3HoAKdzizXLEXDHpBMMKMZes
L1Z5/rCTTJBnw529pQwgW1CQ0Ipo//kJ/BnVz9QFZlkY8avZX+y6b70QxeOMa5rP
sobHqk8U7lN1sQ0VbHzw5AC6cOFBhgmsXMNPkyPGRiH/gpR5FAmaXdbJ0yxlh1Fj
YWWVqpPXlI4iHT61XzMxzQXiihCkSrErnprtgJzrQUB4HYtz4X77/Ssk5pm2mfZM
6+SOT8MVsswrdtzyofuBdQql/uIeIh4Nh/WhZeNhDovCt/Bo+JkabOcLvF4a6NJx
/A9PnK/+Hc1dDlMNPn8OXHJo16gVdmAAkfYCoFY4cYZFPmnOhTYPJAl0uUSplSJq
HvDp5mb89pHfzwuZshw2unAaVvQhDbhSIajnPIjGRs5ZZiA6pAW68625eckJqbuY
buir9fnSD7ImxV8iIC7S9XkV39EvNrf1p0BS7Rglu7rrjMC07AkcEm4zQYTggNYK
JHszeLff61apCHVU7FixMgtsb2rwtZPveToZWO87rVSw13V9JyP+JJnGbXrWCtuz
+sxr96YYnq0pOTfCgG8zl8rqrErHRgG6pcjiv1lwFjGif3mFkWozpt2iroEBlxeA
7IF3Cru7s2VkZbK14fCks+voobDvuLVlm5EEg2bWFDSjU+2e/VZ5COptrHFdr/9h
Y+dhwKSXYKES1lrdknqmtBw9NE2IB5UryCtcBWDTiEzAEoYrVFaUSVZR5tto9m77
C00Zl3avKMx3StHgoN7HjsO071h2lcrUyTcKvOMKtNAUo+vR7/nmc5XAMu3Mynb6
en61fy/j2vzsb6Rr7VwVWKXQJij6YSMCjnEsxzJbl8TmKTrBEXfyugpg6GBmm7F7
JOVqCb3jVs0xS1Z42MVO2AWGck/HEi3SL2rvyN95qcXg9M2t5aSaLfEV62+uB2iZ
lI3MdhTxKB/wFpqQlEyER4u4HC8bYWLnw6WA0DQ7HQnl1vKvwaDPF8IO1k8ETcM1
NBnPMdOgSz+oBZdd9b0vDGu4z3GM8rDO8O0ZUZrQPs9+KK7Zq2sGyIKMgmoA+OW3
DAtRl85SBYaomCTHwRnkNW0N3y/BY+DOkCplT0hhP2GAb0h1F1U4cSjxAY1hLVc1
bQdK+/631bGlr3EkF5TSstuIa7In4YaftdQVdOBz2JDi7U4VmotPwUzwuwuThoSa
A0jOBg1gV7YjwA9ZXIbWJ7sTaFflBKPeO6XDktPkZL7LnpLI5vIvX9tvdufqXipu
d8FtrOLe8BchejlXEgx1fnb62u4kEGZugSihg6UxgzIAYbWrFJySR5YAHCe77LC/
kpmpk9T7jHj4oGR40bk6XW2M27mQva1HXWZTTc28xFuYG+QyeKDx7iIHPCG2MWxd
FB37ovcSmUWCyTB7VI7MKtakqrxEJJJCxj/JuhEfv+zEEUASzrB63bC16/k3Q0Zu
k7qm0VC0EZe0nZVln4/wjKmxOPbwy25/B5zmITeNA8vAsFZaiKU8TBWrTcmVvFaG
zbkJBWmSWS+nlVtOdrtI5T2eGMy2HF4IEj9AubMrO9ewiP9AGHThK/I+IGtjOOCk
ifIAbYggUZwHJYyQr9VjnqV9kF/Zmgux4qN7nipm8oY0EkdnO4YHiYOG/blpIWIA
hTapuvatMOoWmIJn1LIfA3qN8RT5Ypl8wtHeJVWv/4g7/Iwq6xlfFda5ciLM3ZMM
1P+2b53h+4dJKVryvn0+w+LfLWSr3AjM52mXdaFjma08nmj3xUiVRzHoWqgQUBAD
5lzLr3IoU4pwR2QaKcJHaT+PB5LKeiwEgZhv0mstfd2DONvaimFe13izpiQJn3R2
O255vOJh+cLUea24PeTtfveBrYdWd2/Iq4pY1DATdue5tzO0QPwIOi0JM7ZFDXvM
gt3l1Y8saDIerSco0Cj1IyvVE6+oSpt/bJOPOUWo3oOAUr+xOuA5OG4r6A7TJrDt
fHcMME2hUdv50a75kxoi932GjHPf+1CqNa7VrkJx8v3EbNsv9Utkqm9XwxDA3c7m
9j4HU5NR1sREDomPhuEZ9RXkllIFlg0eh+0Yt4tAs0h7RzxdG5bVs5J0+WDVQkMV
7D4F45NtK7LHycWNCPsfCrGGzu2YcsUtTRi1R9Pm4gIC0DauGUSYpj2m4yhQ5ooC
hSkHvMiUWwlWkkPE44VuKWirSSuPLaoM6MhvARRi1qVsOtAIl75LyjYGrCtm4Ozh
01bPcQSfjCbLXlV3vlsp47Lnx+qkIcvWAV2O4LcTW3mp0IGreHsCJSuhx2Y3aCKM
hd0PxFCR69DOlu7CgpQrd9vjv3lZzDC9uyE1m6HAApvin15ptGTys9RvQqxW/tD+
Eh0hrrL8Qoz/JBY+g7FrDuxmUcZKvmMGLmqWKOm5B1MX4dui1yV+3qdmdut9BHmN
s5eRSczUXfZjULutvSXPhV4wKl3NZqNyqGcGb7EuDXZv8Pn81mYnWxmNqKvmjQva
EXsvRDvbawgas07SFqQP3mz5o+oRHbyupfRbbCEIU67N6+u/Evd4NfoHVVw3j37E
d6lEhGz9gr1/AWduORhiwmuC6YVy+KcAMY6UspCKpGYojTo9nfpV4HbdlWCXQrjb
8W/eB7OaC80I6DgaqVCwwQnUEqBVLoDRTYw5yJ+9/bRrBGNnMUHP+q3Q+TbdD/w/
Nw29/4sibfgT5+tzzjD300egzIXxGYGm6f96NpkrjzMkpnCPu7ork8I4vILtUS8O
4PZq9/z8UjKHJtsbaCGo/iKtI/ckZS53UMWHGAaVwuCjFZqofvsGNcGmC7eK+nA2
0yxSIMc3DgLZbEdAxjJZT+AB0HyyqOhiO6s1M5kq6DW89J8gnP3VYTRLDWDqDQay
XqIrAACG8N/wOlnmzfNAweetAAcVzZBdnox4T0bhjPgLyjGG87n+VAz5cXSjssaP
F35Tx/5duhDTRz/UVBZEppu18kLPWE/bgfS9zSDpEJkJ/xBo5nbbOPMIH+gnc/iK
1JfDOj2heWfRb3CkIhBpmU4Rpr5vqjsxGPxqk1wfe4OotOUmE8J6HXOCVZ3iGuX4
isyS0hKP147MOsvSgSaxpda+ZImEhL6CpZbXcaHFQanuLyN+6xV0xV2GMf0/OCbF
E1UbzA/ZgAZ8g0vhZ5IvwcyU43axTeIg0/fP3LKGMa8KTT+1oX+xx6qliiYFfvvz
sW3hdFqZLSFLlRR/FKHQL7B+X85P0BOmYwPGwK/qu0Np7CxyVwXCggrTLbsK4YRL
BlheE7CayBFj2T4bSwrwkIF0BCboddTluEY0IGzavlkD0SfJZEAKgQv9hsaeCW/3
U76fxgYlbB+S812ea+oRYsDQGP3Kktno2xiIOpFM//tbZNM10LSIACbvZg8Z58ms
VVp3OA2Ls+o4jjLL3+TlW+Xs1RtI4zHrF0v53BmgDgzMAw8SQ4ldT5F8Hm5Zrx4k
IsauZvmg1WpGxnRhJ2CJ+VQ4JNotRKfap7xteuxXdK8rZxDaQgqGu9/RohXmt/O9
1uT2yZgNyFqWXlNKtSv3mTezy+1nxd90aPKqC/iXyWnlqKTGvlokNSbNCnpfc6yq
j312uHXXC6QlnY6esnt5wAsApkk12GhB38EF999C1pClFycbpCaq7mSnfDqAofBe
ARMIPzhrEpDOl60hhRJqLj8VTnYLVMwOQ8m0ToQMV8ZeUTVd9GfOrbOUmbyRksII
NS48xLisY3dU9ulNtcU45kr2/TFgZAzJG5AP/eRQduyqavIHRuJOquIS/ncPAh2Z
OHuFIVZ1HGwRvR5ucV4MdqaEFLdjBwPnLhAuFvqFYcmZD/iEBcqvX/bIMaapemIP
Lm2kTIlmAKbFCxeQKjE7G8JT1uaS4qdoSwnLW/DqKIsGKroGks7HVHpXMTOaZVvz
2tBtZNVZi2VmBNwSNmQ0wag9OIVj3SxvOcqs+vz+36U5xGZuToJCe30YgY249mRY
XS+yereqp0HaptsdJuq3UyNVCVGZctQXzW5JZzhiuK8+xuSmvmU/W5Nn257hOS3c
X5n5SEweC/HtHr5TMB6CnWicL3+7WdJHk8BZ7khewIXLM7iOKgv94aO09ft2HpWs
QU2vCtC9XWCtu85n7nlFpPSHvYNWgB3NGxPkBJNjwBJRSAQMeQjMwQMCbdSj06FR
z3O9k2zCK2RrW2yxglRmTCF/jBaw3iKKfyv68iG2MlX1bte8LTfgloxYfAdBN+Ui
MhHuYFwPJ9YMrx2WEG1S48kDkDkLkfFRPUlrz8uO23nXxT2S6d89Xhdt8A3Ba6zZ
8AMn7PYpoDJYYm0BRD4Dd2hiVD+6QHwe58qwElN2Vlg2gzNfWg/8meYAz2rnjZfH
XdZ56eEgRNvZVlnIaA8P32gs1Cd4rsvejHfv11Ny+DRPcwuoKfP0w615IXJBwHs2
WDq77vL29CM6LjWONGvacr6+RsLipKne2yUjpzRw2fnjs6xzYMh5jIbtyHEY8LtN
rNFvOo+8TLeeF+YFeEasQeJi0I2jwAbzHmH+UWA/v7mBShC5iH9md/iKCv57axlX
J5R08FjJKZFoJBHL3T+0ktnP/7LypMalQ4c9cR9gOGliaIKrBWdqaUkFH0NZFiq/
qKmqaJbYrGprNVYsSaqt+G91p4Wh+16vPof/XZlCTJ+6b39Oal3bNh0gtxE+0T7t
D3M307IZGrpejb+CH97pryQSHBrNw65wRguobaXF+rcp4RxbsIqjPVTVwQDVASWf
kuUZhuz5UaoHsLL68s/qIAWK7G9qZZ/T5/u7UhKNTGQcUOzwXfe7PLK2ISOm3lPC
whsTgR1CNHb1SenHicY1+e3IE5a70JTadvn8cYk+aG/1rDn2GRaD+0HJ1iYGE9Vp
cfCU7J34C8jpkeeEViFvUcS9M2qrOZwVdI2Liq8cnxmK/F9iUuQ6++POfBGnjwkY
yJa842LI7nGWmFZRbo7i0dmPqysvyDSDUwm4dVV+whOX3ygCYNEJveEbPaglNFxI
C4bT1aIZ8JvtZwq5IEBcme1vKSe7GKPVmg5dlmWHxAPsWTrK+4eev9kZkLlBxtVC
gMhmuNMuoMQIQ6FoTZxdvADGC7906YGEYjyQEYku8dL8pWu2DToy7qtHanii6KNO
i7waqpqVKeBW3NhxZ94DQf89yQsHIcSOeJMkTtohmb6l6oRcZrBifTfkWsubSjIt
JzowFD7fntvslnqTfUhxGNbLK5X2F0UBmvubb2Wf+5R5VaZBrLLZs5Bo0l0iRJmo
V/IOmjFryBVvOZfGpfrLGK8e8+s0zMCQzI1j7dwcRqH1E6Fc1wqpKYzL94ul7J0r
jg+vaw7i5JjGaQ98n9dxljCyguyie9dodCuiLl+Uy/gQrjgpo82wU1H9g3nEyirY
NH/TBnruVKKkQFbXP2DEUHRYQC8O8ShdA59d+FQVLszfvNLLmKRuryHl3qgg9RlT
wK2PB8NZmkpFQHPXAw3M+EMu+eBdmQOISljEQwTvd6tsj9bSowqFmtKGQPFA3wCW
53VZsQtAzuviWVSVZLN5v4vbfsr5+T03+Q1qBAENjrDp9px0Pe0LrCDUM1e+vETU
dWnhMjXHuZCkHK6POdS0sUGKjzJ6QcNyLtj1j9CinKh7ioV2sfIsIqbZmZTiQuTK
0SDuoIcgr5eHfKUerpgg3Ncu9GDOgy/jVR6gFdEs74Beb6imWiVmvnXm6ELSAeDy
jOYbKnXKZKWHHqsMMEk9fXpoO3fj+TlvGONrc7D7CuGUzlPDBaBwKEnkuXVXQs3N
EDJ9rL4RLRb2KDpx49b73AeZucHQ3BzNR+VcmgEfxoeqVDv++JzQOU5i94nmR/NM
CNAG0CJVOHD81n+8S4sUi0QFRkePTm7VZYYQ3CpzL0wqKZMjBMRVT/7qDSF+e0jW
0b35NlGzpZhRltd8dS8M+RjDteZ/nr+dFhymJuc+ZIY1CH+08ftpYdJyXaFZcUWo
e3mgGYI+B8VLK3Sfjcmfg1ZE69w85oZusSN17Hd1dLO2bajLF3IfU84YHb3PvEAY
ofLQuHLXIpBfpIbuQzePOklDaGrj3MLHDpIpCWDvfYk57Ef2tt86f4fVopr4wku6
rW32YhV0/YlY+HXJglmaPZNeL7YqZLbc2+94OcwKMCQD9nn6SEK71tjVvgcUzTKZ
AKkFM95cvy7y4dL8vSBpV/Vk5WpYeHBs6dAPgBSxbm7OKayIbolVv3+6NsDPGQeG
ld+qjW/alYlN+u8ow7Kp9/4r5fj8iUrsJBGMr+wk5HCuoz+PngAtqOk31XZ5DuK5
YIRxU0DRfsx6xs2/nAo1o9gOj2Z/ToZE963/cJvN4KZfsE2OtoJIM35iKoMlKQIg
GBkhrBeAycCjoCBu3Ntw3YBM27udcnjesbw5kw/3mOtAMtdIpAWtflWg8+hf6aEN
HFeJqKjPA0gchXUV7wQFE9tx5e7pdNrfR1yY9QJEvrXWE/53rcp/1P2G6tqiWFu7
YG503bUyt6RNNmJbH43H0toyJch2TfMHar5nAAZF5FDi4IbLw3b9Hi3B2tD/HVBr
tP5kWlJEFz88PZDzwnnC6VZ+skF+5OPfd+sKirNwIsNvysldRGxxOVKm5+dmq7ZD
qph0mxMtzOivxV8w9eA8Knz4y7Jsq2jvmRxMBLUA0fl6MHu4ysc9fI5kd8CfXk0I
Xz0yeI4oiLG7GwL3/I7xiCM8G+DVS8HdE9IKXQyJVZluSCgauZqpnXMT5XRtnnEN
T/VSXu6xvVb1gfkgrHKQEkFlLMKhhjnnqp99XJ1OXsQLB3yYWAyO5+yazfO+BQVD
d1Wsn3vG5labWGk5EqfkceP926oBtZaBiimuC+h0b8OWtneC9lQ4oCWBjZwUAJQg
XjL+7hdlodnDip+JGH8zPgTclgpt1g9/7ZnvPEeH3brci76Jy8Yy0mNzNH5LPDEN
FW5809hJFQYag0fyQaDrHnFktbhE09q0Q91aFI7/MBYTsBIxqxrGoK9erR2IUqYq
IowbKweOsoAm7SNdHNCFkOG5jRwjvF24DWHhBWvrL0WNmdzqk/bf/9EAHzeeNUeH
BryRzlao10yh71LZP46h36g+KNlNA8DGt6igvToeUKO3dwk7j/l2EIu1h409gZFv
8+R/AFnMtpLS5U+S9/J8n/+Cwo8B2XT3u2wM/VWVZu9Q3pRFvcc0mKOb2H4qcX8v
7anHrhZNVfDQeJMwhWqa+66P/MkSMT/hrgqi7e3yOU9feNhpseQXeTKRn5/8hJHQ
s/9UwiyUMwXR6uhIv2qUJvNDr9bpjRLejP1hrvMvAU0Lq7eDKOEEJUcFf0wFyLB4
55igSbmx6nWsdhUY8r1Ae1v2JrYouFWLiqp6WigABqDwre6u0J6fO8jhxpNDaPka
7LUK3EshW2EpdXtHG3YO0SPrC3WO6LujsHby0XMztPHDerGLrINexN0jFvC6ueA5
26I9P+QGIQwff+awBQdtKzHN/rPpUQPTre5njJNbV6q3PA/xIEYVZfd4oZzT9YZV
nMdcpTYJL0cdb7ozVTCt3Q3zQPHVcsjYmIutyOrU/HmEvLKi462683Vf6O43zQv6
igqyD+/xK9EQhDzaOfpvg4WzRKuVQ3qbTyoaM+C0MKmSCVsQwu+woH888C7uFQgu
kNevsxtCCvFzuRqtEFgnk9rwLbrtqFajTWDOMsXWK+inrKqs+QG+qk+uKMyzp3Rj
j4ujSqoNHqQMCBewqnUIus4n32dD9tZ8fJ05IL9MQWFrsZJEx75eJIwNhH1VcVV8
VdLNwElmKNWu+1safbKnW91Qs29jwA2Wu0Gp1fDLpIEmaCFzy6QTDW409Ak6mNye
cX01zmD16S5ir5qoptJtBOu76H8j5hgjpw17p2RNvzsd28HCKgZHTxLxOXot6af3
Ne2uAk6tMhB1QNpdfun7R2/xgZs61nOeRddcumbHo+Rj91p/JO+bg+JKJaobo3BO
as8HfUqfdg8QzFTc2I9TW3w51T4xm/b48yHM4CDCccGUgT/dbK43+t1+JY0ogMJm
uOSdNhWZnvALr/yBVjf7/GzHpddI5UJsQkoyf7zQqJenS+9NfSGpU/Fh7wm+N5YW
339SZBJlJcrIMGZPlwcoHCAWvKxRtsA1cua5FsWckU+MIaz36YrrI49cmS2LHtZJ
b7katx5Mf2pD74D/mSQJl80ksYETJ+boKsbcvuCTqodSrI3rx5U/Kq9tcVCfVuCt
JeqYOI61lLTZDk9c1SMw90pnG1qvDBAD2Mg5Cfd7ZOMo91KI2Mn9cVOStQwe9Yez
NSeeo3ztiA61Zzx0opTGEwgfuFvLkcnXzvPRga+X1RBrU/5TmYbNWXop5o3O1Tn3
PofLKT49cbCPKuF4XqPkcw7AeXYj1AB8bR5o1BITE96f7jt8E1JaRtBCJZBIrF4Y
bhXB+kw1JmlRfnY/KrceYU7cawIJ5eyZYhc1xdGzVIZWfy4Gdt2k6XxnQhdLqq4e
Zix1bJwHsM1sp6PSOOJSK3nC9r952s2OtKDwdeDs8zU2QgZXGqNQ9G5F5xyb0des
+aZZzlog01uaEiQZHl+PZhK5a7q68IS/uk1K5dd8xuu0dz/++ld2jgT/C4V4+tsT
2RLEDGqt91SmmIVa46En18ABuDzEijn1fnGQTIpMsaQey8vPcGQ1oHvTUXASGCSL
E6P5XRDuXz62c9gp7z2rg8O/bMghCmQq3DOh7zNA9PydSE40w/xe1s5BJ4pMPNT3
VKOESSiqATIwruCKfNW/sOhG21zPAHeqhOsSmNgI3U0woG1WszBrdYDO+WCJvsJs
6uci+OBXW1FneywddDqtxg6nEvUm3gvx4OE1H+8hRs7M7wF2MVOdZITKa9X1Qew6
ZfSEHHaV0aj9iqD9V1SzkobW0KB6NOGCmsfurXK6rPxhXIyx1pVXicnpxuyO/nF6
xgYP5p73iP3ngQuPbSeHBqlxKtcl6+w/HFNLV/wzHqn18PEBjhBhA7wJ2b7cW//x
Cm6oy5fK3LNO8iWepl3LkjnoGAebAw70d/xyNItqR4WSsm9ECHoKWgvCshzFwV6X
2idslih+KWOpFnxtUxGhIpjU3cBPG2mPmCAuHgfNlXf6f988fv7lKKiwW2r2ozc/
6NLcVfl638T7katv0tQFHoDC5YabysYLzKqloBhPXW3Sas8TB2dIqeqWXnbQA8dZ
JurhAkZiYeM4oxhy9APvFQr50l8g7OMW7/nj8E+SMXlPVfj96iFwe5JWQcL/58w3
YJ7ddIZL0ZZmcC0EbkgTQMMpufvtlhvIcGTdofXoZ5Z12SZugpRFi9E6Y49DTf0d
dLW8BjKxFoUfReeKZkGce7R11XoJqNSmLo34qjndLSmF6EOjpRNgG1wOHb+nGZkQ
ewMUZGuyrvcf/YMYikIuH29It/CiMdoLLQyxmLGrdTOwGWvuaN3dVThhFGxI8RU1
HDAWAPd8ncfrDtaUP9yezk/h85MbVTZBdk3bZnB48zc4m8YHJ5V31lgRTp4YqQ1a
zLrRAsPvWHBz+In0Ih0nQJCmFJ2gyBMAQ7ttla0Ci/+HWx40Ly2qWDkT9alN9on1
uS7/+jwDK4dFcOWjAfu4gAA3REbbOTNtk9vCgW3WWq8lJm74/DBYuF6iT5o4i0FG
iY/CSEFP9MORxJrZLwll4pmBMjTy5lYHyW2SGDdmgPSk46GMazrRlNcNGe00ybqR
W/k27FgWXd39YgYgoctOpeBhAHghW59yyGGGHuef9gG02P5XRMg1EX0CAXkVQcec
UcG2LmdhbvPknMKo1dVvTYlfFTGBITXtc8fMIPxK/6Tlg/MaH0I0Z3TqBVqvCQ2V
8+WyDpeUke97vQ309PBAW3Vi/MsQAORmSY3uG8UNiW9i3NhwfEDP5iivTrDhMmfT
YwpplO55F2CC9afHPk1/bJmLEaLp1fLqIvJETAXrCiU3nZfo/Fgjq/Xvhqz6NvKp
oaI+ZAWBnKPi2Oma6/GNdpqzzZAniAraKOOK4Yz4pYswpZchBTaQP3JN+llnPdDp
xNt+VetrCD64G34us8Oquq12GqHBYbqBK7Y3Mm4OVqtLuTF1u2lGL6gDtPxAKwss
EGxrdgv1x5wTwaWU0vMzNyUYcouFC4OA6mCQUatUoDqYI2XTzCmmOhXA3lxJdiRm
q44h4/9ssaq3RvA1A7WoAkoyurrjm18w/SmOqWNm6nkGH/RrBRaBj5vdEofbxCB9
Y8riwnWkPqrrsSspfeIvTXUwU+Oq0B8LLhIz6ap6Lq70Y1168s7Qy1ZaWfETsB7R
YuZ8bdbj0y6rlqCPALvox1OZdT/Shzwzc8N5ha9SBfv2nEhfmauS5YRA+IlCqbM8
aI7UhkIpJhImgIjto0R8JHPWer6V7GKe4Vp381lflf4qWCcO5fk6C+EPBvEfHaRq
37vdJ+xZo9J3NH839SRMcCM9V00W9n4jIrg4dg0ZUPUeDDHUe9AkDvfQ7yWiGrNl
90j2eff3rH4N1KYysGIb0TIQYn6Ftkd0k67HFNDuPt/SAMoAc3mE66DL5/8j3xf7
IBQ/avn3hPfmUOIOnMZuzsrYVIqCI8iId0LtbrfonTUD1Gt8NOccPNzoQeegqhp2
3hi3yu5OsnrF/MR3mHWThaH0cLUQpMM4OrleU2Q3rmwgZpViaC4425JuErU91ppc
7CgdSDkeedjww7fpqAHc9Lt1aQXWAKatpFb46qUO92V0+oJ1npNi/PldBZACUwvd
vSw3jP9uxvLTknci9rqUSVhdPIT+dpAKu6aBGrR24Gl1/f0ch8Z8TfNii/6d9AnJ
54Z91YC/UEANZZjpA6/dj9Z3jYMhXOJxbmZBi2eOFxbMRgnul9lW1EOcNcongy6Y
b9pJroEev/cKkt2JuKen1qrX4rQvIS4igNjxIEBIf4D85jW/a9pP6H9cD0lxAbX0
2BpU1zF3Hz12L2eI6szNcBASOa2wWUPxHczOegqNHkWn/5tJZ4ns8Je0LqxHkwSu
2JGILrm/9nncf+UjHF20ZYIdUkF5gag66lkS2Qfd2up068Gm/eA845juW3t2PSuU
4T0TDypXwMCBaSOpAW3pIffrDYk17tUl4niKM0D0awvxQA3UPPui1aahwD/DsPvg
X30lKLVY2iHCs60+6Pzit++jpEC3GP4I6gzcyoEMeGQ1udXsW8aX7W5wVuMRjYME
+CBA/BIgyjp7Z+h/XTQu9QS3A1wsa9FR2ms5hSh8JHOYFv4EIpqWL4Y48FVZ8Uo5
0XeSyu1GSg44rouwpmE5yOuN4Dy5b0juTPqMlBj5OtvutdMDT7gSvUVHkKLZdSxK
AKy99YzQJS0a5iGp5fQROCKJmmi4E5TcYaJVfeCsTuLfDNpVmOoj3yoBhtPeSJyd
0rS/1uhTpXKfQ5kbBi8k0rZ1XTtGPvzXZ219YqabwjDd0dRrHmTQQCR1C76VFs8S
cE/E2hwohRdSZuzhM1OyK5XIv20MvM8WtXJNFDV7Yq8hjPCoaM/PKh/ndy0YVul3
TSvkd/uEoJ3pOQDE0Zn9gvrdkA7JnxkJq9MLI1ziM/RuEKfB7jeH5vW+psP4FAvc
WijxHtcT/KlbKIi5/UJ3h9HcpcX597sIEQjFGLXJO66Evsf1lycgqHdkzx5lpA+A
8MajzBtQ8OXXsRGNXlhPdhDOcDBwPudXChP0/LLbYHHgHC/HG+q9bVrItQ++5+Dv
zMNm/ZO1vr+P9ZcCkJDVEnIW9JZxHdplUxMY1K1z+f6cThZpFUUpUNYUp9YghCl6
G8yKbAOk0YVULfkgH092cK/W5lesl+QM/NClXyn8UDMsHb1gXOyaiU/qj7jLQlIw
E35dIpcfZHXHvX9Zl9oCf/ZH5x7ml2ESFCbHDpQFC7IlUQ+HVYgf6JhVMINSd6U0
y2LYtWQ3qg+c2ewaLrVRVi7N0DRksTFTYVuiCKf5E0/iplxuzJBxWnp8ZsGrEj7t
kxRblyz+TEY9IJuP/d7v0WF9EYRg6pDHKvHlh1cP6T2Jt2i4bhTi9zh5RmLTYnt6
rMUo8XsBJZS/5EtWivFBazkJDnxOroKAYEJ16dK0Lhn4YFmtl/F310cOLGgebP+t
9Xo5E5XTS3oJgc3cdwZZeinGXgc2bs4nBygR7yWAHycq0uBh72nl4j9kCFqZmrMb
ZkN6G3YzoxlPmB2Sps+/kzKFAJwBRfRlKXlgJ1UHoSDEf0PZ/jSlMXponlK8lG1M
27ioemdqk+LvQBqyajOrBS6KBusB3mkDAuFXrMnyFPS0913/X/J5Y2bNnIWYKf+U
2iUJ28KCnmuMfC/ayNdUCOSxsZ7PEtXmmwdkxjyLeIK7V0sqegX+tGlgDIYerEZ8
lBPiZSmDjk5NqtkDtp6gZmADNT2vrzc1ZOpu1B0CLyr3YLekBjmWjiS7C0S/gUNd
aV0ln9R5jAInKgFzU39vhrODd/NIqBhAgoTwBbPInTGf8xZ7ERU52ETjDXNB72Mw
xYXOHMkcqWlG1FKizpZPJ3XlfZcI4HV8mwPV3Y/poEaZvluKb9Tog7rdiwlPMAyo
lltwYOIZZjnns7t/7ZkTJPtYd28fWZ5VR131r1HCSV5acG8p+P59bTxRb8b2dg8z
lD3Ijy3JqUOGakx9iuSnl3yhVgp1McU83QPboNLytVzaoUGK3s1z8M0cACOHRxrf
8H+CKH/x/7DkU+X9Oup6OhvAI5809ywSXki9kWfauPbO4/LuW2FU92ji8dm+cxVE
o3gylqMWgnApkaQ2/w+p5EABM4A5ZJs/w0hjOMPLJ1zIlNSa7GB8Ukb6090gswfR
jITrAPGy7qwAHUGkOPs+vlHpOGfBSZlQ02eOZ3xxRaZ+3YrDSgBxlnEu8iozVl1k
yTfoKDfg7Y/e/amh7BHcHChOChRCka+uo+aG+B0VFh8=
`pragma protect end_protected
