`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
iJbGtuFxJpqQowlXSap9DSh+qTvhqOCVwtsr1RwwtMpBUQDCw5MKDjfSN+M/ueu5
2JiasDCBPtnrjPiv8eZNcuF4uM49lDrOLE/MWFdWsoPxnzZFEwyWhdQLS9HMphEo
34JMtYI5a1dYILKVQcn7m2v9XCqbbXEVGJeYNSd1ZNQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
PNhVEIZHAFs7yBeEj2xCiKEvhACVVAV5T8QqhvOfO5azmoWM8X7vzHbjZYMT1Djq
SOcCPftYNvy2ktEWjEUYf1o6kQXP/ErTyEDbPN2v9jZ0QygmKcfuhdQrOZ+FGEx1
EptmymiTRnjw01ZnoBztvnHKzDUIkdyFqKgDpDy/RmAL11spH9536Hl2V9Scmrth
D01wuOaA57AP/0+6DLWDjTinBT95QlBbscr76PY+n5+JIQzCcSfGl2qJ3xDEES0T
hG6kE+zCKbS+nArwISQhMqPgYzvUYtOw2JrcEn+WPBWFv1MByh3MZAbCh46ifuDJ
3nuA/zFn1GsAlejWY88ODgedcnWg3CWI6GZTATq4eKzO4y1ASP8v5GEmZm3oWgBH
wtDMwIhOmBLWm38URrWZO0lZIgCoAJYQCk5Fb8OakePxfi8RtVGA11RMX1/7wLGJ
u02ccvTsWLnneF0ZVD1AXsmYt7S/2Kg7/V8I+ZzCvXoyH74zeuI1eTlFPaV2kQLn
yHZcjkF1lC9VQDhVn8vEYMreIW8E4oEt3rjscmanZxgszw6TMkJS4dSrYeNa9nhe
OjnekuwsAB2w1WU5kaG5juWoDdUDqkj0Xg6DiDQMUgN8WAxJkREnuC3/qEs5yHpp
2LKPRoPmw7HUK9UthdPk3mNB9QgE28xrpOGbWUvpbHCY2Q81U2t3K3a4mRp2pppi
WCJoaO72S1XjoV0d3pEo9PFw6S1xCImqIlIFIWS9H4oPi5jwUtGCFSK0BBv0Uqdh
aR2g+iWydNyx7l5Q1EgbMxFohzBC0Bz4vTRsZy5i+4Ez+x6VQGDvpeCmMGVLdyk2
br6RZB2NFkh0VqfWzkFXrJMJZM9AlHhARth0Oq2E+pjDvcW5V9Q40y98ubeOJWst
jCHq8pGXwfRmwvuzggkgHBlRRbb0+rtr1cYWxBlZD90aMism7JBs24u0POK6sat4
NiGdqcF7c5+8se422PStI47OOEVz22l3JifPWq/GHp0T9x4vjUrkhRaOrHdkZm/V
el8wZ+kNaaTXnlmceVpoeoMP3hPy3tIWWbyT43Rim5Jggyp/9YITC3ktTggFiUBb
bZAex5ygklcY3Gt7UoSypS8lEeCv14xEsVMSBeBqNNMpUAj6lJgu1q2JqBaaXKD+
rGmzWcGiE2/2rJyPIf1krMaG0grtTWAyuBQBkaI6YyivtxByD7iJY+hckw+ygCuq
wzMTAM5jM7WGoJUr9T8EKKb5E4lx9T0M+C4gwZ6X45RENG0tVzE1g25Z+nj05Nwd
JzcoPMZpovPkezJjunPD5m9pW/PLDuSiHNiu5fwQ+j4t0d5otHG2foN4omrjaiaY
ZadvUi67zAigqEM0iWIn4B32dN9Wcl4byarHHn3Ri6ZEdfUlyOk+WKR7sRD96voh
8YrjpOsDzjhxx3OnmnQ5nKpoX9YCtD2km8U0tX9zgdVcX1J6va68F/XbL10QUVmH
gCJ8b8z/wz/6UNnpXqU9FsJAjMDLNXILzVSrp+Qye2Zrc8hiu1DmFfTPB+jpgH9q
ssCG2mdJNC+Hi/TVCB8DLIimDYRuykN53w1x6DLcvG+ElJKnXFFKrRXBsjnBj3mK
SyVaerFpmlRiTLyeOnkjjvmjiiVnzbBXVQGslg396GjLx6eq/1ef2MaBtrc617R/
TFcxtc0VP8+VbVgSvalrKKQyQzTwbxD9Z9BSw3MpAvF0HoTjTpT6ouBa09Wipm4Z
ArnnegNu/YNS2YD1dcFnPbBhLFg0vmpU+fo4LvNiWhHx14TBzno7vUFCDWCC1mhx
CMrXUBxfJMHg8QRF2X6zsJZIMh/9saMh2JoN9mYX+8adrQptizhgkXg2cc20raPB
/CIWS+DbJ0hRFy2DVUOEpUdaJnLDzxkiW2dTer7OyHtVsSuoz6vvp/sQIi2K3ENE
FgfIq+CKMEr1Qc5XdZ5FQKdafimIICA+FSvX1vafvDUtJCEIZgWDnQL4Dz3n5Uhd
/rFK5MBPbwplRj9VgRPl1igl/dp7E0gyclayMBOwMbyWYXP+GfGxPf5WMAZ5U06j
o5ueb2h2aILzjRujR7icD1NCNGcwSt4k8fSaPGUvIWhvCaiccVMbgUVpj8L/I4wD
YRW7OeQcmzDG4/W7mCmJkIw0/tI3ODsM5YZVugV7HR+yXoNCjI62af5+04z0p/Sl
dsAB8qKoT4z1fBB7tPeozstiwf1A7zTTvbMCfL6Mx8BRmk8gHnnqswTa5o+V0PQ8
2SBbwk040fhwb2qKIu04c0FgB+GhxmgQa0zUHfUCCD1z8wiA3878jMEwB86SG2DL
NqqQf4ul8tNuxzh0qJPysbHDPS1hApG3oDaZzcyxuV+E6pxPvd1y7v9C67+30mTu
t58fHluKmY014Lo29h6voJh63kZQX7/5/LrvzK8hQqOmJWZyWYFMg14j/kiWgsyS
xltPr2ZLT4BgBrgW1UuOLkiCLA9DnsE7i/N+0hjiIDPbFdgaQnEmu3s/mGJ3GJbz
3alNhuNpxXaDD8SocO4pL/D7I9BzmyPBHnr/mYNi2Jg2eaIsU1ok2oxUUn0wVtBJ
6mYV+O1UAbs5Ww2ddnKkNCKCg8r1vFO4V28se4sou7WqvRIrKkhZ4TxyXqWIqzAY
aOTZMJ+/ciMKnamiiUP5uVHTowDDgrjpq2WNdsMXQxxsNCCGtgENAbGcHKWDp5eE
NX3UoCqEiB/KhkM+VANfVlcnKXo5CtHU6sy1Q5D4iDStil9I6N1ZCKF4iPfUzPOX
X/kzchRaJPjvyT4+OGsf+7p7+GNJc3566XyKg2vMISW17u9mAN1l8/3xvzM2h3qD
fDoZLqxsBf6OysxswKYILthDj34fU1LvZwM5dwAOYTH5Mk6wXe2mI/DoPaTTlIJb
HClKuD5n5I2Y5bna1oLZVE2PEwPTteb9RAVAT/vs3TWKSRdJBxZrZ89h+0bkzsS+
LRWKdwCeHWC74P2yBF+k/B5bfIHrHHwUFfYecCP4WAIORC+0sk5lyt4NSJ8QgVYT
xi1P6T5KbTxvjJRywaOFRGxnwrhJZzIruFxnvkelUGTm52gw580juSfhDL87z/X1
5M6N1KOR5msd8C9SaNCHlgG+w8gzoBeJ6DcSNFD95dqty0zpkGaWIdPfsA4wG203
QTpT8JRUJHFKoizrad4Pt0clL4a+xOAgY++g/RyyYCu+8bnimalpqft/liSrSrsF
DkA7Udt8GSJFhgsNMqsjT42QitsxFh51LH8HNFCnikzHNIzaMqoqxD/ioqsbJoJY
OjONF1C3bvTevR2qk64rxU+Kzi+X2IXTzTUr+SXvaRPA6bYpTgMm0OdNM/gChm5P
TPwmRIPGHVOAU4Z+TecGtx3q+RRodu0dEyKnEOVSmfdgkuQHUdLbtV01oXoqrhL5
JWQ6HziZ5EgTWGZfCGt9seumC0Z4rbuVx2antPIuXH/v2McCvxtAvE8UujUEQEK8
6GDW+zfGIhE2UnzmOo5DRKipMXgFI3xUa+Dntw34wThhlRGpY7n5A2sFvt1L8qnT
USweapZVfy5O5vBsGnwgdMR9ZKXg1UXpOoaQdQAsSQ0Uf2B6WraxZfXxYCRz56eh
AeZx5MYqiVKthHVVex94Iugp6ezQISo4t4fNHWF/YE+erjKjllIvWzt07A2NBgVu
RLPiL68tB5rS31Y4enHcV6LsnehOZZrJvA3iaRC2I8EWGBHMzV5GQr6eEWue0YEb
K3NpmJwhpZB5/kN50E7yCViwbU43gSD84vL8L69PLjdrtV10HW95Qx/upd8ZfxXv
NdB8ZRcyCYCMzh5H69pEZaErpUScewe4dOdpPC/ky2EVHD1jPzyfhY4UNt/8t/e/
3cFQjHUFKfsCNXCLT8MjyXW+xHOHb1bU6QBRBsTISwPlEFVlEiVqS6Z87Zj+0et/
Rvg6XvxkZ/0sm1M7lGPldGgq9AwP/VbM4h5eRJtYxfKkFG45Z2pVozS0Cyiq5k9J
bVT4eVafNcYUP6aDSK6PAyDHHcalh49G7yr95fM3a8dbOMwoVYp36OQz3QIg/gMl
L8DPeK4RWMP5h27UKoAXA7Tlo6b2IbxBTiZd0es7frFRPvIacArAseqAa7hxHDET
8z+3kdV2O/4LvLZYhKHuxrZqPoQetWVq2nm0NoOYddiIemRA+f5tfaR26we4tI7h
7VrFXa3wlvlfjTrD7RoNIrjomOHmABzQ9HYz2ma3rh+m7bvZErYmtRUD9UMWALKM
H8gJsJb3GCJarUMrWXQPwygmLCjxgVlx81TVW2yFN97U96+67170wKD1XNtK8+by
W0/h7r6AZ5IMY8BYHbMk4PtiENRDP3HGW9W/yNSmtnu/zchqaHr4MXWyvY2Awwd2
hn6ZrsEkz6Qfk/HxA8qtiIWs7q9M+9hJHJzfj/rMNWRXBvxUpBmNCTuliHRiYGv0
qFmr4WDrLruSDkGjflbcS2C4CjIAUP4s2AeOBmhSEhd/8RUFRtJ6qwMbD1gNonzC
hANuKpjDQPCkzDCvw9YKvNvJ86uvjLGxxZ/NziLm9zdl+7PW1JaIKpZLHk1aQjcJ
weRcXb54NC9oKFIxiEx/KGmW4pjrxqDU2Z3NZubERNU40kmxrK1vRvFO0n8nEYQg
kj+RWcwQNcEmOe20hfDTuK0U7pjts0POmY5BFWHTnQlMCdizb9t1EqBXBZ0gOvWl
U7xYo+RlQdtlzIuUZ+UbnoSSFJKqxP2BRf3pJgwv8LaNjfRW/gxfXCsAJ2aqZI51
8Mi5/+/8EUHtWTHB/G84/6mfCPuPWiRrhTWwbJr4IOaj4Wpa0MpqUWw4GzsN+tGi
0svc1i2+Vwoy+YS6ldBZMyS8P0qbs3oEf10S0VD5EWDDD7W/YdgZyhGcwd2HJPq8
VrELpefHdEL+DOqdMvWCczr156S/3WyAcqsZgSy85JOBUvK46jy6StwG2cNd7sqs
xvBPupKh1AtuiPtJtAvW35w9pzplM2ecda0/YCgLs/EhkOHkPX0CUR27jhH4mocr
ClvqOc0IqjYVHoKLPmG/djFX1BfNp25AmJJ7d7UX6vi8OdJoNsguVYsFVRBGbcnN
UUah7uAMYLLYvRRO7YY6bRZTsw9MUzOoA+saiqrAGUN0L+ORGrSi0W2tuTyGoDex
yU6kFS1DSCY7/yEPtUffl0m1D58RUQST6m4qBmkUH76XtoIsnafgvErBCoBT+XEH
2srgPoUwtXlx3fBURy0Stlp5rjb++HYtpiWAS23Zww421EDzQkDu1+yZT0xrYB9Z
PQ0Moe5YjFUOQCJ0xYYuoJyasQ2bxdJ9OCCZCzOmK+9RD1Zs/7OML6MzsMDJWsiI
2O8VK13UY79abaUBgB/44j1J5b+nduZ5L2zdPjH63n3QzLZdxnIXhmQdyLaRV+fa
r88fHsn3jmjaYbFtgmO0Enfyb9DROBE86k+QkTvFoGImRRtvkzCZsRfAw4d3vz2m
EYhX5OQuVhORm/Ph6G7p1JlojE5Cjk3hLyrguffJiClTczRfVhfKdsXuvILmisFs
qMRInByIWyz7nJdk17mP5Lkb5Rs6ApVEsEWLgceU87ucvOheJvbEL+H4SPnKaRZ3
XsKn9BpPSveXCY4O5posmbAvvnx4hTg+/akrEn3d0rMSaJMOmTffEy103jPJ3WME
iES648V8KLX9i0M9TTsdl6qzQAoqGp2Vg/BMd8nkiwwc/Ectv2Owboco76tzmVr8
k4PonmEgKrQc2NvKgHb8X5gd4fT5E2AHVcQs0Qb6DvmmL+eZ+gnH61sUgOT9n2ip
KIuxjnDXUx02aZ7hwDEmFlfnrRPAcATT8CFZpOOpl6ZBHY9W4+X5GW7Zsv+yKUH/
wrJzQETGplUeuSPLJ/I3r12t97MkhDUhVveyvFRUmYpTj499eG78dzwWUuhdYRH4
phC4G55QS4BctmPa9vNH0QtyVHu21sdn++y0dntMSEhol6jk9TJODJreZ34e9OLi
jIT08A7+qY6AM+HaxEhn1G4IhIzqImmjvyRlfBMgU09kuy3yfOO3vonfEiGJtfa7
CjtDDEd1KfOtayC8dypVA3mhDLCUJTZO3QW6TJB2IM9kFSsHlGrr4ILQedbDqCG5
kqTahX+QcYYll1/qwKw0qVnC8nQNkJF9Asp0/opuWQgUFShGXlADJu58Ixyz/8I5
e78MeMycPC74QC/hAB+ZQ07KRqYW6WbIPFaCdfWlcE5sMY+v5BW5HRPvZWyUhoZb
Jl/q0mjT3m5YdVb7ZWslwpJ/LeP6Iu0gAwAQoNvRD8KHqFRqdhnkubxvlaUTp9hE
1yLeuGmMiaL4UF8NkRQkTW0tEoRg7YHjE7dtfrGJRPmwyCZZ7eb9zzw+eoUhEqV8
lh9kKgpmNlD34tAh6ANpZiU02T2HhjFA8j736nSATNb0ASmnqH30Wv76z9ZSpUYi
DXxIT921PtzqG1zP/AyK6QQtbayF5eTk9+mxdG6hfO4rmvcm59oJDrLh6bMY8vKK
KcO1p1Tlibjgy7xqOwokMg1vNEJTubbBRuW4hkt3zh6VDgjtUPlrkxAdliybkX5h
uW1XEdKUuxBW7oyTYOj1HZ7ij22O0fyabxtGBZMbF0FI8lQNu2puKIyxapqD/s5w
fvGv1+7TUFe7+oWgzQeQxxot65Vhxj7pYN0u9pVczj/MkAgvJJ9Tx+SWAmHMplue
3gMSxttTi8PUPW9QiMni5vyGtHe1iy3MbfVprYAs1sfdid/gS+yfAGNgJM11g+hR
JIqmIfiv7i5U9GmxKxAw4RF36w4eGaBhkvHODOMPOQefGMwxZE11QSBN6v4JYqE8
H5Qe3cx4QKPaDU93hqJfgeO0A9cRrSwGVsJsvq0lkW1eR7yI2L7OFAosOdNbUP7+
reW7WHRSj85RFGIE5sIJWHaLvzl983Tp0iG7Aqmh/0U6Yhw9p2AFxTmRuMDEtvo5
i6cGY5GZXBDI4NoK6pH5cvV3+NELq0BZetG14oLL44/UovM33uMKyQaCDDggydIF
JfGCH7KgwcDGCwS9pVQkSN6EV/RBLXmcb4xR9KJaRwdp20w9mfc2jnW+o6NdHjPD
XgnSmvaZACFUp1je9yJHR48/fYHtnni4EtsRVfdAsZb/z3bIxAXEB8eYqME1/t9u
FSybcVUiPf8TRYReZ7yB3AkZiuurapK4ItUOyQSmfz1LdLk+Yi3qqU6k/bvYpXDQ
2w43fL2cNobsV83n9TPiLo0GCNmxfS2Awx1KGnoKhyYtV/HRujR3JbUf8ziuWg7V
Un2vCFrp2QaMq9ajp//p/7iy9HlZugLmsNZ8htGLnMMHy5G+X2BsZyPFr4jXp6Z0
Y8uJ/inbz+57QBP/XWX+7QSveCk+ETzFQuVZl/79lZKGYMf1dhJXp4HV97DUe1+U
Comsmq/5PkX7QZBzIMmVIcfV388pyeXEHwXPHoUheqIafTECt0lKbiJ0WiQnl21q
kvaxOj+ncGGu5SLc/YJWf0LJ2lhH52nl8mWWejav8fkaOJQfQjwQ9SIAJFv/dS1C
kHOAm3jYwkrqSHgNK1qgAuvyt+M8rbmuT2LY2P2kj8pw8WV67nr8kFBnSC4PDgzO
3n+KPribLEhgru6rpXKm4e0qBEmvYnQeN987bMwpeMAmDuzucihIx2UKu47kKtHl
xMmzYsreB/lvWjISs8C4aqVARqcE+aWGIV40r2K9L1qL1PZ/lgK9yRFP6x0uEhBj
oBD0lqdChFGSFPzWFeSGbHlgtDl3imgQXkNmxVb1pSIVms4jROXHdHADdrC3ugWq
HNC35ievLTO48+JWQeH6LANyDipN7F08gBVBNRHJ2SAinFJjsdpyHnh021hbztib
Xa1ke2Rvqy5wcVVEBZJ3cbyoP736VSqJ3DW4/rqcsmNMZhPS7awqN7MQPNmPlaaI
23zPTKgcrZPjgcuKZTIgEWXd+DylZfiORo70PCM8nLhX9a08OTMIGM1bSy9tnFzm
fibsG6IE3E1AcxwrzxQE2zcQkYq7G3dcoB7BjWHZR5/hHbSVMGGDQB5mZCv7facN
aR+dUZDt2F4t6KfTt5323zl5AgMRhtx64PRbCom5REjuf49MhJMk4oJxjv4qGdQ6
cqPUu6fXBUHBCAQKctkoUObN85kMs4Zzk7UUblEuEkdveHI0waiMVgFV78X+6ubG
NDtJq5zaNvxNpxcbfEujWxmXiXb1rsP4lIItIooxYA189nJqE+6D2Ql3U7za/uH5
OY4zFO1m9Z5aZ/GIOlIngAE6vwKucqgzKN48EaK85+BX15FDziIxHjsc3uJHBGuO
a39sUJ4Wasru6cm4CnQug4fMxEpF9cxMPjyQHm5ssA8iUnu7Wexc/lkpmMOhFfWe
AcCh3o1oV5qnpfpBoMstXAc5KNsZeZBjwp4VPv++zQCerLluE2vtWtT24d5eluW/
CdnEnYRgxRIr9vQ7XIKi8B/RV1ZYxqZj3Iw/SNkgEPIL3XMvYiOP2xEQYcDxDTVW
4zc/942n8UW/KSdl0gWH0RuGjdFIlkfOFtITuRa0Cf8uyIJLrAvQP05UN3BEQm7K
diH7iPhR/ZAl4dDc+WBf5s1VyrEfkWeumz4OgnflTB9XDx61a87TMvD1rzaw4LVl
1ZFjqauCb6qJxIvJhEhsHD3oj4z7RecyUtw+wj6HRPWnh9clTTsCj9IqNm5D2BU0
HrlFdsJi7FCDvPX6rlpXHqQQ/pidSuWtEwxKHJp06lEl9wfODPwFbhGXulB7fwgP
c+cHj6tUbR3A1kyIyR44vs1LDK5nTYIYCI1YKvo5tw8hcMvCkDmHWkzS7hPj2kPn
uk7dOPBCbZ93NiZZ5aJKVyxe7QH8dAQmJCr98s/tYtZvw8/Gqc6ZzE0/j2UphzDd
56grrVJmgS3DXsbQ6TOrOvKt3gJUYSWkCfG8MDScqon2pjGrJVI5iBWv4FpP1zCl
4GgCia6BYvi1CoNSXApWRYGM26bWBifhCenIRUVgjMog/fnIKtWMELUm7m3eWGOk
xTpFH0dfp7b+KjNaxR20z7c3oKToGiZyFmfpe6KEum3iWWBlPvk9UqXpKPIDiB+M
P+RPJcjZWFHhWGu1K47xTnCV6giLlYSeRzAYa/NwIYMqpxqRHTIwMCilYs2DtyVX
KxbebabRv3SLHfwTtx77dMVuufOgcyMRcDOm7Hoialj4eZsUcOTcuuM9FbCiAFn9
WfJhCzf3opujmmLlQpzBCeCqLZlqW9MzyzOWGmIXAmN16k0FA/DzouV6g156pdlb
vK+BxwFjC0MmFEJ/CV5TrmT+VFJZP7zV4IFubnmb8JYAgBbrodv4pbZ385iB9A1s
HrakuGQV7FE+FOGl7mafeJaExWDiQhZ+9KXOpwZFlMytcMWDbhnaircmWM0X8/8W
UfVxik4grznMTRr+pM89KlVT6/7l2KfHOxXpnRNPG3nAMcpLdVs1E2P4WJsNxX4w
j8vE1JQQkh+c2JsQQqBBDXDma/9pqLrtQEfBQIURAEWlgxjP1t9P/7oxt83sAWek
5ka2NYO3YrxfId0/3EyAo1jlv/PtXKXBgC7xQb/6JLgI7ODOxhCVx1dw0RKJ37+h
lWOaAOhgCUyxuOFOT5/OVV37M24QLXqE2McZryWPowzaAYpLormgdQU5doO8OlNj
SPj7lXshkNzLOk07l33nV+y4HFrBrp7W4lnOcTCN6Pbxsc6VFNZcfCIICCe2lx41
ylFs81E2tXquBlOZYZ+VNhhvqKHJSORfoAixUNE884xusU7wlVM5QI/iPQ8wgooX
gcJ9v6r7+OoHRnX8aseGu6P1b2yunZ7F03k50AQG5i5PecOcawjuVwraTx4M3PKh
5GTRKIdxolr1HqKQClwh4RbWAn+l47ilQTNRKxvZ4U2+CmAigWKj5WJ1t5OHqF4z
dyp3btkXLLCQ4bbBrZN6mVMIu9UyTaneuK3fE8/fZAkJxnxljpWkDZMXYHjvDa14
S7lKJIlXpqA0Y2awj45AoiNUCP+apCucLfHD0Es0fEMLsFVPShZ7uVCnmDIdF7tQ
dw/aRMBwaSau7iWEW8NqTA7TeRe50LD7BXRe/CayIpJs2F2LYAuFCfErilwdJoop
VGke8oAhzn1sF+JlD1eLLUb/hnxeC3VEPQHiclvByQMZT/TKRJlkYL2nTs7kzmgb
4lw6ZOub5/R//W7YdNwGTQXDs1hQA5LFHveYny1+i3eKam9Sr4glZX0vGHkwzLZZ
8KPo0RXyVexhMzYduSJaRAxChIpcO1ZnVk2mlzolo9rBpHt1ziKcIdIpFEuKc/cT
/H6sCr8zU/YpRkoGepxQZ9dKtnlR5XKaCs4psV20K6r9avSCPHUKPZe5iYZfNSMv
tHjcy3sI1OKjuEf6BHS8XUQYfC9xO+ta2VjF/6WJG2N4ROmEU7STjTeyWLZOXBsw
WZrYFbyGi285y5Bgnl29+s6RFVWhmc9P56dKEXBqr5dvPbLbCz8i+OrRQBlDnPWl
hW3m/OQqgUhVfMlZ4F0u9RH8qNaflbwlUrUEBwRMqNRKBKLtjcorbnm5ueY7iYgN
PyY2Ekvs8aS/sO7mWAnh1Uasroy0SbsfVbjSsAirBz1mtj/JTtD2B/3qPadBFQYO
Xp85QQh/g3IkxlD+0mHxr36NYaV/J/P/9tSOKQtQEi+/TNds1wVHhHTYQeERYWz0
kXLyk6JDdTgEs8V0gOwMf74jzRCEiBUzFraPPfbP5g6I81tDCmRgbn5/UBo7IUUW
ALf2WXFALr+c9OplZm5xsgUkoj7d/eO+AKh7v8T6ExG2WQHvP6O5bBGGUyLbefge
yx6/cpYI5Amz6gCN1LDkUZqK8KRiJsJFBgAdNX+D2qJzkCY5iA+upClO6DH1rP19
T/H7jtKP+3iJ4tpRNe9RBIOSyCT7lFMQL2UqJ3Au/he5hrrK1Tn2Qnw9HrVq7mvQ
2Y5AbBNsVPNPv4F6+afSGIHdC3bDVoiZoTHM2H4oRfpA1O4ti19JNl96fsrOSl07
SpZ308931SANaL+/QRmardNcsgvUpiCxJ41NZn80j/JwF0x6G6ij5V58cxk4mI65
+Jm0cUFC2wwbLd7kmMUNTRV/RqLEHeP7ExsbOBZEDkYq748aX2JcOUsW8kidIQVk
RHXU/9VUI7yK0NIL1vLwDEEbgnVBkNdsgVDM3sYCIHFcM5bVdLM9PbSfxh/YhhEO
MI9Y+Acm7f7fXMZuLROy2mv+F+wtSL5EqSZd2Uo170Pxubemy+Wt47QOE1iAn6fS
0zrxMVxhfP1w3adJt6IcZV33WgAg4Ym/Yqm0tgfy1JbnDxrY42wVnMLhjkK1tvEQ
2enOwJSy92UzXuBd7wDhqxXundd5XKnh1buarHDh12OqLuL8hxqe1kl0vtgH8eV+
BxrGfg0hrLpzrV4E8TBM4+AF34vteg5Nn7im92rA0O9XP0PKCSAPtnhpzMs3AqkZ
1noxQKIVEKVbNGX/nOyA3IXpGWwCnIBWHOvXhGa6cZk=
`pragma protect end_protected
