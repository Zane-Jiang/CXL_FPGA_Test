// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
cCdJd44snE+Owb0rfn+wmQGFAWJTOh3ZpBYmkINycyTj8zzvVN9pbmoK8KWJKzr6
zB4im+D6yLCGm9p3lI6e9B++fOsJ1YVWrPNetJ/X1ngzrMt3XqPTKIIhO69+4jK7
8M+7+JS9ys9/iNBxFuVUBuZ+ylqLpHRiCK0tBKQnGG4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10864 )
`pragma protect data_block
c59Ph7d5aorhTvTSGoMvqLyve841MQltOsrsd1jWNeIvl9pvE9QDFxCnMc/SEvP6
LHfKUHMAduu/7u3zjsCrfyx3qXVK1j+vcKV6xGSPmJXgw4G0TF+17JpNid5SmVu3
IjCe8LkAwJWIiRjlJD4r9NzijtcxNlnstsK7yc5WvqZJdxSpriIlnWt00G2vPJqc
9PbtPVlefWwh/YIg4nxFZDMevOvoe+NSncdqdVq/Ps9/ZrwVoyJ6uKkxkrTk2dQJ
LbIMlquBYTm+Xibgk9cQSqzlE3l9x6AuWQZ/wRnYAxQ73pNIBMQsUb1hw+njR3Rc
YBL7r1B6dc03LTjYOE0QkZiBuiwuPVm+Zby+Uqe1MnYq6nC18Prr/yYnhkE3reTn
Llfix1o1dYtmDfs+luhgyIgcMxT7VDoU86Ukbba9WuJecqAzDG5JVv/duTWAv/Sh
wZSOYTw7uRxMT6iijtiDPc9zKcMLDljFq5TN3T/XAwnCleNZfFVg/W4D248vi8l8
yV/z34qXn2ujAFowcbnj2LWVJUUYAh9f02s/+Ri/X1uvuwmHnmLB8Kg+clsF1w0A
zLwwOSo1RvWeKFz6VmhMe0/1qChpcCqVd1Hw3w9K9LCZWv7s+JyOeO2cMEIIwKWq
UMLMkYE89zSD7Yl7Qv0ASg4HkKYnKDRT/qyWlLl0C69juh6BXk8W1q0dXtYqcCvL
BV1YqA4uTOAIB3IcKVX1REsirBKSF+KRmf3Ed5yV9xnKC8N7kjKLijGMFmnhPY8L
hgnGTIUkOufAioC+J4gQMhwKlAqNw2frvUHVgZQsoKFt2Yz6XbfVrvkixJwYmSpY
1IA7VDgHLj9wpcMj/qMjptghzXYG4tf7oJ5C221jkngoMDgZoAUDPvwSYUH7UhNc
0S1PmsToB4pmJZr1T7BPFNkvFFUz6ufLfmRQkYHGkHX5NLg+ED3eCggKJdmFqLLG
cvn5T9OigLyb5fa3o01xvJiwSdn1K7Z/cZSMMBUI3zKLIB4Wzgl7SH5Jm4cLJNsu
LNadzO4WBoBS/2P7vEvOeTZ+PGBXG8hET02ScrefZabhAkIv2IsJfkcEQcp06Kwn
pDYVmOV3ujVObTSNE8BwfLcw+NSr3AwvvjGzM1EmZONSDRhwonP2YH7lGGNjiXiG
h2wKVuto68hFPHRWEU0kOAaDc+6R2qBf/cmBsLRSmjLzttmWkufu/pyCj7QZfZ6c
9veVpDmmWGHqiCx9WUB++LPwTt9mib5TDZINEMBtYoesn8qcf3rzw25MIZkzXtk2
nk5Cz9S3OmoML+kZvb6QHlevQKOZ17lln8twqdZRRih1vj84yx3OwaF0oyS29Fu5
J1SrWbBWO0ZtaxkGjPGZpOJWPQRvtuXQ0VJaAfdFrxju8k9VdgT1qBT49cp5t8fV
yi851TzeAZVyEu0YBfSkRTpl9EzqFtZln6keiBX2XtH4/o/f8dNoq2WotnA8LFDs
Wc3Azt3EdVgsaxYqtxJsDUaVWsMNwBaND5saZ71ynxONShSkv9jBgVor85Z3fRdE
nxmFVpz6+YVTxvKae4fx6rz5/3FMb34G9Vi3axH49NZQl1jke61RmdRrlXT7Dz1d
JkFO9ZDSTGp9camLYpnTW30zNmg574QNVFYPFWUvEcbvFTyK+m26IrbG/+Mw/T+V
wUQAYKtE86MEUXC/l6Q1yHhfTOTLysSFRtXYS3AxteQPCER0QUOtmYwcJXfz6aDr
VqGE1Qs041d2jC8EexmzR5k4AUHbpAJTq+MGImmSCu3OrbstyFubEgmOpcsmNn8c
tx+dfzPYHhdhySuzuf2Zepo4k1IgDocZFKEXnwAAjBJW9aSLeUTO6jgVFvJHYsX/
dUf55mJO/wAZ8tjvOCtKcpwx1n1CfgW6y4Pjrjg1DrJOcL6qiANQrStEfUiCFuRC
HgSEQOXYB8ynIfnmc6lRNejbALUMVzajjAokT4NxakdrkHsw2cj1WLu/F+EEuNUS
+FXN6mfsa6Go0Pfqjlz5R296sdvJXJWrDIAFIAoetw5ZTC0q3Dy+slTDBMSzGauk
DhbEnuRvS02PfEqGPVOV5iIwW8XfhKv64inCQEeyFplgHahxc+DfoRAtzQK4ihp3
hsGRvWXobg0XLfn8ufBTsShcFwCH3fZh8X+g1Nj8LO7Mvgcleb40A+EPhop6Kwls
gFRONpmy8YW12GV7TBW1o3M2IHrJ03cqh7UBJjmLT3lALXn9NI/zdOUn5Xqm5AVl
ooLsczyNYTFZyN6yu2dEpl8kxxbeQVnFYA4/scUhp/+FcUhpQgIHMAgGN5rvhIJ8
/rr4YlhDcNP6O/TwnAnTLq+UOJYvPJDQ4TC8gvuIWEK9ug+jgBHP1YKZW9WX3NmL
ECBN9mcaVGHB0sJGUBcfhcophyOSQvjwWzONdaD2ABeheupXJjBJYwdIZdFEywZj
3kdQ8xG9u4jYbQ3LsoHrYWokFKB4klSiw64wiAPWrh/46EwHGWUJkQEH5VtI3/Uo
Q8ZKil+67qZtUMdeq5mpw1lD7rTznPGhw5dmMjeW545NL0oMEmCZ71BtWnb5q35I
FPOw8qOJ+CnnK/ysmBqFJv8M5d17BImvNat1pHE7M/4cHXKAbIX50NVgRT0DCQ/P
xn2L1orlBXipdLW2P114sVd0bvLFBauiJwmao5BfsEjxmUZ4j+WYtdtXeOFCGgD5
jJOYkge23IE2frhSGGBAYYL4hKpiRk+thGOxxi9ECkuOdYfvfAAtJFttJsbWqQuD
8P/M7TFgjK3wYSe1RGuYrn+hYFL/yZIuxtp49LA28ERMbpAO8ZKE3k5iGdNHozrp
8BtBRNg41M9TWMa2AcYHiEItJ4Z5YsGFb1BPx9B68mvgo3kUrhVwA/6Qui+TPbcD
Xrv9Wj40b7WxKJOAygsfeABYp6BBA3Pqzoxl42trR0XQKmoZ3L6QjjsleidFcCB9
04yofoWlsRMAMEUKZAeDUO+KAwEuTsNCPPcoCcns3///fCHJ0zyMGfuw0m6wVBg/
NTgl7E6BjcbwcjnBlMkCN6LrxXVtX8QnDb6I/WbhQIFm+n5zs6VwJ9B/XnKWJJcY
gxiQ4jFQr5aGiCHJdJaUY7Uj7yTpoc7W6x4pG4sYo0+5InbRBlEXUfhv3neLVRXz
41TJjTLSFELxHO6z58C23riPSHRpLBTfHIo6XKak5JoddZX+1ulzq0FbCRs5Fjxc
0BAlFvMhA17QCRxPL7b8Lj9lgITp2K7iL2Ac5FbSuqOPlpN+f3yulO3WhGc2/xu5
dm2hbwZCP4bJuQlFY/eXXTHJOu7c9rUc1cpwu32mj5mOSuLCI5dWl1v6F+3EG6Sq
GOsJsOzvQ0eIMGchq7LJ2WrNrj0kUx5QXeN8bdLN9jARPO7/iuFb47dpIMeBvC4Z
mw3u8QNPsYKMvGITUPuNH0SxrqF9uxEGmrynD8aIcKKTIaqoURz5VEdN7gsz63PE
cSsqds6tjIeBbPeZkl+KSACFFf+na94kY977f9d2ADTdgSc+UCY4pXSXnOQ2+5OF
+8EsolCqKGj7z9DXPOfMJv9WW3MFbKjbfu6lyVGL3N7YBa22MaqjEN41jT1lKddx
Xi0cBf++tAtr+5UApKLBjdSulLnXI7oRthjK/6PnSxNeatt9Ot0KMuwkvp1FRs4C
4z/ybL8GyCD+lKmVrMWw3z//tqJhD2QSLIbEJnXzcfzFYD/3mFMI/05qJ08w8Mul
/z1DSAOkSasEbfIShvpB0iHwQRzvke3l5lP1heFu7ixfqm+iEAbDdj738YSG6eod
/P+OYdTXpik8JlLwuB7tT6lR5EGcoqxNsgffCf+xPyMpW3jKDG8mgZq1ScPtzdE0
4Rrmc8coIoyhWP48+tzWilfBzqWzEuSZS9qN9KrRB9fDG8ywetYXOeYvmqV7N+kg
j6mi6r10/mib5jj4i5ONd/zvDroriio6F5DWgFlIN2cetP0owj1F6rSFbBa2ZZ0Y
A1plyc/eRMPEuuxqYxcFZkfTEicw8V8r8BCPWencCobkj0qGlbKYmklbOvMtRumr
bZKCHGgQrdOUAjss22REQ3nyOU9gn1B9wpMsHHdJywW3TSUv7N3BonjR5JGQoJc5
2odMpA3X0DzNFYYgUbuajQmVMOVtoIMxAvIluOXN3/jRQGHpjuoFfjf47TQAlkj/
igOV5ueYj9Iw56PI7D788eYKtHwGGbbAj3YUNGj8uwByH+JHeRbVdvUxasezTlxK
W3+9EW4UIO+K4AgBiEDLBYT1LEEZKGD3E9DvzXZXyjDeJpxtVLP+zmNI0O4JI+2Y
WYyD3sFWy2J5Xz8k4oh6MLvIlnDsEIs+FgVdz1b9YZO99qJ+qaE78cblmGwCcfxj
U4tlXcvIGxESINXAam0ieX9Ron67ph4ul7LxFCsfZlidVuOBBajNTkKwY8RNT38D
VCZuLimZ+pIvEdhMgWlMk9rZGgH0gxt0FA/ukJtnwE/6/Bxgonk1jPBPn2JfB8Ec
JwepdTrMNkEuyxgO+ilimJychs9KSw8gNYBAO811TfynvwoAwjOkTEwbJZAg6uRl
J4BYTghQ9IbdmzLoTD62SbRabmFNOrh0CamazvJvx9b2YjuTqvRbf/kbn+ItnK5V
iNi7BWis0cD4dpcOjvMuF2yGeBo49e8bv15u+DqBun+8XuN0x2vvpiHsu/naLIzT
fr5sG8NfzWC5lxr/Kcqv5VWTM6+cUprX0VkEoo3n2rklOehDgPn2dCFVpdo+p3Y/
TB1qhNIMbju+FY9s2nyIpbu3PlKoaiaiuYFmlg+mavjMAcBn0k4vZo44tycrCPHI
Vfe70EFcwwh9sNXOFqwLoABpaEcF1ieg+2VrGvRcWMw9YCpk0eo1WM9VjRwFNuBf
lz9PqdlUDb392OcT8a9+nCqtsp1KqqC7+X+nuZFEsKpwX6RZ6GcM+ZeyAfSijkSO
liZrMIP3BuSi9p+oF7BVEaLN7j2ZVIZ4J6CtUXwfyNUFIFqS5hH+ip2SPSUWjqVY
5RKq/4zAI8J0Zj36XLjDIdRPXVl+izFC6+FcUj0AQA7hbfpvpqKQhZl1poa7OnAs
XtJoI7cgDDg4g8eSqJgi/2ppNBVrKWerW5JII/o8VTSYPa/SGNgC+46wYfy9K0zi
1tKZVGHce+demimSBd7yx2hn54Ale20u5KrekVaoDavB9JFbfhtbmhOtvRkigM6e
JFhRH39WhqbY+n6FETQLtyXXZaAWnow1Kizj5JU8ohuqtOUHOErSteC5hbibhmLE
QrivPraHaw0bvdjJnpo7VSFkbYDOpWDb2oCbGBnVBel1YGxX1V8Smhj1P5t/altE
8EebuxWAe9/fVSbX9s4E4cbQQo+hGOEmpzGQd4vd7HQ9feazCjFT6jDtMU+pWmrK
cMDcwBqCABA8ULd8rzN+1wlNnpQg8YzB1qfj9ClmzSkjRqRd/kg9uZ+qiuCz62KG
VS9wqKsvkVLzRdF1JQ69TtyWl1sqqWzx1lVW4X2fZJZgV/4g7Ppj5Rm4khFnnbrw
iGEAudqdv14kh/IWT31jviPY4aOeSdD+GGWEin4xDWbXQkFbxY9H0r4AZOaU3CUT
TsLYOr5oC9qd4wWABcgdeP2lY4mIykR3zYkqMa1FU+4ff/XUL+aC0ET++/edxvJ0
ecAz7RnoD3AVCeev4z7Apv3Bl+6xWKMmNWQIW3yvDTWzc0tXNdDEUsJo+TlOJUvs
reLQCEYQ1AzVm7v6ihfr2bMU08XwmNtplxFqBC3AESYtfk6oEmXzdkeget2ryccl
PBO+VRUDivwpUhWRDWgkwpROSVBKqj/vIy10jo+tT0QnEghaG9+VFK7epW9xuPk/
hvaUlfAjTQJVKJ7sXI5xB7tPhoHIuM8S7X4UeP1tJijw3cJIkV8rn+s4r1LhC8gT
AZBUp1iP097ya09q4kLTBlGMpw1D3hONu/jAuzo4M0PtWC3uFVFVyroLBegNWJn6
1LSFPa5CdyYgHwIqnFbxKupF0EzBWaInZ1jJa+UYxW2xw+maICoSGN5gNxgcJvDj
4ZMkXJw5EkQ0XWbpb1F2Cq/cGoZ2VlUD6P3FsGAJ5IXYG7X18duG7aAPGREKupQQ
btFVQJ5VDdhwheIAuZX23dUfVWocjuWrx+tklkJwxWkmwgr2E5FIe1oFiRT+HRrT
eX8P4C6LCDmUfGjxYja/iF5mYtOeTLCLSomTioth3vWVBSr0FMEyeKS1zG4utMvr
C/CAB89CNEUdbb16wmTsRMWmWGNlsegve2glbpaZeFDnJRDLWkX8adM6x/xKNmkS
mSF5snYwDvC7o+YpmbmT29k0UbwuF92r4UsGEnPBuNnXggg7Ky48VVhWBMJJPWoK
LB4CQ++zX+5P7BDN167KX2h6DtoWf+2sFTSNX6lZuwDV0J+K7XNMWQzPcp62WIZB
xb1yWjN1Or3tdvTu45bpSxy8+W/WNEi+l1dhiR+Lq/JDLUhx03+z+hRoKJB92aDv
Rk/zDGWL+15hgeFlSD73Xahs/XpkuoY5b+joLDAGX4av4yZ5jJlbzgR/QdaBtMlu
QfXi8t56icvuuxgLMrr8TbjTO+6MkR13qtJCnicq3RmMsZJ3J3JnEJRJI9rlEh7e
Xa51oV0q4fXYEuLixkMnnPOkYhJfM4n3al4GwoHY62R2S9hHkXFJrYL0nm1lufpz
jUI9EOnRYSzQOP71eJYcK2ad35h+L6m4oYfwDQmIWoD6dYVomguWtPe3b+2AH88f
K/P1YCKCtUGE2odUCuivE1wApQDm/TUazRFl9tuvNuAQN5CAblJ0llAPrNl/xiXR
r0w3jbspXJizXIq1yBshX4SLXH6SsbHkUwuxsvW71TNWv7x8x7Fl34kBXX77taAh
vaIHoKFfjq6QzlgMjbJCjnz7hDxTiuZeIsXAALR6rt0JRuZ6PeP2by+AG7XTeMGm
au87eq/Ldbi/p/efr7ryIUY/y7ObhbKqZL1zXiJGjn6Ro5l/h2rp3q/74U/prXCO
4A3VI4DfWr5F1fStXnpDVsehiNGFN2A6f32+Id3xRle2oJzjM1xRCdsDkozKQlTJ
UXd0yG16CI+Ky6OcDxugd15fIoP7akw9HwcNueLJAxxqiCdqlBB9ngZzJL+w/49s
l6jPwyl79S9n0D3RU2WWiia7HLamKJSKTLqik5ysVOCLtR7h6NVOQW8u2DhM9uet
AiWyny9RAH75AjRHCC0ELYLixnr2fV1uEtGirwND96SFqry0nZyApcb6sZCupdYK
moJ6dfPum5IWilXRjDfDrUAZlK7dGqA52QbB7Ifd9SX4lstdGIglAUIe+Xts6Dak
uxu4kU1NxiTEDr2ljTkOcpVCeTaq73ahm/nOOlLmhkgv8p+FUsAksUojmqdA/oq6
wgaoIi6TJNaIBKhIk2RjoLA+5cKl7CjLsY/uv/UyU3aDlXOsPEzSxsWR2Rsx5Kdg
OL4Q4MDHP3yJa2IF+6kKIdpa4zNdkwmGKk3l4XSF8JDdBMVtIW5lu4mL4exsCqut
7hROJKSqODhrvOEfa7Sjv9uIvOOVs5UdQCOw4/1rH0ka4Y2VUjJuLWTw/BKDxy2r
ZA6TJNvfw5Y5PKOquh88LoWe9F/wZYmyxDN3E5h9S0jeImN/A3pqHolBMAsPzuN2
gB8FXMl19ApHjFYAUdJ5MtUX3gxdAaZy1Vy5xTQ/SLBv/DHTvng5I0k18Wi7b7mQ
G7aqZpOBlw8w/l9/+k04NnRYnNgS/yjeIGefwpCnYE3t8gocwaq7c/7BW2F18mQT
Fgf8wQqgzj2SF92GIUw0xFFvdM1B0SQnGJJMdnhlVfBDafnRkiHp6D302dpD1Kvu
l2HaZOlgHpBcpDQZl+RECYLbpnf8llAJrFdRljZq8XZIasACqprbLdl7X40wfD/m
PQo4uCQHzSOHB1GNIUcyJk+MLxBgCnqZ2agZGTduWQHENQRnSbVF5lz8ojEdrz1P
1TqHrcN1KUgmlNEXnCek8yeukw1zXzVgOoAHUOheRghfl+E4iBnX50UOAwU8w6Kq
jeDWfwVHY4joHH1DN8h9TWAbr73WWJruytJy8uGBJw+GEKHkL/kkA17dWH4SVOZz
eB9EmXwF1pKai5H1PlcpcGXPf8TTwJI5fNV7EZzwbsh3nKgFjirXOIBl9tiTuKQt
JOlAOaRqVHbOjtlH3R2zCZAV+yjJ5ziVeiqAS/Ji91J1cxoMlae7rv6ojXYg2d2l
ddJpVVVf6vHoGyTBqba3908FEpZlO74t02QzKbpttwG689SPnnidWRba0TW3kyPL
BnCeoRvFIdpxsN/a3CrfCgq/A+2vM8EILlaInSGs1s89xwlkllH3E7AvH9cT2qyk
UCMmFMcEkuwtdAXhPCAWFXe8i8GIvOcupShLwpT5D7E7Dkszx+fyAbNmbgOYacYl
yYovmsTyhTvMbA5mfThVg6Agz8mLctMCcvyPZJgIQHK4vPJCXvN7Lc1NE6iy78gn
+MI+ZET6YRKmi2WyAGeuxn+Fi9qcuZcZumkiFr1joIBu+8F9Gs91Jild7CmBwE4d
/u8rqgdSaoqhGs8HicdzZaQe+mmBoLdiGdkazxDYx6Cu3VqetXDd1H5SmjqcJXhf
l2VuZHo1/aG639gU9JeSvbQVJwSeOGT08W4ujkf3X9UUHxFQc8dHIVkZKgceCNCj
wqfPqAlBZ4lXDZL02WL4C25oQsxpsXLBj8vidxKeEbZWA2pQWSyFWWdVNDWN1YIQ
J25//JbU04fOIKPdGsZXrU3SuJvHdfjJ0higZpxCsJblY3S0xbXOfaImkBTYylRi
ZTcwN3gwq07uz7Ycu0ISAaADUMISg5HFZ7zoTgkz192tpd/6tEZ6Rwu3o0qUaY/w
udNlJGAHsXkbgM9tmQaU9Ex4kIWjjNTC/Vi5oCSgLNA/8Wtp3Zx0L3FKNwq1OsKY
/l8ZfhOuJ7OMvFP5q+VFvKmuIMLiLVR0KjqLTmbIjT5WYqZ3T4jah+3Cz091vkg6
zF78A5p0fgtbVjFPHQj7Ot6VOePEkciJhqxmjXzm8t0qu+bcI+jxEm7E0J8m7meP
7wIYw1qCcokv7fEjppj1jZC2liz/OjPeRHwzUAIIxh/6oBXySStrLEK4OsvCG6Vw
6KpkG8uCupDnrEEFZoxVBs5ZDk7jMyfftKkVWGB131KxMXQSS0Dg0o26+kpuywmy
ITL3DkCJkUI3IeROJWYr3lKgWlE2eJFRRzAcmp7CRuIQRCETI6PnbMA/emHjDZAr
EUhfJBmD0CCdGKj0GIYBQSlHLHfMUe7+JGFwgkMbdQtWU18zy26xpAIEW9llyRch
N+JHpZtLHrFgDuELUdn0dh9Q2gjt6CK+Zcmm9IpLNJ4dszzw/qOzk29WI+wTyAAm
x36vz26WmZqcf+j6VlyTXhN+PjOBopWCK4cr70HwwM0IuLPq0+iYDM/X0bdAN1Iy
cVVASVpULhXfYk59gWamQfkzbxAiNlcYohzTrLNquDdycU71qjdgZWwsNwxCkIEB
8QZUExOpcW1HYMHr40GUOsyJBW60lGl7UBRlkJx4J8QzaYoWPh5neBqgU19+bWjO
tdWJ547/gDl8TKgHWx40O2q2rfplT9Ts6v539pxP8KHaKlDJLhaXkZmY9umULQ6H
y+3JcdDhISscUchmsZZwod5vZnnEL7RzVc+uVrNXAw7Zd0im32Gb2dNGgGE4efcA
Uq/ODX8iL6TEX3/G8ktvOiNIX0kWwzcSTWPBqrRTwyTbSWGEL1nHNbEyjIH5xigH
sXI5hxpoXvdZymEL6Dp38iiqkiTzzNuCmXWG+DmG8VLOUrc3Z/rdc41pTKJ0US2z
MS0rfSv8iJQp02IlGHZwU5HtTjoy36Pk6g1iE02nvQsVYHaUMCxO4ePIc0zNUVT2
ENf4aOH2OVJ3i/AHW5depsRXM8Mlij3CbZMOTyb9WJsB3XVVDCMI7Cq8Z9hKz5eZ
Lbu1kI3qybK7nYxlJqejLQZBb0UFrzFkmmEvDWgefHE5+vf7L0Og2opg0X9opkGA
Ddnd5eUfVLmxg1pRvCmeSKO2Mz2lpZlcNl42oucIjMxNjaq+AH1Wdg2ILNxDa2M4
38F9ILdq0HwaM+bJwXRQvjdRuAYYX1hyE0nHXk0WJN2JvWNLvvJwQ7AMuHYNBdOT
VP43tkuiJJ2ivnBXfJMF2+wCEfBkEZ5fIoFXQr2CC0mIJ1YrbyfejvBJc3At81f1
9yOkdB9nLLVodPvycNwFgxr4fmx69L27B0hqx1QvZnI5jdR/vorLDYABf8+pukCg
3bfQG5Q6n7tS5bwmMAkPP8ODnkjFamaMgB17CFAiOSIFgTiJ22gTApxjefN17qcy
eKARwlewUf4cNbSJmjk0V7I/NAJxiq1EE5jsQcI4+z8O38fgUd/wJuhRKZQa8vSz
N1sPLrhgJaWyyNU9aBI/ma/l7uZj/qFoZ/A9srbAW7lFNKzFqB4nHBkDOxkGn3/k
kakl9aI6AHr1h5SUqqrrfY8DklAKqolGd3PS32kG+U9OLS5YRY/1ZgCohbWdIu+0
IgZov/tpjC84Jt6q2mGQ9NJ1TpiDa3flUVa5jCfIBxa04FY0aD+Toi04BWZoU2dO
tw1udaYHKSMdWGnmHcqNVbnzqbiDHZMt9U9CJGFdANlgV++JhNFe1qJ0gOWJ2XDD
aBJqD+5aquD613yujAsCThbnvr9sq8RHtoTE5t+OG2IYWbSLqFFv4mwa/865rQ3h
HkBj8/6l7Ci1Fv3ulE6K178MF2JrIGy7U9Ce1lfDaXtTSKHK5QlMItILuSnhdJ4b
VmQSR7re2I7KinJHgS83UGG83oaIKUgkOlV4tVUe1BWNAhZ2nmGNjXORDe3TzXRI
RILbgV4mmKFWoMKK83JSdrwn/ifsGNuWPpIV4Q/PdGadS+UtjrnGzSnelQVhesIA
Z06f6rjJx24yNmERBbgq8WAX9VUlQoPz2y9fcqy/62bEx+Grge21TJXXapqzXCCW
K06xmBDg4AjVrDIuB6g9fqb9gX4KAzVKErBC9rD+jikqqMB4SXYpRXRr2tgjqF60
jpN3Llmejbdgwbw3gzP/l7aeZdhXvUIWHyr+vP6LwtIM4njWfHDnb97pHTdS3Cww
gytztKULDGUPkXdid/CF3DVKOhGoLOjIb3kqXbezNd53dMvShZcfZWg5cMs5QYfq
hHxEcm9G3vg/J1TQxu4ZE+134/aer5x1/SvOSzQDRmqEnSL7lXPFNMh880c0WT2/
Dv+06JIsTLfC4iHefOVuWqT7kw2ke5gvCFjjXVlljAPrOoIqjgHBamLhzaZ3KutL
dJACrHpq4DrjS+8cazp9a18frwMwPXiN5UDofDJRv0qpJrtaimOvNYhdOY73G/eV
5ZkqKv5LAYauExWqDfTkiYxCCfxfgkHkSi3VqGCjOMm7USE+WFOHumLLTzlEoGXi
PsJ1toHlVS5e5fNBf8h6FlHyv5BIwdCAxCNlSmZ5t99KXP2Z9vuha60JIs3tLMDi
d15oMkUxVgTR2dXQCu0Ua69LAFnJUZsHbrceg8rA3/wMwFCwlX17le6VVnbZYjR6
p5GvFdRrtBe7BprtlJwXNokY4PDo1l2uKDWmw3TcsVyaMk+4Egl5xTqI6e3+A/k/
Yu/zwZHlsNnLK6LqlGSu6+A/pPHMlDxsq5GXdnfO+lgrFhvjHpCsArlv6yi7E4cp
lXT5w42UH4scIwOnvYrQoTqnVf404WYLn3aMKc36ErKKdIZnjZpNU76gnMHizsxa
aMSfFaahGNgP9WiDQr0KGrjh6ISXe3JSB/Y225Dteb3lGBPwdHwhsbS5+55z+iYX
OBApMZsU8sZyMNP+53bPJltCZMRR3hJmuEtYE/HiJXg3heC80jW/CzHSIDNZNcry
kxqp76R2Pv48DO6j/ljZIjFnjXeNgzcsLF+qkHigKq9Jdt4OvT4cIBbacweLqVm2
m1A69qYcUVGFuxyFNmzHzlg7k73WzADuUycq/pNYW2MIZBKabv2+Q0Ey8Wiq5Cmj
41yZLu2aaVV2T2ZJMxbLFiiXKBdKKENR1g1KS31sKebIhoxV1Fn77dZRrHfzFsFo
H7JjLaY/Lu9/hIprzpuY6TDbkMmnFkyG9FJ68HURNrXVFgP2gvNpEiq+3T08TDXS
Ro4Tu8q/em3MeuW1cR6H0twIxYVmFm7T+lTEvwUvlX7Mp5nTxRUnS9x7IM7pUmqS
8C55Xc05xKj73tG9DOMmw/mdqVYvjZZH/hWhUpAtcSIluV5EFWEyB26MIEDPNqaL
74H1arg8b6lpJ5p4a0G8vNs5T4e35Db2iJackovgWXmjbHh1KKddfQejMQKItvJV
nn/gboTF8NU0wGo+LE4RQTMAscMkMMNiu6MzdLq+NkBMHyuDEWNQ23BTaNJoB/Nz
Q/AVhW5sFm0ZjZwuLtbGISnCqyIwqjseqJPcKSNlRrJ/li2KEawgPgXBAKRlitYn
k2Qf8dzKXKyzlsdSRTIM+6aNgsuJAQOlV1B7HQl/IKtDk6xQMNLXFN3UxTsEmENK
kU3w3v723YphDtyku7NmPKE8rD0uERvUGT8eWhYMJ0fCZzoFbG4DAHjOH2uZOLHs
+jniZ224reKeLUPRSs2tMLgi86Naqife9F+CiYw+9fHlg8ftuodpHfOVyZxaeIHi
Gmv8ia4VrXZlt3IfuZuqa8BOUkmVJRfsD4xSSCWCExvvzyDctSsvtBHKRPUTngeP
v37y8q1SWjelbnVVhV0A7Wmq2VBEdRxW+ITps8E9GzeXfxdiXOZCUldjJfcbp4NO
cU3Rbrsvj/XXqnnzciP63oRN/l37wbXiLnmIit8dF4ppP9PISleiZifac9UK5Y6l
Ij4YT8/X6XjSeLNt7sqAPcicfZTFRboyyg3bI3cRso/1xskz/DrN8EhO7D0AQ2fH
W2JsJV8C2QCvQNIZT3qgjodYxycGuR+JbUt0mYqV8dXeE8v2qj8WmH4IujZKwRKH
TZ8vfbBxeAL2HACF2tcJLrDIkR6RMnY8d79ovTbdF4SF9mrxD/880I/1Scdx6lJO
DKQLbD/eIUOJT05K2TBiYexC2X9yYHBwkIDJA+ru4Zj+pXaLaVNE0i0IFSwufdxk
XG0JdHzcFCadtyR9zmihiqTOKQ2Z+2rFghbnu4DIZqg8feHRe54KrSTTahKCViz0
edis7dKYU3JlXILTuA69rXHxkR204atgVOyds/htCXZ/QckW54Q7BjmzC86v8sii
kl+js9p9+onQJxpHUKX9CO4R87EKFt8boTmgT7TqIAGAK73R5/EnmiBxCc6d7KIU
9l4SDQuVogNfnJDa9kStwb7Fn1xNAnfldeXpWkoJGJyOsM0nOQEI2bCumaO450Gd
MXqfeTwqKApGbIFDq0wBuUvODHjyjK/ovgYVjeOaiyrLwtGcVjzRuG94e9YbYCP2
SBKkWCDVAudgtgUJjaMLnCR+4oRsq7ibOXfnw/DVWrv402jgcGpD9ImB+l6Ro+x8
17VgevmJBdKOAaB4gl+XZVp+/x/nmLvA/g50Ju8/LRutVfDqwkmOxXJjSr9ZzMVY
aL0/mVophqQxfF4i9gNAY/NuzRZNUCqr2DTX6X83OxBnHCXJGYthE4pD5JeaWjUM
ahn2tiuIG26CCBL/LHgJXwRS64TQSzJlqKPB7ke8gXizxYKg7Ix7XmSoiyC1illx
dyGAL6Nynm324ayAp3tyrmGIV389oGcuZ0IRHxGwR2LgaRsVSUWJHLGQp7q8yrXa
0TPMVKdaazgIXayfwgO/kswGVfTqdLC/zcR5blnphFzZcB7ZCx2ZePi/7uSiNw26
fzW2UDzbNrwHGoLT2eb4ptX5tZSDi255SnA4nuIQt1bvMSx1SsDesf9iJ7EMnYmQ
ZpN5ZyWMQL3ueFnDblRXfnlLAihicVj6FSxeEUMeBjy618dM1tlWJbKLxsyY8pgc
dDxPcOuPmxHWHw5bSj35JFlmknk6DCCpncy4f5Q0jHXMDmOnmO2ROtrQB1NW3Evv
vn2Ykgg7HWhXBTGHGg/xaHnYz6Dzr2bDddl1gAf75XJQxR/V/cqMfC08uhIE1ncj
ZUwI3+PWCYgAsB3jHX+9TBTSkgL6AT1vtvSJkwoBOGYHR9vXBVrO2gXhLW6L4k6e
Y4h991Es9BWFOP7j2CIUOjip33zVHpJG1vnf+SMYQikCW4Ga2BvXF2L/JNXuJCqF
tePJCjnBaRJy+vYLfgX4yLvHgcr29wBknYmIpM/SfTFk1Nh/mchsrUqE0R8IY4k7
fprFplf6Tp8AY6BSPACU3CK6SXXsCpGwO42G10WAOcx6Jqv1KhHB1L49ly9IXUzg
ALQ9qM4DsDfNCT97ADSRXVZDRemmCmy8Wr2HU2dHQFixWnFIz2RSnEQhBmCLT3Hr
xLWs24Sz1aukVL3qejKYCFTXM8dGP6VZCypG8aXH6616N74bmMAktyW58lQeDP34
XPXrFI+HSP8JNzhS0fkFzGX6gePsvvsqyHg/g1TZPJTt5S3Jo/sYmiv7vTWQqdnZ
AbL9E5bByLzsbecuuuMntg==

`pragma protect end_protected
