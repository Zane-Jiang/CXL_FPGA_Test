// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
VqvCCXsXn0AdINsme96AdWzwHlCtEp6m8GZIRodWxPPkBo3MwsndtFaRvTPac/Bn
ausgbADiJneNZSll9CUU8UQIxbVaLwiyUsJkNTNdlUQKeDytmAe6jkapD+orCM3k
o0ta7amzZde0zHiR4parqNXBHy/JNzJBBHuxO6x4J+M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 120464 )
`pragma protect data_block
7DA5caSo57sPt4S7eI7LF30rwHIGYXUvYpzsVCfAuC7Mc2+S/1YT/4BsrcOsYhq3
+9/09pzfwOqvOSEfWbt96eF9MjGkfXEmO/cUahjb5yYXxrJp8GbWZtL/XwTyHl8G
vHO8tfIj07iGipSMQ0ypJYmXnMR3QUR0Msvm1EE0SS4sLeu/nubJLpUxujRoo/8D
AryOmV1T1GJVk9VIXLwM1qqlJZvsyuYg0qBvbErVhH8cMcum8cSCORfJ3sWKVI4K
u6SkYtd691wXIwagpwqKm7HgbgHmcMiIkqd49JMWQkeUVxOBDOuGlWSJpdzild9i
Qkp9aZHt/E+vw2XAsiO7zpoazKvA9qZxVgNpEoD9R9htafxMvPNuKqmq+43UotOt
TwH7en90PK6uRiSu4UHjGZYJl+I1ZneUC+ICX5wM9cm9Gtx/ffrdnYrqEDxkHoTH
tv49cd+xbHHtftgIAmZsVoYRH3dWRvS6qf5Xlmexb07W9DQGPAQJluE3t3ec3foh
CB30IW8TmDYyf9kReM/NE9O5omh4DqV+YlSDVhfkRLsXYCAB889gWZS6WwJDGYQu
KF0YKlSCiey4qAlRuuKYZONn7PDkK6xnR0kHGp+20TS0X5vmTq6kRpTLtZQ0kzaj
0vFwbsGdYedUVhP9y/lSYOyduj1hFuq4FHwpD+YI0K0wRHI22aV4G5eqRQIy9bKx
hWxMh1edsh2rkvUwjaUiVYzl0ZBlx/UPTAjse9P+E+uVculgmiq8l/sp6JQUYd8n
DpDpUL6eePRnzzF7zOgopi656GsUuqT6+ovEKh7ahSl0G/XV9va5QSQAZ9PSRrJF
vy5TBWMTPqLj5OO3yunZOTJ8Hf6ORcISR6SDDSPcgc/lPvCh0Ep3xVxdCbKMIKpg
eWSia/dluMz/Ck7w4GlkQ9AvSXRPotVFg8jcBBmsSEEFhinP56iGR4NmK7JJHZhG
MLlNjP3/06imm4Hf0blQN+9Kykj0IMw/6hCdjK7sWXUDnLijCzmAjSz3MeeO6apa
pDkGrT6QeOP8PHj4/pcplvnAeQa9y/xp7kmxn73gcaIKVUkizUxEocOISM5sOF/j
asYnLKIDGGw1K35ns8DDjdEgdgZb2wxNhB0HhdldoQCUpUMOAD7HYnQQeXU2lH5R
A4NKyiTJKOWttRvhG4Dm/lqbpZZN8H0uGRAcejXIOS9DEJSmgGC1j3Kl88vb8xyf
0yRa74a4nOgZC/0FuWSrzUPtFh6jPlkd89TFSfZrc4hOWh2F1Ek57H6/LMRDlzCU
+FNNG7/aC/nIaZmx6vtEXK4LoLRW16+n0QcilebOOTbEKJKO3NXbH3KqZE2O6Ozm
UXlIcuJM+KKyDzeNV82Frlzscl+Pi3uFPpEXGZNHdKIxx3tmbi/uSVDQc00+a8Hi
/OCZ7MtZy1Z7HoSbIV2ER8gZ2+GdBxqHUQnoQTzXIFYhtFhS4AzFUnEO2/i2rcgD
JdFfcd7WHeSfKpWxDsRdu1cwClq6ZgKLEo/Vxs49EaGzGYaUrRmvJSOagQkoYm1N
PWcTr/4B3V4h31MO3BdPXTo5th+u+XVchv4GRovh8PJR7UoQmdNnabLNh+L8fvk7
HgO0Y0/KKkgVygn1BTXcOO91YlFbZ/VYd3xrMHiEKuICa7YaIY+EBqIFb1m3WZ3a
vq9ltmVgNnNuh/on3h6lNEr4UWGryuFu2QHZrTrC5nxr69jD9B4/eSv7uNXPF2Eq
+zFOMOqXBbgdC6P5Xs9z1K/1GGQnqnDFJUmXbfhnTCEyTff91mc499k9V8wONvg1
mRetviKqRhCosUdT3CbN/XjRP4l29XTcY8dRueTTfa7cRfTV5ihTeZGzxrwZiANw
UmsikXMBByFkfW1szTWir3YxmWDw9lcugLdUVVQMjhjaHVA4VU0WJSiXpU8bIboz
9az44hbxvnjBovhzZiCmBUVVO/vnZbO4ZRZuXIxfMJRiLeZSt/A0cHEjr1buGQT8
kSU9BnUtSNFvC92+DWcOjw5nqdiuSO3jMT0D5CnUGOipypNjIwRFdjSfbQKRGEOu
yY3lAZLLuYI4BaZiJymoZZUE84ngDe7ZB5G6JKGSyTFNQABrbvovo0oBcNp61Jnw
OW5BxwOm0w2rpWrjzSa/DFbEelap5q44g9yDn/HvNGw/iauFdj2Kg/N6GwsUWadV
1UgPYuT/NdyIHKg5DN2nTSfymSYcEl6KKsCASmf7leyXdjQ0A+NlQPZWKYAabHmd
pL4lB9zYbw2LmF0fqafkedUdLnp4/nSmL8Tk6utLf0ooimXIQgq7Sqs58eBWzMW2
9OPTeGFfxsjN39/f4eN1L4Orko2cSGjLfXn3TPYxRGAHVffU9RdwWpSz9KFzIshT
YOqOAcM/u3trh1f1gwDZGqLiTNOjKaiwASRGUWMhRBHWWFnzKAM4M1mcD60zsRwv
KLTryw5fZKAbx/z2X8F6QjrnTSCEZhHljiofT3uHIWsU2TcLmQYq7LbxnjyAQSxI
hMXxE3bDDOBJ/A9mvZlPX3w6OVyN1S30m4HNqWn/lCdVT1d7iq8zvzVhU9l/PNHW
Io0yyRxdKUAVWXYgh4tHG4AmVH1ZUVFFXJI8VYt/DfIHkXOAUrRAOmgGGCjKVs50
GBP64XVatrBHGGfwpO38JRvGzzHjVsftFcO8UzlRSIP1NQL/IwoJpcYS4FMXUIvl
sszDlBCyCeo1M0qaGfdsbNZGxCiV1QYlU9P6MdnUmcNdMJIm+iGDVOOXqJoFoUJY
NHWkwTrHmfSihkLi+1J9gGBH14rKCME8w8uzT7plEdeOfrEnWQQs0gdSX63V9XN4
ebM/Fz81kv2ANaIn0CkmjJ5yqzYt+CkIn28rHqviobcT/st/pMHQA+cwXbLCMk0v
ddZNqg9QPS9HnVOIWBDwU1aXb6LeNNB9rDmt4BQ5v2iXMdytYvcrv2XLxysS4My/
Yx1MuD/WUAH+jtVOkepo1MMaZdfBcB/IsGsjDywIPVovonrtl/Bu07tocVzxRu+e
FqSlMJlUnZmmodEJy9eIqVu30ZRq8e7lhadA0yyLoBkhzV9xOoHy4Q8wFbiSBwMG
E9kgfgi4YsyWMjzbp7Jq3dd2J1iKwH7X5vzY2lceE4Ui2fEtXC1Rjx/yYHtgkUrl
8ejaznwSETqFah21oFvdOMhjRT5YChYY7hZ/CezVp/X4J4Jr/xDGWI8CjZgqU7sN
jHlo8UdOy1d/7lh6461TAf8vzSBNumW2gOYGM2buAR0HX0r3fEHggPZ+ht3BRr2O
O71FCmFCe4UIGbeIIhKSiP9Q91LWiFMjG2ziyJWHA25GiSdlgSGBkE2Draj9w54D
WP5gEsE07ALz45UfsoL0wcvcfrOu2OjSVjLs0QK3rJ4n5fl1XGrvBnuBgFn8hf+Z
VfkdcT9sfBHmWyQ+bwZr2FVme2U64Rur68WM8vHL9BsCD9I/TebuUXcPdL5VPcOi
koo8+LmViWy5hUanYj81tOSrmnZcKgECQW3t1QyTWPhpxyZABceinczErCRk5czX
5YZyO+wbA8/FgofPIcJQ1jCppXhBiZQuhFpKQnp8DwxuEUsXi+GA68r9X75N+eYX
4Uu/dTAZYrjhp5SF1uNhdf6sseh22+SySMj3SAS4sAG7zYe4iIHvvAgafhJ1GuTQ
7C9dGIh6T9Ko3WnRUjjFRKp7t6k2s6ct+jsKzui/GtOaP/ocDbOCfCaIf29HyLit
ZuJKFw+/K/QRygj++ULm6jYVA61mmsX7ek0Pgli6PzZpp40nOCT8DnhW/H8Tycoa
tjXWsP2a+VciKCrrLFyDmZl9XX6VZFwPU/00C5+BnphnNljcgpEE1w/Y+pfAUrLA
s3ShGSV2+YYDNUNPPo/zkAv9y2lW2nedDfGUUgnB+76ZRKDy2Q7psNtY5vQRm7p6
E7vocIsgaIJkbk+OvQHBrUP2uvma5GfdRd3fG3vgnRGOIWcZqbCgJTQYH16kkfw+
ejWz30qjHphWiILqCl6v7y8mEHfWQWLPaPCeQ68en5UZRuc9jByz2zFSnKmiQEuA
OVyxo81yw6ymcQ1HqsjpXhpg/dZ/od1bsGOJsSdBRE+nFAWKOgSmNl50hGZ1QSPs
mlnVu+vGVdLSFehi318rlOGKg23uQDwXe48CebDwIDh13h6Ip/c57rgpeYTfNiGI
I3pb1g4fC5Y6BC/n0WMoOoSY27GALYLyj+4aWiwP7snKbpPxv+brCjZzNETphFXM
GlUjPRYlcv4jj3S9eX2azzzEZyJ87TRWpfIDySIQlQnQBbcQ8T96cz9Gr7Av/ZSv
dfvz0U5WqyF8fjcr7tOj0IbEiisPM4LgTNaBpecQUoiDF7shj/HcePKPovPkex3K
9UJS/DMi3wipitlIeednxmr/5m6lr6QIKSZ61toO2J4czoNxZV9jhkK4ecXDakmJ
Bf7FmZjiXvfddK7xY0yEAOSEE9YyUBKiKs8d0f+fWlEXSXowHgYHkyFyMmFIsUQ3
2UEUQidhw3N9vGykiV8GH8orVf4FJWvspj64f1JjG1nGgk/RC1sGKfvKdokOB4aZ
6pIoe5kI2W7/UNlGVvu1VUkvJ/WBY+9rQbPU4YRKBF+otfF0x6jVfYghIUDx2Ref
KD7Mp6Cq7W5OyzTwxbgxK+XCbuf78+1IzF6p9joDWMYSjY+cjU4162VpDWfHMNsF
osU4gNgJdF+5W9UBYzFK2TfLJQWXv/wXq/qZogwmiTWgQ9C+Y8YbuRqUfNO9qukG
xjowdfQqEtp4Lrxt9KErlSvtQki/rf16EszgJp7AC/gO5qRZJm10iyg2sLoonm3T
6qbZPw2IGNynNcy3udD+nXqYxToTJdzD+DrfxzOU3FYz/FDTzy9nHDX8YmR2xNWc
9Gi5aGbF446CNXdawdrO5wt6cYx6+FtriT4WoNcC4DVyM09WLodmPQAsg6aBNSbF
UId5soA28ceVVUsYd6sveQ6R7/eZytIwmMoJhx9TqXzKE72+VPzeYmJu2tWAF23P
9lpFJKjEjriq8/mSxcHkdpqIBy7GegUG9qk5bIRV9zmxraLuRZgoosF2XHRsV0YM
cCpB6t+Nths4Ee72jwqnWsVgO9V3tmlnss1Osfb5hEKLU5M2uclHyiE2ExOR7K0w
l5OtCQUAyDSc9aWz6td84OMdaI+x907GklR+JWohaBfT3qS+JL844ic2+FAdrPVo
W/2NucZ74x5mIpWUzXBhncTlRcZgPrR6W6kZRUat+NcwMIKXLy8in/w38vzFWs3P
A05sY7XQn41lXnM9P/nkFVyD/b8OrUmVj6i0BU13N4f59lZM4LdpN0uxCcOqrRHq
gfmEpMtsgDucrK/VFhPTNSOwI40i+Naf1lLp9Vjo7ZeCKxo7r0gseTWheVImjaw4
2xHirQKzJIvHPapcEaUPCLNIdIlMJ9kNWEwqKE5KY17pv+C71C6k5vM785/0Yzsn
pbkjhfNkvDM64qVUBm0A43YdL0dIpiGJPTpm5wuomrJlXF1EJyJAIlg57qSC7WMV
KqxJAfAKwURDTx7jdyfmn62qewY2hm74OnI37oKsEYK5GxJTttHSCMKATSB/JxV9
AnmRJFrCfb0v/RRrMns61LmOkPNwC6nTvfj/C8mSIsISfZHocml5TCiARrD+nneR
BxvKGTRIYTknopugikFaZsgsD/UdAoFUHJVriNtDsMiyvfm4tk3rWXN458rqlm4z
qHmhjx+mLLsyUOEzz6dzFlEz4+f3eZ8wbsLUTEHLgGbphliehj6+KaD4ovAnMMAr
A8HP28uoHkL4dYoIGv4EwUa37P15DW759woHdQUOKk6T70fxLBlqVoQ7rCJ/R8V8
QG2K09lyBenWRGXfZQQIlN277cjP+M+b2nMTyrMgon1ntlM4+wZfk+f9lvq8Fh/y
rJPeEmZSLYyzHi+eWy8WqRjW3Dnp0x78kZE4JPpcWS1+0qv8JnuDi7gXjBasSjku
mp6QqNcJMuUaUapv/nLgZWZkKNz1Ze/Ma4+XvVOs1rqBHisLlyHLS31KYBSvOeqk
BnKE4KhYo0PFOGu5IExfl+668kTzbElW0WEbfAROv5Us6t04/zjm1dCCUJw+UlPQ
I7i9sDNAijZl+RJAacZoxKQqZ50LWdq9Cw1gzkBvEqIvFPrlUmK0KIVikMdfITLR
1Z6wYQNMtpReVraMxs2XxyH0rsCUkChkimfvH8mLnEyvzu8sWzRa2Z7aKo4VUMOn
HH8exVst+JUFFB6JOYcsY0L6VFM+5Ua/PqM1+BlE6U1j6mvEqfEuFVvNVoNkuH7c
f+3UyBE+0WdfL7C/Xxdku9H2LVfGxoSaB3Uhj02UqFJsOc9IJNcG9hzL14bBUYX7
v05RRkHS42jp6EuIpvVeDr/Y5XUBqDlBxqutl1hENQZUvALjMKWZ76bTL5nIXQ1G
W3N987XdfZ/qKCI3I5IuR6rWMFTZXRGhG/RjRi9kFkg78fWzk5wAMpInkYdbRfaO
n2qxldaELVfFWLLjcDykA+YoH44F4kRAs9V2YUy9+OXVn+6atS1Em+7G2GF5a4er
RqaKtcDd/7pE36XKY0b1XZ9KgQzignlzaxS+gR4i/5gThX2dyrppa2MDzx9maval
jxJSubjRCG/6Bcccs8u0nyWH+PkeKJz6u8s7psaoSVaGFfZmF+3adHrzK3TfOa2Q
TeIqx4speOAIFv1v93NJrVZjWd8bSwMbc9yH+y0Wrg9yfSBHcfzeo6enMOPMuZQh
zM6qfOV+ROkmx/9FXanci38eu8mECzpLjlOnCqqLK5dbm2HFuZYjmQ9Z5kJD9StU
xI3+ZBQvse7Pb5yvwyMLkX6Ay7e5AYr1hxZ1HtXtzuXxlJOG/lv9AhA0Ppz+LlfD
spZxJrgL0mkML/LDsrcG6GIV+Y7zBhUeNEKXwH6AbgoGmqigks5hKbJWNAwXnWMu
BIidNysN5HvuzRiBTwUnqBfX4EW6vi8FEtYN7wAfNLNvg7oIeOOHdIUYpVcPCH8j
nVSDkzOINyCHj+Vxa0FKsvy8tJWHAn+/v2bVXIj1FN5kQaTesd3EtLGK+Ct5WUCB
mkh9Xw4ViVcyWGUs725M0PyJPbDZntgXTgzMZwYVOVDbNsgzvMKSjtDUowCDC99P
vd8zaiAReuOg4GGc8ifj9/Hjq5pfdbx7ArWAZ09KJcvMi80MvQvq9//VIRrXpno7
oxgOPSEmtimmgCDbSVTa3oKoEewxhV0eFGtdOMPVpQDg8baje//W75eRrcaSvOhC
+k3bg09q1dyEfUZ6B/3ARqs4r+U/jXGoFxdFfcC2d6F6h/DVVGXFDdbF1u8vhCPb
qj7FqWzJsNxq7QGRrxc405Ot7XuBEuvR1F4ItSVTjACrgFwN+eOHcUxKxvRZc6VT
7hHTw+7jB/giviLtTZVYdit9lmO5zge3G1yeN/7NrnEA9n2qPjQtK5XKh9tavWbL
awITsjuegrAg7dT2IzK8qvr2e/MGUwVqXELI0X0V6RS47W2LoNw8vznEPlMHgu15
SnONyvVqjuJ+rrSOC9TggL7jycXrtC+iDh1jtdgNkgd+n4joqLi7QYPmYLfJyuPT
vU1vXb+UgMdOVeTqu3XQlIfolN3jAVWwf41YsNRQqdScJ+vJaBqeicXNuyXGiZgc
/KDj51BKSzwhfvFtPrkazsM+Idzq3dtZCeAcv268A1AO6m4cD4pKlc7VfaqgBAZ7
U5oldOz8z5fYOzn0rn6LQEMp87A6HH0ggabEZCTZ2hDtOZWMgYT8rSRLGPWg4Ry+
tqyU8VlfALOr1bJjzk0zuaWtdI7vC0UnDvK/s5WdXI9j9U4lFxRrzktSmz/K/ryk
hnNKNsGiwway2KZ/DQNoc9u/OliZnUyzoLrH0/RsEbL4KCplhGS5jQOwpFsmdagM
yHdGsLEhAp2mlDwRY42553mTo1OhClDfz8yDc1B/khTS9wY8DunbZpzghlBuflk8
F7rmCa5hE3e9CLVkDH6tgerMPEP9jVut6bvqP8URhhxN1j3uTbQoUO7tcz7hO3a8
l2k3p+9p7NhcppQreGY7kRrb0/agUhob+OhD1kW9KPvHLXlW+FFaKiCkLIjA3Eyb
HgWbBBMDhTzNewArY8QXrWtnlXAdJz8wSrzZ6gZgJCWB2mmDq+MpbaPLL7P+IARy
uNYbelPqnRyllvABx29fyJaRHu+oWro6t+4Akk77lrjzzkYG4/B+IXYOusEoWmiq
q2o0cMXF1YC3aSZZJyQ2oflgdTJwYm1TyxEX9btz9Il7WHLgqdSNIwe55Z2O5vi8
hjg52gvBdJXJVkQcYlaabaFgN4ZyblOUNl1XQ4zu/rWDdVz2YtrXIExFseFNKCHw
MTwrBji4b7gu3cCGVr9N/BG0/z9FF2Kn4Y47TGZDvgtcSTwMTiYkEFISODuA2MhU
OCxicHSKFyOL4w3v9Cj4vnh2R+nx8Mw3GDfAMeT7ORfSe+Y2QfS+3FlYS3/rHrg9
DvoFfW8pIGDqYZN0VD4dL2e1sMvzQg8YEKvIGC/dwI2jKIgPX2K9tkm3v5PJGJxy
iCzQwsG6gvPZUsMCYs48DyqiJQDyNOmU+Dfohj4xcs1qqEhZOClAbirpL9lKIaSn
1EVkBIxdXWTcf1LpeluDTpkLJgxT7uWKwMhYyXkZ/3ypxkCZJLkmbUsSIwR3+pD6
Q1GeFgiH2NwLO7Tn2TdiP+jrXuRUR0jgxctyhmTvO/eq9CsWGzoTaYB7bkvAQKNi
8X1Fzn8W3Rvg1Vnu0hS3yueepOqczy4MT+9erdVghtwW3uG1nph0rU/5b+4dn88M
PFrygAWeZhIKxm7rY4WiscGdNEZUSqaVWT7QPwOnUFz4juzynoUDXk8KNiHlLKbE
wtpTPqa75YxVI7ZsiAoc6RGGmmeDBhLOGhZ0dHY7iBqAV4N86e4gMOWGAFhOLjFp
gZcAIua8sSlJeKQgxcPSaWPFiRKeWX1W3SXTMKxvmZ5AQoIU0xpseFH9sRNzWFMN
wpGy2QdOXKBT2Kgc1QWBoAwzwf8MRpQaKUXeUS6OtbcT5032mJCJGPHQ6hBkJlgf
h5dZ6f/8E/JMttrKFAVG4KwGWGlK1hAzs/Nq2uK1Us11xzwHqEJhO6cGEKy6oSmD
F4VRU2zJ6GzwL9/BCQB3yz6hi5AfN9id3qFv9bf5+RKW6DaANriC5+imMVJVW+D3
M0CRnCigDer+mU9uu7DpbO90NteMIBenpfWT/GkNsjJxQ+ZC10akvqatQhFFGYyl
zaT2fSOCob3qJt20o9gafid3Z5iD3sjZiw7UeQsjFhEXw4x2eogZ7Vsh7iUk7utb
9KV4Uu8i50J8jwiSc97EiA+XPKzYjALOJ5nXxG93/7I2S+VyJNrUPNN2pYze4uiU
cLkvPasmmAwzMYPXmNtXQssBY/MqwzQDpEOS7zZTV9kluNK4eWpHodGxDpQsr2S3
d9kJxvzyAGIcEbGYK9lATZpyZDHPfaurJaab8pXGzRRO/vtyqlXyxh8cVkrLknry
e7wMjBDp/0XZ44xizbIqQxfbFsnMCT1cwl6jTAlc0DaA+2f+wpRzOJTEEE2IHZHl
vvjZ9Cqr8RPfLS+SMSeodSU26K4WxEaUZGArRNgCBwWdvsMh6guTeRztYO33DfQp
bNRq+4Ty+qnzoQOdRWGrqIcutA8l98dchI4poVXL9Ks/rqDYiXIMFlb8bas1dZMd
IWbpIctAi8QCnx2h5UNDq09ibMLa1soUsQcVy56BVorFWl0pnuVm2OPxuGJQ+o0n
OrFuF8XI3FiaZgU8oOL+cHoDQ6ktbsyiJbGZOycguB15lYkaoB3Z+MCOp4YJxZIE
aQzUomUaSmV4HidgJDBf/iWmA+77HpnrzrUBY+iqV2Y7zLVfDGeJsIEvIai++eDJ
cp3lo8cMQnLSuccmh3TXZlyF7SDkDI9Dq0uWWRgZyuEx1FSxYDW7enDRYPgt7EtW
Y4nN2FuFs6Z9Gf5kje+QW+8OABtGi6JTJUAqnnFTL2gjjAG1RleaJQCJO+5OaZmO
sGIltTOw4S+b7BXcnzdiMPYGt8Aeodu+lYpK1zCTIaHY6HZRzNqRASMw4pQjXo01
8DoJmby7/hWSv4WrMcZtrI9Bdt4Xh528GDB8r2jlqV03/agb+D3Ovg4cQyu95E8r
KUTMpclZhn6NJDQ/dKxVFy2+lehZ8qwlAyyLXgmw0+WT8OAmcyxn+WiyCehFFb37
kv7x986EtbzqHHdeLDXVvpOo7VmuFFN9pg0uJaDW87i6G0lg+PIvn4KrCBIlCIm6
lsIiaILr2NKDcTl5wXgyreLNdf1b1OWOWWENUNOeLC8VrxcW5GpGr4Dnq482cbjG
N13PcoqQBJJybWF9ymcEV+S82wvsytDZfVIlyhVBG1f7E7RXXlXx/6mti+xoTYoO
4qYt1z9eqqIrw0FIwuxsKJCqTLtjfjqhcwAtRjNgdkyuZ/zLC4JZT39dkYGnMeIv
+xNFyi+awgv9sbkVnCyuuVU1UY2ii8t6M7Ufq6GOKUTU5xiyI6f5nq9CKTvapZgO
wmbezMejVTkYa/rkcMklb3GQsMRwP0WvgIrJmEslTT1WBqNjoFYGiQMaIj30e8A3
hdBReIq4P3Jyhu7euNswR+dEelWYgw0mti5in8I8bWfB27goIsZGfjJNOKgqTs4K
t3YskNHuXrvP89n1ozQMKZMM9MERqa8lxKAUyf96gwfEyYLtdseD//rUqGxYa/HT
ndbDkhpKll2DWhPgACkXvl05PLwev7LZZ7LLGRz68BOFEKwX5WGYLy2ugaB4dwBE
nzZbIKLTqCeWI+iVT0YA2FOOJsw65KaaB0UIOPcZilvFvYm1qHDsYr8ScZCMQaMG
qlzE1AZXGdOM3CUBHFDtbOkEjF762cHXN6DfVj6fUw66MCkDXoEGd0GG6okSTXgL
vA4KVMfUdAhP6iUgYZXz/ZEuFS0DpQ8fWLM8Qz2V0QOD52/5wt7lsN14pye3S2wd
F8gc2XBPKgimw1oQnJtOWU55sGrkY8IQNYENclxsUQbOEPITCUo6kIBYSvDHdSzY
20d6Ik+J20I/WzOKz5UffW2YzKABk1isvr9ApjlMwQDc9Tw1xuhtnwwb4bVvvLYD
RhOmq+P701fQs/RxxXmu9Imgdol0e6hxQRmCdf6IJbOnMFawj5Vq5MSuFoHUUIYY
bH/IUKL2xi5aZ+Ty+/awo9vqR5JP3qVWvQIWQhDXwH/jWA+5GzG4iXe72qmcl+zd
dGTKFt6/nVh81nOR/89kIp224uBnIZIa/xpoiPm09HG8umqto+Jn+anCGIOvdOu5
jRJq8sX8DZJsJwRcesJELexN6R6jENIskzZm79SZ+pzB7bM9ZDIIO7aviUbEdtEo
lhKij/8CzqwdzMIZZ/dZkPc9rgUw0yA2Tepasrylq+4EFY6jdK8EyvxeG9zt+JqD
SEu2UY+0Vdcma3d3OoZcd8NUPzSgvccQRDic9LlBMCobvfYTfZMkWRxHMQFw8PaM
MABUjyFGf49jcbStbq/+FLiUrWticwG+aZggzYYlAVj/nDofgCm/bh3ExLfvJtrz
59uU8dtchpPH+IETOzMRskeNJi1Gs3+BaPYv0Rmonaj7hFpySMt/hAd8x4iUuvm1
MdFmlL8efeFsKizSyraSaqWspyXdR+WYZKqe90cZxD513gTsw1zwXNUn2lU9RPzm
at9PO4m72anOuD9DLjtt6KjONTA6XBFpZ+0kHQZpLQ/eeZILd5udUqGBs5g040nT
7s9pyZH88HcFPYT0wkHAGuxxYhvkcTFHAgDhcyuqlUh1Q0DYqMXPtCRGmVAKFs4J
wrDSKly7uRRRU00xBg9HkorEm/33wzcMaeawUVigwV4j7BmZSMR7OtbT5ZnikxP4
LslNzWvpD83uZu/RLCIybmhRGEyFcQIlP9D50ZIFL3quJqRbUwFihGHMVeT0WAQy
EUgBnIP6CViUcADXoxmjnRFUo2u0PuQ7019Qejzvd/DJpmn5UYswgeiQG4TmkSbh
th9YvSHdYlGEUW/pAw+v681mYgUtY7VRMLcfOhiSknVGaf+3+xO11YEMMozHWGr3
gsm+0SrwkC4lfyiod11pLrZ+dvsu8o3AlrT7tJi9LF2mwk3jZe/m2WRZmcvgWg0l
mvnrKE64s9P47Qs+E8pKM7Ukxogk0mbBKSRlR18PALUuGbqu+bnD1OGFf9FB4bqh
Hxs/i4E0RP4vBTZwokDU2NpmRjneMkdwJoWjVu7cOPFBuftWcg+LxIbcwyjuhHd7
PHuhJ/9Wedu8QWR81IMPbDnRkucjiwFBj/kmvKy0QZBmz7qu3452R6xqbfVEJilt
xilntaWFWQZ0KpnbaM9gIlF8fjEZimxNmIMq9tSfP3eEfa6ftqb8zmo0qE4XVUmD
90aNH1DxeJm4lsBgIyLzYoDDoQdc1faPiNOIu6HWjCMOYETq8bC0aru9uZOD1mY4
AuQqHSMnn80/YH8r3Gyq9KeAnYF3wHF+5JpsVF0sfKEdSTZEHTMsxoLrNQBggxbn
WNt8XnRh/PulZljoNgFttHLqfNbeXPA072KmqPNTY0XjMkd0N3fKz6RhKVKUtW5+
MSosWJv2T7YzyAISPDVe2koVU7tf2fWlhXoPASdUxcmBjfAsxntk87S3bUkWjSlR
ZwbxLHIHxbcttdyfJ8L5fyoco5mJTRyQ2JBq+069YckfrqzzLa0n0ZGSnttkk1YU
Yyd3HcyiIl10+g7L/D0vykyl8rzfpFaesLYwQcUTNZ0G8GySHuswCOn9C9Xu138W
UHq/ncodZ2SoHb2KH2/N0t3NKWoGztDXoTHXsFKq2IHCoOmFOMGcIfQw3J8pMcOn
JX5upOgno55GNcaJT6cN8ifsiy6TgI9JOiIEUJ07AdpulJW1kYzrReoMfgCSu33m
rCkXa3ZV//a7oU1GZuNkYk+rg1gUnmFBefC8PzzmDsmrFTEKwbqXlxSlRyXbH3kI
j+gXh8Ycj3/OoDkqTOTw4M418I4DfhhHKqlpTt4gipduXgD5ghEmA+k5eSKR7yzO
6IVG8AfIYffIxvp4UefUk/f7w3GJQoZxpnjlFNXjsGXdt48zrMNrcBpTrHPPLRtX
lEzUnqJWpnMf7YBWg80iZMCNx1RFUr+wV1BvJQgnCdlAjoIoEooGCEos/EKiQMBD
ekraQn/mtkYN0j7UwPgCPzMF5KNtX6TAmqPttkFXLLVHeCAs6mrNWEsvMRsXtTgX
AnfzKl5YpySL3H20CSmxqj63QAVXRapeMatcKThVJ8hfx23s/+1CfpEF74r9wuEA
qPmbyA9mKKp29Rtlng2EMCqWE3TI7kS94piA/fcoNnD3YDGmK+nhDuuluTKmatPU
zp+jyRFX+m5C3YPGAE6BFdTmRN1uTwL0a56rsDMST4MmM+HCGprop5KhursR3lI+
V3wRBKfTWL1QNRInLd23VBnkwWmvsUY9A25FUZNLsjN51VMyFcVlxU3VLbcLwJPQ
+I9RInGdkZ7UHMHpCfJhl9XdSsTHHZgwn+yxBFQUFh4Kry/1yTlNK1vduHDwexwk
Mbq0IcZz9C0D/V6WSrbDXOwHUwe9poFudWDmQJBaApf/uvoZ7LGk8PC7hbkPN6do
ggaWuBRl1925eIcUvGn5fn62rpk5n3/FqRyurxVD41qBSrYM41eCScHDg47FWtLi
sZT4OZ1aBJvBlmtGb21yJdv52jMvKxaswdrqz9rebVOhB5zQYnS6w/mnsQTdDW8Q
lTNMBRA9ImuBf1ec3JnuX9RtjHk1MrBD6THqx3oe3Tyl8dt4aUmaBzhYI6iEBuW5
UM3pnPBd1xhoCWlSQ11w24bHyhDA0cc9e9fzliECpi3xecsx7u/3hqJ08fuDw/Bn
QVeJ+8p7d3xm6N96C1nFzbRzbWGH7kCEtvDhqjgIn/FwsuKCV/77g8Tur0F5HyDu
Hnw5owwCwsgehxobRzYljnJg9eum+Ebq/AtpwUDVuERTKmfF1N856oz3fd+WNb9g
oXhgYuIr/fTorJKE42zSnQ6Al7tiggoSRx3OKKDCBeWYB7P0NWwqxlpsZQXHWYUv
d7QueM5Nbk3ccOEtmA7/TgWFNixNNcN5IiRPu0FZ3iWAUxBJ5nFEyneUQABabt/k
vz6sxaU9REC2S0jzvPGzVYfFX8sAv5NOshZMHhyf7tgaARCG/NO96NEq/7CEUPNE
n5AhptHn6Euv6yFRAGCm6Kk108qI+nCisc4Zeszo2DHGvIEOlUjqWGrbfnvXVuwB
/iWeWm+1p1ZaaNkUw283PzwA2WM076xCp1ArTnwSXtTnnO7jrUmHXl9ik2uwiUow
X6BSnfrXQvJZoSVe2Z0uNodbwiFTPBzUSW0QgO6dRU93his+3yfkvWpX4C+/wiHw
MHqJVnpnYKsV9GpWD4HUgq/ADo5yvmGwSYNkkB6IcqGwhxVOHrHb+77+EcqkHG/8
yPoqEGj8M7uew3r8KDRvV//eZZC8/mSv3GalXzdb3xXI1pA4go0wBlZaVIxlsm/b
EEjSfGCvSmQGjLMiBHkwJZIKp3s99BnnB9broTU6FInNpFfoEorS8CU5yYfnDDYz
NAXwPHC8zDBan/AP5ZJKiMqy6aI16QKktxdxQs5EDb8EyvN8VOq1CqVD75a6UMpf
m1qKOgpi76GE/kfF7GmZCRlED1d3kpS9Iq/xBedRjXrtEVO18lNEfSt6FPo22VLF
GqruwEVnNSVDCsyCNPJbeoM1vOgTOLzfHN35tPqbcC4tPfjaxvU/sbN2FUWM5uIZ
QKRuArSv/7ZC/6kdUL/Xds63EJzy77Zmfy7kLLMzmYPtGd5PJDdLNA/ULfMpb2y8
rqHzvfNIDMZcbEEaR+E28hZ+jMM9cfElOrkcbARWt/2naVTBOCkqB/0bPeXTMSA0
77hgV5wlBODGyKrGGZHI54VKp28IY6tvI1kvcgH2uPfkwmEiTD7q6EFvfkGqVxIb
QfKEk7fIeZnlBSQAcM0kP/6Rnyd+lUlotJdbwQ5QDlSl0ZCyS/p0r+3qXhtwMw0/
3ASGGf3FRO96hIyzqRJixHJVIkmnTnLEbeICuIORdOws+v1jfzlb5ut1GMvaNtEW
LofERVxd2vHwY7q5r1YubabbU4ytpWZilr6F2CHXFYDK2uqZor4KEIV7oqwrf9gV
Ye6Q4UAb5EAamqb/G71F1FP6XFjpbheHLMsi2NATfNbog+5nvcUDzH9KjGUTu+pn
n3F+lu8hxwU/j5Ermk6tVlPaBISPf8Sp8vvsbPSloDlW9PiPc/ODkwm3fmLDen0T
Cv9C3Zt2+dLYRy+Bhv3zdw+oxp1maenQPAP3k8+3DZM35G3XoTSPZt7Srj5MqFVm
1n5kJm6H5rAzcq1reoce8j3Lqybnkh9uF0Bt/QjTOG0imStG11VTR38CI2l5CBoe
DmQBYNngTTKzu1Kae48sjbLijuuXDjz24fN3kJhJq4rRkBWyszzoZDmaSvHH6I1b
2v3bEsHRgWgrL7f6ZiGMT9yLcbH/LLS6WmhIpj/RCQNXxoqMBJ6CP8gWvyUIHeuW
pIlL/VBRTOpmFdY9Opz1HzYcLf7DHcor/Ia4ABHJ8kBIjOKxlex9rRqX2Pb/r4uS
WyApb8dtD4qDdm1qm3CquI28HwCb5ZOD50gCkoe3tQG/3R0o5S4cRYbW/oDf/+F1
5P4rBITTJZQuC0mNpTv2D5cQAk7XuYZyqiGRrILb0ulnWG+cbWbuFyYhIclXy2jI
5RJdPtIKaoAbG6GKgffN+w5Gq+gCkqdcDgsWke8c+9XlFkoS+3ft8IdSwfeIY48r
ZThA8piW/eiOHFq5apF9NX7UDkfS9c6ot+XFDt8oJecWKFoS++bDQyZQAGyCq2Ov
UtqxkytLeAixKHUse7bGCvADK6YWQG+T+DxBgzO8oaUtHJOrJZjRF8EZcMdi0CYj
uuI75MWc53H5o+jPuOUCsugV46CYaeCKJJo8cm1nFlXIqgNGszR8KChL2CAGoxhI
nvAWURwF13i5fo9cCH9yxnXKrwgvW6RKDLkxdFr/9crArhTouXJ+t+M1ER6M5IdS
15sRvMvG1EQO88U7JzELjzyTh3s11Zd4azrQ4r+coMOtyANGlB+rUVWAUYp8DYg4
/iVFwRMYGE+jZG2DbKdA62E1RsWlig/FrlgfJEy+n4DBTN2k/iPj+dhUooJ9dTav
hg1mc/+lxqFIx3caClbrZi3l1qt5cqemWhMq9iVcq0PKoYcxFTrvmvhkY2BGkEHV
BsT1JKVh6mHy9BTvfJYBShGPjYwbFbfkerEOlcivs7P+BIk8EBdY0nkCyc0fq9sm
YbK4dlVy8dgI/r9dO2PONAUI3xCmHBmuCfEPTs3J4WflgJgbZLfiEgtvdPJzUQPh
1FdOpBG51uUusfyL7wTfBO3y8i0/2OADmb3sDNqq2jxJNQZGNkioHdtdBbOoUR3L
okHnSWqqUpnzS8hav7jgDf8yS3lGnvNr76iYFFyQ0hAIv02PbjCvf1VDCL8RgH0a
Xa4F164A3JwNiu/qsa4G3/xLmhH8GUmlc0ifnroz63XrtH57ZcGIcD0XM6qBx2qt
KlRxpJWD9xm1FoPIXC+xqVF79l4OxTBsy+vOikaD6mHTzcnlI0rKBSUuHJPbjPFP
uNasQ3JI5dLoCvTTuWo6CDEELpx7afI3aGdwHdREHpTyLRbLoXf8iZrDTllizGpi
s7rDa5dHwSvFMU+zdeRHD4nZ9lHqdIIcH8dVaLdrQ72z77edMgtO/k+lCKyCpvM5
poOzUzslIRBm/ENvCV35OLmj4NhhO2hMOp/tMSXo+Q2AX5Z6Qy26CWWPzFj7LVaw
H7Lrg/+7XuxEU57MxLmTNOr27sqHTLsV+SK4fMpkFRRYD577JV6RsRup38dq2Rw6
NN9mxoanOrMS4c8c2uaXgwx6ovwvgRtactqeE+SqngGRirEwjPuk1IseQmJxhq/Q
4+gD6dBV04JCMg7hFeu+AS1tThQl8XNo3ESzLuJunpYQlSIF0xRiyJnMdxOdrEsG
A0mYmyXF3t0ihlLEuGqKk6ElmLuMl25UOtPmOBS7trsKAIBxfID3n1aZwPSzIFzh
m98jVLZOBwR82+/umtwhdijDmtSMziV7MdPR22nKKRIioJv8GcxAn6V49WBiTO5u
CWlGFuWIyQQzhTJryFGOnqJm5Yg9xEe02NklDzYmhxSnwN2jjTQcIXOwr5B0MViJ
PuFWQZPlYAi5OLocfSDSlHy0MBaQyuQMDeh4xLzt+HJj+cGoVjUNWcJR5ctOFMVu
fJ0D2vO2nxZmc5nCeQLar041b0LK5Auj36D0o+FuANoc92KEVo/Ohz9W8u2KRXXA
MA1SRiuxDfiXSsQ5nmAi1qoMpz2mwBGVgAon5IZ0gMeZRuq1lq+vBeAI8J8tRCMw
AxtQxijaVEmB3g9DkuSGSox/z9Rj38Tw/2/iIGh7RuuYVQV7eOqouP78mZLw1tYC
AYJsFG9RiZ7pq2XjgO8XKamGN1ISjrIkNEyKV5Aw6+4MFBJosd6ttuzprCfzvCZ6
nLAj9zgplDjvptihZWVZASHqGVUuey5LcCSbhfGlszCasRZ5TB0tHCCQUG17+YlB
G72it3+PDocOLGV4YIzCk53pDmbWODvUzFGRq68lzvXZvfTyA0ePf51Y/nnr8mNS
Yn0UrIi5D0pEG8mNTWdzjfOJcsc+quJBabhDl2dDRqsLQIbBrJiSbba7d20ghNKt
LiAZ4FzN6WgZ3ycuVtxIUUBZUr7oksGY+4fCAbvDXK/RJY/rMi6rOjCBJJWga4By
6O8wqhVLQZ3b+MK8ncXyFmm4MS7K1511YYI1X1NkveGWgAzJfj4AGbfdupS6gIpG
d/ZuJTMn0f7QDhm306EgKKlKd1IqUskz7DJBIXTg0qJxbXOkWZlA36jxgnxchVyz
j+NYaJP63QkkMhLzu30cKtAsrGCHBBTSr4SRu4+WvPYqq57JmDxVBnpRzfE7ABFu
AUC9ASYsQ3RGpQkIhEWOYMU/yTwzOtjS83wukBYkfc3NyC8uyVSZ0ikruQHqpVQU
Ck9+1rj71+VbmueHKBdhlq1E9VCWXwM1KXU1O8njW57iq+8yBIb8gT2HRliGrT68
U7CEP1Yjj0yFgFfYf2/EblJf/dGErTWVeNhbFq3c/pIB4FqSWcOyDbnjEKji1KOC
oPbZ0wjp8ca/Ix4jTP2F0NYw9gofR0gn61b1R3pc7fXteUhvhbmup5guvcX88qqh
NL5sUMpKR1POnP0I4gNa5g0FXn0I9DVXUwSkYlHMpjftukLhUDdHGr9q7RTJSltg
HzmSKHpYXw8q4kuPQHcwZQO/6TMh93Xn0BuxDyAxWHYBjpgby6iDNRrizo7/QPz+
pEi5x0R8hn4lt5Nva2yD8FJM9VwQ82lmDEvlkJkURt9roYn1WHJdSzW3jnXZH5So
XJuOSRSYl41zn2CB+ChWBZ3xBPoNHgN3aSj8WuD32v20Rj81RsSjkAtnCx89X6Oi
LFGwq1I5PhuNwP6C5DCEfaBGd18rug8zlmZpJc49EaqyyCEGOjCuZdh0QMDDDYNt
rVeZsalOUCat9JSkyYFOdU+hLc5nHlgcRt6FnLlhpQXnpSYzOFI2EwM95wW4Pyjx
76K12oQv8Ui0LjHXsnsg6Fx9NdJaRAEx2wNSBJPbuSxT4UlimzY5inKiM1dyb5t9
6PECYd0TmvBAKRDzBzhPSg12NzaybmZBgJx3C1iXIsukndx4IoKOsSdPmmV+1/mz
ZH23SFLPT2TLVmaYSDiDUzYj+mEO2blxFenNLcPpgHMkywItH1IKIOufjIWbskDd
Lxc95T7AVmgDSUKkVc1zv0OtP+BEcwM0/TP6tYxTVpc/38xElq4b007dv9dh9LXa
c3zLPdJ2BRqORfLQRjGH/68GhJdn2flT5JLXA89ZcmgXYuL2ue5FkYb6nfJ+8Cvq
8HMw9tAM6MaCv/c17c7WzBdHjE18AR9PZHBFJguf4GhdPiw0V07bFPw8EI1++4To
0zHuRpI3mzP3OtLdznBvlJRf+pO4YOgwns0q4zRrV/LUm+DZEpYLSJIzdZgfwZ6q
T7UcuRz4Lim/lxa+5qcmQCA09EOtrIkXmOZkSRz3rcHxMXcaRVZyMyJMnFAvJHbM
reKep5xcb2ACITQGm+f54K3p78mxDBYXHQ6Keh3ZguENYH6YcIll/wQJCs4WdMaD
kLIaWnNqIDYB5ovuEem/TjlAgPLhjrGcd41xdry+jxj2dnkqCNRGxZBwHBa1YKOu
bxNXYxsrsIogajmdc2+pnNnjlWcREO3tkpo04pHydE4SezT3/DgkNlnfmp5kQVmP
NjjURNQtX0loBwFPMoQGn6YrVkpD8cuBA2gaiYAi71X64YifcQuSFBSsZjp/K38Q
i3/twYaRoRLK4TmEI+X1KLnETIs4l5HrGTuB6bi+vcUB3Ujj7tdobwz2B+tdjZYW
7ZC2kNNpU2Bqp0Z7UzNdNABmMA7KFkUmEpvpWCpGKyO1Au1ALLrA6vFQwK+NJ0sN
d4MX7onZmNfCC6wzf/rU56/SQ75OO3gJXuMFP8mFtmpodqN9PLQxMwa7xSn/mzec
ZWk1ZrDjTdVREGrrqUBQSaZDcmM9gOUwdfGWcnT24DO89CuX5+SV8/0WXEvuZkcc
Zhk/mtJWB3XS9wZ7ySl/sT6lhuxPRoB8gZ6oFNRBqEUOdZBPC28uAhivtqTHWFLX
El0n1kNYjEYZ6e7QL/r3EJ3qfQHynGxZVtORS/yY9EoqwNWgpRHOaNkV51P9/big
AQ23TWwKhDSCmDNtxdKJEbcJnXfJxJMo5rMZy3YQ3roJNV2bwRl+QN54stPUmtAI
1jcHZF+CxzeQxpG83GHbrMMe927EL5qEhr7aARKgvwXcli1/pp4Pf/0zJeVVDGDB
IyEI83knxfmXYsZxnaW7PlIiVdZtpKTkgnnL0nFGY4zFiIUBgftPSoTVeOakhEu1
VKmAmSsM0Ous4rndIPRzRV/oDPjPUnFCat5xiIiLNgMJg7enme1Z138gKaKOoloU
kAc/GOjfn0UH9PUI95nHgW5KKqwH9VNCfQ5jfwA12k4PpL8Ec4/NO0IreA2Rzjo8
u3tAWOawjYOGGZ/vjwa6qz6LaLv84jPoVu+6jbJL5BofSo/57w6C9ch8oygJaulM
lTE9OdsPpHsIInwgIyhMetGWJpCjLpmsc6nTldrDLPGU9vO8cLn22IQCM18bA0Sk
p6SSplr9DMGIQX8lkzKnMPP19PZmnecEYqJmpiPkrW95sHEbBBV0b8YvFFu8fR7U
1eVSVcABcS7cCBzTSUuR8GkD4Ft1Ha9wBADREPzklq3PNR9VHlg+vq7xY2oi57vB
3GcpuoAA3VP5mXl2iWACkciqHZFWsNdeipUoqrQrnwDvmkSD+6qffxlCdg8ylYJs
sUfx/YcA8xt6XLVlTrHtHYdfcOFxe0V7JSr1WrtXX5zYuTBK7YybJKjghbVuE8Z4
S/lKmdydxaDmCyZcGuHT/rAkYmgZgQMyUkTiIPFT/uMMGxKucNHmchgYodDQpyxk
+IDgoyNu/aXxikXA3PnvtRMY/1Jn2qVsEQVSOpxC9BXhhocdu9l1lLytGbi37AJE
qkci/f3ptyLtLD3sT6nOHvcvuRR5U/yqp/DlRst9gkXsXcSHfvXl0u8CrTHiSA8e
Vko11W6+h37S3ji6yjRYuzd66H2pE2AtS4s9p3NFDaCDAwSId1i+Oi0GgMJB2wWm
qxAZ7CLVGYpu9dR7fXfexs8tQ7hAOiZX2pq6uhYTOEp/oRS1UH8DsrPsIqEqwK1r
qHZx0AssvSZIEbn0G6BVoujaKKLXfBEu06XXOXC7gMFOz5gZ7AW0v23CsLqgFJ0/
RpBshUdXJlbmRIv/guS7K+I4W5Pl/oZ+wFdVu7bBmb0t4zWa6C+F8n+Y8f7fvEG2
TgQeH6HoT3SQNe7+5kXJjcbp5CFNHWQ4f1F1SYfisd/BpVYKXTSks55sZzHUWByt
hLku3k1jx1p/rKG0OITJEUzzTpAMrGu+gzGCPwl5tRFZ9zNZQfqiUZKlWaRA8I8R
gWwKe5gJuQKbXja7SSlFMhPeU7EzffeoLCsUKIp3q+yu+dBQV2/nK6IvzXrmAyp9
sKjAMX8s0EZYEabQyFtaTuQnVQqOyPa+C46zzRq8hTN8rQwiyg466KhfWQIL0x2A
CqEJHXIu1H9JOXU23dark4daDwAwtC/qHwiahAEyTq+5AS0GAmyBeY5NgYuGhB33
d4tmsP8AYT459tNR8lfAyn1tYjhZd55g8G6F+f+/4ga8axhYIyjy8kgaO45kK0iU
1PmwQ2TGamHaNCHY2MHlBN1VKD2ObzLtyBfNPT/PymCClBIqKnJ6sEdppzmgGaXR
NXDk+pMRQstsaKBPDWtQa441UuCSOVHCD5X3IiEIoPEfxMDu7Hl74XIYFXA6LOiL
chm1hmm0fkclm8wGSqp8ECQYtmebneb4JJgwPRiZqS9Ro/LUdM8bCvpXdZ1omY9T
5ZxkPSbBJwxoZaR6ff5av0H/b4st3KX33ryKfh/GPW3qRrlx1oKsc8jOLsY0KJ8m
pS3DyP9OJrymG8ysFBm2plAKqUAp6tw2WOybKIJj/djSCYrbmqELFCrQC7IR6BYP
PUdle8zPnrgT3SIsk28W8aGBnk04LSjs6gT/wXlldLoAfmVK8xSorIjUJRpwru9V
9mBx74dNwhWNxwOAK7bX6djZ46gRpN2XOmEpeyEQtR8Eh12Dd355x+g8njyz/jXj
wl6mbEF2aaz3F0N2YjWsf4GhzsC/cO7NlxggmpUnk0Lhq2CbgZFzkJFAyk1MrQIs
Ij7AOhgG8Ycz9LFPItmCuPR02aqT8bLhrk+Z2ZclFv8WEMUGKthuMyNpaduff92j
E/9nD9d8xBsbTd/CyqkegrHYI6MlgBZI6vr71AIsxv+KX6tmP6Z90jpXQcw40gzh
Sfk1d1BGJ447i7j6DPFHTXekNYZxC46DJI4GnwPPrsbq89JK7Ixaqvmd95wfPhGl
XXF3Wn9I1aucvXc4FJZMLKUwHitR9qRUQ6Dc2EUoF3wzBM7WWrfmddtzApqsMZYF
potxpU54qxKRnXvJnVucDJeMRFpyQjCHIC2HWBqmHc1NVeMCWT2oUeObkRTp/b/2
vn6bQeJRocDr7XPBAQfJNSameoS2aixAtot/R0eF0a/j72h7BGLdeKnd3XwuuP7s
37gz2Ce0iQW82JlD1KEcez9RFyW4bIQwqBQJCTRJ7d31zHyuexm8Q8F3hByTfjDu
MZwEsEvuU5EwOQi/EnXN8LsESwI89B6JJBJ/c8ikMiL45AjLmsdbX4LxZ8RNREmW
BBlwJVMPbEgz4ai2ix46erSmLwam9h7cvIgvrqpAqTn6YfcDJpCgbnmfdGCVq6vl
/pZO8By+b2l+oH4mO1DKSIMftqYETX7rSdjtqQUs8JZgS7zHs+xmc4ix/k1SIBoB
1/NK4eCe8zhb/soqsyZCDKyrPN1wvXny/w/SjuANSZE4ACG/SjU6XQQ5+8+vM0T3
LqEcb/C7z2gIBTpf2wivCUGV3Is49DL5e7vYdNMVf+Qdwqf/a+wMGKlV5IPaAFzN
x926LeZ1IXET3tnw6GeCZVuOcxkxwPyRlRaflF0KrSs28NsQshtsutslyprtBFRE
M90B3bBuLDrslpfGSMt8ztBYVC1u6+mmlykUgX5Tn1tU5hQhJlnT5KT/2nSHlcIq
tZHpcYLxjszJy811YJP9OkPl1YQbg5YA9Obv396ZFkv0KEqxsxB176MAAKRZ0zvu
GE5WGoWDeU75/rhS5XsKSX4qgrGvwMAexbzmq5/yl4XIZR9FsYhYDZ/Y9Azpue81
l0hSShX/wjEX469aLUi+23EPEZSvrtZ4W++ZJLoal+Sd+9t4u9lEVwL6b03BYRJP
IevWCa3u8xa9mWI+0S3LjdG0vZ88IIIBsfl6oqro3141qXg7H8qn0YgDfaW2T/oE
zhkjcHQxGkU+wop3epuAHrVm5NmjPcqm7edPgOoGbrQeW9N/2YrH3KVroxYECDx3
FhHhirrv1qVTykid30HGMrGNXK+0JOBQKYNFPWej7Zb1KgOk4BDbHaAuz1eAqp0O
vkWjFNDi0OnqmTHBRDr4mrlzYU0zAKqFXyEsQWkugLSDikgtjN0a+AkajX1ZLLcG
BaNUhM/NdcslnkW4hMP+A9A0uUL8NKeOMfffdB3hY3KkWD/REU0rMiHwHHynRHel
7XjaRvHW2NdRXXCeF6yIGYqpNBgSrPQ9Y3H9QORrJa/MCy2CkGQMiTTj1KTYS7Pw
PytpATMx+Eqh8QHBR4YTzFrL4M+LaQO7vLRFTWkZO9mZDDU6A9sCWnGxnuQEGT8X
uZiloaQlnc3UQse5IMoywWOldjsHBASonnSFig+/XcOE5g2yMRi+JctV5YrrCJno
P0qgb4vkkwf6AlGuLhpv0rpTI9rfguTH+9f1aD1NyY8Wa95bKV0Oi5tug8Gm0R6s
a2OmRqVCDLGAp+/br1MGzpSCALtfllmGfZRabufDsBJl8HmZxGVRG8qyCfn3yqzI
zi1o2f1WHoqzZ0lmgrwkqp7T2rAb7sfrFrcb5VrWzy4FNtI5YhEF2oZza50BC5Dt
o8rWVF8AceY3jhs9H8ApZO7rJkIM4Cn3k0otdNSsAD6ykrjJp5ox6uiF0cjV/+/C
SoZaMOUsgp97q3ZpzkrhwTi9k7cMpRgLVPCXR5Mqvbct/COOhNKeVicKi+Zz4Uhd
9HxO5j1TuVfvo2OIxuNwuQXm2PGxKEidDnici9dLvQGPWh0I28SkiBAy5x4Dqi7/
EE0B8XUz3Vc9XqI+GNV5GnjEwPwT04ExI9mZGRsobjYbqBUmeNqB+iMwFJM4x/m8
D6I/UCW34eDYuZpTAkklK6AFvsspilaD2fUej3PTEuHepHusZDLkKmP0IVmm/if+
KF2rx0QlFvW3nzwVsAYOFYJpPgLVVZib3DjGcVqjaXuGFJP6Qd44JV92PtK0KMuo
fczFLs1/mksyBpLNEqRuymQDNiP6q9GVbvxJtXwWuEInVuj6DVrr/U4tIU9ytd2t
A5Jydx+zCQ7yv5RsMRxT7IAV0brZzZJZ8e+S5dFaBlrWVGv29iwTML6JcwG/3AgL
AGS1G2mUkXsAx3hSN1Zh/Vx9vMe8EWClMw3h5G6Q6c4jQcgrSe4NGcjF2rQeWtzC
McUe9J9CMWr7f6dvgoA6jBsxXmXCR9FpaebZin0nZ0rIvzhzA7Nmyuyy3uMCFJ+w
O+AVCm1o/YQhQ6mjSuSKKURhoD337cvylYPgbDPHqc5pq7eSextVneezMUMq0SBO
8asElQ5EtG8CBlE4BbpHCU1ZonQbnZetYuD+59lDj6ziFLaG8KxHoAEryKwVcJS8
YiydVEnnM6PmeeEyoCtR94/S/NEoxHpKaQESmBiVqai6QTVICiJOVk2WM+SNZ0pK
eNmsMPw70nMBAPYa9vtpN6/mQG4Olc9D+Wt58zG6FM+EliIkHy20LMhf7hWqTQC6
bQoski7sAGcrnSGmJhtFo3t91v7YoPZgUUVAyPn80fteDMkyqiLiubYpDMiVTCHm
iwUIs476qUxV2bYrygLBadOmorx104a5Z7DU0MEJ192ow86NOQ9e6JqdRQq+svpk
pktJJ7/WBQWLc6jMxImja29X3S9p9uTp4s43e8WERwzzxBVP/m8dAsv1u7SJIiVj
RER/6pM7HVl77UQdpquyzWaFOgLNixFu7jOeePO6BSSe1nqALDs4NxpNyrqPtkdC
qzRtqM4JKmIjujmU1pbjmvwnpwksdc4bZ8boNmBTj6wMLn6gV2HH0ziV8QfDNcKB
0+I8dKEwUKfVMJOgsmwflpFbk/WsbqcVJ5FGJpRCYvIimKLyoLsSW+FP8aCVhpNM
j9m+uQlkS9gpowh6i0lq0OogfLlS2gHRut01mT0izAGILfZcyWXc1LwEE9wk7eTy
SKjZG1WecXYF+P6xNE7HsfMMYbR2kxkvmwazItAQDijKo/93RrMYtg51KNajjyQY
CS3Q8eUEdY2SwAOe7DrOLDEM+78d2mYtrynGReNoANCCPjMywTpK0irWfR/CRGI9
3gelYxjHkY5O7ougpwtpKcc1hpuWEhylRIV3s8bo5pwFN/SgsTylVOZ5CLyXbDAf
uXc9nvQHyzPj1i2OX/xRx2WrNHWLowv66WGstOyQKvtjORBuxMZKe9zBzCgTV///
CYvtmcwNaCgGMQ+nE4dQzz+ocQ4ZMTkiayDR4rcJj9vOVxPkD6ISCTHN1J80YPSl
vFo8tDS972UCV7B/AqpBQFdLoBtTeoPNp1mJDXyO2JI9ss14PKbklzM84fspY8vH
29/taayUg69nM0yLJ0ebnr4UBQG7DGXeAsjgA3gOzXvmBfWF/wfgsTUUcqobDcda
y2+nYaO2SCckRHqLyIQWbdMka0pIpajINN48bm5J2duTBiNBNSztDe4Qnu40QwUG
VlUKfsFnVnnDFpf8pemoMrxl5eBakw3Mo6R0YMn4EILvHfyq9gr3xvQyqwaXZYi5
1G02tTW9SE005kTgom0kj6i/RPwE4h/k6BLyG317baDCx9UpE+BjXc9ZEjUK6/CG
fCFEc/uoTQxcf4EcwY0EJj5W2Db9czjRtXzFToMyaDpVhui4h56cRHk3jW0mt9q/
xhOOtQ7/gX0/8dgVuYXtBGkgQFPybi8axnOJiAVPlaa1AjyBX5AQ7biNqrJdkzmY
ZKeEMV9s4HPVWnc0wGb/52uZZPDc/ktbm6b2G+BL2FqldpXis0jG4ABAi8+cfBq1
9Ww/wd9eLk3AmNJM0BN5UdWfhcSJsO2C/ZUykuOyTEUgjEwF6cDmj6CzXQubu9zX
QmnSzXfIXvkdxHt6TA6OpfpJseLKvSDdZF3Gm5ch89xPG24qjB2ot2uRj/ASXill
9qr6Tjlay5niJnZOhzflQqP2heLE5O//qiyp5QBwe+uoqXqZEbZnlpiBqEa0Vr44
IIxjETWdGFFAadXNNndMCogqPMkFi0/E9HG6/jB2mnG1TIllaFVkJKv/boU0u2Nt
mHk27NEPCCbDN5CQdRqvdnAwwY1DoWRViSWdudBrMUmsFxmNV7galLB/0Bsb4qEb
nelfBzzu5gCc4e3J9hSB+jEAwbAsFG/0ZsKxJO+HOrd5Xpthal8vmxBdxxsdnsl3
ZUyY1xrXPGxImvDaDbL8ewzz3tS6GFAjSjOkgtrX8GczfarXFDh7Ri2mgpeCZn9N
6+vvzEf9nV6ecqIRT2CDLeC1P/p6ylX+IVHllITmcqDFhXmPIhVjF550gWepy1te
wxWp8WseVpJNMl+YQx/JIzFK02EOMg/zEmA656XLkokX0b9dbrBim6lFYHKzret/
5XkVAJE9WkWfrI7sy+N5/PJaAydoMampWYPl1RFbrle1C9XNszWx5tAeR5rT9wa5
H1WClSjZjqPg8EHpxclthbLExjlfsYI32Cwi8f9berjqSXpWekEX9HrqSp9ekcsf
Imx8O2PW3Jm94ouAtJhKeR/8O5eh94NrRY9GcwGszN6mgrVOwHab8NL00mz/EZjg
wUCMKMWukmy2kqVIc6TQ3uGJucV9V58NIiKu+24MOzLdYYfoOohZiuLzd/sn/k9u
BxW2QdQ7Eqi7KaWflvPXn69ZwsnWDRCmfYkrEixq/KVIPI/VzLgTiV8HxSEpbYoW
RikFpvsl9NL4yiURMOlAYS+lkaZ9IsKKre1tvc0APGrtk/Nwr8CWj8zK8eTFlxt8
HlocLf93PZBmZAkxon+8xp+h4ZCUR+Fu8lvp7E7JX7IOrDjRb21X1wDW1iY+8+Dc
EohTllT1obXO0y7oO69qHDfwVAx4ce8cGVaa/oG1xQJ9iJA/pkc/qOVhdJTcgXqj
vbOlV9GodIVW71U/TXoY0zONBm9I6S3Q5OkMVXEqoMG9LexcSwb3yh9r+B7jnoMM
W8Uj1HYtwF0AXvEppf54PoNVk0BsEgNpFq3Z4Y6NiHLIKVrmVKIqnICy0+kAhme4
AkHCFsfszpY0bEL/h+XQ6XdBmUUxEABV4uXL0FBOuC4uhauEqlqIDr5/cL3PC51X
rxsmIQ38gzLQGfTv1hv1+noyDNF3zcYnTgmQqIFmtxa50Gx9ghYtJU8IC3u4f5ev
08ScW3D42+uOM3KPqvhB2Mc/32+8JyL86Nv7rDcTLYktXA6nwbw4erWjoP/1E2Ve
lK/3U5HBkZdGg3EUBYyjpXwcv7LxO0sPb+n7MUcUdFWUC6Lj5bM/Z6NGFTdK8BKQ
y/Edren/hFC5s5GrjPHl3nqpSnqvJ6yX4ZfHLLEBLiC5ETGKyaWg60k8OHUuEjuU
KZ8fuZ+M8GEhkSy7vuv1TBbzyjfgBrH9SorYc1GlicfhC0Zjnuuf1tDmNIiha+gw
ttBLa7/jZWUXJCZLiB7fscAnV1esN8OI8AX/1ZO2V48DBllvrXE/lZpMQB1Hm3wP
RtcivHgF9wx3+OINlOV1//0Kw8+/sRXEZbQdNueh/Okag6RK+93Eo2fJOg3T/qeZ
Cra8crwgkF/I9c8Dw2OYm4NdiV/CyvJpCYtDKYFRh1Q7U+ygigSmXQP+hYIvqUDz
C59wjalEetkk0bkYsSDCYbd2zGfeg1CNWuNtW6STG/m1sSEhFJ0gZJbIhR3wlHbt
hIITmYQfjVdVTDrm4mL8Oxx3k8pMY9vDLX61XyYtTduPN3MiXJrTnjuhmPFhzMb8
Nj3PQCVD/PLEj3IfzLhtqiecRfS25r/tEeqvZQjzRrfEOr5C21hwaZtzKZal3DSK
RQNcv0/B2vRfpw1NYz7t4whhvjkjkOrSrK1F6RTuLCOkiW2csSp0PVgE4AUm+Mus
TH1cz1pZP5wkz6VfvottvsBG2COg9NPQO1hraQ0xU41PZhVNTbaYbq4wtQ1rFDQa
v7kRyYGt02wd5S24WKDjgtTVif7FjN3N9Pf8EETmGDXAq2y4QVAsQ5qkwT4S7O8g
icTsuUyOafTVKJWnliL/F98EVE+CGqXLJDxrCs0TBZXaIjUyVoxpRBho2K3hoTfn
tgTqr4aXHS30io17aR82S13htJuMGrCFh0pdpWY/syPZDJLsuAyvNytfIC7L/PwX
qPO3vvZAH7IYTbtRyme2myv0FqzekjyE497f3I9Z6GbOFHrebbZw9sAvOzul8qh+
gYpwlifVbHltU6ryQMmC52SOveNPhHzVZJ7DG8rs3w3IVHlN6/K6RmQ0+hazyw4u
t34MI8SfGnyJJ50hNpl1jhqYmjDcJ8POYOcQF0e9mzIaruwiz+GnMh6Vj/FZd/n2
kB4SiJnmObPp4HdFbBtvLS/Qe/gg5iMpon1++ES4wd8kc1eg7VTET6cyfn5XHus+
NSD17BoRcdL8K0K3z20eNas+G0i+PYq9gYDa0hPWusc75caB4K6+APfkEh+okuk4
n8OOeCOAoq4Xm2PTgd3qJya6aJGRD+D3vSkALpUZxuxvUw0kz6hacHxZTpSXrYmp
ZrRqPGdByVEzmW0A+lXYMolmoB/s1qAeyQWdYz4JA23z+ZNyFVM1jMLy1Fjdomam
Usi53xS5cFJ+Jcn9sAv12Z/lWL/+atq9Lsm6u1v2Qt0z5ijFAEsgNqqB3JiFnGBQ
v50JKrGOn5Cbj8H7thWaYWdLRrO4m9X7KtbQm7ODTvlBRQH08txbqofsnbPfIXW8
NKF4I5RR0BXxB4vq+z1/46HyaqVC7BQlQ3oglygBvaEmXvTSWqjydTEXlaR8wzLh
eeXD6cAALZHiFrDMAN8SQIzi9xMG3Ihuwd3KWzMGIHPVZ7/ZuRhI6x07PuPeXUOK
KS5lC7NIeT1QIalko2Bffsq+CrrOgIKF2f18HTqebAcZECIIzHAw8uzprhX+WK/l
8s51oQrXwia1oD8joCu0B0mXMkseKJFfO1+0K0Et7mBQWvE+huE2tLkV70AUUc6e
O/nYRNcQ6vT3WjaVKThYNewviZ1H9iMD8dVK8SMWVJ5jMHnmE+4ogsAT6C2aELGc
cV+YvfEFUdjWJhA98ub7eogOA1XmGfkWSYCfRr7HtCusmStaw25UegglroaP3b4G
FJeYI5fyaLKHB28hM6kNhBwPIktWzsZLKqFNfhhfqrC61mEBj6gTYWjq1FH1vlZg
ilYOSK23be3o/rozC6kc1TORGcnukiTn57rC1AKP03dCrXEZYU0ZgxI6MAdaPVHR
WQap5oV7A/HoL6DwD4OdmASr9OVN5dtbWDlhqoBQBESbYLz7Yyst9pc/aPKhrAne
eRpaZG6W15KDpj0ds++kX7zfS5e1uVcEEVLpOEKhJsu14nZS5McByYNo9RcNvUoi
8LEbcT8RKDBLKduFqSQp5+qyTbMx+OMeNNDWGai3SkqvBra00vdGGXH2DbSpxd2z
T0CEaSlCQKwKNFeas1AVA1PyXLPgFE8Ou56rebzxmaRhcaUqsZurNoIaVcXbZMmg
w9cc0mdJuL5+wqgilGeyTyXtLjDk1Q6KaaP3YgjjHDUnkdVJeC+4ZRo2hvxi+Grj
3UoZ1lRbvfrGJ9gFWcb85KVUWvmSpmnBhVLPFxpsALUPJAE53EMxXo5cyqIafKyP
zgR1kMOJ4yve2zcyZbDrT+x0sdXK+pa21AvNRZzx5kGnLUtwatAr26VafEgc1ZzS
URcFlPhU/aFXWh/ScCDohwL63CCkv28etxkMFzGkkq0ZzRrxztjAVgKlCXqeddTN
I4pwwxeZMesBMCHH5ZdPX4YwhFyMvaaFGAwQDB/UkG93gGwYjvY8aKDHf7GwQibM
O9vpaN+zEZF55gGARtPNtZdizOGIPVZfV4JVvM/WuWUYu5Gk9u3fYBpGB+1FVvC2
O5kyQ4so1mH/agWd+wVNsgQrlD2qVzUrvr+zV547h8LDwz1jZzrlZeWhSAeqhQCW
M/wDh9MgSEdCxA0XbsGI7VeXwHNj1pDuGrys6fq8BYQW86GpGj52eSG9om/sjcg/
o17Rz4p8ru/59+90NBchCqlKE6OtuP937TNOIj8upjYkIsd7Bh9heDgPpzIytfsG
ltXFGZ85nhF/XMsd2Dy8wCfsfa/eOi/70wX4gHx0oi68rkD0P3nSIysXm99Hjptr
dYFABgbdcZJiGg3AQYybh2r/R3SRDCXEOHKBAa1yxa+wK3TbCeTr9qFUHWQDraTf
tjbxXzXfvKrctf1MQ3fcbXw2UvcG7FhFe5oyrb32gHYSv6qcnSbgKNDP0o1YMxsY
lU3Mv+axzu9iG5u9llp4EqK13eCD299A242talO+WbB9wZrbSm1EjZEoANvanvk1
lC0Q5bsxsZWw3N4pDIW83B+vhU2jMMp+0c1Lf56lkPJiWYYVfevnKY6rukF1KMtK
+i76hw/ApGjv4g/zN3NZfxxvshGhH5Q8Wwf0jASb8mJc3igw7azr7hDN2DQw9R8e
y75Wbwu21f/H2PohJjFfII5PVuZ6eLJSg/qfVOATXQM2hwRprBTYVSrIrg8xf7mJ
zOIOQUtzhcWgvaIFBvrjhU6HX5FWzF6WmQZ+HQKqYvuPA8tXSKJVj2jgfVTYitvZ
TB1fxPWLTwf6NFEwMJHb3d0FVpFX0nap1LWXTnqPjMma95W75FDZgpnxXDyhaH2I
PnmEHYk7YRdcbIpaalqlWIAe0P7AuCcxbsON9TxFoH1Zslv69EKrGoh15QA7Uf7n
XJL0bugwW84oVBLuj/nu16Pv/4ayNj/51NHuIfHQmy6a4xkSDsLDhKs6n04iMRjg
MAbe4Q5xw0ug/Ybhp1ltDwLO7KHBAyiRBq5Pkm1jWlaZcbFabpxATAxnVyeIeB7O
lste+l6nmcFwTmP/5PVMtE54ZymIcAInRh/JpbrRt8WUCkdPP+SXHzslXwdfJHXZ
Z7nKttwdCwaxo/PEeKDedI6duCzjf0AzSCHuTf4uq5Fg1lMEmkYol7g6A5Kxj8x6
VZbzwOjm8L87Mz9cskocVsrQSpSVtY+4VN9NxU0SXshmL5VJtgo0Z0C4fsnlWFuH
BNbAjqOtwxhyaIu9+BrqNEt7MOtQXmGoiC+jbSGnLl1xFypH5uU/HS2RRyTLQIeO
xeldlNQGhE0YO/PrrMM738hF3j5KtsamxPXRsO6EvIcW+FdZCgDT8mX8ZaJvHT4R
4M8hwUe4bWZ7LZ8p27/+NBJ5NuROjTg4zM+07T2NYzXN2HqKm0O5UJ784T3uz2tc
PyEClE1UtVSypmho2CdWOWWnTa4oUv79ZW3amcjFU1hONMb83hHiLwoeqQAFFdT8
q6aCd2IrUeJGMd167HqMV2nsGq1ObCyjrUZD75Ho+drH6ky9O8+9ZV+fLBKmlp8p
uR7osAJgeWvOjPUDhddBvWGawHvi7QzooJPEIfOGYUrD/CB/gSGIatGxyO38RMln
RBCdLDfRwIxr5B5IeEOPX6mStx15dagxOpD8liRX0BJEQhL0psrZ5qn04y36dhEe
HfX6bFD6xtt5yYgFazuxDyig2ttWQBS0VW8Eg2j/Hqkm/JFU3lDSkCgMQjEmJk7P
cMCWns9XuHqg3RO9XlBdjGUQtF8HaCQMnFP1W79To108CWonx4YFHxMs20hCuhuM
cbxBBNcU/G815HHhoUQ/cV53Eli6y19AmHa8eZO5SnVh12DyvLNchrlh0BxHwQ1O
k2YWvU4ecECiWxV0skrkKh35ObzggdEPSItqltNpQCzJX9FUThHClvLNSqjC72+z
BHVM3zllTKqA/G4EfW3RIuxlgb63GyfaX/Ru/mZMeuIh65OS2Q9r/UvjvEEdbmw1
AOpZUaY50YCLb6tPi95iVP7S0Mos4QmB6xxkVhNNSGYJdCCHloqBDk8HgOe7lT0L
vtir5ez16OhOB0LiRFMCXWjT7zGE9k0EUoeqTib2DeKQKcVgTcV7ggK1eHj6/tM0
S+V8Or5WwpZH6puAK+W6z6VCUVFeeqi1lpu0RlmDJ9XYKnnexWctPER7jIckTRc4
0EkVdtbYgK6DF+slw/j4xEnjqRrZorXR91lVsi8yBgx1kVM7ZdIRt0BLLH5jzSm+
gneuTwez0pkgIynK3USHsMp2F9J86IAimlNDbwjsT4cyAR3ina2ySDsRNKXfhnrV
DmzmEcTwCQnMVq+ELu2tysFj/Tvdo7O8w7P1pLquV/L5KjMARmDtBVkEo9aB/bXe
+TjcOt5/0SreRtueFDw1zk4gF2tqY1ISdV5NKDy/ZOBHusJ6C1xNCPDxw8ETMn6f
+PapVcxeYVyTELTzyKBEaSH70mRhEYIJFhWFVt91eBqv9T7FHzWJE/QxLa9920iA
i3xi5VS2Jj+fSJdz7yU3gxrl6RuHRm9ITtmfeWUH83mIyXO7K0nywRT3s9a1i9fV
qUM8GYz4OsuNC6Kox6OPDvxWKlbKk9p5PfFklihtWbMk+qDUcD8ss2OC7aiAWgLc
WsqJhACHilwQymr8MWL4bPZjcBgXyhHQ1hTNcx4yiMbCr1t3vYff/JigNZ/ht4Fo
Cpd4Uud4JPIDG5+14RfMOhB/csIz2evEAoT/2bLVqN9y/Rvvu8hi7RtMG+ReeZA7
pnSOY5nct3dscL5Us+82RydiifF6a4tekx90SJXhuvzYOLHUKmQ1+2MgZsngxZJh
z92F3fE1aX3xRFynU8iakTRVx/KRfpQCISO+wIfxy/Q3ktUprwd/mlrv04qW8+NK
Og7d0OEIJI7XR5T/fdvGTaofKFNZZUhK6fgG34WcDQL4fRIKZ91KR69nogfyU3P8
74/aybh26JQAv7ldHqLWT+os+pWHnbzesUZRsX7IxO5YVvrUZ26LbO8gUIGLr6/Y
TDF1gaClO7LXxwwSLNzywRAuUEQJq2/UPk4JkpS7vSwFJakqpES7dbDCHFV/ktpl
49BWzG4FVZ3alRrWaiUCUb06rPt1PgZRJLcPRBHoS5qYR4gE3G5KgcTxSK19HkAV
WfDRZyLpx5I1WO72KwwoJo2dGthm5VEkGlKBaPXkIoZRz4Te0AF/CldmbmkJ9F9X
MNKLzSuSI0D+K8xMVvKQH/Ya/jHPalKnwJqh11xUKHNf9t6qUXcFZwB18MVIMcyC
qcIZtZhdSM7RTz+oysKMVLaYI8bA4lCJzihi6rkpaJZgSnxG9/z3UC2t+ZDyeuKp
Rtwsc9jozpSdbfDsNnVHhvKRckA0Hyd9sT5NAojAvhkP7LlcIAFqlwFRcl0y5y/1
IxlNKb7LxzFfHmWrXbrpedx0mHgv+36GY4QBmp1ou2w/H/ayjZZWmbEgfV8NiPml
41+o0BEH+EZZvpIIf+M0574Gu6RltWEtalLQQTj8rJgKywh4cmYcC3mKiqkLhkTZ
sErvXXhD0SAo6IB3rnTn3qq1zNvl3eyCEeoBQMQoIepeEzQu6d3EEmEuRSGNAu3g
A7rvq+2Tlt4wqvApf0kIiHDpQuGTmfZa5dn7lP4qX23jU/ZmvAAOh6cLKXwYMC26
K1hOrL3QfJhFGJ2YqL6aLZIZGbAUcTm0ksMkO+jY2aplXn5nSCA2fcjWlA11FjOW
GpotZuBUhomvYt/KfJwAX7OUqBLlFhDzCrpFPZJOcbH7Gz6OGHrcf8WvB+3F1nEX
0B4k3wauCB5zWZyhFoCD7xsocrD/0QrjC3WC02sGPNimUR6YeuSEAgYKudJSJo1v
q5idct30CjE4grB1WphnDZK6Jcaue0DSaw1tBPFKXkkzwz0xvZ0tZvBjvyPCZIWv
O1wYYgc9fmB7JtW7nUsh3o6VvvWqdiVk/hu8Bt0MRQPupJ0YPH7QM1T3ZvUi7N0N
N3W4RJGBy8XzvePPXrWjIg8YjU7VyEvGlmvsBiq63qmzIQLuesoqtKTsNNgfV0e9
LXo3I9Cb6bsTMAYKYU3Qe6882k8lF45oJCr+2uQQbYd1oTyIKOein8DZwtY82j+S
10bdhY9M5yECaljNGKY6rRHPOMQ2M/6814jw+8PxzXhWM9wDCfagg6DQSfnHohql
vktZySqyyDo2iQOEPWRARjl7caE+SXBOfw5obPsDQkZ2d+Atg8Fm9DEFYG5mmT2Q
t2/hWTTisJc6l7UWehwJN5q07pVmXWz9qy73zvKMSyUmPLFerYhJfA9tHkbvGuB1
cvEowOU2Ac4AfiJnbhlEuhUkXKMCCDvjqvweIp7z4iNOi7ezcNDmvPZMkOnGIWr/
d3txNHFii8kWK85qCAWra0cdu/spNEFdgqA3hhB6j1uS64EOh/9IuhuJ9vo8x2NO
meeUVmLeEDq/ww5ZxCJwWARazBbAfaEfHHL/zp6kXYlUy15dKN9BReQkEBe75pTf
vLIxckjJsj5tDDJq2gzl45YsbBN2bPqmVtTtW1tSmPam18oB1vzlAv7yY5xNsOOR
W5WPFYiZODeoHtbu8Q0xumWPqUWfq9zZIWR/qOtLXLsP9TdcR588T/qE2/3XSf0P
5FHhbGG5uvXlGS++oOoV96L2qa42hJAdBvuz/RqeFHjAUgKrqvNPGzWW3DHukXo2
lcWxSPtzdI0sscZcyN6iTVQQDVdoFr+tONLVZ66ToSKCqqwWGmLsmRu2H7YNBy8F
DuoHrm6HsibRcJuFzFp1M/NqNASAAflZvTZiti8A3JA/rfRUBS4eWfCAakg3MnRC
BmcPAxngabUtwGD957my4qSLNasVHZ215foIDG2Id/jmfsmJBU3cGE1XDFs0ZKOF
OfQmir9eNTXGhC6q5eSULyzrFvwxzsjAEzbZjl0Yt8eN3yQbVRmBAalITwVY8NdS
q07ZKYaVRWW2cX8wQqWOzOaIqtpLzHGbZd0RwwxXXRT00SsVMYZs0709gU6k/f6C
MkaxSzblsRUWMrDtRiGw2XmuBsXL+IxiJmyBuIkM71Sa8rwdKrIdiCciLha52l9m
G+jV9H5q7+oMDDo928yHu6gNfJWx283mT8TLJ3uwTV493lJE+4kq5D6KDig/gNU2
D8An8NsSDHhGt52b5mCpSZvJ25j8Q0UgfqqO9kwiksc4oT/H0Sqd8mlOdJVR1Ycm
MeWNlFY4ZEUHVJURYaSTMjims4+thYKuVdz7GcuV69uIIxmp3ZulFHLtMICSkzaz
lIZ9ATP1N146oZnM68GC8AIjnzUonDGSZ/blI7M3xEEW6CpMikHuYKTQE9tQZ7ur
nM8Sb1SkD6HPgcMXvCar3XAyinZSNy3carXx+itKWunY8Sgc19Uu6iDipeZoKCA4
MurlOpgRktPo1pVBVpAZPf6a6qZhn9YoF27v0qivHQUPXCKqQHoEIYur3vqm/lAR
6dTRqH48IgRP8WBEzzhXI7y+2F3ZNfnJNIsznie6Pojfl1iMAnDKr0ZXNFz4vKOZ
zUex5v12Kq8LjqfIfXp9XiyIG2mdDSdWv/7Ue+KyBSAE/NlCnR4u2fpmbRy/R8W4
z2wc4LyFhkotW8caaJ7tQFLGNbE/A5s47fBSMow0EDdD+jUM1yYYUvxa6qciW4Bi
4Vytnn+1/7xNRrJrfp6rDb37fJZCi2o+HQfnIK8AVrwLvD6ViF1/OBCIsbc/udrE
sZWyiE+f3cv7CtVXXnAi/CO2FKSfUdoM6YZ330Yvx6GmSPYIlOZEZ82g1XPUEqSX
/lb6+FPQwyrfjXmZlo8XS2Qg26CEM2c0neFwLR1SmuEqscRr/vZBbjd9gry2pJAf
7i6yTduPQ+Ajg/SCoT7UbEi5XOjfKh/u6huovBx4itg1d/ras6TEvL28VyVG4tXH
VJRIVGM1mjNCBb4aN/iMtTQIAEA60c77iTSAeiArxt+Fc/WvWHvrc+/cecSY9M8H
yOR/C4ziayvyLwgCfoCOYzOrF7P5U+KgpR1UGiO9//OWbqgK/ES6BV0csf0JQJaJ
DBMIQB3eJBRDGIBGwqBxASjQ+doaYQ6CXtviAPwBmdgtOPsZL1WFndeHlPf1abfC
dZTFKY9nfb52AFFoP5m/XZtjsbyVBeL+E3LTEC780kBB6eXfKylqLlOwxwiUgXi2
hHjkF9qbNXlEmiOg5Yt46nHKSZ7v0JP+9mmTkFm839VEZSLPsFGuO4SPVi0Lf40+
gXb9XTmRGVrZ1aUon1AbyfNmTwmr9z1vSV43oRkZZ7uNXgFATcIax22lVEymS0sY
xhIaV398a1kiM/IJ2qif/XeX5AU/xmv/YL+Q4qLxSbi2gTSWyoMrxji2FbAzGlDu
TChHT6qwsmOs41CbTVxxz3V9kItDqWThKYe9mnrsegYJDlrrqzLmDgRTyIhZRSmK
0zGUoGP5FN4PjL5a0YjJx4mU/RIuIU0Z9GQMm9WzAOkE9bRlkKCnIQv6PjbYm47r
BOSNdH3ceGtW1k+xwnqc3z3AxMf5xPNZX9hkl+gae1v13pGWHM6nZ51JQllA1Uv7
Lb4MD3g+eBZUzsH1hVFLmdXmE9ChCy4m9ACtGnn4Y9y0tQds8zgqsmNxF3M8RGHN
sP9YqMQatNtsaXVvNH+dSbzYfErqjMB9I2iGRj0cdxs/pIj7sFApm4kRNQ61KawK
VnnCQTDYZMxPm5fn4xRlVxT68DLOhfJxE3ny18Ck0ihFEwGBRAonWfR9IfiwTrqy
83uoH1EKG5CCLqeqW4odKaQlZUhLp7XlMkJylCAqzYCx2RgfZ/zvdjWkmTeH+pfX
X1jVt6lWmF8y7QS0eIxrFxExzpoiAb0UjAkE4XSXlGkW8ej8kXImMPcV7ZtH0ZAt
cuAyY/wFfWkd6acswYHtOCA/zRZHar+KpwoTNbrZidX+d+iKKEkUvc7+OZLs0Cbl
D41Rbx81OCggMWnabih9+jNZoPEIqt6ZWiMHU3EPrfbY5cGSW3Klz39gYLbQG8aL
yLE+1ylR1sHXHPTdfcLZLlTjTibPURgj+T2wH3FrcIMfxKwWeBX3sqZIbHV4UHME
wpv+iIYm7S1XEz15DycuuhbHFVmnPcsFYfgZkU4eeLuKUWs8jdCQnwZtYwLjktTz
0CjO/OCDkQq0oFrfzcljYDydyifcZkRJ52uCVeZdZ9G9kmbQk7djOBqr5CDL03hJ
N1jTzA0wtzoqNPXR7lj/eRLeNqPSMhP6uGlt66//a3a/eQ8LAgiIhCeAHUsXCt4Z
5qbp3ofh8wB3SYvX+79Ub3/fnDBPJmZD3GJe9cOjwpig9QQpj7SNSQQKsF+0IdLr
F0sW+r8XWONa+9UvcZZj7lXlJzJJIn9E1jeOc6GE0vImpjbMRanxQCfbUmZhY5tY
IlECYVGUU7PsububVLyoSmBPwwzzppVPJJQ/gWirpsvtxcxjKF0SSSOoQX3kHxxR
4ZfOmPeQo9ZK9GmZw3QVF2izbx+AKSzQoZ1kC+dgkA73VSfv41kFYwn6yK0knqWM
WLFvzbIjrgYnEejbYF3cYli+A4dXjrBKKYqG/gXRmlYiFWawWk39eCQNh+KJ+LOQ
Z/+le15PMFouiJ5Nu6Rkftn9yf31tiAx+gHk4VKOMU8ONrThNVIWiWVt/4VNT8A2
JcKyAUI39VHaWN1by/nDiw3I0HaxzoXWa1g9uO4g1V/hMhrTdrsHwUhgvkI+PKvP
yrEKQemXj/QLHuoaScOAHlY1LMEdpJ1B0y8PkBb0QcMqdGAkvvtowR5Z4ahke04e
F9FnUxvfUtXZ7Ez7uxzTq+hetwtYRXbFQPkcfVyu3Y+DO6yo1HvJjNLXH9pRbeAr
MP009O8OKa1P3aO8HstybFL283GydMNzjgD1Ge8oh38hD0DQY3S5AWLn61GyAMUS
t8x2mqbzvikf/jNBTLFLVwGt5b9y8srAbfLJ0hi2C6hDbJpV+UcxqznzsL4wYC8I
ASvBy4PDo4zjtP8D30P2US63D45zWtp5Rz0flpJik6wlA4QL3Hu99QaiyHBtNpvT
HHvlYvLrD1KEfhX3X2FWRFBD85s3zJ/Qf1mEAiL8ybK3/wLj7/E09SRvUCgqVJl+
e/qRwLH8SgL1AOYUZkotpEGH4mVzeFOTwryN4XqNZ17YkHUc00388Mm+11kAblJe
Bf8cZcHTl4rx8XxilzTvKTDkk9Wi++1Hc/3djTic877JDcWO/AAsPJzl8rvKmYDq
MgbAMBcwzawBhhTOBbCgMBAx9jfRAyuK97pnz6CJvzyOwNOh7PikRhnCHQstKgKn
Wrd9lyZQaqCVbjiDN1oPI7iwZx1DiWHkoMbKTxQXW5xq/xo85CZdflYW0UGrGgbZ
+KLHLsAUrzXvVYwfggTagZrdQ8+dp43Q1bYV3wON0/AuH6CudrCQF0xx4AZWhg5I
8p2vP2sPcJ908iEh2bO+KpgWnltTsiexsug4QNkC5zsznFRwSxjLDybSLlDJcIGb
ggGVEL8ZLahB54whWK6V5XIw4BKt65w4oFGDcQt8gBBiSYoHGtZRi+CaEoLTKXhJ
eNy9e+MalTlWTRRYGeBlg0UQeNOgnFBfUK3DHROy4zQ5F6GuvmiSStD1Sd6eaywq
97ndf856x/XhxaSkNBHGX+AW0OAM3lIi8jBv8dv+zBEcdfYe3iFbdTo2JJioImAx
ZTESoDZDq1MIP2q3bukfPhjEDBH8pKunhyPm+VSR24evL0oKNcyqYTiu4fd3rco0
A9JM1e18JZ15kIZCeRY65b+tNYjoQ9dDcrhJ5NxgN6ANp2ix8KqFHfBATWF4wWfa
R3vJ93VT+Rht6DtR1oVz1cEiU688nBRG1xYVfBoK+Fm1G/zhlD6wxLdgAauxVRa3
U4g0X1/ByeFMmprzKwGGf1H8SW/H2aOHB0tbAheIzn0j9Ux7fQ9G87qL86qtvnS8
SdAo+lTIrwckl+icpsNyNO2k6XdYYYVeuebwfMlQYCT4zqdDavZeeuTkXpjSuJ6V
F1nMiHvC31VpN07r6Mnkixg5RIlgTl3Iqbh2YFk3geqtkVu5W27CWwd+KGtQbDIb
wYmYb6AuHQJibGNKcdKQrUDoe0tdWctb3TQMyDyAJobvCkOyaxea7aNpugC+wZeC
nSx6XnWpSVWjTj4HNIu6OWRtjVs5U85VUzqs0VigEn9IIGyVtfrvGqx6iGNuZiAZ
9wExpAMS/4u1dBdEqixY4FfuxzxRCMolEJqX6HWrV78oElcZ/udZ8BkYOdvG7icS
QUcIm7YuuXUN9oR+EO2lzrxE8fjRKJNsMnh8bU9d2d9WpLL5eLcue52n7TAfRrps
ATRFmtN/xs8PidOQyiY6daV66XR3jcaf2J5vp6gjNfao2qFG2+sdR3Wy0DxG9yM7
kgGFvJg9XRsJVuaPzkbTTpHy9e0RfdV3it9AoHxl8gAP06RZXkE9nmBt1nbLpZjB
Sm6rxrHMzVjy2CAk/gM1+pGXLI4SIO0Ac16IPYwEYBN/XY/2B3gvh2zshuXz2clQ
JzZt99r/RpFD8tO6HH0mukG56wBCFkP/rRSlXE5uU2p0zFZoTbG5KgPCYX/IeGeG
Zli1LLhx23Ds/1BXtjEud7xK/0Wa57M666zKK162aL6A78D6D3q7Yr/UzuOxy7It
FpcAj6Ypwyo+0IJ6f2hZGVEB7X1od0PUdbjlgI2/DzUse600raWqIQEKny+A4c91
6axLweAvN7WQTgo/Kz8kcssxPWjUMW/DotYwobT/A56pcrwniRBlfZEGIevpANbV
qQN0ZvU6dpwr68v65vYqi7tVsucSSvEL4Owsy3/djBc9xlB7OQjnz1T3OJka74tD
Ib/mAdDaKaN47axq6CAupPSoIYfgzAhd/Ifxx+iNmDIqrxllDNx+a9BZTkexJCPq
NQglCNGIi/Fut9+CrLRGS4JKNGyWBctCxMDbrapBFWbOrNjFwGZfo86dPRJE/SzQ
VbyZvqyWiG9jpDiHzn3SZQEWO7hBjOuc3JqfvQjNnCGzrHDKMh/vda8QONzhk5gO
lqKjy7BvfsEGDuLvo9M0VBxHCUNpMRXX4lnHJafLWpVhp+adb6YioZzj/+rCMwZp
+S8+FwgciM2IjRr4+ZNHElxrWm8PHllB3VdDOKQqxMvVJCCOM0vTxWFGF1P33h4U
44YbnaKh7IwzRsxMsdiAjLl+APhT00q+ScIoZWeq2bIGoiXPKD2XNwRvKhW5ixaf
MeM3JJ1CCnYLcoi7icigblbi6JwLlnV+6gOWcUupYKDrvosoVe4N7gWtd7NkKmin
PPurTCYh+RDCk30spBCFa4ZeXN3RLreouTLsgXwzagTOvofoGPj2R+vux9QlBJ2M
ykSqM/3mlsSZsK4kmDHj4hxP4ymgi6d72D4YpwombHZ2JRzmmQOuaw+uT5uQUUQu
3SrxuZTJV8fex/7IBkiV7mFD7Tr14KZO4lTd4Eme69acfhGqHJK1INfgTvWaO7Fc
cpcMcEg5JBYn4pmlAUmI3LUcW+QDcgs9o9PlCQ3AKO8L3fV3/oa1mWX4vH44VP8U
DevfX2K9XSR4Izh4j6TZbWuV1OEQHMpBgLvRkgejJuJrIecabu8tMIvF4k6raBCj
m1/Y6FDXX2V1ZzyZ1Hd8x1wMUdVL33f8uPIUB6aTauvTPg+tSGcgA876+YPLDmOl
dqJwIGqxfdjpyhrY6nLKH0dPqk7D/jeVyMXsgd+EjU7BL/G5P6Sr6UgM2vj+gB1+
RCBFuNY8gTPvQr6bsCUKJtG+VQOsZLojKh9poL+YnNakhvwq5sp+0zZGIaKq3BI2
U+Pt5gtl1w9sfCK0bJGFrMW4U9ypZ4Ago8LUGN+79EXi90s52m5XpS9fou+wW8nf
LW7imdWTcVo2JrGZusAnHMQera+wu8NF3rbOsVpf5sx75RPauzPH/2M6V07yxIZa
9NgZDUj+cTAhEmn/IFdsakDPPpAewDL15hkzmWlsxjcmnAnt61fg37Oy2kx1q1kC
nxpaJAmVBOu/xsEjHRxNanW5MtUjgD/k46G2+yWFoOh+O29u0FWhA8wMa+remlyN
ozvDk3Uz4Je4FHvkTAWP5tdbF8cL181UuILxHzl8mZ/v5kRrspvKQIjsDfLtdHdp
3/40x5PI5VDjNOmpDFcL93GSwCegtRMyjd+MklK1JtXgWUUYD5NmdvsdCJX/LDOB
SmE7fJvJplsNVWsNaPlDNFB+YUAbyP4a3zAl2plRdKZGKtLNtrCQzcMqLMyicj0s
kau2+ej4B6PXPLh/HXT74pv+aG76T8Be1YiGgD4v0Jt8MjYE5cywuFoIsSWiOxbw
0EoC0kpZxCfXWugtCrzK77wkZxUpziVmCSAXcXb5chSz+bum9jB2MQi/jRJ9MV6Z
ORkAWOXSUNbjA8abQ3D3S9yLHw6vfD5VUsU7kyt1WOtDTEK/2do7UgG319lN0jE0
A98Y4SeiZeePk2n25Q3Z1RBe3XqJSIQ4bO8E+D+w+pAREMn+jwSHlPg+X5WC9Pq7
U99wYVkbFgMeo81VHnbf1FcOQWQFSlEkP6/rOiRUNtNOTZ2uXBKv0n0ODYpW8oRe
yTrqOD8xcZHUupMoFhgsE4G/tjQbVrolGKp4c4Meda+t3VTf3XFJS3/gpYU/f4cW
aCv6p6WoG7nwOLT+4O9q5zWpEDJg9JvigG9/s5IUSnFgdSH+4aJsfQHA4dYFQzKD
QgqF5N2G8WRAs3Kjd/9fIkaD5JihiWOVRFVAKfo0bC+WBNZG9lnzKdSZWE67jL+L
RMfpBRaKcJlD9WD07xLQvj5KVsy9pQbdxcfRQJ2MfWv+H4TscoHuf/wE91LZzOh6
nhrkbk0Mo1SrP4DJl9vR4Cm6Jf0PC8aMQMW0/6Jny9KP61L6xFRO//v1TpTBX+2F
UzpoZsNu8ADOsx3Ky/+csnGpBOO11J1VLXvjDGLbas+wrk2GtvNK3yIEdrrOiHDU
xSFgHg6pUaH5rV7uCrikjaZ0mPUYxX/f5BJhUm98yWv+qeEPvg0aECXqsUX9YerO
yMhKEpYk+OXiy9Wjn8v7H4Nww2iL0zeif0xg8cRM3AzDQILj/DAgq8d6q/bNe68c
1La94KikmmjS+bhUazni8ucE5Z2WO8fGr65X6BzryQ01fwK69DcbbCRUWIPEVrPn
2/jPmbQnKS9aH9ieiY2EIo5cpnjmrgKYbjnYo0zsk+9BI8t/DN3+ikFvedFcRcKQ
zETi3TdvRIERHFXBraca/Wo/u+8UwNzmEApyzfEbePkxp7F9niZVAQ+pnl+vPWPB
7+0H8Rx4Q4PJ/e44IWGGmFSqeK7Qk75ONEy3GCCPaKOoe+MqifwNUiKCEXKAqUP+
pzVUKk6ITAy+3fjkM/7TN+bXDzsZm10liMAfJk+UEhdQ9Jl83Sa7GD/Lag//olmr
PQka1vxhG+rdzndru+T1Z4xSwcP12HKxZmRfoFqDH667lQ8vwzv/5/mxXr8RussF
lu6wWKyEElKU2y8LUUEJhq6m9G4fU2r+jFVcupFN/wEj8O/v5shxT8im2h9n5dsB
CDphL5oFvhiGOvwZ9hOSqzxY3CnDGKzEW3u7ZmtMnUlsgaJb39rCVopVziMSYBPk
4CVbXoRtsgmJuLXTXW9R+1LDxgHGDg4kuO3aD57UcpChxtkgB3EocoDfAemEXTXM
nLvNohOFi2PNMRGCRsvg8qykeMysdA8vLLkk5TtKd9jREiScurgYhMLIN107B+UM
3EWTN0eEEs/gNdz1etMvFbn9QN5t3MkTCYhgR9bxiZER4UGzBm2YtazaFcDfWToP
JyRNycKmLApVfhcQynOeacjii2xaTu9RrsbBcXYWZmnL8sTdo87NK6h4XvkSvObs
iugLimG3RdJmi9AzQABc5yV1WYPno5lQyNEKjD6j8+jSp/8P7AjQ7aWQnAAY7fGy
0I8zBa00InCr7OuCin0vHERQfkt9DaKYjRh6NhsS1lueF29akALhUclsB8NfTFsP
7Pi1uWO2vcd9COf3H5cC9jV3wnleu6wAYK4wRzcEoEraZTj4dG8sd6zbJCyBZur5
qpTgap7hc1Z8kMjjGozx7SXcfnjykNZYIeqiBFcIVJAVO+eF72YY4PtuHMXvVF76
/sUcf1FlimZxxvRIM6CBTB0m6PcjG56wxvh2D/cLplQ4GYks65mT77n6E3LuaBvI
IGnnEHucHTCLCZt3mpOLdc2JuKkEl9qn0KJahIVOMnxqjkFiaioalODjsVaqETRM
yZDUjjln/Qm4+P22rsNeaY3RtpOxcEdBnm1DAi83CV0f0luDCdq5/wdnPgkZV7T5
VP9QNGPt2iGl3YQxmiN9H27jmUEPwbpJAnY8q2ruLzncGXPDP/lzmSofYCxdJUKe
+VIZYrxHU9xn8sTmPAhdkokq0u84sDQXb9sGQdsyxdSHY0Vrv/11+91LyizP+A7K
8bpB9PUks0o6pDMXrpeSsLY1GjfHvqZIMq/ISnrsIGrvCXF5ouKtt7HVVXjtdbkE
0OoFCnejteoy1s23yP3GP6Q6glZx+yXzu2Nu5ybsuua75TD1wq1pHGfk9Bm2BKh3
Sl9gz8I9vqgGCTXvtqU9quZ520lauxg8oWPEOjrnRuNRW3shjKqiVp9Smfod4e5N
cmRZFUn0WNOtqGQ+oJI4upWI4+VeFL95l7ZrHdqu4GRHpkWQejgKKrYTqRlbVX83
wWPbvgDnN90yWCtxHUoVDh2OTkokDkJCW3UOyyAIzxGLXF3swJBLeZXf30ZcZD8Z
D/NE2Nre47yr5eF2mVR+l0EG4VufZN7CuSTcQJ9VX43RpeWOwWTF5OPrbnqFkbJq
Lfb2B4ZJwbFUUwOb1NXC3x9FKXnLG54vNzgZvuGUS3cHyEj8goMAdWhdfhPH0UdE
ULDj1OZ+SAZtd2LC5AWzhHK2y0JQhXhXbgwo5LeBy2z3cQ4YoXxYRptD2r9ufe9+
etL86y+amoWRHopAL+xG03NDCdqVXgZPXxXxgK5n5bxUCmyT/9J9gMJUgUoxYLE+
UNlEv5T5TXe/8x7vy10Q8IyEVEvJZG6kUPU35Fd+SqJiZFVcK4UApIpWtEHcyYNb
2PNhoOeyJiYWRCqSbO4kBT7ZmNjXrLwx2g5HuADGSWcxUvG9NYC/nLxP5c9ojTRl
IDtEw9k6vubkO4YAD3NR4vTGf9f5RzGJydbI5COAqenEaDTpLRaZGH+XUaCrWYGt
zwcRPHq2TBvDSk0OP8LtGet12omzCh/9liszzEvxlGXDAFDS3g38bb9+cxWiz407
CvztlGzMZLNtAMPCzfn7Aza6s6rF2j7G+pbSeoAzDhuZ98o8CsMS9z+g7/cnBKZq
KUxRNyKfTbNMfyinPGH1jcAmtfFPsPXh95Jl86ZTgWmh/ZPf2/Ppm5HjKPxXGVWl
H4IfI1Bhy2hhDzHvcjv+6efcjVmeHcV7FhnUudrr/nqpJHaqEJ8jsqsxHZ4VP/Mt
scIRVNqoqzbTwHaaEQG+ywZsKb6gmILuhu2ERJKZoShsRecPUjEEch3ziCOE7a/u
OtYaeSzhLqiHyXudMl5I8rQ+rL4J0gnlv9Hj4P5ZcANNpEPUpTZFp7bUpo0I6cU3
+YrMyN+0JnD8eWGJmLZAnDxA4Ivi6PT9A11tqHOlUweW4ZSFcdtFfj468NmKvKOx
2XVCF8CKpgSakqJwZbj++JO5PJpxH0GJZc+k2CRjOCyp9TzPoRpRcV/miKyYOqXq
LOeLFWNUxGRYngU20YCCSRgVy5a+UNi3Orf+x1U+lfzie+KhQ9rR5hPuPsjFyHQC
HIUBqymCKe8YBRdSnEBmhSgBmsuhz09UO2keMVLWzlU1ASdHDvQT8pyvRKkFgJmQ
TtSyn7uOycc+PBwXDTDCc3kpwcp6tq5b5P4hVJbZkDWcZuxNs+ONgN970+4p2r/u
WDud8TJhQvjhHULJQvgPncHxgxtYlC0lNDkBcrS2Zhf5dHVvXF+A6qRQFYxE968M
MjOLATODPvwTaf8pJ6TzZTUPO2jJ7UgFgEAZ9+CvSNzc7tUur+Ex7v9uK8ou4+VI
qB7gnVNaTXng/1rmyuJgqt9LSDdKusZmWSF+muCT5V+F8zlruV3U9vU3w1SxYlmL
TrVWxaO+44+WEKMxXv0u4SSzzu8LzU+OfB3usJUnzDKvo6oOJVRK3v0AtBIF+YOr
8nPHJ80TswTXjdH2b7iVhqnI69aYMXC6ZiI5kN2scvrlZ02yPufGWGFbNNDj17Rl
/k7qFDakVkZ8GCN/Wk2P9RPsiwKnCNe9WdqO8zq7bfrrjfXM082b7lQQZb3MZcIY
XIkICEbXjeqjpXvYI31f7DWWcuAWokeFh35Y2KpQcxgGxC6TZgEKE1r9xGMUY2NR
CphXRK06b9q88Ppp0drtWCPGFxbgMXVpskPQPWYD8c+cmHjLPya9hWSaw6MHC7sM
+Jx23CN+FJqoOGKP3kkCC5mqrDue/axHshUk61E2lKHSjHA29paTzUPb3BPkoaJB
WqNLZlx5+V/+uuonorung1x16itI8K/nCblQC8fMRpn0wa9hyRq23jNn1he22cV6
XAxjSXVtpW+UqIonx+so7pI/mLdishDd+7JlFVRh8zGISX3/pO4X1oNjNYR3CZj/
xWSilnYQmmzCvMcl6EcItTTMDcs/thEeKwpg3D6bJsqoEVPYjGcZJ3rnfNyrjIW8
6ApDl9QnLfb7nYDRSdKNdXxLV0BXTd0iu51crOfUX1mnrU2ck9QfCG4L0rlbxRo5
1sACvnty29vetaN9q8Ff2RFJRS99hm1nCCrOiDozOzdbECVJwpwXQU4QqK4zP8Yu
o+BuPhTp58e6lucspxchMEDE79QHKDm9tX1mMg8utOTJ/Y6Oxf9mvPrdOqdl1+hz
5WdBKT9KTBca6F1RE8bNpgh84oDPw4RmlKW+I9TutOX86GivOg39HqofqNUCf1pY
7XdkD2BEbjvcGiNgOFVp99AlYFlyCH6D59ueVLupA/zH4BjwevYYZ7C4M1qTtjNJ
usyTqixJTyLv46phUPH0pB/W1hUNTnA+f5RylzHLxTRccUadVtFtMdiwm/5LxtAs
awCiCW3Zfm/mVtuq0msFeNDQlYzVB5JKeYGRehhbWJ0X+e6BJl+6C5NtLyYlhMn+
dXvkeN6oT/HaUE2hdOO+SbAEU0gvd92TDkUnqi6RKPTdIHFQvqXN6Ved6mhCDdo3
BnODOZjp7eYZw64lyA9xzk3myABObjc7gGfYDCdsIJkWJyS993Mi7+WJTRpMQUmN
NLSYrtZzOdK0fsCTZOIt2yipMpW5ZwcVkzSKXl9EFB3TJvuwv38yh4wn1CAr1vXJ
cIZd0rrVwrmjPzSCOmA/vzrw3O6Cg+g2jAIorERLV+a/b3XpuVdMfQZZTy5P76MC
XN9aonl8GpuUWdaJbSDeIJY5aw5RCac51bjtmfG+XG8kZkX77qvwN1+U7psVX+qs
e0Q7XGNp47Ku8e6f2wqM6SXx/iNLXzveM0ZFjpGV/zouCDWTbrRTv8PVn7sApQc5
n2sPpAi178WSzAEMOMWWN2YcOyFuwCO7d9B20nM0M0JPDTpIChCX5ZqpvgREK/1O
m66MinlGX7WgaCtOi2GNCLY9F7KMMJKJMB53WXEx2iUAZgHZTc2JtjgGNjZsIlBl
bGKASH+kfMksLYDLn1Yu8b3G1AAWvMbtpyqNbve4cr0w/uKoBoceQ+Fpee2Dv0ue
LjfCsgs+PHNj6KQWT1UNY3Td11Ry9iCnoZoksq2Ae6u3sU3oCM9JIS8xuEVlOdvH
gzoM/Bwes5frcFYWDtUATao6Hb9nB3SqPZEgiJ4v1MAtYvdndAdhpsFUlWtIkLng
H2nxiUwViwufedqbBD14lZSVtMPuhLBf3n5AZ7GuWzy+Wm3uZTVYBMibTekp+xEh
+k4Ys8jtXbuicrz6mOonjI4/30bFjDtWrTGYuJOmLnqvp6T/2yCFOqX53r+Mn8cv
cu6+gabbZ4fxwpmLt/cKKXKs36Cks/YqrC7SjLkGlVx5rTIUeChoas6c2fcVclOL
67G39wKag3OegjDNVy/UFCMopeUIvl/cs6nrw1oBj0gtoqWsGYNBWuKJCpB3pC6+
ekaGATbXHAJL1ZdrC91Rl0tcHZg6xWp7ErH/8Ye0+FLMrh+DJhGk40/E2PoMUAzF
0Qi5jUeaODB4nGsYhBHpIP7oBrPhWdSO1Ls0LcLw68Q5NlFdN4fCwX4AULEP4Lsp
YVG2XPtjAxCzSwN+EnOp+/cK/xKDIr7k6Sm0ZbHiLZYxwq5uj3BVVk+vGdgfG0Fk
xmU53mx7TmslJwpt46BXs2o5+2NOmtiq6IdGdw0XErWUw2qkLqkLUkDRgXJT3n4l
kB5+seQlnRACEEJG6HjcwpnY+Z107hioRbuebFe5i44VJ53J70NrAUaMm4MFL+C/
UUNhLpW9fkrN3Sc53RtRqgM/UOT9w5c8OcLsNWK9cUimIoBo3uKmj3WeXvvbfeMf
YP6LeASWNp6i6CHMnMNRAOfCdouBIjmN99GPaueQy55hPLcosHcY1HThGnewvPRS
Ex7sI9sAdB6VOY6w3fcuVq2CknhRaMUeNhe2qu0ZRHR9kuUWP/sgAajdv0inIM4i
yO/WKgrB8YvABL+XQp2QcIGKuPXw+f4UGyLXxwnzlOyPcYLqWZT2YHnj8DnyVWg3
Mod2yjVUo6uahVxLapSntkWRUKMN7qf9EgdwGE7JQ167hS8+qgNFDAXFE55dQEkf
bDAVj4ouUjU9ibgY/BJbzrPDYVzSKDPb/EkG5A13H/9yfpE4gqoLIHycbgRVcZ1N
VgexpKjlcQTocDKsmyh/8pfxhVhoXS9Qp8EF5hylv5CzQgOPrOIB2kDPH2sa4Ths
lHyUVJK7R0Q2aZz4So/tUhQicHN5UjfiF+SN59VWc9hIWIyeWrcbA6bVBE32mAyY
NjFEbke0M1KlgmBtbH+MUu95LNC316qcOUuKwtpfgXmpRFeqfGPtGCFRJxcrlPN1
/3n2BfFHOxExpMIiB/t6Sdg3DbJTUHIw7rMmQZIHCe8TSIj3LMehjvwMqXHC6HYR
xAIbYPkbWnFnKzsHt8UfpeRghYcQPzkdnnovYndjxtRsP9pfnC5G1sUXeWWot5wY
2u4nNaBNuEnjcSYlR6xkbci50P7GpTBzx8khnefvpA8V0ePT8Wu9l3PAsA7HmF5W
plAzq3AqRQKpD7dwQo1eHLWojAVVMBdG9ru8oFY5PU+01N2vkRYNuJq+VdDBHepc
DfyZyKuCucKPscespK1M7nhak+eE75bfNlhMMBdQf1ucCYDGb2aZjm5mWIAFfMon
qdu49rhJ8V4ULYYGfcjzbdgLIzG0SiTG4wpGsg/zs2FxGI73Tqo5jzb7LxT84odG
6IQwff09YhY6H6QXDcUIqDJEcAA1xj0UXZt7FdIzevhG2iKQEpEsynAiqN+0sCEi
hNhV6KjvroRHYvaJG1KQ96GI4CL1E288/JTmfPPRlGH0JpYrKvHATTElmle6e1B4
tYp5ctjtgGsP/v6iGNlM4zGpP+d0m+DdGuX153cJyCVUKtQywwSe5mZ9xVS/XLYB
tcZOSF5e2XtWR0tBd9/grSXgA/NFMciKI0FvtpCfQ3+VHxgXiO5fvCamwLhy3wCH
Z9ag9lwnoEQtLCL6DYnJx/ZNxYt4R85lEPC3pO9rdk7XRRR/Df66X2shqkrPZ7XX
XfaHOfOwnfbyS4sjBgS+SovVRyRnMFc0jS7EIWFHKi6t5r3AESdT3mh8DDU848L/
QvHQcVer8GYb1+nvD5WZD3oKRvW8B1SV8pnb+rPBzAJtsNFvqK1y/HR6aRq6fTdc
cAtmCPEcRF6mD3O0ZhPmqSZUyfXnXSXfCmS8kysc8Sa2wg6+NElJxM6mt5QEV0Gx
GCtwlByEMXhwtVT7c19aGPMq8CsjsF2klAq1UUg4ptYA3/vvWcsh0I86XVRYbY74
o2CwEva3fFGNihAZ4MP7EIDsObn2oOLmgkVGXY4gQKQjIpIbn/jjcG2ZptAOgOth
Uc/I7me2jHnC4gxbAXybe+tJ2XJREu2AWPmHdSbXwC3rge0Yl9X9bOMDmUBc08Sk
jyRqJuVr38q6Y1hXZJfPV7FLpHEHnfXgGgSYPyawxN1/bpj7FUn0KYabI2d/I50r
n+HufMyek/knyT021e+xL5L8dY1iRQg6I6z4jCejdrYGzql8ZCVRxizxlBZ7437+
rcAo1M7bIUQM07b7owRLUBJCYjuAKVXhU0wzdVT+I67qQ964hKWR40DSsZn5AK+b
zD1gyn9BtysJvMAcxEX/tA4MCg0xrMaA2JAcd2zZU++p8Vty4cy2YtCR/9Fhlgyu
aVMbZg0fsBDRd4KY45K0W4iYq2rqb/Y4DaWZRWVOfVBBqUI0iY41pZs4Qyfru268
APlD5c3XUI7BnXatqFKXpDr2enUxZPn+BxYMQs5qgAeqzNpLN/AN8v2x3tqx+YJU
T4+h7nNet9deAKq/b+EpM1elWHNy71484FjlGzLs+Jz5W7wqFP1tgtd/4ZZli+qB
Li7nqTuv3lIU6pdYca8LKgmPrjU2wrupXJDKQmG9ud9RICZmKspdGq71wlgwAGl5
OSwMMy9QB6enG4yaE8yQ8g9jaJw/vn2yPFDEn6mfgXokMnrUtORYmH7yPUy9de93
qeDlxuZG0rXD6plN1+NeWOX2OcFIFkHXgBFTJ952/rDTEAG3NfD1KK40iU3qvlTn
JmqA6ot3yn9tvfUkaS67l+ea8aAcHQDqPCJAK606dhBI2NeIFAy5jQVLq736nYo2
A5qc7YLz4W0D4ANNhKqsDh1g+2PkEDNrA9YMVnIZEkjPwUnM2+sxp/N5RVCE65qo
Is0/9zULztoU5yCmHx8NF4GfKcqZc6rA3KsHNa2i7+8fyZgqXSY77IDEm0OBNPwv
DYRNPXWzCf/i/4SVh+QgRsKORayo6PvaQ8dgZliIDYreEFyVXinngMacAxgSE2yO
ot0rCwVSj8dhB/5joc+vuohf60amOYuAUA7k4cUA5eQks3oNhK+zsM53KUF8Yvku
fcR2v7cxzon4xGVKs0bi9ma/N2SByQIer5t2Yg/85TKOXz6KE5dRqlhP3aXRp+6b
/pql84iW+xCk9VB/maRV3bb00Nft62QKK8j/VEgDxSSzpej33LGHK2l6LxTniILI
qz6wChAd97oW3wQ27wbAJlvpIs0rsnaR1Rvx1FOLTqH1Tt0wwHVPxutv9EGWTedR
mjaEY0l941lpaRkPzlCCETwVOwfIuIcqu1itR2UeiPyZzKTCSLaXzMJ6LSj4HqMg
E4bjYtai7nRrH2bD2qbL7ePgfNg2laXUG8PhC/vK5lS+pRdt/Sxp/kDK7mTdIBJk
CLhEiJBcTReZUl6COM9so2q7BqcZXI7Db7p767ZOChCmatEczYJ27ZLOMR0w7sJR
n5ewISdy8G+yxVXQIPUoQZDr93I1bmAlimnvDSidOfQqXlAMCZD7f41/W+BEiVjj
Fhe0Tp9bhiC8RuKYy49Tl96zTjJkW54zEDgmyiDgkbm3PgOiTpozEuWqEvZKM/MS
swBbyn5FGTGvdZ+ReqWt3Bo9gQJkND3nBpzJ9IDMa4j2YBdZPljcbULb7vqu0XpY
2P1X87AFEymCPyaAFUxeosdm6w+/5Rs0vYqPc8BIgdzh2BwrRQk3KsINnZLEDmzk
IccWh9sSocDaIRggZw9vqkKucqt41W5CjpiMbXBh6lkVLl519byR+OIegz0oAcml
dgI7xV53zhbmfOL7lwqw8ig8RBRWBJEAKYc+i97C/YL2XsDm68p/1buNqQPxxBLQ
l9Ya5dinYwRwSnJ/OHdztvuZtF6PUylvKyIWaZ9fqKPtXy+cjGXsUKAeqmNBC94e
9bS+SKJV2zNwsj1QJVvl5JYzIJWOognq3us0U2pO9YtbNfxSmn4rpURgcoORrOBf
p8o7XREENumI5c5JRR9L2LoOkQgZ7oRz82dNYXv53JpY4ZBB7dfhX+4LjS7c7CDt
XaVv5socWrgpfJaeBY9qHwpW29N/QLUvkQeAqdDmQF3rUKSXogkGCjI/ZU/ON/zY
CmMn0bw7sIj5yBgn7Qu9sxUCdzZGjyMfWGYRMgV1poDtLNNIs3sgP+4ggO858QsP
lTyM3U5shJV0Lp1VuazSHa+Iv7nc+NovCLfKEoJpyJ4rb3GJsQj+K+SGkvYyoY8I
T5BmUOW/eoIgelrz1Y7i6MZLj6gAaVAqcF904sVmT3leqzlA3UbPwLrzM1n5+pf9
eZ5vDRkbxsVOf/xsTDmZuqpEGdgho8zrqgFXgL8YeVRD6t8X+u/5Xy5cErWSCsew
Ti9P7r+MlJu8F1p/TmRzOPK+9x3n+kgOCMk2rnahU4JVeGoQ6OfaxTAxqkGpTFow
faw3sjBpEuU3ckT9Ed1cNXga5GeZ7UaOgXrGiq6HwxE8/caAPw9I27yZsz7xOOH7
mzmDZZbxoQ7S2uunizQ0TEeYEgKbENetGrl6EtNEPvyYT0Y+nlDpZGie6jxof5VS
bvxFoJf4VZHcfBK8kdn7t752a/FIZ7KhN1s4q0vBxuYgUFpqdy61OufjAOdoRxPe
aj5slZcLsciQr2ZeFq58a0ROWDcb81FpOnXouJRCmZMQD0ZdvqI60oSn6vg5bNXp
QChyR4OULyh4dBeTPr9myKvFJH7p3m59dlMEfIoxKVQAr9sAVHLK7HcaGOcwQEYs
8Nnw8RnGLrpz0Ho7KZ+GP3nHs3SXFx42VD/nq+NjI1bEG/h36r5aotEqK+OyXMb3
pI3us8e4BnVk/zfxv2qLoO6uvJgm7VPOSSNDKXC3NSvPmAeURkPThLP4ptMd4ydE
IgMjfFXXXroC5zDHPExFfPl/PtPZW/AfkQePsxbMRpJlDXpc3hEz7mveTIIJPZam
Lj0gJ3bNMLKQWY1U0ztICzcpU1l0v4vrCwis5wwC0QBgJcxI1MH6bEGiQPxglOv8
E9GuGGKRM8JIikAPXJ6BwC3klKiCQerNqQfHOeh46kBpJiSrPSsF/WEVIODjWRXJ
k8gi09KrOJAJdDnNhecG2mBuRHa3QBAX7mkQ6m9450HzjKCBE6IUZ2W8+hj4uE1R
sKxsy3ix2fyLj/jYl6t9m+i6pp9fKHKRQgOhWDGtIi+e2ef3eHHTtu1fcJJxBNJl
UCG7Eu2m5n/nxxPbdoZHN/5ReT1LaOl9LcpXx6oqnxaVBWmwzubb2dPCc2oHNS/h
TxWjrutEy97nchHhuCwnIaZ4tefpT5u+lnR2aVZZbL/4ER4XnZSNYp2s++iAc8fE
adOopgTD+2TM4dBoAY71lVguPMB77I3gvn2MQqjcFXiKHJkAH09GJiJk8/6j6wq5
XP9wEURQnPXQA+tiWoFinpcsSF16E7gGVe2VSP3WMQMPIYPga822KinyrZIWegyq
AgxR0/l05KW4q10ugaTjLSxkwVU0F8EkYd6zd7Wkq92fXu0KQQ8+wHbDBVwM1SWj
KmZy2jOhfpUmVjgjd7QVsepfLlbaaHM6fRDzFnG55b38pbcOawFq0vvbaDfV1XMf
KyIPJ14eD5dct4fTbORdlKPa0XWMu0vETFvu6gBQWoi+xjY4G+g6LIM4/Z/p97WE
i9tT563kMI7/0jak+wG2APKnVNw7kdUCXYSJrzsdBGY6qaJGCoUpWrwE/QZ7MWrJ
5yyUSEH9rtfjLB6Eb3UBMCkMgrnU9z8XlltZQzvzcAsr3FD8iEJM9YcD36u22H3y
6dC/z1j6rJnrAxxJyxLRvXf5ebEBSbWgBWIes3/PqrThhiLGoXPGiDeH8769oxt4
Grr18RJ9ESciGPdSgLgEa4+B/YHhRbzrvLxX4UX173umvw4CXz7OExDu/eaYd0iS
zRO/B6xEJFzAR/DpinCcFY6ysLMtn63O7DVWDzqQhxvFNFKfDiSqhNwnaVoDDfVZ
LlybqrbYpMZhogOlVL30GWrLPdQC1Naz3cpTswXSNUDoyH/fpIucJEv+FxP79xU8
tDlq9rCQHFU3KZFT04UPX0Li9qUuZkw2z92FhzMj5eA20zNsuAKDWJb+7QRxdOxL
IZ+7JihoQaqMUPTybHgJLCxJmtBnbmuiqEwq3BP2L2tNqUhJAl036TRFKCxsrnXk
k0kF1F+ZCCGfBNCBaOmODdowzaub4eg6AkkRGxFnnHYPyxRdRZeC23zwe8MtL0/Y
xFVZDlYOQfYP1ERia65Byb/yzCNQa+jP+VHqmKDAmxkzrbphT+Ksyqf7F4qGxku4
0Oo6XB5RiIp51a+t0kK8Mzcou0vFjxGFhV5SkvUE67I7XAFLuHEcOCwTP2nXlT8q
C/LbxAU+tdtVG3Kut6/f+eMf2Km6Kal5jIptBqq+ZVAzJw0oOR8+ToMBM89vtp/J
PpEL065Rs755ABu2dBP29k/SfTP4MtO4tEl1wKO6UeMJCqPKJV5Cq/3goS1gXC4c
aeq4dQUrvqRokVDpWSlKcWiBth9OvhmvYZ4ZBHbvpvU8DZw+9eX0ky9i88J463te
NcTV0/VQzNwxwdUVUs7xkjIpEu49fiTGDxJ9OB1AlqVfa0zvSNhBZtcxKy7H5hqq
bfoUdhcUiW+NIYhSI3kfS8wcmW0WfC449o0iLqFQAAePiWItLd3JImuI/G9uYdPf
sFbTkkaWuH2ed+3KkFj+XgvTh7IKcCiB2kOD4ofxKa4SzXcBe48y5cEELzCjwvK+
g9NhQpwF3H8kUqrKB1wlF9No9iaDiNpx3S/5TEU2lrulR1M4MkryjmpQAZ/qV5T9
kE/FItJoVjitlcbZYjZQjwLve6S3hNH8VfBTqFlWE9qJ1xpBUbE80cHEmHtU9TGB
qDVhrwafE90lDGGOxeaRfmd1gE996KQ3PadQtAoe1ezV2Myqq4XfSfQarFcPKBYO
XwOW2EFP2F57f1Gff1977GH1ktRyp/JLdYJzxZ0dVWTZXGPNCgfn6l0vHL4CIkud
0YArNagX/ZCmaje5LGMX7DwGEQ0EXJajEt4JTnk6nXg72yxKcoMswOBzb3pVVdVF
i9+3nazRdW5zhh/ReN1M6xJUywF1eJu4d8X8ZZFXK42wltmqV4/vMilIlP1D7XEO
iGXNn6HfMWRi0xsJlMnNv42Omx24dV3K5czMVuGSUF2XYcZ8zBfBfzo4y2SfOQY3
373C/dHl5/YvAocJ0rcmnjGip/f0bXhn0u5oFU7MiQX/ZvBQ0K38L1Q+sWgT/B7f
+1Ed9OVPvclhoMrkZywjm2ri1vMHSN6KIe+beifnLIEbUIYVoD8UHfbFVYYzIb3K
o16e5CNOY683+lqT5QqLXGbXi1yArNDRGKttsr0yv7TtX8Lf67qfYu3OAowNvOz5
usyLKT9zBGXLsPfqfqLpKfRVhZlbsxLhH4DYAv8tajJ+8ifbKbkjNRRQmv6PQpaP
R5OMqQCfRR8R2An9wXPX4EWqFz1ypjR9aK4gm/DJxCTmIbcUw56eRzwTBqPDaX48
hQgzmU+hap2zZpyr49+LY4eDFGKHGSf8mlLcZFbT28xp8Z0unDEDFBudg8PIsQAW
M+VgLR/t9DGmd6m7OgQdqN6bp3QjtoRiXaBBDfg2fwfa+Cq09ki/jsPb8Q4Z3pRN
tEnGxXsLBDsHcYbIGftnHDMbLv3NMe3qymrmrj/MNoMdrrFI0amNx3FVbwxWbKtP
Uc+/5tNHdcM5079mLyaD/jNtIE7MJowAcVSBFGnxmSitApehE1ludqOg+tNq40Vh
nhPaeq5jOwKbwmYKp1w6zFEfWrrpkPQv/ZOfNuVaRV5rs0NXKYfYkxL0y7Q3eNPv
b5RRe2fkzMPjPu6gQEGcPnoFC0BTLT0RxMqtzjQvvGnxj24tL5HvALzKEJyHgmhP
ujDk99o+gNynOdhl5EGjBtySsJkFjDII9T+/ksPsjhm1ktLM5bd86gOIBL6oL5Bg
+B7QZKYPGYGsUNn5CJowNiOxRXvoeDRIoqv1ODQtVRWJtLiUZ36Dipbt6ak84mwU
nd3CASMhbBFS0SqZPuDiFFpBL4eed58Edpv8pNdp4Ff83oNxaatdm4vxGI9+mfyv
KVqTNPzTy3jWMqLa9beJp4mPAz0X8cjd6qZaUvtGRgKDLprRKgWNMrwkFmht2zmz
lYUBTtjeMjLgvS0Dx9D7whjBC6mC7gWPtoZUITD4vpxZIuMPpOJgkg7eQ6Sd6LIT
c4C/QoBIGB3I8M4gk5i0kx8wqY+8bznnIDQcrwtUlXaumJms2QXph/3CQ7O4TfM+
9oZCg2von59I7HAxn+HXlrEzOO31wl3EUfjJpUz2DmRBevGgd1GOOwKqQou/pmHQ
5P/1GkfYz4ErakZsDcvW0UpswmHkSWJLM8QkbAV0Oy1Ua3g6Tks2tdcZ9HDVeLHq
mekGyRMKsEgQmtKZpFkZgfrxvU0/4qXVOp62Otj3adEpxx6W+2qb8Go2onAV88aj
ar/J1vSQv0ZYm9hwYyGaofTBFRM7DHlIL+WqlLbySOtuzSINEjUIPLxHM4l4+IJY
JyO4/bRYTiN9JSn+xiaskEyOvS+LDITbGe4CweRR3/uP8zoMfG1UATxviTUCpfH+
kufYtH/QBe0pO2G8PmHmbUbs2KMlMafMqvDZrUW3rDyDVqWU3ptN1B/9aTyawShI
4c0di3QzPD1RWWluWBYOIBNL/3GUcw9ZtbYXn5/J8j6rb0hPWm5N7gtUUrNOX/b/
hxFRIaHcZ5tlF7LR6M/jjefZBcTPbSd8tS/BwhsJDtJwLL4c3UGm1s018o3w+VVy
SY6t5gP0KkUUZStUnkzniLA+Avhlm03aRjbXIxFrazdbij4ViTdpq3NahhIYCORd
CLDcVXcViOkpvD2Jp5lQ5azngT+pz3ibPnPLbgaq4HNAM5PgV7BMPE1VW+QhYPIi
1XS2jr7Jvd3n9NltoR3jCDkXerz0bHBIs4KlfsBKLeQ/bR88TVgoKEyMcyFCgr0E
02qtw3xEWD1J2gylRmFBdxqtl0BWSiZmiEozNpuIVdGfs7LZz7aSPcfk4ukwjN05
MfIj+OK61KdJzZPKJZHmKuhwNSPe4TJqfh+pLHEPkZfo+OCGDy80vzJgOTzcToVW
a99dGqLlHXWXmmGoK0/vs625G9LNt1ppXBvEZn7miCL06rXKTuIRbBwrLoGQxb+x
DoQwpE7mjIEmrux9omy8jDwZixMCgYDRS5xPndNJahhZ6Xu9I+eYljSbO7XLqaRC
IfQs4UwQytm9cPklv+rfpNK58sxTxN8uDlSttwxk7it/dfRYdhBmrLQAzLPsC7Bh
1elHo+gHljFDxEal4sDzLjPe7Wc+TKFyyKqjqFfkjkeVKsw5jqOf7I28P7R48k8u
BpDohiZAOuHDdH/pV/b9YVltepJ4s8owv8eUS84UPSoCnwudCFJ0uOBd3yatpTjH
XuS7UzXRZg6Gt+Z2DSk87P1E/0lClHHZbBBYWwt++IYtiGL6OfrMVi+zdhacetm3
gT5aOrdSkzQMsFD2xc4w6vxGZvDoWTiAZPZsxKkM5dwmY/j52WsVNyh7cszgC3IB
iWy3G+fOxJ0/bRYBhLALGMiPIFnz2wjaTmLkANFS1M1hXlsbQ8zjH9QOKTWIE60r
8hJT0gxavQk5PMDjNWEZ6ZbdXh3CALpIruFFmaBdgGCweHp+z/CcXwCofrJCiAOR
gI97V0g/SEjbYKddvIbPnB/9E1kvPD/i1t1uaaHlrezLu2XBKHjZ7HVEY42qKR3R
Aky9tXd2y+2VyGxTQOqqUwQlnQHWe2NIE+V9qm6wLL0yiq8T1OVJ2PtqmUovZIVm
gS06nuHaRYIeNpIeM1A5mCwz5hKUvxGc+dNQUdvIcXP2piCcDNATTAlXp2xNqviq
WAxIW3fkrxa+SzbbV19uqrFfOqtKhwmuQaJsj85tgRJ6C0oYaArEHc6uy9JzQeEH
heW7Ma9wFgbPgWZGpCR+CuLZknLt912ciAhMp2TTtfY3UOmAjiy2l2k5pTIXM7Dc
sVHzeb/FR0AA+Y9zPWSfzSnmNUg54kQNkxaFw59BTRW6693Bnluvt/UcVQ42QTAl
7glYQMzDF5mRTT7pQyyN3LRMklFwfOMfXLf7sMfOv8qhrKGpzzDgFo284y/FulJg
Z3FQYqFkjAhiCVtPP9woOWbhdC9a4c9beDlhjl35aPHSKd2/Vn1frXeI/siUjsWf
/WVs6+i0ubwnYlheqmHO2fuS/2xPaOmrdfekjemQRWV9bsE9hjwD7N6xQHpPYk0R
E5Ki+RNFUM02bnBc3GNUjl+6XPpi3tKYd2mJRkSzJxSiKWmmGJ12Zs7oYQ0S6Ltw
Yn6s8IurLdncRTS3JhQSLJChmf5M1j1iXvpFBeCiNgqQ8sOG5DUId9cZQ8raoY9n
gXKbv/uKZx4nq58B1BsixRr9kH8ZZt5ZwlT0i0gNxWJT8olZPqzoRN+4xVIla+QW
bh7SbvnxyXijbHfaSYu6q0mXFmwTD5YGfzYwoBeBa+vp7UNDCEir4RRZOZuo0nuq
k7p58OsmR1YS85oc9S5blPD4Bta5ZqVsGl7+PMbq/WEje8+ARYWb8LPauo/MjnYh
vm1yrKeY/BR+2zLF6fjZkvBXV6xY3UBalVdv/i7mDWGM6yWhzhRfcOh9E01k7Xic
4FaCXRw2mUmcwUsiaDlq0QlNLmVlwAxZUW9TaUbV0kpejYxk5fWLjzkZ0nq/Q57K
Z/52y4H3lPBWXNNhmlEFZkDRQY7wxbemNysfRL7pOLDKiNk6SZyFSqUAlhwSmZE5
P+BBPFBkvDRXmG1DQ+BTkAQ56QOdh7wf5/0Ch6Y5XILvL5mActz9V6JZPNTDJ6TT
ZnfVDANPJeIxwPKgwByt8L6gwQc4Rdvde64upHAbtYiAWJGFc1iz/sJgr86HiM02
hYrqo5VMzb+Sahc8fnScaiNdopLuHsWYRIXnb/NqPirZ3q3QTmS6r1eNt5n25d0q
B4iYyZVqQJgbdcJVhs4WHqxvSYtCKI3WxDcGGtaTIWDgLhq0NtyeYn2hUxbUzo95
KbDYniGVL4+HuDnhgRwumWyDgGUfc5/YZtUqOf8GQsTteUa5mG75VP2K+q+Jhqbp
RWl7wP0EXL8zJEc3uSyG7ostd4vOx5Nptu5Tu+jFGnBNnJXhNG6dO1dT773QGAgH
RQX6oH7L4hztu0Hv5PAIQkX8hzuwug14gOhFVZm6Ff1vW55VtU2YIFxFUg4dknZC
LaKOzOk+eRPDjPXEtvYST/RBdPAdLXsJtkbMqtcY8m7N8j5pZnj0vbkbcaLXSXgu
+6uM7rgLQl+SGQ0ifnQwoSP9CfL5ehNL9HxCN9Msog+XbDTTHw2vOp86/4Ja0E6f
JhruOD6yWo59nQAIcRnBxT+VKnYOVJSEiYnMyOJ0VaiyWIvFX/uLDwKU69n4XQml
5ezpTLFBaqeWSLvIP5Mlqw8/hctqul/AKWrj/MBoIVMCoiQlVDPbU0lObP+1416M
yYX6ArDgFjZP3S3j/mbpBt5hzU7zVCEZ0X8bCLqSHRPXVWwO+5D0Gb6fKlq08acz
R0PkUhIIqENXf7A9qEJ26S+kwFrsenUIRlEnSpo6s29DL1UfV9a30QucRgUPmPhc
/z9kXBQRqf/a2iPJBvlIttB4UAONXOEtJnKeqgUPjLpyfGKMPDHWCC77DhiDe4mC
NqDDaZIln6l1YiPVbmA7NQX8gSC3LRr5iAFpF0ILu1uwOAtht3ku4F+49Pu0Mdhl
mLLVrsof7FkMYumhI6nfqwqZCuL5kKUKK10eBWZ7sq4xLY9CxIZKAqs8NH1Pkis+
2L7ofchniQgc09B+PAZlcXP2SmNXTs4JbOTxohcoHgczIBtuJYbp7vRBuB8Ewm+V
cLIeUEnMtuyHNJbL4Mnb+v2bOkI95vAeW5VM1HFKkl0puTIR9Knb/eE5Iql7D/Kb
Mx5XhCBGYpRbDq9GX5UzKKaBjneDk1E9GsdmPzOP0xbor/86GTsDOOg9JpzegMoR
7araU8cFmufCmbwxhHrpItD+od+WqP6kLzN68p66rWu0K7sRMdlrf0dz12WxiPE1
qH3fDIQrwVim72l+ZOZ3OWtS2gE+IOzVXn8IB0vT5+0rBOmOQ/fufY03xbesQz2I
i3dOOBYkJSbI0oUIlz8YbuKz3qXvTdPiH7LXso/MrfZF2BHhtxww2/P3ghtF6ZSB
TiaTBcVmC1SEFophP7m4Ea7b1DbvoO3W5a1SFNbH0qexoiNWr7G5REtvhqlIGWWH
K1tWG3xnZdQiybsAmO5YSvz5zvCdThWvp4dJNuYETy0otDEY7us6UkiNtu8GZvJC
38uWNtQ3Fn/mNCP/e5lO2N+NtpKykrm9Unddy2vZV+aZdqwVo9xKbyLTezQYSA61
PMK+AdxCHrvuuimxV8umT2wk6h3Blgc8Mcgw54+zpDP6QSDFuyaEs+WrSmnz3TGy
Mo68Q8VWKZ9iHtOoIYMHeR8CzJlj6+1Nsfk83DMv4CsJdan+u6yi3rbbwxrAQ0CJ
ykGcqu/d5o96eMUk6c10f+GCzTYi5NYVvtdALCiVoPYBg53LpYtvvqUdqrqIgXrN
Up7QsgoH693/TvCc/qZ6d5yB/XF6kvi54ewIfFOA3PNpScPRgNkYkQ2VVn3Gmwfp
nAuDb08+YGGw5WFmWKrxz3ZR1LeETQdR5awbtNrj1alb9t3Xbdj8vi9HebD8qWb3
EC833oDkdR6pLA0X/zzitphrMmc6OtWPRDP7R7Dm9iz/BfhYLtWUVolJzLRpFY5Y
8g6FwyHN5MDsaJYxYYmQ/9cXazH4qs1apNwB/rDB/hRek6Vb5+9nB7lyD2r523uk
HOg1p+UrbAogOgiNwlX8aLT1vCkO96XM0GQ6KpcMVo+nYLqGcoqBIJZGmWOYaRWS
h4fduCTAx2e0y9dvW6Csizp7mWeX5thGz5y27x3v956Y61uF8fk8OXIst1UwaoWX
4ZoLhjDnrz+BD8JsBTs9CzhFMZVbFWVaI27AdgDJS6+7KwFeXYnYe/B5+UrBKyXt
3MxNUMjnkubrZgbTVIiKsvy8RGEPKzb6Q5SrA5z/Wg26brCi2K2LCcscmQePrTW+
Y1ssb4ytYYKFHQu3oEiqzKWDEqaeyVBzXxRv8QC7Rxjj5ClzsOO3I5dVQfBWsKZj
w+uwLpFlDtNPA0gc44jKl9DsAXmE6zCrqvC2wdKIGgOOKMXjmDupeCL4izEv7ptf
y/PrrInLh9xazzrraltvAZKoo7ckTEwh9ux+4UceHcBYx5W4WIxXv+GzzgBAZHw7
cw/Xo6gb3xG0P+c3lvqcLwGj0qsSWe2Sn0ZkpUq+l67ZYfCLUC41CDa+WaejdCd+
BjkpU/2GNm+dF2m8xWVvzQ/s4/j72cSaURJnG058oyaTlwp1lvaQ0YZO4mfKpqBU
+Uwt9bTd3cdlATZ/Jxf5xn0t+9yGZg1GvSvmxy3DLBGF+HxSrj+6q8WxhR8LvpJ+
Kv37cnhZuy+9QKa2sNB3SxudgSgHZJvoS2hnsIVnB/k8FAv/sp+pAjvPEqsXJDr2
ijdV+oFPxt92A6ACzvx3eVVb7GKX5IwBC7AjVySE3rOfut6Xg4mkoi3gRNbtdvBn
i6j4Hwc4mNF6snAa/OMl40YwVP+XUhU83KVO2mZ/vM/sBRLQDB6SGZzzRX72ZfQr
pTV3G3i4gopRaSWm1lokHSPRkpyomoi6CeOs7gkivyhHveXAIbVkWta8q83F83L/
8DQ5AddWsL2pptaXOf2LhcaQjaytUI+eL21kWQ1zsdxXCW1dBZTQz6+uvdjXM2cW
dtjntaQEekTQLAxvgZAeavh/a1exWP3aGvhG5xJjti/XrOqYyuU8a3TMVmYi4Z7Z
jeP9iMS5FHje6bIlDvFn0EQDUlYWEA/yMte5qdXbTD0R3cQwVkOutbygGoxErs7V
KmBS4UjfxZ+7q1g0HNXhCr+pi70UoG7GGkxuLHwk2+Z4xaalmtRS0Z1rp6SWsK7e
jq6wZtpUEIeFvKz+CX2Td3Ahi+ees699anxZ5xnul9O87D3FH9TyN9/xiyZcRFq4
RIIkDtj44Q49jg9wHMyTg0nmJuKVBUzs1u+KMF7Z33GzLUDq4yhSrrSF2/uxHpb4
DgED/s+82bvHUN3zNL6WUx00HMoMYN2WFUt4xrfqFfMdM2raV7G4dti/O0Ly6wIx
UkfIKblLeIiLB9x64REHpo9OZcki/NtLOejiIUc1FGRnv8sutCqi6ELqOK9bx3r8
kJD7nzQpYBZM9l17KO/xCXit4ZAhgIfl5/5+eGLtO3CkwzVjefJtjZRdzwyqEA5l
1ZNmADgLxi116DOoCtBCUzvmSYnURSs0CYRcX35wrT/bo6Y00dXopgW6JyOCUKyF
WRixIWqQ7SQNBPaYzcxyG9XyIKESQ7Hb8pM9xAFNQ4bJdpLFq2cOgw7JwQgRdk7x
FUJ1w6vEnc9vaBlx6zWftzC+Gyu0y8mhhzRP0850Ig2FbWGxqh4cFc/lRDRiy/UO
Tz50aEPBVtRUlYEcSgwUko1yVpmMXBvSRXd9R2neoLd6zZrwirIL/H6cMBhEh6id
SnhQHkYvHFRAHWKqVp6sIprYduXAIJ9Kvj5oIF0EvARHQ6GPAlfB/sYAPn0g5twa
Mb0waBeywoiew0WlNmx04+i5IkHkFTYmn9ZDf4DvcFnnKEGLOM76Y8NWZh2DFdOa
xDIJgOrrcZsNqrO6g4luYEO4vcH1Ji7ydG/7uTG1Sw6yMGwYFO78tO/yZAhcS4DK
DE4SUe0Alb/nwOOIX9eimFufS+1dREYywyd3cJs7Eop359nEJN9b/9lz5adRcHzu
tgU5ba/INbH+7lOzraCzFeQd498IZhg7nxss9+cUoAwYGAJ29nGuII/SZz6ydA1x
q7Pii0eUhC1cDHjf8JLNufaITcCGLKj8sJs0Y1h9DJwECwcntBKtFmico0rZLgSs
AmWFmjj6eh01NcIFv5SaWJPorQYnQNcafhaWIm6w8GPqIH4JVpIqZ0f9CmEV7yIC
kafUYP1x9N90JLm7ZsLqDGONauAdFZfDxHTrIAWW4nejSrh2GiMVwhl75NYC0+AX
9Rio9g+XaDhOFSQKE/KmNVDl3gKZUzZBZ4/qxLeR6X9QeGXFXCMJotQujHJamHVr
XVcXwsYiKdcCZlxMS1QJraA+cGbt6kxmprxTCnQK07qkGx9cpEPRkepKBrw4ODgT
jBKqNQfoMIGVDQIhMMKVsiPV3/nZL13FBZXX2o6FCJO/nj+AAVv7FER8hPSJX8Ch
bTPhAKbEtXfK3HKGg40F8oI5cRU1rfuBozptHkhlu5X6hJPsMkNKijH96dtfKqWc
JmmIAFyKtStZBo0j2uR/+89bFnR8+ZS9MPPjJVSiI6y+Pm6/DdCVNFN5VVOJiHAh
2dyKteyxBrnBSdbut0Q0tNo5h8wRIxnB3pyTt04WAeaAFje5fgpQ7gEFdQoSX4wQ
PkFOzzSGDYtYr2dKaTE8toQHqoVTZ1Pq4iBIdoaT0TfV1nR1gxB7J+djwMz0Pjav
ocvxCJX6Jd+3GPYHG5YG3n7KjN5HvObDYGkMbpdOushyWsFYfcNewHqsQ7XrgU0k
ws5e0khUvMkvIUC92jrxrUM9RQakZygdGaSV8ZOaamG9ItnsxWmlkR9m1OzKOJlL
KLRqcPmxSsJzQVHX0o7i2dI5qAZfPti8KUUGHaxlCv1hgIMkAUnQNEPnsC8nnkDu
CC3DyOCw5T18s37uVDG+GO8upSeiZMYlkhSHWwtoqP40IEeeMrxiS/rPdmiJqZpp
Kuoa7IvPBGrMWtMAQmU+Y8TV50Sx1o5zs1KvAStzUcbPPMykau1p5S3dXnbuGxsH
vv271TIcGz/Qloc4ECbHsKbbKKBjPI4JUugKCQyvTH7BeHzqAQ+UfqIMraMiAlfr
02/R9BRkFAcE6XA8wS4+nGwkA0OoMx9q85kZcVCfBoeMJvCv0RMZWUvZ888jNVYG
ghoX3XlzwuddxtCiKOt1sKy1Jte0YV0dFjBUSbgkE1UIXQBzGNgCGupuheGQeXZB
fsMw64ML4QjeyO7FACvkh1nRSCNJnIv7K+TQWEeHYaruf+dTwGYEvUvQciIsMpRz
gf+mM2R7QXQP69EKwkS2IMvvTw0Vk+hiCW8wcvSGpNn+r5u81I6jHbtZINvZl6zQ
6sNwfFVH8yIcJbGbrcsnXFs8e/1OLrc7BeA/NjRjBQBOVeZkMO37VM6msrnTG3xz
r3vShCpQx/j3QtweDiC2xaJ500yi4r51yMydfEzXG+7mbE5nNhGvwIme7Ay8TRsX
Z5GfnxfIjaW9KprXkgh8FQ0jVKqqNMGgBrSJTRutXUKS0omczT/8qCK/PlDb9Pp7
WdKf9aMyeEUwOtphQaLQ85ZOt1hyaYY/Ew0dEs0vYlDKTHPK1egcbNqr4GjOe0xy
26tN5F1bmFdNl/uBd+7b1XsTyJYEdX5O1Hlkct6riUFHF8CvCBAvkuko3MEc0kUb
uIkgkKSuZZIWawDc+VEShtkH21Dz8s0CtEZvuSexzfADJ5T+UhdaW9PvibAn0o6T
TySvOgmnfdEpHwoq991FFzTsuBVl/fQzmBvnuaJYIF51Y+d1SAWPBdl6HiVCrSzJ
NtfqYMFVVYshtgHSHNZ9LjhtoGY9oECR9WiloQR9NqMi3I/Q1FJG/eiliStnfF2+
SiZoFYo/YouwsZXy8OMEXKQEl8wQ3bw6VZzxd8IITH58zxvbCbnHPJi4r9GFud1r
97GtmrJ6OL5SUcCrK6i4sPX1yapSPAFrjaa425ZgKsfiqRJb5e2RfDLX1Gfl9l92
3UPNRgj+yXKI9ciNiCjgBx0wZSrvxF7glSyBQOI6U9e05UWpjtWjsk8jqHdkkXn6
06rMnTL0u3XveVav5Qm+BjBrPltl9xwO/YitcNZzy9QLCC1Dv7lZGh2Hr/F9UrzS
uAP5bQtZ1iHpZzBzrrwA5CTWWwLPQpvCRxgcIIngrVDnZcVl6LumgS8CgpZPukp5
A4HO5fDsB4u4NKtjyev+UkCgNPEdguWdS84zLTs9hRDzNVkp6oiB/0TgHPEJ2vzq
4OHstY1jc98dekyv9YDescPCR9tHy/6s0KzlYqwRHLDuwc6g/+lC7Z3iyuRaQcGh
5YzVKeq+DBXXloez6nwUVCMSgiRFsJUhlLBNiQfa+kYYtjVnt1ZnkoCZC9XIsjvA
acWfO7lZS+NOjAFLokf5ye4G3PqHo0Io71NYy8qJKAP7tFqpF3btzG/s4mHAPw4i
W6xtZ1DDk75zRNDQ+x/KkGHtcefBSUr+hAMa0XK34yynF5lGvnz+RvGYtW9whoY+
9zDQ6V6y4l44gNhJnkHLrhu2yhkuDeLp2JKdzQS3gUd/FBS7lROlcVm5f7CfY6s3
3X1yGuB+yiolwe60lMOP7koWEHnmDXiAlKRon7n2FhLpp0G6NS4+49XccRDNVJRf
C1WBlhPcBbciTo1LbR3Tht9MHtye8T+iu1fqP0yTXcOM4mtU/h2Xpdenp4FBp9K2
lxFs1wox0O+4bBJ+bv78z4cguyQ7yd4OFfzZyNM4VqRHvPZp62vsm08E/VyXumJ1
0MswHtW30rh/TjlKziWltgF3XzWAZLQdlWmBv4BemwoRXKKad3YmNxOEbz4QpAtK
mhDPNMd+0UzoDqasDunUq3ahO4IZ1lP5cE8fEqZ6/FGj0rPkmOVeb1X59HYxV8rA
irfQIc1nsv73NqxIRRCgMqs4HVUzOo+H59pmUq/be8YDN+naxKjituwqf9Yd/0fO
R1HI73OthzBqKyNk4WK2a3H1Zy2Mei2i91HmCbirq9Fi3/W5Vwhx7fR2rYaVoF7V
d33eDMHXTn+omYp2gBR3lB86OkDDbh6RPaQik+YgNWjIIPRVM5+84aEOWMh8XKl6
kyGmufrIEUeGZPWX4Ey3U6NQb+kD1yEEDoharq/O/v6dk+9XihBqXHe1FDOGRExo
EGFzijkF6G3sYanjTFAkwn8I8FF/ElttO1acRCULJu8wjCbkzr2qCdAPpVQaqIkh
bWVwIqjyLSF5A8LnwXg7fUYpAJsIsGVHSQruUweOoVeBxWvS4syI9wYK0QuU3kl1
isysXvNQgfkt2SXcTRthSFitaBdgg+nULNKP7YMWXOwaMnWKbX2sDS/t/GquIZu9
oQW+bogoajqZzIjri0Qqdp3ARn6CkQDri2PU0No6nGrRt240l1a50UMeDKJ5g4WX
FIe24iCmDkheRv+jNrJ5dV/Ad81NBRPvILC/L7z2pUhY7bL2ELoLa9Lwd2PJ4Cf3
L6w1Gno8lzd0x5jmuY/Y4OEVLfOJyxvkVV3AEu1S3ceV7c6jgheDFjOLHTYL/dKJ
V99Rt0Ro4/6YFMdh4ADNrMDruKeUgSNJiKO+pjvQdVqkWwV0/ZIgVEYgE/zdnHue
G/Hfe96NWFYoZCyBcZC7tfMDAu+ECJNIqPBqfg8dg55Fc51wpluvO2az6XLDmGYL
5djbopdRPZceARbTUsx5XGIZxhgxLmPoMDx/j1igFvFQs9DQxXpAhDPfy4Gr2Q65
Ax+rb5xv9vgEMwbKQRsYG3+imdWe1PEg4/EgnX3qmW11fVjO8nlZVTGo9UyRFTCS
fwB9b9zXkpV8ji50Px52iQX74uRPEPasc2qD1PKEq0dpB/On+ff+hdi/iBLLIXxz
GrjlCLAweZuHRyXwdglKQtp0Y7w6H+ZBOK4ppDobrdeFPfGBe9etropCQMm4gPg9
e/uZIXOd2JDd62+GJWNpKG0HJa20UYyPO2zYSN3pHLNXO7HdiJq1cQ16k55bBYyQ
2aFXEjhV9l6OErG5dvtwhiodObtwvItV+i8XqyrgFd1thq9rJ36tvMTFNlo/Rw6J
xm9OOe93d30R8i/lEzjqZjHDk0DoZ82dh437gvpyGmJz6GoVQOdFWlpLpiJEEgHi
Bhbs6lIik0zxAhA1nH9mXJfrd4cI3SgjwN4vLu5IgBO9kt6aIw8m8mFhprawPpuS
dECOh863xFFKZJBsYzVRNkn1Mc8qR0daLY+CdVXsx+PV1XVpGpjEYFpXh4Dqioxt
60k2XPzDEnv0BJvpq16A6MrK/3SuMpbNvvIgK14KPEyUxEveXN3JfZM364zdstBV
b7n22zv4G7qN6F7Y/dvrDyVyXK1Ffg3WpiIwUukm8Tj90Eo4d4XMx/eWBqO31lLz
8AtJA7ZNHLmfcgJKiQDpZxp4JT/HqSIB8pmX9KxQnSiN/b4f23RAEeJS0XaiLOIF
CZmvIWaoraN3KfixlkcqsOuEwnbMKxJJJpOjNQ3SMUooVayFoVlEmxbL4lKF7AJM
VstVNBhM1YOdegcjw64tqZ2nc0xpYiuCLCyGAZuxStDD6f9ND9WsF4kD7AtirDZN
CRov3iUlFbUhoSFGcZYjqoiT0oZgYvmms0wFgCBI7YUQdYECQBLcSXyIF9ZTh9cj
P9RkQOPb0xU94Z+1Jfieoh0VGUlKvaqHsgTjHEqmMyPoJhQzUbjvawg/cyjbD+S9
EyxplyZxIegOii5ZnYSz0hDdNIhTD+DFspSS1EgDOEjXlEUA/G6mkhsqGWSEK3uC
210z2oLXwOERi2jYLcVdY70O7uBO+cl9+Z8B04GVesrgZrrr4fWfMe9u0vFdcrbZ
PNGTtp12RdfWX/XpTRLmAIYy49VnkX595DFpG/u3CXC4qAQzbg1zSxklIQZoY05d
1m4nGJ1cMi0IP7K1OnWS12LqwbIo6sFxt7xE8XyLAFtv27MuV92KvCf2amIBtm5c
r4JCFOMsR3OQq45mpGWUqtgVORqwqsUxKDcWg6qRM8d69yNKcmqPp5IRyEa5od1A
GF4ibA1hMmHzdEwhBzKVh0aKQL4byqw7PudB6YwlnTGZ6TVDr6oFEB6o1RTMpJod
YNRJNVmMv32WvGVu2bzRy8hf/jcpF41r6xnvxigaaXi0fbeKmxNU4C4CFqktmOAd
voNluU4OFsdl+XkpHnrZtup7r9zehckOCZ4umGfaI1LVFQVW9i+bV4Xdit/1pG7Q
hbjJtaC4tGUkI9A9SjYnYr/f5AmXo/EpRapUren5x1sxU6zEbGA3BFRodn5fMyfA
vNJR2z8TLUDIcrJKosTiNqkCJ+3pKW3VvEzflTOyJoZAMtSt93x/Qdab248Sbevi
NViF0p1BoJmGP6L3pRWsEI0Za8KqmeWsOR9iTF+Pdb8MPiUIQzrw4o7ji9MhQaSl
cpRrgBFHaclwh98Mwe7ycUZTKUcVAXRiniRpbygBcuA8B87d+sRUCHh8IHkOiwY8
PuRJP6nQt/mlPmu6h0VLuuBMlbAgfEK7IMpKh5p+FNWFrdNmiqEq3fUGQzlcr7gi
ERhRT0iJxr0LnyaRuMBweixKjMOWruVAAGGBtTvd2VXGj6/jwPPDXN6HIwEI6Uco
moNqYTc7OjzUcjA3dvx6X04c9K7kkoZE9+flt0dDcyzRFOO15hg2/c3/Fr32vquY
q3z6FlkvgDs4c7dHl4hANAfKgP7j4WXW0pJcTzE0+wofylJulwesSHoXrna9fERn
joDXRWYmUeUUUpBzMuvS3dk0t14+miRB/itY4GwqCYRGSTGLHmEV1sc46ZzWvB3m
jLDVxVjuHnAvyu3kckmxq5wLyh1yYhy1Fa/D6s2+kvs1eI59P98X8hyxSxbOFqm8
kZ3sTJCLQs2Jo9IBDQerPccCtbhIfJUG3h+trUaW/4fi1Ep7zvImiCv5vckUTH5G
S3lAHbqIMnD9R7pZ34sQR6mjOVcoCOffF43Q5PIe7ZcbUkrdtxDaz66VMwkB0pfX
rBbVBCZh+/gG3dsoz11xec93Wa9CDtSXmxPJj1S3QnBX1k30+FEwuQT7BLhpoU2z
qZlfAhQLyH6pfRQRJ3x+2+F38xmSHm9BE+yI5k0PebvQHjIpFC/cJOxpDGGTx+rH
ivwNnC4Xg6Mqn6TXq3sOUZgCS2m/AlGZMnpDvjZR1MszArW+gFduWA7Q/UbyQq4n
98eB1zv4QEXiTMR2Asob8wPLLXmqsiwufDcsvZoAhf4hktzpZSA8iD7Q7qE6D2at
yZGe+9ay+H+YasHHvtQKJlZkzsFn9RGkWLy7+wwztmQqx0E0QZzdlZMNZDAxYTZD
N6mPW+Kx6DrOcb73esWzulf6JT7K2Y97az3Q6K21b6ywVUeMl5Yg5NsnHieVhNNf
YoQPPrB3Oqx+IZqpdFcZFeUxwyziCTbJMt43VloeIwCxZ2zTO0vd4FCx7tJECQ9Q
yY0v3tZzSXody875mlIxvesentOBN/aMU+Ot0PPQC8dAVwUHAQmrpstX0nu2dGa3
tlmTDn7oLwLd+Yt5/6JTGXcXa3koNy+AAph3em+EtUJ+trnlxl7RoNBLySIYSPAb
eSiwa4+lDxTJuqJqMCI5UziY8LrX7b8AnuV3rEEwJsA9HRRpTh4RD5gwVW2RNgxh
2EC+/lSQgZm4m7eW2jHog80KdZQX3Fk/77yUxKZy0gtZHFvNYsDE80aFjZ1u26OD
A+PaX5jsubyR2MysrSGM+56igSqHUacJav0NoBCve3givt037gFYNWpwIXXIPf+7
ySku334KR9WC9fx+8MJPnREIdpQZ4LRF0Vo4yhxxOrL/wWKL+ubVPUdrXDmJNblm
FA/TtoElox1xZARVnaGo1uJnw/Yr4qDqeElMeASl2XK+bAvFZvwgcfwY2E3Eq82M
lN1UeSDSRP1v+LCjyeuVmUiDScB0ZaltiRph8rk+y4DKPsQodnfWTqbm12RfHGly
jLzk4QkwCiEWGH54UFzQZHc73LQIQBsKmQHYiitXdG6SfEC9pAoEQNOZTfIsdiRZ
h+hMJHzej65WyjsBF3P6eH3+M2f7eIltM+/LR+rvb+eBSSmwGv69PeIT7GiZK8RR
imlt1Xvz9MlXJhjSd0jdd+sMxpS8PiDvd9MM0jKzFQQGwXt3grbg0N7ZrVc96mYr
n5mHJJX6dI7n5CZ0cTg546iaZxxwWvySjmRlNMCUBPTrisy0PiW/yzrN/OopleUQ
N1XbRI28VdfmiTBuPP5Av2ddDCy65yCFFbl1Mc7meGe64khf3izoqwz2DjTOKVTI
x6A1kQOp5feDdMIWwlHMWCxUhOUHQ0vgjTWdn0IimJwgeL8wQeuszR328wyXyzac
9bEtIXbccbHbWY4WzjgAWjoq9b2YvDluc98xxSX/G6EY8iw6J0f0xRKyOSnspyqr
dvkTpsTgFAa9chRldoGLssRWAPUWvEoUf8gF6wTsON3F+M4pNej0R11AKBsGP91u
RP+AyogNyQ1O3NfcCixzO1i2NY1Gy2tDWcjqWIoKzFrQlRk+Hx9ZFTej4FqVKc32
YtKQgbvFESJR4oc7tRcYqC53uHxuclyL3u/GyCaUFghT/4g9wgtfW1qh+fel7Abz
ig5DaFdyT9lOqdU0AGVfyTORaXMfCZI4FkYUTTK+v5Jo+XVLGdsHasSChW8RG4ay
GSu6qX9lv8omfM5oWjXtF+7wUw1OnqCa+EUEmhChZINebDeqLxilxKSdvP+xm7Px
B9NJ6nq1u17YutxPlePxCBQwLIWzy5+RgnEV/kk/ykQjCofB819Nac3scYSwHm4h
DKobSNtgePVtDzCgV8xvcDV23CtVOQpM2C3a5HZmdcRP/Y3ODm0aQXJC1zE+ncFr
q12Vt39jIk5AWdtw2IPTwiJYDLr3K6lcrc3xu2lNNc7VVns+XZ0kfdWLrwi3bq2E
Du1nrDihVcJZtaMED0axHwjKvJej11firsmZIo8GSzjorwd0SAKsib5mPDycn6ag
R8HZ1ZcBNzDbcnC5tr1boOB+1sJePTGfnJ+rDJzg/WrYl+eWKJO7xpaKeKD23A5x
Ghmqc2An4qMg/fyGJX6+Q8xm3CEltOUHqLIIJq/SN3zkFbsTZIw+EXz9rvGLI7wi
gvK68ZeE4cgDtKORsiX7koqPilXYE3wRuXpDAecKwD2l85RwtJXjvXZYr+sg7/FM
Zlw7yrRDVGrcwA9UFNL9zzWZ9qoSErqTQ6SGhphaxu2M2xcKIRnTh2NSQQtUVr7f
n4zovKeFHKPhaPs5fwMwYj/WQq3QiVtyKp1VyNwnrntqB4pNkT+LcJ/brHrXyKwa
VLqNtm7CIZ0jzItckXzNN3nH3bdm1bQgxtPvU6QaojxJYynDDU3umweL6wSmoafv
/SWuHle2aGVJ42mxmuC7neiwk2Ll3CWL+gO4GXe5/o/4xwp+Te28VXiJ9FnUqmWd
sSGb5rrX3afI2W4cLIIcsgRLHHLOMwA/Z6f/3ciL0ythA72jzIN9JxRNIvBqeUdN
ul/WVoeY3SzvFD9xd15ZW2aDJE5hb42egtonkcaXN9HwcHObjeFux5VuchWhaPao
1YyFWUWAC48ai7+ncb3CEvN8Fs0MfyPv84yTdHuRzYP6HfXoQRH042i0MWZAB9e9
P+V7Ti85JpIQ3K33H3A3HT9cizV+cptYuTx+bycyWlgwMaXEOYWcbdyyiAqJsM7w
kihOyYgI40KOrcGEng4IwIU1ajL5Bt4KFfNbiXDYPn854IN5KIfk8OBV5b259ZaK
kW1y3TbHQHR1NxjZ8Ifpd3hilDoevki51JrgFGbcFxD04BSOhna4dugRfa4BZE2x
BhyGPGSbOL2nuwrJREVdkazlPXdQv8efKaPiAvfH12sGYXFS4CLbbAg4VUC1ArQS
4JkLwEQrB5GIo5Ib7lyvoxEfHOG9/rSOIn3KOEBsT0EbbRvF/MRkoLFUfKZxyngB
Mbb38S+RBzcwq6bKPHNog4JOfQvFYPXe0UqbXMnKgrTSqF7wJ80MbcsK4pg90PtJ
vJTSfTkl3IUhgKGvgM60OC4V85ybKL06RT65MFF13hKDhhF1xouDcyDH5Sl0RzH6
YVG0Ogp2hErSt5deeQSDNZ4zJAC0P4LxjSHJiMlNFg/7bF9/mJskgwc7s0csmUnR
PkJ1nfDwuMm8yN5ND+cr1m3AyKaUQTpHIvGNiuoIK62XeQsCkCfwUK+RLNuCk/qH
H3wjzU9JPZQ/9rgZAy8POqU4s9ZLUG1xyfuCnm9BHon3TXD4FT9arYDgoLwJ8vCG
+5JzKDYC+WOd0YgkIhsDkoW6ybnFE/3zO1IWPqoXTCwNItzdYF4qVr8b9lbMVRhF
BgK4mdf5NSP6+MQmFIeyAuFZtm+cGdVHdHMkblCTj4kFHsJuOSKR/H6kfw/PWJ+L
vSYtJ/qqbQMESifJlBOs+KU3vB98/bMdN1MlVQG90cZV2PIutJDVDszaHYucu/jl
V8oCnnvKNrYnqec4qA9mMxz9pRmIhW75VrTR8F7cd8IRTJ93qmVPFrws35l+PQyn
KLYpqNIavLyMAJe9WJvNiNcs/LC47f9cIm8ZZG2dq3Cx2V69zrEatqT8vLLMUbSj
xZOt4XO+M83VOfHFZ9DS4pBYwmjzSg+W0o6Liu87Uadruby+7SQo8HPvxxbGLryX
D0TlptUQCrjmuOXatiJ/LK5jepQzUZPntKu0mhgXa3r771+GRcCzycg3cm+fIBxX
v0mNNDb3zZYUezCLwfZ3q+lBrYdQW9xghfJ0m97a1/fzNha+QDQuurBtMsXpNuxT
eW777LqceMqOVOQrFv4u8v5zWHvprjXLuUbULCTYiBAfX5auBR7RWwWs5TSw6P8P
rIpODZ262wG0vYK1nh0MAu2BO0eO522Ka0rjPaLPLB984S3Ow50HEo0AulsQTYuQ
GGDBSAY9mF5pD5dRfuDOlFkBRooWfM5j6Dxthl1NqGtnWjcSvesWOwZuItfg+gJM
K8YTCpnprWpiSV1MuLdWkX6ohy0upG63tc4/Goq8q0ED2IIIcP1+IncSZqq8Jani
YiH0+oGybNqPyDRMnTvj0R48n70Gu95V0b886VZx1peO08mjyG6AHjOzAwJwj34P
LWbX6TA1uPqL/bfywb4yypPt4wueyVmsAZcmuNdwVkqt5aoyNVBT+b+uBDZ0NbPA
pbR2Rz+i4W4ukwY6kFTIfNulb71oWHkIgUy40Lkux84a6SUDMAz6pay5TavUDYGi
8A6eiHe99lBqTDJFf5EUVrg9AMAaqzyKCVRmtTJx50/2aRniAgsO2hCrhu6rYNlA
fl73GF2Oxc029EkJFD3aChvJQ32P5mYxAIrJDbEHwZXubnXdrWMPZNtDQHUlsh6X
8lIroCnAiZ+247YjC6amGHZq0SZVL9rcyTgxJIWd18owJhyUd62skcCraqjK7dIW
YXHFPNjmLv8Tzf25z5j7zlxFSz6OMRzsWhmCKUazyXp8HtbzQyWvFEf7LcJMOsMS
dCvXSm2SR2PY70Xa72F7CK+amdTsMbndmgpDFXBEDzYjTG1OOj4txcugBYKzWenb
xGEDg7VXs9MVO3HN/VJ5Zloe1l1f1uR1MRgRkR7SJoIPUV9PNW0up00Hca5X7TGI
7CWfpfR25g5qF/j5HyiKZQQh+5w1ajQWRkfRqMzGRxMaf6Lz0cs4/LdYaPBH7gRq
uK4uzQCtkVJ0IUZ7sG5FV3bTOe6GXsygtLaGHp6zt0YaPnO0eD5e15aI5PpL0RRA
RkwJ3lttdAhA8Tvn3BBvDxvqd67ilf8UZmjIIsWpCgvxWj3XZ3rY0yUeDj4A6xFI
eHQ/PNWkuX4EUen/m96oJfLiomowwRuAQPWnJRw4MD+MVKOugwUrncJHXoj2C4uE
rqRS11rEBkSlSgRdh6/CWSofSZnfRj1T3TX9G+ciCNI8OK8ucBcw8TccgFbghIvV
sQmrHr/MIfrun5f8V4l249aesoBNdtU6fDZdTmeZTbKJ9uRz+0DANE6ufCfV24/k
HubQoSTjOLvAvGRh8Bf26vELRtGtwwV0PtxEQwUsEqq9QA3OJMvgT3a9OzibIJQV
YyxhaXx8u84u1X5FxhN/8X4bU9Hi5sGtvYYb31wusiOifk2D6DLdcqZMeMLUl6GS
YDHcQdE9eESQjgxFRgyhcnyfJqVX7C0hAB/BN/icptXxsGnunau1PyhCOqQFxfIX
PCe3bimEfyvgZrGCzIkf/w7BNNNcAoLca53eHXrAYJRowyYk9a9cw4LKsGuH9Ai1
bLYET49X9xNw4jR86KAvv6RjGyx7kzEOKzHBvd5aoBoL3UQObbKKJbpIMgU7W11O
0t698rk1/SqLTjD7P5wD9KAfKDEXo216uqeldIBfzr6BUnrR9I5t3g3UdAIMltP5
CndiIzbGPDaweLhl2j6rVWZ350LWrTR9R0tgVYarC1+jX+W+g4Pofn2Ce7pkZHip
Ylej1BADscr/MrMk8FbvkBP4SLOkz5O1HzEGTf5H31+eCuPoCRoTzCZ2VyXKU+pE
mR+ypiGq1o+nmVpKVtkLuAsi2ngZM0JhrCmWziQ9hzqXsoSSmWWNvu20uSUTVZ6z
yVPrGBVii5cGNLJgyXsySlyABYOlSKotkwRVAGJ7TD+AVivknQ59sW5hY3J2miQT
rbfv8CUClG2qjUkuTTUMMF2ee1pGK60sWdZOvv0LwZ5kVInPk1B457JG/j2hS9Ur
UcvzgYg7Yo4HKex+WN2Qo03DngqPjVpRW3/QYdXI5E+N9m3l1W0Ofk5zdHNOY5uC
9zEgy3h1Dxsshegpdtqysi/npHDMApcU11llGklTxDA8xcNE0vyFKTeqpU1UcYSK
se5RAsAmEpg7H8riE/qWSos1HAzovt9TK8Oa2lbMIZGuW0NVT4SkivtPOWHTjeyg
osmEBaeHjCIAd6kryA1nzrZ6weeb4Fo7YlYOJiC0XsTarOiBqK8Ljb3hjv6dnecG
gXAU2xRe/yElUZF2x4W2oqUHvuCzqFhNkw7xCoNxoKxdNbgfAPq50JcsOrs9bVnr
iRO9ZyADH2e1l+P+A5fzn+Ug0wL+94Q6uMnXHmYidZ/U9+gHasJvNW8Sg1YCFl4Z
edE2K99fv2j2OMyk9TA8AxF0eC3WTfcd0YajdhRLd4LYg51+xRSZFyf9sykPozB+
KgCiQgMMV0vP7/VYxSpRqFuh93tThN7k7VL+kb4lZt4Z916BCt+iJULNonAL/Cbx
JyOC96dOxw4NUiFcjtjlMdq69vxNhUQ52664Og056SAv2y4IrjSA/zis+XaLmzlX
JKdIo3/bXdFZphd6TjFHA9RTlubCgrXOq3Ut61OXgy6ub8L4I3c96+P31vZRiWEl
SRyctzRPU0Xk7M1X7ht9jiahLe8seU2RBPjISuJ23eOWeF9xUnPib09w6/AZdGhQ
ngDP8886PPStr/LxIWFmy+MlxbYapIF83pqO3r7VTC3/ZNJjPor0ki0FtExqZVji
Zj5nf3PMMTh5qd/evIPBrbPCqvKNSmPzU9kw+hqJqgP9KTOolCQZXqx+8hbG1S5B
zbuKJvw9dZDUYMMzYceoHcuZLxEZOlQ6NuuiAJ79L98kFGJX5BFdQTtIX3g/gPyZ
CCdj1ZzEYKnLWCejST4yk5QbR3uhXSsBgUOhYGYJ9oVhbyVPyDDF6ChO1aiG4SVq
8KKZ7x/3NMTcAyfmi3yWxacUPy50bYHbPdjTlO0sg7i/cLAcl5b+HIXB49ruKjNp
MVT3EiDnciryJUSGP1eQ8l1weQjSorLCzravrSY4UmcNgQMp4dlwc98Q6cKXHj2/
DN06IJofN/1gGPFFviOZA6Grg3lxqVzl6e+xTV7ngqymt1h4WNduv6RsNsnIhssJ
hIVISFOpG1SEcIgVq8oO1AjmP+JHeEfdAtYgXHe5tJKyiC48gfJlIrPPYJ7te2yZ
nsGtTSbZEjKLa2CGmV0rc7WjAOgScY0QZ3AvVcUJMtagUTmAoBQ7D+9rYc0M9J7s
yu82EblJ5zUZ991hKhI9Gq6XJ3VTgpNH3g03fGt0CRtHwNkhop2uZl+4+0IRVZ+r
8puIgNWylYTwelKTGU/x8/I3P73XUp/OBQhdjKqxwPfzcWbdv5AEAJmSb9G6h31w
VlfDYdybTCiVJei82KxbzAgiqAKIB+ERj5BDLP5KtIQp3ZIled/gID5i08BwniDS
uFxHb3ABwa+4ZGi7DqVXTpiFgBS/L37oh8B66C9pRfgl/pno/CJXrGRp/GS5C94/
6veQB8G/fNvvPc7roap4fQXNrX0H1wViWFJcArDi/d6YsmAzT1KE7k12FmuBA3br
taQftFwF68yl243rbI/CfqP5PC4TWvmi08G/KT6FxngUktDcbLpeg3mwiZCQDS1X
rhTEoVMDhRyNUQDV7TTEC3MDrSEDYpAdPUwTGHUhnDN5ORaEGqtEK2PNzwgNm+9w
P5/cSs8sLLFTDHCq4cJaOteZ3EPb5wXfzdlPH/Ol8x3A9plh8RVfHQUFSTvl2whB
bePW3y4I4LvrVyUvK0Fsqa4qpN/GtvdhEI6/2XMzLBMAQxGC04/tRZZ0DWjLYBH2
CmEUckW1VwieQvjI9BqrwiIv7xrwynb43RHNkvh7mds/jJzosy2cVnLuA6fIxmGo
qv2VhwhVb3Y3r1eynBLJ+CImrN2twzgxpzJhPMaynVLyp3OY1pEysXP2WAmwxKqc
C8iWbik33iIFCpSJ/NhJQ0RpRJ7SgOksZWqxPWRD/mJvR4fCZP1cEQEfx0DyEIyH
yMxyMoWoNCZ+LnW4bSAhSXOx79Inc48ibfOeLiWWNezBGCe1xdVVj43wNtt1mdLO
azGugkQzxUuK4jeJ1/LsHqOsX77s4nsfKXH8mmG5l3x+NNiV8fox2jc7Dh4+mamQ
x4TUIrLEnaaPljaZgVbQ9H7Ds/FRC3VU91TVcw8C6OHB6lgQaD4JezONHJy5LaZD
aHCf6E8AqiOh9kFqZUSTvrO3AAinsphJeRwnb9ag3QvmzobypW4FT6oWyP0boFJ5
dpACSmVCZGa3vhs+r2LYwLuxaBygkea7BjtIKbZlmowVrwH9zCBZpYXy1blndWuQ
Gwy6FFYe+hofMwvz5xLKTsP21GhHNVCZr0MIJooM6eUmPP/DiBbGKrwLpZF3/oda
COBkut6KQn4hjzxMtmAz9MZtryAjoqpOpItfYkw30W3yFodXC8ZAI+2KvpOSnvON
MKKZJQnIsGoGT1Jwv+C0wNpm3HNBDheZu3zDQLiJ/pwBDReA2mnzqjZ56ie1TI/K
74c4E3Ec9knzbptqTF3i9sonvhyCgIfj1Ku0gTffp8QZydOGmAU+tXWcjfvoipqc
EX0DqbENPzfumBeGoe9j+RlAYqHjc+iAqr/sQmPb8ZMkvenyqnysPZFUeZffKUSJ
71OQkDO3V2LoucIKGZHidV3Irifn/LBjXiaiJqeQ66JqUIj2e9FO4x8jxgJilMHB
hX6PlG1hLkEDrsqzkXmugvV0XDBMxkqPsdKGjwuuf2cNKivMxY7HxfyQkpbLWRg9
d7LGmaTE0wVTAFjKfvXsheZJG9mNLs6T7Geq0l++rbFdLVq40DFHS3MzaFb6wzy3
7x892XGG0pwUgB9zLhl0L40DXgpSjGDUwqK2rQGBX6hWWv8wiNsFPt9VI+BRPbw4
Qn73eSThiZSbwhCOcgYdfGfpylZGsJ/Ne8Rm+6Sn7omYZyYwkISY21tALtY+A/bI
6pYvof2IzCOukat5OOsO98l+s5+DjMxjDCyUmmpjnPYnqQuADakiqBZ5NELSSwLv
9S56hFuIi0DGYuSIasczYB6d+kM7cVEr17le1LvKPmyjEwmKheOaRvAODq5RNrne
77dTx8iH5ZUaS9HBzSp1fK6TOfczWrukh9W/pho0hW1jsIIL+Yc0BbxQhmHmx2+A
9Kz3vo+ztWijbEMMqIwfn/xXiYkw8ablsEszZlkIISxMd7YVU6lDNEA40xVdvoLI
nNSgcaKlI0RGmsZPPA/2iz/U0WI2iPpA6pP/WNetP+DHOe+IZfVdFxWIkkaylbIQ
vvDH1kPN/gM27H0zO/5wI2aAXSA1PqD2G3btTP/cmu9HSCtbaxMhnMI2eVMKf5Vs
mlNRcq1D6lDQKUTVCIiBfWbhpPld0M7IyTh6lO5Xp9KEOhexKgrVjnGTb0Xuu9tW
CUjDwTFLK3BSLPv4YDjy+Jf/m1vc6fFOVOlTXm6UiTUyvnpIklEc7g31RBiPaVB0
Lwr+305PmGu4ZazE+oKIZBfN59zNG612RcPlhKlFyWebjQvgbNtiUye6IuqKH5fV
I4KeiZIgHCQysH1HnglbmNismjZSrh55SNej52q663oa2q5wAAYFbterVqq0styf
PnPJxXGuTqleLpF9xDJtbFZIp3pXKUjgTAdrDLOGefg1Owxx/wUH4qcdxhtSo2LH
r920K7a+7DgBTaP5gsfwEiV0ikjJ0gC5iULqwvjzTlPIAVZx/TTkbx4QqRYT+lYH
txg/MONOe2xQyW2B5NiN+CPay8ZD56WKlhDKenrjT8fWbk2l7A6U4sRN02wUsG9k
/B/HxSpcWVR2kwNNOoVHp3REqOFxedJW7WX2HsvxUo+xt8/h39jtcSUPwieLZHu+
I0bMBYzLUuAP6aBW4Odxtq3MpP2RVsMI7veldL66fzgb1dy7fO9hWHBxlKm76l6B
n1YDNuvGh/VF7VEatQc/Yy7UFGw5eyNr5C7XfH8jNI8VgrU3pzkvNsx4koZyCfMo
hj+3cSVZ+k6Pc/R0POpx/mRVbGp9ez+O36yetXDlf8/Va33CcHwZrjbZOfi3uJiY
/3JoF2LUfXQEfjh+QbcS9VGQMubk/FGKL8ibtzfoFLLNwqIKvpDagfALCmxvYeoS
vQ0HV3qnA3/v21gtme+oXSxwo/EbuksvNxAesaMfqO83QLAIohvYz9hsGgVRo3K8
lVHH7E3p/jnJc9et9qadXWHHaKjGcLyluipdm/zDvlbMyQf+VOqIanemfHffAZnN
ZgKyElTz/5B+OQ02PfUGqUcp5IyrJtACY/nnzTMZMYIYasgXhqeY0rrI9LBWyV4/
m3sZG8bUwubErM07MHl/d2ewmSXFmj6J6Jfl5e5ZqiaR+HXO36mCiUrU+pPDnjkJ
lVjg4CFdsjp2bZEmkr6PqCDhYFU6XqC48Q7ergRgf0z5BMRiPe+Y10wsbyoikl1g
yWSsUwNz/IJv4BIviueFmLSY443Ta97cYfgpv5PApAnQATG6PeCR+H5PQ2A0SM4/
5oWIPueCZ/6J/GyUrfV3JvMIqZk5nCjkQNJWfczCFUU+gNkCTtntc2dtUASvMsRz
EFB5Z/BQ1zOTktyFn97V7er9xl2zXjX36GVe9vzVnxWloaicI9ROScnqgmaczwt8
AIgp3c31oKS5tvFzlk+7DDmFZbc21jQ0mtFXUWcsDNqmY85fLc2/QpozPDcN/4Ch
V0rXWhOiTd83YEg7DYjM/nCWcCOme7sUgj7E3GML02JHZMziJeR59jnO1LUYHvEt
bh72X4xXwcv4Df0LRQcmKL0oLSmDjh8vbHI+F9EDRiccIfiCht7edKtvsIngiqFy
MKDTRlBnRhNB4watNC8brHHHgF+WzjiMyq2siMzjKCYHq0uqLUoPzabqfRMY2ult
UR9qmFgBV0kzunXLkQYoD3rk2XiUeAdZQneBA135lsYe1U1LdO4JD9f7F/DgJEn8
VWGIsdWfXX05dPKoNLcAZJS0xUKL2gB2dBD2XcMthI/itIDAPMAGLWhJ9i7BvnDy
zBSESzJUzXDWOfutZk0VmrdhzLDg/2f2VwuiE0tRQCvZlZvVIdOf+Ke7ZagS98fS
bKGG9ut7oXw/ypjhHyeQrivSRQG+iAo+ErpUgVQ9pWRpTyZQOaSZNuwldmvR2zpB
HwTGVbt+JHI25i4iOMabEKONuUybBgG5Kz4zgry9bkFdm7fHXG+K1r4o7XGs8qUH
wOt55DMp7fy1LrTUY9177MJUC7G3+4RYNvYHopMRgYwwR0hiJIcMaOJPp+jMqQRR
hpsP/bB4wbM5ozga5PjEwc7LQTneTa/qc95WxD/EquThAgMFrDZ9NJJEYExUaLUC
TSWqgtnBlzRWEb0YgZy4LprA45AN11c7ETT0T/BCCj7JA0KqP4ruPc2qsOQhWmAn
lCU67JQD7tcsaYSf+Y2WXoCkuTjoMUPjEh0ib35dr+Fro4aBGhi/3iRv4xlw518E
zWozziHxFW2cEoIerIe9ozDQ4Ypq/9RKiMyQfiyEzO3ZtckFJApaO376ePGQImFr
nd1m+FfMBxeVqskDkvJ38NUU24g64ETmTfx4ncJ/4d6eGhvLnovTaOEuKKCL0DaC
lYi/N2oPuXdpHXb3mw6tjC430aATa5uZ6x2ohbSmnkt/gWjBWCyfkTvLOWyMfI0H
a3jRTNI/uGFZkx3aXgdjUDV2NKjoqjDqa2wPaAXeDSIPQbseSi6qc7fzoO51iiCl
BwXZb2r+8sJeNTdFzzyENp/s2rrLOrx8pfCwSRXrpvWSncMh/6qZfx49UxsFm3+r
PQx0/yJBM6QtPY1M2hUvN6yfiOIoVI96EXnVZf9jW/DVn7VNt5ardClU/x6EBGSL
bPFEBX5VbxD0Y+0mXFwGseqhHrYXCuTyfVdMpItAuDQRxCtx1rjhNechxCYuRi8p
//Swbqp6+tnwHZSxuvyiIC9Ybi5jDm8l17z/xn6eF9GYs+sXD0H+RYjlnZkl4XQR
77N8QH4vkCthpb3vk5HkGWPkitj2LssPsrCZu6nwdUYTwSI3nhACUJ2z/vYZzaDa
Sy0mV3NYGniwKEXteA5xDdirTEQvbUpzy3FKhOxH6rjsVkixs1NdSvEhEJQ8Wz8/
fvh/qI/TBLlhYOzn4+4E03F+fqIgzEr863ueYfeHDt5gkSeI20tEtgE9bP4z9dfC
+OqW6s5RbOQ3dzLdcKpmFAvcdNoYO245DuNEKp8xKmLP6e1BXm88RHSxb1O3SbUt
iUxoQPmJXn+twXQsdgyg00kLfTPInXcvjMI/IcU4+v4IiZnn7mP71KRz3wQxtxQ1
3Iqy9VqQLK+FT73Z5dIgN+dbnSGW/fl3b2aJ4YMEU7sZBkXHQ297unX1KD/qVA3+
Q6uWK3NGxc6kvXq1+ZnhAtLGImavnBmS51zZdtlOvQ/B+44wSN3NM83MwBbXuNbE
tJvwb27dpd2ylxmpcbDWd+FOLYr13ef1Q95dyfvTxIBMjrerdMa/HUzYj57VM0kx
J2BoPSshP0Qm3Q9B7t67+3oQdULW7+azR5a0JkRwa2ao3hif+5iHdgeJ2nQWO3Ld
q+D9bFCODYo76sN9Q8PHXWDMCwhDOn0jPdu1bx7B67ECTwx/26T8p9/f0LlESml/
iARWmuVE4t4Pw5jUlBNiP4ocbKp4KyHZqy8jnhWtJQCYnVxIU+4IvY2Y5/8Fql3P
9pfGZI6N9ztm5IWn0UpCKchyd0QZpZZEez81sPK5t1zTbzqtY60miGMxf+7skrKI
30wHNSzVbBAaAu0rO15jLuPIkldYCb7NrCcBc6PrdYPpGn/MuPmgg+vH/BOR7wri
0BWzceCMlHjD81il2upL5TVyVpz5K2zwL7Pi+zEwX/46/D/3HjshRiLjJTXpM0oj
3Ugo4J7S7lBYhjhpBLD0L/blUcjuokbxHGNWhklqkOhWKKULIEHFues3M+AF6PIP
/ygqbUBkPIzxaHuSJfZJugKWP3kBCQRg5dEqL39Hu/nnQjXjXU6lEAqccO7GehHm
l0OspMaHaWbIZQVVWSm5xAG2kI4DJUMfiQtOk9C6SL7gRBsdvelhvNrW2vOW3x4s
Ed8t8dVyhZm5JY7GaXF4KegK+B6clTMP2fYcjAhVUdOiJCWIaVXZ7fLevaJuizZd
dFLijNxc7HnlU0psB5vWiVtjgqI9rV3PwDEB9x1mPn09E69gB/lx8Du2ApLWeOTK
3fB1I0aJpa6L1p/irS42LfXWkzbrdYCcy5v3oU5eTs0Rqsn5qGZbqvQo4KaV38XC
ih7i3NhP/TWxpTxWUqryORZubzsd0IULl7xiNVI2YdamSU5VphIiTuKCh+XowgIM
FKFUaM1Pj/cdfwNCcRWyhdWv4bRCjl02EVoK+cboNedy2oJND7PGW7lvevULF9pJ
hgyNOLqHxRuQzYO3NggsT8tbjzHL/zQCC/Z92J/5HITKDgXnz9u0ftZDtT3HeL4z
wrJ3BYYbIr/stPLublxMdqwdiSNB3LymGncTcXcCK2haY1d4Kf6O817DizRPJ6QY
deFlQkG1h7iU9WJYHN+mfYG6rJiBFhPjhIgSMfec3p6twu4Ha+d9S3SzmQTJWuFq
swDwWi5x/177rpkwTw0LEZX0BoIpR3mFQP7yU6cDBynNZTcYyHO0JyaRdk9vEJfE
IDRK7ph/mb/TVGbVykTzVOfa3PSCesqRd0sMlkuP+oRswtf3Sjeo3nzCtHSJBiGJ
xCGoZE1ovNymEWpzHf8smSR39p9Wohv/KeRZ+vAiUxcty2IOsHxg3W1bkaAmuMuu
0euJmkozKMHqyQ/INNviQG4SuCR3neWPb3/86sTJdF3pUbPpJ2TMmMGy1Z26Oe+Y
KhqK7Mf+9wno7BunvP6PqGELQ9rbVgu2DFrOQYtbd46zMSiV1qkXJd7jbWmaImZj
nFdD5K+c7jmssPdqipGFW+ceo+i9Xf7tdGB2Nw06N9g213zhPA++0TgIf1nwaKRq
kwYKKhKiD6YM3z58YRwEfG+/ZmVILwzmmnTtdlvarmcOBgXNtikZx44BoMjbkkAb
unouD9dBnRssvHL2RkHwxYbpfShXkiNW1ZDKgCyKaaC1CkSyhJQPr58cgAL7G7fr
0GpCbb+VlRKeYsBMNMeGaqL+izyL4YoVHcKFzVBV8m5FBXqPqZXUDik7zPgezkVt
iXrVW6H4EzColTkTd0iqF1M9CG2Z0C3vClHJsM1I6C2EdALZkFyqcYDd1HnwaNl3
GBnZwVx5IP3IyDMhghL0Oc4z1urjssVqEA9foytqvRTojK5huFMgfMqyzwE3+gAp
5W0VotQv6oEmtcFerDr76aJsTFcbqfT+XhNHc1qG5uRelONCrEPutjjDYvvJSCdo
6lhmoLIacw9e2kT2AMK80gd1DMnngC9Q9C1hWWD4dgLkFmF248V5vVaQMvQqURaD
4HWtBZfJ8u/Zuo2LaFP9Yt5FjQfMDBtz45nZ4ks1TlizKw8z5c7QpVLtiz7KyOdk
NCeNvUERwUFRrvq55pYSesm33U6SiFGu3f5N7GW6eEmfSwQQt/JDGDHoi7jT87bH
NtGeXLy5kyDMV8CucHf0pPGUWCvhjeYL7Ggho/NLISwGUOP8KXBP6PIU9rPxZb38
i7znTRY8uQnME6TfOlUv8vel5caWIQbpnevHR/Vkk7keWtpwKiimviC9Mffhg9uC
cpn4QF2VprNr0yggECtlrfv2l7McJTfGXxfZhutJaSqrdJSSuLTYkpKsWIOcCACw
WEQTHP+kXuC9U8WNwwJAlkyD1VfmFtlEH70smIjwz21u2WmJHV2WxwmmbpCDRekR
CC5/y14CP/nbGw3QKct6uZDj20kS+uEIiBzItw2FSfWnWlqrmXk+mGOaobMhOov9
k5+trl7uaTLYngPwJc6apo7bSPOJNfk6qG4kkH1MHLjqUoxv6/7yJVYAplBEIzZa
CWPDMIzt+GmM9K/ekka87/U0XUCPjl3jCbB3eNytJ/WmC9aBxR7bsB/RrEuFbjxu
vtMs0MghI6nbOAyxYg9fYyq6qFVkie0EawQsC9duxi+xmz2FLulsDf1+pDEl9P+l
ljGlbiJeFtSQ7WUqoCcaXEdIgqLMbQX0U+ARS8OjydRcZJENgamDwhvAZYhisCdU
4cW1l8wwFXTrPBRtVUdpi3rWeGXZviRp+mDzoVCfb2UGCTA7jIzBxdxzI2GzJKAY
+lR3W0RC33UBkpM7ySzBpBwSVQWMauahX9UK1nZhPtUp7uDsOd5KnBug2cLjSTHO
YtnFycCezzz/6jA3HO38djp5beT15G4GCEzxwXuFBSz55lygDiD9ZvqE8p4O/pXL
zYdStZktYW9ZnEDtv8lIRIozXYRhqEegnfQ0f4l3uDHRCqiLUcIHFRPPPfGpoNuZ
xpfwGNGS6d/jp5p4zq3B8kJCQeu9JRqLrTz+S7cI+W2SmYVwB4qCMPQOTzKmiIAy
g4aK0gIZ+YEMjtcQGFufBpZNZMVpWcuPggT2TrJGJECjQ5jk08IUBGIlSyHvHoEO
U2fMhazaFFk2OlcWYYajjs4pVWdFOi+dVkCUyi4Mov1ckPGPG/Wuk03tvCMQ7ViQ
WdRSD3aR7F0iqSL/6rQM/Mqf8/ZzdyZvEiHRXNPF7momCZZxVn7hGPFcMXAD8/3k
CbCdVbklIiuXrEqGFoFu5FT7jJDkgIpbIsUsccGgkVZvB9o7525H0M56m2ftOvT5
1QdX4tPkum7Vjna6y5640cJnE8vRcbwRGy61g96k260znPByNoRAfrtLDQcoFGbP
Oo9MYWfqHbx3OFySxoz3RMCEjcds8diSXJjmxWbs/irVu6I4zoVWS/lE+KWptyFu
OegzkEUG3Q0Xk/FJ0B7ENGc4Ea7hepbs/t0g9FHUHuUd8PXRUfKBL1j4LIJ8MHys
umxmodRueukhLreyObC7AKGoGrWwRZF3nAf4XCFl3cyeeGjU3VLE34wbip65MZdR
ypt+20XOKi9krWzhKFf9+L0sxej45hsVtLX53sfjUI/JvHYJJ3OA8X4F3o/bNQSv
3cRKLI5449DGRUFBWt/+2+ZA4HiFN2YXhrLXq4eXv1612YJp77XST5iGNdWJkv5h
503Mk5Er6qrx/Qc7fJNQPtr3+CqRSloc4lrnAArvb5r2a6YbWbRpQKkO3hQKbleR
jTZE1j5yPLE0ifS3IsTcu2H51q6vJx2u2wXS9buwgePxqj4aFoG3rN4/WWp8DZ1X
XR+7T9EaGIO+9JfzNLYwZ0jsO87JAjPuWmPI7HADEFWkMP1mfCjkhQ62SqkBNANN
rwlxGOkLxgNllvdc48xGQ6C7aBVnevT/aeJPjIlGHelfFaFIEu7xW5HzZqla0VfR
iPMelF8F+phAwmUReJp8ilxm0GaW0PPxPQ0bY8eY0j+4dy5cP1m5YK3F96Ua/3gv
NZxaicdPZfnrbO/NWyvVuLc4S2L2FlZqb+vgcVWXFv067C1sOlCbARaF3D5K+1yT
QO06oLgTZ4KAZGxpLpuquEkVpLxyxCtH3xQ1iZzrRvhl9mtNX166Gb7XDtAqhlIq
qxjiUGYUMIF5SZahbhW2LV3C/Y9jZQfLg+KsbNVDbML5+G27amHjuKLU3bzAbEVG
rt9iMbfQzO7Wc1XT6x5hPzmrZRMBn7bhete5nGwXM4lZ5715Lk5F11xhoFdCi1nC
PrgL0V7z7pfeafMbSgs5fWXGfippSbt7bOiaSIPEoarKCKyCe+TboCsWezOwpaLj
MGJa+ULp4QjB1wV4r9FOiswFWXD1O/1khNIAYsufVHAl/UdLfzsdMLj9rjqg7xrE
87UHPQ96bw3x5esvBecpMGBvIKN/fjU+72LDxurih5MztTib99d8q4hNrLEGUFt6
loV9NeKfsQEj1PuUxcH0dp6I6LyYPYPrDx2NPcEcbT/RHrW2fEfsRILuGo029rUv
46w8VKAGpRH2AFEDBX8bVWGhSclNyE6TBVUu7O3Ia/wwe1r2hk02tlZDcEn1RFBW
5zv3T5ZS0Qd/o+/FVFmxAo+jCRQf78c2gKPz8kBGDCi2vpAH6wotfllqA8MiGi0m
rz7JZDEp41b002rSZCA8zEGs4uL17qAahVLH5Rx1YDCZAsIJ6F13aNZHAub8wSYp
HADvlq8VVr20V1FTQCA2ZDY1zc3gLE4kO/s2r8Bz+HxPTZDN5/agx3WtYzmoJQIZ
yLdi6JQrlHjz8evpI3AZfY5IVkhu6qUoibqe5CkHYqUELBJ8HD3m3TBUhwNVISjt
QeuSpdl59aRuCdlDUtHaif7bhIHPfeivh7Nf9NxIkJWC9rEcnU0tGmqDi8TtrJK5
sO0xOEe+aPlCWi6HG6UW9uaii+kTItYnWDsFMm1vWLUgQZ3N9gE9EzfsHtYSI8fq
QSn/K8wkezkvBTKcnNHXepbV7tFMP1PeVndsjyZAj4RmCFL+3uPDA/QahbY/NIXG
YuA48C4LtlcLLWIZUj4EizBOiSsboa0TW4eO+LGPGvvNm5qrQ5BzmcunGyr3MnsR
LIk1TulpAJoSJ1gvbsxZnEXZMBw/qmxTGKSlJ1C8Gm79shbWMNIqAnV3XOziyk6j
d/IOfSpYr79MPc2taac+9Gg/uEl99C3PdGtM29ziRV7UMiav0L36Ckd9emOAzTsK
CDiEQ4qaSwN28lTPew1NVLooSdXJleNjIueaN7WM9cs9NobhTjtQDJUglwFXNBVz
b6Y8NIexmrmEcJc+UqyMtutB9tLz7aAEWO42aVpDAlmyhS5fqaMYkarKoA7ZycKN
QBa2SXKoDJ98iwvS2n7EPlFiCKdrmbn8LWTjqA/eRG4KmXNIY4OmYNLeSHbKk9TO
Wsu/PTmiq+EmCT4/mXbABE3sJ7ohW3FUKQJPk7VuZElv7nG1ZVEYDWDUex02HFdU
E1LDJ240aOmiQeATLSZ+wFxR6zwnmBsIZE8gmLEyrfeOxO+YUkJqqDYDPe0XbVez
TQsszkDsfM2l7ldNmu+VdtzYU4V0LW9G2i0tlS0Totb/YbHDLNFvmf37impz19Hk
jFvhFXHgZphlJVPEkf0MYV52BoBMZ+Pv/3L0AUazyJur5jIkJ9PJXdPaorsI0XJf
k5mHZj5jp6I0lFgwba0RPUIhyaIi/8un2a1ff+Gxt+guYddJYhXMDH15a8j+Miup
uJ6p39DUnYiLtLyIIHC6yeM/myfEo6E1cUD2TveD0Zd5PbwIdum2SK0yKUp9ISPw
2buAjOshikfIEuzmiatvri0KidYT/9kdrsO7bUPyHDWhFAv8UyNpx8El/X5d/ksY
ixFyGW+i+WxYZOfOsgR8lXKS+bapLqsV068GAenGauuzuv72WATFtRExJawFhhxc
aHrFkqRNEmkvVjHgcYZuJ1Tu3ag96W31KKf6nsLpn/PoIzVNx/N2bX4gv/zTWrDq
45yUSH8+PrEJoNmrKPSZvyc4uruul+5X16JQ1o0VtcLPbiC2SXILNfCCdzGBfk1z
WSvPbxI2Np9PnfpKIPQGKYpBo3wuUXwaRa11A3hlWzdypnmK74eC0mfrSqYZJLMV
6y/0Z9xcOlSpdd5U2CcW1SR/VFOtpyiTy6FoLZ8kTPKVw4Ap39q96MJ4v3vlbC8W
LsXScxyqFYgxyF/LPdMPEaaScW51tijLK6gNh6FtqiIQ8ThiGDE0SN55z9kcWD6M
Zq1T0F0/lLhrG/97e+JTkk2Tw9jPlPK0qQv68mQfgSI4cW2pXtMh9BipkO+2Zi6g
ydyZ3OayKoa4XozlqL407rzV2fan6eOSaWOSu38XpNJ8E99quzyXiYyvW8nu41cZ
EZs5qgKvd6fTcI7DV17zsmLts2oFphoxbpsuhsgmaOCQrnmGjSjTmEVZTF5ZHHKx
aUY7Ee7LKVeVN9zFcNBoWjyVRgDqVZg7d2a1B2bPz0ndUk3hxelLIoE5SETEE55V
hsTewah18LpQqbTA+ROscgOJA3ijKBaexPq8BXv5QhTo7dSnEH6ysk44coOaN6NN
Er04uHeFUO6eqnsSIGdGYZrngfhImohLcktx9nFdkh0Aq/XVXOCP4HxRGeGZmq9c
POOqT1uzdwic7Xh85A/XYuzIuhp0O64eBkedFgx0qSAvuj0YiPiX/hhlrXAozBap
qiu6RpWxL03rezUp5/B8pCA+wwdemkbNRLfc70zZitGX5haKtQkgl8Ek+7EHkizb
9IVDr+hbXDj3SSFT5zUQ/oMgxKmc0ri+5hScZLHenbPcIcyM/YbvnwEuQw75yTj2
O0et7VmtkeCxeabj+DMiPnVIOF8XQDSuAdmCNvii+Rr3woqZpX/UzYoS01rpW7yR
GvJBusuzJXvobatalrWUr83732goq75Ys0sFmhRLBOZ2CUV+HR/og6HEzG0HKaCP
DwHmaL5sB7SMbJMTfYqmwYbmB8pgSQGB2nUyFi+DT65RNVPn10lAznl0ULihshTW
2djJ+hGyspQ7edECgwNhsDooKNDP0BrEqdof2ZVzL0yH2Lb1Nxi7ueJTaijFdR6B
rCga+drxc+VFmzwADDy9fp+HKf9PEe3QxLU1laA/TsK2z3Vj5WMBxCkRKRpkpkPG
gUSFWcHwRIKyhKolu01ZywiJ/yGVCTHWdQ783THFaJ6BMDh9Bi2FyYSjbbn3dtqP
seAdl9zSj1PQS7+UpZfLJfT4IkvgSbrYxmSvQfSPzLREvRIUgqkW2lXKyeTz4lfs
U8ywgYrCHcFKUPj+Ckn/2hXeDHAX4p99thIqnTmNzZne8rJ8od6Ux7K6ahtSXtTq
Er4noEO/SQKXcz75a/stOVf5n5PAwzN/9s7HDb0NeMzbtXMESKD1HOK6KYQIk0ny
XwzGKrU6hKhtI3VSZVt9aeUL25PSyyI1kUoIsKbTtGTrHkvQPyUOnRV2jhO17mGH
tgdMmohOyWEj5hSh5XPWAhzG139hKYjZNnVPr6wu4U55CYzxghNsIcZ9BL7R/SEc
Gore9fj8NE0+zpt4+I14p/a3wwW71JuQDrg9O09i8oFiagDIGt2vHGmzLnPtuggL
tQO0iQbxsiH/3B3YNSP6PSYwIvzCbhgeb/eSLF7TUS8LsshzSGkbE8viM6nrn0uF
LkRKY0p4ZBiLWW46ubDzihBiHheABeE7DzutWNR2BTZ1NzozFW5bciv86Bp03O2o
LKizlDLKfrO8NJte5x5SQc2flhNf5e80VrH1G5DNDHV9JpvWhic/aRor9Habp4Qi
XXJH4nMtvYW4oLLKh2rJlCQ2hUlq7UXdxmqglRM+Yq4eIpoekgz4u+77gFmR7N6u
Ihs5GqXOw6aobZQbRIjlyeJO3In4MR83errL7v+1M+T6AdG7Usq6I7dIqdIVFY6G
SZbagKa7s+b6dIs4B6J/4t6UOruq2bBTR8ZdhhQTE+wA39ebHYelELPwjzI8xf0j
n2ziwMIJeGurRb0+5e1qSSUcTv27z4ug+NvPWl45tvObGh2YbIhNOOdbxb5r5RFu
JyJlk3im6yAMbXX+Pg2BsyT5jso/WuPjZJGhhvg7gkmVqVB9zAv5Eepf/tCbHV4t
YA6NeLrhKRSrJQNXvqV2gQDbEe+F8EvPWf1cdE1dh/+jjHtQ88ZOztFU6pl1r1o2
Nj31QdAgA2722t8d8lPAPeGkZO1SamEWM2VLpyKy4ZkBUv8PVbePYA6HCaUIxa/O
wXtNqQNRpGY6UvfKwgyadC8/DaggYPSInZ+G86S5Cw4Jna65N+xihhed+nE445Ox
FKAoN1jCiyCPRYgoxxGs2FgV+PGIYtcC5xVNc2WWzajU+dYt+bv1geZvaLJnZvUK
qLvEabXODxTO8m5kZiYkSo8R1BD8tcUSyz7+rjw54PEcbsFclSkbYj4Zz/GAFdcS
t1ZyiTrLr4EMooFe3loJUzPgdlCtxJULQ5yZCj5Fr0a8bQMmy9Vw6q8Mfcd70//w
tbL2PGmR8GJ1Ud6KokVcaUrr8WD6++FO1xGOx4uCl2GOmOOHyQ8INwOJKrbGaapW
WdgVjTqOOZKO6D6qMm8/dxfIMLJdht7kz4wSqDGtWCukxsDTpAm+uZKDoBh84HWf
ykBVVB9gqoyW4D4FM+JWKCbDOSdx2liVwRFf2svIsHPfwX6RceVztTG6CmAsHhUf
oxKs7IRJLlj87FYjGYOmOOSKpe+1U+iRn5gbWZ5bxXoTrufM/lVhjCXWPFqa5Ezz
1Q5Z6GwPQ1wlVVGkujjjdIXWWwg8xdI7Gnzb/PcAA8HFTpGOzLR2cOws3p6VZJP9
uY4FEdQls1z6nT4n4tXeiD2670NWs5oCVv3eFB5EDO4xdwJy+gpigkp7zc3Pb2X5
4u+BWtBtvsI5oZ/o+TuOCVQAe08/rvxH+O8BYbiqNntUL2aVoJBk2nN/++sDA3w3
pvFYoIbI/TNpTvGnuvii4rE3N8294zrpXpOqCQdtpao5cj2KCHmF2R9BcprDn8NY
JsG8Z01b+R1oSaF7fXUKucW/Ky59LfppL4dYHrX281BSEa7ozkqdD/l6ipB8P1AE
UErfWsEU1uslC35Ym8CqtInEq6x7v1IvJgm1G07UgtsxzEZKgw36JihR+yHADTtY
mc7czzTMwP1yQ05DsCDhHVDZuyJdU3dJ3rSFONAAls1siFRfD+tE2tstfISY1Cet
s//xeUlcyawcOx8gKDvdmoV24cnvL+Ei0vzCPVOiXc/sTpyGodUas/XvStBBoxvQ
w371iMFhDwXpA+TkEvCpWS27+PzAOmuI3U+3RYaVt5yO19M6dJXzBjtv6pkqDjf2
TI6MazfS+e7/UDxLA3bXUF+OUEpCSjDvZFKnvRCFdaBtCMWav5CxVf4/2AIkz9Az
uszShkMs9R1RM09fuDO20iwjgwF/1YOR8g1u8h8aW3qt3liRLiwSvxSByvzf70HL
jJIaHTymc8EUVxitNfapPaeexWeccxQcM+jGqBgKf3ISbdR93HP9EcCACAGPBc0n
0P2AS1uV/9z5VqjQdawmXGhXR2PyBdimRZw6rZjie1nvZ0n6z8Syi//NBYBA8V7F
7d99BJcEuV3N9bUfUaSPIZZvXp4WXfvAQzO7HBO9vDD3RfoyWAy4shBcqxXucI68
XPjL3zp56RpvquElyF6/7oYu+76XZ5oRhOQ4HkkhrvuuJ+sTpD1ullXsG80QVQ6W
cYJnhwVhohRwU8lBmZcm3nbVMtqqM5fNs3vve+iPM6OvNNUcXzON2vUCSGk7XE+i
xECUatiYeqH3KzT8xvmtYTz5i480KL4YEL+ZFMREVnTg89WKuMpG8tT6dSKde/50
ZmUuLB5Pf+bo4dMKpfEfs+224sddNy6trBjtI9Aox0XvZYPq6+zBGB5+lI9AYv2Z
/brqkYzo5ibAT7nCvtWLTTneNa+KE3bA8SXTGyAkI8FailDHyHfz3gmkD2N4Sm3l
c0s5TX391x4Eg/Xabk8y/hRXoJ9l6YxlOnwPoq2wffagS5RZg3t+i1+fIF4L1EgH
TF3VrhxFUfa5f5yQcnTXBOgN81xLYce/9f4BcU1UoQ4qXuGP0A4NpuNZAM5yj/2q
q2Yfgc8UEhZiuJWuRmNexqnG3KQZGRrISKjPAOAoMtM2c/vvE6zKlg/k/23sT3kV
Lwv2li8zeHm+KrSQWUXHiPgbyJEUn5pwUWKnoEx/Q2+sFj79zpu04Em9JNgv42Zu
6Ek+fEFbB/by2bAwovDn6ZPlySHic2YpynMbAp/F4uVE+W2xTq/ar2uz9vR7qtEQ
GdcwdmvO1KfarQ2w6CO88zvJA8hQiRs5Dm6Q19rccgfBDEguFsH8f+DShKtQMOVV
eEC2/Bw0YK9bDanyVL77xlSNQuWqduNAC00R4h7flKgAIkF4MEmjBR6dHUJF8Njl
skpZ37RAlaVWHT66HuvgpFrJlcLC+HMXtcQEnySrEXqcApKtHe/GtlJpXPi3YV7l
F18Laz9NNGHEZKtrj7oQnb+v8mvwtb8jY9F/cRyWa6vB3mmwldAwG+FZJzYPuCvj
doKNX1cDSdmuyERyJH0mILKYnN2K30oTCVFg5AMTnTG22bqSprF1e9mXr6Pdl2dJ
07kVKIgv6lEDyA+Dw96Rv8HIKh+JKrWoA50cwT3LO2u3+Ms1ioqEfH3TSfAp/oUP
c6MaibjtPFV6RGlDGCEzRSDk/zk3RaeW4pMNTsAm7e0g+/PO/ONAmegVSjtvINOF
EhcTi75T6cLg5wRKOJ5zLZR0vWwwCvg8Waj+BW/Xj9dQPX7G+4nfZHs2AVV2wA0R
NNQ5ME/s0eZSXYtM91EPvWm286VDzD+vMqFU1qBhw0H0XFAe6t5xzjwYOD8igSfS
VXTt7fKfH0mNz5d5LD/NvhJURMaj69GxhHpRWBhkl/V8PWnjxMSyZe/TPmx27V6n
1V8FN5wHTP++XO0A6Ekg5n/9sCIPkwEh3VmB1Gw6wZrCjKCNEsU4xTMPpVmyotWv
srtA3AutJG1f1qfpKKs1neI5IRa3YfbrQeBu2iXpM5yHisJ4popv13pA1bVv5M8i
rN+K8x/SbMhOa5lH7qfCJY79yHuv/5cgdsOT91GbdRx81zvtEAMbgySyBMCC85qu
KPqUXV+NF7LCR9sXlU1+YiNsilUzCvoHa51mNg45mAVu5rFCbC7kciL0s0+yDtaV
YqHg9qkMrMwVqHjgj70PXob154jQ05N1gH8wtugkl7/IatwDWbFQhHIMq/GQ2q0E
gObWbmGWC9sGP4/dO8rErbT9BoVq6lo+pWr8vzg5lweJqFhUrBUPa3UInk83R4On
SHeFvoRYQr/75ViUJsPIWSZ2DxQVaGTeUwwVu88VE4Iq5Uv2HwMeKkVRTtrSMwt4
gpm444PTSUgcDwLE72LPUgIlbuucsQCuSgF1VuUioHK/rJp++ikm9Osl79RONym8
OxlkrElh4arihCYpZRBzKT2G4qAGON4CxFPDHz2U45bw70pRaef8trmuugHH7uUX
gFfX21H+RO3k2Nuffp4Bf2mFCcT9qEKIEu2NlNZiRLZnzJ3FjPKabNTFhJZZ3Ua5
4OKOLUPLA1g8dSnDPJf2CAPZXG6/hSMLyNOxGNhSSKkDXzv0vkNMsvrSCfIjQ0RE
8qFm8XvNotMjnoOL3Lvwe5PCYVEvBY0sWJ3saUQDKD3w3Xpx3vX3S8005iSg/OHu
lT1ppKFFATawL83VoqurOVhafvfxiyo8s5EPVIRo/0dz6ZuDrLJTB7CyrRMtDSNp
xee2aZDSR31VzUM6nteQn733CrJA/mJjNXS2OeCWNWFNVoAgIb/4gL6yveGo1axi
0RgzG47op7w4dzpwYCwqJfv4/gVgmZYKb+pHAmnphdF17crMnnMUqgjHVQkCx2Fk
yQ/Q4tu469UP1nvxmf6XWhSqvljydjJlLHLxVQn5cgTUpnxJHWSxz3zLly4EvNHK
ddxMUQaG/ISH8YiOqb03UkE9j/AKFrhjrs1kLCzLQJT4PbA+gbjG0kWoLLq3IL7w
BctVEXNyatQ6f5b4xl9Lp4mWoK77exq7+JYhpYRcDTfSJJwJnYJ4qdD41jwttG8f
6ZKvAO3C7KaVNH3UCpnv6c9qooBrUWTE7AuAn5kuyCmDfyHHf+fubuIWzIL3Z/hG
s8N8rxKls9cxGQHxcF0Z1DE5c0PJq1jstXFkn2vDQNjPoFJSMHgL33jPj/pfySEj
oAgHnJxhJebUPx8W6ruphSlQQ84G5Cujk5RWpFfyJgHqGSqIva/a4rdQP68eJqOM
R0yuwoZ/XFB/W+o39zHFJb8eR5IjFe/bnMSvTpRkZBXyMml6tAVp9IcqXj467hi4
Dp084+vsLHNQmb4ZP78/aoDqveW9X8sLzGd7FZ/VoNw+x1yc7E3HVJJZB1w1KMVI
gwbRTJpahz/zNCJtwdRWWDC75e/qL6Ok3XmPG7VNNb2WcOWyGK1EiqcQZaJi5aH0
H2gm/Kr0yo7l6ITMvKo/5Gt/a1hPNK1uuFXjroBFnCDAjv0/SJ19Ogu3U1R/gqcg
oBBX0fgFFrDhIFk8t6zKo8FM0kfdJmNsIQTvMsdh9XMH2qqgZ6Jm0Xi0QG8Y8kx+
CKRqboUovntwuh0IlcAL9rIi+hHIcNRqG+8km3ZjDoylxRz5UESc91moTy3xrRoa
2kTRiMZl2sMcOsnB4LnLHFXzk09j16MmUMXrMDxg25Qwe9Q64CsDor2AZriKlSkq
ftl1a0TKewBo6i+6bCzrSLLAM+yUjhhVEoVA/u1lyszPz1Ra3R1OPMBhdLke3fj0
A37OHbKQK/9KYCQteUqHNACOB4rWsOqi98HDOCAZJY1QhGLCcgNF43OnWMatZdla
gnwWf59Xb7rWBJfV1y4BKgMx5CjbwPOI5mWmWzakZcl1Wmjpqgks22VrbLNuo5ck
RCKAQ7OyYWgvt5f6vHHCxI/8/2u5BSGLDs7m4bthmCm+MfFRuz1c2FHz2YbsiZcu
OFTyF53Bq9MZA8fWFHBpr0TcJMVf2oQJ9+dLtTFsVV5B4YDg20djcekpHNNGgZct
SyQENU3e0z2FdHCT4sq8uunisi8/yZsnK+0jhhCujGLURS2/0bIus32/IPrdVnRD
5TF2lf49t5RGZDRV4SlNIsn3GmAbw69QWcI+D3g/nO2OtVmzuPpzslM1zrljlCY0
F4GQwm33EyjtXgbeXpFtkaYZ29kVbPgh8FC1G7Bn76z+JNcHEVlXGHG/+PDp5YUZ
g3XTN39i6HfmWRL9V8/86819DzBDcY9ZKeOYvehKz2hhWscxny5nTs57CImlzoYG
/2nKH3C0iXO4rP4WE6pd5Jlhtfry+5wTSbRuwPgtx1QrK8aWwPMfiKtSDPZvn2zK
kE+5sJTz1zFnVt4s6dIbkVSPrM2WEtcs/hFImud0WIkZnBhdrA7QABpw/7JEIM0G
xGKXb32dEZbl7WBv5Np1GFOakeRZ1oLo8dJ6P4R885A4F3S3FzkFU7RvSRCeuJOf
8cv2zRDkpC/VYryBiOJfP6cOCYXSDiLm+s4pY1Ofv33e29Hwk1AUzgldUgCQexX5
kkdjQesetmrnIDveDjV0ej9MDBiKaQR9fPdxJyK4Goq1tpebrSY29qCvU9RZyRTG
84gydBSJZ9J1UVbGaNieKcUKFcjP2b/u/dzWGYeLsrZZ+uv8a4UGt9xgPAVgGJxg
FMaqSCQ8cff3njVcO1B98EaESCM69RpD8rekDfCdUe/ueRaF+J5KtDEQWELIYJ7A
gfwh5XmK0I/P/S69+vGda8Z8DNr8uGkEq1wbJdtxZxhbJjcp2huGTMYtkXK7dXv+
aDA1ntLdU21DmFCd9hE5Q000OidsP9x2vLn6ADwmP0HqZM5hSj78OvVxXvXaI7hr
NHFFOJL5cawXJvTE/Ba7dL/Q5s7ecHIpqPRwZHcTj9KAy9Tzrm9zqgcOBdb0Rx7u
yP+9BMPfDBGRdOkdUcQpqvsLdjSb9/F6y0gE/DiZeWBPsufWpM85DbAmzMLsJ8o/
R3tr4ZRyQklkxCdtUbzSNk7QI7s+vBJmNFI1DVx7sVmT4BUDaDGvrBDQJ34LV21v
bl75n8THtRF4bunmq7KEDCqJkijcrMxU8TS9X0bmWut+6pIv5attt6t/SXeHFfps
iqiw0YmSA4kb+aLJRNrs660XLZfEJHquDL8R8LMPXoKoh1EN6nBGtxYjG6frA6ro
HgS9CqtmRtAakbPHepjww4IDPj6D9+nTBR/TSJg0bypj+ugogixaJXPvr8gAnF+y
hPBNOHliFO2IqLLo2FWFcIiz6prXK1moYQcPUkMZyg+q3/BYuDkRYZseedA/U4YM
f9Bgp9GU4CziQyTK2GAREEtIvAMfLjUv98KWZ10imdFqpWrkWWRixkxhY87t226P
3It9LRtqZj/KswWA5RtfdccTHvu1SZiLAK2KNEf+hs+v2bxhNkNESvGFNLzIfGKK
E7fjKn17A5Q+uoPgNV3u20gSMxvC/cJs3gM4A6TvUihDs0CDj3NL0cFVS/IscbYw
SHXSWpx8uoNvmDAs/YgZX7hjZXdd3WBXh0IhLdl2Pz1KUZGUFVwAKelyIHT9O6v8
5ojXricy80izA4TNknMOp60WOTU1lHkO9EWBWJu56/GBc3ABAPAN0JCOf7xvA4LD
9TqI2nfJrhodEwtL03980DgBHPZPBU9chBQ9yHy7ZGxlB1g09MPFyBOL9ALN1yOG
0BoMSJc48HXOnJSlN5L8uIPpXoAawBD5EoPcvTaCFmdza8e4KKnZfzvp96heJtA7
3s+ifsqSRADx+POHqOqkME9xenT3A5YksmCeMPhJ1W9yUyBW/nppETy48HMrMjDI
AZW97+sQWZ8N1c01RN/UuEhRO69lW34XYesaY+U/qiQ9jENNltSKLt7XnorK46Pw
PKbLda8RG3OnDr5cKAff+7aTOa7iV+FjOTRfK2km4APijI96RTLYEbizK1Zs4v4S
hIjiGVvdToz/xTnxtJKDXOWVeo4aOw/Fq5+wHvrkn9yzgeevTCBh7JDjUVg7sxj5
qEpXHc43ZyEkSOiMUaZmJRox3TNM7WqSQYCJwt3sScTva0zJm5spWzGzGEqhaCLX
7EOQfAlsuNFAdbIjnBV6HQfghDrGmxnMYmKBdq7JwWpCGcabqXeKLcGMfTIfLpYn
v4ayLCXi+x+kukLGGjMC3JjOmTj/RjVUxdgmItspBGqGCFabYdnKbhuH3D5bfUaP
rTAqx9fjN9py01aIRZHU0aGdAko1c4TMYrxOPiXtBukOz5L9vjgW9lKYGJSZ1v+u
v07L9qsIk2nrdTM+dBTMaEGOgqbtk367RE34J4lF/c2zBGqeTS5bzWtpO3a35Z01
2lmP7R1w9cXEShawS2qzTnKPokRlF4H4CCPUv7GaJFDOkZ1d8ZZXRQV/5eqSO40e
3EN5O0GPXayQGAT8614E8RYLtNOdGrXpUE1fbW8e92TnCwIpJ1MMMrT/r/2LHH4k
h/N/yHRel4y6uey0AsLedDhKCHvMnfbIjyiaYzCn/c7qqzvIkCyNFbHARSdIlKvt
/Xwdt10W+g6xb/1bXWfsknlg95jBAVTf6Tsf9Km1xvgmPPQlPmsoIU8MdAZE1+Uu
H9nD4BWpzGg3xtSdpN+smN1TYS5pFBHRFdlPSze+L2AYGfoqjiOP2S25abIIRLUz
trCF0Qr0I/GyzrnwTao3YAFcVkoYmvjmioyWtTcAiG2DrcMVCWo1csqgv3QmtZab
U04iK4NUER8Hfa4xyfG6sSeuo5b0psASiuQv7AHHAvTH5YHag1LpPV1t3N2g9wzD
9ujJ+mudAk2vhT5LEMRAk7t+HTmC2EO/ZZ08EWgYpCVEZA/JhjZD+2NzcZrGsxi9
DwIeeqMwbXsYDJju2Dr8Uou4SV9vT/dqxFrHIM/mOZ+XAffo9gj48g3B/romCXCw
usrCbDjBZN61zda07n3lEBMMcJaBpL1UH9HnkkbaHaCTc87/gxiYaUbtYqV0eXz6
43LUhcm1AxhlvIFyR58HIhxxtYEOlA41bMf6NHVFP/Nkfd9c1rmBxUqwed4y0H6/
ZKZimv1pwGk0rGerjfeYTdSxqdmJJPGiQLf8rS7e8l+S11NncQu1OEiIjUVCXIXp
Ym0/mqx3oihI0ujAOFcbgeaCRq7x1jfzrDFpG3+Rwq1645bGpx8wubdV1NZfdsK9
MTlQLggrC2rMt+vKH5GNrTVB+8Spe2bbMgyJbBVgLO+8gndgprBBRmlaGbN1E2LE
dqcKgGr2BEHIWETF0Pe50gHZ7iSJ8HfRwhtXrKozc5U9LQS03n7gx7I5XtnaIgY/
arLZVpzCq6QpHQRWXthpAF9SvywtiO2ubXqW/vpaOCGP+iwoaSukbkhmSuMblWI6
vjiuayU3+JE1l5EjMmOljsgweXIFDxngjECgBBUA38D6jAhYe25m1fk/pUsIVvlq
BARop3M9V23qrqfamZDy+CwWLCEdzu8trItcjFz44BrKsOJM/ghMUQ72/P2f/wyc
L2EWPV6apJmHgHb9it6DLGbX4FTh009BA4/B8+GrNnO+mACV2EHDDr5k/RG2hcjn
5uVpXMylJ8g0Euj1krSxgL26iLTcpszX1xMThzTnJq/1TljsrA0tojzjGnJp4272
APtrIm4qbpFmZu2ywEUWra/jQYv6cCm/a5a7QqdEIOn5OwfRTzkZoG70sBzZBkXn
dFjT0m+7RwGXux/5dy2gcxEfX6Z5/Rn61RE3qrc7Fxa1E4AHbeEPG7/p/8L+M2Jk
O2BESkkAEy5e19R+BDh+C/vIlBQgtnOcql81qBGfYJ0Khj8leuy/d+7Ee/PgX5UO
8NOflOF39bmQkrQ2tU34WJh+xx3CqEEEapCYSWUkMet5c6sYEZ6+PDjivO/Vcqd3
/QGp5StG3ASncLHgvsCqS6384Yxe2RcRFOcd3EPYoJb+NJThg9b0mPFgyXyp86tn
XsD/96EmUddBfP7UtkaEZyeglL9s7qLq5QedfpcLgQY1IaMPrBg1mQTu0dlo59m1
EIf4qo8HOKN/4qqIr9OjH3X7Gya0wdhEfyvXdpWMkjqEl2muDpOdkBlMl4+zoCRT
vLKliwMre+tTYYablU5mxvGJTaamJiKt7syhEviiobRiKP+DtkZMOmPiQz7Svp0d
+OXD9YtJL1lhW6SXnP8eGxafENKhss8HjFwHIzCuB3OfhMWbkZJn8QqTHvCU2bcu
5vTrR4EJ6tdU6zCZ0E+H8XOXPmA1cohdevwomHiW5ThtXubxF/n7UoGYP+hHCJ49
x38I1RUweOIy6ZBWManPUlNRIsjfELQCDf6eRvKXd5NRglRrI7PCW5srWXQvxtDO
64ezUn7cCbtCMr0KV+2wOLS04uUoXa9cHV5pW+NLDkROtev0r17yXzuABzi1DEIo
hAEdxNlGBKz64PFF30HRq8vIeUpTusgpvLBYXa86B4WwUDp7ly1xCLfcPpXLsmbO
Tv91L52GumFFvI4nzhFVqXu8exagS8LGdwyChgaSMdM7T9X7uPJJsg88AWrjIOMY
UoHo8blqkOha5buqKFu7i8rQ1+HkBbNYKpwuu+K3O/jIUGGjjGMPevRMgWVrnc0E
jUP9OlnpFMs3kwf9UbFY9WzUUWIUBTfw3DsUV/kpu8TGhiBxS8FaPN2/gkra2XdO
/UlOy4rgtNbic+Te1drp33MtAkzXN6o4n9Xb8e/RsFTaMIdOZuVUm+kOxijP3rT5
ncWH2Y+IKwwjk/AmPiuI03pnUqPGWJfkfZfS2Msza7HlY+CGzKR7MMDVmYf0zgi4
8xGGOcAwwiK+/25DGkczIXSAYsnyTsST7gH0QUU3UVweoOnY5UcB12LHv2uOY8rB
uKHCaE3Mlm/ERx1Nt3uWH9t2z0xk6idt74Yi9UW/GeDjoMpqHHYJPNrxKhIOk9Hb
lSSPtJxcn/W8Sd9cnQq4AiHscPLp2SbnHyCfHQD2k/xsqyl8+KSDzzhvyPcn1f4Z
bZdwI9Tu64sQLaIBsT0caXi3oYJIQHJhruj5S30juy/bSSWfrDPT0vjppAZr9y06
5DOu566mbj6LvRjk19ECp2+GDVAhwOT9FsWKdcOq5t1KtyyGoGTNzJwFFSygwNZe
fmtBuR78UJF8JkHiqGK5HKkhv55q3sfI+Xa6RjQefTGemo2FKmdCnKxtf5LZjpYX
PqyAe0vX196bi9fSwZeVuR5yZt/uxfEOUyq52YzxU+giTk/FyC+bbAL4A2lE5TLx
cfrlMcQYpp246GBmtlgZcA2oKyPdIGEkBWylSee8c1v61nqpjA1/qVadt2BVhOta
iydLfvdGpE0RhPs8hTL4fxt3W3R8kCWU8SRqqvV5RCWYypyc8WG/HpnO/fqK1lBK
Whx2OKUMBVDfKjDOZv7toA2RPYoTk0R1RW0KtXGuuKvPgAI94E/kCwFRDF5GV5cQ
58zHz5kawy079pmAEF09ENd83bC4fiOhRw+VWZGkykrtEjw22PFeVZThUhPU2igN
UbP4lxkAQYi0RjDIKabxraliGulhI96aPrZ5/XTJD+wjlHb8taOlqNX9EZT/xEyQ
S6QbZUoGvJjLDsthU439YIlVXV1NwI81QCM9R/jRcrMnoQfNX5tyNtye8DVNiX4p
CWBDSJcU3sKZa2kKuPCn36bNVIkkQPAOKu4hiWtpZ9MDrS5OS4AZaJ3Xg9WhHazE
hEift9rL5zh7WZzNZ4UxdMDK76vpqMA5YeUnmu7OUc9oyLTg8rvP8RNme/GO7kYs
gX1Uy2KYMpxRtiwV0JE6EJkLklrYIeZuWx0KZnAKoO7WVf3jAESgzoOJWKk+YCkS
WbF5bvEMvYimPCmrDSpv5/SYHAe/JqlSpwe1H1wttzr9Uf23x/4S211yGA6nS4HZ
gOyf85EYvvAMoau6eWG4xHGZO6SzLCvZ+oBMIfGdyvmzK6b2tctEBxqJuGS2XbWo
VOLJFsQWfP2XGsEVg7HFFN8t1fZz+XjdzsETKQgyhxpVCpzwT0D/N4XHmr1XhIz0
J5W05njGLoxPNjaNCk4ejtZTMmsPoK3gIhwPmblQah6rQNFb32vhugkbaJ9HzpkJ
Iw8UnKU/IYpfzXCXCVD1g3wcMcjM63KwXnB0brD8ZNFPG1/l3NJ1yh4KlKG3u7fr
MH3jcJxadc8W2FSmsj7yHbbib7fTclGRas5KRu97q27pNUJwhCNuVA9n3jFs+IiC
cZfEHFqfFi/E+/TAubhyUlyvUt6+zkdz1pN0jX/KLowNBDM6x30pqjZYz5N1SV9/
6JirTBNbHHokMY1FQud4by210KZiqXoYs1Ce1d2vmW+7cMLwokfEHbbuid9kmcMy
tr0dvhnrGkpraE36drkRBBCcL0RwsetB/jgbxn/FmQU0w6INtqAKL2iQqWMiJGEe
oOvUku2bNB+hn/72mcaYgQrkLnuK2CternZsISUlSKcRZN6STP/rjaYQeI9I1mJD
qVydoGpqukzCUQM+smp0D14vLkIOE0nM5w0Wu2XaSb9d2s9nVXpwvNww2mQZ121X
xiIQw2jW5CEm9jt7NsVl037yCWNGYJzUaYSY40mDp0zN22d9Png4hWhVRBnmQE5H
05kDzXRAdrhDD5y84lrOIKDrE5k6CrcneZ6XD6IKtwL3ytj4+EQqjhjFQSt/NAmN
t/SQlF++auZ0B0D59UizTWuVhpOWSVIggZo37TLLis4B5dt81hq0wfq4MZvxCPbE
Fzo3Dv5mPynzrHhFwmnmGK6Qgjpmb56LeRCrLbtU3dCNticKWDWFa48TT/tZrIkO
V75kXS/lCZPsESAuie7S+9eGfWpldDAW+uY2Q5BdteJGTReCX9EvYauyGyp8Kxqh
IjYDQqCsLoe4VXRcD5QEgY7HuxxtrFco5fxxD6Yia+tFyiOKJ1gOjEUhNg0B8L1k
H8lKU4Oo34VMqMnzZMvIr/y1uQq5InwHw5ZrbnDQPO042onwKB/zzXI/YGHIiPjK
T+RZBAU5RKulODtYhxsHreJmXWSkS8ixBcopUtI0/BgWAoaICP/cSdMAzmYCkpHK
P/OFiLpgRQ37t6fNvdH1Sjo3LIpYa5CBLF4ZrBi3lUbrVrjejP4P6inH39fX5Qak
IIZTBC4My5Q76IzegAqnI4KuvORnhas6cjEEj18157yK8ZVf5hmN0oVa12v7GdQM
TGqp6F2j59l8zqblAzQcjiU+ytTTB/L6guH0QtlIwdFIPSwz+1bi1wkEImK541bd
mXZ6wwTqgUB1bswEHkCeuUfrtGGmzLfTnfPsyYXej1+Q6/dEypQE6u5dh1SPmfxn
TDp5WqoIsFnRNpfS3CSZvg/f6UGBSJicMTgCWG7rAHo5+93T2XsBGJThIUJlt+R7
7Q7DXgeI8tspkub6V+K4YfpqoHrh8EW7SUmnDvWnk657ZHGkmF8hWaYlr3K0WtIj
5U4jcURahY/HhXFqqLZMfMM+CUJLAJaLpGQdexeMH3QF8Dbvazar0h8T3f+i8qXH
S+gTID8vE3stYzD4Z0nZSNi+wUhPII8+VZaGe7mvWdpoFbVhcoCcATHuhjheQ+mv
BBOHa7FqUEoXZxku2QYUK2Gr+2ScsD4AAV/DaEaCIwlXW6y7ugWrTRYGfBq9G4d7
QgY2T8qaWO8jUHzuzoICxw/uf0OdB6XVxrugO+GAaLxtRWL+RwLAEC0OTiu/fcfu
2Ll4C0NhHu3qXSOGOEpvHSryPv5KMkrJ45YAlT7eIhUu3JVzpi/JSiLs0fWasc2J
Mx2AoCl8O+KD07kl/+hqr9bU+OcW05HGUDUZg8NGs2o901yrbbEQYD/CSIXLjtGi
wzKVZj+DaTyOk9bEPRghBI2BLmRx8/0zRSwixzow4VkiSQ+ERpko623rx1CrCmD5
dLPtc/1wpbY4rK3RdLGeLrvlv3j9P6/2ZycPpjbTMmOcWodjtbp1kph/UeTYCz8O
K7IoIaFitu0nIMbsjNUfmL8iDxnZYsuq631L+bjeciGO1ewYQeOIusUJiR8wkfYv
tbqx9WLFohXitFHkj/kGIMn6Gcd/b1EP1DhLzH6PdvfASaeK4nKykrOQjeCRk+wa
YysFymv89Aeog2MTGkqaAEfswEjREcLzi2f/zCKW8nY0cWC7sGX6mu5QoZJ/A3jb
DwnRkGpLPKoIjDpxQYYi94FftdY5S3710bANBzGdJD+8S5vdX/BAm9gfbrAeTnAa
fyrejfKgmGB9ObUaCL6k0xn5TRC6Y5i7Qj3p00tz7EWLJQW6a+Ft73T4oDjLzIaN
s2CJg9LKxytq/LuUixOHFKcmz3BjSBuI9pHbI9S266wuY3S5I9OsGztiopymMPjN
AkF3KjgvOgi8plWiwyqcTsUJoUm6Fn1RJbEnzQsoBXFPIHTCeCPbhrbOWPSI2vN5
Tn3gxUVVAY8TvKZADgmf7vD4x1jf3EGNzqi1BaPHc0uK8GxI+XGzJYPsT9bLbew8
DRNlgxaK6zagmGh25mRDj9MTpAHLpFnseutnd55Dy3338+U6RPA413WHjtN/P7De
tTCP6v69n0asUyzf+RRcPCYArX5CgICz5A2ZqzAMa8v9eSARJslPz6+OWZPThmvw
pq0HqK7tzQYRk+1Ee5LzEdn9yok5bDe/riJmf8cGS/vrzJ9EWTF0N3OsNwjMP4v3
0MwUsv6PKoUEqlUrl91Pove/VmtSTp6VCmavDSHvUivyiiHkYJG4CJvA1RZyohwa
rwKdSBOZlTcYXJuj3oVhDPNZPEwoqAgIajBOh5HbsMJMroUAKkb0POFdhSxx0sI+
/s0chSGZ03AyHYKE4x2hs5ITv8Bkd/k3Z4oxjQCZi/tYjCvcYZ4MipeIp2HutTNv
jnh6M3fDvDdfsNZYPCCtnllnb/seHN6mQgxnbIPy/QFyksqLjRjZsIRihc/rtIOC
WVVttdVJr19r/4vXBSBo9a760rECT2aHiZT3EjLUR7baPEhI43w8JB6wN85wgS1b
JhD0/hG0LDyDjBkQaH4DMoz7ubWxV4mxmFBXJ7W2WDfASAWTF1c8WOZsIC9k/163
RAV7okfPiGi4nfPtkHBIRuIkHCp3IGsOuI4Q2y6+dAdQI060omhKmlc7AX98fvZt
GsXJbYH9jFNRAChZ6792AAi2RdaIUWDSP4UF9MDfLMXeLS1v3SKwtoSQ6+5WTKN2
p2Z4PGALEBYYwH+VxHHrQBRr2NGUiMB9d0/60/FutLfc/k3PolbUCGNHWcwk8UW4
QF2fiQzebpY6wmS0pSnGnO7QjvRTjmSzsvuruA6j0upaEjLjU9aRj5Q56Sv589zE
xy2HeC5uCK3OBML2vUbKPqHaLXVUP1Q9E0kREAXQhAm6k7w9XjF0jzcawuSnwyzP
WJajh5cV/2K0irFx88mC3G8nBHwUlKI2bn0DIh3eKFfLBVmEoB6xgKbG0a4c2ash
fjhh9mU9I/1NNRMoohcbWaIRMuRyQOAF1X11Y1+FXqn1DCktg9u4EZsCuvMs1Yfd
2VoVRkDQtDnEuLYhVHvOYW1RiStj6lqlFwmcCzxYSOj+aIKDfbrChiB8YcrZiakX
vQ4nBLstBeZRxn+PA0AQUzQ7ym4MiJBO7oMTt7/tGvP0mcTZaNx9ayW2bZP9EVcX
sWIRK3DulUtLT2/z2kFOPwLrnOrl4xNATWVcpkm3+WEoHVYzEwiAlGJgaqIPs0iH
d1AERJ+bWFrWIo3TQJ7LH5eByseELzmpn8hU+Q+UStwML0E3fg09pAVzbO3l0una
8GI/ecICaSLn0m9o3WALkFC5a0nYLfxnrzBrSkZRBVqpULO+n2qH78y9S7pqZI5f
8JVbe7b1Oj5yOpyvO2PWxbLYBw9/W0h1Ty6cOvO3/wYdk9BmtV9AdrxgF5cfDxSV
ib7ptrwlz5wgYkDHHi0olQTwFSNEbE9xjowPaKZ09ckvY/3a3lE8/6oS/5x8FWzY
+cvo7yd3lW3MoBjawlE3mmzc9E3oJhCcgtsH+2ZM3RI+atpGZWl1N/WVRje5EFjR
bqYi1JLOopvoUyXCCTgIjke8h13UZZxxZ2qPv1VDkOfxGzPPBKKYu7IJ5ZLA68gJ
EgfcW906g04GMbmcP5lt5ZTep5ZO4txCX+IfOThFbDhmLu+pJospDiFMrg0xLRxn
Soo+EPcs1RkLsMzCGfa+gT14RMhfHet3d2fDnlqhUjnHutWK8R4GMOt01TDIi2Wq
fvRA4J9pCg7uqhvsuMED3ECpOv/AGFrSFoDZpytsOfMlCtgXKwKQO5e0px3OW6gB
uDH7RMUXXyUxFm9SkcyQcug9Ss0zScjMqOQBoWPiSkpuVvkdnUpD1i4msxWu7V2q
bvS0sW4iEvhB/YclNze+z1pQrldZ4EJpqFt/3el04EDojagrdIM60K/qEEUdB0WE
pI/nGDBSbkE918qTSsi0V6TtBBr2FsDxK43tJUjEMvVtFzZpKb8ohbOePDB3z/tN
ecHz7makKCaMPf7VUe2t+ubUGal7lMJeRgpq4jNu1faE6EHCPVybjM4oL2xfoKTk
fdaSKZ0LpODQHqDDneX54XePtc4KdQo3RHvAdKlkOoFghc9T6BmBBiAJ6l+5LilO
WLUKNJDsR4eyzd1UMO73CvRFoPJnemSKweMcn6daHrfTZCEDhwszi0z67qGAZ4Gb
El1DBz8wazy+XnA6yQnWgbMc8B9qkQrfRenCigrSvHE/tSIwQ19Yp6V8Z32vIs09
uOKudl6gI6bkisIXHA6c1WQQz1mMoE2jkynYEwzn4qvXR3UEthxlzwjAVr+7+2tf
sLwD1Bfz2LMohNUHberEcYuWVMg1ZHkrkIQHLPwnHUf25VMKEOikJPHhExKYIy0q
24GcRQoqmHdC/u3zSgOnRLeazYt08KgxZhas+SKgxWqh14FV9+5VrBOzQzU4iPGL
K5/bDQOb44hs1XVoOMVEA7oCBMHu9+yK1Fou8767LfZoLT0Mrj820k2o4NcxoLqa
Onram4XkGHa/tH+R0onKkGIqCcdKy3uDg558CP/VPTptfB0vrhku8Dj/ABXSi+zP
+5l/2zAgphGSAEYY0FIH5VJaCj+LEFKEe5DYmdPOTodaxv7UUZ3+Z0Vq5MS8xeoe
WL8kNWJjS6jgF/77WknKkxyf9+Xs3SjdrnJD2htUxqQX7NqBWiwa6E8p/qTBN6cr
vRMSDBcdnW6Omg++WNwT1waNY48f3rDtW0ygzEtkBbKxnZW7w9/ewgMrwv7i0yes
7b/X/RwEgpnh04qxrWX+NjX1C3qNOVeo5mm/MliX75yFh7ZbiL950UPC1J4OKnJ4
GJfaEJUqiU0RoIouXFtlK7xyFQgROxFt9inmGTgfh/FN0j6udhJ3HmgcbpR4D8rm
/V7vhP41d40Y/4CGEVI6x2kefsjjkliHo7jf2+FJ4UUij7p/RDO3162/QDyxM8Le
+vj6fkXm6uopM7baTEoJvRqmUq5ykq5pQP29wu052VkpvQXmTSsBv4IXuZEb3lIK
KudOQcIvt3sAQwZ/W3Om4/zyW7gBivseJP3IGeEGNBElejWnuXH2wE3WajIxk8W0
mgHPyUcFsBTfwjdvRqNxSv/cmgWSWrZeU8JAN+a/7h+x9ThN23M8o0JvPYARbxgL
m/qTKP0Je+3uTN8NfvLazFL68vjhkbsyxqQtvZF6fBebLxVr/fua+ZgXa3sg8XF4
UsYPqb2Btxa7BpgB/frU3HyRlcmgJyV+pYYm0hvSNxQ0oA4IWAEL75Yu82nqFbDf
Nu1YQ52XWN10kr7JB34IUewfgy1pyXrltzJbliA1KqKN5iTyCdWjMbwX8l6pb5YV
/PJoLIZ2C1/0+dtlSCNWHxBDRtQ9kfZAjMlrkNIA8PvT5tfqKMu9YothEtaL2WZz
2UNgwMxCX9dWlGb2eRDuZxWgeep/NMwFjYXiZFrANsa5xZ1HVSzAhNjlVzp/hESE
v+F8r5M7eNPTZa67yi33QfRfaDDQ63a0BDDI0uZ7ThxS4fhk8C8S+W2lY0kmOLux
Xfw2n73M17nemi6P1kjoPzdARSiMLt5AM1eGzjUFmR1IKIHI558MJl4b5O9Mgg5i
81ZXkH4UgeK6VdEgB14PNc7S4il+jc3LN7o+aRN6uWvxLYSpUZzRk0HiAMM6ldLu
emcqXAvj9rAMJoLGZQwQf1AwyRqAE8N/j75RLd0iNQiaw1f6qCZAEPEhlp0OlaSV
SC/tg6ABmHPqBpvaIi9TdcP/djncPHWNfygHTuBrnn/5jYnhAeRA+6sugsbQ7E89
wTSiAID8c75BHeNOwna+gEOe1Xq+oPNSGKdr0JPCdJxBNLkvhzq9gfYjwxkDsJO2
GO5RVFt+uhi2Xx/YUGPQ3xVlmw/9fyHUEOCovVZnIW3xxf8uF0V4rOQJzY5r0Z8v
5fXjzZ4ESqu76iM5xPNiimDy6XY6iYbuv+S8GeipCN4YICIFemJSqns/EgLtTktd
7qIhNhKDVZSg+/GDZwgrunyhjJBYW1hB7h6b56MsRAvUOVkx94dnFtNDVDoBgf7k
ypxEeGDfP/sO9DvFmYXZc234D3ZHdHg82+Ilr0wVaOq/dQCyabsW5ojg9jT6PE+l
3/ftqaic/JrNfElTa0lFOIp3Y6NVGK61XSf1zCpuXN+byNJBL2FzuKhI+86Mvk0g
sv7k0xriyXx7cBQBheXG1TltIlTrK8Y9lwgjsqEaAt36cu5sg8EupDoi6sed7IQ1
wyx8TPSR2znYYecn+Hi7KCBIYDR1VtyuOQLwVWcYskQSrGpmA+absPMs1sB/p6TW
/SG9KXOO6L5qge9iofmST0o2a6c5Ayct68b/N6cmodL8qrFaXnuF+hVGVeRNm/vs
MnW+eL+hSHYMImayf4P+Qkorgh/C3LygjAjFcKJfW27AGk30PobQV0zPsPdLfkTF
dHBVvq39QvUxaXBxvJl55/aETbEzZmKIGpBLqGQuiPGAF6aG1YhMWFIQayvlt5j2
SQK8pDq3bAM01ZuXTrse+j3KdKhJJ4TWi/YgrYjVs94VNT4Uw0SaK0u1og5E0tF8
qv6GqcaS/TJ1Ibk9W3ueifqExG5SB906pWqGzIQfrJQpjhLnc85MhWKPDNfJox6F
WwIyjgFDmJMkDdUBTyyna7m1pL8i1feMPHs4iQcb8YXWPlnijXCLKMd8zQl8oMGL
7N3kg5WXxwwP0jN70DeHXzu0v1aXrcRdGpuw8br5q6eA3DkV/MpBxcTbqNSZsdUR
RGjNMHvln2HSU2reFKseFOCuzZxJtSfWKIVTW5fEpe+Rf7IAgbNwe9Ly2gwNliVg
0eg5u2S2423Q5f7U5caTqkfkAx6/tbEPI5w8Pd4D6SYZcMNtUJQ8rAeRYIZk4nGG
707jNUQV3+e9/iQE6ieMeBfaQrW1mDGbJzoTzSRlkezsMPz6jJehxeUHLRXdMQhJ
BYzexmCFYZ6xsaXpvXB2cysQRf5heZd53SzjqQsOlIQDVRW+8r/TETklfQNEH1+6
bVS2F2yljI/NLOdF0vRCJdQ+0yAS8qu7qO+f7hZHJhwj9X2PqtGprObNCQf1tQF6
B07+UN5c8yNxacxcmbEfhJe9sIODXOjwvdCO85uzSzv3aUY1xP4gnvA4gO5XyHXl
eVNAEj3YdlVCnyqRjf5i13tKFirV400tww7kikqaRRnk1oGCRV9h7SgKPvWdaUIl
L6Acmvge6gJ5qzPGAgNoH06PTovuVPithD3WKEkXnbNTS6hg/0fSiG4Y2AJtj6jw
AAJcuItJgACdbVKBbClJgYx0lX14zBBb0nSWm3qGcJDwebwb3lMuwYhXCWo99H+f
ahZAqNYirg+pclgnI/Nluf8TnY46atZOew8EQsfljHlo927TQml9kBEmNbcz7Vi9
xaVKXDjOoqrURfVXeJq+3MdCegv/5Loz11QtT0m5FVWeqNJMRgQvRW1/abMLzfNj
EZKBPL+qNC6xVIE1x/HgOAbj4kS1ItP0dU9xe9wQuNFlDWOQT67z1uRz+wcNysey
FO2/RGCGzYM+UnizB54BzP3MuwuIAVqIofaXGmIYPFVYFCQbZ3PFd3jbTJBpE/nG
G+5NHt/mBduYeXJeK0P3PMXBP19+fhoRNzTfWM8Tkr6jjO+BqdhXbIaDmBxrMlNi
InEFsbxijczASXDQDCUropXjN+6WlC1ChlVHv4nu0E7fiz++bH0XYZrCZu34py9Z
GJVym8h9TzTqcrhDOQoZ106w0UIj4slq1QqR9bk5DkWhF8boDytEYNHlt5sIxVkd
WV4iBrvgdztV66ipe7+QtIKEjvkmkXibzZ0ShgM0rAVvKDkdmo29znYtpNWUj1EM
LeMxmZvXBXEhvIvYjtMbtAxd1ELEvYhOHKMZDWYP0wed4oLI3topKoDWVK3UECd0
AkgrigeY9gyWhN0suaPksvZKhK5uGQ4/GYs8LWOIkwVeaO9wMC1ysP2E+Fe6qpp2
bgMplSEYYeOr5DSPAl9phLHdqZKTsO7Fb8kS6u0yYU8NbzZJEiPl/vLWAO07LGkV
bmstbZvnzX7B5r02MrQ5p8BEXwHi4q4pUxqWrWZkNpapZdnp78YKpTy0bFtNTf2m
V1XToudzguyzHQvEWE1hpyoYZpOWZZ1VSEyRdN+nM/W1knEVHU17CoGzT7vy4CN1
N2CYtu+8RbhfLb5yB5FOsjUBh4+oSBs7NEvTrYDVN/mZcwA/hmYf71eW8o3+AA/a
hHNjwVTEfhgI5MgK2phgKWcWNl7XQt0FpVMo3LY9JJl4y7Ddr2yWAS83K/6cg1O9
Rp2NqN9Oag18tmN7M3xbbpnyTh0RdV06L4UD7To58uBQq4WrKW7qZUaD5aqFrnM1
OU/79/Wchr3GGgMQPNMAtNlIl8uFqq+grcjhTXRBsZ1MwOp9XbrSVyvoEzQqv6zs
pSYXr4LZR/En1mRmRlj0nfiivEyEP12tM8GgACT9MN7Hom/aYuIqKYAUNAU1ignS
XIxYzlH1m6Uwpk7uYeJSkFWQX//KQstjEsacB4fNwwTOYONHOkP3XW6hLtY/AvGK
99Ai3Bk6vfaIGaEyrsLws4VCt6V9ddYPKs+Cm1qDw6053LSNASNeokhQ8KsR87kN
xcEnpa4hgbz09KNQBETEF1ke7mI3a7UAZyvoQyM1N0BK0/oUuTGP1ini/zm3aGQX
T0To8FfI/rrketqXKeYkPvHnSOPGe5dgXsIToB7BOgb670cpeV06xu88WmJhKH0T
L2Nbc7L0eVDcgQl3rGK9SA3MSNv0GYmsgmUGZs/w7m/phxUrqHRnM7ejgdSi6APr
X6imHYRRMQSC7KXtI0sTv2Ro9e1/mxbIKwNqezqeG+SHhSQ5AapVWWMCeV49HJgW
DUjGPrkTuzWajKvRC2Nc3ybuIainAmJ5nDzjm7N4LnCxlYVDsjNzqgpLC7NA7nbG
fIB3lczsSHqjXagkkO7fjG7BLMyoClaB7yDa7xKMZNRmBZNaJwF/85U0NVG/EnxX
EsAn0g5xjBqUdfgpRHWqOrfJ6Jun0mhnWFijvrDv940ovFzLe1RkGhcM4Xk0Fv9o
jyX+JTIw3iND7p4G3061BQtvRSzkN3oyFiAZFhRiPkQTGjuNZ247Vc1+XdNXPRy3
hy8TMUeAknwFkVsTsItea1NMwUX9sgjVTsiae5U8V0/SIc5CvWnzcfrFgqVlzpLR
/8KWq0sNCo5mg1Dg+jM78Z8+uvv8zXSZzmkX8iVFZY8Zpj6+/5lNU5KrkzZjmLdv
0ZhppfXjGl05+lAIUw/RML9VTI//si5hULMwuX2C+ASuxqqkm0qsusuzyTejTGke
vtnAVuaMvYNxjCImVEwy6MVtRgKhK5MNHMxEjiYvIMH/FaYA7rrhrBd8D3H4i8xz
ZWd8r/LSf16iSaYoZUW2iLRdyk9+8AqBNgtnPBC34irEPHEBAAdw1/gT1V78xhVF
bYec0K4OQZftdrBQtQlzQ3fmTNkexJk44kaFAI44FG+lk/EIwPm5Rm9ksTHspD1g
3x9oJEkwSX5F4UCd3iDs0pCewzM+wx0w53FV1U/alyG9OfsgfLmZWTchYpY3V5dS
m9STxGW08f7nRZeGA0p1uYgeavkbSEU1pX+VTj7M6n/f+IChCBrif9KmBUl0PiDO
+sf/5h+Atnem/67lKDxSlATlAjzM40RETaaE7P/egBERkdUo70oLV2aTfVhiquTx
8XfGdkE2rPIe2/WGYdCjkvdwPqXTuYpjyGFS5kNICQ/yHyCK80zlNoThGJCgvEhe
9I+ZHy9G+r0YaheYNeGVMFZTFoCkZUWFW2v3MYQ4VfzoudIuZK1maGc8HR3mrxJr
Smc8egFxA0vM9z6s+FJ1MX9LiT4dW+nlNytF3BRa0aiIpkgvWRUrtlBCGpTg6CPX
tlC7jmkcMHJbtegRVu7/7skOqhEjjJfQ3zm37tzBYluCtUA10cn/9W2o4wiTn/fY
Rzr64c/2wzqUjga7zRL+3eQdBIeodRsYZyqgmUvHJo9DVkvC87EEi23HxxL8W7YS
U6aZCxWId0ryqwY60hheyzZlfCml3ZbseJgld7Ai+/MdXrAcJs4iL5BiP+R7xRWR
vVPmZsXvfpMjI3hxILtgQXkJTfN+AVR+D3jzT0HJi9+B4Ytbgc1d42jHLradlhNI
Hw1vPoI5rumGJ4xIIrVc9rPFzHbqqbuqBDecoM3mJEJvFbnxh7JtV1z5QR9Be7by
DyF12hZ00j/BUbBQWTpuejjrsFwDrYR54HyfOtrgF7TaSrG3rwQ/xMamYr726xmV
EiCMNdAWvkATpYftDYyxsPiX5yII3FE+YByiJ22oMybR4hmqqT5kH2S3fKQ9TeMZ
IiLkSEw+ZRZkdL3t2fgu7ZFF58AZeUQyHDf/rSXK9V1ROLsZpxRzqeTcMcGiCdOJ
XonKs5wGe71nUzRtWCObWQ9Dl6+PbKgY9Sh1zqph6HiqZxqsPajBiqU37tYCmlNK
Lxt2WmcxOtTTNFNgWI86xx5n4psx8BkSUXp4Ad5OnNjcnJaT8wv2/ibRy2glCkMV
hGkGQzI/bgMXQVj/TVvEB2fjiZX5B3koJ/eMfKcS0FU9bh5ExTttxhODmTCUU6ze
wHrXumCBTan1J3g9+RMaEsV83/TVGjKpAU9l7233OMHRCpnbkvIE/yxT0zwIfc4M
gpG4Oz96q+/Fw9B/iyjj63Kf4ASo1lmZU5Sl5hRBFp5o7FueGfNtc7iVMnhljtg5
sv4gUzHVE+LqOeNAzGn2fj6CjBcdLVM+JYSqjOfFy6icn6asvnDF3P2EokbZJZkI
d2scBwu1I1vq0/zyaZo8rhuXw3XymLKz8yACW6FymMO57W/mOhTwvHx3ols/U8q0
ywqBOeAfL8CRh0PPXTt3sHzOEvCnWZCKWwAISCad3K8lKB3z3nMuahEW73QGcm1/
WOeFVfzrUB9/ZVS5opTB98zmFd7eLbQM2CnkPR2EFzIniU/bf9IClhoUtJgjbV3H
w8wZtFxTUZZt5OTVal6HZWMpRwSOyHX0421f1O9vsemxYbJ1xQdZ9iHcypmjSir7
uoJb8fYmmRBkhQnqw/xN+pMyioG7+jPVRj6hbsUPCRG+WVbisW43MVL1VqmR879S
VdLMyKsIBnvbVDyc82x6xpkb5xHu5kvb6HBcmDycZr9Wx4qQAg1MijYfAecCseg6
Ke0ijZDJvIyT2VE49fuEEnfd14PkTiw9TG/S55Cf4HUtBvus11pA8A16NqUoZPbl
Cj6gcA+oG1slyoz4Ay4qfcSl1QrOA+TqLzvALv1LPohE+jtEO4wrSsHhCiJxKF0i
NpoHegDV5tzBwR/EQrhBZJ/YwQb7pln2WsEI2Brbh9DdrLxf4uXNMYHtiFhvN6o4
O71obtaYuRJxiQPMIv+pg+W1jvjbOItm+7N8ZaB0jER5giLI4QGWeCD201ksiwp1
AnttDjfo78lr8BifsCS0789No8cYatUGozLIvnSfieOl6omDI/OkBHbxT+GBR/HH
lNY1Vq9tg1kodKbOqMx0KsQW98k2hbE0+B03Y/Ltby+tiJR2/yMJ4NGuOgINqvt9
pUojZPnYPQrMFJxhprEv46YilmB/qQjYUytXS8gB0AEOmvB/hHdJ1TWWOkCctsLf
DlMyiOK88UQny47WFMmYAhfl8bYOZZZuMwNHthyVSkqKJtR7A0mP9/XfgAhmicvK
1Y5xeQd3YQcfw9WDeeM1mvsPLVV2gJe3PtwDVtB0HgoskYJ5in/gm0iVjN3b3m5Z
VlCMQLMpyE1zWF1dixLutg3O9QiKEepCwEGHQ74abhwZzjiBB7CHmmY6AT/RdFyb
8YjCpFBlI+zejeJTKV2lC+iVsf90ERLPxSU1Y1rqMAoLuqyfgND1sVvYAWhaYcE3
WQqR4HmhWTFq3/UHbT1xzQKItic25C5jEb1EnFVG5hPGZfcDvDK3AiQWcEFr1p6C
A9V1nDNO3ioGiNtQGUXJv8CiUctLOUHQtz73USLfKU3J2GwW4Brap6P4pAQsa9Yv
BbSYBPbE5tvx62zvo8e0KOqS/UIpP2EhFaiq/I9etu+Z86F1pYfMr3eFByf67KGS
z/ijpI98sGisrAWwhPfdXux/0BTtKlWpHWoND5qhX43yl/rpINd2yiXTsSqTmKtU
clVtXOiOCBi1zH+H0EdMtV0VzES5doQ3RYqTGt24Z31TkzfvCWJiK0G/S9eiCkIE
CoCBiGow8BpskGUdVDAM8wLdz16QDiUGkp1OsUNl6B8pfrUATmZ1Xs3EUPz8Ts3k
DhrKrQ0fHjCMEEIIAlRkEhJKbvKAkf8872E//VzawiXXFYCsSfakN9rhqQKjUB0I
Shm9p773AODvNjJgVBls0oE+BSQK+K1rYmCZvS2OzSwjbL6tICXGBe8b1Avqo/UO
1jr6l8VykLK/3uSlN2aJtzjL/WHuTrVbnshZT0zOdfjOb6hGXWgsIo3W4nX9bNlb
dVgd7U/buAydMbE8uA1I5kl5iQSARcnga7xC5GMzqw7uI0LmuyXzylgS09ydnS0c
tUYqY6SXqF3VW2kxm1H39EILomK5MidZI646htFL2mLzFN14NW4xhmCosLpvGMpG
tWE/ld5sv7uj2obe6WE3iE/6hWX1iMVizijcvHFxtHT5Sp2IUShnOutdIcs/VsGV
/ZRdslbWym8bmbuSolnhTWHCZUYw6/p5xoEYRDQxSuYb38lDVLqXeQothgWt6zbX
Dx/06LQCC/3yNX1YzVtDT219QtCSr09xISFfjj44v1FV6xezlrU1gdtfpg00R7Yk
Qx4/pBLQwCXxXUAZVE1HD+QP0n1FJb/PNZ3LOxJrfKrnf1XR1Wwg4qCOfEuTOKcM
3ZOxIk/WvdqK6oZfIaZu9UlGPWMWTXiMnem2cdwi2WTfXVlFFOJBbugM7TqJWSLp
tBdZS/VO3Nxgc0Tt1iWfU4Dpd2I2gxqm71LlFPWLPEcfhza5nfFUxg5lWwI8+OJM
sOEVHjc2HX9/2Tf8qZgod+Z7eg/0P+pyccg1vEEPXMjxAakZ/CShsPZV74Z3mOe1
XdEwS63Nvj4wLsVG5F/bMlvEibzEimHZkpVfBwC11ODP3ardPu1s9PnqvUh7wslz
HOIkgNdVnpQKOvT+c/oLFUJJQpDjsg5+mE4kRNEMu1HcoQqx/aEBrk1XBFh1ED+S
wQ/3SCaaFG0XCzqbxt5qd218Tryv4BSliFLMoeNDnKo/99FO8zGLeUZC5HjM6OVH
yJzevaHZgEUA2qNfx1NHkMvWMdMKIIL1RlLPppHWkmeLOjTutVYVZxCIvC05nUFu
RPAQhW0Jk90wJ6bgvNTnicKgFmTRPiEGLLwYcTabNPnkgZNh7+YYCeNKRU6q1+JH
gaMRD93yjlH/OwP4wuGQEzrZp63KLMCxs4dMrXnGN+nv/sUZkXBFFRXC1JQIb7Iw
q9ZTMrijYzDpvcSI/d6y4wDkFasyI0EWoW6tb4qPM4oQhROWjo6lvWGErU2TNi+P
1w7rGes78QYw11Nu/bN6XNCAmIix+oub6dck/+pqqAS2FjOoxRXpDA1AgkCcAKkb
SkoQ43IGyrn93FF5knxgX8ON+/Qw43n5D1dlpVQXKF9kmzp5Lvv6DqjOHP5aHYGZ
gWZw2NCxvebVseiX63s32pa8ntKxkTvZJF0WCGXFMEMWAYbDjjawPDvELUuFB25b
pbeeWasIsJMaEMicfLkFIOFf55p866m9Mj8YMkAXHhqZt03maPblS+ZjpwVXe/P9
oosyPe6wpHnwQj7xn50kqfpSihqQwwegXC20qQKzol/ESFyjlzweju0toWuAWgBI
NzjzYWwigxU2YDUc5n7PlMVGhzfSCG6J7UQWvgVP4lsG1Vkr/LV1QkIVBfH+xuIF
wxN1wIMmh/TcgPyllZ29/svE+fnR6uNhU2DNRJ7ozqISK8/AqfkiaxJ5Dm0eyhsJ
qWjohKtPrLzILgkGIuzl/2zMG20Vib6sXeAoj9EPZelmBen3+h6GAV61jQyVKi8G
Uhl7keav865VeQrctpnIvcQ2BwSrQRMa0EW+l3HFy8J94/2OpuoCBY/l7vdsb26b
5jjXD3twWf3oZGQP+JZlJSzM/yHEW6odobWHb1McBGymU5Cjh5tN29IZYkSzWVwg
OPeY03yPduHuDSnplJmiFHCv8aYQ7LxXKKL+Jvy+6YhLjhstfwDA0feZ5rypLO59
AJCVIf9hOHAnU2K5/usvgjhLfdCmgyVTb+/07DOAkOpBnB7B+KpPI4cf/kyJZhGA
lvJQ+1+HFI3mnRxanubjKlbtC9RPbAGysU1MCrlOUwBhCI19EqUBAfcFspUbhtVY
MEDm08mCwPJHDfliYCrFP5vHHJIi2xZCHHy+ylCaOr8pMJ+kWDg6IBXQMqGkYr6A
Ijv54b3QUAbshOUIhgYAQ2QckjrARGjuPmnFB9eyzZcDhociin+v8M+QQ+kIXP/1
H0CZmYaiub+QZdWmJuJt9K1mb4Jzxy/ZrtMfXdgzbo2zXuL317/djb5unKVQQGcP
jNaScEDHsy7ri8rOucHJALbw6o+8jp4RWpKy+WXtLlrTaMt9DgrQbV9igr75vKr1
al+k5MFNC0SmRNihmjy/8diALqQi87z51eNhKsgSlY3DVVE2MI7ID6RANDN5lZOt
tQyVU90nPMCF3hAMD2/ihpPUT11pj5YOqc1HowjIKqBXZfqUyoQuopYpch5wtdaN
fnVdvxREsMQ14RSpy6Hy9AALLI8eEWmruTYjvF8osFZTJMPZVY/haVZGjJrEdWFw
DB8LKLrInjBMYP3yCuG7vkyWkyVXCYnmV6xec5qaKfBs7ofTKIrRZUR0Fjd7f6rV
VKuQrr2LggtSxeIE1Cf8Ry049mL3GP3c+7iM5Ec++RXsD/WKhWKawR2So8QVbmlm
SCAPpP///OnPwy3QGvC/tLlHQT60sr8yBCNZg/3B3bdb6tZNbh6LfvooEJhK/jml
xldrqA7Pkv2n4wmADMZIov4XsmKQMMC1YM1Mn1dx4sRS3OgdbRePc9c4z+pRQAYq
C/9Y5RUGMFTXc6R3vSZdlE60DzL3cXl8iahazinaYjFC28fTC+TZYKaG/84hpk9H
E2/DBmLdTgDC3I6XX0Lr54lHa8Tyw4kR4WaBWpXrZwBE3opZKspjlt0JofToe82A
N20Zg+Q4IpqidXJeHcuzhoSe8Ta7E/7PADJT6difl/z2ceIE3MM/zdHYhVKTdyr/
Ah9gqQ3/4Vel/S9hFyJEvlPt7UQLEbAwGOl0RfhjY6LBTjmOFUVHWaQXEibHt9cp
5YeXKdQI9vOFxo32u2MlL3ojSXVxr9Sv6yQfcQxGrH1KLvO6rC1UsKBN15E/HDS4
NOkOmMz6c2rgkKYkfQ1iwWbxzBjqfnAs67t/kixph5O0Opl1oZof6oinTX3/1GYZ
wz4ngpVNaVHgzyWocVhwkzcKTT1K12skz/rsvHF+NDMn9HA/EqAQ2I1Twuwo2A9+
fafl8/cJB6kVEvdsPyvc2xa1MRHMfLnipeyf3T4N+T4Rr++pIMR8zjsd/HBIsne1
xE5DvecwcWWToNo8ImzJLNJdpbqvNW0wHg6Aqyelv1tKEkvQ1+1R09mI0DDTn5LQ
HZ4ycFGOQOBk7nYh0S4z2K6MBgzV34t4Whhxs9nEsS2USse7w1Cbc7/Piy6g4kro
KydHHkQmy7tP30Sz+hNOGT4RwPbwKvXFIUzhAp489r0fcwuXQldFqfGWz4Xp/3ri
Cv7G2OLFpAY+qT1+Gm5ztjPyPMRQLE2GURsRUzJqp6+Py7pX9PtOL5Pes9QPgxvJ
kP67K4rTNWAslDTtuFDRbz4x/ddGcj6bKy+MM5miL8BPJgIgU6yIx2hN5WLNAxz5
J94WaPLYP8Tyi4PDHz54LuW/6C0lc7Lah6dgQkYCfYNWu0f966bmKvZZeFbf2YJV
tFRi/kqfv4kxYuZW8lHo2TQl4zai578zzNRLCN9Sms4o6qqWy+aY8zLY5XiXm6p7
IXFczP/+JzG4MKWofDkp12oN/UQpRgX5LwINl1jWhlc70sviArBvuYceb57uq3Jv
15tE1kgZR7KXW4GjhR+//jHYKFtMllA6WY4ExamBhFX7jdS+VbeiINkpblu79FtM
t1w3NvbklIBeZKMsgmOwFMRBCbQ44Qql1BfbHLtqTOy80YSqFZJymAeEPZb4KPQJ
FrcOWT+m4/HS87imHAnQNO63dSkxXOkzophC2i9k210zlm1MZl4n3v8xX3EOiO4B
03HTHTbgWBijRT7T8D1d65T8wNmBZSMZL/2JL9P2yNr4N3KAFUa/1eSWOwGTtGlo
3WJTrkCGie7Y0f7QhQ/tg2XFOGzlKs5Xi3/itoqzR0YLH/pEbrzLhuzjdd/MOkoM
3MCGsiGYg7dQRWfTr23DI//nS/4glYxV4HTREjJ6fypgQwv91cN3pefy0zeD1SK2
3dL44VWxI77UaDxT92kIBQksdwhkzk5viR5xbPwhrGJQUDgunqDZqtiEKP7Thbav
cOr4dha62XqcdysEqViU9rSxNXaqT6hb321yyXdgmoDP5PRfFMCvqZRFQv/Yl1Ql
y0YtPlPQC7Uw5DNLaZj+bSVrSsOpQia9nx1s/T7klxpLQeqQy1y32nRsK+tlEN8Y
hHAzU1/T9iqeBKV8uy9B1e2qmCiZ2Gv0QqhVCTR79M3A6p1fuOI3el83nrAbKNvu
sEdPTpUG0le3rIOO9ZqwqY2bWzBABKoZqE7SAjYewA/PKEZ5Z4BowKSXVGn51jfU
Qh5C3iv7TE4aeqBcPuuKTqksSlOow76pFVQatbcaNV7Tia7ePg3MlohSXMFmVVhb
cvtKvKH4wEFajt9JCajFKFzC26CV+6Wm98Apnc4eZmy+RyBcC1le7a7UisBQQ/ul
Ta32pl8Ispse/OshuYUfChnKl5mBFuSocMu78KqXmJIWqtQ7slFXoR+YPP/xp0Gl
IHBMBsr/ekssQoJKGd8RLftB+S1/HCymTStzTjscNPglxfHfhcTyl1bc23KjZaBh
VuSxHryhZv8w9loOApefjLc8SgqPJ9s74MFQju48g+kVuPrXavpL8yA8KNPQApP5
IfVVcy8p+iXp477xUubqUKIlk7dvFtAW7eyKo8//YMycH1GxBb9Sgu4VrHKpNkLl
TzAHRXpuEoiZJ3u1SSJy0lJPKdK9wdcd65tbJ1+mfa2sGTcmgXrUpMQJNCGkn6+4
d+yX2JHN4CtskMt8AxYUlJwk4BZuBZrOsOy85TAVDo+OLMZpjjRYeiIZpXriRQjY
JykvxWDL3g0zlkvFlfKDJh3JnuxkDR+2qsnM6zJnnC87agTcmokAwvbUIJrnjIpY
XWJ6giKMrEry3TTOuc6RqdEBTIc9uPHmhUz2FRjy2nHVbs0cHYoDTj4EAXh4fOmo
impBFOmfaT6NeQiaTcoaaUPecz6lbEIHv1rym9hvcgTFlHuWoeppPkH1RQhHFRgP
nv/ATj9WrKl8u7GJ2f1fthckZAEi0iWwhMapPv3FJVjxH93BpWrCozQw77oTUJsW
LlPYWG2AymxFkcgIzhoANbnuRI+VS17fXmH3xuyiGxrdiXyZ8ffJ+eX7qNmIpwlj
4F2HOiBUtI2rJGutlBZ5z7aZiDgQW6jSXtulU1cLxZel8r8nWTrBWOXWB9sso1N0
J7atVf68LVNJ+uEUOrDIhdiC84Nzu3qs9trvdmSO0lPGm2e66TIRHa9q63GkipDB
IUTtX8+3jsUzL93et21mxOW5E9SG1/htTWBhn749Ftcro61Ip7hbgowWGDZw5b8C
PYza8XHHH7MvHNeuhqlbgaHJVA+aeqNcooVn/eOdleY52et8HZLE0frV+rCwysw7
60NRGG/6idViwK24Fko4oL5piUugI3ypgpnR/7c/RJom9eRVIIZR432s93tHkcUY
E1eQLWjb2zbPuv6hQQO8wuspGDFqHvlKWHS/mILBEv5+kUH/2t3l4iqVY7XX4kEl
8ROIZNwS316RM2kjgSaI+Zm3ApG5IgU5OwEKg2mokEdXi6uL3YIDigSyFf1hTAIN
rXPpE2MUfajc0y3AINx6skf4CVpEBAveBO69KFMH8FWgNIVIKJhj6BCmcu8x6hAR
nVjzYfvbh79ZG4Zc/zhhOsz0jWCDY5S/R0gxbvyIN4aQCKMEus6y3mOOnyHcfiwN
QIyc28M6fGbdfd/hVf4vRTyPkfsuayB7GcNh2ZbI4FflENgbfblI7UC5cmKEu7bW
IkjnBjMaPomIolOhY4Oe9R4b8KprYieTKpN6VkHAJctyXb/qRbvl/EvEyaVQ7ZwI
ID6JQ0j9TKCRdIVhPdX+9p+x5QVmgPwiyKi5x3jcO14YEhuV+c47vPN4GvWtet0a
h1g2hJ1R2piEhhIj6vgBrdmkqeygO9Kimv7xU83Xqq1xBgTfOX/dgFSHzxYgXJJq
SnlNjXeMaZRSLxr1Z/1ifAOYr/LkToxZp+mHMGCxvAjNoleaMh3dojtzHTUziEzC
wxP8jeZNC/tesA1sb2EiOxcE66IdcXSoXVcce7YXRdxtyUcT5EbqjKvIG+E15j9v
9janp42Cnb1IFS/AMv3X8xQ9KJgCrvgCRcqKfZnQkragNChaa6Cuh9gON5TcRLLe
+GFDMTrY3vncaGJmaZWkQ5UyI+H6HTL7MoK4VTGQZO2WEhyfRbDjF+clOoKvVljc
KTiycB61AU6leTm0mp+GydjvlsX77wVfI2upXOsbFgtOTU2/j0/UaFeNmX2GK9q+
SgBywXb+yh+apRBN6SENSNG+12fqSchCsgBOrP4FzqUBAEzFBxJp9xzoczvszgUS
UI59vu1F76kAxPU8mnXOTHx3pBUlj099E05JZehgHWImz1wbPb234JYS8uNxkYXc
W47ZpkKP+HNUOXNdGFULU8fwl6bd7ByCXXrrGZxBE5u39pBmBO/F50JAqZlKwRti
4Hx7EYQ3dzxlqPmLEy+Iixa7SOVjnomvJNkxwpkhtit9jEojr8aD0cjaEtQ24viY
pJp/54DieDnvp9N/ABxlAvuZxbqiRZPylV3n/jcvGbxEmejJ/Z43aVNG7nsPYhJu
cZUA9jw4H11OjpgjSoVkPXdB/r3SQlVnWVb3cd5QRv3Ztc8MLM18uHKAvd0uKt6z
zBThYirYp3HoxZd6KrA3sGFIMTgk9Xiwkmm4j4IZISlPDHWpiXBEvLFgB58BJ+99
fZHm9K8m5fJ+O2hGQud2oHZZdgnXEIAtTkxs5YZEr1xOcye+yiADu3voTmIp/fCJ
koSr3Pwjh7DV8nUl50HbMvQSEPzloM4dozsap2u1n1K1blqHpaae71Dxe6og85dm
FjR7hFVwLrSZ+pT9TLgU9+HojwWc6dUw//TQ/GlZcznBN6GSoiPMSj2qY2a1jlH3
xj4VzIJTC+9MPq6qxNXqnEmrSI7UDfftB8M9kLQfjc4t8UV9OunOGu1NOFggaMUL
Gd5njropA7oj7DL70kwXrXGIGKmjU4HQTtQs1zHl20CHzrYmn1pP8lm8zpbrPJct
J36Ket1z50MhUcJoMPMvwI5TFqozAgbyLKomX28r31mJth8kQ2h75f4KjzQ9KHXn
BLZdlB8Zw854QTmmq5CBhfMqltQG2ciairkA3iFwA+fqtM6dw5LBGqujh4H7tItd
wW3FaAbqrlTsR49C9UzD6ggHcZm0HgPZaFQIGawI8Rw41pWGMAMNu5Cmr7MwD3c5
8mH6Wv2jD6ZQG5/CwupF/j33pf7ZjGMkO59NB9vmnqVHLbSv+9O8iNqa+PnT3SdL
xm4K5y6sLjz3txgnNgc4pq0Or2RBaMi9dm17po9mVMZ0yJTPxLUFPPQeNPzNg7cL
tDYQTqSt5LAIf2iPlKRBEB/STsxKOtwEr0wCfjIdasMg6/dEqiR0XraClUAOageA
AZCFeSiT3JZbTict6IHBjjZVa7ymXhTucqLpsyukFnGRUFHX2pAX3lUEnjlPr1JV
iazNPAC9Kgb45BJd2HDbBTGF0sxI+bGOyVhYmTGUqz77qGMFfE7jInAFfxLYLpwN
a4kjt0cK8mAI5bBeSt/RsnAyhFMoCNIMyT11KBGVvTg5OkJdYaGiJ6YTPFW/luNa
wMKrWrZDqixUtIoSnCD4evzVFjx80G+edDuW9tX0PzKB9aMizc0wXqZ725msOoLM
nXglyYvGML3Y71qQUIG16tfZ64f2bPwR5H//Zf+v4OlFakQnLQDxOwpGO61nUKe1
6cYw44J36eZO09yoYuMWmIkE/tkyqvN4QvAR9ClvyCUMjN2D31a4fvZMC+ACDNuE
bqRr+4hGQatime0RbfSUD5eg1cAjpU5GEKVBLbxoVaRQn8FdKkMAEW8HJoxCB0a9
PVnal1f+EnoDOGXyS+TgHG1Q+zZlBQzi7/I6r0k880KSLQk9oKGsfm0NNYA/whi/
XQ7oXtTfeuiGIU/xn2pTP3bLZbTN7LTYcIzxclSpAjpQ9q2IC0yLq6LdeeqrZaeW
ZP6tP6TQtOyBr6qpuMzZSbPyDV0HZtI5899lfy4sduI1LWCIFywL+2KClxbiVyE5
z8n06xbeCJs8f24W1NGY7J7Hat+Xx9ibvcPmAfsvt6wL/21J6VpwzdWoJxwCx/iS
Fa2mbFnqvtOKUJubzCXmxqTiWx/J3C0WZDCUPpeSbYFaDK8QDjFqdEAf6AQMgf1l
W4w2sQBzztc77dNe8f3m5OEgCuVWLlsNx4t6sCMyIhU8X2f0eP7pakad6L1K5/7I
8bBJDG4UFWqtJqsYETlZbb/9xqM/GmTG/W6SJKALly9WNq9Bt9gONOWI7jUiyB/6
ViSvUNlbjwY2LrTd2UOK9VXMRXp+48G+DfKGTG8MxSuR2QN2Jj54ACPJdNzidbVK
l89JJdfSHqh29hC6dhOnLxsgn201ImcIVlObd2bcKvqW+VaFynumzQGRL7T3PcVd
vCwuiNeldDHewHx2VUdu8E1vskNmoonaHerwZZvFhv3jMaNOJp8fUMX8c3w8uR4p
Rse5LED+K63VUCPWwiMv1fYFjtAiLbre8WNOcqaYTAArBLjKPi4lfLMyrt49a6Un
jKoijJnZz3y79keMqIRFenvJ/Z5H1GJ1Ftvo3+FBDmCagdQx/p2pCoE602ZzMLx3
6riCGybtihMxRFxw8nCAQwsnTsG5rP87ChOPJRIasWoINMxQb2sElaCqBuwejz7x
fdedmxly7d8eA8M8VRldeMN0u8O7f34FC+wWqCv3M/c8N231YtMkui6sOG8fvg44
8TiiGAsydUVIuEmbTd6CaZMF9yL9crUHy2gKjrdfYB64ZLZS1QzTP17vCPfx/Ru7
LjFiqnia+3wWZVFUylVV8QzUUY9+DlJRczm5jU3jSZ/4pG+XUPBf3kWgdSmX9c0A
fiTLfswHcFU75dw8mLC7P71bR4aX5SKM8pFs7iGDAeEMhIFJaOrAe4hVW8o+YhMH
TUKBtmQwaFdJ3TgMJafU86UhY7BBjSl68ZOEMNp+vjtMa+r07DLD5RQQDm1eqa7D
KtlI59dIe75ohZEl0Pkpi2hjlkenLgngfXh6iAnm6tCUwnBxs1T8fXXpyk/vGexm
6lX5zj5loKfvSPFyedr/owcj3aSA883LDoc31S4PPUfnvkiej7hChDf5pJajVIUt
tVg0f5u96CYXJEfWpPyJ2Tm6jyPSa6r3STXTsYkF1rIItu6iuBaWrczfoHPoNVWx
2DVUVQYMZEY9HzrXKY9knMXk2feDF/LuGFmJDLqwdB7GEIuvfSO2Rm9lYKjLrKNo
DYctd2P/uU5XmsjZ07UobByGwBayDwEs+LFqQcUh8zJTvflF7H5WsiYYWLF6Qauj
hc4Ip3H8t1WfYqHDmgm0aU87Zn5vp/cQpg1ZFDJB5VNcblTb5GLmmRrbBVIO9Aq6
mpGX+45JXXnPJkBgduwkAY5fl/KxbMFe7WCSY5fJVUegJu6yDTCfLzGYaETEznbo
QIO57oe55wFiyjTn04v8Id9wbFhn2Yv3HIjmBVd5PlJeihc+JuKdxkYC/iHYqIUf
/wnBgqYYsvNiQYB8W8hv/4evTTEqLttG8xlnKazcrPYbUSqyCYAvaQSO8Yx9diY9
XeAjnOvPAcGb0m397MlenGptKbtP6nL8CZeny2fQl19K4lp/ySenKU6vZSib6jc1
30j84a+OHe77K7RgYAmCisqT+tsY2u3a408dNY9QtsaNwewBFgP3jlNaWr21EGVI
Az64x8lqbtjZ7gF/I0CNwgvjJElvPw7nxqm3xAvv7WsJ8ypVtKTgSDGabUT0ZQuh
bxJfDZsz5m/Kk7nGPBVv3tE16f9LF35biDWMl6IBcKiuy4BBh5WdjHIEEkVbALYm
vFJZo0Xmbmd0AfrUXP7hanB22gh2BhlxzfU1Cjjj8qbBw7YIQ/TSAI7hRTilPfc7
2BmhiNF4sJdWSK+qQTYSaSms3UCSSnmGD7xKk7OrHWkRmT2o7aMLS3kp7KF+6DdQ
qEdyfK8wrdiQM1Xx1eTtiZcR84EdW2nzIV7B3Ea9mi02mvyTojngvIzPBqh3S4Be
94Q5M0x9DUuTn69BknmpwWJCp1PQqYyAwnO825cZtx5G2/n7epN5hqyvnOYgcc1G
glDSfFa6XCWzB9/scsfK0davjmVMoQb6QpcmvQwcTidE+yPTa2G3V576GDj/up0y
d9nWTIgtz+wbp1mHPNVERaZputuXoaFbHGYrt6VluG7EEq6S6BGzOyi2uJS7f5Lb
wogF3Zuuw20o0jHIyvXlACRJJeUd+TxVLRCiLbPten0o571JtpWcdH+F502WwiC9
B/B2CAITeRodrVLDr4Ikt5nfgEqxGbBNpayso25HgXnuTPScU+jowBKI/AkP5YaR
LG2r91eMRdJWT5rOgM942ybfkjCSoZOTzIzs7UdfvjOJrMX/B64FgJg7SfZmg6o6
WvHwhh0Mw+mnc+vN3+h4tebcnmagu7oYlvCm969CTPo5UmPCzz8cfeZoLjwzWgiS
79kZznw4Oz0sVlKBBXbyRD+uw4j3jlZ10UThho1fFQW2wRpVZyLLaxGP8l08MMw5
mQ2S5uXXqLimrB/tQzRzg8eD1RNs4FLogXd7Nl23VWbYVz6rBYISBwRNVpj+gFah
CIBFDLBNZdfKQoUFrxG3z/BPFw4QDyVBxENB6pz/CURSCST8b804NEN8kJ8vjNtl
gFLnH/klFUQel5vNnpCl06Xf3c40pUmzEeP/CeLQP9UHXec9H2QLAU3NsFod+ozC
3axW1effPnPpn1MVetRSYvlKyFuFCSqVTonI8sA6+cDUNlW2q57c1iZFT6auxU0a
KsA/FkLUuuS/bR3eiX4Im4OGzaJkOQ2fX+mRU4OJyln43p1ZxxpfvikLgPBzWl94
OisGx52Y2HdiuhoHNOrK1x1EBygXM7ihvAOxhnsqrBWAulawaay+z1mEWYLu48bp
FKpA80ZqEcAPiNOB9wjTgAMOvcszqU9GQuij7+v0Ovee8GHHk5pYI1PSwTeVM0fh
lhurkxktAicaFjT7A16qGaBYcr1c3kaX3Qe6IyfpqWNQCsYVFLKSY1tU5+8GBhRL
WD8PUBokJoPh85BFMsn/ROpLeX0Cwt3RCd+iqNk1sgKPV5zF1sMIXVFDp1m2nQVE
wm4Lr+IOk1YOWqFIUosRksX7SgfC+YzKt9otMu1Dnv9BCI8MeQzXyuJj+e0PCq2V
YVC8l0OLmVzpXN2l2iSJLI9Y89a/1QBOmQ+qXsm+UpAFB2T8A3/7r6OmHWJJ+G7T
26phgg/RPE2t/hrfKhlqRFOLiUYG2I/+Sz5o8c1bAWJ9rmrwaO+DD6RVPv4w0xrh
3JQLe5G+Am+YOl4x4G2VIoh3kv0uy0QacBzXiO87iA67NLygH7yQiojSFzBbcdmg
ZfhxGtTlXMu8LkUz5cU1QNWuK0TTU/yEBs7/csADzFDrEn56YTGWHLBeSk9ZJy85
qMthegKDnyvxBlN9o6/CI4QLmJGMCUSVn6Usq9MMgnwVZMk5n+9uQfJgxNB5HksT
ytfe0je3OCntavtUCJ9McrVGEpKUP3/BuxZmvZK+Dk+5iszjlxq8RMFo+HC6RIa1
PjeczZW00jCb30p9BjuWApW0RBB4ExjoKSBXjHA/9/iWVpXh9uLYDmjM1EHMxmV+
xXYhhTzPeXK2aIJ8wtFiDHqtYSDEqRQdYuVhBS1PCEY6iW7vfQWLYJ9Xuxxc4egV
x+WuijcCFE6M96e9C4noI1T48KcXZa5jaGdvEFXeVKHNXHn5UW+AhwSrJ059ex9Y
AIELEE09jT7/t/DOwjH2fre8hRHyMVVexvbzK235TLzRzCw/IEAHpl3qMc4rRBIK
+rmsLtjZcRN7ZYiNV8HADqiMF+s7KXvK4U/qvSo/He/QGlW6gFHs160EKuVrmxTL
jxBXX1UvdAsqS7fJaPQZ7Sg7RVhFLMj8XUWt65GWxH/lWCcERmPmcr8Xc985kHuA
EAmwTk6+MiTxQXH1d/0y3lbLOxshA7D4quOsAkGKddSbpc5y1q+/fzAAdvPypXKv
kfq6euHeUgEkFs9ltMbAecWJtj5q2xCX8tDmQRME+ybKGG6rmC6bl8ua0iSu0k5w
BHSdEea3YYGB0b2Zw1maSbaKWQJ96d4TEPOKuFfUrejtsz/Z/hpurt8rEPvQkT0b
SQLCkEpKQNSM9+uDCJ9W715fr6nzjCOebP9Ax9Xt2N+UQSO16Zdd7255kbHka8Wi
WwGCERz9h+vwJkfkTZOQ3alKqrC2AmPoeNEvh5bP36tTrCkMBIAZ5gCqkUKZnq8e
vaVLzP7tocDejl7yrpeQdeWB4JYwhg+ns95yJYkdalS/+9I8y03zIKJfccEN7Tce
dokkMVsQeysFmNQI8t+rkQOoH/5NKA8fSkKA5f7uVTYj425mar6NhPuTcBd7Fr3K
p+2m7qPPpQX3xsSC+BHLPlp7TCAx6f/fY42ZH9jDqNv0gBJgg0f5MxknE4AAg3PM
/hlJHPZaX+pF3mbCT8ifCw/INAA+EOBMTWYK1K+0FXLbWaNr/8S/p2mO3zXEg/cJ
8gDELqEA/SEmB7AULstrSuyMxkcOkt5RYM5DlEs69baCq1RFKAfAkVcHEMKNlKlE
efC1ttWhJF7gk+UzwmkWGSzgXb1M03VKfk/5pZEovZv9Y9fuAhzuqVCcMxybWRXv
PHpGiA6M1i/ARSIC0Blr0oLv+fMqgJKctCIYVaMlgRfGxNHHrMETmRWwh8G8ExPs
Jn+pCGxVb2aVpFCAeb+tOZC7ci9GpfDL1JgYbEG/pUaNT0Y3osYVkI8Rxa58JDUJ
eYm92CKEUJ8CrvEwHgnSGi4R5hNQA27uXEOdOtAgmCys1BhRC0DF9rtOYuNylxIx
Ug3qkDAZ8zCd6R5Vz31iyX/KbVFpmj1NP21KiHe38/glhOYJ9dsFnyIe+fRTqIp0
6THEPHTF3MeNl2f3d4S4VB9D8pUaKJFdh7ndTkHxESOmNN6LxN5S5tWjFglItQIL
HbMQWBP8zHCqAehajYPDbCqqtRcG8mAQgaLFyD6XkLkmKV2G0SBVCns0B3/3Enqt
qifmcdMlc1N1Ab/igbLJ1X9ChjFVPALG8qNVU2jGgDCp8Ac9UAGpuCs0y0fz9l8m
ayKauLQ1XG9eN8TcWTw04dt89PcNB/IL81SoNxKEvVWpDKaCLRVQcaia0ntU8t3J
2M4ZjbC41DBzuOkVo5E2fL+ssLcHNlnWK/6XEE6G07HAgz0vF26mkccTX1M5TVnI
Pa3Cu3wceY61IW4KKeE/gi99dpgO5YgVtlLYfRD+bVoGDSkq1eEBmpVCNTLZK9Ze
ec4eRYVWxvdUUTnQS3JHVukJMfDkjvBgsu0ROHp4UIkCpK2qP4nncJfsrj9tn/os
5fq85y8oyFSEIWRD0+CS6kreHFBdbuTN/MhmaegT+f43ZWrd3iv70uaJE3bthqLh
ufSPXPh1vmQN1vPyU7flETZmh8CoWBF8h6R5g7ZWOu4KMVZbhj1YGFSx3h7DDKus
9WnJXI0Svqmxp44d6tBX4ZUMJUTiMdWgis5VC7i70ywyzjqODjQf3ONxQ5T+xa2z
nXK7qw1ruDIi7nKbexCNpfswSR260qG9OviqMS5NyrcvgdEgQuyyngF/ZPsxzeBV
KcHaWbfcvtEHs9B+vg8Tr/NIXmsS6nizpWCXdaH0fJ8h5krsU3bNgE8mEXZpz6Ow
KuWqOLbBNYETJ1wiC5KzhqOFKjEzmKydAG6Isqn9Ggk4MlboxsB4RmfOwHNZRlGd
Z+e9Yg5Ih/v+6rJ9Qw/NIRtkLnDkuhGgrL+zraoTl13i5rbvZcZXGPCb2esFrbXK
hH7wD53UE0jzWl8sYfNzAv8RnyZLDFwKvNsk7ZW+LeGLEMQrqHC4n8O0We6dNGzF
kyycsUmJeQiRJzWMYE542uF+SoWQ69COU0bSsu+d+rTEdkXsKd0jj/FCJ517v+kD
78OC4Ee05iqGK25CzHPztRGhQP2oUpUZCD1rRFrruKvOL+GZKEvNSV1HtuRItBLT
dIX361Z32miZIhlubAXCTLcSkhiaNaC3kddJmk5Wor7HyryxKlXvah085V8ETofG
Z9l9lRU08ItRxggcSuMT2cy0NjS5Kcrkv0urwu77IJX/ZokaLs7qvy+iR7qgoMdR
qmCMT/oWkVNhd2yvyKvoeo+Vj+dqbuFdzwVOFSsWPLI+SAVx66jTVrwRi1o7W95d
i9/oyXCuA2yQ6zLYMLIvO1OEN4EdSrgpweJZUjUkcjUQScIDM54c9B+G0tuAK8DK
QOFAbQ3tn0Y09nB+VqNvxwoJscYw4DPKjvZvb41tskqwsz/Mrj6HPLhRhLeT6nD7
mXZxSgWGFtwahxsnBl9emxpmZL6qP03amAKaPRsmVlctrDdETS4yN2E7vMBmXswo
4vVXz1DtsqGGmwr6YC1Ujadl836b3E476DGoHVf9bXi+gkFYanMCjjZv9vsCP2fT
PVNLKy7kQIROA9ZPP01RM2y1OAf8FBo86gr8ji9Yvq8BzPxHR5xyPbstJklam3js
91AL7msVkwBVbmO/OypLNN5pKaHBqhxdbO/LbN82qldnpCOuQ4cdeFgnlGRdnIak
utYRFi7kXcy9G/c00J6xPZiNNLedGlD88aVh67Diyl8KXdPCIddKo62aQ+j3/j7R
wbJxPhQfdL6v9Ych2w9N0DN3j1UFB2NnmDcJlpXEMSyKKi3c1hItLRX56aI16/HU
KqZh3JEFWURGA+dq06x0/XBFAwX0OZax2mR7Uw4IS/jZ+3uX/FOn7NW/AfpfF2zU
E4L+7L4l8dmP4qhCSUHfiowbNuTprA2quB4Z0fU+Mbzrrd4oshuF40PCa7Cz0ms/
exMAlok/ReBCip4g8o3jTNp7ps/gMBHvKz8McgyiB4p+MHB9KLuc31xI8Zest9Uu
XgRCk6Xwo4OTAP2cRwqiCnslP99fDdIceE58uPXk0h+1XPdoMUdDM6N1q/XVXqYq
uHvZ+yccKJ9GuTD5rezKw0dCsfRiBNCiB3td5YBi0HFx5ZLnGpxIRS74XyPaknDx
rrd6F9PI4tIHRnz3n7siqW/cGWdEIsy13MyVl5q4XjB07IjwmqsitXSv5B3XvG45
ZyGaKv/G7Dg/lf67fTpqjLiMfShfd2jefd1wjBjJ+kq1J0j0VDaA05O5p0pu+axW
eGQdZNbhOhUyXMy5iNgucCUL8gDR1Th4btA4BGl2a3aVlfnL6ehtGTKSQduJY7Eg
DyyXf3YHL+mrtX3EbXyT09pei99DFMS0TCY9CoBTx7pBIzIySdHfydyJViektHK+
JSZ1W61AOBnHANiG1zFG/KlnTySGUI2br/cpxOcB65cuRfGoOucPSsMPwnGTs3Uv
cTYKJFhxKA8gEw+6sOiW7AHIRgOOhoVSakVl1yZOkds3y7Xk8HwzpK2HQ3kLek/U
QEeR3ydlOGOs/ufuIjAhOwUgmKolsHFeyqY+Y7y14cMcJYFZwv46s3g9vDUX26PF
qCp1KHyMM03n6gkwvHGiS4tl+C6N3TI8gWj20auYRQmucNglCjQStY27i5Z6REz2
e8yotf6idnmS8UIG5OQq5mw9VVhSEBYb9HDe2DwFmogdwUEeVNN+Jz7WlNSFmbe7
2wsnpR4E8IrpihLA8vll0oDstd2EXevq3x8+U+2znmFdKA9UF7mNmtrANlUhC1PG
6HmS0Rv2S/vR7a0ApXVmhvSDxkOXKZdq1UsfXD5xA5HAVhwz52M1KDuG7mzWeH43
i0LpG3PFQfdCoZPfnKU/R9plvCZfcBaUBqLOuGb3OLsV0wC28drWq4ZPMTrDQaMX
GKAtBtDiUZpZ9i+hYFiII7Bhy1Y5JIDWxq0L9wL2a49g58pfUrYgfgqWOU0xXqBp
G+9iNOfSFD4++9QG8k2ITb/E0aq4u4Hbgb4yAve/Te+1qHWCujQaeLNjTPCT+6XX
EPZ8lVRlbSDOZO/Ts0c8j7AEzy6IVe7GWXIzCu+Uf+L/kTBnO29RpxnzusOldjor
BcwXzvwzUbxRqsmXySlkRkDjnhQDDVPhFWdHyHPUukEgVtpRt8lqTQJ4j0XBSk/C
GTnGI/x3klMBP2BiDM9GfBArughc2BFFud7v6FUCX31cz1/aG0SLM82UlihrpBKd
AC5/pF2AZRiMH1GwqpQwcLEwetfh9wgsZmFtNpFbGV4hS26BnMIYiKJ+NNHdXZGP
ehmOWgq+dMjrpTZcFruiPWoBHqSQ0ZK0GWwmGKNX6PXoTwUnpoXDbjZhwL4fJtWU
F7GlAzZ7TS5liuo5PmyUZIw3KbBO9FSo1SFCS7qalozQZ+lDmMXv7f11UyJjNGkw
2e4QkAI/WJlEzyb4SHQiGp89ssDqvuF0QDbsVhbspDrC1d8HRVTPHG67tH0wUekn
qn/aVuSWJdETxEIyR6LoRTnhEouoT6hddgvMO1CUE/0WWINTV8uG1fBZSwn1Cf7y
pofbigB/EuwnWnJLalDdJlh+wOUHXGpOqvfmhBFwHyVYjplGyiwX6giqLAMnp+6W
YwNY67pFRFO4IUWcM4UQSWU6l8ioBqYeretreomi24gKy52orB2embhBH3Tq9N9k
k+fdRvHiAHAZqvn/A0/c4utHgdO8QU68rM7R+zuwufgkt68LY+uAHLPPfHzUow73
WIpZLygdQKMNpGw2aQyjx9dF6cQLjQ6fIzWYD3zgjVyiFsEKMrtpsA8JvOq1SoZl
OHIZZvgacHz0O1GAb3/fTehg7ZTYPu85jYhKu9oKzmgEcfoHN64Et2bMmEAzAlE9
rdHVi9wW9u1euoQ+BMhYmZ09MyQErW0CVcu/flJxQlvVL61oD8+HDoom5W2g/1+L
7OH7lxg5m0bYLxFNbI7E89k7/LxVinFxkr0HpbTKr9aiScF6nxDvTT/tZhkRl7y0
ou8pry6SoNJegzXjFZfiovGlKH4CQHcMNNssV/b6ylwbMoS7q23CSC0UiN+liwb2
8KfnCuX9ks1mfZAImZp9FGVLFEbnQiesYSJSd9543ukHh9X3gCj+2cV0MAplYFsN
HTlq0Mf8f5FKrRQC46/gn+75S8W/l6lXN8Td2C3k1bqMPpMjBLyGlt0sOChPmii4
dy9PvNm018NQbJlurr3/sTWkIqMbBKcNnbbC1+OUmBcWIpgTRv6Pi438HWbfuu+r
paJmRkLZjJy/bZyObeeaf05WPAYDXiwDOc4BLGel9E4vbdkUulQBoTnuwlsc0L52
z9CWrJRcMJ+mz5piyURGMZx9dsMvjh+DK1CHBbXIou0gecgBA6c/+7SjVhlAqww9
Pp4FoKn72yo/DfDTgSo5DztyFFuekwOXBZgJq4bZm30ILVdPPp9hwi7WWKSMX/HR
2uSsiAP1h1R4lEYXc9ZH8m6QLdvLstP4QgmSEY1SZUgGJFpUp8triVB9JlDcd/a4
2EYzF52QQBvg9sYHhlaNYewiVoA3aHpaDmqiGhwtp54S0pCheAwUTQ4w1YBAjoJR
CWivcMVzU3Lh2MjJIMNJamsQemwL+rRDLAzWPFOkkwxJYIXzKEAUm9vaIxSMhKFq
oPRBPPOJiuYot7cMlLqPsTtBP7c93rzcmqBW42NpThtPAMKFstJsGXCLlzjZF5VH
JRfSuiyIPbN0kFF6xCHCdSP7gf5ybP0ZSlQ9iwLKio//gEIF+5zzMih2GUDPP/tT
UzVlQKW1g8hHFelpe8DHz6fgh5a0Dz7PiuZdIC/W5ovPfP2VrWplt8KhoMotXNT7
ae/x0iv998qJH2SU1/QwwLT2RG/JHPO7qkHPS04UAOr9L+QaQ+YWNj4BDXMNYlal
YHpiv3gdL5WRodPdpH8BGfHueg4A+KBjjQrdVIKB3ufWoiNUye8MhWW3CJYmqGV1
5FhpzuZMt2e109UVCkyVHKWUfsW2c5F9Z32sgJTI7QYhavkxFxzs1OQV+UPVRGue
McPzeemp1bXFQ8gPUTTMmjZSqHUq+yipXSCKECsxZ3EwTo3CF2OdhpG7q22Ocpwc
JXFHCx3k60ao2DgJ6MHIcvX32TFyCO3V2kGaLXhV3HeejHCYJ94s0dcMWynjOZOJ
C+iGOHNEXUfEfkmbPO1ClwZ+mQWdFWcLfKOLTIa5u9aJ36dYZqLAePnnHokfuCxV
B3Q3jMC4iQg8+BLj70YcsMo19LvcjJ6deyf3E8kGc3ho6DmO3X9glPl1r1djlNAH
9zYC0IadMMVF8BrebQDkOCEjU2orA83y6jIaqc8Knrlr6uyYZl8jSb6xOZrKdmN9
J/ILWZuY6+KhDfNAgjfaboS5j4TwWHbUVsWOLKIjnRHs2FgF/gvEx+pENo61NtZ1
bmZfTAkJ+fudf+nsTPwD6j45IEYys7y9AXXvzK3d3OLFNmbKwFC3MRHXIbAp5AdN
xe/RUE9WypyMUdWwWY2P4NUxSqrbqP5WljtJohWHGHd0cDmwcCwL6mvojLU1IyXA
uLEDxxB6lGqnrMmrz5Eu0AJtz5D3KfMrEkS/0qOxSmTHZgln4kFBds8BnMsz7vWE
FFii/VxVaNKbvfxga7b+mhxAOKH95BaF9WsOr+CPVasbgGf0wgsC9wwKK9A4Dl/Q
zo647MEQXLUPNs8YHyLSAEHbT2mlq22H3N5scO76JELXCA6VwLKBYsS3VYwkTedj
YGxX/+JYNKv39afS5i8WiJAE9dbzSwQx/oa2RQXkGzofJf9M+ffQU7Ay62N+HjDZ
pddxjOA5FJFMJ/lT3zn7hXWtktXUucwUIk3wxvYMt5jvP5zJ8suNeoXcD8Ly3ACe
bsdKCS6comkUXeLEOhKB+yu5j9vcUQyGpLLyfu9x87TQUwTA+R9uahmZnXNPdYaX
5aY1iVN/8f4c05oIzgqmFDboZ8TUN+RT1haiJWSjNS6FLBjS1izCsJHdTcJyfWKU
rYwmSVONWyFhrLI4FEVCJyBvG3ZwiCGda5qPAztPraC02HjwnmMIBzwCqEc5xMPZ
VDY2luCWxPGd8jQX0swlio3UsnIaEc7+d9tGzsuvcA4tonmopBatjML8d+i5QwkM
dfDGsN68seiUBiBsGx3p2Pmv226FeOlZZr6e3DcGGyxz9Tu0oPn44NaZZxBIHas7
nHzvPvfplLFu5ymyli519dYuCWDO6u9YFiJOlc3RZcwonKuw9VFd21svjNEjAbZZ
v40h+c+5wcXHDUXQJ/GuDTO7jJg9mxY4wRFtFA2QAMsp5FmYn7mAc9gquANibsEg
7K0uMNq6Yut3t+7isLttw1wdbsU7c3aNTFl3Umj7mwNFNeWRknvzAQqg1XHNoQyR
eZc29CFFsCeVacEwUjd4S1UolxZqoQsQRTetQ3FhLNz837gebzsHOrQriO9kPddp
ii5c/V7AMaU4lMbimTR+Qur3V1+uCOKAkbaz1OJ1Rrhg52Oq0FLg+DWVc8eWVziT
og4E2byr3WznqqynCGWwMRgGn+6lfIktZwBHAkkN6TxjtkDiqNRFTYpLBfVcCPR9
PCMYbPOlPkazuIAZ/6CsOR0qgQUvwWrXpbXNHEHMkEMDFCzWaxWrvIkiNxGO0dVw
AO2z/8yTJ4VBqkivDaKKdRFtrUFEJXJIBg/rsP7uKkK3V8kPvyPslJDs8BkWDwjV
9X/J5nfS+26+62MDE/pLE0AcLGO3WRvBO18pGs4tLZjf+o4T+kHEy7EvrIW36KHT
G0ueudDhXZ+Tg5FI+iwVnXhf6/xN3XfAwFjlgmrwhl5b4nDca6G8Y6/UytN4ZjF0
13KiW9H9tl/pnIsy4k4dCXZErndStzsU07xrceb2GfZi6KzUp2vxhGoRDULhJHuS
SRtDzzOJaGUvDFLxxeynz1fRtWf4QuIOHtSbWDaVFqozb5kTUZolyc1LFtFT8XkC
BMo/iwpV7BGOLyBdnBUnMaG/PL2LoAnLReKhSlJRUWsg6y5md9XTHip1kW1BaFwH
Ji8c4j0MTFqxHAG6ck9X3ov3mDLVvoRc3JIYxXVBtnsGvveeYapGc2JPQdvp9I8Q
GXN/y4BwnZD388gvZfA0QjQv7qEBkArrxVYYsQZ3MDvNcvhn5ZFTj/C+m9NnFT2y
qCz+22dB8z+ugxaQa3/I5gcPRfdkLd/kyPjOhynM3UMrwCORJasiSbtEl/OtbdM8
zaVi//9dkfDAQngRHKh6cqsSZQR9qLHzWZ+k40fprGloORSbETLic90g3ybP56wO
wcTQeWtKQ8q56PO49u202gVV4Y0YrpbaX3SH2ak07kFXdZ5+tyNV9WFrsAuKAIVl
nv3lIGc2O+1Px/mCym0Gde498rIMRcR4wvt0f5hMUGVYbGLjGEqnMmRp32hDhpKV
goCSPieFRobGFHEda4ucffyxh3sO19TjvFjs4e06ld0FPjR9oljBPjY/eUIe5ABA
wb4yVRYuvi9Yyr2llPUCtE+YpQsSS12i3IttwXGIyTDj74aomMXtCvF9h3m9qBqf
agqkTE8IElfK4ehaPVuCGJgGTVLy4loFVkxKSi0smrg2bGPMkDm+cVJVNFhoCxBW
x7EvlXy2VLNGzyUDcPDIKxcMDaaAzbhpd36uj14rORhELwlcemnhB1h3RaGsJSdI
ea71nmCHDmQpwAje3y6nLUVUyuYXa9Jy7MnFar+Zu7Qo0MVGt6LQAPZsQu7aaH/i
jqFH1pxqXf7U3I7DhESx1c9JfulD+wbIYlxh0PZRFWSKJCJknKGftAh5izfRppIy
dQxT0Yo4NABEQFxycH9VNbmPrjgiz9MyyZggUQ1lphBYODDmSEQBmBS2oCA9DRZf
74rle9W8vaVebkuLT5Y4iK1c5jehcuKXUynyLY75pIGpq5Xi2wHoT7qVJM9rYPPt
196vxjT64e8X7Pea20DxwvvLClqCleIeSIHA2F5YBfJsBkBnJ4t5aE525bmgiR0v
rFffQBUkCF0rIAshantxszAT3BPBbv4swSI++bKJLf8FrQF1ZmTSFkqXvzbJGP2Y
OvxRH9GYXv7AzJ9BJNS8sa+J1f7IfT8xGOP5Y0I+OzFKb3DishpeEDYftZOQzyvG
C5XAVbZ3kFSALuM1u5pytjw3KSURIz8IJD8ZMLsDNO1Qp2Jkf1dmFpWrKsPaoRGQ
+IJUjPJ/zc71rjIi+p0cn+EfDLpYR6RFnWEDEjzVJuy6R4lkyFz1KVN5GsqCKOSQ
073KOINlB3z9ps4HT0YP6mVb6tYCMiK9IEhAEkUcUyBE3Hr2GURRGHtg7LYCXFqy
WvwLlCD5rqGbvFk88vH6c4oVbZzUy7RGzKeJ3buJVE7Yna1FiS0G2I+UfpWHHzOZ
PLNJvqJ0viegDrdpkTAVIDrevBlsD37xbayORIqLInOSQ/QccqlVikRufTQ+aGoC
MSlx+UEOSLHuT/NqpwbXh3d+Y+bOpgt24b6yKAz2rI0vftZutn8eZ5j3MvhsKdCu
CWnpTwHhOGOEN2dUO9wLA3Dk7CYeyNAwovxnN5RxcHlnIWVqo7HTEMpUXHeNk7w2
vqcjbbTZxbPGBa+fAlssmmED6V03YGE61MPKv/a3j+fKUDMJ7GVaKfKB22L7bsMr
2nyms6fnl9QzMWOsPdKrKypfmDRsHDqnUNJgxcrYIspVQlqVMK0pjCMx21ok12Yd
KXtGneWRAEP3XRr9Nenm6+Z7IiMyENTfH/OVL9kc1Qj0EfKZO0U3TeXaqqYbIvCD
gynlFl443Yw5NvrG0WzzHfmMP7PLyhFioC7x5D5+Gc7ETy3HeVyrHKrrw3A0TWzp
/UvHrjR90YDIbwUU62oPk7HCD68YIOJoG1Ib2/6+uasUBs+uGg7/BhivRC5kwEaL
EnU8zyDoZiS5CFnDLwyxAjDSiawaqMrlx2ele2JjzxEFpFSBKXOpvBORSaVwef5l
2ZvfuPf3HJzE0aO+dnTUz7O+CuZ7E/MTnrcgmkDdE9Y9Uoy6CNbArQ7WwhN3mg0V
5DnEbJifo5YhmaT9jrx7PDKgFXUxRAizGEKYHth8DL/Zv72dyHaH9h58thEoWq/5
U78nxo+8KyxMI/TBShJxW2NZy31zaVw/0RrV9yKQZE9z/bDXdDYogeiul7ytLHiO
BF9ApwYZSUvLYx2eG4q3lZuq2WY9p194dEwUAxmb+tQWtrvQ1+0nfTspim/eAOQl
D5MG/4wf46dx17aOcbwlsDyqrKQfNk2dXGZD+DMMT0LocBZS67XCItvlHCkSGNVU
Xm31MIeHS0E7HZe/tzDvmif23oModUgkbJah+uDrZIIPCET70BEga9QlOEOJUr4N
/eitD8h69Xj4uRU6KE3vtsaeiakUPlciFMp5eQApLuWI0jsTIjZuRBd5Sf8IvZlg
hmPVFtRTPMmGNJG/2tUkLXPUa9+glIWCYkobN2XOnYsEEdY0TAed/KCHsz2Sm1vN
tLw9HNqNXRQJ2VywjFj3THD7nqGJNf/sBB1tJ9vF8DBEMeC1nDT0zQbAUogCQvfG
VjF669qqdtt9o0Y4CaD3EE0E68sTwLGnTy8TsrQEOjvQXkbL528l6RWzERSYe7Lv
0WBZNn1t0YIxoDkJmE1MLkin22dD7G4K9ELMvyn6mUUlN7Y65B/LfHGRN12O7jsV
YTVFyQlX5PgLn4YgBQcrnMqa3HIUruCO4CY7NAvZ+T73tCwkdy7cEknSTLYheyYv
2b7wsbQGih+c26oBz9eMgZtG2R3OH8OgvSjMne1N4EPq7OVumIjgyP/cBkDVSdd8
pPxA15TpeXmXcF2+RE9hGhRRvip1NGkxT2KiowJKmoIXDTi6HQkXM5Y5u2Y/kwo9
Jm3QGy2zv7dFOq+xWrGZsnAasl3Sk9wQOEZgvjTTvRHbynNx4AjXfVkiQ26a3cKD
Mmqn800GZM7LDZ89MaukwMaJhYccnbGiumt+Sa3OZMBEVs2DRAU3SpSCljvCAvNT
U+yHIwTHFuyQS4fQhZDFsn/gOkcWfOfNb4+3M9l3HBGOQw1CWEYeGlA1YsYyr2jk
pab2PCZ69bhI4oJ1HTXXwqHxSbj5mQqrAQT780/XjWrkOdUvfnoqCOj8n6yvKrE4
xme3Psq+xp7K/mF+t+r1CBKHx1YbpbZnz/E19vak4awy+QC7AOQQaJDmzy3nxhs8
8Elep8ZVw2G6K0+hgTXEqpd7dkY0eyzWPEM0woP+D36G4vdrmiVph865lc6/2hiV
OH0zBGnRFepFaEb1KJfosnfKd3ybmHlkJ9/hxJt7SXpsr3a4OIFpB8ssaXyIyGKu
f3DxVdh7CGKNufDPCLnzpfTusC20GCb7NsBHVywBYu2bsDC51m0Je/P3KXHq0UHm
EzddhjfZ0Xbyp1I2AQa/rm6lXfDpdVszrdIKNOzWoepOcOc97JeOg8R34WvAnKVt
GGXPcNqNHHhe7vFERjS5+Yx3Rd9CQCsecUMsiL5O//llEMw78gGzUiSGNuoNFKu0
6b9v4CIfsGjHhkWIW+jFUVCUrMQdGFtn8EddugjTZeJkBG5Aw8/mwr7CZaRW5WyZ
CUWC3eDwrjjrjrA0Y+6CWdTrZaecB5Q9t7KWpmhNk5ZBvfQK352/UlCq0I38V0S+
d9WuNKWgp+9re9TjX98Gl649z4VuQZQi0LRo96mo0+KXOG2+Lyxx+sGM0vC4D8k5
eWybh0iiE9c3wisVF9hZNnV3tUkbkiy+vt+HwH/s29iTMnwGMy2LN8fX2MfXw7aa
+Ckepuc8PZLQ1sOEo/jHVccXulqRT5/svxCzTGWdUX0uFRLz7y7m9nPFhF24/M1t
+ddGqKfOJvjMrHFEsnvknCEmf8OWGF5eFLZObJ2wbfI07A1/FZSPDRKWhK9Q1TrX
wLMLCG8tJ8kz8/KChzw4OYUouyBmr0bXK1Q2RmXC3QMkVgLFCwfta+KvCMxMXqfV
3QqUuSyS+MtJnRiodGfi/g6nAKp5wiUdqRJT7DaQTCriXi3w0D0wnq20mc7lEoyG
FivoEnhGFxCzsaMWuYVnDcecoT0fOcHB88HIs4mHap7B0b5SiCqsQSX8BxRPuJxH
HjaYLfnkGG0zu8uDxVjC1zmj2RJZAQ1E//ot7/8i/EuK6/EymnttKhRFu6by7cw2
zL08jTLHkDxreTUTXJVUeW0ZJcv5/r76vCbvu7fyIDLGk/H9M0erp7cVTZa+gre9
OpuYyEHlJzmR0Z/zNMxkya6By/8RZ3DdC/1V0vBiNjGoZ7kX6VLYOEldod0Ufohp
b9xIh814FL7TcO66O6CytZO9LM9oRSgDCt6KaFdCsLhpsa4+HfsN6G9AgBwl0ekN
/D5oTiscuHZPYyQUkaxEpI2otCd/UzzhMv2j1v18iC2jDY+GSgynpV0YT5kEabo6
IrFIBNoVOHgoT6hrv/5F52T2B1k/INHYi+rNmXPNJ/kxeHP0Uz+ujH21wwpYxaTn
UKZTF+TsO++OCrDpHfQJumCWx8KulI0DAQ9VaKWLeNvfJaZ/6VGS361Akux5r+Oh
zm05W469bx8f13WdkdMExmAUyay8drJBW+HIg8egRv6eq066eVfZwYRUVNQnEdfd
MBOd3lADwshpNKROQftqUtpgKnkZ4giddG8l5iPJP1ibLurdNwu9QeMI83Wo0SbA
Tp9XCDka9sj0Me7yoAwXqO5nnDIKi4haU88wJEtIm5cNPPAP0MiXcU/UCBrOE9Mo
bfmDX1wD3eHpT2XeyZQjRJ3XzYQN4B2rpSXrvfx5lZS+vKPqR3V+IsXeDrR0b9QO
XmwueoJWUFIISyakFfK2g1jZwhOQvCuvEs2GzN8djj6TdyPI4/GW796ENDU7x0cr
Gj/mYiOh8rG4NeSOzVjePSR6H+LMXvSfpr32bklAldGEN5M8REHUy61lbdfMKkZE
jws5h1s/OR/Zicu9xcmLOnePW9KiPGG7pgc8Lgkq9decVK3rxdf8n0CMUnffjB58
RgUWQ8wFb7T52eb3uj2pcuhXoDQdULCsDlM2VhU+z23447gj0ZXbyR8RBxwckCaa
eImwr9ZDDC5yR7/S04UjNiYrC2OA05i9SQM0Zs2x9qj9cDL1Zh7CHnMsbeqTOALG
/59ov08wp6Aa07ku2XUc7/vIhmEYtMepf832dMLnlqXYBgWzhdIlJHB3Wv3VD5z+
Ifs3xJF82womdhLHyGnaN8UjzR9hTyk2rwEtAvaxI1CJp37m28blWI9TKtJNoZ6G
zu9/dasnBXovOcIqD/QulqlzPKKLn2j6LIEYkWDn8HDet8PbTdCgRm3FgdrBa3H5
I+4Wa2PeOO6aJiBXhxDOgUexpcws2OZMcGD89DMk8AWyS4d9rMC5/9SiMO1BlCF0
6+qwY0pRaN93FTOMAsz87jSXZq7yZcK1hnTlHO9DMdJs6BXePUVniJsTpWFrVr77
Ft6NwJfEMNWxcvGnpNd6N6t59YzfQpTP/maIiIzkSlAq+/1gTPZ15okXmB1MmnyN
B7aY2vXYDvBfLPD6/FG5xme/lNz7QaVl+S1A3GsvDSSv7TkzyyDi2ChLybsc/s1H
Nf2M9cpPlNGPV5+g5r/C2ux02UqrXEyhXNzmkUBYv9D3LpdBBHqRwJBTy/zBZ67J
aQYbayTlr9fwNUi+CvrUL7Dky28UK0JtOYnVZmfUgg2yVKiho8ezsHzx5wxF1Xqn
wn9a9Z05v88pvVQZjbS1SnQKp/OwfbJ/aXvvOONwT+Nh5XgrbLgvOQQjabk3fRxz
C4x/r/QYbneWLBPaLdSbjezenCOqoBx5rhIji0Z/3J/3NiBUpTxGl0ggHkxkGWVv
vBUZgQO7IpHX9wCi4I6nmq4a66B5nq5aSPId/m5b5E+Yo443YRsDYVHVIRHzFcc3
8sJHuiEfeDuRLMX4+sAFF9HKG1Cilq7WIc79jJCUUqzlrd8kEQ9f/cuzqs4M6jBR
wsGubPiBFeDJflrYTDRdhJn17eFQhV5ykwIbX0D0HSmHvlhOzbWbRAv6+txk7tfY
VDNABXTA80XSmYr8Sr/rg6RFDexPbgazuCyP/IKED8N03FZsaX37P7DBSKYSnoU5
VdPu+QFDhwpoxATFyoA94tvk6ofBOnZTuJqIFBjqFsW+mawbvT9Lf4IaT4MsJRdE
BrS+3OHnzMlFpiZPAwmpG3kA1gYK988EwnuPUuIcGn5l7wo9CQS/JfLjvziFMY53
CTqzFhvRkmlPzAV8+ZsoMYgtA7Y/VT4SpyTIJcdqEVArNU+Z1UfGIKvNLLVyMgAH
Lcz5tDIfleAkCWgdeuqDaLirqLRQ0uh/Na5naRb+bpALX5AzjUNvVJSU27u6I/aq
hDC3yjZ5Bu9R+4lnX7l3Feusms58000q5se/oGOPOT3WhWTGLTDLDG49ZGhs+NhV
b1wVWdXgnyj1DYH0NbobuwUHYgxXhTkbgTUubPHGQ90Ym1WFNHvVEF1rDfOoxidy
NllRQFSDKQmCTowhPdP3y76yx+CVbDxXPugdqOxgJlbiWXnX56uN2iu60A8VSK1v
hYgWJh6w48yRYNNT1jj4c4dSt+z4ukJg7JYKTz3Cghn2U2UNgZjkhr8T3ZzlCrpU
Nu5FGO3kh7gCzJqzgXJzCGmBwMlhaZeDnWqzlczNsiqU3z5lJxm1uWhs8HMRGlTJ
WdIu1w2KoH64x/adC3ZNBjk/7mQV4KjaYdS9jocGjLYbiU7JuLyRFb9HmpXrFgel
crWweXywWqznDY/El42zzMyH7C1Vl62vIQXDzjWgdOvET+UaAgAuih/sHKC1WET7
E/jYtLbljpndD/X5kaw58jzUZwRsjZ1xLTcQ+JLsqgykT3zqAZl45RYpTHvgm8Oe
7ufScVUZXecxHXDuaMe6a5UY3uGfx5mvrjVCftHod3ern2N7V7Yn4fCud1CllgtB
Hzt8F16h+nU59mVr07JLG3ox0GZtYlxeVf4qjwBOMLlcbzmIY54ZYv9gnicyAzB3
2aViTHT6xmA6BYXCOfdjhI3fePDw8Uu93hWcPd8vi861Gdfz7fn46cw/P35qujhs
2BNhhSAt08fAapKFEhMggVPRS7bXHlP2OqRVR6uWOjjg+hNbQgRVh2dNNEgvumBV
HwG84ue0qzjMoEO0fer0zIwwRq+RFx8HkUXbud/kobl610HmQ/LWdjqs7nAvQzEc
rQeQAdtY17Y4ImEqwmpaZlHfeZ0nCPDXga3mfjUqY8zgbpvbdLeuq4VpwEqtUgP6
fbRU6F3Khz2yESXD8T05TfvKvBMqg72LiJgqXd7KFSeHjGXKUMpvwPIapXU3S1li
+i6RLroGqV6XswPSgruYJRvh7CkoO8uUNnX6UZ1ruVO/QLu4fAlN3jWTp4N2mQdq
iMFDAy4yDzw5DGdq4CW1lS3iF6Lo6yIkK4s4roz15P0wglxf4pc0Sf/SWh2SQrZb
wxQwhWVOCD1DweFMcwlPPwxNQzk04scdvDJJYSGwcmPdCQLmiVemcwUlsEbLz2KH
Xeg9yreR81BWyfw5zEXiy1nWl+c/3iCKi8IMz17bLZEiGd3fvX0LcXuoxhhiTa4/
Pn2/w9PiQdbf6LOxZdlsYpB4kOHYp0j+Cvn0VzWi3IDyuOOYtHCRJzroyt9Wv453
SlfcnE57isiNVYjuTiIdwXK0g0frq+8Oj/lo7FJIRRiDXlKiqKonAKl5GcZAYSp6
fkMZOYLs+6kTkgQyiztAuzVWZUFo9JmC34Idg9vc5z8kH6CIZHYTQHjTFxAYjgm6
tGs6q5RSzFRTPexVeWWwWCX3Ku9vO/aeQTPOuufEKOdYVjXqR9qXXRhfGcmhXmTw
U/IX+UxeDlLqT0SHcAfZT92hf8ju3JFwyCNGsXQuNG6cTpoORg1rbPXmN/R4bee2
Aj6HpiL/kksaGzbZdqhC84I+sXve1+liC3X3swB1lp8jpj44amN5Ex+6xBM8pDMJ
zj8MZ2m7/Sv3Rq528avBe7gOKN8f594kJC+bWm/luIlIkBReV1V2oUJ/6wpVj3tc
tqTyaCkTpry/pxufL04g95bLvE4VDYY4m0sbqc5rJ46jKBjVNR8/GCVEKqDuT/+t
VmuPfRkW8QhZODKGazJ56w09B/ZT6yetA7i26KjkyjrC4KT8dfr3fI6QUMQMtMBg
W/lYvB1vLVpCWiCwYBl8ORvh8DtcAeQmLAJ9fbh/hWL0Xfly++MKPG/vXbqj2GpB
aYYPmdWzffT3bydYrVB3AnHrhlhvXqK6/s+wmcKYxfqLowL8DOIgZn8dsm9K/Umt
XVsW8do1LX4hLcN1JIlO3WbGHJmxIbl/Ya9YGF5Ct9Mt9v5C2OuY1CK7cHvClWlR
uk7PZ2uPxmtEKMZT+jGUvyX3SNiylQ1QJM3wJAx8NSI3KIb2CHSGzs/8+QFxzTvi
T5RCpA2tqYkcmVCTlArZRlO4sOUAgvvvzLu/PqPKG2mFAY2EW6AVODC0UV3I/lpu
rwWANpixhf7L/as5R63FbE0wPpnH0IUU8Z5LxKIlfwYjJBQUbsVDwQ9+XkL9l6GM
P4GER/9+aT70MUF4fPW/SPbpdy0i552RXLdHz7HL85FbeTat3An2nLOqlCaHGS3B
8+Ye+68XVQ2tIrnXZ50aij9CYe9axWpnGl7ACo8dHe172OP65XNTZ5wGQKkIU/CT
TYeComMMWBZs1TNvwpiFXZnQ+h2NHjcSqrPnhbiwLj1qTHEMi/tpMbUkd8n+SW2A
Nj4u6dB/lBacOuWWY6hNjvVml1qcXH50rM1vtVIYDGgcnuk7uqqoIewoOQxYc+y2
L1JIzqWkOwqo4DdiI8TcsdzWut/rYNFMe/ZzSMlg8fm1M3SE0iOeY7s9esu5DGN6
0ar1x0hjcuaPqliZ/VBBjk1QwPyYoeWw2u/FJZPMVSZCnnApmnxtLO4ubDgoHKDA
JWcNJQo0cNejULoJwbRQhaTuM10ZGLfqVGC0Y/ZGNd0b0RSo3ZUh/f/mw3zPqvse
yAOMZ2xEbiA+eTxN+DQ+qUyWJXO7tnTtmj6l1prXgWZz/j4y4Qlop4Zk1/vdLvwO
JD80+NOgr3uTErIGvdTe3BWvcrPQHzNU8r/tKVtvVCmzdmlrUMgdlVY2WGiIdB20
UpaBcVWgLHOT2r9n0zeHSZgKryaCUBcFTENdsqam1G2SYtKGCNbZVK9SUR7RNKvC
sLHLEAVjDUdGpj1u4/vumLZAATEXV45+C1dlPISBR8tlWdr5azkDlDdBOhnk+mEF
C048tqj+C5C/UDlH9UenTG25G/zGA/itQBy5An17RNE8hK3rCvjUfMAD22pM4JqG
tCwN+9vzFEJ4JFt7eI9AvAP6VH8Xw70c9Xa3yTc1jwnPp9MhCPi73ZjK35occUHP
O33qNOLx+ai93w2GVCZ6Kl3ffZlbTtIGPRyTjGo2wASWRmHNcrDheZXzlb3H6Qo2
gYlRpL6bh2WulxbHA01UcTm957sfiaHrM9aswDj9Yd3tr1K/aZpS/T3fwh5jNuD/
ypkSuq2wQvYzvx6WhaKkk6EljYJV9U4thoqLVGLmugItGmRO01Q0KQctuAf4fMNb
FHZ6NrQ/OoQFg8mDORVZSril19j7W/PnZKBnGixc0cwj15cULq5PFcErUW5rXw6A
jMAl/stBDKhW3K0qfDjsrDNZViReruYFvFpz08CUF9dOR33n5OSf4SBdLHJqqKsC
XA8G8JYwtVphP/K+1YOMRmAg+aZOmQRH2qrutXh2ZeqgNkwfI6J/qeB8D8quul9M
khj9qIWI9f3P88U4K9MAigRo56kFod34gN6en+TeKazCnEjqVMjZP2jzb3RHbrNs
t+24hXl4GIPlvczAkpxdof2Db4q0Gp4m6dp8iFxja80KFC7ZSZL5BwxoMlMA6JfN
oZNGFDlxeVY596r8g6oQQIDS2TZ/9OCDVVcBr0LM/dJFp8WheGU+uthvgswSJ3QT
TIhVeRs/VGhRaFP8Jz5zMR7/zMU7/tE97Kc/T/onfkRD99IbwZorQTKqaPDaCicn
Ymio9TzqR1qMFJA7Y1xyboj+ZwUgpNpVzfro4ZjCiVYaiXa9IfaU8MLrlwSYo/5a
Ig4iEF067pd7ONbW6aVgeeXol7PxcSAk0lAFEP1XHOFkHR/aH4eN4XCUeHfgP1Xq
NlgdEuUIA9HMYyCZ93saVPT99TsudJ+IOZ/QKdcZ0aZLw7gTBE4PBp2QHWvYIu39
88k8/5r0Q9mns3v05L3izXhj4aUtQWT7mL1DnTuXQYPqgVbWMQUI/YSmXPpCe5Dm
8vea9udpJca28YiMwDk1YC/goqvAW45Dz4a4Aq/5idPefpANK6AIARzm44ySOgBr
3FFQJ4KjJrD3c3BDrfdQp5OQ3AnejqBbpkm8b4+DneB8qo449U01EXcsKGNjKlQf
PpcblSk4p/aDMbiIeKz+xa3np60ZzZI6n5JDBfJYqs/+Sb7j/PDzRMn51Xom+60h
gMfYwsQYZLB4ty21GEV0DICpvTqqmRoWJ+C5pvacekifgC+oOK4hxDXkx768dLRt
KsD1aOTxCmj6630zeSfSwaqQcWKLAGL0+I7IZ9v46gSJYyR5MKXjmDASHzzCBxZh
waZzdaypMbm5j5ExDCTB4usMQ+odtpLQ36D9NXVrxIpobI4cwuG+1gGM9Izj96Eg
IB9GPe74HhKHaZa/4RKTFG5bc1jTKUDwNp+5hCzHsl9zbqUFrnf0+tIPeAP1iQ2x
voWAUA6YKSNpRo3qhmAiqJtzLlOxrNP3vIcKRv5VeJQVXAma61ZyqjxtPe9A5Ije
zDMCG5kMIM8QDhTk0lswq1uyhIHxav1ljAjOtVBpkkwfu31cqUI/G3U5Y3QVsX2x
sLUBJks0DLl5HYibs/Kgy/cH8z5Cknz/xSUVHtUyiWsIam8g1EvOQivUKHalsNp9
hbTr74gwSWlxxH2LmqJ7Oi4nYACsmxDY/7sdaqZjAB0XDzEwC7rUx8Vsw5zkcD1A
PDnNZznXNE2uQeK65zIgFR9ucnoCX1in2PV/W2WvRe8bTzUWeAqDid42T/bDGIsO
Qe9SZU0mHB/ABA/BjIS5dd5u+9RFqb1F2JjWAwlVvIwI0lz3TKxLq/8t8aEvilYr
oFRYFG8JNSSdKVcns6fVxywL7zyH5otRWA/+rF9eMGBtWqfOsTdX4iYG1p1++YwQ
Xv+Sz3ZXHz6lM8tW4OKHrb1MWbmxCbgsU61/m8Xmree5J8xsZbiKbSBA89MYlYZu
PSJJrxO5ydPld23QGNvLIZu3l41XXHZEjBHZW4SWK1MJGY6xJx077MeXO16Nz6tE
nFctcQ4PrOa9rfQlxewobRw/ExdqVTwHy0XBvHQbwbLhmOLQ1Qm0d1MAvaRTTiDG
0O8g2VhFGDjDehwIzk2YDa81C7NVSegKfqqPWnHjh7EmbwTrA/AEay5Vg7G82nIN
O9R3ymqadi0QNBN+2Nxkswlm2OUNwj0c3WU5xNRaVcRehS4fjozbARDFSCPe3ZFg
7O9TH1XucZF12NI9iQClr8Zc2F+S/nQxxqTnEfKWbfcZwODpMfX0L2DzMNiW9aBt
K/yJrn6O2JierDZ7uxiLMwgWuLvespkHI/D+lAAx4I5txGmMRn7/l4Ci0Ie54Pcc
9+XZFlo7Om82xvqmJe6LITvTTtMEdWE7qsZ69z/QY8KEdjP7NowY9dtlc/sFEUM9
VYcGdbhwYizrzRfOj6m/gQfK3HP8ao9ExkWXjRTlLSjPM1g4csGFJzV0ibhKDtfC
bDMa1gJOTqRx+6ZZT8P/OPjVhQF6rB27Z7jiR4QLPW1S1OEO4/X13iKE0LsOQzs0
OnTwDSinS+AW6fyFpAauJN1c9zs6OkOLvrABwVui9spXaVHhusbaF/vCwXODM1jq
IwLOeZIfX/r5DLFkb14K2zeJ4I14mRHAWS8lYR0l4tPS3QNMVeK4LvX2Igch5/0p
WejF5Gbe4f1yjKHXrhjAi9vitILgdA0+krv6GsyHEDioZGvpGeFs4aO2cZrE66i5
Q0V+mvqGNZ2jmjTj6nCBdETv8enoTbqv2vWWTVoWl3i3S3RA8crvaQNGXiq+XrSM
vPSBRLpWwHLjYirisizE06uA5cLNXCD2clnVB7Aty2GZYUOk7HIgeF42kRQIPUcT
u3A2EO6t/03fmcMyhYo6pNK0Wm0M6u/WoPpYGzDlZCK4XBGrndIktAf3r6p54LFE
mvUwvCQctyRZRMmmCcMI0bFKeG6C31JcfUpdxH5/xtEkqCVB3szIG1fAH2DwmrUU
ZAslL0yZ3qMdQLN39n/wJF5AvqpGjXNQ1P3JeIQq4oylfsXAkOJCr7Ik+DbxuL3F
HKooyDbdGve4ilpXDJ6TNvq+U/wFIUnbXUroaOHtn0hncEZosuqyivMfW1MT700T
wCzSCdznMr2fyGpcqDehAL8CMgRhLYpjLkVggcjMonlhqztj08JiebfbgONNYK6I
Cnlc1t4FdmBP2b8KR+/eiWiL8G8g7QkEhNIDrsEfSAWmpbJC2wkND1iqlB00ws/j
OAWisNEYJyKC67dLHgXTIECzBufDyitL051FwjBwtIDUs4kXIXPZs2M9W1CPkKuh
mlfX/ixtfM6Rt3LmjCwKGJhk4R3sS4FLQhDM41Z5jxa1w5g9Kti+0mn0+ESomPb9
iGYWvzw/EKae2iVe5qFbgb1tqO4RFX6EBfew+n2/JDal35ex9+1nD7GfSMsoO13c
Q7xK6WoH3BoN1OQXaDZ14atxIQQR5RrHMko/Y9ly0zQh2LxcMI1KHnOXpZh33e7x
3nR7c4qKzSqar5HC/r26PrBuurR1NVzqueMxHg04zuadDMiCaDDXU5SC+gnX04K/
7QLyY8xyzo5iXPALMbsViFUsRDcxdAZg9RyCbkrSnYaEwGHpvpYeBXCInq7PZF9f
cSmNLkzITBozz+SkIJURAQ+lGonS5YsL7JQkkjMs18Iw6/P6ZLoRC8qIWsQcyZAA
9FbEDmqgQAhj3fXHG1HQVHAeZpaEiN/OUrHqQpcbhw7/qr2qSKMEya3e3hzUVOvq
tLV7oVezrgScvU346tQeQxb1Mu0F8jQI6xzK58Sxs5o5j1HwAi9gob18i9ZpTyz8
vJrSAXdwsTgRui5cNO4d9pMcB/CExrmLGxjxazF1ClumreK6U9MQ4+FHGoPWMNvR
7srQDau2l64HGQFmnnB3fDr4GjW++iubuSOGFBimPa1a0cp01qWskaM6oTGP3WWQ
cqso3BTIIVdooxg7fUvR805mtJw6VJmebZ4zl0M0AJCq2r00u5fMryJRP+LrtHyp
e/YEyO6GXlb1OaL0JGIddZRY54UQi3F0jUWC/UG1ETE1l6EV0rAzKx94W98X+EgY
1q6IRPQjN7Sht8a3gksrzO6/3/2I4orolbSJPULMMG+j++dD13JGvafhCtZXSNVs
HC0NfAUNgft/dWEKdQv9vsC7j2HmOVFHbqCFnwNOC1JQLJl87gUF7m1AIlbvgY9P
ZJyCDuVhvLh/cfkSC37UnZ9figG9GdDGXHqu2VCcTpjmOP83iAWTzJli7TwlRRpZ
ISq+cXlBJeK4UaBgAzN8HpdTp6ntpAbR6d/46xsFjRngBHgA4BK8Om/lPv43sAbq
yNLVoC2A5lbge6WWqxjyzKnmFcuPc4In1BaHTPb6xaEcxgPCnHWBlffu1vqUg1aK
wJSZbiu3CYIWHN3SSs9nbzvfach56j4g8LFqueSEf1EDjyknHD+63JzZchd+qx/t
4YepNJKCoSMpiEh0DWRfXlsib7JdbmhfeWqcryizVa9hl0Oii88YGxwSK8+mvAji
Tl9uC3AD1Ty1iqF4sakKQbxFRpRcq+NTiEmvHUeGTcZCI6rQfQfQdJUTnXy26cyK
/GoBJapty0RFqP42835xyJf8xDYCCJMLtQJEItNaldztA8tSn1KmTV6WHW7iPNXQ
v3G274Bh2M1immwMXZPM4EWtZ4zr3lThGPnHU5UfK/Mik98FsZMAkKpADFEPnHeX
DrYcHdtd98RV5PR/BHVol7hp6rcxThZM+QQo7dIPc0Hn5lEj0uMDrxPA1DJIldcC
cZqtSbuLHPPItZ6agI49gD0IQGWMyHINZ2zzMokNCjv22hpUumYeDsHs+CVLM6yD
9iSqrkCul4GEeAFkcNZvMVT8NJJoY8/KOhy1ZtymmHGW1p+D2aqwlI6Z2dKCSW5n
DahtH5uFyGf25tewIF2JeZ++FnWIFwqvGrG+U3Pvl5w/NNX4k2YRPlPnF5jg56qs
Ez+7g/ORNcmQ2dxTZwzj1yQr66ASmp0f3IAyHBBCofiB7kXh18EwYo23RVqz/M7z
ZrNfsVwS2qjAiFkxblRRAq+e0is7ph/jpZFZKth/gMiqhNk+an55D2W12pOMWS5j
7cXC3NcA/WXUBMkunc0V7FyAElgynioBs+4Vw8K6RGo853kwlljQv0/DqecO+l0B
8HCl+kWWEq7LRop3tkuf5KUGavnUflXunyXH6DDhFMrj+eeRhhaP/wyIY6AN387U
+1kPqcK7jC2mZvUZPxBci+MBlHi24yO3tUGcwT6G3J4fIMNu4wGlBV/cnq7IhjjR
95DJ2WoHrBJ0uJrtecoZ/W2ETcBKQ8yt3ck1vyeYw6iSEusy8UMJB/PdH2046N5D
3H9/XogejUFcXI/o5Qn8XRLfdjUi+lE+15xh+SuuEg1bIGno4hY85ZnPRryJkG5e
010P0IDASB4NyzimwcrvKg9azwfOcumoPpggNio1PgR/i7/gSvvluh1b8ez02qi6
Wpu2FocrRVojzx21OPSil1p3tzwRpG1z67y29yslMrkj9pZazgFpfyJ7oqYHzKRe
G+GFM0Fm8YABsGp2Ze1JuCqtJEJoNrjPPiEJWYmzRUBFRQn52Fgw6QuGtXqg4dVI
IcErbIJSczk0EZcPxigeYdLxOKZz90UhJ721CNIYTI0VYvEdR0Pd26o/W7PvtDry
5aRhc4bmkfM2mzbuIGu3bCCwtAm0xp9QnTdIotFuYKv7QBFY30xpw3BhXS50JpYt
bF2/HE4oUIeBxBaJQvRvU//zOg1S7HxGg5RnT9OFY2Tq7JXoug76pZcx5505x6m2
XoJCzGOMWEZv4vCm0s8KmJs6gfH30j3vAxqMnehcyYmMP8Izo3vPYrM1PsmbskxI
ksMw/69FPgdZUo/BfMYfJcFzwyMbWwNG0TGBhC7LhEovaWHXSbeKWvWsRexuaNan
/AI06nzyq1TJLACKPZDvzOP7cqDSWZbp3Z4ziY6G/vIPLg29aDMCl8ww/qc7Fyxl
l9D9H0kvoeic1iy/ZMEv6qxErnBXQzWOipAmVivvn6TrqRiHhiBzqf9st5lVvdjE
5roaW3MctP7Blk55aj5ODbER3aEJFB1VGqa8CC7NcdPPQjyaXfXYqfwPjOrqbFb6
9dqMcvhnvlp/6dmjGe+zT20zm7C/GygMKOz+vu5ZfHzGiQI4Rkxd9qiVt55ytGEm
iEGoMeYpygSSrhvnwmHX+GZRVYjvBagvruep1dl4+emvuqmJwu3XeqeLkPB8J+W2
uh1cpIKtC+WPh/lWGFc/25/5UYos9aKcr6sLcPsgZC8tSMTJ95CpMck0wYzBQWA7
IOkCNOSKfH6JQwLktS2x7ORirNaxQJH6UeQQ1VqJbmuXM8GRFzeTgY7ZT/Ep7trw
MH8lBGpJc77ge9QfXOOqwFg3KDQNWXFYPzvQ27xDVv8dVCrsSzxEWQkWvdczFj0h
5uvREL6QozOpfmyd7zeu+v9b1HPv2URBRl3F4yy00yWXrDWfmKBB/mgRq5xsoz4E
OZdXHLNhfuP+zqgudAKs3+zIFa/Pw8xvM5TMMcXfIryaGcbXUcDB2PsXL0DYVB1y
gtKR2OY4pEZoCI3fS8tHi4XIUv18FypR0q9gJalt/uNryyX55ByOs3CvjP3Z5WmV
WKtEUuhsO64lgM+fyJpQaluRqTo6xvsT6O/K0uoXCgMUW4iwDRzM/zUoyNc2EMJR
Vsn3nUUPHlQxHgwRMEuiqDiUsOAaZHuV7mDz2cQBp3BmZQflbbuJmRUEysaAPz6/
8IIJO3MupmgbO7F3YCKPjNa1Pr21VWLSTHL30vL2tX4UuMuWuME315gU9tHrGxQX
lxpizDpVCRBAP6Ou8GNdBkoV12oOrKDofZ0uL8GEamafSBSNk3XoL7Pm6zt2/Ub4
Ml2vN3h38nGJQAiqeJHa6hH/NAVslH9+4Z6Ly9L/k1BOIClahKP2HvhQe/ob2+/l
c0DE0SeQqYpckX0pfDX/oyjk9z43s8KytsPOpgCTghK8yjwI1ejthm18a1ulIO1G
cgV4rN5uow9qQd81p7sh8wC5tCbrS4Llf4K9n/mmcK2l9t9ojK+mJB05+eeyEVzg
Q811Squ/vuBJiE4+vd7YTDdKErVIKZBAOAGz+1b9UH319l8rfZFiRmsXsxOa4QZJ
Dvv3HXdZCrZ+mDtJozyBdci4HLfRW7UyCpmt5hmhnmHvxS4oDrkjdMAlEK5A9GAm
nGSo3lWdmNlR9ae8udLhC9KX4s0iXoU+0C+f4eYIzjZgl9pPo/TrP1jKKYYXR/rQ
18hYhu0l6Q9TPym+AorBBwC6bOMYPXQkWa7MLeJdnupJwQH/5BlohNW3btOQa/bZ
CkKfhQSKR4fzRUg7v8RhuaeYy+h3oFxc5lVoT7MsXjm/nZ11Wx2AR5fan8WHKFGu
dDC1IjO6N8PPac7cs/JsErDYuLaanU+ctveySQk4rcs2qQBD15Yz/Bfgr+Yl62n/
SHwNivF1mk3PRx9Y/Hb32UDHXmIMiQvjrFA9WfxG10U55yKZjctEcMZps4KWdXTr
mC6NgGquk32+s4wMYSyeSbTzmVJjMqkMqwbtByoB0suC40PIAKeGrvLCv6TvoOkV
adzwOomHVMVkYFNmQ6Wh2YoiquWlU0DPzrR0sMxHdovVFhJ4WI+nrEpRgEzo5hNl
DhMNJxiUrcFSO4BmGcVu6s63r+OtgtPeR8vHADvNGskMjSnAbIICIZyyzvAjL8FH
xlmStA5FaWAjXb6aJ/TxC0C1Xgighk5TpIPQ7hgil4ABLqRVJNrGXb3hxfhGQLFm
bEvnI/YmfDYwsqLiwtFwTnT8EvC4gy897M4cYC48RAvVjX0fY/yHeteqQUqwWUUI
vP4EFqkR6fWSzgL6G0TE4aN0a3jGJzO/1dTk6FsQ4vLWAVhbkImrQfY+oskEgLlT
ERPYLmE+g+wqoe9Mbx+I3wDmef/GSmpu38i0RnasbwFf5pNIyDLVv/5fJeQCCqBZ
B0A7DP8WnQ+c9K1tMsJjvt0Jijs51Lu7N3zMdY1LODwq/CXRUHc/zYNTkYxexNyr
YBXj6otCmUGZ3TAgvAWIVtfneFxeO+/hQO0Ej0DckziK0pzVPQeSyqn2ZQrYqsi0
PlombPP3SFPXkjCKXMxX4I4zf+OWH/fRlheACEEeC3g3uvY0sNDTxEQnIgkgL194
km7dr30YDCQcqx0D4JeANum+Qrn7ipiTUZLspw67yn5MZ0AWE7IU2hmlcc/wJEoy
PUXf9/nK7xqsPUCbBeksslkMi/7syagNfPNdPODmw0Y7+Ds6Bbkpsdso6Rq3hzTj
5H3bFdNzswtW03wrzYa7wwfMzejyOXbTjpzxHAuNHdzsavmsM+dBhLZhMIFQ6kRS
eTwE8NzLH83fppxtnRFP36vrPleA57cayVJ0pX2q2ytYq5uXu/zlBbyU/Tnl9Txn
OqTEmmrklPffJn/ExhzI47XZDWkAQL/rv4SxLp7goIB4znbOsQO9Zg5gtFZ0nBDl
A4oxcNJ2gesBYHxIBCC82aNhkcKb89sp3wgezVv5tw+9XL25GubI6m0B+ItYTZBS
ppQLd9WGo1OaeSVBtLCgtqUlx0P7bYjcdie/xJsmuiWjlibP34qA4oXHkR9l6ENq
HbHGvMolsHd8kty6ogYxhWCnWPFVbNC09UZJ6gBk2cyrD9KsadH6ddJ9j6MRv4wi
PYcu38x5OVOcOuTCCSXQMZobhe9FdJWAPsSm+Y/mYMCIdb0W+d9yLvwHyvH5OECV
MoOu+fW9Hvv+VW/HxjXY2nIOAIQp12mGEbp3UZJyR3iFgKm9PLtZZD8SJzP8RApX
joqeKJPpJQkgm3BQ93/AVcMYvEKrkEGjkpmF0EljelvGGNrKii49GtSn19OwNhGH
QhpFeyeWUjOweQvFNvm5ojbwKVZMsLhiAgFrCGJXbx5xZQ8F63RPnYNv2pb4HeEM
6SN/MjNo5CbImgeuzcR7iWQdnQtYLBtqezsiZtuVsJrFXud5dBDIweo9IZ9sMqqh
wkGBJPexQWjP+m+uG1RSp0Gi2Q7x1mTrxK7n/I+Np1N8BIozwtSM/ZqBR5pOXqKk
vXo20yN7TK9xOiiyWwPJpVPoBBofkfgIgjdCt6bKASiP20WmkLSbwX5cxbf2O1oJ
MAuO7P0yJZui77bsJdY7Iid1ui2/bDTdclHShc/YQ1p44RkqNU+wUySb/29FH8en
DKvHas7sf07sIyuZpHiozb2xakaiIX/+Tb1Se8dDNYpVMRzdaj3zY+5FPHQQyvVE
lgylgMObHkJod9k2TrV+RgzXmIC400lf1Ji3CPOJQZaCbEba3LkWDXckcajHGPqv
9fKrPrWAs8GH1a1HJYDpmUjGAlBr0yPPlN480BJIIxuzmkFNylDTnJP915KydaNZ
LPf4/I+lA1Wv+Pe8tppDp57ob7Bk6u79/UjbmJQyC5wd6cT5FplwEjoEMNYiQpc9
KM4SgpZOPT2u6OK6azMYgxtx6mKTay4qN9h+c40T73CaCqDA65OJnY2jqWCmaG7l
yxYqDGtXBTR0rV5bX9RlTBbH+feuVAu3D9mYZxBdfN2cbA4tN5pXzqAERDG4vyp1
vcAcQ0Mqbkn62uWnSm8WiKPbw7PgJzDxGs9qL6EgydaYvzSrHNF+iYIRPhxeTYz0
Twnh9IA5HhYH88XRZoIr7iEi1LIS+PQDJobdJdhHI0+751dPPaske2Js0+w95wfJ
ywhVFz1mtJZqVWrWLOkBrzCP8P/ssIPmRaayiNIIFm1/Uetoofjc8w1AwMG6Qxg8
5AvHcnt1zDXbwMTSRhBolNDXhYPSvs0R3qyUeLxPIJchusgm17wOXDz7O3tZc4m6
le8Q4Aqt+VncHT8kw+4Vt6MySeibGwObR0hnN/68Kl3ojwiatl9g+o/ZuepU2GH1
Rzn62/uo2UWA26BPXESE7RAF5YpP8bjW5aKVo6oJfGH7AK0lSkklhjogTTmhwLmz
WqPK8CIZ6oADS/Z1U/bk/2sq+Ldjkgs9iOya8tLtNLCx+095+pxdN6GYCgOPddTD
1YGFYgNl5KBuRGmbRa24J7R9Hjxd2GXVV0qG4Z/AbZlYiHXMUhwp887TWm4F+/BA
ETpsfy/TpURKUEwcLJEwZpxn2f1w+nmRfPaLhJ1rWFG1w7nxj6d+wYL1ShwComTx
1Za+yxO+ZbAzRw7QcPqh2ytyArf71UIk6rAHoaVyIs0svTIxc/HCmhaZb8XWPNR9
2mQtYc+5JtmKbHRzuRsogwyb4P3j7OeRtNVGLkrbraEZfeVANqXOwS4oov/a0HyQ
0rt01wMpooOb9mjdqH5QsU2oPgH8158h6dnqGGob3eHVDrk0KyGHH8JCyr/50j7x
ug0HnugUssDKI8fFheY+772iWI0ZEzhT+HN+0eP9PC/e00V4r9RQNZZ1mCCqMEXX
/2n/4RkgQL340cSlfIpT/2ZwU4h8+TuB6QVr7PTXa54C5bMDfJHA6uE499Jho2AP
0kMVAUxttN9QtiZ3Yjkl6RDqgyA5oqnj7CoCL49jTvSXj5Z0/VNE3873JNkRY5uP
O1xwf7PiEZs22lTO7ciiTkwzu2FtzAUVnfrib1Y5A/LUPD5FTfQAlX8azoRUp0BZ
qA7MBgAFIVvnXCRarZxmvv/uyADdFKj6+5mwicow+YTmIXAJEecZ1wcOc92b4qMq
+qBXtLdZzS3gU6n2K5jbJCabWb+twY2MviluyDtqi8KMPQq72lgP/gaWmcErtph9
LyTjDHtb8drUQ7p9da5rEsPnL0Umfbg2cbDUNc3pR231WXAQSFq4nvtxt+qFjA02
bOPA/f4A8XobY+vHIlacR9zfdyVqn9UEsU82vLrnYX34A7llyceFXsizOPDNgjDK
MkTCal2biAzYlEBdOpCTZj5aYxTKpopVF5JxEYABUn4ZNYCPdpNThO1iDfk/fczS
BR1BE7mF4uKCnNCaPuQg226d/5/iy+JdBhErQ3fBthlEO5+0BBIWANKopaHOcwIi
hpNy1TWud3G0N18FBZlZa9YqOS/wkTDbZUp72nRs9QHT/4HF00QYhoq3F+VpE+wb
uTOpGi2xW13sGp3iGsw9CyehipNjrF5FeT9r3d7+y9S9AYhXln6SUsAw6UaGv9qa
+t5z7AMOlB+SzjdGSKvTsXbAApDgyW7xjHBbX0XyEJsli2+q9/IV4yTc7muAEjM2
Tc2JrZJBYXvHpg7Ls1DizHlXUl+TRg3v5NJQ+92aTpmxvVBbXpCVvliPF56iRPN5
+78SiQUwg51XPBQohOu9qjPj79818gne0ydiUPXc8R5wyRF9qB78axCGAmQc5bgd
jsxi+xdkG2Igl61yOxUqPItC3Tu1GY+JYNRdiZo3hANVBf/+d279No7HeMavt8De
2W3wsh3Bc1jwsvOznNOm/kujJePYdGQApKyPMmSFx6SJmO4DCMVC20PYtUEae/qW
ba/BMiUXMKGwdpZcwPsB/D22bAPPvZ2DTPdbewGmMrBoYmg9sOPW5U96TVaThGie
2uZMwUNM1aMNYuCDEMm6/LgkQuuddut1npYI7DDPiNyEjPrEL93k5pqff8Rp3omX
WBXD9T/VXF/PhjE2qDVCvqP1OQ4/aWhIqQMitEf3Dh9l2qH83+z7K4M3uFypmr5e
v7FmGmVG5gIDOGeNnIFpw+YmybO5XC8JO5XFl063AY4BWmRMFwDE46hVAKDiJXLi
UhEBIZiOA+kyytdT6BEP8w3+A0BDFIr+Ih1MgzLOo7L/PRBpqPs/B/i9VtomqT/f
sqcKr5iVZdQ4YiHEKGNCWMXkOD7DyR7dG/LDGGXceFsRTg9MZ7YB0TNV0qLH941d
6HDNU4s6GcTL5DgEFzx6g+RNKhWeE9xBzA+5717j+wAbOcVlQM76xSRKT8PnQwON
4pCbiCO9+UIuEuIM8zBcn7urY8gdqBZRmB8Lwe8U4EKwmhoIZ3LomYR2Pffbc/5P
cZiH14ckeShIYyLmVQLQHq3R7nl9e5dN/Se2/0rxUo1opbkEO7Y+LmSGVV2gDsB6
OJerfO0+oTlRBKfUSWPxrXE7nx+eBNuaxpqewjOqJ8NSxdBvv02nof/iCOTRBlUh
cWaEnW+3NQ+DgIYiEimw3A/2SiIob3j0D+uvlya+5pme83JdnGhsnoV8nMPezDAs
iLsk08c+GQQWwJfYTSN8fzJV01siNPhfsaU7JWF3WFg50nmkgvFqiGFlVmdgwunk
Hxyqaa2bFJuQ0Wa6DtzJQuww5hrn10BUlifOHHYxDviDwbdB7lhRPL9w1EnRmyez
+rEkZ0TAtfhxBexZqwrPrtMtg8ZaWBZT9cGCJSmdEadnyvsmo0j64Pq9xmG9CdPV
2taU0SC8sz3tra5ihIj+V6r3Yx0u34c6iaYIoOapm/hoNVDBwdkwTyZ+pg5ZIYvr
nbJyQ24kdU4Q5xHozLeJLsXaKsI3uzTo9LAN0g8zJsjvvuTVdJOnprhehehRUnmS
IzdLPri1gEZ5SDHB7ftSGIKN5ey5NGWLg9FGJNf5tY4jT/GUPUMXJijIzJwI7tCq
T5YDe2VSJvthss8NcUP/KlSaus5oySINoQrZ++wIYk9SeJnQ/PODkfBGX2vHdIef
WWwznprr7NEAuQRMVZKNSsgk1GR7hT5CH1bc1yYd8Qc92QpoOHDZx61HMHM8nUqG
GuzucjCyVi838yyuEp3bXxL1TVURU7RUVcNC+7auFfpc72Vn4HudIsbJ74j/SGTh
RyTg4U2unEciS5mG5ShTG2ydaRcJvTYsujyP+ktEi9aykeT9NsPOpdZvy6Uc0y3z
t8YNPv0cm08Z+ySTtsdwheKQepd98+keqodc082ybAWLtxSsgOnXzukmzIhnCVlm
bOso9voVebxFNPUPE6+RB9QrcEwD7KPI8U1WNJ4MtT/BixkmoA6B7/AIUmDyIHor
1W+2gD9ZxPtSIT4B1pdK86zU/N/bqVBElW7evKrt7bvIdzRdmJSHKTLTZZL2fLlU
K1CZXGD9xuycH0HAz8ncZWHGyrUVmnEjcQzNGhkiOA13qvAktyFQGybkLfFT8lQ1
bu/0Ko8P/uXBs36fZ26xdzqmuoNatFYvvfQmFW5uMPcFGwCyKQM8GmHHKfoyD3sS
KTIv2mrRnsjPXe8NxtUwFCkFabhddPqaVmrQxKW5l74/pyb0ewNb03NEQnDU3uCQ
PS/uisjlhZJLnAbbcaac3AKAjEcX9qxn++2LjrIKSckJU0Sv6RIoippQNuDlwUum
OUD3k2EbPS21/REto34ynEh1+k/g24/vg32EYKTMduzpoeX+WDgFuRExFhXNGLBu
rCZ4aA5FQUqqzaKYuH35S/YLQu6wjHF153coEDgNBJdvZnYGV2iElXFDbLQ0mXOS
4ebHtcRLOT/JI6sRN4/hDfH2OdZlTkKucw04v+hVomllN1a8MqijI7ly3vELOk3L
n8gdVsGjKs1HlwqS21/RcNZB+3UPwhNVZmIDO1BUPVuV5ZlfWMQW/GF+hDjPHUUY
g7FOtv5zl9R0VddYjfc3+qz1JCVtAKm+h+Psl56LvcdXCXGpsR+YHLt1QxAX6UCp
Ctu45CGZIv3ei657FUGXCifgpbYM229lVPDXIYT5KKrzb4kOi3RscYQLOf4G+gz8
W5kqvR49UdUQKFli8odYl+cr6H1u9kRKULeJR/3qUiaJivGxZysIWzfgekv7pdUY
dXbnnBQ/QCUJ9ng3PHNgkjAPwnUW/QlNqeqQD9sWsMxoxXg6J2jBau2RPXbHqYwT
5YIdYPYTfm0LbaPIAhXOHKimJkRuF/cbty0v7sgs0WN/B5AHWKbBnjefPyjHFdqw
S7lKQ1dqwU57R6mJccEqx3C5oMwei5G/ktAkQv9oP4z6sGl+eV2tuhgncNyl2/cN
wU9H9UsSQHY0e2BKXiXA7c+GbnsetUei3CSCDdc//StY80t7JUtB2+Bn4DZ2aOiR
biQSfc6BM3nq00cvcPKq4ESl13bn9BBhhzmZH2JbtyePqqgmX6ay95fGdqRg27yA
KuZ3oEg8LvrSW5xUxazajhiujSmKX83wgA+5IFEf6vCDHrFu2wbkBtX79tx/qOmg
SpIswnb1v6pecQidh2saJIiR94GvML3bQrLmsvuqPeo/NOvb/tSufI02new4tLsi
df3ciTAQDcQbvmYomFWadA/FKILpfQs1e2NxygIfmBKDVLQ148KvRiYpOZW8K/6O
j9ZbKmmFtTX2+Fez5tW1ftWeGZHKLXZbA4dlIVugous/6uGLBT4pWf+F9i58C5AJ
EAwPNULxZwc4uoTKPK5YrrHAzIdGmDylXz2CTLM8tcLCf1WDCZT+cRJEAr4C+xnX
aGEeO40PWo9E8hCCH3U40ud/iJVUbfqAhxo+jtSR4ga92YHRy3wVYehf+6kHK/rb
gAkefxmQnHsUrcdvyywn7aoKGQ3kT6yMKlOCb0bCkZa/GRS3LADDMloMPWM2o3nY
Iq1Njmlqpq8cProSR5eHNctMgPtJhPEN+DaXcPR2g3fW1W5T6NZGLyd1mlEMvn3n
DlxdGhxZolks9Uqj5ZfDd83pxaN6pFmJ6D5h0O8yJK/YMAQht5otMhPN4e33Z2pE
+kuqN73qiItyZeqMlT5ZN0Cuhkvlrb6joN/ZXxyS8l1WgqFx5rXYJMZHvLn5kH3k
OLI7u0EoRScE1UwIM8d0h6O9Ee2QMT1ogBmRs/CTCysw+oxIeCxiNUOybqQdwaFv
AG8FMjTQckQgOVkGF2CnioYEnFjC4QY1dbMnQqs67oAgGZyCBdbEHtaFFb/zEdqq
F67Oyo0FZz3SLckgvds9QivouKIAyBlzEhf5fg8ymw6J1hRTB3PxKrpRExCKamlh
7OlA3PbjEKv9W/T0eT60vV0L46WRJ9vr9UCp08rdxSiTX0X3ocypJAW5EJuTZ4+W
kSSL7QMjAQQ4UPoFkSxm4JugYv1ZybJ5vtcgrMOKoe//FDeo6tRHKAIICdn/XmqZ
ozFYaMR8/Zw0q2hngGVpN6kXObHkvmEQgS7K2bIrlFi5ussPUConEzLBRLxhELfd
X9v12kYcnrblnLz8DVp/c2tKMjHcrUqaBuAlgTdANxLTUf8IxpeeLu+UcMR8uBVU
3e2jzS+vT5rKERqkoZnAAFCK3pYyw3uARXWyKFty57JFijvwZqKKwP06NamGHcAU
b5axLbZ2C6NxP83BIUz4jZ8gD2/Nc2PK2702bwSrNEDnUBmar/jJPYxFY0O8zKCM
hCytHi9pDqDBUFsMWZ9jSXxgPWLtIGd95fSUQRubfhGuV16sJ5QEASNn7Z4ww2gN
A3WiMaarmgZu4ekt8zecq1lqalrm5qaO1A+7iEXaOsxzyHiP6sUy6gCnFTPK9Lxy
B6OK9kkZ7Lt9jO+/ybJaveqjgiTh34Hdp1Ce4Ys7KVuF8vXqB5eRNgqphtcGva5m
p2wVGksGZ/XSDPbVyKEZhv3BVmDBeJlCFiibD0RE3iwr1nDdaQgEz0xaYk7fu3ju
B2V8nO/0vZGz2eYETduPUcaWebTGP2BA1L7K5131H6CMpKKwFQeGN+WZ7LMzFyK2
kPrwkZ4XiR7v9MZnTOHjtqusjiOZMESYhKeRrzQcMVjrbxbZ+sF54X6jFc0dVtPM
tr5M6PTeqHVa8u/0LqHqgqPEgfT025U1bEgoozYswtvGnFnXMLLBQlzhj1bRCBtv
TeBqPxIEQZCmRCTXef+2EA/zCXjs7O0B3ytJyvNuaOjneKhCPhVd0w/bquSk4PSv
nr6tXDXwbcpI+8YM3YAtpNe2FyGVwKjUIkmmF5EvupOGn5dqmDhUiQaX5QuBWNxV
to0ijSxaZhDjrkP4UftrqIrwR2Q+PGHMDYy2k/AzlYwHbg+Y7DflaH66pfzKd/PN
ZH8hsA1K9+nnN1UzQyzbB/b4QrQnRrbohkXvDOXTQ4QZrUi7C6qbEzhaCftFuMF/
qxEuhnC+A3D7MwIUsKSCfKcrTjXo9wpDbCQdJvOYO/qZSpxNUK3Im3nPIQ9KiUQ+
oonGOTQ46BzEJA0oXh9+Vl7EuZ9ExnU0Ejjjo7OtIw5umMxt4YgcO/JSStbsH76z
2xBqU1ndNxT/OLx/YQqdF/MuCw549Sk/lyYrAw82ImoFZ8RwKUM6p1f/nBl7Kt5h
OlkFAJ/NHGmr+Am0OAsPo2Ta2+6o9cGmQ7b2xOKPb+Q4QL3txkLfyH1CwaPlgspd
cucgpn+rf7AqiRWLRPdIZXCo3PWWanSS3kuBLRoPDEAcnW0MbcsdIAu5/fP4ZXFB
q4vGd5vRmsJCmSzBlk0RGT/VljNkFssdREAOobwKomfrFRL4hakLSPaeytL23gF3
agfgRNpTkCDPmbflJuLY9Cm/G1PL+hBWNXLBCnTR2c2O3Aq0BDfWOzMx8ccHV92W
5W8C9aziBxTWcFMMMu+6Bz/j/zFpihHff+QYMryTwZaGZ/fnsAQ9eukjaDyZOM/y
npJKexJgjLKUsIfgrpkGg3tcL5OCBnzZQDcIDHGqyfZgARrzob9CSkHTV83La7ek
f4YUhSGhT+bifkthaxluLH1dXffW7RXLidkyq55PKD/AEkduRvk0zfEEKkbuDmTr
ktwkz0QhHYnyMnP5thaCSqOJ/gavMJSWaow39u5k9tH3AKnUjDYHPLF1wZfAUjP7
wVc+ZyA+r4h4GACfD7GgRabtNvZmu8Aa72M1rz8EKXekDT9lSQegmhkkSXkMFIq4
IITCM8jA+VnQvRM3vLAnjUcYWyZEGCmqr8B9XO1wYXvOu82RQAVrtMSCrIycBtUR
tInKXieP5ygQEnbIlK/Z/f3gr1RM939e4/XFY50uwti+U9B4ZueVbyXxdDGNcJRl
RjZ0lH5Vj2VHCcx5o6ksKQyz/XaIsZcl357jVNCkvQt9kEB3+WiSHDKWFNxKUQkQ
KUhk46P/jbit6qURsI+gtl7/CFTBQKyKtkURLZHe+zQPxj2VMMMCnDS/thAaeqO2
8s+W4Q2ygo0vQoRwd/TPPwMjp7FecwyU4atpamOcRp2fGKn6hNJPakGV+hlouitl
KSpMSDoDxr4HF17B/ZCiLhhvluLSRQEd6br24BdnVnvwv9zkppE73bHFFO5icwjw
zN7sqoaB6iLlrPZ+cag48RiV6AqIehEabDkq0bVxHUgj9W7douGfFSOy9N1Wqmxf
gPd13sHA0KtRt8RMmv+lrHu6TnxLjM8K64RlrwzuYeColVL/agn67oLZ0kDMaLNL
Q1TK2wfcYnrsUeomDlqivZGXn5uPkH1QQZdOljL1dIOxIzXem1FstgldWoQ5NF6T
UGrpGpe9DDtxBxkdfcNmjWzns9wImXFhiwMOlP9t3ZqWv11bzJiIoCDM/OUl5Ou1
NHXfTT9JiDPtmjfClmlM8Q20r+GIq4PnbBV88tOknPn+fiPM0Zbt0Lz7J3G393aE
K6/6jeqfhiA1Wk/gJoNWQ75DyldLxzpcujIJ/8/IMMQq9SrydvMMaAqYJeO4Wydt
vKEg084UBPjNL8pQlPbzN4F3w7CoL+2OLW1cbY0bE5uPxh0ZQJuLuRXTCQ5oMqq7
rBpqzAZ7hYniD4pFxsO+OiLJ3vC+4z82eTnbCUj1a5PZ/lB1odAIWvCRKRuDWNP1
/mKXrQKfvGAklSBEoihObKTZDGBtJgjLzy7OmPWWJ/M8lBJbYixNdhqXODuPmBzb
Ct8fWq83GMM6mJNgST8pxzNmBWBb6QscQcVjhtNAM8OFPjg/tB1q6iylkmptU+A9
Kf/DCjT6U5mlNwNJ0s+aE4AnIOfYvsVzwPCefEgmpf32PFxnzqyTQp0mkZVL7lT3
+dlvMffa7R5lEGIyhdbMoO3lRlAlNiPxicAa2xy1hCvmQuO/+l+oe0kPf3ItCah+
EIgHiCW0j0v5BUPI9GpDz+8kytjyFXaqpD3Wt7LKS3Pg0tZW6IvsX7l2JJVh2aiX
j7P0E9D+1z7vm7V7G8mmos9cF7aA8TFBsB+wLcdNUzAmmvSz1OoruzwvslkyuMWK
HGnpIwUS42CMJzsYMG5oCOlcEyeMV6a1L/X5XLdhcn8JoLnaeixqwCk5Z0pW8fsb
NEly6Ix0osRnaDf9bBWGGl2SJljE/BhwDbwxLK3Nhs8RwQ434zEIyMyiAdcayca8
OzJ7dnmsS3SQqwBToxW6aO4w9l7Zct8VaaFDyzfgU2552a2FCZAkzCVDoP5GimuU
VmbHJ3L7X1PxGrCqm7ztES6ImTik/y9isQN8QzbxGSf4QKFGoio++UG/36Sw4FKg
7PgfPbNpCf66aFATmU5jD32FiKGLnC6DRBolPlxnoxDbPOM+2XSluyuJZ/OWk9Ns
DsvRSrE6zrnplyyRU6EZyNmrDhgdZ+8s4zcQIry8ppkfo8bcUqV5uCyr3lW3Ajde
S2bD7d649OM46q34BMlNAGhcEreccLkbBrBUL8amdc9byJNuqZ/N9/HZo2LQwbWu
WiA17RtvMSnrbJCaq6aL2RZg03AM6IzDrBTled3B5V5CheE1Na/nYfTaGFD4HDuI
Pn3Fzaek4XpwU6y5iDZ1uJs1KKZgnXnBoAvWDl59sS+tadiaY4bTdbgeiNVCqbhS
oaFpzXRnYu/W7YsNkxe4cr16ApDZxHTR3knBPscSV6Ik5xrDCZRRg3QP3ojWp3eY
jDJHycbgB4FUCfPPwIDXgmXzspJnTFb90+3G60EHedD0lClQ6r55DHAZ3dCF2ScV
arKpMf6uRnlE4yCQrxxGfPFVoIAqgH6J7WgFhxAc1MeAd/1hkuyqbUs4/J5OiurX
s7BtgZi7zhn2FShOS5jffS+ramS1adbFI0aVKUJnVlq94Hkhf++MjcUyDzi3IVww
l8xhgZgwc8ZONvvT6PGNbbCAprkNfgyielJSmNF9+yB9k7ReuV5MPXaV39AMpOrH
+I8grUYIJ9a/Qf0FSnrLNYa7eI8B83DjsrgbWL/rxm64va9/dR++wenRzv5i+8WH
lw4AZSj3l/ZmQhDbII8e/2LgNy/qw0k8Z9PFswKaLiWc5laOJjwizZppB1t1N9No
LVoPEQKqV5ZYJl4HnAHqh/3GERn886Cf0pji2Q1eAuNFkBpwW/DRKTsZ+hUcS7iI
9jbr8R/DShlebLR4fuzJsrIS7mdRg0R7O3QMtIIu+kQ1nyvq8evhY5yr1Tj+kmEB
fxGcCvJNmvIsYIU2agx1AJBNwkZVJatthE6aKqTRetFo6w2YwO5LosOWVqoo/m/w
oJ+QdqkcPO8fNimegk1KTXGWAhVmS/tXSfItz0/qSymhq1NHMoHQ5K3H7K/ndqb8
oD7GBPmOTy5vaycEcyDZQb4Zve4qiBCSXtIqlqGPxY5TsM31E3dnoBJND4mGU05O
w/omuVMVgwovZE1DNOvJAikepcNWel3cECb0vKJ+U2dakeKxu5bkL+otMySE/0Gs
d+lQD4BrEC9av4A28D3H3jR+j8yZU1dauUBzjcmqsig2lZvjmJz5585fpqYr01rT
+T0v7GpoQL7KpKAmD0iuav/gM2quro2LEki9Z0tpqWfTODdqXNgDYo88nPKdkZuj
O0yziOOv5+quo2demf8H0XNJKs6GqZVs2Iga5C4tlGJNfnITVSqMPtgjHapzefQZ
MlkxbV0olSphifvB9HV9ZkGdKB+O+JT0rpe3e+UbTiePKBokx02qFgKbyjpHks8x
R+2Q7DdBeDHmVW1mao/IIeBt3WD6umO4g9xgnoX8o1IhXNqBqG45FN4HUIvIA3n4
NfGmjCkDq2p4utCaxaiiry9vhJWSBOZqGH7JSU7YKoAd7uYs3re0wu8Ld4ewOzO4
6DsqyWmLWnCR0UgfEY6yM44A13xp2HfvIAhHt7KlsVXILN2sF5ecxoN/J3vchgBi
/pJyG1AfbK9BpOW3IiGH4q3Owcz6oP0OcKj4ETAdkJWEBOsB91h8H9EfYV6hChOx
2HxNlCHOSA2gXuxLbch0W3imQ1xgEdDW79h3Ld43IyugJv0GZBWJu/Ab/c19i18S
dtY7OAcvS9ZX02oi9NvABMBBH8ON0ZqwbIbygb95zyG5rApBYbb6+0i9HzMG4yZi
pabAQ5qnJNrnNa4xeJ4DQw+W2ekca2WtPmhQCjtGPZ4GOnM3gvs4mKiBVynU41hB
Tsxmet61qR/caU0QmYDtz3GCyhDH9BQ6D9UjW73aVA92t6oXRAgNsL1gSipBmvjT
RRfU/qGWj6Ao6hLS4DdI0jeK9IiTinQ6esmssaJD60w1gh7rMe8kTRGfVmjDHVb5
vRPC7ZvrLmdkgQMSnMMjlfzkxsIYMmsFMDlxh4xRBiU=

`pragma protect end_protected
