// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
vBfKfNJwfM/D/VH4ZFRpW2J+11jj4gr+5roN17ZAySpSrfe3kN+enxV8XEyxiVKB
VBtafzbJ2zOGuI9hl0bUzaTrJe3K8vo3VxLh1hGRyzxlNN9pOo/Q0mkScEllZaDQ
yXBINgbF7/ORBrw24L3E3GFvzFqkCArlI32YAc1HjlQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2272 )
`pragma protect data_block
d7/nTl+wtvhTN65AYK877DaURWwhIJyUCQBNEWlVSdTHDzP/3bGuA9NsfypwokG3
DPaPjRU3eQVPLiH9b+aNE9qN2i1nB/zUjYy22aQO2bCwJkBeFHXq52DAeUBL12JY
O2XuRiSwoeWwRdZqZzLYSXjQPhrC9T4UIhXUCE/r3E18Q4UgqY13F3s8jglFVxQz
y5TRwiwm4Yw+QcaeV+EWFHT4EVL8bTp8tnKmHWe3yK144gn/GwEBawfS4xQlRyEF
2yv/8wXAKs89+Us629ybdr6094yNns4dKseDOg1iww38hPIbU1F59gCgMGUNbA6Q
7Sqmw5VE6L+2X957bONEnPuqlgznDTjd8pm7q/OKiDLtufPsXUXvdoAU0EySodGR
n374zwKETd5OVg3kksJJb2Wtfe2/YHdEdXqzMPkGQkvsV53rFNqT3nJpVQQL+ncg
HIVxoJ4wZGMsm9BBGAYZoj357aMhosNqFPw2vNSYgCcQCRAgIosGkbds3Q300kzx
1mdG4QPheOTn1BeAtUqn+TSA6hFf61F3A50qmcWNMTXMGhILQ9Sy4iBjVq/j9Fse
c0d4F9trzsQjlf2VzBdYtwzuTXYTgps9NFRePQIlj3ha87RN1+f+uqjOK78wmvEG
wGI8l4+5zRxoZGhoDWgXLFbjQxfhI5qMTRnl+/YDMYXJ35bIYQoWFYTx74a8RjBq
2Ies482FZrgu91vXPVOsSMzyP8jeN6BZ0DXo3R2Q6trF+TztjXt9vXmsMGnxPjnM
afIxmzcXx3uQu5BYGJRUbd1WneYCttmopFKm/9f37vUhvO2R3sWtVoLmODeW7DzU
1zxHhEvwe2hoKpdaaMTRF6R8F4ffdC79GBN2O8KjnozstBpIGwAPKCfs/nKOu07h
FqfwBwyW0MPEr4tGHdfUJAps42gm4Fsc/wr0DfxcOYe7YIIU/+lwpC9hps5hjPQs
m+2ohG0gBq+RJHriJJ5p+uUl/aWuiGedM+jm3T59yO/jd34JYVWtdwUULSlCqxYv
jJUsjyuuRUrUbN0tCgs87f3fI+gonODMQGPHmsHeNfmVQr6wp16x/8ceCQhXzpXl
TvY9Y3qFEz4SFOxJp6mVKNektjg1x8rIS4GlOYTKsL77lXwVLjabnL/AgzpWQKzn
iozIdLvu0UoDA5kkyQNo32duWagxWQXPafXKsQtwuhZLPQKdI5THa2GVjUH4EI8n
HGTQOCUeZCJIAUXp1Td7QyQk+eog85UfWX+m7sQQfF14I9FHia59oWentP99R4ba
Cs7rC2EZorq8Lth7pXEp47mKvBiS2G9OngeExyAh+Ubk6akRclqz4TX2pFOPlnVx
2CShAQhZF/+por7mK+1+QWuxaPZiE5OkYdt6reE0G3nvTQrU8NL+sQxbXGmobvbe
PpkUTvdrNa17BVYBZS6hwzOuQcR9ePXM9KKVVJV/JasqTHsh9WWQWiNScYlzhJzs
q1+gcMXuPjoxCkaEk5iOQvptWw9CyVD4l526BLrhs93XXzfwgxkWKJk0EeH7ZJiC
zu4H8wCaszNScya1Id7L/zeJmwOuXT/hFPXa5HaGgG+eh0qhjEPnmkVIEEBd0K4O
LAGBYvSstTRRsibAzfUbHTDiu5/xr7Fz72dUx8GpuBgpHrhjL7esNYo37FQAQAys
vt27RRIcHJbQCn53poZrPPs8I6yPMCRdZYVROyAdfI4kmjY+DtO9aZ8VKO9ThB/3
QoiBhrYdjAiJDXXpZj4ag0EwQ8UM9DNE5Y7ZTQ/pqaUEHzeiXln5UwgaKgJ+rdXe
gY1anhl0VeAMQF0we+drZeTkG0Z1MuL4PC1od3ZpKApLIGbmG+lAZHmITr55qjZu
suBxOq21UY/BWYdRou/xq3UG32ZX4qjyEAqREEVoWhftj7oei28TLj6fkAuwC/kq
ZysjhUB32/NjK5H0OBVbt4eemMaKfCp7zX6mdgEEDWjmqZ74JjUD9txPacITEmPx
RBe5AEpsgCruljYsMBj44ystacKCcUCOg+LtG0KYC3e+PMZ1ZL8qb4FYRaWkOOi6
t3LuSDsWLsG/8GmNuYHXKJQZeBhI1yKBzTpuPtQs0OYkVRPrMUDwFyC6YFWXEr/U
6quXGVfF1i2mROaqYBofytgcJCR0eEldDabAZDyOdcNd0p16fbeBg2guaHOZ/f/y
bEbFyVNIkKK271RgYDuFabJgxnac+X8TC8y+/EymuQPKmz36dfGnOYYt5GoocA+S
Ul9PXO/Va5tkwDPtg6qNFusaon3hOuxlJu8z+TIoNOId+k5O1agt5cseG7Q6TDEm
N9xUZVAeQXBnHDzj+G/b9djLCPe7TlNHnGLSXyBxUNDQ89OazRRGsDsoica7LwSV
Nr+/M7jeiOaL4MCNCmOmvqk2P+SBcfPn67RPD4GydGNXdXFuwLUDpanhL3gA5t8B
5bMf01rcUrtu4XRKDQwzhSGqyuyyrMS3nLLM446SmTwwbkB6fmHcE2/u24cKgdM4
PVoPqENbE33GaXZCGMSEJ06LhZ+u/yYfxDZdzLrvwt/qNCAJEttA86a0gOgoXaxB
azkT38A0O7//OzrQpo1Wiaxim8P8nHUFOPlpqx9FqXENDF88TFDuW7HdQqayWOhs
qPhGSGe3mtjQQmGr481NI/dHsz9b73ek5ItndzF2iGEnhsfByFDpLFNjvG+Rdwam
Z3iFjn9n+T+asBjK7pBxTPzb2RSDr5i/GfUWZUomyligJncomVZ7XfPRahTX7t7+
essPGcioaU/Gh8q2wpp4WrLEeP+xshPs/Rb6vhmLXy4lC0wC6vDtvH4vBRKy9XQj
dIfBg2kXQTWATM6e6hFLbjxrlg90UuuwLc5gWZjm9GKxvcGRoijs9qI1XWTiIoKt
OipT6pGlH1/h2OeS/AKNuaPU6jJOTZkDVcxL8zcLijS/aSN8t4vkphK0IdDYPXlZ
FZBu9FduodO1Gc8ROW4TKsLl8/bFmmMzZY+PIGY5OYz9y1yAkAMIWpIDIRRwi5pn
oVLmMcYla2prxga4pJAhug==

`pragma protect end_protected
