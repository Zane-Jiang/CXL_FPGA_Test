// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
s26QQkmExT3QQ7qVhjDy6T4YQcKaHMzIuepFjmHuOHgKWdr1Q8P7zWalZbIr
1f9n1Vx/FcGp9cx0YDsDTBqTUdJoe4bPICHi48q+FGMXNCXeDt1UtZ42J/3u
aH+ajaKpuHkEWvXxY+PPGNjLiovqxRvJnC5v528C5BRs1y/dkU/WQtn30FpG
6Ze9A6ks9QPbwYvh6dMZVsJ8o8yxBA08LKLwCi5IhXqstFrJdELMHAeM9gxB
kfrBsfyNgkDTyXRu/Ygph7OOsr1XTDICswdxLOqtgVC/IN78SGgsWMElAeNr
EhYY9VLevnnWGkFtqoLtyLoaQ3jPtim0aQXkDLAkzQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qZYn1nsFDLIK2acTB+21b17+/WILrFWFKfC2kAyFtZZwYAZVmbTNO8PMoGMG
qkst61syoYzgjokZ70os5hSFaz1owOFeWEgVnGHPieOdm3iuysIZPzZ5OwNb
OeW7DAI9pF1kSAZUa6yuc68rkrg04yJviJhUcwTZftH42UjU8pFQjlUI4oTx
IAmKliD3R+l2xSOtIQKkS/zUPVsxS5HKaWKCyROeFGBmB7c1SEjJ3Dk7Z61q
F+kQxIuDbK7QIWE+mHbn7RPXhECDog8ntoZzg1dx3XvDoGCzNpN8s8DuN+qb
xZOEtqVmboSV726MTa0ZeNaRX11qcQcBabbFeBAu9w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PUBW7zZgi2dBLtdBxmiyzsIEENNKnxI5CXp5Sbn1YY9620LLMG6n3AFCgwNT
EgXXYWZJY+UVm0rX8J4Qoupk+iis7jd/+OVs7S09fbEwcHO6yehBuW+yIL+w
5Xc4Xl8HhEDxHtxRlvWjpJfOcLR6M+c6Q8Vkmr23Y+nsCWi86BbiJEZciO2c
Sm6w3Fm4Id5Edjf1vNm7/IKA6nBeYRJ4gwU34hsY851jVHvOuCS8YygtoqWu
vIVN+TwCR2d/GCp694qZlEdkhsWPQbB3wBAA3PpZ8ECBoMHj2kXekJXAdAPd
PkMXSTK9zFQC8vWl5eppLUtEnqu1vYIkWMmHv3zEwg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eE3PaXqR0+a0i6LAYEI88wuZ0luN0eUi355CZQsiG5+uVwzNh7uIpUVzGYH3
Ax6jpja1fYk9rrrJS5va9jUsaUruXOHyfIPdHtrqehhc/CZgh2/0XCoBhHGv
Bb7cP2g9+e4ZhYU5TFn1ET+ZtQlyUVvKjUOVqSF+jpduaBgvUqA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HQb7UHuphdMG8P6qeRVE8CStG1D3PCO+SMhERhdsCeMme9+MbTtaiYVwYViq
NG5OVKHcRBFlx9kPLnkKgfJQCxqQypAz17A16pYKYpdut12o/nmtNzvNx85H
sOORV/yyuS5ANiJ/65aMypNha56CXbdymD8dQI9OFVhhbj5FkAzHEbH16TCi
PBjKv5TGQ8GHoBCKs4QT6XzGVlSsNw4GxH0yVmK+gHYHWmVKyE5UONWi74O2
dsxHwgzM2rB8VbwiL3zpKqCaW5A2lVsAkSiDELeSAoWCJU3pVNMbzazuhL/3
gfcDzieiaWzhMStt5VuUj53Wr2QhrbP+lYffToClGpof0atj2Cac3hWKQhYJ
8kLpaGJYSJLxJDhCztgOnlGCEolcgH5Jt8cehsTdlbTBYpoheKVYa6et2ZbP
DZzhgDYRVqG/aNrEEqJ/wL/yvwwiH662CpXYjY1Jl3i3X9VSiW9f9nDf11jZ
J+GzcYCd2n/Y6O/WI+jwsK1EDIs+ifEG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CwHFXMKTeQ+qgHMTviGAux2YhG25nLfCYQGgNgqY1ZSj/MbT5HFyUMZTDIFs
H3RAXoJyxu38+VpnkrvCTokmpMn9kg/SZ2yYC5vfPzN+ulyzfPvkFvNH981e
HLAGXAbpCTZ6W1AMzN33eZw6c7Q5Rw86EaCKBMS5eeRUeffUP44=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BuG65+WxFlv9kPSLypoORDgP4JWlZmPCSLQKGhBLIQTNWBaXH+Zvma/Odqu+
VkHlq9sejd38CuCISuRk9epFhOWskfnOYRixW3yWNx/0wfp6sePrZTOPRymt
OBwKOPk0oNPcDbBQeYZwpKez1MlxM4Ms5enh8Pc/I+j2Ngjq89c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
BcT/99/sfYKf0pmH7oJnfRlGbtQ2sFtrZC18PrJJbn0AmDNjjUsdEWA90ZIU
NGN+ioNoN5yLJIifcBhP3yFf1jl+4du3J83vkD2XzbdVFvmQL6fgvmzzDT2W
v0/tAxIK2pylpMq4nPOABEmnxddqXwQMYc/3EuiukTulvvfQatbm7ZVdor9E
otk8L9EMu8/6wO7yuLM5UVvtDDqNyW4WrtRVYwQ0Fqg0lUJzUia+GvcBhJQi
I7oBwTJMNAGuhPIwrZcPFERHOCwZOWsbcnRmzt9evxe1mSO5nCZY/2TD7UO3
wpileVgARRiOF1pDcVjYmxW9dPYBqJdI9dpGev0esoqjNGPqopVQ4/ox4aIo
Yj5KDoNfrSqUZfRDT8dNPSJEVI0HFW65OlTvR1k6cZYsuK0dx4q3h5//OXkD
2MoLxIEQBqnklyZtgExi+qDkgpIHOMb6rpJoo8KB3K9LTKs+cI9i12sx9JfG
mPWuqldoX+dQ/T7dzvMTcr1tzqJQDETNC7H1nW1Vi5SfLrQ1MtaSEhkNIwSL
iqdlM6k3lWHn/ecTyfvltRNN1V1pkmJ6q8GGLW/llYkTo3i+ui65CKMJMmkP
QVm/Xck1iVCXwKY9KGLHSGtHfMbboM2IO3ucyv/y53bFuSm/Aitg7UyvhjTZ
BP9Jjk4N6vSw1pU2j4HRj8joA1A5NYIAdauzNaBT/DeW5n2pEf+IYRoAEG/u
pY9u5zihgEnWiFAmJwjfVwqByByN+kV0FQT1q8/6Ci00m29rFm1YVtMPOs+d
6z3gLvBmmpNH8T7itzpK9NLRALHSUvNLanELePWyjr0kymor+b/qHswYCWcj
Q3AqXlJh9Lj70F/SWU3j8nvezqxALKJYq94fHtn/0YEp51lgU4Og0it5kDLI
qqXGKApyJNPyNqVicOZ2J26SVa0Q/ajlCw4gPQJ5iNToOfpvYcScf4Xl1BAM
DSR5Dep8Ynt2W5bcNhWc2rMlCqZIRVb/DiWudtvaI4c4+NHd48R61I/pCSS2
H8zGATxkHfNlsU9mYMyKsGDbBdFbntKrVxqOLv/DV6ROryE3qNbbbxmwX7Zo
+TWiR+QL1Fe0HYrUHYkzEz1sj9MsEKv8hWEiPKXnoAV2yfN8E/1SZvrBWqSb
rueex//Sl+IlXx+l8tt4k4wuVhIMsaIRB/JROV4lVd+VR/N1PBoyLH42LcKf
nZBIZcR2Tq8QxkRxfh9lEyP68cZObnd0Jh0SYegA8b5MiEkI3XfLB/Iuxk6q
NPo+PvxPoAByNBkaaOmp+1CYLiQJfpDBAbI/9Fr2qAtbL5mKVkBCPgt4iedt
/sA+ykooE4nesn6Ovo/4Ji4iQ0zh1LlUbG/OIlaWikXGMhAd7cT2KU0aBPnJ
NTKXBEEhqD0LAChxhdnChINocCoi2uuZlB4q7llW2foF6qpcnu8szH8of/AW
qw4zXsh4vMX43REMGqCDmnY9Zs7cgpoEgZd6GC+R1pN7kaL1Q8pfhPA4izPJ
pjtmVet7YLIKEIWQammb5W4T3kccKgtik72VygTpthEBHTqLSlb+FhczFNHT
SXVbNmw7KGGOSjRE7mpcHk5d59/Y0oIyil/hQXTdZPHIzQ9Y9tmtookoTAWT
F967ci28SCTNzezhThiiRBfcCi1nSobpUR/9DE+lbApPcwL0UDGEEolDqhly
NtQEFQeKVoRQLvaYEPOOL3tsPNs+fjj9eVeII7B1u7LsiHpoEKiDFA+AKGOM
rPn5oOq8hA==

`pragma protect end_protected
