// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eZ0z12686mfdMl4OTTQrYGFdJ6BbpeNjK0b4v7aBBdIiLGn5bAwO9i5udD8t
PBWt+4eMlmtrsSpK2MYapGRlTGw0C5/iKxX7sSSQ+MMGNBQualrGHVHEVzyZ
/GoIOQXfHcVIdL9yGwE6nuMPS/fxwTw0Bg5toYmcajn9stqRw0guiz1zBKYG
S9JB2FZRBaV+OJyscH3dSH9IdVfPNXOY0FbG3c5d32KRZysccUszIMi7Tqnb
rXUNwmPL9FdL2f6CNbfV61T3ZvgT4m+SdAFctw03JQDz6TlIAtpFzSvuUHlr
tGVFE7qqMQIAk9WMBWPKWMnHTjhuM/KFRZmquC56bw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WMdMLZeX0BWAKXdHz5L6uGlsjFCxPOxvHCCgQ/kNWjPH3PLRid882pl9/fD5
qAdFUSfhVrvj1tgFPzstZHCgZ14ZVHUooyXjLDXGAJE2d7r6AvtHwjztYdte
MovjnV6ScvyovwsPLYIYOX9SDty85XAxMyMLzNjBYfSG8bZ7jzJJbVIhz0Jc
ag6LKpILvR/VJE5LYRVmE4MrATe03uWH7lv4fW6qarBPCZpcq8Cwv19YBZBz
6pxdJLLREK+thKVvkgvjzF/uOOoXXpQPs07ZwLNEnnyIwjlm7xR2mJoqci1s
UYAHnPR05JBe8qC13uM30epCDixUR5dyUcKITI57kg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kE+dZ12rs32wM2Yq327hBOXWqc0lpV7+R33lrEvV3tnfRwHW8N9tHn/YAiS+
Zejp2NwzFO6A6+BeecrozfzwUHw1Vl1DW07duZAo6sMr1rMlDLuuJaVL3QMh
EswUa1wzCYzczfFJizitWR1OLKyEs2k9bjR7Halp3k94OZF1r81pTIfbzFOd
v6H/AOBVCiqKKDtFBz4L++XKKQngNWmp0ZmMwQI3XMpRt8cvNlFojT6f2nwe
Da5JteAWpS1HXCL7e3mV3cdjS0AmbgIY1jesewQsZXKZO3WtqKNiYsFDJXzA
dg16IddnBi9bVxJM45ucHXy8MBSyzlRW0RsPeDrEiw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FwfLAYbP7kuGpHb1I7ECN50V3t0yXuzWuloD25VwRj6dz+Nnhc9L23Jv0Pzz
5AYGPVXHxfipoycWl7ypZoFgH/qpWv4YZP5LsSaz7D5W0BhDnTM6mGmS1J+v
UBkYIFPBi9SPRWMQHmAzLG7jFylVwQ8iuEOYio19d8Peq96GCpY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SC4pWXBajb/avjYVZT0z7QewAlwLOoP9pnQAuJExfCt4KxRs7BsiGj9PLsKk
ZYVYwQOvAw94zztuHdRwoqEtMgLxWoIpLOCNjRZCm6JUgU/lE6xlafqbOj+i
54wLOP3Uscq0SrpY9Ecagh8rVizpUKC6hurvxYmzy9vq9bxQdgtEaTgs/dqU
hQc7IXTJ2itKPemIbOfynK3YdZ29OwOwc1FVG/bRtUBoEKMf+jM6mHPOeXp3
AFfPmMhXaIWJXMgpAqTOMNC/MorC6qvy9B6vSNG0Q3mI6eC2Gs8V3XQHujlg
B6zpCvCWamgMR3pPmwLnDhGb5N/18PLkxiGs45pO1sXI/brgAOlNWh2tskOW
9rLcsqtJAkgFddKebwDuMp6u927vCs0TH6W1ZSYJxUrN/xOcH94vml6Y7gEG
TGk8t4m+x2tMfYqk06OKU3GCx8u9HNAjFwCyGFgqgYSqFY01SYgU/+4DUw6c
oAyK1eoVw5PWVmHhkMZ/0RqiNCUvxs3w


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pLmQbZ8bjmsrWVn3OaTK6oRDNOWqRUvkT1Ozg7/JWFel2WYna/c8WwMCwyZA
G1sv6prsfj0jzTuVs0eCnHnrsXu7WNTtK9Eop5MIvBYoEetEWE3+eEJoFTPd
mOOKT/RdiJlGt1fN8gRp2WPcw+Z4ICuHG+aoW4J9fumJl/Arld0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uSaGvgdiPGXInHjo90T+bpM8pFlSdjUR1hn1HUiBt2xxaYVpaFm47E/pUqV3
WnQb/nNtkXZWWZoALNGk0Ld+vhnxu5kCo8w3s8DKnoLO1iF75J1ft2FOzBrs
mmrlL+SLuqGNoUS3ovEVKKa8GUQeTDJNHQ9C1tbqVCjgOADiiHM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 133136)
`pragma protect data_block
kmR7lTa48xs4Ss0NM3gz7g05N4vNhG46w+KxkefmCyVfof/oVZFHZbE/ZkgV
BcOxTJJIu8Chq0BLcj8f2Xwg2giRY6Ua6PJv/d+J8gSTqxODtCD7OroVhqA8
zLvVUz29/t/ti83k6Q5NKBAh37F4Ews/9fqZye8ZUKEJejNWaoLcGCx95p4E
or7PP8/yrxQYeaEp1S2MMr+0fQM0YV3WaczL2KsNVuqV54nFSAiV96dBioI6
mkuZMo5PwNXt+dCxKv2bdmWTzIUahBanX1nj37HknWkYpw9/Wt54y62kufvx
RqGpnJcFAVOsAIAJ7Lf/K+XQVrwxwbNKU1sPAqauukQyBQ6lIwoZVzuqzk9D
pvpse3n2PlK1YIJ1ULS9S3alXArIc4y/LDzQHW407sSm5fK+ZKoM3lY63CjG
LkLRzvcnHaCSXCWUpT18L7H6PmEWfLjSVSe+3RbeQY538OvJOpgpmFQ8Wfr3
4ZC8dbvJ3DyrVt8Xhw7VZnf1q8LI+kp229Pk+bMCPbVDU1Xo11z+fyaR+ahd
vs6A6tWQxUNr+JdljYdueBTSwtb4nW/Q0u0hMKG/IRZpvbdPjtHiqAvqNqqk
K9XNrqO0tAR4T6snM9HWlYA65abx+6hiiQ7fJrrHqvgyvEOJ2esIBtP3/I4C
kdBOYYLK63vuCcLwcvvKGleKGpBD9j5F/vFy7DZEESbqdjaiPS7rL7qWipyP
i2zq4smBeRdAR7S97Vy6JtiVFhBpcyt9Et0H7TC7tBDNNVfbVa8QqyjJvB1z
BgRqS8ODMY0v/tNWQH0wEWxdqOMdTql463zjWMu76jRvLIbs7wLLg+75NfgX
WDfiwWBQyH1wvIIe0RZ/2d/z/+zlOg5aPSrL5uG2P6tF8fEGWx47dR9SCdEJ
jjhaBnaS0igCaCO3yuNGxf2x6yV9ZPyS64QxMi1q+fe29UfBz55GotjIaMm2
nAmNjmuvjQyFDYhSOrVs1I1cVL+dzFjLuODWK/U4NShElvcmKoew2GB8rjN0
IIEAM1A/X/4Pf3pgJSll4KVK+x9Hr6P2ELJAwnNQhqi2/boFvrlcvw3Sslf1
lUJ8tNIuLvAkuV/+Yy5/ZLAGbdI+at/ItQSl7ZNmqRm5UhUplMvtscyc9CPD
hEbBdDdBnp1gVP/vOkY9b8vOL2R0X8XhytBlRJkngbDVPe2bINZSKtuHAVA6
S7eXwuFl0dzK8HpJiTqoQiGW0LRVuEaIZUR5lNkkRdhy/41fHROdA3INYbnp
IaduR31XW6kobQctF5f/uG1k9LJI5SansQ8P+KReP8Rg7/iYXuPfkU/DQaJx
rFfJodmjeMCqFliRPkhc/bVXpzCqurXvqznLfvmbLQ9tFu/dkQ3xu2TSRh2b
WcFVyLguYsvEziB2x9vB/NNqQnoGZQoQrCIbgzK+jvaOK6A4xc4h1om3Husa
yR63CPRJtNEQnamrS0afXz8xfKGRKuq4DIx86PrWQyrDDsGvNs4/u8grK/Cv
L/SSIvmTbJh/PB8CDBhYTU6vD4JLT+Lf1DiZhZcWZXqLv+HPGkM1Am6UiH+a
YUGSwDPpduERRWck2XS38iYjNjILaLQ+lgUBQFV7h8qO0C183Tt3e0avmG/i
zvDiWhPi+F2UW4Lyak+u+y8wrrKoEfpv1I517ZdBAnvwYFwJyDrAVIJUhKK4
3fzqSYaFgDYI0Kx0B7cHo/3aGuzVL0NZlNVu7cXb0OQS69u3mO3C1HDRpr9k
FtNS0UYUi8/bqTX3lV+J42c66Qpt79DDf28iD+lqSTeIk36k0wZhbd76Htt7
o3HeS3/wbZYfSdBNsaEnbdZKhRlyt6rqObg67qI0oPW3UUYmXz9mhqMe1RjA
MU//pnwQttiAu3b9sqPnooPAqrSe7sen7pAoHlhKUDsza6MTJ+uKYcxLnBf9
geHWHN8G518zd3zAeijQg56WvagOORID6yTi1OTLwoRWxhrJ3wDUYJgdXXur
Qs9AbUH2fjiB/Jw37Msl05UVxOJcdHYrwgGuYm1anTq/T2gsAQocsi92oiCh
Nd5dfK9QF+v+p5llLBYW65CqzVleb8bdXJXqzcEhOqaLctLJ1k0W1+GeKQ30
u9HUus1xxbozkO/E9leN5tH6RZnD9Biax5+vLdzhwJWTWiXaVJa9kKsdaFPx
LnLbhe4EXoEpV84UVSBWFQdgDjP1pGGsAGg5MNcTWX+Y6KxKJ02VGkxwiAzF
dSidvpcucEmDZeFP0tza1YlX/HDADgiBwtsoSqjLXNrubVfQxCj/jrcwMpBt
53gThsJVMTzKmWlrAFdQ3ALlUq5zTjw4qs1lLr15qqkacxv1N7oBj6H6RGE8
cw6OW3NmgE17BbTpc0TqjZXZvhfyEbTmkhOj875/a2J3MzuI8nZsEHtye91t
DCe5wOD/e9f6yJxfXTQ/ilxAwg2n/sYIBk+Ltj5Ylmf0ofZcsvn47NsWFuJb
erTevWrRuGy8O7X0u7EI4k2nNaJ643hTnvCWjr6lXh/q17z/xO35h1q8QP5x
ZDYtGc7JVGaAdZ5mNC/DWGi39iFEDMmgHbxlWFIRXPb45wYQE0JTUZbIidvO
GUn8DdPrbry6urf/YRbxpbfHexutgLZ8J1vhox3i2Bbvy7EhUdTXBn7JztcQ
i5ALtSyLb1R4ICFcBHVxAwH7QjDaZTJFala6HTTJbk4p6OMnDlfRDQsL2tm1
DuHwjjdmJKGKO2Vj1YQp0/Vxle81S5yb+XoTulZEqg2w2rxzxyl+fudPw1Jc
UFv2UnB2dCTHBxPjF1GQLUXfUGdJZInAOY1DHDb87zcYHh0IYNqc5c0XOPeV
j6eXIiovrTmANfzZbPIpE4MkYrcIuAYDGIqmppOg/gqSZzgKwGwriJujTjXy
g1z5fqsq5VHogtZxvYniHhvQfrtStplYRcg9+pdKjOYYsQLfYfQMoEnV+cOp
bkJRMiwpIwa2Z3MD6IoVSuAeRFca/wqbGSNYr4rde1qOgbn73eZEDZw0ntAY
5FmZ0FV/dzMu4Lp0CKCJevh/EDwebKM5tPNovAxGRvy1JFEX2QngwaxCLvEW
sy9alRsd1j//RIQitIzAC26SWi/oCkGaj0APM25cp1uW2WnsSkusWztOV0zk
eGRhtZbqisBzbx2exQ/s0jXOX5i+xKZBHD6UHasr/qjapBg9MKzPGnPPXdkP
ShtxvW2gHDAP8n7EyUUBv2xx53Hxuni++MBs29WifUnL4TPdFLUT1iJ6qjFB
JdAr6eu+Tcf/O3ND2RaDKhCdOl4yb6ZEKcnAHnceaiz5/ib+fUGjP5Jl371Z
dI2i9CQ1IFnnQO5fKgm9fo9lbzzRX6rC8F4UPkAGWciO9Y4Ote9+COMcJHfz
qx4voucBTIXC0R5tHwyHbzlF0AmKBUDG5o4aSxvHj94v/Tov8JtNtezRAIhd
rvHDdYDjrG0KxaEO2W1q4RKvAkD+xBXN1Sgy1zlnngcy7vE0i8GfU8Ki1ccd
cf23DUJ4BuaSkBQAKP/oFOn6oJkAeQpealZwhNh4Snq0YE1ordl0fNg+uVbK
ts86wdb96GzskQwsY14SfK/tOX4o43VSI4d2aSKDkQWKT+uviFGNJDwyZafL
QDN0xStOISVti95Ft+oqSXKnmt7rZmxqAwxtRwZIlpJM4dwua7SCUvCA1Iww
zHL3D4ir8NNzNldef9kCzExV5SFLXxR5XRn0F9T5M6LR6yo+Le2NlPhCdIvj
fkfdub5l3d/R9UiorCYx5mQZIfwNeJ39+ccUbpQTVrtp6Lk1RGb9/bEB9iYm
800LitmFSneunuQKv6aFkktDFFdK5+2VFRGK4Y1Z/2azd2G0vxxbgmFkHJAY
zSoiMDVmANU+E2a2CSRG0CPIKLiO54ZunnII478ONfcfXGAl8GXKwVZSxyUq
EfgGVpwEzFEUvaGD5L43xVVrF+Qi8jOiv4/wP4FnA0QAcZCmPC+ELNTtvNzz
iSv/P8I+FfyGpNuvMpZfs/DPZgGVkyZRIqKQ8R/jStPDO6ncdlh/grtxwwFj
6S8C8nZuc1PBtcPX+FlEHxJ0cKe2F8Io823tDeD13J87eELuY1dfaB8euzbC
qQThbxcYpc6btGs81ETD01UsXmFMcXv+hvUYKOruDprNE2HiWCM3zYpAmiLD
W3z2KltzWqtBIEIO+AbgKzIeijr3l85e1IW2kqBfc7HGm9Eui5KpdZzGNyBO
AHMcMA7KSakW0jn1nudo/2+e/gKdCrHb8kGsrO2aSV/oaAprLWDkVZHE9rHo
9wib2elDgys/t9u483BNs8Ay1wq8YIC/VTlRN9fz0l3xDBI4PVYRitLM/q5S
+c7v9pTCuCFD2/P6/5O3Srrx1pgSlYgOHkezCaRgeerh7wxv89pazWkskyNw
dmj39cqQE0QwHINOpx25IKPv4Vsq2bDMH2TW+GpYfUvT6lhbzYUXSU/JUw/u
65UATfAmguWBCiKOpYaXX2YTbx7DBoXvIVSjweVmozDSec03wvOwRBhyeU7Z
zdNrjoOrqK472q+xPnzg+rNO9eSL+PSFKRbWg0BgFZ782lWzsVYAm6zPI4DA
YzUG0h5PFA+6iUlvUh+JCf6NCFmcZe1+Vr4BorX8usQolGVP+3unWWFEgfcN
Z5YVdcpT0RA+1DNlVWuPb52XFgmYWieYdI+0zbKVei97/zxbI9TxgJ9UIjq0
vIJFjGv6zFRRZ26B6HXljfM1ryI1wNXr+khFMZSUA9PvLMuBCMWR+Vl/gcsq
FNfV5XZJ2MCmsLtPI3QniEGw7f9jWpRONSzz9deQg6RY09JVoJMeelkOKFJH
F4tHQuq8vbF+OWBhDr/uTh8RfaU8aa8HzhBaNGWRJfaXow0swnG7dXo19yT4
52VFCq5GsRqAbTPZOcSnamCBmA9AjC+ylvXqeKQerto6yKeTIzRL6uthq3nC
tAA3RFX60g0/BIZ9X1Ee1PhYJc1/V3aYosU7zQTJJ27+ntM90tRSuLf6+LlT
SufZ9HvdSoHFzqkVGbBZruMLIpGHVpfbK19v+Vrg4FeNhX4OQdPnqpdjehaA
j3FtFbgdd9Cq7PeJTqutC4k1dvH8NKPi5XyPgfVTcW6oLIfYP14IcPzckusn
xRuu3+HzGEB07K40aVPrDzPR1zf7pR9OQZpnQislw7L4KDaDjN69pgbldsnK
ewrxdvFHPUn4obFOpiA2EC7FfO/eMe5hND4lwMkH/evIRPIxduGsa+wVUnSv
R4Zu9ds16xLx/5maSOCzmVrhjLdLdeUFr+FhIfFWQiETynMULXWymcpJH7wG
gx68yJDfTWsfrawvT2xPkTYajRJko0aqNxqieCp3QFj9nNvX74IA1F7UG2bV
Kc9MPG/shsWEiH/RQil+k46htpYeUq9SiYBh3JNzeMIlgz08/pSnWmo5hWZg
WUaczt6EYIsp2EIjSgfGv3sb3BP1qItiJIej7pH1vUI6Knm5hOUu0uz2Anbm
3tjP3k3IacvNzvtMcOHeQjcUttQD+K2tubmmzzCghlu3ECEk0TBWG4BxnwuQ
M4Grjkt0CRAgYboBlGCfqnPft3CUzG1fPig1cP5cSDYzz4xXQ/MUcom0Plh6
yGmNE0sMtVzYjtSYpEjIK4Qsph0EV50a1sUoP9UKFrd9N+maO6yeKH6+j7Ft
/LQHKZFi3V+dQEL9wpgSG6thcEvDTwF5OgUwgMvhhBBtUkhmGufsw7gbbr6S
czCdaVm/PAnA+kzuJ+ZvHPZFIQIIFh4BmzgbZv3AhzgpJqKRARlETb3CA4dx
l9z4TKiTP76d37djnVjlFqR+My9yKQpBbvrj000VHkDYioCBZGVfkGjtkwRy
cTBfHnx63ZjFepZy8JNUuSNVbfX0ipMNOSKt60NhbkGoZbu32nanxqWaHsjU
2tDbngZbYIcNjQSGV1xaP6YDlNTB6K3LKUWbCLkrKWQa04RK6sgZOamEJ0rD
LBj9koyYtIUguPEpA2iePblTenndDdzPG4/0baScWWDkQoxbDeR7NoczOpd5
8r8Chmz6D7HWqugfxUz2r8yuPR3aM6/RlUVzfKfsyNgor1RybJWDR6BNEXdq
ZPtYLlk7kGlpQQg8HfD8ma5OKo9tS4uAV17gi3Mr3jhri1L3x5n8lpSG2Ntg
KA/LR1Z1uTKlmn1chNeNFijKExuA6BHc73bpinKmjd5vOtB0n/35RDPDKShl
BokBLzX98Ob2A3K/TJEoXn/sIB0M0swDT56t7pw1Whgc97TyQlaC1me56bH8
X3ypq17yK24GFyAoOsFZY3uTu0LQ2C/FfWEXbJ0H8UUPn1KFQqg9TRcoUai4
H+dDavoJNVDy0Fg6PSace7ZKm0Kz+8Q/W/u3nAOFVPvvIEht2LxuiEoWFASj
RHY5IaqlwMgiE47EzZFSF+C9GWeAwzEUoEPsIPwbZ+csU58nxzc1lnxsYPHt
hcdG8uqN4YWdbxPh7THJ1of7whUrx9wkjlxn1EsPGydougCbK7tDszyPoID9
gHl7T5fSIIaPJtlxhowBjXzrahCUtndAUTPGdx1Dg58J2cBxdjfGxQg8VOAb
UqonOPq1NfZnAiXO4LUUsmRlZpK9CnN5syCZxFvpL230pJFuJVVRHT1Bggml
8S1zdzxNR098RGWJmFkyLS/ifNuTkBBFSLSBv736D/JPj5W4RPR1VwsFSL//
s/6TdxGyKqcjJ20qpGUyu7ymIiCjt5seAwyn7+suOjnCqLL6Nx6vmLULOyAO
YcKvMcXWtkqd79YZqlnjZryE7+x1NB8JYL7/atSfY2xY6b9Mz3uPI7/w8Zzw
6Xlhqqvv7D4dKw0TerehU4BUwrryjvP0Lpm+48LUblsB5zPkJlrbXb1t4d8J
AY1ThlpnKH2DMYGDWFHiReJCI9hL727GGOn3b9aYgBCQc/XbWHxjnUgiBEN1
oecwCpqhsNWzQX/I798E38JskMclsDSJISlCu5QmB6m3J0YlH0E+VXkuePEE
4qH/BFU44vun97K6tKLWeGB84QXayeZNkJeUGwymOdSUdO9j3HePNJMZYJ/u
IhHDrzF0erKpCEMDHCTxI/mLnqtFDX/Zov+cLrgyNXsZ0TFc7ln46ckXCld9
NkMmrEUxyuLgRejrqooPGIZaFdEmSe5bowdLTn8gui+PV0XOBgCTsvfLvSrN
Oi5SjvliOdsuwTJc4DlJTJO9t42SoacJYWy0CnN7fNlR713kRh0wt9tr/oPt
7JKb0szkNSHdbS/snDE+K+Kkp5QdKc3jS0VwLE0zYGl99YCfQbNNLawkQo1S
mP3BRTigFYuIPo6Gk6iqEOoTYmqJZ8+3clpKA4odOAxqQYvDe/acGOm/Ucko
0BhvnpRHsM+E+ptqjTe2WcsxsxG8J4ENTCDGECThxc83TmflTlLWGPdl5XBT
/J7wduMiAxO/Eyk3XKpetwt0hTIddW1rfSToDYO+LVRfinQaiMLi1YP8jc29
cVbG72pHfWg6+TgkHoIp+gCUTUb5aYY3g5L+hiPUHXnQrL5cZuZ2Ya8bKihS
y/JnuRSFV7/r/YXHN+YlVZ4OwA1PYvr/P6IjNqTDixZBMu5i2J/3Z8Sjj5+I
TU0kbQnet6DdjG9Qe7YBZoRJyPyeIr46/UoEXoO70Wb5uCVC5Ells19noGZ9
Aqrj1+NECG/Jg03/HQalSnQ0YdicGKyk/WiidbYdcQhZbum0HA/EmtlXsIzR
tOCUI30ngSfkJ31/V9Qxmi0HaM3q7zbZZ/ZcgoM9z/h9ADlHPk8YmlbCkkit
U4weZFiBDFxNbwlfvHCkPogm3tAeVzn2sfiYdgvKR/AbMo12LAnxaHKjPVil
6cG8TPrfKI5IkS/fbO+iIvSv0OHl/dVNIRsLG/fh7RicjoD7v0FDPeL00fqK
I0I8VVUOMB9x4/Sa59HWs21hrLHMn2grgtrPd8j2s93EE1EjmkmH5E1ccAyo
5UblT4CB9wLWLG8t63BzuBHxkIe3LpM7jbfMtry9uGD+1JW2ZcpTPnJOvBAt
q2wRSvvSW271s3HSXviTs/KVUzvk827TT0KYz3zitx2XHe4PwnB11/efZTSD
XuXpHSwUK6Aj+EdhkNYmCHglMPEVwbjVD+/C4qC9/Bb43JlxojI+CBEwiyGP
xjR4M7gWw/6+COWWOCuwGzm+kpdO3f1WBSgzKGo8Ay0O3SFkHbGE7SRQKMmG
GduxI+Sqoa/Mg1sHNWY3I/Xd03qtuwa3kt7Qh8rBsAF0sTmO0Q9BeulKaAmv
BAyDCf5LN+KXXie0jrlDcSwyAoIUbv1U8SfRHGlJrTbQBLRKF9co27v4uCpr
5RHmGnUZ9/4a1qYLuNs6SIz9g92N+xvsqCemBmnZ1bdWdcpULDUqiznONvwH
ddWvi9lT/PVdELRW7TrjIKwP78Lg350Yyh8iQ1R5tYfBaDnuh5Vs51QF5jtI
IR4OaEoyiX4psug4fabuxyAjV3X+c4fMUGoPWt0JBRjfQVYJSbK8csGGF30a
skELOZvb0Kh1VADM3fusWLMOEdDI8n3eXtsjkgKaR/q3Yc+2GT/q0dW1gp1y
ROQvyQoggD3LJFv4O7IzabOEDI2VuFxSkuxe9LAi8UayPdhENIBFcIGjOAeP
hU8CgUAN5jmk3EpWR39mKtToKeW9nCqQ8+AQ9bgzJANoYqNBp2ymUb0foiyO
ySulVpUB74ubJ4yo+wgpC/RoCQZgWL0vXSaQjJB+qB3BOt7tVQZ0+cIP8OPi
xbo1qgelimo4z/nK7W2pq5dyqyB23gIc6jrb7LRCHdHZw2EJth2NKQp9w2TJ
Yr0H6BH9tl9DeJvhIFpMTs4ZtHquucO2vjRcAG2xDSIomW1kUXO9YyfRvHH1
++zMP/+C9KONa6rnXLwRjt+jLOqZfNr7Py9GT+ShF2Gsj7IvMu7rhxJVZug1
B7GgLJnHKg+PhIWF03AXWbJP2xZ6JHXcuwxMnPdOXiNn4grhpiK7dPUpBQiS
txJOk/MldALQIEthRN/FNAFPGVDgLYmb1Vs6WDKVW08i/p9oyZNLzF/MxRLQ
yF77SiSqm0aBkeY78OxF8bz7L3eTKNcWTs7N86iyyEE3EPIaFG6sIuw5DLxT
w7Wk18FkDg3yAUPC+3tzUW6ysVkrgYQassVTYRKtUhxaB2OxBlrhoUDh6BSn
sg5x0NwZTYRhwYu7mM8YfatlivboLIQaCB9VByZJVGIYdD8tLfrkDmw5HOY6
n6ZJX8EcGnxpbJWn4R9mJ8GitvHEg8o2/nvZeiBNwmEPEfJZYufYSZxxtVJv
l6UI9ynUc00P1GvfSN/K1ZrHfrMnTCybwcU5okAYCX62nlnzliAlZGkkL6tI
jjvoB9tQrSOas34lghQ6mAWDMdoAKy73oYvXU4GsSsJcifPVR1YWQ4Fky+Ok
JutK2zwU2NHaB3UPE2IE2vDejWyySqjMQ8IAAzzqIx/GrBF/mI/+IOi6dr6D
NFt0ZjJZctmp0Uz4KG//ttPv5K2lA15tPpnAhTr2dqfaVF8PFH68fUVom1w0
lKBa27DWNSrHmoqsHJooGnUVcgKjloDk+mB9O5tR70SAA1dGMELltfh4uHp4
Vp1b9mdCHTrWHDH2mq7YwMEoLM0QhZS7aOb+LhSPD6ea/Iah1Jcp9FYnYIlp
rwIiwNI6COFqjIFcbLMzFN9WjXWWD0bzzHzBW9eiQfJh/SAsXTA9DyT7fakV
o0sOvHk2VEgKWp26m5POW7GlX95pgtVNML8Kq0/w5qCOLxOn2cH35hEgQJ/E
EsF4w7PLty1LNfC4rvTdEiZj1LJqs69cTDdOhfTIdLaZvVgApEyV/W2tH1eU
+63sBYBjy/GMHo7oQBtIvC+EF+6agcBrU/3J03mZfM2veSiqShJ1Nl2Fet9x
HmkY5h5G0p83GWrUf/A7arwoaXPt/QqMz08mN3+CfteHbc4enkYRD2jTXUs0
OwE9yfxQAlY32aZ8CXir61S7P+cGmpPL3yNi4PmjSfzmIKIAamDfFjNK/sT7
cDLgN0PiqC9q3gf2GAV72GJrY7+ffVenXx09PAhaWMPQE693z6+y6G8K7r82
j+DRa5cUQIez7ZzZmwZ6fw6pzHoEgiCggM/0VdbUVqK7oOpnlJ2TSSLGCQpy
3BGT9sQ1L4tyljj1UvzeJ53VOGkNhKkPz3fTzrVIgKThIJuIWaIx9xtZgHHR
lxbT4fz7l/XSl/oHum7KS9S9j52oJD6+JgMoknRZ/a3qYX8/MEhHS164fyEY
ozJEwsqjs/mHbFUK54p7q2DNiGjtOSwgfyGr34mh61aKxy76KUJBvtJ5R4qj
YsTs4MWJSa/SK73Tj1jKSNtC3kV4sPFjoJ5U3EqGGXSGPp1UG8uUYhYcActd
39tQHHa7Z/pjkw/Jr4PeF2fZF6GaKKqvjXkbObpQ8/V2G4RHJHli/T29S7ip
KvfiUbM5IPapr1XIvGeBgJjzDafCc8OhiAll7fqlUREcVylALcc1BP3VFxhI
GuMW/shEfCiTQ7HoRWNI90hiqWgZvgCdLaQgAh02i2ZPYnI8enEkEzZO3+4T
xNd2G0sFN/4QX+l/AsiJV3U1icFLukDHgL5J7WybcMc3cpop5H2XM6pUdLZp
ffTWLZfKTvCC/nEJnNjcEek1TrSsUSciA3jIAgYZ1YwvnUkpFCthW17u88wR
HE42pWjufMrLZFpEMhjEmxUPm6pjPS7DaXVh6738B+IHaiR7te5iZGhy/1sn
XO2IOs9TTMl61QxElH0yCuJaUQaRxvptKBJ63mvTmB5lzQa+4Pq8Dg6hNkms
t64DP7F6ikPaLTMAJHc/MdZXPpPhlPp6AfQ02Tb4iNPwhhk3+E1E2t6NU58f
Zka0NSf80EJZjBPkhMpJuZ6+04GZ0HFMyyQcY714Sk5bXN5MFmzPX34H2y6c
9D1uqZSQi0qntKVEeuul09RULXQbz/ZpyE4PzOD1nHi1wa2GafnxwGSe+wNP
569y9hNSZBCet7gDZ/V5dQOHyWGF9rM4l1pFVnCrt2gc5QmUjO5oWILYWM4Z
6QXIcq0+LpQLOA9w9NA1BYXKPVd9y+OfcH0dskbhdfftEtjk47mTe7qG0lH0
MNrr8wQc5XH1VeHxfheaTzqLyWAxLGqxBQ+TV3YxX6VSa6fEj4JcTAEsCFl1
69NF8g5IgM251GQ5HcwASf3cPWCs2oimvRToboG4jr1PvMLPmhIjajxCZAKf
3oqPcUgHuGUF6FJH1xIgkO50oqp+gwvnw87mo47fXk1HTXtRq0p22ky9Ntwx
EFbKinr8rfpfwe7acpi82Mfvgk5Rxu+rSL78HQpwsc0fzWnRFEssjLnuqZjw
xSYerruJHaPVLQFH8gezDUA4tcceXm19BziatY0wQgi423kCNqLJVa6WNAkz
SECkqiZse5cg36gY5ETg+B2745IifGezkJXhbhpBlvkZFWqYSOzf7VDQT3Bf
lwM32CJpVx2i7/zJynGYGgR1S1eccNzWHyuijTYole9z3oo7vwJgh7IL70/r
Ri1Fujlu/6GytdeLgNr514+4rdoXCeUMQiD7ZdylfCJGGHmP6SF8oTSXSL0U
j5Qi6hEvK5FmoyA1IahczZ2iG8r2HljFWXFWPsDCCnBA3KHQvnQ/dQmbsENq
yabPCtTLe+36rI9Xhy6DC20f3rccQXHX0X3wXFvioAhkxYt9n/RmDsJ3Oad4
gxOy9BWvTVTP4zENCiJM7Qg2S3d1gMtq6zQ+ohvwypMDwbVma8JYm1WONqeM
9wRmzuvVgY+UCjEjhJAGlMHx9pFeeiQO/Fema8PNddF/wJA7xksCJviUOVnU
40M5a1OL2b/BZIT2877jrt/qX2bn9bMhbRMJ3bV2I3Y3wbh0sZohaoRE31ek
LnWkYUibmjfBmVjWsEYDnrLiQhnjWxynWNzchv/OMgEOB1X5UkLuMk83bUKU
parxGJalZScPooUiYM9JbaAZ7hVEXDuigGjd1I9NMkRA5DIsKuQxu6MV4JUG
KqjZhfdWZX/2C8cBX4r4DmV2XT1uHpI3QGtBxls5EjDOq2CgkWquxCsV1FPe
h/JUTm0ezfDliVtwO1UYMGXR7/k7wM3S/AQ5DnskNf5Gq0+VL/5PCEtUm0t7
/t/odviYQO1P0vRI68hw+a93Tq5nvmT2IEfhC9iy6bV5syL5Ik5R3yqCTnz0
cmYEZs6m4r5vkMZigiO61ViK8wOfW8cLhUk/0os6uSE0prrTyKkDMAAfH1w2
HeL/rFrp8/aZFbZdOkPhcTMp+cj0Wv9HMvElsdtErgvYF91fD8kB0lw0U4YR
BwBiVId01vq/qBGO2/rCUc44yTaxdcsJIZDhZU5nJQJPY8Wf8JTe5DzZv5Vs
g66HBqomJREHigPcC4ZOy7zqw5ZpGeb7JUaBomNFPWa9PXftJKcbgb4bw8gU
r/SECWHmbvtpnHBC2YBXKEGeq8LgX//ETVTsb35tRDZfstjXGPkwKNvRhzUp
dSRCugPFU7w2iX0jkIX87VfbwUuuh4F7TZGlTKFaXv8cZx+jmQMCVFoTAYrQ
2MpP5/HxyogA/4Vv5oMJdSvbx4jcpl0Yvs3mA35QjBIiIoYdZXNmLB4SO2ZB
f2yAoSSvshFKvnqISnI1I77HAaXGaRDGDjkNKseAvmj47xjyY6RVaJ9QEh3m
QH08zs1hMtxQ3Qfo1J/GaNbSJkU5UCHr/UidzSTfg8AL5FjY9OQ0iGSarOOL
S6tTSi6HQiLAswh4I8ItfAg4l2CnEHXWFaUY2HlnXPr8698ktjpB2u8+2kc6
DugCv2+8OpawJ/jczJKMN//v3hqIijzboBRmaRbSkDy020akE+SUu7+acARF
t8SedurY/c2YqMEVEqFLLa/d6PwU1mepNLWbZLDFmGecrSbScV/pC9l+zkH8
+85aPFnyzR1RJoh/dX6tDaX4I9zSAH5b0TWkH7ladFkQ5x1xJvNT4E5Qfy3C
UwunZRhhTrWBj+P4Ppn+ixsiU2dafrBv/rrIrjmQqKJg9rtAE4Pbt2uy2UKB
Kd0+EAN9vwbvlr3VAKHdLtfwe+PWfdCLfFKcFNgAIlGyeQ4vAWlHaVvbt/wn
NRMPKZE18QAAFtxB1IQjEGNp9AbVvdFN1IN9xIwGvVyfB2ORACDLO43vVx6k
2QEaAH/GaQ6kb+gI5+gZTQ2+UQBw2XrsvBxxN+EMpz88U2PY74XXF0Sq8Th6
aGDqB8mAIT3l1rjLCQkMhJA52BV7kk22OmDmpJena1tYxV0abFMNYILyvtdb
Bd/PMNBVXK5xsEb1KXIvT8sf0Nq6YH6YDIViO6PqM2G+qw+o18XkROJXHngq
yIqHhB/LNiay6XkRILk1Y000/d99eRvGrqqDslAbUyVeFcPkYF7SiyTOGQRC
ApqBztbXRp5xZOCZx2Blof7mtf978Sg9bgIo4LMCvc334sQt+6YZahKs2r4D
yNx+soMPrWwRlIKkNXzrUwRazq+CipD1RraURrtOBYmtCPCAGenu82i1N1ym
v/Es1MZ2grePTBPhloxPrZk22DPNQ1SJmqsF1XyVtyBVrsAbmvpG8c4xjSKZ
+oEK2byjHEG9JdGIVS+f2KsYJU6k9h7ufvWm3xIGTo8dj6KEUN5xAJdO7qqq
Lqs+phRR1AJF8v7gmJZY6zy4AV/la5h07LGy+inCiNKh3DM7Bl6hsswEm4G/
PNu9g2on1jk3YX1ULwgifQoZDGY4VswfthMlUk+tXtgMYbWGVvFmoquDfSxm
gFNwP7T8Yq5DbD2ajwomp6hcv9cbfvL6QTCYPlaKGAR2gztyU2Uj/6xSOUvY
uHk/TaaOaDDXknFVw+VtsIwrvlcDnmB8MZTJI6S+WrlExnnSce/xC9hNDU7N
5BbKJB2WdGZCCLfaOVIyhyd5vw/2gcaPCaAJ9gQpllzLNvB51d+d+xG0H5MF
BruquOa4W0C1E/0PTdGbD352Y5hAbORBP21EZTUKCX9cE3v5jjSpvm097wUb
5ig5PLDRLvp3oU6qcOlBF4TezL49ulGAQBOOmo0NG91CdOKteO/WMSW+jW+y
Np1gzagHa5P+H94tT5yjXqDkDLW2whDWEpdyYWs0KXIdaNAfLZUq1A+E/aJg
iEo/AKLJ0GNx7k12dF7srHBYqp60ffYq98QyAGxo22JINCdE71Eid4lSEg1i
MkckircFxL/+G+ZGETtgeisp5iXbreo43gQp77CFCqbJiahKc+o+fahdK2aI
maWBXMFqXgCvVgaLG2Z99GsbmnPrHewbOO8UTWO/hcp02xkb4E8WHC2A7o8w
FMoMNnLMSIKyFsn8d9D1WExAB7G1n2gLq+EBs+FCTWglIryPq4JtOJqkMsFH
CfQalaDcmFQoGg8H873dlrkD6SEX+u4ffOh9LWaMkFSOm6HDrJGADnO72jSh
C3O8mbAFrSZEoePW9IO7+UbnkzHEZvE0j0qx8iJ5K4UpQlnp+Og1Mss3w5KS
LjS0DO520Z1AZZX3CH1/dycHA11/PGePDvHF5JZQ83Omb/HWAdEXMIZ9Og2N
fGevHbNILAV4AypVPSfl1BClgoQNjJ4OBgAyx5yMNDzJiQ+/FOISaaYJnaJo
YmXgIgKU6MBquk5LJCMRtXmK4wG18RqFW7Wyn28zxncqo85GQmbII0WkheyT
6v8VppT8+WfUAEP9RlQhvKaDOz85vT9ARYijLyWXYbowF0l47W1phO69oDZ3
9pEU4c0wJMYeHbPdes1HQ+nro4uejwOQb5xlUvsJ6Yzp1y01G030FKk4AKB/
jfgZbZKQtqAWvYWC4r/cbCcjENBg34rLsZxba+r+FRUylRyxFl5XIIg6xmly
9qs1r6zzPNK99OZ3YotsDrIytYH7kGBGM/kF/2+TuzjZO4NE73JCDK6N3YGa
IXKNAupa549/uYr8l9f1jJwfZEJxYCvep7E61SYFfUUyipU0zw6fER7j1KXJ
0uxSFkNlsCRtZGbu/zs/YjadqY7nGNupLp8NNVQq3sAExrrx6OPJi9Oxz1IZ
iuSPxYHRhICMKyD+9EqGZzuHykWCMtmsBhOP3Z4znWoxq4QBOZaaAnh9HO24
oQvaMWDwR20sja9cAF8vZwm04WCnISqpOH20CU2z/DWwoHlkJW4cfonIydvf
B7WDfYfVtXXaTpnMBU5jqJUbBaC3F2wRkdnB5qv1ywDMkPtCq4PA/UJKfXA4
CazctJuxknV9wGlVEpcGUxlsWZfnByjDl6SU25SSmRAKyCjB7xiiJ0i+YeqU
xFG88BQdfeT+s2l1oMcbY3Z+kl5AYvmDaxN8wa26BFKarnn9mQ3lnSertduq
MW/F2+mjE1WtkbuembwUeyYsg8n5qZ96tdFfzK+E+hUM6yjlyjO587BDhx8l
2SZl8IkZgcabEWhmjmfTgbbpnDtbNnlH4KeAjpQKlVV+JCbmjnWPnxFTVap+
rq/Fc5rnY6VLWK9TFkA3ZaiSh283BrJSg/p9iyRo5SAf5mJL2YRk9q+oAzUc
yMI3UZ/5EFsbosKFrDENs70lfk2jNtBFrNRWgHBKiltpCQTvGZwMi+YZCsEY
0kXILuYRwFKY4T42NoOybtuwyRpsGSbHZCORbX0AImZatCFuRIu8tbe6xYck
vNNv324KHZF2LL2muysmYnHqhitRpc/VJ7Udj12QSCCU2k9WmSyM6tepIUNt
CkfVz8No20N9Ux39gTzUPyWKW5HBQmFf/cALr/lFZY6O4svrA6oT84VaFw4+
cnt5tCngDtiboy2JRwf/JeWJskaA5PGd7kWJoypOVmbvaRNOdofFLT1qKcDO
RiVvUpWeat66Iq8k6MtAs+JVg9bDuLO5Yldw52iQZ4J5pNLSSq9VD4aFpL6Q
ISOE9qFDkj08K70uSsKjVDDPmi/EmmMQaf8jLs/C0eOsPDL6b2M87ceunX3l
rQfflkKHI7YwCcQJJhIbyG1GsCJxXgpVcGACKZZzVbEQ290qlLAUxmLrkOPp
p4TgTAdPZWACK10vMl+gzefGugmwbPdfGTNDCc1NeK8gqCsM0qRQ6Ze+FCxv
VGYizmfF/S3eyrppoufX5tecr2lB2FHSrqm/fH6T/imj123Ss7M+SHhvzt3B
J50XULK+FokoDloVDHokVwt/9RGcva0VoorKf5aZWj7MkA4UACgUZTNQ3P5Q
2MJ7H1ViStqx1HmPXk3fli/2m24iVly0l/ga+q0n5OBKTSSN/yUxRruxjFkE
xPBoqxpgj9ANZ0/5HtqUudF/vsa+KNfIh3+i8ptIlQG/86ucSs13DBeB0beR
0SoYa25nJYu2oWbNB+ak06qPRXa0MHzKr7r4+e/lGq41QSD4MkKw1pTN1RTh
irXCuYvjZpMpT3munepJ7L/Lu8jm7xhKfyzasA+lethRG6paGIbMgTDOwPV6
Rk6dBHsVRYggxhDFwGMvGpBfgBBWHi3ORVdqb+mvgmEiitiuxV+MfpZoXk9a
tisSgnD/VxnLmsZdwAlNaJoUxSn8xnHMaZHoRC+U+F4rxewzRGBZ6+n1vpoF
EfAGQ25JX2ZwcLxnKs22QWDuo2L4YOX3+2RsLjH/fLoRmZUHn2U/96PqIGVY
C9sKGArcFEGN1iahkrxuL3mn2YYcFve0k4vBvjjxJv4GdgK98WsWjpwzNhA3
Ej3DzWPzZ65PuG674SRzFIxC9t7gPZjMa7SuYfdSeD7NsCc+l1nHxyEtQnta
RaT9CZfcH/mtR0SjMSzF9rLC1cQxWD93zEHk5lqOkanAAEJvhPJeiUg/vt67
HvPbhnyUn8vJVDOuTpEJQtknzRwHhsUZq430sVV6VkS3ZR+I7Y+bkDK8Wic9
dH0rnOj2mHVT6U4/K2CPPm7mVdY3pU9le+b7/KZeDJJQlFwxHpodedvwOJFO
Ddme+jwSpvI8CuoxS3gtTvVu0RriYEA43FqrP7o6RsnLYDsiDRp3ihWTNll8
c+Sgs2+n/er3lXETwXWvKBXbs1wDRgofAF1YREH3mLPZSAxxRNLaQWkftshS
UXFrHoflPRfoUQr5VoUyQO0ZqO3CHzaHmQ2ps3fuQB0exyZX173zsgaaO7F8
DrESsICXTdMvhe5ptUrrh8fTkBL+uQWLsbbmXjdzHGUW9Y4WMa1p9Uc1aj1u
8m8XF7K5xsXd+6RiIKiMlJ0lBezic7Z2mvvm4qOydf/r68is5HVG79ggZWOb
cY0CTGn2X/ek+P2Gv8EDoBcsg/YhMXA08+wh4Ai/21ilEuVKS2hFq4MH4sEj
mP/beZOA5c7I6nBBvXkI1iJmL01kYrVswTBcveLxfe8WJqykxjSX+oSr5dFH
t1sYTAjZ1VJmG52C2MG4bDuBBKyTavQhS5qlfJtyYX/ud1wVtT8jrwdHsv3K
c4uy+s6ogCP515Lxbsn5PQkUXB3XIS7KDiE5KIEegCk8pC9odsaqLJmzaKzb
k+NG3/ebrC9is7sQjn7Fq0INwNQc6I1zHtf73np61eYzNHDLBhy+QJbwyMxd
aXtzHTqER2u9pFtmM7knp37NYJLXn0ailaZNRbV6cHGubVTytbfFBNdKwTHp
p5G+xzAzIIvoQ5FzmmDHNTVWODlsEmjvdN4FcDscndue/iT0fHfaKAtbOpmB
zPdiztVsZ/0KXC4HFh2YOC5ujOl8GyNXXScs3RwBdYv4Ig11sZrGJ+dhz2Bb
jhnzSVLKq/sae/GOjL7cUnvlJFblS+9Vdv/nzIHYGlth0gVieQrXQryvgmeY
c3ncMeC2tmisN7fkJIPIbdVHmOkQXCxmTPAdC6QmPhwmPYQwZ+vTqk7BqO3I
dB0ix0n6M8sXNVgjoyQw6+JrgQBWXGC0vdRCgCveTk9eVF+/5fn9EQfcwr/Y
LvoLcySCJhiBFHweZ7zLghAKGwYemsMTVSBTswm5+VTHbjfjLeVpufChu4xX
aihOhyRFVIO765qFEzEqBveaFW/x+YgDx3puU40/KyuYSKBsA0quWh8Nov2A
SAnY1Jrg7EMl/V5erXxhhP/q2ICQ7AKcDnR/rT1m63grNSg+ySSru/CYktiV
m2ig52myas50GJlCjIP4e0026qxCZEqbdXBU204i0qRK0ngDuUK7IIFUV6nV
iEsGYND140szEc4e+Ri343bZiN3ibPvpg9rdEsVMN9cwgx09hjDZzNmCOC61
eoLBx3jooAvHOmGlRXAhU1TI6cq11QWeq7mQ3U2HIjKV3Yze0othgoeyu974
IVvLKCTdCbl7jfOeMAPDNjkym2eZr7HWf2lwaunjnr4rK8mYNTi2f1EHBSU7
wXiOxRszc7FTgu4QRLT7EQtDnY1emmfvBPRMUgNdaEVtxMAN0ADdNUjs+Dbk
/vvqgMkju4+dqM3FrOjYmx216dLpRUlJ2H5CKmziL8WSQ4IyTcJSl3yWxt9g
3LbXbicAYgybHqyNhUMDAQLISQZg3VpwwrVhV7PtMnMRIIJy36xjnEbNwN92
dAhjC6zvtCNKiBu1jPV33S6/Pi0xj+MCQT0qtLmoeaBt7OR/pJt4MyBtznlj
ThJftgHtqB9RQPhfwd+1nZtuaDA/80C2+D9bH7jzUW46zQ5o8PDgcCaWIKRz
xBY3SRl/jtHepgDs2WiQuQ1pA1cn50LgDUBUFINboRvwCmPcn+uoaV6U/tbV
hIXaFBej2NmndXp+nKx+Q85jqt4E8pMC5BPNRb6gPoVlu48Ou0k8wT6iSGuF
aWrvZjZNk0fqkECQ48FuhZSW3cfM55TAbL8MfK91AtalAV4G5FIHk24/jzcb
dyopJfJVeLCRF5GlgMOJ4lBcc1/ltRaPGgF/MRhnX7q6iHGToc4UMYXgZP/4
vB8IGOBt1TfzCw7zrCNMBM//OparUDF3K9XVKe3CaT8t2F2m3unHYGpG3Vyi
5jVQTaGlq0dSwC/mq+XndywTYD0swspVm2Zjfi1564aKXLAeklEW6vU7sTM5
bXZxolUw4oXkFx9fMGv7dKu/SmPi/7aSoH+YolyHax8+Z7HfVkUIswDQEOm6
h24gbma5vSqm/NTIZe9vbY3speSL0i0De70jyVXGjGMSYphaNWqsbpRpu6bk
Fu7atbdaa/169539a16051Z8EQ5/xxLqDbFaFqgpkMq3VqqWJgobwA31666R
f0sdQBeaIAwv54GZ/HDjXyK6GNGhzctzDscSokha7m4i/PbivDG68q6oGAKB
0AuMxjpDfe/BcFSyYnlf4Twa/PZvltVrNJQQU6RPxIvet9RXDd4h1D8M3Ygj
hPbvoZDTquQEQM+PUDSJvrki6DHXpXjWKOZogCPa91GEnypu4Gp260Jh/t3v
5dPkAtoWJSjS5IAF5Gp8BhHsg2I9aeakfbaj5wR9zlJsuSN5axI0cEaq4pWz
2O8u8Si9XmCxt8KR3sLSAGTGnuMtbmafFa1KCwvaOuiJj3C/w5/wtnPOMEe9
lptyoutfcKSWqZgV40UWvWE2ALokQDrLL1KEPxyFiYMe+4WGkpyToURND4gY
dlR+L6pFRScg4FGjiqUFzDAy5FGu0nmOB8uWbYyway186Qi/fDzlTdSK87Zq
rWuwYc4ZObfPDI2GI7jTeGn1pSsAoxAufpPpc2F9OD6W8zHlQc9ZU1TjXwfn
ojRh9AUMtl+cA8k7HlHFuWhioRw6VkRCVuh2CH3YzT0jWdcihMQSU4xHiKir
K0Kqvz3obHZUi1I7SRgWfpQlPg0qNaO5r0PtYeQe8T83bD2wbJp4skURDXSP
NqOj8JUWQ47F88MWFG0Q7+swMAdBHSFYi2FpQSH8AAm1c5WAHsUygtgxqhea
dnr46kJJL6xmA667/zUJVs0ounfYOm6JUoCXVlWF2nKP+b457FkAxBu2UAt+
fg+i0C6gNegQdda3ofAHrHYLzScwn+OvY42pcjdR+H2jkeI0ESP+BGLkEoSx
0tePoyjkABb9zJypIYFQEjq3xS3aA1ky8qbmFV2Fo27h6Jc5shTy78lF10zz
3aNVdKHD4fO2zybfzNQUtjs+l/whJiz9XCfqPMSWh3oPBW0KLN1ZA+FfrEG7
6pW+a/rIKnuoWDNt11IheFC2KLCvW7/b+mw3Fs5iMyDmrUF/sb2kBwphKz6a
KuG18hdyg9tFLCFqlxjt0OpvVyZgH4/+gNrSjWWi7jlnWYl5xGtzofe9YWIb
sQTCgfTU0EuCBpi8Xp/5Re1sY1nxff+5fckkBdge4PJLfzpTRTlsonUK4eF1
yEqbLD5uxhSpKIN+IYvjvmRzwlc4CBA85klbVvNVbR6FWgVhsIIfF9mm5wlG
1AZXl9HT+m+j2II1myR0Czx/dH+J+2DKpyPeI8Ld0ZnlG4NpibbLQjJP/RLW
SsSRv5uMbJ3EvC1IMbHHeFZTm8HOf+DMGaAU+zqAesJNKP9/8YxzgDtQBpe0
4EAcqXVpD4yITTk992r4xsL1f1i7fsI5Kzuj5kOP0DSrGe6ESFjng9tY5oSf
wTqOcoLBjZrt/CYdgmkTTDTCyTl6VhdHrOXLTlaYZOnHDKx/q2CjAlM5IFEH
VcrjtLKjEJM585MZQBjRo4HzHKV3zLmIjYlTKz29E12JaYdgZLAsU5ZxwmyK
8q1kvP+W8ZZcmFVUwbnA7sSbAF8KPtI0TX6WB0Dp+iORWzAuL2VYj4btIC8w
eS9U1I21y0M8JgjHGgmZi0BKJENCgfAR1WyXuDcrvkrxaKgC1QkM0F4UARUT
mEb1q2sHmuz9KnMbaD9gjpCh7uK7CdKBDEqwFwRY77QwJ1p4xfRHUdcYW9OX
8rhMeS6bPUACG1ZpWYS7J8Fuf0+hilVEeDNKNITC+ssE1crrcrCZnQR4Q8Gy
391j6bggjx4dRvxc0i4Dd7RoFBQWrCqA9637R78fjHMrjzClqsqaGrrxxHR5
mIcWVUrrJc09YAYgbQm/LJe4IkMi8MZUhFLBM/bNGZmUModbnQs/lEpekzKK
DzF+ePQyMnue9LROiHvP7NxtMxbu9dX0/+9jlQtBLPunKzD9EmhU8yEe3dVX
a0KU+VGzL5hdM83/Cz9jXp6TZPSDLS5NEJnmSHAMAjABUZfelNfeiwFpwJlc
EKkQhb/nNSpCtC0171/k76AQvcnC9cjIGNDvtrpl8W452hOIfvwIabZQU92j
W1fWCm5FYB6hMk5d/IS0223U1CcdM1hGvzazMXIEslS4J78x1opW+V4UwmFC
rpIulq/K4die0F0l4cPpaWOEaR/AmyNmD+9CMV3GV3UiKZSdZctse4E6ZzDY
WTDLZVzKDvoQDl2LXCwt+DgOt3jIsIU/Lw0mCCEYv5EgoZn2dX+wVP/bOY8S
ASyNge63C/+N+hbvCDzUuwiF7sEYaV3VKxBcE4BEQbYZfUSoHTstITHM9rHG
WX99V7mVFcUQuVLz6m1E61NoEy5i/i9YK1QURkuYAgC5L32aPkLe6mIPT9Xb
l/YcIaL15tbLTGSq2HVfzNL+XZMB0xVscWLBmkIoYnO6HnHdRlGC34Ops43E
qxF53TS2sR13uaHl41Wvw0bjPTRA97VkOAYWwYymbHadr1a5qfxC46zvlNkk
nnywVnHVrKOVyExN2ytUbjexSuz6N4O3le/2zS8fpkFPI4K0SOPLtOiIqH2I
0m38qGzWvrTB6IwyKp4WKA7I+20WvSK06xxxSpGgb7wtuQqApYY5HxzwrHyP
Do4QtvHJTtqYZgCBTffnp+u0DrvXvojWqYWrRt0gIcZIynZY3f7Q3/Iuzssc
757wXNI8ssV8z+2+aV6l0Olaw+6geLuFyO+0av5HOsieIoDliLC67XYlZuBc
Qs5jmbshMwJSC3lRAW0hzm2pxdMwOT2RcCounaujpDz7Z1IKktbsvTUMK2i4
juxaBvyWKx+MaUmw7DSTpWcnOQ8PSGwLOejllWdMY74eVr+xhXi1Clz/6R5q
pBsVmMEX6FR3nDpBXR58XO3bdQeAT5BXD2bjzIDIJJ1VyY9qjW26eDGnoQkr
p7ailQVJiuX5WABpGJzyyVdrBkJA+N1b7atvtKlWdbiRJy7tqIGySrkSmvXj
Lwv3vogD1s16k+423hHA7vk3Q+w2wAn41PwJ71t1X5K/v1QGjnrAc0gj7RdX
QpcQPG4vNW7muj37w46ZavbziQHz9jBJpCsMhqhhNK+vzYbYOlHedpzqU2F8
Ju7Q1s3vIKQsalUmCKfT4ogXTeNbO7g+P3jD1nJcg3CnFs3whTWlK/LbBYR2
A2qgwXAfBk4uuZ9iNRuafqe97qKq/ZMxrETcrBQLRI+LEuKx882VlIn4NW29
y6i+da7mpUSFcS71evyHb2tJVXa2Q/Q7OwK2DvlUNTadfifu8wVWiQyzmq8Z
610Gr0IK3yu9NWlCf7nQ4YGbxDDfSx6IvubuK2P5XiWaktuZqUkxXfYE8+qm
bPmSnvmR3QS1f8s2qNmA3uNS2ZrFKHZOhejbhmi7pHDFit2KPtpdxKp1Wcd4
Q4NbJChxM0mB9zIfxfTsiMBlAGyWiaFrV/H0eAkpWME/UbUeZpcIid6GEG/H
uSyun2TFmMeI1+VXBrDlghZitmM8AF2e2iwDWp3ZoAT0fh8HK8wKDi/I0d9K
KFDpIViwXELU5n6FCVpl8l5f3+zlOAc4ivA3ovKuCJJmDmTr65TXB8Wc4gJT
5Uv+ODL9WFt/Y1J4k7Gvh8BqfQ4ng5XO4RWLLqd60qx9Za4/QqjtRrwXzMz1
48K8tbWuGqVo0NeoTrxtcPyEYZ6iYfHQRGQGfe39acIRcaA6wV18dIF2Is7O
by7ruyMWFm3kEit8OHZZKa2C4Wn5moWfV8evjvLDwSazhmZIU9sYaFHmFmFn
SF7R0g8VWLFYfqWUSbFXhiiJD8Lbk4jkc5lnC33rJkVMHXMXOOLk7htvaP06
WQqTb0NQ4puTlnX4hV4UrgDNm71H4/cjtSsjyAsNIQy3rL8+E1ydqJoN7QrX
GCGs9Dhb0nVBnDVLU2Aa+65hzUanZgE1vYGLsBt1cLyL2sQxeBGoHbFbFKv4
oJ1ufKBcNQBfUzaEbQLgc2m2PC0YucJNjmzITGecWgbKCkT0sgRZ6Ub9hHfJ
Rvs7G9PVqfuY6ZXMv0rlgpiHtCQZqHrCn6gER1RJZmefhHfTLJlzdPZ+9N5Z
i4vM07sLJr+sKeP8VzJRO5xr4bqoio5zNYyrl2vVf1fDhgUPsqLG2j87RFnb
ULqOep2Hf+ShlHlXMjfgcGL1A/pUizKOLXcxj0Ge8LITdn20UGMVX6oZCWaU
L7lKOWijQGE2dSJvInQXnehd+xCFZQpHZCN93tClX0MUCECbRV8OiVBKipr2
j3ciNGqx4PWocdJQTgu3S+XtL5p/uZvhYbQh6U2ip0bPRYNDqLJCH07wHr1k
aIxxkW3e3LmUxxdMu7LQnrqa8vFnikv/46lo8ZKhHHu4pC2C75BC2LVmL9aG
oUQwhjcV1j/1pr9jq8Pla3Iss88QGqyUUo1JLRWPEcZGX17KOe2gw86xj1Xr
cLWwe+H9KPhih2sc1CzgY5heBPKBhuJ1sCn97xF5BG8F2VMqSewJHbD3LGHm
AgIPpp2k0PSSay3lfMnlLVOLoH3KzsaMu0WYxMGhaf090aKL3yzVfDTHrQl6
+8ojG2xfUIUz29zTYImK6i+GkrNUgOuPny9xmn3gnSFVn7nPd1bsM5nY7f/t
NBSMZAWNh5AVupvC7wPobwdb/+mqBnsqrw8Ozg08Rz6AN8uAX3Pp2ULLbISe
GdLc/Db/2LqNCRdI2KBkBVs1GkIl5oRBYBhvautV7HkZGCDGoJJNXuIrR8K0
qbxtmFSKDCwfqsod3Fx/r1ExohPVJxYkslowUbmtdPw1P8PilgLqwMgP19Sp
uCbr2T1C5rb+QrodzodQk+N0JVyNI9rAkf6iJKfvFiI2XcyGVg+PINF5gW/g
Pk+aiTkxG7zHdg1UmBCKbAyY56pnd9x1wTdVF3S8asOmEaBw95LuMkV4sb6S
OU4OT4WXEjneNnn9Ue8/tzB5xrHFoeveoUZT5VXQd1ZdcmpCsCnVpYT9Ml0Z
HkwVADsZdUxAXEepc8TnbrdMJQZRdOzooZyETKMVotUT8aE6qlblqQQZAvFE
MRXGiigPi/ox16ssbzszh98prBYiktyKPySE0Pcte+Mjh+Fg9mQasZwWE/LI
LRqW28J9nsNzMbvp9HfS8gcowAeAQwpNAOts9aC3l52EBykbMvW0GX5jxIR3
XRiGnfIJL75lPdiv4NE42OgU/V7HI3UZKZy/aPOGifxjuptsqUlUF5ejtJmM
j77qJyn6RqJtoaFlIhdNBLBpIMpOQZqnhZ9iJXlXjODYIOTPQg8BGNOCeAKr
R50147xVtcCYK0SF4MuHRrcX2GIP/FJyTREdoPDvBfVfPYeqbp7SMCEdxbz7
R6i9yfmV9R7q2cZHYeRb5b2QgdmML8CWNBiAs7pcjeLj3MiV4lOku2aCjHmn
1lYtCi9lQ0pSX2obVL4YYEY0JWcpKkq6MpLidr4R+wD32QT4O/n/SQUaC2kR
rk77CHsyd20eG5BuZYFP+qBP4hnt4S7CAGGaeTkexgTcpjIp6oqbvlS2Efz0
IfBm2WK8I/qSz6feS7tqwLuRwGxo0Y8+loBF5k7pX/btvjh5rKtNKEOQrzHS
3hatEzfyWF3nk76qqLVwHCVlNIycjo4hut+U4hStDubeaSiLUy3v3kZA3s0D
K9wTJEIi8RKKej+NosDOVP1QzY/UQs2Xxb3KNNSVxz5sgTUgIGo1XHom4saK
TIISSK4SGvXHknzbHTyrkjiYzpi/S4iRxgz13png/mjlzTqrP+MTJeVWnLNh
5S24UG+UpwWakMO6ouxPkxTYKqTylt2k5XjAFRC0tddMNUJyzNaX65AXdOR5
YiHLhuEVeRTBnFbumieh0d92xmo1TbOALYX9k8GKXCmhhym7hBX5to/XAuem
8Czi8fxoEt8eIoX6Q/a7GFHYjiITtEZTg7Q0xvg5jJjj3BJ0HXuxdzBjgHLJ
Pi/dm41VCwAmPDKFo3JBR4nlejkA35Qhg6g3DM127eQrsk0X4/O3HNpdhIJR
p+Aj/cfBOBB3QZQlhoaAHxtSWCWoqA/gAPTthIAHbCg78JJ1fG1vPG4ISkhN
YRbUP9KrUYN8Lmcvuq4CuQQYbqkToq+qqdhQFDqS49hrvuWboMpP7JLGfwoi
n+qdgVfeme3DflDxWgB3+h67l74klGd5xWGqfrjob1A2Bss3EwQ+CnVJM0nb
XQgUK7zuQxKY7ckpGFAylO7Igrmy5i4ypxeN6NXRaolxJWXveM5C94XTelum
Xnw86WgDAM73ckbbvndQGU4MvXFRLT9P9qA41hGq5te1xNslhyohUb3NfU/Y
70fXEthd3HCZKysI7P6T7qjBhFVrRObxmrtXh2X4h3tjm8Ko++0o9zosfvNB
KdiA8q5mx44FVxhupVlvrpWPp0UvWSe2N/4Vs018uadiqacbS2+PoKIC4EFA
FjbRurmV8k0RaNG0vA4eds2FsNfvJMZHlH69Ajep9GU7YtHmdHaNLN8LbZXk
r/B/+Ff9LxEO6caIBWxjeSrmgQXlJYU9Jqnqx+gA5bFnKI5pe6PqOlWMObEq
mYTa7GgwVzvzXRusnWH4rR1O1VKYky0jOTV7b4pRYd+UQtyeMeK+ArV3MpP+
6T0wT5SaOb4EWeHDsNsPm1tsfR2kLwoPD7bwDM8kZSRYL4WvqY4V71APQj2v
FBISFOUfQUCxNQWKbCTCvreTpBREpIVJAPii2gok/sBczF25HugmQ+Pa2bE1
IThz6p1/dWWzX2WMZPo+iT91/SXySsNyvUzigHyEZCeJDTn9veOB+H6mbCY+
JLct+Ejh1zVjL/PAV3sbYeHLItbMcvTBHnH2SjMrS9HIlSXKWoZYUtFfaD1s
X2jWgKYILqTe1sUQZUZet/hFvUtwagdy9i8z8ECMP/YFP64xhbE/QkG0OjTl
ihd+Sd8Xfy/Yqvf/rg618O99WtNN72BL2HZ07LEwL+9Tel+BUo8vIIdCqfPY
b3OeIbH9vf4YjKs5SWFAPjx6rIJ/Uense9+LMRHar3DPeOLGpwRsiGQ4CsxN
jrjZWZQAyRDXdBkEsgwpeI637z+k4Z2QbMre1kAWVhllXBaFiFZwzAAn02bM
8UJee8mzh9fky80d96Oqpch3mLYw1groJrGfWnQ3PDaPhg1qI9xpxowfa9KX
pqp2xx8/618dwFZV27rR7BEfu+rbfJ4EkchsCuVGSiyFmBkwednW5ZFwS0PN
efn5u4DlrflgN/SBvZEg0J3TGqJ30Ky4kPgPXXLXk4Ef8RKOQq0gPfk5/W04
TqB1gwE7AStCtUJsQcEbILpMMgasX6RDv77J50zwvLByPREODH7dMZo9yX2a
J11wI4bCDCwH6MyWELUpQC1wZ9CzpZSWk9fk0RKENlpJSEYLlSw+n0t9wtCq
9eOibNj3lzJ0E7w11N0prtOCMkA/UE7H7mcq/Ywy7G8oPJMqqhYzaJe2hdqC
2sHzvRaCDDlHj2UtlNEnLOzhooeUoWxjyRj1VMFsDWtSJf+ktBq/6MtO27HE
gB489vA8JwS7V5u+TppJjscysKJ7c7yiiEZx71Jj+eibFoOaRifzqW3ep5WV
0fct/POpLdt6BQZxK84qH10AEyvYNTb4DPeuMRKZlb1STaPr4BkjqCKfC88k
wVI6cNIFiSVh1gmXEM+OU/UiSZhhratUoS/ksLqoxuEMx55Ls2A+Y/KD0zg7
gLW3uwASfkT6XhbwmgAANLTda1ZpAt99xZuXEdKfqNWtr1LLpBZBA3tdz91e
jAY7486cU7qTew4H6lTXs0jaCvGULac0m/kzBV9edEU2RJfgpZcRL7GauNZv
9bu3M+RkBXfKc/+gC4HQpwJ+vthiz+F++uYsgAVww0o3gb0KvHUX5mrH9XQg
LnwA9FWzzxfNjvCUVRKtagIEQ4AS/yQ6yPkWtf1iLFeOEaOaAOG7JV38Ah9f
GUN0NBLStFbKU/DOJVB3Rx+L2IoUGD8hqsEslUATpiLxdlERlZOKx9jFU8Mq
p0/xsCqF1YllDb8Gr1f8M6xg7t7G3MIDoe/4zFAoyMAmxIp6+QqmYlFD/W4n
X1mEkj3KyrLcDRQXwPZh0tHhEpEThgzzyQr50luEQlEsT1IqHVD1IYp/cQip
cbvuxUkcfZjm7QalMLtBXr+BNsuQF9dsSDhVermZ1jBSgoYOCFFPXmDFwJX5
I+K5IDl0qG7DOYT5V67CBlIygnVRaHFwD1+KZpUyR+dZREJF6t+euVZSE3IP
TPhwx/qm/Z2B4ja6SmsQqcF+j7jU/C4crGFSK+TTKQBt5SZYZnvFtTWJPzIW
6LfrbI8qyEv4Gj67QX8gAZ8WuwqeAkF3YHf4VlrufGXY9ECMsXLvXpfWj4cn
hRGnS6i2YHYd430XkoGKLOWwNpYVkpNk5s318H/qkfNr9fTnvkEjWhhhYk5M
gxEUnvfEpvUbG043pUHbKwjtwmNJYw5oFtmqq5bvSJzF7LzwOHeUhQCb4E5H
xC9XJnlF354rq9bCwCx2v7ag8Nytn4zFnKa7WGcSMlHPqvbZeTvEOqCu5qbi
0lJ2JXE76vcfdxIhnBoHXPcTbIhSgYZfCsvK7nT7KBKEy18zPkMnBc7hGQTS
rrVatd41TKoB0ayb0cCpxzfQ8RzsP6WCRaLaqpyOHXcBlr4kWSk2sP44Xo++
7wNaSVe0fAkpJkKWUotmzyj19Qen72e7U0rHb3a6QvaYVaJhz3Wn1oNUhyi2
MDNFN9TOq4SpXUqmFKJLYueOM6p+rm9sd1XQrZyHTjDUXBMjDbjUXVEkLzbT
dII3BCz65qmPdaqgGCj6mWrAqy40Urlw1rfs0b1VT72jWUvJmhePNRjxyvHV
5JgBfcpt++QIR05zLzeeTpWn4awCRt4B1esDGJgDOzu2+11OtJlnwKyYcK/P
xcFuWazRsA+JlymWSFwjEyh2Pir5HqOqqJc6CEkMMWZkjUNCoFKM9lsKnqGK
wXdy5shugWuWeHDCV1APAMMyOfNQ3Y6QJ2VN4Or4pwt1VMKAA/QYsFICuuIi
vemFVZf2qYfylqdtLqE2bCNRQTZl007cw6WE0CyZJRcoEzLGytpqZXAf0Rcx
aKxGvn/pJnWMbyb+/lKbKgWgCMHwlAaNYbYhrxk9Ynz6G5b+7HXZDZAmCdH+
TYhhQ0oDDttPzuNgpaaiADbzABudWGG1Dqbcmdfe1Ye9Nr196vMCxo8FbaSz
QslpPTc1aWvHMsHczIPy1x1EwEZOxY6xA+jOtfxR30hztO8yhs+Q096ItBX9
9dE5zpehV1/6WbDrAPvJJtBJbLrqJRjiKF95djczPE4zFy0ft/GJ/1JrjVwQ
JfyEc047drGUyhv0mrLlAqBQhpfNSy/WsgvL/yM8MdnMqI3Ddv4hp9d3Sj3y
LjS7l6mRepEAJxpnAZQBYROXV809JHtKxGA82nXxI3JSNY5BVjLb/9xukRuc
Z3BWXqgrlIHWS6/NunNZb+B9eEoVLQevOj3WMb82iyyDLTlF3NrD7V7fAAbQ
yZWRRfGPU63Xg/Mmh4qp5JM7jdZqVyn/uSAvzTr2FAcEFre1bRqHt7KojRNS
7PaW0+Bq6+4EdCdPpqu9WnWvXnO8C4ARXOkaLiYyZSVgX7IWBmA8jwH58Ucs
5ReDidflVge7G2ZfjmaaPDdbQ7VAVGGL0rsNgbUTPLpKlxvuUH9aS6isUt0z
4Nu4gXTFvIsuDH+azsfZSkf+PfWfvivskECV7OdvbQQwMgOpoGuH5lsnMNwb
T1lvN3WfHzeFvFZLPxjfeDLhKEgTJuk1ZQj7/arS+abFLWF6eGJQ3MAapg60
Ln+yJmXkdO0Us+I1S1p6EeJM5coMWiqgVmdBEGAimqj23KYRZGelexFgyefp
I5pKKPN7JfaNakJXH0h3nODjV79WVRmozujXS3vTk0qsPhQ0ghBlqZz0jKWh
ly41wJi1G2dErcfvVzeXFUS2BZvgJBMde6IjzXnBu7/RsGrAm8nvNbdThMv1
CEsh8qNo++QADlEmmPXNjKHifOFiiD/iFMSCEjwNLQIQHe7aNGOYhwybAfEF
aaNgNGkzczzJysrB6UD5/KFv0daUHU2JsIj7swSjpVImvXxkvSB88mjMYGUO
4P84w2N2i6DAF3ItO5xBCAyl/ulHpz76lvEOGp67246K0GIZcZ/hkLXoCNUz
1e5LhIjWFkZHL1PEggIL/amAlgeNDCKaEnseWAyNeaGoBxSMPpVgx536Lf3g
Bmq1eES7EQK1J2yZJR9qqlxuLqnssf0DHZISWvOoPwabI3ZqXaMjQo6Kn/ZJ
GaGPhO5NtT1P8NuVvQw8+Ch8f8m+BScZMush7vB8O5vhFX77ks8kDfYVIsEH
YtlPWDoGCKgR9W7XET5rs8/gmNk9okhmb6sQ5x9FgXZXhTiIo3TN+p7MEzNq
3+MIawJGCTaskKh1wWRMTJSGOMDvYDkVF5WX3kh1F2nvf1hz6En06Oulk4fx
UAYpNc+97P1EwERuuHqpKWAm1CHl8aXTQHB8BK8Zwl5z2olz92+VJFaVwKFU
m/vHOb55PyDthCant9ES8zgeZ18hL55qT48B8qj0BIS43zK7XcLHXfKDGT/k
OS5oRBNCR2P7XNOaAqPFlwS/w1IrE7oDzHYhTEnkKXoCGO2zFq0r6RIpYRE+
gYacp1qoWKmPkV2Kw6cLqIGukIiNXdzfvViNcstpKqUYkwx/A9rXVfgi9F4o
YffX1xqxNIK9F2a5QThxJB5XuoOr9WTjh9Zc7LotQDADB4zJP1u9WNWJ9DRR
3DAT6Lq1KQZ5JCMM7DkeWjvJouW+uDu04gbBS+Wk7V7YHlaCfcH897Kvx3MY
EeKhCttmM/8sfDy0ACO2xmRrgHnKGC0kQrF3qh5k4ogGIwmOWIsOPChZrFd0
IVDzDlJzpE3zDczucNK47OpyU6N4JrHK4JcKoeP5PDYHWDHRTlmo6+lJnxrJ
l1vn6cENFhPpWFgn5BQIERAPhGnfD3dMWBw+TxgaywU41zY2mdvv/HL1kCPx
EXdbU3UeM0j58eA0WWMeixFVVmFIbnn5NEw4du7hwCiNIyivomJ1ks788DsQ
B9hWJt+8DCXjpCUKOidU8F8LZclKA5WixlmNRuZZdrsbPO396idl/WGcn1Cv
7WntanuSn39FaSO4MrpmUDpB3jlmX/A+Dke2hezR3aRzLF91iPR6gKRm/XoX
pjkxtfjqL+LoLhOP6WYJ9bihseYF3LU42ZuxjD5cp/bDNee0TbJexyRlY5ky
3/+aQLoW8W1+xNQxm84AJ9vG8E7ii0rTfpKNPeca1sDAdXEufrLQRo9xovGB
sU8Q4yOdTIHCPJwY0V6HdbGzM0uyIXjJ+qT7bKJeEe5M1teArD0Wdnn+f5er
DK/YEN/VEn1HgtbR+QegdCaI7JvlPLXDiUzWea/Xm6JMgNXlKSFTGX7CjoX+
ZAdCMNht4QwlnBkiKa9zAkQRwgc2qvkLC5AUPaNw3lXzikWYdW5R9C7q1fMo
81kje1vwVykuEsi/Qiphog9ZlOoSS/nUTF/RC5hlfJ7vDx9K11+MoWLsY+Pm
okR3WBxaazXpth/9XpoyLJ03GESRAX1EVvqX/khM8sGZ0/Sx2XoXr67YPi0r
Z7+jaXiaZYr6ot39wBazEBIoqOaKI7/2w6nDZNgXNOTtdF2+vMUcpup7On4j
cOgVzNyk9AHyiXWu857co5dbseyByzsSD4qPFapJ8fQ/FdRBOdNvOUKIT/5x
G/GixKAlbzNJUwyCb8KQ32ln4R13SS8cEJbnveZ47FZyff2ZQOF7Rfeo5FZj
e5pcRQObbF8gVWAJD5np4Vlg7LE18da44YPLsGhOtwpBUwLIKiaS/lcxoED0
JJCiasF6b3g4Jna0VkUEdYKlGCDWkDdkSf+v6tX1NB0U3oh1vmwHCaA/TCFx
kCKKD3Bdnz1JGwO6hdQKaNly86KykongcaVed2dkvSLkAD7AXDmxvd3MFmi7
KU48Hr5a+bPOS/jzy9xIDoRculInVHC4X4OLO6EA97MXzmp/BpBoWcEJoWX5
ckuqVjemwG5UDoYEfIQU5D7DUsjrJrMOVHxNj1CzA1Y7tJz+ixkr/1/f3pJC
fxY3m9sd/7QQIMsC1dem8n09yNZm9kzdjAvyi6S7HI4BFo5VuAcyEoQKIKyR
vEe50lpaj8NCes9jgI0Rpnpg+n+hJYnV7kh3JAq+y8K9TkRBUiopBslTZWO9
E3Q5YPCtCoCLPCPEB5P04yYf38qLCm6jYso9F12EABcxaZNYKqVl/DIT1jXz
jcle3UcIJkcUJsFh2wMUVqEUIVdR0RC0ZAkS5g+XDS4IKG69Cjjk6ZsJr99a
UANxn8wlijuizte0i8jRuCL46LJ21kFBOwvC6wdpxNDrT/RZPskS4LoQQ62w
H65bdlp9fm9z4XL3Yqj3ARnosBu7vDkX8vciKGKBS11xitf+lK5R8uZ2KJU7
7KNPhoV3/TBIpzTLBACNao66KGlrtwtLkV0sTKkwejKpQEBnPfo8ROyvRQAH
5IZgqP3kl6cU5BWFEEqXUlD8eZtqEkmYt5LvcWSJgZD1iEa/4KBIqbj+iEBn
U4xHu4n3LQKGcMVYXuh1DE+limDAeUT4NiJjQwti6tf+OH4z5Xg1vdEjo5jA
D7HddQ4jr6x+U4CW2ZMLy3ygqFNNZutP0uNkWo3PFNXZ6tPEthehrXx4S8kq
25PfavxrJ2g+FvSSF/sI7nre5B+HNOSh5G3QoPGs/GeycM89dLHQXBuBURB6
nk1u/YqBFEFC64cajVL1SoJsbxrw+kPn2pdJgCQyeg4Q5NwVONJYY4TGgQgR
ms6+ZxDKOg4Q4EN+BYCghnLYK5VpVsKKd4brNUYQIDNXt5+jhTcGaZRc2UpP
mc1xBKemP42gmJKZU6c2wrv+2BtmCsKlSuoILsJaIqMfEqQG0MgdUn/iN9HG
6O0HrWbcYrlj4BttpLvqTeGL+6BRrnICTEOiIK6wbawDYYJq4LQuKR/P/z2Y
bluKHrFkuO6SRWMi06FPH6Xt1Nu0ooEfKY6TulUgclS15hl7VJCGg6mdmbMd
72Z13BK9H00t+B4EEWxSJTyBzqMizzRoFLpDU+KDQpt5yPYXEdbMHEPJyqiJ
A9USih6LdoHlDOy+PA71SJRW7S/1nmTOuWAGKZ4MJAaAguj9TwNG1ki2IW5x
XubK8SN0a8wl3/PV4de7ND0BeYJAxSpGyioNWin+hZTgC52G0Q6hMP1Rpmin
OT01IjHMrmJC1rdF9/gJg7HC5PmmFgd6KOVsO0LB7I/3WMuY13X8ifUAW9FC
obeqpXhoSNTPwR9XNta+yDF7UFegVwCpBm+ZJykfrIJcychlscwvbs3XRHvG
8TXXpFvMjO3TjaRr1hJQZp8x1nftFrZghjuFMTNbcD8JHfXn4+KbdCp8W76W
YdJnoJuGtH4Um7jXXFJjlWUmeUBLuVHbZSMkIuVdBdqcr6MwqsJER+ZBPRxe
V+roOKrw7qsLI0pq0k2ySJSi10cXE1RHOZHczfxegU/8h5D6Nwu7zoSIe4Yu
vxkIMv7H/bXWcJ109W/9lmWaUjhu/2DjWmkxtof4eal1d0e6l4p74SvFO6dJ
HW4hSkrxMH5uBrnqSjRpgYqi4zdIGRHOrYU7f7NgxNiwvvP8DmK1sHDiwNlm
CFSBnBNaGCFaK+TLGHrdA5J6Nw27vU1qDwe/SVOsZ20o4pmilgNM4HW65JhN
ot4bBF3LMGjKFRCve9McY4UV4bxGLq0wJa+nf1I0ZE+TFzyCbbQGu0Ill/j+
D1W47iHh7wB/YncPkip1f4ivRRrUmR2Ynn67X0QuwOTBown2z/Q4rDPm4KOp
tHvGKAkuwDFeNnAkBzB6L7V8Zq/H15RQ3ar12GmW/l9spPA5C6EOaW3BjJls
fuc3h7ofxAASsVAnWDBGV+94pWT+4fUEGTFS7XhE1zAAeLizigLJHqoyDElm
k5nS1/wgJwL0qgHgQM0WgzqFkY5PG3cZYywIwctJ0AOmTWBriTXN63kfWCmw
8SGq+Mo+0BbV5UPASc1V6qrEsg2AK7n0SHJ7029I7B86AO6Mm0sf0XaIZGyz
ERV8BII/ItDySDVdqkuvdvvIKt2ma0W0nd9GUNZBvNepNYUGqbUybONvdZm5
iztDEhXlDpqb5+qmguq10y8K3zkZQGZah0G9VDA6YImejM2PwaD6V/owNFh/
ade6KYpbt13AGuiUe6/Vmxgx8HpNAgvVpfuaYNuKsKcgRpSwh6PSC9bTrrjp
kr2wj1wEEoqguvbn3az0FksMmKwFjbqYHmyT5fQQtCXINZCCpGn2YR/3X1kC
SvqaAtk61hKZ+l+KrYZCextYI8+lVumx00tag6lZmIGty1LbFGKHuKZ5CWI8
a1WhjAkLVIKOYtBw59e7TeD4is2+7BCb85DO7P7jTqNH8jgbxXwwgLb05gou
oU2751k6+uNi4R5NQkzeLIH/lind04DyCe5JuHTga6U3icN4/5jL9o+0RiRV
QWH6YHD6mLAREbv8C48+wYD2lB6MzHbrOYPlkCsy3CfbfeYaBJJEVTsvRrU5
wE/qx5TV/pqKCDAczCwqzbxJEm9Do8o72whHd86irR0r1/Ai5QbLKokxvkim
r73FAhCiGmLBNF10fwqGttPhk56L5VowMwmwt0OqfeXnXmZFH5JB3W9vV2W2
IwT4TWgPwLx0HGUFaaztlh130kTS6CeNXAW7hAfrmr0MhD/LAyvgjsr5/KiY
Tm1x2czvGWHxEr5oAVava3CscfZJ1KJ7NWj8Eo20XIIVRuynpN+pySQWeFsx
f6fM3ACq4Y8jVQj+3HUFQnx/SUTBP3TqkSSEGjtHK2f2YdG/6pNy/jzT2tA7
dA4WGRIRxLSpXZ5hOAtTNTo/z6p9v0x9hfr1fB5gt9w90weY0Ny27PjyxuNC
V8cd7C6PKb0ne2kjKI6+4N09CTSK7ucw/j6GaVhD22RE1RIAwYesXSufiB8P
ZxOScCyd9nhNbt6/QyMOLKEHW/PRN/8bjJRNcSm511/+OlTqua7nT8rUcXtv
84Nvb0HkhWF5o4zZ/FkEyZXgZ6M/N9Tt3sfEGCHQ6MY9h7fuMwn5L31/zSTe
uEGqziPIqNODqRyXP6HD9hP4cXOcQr6usEtSsvhZWmczlGucxg6+DzL/iizW
EqT7aC9y3KSuO9ZanGOpdaaFySiB92l3mOayUobNZeZU273x5mgnbgmAnbCQ
3JFGm/Rg4DRAZW4C3LNePsXIB6iMBkHM1Qm5QUaTRB20hhAf9Z6hDxapn8jS
luFRAGdlNAMW8w7y6mJ5oN4tSYhjMNvHTib3CkVkqM5fdjNzPHEo73cxju6M
F+UAH6pI7mjrgllsnKO/8yN6TiMeUI2atKoKZlnf8uxgsaeLpG56G8+9ezx+
ekGiZXuxeAl58mHBtI7ZCsECklSFkCle7sq6oHlJL4LXve/eIWORBVX/gbge
mTHmu7aH5mSDwM2jAyQ+GnhPPXwYWXKcUJGAhc8L3+F25W8ix+zEgeGLkQ3y
BuCAbgNn7udrsrET3cENt8Hvf4Cv4ivFtGQnH7G7bNzgDmDSEc02GtXVdQm1
RRenF0V1dn9iVu7EBQ+UNCY+QbuwcMtKo1YqEBKWOkq3NROQUeD7JKkMDCNJ
SmdOZCt+fmcOFgsEIan13/v3mj1kmfoVNC0vHY3LTwZf6AWrkZDFwERVJXvr
C7///TSRw9uKowSOjrzx6+EqrJT2U4gYHFSq/aL7dliGDKjGzV92Xq7PRmOL
PD3cEWy71vLWUwUwLVEIi2JC00Jo/ziMUtZ0ytQNHLDDNMXigIp+09l9VmMn
JDVIRzaaxwsjhwAfh465cQeHqqaoq7OtitKuO3oF0GbPnVjRHnuBjNedkw6w
zYIquBD8qCxAq5h9dcK4cYDkmnIo9X85TwpaiDunvRR2F4tgPq5MavcS+GjF
WSZPL7r+ChsYITPEHcmzKFirWkIhOH9hes5LPHUzW4NGSP5L/I7xYx8bjuwd
clxibRubYuvNulZWChTSxymcDKJkqtW0pIpYDhkmgF7IX449JzwvSqAbXZkd
DN2Xh3DlBAlzmjny39ulz4ivBKM+oYYy3nrDhz0AvFci8yeUvC5mIUEkxsxD
hjt/W6HUs8TKTR1XdRrT0WUdDvnE2OQkyLAX/I65HKYN/pBxivlEvkcYRqyE
6GhO7hsImkQMuRz7TafUrdDpjiwiYn/uYR/VWBjXhbZP06pWV9Kbfmy/Rjt+
EpHEvUtQJ+GwNSlz2zGDLXbvvJu6mzcHxWgm23koof2gN5A6MTKp0H/Mn4EU
LXWHTjdNrdvwGOHFLkiV86knAdl3QRzfQzhDJJriJHQCTsLV55GSLyRRlmiD
ELh8cSOgOeeeiG7pYYfHZB90VHXC9ius/v8d6dEhh7OgBorDB9DSIOZpBhLQ
mnc5SzbWcmQ0U91pBOxP5e8dkQYua23VguLEGadFIT94F8q1LANQ2ne5RRMk
J6Vony7c0eA4IrTI5t0yGJSJVGVKqgX+jznTve2A7FYj6mitUT+Cz5W3Sl/d
Nvakw7OELy5ayvGmEPVm8Wcv43hG+bLFNlnpDEmSRUdc8w7r/pLL7+2rCI54
c8no+vZpn/09QMSK71eWBquM7O6LGoDIAm5lFSXl7yQgSECrmH776aipSZUw
uHKK6QOM7u0WMXfumtHALIalrfSk6ILtny+Tju7xqdEAt5TJtve/Pn8Yadje
j4DbniJyy4UUTGi6vlwyyA3Xiax55bZrzpNBJoKVfkIuvnTq2ivsGVJwx2Lw
Y6nYpWwRTPJeuS14wXjtcBKEl4iQaD0pumZWSmJ4RNBaw8jMPLZKgFxaT6PQ
Qig5RYZwbl47aHBHKKnIQxM9sSgw1Cwii7PzZ1QQwd24b016Exy6vKfzbvy3
tRgqpw3zhUzu329nIOdTomdi1yb77aV5e1T3JmTePtskaLd0B8clNlhCOiyl
qOnKS1vAuiJcpkycSt00MbAG8u9f1GLdJFiGVB+28NLjq93gJfwGyB6zQip/
9aEHL+nCQaNPe9uQ5AcmPcrNke4O0zVCzNaVerPmU8ZdW6M6nC5GFzYaLc+2
RibhqvHi9byCQw067c5m83weKoex83wa8AlI6jrdYSxVamFPtwXlTMYSyrHU
i0VA4PDK/H18EZ9RXVuoXGwNoddGcJGJevWa/956Z04lk058gZShV18Q7+WH
tlpJwKHmRhzxKYlSjdlW5EUxwugiJzfCfViMFQaoLgtWSMmD1Xmo2emckEAJ
4XY42KUh+v2C4N5jCN3Yo4hn9wh4POTaN5KZ2G86mU/mlXhr38SZOxQx4HJ+
vkc/It2I9LA56/+XsEAjpprTinE2QRSlS+rxq/mgeQOdFzLBW23idTKkTtYN
VtZaW7S3fN1loCPSdTy4wMJ17NRfUCb4VnJNJkGPWVX0nR655+L++gkzwSOx
JRyfklWS/VDSoYUI2J96FpGppiK+Z3zdGUMMl4m/Cbbt6d/0y7m+Uogysvui
Sb6LRrFI+3nWC9B0X55yZZx6mB8p32LBtoKPB0BXQp00CrPKmB7KM9fi3AFD
w1v7dpmb30wGmyich0OFnnGRl9gSpnXP4m2hpUbYjLGsZVnCstC9e6v0xmJ+
0lVhaO6oY9rglLos4GonRsOySKDnA++P76EcQ+I7ZsJeaZkq5NIwDXuHn/+9
2fzoItPBeG5pmUCb2sSXA2fO+HuJalWhwW7Br7O7xbnYgWQO4q8r72Q3EAlA
MkiGDEF0zbUSCaQp0PIQtHmwRTK3HG/E9Kp09BzNurPX4Tt8rf96aI1lgoXK
lV4ZCKWs+mzYDEXo3f/Ncm/nEBLw2732ddrDqSk5TGG7dE3N4q4ZdniwXTur
Cb4LilXXXuOEhs+GDIV/nM+3eAaM5rSG9eu39rpSLR0M79VFlvlQR7Us3b4V
DJ8um0RHNjRPyhayCFVef/oS75quiMSPIlh2U7hgVsd0SEHaqJWMNgJLkj/5
Eskml5zAAlQuDXVQ/WXQgthq+sBnqc6WlgLGHUcKOEbKJhtNyYWAu3KvOw2u
NPxuWnDxlWUXxXiL9jbqa0RoT0Ooo3HrK+wQJFRZN6Sc0S0RFFvQvRTLXZHk
HWRM1BfVzu2izD/GkWMy4GMT7u1wK54eouzB4q9HtLZb2A23Zocn+eMcpTuo
uR1KFfTBOrjXO+jPS5oqSDyASQS2DQFm5QO7ywSf3//QSUVq4Km+J6aEhG4j
1PGdzOBdtUo1jLlGJ7lc51K2pSnJn9EViSR4W6YuJbbJOv4UoUXhxAFpeDXe
sApwZdWXjj+CXkB1Xm8LwoKHGrAfqE1oF6b13SbvIBBl+flrmvpRyodCog59
BNhjYxyBMgVWqurXWcbuusCGIBE0rBqu674Ly2pFYRO3nuJKL8SkSmF00WWz
7ASy+nAMoMooncW19aPExw5GfQPV53DENAmxBXISfnzF2dq+ZmJKtLVQN1MF
+XM7FTHVn+6gPPveL2QujDZzoTM/BVofhRiAiz3HjxGiEZsd8B9R0Ohk1AJ5
uELPcSO92D+EHNn+bsLAGA9XNeCe36BsXqCJFEFQmTjdcMzhFPJuFIX84ypt
/oXG9yxCFoh0NvzL++nWkQ+cjL70ilXVY0ardts1AWgjYUYkOjV4BJs11lUU
cFFYMAyQ/DbFVgfZ6Z+M6Q+RglWfunrN6GCHrBE5VuIXD+s9eWnzjjYrDKA8
Ys2kM7CzkQwI/K+H4E0Ywqbw6oucgxHiK+PSQ917kITGr03AHxVAwO5//nib
SwZDylXdKkRAB4lahDq+zF39CZzYuE4YyLS5iQnmUjPlutiLw+VXNJudUduH
GM4EQeTDqy2SSByv+HmSEHOnDUpOzKClpvFn3Ued/bVvuz4czWgkW26w9waA
IzRTkRPI24OqcFp5R3caZEdYjgDSmfPyt7hxchPfrwNo4ML74ErTYxSFCePv
XLgNsZ4pNL9qfkmYhX4RbP5ODyjsz8WSNHpS4/f04g0cFy02fepj0mS+5v//
o+8I7IeGaWvs0clnK+gyI8p93bPXbd+j1c0y72CmvxoeNkMT2X20Uqbd1bq1
EtwTqz+WEpsYvANcyPtLvxJFSebN4FGmctymI00WQwzuMdvaob/URWjghiMV
tnA3eywFSimaizoajZcZiVmXXnPb6Tn7Jp866pdNU3ZtzYxTh9N/f0TZR2S9
fzb/TEKNt8dgtPNv9EDBSMcjcgAnehyo6c7ceK7ZFlUpufQdSE+B8mEftqWt
euqnam8eBI1FoKwq44pVN95WRgRFFLcseq9wF0b30pDuf+UeeeNeHDUU9FZY
cliHYFVZEzKYBd3maizy8C1DayuMOi1FJVYGdh66X3ojk08LQ83Qa0ZZpVQ2
1cSj1+ZO0ahWL0HzvB2aaB7uF+sXukKIsIr3N28vHrjA7E+vrCPd7HjYNqsc
FHd2uA0juhUIm3ARDrrVC59miP0r+tX9vf0Bg+e/SQb52q01lXAHEKLKqG29
pIqnKdyUO+Z6H0SHkw+bMYXj3D8XV1JCSJz1Ppz0wM2jQQQ+D9GD0ukwzpbh
8TsGl7iV2IuKZKSePRM0XH+7w2laqchxUFDG+GjKKnFHOiDo5AlRyaRWVRc/
dy0Fb0YBP23C49+50lzMFxjtglLppjYPX2+iY+FpR6gQWqP/Lh3NKVOm8WG7
b27nUHdJNDVZQ2HYZLpdvM9dxDCxVx5i4SZrxuTUNu/9MqWteX3wAJ43YIB5
Yv2NiniiZf+ba3a5qwdISXp/0MjvPdYbWtDcSYXs3qnP/toF++eShK+1P3Yb
MHzyihMuOrV1CejoPJsIVn8m5rIGzas4BOsUlTorjv4dWrTKKRr8CmNoe+MV
sOdJ6o0Nbrg3UPm3UfnOGKmy9UZeRV7gX6hXaKjs+/sOxRSe3pzTWg+gnypn
36M4uRrYxtXSsQglueX/qwtpynyenuckOGbQrxkBMT2cVh+vCSkqyQK0EnDU
SuhV1nBZObV2wHJF0lppvBlDohcrq2+o50+G8WcAvUdrBwRBoS8T+XOs7TV2
9Jn7AfmVXGeu5VAjLXeiFlZGnUt5CSrBTtgeC5MBOWhjmawJ1wn1azxF/QOe
a4d4dkX4l3dQQlcKiiMefdnVIJNKM6c8GqSNwd5xTKg2PapahHEitRAVRYNA
oJ1HMGXtxVaVvm91dw+ZnJmtVJ0qKcEZAyGzbmrvvQm/1mHgxvR/6kSXzTIe
dQJSUTxxoVez2pRe0esjErJcFh9AeOMJkkaa1iLOgCjtVWWodnn9J0xc4Z6f
0wQyhyAPXQmsOrhaHlc3eCEPY6Nqy13S/Bygr6XQcnhmskDocqI0ja13KgaG
5otlv/PmL66b9/CLVU9ZeYpai4UBWsJSntLmLzt+Jpu3WshneIKaOLgNs8t2
QfR6jOm7gJr0b+hm5LWkVbTPsCl71yaxAg7X/vHQoQ0KiQ4Ahr01Ht7dB40y
RhlPFMUGQO4qZWnepciVkPwxP2YmDDMIykgkZVBeODFnQLeZQJelf4bFRXtT
UMcOojj6sfY6RAPVBSaws0wn3KkaWKgB5kpkEBj9JajeBQeRz5xVYWPCf4Ag
E1zV8dQs+TW6AEDiawDiT46w3uL1uS2H1xWneyI/vgXSYpfZsVD/X38NsJqW
5Yijtkxib8E9Xg7wA3mV/8+we4RBTyh34WUv5wGNdLd1JEYOV0wXdJIrZypD
Bs0zZn2OjKwEIdpuYfOg6eBFo3KtLj3955DEHg4D4iYCRr7cOzymzVfDediN
aZ/8ZM1WrFBLdsjPfA5WGdIIVyMsA0nXIAArFyFrc+21CKYWnqyVzNTBGnmf
2TGEFq1fEIMc+zMbHYhbM9pZnZhyWZ/TXXZNPn2Onj/BVMqKuUfPNoW4AyDm
UpGoXOvHu9j5lXzfDWQj3qH1pGw28it/4e4VhIZDcDOqU5Su4tmEGVMgcDgm
u5LhFhL6xW7NysG6ntDYSj3DCguq27uHI3p6yKSVd6aWtIlashjibl/ESwTZ
lRaYL6UTNo9/f+NNUoFtYi/FgyMTeExDMJMxS/uBdr8nupSfO2ryHrZSvoF2
qecLmKejDEtXqSzkRFHWZHJYmg7cQNergZvP5xX8OEIaNwpKoZYFVf8BClF+
behCOFXt5DugXVYakEFrIvfe1Byz5KzWAaVBL8xyCAS2hX7E8lhjbIl/YDPS
1QdzfC4hsTk9tl7io6PXWHLVJhkO9zL8hNWaXsKnTCmfw03qeEfvS7K2S8gf
3HHYYFe/EoB864caFwGzVS69/LwPy8+gRuHHAS93TuOQ6jb5UDl4NrkcV8b9
zRPQagMCPh7A+CfTRgeueiP6pEHaEd3whWGDUjO525/KZwMH86Nhj/vB6IhL
3X/JTmYOml3vOAOVaduV6dSPy0eKH01mqsATj+JFUh9/OPHmBoNlsqgh+EYJ
PffpLrHmeYc0QLhu51TuvPjEL2yq/1+DTAlVs5Gs/eTI38PZekCxhLJVWM9d
plZmwLgg2mGIi8eOCfVDbphitAOyyGlTP7BtY+gu3me3Bwm3TqFywuSJBxsX
epMXU8Lo6VDv92szDuIBBPlazJLTTX0tanEfS6QMxArSUWhVzD4CIojhUwWP
vmwBNMI2+Zqlms9AF8k4VG9h9w7Eh/FOSzLN9DfuSb89qPRHXZtzyiquuUPM
VrtvjADMkXStPc241fDnmKDbcdRmvoau+o0gbJGaEYhCwsNLLo9fCGPompgR
OILPmhFHxs/mhthWY50E+xKXi+3BeoJbPVqLtD0K70bhF3ea2oZ4PYLIjxMZ
jGIjCxd6Gyt1tMZu5AMdJ9JMzELaTjRrY59Aq0oRQnn22inVn2EuTOk3Nd5l
EZp0rYJVfWcBKjU/a0texooxcaaHBoqB2elycgZvxNg6N8e0bOkKDlrrwGs2
l2emf8Ky0xYC7qZE+X+obhvseOdTBikvfGZ6sGfFZi36DoE9caSKQ26+0wLa
t5cR0LV9xITtQGPzp1smtxvfCHkZFDYO5wIc+fBwEDZHVsq5o5fyxZ0oapCx
ao8KMHw2b46G+ge20RqcySBrkOvLdBgH5pqf/ClygoxlAAXGEoU8ljj5T591
h2MXxOT6dXSZrOcSly9C/uk5twChtj8C/f0jX4zO3fwjZxzDSVN5QbefuP2/
tx/S9I4R+LMauaXMS4EKpMqurZWOGxoNy7Ng9Gk5SxWPdSTMQvB2dSYMMkdX
oEqMcQWcO3QA0mWp1oeREGmiaVpc+0enQG6pn6wLmrDx5evNURXN9OLwCyWl
m2kCxMFdYUCAfS9H8PaPX5kB0ZGn4bBtXipWBhHUaf3vwLaW/0RZlZiin3Mo
FVeTLbjml7ctcM9z2swFyMXBt0fIkGheu1CuaD8E9D/tV8yGI+cBlzKQzeLd
CbtarXtapGx1WPwmUHmiRy1VvvSALNwlDDw5HnGiSongY/yhs4r7yU3fF9/8
qNFXNCP2zbMJ8kIlTDN8x/FER+U3Ny1y+rJiQRyGIghdlHKiDBFOygxGdTQv
F8i7sDhFZEYFPyTO0g7t42B0/BzkSVX2e9ikdO4Oatf1Mg6JFjKanfV34N3s
BPVwQis5i8nCldrSlV3vcykMrfVtcS9nHA3FGn7XZIfQ9SIe41QnSZ5XQjsA
nbYwdy/PV+XuAJUTT1w0I+/W2CLl/hWdXCAOD0Xixa4yL5owUK/UPyg/kKiN
Fm7WGlJh7WfochQQ8UkPA/wDz9Pal15+HWZam6X6aMbw+Gtn39pzDNh+91Y+
Y6y4DtaINWaifCNYZJergVqSfj9HEtmoAL4hF9p28q4QmPHEapZ/IJiu5slr
fTL8uOdViFoqyUlEPx1Fg8Z61djiUiB3VHCw4Htb/0dB0rgxwXzSu2WtnIOi
nK1oIBgzUeuWEqlMplWNIgPidcGA9ZnNJmsNLuVdN3CjKse1Gp1bnae10ykq
8HSwIfF3DScm4LvoI7Cw6E4VNu+S9okwjWqxvUxaEP6xSn4YKstszdKBu60U
8gborz729x49sacZOS29Uay8Xoofx54jOO7i68aEL7D+7+9TQb/bdIVqjfYa
F4F9Rq3KpDEEvzJ6WO5KLTWcLpd8Hejtl6Q0fTOJVBY5nmLPuD+2LUOuWcUi
Ym0TFV3xkKxOTuVJSRIfcl3cIirNl+GDw8mrXzhx4XIdkWCPH7mOEq4gSuuB
fOdzJt8/ed/JcmJibNRFeSdnTWZRAPH++7IcN6sADkgDYk+ewpcvlk1bTtOW
Ub8TfKTNGa8nrLgpQi8InSI5v9TQRN9T2pVJqKdRcT2G3De/TVvIyLBDKYQL
NDrc1MrqwUaBuEZTIunqszattXYFOGQRW4ZlSpuGF3v1SK32zHVOIRLcJnfk
aWXEB6Xciy5Fmk17coUdNe2wIjezMbTZzWhYb6VivMetRJCnXLAphBVKRBr0
WJ3/GFuEQ9ptLhWfAeUZfO6R8FIeFEPJ+0swEE68qed1lyNu9yooz6dhMU/P
OqPxCyA65fVHnqoJ3ZpOv2Bae7qqnl0AcRFlzhad10R78Z0b9blu/QaGFyw4
yi4wS+GhT76d8euvvwXdliHoE96gt46byYGnmarSMrlBvmReWgJZbXeB+g4+
qtjUZhJuyfUo/rOhp10QLmC1Tgm2ISjKzijm70TdqitCfooms5Vup0vP+Zjw
sweCrPCLukkEDyMMxc77ay+qhoShqJHvexyGUEPC6RKBlWZq+d/7lMIb55pl
oh650jQPPekwXxZQXkJ/6zV97galphW03rZIQ5dA1zRAKsrG3rDu+6amqfJM
Tbb4PHNR0BUVB2OPiqcMMn6lqeyfHNoQ24VktL9XoWDoThwOIz1eqYCtFSTJ
NY/y0NQoaZ68t0Lf4Q5Xx2Zra4BKHnat/MpaMr+SVUn90FV2G2MRUmomd5WS
dad0qKyv2g6McQX+Fsf7lYBbVo3V6GzmEUaHcJr6RxljWzRfkOWRvY10zAcE
/+1/ChGnKVypuIbs9MQYFBy0rMvWLTMQ0KUmknzPVenmcnKgNOrH0dKWMaqH
6Qnd13KK4cYAbSqmcGmoxbXTDCPXgP2eEgy+X5ol4l2ZKWSSqM6rwOKk0MPR
UVbO0dW5TxR5r/YTEvryOT9m01gLLAvMUkGLTZR1JFhZDeE/jiwfqFQc5Hla
YyaZ0JZ6n3qEKsgFTwIVKzLdwo8A5jCXC5qO4fyJBNnFMcf+py+2Ffr9wGJt
iWNmUfMVQqNN02s+SMdcig4OdIP1u7HYWaYGoiGgQOMiBu0eXpwLKiiPbP1e
HYR40lMe9iulop8vleoEo4p9HvRKiB8cnzf9WOiRSpP2xozGu7kFl50EmgoV
yfhX6aaL1YO/BhkPiB+mylzk8cshyRmPCdIJodO3m5JNKwjhRClK7NQ1mbdC
asMDb4B6+pQxPYams1xusUlPHVBXbh/GDdfQ3BGZoxg9JRrJeApGACFMaP0j
pjMjCYGyv7EUCFZ7jX9tuMKoh56Jl/1KEQEjZs6tzC2fGr+QPG3E/dqQTosg
s7aa7CIkycnGFaZJSo1kSCAV2YOCylKkN8wIjDXh1E0mbdVF2vQewNDkIHd3
uM4b18evin1kI4sLysg2gay7y6G0bLE1e3xr73GMMp7onmgsw03/ebLHzuwA
0aiF39AtTaYU2Rb5Rocbc+STDtXhu0w40WR1pU1MWjw0Z963G35cionuX2Ti
5mdL6aSuvK4tDqjdaPh2VyixNLF8PXw+kN6Ft9EHTu/BNzmtSTM+TMSfolwL
wHHY03viJBnsb8tRnL3DT8MYbfzr4636r7Ru9MwLuXkkdyy6ZMd+/RU8CE8Y
RK36ufqY72/nTMXfCAMuSpfbSuXHpHBMIPB0IFtOk9AdR8v2zWQyV77wwobg
GB9VF9ooY2zvEz4EybcCD8Xg8PCbd2VSb6lkfskeW6Gql2KE1wq/OTjNrDBV
jQw13ASHHRNj8C3PHGZpuBm2OXcTYVmkB8g3ubSHbVY10MWrNDzaM3K9Spat
mXHbs0p1tE4LBspCzVtKQUWuyJo30IAvoZFYCPEyZBHwTvugXswpRXSqIXZE
r9kUzg+pzqqd89G+8Fd2ZL+bNnOIPx0vlH4yLj7DjZOJclY7p4Kp9YzCdaG2
WNYa8NgPDODG1cP4AHAbyqjgjDwbpxHBOJ4RnTMA/Vd6m97gTvgXVAS/3juQ
WEATcRgYToTcHPo+NC1QnDK0Fn0VelahrG/TBBrfiYBXmXjkg40EhIE8HmvX
UPIMobzk5KHpE6+w271doyoIquNFg3zLD+LHNOPdLNcFNjt+p4yKdgxCB1ge
yRAT9tBDgtq5aRBf+AY7yTyNpG/CsbFTHEyQKeCuwYbh4GtS9C4+NhIU+Bks
uE1g2iLI/Szl1rJkEcY2alx7/9bPDHJihAhXVvXh+vtCOzO4F7x+lkWmf5/4
/VRXYgFrIWNsPEu4JtNH8hv6kUlbiqdvvC9foxhYJGdsUYSxA4MiO3OtefYp
N6TL8hptX32oC7DUmoIwh34HwxYj62tUaqRdV2t6RxCFlXj/Y1BwyWllchwj
hANh1U+amdXRJIZf/7TIjMuWB9ZzxYYAVD6z0nypNIXPCwWrZ99ta4bb9QFb
H3uk42LjEbW16RsXAq25F3DNa2hu7Lw/i3IBc0oNbAikh23C7CEH29ZkMN15
H20k+byAoiS1qbxlfshIoswQrqEKats+3eyp3jdYA+LrdUrtlUiXaS6+7R+2
SzL2AXDlzA3tXkGhaFpTxGXFr/E9DaE0dhTaixXLos85uDq4aUT/JEZ9rYQR
fMPGSRLLy03ZwfW0xdDFOBFimZbVHuS3ut37+rJaRajksCxqVHqq3bC5+L/6
YBfdBADR/subfTqfEPU/Y6ajMIi9Qpp/CbMukTVNoE6hZPjD4rAwIb88mlRQ
HoswIa4QB/lOs5kVYJAZfzZR2oZU4hk1gsyJSEdS3gfQtdhji6Dze1qwhPYO
RcpBeKYVypKDslBeQ/imute5rzJQ3aSA7k7vwdmJkyLHprqgfNbqiAhZ2IQg
9DYy4VhyuHFdpDbOwr4hAAa532lAs9PawDpkkBK18rDdiz2bpLCjr1g0Hd2E
vF0WPXvsk5okxCbF6HjyKK/NluH2jicwmxzraGUJ992wkJ20QWN9lJW8Mw6M
e7Wo6BCoPZ/wcT+tbtVhk/bNyBNDeEDsS4HG/qA5c2hK4xT+ju0WNGkap69u
twQVwtrW3eCfjuCAfVstexWuk4Sinay77fSD7L8Ci705V+P5RocuPpurZ08/
Z0l+sVhTub9YRQMMAzyjwnSzMDZ8nAtXjE80NEIFNCb2yj9d2CvXu0d8KqOJ
WGxmL94aDc42QVabF16p9a3ddTUbQsCTc2NfC7/GL8/vw44psSunb4SYY86o
1r0OGKJ/IQ4OFf38t6T4xRS76oW8J7vNC2KTcuQ3FwoAoJqnfGS+H2d6CoU9
GVEh4SShi67TAVJqotNsDi4D8k+SfDv0TwtIkGIXjib7Yp67UB3Dpt3Hqr9b
mz4QAOagAFPLieSD6I3xK1GadduI4OOwA+W1XcowJFhVVWzVFJML0UfB8h4q
ztwzJPstmB0eHaj3fc4H27Qbu0o4EA3xacUN46H+9mXwv7wv1r7LbkAij+yu
53EGkI7TILCuw0Y7InXTCDm52/JPJB3LdhnuHVJfhAzieOtqrmO/o5hmtswN
4uuHzzRaPfuGRNPmQU3U2IGTvyxPoXnfdt8ysjmNt701XbQeIJukcwBV/Ir/
/tHws38fLTd3MhUivosMLikpWpqbkcmNXin/N8pBVpNp+ekk5m8R3kKSCWik
gvVkmYdoUFPVxsehjPiGg7zkYbskiNiy2ONgOMhUanK1SRKASxAGRET/aBzG
lIrG49FmNYEr/NJgnGP6rQRgLCZjLlWGzy6Nn+YETThYKD85rWaxpaKwQTyF
sBRyBorpjvdxLUVHyRt1x62Z2Vdqm5JGpNm3IYcWPXaclqif/BrEiKv6vfVA
VHc/welGoNpWBY/nVR8gK0iV7y1C0H0I2wS/fFjWglhYoDaZnXW3VEJpgP6t
Ba+yWnoA1Arz7pIuKpjPu99bAr+cR5wBmuRYQn1pXRmNsVDDiYXqLj88uPiB
uTRnWaLtMT9QE1LwioU5K1kGhUdBayGO0dYX6ideE/ITCHLbSOSbd8ENil8L
m+kyH+hQI+a7CR8I8H9UFXEq3O9bNZgbJqnheORiTg5Gc+UWOBatR/8rsshO
xSRYNrBb26X/eBLjm4ANHWIlZmti0D/cSkagyqcRQfUcZDqB5WuVId3tT7nh
T2FoFZKH53EtTIwhC7/m6rf0Orgpw/mdJeXIXfZtKIWFSOz5Dg5pZJDukZX6
FNOCoAd5stu4xe+2TlYuhDJNOxcSUgrUXo3rvxXf9N7LhQzedCzRL8Epu6R4
0EvIFJdH7ipEsoavBjnkpQzSubekqLdrBqjkW/JbFNsoW2rIbzX7n5vcfnl4
vtCcv1ZdXy/i/zkE+kCZHLO1OrLW8S+1XY61jYlsKLnO9+vUiZs3I5nCst1k
Wp6Ow1m9fmlnI3HmsG9LaahJMHr5oIswltMHzG1FAurAf6ojNimPvjbhrnIR
5waAWavNHaLpxfbK5ywE8ZuZogPsokJkgKDCtzxmCQI0Ocw7gF6saftfyc+E
n07BEiWkR6w4/m63THR7CS6vpOJnq/NvMsV89lywjPjhESN2iHKwyaxbR//U
+IL9bF1OX0uOamTjeZKAI1Jcp5lxkFeaOTqeo5p3tR+w+g+WlPVE452Y5nmQ
l5jHD+1DhG+xB0/3hsNP2OMl9baerMU9cpvYVQeevxMmzGk83POtAGLM00eC
XONfdzHDVDZyuQk+FUlTP8glxGJLbmSz8LXRKtlMkdv6FMw7X563tX72ligK
mXDn3Ql34M9NhoquYe8Xq4/TJW+wsPTeLzVbF5Bwf4jp9T6MPtknyUQY0Wz8
mP/2yz3dNKw5d/nlztBf4iLVpNreSkLBmpDTkLtm3tjLdcGfdUXM2tT3sdRz
SgtbRF6fVoOmic3rtOgFignPrrdzRF/z5958HSYVAkyVLvdhieB9FB9THrqC
GsU1ySTgSwy3GXCHPCBmEYeQQduNe/5+QDTOEC7xavQRm7m7xzwjCna1vByv
w0I4EriC3zm8AYmda0DpZCd6QRjyFXEbWU4FW02eIg7uDzJI2P+A9zbdHrQB
IXUWNgpi3/VPiHwUy5Tj95yp4V+hzYV8waGDyagHu2aFBhNZo8sUrIZaGrea
MJOPVghSNcThyPVkAp5tGDaZNoFIvs3iOx03keokiEQKzwPM/4xxasR4JQzx
QoaizCtesooE7oXkgfcApfvSO06EavDdbJVR8msZfQMrwmPr27e4FLC9faWf
3PI7IZyugX/07pko/pGwxNIRcBSJ4nAIhWGbQVrSt93NztTtCf17S0sfyw4m
XDmBqMZ/J2BB7Zikd2ag5S93IW+mCYybTriB/acA28/mQl3t28mvcnIP+z/S
kH1RITzKZm/oHQQEi6vJoM/y1ERaC5l7ZrUL7TUGkJJi3KT6kJs2Je4O2bU2
EKzE6UXJvm/lunaHLL9HSV6DcQ22sPQyfYXSBUrdKU26pMs4+qbGw2sagf4y
dsEpOzzJosP1KCvAFgw2V6TsnAcmBHVsNoA/X4wrmPSgWc/RledI8JDZjiQw
KtPM2fez4qQXoPk9J8WSFE4awEfjinCMSDvyrZ152pBNHtlaxuyww+RpSbIa
ZUUcqIjop0O1afyPzhmmD3TE3JC0obTa7JwDz5jWB7nCxXO6Q63P8vQuM05m
gWXSi0tfyGUiKuWHdxOXFiM9iEOOoOy/NQWWVEoAEaF5rnRvfMHbkPSpjHvd
pf7tX3yt1U5fQKU1TLt73rHJKAfGe+g9gIqfGhnLmpVE+ZYB2L9JLM9yO2yB
Sppe4r1MPSQlm5Un3hDNVQD5vFBhm4vRhp3FushjlAt7/ebPKUZ/rW056aLM
fiaSZEqOlQINjagcMOUAqEw+7izWURv0cFaw07vNVRhxm5PxCbE/0jT39fQX
12UhrzewmzzhsAZ+72IG9FoILjhdupcxghyGUxcSlD2W79IsWwFZJ2mvkvlX
suomSqIte/WaHvillIRANZzsV5PzMpCfgVCKrrtEskkooc/kpB8gVQ+pZrGm
fTxYMHbhCppnMvX6ETZLeLw/dN9vD58IWus/+b0tH3e97ZeEEdZC3v38SHfV
iUi052CGGkYBgJzbxudNePBfK92T+Y5iuZNbBPmHZOZ3mvSRxCmtTQbvaWfK
GG5gEgFyTVst1dQlGzyRBRg6FQN/4rIpzTzcgFiwZxJyUL0M/o7iAkClI+oQ
ZO7Rf8/f3Sdw3JHhPN9pRHewEiyW7nkYwejV4MXMtXlXfYEViQx4LVp48Jbg
Y9tLigXdTfUQHEoPzJq3qcL8KiODd+rd5cHskrhx+x/xe0YSHsSNw1bRDbm3
x8lFSiXHT/3wh5i0pV6oVmhAUDaqWHzvyI7ETJT9ofz2RuM/d+Qb2kWmA7Mc
C+sGvxnqMu7cASpSDKh6axHMe6PakEzvlTPJtifXWqCqILvs2gXGTrmZup66
17DsHGl4Y5PUzrD/qezm6hFf1kf4x103TcIVv3Sg1jnQcnztXbvc42mHjoDn
dt92o672wmbW/27Fi0t5EKZg3faOfjOn/kiEN4XrSkg4R0p+AjJ2+pqL68A5
VJtXnPfK1xNyNaYL8npVLvhX016SzkbJbsJStLq3AVkBbVfKcECInuP3NXsZ
ZxF2CXjuMsPtHI15XYoW1Igx3Sl7g8QcD9wWmMx8N4rDOe3zsznx/wWTCz6+
qiALPkDET9nlqg9zsWQomdHhthNHvLzxInwi8kfUWtm5jIC+bRg8O7M7hbi4
ZYumNr2IR66oiHW9AorxdF+BAs2Uct/IUIRplgIiJzhdn1bC2g1CrkhfxMRv
w+7MkPVXgJpmBLra3X0YBCTmyb5Qa7BOCRQSJKkLbnParr7ubaCQ8OZ4nNSI
+8JasqOba7wqOpKDMddWwYF/sH4wwfkOKVxPQCbjrPEM/6yn7pmAroFm6h30
dGP8lMJYctz2oR7hs98QbwIO1J9Bf8yZzPdvraOPZLZ+U76Yrav7cYf+0OEg
Sr7eMc64ng7LsntMrnIR8ieqfr05kGK3+PUCZr6eFOiSnqRvu6frAp0OQJVB
YJwaLj7HemMvpIZiTNaDvpiqz6syz/NrDJZKJb/OpFmE2j6iHI3tfihO+mbZ
aQO3nAWWXkaCCIMXbTcnvLDHsWTzNB/rPH2dfgH7EwUM9JPuBUWYs9ORtnCG
qvsgXiOhkMO7ZvLeM6EvGqvxPgY9Sb2+obWT2BbNGEK+qJ8Ip4DmTTsvpp4r
+CZOJ0QnGjngH6vONWqPE1Yf0uNgaJNs1KzOJfq7MVjEFMEKMlTGZPObL7qX
ofv4FedRNgBbQAZ4R+geONVmHXhMIFBZJ2rzCUN4siOTPBU1buFHTybh6aq5
diGmhbXSACmpZTX1/i8obsFxYOyFFD8x8oIzsNcSxACikl9EOduP4e/tMKSZ
AChw2vC/xhm3JpK0S+ARrWaW1DJsPfgf3md0JvSrw7sZEtnU8OK3gxBF3QCV
cPePKG/62PRbslGoK75SSZrx1Wu8XqAwo0fk23E3NyDXoeKzvT5xk+13AH0+
AosaF6daCFNkivDzmV46V84QzWceQd6InNHnZ/agcKvbqrgUm/3IfJzGM3cA
InvuJqXl038xRwI2+m4lJNebXvdmKNXsMbQzdKsPi60TmO8cSa36IZN2bDCm
UGDMczPh484NI+R1J3PnmJLRel9QGHOj8UUPiH3bULZGifCb9gPzjhgaqPX6
JsHsqxH1CA/IsBM0iL6NbhiXPNrAbkos4IbaF4t9kqdWT86CsVuA4e1lFlxY
+8Psm1mJeFX4UdJbmMoRtE0pqAQ5zNnZA9LsTwIbGMru7onl3GJPHs2KJ+y1
zULllQp6KNvNROovStvU6XEsR4IZxY3r3/jgodpCjbND2UQkMVrv/dQIEBbA
ZEYki/EADPfcdz9+kjKZyokjhMj8FphtDm8/TCq3kW5DqtQqyk9j6IP/LlkP
DGI6iHp5h1S5psnqATij1aAdEfH8+tgstKjg5QajQuCrE95DnwhQZPbw+SHT
MXQkA0M10QFdcvOxN6dfzQHoa2AplXzKtba64HBiAsAECNurdWwdaOjQWFhI
NYXHifN8bsoUSan5ojgGPOgJLGsxY299YUBSyg1dYwE0SWBGJ3uiSIQReO2x
Gcrco9x/j/n4W5/WP0EfydqfZslEoSCKieavcNZO0d1gbHUUr+hger1jBjAu
5AbCR5+T1nzhNzT0VqErfFOy4luclrotvRjvt7jHHTuwfGadOIxPzojZg37K
/yNsXdCjpybQIRCps6NjKpX6jVI0ujzoMcQy1EAh0ZySyeq1QeSxM3mpKAhN
r8QM4RJz46NsrX6d/qBKIHmbNrEVwt7EVb6WnubLjtgEIgEGFjivWhYL+Xu4
HgOuzKmObSmnickqyArupCREuEPljKPXjN3oDvnCRCmRTVG84eJ/Qx2LASS6
rRibRkGYmX+PkfyGnk/fkPbCs86gK425U8KTqhGcNozuBQyvkzi4A0lIkcdY
DlyGwxowlgtPBNC1c7xF3jlgDiDueo7ATXYpDmMPjSHnogWmLtoKJiCiMeu5
6lilZIAUVuuLvPMQJ2bSrOtFX7X8qIV5mhSAlJbIJlvSkqlNeHCTtEOVYHRN
A1sqr9TZya1K/UQnF7RLdadra5OBbNjaaenSKOOgPwWbfeW1JKbxtnS0ZxCL
kbT8L5LEl3uBfmznM9Gitz9Pogon19BH4+ACarYV8hBYQeHGNVWCxi2/j3iu
XLjHZQRAfALzQgkQ1PYNGxbZKo46k7S0R9iOEY63xT1gdUQpKPQPPowJEz2D
zAljPPKQVp42JINkHtrTmKAYhAPjJbgAjqWbOEzaPP+4hIpCTXh2zaw1+7Ej
NkUFqclfy7hWwL2MXdua5cG+Vqd5H0BcN7hjx52PUjV5fbC3IdddFqsCzl7d
jzlSCVDNZUusX3hADD8D65YRC89I9AHVuPlVq044lkGxwlBQM7a8upIg5O3e
Md0ZAsvgCtZOltl1NtsIPJinpru9V55WbsTbugHjqje904xMqk2Kv2LVLun/
IGi40NK3Lc/OA9cAr08UA6AHF9jFVlvforijTx8MVyZdF5YCZr0nvc7WZedu
Gv1Dd7kqjl7F6ob9yVEegNzXHql6IkwCo4CHnuRFV1aOkvBW/aA1HBgu/KoF
+2aGvkFoedINubCLkXj6C9ND6w3pWHHKF/qQh0a6+4vQhi5kjVq+gxgjNQS9
WTmGCybyVA/GkBgs1ITQtm93PCiE/edhz23pWsdAfgovLmoTK7CUY6mHu5/U
filuvZeo8o424AEQ5QwdBnrD9JoNgz/mXNaE5wUAE6GTk961UEK8tLeZ4XN+
kFggt9G2aPrCfOyFtIssAPpyVFYC6V+7JYI0MTERfgjV42piwqiBcfk7Ftv3
ctab/lFHGTQj69M8DxMXwFeutyxF4UExRRcn5tKMeXvr+8nJjRcol1s0ZieZ
Vl9E6WBSM8duOsvKNLZ8h4p4iig0CKKt+88stRbKZrKicPywdZpP91t/8aOl
yvqSD1lTc+Hf9w1yOPejBOyayZGBtk1Je0GBA71OAKrR4x8ny8SeaRs1M5wX
DRmvTACqzxPG3C83vZLvGAySED3a7acW8zbyAL6wr3geFnr0bLY/rUf54MoY
LiMtEs/ilAIkWKbgX2rTUMDs27nk5MjrWeBUuSS28b/4Cmc/iPaHt1KQ6gXb
enOf0zkkURozdHZY8GZrwv6xbI2EHqtB2rc/d9zeJs+jRZHQWadgT3m4beod
vWBPxdagrerNDuiM8jPxAr/IRDiH6v/keTIynZhEFrqkn3p2VfaW+VxQDw9M
kH9k70+rUCAPLnyRglJ9KcPyz3v6ncDEycpeYBXzEN2o+cr9hXA7QQQoo7V/
LlUv5hDaVk9/QYeQMvqIaV0PFmLx2SEoppzcX123JMJ/2r6F/kU5RuDN/YIA
1rrDg5DkvuZeBcwcWYLyShLybG70wvULQjNd7Fnxf7qLpyHqOZlwSCOW2v4C
5zafY6roSCw0lfbXKPWpG55VCXZZhBewmnwZj+APsv59FWLCdOAluxcfvVew
CB/0CTYWcXpPXIlXNcWClgOS67b3N7v3FGMdksXY2Ebw3ipNNWIdMkcAxJC+
JqIO6s0tllt4+FB/6GDmRYtTzVcg9gKxkIR0Wem/gYNML5xri48u0Jw9md6t
yxP/9S6zI4DbFHlKN5QejvHab5B2keiCJ/OOI8x4YL0eBJIAaarp64zp0M6R
e4yBRED8yefZ/2BwJxz/Fc/I6vAuzIHbLMNQYCCXHqT0oHGt0a7bFdk28Di/
3YlzDHgIZpfcqY8R5pS4IzFCgxi00lGjae56E1/RcCNopge8xGCsfhgccDLz
JDwNWbRSpKrWOXhdkUysyNzPGvfnVCXPrNkWG0gJgBQjLBDtlUcrtTd1wgGj
aq8movenSqC/LRvfKgA9Y5H4bFAV+F7dugO2Wxj7PTLuHwn9dQWept8m4uzK
sBn9UB4frBTg8NJu2Z8Eq6s4wftTdqDFIZe4cltOcgTUKCYdgmBiUFMxLId5
5qagSlKZ4qqEdaahYRtY+rklM2U+nO1XaR8MT1HEk94CpvUoN5giUpeiKQbf
4CeqRUzfGcXcCJYqzFzLdGFtZer7dyyNNK32yZ1LgEaj1Z8HqBGBxGAJG1Fb
iQXiLZro4h79sACjAPUq3rhhIH/xp1rw6Tc0UzcHg6FLVExyo6k/H7X9RyM9
S+jlPLDpMx5QBObjOY5m8WaIqogwvrD5B+qFaz9EUbxHZcxjtciTfLc0T0Zi
sMgBt+PuSD+xak9ex5PyMCyEhydu/Dcm7w7hXGzxwb9dIZXM7I/jOIvzqjQX
CMz4ixU/gQCx3uE1M8b2neeYFXuyZtwxCj91eHGExYD5XKvyO2uTdLjZBzZD
glZElPBQMzUCL8y+OON8z1oJtI9xVNVr0U+RUkSHuL2zo8bC3Klgoqnw0wFT
3DR+bsQtgA2OCdbjaykljaRcihEgUWRRZE7MSaegSdwPMLj33AkINaEX15OP
sRBujr2L5BegYvGTh3THao+BrCOC9kR7/DdBPhLunv13L0e6JQbD5pq+/YlY
CnzFBZwUJFI+F5mGW2f3Q+mkcMafaVvjVwV5idcLE/fw/p3FaSzho9uMvqUP
t8xwBHCLafgbF+NUXDnyKR26ne0yX4uA5rHSpMeHi+9pNmZEYby5/BzeDJ2/
3iRktdP8oe6TBVU4y76jOKE8ThLrtTRndPN3RHPNSU56Owme89Knm16QiUvZ
NUYLc3WgNG+1n2s0n7EcU+L/CWY8IFEFnnJrkZEvqNNdRRatuRlvj7snIjRj
pCinmE+nChMvnrqHLuwa414Ej17t+DaikDmmFG/r0QnE5nFutoiz/n77ztoR
fV2RQHFFRwE85ovqH55gXVk8AgR31gRYfBGm0tJ7u7kH7m+0DKl0lOJYyqFM
tZcjQi56bDbsIelWq/DW3sOUJU/L2+f72KMnA9chWFy2RPIuX/jzIOAMvCj7
5WxX9zkaenMsFtG5ypmIJRuRlzF3mHpJJA6wddcfKtLtoE9aXahIY10BZN6k
bpQ4vA9Pzivt1Pggf7lqIe9mTRw/1xzEy6lVFrKDPC4GMJNvAmTU7C32L2lI
d7KQxtbHbEIktp5YvsMMd3lvgYznhL34i1s8dWOjUUlBw7A6EzURABMGA1Jf
DXatgqT3qzujtAqbAIHQJLaoVe2rwvBJYK674EsXt94idRodhf+dQyt7BEwb
6beUdU73YZFunUKaAO79yib+VfHJMll2G7R5AsiiuoWDlQDXApYRDC1LkIk+
OGJx2LEyXBICzXa025mGt2RiGYS2X0AXtFUbgSi70eQqKY5oNLDfo00FVmXM
pJcnfcvbYxl7aMfVEqQsp0U3PLWEiPL3U4DHrCpN+sxkoVoeUExnUvGSg3HX
5smzsn75HJXYrhmazm5CojFmmJTBpDb66qIN72Sho7zKBOb2r7UeeA7wqQtv
nZq09oc5lgXHcMjTb540oHoiNFHudJz6QN6It+IAzYUyyrjlQX3gTw+frUyj
PLH2EyWxE0wisgjMEldSWOBE8rFVlW3EgRHyXQauTQoM/kKXrdLxvTuW3uGd
OFFWxWaFTTYomeC5xi5n+wFlJn0kBa6ELzUERxH+VJL+0M2+E6iyHkYF2p5U
X8kImeGuTgIWWfpa3lTAK/ZI8sMF+F7hejYoAN2DajOAvsCQ/QvLqnZMQKZx
wE6zBu4s2Z3mGZ3c0ytKZ5am6UJ9Pabm7UaNtk7SA1RHXeoQDRwwAkNjUU4K
9nX6f9/Lo2VgTmMRhapXmfqVzy7iEE3Fjq0KhEsyf5rYaUGLKY+ENHFqYTGW
ipH8zxzoaJwF1bpV5HSDbz+8Ec/9LVD5/csE601VMoEC6zImMtcfLXTmt7NZ
a27dhOYef2nr7EUnNq3U3fUulsfXeprDEcLpAXGeRDE6mK/y/D0QTVhGdCqG
ecCE1xGZPgk5DBfVgAWUMA6435zJTZWDqz2lj0C4ZNoi8z8UbJ3MKxEtwF8k
5BwZ91FXRd/muvxOfIkQeJCwYTk8sxxWwO38ry3a1x3bTQcjLotla9L/jgEZ
QacHr/Ch34il40FWOjEsJeFf9IXJRnSPKQUICxB+rF6UHKC/SK8EE8WvUn5t
ge3mYs8iu2M55FHMrY47D3G8yvcbI1oYMi7Sn6WAlv1SCP8wT0qgEzGy9YyP
e3FJJZMFDdpNvkm0nKoY2MZunwnLTQWHaot+WOm+XtYbTLpP6R0zH60xlp+q
0TfTPmkxjbwR2g5PaKs3TK7833Ngzd1abmwis3uJvcGAIzCud/Q/ESRAu1o/
YeicoVZeSCHE00UlhP5b5TGWfbNx6pEO+aFzooStTfE0hMmEWse6gHs6uDk5
Q+kPPutUBYKG+7A44kWbW3skQxjutu5QGcW+elQtC/L10VyTiAZ7a52Zja6D
vH+PSy6qJEIrx4HGYCW3a6AEW4qi6rv9j4mkX+jSFTp9kPOkJHMNHbPGlPLV
YxxUA68VqwfDNyjOiw/vLkcsoSKaahX2k14DZcWIkh/igDGzBlGuZPZwGMsq
wXYFHDSE5UukpBxh4XCF2aib3taQ9u5XUcuvNYhrfxsEYx/TpGAHULkEyhwl
2caG3JkKgKQFR4PpjPYgm0OY/QMhpOUvFnx8kTcWX/9lhxYzvYG0+dJ8Ftlt
zes3lDZ6K/l5Kz4zDChsut0PJ1nOC/6/v5/m3urZKFMaJtqQ1GoUx5tqPJ9r
Q1eK9E+V+0qXYghD4lYZbS0YsWHcfZzYKQd6sDetgVULeHpWwZJeoib/SJ7x
fcu8Bc+eM1ACvWHOscS0w5awQgOUAxvxGSLDyQcQLU1v+AqPEGx/oFJB4cTn
NsbKxun0XEPp7OcRJ0dC8Q6hMhPxDNRr5i/AsIIlekjsxvTG65qbiA5wYJBb
w4AAvy9q3dXIpYvHHQlZmTDNKrENNMvzjJG/s67Vzck0ASWluMPH9r9ca973
4QzXdLPPeYvQHioCBY5Yz/TJ8WLj7+ahwWqh9q202zrvp0GuvsY7NOCgbP91
5UvJGZYkASeExvcQsZGmnQxngE+Tbt8p+uZlBoQatysB1vmMRpQLxxsIlGD4
cbErARCX4S1WTHiUGMK/Qkjye3xJUwpPx1UqlG34vHhG3iqDy5s4mVbCa7Ay
SRetHzOvTTT1fPEamV8c9KDCo2tJxM0uZsR3puA7QOUQIGLeVtTZR/jZTQWO
tpftcdo2L5oLMuPrUSrQFJ8pZlHEQSof9hDJ6+wutEvapeur3B9gPw8pITfB
QLP/RTIv38eCj9zzzWNLg/SaMvGmPcnLvVCdqrgEDRPdgFz5b/bmvRvH2B4A
R/P+GxZWXVD0YG9jfwDm8kClf6jV8Py/q4jooSoWGdy+Lt/fuOfpg3uLHW2v
+1iTSAxf4Vd7yAcKDF1XmMWbjRA6KjJkhcmtmXeKII0gzGKlYLoVs4wXHG8A
U2bZ3dvIp0hq/0IBYlO1RX+DahyDoXI8g1GgTGnHsrXeCbrpXheq5E3KIQzK
i8rvNWYEkpN5SQfDO1qATuOQ4FOZGE19aUZvHN/sJREbb5rQKmaPvHnGCK+0
vHxnDal+8cSLSZIFat3R3t0AeWFB5LFMI+YNtI1GpPjhR2mrZFtbl0YGsCAb
ip/rvEC+3NyzBDM2MMJs80LJWLq01ri6U0NxSk716X+zcKlq3ZWrnlXe6yV3
HQju7ttAKReHdZHnmZrlAT4UsinPIlaiQe/TqdC93H5gP4ld5eKZ0xYf6Tr5
fPqhqrDJWGbtfjcpbIz+BW8pzmx66WofyAyfK3QYYUipMtDzXVMGj3twRkZk
M3BFFtM2XmwuCmlzZMzqHVAZPP9HkdF5q4cNZoTeJoIbkgGIUgJygKz3+/Nt
whocjjU/nfx3vCtSpU/NzwO/q8/i0ugXnTvJMMWRkQKAbbWNlfoBXF7d/dFd
OQdyBe7wt1WU46Pln6L1ScQEVMIi5AYlMbeXhtZbBnVVt7fqExykt44pqHue
d68rIsFL+bMwKvLbBD2hINIZQ0Qz9V6gt6AaHGvbqZwPuWb31mzcalhUOtIP
FuOg5yFTXFh+UwZnbEqRGKA4ez1QBSdsSqx1JCjjO798Ug8ITAUxs3LlKJA6
N43kryhFo5zvM9Jm0bHOyOeIQ7eI2Ok7xTvogX0U13YwOeLkmmRr4dmSLFYp
VT2AGY935SMYo6vMwS0gtCnCv7AQ+hUNH1aKz2dfIKbggOiE9qbeWQ1P5OZq
ELmNuPf3D6rjAZMGmsdJm9y6V+7/m38CgiMIwjUh8HjlBjznlC1FHyqEqRq1
LDBMzFA5NohZDIyNVwmWRasKLxczA/AiJqyHeDiGKrVIftTc5LfztMpCyQja
zW1I4inKbdw3pn9SQOjlL1RdLL0ZDCkcxeaBsDhU9AyG3p5l6rYflD22h84m
uKGp/OVlTTyH00+jo5QcgX70H//v82mMhfRLzp9aMFBRkKbmY1qOtnzNQ5wS
iXpmmS3Qs2qJa8/jrDvNHkSc533fHW3/opUoA4GmT/s3T4i4lN2EEzpJDaQE
/GgGgXAFjX/aVUSiqI0egsVLnyPM7YX72LaRi21n5H2TS9HdaqVRS0qbkQ8c
N5hBI8/t4BRyykMmUxF1bwIl2LLCHXpHekb8APQHV3kccJqW2+cEtZBbPhG6
KrVcAxPLZ312yG2oiN5CnAGvnNipjMnCqUZzpEXjw9MUB4rvCHeZ9k8ytuNI
qPgiD9z6UaSy9P1rL129wjLj4ke8iSK+7vXZts0Hw7MhecX3+NJNnOcXrTvD
lyOmJsed/kHE7MMklPp+sogg4CeYv+VCCiV7+G7eitOBVc7ioFhcSe4flDDA
P2qrO9J1qy5uBiy22nnJ5onL5KWVJCxqWXBwAMywQUALn9LYEm8IwG1gvTJC
EJHqsxeZ5WIfhMR1u26TEBAqyd75eL260GhJUULe18zWFkhycVCATCcsqe43
dDDinpaIrkctYqxYWFkLxPjveLk0ivkqSNh+k3GeDYdSpKUQagIgpaWEsjN4
ock53sJjhpXVOu34csymLrPVueUYfBFYqFm6Aj/TMP2TYBJddlvhkC5ZXSLN
PLfksnrvavmU30FBZ+i72cwGSynFaOrIFJnsGwGG3xOGGS0WyA4YHt9CaU4E
gzdFupobjz63EwLl0Cwn5PAZ5kVV0+rg9efE05qG2JRDI9IqGOlkytFT1DGR
bGjSiluPDidMuXcj2hkvdhpQg1Iy9zU3D7EGXfWWbbcFPTKrzoOIC0tHxfR4
pG3V0lY2JE20L6OfGupsUvZ+rFlcvijPKe1lg1ESV+NNQQHcfPFRr0PshXQP
VaSjp05L9tzAi/2YdvM9/Cq1SPGlNQT/l8kXY/lSfM0COMdNTtMOpw6/KJwa
nnqAhreAdnjzA2ISGDtq9CviWT/l+AdOKnlodyyYkVMNxcgIlH1LcVtrmCLi
zOdyiLT7HdIPAgPDL95aBXk6ywD8sFzMRcb26/iRXlxdKP4tkO+QKCp31731
BdRa2ChOr3/twoXGJKwjA81dvgvllvFL0nLSX580g/2FrP1c5XHJL41Nfu9m
sWd6AZ6jPdja0B3YH9IzmBJ4QxBXtDbqNhrmlLOiL5RHfB+jasDcjSCbBEme
Kj8K1/hYlpx4bY1tPolU+Yqv3mmuQZisWgA/CEaVv+wdG0ydKWUsU7Pbvmg1
AMV5o3GC3XSGqKmYVMt2YW6iukAJCThl5bcG7cUl0kRrcoMvbvG2yHVEggED
7p4Du0wE+zS0rbH9KWfIJ0fAs1+cO6C1lSKybH1BwJU9VlOz7mKgSlUw+jAz
i5sU54f53xcqWRtkJ0ygEgi6xvDhEun+LXBvBoq2L1bbUwY9OaSawb3f+NsZ
LtOTmmxTOnu0IQJ4aU+VzaIte71fjeXs8C8e7OF2Qxp1noLRjHSEIg0WFHO5
EFCBp7lE/gWFKod/w52YTk/PAs9Iecyq3w3fUD2ZSQ5x/C1qdmgSk8SGDhcO
rhvF82H0DyCLiiniMmwE2Nz/xTLd85sxm534pUnAepYPjqD5wF/nuMbo03Lz
aXrOkv2nDkvfX0ybWd4IxtBW2CNisZekgcEeVCJZP03TJe7jorSKF491BT9f
/DYeUEXSYyxVOfLFbMFswRPcsBzpafTvtEAkpN/uHnJ5dwcnHk3zbDb38EFX
0pfdzaxU8PuNBpyPdGesBjKKSUvxNc1j1vGl54hRfjEn1413vfna15BTSFij
h94QVm1XPotU9HrW/62nUlgxksnY52t+2Or2cXNM0FJgDFjkcyOrWh2AecLd
e3ryt6UGis8tko1X77yZggUAFUio8xlMNqk1XRdHzJAdim5zQD6jwrg+1+D+
agO4rJIMrR2ON9rwCBRN7JWpqyhi7PdZRSk6PgjnCGH/vx8vm6pOZ8Val7Sg
Ba+7F+8VcqkAmp0TwV/j9lPxWfY29246pMmtSwW2ZCpUBBrpg7lml6eNwynK
FlQcbxaPeH9q+CKYzMBS4rxhTC9vHweEpgVGFQYl88z+Nv+YXt7eFk7K62LC
UkkUOl3lNI/EzzeLbKEeStgb+V9GRWevzTmNe3FkAeeJ3mK3LyWSi3BFE3+D
Mod+iaYFKkTFUy0GUzcljmZ9bBxHVbxBV+XxuIaLPJWWEHuhCNsBOCQ2emp1
HsX80dvXvoaRVhuuxB/PmfQN7dejXBkjhc4d8UTIMK+rC4wQ8Zz6cLd784Ce
w/GoR3HnlRdpT729ja/geK+AWqhcjc8B7ARdS3rCpHsrzQnQnOgExRRNqYwi
uhefCXhrRReTu6MvtfrwCS2uROojkJOy6zl9EyMhbYEvqVodqzFNROrMadan
G56L/FGzcdM7Bg3UYzUae/yuxBz/PKaN7wfT544+OmiQDo9scR+7ujPrZE4/
82lmzPYMqn1iuJQjQ7wXz9ox2ec7we6Tf7KuzxErAkElanjdB9bwnpb7NtTA
xH3jnO0iC0InEoVbf2KwdEHKuc1T+vZWRHbksg6JZpqxbrOrxRz1vlsGarGo
6xwJzCFfj0upCTN9/tiJ5v8hCCLmiKixS5fcwwJgTKEy6A1knv16sNmAkRPI
0nzaTsYlLShJ8GqF/PbgoZs7wXq5ad2lJHs89ROqdGq96lyA1dru0dEHC5wC
uEZofkIpvGCtdJfpWSZYoppKYVQ9eQqwjXcxVRS1zS2s5yG7M1wQMxT3w+Cy
GiWQGvzXxMzAgRxoZ1T9thn0ZHTuUaxbnhQDMWvRRJ9OcEBR3r0weGZGpSA/
Y2+TyURFgJqhYxft7q2/vAXe1LaoKb76Cw7gCkXlV60cOikaTlrmziK+swys
tCo5WOBvDJXvyyJzLK4whNWNzyXa7joXwSAP5yD7pKFa/I+lT1rjKHaaSJDZ
Sgn103snMa0J+cxWNFzpEkCjO9oUaW8YiJn93hhxyCFXDtCxC2p1HpThDC7n
whlkSVQkB3O5Lg8JFGAbER9+CO0T5YqlowDrGvnrg8Ogm+DUOnq60fn3XyAD
XDHoqy4q8vjdM0JFbkadb8wzj7cm4oN6p0R6DOnAZWbd9xNY242KA+2ei/h8
aRWRgcz4tgIBv0+p3VhuiTfGFI8eCL/lcTv1eGKK3lttiQeuobu4QRCUPN0r
dnNgVf1ylAUU7RKqjsqs/LOWj4iFkihqA7DxTzMAS0K6O5TrrEoQjSQWYCS1
WO5d/NBbWkLBS/ewvWzRBJgbQWS8k6cORV5aK/fo9RjtB4Jaj5ITtPO/0jCV
w7qc/0ANpHxOYsJF4VaiUfTIiD4wGpdCwDsssqGPDcUunuR/nPpmR5g+qzIR
nPZlV6zHzUVGlXpJ5mlPxlmvpQWZC0ca8cTRxKaFSIK+t5x7Yvyci5nirjFw
xLwReK+6iKBnptr4MR7NTCVmMW2UcF/vAjPHMJp9NPVPAi0klZi/J6Y6YCeY
x+Bzkx522mWsvySWz2dNtzTjglu9S89USgm6WXs6jCVvp8IQ3zAB7aOnGfX7
/ABxwzrz5SyvSDXZjrXlByoEki7xCsA2azIJMjX1jzjh7drQB/py+vdOBm/k
kU71N0o4iQIigl5J7h+AEim2WTt+u8+KMzR/MEWAPA9Sc+9yL2cx35y+SKbA
hQcrbi/SjWVjBiOFosR698VLJfW6C4b8scn9PFuwt/rwhHZSTMnNlx17HL0k
+COokQ5NAv3vt6zktqwnk7TeaHOkSvhwYZtpSIBhuw21Sie1rNzJ3FrtZlXj
+LeGVfdVa7lxMLBpypaAJmkBW6SpXbM7Ak0faXWnV13J9kbmV8/anEDRAlfU
kIah2YA/xSziR/BwTjT09ZH5Cjvyg5clRQELpgRYDTd4lwvpIvRNn4xCB81e
uYQFMzYmsZMZOiZyrm1S7egtnYQxz0tij6x7BPdyEi/reFu5CnGL/3YJBdOe
b8+b5PN1rx1ff3LZ3Yf1W2WRhTq9aI77IjelXg6upzLHSEzJa+GUgMPyxEUo
gqyYWjY5EbxL3Liw35rndk190M9jsBVT+4zZrTbIToEHJpJ8f9O68PQihJZA
nqnXnY0rIePu6znxi7LCfx4muo/AFuNRXz9lAaBwXzodS0HTOqaq1H7wJA1q
Oaq06ikEpDqFbCh/x3/OD6DRAHWxJKJSV2TTVahopB+iCHzC4qSU4Sgz7hIZ
H+vUx86YokU4mRulstASxrpXpY5T7LNHLFkJEIPTtFMwFS7WOQk1TbYfA2RK
pXMFeUxiXSuszJ6DRtdDPC+fZaemQFgyxckoz9dMDLJ4XOWGKKS6QnFEe/dp
dtnHLCrWo7QSyfEyWOyssLXzjTd7RpUx+RJ0kPdUI1e+lyvszSeT6Y+1F5Qw
EzYa7LPxFR5xEuob2WxbcCbGg6h5dMqQG3UanKGTpyWKx7Iy15YkXzBVVOPK
tImAvfsfoKlQg3wVe+fWTjZXMBNQGxoLEH3CTbZwVU4q40UTTLXMt40BMzOy
1350BHgyxcrNtNFnnmZKCUat6rDuOC9PdbbwTgAuN/EP0f2IE4+UqBe3h+wN
591UZfUgQ8ap5QUynSQqCeaZWVZJTJ05UzM0oRX5+BzLD1mUvL6js2mdNIMv
9hjT1HkF29ta882sOtbp758nm8BBC1Az/n3R4fL+q3DLTgNuoKYGIo9ed2xJ
6vb8azcfHcX8m/o6nJgt6jPbcgpHpG26W/ZW4mCWKMS239ucPQ31Rtk9X3My
q5Hn2RCq4Xn0wkkDEHEqzh/h2aqD5mI23RyPbJkLPZ9PkeHQWwT1p0ay8aeq
8qkWEZpIEPeuz+a3iMsQUFYVaJqNT0ri2nRPWPrPGrMX0B0djyAsr6BcpmWc
U3XbIL1Yum35umA/0mRsITyRg70IbqcWUFssEJt7Ih6rQthzCNN0/dND0sB+
KbWvu6Rc9nFdHAb2Ym8mKkxgvhHlDQwyBaVr6vWNRq4ZatlzlZg8gizNF28j
E+xKffLOo89N0CJ2TjCsmZnf3uPZVGzC1Fn1/E4syYWB3RLTjqZAYzHBfP+Y
qutY+oZOra7zrx6EN3i+U2DVjN8fUw7VresAropPu/lhSn2ECzb/xq5xPlR9
8jH6YSeXyWXAPht2KdUb9uqPfMtha80quwjjusr3k5Jg+/7sYKiPFtQczUAI
QWHIavBasEL0f68AzSRYXKbD59rkKys3//FeAJO8BmvgI52dEQ+Fajloo8ug
ra4LMC3vgzvyE3/xZ8/XXF9cr8x89alJo6A//QSM3MSZkQEZUaJyetoDtXWq
OvMGiZ3CksDqAxVC4MT5uC3A6Eb/Pvge0KjF5tvYtVyFt9scQ9SDEzdGaEzw
/cUSMAw+EicH/Q5LSaiD7/xGPvnyjGNR6DASGqci1Ai7atR2JwFd4tHg5WuA
g0xiy6N3gm3x3ohO3M2T+1oJxg/+dsVWh24rmABjXt5cAxQUCvb0TYm+WP1R
T9hun0hHAZm2QcvMqF9X4M0Dz+0+oSToA+qxtnrxkmvfb8c9luMikA7hAPtz
OiXcpCg1xhsqMn23IIfFH/gYo9LFzpfoZV8LJGnD0svnkue1BejlYr6o2wKr
QyDG74ptRWEfrr0hxdDllYL2f6sOM9M64f3NFfnd0h6hFlsOEzhKOcHFBMSL
XtkmS1XP7Vu9wLTrh+dEo32HsPJyPxqwb5NqXleAkA9NOj4ehcLOBZTYY50L
eAz+Kk6aNPvgAI8neScypg/ad7FbvB4eP+DSM5mwuPuV/2PC58JQB0uFSUYW
y0YwQEs7zieVLfsoycrCIWFqrO9hszfFRPtKd54lwF4bytG+UXhdBWfwaa59
fmigwwdRH4BwGZNeS0Dy25Mo51FhrQty7yVXW8tOEoNNOTeKFuFwWHYxZfn4
OIfZh1Ifz86Fy18cVIIkCE50W1J/4iq9EjUJppVqrKaNgSuzSD1As/bwon2U
q49rur0SWtQ4SFHvREwakD9zfufG3TltaZmGHU7csHlu5tO6mIdu91KJHSkX
KwAHCxXP7PwEl8grbazvFEVliFoaTU6TMcB+xlKJh4TrZZphZfBNJzV/HN6M
uYYur26vGowrCDASdK8Masfxhhoopl5eslWS3Ck8ulO+MEFBRKkQRFr4IgMw
R5QjBDIwHnmJ74H8HN7ioIAoaOyN9++XhxplU0x7u4GV5AErBVd/9aVqfh0S
BVr3UqFocwVfiawngfASjuEVI1+ZXR8TFKAfesMqpJMjsyO3So5bdZGhGtMh
KGU3ttZUZWwy/XZ1tkO6UmW22rQiZR/XcsqTQmGbJybK3SIAmqVeQ3zaYdHY
S4LfXK/wkxeqUKzSvLYiuP/IOrrRREPqhp4ctnoVYX7tzmr5sEka23jnTg1o
qbrpBoIUPVKmJBRLtVbylgBQVanRYz1SFKOiK/wylYQsg5UqD4o0mjwa98+c
4331BrBCxnNPDueUoo+c2a2dV6rSMfWhBXO6XaTqPBJ0B/zeIF1+jKTRLySE
uP6P14GVcOm8HyXV0eBz2llOx3JEu4jlhQzlYrZwaBiGtDY5eIxnQqTaCEhq
KtJ4H75PhinoYztZIaJ2iwueKK7h0Z6rWjL/IgzrbEgqcoE7hl1zSO2GrMkq
taB34H6J1cKJQ2jijZfsrUjwNM43dHLwtX3M8eQYOJjQin9BhDpBAAiOBWZX
6J2QB33R5kGEhTsMnMmbUjfLHye2alH7X7ajVqFVvtObgYtIzZRVZ0mkBKsH
kfmh58bUhWJi4AHEtANjPOT04ZiVTZoruKN9i4VWxrZXqStjprUbRA8YWEIe
RsEvLOHHf7uxhki5GMFi7cDbR805pdBtXFeAKu1yI10gRv1jfGhHf6JvaAKL
SLh+GlBqSqrrF3E2LFlJBYlK4rrfMSO/rXMex/KwtVaH369dacsmuUVL7V8m
dONBseMyfkjr9q2Z5vgvYAIo4WGWzlPSzew/oGhqwBah75t9PnjKG07DrGmj
6vD3LDxjCgqROph7FDAqC0RjHspBvtwBmcZrv94GQ8sGmyJh2UZP/iek7g2A
6Cp+7FBT/LCvopwRHItlBymSfDbUBs0PiYHoFf4aM44MJCAk9hPjm/NaFt0p
XB1Xz0YiujLdO6sZQKWkf9weOaOvYM0H3JdNl4mNH61/ng6GJ1TXlLWDCh1A
jKQ+bwwOBYjXnBWXttQ0VN3BNW0ZojFiJ9P6eZfsqObymeqK3t9pQuODbT9f
9eNY4Y+ikHcBzHLJ5u8KzkrTr/QgycQSXPyVnDIfQc4li1AICr2U0v3+6XNh
U2O+7k7Z0CCtjzlH0Ss3UpwKNjU3eY1M4OWmcGWDTvfV60HOgFFcCrVFCat7
+qOjT2JvKitz2QlHET7453BTV5DvXZ26Kbi2+PNo3ZnIxFhQ4eLUO0veKGEy
7y5aAVAOQDqWiV6aNVn38eHQ8tZ2ZYaG9YP5vyQui01aiNmSxJGDQn84zgOk
HCvwFm0ih8G9MF0EZgsKVGpqT1DW9oyo759sCILMERmHOn6xlykAgav3lHFN
GyGATx/La8dklkWx9aLEairtgjzmPZvhBJ5N3Aq2LKppVMDEktUiT0pn4rex
PgPz48gQspqdoU8lSxKBRjZlKNFz94/NoIyQg72TMv8E+0lSlljqT7BHN5Mn
jcVlZIANhagfBewevzwQn9JPeFg0EbYJSVw6C31l3WCWHw+U/bwdlsEq6X0k
tj9U1Ldth9dM9idOaeWXJu7GIrstNGveeL2h+FpaGRSHFXeGTkLPbbSDz3lH
Sk1xgskwL2iBimZCV8a9/ascGpIqz/AT1wdm/oVZK97SIJd24QjOiRQGZA5V
ZZ3IevlX7jLB44skjwOEMUIlkrdglVfzkptXyhHLKNweIR/fTo1osepUu2BY
0sVuejP0IipVDXk84kTo4AXwiuxAirhojIg7rm4VZWLCd305MqhmfU1CFYcr
bfNjE+bHR+aM+kd/mLg/HDKVvnAZ3OmR7WPAIC8mlpgLJtiON3h997bREMKc
HWtNar4/sCUF7hbrHupdxsnj5YUiu/UNYiTeHA+5HvGMDVUrQ+/OBcKteXGQ
3GczQe6jOViNW+U068HjV2ULzt7fHgHyOJi/ZG4BbbOP79h5U+ZPa+ECqfQn
1skC6JJFguot6Yo62duh8RkvEvOKo0Fvq93nECcLwn7PBxsFR25F8jPbV/Av
HM0kOcCuakmhRSyX0ntcgd/5/G3b5BWh8vsnsXzmkAXBC60xWPvKH54QWpyA
F5rVoktQ1BCAWP7a2w6j2vxvd1dWFykKFXYj8mNslHN2c33BnHBi4DKxxnC5
a2NwPG6x5NjQLEz2Be/kC9AdAt6VcSiCza+6QJ3MWp2SOYhKsvyj/rviIDAu
A+RacbW/53q0RkcGBgrO0xVz3lbDa1byNYLje0CiXu0lxb1prLQxRGhuk5Vn
s04T+zhXVgch9JL9opsWoe+xIv77v2xJ962NFkt7FKE7Tlzr3KVrDz0wZSBq
uWqWWNPZ/mcJvwX3w62Wg55pdR+wrR8MRWgP5ak3dtO1s2gI3N5zxJnRJC9O
AcsLckex7tUkQ3BD3C0/F5iiQuZ7PV5LHCjTG25lxirz5QzOs3/+cUBBwq3N
whWUdiFsIXD2DHPUrO03KzhWhkJTqPnEeA3TaBKZnvobs+IcOOUYWLaALwmH
UkktH7ufVocJoOxirWMQ8PZV1K6fd19Gkol5UQOUeOHKYvwGKxcBZ7jZ5wyk
/SMi60YUieEH2RgETwduEivoReWYqYEV82E/796bKZuc960Sm9/+wZbtVO5b
q1zfJ8dLcW2fGDS60UuyRASJ17OzaGK3VQ2dVcGKU5yICjYc42QdQsg4YFL9
pxLdNEpOgfp3wieDori146MKaxn6YYRt8+zzocZ0nk5s8+TQzy3EV8wabsnM
tFPkBv+B7UDpBJqIIxJbrfEGNqVRxMENUvrlyOWuj2EiLpUD1sSgu++LsNCb
P6Me/tlRD7iVn88o+AduPzJiUTt5OQrW+g4A2E2y+Q/bFQ9yyIQBaCadqXiW
kC4nyfnUbxd6QxBcoFmGEFw+517MhiJxKcd3McHTrVl7sCTkHc2o3MPE/fEb
3fU4v+BgTv39GSxYYvGsZ8DU3Tq0SkcSrNhMwV+oNOKVNlaIvcXXmlzitQ4f
ZAm6DmE/37AButzqLVDFR9eYIOT8ukqN92SlSqoJEFtpPJr3uxIRpuSkG3NL
M4JjIbXCDK/sHvA7Eb/LWpYx+K0JMX5KT8NfktKpCX4/vf4pBkWiMaKHYEps
wIPtTd97fDQdawEHfUJCrjn1pdHMo/VwnOTwmT94E054BFjpj7eJE8rg4VQc
PfuMACMPMgC95Vr7fO5caquzQOm20i+piszCoKpPDsy4PT5YW814yLxMLynW
8l94/TykHIdWpd3sqqqFwazQvDqq4CYQD0JLmfk7Jhgk6a6JtaqB9UAF/hpM
hhvGttjY5l1H82y8ThdMBk6nSTjd8+YiKyBM3hBIIbPADgKkiH14Z45W1+AH
eNNcbHC7gsokN8GOcPsHR9rIHj0zXJIiAG3AK2CNvX4EDRz02fc4jqS3wKEk
Yql4hmFFjSB67fOS6jfHBYp7sCYAjHgmjsMxIKhRpqwW1FRNYAKH/Ye1qOXJ
G5VkNEyaps9lXykXv++2tJyT0rR3a9LfFxwL3vNpE4kFsys6awRxwmTcjH74
ZyrWf9ggYrP/5/tz+gqTbEJofdtnasoWNAMwXrAyYzgZn7MRUBcPakmsEh7a
n1/MdMZEDnc6qszFIgqrAcWvnFHOnM2SmKwCRb50sd4E4vaeER8sN9/9aWOv
eiG00/qeW7Pusb99O6ITZQDZr5wadfkg43ZFKw1Bsaa5YJ416RUVzqlvb5Hy
9s9h5F5d5Xcl6AMb2UbU0UfxzRnoX1D+RWOFMqbOxpJGcp5I0f7S0sNIaRFb
JNHGEwH5fNftiFD5ZM1DTo6/QfgvQPBH/uQ4EX5f5DcM1TI4Voxn9xKtB2+w
lgQTNCuky3g3kCQctG0PoOv0TuKmh7rhfGrY101vfhexnB4cP1sOQ4bFl1vy
kCHmML/Gikwyi8sBNyedvaN5VabVFpMWdxQljxrSHpOAaVZMB221rSW34gdN
wfedLcO7UU7grVnzMqcCm+Cu4bq3/UXkIkgH3otZmY9qz6o5Mw1jM1NiNwK0
9GCKuN7Dp+Rul/GG5iVz1V+UUyOyxXxhqbfBgBMas5X27KEJ2QB1aJgzk7SH
31oXwBCAv+JXD5BtTN4EvdzeeE9umLvfD81hiOsfkXuuoPmHQ4X6v+v+STkX
kPhfK8bGpqFCTzvtT9HOWzCzl7Y0Xo4LTA6NOdI3D8KlqiHonvRop4qBaKOf
kDgjJIcEk7a7LSJ91u2VVBDC1dx8wgLuLsD0icPqvXW/8BWyVfBsunoN7T6j
CzHqNtqhgPhb/FRAXHilKotLSpWAAMCzVFnl4Thz3hcG8shjm/5SIdbXV/tR
5dGn3J0JQxTrFq7OPXOfdlewhHUur5APZQdz6iMAfFKnx5jyfx31ynjQq6wj
5HNjt2KSSjzx0RaJZu7JduqNFlwVk2oH0iJg9imDrXy4sL9pjlKn5nOJCGhl
wNBOfhAcBsG7vu6nLdEgU4CwNxWpGqVZkXfxz3k2WUqVBFrIrupX4pU4PYPB
hfuIGPDHW7IUL6YHRnj4AKslIvKOa25Q4VjsnYm3shWgJUEJCOLgPHO9IpL4
93Hb7eGW2feCK+WCx6W3BGryRKGZ/CZidNjLsYRTpeSQFdOn+xiQm66NRLho
ALmmT0Co/9bhLc3vUPmR3gkfz2LJdwF/7j9rlWUWMFXhL8tDphMIx5eVRoM3
dPIGr/8AuXSBM0p9V/5LjBpESX4Fy2R0g5awg0wcDpJyYVKs332ke4WXsM+X
TIPjj6VP8ZxZPNCu6xVYYSrbc/fom7ATdgYxUi2veYzsU16FjjkzxnTY1Z08
WpzogYIduX+B9wJI//yXO9VkkEn1vkJBhjfdUEo1RllAMYaSnIGnidQ5ZZMg
sVi8GlIhxAek1HQlXpWmMBmSCFEEWkOdFKejvVrGBngg9skMseJGY0wHq4aH
3+S3Wu2DrIccvJjjD0i9gLw/WIiDoKJVWqNTINg5ZZlxtAlxu4SXTZDK7KKP
zOj4vaBYAZmVpKIfemm8ECYPhtnhurvx4KiDO8YGlLjktTSHCpWIerAX63qN
PO9RPMIdrKkiqbtZb7RVQ4Ow2ndktLkpJNq9uXHJxiII/DTbBd4UolMmk9LC
tYVqpWr5PXNXOAcjKUnZ8+/14UigWpREtGUJORvkoIPVoCIJbIXVPtopZlm2
62YeAb6z/moLhBDt4UA8sFo95Hhndc7E+hk6NjaczYGV3xfXUhk0tuNRqrm7
H6QNBTWRo/m/s9w6WCzwY0sZMwxIkelIOAsUqcu6lTj64wsNFkEHmdJmR1gi
glhRIbEgUe00ygGBBqDibkzwF7VWTmDJtDBnv8jjBlevZYKtPfWPeNmK/Q2i
N6zQgCYyay03qFfO29cwfSeJ1V5u7x94Fwb1kMeL0E7J12YDZUDfxa9Nrh8y
85xvKsYI6dxkTI2VOywM0i/cEcy6c7gA8zrRjAsqFGU/lZRY+SG4efgExhGj
/bDcInB8tRIzyd2RQ8JDC9hbCUwOqL4kU1dbJYByl8dcCwdzXC6nMMLbCeuV
uaA17c+095fOpGkPaUXCmVNaaOV1WOEC/FsNqSfXk5ahFwcyEM9BjW/rMt3u
BVYzy8ArAgmCscGgkQ+YDUDqCpqK+27QqfpRXvbuIWbDnqv/3nuBNBFMSX0l
9ll9qydwxZdfKNKq0pd+5nHak/a8fgXCMdUcre1XdLBPaRlFgEMz+2eQhHZN
IEoElOAunCDle52W18XJezdvnP7dB7vteWQn/ATbC8hefMxcaF+R2NXoPkU4
OEwF9UnP85f9IFHQAz+SUtb9ZmnKYUI6HNfDWJw3bYT8U4yANMPAST2aNxNh
5PvJK4GEz8bPmyz1JO97GRAY6Kj3MKnWf67bbz59r7GlH6Jo/4Ff1j5V2C1N
0AGjU972MEH4/Ojb8K9DeX+5iDho/+oAi+abB1l0DFP3dmAm8/jHWyXswxKC
E4U9WIriAMV+3f0BYQD1X3SiXZqA0n+N+0OkxkC6SqKgYsvzZ0TUPg73bTaO
06+eu7SHqI0er9ifK5j2ecn5Rs4Nk9qNhsSS4vq6sxXMlQxAwFZNBB+Sogus
ZTI+1DRNIl0MU9bjD/51Agid7iIsG2Jz3rcyTZfepJXpcKAfYQTx1+cQmKG3
0FZH7Iupigk1iAzIrgT6rwyaDYlSmEHsBAEFcN8JD8ZFH/kQ6e7WMcPn38EZ
l9BqsERrboI+dMmJdKxDn86rWUzVP8qhKJ7mclJ7HaQtwJFn+r95Y88E0LZl
tGDjRq4Mq2u/01A+PO4UL4FL8CnrMdomw1C/V3Kq06/CldCg0y0yT+VzIIiI
Qjkg5/jw/mZIOkVVRj8w1wcyO/pdidTqQ1ccRIon8z9Bs3RI/Sf5bK3ezdIt
E5zJ28ozuwAeSjdcqISTy1RIEKdLKFFiOFxrqSnm7j7xdLMN5ITOaD3YJYp3
O7pqDDKYk8CNK3fAoVtPIKrOah97wQpWW+PjHcHwys0FjFnSIctzEbf2fF4a
haIxYAhVTZQb5HoVWSBvTi6M4PIa4TftL+hgIUfnCbnk9J38EDtqrphBXW4Y
xt4V849rrpFznRs61hAsfEmxD29neiwzLK2hFtgDw/D11HjfImNw7aMt+VxK
fR/G5CtCke/A7ztt9aj3zd8xgEUSUrIS3LHSI4oRKPIN0RGBEKRCCV7PW/pE
RDAPv1TDx+2/l06MLKC3j8g42cGzU37CePdDip58efUTi78uGDleE/YF3c+n
IMPsd852FfgiwkILgwcX0dkPSRiDJFcHYfLqyUhmRIeSEblAjlXZzy9PyADl
SXA2nfoq2vbQ0zidObN1hgMakoxX0IalkxWEBocSz8WLKQv9rjczO4cr65Hf
8GBVJJ0lYRbaNRxwaRuGcxhlXjBftXjIe5JorXnzq4GblzHmQedAdzcdicMh
FyJjwe3LVjNZtIxFIVG3+JpqlUNdm2pBGSkS6rBidDES/iEu631BD6l5EYyV
HcMX1aKomSb5TC53Ggdj6Ip+cjvP9tZi+02pTq24FmiONRN93445mAWCPTeL
ewv/Nuje7u8Hz088RjuvhPX3daNsg6GqezgzmHDj9plNsVBTJoqlD//jrYKT
3FV2xFrTrSTlZjivsnzPCYKMYYr6kIGw9N7UQY6Qp1tCkKUjbVvkBBSIelpr
nOIBrv3WBoySkyLJ+ok8mcojsqXcxA6o8qVJ4PRstti0xDk/Sd6sDm6VHc/D
G513o4cR0Tzn+5Fa6B3rLKSvAMWVE2l5wYBNNFrniXvO9EhZeCI2JtN1/jOA
IWikikGcmEXmxuPFctNDgXoiWdRvCvQUDh0YEzvW378blJ9MnDiLr0Lo9QhV
trXquc0tPvtd3Ndm+vKfndtunukz1A47WNS1CRZ8QmYArKnmwpN4Qq4lssS4
KFwW7d2MaXzl7OXRCKYUBdrj2Og4csKgJHLWlrJGlR+xL8wd9MrtNOO63gZj
WctyxB8LFMmGSHZRdP7YP+RoYeROH6TkaRT/WcEUMkYs281Qb2b6SuyxdNsp
AwBAGm6ZEmZIoWca9xssUYbDGrWdLkv76mv9JpWGJ0W9AqvwC05PqZPEhB2z
zwCSvC08Kr7IKXSpOLidS2fqRccuvtno/71I6rq44w5xdigFCT0v6t3OKdHf
KwP+FDG61ijDmh1PRqiwZUs47j87yDyK2OZyPRdcXIvFelwR5hoid/R4Vve+
ghauuNOtKzCWHs09zO4zxuSfiUQr/wSpUwb4IsFgyaKjfRizNvYxNepX7eZx
G6BTGEaOvF0/IPp9wx2wFT1bIV7plPIyBWlwPi8n8ENwLh4GxbmgvONMI7j8
dbnHIlQg4axtm1spcCBd4CljdeCEFy7u/j1R1+d+jHs8cTHFWjR4YDbZbM/I
ZyCVmjx+dtg/nFElF8LQKH9sAfNOp6lEhb6YNFekj2oWSHEMprB9esANGwbQ
CJ13eamk5LHXatH/uwKU/5ep8tIdaX6WM1YvNuygr3Y6acEVfGYOqn6tsblZ
6f9mwHFp6FrAjOhW//bhF9av9Hi7Poz9b28+3de1MYmInoJU6phXCKpQlVMx
eP+i7OVjvtytixZIq8RuCXVh1wz6bFia+b/4h1u2I6Zt+yk6cthFV2BChEgq
5VEoySFoVehc1dQbX6DUM1uyDE/fdTYtrWeuBUFlklOmaeLIiQvuA+sRcQeK
xnX9AWnPUFj09d1Fsg21HkxII9FFDVcYHcz0fwyOxFuHe92kStBjO1CnosPf
4p7utVozYYuZBhFwRSqBhhYcZnzOkcnZgVLbAr8tFkeKwrXv4rQ6Mk6y9POp
bWy5e5QiI0ncgsR/V1F1czn+2kTmeknQzhxZbcTl8uL2bOivZjd4aPnoZ+iz
empa714u5RLp+B/2kLHB/1RvWwVIqVvcVr3ea4Czz0sLWGESoId0l33rDR70
hfRjCYANFmSKH7BxdB9HReZQqwvXicQaQHupYz2xgkv3nxSvLEe0V8OGks8k
G7iNn61d8XHxD4tzfPVVwEQ0de4Ivdvm+eeUGbIDUEY+11SbIX3/dtfFLgNb
NIhyYeuDpk48EHOOe87I2OXOi1w3MwgnzzT0N98XFNRqaaJeEUP/Zdg3wHEE
6wsad2v+GL1JotpqegLPsEi2MUhHw5TuWGWXORWkwipXxqI0beg6+zEG5Ogz
Kk6EBtvicms0HZFXpZLMJG/OWnh4qQngLZj3UPxoj8Aq5Dg7eOsa7P9UhzMG
iv90XI8SIKK5Pu/udrAf0YymkFFDTfDklWD1mG1spm2ZsWccyT2K+aT28RVi
5tsd3gsX5hpWsUSuNsrrUux2wjSyr0AbqWxCyBMiVEOiIVn8ZTBQw39d6/2N
1sCn9cYtTlDLTHFH9PPxTaKPCTvYXByt8hXrMx0SPkwjyQe7x2E4v5INjwqL
Ke0N12j7+Pm3xYEBE6KSv6Hz1v6qgfJsY8guSfRnzV5KCkti+c/Yo9Gq1mbL
1Ui7pciObZPKyPcal7QcIAX4JB0gd4eDnXo4eHvRiqa7VE27fTHOiNsWBC4n
z+CQYiXFkDCZPSyKkVj9nze/lRShZRccf2hnrXRZDYMCOP18AQXRsyDyNF4g
yz1FuLLCPoagutKHSQQVMUwEiBdSWOsK5oXbPl3qoQxz2Fjtp+85QbRGBgQL
MFUS0za3DA9aCBtlVX+H6iIgP1w5LQ4FCz/eBqt87exCT6j7O67o11+AnExS
kr7FV27uAu1SILzTGtl82zx1iKkSUVtKhXPaTRIBpZZaJ5jdBRnoW9ijCBf4
HeNGeagjGH2wyoKi0n+w/a8VyRLTpvnR+CWChMgy9HihfMlTFoEHFqUbi7Ca
yIpNnbAE8JkMHO4+pDuhgJZ7OAYBvhGlzXP45ulNipD6Gp0/QQcWR394oK0i
ZyLHyefrIezjYABqy1CqHTGdNnbB88ybBjaG4XIySIyQt7ZV0b9/3QKKfJXd
WHPDiWdbVQBqNSOTKSxnjI1QlVkD0i00BFKodCIMz6cq9esAzlcdmIEYJ5K+
aFjTX78PSzlusnWz6ZbrPU8r9a+Ifqwrit4Ks6Z2g1gdFZ8os3oyr+dq2WqC
EQBKicRN+7aTwv6ybjHGluWqt6uXlZng1KnhQ+V77bDl7+5Vxx/yEkXQBmY4
JGk/adXL7dlFF4jndAbe2wc06IasYoGkUdXxpVOIPmLOtVr28dPsGuVdc09a
daz1BECmYG850pD/rFQhS8j/a6cSPWs3CInxrnnhYSLfVVVs48Uvy3dEXFtd
ikQEDO8SaPsM5bVHZ4dhlPaUbYXZDZ3i/9lmE9lQb5inaTQPo4t7fZitFSQ+
kSV68ihKb4zG89MPXtW5sEpyZdLYA1vaREaBaq2sahTKDDmATs0gJHUU9ULe
+KNFwouR6LeOjelrIq4x5Gdt3bQ5VYMJGqmWC+FZVnTmUnxDLeSN2jKzd67B
/3HdB+xIeFrpdeUs96/vv7DqQhV9/ywcw13w3ZwzgPxV+uP/st3BLkZ55PgH
wHxzn3EuheywkBI5XJQyGIrl2mgBiURse7pEU/xEtqs6jwUPKgHPLZQRYR8M
J2+xbeOYAlKZe9LH3xqXEHDukijvQzeRfnP3NeTICm2i+RODu5kteQUf8sgu
tRVC1jySuvSR1keIslLyH3dIDOCmAFy79PObF45+Ft6XA65n97tpN2G2U2uP
99wUb5W0qqYbdjR8oEZASCMlHY+2/bgGLUcaagjAULJMHgg4xCptaHnl0s65
XtozwiYpQUyuVMm0zvIIDJcGJGuHpY2GrkhjCy+3kNSa44zhyNuLXlwi1A2p
BDY0KbH9RmAV8F1ENU7IX7v3VrkzhHTtXxFjknm3JTTCrJvh8HC3KX5P64QC
Twwarn6Er5Z3McNDOr6rta614A5BmGoqHnr0SUx9z6TDKF9+mbohlK5hNtZh
REVDyGewSdUl8XljaexScadFq0NxwDhnd0IMVbFMGkyIWVJPsVRE1HZL7Q2w
ouHfZ8bUVWdSl36df260ZHyga4Ge38WrzNe3pVWcq2E7qrqVB3emYoGr6+Cx
YN8ub4SM/kO9ggIuT/Z9z4PlPmsdiDMDSPNInYoF6mWmN8bfcuZ0OxUFgYuQ
rHLR5rBNIuJ8mKOC0TAV9Y8GqCcmN6RO8TVU9Ug1CUaYT6PjQe1YlYmHqYcO
ocSZE88YRmgQD9o5I4Qjv7BoY/l+0L/WwNKjcyE6ySHxeyTVGS9mg0Xgokur
o09BNM8YMEmCQxjeD0zKcEskIenPTDm9rIGeJXNyMbkEpDYa48R2M8E5Tu3M
qLuAxdqd0lA1qtzJyoCk9MYQzX2WXRzSuhGj5VEWDH9qCU5nMpR8IqN3DpwZ
Gzbe6hScPUrnDspn6VYRD7WSQ5Oj92dJMuBt4lqBbrh27He2PwR14jVob4HQ
RdEpH3dQ+ysqx2UbfUmV8GnzmAC/hNInp7O7io1Vxved//Y1jKs69R1mMoMY
UERIaB+kUBE99PMpKVLbUSd+Q+XGhWIIjzizWPNQMu59aAngvFE3oJyUyaer
+UTnbOP3OZecWe9cCuZsVLz8bRNjQQWO/RMSePubT42HKl9i1LRLeiixWH8q
KZ1jsrIVqY7aqOvqfJkzuO5x7WBuR1Tuisnl+wurQmf1EBoZqWalI6r90hkp
+z9llLx9Gwy9plE1q6mN0pGBMYyXedS/FfZZCz/YV5wFrXv+oiN+WmA6NG3+
aUt61J0TyXFANzOnJ+Rw2DmsaGiUjmed4x0eRicYo5ZsabiCeNzhTQUw/u2E
8H+L57lpLabdgbvHi1FVu2sI1WYZa9af/r1DDDghwL+FrbdaN0tVLP4sYTp0
zBbXHV3ZgCQD/WqYd2i75SiNu7RJAxhir6vchsU2VrSAeFjAunYC7FVRBAOj
coZcjd6iPWSKMWN5tQmJkVnZRXWbhjD+9sQE/S1tW0An1SlyZz8iEUYWHwft
n8QmdKe6SxpumZYlwjzc4ofaLpT6M/CqIKu+G9jK6rMqAm1T5C32mut06AzU
wnfRW4n36kBDbLOje2hvDZHwSRDXpwWfKtqoq56+mU9H3xsc7GsP4a9mAIAl
WAoQKUWpCgBs1uNZmGYJWTA67o9jqwY4jYcDWAHLtfpw5rHeB2BL/gdDr1XV
9D0Lb0nHDm/5bKFOSQpbWa6Yh0s2n7+7cUL6koKYEY8kAcZlYLODnJ2Iblvt
B6VzA0F6yCOPlYz3O+X+/D8AW/gXSZhtC1lsV//74n5uhdJHkHil0zJs9TFX
4ut7BG6aZKUs3vDSI80wxGaZS2TvZgxOdBI+GpZs41P0L9IVSL1Q7IFRxUri
xGQINzz7ihyITWaVoXJ9OxScd49W1NnVUG0gg6gAnW8qPEHS5oWmi9aktJTh
+H5pHpDpfQtqnrpOzVlwmER+eGhjqpzv0CmJH704Ht6MLw4myytNUPPkHuL9
W5qRjofQp+j1zIXwVMJIiEEtGu/vDilcS3q9kvB3OS1YBLVVSuh/Yh7WPosc
Zjuk9rN5gV782aOkkxKPqFmrP13nNg8gV1MaMRq5F6KIgMyqqnSOCOh0Ob/y
A7ucMdpqmt8OOE6S6yHa1B1fRXjPY7ZZRlmxM6HMSKy+xEuxCOPJAwO5179N
VhE81xNjPf/j36q6GP6b2AeRzGnajcdVAP+h2vHi3ZYbK5vrWGZ5nUrPj8g+
Vwgxi0u20OZ/nmTZBolHjBWyfL5fRvXlv4Zno+aKmYIo2iT4m3Q0Knj0dVfB
lCjr3DKnlcqc59RVEHft7OdCw7lwBB/ABoY4uUTRmAXYKefW7GVou+HBmARU
0n/K8HZrrvNFBS3ySREYZ7T7Sig4W91KDiqSQZG7HmxHg7ypqL6oNRfXhCnE
4qm/PWMKZzbDnsLZTvkztB0h8DEpc75ijoeaCOEmhjAJRBQknv9ELNADZMhR
ws11swSR0giZ2ae0kzF4w+HjyfBcA8oDtsBZArWJjClldpuxmljToqNRNnlA
EmbA3wPS2HO3Aa/sVwZeuRzsg0NRjEKsp16GcYVmzyOY4Fhrs/uSiX42WXYB
HjwejKfCd97xJdxvZkh1+49/ABVG8SuMTHSEUeOXsUc9w9ZcuMRNXcHw2p52
h6oIWg2n8KUH6Cl6xCS86ojehfCerhWNzVn1yYcaljGXkDI0Ki+BxQogvF0S
wNYdV+ihf5ZOEWVNRc4PW++ltMIlAYcyI0FI+Ik9LfLjzTpZPFjldtaPq2kA
PUPnjWSoeLVJZyVvowdFEkuo5Y+MxU54v4dY0BEWzfeSckK38qm08f1TEe75
IFWqaFFFgvMnxF2Bl4tZ4+/Y/THV2v+aK0gEob1Zgh4YoMP9zKK9lmNhW2zV
7tKpVWWge52+CQO3ne+fVYDvPHJ+8Ngdyd4h8JS9oYKN6+XGhNARaWEr8icE
axFxoLHKC3nCwHHmpOdPwiCz3+U9/RD27Ah4WKlezvQCbhE/oic5/+pCA9mM
bu0GMmtSyxi+BZBzKpQV7LndRvHXWHyKTYYdPcQupI1ND+KR5oYtoD4UVsd4
sJoU16HpWUvT+CU11/DSCPbXApWxAkSeUNt+vDO0uyDODTLF7AQkg8SZpygJ
fQjKg/Joq9Iy62WFJiru6mQFQnfMory/tWujuwB29k+2XaCW1AyX6zPFsVQz
0dOvBXDvSXbH0ARyJDYWV8m42+H8d+9puNuYFCBLZO2u/DIzm4wH4kMnWzdr
cksBChrQ3FuT37Wl+ygv9fmmy7u+Zntq8+I+x8OhyCp5RAk70GEHhckeQcD0
2KJXO5iHnSO55ZlbF/lfy3z1HCgcYaa7Up8PUWqocxrBuSb7QdODbPrD8SY/
lIwjZE7/Osmk/+rWee1t/kViZPo8sLF/kcLLA3D3oUlvSsh9/6qYA0n4mRR3
m7l5KbP+kLZMTStZ4YunuztywcP5V9Z1rqblhchFES9BcZkbNK8yjHc2LNhW
7iDt5F89VDiVAfAg154bLuH8pGBQYNKx/A1wuGK7IO6U0qCUyCA4S3mMUwBN
BfQVPbTIt6HEQRcIbuKmULKXmAZpJjgDmumeviOjAhxsy/69MXgIEaf36+8N
gSWe/pnDy3yUYenClwXvFCt2sGXvwqquJPzXHn29akb2wZtDFfzcHGZgI1JY
ZlbT6offsiQmNEgvt69rC2FW9rHSG2SYUVDgYgVG8qPdFYYYtYdtjLl47x5b
V+XsAyyvSADFZ+bN+9gq+cKu17REpgz1q9fzQGPV9UZiOAfrO2T5xHWlqMFo
pIkMXGKokbt+HV1LPM12rwvX2lyGgSAyukjlE0sk3j6zQs0FrzGkXDkIAoY+
vsxeYIsI7Ue4qiUbCEAzRsbM+nRqfH0quXGN1n21yu+PU0eILrPGHjqYSrsW
1YvxGvr/lQFAkDZlI0roqViTNo5HebhbvLKEevpaZrLRbcdRCPn+u58IT6L2
4KUlBpkL/xYyg/w0snGCpsIsCEazNrAnUNvhaIL/L9icOiP1F/oO/dqZXkDO
akVoL1rfHw0A1S+Gf7eOYIsgJuSGD2fq1XZpcT7RFqpUWCcAAJIcHOJIAw9F
j1+RiYoLjrs3YZ3JiwG3hFwBqCUijVWEW1VBMLJdiS2o6RBoFMg02h1ZUrg3
ViwdE8MwNucErbVaoB/nBlvauoDNenBehmP2Bys0ho8NigzcqAiQjsHWGP+c
rhv2nQW/hABGach7KlOR/iGeoj15VfyJTUUUTYDAW8pxxl7Nf0eOA7P2Q6DZ
/73FJ3FflyXzsjMeUOPUjL8AQq6vOH7HHk9JbkKoIdOnQuf+C2CGH12vcQyf
+/VpgvNQRYirw8txxWH6e/aCMP2NoEb5yFU6RtxcxAPJVZ+yeHDl9cDJsGTh
bY42nH8Uvg6DZH3Qe/KAHClhpe43c0NS/T4MdY0Hb4wMHhPI43OtmJ48nbue
mee1TM/fxQm2YcjwMynpzQhokzBt/WpVKm6riIz61K29gShvPDmVFmeRD8hm
q8xjT9B8BGR4WeOketKWbb/0P9bjjWJE3AJc3mxTkjXJNy3tJzyAIMLzecP4
rGWsIqdKY+O5Jk6D89o/U5dvcj/8uY/8qYUeu2kZEsQBMecilXKaYgxa6v+z
aT+0uirIjrgWmAJxIdz9iBsDpebzMQKPExdWoV0aYtr28haeysQbkrsYqOn9
U7l9QrxaIOluv7CfSr3EQBrYtf/rIjrVX98DUHoRXrt+gwzdQ1Krs4eDPcL/
QFcg9oQiJxY6APsJ9XcIf79cY41x3WbMAYgiZRTWfpUTvjcg2pbzCoBd8Ko5
57AZ8YGo6rW6gh8GrJ2e68YCHRhqAZaeoYPNONOI6gmOXRZfTIx3G1D4sI2B
JtTSdnOxMv8GS0VrzreyTSH11Lz4iJ83JzvEmaKAaBR+vg51ooCPwjUozk7u
w+O6xCS+3ttGt1zfyMIhazxKuaZ3SmgltefQENkJvkJzd8jA15KhodWAW9tj
SZtFOlhQj7Qu2KhltZeZn/iQ+JeGsc632qhJ8IMklT5Yy4q7TA7AT/XKFw16
FxQp5wmVg2/R+yf+JgIS/6+Nk0z0MtqVCs7HZE5ywQfPxCnQ+bH4AGc+OPl9
GhVqAJyj5Jo7hgawyheXE4O88fXrzLxF9GR5afy6akq/HzPvUFjcU4p6vAY4
/ZUAyjZXSSkuxb1aUrB+k3kP47JgtPgVBsWcYS5dr/ZcVWa/8c2g68LdFMMC
8i5+SUU3piJBLxU7lyBd1RioCSH6WVWW8JPrOmiXWnaTmliRaedH10BKIf41
6xgZ4uQjgywzBbBTowxbp6g2yZd3c47WuaWpEPG6ICKfNOJoqlLlAuo0C7jw
PV+ccbudNgaMCnTuGtMqtZaR15wOdCYF8L6DCH5zUv5X2Qyh2vP0wmyYdv8r
8uPIzu5Cb+BmXwKlT0E5EYrFoaAeVTsJ3tht4Q6273D6tabnVIq0wUwM37Lb
qxKQ5f9CXXkZt0We3zycS1xUKTpvW/7BYdaGMHGvlhXbFyTVlQcjW1ey+Bjz
YSgpMWxyeb+V1BNsMS+piygz135DM8DDU2z5wWG86UoYuOUMW6iVvIEmDvfM
T/oh9D44pJoHgG7Qr8Ac3CQMRNrE+aISw0ThBAfhamvr3qKRPm9pQ0VzkvGq
58SVJQdQNYF8qDSwvy8U5QsqXwsaqkKv9SkGPjyb4WosxTDmlsTsx1M4b3YK
uIan4FULR9HHxLevioB8yvE2/LSRTgp0nf3wmPeseiYIao/Q+SwXF0+/lU38
lOpxLXzhEjdunxvwATw/yGiDJxG9bZd6u6sMQA/i21yZF4K9NxefyPUZepFE
Q412u1nTUo6ULEiTLN0DpOQjy84yzdPpS/v1nWdztw0dbRHGiZpgbHk31heG
qe8esC0r9/c87pwiaHYyVYeRapd3S+qJjc155g4pMyfmGD7zvvIh/q7wLAXC
qpxKdeJLbj2EqFEvgfIUaeRau32JCP8fw4hhpSKs5afJbwJ3HNSmhpPf6Pda
73Ja+c/ek/waQqy3mTVaHGsDAcERaMWrhZNw8xIdg7X+BFfzANfwDnIwaXHW
iUhgP7eBGz+J2m3ssEC3pJTjxjMIpibuc7ymDdTJxeiXrSrPmMwL6zbyQKr0
safp8Y9GY3VrkoLoN8dc8xbnb5WZrtNx3ztW6oRVZqRkFWE7fZOjo20+ZcnF
StnpiAZiWroagceejziYyvYeK8uTB4nSMgjxqrHPLPEcWtr+t6lbsCitCqKm
flIDt+gbdJpAqD4gBixb7SowDGTN55XjG3+zz3q8gg0Y1/QbNQeTYb2FKVpQ
zzSlho0aFEs2iPN+/0VBR5fr2K5oilNqDFoixlUPq0ycmjs0brqZSMwvEpPX
0eYkmoxZByLpAEUQ8ZI0gT4PEzua0YfhI9BW6zYpSqiNG2zjxb/ywDc2lde3
QaTzYFyFOKwPXGLGJo4faaXHe9M57r006KPggvKnqx3LtzOsXrtOMQmITtdo
NP7vCta4+XjJgpWWwkEezPCpAwgnTZ/3D9PrYwlqCvaQAztBnryJneAkGSV0
ds8P00ykj0xAbZHUL06ILj4iOZsbKwLsCDOdAH/bd66VRRqL+ZrNsbyd/O80
FtZ8KnENXzbdsExXAcEByqTP7miU+wBYMudzd1LnGh5CHcSnnQVyTOsIST/S
8QoY3vogsuzXwVY4AKKuIjTCLARJDHRJ03en6na3iYGzHWQmrS7fOXz4mqcC
hKgWNMccdiB3VVLBilXIL89KBWJQITh4iER7jlLpPMKLdQvhe1FPs260f4Qj
2b9ZEqxv/D3tmMfGPdfmQXdGcNuw1ZfDeJ0aIlp3AKPuBJ7amjwPmwZFypCf
Dd5JIygMxz3Jm99lWSwJExcodHH2DuluzJJjvlytivG3R6o1VGDlzr4tihNX
JlwsRSiyG5AZIWYHtKTyNlSWqWVgpC/ij87ninCO1sLpMe1G90h2uo7WMcog
5Bw7ExP6tME9eadqwgbvJgoiA+/M8F22sdcQI9ADcacptZTjLDBKhKgelApT
ushE0VWOMYpz6BYgqoo4VSU8rBih43ERama1uaRNtSQCwBFHTZLsBAX1yaIi
lt/Bct+++uQk70x8ORlyFTuobyGgoNt4Vp80hz4Iq07wGYa41gBdbZ3yWMbi
+4yHXEHScQo0bx9iGZcxEpM+QlJyy8LbarT4kJzmuK2IsSdFhbJWF3BliwGu
R83cawU1IqscUOe0kpAv8sIcDRAXfOcXJsRsnkiYziH8Upe4KlSuo3JR5V2Z
YINTR/ytP92yYoplDIZJpDE+6ReH71YXjuPQDA+anp53QsbYA5OMOmrHIUlH
VbumFX+Dl+JDV1WWKrg2sMJtZK5bcGLs1z1sprgUDkbberlvGxvy52ZmJpUC
iOg4xdXC2Mmpa/uE8yDIcEq43tkdaiiIJ8I+YJaHujDQPggpE7+G9U+jMPUW
ZRd2cx9oUumu3FrWEuk3VdXxTPKWqsnmbpBB9CiS9c82xjf22Oj/WyVpykFN
CN/K6grzCwv0o7Z2MeqQMIK3ny1/DfUsUwWUshKrObjrMRfGg+NVHfbrrHnO
s2yVhwO5Erd4UznPEDc54lKswJzddx1yjnUOsM10uDhRfM60YvKrlA50ZGwK
9ybWpxvMiMYQ3Ccqz2vBahnIlvtfrUnQfZZqOUp11R+HiIGBL2voodtP2SdW
YDpY1IeC1ZJK7iXufwNHu6yZzJV6uALw64NNIsgUppVSXhy+mTxfDy6k5bhE
K1YSFmfPob0ck9jZfIwhPjSElXL6SAaTbR/ADp6KAjAeF1oaEfEiizHJkbtZ
E58bWPRlmqK+yP1lHXTdagEO/EnC1XUnq7v8hc9irViuMwYx61DNr2yUCewQ
3yVzbdotwZiYtj5tU+ZPSS7J3qhxziPsPVfi07VA2BkVNNwL6URaJlmq4s8x
jGHJvEb1/lafalH4A8Q5mPyvwoYSOrcNtacE27M8HaFUWAosdtFs4oGbt2M6
NJATu6GLc/1+lsrSHJo5g/GSLrGm4MrO6ti7svpUT5zJvAwgMgFAmEcqlPOC
Qbe4gLhnjh9dhN0mAgH5FQGC9FLH9Cte81j5em9mxVo/OPDV5GXSt/NtbNzt
1V5BlRy2kh/FvQsgSgDzkJef2VDu0EyBVV2mCoE9diZYyWPo9GpWsnjInEeC
ts/aZeqkINk2n2D3n2ERgUJdqNZ2KYaezW4VeYm5qNfPQGGjLsAhDhF3qrD2
WSBWgGRh9d1RNoIZIKXvG9HTMd2A2Si/odiw1L4aHxCLhPtSdRn7mFU4J4MQ
NNhCfD5NOvidutQltVdwokhPZWTEleKmHU3Ylxpd92z5GpgYem6HO3zSEpST
37/9uUgi7WJ5U1GV0JXJN586EogsVaiIGlN4vkQVrBprHMrt3QBRdr6ITrR7
Rjgn8lPl5zgVYOgqmWlHulWZUf84NHfu2fl81Yhq3oKNSjFpZNtJUmfkoTJx
aLONWIu98c1sYdKJssH9pxt0b0cUTXz3ADicX0O4b1UHAwcNrFL34wJ4MRA7
/UM+NzD4ayJbnF+O22QEoYvUI2yHd9euEx31iXdjeiRTY60Ern973KvFkRXC
wV8DC2FldhaKx2IteFEm+zA/e71ln/sopTpdOku75eMZBO1p+d2d3s3RCKwQ
F34GNoaRUV2jY8/EHR388fIELpYse3tGzHKt4mpDtcrBslDiOCHhNj0QEm5e
Ox295YU3rhta+28ZkJPay4VYqOtiEPYyto4vAZVhVJPRIKwUJSXt0Z66GE1m
sOuGgrhhExX+LKTTvDnfZOdp/XcQzuz6QRqxrGBSigf/xB4fgY7OpLA7kl/x
ilZiZP5/8wzjtn4jzJCRCVz/2V8eiqnDl/L3rv82wcbJ5evac5qMuoB3p4z0
4EdW9YfcOIwWlfBCGRES/jjuQIHvu+9TLTeVSxAhM81VOiYukCFHDcA+A10X
9GkWFXraGLVbPLuITG6jNm8zyigtiFaIdRGYns8JF3fnR0/WM7AoNmPYD/oB
MEop/rNzy+TPVCcXmLJmxelpxVG6OY9aJjqshFdw9/z9oZtw4TIv2mcdl1dH
wEckogMute3y1L5H9lf8TMdSJFdoz/C84eIxgvyEHATsG9YXgbYRUHiPEF0X
g0CqBM09M7PBZs00hLx7+zTVsETvOxH5iE+QQBq+DQuSNsWOLE9dzJx1ID98
/yXKn42ec1FsGHwZSJNuslIRYggqcpV79Lrb9834HjVRxUCzZ7JNck1F2HXv
79TaEnobRwfSoL5N9Wqy3LQzgi2/G6Hcs4yf2RmXfo1wFIHORfwZxAtuRs2m
ertk8/Zwp+7YKThZJ7vsWrN5Kv+/iEz/IWoq3KdYJdwww1y1btbr0TfATZ7q
TJ06Qycy2jA5aDXA9NK3eHM06mlhSlNpd35UkEscGXsKcZFz1K5dbAyKXDb0
op8ouiT+CEUi4FC18g6SWUJSrXW42GCIA+EUnRzbH2xUgwy/vaLuMtuCw5Za
QwPEc1dhuvdeBUT3uRiJUhrpT940+pC/yVuu9U/LP9Zuo7ZSK0o2MvP2c6Zd
Fn8dNQzZyyHeidnxRyBu7ZtDoqfr/4Ip4nH6KqJw+wAk+2K6DWKeXWqHf5CK
3P346HO4Mb6OR0pT8zl4YE8463ENKHsW8Ag5zYN6W5UvdZFN0HIa4CkDOV69
coTLaRBtSHWkwC8Z6zWXpqC5zB1G3W37XrtzZK9SAc2vkFg5a8pyDPmCCB7O
KnEMEVRySj3a+yQur53dRwcsTfJNxTkMTkA2VDWtZnVQbIhf+ZT14i/IlSRW
35uTw98PBcVJOIn89AAHHaZn9lVu3eEPC+8K63rKt5O9o7VBuBdY3BznPSEe
RWLGIjN+hJ8R6Sbvzy6mvi6mjuR/PeaqjaQR99sXX5/Mxa8pDEzlmMZNYM9T
/wVBBh/W2Gbc4YdT8Q0wh/OmOv7Ik6k+uW3EcVFEREuq21BFhk0zpTyZOYsH
6k0mRi+Op3A0H4nv6zobBTYvW4W7c2LpmR0GTzBHA9tv0Q054Gh0tWow85RI
Uy65q3xwtfg34FpBQhKbbFe3oHnBxrfosmpJW0ET/F6xuwdnPeHQimc8J6tk
DCsR4HOwyOxnA/ntffMXIDsFzrzq0fzxp09ciXTR52tyO3LOqEV8luzP1pNX
LWGj7dTTTjPegDVad5yUBMHjLLmUVTDHTPi+Yo71F5bInbHq1HWZpF5NiepH
jwy55mf9Wm7mjJZB5brC30Lx+UxFqNiIaQK+ZBes7gTxkUzOQsm46ZRH9OPD
cChYCaNcp8lQcGVf3mhGKkK/5onFX55ZQzvPbAe+EEBSohVY6JcFXoGx6m3K
7gZxC8sWePwCbusTn9ha/mSZc2qzVauna2HIHBkX95ICwPCh2nTMKmZhZ5OX
kuNMFXpL8FWGOVEy18DbxJMJM4GhBBaHF7WPFOqvVHXsMl5vrDQ8uGkgtXej
MCsudCcKrKGVxnN4kUJD7oNnZBrDk7QIsYbdipt3G5/H+sfDssqvA597ozj8
hylgJIXFFSjktRUZ/n1sUnMFeppCj3qPL37zBryxNvvSBg5KItcZZrdq275v
+4JoBbaDIUVPdmT+7FpZJcbebvltgQLO42kTXCe0PLgpvRv1QL0MBydv/7SY
LwigAMKIDa7eREzhxmPmxNMT4ZKdt49l68onGNyDIf4uiAB4OuMEolQqvNxF
24OMcAayK8I7q5XWnEZRkgoyUwsMUE7JgPbs+CND+di9JLKxmBxSwBpiY09l
20rTpJdmN6Eu9Tt0GVKqp4y1lAgaTL6azRaVrcEOKQgWFPaYTLKb1r1ow+pP
OwLy5Aa/6wT7WFx9mYzrugZjiZ4z/TDhq2dl2ueAhwMzF4LzcBsn0URIdsIE
6Hu4fyszNCGj9Yu6VMgHt9QDc6rEgC3n1K6No6ndncloeFk6CZZicTwIPo8s
WVGNsejMsnTW6IjVNJ3Hf7OzvFguIx+mtXNNvPd38KBYDSam77p1PhzR1rOt
NkTHMkRkqsu8rflTj2xxiDBVWuTJ8tuxl0rBy5wxZIWbU3McDyPHC4fDlyZn
P8fik60gEAMkch9GCY/taxJCqRVulkKVkNEgLf/xoYcd8axTDeZiJHaWYsRi
Lb8EeR/i7ZeklAqBDmM8uYdeFSAhyMHD7AGF3X7gygEUSkweqfD/O0jwTK7I
SMyHR/+3oOHmUKPhmZEwiJvP10MnOCU9BTVQ9w4vSX3vF9h5SMlS32qPLfv/
YdSwS/4bl/RcKuZRH9DxupHk8tJyJFqnHpWO19sStX4q4sfxEOItt0Pk61dT
LwVAugoOb12/ZU29XHyDYMlbpOwpofYMtoWs0E51wP8ujbLxctRgFVN1Yc1j
EiCp3Mf4LW6s19YHwlg50uLfB+BlOhloby1VOAoVtWJBnwUK4bkUsFeufyWG
Q/Ha3CDVvd0AxSxImFhKjvuE9CsgD0xunSGCE6BOVhh4aalQ3VTOTEVc1t/s
v/kytI+H5+oYA4Eeoo+GvbJHOhqbtYe6dgi0LXF6Lud4bLYXiSOY8Hk45b9W
NMEqCW2Dz5aULGRnwNXf+pbs6+VTL6heurlIWBtJcVRwGtTt9Z691K+DNpx+
jj2XSbgiiF4+l/f3MRQamywBdxPUnYPWMwV2CPiN7Th7b1t3rdOSj+I2L3o3
IWCf6nddsO3X20YcOQGBy2aGWhMlq9p90Shi9Bx2SvUKYq6FkkC2tbDgHS9d
vIL1qPGqAdHWVkpu+kz1vcglcrH7DNDZnlXmlFbPChGI0uQttgNyBFg2hQFY
Uo2IF5svyC2iD+r5tlClnvksshAB8jJThZRX3N8v1dDWVmXQC2G0sI0S5PL6
z8MSWBHBTur2jOO2TrMn+RVf+rEGwXW1IXMmoR+/AIBsgWDtZ+oXAuWUY0tz
arw0HXxRi7y1HDdbt6vDJGU/YUxT676zfdhqpKOAzXTtecrp7BGYwKq2wOxQ
9UNtXMrBzcTwVHBKD15AbOxwu092fuSR6bn9nnwACKlj00BBqM1BiJidU/UU
sT0oKsPU5hK2t9RvNaXda6KC1Q78auWFNC22uzdyo6sn7gfU41bvFrz64+WF
nQOuCGeCANZBAVoQqomNSspF1jDyXztVeqBexDyeZPGBOXgDCGHcEt98eekT
+XkLf0XPOCGNTVnyWtUnNziXEu2GS9q1tKn2byO38M91QPkXNHMU4rqQgMQ6
tsLclTI4evqt5wMcv07/kprjtN140ivgDELeFNeazJEc8DMpjXyUeBa75Cv9
qfLDfEamo0EBsD1wjAFcUMmMsfn6iW/DCcXg5bVY/Aiy78C9llrPpw+nqjCi
F8NEtTwfcEis4FUTAJS8lwUOT21wJXAeWpNdHLn2/ASDjmENcNPX8gbH47Jx
GynF+wsSyVQjcpbSXkzLWUjgMzDAtYwkZuXJ0UeuiGVxuw+cqoqd3V7oQSjv
AstkI9vVtMLDV59mCEq2BKnbUuSua5gXeUkkMejIm9mP9/SK7wKDXfbCthKE
CrOCDHy7EyLpKmZn1BM2S/EVeqgIeEMqocAP83o/jhK6lNcLgnCpOs8w2tLQ
QvA6o93Brrc5CPB/jIyPf0zRSoUnfLZ5qIFfYxjtft9hgO53JW5wCHdP+Zrm
2vE/fXGgyOgGscDDsAQGm4MngFKcHvAGiPKc+3Zh0OxGxGM58UEQ0HymBs6q
IxfjAv5Oce1ZuWR5x7XvJ9ujABCW7xXZgsq/ly0N4xeQsEw9MsK0NowtFddG
kHJw//Dt1Qqw79jGvvliK5rpP5cU/Jgk3WChTxuGoEsygqI5YqI8R0sVRO6w
+0S4U692GUTOCz2exTbtTKwmsk2XhEQwluEtxpWNnz3zztruaSLksQ2czw2h
jESCiyZ6kFNGc6NeO2PW2rpgDPbhoOJimjJVDqmJt/ojQsyVML9JLz1ThTj4
zWyBBpRD/UkjxtzjB984KfAsHnzCD90z6vYtOtNrmyMgn/MsdjoTl9C1FMYO
Yfhli443c67PGsaOrCsvtRknjtevOMowaHHoSq4/PyWCAHorvNbroxDEutg+
gAwPjnOAXuj51SFWMoye7w6tr5O/2OGePMZBS36fN2Q++Ar/1pxJptvzrq4m
MS9sdfnPYNvTw1+GpABHrnvORZwIOlkavicjDvAqFJmv4cMXH+mW3cvZWTXp
8Qe3mrOsreYLZEJYzZufELTSXDEd5KeUrzsl1GSsFqgvzva6GfI9WDSNjDiL
eAEVsn+IQ6xJG765ctoyNbvY1bembcXupwiPpw9FyC4fIAzAkl1Rg2QvBozF
g6C9OLzM1aVDyyAdgwN6ugVqD9+ARS4zuX0LgZGTBVuUz25jJMrmWdi/9kTT
ZXptqmO+pbnlvnYAZoy6mPWETeGyM4huO3RaygGpuGUA8rFl1f2Kxtiwsmgi
ESNCCuUEWCk1P6tNlX2bb3cZh5RGkiOwIMZyddL9riRphZWn0fWxb2YdRbX7
R2FkWbUO/w3G+Bz/wv5TnhNe37P6xnST8QlN29e3BRaubabfJC9hcomD5JW1
NYS+4kqx2yGZIdMV7LiPOvTGVfIWtSGBlmUj/mEg/LjQJLPUIx8wMUxjmHWK
prhSg3W5ZTICT2lGbnQZ2frtyOpS9i2rHOxPOqsGnXkfu0sX/9pvo3LP/6Ag
PV7EPuMpqBzjbFt0zN6HVxrFPTgnxp51CDrL11wiMv43J40gRyoSTKQ9poXP
RfLjZ/Fxh0Kpv2JHNNA8voIuAkhNoYoOpC19a9wkgmVF/k9BsewfL0dW0evX
ZkspHNlPGvVctkNiYLFEVIueFDc7DvgFXXLIjGffZdxyzlDAeH9gLFttjEHk
ELSU8E1/WdlT9l+XxN+mUmDWFWZiO8jqx6u5dkWxZ0np/6aj3PNNMv+5C9Fu
Rwt92KYgMryiq+KLcEPnKMG0jglhB2Sit1I759wpNIzKZULihzBuNS/UpGEk
xlvpdkZ2P4rWC+qkbpN9wpNyatu8yIFuPgmtYafX021Z0rAR9U3MBbKDxXGA
vjFzPShz9kCgWIl7GCElOkTqtgryFpGGPZwd2n4yghpUTjSiAJAboenxPMhO
Zgv1r98gbZXgxCZSGzNAMLtEyz/DS5jtdVft0VejU69Z/NHA5xPpHrtcbH5F
BjUPVslQ+EktSsrCjB9QHJqXTMkP5Qmmupn8s7vLu0Rr33EaZlnEOJb8KlUZ
uC0gPV0jwMYFP0K0nr/ilWq6Jvy+TeDK0vxjQmPNf3hRRrq3KsLU6XQNWVtX
ADwnQY+injdzyLEAqVH3uu/CpNUzRv1QoB+a0Me4LIDIiSpis5np/4j0Lqcz
VU/4DQKJwmurYZh7L5q6GoeJS4UttkpaU/fOf8LKFpgJBF5MX5/ua6ziCBQ4
W8wzStrYQ02oJmL4IgOCV/fGmQr+hEzNmswXQhA4GNt4RAyz7xcbsqCQd06r
IC+B7tpqlIL6XbtDKneB6vHQYc21nRBYlR0orlWH2WMiuW5sN8j7KMOVZmS5
yx8yfGLVZA6BtRpO9caTLH+//xkkNrfjSJj0yfIQd2BmkK0IIxBAAcFvPu7G
eMRkRFHgK5M7utBGxj4obCe0UX6/ULrJ3LT7m/udzXf2w9Dl2aEIYCBuoMzA
krLi8HJWduxEJ5VOYYOTy3W7Z2Vos3NUHYH0NJVFKILZOXbqNHbG9bWIYe7r
rghYIilA8TMpVrR74NaSn8DZSOTKB+moF2cQ0sAQ1NSYUOX0CZaxI1nDcy0s
X+rf5IfZiuUopr5Kg787iPVsJ7LYM62cjFcnr4ZMIvcwQshBI6C3xp8m4ZmB
CoiUTHOcSRtsi/7OYKr85apYGVhg/9PPr14dDhYDY7aUSLaYi9JqigOCZ9p2
fgiVC4wcZRQBOyOnDvWCpNfQvXtnnF/Vy+MGveHcPESc+ZquyM6LUhNtuRzL
MG/wOixrJD4174Cgf2/RrEPARCkcDpVmJ5zzozmYsvs5iD6CsV4vVtTlcxIr
bq7b64urw6Gy9mrxqUrV959vnBNiKYTSqURTpA7HZ60t+gVPZRWd6aqw3h0S
9RzWqXKA3DaPG4jDeqWBiy7jKZSBo4SEjfl420h8eTuX2po6ze4Yu3df8hR0
hcj0hAx9SMJr1tcvQYOSqEqkKUANnO/fEOqHvxNLmTBpQSxgvrLsM8LA7s3O
ox4NGmGrwElpSu993+/Di81Q1QB69ie2psQ/9AexjW63x5HWslrMHdEtGlZo
B9XKqqaBgihnAI/ixLQSN7T4pqjYOuC7Mb7qkvVw65wdSp0XZ8Ukkp0uyFoO
jSlDBgrLECgnHCad+mVQ3rAdu1AfrioCh4Jmckp7BC6fOyDTwedlxDzIPTtv
IcGbJ7xJn3ghj37l1IpsqUp242+bWjDs95jmDCXUh9ncPwJytzu4tjfRdOto
YVDQUy9UTZGBHs7m7IY2HHDMz9G38e1PVY8CIY9g5nw9XonVm1dTXXlqKeG4
bdSswGEGHZweK6Fx081KiZP0GOavwJ8YAfv68PfqN00HKrKrX7kb8i3hqhXs
JlXZvcU1KwPcVbT8slejUaJxcqOy7gzH65uKM8b1nrRDH5+JETjsVI9XyZOQ
L37WUUqZz78DqA1yll5w9/T3Q7cGRTr1GwDqeLdi8d20b3l9LT9tAAPEWrsB
NUGK8nU6DSeTm5S+t5ap+dHdnC4EUvGst9lyzk+2K0x3ceLAuMMfeIkiglSS
1SYD7oHrxxUIcdFOtV5eXAh6i5x4Nd9WJLrnOdp7jomyH5s4XZRXNu4rIFR/
7KVXlY8stZGrVIBEMQ6OCXYAI2njyOYydPWSNiJgFp8oRnOKX0HsZ1u7rkaM
k03zw5wnAqfdouTXp1rGTovhlWBtXXD2HBWsweAnJL/ekrrSKBKjXEqk1U6N
cm5SLYdSBXBtMxsBfw9zQL9waleEOcz7BLo3SEZ1r8RUMfFWLX8mEvy2Gm6w
mLnmeTiNZ6VOhjFH0j8O0hPf2h+5yxrq+ZJtd5qTk3rjjk4Smbp+yzjZKnWk
Bq0swRlueN8n/QVWgwWAqIGaODalOBlktWfs100OlFdZ5VDTmLXe+ps2bNM6
M7vsRaX5OR3yY5ezTmVZo3l5PZDjFd33BlpqYgUYbjYRFfKxiRdr6hvQeQl7
SYUSICcYix5GNbloQ+6NUtWn9hLHXJE1mKWTMh99sT14/YhaQRN6dThCKreB
VRIl5jn+p56Hc5DIWKG6F+5hrXfpcL8469B/bNesixQzPNyhCXS4TGXbrByg
iOc/7prpyf3WMHqKV+7UJhxWe/zMGJ9dcp8cXyjlIAAWXKaVx9LxRzuUT7eW
GT253ow0aMHFmvFDVBdTQHQefslnb8N04mz6ejeATTwXR2fk1sSvqG6yPCio
G2KjISxJGinJdSOxYXY8BFvVAei3GOIDp+fesQjvZg+8G1V8wncxvaqx1Kxi
xoOzZ99KXMasV8lJ9n7cDjmuRwCovjyKGfB9+58ipbdq3VEBGuPihhLTEE+y
zUmEiPGBisqEkRxCq+M5lNxGkpPHtz0rq7G+nYsYd45mZ6DvyksNrmlTS04H
l11C1A9/AZQM4RGzYte6Agd1TyP84w8aFMRzhdmOAQY23QTtTE+DixWf9zkG
JE2HdNHFs2NkBboI6Txy6ePCtnEhs1bhyCZ4ssNlnX09sNopPiTqkcEjsWfQ
0DVxWfXQ8pAB7jTfXtj8zHOtOTYxmN8Y+ERa/va1CZkT2CtNdreje4opfAhv
+a3JqwACh7Xc8N7HH9iDseEkMYTxVwmUHycpkVg6+nyI9xbq8TsGPPFwPg5y
PEAYs5Rsk2i4amKT+VZ019I0omzFqJe5nKnEiXck3bXyLMjTgypN9ZPjuC0F
kpG+RPX6jOvzSOWStiDcT0BJ1kcliqUZm9Mx1TeiX/v+UKtHUHGmdt7uRrUL
Py+fb469HI1g3xputiJaKM1px9rn8SH3NN+TRn5539sniXW4nDAl9gE/pn3+
M0skt0Y/jw/mbYpatukgR7ghqbcK0Jl4BWopXh6cMYtb2ubIuq1FyixggEFH
YTYFclgKPi5P7RE+VZAED1S555ywbLjaqy4agIbPAywGYXLyST/FjA5lJOkv
FaA/IaQ6YR8jrPRtA9Smuv+MH9Iht8Mdd3w2LNrtckSX1zJFxZJH6KYFtSU3
Q7VDvke0g6uCTrd0oja85+oX9DfV73OEJPjEVNNPQqptpkg4PfmS14i9yyzH
U/jJuNgptHHXc0/5EZtCur2spZZ8vaga9poTXlZcXk9GjxgAgNDQUwvNHRqk
uUsuGmWzXnvNmF0tIyaN7VOvgs6aczoDKuWSBYMAtHEO+xdicL2w41XTbzJg
87Bmz+LV7NaD5p2OuJmuZ3tzoUtF5WoWDqUM77IquXqUjJkIfH5/GSCcye+Q
bge8nH7q/sxJVkxQn6XsNVNDmd9btAJBLCaNku8IUHQ5vMILIvOam5zhlX70
2eKLUD5P9c/G08wbjig2GYEs10TvqGFVr0MsryUV3hzXGjIz8H6PpPoGQfJv
souDlT2zye4Lm35Lq/38B5fVm56PFLXemDm3HX5CaiA7AimOodcqPg92j3xN
YXNGX5tzTPSwqhoKd2FN9v0FVzrVH/i9HTz2FWQrYMIvRTHpmYAmTRAoTKML
c6Q0zAmyuWKfjzWhz+c66I+nmi3oQaxPRqruMym6LIuU5s87l9uCMjd4OGz3
G9CfEhnAeZCy3/76PpcHj10PzzyKj+T+IIQQtOH5cz5YqwN5nNnfz3tjnzGc
Y+nOuwOT+JdPSwpcNTRM/HXK0GM9eKPy3CowW01RQL2tVqOg2Jt3bm4SCZtu
r8Mv/iJ0PKwR+EQnZiKRtthfjc1TSAbNwCNQTY4pUXb7uzXISkfHss0kK1KL
GzY+PZNjktpJeilvnwCR7ndT/qTZWdSdHNFbkLbw1MwPxKxVvmTrFishL3sB
f+TogLFlTlcjlFna7Bv/9W2eOa6P50Z2LugxVLctHokBC2WvqIs/DRjiCQ2K
VdDlX0T35rwHHOPSzjlmbDvXEsrljJYxDgA2k/v+dcWVdJfJBxdDN0k9zgpP
fQAepxVmVJ49m59zCXAWTemFP/sCv1+y+JmefBdRQFgGaMQUkGoXbNwep1yP
1/DkvFN4KcSHppNI4SGLqtkEI7+s98PZ+FzTjfmoTO+zq/V/lWSlpz0nddSU
E2X6i1uw0iCkr9cfzDBY1fyONMuluCk9iIy8MHWA30vmPeDnOxW2yzz09N+j
bGXLP30pxvFM4kKq7EDEfvWUxwtAGqHrwsMcdD39ht/0w5AbstdCvDel4NgX
tp2UhXM7IGNCrZzuWR0cUA4FB6sW/VvR0u2rGVSG6RaIduSS5A94AippN0NK
DS7UXlTW2+4YiX9Kkw8Yl+fHUMq+WN7qu1pBDGKHjLToXFCH2FcpoL4oJbsH
SjgQz/EvQfGxpQ8TWZl54xX43TBEQx6cRwHACy2BeSlB5AN3EPDWL7iGqX5Y
/3CI8/SsF/kjW/MKlx4CadC7h2KA1oR/KbU0rt7lTSTDDVNWmWGIqNZl5y2g
Zll6iYMJad40FhcbiMW9SExbNHPHFnjP8PQuHKkEL5eQ7JWmxMxB9//si8Jj
Rh0duDKJyKSmThkgC66xI+6b5FyMFbAGuRwiYNGQ7/XIeO72NZGvY8gkKYpN
qRvDbWQgx7IDzcWSCWkdwiHfDPV68Y8y6BWaQ6mtj3lB14wM/Ar58fpZnqdH
wCBC47GOux8cz13VuUpSdCEun7abfVxpVio3aIQu9JFGjGDP9KJl+j+Wwsb9
sQiFVUUZBxNrtL657oakcIhAQupLPKQQ2909E4in9duywtQm0QKcCxfQa75D
j/TABOiVQB+0PT023fFuJ4xC05zjiO7qgHA8QXlUpgxrnYKPcAO/vRZ+d5v/
yb6/WCB248TvhXyZndiD4xuB+cCBN3Q/FgzQUz1ILbWAVDzOCmR/F2YGrRxG
ffIEhnfVfuHXRdSPUbFV8CyOXUF0qJwHXwbQQzuSZ89lrLPXWRPIkKn4EedZ
Ne7Npo+oyW0NFFDPqWuS8y67IlaiBww9W29i5eEFIvW80JuYdVIUXPdRCPo1
abcsBsxYy5K4cuv6MrQNy+KYlsVL58yV16j8fiOF5be5x7Fv8qGbhPwGcTom
k8n96R4wrY0Q25zr+fLk8y4v7kk3C6GcxOWCsighR4sMM+a0QPLceLdXNtYP
hlJTDTChbjFgqjZrMg1tD7gXr9ylDdjfWp9ni5ZcuuThQIbNJWf2AF1JNfaP
EgheIbEKBP1N5qh6Voc6dbfmRUjOpEVEMP+Jaxs0qlGeCE9q1klH34KzJqmq
w4PUIVTDAjCCJdPDbckaXd3ym5pYslhktxIPPeVB1+fw/CY9Pr6LJ0Rp6UQU
WxSSgx9WsayCiZsppPgkZjHlZsoPTzZv91Xb45Fhyqw5fPVsyRbd1Nd2DERO
ZdmmlA51lW76TaVaLCNnawaKgCzCTeWKf4aMh+b39XouGcqiuk6/9c0dNIzz
OkDYw7t5+e1HQLA1zYlgfpySrDivoRrWkxt1lh1uC7nf462psm/JU8YK/H50
gJTJiuQq9oH4PB9/pmyCIml7Iaxye7HGbYcEuCgLDv4sTzdSm4Pmcr/9U4Fc
/oRjMuM+V25SpUwggy10vWpcNRGkAUVVhidEXr9I/KsSPDQ0L0Jb/SacAykN
bWmXFQ7nfRw9q9iBPYPb1h1ErNGsZFK4CyLv2Z9sUry7sKtvtByf1BLejIXl
PaMXCG5QBB5XIJFDbKuoRMYqJLlaY+HI9ty3kZ+K5uKDyX3LolG9qT3Oac22
1XQ5sZyJnWHYNl569iqmYR0QqN+hyLkRGHUEZwRpHf6TgNc3fpTKxrW0pqKZ
x/AjpqjFqTPJiQA99a/7Wdt7WrZWi4CL5s9P+UAXp2UqO0IEanBQReBuq1WX
JdAkkquhVp8hrOhJAhXkHTQBipPQs5VsLC0y6fKipT5ZKxHGvYiMNWV3pWXN
XcDf24T8LBU0cc9eLHLSl53HoQgbsvze2VY7BcU5BqfdkLiv6W0ta53+0ZUB
fql2A2eWxboKz+vzUQ1LIgZ/K7QpcEp6nu4yxD4ifLk6c4ikdKZv8VUn9cmB
WZQejUGyYs2N2C585hLg8vtPy8kPqtNE0X4G1xvh1pWOwiYM8leJdEBbaCGP
c1y1Pj6ymNFuOHaOVGN3sKtggPIbqqwI2yEF5y9F/Y8NyEMbnlTx/S57FoyO
EcR7RdO2QfKYyu821oKURWg6kZ7pM8UdB1BoQWbN81LSN1pYeI6rPjdpIKIe
URleBgtFPF4sy1B4kF9Xg7efz1vP/l4raSAiLNagFz+ZER8u2zDtk6fZOGUt
iBiabpdtJcjumz+h2GqwybFrzae0IdniUG3iZ1NKezyNuv8m6MvGOT1fFB56
wfnIu7i4hwXHje49/WW1yGUSW9h4X2LK0Ya4f2rHRge6mDzSHGfP0r08BIW5
mK4olG6Oxt5ow+vzMWPd0mIHXs/zqHfE3UU4QrFMLB/eaNvkwMHvXP5/5Gwx
B3f5BqWs0Vq1u9/ST5Xc4o8Np6Dudt+zxzo50YbuTZFNA1ORTXbUTihp4zzd
FUAztSahWaLroDB8Unvxjidb3+GPtfMQXeSBUvDlDF5VQlcZq2BrWkQ4BWXm
ZvaOjxnPS78RK+LY43f81ahFHJiEjD4knAySBq9wy1pn5JEPD8/kpyeO7/P9
vOtcIHDdvUti7ZajHKhcoZxDALLduJ15e3IJ7gEVezR7TjCtXtNbYVk5ETkM
I436ru51oViNp2N/tDAZ0xXkoCkmEnBO4EWaUzFWFRH++o3TrE6sDI1dthsV
5gCIx5Z+lmjOBHsImxhgYashXz/6Q0fg9X75Q8/Z/eoGNNFS61ZOtxXdZhO5
g7uNGVSLu+aNcSQkZaP6Bwo3dMxyI7zq2F0MGmqSc2PGHDkjtDudskT0NBKi
KVbhbNbiYiafWPjKw89ghY+MwNng1H42J6kq/DM9/LmQtEDXeh9wsxn7qxlP
bd5zyNlgmPrDE5OYNWctjheKudS7JW4VvX1Q1o7BnAO/uPvBKd9vUgBws3Pu
FrWDJpwq17+XdMP0tGvUQlFSRkD52jJSqLZ/OSvi7KcwavWtvSffES17U0kT
ahAJWg39+68jFEqdGwpPJ2CFJKkISi1YjHKMyjdQIVSRwoE5WjRk8QX5v3RU
tn/qoYHkYn3lXANvGKzqIM5ZVhv+cuThCL0u4u3Xf3Z7yw6ZaxVSjHW9JLt/
kqeucEhhuYBJNgCe6yT8q+lEhLQ1zUvqrrSR7GyGIXvZ8JyMcQgVn0YhoxD1
yDViize9Q+SfHmcZUAPVjrsl99MOAfS3nLEgBAHWJR+vRcwbELtKJPmBvjzb
Lltfny/vNLHwOAtn7a/EF3Y+7HBKPEY+/u1uQAUrOJ3LHTD0ltj2EGoYBJcu
iVlDpVnjI9iNNEFmNkfQJm/b4s1tYhFlqte5u5tub8kFExq7vJVPzv3pd6X7
KWQZCBDm+fFchWKX4ExacVoil1rQ+4AsgYnH6lFcPEbo+jHEEJ+84dGaDcy1
6iwrDNLyTT+Czv+TWmhX5i0WgDlw7z4ElRL0KoaWaVFLToMwb4x211t5ScgI
2d7kTZOqQN6+YJAby5VxlO4SbZn6Hyl+ydSDQbjGqwwgMHxztICwoNqgkQWB
eGRP3IQvxDMnUphdcYD5jm7yzDd7HzQdlWkoMuitGJfdWnYgr6tSHdopm4/b
6JH1g/9BRrosUdUN0VfE2Es0IWjYZ0kFUsHXUcKWCuzkUTV4302VQRu8Yzrn
vtqK+V8bUSd+oJmYkftVnRjGib/wSOKX7x9oZZsPBtbtIW7TZu7tnyjqqBVK
3kvXKNH+sr9iukjpSHhcC4VnGHLgNFsr6C9czVTGV3+7QrheP1tH/ADu/2oF
mvOK4yq0ZZkvQPlOIpsSMfSJQLfEaGn7UDYHeMZzUxA8smKzJk6O+dJ+VAje
zEb08LOemjBG+hdCz5WOXbCSP1cuTQFgb7AE1pgJpUHk362EUiQvyk3jvdMw
WJi0eUGr1H4NUpJrGuJ/bYstIHEtQP9oOZhLvGprRSUmAXCfxAdX7A47rstm
NaEhPctBXB7+5IsiVMbXklD9Jeq6zGPBeCXVFcqN09pb89oMlfRogs2eQ4Ci
3NIs/7t2+j70DXHddGjZduuGmsOQWHn+gV2p4NUt4sRqZzwbdxYs038LRfPx
3ccbjVRyUCMoPZUMU3DzdXdM4yrVMMmI1cDvihzfPgODLVp+GbKkdVS2yl/R
QMLDexP73TfJQFNQUL8BnKcG3AucaeVdpOBQCCgd9Suc5qIGPTGtkfQlQxP+
9BJ4FfBt5nXRYDW9r/amWnPsEvpacljohADk8GS+2Y3l0gIHPE8nKc3VVZa7
dr5eUGEkZ8HuukFyP/IKygu89V29xjNdUooDvde9VBS5RV5FGpWVbw4eScTy
TNbr1BaREBV3zWv6yYsbVVhg3OQfErl2+HSB1o0F4wY9RhVxueCE1bhuAsjH
FraK/+ulCdAwC6BcIhtJhblhXNztzVkGQlL0sHlh6jRd8gn8TkAvBcEvQEP3
3rFMsm+Tmzrd8adFLh41aN4klPZBQvtze8rL4JFqeiNqltARU5/yJ7FVCinU
A/VeTtzEPF6zaZK8vI6XiN0C511tyYGHIMZEP+YKX3TweHPZT1CC776nMgv8
bIvJ26X2LlUirVconoxHpKmFOwlzImiOIv6PFkXOoPa6Kf18O0ZIryo5t0qy
DqUU9gMsqlCSF1XDqUxhxZsIRJaPFJTw1YkgPKtEijYUAnReMtlzkOxLve5O
fvZflUQKMYmq27JeY/LqebSkCMyVXPTGSul9uSFelyNEql66geLgyQVN8T13
fNIEV2ALJ0aKOSVsnCQW1K3ds2M8vxLgXK3toath3wsTqXa/1Axo2X09LtoK
DiQWY8a2IElRkvzuHKVRnGNq0IRerm8yvr/Qsqqj1KxVrpr84Mvfhm1JrM7W
QYcLmP6KpKiOhQGUdGxop/qYKGdkPnkRgx4tTcwPULt49eEvvgj24ut+rTeA
ZPOJ+f2bmQch2BrTmf1If10EB4BqK4HTl0i6LbQmShacPzdfh6ld1ukMmtka
6LxLjAfCW4kBdcygEoAdtFQqeOEAe3mmLlab3JfPnbOIyu9IYRzu3kw/xSY7
q8vSegJzXEZJhf1l0SGWRc5n6rtlx1FG0O32En40X+EaTjmyw10eDbG6z8s+
lb8jfL7rZwbe4dm0Gw3uGZgW1+Zr5OcrhyT0Q/vpTTWjDtK0VVYkXd2b7ige
IhFQapPksWLdJ6Gz+RJnE4/rLEzXULKGLnYx1bWjcdlbNdZD8Gfd4j3r3q66
2qukYz/ibNK3xdJdeWw/M4601YnMRH29trBrmF3YKzEzl33+pWnC1uBrv/L2
stGsy2aQQh7J8/J6LITGbhqaF+CJb6Szag3E32kyMxz1zIv2OBlXNSAcgqXw
7kCApZHYTgpSRtD8ExOd63zBRnCOAfVYvuXdiiWxeDfEKQIN4ylbRWcQVd9k
Cw3fBfk2PZ4m9VOOJsKG53b1M1oUUEMQ2UMczZpXJkIdSO7pqk3aWToGJnY7
lr1IEtgfxqgubJeEbbAaFCv49eWhdsUJbnzSDIdCNnVCtb3GUTA3dcRJykgM
AsTZcgPNlAtubZR/X28m4/tTh5+c60G56Qbprt3csiqKZVzcEYV4IMS0jyY/
y6H8NqixI9DlHBKlk6HobpHUS5l45sThoVrFbOMWM743IWx2TG6+WuxUB4Kh
TePOKI42miLV03bVp03nb83qesFE0+4wdJniNq/1zN5GS3Ymxdhgy0WXDesP
nvVmRMscLyvmadanaaA5hPpqZxw6Wpqy7tD7O//OqJYYOPHTI0gt+bB03Jbc
U3B6eaWA4xQixcRpNuC3QJV68Dgm8cFNaF9SWcrHdj1f/aJem+zyGVFAxikr
PWaW0bkJe1f2e3HzAvDjMwHPdd1maTKrCypdSfsbwHYBBlK8SAqFbl7/+r+c
h0Wirl5g1gctTau5ZwuuT6vjoAK1Yh9ucUo/iw3CUn2aLswet6/2h5qGLCku
BAJsJIW52as1eGy/csKSOKd39lMf2rRaBAOx+hLnexvqT+cAN09AB0mcmZ3f
zBjjKNDNUTKjA/qUDs3G2x6YdnJl3ddj5iiFRh+4tGGZiMEy3Qp9IWUdHnxX
eRaTlfN8NCO6+13mHyQpyz+UBEnOhHbnQ7H4uF2hYEWgOf/G85jtQn2lQTGX
C8I6R1gpClNSrtrvVk83pW8IGbtH+l+OIM1LlXAtKX/UYS0Ak9mRWVNm2mcP
3insWk0PpWMsYYjGW8Ici9/A40EgSIZZcRkWwneVoxcRaHV3p09nIWRKw0dD
NsoP0424G/dKeT7htvaBY0GOAf7Pgsgef1rL2x7clwczW6B4UCGm81EcbMYE
rLoFMjSlccOnM16zx+88Kv/BR0JUSLIStxekXIP/fJOYQfEkirOQ+W6hT1//
xEq5uKGyAY3NHTggveUOBRaYpSH6EkuYGl3AUgHF8ZOJ4jX3cZiwYglRR2m1
HpGdwamHCr9XNP/nE+olBzp7e59sqdxOGsLg09ORR8nJZ76v0AAZ7IfGWCs4
51NE2LklWYz+spGvsXcn/2YQn9EjtzZHft2bLwA0xaD53PZvfVjScjFJ8ihF
C2PwYPgDfrD1p8mRxp7f9K9dfJCmAiQiXy/4YDS4M6h7pfQpR27zzFcnMx30
8m9JqM6CzWVmiQnWkeW4czm6zvlNx4laFPQGN87TlIzCkc6KdsoTGD+G/0xz
KLlKuOomCZ0E1TOTi2R8qidS0cG5yvGKvLoBDy8uF5lpVH+f537DPDkGCsIf
ZNwOd2KT5Cxh6FgL3uVvxdUnMB4Y2NeL25DuYV/ArTZ9PNmNRdK4/bPSW1fa
S3CKWgk3CksEGq2m2sSKAy4+tWkbkXrC/x9X182BlPZsedYisPxC8JOAKI6C
e43wWy0PusidML6A6ElsG6OcbTOJuabEpzvNn7/kjpMvg7okmt3Ss4F+cj6n
eFfYc/MFrPaktxbchFly2TbhWjr5znnyvPvl5ec6rol6RonR8TxZLfF82e/a
lAYM4sxrsFyXWQeC+s3f1uDPhTqBInkMa9v+Ui/h/PS18Bi5y+HWY97dQOH8
xwBnPZt3GfsetatY42IngIIr6gC4RVSVTMFeYW4zIhQf+HUqmGXiVLb7wTE/
OU0irB2nY9JacRbmzHfP+v+bzqXhXzl5uu3ZqI7PYLuaEO9j6t/svCD3GIUt
BqVg+aoks8uISsNyspzS/F6rAPyJS6JjZ9/bIjNonFK/TsNfOCNqtZi+58t6
0QzdoaAO0tQNTHn34uIYdW8qqnsqgY91+FKhGEzJC9UZ6zFNiNpy/OU5ef52
MBso38xrFzrQEQ6+cqKbyrBxfXXabIHOB+kNeeCFk1LCnksthj9yyUXZIZ2/
8e1RRuUKcYnI5pYVkskOD05KDkrQx0JTMBkGh6/L6r09/XupoLcgmq4UvTGO
aUdgUZ51y3EXizGU+ENqszSMk3eOdN2NvZ447LKmix/5Sx30VlCpbnOkY6Rm
mBN3m3oWwX9zmTnwili1obpwivGURmkqFErWmBa1q3cPGSBJvoVOaTxUGP3I
Mt8OkOD2smLuZWjw9l19LEc0XeICBDQK4XS9ogspYPdk4MB5Rrob3g34i5bn
qs0dAOpsWsPsrFHHufcfy3at2ciQKQzLD9pRQFuRntRsTt9i0XG5wO0sIjJi
F7++O83qgEY6R9izwtOtM10pcJCj4oEy3ZQIV6wTGtsMstPkQwftGfq+e7cj
/qdT4gDBBapGfd8iRvG59eep2Lk2j2A4GaLSSVMXTIsE7BarC9B6TOMG6fMU
tVbdEo70T+cH2ua37yw8pX9/YGEYaUrL1Skwi+vi3lyIt77zhE3riImaA3Sq
62VXGhw3zSouJGggZoTUTggeQ4N2vhE/bFf+BmYtbBtleESuWNJ29ne2NAhG
m+PqAHo/spV8tkQqk4KsJLkdytNWWeQP08hXdyxAt6OW/odZ6XlyuGbokBR5
L2HVSfMDZEPDmpU+51c6Q8IWQUYa+Xb/yrP5hZLXfxwOwulwDsmVtcToaNL6
W8gkYVEY5sXNe2OIEnGji/XepiVOOL0b9y0d9CyNnIp3nG/ubG1Mu6nzQeap
f2gtZXoViZ/gGV4GEkHhYUY5MNUyiipQSFjb/dreH/dQ92iYNJ3I4itM2ORA
kp+lpfEN8pF4P1LsKju9WxaV0sLOIJZFzg11pOF4+BwHJtmwHKUfcdUnOALo
JsHFqLn9V5WZ22IGVXpgADPmY/5kAqOx5Cc0Aa/QDimoJM9A/ieK1vP3ryeU
Y+TYnyUcPITfAB934ZWDUeeB0kU7YgmKvvy4SsywdaY+eyurElI+pNCQYguU
OW/G8dImFN+9u3PPiF+fZZrW3K9anPX0RLFex8kd6u9t1yKLHy15fg6fihyA
nUj1KO45ZQZiqgH1CeDz9/S+zRK2u3xBE3B8a6IviBTRSW5ti5n1KPZgICIw
UhgBoKmkFIpaye0jKxsuEqN9FHsJV8IuRZsD5F77s+nuN/LET4+5HuI7DszD
RKFXRDf4nR2g+inOVVm38ayWF72FqaQGMUE/ez2GVZXUdAmrqOM/kZiu2Tnr
by2fMlID+5PZ2jx8KtNfabdstqWnIUCr5oSXYBX5IYnrORPTRs0Aa0T7mWvx
xnb3C8iLaF4KHXnV1YO1GxynfOuF/yIlXCrbS+nJEZNCes9RP1P9bEJZmW5s
nF6jjq5LmJ9QbTt5S0XU+NFXJID7KZoewSVt3l6N5Jywpnpz3ToB0xxar3YE
otVmHq+M6TdkD2JeXPJ3Xj6wWp5BShVqOwPOgHa3ovDOCZ75t9BaGiqeiGct
B01+30l7q6pdeviXSWKpufQKMIhro/u9I2J6/LE1pfodZDEnfzYgnzOH44p5
65gmMUnhs9hQFgJysh3KcddP7uVUCaKt7fw5TKLg255EGp8W9qjeAgYaXNbS
XNsPc9hSmH7MNsQ7q2a+7EIgld8KyZ2h/HfgLH9btJ1qDgsBoU7nmtURYzfv
+vohJgnH8vhgSMVfMj8eJDqdLeJAckPR4WCzzpO16LQe/w5JAR8xIhvpJaa/
9oHGDqO+7oJB9xydH+a4ncz8PbzSfp9qzP5XvBfGJl2kliM+BV8xAS20A3sH
EfQcPLMPRKNtWK/rBWOwa7FADoNxD6OKbSwPh8VcPwph9F4OIAtaJC+m2cs8
ofzUAOw8oeCWCI+bCMKIh41OuGJmKTpJL/rI4+o6LcPmp1ZoXN62XK/uoEhk
fY6rLweTMQCZr26YXcHY2yLOwIhMq8WWrNzGIkmUOnut2C/Mmh3Qgi0DXLoJ
zbZPCgzgaADNKUPUg//8gWEylQ9CkcPpSseD/kjp1f7YsoDKqmZ7YXhhYiP3
Ld8mpMlkfQTx5p2goItSNLzto5QuCmeeG2jYNHt9P42aM38oBvA5a3Zd7JGo
OjIffs134dptECtSvfOtZapiBaw88Y5xP26mW9lFO1i/N60uUhL7IE1Osjn3
uirEgyOkiH8r+FL4jSZ9PJAv54NFpLxhqT+sfWnwGsEuoiDiVwg/dkD2CRND
alWDTfLYjw8CRMlbqn7BvJlRuXLhJ93PhTHVRuYOl/1kOASGIVAZRnzmc0Sc
/EUA6sVw795aIfOnifZ5DX9jLKun1INiJmEH7writ5VReIGnj7rEH8uvN3jn
5nUHBUHoloU8iRGEe18HAwT9EO9pjnuGhjSFZMDCh3cAjxwvsev41vuBGxvt
K9kNefNvizfdu0vwic9g63eFx8ioz7IQgCTgXgbZ3rDcGT46RJqW87L64BL1
LotayUG7r65IMgRT/DExuYduYoM7RomHzV/f48J+SI+qctqgxIrdYR2XAReX
6IA4BH+J4lhQMYZdlx62cKWnBxovv7fqaVbS58j+txvL4MAE6pm2VsqjQ9/w
xGtZBeFNnOEoJgRoZiSuEssl9iZsHeijHqULdBE/XhmMEwmWElGYpYxrWUX5
zShxTpAamYA6gfPvQ6xz2YJcbdEwmwW6IeBAln/5RiywEEFuE7kNCbtjvvv2
gBEZnZwIT7z6y2YFiKqaUEE8w0AMnofWX2gLMQiFDtLa1hWii1weSsS6HJGa
bSAoEW7y6UitFxx3zGL5BfmVwBfzaXeQfu+F1Fo4OfL3sEb502NvZQfJOHew
UDzxF3o34DUFSRpS75O0LkT1q/EBxOnfxzVM7n1gFiEsiqqsnDQsQEZyT4L3
f7cJoQBk1/W0HZ+bevq0QOohUTU0NNaURQmtjSDgQYlhrsl7x2lmJBNpZA0f
azZZCGLVNKUY7SzzQrO50lGhN8l1axBI79idKN+gG5zDLk4n36zVgIh3LW/f
ntUjw/Sx9U6b0v7u8FVWTe1ZlexYAenbwTsjaGw2OheLGek+VnTjjK5iJn6Y
gEEAKFebBmLkgcvv6k87kyCjr1yUpUgaRCTIoDd/nTC937Uzi56+EnAWkJh7
y8jbiXrhK1vCZ/oY4NkkEWQER6G1/GEIHUx9B/YY6Sg9UEft9wqYn5By9uQ5
yzyqU36R0VWvtb0Z1N+PB07cljaXekpLVReNlyPEa3uQwDm7v8gUJaRsrBbj
dT86kQLHil5/AUYr64Sy+3Xz0nZOMHO7QSrORapySYVsi0GcRU/1tkCmIYWC
7JTgywuwck9acvqGMmMSqlPiB+H2lT9IbCGO531tIQeJM73zTG7gtVk+MtXo
+Didlx6sAIYc+NNsFUNNNqjp8Svu+MZARMiL55TSkUk61ThnDVQJWR+pv+H4
Ubb7wPg+uyQQr1wAKOiBDPg1ywbTeG46qNn6nrLEqa9i2itx8A4i9g/Zu712
ve1EP+xbt9+HXHakYK0T1ceCEk1PLwNQuOQjuMPOOGW878tMNNZ+S7dJAlQZ
8AoQ4alzh+YupEouWdkbMdgLejtYuWBgZMeRhNiNrm3+Q9ebTZVArCN0J8Wk
g8oUblhO+QUVfZh0+ynLGYMn+3EjwHkwo4xfTpgSYRhNbtGFDy4YBIwRZ6FA
9yc2f/Qwd0mEOYxqj8ddNKNY4lhCX2AmoIv54z6tGbRaaqddaSWr+6j536eI
s9uEMtSwVcKPxtewvOIvj4IPPDp4tQR4OjFWb8biDsOXmK2/qP71CrTjW+JM
a9tCeH98O84AxgpyDX0HJu/Qg5WUyHDGlNUWogqkYqIeFaYP3F8CjAdN5hQW
P0BXpxYQRPIqiapdsvXpPCMjAfxYBBp1hiHeOcoLp9ZIOXhuLZJ+dFWDsdeM
KFiaFJ/P9i8jaO8NlD8MXlvR3zOZ+iNEfMv7B+ApyML12q2THBwfUACTc3AA
dyNb5GBLBDRe/RRTPBzopixt8JHGHV3gyNKe2UIqwqRTsEpcbhyStUQs7omF
qy2NhPhcXpEp21X1zzeTUP8pgI8vCYHzz7Weiq9HJlTOwutBeF9mCMYhklgA
gjjLhtngFUbWgtAxIzl5GcvQ1e6vQj+Dx2oBBbQ0TfhVfimXnZ/QvtNRePgt
bB+EZM2lDqkzE3eCbU+PlfuOIgnsnJhw9oN0MKjeIFuq6fGRByTEYZvxzaBf
9F/GfD033qIi9KADHb5KaVae/Pse0XFmHCvlWEqFFX/d/uamZL3ScelrKd1v
AI8MEpZkzYP5DaXBAlTJ1faXjcZc2aTxVrBaPqysX6xC6CaVwtym31/+5DVa
4WbnSTVgA1IYN3433Pf4af5RFCcU6+8EZ2EiN8QOxMpZCyeTVqkEQTJwx+q2
OleFra5UterC55NborWFQMxVo2eJA8Froe/O4AYGnLz47VIGENXFC+GpfWMh
JzWhDEWIj0dQOnB0sZtYaCzNZ+XlqnNopc9rix/nU7JHMkmdaVdmmXmqY2Ut
KFMy3EVzr0vYcj1xpRdPoeChBauzsbeqG01keoVuaHcrHH8pUZ0whAUS2AFQ
AKLfh1673Pup0hY/95JjQLM/FEcOZk2+7N+TA3v+Qfv/2GxlNDEWA8jBnsFN
V+xM9By4lCbc/UbXDaWiNxrnInQOczI78ivtS+8lknn76MVGVVqY4UsYfdf+
MS8p1BgQifBK20cjJdHKHtUXW5ibwI9ddPMB6HxvF58XK11DuumYnpEghCum
qH4d4QyrVKaxa4daNPb09H04rMPm6fPpYZscCbAth+xondxfLLpFBurrQUOL
7V4CFax0fjJiQWOF5r+J3EHCZL6yYDAHtj35b9BK/WZLE1UXoKq+1qA9WuKD
5IOPo+/tFo+jFLaD4+73nkS9YX1ZyuPFhuHIqMVTVHTsWOH/vLLVGFt+xYSk
zpxo+PWsbyJbkhZRNy9XiaopYI2dyFiNYAG7fh8qwoKBwUTYERmU8DBFEKxU
sjRrMvkzR3ylSTNBF/qGKeMDMjW8paE6DBVTfp+K99C+OT2eAtUrsj3YrLxw
f99bPTZvLDBa+H7C+3GAxWpvG/CzWAujxP9nyWr3cWYDtsy9XFYuKBpEthXV
v3tzEaB7NDgdGOg8g8rQsvdzRWlYqkKHcDHPa/1p81o5d0/Dn4nL/2uM2RLk
+HujxsYTwCmtWtbhBKue2uoPnGap1ssTMKu377p4Fe/DXFq4zBS4CX+iba00
H1R6vt0qqQA4mr03Nb84own+2TIpUKce31X0R61BxlYcL7y5fNg63jRGg5sI
a40bKC/Jmh3Nx8YJ5K8MuwAlSZWuneg7zGQPjdY7f/a9+ZFhTRtDnCzMkUSk
KiGMdFfbpn309NBSdZkDZEDuKZvDbOyY/Qs9s+f1/sK6Ztr2t2QyMir894v4
Y6GyKefbOyLmtxc/SIWeOyTA4/Dy85Ro1tTl4aC2OSajzUanVVg+GTSVImNE
XbZV9z6s7kWA0LYmrMeOix6BGkrfvnVhtUpp3L9gFiAJvn0e47P3qd7PlpnZ
aXaKByNHDHh+ZO7NtD8g3ahH/X4bzYdrUjrB41lB5k1MsoK+oXxYxEvOvQN9
S6TAUY2DVQTelzArh8MaDXAu/9EVY8ayJmJ3oDXSB7Wqpttl+HgvLuBAksOi
4kBmm8NmEFkzliRwHZhT/APrXHWQMiNRggkdQ6pfwsV1ADRL6llCROxyvBW3
gMhXB6pX+btOmMTigoQ0SdsO8zVZDOjEXH2M8931v+WZNmghultve1PDq9ko
CX7kJ5bCSwzrqNqldoofR6QWG1Cs7l+tnITUbuwNxGXK4PMHCti0KXYRy4Qs
Ix6m1s5kmNJblxk7Z5fB7kOBCmXv1icpmTRNkEUgrKUO0n5EAnSija2hCZjK
1ccFt8rm0HRgDvxZYzwHswNknyN21K9qMCz9AH4L0c1CvMSlychMrfMuVY8Q
14/v314v7SYHCqnccwJtO60nUgmpGw4vRZdoUQbZ0j1dSTIPDBYr7nPgOSqr
2AIzWyUnETSQ1yH7s/J/q50V5cvsbHrdGIyISzKu0iiPNlvXEnigyt+83bpw
vr7gvBecaLqkOPV1OD5P77hL+xqDGNd5cwiYaZHyD5FCEJT90NaFeF3UmtVm
ZWn/1rnYvIexJY7omPd7ecY9UBliU3Cd6/yM5jkrfDvYReROQL4DlXJ8Qne3
HexJcB2CuK4nRxOjMD9KYDq1g5iAbIPJDn2QdntzVVSt7WS61ePWc6Mlw8Yf
3LPf8HYX439fFwCNky771LU82pJRzhtu4vdgTXWiLo1DV3AuV94fHJ3QrMlD
gnAZslRyrtVxuXfUBWmzQtiK/B5XjRzhcFAn9PNEqpyvWiAWL5LgHZBJ7BLs
dg+kI/+V+qUYcYzgR5olS29etVZ9WOeChHpXz7oLRC/ZWuII5cLW1nB3iQA1
ZVbjKEsH+S5UKANjcA/9O77BEehTqYeR4ekTkjrKlrOoJVn+dIjgkimft7nA
lSOZE7r472wu33dtVwHBvpPbrpjnai6MjHAxb7A0KhHvUeiHyUhuZkjW2LES
JK57JxqctJApgyKZT5KNBksTw1ZlStQvM4e4lXL2EsMRpFONESOz1zE86LQQ
v9Xt87KkV+cdDN4cfUwzg/dXCIFP6K6o/Wqfii7Fp9LIGhPo5FKzkZA6b0EK
iFdBaYLRplbgDon7AF78Y+b75GMrUyiWaHqIkKQEvwCbEMuD1zJ3F/HulIA9
etiXxBVGRtg4HbnZJIkK4UZYlhGvgASsbswikuTi83S7BO06p7nzTVzpX4yf
AZp1RwmB4BBU1FwyeVKVI+R8RrcWcmSt4/p7ZE9SCOOkdzyFregnNGfgmqAl
2OhPSsHcm4NDJ32biGhPTk/YeI1g+XSt58XWOy8gmj7i4L9NPMYSwfFu/bln
qAanTSL1SeWhtPI7I1nCtDxv76qtn71BRSQnG16oU40ThQpx2gD1nv7uGY2j
1htwJoPFaaTMndAAbqGZl0+LkawjDUeAoaIkV4b+pSWSVlcUDlY3sKIlWqpR
tWQAsjgoA2tmhPJpWI11uE/G5pXB10dtkAXfn/e7owUjwQtwhgm6Clqk0Pas
dItj/QiDL3P4zltd1SEGLnDfUdtypA2WWSbpmJA7YEDPxnrbxumnqzNo8XK+
O0xeLIuuh64tbuf7ErX7E6gX2uTL/YTlGEUQm7OmYdzAOtd2tAP3WE1xiHRD
TwlsIsNpp22vOkkThJ0xB/FZcEFahR6I4A9eMyOfKKL/6aZTjqbMklK4A2Wb
aPo0tgQ6P+7Pmq97UstTgf7P/APkOSQOgaydamHegQvaabYow/V9YPCuaJzl
qAWYcfnFfE6oELsDBF6l99FHv2pAS5gGn1l/oTk7rdwsukBhbXWpnx/zJFhd
WUYI8xQxcqc69PPcLOWcbybS7qs/V0hAr43Dr2CdZwprV4E6r2lKftwsDd8c
MLIFo3aQDw89lokvKZZFxheoVcKqOJOPiUCbD5f+/P+5RI0D4wTEFkFlgt/j
OG8iTJ6XMyhI0NRkfRv2OFZ2mPy7kMRI4W40s7Cudo228wYTgFbGMlCmrtqS
rb+01aOjx+3z+vNGDhlOvfwJysncCzbMp5eHBUEUHJeuRVOAbpKbPSpFltl1
d3ug+xubdynGAYP1pPOaPjNRWUscUXUGMNXpWm9QsQqrmF8rnIBMTjt0pPrD
buE2VbFLq6b5WBurD/dLejo9FZft7qk4VpoKE3s3kdP7qTKronpBi1G08czF
tI59Pjs28ZEMkRhSiZLsEVFOL/q48ujvB1LcDN6wKixAtDB/DKnMmxMp/Scc
xHhGsJ/XQIn5AVCOB7oZ/2wDR1V5YPIHjPrg0RqhwrqUsb6+h8ikrsHDcPBC
lNd3sL75oKrPoUaLxVRh/Ocm/gxBEYGbknwTCk7LMAcJORXM5EoTwmcw1s/5
CmiK9J72MqV3nnRkz/xoe/4lI0aNqzgQRWEAp5yK5c/b392IbwGqaBkwrHjP
YYJ89ixSOyY5i/D9m7SvRpwEqC45dz+iO/34UHZqSvZ5KpRMQa4QjFc5aJ+z
5aND9HePTD3Ly/LmlSHnko/0o+bALMG2sStW4AphneQbqVgchU3k+CTpnTzc
pTs2W9QakfLDXsb4sRVV3yElpBQk4HdpsvFYMu5DGua5wyAe3ETxs19YMj47
Z3KVJJyXgsent1pHySftV1KQV7hZPVrb7pWD0DLf3nJ7V/hP364dxcJONoUV
Qe1ebXUBAIyS/jIquaoeNhg4LG2r1LUnCaRKqrC2ea2e0+5/y6d/FHxiCHxZ
yu8c8Keex/ipxzuDwUylBtURWFxknZQzIVXe9PO6xjB95cL347Q6Z1GkD3mx
byKkplFc9b8Vc0/fz0vzaKJxgYkLzMX3jJ+Rwh8WDkImI5OXscrZB57STYc4
O6A+DTNTExa5VzqTKTVbXu6Wzl9ir/GS4qsVwUVSaUlO2uUsjgPkIJxKzu2/
Zuzgf0rnez0r49SuBkfECGY5gUTtIbDkMVaqtV+xSjTbFZU2TsvKs8iM5iYc
Vf1mzP2luvRR5NECTAGgZH/PY0OtSQq7GCM/E14XF3zIE5xlk1lZVcYnfIBd
E2Z/bc3g0Ii5tJdeVWvl7CmycrGfKAlEG2TSmwYlLPr10V7257qLiWTzSD7o
g5vUyOPSj7dVbjuqDfZO0rinlKcklKHh2yUaUilRRmADJ3tIJ3uZKNpn89iD
QpiJV4kbWPuljCGRqMVHMZ5aINahV6jZRMLDvohPHMkCGAcCKQiZ9Qjf4Fs9
vPgF6DlP7jOK9100125+vkZDznOILnCrK15dUGYhyBUgNeBic57AwOTV/rJw
6ciaUld6Kjl4Qh+rKByK4rmaQxaigWphASnw48H3DwOAkpzfjnNxmPIfxYcZ
kLPiSMpYSCfdEGyn6YgMQhYNarsAVJqpCnOvwNw/p4oJBdzdYnTXps3Fp31e
UsWz9w8AlanZ03OucV/Tywj1DCtnhC7E6T4j1w3Zl58e9r6YgZIJ5dZb2UrY
bqANOjDU2qLjiFpgzsEwS+l0VPgVcxT2lceYovXP0qY1f3grH0pDK5pq4hRQ
vpxFYxIubZhN3TpuNNr778r/IfHeCCRFQxHAzbcXq/D1gMoaapi3KGZ8YFPA
UD4b4+qpn164I/3CEmxO6ECC1bAUUS+D2xDmrtsriLVbzEXVXm2C0hUUmlXX
fdanvXp92dHEYjU5Z9GoCCqM1XBJWWnTTLE74Lwe7GF9O5Bc7wFBEz1BlXq3
eGSnm2yIlec0xyXRTJhtRoYXJLzmhVb8fRBt+ewrmIlRXbIQrlW/1P8CwcKE
txenvQ7PNjNgW371tzrQUUl5tQwzxavXOYFoV5xiIwAKaKoV0u+YRNxN6Ng5
Fn/oIm83aidrJXMYRbSD8G3B9HnZUd6gD7suIRlFH3W3xCRh5jmp4h9wDpO5
7T/e3r2fal4M4uKCkIyhu4MeQ86HT9XmytCk0xTQgJ7AzgNZus9GPY6EYGPp
MNXKQwU7O/Gwk7kduiN/jTrMq1iEUQA/jh0YYArIsGsC8R8octeSNXEy5ppU
xXEafczkc9c9A3ruxTXQ2LDtvHvKDlz1h9BibXeazhixMDuIjm4VT9vsVWQQ
siBVIpCohLYB0nUXh3kVSTOub0IwP/oxs5KlE6395YgX4AKz8g+OPSSX8HU4
6NLPRXcGaefsOyWe/0SFpEpMWn6o7LP0z1VWbOItpHEHkjauUP3FbkXCHyUD
4pKJyLbXCGGHowDpYpIiPyQ61FthiinRgo2FCSsoU+cyIhz2PTI3BIsrynrp
+WGUmXzC4TCE8yHBwSkM2WNIHZbQLoX7JuxZIIC+ET6SN8sgQf+298tXPx4a
m3h90pHs2rxhOaGpPnDyKx5OO2lkafj0nT1EDVuBfUw0zR5Laz07wctgThh4
co378Lq9oIo4bvZuZcdyFulEZVcBRjt/Ip+mYe0ut6Vo427RRBtrIb2GZLJF
bGrEg65+2p3qODEvtq2tCD3Avzy3mP/g4fMfNHyl6R2V4M2e52PvxBc9/LY3
AOTO+qIpeHQLi/o3YxpJjnp5QmwLmi3VFNiCEiyBe1PKnsPub6qz7rzNQzFq
gYBEKxwQYL5DZEyqVY6o0Axzort4Zyh07J4MZwxRtONLP6ERnG9VBxt2BePM
lv0rIVZj7FTi4v5cC35ADLq6cbqKI9df340/exJZ2UuDfNXQBopQFW5WzCUT
5wLzR2RSCKdC6ecGqFZeLc24CixuB0hDrkydZzJLh6kX5pDSDT+zIq2B+OGc
FV7xGtcvbHctvUxoTJsdt5QlXotNSBl+IuneV+kgA4Q9esv0dnFS8h0hP2an
3Yu+z8KBGCuqWXavMz16lofSdK7AieqapHMfiNh7otyZ6s2MCaRqaJ3LBbvJ
ks8L1m1rneK0dqpE/XIS+pExoDuK926zoLYPc9TAjMESndbPQlHFcgTusOft
8yIBIs30U+aeb2B9BA9zeIrbdwC6KMqO29qfwSBPgWXDHE7C5OzTwZB0aEJd
jh2sq/LaC1s254lSGFmmADE6vOgFzXkceeYh24610cj+h7Y4xB01AUpMhlh8
FYOTQc4FnIlKF/OfIGhnmWgUyk2yJEMD1mPZF1QyGVLD3AMJIf8MvPFKe5rE
+zChtIGqizcBddibTkIqN+xqFJFqG8VqSB0zkSyGCuNOjJLDryTInuUnUdal
b/WPP7larmXDajS0Yy+Em4q/aO05zrDmyPKE7Pt+IqX3ZuRuiDVsAVPFMr3V
9jK31YqL9W2lDLSbelXu3R5oD0rVR2T+bedgq9P8TdfPs3l7YwlMA1/BDFA1
QYqDUOZZDj9Ta8KNxXOjTXmnobL9IFTurcFF3ZqCElpFVjm1vBbFeaaLEJHq
5pVYJomoJWroS7MRzIYuZjHdFdvqo0UrAWiCKyvaG/9s8UZj9KSPM2PReG+h
2DmM9PUhfxckmo30sP5083qJTwdqSIK9zRPhKUzaH2LkZmvV4g7T4hSMKXfG
rPbLOZiVNW/P5DVqQivK8X/y7fPcmKqbg5zi0Se5m522h/A3rYdIGPO/XoRk
k0F+vOv6qBuCiO9bchhU6BnpZ2BZgrqLAzc9dcaZSTigaoLpK6cQ8cUbkvpE
1gpU6onY+HrjvgvVDiLGYJlWwK5h4aj7Dxg5MXN+M3Lxq02sLbj1SmraiHdi
AnOeDY0fveu3UoYdYw8rqjmSzM0aTFbvvEm1R2i5ThOH2+//lrMO16wTQvsS
yKkDx8Au04PCHF2K+RdJZJouPrnp/z9Yyi0dqHSa395lKOB6h7+ukNlnADXW
f8UrAvS1hEKyKVZeXApY+5Rr5t8zafnxOm7EuB3ylzxmXfXhReDb2h5iMOWS
mmbxsWBRenj4ZTyrW0oxmGwNVp5eBeetMzGggjTy1U3QUch4QltLtq5iikIu
iPOA/tqwFnsrENGv7z93TPBM+cV2lYDWykAdhlrTfRP5AD0Gn17SDFRxFF08
uNKzCNwolJVCnL8xxizzhBZTM5IY7Ve1epM5ZNRMeamu8cRPYKZXUmigmKzh
inybaVIB67V8wWY3pL1CEIGZQNTUDEPS8niG8nYiGo/v/0OB6IlfN0h+7qct
6XOOFJBLo04N/5XvGJpV/0Cbq32TrRw4bl6T6Lhpqj/uHm1e9AsChOXPGM6n
sACpPbePpnAhCP2wt5bvKNjr74tEUyoTUEstqIYOw05jieY6z20yyDxFp4+b
Nqr7aQMyUMfrXtbnvJCpA9YbgW1ig/aSrt/o9I1Z0RIQ8kCHJ7Hm4hSC6SuN
1ORoLaEpRvDhXfCTtZXqN1YJvQJS38o2ha8MiwcQs1scv8J8XgY/ExcXDnIG
q/vkuerj1SqCtZ1iRsm/wQUZRt97vJwrhv4l79NH0NqlArBRk25/FAsygeen
b+JSoFqqdC7SaBkuUVgzr/99Z/hU2uZ0i9e8JfX00TpD8e+NsnXAR7zJDBVN
D2w8MGvMGP8B2xR8cJuLsuVn3rFtcDLd1I9vup9HeG6IHlTBHa+rJJ2+Tubd
Eyy/8wYF4jbpt/bBnc6c0UlsoyvAsOWKFGvErvVMpGyN2NVFJQMr8Env8QRf
UkxkWSvtnU9DsKd9U5etkaoAfmm1gpPcOlY3uznH+X9p8dtHjXa4t/U9gxDp
hVpIf9uuXz4dh/nbSZrOpEX9AMQ6EiBZod4zf7KJCWCDls3zNDw/1CmgATgr
1JEUEI6pfi3+JHcbib2DVhUQ36Qji9yY9QYgzXV77UxbvkZIVQcjQziXFEKN
Gsn4ZlZK2GdvkfZYheLlQuHcNyiWpi5MYJ8Mp08vUKXNJc6zNUIWT+eiLONa
QdAiddagNh12vXKLRh80IdGIAFCV4uxS57I0TxhD67oyRXMQDteEaBpi91iy
eqb7sQXa2ALv+UuJ8CiK77GDn0ksTXuThhDonqsXc4qTeAdfxgQRxSCrHZNY
b8yuu3FnZSpnD/Bx5s/IYfA1Va3iJzEVjaFe6EP+2Fb/T0rnyJSwG+EYqava
FKVEqEkTThTq9js12qHXkz0nzugLbDhaMxu8EgiJr3fB5dihjmQEj196mJVz
7NsHLCwZrz56XCm8xeqMIuzgteF26/9jSS1CXT9YyRG7kBGlxzuF7r+k0PVX
X0cQeSCinglislJ4Xb13SnAOTWSVw+9v03TJgBiW/uRfce8idbj6F+XZWcoE
IANy4OJOM0MyGI1WhvXsct7gTEAsbKWA1sByz054ZVRg28XfuVfN3eckZqaa
R+5sPB9N0eRk1MEMAmZG2RK0Qhx0Qy573CRTc2aIWXfy4Ffvf2pm0MnJBMuk
pKe1GnKJkF56ubvC71gkvufWfZVpsvDGyctRxZ6wbgFAOtYgwTTpu1QqGLtY
DcBDs0mpKUJjeYyz9feA5KCANvQtyYJBVbokLda148EYnDnMn398uC6mWLKu
RhzWubJj1mA6h7aF2eVdhFzO9HqPzlaxnuBesfU+Z30bbPyrv/l0aRluiVtz
Tq72UDoJN3xhwfJSkH5gWZx9Qc9Q/l8gRk4hqY+ce4x4hvsWlUUpAtJ3gU70
shIUCMAjdRn2yjkWIYrH4G8Faho5J1Su+0STBKmbB1bbl/pIDRRWNzT6D8SS
xwIXOVHTIFXHXrq5HLdL4MBJGSOABczZmLLRQzCvxeHk8NFj2RP4OS+YjWAF
AaTgMumK9cA6b/H/3t4YIT3d0oWMwH+VaizXGYS02XcAYTfv6u8GhlxcEOF4
i9YBI0kPuJjDBNQq0thQzbw7/wVm3QxX1nnPgKIGl2y1AkZfX0i1BXeVgfk2
lbtIt6ELG92s8D57I0xs9sJTktjYpdWha1jbpJ3iDqMyb/jyuka/iNMnByy6
cyHZvjCpR0R5reFqZ5cP2sAtLuVYaprHPwqehNG6rnNiOyYY+PZQS1LvpMD/
N8S5aMY3ouQnVjFxEPzptw3Vz1mHIPTPi11HwDEGD/62cy0IRvnB8/iastXe
sHFi8Pc3G2GlXi2nNW6XLTI37YwHl1K8yAVAXblWzaKO5YB7Cg5uUG3ip3A2
awyiMgVEr2M6J3kRtbMDfZbUvgif35/rudW3S0sah/7xsRJs54ZMRqDTe9oA
8al6YZRRn6QWc5WDNu7JQjBPShkxIV9t1eISMtHosELKtxnys4tj4DTWIDYO
ZRyqsweGmCpdg8fhj2sLnPkECdOZDwce2qC5PmhSbTjPrNX/0SfPOB8mawnx
k8X9Iv6Y1bOwyYIByLD2GK1BfBYimdIC5fxFa+qL8+wlVDIX91vqW7kR3jQM
nhxjNjOHQIZCfpiRuekNlHDLUcRFBzPIVGl/smsecpQ6ZvK1N9+js6qdTu6x
b49zuAiB8nWsG6AuiYOfR7876jff1y2jyVXK3CR2P9DroUmpL/VQAx4ae3B2
Y3YBnrAOdGh7EsvZs94d9WtafD+zvVd1cXt2jLtV9hPRbTTWyvMpwaz9KCYm
Z2FAtmDpboaZ15qk9fH+r2/gMK2DQc9VKUGArtwwxxDI9/g/xJrk0fitlHfl
z6X/CeTld2di2MmQfHm1HDSPu6Boqo2Yu7yVhz489o/BAs3jmUBQ59UF2g4w
EOxTiEhGPXjGKhIqXrItWG6dkKRDZ4jNfY0WJszedQ0LNVaDcejs6QwyHiaW
LWRF90Nla+AW2+Ix179rQcKxh7tGFSxkt422J5RlOLeMA8MKu/Jr3Ikd3fJC
TeV8Pz4pQ86FV4bAiNNetbSX5p1BYbmPt/CmAO7h0Wfhvd4e4ty1b+tkcgyH
s1RhmWasvxvWJJsDfCOlMVviLdjoeld/ERCimlqkFnV5E3DwsW4GxA6NBBHr
cN8iezuvpqdUGv3XFECxHaUuhJkgdjz6ciXTEQoGGT00la1OSMCw/GHkv+yE
IpCRn3tPxF7gSSWL1LueuH/X9fv+lP2wtPL8KmAk+TDlw9yXNUwvJKlsZYs4
yjp3ULeHBTxAfvOO2+UQBVf201mSq0h927vNJri1vQvAq/h75fLqp/ujDFkD
3xSkTs/+NkxAhAQ+uQX/5q4TUjKiaINBRYcjpDIvA17ydBvysug8kEHZmuW4
2QWpzh/cN+/KU/NmFHRz2CjUVCbJZp3gC5ZKGdzdekAoMR3/zCDHo38v1JVR
GfIXXhdU/zWqWEDUlHP73QYkAhjPjw8DhcHk+/aADFvDaaz4qAS4F4KTWMcG
vBg34Nwte8647Iz3yF1x02myvtybKFgVtuT80/3esdpygeidjQrprAbIK2RZ
SWtM/pzv2wZJlpZG+3dnkA2YdGjyPAfTOvJdaiAW0/KCL5NFAt9f4TJeMTRm
LP50zJEZYNRTook91mP6zDxvG9tlffiqJFKmJ7jOcLLBna1iwhZatEch6+C3
HsJtvwWgmQho6Av+BOxU/yXnuyPtxS+xat10ANc6gE0zyDYSPRKIJDWgiR18
5j3X4KOFcJBqNEvez7rRo8bMI51e1leBs+Z9uRhaMI+RRzATxD1cbGCqLM8R
ZVUJ7bPwk5duJlwF1SerGzQIBKdkExz1mAaJln5824/xJdlHWP84LGfI2J8X
yNooSJnLBft5sJcIRUdNxNhu6wNGYtDzoNQZRjKWrKUc5Hk/Q0l1g9P2+5RS
oyX8d7GcSM829z29FZ/uHVkyVZdXdb6pui+5+Hu+gIUNqv+uaxojhgMGEt6o
ij/bpj2HjFQAc1qzhQeglwthk9nmj47i25QFJmJ4VBoNtEYW/9ikvsFVp8mt
Hj1U4sKUEYuTtBwoClpsoQQZeUSNjGgNH7coNN9FD3mkq81S9+OkIBZPBYqC
hBiixGMdHunJcZNTdJpEtIaip3AV5cshv36PCApSnp9fv1dHrpJS2gRrJFYW
2EiCvL6O7wjW7UI8nqwVAqmOcDdLj6PLLgzEgks3Lh5rHrBtLWasTPLABNHM
k18bH/gZl/lJOEGg8uRIMYlmCf19FpcycG7oMK0T2yY5vW0W79UkEH9HIKhW
Ue8ZAnUWTOPjIER41IzYEXu/83HrW/kHgxecLvO0yKY7GZZDkHZKw3A7TuSA
K1LKZcN/MYehYCtc5JQs1QXbLS8a/DwsPp6/SaNdWxUtHPwQtCdCz8U9U1eG
d70nXmHHXka5RMTen+TWqKcXy5lyiFGKR6Tv2coJKLOz7gBLhqkWgkgbocjN
4/7LSP6pHPpiAiRdv/JkLFfsgAwVL3VZMisL2cfZFufMxnv3Pp3XMEGEvq6e
joZ3xrQhOvVO2cG1s/szr52NA1aCfB5F/Fil3hD35RZ1UtemsN0YEUBMnxLP
FceKzpx1tOf+jqSUPC9u3C1NMF1qZtsE1k574JgycirunsSl1n/z6hMPaCmC
9+CWkDS1fPNiN3UqPNgMIDigfLXT+zjEBZrhPTgr/t5EMi8IUzE70HUoGFtn
Fx7XqvdzSKOYokx3BdMtPOGpS6RSOW5/NZhy+6a6x3qLUnafXkr59o7OSmu+
cc/vmB+VTzbSP4VcnfMOuKYqCarR1WHsTzziDPLl2uGDzaisb3n8VK3o/zo2
h6ec57815tVHwenQlmDvjCiax+dO8GLefufqWutQDidmcOARNifJJyXcQyi2
XJ+lpVlEonleeCYYUpq8wyp6iuWIaP4WzVJCnc0c4GZgvqAn9IG17Fop0+OK
GnE7RUZVshu40cEeW0FKEQjwh8WY8CCWvPo42PK3zUYpFDInVUDW02qtZFLx
Trm13Bhx4X7gC50esBq2sRr3Zh9mysObW2T1OMTfrI+VV4LMWCxtwusVp6V7
jtXhvctNLC8fLF7alUhJFY6CmEVHNpIhmj0ORkRACCSDpPB2nPmpc6LMoes6
xt/AYH0v5ZqxpFC9hNV6oDG/+fOXFGgNvy8DXkr7yQNe5qykcfBermpdD/cQ
zxwOYvuU8f5Fl9mz1UiJvzQnVKIp5TWoeoRT/lu3QbtA0Rv77ZvtnKIoIPM2
EESv5FNNXeP7pF3ezheJ7a8We7VMl5Z0k6HspyyWn1ludSEs+xAjcqt0Cv7M
wznhh8jCgYQ653Shrrsh4sR2ER4fhGz1kMMcVrdaxUIORVEL3WmMnQqHzTBc
Lqfa7PBCmDN0DwgKfqajBUxPc9tir+QgvlwafeF7RWWZn4RDXubHokyLhIy8
cSU+zzRiO6hAkJyn10ZepZB6YslfrL/lTSVCJ4cntGDe8vid7Ii7qQkggK3H
Qn44pxFWVM9ffbfmA+Ic2mTu2JOQax4+SOTE6rwaBaKlrA1/ZIdhDsqM1YCs
Dk8fnyJjg8slDsh0kcFIFENX071dgaXBlJcN/SUu7RFav5ctmQ9RAuzM1ChG
E1F3kjVYAP8afikDxbNCla/FISxZJQBS6ctQ46vomwyRWgYLn9PGXP65eQ8D
y3uML2+eHVJJYIN+MhiRZQddTvod5CwqF3F4mDVw2NYYxdFUrWupG5kheLW7
kpGATZXMsgyyGYI75cVkSVQvzqO7nb3PQijdFoP+4TWTGVV7bu+sgRYwyzYc
rAukg7AX5IHCN0sZgmTWH8Zwp19t4DzS3NOEKdY5yj4SKN9aWHH6JMAQg2lu
GwNetY/ZY+gh1zAaTTiKUk6cYoRnqx9Yf/iAkacZzDEFnMBJXfAJ6Qkz4F4B
0Jky8427nyErgpZk5/TAKnj6ibqIcQlNs2aZvAzA9I8CeLgM1u32q1Sv/rJ/
QE/OnII4IqwLSHc9rX/zcCKjpfiTnjZ1YGWo99iZqVoYbmIrNKpnv+JlPt4Y
n07ExX361QC/c8dKW3VeQC+Z7Zw8T4iJkAwU78cRDYILS5ENE6GQY3tceLdG
a94Pbg8PW13lnpTXZLGGAOFPDHgR8VwgnWyQKqgcd/dw7YXln0xjTBj4YLDy
9oQkhYPYnJZmepQg8+xYlH0qG7pU3nGwS+4kKmySJmANhkJzlJcQUK/MdSST
NpVHFYQZ+sT+h/IhMuD7u5NO5eL9TDgwR0UJco81PonHNTEfgJbRd2vft19k
0PHxRObt2TlTmMYgKiq0o7aMcANWSEH15fzipz2Y90MuUAoQtL9Pa2q4fABs
kGtnfuWrpyu0xjeEN77i1qQMviSq4qD1UJpu5Lza3IOPywv8nEvVbgvUR9P/
5fuC2Zy8E0gsEZ/+Jvuu6Jt8G15JnitejrzILSIwVb5LKnLfDLayBAg2Zx8e
CFpknzsWanGTNGQguSkdAo7d123lT6ajKNzCcYFZt0Kz3YuUktUq39izekm3
h5u25UZDDlV6htDF++DJJa8zH6OIQ4CmU2HBm/EfBilkd+eriAB+qbJBNG48
phjoaF+sgJnOe2bH+9QZxRtoaWFssJxBr2HkqtL5r41nW77Wj3V0d0KFK6BO
oKzzRfPUtwze/4YPitX6qyvVISRjSXv9ESNrehjuM1mU5si5looivuzanSvC
cSXRGRkZZBqJb1g+h2Hwwe3w7YEU9uxUvEhNJ7SM8xxP/lEJMgJk3G/o1CWU
PGt6Bp0GhPbSGSm8stnnSqpccnDA79k2F19+zwpj+bGloWPhZQiuGHWeG8A/
olfxTfjdm4sk8ZP1n2o+paZMyRaIfZNC/azigOhN9E/85Ld/fyPzDFfgRuGW
loZS4y0M2EQ8uVbhDaBT104RhzCJ34Y2rK0rXwdRkluLtxbQNKqOGi7SMsX9
xSm1Af8pD/f+obakAPdryz6Zh5UKhYSeBd0zXgpai6i5T38UaSRCTGS21J0Q
KeeVN1J/AzIa5n5YZEz3vZslOWxkGfvuhMpo3fTOjyfP0iYO8zLX5awBqb4L
tPtgYe8vJIg8SSF6OvidmRPS/WCAU5P1BNOQnz7XcfVn0YEOZT0vZKEZzqI/
UwCpQcOdjnMtij0ox5peyt3MhrYT3U4oRu/pO0Z7+RNtOVkQkzqBEkohHDP1
yuJN9+eaS4yF6VOkqvgy5epcqgm9/THgj/5TJiP+nuiRnNXY1r8DUCJ7kin9
rfuClZm1I+KB1INpkgC9Gr8e4ot6VU2Sug5LFImqtvvI9NOM3e6y1pVek83C
SjTX9g2X918CrR4TvJ6oWBYIut7rzSj4yJEZ7vbq47/V6yD8YvctstfmpV3Q
chDdTdZUoC8kFbmjJxD1QX3lOftWFUfBiotWlSd8jCwEoFYBat2Xzn9qOQSk
CUyOcUHiP3mKFm6uXqUQEmtXAyiiCsWnb2CK3K24yzSwi9WyeVFtGaS4oTck
QiJsbSxGqrlTy+lmaqAihvc664S3FpCJnwQiWaxA3uzFLMGO9f59tFFICJHe
j6m9JI74h82gozBqQFtsLwmTqw3IH5D5yJ74zUep7qSWG5fzxVW9vWNqK6cc
+wDiQaaubLKTXB5JLy6sA4Qzzw3XDo3K42GxeuvZwaNEL7vAZQomzd/F8Lrq
6YZFREdZWTdCjQ8ESoB8e2R8SjNoKMhzvfTdK+6muTu9xgbbaW3BXdO+pSCj
OjVazbaZaN/x8XmtH5W30J2OeZnjbf8bi36H3bKwNDxYR/iTsjVauclo1oV1
gQLA81Dl16ywR2d8sPUgeNnxZ2CAS/DyPQ2ScHq5YAmJ1OmDXY/+/0Sqz+ka
yIzwcgHV4JZxVS/IjfJdcE3O8qk4mYF4U3GN9HZIjkv8fKQgVBB2K6YXTh3j
uZwrelUoxg3rhWTow5VjZYxPaX6nfpSa4tHQQ2q2Ko1uSflMIkEFr96e8Luf
3ID3Abt7XiP9UDGA9rcOuF4pIRU6BT/T5KHdGjjPGPxRh5Wr0Sa5X+aaUO8k
yliHAmM20ZDgg9S3C2Sel8f3bfHwXRJutkHe3/l8ow81d1m0dmQ3uWeMOQW9
EtA6TbBOt1BxddCS/kT0XreGLETclWNcNvYflvRlkyNS4vsPGxTDzudSnUxF
WiJeGZvOdf4E0AJQoRW2VOOtyI+1pXzIbd9DWK0M5JLRyz6lx/wkfq0jO8Xc
BTO2b66LCsxtM+uwtEEGuJ2ykTcXlqPmBVQ7kfPFHFnzcwiFe6Fd6hJL+uwz
H75jZweP7TW5AOgbjgHLEOLJQQR84eaFv6pN2HpQov2bu5fLW1k267Sn/Txf
LLt16KNtdYnR5gbcuF7lFiDHF9R1tyobVOTqLRgENRWkXb7OGTjdsaTQrquc
3lJVQYMKKG+nsSMxhIRRwUJsN82VxkmeP8HIjqBFThnw5tONcjK9rV5EVEbj
ioOklTpZS28+OFT7OxMtzzflkh6ci/67ISNB7HItW1HzHt1jkKVYAzeJvlJv
mfk0MQQmHW7tSRNF5ZVbVUtkfVauHUxvTxkPNutBl+Lm7paayoGMR9SB5nxc
0SmcOAi+Q4MKzvFWQH7ZrhIe5rAJ+0hznsY6fO+OId/+33f5nXbsRcyMXdLs
dEIjUvg7nKNrE2lDkx3Q63JuRIzZaoaYSNBsrwzn/Xl+5c+AaBt6D+ap2inf
4XdS7TbunJwvaMOwkdN93b5RTZc8sFb7kp+C2bS/GZnK8qAoXa7/QuzZW4Z/
nDFh0+9b3tj5ZpAPJmwnlyrqwwyXGRn6wLmbdjJURyWWfdVxRifeU7mfEuJ+
g8OI1zRdppgkFnA6PcdPcLwiGSvSRf7wjp8IDg/dk3sZjgrKE5Lpv7FaIuEf
VNzrg5llk8O2vBenWrFCkwd73kc9C1ybH4sQIGxHU3Ml/O/3Ut9yefJ6PF0I
4KAIh7s7L/So6AY9iL4SPeqJjQpYq2aJ7+Wit1ZYDCl3LnVpF+UQl9gDPast
wJbZ/RntQd0QLQvIdkZPkFRrYZo3Xse7YNkL/Z/qieAwHSWieP3w6CPtMwLH
Ylqzg0MIVAuYY5c9lhGUfpvXEx/hvciMZ9ru9yhTUTQZ0YVxUFo/TmMcBHCU
cs1cBQlX/t8kc2kvkakbRB8BRnw+u0UWFotKulDjbv16FKPeLTHNcjw7V8Fb
Q++osgkZNoiuQUiKHMqY5pALjZ4N/DQfYE4t+/tGT5otpyVHDsLTTpD1nBCf
x48ZHy2zoBp7dv3DSH8ll0uucjM2mANYtuM1kgaaBzCHWaGe2AZnz5j+j33S
fxVNitd6zx+LKeTXaSCQOQu9eCjnzUFib95LQT9Ls1DvJOr+ITQjNJKPhiZ3
TkSVvtQmHg2Z4lPRQVbMntdJcB/kRRRIH9R1zyfvhsB0dbJFaM0jV8iUpwQj
IdPPkXJS8MIH83ZtnNJXt6sHwCQoJFSyXpnz336f205wczeF+RvcaWWhVL4L
iTeaPl7qrbSUskHlVBGm+BfoRgd8IlqrH9wcPhCWV2JrRokhIeUKLixxyIrF
/UpizIO6ccjlKiQkN7JCqTyJifvDdl04n04+Ew86Ixc3+4HzVBkZ3BONXXO0
I7sYL6BHYwvt4B3iQVULJg5bNzPsWQX/OXXa5oQaKBQYzZragKJcFCIf2XSr
XLjnD41bS4ZwOle3wMaypXQCld9kG84HpgLmUngMKHsczBgFrSUUnMWE3BOH
TxY/YIrTWuoTDM9paohXw4THAvRvGhbi9aYPcqF2QZe4TerZ0Oo5wCocJHzp
JgOaMbEv+LXQzTDcvyTQ7pWkcXxXBh6UQe2CRXwodWqGS/Fu0RTAStnm7nDM
AuEjFwRorhfb0raKJQ2bwumLgg1muPbphKoygjqUf7E/BTKT9YjrLwS3yyMh
SNejkIjXUKyblI4XZgtl4S6KgV2hQVLhwI40Hhp8BnwrZUu8DO95LPvUQOwD
qAzK453hE0lO1vghbVqkj7zBCPOfpSbby4md/YgiICSUClzodTEa8oCOciq1
tnSyWhmvnaOHqZv4gN8YFYY24ssSSCdwZqnx45odCtVHL2i/EU3zw65bZulO
UjAyFG4IfMZbUnfkqN4OgBNsChoQbrs9mMuhNuYpuLfPsls69BHknAky227K
7p5rqpAzm+nqZkBeOTeYPLFPmqgEL0+9Dpchu3EucYCHowtI9g0b82Klxz6q
lRpyCeylPpJJWNGBqNprpfvL/0gRtQwsxBeSmN76mN392MjBOM4LehYto8KF
hYKFdb25RjH2pJqhFthN96bpqKCc4WholSq/CQIphIoQa6AtrKBlykrVhaam
WtUkP6maDTFwZnm8FWCZ1Mo52KJGeDl9DvMoz8f7BcL7IGa7dZvzx26eZFQ7
LIBWC174mHx2HSYLfMuqO6gtUEcfD1qFW8NoW5tCq5hbGS7M8r8K0KXt5sWW
axZqMrA7P8PXNAIXIqocmQISkDUtKMoR8QZtBL2NQA7i7FQo+ijbIdAwNeNh
WyccJ7/zLPwcQ1v2MV+8UzXtZ/85el1CE5qD3ndasTe2+vjAgo33Gr4RcaNG
eKLYBdDEFwLN1LbUwxEEkZifvjinw68Pow3bV5RqCEdZrpM4+N8tpz+6+Q88
K4XN5LdqQ998WkJVQ3T1s2uPILI+DXdIwMwVQB+D8TE7m9ylIz4CwrN0AE8C
ILu20uQzsz2jWIyPlNrbLA/An9RxzANkoyVPq9D1/1xxhIQDmdVgSq25YKoI
2ReJXtx3ZeonrCNgOb0mvhOVQpkl0yJ2YTqUaHtiSLyZ7oYD/X8qYh6TAIQS
r+vYvKOCtQyQXQ6mihMMUpj3qJdOXxA1UEAOJkYYYLfql7cSwjetWvt6YiHr
CJKIJifX1VcE+tzKYYgH/bBrMcS1n+8fy3OsM+kPyuP979hpUIkkkQDgwAoB
fW219lvE2sjKzRj6e9JY7TJDWY+SVybLFrtwjHltxz9avTkd1zRzqd59yTnt
fnPYi66Xoch0jH2iDinOx8f0LKvQ/6ymxlWzR0mZudaFiGQF3MnuiXGFrls7
gU+I8QI8nkrmehfkgfMdj6jcE3StB8iByHGaO+TvvkbO+W+KegJEHlRrYjxt
8P0QPm/D+Ch5vyHG6VAn5XGIzvdhN/eS80BuBdhY/wB+QWpqUprQrlFAhEn0
PqtzH5+rvEMVwlPIgx2lXqCtXC0HM7RsKAv+/pUp+zmgnwWGyUrU09vHwlly
fCG778iOvfNFOELlhiKOfeb++LsvaTs9ko7pz03cZeAZS+FxBqfEJchoSyqR
s0yWCXl2fEEZk1pla44eO4mlgrUwZ2/yv5rCnmevFDhY5Z9f8h4os6frQr1y
Am73IT6KKWlNP96qbSH6cGKNPgBNhnf0RycZwp5T62ci45X/fb8FvQC0VqwP
f79PFSeMIKZGru8Zk9ok/YbobP8RLcHv0YQ+gAhfrvr/x40fQeePniGjl3RX
QsB/7lSlPHFSCvlAe+fZBbzTf5L4y6NAksTu2TlG/GJUvbn2+c1ELVUlGmY+
c/V5drZcdvKti/5V0IkY9BuI9HjwyhHuTg2jGzBv5YskBibk9X5forGPmyhV
uagVL2ynkQaHPjy3o7wjQKjTEdOhv+rMSUOiNYmPqk36yY5qayNcisBBHcxl
xTD/cB9jimABqRSeH4ae4ugGEk+fMu7/mNvyO4g6XjnkxY5tTQPpAJASgTF8
oB8fQvGDaTDemYxKTTddHIBu+ViJ8zFotmuENwT+2/2J61y8JDnGAteRDWrG
08ekPWkZHSD+53R0GBAigoHFLdyrB9Cb6Yc6wcOULskPrBCM4d2FygI8Bm6f
koW8u4nwMeXryAsVXzlw5fmN7PrOaRAkX7DdHKX4pbESf0V0+B7p8e/h9FKG
zPQAp0b/RhlY2hf72Xxcl7JbUktEifZJWaBQlTohYzOmaRPNuIWGgz+ej9oY
M1T7nIdqd4suayBFcN33mHUAafP9UD/8aIsMS2D5mhycuSZwSg8jYibWJJeG
3vl9EV+tmVuRoXUBA8xv+6lbNjNVURkIrGN7p0C9PG8oqfD6QOGb/ZgFJb+b
l4IN1RIxwcLUSN3AXRcNSNal1f2ORsZBUOdoCn10K3gr/Ma6cbAMU8PwoGJN
qZMCnDsPBtssoF2Y0yiga6viuBk6u0BuY0/WC2aPNGrTyKv/T843H1OMtQB5
0uVkTJ84yyGsjpsJITCnbPQPAUizca6kwsqAURlmO7HGSCDlpAYpzSfYNQf4
bB91uY9Ko7R8E1WmFkfh6CdimqLVcGw2TgGgGLcV7N8+DpC+OD1bsLUfaRuU
PpLfXzHbQyq6G1DxhAdaxZ7iTCr2KJ7/7Kn0q5g1asX2t2kjYtcYjUEqzSI0
MCw4x8OJpj1PswjX/Gt04YoM7/+3eFgvLX7fJRRGJhZSEaiNVq/wyLtozo4v
zBk+EaLKeslrweoCdCWQ1UcpTc0gjVq7rHdWF6+6RhRf3VMjYArbKZ564LsH
ya1lETIB9gRLEL67nsxtI5R3FEANIi0wvHG/x0wTchumF+CgroxG1nwi+USe
UG7OIRKeNCryEgU8uke6F2IzDhqKBbYhqzsjN8VepIkWIrf5Z0cX6QXBR6db
uVnFmjk1xNeCfe8rCA95/4olL9Cn3TdKVyDX0Steh/mYK162wFvUrPAEKGX1
GiPicTbuXQA7LQdxNCKmdJvZ5kri+O3DxGAf1T/JInfFq5SXN1kat026oKI8
6P1UpAIcEfjSmtey+AmtWr7YSdKPSqsQfRRmqR31megYMioJ9adJZXYmNOYT
9zWtnsPljpSB7o6PHrTNf8HVn+IG/AddmlKbwffAktRa6dWMb0XB8Pld2ewl
Li/8SDPVTSSkiFOSUCYJp1CxNQPYvMn7mINCB1tG6YequxY9ir3yVG+IDOWP
9mlYUH7X/Xf331OUSlDiewo2gFeE5FuDfJOvtvH3l/nBlH2Zh5C7KD6DS4Bk
x8A6mwzRQKD22YyVWzgg8Kf6LUuP+arkUYH+2L2xpj4OwYkzVk/37j8Esq0s
zs0NVTTcIxx5jmPMU6kma11N+0ya6PeoqkXXIp2F/CPfmcs/rtej7aLXkYma
dXsyyndKk82uhrjTOfkLxYwd+7H8zoPaXe7j9uH3Lmoh5cf3QsCCJAEKb3+Q
nmjMbnpxZ+9MCxuB7HHvpO2vBPLwbnjVEm8UCz/brI4GGf7qUcbwLy9Ty6Du
aYL5bRXVaGCNXAgsYOt6t5dBHBEk5RMLA/ixIrZN3mttPGHWNjFLJwatGVO5
LpSsI2oeyk1Yx9FbGTVY+FJjBkZrXZHTzzkwuXZZWRW1+wflZLd04Kv1NNG5
8Am45ZYIt6IBbPYafhkF/8uvjLJkvmrmeYmeOU0Ui1LxCXWhtzfEIfRTg68z
Jacj/uEXiDiCIFhcO8G72fNl+g7b4BAMxeW7uVDiXowH5027Mq0Z1loGZ+Zg
0ePYC8jpJB/0h541d2zLfUGzW3lpvIYMOs9OCKA+If2E5SciNdlDny59TaEh
p8y8X2/ealfwpjrhEe3C6ksJLvNX7nzYDfG14GzoBQjXuSmj/s1BhFpj4v8z
rLUgbNwWjv8NgUi6dgh0S3Kay2e9bbOoVI9iLErwqAwyqmqpu3W8fkb/D0ct
GsIa5fs38neRRrs8Xzl58aCWXX+bRKyn7eRWeHZk0zp1e5hqpLLss805YD0x
FPn1bs19ppW0NzHGJYCB91AnHCGKFj0hanrol244D1WdwGCjJIFdpFfPzEhT
ot9Jq4svaxg9gw99aYrrZz1Y0o26QHT4ehNgkzPvyvWOfN2h74kvJhJ0fvqv
yDKxwdCv2FbL7X8hfKBNmpJwXLSemcaDWmu3dBTst6MNVGVjQsaq1rl0yriE
EkeNZv4+20H9lRqzky6FkBzgEhVVDSJJBaIPRUpOOC+6wXtEP56FdMQZ+G2e
O+BibBjj8vm6V+DV77tt3ztNBf6JQfE6LkSmpzKb7AgodXifJflyzEWH3hyP
1u7PQ+7NuFqTRK3+cKnf0TlwI8wtOwvXFM/OtWv1+mJkfQG4qfxCM3RH6MG6
ooLgOZ/qoa6jUBhC2F4VEJzXsXdbdabaxMcWOJJpLIGIL9jn9/Poztqei9lR
aN/MtmTWE7jGWCbn8BlGFjdZut6qh3J2JL7Pn4y60Am1AjYvci+KFOmT1mNf
gJUgluR5Qp3/ekysQIGd7pPcJm4UWZdNrChZFKH+Mgfm9wwyKeOHvyuO+Tsp
XZ7UahmQDGEpHHbEMGBQ/zy+fGsLvfv0uDpSkq7s9vRGi7umFUq2qMiiFptf
rHwWMfNKRGvt7nF0rHlD5V09NX5IcXrnFv65YJ2U0f/29XTxsfNHE8HI4u6f
1n7YfATEhNJFZMp3HJKLBlUUdhSndIKfwLw2xACk9LW38CsLQMIbFcIvU66Y
L2LXhTI0ZxYP7jxY2sNRO8PJWDCrWcIDLg6pIKvqbSmSC9CSsaq+xtjQcTDg
VGQrfCoGi6dyrJyg08qDF4sCH1IcgiVkZQiH1aNmq8WZ3SGHe6aIcP0GIhfw
EocpXR6iJ7tcflaEh5stEi0GFPotCJSEMtgdfWYZS6nUvyGiSTeD5KpHKz+q
D10egKjCf28Sppbcp2WYYR+GHFKNhTgG78cNYawlO6KnLKWiaJIEeJLVACre
0q/dAh1aGjWObSKKFJdsHov2M9/AdnIB8G48cKKt+Q/R+tc92P1ybn+12wxR
2v97UlGodPKZ5h3J9QKDjZ1EnVKn1kCqLo0hedlL6g5svmDrFIleNAYKgLFL
dygWz9p+KBtH4eGBtWEbRmV1Mu156PBU0XOr5SBzkdiJinlPUmvHMcNEzijc
it7RXFJPu/UQUBdZ0dMSJj+OZqb97NkQDXH3r5zyyNBeHZzv2ITMLjH03vL+
XcOBRR35AwhljXPbIL/bfPG68Jp5HxyDGJhbK1+UO3D9i9vz7Ojz3tiI7T3J
ql4wGpWP0ODubDd669rssWEPvjCcWE25SEyVz98algWQ22vF5T4x7+EBKWpy
M5N7ZP0p6gXcdGcjQxLWzSnPy4hNWXW20xa/XJf7o1dBCxULWjow6nWiR/1L
5mzPZz2Uo9uFRE5zk/z30oyXqAzEv9AkdDyt7p6b8weBevtSMaERIID1zbCO
N+WnlHYeizi/EJi1xzth5BqExj+7ETxsGhlYr5IBlsVYvvNmtAhTLfrSfTd7
OU810AqndDittxO4B1NvJgo+gq6sdZpv9lgQwEz+kXqhcwy8y+4B1swR7mgH
8kDnNfwCxdZXnP89rlDe5KcLo6NHcuUfI8vJAFEHF9/GSqfLK09TNrAhrKoR
63gxlkYHdmee3kcgNcETnYp9QbBq7U82eZJ5bRcs8oi+cZhSqZl/OQOvIkJQ
R3RVUf79LSpjaC5GAaKF2CaaRzZlXQeRo1u7uix5XqZmx5I9uLfddJHztZA0
PrZOA8EKC++1JP9b+gCvJQ1XZr81rPeG62xBC1YYA+8lMDhBx3906YwvV15N
iWvuplMemn23BtiHRA9pELwXzR0QEq1axTH8sBDSJ4OXbm46BCVjBPnVPZAI
wBdKvDFJnp10nFa0qOisx3s49h6JC+7fHVVqp3Tew/yn4EAWcdxNTDVANdOk
BiHcUPT0uL6BsvcblOUQrx07FGm3Mgnr92Vx6oCGnqUItUFjUnHMSFiSXCLb
a3vwuJU/gUJBrqJ1EJx9AnG1PYQMGsPDbghE28mIzCydmCZDs3ykn0iwvRqm
TJmGvw3Dei4rYqlLMAhnHBpRjIf/G0Dn0OSivjqdjJf4b3UsZ3wAdAsNsG7K
YfH5bBTasrGAR2kXbMMenDJBN7czdREq62URbfcY5H4HU3sIBf7j5SgAv78G
WONQYKuic9PkB5Y3l4nO39J0UwtSIsXiGvRuT6gV6AZvbwLvC1VOXGJlhCBd
Mj0smAtpgGA8UgVT1FZeFTEoK+olL5Ns3ELdFsmTwPD9/DIoHUtaycm9qana
fA5JFryJBVlG8KeKRKZ44Yvbdv0IPrmZ5pttQTkjS9gJ6xevG0birSvkg5AU
/6xh/jehPFeUYLvzB6oYOKiSXbyZx9aH2UJNT+fU79hX25MaRq0FiAnyjHZ9
6CJopGN70QUnTNsfUqq5oHFSL9sWmav7rfvWVKUWToeHNghsyIkjYU+Puctu
TGj8BHv8B83yqPhzxPitMv1PO8sZBgxywBUUO5VyGy/8Yayyh8puoFOkPCgF
FsFsL8ExIu374mFBILYdLVjCrhRKu8DZiTKdu8bAXL2jj19lH1EfdOOvh/WI
OVzR11jpl8DJxaZC3tfKc6Semr6aWyh3nnShO2wOtCt6SJacV2y/auGa7gjD
LYIw93kYoEQsMtw1eaXWWIBebUWKd2QP489uaLegspHYthIC57Gy838BGtX8
9WyfqtlrTcL7mql7+mVLyn/miBC5z8sWWf/yfGi4fOekhX19+dls08+CLmRE
9DHg88rDh8/a0a4K60oHvJX0fsDIIfWE3fJUPle/otx2vYOLBwWGmyOTbv69
KlLaww4XXVeQKZ4gx5d0Py5/Xd/RmD3XflD6ebpqIrmBxXCPoxxEcK+Mqgnc
1ROvgMGIeaekoyzu6lTH1jKto+4xUy64qey5Bxuvyx1d6NteITR+bwRtjgnb
X1Qw23DDteJADHxARxogstiIxVJ+4ry2KO5Q8Tx/4g7q9u23CnhVXO7fUqyl
GuINIC8m+uz9WWEAXhZAz/MX6EJlkehHGib448Cl0m2Z/RutsgeEAAPfFx3o
LXI5d8d/+Dqxp2Eln6t1GOYQT8HPOBMZqxFPgVsyOEYPtiohMD5F6/GyGZ+N
aeyRHKg1yPew0LUpbcRpRWWxoroYMqXTSM+pt4MIG/Y30HmCcjTjjE3Iawca
72by2RTpRgJp26wBnl3UvOas6kZfBjIU8EmL5EroLXuJPyMtmnHNbtbeCBxy
rEkkTDn+Bki6d9OE5/DkxwxLC4v8YVH8IFZHlZNVvl3o6BYzFAW8NsGgVQB0
n/qwOXj4ZWyhAD3C995FpreMgiA52UbsrjvopigRz/vZ/pXnWRLIBj/paLk4
6Xgq3xuSiTmBDHM0MG1J1NGvcS5d33lHq/nZKSBjlsIpgcmsef6fFAamvTUd
i8HJEQbk0Jag0e4b94C9IUTQtwfxCxQQmzhGl0GLz4xbzy7Gq0dojdHeTclB
e5So3upUAjDm6r1briaGSJUuzN76mGZSu0Ta5Iy89x/sh21vl82TNwRQwQIw
ENcz4vBrhD9qyMjHdX+G3cmzaX4/+EWBtcWn9wN4sHdDU0hcCeUtNUV74a/e
KW9bxE57+Oiv0wQC2GA+EI2GewS2SAo1KN1wNX8wIPMZq6fqRqDs6Sh8ApA1
mrXk8kL4W0UUnQEJ1tf4IcBKdkVw5+kk0bZf1wu9S0sEV/lNAalH6jVZvM0o
zQnuCnzbOjRvK5H5gSamHPVCYFmhMQlnw+VCIM9qUEsIYg3YCwRd+ZPkHal6
Chr+LKxJYzMwx/gghwePXCjZ8BwPfDB7hMT0Qn3DKweMev6wpuyarA0u2xcd
/x/YPKIZWIeWcZkf186vRBD3tDIpYrAaLvCATjvOBIj5ZWkZ1O750dWcTcAt
79bJZYS7eRDuSXrsKQ6B4ZHyR5IQVinuhGJim7t0sE9LQTXhpYzELfal0g5O
Lr/U/qo1la5h6sVznZ1S4/hyo7RlZFuW0KyV2lv0JX82+0hOiIp8M2bfUyyy
r7PqtvJ5JqqZSE3mW6UKfLVweyVdIX9awQCu09N0k8FV7ChRjteBENqHbh7/
M3hjQyckJovwgS1M4pBuBuDRDbBvqlKIXqjnctqNYBY532YZDROl4jXAtHYq
6XxJcYxc13SkJqZh8KJKUF77OWT2FxZynAIF2P2LGUyuKB4UC2sZdfkLSTE1
yZg8uZjyXBgzAoMv71PViw7AFGnWPWWGwxpQLkoU58BFEH90lnYiU/ppfhr0
KnR/+c9bwGUIwI951FLJ1eOKHp3kbkE6co5N81BfH50JvdKjbf7z9msCyib5
h5khg5Jv3VTrEdji/1MuHW0qDSDv0/WGOnglywABMpH5CN5k4mj+fxIJUbpy
eGvj4QPjN2atvta8cSZgR4hauFlOTKljBP4cJLs9X364+uF+SOLi0fq847zb
dSd+6cXGVyAyQ1SwSiKvoGwZ8P8Lfd/IaaWLDl5u8oUD1U+zPGSFmczCDNix
ub/cDAPum1qvONTj4d3hsVuoRUFvMK8KjFL/Q7GmQDfPdsnhyapDbJ1birNC
Jv7eDTrNCxFXnobux7l55rdkkaEqMr/X5kKBDQFG9Vxj2JmNIUmrMwIJc0nJ
lt7MsOo2vIvOqBRdZsYUHN6cOKAowGwvri/U3Ao4avgVLjRK+56FYvqCk7Hq
S5c5VfGNgbaNrm4K3WzRBhH82WRAq+coE90NlpaEYElcNwfnT2T/HscEbcuR
0McIwAXwJxROzT/ttn1gIuax07NbNms8KceE8CzqpUeam1tXndl507GIW8nI
lMfRrxBiniHasDOgC6bCIgFRkDCxztsyXhQED3h7agzL4zsO/1UZIZpVxcPz
z1bpBCJT7pI/urZHL18FJykZBoF6rRBU2eWaVQNgYw5gykrUUOh0mf6EL6bb
xz2qDYC5sn4HRiS9yDJq4tqlSrHgAZGwsSeNMG/aYt0cV6Z8OosWeyN4yXpa
wfCb9T3hxH1H5jOkqXoWdXEsnMPNOWWBopFjF+XUY5h8EJp3SraSq+ODS1AO
IHRaiV337i6ZRt72qdOlhBQi8dcLUcWcJUqQRv7TV7vhVXAbEWUmTH8nkWXj
kIIKLfL0IL3jMVFkE6ap80tNORmONJEkBOq7sZebJjl0WRspdOkSz/SBD5rz
945NYAa9IQGxNxQ407QTeWrRDrMzS9yOIIlovll0pYQvevzxaUnNoQ7qi3kQ
VGE4pn/iMnwq/loveoeyeYwLvpF2g5tAWLfZcOV/ri8Bmgs8G/4G2PqbUbx0
x5A/PQSY6RGVemPkhNvamwArEVASkCufZ0W6NvJusJYDT3d04VLuNUJwi7zb
SzwzZkl6SFz8sinKv/PmT3SsC8tkFAezi4ziDbE5LnvB10UtIjSELaEOvogG
67MZj4MqrJb/yLy3ZHWHO1xyaHSkrbHCzJnLlc/7CEqYO1LKIwnZTT7FueYm
frbWgSIBNRg0S6RXlbBx2pJUJiWdft54BKLeCC3R22uS6jDzXU66BvqNTrB5
noOzt1oxTA65/p8cN63bD52B8hKaAQpcoDvD6iffAKwiplRYdvJhaOkRos1a
O9FCioyRyips+fA657/5exanTQT0yGBVtqlLj69z7rNgXLWC3ha7NNwMnkF+
nIeRck/4/VpLRa7X01inTv6n/CmhtZD8SJj2nExZ1UX/siIaVkoz7w/Maspv
V8IIHApFz8Xw0CmRp92Em4CKgFcu2deDf/O3pZzicEfwWSlevmW5UQNgQMzg
b41MeywA3rnImArGp7uouzSLo1vwxdqf3hgcLwf3GiNj3qZmQyEsaYsBzznp
Zy23hwrsRoHpn4wZZpUlrObOon3Zj/Sf7nRtLvNaGHe3WEWoXZ6EUAJr4auO
XM2qGGv70XGnWWtx38WJhIE2EUSpWYFXPNKfBhEdfexosxG3c5XKZFd9qQZ8
2OYL2yzfIDtMBQnNDUifh3/4bBZhBHlHEn99m72x6SeCltzzTu99Q/yEL/AI
8I9OlTpn8+O0AnTHFC0Nr6VfqVztMGD1duJXfn/Ue3dAP76hamzvTz4s73Hv
w+UETWwgeqdFwCuaiKzdVhYEAdkEXtqdTVUMSFmks5oyCvXs7GN3BSCHn9ve
gb1NBOYdcOHDYD2BtveVtzNoTUPEiAIEAFLb4XiTTpDIWGtesatQrRXblj8y
rsgDYqvrJt7thMrJep3kZ2d5n0GiKN8HcgK/W5bzT3CmQ738h9olcmk8bBH/
g5i+xTwPkHXCPRdphHsfUhjS3jQYr8i8VF/VemgDPE9fA5+X9nT74qwG3T56
a7dKZyL92rZBQx9e22YOWkdqet3gFqtQl1uYXQOcSmAE90nxE9urT/1vN1QM
UPDhnacZ8vbRvTWBwyKd+YMGELlI6LPmdhMUwt4TPoFOjfJuDtwGIQP3qMlI
ItYEjg1iGoQ33SAzxJLIe8tE96tTnfwcR8U9CI3LWjLVNneWr5JYOr7AMCLo
dSzKSzZKEPmyC9wTDwRyarySlNQ/aGxtBBTUVDyuc0+vvPaGb5Ka333J9mHV
dsNDZg8z+9aDTMGsVmXyNOufzJHnLbSPaIoH7sd8LC2ZVqXd2ApSNvb/WnTS
ZIN/Gt0pIB7KEcmBZfkldmV5tmwTkgAxYhLZTkD5DSx9s3JkA8v9ulZV3Xux
Akm07dq/5ebHvR24lmzwG4AwYhS8T88P7BHQzS9mGH05R9+DBh5XY4ECkWQE
BDjKa8g/bcjyhchvSHizV5BYyxwsUL58uTPHhimSdlb+erPZQv5YjfTGPBGZ
ZBsbJGoYsPt15Df5p3x/vaH7/l6xwaOVjuYOP5Ot3M5Wtf/YFfPIKFORnNwv
tRdYCKYwixVqTlsANJDzUw1u4k5D2WAglH9wzhDCj/MC6mxP4wzdOcYFvtNF
g77+wUMhLvBmrmO+lcX8P4OM+Mk9jxxrDKAzhxSsa6eOTNsh8J/2WJPxij7P
S0P5IDu0shmXw7oLqG3ExmbcK96lKUWqDLJIhV3wI8JFB0v5TKELIB7YBDND
TqzHVlWZUiu2QlVZTgQEeZvSDkIDl7HVmm2AQV7qo8IPmLgeyumNfH/20AND
OE/aPRUb6rbEZTlSJtWKDnw1SpPQd3xF8FMcw3W7xQC2o7IFPQTS/u8p2+X3
EBNGgNqVym4g961kTwqKUwXpUXKWiduHPRwbxuuQ4F6+xWzZB2vzm9Ogvi2R
ws0SvufCDphKXjTu54VpYNcxbz80x6UxXyUeebqRUwae/vkKVAxhrmZ8tV3J
4ErFQVMYuixPV6AT4NkX70Lu7fGrhdYVXsNR9OjxtcMNqYz3SPxfuoBKAMjF
Yj7X4N3Ibr2EIpoALlYUfcPXeiHfl/MkbKrKtujdjGupMr+iGbfZeE9RjS3c
paEBTOHUTGvwyy60vx44CiOP9YshLJuMEWou0LwM7v/KBO6q8utEbTiuF1zj
tgjFZqQoF8KUGzTTxZZY23ucxnxJgWKmwofDK8JAX1TFABS2j3CZDcZ5lzfe
35d+LK3TWo+j7sgLi0+lRpYwT+dTHCJYjNyBastT/Cls01OfEdvdLtSQKJ5P
2ek6YEP6YlDDeF6KfRPs0s5l1iHWopHfsD2RAzGaQF1T6I7TpVml0by0Drm1
obSMUyaXGVL72MoB78X88Of3IqM8bzQYIk/505NhM+Tm6xcsPjc+Vp2XI30C
nmRVQ3751hQEv98aI+QW0hyxX9GJ/kbwZuU0E28aAjLa6iPE5rIM4x9Pr/FH
/THV5vpatx4l/r/JZKkWy70/H5nvv/N2+SYs7jvc1OW0w17JfsiTvWIcYjkk
DqTT70+EqlwYVVa9WgwlmcXRAx4T0PAKMqbn9mzX3qIW0xfQ+HWRagAhxf1E
dpumpnStsvYZa21AddX1Lto09g1BNODAIfxALoKvP3AoMRSX5RghE+KIUHte
dK/6iDz0yi/pTcGmDGZyc3njXqp8W3l+4H49augrx5+G29FT8B5dKgmXFV+G
JJtlulHUG5F6S6fgxlDwqi6HNsefpFOPr71uzylRamqCDW6HpbUDDcxDADDy
i8tLpe2QWchuwa6ZSDQKIOgrmm1cY3oMJofZv4gL5+hQjk4hLG/fmFChPUqQ
p+jSZNnH4pgm6+caCwP0bLy3JPfzECWo1qed+Oxze1asZ0rHP2pRsE9r3t8I
UkFLG7feCcHIjke0JnFCXDd6XzBUIU0k3iDVGnkzvvBGsJ5f1mGv1onhdOla
/pqasnVxGuNLn47vZt97kyhJwZTTTECRpS3Xi4aWFKFdeO+nFyuJVxOAPOPQ
0Hth2LQzIPLEvM+7+4999GRm6TcQtFPCFycMKgk7cfazZk+tj1z41LlvZRR2
X6eJrzO9rMNs3JxDBiVEQCFAtYwf+yHearjfvFEvFIbEV15d1Q00p616qSnX
tcI3uO80vr/d4oT2LbQKoTL1koEtIlD7bLsmyUt83iBnH9tBGsBHpXMKTYwQ
vM3Naw+lpZ+KESYX+n9o0lx3atEmgEq/wQAekBA1ROubNWBHmQBI+Kb/3sJT
UHrzU1/bjszh+WELhVBmb2Rj2s3OuGYGpTMlJ8H3tp9DO1hALuv/1blFbEk4
LfNoCpFWMvjce7dYPJgig6Dq68HF+2CSgrlBJrjGUEknDlb4MqYbdv4uEDeS
VXrhJ/YoYXiaLL53Qj6Eig54yIW2V9+JhbXFiVLLweE651R/5fbo5IVom+JV
A5WLzyd9gTjakECKRz4Gf5FNFsybPhIeCX6UYCSSllSWhbg+ddCtEw+psOpl
+hxUKxHK1UmjyRCyJ2wPOIepnEGRYeZTA8YNX2TxTtpgWMD6843yfyiaBqk4
19XA3vT013mIGUOWvEdvS+niF3YiJD4RWDPdpd9uGOPy+FsXPRf0pS976B0j
F7e/vvSAYEZmSGc7WVVIf8CXAJJukg/ftRnPCIOmEJXGNyPlqYsyUljHfvx3
+lrzSLRBgCcpWq+bhIDB4VSBxx6V5ZUTaRrCANiHLda0nL1wmMHteZBdPARj
rqnPzZrW0w9VL5XXxZZ4cHGXaGhGN017sOxbXhC8ZHd/+6yrdRMILWbwPsMj
GDWCKYN51aUfg2hlSBL+xJJHx3PWLpHwZxqCjD1byLALEb1bVzyip/HLUUjy
VHObD/uLrY9yMtLHWINzpRRtoeqcfVuHsTz98ut7ryLbpL5u5/TKK3zx+9in
huKmOUyWVMIZ8TRHwIz9DPHwJ0XEAged7z3JZ3DfTwURQ1wkVdyuLHHNZvi5
n895CtIew1XwHF5ogwvo2vBLrKhf7ioPjgVOEkg8y7fa36ZdJV9pWiAlSTds
IQesE7U5PKVR1nWdrIDqYEzalFMyM/bbgLKs1z7qiK9pRhEgaVDxPzEUyDBu
rtTQT5ZE9dUcivDkjz83rnpAQmnCQEa1kuIwO74i28ifNGNzM38LmTzytgH/
mB0HSaaOUA4uU2ecWpzjBNYf2a+aoQKaInPZBMqLXI863P4C5zhunJ2IEXWk
owhrGDvXFq1/pOUdJYndkFghI+occYhuLx97DaYaRt9DE9DbOOiogx/+kggI
Lrf0QJWVMwAy02wsWkXbKxyeRbh6WVkgvtkyH0T9riqLvtilfAb85HXsKmyO
CTF1oFe+P1gCpOP02CAPl3No759zyMI65lutFv7fhEbdb7CS++wJiXsYwgzi
mRdooRDf36Q4hgRI0d99ERuE18gzl9mgMy9V+C3+yS/gq2pl7ohESk5grVZo
2g05fYAfABCc3LPzFD2Xxb2IRW8G9gZD/3HK9W+16W7/slJCnpiWJVGtNON0
Yf6wni2YMF14MnAKyNazBXf3FqNA9kmnMf2Bj8yRx0Ev3toFFUAC1iGPyDZU
bJn2aiDycoL3tazC+RZQtBCYeLc/omly2NU18w1c/oAggcGiQ75qNzuz9IlE
upEQAum3GJkckxFCoHjzjRf6uiP7LaojYFxbAu8c/I7zRkX8UYt6rLfiYwWh
p+u3oxBCIOuy50pTbqjRuxkblFJL7EgyUw7Wxe63a4pirJrnzuC1ijYJUZ7R
uEbM4GLlDF9P6fLzt4yHef8+Tmw/Gawo3pQSmaWkg8e1DzWIuKSFc9ijgVR1
klk+BT021zHJG9hRvqyj92i/XnVbOI/yU23bx5QGmZmP20EpArxE0B0EA9A5
ojNZBHQkE/etAvQkzDUD9u27lD5pMQwRZQf7Y0O0Xibc0qlT7YP0dN87/0NM
wuqhqBJqPZx8NLoq6gq6L1U9p2Ky3Inu81gfrLfeza/1gfc2Kpw0R36FjGVU
OIrhueBSPK4Vgp7DSqQG5FtVEH8fU4om39zqvKRqEqeh2tLvkaUFYgtV6H1l
5eEdndVYPSaVa9Buwm1Jig55b8ykkSbLu2aHcLAecAP5cbjm8Dytr9sO1h1E
vF81CdSzJ6rrbnDIfRfPkzCw5D4BHxrGRpvYjuxNqdNeyESiFWDqjkEOnup+
1zuy/Sa6NPMb99kq9urVGFI1uItd8EoE1YJxUOzMQnwwmgj4lI4/LZChyqq1
iCB4W1QinB2N4E1BROSLKpsBzaOYpgQhtcW4nxzVmmMCk4637aWj7Ylpwqbh
wKsQZnd9rYLKVfDYIrIsKe6yIRR1CoWkEr0kfLHxr+u1Wo5B3EZ878uoP0qO
YSGyTGWktjKxe6ODRYXnwXYdsM0Kpt+dVa8V1qpY8JE3yHnefC2K5Jx9oDtQ
oSr3005Z+Lh3UlmurTBPtxp3LnUrY6Kg/RNXTt8fP9dPTLAxt12SHBqYADdf
CZzOoEEIa3kgVD2KMWeaGrUxmPif8bSHXf/hpqx3+VHxZrw3KksNRr66AMmR
K9oAZonuSZcYVctNVatrGgyQ4KJdsB6+5FEMVhV8c2eAWpv3ndbpXklS3Zqs
c41BOoi2gLqwdXm45ZCjh1GqPhgbbc00oTX3YFEZFXPT/YnYocTp7S0AexPQ
kGCFPPT0WfslL/XZlEE/lTPn3qKEVDKHSMgvKvOcmBDr3uLmVvZ/BFkjhzwN
kQ0d5p/IY0RhkawsqcgRfWd+tMgwV/Xj+2Xdvi2usYbewCoHBl3bSNXmSSI1
hctjvC/ft8UvlexaNJxPMmA5u9RDqJ9Nc06TCuTGuQflo498j8v4OEmwqrN1
ltFE8SnXeKBBlFEAz85OUSM6TxgEAGfvGIFFrwnMAVVGMsryZ2hv281++Bac
81gjT2/1IlJ3qwnPdOpgyLeGW31MwxG7d+0gcGJNpfBo7+H/Tg2IYuINX08R
zqn8mwV0q6uKxsf5Wyf6AU+YCG7dz/PuYoXJNOU8TjbtvP+pOUMt8jfzN+kj
5Efnphv4TVski1tRu2hG25E5J+8B1F6efOZpmN1ySJRZxLmAqP7LxPKwOXhD
BLNZ88dWgBoz4JKwKJOMP/4vIfm326YNBo8uYjHviwLvyDjFf5kJRvXPGWcU
NRKOU+qwH0TN5zBXgYI9lCwd+j4+3bPHJiRcTJjoqXWu4TYh40zvblJYq7bv
7LiSknjQoXZ59+68jPht3pcqyZVlCxjV+lmFtmgrDjks0VEq3jpwke7Nbz2u
VeGGaIKo4npO9eeZz05s6RAZI+MmiI6ailfj+fPtGMhd0SuLhO9hCF2ZSURM
8YGLWJxgw040ZpmS02+3Mhf+z3Ie7bEnUAHdtcx96Ll8aoMukAISz15MPKWt
vOSrhmydo5zv6DkSp5HT9KUK6GUWN0EvVHJt2w3FfECkUueojcRtQN6/P5Dz
+Lt5Rc95S50nKlTa4VlLM6sMPBvT8NfjvnqOIGtQahvGzJ9nMVgIvxzLFwg3
BzaybzYhcxMUeAw8r/rlXmL275jV4x+N+tmCdCu5jW0VPu82NjuchK13L2Gz
dPTAHEdp4Wxdj64NAkxoUsu5dUlzp2Jfbjf1EdqiM+MTE/M3r7tWlPKRC3gT
sb5qg/Aoq0g0m9p7KC/Rip2KopS4k2k+5AjYPnP4SSEEFkx093fSez8tkg6E
NUqhB1QxBY1pXXUXJVwA39/LUtVxz85ys5IhKb+azcrWiYOzM2YrNucmS4Nz
9rn5CCWktqfEtsqC93/W3KSrsmMeWQZIc2q8IotO0oDY+xIYMui2OvXKgbcl
gNMVfxOEgEoxT7U0RXXfZiXRMM+FcOhz1cj05oCMfN7NG9pGTOS/3uVWz06j
tVpHwkPtsvRQNsE6EKn8mdqU5bO5WuH0opjYL7bCsBQN+d2mTd/fYtfXeQ6/
KCM7yL3TsfZzYb+RMLwdybESw+qmAV2TbNuc78iAdujkyIjRJAUZddZXGfOv
2Vo23qufGp6DjvDQRUyHg2r6Yyms9SLynnMW+qKMtOgYJqX/T75zPYiWunes
EYa6gbM9z0wQB88gYQrqGpVKUIQh/76eaPdemosTVals6416yIFz47kykqQY
JJxz25Nc5LjPJ+HjHgvm+i46cdZ7LONFmSdL+FABU1WfCA01QXYJL0yPnrng
Ru611y16iHOlJOEqottoOZjz0yYI/wCx3cgab/REqNZOwlqcuJyqI/TOwUZj
c10zcWNDhA1APc9JnRskGu1DEXoazahVjRTk/kGTSBsmrpD/yzibdwmhnZge
crjZVyDgQSAQbR+QMGoH1a08IqZ40oxLbNvjPmJfmrYd+4RtU94nLUjHMHgb
eoZh1nI6F3HFZEmtCmefUE+f0qu7rVPlvT4uTWY5quqwHUjngTUr8qN6nQG4
na6uxWFNDWZV277D8OsXui21V2i4JFc0inOTCPE4ERl6Sw82xb3Qhwh4ziD+
o3kYXUZV1EtQHeSx1k/CgNiSGJ5BReK0XJNieX5SXYyXgOeMV7IcgtSSxlYM
tH1VSbJtaI4J1K+O75y7A5TpZ1S/ZL7JWZg+y9OXPIWhTb8RYOZnUAfTa0HD
WMmZ4HS6uqRixgzQ+KhGfw8Bu3wpGiWOpQWnE9uNGhVE2p1wlnQGa5jTT5zs
ZjoFvWVZR+9DhhX2c8QG4zw8EPIB+rjrTXjwjWB2TZCYR/nCOq1jDjGPcYy6
YY5hkAx8wf4f9tAIU3kkqK8tk331ZuyjtMOET8S2DCRv8kUfB/NhY5bWkxPE
09c2SXOcogOvYJawg/4Uc031qLs+qZO9O7F1Q/UV/sSgNuOy2+wLqZ8ONr1I
YGAT7LtVbVfHLVuV04RQjSeT2wt/sBqYJbhWZIsBjRL7SuRBPAvR6AzJ7uEk
BDu18YjBpK5tmV7UqESD0dXBcQMznO4zs7SJrGZJukRXNdD0ViwSDjBVXUHF
56udHxZjEniWJuXNCBPdJ6bjtycZ8o1fxJc5exZKSuy42cjN7FETsv/KPTyp
R9FSglp7EXhHwv1SgaeYyECoVeBGIKFfVqjdYfWWfRB7Jclgl76YyuvbODav
fkwuyEb5AitG5Rk29fk36ocv8Fs+RQVcV4fJaSf1XrKsaRiRAfihzQaJeMrQ
02GXiq7gUR7IB2OGPU4UNp/d4Ry9k9i1DpkF64xkvLCLgIAnR0KaLaE466U6
SjMVEpfMR4qBvDYwBC3GN9vof3cr/bJwX8Z4wLDq3P5vZxlifCsf6ZEiVxJE
N1Q5f3Jg55oJrNWPM4UW+TV6zgDJQm99Wkg0nZn7L9mLc7cRel35moiWckBw
PvTYHZ5zbJDSmbltbNraPKFxelw3iWhzy8ZnNxyPgfsNTNEqcPgXOVmLJ+4u
Tu8PMoixGIHKZz02BAMdb1f+8uIF3bpaXFuJlsCyphvOgyhuS7J5bb0gjqoR
FG4kabnVBQrIRwHZzwoO16yWdO1pC85Ezv9fcgmvjqroMdViELT852GUiY2S
F2O9uhTZcN8AhY3gdr6sSA0tmz1nEXjzK+aQQ5E/0KjxgqR0qXM55fiYOBbP
JLLDKseNrgciSbV8lBGy/iBm/p1MLcs1wmg81/u3z5mpMg2DAxbaFApitPzh
D3INXvQLfCK3SLhFTMV+E71Ruz2mNi/AlBm0G3I3+MJWIj/2/IrtLZvhGCYP
ZvKNyosKmIQ9apGAwME46Ah0LwsF9ccCsdKJxWe3YElv3ASG5ANaU5GCsBni
+N+sGjtB5rDMvkheDXw6AA7qikHOUcPPAD5YTGCuuvDZbr+drfPys9t1HMeZ
hPVW3AaORRkBnft2iyFxj6CK5sSfObxDikJpwZ048Wp1ekjXX7hlhcH+Bk7s
VvRP7wY+TSKeg+jWiUtWP6X7oIsbLoDEGI5nPhTB1nw6xuyngpd9j1D/yrCt
jPjwMjr2X5Zp3GwD14OjJlL4e+Z1GrexA9MebWmPvF755v2OXhTO+Dbt2dgB
ca4AcEx8yOCfZNgQzDK05Sjgz0WSM7IMrCzt16yqK9qGWcKk7AxiTKyx6NYO
6fZdt0hQg/B/ojNKQPeweAD4gHOyrZMUMGhOItKFlSWGB34lu6h1Zn23EMhF
y8SVyUoBRCkUTBKVrBJllusnHNTopAUEUOzGJH+doKf8i7+/RZaIkTlBgdLt
AOBpGvqeGMlGBwJ4mYgfMzFqIR2peyGaIyBF3BgzWzHOOcrreO5xqiibn8no
00Z6H7sDWQ8PCREGLtWuqK7ofmOCoHxqC4AnCE+cO3he0wsoEOxwTV5gE6u/
D+C9bHOqDBamsBQDMXkjuk1ziTZm34iy0ldYDtR1lOjZ9Wz0r6O0AnSGuUXM
Lz4l6iedp49pOI65KYZmX1WQOiheZUS98O+rWHpEasPDdAd7Ms0F3tR4F+82
5ZcVptILqEuYZh/BHyPky668xLAmZU4GUcGpovUobjfpxXxSXeg9+Ku164ww
ABt4cx0+qA3uS9vASbvtMVTamXG+nYRLr5d4BXMUWI3ZqnY/YsmEo1bdScdl
eqat69L2rx0WUv+FVGBxsqY6+ZK0kwJLOjVU/ixDyVgfUwkiuRtbnePk8qkK
py/irdYfPoh+P5F036USmaaMHuXy6ALE3tXn7ryvY0/36+R52g2vaX63Xm3T
TjZsqu/t8Z5ybVdxv/VrVcko6AyZWQeNmmOXmOVGhhkZFuigDNqw60w8aNah
6CCB/QiCGPaRcbDuGH7Qn1wIHE+Are2TWEHhKPpMuGIBvpaWKgybZp89AXEk
T78yIcyP0uxANSDw4uGe/oXoPnqsSfqhrbN6a/BPtmoGnacxga+TQq4g1DQD
ZG+wVaefdHMR85Bx9VAzWXjOzwsHMnjmNWXak8l1l8XnUWlRovExX5Nla3Iy
/VHdS3SsDzTqwhoNxagUJjKOCMZQTuTsATnvtdf/oJFiZ9i4dD293IsRFSF2
rMvS5KytKGQP3HfAf7Zu6TVloFgOlLlO3qPSyc3m9SOUVB9xQD1BGbeWcHG0
FksU3Kv0JKsyMB881IksUpcm35uLCGQscstcySbBkwBzSJohYAAOGcEKlm2G
02DSX5qWdqxBXcUlPo3y2fVzVOghToRcuoL/eKWeEDzEwWCOe//Iw12IR+1X
iSEYuyWSE/ZWc3r5z/iIeO5xHPEcxvp6Iuu262vZZeqczxbmRYQhnn4I4MNc
t46gjx2KK+sLdyZ/WFi6i9PEq5WlVDh3O5oW5zAUCDAJ6TnmLjyRZcMO+Od/
p9G01SAswsmL8TgTIjZsV9VXS8x1mruTsnKnYAZm5Ss7dTHGaP5CIbOT0jo1
EXu1w1KFlmEICtW/0uxmE3ZOc/tUGprg32OoLDt+cIcjuNqz+dC50VfcygbR
rU8Ij6ZRzNEyovHkpgfKIlJjWbS2ptUv8x8mc/IuRyoYlLzsZ8o61xp/M21c
jc2kbUxZ2tFTQHVpl1k4ml9HMv8GZZirgM9jyeUMEUcwDHM0ddEMojJgIWgv
e6ihMigicCh/KHOJf+apphZz2IHG68XJyMRJc4KE4RzeOpKajjLMxX5PuKbG
g+Yh1L5ObvZsSRJhUbxDzSxCAzjZnGAALajmMELl7fiYIGYZJXIPQKCUlrTd
5R2sw4a7snbLRZT1cjD0ei5eSDE+ENg+Ese9srgwQUwFCs2ny/hiHJLTDO5E
FhmlZij1DFMJQsaXrrU6sCu/VMJ+4tqIMtN+YzR3zA6sE254wFUmUM0ZTj7h
cvYpk+ueb/bgtexzdvXLQHZyjBi5XVwFW7zRHTxfeeMdQrz1A1/PtHiATFc0
qyP5oGBCtpWt37jLvQ6yNFeXgQDjwQ/sks1nlR14BNRhq2YQ/UERyEMESpRb
ep09yzm+X4hUqTV2TVdOySLK+bgaL3U/SLkDTh4CBAXS92IcKZSNSVeDsr0u
QyygjzIjEXoR7q77cmcdIG2AjWqTzmqdkoeEP+wTQqs7TKqjurEJksyeR7xc
HZE6oAz6cFuAXutA87zLkrIhkHU8AzCEQriPfQN3RJx/WPrv8E/ySlBWJxUP
6czuKGCOcj/M5qITNPDa+Vs2XTwBpFL+AN1y5iC6mLoO04yMaaPfn/Sd7JBO
D78G8yAkXlZLF7Aa3szMeo2EHYTzZKAnjS75On1hC6znlKbPBl0PAKphBx7F
Q6p+DpTjlWir++qeiV2FXpW9Du3xQ1FtZOb25flcpIjkKzqZmZftG224aRvb
NoyNWmUXu75gykLfCpbBafpKNHe7XYM+S0+xJPbYhLyygG24hqcCXzBhKwYN
jgj9EtOtrkvz2ktKiJFCzlVtf6H/wAZ4N6pYKD0ypgs6zax6PE43digQWoIJ
YWlGxpLfPVMvz2sP1+rmrAgrwWwDNz40R09leyfkJdbAGvjZ0lvt5g5UBcEz
ELL+YwQjEzaFrX/anVKtoKwBUkWlJQghAVAMv/tzstSFAm3uiz3BHgR9sHhb
8Am5FgolGheu1C0176aScPKTdaPsvF6grcSoh3cP+UfXd6xWxI24AQgBVZAv
cwbnAzYecpRy0OElFTPQXfybkTWgxNfvk0C1bI9p8NzmvNcb15j8bNk2sRps
eDfuCxNEWhTas9m5jAnUx5WE8oVrfLly1xH5J/ZBZrVcCQst95lwKHVBy48L
21t2ODVV+inZNKvhEXmKiASX/tWSi5bIEzlGfojR8nGrCHquSXjaIjquteH3
juOT13W9XwTrOpzheQWY1JO5b2egA0E64HZLOfkvM2+7cjDU8RjsyG+kfFcR
DY/mWjZeriX5rqtuMZzTNwrod8gARO34Dp558RGKi5vv/tcw5lidyBRjTkTW
KmGQk9Z99sF/BkNVU13Y2q2CYwDwNKLQkBd3JLiAiTEFROIWKR4oR3P57JHZ
H4/gDq7dvkzAaT2hpqX7m83Yb7fogWGLRzvJ7D/1F7BJjDJDZRtzOw6HCY3g
7Ukx15RVjfUGWTCHgLkL21ic1sjezBj2FaoI+Qx09CGc6LlwpP9j3o5A94by
KOID0ANAtTpNZmRSQ72zQKuDLHm06E73lVPNaNbhzUfS+NnFQEM32lrkDmrP
IKverbKdV/jhaEXpdTDISVsKFsiLkh0ZdOohe/66/GPCzoxNMqdSAwX0eMae
F82VX/XU+32sWZ3SyTOrEQZLiQkSOw+Clj0r+F2wvbXggdR9QcjobYQwx+R4
TwbxGKan7F2CYMqHH202P/GS4TXAemywUFqyRDmnuNCJcThcBi5FrXYrU+Og
/zWLStrdLcbtDsAz72PiuTPANywGzOtvYnyF4SoJjmb3xfUqfkiemVKDKA3k
j/4wSh5zGnSWoHPwHWrKwpDU6FFTRd0H/D46jjTAt/13TzZD3ssH3knpA51E
wZQUr4zoELpsEr2FCawKDTCTgQuXddUeN2kge3a/wN7DUuHIe4OHXdWjIoXs
2jSPxUpozrwKqNiF2b0cJhkHeYipO4JEi3pGQcV5gMtwHfIZyjs5hEBcidRU
97Q2NRZ5BKK5Al4YvjknX3NCyKCJA+v0VDVubWTIhZKez1s7N6wb3bxXCOS3
imSvicritMlMwAv/uVcIaw+BuLkwGRFNR11TQWzRL/tdUBfaNDb/MNQBkv/4
4ViLo85mQ0P6arImNjPDqo0yA30veDbCB1IdWVimnwABjQDPX4GUJnbXD8g1
JydnX7pIxtolQuHILHFCy7cgc8PZIQIVTS687H/MJ+FWGFNx73y4ZjScfQmP
Jnkity+bcP5QnX1wnmaRirTT/WCnBRiaPtBgZhoQrxRSqf4P24Lunvstp7lx
azbKgT7awbzhlSzOyXxW1fOkmKErPC2piba1Ah9B5zdj9vGESfAZnig7IkVP
mGe8dxmsFtcD5SRjGOMUiPxIt26UYhfmaevpwEWINEAhWgr80BZ7ENcXpb8D
rGXpwd72Kh1cIyRDJWsCGRBQF/lT8KKOERrDzKC5VWTcLguGq1p7nsvyk160
NjikXz6o2CS2DfBszN8SUrrpS4GffdWX4GG4S4VfnjLwCOoimYqJF+Y4f0id
YkDscqkA4R2p9MWfbqQfF72sV7nJdzTVzStJbe9RNbpyVlA+ML2H0uy6cL6c
8a7RK/UxjDPga2s4j8b1HabZcARxJ2GG+8KyxHQYezTnAhhDuSkkAtUlLEYF
bbz4Xj6TKcqgjxzc8MeGQd7efqcPJpHDYWhO/SvOuM+T218OWsLsO4zZL3XV
DmV1ZePka9J36hjyBUOjxpI+5ZZWIG0gFhbDOuYUokGtAioFfrS6VzgbkDuz
UZAFtdPwN2gDmAi6tYf5MSxNrhH/yFPK6KOTrdxuZAhpFrlYm3liaaNr2Nth
Wfr35gIW9sCI8tEVP9adB9W0r2r0M+Jng0W/ngLOdi3YYpomtp1ADZedeG3/
wXiNXDwIaxqPVcFp2/Kvw//fjuO32QXV/w3qNRopG2XMu81kI8UEsBolEIF8
GfsL0RKkULMbOnBGy3uAsn+gu46kMz/nYuWxLJHGLLiheBUGpthDWJZUUzPu
JFw9dCMWyYH6XyGD7HBXzvYGW9+otyfBLUoYnEbBbo9KQfvEAcoKpjz3GpQj
j8gb/fxP8iYBnFATEVH+uK6kqz6ulm/iTlScSlvmuenVQbm3CU3R0/CVUsPs
vgN3cRRa1XJhCNx4YP9HxEyMlUbQuY7/+r8bAJEzA5gsi30yV+W/dVMDmo2/
ygzUFIksysQ4eRunSXDg/fWxMXWlFCKMTDTEkkWFTwcZMiGeX2+zt7bNFyf8
fM9I8mw4NwRNVyLg9M+vBy7vxKrJ1CU98cuy6Rx64CQ+8sm474HMWiowtvHm
3tDAeGgHZXto78S56r/Dc8WnGja/FmfDfgfPKQ296hD10e0TozL/jk99rt+/
r3ULTuNtn1FtB8vRT4isDdEcSiJMgycPM+3Dqrml9vi+9SHDsG8s6FsAt0WM
t49GzJNAjpD4d9hIfIID9QluAtylMLSgAzphmSj+lryDY5BSTytZB6TmVSx/
lNUC9Y6fjiPepuQO9/+jNw4U6EXI0xwpt7lb87I8Ti76lO/jzZ8Q4kRIV1lg
usaZcsfW40KEaTvv0uAUEghypPlwPGbzlSR6DIPekq/yW1j5qLpEQLSvLgpq
PbxkfUzGsTHkdEmqyXWaZ+8fjFD2h22MLbgTyQUCtntEUZaWnYUZ+I7bZU+D
m2axPj18r6xCfQv2nPHMPsD10/D7MEijgtEwllyXIo6nWlw7qxzfMIvm+Eb9
Ti3qaf4kaWrdlwwqrCxI8dVAi1YsfKH8Jb2L0EcPMZFPWOWHC9Yo5OSmh+Ny
HvAdhTGIrH8/zk441O/jpetL3ZJII37vyw8OMDUAu4/RASXsC2VSwcXPbfdo
rh1G9kb5J+1jIpEXjEG21dBecloVVjXBOkKVeWenxUsJq0DW44O7LgZlIuLg
192QEG9oSRvPuE3nlK8NPaGb3FxIAZ4XhRWg1RuD5fU2We/WFIOTB7DvwDEi
7hhzgBPrWzVdAfpjfMwbY6DIavnHCAPctVyscxlH960uM3t6VG4KiE6z5YDn
BHDiTNxhu8/kwOLipf0lipyfd/u5LTP1pLeWJLi6NebWQ7YqZeYxRXzZGTHV
bdW4Y6TtmvskIL8ZduSeqT5YxvYYzJFhrTnTfdo2totC/IO49mtfnCT9n/ay
wW0AZZhfvTNzEjvQBSANofmU0v8GLiAv5OVMvJ6ah2sm5GPdazblZlOY3Z/Z
WdDWmx3lI/iAfIMMh+z6tZrM4SkIFV32QmIs279b3Qq7MDVwEIZ4G/ufiIKK
raNSEfes/kqLRf5pqzDnf0BXpBaJyN5HPofkpeDIbc/NbGZ95mrhHN7frAyE
lENehMZZvJ9yHcV+qf1khK5dc2rEKQae5gEYgabJJQgKceMSMv4Qv4L+1ped
PkQHCeHY1NMg2On0b4PIMT/0wmpblVovHpG9+6F259JPdn3aaw71HkPJbd+s
bcVkWNv38gxchMsoeUVmJ/NlE7gK2yW8Wff98/OQknDge2Bmek525IJZ87IO
01lkD/LC6GD96jTyaU1fqwn5PLsRXP+MxPSwny34w/B7HJgAOf6R6xCJcLUN
EE35+hplc/GBxADiUMsGoh6haWCmx7d4qVCX1zl0nOyFg2t50GW5L/YPEJOT
BDQHSPn+4Bj3Nf3xXmfcRiISGKlQEfvjCo+eXqxTU9Ne23EgvILnS2sWHkCG
MMjsWQGNXlIK+Fu+qa7+tL4LoOqZIsIhXjmC4v7qYr7UVcYZgLueos00zOuu
FuLRsaWckKhF3izMoyZyymtZI+dHbw9RrJAtYoVdwGVzH35DtCyVGARMePYo
jocT4jHXMuIhmva1LSzYKNqMRHYg6AagFzt9858fENmvzun8ogI8cvyhyGIy
WfTG46wD2IUyVBzScK5Drs5eQ4TaaXSjpXNu/UFlZc0r7EyKZSF0hkN/OcHq
h0dFMHeWL91VM09ElvfreudNlqTR4glXjwA7Q2LksW/KWudinI0/c7g6+tnw
yWpdpSQECBSdHXlpKcwJ2TVBlnGq+1LogvriyTlkxOFBNzFS71Bm74sal4zV
5IBA9QuQCgnfkBqwz1c+kDkQSorjUy9wpGQCy+QLhDPCRAyRdQtPzUCFRCQv
4+GgHIeBVE/OJTMtu+1J8Q3rjG5juGagtBYekbn1E0bqe8aAjEesJDxIBO2M
yJFHYyIzhVIfI09e04iax4DxmtL+OmNVRUggPr4crPlCxxwbwOEHYozzgsm7
0/IJjN+ob0Q3rsHICJxAbWpqXaJpBAl6V1QkFVvOo9Uc+GzMZRzO71gXd8h/
KEinLT2MvffFs3fomlvte83ha4DLd3zWTeeF0MMLUH35+H0Mq1mV+DKuUJ4l
KMNjgWcCcpncyzJfIzPVPZcuViIiVuufLzeeb17I8lBstDRCg7WGXln4PxAd
F0PaHcgpK6j++wKjyluhIbC6S1zfZOaooF0q4chd0G+g1c4eClg3PjeqvphD
CAbVnmGAL4VGCF2uU8KqVJ76kjgd7ks5ySk5cGDv4ZPEzLJ4fdElgI4gIYun
UXt97At3GLa7T9UfPJftY8ozmInLvU9rMaP42/icnr/r/b1PrwFu9tnnAn37
fNaPrGUKh6/MjCSLKpsz4rdAiRkAWB0RdH/ah6AWAEe2Umst2xWVt59J0UYg
C84yQgJKLqkC/eu0Y7ZnwrUwNJdkWYPpXeSJO7BBQN0bmHTBIJvOKj936QlY
LCq5yjj9xxItSNITlzhNU8+YZV6zNITg7YbPxSyGGXDakxguhu8twuCZ6Ia+
/zxBeTExf5IaZQVXg1xAtmYgPn4VwOetkqB71cLxScPYhbeZWJC0A7asd4pA
tLVatsgb3SgcXn3frR+GGsa+y5EyuUHNP2xeJ8HaojFVTHf8IWSkFElJhFsV
oGTU4K6SfWFyUDWQbJrurGQ41QlPYK5hAaTtmGmzZhTu6eMXlxf3ajGmKTaO
i+5O9Er2Wu2MX6opQDMHRzPWPGaxqNS3FJNMEjqiOj4EQ04g/PNayeDzO9YN
RBOW3uPXctaMwR7JKBFbwBs6NTdIBjHIQW/dC6MT47P6LS1Z2EpPS42yvGeF
tPj2LutBrpF9M+behHGrq4m4Iy+ZlmIt/c8e7PVt93ujX2KcZkOHRh4HCCnV
WJbSRTHt/+09WQANB617o3Yt+Pm9kZooxtM5131PIJDDfKrDCtoGcZUR237h
8DxCcgaK/hBNtkwSQQTCqK7UrE2seM8bFifVlQXqFASsPMFHNWhu8IWOkXzR
Qeos0zFYk2Sw+Ii0YTACda/ZI3euzqPnli3Jp3A+bFgC1xSLlJ+ufPk9N+9I
gwCKL5E2IhS2LkcKJMJ2eu6CaMhFDq8Q73PWLF9EFF1vg4v2Tb9oM2E51WHP
y/Sr6m+txk9FlFWp0yNWw2IOznL0h0D/9PMJs5EMLsZbGj2Ff5WZXIDbqGRk
m02b5M/LG3lQWZHi8PU3wZVQoTHfKxmt/iZDtkZNV75rDNituHSbiP1IbHUJ
fh5v+hZMcWKSsd+o+yfORdywPWkifpd6JGMs6zfOW8IpHkcznuFMyhx4u4cW
rdNRZsVpD2Rnb4B4CCqDCw9pIpz/EXPTyUOUB7/C/WPjycocou4RibtQ0QHq
Q80sCy9eOF6/LX99wPFz7oZZUgl3YATxf+QhrpZuoP6uq5OfJlZCUEaH+jlA
j1trkd1KTBQ4ldL/5kE27mu+MtQFDZhoiLpdq1JXpezJKRoedelRqjsGpVUz
lnNeGBy/+zked69dmEAg0yF9Ue10gbwPnFvGaYKXnmuYtWK25fvBMsFGQkZg
afw/6609K4iOV8K91+en6Bnh8+mVCXXvqz9tlBBqiXSC9LWCOylNeE2L7Rv1
zWBQbZMAd9Uz/Jpu/Rq4kPGsqMCMrDnkb9DUjAg3uX52X2ghlPmdlJsxtreO
K266RNM/TyjScXhKF+/OHwfls6ZYEWUKAsIJy4uqgZjy8ETH23x8K5pkHXjj
Cuj0okcHgd9y27lne03H7U7uD9JaDuzb0DdoFJaOrBkt6rKNgEr2nX7rj8cX
JH1i566S9+SBB48Vjlt4Ffqi8MM8iPwpCexy6XrFwMBCCGzIr9IcOrY12rpu
NnFMNilFscgi8dhi8s45SGdgkYUAP1ExzNeP1E5R2oUEVfKN3pWji+fqmLLS
6VoNqvLZO/OFcWMzqXfkkYM2wpc7wPy7KNaeeuYVhLp/1McJX0CeaGKqqGcM
T+4QOb/eN10hiPIjj3Z1gGZpn3ejp994xYSF9e8aFwK6de4pJyYj8J3CETq0
fD8N5ufPubvXH6ToMtbTP0WdVm7LidwzRMkLtk1lZZ9firb2pGFboIpnkDa4
sMsXDag/7Ik1j9SU3OxydFMAMzDmP3kEYbDIb6oaYjJawMUDgIFmujqsVpqA
BlcMNebGaWc2PfaDvDxIQk/tz/6py188iEcJT+QrFtVINM2XuL+5/KjpJNdj
FrCPJbeZZYz9sAxVg5n55GKI33WXnfTdeuGFaGzM60zJy6YDfDs2t8N4uMJd
GmVf9hgltK1px+dx3TQx0QJ1CQJB964pcig+IWd9MpHu+QlN3kR9j11AmGnc
18BOkkL0Mr8IYsimpjBtCcMECqweCqftMBJMA5EHTk+I7Hqjh/IZJsFIJ65x
uNU+LgQf98n/N29sJwJw7kxIKAE7P3+JIuWcoXq0OWWwYMOOtoVse5r2kOvx
4QEVRyUz2uUr2MQYkHp9GKqLYXVmDrY4i6KDjJoEdntOo+t9qvZ7wOA8fNoz
vLYI97p/EKbHNyhdWihastQLLco+NXIpm5AbW85sn5oqwVkasWsCXHoBv8UV
XXC55pi+xOJ4aFGzr3v0fEVxxMjQnfSs0VDxn7USQcFaAigPfm/dstYKUjbE
V7Fz8FmNdvZLFwsOq6xeTxR9gvjxgH6uy31v6ue8LgDVSmSfaf76YBNKEpy+
FDCEDWrIrRK56Ph+dJ5JJY6Mq9DnL2ytBT2S3ReTNaBkiFsWgg89H+98uIJ6
mM6xewMc3/C9JaPwS3UYFNHxBCRB+ceMdObFxh568e8ICVE37aNo1qFNidSQ
OEbxWP466FICfGys02lOc234QxeMdQR1Wsty767cqUb+Q01ktqjB0ZzbiRUj
EJxQLipR2dOmLIAMXvr/HX8Vw9haH0bgaR64YYi4kMmUqSeqJO3aKUuiVSVt
WzwbjhnK67TZ7Lm94mQhS5HBk9FP2fDTql64GldaBgNqRRrDkOCjCQzPVw1+
tAX6qkfnEq91ppE5RHndIqEoNgX8sJd0zarc0qvxYL+JvKyUWEtqOl4tSX0L
1oKYrlq48hw0Kh92w4wOTo9z6shOfnD69yExiAE5f8NSYxu6XwuB5rOlNWA8
b+9XDABQmulLdSH5Qfvj+vfJeJAUN4RLr6eRTfZR7+K9EFk0seiUJS7LyXY9
qzW+/WPw+st2fytqzWZ/8XybkFS3ifoKI1HuLL3khtV6GUb/LXTdj6uezQMM
LXeU/YwuuWeCFoNxVeI1SLwCrN7gPKm5xXKjsnkBjdugnSMqqwBEyVYIwcQ5
1XnH8vdvkpB1E/FIjWhLfqk8NWVij7GZDs6PqGKMK3xjSfakLQwPV5vTwpO1
89a8+cTLrPBtFqK5SBExPtHRkGviIyRFWdQd4ozAWGodV8cZj0K+UXC2YPDg
qvWLFsNUAZ1CdbzInZmABPj+//NuCCh/l7KI4+n1JGtFyzyIydF/5nvfnq3R
7DVLusdao4RD5WM5c8Qt/ATSq7BkpEZUYtuYqqJbDFvgG8zOBnDjo8D60rxO
ASW/NRXSekZGtIkWoaop+tROw7ikZ2IA/mcU/pH1KBtAFqhAxcBAMT0iStFA
Uy0by+OFqpTrJpOd4EYnvnhX5bfEmrB8s2rLP5CFCfFxT+x2wwKJdZ7box4e
sZXFSTYOH3xwF0Fee1FX2MGEcp/WtOOHTcPEPV524Ban37P87XvWn6cydxJ7
zmuq0T7MQY20i73FomGQwOuvRIMy0OHXD8I4ntx7fwvhuuiWC9f1dAdCU3z9
VTDWUR5FQVM47pJ1BeC/GbWAJuPanvDxbO4zH5LCIXBycBTCB/taMSF4rFrH
V1VQmh+2svZcPgJfoXXBsExJltOdVmp7CtBM4xRfvIcARfsX8qWxYg5XDe8g
kaXW9iWRkvrmTIJZuqlXA4CRZ9l8OtOHl+1GBCrmd15gghMyWoFUCyXzS3Zy
nyb0wEBPYIFQ/4c+YDE9+we2GeqOsXuUdpzavE9zp8Z2TMR+OiThQbuLfDdg
pCUu2ok/aMxJ96x2p1pEIfIGYGjRsk60D/Zqb1DNO8l5NKSCnHGkBpCYBjw4
bkaVEhjv+bOoVFuE9ImHOnW4E15HkWTQ86FQ3tLuV5Tsv98fHzZLozmqciKi
rgQmwusQQ5MF88BEuch6N4vBTDtVp6JIocR6RtDuS51ODzRZiZFFZiun9L5z
UOmKDa9oWz2co7i6TV0e0O/8Hv4TrvSEWxFL+wXrZ0ACmovCaTCOuPYnt24A
SGBfZVnWO2ExgCFw2xz/zpmGnFNS/M/qIiYFx/xgqGLOVL+cdWU/0MmGf9rT
sy8NPM9lo/s1alsE/sdePH07gJkDzQAcf5unefkowPU7F6hWZFNRA2WpQw0a
jK0Jsf32YzpxMFdKYXyvsqfwobxAVJzxhJyjft06lt+2eNlNEEIh8AxymJjj
NDf+SGpSFUT1HYaNxtTdm765jOHhl7D8CP62letZ2r2OT4uEpr1xYPvMFFwz
4qsc3RaSX0FgKrmTn1H2fH5vc9Qp08OgaoLAI7dkDnuZhdEUK546usmOI9hN
mvm43EZ/RJLWe8/lqK1GaBJihtwWx9wA3G7YqkgJ5vPLXRrl90q1J3k/bL4l
81gE3JJELTUJLWWOwjyi7CMPeeERzV0ssYMopST87XvhE7myJ6ExzUW9u0eH
sOYGlhl5waQTL/OC/Da7z9DLB0X0vGMeBfjmaoUf+HB67YG+9Q1jUvJS04fW
qYxGkh/MxnGnWE8dJFxmM51a1Bky2d2aW+gJ5/B/5/1C0TFcz8My+0XXExXb
kLITP53OkvOuVsATn8Rfy3S6SXLwTQdubITG+DkCGyx60gYIvBVhQmN+YN4V
K8gQsxDecsSzjL2jOfcnW/Jb2RWLg6APompu58tlRYcPG55wkXogFQIo4P9s
zDuWrPYEwqxMOliOkW3YUgIlhzy3jBQgk/qtqDAAxYmZiRpQ8w3OOvw/9AEs
11MnI1fLDMcRgvAykSmAsaZF5ZNDWEWihgQTcRjrANOagTXQv/NxIWherHtz
TPB1ERS4hoLWoxfx/y+c1TY+2ri2YsU8gkeHwQGX6xIjGGMpgjf26Kp3SBpB
JW9QWIcPV/2CfkPObGSYpSSZHxlf4rVPUSiVXCgsYMfLXhOF92HF16979iQ8
GmJsR3F+saYpUMyOFb6x9GMk42ybV8kTdv9p7Ulf5klv1vr3jZIfd48Arpv9
t4KmPiNgM2+rJOcUlfVBfrWkNUNJH+i1PdReDXVB/4D1235ZovAAR+Bxh+xT
bg7lnd0aMpPpxa0phIdHU2WLBcu/5NX2WSbMSHpteKSuL6zusBihZEf9rt8z
owHWWrlGZ7Y3fn9vJel/LUKU2qa2ztfgV2ZqKn7oR71FpOV3nLSy8ZVrnFHS
EFydGfL4Wcoor2A6APvbFRp2Vba+qBhp/IxyHwgTw5YJppKzU4nK5KW1SJ+X
Szwu33DEKg4eQxcKEMnuG8ZZKSzvbqkIu/WDaFQR/tCVyhcqv1fjwlVIiXI2
OmpLs2mpPUtRnO8aSh5qsa13ClWCTNokgkKnrYtUvr+lIQj/BisCpwJspKa0
vgFYqDt0vNkiJIPPghrGTYtUFVWiZ7+oTJ2vYrz24Vfs8ctwgAj9u+BXHS2Y
igo3j+YvHNS+BE3KuqEefHa3mMMqFctIi1npA8Q8u6Thc00a7BhT+AgWu9M7
akzst1jHdYCFbBznJIx5c3l/Ih57IWOdKgkP18s+TyR6RHTT3B1rSFZ+lnXK
JJ1DqJJ10BWZcsKiWo6F6by7IsHUyStQMPkxBs2EcNbSGa/4zrD6cd8TCPhT
R0KA2MykFseR3hFv+Jns9z41ST1WotEVlHzsOVmSsuSnyAozaEYJUb2bNQqh
XFFDUAcN9cKiJNFCAQ104+5Ne8e07I/wFRtL19s90SW2U4FCMmVidxhA+t/2
JIQciEHL0nO7S7OOwa7QLnPOYMorMiU5NZ8nPKqzsVl2/DPAUMUyB+bXvohH
NVu2AhnHUIDk/H6FM9T3lBNHcQPdobIzCRJBhc3dw5kaqzx4Qnypcmo293dK
ZnOvTI6/UuwwahBxQSwouRPmoz1xVEAug5vK42bpCWfbrduEks1soGlV3Uef
uDJib8qgYWJptoN0fO0P64K9awG2TCkFk1rruIsmdqdieXsi8MR/pHeMgf6a
FnQvTza6l8GQlOwTy+NnCnf9fRO4W3JrvN2JSC6EU7Fg9sP+uE0Ji86PLe6H
RiS34Qzghre+SL7LcS2neT7va5b03jJxVZo3Dz0T3xYLGqA5ncXFsu5ioqoP
5TDrR/ILt16QTauuJ585R+F0WAesc6PZmWH8VZ9HoS5U7387qkQsNYyVfd9o
02J6H346pp6vrAJVF9CGVDx9YFDWB4OpcpQxc/1nhbPFrUaU9lghIzlMSnkp
YsJf6x8qckLF86OKVxS2Ge0gKNe+Y5O8WIXmK2i7ZYLXWgPjQ5VORudRbBjC
ZJpnulxCu+AmRznR9XcnUP1HmgHIi9XgEp9fd98TWbMATqerILl/85EFe4NS
H4lNcKaHnRKGKFqcmtNv9nXdOHCiyXdrXutIS5OqpK+uB71DFTpvTyRd1vy7
aeGrRVbpT/JKqaHFsGMV3bR7JGmASMVPjo7bW5D6r0tijaqF+Al8vg9ys+hV
1S/FqvwSjVm3SuSDdfxu17p49PvB9smIT//Fb8tQ9T4hQikmBrrGyBXxQcTN
XY5TsYEj5bOQH7iDBElsLyeC6BlP3YLDhJcRsSqiAZq+sDJ84YwhNe4jBUn3
C2rJy6TwEwMxPSR7h1UNBsmLL6AY3zpnQORQUtmDlKOao0X6+PH1OJdNmv0A
jbNbloqTgQrLgMUMe4wdyISuBaXiTOjNoskS3dFWvRwnlrT7e/gAD/4vo8Ak
CqKrJ5JprlO1+xSSs2cFXNIenUc9cf17Evf9Td9xfrXW7B2ghvW/IlLtQ5Z4
1MqTEtL1+OMiNj5PB+pUUjj+cx8Mbv4LYLJbY+vkgdjsWcvo9KLXMnsBbygN
U65HsNNit0UOxnjrR+0bEe8ELy2CLzP6pN0xhOj/R8WP9L8fx3twGZKWLCD8
Bl9+IW3U3oqo+bqVhonXtX7O246DRvBOU8y+jrcQ4RdixrFWZsHodW1VFbCo
OMbbuyfKCmQiDxAA0Ya/WCaZbx1MuJ922K7iXQVpXywESsEUAktFxmqijvLa
QFwTmAwXrXYXGPIpW13sEKysThvohSvTjHu9lb/Q2zX75SFeVLuageumiQdZ
mCHyQAjcwBPGSV2RBN7k/sshTQYGtMvhoUA5adeAqD9HnYFe74AUYFQPEeIV
GsUnwkhaO5YrJGWAZ6Xsl1Alg+KCtUelJSozuelVRe5GumME//DPvIoxw6Rc
TrAOK1qbNlcRXTYMMr3I5l3iYL4y9S+yDIMYBDV8ezcfGSwWFK4C2EN4rCFU
6mwbdP8av317ZxDYPjQfb069zNebSDjN0ELsPuDSgoGQzB2vr1IEcOGxVI6C
4dExWIlFTSwuwjHmpDN0eoPJYkR8mNssrMmL7UyUxzXbLaeZcoCeWUBTufPu
J9Z/YKHp0uAp/y/iF7A/BEyG5LMXKroPesGciPfA1iCRwYc+CTGAY3GApMNq
FeVBUsAvkr2nX2ew6n8GP0aa1AZHyJ2uoAZOnzUlUd+MsB8smbrxT2A0e9Ni
feilFnfqcke+/LKPW61l7F5E1cs6zFyobpaW8UQt1GyhvzeFo01+BEywnbv8
i2tSd4yWNSoj3wvuaWa1twlZ6Fb8xJ/oNi19pmQOLcSalF3su8J7DviyiTEz
g5JENH5DVs+2zRQUI2SiMGcSvBufnl+mY6eN8gOmFcR0qwIzEuq++z237MBd
g3+aqDg4hgzuFChJ8hdDpTNwqk6urQZx0HrHnnIak5ysBy4KsNLJ0vM+E6mu
cUz58hq1e/zV5NcKUjCSMSvFFJ1sv0E2qCrb0PtFgGeaMGBeCrMfQBdGl7Xl
Lx2kSOi+YTqL1Ya/ty5EDiuwGvUWvk+b+IEaiWaVmcn8etx6ldxbjxEoBldy
Nx92OqYIGzpvvtDb/Tm9k2C5UJ2+rYDEGwUoBT6/C7QAoQ1YmQ4C6vv3tsIR
ujcZR2Jfk0FWfuWrpvTxd2/RHo3GhVXqMrpYalvA1coq3RIUCtodj69lm0i0
RoogeEjQI7HZN78Lp1kWDHNap3//a8HQMvPj4nIvmG3gx6eTVX0lW7aACTco
jlmUR+6HyZRMNqQJB/Sm2LmAHbx4tJTgSeDvI1OvSA1dLq9sKsN0gA+ZJd51
SIQt6ewuIcgqLTPffRL529EC92OahD7bLPnniOlA1AnznJfwrNZFXHiik+fB
oEfm8YPqiIaBAsgvPiwlL207Qn0AwpOIMYPl8DQrYe8ydR3kbcglpomTjP2/
z93GuJc3qYGjNP9mqlFkedkd+otY3xD/+BIAdt2eVyG+gBA6I3Lii/7ODevz
f5PSAkVRHvSZxT/KaoZeYWITiyGJYcohsvzGO1mEGXKxrGUH+mAnw1eAWk14
loemWtNa1MydaOUQjHbztd8kBLesUAjg8wRtDBIwk8/0h8h1j5KiaJMa3d2u
AmVNJLKTu28Xhqne+h58i1VwkicFwntnMfDYzpTJyh9P6v882Px/r6N9iDM6
E7LujL9A8iPHlTrU9EB0EQkUDQMAvHiLwv/2T868rHMFLy/pDhL6RsOxMfmh
TSBfLVVrPFN7JX1rlhfUhlEo7r0ph2GkSEi77tOQSCjNJuLOBlRAJTiRNh19
BfW62XlibEm4J9nu/UWaiHn3D4ea+vDoGcTBF+UWWBkixWMsiPDaCq2ndesz
Y2bbxkhbtQz4cd5wzWty+qs+hkXHNGQAOAU3KAg3BBDaA6qtKtTlyU4+bS6B
j25lNTcf4Bg4GwTCcUYIfr4ZdbZreirS21MPXgezM5f8objqDhuW5/eFqNZ+
cCpd9VXnlYjBIaL+wZ4maDfpG6QpHvn52JteK3Cy9K1SZcUQutTIr3rJgvyJ
cFQHO79RAYxWKM5f/ly7m/FR6YAvMsg+iBffA0F26ti7q6dkznOSloi9MCB4
MUzIL+ggyAw9YUhA0Svw0uaGjhhtYmZskWFOUwwODIvLZfrSC8rzlKDmbp84
0i0h1jl577+QH1O4fBCzqnxMlEpvyGwUpsyZEjKnXxGG45MSL2T82ItKjiQc
ecK9YRgX9x13vuk0QDESM89KgpAv7BHIGXzlVmFkbuGJ5UchYQz5EpKULzyL
cy0zbfTH3gb/Ee5Ly46rnMnGxc4QS06lGkchveqvt1Td9TcUZedNaey2ZeWu
5XCwUrafFEK5t//rW2NJHM5dobbyoM7li467ItdIbRfvq8/S5eFpLofSD5YM
cyLl2Tk787SpyCou7eb0GUKc/yn7/rC5C7XoCI3t/weG0OF1Q0tNacbBKqS1
UVLWtCv/7yNF8I5BUSM0TJvO6QSGLhAGOx1BkbC+bPi9SyXYXv6ymRNl8DUo
t/0AHm8aKHv2heGMDc6TXZG3sPrYlW9+G2ycLUKfOJdw0HYoJtNNRlTGwK+I
2omwTvCckA2doUwlwvkaGZbwJPu2nzXGwgiZRxEHSJlKqSKq0BemPQy2nwJQ
PLXwW4l05tljS0y8BQEmEmQ2s3NJ8OL/yrYAuCWhQAWi8eAxeVmbqI4DzEJq
zerIXwOs3nJzJZi1yMWObM07bwkzZR4G/0ygfmvbOkBu5ftr/0tmoypYn8zR
9xzzDLqCzD6VAXAaKIprP8y1e38NrR+YpuKvLqxwXm6AXl/1IZi7+Bj+Vb82
t7Yz+FvWo0jlVkk1ObmgxYTUUP+XH0YR/dWWMOprfcH4DaMlEBFnWlxoTRU9
jNXtr+L6Sbv0LO4B+CPBuwMz0wrg+hAOW+4+r4CtTLxc6VFyq0Qc21EVRHeb
c9eGqHVqk41oatexhzUq4tjYOkBC2zylB3aanExyBDyHWBz3XyDTtoMfzwC9
rM7lqD2xBOI4JIpt545ITciMvRfbRMm469R4nVdirP5qROW/Ib9wIXlS/2hZ
UI810zUm1wEBGBSRqT4MwnPNvDuoeXwuMgLNuholj4oCFnr7e83og2OmzxjN
HS8ie5Z8+A2iq8lN5Q0WRkQE9Cyx/1oMwiWTmSEhhNJ7wEzAA9f/S78fqNcV
XlfbVi7AfpMjP93/OUxIwAof324AjaRyltzqTaY0JsW+dXu2Gc/juSQNQG7p
d9rLvpeisguKAgCCpeRWqI//oUkPpyKvJNGL++a05IzMK1rYH+L70UY6usTT
eXEy428yn4vtyEKXCWlDiis+mCwvMKPeCsQies3RWoKhW8BHXEXOfoyGroXy
2XV1UU1Uq2RzXk673PxrNd3TfZohiMX6x6FU/9wiyOhDM6DvdXdm3cWpJ4Qr
ZR8h6OjjzlT4K5L8wzBdjXnU57XYSyg+Bpcy8oYwywmQlp35lpskt6tVKOIu
C4qoUPwLZYL4lWb5cf9d4V2qca6T98asYKWvUzTXumbX+Tr24NH6hU/nwO2P
2E8Db9IdCVaEoux6scbBbKEejGoSoGVK2ax6dFPlM8KQJ4b2sTXkTECIOtju
CtxBg/ZSCa9qjf4thE5UDpF0YgiAkBLYuEQpzjJPWBmpMyiKXB/QmB0/3/uU
TsJgWS1F8hsQGSLU1G2O/B608+TF3dX5RN/DkJNH3OBWT49LbkkHfLn06t44
gugAMbHLOefQLb5QhNKN8YJy4UzznB4kqUsK10vAHI00YvKAib9x0zjKvdq3
CPYIL8mdPI20YP3GMy7GSr9Hi2u6mD8OkAgzIRNq1UmK2wAh8kRo9pGceSKr
LNgCSbAUfsV0a0tLXNWPOW+U57EIfgn3aJ3v0FqB/JjVRnEHDNqTa+ywKlNe
ZfMXRJ/8ty68eGL+dEB8f/KSc21c30gIpc9KyBQ50TqfqrTa5HZec0os344t
d1zwMXW41lqABe8VrB+ECZzn1lPfHd5SpL0+LLRQpIF204TdqHfkeweVt/Jw
CHt1Vnlj0MpzGzZw0jRo4VGln+fjBRAPRSrDJMTPQbVEWiuAro/awpA56Mqg
g3ay+LNvZMfHiLmYW0nbWCz+9g9lmrjEhQDMjOpaAYMQYk4j0yCV6Md4tu5L
/9Ayy13a3PZMip/ktpvocT1065ihmkT187wLWPfLja7NSKOilq9WZ5vGNiap
z71VkdZlF6VmsIAo+nQVKEb7FMz2zp8A3MxVS+WDUoo2G6ebHT9N33ZVegEn
Qai0AKKzbyVApiEDjgSLEDvGjGvaPkYbYYAGY3csbI4NDIflWV1nNZO1uWqJ
lquJcDi/1OCSMeD6NMY/WEA5V8nEkn5/sVbUEraamq+TtwYfuewhLZbMlFGt
nckIYojxCP2VLA2J4Vnk5G0XuN+qApOgKdib4LFf4+RftBkTWCADlDd/L280
yHEDjVr1ILHmFf2k0D5uGMqseyFA9r57yMeVhMK9EodhS4OFCWQ4OUHSVhWn
of8cgEUOtQ1d+ooOxQx3lnU8Fs/aO036jwS37HHtWogzVz2i9BONZ6tzPokR
SZyyKOvng2r7dX80hNgt/6w3EbTTzHKZ+hQ4bFe/lYOjgOWgTT09AGKd84C9
l6LanNPM724Y4GDNB2AB4Is0ZyxitcSn8Ue5PebORQRRU0wxKpmiV1q3/Vzz
Awrfc2rgSOFoFkuAmwJsPAd+kYTp6K2Exe4J00RRrCLw7wPT5XK6MWQT2UfA
p27IEYcbzZywD1vDMgOlg7xGw+krlYc4dWfFCINLYTLjI9bEJ2bnSNPCP/zF
J6qMMXZQ3bzYJPPXbo8XWcXBL9xSpt4Ikj5DvuSHl4kpFZaHx7Rvun5Dcr0b
RKqd6qN7wr3dcir7VM2Qm3izmefz2BBrEXFJqFyatueh2p4IvhMc2VQDmCwn
X1uQVtyPLK9bxcsG2N2nwh5aQtiKYnrykJ4VUoCE+Ft+OuRWxx9UypeG1CSO
zBSquGwShs90/abJDbqYTtBg1JlmJgOAnUfKxdlSdqNjPo94JNbjgzfqYb0p
3CPL0nOzBBpol8pPA22SawPjXdcsuBuacU4YHSfODACdRSJU+Yglu+oNVcZc
NHQcIOia4/cW0ytIF6COJLAo3POgycRuE8PA7RkhC+zR1DzVW5EKxw7BU+4W
wNPvehNVhHKTPraN3FqQoKx2nfVYAiPhi1dJy7Xqb7Lw2c/0+2J/Q21f/PZv
0c672KqNAS3YcnFle5PVNDMtoKkBD4Fscuy9UEVoRE46/S+fAg/wjw2zGPNx
xdFysvRO3I3t6Mqt8HJ1/oI6xt2MSPg0Q9M/7OQ/MPXimlKWJaygwcQQJbT0
cXIKSp/Qi9hyPi1fCw9I1O10pRMKcx+cMFEY7dw+5v9TQiwjB/7ZOiEJJS5g
J91opnOJ1j2FLw5LyHNJd5iT3xFDVlvWVraVXFE45gmO8o6WY1laHCm1kAzj
j2I9kCpm3GVB8jXh7/nK4L2JT0hFhg6cutKVbr0gPzkkOKSJsfuB4T4AEXDF
seUcYvUSeMlea0SG1884TYmjfxhK0VNE/3nthCxvbbOvl0dHJnsyqx69SRuz
S7yVEl8vePbOYLfbavqwOvg9Hdv7zCHx/1xno37TGr+9+1ioUiBiJ2sn/2ZG
wW5PmQ+KMFgFrRIPoV7Kb0MpUZ0SGKJTxGw253TF3Tiey85MKMpg8Iwimk6t
xsFP+nKykcCAmodNnwp8ROWbQmM//mpWlRTc76fVqk7U13u7VMxbvi8VkHJK
xmGBbqyk6q+1OCbHu5w66nstiSoPQwQsRPt0wfsNmZLKR4YJLyweBPuQwnb2
ljDuwrgoM1ntBlxldTbTFyCgbqABiyy3x4pXGkeMcSv3rCTUqc4dzzk78pzK
van10p0ceN4UGOQuzDh0VSb18qK7pz0gjpQe8i5o1FpYaQLP4aPdk1lO0Ag6
q4uvfC+7wowxNijabJSqAGR55lStdYyjzQ58NJA9kiavUwkbVPnbSB7ZhhL+
DVNbUC13iEtGWHli75+i9fs/+LVL5PJku0B7ygGDD6lL+2p4ZD08VZWL4Cmy
ZzR+3U5CviMZokVOMtt+msIwUjEFOd97KOniYLio9H+ke+u6AG+y6kx8iFxT
nEYpDnkVcnIQb6KL5N6jlmJ2c1fiHB5slVADjiAr3G9UeqCmhSMiVwttgW/V
Npxn+iHQ2dVe31Foz/OPnW7ICaxvw7DwnuUmZuWbokXmThQurrEv7m58mme1
bbm4jqPHeOLcI0loAIvERkV3qzZk90kde3+i5eaZP1mFd1qbUGTDlEEXgX/D
7RkTncEgWWhqTU8ONgbV+yjzEjTBQp300guE66re90Qszu+aQFRl9SLe03WC
mQ6OlO8uf6oXuCMAG5IWiMzB4YubwAFh+sm2K0yvZg9ZAa4hA0XG7/JyqtlS
uBoDjTcnUGw3sdKPLBnhPspBLlyZ1Ppon/gtcxioEENhcYNiq4RitOHRisbA
+R+RBj+NAT3qHXOGZWBh0eR2APLFuV5WK/lzc8E9cmCqfSQXy5Ts3Y0f2cuj
yCMNdeeNxkqJh7I2MZByIZx3njunf9Hwj7j0ZgLdvWwBI5DrQcijoDQTwdzZ
FvZZ/ZI7RTC6MatGGVsBkIUrEkVxxIo3jIEGd2zkKXAsDIrCZ2dkGU9Hl70J
tBYk4ql8FZjSxHYFNXiis+mYQar893lxOmuOH3NEG5GKiQE+LabAJ5HqdqII
GbXC8uNQCJC3ogz49d93vJ/eIQfqwI2nJwmaIhEkuCjwDuyQakPCpM7J1KJL
AiqYNnGp0oRCNJ8QNTlzHxLSEpxFx2Y7oPhve98aP0rJGtKSRj0ZsXa8T4bH
vrAGYyV0tkC6CYyNsad4rKzgtR+0Y2zZC+x9LvsUhUPGMC5GS43oyc9u85OJ
wClHspVUY5O/J4bHL0IV+AS8myfUcmGpDWdEUsEw3YlImTxVF5dGex92Tqbn
uLIu9kDE5CBz2/CY0WlpTGCMT6ss6gU080DP92ZZyIzOAZFujOP10BjReys5
ZWJAEzq4TJ3VKks5xNxxa5MeP6y/7Ka9fkd2yYQCA6VqPyQZP81G6RAfN1vE
QkITXH++MbcIHnpbYI3weh/Oncw1bvI/iYzmpNOUw9f+nmI1dIhjp8d3ewey
QTU6Rg6Vgeto20U5wwIDbw7c0Wll34/2AkTKEjlEIo+7cWG32h5M74b9bm/z
93tFx6iw5x+8FsuddUVzm6a9d6fWRB2sD6uKjKhelUSwAr6N9vt92p6lUsGS
aNjpQ/Z8OiUTMwgQelPGk3BgLwPRA9uo8l3PJZ5WeTbA57S5zrh6rRsPaC5R
xKtNOixQ8ZYzWMYFTV4zaus0c6UJXxKfMeIG6yi7QcfLtvDElU2Qu5SP2AAl
6cm6CFLoHwOpBifKckMo+F+/Td00TfV73CjqPOO/2+8EfavY+SjWNsf/2zpY
4vF3Pk2D84SADJlpFflyC0tfEmtzMuxunNwUSZBGIBuwoJ7BokA8MpY2DoG1
C0tuPcFpTRa5eP4ZxzPS8OHRj3dhcxbuL9LebA9U0UEErYxeFDSryGogG+4v
fP1k8u/BQaL9IQb0o9dPVVupIihAvhIvvK5shKaT7B3Wuh7Trgwfvk/KeKUM
ogfkcooyifwQNSeBdRqHiRN+ft1+SlvhEYE8n6j1Lnsmu4LA6cQAkUzrlFrY
gvmVTQiVzBIWJ7LDzHJiOrz7XsFGHzfoWvafrIoCpSXIuU+JK/JfB3DodGd+
bWGKMq4thj/KeWQZ8gtLOglAGDwLaQGSbhwGNRnsj76Qraq5MDkOpDS2sUj9
nnfRsEIkt61gY66+dAk8B0lKt/6sCQVGPnCPoM5MrhHlFUrz3c3/9x7GWJDc
Td1QJ7qYZDHuIRFPe/m5AVo4GhdrFKtA6Pndo5jOu8mHPgx2e6UWhY7o+B3U
mgl7EondxeZidZpfHK95J4B7AMKDjq+B4VW5nteqCsIqot9V9DpptJYCEqYc
168SFbFPjo8IR43pXnro9MIU/UeJn/VH0rx0cPjday0LvrqXgtNdEI4uVAO/
7h3RncE7j2iL46D28t64UVy1GaFKLU2thYy0G5TGguEX/jRQn0Qo9pvNHdBE
8vq7z64XdB2wqrNlMyH222EXygGBeaFPyJPkuW1CjLvbsCp980ztaFNFHYYe
YpN5ALaihkUmkFBAKlRnQn+YGTDzc4spNzM0UQs+xjai5LqjmQkC9DdV4OUn
BHUv0ewVIQHJuGUejMbo0rLz2cO8L22SQsgEKk4JUa5hOxLJdZiDmsVwKget
3fA7xULe5zW3hEFwosis4JwWylI8vN8kKlAHowq5e37jXDWPYn1hI8jfUmKv
rMIQYE0nkbkICgW5oq0xWPnerY3roqh1LUINedPODlCh1hEP6dTxvZq6NkKH
+S6/lIWG35oAk+Q2l1d4L+bHmnENn66KWOdApAalxWGL6oOn/zOS5robcWzJ
fcelB4MG+fByOLgr/G+vwCuOlNaQYHmduNk8ed8jMKUuM06ROkD7uMO0BzTm
SUkYBxNt1MzKe4huyrPxDOdvr+AhIyNsO9fPJ94bgi1ShL7Hdr+QTtl6b4Zw
WMZvimyMcX96bEm/S8yredqZrzAh4iRGLtFkaBrzTQRddOvyBVnaEVmcKeK4
I1sefXKZ3qyHduLeRFJWsRM9ifSzQz1cZ5aHrG7y1sBrKQ4EG1kUB6J7+I5Y
pH83Xknr1mzTYQI3dY8LJGJBKjh9V1JOtZiJagfgp8h1CR9sh7r0sDDFaK2S
ErGss43ybh1w/fUqc205SUttHDe1MXVYDmz0umMuw/PApIgO9sbk9hS/BuLM
RAtmSBQs7csq0+JLhZ+uvDeu3veWVxpohaZPb8+y2W/M5+WovjfkBGF6cPtL
O0d+O1F57ejJISEM3VPMczfCrjOgwgDqilfQtoKfEHmjvJZFpSEaO3seE0Jo
v/2P0onFqgCwZh7ae8Lfb2VHGReu06BThcF9mNrJBgVZREE5zfVl2T0j8ICw
dP00FaAl71Yy1NKG8XeGgmHEspG/G+o7X38T6bqKUsmcdoHeoxAyqDot1ani
e2b8C4H+FA2Cur2KdESsbAp6TGluXRpdUbGT+LhxMhohbsTGqipFBXg59oUm
+rrQXr7Rb5D9ndVwJtRieZgmA80VljIqZ/P4OgjPzPaLONDgyr/UpHWmQt+0
B48e9puVCqGfgnFlZ6Jzpksyravk0LwxJl6kj4v5oe47CCK6YLU1FbcrbxFB
XIovuUkQ1GDGpPHfxXMIS4zi7qCm9myoLOTWg/Kqg63sN3/pU38apq7OR4v8
c8BZOwvn6R6iezxa6esGToQKCOETT/l6zHFskorZHA48RsWwJa+hSS34DWvA
H9zu7NA8z2L2QTmfudRcHT4gS4u76rINEWeqp32yrWnz/Etq1anuUF5mZ8u0
dVsQgzk7HoPRRduKAC+8jyTeZz9UUAAmIDLfnbRudIRtBGi/5Xhe8hiXBbkT
x5gD25q6GJ/zt/r+Dgp7YolGqRh4S+WydvsmZxaDNTwMBntn/n8f7ATYps3V
bvC9jyxtRBF8G4NxDTjp27EsdbPftTo5FUewI/JlfTPEB7nGR1eaO4kiQlHQ
uDjzLpngq5Qt8WCfgT9REjJS1Sx64uWKqgB04+nypsHP7SELzj1ZCtycfVKG
hnXgiWVrN2JyOKynemzA/RPooirFsnWtxhPjIA9p6idU5ddgXj6/hP3eInYe
bIg5cCX5m6W3shh1//srToKXdGGSwrOdkf26NzOqERj8AqwqVw3p3x9knlyl
d3mPDlOJcIYWUjgOBmBNCE/03H954Xxr921St3O35QFyS6LCRR2jfXk70zAG
aqbnfktho9gXFBZWRxbQSelA1ulq3flLLvXZGQ4QsIlvNVn3bl1UwHtYDLT9
smPImozZ52UpBXZdMKDIXzce3sB4EF9LofnGBP4qSFKF3Uuic+6CMvThtfe0
WPVVVlh9fYwnd/xMVjVTYGIJHIC4P59dWiozK8CE5TgTGZz3H4IjaKV1AWeC
GggOslbNkx9pvUFqqdhgATI5lgBYmGGFwk+BWwJEULXOZR4kcLjtdlbxQUft
KGu+fWTEAOZ5s/3lbzxLhX9Mk2I4I8hhILEFML0vXneQIb4e2NmnweSQC6LH
V7zmy+/IQOhdFmIWu9qK9AL4jp3Mgsdj7LCIF3Ks9yD2TCSXUUJHSakT19V+
du5hcGbMZ4xilWVstaLi4vgsYv+4mjUvK9n3jhiXEfGVc96ArMa+9KV4rEvq
mVLbqZ4RTonXrPLSpHLCoiT9oRW5Sm7oBFFkpGIZhg+PdXG7qVIeQ/coNhYZ
l/wsw7WE55AnpruAMdFdcY8WNbc6aGy6us0N4J9aVHe3eyi6JPxySkuSyKXG
7bV5gaKMvjxmFLdGpOjrpPhf/6w4/ckswQYqvonPB+Bs/103KaRJrMHUKhKj
tu7dK/nF+y7ANypQgtirKVZuaAcQsaIbcHwWX1LPJL1+SWZHXwZ1Tq0CNmmU
++HnkyR1qyle8VJ6TuFZ8IamaQ+MCRXKQMzy8pNDW0jsatZRQgdvi5bs4hSm
dLBBqQI/YPY4nx4z3quzuH8IuFfcj7wqYvxaruvanzf8dw+Mblf34hWR8+DW
gTsr/XeepzbZSvTRNFB3w6Iw47LGhWxKMea7oeDm1aMNvS+/f/J4PZfnNLfs
9SJiVCzhBQp0iROvO13fbfqSy7wgEz2KLpKG5jMOGpyoPQOuNTn4013RvpY/
Q86z98zR1OXxEUzo1Oi4rCbV4WmtKYuaDXJD7bUW+CUBNzuVKu//dhL3YmNm
ObRKNLNHCMQtbeBIB+QXfpwvXPBQdsKVb/BI1nd0EWcdsmq7Cp/j0Yu7j9o1
4eagdBICBQF/bbze/m2DJf1iQdwZxKcaN8us3yEZt0dp1ubXZsjFymgYWOL9
kS0AhottpGUoEAGJUBQZpKlHKjzyUQvksPp3+umnvWUGdkEH9jeZtbg9yXYC
nPTB6MdqrR+eBS0kPtt6YfyMwriQK94z0hkCw+r3diJVmmYxNwL8dDn9MVkI
DgsV6GXD8eeSAPLOYjo0jl9rG38zi6m8RMtT6TFs/ydWnHdPP168PlLwWNjv
B8mILKMMW6ufrKxMh7QAVDyoVxqVJDYfwd6IE614sDdNY9oFUo+mbNffnhfv
OgPvtT3VMFQT++tIPRLi9DZKErhuLatIovTam5nCnWP462Wg+X9KxylwHEbK
PXrFoB/6iwYRrkJwxbG0wJTaNygGl3qInBPtY6DnkP6FH9Yv2xcntAOijyQu
iTSvbj9/F/DLsHE31ojZU+AiP73cBLJVmoNpCnMd/nO+NoA+RKvs1aV6taZX
HskH+s4RWUS/MZ6+iNUlUYvP9z9cvBboLMBcMq9Az9Ie8zii+N6b/d8wpM1W
Gsp9lv6PP7q0zQf/54iLYi0e/oZG3kPg61rdAY0kEvOG6SDLrDu02m1pTXoz
+DGY/kAt05lUDwl9RgjLekNocrPXIOe/+vCy4RwhLMZXim9JQYZZwZEhfzea
IqJM005pOZuqX/bISynwLAE0rJnGHSZD3uzJymM/P03nMm73soMiDx1hJDoS
bf6T2zd+F8R1YdRiV0JWOaZ/KavPSMpG2khH9W4DbGw1/BO3mCzHAp02LGMu
Tx89225cgIFP6rv2cSfZvWJqCRdVutTTlQGaK6Sy52nMPp+DnoApBIxTINcT
d9N1rAVKFfqD2Kgn9RPhb+5IMxZjj/1mg7gIb82XzN7hkUa3buAy3GFvotO0
GH3Ln7CHqMc6Kfa2kv17bjZpzRz2shzs2uzB3BFAhlQLd1QbleyiEDPnoVQp
BMpU0xixzDMG9cofUs/0leRU3UFaGwmJ3+QhKU50zRyZ83uAmQlwDTayeiS+
I6h4CF+5EmE9vXdKzeRrKl0wc34seI9unuwdwdFotPJFAdXEmHWGTL/amv0W
0XQvjq8K3r6X9jA6efXmKP7A5HckDRBypg2/JScc9pdAJXp+IraNKBPASaTq
gh8fX26V8Zel/HDsIjb2oETNLHR5+GwIBiORGP87Y4l4fkTq+fNTZYmfgkb3
szY5FVqAfCbq3M15EqcFP5s9BUU/31rdL2FazzRYg2OQXA5z2iOHzExIZYT3
ZDP22p4ynMgSTHoe0VPnoERa9SYytxGd8gJZ9EyrSuauAQVT/0woFEnF7nMm
qI5wlLKHuC58nFKS+1wvLmyq0tokoFRtWBDZE8WEboavbGuEzlHVnqRVl2/+
gq3jCjsHpbz1r9FR82Se5CdYTdCIHEnHuF2b7X6slEpDmZu3j71ntDPYgemV
NzdlyKbCy9sGSLYGngFChmjQtZo5qBG74ucT1AGVL/hJASK+jP1L7rkCq4W+
81f61IYFTFtBme8vqjdVxs2auQ+7dRzlF5MHeyu0MkprnTP4XIZXh0+Tsec9
Pzr7OVrtADeF3qE76KfSjox3Z74CkPb2cRyRr51gcGFiZv+0Gv541UPzpEpU
bbwAfI0/ONolPz8dnInITOn1z2e2ojLV11FMLssWKvrQMyYrmPXirhPB/ZVg
wYvn5cgLR1m++N6JiOACuDE7nRbUGLMZAYL3juvl88GnRMCiofNJMt+rESjh
KdbPj56doqTk1JEXA2wNN9bQZGwvgY3EVoJdmCbIK6LVce1YzM7S5bvDiRuO
pn3eUAR5mVHPd5gGbzqjwOmFbfehMiy/FtUO9Mf/9IU9QOW5QtWHEAK+7Xcu
hbSf0vc0YxpcRwUOvJa9uaemrN4rNlhZTT7GwbM8Yqa92p/qKcLckK4m4tJy
C/7YWQHiZiTAjAadbdw8tQp+ew6tYuZkYHe9deU1lUro1oYLLMh+j9gyYWDn
fXPTrihvSRSQadV38gmYQ32pgMUVYDjm4PdzCin4K8Wpilf/YL8RK2+e1o4j
l8hufQcGDxfrv8kFUbz37KjM1eoC+BYFJJ0X8Uk/9YxUP5gka63/x6dACHNq
qBk4RTEZ9S9nq8YdjG2l15Mwy01U0e+4btNB0nFZFyd0V6aC2i1M5e3rZT1z
akEuLEDo4gPBzomFnXXtxTphYG2m6T2psB7NwkIdmtAdWCUPbIJCEZsOPnXR
lRX1It4qrGc5SB6ruYsBgNng5mxtkPpHbJcicH3b1jhImwCcf5ZwmxPRCVEH
ApQ28ke+nLfHR9JNtqAhJz4aFZBKtk5jxlqK2Mcs0V35rgWjOEubr08i7qil
4Z5f1QdK8vgWt9QWp/9Lvof8WyxlMkrd3WXjo4gWSCLOm0OQD2Wo860Tv7yf
3gBA03y/EyAi7IKKqHbvwhg38BCN/3ckKDQmDYmnv+oO0/KKddFdOW3KioVh
pKvqCM5BWhM7Ks683g3R0pbuWqdqG1aiWGzOIMoyrYnoynh3r8b8w+0LjiZs
TQdViNLLg0jBxzIapAfoGQn97LWeJLwHaVHE7pqz10R8cWcnwyXcnCariHRy
o+Wh3eUMFAIWP9P8tzwjT54J3SDqfDabCfP34b/Sem1XstJvUx5VT2D6lME0
SqodbFwbH0XKzCvOJAsVUcTh169pg3YGY9dKEI2wd4jH4sA/hopbiscUPz/M
4QjHZsK8MaqdJqtuEZKkcCAjgdbLcpWCiYw109le4uf3/XaZ6AvfiM2cF850
sHUx2raV6nQHA1HWoFZkGrnrccRhPe32nzMAzV0Po/hfXjItdCimweeSKhcF
iHaAju+TSF/Wgqr6gHLsmbb7FVSnbh5fnjxZizI8n9bx1L4hzxObO5eXXkFr
IRu5ZCJyyr45uAwLPs8hJzNyNeJLkdFJWcSQBhB/aKrfVhz+JM8eZvAWXht6
BhyCEp2ZKRD9T1F705dZKfeU/UimB/OG1+YTJWDZD8cFw4CXDL3dcabmSV0y
4nVcHZeYikBOkmhTWVKud2RbLKmMf4plXfQKHIj7m6cKHUzE2H+xvv1bKNB9
jkW3ww3oZM9+0KhcaPKlURAnURZN/9fBbWioV1bUBsf584Z/aeDZHYIMQbJ0
BAgCtYalU3adOy6WL2Lp9S6HpcLj9mlwVxPuKqbc9KJm2OP6NvqFiWFcuzh1
+lUdYc2p8BVL3c9WlkPiduyu+1pBfXzs9Sjtij+zvXKVZem7KIRUxmEl6u2X
NmkVood9i9G16tJX9eZmfETDLjLf/OzGmIYh6HckaPzU4DaNG9Ey/rsPVc1Y
I8EblhAwYC0Y8Geco3j/vIIejOhXsTQV/JtdnuaP7plsM38SOY9Ye4KPiyGv
MMYGzOdvBX9+nU9MfTW4mXcaYKQMV82q3VHx8FJP3KoyZgn6D6MjK/e7qgNP
q0z9jMS5BASLRAssCHAPVfPETXjQS0FxWYWJTwLCzM36PG+QB3UVHnT/uE1r
sZMHLt27mDmA0vYq3M1xDkxj8KzX3B+BVPgzMeUBlZh9r/WwrdizY3YW0MPJ
zsATFYiMnTA9AowRRIRqnv9tK6Nej4Ur3KjWfsVj0eJCe9+y8/QFvfCdhGyE
klhgBrvNupk/fGkAZ0KcSBmWEjrNZwg5SCu856PBIwC2UpbsMHx2hftbjdKv
xYh2ynp0K4SgtksJwG4Br+tgfGljANPNwpd6+yzGRwzmtkRmacm0WEm7ra7C
Ugea6SqkBWVXpXnaWdbtqJP41NspJ6WlQZPBXW9MBbNWLKXkvEL9VKOqvHPk
LwB43Lh2xFx1sv32OZHWQwPfyDNydCU/Pw4H0z8Reg5K7quOit0IWC068jDz
b2FwyLU2GHvsYHMofJbNXmuWrZ5tKdNryG2CBsEDmmqbo+L2Oa7i6swVW0WV
qvyLpjRJTm/0CeCARy4a7fcqnq9FfnZsJXIZu9f/NvJFUiah81KZwJ5vxtB8
REaIeHCOE6jLChR7r67zY0Hk6dWriWb5UPOo2y+kkn3FxaBHjPKGCBgxVC18
Fu+ZGxU29eroG8X++HcAkoutORlUBEUQrlaqwUkDf47RgFxQQORX4Dh8F5jE
tcKILK5aFvvKGTpzJamdVk5MF3SmzLVxxjtqYdJ5kHqTzageyOHjlZ2MFwPq
1++MKG2wi+QOIi7MudXJllZRS0Qd5kBKXI8gunDpgCNJ2xD3EwqZn3Ftp2nn
1UNYvdR7kmV5R2SdqHxp7o53yZ0V7RkSXpT/3pUSHWX+yur06KzXe9ZCHkvJ
TIyf/VSeAMSJkxwd94bXeT5VGUcCLwbWI7RTPJSPTMb3qAaxv8zUykEA7Tgp
x5S06iYwT2v2oOmvWAgpGjuzYUGfK7sO2QcqnxUL5TnRJXTKj8uNS64PpE0k
FRs3hMQa3sS2gCUwZfoNxkNPTyaC48lDNRCmmMT7sZkeYghtdfoo1QktuzCG
Te8SPz1dC43QJ12WB2DJXksYpZWGNLD/XYV/g/0UCzfeflm//Wl9PS2/Z38w
P0UZ9MtY7WTIdYkrUoEfPJSA3e1ohUDOh1RDOhRIDizRGXYlFy/4tbQIPJrx
RYKWeFBOECq2i9HaxP+Ah/eHE6SVlf4DfrJqoPCiZ7oJY2ZD9h1+Rl/Einz8
mz7XqJPrYyfCkwNmWNPiIiMti3gt24kUQNBRhyrZdnwKPsWjOzt1f72yN1Zk
nnols4oql7WTKyt5SkLm2Fv9eSPJ+AMDGiaK2T3Tm9I9WOHkEBcx7D6A0wN9
+CcLweQpwlLpzjSDO0NYGR3EIoIH2xSFNSHKWV+kPG+QjnIAexqKeXxKeNeY
+xBnXX7wBTLh8pCDGx+5L4Z2aYyIVuHljBCJ5KmkfST5WEgI0iY2nmuy/NQ6
dY9S1/2oLWDIa0VqJyzBzibNihpBKXSIy9TPP7ATpX5IeTl0ab/dtQS6drXg
F5NfMxUZqI73e+s25NW5etLtNEO8w+ML3tdnKKBDbTmwXnxV20BH4gJHimlr
j3GLE7BO+vn9j/nfkf5gyhsyVfbDfc19UCOyzmm9ykJX+acdQByZeEIhY4wY
qrrsSqrXQTeNwZU0w7OxcTDLp1cdaDtY65bjLBcFqk6NZaKkJSpx+ujw1clH
xEiqNHlAu2uSUFAKoLDplS5Cc5sVOJUtEJwJYOboMAPdMQh798HtAIjw7Od5
B06QYfR7WrcDgJoagrmYSslPsDtDcnoKunFM1WsbY4Df1i0cSk4CMNdiqosF
G613hwthVyzTPc6Hy3NVwx5ULIiNNBkePHsh1aezNEj2g2Dwu2tfDeWz/wDI
IHLu9ZiyBeyaJENNXAL6zewe25ZzxWmoFK99ulHEXCY1b2aLlmEgWKJfJKui
I7UyMV43l8RSs9tSF8Mi+D/JMMtUFKJbshrBRVzijkZ0DHLJSXoCOXLQrwGI
lLKVRWNEn0UMsWNqidxU5fp81RrpBuQeBatN67kE6Wk1vBdcmu8R88sdtL8K
IOZ/4G1MF8NoywKWr+CKGN5pIidhtj/o9kV+amSDB7blbQFR6kW4e8v4x6X9
y3SP6UccR69CCZe3bpyUPF03OTMUDLutFMAzMULvQ2RtSDsN4/uMzS0kPhOg
N4xTQfKF+p0j4RqOXmtcCeSrSKoP6STLN1Sm98Pwup/TPn6wyTYXxNcoz8WA
9tjlPDObP7zGR5kR75ZMf9QgG81EedmRDrqR9XAkgNZiOTQbWUIyP8+lr+Bw
VuQR0wnYs1jrPzP3fn1IPJ/RMwqrEjWDPziGbH9kBlU1O3j1yla+fbnrbGZX
rU8iEpklVZcvn65JdLQh8QFkabXHReav9HlG8WiKM4gWoqrZLh+jaXKsCP/6
NM9KV3/95MuDlsSAtb1yNUIsOaT12XZ3Ko1lqtYUEm2QKPPgXA3RdszbQYgQ
zy8xe+ca+jla7Vn63p2wprY0+TC9YjkJVc0VH6Vgtd45MJ6eGBhqKful+foF
KML5RTOgIabIomajnsjdZOvppe06vW1bwJouexc1DgySAvsfZ3aQ/ktcxtoC
OAbKqzTY09qsifqlI4KwJyVhucyM+tYqcpBUbxqHTLhbn1qszvPSEckE7ty5
qeF5Fow+bv92+PUvv6SNh+i2Z6LVIa29wcKdlSg89+DMDe6P6RwO4vDc6O7X
ySbJKIv0PY2GHqNc02oQ3PQFJK8CYVCJUp2a1PlnvfM60+aqbWQX9fEcFChd
5IvpqlpEFYyc211hJ0rxjWKpKMA0XR8nlxH1lTEZWy7vBxEbpirxADWyIz5w
SU0HKjizbHvzUYI3Eg9ZquiZN+FaP37pBqOPKWy3vdrbLe2bRlRjqvLG4pw6
TO9gWD7QBHVP2pI6r9NB5OqgSl7cw2wKZUwa8zsnfFPOhSWwDtDoR8/ZlCBX
Y4SX5Q+GqYqXg2XlRV3fU3fo0FgjPTEpQv0Y+ughsu9f4AoYqBZut9HL3aoe
MHaYdYdbZYIYfjZ9pamf69EvByL1rWHui3Ze2TpUiGKweuuW2SEK0qTB/3G8
R8J90dbqPk/V+V3mK5os34QNjL87f4+7/9R3PAoUC5czTbkbCR3TykiS3JpD
zyPKB7gR30f0uDfPZjtZrnrTQx2Gwq1W8mzsXxV1m49glQ9ILF4SjduY82k7
Id2cngdX4FvO8V3EudZukoQz3DDG8K5JSad+DPm5RJ6OJLYh7hsrKhjNjzoX
QtQmMhb835g93DTZJ0i4oWMK7nmrLe8xuo8klvOyOg0phm1hmYzJXNHoeHfr
hLyw5se4XVWgSFj8RCjA8DbFFJcrIqgzK1nTbcDIvoZKNwkhB/HYvm02wpv3
l1+2QGmDB8hl7s8R2bR3OTtPSP4UC0QzLGomDv6pJMyVf5X+r5Du/DKVAr0J
SyOzYwvMf7RBOpr6SfYz8nbsvx39S8MqaGRP+o5Y9BD7k+4U11qfg6svg1U7
km6xEKl+Jj54eVnCA8ORbSail+/D0z6L6qdNqQ/+SzsTRyUPcgYAhFuKCdY0
vqD5lQkBcIu5xNs73zCzwZJMzYQ+Y6AfmODz6JyPdmRjpQY7LXghTbanxfAB
jTfs72QquShIssMOMD/Q6H/3Le4okUaRCZraHPydBFZuu8vMI3o9rnTSmjAN
d/+kmR+jpVJJlAnLRZKF6ADGVvV40JUGCqwEY3D6nq2hQkW5SopIOXYqCrua
JzN39JOeHMv+2WokcvUffyceNQDXrn2nyXcvjOgHXpQ6SktavuRoDr9HC4Mz
b7hSDOMqk5nJGlpnGQI+zRLRSAtkFw2HAeY6kPRnE5sOEg4/Oj7OpDYn7kkp
ShjArrFscUau/zJsMY/hFB0zVy9SpJteSyloaAHIJ2dTmTtXK5yDHWyEML7k
0DXyvGZO1jMgtqyW1foB/Cg0DsWJWYsYjd572qxNfQOAHXnp4vcuX14+Wab6
BFrj/SqU+v1yKxraOiXE5uGPL0eRGIqdVSVNig/ANEE5963OpC5515mUlI1X
vaB/ah9A6qfW14ozVE+nuElnGoVeqVpvKVUoeLukzE76tGVMGE+M+YnAuYEK
pC2tvhCIZ42PgwQ0bwKtvRlTTHEMbepRwMr5U2cKNRHWyh2/ZMol2JcfqylN
Q5i0brQdtq0/WYmi2tA2D5RdplrL+ofJCzbJpV7jTCktNoE9Zq7bJc3mMr88
Trv82hk+MzHCwdOdyG2R5/u4paT6Vld0rSIUR+52eZhl9+dd/V7u/XAB0FM5
kpeflIM1OReqHOOINgYUrA9E3o1IjiN6DbPP4MdbDlyUQsFNyVGnldbVOfM8
/r4iXwtdslkX+N6QHTxzuqbJXJwLdJr26YTblEqYGMnXsquAdawX/oRt93fz
WVrPqnPXBuKpfNo8lx3A9V84ye+NRTFikkpD3VkXXB1CG36IwnjTdUGFc6eK
xnZ2SNYSFO2hHIhDmDAq+L3Iznh2z6T9lwbaQhrvBOmusgByA6Ig+RPAcMIz
6g0r9CVOYEkphs/tz+5SBGAUeEhIBV6x9pWeTL+cTLVqTESCn4UTwsi5Onr5
63m4GmNkea9xcGTvIHhP0ffuOYvsvYBPeo7G53iLaNmeiCiHOp3vkR1QoYGs
bcDoe7WhgW5SAoCN+sM5ozivdGU9F2PgOALKIy14v3ji6AGCPQT54QDmx3+x
HniY3tT13zgvN1AcFl7Zwo05QSuxIC5iEJ8x6oLLLFevrRQnCGcSWZbMcrm7
fkpWwuaGBaWXhtD5lSPBdp9sHtxDSVKxtZggUKO4R5ux/3b0HxOahh0vSVKp
jpSfHbIBg0cHPO9T2nXPJ4Na1cXw1kGtm7qdznn9Y9/IE2ju2wRTO3x/lgXA
v16jONlAtJfbKAUH6k4DJCY2IdC0PqyOfh5/0Jok7NqjLcWVgXqFbel1hq6z
f6hfFgeQP/oIGVoJZtrh4mDzqJRQlOq3TgANWfP+jU9KUvg09IQhtD6oCy6C
nBgaOaTt+lx+dEa52o3uo4CPIkmyVaqzdqhw3HM0MbAuBNx7pIuNLbIIBeI1
GyBgN5//SVN93jdTwLvRstE4n14UDPDtY5cjVJoHjE/81aBiHtg3i8X10CyK
PDFyoIXYcp7+04W3Qt6n8Z4AOyWpKDwvx69MDMvJ3TETyO34El6eCcedxM4v
0S1b2w+yaBl0euWCNUqb1gAa0BGI3IURV2taiFh1h/hTRpUyemsl7qIlZ6Wn
p2bvIt5nksW4o45mZQmQjK8CLeJce7MSHeikSd1WfuNM2whPPxhd6Urklu4a
uMm+BZ98CcoTDREKjzpWjG20tKd2/s/kh/iszQAuOKQnwNXa1XkpHJJa0AxW
JeU+Rx/OCrCno5T+6KF7XwkUAmRNoyVUWWMQ0+cXH43iz62EU/ZS2d5Ad/xu
jksESZcQ6uQjir477pONSnx/5qMDcq1996QsXVLeoBVLC2FSrVW/H3uYJupK
s1c7nqqmUXys4OVFKrJUzRtAiowJYbAlp3e53zzvdMaoz5jHawwwD0L6Az20
M/yGM4vgB1rg57A8aIn3WPBXc3YTA4KmIdBIT3wKbHjNfEMoSlj/uFCBVSY6
cuhrL04X08lCicoaQ14zmoEeNSSiNdYw4ZyQx03IzzsVvCgqmis4FuueCdbn
WYwXnpOEQCEYhamvbuG9ld/U5lHmKYAVX/cqSgdDxqSAYIXUO5cOhqilVKim
Qhy7snFcx6Rkk0EUIR00OJfu0jSFgrlpBWEE/KeQQRNkao6JdU0SJUrswDpc
Nrq1w2FelQ+84r6x+Y2ftEvUp6kZkimo8QicsxkGwcsJW/oMDkYbCS1IbhkR
f8TlEAeZl9ozflX8L8rS1ge7dlhWhYKal5+1/X32XjkhsJBsG3+HhidsXIrf
a/BCbFdxOcrV2kemWFRt9v2AEv7CyfSp7ZGGOXmWMldKdmVemeAumXdFPrBY
m5yjzZu+1MTjJS8zeUrRm6MxeoPc4rmfY/8wcfRqZALZ+ib0zZ7Cn4E+mkld
IC/hc0jBMVmeoD+ps83CQIGCG7IVG16wSw9+Demp1SJX3VhyBmnk73Yy9EY5
DK60T9bv7XIwU0EMVqmVJDhbyenA9tmMPmYZmSAYrXZnDTxZRgnQTU04vfb0
+B7uSaa19LHRyc+SXkLa4sR0FWHGMjI82clWxNCdWiJDAmKDomj6lOqGh7fa
85b2B0Jb0oBBvZP4o+K/z8xJ596YjPDsv1vmIFNdTzcxRkYlOZ1jsLovv6/w
j58hN7gEMZ3ZwXra57Iv1KfUlKLCXX4TED1v1toCTv6iQcszfVh5z+nigez9
9iQUq/ibmrDkaQBVOXT6M6oVknyjLAOmDAu7lDzEkTMfBrjI+OXUnWVWfFdg
5GNCqagFm1Z1hE/gOXhEOLaIYNvOhQ7elBx6erVdIibfzeBaTS9WL0bPQXCG
nHpTccR6nV2Y/4Di+J+riO1uetOdUVvriP0kSXxQeRTiaL2bWJSNuOGxVPj8
dncu6urKHQh7Kos8wJEShtTLfBG8/qfueEVINgCcOCJq50vEDHqr803ZpUbu
a72gvVeoJ116sKOpVL2VI1CfzWVo/ONiA5hnk3L5PrYp865V53Q+6SiWW7jZ
xpdqAvXqkhEcmqtvzoB4zP+GHNEXJcnX7ELcZh1/trDANSpET7ThID7KjuWX
2QfYf0k0RweBgnhUBxzf5f6BbXe+fQgz3CPx2oIhPdnyL7qtuIg4x5BbjYPy
0i+PFcZCgsyI6rKDYRQudevJEgw2kqNandZEJTMnL5xFa4HXlgPKHDfHkgBv
uimK8w0Byzj2Zzf4FBBe02yB+mibhv7pB9uSLjfP68s5V8SX69dTB5XMFfs2
U9+TuT4IDelhNGAsFC62CZiR18CXkmnxJiXVtRiNOk1KS0TlBOzu3OnrZtHN
l96aFHacYnrhWZtTkodttFBOMQu7Ug2dFrlXtkZgnGDRs1h8d2y4Rwtyk524
hM+LYr/rP+ywkgIXw8EcqGTPp8NFBU6n1g20P+arl63kICu6G9L2MwfOtcrd
QnWtQVDSVK9TBG+mg/bUyTALZgT8nIcB5ujnG7Og4MkqMpQ2bOCpJmdSTfaF
kf6TuTaE2Rvnk/ch4jR+Rpx0zIy1V29e1QXEJB8sWaGTBvJXsORkWHyMxGFh
gUeXFyGkFli7vPaDALHADB4uUVPrT290zi3ZhVtOmrtWBvH3x3WBdZLB9fpf
fkMf0IiJr47YRi3CCm8tIXc6JWQBcrIM46SLDAmLybY3MY1UmijJ3nxNOGq4
6lFEzUWg1dOAwm3GRPpr+FSpsjsfZpdEpzIO0mHWdUQmXx1H22HDZE+LUtqt
yzNbe6nFYC7xW/y/1TgSHuIBVaSMO8SIXdIOSXQMQrZ1zewud+kZXJ3gYYHO
M+bN77pmUD0Xw2+fHQ3nnj9lfSCXWjhxuAhJoz7wzXyO1HEDIMhJwXmtRl+m
ptgqU2KDN03wB7FTBtInWt/HufWLvzRAttudaVzMjPbTUJS1Fn8BcYeRcVm8
8E2k9JxMpKxjFgqAn9z0bDNAEzi0B1So6sWqrQPLIbMkBrQuX5o6vm9lgNLW
zqf98h9znYASFgwOpAwkT/NdsJ9uQZqlM1ktsehGusRn2sksFg7ocPSah6Ci
aJ4cjLfmfEgwfeAnMGfMC97qqO04QLp7ZXukzSOoYPaP7gLFy4fWJqg7dKoJ
izpxPoMt54XXwN5tsRNTSfB94LXCppEhLwv2ftzz84P8JctyY1YNnChOOVcS
GY8uynwamIh0y1TDGRakwbJBneKH7eow+mSjaTzRVP1qq6vP1KyPF8uDhfEX
z9yW5Q8JKNLNuMBZst88fX+qLEY54z5bxMfDk24H2gUZpB9w79jW80T+fI4h
KDtQbsl6YcEs1lWqcCtzBO4yBn4uLtzEvBwCdLUEVc1lv6CbTKcCVu59KSJW
Morx64+p7tiF9g4uGNVfTfRrTN6SMwOYprdroGUXQesPpVP5cepImjMV1bU8
TXQ7GLXnoBRA+EW/rcDRoMcBQaww3MynvOynu0/AXhelVDw5sh/7VKTPs0QF
PvDF3UBhVyfllzdMJFSALlie/uY2AggVuWOeX2qQA+0aQ7Cr62uCSqDdyQeF
RB1AOBL2NaYceGPSFESX2Q71RnSWjVX2mCc0BlGWBj/CZyHmLzhuiSlI6xXb
O84s4d/M091PyODTIc0X03R+SVpJot5ci8fRJlKoxNPUSKjkne6h+Zj2uXmP
iS7PA7crmFlnZHnBpFjFzG4U+qC7v9vm6cc9XNx12zXeM1e+1435YlH5G1jH
kjPsmCV7mKu8dwkcz6m9yfvFaoCY1QcePLN6fLTwup2nAZaJJNym9g/nxPTI
oYTA0VslWKj7u2Rta7TtLXisdZfKD/xbTRRW18Vaio0yjkziksIB8/2G1imv
YDon+FnfckFc4JlwMxlnPpDdHPg1T96css6sph8xMrqqhN+fybHyWkL5D4Lv
bDD/GXN++QxpnkUnLMw3syZzUfvuygvUlodhTPNF3Ikm9zAR2+KxGF65lQSa
pXZvoHQTWQ0enx25ZDVlOGlLACbX7lzUN4lDZh5K2Fz3Uu2Y4I0268W+YjLk
col2Sr+m0jihJSxG69xe25zZVZpSoUMqST1RHGcUsJWCZB0N+JZoI7ZaO1XE
8ZYehZs368yWUbZzXG2HYw4SZdZsM9a9JkQ1vIgcF3YU3f6s1cN9ZN+SeFWi
HHr3Sgw1u/iL2ZecUwKuffniOs5XZCRhlMGbLnI6w6Ku7c9U2Rn9rRvdEyb0
eAgQumF+6LuccC90AbJcPcr3s/+sL0A0icbIj8TQIdLpcus58p0C31/bFB0f
CyjA8gmGsLUlG4Ic2WWntY2HU0cQhcoQro4eDaxUMsdSRbwhLyKxsiCtN5Am
YggXUamZ6+UUQbChf6pVafrKj8G/7PsRiD9/cwpWD8o+GKbiU3Fi6AOzrzm3
3ohoutGCw+GnWmUmg2li6YGA9M3YOv4P+XEHJbfaBP28XtuY4vCKqcCqNrfy
WroQL9wxYRle/vOAX2H9Jx6UABvhAea1p59wMFlGBkCDLbNAHMni6e43gtRO
nQbT5WPeT8dpXN0eAx0MM3peC4JKdIjANNPrXzYq1DNWfb8eTDy50nT6QC1r
iXEHUGCWIEx0MldqcxIEmgg2UMfu7oW5jDuR2+Y1VBKk5QtlvgZI/EG0sBue
zuPWrcoxxW/N4xuXFZXvsUfRlLs1QWiPU/6lea1oedeHj1bsjowHrH2uRdQp
FXDhjlbC41HeLNIsSu95peYhyrtSOOdLPRUfYmbZg21AboTGdufkszV2tpUQ
jseMerQETGgK4KiZUsdieuhyqZWQPxcnC5Tz1+IVsyRuxb1xteUBgxswHwgA
jHe048djBDLSzb20vMiGDGiP3X+5oJ1HFRpz64FpfMVwfklt+v8NSxV+u7Pj
ZLrvSHJZHO0njOWnQoFK/5prPCYaghIdjqCjkBiXjV0QjrjNxYb/7Pxx0a8a
dPcugyysZstuC9rvigxqDAlCaEoAtQilwUtyl1rFzD/d2EVVfFtgQG8cJUz6
ILImqVMfTnMlJeyBFyuiM3V25L23MGaaTSWgLOyvbwY8geEpzkl7l9LrUNZ0
cs9ernm8+Nh0+9iGcEMvFImF308X3W4yRq2+GaxCvsKoPGzbzA/OfQh3v17x
xxqGr6gMp2Fw5TbbILQUQWlhweMpTVSgNmK9iP7DN4xpbqERIjh/38cyIBCQ
NB3QKo+RGnAXZDA1/dhANBbnet+5VGVrN1xQgY/k0PlgSvqPg3+g9NkCakbB
UnfoQF8FkZo6u5qrRrYhanR2AfreJ0V4RAEH00DPgcWZoIEJZ7CmEhM8WN5l
rdl5woLL0AZ1zhk8bBj7aRgNOFVF8YPtudVf4ncuQLHFxAfg636T05m/2a95
3qKD6OL0V/yIGJqEI+LVFeyZwbeIG7wqwGqTnRF/gLbC/UFh9e3kzB0LaDrD
3NFdoU+cuA5T4Ut+qg9fZAl1xJ2DfL1oEiWkePWYSdA7L0LJNYT9umuOIzdP
aunSf0/yKm0kJk/MxylggkqUzpzUaeGD/JTGkUUa2gUCegGPztbC8hJeReGt
7JmIwddsm1l+dUkBteExg+CdRsxL14/sb5UYF1hHYBHsPlwOzyNNnyrUGlzs
FQy7KC+gyYhtiuCNA6tbdgrOpykA/Xsd3QxL70UiecNlipR0C9q9dyuMKiB2
gfGMm8a0NR2zOufhRKzjXd51iLXP9qToA3mCbQF5zHBsrw64I3EP6TF8SS6l
3nD/e3KLQwJ9hXsuzRpK0pd0md2sbOs4qqwp4Tym+0njByC01Q4LCevGl9CY
LIkYPJOKmRKhiS0TcmidvlsK4n1V83jkjE5P/V8ECpCSzZ/Pi5rqvzxAgI5N
sPpR5AJ/Lq8oqPLENIQDLyLckhWfhnMCBgRhSNidVV8VrmUD8trHr5VNm8CD
elXHWquRTrAnyx94vQJSk7SfOYcpFu9rJR0kVZXCQErbwArSdrq6J4xH2LE0
1hP9DNQf0eH8g9bLeOnF/dpRvPvCMFRTJwBq4MjE65VdllGTjks+d4EvTH5B
Uk+Nt6nQRZIAso0f9d70y/4oy/g3QaQM866m1gGZCADdPiT6BJBvLzbQrtOn
V2M01K0rqnhFuvzS873Nm0R6+klVG0xU94JYY4en8wJOz2tCAyHsvLBKTU3a
H20rF/shZMi2kbk6rcijBarCvG32Rsg36ng6OHsyZMGW4tXTQeS20oWiInrU
1qsZQtvlG5JrY/8Pi7njrSse3j500FmDhfnVlkWsZWCzLnovC50dtrwLogvC
o7hXLyU7ZkaG4u/BQvLpJa511zasvPBMG9IO18bmSKFsEMrYon6UsKAEPsjv
igT6qH8isUrvzDemwb0+OfPX7i4FbwUyzAgHzBEp7HcnqvDP6WKQYpeNuYMO
Uxb8ZPclbClp5ZhRfoFBKJxmte+l+C5XxpstbLidVLUTpsM9eniDvFI48N6t
ACnudFWeRWzf4wlfIAaLbQW42Fgk3XtmOm2dP5Arxw1XgR27y4sCZFzxUzHy
3T5r9e9tu5tIo3KCOLhmHwB8O0Vbz7QQojh1r1zx9G1d45vUyLhR4H1ozr7r
t6hnVXNutzLe7OuqdcT+RNXc+R/AMKwmXYKhXTKjrFyRZV8QjYy4X60ctwCg
Y2ZN0/3UhoO2dicEtqY4OwnKaa3A6ObquofkD7BM+LOgQ25pZbAfGeZtqwFT
YGEay6UeRMwxzSKBoNWz8hRoJde2QDiJnB+kihN7JEUrH+wLlF7JQjKwV2Pw
AFx2BQB6bhQ1n7UYeu5kQ6/SvqIiLBCG3rDWpEYMkJI6o/ghJZxnna/dq0se
zsmwW2KZcEonCdRBi9sN2rr2bGH954SseZx7NYBbBW0WXWuyZjJd30sg4W2V
BpQXmg1zigExhNNoQTTg5BRccyWXPcQ71psmaeQbwNoWCubHUTbwUJ8jT6NY
HY8EdhSEJZdM2NGXSIwQFOuSm4W+Y+XZezetrRiSUZdv4chSdg9dm7Zn47Rb
wllkvSiwsic5aCF6BDRp+Ly+EyJRtwbsVrg/ETpPlZk8o5rouLsmPFX31/Cm
OAwA0PUN/ph7fZPTbqa5ybZN0gUbqFpgIoptUZoqZdEVhDP2K8fUJvkJ+3TA
cNwb9gYjrb6Mux6j/9rvodomlKdCkwbXSYaW/ecDL/lGb93/h5AuCX6tDQ7r
UPfXYWwFkot046DG+oz9Ryy25W4G+5RtJtn1wBUxz5Han+a0fz8ghK9bafjA
I62smxJOAnm6ZP5mLZmcZdyFJz8NMRrYnHAAhz95e2Gn5bLAEYUb66XcLwWa
JDqhflZqFNRbvqH0PXOmlc1bm8c3qmEO4iHHOaaupuYVKOIXvS8voahC1lsU
LEoVHXBjfjEhTt08jMTB8MlDTZW4dt4itI7nCd9OChzdVFBzUG1sYY0VZqex
ZEJLIoo5IAe5kKNac58stiDaQdtKQGS+957ymRP0Pm24tS5IPRHqWan5sBrB
2FNTwNvEzMBzLXWMD0hwQniDomhKRiyfo4gLrGbuI451Tx+R0C8D8kRvZ3pl
cn4ANntym/MqZXojLfSF7JZQ6lgyA8dNogSu6Xfnu+FuWQW3+fsyC238SFQB
HEhnliJYyWOu8qPnFD+6rcBvsmDlBt5GJnstJ+8LSHEWnJIelUE9yxAYTpLm
dj4doWXaNcKaLqU0gMYTy302lUJi2Okj36zaNrs08vyTnF6ilXQC9GGZRFGz
bdpgLrMIOCiPwU6DElGV/ZA80eqwWivuRLE3sucEEgVxQO1BHLdkaXrO8pgN
3qryTy+F90JnD3ZoHejIyD8GzQzZPiW5weZ/SmPHn/Uv8GTWkJFTqT9cHpxQ
Oe3SxxNF8v92tV7KTvdK0U5NhTyfaInhz0k=

`pragma protect end_protected
