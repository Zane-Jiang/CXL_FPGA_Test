`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
occubqmOff0HS7vTgg8k2Z/Nnk/jc3MUra3+SFbhYVJBT55HihmjvK3XOD1zhTH5
gCVARfghcUxpO9riA21RAr+uKienrUa00cxJGCMZegASHdHiHPWmS8BQ1i/NFodM
PV9ykTePa5ab+4ha0YTw3QmIB1pwy++vB/wLUGdTECI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 57744), data_block
kYq5CZuzY+uk5dI26LWf0WARlb3M7n1MiK1u9vGNGhEP30B05DrnEdAJ3jRltU4+
Y913DqKPhfhAbat8oO1twi/Qv6IGiFiPLqaShU6OwbbQ4h/UCgGT639gVy6BH9XL
YKB6LFGh9t5gWKAHSmUe2l64n/vWpMgDF61HYbAajeyRJPSs0q3bFQyjk7GxdVFX
MRN+CQLV94FoenQzK2j2dxH066iDRlO14Ql/Dj6wq1en7SR70y7cLX3t1i7DNXEK
Fvbso9XELNq7q7QtVOW+EwyX1fR3y/IyIvaNO1G8Di1O4pwAyrV+3mFFdHxz7tor
NA0219iHoYwAglCplv60XSU2ao0G8vjaoxT8X7gywDY/hgjcfmQPi/nIy2ot7KbE
HJ5ggtFwACP6xlP/AyprX5pj+bJNoyoR3EoPcePU+b+UdgIRpIJ9xAmINFog92S3
G/GjpAA2g6hwe472yLaqPLnTWjnyYOF19njcVubOWyMoJK+AJ6QDhSBgTiawZ5/y
WEsxj9RzMbALSwMA78z3YZnx1OF2r8nUf2ZR3/UWLUbMDKLxPyQDWP9WSBMOVdj5
FKVwfBmcydAOo96bGsJ+/kROmEU9umb2SQIBUKl95rF+lki68/2fTtAi2xlr6hon
4nAscFujQCe8YzjCxrZXPwh2vTs9CVmnZMMJ2KXXajwBmlKizhjGkvDn1xeDdwl+
GUo+xcvXgkmbmC+z1tuqhb1dj0L0gxgG5IxLtpEZ+PBGtZoPHmtQ4rvg3IX5/8zm
RsFlBvycl4zmBv8GD0r1B575U4KFgygVp7ZP5AA/gTnpRoeVD3arQgItkj6WbnN/
Qggw1L99Z9Q6t95ODVAzIpIZyQ6GwStdxjfT+zwbTBF7Vb+He/4BgCT2T0dED4yK
NjYMn+lHVdoyOsTQgmk6s81CpusfoE0uBxfzT4tXZ96nXlJIFejxpZ7COWvvIu0M
4CrrjY/f30GIMRNKPpJapu1rA4d/IM/JhK73FfKmzca//0HmIQrpeFoCYUpdWBfP
d8bw655WSDcdU7uNz//vKrWhCCRtnxiwgCCCjiegKcevFagOnqZaruUMAIMfSNOx
jHCFuSZJvtqvC3BD4nSIxlT7fzNGOMDmLSeN1nV0U5KbI/2sidOYN+/l5eG9m8eI
myJcnnVkoDvO2Mh9CpoJ/q+XQNZz61tuWUcuMf93QdZ7cRoAN3XaVcA0qNj5wEbr
YQeT4z4u9/EQE1EWpiW1AaM97agPxRj1MEdESAXb0BaZSPTsnSeKE/aRTKIN3RUs
DE5K9KQDlzdJKj4cBrrwcWKlkrbZYAdKJLVAl457pQG1oj4bSjRaS4XPWLlhDALW
7BmmCteRhnJXI7/Ur6IaYUciu9GYWmE05S8f5abU7TVOGWbjSXNuDCA0nXSrVNdI
IcjIyXvaDSk9SUKKHEybQwFeLYPdgiZC886kAjSDV0yLyyM9oJQFFdlLyaKMb/ER
iFtIuXSfKBFBxJ93gWNtHzsDaiOvGO/JWHFFYJtiEoR1kk5wedkP7gfm6MhBsaOH
a1Qr48hmPhcHmAFL/hEAxSTN1ZnRhVkTw0dtLz40EG6Y0MoHM4qCdxQUzMFQuH8s
Q92/a/+EaSWz+NnRGkeqxWbmpUaDQHQIgyxtoVH4H0rRZt07tGwOrmdtNsiwvZOR
g/O7ZEwc+/aTpDRnU24gqJDFPf6dAF7tsRqfxqOKFvGhmlfS0PjUKo6p1Mtc0oKB
6w+XLXDlHjtYRriuUf+jE+wMl98lG8u9sDzupUpaUpdQAlYhSOT+4/CMEoTbJVl/
61Kkk7sm84mqvTtQzpZBOrz+SAvfg5mEIUXdnao6EQdZ4ct2zjd1fk8jsZGai40q
IptpkYTeMZfkm3GgrZ72qGG5j1LOoeM6GgTbTg0gbZnoGdg57OBxlTa085BykKWK
DNFXy93QWntoT7iDnkAmTvqOi74SzDpkhyWotM+27juZYLW4KsjZVsvaZEKF1jBS
Rn9jdZohuSNMzAWt2u+7XlXoscFBoryQugGw+gPMEqfPpm8oURc4EiLsHHphKbH2
KCU0Sxco/QUhxbK/QWt0xBNLOh9QnKcRJvo2YKOyD2fZ5e0ZATcxF6eesHToYpEJ
s5AsANH3oPZvgpwq98YTetYnpviVVr3cNgYrSltYn5wuDpBj5xVaNiGfMQzimiqw
QjG9L8TdztBVFwy9uE+4w6h7iiP/8zEXHccvDlHCiP3RSGsYkLGZfx20k6cHaJW1
X6Vo8BFRV20wUiPRYwzgaFq1Gr2PF/D0JpvPW5p9Cv0s5Jwj7GdgA/Wu2+ZIa8x4
nYURnj5XN2zOsTGhjLMOyjRbOTGnQzCBBqIt/NJvZw2qwIA/Fn1Jd5NoeZthnv/7
tKGscYiA0QXygFLKoEtCy5G8xMU8ZWGddnHO4kSP04I5YjRFSjXmTsyxpT7rfdQI
+paGqsX9VSmW8kfb+UCGcutWHZTSwucn8Mj1XmyfHexVs+GnJH9bdE9XDb3nco8e
P2RhenItW9hVr20lSpFeqPVtfmfzOkSnpO/Xwib43U9ghFOWKdUVsnAbKHSAB9kq
X8tR7Gf+SW716Ef0Os/CvsTrS4qniVQnFigHzymLUL0XccxgTlORVOKRaq1UbBUv
09uElUkQ+DboahGE35rUhbtPf7aw415IomQAkbibqXCjzwIEBxjo2XMPE7DtjjZu
k571kF4N8wTlffmEpDhHhyN4MVIx8HIHJK86Flnge1PYjfKaOu5+4VDa/u1KqBEo
Helzo6el9zz1v9xQeGZ4PT2AdT1vZ5aXtdqTjzrLnyQl+E4gDNRds7EJtX+S42h3
/KZvLADk/XTSmtPkAObZKZPDe+kIHA+2nzPAuz24ZBaHbRnpv8wpgU1DUbknpAUI
tvboF04RmrFWQ054LzMcv2RUDXW1SbV+Pg/zCsGsAdX6D26powDcXbXvVbyleNp9
TB/e/8S1uuPB7GWZJaAuEqNFDampJyMU7ZXH8LBkTaRgLXnTvlk2OdGWziGsmm7c
dop0GNNDYi6i5SRIIRalub1Dc79AtWA6/qZDWUaywK232APeJRZ/BphBq/8tTaml
RNGZabqR1ubXOzxbd60L9rR2K75vD6R+HYI5purOWw8fL5Gp8NaWSnQ3h69pqUrt
dsr14BHRYLFL+32fb9ZTlmXg9HSCowJjvpQESTeQqLBZj8UMnrED8KKn735YB6lg
fwhZ9oUJ/UD1N86Eq4bo0I7/1R2lUQZrK+vXJqQ07YFw+C9grNI0ZI8GUX/mWDme
fq0oTbO7EAErXs7HmphwMOTT7+3iva2JgzKN/pVpGWfdJB5MKYJaLq+AhD+58701
OjDP0KeMECAMWzB8GSkPrYXEi0L5zUwrZ6G3TPNum8UPkoxWglqXFYpYc6+MOYLQ
/T/Jj+N4ywnqJC8/JIKKgak42+qzibXvb67F8GU/hcx4VIOhyuzmRLX8UsmpzYZU
4Url0Bnq9ibwGQ58lehRCWYcSMUOQ1Q6Vt8DAhejCLEcRlx0cGGqs/1jchr87U9c
pIH7gCsP7FOb4WrxR4YDlU7+316PpML2EN8V1SJyQAo0nLLUXa20IUtC6cOHF1SX
Yckuv4k0XBw4pLV4wmcU/TcXBZbOImeW0ytU0DLWy82/VRei+DhPpdpj0XubZpSv
5Yh42xB9HKQqgNJp3ZsxOBzjFFjxCOyJOHhxUJG+5GO1/RDewI9P0ZDwdd0AS1U2
1ezLB0qS/zPNQtcehHrsPl3sbi8CgfJwcQGVuHsYboBmZBFkkZbThyJqREOsQiKQ
zqxpVsK8k4fXjmWamsu8YwzXSps6rTB+aClPj2POyqqb3g2fZKb2bzG90bngEFOH
iaRMoaAFUHFHNZnjv3aWwxyi22z/OkUobC7CX5XX4mTaZCZdQaPawHe6wAq1bwSd
xjTi1jomC4vLJqRwrdgWe6Fidrri67z82FVdIOZjcVCPzkJeA25zkUAqvCiIdxYZ
P76iLWyC3fWpPhJbVBxroTarjjBSBZV3WlpaRtTQLoxEU6Eg6FcsBZbNFceMavT6
FQ87lTeE0PveowfeUukvrwEebNy9t/agrnwcdJqFhjt//i/PfLfnw+5h9YWzqfMp
y2H6txpUE05+ptfrA3HQ7X93Fb9qf9ueZ8Zg4kPdpmW74pRb70O8hE06R4eCWYRv
WfUKZHB+1xI2x6hFRUyLEaLTyZAKI7FEFmSKkzwADT5sGSBe5DPhtMzBWuqNKoFY
Bv56FqTUbnfYMd2Jl4jcE31mqltxcAvpM0db+DF8wY0ympPF8wa28t0uNkNrKQEX
G59DfsxLO2uGVFYaPIZTEpU4XUR0DrafAfa3jvvBttD7uDtizaoREfTZGZIAL7lo
6SRQDg8lOy+16C5f6GDQCOdMyjhXSraT/f72yWBalOiTY48CL7q4H9qMRv4RdXUk
tbYDxmJn0hzjtYKaQx0lZ6rgkQBvgC9iEgfq3oscr7PRsosHIVDhWREuJ6vgOQOy
bb+qd/TausOcCZ4r51q7AZYOGHdtdwI2cJo9DmI45o6QdvHXvIYumXvuO4QXvds4
GQ8X6zkbDI8J8LmZHCz+O1FN/U/pz0jetTEl9lwIxk5j7eB/KRNwc1Ex/6+d8JYJ
/Psy9O6tAt+OR9P0JTF6FdkuktKwq0jqQ1x34gnU5cGbIITFnmDTzfsp9/ncryJt
9dQSk2Jp3L9XpKNtS1ugt92vlucUtaQ/vsEQ6k4rT4VNi/lQ3WmjLbT841NJqdCe
zu/SivCGxBL4MdcQP+92CL81P2y0y4JRg5A6sb33hyoaHxVA/hicjrTIXB3u+Y6d
K8z/6XPgjzSABnCxQsasffQ9ZGwiZXAPKe2S6kKI+pk0saFMwVNPk2y2q6HPhN5D
g9U880ab3mKkdiqt3ILi5VJyfQnT1YDDtbD/cJ1aS1yGOiz6335N9E1bYR2ghzus
EoAG/Learww6TzTqOkdwOQjLtHpOGNJj099WUoAdNLufpOyAnmpp1LyQq8mnNtec
As99+qwh8BsFdmUg8ZdNtZGzorukq7Y/IGlbz2aW0tVHXH2gtSiru3DkvmtFupwm
7GpcCI3/j+Ixx3TCOM+OVjpM3uL3tcCHAmV1M/oAPGEQVibx1Y73jWvK8/s6kHpa
V7bW2Bme29Yz8qe2KAavDpRaiNSaT0WcFaVVgCKHfpydKDp0yPCCfwNYsY5mpRmm
H3Vs4wVDjPcUQ383h7rP385lhNhcZKOBJxRL8LEgZa74CqVqN23vIsLvRIlZBowU
+ZkeTmnTCaY56rnB6XDMSNYUP+7DbNqZgwo1Yp8m9NLdoR5hpHzGBlTkyLGKmT7a
4Zh4gplvIlVyGJ/EUGtVf22uiBXyoiK0FlEzEyxxl9U6vOH4ihCil/y8aVjRtDNF
H35aTpuYum6dZDOXeTfSo7EDXjhR1vE8B5syl5fOhvbNwsgycW4MAesHXQxJJTqZ
kHnph4AXvz17iqgaUdiyla0KfNTHHLwheLwIvkyd/jy4Vm8W6NRtZZU8YHY7Bl4d
J221j32D2wlyRlLbXemZx57MxImnuiCfzJIpfx5JDgOZzC2OILB218ed+JjYeq8d
g455/zgiM5M3/abM6YYgpZ+RZRyaFWNeJdyCMob5wE9b70tL8XQ6Ey3NqwY51iZV
Lx8L9i2s+e31dTMDS+tBmLdJKk8Nk870nz/ySmWYD2je10HYLeTeDHsPcjZWtrgu
74iOpSaGJ3di0ledFJWwoXJHyyHuMMNb4m92Da+lJJb3MaUl0i8twcnfAnOQEWr5
MxHUWlkF0EKHSll436vI0ZynMQB+M3uRFtIEZammoF7nFQo9gEyXeA6BOCNf94+e
UJcJO8xmbwWWQ68szCOEuZCBMrpoCWAD00DVMcvZn+VdUzgVmwlDv/mYbvUgBb9T
t183azkWmP0AGgKSKYWolwnN3J/9wvLy8kfclLbmRBFETgtEWV40FMMwKdK/2hvF
0L2aSZ11N/gtZMxwbzmPOX0+v2C8mg9vQ/cBdXvBEBxfYH41RsV7OUtg0RSH2kvP
QCNXvzjFKYgUcDFWJ2fp5yqYY/Jn7yLM+Yz6aCuqjt9TidgjDxsPA2uLpgpaQNwg
Ew6H/dsbCprF9K9qsxgEa+ODh8Ui5VIx0sMjA6E7TYYg0ksA3FXsgL1nc0d1rq7c
cUfLpHiCxjgTNG2r3jhWZV0uSrQzufhtNa+Si1qoVOYaeY5ADbHSCqLHMPbvyoHr
5QxsLQ+JTv2qhYwxUoS81deRK5EYxvYzC+bCO4X0r73WwlZmjiAUUn1gTgIuIpmj
aK1nbTx/o/44HgsQtxOoKnmBet8VQz8oE3RIYsQXXAIbzuYEGYO31mGcifzpw7KK
uQk3tYCV5w0bqSvK77z+s4TzZlkKCco0q4PGNlyc5e1PExSLNJuPNFefDXTN1hYN
C/2UauP/oE0Xm+z9l28p0+z+5+A21o8c1ioRHzCDMgVtNjWTklDziH9DFCkbY0v9
8yjWIysHeaCru3FM8cPTVBgOfU0wtLMX/SaWwXLfXK2/lho+Y/NcDyXMBFdMu75c
ZLMpG0P5BBaMVIOwRZbGNWN61/Ssad/BW6ruQvk5p2vWyNY72vwiFRku//2ibE7p
tq/4JLboV2hP2IQbdVApShjZxS/M81eEK2A/QG7Fo8gPkAeOeDyjzRGt7rTie/nB
spTsnwvOrKrt52q2C1C0YL2PaBmhCMgJv1D9qwVZP8Xk5z6pLzxYJkXk9qj18Mim
azXnIImL2KdwTI/eDxFhctSFysjbCaEgfGReahxicK/waq3ZNMpvPpN523MF5IKT
Ohpo85gXbEB8lYy4DUbVCmCP94VLqgr5usqieXpnveQq7m7z7R5gxrVJJL2FrSuK
KLuR4uJF8jqR3sq5cFi5JSQOy5jBbtBOO4xB4tq5tyz1RIhvv+YvP/Jj3lPPfBfV
Vk5ZBYIuBflIYnSwV+OLdX1gKsBkO5RnMRxiQhJryK8JZln3WjYn9rV8kE2YImv6
rHbCoixLNdFaROlqQXMVTUlQZGIX2jK67lzw4OlqPHoxEtD4DVQlwZ/7+AP2xpfZ
2KSP6D38KnEpnBrwRyadnRNplzQzPLKp2P6X5mq/jDzcb3ff59hygMf2gWQLncgQ
J/AyRC0MioR9GOrr9oDo3lK7JEzvfWflkih8hMwLCqvCOhazo3G4pwuZvrAAEMtA
sydRAiMygPsyReBQBV8HlH7MjVduuL6bJkCulWSmtpWSfLHcO7kddziDVIovwZUA
f8+TUz+A6F52uJD7GLwdJqkd5CquH7ihCyURzzMFk5BRBZp+StnTHkDL8Y0H2Lmi
DsTcjbglRY1wtAS/8nvMzv+FjaAkgs/PYCdz09EtwcTFR6X2jiH8uJp/znz6znpV
c2Qm5P4Ei5j5YQ1UFkPm11OnRTK55AVeG2511ACakGDIQkWDWqSaB9nOuWIJj2GL
Ec2JmUBeE7rmiWenSrzra2K4qNVBFViOxSdjS4UH8dIyxeiWTv9CqfceiLMwZwDU
zyLCGuEtY/eo+DZHGLG6IQqmv8Vf5LWoeoeKBgHuq4NvT170iPeR62iBapY+PW6x
DaJ2y9D1upRZTORFT/R2YteGqlYmOVko6Yxfi52oaPOYKFENu5ObYOC6oJoWIwaL
eFPeHbdwX7AMmDp2eu8jDT8ZMbFvPCVVXvNpCMEvYsBDv5tm9owbsEgEepYqWHQ+
UJXTL+4IJjNnUSU3nZDScMTW0K6EqGdfC84QISYsTvoboY3kpy9TkxOUBH427AIu
6NPWc0n3E6BSy5oJOTy0GPFg90/svTA7mmnUMr5pUJ0/00Ul7ZF9dOftbPJ7JXvy
+XPBbPQQ5LfyuZLdTm/gt2n+65d75yTPemTIPA9g+7YK1Ztg8dUljVannbGvUYcX
l350BZ2C9qI4zdGVgnQ7VpQFpe6psJmy9sD8g7ejED5i2/isWjv5exckGI6fvufn
Gde8h/UBcMheGSeiozChdPpq5bY6rrkdhG0vFQ9geMwsp7HaWJvpO/kQo8j4E/tP
r+CObVCO4GkrBG+5s2TnI7X7G61Lf70J8xg9c0Q1l4kLanAZqcL/x/9lpDkXXDEd
p6wWlSUruHXtMwO6I4h/8n2Fi3BD+kNXvoDzvDHoK667ATaQUFSdES/eh5OM8F9Y
me2NLCSrmK79+nbOBw0MQJTKWeKyN2EmN2i60OW9gckCgMcvYVACf3Mj3au0KK96
yMs6e+pLMJkT0TtWyxgy4h1A2o7IcyURcZ/EPgDln3oiulcajdto/VYFi6omPHd2
IH+XtVfWkzgkZF7kVyJaJGayVkXZyF7HmXZ5CMrDTXCAfWhXerwg1dOQShl0e9UZ
lJLoPMafhlD1DtiHEO4Uv22O0HtCXmGfqNLcesfsLCzuEdch+e9UAiclSwlz3g8w
4JMwlzYFC2lZ7eHS/11qtUGVeKlE72qbboiPdIPuDrQzcQ67cErSCPaXQ2r0yaJ0
fViJFKIAVltvB2PzOge5GvBccfXB1d00WOx+E2HT5Vd4tdmE9ARrKsCjoc/YWxh/
RBsrAJ+5S9OwnpX2iA4p4blqOASetmM0+A3f0gUco/0IZNVQN36ZgCcCQBdlBNWd
AmzPSOIuyk8NLX3qRh0lZbTkODH4AJ1oHngbOCWyNQ+eGkAay8mGqZIhm6pdqxiS
LPmkKpd3Qf5oPsZcEyR93Ydcfexh0NHIlA9FwCrZV8tC5kQ1bRJrZV5BaqnmOaX9
e03vgVoG9V+eMJmu8dGVqN5uGJngOEVvjni3HlvfeFTkvFRuwm3nsIJZqHl/PbAP
l7e2KzwLwMc0I3w1LwyqkhDPZ55P800OOtpN3+XQJX16wNzv2BRxxG+Tm41vPwnq
A6cN6Rqyk35yAIEZjcITzqPeHa1+79gOccN6PRwiEdHUEoMakNeV9jrOdruKvf7S
VqFQx/Uw3wiXlqYwxmP/XWjLZZ3Mnp9CqgPlBa+4h5WbKfvEIbU8MK4yfcFfApN9
TOFmUf7zZMLtf5TQKvwA6WwCSpj6fdPqZViYmzW59DfWUqn8tZMF6qWsjPArdt80
H8NgCWJ+YRGYrrjS8JtdoVpLy2CDrkAPVSzUeOw5KRUpnp+tdA2ZGWz7uszTPEwQ
G5C6MyFOsAyzfCmY3KZOGqwj2ltABtHBdeMhWHDq4EA7ncH5PtjFMGFL8jsRueTw
LDcqJoPW9lH6p/UEDdYfXmoKqcP2Ry6myWz91MBa/6LoncrMgoG7RbhQmeYdnHzt
j8AxVCKfgESvUWEDgCjqNPS0rePTDKuTW9y/DFLFHsApZAMmgdKg6jPt/pmcpmJD
sfkisg/LJPVMnXf6/jJPy99/RPUS1iCuijBmd/AS5H4/kSD3mkO9wFChNQZlWfJC
S/Ajfb1HOTnGgIyqBFQQke0FvbedLybe9STUy7+vjl4MB0K0cK7jOuNwd5L1FrvL
LIDpEY+pnGhI+ztM2cXYRuehtMg7j3spVdFy1GoiXpJ7ZZDcOFN1iAKBiG3u9vTy
iIi8JZpWjYP/uy4mXB6bev4JWUkuwF+UnvMnVGYhyQGm/+6Z8ueGSMDwyxgPpYZv
BDEWGGh0hx2Y62VVrTkMG+jJB9fpmuWvUjTG8qj0YNQZZ1hSj6By3fL55O6dkFzS
w0pDrQx3PYschLT6sNarwXiSmIgKceJBz1piniyrao+eJ5pcNoYlVnyVwgM1ljRD
VQYt7BU49PXifAXP6R3sTt+DcdbtxNQE7UfcIn0F+48oB+N6b4HseuFqUZcVBkon
hC7AZL4ZqtXUIfzrcFVcgQ4IE2w9o1JVb4mHSjj3skFFjlOVDMXATK1Abm/Yzyc9
ZlZu5PwY3q0FFK06vVU2M1rvP1HJzegsp6uMf1QrZyG4bnDrtEkt/Jw+I37DJajj
cr0VG3GbIX+jAdFY3dw5FPjTOKo6LL0WMYh+bC8cFdtu+zhBQk7BRR8lUBCTfJ+w
5O2ASanCTPHPnd5DMMSNOlvRV4PWfqjZ+7Lz4oiIDfAE+aJYJa0MVZiac/S/g+Vp
syOhwRVn5qNH7CzkyIvxMv6JBSdb9jK31AnaMrOj41/nU8c29TZkBuxOH7q5HsWt
tczS1KTIxCindAGCSzSc2hV0zdZBQ+cc/+Wz/zXz0UtisgbA2Naz/8i8A8JcUkWz
wRZ0IokKd4Dl+JhrNthl/WUwYDJafHCDa/wuqxP3r0Llsy2HIh6aZ9Qnf5jXhY3a
TV5DuYRwRhqY70ygOed9MAFMSYYrYPR5XCsLWwB0j8e/20V5gQ+iClp68DaHyqUE
0mUfRNScpXymiFym09WvJdLvOvQ4s+lGAfxV0TvdQjn0lFGTVopttTHlrzm7vmDR
Y8Hqav5YUzdaGBs9XH5AQfhKXw+8UqjgREB6LeokUnxBoUZkqshp3SEqYqpzQCrr
DnE51oE51gJ26AFG4/uoZXbuy3IGUOAdhyMxHkspO7AfNnWZaWikLVAJI/ZoPjku
IYpuolx1uYJSzQH31tIVtBqvL1Fmzvima9wag9+GaH96hUabMaQlOsUL+tYKtvql
htA9cQVU+d0v+k8fL66xFyqqX8EdamGOt4Uj6NKgBC1jrPr1LwYI7tdQLcWzLSOT
CJ2vkAPHcJ7tXBJGp9lL/b2Jfz3Ftt2brCrhqUK4Ytas2ylMn3HezSlFi/Rdqxrr
N8VD39tMOMa/YgJdSEpJwRF/kq3FmJLFmSZ8p+aH8KMiBiydAX87CMj+a9DvgjHx
TrIFaXhRXGcDWBfLgNfzjB6Nggu+cKk3r9Ob5oBnifh7JBAJLLfLgbiYEhsWQv7S
CXDjh6QGGEZagI+gT1CUt+IcPVDl9HOphQ2eAxkRn5rwzU/cgJkL0A86Zl/Akbqd
YWYNXlIDMphF3FMBHQp+tmrR02tBh7W0umq7JpmnCzIX367+HH5ua4QhuW148IQ/
Rc4dVsc7HEeqk3388hEWE1VmPqRfNfI/o/QFIzOHOLdsM2pBUHvJCiRwwNdYdy2/
sKuBwazIvErShxk3xJWYszoj9Sctow4MJWcwz5+UDwIyvasnKofwf/qZ2WTWHP7k
ODKsXYhDuq7/F6ue5d8xdq7RVW0IgYQlgru7PHsB3c407JItf0GlLvdmTodsbisY
UArKK+iO2FBH6us3qSyFVj3WR69Jb+42rzf1iX8szLb25Upjw1g/DtzXITQwrIp2
yEzLwO4j3egneEuaagaWj5rdi1UtmJ7thl5ud1TYj2tTw0F4HCb85ZbcjP+ZGeEl
OKHd7sc46jbt9d4wXM5e0Qsb2w9c1AcGp+aeF4kQI6Rrzb4iNaFl8QtaC7UTapci
WDlgLvGdpBp54Yr8eTC75za3gl/jKWo27ISE/OSKForQiLiduMxQxDVuvqoLFwpU
fww1OSJsgRjGqu9PZFDLp4rTP5Tk0TJUZt15ll5V3DAqVs76GjYWlyjGMpmLV4if
QIEmykOiC0gjn2GnahqvXEbOou0vCRD9mHQWYt9N4zQXSr+MuWYCKxU7DmZWDcYB
uILhPjjpjRlBFh4KebEfw5wTbpAD0JV7RDYEtMo+kitXFYtmzsPJadtPzfq/RXxe
P/1j50/vO5bExhZ6fN9rfTGRYyfQE02iTueyFtCJMabgRb7qTnDEuO93cza2VEBC
gZ8uJ1genraL6KY31OGiayu75XlxIuKEhrtLbxv/KwfFJKAVDyJBkBquWebw8HdS
0QTeZ8C1kT3xCaUJAQLXMdvG8jrtqXCA85jQ8GMw0BLj9WfHqrdMiDNNyGOASpOK
B+gJgwijYGivnnNFOBV6nJ/VVG67tbZawfRZM+Se5vRDYK0ZRMpduBucS2SwqYaV
ilgKgafOZdYGHDpYNCV1/woR5ODlnFTgUg9AI2xBRK7A2aMtydLVD4hvZSCArBSk
ZeTqn4EpnlYoECQvsMjOO7ThO8NYclw9voVXLKFZLG9V8LA3Le1hvuq4W+6NqFah
6IOxREZpMI8x8oJDld1FVYh2za8eM1GoWorvBdqOpWZsyozXH3JVEDW6Um1ObvQN
pzbvf0+7VkpYlsePAoKY+C0nSPSaSb6oi9PHgxo1K0zlBiULVV1BdW/IQjMVi2Lg
UYrQXkJcAAxgZAG9a6RZfPNrZDfEj2QeRGPmrqBvpAdlmSglQn7ptIE94XIIOPN5
GA/Y0z5r+I7Pgte/lafIdyP+nfxoUYkq64xXXR5di+o4ss3/EoBmsdXmY2rYSRlI
hW25atHK0PnyOUNGsLosyb8lZ822Q8R6TNS1SIU3HInE9blp+HMpP57Naip09P/U
N4wbtouDu4JMcExaQMiqsKTgvDKEFSHv7AaAeMnOoxRqgtMjmWYvjge+UWfEAwJK
Tu6pcwhmBZNjwNNy+P0to+7xlX26ByJWRIFkWnnS4xiJW0Skq0SQvwxuggdbtiMl
RtW0PHR/gLpHr9eFbqPNqc0aRfVipTPUQKfyk/nNqhEduej/LyBb0rsUNrYYHyqI
GQxsy+JL6ngZ3YK7pguVqEUrH3vX5D+oZt2KKm1tHB/hcxHQrq+21qsqs9vYtAqk
F5HGbK7AOrOa9o/8XmKN7bgdg+KgKP8dAeJLv69wqtQWjXTNR+g31aHC3WodYRZh
1xOPMqgF9A7hrgVpGNUrIF7xqHRclFCLlZVyJbl41EC0lXLm+RN2WmolTGLdUBZH
iUG14jxPuH1TEoCq+8j9risvlEPwcS4dFW9FDtZwAP5/j/tXHg1XeLMwYl7vwegi
rrnU1E4GgsIXltBfXmqG2YbMlauWiYVkaAIwg8T66W5HAPFraQGY3uDlYtlMVVD4
8yt01v8wlWX10IH8FsGWiYBAdYolH7+8T3UXHEouXibmN0rfFdJS3hrVTaPRqJG1
BB3vf08DhT9b6RwzMGY6cUxgwuUgQOjjdJ1Ft6D99cmU3i6+tirtnYd9kE9eNAN2
9vOA5HnbS5frAHBTWPij3ssWEnmxyx5CXCd+IvkxvDFwuM38Y5pJKtBg/314QGXM
kf8mQkARxl5THKfTzC4Yr2bxAtEEep/OrN8LO1ED+fQa2j9JibX1ldk9hQsKy9dY
ytfWRzT9KoCNqxBvSUMe0HWY4d+la/91bQ60sLi26nIArb6pn6ktPtLDffDX2NmZ
mpaXS0hDKxEbSRMbycitSjSaRQri9zio9am6sm+rDP+ZoZVArBFVl396+nNz7B+8
PIMh5iekBaHbQCz+1V8CH9y/Aq9sdKVv6MZ8jrZBZzp2K8UgonHoLqbhYQFHIu7e
+QAlyiR2CwtCwFzZPbr0pa93OhO/qdSKtKNvvRj1O2DO2wkQuj/PLDez6jcvuQ7V
WUz8WuYzO0gDYFfJ8FlukXFhH9S63qhgj1rgG6xILDGRzvEvu7f7kZ2Dr8V6Y2oy
SBdV8jonJcmikI/19fvaPUOvnc84L7mugtdHQInlgEY1ToaltEbJNyzEHGiwOFTz
u1BeGjQrUZA4Ksa2fN9djbq5QpBSK+6HcjVMwbrXju8N7p4AlBiAqUjrOqGxl+6j
asmdK1HUu4rA8tzGwX19iWifQ1f+1F2/ZUpdi2fh/hN/CbCLM9LbFxyUDQv6mBmz
vMS1OmubzjXoFXvRVyzmbU0xv+GO6Szd5I/MPJQal/6pUHzaO17GJco1x3tcLqGz
UTWzTEPwKfig2cGGrkOB/uJO9O7Vfq80JJTV8n0LXxLKZs7fH1aqPJQUhnV53x45
DyK8IMtkvIc6kkcZ3D8nDdAdbpaqI6pUiZ+7z42p2N6BTLqkcGLj3df/cwsni7eF
vutlrq2HC+f8/1j0HP7iDyZhytkJ7g2SwIVHGdkNKFb6zHFaMwJVUfBJrBW5A/CG
pnflRgVe99gBS9aDtQhG3xOFplq+MzKYpxFw63z+69jtiZyzRsFRNRsqWAruGkKt
UXjBVgDQTWDlyPmj4ff0xxnbXe7hfNetO5CazCuO310XQk+3WJOpzuafw+JE72+F
A93I9/UOa+nuhyLQ/sdX+mckWvg1EccPpsfGAqiRYHu3zK1dwqThVqrTjMv+CvAK
+eg/w6kO6QxbJ9opT0KDQ506qNL444mt3FQmIkPG/yj3Gf50QxDoZKnhgscnPR7Q
69pMH5YsUJGVxUd1QoLury+bucn7yxi4XjmnGtH4pdQlo3QD0ck/0ShUsAtupYBq
9k09C/DgCFwF4BeTDmh5fSQeih2tCsk2dDLVo+9ndZyxveKj7f2QkAnTWMiuNzDE
KvqWb7W5qgvZuES6NWbXgNP39TKTPB5R2oCyFvnMmhTd7mzqosOl5OJCoyi4bzOb
LwBnasYeQCADibQ9seCZDphVGIQWhUt0EgTcn4lwWVPx8BoZLHrpQpnA68Auafqb
P1bN/fM1ieHwA5ZB+wUTV/HFLVFSS8meBibRbSC4IWQkp5V/n60dI9q0G4VhTgtO
bTYwP+dPqvffStna6HCw3crkVY+AtFsJ+lZbqJGKXu/gO48PbsAYBp/E7WHiDK8F
mWcYGKyAP7O+whUm7EFgo2/x25cKvqa1sEk9wVcpjw4HbAaQMiIla94CTfjMTiOH
YblIV4/dtPtH5Y/2wo7nsC5nC76elfqBetLKEQvvdw5E+Ei03Mnj5Yk+ZKwArjqb
6uDdUCeHA+w/rrQoZptFORCrwiICT2mFayqNWyBJFhP9lpQXMyvoDbKCHhAlvDjV
cWMwjZlUG7SH196NBqhECbBj3by0vcr8Y+lyWfX7ddFOdh2rWW6C4rt5fV/ImmJH
bFi3aTIs+ndSqlTn5R2TsrN/jnP4EOUO7ulS/kiw1GTkIoKCY48wEWgfplQUxVo8
sTc+EHaCAShTeG8CHQZgb2PoiyXp7npx61MJXfbZuvmk9fjlHUY6b/kxyZMhW6nW
0R1qz8qHn4k9sLd92t3dgvE91V1n4DvAtATaUa0zSregIsRIcVQXmv1I4JPgSSpI
XVg3He3HAaeEalsbvUUQEf9F6/X9Inp4BXCxwxLggvNF4C55PEFfUkVk9aWz9lPx
GkM8zT9fMyvYvoubVmViMcU8LdDuQ5PvdOKpwuGY5oJVrUGusMVyxuXxFCE/30I2
fMEueiRUpHuEQPLY7f0XTRA5YXOT/nMBZ/Rxqxuhi3xXrBFZaMv/Xrldu4LPgxft
hndZvMlMLv+4q09rXnCxrJPKo5proeGWijnnm8W5C3pNu/iazlhvXcDS71p9e9Pc
azftblGhViX14C5CJys41NPTOeSEpi5JKsxZn+2vKKBWXWGci1oVchaUbW4ssCqt
4EbiMydOSbDiRzoZWJvUFmFwjivB9pPG6LyOgUkHslLnq4jFJB3GN1fTwqRMbVUd
RdXHQ9pJB/FZ0Dahi3YPAWOgQenyRklUtmOXx2ePK6vmWlN8/haAp3rPOX26vihq
oCGAUg4vq0jzrkUTdzyLrMQ39cwZ9iD5ZkmEIwtUF+3dEdXan62dklBvD/lIsuR2
kaCXrx1Qb7WVHWTKBDqrIKdai+qPZjAC+SbEz79RlGsPftcCSBTZnMa7OGAl721n
A4itStxKTzydr61Du4LkW7T8eRRq5CMLqMhZPLEvuaoVE/32ecrSyyjbmrhj5JqW
BjWbKSiZL/xC2v5Ya5OLEkqdmWmkiCWc+yI1frZe7gVbqC9uhyQYFjqEHWpwpp7m
wRoWtbz/yMh5mm2l01kIhaG4u40dATxOVPufxiT/uheRl7+cV27WJzxLR/JTy5e/
pQbAapBPaor7+o4wCS3ks7I+P66ROMNvgMeSSm89zNPrCv1CJmIyfDFNTPGO0Suv
yn7V6oALYRLPsg+HbsqOIMOMi7JBF8ggEX9d36A4YgPEXGZNmotM00NNM314tIQq
jkR2XNnx1nFNGQiFk004KIRqF/v0sV+RAO/FLWPubNMhZ5OaIt52fwe6beKX+F1G
PP+b9ipaxa8deAKMB9/K9/q85HrMqJsDuStiXzw8zMCstsUUt8WMwfa0P6xFUZt9
V4vYSHYHyUiuIy4y401pLHxDR5X/dg2YNjvXrF5WGyk2B8mXfI/OZ0oCRQGeoFGd
NBjrfiyfe3hhrtknByPgSlG6HOj7JvvE3fjStmIHOK84fuiQg5MWgZLajzH1n4br
h0C9T4oIOWyZscQdHgi1gdZ464s2v1eDga+3xO+GH5yAjjf4lfK8Kz50X/TaTJT3
BqQ3whY+3sc7ydVjSKWa3T7H042z2wnujB1x6lFIQTjlyGtpluInAmXivRDtmpA4
L2KTY6E123jDeaHk41OWkXvnymrejmnsbJ8w/XOR7ycq9U8SNbQ+4lbWTBadDhQR
novgZdKhCyjs4/s3KTIZct261wBrPTm4jsdjDT5ZFNUq+bo1rmH8cjd7uRo+Gcax
e8iSPKlni4/rFYxuBYl7sGwqikCxToKxIFYaMs9ZT2PKTYscxnZZMcuoDVkhy2uE
c5lEYIJ0y2yb8DtsVPc+PoT3Oo+SyM0oovkkezZMzzVPBsgO5nSJsfDBxifZa7sM
aYro8CzAPM3b3nNy/gI1vm20Z8Jt4FMD5h5oQXNOrgh6qWWV8HQFSFgyUIf0DrlD
i4Jj/vIV4r1641HJYn4xBVJ2FdfactYUh6Bvn1v2ea/mzFkPZ7V0yTWTYfO5A9Ui
m/lgjZXN+dIVKNsJUqdPvbsHmS59OUny/Vogqn1RyNMQ1J4rfp6InOVoh1EFpTuH
Y6GKTZw/4CrA0ricSgzWojE0MIx1M3ueS0hP7+gIGC0DF6s4tKxD6kImcZy/Ipkw
9/wFEmA6mXHi87lDeyRZWQ7cYXFcSPc0EZAH8xUaRvp8S69KEwbYp4Q4Wk3xka6b
3WOJjW3WjUvFb+ajtwl64ZyurSIXrsJCGfXKbfF3noyTy1vdErCyMn5+Ho00VZWm
WQJiGq8lVyISSf7vzgRzh87bEp6FniHOFIyYT5sEMdHChf00V9kuUcRGp3XcE66C
2a4rNWYkrBTCUSgfsMOPg4fmdqTJuDr4bAd2VqnOi6AucCQJlhvmRQrG9mcua9rY
nwG/L7wdw5iVYyLBgScA2qGX3IBZsiTloL322Xe7rHGviBJe+hAkcszKErY3/OGg
qSab5BT2wVHqFppJfTLEX8Vv2e5D9RE9CgD/c87AGHzxwquhsISa5k55QH2KehzD
O4sTZwhSwOajzLIgYPHDAeWrp7FTFeRu42fujZ2Cv9LVeKCd4xdrqYc3X1CEQf14
FuRSgDRe12krlbIdifsHz8hASQCzGWPa4BTk3ZkEyRjZ42b1RrN/lMOS6GzGtjUE
H7j9QY3j0e9NBqBupyjVfmkm9ZFO224Eo6AofQLFjfzOFTOYmNqDzvVO4cB0LupZ
zrSIr9kSoo70hsN/hq5UpIwwNSgG9BplsphVfKHY/ZzSGKcQtrsFgO23o7OJesD8
Oo0Db2TXfmQXoXUZa8BNICZEKpTojyIw1kl2AESqD4IuJYwzxcM17gNK2PaUSf0f
PZ/RhSkCdg/EQG5+lQHSj5sJIRIVmcT3/k+Ncn/gIkzOAKRDpu6a9zBiMQiif3C+
Ydx9YP4MliD+9onQjte2pys+9rTDo1vRtqVfTjwQF3ZW3xSRHIroWVdGZUBTEGAK
8t9StMmHnJx5WmCp3OTWbG/V8j4d6F0ClhfaDw1bc2qvNuEAWKtUsRvGsvMaNQK7
DtlI+BuPiKF2OFYLgh3cnp5E6ihvMTFE4m4aIXocEpi3F8jC8H1on86oeYdZLcbP
yw8AxmOaH/neKy22/bBKGw+FMCfP9VvyouaaR9I6CRX9Epsrn4LbP7/uFoNrCFTr
qqUv3AmOVJSGFEhaLD73nNQ0S9+yq56+zyd4z3+sxpLjSmMtRbDmJhJ3uSPrhMCR
P/4ounIUmKj4iQGMDKfrdHiF3ZLxu4Cp3zWYTpraddy22TJND5lhqBOl9rRm2LWt
Wk0aKkrzYgKO612XnwLQrIM1CWqIV9HN4iCqafhyiGuJx1BDJiX+yanqAlEe3KCp
JT6+RKZjcL67E/5VRp89wMxhcFCWQ5IJlOlOB3MhG2Rrd3c6gFCT0Fict9W7itya
9OLiaxwkeUo/aEas8vg9spS7GY6JbMXt+vXemya3TbDi2nRLxqZNPRV28wMnBEyV
m/xnfD3gxA43HHXpJA5fqSB/5RdOXbh6yuq1tO73V/LcO5ucv3DoHVRLb+eWOAGj
fqqm1dRkdPI/9AMEUllTtCsrxOGE9NCA7iFGzqCOwAtCNUDX/XOGtYog2XyWN9cC
SG11brA3QY6wjKko/6VqAU4rcKaFdPXjpDth0uDSno0PN8Ba2IoRHGi2mEBMjnPn
uXbY++wC9CgkzpsgvAceayi2o2TArVBlJFGYy7BI/bNHtryiLqCmzuwhTtcH1tDt
fa2SyutabONWZ0Td3QAfVWKn5/ISauuqR2kH4HJAaYvWnfq+2JtNGW/6ICpjobln
wdFdrUt6W3iepAosK+BaXhRw+5huE3SEcRPgmGgUQrONh3LjwYGZWzJmtq1TystM
d82sIwUCoDMuFL/WTBRVemTY/E68jwol7/5Ubequ+N8At592RXz4cU0HWRIvAdvL
1lUZRqfO6VCB69A3RjV8hjW6eE9dW395yjV4ZLksPXSsiIv1LoD1mOAXKSyMUUTD
d6GaT3aa+G+e9XK0K/G51YM+NBRtbPXIepWoxwO8L2eWgqIKQUjEDWvbnvnY2IX6
2hnU4SXtB4dz5payCn2FHHaZyflSMmG8NB1AXD8y+cpnmAe4IKotyV73wpYcPLTJ
gF7YN00NlD1ApDhr0sN+HGqcUP8PFTRXhhO3t+Y0PFsM0PpfPK/obss/GYyCi1yS
LjYg9JqrvCZKVgwUc31D2rbAkjq7Ra7etdNbMNMALTPGFR8pt2t0FL3knbVc7uMu
KsoPW0NVdSHDcsMo4SamsW3zFpDMPAG+S6W2lxNwcYlesFWEqM8nEEx3WHbB6k5c
cr7X5AMK0MPwjsaRCUrxPBIs6tbVGLm82bziH95RB2wVZQOPHCAVjZaWBKbVqe7d
1ssQokBo4SnihzYgfAxxAa+uiFYoglUCj3fgQ9LwMwm/Hk77+zGA7xl6shpzoVu7
ac/jCdgFmradBBv4QUeJl2dyBU98homlbLLlR2hnYpofCPdVztRCINzGW2TfFVhT
c1IZgQBAAlJL0gnWrHxkHePT3K1IvbtOZyjLB8InOXTO0MKYmBNMBoMBBHK9QWTy
RUO9W5FsDPph9Z64Dmknm7GPQxJ/gE3voeWOwyUNzAJ1AKDzaUD8Hpe3e9/UANeB
HB2WUvcwlkUGIK/2Sac60WUXvHSFtkN9eWCFsyM+TAycQSbuzQ6cN96djyusfOr4
1w3LSYkzT4xvjSxgBzWGUSnAHXzluPQN/ikSmcBDRF8ZSdgECwbI0YjAmfREekwH
99LC8dhdZ4aMVu9qrVd22Um6r1V1ICpL8urupXD71Z7u9Shc+VVajPitHqfmBSeO
smp1fuuBH0kI+HAQ49OD8KXc77uETWPWZ+mKCSKjxkTYRNysBhuIgzEObb+UUjWr
Y86v2StYXHa84GpgtYewTNBfzfbm3y4K0kiphBgc5MpzkXteI3EPcJcK7m880rV1
l8iiKPcISzSxA6G2dcfGqf88xd41N0zP4aFBHEiIzt8J5KRD3r8b+sWDJrljntXr
0rK5fAoO8sHgdQfAWlMAk88NrduNH9qSkLg/90cJCUwOtuzJ0rvgK2mEqdHV0br2
+1PgEVApKbFMHNpd6wz0PHo/3hV7Qu1JhENXBhIN/C+LZAX9fCQwENpf6qFPvqtR
kv+lCZkP/4934iimMxa1Q8pQ/Z+9Kev71wp4HL1Ae7b8V4sHimG3MYIRH6DGR1UW
mOh+g1N/gp27f+2QxKDhOkBjR2oJLez33misdxb4om8lEBBEULOPrB6qyedXXLMR
wpuNKhz5YZKCfLG5VAJfUuTjyOWTn/AMYg2EQyoAklCMXW5Tek3XU7KZx/booabY
nQADTZ540z45htOQ7k/OtEMcq1Iz7lJVvLZtQPb/bNk7CPi2PdzOeXxN0MZeA/d0
829tGuCBjmYmegxj08LW9ViHGomTA1G2sybTI2dVmqLqnFSBySwW9K2H7hA8QLYQ
OjeHsK+ZVEKesUTt1VXixpTqM/lsTcmj7HflSHIY0eaUHJkzgGOMLKmoq1JaRZws
TgKchfSxgetxK9zNEL/KrQlzJzapTfZHVKcUfMJmbSla4qDRYw44w3hLRIukw6zM
viH1h/gB8fx2idbgmd2OnGi0/iarqUmwftSY4saOmn0w78Egnr99QhuVY9PuYByV
dYeDCKRQXCjaN8rJFeQMAredAzh6e0gav+BApV2bhIU1OChcNtqrjN1sjycGfFzo
MLamHW985EOd9Mb/13Sht/cJbENXKJXMirV0w3TBsXRqDy+5jYTmA5Q+eaFmlO8b
nq0j0P+iNEQXpvIjcWp17iEsnzJbjM+dkorfszFIKMshThJYUW9Y7oDMEVci4Rk8
nkAf9dO11aCUZalMyLrv6Bbo5qM7g+lDNPmy3P7y54qI3aC3s9lxhvoI6AgY4EDu
1DtnS10beV946fEyA/hPgdYHBWAuqHyZAgApU8yXwUqADmdDHywrB5avsne87mFd
M6EuxKEBCg+H99rm3fA6nLV1cKYUVcwjVnHkGiirbTT4B3/bFqqgbSSqmXPN/jPb
YAPlUXwBB4F+oWhUoRU3t7rXUMEVkJYdFBsJEjSIXDL8yykbujIJbKOUV71xiIE8
+9Tx0uMgQtB6Dv2xZd2KitvOMrslERM9TOsnSaqNkatqs8wc6WJVed6u09XE6ab1
ZucNWhIvyUtrzSW0WCdgySeoBLhsdf46l5NyX6lFLvQgG7lZMMghDYiVBNMS8QjS
GSwYIVS9uFOA20omj6BJpUL7nGmis7t0q9cgDsPJyxx6azuW9LLujyWsy2HjSbRC
u+GrPDFQhMov0s6FypKZZVTSgddujw8GHipFCpx7eWUANRnGOB/T155HH7kC4J01
WxsBVcYarqg57yAUUYtDASrjF8D790wU1amAFEIrhTWdNXQ84IlOo0PP6SF9RLqd
KFWaC1D39q5PTUQX2stZ8kTOoeWf3WiYovUC4iYB/+b48G43yhRuCUBpNaW7NTQN
nGbd7fz7Lo+io4kFrXB7ZfUVNBUw4UU+3X42+JlH4b+ReVF3IB8pOJL/mSHLpFhk
eGHHbkqU2V8UJSvBx1tH8YDGJBy+a/2yKaaqTnhi68eAVfw8O90oj6BL49o23Rzb
GlPu3Ynf62emjJ+y15Jf4WW+sEs6VcGYfv6m2bcJEVZ6xM0kZ2hkofUgYuSonriZ
dBqKyhQuRH2p/RQo+haG/aa47OlyBlAgiVEAgnuuT/46QZXy/PPlitt287BpEe0p
jMDG9KfMHJOPYo1TOtbg9OHn1Cm64m8+EUkRK6PwT4KK2IdlYTrVpvmmb097lr5a
eqOWmfcgzSWpnqorW2tI51oJhhLbD5jf9vGMURyHIeg2u/NZEQ5xkAfO3RkxxTWx
eessHvJvt4pXCJx/4Fks49xPYwI9lUEI7Ste21qhLFzI6gX2k5JH4vvmhdGIv3Yo
DyesgwijlmKw1ZxSWBYDmhXdQA/+qW1TMlZB3wSFdz/szmbNVGd2WEwjLkpRvblM
qmmyKTpPKe6jPYTONlV0n8RXFIFRTt2LdeIciGwIuYopmxnFRQCRK4WWYG696diX
EBpBvLOaUftPtuiv6lBizZzKXiPrAOGggnRimqICMSaSHSdU1BEvJ93XAtgXTYHO
B/RQbiCVupgkPJKxldnOVhLIz0m7PjA9wICWUmPRDM/BNoJZntOmq2ieT5NL8ebj
QM44X5W12bwgoI+mFJmXErJrCGwXHOLHA+Cv0iwgX2PnJKj9wIraYL1ne9MRxXkh
kCJ75c2c+Wzm696Zpt+LPxDY3cCRg/I7rcEcDpajBEk99Hcyh9h5QXEwnCHf4HK8
Ko32crRwyrz2XA88uSbX2HkVDd0kFDJD3YhqSwOoE2VCBryN57x2/8QczDBXRxdf
AW/BBAapj29NbF6+10FrfK61e6l5+opWOU/uvyUaM+f98RTDz3tk6AzpZVqBkL2i
p1XLcORi832Nha19anJv3Xu2S6fRN+EeJmvUExeART4ggsz238kyMhY5m6s6B5ON
X5nC4E44fDDarIRUIZVzaOjwzGmGrExPU3olMtI3w2VpzE2cnmwyzBQK7mTaSEwr
gTiIet9Hh+SAIbLStOmYWHta82KjIhEk4W6g3ubuT3c17CNl1vUBHUcyLszkxFtV
G8zkHqu1JYNpNmGSsPld6AtrCq1SANw647F+LIVM2lfmebcweawJjrqr8mTugzTR
Rds/p1UqN0YQ3R1JPJu9p6zofX5ADJKQmmIRA4/HiyojAQ3hclQXIkBJP7v0woAT
UC4j6M/0Hn6qlacaVn4bKT2XTSh3REMqT76HNVidcbBkQl4cS1sKo3V6OkxrS2ds
Lmxhn4ZPc0V9tJBfKV92uGDR8jKnYzWdjtF6DWnjb4w7feWJZ3xlZJyd3cFpJaky
UY7X7siW2MRI41LBWaQr5O1QNkYreIVobSVCZ80BF+gKweUNLcAaWmmNmKYVkuNs
qc3PzMccdevVKrF83VGySEdvzghbdvAaQIUZGm/9+NRmCFRnzlTjFkmfdk080Dja
eLTZqqnLmPF/wHL/B8NNxbC7gcVYZdXQ/EYM+i8G/YPVCvevgjUuuTHcLB0w5LYl
YyTEQ51clvqhExv7Y701bDikOrRZFcv4K5CP5vHomlzSlKsHvRLkzA5zbYkxF7Ba
dIK72nCoJxQSbWMh+N3J7fIBUSaUZ3ZgocXZ1dCNiBrdja4EAitwezY65tJonU+8
ho1rngEFf9Dkndx6Wl2mrwJfKBZr2mxD8boOM9FGxvfPDzT2jWtvMoHE6PYby1bT
b8zpC+G37+aW7/o/VYImounKYGn1oVb0JjGgfrf/7vFXwZpiuW8Czno7u7+IYb8b
s+X7fpn3JFMFZMCqiqCZL5C7zCvBjj44gmbrixkf1ooooV4IP9pMgt4Z3i1ZM1P1
BqYGLiL327iMW27+M4MtCOTIzlZPOijq49ZIFo8Es8RxonQBWjxJIp+f6HLym+7j
jZJKkl2naodZJsl7/amu1S8ECG4STdETcjeGiX8n4NC8eAy6Ju08ts4ROXMAF4+R
wImB6wQqqHpSIfHeRmlg4Tb5cl6BWUTNRAF9YrryBhk2qdhyvEju8gk65ont/C+b
sbsAbZ2Dx76/pmtgrx4NajceBnmbWCzR8Eij1ZV4gZotqwRlMyYuAnYio4e+0voJ
9PATimNXC+WmWSkyVKQkBaoNQezR8Klzj0sDdpWktOT1qFYd0p85w0tEQbHdJTgN
iY+qSupNBkmKAJH5UrlyDkyi0Vp79u6nwU7+fxCNcfsUX1IzDGz3vnwzWT7KAy06
F94L4GhgAXWPSp+ObjehiLGhuPNL4Iz5d7E3GluFJnrMtQHPw6ovSVqBi2ptF+pg
hs1yL2sUHjqFpzkPduNxnAVsJPkcntf/PfT0c3ulNRQmCx+HW0ymHj/VWXgQKR46
f0/vD6c+AskC3i4UYK6OW04XwkLna1SH6SOiX5YOz6lwqIGC1kCxJTxQJWoBNS8N
tfki3ynaDIj4ox4nOHZLRQ7p6QfWahZVNJLQSQ7b2Wzrpykj/XWLUKtD6VDh0wZQ
nQC0JosmCCDy7uh0BZOZLZA+hM+qEqicfELXVkfvHLQ9BuWxfyuL0A4/zOnKoUHq
LoJkXUVZ/NYXuUFVJPr3Av9f0oWVh+Xg71cAHn13fR5zlg3KPCR9K+KipgfKYE8p
kdhzjxEMjcpz9mDMDF81sjgI9y7XmWktQECb06XgibYST8oz/JhRF7hl7Nbsuzi1
qPM5qNdBGoWc3h4qMY4epJbPehf0M6biq+ySok+g5q1O4WxqpNwZ1P7km2LrzUGz
H9rSrZPEZ0qsdMFlPr/TFOLh84B7kqZMcvnEYiPuH0v/f9G3lJOeZoYyNgxkePF0
uq8SVwgtcwBrYKbMg31cjj7zM/MRBCX4HJaQNH+f9E0EaoLygf0BsUmVE/vCbxjK
HiV1JpZ2/ee33M3B1N5JnWTo20NkD8Ofhr/wnd9BZ8M9vturQRzcKffdn/PbtaPZ
gQapy7Zv6TzcAErT10rsTsHx/iCi1oTrI5huBNtow+Pi05NQHL9byrt5FXH/Fvk1
Lv5tNPOoDarUqsVBmbdgspv2/VVW0AtavP6uxG4nZZRh9l8mE0mivjvT0tjoOzXI
bbuc5GnxjKaNI2jUZNC8veq+VS7P6pmvdNGwfqaIVIv2odJv4Fs+43QdZudjq4KY
QcUmsoidaDFRkB0iR1Yke/06LhAs69zhX4kx4uFcNQcs4SHuxE07cqy/Gx6IsSWo
qJR4is59Kuv9cNTIgwJr0Rh3VKeTk7+i3WWqdBognVb3TzR4z9x6HIpYAdKfxZl4
ErnzVSZH1HSKaHikehrqTVbPtz1u3uO1thMV4blS7m4umwZ5gzEK2dypzh84G75F
locWJZga1v0FxOHwABiyX/1J0hhUTVcgLcEkr4U8TIJu8vbzmj4LJzcoqV7jI2Xh
7g63LLVXRpysbFWO5ZUCsu3UsADEbHAu48XARtpWja6T6zl4lqpa5N80U2keFZPN
2ugK5rxDE+r/YK049h1XIcMF4wk7JN8fwBUxoC7ErZs5WyP47uHsc/BkxjrQwwa7
T673abPIv9Pa3FDQ5tmOVUwmVqeHMOx6pSXdqp/Sns0xsH9t68Cv/Xo6HS7xDN0j
flqPo614NrBMB/p0R4wgNEQ3bRnoW6WVpQCYzZ6IIP0YnYYeTs4NuUpzlqyewTvM
ocY6Ke/NxUt46NB4KqcG8mo2ucnF6ZQzrt5WKjANtgohK0WW/rYQipKS0kpT9D8Y
udq+XkrmC9+WuCM4wYQacvy+XoQbNO542FdXd32ooQlaHmNLpXZRVqFKPE6uBBlW
20QrKNu7YgmvizJULr867FO4A20IHkRnWFhZNbydK/c558FpARmSGcRbcB+VlKp3
QXnImUfsAAjIRZ1Iy7L8QksP6HL26RD9k7fUIyYiSNAXQil6kimf97l3NEx6cC7G
yMXI2bobM+1eJCxcTAFu5egZ4c6wfVmpYRxRJGwvsrBbkI/Dswn5V3K9w3rdB1VN
Ke7yHcxrhf8i/5r+Id1NLxro1mMCDskiXzzkn9fvKE9eiVE9EH9kIksF3nqOMJX/
nApVpbb5yD7qFLhV8BmBLI1JMqeSdZ0ukhPhLSjxpAu5gB9GdDCOeKeTZxLuoPBS
PDDPYsQp9iTi9maIrNChvlb4tLPq3nkKkE7sqOLHIdiZgYwIGC7WU7fjoDAR9e+0
vEn2uiDNIjtzn7RGfplijoLtok/NzcIzWZ/HMv+HdEVuClZ1y/jlSe3C6z3SyXly
1kNPUfK7MEHnPfxho/R5GGEp3AAYM2wJeff2Ysbo2VcXm3NFy5umJxBzi2urf92s
4OtGHesuF2cotPR1tD9s0g0xsK4fLshAyPspJDKS3ECrpvSrmlv3Zjbhin+BYM4a
koZBAEHi4Vmyh166Ps2c+CETic9mCq4DogcAbeW1sn5Bze8Y2behQ2Sye6xnjBon
vVGyXM5+WJf1hon66WanbjYWXpcHl8ZC9Czc9f+1pA/KOVl3bEurAzGOcNbZd3Gd
2qu0Kzf1Azp3qOtdV5OxdoLU9Dud+eWWadMvvjRhJq9hG2VBHH/hKhfOYI2vRi9w
zpkvOb/8nfrpj1ZNA7X41xSniyN8y2dpw35evnIeoKMGLFZPUYZvhdRTLZ5haTou
o8qYrIZqfbPflVcDkJwBy0mYE53MnATxsVWFxazKeittTEKmfxOFIfTrVIDFzJrw
eIYXZG+jw7g20fpDJhfy4nm4OB2fHwjI1HPaFNI1AAyfp5ukUGzo6tesEiCM+FMu
3y74N5ZH0tz5Z1Av90fOEfBzLwUGlAwtV3wN4gXXPF6EI6S5TPv3V3Me6FSGbyjA
F7rhhdUANeHTQ/g6Xs+M1k3Avbd2v46OPEXyG9Op47de+hRQlm6rcLuZQmhqxYDL
BbL367xX3TzEMjCO/OabaLHUmkL3Wp1NiW26oK2+3DSY7ZiVkCxbrcH/19ioEQ18
MYy6yIMtoRafSikmy7FbHrgD0nd+5rm4FnfVS6bGk0gWrXlWE+ZN2FjnZ3TyKZYI
sGWBJKPVAWJPdfhzBANFXxn/IKpGqo1o1bVWSqJ/jiECnh5mVzIcAKTqz+u8oxxG
7+ZLEt5Mc5yuZoxnkeKlvARWpbFIrcdP02VFdYprIpziKN2i0R6ZCFHdqDmwOS40
nLVgTAFMhbX8AGMRjmU7lOVNQ3uFSdTnDt6ejQILqPEWNdtnR1GZy4O5OirFADvi
GJA8hscyKYLLVUB2PgSdZgN8zzGo58U6tKOczB74FQJBkJRBmANu8aYKpdvcOIxV
hjvVxZulFPxYYnFVnU5xvn+qrd//FA/MNEOtvay+nxmLfHOp6F4ibiOMHUXhSIq7
zA+nClLYUmQzh8t3ttH6ZvKVUG3RYKTXk7k4IXW3IOlvc2LkDbR9PCOsVVDsbYs9
lpK3jOZvbJFtA168mQDZtkMfFEftwLevHWgNAEDIJRDu7YFjgTGbiMeVP3ZTBHoQ
jpx+KeviTVPfMkm9Z3Y05RMyICPSgDE6eVFtqMVIh+UqzOGKOP1TVbnuZXckH7zA
tYC/Q6wl5MUNpmlA6RHkKt/13PT85N1U3dCE35GtdcU50gKbcuOruPl5DHPERFdU
KdlfEn88A8LG/WrPQ1uQxh6+tSi2h8cPEXu/i/PQxArlnfAUd1OEmIjcrad2lAwP
BoK2X/lZv/dpQ4PrdePCiPU1P9V9PjgZ9X8YMlfI/CSMPMiZ+rjM2TljEDox56FE
hSWSQM+xmy7cqCDcQyKfK9nMvwqwCx+HPJ/GRzQQUc9S2UEZt5vGrveSSIQl2bQs
PbJ9hh52TjPFXIWt1gCHDFTmHjU11SVMO3H0Lc83eqK3tQvVbuC9mELq88GiFzSH
Clj2BZJ4h0bGKAMSRXbqm41sxJ6USWRYdIOzRk6dYJ0v7ULHsOcEQ8r87UoIDH36
fezmunoEawFzcPu0VHnlEcDWXae/Yd1vV2kkuavA/PCRR7nw8WuY7Lzhwmz14UgX
mXsYEznSHZyAjf63YhKvA3KUUJHY8SE2TPYEjDCqs5IQ0rx9GhPTA1SdmEW/fxN5
RVYqrXa0bJOylF+kkl3AujM4DA6xLZoQ1ehIBrPNsjisjIyAW/xXmLG0SpiAyo7b
5hx10+uauhYnWCOGv8UkPW2/2l7EPNur72x56luF/xmu12e9XwCT/xTcpL6uPplX
i2vli9Oa9haYTWBlqDtKLJSbfGKZtND89O3dFonYTJjgVLwVouoPKTxJcJBdvWNk
DHrUs1RS0d6ag5sxCgxDPPNhK+fUrR/Tr5XaLtsIsLAx0MYB4UjLzYASIYODt+P1
Toz8B1kt7R3WeU9i4Xo801qjxinliBu+TUG6JNVunwFjBYJ6WdvJN7qN8sA3W2JP
9hkPvcKlpVqVoFNJmF0YiF5lYV9fou5sDBbKEmLFjlMvKD0R40m1U5/8DByrisue
Z0sHxvb3XcwdVMYQZKc2h4Dyru3CPTA1YeZYpRlhbzvSdkxBtVnpuJNuNku9An2t
F0xKgeSUcc/jJ90EpnTkjnbHHIg3QhXbYp9OVqLNBN/sO/JPOV6INf3aIVCL6A/V
gKqJz29HC+LwdPD38JouvqTEaaesUkazAVZCRGyMgR6dar3076XIw74ENayGYYYj
vQyiBcx6I6LCANBw+r4KJd1D47UEduqxrL5MImWxwjeRio3wDOz1yFqQPwknpeOm
2ylu/+fQak30QYMLHwTHLo+yLI8coAPjxdZtIlZXCMNumMUFNQx2NQYJr1thBbSO
nA9IaidWvhsV+IYWWDuoyFMGAGJzJ14jcQMeemJTBij4ZqoNTvHMIeI9wiL37Yf6
Tl0bq8Cgk+R3XQgx6bGzLcjo23BAJCFcggZeNAXt3hf6UWTqlvdQgKpH8ATB7ozX
c9PtWG2mHP48lfE79u/tVykpzSwEjG4nlYZQL8M1B1dmnhFWsOhIfrnJ0IkTUx+6
eqIBax/ZR4Iiut1syFG46cYabxBw1Nbc9iFgAzxobs2DiDT6A/3s7U5DASUkKoTt
FO/jmpPxJLUGOu6kCxJByPonwMve+kRmwXpeET3go/ZszXsJzmElwq/8lO2b7UCN
btN0k/eSk8scUrGvHv9SAQHpcpeljFrBAdTClr4FsejbvpqgikbmAiQ5V9Z02UFf
6Us/MnGHcR/9kyuWroPgm6QE+OUMQ4AAhuya3mM/LzZq8RVWaWFsyJ/bAeQs+Cbb
kWzKjWITgSIUovGZU/r8fsDA5vWImp3AKjtobg7Ev9wxViAT6KGnOMtM14VZscza
OChtqfEJp9k7hDNmraxjtNLx3SEvgrR1tAOHwRTKhpfpvOh0+GjEWONSMCJOW2ao
CaWwfocUKC1y8RrymXI87VqHoa0bOJMGvx9dQXP0etmtV9nwjXkFYgDQAnSNMI5U
4znyWPbOj1y5ablbxMpStxopy8K78nu8Wt0w7ik8Z9R04dnQu1FVPKnNi3Kkrvd+
3u/w3bFNeFUkRYplvcY9W/MAth03KnK8fLBtN6mPFU/ErLErnbhz4jjSarFWtMnl
1UZBcxZ0ehMHBamoYi9icq3S6m3Fz6I31ki1VXI3gyJlwWsXdK8rUX9M6gUnZQdv
U8a1Y0vI4Z0AHKVgKoF69qFkLgijh2NabzYB8ppuVBwNfNysJiDUGBip0O08yVVn
iw72XDvrbyQv+0Si0qoo96PDJFryEoIYhLecl6wqnEz3ldRd0j78SoK2KV4+m+JL
gopWsQqSpBUSKnXDQn9C4oiME09F7RBTDmzSRriO9xvNJ2VLLcRE3yVut7H37MBs
WYr7JWNRXKxBu08hrvFIx6Bm83usjhCWk4G/iPIh9gxwigYGjMCGZhAQ5l+r2pE3
Q8WdIIWtCjF0QU/g2Gy8PqatwHp16dxfldIZfGmE9Kbk4ZMVXl01DXdWtXwb4Q7I
uPVlCH0PyDRepw/l2qVfFD8ZuslFGpp0rq3Q/bA+9C91si5TeFcIQPOarhGtz8C7
rgIVX9HT4IAWIh2rpw8OaI0/uGQedk7FSYbL+qVKFmK1pbPyPbbjBl1LvqOiD9qK
MVHS7upeq1r4ofU0MKOHJy1Ih4gPqHuFjxsnWtg0tCn8Ga14oepzZbzVe23Tja6b
/iMrWuYuP9yN5TT+ABOUR8ichAqkagvbjhXKCoFD1g4NtPUk5/0v5UPCCXeLvm5S
+oUquvHUR0t1I/Lw8VCEjgDNKApwale/k12vFwVMNCUWqVfVIDzsqbEwRZrh+Q5k
wOWx42sKndJrc9tfZpJK8anA9SNZ5FrDDqxDunzfRP2yWvZxm4i9lH0VZhT0ce8k
+kNNcRjdgdk76C68iEsSLPz/fUN1gBwbw6hyp7fIOqKbUj+RzgFf5N8dUeNPyODA
EQ0J+vmjEm/07S878L+iMDvO7gaKhpfj96ejiU4vAR+5HonzB7NLVKt4WhgHB1Ia
mlIBsNcK+Fcv11s+6Jyqk43kZ+wd5FI9tUJIcY0MxY5JfELnx+K5NNt8WuHqA0Pa
eoMCpy3Bc9X1Ysa85yQhx4eL7MSgJu+sB0tLzbHDS3RyjB0KgklqgJrazDwrXwpY
pR4q1VN3o0Y4eO1SNwVCfHCYukMDzHZ4mt3gJ5CNQbNZMsCw1StN+DAGGTBtIhjf
nYn3JMvuB5qH2x7smQY8jJ3et9F43PG2YLx3j0DLQmXIWufpnGdcwFPN6JqaTR/e
M14Q1k3PfNevQQoMLlL5td51BM48iBI+6E8UEEH+ozhIkHNGXZQizJpUipTM1pr3
XPpwWEzTNQ8aGsUYWQr9wS6xvyPwZRuMh2r827r17mCIyjH01qtqIoXUh+D9kU7R
ABz6UKLa2dr0lWu+nT4AHcd5PM56KpAfNGNveA7gyTEKzPd7jmzJ+9w/Wwc9mL4A
FSSkC7WsUaheOg5N+7BJtxClDQCXT5oNQ/+XYny4hB9y/S610eYcajKYIGTNP3Pn
IO+RgudiqA5nQkcxB0fuho9WswTTcmQsrLztu+SZcHSs3c0N8ArcDkjDN+99EwvE
T1FYMBu9LFQHsIholBsVB3K98tHWcQ1xDCBmQhl6vl+nqxCeIA2fh83WaombHlsa
5EGvFromdZjottVewiq8/Ej11S/oLS76lACsFvJ5GYgkWNX+98QcFEg14cCB/jBI
vF4DBLVoN2gL1SwfwRvK7hyDK01gx9CUAmv9S3ChCz5ryDyrEve6yy8DYyRVcagk
hpRzptcpj+EPP6kDlc7/9CoQw6AKiU9Vp5Wmjy9xVqhFtpGY8F4IJUwPlYjcf1TI
8WYJyG7QS+bTyaU5lyhkxJAf+vBnCPCKbbL/PEciyBRtI3e/keagTbL9D086Vr1H
5deL8U0vBfCLtic9S7d6PFrIPl8QcsPz22QUovHQU6zA7SbTqmKUQXpFuhmixKFq
9iekkLGXLkwfjoipAtcqqCUpuovWNOrbtOLlBKhlwsJlVy4BavjMQ1AYcQPrr2Ru
Hb1rMhYD8c21ztUkEnimwEM0S4lWBh9KSnWKFGguFVQk6OG0IANF2ZSTusOxoFVT
3pQ37kgGxuIjgoxtrSWTv9e49pMJJ4UO92NYsTDoiet/OXST/tZueLpoAjC2pTKL
grRjRWCO/W+6aa7UPtebVVbqMv3C+BVPx101GXlNudCSSozwXwjMppWjRsVuGnZr
/mRrlaeX4DD7zDc2+KS/hTv0Dzy4QDCLkjKyWGGa+YAeGTtl+rlI4kGqDlQayeL4
7pFoCTl7c9JRRk7rWEvnfm/IHEK2LJktTUxskEffOFjZ1AJw3CSoamKV+jNZDo1i
YKjJAUpH7irQRe9fyEkQR+1S4jVVQVn9jIjQ47J7MWXkf02068m6OiZ6xggr022/
7835qpGsRKqTm8sG/4w4WXzmxtBpst87wSAc1zN+EVIFeUaUnNYG7I5OizTFkp9P
x16OILd0SN+KtyI9/6vJW+ZIOmwCVcTgDxBz5Qy7OpEmvzp+2BxKkO+dQ6pQ8MxF
XYvoKr/m2tDsG7Lt3SrFVVjrvT2SUFtUpZ0pkM6Qsx1P1Ug7aiujvgmEsgMKoxBn
7ztFUQ73Q+JfG8lrtZKiLAsZEVrq1h4HQLwsCF7DeYgGj6Lq3JnkWuRSAvMkWCZX
Jn6e/oIBzZEbTbVXQWcirp4+ZN1o7T4Zi133hiZJJ6BOomg8x00KgMpyMMkdVZhB
Zs6reZQfR8t2uOsaV5SSg3XDDXuv/CoMQYXjR9CWNFMsV27+vu084mqph6lTIaH7
/br8nk0BEoqDLCVqbPIIB3u7vQVUJL6Qr3nxzyWt7E8c2afXcWUkNjfg+Bx0LB90
2V66eFXXGFu67YzhlnjoebUv2uMCfAa5hxmrpFtOtuyXdZszlZsIwae8hlSnRwny
80bipPJY1p3pKzVVDVOESyQ9ideHnSBDpFO4fmgGNOuSed6O8tb79KRcvxNkIzrS
gpgie5CmT3bERhlzTBPP8ps+FXaPWy7fjXsYTS7kxdR5UvJCJdpI31iX1bESBS+k
8I3cf92UHhzGBB7A0GasXuAJkrG1wv6AH+bs0iLZWheL7Vn9VL7jH46t/je1INX9
uVeOFd9rNA+i239/tc8XjXg8tCEfM7syvPxfuCBizOCIwSPQ834gM9kqF5ic24L2
H19nWKrfcE/iLIEsi0kxPfalxfRxuNO/DHuLck52R31k67oucswrjNa8eG5h4rbi
Bl3df6oFwIBjsHnBeKG6kcPyQ1vN7y8OXwWZl6xShBqIbqUb5ExPSX+nENBwt7aK
64OHyFEWiAmT8zsmukY4cawc9rd0GZ6aEim4rKnqndH2DUqHQ3dUsQoX1o20/mSb
B6h9qUZmA+MLpSUpzhghZyg4Isd81SZrLX8YvBFP52GLmCein2yU4K4SBZj8NkuR
ho5Y6VIor6xpFtT30/LXj/5wt2p+RhSK/ZghJt1CVziehsxDLy47zGJM2Mf3aXfp
TSZrUjfwPigJZGhPFvkmvVOpDVLhmCtxZjyy40EE4s7ONFlF28uZ3zM/AQiL0SqM
M2RcKrRcx9SerGtcAwfyXYRNruGkErh2E/2HpwJEE8kSYRWdmu5xRZK+iCaOKhSS
MOHqx/WQrBzqmfvbc12+Opur8t108PvROo+gBkAp7rZCsWioh66QNkj+/jxCjFte
uZhAyvrh6t4mjzBYPV5VQSx51JgjVuDOTha5xyrO5m2YVqpzMVn8luvxMWF88yZ1
8MgF+qbWAhRrmR+Qdg1KyoCQCT99IGBbV4d/9H755PbglHU1qWsv+sGKZqQd7HvP
pwB62xzwMixMC0iJQbVovAE6DnQJisDKMrM5g6+6Jz3ROrDlCnyH5HYoNsM8WCKa
tnwVltPrG4/xuWq1pEkb3QOaszPHLcPvTklFwjLxV/gMvjirXob2uCdJzOp1MNTP
3oG4pZYj52i5KzSAeGGFAR/Ipnzvzdd4BVfGWdFcbqJY03G+DptV+Vfey+06udl3
KyhY7/BB9kfdAvFJAKYyNyvXtJrU7T1PNWYZ/1VX2J+QHF2M6+fc6UokY78iIr8z
LeeQuTb/ejHrxshcNoQYOFGDYVmaNZRyUWMjJzMcrpyD3HMLgk1qRpYfXtNyz2xJ
Q3jho5Ibxr4YhTKXbbgT8EZkeXHZFQ1R77f2CZQbv8tDpxAvUJWncy37Z1GIDZn0
rWn3kH9xpl7TNaT5lQTOh+HqA49UomCftmweYQgCv00yB3kabTfrYLhRMbzWzVGl
xEpfj7AqkDhhNxa4hX80/bBz7CiRtKtykqu5r3/tSaerCdAnjWwyAfluQu48fomR
Pnj7eiJWn+FSW9X1luYuF6wg6646XgR6pXbobgHvFCscbmteBFeCxqMVjAK12Llx
Y8ENU4WkAjftrcwD+PPk642vF5zBaMJMa740HnwEJ3kGh+WQ7gsdxjXB3Vpd7r1Q
x5pYOIqo2r3zYUiRUsMZ+LtnP9mJMQu4O1reEAgYMsFQ34IZ81F+VrlueKH7Qv+l
ysYgs3i9D/j2szZtlEoMm4XhAc7PI1vklWuT5aWJugRMoMrXuK4JTFz4fTdIRoQy
i4T35n77Myg523aVDy3v2ApA8wEiJhgsaDYv/AtZCt17q1tflQx7jsm0FBXeqqU7
9+ixNMfeTp1n0KQYDG7463mbGl9BgZuaF1Rp1422egELCe5fYyBZ2lMzRSNgLFa7
bUkgGiKr0UnsyAUhipTaM1TbS5l4Ht97us1cIYbBstHCP8CEpZeH3S1CsuDqltkd
gMS8D7ecwIo/RIIuFvCrofCZVn4+7UAGD5AY9ZKc4ZRdGSiFcObN/k62R3+j6GZP
FE7aDVxTMSnaa5yVnQZHhzkGj6u/o+jSqGQ3XcZETkobJQqe+RrxDH4F9ZMiYc94
7FxjcnmH6OXahH8ZC77FC7w7kVuh9mGwQIsncy05n2i0yKUQyl+2EbXJlFxTaQhH
BUhkuy5AWq5Ye5fLs7pbIafPG994NBQcGLgukxh1oGF/lpsxuekDrQNW4hYG5PiM
KTjGYy1dGyfs/O9jEMq7492oyJyUY6QafkkBPNlh1di3D0uZKSgkrqqVENJKxDtn
rfjf8kVeKxI5oMZrem6PKcioFvp1cDu4w5U9pxTwY3HVGPWg9Nh1yt0B6ALDxInX
oJD/ax5mcf+Hj4N8bFG8n3TS7Nj6l/77kmB0c3+js9dzMFnXFuZEsDaqABQo/uG7
Gwz0vIDF6Xefj7PMmxQf1QyS8Ge61c0grzLfPbIYm9Ytv6mZ0MM29BHVjds709vr
jXAbG22PojPF5S2jWAqUsHXv3Np6cJwHY394z7OWSO7v24X69v3EbAQZ3d6YJR6a
EwCULFcC/1DlShUGQNaROe4Ynthqmj0DBO285+/CR52BWcOC0E0MDh/FBfpXxZQt
i9Vj0bAQBvaQvtqewfBxwnYRHpGsDlFHAKCbeODE3M8Z9bMjNinnPPF6+qDxVGyy
Ozyy2CEaeuyYdtKH4oIlTlv8DAj3G7z9u5UblYgzf4JvY8B6bFvdI/goMwz4Y3Jl
zqYHJsDS9BTQ1guHjl8uPbXZSRPo4MNG5dL0uyVu6zdgGwubA47hPo4SGTKJf0Zf
jwk3Zd085AwRMWche0Fh/4ZJyjNft48ngL5eoMYL/nhxsrAllDwUAoxgrxnWv1C7
hGdDGxVm/b1srUDhb4R19pRxnhYeb+v62MKKCq5ojhXZHWjyH44+EQbAXLB+Qx68
uec6W2TB4fsSapRU4cF2rTgnkPPBuTijdfv+xwmWZ6ZvS6dN33rpF2kPRh2Ze8PE
MJvLA7kIrhVut0+sY9VsVkh4CSCRUgzEbZRySmCqvKgdth90xb92M452BdclKNsy
mmYiZjuswAxhCGiBt6ma1sXgNnFgLkG29r+AU1NQEUwqh9Gi7FplPeb+DP0we96z
NbhzI8SIUA8UzbUxCbVKqQeNv6DsY3OE00jVe4W64oITQP/S7CbsFZ8ioD04jjty
tmsjY//9NmDIiH1DGkNH7HvAQoMjmgwnM5pLcorNtRYnRXl3IQ/fOswP5TAIgcrG
ARHIG3ImhMwsTApOJ2U2zMbZIrIvAgoz7CYCZoDAdErL/ucrhzgiA0L7GL7fzE5+
KHQ4CnyQQPy/GUZNvST4nUDgh9MWWBUobryh1FP4GszDUGjNfiQz38J4cc7DPftc
Z47fVIxivifl1Bej0LPyz9b78vYzNzRV+3YI5AkBF+f8JQH2ZdfxYi85IoPFYuml
AHYfLvRhTHqIeBXeMNOglozBqNEUb3hTGLo0XwGMSGhHuIRZCDka0SeP9oyM9BrD
NGNTi1sDfymnkE80EmkTvKl1J6Kxs4glocopscx1TaiXEQtNGF+5QJc+X4NNkFIv
FmbdIbkmgzN1D2MBGW/QVS6AEVFwYU/2NGslEAgCStBKpRrZ9uUebgeKAumSqLBt
8xC1VbXNIW3QoHl2z0J1N8X5/7HGjVBYOdr01qS3ZFiKaiqH/k18D3qqpzasFlLN
3mQM5UsnOE2vcACTMrrYH9ieN7dEETMBceeXPE+7frM3srG8cL2ZoVSHAzL2Ql2D
gOkyCMSAAdYb8aoU+gLgYJfssRQirQzq46iLZbX7R4mQY441A36eEY8HeRK1nh2b
KuBdhH+YKAIDR0B2MaI6c3a0ZxZy3mZEIrUhUQvP1WIT0PxJhHU06hobGf5PZSq6
UNr5XwJKcDjOaZqBpue2vG17mVtJRv67oHD1PwBClbiGnvtNY03gi801LiH/1Dbz
dWKNBsSvxPNA5UPhGSIVBGlLM3ZWwiDbRiaXWiVy+oPB6UAOzY15I3H7W0lciNOV
QsQ2ijMLV70tPjrPUq6ieTLyj6VBeDfcSL0to1oFSsQuwy7rCxFRcieosAJAAmFC
YdBSoDlgMev8KAloK8qowA7ucJrv+/EZVOn8MjW/istLdHCa2mI6mPmkVVxHO56C
TWcRyMGotXfouYHi3EfPPTnjw/Tcjf6E+DXH5qbUogsnmlu/BP3HihVce5hDynca
40EJo28U1cazEyR7J/MudbiSQAwQHOM/Of2nqaI5jZeevJRh1700J40favYBBKVG
X4Kwn+FTgxufqoIjLrvbQc793rKtCfMenMfrHYqIObQKaFVjxPwAubofplfWgNBu
fx8M2+HCRSCuZQ7dE9+Vf5TtdhMtvWURmyOgj8UJ4DKVDaHRKbGzbD2gp5b2+SNT
8iHIpE6JhEks8EFg88/158Mzf6wCyIS5fDlhWbJST97jnAbbYanNsS/RMicGYk6A
ne7aP1+vnY3m/qWYYJHP695nVk7cJ1A4PWBQx8M6uvzO4b35QZuq8AJ1etw2jsT/
crAZXEGFjy6J4kwdy9d+MtN9MGyy1MHLSppHHlkb3/Zb/fQX0+VToeWzaaDBYu4L
g1cHPB39q/CTlD7hmTjdy3CuuwPtmUwYorcNAPsFg4IDnoVb+TOvUZ9Erf7X/amd
/5MQ4rtNbo/WnXraNJnNJGd1nAoU/lKW2ZUsqagDPbwwmmiq+Q7yXP1BxylbGitN
+fdsmK/HvT6wvnMSkQDR6q5ZGCahPqQIdYz05VZ3md+eirEkLo6UsUxma7CefWnf
1wKKfh3JqnLfR625V/4jAF6zH6vAz+sMQgfbgDi0tDuKeikYxp4o68F5YmgQXV1e
Tpb6TfL+ykaKinZ2KaO2pZDRQ9D7SFHsHApZTJHzTKgqLKYGLZrRSc18AMhi4Riw
+lCfI9vco4FDU/Udd/CHhBjH5vVi+wg/4W0ShUER/OJZGRFSA/WEP8Nwpsv/Y9vp
jNW+YYFzRc1vLYQoT6oGO6jrvFOt1tVQH54F3Yj2e7cuHUu6nI+on4irkRgP9nAd
knIs4Cmq12BhiuLQvvE+0gdL0Zp3hMGD3crp1ieCXpjwU09oKlAz7WI6IecMOfn3
T18bChTkjPVCHDVvohsOJa+VPt1dHVNWtQezOMjcWleA10Qxx7RwMWDeieULfLSW
pp3ujVj0a0bekxKjwOlLRC3DMvFxojrwnftc8cDlNUNrZQw0j7UjolXU8cufCeAs
acAEKKihIvlIOcPVh+9jLWhD8fzeqUih3O1+kQkSy+/lzr8coMZ3YmTf1zPTw+tL
zXMinU16fDM/6Ocq0x9CnC0uZioipipw1L6986uHewpRioQn8z57aHx2wZPX+/LY
Bzr2YoTH8EH33KgFjjdEqcwk52aHDo89r0H2cWwMRJbVTDsLFx9kcCOu4wSyT2FH
QdJz5Gh6E0Bba16DoN75pmD/TNvEu40AI6+D7U+bdcliJnj9XFtbx1b2smEPmUGC
oU+5Gcs1w4yIM/I2Igwvp8Xp3D4FAmQ2FfjRTymvTlLAEVs6fBDhG+EnE1ZBW1p5
BD5l5UDt6WlhZJq4QAd+vpvila4t9xAI9ehsNRKLKfI6GnGKvLIf3QskSKzAYOk3
WyemrRoAJ9de9GDTKDgC4w1VuV1qzds5U7O0Cp41UQ4N6cehUB2UB6/unApSkkXt
Qlh32BNRBeigjNj1hPWDCupfA8ao4pM0ObZCaiMww8pTYGIGJAM9gIR+KvdMcXYu
FqExBCJEp3jTWjps6LtzowhlJrxXZFYCVJfK8orrcte0c2HxAPGfy35m5eMsTl+Z
4ZKwLEiqsU9HbzFOycJMxS/YMcNk3s5+aizmqSUyk0xokGRzbhhrNLOrCBN4CGNE
fC93TbPAwkhzOQWkS48fIbgW2dPdbtX3chliI3EjNEDj3bt3K9rkJNgp7+GM/Tkn
LJtKXbvVSw1GNbatte/45PFEUl8gFU/Gs5UouB/weOqxxWzSQOFXaMfGr7ufiExD
47eFNIHLfN8lOjNk0D6nfKvrMBXb7yRfPk+fdWl322t+3k9CoINtEd8HvGE4/pT3
oHlQ5Zm8b6SlBREUpsES+UEJ8i+cH4gTbUlwy2uSPpn+/SM3JNq48I1UQwxv7ElE
uJjj1dQFVWZ2M6CqjDRMrUz2mlF0jXu6+EIJ+TD23s0154teysa3RzPQvvFFw1eg
tDziJm4vZbSGJqkzhOiMwk9poJo/eCFxM8HWRsuOQNHrkdEEQo1VOSW4UQZXFIyN
5gW480YMaSforG9A5JWZl+b9961RnpLBO9IQMvjw57x/f2ekd8SovOBSwsPrTX6J
lXedy3S3Ku3kVefKGIfiFXFk9wD6j3MkCKuLavh1CqQV2zY8SPhIJtW1sNGCdVwe
S8sR0BpWkgOWJdwsmnp6bdjhc9xfWHUxXWMElJElQQriNqVhrGt57o/vVquiUfPM
Otvf8F6SW/Ao4vJCc+kaaAuqb2VNqNTr4JZPgLY7zClIl474ri/HgbGixmkUNh/O
tL+wzSNYe0Ur9ca8gK7LqKEhv8ND3qdq6jJdeGeOMCQ+NI3uuLIOVC4TP2LDBnmZ
S1pjsTaoXDJHpMJT8ecEfBI7rwSFM5/c1ucxGR6AtY/gCP4R0CaiFeaQgjOgR5wf
4HsRNlsTgmXOc0qguHGWnHIc+E3BgbHti9XoqmjcgeSi44s8WlTMkThBogGPG6F7
n95REpQ70XkvMB6Z33jDGrmwHk+pS/EKB8JcOBmUuKe6SDWq24EPpR1SB0wULKb6
UqV6K3vls9fh0M8ccODOK24sbPmQ2RPWfjnPVaZDKnfZx7MxU2tQQ8V/vkhJqL1U
MVJzW/U5xlZvd5zvcRK/0dQBha+AsTAjaytxU0BLmeY12f/+d0TyeawFhB3XoQjJ
sisSGWg7yc65ehAdxOyNs8oz0ErgRs0A6dPSaqQ7/9DYVS3l6qtt+emBVENEWO/d
G6x7tCqDJ8nTMGol/GS4uu/rwCviyE31tnTLTkWoGcx4xtUQrHDrt6bpg0zma4Mn
5dzGlsLoNZPD1b2Wpz2+cb7QrGiwZcG6iWxmofi5IPTYzqWdqXFQLVFOA42XUYnj
qmNArJ+pQJQMn4B2EHd0mJJS2ijveBqEa/fU0SEMhFG2QFRrblPLmYY1EYon/R5K
vbkHMsuAdNmJf0OWZES0uQmN+dPwl5EFGYGn/1n8o2qyoT++9PpJxY/PrTuoNh4O
zgPjkUGoy+iyINPmYgO+Sd9hCVpCN2PlmZFhST7a7SbrmHkO8Xikrxec+C+/6SF3
hzK/H21PMRPbt1ljwBSi4bc75LB0xdof2oY2aEPTtADoHEnVimTed/BZV9AR/H+n
MZ2HtZchTZ8t+vli2ejhjhpOafj18bzuybEHG+593wNawtA2RHEverxdkFiZRAgz
HWRGUbLTf9hq2/rMjmJs3UlFR5qpr2l4bsaZ8Mfiqoq2ISCvXEmd9wDk46W609Xa
69w1QakfvIdr8QPJOEZ/V5bOf0FzwFs6Feme3JaNwMyYn/8xW8J96byp9+QpfyWF
ikd0kEjSPX9d/ClpY/TuaydyVO5PzI3i5eG2mFZEe/qMLdHbrAQyuipZgFt+RWO3
7nZPm6WHt0lukPu2P2mgIk7VsiGpYxEFzV2Fa09ZT/lI3ELYjfSOVLwZyNsWBWw4
/VUQ0xsiKxuzapMJ+5F6yvFnwoBjwX5WtgEkuZwGEQLeOl6DBFkabLQjwS2mm94T
ySiC5yX6pc1qirOS8Eegb93+isBw70Gi9zNUBWZr+uNTAtw/fozjMwg7nbOF+t3E
1tkipefAzpHciGrJEiqv8La5LGr+dcytkCLkMnwe9EmVM/0HbFTf+acJSstoS011
0kY2Qtd2oadetJdQAZ3V8TfS1N93TAXkalkXN5GgpCTyJE+q9GcxDPvbQ6slryR0
hjqnZhlOXqby3Gnxex/YZLGoccWM4i//tfkCEEEEUR52qiRU3w9EXJSek9ER4U/R
nJQyWdslkdaQlM99CePsUs9Q2GHy6UBYXZJGZAA5EFbhf8jcUh2TOVy9tihucKEu
85x0XG8CiSkwtIB8e5k4vTF7wxww6LIt7c0mKK1jE4uiKzIWLF+B9NuwYCxEjVHM
aebfFjXsr7jYoLN3nPmIUQFMRwH6f6X9agS5rJTvSZ4sA/1zoykDLev320ryx0or
5ydooWHSk9jKgWSeUKgWEc0x9AHH3DER+/mwqTe/0KGnuirGWdENe4rYU2e+PXYA
RHAbacozzavsvGb9zGTG4ONse5cJmwY2/Unma44tWbDrEFivZLGAfCYBVxmFnsfn
WBs3s+zpuGpIaG3+KG85nO8Ak5hGMHAYegJcMqvLqGo+QFiZeXKRv1Nz0t3pnClx
i4Ol0LvlFHFC2+Pjxkt0syblv5wOV7tr/mPoMusu13ehUAcq1xffFTI06ImKthsU
DsPd9hXgHek6V1FiXG+8QxGHxTjcd1J/qqh3fUY3mJFwxDmOUDStifuMrrrVF6aa
XaWtJmwk25uAUAvliTrTGcmK1f5WememhGYeVfVOJkLj8fgYmg+6lWFfH7g7zkQm
XEYUkeV1Q177EYelakukLELoIuIgeFmqWxotA9Y7n7+3kRP+Ci2/FZ/iFx4Aq+vt
QR8G3VVnl6UPR7gqBoYk0FYDWQdXMmACHb1uG1val/rMpyScFm4+uLS07rPZxmXt
FhxdQvT3IyH0Pgros7cIWU8LWezucgQgVBnJCIsoo6fdKVdODOQrvI2RDU3RWOzY
dCkVA1lUi3I3jbkNDAkgFPVoBqr7g4thda8FasUfDRh/SniPCo5EqZwRkkUkv3wN
ww1elKF/XAjDNim+3uUkPu165JT4lcgII2Uy3Gr03h4DFb0Aid9c0Lv0cvyEkkVn
9jQbByrkIvqw1N8YS93QX0A+k9BEdSZqvm+Fu4XZBNcbMHRH2uH5HYh1GR4XR4Je
B7pQU43i6NiG1uslZrer7rJSoiKmMprE4r6Gv+mJfK4TX3uOaZN5wqrAuL33hQSy
lQgI4EP21hT6xhBVUrSlRWyk/B5ArmwzZjKXjJGvG1qSDg3U+NxvMRd+eL5nOmos
o2SIqjFUQFD2NXcqew1YRgn9AcrGUaFcxN9oplWQMx1MQL8XQm9TgGuwO/GWaOJA
UDnVZp/Rk7X6mSmwas999PVcq0vGZkNOK+ocOhCJKJFSLfT6xG4qrDye8sc5kPsj
6fu9flihHkv7VOffi+ISztfIavYgoKg51eEkYstsNATImQPxwX8HRwO4T+TOC62t
VxZW09fBX3wfbhuuB699ZMOU5PuzexA8Y8j6o1rMiXJTA1pvTXon/Wh+mOHneY2Y
nP9nBI/WvHNX++IKDfHcN8atX2NT6D/BPgGtdYFdvkIrjq+Ilyk7CfQ+Iov4JorW
Lhf4WnF7Z0NGJlhq1Bb7mfvVesWTSfxRjTnRIRdGKsr+Wcf73bLh6aitk1dDGIde
9zq1ZLhyndLheKl7VEt+xaojIlr7SELZ03MTtstiJr8Rm7Ci0dM91ulcvIBr58we
a6VlNe6dBv8rZfeHethr8Q1Ud5/rFHB+DsMC+vGRs4b8k6DdSFEpc4KBwx0mjT8o
xRh1gtxEfN8big9r8bEbSyT1TqJrpYZmpyigRlkq4+gZ+vITJIWJmHjfx+KN7qEW
M18cSJIAa09yd9fpM/UAqEnquxLLWNyPZ1LaTEl0I16T/gT4kAV0p6aGZPiw4Zsj
uYln/91uOj/Ub1dUShXJXYQkldILLE2dn5KQTkI388a+gBhztkdtsMSnCVFTxKND
/lyXJdGyjCbPn6aKE/qTp4ESJXNo+mQJo2WCq3xNeYrmEStifBaDKobeKtnUeObC
xJIE0UOG39+qAMyWolkN8RlkIaBHP11RhwGfZXoesIVtgXUyZ59dIjhWNpZ+9q/L
jXCq/YBQKeIuVXJiGepViJ6FoFOa8NJqKm1ootHYU6N2/rptpwnXRVkWdLGfk6Sq
mfs9Xb3SLfqx1kz/cteGDqcbCbbbVXxo7kfTCgcu83Qrn2ezPZ3dTTDUT+kGNpMf
4QxHWAShDeRPujRb3N7P6X6qq3VSOK+jQ0GZ27UEN0UmQzcJzpUOj3z2vRHROG4U
q9fzUMwgi7g0r89CLa3u+OIRJ4zc1aqdkL1XjVrTiNNXsYlS0SQZU0CfLl/HQp4X
OJKpH2bXp03A9SsfHXdlyyYyaO0aGh3KeLO9CIaCWqBQsCXzd8rh6v1bfSjAiU5m
ZMqGwQ5q7slokVl93gJcpIcdG/PlgZpCaL+KXGKCAuQ6JTaZ+MTtKuBl0li1xTEM
HzNHtBKfDR5JxXXlByVL1eAG2xjbBpn70kNDcrlCJOdbS4Kdkf5Rvjh8bWSyQnLV
Bx+y78+ZPpFam73WxuZl2RHShcKqCIprCSunczRlSH8KfgsLdFsMQw3YLO32VoDJ
6vckQ9OBZD5XqbzLDurc0s0/pLX2e+xNdh0tq0vgqgP2axCD/HLcH6EW5PPJhMF/
LpRG/OQb1b4DK1bQEppuPr+FSv8+oSm9LFgRqYRJnFaRmhW+JjmVvyCr5CfFksN3
qpRlO+uZSfx+Zz+s5iQg/Q6RYMHaMfblZa6bXsAUSJsC5Aw//Dw/vmMNoEOxB2zz
EoVIlnJV5vrlle4pUWUqz4AM9YAK9oDqoIGRgAMpIz3OnBrLkktFd++bAbagXKpD
z1EYtn03OLzAlst7C9jLUkO7yg1MtLiUAtxyTVQIbMUcrhleFHiN986NkYNKOOjW
IM93fTRzh9xxKmtIIV36sC1Nb+t1Lh9bpRV+83TY94zGRo22TMyYIVjin7pdbhyF
a679+aQb87PZRVrrIzfNA2N7jv/uamcQIyVjwQ029KGj7YYx7rGnmThIghQg5gN8
qx0S+CTle9RDNUwoujIflxLmaiQHJsbu9NXymrsox/LvRemxPapfSnAzF/FP8HZV
o27FubOUtlML2vH0gdVF0l9Oim/aBZISUmasnQHwrj28Q0uK8Sc3sPmJF530OOCa
a7leeTeI9pM3Ojs7ywLvniHT2vxkXJFNvpn/SVZJnue4Uk+cDGHI80nO7w+JU6wW
hOZbthuZwvTS+mJGPsG2LFrR1iPMDIs05dMKn+wgq5PITPQ+9ouryMPvxcLR3H4t
EveZajrlWOHrb2enRNeZ+CaZqR1DoL8xSiwTZO2D6Psgs9i3V8wUet/XqgnqYIQY
eurBEfXtQJ+RSLuOe1cZCLDOCmKa0Qb9IMl6lqUTodkntOu28Jlag5Um+D3KFdzt
MnIE/6ic19o0mO0uTzZMYFsDpJLuMy83Yd7BwZjFV8HxiYVFlc2bM3nbfJsd18ZD
SBRX77OzxJHB/w4ZemwuzmAeI5PGGWIN0xkOzGxRzjCCy72y/bHP7i1SxX+OXQaS
Ty7Xuluhhh4VJEzBz2uZJj7rPsyM65D9ZQMvb4nR0m1G6VAFiHZnLURKXJn5uDql
qPpekVuaMQZHQDRUa3wYLnGuTEDqkCbyLouFmSLBsEQctEHqOUH8CK/77aBXmn3S
KZA5zaVhe4d+DcszbAh3BhhvhjKxucYMvk1vagSG3tNX9G02J6nJW8+6cZ0W54Ol
z9ugKPeaAPQEFIUbbFPX3FQkcIde31eL5NxbyaeeOqatv0jqUuWPyw3VwxGLgyh3
1M/Nk02Ls41K/tZpvf6KT5ldqV6yRJZ5JFc+5CYps7YxhC4xFFYePEMlFZmZA3Ss
KhgAVf2Z8FBd16qJbIvQLcMgX89Z9tUY2/VZnysYf24jVwPa6fHN2EvH+cZet44i
ceyJu5FmvyJeJXG6/EpVWw7KE5ixoCRmpRzfBHQHmqqbu1BSepqu5sSZi0dlJfHp
uwJgsBhIiUY6YfuRtcsrXnWltjQKYv1MhSYUJk/9cn/mq9JpxjTx8s7xbbwx8mi7
MZ1zLbXa7kNA2VSMDPIL+/vPm1xDwIoi+aAaljXH2/mbNTsmBuO6NBk+gizT4Q6h
Ieyb6OZWgPpJb54qUl3EA0zw+7XO9vn9iRYFuQtmnKLe23+mPFFfzaJfMPl4DgPm
bZhZEYmCEUzGgfzU21rJMcTBUFfvDJgZ/S+PtDP0UhRbOA3z6EIcpCQc5bZP43f8
hmlUCWrWfYI53Vd87TtwVh6Hu1+Z2tR3/74AraDhjU8zJXhsttsrBFeoqW8Xz/vO
R0CnbYpGbTghm6LmDeCcTWz7P7MZ/Sy82WEV9N4A8bOyRBY3y7zqJ3m8MUSGam44
Pgq8tdSbMI85pFJvDsFQxscRVdGnNTco0UlcypS42lIj6jG4/CWlJR2muQJjBQoO
/DAZvPDyQvvGGzZ2W9s8EXyogf0e/9OAjRtPNbRIz1SVD9ioFrL8R2I953M/R9g/
EPFHYD3Yl+lz1j3bpD8icI5zVgxgk+9+2nh3rBJPhO2iN368nlG98kAaSNilkkGr
VHG2+B/LA3P8ikEdNn6roOxstxdbZsUS/2yWPsV9O8rAJ3EjWnqhnGwfztadaFBw
fTMus14et7tyzwFI7brNvaNQUnseKaIuytL2kGgYdcUdu0pPsIZT0JHHftimZKAT
MwCX76YksDgXGPPLjr9fxTxDfg5GDXWCP+66sA2VaQwP5z1FrAHuiazuqAR+702e
Y6mWbh7XLjClL6/5p8++purevGOIEt6Fu2OH+H6GdItdmXs1Eb4ZZn+bM8SN5Tt0
4rABZF/gKhLimKRJRKPF4IiSWGLL3Gvz9XplS6JgyFfZ/QbZGsyulJ8g9OUSBq5Q
puHp5FSeNdYUQujTP3YF460cm087wFk9v2hKcqpgrTWwF4jQYtlXKWkJ7gdYOdIr
jKxtXpuedUCMGOWg2KTRCHouQ252rdzZ1+I9n8yNqCKuaRqTE91QFAyRPj804nWx
SGv4bXgDhgmBM4th5IIPMG/EmAGGPiR+POyYp7SjeAnkiAjoqmsDRxNZqKcRRceU
Ua3haCT4P5kaeNCTmtiN5R5tFAespIvqbO7TudARmPWTVn/vadmo8jY8IDyVr60n
2rNzvGTgLRTE7dvipYGd0jbsT0KRSu4SpthNeeJn+ZK0PlMjDsbd2NjdI4f3RU9O
afZP4QXU4xPBP7r0xWKUG3W52Cy7vS2+g584Q/UDBDnD7luffGuvShHkZEKNx9yS
4bKV9gFFFG0HTspCRV2ebhAXiFkW8Tqmh/FLb1OYm+LlWPPVRUzilR9bBtEOPeC4
aAbHWX3ne3dAa+MwBaWIVZfF1ign3mJE32JQwTXZf/Hu58utX4D+8gjQKCdNqU/W
pQprhI4UymekV7A0AnzCW2bFoE/RMVF+oyvd+VxCos0dUFbhDUobOHw0F9+f9gLD
NW3hnsPNR8mIMrVw+PR8EiGYA7+PQGauQx9eM9BtWAXcPT2n5P981Kw4y8YAa4fU
unFtnvO96TOvfBjtimUIlp5vBmTf85Gdqyq5/XH+PTuKJiXZCRUlGsmgb0L9pa23
jY4vlPhYBp4pIUz+otgADl4+YcH9YcBn8mrBLJfZOGkCIW5fUPsr++mvwvoLa3oP
m+XoOCpgekyUAwst92yRD8v3Yy0vFRutYRKgkwdlPYVcigFCpCBl2AF93dqRevYh
ThQDYESmpZLkmHUJ21X5wrJ3DJwniG5xtSKyMqHDF8wJhE08l+sfHca5AaChZ/pR
Pu/EJKR4nzN295HRWj04lc5GxVTSQa7xbFgTwaKu9Bm8m9hkjhf0mpHZkZ0DfG+x
+HbuSvD7FCqK8phhyqo2gHyBsukx8dFSs3aQ/fpBUPVU1KwWvtgXhxc4xdW5Mkfw
RPBzG2g66onmYi8TcrNHOO0BI0xH+ez2mG5/Jh/djF3zwpzCgl6cQkgQA7TcS/Eo
A2zGurnuWlUZFrvCYykis2FSdc2eqXHC0uSDLPAJxrz6LJFP7sVtgzqSLnHtyM3a
RbUHrH/HzjgxEqfpOzXmiTQYbJ8JdvIq3F1V6ys9YXjw5GTtkMAwWtp1W/M3cvXC
GOkxOtxgsyTfzy+BgnPzKAKzNSqcd/kL161XoR91swJQguPiW5Lo3XATwm9Oc6va
twWza7tN6AWFzDLyaAMKWLT1tF416ujD7qpzIMBKW+oWTschuUXp8m3W7Y0dFvEd
a2uu1+PgZDWOOZGJQ0qBam3jbftwDU3cML/pnneugcIArvBwrUyvQGyFBGnxNGBh
fRT0RPwqJ+LaPGpS59tcfsGJtG28dhanv0EvvYQQCr8022sxCHhcuRYYr+FWhWF0
4MZD91htfCyIkNFI0ZxLs1Bv/wHkXVkKYFRjIGZgJFY/KIouZxpUrlpjSgDqQp89
lAVJdULJZXsGjapN3KMvuPPsA/0bBG33/1EpJUmomNzfrec0kAXb1XdDgwNVWBmJ
22oqdoGXDqurCCipksGYmI4VTTlmPtiHV/C+My2rBGozISE+I7ZbuOiywiGcQxCc
JbmiCdTdCkMqFi7fWbA+UXx65aawW31Wi/Hp4e9+ZVjvIlakElJ/Lkc5eJ9yKmgv
3qNOVuc53L0ek6PvQm3jBqdRU7thUJ3OI6shKzIeqwzPsh0keGAE9LwbQF6PEbqN
1WkoBWvdYjwjIOc9+jCjXOd12wvnzdvHC9o1UuO8V8B4tOnuVxkWD3DOL+PdCpnn
EG8LYVg6ZeBX8B8khbWHL3Gu0/fZ5vZ88aAO/YKkzKQ8u2ipyNKvkgz34aayrAJr
oZ3X2PCsAPN4J6aLgddOCCBw/MnrUfKmKc5p3D0au22GcM2zK3cIpcqhrynfYnu6
b1K/Tl13URMWjRFsUjPn2yWJ+IrI2YuubInmDo+1lvqvMiyj2cBjGXvGEw5wmiUt
Ze6a4ykwqv867rgdfepUdiMWCG7r+/7iRhxKKR2fas3fX8BzgLm2vYPH68PeSmQV
r7z5JbTTBozTwHjeDqQ5TfKHqwHeAQvp2sHquIU1Mvew+zcXV1AK+ir35JHKcWpC
dUOC/0QkRjBjyb0+vvBrQLnTEdcdwIzjPknrA9PiZAJOYIhCa1WgyvqoBJeXEZ7K
uEoddsIu8GOaZIgBsXL25DbXmhhCWvYjKOwshchSyuKSgg1aWu2wunN3aoO3/Z5i
g4kQap4aJ6ShjR3a89jLPxyKegx/QCg/bMJ9wbw0LpXapXHP0qu1ELxDxYgorCVM
5fTEkY0jhkk/OtCPdg+ZRuS2Y5ZSJ8Pb/cyGAMQKrxpiBxxkFON9cys21Oxc6qZR
lfwg0nfUXpQnXS9PiUuHPZwIgj8CmSfWjJkTzIgr3GFZlIM4ZKoYkfLP1lH9ZHXG
Z7dAmUU4WMlqkQ14HwO6eEJNU9UkA4ieg/HnufmiOCNj6cgO7pDnUFr6ibBE51dy
opXIe22+vObvvwwy04hxpAxHzwnpnEBJQAcya3PyGChmh/tlwWdaNplqU8EAU+Ce
1zL+cpujdTUzaPnmKyGSZM+UrPitUoNfUuUgKxLVQShRZarOR9gMMIU7g2UNxcmE
Khfeq48Sjkx1EDe67IlWBq9WmP/lK2lZYUzaR9L3jJ2IRUNj30aWOnO7CFz3d0/S
qUA8ylXL+COHI27vSHqknOgaNf0A2xzmo2wBFoInBkGOGr05l3x3IxCD85Fn6k8S
Sgp9CNqM/67uBvRHGBeflRWVxX9TjBs8hWn9Bz7ZQ8+1qbA03/gD7H/Aw+JkGLyt
ony1t0cipoTEvMwYanxsmzfj20RnT7PXacfW/BpsnUSkbeiBp5hg7yrA/cFOCGif
Woj2JzUdR+5Rz2AL5c3HdyCajylqBsBXZwR1m1xI1fhcSnGe5j8ITVroVs7ZYZTZ
8RW5hLQ/Gv9h38oPxcwsN4I3ad86c8VFni4KD3ai1PRW0tVCjcB5s5mGNqVmjCpb
ShGZowfTu6nAvGclhCDHDVJMdoP/HWRFt/ZdPv9AdjnTPVw9YrZ/TYk9A6yCc1sT
laRqN+PKdZUFv1QesOEe2eslZCDSiTwK14DH1JwBhFMkgoUeXxjk7UOvWjJX3brq
Wt1EUzxYRIUId2Tz8TtmInJqxLokAtvvupx91uG1Nge2Md+33yXaHKk2p1MZtidH
GSMLYkmtbGIuXK6MBlhd2rL9zDQRJ/wDdYhwevPoBgMcruI00S9Py2jC8Mm9Xv6r
w4lF535rcA35kKIROZc8z+8BrS7q/KOOSsnUBLzl6ex3RsRDB9V143OAhktMs2jf
PiPqq0oDqd0RBoTZLoDfkDsCF8x+JkhQEJHZ9SyxPapEaK+sz/5mMyGNkQRc/Fl/
bJdu/OvzwrO94RntC48n9uJps1cUxyFat/4zBdGrWhW1K+KV9QclShpUgQe80zlB
m/d/6YfSr4I98g0jwWG8OCeuN3yAa1g7dvBiL10VOc06PUGBI/MZlEEBG3hZ0kL5
hkVMOpjWZUODr3uT0xQU7soH4dG9m3Jyu/gvhIPUOty4cum1LJ4FhsfqimAf5MJ6
49/3xwGhtNbhWclfzL5vn6Hk6Nz9FOX9mWJTpd6IepcYBHajTI+lMT/CspKoHMp7
CETB/ZtsH2jDBagm5p/oRMi7LVezt/5M6FxtDwEpg8SjVEkv5yrjVxGotRETDcVU
R/tH/iDfNpZ0SZbL04O3kTt72Y/5sjkwqsRK1FA/bYu9ZkG0M9IcVByQhUDhIdyi
GxnDV95FEbNKzpWQR/mJCZjSPkjiF86wzPHewxYiqJYYZdIUqWVLuLjTxEvf9ZCs
fAeQt0P5BFlqSBkNJxNTV1rgRvJLsdQw50LCS6nuPuVGVOiTqqfX6Y+qino/bRJ7
+bBIsX7L7hWx60BI/8z86mXrEZ81FWsUcoaCW3eu8nt2S2949xS29Xrg8U/rElPd
Fc6vS7UNP3TAwiB1uPSlyLtT6Mg82lAP0Lhy+NhgaGXoLq6aBFrLoaelhfvx1onm
vApOoKVkm+yu0oEI8J4ANhIfRu3T5lauBmraFDQsj24BHuMfv6n7HAQPiGrhUwcU
iL5cWWDGbNIWRlB2/WHZRu0SAOab23ZdOTQ7ywQRO5ZKzNxzQ9IpxVRhjGf81rW7
nhMzgqKKkhktI0ROyZUPsnZEL1J93WN/92yLHbV+elpAC2LrDVz+ERZEgfRqJXCv
Tf7cFD1q9Zim1EhjZamKgzWRq0YxGkjj/2U33e0u2rwai3kWTX2/z/psrvjOp5M9
eIsVb1Ap7bVmdh9mcvMjFemvrRh96sNgfGLzFDpmeSqSwjh1rKSL2q/rVRBJ0o/H
SP8RQltEuF4VYSZ4Ypi3utMpnE/mEOhMYVL7HCLGi32qm3T4sD5m1WAzLPtvBBuG
KbLogKnwwHWEabRUNSTNSP0qTxmyOoR9dVU04+xSNyOssX1DUslE0gPwt1cnwINN
2gH6lBAmhLIsIzxhDQs8Sg/NbRWMl89RVx+4C0Sl7Fj+z8EwvUIswrxXZZEuOBz4
lV7EQB/yg5VzLsLIijqkbbwJGsEPI9A/z7akDvY7PsX2YB/xqc071eL0AzDDmdCu
pcd2utziHHiLWkgzZo+hEVZVQP9nH9DzDCZ7Z/MfgH6KJyPfMin+RyNLWD9XkoGg
BT2dGd5dT9Tsaq40fwZ+BmKAoX4fN0aO3w6sviIplqpevG/GuT1c9O4W7rQwV8O+
oI/EH1M7+e18HOSrPy1R4KCjkp0X+C5/J4S3g4+B9mBzAlbam8w4ozSZvxjgN5F8
OD8T30fXzJe3+lyyEL9YT8GbehElZUv9MY8xe4gz3e/wFa/8eFDNzc+As5uqspXQ
/BbMY1Ff+TedKu5dD2BN1Rh5KKmCvIQ5KeiNIvq+7VF9CYY3NxYfzmX7dHmLGcSl
BLtwWRun3Rxj7pe8AChggCzXMtd0+tjnA5Usd3TbpN31QTUbmMSuVr2d5sscDiq/
wkzAgVANU0Q6vYZCFO7CpnXJ42x7+wWIQHpVXWdQXY/YN7YTxW6hAi1Iiv4+vrbR
fLG53mDJFuVPdb2xXXci5Fo3oO39OrLAx4nyTQNgAu+DByexDUjfinTsUYO8qzZt
mEOK2wYpzz1rY3EGfs5RCSeBRaXjzOkLO6rw2lcu6073nnu6cBGOgh8tzeeAXMQu
KENoTJvS2mds4jaVZIWQVBRccfEQz4iLh5/JWxEGX3mAZVeGvw1Z9CrKHJqf56rb
c5d5GEnzRFNNm/bPFp8kiA7smg8AzTVai9VW8+CMZ4SY2gHjMSHQsHTBQ3O0cV+u
92CUEnlujtGkJxx6INwMQ7T/8q5wnj970SGZ//t4TJmlROWRBaiYgmBJY2FkycVo
G+FRb7Xvf9tf+ysrsC99ansIWbDrVLrcBiduScvteImBYukfT2nbXnCs8sO5MRh3
AHjQmORBgJvgXWUKZNBc/MyqPrGdwYYLGslcCWAFMSz66/rFaIuf5SxN4CgJTAGQ
NblVPRifU+ML3C/YWX+UnmwQShtkFOc360XKHtxhSAbe2QHnR7b8jb4qsy+HiMV9
B7xJo6pDlyNV1KX0GqycuMMsZG9NEdM/LQivviVdbX0fXeeYse0X9ECHsquNz36Z
TLIj7zD0q71s+XrRXfY2m3PYEmZAMQxpwbBCTTYn3BKbERN0sF+tUeV0aUCq9wWT
gfiCEAP2OdW9SdEe2fRS/mDXhwRh3T0EXU+WFwHoamYX+dgsmy/wzB1gKZdzU1rq
94olhwn5C5h94SCsnB52j6lM3jaUgGz4MPciUkgl6soOpiuO2q9iWj4PydKg5H0O
es6yQ70+u8kb6USDpS2aJqDjLIoG4s8yxKNxFyQ0iyLAEZjN3KpEqYe2YuHYX4NW
qr3/+2vMk87GNnxigI4L/mlDenBPxpYKSTPmx7n41BJlQmzH/eHlscSw++cKGgyf
307UJvGfffjnoJkjbUXgNZWqpUlo5Xt6bWwL8dB8P7vNykZhARDNPWvpeO/dpMLf
GViJ/aHRUQ+Vo0eAeF7OVP8uNz7l9enl12CGk1lb4TlFBhsD5UPw97zZa+u+Afln
5ffNiPyadBuq/urH7f+ivoSwjise7Q51XqFHklEdcr6Qo8LVdrH35Qb9C/u8f52t
/xMJV6lmnrqJemfWet+ZygfiVbzqawnsimjeFFEHv/qwgYvIOHvhQhkUJ7z2yjRl
YD1F8xll9KRWJ1WLlcR1UP2a4Orn7Uy8AOMh6zq7VcuFYUG2ys9zOBlmWHgpcNn+
WLSsF7wXmBtgN6JXVBV7l7PXrOCdzawUvOdfzloveXWNgooiUl0aUD+1tLhaiivX
KoCfJCMB5JoXLFkwuE7SGCi6+4JuFZ3oz31CPewYpktoIaUu6n/kZzz4hcAw6677
CUcQqgviBmAHb5VUihDWAyw7NLcybI5AptbttEXGOAhRoG5Z3eHOYVkG/BMOtabA
rNVCzcycYtsPCGbZvN6KqnErCmtArIMOEuCnSL3tg6L642EirkdLMIPnrfnE+FUG
vGgMRZKQ921bTJKBn60HWczsJIeeZg7H5RfBEgGaX/VcBnvsIahRacRG8AZCdxhm
yAVuPsAalminwllNQj63Ze7v1oueDyAVEBRjczlqTA2+FTuV441y2UlY7OIgjkuY
aUGPy5HnJe6//xyYDDpJAxOQqTobIsuoTOvg1ABCQnY0m7o2hOC45guby4KN/9zM
hl3IJiBIHtfOqu22quJ49PAbTYWzJiAzAzlU4cBzVW+PLpHuUMDqaCN1QpYh4K9a
ldcrNZTmdsJ2f1nE8HH8W0e/LdFmK3gEzd9QxugERGhvOQ+LwycjE/OcI9Z8xH0Z
64vo0tX1SsTbczB/ZBcWpWJNIqSRaU7k+IejJheVPIkXlHAajS3ZDakI3XY5oNlQ
iIMr+qcHQWV1URCpKy0Sg/yX/lGa0kN0pP8T66MOhoJXufODSCU4uCO9oq/DaBAM
gI6bLN8lWFxIRjUOR+/kvDfmUp335yTfCNjIz61zB2IhdXFSNZnvdLlUcnmE7ip9
Z5WUFXO7xxHBL8dCgVfsgdIsfV4mv42KUzkBtgTVszpokQii2lxBspxWiNe+RsIv
EY/G+qM7vIhvP+aqibK17M6B3yl7b/l67bctjUMbx6YrlY3lhCJsI4Ftyzr3osV3
DhXV0YN+puGfxVy51CmleCe1FGUucIpBqajpCqESYAfZ6nzizWYPu9mdQgAQUHUm
+vc5ZsrDj6QGcPDfkGSaaKWLfeN9RaiIMROuqSX+J61sAZe53NK1qBAIFKaCZyXi
XNyuL8I3M3mQGzQzGhc+w6qOfJGZUbdpUkp3msut71UAycRXDwmSqGxXlGoMuYM5
F3fa3dzP3HGvC7nv1SUYXDMWm3rKGuhTgFVBgoULEvNTvpgMqNw7GuKMlUj6rau2
FkPvxlIL5mVlEyRMVot177sJYpK0scc4ys05OSffAXrYdMpg4MV8nfWoWLPR0WPn
mqR/k4rBZ5PGTLyiq4YtTbf66gCLpcb5XVz4H1kYANcbIi5wvalMNdXQN1+shBxM
aX7JOPlJV/+k7yaJ4+kF8UtJebFUjZCRBgJ9xY4Y+MdW5z4mgrc4WJwW86feBh92
By46BrwE379wWk2VWgawMUsWfjF3q7Kg5NN1hETm4TtprolKAB8/YTxdji7ZN9yu
ZrD7eR//fj5AKmJvdY0JRI1xJ5Mkp1gBU4kkSY8PJFDal2oJ6/ruUgTa+Z42Ywpo
i3O0tJ/Ol4DATdmI2KwKlFZqp/oOsTuXwVxw8plQPlZFCpPjeiFi3DpZQQoaQflB
jxDvkBS3rIrlfpUWC5Tgn+CanQ2EP7RFMhZ5uUGal+Qt4Q/npNZOFh8pZlBIliZD
Zb2TVJ5W9ggH/his1PGNjdF5EeI4zF/ldxrD4Q/nVdCXD328gBrFiVDScKhTzLAz
4AGL08DqWfgjwNpnkibY59mPtwe0ZvNbfF3mp35bVc3bxx7q06UuXFHuIjrvUrFs
NZQroGrPTjDmT0Ewoq+VpRA/zLA0aQnTWFRpuWDyxmoOqX4XEPIoeHxY225DzY0I
UTzDBQvlIXJyME87W5ABGU2KnAsP45885iBOhyIrt6LZJg0iivynMItN7/9Hhs4P
MaSK8sQ3KfcZ45OWSiZKdmohPGQmvuovGuV1ThvKC7B4PtxgrWtklIOXGd//fcqF
v68GBiI0qyBs7otJwgKEPcD5rB1HC5PkZ8hhORJzzRbe3Z3YS83ht51xSgt95AGi
NeCsgaKMQvKoQGw3DoIb7gr6TMpWV0SNPpneXqPozCp05zBwpB00AHE2l77VaP5o
K2z2BdID3I7XfUNcEnrUOlMIkOfz4pzDW6jaanOfQZ9nq9DZkj8D1qiJ/SpBEA/i
QqpmXBh0ISV0w/49nz83xuRP5ufC/YSFVVAb6cJPcAczJhJkzHOerxGnW9IpT2fp
UBbLtQ9+csv2/mXqOI1inaoAwYvu7uNq+YrbGAs444+5kvFQJJKJ2XtaIpK4b6aZ
VATmcYHeL5VirXiOR7Urm+oNTUku9XBKH5//9nldovtogF7y49r9alyCBIF84ezT
1UhVToHgApwDmchrr1tkqBLObQDy04SV2nFfNeQo07nxkrh0xK6S9TgLB2ow0aSi
WbeRObUkoihtkb5jrEJPJxAT42wyylaJ4aT/kFOL4JP2RwRODj0JR0Mg7p8yZWOe
aatZVMQuehTFa6NQVHhXcAHIyQsPWgymAmYD5ijwRDJM8osnX2GGIwD8tTqt51MK
nGfivL26PsyNmFSwtQsJQFfQzAXXbPQGqLn7NXhrFUgd4hl3rS3kfN/sUHonDLC+
SoOGjdVbc44Rh+VsLsX4Lv1PTY1JphKR64sNlpkipu1sCkKdjyYwwKv6lsW/VNyu
l88wr0hBPrWG/lStn9m65F2jgcJe0ls2LQAusmYsjjx0rPR0RM9LQ88bbyJ71wjB
Q10ZAVQtFpTdBaIPkEULS0sgTdX+YrRbYL7vlCiGQy54ObH+D+qwITurCdnSA5VZ
W4I6/UBlMboMu+cYuPgejkZDijPnF6wtAS7tPb/anaH21ww89dDUAPbjNC5wsl2D
6xgK2OP4fh2SB+35UqCsXqm77drKeXGLWOIJJb+PSEifIAyKHK/LaaNICsEl+fog
xrE3wRStoGPJfs1JFZCIqq9MstJ72vGWrly+L/A4oznd0Xgmtg0krozc9tb0cT+M
YUfBTkwg/Yg9VN9VOIt6yKnrkTAA/Tc/MJAxgeShkhNb8Mq32yyEmaxu08ub7/hH
udL8xGZ9Il4va74/wIegjdYJMez5ZGvZdheKv05//vNKgqebef+Z+1KiCepVEioy
EgS2tg9lFfAwpk/uPuuMjzHo9GwDmzQjOfpn8yYYsWCicBbUCdgKybR7xKLLBd5V
y0l+HNMorUqhOpp68gHnW85TZuTA94GPeNPDCf+KgYSpCG6Ezs6RNXj/QOMi9c5i
yp2K2+XQqAGoRnzS/MKg5Wz/5I0WME6xUKZj1+RoPwS7R9K5UBIBXgqg6TCBOnGq
GmiMIC9LFkn2of7UGYNhKJf7OjWnbMpRlWuy7mbvMjos8uVryKbcvEVERowL2jV/
kAw1Iqd3gUeuMTTf+wsNgsJfmCuZyGcoGJaB953+HBhIBeNja8HDrglhLb9+tqjP
VgJ11yK9J2H0sr/8JOofZMAib0yABUMVKMeWKIs8wh+QwrpFHOe8NTbAUWrYRdVx
tGzO/D0QSYUguV3CJyK4dERzn8CQnl4Kw19Zqa3XLTicQMAcMQ0+KMOS2MSzFuOK
PO0aempRZll+fqUdtD8xIQ8yCsbCh15Iss0dCdV+oa+DLYAIF3WtmEtNC/iiIwG+
D84PWbZOoHmc/pez1y9yEDFZPBFHvjzVpxhH5F9zSpWu/I2CPPl8rjDt0HSsQ8aR
y48A1O3HN7xUMdAAsT+LbpI7hNnjp2mCc8DGjER7Izlf5yZwo+ocHZi16dFVQ08K
GeYFNbFkhwoFZKhrIAVNAXdk7/HgK2ck/mXhDAn0pCSB13Y9G/+6LR5utJ4ZZ2KQ
qNWnig9DIWtTTzezbZc8hy8f9B+FghGqVXmbhb+ysW7GdaLf3u2sjshJIEAlNp44
WRuXldNM4IC8mSC471K02UUxEa8iMrmpnyID7tZs6dB5pMxcpbTaLZFCB4tynhII
LtEb3glB+lOiXMq5zAc7IJbs+Ead7AKOy5TYZRDCy1YtIS4RhWMxPqNXdobgOq7B
7Jt/aNm+6A5sxSU7VFFT5fK5iHCOFedeTC97V3+AhJikyGL3Z2IbjWil0Mu0bw51
gC630a1ve6enqsFzVlK0HfRkHA0LDPvdaiCOmogmjbaG7AfhAnbOTXJx7W2+hqMB
Zik8CqqrARqo7ojTtlZy051iDJO5P2k12YFRPRrJ5dbXfdaNPMD8HlsFnWqmOL51
BCmi0SpVSjTXoSJzUt0c42DNOEmT0fAaTnldkNMjLQzjAx7W6WWFgFJRkq5vlWOy
q/cxO79iJLw/p9RNV4stYpePFlkw9k5CUpOJ0WPUJkj+J9z8CtSrcRCp5kOKMDkx
STdfs2tnUz0j7VyQk2ab6ajebsWaRjCubYJGGn9u9jd2sak6yEPkVmbSUII5Ij8Z
STOcv8bVb5BWMotDnEB14PM9PSNLQ5u/cz8k/fDgDHSyf296zfNJkZBBXCKHUMeK
yHp3GcGkVn8XnuKH6pkMgbJ5j6RVAiesOf4D2spI8aF493y8E/L6F3A/l0lwRnrJ
hYT/uG9BUAMVV2s2A2BiHtMNLBwCM4q/Scn63059GzPHnPXG1yAB4bQwTadhG5oQ
KknuEYJVea6Yrai2YV5KGgI6cJqKkNEFxqLswVmhg1jXyWZnnEBJFp9abpTVF/2J
FXISJUyJeJnodskjKacu/pUq+fZIZTYhTo9J8Tyxx06ebxnWzLGeWlOetLXo+E6M
bi3/IXOZwiPCjWgYErKCA4rTVRQ6y+5A/SPzfdTl3UaG1xougFbwKQ0ABn3HG1J9
qjNXOdpEXGWFq5+a5cUWC59ZrSRpIBeMJ/NuMFD1RoKXtvHBvDj4Faj3IG+kYt3+
q/FYfOPG1nlcC07fwH+bFbyjAPd8S8ROKzxnNWrMfVtu1kdZ/Jf5EBSEs00p/RDM
Zr/3BSk/rE1IpuTRJvBULWk7MHiuQGw/AXkC2cheqr1XcOEjGYYQLwRoA7YE00kI
LQs64kFSESVBFyMUQ7K+E/QZvWTZ/qI/MaO4+kaooP8MzVz7St2RbCSGtSuhFU9t
If4C4XnuGjEujsSEQefmnQK8fmswVva1ldDcP0fFQ9kHsK0BSdRZbpy9ugupVlWh
W8iSCJzC+10pGyn6sJNRnJpgivGj7JJ1rpgzBndzfqZd1mY92HIaVwQrZjTeRlTU
WYT+1BFRGWC7ReUohfrnNVmmIq8/Ly5lhG9EblVAm0tNbKLfc4H2i8rjHMvRMMA0
b7yKYISV9GbBzHiNb36ILhWdERZ1zpvxXO+SsP+ECTqBm1DrkKFuiPICFLObA/IR
+szpLU21dH4Jhr+8NuzQSuFb2S6cO5fByUv1EwEjsQO5bGFXegoaQiFiKHf8nXVD
15tA5f/ZiqBKeUR32FntlZY5lcqN7BreNQMB5cMvVeZUlZkoOuy7zNLtdKFHdM1A
e9ykS7n8TIcZtebjq1cD0cB7eyAfCeYE9ovB9lCYJ99kKGdHFOafs5mDgCqTX3WW
cUFNyOcaEU2z9dOfMjplFg73uh9ISnsJESZIU5AuQTI0967kXMsUIibUpdLe6C+i
CrIyAHxMTn+FvJktnU8zmeUDdeFezDIe3zaEP6Enkc1GEAlcNS+jEmLVS3Se6P2E
rRcxj4VUOgyPhVHw/7i1MF5uIpcHfU7xC78S6I9QfYSy4zJxBbZkSwc6HXmhvDdK
z3yFv2AEEGS92fEHrliYQDIRFkFqpfWhvbutwAm/kUcYL8MhLhDVJJC3142S+1le
15GRxU4XffUWuPxyz79fiTOyb98+dEBh38SOxGDy60LC6yiLVAWEsiJ1h1MVf7El
2j89WRGmUtY7IAURIao0TFY6K/305uFVKvddui7UW4qPhtU0pnpcIy01/SMLy/4L
WJVQF+jmSdORrZdhDS6z7ZZocMRYOimeewMX04KPykycyMtHQRQU26XrPeRqt0y4
GGy8nQp2adYz6yKkqDhPpseqqvfWksKDr8O0x37XNCDIF0S5l4orzt8HLG1wxBdr
m38nuiIC1LhPtomeiwxHW8cP7G/luKaE7klzBPHF8aUkCpvzgvQ1lV/hHXojzwXo
EcJS79Rqi/3m+l3a9kp1mBliDjll9df6J+4lDJlC4pKG1UBdftZe+bTdIs5gG4C9
1Y+Oyk+J+VYrRRUjBYvwqsfiKbuMTNALWBpjdSPIyyaK4BgV/GOGag67h1h9theN
8RSGuc/7kPIu+e94HFvQ0PhJMrEeCKvEarP+Jnx40YpyftnPoQvByQ6/m0N/uWIx
DuUGgmWHGDTsuInKL8E88+pxgu5Kq2yB/cUuSK4KWOxHSopRTgsya3L/9d5jzud0
GafOGlXk0s8X0xbqntt+BemWqlYHWFA9KPYXaCmUW0iAfDOAn8VsngWYbbE/nGhU
g/njwQGH2X++IV7e1DyQT+xnq68ZY0B7qGinMpxtdBV1UiZSxzyeNi3xEgCxiAba
T2nWPOmnpo5es6hLbhAKWG4t/dG9OVAwX+EzfJYMvgYN3+VjgG4h+6XCpRaAQsgF
VbbyR46tlkF7TXBCvD+cP0wWnvLLHxsWAcoVIBqan8ihTqMj9KgYIDfcQjow2R+A
pRm9BvudvXFrHTgQaV+no1ISlkH0iYeKWoDgDRGfrrcjo2K+sUuuJWHaMzDl8EU9
TUOwAtgd9jcQsL6b3Hew6q5qRO085KQ1Et7H3i506AKoOmDv/E3B5XM1sPak2fVg
Y1R20e8Ig13aG+Xt4OFnZ/iZjo2LtBeXErVIaMqaBQMAK2vffesA8Y+kiF3YjSHA
xlMaxOEfDX1uTOcJ4r7SIAaRv1FHELP9IBvT6V9993ncDhRSyAMpTJG+uIWUCYVn
YUws7dlQzyfjHYWaUU/THfsi318Rnz8n4xDbhaQ1VCuS8ircK9bhfSqgZOpYqfuF
rxuGHbg2CB7Odgg3JNu0AdQYYodp10SWqKzTdTzJBazCUAmD6EvS28w1CMrBkwJR
C37b2kIRIcsjfvst4Xf2HD4NnLOt33zOOfkodWtAg2IG3ByK8j//Z06gZ/I5sVqs
Yt0iwqojlof0tXKna/mO7rQD1ADWusK4aU06AOUpU3vmBTtOLfbuTPgRB9XUZGrW
UC7AcEX4qL9s4iVfFDwees5nOrMqDVeKTTG3X8w+T4KDw9KRdrlG472HuhnbtJdI
B7lYhWnXMq9DKNoEoGU4nqEXI/LJ4h6ltmEOiEN1hnwmmWuBfLYnstu+2GYGYICv
g5+4bbuJmt9pPvxsTi72Ai8fJ3BRgBtdu/cXxRm2hrm587VN0FScbalviic2J5vb
xQ1dymtELuoTQQdzLFu0isoYEH6wQ0EAynZWuSC8NgEE+e39YULgOgpay8geO1Uj
KY7a1rwAk1offMKQABcurtKngG9z+1FMqjm4x6gs/bvwUX+AWxDBbl8YN+udKtU6
ouYhCExQ/WP6qFANr7Xsyd1TvT5TUkn3rd0gKKXZhdr1EBXLLZQ1P/i5LIw8WDjN
37gOvJBOnn/0qsqlSy7/qLNuafI+L8XOpwtxddssAQfTTIKMflJhyxrvZKQPEpmJ
z8Xs0uKJVfjCEYM4JskOAsf8dfFqo/t8MU6uvhnqNDY365NQjuSzHKDgAlXhfI2w
ZWQtgRwzgj/4Hyhaz82k9yL1G3rHPBtjb4ZgIQG+0nyASXwewQqxtU/TjGqtk3Oo
oKpyhDqdTi1hV5Tb4Bdn48gmQRnLQaQREfYXzvAxtWxKR+5e/ZxtQrwc7kFGaOOa
3KsbgY+nFruuRV0Jc+kh4Ri3HqDEmea49eyfjx1R12cxIFXATxc6snnVjImI5sOZ
Yo9JEnSHBMQjYvbtDVieeREtVAWTKGOzPi7SlWfvXiWGzd3RK//DTgF6aevknH1+
q6h+5xGq7JefL0JPagWZHYyia5oEMVfmx6aYjRq9mmzr/SsZYV1c8ZyOjBPYVUee
qXiyRgpK2vHWAA/OC2G5UQ8QUUIbQvxLBP3ywp1yiTwNzULWu/kh9/FmPwE7Oi5z
7+zCLonxs93X8iOqWEXgCmN7Xm0u9zUIJJ77eZQadGiaOqkkOtS6fXmTHHqSB96w
Z6kfYWqz3kKZ0cPR8O/v9I+kdpQ8epy/wmkRA6VMVeE4Zy5wMK2piTyVWQJV/sLC
QcyE9Z03JrG/3Y9W5Li9YRs5e/3DqUKRqRQg1r2FrvQaMx6L7JWs9IBAysK18LEz
tEt0wPeWntRkWPn6XTE+ZrYIjzyHoMTcdB1VJOrXAXuM7054ehrNxMrh9UmBqtBr
5Y2vpb24ZQ0/FyVEcUpQFN/Cizrq6mbzQwhxqmIITgd34/WdfmWk2q4ggl1wYYCc
Qh+qQo7dY79BK2Va3zl777Gs4gFKrNQ1uXTyd9WGB1W0R1ahIBbYM65TSO4+dEFE
I/gAwtGIl45vRkdR8mOov3mYEFfazu4klW36XEBdt1IjaJlRSk/LE7tyxTulcu8v
Vbw+fxOiMwwNBjYMpleYyk0XYCI2pYHXj247F+Q/WTnkPAmPcFZtuJgixWwPZibQ
rB9TY0UaCXPoTFptzduMjutd47i5bGqH68FhJwgWk4r6bM+iwNC2G9tqJYf/Pap5
rTffIpEx+CG3uW1UTrqPgT0XNB+/ZO+xRi6spkS3Wq1MO4c84ACycGMlVi4wK8hI
X+oBwC+rRXZNyL4N/242YzU7NlLGvRN6mIxDEXf/BEqixqVswOh/RNl5WQbbhVIF
E2rDY0blFTKulUuoDZtBZoMO6NvGo+hnWVmb+D06RWTR85VaZ0NG9VfeBlok6IjB
oSuFQUHD4Fz+ZdElBIbRMHa1EuhhAvPOoWj8wLWCxO3XSt2Z5sDdX6p44RE/84x5
JZUS1V9ghvkTJUHqVRz1PD+wt9C0d9sxYsV6xcj+xodEh+3VOPprXvPuNJSABEEU
E9F6vZi6saH3AKL1dLrgqdUtT4uswVkgzglSvZE52ObepCtrN1/bB3CUvMqmv6Cf
Id4dqOrZmn9EtPRIzXjpy8bNiiK379aPgU82sLQ4khdnDZy+qqYF0BSoFa3CYHmV
HO+kN1cSzTvFOJQC6GItbSyy+0pcNiJ8pqqIfVSTh37FqoNMTyncfXitNlqzHOYt
1CD0sbcvgocdD8Gb6fMulUwBTUfD1XUWolp/VkYgW/9DKQTT4uwZLQNiee4IoSd7
AX6v33UULU0m8e9HNiySM7YKpMJIhiU0Xh7AjMI09TvhKwzYj8ft1ZfiMcWNfMK1
Qlxfe/gEq/KkpNUvxwHnXbd4jh0zroC23Uwpi1vF1rciTneUNXfbe4l2XuB4jAhh
ZiDEo/SEvFQqEK+ihZPuPg4rFr3gcEDOuGy2n/gdlVrjswXando10pGg8Hwmo36f
3PJ6XQxyi3fbd7jNNj6KzbwjtgAuiLdg8RhnDRY4OycnHjCzscBPOqAyk+3Jb5rD
YaicBtViKWvTALXU0er9EvQ41KCTfFlQ2gcXjOTBnJxla8mcigTTA74ZDHR7b17J
pa/bOTh5+UpeM8M5IpyVTsp6z8DSmEXadFjSrf+QeLvM0n5K4PP+UPP+D7jZsrW1
vI2x190M5kDaA+fwJE8kkNJLicFnkZdQcqlf+gIuO4rqMJqLCGl2E3MQLXO4UmDp
8IgGtcz3qL3FVLKyuMaObFqr31oEh7gwTblkLPWhzsvoQzMo2SGJrubm2FFw5C0W
FAVWOD9qs9A8w1nE/0yqxOx9EG/iB64OY00MhtqCh/dkBscinzhRqaIuB6eFJe0e
Yq1sOVbFiyNPyG5NEiGA67AhbJFIPCCNL2botIVkQLVL87J1E4Z9dAwYa+GUNYOr
A74NZi57IN1pByjonDwmsYPAO8LhEg925ZXrQ/HDgrCJClbXWzfuYnoadHlMKUck
hefVLKZ9X9hdMQo7DrYnUa04sc3WxWyoGKh7rI1guHplzbOawKoYsaasS7APtQj3
d+Cg6y05BIjD8UAabEcVfNXtd+Bxptqwbxd9p4xyOYBKqariyknTMmW+pHS96mP7
CxVY6Ue2tQ7NG3HNhhsE2UXzFnpggYUWWzaYb70Mf3hIt2crSAPjtnJKnPrbG95A
xTuW1vCkSn+TkBXYUvy3vjI7ox1PblyAp4k9TbTfN5omudK+HZFAp3P1d7r1s+Yd
1+/I+FaclgPp9kI9aoZQUV1d70INQcAVor1kg5o3yrSWXEdlYwPXhVvz+G97Fmjx
Zajty072OhBFlbRzPhusmE5RAHbk2dWvRnCw7r/oiRhKdYFinVg84+WDf0C5uPwP
+WBeqCt7UE8n2gT9yGnuyUV+wdzzn7CcvSKuiCXOEvIsgpIcJJ3PTRvMF0wz++SD
31W6YJ0E+burZ9pIFT9kNvIAp1Fghil0joXtnWUuYtDK2a2GMPdtooSvmCFm+r7E
TJKMuvyzbwVxH5T6+fA37mK8Mu+1eNP3rs+wvIo1KCU7G0lktt5uK4Lu46palzi8
7rUNmqEwvUXL6eKnB4HpHOPmLkGLVs6fWxzureEGTDId2nSrUdNNZmd20aWNx2g6
C7fKUsN/krr02bfqsRRUx/GDctfpc3HaUy/TMkpY4i6DYNoXmJbLvPcKiaDE3exr
n7I0VxWKo8dXvgORB4O+C7Qv8Bxu1dRmNoaDbVKHyD8nObW4u1sCKpd230B6NZZR
lAtMsaPn4K+wQ5Jt36Vf9NJLa/ut6l+Gnt62zzCA/mZth/gyALCqzVblwN8JulgY
53iYjOfRFiha0FEIFW9SrZ3l5HhWKUNnroOYBoFQCxL5+YlgPHbFffkcHXQ7TGSU
ZkXueNNXg8HAOizmax8/1LUMQGiKrnBEbpZPoHM/54BBxvJG7jWdJ4+Fp1lP8+dD
aTjyUCXMXGPC/Cj1GNKYa6/BzORh20DHI1Ej8QSJape+kdJpXZ2QG0OK7Ho4x3TB
6LiVnuwXZ1TfBafXkawx7HAJHxBaOMbc4M/2cWn2xMGDTnkrGjFKOBy/r66xIlu0
GzG+DbldLZuA+MQUZNG+vJEQULsxKb56tOemfxUHRYH21S7zGO8QoknPC6qodKdY
C0OYQUaX8i6y1U8IxGnj+3ZpuhxD9u1MuEftSwvitL9476zVWyoPysGH+5mnrPLl
67MYB8h8mfPVWB9Jzf3OEgumdH44tJA00pm6OuKwj3tv2DOnRBLLzLMWfxiA1bl1
tnyhkhga3mNP05fI/SIJSGeTScWbR4VRBnXEqqqiJRKap2NtY/0rzV42S6+b24Zf
HN2HeBKymUHqIMHpd3C5nRNfW6lDCczWa3Zj+0FwbW5NcMoW4CowEqTcCLsNNzEX
9HK5ZHHEXBNLq3GAcQKk34DiBy34DzXftoUhZuC4eaa9atts985/A3GvARTkeGXy
BiWx3YKBTfnm3g5GV0K8d6xHByp6504O0nru+rrMbQHFznCZyFhgPIDoL/9szftE
+m266dXCPCMJVoilbl0b6x0BbUzTMzGlnzV4PbLrXrzpaKwMwXFDchXp4tR3VA+6
EWyLMSNyu8inwbgJbfIJgQO424y0LpUe6TV7clwMGWlSfyQ/aK3El19j2uUoUPsd
c+PAT5MsSlDvgzqqifFC8E4tXv2jKrgo3BUapI0vISLSEmXnRkokwMzvGejq4hO/
nWSA+/kmkQ8GIxuJljbJ94iUfEyjmZB6Y56irUnK4s9TG/YP1rzEHqqJ+N15mlto
yADRSvmQts/Z+UJ8HqNaJbUGB0EUvi7PmtAqSb65zSTnFslzisgK1TECHpKqRdx4
7RYfteMckTfzuh7deM6DOQtDI062RtW2LUzk+1nkXAqk2sONd1yf4xyaqHNhsrBc
SXEgtGQ/5lipHA1Y3hVF/Kjn9L410M3R7olCTVVcYKYem5k+y6q5MOloJp9GpAKd
1qufZ3bjBFox9vsVaH9UUBykCMS2EI/Px0/dqThWyaIYHJA9E3g9iK0AeD1eYBLs
cC9py7hy+72RBkavtZp0ZKUyjNRs1UpOmUsnkPnJVsO1TOYGTvXiMe2jCzzNZRJ8
SP8EVZUSpeX/md+1NnKPOeQ/da/DZrGt2VxDWIFAjngSwMXH4Ij+ff2xA54ShNWr
pVbZ8Oi2CqUkOGm1IH8BEYdjH6AyTP4xtd83CVemHl7GKMFPZ7rMl8Cw4SZ0A3/a
Cssd6XY7w7tU2DDwPebflmHifnnzacQm02xb/FM5odTDDxybIItWdChc29A8HyVF
uEwcFdBe3cSeGiRiVknm5xyzhmDmLOGbF/gDRbbuatGLh7K1UFhdF5qO06gAOwKW
9g1dqaw38ksM+M4aO1AHICNHxLJ3uPBol9xkfnvblhi7OypyTRqg8YEbnlipvvQZ
BwCcKu/3bFDMldUS2gxGOnQ3UGrDNQ4ULwB15bGlT4uj4/7/r3b20jzlSR/Klsyx
R5udcfZm1mwg5KQRZHj2VosOJlbjdHwLZcFSgB2DK8uaRCdppbEMUg9IdV3HTv6i
p9nTTdwDrKHZG2vTnXZ5KYvCiUC1QCdtLNLyXJKut/wSuYjS0Wg+VqXyoKl7Wttq
7TS8YVUcl8xjWcE6eH1J1zZfz8sPapuUh82t/fR9GqndoSZJfBqxeLM+bso/uh9f
Rz3TAyhcmNKxDu+wIk0dsQP7T/1xbpiX9rnT1Tkkh+bS77+kFKqmmfpijO2xZ+5h
u9MLbGa2aQvWrXmWITh1AA9W1Sd+3cCtRBvjuxZgHV3mxFVyoIuiVOR9km+hIki+
UUZ4H1RUVRgoR+PCzP74hVuPNoWiH2NvphBKM1/7HvErmv4V7CzGoq46lvLkv8QW
eThHqvevabkoC35heM4PwYd7sakrNKtDEUkpdkGuC271NsZl9NIT3MyjC/WSwWsV
PX0l9gijT3s/8erf86L54HLO744ClYysyOpLDhCLOHuwwruIAPsuOW6SRk/Y6LeY
inQXpmfj7vdUpq6O+NyowkhsNpfnDaCrJLX8QqNHETtfxCyDsJK5OY/jDY0o1Rac
F3wBoKPSsn4pbFk4Dz3FQCrsjbgAtfyu7yO3XFxVDDdGUfpoUYNmupvazktc0OmR
XZkiwzCyCtEOEtbyhZdkJLBgHssvAjbw/TF4VoDUkqN+0GWJUjd/N2VZgXlpc6On
5RlhvBLdRzbmNnT6Vj1Hr2J9ag1RE24ifW8sKAaUyxWAjiObgMsf0x4aRl8HD5AU
4PuoBR2tga4wwx1PLUGSjbVdxsgrRqM9zEwL5EaKEQDpd8O/7r7xzS6qUdmPNdOQ
cU4/TTCjtKWAZ4dkpbXq+LLQezMUhym4fk9XuPTkGO87516D3Qac8kk9jPoUqkcU
/QQdxeR47Zu9Hqmypz6KhZRUQGHDjLT4Qo+oG3m9sw19mqrPD6hZP6S4ZSQDkgxb
lSPLB1Y9BY5MZkZnoK4F64eHIiZN9Fev7SSGjZHRu4C2/ObogQ6zU28wjHzRYDsQ
ldEpaSqsp4u76pwwCUy9IvMt6inpLiOCmdYRm5/cBTs3CcQYq+hKYGPT+PnDYoiU
Rj12Cj2Mbui7CuumeMd4Y+9R+LnHyFuz9CFIVQkXCfeKfszNq3jmtU8jlDOdhnKN
5yqscItk+1N8IHzG1pe7ON8NKIlXXf5OcZd6E+ANmae+zBmlCbf392o9IZ2r3R/i
aQFVOApa0TqLOVef3/OVJFrq+BtkBbbsZGQHlNJPOccd4IrJsLec6B2z9tDv6H5q
LSNydt6mJ5vrXf0JQrY/2wGykaHNjPZbQ1C5TSD15lGbvK5wfrOXMs5DFvwOYW+X
CVypbZHmHrgBK9YRhKfEUBILnBDDxX8ZEpmabDiPIbGgIIf5bcWFrFP1zC5TaUyf
bMWBFnrcj+urJ+2tnguL27s3Ujg2wx9kN6GGAri2/ACzO/sreZGwKS4gzRUIabIr
kzLFTuleyhjZMX+2U48foc5E8KuW7nE+SYpZmu9p8Ear3Zibpw2F1SXyePI9y+A0
u29phHOqtHHGe0x2URHqLGijjecpioLM3I0pUOowmn2HWIDGNU2xSET2GXaENVFp
dVKfzlRqMIWIJznQgthW9vBN9FoN3cw58bwW48J2H73t/86SwN8JZzEchJL/fKJH
i1nZ0pCqVzQ/AsY2MH53BUzM+tdqLI4wwV3RdJ5DAsTkzM8YYt1xis3qTp4XW87q
QeVtU6I2zEYFH4Gw4Te1B0WjLExEBbpVTub3BHD7T68yNZgnM+ozLoaOi8n8y7BR
wxzhm/eWWrzcC+qYy43uulZYH3pArxGUnpZROP8NkDZ0kHhYc3NRJ80ntn+gduEg
ZW/uqwXy1R2Qx6jvpFC8izkNfWnDahHXZL/5ijXdXzsYL2iYCB4sb1GxvQYpJYFB
TyZP++H4YvksqvFIfum9zBd+aM5nREgLFoT1KmT2/sPU3hquNoQarDyHcUA8g6vp
naHLrJ49Kjj/f4SYzq1kFq34kU8psZ2Xf7wHlTP0nhb5el5je54aMNly4P/puiJl
Nxd1e4c9ak03WnNmi9Gubvbdbu+m4Qae71h75v2wWhFWzQ3XQfScaWUr5Fqow6Tc
o932QDSP05JcMs+FUXRQBOBCg94RwjesLuqW2m8/h/2VYOc3CJmwiWPgV5Y0PeLL
aQ6nJWrfdXOr04PytlOJWCm/rsRZMpSRbryWXGBt0U5gF6on/w5wXDU9nBXgMFvh
joLq4vV9mNWAxMkq7JO+qwgo2pkq0Q7TpcXtoQffDju+U6ySBY1QnkOK3fvjxgCa
GItc4/dJOGIwNel6U0zGEXq6XB9/1uvmVwHUz3NNQBQ5X3t8ReVgKH5n9Af4KY3D
nTOIFt4Kt8kqeypoBM+MITQfyamUdqndCp9rmYBjaIUZ1YwhKmPR5m1J267NqH1b
K3o+aCUozETnFMJfJrclEelcllFEVefCw9IlrmQvAmsiNotmiMRfaD5Wqj1dlw6z
epJRvb6y6ZHGC8gdjOf6dNOhD7eHSuq6Bb/km9ru3W5SLzEI822VlA4Hu9Xb+ymj
XLDhx655N6lYGDZTuxMdqrAAqsba299nkCA4nRLNPiuN5oxzLu5XQqjzEXiSPvox
gnMERbOYzVITTbC0FkZAB1+w4owQdSw55/pKgKzLt8KxuPJOXP/LieRX38Pzc0vC
719sreE2uvWE/kvR6qHvmnsLCc3RVcp+peo4nznjizdHpUf6shN2skszguSdnWHZ
d/BrodUyNrORK6jmb3K5HOmWkXfMkIBRCXJud+dOEdUVCPdLX/dm8/sB/65zWTMB
9VR9jnWO2a8VuA3R3BzCZ4EcxHwGKbtENePIHhvQScRHE6BFNyqzBZCg2HX3RyhZ
juyCcTvxZKoqa2BUvhbF9o0xWZ32cXGESy51NSWKuklVe0ae986KTPmgFGDztO/B
bomM2zCddcwTTXElu9DhZGYvEwCoY1/hl4WVDTeIdOQZMG1jVPbBJW1xGlJ6RfrE
lXC86cjqAWGgYq046P0lMy7psJ/tqpmcMwB1pNAKa91DmmTrh0hWX0ouFJHpDznj
R8ZOy1wOeMHzABA76k65qzCgUVtlJ/NSGtxXClFxRJ64dLEPBK55t6fIEk3yWROt
vIZb/4DeY6EEInjYukGZ6SfFekhX2jSrJ58h4tn1ZNSbxHFHk3tQMGL2gbHw3dPR
LFkUmw8ZPtZ/IBFKZn4k2ZPMrqSQ1KhDxf1MDwYU2qk+VUpWA95mirAgfNTAuJKC
epstrzgpf1/WYWX45JPw4Uj5laGp3cA1cvzEOzfqLW69HsWCuymVyy/YmKkRB6eQ
kyN3+swFXlnOKRoXPzbHOvX9HN1+Ldimy07mEjiaAtSywZhZGgPAR/D6ziW0yxxe
PBf/rHzr7RqbtuB2enJTeRXt1oPAQmLMCesyc9/jYtMUecbqieRP7gCrWPnDc1c1
ITUBo1IhFTiZAVzMWkWEc4lbKcO5Pf+BEd88p/I9OsGGpjF12ERPJ4GldvecJmsT
oFjShHeQCBYQJ4+CdQ/+EDDedWINaAnL71+JDFOm7i/q9tnSHJu0OBgRMtXNC7qw
OS9eOgdQirNG2Mvm6bMObEA1NzpQoy5DIXD4lzdKMS3nkewt9ARYjfz9pQKnB9ce
I56A1oJuHJec3OmSHqwSeMlGFm9UeB0cPX/WWFTDx+b+e2tlM1a/P+Dqsg8m5O44
PRyae3+teViEO+TOB0MxvTp4X/qCx1dtX9Oir6wr9utvB2r4hbdfvTkwlNE7YPRg
UR8ZztjLngWtDDgk1ErSlILOCFhRPTBIXYBGPhkuuoNNRhw6NZU2gQ3UjXn8nxrt
FtqUxq5Ls0BhZFqwMMtBsOq+N4AJ0FeZyrBuKNNnSjPMsSuOstW1YlbToijms25+
29WPhwdmzs509J+Oc6vvWzwtwSQzJykMcxNrv7yL67bSmwX450O+HqSnYYhYSFg5
DvZDAXgk70p4RqgacwEYaowerjgmqzqkCbC2uyFMMLpHB/kiSeIUBhBGDOMvPpkO
xes+MlPUwR5yXxyIrOVnocKvGbz/x+sxRyp9/m2aFFgC1FlPLnp3eXl5IKbmioJM
DFreg71Y6dIIDeTOrezSI1UdJH6X/JbgF3ysfJArz6iBLZdK4dV5V7vg5jPKtTLe
6PKsSb1qozIZJEkFQm2UP8sazOn9YnRGC6hIk4CCyr8rhzJ7VYy7AzXYyNpVZw9t
QluXsECuEFLzzs32hwuwhsZ2DCLu6q6IgeibEQ0Df7c19AsBoG7vMh4YVgyvvS6z
ymC66Au0k/vv0o8HMegF4C86l/jJ38HpiOBTACzBCj/o9as3DsAn/B8gtf6txPMX
HF3mkOd2O4T4exAzOodi6GkWx7i2RBUpeqjewHL/5Wv9bztrn/MNOZqeWnPoHmxf
4rNhXIt/zcaaZ3AUuM9/c7AxDulMXnFIg7W591CfibUhuu13qpwehX7SX3feWmWo
QcV6oQX1bqy6eDXzlPzJoPqvV9zVR2YwMEMxJnClyaLpC4l6gUbjT812lq2iU+tH
nx63d7fYTeO5VXqiEdJqZBEdaOFJbK2mj2N8FxymeIflzCI95LrH8qeIPR4rcfuW
9TtqeBiyAZqAURV0cV5CfTR6SRsGJ+mgi4Jc4tYjSTEJPYYEqkg6Je5uVao+yZrT
95KvZ0qyMtWViOS/flpgGjfo3uZcYKjD6ILk/DvmoE+mqhXZTE5TXeADw1p5Te3b
WE26uQ4wgPUGC3g4BY4BAxz1BB0zYwWrQjpO4Dg2CgjwKKVvuWlY4EjHUMlYruqf
ZBfSzUovPWZH55ZO+BwTtZxVCcrpvSSYiqKzNb46vzpqsdyyD8hfYmghiDS2EGuD
g9DFOpIkH2QPWg8MA0dLBmXVLVOnmuYE2+8TpCpySeDVGyylY1ql4nPJkhtyKpI4
0xv4GqKNr1N/2Fzfd+3cW+CcpFu/6aT9uUty0uEPQatwYengq9lq/XURO7nGzF6M
6aBSJBSARFVSAub87Wqm22Hf36KG8nnbL2UybaNGMH4QiKtj9BmDIxbTYUiACXXX
7zk/rFnRSW16gP5RqrOvYpvtBb52XXF4puRae+jGOaSHT8LppxeCkd3v0pHl2dhx
9PSciPzC2wD1iUygvai0Wex1YrXddgUQCFlFI0DW/QNac4ae4/RTMCdtiR7ejqft
9Xwg2ZvgbTvFl7aGh8dX9tkf02ZR4j5HJcR554HbubkWPYaZDoCUXLjnqImjR64u
Odf4kImiq8JXKKZyUHQnUq+8jy2P8Y8fK8Hcykn6aN4wlgjuwqjhejdlXG6XTg0G
PAcLtpVVSeYiRDJ7Givn+kjOnVf8wNcTDMCaxLHdtNs6NyIVaJLGkFOUWXcj8k4n
xBO3pbbbp/GP3slZrJb+buiiSD5ZQudLG3IIwnQYE9gVpDDKyqqCjmkR2GMn5gFu
IOyrrdERcXtGEhIhz/1RyCOlUcNncGP8cNYFqdrgg6HN19fFDCWXxh5XhV9k8AsZ
UGQLt0MIGYVLYj0PCCjcuqy5QzmktJLEolCaAa4fp0g+eLtWE/ab94udeDWhHBpb
s+qbr+LJ9MlzPoBzPZH+Rl0rDI+BMUHufJAksuO7u824IFfRS1LflVfs1axTrGHz
XSYdkQP3cZty9DL6ZSBa79eQw6GRQjWd9VxBRKEhqzBa5owR22t8T0hr35uVq4Ry
YnuYXh7CzRvUq3pIeZBdHXiSmccBow1mLjbjkfrB3bVWjm5/sxVOfmckkO8ofm6k
wPmpG6G7LEHXPDyc8w+qxV9Lf+f4VQ6rYbF5FqQ5HPQESTaLuP9ntxsw12A6pf4m
yWkLpPjd/462kPW8xFTEgUPU6cyv809jEGtrNFrVDg/G4yyP18LfJJCvMBdVT3F0
fZg6H1WaFTguiSIPJhkbSGVHMz8ViZdNc80X7Ow5ygtikkPEZD15N0IH8JzjD7KI
BJhOm4pbqX+DJBfA3aa21r4PyQ/KXuIbJY6wtwR4LFz4g9Nne9+BHUjbUSBcDZJb
0cONGA+xcgwUwsXJ5CAVy5DL57+g1dEAx4qoK0xaynE1NxfXI7n1xWCrw5wIgEwp
3WLuUIy7W0vnRCViDqpsflTIPFHP3yekkwYbYdUQK4vZvVZdJe7PI2Nhrz1vRWep
Vy50+/sloOSsa3hdvmWsyponP4N2IUe9mkVSEVFBQyRSS2iLBIqu+g/NWSto8flq
9JxENF6hibSszYZ6rrH/habOCjx8vZvggCbj+H44elFDoc1EexEt4WcoRcKim5dm
fhZPeaAPR5R7EFRKauMbRVGSryhUo1zTjTNdn11TKIEW3DWbrZY6Q2i5oHY/djxg
LyJMUj8MiJrar8vyDXHS8pnMPSVXvPrXZGmVN2mymjtvgMlqUiRPI0knqsYJQlkT
3CyRR7LpCeICM6FsV/Fowo0BLaHLVBX1OHLFqg+EcdjQkpggg8sHEAGJA8irq89w
vIduif4vWieWC0SIq7ap3v95v1xmFUAqEHz4JyebhX+J5IlUHNeHuN9gVTd0mn7V
e+8tz3OxWGjqoDmNuurzVKa2Y8AyqVSvSrr54Ug+wpFPjE0b9DlUSPUDyjafU+wu
Gfz1zO0muytzF7beyp9k4lHcNvjiN4Nt1WMp2KIcwLEBIZVulQV5YANR/4ObxQG5
zzM0etp+njc9aXqAXFDtFdMvmXcvXOP0wQ/gSiztlI3DJZQR4vN9u60EMNEHLDvj
FwW8KWnl4GWSkJRrtJ5vvBMVri+LPZRtLWDxZpinsPH+UvxUYcBys1Ojn4LcB1rd
6xIMlpTByuLEpnzpv3JAC+xRkQSbD488JGuqZMxlKqvaFVVCE7TjJCE0YEoDbWxf
fqBXmjclFspzc3lTvCVNtifmbh007tSSPeXG6xPmjISSVK33WKhQ5GolnOTO8sGX
G7UTvZuK7YClzH/yxVz57hazx6EcCXN0MkfT20GsfXTXD0yWTVH12fK6w5vaaH4B
jQxyD5/GtUw/7nIPRL2UhRPVeBugjlrXSqNOH7NTprFwlS1T3ZtBToL57v7N0oAv
2ILv5M6qIEbri3e+5pa3Q9oFjbwsux8t/2i2+DFvgsp0UXsHNEDyHc0tl3veMLUh
j//cXkMC3ABB27MCNgKnX+Pq3RzauyesbGEUlbjj54Aa0FAf8My2MaOM+UL5r79p
bSS5CJqWr7MbPJX7Hv4ebq9t0Vci+/qLXMoh+eQrLt8Us1BGAk0z+ECrEISazQc9
EQ8jr2u1BaVF+Af8w8/AfNwFtocnSXQZg3LhurGj6mIji2GcVqpi31rK9gsPwcUC
sElYurPKT1QzT930jj2nB1uV8+VUEWhBtjjMtgWO/pNKTBvVgq4uaIBTeJa4ux6o
jMB6UOmZGektDFqCVdFBCN11+9SjsgJcoRx0AxGPenZuEuy3EgpbzwJN1DTzm3T7
8q9qH0XUtLF2h9hstA/vb5f9bXx0O80BGdtFGntR+4JGJoNh7SgaIkjlq8VJbz7T
GmdpjjwhyFJJFYKcbljPYg9lvAsTTbk5LxdRYPt+01uJGLWPblOoCXd4z1+cx83s
E6HmrBPvwa+31ybu/9M7yG4P2jKyNk9yst750jAazD7Jna8Z7/UM8opEWdoduzDJ
LgWKOs7AkNB7aNxUzaBRamj9W1tOriYBss9CKtVuKj1xwSocabRMeio8hpjHWd6n
lmQEbBwS+0tFqBtwCO+kLIVf96dnvn4VPhs/GAoKHosQvzTud6823HgkpTSWQ06W
OrbLjwIKnqdKQhSuk5IN/wjhfbPxc8bSMH80Mrv+K01q6LSVsJMUYhjHbTwF9DnE
96GBJDRtGAf3sjSscm+JrozJ8ru2gTYi3y/bwnBSzosTF3VX0HuLzDSO0qhCRZQb
/2mDIEC0iJrHwkHk8HMKxvkW66wYw7dHZky3z/f0wXB4MraySoCIPEusK/ZdAH+2
8r7FVYm0w4pt2Hz/JhwChEQrr4384fNll84a0xSiaTa+XDsOtrWMLnreuBUgd1AT
lXkM6sqi4JM9b7zYsBMDDTcP4E41WwRUBLevXnFrV/b1FN+AZvbBxNnSsZLdQOoX
dz+qcUh7N0Uv4CUyxv2abEWs3qYzBzDKe7nvBpAWwNI702pDw3OJrPEaz+0ZZtOl
4G4FugXZ9JCO/FrTf80Y3cpNTDwH02+0YYIPiSZjUyv6mEHRxbX+g6skGa4rBAH5
XXNj07f4ByIbukpeIokmdT/wwM4pZZXjXVxviFJmDVtS/+SCsR87dl6miYGlx5xn
6i6F6X16D5U78jxBe59ZvJtTXUP+5Fv6g2SN2L5e/l5LI179l/nho8UB5C6mSIEa
7NVUBYwZpBL35FRLSQR/DFuxXNGw55QYxIDd8g2UFLuoP01xb0lx04Lyu3rSHXe8
15H/X7xBikdPbIwhmhuP8OkNryzGlZwEcaxlXmZ82QIOKuRXWJQATkGJygJ7TxIN
Ik+1ZrAO8SR2br60g7ekhjcgNOzZ85MRHXrjV2XncDWX6d6jDo7hAgbqCz2zqyZV
UEGCZrICEtzXwRWJmx+2Ojq9w30QnCoHDsbFNtqg+IcQejw3dHjelGP6kN4LEyky
ibQvxk8dBO8NH/8rggxBO6m7WNO5t04WzOK5NghxtqKr0IUpXwRVz5OEGN54z9dz
q1sC8AxNlISCa0QM2AIcBMSoPb+NPm+ZXuixi6GltWDf6tu91Y0LMC4BPWuoMs0h
5b9CMRE46YETUi3TMR5Y9H+/oyxonp2mEESjo2sarANFpkzIqRYPN6evLCuMhYY1
+vx4rdyrZCkxnRbWF+vWFWx9Hb+cOkTk8SO95S31tZnvHXHRiSNFaynWCmIWEwhr
4gqnmLKERGD4LhR1glz7GjlKN4BpwdEl4j6iOCwpr9XivUl/hNKdZKsaJwUIsF7w
P9uiZMUjuD0CYLl4QQAV4xsQCrNloNDG6QGX7yY8igVDKtFIcHpR2/ZRx3VjHRL/
VN2tstC3dG8yusBOdd1b+ud1KOzgqqXM26aXOdpSWtgB1kzRwSA+dcIqgmqo0knn
9utpqHtUJ20A1LNgFvOZoIysxqe4O/5laIfCPcW2m4kIbP/mofZeL2ay4B2lpA3Y
1SlFoSggmavTC66Q9edg2gGs0YD5iDx1nMIFld4kDHSVJFxNmi4HEL3aC/49VP3V
JTXynvDjmLGettPW/tB/nA6HBbhQW3wULeC0K3TOQBLD9fEIAhq9bAOg6641uC5j
mY6O4o+QNSRaVKP/MU+kD5XD2EzFLyypwJpdLET2JQb2kdZKOFTGYpi/09oFmGPw
NXCyh76iAbIanKCnjFZrbTQAkbqmhD8F/paB6WfUGsxEFEQEBIdIiEyyVNJ0AUB5
ANZsLpZjnnxLFzzP3QSJGV+tpZge1xHauzZYFWAm8922KzHm5e2f+otY+p3WxOkE
uoiLAhDY7sisW+TpZ+5QVBPu/rpAHbVgohpqpg6bwxcY29Y+DXnxKSGW2sCxN1Eg
0RX3Qv5oXyoXoMD82lJezzTCgUpAY7pczJQqQK9Uwh+rQ6vfSzAf58GvQKs4BFtQ
ASQDhmz0KDDqYeKicKZNokIZjxNtG+hMOQ9ytNKcoobT7QsAPY8BXB7vJ4c4FUsk
g+qvY2m6ogCQEwpzvpjzlwOATue2yva6WQLOKMc/LYt7XE4oqdo4oQd8Pkuu5q8t
flQ3WrMebrB/SYmDft5n9Qpk7JOAMh9nZOBgFcHeK+/Vf+EkGKKK4jxGhS0r9JaM
5BPxiQEJDXh9EHbleXKiwP1yqmsMNqn0GbnRW9ZZQsDqigE305TDUn3rvpMc5gQn
98DG9vLBrL/P0tSw/8tM85r8aa8Wklp+vpZ7ECpSB/HPemNeEF4M/v46zfnAEm9P
ykjqZ4/zWit1s2lfNlVWtXBqlo1jcqnvLsJkSpkoWq0gujjUHgRQDmXIITtTktqa
cKeH7wBs7Q6dENPOrmJ9ai+9vx+4Nz2r8FkPOoMAvsob5b/lZlONiCddLezQrF3j
DWpVRgUy48D4IXf5SZyEFJ8vTiICsygQadcqkclz9Xzjdje9F2aSHEZtMez34xj/
FWmx0puz6cJFt+sjTsXjEEV9HAESAr/nk1yQ7/ib/kFNTt1Xh0YE5sKopz825zL8
q+hFf8jidNd1ZsAYVcqaJXFCoBlKJ3GsFqzcCpMb+uKkXqFHr2XDe6RHaarAZQ8B
JgIZ6suYZOuy6lCumnhle4jT4kRybpYk7snGo4Dk5SFeM1ldnWsi7GQ/XkP5rSm2
FOixaaS5L8wM0iXKsgDAMi/MF+jEE4m0mpl/6ZiGspW17TH4LIoY2ji10mz4IgLy
4umtcySURy9sj0M6/BwhFJOLeSuMIJ5Io+TlbkrS7nmSIln8zdPh8poCmalfuzzv
dKxLV+3VeO31IpMJVHM4A/2GZGavZd4Bp79VAuvFoTa2p4EjHG511U7MzPpd2rvh
QWXV+Wt29R8/vU7OMSXjJEGrbhZzjZ74DnHVZCYZSrnimsXaDsrOG1HWOpJjb/ia
qMGmp4wRWH+H9CdXrvZBEbeu3/3nT22fZyn4UAXzjFMZKKhNed0c2kepMzw4Gh88
fauVBWVpSdefJZybbeK9cju0x5/dJ5BI8cJXfEOTNrk0GNjhS12eXHXmzjRicx6k
f/gWDwBZhvb0vGaeXtYq4mT56LVtLF0koKyAu/hUnHs4XRdGICdzYkB/FYM6MHIp
6v6syDvdYJiBxZddH6oGP+Twkmmc1A/4TV4IU8f+642P/Nxvbetiiq3HbdfAaSdx
9SLU1/y/h2GM6K/1O0s+uxEE7JcFKkWIHilkx+gRZ9Bf0DaQxTp77EnxBA4vtlJ+
d39Yjtg6etJbm1h7x9hBOgn+TeMPZvo+D83vjCao+jf+Vp3xsZfOFlRLNpPfWlNs
ADOHx5lcxcZxEItKVXVKgVN/nOrdV7lsflf+EnUDJNvXijfAEFGLwG4DsNOrzsQ5
RISTn0UBBTV49tX9286pvzpwyl/N0ljTtsxGBTYHzB/zDxlrSaQPGMXxak+IONq1
QLA/Pi31NcGpJf6la+To9RqKJYBk8wf5f3ZrvNZXuA+9AJZn26GG+kpFk+qI6Gtt
qQlmchucvinP9T7Gd/wE7vBMXOY1VISjM3Lt5VQEpGq99RI9mLCMJLxulKIB9h5j
duvHBN84mS8y3BXPwhXqQu6+zUlYVVcTsaw3gLeKNzg/owG/DvV44ZZqf7tjt+RF
CRQkglh923VaoloST2r2vckapHxTPgU9bgUvBbopslsNcfTM2ffDceu1p7CdV9Mk
q4Qezd7W8WW+dVVSIP9UFU6VarrQNbI70SyQg/3mk3YG6fS5PP5ZG8mPuJEylNX/
FXHvQsadd311e3IJRVJdNviQ+x0rStebd/Enyk5ypgT8qmCx9LqQYxsCFIoC7cUj
EcIz31cRuHEbQmLc4b6n9yi26mNkNdMKkwtncN27xgOwhCbQdY12s6Kodp7LeSE+
CYyWDQxhagPLhsjx4TknE7J/Ol2VuvM52eLxeYzYomSOP2zn5GQDyVYii7e2zbMy
xsP5k8ua9/TWuBVCMNnQP83FPce27YgJVQq2rdWFTLmPLAqi+/FXm3SB6zS4VVCC
JE5DHfUFKsXO0kGjG4G5uuodbfcexETatYBQAZr2LovroL6z8d+0MiG2K9EE/vXP
coClR4TDeFAIcpW/dv/qZx+Cr95DU/yFLN8jgIsUiTAJzxLlMNTTlkjSxYEkmmlk
pCwjT2Ku/Ealr4evimNYC6/MLRXKNfoHHCjXvkt7qBpcxOhKK/zkyf1/oI0MUZ6x
w4gAdz2vmxM1FYJe1jHCgZIbEs+DaV+gE5NcKF6GXzHPEGJiebGe78CVqJwQzkgV
s+NWmoya2W4GEZ60iQeHdvCVN7Tvk1AgEr/wPLxoPs6vy+Jb6FK/XTpB221o/4AL
6nHJ2qux07r04WnWC6Q+AJSRg+ZbdkI0RpfwAGnNQSSZ0iQyGCbBw+YPrd3NVJIO
lNN/TwZmIKPtsEbhybmvECuF+IN/dK0pqMgETSsauLr7n0hqw1NMHLXx2XVnYyL/
UwCuEQe03HC1yC66ytYJ2IzhfveuNNpzU9om3LvXAgl6mmhGfQU7dv2MjKWceRxZ
k5o5TCXpttKPUlQMqLlueK61BAuobmYrdoA459Lw51lI5otw9Bft3tW+fdKXkg4B
QWWhRqC5BVCqH5JvYga1rCtdiRttvOVQ2eHrqDMM3IAiBGY2ep/55XRIgPwJv7kS
GD5JjCrOYl7Bzwx6DK3U2OQF7XYUnPP/UhhjP9poVDP61/hjI4KXChZ9rMqKKvVe
/fI5s5KYdss+5lfwHyw++1UADDcunKO4rphRpCeD0YwpWsl8U3Jrs9fajgijLJdW
zDGWZecXutIUQ0BAVQH+uEV9pTc1tFLqiA74hp1edDpoAnfe7RZ0wa46uwkm/K3l
JnUmjxiGSNDx13r+ER17+cyIyDTlcZuINE3O8DOKYPS3KG00xQGYqr6d1MWSru8k
J9AdNS5OQWi4+Ad1lqi03Y66iGkenlfWLP633S2OAcymi5l7Z3tv/MEkMEMTT+8p
xIJ4WdBxXYY8CkC/3UHGjOMUjSrnS6/nbM8cKWdPYAOPglK9JFAgERF4FEZ1RydW
D/SyZlfh/OnhAKDxQmobzjrFmjfD51Y9ADBub0FGZYZGg4UfE+s4ASTdD035/ZcH
agwHPFvDcjHC6Vwc9aXUFnvkDWpArdpVk+BQ6trdV8+jhQ9saBaBEtkwQ/idWcWx
9X/Ld+HfgsW1xZ9EP++3NCifnEz7CfSP5+pj2JN6OsC93kswwMVIA+0XkpyFi4Jo
fP75W1muoq/nXVdRp47zPc40noY+WbiVLpLjwaV4/w6JU6xGbc7kd4MhgNyi0IBt
jJ+5tit0Ty1d3lwAmwdq/Wjm/zGdwzCtiHtvRE3pS0DDimIvYBfGHUHN6sN3RFi/
EYMZYVPvH+yzO2df3b24p7j3dnvs6lmmnpyjhfcbUmsyc1+pKVEdT045K8ewecLR
pb6vpNkRv2nYLoLQcGB6fzbJvCBqIS/Y5mqt9h420PyqCbrcDb8VsEGehkRlk6Kb
48l5dUWbKNKG3WvUyhZboHcyCenbpY+xsLfsBQye81YG8pa5kELiflQyD+R4b6lv
/rQaVeCYuPuZdO5W1FQZucNnJDDfgwewXgMAGtk2LIDi0dYWBIwrOB2yJcVH3vwr
kasisl8iH8hkOxviHM7ka4bYC7tejWRNZjhLrQrde8BfaK/Qq9ChvIbjGo78vJ6w
KQrrHUjAbgaLAGM9QlFlotVkHcCG8Bnh9FfCT7AbT95XegsA27lWaeC8zurt9JgS
vX8DzK4WddiuoxQlKcjIZ/OLAKSWBXsW0iDzk57YL01HnK4d6JFq2Ka9pIuH+Pey
ewrfzuD+bsevCNMiTXdn48NzLvOUqNIeNFzUZ6pV4iNtMMX9zwP6M4HoZ3trcBXJ
dR+Ll3UuTqOCZrGS0kjul2Y8cTt+zdk6iXId+l+IanDoRrvnx3U6Kl6ixpOt/x+2
JwssVQQ9BAk6aCw0ScrTDpFtW7HGarUW5y24gUbT0wC26doTf2Af0cBdP0r5mzKu
/+oP26fTxvoKnvnqTNZ4U5U/6VSpFiI8Xg2Y6Rl6g35mucE8eBR5VLeTlE5b93wA
m8n39Co1kjDtr7o9gKN3a8tqM4sZUg+/0/3yeMNonL54AHxH97dmrkemoVHRZ4Up
YmDOnld/y0x0IyNe32H+gdXT72+I7EtFcjoxa081i+eR+RUFLvfFR8BvsNPa4D6C
QitxuNJZnUWVJYsLKnp4okdG3ZaU50JF0J44lQ1Q92VCgyVzcV6qdPddsw7g3H4X
rkXfelqoLqUFA9K4g5Oa+v21foYD9uSmG54TZbuj42rmWT1RxuQhaUNh7lKwNOgj
9Pxssu82Wvml0YBlJNq0UcLNuAT5yRbrgGkw7eaLPBE3XSxKeYP7m1/Y4RXQJh+n
wGFb+JPcHOx4bE+moeD0P9z2w7y57DvOflmoulyz/jocS+VucM0UqeL1tJjfVE6D
gmbPCJJ/R26SRJjwkX2mW89Rs81Eme7i9B8AMYHAsPlhmgEPZPnjM82VWKyguI2/
JCab/ACOITtgx1R1jlO1QlT9f2JZRDLfBCj5N6Xy3pDDd8rHUkrgZwRYzUHJO+tu
3JDqy9rjcqgiXZkGemI7j3vPqFaFHwx3A4CQmp5lZ6xWQr0Qz0JUKkdc8h7l055b
MrjeEW6I3tarqai/eOf5UEz5SpOLTkgQ7bXrZyOrPRuZYkgnsRIRAjW5/cS+1P9W
Qwd7ZSCOZQ96dAtmtK1rHbQriyP5abf62t6OEyaWOkhX7CAasTDatYxsCdBJhzt4
Iwl/tahIKGlZXeL8tYtSgfvVey6kXynPqYckV7LeyC6qrHjNBZzZGFaLnMSQDrZB
`pragma protect end_protected
