// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
u+3ptzhp6PFjKDHWV4Mp5L9uWyKH+DIav7OpS3Ui2URX6hNzHP0UeYNIDvYcZb3g
B5F6bCKx8XDvXeBGxDFLpYOKV+bh0rlwveOudASUkvpVmVCZbkIRxt6cuKrn64Ec
SggOcbu7PfYkbyIWFMJ5LUYnlhTfJgpw8+qG4QNk/0w=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 81456 )
`pragma protect data_block
PrJmAEPk/4jGUsUgPfAe6oYcRGkSSwl4IE9Do/Rqln9c3EMfcFISOtp8068wiR1e
tjcYxYLxy6NOteCrzOJc441jb/mooK+UwPfCj5bhecNyMLZi2ZDyDS8jofVZMcsg
eawMpnipugI/lwSujQl4fy3QAYfXVKMt2ShFoybM/5d8wU4pfAGiFjZiutuYeQxP
6zbKM6MIl9vCJtA0VsDIQFvutIzQmr6/So3a9ClhBPH9zPHQSTEOWZuhCVlWsPsS
1FCGpIk4c5ga/NtorKPgKwscx0mYiTUWXibiAUOqLk38eclNB9KXg01A5oCgslFX
q1eIUR/mfzYSiVCZcquTyC6U6SbUeaDGVCyeBEHlsRA4u2zlEmMkq8xfsU68T6Gs
ofYOgYD06vVtetxCATLUlooa9wXmJX0KpVoyW9aBk91Tiv3pGeFge9QiDp2QFaJZ
YkLikBMRticsu7z4Bx84dse+l7g6Gytin/fX+GLJIr7RU+XDX/19/rUlqzkse63U
jzX78eRnJaGQh51SpNOimbrVTQiuRC4nRBBZTw/EtMhzBZlXPaZ2ajejeyYz8rQ1
j2HC2zDdKd9Gm6LPLDOt1Pi9UoMqw6+nsSUNAskPgHuJEGrlv7Bhyp6t9kysTp+5
iV85vqLvb1ViZsYJ473BhnoDjxTMhN6ZcXVdVdnMxay7moCmwEuueLcX/bH5ewcH
SfOqezdQpkMUjlksnRNT+ipBbemfEKEbip4JCATJdIxY15EWlo4IhfUB0oiTuwUS
+4hihGgQ4BOtnwB1T9GO0qot7zPRL4+5a3Vg/n7Q12GANjRPXcr+zyT6zjnmwxPn
0ikuiKE/OF68ZPkn8QYurgafQOLj5ak8lf2NsSi5W2+bIGW3T1WyYLUrkQ2rl7Yf
BynMRAgTmmv9L3GHb+K85urhRINPmCxOzrusya0+vb7wuchecPAYFS1JMV6bet3P
qsmItZQzwdYevx/doxXB4NEA6/0vD3CD0pPWHzy2YDFjOGNCoGniYteMhp08OwEs
ojM9uVkyeqbq7RveLr23H0nLdXqiWH6mh+NXoy8pICbbxEkA1Cce5fYTLhlXxiZp
+hSDk/qbmwTDU3hSlc/uQXVKB6uZi2qMV8jY4OP8y3qyiSHX93DtA62hvOqPDu+m
BczGRuyqNb9lC+kK/QAvQMALcFCCHlsjWv0/Vzzs4AFOUMgOgHI4QjrWMCdEOaFz
7QCyJbpYPfPNglZPttWJwCBmVO4ZAv00TwlR19EWFsMZZaJlSwe7T/TdQDMloH8S
5XluMw1lt7of5drsgsxTwyRW4hw2eO+atk72W5o9ahJpEzKWQUQGdjb0pxnAnDsY
GwQiEqelEyMOA+TQE13vLKvRpcM41DtY7CWcPWA/t4LxPsq2r53vpFiz/BXqiqrl
aXosMTg9FYygXrsSyhYqQdduELsqOSNg/IjkLeL25JGrNQu3MkH9Bh2iX8yJQZlq
R7k90p4PZ6CX6RHXT84vIgacwvm8KYq0os4emHSFcEe6BNUc3tTuKXbeMIiwhGne
8XFluVe531ZRtgPfpXPNXZaLF6bLdBLvbcVaOJsWSWBCbRYBX+WZLl+rJlg3hyWe
lm7qclIrsY9n4z14iVD18qTmBlD9RB9YozDYIHF1m/4ecaFwIMmwAd1MoC/aFKQD
L1QaLKflgQyarHCOmzEmW/sWviF6lyEm7fAJsd+B5Jb8mjA2Nb0IoJrn2VaN4MtC
/JscsY7ITJ4TJwjfNi+rLY4plzZ4SYihqzdCERIAeZIryZ5+STduSnvyyqVPE54R
QUdUH4Tdm9wzCNfB9kD5ycBqnybaaaogfF8zaHOrVpLklFLooQWcQ/2pNPRu3/PE
3638pd/3/R3BLEmW7lKqr2HdMWw+LuLGAwjtbNR8Ej2x0eHvMbjJy+9zwdPjCIke
nKlxHLw6qLe2aEGJvYcMZUXD30h2WkNnOodRkjyoybq4nTr5xPnwzHjyDQZMNNyg
RDkKzr6f990cm/x9ztZYXkP54jX8aDtQFLNOsig4NcOQsSfzNFCq6jK0CfM8XLlS
7+osNbN5rftpHDuZGufqrUYNNr5w0GFei+vNjK6IqwnUmHFVA+TWqA8sOIVBAnfg
NuXu6utGeXF9D2vMIqamJ9xqq1rKcI7lb+GHcSlTdpBD1OzyCixEmePwcohjr3nA
asPvm/lq/3AKTgW+oVtmf0hH/RaeOkmaRwMLiEmqCz4GoxMAMd14QOLnM+rt/N1m
W1XDK/d/Nl9XoVyO1BQboH0kSO27PQtKH0i06ZyiwwDJs9O8ZrIzWBhC+HdiY1ia
fD77ydIXVFoXDfF2167+ZsXk8TxzKgGwUHp49m2soz20IICX+oUWVz+s8cQaCCmG
2iy0VkdtRT9nf7WomEGYvmXthwrHminw/KXlHDBajWkxTfm8AJA9PtgAOlWatJ3S
IfX00wteGj0bWyzWVwcGsQM1+3lwKL9YlZxEk8An+FEeMmMUfcsB7mTo6kDT0ojh
yfZ4XIXUcZTfD50DFMBOP3kTJVXjsahpVY2wN/7xbDx8HYW5W9NE1/yPeYMSTGIX
wvOWiVarB1e2OW9el6iN75zGmnGxS9P2Y+8WxRb0kJkU2br82EYBtGXHDbtBF1DF
yxiyu796ZTkuGwPp2N6G90sIBSHaavOKUv90WCKFBLkVcsan+bsfunDhavIozHYz
Co9D6TRUA/Qgl9qMyh5gjNHwVW2nmEu6Mw2GQ3vXuF3aKAsPLTr/v7sF+atGwqBb
7ASRaVHe/VdzzTZcGqjeIocW0r+hair9H67yjgB/komFbBeMu08f2EsE4e+MPHjI
KJChFxXfUqDcIICGKD+PyE4oOsKIBRkyKAEYbcXPjthvLPnjbfetdq0QWz4IP3HV
zNj/CWSglY/cCtu8rCIwVl+EzAgUF9KLEaNatvfYGrYOmj0+XmHMP3Dq4QOy0q2O
T674412YK2uCrvp7YirebZqGzF+p/w4T86g4WIiW1NrTbI3Ty4kr03dtjCd/YNwU
4sA8F9AxHuDEFdJbJxvcfEmYoAk4B/hDHbehTZ4mk+zH3LnJCtXWqB0WvGTTGoLy
RIezZjQmDn7N9mtyLeTUM85NZMbpqQTgtKShSqwnPaIbZLUUyLZJexKpD9TL9szL
tUOZaFGQ3X68AJyGMWb6EUXeVF35BemSDSd36BU6U7ihrTlNwbz9U7qzsgUBaCSg
DrMDeSYpTpd6T/krFjmEgaF22B3I0Yjr1H8eRD3b9TgH6yLUjbsWdtpELIk3RYdM
7C1gOnPQjTMIL6SrrC1hpq97TrumOwgO+Publ4By6k8MzT2AR4n5YcW6dFtHsx6g
RpZuduw4o9Z4T/w8pt26BuwOlpwJ2aTJJM99TIm6ZoVLwTSAwAgl+EK9UV8wShlU
Xc4Uqdf7PTfg7sMX0DxzrGsXiRTx/tr9nAcx58AdkhrXkXKAYg9ehgtrvPHYVdhL
uYM2zR6tylEEvHpVUORqWKvdB5FlLEgpubVPux2kmqLZTZIDx17OAw8KB4v4rp1d
Dp+0e21wJ0KTl+XfeosDo1el3SrbGCZrw09i6IzCDYziAnQc0EX37jjM2PLq733D
nr0kyZZ1414vYnaqIZ/4OX/EM4V7Y+Yb+RuSbnF4aSh22ERNSIJM5c5zLoxAZKe5
oySwkeXtD8qPC73z6dwnmKLlxfTk8WY3h6R0VqI/TgyNuG4G8WoYOgafGrnP4Wig
fEky7q5uriWlwsiOn1qTXbSfJuiwM9Rip9DEyFtZjshnI5xE9ZoK7pCOoe5Wgk51
1cx50dD8EfGca81IPKAjOrJeVh82wCVViNDgsT26ps0UdKWRBB8kGJpaye+z2qYf
EuORTmV/B859+V1Lav1cXc/5P95ncFxaDFoT3sNcOAyHF8uZIh0IQgo/l0JWYyRg
BTMI7QJ7vCFdaHOf/wPUoNCWDl1rv7ew96RsWrPHpILmuxiwz4dV2Zl8qZNh3AYt
TluoUfOPe0dM2LLQ8WkRpQhFPhxDWWIkGgynG39Xz5OCvbdY6TqbKbSaySjXT949
S7c42CoLm8d5NzN2fXHc8jpQS7GwZfJKxqgDS9BHYVmxx4Tlcdd9l6Ps3oDg2Bp7
5OcWAnKAmy+V4VsZxNg/BWxLv679wFOsOjQhDM1b4tZ5douNzkjaSXpkfEW4Ia8D
At23RlhZlk7o0Xh6a3jlkCQb89gT7rTmO7NBPzMWpA0nDW3cLQLHlSrc7EsLFG1p
JEXBql5jq39Jj5KXFFebSG7FKyi5PMlns++sD6tXOuv82HcLZjX4QoZgpPV/nfAY
KWGrMuOptUujcBAfPuqCs5Cl/Q8rJBrFPONWJ9Xv5Psxvo5z7qHt75TEYucf/Jdb
Q4tJNjUG+sqUnJVaCOb4EdaGwGx8nHZfX1k7p4I0BIr2PmNRUBRUjh0Og86DpMS7
0RbxBYuzQ75e01ZtBsRmPx4jWt4kV/ZJJ8NzuVcfPLiyc7OOD3BVL2GUScHxP8NY
VxiSdFzvr0mUCP3izldmuahDqU9JTBaobQYDe269HlF6CYAGPbokUdgOXyYDvOiw
ph/Z7FMuGVSPb4qC0xAk7R9vfND2ONlX0UxoA+I+Atq4DNhHebp6BekAXxWkHE60
x9tb0W87tLJp07Uf3S5irvO14Kyg4/TYiEceBjALaGpTEN0Tz0D9DXG4GNPK4Voj
liwt6nd91krBgKr9kXWSeFBaMQ8okroFadtJqzd1AFOiAemj2OPT5O/voijDbfoC
Kd2VtyojYP3Iw6l19Ria2TxnWy5Ut+eqps3AS/BQNQH6iz8Z5coF1DLmk5G09XEC
we2zhau6+q+LPdZA8ZDbwkNQQe8RK1QDlE51OINoqMWtdW4uN1BYYB6MqHYauizq
4/Rh8JbhI01RSf1R/XST9ekUQvOU9nUNfUrPQsriaQwenEF3/e1aIrXVDRkKP2mV
dzklKTSSO/gpA+M47OmDt4vChCztBIAvA4A+jW2mCAGSqsB4sNJcuf/9ocn6uuBu
H6FvyU/L0SVJJBnhzumCfXNd+i1q/NRn9PG94UQh3VOK7YeBlAf5A1cfz+ohJcai
3s2z3cKcGYHIABkRTOIoDU17SD1w3UMLK5UySS/m5wmCX7hJhhFP/+ANRJ/OkoZW
UeaLoU8hdX7NyStTF/RUjSLB7xETB6ALMNz6Aav4Jy1EWu88ionCXQQZ+ycY+9zY
lPp9J7iftkYNPYZZpq6o7RPh3ASWCIC3swCpxljfzfk/LYxXInKRMN9rwT3OjwRv
AcFbGyUc0ejqqyKNBnFu8ZVwdkjjSG+JRgFRddZpYbLylL7RK0CwwIs/w5D/2Ql7
IQzujPyhbmD2ftOSczH5Om4XkqeiHvgedDEQ69kyQOl6SSGRfVsB+cVL2+RkySjv
Vx9GUhWx5uov9XHanRLj5ODCEqyUqVjPcNY8GuFkFxrGfwCMJZpkP0BJMnXsASd5
WH0dJ193qA2rV3l55iINh8o/5HgtuJvKCmWz1eq0xpWmJGXmzkjriOLbRShzXCuV
m0pMMXqaXIWkUu9Ld6l3fl0qq5k3SWpo9sZ2pZ/axrKmTa24d55hqhyB3fdTcMpy
edD6acnAB9Q6i5M1eZ7n06hulAdQmzf1p+/9nGo1LL0/4x+oIFznangLKcAW8era
gaytPIT5oOqoOa9rm9neO4w1/7DgxF2EhjlR8PRyFRva7M686inCHBzJpEvK0M3E
uy1R5Ofks9gYmP4MSPKOBs8bePhf4mk1VcN6AjTCNr6zcBFyHWQX0gVe3YzRBRIC
agWffT0SBgnHWxNZ6TLFqo3kkZocpx2PRnY5yRRJxuksq98mXNkB//z8OKXEqJj6
wPmsxUykbV0HviEciP30JAff4R8+jhmv1Tf+yCTwxs45Tz7jL++ThfekUC9SNYg0
GAxqS9uS7VKBkO8ecQGwjI7zbtihf2ZuzG7aweRNT8xj6ukCtBxnW/7wBLlggmwZ
TK5z5BrVOwTo5pmSHrzRXKmmmKun4yetPme9UoTi3Sd2Icheo0N1nSZP7IcfSupg
oHl9YAy7N4HOjbsovXqr3qzNMoQvvVgFCwPs+/m4VCry+wmpjEJPZqVhu0zQpuZv
NKkv/NycF0k2WiE313svttRwXogdaf5CYn0WQ5B0KA+53EDkIfLeiD9fipSxPlE/
EOC1RtVCWWcFCucNZbRGh1wwsOLkx9DcNgqhrfUO5VVZJlUIp2BM/R9UxMuQqBlO
8yj9PRYv+5mXVClhsWk0fwQfirtyLip4/i9QIbRLTgn+Q5FPn4CHHAewZNn+mr/k
uCPI8pzyvCkvHchp/Ao24zFjWDGRNJp9VByv3TxjLU77qP9897eh8bX6YzLofY5z
v/OG4rT6FZq4+A/Swtjef2RHav0aKFcEJP2pdYEnexgc0U2hEXF9bMmInLAPLO4+
gzT25qbH7b+e8JnD29kCdYDWaY4LlpHX4RFVsKMt2Kn1cXUgVwhPvafzapVS1L+R
w3fTbR6ndd69epXluQ/cp78JrKltXxYS5h0kzVLYzDh+vXO89Y6h3Ab3QYXhKtIb
TaX9nM01fO8gOSHJW+ME3ww2rKduqc10uyNjENbq2C0pK6lNRG0yxrDx1nYdZOx3
/Ois07YmBYvzJ99QgHwEW9y+NTLp+J03ejqEAX9qo5fB2UkChDmsiGbWPRXmxzjD
3zSlFrlNuHoVwbE7OiFlnru9lOEd3Ry+Vq6aOcXIrcaKjiEq/lJhOyBN/QIfAxvv
3DjupskCZDyOwIkpqPI0aaRAVXYXPDnDgoQ/Crz1FyfEdcgM8R+cwLI6oBt5fe+o
NJ9xf7QTtVsYc/0kclaveqIajkfYhsQSDTZrDd0l552s7xP9mdqVLqPfzsrpGReA
23jM2THcK6lZRC4vka64FZW7R0UE1brQAyw0bX7lFct6h03w6DdiayI9C+MOBpQn
1c9epmngOwulXQq53b3PvLjnNyJtDWkxp2nUAQkVfWRAkPv67C9X7wg1bh1lTf2p
a58cGXPlUNYYAxHHf96LstEvrjuuw84LbfSAzDq3ZBbggqT00X1VwRbo51gmTEXB
7Jua+xoZfP/QsbwfC/1uF0Th9WErDel4PTeS8pcnwXFWeKjwXUxfqhL0FFv6RXlm
4Moi+Wr0dLX90mAWQez1OFtvOqGLG80Z7Q/rPnn4Y25P0cDtiYNp4+NnQIwS+i89
fRJ80b8Df4kgbJxOiLEa1scapx3tZ5tszuSCif1rVfLd8XA/83CZbAgXZYxp0dWA
9dohLIKDbE1nK5T5VJLZiLAl/qvzD8+IDAu/626c6bhbktJDNifB8qI/mil/VDYL
NV3p4ks2bjszbTI8Ods/b4NmPFJgPRWJtzdds/kuTZF70vYUm3imZu0FkbGMDdM5
MzpYf2lRRpQspE5+Od/eCs3TMdRAR63gz2OXZOOEaouPNjL5RTrdDXTGt2PrciZ/
aqhkKfqM4PPjvyV7yOaBCu9vDE6Bnh6nUtcjUhOxDxFPXoAwqoUEol784C8wb+++
hXncRupgW4lSESbssTf7fLV2x2ksoy5VD2fxflsijuxbBJzwXfHlcvoouRbEzn/L
Wc91rF7HYoHeP6JbLs0/WkPg4ddWLmkeqf/fyEtvMJqd3go7YT/PxvKZtgtZJXGW
XcVcan68xm1QSe6pNMQkwHHwb4Zu0u4pvKA/Nfq9ssKuoqtsZdwA+0LUFdulzko8
/JP/KSnMFyr1jxgvOVsJEkGdQJeh7JVqIPFCorOGQBhMI2mxCet+YhUCReH792Lr
arA7F/ttsI91Mw+k+31okTBtBy26yRnu1Ql+tsngUx846+vw8kbX1eI89qbF+vU4
MkuQ9E6eVKH4x1mAM1b48cR5bK5ZHMZnhkvufcBu9Tfv2e9KFe551/8Y5yx3KsSE
3Z5hDz92jSs9lhp0/zj8Rrhj+ucLJkYVdIgsv2c8uChtCfj2/qeh1UJj2iq6bOun
Czp77femQx/s5NJfbII4VEkRdAHRUMjVZkuKhgSStOZ2MYQb7S4uvNIs8Vvld0bJ
K0GJgPBCYbDWcssTPO6B6VWzbfl7XRUNKOXSBR7oYCglOrP3fd7w/Wy8uXUdI6UC
4wHMZFnVDzDR4kM9R9wa7nkd09veI8pqMPmm8Ks23DGdgDF+jJrbDABNCgSnP3Wb
8wmYv5oRZhujgwLxfvcmjnYWc92Il4MnHFIt5EWSGQkYSvNBa8iMrtopzDx0NkdE
crkwKIduV/NPUumHGxeOaiD/9MrFN7uZKKrOyc0guuS1cYigrzlZ0LwTUhOHKCjH
AbW4Y/5F/fVcEi1SKtNm9vv769VUuTPgPI1evx4BQ8m1j3nqvQsVpnowH/Wyd5Lo
JfppjdZIacn7SWvUcIi6t2wQCr05Tp7s3yrzA4E/E4RV6AhTqE72dkESE43PbIfw
vFPpTBYrOhOFTmxqumBczJa/gye8nfXkAyNKbTfOcyP9XGHCtjp1cNZ/oEL2qw4r
MGP2S8Z6cvGnoFyDoIz4y5C1TFdSIV+RJ6nig9jnUEvIitVpw5XswlYmHi+p17dL
wSb+ClkSI5v+p6wOUIZNne0I1QUWzXh1eiycXoXmMI/Pj9osKeBY5fURBphOwuGe
H2kqEu98MNSEXyryQB6Zw99qB4/0LTd5oq27n8WTtuENt7Q2UYuZUhL8vHrRUGtK
pjxYFGpEOM4/dNOuifzS7EDU8v5N964hoEJgJHfucosGyzpP05QNW0GbktCl2NZg
gkOiscxpd+WYFhbgYL6bnoM0W+bUSk/5/owChaRMa8Xna+3BwVysSk9lpAmUJSk7
CxlCXdumFyg7Si1Sj5nFxktUTca8bDcJJ5AT/MOyvtlh2Yfx6ZnHKKFtk5fd2G1v
/Psu+7CFdEgxNAa2/G/LpDMGbOO/93U5OoaYk9PI/RD5XCsymfqRydWv0f9nyMzq
PDdmFJvLBVypCTCcVhxvfVRNblAt0khkXcZ90HHdVCnSWlpcw65leyNjIZ45ceU3
FhOA60nwTJy+zYCgVrPX+PBib/zfDEoFBvSQYaK/yQqC6aXYopWVpxe8vIAaqIHA
evzCAun+H1sUHomMsheAOOocNu6TG/8wTp0HXSyTG/5PyiaFwIDMJyIsk5rrx+eY
WzIxCuMbqQCakghrVB1mAxyykYZKCpHCyVU4+aTQbVFQ+ZLpKfprJfwZpAFovQaJ
wgRSqFtDZypkbpDxEz0SO4iZUhTFE+tZnmUVh97LeuWAOegcxI+JXFD8mKz4OF5U
NtLdxVgZxH87k4os/416PEdzZyH36pj7KPt2SzxkOsVY7jcVrWLR/27ekJoFxDBD
B9H9kqsKoRVgEYoTA+a1dpxUanCiCnAQ9DAyzVfwCgooL6qZD3weoNTcGUb7fAhC
KuO5JBxNkAyBsMOEZS8m03uYYS5ySH28JcWEpClMZkDCngDcYkcrmNf39gdDbxoX
prWphK/GI/nJCtAQadPd0y9SoTiksMYokMDRHUuRJpMJqXZGvTW9qVT6fS6IrVXS
0j7C4DyXH0vzy7XsgCfQHLCUd+8Rjty8TA9okEen+xyAaOlJpPVOEOKN/0RhuvaG
VmhzxCcCrDOAYr0NnrevRPZDS67Vbzv/iUY87vtclXb4hvCckz1OS+DTG/PmUUd0
oWyDgQ+J6Ci102n7VTNmamrUbSzSFv0+jGGY5wJCNdWxyN6U3Vk6UyeRYcod39mN
ZtdzqDKHj5s86HNgEiCR1qNIljnRaBCtccz+79Z7u1XshtuJUIdUpq35W7ALldjA
RPAqMY7zycTo7X7cxetb12hn2hdylRJHE0Defo+5Mn5Qy0cS/SuTk05wSWpW2vrx
kk6zVvEdVC9JFjSez9W7j6ZR/D7CxgANgzNtGnIVrPckDV/rctoDk9EH1qEC2PJY
IKs5ee5U+s63ga5pH4pJvNmrFVft7u3s8vpWtFJureFylytrqHsZ19tj5b1t6+Hh
gNzNQwNwyxMgLI5rEbqGMKtQpjBM5uM/05iox5Q1Rh3f8sDcjQm2jp2edwLfl7A4
ip7L7lOQMgSIaiATwT3dxUG0Ooh2XvFFt7QrVYYXAei95LtbZX/Lg0sII5KGfnPL
XiImk1FupLgE2bz2QYDtwRppzvCN1c4k7ByTlFclJ0Y6e4u7LAhBa9rSLkUa2J3q
0MzXU60Gi91SpLB91s5SlvP0fuEJ1DzGmqqsbpyHV706N1adBHbyGq8+rxSpcGIT
0aJrL13s6PlqURRdO4mlk/U3WCeEuW1Zk7Gvrf7K/0N6SJVsZsTDoZ1QYcvORmZ7
qfwkh1RRwvNA7F2V5ki25zNIiXCxiU05mLdoDMz/ndKM//3MFWDzgse0g/uTDPyQ
pVW6okZN2qKomXJA1MQY8qfhWOOXtKm8hX6WGqk8AB3eU0iXX37PlCk3xXzai8R/
+8CMerJATmHV8Eo1kgDKT/NfMIfUaYAUiYMHde0aM2tT9CrZoNcJ9AaFQ3tT19w6
lOIqA/xQjBlWrGacT7pWDlqjPjzgr+imCpmvThgmedaR0uyTymuJCUAUsyLbotns
C3SuEUYZ3YAHkusY+8rrpoVpd0vppdMSpgIsvUic3QwTkEzzSHqfOt3sAMearmiX
3r8v1JRFq0QJ1TyfOXON3GnLLE5kxwyU+mUBSAvD6RkOq5tudXBTT0C1Z+41xTW3
hCzlSO8Q7XzEhA9QAwFTPNHTQPO3GJVIvEOHW7phnPS4v+34j7S3IZ0zlkK0rFcn
OXw9Wmud3WTojHALS+SJ30Ltf9rfYLtgzugfftJMMPANY7+aLUU7LtT4xs9aSfeG
/ujKeNdkpzZVQ+buZ9X8YnPGEXMp3Gwe6EGnBo3EcY3mqlluwjxekfKGTCk6Ia5U
McPIr6PW6CqetgE6fPa/TdeIHEipqo8dEYNC8i2Pz+X/lzVwXZprNInrFtg5cCER
LUs7Nh97WjLkNFdnSWdjIRy6rXU1bMXWQVXiYbgeeerqGVm85ayvzTT+DN1fh/S3
3bpHalZf6s7HQsgEH7NiTO7Lzr1UmKNwlRz+J5b6FAD03VNRZ/L60fla5wzqTAf8
N4JqGyuCaABa8vmnIMZQ2BTO6AC5U4Qtpud0wtQVBFiwVPmM5wo8JERzIBwEG6gT
l/vV9tF720Krqq7sSju/YdfIOaIM6NtCBxoZnuhfBqcNEuKuZqG/dW9yP5PELTkQ
20ATBIOX3b+SZixRnwjo4S47fMwcnOBv3nfOw8qjHx/6IrrYnoLB+Eh+HAIalY3R
u4CmqOXRpdYCJPTxltR5Dg9o0r8NBvUnUeDyhr+cEeJXS6c9l1t4HZGQUfLKZQSJ
sWQosVXv8bkg84uUhN2cyO2j/ereWE0PstHzziUnuKNmbLkMAgKwb2cl2uRCY8Ay
xZDhGc1zF4mNY+kxjpqTyaTb9O2hfCCckSgKt5fn2JqKHbypFwMOa8bJP8K4VKdk
MqC7j9IQdHiNriyzTlWMJFqwEa4PLrGAPm4T89RYZPLFxUNx4hyYDcxqsJG1VQNr
a/U3im/XQDER4SG0hznd+9OFwBYXW/X6pIVBCmnqHFtpoW41wjgZLGm6t7JZ6X3o
nujjOdjG8Gbzxusw3MM8DKTs0ZGax5VTSZlaNH/g6i4o4l6kPevwN72ozxpcpRt6
pdtFPw5uEx7MtF8BTWAH+USvFfp1+CK6bMJK00She+oq8yPU6sOSMiaG/oUXX3rJ
gPoTI081d5Ga1QgzY50IqC06oNNbLUv9U8UWl8RS+ZV+LxQKnM05pJjQhtppsn6H
Ia3CvmW+trUmBqGkS1C4A+HaatLENYNjTQV9Cwe5k1GHcpS7Hh+7onkiKsaOfm5+
E/uqavI6dQeP9fR3obxbDvhifhlnRHs201DzeL8I/D3lO4mtnJ5ofaQ/ZWcdJJD3
tSyREKdmy/Hg7fDj/UMPVQm5mHEBpAlMyQJQby7MwjQfo3CSvjxTsyapMvEzzTuN
9D5GiT7vkUsXKM2C+jLlKfAcPbe1MSiVnAf2SqDqbXj46h3/Iyxef9Xdl4Fn06Y+
JKYpe/RWtCmwbPkrDuYc5H2PLi54Adt6dpLK1/dsLuOxTnMz2e5SC5EITratskrV
NbdZV6fFVHkzp9Mi+NyXC+2JTOrA60WY35totOJ+wikK0IatKQmJ+7sj9LQGHRun
zIp/dmwrg58vwTqe/C/95ccR4QH39j725LWbwdlZm4Q2d/EC6LO9Tj0EBINcaEsD
/W1pH8I3rnN1j/5A6eMFPyD4HaYbBRYdkcwrtMr9ZXpPmHW/J4qhS+Bmewtz2gl/
Ric8jJy9ZHEK0jQkaL94u3v4efZZyK/Crkt3sTrRPrYIuZ64WW1hvn56xqNGqp2c
7Yai2uebrh204fs8r0Kw0v0Oisyrarz/GyrGg1XxcYWExc8zBS/FAS3F5w2Mz1XX
aYTM6iRVnYd6M5f6G8ER+AuRz1zXpq+IaWtt7AP9s7mH1d4whJPSECbg40KZvSf9
IsBNninqzUpNlMhCPlPQb9pT3AT4dvBBlALSs/OBD8lb0b64/sZBWpQam8Cz2YxN
btAjZ0WxYsyueX/DUzwQ9eQd2nfQ+U7JdUKCLVRTig+Z5Prx7a5Up4MjuXE6Pmcc
z3Oo/HoxdW8aDwNsSA59Yzjgz0eFly+6j0RIS10Yp/32tO1x+9tMF5Ndqczbi1R2
DkZ34TGqWHRw8oJnu0ZaDtWX5Fr1sdqM8l1qQGnU5KHj66kLvE0ScfSGHOe5OwH3
WL6NMHwYvwh0yh9/v3Si+OZwLWq7jx/FAZSHvm+Sntu4dPGX8XfAwg90nfuPmqvA
U9zBJPDDDqdSfnWDVpDQWwvZKbDlNlvRCGRbqcu5AdI4QHUUxO/94nwOgd0qqOns
00fMo9i23LsZbocNOIWDJD4N5miSPljsRTYDsieC/xC/sU82IhDKZPhHMuNBhltR
9GkkqyH0KJUTlu9NlwOcNYY2AMy92D4LF7q7URPnCETMjaWQN9/UIkYiPPZRVifS
BQb647GAoxJmSU1eVG5wDe81p+wIwpMXidTlwQi/D1HAxEByT+8/mEjUASnFzHmr
0Grx9HJk1ks1oGR08F+xq9QoJwnZA51PtgX/kqM6PchjsRJGXEW+aP4L3IzYXCR/
q9rdx+p4Of/72sws/Wo7VIvvCn7pIYOMe4JiAdGCrHensRwWE470+8rnwLQkq2gw
eQtJibClBzcHtfmsM6Cbb4y3FNyMPg+EWNKMalhp5ZQwyhdrQoXiB/eO6LAOYygm
dqbQ7OfObk5gzFV9EjuyfFIvpQXMEkxhX9jBYoI7la31LfjY7AOO+J/05YkxQVDe
Vj3us9VBgIL9c36wZGPsGdsyOsxL8zvzQ0wt5dbJHS6CCCfWhwbTyGFZ3Qd2bSva
g3KDRqE1TFyjMN3UcUtrU3X2kItft15ISJopvFHmPUC0kFxK0sUqFxBorettvwdM
RaSdBuJMt9taAH5fehRbSKDvUIwtVcQ6RIpBUWyMzIs1LZyrOVSrFe+MfnlYCHUT
EVBZXnxL3OI/u7hj48vOJQeEr0VfX2FVy3oc/y6GSlzxxfRxZNZlR7JnRR1n9hRv
m8zp79I57r5O0S2XIerbIOjr6i15kiEDcx9G2S6axAYRr/A5lleaL/TzvlElBUcy
Uychp4+sip4EBUm6Hzt/Ncb4k6p4jNjJVqnom5LOLTTRrOpbOLA7SB9AYBhRwxvi
kSVJoN650dFlZpypl50UXk2tx/7RW0JBZ9c76xJz1cvStcVzRpcGu0LQFDqIg6VX
JBXiZcerq37rb3gFBMzsqXDt97fc6bfqA87OCe6WvDe7wQLMIGpDQZQD3nE66IIo
UZ/Se7jrS3I8C20gy+0tP4UoCeLpPB3gRlucfCY/8iNZ7L92CzeAyv7/WWCpmaYD
JODmW+DyFFuW6nQ0aJ7VJNFECpp/joXf7ERE5wTw1jU1kwOdPPqgweUnkrLBia0T
Vq0z66nQ/GH3qBSSnSkpQFw1dqd3p4s/pOm81pxtiQ/2GQwZNUWDu+nsyFnW9jLr
yUAGo4ZrFHXGhVYRJV/zWYzTXxe5KXAelf7jVlbClIvBXnb+aiUpLBjfAIyHxiOd
84/ruV0Vc/28kfqsJTFCnVxs7kIiRIqkxV1ptA4v0vu88s754VjL69P3gzU/9HwK
RsSNR7mP0prkMgKepadfxd46EZq83UxMmaIc0iStVQaxTcYVNKt0jlSCVpD20GY/
EPdEnVhndicSQkhdmPPkFQSRKFRXHJBdLF4MDFT5MxoGOXWjDrAcNOvMFHu9iKkv
dSr8NvIOu4ToVrwP6pQCrHkE6mr2NifFW0pG3x1WW6Aj+fQnyPL7IHsLP/Yl4JK5
a9iZ0e5WgZ8pvrw8sfiUDEkX32dIfEVWC9vbFsxTw2vAh4TlhORE+xBltLZeuUHq
8biY8x/8C5D1BM4qu/uhO15nME69R3F31z+o3697DfF3g1/BqtYaAB2Li8zuMdLb
PDPWKMigkk2PQ2PikJgZhcTz7I9xIpHv36auvTh0GMxfrAxtoXBjzmaHAkW7Aq2N
E+RzTKQ2W2c0+jq/y8Fl1C6pvkwnW7iWsuF9KGrzILOqISv3ffWirgrbstxJbAzu
Sj0VL4eUEp8yBistF7e/WA8FWLaAgE580mkm17qD4WtyfLNr3ElCg6l2HdJhaPOL
mPAr0tYdz46POAp38n6yftk+B6BbD1ba00B/i1viSwEc7TDCjCrfOylfop39tiZ2
ysVe/WjinYeEsEjBlH52YCw46O0q2UuY8T+xpJ498BzXPCJ5oT5AVUEiIEiIU4XF
NLhJeLuwXx+YnrbTQJId0ANKprNdNNORos3eTI401fMKbHAXXScYhUlhzg/MINcA
YKGu6ggBz1zjDCQrfNrspbQ8ZJvNWnXbztUmWNqZWJy7F5sjQda5r3qBsI9ogdbL
hfnxQWXlSpmT6howeM28pJtD9lepX8NZe7M4VEnYZU5VbFAXDDXpY/EVO6iJKcTU
2BYXWhsRUzFXcbMhKC1KtKMvo8rkD1qAcNg1lt2vqIOf+gEcGkjedhceAKzE0qfh
BhohPqzLiH9yVcCpcJwX7gE7bqG1uL5B0FRl89eAj/amW5niIzpf/K0P8JPagv5n
H37ixiTAyKA0UIsUw1WJmlLbwNO+frOLtG3oNLY5vgOrIr7Lc9PyvXnglVyIgsmv
tCNas2ji9UCuZYVsyJEdqv88kLmYHP0J1VOXSE/ew6kE3FVYGj7ve1YBBXJ9/yJC
6xQh9MgKesElHZ3LIfkMQQVPH8qbVApUc2pEn/4wMdXfhZ8jJzhKVgnhwHR4H1dy
3H/SLA/cpKFcVhx6yXt9szHOhV37B8KeODvkuIS6rwKoZRj3wfbV3VjGw9MpYq3i
MIkKosKTuR+IxNx+Bg8NKn7zNFxwwUq678HLPdPBNNxnFAcQdRkHmKqtbMgmAJhc
D5ahxq7w1RePq54yN2K87XvCfmYwHFhD8YKzljPBOTZowdoztLDBFHRHXo03IPD4
8gZSEAb/dCFmx5+f/ajUc/4iovopQzH3WMwBX2DkV84D4uMMbCrXA+hqsmRyUS5r
lCjxiZtOMP2+A9fbMqrGL/qwg/k445YZVB97O45CbyW9DZfhOKqaoxPOBKgpjI0I
fTnAJAyHFD0k/NsyCdW3O8tlF+JTKxnlzfzoGQr8BPxtl91tvPxaspVrqNcsXNSX
dnsNq8bGAR6ZP2bzZhl7Yz4PnVIo56MIw6iVMh7OV+eCfli7NntSzAmi0xatuT++
WPi9z5QPs7fE20MvkcqSlmygqxV1f/xDgjgHsQtHjya7SL3DUPPuZ8odtQRfo5jp
dBVDU3RA61qZo9/ZMTiHFIx4YwrEoxiPWCeenHouPiFuHPhPQd8KxR5JOHOKeTn3
m5vI3ZesqJHYPY936N4/CeB/yqjpTAD8mSq9jxWPZziD8nlFHtATRq1bHEmrAznU
b+90NlYCCpGP3vUJ0PDgSHayayenK8fqHnBosinJ58TmpQucNFbj8FXYrXWAwS7G
IbfH5B3TIaAJ/c2pfJaol08vVWIM+Dbw4dXzlX9+5mC1x3isiC26wboYZobQQFrS
kOpTWhhL3fos1iRqpqD0RDUS1dQ7WuU/Q+5N37Q7YLiILNKspCPooeznUYscCc61
8Ynq7ccdXVUwgPiagIfD6Un2StKxlu4Iup8q7vGcT+6ec1+I4S8+h+cKn7tfwb5v
fqgSV3+3NP3ab+N28X0HFwdFsekQXa3eauz7yFu270+2Kg7Amn7NOC4rHbnGUBIp
d+jowM734zX9V2/0jlvgu+lIQU5BTnRcl/GRDQqVEQB4AwtJD9brNemAMbE+lPEd
tAoT1WR9rSzUODssyinAtKj3LA80FExOQodPiELrrYhe+xfiuMkFSzYoZKoHMdw7
+t9M6fKMb90ETFsD0yJkk7AyycPSXkyMhCXZQ+AtU8BDK5zgSm60mWBsY4WJ+CFx
PUKV1kdd9pO6jhhUHOsqRwJOqUuOTa8iILkoJ64XDL7YmI7do060AMogl472+KG2
jzrIiS1oDPGrjPJ1dsh91QKCIJFlkcL8kYSKTZKzww9nQEoYQcFDBym/zfXkKUx5
QEhXL6PJb9c8rfbDt+rUM84f5tOuRgVHp+doyRorKqrIDIP67ZkAnk/IxKVkS7L1
wD3lOshcY9Q/4t1wEjGLA9fTuOIOnyHBRB6Tut6vLVApYGs6dryMIVOyGST2XR6A
VPu6OXTfVLIaJ3HDCxlOpZ+UF7i/pR0UNvFiyglCTqyFUCjCD5TL1m3EYllyCcYW
ReP96eeAqMFPYSAmm687U8i1sKaMRkmvaHd6iZKLRm6MSWmXMIasbYwM+Etl+Wox
30IRh/88uP4jUD6a6yf/NNDZX6VG7Cd4OFH/PLVnvYqV9wR0CK+zYeOnaMeOg42q
ls15jgu38s/tE6G1jqmUmdI8vp4paMt6YoKlpaW80LGbZMFKYcMYbg2jhaGY5504
mRPB0bHULFkgxtw2dNkf2n/priEOPbGm09JiAGYhJPTaQTAotlz5ukfHiaI4Ucsm
bKyIvdk/HDmFEQ6sShmkjAuVH78xzu311LVVEvYU2qbKsMOw33m9HIdKYZvihyyp
bROtpwX7OtyO9qPln8I18FoKZKhf9FY897WyDmDa/ImeEhmcYtVcX6Ky4TpENRKq
1KPN06JAz1fcanW96CWtniBGJF4VGt27FrRdz6keUt/9X8FkKa6UhZziXcaKxAl3
MEfyJb8gPFfvuQHflIFIyN4TU00Gp+3ZgMAPCxDlJ5etEA9WIXKjZD/JlfT1Kos7
8msJeCIN034QFpxQlLONikoG7SVdwvLTbf4aFd5sqA2ph1w4nAJ37BxVGmtyrggZ
Lnd5RBKUT6qv04fIl71vZKArqB9V0AL+8aufbN3wKAa9S3JElAmFybCJAW1/tsFz
6/79QFFAAzCXOJGATK3WWpz4NVWlo4c/uHue0IyOVDA5KQdBAloNb8enIES2fBtV
fYU9ofJPk75RaKGI0z17jCkHIgxFtpMqIrVFw5bfXo5SY8TWrjnfAbK0ySraXWx9
ikGEk54qkR1rF3xUensERbVlBpHXUBKmbRajp7uLvjAU83Rgydgkb+BNQrb2oa2R
oFx1vUfz246yDRQCLcUAWthyJ9haBxQ0udlzaz0M7McqBKRHdtswZf00aUt+rtgt
FyyE1waJL6pHhGwop0qiCT7J1wjvXCsp+wtF9TXZJk4cPdx2rGQpH6XObLDb2h4F
Z/AeHRpEGnNqpaXaIveeKaaFZ6phRL1hquyxSTmWj9BsN+bMuBzFTdvyPT+Rw6Yr
cinFlB/cVM4H3km6hESTKwKslZE7ljP6+HdqRzM1pbTsCoDcVyPwmixqKqpITshM
OUSqQxfn1rZP8CtCtVvMESwq5Ylc22sj6YdIDXl1WdDlyD/MkYfty/7iT1z0u9iT
u6AEFWKLc1j5knIR5eVN0NXfIchCSLnMy07SLY8jZJ5oWbrCXRxCUOEuaq7RlCXP
9/NxIbdF9y/SX4K9InGo4wrkeww7lYcepxxi5NKtvwT71ZeafVfP5mbUh9nfdEFZ
ql7aANZE/9TpKDUOz3cZyD/W7ib1oigIBuRoaw8dgDNrq/pvwVzknug3C/DkclIg
eEWpmhZZTffbytYS40hCfp3egLWOxPmF5moAQhlJS+9VSuSRF7V1gmCT11vd0gCG
kJVUEyfJZc+k9K5JV7XjvY63hlmAa1J58eAZ+X8fbidM3gWdRxD7M+812YxiDy6q
wXNt3S3ik0+4odTeCtNsMnMqJgfK3wVdEhRYIRyZWEo5lTUO9xLqo6/c+HBOKtvn
Sfkgo6OLPbS6z/RQRCexXGfKeLbJC8yCxugyXRMQNTpAkqua2UcyOsUdaHLVj0MI
YZeOwHXe3aqPQvH7fg55JKwV6IIBO3TFyPxZxr6ZXCkVgqPrVq2M+3zBfOpORwdp
NCwyVhuEd8phMnTACmnvtkpkI4BATTD+8KsH1fOnfB2LR4HP0fKnd7UNsYEWlFR8
e5OO875wPgO1JrtKFYVC3LqxBX7l+mM/luTbS3Ei1Ky4mxP0/QnwakMEIplNkL96
JiIDlZ1lF5RC4QlxRhVSHpuiRIx0s7613VuhCYzylweAfesmu5NSz9DS9JwCrLWC
aYIsJhOwedWLklPJAtqQ79nfZqeMYa8zLOeJ+xZjMjzHvfmPjrSni63dJMNRNbpv
xtQ12HADcf9z92fGJXZK+v7CY2j0X/Tz2RSIpfiZGgPnm+FibKG7nNGby6U58aCz
1+9We+16zm337KmctSTIWaO5znxlIg80TcDtiVYUBQVsF29gcRcz7cmPjvVBVH1G
+NB6qlmCUlocP3s6Y0DMbt52y3zX5Vd9a1Ejil9IGZ6SefOh3Ylnre0261ZPadqb
A13qrqIB9lNs9MNdjwBQ/lnwpJnut/H8RKeOjNZV/qfXjM8pSkwlv4eQeUwkKQBB
R6sJCiLswGBA1tBi4kE1oI6mMqj7yF8h28+kejeZLOftEUC3mPQoC1FhMHyfcxDL
ycTK5DWvRw3zoizZ3HRktMQmSWQ8fWf7O7y1g4Gn4PGx1byncbKo2iDtIAUNyENP
q0Xh0gJySS/caZPsSOVJCS1cbP/neDNtiwkKC3DfbSX7GlW1iCYouPAKib5crv/H
+0MExiCeFkZIdduRFz6NVw9oD2231d0w+lPCPytL6g7xD7Jura1QgR4R9eOqqOdN
zPpBMVt7WuCg9xCO2XL1Wd91taE6LRB/sSAgs9RLHWXAfjuhUilJ6Dr4yZgWpYmY
ts1i5+sIRvJbga4A3qV4JaBS5iXFj+Og1dGodw40K3DDkzxXxBPht4Foa+vSk3AK
JGzWbdgSPs5EwTwk0Pi/ycoolPsuFUXQsNQ4dNz49dSyk+5EHpyIa+wYsDGrJzqZ
pAf8aC/lIpwwM5sUC7P5QVOTezADGTAS8pjz3MQFL9LCY8mnt/7w4MgQtEdAckef
xU3yrPZyeeK8mPuGX2ebKpn/MaCUhUKdtTRXT2SdPdbnJM834T3t5ckyFu+LRqFe
HWVfu1M+rM8ZfvCizA2dKZo9+eFgO/zg8x4ZEY80sdOZ0ieXFwhNwlTE6N2lZcrT
EAIqN4zyjmW56IfldJkxcWse4fzrmiGY7tTtDqDaJ5SAMEYYIHfrmNEXg9cZsJcC
U6GwYXFL58rQfJsjI1PFOHlezSPFes09jDe2ny9+Vlmv+LGKMusk3aD4jrhNfybX
4wtv7g/F5uOrxLiChiZNfbPc2H9IQVO0m41Y6z8l549RrvkneOflawHdvLfk0mNl
LPKhNuNJ1L1G2lCExE2FdbvL711CJdV1kHKn/Iu23H3uDVV9RQRqYLCzQPdi/A8u
7J4I8j+kQ+TRgupw2uU7UethggtuNAOq7AoVbrNVeGef6Aq3J5gkqdWvgBBvHTc3
/ordg2MabZR9NTVzcXveA4USzsbx76CmFAA7r4R8FVyA8LnoMb8btHm5m8UL7Yn3
cI2VMvoRuy/5t1MarvwqW53wLXxO4y8Zbd+oVice61JWP6Dlo+65uRJJ84GkfzBB
BsovGe46CUCAoSrStrdMTv3xwW1J87ds1tDOTOUJBl+KhlnN6l7el7u571z00mzt
4BUyd7bizZge9Np0lhaB3/fiyombMHoTkXS/8lbKhxOuYDRTP5GS46loSUG4kcGk
vN6EPK/gCK6MJM5aCoF8/jI1BoDMPdEpZAZC1UC7DcXLhclAx5rTzcRRYmejJ2rJ
DS77NYXn3p/gp/5blhA4Rk2/u9MljqIlVRH3lM0bwNHb2xaawf6fUkvDlniI31L6
Yww/ewOJXLyMXiuOG6N7kgQ7QLJHy3WoIVUhNJjYRX03E38YoF9KNw70z+hEUR8i
zaCvwx+Q/ufc3t0pccEo34/8MXNyQoEOQD1KFcARTXVaNkztepnd+sR9fkXyTD/+
UcK+SUfV09frHiZDVijxElVYbEIDmcog02xtUPukBH9ZwT/BNXVsD6t6Q8ec7bti
WxXWwjTcrKu80evqlE9TysMyFDcbNIcxPkajGgnxu81Hg0OuAP90XomUZkFW4mzb
7JhxvmELRl5rmfhdOg1yBuBXvrCyT9pFnU1WYqScaKhJ5OfnNYOfUs4LZZflKY+1
Vr8UN+pVeiCtPqo49gHxP57FpFAYfpIsjJ+gANxkgF2K/0LwEgXWTkugwaZ5VLH7
1i4TUalJnUwH+FGOm0zMgN4lFMP28+/MchYa2M0moUWAIUZVXyZkW0lgUnQDnXM6
4embR8l/fG7+GtkqIJyNhahPT8vRn1Thtea4kOvTjntX6Ac6Ht4e7YWn3OfWXYES
+U3ng7xqBmKUSK+aSS/c9vCvuumlfRaw+FIpEzbXiY1ATw2y7LcO0tkLH8hPcpDm
UAreDo5GPnZjAs4mrVw2WJL+xwrQI6S0kqKWnsuDFGfvYOQJH2MHUMeA3/w3vWfD
jSrhiqtyfZLlQqXabgV/5m+f5MBH7nyZM7q/4k/Z+hTEbBvtOmBvqhguTBZZLgbY
nRUoGjVYvoE8uJ0XfFZyK0Tgp8cRQWY+bbKmcS5ydBBgXttEYCSpU+AIVY9+Kc9B
0UfEpq34dZTg3L9CSJsEWfyFssDzjos7goUmHlCBAf4DrJuSiGQq3k+8gGAmXC7C
MZWGpL7KvdatI++9n9EEWJlyWDsHP5x+tJcbrht6X3fsuBJWH20p7/0AcJLAgGWi
81JtLsOGWsuViOipWN6RBFbYH0IXz5bc3blzDVWFj2KHOc2kNajLABYRyhzcXBC0
J3b7rWo53tFq55Hn4b0dzTRl8mc0PU8hNhO9GyzzSTeSBdt00xOA0fpMC4dfvaC/
TO5hdOdRFkOSrxZHtKQNGVqLbbyx8/fGWsT5YEEZ1VmudOmzsrzRBRWGx4wmWc2b
csHDVMLOTvm6jN/iNPsiocnD4g3tdc4YjjXxun4b6W+AfJTiF0H3C6cTnznQ184G
loZ6HsbylBcHOUG7Ef+rkqpE1AmqGhwIYllP49Uu1jcSrtuQrQrTkkai73JFV8uU
9YYRhrT1DJHCm9Y6FiKWR/8BFF87MBmjfmEIeiAMvev4chgCcepB8SA9qQhGWTjs
5biJ5CDIGBPAnqNlgkMMFze3DCthtOQLWc1+05XdDPBsSeZ7gdJU/GUB67+SOMyN
vVSggKj7gsbdOIIsHu/2gbfhAT5Rx+BGr9rG0r+JSlfSEBSRpeADXI4irRaHFcyM
HdM+eST1jn9TDOaN9NBKl+fA+3R8xcH2+KRYy6ys/MRe1HqGQiL1JX1NNT+Z+6OQ
8k1v2tTvXdfRKosXRQ+pSk06Fi27W3vqawV4FIcscRum9KuXDD72XA87p4/8AlsJ
ZDvHLiRzHMnpBcw/dK9jw7XSJJcP6Dqw5UVPnAXmNVNgziyWaGhY1QXcu9Hn2lyL
s5L8TjZaM49hTgqrp08PdbXA+CCe/tqrT36u6ogkJGOhYTXK4GCr8bOBAgOFyZC2
LsKGkRBVTclLbUidTN+Mf00o5CeG2OD0Kw9YttpPA3YcdCTiuvFNHCp4Y226LKNO
+1GiaEBZFsWT77S2sRchhsjvT/dZmjltQN2CnLXFUWZzdbkoL0v5igZBJd8/w8fS
/+E2WCVEt+FmR4KjGYBEV6z9exuy88otpsFTklv1b/mINccET1YGRrOEicn3tenP
I2j6Cz5LTn46ODrsJzMvufBboSncNql3Z6rGq38uRBhpM8oxTGttJlBq4xaYSDFq
CVY7bTKBs3M6iZ836WHY0HkE3BDzzqKqx9tAcFD+8r1I79aKtAILAGe8pC3OJEW9
vFdgnYcKEVcDXTRASF1iDD5JH4yXYiuZMxqYTp++6nDEGiWKx2CHzqnpRYSINzH7
bmM05nk9eSYB68TnCvJ1Aw+uJpqDk3QkT4ykZJrrajB3HPNrq3vTMS1moZQnumec
NxmA2eXTR2IIyz46YxtnUz0ZJPD4rKfgxdRRhQR2vrsQxG0hSyybjiz7nZyt27kS
N0VP3Zby488rWKksAVdvp0rrVRrP0h7fUB4to+beU3nF2SiEQ0iFehSgPj1HvJun
4mHbyFk4H/bzx+TGVu1AaNSCEdIefUwhrjzyPtuiMuTRdlN3bGF0czZU4UbIPFQ8
Wri0BTRCIq3u0csQLRcHnNXsETeQutS9S1I7RiPPrPaIXd/n039RG6TL2YElMhVB
4SCrwbgkHuZ8xou0Ym+a/GtBpJ/THaq+EnvocrXuatdRDYitBGTsgEWOLyTWDnBm
kSWelX/FOUOk+ZpYF74gcI8ulFXsJHL8eMdRNlCbuyUe8l+4gTfXHRhzVx645u3H
qjv1NVkhQOTvA5yS5rQpZd7GN8ZTuH9jDbB5azuFvbNo3dRKbzqy1EWXBg0P4RBW
JJP01Nx8bts9YOJ4VR12Qu8lH9sHPgaiMQMv1T0C+uM1zmYMgB6QxazAup8zZtno
utqg0k3jWmePcP9K451bvX7BgT8Iuw4SmZdtJjdREBwwq2IMrpb5ixD+8Anns+iR
MbM1rYhltxMWpdAVL9bDvKVlOfKsOSsADmwRcOHbTimVC9K+Zg5R8V4+wgAF2piN
OMQqrZzt7F9/qRvVV3JY5qyn9sQ2gFzbC35BBKaX7T/Js38FrBEGdJSAvs+tTVJt
6kddGMB6ydW67B6HkdttQ190HYQ+ZMKgH+fW17N4t/jr5PnHI1U3Y4D6XU5xz7hk
L1zEK/KGwtMYLJcpegynEZIDdR4wSxwsk+upBrs602RjfN4NaLcKTgQoqEPeJOLo
5fOd72T3xEkvyMCAEtR7gyhO9iC8WwEHKCGl/vj8XzaLlovloQW7lCfB1Sp4p6pI
8EWgtNoaD+8oQIBYyT9vypkByjs6RixNEMe5YMXxggLnGau7fncKBz/T1lMiqnht
UoLJS3TWxxh4WR8vWcpiREbTL0kKWE1RWxIg3P6qdI8AB4lbJvxm34xfMtANL/jY
VzpyiOygRLE7gpL7DeNHxazzy27YDd5vmECktzkLFef6GViUW3B/nyIJqPsp76WW
r9NvZQvcV5ruTIZUAAOgbel5K2knyhQ36BS5py7oDJA0B4hx7F/Q+rcSVrhWNqBP
aLepdQrSYbm+GFffzndm7m4s3tqGFHyl18PHZ47ymZ9K1uOOm6sAM+uj16vImn4b
uylwX+zvuu9JaQGkvQ2cO/TBVBejz11Qzbs4DtONrBPPD6UkwUFwyuJ1jDLpO+tV
m+pT7J0LDSxUzVsqKwQa5er9NS8qpzgLAVTxsiP1miSl//WyKIje8Uc3Rzf4snY7
NeJP2xCsbpwWPTsFOjoWNJgHsRB3aD+tV6GPzmxsGgj6IuKvjtUWd7GdrIivXc7h
AI8pbFXq+8MO4V7U/6k6SI3VwmU2gQAmTjAkbHb0QLoXLJTfIVm/ssG/q0TM0dEe
dqcND9ZhEy2+iZvtyelMWlOqTN/XJsv3cVOYR5oNhkYT/U4j+qVOC7seZjMfTzm5
J33w4Zf9kqvjF+OPimleY1xzJ+EtiwwP5XcM8rc7ZtfCD4h7juVMljaQx7d3Mjx4
M9XBX3EBFvld1kzKvNq63ZL+xY+K4mUQOxuN3GHwglMj4IjoAcNISazMpguiFbKv
QxGymQ1fmAVGmBUbWyUaqkrOb4nn/OmVS0fD8yxV9UzgLhQSn/vdmEpmhjWf+LDo
cTzaGH+ExY376YnE1A98PKsQtRoOzXPYdxunoR+zBGZomkdLeCABVen+m7RizKEn
l6z8jYuaS9pvtaLSbrfZTegJ32vnL+OtiSq6l5J+thbVnShWOl2Op+vfXtdYxf+7
MRldri1/kSbxznNxnu9nuihccou9FhoFzNYvBv+BbCPockhBbhRGQKmpu0he5RKK
YcZ7Ax7X/QDc30amW2jrr408XHe3HWdS4nVTeL43hFuaitibheGnX42+HMI6CkGK
8TSLG0G47GVfzmZi5Vg/XTARSAhZAF1I/kjlEsv+XuvFXAV2SURUOEGDEQ2j9BtS
do4QI2T/tXEBeSsRlrFwubOPANfUQS3MdltBUUXopDQMbdyEExtzIRNLiYfqct3/
mCG8qbjm//0ancEoq9DE0vsRlQX3gZQvNZwzjMx0shYEMe84ypipjedgYYnSdw/W
XEzmEwTcQOm84cq8Zsvb5IYJO7xPCTtPE2wWquJAfRqcSBt4rPbfFvW35QMWESba
PAnMnmmguMNRTWd/otajUyCvIAwJYVVgnlQZGxSNQQeKZ8WKSpXEGtIM40p/nJ1O
qgfgMDgKvSNahG93LvuTb40UlTDShM9o5+A80RACkBRKI+Qi9PwEB1g+D+ea/MDS
J1RK4IS5wgW7n6CTZbNM2m56PwIEhmRzPhcJSBoxOvcWFvQKl5+jTN4Wdyd7bZ+r
GjGExxuL2h4Lhzlaur9PfUxWTa4cbTlaFubJ6PS5ctcHsvlHOGVbohMKQq/50K4K
RTJLFb3AROfHS/2ZI4F7WfWPoNcbguCCOZaojx2Pbihg+cm1c1VKsTm2AG0bSOua
roWOZ/veAUux/try0Ol5FXXzmnd7HOwSjy2BJiT3sWHi0Uk4SSZfvgKBNUFe23aT
eE2yynXR6hJk9hCHsaHqHl6IUD95sKQTh7tfWjxYkkIdpp+QgtBHdm9XyjmcOcfE
Np/RtPtOAhw6VS4PJZQpnQGT5LNrxe+3xxRmkkh0sg+/MWLPHR4129nskQ+wp+aB
jTOb1VXRspHHNOb2vtDsLsXyD3Ab2xz1EsSjJR7o/0QNkIgVaDZHPrT5pOiNu/2R
QZn48+TKKzHyMFCQ6HrCy0y9tBzARYA1XlbhqPz9XU11eqEU2055D0cjsl84PS2V
rI26WrPRpl4bTLRoa6MG88o0CYdUqc9cbQCDSRtB0jAi6jtNrLjb7ZGA4DYVILm6
LhctB5DEGOJN+KvyPa/5OVYAP3mxnnM+CrTL6KWM/AkwGG0r6vfx07rFTxlIZAfs
nk0Q84Aa/0o2JVIWkKmG+UYtggvkKVpqf5VIoYgentLBDPzd37s2lWfHC7k4YdHv
wynMdpc2lEdHXnat6ZQJmQKRQ7rpGD/NYq7OJe4e/kIPRoPV9iHtbt4ssfRsj7Ga
Vk3ES8AbgCFDyeX2VEO71zYeVxT9/tHso1J6YGje8R5bQpS4w7EpMdiDAMUL1eft
z8SbQw4qWneyThSg1200O7KW93+QBYVbKlGvtrXeFp/HyHIddfF5LPwR9/7CrPWB
GV6+AAMGDbDOuIrNxCceNYrV+3HT2De0yoYOyglbl/sJJi6hkfx8vb6n28dAtcQc
UvrXou/62YECFKscXhK30uzQLOlfiuq94h2gBcjF86mjoNCq1JW69/t5gEzeAeob
tB0RMLrAJP6Pilr55QUUngR/J0sgPLY7KSc3WMKyMQWfVrwqXmC9KC2hC8kzwHCV
/UYPvlIXc4JYKKo/nYEi3SaRrBrypzTPu4dUjJVT7AsYyAE7//aI+rr4HqSkESBB
vLDiGKVSdGcaQ9zX/kq206bgZFtWRd449C7Q96PWIm7baLv8FjINzHMVYnvXS57a
6QXcBQvccYKQ9y2PQyE8WkAN9XT3Y3ISnOHu5XeIC/4Xhu7Q79EHiDZjvctJOurl
2cAjVAl2gWXPQmWILeRgNV4VYOAzcPRZQ7zgJigFLzd9ztslmeG1PEV+RJ/m2Zn3
BdiWqosDMmrEWWwUlBCpzAEcTsDop+nUhAyva/rz0BaVzOJMP/5SH+NJbmO8W3NJ
75kydQe6QU1agWhA9NHyFWGLUR/cil73o4t4BcRsQoA7exdn7Yd5zQ9KqxB/oav4
5CmXxUGX9wgZFf5WOeFaGI+BF2VlnBB4rNzBSa/cdo5lQU5OTX4vpo1z1DRGJvVJ
AylOH6Wc6UNH8aSNTpF/ojHyP8qtDvOeVZugaTUXNGgCQXOukske33e8YFxsFeNj
t+gWXnaIrd1G/eahQ9coXUR3hDBJndxLrH7Djrao9znMCDwYHPit6MPqxcCtTh0R
tK4V5MWrFLsIU11qWXNCEov9qXWChrbV2FO4kgz287K1au6olA74DKlHdPt8mKdv
raWA/2CuJhQzsCcP85MpSrVQTldSyTEZEdKdzxhrGLYQ2xe9L5uTrHptgK6w1kSZ
hGUlg+hkNEjnYCCpcXOkvSaZZo5PyRfUqZXKB/2y4zg6j9NaWOvenTvuYXKFF5IZ
MgyyEr+ZGkrBud/Ghex4pYvrPjnFWipeDQs6rjLY/a/raMCZ7b7RlMGyd7/auhZn
J5IqyDcRl6TN9WuNE6lQr7XUG4pkLD50ClJq1+9kaMIsBYrXZrBZ4JIqSfYKH+F+
9qFhQ4S33w+qfD2DtEV4ovlmkbFXly90BhNGffZSxLYD0WabYeanlSav0uNEsTW2
AXf/lQ72bzp+/sPOw/smPLEIzTeThBanOSSaGixvU6U0LkOlbqqEuRyxsJbjDIGk
N3YxeuZ0NmsTxDqvU3ss9e/Rs+DkTbmjTlpOtzLvoa4uueqrvCJskvedQAvBoNiV
A3lNgYUt6xPchJDqE/U8tdlo2qPI1GRAJd3S6aL5Hv790C//+EclXM4ImdbUk6AM
KXZ5e7WYvVvba9JsaeOpGkI2wrcbKbYuvIE9QalK8xVethDEZZeLQwuzuLHZI3Xu
UUm5H6d/mmHnJV74ilxr0cG7JgbeSgiERKOXYZ96sUY2gSBJWjkIp80vSuOh68FQ
QYsBU4fUXXEhEa51odatvkLKmlO6U0iwaMLHa6yHMHwdD113wI3eIqy2b+wlqSQM
CGC2jlMmxQVHTxY4rVdKb03HUGvv0saRfvrEmIBiXkHPlrN2D+avvmFXFGg3RyRf
vHvl6qJ8zy3xR0jjfxQQ4PzBxTqcGtR/buI/b1Z4o3hFkOQfavX5210783V1tsZU
XidfUy3PBC3WFTyg4PGc9bAmJLDWs7qMnPWVq3L9GOOof2Oykxv8kOwPQRYuOCn1
50ERWrzsj1nV9/bmXmu1140OMuvA0eVERHhYThdW0AyeoHE2jaLoDjfxK7rY1foF
C7fzHLsArtVxiOS4gNGs30y5LYkfs7A/ROFId3u6FS1PsYnby82Ggr26UJfYB2DL
Y1ShN/oJlEyelfU6NMwOd6aPJ7Em+rXNOsPuRN83aGaqQz9gO94YYLMXvJkiadxI
LFZsXLN6JvZg6iSu/n8asp2IFDU1usxnU3x/Wzcay2nBz7h92qke5opsfyATjJ+J
0AbFiNaJYb6j7u80wvD7jEUamqHKwz3zBmjwTvdcvlCB4qWMeDh45OYfDudiQSDN
E5PlDc1P0MZMBymzp+744tXbxbz/FI4sghXrwpDhwZI8HJ/GbpIkDNmqKrJ0lMMo
Kjr+XOwKdYfMXJ9FuyPmOP+Yhf9IBaNA+ykgW/pfWtqkZoGpneEO7WDKtemudEZu
1e6u9HB/O/oCyhmlXUUtiLLC6emZ4jH8a4SFkICOdwGD7BQ0dWbjGVGKBn7rQO51
gCWlhHCK2PFH+X/3KlYvWQJH8Agk8IBe18tBJ26REXo8MAW7CwjSbekWJn6o7qb2
sMA0HsdCcqxsdfF+OzROilk53eAWAI1Szqm8ZHq6/y3H5GXz206ZPKoQwKgVAWTV
igLkeSKlcPyOhSC3Fku0BRGGq8UejDmBLcawCdPfWrzUPqkWf8fZNPVjW79N/xQj
17wyzJgHBjDdp6O8pm4PZoXPTURjbm8FlCFKcwzqLxaiCGO4eyHE6w+7D7+UPDCJ
TqjRhbJ3fD2fj/K0GnnC1R2iDaqGwSSD9OI4lW/aAe4z/sTQeZvs+vpBlo/OR2UU
AeV2/U2RnLC9jRHNhXGUW3G572DUfST8T1s8lM5dNtqx/chCRlA8LFBWmzTPFshr
iiVAzTVpo24OE+6IaRFRTtzY1p8sDPxoKN4DUNC3HgDy6TK58m/kiDBTbvPjQClb
cazUt8tB0Gif88Hta50iR3E/P61EJ+YJLwJM67pkc3e+W524t/QOPgqg7KfDsVol
hJ0QWknSjPB2TLicpxYPntap0JwLHSLlVotBYmPb+rJ4Ogk/3hg+RC7Xik22HWFw
VMsykNaLhm9kil0P3IwWStsvcaKa/O39L/+AtyxpnTUF9zk4/sFRATP3ysEOohVr
p/ZgHRbLkruDXSEoQE8GPCJbptSAXtnc40WvjU6sTZf1wC1lLKWPY8b3UM6TpHuV
E5VkSraaERzCCE92/TD+L72OKw6aljjMBXu99Bw6OB+YeiVaSIDxl2bZrs1Qswyo
eYe49EBLGVzlRflEZ8Jtqe3GR04iy4hFmcPS9iOVejTUVgG+dQIRGvwG9o/CMDDw
k6r0hO9CvG60Q4WaiNz2AnJpdZFHYVhiu+IX0oCyZ1c8ZDG9tBoh0OhPMX3l0N50
WOYdR5aRhLk36c09Ss66pvG9BlAclH9G4MP7gelkMaquCJOUebOC2Gk5sV5gxLWz
0cmoUN9MyGRgQ48khuuzmZBEX2MgOIuae4OqVVzOGvpDGYaExGbhlx4EkxAzKb+M
zk923/yZW7K0S0R1BWM0TecMqUfNSzPosVCogPXdSH3q1hii+jRnWa943ocyAg8c
0thVdTLGFxoryN2Xl/NQi2CXfwHyYxxhhoR4VL7QuxzX+TQWiXiDP2coJ4S72tsT
afuIUbftFCixeyHhcPGPSMcWe8/DX+qAGiyxdAjtUHlvOq5dgIvUvmdtHF1ON0HF
8/1cawRUhTCX5/ClZ0S2kEnW1WbiqxCnmIPIarrMLAabEUJrJ9+CzIVbpkhRHhby
9qFivBdCJNjaRHTHz2/jkBa+RHgVJYlv0VbYS2xePuKSr2B00sLqmXfiHV0v0fBl
uNLXENtf3/nXXa5054GizHsgKYoo2tTMa6IupPDoRJwK14kg01HDjcI7goYqbOI2
oPHfqVj1ct9NJz8yj++UBNbuLGMY1s/5VL6KOaJ7n6miLvLPMvibTBkkVpYAdS0m
+Dg4eswi25/L5TK8TI4DzANRFE2Sc+XWjDPg5AsgpRp0gYH1njaFskcBRPMIcDLI
qgmUMIfWfCG2cp3u07Djrc+VaQX1M6cX1ix42wt4eR2vyuJn/Hk4CB1eXquFrYOv
y2Z6K4/ZCh58ta+7o3zHwZgFo8LUFoyJ3TikCI79409TL6rVPnq22P/8khTCON8A
je9MgVxCl4JrKRYxU0EqTrkvGfsTtW/3F0qjINJ5NNbcPi0H/WX/VljmF7NrX+4t
UsGWuPqUjfNc5De3DvOCxYrHose8Hp1o0nlNoIRH7wiBQIHISI7cyawCp90t1AKV
86PQJ+SEA4icOQ391OIJxBBs4ks4bEAYxnGnVTES1n5/bRoA5JL/sd/SpsJgV5+6
yhPiorXhrxmEPUgjgS0muFoMxtueY5iPQrSbMvlvh2cF3o6leDCIaRHnfs/KqGPX
NfuO7JJ5aBJdrhKZQTiXML3WhewIM0zP0NcX1Mi90tK3i9c8U1mJjyK3YoNYUckN
yiiY8UM7d2SN78LiBDd2fscjcnyIlagi7kOUCGG/zwx03wMR7lyjTkUluk0RYxs3
+4+6czIWLe01mi9Bg8LmA6pkLbW8HNE55ajuLff88V6gFL8sc3S9PeUK5zuNp7i5
FaXZ3JJbep40r3WiGszRxZHju3h+UxAqqPzUqcs65ZaIy9N6GsAaiToB1bI1gnPY
ZUz/12IhrJva+tJw03ocGqAvkkEH4Fd6TFcFqAWj+55Seosz55V2wwtXQrhCMneu
L2lTMPsrogUVdg4a8ypfXlTIYm5DT13yl8lL6FsKoKfhCy0e5xlaXL41o/iIdekL
xLjcqTL9mMzglT/9MVaO0X72sU/UrXheBUTMdxgWl8l5m1cI17o1ci0DSqhW+UZt
+7P62DCk511D2Kkl8S4annAzUdS8cdOLNImWmOGnO3M0Fb78jXTuORa/OyiPA7k/
eTKQC2gW1UnofWE4pzLxmowehGX8UwyoOu5NMW+pc3LpoMIz3By+dO1leEAlN+Mj
yckBSisTDzVux/hiHjD+EOT6G5/fyqgj74dAKrTZ4YNjulQ6x8iGt+a1TLOON8Xj
e2sLKTUc0tGmPvh3YxcVfWV+r9h/I0wk8/+zWmQYGTyGICVFNXBWye59nGm5/KsY
wGgdJhJYzfzEXhV6HdXGo2YBjfbXZMSti64cC6J6u8kNdvnusgprTAurdiY69XnR
W3cPIJ/26P7pi+cRzLk6ou02ynvCI/0CG+pd5pusLAgMtuLPjBALt8B1UYreuXE2
8q+Q7gT5si5sW5OQiKj9Sk5y6yUsy6AOS+6geUKNejznsjnZhacf1QAyGN+TbPf0
newVtTOEP03yIxj6oomUwgom3z2JD1R/Whlub3aI/KmO9Pw9gr5zJOQ8YOop4qBN
rnztRSvySaO9XLDu9qx8Kbdy+KIVlRZDCcgIAbTY2mt66aownFKhMoRxcHDpwkXM
w2qYmVyhiSrcFpT4jHDNRuJSmQrQ7pyXQF5KS/4WmH1xMZTmpydhGWeWAoEjzdF6
Z6yn47ntYeGi2SEzb1gdVDqeZf67h0VCNrDOEZmztYWKSqNGSS31oY9Wxfn90ZBK
wGOA7/iZGvzSalcXITTU2jAZW5fJmWJ4w7RZUGz/hJIZtCQszA7jxJDLLB/o4tua
LYxDsa5Gnh1X9ps/haZVFeKiOIREN4BE+TYoW8n/p4Y6gitjt3LFcwXRqQQ+iOVL
1tLtyU8VM9JJ/M6MAP5cFQcWZsNq2Tc8Zs8KKk8EJsZsTfn5XYvWGFhiTEkydYhW
Ocotx36dDrQidAlYXfowWT69dQvWu7zg7xZ8eqeAVSUONq1ZXoV0VmBWIWS8zw4C
my50k0nfD1E5A3mT8wyH8C8KDVAcrcfZtFrOJSDGFc78hzjZ4JG+djPMYv9O6sr/
LGgQuMQLvH08zLF4KbbwbVQnISu4L3ckD1dZ2sNRb2LWISbcStRf1vZmdByO/MDG
rqHcJU2A/OrBbZ3Jl+OqDIyDFdXx7bDIRnC7XJ7+Pb8zoUehCeLUtX0YF7HO5sXO
vgnR+u92rgRQQa6D18wlRLtP2FWJ0+CKzgJO+foYhQYD2BWv1CRwwCIHBVCDJ4Xr
AaE8TxwNGK6AwMhytMcdAtZATlaJmjjN+xujTPVCxcmSGe7oPp0nzYMOD3Z3uzH9
C9QbdKqLCffSzp33EUh1MFvsG/z1ZJw1Bb9BRF77DoewlhGsWK4nRGP+rKW2azLv
ezz4L3YFHDLJc9IeSG8WDusfUTprns66UTa7unhWTCYGWML+vtaXhfiwAg7xz3lE
Ho859eg8OFd3QcF8c/eZwiNUf4Ee9b8jcyZHhsIPMrl/iS8tQmIbpwhATpjjiFpY
jBzs4Cmf6BdQUcSs3pVC5apXxibagDTJz9Sga1SVqZYrJAJb4busKq0anVWxFo9J
j//BhST1mHlNYrvLwqcMRigTrP0BcOaS/BDT2y5p0iCTF8fCIcqgl/10+uqLn7ec
wHrU1sNFWStDoE6c/KUBLPX4GdrTxaxEtOgTKxjVc6nFbI2CKGQV0YlBbmKT2MA5
hmDRlQy0L0PkQpJ50aD8DEhskjcP5Y8POErGLk3Fd/INfi0huO9kYrURApzDvZcj
Z9cR1ONmLWN+Z1jDeiLyQAZSIpsrOQGQwS1I47GSGbRYCe5zTJf7+1HVuUc5g5bf
8sOcki8NOKBLlnG0uHAhwCUQeJY2fLLAJZ2n9DqmaycpWUbaTe36EdkwBx310qBz
6wyIlz6ZYT0zKWbW0DhcR8i07nYmKbwqz93AWa/tAxbmVegMR3UOgyqHQjp25VX2
6ttmyp0upp8FFraWcfJCeOUL8SVZyy7cP29NGhyBBVI76G/NPCq5I0A9TNBepocn
s4n6OSShf78A0m5WapfwgW+3HZe7z/zaAG5w/0bug+qX/HDfBEv/3PGHtk2T0Zej
qIjbABH5f/3M+stZtXD85cVsbR34MeBahGC0aXio1ye88zBx3vpnNdlRIhMZbvup
HcTlHrYBcpx/LTBD6wx5TpQto8BLAG/V+82d+XvUEzZx/0DutpK61cfSlS/D4kFD
W8Oz1nu+ee5DVbsdYa4VJOQeqB0VSHIAxkObZ1Qsl1bnxFNEHudCfEzYoaMc1fT5
k82CKJISONIZ52enEN770B1mZrIeSth/fuw+40gxocwYBjvlAlGOH3lz81jzG1O7
xr8mHfrYmay9bSbYAByEw8HAUU0i9VrHn36VimRIYufkmTLiR0dCGvRotLiKiSwu
GUI5TXKIOMgvkxGepZheUVp+fqjHwCK/XNYBWMl6G+t8csT1BnbAJB2I0bHfRyJ5
onxJ2Ez5QmRrVX5j3BLMc7DxhVTy/r4vnKcakbbp7lul4pehkxf2HU0fmWx7TtWG
Rit2TBejePXOvfSbJGIh4qNNXjlbdu1l8GMYUB1epEEWA15iDFK3SA2YhU8oW2+R
d1bffZnWJelMKzXal+mZtUeN5jtlAUa2/BIyx6HNI+gUHQXuTYaZhZYG51T0aLZj
4bcQ3mTVcndzDfHWsRE0xfRaoQl6SkXY+tCSRfo1ucupcgVm3Tx0yed58TCnlviJ
OTEXIuKx8/2T3UWhVxZEHCK+WwD1fC/TSrCoWJ0ZtkJnls8y8wcpwTwsojyp1Zyw
rq4175Q/MO71hm1XNUxBCT9eTHPdARcNca2eJz8ybHysKm/5W/zZ0oWTKhUFJyip
G0h62w/ml6QxK1BLDBudDsChOYv8isXKCTZBRL5aoi3QA4Oyyb4uX2rZnBSqBrQJ
H4jDqVZkiE0gPgcilZjwzooY9WOpsjfSsGsFWZPlNsdp+xFTLxkGTpVCH09lcef0
UJ4llncujb6TkxZ5spMrjbVmvdZA9MRc3PEWQ5m+XCGMj2B3cTOXKNrxlKjPyKwz
eaVY+iGJiz/gfpUHhxu63Izsg9AFuS39L4+rMYX2knbWOLQWfIHdd4c0DjoUPhnS
EFaAXnPr2QsQFieS0oM1xoe/qF1cmJtQDTgUhKcGUBVXWMVkabCNfKhP8ScHd4b7
cbJ37BbQwXZhrP0LWksXv8GwmNjIsBghUGkV8vja2vA1inNV6JynvfJDLK9JTIhM
kRaZoWaqSnY1cATpbQZLRorSgO9CpCKoj+hFWxKhYAkH90J+PbJJY2x5QCyIIw+8
ZzGaJfBu305CxPHnRx95QwKw3Bt76cl3iWyGEPzkheJ0eB6iroufo8+yV0mbvsOc
8rLiHJf64CVxCUo1g/EoIYlRHJZLJNSY8+7BokMOhXue50Z3906kW3db5P6q53Am
+8qyCJap0X1znL2zcw3EljrS7kDfTflla7ZtkzRAAlzNoXeESiA2t78KCkCxZhka
zv+PycGeh+46AShlWcxJYMONZL2hF4c7xHbX4eOlDQDOEcbhAprLuMphHfCuTrVT
ABazPzyTeJdPcqwY4t5dHEd9PESMXmN2s8xJqF4mGM17YnnmIvrLb/rwsrxPV4f7
xqSFS97ftwB0xQiX6AmwiclwfRkstp8nG/8JY/xP4txpyGkQFHTv5ftwNA+7kX0b
G6aYFYPOt0KukvT7zSw77DIUikhw1rWDlB5Cn5PX1NkJxINMMxLiyAJSD9sRDQ9L
9a/HLKPOYJCpHIGb5ftMybQTG6N9J6X7GhnNxjGNpUDEo6+YQho1cm0szRKufj88
vEnmr6QQQ/lXLqYJabVooSnC36Psxbtva74vI0LJK9LF4mIdCK/rZRryreftmecs
+KzqvT92kc5/X0jirVDsiKoplo7CRmNH8QEGMvkgv4C3+wxKrkh3D/u01UzXXdBK
x4NEvZyddo+3kHJUUokXGqP+0LU6GhMiYUv5x8/ut6W+M+N2rGS9vja4ogTfbw0W
iBG/Lwo5mFhdaPCs5tpq9XuuOadbXSK+Tfm9idY0c81pvERAJn+eKfvkECfqlP8l
OEGQBrkLpZ+LE8jEc4c0ArC+5Z8FhVibNzlXJPQQERm54biZrw3oyu3DEArU4WUl
K1ko0wgfBaxuF1xymph7oow4XOpf+eK5cQ32AVk37HLA5hQfZSkcpkmDCgOIagDJ
6PwnADzsm+nKePf1ciCpx58c+DCKu1CJ/cy6f/RVaGb9g72pHRK72T4jmb57/xG2
0eDJ9VCd6AkGRcy1eRzElFh5hyRjynYnFm0KMyaHgtGSsiglDiLD3p6qCFSJyIU/
O3tHWXPnD2JpgHdMftVjYyxoLuBNWFEX3zt4ziAFJzm8iKaDD07r9ebCaFZhiZV9
5cMfQPiEyVCS5MzYi+yG5Ir3J2n+nVv/dhRTT3M4zdYUR9cJ8YK8gT7dQ4quuh6I
tVtmsiV+KEsIr/D20xaJFjPlmj2Ns8L41L4nN+TRvcIR2kg9qD0bWS7TNAQIXmCs
YWx47STilCaRKkLuleMb9ZPwATCjeAbLQ2a3lJzONEGzOu64PwHTUIvfoSsnKcfj
kiEerLJTBw3TPSLM/8Wc6Of2b/mNlXh/CC8ohEzhDn7RAqFeQUPzJHi4LhGt8uAe
Lqadz+otCHL9sa+RYmeqKmFCRNKV+c23/6Atygx2srBuQAjx1FUD1yj2QTK+a0CA
NYkImrKXX7VGeHJGfqYk3xPVqTON3PzzlP8v9giKpzCZW5jw72LK/j6pFCJELdNn
OQboa1eZDrgZUTnhXXxFB6Q66EvwpMgNb+a7JgDJgJtthBUr83wom6gyD/Gt8/9g
wR17vGdS0QH2S/qOXzQZW7i0HD6lQQwyNQWW9XSU5Eyv3x/Dtdodwl2rwILPpQ+A
fPQSWsqAUyHhPlh8FUpzj5Z9e4VW+om6gJ5XZK3qB7WEvY1LISq35x/Y9rMdJQER
9BEHw94wNrnkUUL+CsJyeobYYLYJmLyP71s1pmt/hsl4Fg9RlIgUUYhnEe7c8UEs
chIEtWhfOKLpD7UTtaAxa6qq2O0jjPvuwmt8ZhOgpFtImb8oVdRQpg/7/Hqp7pb0
o2bw4F9QT7qBiHQ1935MLcPryttkNgw1Ugx1mvAzxpZWTe6/7QnEU/9t2Mh9fKg4
0RTt1RAmcW7yha28qwOLtGfO9p2Cy+qKW79wIENUuDpoZMrUqy+0DUZeE2HlJ94k
V2mvZp/5X6kg0tITSivA/J80R6Sebe0QLEOzt5cEb8GJvo0+hv+saPnVmqxAUf1r
UG6l4hbyMkkGNw+snoFGuVFyMpotwcgFXFHVGz4Q9JcWuNLRpi9bTuYuBO4aehLm
icgDVGtX1C7Ym8MRd3YqwQCKjCCpu95Wntuswc73ndPZw3dn7teelZT9hLMAq2JC
PNNE4c0KZirmOzTVfHeaGFBSpXDP73pF/QKaj/C3FnemXeJLlA0U1P6+JAk+yd9T
akddEvFa0V/3NBQjdNfzsmvtLq1o9Qq8KmprS1yB5GhetedqFVhaeeWEsiKahngZ
n5cPQGrF6i7ZtR1aqb7qicqlbCLuiFqGXBQCNBe27W+bRLZwPmC5isLnE7m7416C
BGuvu1jv4R3Kb+Zn4t6+rYKU/Rdldwj3r1RnW7JzNntrkWNj3pusmeUf+G8I6Eb4
PKTmqUMAYGi06AWa2FN+EO9xmcBQPR0rZRzt5O33KqH9wQL/cGRkYADG4pNd6EP4
RrkJh2Qhj1ukOoXi4wqdObSRxGjolhjKsrRaJ5lyakXEBhOaNR4M11VvJAMeksxv
0IHhvJMBaDRiBL30Svs0QNMFoY8WGqUfhT/B+UhnkS8N0K9pJnkAVd8MK/0/aNZE
2Jb9JKLNL4DXeI5zR3ngUr79EJ8CR/RmuH49h0sEdTVv0J0v221vEGzhk/lyYbFe
UQXJ0ZS3jY5d9lW+LAIkR4BGUt4hNSc+vSfxEKY/Ux0lfdpEqgkir5YuYlSFd5S6
TEKaKHzc9+nJUX+qRdu3TYuV93OdbDl/HBZL5MT5RucHf2UJMGROxq992A/RHVKO
xPNl9oci7vaGvmmCB93nwlt+iCGLZZntPsaVdvJ1U63hGHALHrzhljuR/8TnSjyU
sqwJORk5fRzMNxiVqC1SZtz/55WfQ0QUdmnHVxnh9Yw6ebV6iA+8lSZftIIdeJVM
YCqFOXwN851mJlstdkythNqBVEAXKYIqbT9EFSfv4UHkgUJXfZW/gSOYSNFOasba
OeNMcG+qiWUjLgzVerwS7Zje2eChbszFbgRUx+tf4oYL8CYCLFh1LhfSUwvbcm2j
BOVpFOB328RC8fA9z07BGGfANFz542PXwhPgLjZoLqmKwVz3xj+6AYHhrNRwuJ4O
hIejvUQLy9vAtnP5o3GjYuIp/vl6wJat6vNTvADZkHMs9iU/x+x/J1U8o6naYltM
rV2BTIlOJqYUhv0dB5XnG4ue9rPZrk9+2gJPTrqgqbDCv8vheytup4yr0slsUrgs
eWHy7KNpxoJlFygqwuVabU3+1Me5aF83lKJLEmJzeL303rWWDJPsY5IO1Nkb5xC6
ub6uQ/Ipo30LBYu9P1kSTNSCo3iqb+WwNLJO4VRgNZi3G8MWLWCdMnmfCyX6igrt
vBHqbqGxpC7M1u+PU8ou8fqWWTxrKLmnqWUWaeIG73v9zlbhcB9gALZDUxUW/2Da
LbUglM4KqGSGYPyj3lic6AsNV81+/zIAMFSBdv884T2qh2kkzDWgAokC7g4zses2
MKbnZzQdaSZIwF+J3m8o4mEdMMremnWE6Q+7gN6oXboY8zcEX0F141h/wIhds50A
+LE5HqKaF46fZsntqLbSZYSerEWniHgL0S6bJYVy3gsq2Y6B9zT4mbojmonW6yPU
jNwTaren84fye0AWocEhx8PiLzOB0jY4LSJ1cnUHxyM/FI3Mcy49q+z8U4egZ4DB
R7vckE/xZdPQZ5+boF3aZr/TScGw4BmYrTyvPAnHbyHWmXzzbzHaZlEAfur6dLHM
RHGgv73BaQo6teIts6CbfTK6c5KeI2jvn2Ns3fPW2AmNAlwtw1cSoirWm+xq+VJB
E6uuvR/a0BL/rxi853NlFUsnsD/5R68Vp5g6UdmZR9YopTkt64DAEMwN0MpAkuGf
pL6cYKqZf4Kp8pTISVzhKOCOq/1vwHOwfB/XYQUJwq7AJdZYcq3ltlOETebgMMUf
7OefWDXENVZbE4l2Du/4/BwLbuU8CyxAx78eSux3kvXtgN07LXyRj9WfOfin7M43
Qorc9nD9401b1A740L4/T0Q1qX2hE/RKzlMuStT63Gz8UYpdv3kZwMDf3hxNnJor
gactJEXETSDZxntuYGp2/dRs7DA0o9yp7wx+V/CulFiJwpg5kKNwtZZwyQ5mnsV8
w3UPLiLTJ6G75chMOi5SXasEr4btBTpxAJoylS3fpCA1j0aAXosFyet7qUxekQPa
P+9XVYSP6tcvInTmKarFuuff19RHjtMJZ1VqD5YPVLnJPsSY7gAJRqisscuNPV2P
12iDDNrTZqsbUgeULa615dHLyyU0BO6un8K9eCJknztGkT9jFUjZnKhwr+30YBhP
fm7YktvhH28TTdhLipMOvbbFD8F5s3goOky+Ih9Em0jvRQZje31Lh01FqXaQ2pVr
tfzhJsVl6B+hob8iAmShXq5VNu65pLj8Am1fssYtPH1i2OzQeLb0d6UVR3DMTWTg
1uAEy6UIKABD7FRiyNadiZVKlVqqm7nqOenOljNXv5OOIYZG+0zxlpwSmsFEO6tQ
8vpobAN5guIyfmgo275giqT0sT3f/QdbpfHArmpI6mwdw4UdUyldBFfqSQ/ywLyg
r3JbDc+qRvObKoD5Eb17zlVCEYyDXk999t7VF1GSR5zz37O8hTbkLuKezKgWaMou
IrRh5OFqos2wZQXZkLAWUT3axE2ooNleaWmiZCpaSMhXZYnN9mRMoGgDIUzsRU6j
umFjrE97F9N4q3ubut4y3DGb9At1u2j3jgdP537pe8KDTTMyYbrD7nktL2uiGYH8
FiL8xsBsV4YIEQzDHZYlMysN31kDbcBVy+umnNsBruciLMLSw7JA1x9il1Oj1IcC
Ep6Mgv/MNshypTc/TdVwItka4rG4MPxP9cFNXzbxNKeB+efmb9QZaIUfoaITxtx1
c4xbbiO6tjHqo5a/BZh9Xxgd8GX9L/AwecGfbIm9lxrIwfw2x4gkQzJxnuOBBfAL
g9OvOjpyrsnkz8Z08+a2mfcnlDzjgVYiQ5WUcjAf72SngRri3UvLx+nMRXWo/j7f
AiCSV07A0QxZh/Gf71vVjAhmGo4S75C6FofxrMVDS/sDOSKkZnkK5AsUAFeHyUND
JAUK+Kf1v/3xx2Xag6YJBL6uTdvBnmUH7EoQCxvuNTaDKzmN5n8IIQQa1QRonBxo
ImVMTYWWuiga1p1SDuRuHz0GjJSOiDT6M1Jw5k12u10yPIPXAWC0HrP+MGmBbnkF
GzgVPv0/SECEBiNgPAUkkOPyPuuVJv2bUlx6xfsJZjnhE/RHCEt6PHNjplEmGcrY
SKTZXiDaH3HjZX/wR4jjqr7EdNSMC1tinn7rB/yH13fJN2tJSk4qdnTM3aXr/D+g
zDQesWhnANYwjJck0L77rBTDt/htuoft2d+Y+0hyiUAi9ofw+zzAae2O2Toxvb+e
kf6OVSgYe1ri6gI8PR9t0sIdMw7vPfVQ0DZCvilkp1/3Axhy8kYKSjQEj5ZhT4VA
MFBkzMGY/UIgUM3kNVhUjvc0yI2FSK4wJZPaN8gSbGgNBtQ2vlKb/a0rHzDjVXWf
q2jot+ru6oQj4Pu8YdZeh17pw3w65TjAaXIyHOmt2UXyegQ93nZFpTI8ujOte7yH
g20mcYomYAh90Hyhw+cL4cbkt7AvWUoi/YS+XNUX8/g5X96rncnnzuHwftN3gFSW
kou64zFd0UuIDzBk8+OXgMRxOBLhN4hUmiozjO0/ng6SVyZpFPMBuliK+BofVZsW
au5gl8z6axil0Cie/QUhjAbC55i2WmYVSjw+f3+dwd+vI9f/FcJ82Te70u1vCsnU
TxXyF4ELfdGp4snOnK/v29xQIXLQucBp//y9r+4vxCuykODxiS33HSkj6poZYof9
SIKVH194XBBTwYvdhCUMJ4v2rq+bZMxfry+mEJwLUg9wLTfJnjTpQu5tIcwg1aI9
oguZEuICCvNhlsqsID0BFnaxwCx/ruFk9iywRp+7XleFDx3ziRglma/uoQwAXApP
34wZSM3oOu6cNqegMidSvAPRPzzAZsgD+3Py/j4SDM/SuFA/gRkYc0SPlOM7ODUu
F7DtBI3MmeEBOlKZ18fth+xhHPLKlSC6+OajCpsGZcb5t4pmJ6T3s6NoTGNuCwTN
78oEwVTK2vdBdKBBLEyyOnPKKLxWRrpHr8bUmsT6dDpWw4+sC/in24M+KWHc/AJT
yrThwSsx812JsUeSS9CpORXCOgDuPSCMSjZDiR/Zv9eL/aPi0XHqKKqn9J4jytnH
oYBv5uQfLDHk5oYJXD03UbzQ59AQQPy4l4TIDxl1EPvNnzeTrBslO+V1kxR40js/
w7zku/mwY0zssqb8K4yqjIQ3UBA2x3H3gpZf+Biwh8wtPUt+XogH8tKXEw7No0sG
/nPqK18Z9jzq+5L6S+NH8iZKbCuprR/bTXxbzfiUkTUaWfsSkDYdO1N9K1rjD4Qg
Z8pI8pUlitPqHBzFghZNVqhrXv4ir6ACF0BYHtkm3xnEn2peS8quNuOURUwSXjLi
Ma9CFfxF1tT8FtGIXlQn/sCfm8ykm4Mqkc+syoN+52eSkuOH6kgPIyHNllLJUfXe
PsiEbTbdQu2vvsdyyhVlQmV79+dA6QXZnsM3c/a6lMD0YEwX2D36ZRaI++z6hAfS
+ByYLAwuDq2wYbIdhXdM4/QaxEi1a3sHESUFofdD6OJhsxdCOQngWZQFj79c13k5
hKVz88FLIQl2Ba29ogAWfdinX31tthUm7RDC1zdD9/xw7PrHXa7G5dqE17/+vDda
uWx4SsmM/FScRUE+YnBs8InmLd7/3huA+VGtkpn8iphDPH8SF5mugTEXd3yoznvy
wb+PZZylkWKLe04ZaNAVEr9ANcrDzaeU3t1XKGlLwr8O1Zz2iRSpP9fmsLo4aAag
LX1Ot7w/h1L35xMtL7aoNbiCppFa5xb85mY5MfmZz4/zgVHb1ReJmmUJPhcgUlec
FjkyDr3x35M4DOzImQPwXNRkPJfYqec04ALBptT+OrZHy22IjwY/eo2nxD8EqVD3
i9bLSOUNJ73TJBlz7TZveRZfdPlaDBkQ0R07cxhYx/U1I6kdvJoNOxsiJ4f4dWyn
cwj17YlOEa8gNNnJ5LYr9gqyvqcsA+NR0vVMg+cEp06v5miXW0v4FK5BIqsd2Fih
sjiRcqwrF5SNOIIP9iddj77E7dzSu5AdYkHH/Xph830q9rwVMMN8fbxXWCse5iIW
LlRWaze6Jj5b0tGmWtO8DMePVW4UKE7R9iBYoDsldBJaIW3FiaZmdRJc/Ys+qhqL
LcGBLy5iC0+opHOtG7v3Iy5LCMKRC4DKKZlzL/4HzOqWRdV4YdIC69uwcNngEsHh
3Q97WyJ+zoe/jiCR6JHEropIFQqOdH0dBeinOlxGZ5rCwjfW0bRC1nrWAQQ/2vz2
jbWfTXXaLLsOfcbrrl5V+5mPhTNMpfJPTByNU8Qgvh1I4Dtud7QRrxsnX26qTBeI
MiF7E3W3EeMfAJSKP6kWkWO0y/FPHC8eB+G3sKKpM9X9O5zKr7Qm90kHQFVMQRzp
kyOjv1s/R+UJV10X8pCiM0gf6JXIzoSVMiTBXS+SqQnCr/iEDGccLxnAU9E4cvP5
cUxPDGaC1y3IcRA0m9Hu2sm8wnz2OuZUb3JNGitx52trqycQK+Lovb7PiHVYBH2U
zfnGXEh2aP3Kn0iL27RjMnKM70DoU9E3K6aP1umeudXN7wU4YUj0HBBHC1rEumOu
GX88kpB1JVf5T49Y4dIr0+N8GKDr8+3zBRMFqMSGpCipwe2fpWgSR61ymsw2MSKi
UnyG4kEeVWb1HUVtGXFEcTYKuli9Io6n26m4E+mtXeUGJDiZ8iIfyeNC5qPfeOMq
4n+88NqCItOPrxcH7emRgY12vF3KvUd5YgN4sIyH1Xcp67zcG7yucxYFRLcexo6B
A8u494c5TrdgHvsD8zRQFY5rEN0uv14B+/aiGrVLUqd+IPNGvZLFc7ARxSruCntx
aMx9a9VoJkD0VbLnUzlrXppfkXAgwYJXWFq+G1CMNv6HWbxdolJxaj4VWv+b2IFJ
OpasnoP1yMs4apT/NQtu/ie53RpUhs2lZ0u0nEpAiaRPD3YchirgH7W0cZygLVOb
OIO0fbLg8dSL5YGXWLFVEnsMwnR+ulbOii0tyFH3Ixd8I093DRdTVap8W7uCQp+L
Huka8LSxuWSruO37Y6lGPf9zK1c5TSUMoRedM0IXtFFUkeQfkyoiwXYxDMVmU+zF
qHuV9iK0VPjxTzBYZHNzx/d+/tgBfTpE+PMAyiNvfvLiLKc3nWUChwGIMtUnKzL0
W/VtHm0Twfc69He7SoKhng1v+pigvAhPIAlXK4t1VuiLgDVBhL9N1gaDMBCYKrs1
pQntoEckPyo0CRVxfmIumABLardvM49fX3JbAGbK0dQdCtJfSt7CI5pEhUB/PLso
pW2jHzK/9l+fuz1cSM3lXkMoy65es4iKS3Rr+KH7TgH6lI6dYNjVRPxG8yYe4i4N
ytx5EEUgboXqSFfFwrJQ3YsX/xzqb0h/++Wto8cV95NyQXsOto9GInwhbr8VwvFB
p8JwX8zpWVS10Ltw5oNxI575HKsY4cQqD1Jpxm8UV1xXSPPjgqcOLLQBPTYzwSyB
NmArznwDsZSWKy5OyJ2Yn9ewAklxBIr7NpRqgFiBRtAGrVZ83fI0l4xtehJVN7pF
eQdWKjDpjySCQc0SswtUAI5fA+y3WxrJy1oB6zoICr2/sMA3QR1xnFenRrCdT9hk
HkhoM0a9u6CjAGaDP3XH8KYPE0hqs43QacXGyNuz2vT8tYctQexBnMMFvKEnZS6A
sYXNublPi5J4tv6CYfdgOc5FYjGMeklwXYSdkF/oAz8IZYsnsk4YPo2OS7RNjtpz
lO7KuJYtrJEMCmoseYn5/awHyRfuBV1LVfUlambVqf5eVi8f2/LW148w6nQvZxWI
vXJBGVnrsP+wYy2Gm8wOBjTkYWOK3u77UywJ6bhB3b//j7L7QTRYpkXrymDN2V7A
VtLg57SELKxYdl588vWbOCfwE5IQSuduWcV7r2dRVRV5ZByaNbs3t36XpjAp1Ro5
1xcvOyqKMfO6Kv3+3GMaoFEP1Mjmjz9Aip/i94D77V66P4JdTbEgRk7jYFxpbw6R
ggO2kSGdFfRkJi0R5hcblq7ePW9QSnHbZRguOqeWEa4wpC8PFRtpjkXpA8UwUDzv
mhZP4M/D+mzdVPdd8YOCLYNsGMMTsw4vbqD1G0cawIzKPcVyH3GJ6nIhmdSiUgo+
UC/FTuRQuWRmJqS0VxC9Bobs6Uc8BJ8+5cHUaSfOQCp3RRrwFV/ax8qRtXu7WJT8
jmvZC2f7LLq3VKHq7bxJmojC06FVZPiPjQH+c+82+GLM/cefiPxMkTEyoF7J7Vvb
qLmmm7g9G/Jtmv84io8evZXZBBexxC9xZ0K/XoXviZY/Sw7zyjUoOkCyDCaNnK+p
y/kiwQ0ASaZJ/1G+X63lw4nAtmWeBHrhyxEkMuzTYZTkKeKSQpWCR0adjSUuY4p3
zt3XEmvORQ3S1cv0yQ1mh8AhAM6KeeCcyJUigox1dU3POSJk6yQ/5j+2cO7A+u0l
ZJ11m42YooO7gY1RuVf2J82owgRIHGxTfxIO1EXMslxXgXTAxjt7HicfA6nztcXw
5ERvxuWdg/+01OnxqOIs0VPvgZ1o3AcVeDEnEGr7/3lzvL1gA+ONpKeNrAJKYKMU
R/u3hbTC67twkzSenchPS5NB8kMVpCAoD/W5qU1RIJxulMpv03vBohzdlUMs0eZu
GvIf36hRPgvVYABXQ/7TA3syIUJnEepeEJ68/kxd1ChYeL8POomkjy8BJ3bD08wA
Bmlp0sY/DxENHmxq8nXaTUyshOiafSnBI2xvBEL1pluAJJcy+FN/Jd17eV5ph5YN
n8DdG+CywLixCw/crUw8ElrTsCS6TOeqNGweu3TXycUY6MaA5uuLthuikWj3igLs
vtmO4bgkpWrC58SlxWawz9BQCv262JGkXBIw/Z9HP74TuwPnnaPxiSggbRy6R/Sa
oLKKMD6hxL6RBZraW7x9+eGm1i/9vEsFzYRHoRvT31UhezdSYZuE7+xqZsboXirb
XWfrJPf7Sy7EyZwccQ7KPHJmk2+i5/9t1gxQHpj17bLFY1hIBvkiJ0DWGaioRM8D
4skgn7V4F6bnBgo8zzUVZIoE8Z+Z/rpmGVKqSXIGkIwbNQ47tCgv6GOTQVVFbhAb
jUPHEhklmXD2lCmAGhqDJGWBaNQETKQJSxyd0Buo6dFZxgtqdMg77xTSvDHKjgn0
edRXYBDDMklQTnRS5/sTTtOJNLSXIDwRVHn3HytYY9It0Wseq4FS+OBz5qpTdFbG
MoVRKYfgyy9nzezZ0uUUaRZpQ4treHRVeptggBisgMCgJA/tnVG74Xr3WXl4oPPV
tNQJUTwrI2YkiqcoxPExGU1Nuko9nx+zfrEsEPuIHOvMvVbYwCoHccSHzrrij2gD
+rZWjkrGKdBD394NMzzjbwpHG031uDzJsfvtWrPuEKS1JRUUpDgbIJ3DDIfX1z/A
yo5Nf/G7IZkE16+SJun4CT/LCKAAyxUPOnMF5AKf6jGNwjfl0a9AtSGFowFzqBpW
L3uwsjku2Ku+tZpH9cmHgDaMBXg2H2A9jbaIufnMtxWjNn/NvXYS80iUoAuxM9AY
lVWrWivXuxcXi0FwPqsbE1wKHkJGXl4v/DinQq2htzbOi2TE1yc0mPLn3zeKO8e2
G+/Ms+Ncm13/tHmpxYIbYITYQiJ7+bFDD6yWND7DB5/CVwQb65YVn5n69tKuI+tD
gjZfBzLmU0tdDlViH4o0I7bePPW5GCjUVSin7dLqoqTtTICupWXWi+rSYuCu9DsT
Gm5zFrpt6qwOFSvLw/Mq67ERjYjXAXsyUlsPQhbM6Mc1aWUgp8NGJ7a1yXqUso0w
BdStdFBGntLFltLnQb+LC9Nn9mNua/7dTJb3E+HLk+jxOeT8cXwcR2gQxKT7Sm12
3bzpr/upgN5Fz66w+Qow9mpYVikBXZXN1ykx3C6UvaHsESUWRR7QQSjfj0KF1ht9
caAa1xibTKNxrCAuq/VQ4ugYdFMKNmrbesBxq4Hm9qNdsfjz7RW/SC+NetyrwB3I
w4crXcTbdZnbW+Aka4Cwh71ZFuuhE28Axk11NC2kyKmIwyNFEI7W2UfC5Y49K8jQ
Fz5EBbnBfK4cbtHkVBei3v7VLfAcM5OphUx0JdmG5yI+psKuO20uqmQ1ZgS5chTm
6O5bRPZykb68QrCNMHE4pPW2mIozk7q6VkVZMC0V0Wnt7OFRocuuHGVW6On+mQlZ
c8sJcnhpH71aMywRP4wP5IG6juCfIYNHSW25ezImunJCIOt6rBLk9oXtHtbUM75v
6/BuHFL1EIJ/MyK3JPzyWOe0giJ1JWG0yzaJp54JtqnCy62d+PldkJUj6IejqE+c
/3j5YnKe/i9iPOpEvi+9+6cwESL0mzr/3syZ4UFVNV0eW8ONc44vbIGr74ytAYHz
Ps8yHLjt1axSjKBTJoVez35VU+/H6+uv3oE3MVxSf+2YxIIyBSlvPrDNj8XXZOh3
InR2+SOZjgGsj76NtWJ9/T3vqSmMO9KBAQnh1w4x684XaurS88HJ/YxQIiYV4uF9
1kpCbleaWubgIN6EtkHCI2Zhd+pGP6HZeOd+2OmBdrIiV/4NlhPPYgdl5xvW8GOe
zw4PuDr4eEnHtVzCkEk8iHnbZuBQYqVKNj/yoSFj2kIOr/1rYfw2+jsI/HIwKPmQ
RYsOtwSQHInHFiUCjYPo+cSs+lSP0eCore6jgE+ck4sFGqVOigLX8veQaGgooeV7
5UQFbL2JM1TwWj453dmpf1gLoRy7lA0FRQwbGm3MEj4lIluD4W7wvZqu8/f6Vrqh
5RyTpFpa1KuZhlw4BwydxQUJ7/yurcnBJIRbPX7ed+4EAnxtQvailqPzoIgCFffm
JDBNrUsIBrSLjvzEtrhlvhHFsZScV40Ko1HMxcOUAX8Gv7pjwqkZ3NXV7xLGZjnQ
hDyTjpW8UPTEqmeAteh41JRWsaKMAY6WqbVtFkbwxoVvQXj1qxdsI+yJ0Wbbf8CR
cjAji7/dvH5x9QchSl/n7PHW5bqmw24qaVI0j3OYI92AipNUkVqF7TGtsDLME/0l
SUG63kUJcXplXfcjCsUFW8q/lXEIVen8d0GE4v/SDpd34BwJbg2BS8t0DJFU2I6c
IHxuhFCJuVEZ75bk/DD5ZNxea9ro+dke9j68QQrBCCsEC4hE2f4B9a5IGzntnrMn
6AVPFqgWSC/9upJ4RRGsiTu+5n7NY2KgA1Sfxjdh+TtHO/8145Is0JtGAa8zX6ah
nJNiyYfeCbtmUaAU3b6RpdHdy5tmPmCvMeCmyrZi0jpsP+VKVdFhWYgMFH07tOPL
06jTQPCm9AJF75Rjyu3rm8eLeU9RVLSIMdOvi/9Q011cKWuXzixy8nQefpoZ/gJa
mwPLCuZNGRTbvflj8zF7NI6D+t0+Mumc8uk1cq238MjJS+Z3esZ3hVS4lOlk4eDT
vzxAEvpkSjNuzUmu0cOVSGkzqq0s9xOJ9vM6KWAwNbqJFGlMa7I0GcWLuyew6xio
k0+zzLJ2f/nB73raZN7H5s67gaKRUeWxWw+PdaVvRHDQgiTPDjaTWSOSs3lIev0L
tPA9R8o21AqFYBcB/de2jcP6FOY43b2JOV7wGDfBodSMLp8RdSqojiMNXn6UNJOk
Gw28VnDOnGqZxgUflf/xVkL7h5PwxmUwRBhnNo5I9UJkzJZTXxoEdVanOU+K10nw
aVeaBg96eZ6m5DsKb6Q/KtOrc5SU7pF+Pg2MTYOnROyiEyvUrCON4qI7XY0cFEq+
l1BsbY4bLkB4p+H1enzDOtl9Iow4J2EsFQtfgkV0QQqELPT6t3dtFQsIjSo7aB8l
FmuYi6FYA9t5wQI63jx7+HQoDawN4nwclfgk979N2KOnS0JiVFjEk43+0bmhDdno
+b1T3xGjycH8B1ua2V+OTpCvDN7JzSvhHzJHsbhwlRaRSBzshA9kLPrQDStV7A/f
UHot6AH7j+G0INXuA+3hCS2Z5THTSXd4cCopLywuuUBgw3Nl7+2SZ5u9uqc8eNwq
U6zEIPyZZxU4BYM3lmKce+U+MFDyAoVcV9PWIqUBUNDBSLE7T84JFrsasZ9DmgZe
cpBEcQF5UsL1YzcXahcpShR8vVuSDo9cw8tmZfjPoCV2rcLpvlNTEScOAbs5TIRA
1JikFaxdFEdK7daIHB8GKCRINDbm9vZb07m3UF2H7FcVVf4DGP3NqyJVeyojOVUR
Ssn0k3wgXdsfKl57M7m3scsfP/5UENENN14eamC3hCpWqwNeitSTLMmvi17axo++
MFczoZwzT2q4gf7mB0ilTDgLTWpMetJwNaPaycqY5wJTJTbHuI+Ob0YxpVv6/unD
bM6fk4MzIb8NnN5J14wFAsxMbTsy90VaSwlbgnEyXct7Zeq/LzOLXWKMyGH9TPpx
3UYKCac1urvpI3moKyZVUn4MZt6a06ErNjR1IUCSljWbwmG6Aars+mUvuKrOIB+p
j6eLb8Dngeuq80qLTjS5TEI1yOny2hqVqEKV0igqlC8G2Fb2yZU7DaqV56xHsjwL
Q4MuyqFhAnEivKhZgKuo+7zz1JlJnQLEFBk4+UJV6GZbr5VnPBFrh6WDgvoyQLtG
BmsGYvYudgsIEz1JV2nwN9Cgl8Ox7tmlqHIMFs/1n9wxrf0tWMlocnyWLdanavN+
6YHmb9iBLw4YlFA5wspshyEFtkDFtU+XzV+OkYlN5Rwms3EzBx7tAmFGcLon0HZn
xic9HBaOOB+kfSpU5KmMCtvxABFq3rlTGjiR3EKDAwsfXSloLWGlMJic5zqpHpso
S3PO717iPsEpjglAhvjqdOkPb4d6jA25dVJnn3fzVK126aKKnO3ssdM9C0IOIRbi
qAdUECk5Ur2pHD+dpRii8dAx2/J7OmyhPqEZkeZuJgQrJCuQYZmgNO64cMCq8KLb
3qBlpYdi5CEUbHQtcxlvvc8KaVY9DEVd96/4fKjuZ054kz3Ff+/T+zOG0Hnkvu77
Tf43xB1by3iWS83LE8q9KulBpD+y5J5+6ZfOioFklbE2/zPzHgKhpxU3rZ30v/+7
3in6Mv5GIqkYSiTvk6I2MtwEPKHDM8R6P2vueXh8EeqF7pc+O52ApPgUJoicFYpc
J4FBHnRWq1FUhipOphKaap2wVbbE31R/jrh3fjChSYU99Q8YguLArf3b1aRCP1Xf
vLUuynQVwSbzG3Ec8zxofrS9BcO7gxaTLZPXu+sMnS4X4k8xAcFawUGHaVIaAL/O
0nWfGCpPSnz4/FXgQYoEpwsCvYQtZBeWxPV+gYgdnXiCVBK1RP/8UF+9EZG2yrFc
yJQc/qHfTUIEGpYhjkcTuLuJyOXImEBRa2F3ghQFEMWX+r6I4ZhSjnzLzW+PSTk2
95TXl1fBUEmY830iBj99x5VNmpkKSe5Y/Np+yrJKGAciSXD/TLlbn6Ry8Z50cLDx
LDltlrx4XG4nrafmo5YOo7sApRBQVZhRg1mIa2E05T7b8vW+/xth9z5+uzhTxpIO
RAHDxCOsmOYAWnH9Vp7pR6rrMzQmK2gmLBy7wzY8ETiOH8FAnMSCc5rl0lwmM69r
46FJuo6LLjYY5zvitv/eTgvIP2L5qHTSmx1fOMB5Yaa9eU1Ak3+DUihE1Bq+nOAr
9WxaXu/nmqM2CrvS6J7Bs7iTwhbuHUilSProU9ms8hL/IgVUk2R9lbKho/MuTV8F
y20dAfPnbdmrfTdF+NMsbz67DmQ8u1LlBTjkzQGpagfWht+ZzZi5RUEvsuLkVtP2
vwoIEMfLt67fBg2owtjYBcQpTRI/HTOYTZfBWvydHhNgPYsrS28msmK31VK/eU1T
eblD5oGHmtHoXtTstk96lsb7XqqjD/PkM9JUGgkZsvrzj3BztQB5i9/CVky3pAW+
5Mgpncr20SRQ07Ka9rO88MP0XRMFPYL4c7IQyuzaEKIZdFGzuahBo7cZ49BPpi5o
uwiDHLZZzIW5LKVfAEmUD1XaE0jWyXq5geZ21bwyOgLtqHVRn3DpQSVpWdXPat+G
iSiqd3fgJGueqYnMa24MCQ8eyuDPl/L3tOcgfz6dRRy7pPdJw8DLmVZv2NhkH4fO
g71V6PBxVQjMgyB8Ibm1k4RWIW2ZgMg/zsLzj76xc/FQqfkhkjtjELZW9Du4Bzpa
t4hCR2M6ngNE5LwNqICpFutSoDTjysDQdBrDwzDkyPqg9Yx6tghDlO27f7ZfUZzX
ZGyIxI1Fr8OzwBRDFr4+KtNh2xB5BUxsmnbO8CQHKpeLsL8+1bumuo3eqac6Ka9R
kDPsxkZWSwQGCsh25V9e7LFj9tggB+g2RdjbdU+kSW1tOW6KTWX7lzf13MYeaA5l
uvQOriWlFMMW+oHhyOLhu3QlFCHDFAvKreimuN8bD2BXvcFe2GEMi7ybQAuSHI8t
qbhpxsXLRc9bOti77u60/Dq85BZrJaYa7Hgiv8/BtxWh3AXyDNL+EgYnfZ7TgmXZ
SEZVi+/pwlMa6wYX8GBqZUscAJAz8J0CeNqbttYkqLkTIa/mDEBkyJFquUXu/5av
VixvuPMHCAhz04Ntlb/oWjVVrQf9p2dLWkMEqjZtE9/qlKOj540dlEGiiZX654mQ
U1d5FKrJB1V/4Z3SZF0LYxXnAwq7yGHFHJjvp15E1JkVBx6/kyr3KYRThnTCzN02
B7yR5RaE334JsWa0ujNHJZEl4+Cx6dI+EBPPV/Cv2d+lCukjkjYA1sbZYkxt2z02
28VwyuJUfS1l2vUq5+waoVCr+ieHlsCc4FGT+8jaTjAvdlti6GtUBt/blhElF2YU
7AzUHBxz4qELBjpACCsc9dKml5lhmVaWlHbe5EBOux91J/hMYHwsYsO/C+8iHh/E
m6tEKi1B29+rMIApybAPErJsIzbg3Z3Ttepbv5DMbSaHV9bb3u0gkeU53SiLhV3Y
zb52xzXZB+swhPabDfuvJFrioYiD6KI5LRpj+vyU23KD5qWt+hQn9ienI4RJqgjM
ereRqsb22zNB+i9nKG+g0RKMT2XXNqzWgaayAlz93eSNA4OIgr/CGoTrku8n4YMx
CoZB6BYPDPNcPE1sKbWUOgy194pTJlOHGMH8wnu1Z16v9fC9KQGx8OkNiQGdVZea
PiXP7cKqv/PuX7itwUFJY00vlTO9D462/2PRTLYxkf87unvXj5iH0Bc084zyo0bR
jjDQtCD63qalr1jmaEkBEFQEYtNV6hQepWDc5YeqL+LQRryiHIaowKznTK3kOrHq
IFpAyBI8SRaGT4tLBSZCvr+ZupnhBXiwDZ5HuXtWEzt6rl8/A4DHfeiePYcaqn69
0s7zERhOmsQh5toG4z/kXKFQXbZJR6hP0BFrAglcLtbWJvEL15nymDAhuhK00gJq
1MvvaRLv0rIOt7gbw0mR3QudECDD/dadgi/ZYTCtEMenTs/5QroaQ/haoGZazofB
R8HcWe3PliN7on/W2lVWq/821bT1FliCexZKCslkzObg3cxZJcEc/cN7WcMpcz7j
Ow2xv0NFCb1VOyhAxXWbNyqoHQP4+YzdcCtek58PN3KJHeJwYrZRKWOGfVTZbABq
z18o5xwuWagoKLN3NllMJTxuvf2khIOTUFKBG+Ax0S5mxNLa0EzWNAEl1272+4IK
nLFdlCAH1ce8EpbkBO6EkU5OI57j0Xjf78u9Aqq8Lyx8pHxV3HjAfxPQtc66NucI
O01j1fV6Dftx45VDToY45+lOeeBdAq3Qt6Xh93Ylsf/i8oABWeOnuxHSGTIYCtDb
5ZWxo9Xj+qm4EOnzITm0TadYNOeGSfutjlESaGVOI5Ci82mQy9alN9xpaxwhXPbL
V/4u92oSrq/LwAKa87jB29dCKk1/n6uWvUUF141VQ9fLMrd14FIX4RgI7UUQOh3T
86leF4/+Rh6jVsR+wmbJmo1M0z7UozwesaPh1VgcfTiqcs3+3e7aIca4D+WKeAhp
T22Bg/5fEMH4xf5xn5DLOpS1ftW2BUhKKJ5gdAY5jRGiB+N3uZr0f2MxD3I5cFPG
Z+YZq1ixacrLAqNmVeQW0GhFZ8P+QzOUlnTKf8paCd+9eEjk5Sc/SLVLYcKX0Rsj
ZnEIZ4lePidoluNLgwB18nOMkwiO6CSvKTrcbHNXFBORsEl8+5UlTid20LJHQ08D
l3OEaTIUKl9VIUUtBG4PVfUYVedq/3kz68VAIuLnAeS9UG5iJG81+gFX+4J7P19m
b/uKk2PZDiCKhKPnD3SudDEoGD0ki/27ugLwEG1GmZefh+MtAv0aznXR8RTDe8le
NuYrYZE6VF61EDWLuRAS3b6wQ1rXV5fszn7+lE+68eEpbAgjw3J28Hk3aqUG1NYY
oC3oOtNyPA9WMS23zmIfVd9sOBhTIGTiYPeztKyWsebdcz3SFJweBQte/1k3CDTo
fZf6D0kUTuQkmUSphwim3iL+B5LMvxqRGBTzsjsRNLPM4MZ6GwRcly8MJPFsWV2T
OXPZKYezGCpS0uQUqx4xmcaD0vFs8oB0CM1V5yqzKSGWHm829oA0FpSBZ6AhB0Br
ooJkD3yfkE3F0lJKRt5zxbkDen3Vg1/urjBd5Glx819oOAJDfbEUwY6qlPtZjVVi
zp3PWwrUjlubBfExEX4J3i3XArsa8loJByHDteVOG/vVN9ksxBpbvWbY8rvLa2fs
HILF5R6tCwx5IbRqefGuH1z50bclP0mahIuXA76n2UVgSENLrXFrcpWQG5wbhqCn
tGZomdrimN6vUOm0tFHPfhO1mOawLQaAHG1fqvwDYgujTCTP4bVBkogfV0615ARw
H9EJ7oKunK3fgMkYdV3O23zmR3IUMkcrkIZZfp74KBTdasKWaecm8mBpVvYL5HO8
fSDRwyhaLTwAik2N0F2GdHyfuqT/sjpIzjkoLDZOMcx5OtRKbdoT3G/INZaisqlL
SrFlFMV/SodH7HLaZrMW+DH6dVaTM2ciPuobJ0aEkRXndCzyNrXkzrlgwic8f8Ir
mnav/y2bEvEdUY425lxmIGzdGGo5lHU/wnC+86jVVnzeHK76+4J4ecaLXhiWxSdW
qbZKXZWJodCQNpOnVGItWXW3L8j3UxVygQLHtinbzi6Ss/3gIXdbcSWQjfkzFsuw
NWSnauA5aTMoFOcz+TzsIFg/ahM0EHdbFUP5EGxJ4V4BPn/aattg5IrnQAkA4I0C
TQ97gifflrhEVS0xFXcAR7hzVJtwOWm4h2cNUBtbz1Flg2GYR2KM9aKgYmeq98MC
llaBiAbhfhG3c5AdT2CJmRHGgCBvFh/rwyZCWChSW1aMUt7whoPgGYqcEdRr3hAG
G1/V6E1lS6d71aYzMKlfA8tw48eWvawY3i/LtH06rtPMXIMcYHC4cZOZ6IZ75/KA
f1n/BXqFvKp8vegnKtzX+2l50qCFGpS2B61H/ScRD0RItuYXOLCGe7CYXH5ZzaQE
bvNwpQMtJnO1tmF+MS63Yq+cx89yI6VzspF1sb0mg7V+4iaN8de24PoP5sxC4z+u
wSV0E3TXu42E2Lxoj4lW/DajwIImeaocWhgewXWl24nk9uipOvBtUgnGhUZEit98
WRRvNBZRcGZgq06eL/u2X2TpK1ZQz1zW85wO3u/Ec5YU7qSQquGZ19p7EknQm/IO
+GEaZL8pa/OwmBwE65OGDS5HP1DEE5mwZ09HOSHbPAiC7xE3rMhtnSeq3K3wYO07
pd/93Oo/fZIpRr+0ljQ/kK4ekCHgr4NJ+rbyDxv8gGme0IdqCJ68RU43KLTatc1o
CejjU8Ny5bJv/Uk/Yvtftc7jNbnRm2isvV9k40rpSMTCTVlEr1N9jMF4QfYsxKqu
ZlPCLS2Zz4lhYIfm/VJrEB9GAbxzocvnZbnMApBnK3e1h5WNPY2UKt017/Y1hCiB
5xpM53Rjz2rPgF/Qnw/rrePNeIB3ceimJjipMt1oM5x4EHt/PScfXBvaDbY+W05l
ZSx1sSEXFORkfAgngtIfKRAzb/tAvCAY3tNRh8PmTXa6CKaphPS4RObRuY8IyEWk
eG8rG7vzJyZZsnxKhwA8mSCTTfErHklqHOSqLROqozv7Ads9Ymh9PXegTIHUqKKA
XXVnSTDStBIaTuZpa92m1fHoAA4FMQJGpRDqJ6Bu/6f9BpF2xt/8smNcqMiNw9C5
sAq6mwnChLcnOvRrJ5aLsenziViWX9RS7OclrydKogPPazx74G+FFEejby/qqeJp
3RlOp29ha4oZpiIKbpLkZxDwjBZhjRtXrVs1OqkN46GAlLVRiOjeUzZguM3/OU14
zu91g5oUVS8rX2Py/yav9oN9+KBI52ABYXvP6r8r98m59BsE7cF2WQYdwsC6zryl
KPg0Od45/p0urhQiNNNAJuo4zbutfS4Q2bvtKRsFJl1Q1wYiSiojoSV/7blmHtu7
h6ZhgJ3aO/0orxjLitvkkntzJ32egvSvFVxt61zvwYU9rdPb1SC7ztoaVYzJp+C1
5HyuhJirMjmdi0XXbu+SkxPrQWAkB2MEqjCDv/lQ2w1uwtLqzKE86rz0oxW6baL3
i2w8Igqs/tWgpasrWO5V1Q23+Z0Yd+LZ8SwA/AkNbNN34OfkirViUh+dPsTji6/C
YFWMqKWIyajAItKlLaeY3wwyRwskPPLMNpyzLlK5amkk+mVC3Yzng0DKGAAk8cbf
zLzVqsAI/ECmzUjo57Dz1lS+3cnT6v8mx7cDvvhDVHE+ZZS1dfbGvrsNmm6dOsFS
jOyKggRGm5jE4yd+Tw15QFqJuCR3ltfFTYO/WVpqNwMKv7ypvonjFX2o0NWK0KDt
QBQ4YzLJGySoDTSwKfoZH9HHeKoqlPbEMNSfohZ3fq+W8xgHatc0+W7ri6nTJmY2
x0p1ubRs/Iq8O6RRcoEbhMMFhu8wEcmQJgJHy4/LJWwoy2CpP8IGh4kAboSCsnRF
7Ii4TOYAfD1RZI38uuwKYfpeLB4qUuM+ZnZnDbwOt+IsBqcGpDDwOfblWNwRASCK
xu41K2seqNj1p/N2xwsUvR6MgXOBArW6894p3bkJqcYDI6MxvmJK82/2fdeISBAy
sgCQ8RlPeSKplkHKEWOx9S+7uQOIAk+4BCRbvETrfaAGvfsL9FukCFyBviqBqX/8
O9twB0G/KDOeK6ku03BNXTmKgO5bTWJtY63I56ucyHpjgy0jRqUbLOOvva36dNCM
OaaJJVtK3ROmPpamhX/CfwoWaapnZ3IdGi6uycX2/C5Zgl6aUcCMY6LIeiX38CVu
oXEerTyakzUYuH9Qm9P5NPJHrumaAyFU6/Kld5sPIUCh/1fcOLrmdbOP26LNlWZ4
Yp9qfOJ9dwwrBcXtx9JlC+mzQn0TbdX+IIOdqW5KMidDmIWMkfnUc4+YSYZSkQtp
CFjRr7jt6RGy0LbTcKIX9vAOeRF8uu71sKuATSPavsg+38B62hofbTni37fumoYQ
hgXTWiSUtmIvinDFK3MsBmXjHtqu4GNoMXf/ffeqrPxRmEFZYJGJSrUurlgGJKi3
NVJhdi7QDDHVUuPT0KEFj8y+vPFMKqbXVvPhlA8CozklhNQuLlxlVW2nsTRT/laE
p+0H8GTnPLMgKhWoHJMpwsEHBDALPKRYyZz3YLCNKwHC1BEwfs+e0QjDHoXGopTY
cuTKmaXRgGsuf1w4Nu8bxptcUn56CHn7aT8UaJwCdPvWaE2A+Zp62iQFy44noNtj
xF3sOg9lQOzPH3+QbTblthmnEydiot4HYGOe3FDqkmmsuvOHmA7Qgo1jo0YgtFB5
3O98CndZcyLmdiRoO0DV48zaD/HngmO9wNQNJ/Y1J5uNg8goimRYBuqWo9QGbTyp
a1PcZLhUxOXRPT49YNPUUFUUowliCo2UhGQ6ZeSEkqFS5idmWnREdtzo3UgyHyIB
YU/0eXCVBwkPDvtYsue5WJKvmtsatDz4hIm6SGK0RRSJlEfj0JVnKTS6kUYk+Pma
aC+1L3YZX8jtVglqmCUpbHr5Rq9eSSBqTMNzvlqrJeuLd4ckZYFNKosyHCJf2EZ8
IdQ8GaJuCc6ikA5IWlQAKaPglzxJKOAhdV9XFxdSqH2swMGKOCHOI6FubE9lmtVc
hbhlj398Ozk08NEcdGCsYtF3djA1R+JsUcLg9E11ih6wS/2EJ+MaS1f7JSbE5soC
GP3n5LjYkHyAd5r8EWRMbqUnqgvzJ1GFPqbt/s3QRvlxSDJpAmznS+KRzQWSnmfq
QmfKW/6g7IhuyKeTRxqRXFrjGkpY9Fdb7WUaxnLwGqyWgKpxPNxreRTi4J/g451k
t+/d+LfxWzeKJ5UMedy0JYyKN711hBovQQxNM2v2Mp2OzQPYHL+EJL4hAzn5Iv6m
ZHXVP5FYwxw5v433LHBuAYbaKD6yWyq0dJZZfhajbPPmSxqRvX/KdzQTilXVeWhh
JYhE37feIzsq8zK/YBX6FJEbR1lvXCYguDgj89C4Lbq3hgzwtukGkwdEkEJaElwd
TjYQwmKJZyWX1QD0pwM7leInpcO7d9O0hP3/FzemuqPkvMEiSD+a/wQ95Dqjjez8
MlrjnxZ9etwLSGuTY5BiTz0kW/GXZ7RX1Tgh3nX+3BAt46Rxa0FbPqSRrB9rfTVi
ktbPH+XJcSulPMAPab3IimlSwok1NJ82ZlCko7gnGIreZoayphNW+jCMjmQV1B3m
x2kdxZ9ruVCZ6QQ+W7Ybi+g1qkHyifhXkseygnsNOKhNUKL3td1KMNlqpT6Tchdz
uGTMu6rj7RTKZJw46hcRs9lzJjW92kU1ASFGoz2ZUjJTauMFQByL63zPA92jRQA7
X70Kg9Exh+O+8Ze555DBXml1iuucy7UD+JfWjrCmHrRLCZ/YEsQ+1FiSJwdiPcXZ
KegiDFIOcG6qAbnL8OzOEg70BffXBwSJ8NNA0EzPcriJRRK/1aNtrVKo9vey+s4t
owAQQua1gLouwLxyLJvbSy7EK9jlnPEI9/7n0Tn3b/fjbkE5KqbkYiKiebgyF4SM
JJskJQija1NDfAHd9dEXStVxIpYALURA/P6TuytwqkgrSBQq5ogINNhHhkrynw/Q
9FU0N1qed+akuayGQqfQDvqhfvl7yyXvNEyL2Synh6gRHyUNhlHn2uA9gM5ErFuZ
l74A4yPl9L0FGCPp65Wmt5oe15esjZZwmoKdCquD9S16/Rwq8F8XW9zjbe6iG9DW
IQFl4Almexeqix3hG6NeiZuOyhhxwblmU9sbNwWmeDMBKNPUEFDkZ2N5L9zHSrG5
j22dcSFm2GWivh9iKWL9QTIqPGrIvTo7JecnlfmWw+eGIGDbsmPprBXLFVqdIl6I
2BcKvr0SAUigKotbVy5Q4zGJ++T5Npl/jLYV3U/axBotmTH5vEpDaCG/zhsf9d1N
LIApcHrvX4mm9fNgGMRe+b0NlzvZieoRDz4GMCzcRLiO3XLJbMWcB9tdTbk1UvQb
aPnyJVqa+MMQVntSOwis7oEwRR3N0z4rUY1Iy1IBbn1hLaWViFOF4uPv+NMA6HXm
xUE2iCyzXjX9ARq+b3s1Ez0IplrQE3urbg3SZiwQI06gT0hLrTw5+tBx/Bw11Rvg
8NlOnT41PYdD1G0McYOW/rB1PNRzf3KwgkdLNSPlS3xwazIkB/vgTH4Kd7UpDxft
QeYX4kO6ZILhxMHlwyE4GwEt3ngHdGHQcXXHocOdHqnYV5O3vqayyIaFL6sUPLiL
7dIrK9yl2KT8bSpDdb1j5WH3kdEMu+v5S2aghWVknnTPBaP8YcpIj6FjoFcmk47V
mMtKcroTDK9cfZgUWUiqGoBAUiWi3qZfhWhtXEKhrKp3Qx1he9cEcDsaTGKJjqjH
IZSYOqdcBxxcyNpsfsXXCIJ5Vjb30WFqJK5FwMAr8SalT0K1io1vaXzYM6kjmccX
k9tJ024i4xybZC0M3IW/w3XM+a+tuKvhXnzofitm943RPxSTGhFbyPbyDr3M5FEZ
3JB6a/gJFmstRPTAg/1ITLG8I5WrszTkDn1eQCdu7hnnZ7U62nea4cKuSOesZqni
liJVTp1XIhfZ4oAhUPqnbeX/eATWo5xrDW4MHUKbEBs/tgTmd0eUoMMIb15efrFZ
2Q3tCbOedUKxaMxvWEVFD5KbiZ5JmcJDVDZsMYXH+r61GlBOBAMJNCCTZdwGEbyh
oljZSyB/mGfJiWmfdG92gVFp9/gCX48QCI68k7SUfj1DXmGe51ku28NOUperDy0Q
401SyN8GouJigJaagP9BiU1GrouYpEQSa4ew05ZBzaNx557+fm6AQ+0MVlcuzNs7
omvJ79A3560o1RMMyGnYUQiB8rN9luqeyV0+wzhLgdvLH4iZEBJ5Q6rN/nY/mg6N
WC62lIKLkavmwzPkKQqPtjuFRwrGTfWgFv/J3mAdsZFg6l9IRuOATlcXbD3GBL1o
eQFW8NV7L2M0qQ+9O9G8Y9bk20IGwRWSTvDzkX+XvgweRlQiNAA3pXlB31owtooE
piUalSg7QNsGS4g6KiAESazCLoL1pp97X42Yf6GnDu9KHI6VpssB+zVglUu9bzwG
pmLrnMiGDcaBLgbUhpUjEqRN/wqDQeHXd+b1YURZ61Pma1zfPEW6Xmevq+DGae+a
eDIKasWYyPf+/uMlNj9iEF5yO6qj5PoTiyJuQ7YrhapOk31CohuqFjxLtTGH5sgU
V6hb7i3ObLkXjTQgIOSc3ns6Et7C5E4jpB3TIniVsx+LlP8RqAa3YYsqa9KBimqX
JBjjwAqjsBNSsgiqCT+jYY5UuGBz76L8FKdE4zTjuR/25lWmmWsJ0JKeu/GHAeSD
Y+0pvfPywf+3WqQgtLw1j31JqicPod/pbxO+x71HLM6QB+4MYTzBXCJr7+dE9IBW
oABT6pucCdYyqBb+y66jcf3W5a0OtW2+APOpU6RjGoipezIJRMB6RxE9hwVqfi3/
/lRQFDad+wfhOGu7wukAStVlfjHHxkjJeF6nfDf/xCiEhYHRU+XmALRzWzdUJgmR
Nl2EoUjurq0YH6DX5XrcSLeafXYeVS04UR9/01SdaoOgx6U54JLIR1JmKIbxEbkE
hohza8wDG98bJCmqm5gDkih2MNo/QJ2ZnqMlBNtJ0Cum6hD9ipeiFVWNO3nJS/fQ
Dggk9ySod37yIesHgH722bLL2izfk6KIrvFxk2DkwR2uiJ0oxCSUhmSSux84Iwpa
BDqPmV2YD21Gx8Gi+OaB2tUw2z2e0QGvCg6I32vKmBJLtIj8GLPfQdu/AefHRjuW
NfcvYpDqBFBz9Sjqmomvm5UWiqjmM552WCU8ToZ7fmBD/QKmDzP5/1etEGFSudmm
rrBVB+487AM9voqhLgnU52wFfpoLQu8OdqBgp/aAG7CaF77a3porbljVGGZUKpsx
iKDfmThkVMQLGuoiHeWfilbw+i62pFGtf+9ovdgcHftkupK/cdFpnZljFpR7KMLD
qln5Cz6CDqGZ+ZOH7cLjpmbdB4wnj91j14bnCTQpcOn5f71Vz0jUu+JOlyc0s7Cg
BnHHsqQxu37Hvb/HUCKjaj3fK0nPrABqftxOsfSfmI2PBSq+eWF6uobzZzegrAtL
iF04oqGMeoh2O7KsIyBT8s4+Jt2UjfP7ShRn9rAlFi0sjRZonVFT4kd3x3zaqpUv
LK+ZCwKECAMt796B3ZtQ1vkzbSR0funmeR1wKreRFBBbPQIj7vs/U59VAms6NXRB
ELjHyVWlMSYtkW9WmbiKDVUWZmWW+8gULYAinlztMLxjnKMT8loa9fD6ASlCBJnp
Gjn78bzgK0od4ItS4eH8Rx9TwvFGuCMoq0FFmUc0dHGjS15FnlZ1uglfCroRrA6G
5ocRUQECpmUT1BOamOa86CXbyWz4MIW8tdsaYIShkouWs9O0iKGdJPOj5pjdZOnp
XB/leaitJpJ9lD9+rDz9omfzpj/omG7YwL4mdX4h1LfRtKYVwl4kVIMp45dfBQlB
pg9r7sgleoCHY3si6zmMkRQCVZZhcKPuApNvgxEaCjecz+Hk4Od8bFqz4Tf4PLZT
nGlD5wJ+dchKk/A222rzWXtdrFZhG/GElVal3QdTc5agY6YuanGrtJ6CqNXYs8dN
2qrzSFg3cHTxpNC1SEiIgkYFALk2fXbdmRPkHCcInz3+7G5W9QVNa1vMzk4BuhQP
7BbYCgwFinQe6rjGsqwkkcR15IwrTcM/WgxS3YdslZw4/EWO5T1ASwaYMHIGfvWl
yaaUAcYUIkwSmDJpqRD6DuCk8J4Rk/uY5/G08MRiQniaF3kT+Nk6EXptFg+nwovW
CpzsesUoTw8pr6P6aIIH9mARRkpbmjdYAvPFX3kFDUyy8OumngCD3rh8DZXRN2tg
o+Kwqg8i6yaAyHyuc0V6aK0d5IJxih5vJKFwp+hNX+lhw+jCSVPCyKxqRrvht3li
Dmp1yrUXkI5mlOm679erhb3/PI2z26tA5U7YEsOCAUBbNniIuIjp4FmWALjVyUuj
qyUYIR/Y5fP0iUsBKRQCQkak1VVnzOWv/RwwnQecssyoXw9Pbs71S8Mh/duwc2U8
SxK8nZo5Me/NEHW1eowXL369B6BQd9IGkRUXcJNQeBfaGh8zb9V0OVVY8VQK4/ti
FCReYq7phYDIXigfWQQZMPxsobwyOcWlekQTVXfpNzZinC7WRfAiDdTeQjMFzhcb
KsbGsAx6ZiUbF2Pb9uJwDCg+uqHGi58peP8c4s1QgXCpP8tWgDU97ZxWN6s+Cxpt
10nMJc+HBSAipd73+nAy2WJG8BUuwNtKx07XcnOHhbmbqTqHiERnClhlIydPAiqa
IX2ZsTgC3wm1/t57UaWU1z3DUFmdkR9GFpXDIxPiI1Pd0R2uDVVE64ZVnSVgOXV/
ahz3CksD8ZaGM5hMQ4JvK4MU6FM/FnpRJ9KSiLr5pf6LJp9tJrP+P5xCdF/KYhl/
xKm9xdsMFz9XaD0Zc9b5zVqClwOluz3qwaGFmp0I4YPImT3yUHjzrjrgLotmwvNS
QeAWcGA/kjeXwIpri22LTaxGUizFLgUwexcFnUCIYfwgikwBsZmAINVWh4A0Sq/P
MxesJjiarJDOlpFNbo11FjlQLSzSuSr0s0hb/ALPY8j3twAe8cw7EftCiCx17z/K
t5obVRW1EI9vie8ey5kPKmujYonfTUDbFUm85X6A8nLxDP1qRWn0611dSTp5GoZe
ma52OHGTzyG80jK8Gi8NjoC8S5q6mxHbqogX2IPI7rqMQ2HA8y+OMtQ5KO0R2d4M
4J2RuCrXHITbJHzyumjDfMI0XEet6w0MF1gMy/H+Eh+BjcmZhM4XPUxs7da5n5xI
+M2p9M3RSGI2NiK4uXjyDp4G7LRWyfNw8j7EWLMw/q3g10i2WIE2z1OaMHNne6VB
QKH3O/roLEMFDaAnIpw5YcYDMrukSVwAIc7JIB3IQkrcP1+62+ICNR1QHmXtmbpA
BcGMTlnVtWcrySxp2rSfdrACAzLI/3SPM27hBvSws7e0ZBPzIwu9MhLN2EC8fx1J
0AhZaEsN/jpuOK7hYLvTCpMYbNe+GTXgdKAMARgK8gRRvdxaWGII86qO/dzXSZjH
gh+2cDmNDM16dxbufegG1R6pDvZDYTpYin7F7dWodWSXcjzKI4bs59xP4N4bjCax
aGc1lXe4/77V3bbgR5Jgm+RXLxdgYXQt2lVLlDxujFl+HYKF9BQd5muuL3/1tEev
mE3g3e4j3C9wMnXxom5Wjb2DLKD2yQ3m5S4Zv2HzRr64ZzMdjX+FC0fKxC8sxki4
jDhZsyFgyshkRBadxxmRQmX4PUMkAN8vBbuuFC1R3bMaSbuoQ/24Qol1OZQYs2oO
JgqdGhXlH3zLGYtx0ONVjEUUzvgEqDzNBBQ0pWQJr3JvM+knClySDh2Qu8mbMdlY
BgnMppjlbwfkzncWEy9YljMHkylBj0b9RoiPOtWnSq4lx9nwFqNUARHjn6cOZij4
eaLMlgLanH/No8rTRjn6on1QbQ4aPL676ITDKfvt3X6F8PqIXFn4k2aZ6axvRfAk
tAWIGBG3m0nlHnFReVs6NS4TcvTS1NDN5A45OCkyCi30Ym9ED5DMsLe8k0dtc6+W
QzP1eRXY5E+9+tHUrDGkpNvinxNR9jtnYKOOsP5X8NuS2nYZTamjTS4+vR0EvC3v
g8XSAqYjY1zE/5klcbI+l7LuR0hMKiCtA9fPjczJkp+Z7HiMMnNNvSZE5q4UYczL
AzK4+34m7Gh5qPe3k5SE74FUNlhO4n0ro2KM3Ecq5C0e13dZbFseAUMR7SCZXKT1
G4vcv90FNiCdShhj/jLSeQxt8MrU7pvvQfanSNIUbdDaBFtLCrKpWLnSg78RtGTD
YvBhVlCx6XA+HMp+1iS+mRxQZZxLdmb3y6Td+vwYFaB+OuOwhyX4ZlTZiWJvfAae
0Dtu2JypQo8+6WLF90TLRK+ZaBBDM9RD6Ju7iEOVaBRnHb1dhdjw5PSwl4nriAVR
9XbetNg/1pXfGnEkX7rzLplqu/AzCLUSzpknqvQ/Mv+hA94TH0IEJObqoXCRfME2
5wSlkMpr3pRrm2NXRI4Jcy8I9qn+tNVxYFXx+weBKb2PU//5NY8YOlwjRTF53NOS
Y/CJhX11xbfQjdpCkvk/X70MtMBiAaGas5+ClhGSRpfFD+p7Jcar7nZmQVdJIdYf
mBoa5yFQm0eT7STNMYX/fbrKOW1dxntvF7Elxrc+n48hqfE2ql1dVuS7LQiZ3you
vb+XB29brZ5nuVEOFHNSTEos8yHZKeKxT0aPfiPfLBwd4+euWwMbwXhT6CnPNkFF
XCP39j5141OfqoTH0w0w+0xHtcrtiaV/Bg/7OyiEC1ugQq8GQbW9V1BKiyKcofm6
imJuOQiuN2VwCZDzHQ+nZBHtr+5loPCVarwtuvTJmYeSWia/wikXLKlgE3xeLrSu
NecCx6jRKisN6N8/W1JkbEfDP5HiDpnBAq8teUjhPOSwEymGosHXjpSd4U8/RnfI
KYyYKbPr08XoSMkn/s672nYvDxa16G5QABcQbv6EO0hsDj4Iuzrul/zYWZiIMTgP
GjM0aFCU+42VngTHQWYZ0qGDLlLTipK62HFkqxbXFdOtTqy/T3pc1ub09rafVhbV
gqvImUYvnTSRNMsiDeABBkjhoU5iJVj5vocwWL3O46Ql2e/UsF5hFJhBWwDjHHTH
lTvDpC/6Kjj+d+m6bbk+lhcsdHDvveQ2hBmcUe/xLTehu3aLQwN4P22bue/PjLEZ
37xfgczjFEIrymymoEDyz/fwVVt2CoNLHNSgnukcYurrU++zEhLW+nUuN+TD0NiM
ktxFd1sMAI2+63NgHyaI2QpQ11oNHbEB6OEdU20hVLFpCsz6VM2lSMvpd+SK/CTN
JCN+jlJT3CjUKc74mZNkP73ecfSV84jLM3skY/8NWhZm4m2Ailt35Wz3GrsgWW3H
eGF47tA0ByLq2rot08iqZiXzOF7m18pcW2KIfSgbXnTnmD6STJBQc6nSmvi2M/hN
wPb5K4XrwCt8xf3xw/AbvRT0cYvpsOhPSTTL34++4Rwbvxj46J2M0UOj0rsmxMdg
jgYHH01gH3wgSo7vW/HFHGsClCLcZ+ZxsnHqCiMDOjsqoRcnpptpyojN8GFIa8+I
Nt9YUJDWXqLfgfFF12CHJ43AWn1C1ZKZLv45d4BedW6kPPMQiMgsw++Frp8oQ6Nt
dJXyUhXKNoBPVWEYSZ2jc1LdY84y5Sf35ZFq392jAMhxAsm93JtDJJLbo2ZQHMBw
Z+oTYXbkwQCOiEalLfEyk+RJ41oZF6NLRnEN9TvlQFmAf6n2NZ24rgX3TJDLPu5M
xJxo2GgEbmqZpoB4oQ5olQ0QSPlRg3sA+M6jTc6rdHjGKJWsDo0ebY0/iE6AL6+N
F21ShHNrqetRCfal6XegvrvAeMBFngiHIb6DkXWFjrr/12pq46E5RwcyhvnlWwis
KqZHD6eNflfVZaBxUJN4uZHSRjDmfU4wdWZZAQEPC2MYp2dCUnhzHd/gEXi5/M7N
sCb/O13oDDA1og4Kq35JWa+eyG11YMAnIEnFgWufXu23pm9mRgwoaEODRyCjW2xR
njgRblZ0oGzC1ZGMTnLdOHqwNg0PEKzb6PzhS/ahfEjrpxwQPXE3ENHhXExc2LHK
BxR3RYlEXglXR6sJkTmwgCaLHQ4KTzWhNxjZ0k9a08LuwjWuiG9NptDNwKatf4CQ
CncIJKfXS6AvYUu6eiGgvNJg7GuhpE98gzZQ5M0xWGng6hLjFj3tmO855yFxO2bx
36xcUaBS3pzsOl8Vhv205CxHiNkZCN8Q5Cd7E+cMoqPiUCgcaa8VCUyEtRiiJ2jz
SwGn0XWYUtRdW241J5Y6oaUU81CW6qnLukL6TF3J0j6Xazyg21jdhCS53Lwvpg/w
6VdBDkLjdW2uEJtlC+IQg5d95OzcyLmZZ9FYBJrAMnyZw8RuUcGZ56rLcegt+gT/
tLj7lw+IxwUcVNhU1sIZW1BH7AhhsncbckFzvx4fijFQi0QofncgoUQ2iXe+GGU5
+TGNfuOgdkjxz2V9IwgxTPDE7WYWEq2exOg9kpux+6eIoZu0y/DodjnCU9MloTWP
/f3i9dgU/dJKrziiUptipx6Gi/3Xjz3e+6UFVNVZjUv/Ga57sIskFW7mdc7q8qea
D9rreYImaOIxoFwhQbcT/uKI5Bu+BH7YyBh1MLLmQ7coWFeqcIXxSiMyt30VALsx
11Hi1jJgLirGZ0SbAywZ5dAC7rA/LQTy7IwRIxvfonQ4zLVZ0RQla3MQdEdgo9WQ
jTTFRHcyIV3TApC/evEk+D6RaekFHnfjZMSzr3eDYqdAxO+IJPV8N+cqTit/+W6M
7XUOlCO3WUP7b1AqkgZOti/flVnXjrnJLMA/PY27+nREZH+tw/aaFdlIhbdp38DM
Wd3Gnpgyz1nB/L59BBuUsZQMnvnJCfI1YkYXVL//7ZdV0Ur1lZ9Hq2h2xmSBxIFr
FpK2cxDLRQObTI2aNBt7asi9Ijt0DtvSs2eG6iCKEB5nwKoY1eEloXvPn7HI9SWC
FYrAg+3gz+4f2QTFRKjAQOqnS0d7RSFD/YlLNRhQ88tWlFf8h7Q55kZrOHmDDMwL
0zQKYLm1fo1kuOAagEWHHpZKg5sdGKKPAyaHkWXL43xUNNl1UgC5iaR8V5IXJMfk
FYI4oatF1VNLLlh1Ivw++EtrbFEvz4fROvJOL9XlExNS5pBCIZQysuiflL7sBacs
s+mzCYlgUdhwiEZza9FyHSAp/4xhQmxZBbmBJYbMx5DF9sPgNp+Tq0PhqyoT2JCA
Xqkv1eTKg4IPCwQvucYwCm5XW0fAQDuUiKFahcAAOiOk5Iz4DPfLgbkULWEeGzW/
yXdabs/2ytNxrEMQ6T7MGkuS2zz7BNF+h+vixYl2K4slmgBqsi76VzbxQacQ8E1K
03do6IvZKCpTP1iTc5ZltJ763E+ZkUrs89XSFe1C/xz6JOYCgXofa3HEuIhKqYO1
Bc6yfFnCEAgVCmaYFL87FpicRJtPBNh0QCU54+k5gWwVywbhUgMmVWSNZA+YItKk
hPAhjAkP99zF0+tnRO0qSkZjPt411F5V4N4PCIVjdC7MI7P/pOlNC5FB/np7jelk
E/t3hXMGmVYv6x/CYDgNVu+7VoVtKjBQ8yTI2U+l+j+psJEFGSxBo7/1VH5wAoCN
9yKQ2woBFjWTViNW1jSH6ojVeKrfuwAXR5PHHpg8sdE564Gq8JOUXhq01HwobDWC
vBUq1fRf3NnzLnGoHROwVkodwRJGkjNYMDbU+XJI86Q1HhLAPuejAypjuEYh16cX
/bu+8Zdgr7F2rAAmojhga0+bmha/8qh7OzvqP3HbuJAPtHp7xsiIJ6oOu5CIaa98
FKrrXndjBhLhynkBs+zBkwULh03n468Aldj4ixOxGJvWIs/XrRUjP8gGSGt4SA2E
GY5hIDPItk9158cnpyFEor7LFQmcBV7/ht8KPlnFFxdGF0vFfMF1GxEoR1pzxZBY
hW3TMXEV8UlE4Z9h2yaTRw5S0OhFYgzANiLHHwoVTK/bDfUnGcncFTL+f6lKk4mt
SM1Iy24UTCJi6den/sxAjJXh7alcIehxYo4/hPMf6WFhQvNkWBKpJSyu8S/tEaJ+
s78IYIO8Omay4Ggy0zf/DqSZl7NzVlmGb8T64kNOu9/cL9CpCHbWwbSMQSBiUhAD
08ubVZrFkFnHT3zwNgRJv7qTNm9+yLTzBWLkS15nMSVgm88axVBXOqkZ1M3aJSFM
b0BRLT21oxPgMwmBlibGoPqo6NQTEGM01ytY4ixHjRhoh+d5gEeUb85Cs3Zh81+I
FSIQUi1A9+dC+nuQnh6TpjDgh9teC71qYiqI+0OY4bxpg21vo01zsd3MJGpbwVnc
0ywzQ1wvIvfMMr49CgsGXoZ8yc6w+UkEoNqI1AXB53J31GDavGqCma0ZfHnZQ5fB
CmY+xjpH5T0aaeiMwjrcnisScSV5q+yH+ptblo0sHxzMuT7CIhR6e2sM1Z9Gl14W
1su3TiAGfmK1W2zLu5K+B85ydFVHNdYqTjku3aTVlGbmHKpt5xaGsoul4N+C7nml
+e5v3gbQ7mabVYvvljzWfBxz/IZcJJNjPpOnFwpHfeuXFYKmz12mDK/Edm7kX9NQ
Ad4xn+Xg/Bqm7yiVcdHXt0dlng0qtQ2HJ/UVw8F8lI42S0wHawYojiJfDxVt4XDz
0n5u3dc8qOWVuXc5EBNAvMTtxkv8t3nbXauAr7L+XRYdtS6z20sqxBDQU9Fvfpx3
wcbh71QCnIFVDq+EPdLFIBtXjrK2jU5D9iYXjkriWlg7oEVYXtFFB+oqwoDgIm2n
hk4EgINHsUqX/+hGi/xUQagYV4SuWHhSKscABp+/JUL1RDkm4LNgHQfTj2bAR6n5
3f6zNawppuiaZvo99dMp0oEH+oWJOJ/Zuc85aHa9S+2iHpEyLNFs2BplgQgE91Z4
XDYgb8xbUoq6PIZvbkfrKLiWAoeag8taYoN1M4jmACB9IiXd3XiJSvrz28YNdQDG
2okJeJaMlQKvGpjeYuYhC2EB+UqjWia111KGwtrk39K8mD2CbT4sHOpDzEyi0Paq
doUMvAqKYftYoO7FO0bPQmFhJ9vOYvwTy280xa1B9ZzGvnno0NEQAY+NvRiK0YLd
DSboJo9hA/H43tJmeCtuQuEhuvv95siVDGpsdFJ49kCKIraMpoEm+NUnUByNVoWw
EDXooOwUnvZ2Nch4qbiD5siUabKd5tcCvNDz+KxHD5XD/3RwzqvezWutka0TZfDn
R6CO6sSeeeT+st8QaNWt/q9pUffp0Yb9vNQcNN6kdIymquBlQJtLRIwch9C6d7jw
uQjuNuzFLwTW5vN1sEBGfTGc+Yy7kAuktrPrDQRwWaJdusmpwDUseKdoXYE+kN29
EDaqaYw1uK8l8OyzvYQkU/fBAgzwrsDi0JxcHQt7WpqgwAu8sTpHefNlHyo0P4m/
YdZD+GbDsSUIaYGu99azMKhJYzarPsMMkjDsech8Bue32QTUNrH/PN+wN3kzaOhZ
SZvD7iBnld+2N+QRcpgwfj1Mh5Y1XKzf/n3sdFfWq3l3i4Hv8T1fgQ+5QYUX8tC1
j4wGCpQ42DqsllIXKD4ULgavC8DC6m2lB1YUkK+j7ovtTcDFbA7J735F/iCekKce
+OgOb6LMHOtCMgs5D/OQRm3eVlsOOi9Aw4oS91Kw7G0bltjgA9aii0KqItjaAZ9B
nQyJtd7aXPi89f2lQBAP9e1hvx9kPgp3xAzeAB+OBtO87r9GQRXc2QHRn0gXyjdh
wNGIw88sFdOCkbb4+gtiGLsB0YkBIdoMTmIJXjYCus6y3nNmXf44LH71ky8NJcFK
oEhqGdCrYQFtjvOrCbrWzxlTH16PFLY9+8zUIONKFGG7DD9oajz823usAzB3stUE
2876qr0lVykXX6mG7TAC5umYhSVBvtUQ+4QC2iiX5Ve1K/8x5WkV7eIwz00kxdKc
4F3BtIj8d8Ewih5r4qm/SeKshqzFi5zmu2PdjvC8mcKVkZsgRVr/usiqOhkLZTLn
3ffiH5lKb4RsudZAa5f+zCM9xJKZkgPifH/yvfswRwkZm72SD8N3mNMmO6vW9Pbo
mqp/N4U3MmMrwh4pBb89Owavekin4p6+U7tlgkongfQzNl/Iq1nQIaL31TzBhML3
QTujOKsBUcI8cExe6WauvQKopfzbtwdniTqo9T6cVzm05uzydwDhkprPYQPd/aMy
8uJz+EeN4cq5mITbvXbACVO6DVtFnfnWr99/8CqB+78CSqpfz/KpWQcr81ROtbdC
sHxX05+9TmXBtj/I6W0vs5tp+wlM81H3oLgjBWWa9sDKTMotw+/poGHmXcoaq4FQ
whV7Atc/zppc1GaaQVKTfRZtdzgJipP8s6+vQXMbkA/P7E7IX/inc55LJMolRiWV
MGHZrlKa1/H1SBASYidLx2VDd++8XTVwaGlSMq11rmRmHGog+2VDKxODsMj/O5Po
T/hQ2YCVA3gyc9o6OxsXkG6SOSWOq6BWeJRhKN4empM/5Px52cKStfb8C1E9dx3C
dkvsyqSFwT+lWJGCTLaQSNco/Oejlr2RAzRsdKdL5gPRBgwRIMd2Vblgd1HpBVKz
7ElsOnCazg4fh+he1JZT0wEfptjL5uXal7XSPnzyOWf/hffHLw6aShFU12ZLoDA1
pnQzQcL/1hoJBUTzjTbA7382zzkCoZ7ap+9dkHeSuRe/UUZG2SN3LwUX9xcxUxU8
/q2hx0+A+hwKkWz01qTdmFm89VYptadzEkSQoLATPTi+nyMnAdrOGdxU8Pr3CrM2
v863yWClZwQKpJkPIRZUbU8tOwFZ5biGgV5Nt+CwPcHNN3DskrArx0K0NUhaIStP
P7i2GlzQj6/r7+fLYzbJC+heHglA2qI+TAtkkCBuY+0HgsAzs4WgQOd/eROejeiZ
V99kjOwi7fp2LVQYREp23NNC88iMoJ9cc2K84gnvUxvkBvcaHAplIB6bGQWv/AYC
kwPwWdSiL9WLuKxjgOE1wAKZHz8LXjx/H+Qj3lEyY9Oerkij2mJN4fG2EWJ5wqCU
n1upvHTAdqASvKzNj9fjEFXProUwI9mNMEUqq6mRGjHtS4S9XbJNQzeTNUYoIN3O
mjC9SPiDEsLOcCopoxWRADEr1sQRiDgq+quG466fv1fIpd+5eop2yMXwhVbpYmZh
LNTbGduX1uY7iEiDbeEW20H0U4IxbHuTsH7KIlVJoPZyNN+b0F8B4MKr0M2yrf6l
hWCEgrlTuDdBEpP4Hu1JhKfNLYcH1nQhnqCcOAu680mUBBygxLAdMBTstu03/dVI
ZUhBpTkZnUn51NPp1ZEm4OdLaWUJemliXo5FjNYhRC8Df9tB+DX7Qol2bi/bYJf8
VEB+2KLR0Py58mex4orozS5guv+W26ESr12rpRzWhwJ+K4gOmqduFdxHG49xRcjj
qKj5OESdjNDMPG7cixDu5aQg8GnoUhyOtjosn7Nsb7St7rzQc7F96ny57D8WqsvX
uKRHDrT5uPI+LTHytWvJnMnfWMJvNUf/XWltPMLyi7AOOnYPA/grECtr5Bbmqlne
59n4Oaq8amPwj1ln7euR8yWd+4rXxp/Thm7Bb0mjS/zikJLmTUVPEQIwuSVRfftg
ekZrKdhZ2BX9Cyanjahfv/m+mL7BIRlAAc97WT+P6fjIxEqtoOUQ3kBHBdnL9eEs
tibx7biT9jAc1c2J7Nb9/Zs6dNrmsco4kf6ItNMiVGfm7MizDGJIFToqfcoPPhCT
p1zeg+MuTKFpszaym5xSsWpvDHsvU9l0UWWS8/IURH4LWYXpIApZVPb55YX+vYTU
PQrjzyDaa9kDUKMyJNgRbRdK+S2up3yScS1Xi9ic/dGHjbGUk/H7IqFZBPn+azDV
YrjkoQkS4Hz9Ai+CaNtJwStY1pxw9tWXNVxpbBZW1y5F5yxkUcbV1iU4GUR03QQ9
bctboWm4TA8c/fxUMYE915BvvVLOrSYmij4ny4pN/IoHQ5o9m9chQQFSOebbF6BV
xopj1g2TtPCHay2FC0zXbST3Ax2+gx4WS54r/he3z+n9QjhCJMG7U++uVAITFJZh
H3E25F20MH+eeUHAWdfbw4osB5vOsk+UAV0x8Um/Q8IZ3BdGFCuXbKUQDxU7uQsj
tuLQKkEEr2X5zqcVVQxddiAjxGxR/Ta6hQ0GmxACLH8lCxYskBOQCiFUdfL/QhaY
xVDd4mrybI3qRP6l2gToaq2JekKXZcAkzxvef5AA/Jjn/pZM1ZS1IJ/E/Je4vRsk
cc92/Gd+O5CFnW10t7BXlJGCSbZbW5Q6fdIL7J7Y98RHtkW6FLdxc/MUL/EjUhI9
nwfGv8/TU1m5E+HAHozV5tWmPGi/GUAwR1QqqmODnZ0FVFjAwv72MI3kmkTIABA1
NJcOaQXwTvOqK1aJyiZFDyp0yq27ZYT2OKhPaB91NHVMyoMqUYsJH4zVOS/px9GT
Df6ttJOnEeMcKrydF9n2uygTpFOgT2Uke80siI/3Z3yYga6sqxA7RxiqqWH5dcFi
sv8UrmnutrWecW66jQp9ioMzJdKzJLcjipQLycCvWPekLGaXi9K6rNYXb+TIU2pH
Bmmuoz0SotXA2t/OiTlKsSpjXs7QW34z7w6btT5Jg3YXL3WHWFCadLcP452YHWWJ
qXbTKscA1pqhah7f/B4Mb+yiKdCW/bGsSu+oinf7DgGi+KOkD5D7COliEe4J09RX
+SHFsrT9rZSPyJ3ceinXMqU33Ef9i0KrKlJpcrWI00Rspx+YWfwn2vQJmAxM0koK
zwV5UjYs9vRKp3IjA5pLK8CogwwIXiRNCVFI85ESpP5pethmxvHQJDs/fiSlNEMr
QItoEfyQhtKuGSjodhvAkB21jr0uQ46CTmnz4VqffLkE7183ib4n4jOsZW8rPi1I
22/U8y3Epv/js/fSGa2A+paTL4ooYIvS+WTE6WP4CdRQ6H1sVMwyoZKhuavElTCt
EXKGokmpR+WjdwuujPRGjmw6ElsPesq8ulc2Qd6tiesPyjGR9Tu1pH6EbfazDTQS
m5TWsU9IeYDRtt/qwJtCfbyE7WKdBEJucCw/In/8nHfccjarnoEN5tmPWNChyGd/
eZIpamsEGCA/ptuGuwgBUKDBC3fuOoeGYzaEWphXmv6D96OPv2qmfvt0xkEd5kSo
/odiSqMPVDgMOlB8dkhdjv67DvDHyA6yMaAU8RWls/tK7NSr4zIr3ytD4OBN6glr
qJwXuLGg3kv8rLkX1Kf+Q1/N6HZCmp2KOUiHBfk7iPuXbhKCtvNyo51r3FPAUYVM
sY9zHKOYASkmjMBJRu5aab02VXBji7nG/JNXTeP9o4jAYvJAnaoQyvZJW+mGrhGO
YX8rOp/zvfhZH92MPuNJYbhoQvOjCtaBcyO9F3MMj4vzMT3Rr2O0YVAqkUAohrHt
tlboWHD+SPIRz8RB04ngZdA0wzTcsjCdZMwh7JqCIBCieC68SNPz/x1JuPYWl6W6
D2GTaq2wYCFBz3ntBqXaAZ3hkNM4ZDqpyKOK8qHwMFHrpyAfybNaAdRU2IIUbCtF
5HCBN6oZoT0u7VLgoYIAaKXDsALmWRJ1e2ehLXjDOwhgc710faL8UItx9cH41GFz
08sRWxaK8GN4Q4j+ZPssrVvJLN4Vzgq4BFXYeRCjgOt5x3GJD9Rgu1mL6GjLXlo1
OWU8KtHqWlOuEFAcISYHvUqIuZj9aI/u4feLIyi56Bs136HZSfLoo6P2tVzX06po
yoAPjvt48dlMaOmOWq/el+OwJun7MP9NWEHLY+SZoe01UwP36wuFg2cnGV0XKErV
VhIrJ7kjBOCIvcTQ5buD6CH8422ypLLKKbDG2toDYa2Rpur2A6ppUGpqhRs711Od
K53hgVf9298kg1Uh/wx/u7rIf+FaYbU4Z8w6uKq4DkUbTkRpVPXE9if7QdHnZydG
uUbeZBkn2Bs9xrQLDuSIogYjHADQwMcHBh7SIttGZ+KHGOGvJYSIxL2AB7k76A7K
3YCTofRY2jzq3ZpnxVcN2gX/156Kma0etZRJzXIVMk/blyLWAHGr7v92mHw17IAp
Bx62QsHNRG+qOBDZMai/tkVLQ4DlxTGgOgdYpiGPOSg2SWzow10/SAXANIyI33zA
/oDZarkBQiwQWyeON9S/l5f940gZ7TTICFdrGNdVOKKTb8HxWSkD3RqY+PMHo8ln
BEV2auPDUvC80yoOBLEkVYFHqohKbRpghCtMZQRPSFTCsysfesuT9PjdihCXO4+y
Gs320CzIeMj64D3nacUws9R2OpNSGB1qwsHol1QFNZVW+NJN0+8wGfl7FVoQM9/A
6USv8bLgrux1ivrhwo+0RwgcYknNm+sO558mEPQCZp9CajYPXGppnG9b6tVishfa
B7ydE4Y2j0xin8oucInMInisqxFHkVgU7sE/mgjW0F2+Z1jwFdnp619n742s1W0+
cWA5HkAMmFI9/E7lEUyN3chkyZ1uHwzP1Vz4gV3A+p3+l3IYaTTllrJHXVAdbDYu
TYTTVp4ix4pKoO2TBOvwk3bWZBSHHafx+rqb+KMf52CsTLxGZja+qC7gnjq8QXTp
7rtDa47Xp7NmL3uBFNpnFZtDDNFZe/h0d9TJe69fH86qGd+M9TXsoxIZiOcFlGTt
3u8X8lkqawxWQMkjo1dp8SeMXQZPtXNGp9Jahu3/b/wiS0D3Xcw+W6LaOBNNq3QC
UlBcL1olbqvtB4bc6LIaEfLuwbD8z50UlZ0UoiQRn5WudnOeDthWw8xuLAYJG6X5
dSdSXmE2pVlC9VOPqgv6jYUj1gFbJ0Htwa66tdEKhpZxHBawRb4LjBTgpuH3PtXQ
HoahnqiA0KqwietCSG6p4NI/fQsgeLZO6TKyjjtHCnAUcpL2EdU73bOp/kXxmgSR
RjW6OTjgR/hzC3cOSydHyN11jbSSeMY5OBpHaaIYHunVqrKR0IMIBaKOdmg3vO/G
Zt3faVyThnavnnPYz416w9OyRbwMCc29Wisn6bKTGAXur3PZRXAnK3Ptgx4rV1Tv
+/ftL+pZZdsns9cfzUi+ggu2l+ppwkdu+vVNFORPu5Y9dVR9faGedsUz7KSwRmd1
OV1DtjQFLPqp4IUUWmp8GpXQltJK+SdVAx7orcGoHMPgv5tR4LaLIubDgYDxx3Cd
u4X1aq0GvVgRRUZWwToDENwyYjosNJ/TOOqdlz8fqOIcNPSLkCHz8SVaj8bkdRwO
+C+pNcWByFsxaNM9ltHSB9SzuaR+8U9922GnsInC2MXIsPGiTiheg/shW5G7Qe/Y
7PRzy9n2DHpQSh6xidjZUchTq/ktlrbYnxlDCIF4xocFu3OVdUOWcJfATCODHnOU
hAG1eE1D+KfBWgvf/DIm1Vh04egFHKFE6W1rUCKoEgNjXipv7I48NHVLVlIN6NDw
gLE5pUnyhDSfNunRMVQNk5MBxn8Hn9s0vXxLlhxQf4J/VVADHUKD4+8c4ipiHOhY
BgCVTVSktHXP0Y4kdSVtZdpgJcr0ankSuKzZC04/kzIgm+Pm8L4lrKJ3bhaux8BG
GduNezUH76YsDCoKbgf2VXbMBJtaVOuKr3YzvEerNM8868DcSIil/pQfAoAln2e6
xG5lUEq+WSoI15Jo3KTBwihlIZUnNxBXhPiwsorhvHMIs7F9W42fkliPGnRwy6p1
L2n//3r4MgHhxSTG+8q22K0lVjFSJtFuDRw2N50aV3EkWJcQx7ZDjBf2/nxxBl83
ut3rrhc/NCLQ17u+NH9xqdm2vvrnW31FwcStZbOtZrO5lRGerrfOYI7b6I4gtiUk
KVplItf5FOUfTyKTNMMaKiSrep+Jz8ngvbcwcmH1m9GNXGkD64/Q00XVQkdU3S+s
cDD6SAm4sdxzUsu1Xj/LV5pRzBhCEjF7bnK9rrlV7xxOZS6NUghZaVgvEBHK8Ggx
dBTyq9kwf19j3DL9nbwZ8eVRGsG98B8WQDGZmu9R13bk0uAsNcEPbvmKROtxKjxM
KHnKHxmLmoeHp60eftzyrbxd6UOQD/YvYCHVeYCYHaiJ+tpN3DujRRX03i9gbSIF
ZN2t1hru0Olgv6XRAWZ2cXSGXKC9PZnGlC1M1sGc7Nrh+YCEaz7CjEDo0LHzJt3n
6OKISKsSeJnzqHAl7LRckx7mSwQ6H8y85hBKeVhSl8iQfazNAoFY97LP++YAeGWP
QckJV7DLjrzyVbgWvbjgAn41ssUOHjElC0/T3njSguYeCQPDMqQM64JsmU+I9I8L
zn6qhXr6TLdzZwgvdsAM86RAJvY762KNsHAa3cXNJN4ZaMgWxDQ4gVCoCvqo7Ee/
ZKd0SBvH3rfCA1oTgXhktzt28dPuqbKy51qInTRZoA520RkWLEEARBCq1ubQd6YG
+708MTfriPSJ8dinNEWFq9Xr1wj7fE7fa3DzOf8ODL/2USp8zeYHVYwfSEB3IIiv
LxCAggJ+tu0Dz38cst7vyJFKKddd/ynlRqpALXlI/Cl4hOWbkkuasuFVYlKmOs5G
ESAzrkd0sMro8M0MlggiWamC7uGS7HQRv37ZYVogJGjisTcnLyVPnGwZlWX1hjiP
sazVz4JQGt/bmzhHdf5mdg6t2uznRVQwI/PBARoqYqc9kEpkKeIebf2NeVRHld4x
hhG6kcrBUwtbugDBFpysZf1pT4pOYS7+62tnnjAoAEqFOe7Hr/q8SwjlqNUVh7PQ
sBEa8FR+JHWgomiEBcKNTKIrFkBbX5LqFX/0mVQvQKV9eab7IGlNHfEXPGsecDae
LM+HwbqEp82NJeG8A0vldtzmF1I6CVpLa2bxKhXDewM7RAgjbuydMNP1ws0bcLRX
YgaZMzB7URoOr7/25UzXDLZwAmBpgbiMPjd9ZAq1NPsAL3oCkqwuXIm4ugBka+f0
rpu9VX65z/xPFYWXftXfrH7GBX1aYgUlws8vpkP9wNlXzimFgoBN2fhcrYzgsx9E
cXtZluyliaTCOs0a4fPvt6vTvK+GR92GkNVhlCQkJgoec3xxDTwkhh0+a3FLAGxG
uya7tc3BB+UpfSB5MpvNDxpaIS27R+glg+/x4CCUgDo1ZPiFo/tu2a3KPGQG+jVi
/Albk79v/90+wbXhwowZc1juZeyotXBCDhnBIk2PfoxmT0P9mO9QkcXPmAHBt/g5
3cTAfA4k5kIW2jdjlJlkuUl2QUnFOCwKXeeWIWmgdLRkv3bcaVAS+9Faqrrcihlh
i9waL4mS8cPbnyhGrYhVBIWJbPK9bGLlFJuwJgSMcxABe1287rHRbxqaJH9UBHLD
HgV00CNg63cDo6U2wA+dpiG1VlV1kegCgkS7UTu3+FfImToaZVnJRp4iPykcYy+E
WHe1zD82iL9fr62RPpnjMYdrWS6y56+T4w/lo42sKZAubV375Cj5DtNuoZ9FH29N
pvsBX9yCwCufUDwpLeGhkaOl2pM+qGivj3kSS5Yy/d66FcDFyiJUbevzX3k7j5OI
Nq25TeXUz1277YDwjXNpj26/kh9daSu9emDE14jFqsYDV9fulmoOKUq8vFRrT4h7
WmuK/noDv9NnYux5ffiXNZFxuglckFL3jNoxQ4ezPEKORfW/hQ7qdxULqCDgnNkv
s441LpBbiJntPXYhhW+Saf6+rk//5mXAe8MEgSaynMiE3kDMY0EHNhZz8kDgapwJ
TkiE2UNRYeulCy4eymITfVG208PAdsB99xEJR0pdcqp8fXAx5ITtKq71TnRPLfEt
z56AtuAKrWajhnncDQh7B1PdwOL/rprhHC573vmi6EVFeXK94DCT6ZlrCxGfGQrE
4X4GnfcABenqUU81W8xZAD7rXvaTofgzBv6oITb4hsmbd+hokO6+AQ+KifzC15o5
8885pP8nrgek92z03STYpa2HV+equOBbIAvglyP4pJv52+pb4R01qVT4M0ARoe2H
7Pg8wajpEZX9vU4JvJBDH2V6YVZlWjas/TJCdGN9PYbZG1bwOE+EJou2oJ9o/PZ8
r/IS7mwRzbMHPMqUHBNiAS5zLfV6MMVqiNYJuCL1AkDzEOlMQ3b5fPMuIjhOPWpK
31nJKgMu4PGPd+/JvZGYss2MxjdsGzR+MjdwHqaue7b5nzWTJCgPA8MqFpXTkzEg
l47LVLEdG+v7guzq9YkecIBp4V1boKLcGS8EWpLPuFgt7Y4B55ewFfjq8mQ4nopt
lfK9ZBq42SIFaU9ggdgA4aIkJMVFrRrooyp2IKC4XFqC+oD2R/ahYZCkG6tiMwfU
dW7dB73lEEnbo2pfX0Vy8dASG5ElwPBlywsva1LHpOXKdBUkXCLb0QDiUJEveCaZ
LMh9t3/txMUQtfr3MPl8oU/WQEAzZF2CFBn4wcAWXHYNsrGRXqrsA+zKjHL7/hDg
8auB5rjRPtiiKVtw7FZe/IddMHxX8hVzR6ZwyhtXI2w18iCWPJoIgv3AOqYJ2t33
nOcxWdsWnMF1wg62sSzrKQyB3gLRW50xgwcZB55CDexMH1APdGPc6zVWaMSYCfYw
kOD5iPOUUpy+8K7UEvFclOagKDgzsPInXW09TMJIord6pDt7gECeT0hrl8yrrcZA
zVvcu5JEj3XVy2r0FFrKAgexQtizbFJNfVsHIXZogKk8JGUcuORCKN539syLjppl
XeKcgv5rF0fVILX8XdVK9IY9DczcP6cOUhskGj2l08JKVuLRXqqfYHnqgUgoAxMf
j9xg59xEG+7IomOhm17g0jWF2Xch18pzDoaC6A7pp85XzL1GfCoCaMIuMr2QlhCP
L1A60G4wzI9tJTAOOeHywiMsoFww5wjVwuJdToIgcLsKJOdukNVlYHglAu97Xg8S
qhIHpJ43v/gaLHWEQ70A9LAP8VW04Pjwt80z3uJEcjdTWW4Hk+PdZc+q6Lww0J5T
Qpna32FGBUaMD11OAfA1Dp76K27dyePJ9uN0NxisOhZ5PqegsiojRLJs7yfeBu/a
eIUehBsw/IO9uJrr/V5Xkz/RWS2KKKGwsovegzsGhh1OqBvQkIfcfO1eBkwmVmZ+
wfDvAP2hDEEtXKO7IhhhEoSq9C0+vkwRVkm8mQAwDA5OCyBT42F1gDEE6zMAT/Ih
hU+AQFMtKCw3sxpDP96+IkxS2EMkWibFhY3Rsdn/nQs4FdeBLQpiN0CCMbcfFbfb
L2Y4KhKTYCy0AM13GUE+hDzW2dXEDT+5p2cZyeMiydDGqC0nECaKesRoYc5AJSW9
HggCk8wFsUJSqNmYNOuKZapgTzaJx9Ya9sj50qdtbPDN72fujuyrNODDnTNJ47xG
qbA/uiHGcOqiDLIWNKsGoe092mcUHlwWaWn+IPHc996TgsvoXlT5uJ+rovmKOQc/
vYrfAEZcBRDtcdSMS3Ja56BOtDBcdKdsyMf5yhAoKS6gfUV8VKYk5meuTXXwyRfN
ueSMNPd/SqZ204/NYtKwPQi6RWPnQJIbWnOkwF/Hn/HHh4G/oRCS3/GMLSfCeD2h
OxqUV17gFuVLSupw8+uoI8pA/UVJeoPzqApPMo3nadm3wJcQOho+B/L+By7pSFao
q0ucV+ubOcdhUr0jYH7PqmE/dW2PtUW5uyOflNYZfnsikLq8khQDmF/9ePiaw4Mr
P7w8602ebzxzyuELk+5x8ecSMGprCM/zY1nfh85Mqp0bolzCWetQ/LloSWzzz5WJ
37ZWQXMIA1pJdEp69biRBqsGtGERigbJZEPTO4Oo9wraUEWpkEp21DfUHx7CyNzf
r8JjGevpY36vYlwkfw1ABiMXl/l6VxblHFzRfCfTehqoqTR/T1HeJ6D62rLiF4ga
0zcCteDEM2byIpuICynm57dMI1Mcx1iiP+ZLRzSnZmmapyq5NE2TjRdKuLFVap3Y
iRrO8nUBVDFDd009NU756swfHflQ51z6kicDopy/IDkTgdzw4vYiiLwXjE7jx7yH
snCmlMhmqhU2ogPUtf4UT3yNEaNKe/ESGREkPHR6JN3FrLymVnB/7C+2jB1/Reks
uWLRHS9DaW2OUw2CHdpFR/Z5//NW9MTGC3/dOijkNbF52BpmpdHQUadoZ7S23vLY
GgUoSYCVlUphtC9OcMW6u2D5nWjEKy8yXbub0bfPr5SDYXFpLLbqEGK8GK8i6uvg
mfQnZHAz9iAgWj53QzeHoIEWqrYxiAWT6EEQwZf1bUJdtBPQqJtbedYWGOe7eVVa
imCFsXbAiVV6cBi0qNemxyfZGN4h9rPUP92MLE0nuq/QMW/w1pI3d5tZxRlPzh5m
PAjBW+xg+u2TpPxSNh1+8RGJPDv5QS6mWGJkP7/8p6tjunJhRa0B9VUuXguZORrV
5zN+gysJF1qS4OOekBio4F+FkmQ4IoxTw8fOt/Xus2cPiRcBdyHGXpzvkdbnmnqd
WFrQlezrTkRyYHRlIoXmhnnpbGFfia+syuJG27q2gy6pp/l9aap/IueywTskXmV9
TjChsF3jGA8yXoV7i01QJw70Ov19HJvQh5fZOA3k/CcHMEXFg6uz2FWkzSj5WQNb
O5xxC45XEZOIMEh0S/9O6jx4qaOf6oleIAzUECpJ4P+uJBDVSmLvwyRBWXGAfL7a
MCCT8XpWRs+IYI1QolBaSjWs7u3/xdW9gpZVlhG9lWdVipdErg72q2NezgTmjDlU
H/2fbfMQ9MTgbCZjV3zILcEOyLsLcD8xI+2+PO2wHxNyVamgC/UTngSdBk7cunJx
bCzVJn02HllaBmxg7IY6fQdUgqdxj4JPKoj095zEookyGmZ2VejV2Sq7AROFLOly
rXn0wd4cZdocoHITRqaUO5BlunLagUR6x9WJK03YAALqMlAvFUNW2fd1YPKTpwhf
jRaWu+cVl3+etnUwTS+qET+JUxekDknPjPZqgd9QkGPCx07P6DR7ZvW1AAAEC8+b
iNcdQTi8dvggCC7zXIiq4qMHfi959rnGF+mYYa23NmOQBDZTH5AV5xyqrP5QBxRv
K1+RzWlMejGfF29hOp4qHzqQG7EHqEmB0IbEU7dOYX9IoRq+6TlZk8c8gKhW4xKp
Pj4fkCTGnAw306KrWchPlzwfVTjUKvCRgDBx6x0coFocnNZUrf3lVkplkYFKAyqw
JCN1dYWpSTFUNam+4BtcyS8+e/XqdHCQHSwdE16ZkBsmmHK/prlJgG3VEqxas5pY
Nblj1iHmrNVRBnCTY2ah5r+08ufAKOpF5s7sAtNsnw20aOoZerTTCkvX1YtrB6vp
pQqMWqH+38nk4xGMSpWSMBT9Gcm0qF5EZWJUV3Hi4AhG8flSD2Dn1lgA4OlzrPYk
WqdbOxLZ8CMjrWThdQBkzoBttIM0DuPODLPtz7SbCcg+Xs7IXCLxzSRFCHWV5qbb
1Srektv2nhRQmMIVeoN9AAW7vjFg3LVCCQZ173fISLU88WN7rmHqOOr4m40yrf7l
t6SEU2xDXDPLT3D3v0beWvYNCjWGbgklKUAzGt/ymwzZtb8wEiaVKgtP7pD+KqaC
K0C47IPIalbpblnEOVb1nuFxB382fSSop+JdoN+MvPBPUrbEMBEIUCVo+hBYg+v3
y7x4VfZN5+vWCR6/6PBpNRHfZ5Gfo17wAYk9t9GeNO2BGBI5AS8yp+hTW57eNJvM
/4HqdmORT1R9INWFbVlA8eFlqP8e4nOZ2SkAmz//RePMp1G0ehUwHjSUnTrVu07e
OpcDx+RxZic07MgCfH7f7vF2p4WjL/THqgMP46nNVlR9ZrIsU7KLjrd05LeijunU
Kld6IqF310fKKHYFfII/Ivb2RPTnhaHVTKl6Bt/KHOExxGQFNkUSD3SGXdtHCvVK
6dU2lMg8Ko0Ieo9NmGnDFUZUVAFxEMvq9pAtsQxcqPW23HtOYQHACQ7qv2QCWS4P
8Gf3Ddl03CSjsk/XfnVqDr3MUXQxmOnPu9mncFnnhdZhXHHLFn2GNByOqru/alxH
tkD/+fC1+BUcuM0pY8n1ito7oJyTqzDV0Mc4R+9gDbjAFcxS9RO1Wt6jE9RJn5eY
48XifcLLrbFW96nApHl1srJjxLcyXTTw8asV6XkSTNbsYBIhvJ/xoQhl+UdbA9y4
J3Pn9jGaaLXX/BI33KKYeGa3pKJnlSMYTR7lQYa7umgZjj+d0yVgfJHQVNn9EIFd
PYfE8FxUsnyVWj2msFCZCrnbBwDwW82WG60Bg12kT4BF3BEIN3yX2z3JnDOGUfFa
ozORuoFeU6Pr+AlLJFycAggBKK2hAfL1SoJMFpCKeX2xl/8jz56OFNOGlUPjKAN/
c608dPurJIZg45GE0x0exnhaqJM2v4yTE9CJkW6yRBNpFp5OySUO0jbwwjLJmAHK
o5YSI8riTkr+S0lAdl9LtGyRbuztuLyJEwJHLMynYj24uo1RRdb+7Sb586Nxx8MU
a3gk7xYc7Y/us20y+0lTGJvSUgOlevoAmkj8/f3sZka6CSXLoGnlQ1w3PdJ4sExt
YsomQw1oblE4gIeQ+Fx3T/sB5HxdKbDsU5R9PsVYF+ZdbD7ggtlW6KNgsCdOlLCJ
kF7Le9hs45TZgd1Pmb2/5aWDmDQQfTQwhvX37Uxx1q1cFJRrR5kdr3lBBie612VF
AiDTaRIxgxJDNfsF5CHmWWprrC9meCelfqPbYlEuJ7/DA8hSEF6YY26OSt9pYBcn
TIwXi4Lwld3en/tfZLe3UvMkcpwOUO6oA1OIy3201ciMMvL++/rRIeA/o753FErZ
t93KVasw66CDRiUQrHkYaFZy0WN2mXTXf79xP5OjZ6eYcFOuBAEka4v6UCrGZm+R
q4ZtwIEO/SlXnuQAadTZ12evqs/mmg/v0+nxrnuweU5RTJjnM9FZ5/Qbkf+t3Q9o
dWpKaeuvG3Fupj9Hufe84HeCvM62KOJ0A59Is6e9V72ub2g7lyn/gU6dd9bmUEBf
XNhvI6UzCvq03dYDoxmoyl8ib4rOebyslJNcPuebexmyT7/XkVuMs9VI+mUHAhOz
lBTbjzXFBmLuyC+3mKl1+Ds18bAgLhexmOXTtM6aSJFMELirDBDVxkbJ8+YKkY/m
YJ2n9O+lqN07O8yDDybiO/1GUac/IJer8wXPMXArdglRdd67wnGJJwijMzchN16y
7L8/r9QIWFvOrzVft8bKNGYo+fc7hFTLDxH57GdpVhdXCOnEOS15JjvMYwGwVwcA
Iwi3ZFkZCehWYXJXXYoqyFK1X19gWSCAxPPKb8BUC8BUG3wRlaQiwBA1oyejeLmy
tmfY8Po2niL9WsvWUBhnQH//N10jSqcZANo6WqVf68jnoOEoCofE1Me/5LHUDPHR
9Mf5VAVBnitEHP5EM4VmY/HNbZBWLSVZUL1tDPGUnqYsHVHk0pzKr6R2HK2xWej/
p/bY6HNBJiexA5TOkHQOofQEZD1dLpUP2uww6Ts/lPTEMDiHQiC1BDLl2yCNgeaI
OXazeM8GaZZ4PRqNT8FSz7QhLd3w3NUJpI4a+R6fvKbDwLJDndlbQ3dpy0WkSJQe
IppJxEJdlz2HuU3TTCytyiQhrcC2NunaVYrJZ13klz6Xc/Pv1xlApbXNIdyKU8IT
p6bbpSYkb629qgcnIszPRSuHz5vWMOMbtGB4LBmiDPtR2IWBjbnmQCN6jkbpdYlQ
WAsoiMFDlqsYtixeFfb5cZijN+CcNuXrypiLGHmss7dMDeMgPGjJC3fEuBWL2Lwk
o6RRqv14gwUMBpOHXNDUARQN/mKQiOcN7guQGqUEeA0onqjxH6IXg6/ygudfxplO
3EKV5qshMDx7C8TM1F+wREEAvSylmUKTOqvC1KZb6coiyzHW4bJtlHpPIku6w+Jp
5XwfOMrN6ugsKlkWLYHj1Aw+niI5F9x4BHd0LTD7LpRkarW3Rqahm9LAT/gO1FzC
oIC/ZZhoHgGygdIy1hBtlwLWSkBw3TZI7EdWst5MDtXBjuUdKaIL8Ukm6dQap9P7
/it2yqJtCWtKbuOPbQyZH4CZZG8ai+LSbJZKfmaKV+JlW/ol7P25RjSa1Niuv0vy
EmPQ9tmTAlFLRYSa0lf3T1yPhp0b6S5bDbg6jRpofVMugfxzIwQ7N4Pr+PZK4wBb
ATpMosIgYKW3N4CTMU43Uhc9iuPGRLNJ9z+0sK5etbdEX9sL89CCuowClcYzOCbD
5n1FuERCZe/jDsdiBkda+5dAHAtEfuw7o86IJGKzjrRddUzYO/y4SM8kurLAzFvF
wWzdCgRmKZ3P15Lv4s4jIwCbDlOTuZnS7ivtXve12yeJaC1Y+oVKzlO6OLzp7ezL
MYoLFOCbjvWamFXF6fwTDq+K/m2FhSuYq8Q4xuy4JaFljmm2JsP3L9csqIe7ak9T
/BPPwWjf1YvlF8a6/Lu5oztwwR3DMrNExIKN4N9R8fUogosxS2eRRmw2KTdzF0ux
UC3pXMGdQAkacxhId6MA2725rL8QjlHmrEQK9a0WbHLS6HGR5tBkSDc0kZTbfvtq
e6xjqmNydT+oDe9bfCj/jasE7DTyNtVvrNNYKiRcU4JNsLw+OFvNrZDLrH+ik/RZ
BD/2dTZHMHrYUZVL2ZZqbgrRzTn7KZFDaYr42LxhPu6pFutkk/CPmeTCmrDLhLCB
IbxbAHDY1HYwoSQmDDMUHv5WHjhLOYHv2VR0waZnGEykRMXO/EibxkNCH9eEjVic
WAW5q22AMG/TpnZk/0tlyjnnOTm/iRwbAv80OJsG5H284QSJUkmDhUjMRF3m8wWU
/pCTm0wsaUeKYYuRla3qBgxeaPU/c7kYni+VuMoKkNhUOc/KbVZu53l0t6vLKPUE
1a4H6liFAM2/cANtFLUXqqWIag9psCpQ+F9977uChLHyN2HMbsw11PfqQiCFFhn2
hFG1f3Irr79cgEnMYDfZwvzYNJqd58zEicEnbKn4qcZwVePLR/e0qP6cmk3cGlM1
nNZp8VuMVnTb3zfjdg3Q6WaZa3e68wJYUfN5UTMsc/zfw3NPV6y/zdFi3k6KgYs9
lYjYJAY4wKsNXYYl2h32n2beiZ4lpZ6u2eN7Bj+dmhLJ45POI4i+8Yy2GnmlcE2m
3/Zv895B9Q3hXbY9pOvSSVDT5kvFCxblmjELWyshECmkeKxFU1hJ7q2hskQWtwym
snL7NEGwlro/PjuXElhbUqf/tZLsFBoCxYT47KaRkUN80Wzip+pX6Zbt1j6GusU7
J0kFaQ2+pLKRCGR+xiOah8rVZDiicrcJLv5VKKQStlCjSOEDxOeosNXANU/gjPhO
S2Bpa5fE/M2i+pCUEmmkhwXFiu+DPVsRdo89vGbs6QQUDBGr/rdL5w4lfRDnXvKb
jyVTK/I4AAhQVpT3Uw9I7gAo5Nbz5Bksg97ydvPjLbEospLZRRWJl3HKz4n6ZMca
UcbrQqsKVw+UG8xvGb4RZDnzGWk3AFa5PEDKFQEplvCSVdikVdLwY0ddmAe2CpTx
YPhAjlSZI2Nm4u6HebZLjvMMFwLLKEqCKhINMZkzEl2R9RvAYrxC3fodAj3hQQKe
iPAlpGqgGjQ9yAx2/qdLFesM1WYpJHl3pJZ35riqftDdVTgYJynhgDpl8TrfVP4c
vzwtDeGhCe1ONij1NidYekM4t3PudE+VxgOAiJGeAggMRL8pil2mC04D38qPDYAb
keTFK+1RT3X+H5bZ8E/8WyAmgmQo21GnVZx3fQlKLT5bknOBoL5AEBdJklVVJz1Y
kn612IorHgsAoR0T6I1/Swvj/SUdv3SoLuvZ2GwyXEabvXPvGgt4KYLmrZrkhpMA
MbVbvfabdqt75nClWcaa/Bo3MbqHz+BPFtXt7mk5h/ZzeWdMHB0M+UFmqAWFKF8X
xD2/h+pSYjCVMd5WMT+d4PJKL/TKJesJMUt2ppLa98UXdMvscZoTq61tx9pTQfMU
rcDWdDpyGdcpD+CAPaHvthsY/H5JmWxOWBdlwTvgKUZBiOMEvhYfeswByvkKIVwz
2/ldUB3HtcztK9veb2jmRTRLE5fkmriTqgPyxHWyWZaJl/gLUyWpaN1QdLlz5sUJ
vTaFfQ+lUhErb+ONSRbMdVuQXM3nbagyoMae08AK+fhvNBPAo0muGtCAyoEU6yl6
kH+gbE3mqU2yv2cLO1TeLVrOInJULMgfp6k8pGxoJwYmpfo4JO44H5YnKfYl5oYX
mjmd/MJ7MPDadEBbDGBZBcgf1feKU3GDMjbeb3+v/DbAKeKNcYbz262ehFRTEIGq
kEYyLtc8p7l0QtjqH/iBIWfIeAJEY4vC1qaMhAt+TXZ5nhLs6Wh58FJH0DILVU1H
Yz2eLaL/vnUG8/iXId64d+EL9zzAYWDyIZb9PL01l27NBimDOXd36GMuXNlK+8RF
pS0qYWKzattIxcBblI7sP1JYXkpa3B9+KPyzncueeDGlaJdJjOv1TAUG/5DLmJPO
lNYfWr9Q/7wsrqE4rTN6C8WcwpoW/rrGc3X6sYFC36sFSg9C3WQGxD8haTU4JCvE
15hO8w0bMC9+gKJMbnMs5vmMVQVqO7jd4rvWF3bsZodUc7rVj2SXGq+hbaIQDvBF
mnIfT2QcCLZn/vEJ6a3FkyUuzl3D1M/ifUCAJDHeeAuShyCI65ezouE/W1drrPra
ltZ6Wnd+GaxkIAZQfdFL2iDpp8lxGSDNQXuG0m5A4A4+7LftXGKALg+n1boEa2lZ
AU1CGgdqoP9zSFIA8+4F7v63+ghVJHRSe2/PRYB918+ByyOcl3ZJHTv2hYYgrCou
D/q/II1Wz/5M74hsCwubTqq2i8vJwCQ4N/LMEF6/A8hRuNR8tsle21V56kbfyCYw
0Wfy5ZIKUau0mSmokf7LAM3kzz2NrxJB5mFeWIfU80Fe20pKDDLrNxx+SHdAH4dv
ecjNE+2Ts+vMmiyZdWvp09d9bQsrTl08dcATI0749LK8eumqO5krJ9aMsLettWTq
LHTezj1Q7rLF8n0tbdu/l+TOSBq5wZj/7BfiBas16dbKZQZRBGtSwy2A3XWR8+rC
DZoCIXgIgbMRJFSXcDV6Z6E4k345KF+TMRd6uaR9sf1W26aXnHdEOIMWUYxnWrdH
sPMkEWHOyzpvgtljJ2a48Wg1Hdl4P72fQW0DGjsohlnhG4pF2DDJjHptLh1DfKeU
SRZ7hsKNenmIBBwoLmNcRqB+LsNNuznEFi1f8PtqOG+Pm6zJeORzYr4Vnii9JuaU
dj1ki0d8mqXEM9tfUS41ykqjEKkCRHOaylvNKSXbTuRnyo5AOZGpjyjWpf5z7zlx
R+Bimlpyn8Ey+OiwWyVez2B3CLELNdsXWuD8qLOd4xFPH6X+y2rtcXBiuqyf8CbS
9TF4CsJn2n1eU0ueAdT9ocndDCl/eL2qNCTCj/u8cIugq80r4QAQJ3KPyEbzxlQG
okW86xgSgXMlahZ/BDgwnpXirbW1Anr/cWcQAW3hjT6hJdrhZKDxCNeRwmBXu0le
seYGsq6ctZCvCkhi93Wx9rHz220AL3TJCU98Ni1J8IGN9NbbbUwt2r140h3XJg/t
2P45XPwQUt/ARqhdAwHujE/cGbzVqxCd0Y5t9nRd2OW6A3BAp6Us8DhngCNr/FIO
RzSmLno/jmNiAk8U7LRaArzGky+1qiN7nlWr31Xun3ixvKtUanPx+ZCrgSW9rXSk
oyyjHWOCkxqlaWPh3vJsBNA+FEAtjB9AASoR3D1KnMpk2+RUTrnw/zH99xQ+M+rb
wRS9vMkwZKkUlrQNPtLDt7AU7WmnH/lOupf2O6Y9fj3KbPTiRvV5jly01alqqF8H
Yw6xhaHK3ZlvD7yGc/ZxiZPFcnMDIH01Gyo9g/HhWwLNNkJcbhgRjUFK/ncMGYGn
wUISjbUYoUhuxRaTc458AoGGdjSDol1htbLDhF8YTL0K9dAiub/3L42ud48nldrV
BfXhD5f7IrTKWy67iwk2T8m3wotBYZmqjh2E7ROQA7nHba7tzxEiSZLG+AFhK07C
2xUKj41z/66eo6FesDfS3meXxl2xZ49NN2t+6QEOjXCuhrPQQxE/xAYpwrfL3Mhj
5gXUyggmQfLNfub11NydCWHjfgKOnPkOUrTSG3sbsPHqHpm3nIuxUm9Q1SyB/cov
RbMaM2F19EuSif7VlLV3pkGWOTiRTe6RHz1UkSpLIIFO9tqt3cqeQaeOtW3XSwIF
cTz+uPOpkXh+yPYMpJJzbJYTulG4tiAfv1lghmX8xug6XnjYli/hfJGyUrGg1pQN
EssrMhy0XOZcozLR4a73JyPnQ6197vy8ByVI5wC9v70z0ibtSzVmg+INQKHuTr6+
X0zB5mc1CqDH+IdCObk5avn54q7JoIX0vUVkCjhk72VrRFSFY29F5sIreMmSyE81
P7MmRId/09x1DFk64njiASTkf6bYTisZvjwo3czSjkvSv12Ka+z9kdCTE/2g2NWI
he7Znl4TONzpvBJb8sU8DwirTFu+d8fiFYyaZvKjZMbfAKeESIineX1D2N9Pb9se
xYi+aetVd4mTbjliAcgFoUTuJrD9vODxSGzbuHv6y7iwnW1Iirn+Nw+/v0oNysKZ
EE2ucn+rIBK8/5q4vPGylyIW0ZkB1g4HTaGeKm28mSs9S4MYtT1Em5X7eDksmNE1
g8aStnXRpb/C7V5zf0oi5EjmRBRpPSjaVMpDE30mTuSYJwlLhaexeSmmEZh3j5DA
FlVyhYJHW3aPZ5K4p86fqn9LCWjlyrs363ae3NnU0ocRrb8Fpy/EkautGZ9Xoj9T
jyY35HP43Yfkdi/ApfT8UbcCmgowd+b9NZdFAICax29vdka3lapdi+oQQHCAzkoe
BwJja7HusnGSLm62dgG6Jnxgwdqx60Q6uFUlTgRwjp2TXdfzsK5wMHLMCbrHMtX0
M1c6k+GVOAuitG8gBKA4S6+gxzJ4AEMJTb1t8Dbc/Rd5ZJyIS8PHeTIaTrkSVVLG
gJxMnkbgQH0NzTosiVdJ09qy5VhMQXXw6hN0Jb3PhFEB+Su0H+Ngu0VuYRtJn5XT
sbV8HacgYtWkyk2uxbPZF6k8Q/1ewQ0WNZKhfws/IIaI3XWJn89YOFa8NQk2tXAO
gEpc5k2iLc4hh/GZlqUXeRza010iCvlON9Na+C+LM9z7zZ7hFGnNqzZ4xhR+eAWM
vV3oTpT8YSXZ3YR1F34OvwvzcInSWnGueq/fDcJhiN/g3C4Ksv551BIbWl7MCJg9
+JF1lGEoVqqM6GsUCrhiuj0P7FWxC1E/8uchCu0lhdZn3hbyDy57jxLVpZVh0Yoy
POFLYT2xOjWeCH2oMqqvl9/JPLRiUT5tX1JYHzCgVe6AmOhRDzn3Gto0G0uIx5ff
KCb/GQQ5f/qYZyR0j0UffWoW7dj4DYhrxz+s3ZB+gJVm6LoS24oyDbMn5KzS0+wc
3u3bbhl4z1pHjjNxe+BCJFHl4JGiwqrWJDYovFe7j6kjPDyoOsVUXXaYIYzoMSXI
nuTanycPDIA2btPFTsMfynuxoBzg5M5C5eN6fSINtn6U0igdYztYR8l9YritcDGQ
YIhgoezla4P9UtMOLJ3wqfVIeiquraArmZLxoYS5fBBAH3JjzWKvFtFGfpcgU+zl
BfhkdDmXxarE7zgnh7a4xqgWcCH7V4s6C9F3uX2wivNmsAf1s/bD4Ib3timA5z3S
q0GA2y1y2VuurL6WdMs3dnaPPHbEMzlLI+f6wHPXutAQ8oRYQYJgst4IUDX1pbw1
dJ4sPNmhFDcuHReQC/D/bILQ8y/cQGKPcst5qsmQ4wGpVhNZEaKzLtMQcj5v916R
3+TegMZkPAS3FBTvYfZrSP4ZAmMljsjEIbY03akIUUBjJClG5LadEFjE1eKFM10v
ee5wlQw+VORJJb7GF3K9BhWG+IfZsn4uWPkJGva/OmWpaxF+se55AXOyidZtbBsQ
1HCsDEZpuLafSlXx1/4dKmnDowSqhCRa6QBvzj3xFgcEpJMRscTj+qgyU5biFW7B
fNJdNzBwwOQ1GE4HEUjgK9e0d6OusfnbOH0OXadsIbUzv/m6QR7keHK78OPO2ggT
1HjaV94vTwl7SRYqJqw0iZzFWPisZzYvAzhlDeyD555bHs5MZ3GcdYCa1kIrE0OF
zgBEIJbS/aGUE5wIBNh8uhrdMVY0U9AtQChVyk3ANBvD8/B1ld44xdKSjZ16iwZj
FEStKUZ5B5G6r0jdcHFd0+DZFi2ESAxs/vjQ4oUpioF00l5/e2VW1rCfIZH4Wvm7
njF2mwhMpQgxxR1PRxKj2M877G4CKJi7HxTMeH4eAlecNkWezSrGzpPKWmJ+nPc3
93rQ9XnoSrck8ip5QqZQ2FmDiFJUkCY/kHVQ5pN2BoxY6PT2IDGYaPs3gDumtepk
+sC1qNojJaoKD2nPGOuN4zOdZMntKqeEUAbm+aDv36P4Uv5ZT5g3csdf6du513p5
vAcCqvF57H3uMLqz9Y7RLL9sqLWiY5SDgyfrAEIfro+uXo/J7KsRbJ21Mfc19+3G
nv9ZBLxAbqYoKrYTjMGQJEGEyA2RoenCQnx2cOQi3+ljzd8Y/kGyCYri994RrOGq
AjaPzr0WK0/gM5RD5yYzSa2zVZ2iCK9c++LjMcIYxQy3btXMKCBT/JihImTouyXN
cuw5V5Oax/x0VB4KaGityD4+ZNIdwvuog6PIqskJO7Gj+TrVrcoYZOW4oHcmLtMl
RBmI3ve2EMaNgnUM3fUD/Ow7tfV7aC6lLSf906NnvWuuumdW5IHVE3YEtknogATi
QHvGI7lfnsx6QHXGtNiVUscWHZcXBsMGbYqZs6nynRoKfJMR6wIAEWs3RuBXp/tv
R49sP6gx5icbBTovrIpI/IgS+mXThAyZJsJSXHYGed97NxuohrXdoujs+Uc6MzSU
+va3jf5kUSDLHALceYc2SkxVfqJmYf8sLTZTZ2qgowV7O0j4U2diKPxdoWdbeY82
jrqk0aW0tni51isZIOT8IBcmnnBWy+Q3IYNBKI9BDxqdoUvGAI8W1VECzBw4jvFP
lzB9UwdFCAPBe0WKCMThqFSxYvtI5IUAqJfTN1YmSD2krJEQG5+B/Ft26+B+H4Wt
Hd6w210Qe8+CdBa4ZpiRTI5jCeCZ2kQBIayBYVhvKEuw2udiRaHkAKQj2Wq+JqHR
Fm24tQpYwnU0tU+GqOlpRg0DoErLznQ2L8yopOt9JCoPOV/d2rMpjaKr7RGLhjr5
Syob8K3hQUqQxk6KIAcY4wcFOgEYzuEqBu1Nzvxyu5a4Y9XF3nFjooXbhNLU4O5a
n2Tmv9Nh5fK7QCP7v8DnyqX8hCn/Ky8DtCYHjSf5nlPhM4nZ4VqHAjDRrvJLxCZ8
jRlbi0WpPbWtZHHIa5qW4ER7w/0QxmpHP97NXFDc4j9cbUubsvLIfSCZD81SJ3uE
M4/Ezc+jzOvTw47xrpYGGiMUjGzds06qZrDh0OFI6GehdWBenKYOWVdI1QCIUm2+
iwF1SCw0vkNDfh81+0wZTA9orPZAO9Bit+ppYscuOlgUk/H6VUbjdlZfJu0LQBSF
1IEqx5sIuee2Ud6mMhhlTjFgE14o2PKf3W283EIPi2dDe0UIDwaDYznMyAV2ZOGL
h2jlXc9Yqyjvw7ciUkuAPJZG8nwH2Xzyhw68jmB975LiTNLytN1+q5aSZSYgvWjU
rxHwOGy1vHOYodXAmD4dj8xz6ZvR6uzgf/HE/iU/qBpn8pWdWKzz8xkt8iVI3on8
lzu9bm2rn036lSCmZqY6qkZq6LYEj1eYUhSq7el+Npx/vtLHq96dQvUl4wKdQf5i
ILuZoviMmkpoFENZgfjzq/3gppdf48wjKLD0y6B13JS1L83QTpXolghOdgWlnyjX
XYCgYYtqbUmcRWWQOfjPsL/QHtry4qYYlAlmLb7R9BJlKgXMpiBrLgSGae0sPtSg
WRU332eFeqx2yQ612rGQZo/r0F0RKUsOGFBeH4tSeKCX/2aS+tSzFe1IIE9syvU7
8nMc5UDcrdgGnn/6USjdI2vsQMgL3ocx5/XGZ2mvXo7ommyCyrE8SWWt/mRfRyUG
B90LDxlvamnPtvmke+ugTRuUsN1iv5ZYk6j5aAqH01vyjr7zD0XBZyLeX5lNaTbH
bpqC0OfFQ5aEOnMl1V/minXfvY8xA3BS4gOb25c0Ujxv5vsITZHP/xz3Og504U89
YJI58ifRW4K24Hy1Ceqz0KNoC7M+aZ82TgMxw3qazTJNvAyi1g6r0hsU1JN6PVkP
f8BPvgA25BjTDGMteD7/JWrxu9lRohI5EB4S5JhFmy930yJiOh1WUikF9HFkni8C
HW6sMhGc9LHpusPsfh9FLp86CXhmZKr8K1iy5yVLZq6sGzxRP5/aHfR27173R3A7
wAs05k4EESzTOn0zhA72eODShf387k5WJwZQ7cQeyYK/mBTE4VUagTVik+m6crnk
1TM/y4WJGYKtmM1zSta8c7Rg2LgWDxJmp8v2vWDMRlQJMj9KNXhdGUO9I2RIqiWs
bMyUsYGqb6RZQIeo1rogi/INEPkwGDNMYZf/tcjrR+ElgjWgsiyWswQH1gwaHNHc
AXvfKlkKNPoksYDRGATIzp39v5U/WRbOioMoCwzFFhFeORAB+CAiLz9xYcc1Y4zx
wlTYgmhXNcUMryLWBYgWxZqFoZBNUGtqGoorESLHcowC0kwpFCF6dHjVKxUUpe5y
jzcrg7j4FVIfp8DQS4Lba7r2DuJEjYKu32oY2ZMPr3Z9fpBdNYpfouAkmBMWxwTK
NSeQFy59pF9R+i/1w7J5Z78F0ZanTmY81VcYOI05kcp1m/eRI/vojaZsZ5sUN5My
E37jrug/BeQ0c/W2wQKLlTeLhUyr7K5ycEJVa8Cvki6RYM+1kr/bHmS89ZpCTbc9
H5yxUGvXfk7bsoiD+9mXMdjpEYrUSvlWybkTpqKrhkkgh31pPQucmEzyMygG6V07
L0CGyFTfxDiUGKg14h3xpO+MTWRXNMaLJzwpI+7EBPOcLhWrVAF6wxlm6bwW37U9
AOFUbA3XKfBJuiGj73+k+6HL1or6nYfBk5EqoVJDF/tXt8msatZUlBxaa2Vw7Inm
OracRnMua5NGl1NMhlJfqvt7Fc6p1LrWCGXtxnkesdTqanrmC/jJ512Nk6Vv+sc9
thgPwCDAHPMoOb0ri8e43NeojhYtMCS30bMHcwCQmGw76hqm58OP3IJoIcXVuOb5
uCjwyBhKi0HaNavQz7cRDd+PiwYNtMCU00j+FjchPtYg8RDiTbl+9RIxMP/9T2yJ
y35THRY3AwfRI5X9VpbduznbqY9Mqaxf1zLxlLc1P3mf1T2IkgqLl6jnpakkg6m4
QiIIVwGfd325LqtjMKBLYJlvcavb2TNOzhfVFt+R0rp13Xjej9xJdCQ5rsuaFDZ+
Ul0O4LotyJmBu2Kd5Tzc+0Hgi/qSktZB46Suv16d481alEhlElfHDDnrjyXegaOo
n1OTMV5rPGkAwaexJL34OzO1P8oGltRb/pC2LRSKu0BVHr/DTWJxiHlp7woNxoLC
1AcLCaePLwIZS3ZbTklnS3D3zeALXIDr6otL27FOr2UU+w2mjFHDh5V9I1NQoOBx
jHwB4+YtzJ1gHHEmxUYrSTZyw2jBUk57xHPfdqsjRy6GUJ5gSelbNyp8tVVFi107
Lb7zcFhh+OpBWMICBgrkKtX1WkzCeJUDsRG5sIRjBsOVZh3QsCuom59sT1vfPPHb
8NL03XQcgCSsrMm0keMsINl+pdBMkqV1JDa4hzW78VwoJw5PWEo/L20iAYsqQOF3
Sd7nSVRD5Gtl923zI+SPK0aJJ14FCMi9FhJAi1r2w/stJ6IS3x+NdqvK9UVMOKxU
SUkqfjvuXboKJhnR0Ro3TdgeFqsKNlbcKpiw2DqYMntqjz9Rp7+c2lOt2M87aBTd
Kt8FuTbOuet150tPo1Q51VJGLicVj2vHQbMD0db042DH3+zYffPAUHlFWIBADA5K
+WHgVEoQzU/0H9a1ArnjQcz0jv+hGUbekxG2LVOPLcLbJ8IfHJchI2VcoOLrhzrl
IhRqmGTFqEJR/y0nowq7eeMxN8wl7rzK+HQ8xCjnsaSheU10TTm/khXzC6NflT8R
/M56qNQyRD7vh+gPwk5rL3u5X9SDOwDZ9m+fJCy4Z5W08cIvf5J2soZ8aSw6OZEb
g1YjjNJRYuAm7RgJ2yfUsEJVrlXK26JG3ZMpoQOw5XucqyrVBkc5O2laoQIW90O3
55gYfKzskJeEiy2uWT6iEa5Cdq4nOIfvrLozaeSYsdcB5TmVRUond13AT5htbSpq
K08YJ5t7KBJj/jDxtFOot5JysuB+DZdfeaYNBF22fgIVDuBEpbgADrdLHUtzZyRb
QB+AUqdhKLkD4H3gDuo9E0lJ+ou4Tbt0CCKe0jkYdUVqZ1AIFDjNbR0hM04VXSQC
H/VRjlsxY78Sm/szY9YkJALZSG5ZGW+J8168ziTz+RW70UVgoxLikUE6sI06YUh3
vpiBarJZl8BMaiSNb2E3lm0Nm9vmNcZGPmMBFuDTQkzQbYfF7TsnFsVnvuDOCEHq
8sGg18rxYBFIeWdVdmdlvtWrVsMDbSHD1UXh2hBh8DVTgmwZ3EtlZxWEA20YkyGj
xAQSr85l8kQn/Z5hDg+wJG+b5qm9wCqngdpL2rrQKZZwnbhVVmJc6ejxD7AM9oEF
932Cs+uI998aiWggE8zIqBHXmNE4VqcjjPlODnMriI4Ya0GiPpVAEfHyjEeZlr9t
Xwwp+ZqHmwck8bOrQUeFvq51JMX1ZaZOYAiLZ12TbFTafo2uPfOBiQ1RiyIjAF7o
zlMcN20KwFwCR8Gwv9Wh/f5/Utk7ecr8rXAxSr/chngH88ymZKY7P7hH54SoSaTV
qRnQZyk2+RTVhouk0giX+S2gWO348TMhf73gKJ9Wabq6yOH0g2Vj0UiZox0jRXG/
GfA3GQMXHsVeLS+X7hew3kx3vGVr3v3RcTsOvnHmJMpPUKIXd4m5IQuWzH3cNY/0
3Kvch7+P1m/t+c77VFbFPg08DsmL6Acbp3RogwqOVEpObfiKOcdkexEUrcyuLgRf
yxh5ZkZrL+q6C2iY8kFW6mv+H/lwaOmkSVWTYg+wRRr/BDcJ2VKddm0NOSD8z05o
5ZyciG7kexzeMs9ll2oWgiUn5awfUgSHVPB5Y45OKZJgtQEsxfZavQNHcDTay8+g
goWz5VSzWy2lwH8lOuLUuxIoJAG9mWThYN/2uAvEAX+v+KVfJptuzBPUShYitcRl
rb5mrwlCK5JABemPd/0KrWFvraJEUfLMutJUG4YgK4OFDhPIl6w6iHhQdY9O0p1y
+2jL9e5elhD5TccqIJY7Wya99ImAj4fQ+kJyX/iejrSPt9BoH4IJZZFdQrPcQozM
hTPs1Qd3Q97JV5GgRRkXKxTV2NYvZge8LRk44a3y2j7NfEB8EIejR/f2r7GfgGGz
NBOKYzEkcoDPGRKt2G/iolX9X+dqXVAHKshzHQAtQhUs6vjOzZlb/3swiWP8BWNo
zZtV6mUrzDvtSRwI1XJBhmX0v83gOj92glCHZ3mho6C6oAtFjz7GSpSulHsC9txN
IcNjSfGtpDxLGW5xTnaYEj3tFCSManMu55wK6N+Q1gVr6PO0cXk5q6wePqTvjXC9
mEjhH40/WiwS/ZbGQZoSmZgHaeaokJkzJPIo4xSHMRjCwwc3egOawtPQH0U9dOlH
Tmuwg5YQQWBNeKXixU8rqALT4Se2zWQDiBxHGTHHaQbAS2aGmoGWWfPQ+x/T48Xw
VpAXaOpC6NE96e2PA7jk26e5+QX8oHxoVf59oG/rlvOiqXkGXcAIULn0E25boxSr
6sHDiHTltK1junb/bixzjxFLgmd1WDOoFyL5ZbZxkLTB23JU2Yxguddgc4JwABst
WPvhw2Si3nQGFoUo8JIMgQN+fUuQxL/LgZPbQWfSBfbJbdxGXXvZQScADkVyP/hc
1aw6yHn4Mh7mFuRK9N1K9sg96Uzbovmp2k6w6PCOXAdAR2FRyX5wCf5vg285Xash
Vk7jVgJ1fRhGqLZwgXxFuS8fz2gzE0p5s6MXUvr69RISyx2xQX8RcwNewJA9Fwd5
Mxa+OQBCijtzAtd9JAnZS28DBVegBi4nN2CF8jNdZECERWzfrTuhUlLWSo3mToE+
TeaatvJGvTGu38b99ailul1dEfhmT2NcgDOIIQHMruPBH2mCqZDyT5iR0S3lXuAD
G9YufNoWv/e9iOeC6bYydSTmwHn30w+va58iAEzX/OUrJJcZgAgDQBZrQe2pT6no
xFUY0xNrJYVi+0rk5HbAux28VeiHnFGISXtiWJ5Hcp2f6rvxiIU3Iu9/dmQllrs6
J9ZL6g2/4rbiz9viX2Vz2ofu65eIPWrPt0xfsJzCkxgrUD3tkpHYZC/LIdHMLKCm
YasfHBSXc2KyqqSV7GxFcMiUQxijyVUQCuHVHv/iclTqxM2LYipfoMACg9xSFeHg
u+pPEreYD3uB/DVTcgaCAAqSBBoZ25Mx/zy6Ui+pBL4MWPDUpEvCcbXQLMEjNYz4
T+0VYcot5rQCuSgDiIy/EQunNTXzabaFH9L/4QdA3dpK3X8vtbaTy8w49Y7mYGFt
KpQ/rwgJa6aFn+HTFTsuKj2vy2t40xfNxRoRtVDRRz323VwxMdZdnDQrreXwgMxk
LgTao6BIU6R9hLGenQaaVEdAwsNPDaDDBLz106fFKzOeVymEjLphYUKpVchO6hHE
4f511ax82P2A2KiZomuSG6SEWQg4p4baB6fygSb1TFXbxxKkYEnuIzTLwZfJJ2sM
C0VR7MUO7pz2s+Z4U+EH2MsaELXwYYHRjaS0mslfLUiVjP79UMAZJzmoU2WLYxQ7
sRYgIqI8Vq27cGxv3XgmNR1KMyiZNA67E/b3S0iEkM5ALQocdgPeKDQAeAjvEypn
tZ1+9mKCQoLBw/5PKcv53Lde7Rkn0/om++ytIDXVRpYu/gok9Ck+IScdugXL6o7q
Yo3ii+kqRWuyd7EH2IboAcf+qOB7BSPLdne/N4I//v63Kbpwr3lyU+t+H0YseGtW
+eu9WN5B4A54+5vbXpQ9koz2xLg6WOJ0JvmVkmp3Zu9HATl+px4MxXI/lusvtHWv
XLLNK3MAd0fqqiHqcBU29hIwqbkdKC0bzn9qQL9BF2hU2pC6wVTga8o2sQUfvx/6
IimX1rShSDK+jCAUKCUmqw81g/p9gC5Vf09wY0rsHj3ddcwhkQNCMeyCI6t//JvS
c3yD7nMwTZrxz4dRW5y5hTFlauayAMHoXV0ELrkknvGR1vdDOqaQwKtm0hbqAHNq
ioNhulGkY5PX6PXQik3r5DnZjDh+Y2iZdOsZs/50P0LdqQifK2sP9rghgjATZ23W
0IR/uIqTH51mcFhwkGCskcpQcmADenWxjszWJJT7BH/CRKdpc9zF2dQ50HpnfSdh
IIhFX/hp7SLA0yhpKVl65ov1YuOBJfLwNSYHYeMU4BXafLIiub4iuwp59sOTEYJH
3487WwGkhxsZNNoGr9sbAIMv+U10pi5OGYAt5K36klmktl1iCi4oe4zAUc74Elno
rPZLjSvkhv3P61MJxi1PKE8so97Stejq1S9f4gtkNyzXJxpaMMIZZ1IJVGlwX4EP
B6EJCCZs0CUOHOkZIJfyETMzBx9QaWrtTfs7En7nfX5tAC4FWNQNqtdBlLAZPPhE
AQiy3NzQ8gUPrqdipYnGGBJwkv2lxLQqYVjZlpXeNZ/kKrg5cUPGC3EmpiBIE+jz
24sJCEF9gp2Wiiik/OUy6zkwndrYEsgam+fiEB4AqMFqZiNFboGrqdDCu4WWdmFi
WopaRR+EuYEn80GbMySK5j6Je+unJAM6gzTT888YC1AbWXun9QtbEOjT599TOy+b
dPS02bSoUhrikqiAJik+9JVcTjEpFiAXhHQEu4tvX9nsCxWt2dYdNySAT757Y5n5
n+r8Qtx5xIcX4BdKHx9WIbSscVcHVv+HHfz3e97iP35wEjuVFFvoOZ5Xky3uJ+/f
CMOnllB+jFCayiIjEM+0CE3QqAya6D60PKjF0EKmE0X4ON9ncllWrlVNIM6Da2vm
9Fh5AlGSUV4X8Mn0sJWk9KrUIksjP6jNAcrpx+TZiu6fMo9Dj0WDRPVmFebg0qHP
Aw+UbZAEN8voIffqYMnOM+bqQs07g9JTjq+8Abk6SLOlVEd7OrBA0BipWz8lDRzo
ZzqnVaicz2ZMclSjAzPb1zLDGK4BPJkN1y7AohzxHteq+X9/+IreTU4rmSbzgS2b
fSX1iUiLT0BRW/JDA55ociAc+Nf7tDan7Cc1evLay8t7vm19xPDO6fV7YhCMEoju
Q71SXn9WVRR9qzRhvYMoAwd/GHg53Jp7CEOv936IYsaTM5MJ7xhqkWtFHnHmEuK5
cu9poze3yp0h6CImhh5jy9CYjBaYWOrWVbSGXiZItrt8lj4MSuotM5igfxwcFzNN
UtTWO5NuAD3YG3ysHgzE6BVIMavwR2AjF7ndAlGMU3ZiJkKWd69x773FsspeX9eA
WodJ4LqkhbXO/erjyWSwztXfQTgHEgY8pFAWxg+T2Yd+ZvXHWrGTAphxxCjobDZJ
UOp3NVEm3uuLqeLDcj/ZFT40mZ5mRROLSCsbDQESw9lmXytJW7lbaB9fhn5vkgqR
xC8o3YUaIUH7n5an8rKYVB5pjJ4Fg4za1Ds01LNOC+sVbQtp0nkP2ddpzIQrgctM
NOKdLH5MytG4tpxGOFyC2olXNLIGJLthABTIFTcQUVmCHpSI6fIE5o/c92lw4BSX
hfPQJgff3UBx6B6nM84/jbyKCLCxghbEx6yubk3s9M3Xa+R3vnWmcSm65EzojSRM
ZXShZIYVw49UPeTZEEjMYwbUti3o3XkvLrtekAzyR3C/dAT7FPeki5y5eFbOBk3f
Y/TlejRq6zoIyZNzyxKbPnGUTsl/MFZt5TwBzsfVPP7UYQscz8d4g30uuk2Vh595
YOR7K8eq228eaQWagslBgj/4+6ovcySjhLDj8kpj+VumEvMBY2mbGYgZOQ3OzTMD
IlWSfF7iOIbo0VC4kds4+c+MPdnqufqRZhtxPqmr4pKG31XbQhVpcun7vx5SRySU
ayBuDJ23Xkbr1FQMNUcemgRg2FBy06HcJRcocaXnit4f0LEJrfP7JWCQ32S3BvnY
ItJubIvjU860pfWJJD2M7g3W5YrZPEsD9AI6Iyysp81fcglXWMDmw5BAY78ZVzi9
VBu3lRkHrXVoQt+7iDN4q8y90fRD0tpGOqSoKfAsUPY6LnXpRftHK0wsArtHq0vy
PYEAuD9oc0zHrMweeoHPThpaFPbduCKoc0qngSU64AHT2BZ005jMLScsToegD6Nv
UzffFQMkuKg4j1TXzJyQSCDke+l7SEG2E8pONZm9VYlzIYIEzlLgPwd6i14ZmL+I
BcxRozXyhQKRwR4qCR53iSRyS1fNy4uXHquzeiZzCWY5ViRb3ir1VytgrIBvB76u
/5J4wZt1/m4x5PATJFUYLyhzaPnpgLD2uh4eKJKfBY54KxBDagkx/7CXRC1Pco4X
wANoAHa/gjrUNLBz58AInRdACSWs64L0bA9MqGbvnA8GzO9K070gsnOAJ8HBqzoJ
JKDQ59R0ro73ZRd6sqk8N5F553QQIdJE6k2wRKmhxp142uuTwUe4Tzy6LZ2biIUw
7ClDvjwZXECzpmR4JADdMc1lbvJJ5afOb7Y5ko5IVje9npzDdasQUaHX7uvCybzM
Z+eRw64YB4tQQaUDSZF5vUBpSIxlhWnY5Vbj+78HUZiRdtR0Owx9VvVcPOAKOv08
bgKzBHn4WNIBp9tJ6flmoZgyrxfjnsREc0wOWkIXw5SOkPzIDm42gh68d2I7fH7P
7zQHJy+TBDJsTrYUgUeHz5Z1M1dMiehSyubM7ZXfqIfRV6Y2bmcpwio8GH2HoAVN
lfLMdv3WZiyqf6jxZaxWMzHbd7Zg2xZfeMbqW9dVCl/fC/DsSLCMF/V8Ifm2RjMy
v25kWBA2gdGNZwobgwXHprxhh9qhZwgKJOF+erCPaIi62bzfnPj8fG8O/meXDfLX
2Mv8Auoa+1mmtSJsUryxHlKidD8x85um4lK4MhlBTzCG3QGTHUz+WK+6/XSFFfUX
4oSJJllmWA3KgA9UxfqwzRs3e539MJ8w26BTOzD7LsDwlHnlBctQrAh/8X55etxB
O1vyd7xE69JzbKVmw6hjixVdJe1bmSp2NwZUB0bSUT/3V9RI9WmoKTQGBH+qqFFP
iTWOuy0jZGqzalrx8q9gNm1p8rbdS48jEjrwnMx1nuO2BuI010t9PXSRXX87O6yi
zG8ZpdYN5bncs/TSteAwFrJGX6Qka9F/fw3ObRyaZslv0GQbeJcPo5HHXrM+CoC2
V9WLUd84hDhr6JD0GEDRBJGRMRmZTW8NTxgKSBp4A90X2JNUmHi1vd16k/Bo73hV
bUcv0Dx4PawXwqYUNRPC9wfP/tAKnztxvPn6m24Ixg99MLVcDbLuuaIB9ZXaOiYP
JUvO4VRTlyD0rxFaVq+7PCrLG7USOjFU4Eu1BNekezfsFrt745gLo11kna9Dyfxy
6ZqCy90sUinIaGMvX0RC4+dVl7Uovr0YlrZpurt0C6ipraYkhiVtrVxbU0hfdS0o
iV/CetNVWyWDHnGH+4MZubgm5tpSxaxRzU4LLiD5KqeZUfIq5xpjhZnOoXFYZT3t
E/59xU3uY/NdI6AOgSxBj3FWzAk49e+sjKla3ExC4BsbhtmKnvLBOfr0K0b0uZco
u9z2mr1yk1BkMfCYpiwDBCnR8ZaK5k43IQTR9LUEcapEnAH7X29ARQggqkp4iHsz
B1bMZCoZZbA0og9TPbMtGSNU/znl1bI0Lec/lImWgeGSe7BQKCRUcHkCLWL9Iicp
gIh5/8kY/up3jqOAxTCl2MTFp1GbUDH0vl1NZFzp2Wcd9xqmWYzPSMr3y0Qw9I2k
25J+GdoEmbY+1GKblgl1R0WsZRar0UaKUTskidcaqMfoRnwvQfgdZWfNeTOsu4Up
V3oWybWOw7BXa7URYQj5GWkek5qbyded+PWrEK9Db1O8QFuWpd7HIK9yecB8ETHC
Qbtw0JEKXxMCDtNZuRDsigegx6k0s2MDG8ncEAj1s3G4vY4ErFbYYQ0ulE32CJWX
+m0skYIiBGOZ2P2WtHaoPhnCGyvxxdKHWdwue1BqSm//ElXct1WOxDe0HCu54hs1
h62SOIURgiS+sLa43KYyV75i9oCVfeWkRP6rwLMIXqwtfGSkemY8mYnk5gTWWL6z
rtazk8UJ2om23XrGUDzfIaFHvDGJQfiE6POH6Xjhrdv+r2EvYXmT+Xu0/t/Wr+zY
UeQcasTs+aeEJTQE25mmNjDYhIE6ANhg7RGj8e0lqBMlLmM61yHQWc3soA8tDkUR
n2lYbVuFa6HCVDDoI/Fz/Bh3MKFY9xJc8sWS/FTwYvBe+v+gXmMctlfe0U7r5flv
3wyRFilvPYnlVHNqXhlRs7U79vhe1K67pVHQ1VghuRxoPwOZKUqNCGf4OFuk29PG
uQg1lquAg+z+fc3SNCK8+5UbOJU4dtvtKyZXhzFjn6tBvh8D+NWwlPpfUcroHrfi
esJ0GRVHQpw/EdlJ28J83yezmIPJCgpnVIRKh1kd5UM8vsjBMjCDLCQjeRVF9cNA
+oRwjt2ixnyIHKtesPPK1BrdvlJR5TFkX3TQLG1lvkNgrnTVf6H6jhZzZqQiDJL/
cbKvGzq7J/RxGXTDRV98mXKaggxrZck3Wym2qRjp2aWwGnFPdJTPsJAyhOp7DAz5
nYfeBCEaesgUbej1jlhRVjRAr7LoSDuAiQWjeqNB6KACEA+aSFj2T/7+s57o7svL
+0qF8KmrjW244YA+aImS4JKGmS9iFKdB4tiw3vUIsy254T7UV6IV7WqvaOg/kw5n
rTGfVU82xD35bxSsobMKyzAnYnyaUZNOBtnjUtI+3DfIfaZaZP1hnL3sP0NQuwPz
CkkSLE3pEkNrL1UMMI6p4mQKAdBftjrOGlg0o0Fc352gwQI9MWImdUcA9wvVjFLO
HorTgsfsVjCSJ+MsRfZH56yeW9ewKymBjP3YQ2zrNf4dnO4UJ9xrqHvpnNtt41K+
OK/wmeurhg2P99o8YvCvt59Ux+eCfJvLst33Ujw4COBccLxOdjZM0adG+MyPmEU3
ONbTEjp+yyZKr+FOtUxbIvISvL59iLxCMhaWcFvO2Ak5in7PtqRNxhRMVOQOD2pa
jVz2h40UBQZg4k4cyM8UvzayBVwUwS3qgViQtrd7ccq4ZuaTcBl0tVucTps8RXK6
tH5c6fv8nksaiZTt33/ntJIhpmWS/OYGojp8pK1GO1r9babmBbkBQVR1UZeUnXrs
RvkDiqTuwrDs98g7ljaheeFAy4k6MA/DtfyTdJqubD8CYGS8AkLTP3WpFVcNIl2w
HMxsF2TgPafgqef6tdq01qEALTwx9yBkMcZQxxflzLZWU8oz2Pf+HCANzQdrMXCW
Jv1fFDdW0LeP6JzDsrCA9XzStvxQfO3i2XJatYBRupvLVHyylN9NciFlJilLlhx4
h0QlY843bNzH9lXMXUGxqAn6Ct3sW+GgwC/jfgvWBK3stmFddhOhO8ckPueFxMSW
aAkxRAlzpw48AuAtazYyLRXyXyjevVUhivrMviTEr1/puroFJ4nLhdch1RIOU1EM
bAJb5LISwH5opgAyjbW8+qPrGYOUVhr7FjC7G6h/rXDYrd0QczyUB20OoKMa+rae
K/d6avHdemlxGG8DpZe4Arrt/okdQXntrj9L6t8LFG7GtGzH0CdSdERWLsZZzKFa
HL+y40lPE2h4cM7TY/HOmm9wsyMJhlheLzhkz4fUWmLWwueVfWk7aCdmfkRL4egg
fMWmWfkDDGgyC5H5ah9S6HpdUreONgUpMZlGyCeAn/V3nwd02DSCEKroKAHtjIl4
wIvlwLZRY1+8zLi0zPe5iTrNumBU1lzmH7fdqKeFVVxxcWYINPontGLqc7y+2mBc
DZP/VOUlqMvwAZuIVkIFW/s6icZgsMdVUSe2a+aiXx4kLTOS64DHgKa5R7IwZwJj
PWK1nrDyBSu81eO0dhtTykOCWCpNJ6fYDt5x4kGWosSOsQbqgxQFUBRXhkgnMNAN
/TjpTtXUrvlZeJOEVwXpr8XXaJ1xeEjXt7rF8375NBRkWWoq5IjhaA+TP/8pa578
VLJmsiw16br6MsoUSEukbo4lFbCbfYpcXqxi9uoYvGAe6SEzBN4HeXFZ4Djis4t6
va9Qream3/qggRFOcT2LtZYOvRiz3PhFniqRlLJBsm0CyslLmUgy3J94zg+tNg+q
D3GFxsm4lxleivglkTpKnoLZlSbh6n3nrEfAbSG/XG4nCJGdeUz1LZOtSWW82/RX
6hXAnq5hzwmHlDEtExLgL4vdhORNsIWb6uk/643Cpn7n93hvh0Gq0VYzkluE0Xzk
+a2VY308gl8mJWtQqM1ynsXKjKZdjH8FBihAj72LVtRAMjAvluiTdzoyvhm3DMrC
NcIRMaK/kYjADQCZFAPewYe7KbTnYbUglVTdecIpTxgXHZG9xV0GPcSflJZDzs5J
w9sphsda65dgvDZ6hLhMVrrclLIQzJ6++gGgkmTaxPhg3Lf5cW+tFkxVlWqWKbzV
50E0g6WV0wmkgOt5qq9zSg7IeWkWqOAqYBUGUVzubr7Dn4dERasDFKHzIxksg/Q1
ZhR/s3h8Bp0nzSNrIOVJu+//6fnzcgmTMn32HDK3kn6RkR7b5DGSwjS1nOFMR0KS
+q2T+v84NQHTmYWn6YGe7NCiWXcrZmHzBQvn7Ki+TwAg0vHHDvmanaF6ndnwLGuo
7zvma+a0rOrPLMyToSqzvMmpR+FjzvPW2/DOyt7CGnrNHxjxGY4B5rbUBVGdOG97
Yw5T57iulzQ/iIdvSq04N4CVDgTyP1lBr8Up935+GYphK6F+t95wWzC7vE1AH37/
0g30bR/RGJyaLkjmLopGfE20OEwnDqFUyJbWfZl9KuF58OTQCI2NqZnhF+Y1khbO
p8ntyC0Mlp49yCH+83glkBj7co26Q9CPlbrZCRM47NhWkOVq8Jd3eNf6TSRf+RJz
J1P+4LKukZf6kBiWaf12lmXMcvMfkMoyHiqSzZebIm+NhzXcZVsvSqpw1HrCndV8
555/Q5IJ1YMgWzNkRiheMST0f4D0UOD2ndAJw7lmeZOLavPDwR6PfriyRVhyqNUh
lPNh1YyjKqoazMbowvStvmU26+8RdBvL/kr8qrq3pkdvAfecSHjQG1fdcTEsZtAg
lacbRv368En0SZAVuw62dWWfJYS4D88KY8MWQlmz8iopAJZ3AGCsOZfdJOsF1++w
rKZzVXdPueoShPEsnFbfTSsekenmDw6UreIXBQG9XcvCdA8JKJwh1ScqZ07ERf1P
LTN2PeD8xwHYioqpBh1m6ADI0+Sa22LxbXKpoE3XHTZO8Mo+osrU8KRKml55gg06
UE4enJs/xhOUkYL9tDKQcWJ6IJ4RmskMOK2LHkob8t7/CcAgQm9RLE2XJEtAnH+s
kHy0Aylytw1wpyO6GYV+TvUpF74P4qi3qXzjsvd3p5ydQKteUR0wIFtVmnMVA6JM
Y9ZEKQ7JquN0UyDCrulE2KnEgGlaoJy5fl52Nt5vO9oHOraLEtiefnnfu60JuuRA
7D7hwWTHeINU/6YvpeJjkI9YBVqmrpIBGBILQoFLCMnswwKgzFpprWIwOYhbP2H/
VRKPrIIHlcAGQt5ssE1r8+0I3J0rPfzPBIZ9iaV/gBDgprG7eoHAQq3qqpIpumQ6
Imne6UvNepwx5bo4bmLAHvMR0neLPMCYY8U4nIkhFzvfy2PVuqjCi9UIwJIcz92s
gWQlLHu5ThDw0+ZS4vqyGg0KS8A9OiuO6/fyFSTOSOfiWP6yaJkeZAj8eJ60FwCT
cxLoySNdlMhunNG3NadMMmUf6hOwo0++A0l4gV0iDQ7nsw38Pgq9XaNs5QVOJjos
BhGZkKFC1tMgeegJ1zkV3wgIHtnxLn4/P3zT+I8AckaFzdPMynYtGAwADDu9RN3K
GThTb3NEFv3SPUe65zMvylsg9Aa/RMCMuYvUSSYiOWbeI02tT1b8YpExX3XMRPgE
HF22MaHScY0YLVF6xyGZHqFytFt+TD7tPtJYXCPKT7dZ4se1d6V0SWdZEWgqclch
hQdo0Ac9u6Z2KvXZaG0J/slFVB0qiKY0BOpk8cbk/3hJQpz2hDH3MIaIZP/cEIlu
RXeu84aU3o8s/wgPS6ah1POHjWFvvXr4e4m7pgcpfiRk4JOGmpWZ5edhjbetlCiB
dD0J1TDHhgKbUcTiYfETRD2WrguvodwVZ06kxsheQ1quWtenEWzWQvoU8QCPFSqO
pN5QTN6ImDUXDK3q+jr/FKEAPHhSmoSKYFQTecsPVWiPLM0SUOnmx8+Qoa+LqdoU
Nc7lEbN2uVFJwigTeMDZlNC5h4hA3fXjg59vCA9MiFfdtEK3uIzbd1uQDkAincdr
I3WSh7XPeHekx3YrEE67jEdBgaLQLEWiqneORnEV4IyqDT9xlkm7SZ04LHa5Ydux
Jyg7KQPiLdgfM+mFGVYO0ZcxbpsNqHW14Zi3lzw4UH/fJGMwMZ5r5I22iNo9Ml+t
NILY9E8hg2QiNjuKQoCSy18oIfZqWWXBdPnUNO/3S2/hrdY0kF3ZCybllg0Vr88k
n7Ozf4uZgLC6D9ZmwGMHXbqFose6BizTY+fJPuNOqdJoTL847lMOThdUvURua//Y
32uFjZd7x4gHiVR0KPGSOdIV9xwnWKxBzrLCf48nsVtpgtDpEkVN6K0eEIKkg3oG
I78QG0bgrbsruVPdZ8iJzTK38J9VHhl7KlRx7JaLjuWEqx8mPCTIX421sN5oEr1s
J1j2RMQURHsdwUHTNr2VVDyTS7vqJBY9+xKb7OPEEDx5a8MMa26qE+AUwkn+i2Qs
krrPxAApRtkfnn1RESmC/4bd4zoDOYBfMdhwj6mQtkRnxnVln2j6RkGvLsomgR+g
2scuZIc0CPnPy3HwYrZSJzsrSK+4VUmtIkyHxmSR7cI02f+NwSwlr5YOCcpOEMm3
HEsZ6F4X6XsEEH+mhAmwd8m4zKXPpr9YJ/7919FQcFfLG+RM1QXUcs51+prKVkal
arV3QMYvh30mhKt5tgq43wSxcEf2FQPjvN1iqOvnWK7UgXqHmsLpysrBAMD8ouq2
ErM4phua4XMd6T4ro7OQu0yYKFpDpedVz+S2gJ/0UCSwxfp+fJmIGzmns0Qwu8dO
EQ01LnMEa3zfFvAC9TwBKjhGdhcWgwlQiSueKUaVqdRfrToQuVetCgGJa0B4erga
NoVINSYR2Oq4C63EUrcroLwvdbVb2ollKt7kJyEvj8Pg8bd7ROfQnQpEeixOpBoW
LXSU+F/udbtkbLgdrv1PWwoK+iisSGtODgz8X85gH0FtCO8XIx5cSUjqGN8QO7c8
Uh/9AnMDQ6uRpoXxYUtn140K9MqmRFeaqh5FG8CVuigyoXGwN4yqfy2Z/twboFgs
O2Fv1o69JNpJqXaK6z00PkZbISWQVUOE0tBjFLROYXC+2zMQgSS6BcL06DZIXafV
+mr0aOOLPUfDJvey/zvbnQxPHKUaN/I3oQp6BUDSEUBhBbVmnplGL0vFsirArbWu
eR/n+tyJDMiSgpk0kpOUsLZgJe7R2XOLX991Hyh1+3sE+ITwZSQ3dVdhgBHdh/44
lKbi2mV5AlkEbo5KJjA9aeYvgdFwje4PMdk7TrVVviEgnRd4fNr9yGLPqbH0etC2
rjFX1TfqblK0q61IpfBz6aD3D2ENzBs+1aKiWFWRd5mXheLXxHYBG08vtEmld3c7
ddyOECQUGSLJ0jO/Om4IHhAM/2Q6clwzF56MTH3sqcWJJqNVQOciAiijoK70YUK8
WDT51+Hk2xJSpIizy5HpABoVbx7J7n3ExVgedldGMX8tctbVO1lOW3F9mVa8N8/m
qmqFerbCvsgrjW70DlFAi/n7puKLNQ4jbqsX5I/vCeVAPMnBeFf0Lk+v8LZf8Pba
5IK+PtVt8NPMKWwEvELRzVzN6IMEbNzHYBGho2BM4iJHFW/mMbjvY4ZY4V5/2Yqf
be+maq8dFp7UHO5aH3cDebR+WTX9JdA3VmjWcRr3naaL5NXMUqCICLVLsy7mewZ6
SNKZmGi5BRFPoXjoFn023CQqOcjSYPTQGob56nI61/0JpSj68uTaCL0jmA+Hs4lX
7QirSlC+WfGevjeBy26DHV51dijHssfhbzaEiET58QsZA4GO1ugCzx1t3+llnTYq
IycWwlbFgXSbBLh1arQrXLBS/QJm5GWwXQA7NOhzkonP/SjdyLo3+KLnnsmrpWmW
/yX4N7hXcTyj8mqRIshniL8aJftiCMCkxApW7Mhlrs+m5md/MiNiWSMUlA8H4vN6
/Zyy4tbXuXfIJB63AKQKPuSQy9vO49Aclt0pbQkE/qXTUiK1rIGJvX36QIZtlfQ6
wy/QWeWsm6/4Hs2gJE2OUnyH2TvN+eQdxSXqvdIaDbu2Qz4bQ7vGJ5Rokc1s5yG0
Z5v+4oWhVglchvCy/8RVw6NVsOSunMvPmVpz8uOspJhHr0J6al3DZJUh5UW79Iii
7XhhH44WPWacs1DEBbsEiilEUMp4D/NmLY5kgB3+80sBge2cO+oqB4PEBeq1dtPo
cXMyWTivRMwIb6kIkeTcVLC9eI83T7SuGgMaBVuMb4p5fLbC4gf+uZBG5Ei1P0le
cBkPfdrx7QKsh2l80q3t2NiUxx05xlZQI9Q9wXO0pyBdiZU9QhRwbynGxc6rEGbt
QeZDnzcKNOyGHiI0a6d6W9wHgvsI0VhSzBzXEs6p6ZDoMqOImwM9Z2rx5l65SGAt
jJCGl46E+AFmW0gXq1506gFmCpOfP8jSGpc+yYesA8UD6D+wDRiXTuvjJjHp4hFd
judnhD2XOOjrLp3IdYLmqQcFZNXBdZENDGpcz9mKOMwMSuwr4Hq6VRyFIJK07DXj
Lj+XtZq8vGusr6Nh5tRosE+yTHlHagH1RSqTaiagu187uvbw+ciwTJ02lCy36qfA
/k+qkkbC5gqjgstYaZU2T+o8jw8craakdzLwJFZ1FEpfdV0tRi8z41vTBk1lvcg5
X/HYt2r+mg75VOwKOGSey5OHBVE3NV0s02mzRH2CfJR4MWSIWPIF+JhR0tPcohJC
LIRHeYrXNX4WEbmy+mHxAQM0us5r75coV/7FeFEONUu6EIvg7BqyjzGIYwVpAEgz
fmNImTcY0n3k93Ut9IG0KltMZB8qvEkBVjET8vGGR8GEKfDdX2ccBIdHorcn1+SG
v/6OyPNh8p6e49s57SsYxyUBUqW5ITScbrREwX2rrCnRoKrYcJfmYqE3lNHqgnE4
9cevt37kQkOK92kCgJOnLM66McqxUdys58sRLMkEy2baMnmwDms8Eoz4XA3A6B58
o9M1x95tVnUxECZolqaKqeyvHDjyvj4aAphbknBJWz573jcffDOJfhV9ZAHQ8759
9Z8StnwwKM4Ba8yDbeLlSZGrp00q5gjhs9s/LLTxUT/6fgdUPp7v0CtrzeHzliiD
cIec3SijW0g7wFeDV2B14FJvQ6h9kYsECVMWoMfwF9gqxjpI9zEU3p+s6TebDbiE
MxfD/HRUrA14tt3wtiDGHw2ldQJYwq1pfLZ+kICNqNeTsUnKY7jHbFaboky+LFdf
G5BnOtcoudRS16K04yMIg77L6UR8+xnusSegUgy90t/uqkC51GLf2nyrfXPjt1ey
Sg6m30sWIwn/Zc3J1WySuevL3VziXFhgYBYtgf8WhYF3raMQ2c6QRtFfJhGrPwdQ
cSt9NWJZomxAwhOq5iqFmHZmcxW0HZFqOXkC2YkhRyknjEP1zubfEzLXA6O0mbLr
3CGpXj7NtTJ3BPEW/sn5vJzffHe1eWZgwS7wBR9ZEoU2hXjeLULqb9HEGTwsX8q7
kIHuoU1K1j/Lxdtgj0LUqYWoAJTOAMzrDAQHAG3LTeTXJc0Ua/bJhm8M8kY4G/bU
rw0oeKGmd4o9tu+gB053sCrgz3MQTF5nmJ4VgNwsnvPHMH2IEZJXQ2CsPgKy0P+u
h10qaBqlOWNCGuknmnt5JGOJSDkBaFfXCNAOjIHe7kFBLfY4SXORtUkJXOLCuEo9
Rj1p+v1WZpxEPBW/wmq4nAf0PaCwZMtxV1oBcOF3qq8WyXkYTeggU4b7boP7a8h3
OgzL8pbb1ehivAWiTZ4gD+slvNSC8JUC2GqgiUt+bErxWcMmO+0h+Wec1paiIJZP
5yYbV9QUtRSqGAcZcHuae8aTfQhR7YeUFBhYs44+8h+QUKKtR88r9qYAucNNFpB0
EwxKSnEe5Hh16vRlpa+Ivpx0K+liYquiHfto68vcKgoJj3Nh1S/k58B5iC90MfPW
jgX9AsBqbrjYvpugSoFKw1Q0CvpD02BRdnDyEYdyWbPtf1m5IJxCXLY44qgz+xhN
MbM1oV+sC39mTDyY/OATwqbGmrwTDXpqepfaDr3twhFLMt165dKzWLKKFlb5BZXt
wlhGunmDPi9TREogLUUQRKjVccYHgYqb68/f3uUPOVi4aM/s5jS40rQ/u/HiV5Mp
F+E6SxDz/GTuH/i0+zZ9lsCyl2n6I3EeQutCR9kZItnD8M7+ex/v6AIoUzoGTn6h
WUe3skFPUX3HWe6yQS7zQZXsVMDXXjMzAv1okBPbZwpMxPRixxczSSr70SSsMlpE
3WHpNjBkHhD1swF65ghRX06g1xcv5osY66V595/gvpd3YUM3L+TE4Fsx+GEQosTT
YEwlX5DIyak/W1pZyrVHAkwESkqRH+bBva7I6NOMgHr2lT1F+kr0q6GG6ZZHhGaG
oqqr4P5oMPlzrUsLqXLaVgue7MaXqjIQYuOFJ6HYpFY5CYgfOZ0Y4YQAFTmgrs5/
BEe2Zj+uVal4vZUwUC//cemUexM0N5mxEtP/lxq0H+eCLmYhVDm0l+1QwaQkyxDF
WcMuZgQIz+tEM64/QF7lYYQLbdFwPw9PHg04YwIPUcv75GoT85HrzVcanSws9ZTJ
wz6Ct2103DF0EpvT7geTxXbOIX8pZSVgl2QdWjA02Hj7VUGTLU8Kf54Tu0epnrzZ
9zC5jO36G0wJpSG9XlcN/XXt1OtSMIW2Tlpvinu9/SHmbpHQRVVajpoLYj4rXdq5
0tflgphcAhy33eADg6VIhkChEYVmDi9WzF6kl9XL8A5AKgIX9zaNsJ0CnDJ0C50+
cnvRBGXiQA+44ThdG6OVLImydFBSutf5NcAdiDvdN9dzQaTE2DS+r1CCfC0Zh40T
2nJzCK53bD7yRs/DUviIMyrx9oTLFZMiuOwWL3xq3EZPXSDlBAPOM+e7s/KWzKqD
Gw5RdEx7pBWfQR7SeU364WQmN2NuMqtgZwSxdlUsSXrudVXB4mMoMyDBAVHEQemh
+1aXBwuT1ZMeIZUrZHDjxxMxXmQ5tZvfrIjI48v+MpFtd+AZE2kFOiEMjbMp0gAh
1eV5e4KQLSvAIryJ+WjzL3q8XxNaOfeefg5kXVj9rIXGTHvGLWm+HEg+nXr2bKbr
6ATQiJrWMTD9RswjBOwS3yQyjEUSuo0V7D24QZF7GXaUDLY5Xz27QJlXLAJzpwI2
rPAMGPSwxn5/Za8yK2RMRfZW11Xmp+kHYPl2jUIUJq24lMnMP498on77HN/cGBEv
suehufPMKlw3LsC+bUn6kVNFzdK6SsGL/CpWBcdBKrEljdIXFb8u9GAn5JjhYJRO
TJZrf0WYs1Y62XZWRwFsQ+Tk5dbecZq23mNv2CDynSuIBo/PGi/bmZrwu3nhKCaA
Y7VDyZSi3snP7BNa5F0JT86J9LudY6p22GZ9GVVUJF6yfnHTS0WY/aq6JUYcywao
BQiSytXUbJy1htAGn9FKJw2kB0BD5mCHMWAFfPPBn3W9nCYgfyjR6KkileSk3swL
iTRS6T2o28BYDbofWH/sIWOmxMfgM8MA1b/ay9tE3YZ6y8h1aVKcucDLgcw6DfJD
HsTlTBl16y1sx5XmNXze7nUw275uU5Q2SAVNbnXM8yq3eaW/DxtJHPyW4x9QHtHi
hQ4mTD++ckGHkg4NkkTSo/uAfHOV0onQ2DTqDBXa3ndU5cm6LlnK0YDxABrrxBO8
daDSk9hibspJqFC32WkzaVsUG/wa2flpLIHGZfj2WhArywmNkGKdKuU1GDw83/cE
F7A9AFK2qwUqLEh44jG74bIWJoqpz95mKeJWeGj2/+A5ERgXx2JdxdxFAs/0kYCs
Q25kle1vwOhqhgcWv1KuRuO2174cFLiYuK6Yjxt4xm6cgI6g0OMYoClivQJCHln3
nRfVXQ0JZb9LVoyAoTDjmrwfYaE9YOXcWwP/tACnDGmHykUJgyyoMBjdtsWB/zZb
O+U0QfY06psQaatBr0xBTzZC8r0vVytJ89ButiMKz5KmdcqAOgpqDwpItolj9iGx
pFJc35ieurxz2qU6KnsEwENU/PCTCgSM38DnmMWzSTTNmORoW5tl8LpgEWmQa+Wv
WMLdTOpdMbCi0/SEvIgWkaPaQkdMroOWeLL7lGjS8ahXbE5zVrsd4+w05dlZIIQF
jCelb7DkaLKWjf8Lw1VK+XLCrkpyEkk6u1vdYci0ImxYXqwQ8++5c2BpxlnIHZf2
zzRfSE4aPcMrYKuiU93K0cKGS5ea/+uIjRaNavtEWHQKPua1vXoHb4CqUBtfDGkC
lbOK18ja9CiUYjfyCwC1rscEKMMypSQ1qOhwM0YOB1jqUtRQo+iBKz/qpF4dKAfJ
tDf9O7qInHmAH8fWdEeXrQD9SEb4f9gsdKb/JtF7TyFbAvS3tlD9CixV4dzGMmGB
g6cGVNK62OR5uf1ETShnQLimTQF/JKo8wnil3isIkX0qoVznn7SkIviIg6a0Ocn9
UiEE12jGRVLqBpPVw2sJler9MTx+6ZoIfZam8RpYq97izqOXOEHQaYDRtzU7UfIP
YOjgasxba9lbJKNtkUH428au/rPGbjIvB753+nWo6yXa9bRMILp2XnTABAa0pRPF
ikJz3VDShWNOgg/53slE8kndPwue9I8FoemzbMnvxOlRrqQ6dXMzZuxP/Wg7p1yt
Jcldx1V0s1UIx3xmbBTzDlisnmBl0u+P5BKVO/6Nli5D5jSfNhqfyrFjAOT+OGdy
Eh8sSTegwIYiIcuUTv9QEphKYcTltvrzMCVTmX/+G/TMntp946K8Gk2Y0751ICnt
6UTWKTLk2jTM1hIG4VtT7osYogZDr57km+mgFd/xZxWIJtT2DYNSi2DC4Ycp5AoQ
7MYoQh0akriDyiByxrK4EveR7DX/lT93TJwnErwxIlLmv/M20Oso6NvDBKWprrud
uL3/fYdwbi6Q8/hfzH2Plrzdn0QHZAZATg9VuKOEO2Xh2kIs24je6fYbrNATiEc3

`pragma protect end_protected
