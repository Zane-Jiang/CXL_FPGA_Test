// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
dIzvxHYGN66vuOUKri7B7Ls5odt4YYmuhGRN5XdCPP/4aNd3E785pua/3IKGkatU0H+FUFcORqjM
YKQKVp7j0fsLTOM5ZCd9uBMA+jdV/S+hNliv5Yfdbbix1iB3+t9n1t+uJ5HNkJ2Hbsf55rdIMaDe
mWd7F24DAqbZ1HWVoiW4iomQQv2v1uvMSo/Fa5zIDnA6taZu5lA+aO5lVrPgohVYuJmOlK0SpBRZ
mseLJ5jbzCJDXMos3+J+y3MeN+XYXHNgSkKh5+JXa8xiUxtZEG2MQ8Q8hWN20QXdt//c5zp7BbeC
I6qYphVrGUkF2efGF/yPABkNCNRU++ZeW8Mc2A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8544)
LRk6cHYnyxw69dDZ+bsbfMrYdLW2OsNyUucIda++Dxr7TGLPKL0x836jdRQcy/CUfuxlx7yZ+vLe
OQwGgu2ecz85vvf73bx39fRaBtzvMJkklQd4kVcIMDbkiLcOECcgZiFvDyINxOf4FpUJUheg2LJ8
wjlM3HPoAtbmGn76Ie0CJ4HqLSfWQOP8xyJt9NuPz4RtOhtAE8SR3IIWOEDgyrEgHmRgLErThovY
azBxPSksb1zREwSV3SeUKSIDs6ccgGT3nyFPYBO76YV7EovtxIDSpYyODsC//NNGaAq8iCfoEOQo
9Js/O8BUf39uX7FU9E3Jis5Q59twINiGOPDGbR1HW47awfbFa1X7WHJuRpZS5oQ4Cm/zmwqTAG82
Ryp3AQVz/5oU/00OzYnSS8h6JlR3E2ncdiR72iMuHRIIHp/et2kUdHnxT28hgQaUdTEwLWVEIzfR
zwhcABntgczXOmb70Q4lGqIFhsITH54OPFDco+EWIWBeOEKecE9T24qJpSA57mfja3DM2W2BOKt3
EcvYmrQMma1MfALUDeizg6wMKKuibLHdP8dmjC5V17W+rbMjjLdA50g/jfcLAeIZ6fD3tGNDJOol
ekE2SBm2K9VAi4d3SvsZTqyqcHy7jtBYBnc9qPKV9I8vPUZxxvq92e4NDgI1Z6thf29ZKRTeZ12Z
Yb/Ibfr/FDb3xO1C0exelIArwa0U2Vwvvrmwh979vdJvycJX/2I8FTLQddqdM/nwaVHSw0QYsd4i
i8+cytzBO+5s6saA5DU8HsSBSjrpCvSjcEUMpS9ANkA6GKq3Sc3mH2tpv3sNzyvaO0jKUA1gUycD
BOZgYPCjtDlifIU7+oI9L+g//5SWGehY9sxNcQfw3E/djWUvJ//r5o9TXAlcN6ccFS2sAs7on7Sv
Vg60Tvs0OTJikuVPWWWcVlDUBzkCwQ0lx6jX3SjdnS5SODojlrR1OiPdFpJ1l3l2AD3qek9ICEz4
mltLPjpQUF71CzXrJE+ViddwWCVpw3/aM1BwwR5XzjLuufTptVE9HbPLjhvLtcz5fP/eqdZJZmUn
MLf5vOl2U9ZO8T6T+afB9ED/KTfhPkAJZy5oVGmRO4KgyZipWM1S/21MUDcy1tBfNCauUipyi67F
hGdACPUZDsqMbyS5xoR47qykFTRP1g1XAkOXV0SFPuXW95CE/lWS+uRHUt+/7Hm/eCSf55WVHtm7
5yQmpwcK2NLo9vH9IjEe+BZ+4R+tYGAbj7WD9R9dN+O2h3PY3lLdW/9OShPUXaWoSler7DZAhJcJ
v0Gpuh3RulK8ukpKMTqO6FhRadd3cB+5ljei9Cja/wPYPC+zuBEMs0a5V4iGFcTY+E1l5alSAwfa
20Os5EVtnRISvSbIpMDY+0TcBtQo8QlzATqOjj/k+JHDh94suK3eBFm+AHtR1y6McM5NXv822b1P
tedG6nsjttH5GhPCrdHmGY5NpHEZRpqW3YDvrz5GTZDf+N39khLMkmvpOQ2qQCCDL8Wy2KHihfNU
kJKPQRxShjULWoj/6aSHzFO7G6UksoT9sknNnR4Nqwmsg91P4oKnay55M3yMlW1B9ERIJpQFwDir
ab2zgHs1Hun5JEwcozqax6aLflEsaavbQhaLwNQQ5H+Q8XIYFPCmD0maX0viPfmDGMPih+leBYUq
VixkO0M0Ds+JZzxaFEKwT8slOkdd4SQ2o1e6SLdV9F5dexVx/pNN4UYlgRMDxLBWqxP0QVJSdeCV
W4s+mjzeVXIMBWUAQXtTCjMEStN8XYWGMF0VFjoELrbxL4fncwS8XNITzt0jzxawY0oWmko3sLzF
T0pKgLmiktAExOxyq4eqG5+b0E2jZDqGW96uH9YJcERlRkKqXdUP5uWdPJZZpzwtlJrG19qN5yHJ
FhJffBkFO6cyQz7nzKzTL3jYP0oM8Hxv/t94CmMdsRdUSzaYTLvoi+rGnDcrrpQYCZ7Q59peJ+zb
o7Cl5asuzsMMFzCNS9jAXHxaQNOSenF7Gvm2Xc3acpVweVCPPAFwvOuP/tGW+lbKmNjU+R678ZIw
O2OWpDx6qSxSz+RqRrEe777qaXOd9AQ7bcBT0m4DBUmfiVrxOxF889jcghoVw8XphKB+z+yWWk/F
MxQ5aSRFJax2Ouv7q8wuW1UlaJ+YCAXCC1KCXQTbjWrke6dyHKgv6Zjs2mrA4m0qj8u9ilcdQKgs
Z358x1AHiUvQil8QodyRh2f1lPBj6COyv1ixBurZK+T3QPDQeAGMAODtEHWq7+Z9fgDeJcCnhJwu
GrRaFeiSJu1wufC2tu3rO3SIcbtuQZU7QU5rjdmivQiTBcTSX0YDtSxpn31Pzkd3wdt5KTG/k2Kh
UxcPgVDNTRWPtz3mKzZV7B/hPKfDV0yE8hnKclVp9qZSn/aK8/VlL6x0ULsKTars7+tF18RnCJsB
cWBwe7wuOcnIYukdsS0ysnL1aEoeWtcwU3NqjcixF9fTIkKSAwzJtK7sFw7GnJ4GXEnCPDqzIVW4
yrXooZMp+Qp/pi+YRYydobxhGyyGImfAzcbI9MAc7JbvYya6X3UFkWYVKHJoXMQkSTTarXLiiP1T
pytpnEDSgDeBchFayqYdreDHEwsZ1gp0miVk62U91xZ7Z3RrSVsTOpoqkeeDOH/mqNZtYzKC015d
sHpVjKhuYcLTWtm0OIKePXsfKBI3dCLgOeGZzP93nK20MvNHqqcyN23CFqvbmxeWlrWGAI6Gdc93
dBpi7P/G9PqN49m8XppOrgzvZA+3AV4QDuf1vKkp4x0psTneHjGoTu3pvFch2ABp06XkWrRuk3x6
KFjpuC7RZZ0I9TJQ993juB+uXwW8bJ4NgFC+bMnZIkQN5WvLMMmu1jXsaNZcMSZu3A3XHPYuuwpM
0aL58Gu/LQMEYuv6+MQf5b9vPlJp2xUKYYMAEIKw81j+C6ZzuySck6RYtJJKxZBD6ENLAfVWh0n7
LsrjrHXSJhw6sqw2f0z0h/KXwfaD+FUU7llaRmKy+UsPhx1tunkOoWy1Jhwo+nVnNzHf/VMH9hZO
N8YNOyXqaPnM8aypxJpjHUatZwjNHapjtb1l3Es04G+u3NS2RjDmOH88JhTzj+D7kVvZ/7i31J0/
SrMkANKPTQQdP4pvElRe0X2pyxjjWuid1qZ9n8foU6kjPf6plJ1AcRO7HAnrokuZLZTXmmwgrCHa
wBCC8fsgwHrr1YOZN2ncP5FGzWfb+v2161D9dNeGd3vER33XtKeU4tQXLk5OcmoLJ1jF7AgjRrPI
maNIzDcDl2+jXU+9ASLRUcJdpnDS3dFJJTgkRo2d+GQ7gvPXrjDmq2ZlYCWx0g/qEKXqoc6caiVB
QLR5dNLJI/NNsEQJWoSEWm0nTbXtz1JsOedXCE9+Au43KsrDyvoXKY49B+aG9ELjn0Gtm5R4xHlV
jAsv4Zi9Yhvr5tw8Iqb3URSViaMwIfY1LZDFhRlA1LcCmQW1uwMklYjGI8HmMQudxky6GkPBKWS9
kIMSuuL7dCDpES90OKRItmDN0z7P0bCs3PV/QY2ZDKfpaLmfXBQ5AZKkGhwoszCLV3itdZ66MD1u
mM4AfJbzCWZ2Kt92sZ/es4c6pu2qG5ISlt4CFWyFd7hQBFNr7o7o3L46yIJVc8YulwfYG+rIKGgB
1p5+QzI1kWPxAgIZ4j2qha8FkOncjU2k4QmoU3JR5onfsK37NPJ8HTT/NFcsHnWpGFC85WfzVx7d
A68xnWoEae5UfxwNKCJTrbyNNZHxN2gTOYubsvgymSuntplMHLp4v1BqKRI87u7NZeGSqE6U+BuM
QwVDAE2xFInKijs2OIH84py7i0yhse2m+TcvNd29425adYD17395QrgPAdbB/hhzOMBeGbWFkqRl
Ao0YHd3Pig8qRHhoMSAtZPKhVqcW00/MxZOxo2dcq4dwCeJCihYvVqTPgZP0r7ryFXnhbB6GY62A
IPyxMmuBt5xPoCLsr/3n/1N8OSyqKpNge3PAEJctxlhAowJcgH98BZfTd79FGqAtfxEJxh5hL+K7
MwNx8oBm46X9XeyOKzyfMjT1c02RvpsYujVzFWVAa3gPAd0K8rXgRM9a+4V8vBuz6zIR7BlQWPXz
50QnvuumTg8n+cqPoJI88ehUoOFK4bLdS6crNnqmUMV9nbg+y17FHI0utp7XFRFlMvI2rObJdi1q
Dg3/Z22oub6bvkUvBPde+x+NdJWAJpWFVAdrlXp2BXpJhkeqdJ0nB4OrsmX7FcXKUgTbHUWqOJ6j
yHm4T7oxC7TvCU5JFEgLjKB794uTy3vWKyx/5R5B3ruxRL992h9wW3EsyBD0oY013iaSIPbY7EZ6
YWaTENFM191Va0MPspmEkwZGXN+xdcXsEOesxTcQHj9EOyvLfagrTNb1zMQyLX7HGzDnKR4RYrKu
7HAWcYt0RnsVAnPloTIRFiJf0mP93stuy280CZ5tpYX3C2Bm78e3/wu+23PoiEG8UeKBI9FMrf91
m1UFJpcIBmhSiqdz6A78Xs972zbZWuZDVDgdwzdcl4PoJMgFh3SxJmhdKaCw4n9ffjWcAl53Mu6W
W2Ka07Xzxc8OHQYfjpFJu5rroRZWNWGz7+qslQXgRpVPc8nAMG+JvNJ1L0XSrgWyaxgO7bUqjWfJ
7cC/rzmWrNZ/MT4Z+uMsUpogbBjtVlxm6JCRgiSQ/fnp0pUni2K9X7MZvZxBADoM16CzniHeeGSX
AbMKcEzts0KXclJrVC0Ww0GPaYQ9UFqVlX3/PRaAOLtYytkor5IGlA5PoemJ3LXtQ6eNmonChnkV
aWa7MbTPNjDYqhj2w4b0g54F3BiuV6+mjyj/ifw+jBHB5V626YGGCv0mYfbEU4WFxYr3PZSbQrNd
pLxVDgA1LKlEJKO6+MPmjM8KIEbEVJT7IGAdd4AxaOw5XB/zR38OaDPXl4rCTzAtR9jqhCgGHlEw
Vm2LYqYU0o3vw2xWTdkXIzb84t80ySUJzxEoNbKmrKbj3WKedE09fkygPuzf1OctHAMZ5W4d/0ym
S+eUZCe93llmEEdkaX7sXdtOrctplX3vgEtdPjc5QiFcph0TPnK6C/S80LByQknaqzKNEWYTBRfu
fhXap4ko1fpBdP8OV1Zj3OuErAHxNeRCeAy87sTeVpGLfwpsoSV83MZX8Tj9r0Yzr9bE6gLXlte1
g3ALtE1Dh+fOB3yCGAGh8wBtqFkAdCOAJuh/b5mTPGpsx2dkuNMfr56EBl/bCvHJAIWRC5uSz8Lf
2nldPs1qMpUcR1ege3nCJr2D2CUayFMz9bzAlEzZipIyZQjABacJH8wvjZHS8UO+kG+snY86e6bB
COBL8FYVUYm8UL+xLNHl5+BOwDqfHjUH17Ms0RBUM74fpUJwY93S2zwL9MuuiYZroC7G3I/DssGv
ufAHJcVvITTmmdxeAbv8nLdyt1gmoEyZJo1Fbb3ybjT872Uk4kMKCyH4Op+N6wmbUN0drsHkWRIg
O+IkCm8T/t/JbFSVbeYSq3mhgoMBL4/iCvWOdfnaal/GGNwRyHfrWynDulgVXHMFcGS1Nxp2dhJM
LWz4z/HO0uwZYltoKC3HGuuscdlPznfkEsMUWv/1HiL3u+umpRl2LUxElUkiy0znp1w2RYqLBZ2R
Zmf0QRpB01DsDDAZZgsdRiuNjCrdcGeFPfabuvSVJAxkTOY2gOjAScbK3zJieh8Ij+8OmeeXbWeZ
CE/tCMcUHptq/dwqvdBi7mxHYLCkl8iI2++cx0z6lw6aOHi0YAt22i2VHBGCT8Hb+s4++SYJ+5DS
D4cYyTDAcazeI4WgZCjEQOwy3X3CEf2I48s1C0HqdpNoZhTV+9Hfi2sI6IpSnmIMxmPT1MwHgreU
VGnFlUt8/Uc5SLSzKyhRsqlND0Le46jWUzh5RyfSH0I8dabR20nymgCY1SsMLJIx8hh67Y9ZaPzh
EVW94Xnlm0fuU9m14fuOZ0SLUruQiaqLNa13NWT8CwbWX9OCapDx2KdhVn5CA/dRJWv3x4TKcMkX
gKqM7+f90m1H0TrILAVKjBEvgybDxAqTtD7umsD/een1uEkAM8zxV/sQ5elMesdv9BhbgEh8x/K7
FFoXyFjUNSuji5IUaTONKn/I1rTRH4zIdkgkdZEjEPSDIFlZ1OUwj3dANRuzXdBW3OfmhEry8wpy
Own2KvRpkL68pWOfmz7xjGo856IuZ+zOpKSDo/gCyNrWd1bz2ZyvEvTThSquezHlKbPpwd9Feoh3
cMDCLMecmDw8Di8FGX18+UOU7WBiwTw833uYFijEEThxPcjUbLr/Vwt3S7SYdnYyoayV6rSXtrUV
COLLS4d4lu2uoDOXAzfsH0DYKHKcJycjE+DfqX68tJTNFPfGi0CIoefUxp+5B6g/mTqXplJ89REE
cVKT+Le1qXh3X5COZTENVC8CAcP8mGh1W4d0YXdsYcxWLxcD5rSYkDlWKB314n1wDiGdMor3KrEX
7PqV6r2Pgwiw4RpbP8pNwJxRUDy41gcvcCnqT8917Ugv4opDKqdysfIGZe5Vw9y7gzKj3MN0BFjR
FUIISNuWJS206JUNJaZmbkx2hGSowKp3QVuamdQBZyiWZxPURKOsnhu5O8ZUzCEdSqTL5OBNohdX
1f+m/emmp5Twuf0v4OyAQpHQHsyV+5of1jRFDLJjovwTdJsXmCHHjY+lyPLpO8Bu5Z3mHsSmjImb
VYqXF+0iffTDFNWJYCrAWIAGcxgGlg2HJ+S+hxH6qnFxT/MtuaGylT4j9cF9VKEzK4hBWi8IDxfX
0N/sGRanWEh5fReNaWPvdxPi3SNDo8fw8p4QYu6OwXdY+7bllifA3Q4vDCbw8HPM8O3VLC96UAAG
XOupM5Spts1t/zsBiMZM0JBJfjQzDQK5g19H2P0qd643M2s4WDw4B1pYyNY0D5KkuNXE63+RK6JV
l5NC4wUOVHXZBMEw+6TW3Nx60aq5aqWllJqDI+V++2MTtJNu3Q8y7ndgEnlfOCRGUte74LRHhanQ
Ap998dCs2CpXk6Oj3tgMpE/ZK9dWr4ISk1gULQdUqlsxnTU2/8QLZxqTJaIn3D0Cy/Gvy7cJ7dbn
ui1mOmvrYCq+iBbmhqkNKAh2hGMmj1vSpKPWIHX0fBYNEW/8m+XCScVfD3gzYwuJP0R+xHWsNqLL
OguWkmaU8Pkn9KnFUknAZe4DjJOPtNP6wnRZUBQJ9A6KMqXqLv8obSdhnVF+7/73MY6dPPom7M1U
BAasftUwXXqSu2rkGLYVFl5e8PBbVelcGY4iVEOgjAvmba/qnvtW3bRztF+n18BgH6F14DKhp4H8
dtSQs5bl4URP3tIQoeg5BLtLx9khX8b7mk2cRR0F/kIaR/pGP3MdaqMkwMUuvQSEW0dcadYC6Pk3
ozUnh16MB8oQUi5prL2QBpHENmUvFK4ImbyW99mOko1anHGCjPc8vus39ixmli8tAYNIp8Zt3btA
tE/cG+jMh3g/RxecToZ1ODrGrwgCxxDwKyA1aTPTqDz2lLZBe/yddrODpqnLreqj8FHP/1G/vAbf
asWPoCBS54y3etAyOuOxGnbYmvjxYtkgT4AleNI9Mvc4PCdoukilZ/Cqb4msGHKB4otZa4be5BkQ
amqb0Yn3ZGeyl6+PdnQL++nLvugiDnBaPXLK5WATAl0cjv5dIPZmBqacpwqRHhGFQKbNgeHjb1KF
CCb6WruHAV1aOBx3CZYAYcVW9ogAtP/UFCEM20nNs3dkHI+GC9QnUZ2OQLBAg228ab83g4x4MHsV
8o8aQB8+UR8bbVATj5IHWoR+uKKqMhhGvWo8gYZiToA242a5rWXr+szU27Q+eXSCUxwpAfoR+mlg
n64C9r7+vfcWO9T1Th3ZNvR8OPOOH3q4dCDFuoQCXoSPSQLUB2065uIssDpWqH6+sSV8Xz7YSxhG
JKQJdEFTN3yKodb6BLiemXl3rltYGsE7iqvhdx/sAHlmUhYfEUiB8tJl1mp7Zj9iGnmrchMYH38n
3WsERoMl0vLFGtICeWD5H5xp1wUW8bC4LmKqOgrvIECmRcDcYUuXtUAoyWMU558y2l4XraBBRBT9
GznkWgLLJ0Ok1adhCdYBz/PS/ZmWRZaqup/bj7p6eM0TMo66v6ZcdRSLdurq8Dn1462uTZ56COf6
39W8elXyfgR18pW07Px8uWBJNVpTQDFMmnRTVy1F/B9pEf0l9VKKCcDJvTN5WBXTIF3JZ8+ELNin
DTY+R94p5yfLjIR7AcQWg3d7trblDI0FqNOTliHKc7FM2QHwe11Vjcxrl1USc40C0s/zejuFXw6W
KbioEWQnwfAu8ORDNQCIjWuxyrHg3QHcSWPwe8HOMGUKepedxd5tU6UbPmKbN4wcPBeUDovdmSNu
ZHuJNe3EnsPWoWYSstFAb2LTn9xv8+D7VekkuEIlwhXZgmAO1E240OZZJG+Ot4Nj7bMrgmEXsqb6
iOah/mq0/7ioc5XSWNsEWlG2LYdbnJJ/A0/R39sD7O+gT37SD7w1R6A1M7FDHjRmv2BQlr+NaOLc
DZLLcFrBvEbzlcqTOoLldMpOQa03gTjtdFnvAAaRoMMt2wM53/5/2ElnMRS9VQhtN+DTYKWBlhqZ
Y0Vtn8dF6XIMbkU+7Cy+yRP0Jccm8vebzkoNcZst9rTIn6E3HX996sTv56Lcv7AV/GzvnjsZEDac
H5Z39a2gPE+FbgRMMGVdq+scLGvVgVNmt2pc883GSBik3DfDU2S4lCkFcUIlP/tLCawNNgm64ane
wK0+IgnXV9wrHg86cW4gVYFFqGi1ePb0oOT4yHvnlw7UhYBY8KbgKbndkWYpNrPBD/NvtvJlg44e
s9qWojnHaO9Vx40Qd2NxpiUBYvkQmqyyg+nSBc2KMVXGsUP+tHHKvQg58zYteGWlb3hOylBtmtuy
R/lsnf8dvamkb81k712XJBUi6Q63h5Y0dMehmVBBidpl1noioZPEbsPiJqPRY9h61AHn6e8ENPj/
8QROdXJD5E8s7Hro/unz+Mr4GCDzpXG13gtrgrxwokEP7UHksgeIDGFEk8oYFLufZKaIh+tvikmt
Cz8uHyb74HLOww3Ti/lxN/1Ba2o9/o7BYScoxlIgN/KfABooTUFdi6qNO9atkTdqMJFfOZXvavwt
IN6+uIPAL9hpMKc+2WqRaUcviFFDu51WCdIbXJyGZ9nqQ15qiTNKfxPkWrRMOvdAuvd3a79ceuG1
khUI4KzO316U+OnVXJWxOw98Q7g8C2/jMq6pQFqeA5aSGNRmPPQ0h+Oy7w3BJEYjHyLmDehO0ADc
nPWA3V+ahqlSeLLgxkEF22waY2h2sdzMwFf+DX4nypUv4R8LMjCP8o4rREFSTS7GkY9Rjmnbw8Zw
IIF40kVs+MNPTfG7VW/aJIh9I8QWhshvOIBcimVekkrihZfYSviMK7AY8kWyDqCdwRZm9dXiLVwp
HsRMcoFXBsnyMJjIcE/AvVHOTCMJciuivrLm+zUzld8mgw69OtA4LJE62kYMvAYbZgHv5qQUpgpN
Vfx/W1tAj5lHE9xvZZrenuPdICT5CeS3T5bfCCfoHYqwxxgUUBaOo1lnWUcdTYhy+b0TnyPYWRfk
DfB1VcCtPsIi78D/cL03SKZg4mHXP/DfZdQySgRc3p1FjVTl5B8sVe5dg515JIJTw+p11XQic9QA
sOIyzdDO97JXFhFsvG7bQLZeZEssEsOOa/IjLd9KdcUZYHQejIIdR93ZB14PCLZg3B7yPuYIODOe
HpxUSF10Rxyo5+rVxZnVbwkL8ITvmAfX2nXHvKUXGWDX8YrtMGqOaR1v63bpbFhcTilkfrPQwN69
ZJM/eTuyHPNjvkKH5RqmxgOYcRbj1UPt27vAzPBgciDrYgSNNzlMQ//gsyXc6PyHE+/QJdVNXivE
geCUcb7J2rdLFF56PhIFFbK3ud2YkbY/CuHA8nmy4GE9n6/SSSisGtiKS6szE6fqaCAeqkgnWD30
noYHlkRBjZSzM4UFpg+2oHsGTkcbwh1ELvWZqORdH6BCfrSMW4O09v/AZnNSYA3c1HCfEvu6eLbQ
WJsb664ckahAWtITz9mr6NoYm9f3T7nGohVhoAuQBw8VwO64U923GOKOLpIUCaYqWGkOQNwVeWZA
GU5fa8yGHCu3iJeYp6enofFy4O+8Xk3E25XSj88C8ra6cnyIdAei7nsWaslANsENz/LWK1SyzYor
uFwBBDdvbQjvBJUanpWRQhy3kAP16zASU4rp67ZI1xYnCfED+k3/cPPqK7u6oN1/Uuy+q+q7uKkP
gJtcPaXt/Juzb5ysoCmwgjrIsk2/Mpkjbaz23kyWrM1zMMIezy60fJDjrTeiw8O9sKHxgg/JR1JH
8yaDQAbcwVrvPEhAHt+pjZkJFN4HYK2l/oZ58AyA+HU4cj5zetHg9Qv8dzCQfZjyiw7pVRffc5Iv
kjGA3JHcE4RuvbYM9OGsiM7Zm5BD4nzJcMy9cZ/nGXWbSftJj/vlyWFqWn9Lc5vGl7QAdTSxrt8F
Dm3BGoBsz32TcAOjf8WsJKNLShKx0NKjBPoPzy3YNsBgsZbhU5PwGhseAfovWXtfvswnd7f4nztm
pOeynKtsZS7rtXRobyKN8W6tcxJXSZ+U1qtUWo/qAHn52zBKyI66K3L0UJ+fXoK4kOSrOChVbLIu
gCy8hcpQFce6NJf8wY8EwEK/D55nrNQi2Eh8qSQ+foDqm1Rtqr0c8goH8z/mO9Y/F3wg8Yg6ro6n
EbqB0fDfh8zmyeikfxgXtlBUsg9vH6gJXtPRulZq/dzUn12erXcTtE7Rk++BD/vzfc5YxhVAMZkK
Cz8cMLFBoHnOUi5V55190Bzch1HwvMrE2zOHi7vr5+gfzV3S8ObTSyYNIwX13+gAO0lMK/Ab2Mo2
Izn23y065Kr+BZixekZcSsAnIvYvn/J9Yk1HqbCT7jV7DLAaUlbW1o5sKXzgDZkUsDyAOg2OCCyI
8Gdr36CkvZ42sXY6LCkdChUsYLWG1fzYkA5+w8G2NykCNkAhPsx58woqYVlo6J3KJyCa5j4l/847
WtmKCZS/7kxRiEOqcE5mDNQT1TM8zsZar5HRtuuIhqqHOd5ndAbVg3exzvMsVnoH3dZyzwGRI9B9
7XPoyVUv22W3+YkzTWF+Z6/entUjRgz/EscP7LBzxN5vC6GAQozK0OEw469IBWK5QyOZqZqubRWD
B6155ARrcdJMBPxtwjbc7cR/ICofovI9D0yAs9ab2ExfbcovOcvr3yBtRjCMjoKdOD3o6rKbm3rO
AaN0gp0rvPG9uBEs334z7Ntbt6jyMjyLvNG+/Twz35cJBwKnBt0EDu9UDpHzYuXNrqeOY+CxpuoD
AC0EmgvZo3PUafMzpsfgyg91o2+HIOtB49GvvgelFVbzE3yIIydIqr8s//JWe/D89Kt5
`pragma protect end_protected
