// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RuFUSH24Gtcdsa++rRx8izpEUvxfVml+UqDMEXJ/R0jvFSDaYVY5dcsbyy6o
yNxisxH6hTnY3lSJED7fOKjQ4NJ9yOcynqK2N+uRO29kOoMfJWCA2viWkeFe
Bam/7ck+DhKdLvnNJh0/9XrkAcC7YT4P93OlujfJkOGmZ7CzQrOnBF+tTPNQ
jE65yAyP08g9s4lfnHNQ1PqqQ5e1QXGxMrUjIlixbPtlHA7Wh21rw4B6Bl4m
bYheQOkNuiXtoOvm1j82SykkQInRGRdi/ftRAR6Bq4R9rOSavqcoafkn7cGh
Hu0kIiNEoIB60XOh2aIJrhlKvQ3tej+O6wPF/FYZTA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N9E3n8Wuc4NoRCMTyeJRi86Pp+jb7sNYUKB/qAo9Hp/l21AXlmBULvTCZW1V
9Ir+JMknA0xBIT9zSy62Z8P/JxwCZ0VJidUR7DNYASP0eou7KgDJ9FTQxf12
E0qhOorE28wdqxBxa3Tmr/7Cd12Tb1efVPYR5XqCUsn7b+eCKEuyEYogx8p+
L+Mdg8hzv1BtE0ToYweBE9FiE5bvE2OYzVp4wx0M4bNl/KV82UFdbknz/wIj
0ul6PtaYHrFt2kozPFQVpz3H11N6qAf8EJoQKD4pZW/5+p/LNt7IEn4H4BWA
E7PDgBH/JIqTAY0A41qqNDJMvkqrCU6roIgINBF89g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HG+2jKPlABZ49Ech6YF2MWDjmL/oF330NDEq+EFkxrhhSnRJqzVvGUMtBK64
oirMxpS+r1dbAuuBnN2zm8oHTkYs2EPTGYU08iWNGyfKwStmyg5Xidk7thnL
yM09ZWDdQMmL+XqDK8Q6Dk9zpbOp+xdtMbr4jTPwKq8Xwl4OEde6JLPTJcTi
1kp+CFoZs2Q219y+IKdLQ/Orfu6MXlYyXs0tkTpp1y5eEPAFA59kBtbT1Z6N
PDI2kO6QsBAe+EriDSYq4HS9Njln8fPcLV4PQK3hgv/gowKpwJzYx3P7WT13
qPkYJSHxkYwqdwicQyly0BLEOXrtKUlsTPr/DIOK5g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JSMMeuixblsBkRgvG2FEIB3G0aO22boVxKF6+LTvUKF/vm5A/1Mhuipx7/9/
/NB0Ei2KrPnYKui9rpNC9f9b9V/hQHxRH1D1IJKdpQYO8zasLaNHqdiH6lqP
A98M6lP9hamkSRuGG07F/4Ql/ESIVutUdfFc27ZJ9zQQC7bSrLU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IWs6eMd/lEA1Vm569xeROLO2YiINW5IxQhQ6AD8iuPVL1FjrWSuQtHWiXqQV
Uqb1vxEjvmy1HYKiAXRQPopNlqLhmtc8qN0DvOZV0aGPSKM/bnTfAq96nkLr
VE7B/67MT10KGgx6Ih9sz3RMsF35NymWXe6D4hzahoaVREQD5Efb/XmyPBQS
SCY9uw94qzs2n/VLshJCw9cZmkFzQF0WH0WORraJgDBP4VyuKFhKc2LrNA+H
PYG5J8A2cwCuGiLItqSEEMkqjeXRziWdOMSZsdcx4/ihs5D5ubGX45Z7cgpf
6CpWMnj/9Fvz+5KMu6L4s5xP9ydYKV8F7WTP8MjM6jF8hhi+cnmgDLu869Y1
IzS+6hY+1CNC+7Ior5MMRJTEAo0u+biNsKTDbzelrAv188orkJ+fwm6EAVhb
M1InE/vGqL9YG//IDLhr7iJwRgH7lvtRCWFHTBNftddBZ8a7hmgjyxcEpzVM
wNDVeJDgFBwLpQYltIIHEg3hSi0W2MmC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sY0eW1mIU6kFPlM0yG9pt0Z8qdl8N9Jy0Kjw6J/iDTc0dMmEccDm1ktd9C28
2CSOZ3q8XU+JvPL2DSisxTzqfZXSO71EfUrktRJslahQwvjIxV06AgQkz0SP
M2KTZXf2ZlZGeGwLHWnHR2Y2ozY3xVL09nd0z9bvTFtbMLO5hjY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LS6nkoWXu1MbdkVEiTW7nEwSyqCWB2TEU5YsvOCiZaZwxqaHDZ+PFnlFZEIg
cZQJ02IirynRFh3BiNSl4A+SJexaQR4bmkSF91bom1UaUBJXL+rXiLcuGFrN
GrP4KTQcsAHl11TaavsdUTLDIxJG8U3ZI11MKo6mpBHHbTls3nI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23504)
`pragma protect data_block
EcOyINng3GyGvyXxoUEc4NYHIv9S+Ns58E5M4miWE+8TUTSq4LQT+WY4njpw
0s9QlHxLwKx5lqj8InpOtqae/WYaV01X0MMdZWtNUHP7RXNwk4oYYNj3nlf3
TWfghZNiLR0pnvCKCGsT+3h0007g3IpuumCocloA3imr3HXhqIhm/OHRLsph
cak2vs8ztUeFwvxqvH6yXRgqAdUrAJLJS7FTR0MrUyMTuP/B5itgeG9jo3/b
qamkjAcc4gfifOsR/MdZ4+IRyJThzN/kmtKWphrRoTWjtT45wKZgKcnkwp3d
G8ieEqcPt3eWPKQjWx+m1UfcHysBnYn/OSpCBPrTXermt0nvAcvrk7wx36wj
LYs3NTP6JqSChxdvyW4b+dKUGKvNpNcIar40xPnd+Y/IaOFDQusGj1DHTZld
qn/fIsEb2VDyoDnbLXuMcz0Ehxde/PzJryAAe+dRjXEIUPIklYj+2Cwui60/
i0+jxviMqO9NMz/dByz//SHd2hHCB7qQxpEcEiZigmbsGEgfivLMYrvqDGN4
//zgj/e7wogvKJdrbQ+uqIuFeahPeofizuZV8LKlr0PotFgm5fOUjonKq1TS
sJoEldJoMQPQAWmjQzdilgOM7PRWbuM0p5Bw5WPMAEHyOPlvkEMGnVe+r/ep
tSQoMJ6LLY2JtByQZegKIPLwpwpN1WaLiWxWCXfkfC+H3YCGhsnMlNdoElv9
Q5esfpKV9UWIk42g7hiHFr1OQw3K6wU/MbKvnOrdix3vzWH9r8PMIo2SYbSl
XwYWnw7Ow5cZ8sZbPKF5gE/7VMJ7jGZC4PlPyVd7f/k+B7sh4WNWf+IyeF3z
qCqljS9cBGAVfZjhwKaVnkpsdcKTSu3k46k7uPzaPcObc91nP3rj2ea/2Zcd
VsRZXlgVIVzLajgyIWyU6fufjAZZtAD42WmZGozLO4Ng0ZJwavNHUjRswJjB
C0bBlusz1A+GN3tWFU5fi3PW7r8LDpbINWU4AAuif8b3zUl0n/o+XCUwAidq
KqYSo7gSoKwROMBPUpsDbgtIPTFCxIWoRJpU6JKsglAlm3uE+1UtatLJDiM9
YifND9Rptc8thVpaIqdpl+kVDIQWTqOLioBN5NCcNM6QT+N//UAER0gKgFLE
59LskrBGAvEHh/EvhVMemkBzqR7KE5Cz6pSaXZ2fyPpaZfIsT6wfLv5GDQsY
yZ5w0MZKkoD2HFMJFHAjsBBpY9kI2KDR0gpsY2uR+JMEwW6aZoyTqPGYswpc
O75Vvb8hPlvKXnGhcOgOlQSzCR+5zKw6yfpKAULFdTi/ccTBRsVqo7RGFLOe
P47jIqyQDT+Nhoy9GEdhuXPb2Mpqjr07JnO8oEKSCde3MPn1lEdlnKGN8Dsg
KqGGk0zEK5kPSO1LVOi0y+HCl0V73uGGE+pmoyC9EgIHF/7G6rjiUkQ3xPvt
bDlFRFpSsI3UdxwMGDqk56m9DCewqyx50Awy7t6AgE7sjkWm+daaqtaNC/GY
Dh9qhqV0vCNqe41vWBTkE42Ig3X/nJxLZRPlLIjaMLdEwttYM4XWZOMaFsfq
TfpAkNm0V+MH8Ze6sv/fX2SHTrfM2uu2i14v2ztLpHLku25JTKYH/dM1WFo9
PIDpS+MAjTH0K48zG1Bth2o+taOBIT1Kug+aUUPML2teB5IurwfKDqgwWs5H
Yn5uuCPSu6wpSoc3MEAEE3C879tOpDb2oxH71Gf3Z+t0xUnJM/MsHtxX2SFV
nCHZKwwyjyufC6ON2LFUnThI8zuWtOjB2r3T4x6R8b0KPeFsNOi7jbl0dkbr
0tS2y+Mizyy1USktV0vKxkQuHo1Y4HkXFHibLabzdwa5WBzj44BbwWCO50tv
4dXtupCoP7CZmqUMtBAsORDROg4sMie6A96fmp57Exarjrjpb5yx9whYqhOT
6XzOcS7i2FldbCpU4icCZvX/mcPzVLaAmMSoh7WqSQahhPBaGy749TMBDdXG
/REqeGHvbFzpUelWQF5Xo1zPN0huBD6GpNGrj9UaYw2oipcTz/fAYiDJCajf
eVd01bEkH5xDBdnlbNujKdY/rO1luJHE2GmanGW47hghAnKvB1VC5cQPTmfd
u29xg9CFZq249x2nhWLMMdKvJdKKhdm3+mZALLfkCYTqOKoEmm4PKFxLiePY
wO08oCA9fqR7vC80G5eiBgV85dfAQNhdEz5NTj7ij6I426FYHZxc74ZLDCcU
L04VsXlrssoStnOPvPfUdqFUzFud3CffSQ1/IiyfLh7oEVvrMgrbIHdBH8KG
bAFXrR2SC8bVgu5ze+s6cFwPHw7GlkIwZRqoUUPBkaA+lCfbasbDXiox5H2y
oEAU4DVFzQsviU5/1fhljXK2N2KaTi+zyqUeZVBJo7lpGu+mGcDfligIjcFl
YjYVuHbLnlwARgXYDmMWMpLDUf65flZqeILPBGArFoeP/ogNNIAbsYMsd119
VKGTfTQynIDfAf8Ddjttx9brJvCFrPf0vazdfZoCgZqejPo7Yd5BcK0DKPyS
C3fhXoVMFBCl+somGTpM9p03/AMr1N5UusHY7JOvA2kFYjfM3F6hxIowXLTx
pPv0xUGoP4fG3CbILgbMYdmVo8QVC2vRTz+VgFN/1fmZRAGDbBKUpfGPGY31
NjHBSlzrTi2Z2R2SvCqeWK35dLL8benQBEUfIG8psA+FFnTKmo5Undzc3QKX
Ve5rmWGvD7xNKpF/kymwCN7C3HOid8WlTPtjc+tbIDhjaZj7zyRQpVWqauty
LOMGB4aJB0TrloZdysqEP1dsI0qhLWJUxORnhER2OJXfaze4GfElSO4wchj9
imuRhKY+SAZWJxNkKU4xVEeBkBx5y0QlBH98nt7vT9LkvahheDTwsPKO7O31
25k9rZpX7GgMaINyr16zBgwmvIsw8NXA+ngdoHLRWTzfgyDHlfjg7vDauuMV
T9bBoZtWpF86CaQBmz0mL99/iTNd1C7xTDJA7kUOVaxnf/bNiUexvfGBDNnZ
6A3XbOyZbcC49Kv1Iihq7bqPJF5bLLB31sdQaE4pPAf+Z1I6xkIhuUirtC//
Dtk0rbaEunqWbA0aFg9wbIF3ZbNjVFVMiIJ0bAxyz8wgAC/pLVmg1jjTeC1+
w0pWXfnE4OkqF6u627ryGJHVct85Qdqp7JX7+2NTfEc60n6rUutHvcVfO+9+
Sw/j+K1hYXHw++B7nMNZRxtvBUXnCxcd5ny2OQTLKZXvWRT+XYQ7xw+cwgje
NRHMXWIIvPEEkRTcGEI+yPMsih5jsvV/1LOtudXY9I0xoV0zBBryedMLRVuV
LW9YR4fFfObPov7Es0Ie+iHcj8YoFEHpk1WH2PypZsT52E1pvMr5XdhlS1PP
L7WBfWp+iXQK0BEHdEE1qku3ekbHH6VyZQrZSd7Gwr8p+TzNVR91nN1KT7Wr
RsdSv0oAEur2blVl6TG8PI4NEB+iWNDFBlY7ifZagrsY99/Uh+r8NFxVbUMB
Eq+koWI48v5kl8ZXzz6qdGDPxSu3i3TkOGlupDxwjdKzHkp5Cj65J/2Z90Ez
gmXWzPCZVOXgNxyuVGA6YECm/1um3oFgoziJSNULbe+DPVNp7CXZh8yOxPAE
lWlg7t777dD9pdHeK+fGL1Y7b3W53FlsxkwGwGaE7ILarjBy7XwH5J/9DEih
JpXPTHk+JRoD1jXLQkgGANEtjqwBvqrEqq2U+LLYRamTaDrJaJOrxi3KGEoN
PKFQpCvNiP9L7T/SxRPt+83KQoydbWOxgizR0vC/2TFklL7FFZV1x/M9EkLq
MLgmU8sh5HxsWvTRZatwBEDwOkL+o/bzX4ZK+v6VHe+RmTR/t6ATUkK2g928
WdnzBX7i0WxUpiYHOgqc+Bsr0SrCnvMsXOLqwO7fTAgmvf1aaTZJZTmi2OPr
8c3+z+3n3QuyaOfjGX/g79amSDqcp4+e92rr7yiwPqVq3ztVSR+zeQ4iTxJc
v63/pOaQf8uzodMK4M9ZKuucZsD6JZzcW9Zkg46SBaSMpC9WaGz3KXWMmlTk
2/P2EiDdwFSpCfwyWXJsa8ksI2CI2ONxcO0YW71EHT5RYQm/YhODpXY/D6mo
vG3So5Z35ttFOkeM6a+jucPW/kfblHApJpoxRIKkCf9B7rOM/CjX9OQ7w/PE
cyE/vBcuEn9MSzw/SvHG4A03+Ic3AQY2wYyelDd5cHALedeFBnFwYvvMOzy6
521V+xNCMl+x382YgsjDeHRuGhfU4c+/qDftv9fHVozRFbRjI7wYD/GIrz1N
4x1e6GUt5i4G46RSalr/EhTASME4yBaa4YPSqYrf2PGDOmZNMIRZyZYueSBd
1Kw6VFoXRT5gyRA8FVegVYynZAOgggk/qU4Vx9pvu8hXJbMGJHzWRZLL37pB
M938h6vVXya57kOtKLiRo8qDqpBeyOZo9oUViB8ZubeUsVeWcxsWL/e4kCyD
FT+c5NaJ1BpAHA241OLm9P8Fu9Tm/0BQbuJyIvYvanny+ZCa+PO+Y9yTvd66
7PDCy96zudo1Ei1av3uf7dota/1+pYH/9sVrVNJadVKIln75TqIDNN3alBUK
oHyV7Lg+gU9Uu/UZGTSr60ZzUXYVSolhS7j7OI9oaB4Yo4CtlTN4gMp1nHNF
PiGp5l3/yZb3G81pGVLGsSOFo9MNZ3+e/fMIZiZ9YV8MwpWFdEUOFnT0xPjd
RTAB9419BGKr0M2OWmgc+GMT6uMxoCRFp3etfjCnKKs2BN0Q2VNHi/130KFq
oIc/dzTjma/BDE4HSF1a9QCrnoX3/InHamNzmMUSpRH7XwLpwGzkFMBjjlBf
jGzQNyah/Q1Ad39QVNPpJgp9ogR+QIH3wlsmeRpeMhPDbo55pUQ9tzW0xQCC
+5V0Nkfh1RXBUpVV0Wpp/n/voX7MTQoRCKnJhr1iqJTcOCKrY5wHLr7BqraS
Zlc394PswAqliS7vuAJnkCKtT4Lyo+mmFMuwqibX4v5EfUva5jLXDjo0L1hC
Nms9qJiIsTSsQpsiuW4cF/Ncs8BeNilhlFWNi2Hj2alOK5oIo+EBPutwvvzp
Vw1NzzqFdoD0V+lC7ZiM1VfTOThlKNYs7x9IvqK9lMoeEdnpKy3p5jES9itH
tTMvQ6An8Il1SZ8ne25/n/Xhh9DpF+ulLKZvUShSjnjGoybTgOL3JbnnhakH
6ixndTqYMjUT1j+CXxQj73X7V14Wa8WJQfKwa1DOLz/5c/hI/md2Zw24a1Db
VZfA/S2AnZ9PFRdkK/N4k6zoAFmNYYQrrGOaR0tR+Bcxitjov959J7JtxnQQ
pwTVS+XHBtbTUqBgnVoV+qvBV48gn5rbiJB81fk54Wqe8EaRVOccrsDgdyFd
57+bEJPCKnEQdVCZX/i6jQ4PMXezGYqjnU0WtdsMF4emOgcVtIIEXFe/pi0X
cw15N/D46EXDXVon9pWfmP3llrHULYiOR61W7VWiPiNWXO3Zm5i3ToRfJDdT
k0fYQhtxZdUrTxFK2TPli8IObSZZhFn2zZPNxRVIQU1bpXtEOhXArSTyoWRX
M+nuKdu6HSldek3llw+BgP5x6DAqbQbYjwak7r7UReOuZsqaGUBTk9rG/Fx5
ajShvCYuQTpdmMCg4Pm3M8lorT5C/95sgA+0ZxiLVROzBVi23J+2XQIXkyZS
gtapTz8vIHSq/sKhVccfedeJp1XpBosv1VYftm76NXia0HHPKEMjHs2rkU3S
15PQgQrwYUk38+tB/f/ACXPnnh1gqYzSheXsqgg3r6i9J254ZL9w1yk8jfue
YtcjybS1hWKNKJSWNdnXcSM5jk1188ezc5yveXI1IYCi18vr4Q5rQrB8b9sV
S5KrKY18zp6n/RiqGeS/pwV8BDk0YrbRMf7cnx7uWc3ukXfpnCL5BcGJiTIK
Ro9e3xqOZnX60p00vypz8eHZDxi91Q/SY3PdVKmzh5KgsWP2YUMuJAxTgCCV
KTucL87GXRo/0rgM34A9yLe+SyJwuHy6Yr8x1k5So48PxabMeqyAkr5R/Mt0
d1FmxCH+TnIj1KbpyvwjeKONDweGbP3f2CqFof42CbY7WNTaP2Y9IAxF6AgB
r558+zD+znHj0DIGXNWIkUcLFNOh0qDigAOwx0KNM6Np07r/I6h/ldlzaDrs
XyY184E0GZpwq9ucR5JKhs9n5j4L3t4ro2F1oMSDUCc9rvKivIFF/VKo8Fak
dBgqCwjwiX3S7Yyf+XHak5wxbogZVqTKCJdNDtNqhU1P4uW2BLYUVH4+dH2I
fzCkuavYFLh14wXntABJOKuXf2HUX9h7X0Zlu4qLzthATozyewhIdnYhOuYO
6P/5+Wzgc450ZUi5g7UkqguD5dVPc3t7hzrK8X4ho9JdAZVwEmVYdbbIKO9S
fhwzuFH9vTUUiFNtrY/GyoaOhJ+pA2H+VYzDjeDlt9uKx+Q/JsaJ13ujkr0j
q7BPCgxsICB7thribFSExsQDpszzevECwz4Zi/PEQi5RzFlksMHoSZ4zIOEf
KSBXSUd+cyEWIj60mwvj5cFYT7smiMkN5Ntj1tM3J6nW/RwqZ/lDF8vOv0c2
c1BvB1BysFNP51ClFcBcnJGXatxbIPV49Wcu/l4LrdHrYWqwpZrv4oHy9c2b
Rir/ShC45XSKBT//UUDgmg+zOUydIuEBQrcTNjZvb/0MR8o66LsrqIUMvgq0
4CTeiEH48AVYIq+CVouA+m4aDkR2f/PETQLVMfAtpQn4+RP1sGI5QQdcCABo
FNDYYWT9huLmzFaz+R53EoVfFIE7hkT0SgtsP9nV+/1PwnP8vfZY51E0MW1t
EYCSeYVDfSsqWk23c2/uSGjYiPaGecZg49XPA/+plmM3m5vvxvifzSKxvETq
bw74f6mmoCXL+BwLojrKvOA3E9eHHOq5d3O7XluXfZ2qzRW1hGwN/23b9bx1
mKlP0f+CMfQ/Rn0X9gq2brOPg05En1oXdvItP+Rjy/B1vOKgg19N5h244/oe
HVju7/+jYi6Lms+tze91zoGXZXvGDl8l0LQGDfWrO4XHxYF+cJIwOhXDTGKh
12hPkYjlkYq29CxqAS8kSjShxDh223sKKHwV8CErAZReW8RV5BXZIYNPQzGz
/2QXh+WpXIGFb19OX3IgZzYUD1omEErzmigw8qlWcRwa7OmuL32aOQU+bjeT
eGWls98ysccyeapo1+3Q1S3JsaUJDgL6hCHvw2AB7HWOXOf5AELHM52GqGRT
ZKGlexVB22301UD1A8KO0yhAPI477gqoLAYR1ozQ03fxQ3CX4elRoD4k8Cry
byMi1C6xESV16d2s7PDWH6XUgSn3Srpp4JywRC+3YK6zGe60+jTrZ165Xmnm
5A6wgWUHzEptmTnTcAE1uiNWAYdDHCbzisvBBmAsQ3iCtPzZiQOox/0f5CcV
QUI956tlLeu8+/+GUAQJ+PfNGlz5gBqYh//h0ClU0kP5+axsYhx6YPGQECym
gYYWdU4BA1E5dWpmpRfRYYB+2VF5DbQskarxVdaw/82vYLuPoGMxnHU01BuO
SniI8w6ixiHsxWaeAKCRHXtzo0TsaN38wQRb0SX+KAufWY3aHDKuicqErDAS
pwRo9CuRNin19ogdEMAFdbQQInOa4e68fkPD3ZG/sL/0Yp+FARBwLjfym4iq
NK3nbwKo/m+Hhr/YMkde0ww+4f98AIG5gI0nCnfNx5R2rm+LVDidH08xJjb6
GFh62hhYHRlVgQt4KS9mSIPv4iO5L0pf2a56o9oyfjvOvy+sUFjxTOBqV+3l
RLM9B5WKC2oAhNgk1FyKn6B/tfnO86EjjyGm/be7hsypVyKRCcYzmnT/w397
P3lHbIfNYW6RJfbSIBLe/TejJNdGJAsBDp3CxNB1pTB8q4oN3TyclhE8Zo1e
fcoGO0VUrhvzHor6x0+pkUzKNLXEAgB7hcaFfrgueXJKDLk6yYLeqT+IvR2n
02lsYPnf7c7qWVME9gZV7DyLu6rIe4+OYkmhQSIJ6h6AxDETLay1t40aK000
DO1I1/HMCesvHbDULwS/SSCIOpJ896mznGZ1ZYaFDvWlKkH+Y5wO7asEhNGi
ZvF2VL2jTvMh7aovOAa1PCpd0TU9470K4l/+627T1xLif3ru2txg7yNqlAw7
FojQMVtHdNY2AW5GQM2fyF7lJlsB/jB33DVU9pQ6PrkU4/3bOAtL91yt3tww
Psj5YEFLIhpuZuiFINrwro1uRt1sy5Q2MXUi7Ee94R4TMd0ARGxCZCpQAIF2
2OT4l5QSi1KvLp7DjmzlwEAgwkFfxzil+/Qe7cdqRtlLzpgDeI6IKSzMBnyD
P+uyrAdG53eF0XWYLUBLzr4NhqjnUTnbK4EU/YfyM/CoeQ7zAywK3VQfmxeN
NRbFaYss7ofeeAv++MOQKTLXErvIAbgbr392iDfI0c2JNwR9UcYzYDQmTTPr
VHOahJResDQQWxnqwKMh/YDWRkhlzSesxeBUAOyNmwBrPQVMKw3q9wgoy9QS
lC9Pa6PF2NWgzdt5/3ymT7AiOuMq5yMaI+FSY25eiHzIz/1GMLwb+2ZsZA8H
udVyyU+1XCpGIzL/5CQk+Z1bHrAxyjnQKAq1KrjrmSY0Zs9pjC+DTIpU9W5h
0O9ny5jEGARHiMr/ncH8qzCY2cSwBC3I8i9cqfairkZumIBSnC8IkxpDh/Up
0R9tHMVgw5+3YJilpiUSSEahd9IW+SrFlg6N2I072cvP1xHc2QmcUaXvYGQQ
F47WGSz68qPjhdP6NEWGRGZjzvdnFZhj+l5406wnjoYfqXMceGVf1i4/5QRU
zB0nDB5SVY05Cnx2bKqBwplJA7AeYX67SanmDwY8SnZYoqOXU7F09m8fU1p0
Fl+IrmgJHXFGF8EBI6JG5tnzUMwA/QH/XQBrfG7XEZfYEHUS6rElkYg3r1yC
lxXPxE9np572iyCj/zNuLrAT50MGHdHIZwMrmzupB6yfHetldUpma5xBpUAq
+pvKVHov77sBmpg+Ch2rkF9b2BpEIpW9vDra6xI30OoHbKI1sXfjkgO0hKXN
o5yytxu13EIU8WxPzgTJRjG4zRT9PG92ywTZhH8LB9QPDSmvHCZS1wRHqaJ3
AhoiOZMIDQpsE7XddT8dKhahctFapd0uqb4o997fiOKtTPBeMjrpxKg4/EuE
fn0PkDf9B6iP476jBzIHfM8MmdTkYw8fXPuBi+2iMg6h5cgVgt+svJ/GJ0rD
2BjSc0331NAnlKxpuzENqmVUq1LA78aP7DLkz6iK1i6hEPN7KBw+tJwJO2Wd
RFa2LPM74ugvocst8JFf+JhPxBE7uePQrwtHBBsp3yVl28BtQ0otGPFz4m2l
k1ufUra07MMEI2oEHnQak2K7oMdR4O4cwjJVppWfCiMs6BoGQxWmcjEXz2CW
O8v9uMfoHamcCucR0688FVsfeuvp7wAOm2XTFLouTOrzzqlspu0RMKm3huzx
ILYenAImgQpGWXtwuMY+Zo3Zzk/JifGkeGtzYHg0CSuv4LVcsI09UivpXmcA
0Xbv2LAs623XcfOYvz241lVXtuKjRIkc5/nvOc4KVFRxHH+d4118VegvveYr
FAQCwkfsw2AoLCBBjhUEHTu2VHhy6XqSk/13MTHymxKrH1zXJR927HUskC91
3yyNiB4iC7vlc4ZNMhqtJxWyL25Pudjke4xrvVps81nzXJ8vI3yIHcyvI/qD
igXWVafhr/fYl9GQaX9FKkUHK4fClEyMOrPlTqWl388xswqFZ0eRldHGVDOV
ZnXGkmUX8JgVIXr+sUUTHszN+lSPnUoJmcO+lx2xJyh3RFha3po68UrXaj7T
7ySH3oFBoQROohh0AuCfsJ8zeiaEd9+eliBe66TJGntihveSVu2NwXLC6F/A
/1sp0LOL8LnCi7Immzcm1SM9cqGYUOeGHV3bfWKzBSNx7r5H6GaogfXxVECH
4oMPQ1aaqBaUCbkFInzgxHl178jrCJVvGTIcqAwhkY3yvFF8xxwa61DeBzXP
OQ/4la6Xb09n5obx/JqJx0b494ZlCFjmFyCtD+VWliojRVMj2AJNZjF0OAba
Q6iRMSWRfKAaUrGge4lJzQWgGrkNU8loINvuA2aXLsTUYeJl9qmIqeqPk7K5
kDTp0npwqx9wPTgppuKe+QMu3vkqcZoMRkA+HBxZZH9j7ogCzhmvDwc/ZMYw
wKWtHb+n5JDgXtc7rfhmYZ2gIAjWs3KDpecSL++tIML8F3iuWtzKMA2v9eme
DHhv0f/E7MRwopmmWANanFVgbI7lS+reIQ+P6z9KX0g2Now1SmDNBw4X0Lhk
4TDQFZeY48GDeLBLWL8whQOP6n/MixEW2sWe8eU56n9kAaY/SshvscWMgz38
BLsuSoRozeUAVd49A5tSBE666nEbyHr8HEMsbGPfqhfRX2e7cUq/JUCxHbNI
kT4h9OnwQLU+crK+yrZbHd7+UULdQWK0tq2SJ/s+XKlmuY7q6c1tOGO9UgGM
tinqO/Iy2QINkozZwt9vxFh/WDPcEY+H/9MsyY+DMeJtagb8pE1UwzBGdv/a
f/0Ya0NQ86LxEnMfvnBN8F+pUfG90QHZZ+GUBuUKJsEmdKZz3yWf+DonY0au
4UimRmfzBey4YHvNQSY0zZv7AtRZZW/OO4C6kWwgxbCbu63VImlWiBxiiANT
fG/0tRDN3YwKIw04DOMFUmS4OipcLq3T9woib2nyVP6qJzVTxbG3zhJOjsIL
xjtu1RqWMUIQVAIj5jhSDjyYg+hqvtoel2GRdaCm7nEC0J6Ma7a1N0077MtX
33D3FeoLZWZYF9HF9QxykoF+QMgNNORCvIuYYVovpI+HQfNQ/FNjs5KQTEhm
uKk7JS0bkhHfB2PEUNOBG9HKGYPlCXnhGuXobHjmmzAQryHkQkwiWUwIXXT+
YHdrbKUucBcxv9pDdQld2BXlUPCTdGTc2fxw9c4F6zzqggXfTGZggVfG9J/K
93vf///s4H3yoIon8cH6gmaXqa4BVY87x8zNRJaWn75ceyBHYzLP072j1iBU
0NESxHX1XNVEz9bcEBnSJWfclVqJfEMoaaiN+5EKxeTkeXatlXttoGgyMBIL
YPjbfVp5qorpGeUeone7xQsE03Hn3iIMux1r53yzpgQSuCAVSxIsekITUksc
p0VhL75iTGMSBbLabOCFPUBQHGrU8WkL/gasUUVwQQfnHWQN1ua8FCjBz/wU
V/H5CYP6aF35cM+s2XWQbnCspQR7+r/OF0eKJmDjeqVd2zL6JZRuvz/IS884
OSP/GhTHHZbhnOzl7DDu+QyWlDqOxT7+GrAGKoIxMo/fMru/zJdYpxN/WuP/
ReNOTiMu0tlk5lpQXqYO0srNkdzdlSig2fUFpOWgcPG4iaaW26j4eXjCN0ji
6cTvUFBNBd4aOm5hMog6DeE9H7vS25BxK1XqvW+YuDiO9e8z4z3A6MnAKV4Y
ubrYLyoU2IcACBMq+H/HH8484nhqZhKflg0Ez+TWLanK55mGOxy37BJD8cSq
tLAX3BiqChTJKB8z4g8FuzOyOb8cD+mP+i3B0sLlEVbPcM2J+rlEluQV9oPb
M0id5CB96QCG9zBBNmeEciGKgTzZV3ZzSN0dgqpYmw3zYtH5JCfjmAECP15a
SqcB+ksdjJMJ/XUIe+403okaA6QzhakJPsmL95YCO6lIGjPIOTjdQNphg0DZ
ojU085Rtjkn2zn04/wS18UA+laJ/zseHdr/BZACikXmo236bqxfdFyaJXJ1v
6b+rY+6UlecyqIgUBKk4/lCgavs2joSsUhN/9jrolJm25AqF3sJ+2qiczRbD
S2eWMnGVYlptt4IsIwjkJkwSi4moKzBCheBFGdxHQI0jQQ5pkoz/KMwTUmm0
fvJEcn14IDvEeSMrumJa9SY3l6yw1wTpHWcaehZMv/ZHclYdLnA3HXsabw3g
Kqv9o61L62Z2J1CmYysmducFbgJlmV+APjXJtbLj3wZYy8fc9mfinl7cIzEo
p6Eu0zwQ9qcMzfFB+AkwXZ2rEOtO2ws323+T6bJo3v3KuARO5VWWo1WrZUfx
pvzDhpIjcNMV0jBhUKYMgrwA2xKB0977xIyqmbnLtopJClUdmbchYYPi/gHS
adLtHWGy2P9Vru0VHtXOVAXmJOonWPs2UaoK0M60yqdiY0PsCSgBtu0I1pyO
iNHlaHECRVvbl5TwdWFBejcp5tPpkCyZ0JHPTMZkm6kGMFDQbO/Ev8axRIDI
e1deKObOO/fjjb3XYalR9ICqwVp0alDmTxXC8LYdwNXlk79x9rGK3Zq99k7/
M4opQ4LR+Sd0BMaCByQ7TF80ph+x46P96+ptQUokMCmoHjVg5dJI3DydOrP4
3OUiJkFu+HKQ6W15VmqT0EpYuZaYxRTVZrZhs9I49WqXwOlAvbXdpPiYHHi8
u5iQh9Vd6vVyZKCa6KadaVtjI2NFSc7AROIXvjamqYxSsGqxErzaio9nVO9+
alMN8qZuBZkJCSoNKAcEXHdicDg26twn7JJUwLHVucVNE9oBm8GzQY6uorfb
cO8rAJwf1DSVK8CraO2+4IFGeKgH1bMMyUrHRDu160YVrVjsCwM8QLBZmY9Y
V2GdsD7Jsn0I62lGTOIYvBWxFrTkru3dNdtl+QEG5vF4BlmcZmIbGtwT5Yy8
JLXz6h8r2eTWB+KJmxwb6uB9IAXmepAVyZ43s0jMF/Bgy7KiKo+3KVu5DqLr
WsS4FCgucjlXM6p/d4B0g6S56b5j5Bjirsvr/KYICbyBQnmMhjb24VE2AMm9
o55yIRCOFjxmf+kungAz+UR67/qrDt27hnJkFCSfufNqiPlI4cfgLJMYEhCR
vrlAQMZ7AQfbt3G239GpJmpHMGvGxDWn3x4tXBZNKBWVclOSnLC7HdFHfDh7
j9zzeYRDzUKUTvj5RIkoSEHbqYJRqB2738yd40YMhBnlrpyu2R9ADwMqIhAe
fQWQhsxwPx3ZiWOv8lENddNohW6AeZ1gjEMWIAQaDPZIyiSwMRWZgL9S26zz
vFiRXhrwnC6fW76RB96vHv343YzComhQWMd6GBqlvZi9YhDUxaa8jjVSfV5l
6vTDDFEdjBqSCzXHHXnAfUn5mgTmM3fCAKA7BVCIpth7cALxKNRfn22aS09d
F2Pl59ZTcDCsR6eJEes0lXEYniruNbVOmzp6t3mXoC6VE+jPaVT7TfmaZpio
Ve1UOjCD+9ZalgjMR4CFR0yJ5+3mMpDk6uCiN7XK/nHuWemi3fMzC8iutvha
hn2adtrDdiyYXEx0/qKxckgFaVgd238rQiuVCFiprR4VXgtaF0X8MaB6uLFo
lcr+WeaADQ4+GirJuD0z3GeqEkyK9c0KEoQu4iltBULlBbbEj4Cm6H6BYaxC
maFg1Xm+Xuy3F2J46PI05hcGpujW8PhgKDZUk1bSBycuE+Wm9PIPHDdQ2a9g
z6O/Ry1iJZAMdKcz9/vW3mWu7oHbLGkJrhn6aaoOyjht21YmmXq4bPUrr6dv
/+vcJGNpvG6eTN7GxKwJVj03gmU32r75qvnnQ3LKEdwgRIfNefFd4R/zZ1tR
2onNBDXmoI1BWLypRopizCm7a+3fbbWOX3+b/l1dfRb8dplQvUwoooIzim16
y0S+iIS0ivMIs8E2BsRGNhgUcK74wQDpLDwIXIVG/empd/6cQcUvKPj8YbIT
JW75diEF+ufPspKHFwBBhILrRAPYB4rpyB4Ci28JcIsrhZdYa3BWCRNSrrXa
VjTDQF3PdonoTxGj+tPBqUHBiAMiX98FDM0XXrvVbxd834aOHrIMi0Cf6N8V
zr2C8Tu+tfSzDCpbueNTsan/DVf9k2lXdBsNQBru1MH2OYRwh20cEcd/X2ku
XcoiayG1i+Ukd/SSer+8drJwDMHS9jkDoKUIyvOlhSgUKUjTtbNdRf0Cb9Oo
0z3q9ODww9Z9iFcmCeAOw3i/su+/FupWSHGrkNm2kxu/4k9/qbEwdU1K8+Ul
xEyKhbAzzlLzdFuj/BKm6ovXYszEOPWakYJLSTH/t6LVRVgvJyOB0zrMn3Ol
6q6OVm4vj22yEgO/PQQ6xDYG1WjcUV7lfe2mm2lI1Y4H2OeJLMfrgJzcXN5J
AR8xsobBsUbMUmaB++qdc+k0YPV/ZtYsVQTRLAgU0e9+7BdobK+NvXZ/lw2U
wEE3S30GIDNEx6Wf/NcFNYHr7H3S2yHup5qS4Em8vJV+ZJT1bQsCY3LtZpxI
zG9CT0lnu2AFU8W6u4DOvMYy56msmK2CJOxysSlw8kqgohlp99rXD6CoNYtH
LYyl1/FKsmRqLZDmPME8RI1znaubpNKVIs1afm8QIELgUn8AQbjiMAvD8fG5
We2hxQ7guBMegcG8Sh+jfSUY308Maf41ngvDB2vfBK0PAGMS5S6rE1Nl1Q+1
g6TaM/J0FGeML8ck6Z1+Pu45pSjzSaorH06HWrqn3Z68lQdzhyFiPL6x03gF
8ZiA4CP9jmKY1qPDFI6bW0a3cKuwUB1UmiHU3CHB1lYQBuqwDONclfqa6Hxd
NXunUXI8v4GYOfc9iQRggZR1NnoEcs3s4K49eY5AJsoVsCCxDjBjKlzkukok
kt4eeNPA9Rb9JYhbaM43ya/73pHTACOog0eaA7T2kPGdpzTgvQIAqrKK1FU5
aOqzCPGgP7am0lw3XwCDwmsZyC2pw2GKkR2uc1sB9BvhXUuxsB6WZZOymlkv
uC0YJW/hZDKCu/Ad5JER5/esgd9Te+8o0k/z0dRgup2YqhD7GixJeHBMYKZC
wbLO7WE2phIUIsLen/lw0lEmD4BXqracsLHgEQ2nWqkd7KULoattRnDtmwL3
KzkxOxCUySHU0a2WFK/Ebk2VgcAsZsju77tVuNcmcDyRTFe0nsCqoyTy6X2i
Yu2FTrF30BTxCevBiNm+tn8HdaOgHK7Bla41lwiJqrcVon0pYdDENNUBwaWy
hU6Tvxc62N78iM2dYnQPxvgSCuUnmAtBPmad9LjlEVEqDqkgS0rtLaoL/RGf
hohP4g4fHz0dOVCWWRQJjR020aFmr4T1oPtXqRXoU1GfBmLssqzULYlUlwHw
tKyU8J1wsy4KhOVUiiuOeSOi1ptchv4hgGyK3TarH8MoKIgR4rC2o+OED+Z3
pTElFVTLnFWroXPyaZwzzB4iC4ADiVkKQZM5rpT4i4Gs9e8q7dZtigN+ukHT
owI+aCJq/EA2dlwxVXZSCTB5Ia3S4S8jgBaLfKk4/ptLLfSmoCVNuXSABbQf
Bddhx7dJ27BKvs72D8rwL3VcVpHkp37ld+vRNkIVE+zj9i0ahZubm/ePB9AB
AnWN4mUt2mEWwr0ta8E2pgTf8nRLYtEQo0C8wTMNfmjCxdCzIG7s9GGvGfzq
CKRW7WYkT2DWdndlLPwEuPG7s0J15MQ3UyayqusPRsfpd/YTfDdh3tQveCK6
wkiyt354/OTfYmWUJRJZDVRmfUN6xVp4yJ2FsqzjXOvRsx7bIZCjd6Rcj7zz
H9a7A0MHgbY9+mqN0egoEqtHV+LT6yWc0AbDt7va7WcyRwb66GxUrqfqA5GR
vmlDTafVkaDWqmVcIznrQFG9a22pqIwU3XvEPB8tYeBvlubzZPWVxNddalI2
cXz7HdTSbIr912dAKaoR7fBUonYdUOnSb+kKsbloX4M6LroFoSNxCpx66CmB
yQ0uHiLUW6UW5V3UwfCuDQ7Hp+d9v/Ffhc2pn1WMuDz5H8ILWaH55yIk7kJm
o8L2LPE/RqpNfCw9KQtKSrioJdo/DdLaVQQTjR/+0rBo5b1ulXfg1Jf/GNKM
59x8lZJk2/jUPRGiE6B9FTwC3o/kCLw/Sz4B9BXgDXmb/mKHBESkUVHvS/mk
CCHkESb42ZcTLX/QYXWsOUByOdAjDfZJqBXM0zPZKHH9gL2Tunw2om54kDu7
k8Lxi7Wx5MLo/kWEybSPN3pu0jjeNkhty8WG/3vgXMlCOiqgEV6DY1EBxHLh
kgc7MPeewpNl87a/dl9FeNK+SdhmtQD7LVDAUEPK1uG6fGNaXYSlSP9VOxgn
DVmiZOVFQJe/QdQRZAab/CTkDCR046QPWv29cae9YdFNGxzPcTh3z5M2jKZ0
t10a3YSNL9DNMhZXFgP5fAD+pflkcxv4iwVNN/mdWhjmtaOetln8AXCFOPaC
9X+BIu1FeisVJ//sRFfdW5CmzP8DLLxHpQ8Y2vo/TB2V3htcWS9TNBcfyhfo
invf1W2cMWTojARsAgR7fmNWOYa6mHic/lY6h6V/cSQIS16T0Lhu0Opa2ben
xZcJ7NRBNxBaR703HQiRCpEoDvBn0SqyD9iaSAgKIiJGQvWImo3QS8knLXK+
snrrBJqWx3G4JYnQo9yY2mVQjjXd6HVXkzVrioMJlBZy4+YHyvCvb4yK7gKq
ZQ480W8njGs7e+VuKtu2lKSvTIt7fYH8rbyK9GRKjx8aj2kKYJ0HBy7D3tJb
aQ8oo1qg0UpG1coui5TZ50VklgWsSN3PnJjawE7egY3TRXemXEW+G2+m2x79
9k8TAg8y8nAO6Xq0FQpLiLFFBNxSLMDnAo+u38lAoBuiY98SAzAsqpSYBcVW
gaczFnyoc38QBEu1HSdLg0h04iwKo2DWd9kSRA75Cx4SIMSa6rSou6b9xLL5
QjnbN4a6eOFa2VBuIGjlFLBQWCOb80FuuTDVpBnSGjY+vpzFr33dYwhZSKRA
NZJNF0XI3B9IONjmkvjW5lwqDs4SxLzkmFVM5OuaIFiX3CaTW5Rz7D4qNw23
bmFBL59egka5tCxd0uaF2+GBIyNxuAhpkH7ZSDrA5Sob+sgZfDFHjFoo13yA
dxo+q1OvanaVWStM+vZyO3UmlqISjfb5+sp12C+DflUGmhcKWZfZyQQfl3Pl
XBL3XWMUY8wYe1PjQo7BMNaRTt6XKQ/fUDECCugjfRtkOnrh6uZxC4EZhVmj
8G2eHkFhX4uGWYa1SIZ837Y/F2CKEqQjPbBmCeMz98vPSReG1ClVJ7WIePwj
RlvNVJvll8fDIVWObqO5zO1U+acjsysuntSgC/ADGB+89gQ+FqlqsELwaYdo
L1c3UJAXd74PfRJkvHKtAmdtjbhxaUiWuVwvvPqXqZZaRqjpvSKzda3/dNhl
7ZpfoRHXf5B+bGnqIDd68bdKzMpzAUcy/bQNYyL8alQMUiECFAz3CN63bRAl
DT9MYLio+fFrcwCvuzXuR9OTVpybHHLtlPpRzuj3QjJm7Eu9dQqsWXNdw/pM
Xkk0EQjwkl/TejtyVrYUPgkcMYchKyAXUarhSoOo6MzLhy/dKl3arOlTO4S8
PXDwPglWuB6QLo4NnuTIP5HOAdX5/4kXZZql8hh4Fnhph7VnmhOtegs0fVAg
+JIdCDCV89aMKAHBdpxfxjU+oS+wn4Qpgj3cfQ+uCmjkpkeuYpEghahjh/2n
afREvdVHOXq621vdIJ+EGzeCQ2dzohvjH9wcSb3yqq3UMXq4kg5xX/vUHVQb
gKsjMmROt3WMaa6uqxh3L1wapuj0F+8dLQkcKN9Q/xLWJH0BD/uQOWORsGVQ
Lri72SPr4kZdKBnYmTtVbuo4KcN279xex0iFHEOuSZpz79autHgRx4hj9jnY
7ZcxNpr5EFpKeS10FqAhh3G39GguQCWxO5MmRA62KftLuwNItYuGA6X8aoww
d+FDFFA2GWsrPWpGsyJtqmL/HB8ZT18TxJdV6b05i5/AJjS8l9RI0OLW7sfg
7X/JmZwJRaY+yKS3IvZVKzeYWxA/Hu2mwjsXtUCDvH3rpoyl38YmkWecgfcW
ku2jcHppGLcvjXMmOStPvUUdEvOWh676vaJcaou9E1w6j1XSQll6RpCVO5M/
IuiF1DKqx8Omlx6u81mHwCq62OECyo3SytXZqycj0XxOAOo2RyLa4pGFvuRC
LdL72OinFiDyB8qtOWe/29fgjmTC39y4O9J98e2ZX3BHDIWI4QQvQxxIr+CP
GYZz2Z7UHuM+j2ufe2X89Prjk8s/FQ9GQORjkDI75huPdK6/hPTGYTt73Vqv
esB0JE4s0LuYlS8h27iO0fIZaKyqNUkSe91zZqRdQWbFVXlIHM6HKl9aaYv5
smqEeXs68QHPiqXxi+wS0FAy3nxrdzTg0pFIwS0VspwLAZTWWdYRFyxbKvzZ
gS7so2ZHRI0mNxGXxyQ9P/iRsBPlenR6voaM/04qWg0Vq1c2IpZkoBk91AOp
M6CfT8rPUzT2u3jX0avYbxg56m05x6DvGvmwq/0XI1yWcIkciYHgAeomNcx0
YlGHoST+zneBZtw4W4HJv8UtcbaxNH0J+eYNrSE41X2vdPSRe/A3a9GaqDdn
0DeRruCd2uNsaaXxETBPo3ax4++OFa/V/yzo4a0zpzqFxPnYvZ3XkkRRKhYF
MktHg/5KD8VAE1YhefpKHMi9MIH01QVbYFqMY1fzMAgGkuypNJWGDxh+kD2I
HesGEhasF845WebLdo6rTkUraXM43aF/lRjY4k+E4d9UYbtWGzl4H/sl2ohH
/yfXwU2D1JYar0tDakFUWrX6CsfFFCpE+m3PMkwmRyIpVM3uEKEXAPAUh7yt
E/td82Q0p9tW0rfU9QpahrDLPcoM2FfkeqpqAVKFx863cfAlNX6DuOHvEadn
r601bFgxpZkMG2sp0jbiY3QOl4wJdZmQ7MNwJJqHsQI5SW3MCXlurxkpK8Or
AL1Pp5n/JftR9ECjIfzkD1aLgciFzow1JBGgCI3N1t0Ws/Fgbyk5zaVlxhfk
mhyeovmWkVA9ScThoBWEa+aAuMTVTeKd4YB//7Ny/rf2nXeReaN4dZUqLf9H
tKGPtkzbrUt3kk7EqBwqmfi6rtU8rC9ZtoILiC8f/mP+iapfp7r1wMMCbumN
9uqjHj7kWu1pNM61OYjtwblQwwdKiRvBWgJoqrqj9eqrdymqSsBUYw1IOzX5
Q8RqaojJ6asry+S+fgsj5zNXi5gvwmDNoKwl3W2i8pv+a15Y6KSrkNoegGzo
/2JSbckyFN11DqKC5xm9pEO9JyhNIhd1qnBr4oJL30Wk5dgC1Pj3mC8bJxJ3
N354I9rmaMfHE3GeQcGnYFbuiHxxiri5aJGvIDIfvtMrpEoZsDOo053oT4lp
zICRIYKWoX80AhIe2Ry7WyAFsuMeuPDtNnuNK8YZmIVA9s9MPo8NjbygZamf
nxluwqdAlwORhIIOuJRaUaO7WZEC4BTszybpI4k6L5asi4D9oKoIg3n+bAFd
tTVFELRwV/zfrUM8LgdVHyRoeQL9g0K7EN3T2eSC40bT08HYqvSXLgD+srHi
Z2IRqatlhLUDBEsANsimj0a9aK3L/7KOKtJO26jA2PHNbfPKwJ32utHup03U
EuVuEMz9b0DbbLRBV6moqhsORJghnrgEjEBhogHCqs1MFtY6WjZWfygjZrMb
dsEB5W71Ot3NZ/Tmtg8GhQ26qWbOziVIsqR5JUg+jNAm9NB0Wn91C9GQ0d2q
q//HR/dtYTxtz6W2gLCcIMLqsdTJx5U4pkzU44ffFIUNvN6QfWRwHGxo8esr
UpxPgCCrFaBybVLiYXGePw4iqyNlBP+jm5ICJ6ExE0uCIijmQS0lCVol0J5Y
LxmCJNZxpC4jqdsvLlXF49zPTvFZZMOpJNEK4BvkHel1a9N0pxkRhmaA2qfi
tBToxQQomUuwt/A9bW4Ar7MLpKS2DSIJuuTM+gAjC59Up/GETDfAuGuU1/TS
M2rXaE3knCXMtEHSET5dfXWOCDJ+696flyWu587pbJecp1ejQF8cGfvOhWXX
yPTp5PWwZtQj8mfrE7YREweYejTY6SH9PwoWAZK5KChHW+l9ILtzohbkpeOf
1Ht5Lx6U8+iLQgMBNvAE3SE3XvKwUAw8vYzcIjYf8fqpL2DUmzQt/abNmgi/
HzjQ6OLzb5paZ9aVwCT3NNKLeyl99e9XABVuI5jZbxbEON1I8mR51jRGUQM7
sBn6LTRPl9F0F0rrSaYs8BSdUuC219CJ4lhCTPomJjPNbx0abURebsL1pwlv
eZPs0KSlaNcRHuxZTofxOasiRJlCPzCdvyGpydNAlaDhloBNDs1Zo96xzhs7
bwFxbuBLlgj0AFFSDZnE/euuNV4CIjrgYkzuJCijTo4oj71mIT3Y5osazdc2
r2WdJs8gMJHu70Fv83GemqFpUNqjT/83pxIliLcdWRijE6hFmG4OXuKKUp9g
FY2W5eHDmDk77/1tX5d3zItOUyo1uhPOGB66b+RbdT2ycbCjc8xeVe7IZdKo
1oyuFbir8AlSjvdhsscze6lPN0t3/4BH4H5wjm7fZ1pc9yOtHqtBrowfzHlE
UZtsJc0v821kmULM+KkUdsOt4X6KOM4Utm2Yj/Ssoxg2CK+JAcr3DpvW0gGO
vye86Q3a6Aywm6TiWzsTDbEPPmIYphU5e3tGKPok8N2T38vWv+VUXqpRW74W
oPCYku6J4c+Bcg2xPOGeMyUKo5tZoHPE2A57TKTNdGG+bZlOX2sIcPmCNrlK
De2y/6nipNBRF34jOps2Klh5Gf2N6j/mGUxXgWv2vEceplS+DdLxMxJAgc3s
7RotIWjkbTJr5VxBD0jth+6nsxk2G4fwXarWvU0Anh75nJ94vR6mTBdP2xPD
1qIpPD7O3m3iww7AIf9UHFxwvwKGVWC7jdawuJSqydyHHXdtg1ucNpZwgRjO
rV+X2c/u8oAGA7YYVuSFhbTZv6G0H/FSKrcLvduO1Yz2htGwI43lu0DvTnZd
GhWcK/kWpSLrgC8mMl5SbMmpJ5JjhPz4gkKN40VF8BGI1gS+njqLPKOa27fx
WTilzINmB9FQoGyYptxejU7rbg3+mxUJ2VeVh2fpgIr1pZC9ab+m8blBMrNK
Z2gr1KB0mPqHVYuEfw5SAaXh/wzoVytNzM17wyFSFwglumjUGj6XRnBWZrwU
A2A1oM6KXlaO9x1sAa3eYY4arE9PZC9z/Ubz9e8Z2JxI+GXv1FGSvoIJpIRK
it1y/B8f+58O8UdJ3yuOYNRHaT9u8VerEzC4mHOq89mGJUgbvJTgBbvRGRIa
KjYQk6dtIK/ZX4v81gKWztDAgPS9KfNjpyRDAJ5J/51AiFW4MjsEjF23E+6r
tR5IZDN527EHNhdCoHT8mVpbDUm8sxkz9humg8fBU9jjcHRgqk/VXhFx1Pcz
tY56IX4xtaJyi3QSXkSJObpQuZaFG+GUF+Wocj9Y4KHvrGXyXhSsvpnR6mGV
03+yAFxOWoWhT3x/zIG1M5QQ13ImNKofJ/zk+8C3D9ixgOL8ikDhNhtOYElM
fo1EPzXeb8qOJ39Urla73XelH2FmK/3jdxUkChDX8DYzDQS99G5jVOGC1J1S
Au1rnBX/+vJugDxuJEMUm42ZlZZsKuOvIm8c6YzYRAzyutUv8QQFSkuKBDHH
tmAqSqjh+wtaIR2cUUPj3o05mQYworqrdN4WTXaPLVsyC94wSzV/MGeBLpEQ
F4lR2abgoMdjqT7yjYMt1oddxHGb9qlX2r86TEe1LihXQYjybmzFk0OGZauy
6RsZS4E8frERZppkLBzHFC9ik8QFmTeD0eFIrWfnU+PM+e/H94sHOhsqshWz
kDX8rEVn2Gk3u0yuktZo3cVd2Y5OepIWoGPl7w6wUyNZF8pv/088TAkjiL7X
AC+/hZxpFkjzxnvtDtxYgsjHBRfYJP92ormCCF8TnaN+hyO46QXCUUwh81U4
kFt1ffBgk60PGHnNhaIMcRv/Q2zVCTUN9w6ojx2IGS3gc8fiWhsrlZbKCk/o
/5/9V4o4hDcQHgk+aKDJ0KZtHZYg+q91pd4XGPDZeeWbDwnfvUHrJipZavE4
HE9Wob0O8F0Iuet4iAw4Rl6XRHVaLUSPRFNYCMCLtsqVqWVPCabllFU3F2zi
DQeDMvbyh5i8bb09Jb2g+2RXXJWGkxalxxevtq9HgP0CsJZCPzpbhAFWM7sl
rq4v6+lNk4cihHRfRkakEXvhaLhb4IBGSP2kg6aNu+BlGh3e4i52lIUED1bG
M3xQ9hmc4DvUE/pW93bzMNMt14+2NnHhFAfShuAWvt7y6umInyOR5zm+uZk8
eXz4z/JOkqPJYxF6c9bo4631SlGEas9Hqbv9wt1WhKimmwstc7UA+7Lxnmfl
Yb4ciXTOMCmxOyuIMXKJRo02C1LlFw2YnRRgAwKAuQ9I0DiJA2JWt7+tav+l
NY50R/LCjClGngeIA2EGMDsds5AhzeI5ojKvi0Phe+sTKW+6reypIfdFBYTF
thEQMkSkqUCKDwAQuZSA1PcXEZthlg151ANNFPj1Qo4ef+NSTn191cN3mUnf
pPPg6SQUCXZ+YvlMF52e2t5i/WRAbu4kR7maCWPuWmxY/EPEc4u2b2u/hb5A
OB8ZySprnS6tQO2/sjF6paViNp52lZKfTjXc9mKUaCsNu7Nmze2TdN+FCmMx
TCwiEwtSnasNKvhN1PZenPANV150ORJmCycKBk9t3TIuHVk8R5ODZIjWmiKM
LBq+ZsT3WNOm4/tghBqbClkyMex3EbTqIsi2bDFL1Zbg3pLL+S/yYErmLuRk
fLBZUrMEQbvej66BM+wcKxtv+34R0JOyuadeZuHt+QOC3//0yMNdvPLi+MvQ
GemkIqtfbjSoAnXeAR9WVPSBpL2EtrwQ/D9ITKODG6ih9iio3seuuL89lnH4
4vfHfFr0jW/egtjXoESK248sEzGdvKc77tNGT5yK9A9lp6deIJXp4Ji94vjQ
KGGK/q3L4ZYMQ7vd8U5yZ//5jb8PYQxT7IvV5h45VQ882nPalqMTcfCj0wLJ
92IEpWoCf7MzyC3wrBwqLW6C6cZ9lnjl1KylfbfS5y9tginWvi19ybjgb6G0
2RmvBi61k55TkoeGca0j/0hLVvzoBD8qnbJLYfOfg8p9Y2nruzeBrePvATQ/
E6GA8j6cYawa+OYavr1gXKQ47b60Ng6LDT42xEbmdRS1oI9z7M86DXgpSLkg
17ENsErVQ2iahf4LLSs3cUbRrZ/8REQOcHC17SwLAmifj37QT0NfD/R8xB4T
UozifHxHkiuBl0nVxXpTfCJ33BZppMCpwV2MqgExByT5bih5kzGCDNbmlBDQ
aHB+ClrmhYBMUtvwFslJwAgEiM8/KLzO7n6qJnX0tBt9EQIO4XIFOn5mR1E/
GICij5kRtESHfbsICFYEYj2RVUdrM6oZevo98hSlfo7UbzqE8FaOkjkdiCQr
F1nY37kpyC6MmhgCuMqXxL7Ybwlz80DAYfa2SgvWU/XS+HRws8cQ38D1mSYA
adFasJ0Axg02dLm2cNfflcyyVXC9hy/3BFdsT7CvZPZPjDzwrc+dA+X32NYF
1QkPpWCShR7TbJXzZjt0JQ3MGw2gTf5v07v31Et9M+O135FRnhxWWTD4guTr
ASn632VlVOGPsIdeMB87tGHkwvjhL2QhYhFJh3qPT33xAJz2dR9G1gzWi3Gu
uLfO03B2nkrHDJGgCpLlWTydCQNd8TCjwtqqDEYSPMGy087Wx/8VE0F0D/YP
58Pg4LpK9ThtGt3bilXzwNllC632n2BiySMtRaZQ1NpMPl+Xh8TL2QiYL5Vj
wJPHNZxvU9vf0AHDGCLqdKnpmOgrvDEtU1JZqnwV/24VujQxZH8tcJE0U9Gy
QF5g0WkY5oR7Zjgp8FNiMXHFPKEKS1PMN6nRzd26q1gtIkq9/hFQQVYOenTG
TmEKAv6wvbZqHdaCTJHxm6PGUKrYGi2fqGD/AL3GgoMkeVuprqA0IBnQ5Gx6
44eaApt+F65pQwE4LPDQJ5dWfk1kz+a379bKNhEnXaAD+mbkAskK8pFmZV+a
3bOU04H+VAQmh0XLUW24/WeWICa5UPyXy0lftTeTh49G0ecktCDb5zrp0ZfC
+ylTBm7O2f9WoqWvl5ydozM1x1Gs0Zbp9oZC/LePwiMpH1zI3rQON8g6Cddr
3yvCR+YwKYdQJo/9tYwPZF6Laby084SIV/UN0z1GLQdoPEnBx6sRduVAaFsg
qki8f6KbSiHDa9IpmY5/2YBbF7+L7ZxGSQXJZwIYmaCpho7VcrrXsee3xICF
iFhz79x9J40BHtNcn1pyqLImkp+ksSBHleNbhia3tLc0GEC2dy9T3QA4EbRA
eg/orKfAcTklL8ii74refkG5puA7O8AeVs4DJR0c1kovyLJd8sKFJmzlc9s/
S0jOeGRrG0OxZC59CNqBv0DzZgamfip1F+MY7VAC+wUz2iUlsShN36lkIzHD
KnsfUXIMcknXnpucSSKk6yT6uUUD47eDIAJyvuOAw/AK3JGxsvX1QRk1DKeM
PhifmzGBOdpYbJIS7LcKed8YsdsfwZiXimi8IoUtDzmoDso54fOsbmHo/TcR
x+xRIykTPycknfKcGmJE/D6O7MV5Le+gAJy8ceRU1cnY7+rumJW8nZ7rIR8r
KX4laBPhcSjL0hBeTM5sK/pIJdRuXAS5tEhGCvRvabvyjMIlefWeQe1cCBQl
MhvYpHUg+xhtmVbUIIud6zT/iEMd0uidJ+K/pV7CxvdQi8k22JXG/sl6mqFy
Nu3GYo5DTvJQ/NmL2h9yXP1yaYo9Ejx3A4M/JQwd7NBhqPmkdOLyCb8EURXB
nM0GJ2yCLGGWEDT4H3F9RVvu+G5TUQ9Emn5ywMQqO+7MrPO2wXRlnU9g0lBc
oDiGC9JQEzu/+c0z5eRRNmWUKXwuaHl24sCojOJWjBpNsChZF3E1niP9+xgb
qWRwxW9xcxKKN5k30Hhb0nvrgfaMK+vrrG3LCRLcE3OR96rAM0jMT0iieklw
aBsF5QKDXyjp9B+ey4AkYXugka+KYtMeumiKgA4e4HIeWxa5hnZvpG5KB98m
EIJJy+APcxJ2M+J0IY41jz6BYayyhdo45AJ1veF4oG0kFDmaChkgivIVwvTc
c0fwCZQF+P5S95Rjztz0z0UFH2Uvz8Lo/ByenDEaL+K8XDWk5PPGY8/C27GR
iHi7eg+DCr2TV3BuUe+7q0G+cEm1pziYhJlGXiRfGyoxtpd4VeDBb4mmNU9t
y4SFNTBRG+gIgkJLYWBpThsr/0wjciP6KD8DgWjRxnY2HCPiF7TcUNoOLYw5
xoKOJUdS+0tbXT1rktt59FpxiTuFOrlPV4m+ZDxIaqTWuXw63O/DBq0aF2Qv
XIeufB6F9RVF0Z0RcV1ZHoCE9Bnf35imhHeVvUqmphGOmalEEYLXM9tifGbt
CLclTaqEDarrb3Tk+V2lRZwX57sHz5GIA48H90LSLrjmMouWXJfD4Ml/aojW
BJwEp3gdcRqFgZ6V0Nf0eG2hNWw0/sp+5IxqfRlIacMf6midt8Cc7UPF+2AD
hphkgxYMi7GyrnjNWQVPYdo/nCfPThsDLHOYR4RFvuGpXzqGB1CEuN9SOqWf
cnXpbiP4khmWqkIqdNfqd+GbzWS8Oibl3OtGG1rAvttPpw+X+ZIVayqjMtvb
F19pJYlCDQ2gVxbvdrsLtvUOtfFBGBQW0A1InJlDfA1FR/PMysvCtJkNZ4IA
sG/Uv/1cBYJYp7gGLB4MSMKwgpwOOaAV2aWCOBPWT1s+6i/13QimjQCR1gY9
2yVwYCJoMOdgT5iKEU2SaN/vENf8tS7SwDpFi69MlM6/bbdJNZxnoQl2w9XU
nXV9LjpOrI5WMLjGT8N2uOD1EvJj60zU80OjD6kZhD8GwWlIuY521YJxUnr8
gnqR6aUHOwBhwuwNRspgO0kJPGa9i7uRaaVm6aP4XqNhahW4Eg3FPevZX/sV
+6gMzYNC0Lv35BLL5paqm6fNoe2VdAZkPItHkfN/4bKMv5Cr+qN+qpaQVjQJ
q6EnSV4RLJ4s0mjnFH+Hz3nzlbuYu46MSxPK0aze+6/QJPgWmMFeki7LoJl9
uLu9o8g+d5KVvnH8Kzri9OYJf1YaxaYwsTPc4VNK5F5eSt6VZzX5iofxYN2y
W4awWvngYX/FFk7dLkcpDZ5BSvZ7iLqJXlvK+qm05KUoeaaIG+tt3rEtty3R
SONtXnTe7kdeWqvRdpEhmwJ5sYWA7gC8H9P4fgcBIXb1W6H/cihtkTJfmzhR
uJFm51J9QvlUUOunb2HnFK1r7OI/Qq/VBdhQqeUCgcFJciwEpR/70ZUU+Q7z
l59xS7dEHdjHa5CTxbv8f/x2vptxCwb+Fp2Mu5yc/lNRKWLj+6S9PnBVThiy
bK+yQpZOBwU9tDDs7FwQyHXZotot8kVOtIk6ySjgCD1IUpyrFrk6CqG21wKG
/qHk/5dvt97aBmxfnUalR+8kTzWNJf17h6l9VTQPiQ4Cach9aFTEpNWPLghQ
O99odX6YpKbFYOnlvsbbBAOnJSkVbaWrkuVzAcnahPtchmmtO3MUCo4XTMg4
cbauwlFqpEM4O+H+cvBHS6s19hd6Rf6y7Mkg+y9g7rWmidSXQl3PKiHkG/I+
h/SzdOpS47w1I/Ly8b5IFjrKNFQiQ0zwpy5VzbBrvzm8ztrBIfBk9OMUR+Yn
PpzqhL3sHsSItDQN6SAnwwufnqMT1MLpZAqnjXoJI8+Nl4p7NGOW33D0cMJL
/rwNg1Rf0py2mGD3aSYT55rudJ54sy6V5pj0hkhRQuH4BN2jw9tXglpbxm/z
i1SYZq/1coL6/INZb49lF0tzvFylju0xIqdg4cyAiCKhJd1dQlw/fhwvFaz8
g1HkKRkb+psuKnBWqVRtFo/tOL39q44KYryJJpp0s80N1iHIZlQD1KBU5u0q
CUWm2xKrESPLCjxjob8JDeRevkGe7kFBNyzW687rlbw63KVt2XlUaUJTJAV4
nrPuJ+yK16XkCv+kBq1U+ewbgLXTuBLuw4gpAoY88GkdeuIJi5SPp2MlROhH
dB/wOk+joko0B6qgXfF1s6yhvW5OlMoPgXjeRtUQSQhKQr1y841wWuOpRntf
nE/86ze33UxjkpNLWLczG7mwksHtaR2DxPMSMeg3sEZ2MCjNA4ntkZtvM6pA
xv3woMbA4T4sLGuKBH7s7rop3iFfEvg8zOoE3kgjzVkm1ncBkxWkEiRiSuTZ
ZXA4pXQIkkM+HiOJuVqKivqA8QebxLr8IAKqHt0Obil1bvB3RKuUZjCzhsp0
8y67T0uJDsGgKKNtWrhNQXxpeLmjXhI59CMaBRg+0h4j3ZNMPNCgVz9eDx3Y
4Eg8yPM2lvoUCnKAzj7u/E1cjZvSPuCoI1I3H5Dx2F6WbuWKt99LPJCtxcHx
bHm3hSuizLzxoBVF94NMk4k8a1FWCyru86C4yQ0rH9Ai8X4ynD5B9PqGg/QT
NGHCWS9+KkMOvXkISpPrS2S2fy/pXvHxEPBpytUjdNduijgq81IXYJyKn+lL
/9J4dzPxowmfPLBnvd4f8gsXbXErNjFDUpDb5jk7UnJVrQQMR/dvWLFEeeE8
p+hw1FLgIVrR8bqqiV3N5i7gAt0q5KUcpaPUCQZXK0N9Js7UwOaZFDWwrDPe
klwjoYOp1mcnhrtB4MHkLG7xiU9QwziqLmxZzRnvPs917MmXxZ/TCKi6REDi
y/PrjXumBN/AnYR3XmhxZGRUmjbJosSOUymcKwwj+yBzgUksIAH3Dh6WUNby
e2AFlPOAMp+JQaZou8dCjnm/mr7+yMZxb1oN5Z+tHuOtfPb1d/Nmp+h3NIv8
7/FRfMTvgFJWNvdyTMynsxWz8XFGmM2eN+Ec9WaalEJzvDXRP2w2MlDOu7yV
Efw1p2cWL8bW/zKHCOYz5Qv2+r6x8kQsCNe7dtnqSY6SDfcIYzmp1RCw2Ek7
N10i6q7yNmUONR6+MCCoJUwQFkq4JpnOo0afnYbpALcRn9rFM9CJB22HAF6r
VfcQKJ+nUwIUEgVvpLbkXRhkjaVEmW65k0OqqHe0hxwMBWxyH6S5tsXd4Bth
sYrT5IrzCSCICy+PCssdcSNrnWKeCWcjEy1+7KNPLPINcwR/5cNSgha9WM65
hej3VPknYfWAU+XaYIuELvnTcpuhyYnaj3sJQH+XyekhmNn8x/UD8w1mKwsI
F39SFEe0+xQi/gElMgYI9ceFw2+FBYpM7YKwr2xdmdBFMJRNfHx+8RW07owY
n1WAD+jPUNpTGxuOMbzk7NZlC5mA6BHJjjNTXfmy7/9DUkU5tAP5QMkTS0f+
xFJ79Co6cBmZwINjYsd4u8dUTw8BZ19ULHq1FVJAI94aeQN4mXs/tcu5xKxJ
TzSDz7mGmCJQh8Cvcgt1ulrzyjdQA9maOcGVRfYhqnF4O+eDpGOHJB+mMaVg
no+pg/jN0JEt/BrpTNIkhXgVqz2njxfZlRVrz/G7qdGDQt/egfoQ/Uk31DET
xqSbM2CK+m0CLjsQElwnffAbjz2IoH/9dUyu6wF1WOeYG/fjmyMWLx/v1bll
uefkt+86mWE2zgZdxKCE+6ve9od7K+QfvnqTlqqhr0waL6S7T4CUe/tMWS8y
idfZN9q8qtnCgu29eT8kiG3ZhTpsUM969m64aiYL8fQSXDEML/4GyUNW3OBb
bLQNLXfmbkEWXJCgY/+zKccUWW+kUOMMQPND6U3r77NCmfe61oC0yz0SU0Kz
v5jV0msH/onv1M7OwnwjWSp6Wnp0ntAkgoF8/VyxLV4ViF8WkKgwlIWdn04H
LpTZthxuZM11Bgf8ylI5DqH0m4i9o+W56t+ssy2bAeb9/PVNS/nTZoLkaYZn
uiKwHlzNwFjbrFHEZ5oAHu/ly0+Krk/3uzxn8jtbjLrWxisx8iKcdvBqpe67
scrEgkaQVTRT59gC5V9AX7VqJEuVy3bg5Yy4vWW9WU/gGSqizykhwub5O3DT
XDns5bJvX0QL2aQb+K37pzfq342OgojPp5COCwzK9WVOukeHu/e9mCIHLHls
GOj81SE+z3fNgH2YVO/CbYY3KwLpRyxGWV60WrlueURmMznM/OIPRb2aZbsT
XUuYueqS9goXu0d5tQiZORg8hh1qLoKmT6spycWbuoXJze8HYVGvrZkRbseu
MhLB57+CDCasi86nEw+RPGKyoT/v08km2gpYc2CLoghZwSk3BVXToaLxbZ18
4P+ZmZPyIqn3+YJeWhMQg2HhCJhsUYBmu/VIZF+ShGCM6PCiPOzyazRBuFrP
TH/KsaAroKRIymGh4KBv/YIU20eWXPaIqyZSVd+5fKA1fKB/Zee45iZkNznt
fqcEOfcSIqpCGUSLyXxGYsnSdB8MeJb2KItBxCeoQzS3FesUuwUzt6/QkV6h
BxlQ/NRtNhmFLjl14Q3X2MUJVY5KxYjwWj5vbPoC7LstGRkfWEg1OI3alGw+
CRA2dwPOtBcKzT1sw6eHvIkMG8YIsHyFYaNsgg368Wtd630U8jPczE3o2mjg
fIxCIBOsJMWrahifRcQzckEB51ZXNE/EtAFg7gxPkSxg7aBVQQRUHyes1Y1K
9kDWC/XXnyRISBuUbJ7F4TER3+bWm6HkCj3ix2q4zmLfgx7pRkAF86lQPs9V
4gG7thP1/As1U3Y2yUhEXTSlG6aN8EtYu4XxLJi6cA7Ghi6xfBicmsFWP5H2
Bm4PgvUExQ5ZTO/RSyQDE317ikG5WGKUECrdJzCVqcj0gpM8ZL2CZxz4msQW
kvX95i3/ppTM02t3vN8LBl4HPA92qQx4TIxnbog3Uv/EDtEB6mRyE3EQMY3x
mtoyNLbjA2RnOnrTmgAbvJye7u2Lx3A5RNr6XiC0hQj0MEhKMUjJ7o/6J37f
a52/bdcA31vgib3l+KjnEqn7f79r/7W1z0/92Ufkka0fZ0JIZStpJq1xpQGa
xJGA4LFJ8exW/syjNmttVKz3jcswneilC/DPM9DsSx8gcZAswHqcL7ZGZCb9
HkV5eVIwYnxOYWPQWs2tiDPtr7viz99pRcD99aALW9baLlA2DCgJI3YvgFvP
D+GUn1i3NO2VTNWwYpVD8TNLfTjko5fc0jMD2D7KU0CoFZdqip/8Rgh6yOAi
btdQRuTYIXpbHJPp1qmSoo1ZODVLmyfLb+N9xhSe7DodNa2KjtKm9otWIjJr
DlXOkJijGyNWEtJ1CMFU2que4/kTnSRSAap26OZueEcSkfJ8yQ41Vff9Hp+m
RXUW/H5OEt6zNSwnbhOt4aHCCgNAu/MdrljvXO6KiM7BgiQImUkhk6N43OjV
8hPX+SSQ3FWeXSu5Icg27gPoBFLqfl0j/WHzWja1Fa5VlnZsXGz9WjnISqR7
ae2KaZBwkrtlKPv6QMGvZ8/RZthU1E/naXtpZ8PEputZKrFIL2EEAm3rJHeD
yOQLMT5R2nW8Mr6cFhpe3Apu6lgWLMzAiegB8D2Xyx5wsR+u6UpI/FtPExlA
+N0YOwYLfZJbzzwdnMSfoK/zNjRX8t/ncDpLwiFT8FWtucLQrAgkuhcIjXPg
tkGN183U01gm5Ki/45s4hCF0YBwGHpuFMD8S7dVM1aFOgv3vpZkNbHJupxtV
NlSplAOsfsHtg6LhBcHFmog8Lhr1Wgk4LqieOF3rq3VUINdrd8qkNiatgnza
eP8uRbkAq+7hcjyHAUrsuAYVU0e2BYugPK8s0K7acrDJKkblTy+W/w8FiHkd
8XGmrncZ5BewYqj+J8xItJA4SGQLqPwa5Wm1wdLh7Jq0NIgGmHlcK4kCopUc
ZytXozH6BCpRlPPiiyye0LtJf3+oVZ/KXv16fjPpG5PZxrGh4PAyl2aVPMKX
GWIfIsP45qvtdeyrChcZeUj5rQC8gE8TT9jBfAvCdJzo/9p8xYbdJt3/Rti0
744kgFTM2NwVYcWJya8aC3YOP3GBsRuTLUnwY/rtCwN8kOGKoi1XN3LG+RPb
3GQbxBCIHDKXarzCDXi1LyV8GxtGopMIU4tIafmEjS99Z75hm/7z8SWwfTRW
NdagwoUuMWlipGQclDU3KuMaffeTXoQvziCykh4MFzlxBezSb4mFGxeiT49h
wO45/2uNy3T9tK4WzqqfwL3p66gLw2KOcPtJobKP6W/vKmNmQ+Epc5q8Lp4g
FiEwikQhflOLhk2vCfTRzxgPo9rbgZS3SOofOHtahIlyKwShdb8cWyG8AZes
Xm4exaQpP43A/PWRVV4MnpC04L0L02hsKPqtpoP+xR7Iv99j4gLExwi6KRLg
c5gtAHTwTOCkIBgV6HL2Wa1yOc2kKgd7QCK9V8XCGJ3QLFLjSMETdJYvizyO
vpABpLHm23o+G+hFNq7CUmWi1dLf35yDaJAUy++8CsoaY34ka29xTHJNa6BM
Std3/CrHOqCW5lMJEXBHcNcDeY0XgoG0ERO7Kq+czZdRAomCK+Qq0HpGC4eR
8PXtsbGgSKlVFCFKHxTRcbv0BMxzqe1KAXcZKQo88EPIwE4yFrRqDTsULQnM
YZkU8eflh4vgDuvRnFK+/CRVwCFMr+9XH1IZg7LnStBbqiQlCS4SDVJ91hKK
EyetnqUTjL8Q1HMugILm6IyQbUHgse4xmhqyY3nSwciuERqdJDkuVZp04Whv
2pxaNVleiXJWQ4Jix7Hp97IHQuu6zY0W1P/bwipFOSijTPTx0tvkKES2YQxM
ml598temEPracyb9L3s=

`pragma protect end_protected
