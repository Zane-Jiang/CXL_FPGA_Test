// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
fQV8OJHBk7tT2ha/DoFM60GgQ4AmxEguHhw0bYhCqlBMuuyZ4Hc8RIb/AKWzKcrH
naSXFxRzBUy+HhXKGTSXzgI6oB3cRhrCokv8Cdr8x42lDsnMvmFIrkKYTET8/tjL
TNbe/KqODJnCpMhItRowJMgDMTssGHXEPfZzBZg9pG8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9680 )
`pragma protect data_block
CQYtjdnk0RkS5WU1iI2mDTyzXlVYLDMJgYDUoZAcYwetvg5lasY54/3Oofv70HyD
lOHV56b9sip5ZZXDiveWYZn9513qFiw5Hr98u5cY87OhihQjqsP1Uekdr5njv+z8
hUMOYBcFjf3tIvVtWgCE46jJD10B705CljHhzV+SPSAQSOiE0ADVnWZLNtbaLLtD
Kqre4untsuMbwk4HzWzW7HZ1E5V40NuMoK67nl3562BecQPv7gs9k13yeTVoHivu
ukAijIXpNkXqm4FW+ZMkSGgg4Hu8fcZmCvUuw2mMqkj6J4DO9IJXJVY6t7ViJlD7
oI0/mjX8rcinbAUSWYA/2YXEoy8QYllUsqrMjvH51JpsjjmZIxe9upVuQwCrMWPo
45zY3+4E5ElUDVAnCVqJiF//yq5+yFsejlOr2u9YeSv2Lt6BIKjmsgywvPDcf/Cn
EMEi3rlFeDhjRWUCcn0Vu8zBxYW2+TD/sczXmzcLATzFBrybVBjDg6gLOrLRYNtF
gkVbdzLQXwuiCpEYuFZ4kyoYpFnq0+lLkVy8HiZJd0JxnnlDnMXHgW1pukDYdHAP
PJjy9jHhDnj3q/4xonaOrwUgLlnpdPaHvj6G9XjsjMxy53NPDxK+JUhf1BKklvaG
SXaCxx8w1IdpRm9P9bQL5c2WGDvsWNH9r1tekQojd3kXCofP6f0PmUKPxrHCzNNY
d2pcP9ncogEdDoNARwGhZDJeyreXpIDKlLzikf342pPboEYHgeeZ9Hn7SUZJo4JI
GboV3bxdLquTADAnbLEMwgA7m5jYSvjqmNMGMCCzTM4iuGupPx9A4pH7vH3P0naN
LmiqZMW2WGicqRUEhz1z3F2wnatdxBPmfugm1hzJPQiMqoaUh2XZTJEGY0IgKymw
911IQ8mkSMuqNnQi5GhE1nAIYx156amlw3yuPVTj2zoa1W8qVGDgOX5KfhOJ+YFl
oyyPp3dFzTw+DWLFjA8OW55nOXGN1SxMbS8RK8oQc6cGHQlTAtasuwPAP6kEnYrF
WRrK8pCwlHQUKjvDRtjgCNS5YlWzmfW5ALa6YjO0idj4GjaiYXV+BGUnXvHs+T/A
Itptjt9Po84U2WIEBHquG8n+zbNIisIXXu7zjc3TPIOnOn8an3sbNpMhJGcr4oZb
jBkwOHp8Z6oYwUMjCry/BLS3hh77LyNjHytcnS/i486W78+qM07DS2ciAIvB+VCn
xJ1LbCIo/rz09QMvg2SRgWur/VGxMytSaylfcTP3UOAcFJQJKHFupc9X+6nj8gVw
Ka5Nq8WsDu1Q9iz5vKcCqVz/kLVyOao8k171+ITfWVtw72D/V98V6UkgCTX5QAP9
FKrYxwFVnqS2tJ8pwKGrE8B22aStmdi7aONPy4y3NexJ1tz/uoxOYg26FUnNutvI
5cjj3/NkHmWq1eDb1XBX8dzF57/47iPW0Rj4fTKy/x7AoZ9VF0bOXab6I2e5uuot
3yxzcPgNpXfL+ZHctOKwi0w6ZmUjff2CA9vSaR229Lwgw52g31pV/iWzq0PGZDP1
us20YsT5P3JbytqKgzU7+LI98Bj5vdE8pC8vUu8Nj4WZuwYzQPw/eVWA11Wv4xiq
4bx/t9mvblzyXS5GWYEotJuidJEeGyeTp9V/gxThI2qyR6LR7A51oPcnTXwKtlI8
w7vlwQNuYUN9SCJ7YP9+0eBHW4v4w47lIrtpu7TUZAc5W/fnTXl8ZfOkHlmITzpj
VDdb3+jFjgVZvm4KM3ko/IpVygL/OGu4m06W2xRHNLX1GFCZJdHOeX3g7nOrYKGd
q5LGfRRRyzgFQYBq3E8/8NGufAzCGLFPkdPmxCXtWP6RPaFbbpjb4d+M8OZQkkrA
mMCUrOo7iKx9PyEbg3OzbKA245pI3gAhNaED8RbvpEO7gykYsK+dpir1iLl1S7GG
zpYqYM26aLpC04F6NOKF+MftrrFU+PVrDOeLh0AjeAOae38Lvj0TbXQB5BsbvCsG
m8IbNTJ7UQ7gEJ/KtJPcb0ukFec4l5xytiu6ATKSj4u12UXUuUnHeYp+EQ268PS/
T5xfcuMf4ZRpFv6CQUC1QwsuTuYFFCuIyGCRmd/KxSYsj8fRJWjfqBhZCZnRUoQ4
WmEXQReKXQobo92gJhIiXSszOlcLkrflBEYgHBcIbSwtTiRE2ON8StL62eOctvqD
M9cyeXZFJ6l3U2AwzqIiT9I3Aks9R19Ejh3D2ymro0WzuCcnuVdR9VwL8YBKMhOw
PBdd8AXvdJGpG9YlVwl0AWFrjV6y0uEfxEZsqlGn+kUk/cDjziEptos86cx8XsES
JKC9xlvFzkSQhDR090ZqXemQVm4k91agdEe/C4HTtSIvGFWPH7aoYp/EsgfmPZ5w
3kPvX4+//4g9a8RQIasv6OXCCF0YpsWadqGZcC+vMTen5XMKkjAcTfTCQMtCWL3T
L+0fH/JOGgYse0Yv9nswLuRPFJS7r6tSEByOCgdLvLdYTbcSb6FUGfgZERlkX/TD
7pM9fP8xicRaYSMVr40J6F7hYxjp1LmmI5QyauyXPOmk2/vnlEMBCB45jEQuiPwf
qC9vKODvvauKOuY0vW9kL64X8Mb8Z632ir9ZzoG3V16Ry9v4rxmtg7IDfdv5oiFK
huv0CKsfj9gnMjwOFvsRw8g5Qr7k1cySbZyEg8E5dUnisZaT0BWwoDN4urSyV1bM
+3oo0X+KPfRYw3mW/qezg3CC4DU51Uqt0tFog1dtBcTegraWrzYOuP3QqS+i5AK2
VqxIC+d3gP3X0gEjwfkWLUu3HaldP2EaWMdZ8f/H5lhb8xdZ5FXHAaik0jDja/Io
qNGMLBFq0rcRzfSazYwIUSgy38nE0ziTYlL1pidacfYLvzu/cfN+EdoDzfi4U6El
I/epDrJxH9YwmrCDznLSnKmlUQpN54PzZ9WtBmloJw3ecAct8jMvDj/TFJbJxxTt
DrTT4ZwD3Zl/pArsI1xaEXDziG60L3QTgLJgJI0+5TGMxfYOzapnA5QX9tewzaST
9xzXcGxp0TnUsUNaLB/o1safxD8vHzO5ZlqdFa+COmy5wCJqO8qOL2lianDnf9pR
n1r+diRjJkS2jqZ980qurKD3SsZMCLZ3m9NDJspusZBSAbTv4+6IRErFgUFKQ1TB
QmSRn7DA6Qx4ZjQ6LMdQawXL0nEdATyW4DNCRS5wyolkGUO09MzH9/YsdFtfQTX4
ZnoF0RWtr5oga4aMScTi7KTf2J1p4gT8BX7wri+D0hdqeEETGUXBv+qLuaXZSozc
dUUSdfXJm1S1Bik4txrO5uAw91PTIOwAsu12pQBXckIqdXFNRpSvnnoqVO7GM02s
tfEP3mvRlJ9U4E7UGus5VXlKmhZyDUphzZxaCg363CcKVMSvC+ROZAcyV/wd3JPG
hcCVyaY3BhSYG1JQk7QcSYk3sAdnG7GTNztvp7j4ST1JPXGf5wllYGKoQppvJEe4
MmqXwHyzgGYLmqlSgx0E5C4BT12CN9qnvAHK9hLb1G9kvJRNefhc5Ys6YRB3QpSz
FPMBwlAMU59+pxYLDqMFRtG0F17ZBCDMpLw1YYcm6Ar1hv8tci/QIuAGvJ+jjCAJ
okEe+85d0FmWcUc7NSEzepsaVfcQqZqjZodQhG3G/dCeDml5FdQJ/BvJtGH3ZNh3
aHB39x7aZ07AvbxdiWSFC2CsTPIOMreSLm5Qwd0ueEmTd3FoKJz6Kz5E8myuJvC+
Qx4fXSbfs0T4BX03FrmIp/N0semMmSMuNTPdxQUqnIPNwityVX8nnjJcK3qzpMrZ
YuXccwbbmIqkx/kKm+Nm/Bfuc5iSCz9TGzh6VHpBcff3KXeG0s9b27/IiTmdoL9w
JtGxK4IX1CiQsAT0DuQDocDQEpDqIO863+D+luuuUrba4qyubQ7lhCunXXDGN8pL
UpYKx3g/nSD76Jeqae775XfbGv9bge7tg7ap/A2hDir/qGdNbKyM/Q7TW7r+nEOo
9ybc5NjYLT699FZdts1ibukn95rApyvaX9+5ekgSw6G76ztkd8YqYyczQYFF+w5P
iQ2/Ebal32XKWqfyP4q+LgW7MHQ5+4G/ef4ikLT5mDZd0N3TEIvTdXC2DQfktdSx
PowBrGXTjvAbv0/3widwCBcT/F1o4D/GNOMjLr432xzt8uz1DWX+ZuYA1hoVEl9E
Ep27YYPBM7vy13xYOLCzQJ47+5xPu0PaarbS9c21EaXjIiqDj4d3ChyCbgEYKFXQ
AYmEXIj8r7b4/urxGzwt6eUg1qeygNyAhvA2XjrEEnQmx4QTPGHjooiEkieB0C/g
pUBssxc7ScYK6PYv8TfBVTdHlSzFwEuzeTgZgmSCdM6VoVu2vzMa6dkROaK/HxSR
hSef6xt744SsnGUAmgvQ99PgehvSuvEoOjVm77g3U1Hi0Kn92ygn+UtY7BxtR47u
JV0YiSoLLgvEq2ksPxfYuASi+WhxrFC/Zavjt64W3RIVguFxeiCJ+Jl5pNqeINLv
/Rb0CrldS5YLodv7bp1if9WAiaZON1ls4aChzw5nFmlIbZ19qhVYRs7MorHSIEO5
PJi+PbL5VbKhhUzqkyl4acIhGTcOUSstNavBQ7N+JWwZXLp0avfpKfUsIgMhicW6
Q8ackbp2pp8GsRr2q8/HzZRgVvQI7BlkX71e4/ahdr+J6nyi25j2uaWznXprfNjn
gz7L8niZWou/vQ88zmeDMMz67SVULmCcHFJJlNDVWqfrxwfWnuUEF4qUZ+uGoOaT
6BIGi3FfbKH2Q7wzgYJsJXE7hTheOsIsj8WluaY1plYiYB6jHabiwlni2CQdgY1v
TsxbeeMwb/1/+UnIyHtOtCPiWcXNVlgRneLONsxDSyONXiTj+O8evbLb4sAcKavE
Sw3U4GnilFJkZnjbtdwwHoSbr5ZxYzGw/SiDj4/IlVYgH1XSckl2U4tv7cMWHCBY
Q0v7Zw+fI50tCOjlqHV9sma0XKeUM9csyL5j/gizDCMNIekBzgeVJHwoAAy6dn8l
90JjsrOLOsCQbZBeNHxI7CMvdunnXd2i/ETNJNwgE7+Zu8PKcNVugVaiBUVLZZHN
0rOx0bn14OnKqEsN9fpeXYy3m5MnFFxNdjAF2mSiSYg9NjQHBwl4pL6ptBENdvUl
RP9f0K66ytR3wRArLQ/37JOUFYrTZj6CeWVZmgSyFmuuNFsCUZv9IRr2SMdBtuNO
y2F83TDhy1Ct8tLd6aNX0MYryP2X8wnVPUmndC/IlFW0JvJggc4OP3m1bMaKx9m8
4eiElQqKbwvegaJppkhtvCvPLn/YOlHyQnVmArUCJXQRJx2z2ffKzu9gh1FZKlcB
pOglM2oi36uHBskuW28ZzCXkAfQm7Dk43qUl4/Fa0+aS0lucVfLhWsEI1tGFsyNC
jIiDmJXC22+whkWAHMzEum5cA5zSlZ/bdHLrLBIZpPvMMDaI17hSKUcpLLviD4jA
UMB4bbPtRetfYc0m693iRJYTaEnsuRk2OxwToUEgszJktyPtH/j7mA92wpVXaj5b
j8CBPuC3UN5nVGUSPOFt4qb7w54wUtcEzkkeceWLxdEnzViflDHzrt+fD2cBWxlF
7oMUDUDNjb+Yd80f17gxF+7kQS71tYby2wAsagN0ny4o4fhkbeeCdt4YWj2BkanW
zcIWQVpPTc/bSIOPip+DOROzHN7Y9y/UYAUjCbaTNkEWZA0+aitWHikx9XUmmPbG
2brZ0P4mAflzhHrGKB6rJl5l+Atqa6/im3vi8ZYwlG4Guyp7mHfFxj2PUkfDehgU
6WSBOQ0B9390Z+baubPW+IGQ9TSBiAYE58QbxO4fjTmE3MGdabMWHNjWhumH70+C
jCqvpHgrfA616PNUDz9bQYZxH3mSNI4nWo7475wo5HYWnoD6pELVx+VGhDYFsmjr
1Bx484mmPCwRF8DLhpxDExWcU5w9dy0mEFYhLY/aRfWmDbfIMiSzXYzy7uWcYt6h
ragZ4w3h82kzSVb4tFSbNrl/35sMuqAvwR2j/PuWDtM8q041WbJfQAp6IcgNL+ID
2SYVCk5+lDL0C1gCI2P62I4fKVKGVSWDgasiQu+J0NlfPGb3TvymnDpvvK47uGyu
uZkFrPEsuKRKqFUR4VvlVFuyUoCrKxRtq3bOfC8T3RDkL8ZLiyhM9iipUpjyMd1+
mkPp90iMTR+qBRTKWeVFuAvRhbOsl8LyGxpn0D7vky6ketc0jsDaEc5ksDs95Inz
19zGfgeoReb/4N/3hZHWHo7QL/nUqRpRRjxT+719U0sjVwdhYhHUTKHy+s4oPCyG
r3w24xw/e7KHjQnYXgMqFW/FeYEFU0hkoRTetm2gbU/LWgcHYYTNx1gt05wVruho
ItLNtRGbQQpZTTgCLOyj52ank93PXUl5hQUWa0xQiN/4QCS2jtuCdEk+/8r5dR4b
I5Tf836gP9z510OsEWiKkeDCwrbDLZK2cf5qrxlexMYwqXHjbwgLqKyAc6WwLbeP
oMl9NnqAvv0eSSSsjh76egdmE6Nlgh26lkiNzbVZAvAu0IdBHI83bmk3VEjkuyci
nm2jr6ofi27eM/65iqHr31fQwRlfdTbfgvAPaqhPpIU6+YTCIqU2/u8Y1MGBWFDO
u9R5b2ouPwOulMxkUhXD09oReppiQvWoVmiX+MCoOaCUk1zRKUBA6HMwp+fQupHt
Ce9CE1nBone/CMlk9XTidTJpR2jgRTRviNCjAtYPnyT1Db+6R8PHLdr+YRVb0C9y
RI+DlkxEhDPvKLTDyopvE8h60obZ/lELk69R70U5+ZG5cKQhvYAZTf29ugUdadE+
Xw3JWVTzum/2M/LYE0QqXk4fsg+wJQfv5HSZhOo7kov/oMzCjkhMT+Mq4bX40OmZ
l2YiyIx/9rZkAl8AjNd48jOQK9ahJFIWeNkLGnoc14UpOxwEaHC8I/62e5IGbBqi
FjiZVAhKM3jjw1vpz3sZDI/8wG2EL5W43/TF44ONlqH1L4c2o2CxFKYWsPGhb8xj
pzBaUWzyY0nVSsQY6HklN8uXpx4m8/AxcKMfk2yorfvasOxfgxGLPiKJTW7d++Kj
g/ZEsAVwBQryjGGQNTbbiPFm9oEeCDuFcWuPClHZI4K01d5UuH6YdeOKA6d+8phX
vresYyOBn5pCEv7UYz47IEdPC/jL606zjGGnsUO6bHUZkHm8wNAxM+LkIaoXiwT8
FEaGKtwmN0fdPH56sUbFWJR0suCvIp4dgO0CUj6ynvPp0JZccq8hYGWEUwHw/9HZ
UmiYr+OLOr2lxaauyCwkuamovkWPeDNYTzbs69tHcgEdftGJnFAc4fQLplIABulg
RJNRFh9zBfrQrb6jqLpIvEVLXoBXTJuOkVFY0FvWDM28lOawejky3I5q8LsSUk1R
CjIIzmf9y7IBCJzNtnM6oRouu/onmINvPF7ihb2+IwE1gwW3IZpkrinBl7bWTiQx
0+nBBq1+9DD40th4DInKeei8ALk2zq2fte2KlfeX5j8neZQ8vNm2Lxivzgd3Fxom
b5D0uN7/iCLBqdtm7pgvEqZ/yUjlRnX8D143VDv99uCWCSmfbSHnmKof33Is1n1q
Vw0krUNII9lJLH0ruGMpwMlbJC+ZiMSaXLc4NUuqyz+NCc4hoH7o28OhhuiP0RUj
LFME91wt3P4haLIa8I95piJvc1a8IYSDTDmMx3uv8a3lxNCIpOhVGUShjdI6KSP7
/3XdHq6xBhQ71/+dwLMWW/6I2y4ELEI/6cSaXyNAIioGzCOBLjq3tYkr+rx59t1A
eIjaKvbDQ1NzPArQuvYc2d+5Yty1puw8WTrEnBWo6TgWpNI//Eis7WGyv1b8HqIx
Un0GcVhPKNrWXIDFQ8xB/Yr/w7DtB6sa4Nj0wlm/AozuuuXWnHYF3OvJQu3rfdx7
4jdwFlcLDqPzxds8hHZAM1HrLEzBP0yNVnwH0d+OyEBomNWUWMVqRKk2jCVu/vV6
R4uxUtJ160k/qIvMcQUHhWssptiJZDWrt7v+cGGeLgqtwewSjhSS4ezYMb+lkzBh
MJtDG6tPYJVPCYuNSODex4OrffO3bNBBBlTwcqjISpO6jla4xTnlVwtz9clLIx57
/Rr+5m5Qlu2CxHWJVZR/s32sYDvkNgAgCc23XMyQ38bK0unpDe9EQgo4DQc5iCm7
Kl/TAxR0eqCkr+c9D9f3w1gqMFVSv+aRNjMZ6rco3kEtCbe6GoM3UaxKZyjijt+v
uU4e2AP8Myr0pvxEJ1TYqjWXZkA3HYKX1Rr2Je6cqvPmZw1xdYXicL4UHXbSZjqK
yXBQRHsh4y5HdvqIcOVw/YESf+vVv9VMYOw7xHxDaeb85ob2a3G9/odj25moxVS+
YoHCxR6HHP+E+7tLNtRrYNMEsxdgtJsTCL66xprBmSIu4A0SjLeZV4nOx2cBmwhS
9annBK+RZUPjQr1FiO5tlNsWl1mQ7VikwsnIdzIRVF8PG3DHtqEsn7IjtSTxI6St
nYg+VK9SG5wRiPd75XzcFPvaX8DkkCW3s/+mpfD0PCaeC3tHfZWb6RRbzmLUEALk
GttmJVmCWZl5wNw2yacWE/oS0vJNiCygEtPTof80/NnIIkZuZXAqfoiqHqE52zYB
KAlr4cB1yHbdIoyUyiJz3GHSiyDNGaS+jakUQH3XvyGu5qC6K/kAAS97MKLCg3Vy
vlQWzI/HnSulq1Du835Ipbq76lfgtWB3MkcZL7cZL+7AuRciTF1cb8TsO2982c9I
WpdKYZ92WbORKtPTr207/xZXt6tyThbEYzZ5u6Ym3/m8bVG6ymz1dLKBU+r/VOtC
D9wf4/jVHzWiRHQtmI2xBhYwHAcHbKgzL4OCzal/bUkxMKV4zurVrTGvBQ+B9Zyp
9wdzAGRG3meO59hGvWS3F09lJqEicmur7h4JAoiZvMprM9Ddf07YwYuDk0Cw2c89
ME4hl0LHvvvLEdBEzncWCDorZ9T+aZRom5UjVYWXQ+ujQ7JmQKN5i+q18wlbADAz
DoQP4fkyhOFUBAU/uLc9o1oPtB4OolFafovrjFtJSoK5u4f5oUZjSXC8Hr50XiFa
Sum7Hzke9Tbm51XUFeuliZD/fN3VfkyB9xrILPF8/0wFl+BZC8jwFnG5mTvAqbd7
GP/MxKU+5c2zd8XDHzpNAMDE5/0988z4+4CZdo3FSQ8XvyESreAq0KHkzatIurhU
Gt4hu2oOPyoJDrX+qrAV2g6DE0QQ3OkWb6xX7ADlf/dssbmiYq6coefEjvOjFDA+
WIO6Gl6NEUrAlK++Vc5HpFnOMPFbI77bVRMJD/yslGeyenBQbIBd0wDB8hd2BkOr
gypAHSwuAw6Wrm//6anc3nW7IEC4OGRXC3ms52HDdPQHDvAzMSC220JCQGh8MuQN
xA9aRDDxSx4pzYmednaE3K22U8mFpBZqbbmLaUE9MeO52Fs2N1m000D7SSZxVVeE
9BBjILO6WRmVcL2FMwaM2ESJDbcHZUKC99hZGvvheNrlFh7+pIhaPuC1rtqnA+RO
j8wFByeboAOpifKlLBLdq1yCVyKmLy+6P6I7OYauTHgdov1sbsIICU521Vyesptz
CIF5CCvKUxeoiPaanjSSVzyjvIusBITBMbwGMXzTUZjfprh47BCA7HmtPKQ/6bkW
CZWNMYRyQjmXBMC1az6TTgFf5G1+pxI+jmoU4IRarKpkfCVXVirpvkyyXd8NHuPg
sz7X3gJoLQWWYi+8KRJmEAAbu81QNfW6KMhPUcIONND+B3YLN0nIlo5ye3Tx8Maw
NGyC3tSR9BYxGNkV7qd42AhXnl2lm4u5/A7ST7udz6REJX9/h8RHHSBSOCrU6VFA
R2Uj73iTsdQEctBPWu30Rya4mgBDSK9IehcTskMfBiSDh3RLzS3GjQKLo/RQKKqj
+1x2qhB3IKkpGXaqk7ljet4tRqz1YaaEwnwteu8gJRAlzCmOVFZBN7tkusYa4WKW
k69v2NNfZLTWBDpXY21qNSFqYdEM6z8gmDzIO2g7PC6C3/I0eNHh3QXbSOcuLjhr
J3/vIDgCaxgot/HToXY3eLwWapq4uh22dtexPfz5zQEeHw7tkskEJcqImd6LRtaf
YEC0b13B3s2afIv8iprAr4hq/A4K/GQAQjfFQGLqrN+Osr1MkQI9HO/OuC9oXkrJ
coIY4Lxm73+zMAdgzs8BEfQlFmEJzXq4xCHoa1zkQlvXCbHqAUHXZdqtSnR32aKT
VoXlsd4za/YL7N9UTT1LvHpHVDUzZYWyg9IdbifzLQac2EGg+ga4sfMVs7MdbaLM
0YsPCULWpGndc4vBIZdBvkm7lAIvkaAA3Ovex0+OOHz1HPhSBLiBFIROod0nQauO
hKiMGSIEx+e9/jRLNKfEhMCh6HpsunJEfLIor7O2yjEfRsFC0JP3RsvZMSjjCob9
yq2kcvO5JYNDqTeeHq7xJDpNFRumA070X9JI+sunbM+fyARr2XWYBLZgOeHnbOBG
FvZfJVzB1EiOf273mR8Ib1OuBuebLLxLcmuivjHvuy9OsO5LZY0APhqk9Pa10+6k
BTBV9qD+6EGQUDG/8NlXSSXUc5oQKj5RQO9jnfxIAjJzWu2Jl4WtvObk0Mt4G+2e
MyBLkPcboVxI0kQMbbCVtsHT7kVSirnhjGh229OltMzjwS7qSwGPrjQgCWesv6eF
inzj02hbbEDoYas9H9EEgJ+NSwEf9J2v5fBcxfZ0+tVKtmRFaQShT/6mIvEST6c1
exANdQsyoK2gut+FALyzmJP8bJYw8xhuFZVhJwkQQ9eCDbTFMXhjt6wF+HvJmUen
vlrfuA3lI3MA8jJU3TMrvrQFC4BW7sptnujbiBCz1OlbyE7lCGle02CrxX+aBqjX
jtL2j7R3H37IlOhaZ2+hbBO6Wq7VuCOuAM0Rk59N0Klh++cClcffL9ChF5J6buA8
RBR/PF2atvbB06pipBWChSfPEXbkV+g56mUFO9tDXCSzsJfgj6PwJRDlHx9VZxFB
WAVVC0RgdgPLYkSGMj2GvT6m3u+KeWssmEXr+qrkPmDS7Ogj9IDeg6kZrk8TeeML
fKLCEb9KORHKkApt1tL8sBOtIcwe6Y/TElxE9b3Rx+RMTCnsYZWP3LLEJ8XdeNCR
JEkqrpHaaaQ4cmpphivvrbb/CHmwr1UMLyMCzPvtAl2S4bwOoUrQYlIKLf1mWlk5
yuONEwD8wj23A5714aISyhlj49l4gQrS4YBd52g59hsvRv1Fwnnf2f735xWOUzJh
uGzteSHs8spn+D3duaufKfgexjRqNTGZ5x1o6gurVz7AAVsV+/duykZQsKIZwKr9
zo1kRJ6pqhCJ+aNyiEMXJ5cttH+H/yoFp+mVY7xFYhAVIbYg3P4AwhX6nX4hgGHp
JGNCMvIckQefPz6q9BtXb4mV4mPv35rPD364u7Gh8e4VOXsJA/b5E0yNmKL7Tx90
wo1DYR0sxhLsCBhCt7UQ5hADJmwV4jCm+b3GbJTZDTdwHlkKCnck9lEAzdP7gdXz
TgXv961x8euVAQ0HiqtDqfM+wOo+uDpLKhqsvuadmlE0JC4lQKGOB63X/i2AI+yW
X9/GpNvXgXdPDtFWYV30GMWrG44sBRsJqOq7iir6w7ekMHAz59izGnxw0hX0gSl7
NPuC2Davj9ohaUi6AqzKH7JXHxvIgS1jM/G+7+lrowMGyaf4swN4pimRn35LlTLg
9z2HEmtD5oqk0A4uPT7vgQ39sPr6+ph1d0G30RrRkG1ZosKBz7yNd8eR2GX6OTrN
1jD7YXA3NUHdJqlZqb1A3NCMQ6UzCF1gS2ARGDTcUuIX7YcqgktqPNaEGRpl2OIH
qsUa98CwV5umZ17pHFOkMkRIIMLZCe4Tr1X63RJodUhQKjSasRx10wq2fPF2Gmka
/4PqFFGegOvE7VTniLN6alhJCGADqCbtlx/ExA1MAeUF/aKU7ZwEshD9nUEduc/e
5iIsFRF5280J7y27xuriTbMlOlaXbEV2KFWhV41XZCwHTM1yUz21hSyQ57hKu+/7
kCc6jehK13+M0VmXXANBaeM5Tn0zFJ22QF8d97IMwQt/xZFmfMsvpSQjJCA8jdRy
LcqrydUzZd6+Y8LEaHTJ2zHWExEe5hAgq+ytTRQAJZ0AJnZUaFFJ7YZK5h6wIPr+
nz1Uw2ZMgevpMI1abIsDzfeU1ei3mTT+sx+UyXS0Dm7aopSAs8+FvLdjq1mPg3rP
5hiVAq2F02VffN69QgnCmc15/HRKdb+SQFyxhnx7naE2LGeMr8IhhIuOjmT43mO/
u90+d7/fo0cRKeSQQWbgLeuCUL1AJTLNUgHHRCTmQJMmYLPqEkafzc10EWgs76JQ
W20DXgda1YgnlVoUitzTgqXRHBHPt7Gcp6PUetslXYAWB8AFUJ3nM/Xl4YzCvgvS
81DddybyQMWnb38LyRoRseEarrjHoDAP6XuJWHHQRnpeGxDVV3bQl8up5F/AeNBk
kyEfMN1thzE/bFloL4WAE5myV3ROciBVd9r5kqmqsT4DGciO+AVAKH6AdLOmku44
eWQSscEdtkBwdAWGCnkfULOMtEiHmPBuit4xk66anPYVThrV1y7IFtsidHxFwLGJ
sx/PGpvCrbDm9Smp+EG8ARTJkm2BWanNowlRX5LTKeWyr287+qonBMv9wJ1kUHNl
qE9iC70gI3yBGSQZl/+Lyg2TES0PQcdAfID+U6mnPn+7qD5cUpzexuexrtdtUS0q
3yOIkE9rVIndnm8KLRHkquVzT2VpX7noFWY4/br8ksB+aGUHhQAO5snRzkAAA4gR
16V0o5JZ9Ny0Vo4mBh1GSDC+HmTki5d+CV2TkVMl8chvycrWxeNnkxF10FOYTyG7
BG5dgaIrowiB8Day/E48eF2J5m6Umpnmhv7xim3ZQVQyMKpRgiZ0t9h1J01ebyGM
yKl7dIk0Mv7Cz2kpRdRSD7+PbbLgmw8H3OKitLNqWRE=

`pragma protect end_protected
