// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mjS3OOOYA7nqlibUdh61XuMullUdWfjMMsJ/EgwVqmSShwVRuOlMuD+mdIED
jkqlN3En4iJ0N7g5/X9h9FkhjKQcNIzSxtoTFXuOmnPCWl55m2TOVrN0HSpd
a4hi6Y7AlssUZD7jNRpQbpsig2iCU5r96Wd2aI09qhx3pRULPrzFFF5PhGXC
PmBiV6HOl2yEY1gQaCRWvZaZpjO04Mv8XjSPkmuyhpV7YTzvbVIJRfE4eYeL
BBmCS025AaAbzUFZpekI97CsduqprayoE82XL0apRi5VG7f13fDQWWJc0kb7
N9RYyH3cE3WBXUI6ZWc76G/932LN2qq0/NlblEfbQg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YMQxe5uSnZ1evNGoHmafXWfAEmvyoa839Mv3Ve8pfk6+J45kUV7jexsmy5dt
kKsfHGmxuYDOF7cOg6D4/hAfFfeilNMAAgM0RmHBwkjDA0jmQp5L/Mf1KU3A
QiDCvhKFlEOntCS0MnpxjAg43Affg6gesyhpkzyNBa6wijfjl+ojfyeMP5TE
LpPD1PSlOFxnde4Bh6qty+URhRUWSspHfVKXQseNLIkFmW56vnuLDKntU3Gz
96IjfgSwdbyVyEfgRwRHlNNerHT9aZvQpNlOwGN8XZIB6z+9ZQAbERI9h8IV
L2yHliKawJsAhck3XuENevfn+3Uzb6wzL2c80JCDsA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b0r2HStdp+ehlSs+HkdZ8CxXi8KSHexINVg2MfxLxDEZYkJ0RqHKZ+jV8HQe
mE4nSQT3Nd4Mo/vjfOlrk7ygMgoUmhs8ACJeTjpNJg0AecVGQKH432XgxizH
4xH+I09SS7aZXE3+DT77hZPeINR5O/Bc6TWBiQtqANRZCygP9qzburfD6O4t
oknxlee9eGtCAfrVTll9qg7Ghjx47YdITrQB1c/vg4YQbNShvsNpEAgzoy3t
CvFCaEBUFKEkOicBlizgBy8LOl/1fU8o01CrIP6Xba1dc5Hlr9qmdcUd2xMB
shYrHc4Up8bxRQmNH8p3uiXU0xrMCUUYf+0PoebkcA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oA95jmsV74beir+vQDY82LXvun7tCvt+AkpUvwiHBQHA1cNNDYFnkut9O7HI
aFmauRVrRsxjMtKZKd5yrb4MeJzCKSRSZeaFhdS6EjizbeXdTAsGEv9U/gTC
h34eBr5wzjXEP+hkGh45EvMiLaJ4e+snPj+wJSDnPe3oe0xPTiI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
iOKqdKaipBaU3m5/w7aL4bcFlz6q2kzc9hX1EG9Uw3VLdysxbxtjRKlc5AOj
gRGY20GPPoRSdsmpxAZw7eKXZP2R49L1oyadKhedzhizU+F4Ec7JzjfK/ZXU
Dk29Z0cWGBTg7jW6ejIGFhsw07VcMEBAW6pf7TtwR+Dcct4iD5PWsBIH4KXa
oGCXWcIEkKijUkamwYfvuN2ic41pnA2/WwPSUrcHXKGtqDeUdEA9mL5236cg
YkIIGX3ffA2h2oPqTi9ccnCG4dxReOB4FH+2CuEWmTAPJz628HExYuE2SRa4
5b4QB7BXTkBve51wK9GY4kQVn8Fc5uoMc8P932WaGxcUH4odquG/98ltPhZp
Asw3Yz4hRl0F0vAU5BiHARxeY1N5RnU0sM+nzSX0c7oezEcIK1GWWuTOCDFG
IHzbfPgkipXjLgSQMYRduhK0Wzty+asfNTOZABbtWIpTG41uGewKI4hieGpP
7N57HErfUIiPsHw3PvCJBdR7sqH0U0Sb


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ha6YeXPGE/zTyWlo6vAqEbRPHAsecrFldRN0FSf15PzjznjPohU92k7kqqPw
bTszG9WRvMw3UpSGJW7xr6OWrX/nBKQwYfi1vbmt6kC6e+x9+Ob7R6wPxHxH
xYOP6km7RTa24sBSuNPHLD9oR0rMrfO2KPrgckcs2inH76i1yK4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HpbmXlyAwa/X3K7g+yeOLBHTTwJVvGT3rig82Z1EQyi+fr7Ru336srkeLxH4
QalR4ioc198oIHxnwRA1ZZEOmyV0t65/5AfHfofRMTELbu9fVTNDXc6pi1V1
rLgTVMFOJgVMpOLh7j3O2fb+XQJ7n4EOx1tmcYtBmwh1Mr1G99c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
BSPJfQrJ5bwljT7VcLkG5vUY507ZM5hNa2FaNNLC+clkKULtU2D0XJvZREjF
57f082R8JuwCIBP/SX2HaXpW6hTaEuD5EFOyY4vtlqbqxf4dUiR2Tuj7jz/h
+qaQq2TP1owrT0EXxH0T/B7qg4bdgsYdDuCDwjQLGv6c6ozwGVwDX4bTBuHV
2XNBwr84UgblpTZ8STgzs0VPq+CBYRlx7VQRo/lBWwKMvXlyEERiPa/bzvac
EC72Grrho/aQXXEXso7lMrwJ5I5+Sx4M/hecRMnaNky2Ua38DCNsG071tOzT
C/SuqEL9sdUm6EkXUIsMKATov3NL7yjQdXyzmzD+/qqIeO5i4UgBzTozZDPU
V0L6Fwo5Mshb337bbXOmLTPnEH0P+/O0c9qkSY87k8kLiajxUDBwlRv17dmr
nxL9osV9z/XKGYAX+88Gz/544xr4n0mnaamQWEjJ6z5zO0amL9gJJl5XNrPd
1oc3qHdMMVB5XwABCgAYKz8fAqThqJKeAltcIX4bJ07xCU7olXstQq2q8+Kw
Zme2cAduy+9huMOY1fDTrGkOP5qF3hiI/zIqPCNvxOrEEXEIngf61hFlqQ8c
cL6P5bWN9v9/Ze2evtEir2PB+3DeHbmuY2FFxuRcnKGlBPGZAjHeXBZyp88c
iDRjDMYVsUKKG2XaeiqamAkP89n3CwlqzzR6IOxuCGWyZKiZTp6Iih+OWLvo
NOxrsnBIOyP/QPGVYb0zIFD+zf+sfTqAz0Ok9JyFOxqTSm3DubLcGxqUfbyh
I+aonzFjaYth2IkB4Q6Ylvv48XHUqsdxN/Xfmt2CmHmW+olobwdjcK2/2JPO
AhGIHNCOS7nzTC0efeYdReriKdApzX4hR570PQg5UXA1oPlGbggAo6CF6V/c
X2l5mD0tW6D4oBFtBoyZ54XMe8Kgz8jy6GjQJtBs8XeWYxuYDpqoN3GSHTO4
pnOjrvcV9gTUWt7niJKcpe2SeWOAXpq+T8OHb47UkVXbybqn7hJWZJPv/b3D
hswbpVYE10B2qWA9g1ffXNHSLZj5Rcwp2Gy9gBSEa01d+QiDMoDprvT33Eh0
7DKFsDbRv9bz4JumFazhGC44RoLoK8PqQoX7xnDdV5hc7CbYJ5e6mPrQWE0X
f5d5uLQwk915f+btm7xwZm6Ka3TH9ZfZvd08CqLjC+3o8lCNILlk55Z23dy2
wSIMTD5Us8UobE4cwTM/fHzoqvqDtyLt4SRDmTpdb7Q4WfgUBusFOshmRTDY
s1P7ub8yFq8GiAMX6kS2HC/8Rrqdf6R6kIPg+KKCGECtfj4tcMvIt1x2EmxR
S3/il/ETADmh2asIFyYFN6nUoMwiQOAEulBqDdF066LaMWq/O4erSS/TTD2s
+1VOWY+1uGCCDEeco5ITDBpMaj5h1d5Ssc4pf0FK/iIQDKgnMfvGIpZ8Oa/Y
UfZjNasFHgNm0WufSakc5qm69GKRByUFkjL+D55MlI6eu9xIlI2l1rnmRda/
1wL//3O9RWLSvK9/x55ayNGiOv8fdFEl95SFHN6RT2/G0W/Vk5t71LHkPwRl
B+o95kX1os3H6po2qZxLnRw/vJ546M/msMa60RbW1mkoMliCZhDlvaM7hcLL
PBmritz578CbmzOvgCb5HOj7VOLmdNPPFlctCrbAEaB7Bfre4z8IgYKXzMNo
Z7h8hVaeo+0fktGEH6TfwQ7fq5QpUglnumtkX3IcAiMfHFau/GmE4QUTiDDi
XVxYqjB/gSXhocg/rkm5+m3koGiedH5LVx5aDpdsS2xQqEsIW4eZ4iewvJsn
1nVD5sGD+gZaJdHQsz0a4SDniAdxEgVblisJuHypCZEMFs+mbu/+CjNe6Ks/
5NtN+PaSkH5kHTiltNx862ZSVxMkcsIkqbmlabg67hDjSRIP34DelW/J6iwT
bmWQSiImVm4eFjrjGzSuw8yyFZHTNAti+4i4ZD1ES+XTLedQ+QbM4jdl9vR3
jqFBQE7LJ/6ks7lmp2E1Ff41o7KBXPf5KTRAcauuadIfkjoL6QZhjhKfzVKq
yly7tJZmyhQ9MIbuiz5QpR/jf6qEvDiq/wBuIwwuNa2sBDlsWYye6eDWOqUE
JTpxpW+llyDdwV/AbaRdsH3p8legm1SL9qJQbxh4aQmFBorN49lRd4IiOLCH
97R/URHEFIATRrnx41t81s22zcvAVYV1fufTfjPNdSXx6tpHaHJ6kyNusWmL
RerMlgPtcsHrUoxlTnPCOHsDIJa3yDZeZXxe4KhwAZfshQoJdtYgWeR8zLcW
olOYPPRO/qivVqyPtbqTSzrqLaBVphgT84pLF4Zy9o75gSNrz+G5/vK6Lz7n
jAUVyF4g/DuJDmTz7aEp8ePxwHDphVyqIGPzRhNeC/iBmCzBNRa1+wcoSjg0
+DiNUd2EHLMwcH+IEgNYzvDhknYWWW6WSVzQnIKFiCGST/4KgsWElv+9FSzA
6rKLBTDxApmv561bjj6Reo6B0Exag2oYp6N/Ngrh+eqfvyB5f6UgaQfk3ZR9
1PpifdO+Ewy9ZCNKvLeknjZ1F7+FzunaYp+RA2f7eEIbUJ3TbTv9qNXY9BwG
hDDFh07J5YpV04MIKh414mJaAOarhfSTw89jPTaKNsYhlA0PRbq20r8FO9DA
zhxOxZ4kCuwIsh3TUjb+ifeGAA26XivyLwmDzqw3o4MaYyf2UywOKl7+//aM
XzGuvf+p4CNM5CAVon5uuXW4TKDBMbyhc67P3a5y6DpycbSRS9p63Skvx60r
Hkt4BN6MAQDhfmxAr9lQ0/8xEJwKuxd0r6fDohPr/e8xkgy7eyRbifGzshhd
SOAUSiGp6j12Ze5pr2ZhVn4+YM+BJR8vYskftZFdmtrImumdPPrzBi9biJjn
ga8AwkKuWhwGSp7bIh20Yez9+QmcTeheDDnkcycYL8O/cCpRA+p5Sur/6IHV
JaX8joGsTAV1aCeaGQoU97JJ5W+yhDkb9T+xNn/Xzks14aWaoNuQBQ1+RKz0
/8/R13OJbKC0Q56SURer3Lj8QJMKLvGT0ndFUOipQZR/d49DOPA1MrtowRwM
iKG6Hb+W1OqDfQ/fCmIaVs2jrgKcdbULrBNVUwnyY4k3wHjqaZ28FErqZfkY
bQ4Og1Orajm1rnmF+tdH7K3zS1kkvCVawJ5y5lf0niL9ywpUfKXbfm4tpxf1
lNdlm7AOZi7anLcJ0IkXTLVARJqDU3gFiZpP2OEI0Ryj3eQVq0Es2jUlckV6
aNveMrSaJN1EKZ7cEm9iNxlU6MOTyBNKKr5pEHFbB50hevsu4x9Pg/esEHlQ
0yHhvDTJrUbMSCqR6N6pI6YGcWCWAmF67cUI7oWrHmsdUMiowZ9F7u+IdEj1
xRJ4G1ObN+Yt3tcqxmL4M8pb4Sd7vUC0mLSlE0zZ08/P2QgKGA6u/znKWwm6
EPb9s9naHZg9Hj9Q/o6YfvmSfh6Ib9rQucS0squObMGKc7gqMcjIFKkPh0pf
loRQ05xxSRwWz2nEKNqfVkLRnQjZNtki9pi6uhbDhAgREDDH6wqAcBO12nOT
/CTES3Ix9tvgV8buxizYw/DVe8hRMCdrzFKaXczDfg/2Gri2FlXIPMjPbsyk
2aK8lwV5KmhClFZOtF9aS4EBTCcreayRqjPpIPlROu1rt5V6v+h39gfBHpth
UJ96xg1H6Mff4HITz2ijv7GxEHJZK15FdjmA8quIUja/1GahVRyA

`pragma protect end_protected
