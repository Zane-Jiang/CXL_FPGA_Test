`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
NzyN3jkDex6ua6eNiCRc8kR+j/c1n2xI2KhU+3s9fGKJGg8dmsym1nfQ16BFGNsO
ON0jgYjxq+o1JD8gV7TU2ESBRY22ZeMRrg145Ba4snxXFtblTG+K6bpsKzg9YnPS
8AQzMN91F0dHlk/Y7KJZ/7s6YzYXPfqOvBqoLbIVkBA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
DaMY+SDRRAuuRVJFg9MQwLMaWqefK53lqDMAP12nynt4VK7BXstzxRweovZBHIMY
4aUVnjSjiXl3kF2w/e9JzdqoyreDMKCM71ibIYnorlS4RJHpbBGdgn3t/8RSiNto
BJv9lwtbvWATwGEbydKc5pyHOOYKMJCgMa0qkmB5lAcKVkmIVedDwyis+pFI395a
knfHskA83yb5y3q4Opog2yo8A6Eof0hs/L7IHuSXUZAxLnG2rEeJOqFRkU0J7yhz
PDtiewvPbzjbv0byFy/zX72NFvCI5JHw0s2M1iP9tk/NJ+4/BgUiZ8YlN+eW6iVE
SmPUBcfwHR+OQXDVSDGNAo2ulI75jBOafPKyiky84rOn4K0n5riFA761PdKNA+RB
BVq7qA9JDMMDAx5WGIdqOclA3F67LQAYtScNWIsfQpbM3Jv3pCfW1Yfsa/lDWQpR
8I6mPnjWJ/bSeX2JHv6tGZ7Bg0ursfnj7aQUJfhldkaeCAAcsayOFv3v5O8p3967
Iimh82eYa1lqYLUgV4cvVQ0El1NSuSGQ02q8rw7Ea29+6HtPiMGmS3ghPwZzuuG3
vKvBzRYQLOylXU8XS/pBs1tWTrgVJq1rKJgsQIDxfcJ1lnF8nJCwwQ3FR4Ww5pTK
UnkP8QtuiE4i90xQ+pQ51KgDDHnv4iz2X8QXUz4WWaqYBKG23NtMZXPVtH9aHP34
lNULjpEQcpu1R4g2+zwkbcZLGmVPJ2d9PRg12YqyTuYzvxdQJ1JV4ESQmFF0gnJE
Tnv2rTCNk7rMeBfkNHxsCzkvj4iFF9uQwiqISPqg3gyc3qTphiIzxXfrjtiTcXN8
45uWZIaK/em34EV4Nm7+9/NAyo1uYOt4f90yRAhIvUXwrkUQTO9wXxqhK2bqheCP
gg13GOpS/t5qdF5ekA+KP0Lw/0mN0p5JeaNDmh5fRmyevjVsdOXFXDVj8akJT32V
j3VidB9PH64j5B/nsdNFmkrf2u7GXM5HfnaF5pLH3l/v+K7T5d2BJW7MDGUPwKZ3
DWb2oNSjCtm4NwzPvOiZDBz8lZ/2GvJ6PQg6TAIKAsZkaZx1X45mWDZH5+WOuY2K
qOy6qvphGAnwZwLNCDB/9xL/MNp1ZH1+toTrDYePmk6GszUk20k9Y7DHO5pv937u
ADSP/vRcermdQaRXG70XMvbem5NdV0mK6ToESd7xDa2B8PFaycUJrJl4IZz+cLZa
s+cjFSwNrm1L2JSqK1IPOHWQFeKjwcccMTVvPybWuYBqBvbgkLGCtUfuaUXC4mfi
KJmSkfUpCOMRhM/sqU4jDcuKZJxRiJYNEG1CgqzzcdeYH5xnoIDE8j9hMpkcO15O
oPPww9tbK2tsvoJrzi0hx/SDoqHlrWHBFc0BWC/izqmRsFuLBHQmkTetZ9X4qx2K
x+81Un5bzBVUgsaVQ8rpSks/z+fa7liN4Pc/JfTZWTPFBAABiP/TXuyxRNu6g+KB
17cmEFXHfZF6NPgZB7AySfVAOjTCdCGfiOYFrWZWVXZVjnCw4MAUPN4+gflKTVmi
Mvy5Ix1Hg1kGDGZToICH+SDeCeRdUi4wXI6MVeF25V1P1wLOhESPLEbT+TNEZf5f
bYg8saxr5GG/cYtl03STg1CZwca6YyPGYSjDf5ItrEHAxwWD3o9J9Y9eBAUR0Vm7
NTxKTGHWLZrKmlDWYOxuJqq4cOaunS9uKWZiP4DlyMZZPZgouFozR+qMALc4T+iQ
5Iv02/WozhhuIkRKhWHP5Dfw4U8aV6k/nThsIqpZmUZPsfS2c4Wymu9Pbez9T9j7
WtVoeOtOpUfxWPtDTmt8EJmIK5LMzOareg+r29IwHmI34ngTtnWtShnoKSQJ2E8B
LuSU7VedNWjS4LBh9OLG3PdO81+siW4C7xDmSh4dHYoL7mGgbilERJXYR6GZa+A/
CReZvr3bvyCP871h241ow7RXkO4HLcPIDrVwJuBiBnVkYORIJsQL5mIhgRCSIRq6
YPWuR+wS3K+zU8Af6okl2BxbT8n9ot/I5fgqzAJO7DjF6pS3tDuvt43OVFInQwMW
S8Il02jMb439WK8E3WurW2IP4kp4jCHlYEA6qrA7tTICm4WCTI9m/lQxnB1cGOgs
SUj39o8ot68YIJMItB1ds1wlpmHlLq4qwrPCvWwe1YyTLoZg9eVjQkfxCw81asU4
B77NsZX4B+dCoWmbJWjnaw5TFu+AQ5gplxBUTsO22r8PrmbIbO/SFMcALFK17qe1
VePqXLgHzzYaIp6Tye6feYqidXj1NNdAGFFbnrZv8L8FBEv3ANoKb+mbwGfXyr6Q
0drlMS7AUCLVLTQsD3wCD4ROYvypHKsYD62gqjkNvdeTdPsF9k83Q4G6VozJAFCc
BWU4hMyeR5WJCIxV60VaXLnETaa4SsMfAr7QuJi95yxwI+ufrd/me4EGLcGkhjoo
5eLx01rqIwmo9WfItLiZCcmZoFFaMLm+cHOD+UZhbZUlVtDM/ZywVyzES+JmuEaT
yifiCIjfDtVtUY8TtooiPu07g1USPynGpAdGgtjtQLONONnS1v4l3ybEvMYyqY8k
feom1WwDgBX2FsmISugAaucn7or3fGDzXz++z494Gl+t18X0YtnM/w8N69qEp+W1
dRPkL2L327utV78WbttRu+pYDmpMQk65VdDZKfnI+82ywR/rrlzIY+h063Ed47wQ
DpyzEx0Excto9tQVv3k7/TvXNC/oy+YLbzt93vx50qa2L5RMm0racQYJRt6Y7eMc
oMn4EGnFyAcEecZ4lI7wNX6906Z6abqhwHSeztdSjp3RMc093+uWNcS0lihejdzC
upjRbvbBCMAwZz5Xq31t3rA3lWdQESXYiOHc5OqmdHfDu86i1ZdCS2eXhKKK8Zyw
Ro/BaYqvs6x/RlLdOev7jts1zLfQnutEHrV2nR1rfAriJMSiNI2b1Ba0EzmuBSN4
xT54DX4CIExk5b0q+dSEfd2FclcLE9IrknpF4SnvCBTeZAXrTRc/Jx06RlEqpyFX
L6DHqP0x0Aw9ni73Fg1pfq4yF6VviByWAKFdbecVlUxt+3P7/nP1tr2F0zpPtHvC
2A1qZKPlz3ElwQcPmteq0mvV99Ar/bGGcXc8rVXDeMJa5iqtGW50q8cijSpKanVe
csnkT9f8SaU449/46tMx8EKOdImGkrQ3387VZQr+1ICvVj0j28qBN2XKgSkMOK5y
ITD5Zw0JJRZ5hJHf8I9HoEMTqnxZusrHx2A7UlX60XQE2nCD0iEYiwcPkj6Mp3WS
7wnjcN/hvPXc3RHT7oplny/PEIosuiZsPwVjMvlVtBSRyfW7YbsS04xfJAO4eJ9T
U3SulCNn9p4iQzCMkdxBglP0ad7QSftP8Gvnu37yG5alCf6X5zGUqJYAMqkBRSh5
Q9DyhBJWi76WO0oI8Tni67v/4J+r6QuEaxFEG5PSaGwSGIp0tBl63Pe3iVUNh6aD
W35PfJKTHXXmFlo89kOetG3N3cbQFpRyJ5ms3owieNTzpMTEQhCVR/oLzeE1CCIk
C57jFpSBO45r04bp0FUvdtG54Y7rvMjwK0EQ053fmet6QGnJZaU8joC0Sjz9Jdbn
GSPjfO/5WouNVSmUA5XCAPPl6HuW+ub/6rcmJpaLP+CWQyb5a82+tipozZD2U/3P
zsiyep7PuMxi16MyqWOtulzeYyyTSClgdWMhHdn/Fe3c5NJO8Go78dJYFO/+TdO3
nkGJYFE07F9NUxM07s0JHyariR3/sPIUvQwx15bjE2CMVeb9BzWN4H4zdkRhsRCl
1PDQMzZ4BGVfkxFLxzm1nlkkWiSKbCns9IfguBrXzSn2CzmECw2cFl8Ql5O3waR2
CUS+HLaeYiqRtd1QvQMjJ5ofYj2v1FuOPX6N4+D91YAAlQrzwmOuqMiZyqANUpLv
bhfUhzP80oNaL8qt6ggHz5kLZCSzQLtd7n+ztda4mIAc2qH9rQ1osZZrsYr++emA
r8yozDgQZP4GJV7MVnz9K5X+k05HDBa4FJ2EUfVem+GCoQGZPCVVijEb7qUW9PyU
CemOO+yIuA4/F292KXDUEwfT/Zmzc83u8Kbwxj+b2A0rzw865EYagvh1u1m6IMdv
jBPW150BObrHc4L5kpGwg2HsQRi9Mi4I1GygS0M5j5kfDBlh4VesSmSK5Ek/BHoJ
+ONAyZ3euxXB51UZ0WxwPNLC4Rk3V7Pp5nbh2kZmIRGsFNIYUZecINN5ESazhnjc
iFgN4GlZzFgz/fjrnwtWRCt6gGvXZ4q3OnNfTXanUY45zeoqA8qUN36SLZCLdmxh
oQ9cDsT+5839EjYGLz1zQ3oXOwd9pqXLXmaKiCm2647o6cMCm7K2XL9PpyuJXLWd
EPyGwaDYvXPPrmwG/oJCiCjlbEu9dJwi5/LZxy5U8DZBthj4Po0pSpZZgrWgRe5a
8aEvQi6yGqDTEzPh77jJN62OGtOr8ZkqzPgwMlXKm4PU8unJN4XsKUt2Zwtgwbzd
fOWU7zejZlQeAv9y8qJQqX+tUkSN7a1c/uTZ+Ca3Gm54xNvAwEZQh/dpFZ2qhtXL
1uACZYgvagdP9swIORq97jqeHikhcmLAb/LJjkfbeJcDhU0fTVp9Jyjzeh3Y89Fm
qmd3rpLF5ViGiafUstbW7Ua+DOO5jg5IqMT7g0GfRPNbZRvHmEBptIcxKOoPlX1s
8dUrNgxIUhQryBbKge7Vatpes9InHGUYx12xU8w9A83N1JypSMXu4yvJXPN/TKa4
f6XCX6HxFCAi7knZ8JbOCeZwB0JCLfuEySMAAaWTFKNqwldhWnBPZM3XtyNh8Jp3
DuoozgZV122cZkMXGMpA9Npqei/BRcE1Ue43C+TjuEcIyjBvZbb4ffywhHx5Kf5T
+dOHhGOf7TDFaWf93zawe/Si/LgMnWyzxIlWf6bKJziAv4R4sOanZEaxDfZ8q7xB
MsORgSW7gT8oTR52j6J8MSh2wNCbBeKpasrgh45aPt7ZPfDPm8nPSpqp690BEOvc
rOEyTVzxz9nF16IgqYxFbdYCyVZeiqgDK9dcBdkZW1mQGlbxVADLVQO37Ma8muvj
g+8Bft6bO8bOzMzbi9r08/KG66rL3sBCuRupbgK4agbUqwA4z6eaBK71CeGi1Que
D/+5P2Xfnadci9QVcpJWa2ILDBnbCKNQPE8R1WF4TQbDk8QX/us/6XYT2qS2Y6eF
q/n4ORizqi2xYnZiliWdlbNPBW3RmCZsJiYvx8cWIt393YhtRFujboOr93395vIy
aE4aEtNk9MzulZ+UQ71FeFeYQ6D4FW8j0QSusVHALdcua1/wdReT1NG72pqINeeS
euLDeR3e+SZhCTABfG9EzpxLp1Gc7W8UTnDHFucnhIL7YujhqXDbx7oMc8OKyHvq
IhPws2VqZwnyJXFUJ1cvFwycglV8R24GfJY70CgwK8txUdJeqLbSgEgPakFPc+7f
XGn1eJmeNFUBiZSEQZE2V5Dcl/80s4pmvi+Uf4y/x+CdH+LEiR7OPk5WTj7Vwdc+
tbSIsWYez9yQKs1Q6oxB/34MzDz8e8lpH3wn+Wb3V41ka9cIa2xE4dLEfMLm1nxT
BOiTTpXN4931aOh0xcxsLFJVv/HAh6UhDSGh/dU4TZrRX2W/LhxPwD+UKo+8A31H
cz08st5uWw4304FkvYI6ojlcljuCM9AhCD2Sy1+b3X9ll0nsxdsrwydItab+b92u
hkt3R6b26V5CmfisKD4JJivI/5EBODi4EPWrZdLKWYqL3DRPCM6GbJv6EW5xnl8H
ZGtHU5f2A8h8iZW8Zo9g/NIiSxX2wmlNJ4CHeBt4ztLucM4Uq0M4DMvBW89GhP1n
Ijt0DwS+SyakvvHDs9h4Q3eREFAdt9eSt7xujYHjoZvI3c9mVBIA11G+YilYXdxP
PwfrZLFK4Sr3VNMCEudksKKrlA9lAOiM80L9568SqrB3iprTHFoKR63+6fMyxwCR
B4u+0022VVhU8Oob7/ZzsIPScTag3yoGWoAJktboaxDr9egplWAD+I5QPTPcTlRW
PSC3E2E5Ew0IBbjsJ7/zcExRf7b5ypMjdqdPZAzxrCK6I0j4g/6JsgUxZFezrG6F
N1+7bNtzz67BDk+1teIjgEneBJeFSRGpz8Dc2+aEx5UUZt8JZin7tanAWbppzxdT
a/jmAoTwcTaK83k+sG7BObd5+zXhuIhb4acpuH9+KQcEXcaViaRfNh+7Y2L8BpT9
Lh822yh2tg3icr1SMPrtaLLuCFGxTaKw4VskHvr7HVTTfNzeDGSIJahNhga7PKcT
y2t+9J+a0SNF9eE+SGYZ5sjorhbVqeVkCzg/0LqLIRSE2VMaA6Fi3LwfvvzrVBpl
pmF1lXMaX5N0HrA8B04YjCIV2qcK+CIHy96wS367nqH8s8m417IRD5/bpCbwJTyV
5oxeqGUDOuo8PCfaRRQXsjqv8VICWRr30sYFvdIwX7aBqtRnwKbrW51dGR0LPf1Y
1TctMVvx3vDeN/VX4PSMAi9Au8+uCZdIGqbzx9GcRzdvCGj748LV5wtysXpWuVJP
JGdTRmvcwsim+naQ175VDiJazoYu1fktXwE02JtfQ0L4MmQrR8Me782qMKjY/B/5
kSiYdQApln6wuYw3XS/3BCSJztSAP9BqbBmd+YodeBijMGfpbs+u9AKvJUGPmFtZ
AnVaa+MjmKTAF6OI77Zv2O+P26gOEjZtIpeBuXUQm7hUtzI9PiXVR2NIG0ESH+ix
l7prOam23YHfUl3rrXc912CXxgNNUye2ccXCY3fGUDhG7DMw+egvnKF6kmVDqhxy
9xUbSommZvRbe8690q0HsSKYuseFnxkrzJfWDjf/iyW+LIGGTe9Op7AIm0im3TWu
ojD8Uo/aUGyOPLjZDNiLNn4ELhahlUdL2L3Mxjy/pJWHqC5GOSa9iNv6z1YEe2in
0y5QTZ79QVlM7fD+4m+Kf5KigsXRipOSVXnZGmTAkBSxzWrfaPhvgpZsDgHez68u
j5Ojso2DqY7ls6U/rwPo0+LfmyNUos9Z/8K/K7EFRiGMqvClglW7v16F/OlLgaz4
L1kHlksiDXBnhacU6RJJRvT2sAIEjshjV6N0qOjlmcPE+3AqagnOBlxoTxSm86ma
HDl8hpUiG0r+HXm+Ohn/hJo4D25ZG1ZS7HbChcEs7jtNCfZUlhMjJqoWv5RmgMvf
Ww5n0iVFjgbFd2dAM6zAQmNqVeL40CYlc8s7S97P+Rx4IF2fIiWCcWDDGOqGX90/
Tyg2uTCvgl8O7iosmYqkVJ8/RCV7BVwwUieZA7GtDkufX5eCyeRTUahM1RlKwlPO
ePpYSw5dCb0PjAItsXuKGctjbaYWZmRepYXMW68dd8FualXZkFMEB/uJarV86CTN
zY3dwh81j4li0KtoUYtaxLuJP2M1Qn0fu3BNJ+Mk9fAW/9rDpUWwtyQEd1m1YV2g
atJWniQ7PBtdemTa30H9AhhAUeUjhB39nMpBIP8/uYmR6lYQtcpU09x4gWl/7uxC
8UVRwh7xmhuBx/c/Q2odxRGqS3yfSHG22UupBoX1pNdpmDMYunPDVXxHsYzm8zrE
AVUDUpG2KZNXAghupxc44eq/JxnmW262gkWuDj3uE3HveSGYqhGLFcbBq2myL9Jf
Q5g6fXnSz0cjBbAXlHV7fBD7STwaXMPW579Bsryd7mFhMAh3qhGgd9dd6+TBK5F3
Q7HfA02xJoQP7SH8pHQmtckDD12xRIajStfrP3RSWV15sS/prYmEXtLgKEZp1NvD
GS8WBxS9p/S1XFWCW+GQMYZ9YmOiqsu9f6atmAuHToyaAUUZWiAcRHiX9Az5dNDZ
WbRElGwzarE/Fc7lE/Z1/fFtIxrx4lSrFkZzPUFYe5Zinpb4Ml8DAihLlT/E98h1
S2Cx9Qz0CYIlM/5g3oNgQiL8LblURAdBO8iv7woKsFb22kdsO/uM30XhaTe3Dn5C
aUPYL0Vok1THR3INDp8yFDn723EZUq0MZVuRMckRQWQzWFYY4i/cZ4aC99oV7FLf
5nmwWPOSdTVoSVu5f/IrlusXX/WGKASbBcL0pALksSYg7kX3lpuepRS3NxVziTZu
84iWRybrmF9+SjUDbebvYKsdmeVA0oCazjs86Nu5jJWF1TW83ppTpV2Ril6s/jDg
qzZR6TC64Ct2Ap764Yu/cHF/olNaQZWYZOZPsnO2FsO+CXnmws8XBuQpJF2eeJ7K
ja1KCJWKBeDeOOcgTc9xnFCiZAf6uCzzYxd6QuIaXZoH+FA91ydqFa7J8aVnfMW9
NFbcpw8vt4RyHJL9jDFvkZkSm46s+UrgOAPSI55HW7XsSuYNupEdR5uMilie8Wj1
sqVsDNE6Cvy/UG23drd0G0jb6MBhJ8J5eCacDgqVxDS66/qslf29ncZ54Nut9P5p
Fh7AZVyziNUdpE5aZAygYXhYKIPOOqs/np0yqmNuf2gc/zPAhy6Bwl3te+xrMLax
iqsTN6rwYNO6UwBvzOqYNaxIQGgzrkKe/9rqmnqFE4f3hUArm3lLc9Z1oU6KNNKT
fMEOPfZRMcq/kDOPtJEN0rjdmJkkVjgeP/aTamuDqQqU4GZ8CHIM56kufb0HiDkJ
2KFUf76J1KP6iGEkqY0SMQG+4QRA9arEm0rzJzDmfOPWUh9qz65yuNklbXuXDb7y
89mB6Op8JWgv+GgOarmluHgw1e9F+w5GujAXePYZPlBvufo+svZ3Tk4HqSPsYgaa
G4jSo/3l1wrXMrdoKFGsChh5+6hp5t/0pKyCcwpLjSYr7U033okGvXc949S+PsGz
RRGCZhlUXC+okFDrQih+09mQEk2D2XMEo9tTzBYB6khO53ZQ4DrOGkPXPTDR9jBX
X8wyjZlfhZfkFN5HOTnn3QIayZgmIz+kX5JwZ9OUyUlmz7n5LZvTwvMQ6pmI+vuQ
PxhC25Fngsqe3XbC6ftWwXxf6hdWH2uHjUFmDSMy98TJ4JUIr/pQktBOW6ckjQw3
0mzFKt5WsjdOrmb5XR3YoUOsEnmLhUphSFU447S01JTabiXtTex48oHVm3lCYYQ5
Lx93yLy/Pc/SewrS1NsajlAT7qsKdvUWr4d6D+yxhbUtVNUBhD6VfnPAfkCw4f+G
kBfuC33z1OkK58qxoPePhNLTo4u4JoQaOJln8M9ciZylwPxFZiF8PCv+bB0dMy0+
qalafbvoM1WSm7DoBGtk1Vs0D9kGI6Bn/MHSayBruwB0t99CpHDE4FNdSJnJdmRX
Tuw1LJqgjBNcfDl4TdnP3xRCeo6jDkB24u+QbIe0QBHNW6NQzk+xvtJXxsphlY1D
ajZHUWeyo10RaWi9D+6EPG3gT8abktPCOLQsQ9raxdA0QLdMiiPQH0GhpPjAfLJD
NX4FJQgW73Cbfd1upFdZnyGdzb6rLeJAaF5WaBFEd+PFkVEYevfh1NNNVruAFRel
RYqawmc05mIL3Z83iOBljsIiTmU7OD5L06cwzpfK6uyBeN5lcVEujh1t1Dpy9Y5r
j7hKvNn8TsGRCxH9FB9pmnLDfBLSWTbWXnGKV+ILrUtVMrTvfbPhZ7oiblU7GK7m
xPJQRnR9Xp4UqeMkk4M6h4KgFIOnLKvd/RAJIC7aFrwV53I02ciIy8iDPTFHdbDQ
V8UuUzlEi9ERhSRKapIkJOhm+VMn/rKUZzL4dQ6pO3E/xQSMeifoCwDndh2wbJED
g+vT7kxFBUkxvBcwb8XOSljIgIr8QB+dYum1Vz3NCXhhHzkGA+ioq9KwybsuvZ14
thGKVlzX/PbdhJ29F/Xk/KPLCVcRjNm3rVciEtN8zciVVsKncWnNNpn0g6tissOw
lrdcwrYjyGQBzI9TwRHpXPmXpR36TjiMn0FVVEXNATrYo5pxy+BdOyqDrsUTYeuz
I8LjrJpSzVsQobWlF56+8Ax71TbobLZksHvhXW1cau3WfoCMELIA9hcZpLYEFCDY
OUeo4YO2usg0CYh4ReyDaq+VSTp9yNRbLSY+nK+LqNS4QntBLdhe2Vyx5DDY8qdh
9SU/zbh9BzLmYGuOk0dL2KTyWpST/hUnBnBSav+k5j3mDcZruJkBo6OFHx8nIrXC
jCBZ18SSuUuTBQ/oUDMLqOfNbTE7vJtXOjZrsYYg+8t0haORfI5b62zkJL5dYbSN
KvfFqpaFV8cl8PRoIjZiPdZSj82sipgczI3urb53Q1mV511ud7MwBee62iFAbeC6
orqtTtIE+qrrVxloyOw6w+VxMlqLt4UaD9ZvQ1zrmNRBhywAgu8tJgQNnKUX76c+
Vtat80T87hI/RY9/IwjVSGj4RM9oV0y0KAu0q0mRDvU9jCraHqdH5VXwig47A27t
pAa/8AkAfyYwIDH7c9loBMKQDEdAYeF5nwOzNmC+2HI0+17SuY636iKbTQVgPrW8
V7seCzQ2rgTRCTirbUihX+PZjBOj6+yAtqcXflxlmnP65murE3K1Wl5a666h5TTx
PIJ4T2kLED2HjgBhMlf5Cv3kgcgFsmJrNpHA0Fvq1BTMRD9UpuLmK6tfn7WUVtEf
ItPz1pot+jovdw1KNSDdFKniIG4SRzAL9T8CgB1wgbdovvalEnqpJUdm/caU/mhw
PBN2d2w4dNBC4VAXUVXc7v8Dxj5GqN6T9RRqjaQLR36MFQj9rGNdWNnWOHwU8Uc+
x/ZCRy21S+MTd5W+OmMn2VnlTV/FeiE38twCUCLvipY9o0kB5NBo7X6FczghVuqE
Yi2uhnO0CQyKc306z4MQfKPxHVIcPX55jDSlGdLVz+uaOUBqbI2HJsuGQXe8yxRG
yht/Opo9RnGklcSaIoF1cfOj5y3ba43za1q7LURrXMimR1TlPu9ibDNJowkf0xMn
p2GuufHjmsTAsln6m6i0sJX6Mr2PVuyWeENVDZgLvwN+MOeI0tURz/pOeaQkfJ6l
/57NnJN7lZl1h2wd0dSBTcvXqmB152SVTKhna7FnRzi75hYF+v330AhpHr6mIy9l
EXrYodfBQ83lNkeBJ0/MVSGzmOJCrvVyc4mP7aZhJtFFWBO+E6IgxKtstdtB9AwZ
n9XPHZQAUSKEtUOe6aCafVEWQY73wL/lvDwP22FVyy5jNkIzWG7EkLi/WDDUEfyV
DHsZZC3C5NdCXq0cACpXp22LyUr81TACWrROK1e1yaM8/hJAhfRidS7IRfqHi2Vf
82pjZhOxA1IDFYbXv+tSI6dgmBbYZVQlgTKeztoejm1uMARngzFA1kRwBwfkFBHg
YA4IP/iE68qGV28f99M20F5v4kKIra3h9eGBI1z0x6l129lPL+JJJ+w6nTOQoaBp
guYAuZkruvp9kcfyKx6wO472atgMXCCKN3eFGI/nlxC3Aw/Hdw60CAB6L1Wh16CD
szjFNMpMCjOPhhvsTzvFc4c00x5f4dWIoNfF4azbVVHSpHx9OIhiofuin3QQ0hSG
n4xopHBG0vwq7UhFHHB7E/qaoXUdUV1yzBD2qU42u8Y=
`pragma protect end_protected
