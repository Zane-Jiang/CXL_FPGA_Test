`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Y6CNXwD1reNleXHN8i2oNGU+0wXBgfLEcia9qefiyrEfXM8FIIadnsPKyPH0liyA
czjw2CuJ+QJUZwWo4n1eyhdrtLAZhpUj/wYpLXGZRgWCuEhc3iXl8jnC9JwkGsYo
kEM99SLXWe0Nk02u9y2QcpRDVi5apayhOiRogsaXMUw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4688), data_block
EOqn8LRda1n+IRmkaU/rVMhWIyNuSFhjo/NQ910NnPmVt0RjpHNzfLkROYbauuk0
JtNGAKeBCST5pIHiHIfJ6SeRcpVIMhBuLBkSCYBDIrz/5bs0nbtpKH2BaGhdCy9j
GUMNSrGJ6HajWMiGx1q5aVL/Graz/50kWMmghbly78V4ffjGF7obHe9PyRWTWUEu
3h3CG6eVkjTIMwnEGmybO6Kb1LBCXpnD/A4Fh8h0daVQyIRTRhnLvLFxkLwyCVjI
1L/i6xws7qvAUm0Js2sO4NQBy2fJ2mY2cAlUZDKQDbbSJuggb/uEu+6cjeZ4vyWI
8vchJxH6yhJb5UKRnM7yec7nXLevEZjErH/Al/icj5r1T/4R6XbZuXBPqtAgN1Bq
B+L5cdXEF+RGYrPEcIQLdEwLl33foA+RLxS3K5UgqM+R8vzmMW3qBZ1W+sTIbEwp
DTIEj8ql2UUwDX99dbOJrZstfEcrk+rDHoiLpu2qH7H9H6XRqe6BubmbLl5OvQTB
m2I883znN3VC3ngAhX8E+sdM7m/OoYomvcDfxB70ixVSVecxB2EWDAbbVzt0+UtV
kaodIBTIw6X940YDD9NGHn8OZv95UWqb2p7I9vRiKFCbSWpHlMOtI10kJ8CvELxA
UkYDrfyF07igUN7NaCC+ij7f56SfJGX7UiQ7v9awD212NGhKreS6XoqA0Hm/x6QJ
hnGALsr76lkbQ/gWuLVlByTWESN/9k/p2IyZmxd4D3voBBKserjkmkEaHaPGzGSR
XYQ4to4Y/8FYtAeSvv1NXmRvv1O9V9KmC5qRLAlNTHLL3Dkft7MPuTWhu9/iB3Av
aXRTrSDYwW41Xo52k76PIY3ajmyW2lHuxWstJenKp7mVYxmxmkWwLpThpsFY6PaC
pb+07iXCKCvRYN/AdfbH+ucGGX6tHh9bCC0RdQdtHf/SffblhRIA9EP/nhD2ZKsL
+ou9w7OrXAOZLiTEKGKL8xi5uKtM5nXvIpds6gRA7hpoLSyqHFWs3PqSeCXYNcas
73H4EZLr1PuWvWebRyHUt9PBeVp2VHmGHjlPaLE8p+NsIOvnj8zMszbKSJNpdQjJ
3NIHcmnFp838ZQ3uuwUkW98FpSvCSN5lqGoPVtUH9SZF7/zLQIVKd1nyF15cYJya
RxCfiBwqPaN1qRRXqH2QRp/w7XH0mtv/y8nulD6RtRC4Dk9x/2pIWQjdjLoewux2
jytbvjhxglvVnHUjnQHcGP1TLVclYFbdlY5FpmXg+/XubMP9iO7irbX4pO6ARV9t
TbFmB9Zq4TpHeysw2aL3i7KtOlJeCcJp6L1ftLD403NkFDVFxs8SwEMiEFHLAMiS
JrIIYqF0YYEq+rvUO/e8pNdLQC6gDwnXPUwN7FupuzuP+ziEjhrlpB9mrnu78Hy+
R8dMkTFPZFTDtEdXKG4lH9AlNQTiinYiYdwh/LHgbdeKeNMXjE1i04QwxqElTOj8
5/zRFXkGhdmbXJgS+Yeu/kDechoFvtoYQZajlF7JLYTfPmENJUKzYZJHW4h2VJ+w
IuxSWL+RCvG4lFbl1/HaMiiWAiV1R8uUdJkRg70NhWOdo8N6zi7K+QNmTGnXx63P
CnMWBM9n4WqFPLVMXxrszuhGIkWpKQRFSRdHyyfFevb866grGcDTDivKN3tDXkia
SBk2VKOOkhD7wccaF98FJEMf6L/uTo2EuXJnz73dlGjzDlzpMaV1e3rctg6T3NKc
bqcHVdN3nSzQjiRLlTyLlY46gKa11Xpcbn46R0l8NrwaAj2VBd+YjHsvHIFn70H4
xGHZlsmedkxzjluP1NOyKtWpaBOTUlfU+/l4VsMjZRlzDuBZgRk3aoDNxrBqRgJp
njKJ3lJeFbeExXlefrn79XD3Y6j/H2O4I0TU6IiwgiazcPh5+E/vyi1qQUjMCtr3
FjhHhZP55egsGgrphbBUz0NWiYLHWmA7VB6HKsnyri3a4O3G7acmaNn0i1g/+Pcl
qc65C1yl9FlQqi5NOBKiX4G0BC1pjVtWwBIMktsRLi4wswLblTh/Pz0mtcM5UQzU
uE8Kel6p67vMFrSgEFZEXpOh6PkYhAaUeBPdFOiX37UMPE+Gc/lasV8AxG/6W/I3
JVs3W7SRCxd7K6eBIZzVTFCyc/Jj5nxTwv9LA5hiB5UDcY1hLMqiVK0MvCYQMmXa
DCQBZB49/xI2mtA1ta/rX0XtBjZPuHzvr/6Z7U5dBbx3/+5tMErg6nHYUs8lpJN2
DHOPzRABeSdmyQXs0NRCL0rtpXFwSyon5nEPiyuS7FWKVWnoYZZQv2Mf40clvUPB
N+QkJoaYpshVsUcTF2NigTgncKUgr9H7VExfHXKvNnDZ0t4TsIRKSFIt044jaSMU
HnYC03osgrPM0jLzjHyFm8wZM/eXmiW+/bZMXz7zi7BQw+cSt1g3IbQ+VjCS6XMk
JnYpR+aorx7ddcIvhgyTyDA/78zH93DdF8+xx+EWSHI3NwKNvSG0L/xZJcCNfmiI
YuTq4oNX3l/0NHCTgz58EsDqjJX96jenWLWHDklhpJ6JassJLvUiwh9+VdL65JxO
jJMXqCEVZ9iqbQdu3ndi1VJtKmNLdWK/giG7RBbaahDWX/flTxpDmMjNT2W4+TZF
hFN5NCSN4txjzWR8IyVMgIjADs9j0Bskz//2wWPhnzOaXiYGD1jA2bZFMqYKeopQ
Rie9CNel+AYWXy1qx8MdkoQo2gp+DCDBW2nPmP0Gjsbckwonin6yPGQvQmvozTMp
1JUYciPSpw/kkbmK5SSxoy3p9SsS3DfNLmOu44cP28CoBscL3zJewekUU68PmXkr
cuwGxQQHUGdXp4scAWt5qWwEETOaDfY7lQHjMSeWudNXkjSVy9IFwrCwCwKuWQV1
qJEffhZ5VLxC+TpRvTtn37YglBnzPYbrqD4cWOKL12NmAi6DfdpqYEc8ndaUf+/Z
W9s1RzSmhGPy/uYefXZM+nNM40Z4cxHiUGQI7HmXacW/EG+vX00K/GK2aeU7MVcY
7vUWArIgShTBgxUYlDFcGqPzs0BfhAhIN5gpFRmmtBTAiZxqsAMRBz/zYLo7W6in
e5igy49VVcDFZizZa4LYJLRbjFtXV9Fc9uXFZV9SN2B3PqgVNokjMiuVs6zG3JwL
E/4t9/0dz50EsOsvfqefuqB1LJjytzDSNjJcdv1AOINPiooR4SYoKptRQKztJCPP
6qKvk/gu5kqHve41tfam4CA/8w1VP+b1ggLLVycT6CooG+OfD91YNySi3bFQNIo5
mdnynlQvw9xK4g9HGys+jovODmsR8rNkUgYUBJtj+eNq0/lksHUkH09FTVqcCQrP
hnuazDiklxrXpHaktTTlQA12IAnr2X9dAi4zOv31AadDCyZFS85fAIf9FeZUfSp6
QXvYL91GpAkZ19EXkflXmaSyBPE66JxPChbzkhWGAvHlSKc6JfFh2kU4qFTA6aoy
riSq0qzKCyoqU2sqA+9e/Gyvju3nPS7dNVYod2SfQJlk7hHVwgdSyHyznNIiDFyy
jTO0uJpWg9QBAylwBqJA14GUutT/dMi7aRfjVXPMTCl0PYMfFsLtIZtCDnwXWBhv
GF0HkNQT6xNGLkGXLQNgxhWWJ2mrj/xtzPW62YpBjaFarbR4bP35kLqJ5XUiKz2B
Vf0N9qGADm1zsWhe8EzBW3vd6JX3JOHCw4dbFbXAKcitFSsqwPeNu8CIoujLq6j9
Vyqn12L7lZF1cKywi2cV4HpWTAJKcuvx/qtjWK3UVsS5F2aQLy2M+eMaRZGqgFtA
UNqdodiLDqzRfiLA1nRB86Y0SbcFOzBcDZF6WhMq4PS9m+qYmba9YeBq60caXqE1
5alTh8o5pPDM2FwQaQKAO7YlHjIT/PjYVOyMrOYR2zQJfiE7sPdSQESr3/jOBKbX
YS1IzYtkqaK1qI228T3hgEjwAkOUI8GJXqJTdFfxi1dWE3yM5LQvn/CB/tC9aEZa
dJjA1sirWTOPtwGbXHfEC0VDKImLLzNDIYEColcDfmsOOYJXrVfnVWFbN+9skJel
lOMu2txV2EcUuFWL+PqLPulT33KrVizZ6uzSY54A2fTDM/mrIZTIlr3IZvQjCOXU
Z2WjJHhoQWNKGlMwdhC0Ad4Dg/QBDlIDsv/sf2eTLg5bOLRzi7M86kRNAQ5R3368
AnbOKkGQ5tJZYnkqbrtZcaGgcduC+FVolAD3PQHVg6e+uQ0IwKQ9+MexVNe9NGYM
JHFbZjHt1PlZ5c7tHlR78m/aozLmR0AXvib368nnEq3cJaLn6Uj6v33X3AKZbyqQ
OXpkWOi9fGW/jlPMVQCSXd8Eu1g2nuNBHC2x3hqdKFo9CBNjBTasSiGyOfok6kdO
RkhALLnQsw3DdsB4PYxEH8QK5e7JHwhui7CDB7A9F1ujt/CaLGmJdW/odZVoSoHV
oF89C/c1bHugMdO+iCVIAqEewaK65T4NDkrJF8v7lN41M0Y+Sn1o4HKseWwTnKFQ
jm36Rzg7Fy5YWAnkHg5q2i44K59XY+BTVy70x55KOax25RDJGZNkiImWl0RDQ5ue
mwy22K3cs+EwUHBuiZ7jQz1sfQhkhcc/S0d4uJt9eEEyd8FLsSjxHJh5xE/89NUB
LP2vwNK4pUpQSEFz6KGecB8qiSCMATfdgFqY8iC4yluyPDmHuyH4PGeLhb4BD6db
+dKetVspTD+FYw8ib8XNbSnVnof2uJV286kJbGnM+eJ7m+TAXZnP6z1vSDJrhTJ0
eyDdZdQmFZKOkW8lh76DRibtwTJUF76O33mzyGFVw11YVqPuMH2GgWuvysecatoQ
arbEesdqqnrj9CND9+rkqmGzUs6cVO/SY4Vj9O/UQLUz4hfr12MGvlWHySs/Hbhq
LbKGxf5PQZ/HwmsFI79tqN0twPyQvyKDkIbx+pgqESpuHqk1pGimeMkNBhvB1xrP
85x5jrozG1YnNRrYhdWzCTdav6AJ7sgwvrWl0u9PqD3bfyjV7tmbfU4kcSeYrTOz
2+tT9QCFLCw/qgPatPPQqIgIaUHilmu/Efyjt9gHSBlKUPedUXbWbOUuIU1n8iiU
rmoXHMQ0xafNA5QvzZylC2gYUtp9lyrfZzWZ1HO4lNVPpH6t20u8s+7RGKo5qKVK
fzE7zCifGzHd4cZDdfmltZ6e6B4MQrWavOlK9NNpwFNIT7oVcLn9c+D3BBRhklKH
QXXeB6L/2xEywbz/qn0AzV2f7MsyqUx6Gb1lO7vNXh51KdcK4a1l3YvBHLT31JlA
/OgxMx+3jPOsal4osODoGhKIydLmOsNZEArLoA6954Zp+nEBj6g5TRsstzIF/+nj
kigGv3+vlWDMSzOO5+aEDR0lTT5+e3yQxAzEicUiKil9BBohAT0nUgggDA7U5mav
gedXHv/EXyejJc7mfGqV1lIVrEibjuTwiW8lHbCsMaXWpIB1B1KMLIRlL2TgegDm
64D2+DztNZVYMKOUBj5b5RWcvd+5w7TYarNxVzeCNH2tnvDLzOiqJIFImfiQhTkR
cBtem07JnD2074nYSDQTrVqpbikUhRJCq1DdJJJ8MWKJwVuDs0OUdjzTgAurCGkl
JrHMTSY2fiP4cDUSQsLdToh/dFMoJ8fQloOUpfiEl/3DRX/Z3HGiQZdtDixF9wo7
NY8EFc7+IBNLaRqs6z6qFw9MJGEQQ+itdcCNvDgG5OX+tnZq9xSYkTr531jRMARZ
N4yganIpR8NLhvqbPbiBwvbVPVGAbDqoH6HhwgMcjsN8JZ79jac2GAz1qSZzsg+T
/H5+67KKULLzMMXjwCBIw7UShoM8LACk9awsREJyNR4LriIDlIcUILWk90cseDN/
XMBTnzGTRd9cRcbWo0E7aJrIC6As1aq9MlHT/3+iN6pbt/uIQfvneCk4IOYt3Ybc
byL9o3j9J4woRi0sHeqOjxN9gUun7QryxaHfPBt+AFXqELzs7Jml+TFNu3v/Khwb
Do3AEx5Fp19nupnfFPqXxzxBXCSrMn4NFQXd6CX5cgLJdfUZEdzOJn1XSnicVCZz
c5S5pDda9Xw3akmyFjU1nhQxbaPkd8BG66QACvWUvQ8a6Sc4MuWGiAfbttc0jfNX
ZITbXgZurPZa83t5CBfmOs4i3ZkRbLmc9wr791nnfosq3Kb3/vSq4wpvqL6xzAvf
/Mo2hprOMrkwt0VLh+HWNoWjqirE5eVTckANck5ANa7KxUrGl7t/AhWXV943aDSy
rE+7YWDA5gmb8d8HCbRiQQNf7xaSYVN0F/Nq3RcxCPo=
`pragma protect end_protected
