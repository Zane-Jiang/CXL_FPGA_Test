// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EySu34sGg2hn2CwqCeWRzBQ5PPHTjyqTAdC+9lgIUGEpZRTKngLCFOkws607
NEahrBxWLFd4hIAAlswxPX4FLw9s8bbNQR1ET17BTi69TLFOIy7xo8v9L67s
Zni77kL45OqY26QcrnDzUEVX618NadkGV1aPxbtO6I3WDry5VF7nGRR1AZV5
ZQdyRamVbuOZ9G+TsSQJqT5fUaaXF4CWawD6qC3KuXlfCfJlHBsfAnlqCUdO
QrNkyqIvVEz3OZRoCxggRfha/014ltz7RsiHATm1m2ui5stJkUJn/E4ssTpB
YwDP+PHPDK7UcqPFMsRrKeuuRFP4B+r4onMegjSVGg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LFFi4uOqPR+muU7hF4ByA0hkf+EAdV4W2/iENCiyoDNRl/otvZC9vTNZS5XV
wMWTdoaeU9fsFe6SwNhFvgjETd2OS46wlgVkQoceZJMn0yh5Le5/2hnQYfx2
xzmoo0ymMNVF5Ud2CdyRvmyR5d+WhgvO1YwAYBvgHPbRZ0JsXgLqy33Hqw+y
Uhsxbrs/pEqasdLJZhF1Tejkmfv7RMOrjtMz0pTAcelkak/Qbaxwk7Fy32Ly
l/XX/WgMULK4SZItHLRVzyWFpn/BxTLl3QLRDDKiAJlccJVpKg0kPoeCKMQ7
XK4tIyt3jsRLzFcTUeBwi2cCJneSVjACnbWkiIs5zA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
puxNlV7mZatK50hcqHo1GE2LLbhcgT4FaJvtPsclGRM3BT+9jNs/R2yU3cQP
HwdvFqQjE4163hEiDMDnwdbWUXGuuvUUOYnwmu2QimIb5zxNxtryZRT4heME
l1YNcqwg1hCZaKfwzOwnkTyyTX+7KTxPXkzwUHlRx+ql5RQgmXQegt0+b0x0
qdtzh88uORbdK6T9nUYx3ksxlAfvAISv4qf1k6AfebJ3mZQOi+3eG1ClljSP
HN9SbZ1gGrPmRY7kFFPQlGUOH/JC7tHidwx2iinrrCJycI27vSTj1YDYozAG
YEvnSCMbm7h1TbY3alajqLNVHm4wYdKWhMm2stF1bQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
An3JsQ5MFSgOoDdtfILkp+EZUMlYDhfAC4xVrDQYQSmDmaj5CzXZhIh6Zr5z
WyTj/KxXJ/cXRsJPm3AMtpdzrNOKjEeg0+doFuyw2qlVOnK7O+eH3Ec9v1iE
dayjN51/LW0YK3sKemEubJLO9SISdkEZL25UmKpqKQuyalaZJN0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wWoBrmeT/xIGXXrgF1Ne+gk9JLxpbX5T6uH96YvYepMrCAsyO8TgOfv6guLk
I6SMHie2NMtmbp3HC5myn0Bcw6GSApsus9RtgK52IA2VDvG5Ga3zaudCZSWD
VP6aFVqgdVRxmFbEl6tQNS1M1aGXYeLtfjNude+QXSfXdUGBkE8nzrNBmdVX
Joj9FU/CDds7H0eNxI15UtuiEcFvU8zZoZgSJ7t6sHcj+TPL4QwcdMpR+0Ez
Srh3WCuHDNbsIMzz37ZfJJx2KgANb5+eHC5+SIJ7pwt2eKX/ap5caryw4VqX
ssvlQHDEBjM2foglxqfjvKqvJUxLX63HtCQWMecyJVI6d0oNTvkr0lPtLYhF
hPDgSxIy1jKU+Uaf+bOPdMrHa0enry9YGewOKANmtin2nxFIoTK6hxJFCbkY
nuloZMlVqoe/fl2fIYf25XvT8E1SCB9t/znvF0zJjIWKRsmKrqVduvmi6K7d
nlIgtRZtosZUneVqI46IsoFoKbIYMqCj


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HZLS0fSW43LU5EeeOWqbmZjXmNvYD8t7d3WvEbI3+vQFOdJsDTVclaznFRCo
oSTeL12ttewcilP8dqNSD6grvhs6kuBxFZxlJBfJ1BFwyEIrN8CKP5cKj4ol
ZwsyiksQFjmFd0YKIwtOqpfLPXEaYSFptKxek+VWUSU1vdo1qaM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kSPneQBAqw5hZS3odYjDy8YSRvW4h2BG4rpP+BFVALLcfO1YrPRz+EbqRWSb
H7O5VfWupJg9pLEQ1pUzMI16IKlRxeKSg0IxUVZVW+3OL/oooKqMOzCKqTmW
8EyFeHTloF2p4HhLCL7kh31E8cXYiLEyGvf0ttFSvEmSSH3ffdQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
hYkIt3Ppr5BHUMf1tbXzxrMRXT0Vh/21hEuu45qD+SCnSjWqxdEY4seN91aJ
ppNkH7jHMh0WojxCDmtWtwSPTHINthESjdHMqJESdVM8LUt/HxkTeG9sWs5r
paSssdYOyNorOE8sMheyUVv/6MBizh71ogIQmRVY5A4uWEsB+bi+ZSo6jboW
VHCRITRQES/DP0qRjDwLLM3r/fDJuZZ1Eam9rWzADS0fwgBvaw/yYrwq1QYs
ZoUKw7uoMQyisQ08tAGYeRXoQ6NJCbaBpYyceiKlCaAZDlRhiq64dyN9CzfY
mBE16zkqwx6dtnms4pZ6IuRzrbvormzOnx4U4u/QSYnhgsfMN/aYzK2O8Gne
v/A0pXjzS0qGga6QhgZtcp9LqA9hr69bjTxAEJ0D6TBT/993qzjxg4XyHpHz
3H4WBOg02CCC6s6K51jY0e07aD/7+k6+ydNpX3gozSUujZyOnefyrDxRrDU2
7sSHmtvhxFAVUGONu2+jA+EgQ15UcTtm4Sz1EVoK5gG0k/NUjg5Rf2ZwtN5K
71ndiQWEg91/67ZOqsgm7wR+zx4XnhTIEBlHhtMiqCTTcym0kUrppsmgoVgM
cpoIQc93jbWq1RS1tFB3wGIl0JYIfKkC8v82Ua0XmgGmhy94VUnXTkA8/8pp
EVIPgkxcg+/RMoyFD5vnXlDlBSw+5h9DzqsImnKO49mAOMranVbHfWJ9BDJM
Y5sTtCNRZpESpRdY+wy9jHDCAuwyKDHPtzf9GGwdCul4pxiBr+uFhyb9AV5I
bqpan9A/lpSlXpSrmkZUtg8qT32DFfRphi/po5PzRG21J+Ck9cauTO0jrvtd
FZkDeVcSIX098IJWer3PxSgnMMBSfTv8FUrbu+lgAdhBHKoGftCkvOyHlRBE
MtxueLf0/QtylJ09gL7xVzARdRDCq/jQAF8iBIFJcbJ8T0sE3p8CclnCofBj
ntCrN7z1xhvxzdfBNLFeTn3ahovN0+2w1/UV4TLNZ0niRbcT4P3nv/Ysd1qP
MI5uijmZsdE44JAHKV/lktChcywrThUrTR5s8rcQ9w952znXgkGtB2PIItcg
5oAUlnvc1CX2pa98ESeXDUzlBWdpzrCwLg1N0IooXYVF3fWaT+VKjcRqOwsn
xeunBzqPV+dVxWWhNc4UOW+Cjo0h5u9tRWuHAD239e8sJdvJ3vbNzExCo5BU
+Wsk1Jb1VyxEMXQ2rEDlclNhzn+6b7KV8f/17XAGUeydfFtrind/1LaRBcmz
io1X7nyjOsEfWMqYz/dFho4yuT1nFsowVOb51S9XU4SlBDWvV7uqg7N0H+ft
Ad3u9hPeB6KeZ+XnF1jZrxKPD/AtDDI5z9vEdodWssXy8g==

`pragma protect end_protected
