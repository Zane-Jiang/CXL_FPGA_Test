// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
bs7ilpCY9mJa6XtEV4uu25zDRFbzOELmzy45OWbwXOlxO0L4fX4kwBqumg2P6Ono
zQsQIjB2Lrhw6JF8U48CCXWTaIW7FfemKh7er8dg1lv+hvY5csIruLDQ3YL3vA3c
H9SnWd5JL38eaqaEJoghoVSEysLktz+h5JCiZY/Xci2RH0vTE/TLXg==
//pragma protect end_key_block
//pragma protect digest_block
J0hbM2Bua3QLEI6YUG8hN7ukvW0=
//pragma protect end_digest_block
//pragma protect data_block
yCQ4t+5FIHOAn3vqehjJF5rhGmT4Hp+Lcz/UklAqnRPDbZvtQFicTLyG/x2OjkHr
kMwEeAzJOHg/Mtbp76jMZKOYvR5tL/fJQCXWbk8OeU9kmJfrepo05s3q2Zqn8GS4
ZwdtTkHmue0H+7Hi8rI1xiDy6yY+REV2lFXlzXfpMdTjCu71diJFEv2FXtIouq6c
rPvOdpR9lKfp2j+hqWzSE7C/mj8CXQ1L4MyphGV5QkcJADVMrZGR99PfGUR1Cclz
ORy7hxBEQR3VCDvlM2/jj5wXovyzCpoLfQF0XR8Xnn5NzYInM0a9uuSxNb9sGZus
s4qxPio463u+9AWVvCKpT3+pfLtPf9hsrvtCnkHucuat5JPL1Drl+X39HZz6nArA
IOZUiux9StMqvmKdfAtj72QGXkHCqYbRlcfZ98HeAzYaLxA3RZS3tLnaH5PhkkBI
riYeiVQzBW00/+JQzkNcnIZPQtbGtQPx4QFxGcS4mDY76Mo2iWUDnkkm+AQaoqpg
MjgGxz4DISVuAUXbx37g864plT0BrP6Z6TtP/SaAhS559DrPn2cptuOwTEu1FuVi
Ibsr7aKW5x2LHjTUPFwFVjUR2wSn8T69EB1LeezA2Nr1i8CSvHCtOuZq/BoaKzKJ
8Mqe5/cvL7UitTEEMQMZlGFdm2VhaT1T58bx+2+uAWIw8OsNyeBA9SfXpXOovP1T
RpHWkwvFcm45ad5QpgpCmqNLR2MY0BmIXNd61QaqETPo877dj63qpILIDb84uQNS
YO0rYcx6myVBN6igo2ySfnWLhll5ClC23t+y9sqVaTj0eXPGkEZOC4ldn7mJrRyb
2a/pHkBHX2XQLpaIcatGhPjvN0QBSrSPBN/Lh9Xq8uNIB/56znyFVmNmcrhvUs28
XiC0zRXHMRrb8ZpxfWenJeyfVdR3e9e6L/OU3qw0sZY39VwSmAdhdmcOxd4KPo58
qNaBtyihmo7HIPV/i7NIjMLO5QU96+W/C90y0LqQR9HoXhz/BANnFlTdsXbRBB7G
P3u0YZKsA/eaXqaAj0aOQY+AJW4x6EkVWZIym69fi6s5NSFlMeN49Q6jwuvjqmgc
ONzSHZixznYZPeHNtYS3CH/rSY08KTTJyCiB8+DyLrallETVUhyocFjyHJekgelh
XwN7K8y6FXBNOUQMaqUgR6xPObFyfij+iOvS+zNcO8CdbP+uc6qgryZWQzqZoqqP
IocLDvf2ShySCdxN5YmCX2oqBNvMWaKdxJftRq3ARnLUoQcDebVo3yJjdAMLZ5za
ld4SeHneVDTOOionrvdINxhi391zgTxjijjmKNuwPX7gnHfuL5PibV1R2lPxzIYl
76ujOSwXLDGsnblpXwlTL6zjh3lTbqE3QvRtM68oRR5htMZ/sN2nx4DK02ucy8Pk
gvl9jY1T2VF/3PXL7FNPjWnCbtCFQwtqkq9MRLz7UQH3aHEaV2UIf44fWbkY5VDS
yKHkxpJCXaGqirozE5qBh1qA8Qg+M4+HSPInW5jvQ3+RUH/dlKR8Vdn+Zvv3wQnl
zaPT4eykv41ZuwBgaJQyGUKu/SHd19dGOTBRv4AXNfgG2YTZYTvzMXRaoM2Ncolw
CDpPI/kHyiDR7rfV/oNR297tWYb+6senF6JEg7dOwGFXLeakpRGOm2hEPBtLbUoI
tVuoPZYCOEnTu7vzRTCraJ6R77xpSAmAQ/7jEpu3dvmjEc/jTiMKLkBI70IA/zvz
06V7qH0ZX89FH/4YOpKhFO8BRAo/EU97++7KjdZRASw8fW6Ju3rfC4DjLB86Y8xZ
Z3H4tcR4c9BFtE2riYgSGv6ZF4I/o1XSTfuPFxqlGPOX/Ox90+xOuaV0o4tifQTY
jyjhb+NvIpXuYe+SwK8/E1/wl3ybF8JZVilyLa92mh0b1Hhl6f48kiSs5LoSNN4s
1OwXVrRKTDnjJt4rWN4OL+KwgLEkVUVYvTQ5ehbNxzFJ511m3YROZTG2sVDWNYP2
UNxTL0DsMQtHUgGoW8078nnPb4pFonw5+eF7VGRfIzWpukUuLFPfM8DWW/bV+Uqt
ngL/+zltC7/DZf8WrF+01+5X2q5p685tlSwSgSd9Ni/qZUsVlrQkdKXf8uWxDIqC
Khs11OXzLqzBy6B1U06Q7p9Pw8awIhdYWMaNrGAeCILdO7ts7uaSRZ//nfmrtoZ6
KQ+5SJLNY1QneJnvZixK/cL/kv1ZaBEUsKEJUXMkl6iZo/juj24Xfu/E7/uxNjxP
8UWJnsqeUEAI39q96HHeZmY/X16Yv4xD0M9FX/633uu47gdFPr7lxLraUHkh9aXZ
BYJXKIhhhXc4b1lSMELrRyU8ADlYy1e2x0waiumk2RPet24pRnb8AW/z4Ui31QA7
iVjXI5bAIfI/SoFxvnuEbgKkrkDBC/MwTevvHP0PJBdH+f8ymJdeg4zehd5oRRsN
UM4uYAEF4MeIxttcLN3ujnumgMmNcNjpcVkJVYIhwsnX61xTkIHREuYYdvMsavpe
siuBf6NhY2FtHibMD70G1/kIcVJo+tHVeKz2NVbOCdq7rViW99QvOyf5fjhm25pE
+zxzkpq1+klMcxgxOpkvwaiWVyi9F3ssej2tyK/tfZ1rA292PYXrtovi3OoX+0zn
H/paBOpwjLkf6eKy/4dMKi/BeCughYUQcDLuh/Lw8eNG+qnmkMOyia8eB1jiZZXE
6Rj2PXqthhFTXHufMV7HUtKd4RDv7UaOXrmPKXPIoAXTLsj2XJS+0vcvEoXdNBJD
R2VpHAerJC7nDYrGCkChUR4Q/OPgEl9YMOIdQjqxXmSxpejov9kaRzyYxEJmBzcN
4IFNkJi+qHxdH7dV5QKJTKW0ZrQJgViiAAGFkaru/IO0vfuiNWprIu+qfKqiPKmr
uuqLYJUNq7MUWmqYujn4hTY39KLSIz+sVPe8tTmc6QpRlG+vanajRNwtn/GDUmE8
tDaKDcqoQDBgx64hO1xnpyWAMH7BFiWr20xVLwPoOSPECvjGc9UUX7g/huE5isyv
9OqafR9hQSczNjDJklSHPBzo5YM0HobutqFuePUf6G/z9yKYPlLLRcU+iapPn09M
mU9iQzVKpMhrjloVLb0Kias/GnsLC+plxv4a0+uNu6CA11NJIX6TA43/esyvTnI0
Ce7r3anAWyI3tMjFgXCYSMe8cqylJjkZWU2dwU0OjRnfwBjgxw4MykwR6xNpuJvr
zF8cCGxxQ4ySt6JsVA/gSP8QNjnp7Da0How84mRXJPqFhCD8AVTgY5hrOErjbVfE
SX1YKXPRqMRC3JLOOLXX0QbjAtpYk5xqAWW1Eli2b3xiqZYCFRQDOIvheVC3AXOZ
UZVHGOBe+snYnTjQU8c9J+1l0yKQYiyl9bbo9sPge40OEjWDWX83zXoeaQFPTY37
qxU4bOTJHYmGEbe6ZWMKLpStkDSXo6t4xFqZBIEmsoR2/N9vSuyIdYJH2aGn4soS
rQoDFYOWj7m/7xLSp9HyK+Rznrg35eLgT/NDfFaSrF6Uh83OX4WbNZeL9S3CbQ/T
RE9Jpct0fbU3/RhDuRg4m/6PqaAQF2goI248HP4NJKsAbSiK5NmRaxDM//e+krDc
O5DohNZLxET+P4fwdGCd7MbBVmVaupKurh1qHeP3Jfjuuu7yqRWSFagdWXopdb0r
bsEqX+tEr4vOA7ZsCq+CXPYuMDTVnkJZfp0fqOYSLUhYfAzUJM9QANXIHsdy7Acm
9QZZl2R70V6cV6i5rQUyqfatmGkCbjml9R8HwwNOoMLIT77Gjf9wDJ62M+p8jhQe
GQF6AWsd9wr/Dfgi0Rf/1Bykd3LIXzUkMORPujScJbQnWCZXxedSTkLg9jvH88v1
Z+YbhzHxEzi8w7tX6AK8gEAEf9y/QhOV1vllj6csxSUvN5d6YZY4hY2yD259dMmN
+M9WTkG7qPKDT2SFbAkvZYkAH7VIFkTn21FH/M/k2Q3In0f6nDIBLnqmdcgNE7OI
0rboHsqJnPeqLRAy02rSXntj2/nzvjOHqlK93s9+gw77ejLPyZP9DOjioBWQOO+Q
R0C0up9/VzsjWnVrjeIdb8HeguUvq3TJolBQEgfQwcxtybbWqHquiy+B7vjiy23J
RNuKaaL+Wyun7jKaPwDWsYXyKagi5Cbkimb8iyqIGz1XqE5al7XqVUUWfhVfpQHe
dvggtkIeL36mYP+TRQSxUt2tAjcyT2eKGumA2nfwVlCwF6YbIz1swo4Q67waYew+
mbw2Bm4JX6c02EFdBsGsMY6TmEWorKZh81wnyRo091BvNfUteAWnD/J6YEJW5Y3V
73nzuBgHAUwy5DiG6vg/Ezabj4rqTuTCTDmFJZuAISrsIZ2ue0RnYGgQ7UryYsI6
qMQT8PYw6bloAub1N/exo935Avna5kDM8xQuD5Aqehd20Zqy5oBJ/+XKBe6T3ROD
N5hGfRNFICJEH/euFPHopIKkI+C3TGIwNk5TS7mPuZ84R/8G5icQfSfINROVdKxo
eAJzuLwK1x4HWrGZkzbiezxClT3gaRyd6hZuDiOBFTzhwRChrcuLfP5uHPVIRK2+
XWs1wiHjGvLE4Pf8guqnt+ak3JA6yXb1pG0iDxSsRzMIBDsFsgu30T2l5HYl8ZOt
QdJCsn2u0NWzkjq6rnZD4rVQJYB/yAJ7Zzey4QesSr+coXt5FVsqj5d2pG73wXDe
KawUqaqmX0I2A+tI1X/DUJ90dPtkpThEk+g5Ic5Bfd+UNKJk5xJeCgcApvVf7YTW
58bS+AHB3iujRBdJ9itYjaUjQkkLGUVo5vCVdC3nB+vn43G6Grk9//0UlgpOA6lp
oaUkJbWPz1luqTAzzRfbAQLgc7ryyjqHBdo05EUoCW5DlD/mmMYOwlUNaK5hqjZH
TkFQU7OvZ0imS9lHfd/QQigrUcomCrLLzgk30XoMSbyGwyKZSH4WTw3gBO7bzmK4
UDW/ulWIg5JqO77tZSP3BrNArtrCoO3eZiCUzHtw4hEuiSCYj5gdpIW0FHMLrnGl
h2rM4J0kZPjBYs4HF1j5TbnAZbuD4M8bDrC9q/qZg0rX5L1wnFFuL14kgetJnEAL
p8oRzTjHbd9V2jaBxzX/H2DwVcDEEyAiIgRaIlFq6C2Ue3tFDmYfMQsf7gX4qh7Q
wHDrHASXnucbtIP6RW01/2Mwm7TblYXCKCYUQUFGx6RRkylBLSHqm/f2mj3h3j72
3W/BpQKRHef62kiBZ6zL90hB02Quf5PImqNxjnbRX2TTXwx+Nu5N1gIepzH3A+gn
6KAzBSarQGv1r8ynQAocl7F32G+S5WpNyldM68TALppaSlwcVcfF8gJGyQ+Zx7We
AoWU70B+6quUayAmnlDXYAKFW4TAdLufJI8X6VL1PPm0942saKsf4iQ0b6paGu/G
L8W3HhUh/KdA+EeAwiHwkzcnQEpcB9Pb76NZFiz2HCENSUM8xIo3UV7gCfmDrD+m
n12uL0bRFNHuvPLJT1zYbnyaZ5kgWU1t/mXtbWHn0g3HYSeVfxdsrNbm1NMZWVbl
uBXkMSefM0DFEPvFUEvYMkwMHQUPP2AzyPKCWte30qFIUyTXQUt0qrWeeXnUmQ9m
YcE9WDNyiBhksUzYSaFjJJoti91iGBkj4/kk49clB+LWuwSpr+ICi8TDq3Qdd8f3
IfP2dJAays22xGGgoGJVK9x1Hvgp8hzF8xs7DN6B3Y2XxPt3Z/IxPruwX+K/ZUKD
9KbteZo27ebX7rTUo3OJFrNo2Z/K1oIefzq5VFJE8DCYcpYcNFBIRJSfoZhgRPQy
XoSTnNW6z5fL2MOZj6ipXAeYtoetO+aRBemdpD+uPgjXw7n2ycpgzuZw/nbLUBQI
/uG+ByPG1g6zax3jS2Jbj87GGnVve+6RcznHjQHLrNJgI3YtFzhzMQQ0iGCe3NUP
bLbm5XiGXUgzsnew8PRGPREe/WyY75e+aYm6kgm9eyTTXfkhVyYPe9FV+MN4rfuM
M4r/5NDm8bcblfvqwMw7zcChT8/R9SzhPuckI3OkvJAv6TkFfgMGOJyiMIZAhTLF
9ul/i16c0gvxsA+43OQP/dioOLZeSvXHpVYg04/7BawlWZUItBV+WTPF/JpV/yoM
zy0ZqBDzQQLWocopqwP5xoYkvUcpjMX6qItDuT0h6vz1f9GaYFXb2D+1XUCIEGGV
VxXuVV0ANA/mxwZ72Rb8HDz31I+QXzkUg+Sbq3mj7yAyYj05no/nuBjyHRj/U1zC
hySXQXSQg5PoAbm76w9Fc+VLYhRuw0o659nBCgCEhbBk5nsWvmrrAwtLd2wagwrD
SqHZhGJxtsshRgpRb3eqfa+ALT2FJWOU5UMbLAhdVRnA0EGh2KXu61yWpcGVFXCf
BkybBfG7QyrLF3zdSIDZ4myq5UhNDLLMIpEXyrX5V9PsGG+0tIOBmvexNbvX9NYc
Ef7x7fWnNyf/Zysshq0bXwoJKdb0BFXK+PHPpmnGFRfJlN4Bhp96Pz+LvmzWae2a
WvFFVHULGxm0ngdr2HuzWGCHVGI5QYhZhvkEUA7Ffta5Q5oFZfbCI+PyQfbXrmCd
mEYarR6qQx4GHRjsl+QjrmF+PwJwRCjZFvza0U8LpynO0tADJOvnfSI+ZE+dxe8k
tm/YaazJFNehQgQ+mIJfxDJxkKoK7FgjZXmPcz954752b7LqppTtbbkudzIFUZvi
naPMDE1ypCiynCyQYOIVdg4mpd1T5hhbDKgGT5GvL6R2yKB7I00u80gMkH7wCKaX
qzYIMPoq3WLVuE9F6grgfPsTNFPp6d1svDmbJ13GDAyvDuilY6K+VcNALBDxCEsc
/ZwaeznOB67G1kQGd45dasY3OLKAMMTTH0wRqLliAwcTKkYNX3G8ZP6J2Ng+UOUZ
g22+2wKhKzX5qTIZlLv1CiUxPtBvynIPJo/Jol7K0Ks89UHG4hA3kigreDhcv+2/
TAmz/7FIQntBFp3Y2DtOqk6LTDERghi9Oj/a2LSVvwIiu4FrQOJz+0qeXjK5FFFz
M6YSTewzL46dvxzDVDTYuaqFghtlwDnpenaR8r1Jlz0jgCdc4BW+lw9SJkdp977t
I17NINp2E+HQKCGqGtGEIyhtfc177QP8UOCKO8+71Z85aUXnZHBcu0VTCDwQ5K/g
4wd1Z1JAA5IBG2IrHEnC0kD+vcOU3WgG9kuylCALuNeaxIJ9/9L/AYiiMB3t3X9o
AxfZ+jXzoJKELM5m9a9VFj9JLCFbygeiQzrz/ZqOLsCqMvSFYxxb8LN5VEU5qj2g
JWbv/ZVCK1k6xkMLO8tuKytKeCcwW+ubBKJLM+h+T1goALiBDTQE7WjMLnnPTMgY
VW0pRqEfe4V5h1qqp6toQXCiz8cvhOEWK4ubAsMIg9ONR3fJIUKc9jD5dIeBTfoV
E4LRsHjhh1wdMW11C04bvw+7L5/BiplTm9qhjcqZJQWvwK5VIIf23ckcKRGNVsAL
q6f0Tvnn5mq7YyIcs4FtEAUA/eyusswf8R2MB4nej+pjT/eoeTOuUQMqUnzy6EHv
KezDQ7A8AbcbykE9DDaUNopKu7QiHQM3XUmPHzKbLQ1ZSv/K/Hx4pnqETU7HZGSe
iu7a4bWGUJENDwBNcsSW2ZNMGftes/LM0GTe3ZYex/UhSPM+ZYmvW/+QmaWfi7V0
/Uqx4xKoiUc4cGOgK3EfJTYSx5/rfle9k15QLLFKI4HcY6OqnPKOuuueBy/iIb3i
hldQT8QygIUcwChQqnHdqDJKMeM0LO+S2BgWT0CGY36LyhVLDIwZXC1oyISx435r
wan+gQe2On4DC4aF11Gpbwl2CWiQdV5KGLFqvG4ahqK6JuAfUbuKY8zfFrnA+pEU
AuMhwHS9d7G87dKa66BtkPUPFcym8nynfGQHLWKxA0vnU/MmYeo80PqSFMWxhL8X
aZ97xBLe/UgplsmBa1C7c/fvaiZBnjTqSIirUIAJzqWoTqJqlxWEE53SV/hryy/9
P0A82DUpxlqWcsusKw0oF7yr91oywh+PN/qnRhLOeZ9s6s1LfgTQyTpcaqmHmXul
t0lYk5FPwVHWRhYmkydWGSx5/iG0zVzejjr/bIR/VE35rRCmDamMbJEixOTqJo2N
KNrL/ZNanMXFRmNjC/x+SDvRe1PYMNdXMqo4JJHZTpvD8c+tHFG2Qbjq+nxcrl3J
PXo7NmSCBWGJuwi1YYI/N8i2A2T8utjyi6ciOdjURLortDOrugw57WtlquUzgm5p
AyV4w9O7dGWcjZh4+wOBOrqD9iWcrvuEmTFeSF4AjJhgTXciTbeHX0z1/0sOfjWr
+78Kw+susDvgRUkynGQHu0uaVu2UrV35qznKMBi+rJjiiOcTPXFJve638fe6iCl9
S3KuuqiA9ARXTSXvF3XsvM0uATNCZv3AYdWfYrXoUWMMXBp5UsfICcaha7xGMSkI
T4wK7xIA0u3M6hurAzPodt4qaVPQJIcUA0kZVT5WZ1DDBeP0JlEYtegXnb2o5dyF
zVeWFxdWAPvr5HyRR+Lf19mIAsZEEKPbA/zR/NXhxLS9p0Hl7gYhSxZMXLLFIiNm
IskLFYv927q+jOavFVRLp6h+rUAO0pFWY+yRrdg49AHlzExXsIfm1fJxc1DmGFwo
kYsuWZTaWjtSV53PYGJRjjgi9qznl3O67YpIKzQuwOCkaewYmHEQdZ3qbQvo4SV4
pLTl7Zwe/77ERUvS9asTM04JSNcZ2VoxeYYK2Xa7mD/v2GhmpGHs4EjK5psSwnU+
fsGTGCTHZfn9NlrJ9jt9w4kOogqCxBJDr35iNe3sIyLnIlgtIIgFopYJAuMUI8gI
O2jnZnVYt7YBAy31kak5zmBNBronFWCaJFR0zchIeUf+u8A3SCRxVE6da7z7uGET
/MSLk8PsIkHmv/1A1pCD747bHzogxY5i44fUDGu8FrLK25d3ABvx13vZ6kbXL0lZ
Ppnpl6wkF2ylu5Q+VGUhAGBbnUpG48gdLBn2n+Blt9ZYs2LZwB67/PJl3iIcBOok
hVEb6LgPnu9ikGzw9O38bsgquAu1Nt6aXEziYAlX4CRPthjA2j4tAKChHlfliFO+
+rltSvYbF9lNeRICla0sqTuIzH9VKucxHlraJzpQt1TxAW/SLMT2crta+B0Lq619
CjW/bNW2VRxiCB2GSMJ76Dn1YVUIFHRmGGad54weDHm+SnvZWbhblAHR+2chzojJ
I6OFA6/i9Z32sr8BMmYDZgzQcxRYpVJmzn1Dtje2wDAchiyDn1Rd+us0qRVoJcOT
6AELrGPoBmEa+jn4DzAOvU03z3X8LG73+yuazU36brZMxbPEvsI6PqEcxKLyjmMa
v1BvxB2n+4nWADhEHVmljnT174c4/MJjjVb2KO6qdr+YNVpm4M5eiNyF0dUAE09h
10OKTecDv8d+uAp5gEQZ3+8T+SjRVdrpKKXc7Ul3oCEfgHwjm+aRKDHnQQ7UN2qA
oCquL/mlwNTbJr8UnVMnlD41zgMOI1lJCenTGijc7tOa0Adqhclm33ph/p2A08oZ
cUKqqDjwII/BzlEm4l+i1l9aVHSgzPju9S6E1xQ96QuNCD+PAmi/mj3EeMk+Pahc
sxj8DHk3r/nHVaqzKC1cBOOwbwgE8jo7T6nTY+AmkWpl8MixzQs2brb1gHLSbNUx
bUTz3eWDBAPpQ+O0D/Kb+F3SHfHBm/PgOUTUiOfz1xds90o49D57AoGrFbipkTEw
Ak90taELMSg6XnP8N0jvd8MsqezsaNxPet8b/08+lqHQSRB759bhD8PvB0mgiFdc
jhGjuzRIOk2Amsrfw4Wj7sIfcWMgPV4RbhQ4Q2O7NFfMv4z13ZchOWHxRZIwp0Wm
N5wP+Qegm4PZFG7mnC/wf5/c5iYDr9kfxGu7Is2Ibi+aRrZV0u8rt1WTjefNo2rS
ERHVaPdOd2HkMbY5XqsAppLl/z7YlCE3bQe2iVz1XapYcKxpMsIAM/lpKr1MDou8
HbLUCfKA6Yq9GuwIGzhIO49CnvWdu/PybJep8vc0ixSgHrR21R/u3HtAhyRdpxG6
Q4+o8iQjBeNGBFJECV0+NRYjVsfuP311SzxcyYW+TB6QAcOSeFtt/S9c1CSGQabQ
VF89/aJzMBG5I0PbY/jM2RnzsYpeZtIa8nWcfe5YXkiCfZtiNLnRDWHZz5FLfB4T
/XJ9H5XpA6IIRvKy0eFL53DCbfJYu0glEkkq1FhzPN4b69Gz0ourhB7WPEygDx0Y
293yY1AEWSVIeCXNmVoHE1o+vCUFEbwzSnEX6iXG15hN5vbF8IpwiiGA5D4kv4Nn
GRIkpsiFIcPh4T+pnNVePP/r1Wgw+GTRtcM5pEFTD9deJcvsA9SlSIGQCzgxhvJ0
tBmOWk8N6Xj06+XPA88JPQn09mhXBwYE27ojxJE+T4YpVXWeuRFlHbKkczWR96u8
FAccR4J8A501ElTkUe+X3mTjUzWV7W4n/BdMTG+66/BiM1kD7S71nY5KwC7XD4zW
I+XaV0KJ5uTQtdGMitXZHGivpoDNWuA+7NOULK4wnb4KYLfsyD2p6W2PKr5nftnp
Uac2VJSypYXuwsJnckPZhp74i6K8ECBKcmeBKNywP2GMcmXDt5P4FpBKZ/Ya02LT
kqSuRBOkaL3MQ9DvQofXP0lg7boP5ERTajcqvazrvI0F6xwjE/74h5w33+DA61GZ
QlztCKS1+kR/GtvNNcpY6xdbmqlqoVinbkvYQ/tbdiwsi3Ak4yGpBvr3Yx86azXw
/Owj8INjTLUVyzC+yl0NrYSD7fL4vV7X2x6XJDk+MGCDub8MB7hsz2hInZf05u87
dPiDjrUdwvoPt5QsOooNazV8591En/GyUAttCgcqO5okItCP4ENyrlkROfy3QB84
WcsRxVXpXay3EvCVKwJVbIEZxZ4ySv9Q1NZiPqzIiGtXteVXheIVxXRkFhatKekU
WVjefs1KJheLZOQVM8wteFKTGT8kyPSwZfUsi42gQuGAsdOykqTCWePsqxYleXmo
KbGaTle7BxQB8+usvUSiFacy8cGH2hbBqqEuj7pfT1WfWG3Io5prTF2T7MzKzLKM
nmqO2sMIcyEKavGeK66CbJanEKf1NcBOTKHVQiGbQX6G3fZzIVJbTNWPAQTC8AKp
8HESL9XSpk4ZKH8f9GlSthbMVXMhUil0HqK/xV2Xc+9u1nFP/triviOobt950IiT
Tk9ifApvAdo190dHESJTrYSGEHE+JNlHMB57R81UOjUyD6M6rpSHtNqTUA5nceZU
6KXyqXAZveEZXl9rMaKcS25M3dJSXhTPBC1JXQDZaBUjmMNt08uwj0j6IjyHW0iE
xwET5a4aUDyfaNrkGmPO4MOfJYu53SIVluoqVVj6JLh2t2GDtlIFUrxrQoaylZbg
7cDCFbI5SIZ/XbRacOIvgA5yDbC6lDUZVHzZjMqb4IOt6gtG62BAAj25AV79QRn8
wU0NkBYuolJhSELukNMdiznk3VDaB2ZiEW2vGI5f45A7LxtEAYGmPvIqkddg+4GU
+6RpqnLknhjS8hFU+xI/YfKstYM3fXhfQIEvBio8S8IBzCa/Vp1UEqLx891retNK
hjhYu4Semgon6/rIryS1vsJ+MHspOJf1GNm7cgwwrXqvAeofvF5NGl8RZd3v53E+
PTXLi4jh40hAHASKAirzDosbI+QUxkvk5jQ95TsDzg+nONlroS5HDqpv72bCUxVv
vzWCJ13QBmLWWd61QECDnnFK57JU/G/5MJBHl0XfrpRz6sJFYoRyLb1EXCybBxOG
DflqZtcDVrrKkiFxCNIXvN/uJrakf6vyMW7b931clt8ciYCob7mmqQXm4g+C25HV
YsnYfvsYUNbMksjw89uJx3bzEtkUJydx+RctwxYTlIXfPzYlVmeXXxEM3wJ7xVpl
5F9zABjEaGzeSEW0vOjrbOG30J1cuQ+9HcpBHxHYvGWgLnw1vm2R4Fib4+1Ag0Pz
GvswQj7Nt8UaQ9Zrgv6mZvCUVd/8VztfxIPi6rpSQWtJgrkiLkpm5gUZmfC5vb08
GOpkZe/KFVzLamxxajBCOA9/EQXODMHXLCr+fdNR8Dxep3jyWbxJzeaAEq+qVafv
lNwFO57yBmVT4AjG0cqLP8QRvRqoXKNFxk3A/gXed/ci30Yu6zHxXPw+N9UngKIB
VjBHN5oiInNIVCzKVl7y0cxl0QgPUdy5tljJQ5Bi9uxrMTLoKmo4VOKIbQpNcM0P
XwXNYix6+nijp60jh4anPs2fmupZHBo2uFTTkBZn608QfIltFfapJ2VWA+9e6hiE
wQf2Idz7WxpXa1eRYjZ0q+jjPW7UrYDoAcBE2OKYq2CYDFciR+xF8BGq7aXYOwbg
raOu7PgfsosC1wPlxunMGBoEB06WBuq8OUyblZod8LBeV+k6WAijes4Q4r+pI9F5
VHjUPRftmgHvNFFowCJu4G3nS0a8wNQB2cTxAFz42DCC1Ld5uiFm+V100cZ6rdse
Z3kR9uYz7XwDBham9TFN1NJEIC3VOqWJfolvzp1N1hWPa/HknDT/mA+y8NBlXGjG
AmgIOun6yjmD0+8w65FVaQG4vAxgfBVAy2wKASPIUmQ946+jvs0XhwBTcGXdT9Fn
vfztF2I33xvmhVH2xVBw9d8Ea9HiMrisL77/pmS/5xImWjmMfqGO8yx3MuCIRiaK
1rZQ6yRjP1B5jT5+gh95j6QEy9ipCWxK9EMhhp1Ad6cu+tUpMV9yDVcpDHRTQ/hc
eDVhG9TEqSKuKQa+OskzrZdkyktGp8BzQ92wfG4soJHjcSOoOrW4aEtLMneDwOxa
q61nSHnOUu6PdCA5SyOMFM4HbuBEX4fIxGHcYXbVv5qO8cxOAt6fOJPCLVpzuxr7
tPzuEh6bBY6wb7TEpVoUg+yn2LiTffkxMewRzf4sOsAqaZEx/tTajlDSd0XUtLBa
b6NSTBl6zolMcpHsAICWME8M1ZGamvIk1iV0pMpGwmiGzCIzmFBceaVmWHMsZnBB
ea1RU/s0Ee/ZhoCFHuAgQ42lGxsVa88h3N6dO/MNg00+zRLT0WDLz27Zxh4qZ78v
RqvNL6lxKDDYWWpeXMx5AA==
//pragma protect end_data_block
//pragma protect digest_block
fMPUpWd4knTTlTt2tzENxpQGb/Q=
//pragma protect end_digest_block
//pragma protect end_protected
