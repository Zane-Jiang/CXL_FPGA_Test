// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
05IgxvVpvjQgPkZhC04tXXPP7niWEOtvVBXMA9tRvCABRzIP+iP2B1gSKM7J
dNtzyhO79Yayh67vGvx4nOsAY9paKNcsonzjImQQAHuKuwJJahNuN2QDsJle
xOvusbLDM9mVOlnuJU5MShelqvjxRLNr3cXgrZGMiZE9IkRH0sJkVSCFi4fL
Wq9usH5E57NKmok6e+YPXrsjDuaV5d+qrbyKSWrkcqbdT00w9UZFrRg4G73l
ONdaK5uaC63Odst18yfcO7r8Ua0mYtIjuNKYE9XDldShWjL/4H58RZwJkXR3
c2p7ieUrXFaLtDVQThaDHQuCLcqZHmQDyWdMOtHN+w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YBkAUgngaueLOz1SkkI4CFW9Fq80e6WtZjpE8MhOAYPpMLXxjU3+d0FwOGui
YlSAftdXJfwFGom+BK8nGf2aUsNX25sLVrnYVfQZ7A/FjymRFXbHLI3IwjvX
1NIjwKaGoL6g52WhRTEYxvMWuMNntLWs1YPONx+dw8Xt9uXu0WwZI3rYau+K
O3KFi5hTDcGs9AwCcTxWbJ71/sFVycwdoNnB105mi2lYnyesqNSWdAzd3OsQ
Qff3sqFsbCKiBAaFhqy2UftbZuT6MkmHKgbX4RpGgJxJq4Az8emHZgPRGDDU
9RzJY/nrR2GzxDXr32HGACGSIgMy3MxFN3B/C14uww==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gT82lWvJ5uXbyrRtqFK0CXIYjf6bO79Vk1GyHxNFsKjGbi6UpVB82WffHwu0
rGqE+Gq80xEX3gJtC2sFJM9Zkdj+dNngHhoqd+aZvEBCXgS16xgWHrdcEeQu
VAR9Kveh2brj/vP0ugCeQbtmWad0VUFBH/kJV8d1tGca8W0DrIQ5SvSGqWVs
rc8z2m9CA0a1w6dd5LRjvS30rYVkkHAXCUzkHpnf7b2OJjxxQwBmPdZUfhvr
DYBf6lds9J51qrTRYtBV0X7aHWNK7dsCczoRi4EyN5hadDGjan+rsABu+NbI
wCzmodtMInOAkragBaw/xFnP3N51O6AJUTehpbhNuQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TVvGXo0YZmWpLaC4U0UT4KNjN5JOzS7VkjxJ+3lgBojlAYU3IBgm8ViTz9Ka
diB0qt6gYUTwBgcdHrdmmM2hPDosPoKNMbUlAUo686RTzZpU4PgfPPKePBjM
jIRCRxhH3hJJPRL7HuxWKVeL39+u377CBvtIJGZHfUuBQMPuGU4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SyhAif4mLdwws0yBtB1eWRs9frqkyaIvjWDjtFYwfsVqlepeaQE7XLHsnYqP
G8Iqqm6PqSeILms6RSi8f+9jn89SlxGh45Nk22szOsEsA01QQFcfYRDoeVU3
SnMJHjdQjjXfxjJmXi05LDq9t7NJZssm1AQ6ywgZWPkvB7aA3CvaJbgJuKia
uoTvL/eb3MVtTi1rymukvqH+x0lxP30GS21kp7htYxd2C7y2B541Fhr87Ozm
U9aS4QWG4gTHeDOr5CyjdHIX4HPycNNSMrwvuZjwqmU2nf6jS5PwLyU0fdX1
HfIYjdFEM6NVRa2BEa1Z9TA0hnWd8QeyqN9/+e36dHdRHhadzl1NnB7QCiB2
2CB3cXDEYUQCZTaSDfhcrIPwqJ2AlQQsPH6EXCxVbomMwutT1012XqF3eNc8
J58hGH8dNQsP3qk9ovPdZhh5u7F/IPmXeXILDp2mm5Ud67ehgUV0oySVpUQ0
kieH/GCLbTLYu0ZS89NVJR2nVHBxlacA


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ktn1lsGDVSGhuAybARvZV3B9anQ+OGkljslKGApnydxGn0jqBHlxSnUU0XOR
ySII2nAu/xsgw2miRbs5fFsrzDSgd5uyKd9szlH95J6oFZA64epBFSc6JcUW
3k9yCcTI+tlYcsffqwBKJ1FWf/kGTojJSQ0omq6SJmnY1GoZvZA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lyuYHlH2dW8Z428msoE/gpzHdICwoJ5a3d4s1BYZxfPFzWyEiva64DTyxTj3
k25t9hYGB8biKHSYl9efC+wDdn59K3HYOfT5xX7EYaKNgbU3LCAuG9p3wgIv
yHX7ZfNRVrZma5wHcWJjLsV46nQHb9wmr2/prFzzfWQJIM48qos=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1024)
`pragma protect data_block
cL5ZuZVwFbmOsbp9YCIUXIC6lnL1lJ6Ca6fcoO0+PTAA+shmCTHqmpwVy2uk
AUXFY3+pXFV3oveoiYi0k8sOkBkv8xlcQlmSkokNUr9UaYqt1QDdAFEZgUWR
5ZJZxadr7Zc/qzJ+Wud1WqtPU4skgZLHsObcD0vPjbBpwpPaZbKHnG7h5Bol
RpWWpTXCTaAzbPejxSKEY3ufQltuR6LO3ug2c36G3efYVIejaqUMcf5kOsn8
qDUv/orZv4VlfVwMnqSVAOKgj2dPpKv2ziM7aWiKgtPCamcSN9vkXpWHHYb7
SgMGtv8bUfmbUh+2AD3Epigho6WGOPD5S3T7oGtCzuc+WlwOUK+rfZCfsfVI
3kA2xg+IMOdya5n3Ln/hcdXAPgmunW/dEGGhMYVvcBDEk+wM1V3c9vz6zI60
ImRUQsoJZflAHX+kSt6B8xjhEWiPniARgpNDm5E9Ika2107u+cK84C6Nq+Nl
Vxbf4AcCIuaZbMsRyS1P02l7Pc+AL+okHMrZHapMzY6lXT1bRdXDFxUxxERR
H9xd1gBsnCzuiISrWJd7X7yHoQvoYnRX1Udnren3aFDBGEIZD1CsMOSmLcGX
3Huz8LngA0kkhU5m7pIA6LZqIxtYr8NalUStUTFlTX9o1KOfbf+e05rM2uPH
DZK/uI4UilUygTyQ3WLeFK0SEXlR2lB6VZX4xHMavNfm6QqPZbmzUhC9rdOd
xaK6P3wTJhJ19+9QoMRJnpMDqG2KMCQgCXG7OLXK1cuIL3o8E00+zFy5eWVo
Vm6S6xDZ0rc3IOQ8vu4fdUQDBE8ftO9qPzuA1ESvfKDl/0hdYxLeogdV3ghO
/jPgbm/vwGnYrTfirBKkPoaFGiTde3e+Mg1WAJlk3Y9Da63cnww1UWuWgG7A
23M5VKYddxsRCNVYDMYuB+sDIBpOD2O6MEd34Qv6rQbvAoGDq/wMPLXXEVYq
uHqhInvEXMaxfTGaxpHVCfAJnTBTGTrrk2HLS12WIFG4q3+kAvw7ZqDc5wcN
1mu0g2c2HhMtd9hoaumeFp9Go+hL93pjGaPJxdrTtSZGji9k9+9KXYl/dNLZ
7BmRXRlFNQATAyaUH8tXOHBNw5DPGIRjNaNQMsw4dohr/bfZUrxKOczWSSpL
/tMPJ5PrRQIxqy5AqTo+MudXk8zVy2F4jv7nw5fcUQpc7fOxHhEIGALWBgNE
6qov4KZ5wRxAaSz700KsCql8pVRLnHTRoJbKBq6KR/cl4ROFwgt9IS2vcbDu
yW+ChV3E5DRiOP679znkKe+UMBPPwqPl6E0UUP/8F46PuIuK0lGSmrW0VGCL
53FVzOvdgiA1No61YQ3Q6TS9rZ1n0Y/BW6q3xME/aSQaKA==

`pragma protect end_protected
