// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qR2IQpLMSKXzOAStyHpIa/hIUbwgTFd/zL5KAdmvQg9QeK284MNNN1nZO8B/
dEkKH2gHJEPcb1l/Sso1h3OeTzLU/iBVf7KHInyA0BB7RfbM+4P8WNauVemf
vmhi21swHqCKiGklRdnwgaheYB7MzwoyNEGSNXCXll9fV6RVumzGEL1yKJN5
eV5Y5hBrhrUruVej0b578Byq7AVOLtR2jCBRQjm8FV2+xRl2YLH1lD39B/d6
HhbofQWr9R9gJCLGS8XlkXwOGGbFBwkVB9GPYBFf2HohWSk1NjzzFUed6BUG
FYTS8Wxm11G/7ZLmuoPx5V4ZSbtgZ0jwObKJ8n57MQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PY46sPmkksSGaoP1tQSduRg8KmywM3zDdMvWPeUDblIRaf1WCKttkxhONT45
N5e0EZvtJyoorxsq60thCp99eZjaxrcxn5aAzcurrW5UMu81Kl4vyyBKGT6+
yF5QRjgOFjR4fkLcbj4yhR9sU3ES1jBk3Of7iD8iCdwRJsQka9o1Nt3SgCmj
bSC0zjKb0i0RBILaVkJsofmBqRusfNzN5kChVTZ51C5NKcK6loQIKZjoVOFb
3TnxowbA0Wk0EvN6RueKG0aZaDvMblV/B6dzPhvoxGFOb9kEaHsRA02FsKar
K9VwoAnoVuy8TlnfbHXEI37L2iET33la3IyGi2weiA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c7tOscDsg2WNp4+viX241NE0VfJI3QrMjHJErxnWmQdAY40OSAjaPAgF5KVO
ZzxPBFM3iB50jDi6VEOn3+v3+/4KNo8iD2XVe3iB+bqXQ9DUcZKXtk17ECjE
W/d6VfzqMmd5JyTV9O1ZYkeYN73F4TKTmQC39MyYb6YDrZcljpk9RHldC2nz
WU/ALmL8b0vK3jbYL5EMXBUO2i2i0yuinlU2szMOIxZmfmHeLeAS8Z2GDpZr
Kk6IZxAlq2LYU71svxA64ALnfBDtbT3HYz4ZSzTH0nxunYKu5Nmptc7QM+64
cr0sBK978yncw+/hfcmk1XTcXkr6nI8htvg0aZkTsg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HU/euiZfYPENpoVuvCI+dU/YCQmoze5s36Z1p6VJc9ABKIHGMEP1G/b272da
mRt2vhxvNfHWfAFEbu9eKbYEHbd4Bu5gIXrhXtY1uBLrVo/K9cmrMJcoHyLt
Z94qd6YR3yFROauqiQHKlQYcVKUYBrCr7F8ox3ZxhRVye0WzX00=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
u8H2jwu0Iq53NJ9acy/oHULSqlrFJ7pB3sPq8PnQ9Qh1sDMYLgstFy2SEn71
Tr2m1mECjDt5SAiYiCSkRf1tegWQ0G0OkA8MFvZSBQPpaJH0NAi4Xi2qCM6R
sOEyRE7VMzmO4bKUgoHWl/FFFhLobKgiYqSEgT2qvBA8dvNXJ8M7KC63SLX1
rllQzhhEni4twEwiIWwrTEfUWzZlQSejKP1MUgkdZC21MCZsDadJ7ovNUI+I
r0gQR9g8eRVTpzeX0kPBnh8+joaVkgLAu1jcVh2/OGR1EWQiEb4OJzTkk1nh
fuNQBOysubVE9kGcnw8ciaXWMeyUAWAvcHKFDzpcBTSt7KIpxogtR7QNDJ4V
ufdCdPihMRzQyuLiwoY6EW40VQndmt/qfmlLfbwxvqDNJPPVgtyn7bGayH+u
epPvpStHZ9hoHwt+OOzfZCx80Vw8hl+zKqQ3SD6O82X0ptQStZq0PRcDclsR
u/q2ZPM9wmLzg4Kq602qd5SAvp7JrXyz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QSHgz4LSoLvISbtaYtqIfb8vWut0YIBIZ0W3tCO8a4mDiVzr0Xc4A3t3ZkSu
Uzg8Cefr5zWc334kRb5ic0HeCWuhZquqHU/GZ3ibNV4jygN5Sh/Q9gfHoo1q
O45cGgQUzeL/mV8+i6QX5QzPaOifc9f9gAAKqn/7r84SjoBV/nc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JI7iYfqkuATLp7tDCWFYQZFBT2pX7hITTVujRKCwxfwJnmInpgZr7anqjadH
xd9ovZKaIC1dCIhms6F+DV+IOUr3juHrGU0jxlRZVzXshmkwt42EghK0BDoK
JSJ478EdjsOHt0E+4FAy5D5ZkAZDaF3eaybbLZnxred9yhRuk1Q=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7056)
`pragma protect data_block
hWywvQ/YljbAfpzec3Ktl8i1mWm7KnCzGTfaEk/BIw4/xwEk9oGxNfUUZvcL
rd0J++8UAcgK0L9Hu9A2Lunpin1rfXNlvsmhdEA2CV+n2XzgwD2I0bDQORCH
g/Xs/W3YXns8hu/gpv5VuIoBIkgrzoHMYU5E+QYeD5TcytjOY94Nf/ewYCRV
5+YrXDRonYnES64IqT1AICD1zyBLCJUt9ZmBEG/UyjUAQhougC+dfoDMpPqt
UaKNRAvotLr18ZP77iSTwGe/X9SKYvnOjn7e+SMEBzU3uJMxfUcxtotDuTG8
qM/63aMM0Wg6mx/sDeXkzp5UBca7wQDgqJqQ0DWYMMsIy+aJPuCCZiw9nCfh
XBNnV/e3Wkfc3QJh/rR0Zdo1hO56yopsYg2bq53Cpau4V6WIsrz6xVWdBcoJ
Fo8PUQZmokySysGSAbpI2VgOs/3IjtsoW8dAlrPwgKEJQlqT1KjQ7WOc0VxI
zocmxqwfwOhYHBlBNm0NOuj5VFnI5wR7kKG3b6yJDpPYpkTxEo7FzXIQvTwP
ebEVCORR2TJ0wg5szfAt+F9dBXbzvixAJalAqaVF+EuqP9O2GJY+kFl859hZ
lxzUsumml6WJU29X6ryP9WEwrUQeJYfqt7Iyq3xEwxuuhWmqE+R4zu19AnaH
BYGqgPa+uNGMaX44m/r3mG57rmdzWgfuO1CU2yC6WvcOdeVt38VRyFnhH0FE
AGNbo7HH5WtW/J39oH0Qy4eo08XP4UFxSGOcjPfxnI3hIMEjTRkglzZ5/n33
8T641iPNvIkP/vLQkinbyUOqLPq7scZF4yya9BI9faiExo38Bu2Uef9u8NaS
26Abr/MaM9mfgWIvnbN7akeQA2iFkfM4jquRM68BpVqzTApf8LQK7yCD+9e2
UlN7ZwDz094dp2MPWzBReqdZbSG0HwYPImTxUYCLAEXkvm8wsR+OsF8tNkkc
CMv94LevDrqaEtzhIZpj01hqNgpIBDCVTezn+swZgSANTOhEoxFFIinzFXXU
GOTx/tLBdg2lZaIfZQntHcC++OmyyobWufr3Np8vpkjwpjNCFe+Ib5uPPv5q
xco1W1+DMuq4mD+7jC9ZkKbavk4mtLD1XbTNPn2Jae25bLfP5Ok5+iwwLsWr
dcNScUw+N4jBf7A2pyuTZcJT7gdgnihAWY2uEFBp0MPCTlZIFuLOELIeM4RP
EtnJeiyaYZjLuNDlQaewdamjQVxpt/jw6/iKIyJ33wHE/c41nCQ6x5aq571j
aikL04+GTEgsRWAjCMUF7PXf3XPPtuFE40vCFIyusU6Nepnkhu4vldH3PllF
384uGbSZU12p19obh2VX+B/moDOpd+CoXKvaUcmB7jcwK60y/bo7pmgjliPT
GQtxa7CfyLkubSr+AELeI4Q39qPlEZUkCBWk5+mKRtV9s2WLGGtAcZ2n+3z2
JXbHDe/xxXnOFhPfKVuSgKnIpaR5NdGG/MTQht5flcYjylQFgx4CQIHElfyq
53y6m792JumKSj04IWAo4rlXb6GhbIOJHlLj31oKwUTsEt9STimtfgipIz9N
HSlgagIgjPdBEHw4FiWZN/zkdOoa0oig6qQ21eJ2cpP7eqdBzmz3okHgWEDO
OA1GZ/yIcMKFTN0v5G/WClQwHicq6F6GBFGP/ESZaG5ydjUUq7VitVl+OALI
TSBU6Rad0Bvbz49K5YL/WayGaxOiOiZ7xZObvruS31xBRN7BWWsmDkPOFWcE
hdz+Oly9/e2RQ3vikalQGTu4TUYpW/rfkgLvzwSV03u85A/ohOYtfTVn4gty
vi83HEiRf6aQY74yBKs9eTdr9t5/aMR4843mBOO1LcNGxNCoYGTnIrsXzPnt
3cBd9ib0GLw2oMCercGd2dTquB+dyajm+NdEb7bx3S69DN5jAyIc9N8WqAbL
G2n2JUOUU75HIXPJ0bPUQC7rOPTHyTIvYLAKne55J1+b783Z7zjGY7v2wPRg
kga7c7m+Etq3QUlTGDd7VeSTX4ei6p11SY00P/bPGcgZpYL0sPw7xXHAMsR4
EUhmwvD5fbq+KKkGAFJXfJGY58J0DybLrJ05ULwFgH7Gvj+6gqfldHwL1HvY
BYhaPVPNWW10fZwZT9Xq8WUus3axZuen+2D5/tv21TzIATleGpuYSUj9ssa6
dFLatC7eX0i16RMFxJicIhFfgHEomE4pezSKWOtezJhZWRSw9mqifDFJxWBD
gdoGhAOLGH9xwVvuzpxiZcNtEzfZW5pgzz0xqCmHK/yW8UtN9u1055Pl10ch
xgUiaiesMwEiwlseZFKK3yKJ82p5TXNV/SgwuBFS0Jxt2AxHEb/6+UFW3p1r
5eztE6OzF7ue5S6x2yZXM4uSrfvX2U586ciwRnKsgw9eMMZcCwAxIWJ4HVjk
rz64H6IIpSS6N6rsevJJ9jUH/jVO7BUQCOUGvyots7yFAeIhE4eG+71BUPGH
i7Bo+VlyDWJmCaXvwfSgC1iz+lrSJ50rQx9h4Zi8hp8aAnzoz1672VtS69z/
CzWMkilhtTm2yl+XLd6CuOIj+9daDN1ajHFxmGo9VbsjGbLfiOzztbW+IZPi
HRgjP3pPeQXRUJqEnqw3E6aDAN67wtawbU/og7PDPSlC+8YHTF01tLLmZyj8
a9/DH5rUtRNH9Mh8zTyOA7mBgvUXRilSXGlsnIPi22diiflm6p0PKu4/+/7p
mRs9pPq5hIJhWorwQHy4jPv5CX20tRidYTgrVVvMeJMJJjjAaboK8lWnipLS
ogqZzDLt6Zd31+wOe3x3itt8uJkGcqqBK7dxWk1IDexfd4TIHE1tXuDvObVJ
ztqQ7s1/gZDushmf5dtJyo86gLczs3CGokYOwKxB1Kkil6XvRQhdkYSwxqCI
zWhi88MGQmNpD2FFJ8GvJyYvnxuYwBySV1ouIbQ13NY4kwhPzk38ngqci9KL
FdS6HVEndkDXJCRYNgkR3yXcatqGHiApSncsnls1QFUKprl5n9z1LVMA+jG6
eOnbYhaNrCyYRsPfOoPoeRx8DBv83AXQQbFhOe1651UeME5tYVGDlzMll7mC
SKNyJdci0VnI+8ML/lOI4tnh+9V/48h37cButXy1+4C3ksung7+fF4jJA6sN
pTwhvrc54DYQIv51PBKn/AU4xqXsTKP8B034FFbs8avmnnqJ+WziUkL2W0Gr
TStWtWdFEEyK6q+YeeVvv1M2Q5xANbORUJ/N4dcAfKI/iTFhK1arifSzpYQ/
X4k/BQZpTHoZJTVkAkvUeNZSQkHz8mpXADTpJQ4pSQKtoMjvpRVZ8J/FAgHT
DfDYOJBjGl2KrLFkUKi+XHr6Yt9UDtgonop6edh7CnRF548y4CZ4EQgepeGf
aP3AMtLTm+IJaObvUqx1Q+O82fv8doLacc5ZuVlEuqTmU+A6+yTfIwqlrbbT
+W+MqXT1SM6M/1Nhik9U5/7PioZQ6N50VagTjv6Eo1zprXuXuRVHPk3RusSG
OowvJAQNV5a3RB3HbZnDpsRw6kBeUexfJybTmqEY9r6vE+kX+lE3RQhKGjt9
EOjeKP/3Thh/rM9xN2f/62kA/OzyLBCwG2rq0DyndH4zurhU91Og7L8gING3
hywn3tTE92lc0RdXDhhl+t5lOtl3AykRLBvHV8fSCwiIcL5jhuTJSNxXyVlL
114UMVqe9HFAw+nB/xnlMNHmSEBrL+wyEQGBvsi7ieH8lFuELd/dZk8bSOQF
0pq68sKIRffaFQzUsuMWzflhqVGlsiLAQgmzEBfm8lIQ7McOwd6EH9E7WuVj
VUKwncNlKD8XIsGT7xbqUU6ZQj53UM6ydFQIII04cRoUlimvw/RRCZcPcVkv
u0o/fnXCMDNfIRNhjGeFFtuHV5NauDFcGq4IefCqnnExBWPuSQJx6Qs9CBS1
kRg2pEYnf7KcT3vqzmbuCbNVA8yn5RN8jBxk/41T+4UK9KBZuC3sTzxupZL3
3ioBwHgadthtKGCPsmanV+MWVvVLuDP3UPhWCZqXqgrL1UjhYwi7wa7VUlrv
MBAOfFU5jza7jChDhVfaeigb5oU6OsYzAXlRvfSwGDA1jnod2OysBr+EGLYD
7Wv7mi7TJTeA6WY40LOwY1GZtbRn8yaIuQ4cPdBBWIlJ5jIKT8f/XR1pYeDZ
nC0OL6/o3J418UKOKHapNwTakWqgpCIqcfujFf9a9ucRHvhTV8in5jgQcKIE
q3VyvqgAnqJUUnweG6iDYyZRikG9+jiIPvMuFUE71BAo6PGxh44B41Alsfve
9TpCZfqxzV1MzQpKKBjjclr9FMIM5XphyA2ZsuF5Ei1JYBhBpahOn1HAIzLG
kjnMxRC5gvoB8F039VFSbc5QhYONALUMENAPGea/TKnBBqg1ME5LKbQvoVYA
SL7lauZdQHFdGns/d/v1n+goSZC4cxz1x/5nziRHVJWNvjWMfYozbXmckQyw
Dl/LID/Coxd3C0N2VeX23Y3mH0uSHYtwmgUQ2wcRL/pOCLQUSu3/Qh/UWEzF
Ngrz+4XRrkjF9v/CCmJl7IsyhLZ7IZR9SaePZktwlyPXhykokL/wJuzqAsn+
SvbkFzIYBdeoJLFfcOd5wS7NSAJbmYNl4zbCn/OH3OKNYuHbxSwNMayZgtrW
TS9zuOxPtzBQAuJIScKGyCb9JHrxEoEyuba/cBIkUqNsJ5WmQ7dhoBw3y40j
tTxE9xrreni7BSJrNJBH+4VDWSF2Ydil4oq1gXNZOZX5HJTELwejRJVn7Ic6
5lFQ9mBhKwR2WnOxz9xNtzxZiWy+KjK1AA+iyRRICOK7SGZvr4FVSz7aw0+j
XbSvPsHibxow1A6cLATB2a4vNg7J2l0aO3rV4FjXt5ujMx3nDDAyN8MT4O4Q
z2kp7w4k9rpwh6w/zxiP/GdYD6bpccZSc3Pz5lBPpbsob46dQEGOwvwUCvp0
9gFrtpZlOi55uJOrcHTtdBaQm5m6qPky/Dj2ThIMbwbSxeTLnsxBhxgNwN/Z
rJ0dyLSbxdN7IVnD8Q5UOjpD65bT4NqE0Foo9L8CL/ITZxlxlyDOBmfSZO1a
iIbyJ63AfQWM+WBQQ1pBXWnaGbRVq7YRVweYtSKqPeYYjlVfjpuy/E8wzLeQ
62PMJIShi8qhjf57OafCJCpPwYypXoS2OQScvkJVKwRiCjtkxil2bdihKBrg
UOmmeA2AIcadHpMXlVpwRAcxWO2Eam3W1qoSWJ0vyXUnxb8nkZWbaJNT8cP6
MoltpDYs13iv6alF/cDcFjFS8pAlx/zG/8GY+6qRRHxlA6T1l5e+1xytErmb
gokx/IV7WtbIB4coy5LYIVijXZGLBMqsQkKXeSnZm4agFR2xG0zFsA9bKCUM
mJv9qdKPHiuB8uP3SrKCWhGLSq5Mj5GctwuMn2vDxe+hJRHylAJtjOxJ3Wxq
tDi7Uncj/Yrg1XeI/WhHh5DkNnZgWNiQuWcCswFQOItXhh1pdCbLyHKkvlNO
QmYZ2Ms+oT2RNh/IVWHcqtz5uYe+00I+TiM6aCR5+9DlN9qGWVebAYmRzJ3v
ksoMTXZRrrpasIcaZ1o+rdZ2XVlS1IcsxyAUf7k5Qu83NY01tACU+4uEz5e7
b6vP9w58b7CqNUitP8JwyzvEFwQJjBnc7HuQOaqzsoW6YpCkPDh98bo8kj6B
R2HCul1fJGMYpmrzTPRW1SkP/JLGPx2WLMY7TSVrRwjwxQtbZjCySxCKMwAR
nF3hh5qTN/aI6758JCb9m/uRAi5crxeHqzIh/bZegj8GOZeB+md0Frdf4cUt
uVe51JSdNCGz12r8qPAh8agUMLrLvHflTtXO6ve3mUYacQYN0AyG8TDpmOM1
Ggf9K4sYipC4CsudMtkLoKLqwlgdW1IU2Z2m1srArsSEVw3TWZFKbdOVgnGc
0r9NGXACt9Av4P3MkwhfC8ovBdw5CAWtBVNEkt/44GyqDwRkNRCeDA6H89FI
lHE6S4H4NENNv4OHzuiF37mdUEI+oLw7BvioRfsUKXFHgcOocYWfb4ejlPPg
FcGu/sFQFXTZqfbZHfs97m/5QVafqSK893wBPp322xjsy1OvIuOf6srEstsf
Ymm4GqWnewZVajyPMI9PiTDie4YPYDeZp1FIEAEvwq519G2DWRQpG/PTzkAc
pVIHan+orautR7J6uPYtwQUvwUCYq4nuIyAWpZR1/Iyk3LkDikeAXQyZOnOy
k/uPkj5KyUi3GmjH/PfA+0PTNcO/nCAjzg50ax6MZhZwtsSHgCGSy7ZZdHc5
vukELlFH3LeytjmFdEUtdmHskl1BevB/NknX8pMwqeE2Z+OLCMWX2vBMNAbm
hbdR6ycakNX/2FFjNnmLUtzdakZ3rgRIygeoFd5y2mKMOFNTf+NhTOS1bMOz
Hlonj7t3/J+TiHxFoHms41jyAvOhlfnyskpIU+FFucxxb+iGIiSPvIv5ZK+W
2EdiIRPbpH0JzGJB++Ezb4cWuUyGqExo73Kt1lW5nxbp8CqucTSaMIYyMMzQ
OIRbUt3XPKHK87m6RCl83BpTbYMQUjtJACk8mYYibsqEeNpPjPmIRIEr4lsD
dqTwkhz0+L70YkKi1XPHxvhrXbJ/1MYcenC29jgECHdp460dZXfa/XUS6zap
rriXayUiY9nqdUtDogpE2TDvyxzWEF0DDP6zUY0RXVVBR0+2xtyB+03j5ILv
C9sywObH54rwocuv6v0W0/MLLbnyB3lqrqvXz2fC56388TpUYBAgcGrWDUw9
OCRzPyKP35sx6VOs2xrjGAAkCV1tJdJRiTFOq6rmVUN3N7n0LHSploT2z40a
H9sjcXHMEln470F3Qmfs2VmDIh2bY+hJetxYDhVm4wK1GyJvKyPKuY2a04RH
2bE1VPvE+51TL5aG75d6FgWzUQDRAr5QocKDAwwCwH0kN7NgSGPiNUvqs2rw
akGJlqt5qNd/sCGoY4lxQwRT85Vyye1j71tsm/lHtdYAj88k7jaKhTF9YPrX
4HRIg1+zOl4IByCHbVFaOT4g1uMwSg9BEAA+Oy7w/9GOmQ+n7BKrQuaxxWj5
pjuzP4fvzxAZHYxryV10vePmOPM7eZfiY3ALt4OsElm5BpPibCFcPLCwbnNb
S58OgfoAmUeGNTg9O+to6/wYOPdqECYeiZys+9TbcXtAr4Chzzg8by06xfkJ
HVRE7P+WPACIy4N4jYyixIpIwpBU0VKirvOSSoBVcDyo5i3E5eI1/5gTdxyV
vxlb9+VBGCdnwRIANMjvBQa7MZqxmemQcBGOit9yefohud2x/O54ESa8JstI
CVfM4xV8tQTRDV3LBOrEQjSFUBLUYtlSaFyA+I6TCeuMg5FcmhOB8ULobqlz
dTMQL9dxRmOhwgA5OFIZsDgRHnnYu72EFC7L71pkkDdtZt2n/+OLxKylk/iJ
AChSuKjtJxfKjrnUPokuaqXg43qpBoDfmJnJV5x4+ajmXkeoi+01gLb3EJiU
WTPXPfgY5hm2QtSjtPlsHoEdJAWe4xdu1IQwC1Lr2F4RYoezeC6aXtXqACif
BD5lfopn25A9juUKowZ/U8e1bB9LGYEIALGaoOA234C/8rWfG+Wfow19YQ6S
9fh5k79IfFzdTwRX/K6c14v90vzdeCqyPuxsLMLeBSopRHp+Onfg20uXGCSo
/Yzt3aQRjYm6OgEm/QK0+g3MPh5CLNQXH7eERWNBdeRVmfCxdulpjOh8nIjO
FGLt4IugsDE2WqghpY13c6Ns302mGcNnxdUIy7wb7oZjevmIV4IC8lsecaBV
+IMAwen9DJoS80PGgqt8Wgp0fmN0phuK2JuA7YIUx5qbUHoRY8SIcAGhbQw8
kKwtjex99WHDymifqIqQ3fLrC9VxQH+ithGhG6md4X3NHZp4L3wFnCkuWv7Y
U1PbfVprctRV2MuUvLSuOTCgSjw+vjobM99DWba2RR6EiykarqLxMgxNyMoO
/PUAO2QNt90+GjRHQ+HUahhy2eM1rXRHtT/pNWDQ3ssAz9ld4MwGhDhN3P/o
LmyVxSTjdQ9BN6NSeAUrCEyIMI1jbARlqIA6VdEitQ/n2ZupEV+FzVZqiNbU
7O1Eta7xcUzUIk2Ewj7CBm3CtGiPEplGqJa6T0MjJzreHI4/gOM3pZmFjJVC
F3kMPgA1pEHUM4iyC0HWLn0VtqX/Ktck399u/tfq+jgwp2rBneCl8osNW+1K
8j/235nq+ozl3IxgaabXQeSMnvYDzPwjGHl1WFcoCA7olr6fJ5DMiVR9uZVh
L7T9tV1j79/Ufp8FJQG6iEjDXYGuYkIvQUfJhi4bgI9CnLJybh+JRONahx07
ADdow5Z6tI4dxL2VjGTmfvNiorcrkDFkSD4Eg1wC54nk2CX6/d1/PkYz0UPP
+2gB/Ii3KsAC0hb6IlBM8Wazpxu7rtb6MzPTP4ILQfVe6IKCDq0PZJkTShEt
Flb6nEUkVjWYaAlx6vTovYfIXnEc+KRDqoPsgJzwK2YW0s7b/90c4KApR9Cs
y6U5bxiEZd4zVM0s5je1437a6hf7b33fyNqkuOPQidQnQ3t8zJAeow6WQYa+
z3E3jJf/zDOHyNfOuws4EqVPKJqwvsebMuTtdlEL+ZAgaZkcgdLgSY3ZnD6p
GouR8rTzHfgfUvd44tQ6ozXZLI5uWf/ogWmPfU2vWKZmSAQMUksCPfZwP7Ue
nzv1FbAZjaTrP8ewEW3GyWx/f+nddCIg+YJ6e3AthtY/oS4vH5dOod4jzDw4
jj3hSQfS/OeC7j9TpSQjitwa2/riZN8XrudVxhvqt9+vqymPN6cCjNbZUxhK
DG/dSRtjCxfPrFAfOYGSx5vmsURcgMOx8YUTD20vVhfAUXvgfb9uCADUB4Zn
/Z/oGMIiviVhCnQUOqbpJt5PJdHqeUcNjx4dIOO0H0TnQvAtg+rLOOfs4D69
4bON+4gJSI5DrILYJInB22psvcWKrGlOOH4xhYu6q+1PXoRCmvU8xFNV8PPA
sxc1iOPkNfY3vi5OsXbWlR/xVUEqju91xRHPFeSA1LRL5TF6xdJbzMRgsBm4
4b+sBfHqfQo7joNqLzYaf4au9Ib/MMiKz69kHgpq5BOmmHvrKZ7CbINlqsfr
OTIhnYbt5wJ9s3vyPjMxTabKcifnt6wTM0rZQIO1ER+BhPkKdW/5wzjMHxNx
OsU7yxca4Si9XoSfij8iGkaV6lrR3t4y5X//iOGZbRVQKCsCSqGtsiwVLhc7
NVgaABO/3lcXLq7lusbVqHOhdHDyByBoIK2qK/N4qfbXatWaELIRtwf60C91
syqz5yELztuOiUrpB3HZR4CY4J35aZKmzYt7g6yrHWvUv3qwxOH4ISy+9ujT
IbCwcvXujyZJNwrXTFQNnoJnqxgNRBlaLYUytmKzHYdWC/11HjHAROrBmB+t
hw+XBi6CNNhq2E1zcKOEo06zIZH70bLNajE2lMt/FyAnA9A1

`pragma protect end_protected
