// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qOANQ+s6S3VOt1L6DFHmAJFydL+j4RRP11sjxi0Op18teNUP83OR/BMZnVJ3tIF7gLkMRXxi6P1i
BqvXFzZQkrprP2AiroCU5TMXCvh3QlAkVLmVOa+IFDdilg1EYdF1EYgJZoxGAsOZ3hWHxBhz78sU
vElvhtdvU2NaR2GOsuW7eShvv8uDIUq596GLT80gF2W7UlxuiXWXjWJ6nLGFBqYmLJ0m+5edDG6T
JvMLvgaKv0JdxOl6bSSp2nn3hgmImPldf109yToroYPWWLy0oZcZj0BkV6ONUSip9cGdAwH+CBUk
fLvfom8J2ekXfN+rTztwARMEpHQ2F33CaqHn5w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 46352)
QYrAYzjhUZd7Stq/yfptoGcI8BjuNb8WyGnxij6R29z1ldg7A3rdcAp2GiwWUFuilDrKQTZYHlgK
/DRMfX+jFPFWMeVGTbLpip2ou/YoajR3V/zwbCtRSIKwuBbOUtCE1mRXEhCTftgGU6LusJ7+oUev
yi+sGvN7GV066LhSbD+Nf3k4BJvCdWEzmqLbUOQ4AuSC5o74RREfUtzYFBaq1oBQY8wQTt/a0N3i
tVdlS5dlb2Vnv0FmofpONgMvqoJ25QFcoMlUsM1G/PFWCc6dFMFR0v/oCptsg21/muT0Vdgy461l
27Zw50mNcaec/3mRyybmyPxeCvbJmrUdDMQPxeMDVKomFO0tkagkFswLRVF8zfxTgrVeAjnzJddy
Wd/nJqIjoo35rIWY0QD0wfMQitQvrPWqhsTP/hUYoObKWQqx1jYDZX7G8qtbxdhzuQPfgQOUE7gh
SF3jQgf64lZLT5b/7jmpFrNQY39ZH0GOcdG6Dc0XXn3s5pwuROOKeIgb7NR5BIim8h1zVmXP+uf+
8f+5TvIMQPiawnNipsU85QtNmwKRR3H24CAZgifir5IjRRj2vJM6zcdR/OJZqKgl9LS/LputQC71
WbdRf7XvrSMFDgT+QXEVQUeI6BCec/JrfyYlXWP0v8T5YhzHlsZopNvhzEhSgjr+GE7SVBJDrlB3
PohC8MhSZxG8tcp91uNs/STdeKpmZD2644vAZXAP/hu8ntEX1o8ZsbQ204T0VMvC+cHxmyVcq7L1
QTicf8dAZ3PXDKABAx9EufrPSkJGO+S7oBZOqbDoFrMDCrNuXJWCzoePlx2naELkAvSLQVqM6rmg
CgOCGkjgZYi7D09WWz/e1GaI1prkcSiMPGfE78XywKYJ4gzShAFuzqCMsxJNW1iUuk3NNMOlKgba
TnCIeeJV5/YwXBPkbP0eXopJDB1YCpVBeiHpXPQPFxOGkfqXuYbiHikKGtOthHTWRuBVRttasm5F
eXpSz1x68fbxaWpL0/V08Gwk1orOHeirCJqUhBOwkUaCM9CwE/AvUx5qwvPu8lieOUGxAG6jtmoh
zVvsVWzvbQF8uJeJFih1/gW6aAPvp+77ixt6qLCIS16F3D17nPg9URq/IgoI3VXxyNgnzfWBuQe9
5R0tbulSN7hmhZk97bNykbZGHc8H/yLNEj+1dM3jHs87iPwe+5Vs3ptvuy31HqM7Pz309AEUNRay
Egwg6YfG89CtEfa/FVn/CoG2O12PsZkHqxWwVWcdiIwi4IRJ+DOILwuKdsei7ULTYONs8l+/v4ii
BH9VSTURPWPh62Kv1/4bipp3YPLJTwNGEGJzLh5NHtUvmaO+qib2MIyinmTiYvSbqg5y7Ed0TESE
cuoKo0lyVlBg1jUuhwm5vP0px5OYxs2Q/WrCp8kWkQuU+eXYgiKludz/3DioJvZiWiQlQbs9+c7t
qhqD4jTDcuTAHuAXGgogQsN26i+1UKJ1jS3KlGDHoQL6auCo33qLNR5jWGs8tIdaYUeQAy/lQcST
DRXZEAfiXquOEzGShMhEEnekP5dxA7nnZsFRro47Yl/kPtGy6CBQQSVZ3lskMliguFgusslx0bXB
5eFlvr3KGzXQ+YHcdKAZu6oP079mVvraRq20JesWME0HIaAHAQLyBqt7R0DWnD8rbbcIsHqtz5f4
pYYpjCUSzw3386cxLBuF27ojHg2p2JjaDjSpYciNAUtTjyak2DufOzgQziCJPTck907X69xFYWgt
LbHWbdzlBaxgIQPCGTkMjIk+ksgly0af+9hRVP6EWfVQn5fUTz6JJMBqLPMoJFptTpV9lH71w7iJ
vNMWrfd96aoWQda7vqLAWdig7tR5wKMOnDqnOtQu0w1AVFRJBRifOrLR2YIxX06K5e6ex+zUU64R
2daRKH3tK0rDtgWWBdi87SEQy6Lb2L1U0CtYuRWVHN2iQ5pcZ9qqPDRLv+32ExguEowU5XzlciKN
HltbBa0zIUzFyU8+tlIB+b5IMCvhBCCUQkr0wbSkKLfZjUXj4kxXwL0YKFBBr7/ikPczs4sZK2Pu
QmdNE7pDhv9DrxXaCFWfhLpCVOUNzZdFDuaCaJ5/Zo5y/O1qDhxMTQ7pgkeJxMbHth1CxorMQh5h
Eub5hud1PGhij+wf4iJOO88RBozQEJI7DWHD51uVaAgl1pNt+PNphZ56CpTaSwunRld2u2M9hhCM
UeSyyZX44hIuH+83iuWP+OnX0th+5nyYyZvjv+CpbtCLUEuImJwfIrB1NVTX5KSq4VURwWZpiycb
+MjHf5O42ci4+WFIb0TxThVaMNrwayKj+4M83E6SgRDyiWO7aa2mZpPnWqQnyC9qcbpi4hXy1/1Y
p8fLNhcV0KS7efLDDhAc5qbV1sxadhM1Fd55eufcdU+WZp7JQvzaygxz9IRKP4dHuPxQJnfQ7WtT
K+4zuL+yYGaGFpYknfQvwvMqmkD0KuATyVde2PC8YvSbFokP8BxoJ74E7OEV4ZM1IP8ZKe12D0q/
RIF/+rrMBUBAc/v5OeokmSeYHSfMIDWN9Ih42OQfbCi8lF8zWGsm0nnQED1PtUWKhUZVwC0ltZ7v
3rpQAR11ZuzSutelaYasMrxuqzGFix82k+p3Y51lnDGNuqZ/q44EwdqAgGoT/1MOcrqaINhDz+1D
RwE1iMm48u48clL6j2eFzgIUTeXN+ODg2NgSFhp0DzMbZaAY5baHDdrCdk+pr4lUb+gw/34mQzK4
9rNxXQv/kcnqGMfxTz/ehaN9sQzkhjNIlrft86jxmfYpsrRIOQDAo32xEBciNmfbE8CVJKWnzalC
NUe6yedhVfQRv5jEOP+2sWzhhrIhQBly8dkDUlFE85eg+8Xi8hv0aYPhWd+wyg1JPoTClK8VveET
Pxssox/hleV6JqpxB67sXLwk8ll9w0djwIf5nW8gnThe5B6Z3VbzipN8nZZH8Wyyo3f4IWE3OL9n
yF4Uw59+2B5oM44z92B5BtmukBTNrj3fQX41WMxhw6n+vobPsjdP48aYxI2KQvzehsA2Oe5xudDi
aBHTitxkQOGywIE0W1796l1hI2Zsv/0WYx3x87cB5Az1eS8VRPM39SeQz1DjHWJmzprYVS0K1xP4
NtwCrEVyaxzYRHZD6izr84GCBPrLahgnbXwGU/P0W06lyv10o93eNdGwoBxSwPcND7DsaPLyt0yw
LJmDfHXrWocWn4MG9n9/XHjMxHCj9WEtDCnCWvOBrfWQMaUP5UnjlgS1HlLqjYeY9lo+R0zevil8
5ZsHHhLwa/6kO7FDdYREJdWBz6FJ+5j3tyIqpz4XKR6Xynwzj1ZkNQiCev+K9bciUpeNV2pL+Qx7
8EE0mmzrpuHgQ6J93uVI8Kp6DBBGRsj/hy087XGwWKxJo+PAe3kjsMHFAuxWGMrQlcQi2mpDh9bR
S00HvU6gYILm4ESrsB+QAKCfbarXm//K0JVXmuCWKT+LcnSj9RcIFFyCsm3sKfHiHZPjsUbjUOOh
whAfmBxKFUcpQ+u3oKHyxAeuyZ4BNrQzifQdbjydKsM7K6aAOoBt64ZTXm1Et0ZP5u1SgoT5tFxj
7xU9rXR5awiFbSTxjiYoaNNOzmznY+nuFoFzZWYVNRS8ouF/OS1UgfdDg3L0pl4zVjIaSMhyO2kw
hE8SxJy+m+gNxwss66bemCaL3xOe7MrviA5wzYR0xDm/zbndZQuG0634BXQIfr+wg1xR2iJiPrYg
Jb6kZRWc6Dru3K2v65CMlhzMQznvs6QFXyrFuQA904nL7Kc7zs70Jev/lyaSTvY0ceXG2GdT31FG
ZH8pONWME6tog4wHGMeIQTtia/9y8xaeXcx334PmIrM16T7zHSzi1dSQ3z0/OfInOvIHSnxlaGez
g7H9EWkdP8XQjCZQ7dcus3rdx7Deu8fy0HXUYkz8bfPZ/dnoeiSeUViODRDIgd/G5D6kPNnS+YzJ
1Ls0zpdCqKD0GELqv1zdT6f9qjkjl/gMsimhnvVFZ9XYlh2KCLhapzTYwVT8d5qM0pmADM8MbhyE
RR5FED28yGMe5L3C/HnvCfwMLgJCtq3kPNEqrkNZn3/WfJHqAQSzAiGoDpHsPdcl8at7WMug0TCT
aj5yi7y1chqKCSdtY1fmBkrbQ0+d0GCttAvG6W4mtiDz5AgzcRqV0/aw/TxRjDMmUsLtgwcPiayU
bCl5PjjXNR/7dZxafw1u+fGS6VjO+6o9JG9E1sSx/xKzxscG87kePF4TyvuV4IiVcAN/fCD/lBBm
1AyzPHTU1SfwCdZVyranQVZenwHcGugY6O/PU4AuHddg5B+k+iwYMWUzUyo3mOdJsXiI4nKuNmCV
Hp9aTwVD2daXG4bMJhC/utBGEgKFOThrxnbzdLdDmDdrBh9AWqr18cgItzVyYsiAiNLxpYb6U/oM
4shN4eMMPO94r+3Hi0MjZIbnupVSZxX950rLeh3A4AV8WS6tPeGQ5TQnIDCFbbte0X95Vz6QddBG
Xjev2fmp4lNNV/8dxukHirGs2yGnT1yp1msuKzuV2vjrfIhZPqZ3T9mOv77csOZ+9ZQ7xz7q/Mgz
q6KYdUUaChP2SwiwuRVCXZWxpnAuONUufLo0gI1riJ3/bFPvqHVeqN8c4cAV9XGwNzDlXcwURrXc
FUQU+VPKvPAkrvXr0ZXp2quGo9tweR6o2M6gHXjB6wHs7DTnnMIJpkg4TNgO5WTZ5BOdwdabUVQm
e+N1HqY+LbjmcuPHrHEabeRUcNgToT9rZuzU4Oy+tuDPbR5GQrgdO/RKatZ5x3Nt0j7iymdjL+Yf
l+BQ9eweV7Dh4KuShCYQXx32RtkHKAoPG/c+/4pJHB3RZYsGiYCTD6y0Cnh2C940wZUltrLVvv5m
bAShLF5LuGfr1KTj0VJIp93Yic32QJJB4Yf7bRRZV8bk7wdMBxUC6MRv0rcToY090g50RS5AuaHN
kMyUYWYr3SD8GIgDo1ZOTtC7gUrAu2uGCZUFDZ7/QOz5XndWCVe2ZCq//HI84GzLc+k1Bug6QqRC
kunUX0IpESrWWASF2rLtM4AeRP2gR7t5LtJ2icfsdFd27pIqnCzFrUuOhXnnSmimTonPGPYifhgf
l/kMdUfc0/EQbtFN7mFRXJ0PGy7SJG3qytOUHjgQzvkCWccPxXl5lebnqYeRt6vmgdHii7H525qm
TfXnR8XgxRr3Q//o9+oAaBrCVEln3F3vpziB6DPkkS6AhIdVkNiwT+/nKN3MtDaWsGaMgagsZb+v
WnRn/dp0DvzcOHe3mUnQBUgLur9iDxrtBOZOdpqovQ3if3WQj2szORB9HhPYFLIL6bpLZGqdfJSg
sqx5+J59eefyBdhplqIuk++PX5s5XKwQxefdfAm/gPj/2PQ20A2ZPOJIx02y1xAZJgfdpcnUbOb1
0fFYky3za/T6AKIMN3s6+IIWDUWMNXh2wokPSq1LM/XcIsYks/CpkgBo9RF3obB9ycqvGKeMmGSB
5sFiDVcMIa8wLmYltNoRDEjEcgNQlzbsbiHqEAKRqA0bPrrCnZvqOaK/MiH3gMqulRrlbgPQDAe3
tx80FYIK+pr1H+gB60VV/d2Bw1Aglz3TmzVDIajXmzmUNO+PLdvtGqIXG7bkK+3XcVEtvCgUcPYM
BlIWCqrhiOZeujPEKTM01XmjiffJArkIXvcN+lk8PBPox2LZsFDYdwMO/obigGs594dCxLdalAmq
gxcBkwTzH4MSC8WGFoH5scp6FHX1cq+DS9+xk8bqdKIGzCPpFOY1Hm0jqwbiUCp2vzbV0fwhAkyl
apWPVejDs0HsfqvIRxtEVAUZ9i3NtNl7PRoT8AfAO06g6sbYWYY9gbOmdAJt3/K6uw6PLPiTrlx3
6SruJnzNA37N4fH8JRsuUN9tLLpr0LrW5ZkV5Cs5FAuiRcOaNnBTdoIR14CmV7UyK/fnQ0Qex8+K
YC1gDjSGhluy1dhSZrC6J+TOxKhRn+4wus0nzuL9GUz1C3eAwm9/7TBBNhB0mJqDrMxE7WyEilD4
4M/shUakEAjq0N0JF8vZbEldwZ88YPSbSYoCY5CjVGsIhZmA54M9UcsCv3Iu2DfKc6qxOuebBt1q
izQCQ8BgxBPSoGxDUsYnuq44SvDRsXXFokAKsHE5CmeiziZ2e0F3UZID9dD68tPJ/Tnw0mvCsvVz
7uZdZAZFEoVWyFD74OjjD6YjrdyQGeuJN3Wnmln/M5q83U48F57A4sKYIHvhWKg8yl1hmtfeGKNi
Iz393R82DP+5WDWqNXIjaex7d0oxu35SXhyhLV/tgiu1igrGpgFgFi+DltXF4i8oDxxU6ZK0gnAH
lp7jHIJ0mSJ5RPZ0uErqizks/h5ydTgpv72xDWk6p/5A+liGftbKjubieB84MLomCXpf4Oj4i+q8
3yyEd5VF+k59QLTqm8uyaQNhDlcqxaiCulzDEM1nvm1+BXyjcxRCmCi4GfvnQF3xwrK8+UaJteoV
2Buq6LxOgVrwFOhkMJqAPGhv9WPiB4wUozweO3EcAEcs+u+ZGVAakRuY6hq1dO/DVj6a5PtQZgZb
a7gVPbo/DqZC9/DMt/ww5380wLy5nh3qHdOgOxXAwiw/zY0k3AGhq3+CCmsH5P54Jer8Dyk/PKnu
h1xqrCnb4WdkhE/LeI0zt4Zq+0GomviV0t8j0dUOFvIcU/Mf7ZX4YY0VRbDuRFCXP9o26PZ7lSXB
TxZI7YA5UWQS7UhcXIsFS2Lpi9nkdjgRVjiWqWgHVCAnoM1mJSW+3sEZxeA5f7KwnXCDpiAj/GuH
zoaLbuNOhALARx5CPvFKV8C6RR7aYXtFBtJAFPLXs1sAGoBN/AfTXZiJtF/sfXzc3IZr9rM+oua9
sjPMGdc7yGtpSH0KbmvUFgtL0BJhHz2sinlwRvUapl+LuNJgXUL77BfpWItceBpsINPm6zKdIkDZ
mxl+QYikYsVZiVaTxGgMLMM8kkUH8BApghjgt4v5bI1qKRNB0NQPHOIWBP0NrlzEii81WhFmVgZ+
h02Oy9vneHKd/EwcwdTZwZrliGGxtfKjgfq6P0+yJ6MWX5alvA8pUCvEb96cwA5xpCFoCq9uX8gi
H978SycgsMKeo9Zqyqgki9xd1hLwKVWE1z6aOWWU3kjNYt6hTWFO5j3ABSbLyFpYhLpZ35bdyZMI
6R6Bmu+Vj9wgAyxDTdZfS29v2iHRVel3Wpcw4/ePeaAEUJwGuDx2Kx9TG+u48L+K0lDl+BfCh1Hu
YeBRxlz1oNQD/FabQuQ1BjRPrXt6TTkxyDlU9a3tx/Q/nSISV2DW4KjrOGzlSWLXA/x64pUomUSe
W7C9pT3p7UHxYhz3JtJRLUk/mV9dZyPjvTNy2ku35UsVKTtHaDGTSH5WW5CXyBOfNDuso0yv7zTN
Zn8Pa+KSAp2EqBTIGmf9oHX78YzBHcsfQntXOK+z4fGEGVQumY/pVX+W+FWRV4q871CNfki/VJrP
IMboWOJpHX1rpSI41J8KZembnXWqdEyIXseCgEv0XSK3c3MuxZGHmQuTHK4+NYJdBpv1L8so+M7G
uAke5pPE+JOaz+7EqLAUw+bWPG4nmb0nfY1a93bv74An30ZgwyjgnJhru2i6injLUkYVkCVxcNIu
Rcl+E6+yDSZRA5at+J6fNOcJ8caU037XOp6s/JBJYhqmRV6t9fHecFP1nfEvipTyXvZ65iRAEqZr
G176M1tDV8jbopEzGS8qm5qfYurN1kiIKq6esL+cO9dSvRv0ui8hRhDQvgW6xB0XptwuybBV+Nyj
m5WWcOlqk5EY7PqTgE0gYKt8gaC79NppKRKPcbhINyaiByAAlikVnA4vTKu1lR3diPiNubIi8Uho
iXU3oqzZU905lcW/KNu1H1yX/dEeQE3EWQ+MIawNSNgECULbnrxQT4cOvt3EBe+QE0+Ek/xbBFFO
pZoKYlYKbSjN0aIwwsANnEurIchHSNVnwsdF/1oMO01GMQ//Qt1Tw/HKyrIZVCKZ6trVPxKgABna
T81blnOPFHftZa3GScNR07DH9JokQQ/Z1plx18Q27wUQStHK59Bc0/7o5Em9WEc/TolvHw8+EQr4
DcqQxT/HeHwr578WgN6O+PMa+2rI+MQe2jLaDklXZU0/1O9VXgyUpac+/CeoEXudyVKmSdP5B4Wc
lBLz8rx9UOyRATci0vbJnlNLhHEv1CmnpkPw3zUJNb3/X//uMcLvOMLWVgI3UH9Obi4he+DNmGom
ftKcTFMgM0l03dRw2BRDnG/V9q0FTJuD9LlJih2GopLE4ZuCy6n2iepEUiIbnObClbuEbvbdt6ZV
0+aPE+0RLpUBGHXvJMuFyGO91HAt+DZ5Mxv0i9mEVVno/JoFytv0xdJ9VEuU+tgx17A2OfzDMCeB
l1/xmK84ghQKfW0M88aE/xL/VFJZPd3ifFQ1gzNCTENS/g4Lls0SjKjCwTlLehCIPq9XOEAxsqff
pEdRmRrTnm6ou0HLgIWzAKl/apWhR7O2UywHzOxxUGowob1mAJad4D+cTH6q1zP7SGZv6bVXKmQE
MFVQ7QAN8MfpnU09ABhAtNulLcxiWHZCcUMVJTjcE35GlXcdrhod+M9Q0dFpFODKhUL2fbyAXov7
OapEUgnvVHa9HPgZRnDah4eagGUd+um8oBxC0pG3yF6QyoeN/nDYwS+h+P0bvEb+3YruqWAKTM+G
99Tsf9tpOCN0sBCuRCF5eWAEKXccVPXCJFLGbOY1X3XLZSOAfMRjTccI9kJJEWK8k3shaFctN+T4
lAEflp+t1vPS2geQq0/mmN93TUU/dWCDCsYrb3aGCViwn0Rs0cub4fT9dbtWfp3KfMIcQl4uKjRT
ZCXEnQxSG4GbiMASpgSJdiFGyuqODjBgrMT1HgQWbLOujhvNFzxhe9Sr1VtKMP2WKS8Pc8hQu8rq
OiRPygLSXBwUdeEkLpCdWtDrNAD57Wgt/nZxI7KvayJ0Pv9rcV0IHmVjAllHN2itMWODk0f9VZn6
7zqkr4ZkvTWTSlYRAaQBizS3auzxntF6eZXdHJfRhbYMw/sxYOCkpC9VMQFaSiNJlbl9J/NA0j9J
+qzSFpwy81NYyQyFvnlviSG41pmw4Whbb3DsiRIUEYQy3tBh4dElUGnjVAorVHqDzANFINhth8Wh
8Z6VSrBJlQcUU+lqi577J6nCB8daYKyPgpM7FoZm4bUqeXZAdaHtDxJVnV7CL1AckdsaALlor4Qe
dIWSKkn3GjB4MOZ1wr+GfWF8q+mx8N3TSXV0gY/ict0PRZFKegMv1/ehW4J6rQRiH2BbgtsuSibZ
AOSQwqdoIRqcVJx+7gGH/i+A3300HxLtkUXsRuM9OezahdQNAJd/TjVLq1x+RXFPhup3f7A9Lymf
dHv0M3AJK9ECX1mRe08rrnto9KXqRWS0pLlZ7+qsI8xTihDOH6wzZZ8mTvB1K3KinRFuI4iQsJus
Jb5iB/6tsurMNJz9yNxzASVWhjv7B7ISmaLD5UwdT1BHwVQ5EHMAo5Wh71rNKtiUl+Rj+J3+wqIs
v7mJoNIuV1I3pu/igrG8C91c6MNdYbpehKsFMGWE4PaUf3sd6VdBGvFmrvTUVbWnA25bsAXjG4Nq
QfdkDMDi3rS8eRwRmaDG3nNdjH6YtNz5Oxt4miZx2971Lmv/yPKhMI/2YQGps+rh1B8JiYPpi6PO
yibUfsymQ4rjMevnxigff55fULVSrOlGzKURd+BoOTEXF49s4rAM8BzUcvjKX0mcxN2paC1ifLKM
GxImZJSIMrcbhitokmrJ/1ihbspmlTclnd3voBSkXOJwVcFVfzpCyzfGve8uSXki6coHUjbj45Ng
3aaTEyUEn1P4i6Wx0MsFKbZGKHusGW84FCCqN03TwVWUSm3e1icM6ChcBkZYl0FoZ67dgPTGnCdm
5eX5ZjX5azXNMs5PGNjLmoL2czV+KAWWwMqLO+TfClQxDj00Voi0HfgxxI1AiGrgMj2sHbbTd2EH
QNRAvki/rylccoVXh0r060j0OabpZxrpOXXy6fax2/3HXBqtMhYXJf2tpIalng34yzVYcVMs3EES
eX/HL5k+CHVv/gEG7R0tS7lNR8U4kYhhH0h4b1fjUHA1qF6PFafwy+lr5Jltl3Zy2OZK0kGGaLby
h61gER6XMuLwBT7lc3Nt4YCoR/xfp4yxYuQH6k86Rvqz0vR2hM8qpTGnIQwoGJrH1EZvpQJgT5Aq
BkVrTPhxQLB49nx23bWEnVtUM16QnVZv2qVdJuOSu4OVBELNjMOEux1zYo1C+fYBlWdXOPulc5IL
U2c2TzJNUrhyjUMjarLSyJG4tiEyoA+iuLNqRXMWe5YLw+HRdZ6UzUzOKcutqx0Bw2lQleTHNkmQ
201VMe7gdPBX15e9GmEU8l1mfBGMfpSxa82kP1ldgOlJV7Pud47pEc8J4rnbjTSCvq0q19gDvGh1
2YH2QoRhg0knAQFUHONoB7A/BiAZ+hYs54lUdaCuN4i/MiOHjR+mkEsI8cXO4sH/eF16MDnZ6vBI
PgSqB8JaopYJxgOEvh3Z3t7MykHa7Cl7WF78Yy5FmyzVxENtEVbuapuGK+vSAL2G3FeiFafJdno0
YHb2U9AxMIxGpWvQI1XGVWd36nEO0AyMQr/ja1A0SvkdfWYtB97aC32L4tvZJrz8U19rGvWoqLuv
g42NQDdXT85mvBlaWWWJVjDF0rFa2vyyUVvOlNqJuGOiT6AO0Hgl2COFBBWlUSWBhbnbxKsf604T
Pn3+Ftj7dRJvdi59g3UgAQinfc4Hp1yr50MlSSUr8mUJ0KZ3T2huPj+g4ErhXzs0Hc2xAi/PmtX8
UaXCzSoUrlA0V4+6KtSrgpgkNJcoeAS2+3qO/zIVIk9nQySGe6o2AYCKbr040S8yQn+bCZFgviEH
p0aS8irkwJVOELYt6VUsqQjQboRCu11GEiGVRggjicjms14wGDCvo72ybtY0Zf9ryxd3QOrxRv8K
TtMoK2O+lnG7rn3jGAW9g1effDTDVz7POFYToijE6gr1pujAS3RTb5D9TIaAX93AcB7VUVxNHHP0
BdHk/XksErrinY32vdLcIgdcPLkkME8QPTorgEZVrhnQcDrK9IZwGyUIMzCpyhX1GPT6I3pyGHRe
zVhio7086NwbcoLwWgplIqCN+3o98kxF3/CwOiYCSbtxDLdyoltQWc22d3YvbUhGi/A2ObKrAmmw
S10MkvQCyKTV2fDFWzvxIIPp3f1PPda/LX/Qc8TISoxjWaL0HaBdU4GFLeaVWemhoomlCagyrDYH
KW9dB+g0v//hFWTjR0Ostey0Pbbu8w1YQJF4VdVul7hUiFlhcVKLMRacDQxt2lZ3pvXpB8K+Emed
bJh7Wtqbhp2ikDMtij4PoUO7ow5U/ZACGAGhgwtdOoIo6e2YWgdivWrYeCXUP5lFcEbxvds5wqgy
3rtndMVVJmM7a5gF+XgciJBh8CEvBMokgIwF06veW+FIoHX/n9juRafJihOdYcxwhExq8Xiai06u
eusIetb0sSqu/SDDE0EQfhnqGacuopZI7AXvKnNaG6prPP0YEjcxYqhOuAv486We1kIHwmP7IGO9
FFRvpX8Vczb0i+ykzcItwOSmWdlnN6IjdlYLNTF7mex02hV+pRWBGo95wbHtfZ2+hDLiG5j9zObJ
nkhE/Mk7wlzDPx+i/DWyc9z89oGTw2A1gQw3DK4w1vkuBfzwrpTYYpgiQkR9wTjBfboFbifDtuYh
aYbnCcx/YWdCKXNVt0ogCEZcN9DNge7KOZQ/GHLcdcZUUFW8McqfA1H73Eh5M8z7nZIeV/rZ9E/N
/MXjtcivUTMox81f4P2xqJhhNTXeOJEKxHA2AT24hYSTG7NMTAINsQdYlfRZv1C8aKx2ZCi2dF6M
u0poa2Ii2kS62XHyi0r22JHSWQ1ai9/T288IilB2jo9F3ebw39J3W4ZMOP+NPeZzPsDVptfDzhFf
WqeO/Z3B2pxe1fIAoJeEA7tMcg/F01LfJm8IooP/DshzlLMoU5Zw/JrQOT8AIbWI8+vQN+sisYuF
bWuc3JjjITsE/QVFmY2ku/70XZbjxf7iLAn3sJbQnHnkUfvGCNfyn5XNirMiMj4SWF5uUNnOJ5dB
acMca1rOoxyd7Y012qDklq3RpRig2LS8h5S5T5bLW2/K8tYrzoa9MgpAER+TKAcgVtKOdUwfOaJ2
yXhwUiUpgp0LruFKke7ahDoK3yWtaR28NjlgwIkuvtey+fgeJseVevD4/4lVC5bBSaiBb8M6YhDC
+gsAuUIgkbWtLx5jKJ59TFaYSLQHm2kguRqBv4mPv7/mwrPsYLY1hy5xNvIKRcqjGOcKMYraTI72
c7K0iIxTcYvTcmXHqzwwU1L0gwLBs/H59DvvjBwLJLW4THQJaFTiiI0zmSEWLO6ltx8S2bdfeHwM
B0RulLjB+UkA44sqCNs4ztaCuLbZwRhgO0tD76TDGys769upgH+lVRMhA3rvDrNgMO90AEIcQBYk
dY+f4D/57PgZ3NzEs6wdoYhKtwf/DmqxAEzTj25Oeu6LrMnihO26DC0CbyWu2Ld1wPZvFc1z+z0A
zl7c95ueKFR6URDAGHI1dqegre2dn6gS1YnRY2ztGExrYwp7euQtE0342wu5hrxuOtt2kt/TEK/+
dtA/cZplFw6t2Q7LfxuJeEv6WS6n1PcRe+vjSPU6o6PNvcvm2aO2wzMUz9s9Ea2cRbkhRdvkdMIe
Q33GqGH9PDiC0V8+RBQQxLWqSRMHz6T1xIH2cyhhLdLbss+EYDprCpd5iKaif5lIEKOg3EShDEwC
0aM4J2aXj/n2C186XDGKt8QVsV0V386nurjhwAoGSppmeEYjYBjRTrmyu/SpnJl4iY3ryoh6siTF
j/gw2mX7LY/cTqmW/Uo19YyDIq8JXoc/oAKlz0rquD4CsuuRlDH+fBiwNMENpURTlbPpuEzRLVOL
XXgS5a3nItjsbxD4mZd5cZMJ+Te9F/w0HWensDEUa4vYzqw8S/q7Iu+J0nTIhgpizgsg5oKbJi6V
r/WpCerFg3suq5y8TFe+C9KiYlVa+0v9nM3zpdjJ1ZVvsa3SHcy7Y9TjWlLqCy0WF9IJ7fkkr+Js
pNT8xoVfxCa4Kp0jfSmv5Io7qHLcL0OzBuQp4P6nVxUOp3Q7ziPzRGIgqJ3eFnWEoW+ugSa3Xkcf
RPn9YI5BzhXJ0AcXmaYofnJ8B/ChMf3cxPMutWdl23hINZ/uUEOzafEPp2DMAKamCynB+Z3ZUx5c
M8Pz0fk05wd4CYvy5NtEX9RU5WVzRbGHB/qs4onBkZdnnT2TwQ3LJqoC6YhFaDbKvJsVPdCEpqEl
LssL4Njp59vOT6ASI+A+gLv1vjxWWzVsjhPiiZR19pboVpageyMxRaW4pEmXsqRpadf/4mYWMjfD
do+lqG0GHAjDGwXVFY8lk4YmhwAX/ycm285j4AvXehRzfSQjnifjJ65sgLaoNUN0YNPXxc8vMfA5
53c8XO6TOgHh4xRfalcc6TYu+MpLg6CUE2LFWoIQHrJneAFiwporpMYA7R+OAcgWUwT+R1p3CNyh
Up42F8OYQk4vK/G9j2fjjPAGHW60BQ5nAAlaJP1HfQQph/jzhdfZe83MXyKNPEl/M2hw05x78rDl
rIlxMW9Vc+EirKvZE6QZTI8le860xMlIqMt6eWtMhFXrghBnzHSIAfdJexGstQFae+XGChe6biiw
YxD6BAWu9iCuSIckBCKXGnNtr+CygkLKEHdoQozYlc294r+HqBrGzsQvmOCnTcfYDEueBhNM71XT
oYgo9+aRhdeTW91GyU0Fszyd7Z5Nslh9MZB0x9tcZ+D+i8i5y4ImQhOfZdZ7lbdxrASTkrVFs1m6
KuZkapB9ahNtkodwJI0WbFrx09anDnx2TUL8MfcFJb52zIgkup1nIKwQhko8EK0oheJwpEdnGVL3
yNCFfTCaWYZn2Ix5Ce5XPb8bTSu23xPKECClI9FggsEo3GBmS030YOvSE9QKQgrbqfzkQaYi92Ii
k3xS8/m8ZDCcf/gi083oB6FAHHqhF0DMHjRVxZB7HnJ6EWX1K0f6Y68F2404y45NL3SQ6ZGCb3OT
YI09yzBbPgfHv73L1G3jgf4bfFnURv2biKNXEaK5DRfNG86OdQmMnFUT3Aw1ESLKm+P+SdR1ZvFP
UcNLg8AL79hnNM7YnZqoxSn9HZUkPZYBbsdvBQhVwSfin7kvYLQqCRgP09SgJU8FfMOTJlG4nkaI
TPSyaJ9RR8OQY2NwKE0PyMpo33nHPK9e+cbWB6S8qHoEQt5zgIjMxJB8Zhxwr3sKTLYnTPaUmxaH
Rczl9i8BgbZRi9b62bbYFKKRFg3/VOoNEeAF6pqnMCr7Mt+NACr0CukkZwFVMMlHltQuvfSDz4EB
KXDP3/8RRoa7UJ3R8ILx2O65s+hnf912OBfMTsFQrsaWsPBlfNUYbt/N/XSefZNUDfoAVPpwwHGu
LeTqnRSTPVqC9cFkdeIaTBoWlkNhEq17n0y07ePTMnywTdhlFMPtqlfqoadyrnCX2htmh4cUl6zb
4l/bnCinvZUuV5PrlkD2pqIhcPo/dvkUSxF4pWe/0OUlfG1MkfPufA5EdoU/refvvhD+e8uu7tWK
K841uNanB99KTczZ0oBTQTMbM6qiKfYGuIKGEf9VM2r8J7rnqeTmXGrlgIi31hTz2ei2vyUsP4UG
ajZXHxuJeHf3/A5xdFWVt3FB/YaBWOmjYpcf7Vee8D139teyNN9lDA2YVZI+haH3zaha19YxstBM
/ijErt8/7cGFTHO7ki7Ofy/nMUz8WLY74TQktFuS0Ysxt7KDpJ/ejE8WOMroWi9rlR4c0qqHoQFn
h68ElSu9tm1IXM93QqoGgofudDN/kr6AyRnZQLAqnbebkpxO/ozar1fwX0627VdXdV9YGT2l3JBP
c13HJRBIClIYrlk6plZb8oGP5suTAzA+GgxlQVdPRKb/Ox7UPS+BL+WjmWOUdH4VLna4OjijONrJ
mv4htu9zYO8pVB+C3pmV0DFpDnGZGsBnQoK/8cV4gPIpbvzMRhm7YBqttXyJRdXTy9mg3uGiG0TA
rSuJ42NhHo9tKTlKlxzwhiyYmP4/nuFWjCqZm3RuaTVh5PIGbZPGmNHjyujjGBXoZUg7pjgauKB5
YIcTvvGGZrgiNy2+iJCL5KHcmciAx8ZoSwMKEIeEbMTBUUCcCFnJQzgp+BAEUA4FEbeDGs2/pR8N
IBtek2eaneMq3XYJhxbkLMfZccKghK1TqUDwjjo1mUIEMLWNIDULzvejy0xIBNFwEf7UHmNIF6N4
o2mHMwBC6kxIyAUnFtTveadtyL0IQeEbwaGOhMSaJuCaq0E62SccAGhqiUCVo16PK0qce1JhJw6r
4wQDV8lhmI9o9drP4aZtJsLzEiP6mJdr5Fq+Lng537PZEmadsQLPgek4e9sYGiwadhUX0XUqQ6Sg
8Y2Yg8VolFHI7tID74ssS89BmfdXDyrhGZji93LNTIeFjrYLyHMZTY8jB8eNhP1UrhlVMvTVBmz5
tJA5d7aCsTG+bhJbFv99/H8LRiGdEIQpjykSQtHxnM4VzX54kOxaTRAY6IUmiWIw2Xm/nW1nsmgC
D0sLw8tSTZmSi8EDQUdR8yI+wt7T3S1IuJC9FZs+WopG6ASz2eNMeWMMfxkdBKgB4tHvC8XPYatR
NYH0yW0liDyxF1hJGOru3G/qrHiZ2ZI0w4lI3VZ32hMyNWSaHUNlRc7VfRuRX2OQdL4CrdVKlkVa
7uW+lNCBAcwJTqRIodk/Mw3WvoWVoj0CYFygJfpDps7qQ4Z+XUVMkBGKwDM1hYS4yuEOa5WHmQVu
PoKbe/OrMCx9NEfolL40r/4VLdNEZDDKEYM59TkFZTr7QQTakvtu4BxZ5PNdDkQoGVUy13/8Chju
/3DE3Om95IkXxmv8y4Vya0yoCe6UUXJFKgYoGZrqLs+g2jNFoeWqTm9hAdPOirSBhM4SR9ZgCSUx
r5ji3vekyRnULw87OvHdGGF796iy6xwLxpSnqK1luPCfPwp880sgsgLv9Ps80wSUJMRK7lanhwGl
uKeQynA5Ifhn4y2/EB4mqgIoBH2/lVRh87M3rUMz+6rPs8JSexzhEIq/LnuhPIQz8o0paHGSBE0Q
e9a5TIaH05sdEFjDbGpuDpIn0bKSddp4n+9z76Va2JdJyceaTsRaOE/g0MpL+zIw1dEVErRzzmRb
ehryLsE4m3S6pupNEsbU1WcU8H+x8NZctmeQIYBX8h+hGRMR5OiOMd3iKnMey3vmQEGcaWXsQMSh
qAgLjsF4BbxRJ74Hd6f6VGvWS5f9DMTfm5Bp6yYbKX5GbG4vlMYnZ6d4NMCzGMkKlVKEdAkGQzpx
HUt0fIHG+ER0F15+uAPo/spZCLkbosqDYx7I6zTEM1SyI9x7DOS3CPgI3KmH6m+hWMEdibsO+SSV
GYZFAgtp0DamxY9KUwgcIpyXM2j1Jy5bu24CpouhltVZbnY1/2cnBKMa2+9KmCnccItnvoo15gdO
cI23meUVbyNDoTipR5Bak1YhDFHu6fgUT1ITlGrZJ5SCglou//p63TdjBN1Pb5TovTyN7fRYkQ0h
9prenMmXKYalgJ4TouxPp4JgDWFmAVTEaZ3vdERULDtu/gqbEuHmeuF4FJPtVkzB14wIuYEXsVyU
g3Wo7Z3FX35xYGbqZo5QTn4xxD1jqqWQzg7DNZZzBMo7iaHSNb++FxVHzsAwRgu5aol7qUE1E8c4
ulG85V5bfLRp8WhknkWNcHFz6I+7fQDE5YM8D5Vy2Md2HkWDvpWu1bDSxG0YBj8YGi0pB3OZ5WUd
p2zW9Z2oftnXdDKf+CfNfejA2gT7lES2B92eI1iw5veBL4wGiY4TxvuQ/MjZaM/fOPhxmE4Ptokx
wqnhyVefnuTiMFo7HUIEYSMPRTtPzGhtXCEqE1rFC36hyz9IIhUWq1KSUua18yMWLP2mnFC098zE
OgrnXQ3Z+wfQHSJKznMF5H8ItuWGaGYmB8enW5gTiL++jfTkDvuS1a/lCRMlW7M3p4JVx4gL5kRL
onksUTrEh/S5Ho2+OPvY+ibghRQ+sy9X7KbITJzTkh58O1jKfs5jnqv7umZ8mz7SIKMrsLgp8NpD
r658ZWOsLoYh9LXSIaEmE4efaaSXxsa5gxY7nF3xwPVa8icGKKZsxsRT411Vb4az2NCDmd5IU3ON
8ukX2LYfIrofW/je6HGTA4L0n6JMPoNwRAv6rLebLxL3wa2anTTkQQUdRHWnFtuWUPGn1DP41Hqd
p851teUAgT0cPkFApQlHAQz+nneKex/9qoz2APjZahftIIkKwZiYJjPSVIAtWrxrLxBWluGIqipu
gUw7CtYhKPEO50s6J5DT31Atq+kQOP4Ovxms6BqTeOONTU6uRArX9eBkgoKV/FMfK5xHquL1bmu/
O6Mq0FglQD/nuph5rWuGJabk852Uh/3rPM47tqLyj9IscH1w9Bk70WJtcxT4o9CcELqHH6m2nNTy
njArOya3u3l5z/oNju+BpULhxAoHqhAB5e4zn1mdBN+hGGM2eKx8A23f2dRAT73vtzG1wOKOu8/S
zyiljndFlzP5+UQ5eiNaG/q67KRmF7sL3aszu3XRaTsy4MtamqFJS3MGBic8s4dgqEE5xmZKfX1w
4Mgq7VHaEm3zKO1To1ezmNir99eq9d8CrqTdlrMM+aZvDMZoUFlbFY0A/pXVBDsIvI3LjvrPkHht
4M+VT6KSPPvsOKtDov8LJ2pjniaxNAxsoqaR6Wiu1b/UA1gOcMsuzQFlOe4RcW/yguJ4X39Ucw40
/c4pOgcGoQF5MctAtJ2Ht/72YSskWzrj+YlKlIcCko82u3qZSRNUlauEMbzDdQRBhDxbghq3vo7Q
//vVpoptq3MsKjgpWpKHHVxMDHJHrHh2umVGhi4gBlouijnX9H8D5kL4Xotwd+BV2oVtKIuRCZsT
mfiSVCxlGAWAWmGv9E+VKXToGeK266KKlGoLCbFVHixd60o7FTd+/a8twlxaSW31pOjqf3xjGJi2
NwYTBEJEPWfNOCi9moJB8hJZC3YsVZ6iN+udJX5gRSdx8ud4RpQNteeeuBtHbP1bMxOxmliUkoaj
r5R4HzMemQpnqLBeHJLrrho4nr/BCbuatjx8CY6hGZC+Sgq4iy0ffeLbTxwmQe67TBUeN3sCT4De
CIK0yAsDL7bAYYaGnqAhkA/d9TUrtIQaiOY3IvONDexPDn2ZtAkDnD+yfL8d/Gk7zVSQYhvag9ag
IK/fY64QmPPHXi35JnMLPLKlQBFDDtMMnr8r3T3RAxrfsiGBDHr3kh++sZf0i19mRyiP5QwAnTwO
7COa0TigRq4jmUtn3zVqbl59IJ4qYIez44w7w66P1shW2WcJawoE+Y1DEG04nJ5OJWHZdk2NRyYc
scs1TJ8bVnnvLMxmD0EykfYQbgu+aXXidZBeL8Ci5CLp+44Kk6qcZxJbTUUBACPqLVOopGuCmfIa
/r9LGgoMrYPdjM0o3J80KWGjvqtVoGXxSxzUvKfbbkkx+4xuruTmLUDw+kzKgeQmhwfasdXtFw+w
HzuY9sNzX5GYA3RN1MjT1l6W4/hsVDKFbQyS2faP/qEjjm5xnZ89FzCBAkSDKVU+XnsIaLBpVSQL
UX4FDIKv+WZJFY+ckUYCQNh85kKElMprtKsegbY2BjWFzua7igS/gQh9WZCFEY+IzJqrUhX53LWe
pwOF9+y9uaZ5BTr08aaqkBKVf6pwefQBsElUhVViJOpvQouLNAPnXm5GBpdKG+WQhj/jhePgIqXd
5QbUVv5xJTBoaha0wvjHDxyCcB1GAbIfrnHaubdSqKog0mFJMrua+vmYJXag1jBIF8i01q12cEh7
rbAbbWERAJf/BM5HKXIDqKWi6KXaMUJcGV6yLGOdnk2cCl3d9n88e9SXlQXIw2rBaWmYco30sfsK
NAtjahEXNcSvU/qmALDiEYHbGIOOJJwDGQELf8I8lZqJGqIcUSz7bHSleAEqZ9M751IT3tpNJuaH
bUa7pI551gxORZl1kdi5P/tU8VRTrHiD3GBWT3eSnGGhBOb9k9fMgxmdYD1MJvcoyKYPiQYNwrF4
gx+DBC10yc/HhQex9XFv5N2zEtm51Pd1S9wn4FjZrU3+S7ucA5mWD7wZ9fjdILYqLiM6XMbFVjXH
IbT94knaaXB7mLhohCZCRJK9enMa826K/TsBUcO2tgJnWlewlJFqUTzJcxM3+qBgSrHEXOlB72Rk
g/tAybE/MUYeqDFRVU+v31leYsvdy6SZv52bryT8v/FseE7Dw8hxFoFQSxXxEvuijyHMCfn6El0v
dNLvEJkQFwNaVgB3b1xACTjOxnjPI9au3z27D3jnJKyGWFyIepKdPmXxHQeDRt8w8F0HPU6vmFTY
hCEOzlCLpuZn5/5Mb6KMypOP7of70ryCiahM35RRzVzCb/+NO/j2azaPYSDildxK0pu1ce411bEt
M5rADj7xTJRWGwofIgQ20uN+d35CtWk9XR3AV9SWV8B+u91ANCV1PqAkDiU1nbIbYkuQsNUwZRzt
U+Y2KPeYoX15lnPxoDk5HDv7SBtpfpazcTdYGFZB7UzqzFguWNDkRc2nHzrorYDeFjVm60bykc0z
MCvTSafk7zKJA3t0GIRbHW05usAf0ouC93/5e7HMeZh5rRE+119Q1V4b5ho/v4SHcyjmfdE7NIbT
JmqH5AYAEqbr1N93RNQ1zx3GbloiVoXIu5G8OPVTcQvftpy1c8KTZfQEVYXV0YENXNTrwn4Sb6HW
75EbCKV6dTXb8QnNe0baYPf5/g+26mtyx9wmcCjIJHAf3QvQQBYPZ7t+sES6SWKHb0PwNEiASEhn
QsRfd7xONSUcDx58n0NdQiuhD5V5SYkWONE2r7jJalkN1/n+M1kiroKwjdl4QhCHJV7eFGurDQUU
uHWIjZ+R6vcc6QirMEaXzo8kdyFcXPfKtpMNXWv/YRtXIluv5y3p310TpLk5IO0MLKyy5PNw4mz1
G5un2xFqAYcy2EDOChbw+96Xn7T0q6ZAUsl2uTqJMqLzucvFv1I44HKzXD+IWctSvbOkRIH+oX//
H1Z7lH+PDL+n9Xdc3K8NyaaIrhhKMTz/EUp9GhL9VqU2GipEisnvCprQsRzGREKbDE8MdfKFj+oH
fkJGh95+zWOMiiGc2RJt9m+sD6jM0cUY7rddja/6RBvm2/ANsBAQyeRW3/P94Y/04WWLS1G3nicx
PX4LzZ3F5CLkVtSDiYVPggIrWXoI4PaHy4BG/BHGzVSkt/a6IXHd2u+qlHHQJxlS2HRSxwD+aH73
OEmbcSKX5wV/Ns7kPQ92ClmgW61dMaU23bRwERgkapk29HK566J2mT95UHb/75iMjMFFFeo3zzfs
Ete0LIk5uL9/IYLtFkWpu6yEW/bP/Yvzm+EXNJpr8YIX47h6Ty+uGs4BMW8asvPIWov1Cdsi83tw
CjWJ7TzGz7HZUU9MtAzbZzwHibQtiEfHFmEzJoYuOYS9Gv16wWy10gEbjLW1+EwrkGDkrlZcqf8J
YL2G/GLqflzkS+i/aoOLYRAEnuqzp2R6GNKJQVzUaHzGTBHcxJMfbR4fNrXQaP+zTi/vgiEay8oX
mvkDRPt2+aLXxVadqac9qdC42DEZD3d5H9OgFEdNAXwPf49OF7Z6bG/Jp28+laU+D/02paYypE0I
jEohKispibKV6UynV1Z2plUNbGg6OAQrdkrrzWMr/Qosb+/DBAs5xsJHKs+bgLW/U09eYHsEvTC3
E9ctNdfAzmZvQ10UBMFQZ+ggJl0SYmwDJXoa5nyd/0C/g0ogXnU4z06Zxq9rdyiP1aBmf3rAvVRr
PIrq3Slu0jRccQbaZaVLOsqc2EbH48o+KhQhhceQ31kbc1f+aceCdTE2fvuHWp8x52j6N3sxXxyb
dz2t5oNyAie6FVZ1OxUUmNdmGc7cSiTiKx/QtgJOghuMNDH8s6cIsZmlUA+k20q2LvDg684VUysG
ANifg/3vXTzPtkE/0JV8vNe7P+H+yRP2UHdZ3qROptCPtaDxAzS2FJlXbmG9uDaXhvDQAwM6aZqo
WLWKQMm+0gsO2iup3cO93tH7QBEBrkaK7on2Tv/euXGHBuemHS0ojXJnvr81YYcwL6meX5kH+Axm
U243BXaj3x28AIh020xylC913VuAKYPETLAgm92fDg6ZVtZ2FzxJccLbndBAFt0HPbzqo+RaPPQs
EmAZ6VSBW2/lTK9E0t+nATJhsrNoAI2oq6RrCNNjpMDQn3Bv/VUh79YCXtYIOKvM8JZ6pczdSMWW
1lGvhjJuwI/ESdY9dfUyl6KyOBiz72W3wUstt3oS0pXZ+SedJwtdXxzLoJvg8GLnXxsgNe+E5oMm
LnaSI9oYhPRJ3rC7gVYgbXZjJG18+oqvbEMrIUVCAY7klAwNFwUJnrWgMMnWRGZ2teggiy35wjTH
QeUFY57iquOfn3HqOpCrW8dEe/WmbfDQK7Pv0i43ZBAo27ngr0yYqIfZ/jj21fR2hEoEpsYsVXDG
c4RCwn3dvM8mrLQ5IBVh8qFSBWILXRxuSR4wktirXUq3nn0wuFkKU3E1eP/KbIF/OKxns0bVV94G
cSANSD8Y/IDAT+lZG3YjZWdIn2/46MPw8oKeyOj57lTBB2D6p3Uh8w6/78Cs6jab5Cihv7+s0m1Q
qSaXG+NsEqEbMxaJ0QryHWC/qHlOCowuwpyCKajFYoyPlPyGBZs4ItP0qNdDwLOGndjvTiNakxFu
3yy0yA2Hgp0VUze8Q5vIrRpF/eypox0aPqfJIVDzrnvf06aHTxHhKT9HV9Rn4JmgNaD2Rbbr250l
i3UThO2RaIpZpr1a/ASmtRvxKIr3os9epf8fgI7V9y+D/+GR4BvIsyATiIjm0ZBfCFcu7cMHeLKN
Q+Dek0TTJDCenjrnPQir1l6hty2pj9F+vi1AAEMp7IpZES48QJOvRMJHZzlwd0inqsbY0eXTVOBY
okWQPI4zyhJaFZfQlM8JZztoI6kRLT9vRErWllaC4WU9qL+JBQ8Lu3awj66+wcY8JtjQ7a9mclGW
oROGNJ/Yqr6L4w5khQkdPoT3Ke1tcWq41xxeBsWf5zacCTvqmnLbsnJ82Owq5ge/VGEm8Ir1Nohm
FECFfzM1MMsL4oV6l2DltaRgFMr6nUC2hDCRul6Tejy+s7BgbFneoUwL+0W10j2JBp9K44p2MzD+
9wAJ1vcgcjtXZdYTN5QzwFg3UED0dFHxrSWTmdkghQRb0iEufp0RHqADj4KAG431+W0ApykWnSwg
QonvCfhJrvIvPg8iBsiRPp3E9oWW36kjF02fLItswZfdhtI0LL3QASAKQsf2bObwsQCyfSHLm28o
wTrCT6SU5kUe1ryYWTsYF700Tls3lggCUKpt4BGMte/zg0KZ7xViJ4UkoEU+GhiMe4f0hzzQcEdF
sc2d50394pCfVlymBt7T1XGAFHC8FqryjCb6dg71XwtzYsPAoSnaMM/A5gqYBQvzkCIV2EV50EpC
1uXC8rK79q8wg3yJZf1npa1pdvIljFwPK4DQs8Ig0YeV5NmIP+dl1kIbLbR+NnU7SixTc5pvlrns
71C61WUoXtuOj6g+fTz8wyQkMp/O2dWklzvSqleVlB9DrzuDBG9CastK+c3OlIbCc5UicS2KoE+A
S92n0dN4VHpcvok9nJb+JsC3fRUDLUzqKhuPrTy5j2ZTnKq8xeQW2M3BRpsVwNHHrI+88JpMb5xm
h9W08XqvkUL4wZadAnuM3U1J7BotX/kPxAsTKTFsyyOtot17kHTACv1OPa7hZfV4dMjkK+iFRjlM
XYW8At5Wod4bui7YLWTz0brd+skBlLlXX7mn6bU/OMzPgYL3zPEGqI44TMkVJkWarXXLuPzO75zV
dzWFyd/xUcmH3oHi1Waq7/6E4A3PTA5NZmwtitXmJdmaYMmbPH4ei5NwWkHXoyjOojlpej6afG++
QS1qmw1pFRpqr1a55LdpjzINDDdDHXl0YzRGppCSI6Mg8WNWGbjwmeT840ueHcO1/lhcBDiF38Mn
mMsh1w/OK9BueoxFs7YiMxVaQl/HusdeeLqY4weS+wrb6Mis+pyR98fGlm7vFJEEyZQxRDr3CHwH
dvoaav7kN4RnM6f+GEe5z37/0RSxTGh90tEADUpd3I641a0dQo/lbJq1fjS7lG9gE+j/lYK1Sp+F
Daabwr/jH8QEaNWlIlP64Qlvm/+PvfoQ8z1v3N/0xsukZ66gVBRqLVyP8O6kUnjUVKMkHkkA+wP3
nW2v/yaHpZaAH7M1L+AyszaC6EYetNykUL70qBVmiiNPm9JcEiApqOLFj2/XGdvbHBaybzUS3D2H
aqFd7DzZVNSPqDpFdMYfKCkWM5A4NjWuqxwunI0i33Qith5cTUl0+TDW2yptgs07KUn4L+em9smB
/jzk4XtAUX/BM5KhLklMDvxhghi5w8p/Ji2Yttw/DiOcNj/g0A3N6WrffQD77W7ZVgFiErGD/aL4
iwAhaRJLkL9jRFRt7CyRfS4y3CYmQKBDPaBB6m3FMciLSft3zc9MZ4JTTElSnni9Ig3BpACqWbVZ
HMe+GDyRRs/eccMeuFDvOZTsxyFlRKhuPVvfHY28+FPofqXjXe3NKDCKSM/N0Cp1JHTjQKgL7eYi
h2MbLKGuSlrp97nt63vraFdKiaxVTpp1YW0WqoogPBiXXlx+kHb7m+1hsp/Tff0ChDePi0vN1hVn
/l6KozLnwpvS/7DoM8Wzdcdq00y2DWW9LYFiojLfm9HSAzyDjI1VhHP/ciGqy1xE+wQUj7Oj6poD
iO+VaN2a/+K6LRrxVawUABOQwl8scBahSrEGm+/qhOMzFktpxkTqrW8mxbdPIqZ6c2L8R9W36c7g
ck9lCb3XpJYBA9ReGU6c/SjGZKXFG0HHORw6KbKgGQ7GUm/R0fdkjiMCTmQhzniNCy5GV/Oi7Ouq
nOfm8rzvSpSXnP+kHeDZkeaNWJKppfX0791LMeDuZlSron1u2Pd/nxs35Kb2hJesp3cRve+hAjWg
t6VfltrOsAYVg0MNXlPuh8rOVFr17T7nZg55/BIHC/OI2U/CCoG4syl1HKg2ZqJ7btpgCcb/+2v5
RwJIDOKfpY4QH6LM4Pl+QhrQwFaUB/48zIkitq8TYZXMVIersnSrYwCusRdHCPHS9a5DjEZ6HZnR
T7mSD//6lwmJcUEJf/zKgLmAWHYOeXp7AwsVY/E+7JOEDmVna4nx8qyzmmIpDffLH664vYmJvz/+
SavhVSi+Gif8kjA6ZXhN4J78Y4icW0y4YbIMMd2vJM+hY3b+RZqXQvA1kX0DK4UySgWD0+noErUQ
iXlSlYsMHGNscPydyGTgXtfC/u0y0t96WrMzZdBDvA5ZGGPoccRoDqXhRPFS/dvTQxg+EwHaU91L
yWG+pcVmePeZq938b93O5c8ZoexRmpSzuED0TRtSdQ2gCPASqoEtMuT0ILnlX/j/gotk7yJVhPwx
dVEVQntzPHCjpU06m5uHd3104RgmnUDd2FQts5IWpIvCHwU8hJNVfoti8qv6MDOuCk3YlqcbUvnN
tQkX49vw9lrX0Xnpgyckzgb0+wMc2p80S6osfE/2p/8xXUAr1jVOoAKeNKViK9EqL+3VmEdfBxo+
xLvNmWrX7B8g7qOn7uEvHg9ZmPN2NDFguBhbmjqesLeAa/mAP9CIAgesWHZIIwKOxmU5HmwDhzgZ
SZdPpBiNY0HbxmJ1t7P/tRRYFrFZ06SbulZIfpmxfAqgKKFciM+uc9yf5Xh00qGV2CED1dk+8KoC
c3eBCIEW2PhrPeltTMLnN2c+Pij8RdOKkV+CrjxUnpGPWo7FUBfjwqrKPA+ETNc70Cpf8+YEDMnt
KV7MRZaHzvMeBlL715x0DMxBCK0Ly5Tf6/zv/n5Y7Q8qrT7uRmMg8sv6/NB3Of11Iqo21jKBnTjr
CzOOeCLtmd4sncuwckGq4HrTagOQAH3jmJtD4gGaZyNTFy+IZSNibQ2KheXxwEzigBUkoRUmEXM9
P4gV/lN8iCGuy9HMKEF5pUWBDo0gRaHlgddnywlnWhBdOzqNhTN+pbgJy8AgFDWS6bgF4PNEEQsY
1zfCJ1xi5461B4CkUE8lhhtUZLN6bf075YHmferPSPSa8YC/PyQp+nW1T4yjWYJ5rbXzTjrGbl0y
ltofWdDJ5dzZfwnjCThuWWavnLRsBu0hDOGN3kxl1CamvP5OEL4EH18w8VSyPEMAPO8yKPlmRP4M
CVGL6rWoJcEkDchX34nyHVrigzNGg5vIF6vmMKfhTNYNhiwliUvDwnc8JkKAzTQmV4CKRuEdQwhB
LXFYSLLxTn1dBhv2ou6BxNdDaVK6ygn/DXBEG1cRaf1Y864Dy7dx1BmMSeKHs+fE1q2z9Z5vg7/e
5qf9Zd6A0OlAkST3RvMHaMiuimGoyXLVkV70juF9n254ftwdSd/DLTCNm3TkQ/kpNGyoF9qr4nxN
ZTZOCHss7fazvooJRoE8i+y/qfvsG7FPTDSYmH7hHYAwkW9hHtGJN6Rg8f5AeJTKApo6v/DV8T/n
QetIx61GZ1bpI2r/xDL0yGqGdGdjn+IKVP6YmGazgff2RPvdCQKEq62y4wTrsTcGcA4TGjCaeCED
pkjUKu+No73RQujWtpm0lIekbfxhD5oLeKcLD8NUKwuK3mLJR9HR/sU0AfwtqbXlrIxsu0wFcDeR
FwHsgGbSvYrCFh322RyoOjDTAHnoQAEGWWB89OBdREsWdS6o0Buqqf6wnE2ZlAUSp1ztkmyWSwM7
8gdQeQKpfrE7nvZUq6UMHhc6JKFe0uiz5NGDOxie0qugplFpe/4c0DMkstb2un3wRNVg1BU4BVoL
9qQIMEJ0pvftO5XA7y+Huvas2h7ngIBKNi4VAa8y9w6paTIY7RqD0cARkjP7STZGTxofXD1LuyRQ
GvrU2E+PgMVKMqykXWgi+2/Sct3dFudKj4pJ/jy38Sm8LQAQSICL0VvPuFeuzYvmwpyVTo0mN87s
f1dYd4YpMxxkBh+HsazLhFkm1ElbASBgzh8/cfY/1pmzO6vnpbzbaUDLhFMmF1nwJaVdUh7AxD49
lOJ8vY4QP1FfttkLIsoBh3y2al5MuV149vcNc2Sy5hJby1L5FFpl+nFgXYgbeneMbQOKkyg0IHkR
anga7qaMU8T0v47rpsSzJNxL6fxwRomBNK0y5RVX8L1sr6sR7u8jWUwO9/8QaAEPHresSgt2hy42
7sZxu4PBOy2LaRfJbApuNtJ1dOnA3fb6Uha/0+lclxg1mrk7lH1pMMZ57w2Nq52VK8MJrtU0HdE/
v6zg2Glm3KYzD/ybB12qpEBLPR2HGoUwH9Vfoi8lUOVIfdBYjDFHLWGaGBEy8HHLptbok0ZpNyMH
noRt0I5L2pAxbYZObzIs5vp+F7DjrNlSlcA+9JIYTsREHrqW2HcPefAPR3ZUhHvmv6gqbMh3As0b
dtZ3dpU3sbYb2rNAa1992PBVHSCvTvTHxGVerCTsBDoRRmiSK++3F7EuhoxNy+BBTbmoVuLFSBqX
Tr+85+WyvrPLWmjP6jpcJn5Sd1b9GgywtLLrY4fJZKM1855p7VwO0L5ZBlsAv/7tTQB8oMyfwl8s
13XzSN87oRfLOsowx3Yo7GMOPEBTYFs8Ejtq5WXVycMM9nS2yXTWw2OTiQStieKjm83+A1AJxVt2
pyqa/aGW/NhmRUgkSefut5A2LOG3cZm+yNAnovRi1JMm9CusLM1gWwPE7GyeihfVxpj+5vXT3ECY
L8kScYZnjKiMQESmciJ+tJuHwGE+RKsuBvApFQ8cGbdEpERScAS2Ts9WZjmzE/28vHp2HEOh3yCW
vO8u2A/xkGIR2cXETg/GTs1WRLP5n0h5JgzqshBMgnS/EC9JHYWdvT4cESenLneN+NkPmHEPB+UN
PCTIfSe/TwPwqIlb5uYlOkPyVDCLyrzQ882PqTDtO5G+Nixijq5ooMKRiDC0reJn6Agc0F5d3T56
sOTamA5gZSSJTecNBeMLQtInaBIkeEqGWGbmbCnZmT1LzA6yL26f996UokLlvLR1vzZ7Q197AAq4
QJztmkWGAV0MMnFr/VjnU24YLjkcFnvAupyczOZZoFX5t9SNoKGLHN6+Xd7F+HbF4Gb2ZjCVB4EM
+jSZvigH0udytZOVDC3TdIf1PkKR86/p61RRyxKOohCf7R7tl1xWPxH6kA2aavYjqqm1iPoGXxst
Ze/61xo5GzJl77xFfzyPfuS1enDQPckXqNKkA0QNxlhq08IZAlpV9bMnsIIY7XI8/X/kMNF5EDN6
4TOYFsuezxXtDIFImvw2PT+bvmj4Fr9RJwYNPB7CxebAteuOWD2IIdoDb1RSa/nSN5CJ52ecGMsb
Qni6X68g5P4yiZY+XgIlamigyK4LyKLQRPcwiVIt94Sl/cPP1BifLRj3f6ZaEqflj3fELtRU2ISt
Agb36AKxLIVTApH7jpCSppa69qyCCwrvwMRH9LLbm7xy+Sf5nsAxQOly2+BRiMPr/Vj/fNlkFJnY
BcxfDBE+QJA9XjGdzl/apgpfxvrTagH65tVKEyPMRPkPD5+NsJbkW3wfJI9r1GM56Gi87B8Vk0qa
tmV1BribgjD9snLi4TX8ISN78R6mo47vLsdFd97WALcIfNMvolFycoe2XM+nFLFu+oZzAW46Sg1S
nEo7A8Ge/ZMSKDmj1j0w/TAJVHtnyCmMnIz8W0puO168Ffcq/t6w3cxYQTtTqGlkAGf1ew91rrmo
N1fqCgcleCHv0s1udh8bv53JZxmADsXpXMkZ0l224+nzch1ODOrYjna/8lI+La2lN8izPj7UDdYA
r6f854+46grJ9nwAME0eXi3je5Iol/nlk/iUGBiwIf+l4rX4kdLz6ASh/TJ6cszq5mP1EmiDeEXH
C45LAl1Z3ZGTZge0byic/8WgDI5FtADNP1+Lpiee0fkP8Rk5/Bv8Pz8w3Gn1m6Doo8j15HWR/peh
11PcZ+crS0drrFomK/UhP1Vl4TueKf9Z63kPchw+gdSEb0hls/PWc0rKSqrVtDae98mSA/Bu7qoU
AjBaFk6bo/QcydCpTv8y9FcEgkCQK4K1LZo1zt/+PE+m35d3PELJSNJHAYqsP/9p+vs3Y8svWr+5
+CB5x3jC+wNkPO5wk5BrEwsLL7Tex9s5fAEeM0Ho1zmF2xeF9tf8Qy7GIRdxVBQsOY4HQNAOObLE
5Xy+kcog4fyiskmT5y6uD6MGyX5h6ZPo0Ugl06E0XSvkyujA4bQ8t8j6Xgp0AsS/SfGy2Q09zeUp
mtVVgnDGl9WelSlfydLsYWBvztwt4TGu1xqMvXLYCMpqvZ0zyVbp8EiLZ3SontlRU9OxTe1dZYkg
suvpsRHZmA1tMa9jVOglDrrJzizpaNBL9dXkLJhLM6lSimY/2Gg0H9+h1IRW+Qqqpcaxgy39Mr7K
W9YUMfkFe8lihO7fE/3WaaPA4SGyMVuaGtNHL23cnEZII0ugIVk8taE+FpoWIu+yXoyMJD0H5Fnv
HWaD/LCAeaU5JcNCjoLAylRU6ib2LGMsRZ5tOjBEjQ45bYrlkiM1ynPOD3qUzs05N5pVbHD5TsZG
fDOhx40p20VtW6e6eeBbCS+qyXVePBbw3KK7cQnDnC78qJJenAf6Mr+C4jKuIXJhKuP3r9ZZy2yv
nz9uvvEKWt0Iikc5wBC8k1F/AWp+J2+aioM3FyT/ZtQNfa28yedT0ukThCDG6WkzXjS5s6+SiA9L
zG6eBbbzC2Xy7wUQumUQUpCIDEn5qFyxTPrFOfNlseLpO5hDL258p8yi7Rstlzoh56yWbCgZbir9
sxxJzizH9irNBgHYVP8tB40yk2BHPnUiY8SU/eEhzxrU55oI7B6jHMYNipVj4QmQy/+fdmbC56Kn
uBY/O3KnYVU0qV6Jy+ud4oyiCFbEYY/FgccBjCYsmyeFEXbBLjuy6oBYBanbDhNrdYGPoCQAo0WP
oPO3ihmp6q4+/J8wo7SAD0JMsUJObpOIGooHuKljp7QWO4CRpfCKIcbm8ILqZLXWQvQ97fnYKz3I
CiOtHvcbFW4cgNvX+vDMSrS1wAJlWygS9SINEY/sqdJrx9JtnSBvpQ/pTqRMQmUmtXvj9o/0nnmt
6yt5siRe4OM0Q3b87ugW6/B1lJBYIgpE9p/V7PXBaF+lem11/BlfaaZ2rIPVNG5M8dAR2wYlSDLR
SHuDBo0bRbm/ErnCBkFpSYBIyUkiXT691XYBCga0u7WorbLAIQZTP6pBoroWpEsFF80mtfR4f4pg
PNjBvM++JFeaI4mDgGXZUSakN8ClUvrtrEjJxhKl1iQ9h+oRpRUznBdWCHPCd4xXrJKbXOhsrXyp
sFH4AS54RpKKgQllZnuEy5+ZqBgUvYK82rHhiNBsl+IRHGKsHAUYDZ34dFGJJEwM2YT4+YIOnuuA
mU7eULG+C/ynnA6/PoWXrA/TDbKywvvnpilIBk9ViI1krmnY0DBn61z8upUDYXjVaQ994n57kmfl
SQ4mCmiAQNvB/C+jm4jgNLcGGB5RzPNh44xyeF9/MiEeIskHjNzl4Kf5cJ6r8+kJtAwD910uVzL5
eKj26240P19PCFqRmIhH97IDwkfgMs2V7IH6LeNwOfpEsEPZF/cVAkg7tIbpWHz48r3chPBO+9RP
Lw9C4He6h8m1HT4WbRkqTzZ7Vtm4vSHs+1SO0Qx131kWjjAysx/uATbsl96HOxvhFBWXyihU3ys3
up9OOsU+aRWBekumX0tLz9L8IXX6HQWBUdaHsCJ2Zc//ldd+MAJHt0fS1QENsnsjQuDRhaRyJn+J
58Mx51A0PnFsyiPZtFolWKCT9tFeVDo65sfqxe1JqqekmxRwsAf0l+LmrdjEdUalI+EfuL1zklrf
CvTLNcAz+YL6/moriauDwUmQ+gbzWSZgaCLHr79X3aRn0XcJoCfPdbv0n3rTku6/b5ingnI32+yV
ahTkaGgiFwIpT4HqXy43SiyyDvd2XZ+7QnSZ8ZLmwfZyumLKY4AMIwMHR5x36HgRcdyaIKpajBNC
4jYWo3aaQuhQAvobjzwBCvI2wdlwxy9vaxV+tA5ZqMaiMEoLC0jvELFgOwBPVdFWF/ZQFCqH4zg0
ffHA2DdwSrRHaNbXi2NtGt9QWl9FxKPkKgTgE9Ygv9+VE2Pp8CtDQAD+ZZqXs7ZI1OBw/d7Visbr
buWFVuor0dq+se+l4Xhg7q7tCm0jWDH22XxCNhoPkDPlkC7TaLm+hZIK8djpTnwxk2sRoYKsSXMY
7ZLmL+GDTnEV0ISH6uWlxpLYWDeWIZ5gBayruSxFUpAUtu0huoQmAei8InOoYeXvpnWUxXyL5M25
CPF685UE7VKRrf02Lm09hCQHINf7YUEwZOfkyPxGfdXZeH1f5lCIpwT/dBVwBXjAIU35/koy/6Zi
5NhTPGQlqa84SPT+ReamUdYiqjL2v2sZ4Kc2tLuhWfPpI1+OvF2BX2UV6dI1Manu0xzHwayxOKUI
wL64tVS2qTKWuC68i4cu8GGf2hSg6v5hoKIN8RMFBW6cJiX6UJcCMERWiU1LsZWmykIYk2FkTUgd
37n5WEd4L4tkdfPh5z98qnoGOuKSPUcErPbINKhCyBLS3nOAypjWn1RgZxj+85lLwEjt2EoNo16Q
sRn/gwq9467AScGAWUe1CNCC8N8Y4tcjnHZclpE6gZ3MhRE2SbM9NRYB86je/Fa1b+MBe7AW4Gv5
ipU1/MaAP0X0GcGheom+vMiOAn+CjWr7WX9mWb89N6g5jUh0LcN0Tn751Qgn+IhR7Sm3Pw2HMZGv
hprQWtyz/mMaIJDxrfPiFFRcN4GD6egrxIYwMetF4zF0JM+e3UEhZXbed99PTN2nddWVcVU+Chhm
Z9+KeCMIeDNxpaV6dzLAmGCL5+TD89wOD9Pq9fDRSE841QyMqvsrN/l3u75YUyFBh89MWMTLaFL1
3gRg0hLL5hZ/Is7zAQ54mm9BdhPcRjkMLcmK76LIxdO5Sft+YbZlVpTE5sV0XMTjTXYi+xo6m+ga
clFJb5HjF/VkN5z0S/jW69R+pnJ6zEVIQhjETZ4HQAwUqXM93yWZVyUnYPNqy/3JDJ1on8MFEfBf
wMAkEmTMz83SvvyEIpZmO4DS9/T1xragKVkPFDEi/3Z2249ltvmcU07zSVcWK9PGPJ58b91b/I5d
mA3NJkvC3yy2huY/vmHq8fmwOr2bysshFWVV0dcpYBKyqkrLNINfgzYd66H0N6QPUtAVp1/G1jdK
bCOpRCfDYls9IzNmcsA0uQ3PJ9rJ8u0q02HbBqcVCTeNPbSxugGmgz58xCt+PrQjgN7XlYUxtwOg
3FfWAiHorxziM7SdfWRjvbQa+8jrivO6NxJ5GkEQrxqpqO8XSUwF8VsgYz48zmlPIOw3mzpG5yBj
P4aMx/WxkVjnGn2ypOsTLhYegRFIC4FwmVnjn8N01O9hIwktR/QsF1s/lpXqKTjmRDv4gHDozwyt
Q7d4B2FWVarecBhQP9a49E3UjShb1/HVyhRPtnjCXetdQ3Xef+wwXot9EUNbicmbTF/UP2qVuM4W
ppK/qtlvwGUr+JMClN1KY6jSjiBz/O1Vgk8SnGNs9pFt4hYhiWQTD7+G4g+SM8Io/+UWSoamqFN3
9LAQ0g75fWZTpJrnJ49frI/6mBg+ehfJG1tOkeJUgDJjz6gVEYlhMFcsHBtkXRft6lEojSzsXRI4
L4Dl0iPEljAf8D8Dryd5ka25dc7g0r+5U1oztnGUZHWzqfW2K0FXTez9Tepuz3Qp2sYcOqHpLAfH
MxuawS4Vef+TR+uoDd5L7HFhmvKTZ42/FgXRYwqBMRBeFZy1Kb8UTa/9UwruEHXrGqxXVUQBb+gN
rYrKLydIR4qsUqmklIqoATEMFkS+5pnJ3a/Lb2onLsdJqEXzxwFtMn9C1Xg2Bmg4xTmAmrORWuH4
WZWo070/0lKIuDwzls28/hGWUV38sIo3i7RGavp6/fgXSZbDcez/mrmQy0Ec2Rhc6yzfOoI2hR8P
oLKTGvdd6AbfH28wgVqIgPatFHMcYHo9K6GWrmw29qWa7xxgaXmngrHrRu2FjPKLfmmHz0bA2Up9
1U/UnHLWisg6zXO90P/RhIvG/gnsW2N4PllUitWWH/CmrFPa0X3bfbOJq/FW9wX03dEs+TUuMzxb
5mA4RKIYzbW7R0HXCKMvakt3N060O8PGnbQdUcqtuWKyjz5nYzXWplIxTT3WY6s3ZoBIpVmUaXOY
/adekx/cxf1S5xEG6SkP8xn8ZVUVOIqTLbM/X8HWe13ak+ymcfroXoRJXvtyLCn5YwDef+Lgjx9S
WHHZkTobH+Il6pPD8xpJrSfk6WadCoHYYbuXQCClyTr85jemGzzrDzVmM9eJO6ewv1c6Hv5pgbzF
kFqDjQJjSBWzO2I6spU8OUTwtHdo8/nAbJXQeKCw98Xrzv9ZN2OOk9V9D7ZmQEBGq9TJCSuQjhGb
56UTPcDrZCSgO6ir4DtE+eJNJDKSDq6H2wdR6dKZVOEyzlSFOb8nSVbO37rEjrllBT+h2r5XF5Ni
xRmK1Au+OkbXq9hfno2I9+xha11WsZGO6GdRAZ3fYCUt8IA87o3Yha4bEYwH9gy76NfwLDhzoN/D
YSgbhTNKwL8Bqow55xHRoBVW0VV0trpIG3Pg6cS7g4Mn2ouI/WuzDcn6lqeT/JAasd3eAqTn5o4J
ZqAXCokzy6/5/Zpsl6pDzgsK2V4JIEtLLTtheVO8y1gCY7SpNGBqYH4QbndNohamG5TUZaTlzQfc
br8zuwTkjU79Eg0UnzEFUdiihYB0kLQDHADCLJ/7iJCpoIDOTX692YkOdC0V2MPi5GUTLhyIg1s1
HBItsiIZyDSOeEmSRtDc38xQucLgF3uuFL029DCqcfYaEFDOcmG/0fI9ZDENoIyHccOtGpoOqyZ1
V2KwtjsbZtbyJVBTx9m064yMRgVWxhDIlJr+5rJnnufWnd6D6Xxkx9dLfUPmgoPoMT17zFU+9lyG
yBRxNRgj64BHU/pdgENaamPOINkor/gO8rBsAQ4EGfmN7+5xKhLzF9kl1GMNIHjsr4y2+WsdMnQP
vPeBCOqm4yUbh+g5MJZJSnYGmDnUBHlj6mc2Y6quezXqB1ApZvPwUetPUKRw+90b5QrwEC01EvcP
ExdICr/Q+FiMYP7vjXPO5bQtqNS3wwPvTGeP3ayk4sZ/4b+itRzY0/02qPodqIg+VfqQ4cQqJ4hJ
JN3U0DgHt9syNbfpUs3GBa4ep/OPnmituynVat7xUEAXz1bfZVQn0F06/5pz2HcSuEHNMQU5QPXM
WehUCN/6gMuqVP31Uby5ln7+iZ9CD6XkKlsgYU9f4g51tN/5tctLQWLLRc9HxuOSk9g5y9d1US9u
WB2SU13ugVU5bpsg1LvdtFpS+AXSrJe17c6+tVB1ShYwq7genWnmVBmFdMADyZQQjUfv9H9O0QT+
l+YixP0ekj5l5SUOcfipRNYC7Pp4fgH8OYCmCS11V2vVUcG0TbgLWIk2cfVE0S5IWT3jqz+yvc6G
13wyxV33Jhv6e3eIYO5Obqf6Umh6RVJpJsJJGMsgr3m7kdsHJDhkrIwCVNHsWsg7ZjFrOXy7gO0h
DJDICnNxFqh2dKzqCH4+kgEiMMOi2esLdRsS1NHbPm3L0URDrSa3SDA0KSHr5DKQFKo/uFZq5jJJ
x6bQ/ZmdFEgu+61EjnAWrdmnnu1AeDNemeMbyF6BcetWQx4D7MKDu52FrqBTtHgfFeu8GkCtzvbI
q6HzmsEbWxbgVwu8E+ffaszNvPf2z44CxlAoukMakwN/7izm4Pbs41QxoxEgvnOmIt7ubKYyUb8g
jkAn7Xy7It/ttj0ytqdOXWqTWA36rxPk1qQ0Bx8ycJqfXFq/CTYySQX1f6IGvzTxuQkJFYg9cR4S
JXI0+KXs4DOR5yYk+ByHEwyT9hWn/J18Dh5uCIo3UXeWEcoe4QtPz2hnPpn22DKHD9lBerz6GFc8
Op1ssxl8E6p+z4ACQlKC04HKp/U8Xa1H+OWxalz5rvvVzlOxQnzcRfvhnxYDUOru++HAu81JNVdT
2TvjNVGLXmB5rca9WC+W/Ae5RQaKmXWXwSbpCqBsDKExgTJCHaKqKRL/JXDHYbjGKCGMDfW7cItr
xoov1Rb81x/xmEIQvHSMAhGNRMluMIfza/0C0J120/Ta+C4c2sx/nUuILj4JRlCncpC3GHPsQ6z4
Uzfn5EA6g6CDesjzgliFbrZTPmQcO84cNsrUMStGAmvFOnE1DpudXhBYNb8nJeoxGktX8i2nkzJp
UPb7kwGyAMYXO0AWhn1KQw9jE4SvqQLbLsJYerscpaGVxFNf6O/UUtRVC9GQ6Uha83bfWg1FTnlg
EDpFthxmK2k4prfb8BMDeTbKxmsxZ1NjJXK6MUviO8zJoL6wAxXuY1zWVS9sPrrD4jBCUGTVzoku
/pBMFyOTaAGMmZa9wQmWIV/lQHPKzzvmAXtoXEysPwiWJS/U88+Y+Rz/U3mQI/YMDPgrSUd8b/2Q
qT87voJiumGD3fa51/Epgfd7KKTd8pG1Nq4BF/aFiVskBXZOB4/ItH3WVp0ZyQIUokBhsVKVgk88
v07jtex/CU/htGiC269OdCBB5JVv0rTHpganQj3VKSBj0RB66CQ8D9VWhKav0j8sEQaZydA2xyen
pubbRGJSu5g53sg2Yo62C5enGpIeFn2ZLcRfkJp6h2HjSnOVKL6EqRJC03zoOJs4IR8I6VLZ++1i
94wNrOH9w/QYObWVM0KoFPcFvThGrmnxjQE2vsCCIDhHuLdj9Zpc0JtpjFOdvJUai2GQ0Xr+LTv+
qfC3QzbPjd+MHOgQ9ZUNnIJQdZ7BC9j2E/WEsJVB/zZmwm2dkZddYshEyEVmmnn7gUCpFipac/md
28Z9wJUxSgtZV6a0KhvxPqHP5z8nE6tOvi6AuyAktjjux/RpuVsuoTgPhTZePrhF7IGC25kkppyn
Ex9Jt6KGUA/WoBEjgWjJYLo7wJopGQHiI2z1QQYNtM27uQE+adKACU8vqswR3PzB8aS9lAjEUbsn
JOcrZH+QCGDOW/YRd03TctZHw4Mko8kVy6W0YZc9coo+gJP82ydBwz6WbOv6rquTQUo4rYervNlE
3mxTYzLumeaUVeH3PAMi0/njx4WOCId8iweE/tS2saCjYtN+wRcwJ/z0bEoCrJH1msvsfgMNVUtv
J+hzVx6LYKJouzozL/2SqPYEsF0rCboqSA1KyQqWR55tXXGkhI8e41cU7kTsTDtXBzYN6d9oTBYr
bht5FPLb7+ZdZj7Ln0kQ+rxYAnqQLWYNDdrmmPd4cN9bNbalCGBUKa/lZAbI92ZOGVyueSMAfBvW
5eQtQqdK8wwdwYR/hENnw9r/Birqx5c7ZiGHUKN7y2fqFSyB8UHhko5goNdQm2jmf9auxn+km/Kl
WLufyTrWD9jwytgnRw5xAnUP9AzQYx1Hxey7kn8a7g/X6v579xQkbUqi1OVszDyvQy8vi/bNQHKP
XUo7YR4E9bRwj3tzCh+fEyPiy8zsXKCR3JzLXncUAbAjPBInd8S4gr8LFaab3Qgoqs/v9A6k9R7F
yMQosZBm2tJJCyn9i5yLiuygoCQgLDECrvCi922V9MCqIJYBKyxLi6YnXtoCTvdqNcCClnPNfZN4
/Gc4qsTI/1Dr9zrRlYeKG7Cq+SbfnE3x4FUtXtrMzLCuu1jDRqiO0xjZe+lapn0PO5u6xnRAcYdd
icqNQSHpk2+B4dj4p8lYaS1WGWZy71yF3J6ZJ//C/5rTgDbhrSF+2YDDnu38UbWNdGYDWXqZB0DV
XyExJQAC+XYF8xNlUUX3ZNMSjh2kyopYTzLCqUQXHTabviC577IeUE/enIU6OvJz51uUw0tcluav
1Hn2B8PN6+zA9W8nN0/Bjq1rP90gUotmGmhGevKVnBWMzwv/Euc6BkAu2c78BSYiS9Z798BfWtcW
yNoCxb3K/8NWZVuaU5uJ7ri7q2nNB5uB9+X4bxEGol6tQ3LlVBABiQ2Zyh0qgcMszLXw72E/yo35
S8JNvu44+jpua+z+GPm0kIpaTihATmiTh1frxDCAhXzHNP8sYohl35K+8l4Pqo8V+qb04R39Nh2i
lxKCMJHKOo1xEqAK32OQzh7LuLRlHSWh3lSAMM/O94k4RLdKKvaWoQyVzNV6y8pHGfdEJ6qEjkc6
YhPf8hrtoBWkSBGBxL8CoTDbl8HXu0gojMqWIpJlS2uth4+p1S1H/rifO1wpKjdmnOFjEOAXy8qK
2tnM0BXXCjuNKM2XQqNRRtwNtBNLrR+qbaSQKkvvaAjz1VmNc6gp8rsCa737TvKuGwFqnZpirmXW
dyryW0JsGpHmuXv2Zz5f1eNyj0Nazi2VaxOHgjYYbYtwoM01i/Ju3gAgXYq0tSco6aaIsoGA4Dxl
VX0QWBPUiBY1z0ovM+75VeWaBD53rRkjSNmKUVoOzq+Pjqn6fT4sGnku+5EN4qT9xARsp8bVjAtm
Tgh++TPKV0Fy+d143u3wz579OB74sU4eR0w9FV0Ik+2eh5Ao5QB4OaoWXnG0KLnoSlg0fQxKrFwf
46cTKDlJ10e2uDR73QdjFz9IPfyCwCzTRdvWZQiYpkNmBuiKXULKZz1c0+1NuaWrXNXCZHrVXsFM
Xywsl0BikFPmDyp15lcZ9qmhbbZYbxL9wzm/E5oDyVCmmZXklczBdmz2BtLCpAXDjNfVdrTIO8eT
ggsBpfiQqiBUXT0sXCujQBgMna9ylUilrsNpIfkIF4D9bNGm5oHrXGNDP44vjL2mY0KzfO4tmjgF
473IOuLEXpoTjBRqCADAQzCFmm2OX6FOgj2uEqn+GlRycfsoK9ADE9Ggsx0dS3Mw7hne516CNULZ
KZ6M8XA3fhsGjCpHp4Gb/Oald7HqWz5oBbRda9TUmH3rvMrCau4Tlm4c2bl/pz42FSMgyPTw0o3Y
q6MkrJkTf/2QhTHectJFTNPsWtGWb7HABQJM64vbSRGOmZGBQVAzifaX0JyAeLPIJiP9WDTf3+Y0
sHPICd9CnFVBakCqa7eoNQhgz/qRt2rWy8LSeKZZR1GUG4ZscxI/B0pGOurATPcw+10+CTtiKvXM
5EcT4j9RTXWs/jtI1HDsQgotPv8xosWOJx9aGf+ATwCvhuuKI3U9+ussGI3qkqzaTuK75kM3xCKe
ExXqAvCz7IAj/gcGEcjL8y9ftjZq8ZxP62iuw6hIL2hpsOUvLX96A7ZeqlYMA7uQ83GMfEzBtYE0
psVb7/x+AC5rvxsv35oqOYQ9qkjG30+pUYLhMUVZCl7vIQrwaFZATVXyAnceiJW+Sgz1MtlAjELB
xuXUj53Xc2e3dYponNF6YUXJ4TXIPtRi8vQVeIzDdUW5t7eJGkXUagdnnGwRuUr/rFP9Y1DRP724
YeL35ve/PIQmC5BaSfDvyVVFQcsUnySpyjiW/bD4Xru8gIyckDzwmkayA5ws7A1PctLJSqSFeeQs
67AN4xjBVeaNBhLQfJZrxrXUHwwm3FH2gl+py57OnmEg7PfVrza7uFcxAGIHeWK/w77yUZo4K3Wx
LxkpDR4Ry3m2mgvmfsXohqRk9KiHexcbJhDZutT1CgnT2fy6F/wuuJF3+0SVAnvVqHRQY8+Z7m+9
rKh9gLm7OeVM7ZECrNasM+MvOmcKjUcO+9mS4yyH9szn2QAEpJy7qAWMZPsivxe6pi+srsUrmmPR
T2xD4PUNhQMVC4peLxYTbIqm4JXLrIC0BVTJm4q3r9GYMwMtcKTd6DgMDSK4RsGjI4I7KmPIeoSP
oGdt5L7GLPJcS45Ng+BRosbZBa4nJug0VJvijQQHLUMbPx73FLM9PzHdXhoftI2zAHzQ2vfB9bmb
cEiVGFiF7wKfh9htVh2sS1zblhHfeHR/P53I4dBCXJod09adF0DYOCLOlBU8gN52r+9uUjwU4EoS
oFi/WM/bExGaTaa2p2LWRjyuiqTXJtGSUqf8wNDZ8/O5IfVoTNUPcYxQvCMpj51CCcGz0Dx4seqr
l2IWIbW64b62ZmdcjO9WlsQnmjxfnkyFkZM87AeRHaMKaliD4aDK9nx5v8kdMRkh2tqJGmUicaQd
szteNx0GCwwjJyc4GMESOy0hO+UeOguq/4LcX2pNNAA88Q+l1Gcr59xDXujZg6mwhZJTopRAzxeV
TXiH3eC60y2pgTi7pkxGjBBdtEZvOIxUj0GgyPGcCtn0OuRhSy0J9xLloy4vehHDzYBGQTqd/x1o
KryPIp6b7zltpjpqUDf8Yc6JPC1rdJjxnvKFoao3d0utMTabVv27zyR172QaSC8gqP3oUGKm2L1r
TxMM96v8JvVp5tRHnNWPindr6KAsce08lV0LwazxPUEggJr47af7Sa2DN4L/7K/4OSQk4KcCuIvv
Fx/D1ONDKJUnlDVneimYIdPz3d8Pa4Ggnu/ab/4SOT+WG7JY+5HbsmbSWd398p8qtd5ZpMb59y+3
2sQDcF47tGLYE4bG3qfnQbFfIilrtM9zG8lEYwnpKbZiNGKIjAF9peHQcCGwcf1u+kL+dqhRuTDY
7t09mmn56k8iPwVTe25Ei3rwl8LKb9p2PS4EOnSI4Wd1RIDXJVpocut040NGOGPRtC1hC42Zgfag
is/LbpHsueC50VErP/i71Guy1Lu2KMR3N/KdlTvMWpp9pDMI7lCVA9c2reEM9u/A+S4hwAZLQ5fW
fi0VN+X6BOL7lCkdufACyhRfwGHX4/7bYor4PMvNUZ7z8Za3JnWT4kBjAYV2qDCnxuNR0DuxuE4y
4P3ZYIehnRVPvIXjWwkLw/NO4wRGM4AhXVneU6OYCGKtzRVTmP8ftmuI81zJv8Fjkvj7SKxrXLfW
OBAqVPrrKBH+r1IQKpmPLAD8BNgD/ih8hF7B81gIue5BJIZz5xcA3nS6h+GhfSW+55jiDnMnQDlD
S4CU7PQL1bW5PNRtCn5bZgq3W0lRJruqcpR8xGWAjZdi1zXztEGHF6gbtTJMYxWnwDUxyCd4MehY
OQWwTPs27O+DIupNy7WDMOUW85YNpa0sjEjvjA96BNfWEXcYFN13GrOHVjSnzzbeIZRgzQiCKQmJ
BaXUxcr/MUfh61/uzphwafmrCwU3ERM3ApbQYB06TdL2WB8w+15MDDraIqb2f9z5SEfaoY+e+6Zp
QVfkhhFBmjIaas+Ac86quNSRdC9aqZZjO9me1jRe6I1w272LEE2bDQLd+kRB32v/pUxbrZp/sasZ
o5wHY3VjWzt39HEjQNfuV0x66Ch6R3EZfNAsEV3Pg5OMS60xhJqL/dn1v2a64ZYodqlGvQ1FLZQc
3fDVdfDM197TpJS/ZjgInIjWJiZWN0PqPx6VzkcqC7m1G73AetbOKusWGHZ8Z3fEGAfInTqt4K7h
BWh1Zqblb1MMDjEirA/Qp5to2VVfM3OoTBlSN33xEb4FhF/uGn4G3Po6zfOjhrP0hZmWw6HJY457
ePj4GPN/YLYW+kGDolkMO9aXedotZA7Qg3fX4KuH/Mhi0d2Z1OnqftZO1KNHupY/xwpRMwxCaDaJ
f+VZOIvdFIJPdfkyiRUul6S5GOJEo+okcKgEHlRzqcwveSrMuGklGBJJBK6V9Dv16Pmkk1kPNhpI
B/vwXkieUJX/I6scPImkIn1J2va4e2LHB6mQ9YOs4dJ2V2tUHcSjnkMw5QgBtsoDNZtp1OKemFWR
45XmrQEGDZAZzGsenGvLSR7bCSZ1g3ctznAkCxJzYRtXI11niTBTgnEiLBj09NPp3uHVYx6A50Xo
1V9wJ/Qp/5aG6xA9ETezsS/LKhndZ+WTrscE/VDRPKTFsCaXfMoc4b2h5nD3miUyCFS4FR828TWF
d0b7kfY7YD92QmUrOl4IW9xUba696uwELgfjwk+TkO2CzHNN8nbXPLcJcbx595hOb7MzVSVss5VU
jLViAGJAySPdYb7xQqmQKUYnfVZRYq9dtNWvD/7xDbgLxpG0VU6d/85cqdxmaneQSqsajrokiixC
8vyTnbe1FH80FziDsLVugwf6OlKwD5TuM5G3FWy0x5jhIJPZflaPBiuvkBjWeEhWjkx99yqusbAZ
QDaxE2EuGrqeGjqneq4Epe2pVKRqcUMbcJ1yFNkEBCw+pkoL78odHsQL7jJKYpc6JmCwC4vC9yuJ
y4KJPX20d9APcknz6bIUFPC1MPGDq3H2o7q/JaVvzxOROoN5BPE9HzXWF83k6BtUL0v2Nr+XDwHt
hUKilQnU6iTxae914DeBDEgUB44RZTgn3GNpETh5tHhLEiN4w0Qs2c308o7hbjbnpDI6CzvaNzrh
C5EpW2qk9nYH9TLA/sIqq6D2gNpzxMSQIvAkv2usjEWviSX6eRACYG+63Oq8tq/0owQmcdJswlW0
JiTD3ucBsXc+30fM8gWaoc9lnnsqgMj5ary8SwXf59xeBtZes86wer+gOk0t+OdSMZXraSrEkLOI
jiguitn+KhrudHCmexI/TLHVPBrTt221JdWnfwCsgdY4tfvbZ5q02orgoYGIKrXOTgpTCxdv0DMI
kj/WOJc83LyaD4HIjnUvQ8qM+eIR3yBru9Y2fMEcSflsTCM+DyEqEYvj4cfnaF8wOPChFL00D3We
F6RYMaR+jE0HfAM6zBcXXZhPLir8/D56/ZKCutQA91zkEDhRrn97rEGrceYsfDdbH1vrWCmnT7G0
I93J2ZvEWc5j5DEurqlfxopVPkjO7Qq7LlTgHJ8EySXbJrj1B43Si7p9BQcoEjPINSL7+fKbDLHp
YT7OlxaREX1pCltB76d8b9uFfqW9iNCURnF1vpGl9r9bufdd6VgJXKNvWxz0Gpn2nyGaiB2qQxHB
Ch71EINeszQQOrJMmQvbRRzvfpZWL2WJWzf4644dzoMEjxz62c+10kTJsoWkT0LKM10QVHQS0M2J
FEqfHkNA3WMjTEsBD5hOmqeVOxspGMsxd408ygaHF3IwU4R7YDiGpJpQGcCK1kZe/DZ6yslKg0/K
zRtH5xIqVVsbLuyvNxXZ3MBb871ht/x3qw7d9D12ezNLLvl2mUVNUg/A1bg7u+s8I83Z/iZBvnKi
FNQHyDMAsuSPRJRdtnoXM0Fm4k50PdErBobCWzj5ZBj7FOxA7Et7jRdz3TG2wYZ5M6H99+evCDof
oUUeB+wvpYEHTVQ6RfCfWZ2PHgPuOLNNbwFF78ayaiOpRQqDYNrUD+wlYxc0bWrjsrfuH8yVmaf7
JJkWeeI+SR8i3xhtZ6wT2YK8DT2ViD5e8/qFwjdVeSU7Hj62o1bdV5OWVMjsB7nIZCsvABxbGRtp
/jh9AB64bK7fgD/ZnWuhSv9L4jR3jIRfGlatBM3LcCZlM++lEkV8TZDdCA+KygThll3WgmYliU1f
CBLzsEMbesltkeXtNohtnlrvE91+wJJS3e4hHKR6HIC+lXglp7LS/MQDRguJ1n5thyw3GESSYOJl
A2t+0MhRZS21LyQGRET1f55x8nuDyWnDsmBIilDgSGP2OfLrJRGgljyyfu7dPrXqrYID55XBPGED
j+36p9cBt2dCKrWsnSPX5jS/z/j2KCMgTHxGzNLZkjkmzy8x1dWCz7xt+MvEBpc+3BPije43w6Pq
FR6AZiNCcQl6vCVPvf2VSiTvE1BZIq1EhWUieEpNORewb4bd8CA5W58tPtIhiQUm/9kY8pRv1odN
zjBvf461YplMzDMSUIIZJK78W2EoE575CZCXVG188Bor48qkcY/d898IT+Uc341dMIOdam7oZSrT
XOku8AadLZy51LBTQuFTX9xks98pgJH48bRA08yAPKkJ65sqQwqKh968wG/SKhlbFmU+xtHfV2fw
k40rG6ujPq1E1SMoj92IKC/kUrjn3Td4lhOmILet1hBA83WS/5wc3VOKMVySzQuJ/GeS2LEaD8Bj
41frYIc4i3voZqnWcKd5pUPfp5asBul3AHfH8XWGeLwKNTTkdgEkQK9HHdlmLGB4AX7M+ovtuPCv
N62Mu2YD/mKcWeMhuPsODZ6CMYZe0nCzpckB3jLBORVo7m+Eh8QbbyXSrLBFmazKe0QNtDdV98wD
+v7UZU3ZcOAA+j8USaTkcMTHQIn2nJvvKunMZjwk2I4/VHNld+Hmv3mp4XMbs12okYhW6NIatK3u
lnSjjCkaunbk00c2ImkhAKgyhccjhxzSq7wUtvM1SHQud8RgIp35K57/zHwsuIzKwEzyVz8MaAAu
X9em35K28zHNR9cs3j6KUG/UxENh7kieRTokZMdhFJAXXu0mPnRAlM/z11DKVmYB5ppwYMaxTYN0
BqlPRagsBsDmUgaX+ZZnkvw8WviTUxTia0ytZhBT9hHhmI2PcFo+6q1ErPFJvCDdGv/kUTNLteWo
3v5q1C9cRRDyw47PPEgqasvD4TLKL8+yNh2LXXPwxrdkvcdMOvhw2CMf+tL8jbyPQGiYCGUfHQXT
J6pnY79tY7AZcAL2CvHnj3ek6c4ItPw2zsLfygxQEJUDKJl12tWs957LzJt4BGxqF8bfLeb/XUyT
9egw6SSO5DBOSg1L6w+xPWfp7AedHgod9yqwtBiefFadb2mtY8tVjY7vMop1dV2Yo5T1lyIshe8w
IogAsWJLczERHaOz9QABwT7WTqWlSwHGMvp97vvB00z7NgBVHDbpBiCi2RoQImspSzlQ6sdRTAUU
a5kV+D91ukg2iswb+McihRGUXDp69g7RNWxJ44SrJHk1r4JtyLw9gr3vz4Mio7quY+Vxl3nghAGR
T8QGkOUFc5qnrRmzh4s8WGhxcAjPZ8PiedBvJg2M9fjCka4NBnQUyC2wW3r3/woyMWiGYydZES8t
LMgeI6YAfzWCeal94XAuW6y/LyeJnSGmKRGBKp7Y/heHJdDkvzYXsFT34C5t8yQvbcpZYZZyhZYl
zAEY1UKab1UTNO2y0dk5qQyAkbNx0k9BvD4z8QQmc84eXWGBQabIkmkRjaplFiyy76ondRjFwJuc
5KXMQgmSvSIQCt9pbRw58pXxjar/MvHLRhQajoSRQKTeR9OdO2gXamooLBOveL5Wj1FLgvMa08/q
tv+hek4ioIVRDT2TH+HLmURHMxS/ij8cl48IZxPZ4xWuXP+3wskHx1K4QyhIeYtMs3X5o9sD8ipF
7bv5+WAlT/tGb+GtMQY9mfaJqnwl6RfHKsfXLbgpIpx92e77IqnnP6S0S5Y9UeOtt+2CXyB6IVU0
camzEZs2bBWeayHEpWdebGa3JC2Q+pJBFhYSc1X2smzA98hwwX+n8qFJbtVsG5GfLbr63MFSHH6S
wEMiGQYveA6LHUxbFFchs2su7VTmIbIg2T/tjC/aW/Gj2oQ5m2bqs7QE5EC9k3jYdgLnCVJZ5rXh
pTtGV+fG9i9yQ9vR7BgW2W9PfT7PjSq05CcdHBTWZI1y1aqWRleyl/qqhqC1Rx4Bo8GTm5YOJx9f
QFDMufZJs6d2LJuldI9o/XsoiX0aVZ4S7MzD2EwPBCvMaHBfiua4a9AdSwX/nknU4Z3Er60KIzZS
HeITPZ1U/bBMqCsdNWy+QTRKrrVciE4OQIfEBq7wO6n75IpPlRYq+cN75xqc/U4r0HsItZ4LjDRS
SYmtj+pTmNRSIa5fGVOz0J8OhqJOHQZ7+yNHEqTOQS/tBwAZ9ZLRtSmPOjnTNSiVx/hvCjQLlqfC
2R6RVSd/6IhmNiDP1W6e+syXb+I+jWT0zIJg8msiElvqyCxiF+VF+qvutDQKyTPZKl6yI/sSNOz3
zQMLPsUXjpyjulC7p5Y08yPVTWomHQIW+QTxQ5Xzvv3qMWGYb9ppggQbYiqhMJ8jHdQ+9Yw/BXHd
HGmgsMSi5qkx3eBN+gDWwGZO6fFJZOhNxU/iYiFLfEGoRZtlLn4xNxv2RjCTaMsHyaVNSGLtLVmM
aQC+XN3y2wfWXEmSY7CsUvv0XRgZBQnUxrr1InwX40ErcV1m+U2pnc9qhBfmS7TTVUNANpYA729u
nIYAC9qmZTIYpx7apNRqq5YSSXjgnMhCu+3XtZdfRyVziE4FfZocak5X5uMozedkNQrV9aR+kH8P
oYqnHt71K3nm8z5PC3ixRZ8T7ArUx4Yg12/2IZrHaACarz9+09X2UmmWCHQbqKjh2eMnD4xJz7Qo
zDZ5a0L+GTiTgYpXDc+C5KQitR0VysFQ2PZubmrdybdB26dwk+U4QCvQQi1Ffs2hBmTQ/E1dkEPZ
SWoxzF1dxoNUapwP5xNgyfRigWdi8RSYSQLlAVo+omII4lQzEEV3Ix6Rj83e3JPA8erG1SZ6FBvT
HoUHETYUGwrMf6G2QXqX0hqWj5GQB7vt7WbMtboK+lkKyGsjVUxhKqZlh34K/JjSfNCFF6Mti05u
pjiDk2PELNIe2p5b6n/t8Y2KzpJGVfmGNRipGsozlQNU2McKaJP/Jx4hbXBzVDZbPlNh8Dx+xGeK
RUx5jTs5zsDrgmNHnW32rNiAMRSmyYO3fvopo+yD9QFTBJn70xWNiZIMD03c7ZY/Cmdn8o8zf03G
pOhsqCgr7w1mZZJZOxpma3tGzNZsLV7OW7FEFksuYTpLxs49sv0tvVkRhno16Ys84h5Jr4HwT1yf
YVo5BswsBOSmpXZ2sjMQP+JFTLjUmTt35H6gXsVi5WyvPb6ZqoyZTOAw1LljwPCDctbBDY0jgfhZ
GMvHZcVMrLQStVyJBzVkwYxuepmaSoRxxyUqGkndg0zZ+BdxEAn8PoCf60g/WAlX9D3vhbSwRV4U
Cjs0cLSktU0l8IxPTo/KqSKRqz4oKqcsPcXVTfPsv2ToyDSCYruecKB4+4tjrd/SYxayrjPi8ufx
n7vID4LofmF5BIKVNpo3kCU94o8BleN+kIpT7QcyjGmxrvaOATqM7ujiZX9xWvqw0s9CRGGy3xqK
FZa5PXumb0m7criDCGb6poBVowiVXE9FsPjHV4Hq9rY6hbHRgMq8R3JuJHTBDMP5ABS+Th6SllTy
mxIdothb0mj/xfzJpa9QAJ+QnuyFUGIDKmI7vnscdiCvMyfGmkkObV0QFIjrKFsgKDXB4DyqN+4k
FSkEXtxua3dIB5/OBTih7cBB7XzC9juzsSLLeYtgdz+epBz8auENBmcEdAp+3pGEhOUuc2CkaKqj
pNprM/C++DCcVO8sJx7p5SG0llRKprBJ6XCz7fQ/cI+rUrB2A0BZaw0dDMPOcy2o9uA0BDPaq/6Y
pp+N4ZRerUkKamyV9SZHHoLA4s6ogKyhiA8Z+LiChM6IowZwK3KbXBu7pERJ9cmlFc6w+TPnYrpX
w7CbgSrEkKnxiLj+p5V9/jmXh2c/as6v3/XjRAgnYtK1dx7EOGlregzhvB6fsprYEpLXcvgXHSDS
Hq4YSyDdI5+oK87cmYGD669Yen6OTeGBEXxetMMuQQdRbGW0et//UAbfIJtFxKVHWYiY2itAcR1A
h/A/A01P7GInoU5vcAd84Ph55GyKpC/tzVRtudTa3SLKL/G9me/PmdtMDEOlk9b0fkVqP/+T0+Tq
RH9bmjquLu1aW0njP/O0zUDtrmIX9AqPZAxK25rtGksbSHkEN6EGsLf4UlWX0nJSz+2+z0Q5sHIK
1dQvL3sKCnMDpHsuOwmTAJfc/VrBsOBQ+H3yBGEZEdD7OKViWKizpjpotb8KUv46KqdoEQUoZJbY
6yvsQpWRKm7WTEoef6DKPJQTYKQwyYlHNd28nlCBMnlVfXvJyRHr33pjyS4ztRLP7tya8GiRLT8c
zUul0b8qmNYNa9fEdTWgNYnPVMlQ+bqABFOynM1Jex+cizgjcz3MLY/ZJ3WKLx5EbdwYl4wS9lOq
Q/+ixdleRJDd4UwY/RfYN5vmdCX176qz0UJTgMEY53tt5NM2/l2oW3aQjEdVo05+enJtihDoktA+
TdU4Y7CNPMQjjQ0XoxEXLIlx2rpKJmSVRK30gf/Qq5rZe3WsHNmJcEtE63u8u38zxv/mnkc3Z9g9
kGWtf0ZPbTrtUPqwH/HM9lb00+BDNobWi3m8r82ypJnrQfBZK3Vei4ZA15eOxYjLoJ3dhoFVv20T
79tVM1cnX2TeI9u97dkThy4KWxpVVNr0Zs5RktBXBHFMjdSBU2CB5JZmDkjPB6uyUmypxvdf9w3T
PboYd7omLzznuWtrll7sR1z4UkQoQZmKjfgA7yp4fpB2S1QjJG4D+YwHOEubspD1UVrMQ4IKhOiq
cB0tugEQFaXgownA7vHpGh5r6eu83T8v8g5C52H5AtcDZ3R8biDw1F7Gy/zhHLMTtM/lt+oZ6gGQ
eGtZf9LPptv+rnK6cloxLOEemwH133N86vmchoDLydTugXKnY0Udl0IvpiZE/FERTuK6ojoPjaSc
mMMHProjRZLux3Mj5yM603hsM/1sdWscglD8Sygmg5q6uOXmca2Qvi7PdXylQ3OjChXlYLgwo93o
q3racSx4KTJLzgP9Vieqw+3cM5Lyn8tuYjSIa2+TcR4iWi0Y7/Yb/ofPVICg/XybbwXWbZJ3iD4i
97n0s7+15X1Rqldc56R8kvX/mGnvrSIBbHDy02H34UeK+/ChIA5UA4Gg+gcSGeN+Om5Fmrhvurdn
j18ReUhklFBAABcm65MkhR3txaqGtXmkMdjhQfG1vxfTUJe1ifKLxKjkX0MluLER0pllD21eyoOZ
xbwr7Jl5CjVdUO9KgybB9RpH6hNkkfpVffeSFVjGJL6gExcwpiMJJVgOWbhZqWafuHte8KjDzSLl
OZz+AWCXyQ6kPVdXVeXrfsvoWVW/fQSZHu5M9TGlHPWEMJgpb6SjDMf45y8Jcc50X1NO4uXMVQu6
qLsliEGj/lKRqsTiT6xcFUwHMhcUGPSyFlHGApfF7TXcqYmpzXKhDboiyuHr1W6h56mUQdMqQuRs
glLURH4+tiSP/5vBYt2Yrdi3UQZQMrqrsaYQ3Ok8OW+Vq7SzGJMvvJ5FCMd6cz7TlP19FYkbrzq8
IWk1nbtN4xmGrVcdvQ3FEY/hhwicbFM0kT2N8HM1rLoC20CwOwwPbdjM4e1Un+k43jUT3xcQxrgy
CdpHlZxgJAIbQnwd1Y4qaYp4Gxv8X7TbZDGrKARg2+5rEIWhexvcPJAb0ewTQ9QNv9I6P6bucotL
A8A3hcBOs8UF/RC5gcsMWqTJfD4lD7kI7qZyEMGIiw+Ol1VANuM4JYy8uzOU3vhm8PQxfI6vy5s+
2In/AHzhou+2Jeu5d6287saRHb9kEij8LKyb2IAHS4pqn0RRvtAcsxYyDB2Vzs7Hy9KS+nYqf8Md
6NlZytlhITfjLd1S78LSNg2Jxm1ZIlYmSrlKouMC/R3CS6dm7m/g+0qszHgkCNDIGeOC1D3VhwVG
rMwARIzgWyUlzjCyfRVtEdWgW1WMORgtTterVZo1QKwb/NPydWbOOqPDFKsvXQD47dY+VlG73O5B
bjkYIZ99oBSXsoqyWNUvqiHAL/AqJKMspERQu7KN1XYA7VLEvbZEh8Cpr42VfY1WBI2zuBCXmQOJ
KTXrhm+HBdN/7XrNRNOZ87L2z4ICpmmObFDxWndk7mJU4qzdHKcKT2+rBKPj24n3DfNxevy/oCDn
06B8MrWgDm0MLfXVo5eXQ8My3EKs3BoQ+nLXtb0Y91f3VKXXKQvuZu8OxNB61sFScs/5vcOpeH6m
hv2B4aUlGwhWGm4rM6Jbw4iMCUkZM3P8sX50v7bEvJWLFm2BXU6yQUPWRybb4JoZ+DtKGOPRiejA
OdElSfx9dAwuVLnvfFvZkm6WlstiBg0j22TCEqcvKCa3Io0F3IslQICF2Aj6zNNg8EWI1olzwv9l
FaP1eHuAs92Q47o68kWRoli/u/5ay57CCYmMII5HkBEibxaZFGuZls7pS/i9cfonZ6nG725nmHuF
oBW36L7BsjJfX8Q+zYeMRek9yf6T2mjM0gyBzQr709A6DI1rqSBfGnEEp4aLZxeRInyHwF0aLcna
HMJQKoVpsMFfonvhszCnfiV3pvPgyAGczv1ed8NDvT+ftQ0OBRlkaIoMy2g0Mm+8hUSapbxRFsQo
lecdfwHPuOm00Uq8EPRuELlFCQpa5qfSNMQflZjcGb0vrcQnp6NBgH2ETpBDNQjU2BvfvTSBLBr+
CNDRr4JsjhRwL97MCmf5T44UbNgZFvmMRMzHvSmHJsxkIxUfNlSq18ItKBMRInklWmXXITFnsBeX
jaqrvc8aZ2ogSoy9jeg2DcsmcH8/lcVYQ6gAvoAdaO7DAuloNptT2mSsBFBkp7D5cHYM70DHHS6k
16FXkooxb83BXFM04EpaQfr6QP3xPTHRJY/yowgZ1b7PHkoayucnXyCeQwarWbqKp72XTOa02uPi
tSDSCE5hO3YBYHkNPb1bhJu40G2djbJTMNDVYjPFKKelKpY2ryBYTM2g5dgJAMuHcglqqS5Q6ueN
YUJvvyuj3a18M5CAf+Dqz2vW90PckIASlEsDnHEblPqqcpBv/Wg7N1Bkeff43G+IFday2wPwW2G4
7uqLuXVByTRxNz2KYInaZfQyPEiieVPGL5vyLfYsnHbD9eChnS35pQlIlY898AjkeoVmjFfLoCgr
I5x8mJSL32A9ERHXwYh10oApeIp+FMD1ZrJ5O8tu1QD0HKmULyyMv9dmmeoU9tEyUPtggP3A7O4u
kNdSBCl0xlv9CF2stFCf6FipX5s5v6szMuhjayCot22SAFfVC1R5GMiBm7uzMznzpMmkf71H3Epb
L01fzL4oLfLK9H8hCgbTDHlRWGfEloJeaIKhSADhq2HsN/ft3mmbxmaD3/z+2EBlI+7i6DGCHK/T
16UgOCE4JiCYeM1jHYAcc/HV3Da9aR9dxOzdpstbDo4uOK9rWdBJuj2pzshs4QFOns3pl9MuR4IV
1DGje2/XYdSKgW371yryWmpW2qO5joDe7hU1V0mh1Xhc4ms+puLqoAGlG9FF6zSW1kJakABZDHXY
TmuzjZq5tFBf+7KrbJ8zyXEFn6N9x3kf+R2EUs5i8gCrlpMADuMigO88hBlsWqmgSAzuHLerAq6W
B0BFLCYK4EFxXMAvetKdDi0MR0AwGFg8FEVg3JzCoxjhFRECSL5p4hEncIptB+Q0LA+/ngS0seft
+O92RsnS29+SABzHZyQNz+H7Hg7NdjJUdIG4QUBEZxhf4mi12MFWVoZeeW1f7N2W8mlDQ5ZRBCq7
0bqd3zzue/aEaZPV1EdvWtXPax+lwCz+O9LeArnJafizjwc7+OCi3niergkU8TxhuCXZgUuJf3VQ
HlOWrwFquo15QZTU45eusdRnEPkFSIf5bvpg++ZR22tme1KT21vnn2d5esRpkBvJXjFXhFb89vxj
S+U01mJAlJLXcHkzR21Ln5xiSUAfX+exoW6Si7/0ibp192yYrCrg1jPXVDx/080Yg9QO5vgLVr3u
ci85hgg8QRCMJ3PEFaIBoEVMvDwipREQN64sYpx7R+VeEq8SF0l+LgTkzvQV3ws99AMjrMyNjq5r
YdzJpQWHd9tCQNXD0s7ibSEztfCy7AdjuIXE7awTYYmX/Eoy3h8iohxnMRWbHFvu+EQHXSAyJfSJ
G27u6j9UY9qTw7BDWz2LKYGIxYwUoXbNIQQcwMmhnIz4FsyZ5Q2xmc0CTjp98h8OoCzhCq416zAj
2ftqq0XFk9Pv+Oc0p9Iee82jqiQFy7juG90HOLtFq5VFThwnYjm2Ma7Kll0MvUaRrYHz5Eyzc1at
5tUp2jX9eR+04UvYYahcL6s+UEhW+wCKpFHDtFsrDaGL0N+fc2dqNg+I4OP63OPMNYUWX6kgy9XK
Uh328Bf5Oof4KNu3qT0TKAg4BV3C2Szf4EgSIu634FNmA7ivP9E8gbQ8O14bp7zZVVyk81tbEsrh
yH/lq2ujRzuZgI4pbZaaHIoaDCChWxvAPDTYdFbQQxrQgBSzwdytvqQE84riE5C7CkBclsbpGeuR
3MDNvsI3e8WSoUKK1SoLUYeeSbdZPGCk+72iJPeKAylrjBOotlUQMmSgAU+fydQD1djMwNAMwHPj
4QDEQOBweRx19ee53LkYZKYRIOhCKDReeCBF5dq+gWJi6mM9PMoFR7ZZe+Wh+nSQH7pI91sTVe08
GmUkA2XjuSDWD4TeTavTSDFzuaJFicNhAU5JH7t36bNSNw4dsEW6gLiPfyW6Soyzm4ARYdwHlDvN
lu7qKOVkZEVsZgMHwTYpXqAwAiLDQ130/cqxlLD+sjkV9GiymQMwGHo4Ec++NNHXGHLqp7cxGSRw
iyVFlrhjTpg2SCf7npGjFVKnlG7YzXoBSLkDqq9HZLn32eKHnI1O+9BMOI/woPf2HjcPakrIwR4N
DUtVDdHgCh93C7vu4UCWlwwez05ku+o9jLfVgRjS3vCUvWF6CFKGigs06U2SG6NAiEPIX37fbdC6
o2rkbmFDjSDS5LUDNh7E6FbLB9ZBIYaMSLbPSXOAISrYZZJxkN2WoRPN/P8ZoQ84K5/AHuN1Ai00
qitQUwkaGy5a6diz/hFghuFZJC2z7iwSv0Sv3nwihUmljq2CqH2tiEIXfRs9Qc9aRbwVWUt3AKrK
hPBbxc1mRRmJ9WhlNLGLEsogbCySjVfyQ+rRJs4kuGD0E6TMyB+8ho4fo7/csQyuL3vpZ33WOm0I
3SfbsddjiiVerfTL5iQ7VUHcaaeWELF4u36trXsKDJP2hOT8vQoI/hLB9cu5T0GnxNbjsNhkJ+Tg
1P2s4J/KHGhH6kI10q5YoiBmtSkK+85zs9CtREYvp3JbZn3876rNNBvk+KySouTXKxEQnzbDYXgI
vEHDRDTUdpN3jDZq1VV6rTDaHg32ax9EP6U7SNPz1CJd8AuebpUQjHqbGkue4tP9sb8m6qwO1YjD
b+YgNEWj2rqBCNY9eyzRUWE7+yAl2o7V1w2+QWjde0QfgTYw4ysf55FUGVPqU7tuxh4L542JD0H2
eJbFdtc8Qi/ivH4KMaDTtb+ZGBjDArWKxFUL8fWpG9aU6Dx6ukTeCAE12px39p0qQjXlzy8rvk8G
maVucmN6/PdviB20oE6Fbyvou6LXFjU4pZR1YzbgdjNqE73gwWDFmNqcxoNDnBcvRSWZamI9TXTC
S8y26PhFhocydTbeHxs9waCy9nZYnkBPHsUB3N3Os+sevDi9V9jfcEwezl4XFFNB+ZcgF4HU/XZG
QEVjecDK82RAqqxBsIKlkEvnDtnzRNewi7s8F0uLte66U0qfT0T/wwaxv+Lw7D0rStSDNhJtxlAF
mgVmvV5A9FQmUXZCUTVmzA+qCEnAbFryCnVYb9kkYj6eYm94NLxXcfJwbOl1Iz++zmXkoG5FpXad
LWzYM7JmlNwcELnyhWEofvhwmCSZ6gBQ6P7kLo6ZxjXVgvBHJTxn1nepuKW3O2oTm5hBW0dutXal
LkJZS6MxWDC+2KCP+IbxCqLWDlEJROzUJiY0HYU7dIIs9S5XLNgyoxgRxuU2Wohfc0du96CJ2+Gv
HhpQW8B2yUFzeW9lg8zb2aZONFQVWV/n6STDIcZmIUNND2AS1jMTwZAaUd0Vd8rV/4kAvCJXtmFm
3o5ED+8aeQiXnnMrt/9Ug79v71D002CGsSLaIRnhblTUSUVKpepeP9RcqQLMfAduHee1Nkdi6at2
O4Qxaagj+6Z+Wr+QWg+siNfpTvkP8ufL0ItcXXcwmxwSows80bjt4rJ7NqV9xdvxzcAWqMhypMzh
mYIxaGLU8fhZ2lfVxIHEqi88mMFsAKhY+EbDAVLrPHvaVS1FGLWDHnBptx2EgBeB/Umrnl+uSmIS
SBuHoMNCPkTpl4pqmCqNk7p8QIoL0TdC0zTX0Sf6+zwHnslQQXY9ME55WWye6/cyRNE95MedQNSm
bmIOTqYpU6WZS6HcUSQ6XMkuKZk6dKIlnjglvhopW3KvXnfjUR+NBOwNSEmcycA3qiCY4b9/qCz5
iC5KLpI9Uj4xQj7R4oPkrH3kH9DDRgnFXob0VNzZ//zfeDcBpKtebpV1ZJ7U6sI12ap2Z6s22duO
mCNYuZXfKPa0OVZI+vwjSdTclFyjxY38YQJnlGRx3PwJ1JUlzwA2GTgVOyS4xywIcFMTYKmB3Mhz
pOhMOPcTQ7q/bGQtKTQVTNSKoT+8k65RqjPgoGZNQiCHGWqX3ecWh9rVwb6rhRyN9FkXilUTInsP
L+MRwC1jTV4riQpqex955i8xOpDCDMaT+yUcGRxiUNKd5F22NjUV6PA06JpeAX4o5luUSKBMM9qJ
I9rtRUdRcxgoPlfH4bS6Xc1SQ3pOV3EBSTRRjbQyFGjRX1Hr2138if4PErbDvERCaCX213GyJfxE
ov3Z6EB9zU8UJIGfr06I0tVTsoVygQP8ukbUpBf87cj+I1BAav6P8ViNT5ee8wY3PycNRepb9dU9
m0iMarIUGsdtomEVekEXxK2FR9or6RuMxtshOARWQcybj5hobskkKkC/zSO5iFWOzcjSthGVqo7h
ymSZqiWGsboS1JWo6+FKnvQmw+s/F58is5NBh88Ypfk5Gr6nLr1hzev2UPjOdijVihOAlsfRWEOA
Nc6ATVrRa+EDuEZ+1NMU3YXl9pdI2GZiGmSxU/Gi7NbdRL/pI6P83t8D7kjGdV6X1dFGdV7U9P04
rrDRVNO0rKgj7tc6+80jj7803UdEcPc/3F43ALhA4y8k1FXiXw2JjaxblFJuGxuGDCO6nJQA0GoZ
pSvKweb3RJ0iRcauTDlIcJf6qd6ysAX2xc00Cg1/3VlzbV+AJHVX1Ftq+bXHTX/eKp52dQ9z+yh0
WuzpXJFsT+aCysfhKhdtOOgnlIbphCP08RC2ADgZddvmevQvA+FfmBhMn1G9HB2WFoz7z+nKfRcW
BEAdQF286v7HFY0fKSZMnXf8E+vph/TpEPBFfAMXmC0of6qCBXmDZjRToTM+gFy2RXHWCJ1Ph829
VperlarbIorBRU6ucvvuagcI1jdCGZ+d8OoWXrr4JaL5QA0ko+/sPU5uLXGWjf2LCQhvyEGhwSxT
JK2OhgSx9/XBWv45dQcRMsJ55u8V8+9qqgbG4y45uEhgrSUJXzTSg4s7/oTVzW90OOU4ieoSyU5p
nJDsgn4/o8Lqs/+BXd9zdsjMPGOR39QwnGXSGCmuLpFrhWIGufVyO7RSSm1sL4b7Tbdyn9S7ytLW
p1X84x6XW2WtNa7bfXaG6snFbNV/0ZNpiCpkuJEBNe9GAH7zFo9oBcwzmfxeqX6cuc0JVUCh81C2
wSVNHzibdx59/Rj2Q0Df+zJ2tgoxm9y595ucivMU4FU3/mvzKmdaIes+YJdHPQxss9MQAx8tuftS
/m+UwoMNXvicMUDE+q8PTXNS7LCH4xgIvOtxeeobH+Z7Dz+6jicQKvc18odn+TdrTnruPWME7Bk9
efjdRNxY0xJ6GGDNbCX2E2wrU12kZd86Q/NS/zxbISd3JVbAYo9LKBe8HCgHYc8YFDmSvTSiS7U8
8U+i+4ZUz30kJnyvM/hc0ACqq/m52TBHmVrXB0lOtMZYKB2aZadUEGF6nqfBsAtAlj0xpydbZlvy
wrygesqVzZ9g1DAPFCSFd8eRsF+yAcp7/VmJemopzYiZRKy1D2bMCF9yRe7scLML6i2UyFUA4ENa
jGyI+4iF9By3FKk+LKYKBa8tEiM2uAc0XF+QUtau9lkYffSUV7EiOS1ktaD1IVcj5DBnauOv3y+m
CSctgomJqFLUKoZOsg9m2EqEHOZXF8pn0fzQMWXElDdfoL0KuksecXCwCV5fpnJ1+tJsqGWukg2s
v6Xo/x4yZIgQ/SfdytwxAxEXd2Hqmr1vOkmmDxiWCugaVq1Jfxf0ETUSp3poJXWAyM2B/ViKF/x1
7hzNqGkvH4GH3TBg0ckYqE/xoJtEv2zDzanUFVMwVqzNEy6+0CgENI95eZRA+pE/ByE9cAYGtBh4
S3JVYJz+cEHCUA3Q3Oi1OyiOfi6DIF25SAL5JsyHcHG4tXdZFuFqP1P/1rw78rjd2+d+AI0qdzCX
O0X2twHxst8M3Hqt1GCzplfdApoXYBx8a4YnZPHgky4cAocuCn0uZjhmBhP0ymxf9dRaKLuyWmt8
NgZT+pVi5dYhYAFJBwDHGWo4BRtVaPjT6Bcb9/IVyucxXke3ZpLjOXtxYjoxtwks44ZAmfzLAp4W
7nc0jRw4Y2F6h6cqstz5SFargLPt7WE0Lj6qdUwG9cCdVzF3CvOYg3yP3wZz5lytV+GuY0DbQLP4
xnohyJ8ZbcY0NFHjJtdHzv7QvS5rvHU7o3hCEadYans3h/nKowUuqg/tNEwNv+fQPABG2NR24myh
Dz6yGgTXxm8/h2GjzI0Iso23z89myxQNeWHtLzppIjA0i+9DjJZD7VxTNAAE0bw6Qb9VUEi8Na9c
iJj0/IhUBlYiXf9EEY5dRdJeX0AmORpKc2YZO69jFNYInJ09OOv7KgPdSkPByp6LlhUPPwZX62S3
LOlj8VWs6R/UUVbrq5tWUfats9a/P71eV919kuBZZd2Ulndq5mU8GKw5ox6Tdaru9yk7FgBe7n/w
eQj6dmTny/9b8sqAdomgWZcBhz5PY3LbFdelX65ZobQp9XBPzc8SaELsyzhXK4qWcO5sDYZz9Jc0
XPXN1lsYuW9n7rN0Y1Bg3v/PBTcWmRxC9fY+zYRWPOfldhDCRwEa/NzcyNPwnEwG4SANNLX71xfp
h40xDK3DJ8VPG5yiZ346mjAPg0ni+tkj2Cq0PY51B8ccKMUas0gV480Wl3wj40+Q2Asbcf0gSlG9
qugjqKOb91XW0pqXmNZ0wU2ZcHaQQd3zIMyUHg4TfFhQ6XjKGx12ABblkHfIZKPvI9lvhGm+1Piq
pdXxFA6eb9LpfPCZOsIC+z6C5d65dwql9NBtuwN9AZy7ja9KQenWwoIO1b7XV1p1QnzeZVaDOqZQ
6e0MkzAnuGoL6FLSIZDGZMWDXpPofy7WN3mCpjhjQTF5bAz6EOiFnCnueIrY6UaiGl9PF7xoILeZ
KNAbSYeWzLtgLEM4X6kjbSgKO8qVw2+oCSOBcmhxR8Pz5c880e+TjDO6Jq5QFCPUrCI6loM+zh/H
/ZrYJ5MJX/seP9SK1myUIqbb5F3yLm1h05tYj8WxkfbM1+YH+QW4WJQoB4QcXj9VAJb+FtR/fRm7
CRRE1BNmykUrBF+4UvyxLm6GeCq6vD+YW5F27hCp3Ew9l1+wl6KSGVzYxemCMmDiSApEpwCJB/VJ
2JRXfmyDj+tzr2NrtuktJIjfEvy42TRafl53USdRqkj4RyuwRkrrRIkq2FWuMh/zc0SokltvOcH7
9SYXkDWgaH86l2JZTYWXBQ9LmvtcRQ8bfUgjsM4C+a4DcXGcPALaGbikIi3aeci5kC8AoGI5jr4n
TD0aE9uT37zNkGUgAIXrfswIHfb9tYUsmG7LGVc9Y52pWbfIKnnlFqamtWTsT+h5Zu7opg+OK5EO
woBXuubPcsIaJKK6X91EjnvFwwv1kbtUHiftZYw1bOJ3nDxtVBhImCTzGaxd8nOrNJjtu23Bk82A
xPsYNaPZ66Sk4EFaDWh0B4nRjWOxcpIBnsKfkoEw7urBa16LLmyP9dGuu1n23OL6YFvilCvkOjRe
Uc7LavyZyPWDyyKDJ2w/JFU6DyOgL2ydDVTnOyBFDw6UWggnmQJNXTkMyELETqC3v1U0eCkEn0oC
g+XJVC9b8mTAzGMaLzuiVcKahcI0XQ3rV6D2K+zYQw9ZcjGMoCbXzRx+8l2hX3ATaUz5YEzi+aGO
plT8OFhOGN+Hot+ohHQbwwPc8Z0i0bqHEXkaMraa6dlCk/kM2DoC7z9Ug9x95JRv5geTwUiWV6qV
FMuzdjCzWv0QxxHiIF9oHtJRG73wK6EDYHtioqfNwtAsoADhBgVwZ5MCZgBYaa5rypdkqdIFXGFq
UkO5tjnIZonc9Oxf5bkIct/hrvWP8Q6YuAby7CQWkIEjCIA/X8pPLTBPrp5T/1BRyz2bYeGT6SXX
nw/5TYZ+lD3HFIAuaLXdt9j8qXkuKvCGZj9B1DbY5z3N6y6xV+H1L/hs8Z+9uNYMXd06M91P2vil
Bva0ElCexe2jMygakHGDMiGAdzM3FjhSPAcxlaNNimRfe7IrZtBA1MD0TmvDjY283+ZG4DZzXO++
zYgToL3gL6e4UQDxGh2XcS9ViVh4y1N+2Zy8egy1VDhXGcZaPiUfgRMDi0rkkO8YBEahJdpvq/JB
HRH37NegMaYFcLoqIeayDHTKcNyWnW+WNcEUwnro0jHwqOfYLfErraiOndO8qFPQ+Np3fq5iQiG2
AZYoK8/fFbrEvtAKIYXacNh3eeaas8pqfohJahporR+0LZb0xWu9Yf1PCyX6JzRBh7M8VnSj1gOQ
IEaoW7Z3bruC2TQjBZe1msFqBN1BiRaE5jtpaPIvIjzSm8pe/jJokYtnQXNdWu/qAEonlOzAkceM
IVUVlA5FBSo/MK325lWa6G2HiqHNY1qMQ3Lki8RfgJhsF+PRClUE4cm7k/tXaSivdGL9MyHTPm7U
tTWrDSovhrSkz1ik0frUlIclC0RnMjfVIN1WatuNztXADY/D+35uMk47fbddzH/sfivFwfLIXlUB
lRhBqZK5cDJAiCZAP3ok4lBoGvP/gP/kVk8s1066QN4Lr0b1ckF3ljKynjg3oF8wSdK+TRhF8RRQ
FiG89gcy+l8SjJnMc1y41087kwTmnivL9fPgvI2DLSPzwkcDFEYKjk8trFPUy0mmM89PJrmOWvn+
3tfX+82xPmv0xUEHnYzbWNiAFjdOu+n7WV718H50RKr15HGWltxNdFYI6qdWsQ6MvwqGimSLIHg7
jlhtj+G32qW9nle69X5JaWhs/jbCNnWkTCyCm9S9dkWaN+w3J1nmygL8b15Y7mIIQHBMIFgGjQ8r
DLeCaUlNo+cyP+dlRHhq7BUtZ/icqKxZq6xrgIhWAnwQU8DdDV+iNlZnidsV79lERZQYFg1SoEpm
IzZ0JB1xpGOR31ot8My5YlZceIIOF2vx924QHkLXzK+i4kPJME3Iy7VlXFZkZFAhuPzJjrOpIjU9
ywxcGJYAs+zBwzUCn2d0mWd/rM0+3dGEmrsWJhlEaQ3qO4RiImaUN4+O37A2T4zzXGIa37HyvKl4
kaopHqMvTSfBEniOpQjdVcIz5bTJL3sUS89wRPpJcHTNUS5bM0e97li2nT1cEAuTBxRMFbUib6wZ
uXGR+k/M3ZXVGToipAi5ZRhnATdKJGkH/rhorg7yLx4bCx1cjjsAlg6eB79UyVtLtlGk8mnCtKGg
NYLqT1E7dBmvTeaZzqU7gV+8xlj1SbuYZyTR/zA6divf6SHQaywz3GGFLBkAv+QZxy1eSbJQXigh
mUQFtQehhrrq4lWhKflGoAjROCwjp4OefSO/QycntwUfeRnwhcyGFAB+0U8eRb4Rkv8WXq7tWXhF
3MA504u+EREwZPwZj9Hfnu31DjAZgRZjbdQo92o1siI7iPb8VnY1IVt8osH0iqpCUFNM8jNxrlJf
31eTcLkR9MwDgrNkKeAg/7tRFRpsIi7Hps0rkI9PcOsIBQH27ePdfQqRB9SkjQOAAgYqf+FsxYI3
wBzTMDSzTldgR4s6LWDJyayBOTjB+COTL26pwB128dslD7y1gGSs8wHakdJl4Hjo3Wpuyo6vSrJL
PwXyD3X7oPOtKA2kKHkKcvpQWmmlc5JkTtyyZLxFgu0Xro6ZtldoN96O3LnwcEYZibsuII6nhSoD
SpigjD7scHMQhF40q8LWWy16Fca0mVVC83R+sVHiKEUVlW315UuDYzsr9NuWbIFM7NQGF7Ezz62f
hEUIhwblK2jjn9I6QyULTwZlI78BtonGQmGXgmG0Zk4DV6dEvb3YvrOweuLAMfXc51ezSpRUkAeS
P8dnnNIYSDBjokP+oVJ78NC8jy9mPTf5a12MXY92Cfn6b8utcEgKUIuf5//oi9zxUP7gnaPEBh9A
sOcX1R9wPQu0hKBx5GWM8sRdo/FVXOWTBnNjwfZD5ZtALUSpneC1TWg2mioDeVRRJgrFcALdMZle
IfJQZpXEQLn6ZwU5218RkchK2JsuXGSwi2yL35OJJ7rEUX6nlLS73aM+LB30pMN1HDDOY6G3vtO9
0fTrliUyqZL+/31uhgufYfrbmFLHsc/Gcu1Ez3mk2x6g+LIeRu/+ZiN5xUFyjFs+wR8Xev//5WKr
cqJiLYloSHMXVBxcRXX2VgmLO3XWa2AxuiqhMjkir490rWx0km7lAWoo4vDxYdZen4qE+YCnFhuu
yLmJj46L4nfVVI9ufxFAipKP/ZMdN7Lgv3DSw8XVZeuNTE6+cweS43q7twtCJxNRtMK6LXwDTWqm
DtcS5ZZhb9pxpGF5PoLokAJvW8ZB++4aG7hQwzOZojYUk7/WVsCmUk45zZR9bHmv5WcR25LWhkgy
feE3BIJr6eUdXMQpmArYhsUrEogebEFdWU0oN2H27vKJr4dtO90xlr+HOT+aGVdqOUNgMGuCEuW2
ENTeteOWK+dVbFAvZtf7cFXDxPLS88+KSmeG/BkKPPj337a8FUfaj2pS49Iy1EU8wMKA6XweJVFe
6W8IjkPLwXxE6mz2hoMm9aviksrfk1qG4Q4ThrZpxe9xoJZpw7BCN2yIuJeyYWkti04ienIRGww+
dkYJHmMYyiRpEwGwWoKJpYNP4RXzDhm5FTJeiDb3Ba8ghtU8iqTjpnvKd23rb6Nx/PrTw6Bj4BEL
ZEB/H2A16DuVj7mFtluxebJ5xjMx/vlHnVElB/cNQIZAEJ3UnFgg4FLkCVn0SOYb52aMtHGoCBBO
o0UPWqnzJGBi9bAhVZU9bh6/TCP2FX/GZgKx8uUjxoyekt/ZTbQ8lb2mfh+5NXkyPFpscnMqygHo
w/3gwOosATTI52XooW7DgSyNwW84g20gtdPAbhXMXpRxx47WCbraUCbHNoxqFw6QMbjDOeDQeAOe
7nJs0x8GntrI0WGLSI7zHEdPhqVVS5jSyf/XajXcC+NsWL8CB6zRpJS6pj0g0KkS+VWOewvBuOtB
dn9xq3plGKHXHWM2WvIdiCgB2G3wcysRkLp1dpKVvyj0zez3dUJ5xOfQVkm0flfcMdtyOVGEdB6H
XgjXPnXs2Td3mwQS896KZaWpZXzkaMKcRzk++8TyzMw9rnFPRbKBfSgfHZtMR8zsMKnZyEAcoI5d
b3Y7+mexVoUkWLgl2VH624ndlu7/Fz3znh0iyvE/l1VSkAZFeHj5Sc4G+fkjFb4sFi43LgpGjhCx
f6T0QCTYPO4bCP6xN2uk1RwvkIh65Ap+AA6teZrcC7jzvM+hldPHTIxRglnVSGqL12PuLp6j7+Sc
5L8RlcHFjTsZzA8qn8lhHOe3ZJMWv5N4Shmt+kcWkxMcT1XiEfVSXuhOpRX5s4ET9pnnwODt/EQu
JeJ5BItrj+aS9GseXRLMqIMBXFf4tOy7pW2XhNT/yL7FNN+MG4v0UAFC1JSm5EZSY3GD89c5xudz
bzHIq/DXKgJKjYRsxnEA8s8l5rKjw+uaq8k42BlgONiaFzjGXlPSW36zZJzO6i/iSPFDGnk2VlId
Arp57Y0C4BrSInquDTx6eQEw3L44IJ5MGTjsdd1ODeMJkQZGDLtWbOSHPAOxtECi24LO032imUB4
moOmDlMh4zoYnoMzOh3Z3RAhUQzNHNzbxuMP2I+rVJxxuMZ7TaBeYNkEp9CiuVlNFjgy3gX5wamo
Yp0j1Ei2vmXeU/upgRaSLxr1m2aJHIImxbW+iiNcWKkfCCFqf0rKPbcZUnP1ZT9PANNuUQZZfpC3
ORrZaS6Nmfg0Z/KvbN+JD95CF965NUp52aHR94O6/1v+3SoTfBjh95kJmkrQBSjWPyMB6OAZC8Xx
VvaTWuijpKVzkaQJhHHFDvkMrtCshdQnpAy+cDwuhMTGBKJeBEVufGxxGvCSjkQxnAzfKDocygP+
fz6itAn0Irfc84fuV0XmRpETRhIJT15I9U3FGdhtJZ2rfhGDbIokqaZ7nBz605AkjKQNpLAfyn8f
ZlDncnwpYj3GMwouPThEXqaHvvWStZdrP9zjiGH8YY8sbEVdvOLDXNqz7ML2idCrc2dfB0WfT04A
IPCk81P94Cr+FjvNd2gOHlCqGbmuZHenGeaNyh3uvMX87QFVRAXopgkkJy0ImHmEXsP8cZwuUqVs
yjUx3+y7hT6fKFXJZya9tTsgjyzLRLSZAicPQzRV8pQGxxD+ekfx967FRSiWOV1Pp65O7x/ZMl/h
LURJnPHyhQcjkKpRGKvFgtUEEhKqYAG71gusVjnN8GegC5pwNmCh5tantq3bIpyV2eQby+ibFdiV
HXqzHn4OwTRT0c8K4AycZq+2sOB0xDnpw9+NvJyWygbGe3vgbwUyxF3D+N2AR95j+vbEnVGpGVVt
0M6zds54meTjue4l8crLNl4hvoUicDtHqvE4RoeUV06n2j0If+ByXQmDfdJO5CfDn+qmmwShyCOG
jd/N3MEWiRifHSpXGaagDktwso6kNltblbwSC6lV3Uqyr4yZykuajNDXa3Tb6dvmZt2rXLcafCBo
yWtxNdQw33l3d0zRkruf1jr3Pt9a3Puuzdn1NxL26N7f8i3KCoMSTNOpWmCnHhu29qfz5mTrYCj9
Dm5OszKnNpi7FbK/whSX2wx/6mwegHffXtHmZhu96n3C0Y4jNhBicRifXgAShfLbO/9xqbtsBLI+
KFC/3l+56NUBhoRtghlI81QOWaOHOHipUSpTvuxFIdMZ7PjqL6AEqtJ6imZfcgrBr+PyUoPzBO8z
/XqLu6RPGG+nOa6Hb4VlNhxn4WWQZZ0ful2GAb64qLaLfTc9IhnrwUk31+LxkSTDpC2O+lbo5c0K
9yF0U1XHlp7W4TEah+nVnU2dS8TZ/8OPHEuu4KipBazzJcExFQ+FEhL2x6GAR2THl22fz378FJ9y
+3Nh2Fg1Qa9sXrVAZIhVd8VbBwoRpgdkwpD7TH5XCrnEPwRSR/aaWwQz/rDXmBLLbw+eCIbYCz0r
05NMpxT1xKThSvDNfij4l+S5NzbcrhI42e1aSH8wC8zGJ4TkZJDxRjJZ8sxhP+8MH1wfEeBvHlVg
rkig+ViCvyM8mvnTXuAYl24g2YZWOtVbyFXkaU84mKZK0Hk9eFqS5CcPeHBroYPHd9QyPY0m2mGR
qmnUV72fqrU5VEqerTVsCTjj1UaQazI2IMXSIQGEFNmQfC9SGdYC9b439Slph1bTpUzcKnGQjhzC
cKnebBzyOxCo0ykO9bj9zZEKGBB5orznfruObwOONmN37F7phiB0OCKDe02P6uvKU+MBenJBaur9
LSZimxlRHTUDynU2B42KAOtvTcxgYZItBx5pa6sGR8wgvMkIJoQywxbORY54OeoLQLTXThGxNDbH
iXtUZzeAC0C3JtGxwWFqS7X4D5hg37FwzUmbzscaPDA+IUUe4peVsWW00HgWhhufL4jJtcvpjabN
s8WkxPBevmN8xLX8XqUAmVepGvcWvgWbBU60UzSliSJwIM+AhK0TDhnLZVB5IFff6aKzYW1T/Iu7
lbrEvYac6nim9hvZmeQStGjHuGtYgxKS1IAPBCwAJI8C4b5r3nz25VJrc8Qbfiag6yLnXio+mp19
ZUQ8xk8IJx5elhP44kDRHEQras3uhd/dcnNfu6QIWUddElzUKHOLGDlOHMawUiU8bxnEWdScRaI3
7Z9P32JOLbpL4cBdxtgDcTDyPQTj4FvG7mRhQ+9cYr1VfMQlQpedtON8PWd0mg0eBeepsWLPzBXU
sDymkfZaOUtnR4WRtw5VfLpj2UmALJrVI2EegkEUFRXUE+m+kul7BU1VyhFYMPkIUsvtFkHYRn2i
RqrCQmE8KlO61NL2ib9D1x1zLEjSIT8De82RyekLxqzFQRNO7wmlUx6RFygGexlMl8qk/0MWpdOE
2eJShtxM4fLIokE=
`pragma protect end_protected
