// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
bShhf23gnSVGP/mtKdjuNX/7RLMhjg1aAcFdVoELHRD49/temorIifm1rfOjn6zk
dJ3UHREWb+QfrgTlzQB0GOFEavl+nK3H7DfQhup2A4iqMld/kowg95nBfvvJqUkz
Iafhu+lMsqMgQxIid6PDGHPshI8Aa2LiHM9Y7AqKojQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5040 )
`pragma protect data_block
1xuDjyctXprHlJJ95VspsLJSqlZN1Sz5OZOE2wRcLOfQUXhGiYGjze5uI7JOkiH0
EIoi1/BDsliR6n59kK037KgJ2Ddb++CFqGuQ2NWLrlcvP4xzjnvuOMCM3iiS14PB
dgOjNBtUaQbtdlsOgI5MvjW8qnyftKTcXBy0ieJ5hzKQgb8u0cdbwumV1S562Hij
06fHQ6Udkp06e0pvAlua5TCWQS+9w7s2xU3zJX+i+ABz2DfofLyjbXlafzDxW4Rk
he3XYHuzMZWgXYe+zOriQsHrfOlbLKjDnZLCr99azn0/AS1zu0MW+YHqonyZQ/52
IMmzpN0bKB1BLVjkZOVxVsZOOj9+4v2aBRK8uGh66LC2iguxG2wdgnNkk4M6m8DX
dZ/vh3/w7egvo1WBAEF8SxsrFZghZL4K7gmNgDyE7+L8DMIBBeO9QETg557s0V8x
3qtOpgGR2yCL6VS+e/yfRwX+xWjKMAlmX17mZmgdI0Ptxu7cdY69p7BF5nCp2ngT
tgPungm/UIpdeyVS983NEoPGcQMgj9LJS3EJB6NOD9eZGQSWByDBDlJpzgWd/bdD
MeP03n967aMbxXqJJztu6zLdkQoWK8Oct5qaFWjZOrDpFUKtN7RLzpEA/x8AizOa
vt7peSvhFxIptYl8SGV120y2yBisTFOWdQ/a6mgZzDJDRBqm5ms8z+EeY/fG5dfE
VDhKXopteYliK7e3I8UcJb0QpM7eeeYtcimMHKKSQGbKqAZt9u8PS/z708nd+JxY
cjQjIJk0b15umPHySwPJuodV19HjYHowEmDaKo6uCc50mp8AuWd7JpTNgNH/IvnJ
OHgt+3oGCKSix1Ep28l6q/YVlbukrslrrJunLRxJGkkeJkUxWjlvInH7cmGB3rQd
j5ifzqD0gOeNd4mjxsV67uicJBsM1XU3TRhiyM5eEHyEmbqMiuHQbrlwKFavgo4d
hhO9LjKrgRjLRdp5wWhUCE5RycD3h3d7Wd4YZbu366R+rKjWqx24VAbm4w4s/b3l
I/7bJCnJuWRJDRr3Xah+Qtjyqqgq8H9rBFcGmAnK6AS0qdnvG1S4kUIPkWFH8XdC
8wRwlQA4gjUO8Z/oN9KMG3GlSlnlDxlfGgbR2Iyd0+gKU0ZatzzHw4l6Vmiq+LFv
30Jd4qhnlrGH8gs0onTHv6b9Zuv19aC/BpWLOuXEAd7x0QsIWaDD4mLDj9EdXIT3
clIRin2zdIaU3A2eKApuaLldLJULdTZVuGgGyM5+0U4rTb8f8717jJhfqX0YtR5C
YgzqjovfT7SQv4iurU8qmVhBTTWIUpMe3CfkqQKXqx2/cI+cvrlfZFmqf06bVGcy
ZNCLGpFaCF5K+pFNAuN+A0yr0JRH1IAr8/Wt9d3qThjhPFXo/QihdZqMexhZKRc2
Q4fs6Rq5EsZlIx9d67fW/QoTj+fNotfo+oHrtnq03dEsodAgW4AfUJ1MHLN6dzas
bS0sMkwBWUJhX8Ia5Arkp1UJpsH6CO77F0Mgsly7dXYYP3fEOxaJpIwN9vZKA7I2
OsBBbg3r55q73ezxCjePUbb/WM5UGQDVimg2soafnzLQG8nQI6qPkX8o7YRYYcvn
SCl4uQEYCpl6v9fv3gZmVfgi60ZAgByhlYc82uuQBSa46DZ7nVPdM5dSpuufsb6G
dglYgLiFL6O8PUhpGy9AL97sYxxoWgSxHwp07fNxGlqYmEFJj0CsQzyljoj/jjxb
WPJndOzX5oyUydPFbCqsnSP3VKJGpylpNVwaR+Z3QEZp/zx+oyJ0A1xB2o+sycMP
0GigDgCrBQPKccDkqNw0Ur2M8SiFBydUoxs57/Xe10/goU0XvEmnhTzZV9niDa/6
GgA8BJkAsZ6cO9kyHb1TJXHjlL987BMXicfs71+jXsBVdw6ZVnqL16EfYuXJEUf+
favEq+P1GxG8fXBPW8J45bZNAuvvhyjcPKm1Y51xNY9+aB9O3dUTy2WEyLZOrQxM
e9ePL9rju1+v1BnjxR6l/T59oheKkzyjB8GsrVTXFy88BGVx/5x7Ik1Z74i3n3f2
2TAiWDP7/GsEQgfmKmaOZYwFs98qHM+DC/7VmN5NQ6YIHEFtTFMxkv05WK/8n5sp
+eBM6D1ZeXvCZCMX3uI+7Ofq9E1VTqDKmzlJGmKRhUH8VI2CDvtOtXQhG73lsPvT
/1nMRrZrO6ALN6GNsUQQJR0zAfIx6CQ1r4slhU17GNUoeC0NbakUICetQ0MBHwwW
y//bdg3BQYATVfIZkZSEecQel1uNTAPV6j3/uPEGzkDYywidpV3T9YjR9ygFpJym
KKRKwZPkY7EQxRXqL9TwqZGYfvEuVvSv+/XT5qw6M1gPws1HRG3BfLORo2QwYvja
UHIVAlmwCQwY30Adl0L5dgmcwdMURWJIMwYDkhDIxz47ZBdqL6GLA4ns7eKPQd00
8o8ghjTLvScBLsrRMoFFugqji/gFllIbMpPQOhfZU49iFlRreBLHpbxcIw2hFixk
aRXmF52EjAyrY7rqYr/m7wfiUzC3dXMMiDoo7v3WAgeZZM7CBmYHVstk1yBhD4Kz
T0LTI16l1U5GIVP1bvwKSr+/aNTdvlbrihgdMGUsUHj9NGCO1A1YAo93LjLLEb/Q
K2aUXvwS07xBy5ag1tIkFhqHm6F7JN+xbECbBPk/ai2aTsuw51oaFh+guqjnjM3b
kDpaqz2aQXQGTyDuR2n6ke5usqo7PoHK2lPatwxS3CgqX8ez3ISYG/EylAGyAXXN
eHp8Qe8CaadnB0FIpYuLVi2mACWdIWAzbVgyfS7RA6Z+Q0d1Cwdj3XW3G3527txj
YhjmEzGtqA8hs3sXOHTO07GbNIZ9ddcvKYpAktfwhiw6RTh3keSyQQZ5a6aBV1nH
BeSZbDV67NHNo0myGrT/bOlqKb9KTW2T0M3uZM9e8PPAv9NhduXJHhGvT88junug
7XTtkfRA9xtC1cASt9eOC4nC2l8LUxvTdpw7XId9VDiqjWnCJSoAybZw5VKsiVSJ
/3C/R9PrbiMlzufR9+9XAGhr6lM6lQS0OVx2JxS1kr5TEEYJi0QbKThfg4JbUYNI
L202UKDnyGKrMc1Toc17jJ3B8/vE/polETMuFwS99CJ2esBJlXk79XiiYHbzQg3/
f2aiDGA5XlcW7XjJqdGJXmRApx5hyKPE2h0ZhT9mr0DanHD+U7NhA3WdTJk/461B
9Bkh3sCcmud0xgOiiafPF5CNJpH+uciW6N8fKXOUQGbDYlbHhWHazkzdGb5Drv+J
GaXseVFMeWFH8kPPp2zqcLGvdIaPyzhbhQhZwdreqpaoVRN5EeW6Sq0A152JXmMv
XvwGDnnSZp3/3WBZihJ0fB/UbS6UTwMjbeLgnY9/YxTgVkzItzN6er7Zf52Yb8E2
kgB7t9ZShg/kz10svFEng/VJY3Ws2NXFJRxJM+ds3fDREaQEueG13PH9LUuRpo1R
FqOCU7px/z5H+raHwUAsKI2AWc7JlYlMhgNwK/ifnywUFSQoCK1SSv4YFDVzm/kY
RvQ83NoKYovKcKPi8RcTuPpseGcrISENm7XN5mXx5PCZ0+ODsDJH5QR/z+XX6Phy
OpS+up+d6gOhpdDTbpMtu+Sc4S9GM6O8njHernkwaXmZF0igSIQDARAFVoJu1SHG
tNQQFJ/Fu+6JOCuTAJrGNwbaJ70O0QEmLnST9L2SN+/oFVgVroX23Q/F5y6iqwhp
8QO2GX3FONnmNg/dTyAbUXZ117/NV5N7tpem76mShud4+yB8cm/1gr9U5rQvSogn
RrxdVhvOJHBYdViKMerLKf5NipwZN0jYqmHnm0cWXq0ip7YEuEOwV/HBt6WY2CAl
nG48PU7ETXKZ9UmoIoboMP0CLEHZVeDP5wM3L2gIz+gMybl6K6gJ+vbTKezxiXPx
8OpoGvMqiUWab8OA9sxo8bYXcEbVAnQlUnpPmjsmoSkryfP+TyNzNSf1Hb8ZKq1g
TDbTN5pjAfcL+/7CAZuKiGEjlTphUIWyHK0SdyLf0hf7gWOF19tM2CAwaATv/Lx7
m61fa1WJzowUT32wjv1Lh0Ag29F7GsIAwjTLWABw/6zne0lmKyEdOqfJ+Q6YqNGg
uLnReAuDar4+INbkAa8qzpPWF/O8EtLIyEsF6oBSPNd/1NRVoXFEE9lMOr+HTK7n
ndOu0yHvh8ThYT+J26qzs0bk5JRp5dad1ZrdFoL0KYjBN1ctEK6j7LnGZA1pIra5
3er4zlK9pYgYAQISyyvgO05hDjCKXl5+ZiWcwrQB4lcNqz4V2GyvmCtA+7XgziAB
SmnLRRgux+qakIJIm94ere4PuUDMc63zV+otVkxO+iK8spPmV+IjoLuaTnIMpwpT
uh1f2Y4GP6IJAzOxiaLTK6JL/pN+u2NckEwdja4pVpcHiT7mn3DCCFFgKU0I8xPl
AQzN6OG1Kr/oEv9FXWCfy6xUGCb3QNUrbPR010Ed8gQslYcONSDW2tkgu7jjte9L
YtsCwV9X4uzR+MKHPKQ7hjJdu+DpJaGydYHV/uHtEkyIKmDxZQxdF75cWwGYn5FW
dEwJ3gD/DCGvg2Dt0ZBvP5J1YL/WCMmKJ5NkT3aI+WuZmVY1o/G1EyNKtHmE1XUD
KpgCfEEhOburcKpTN+W2tfTSP1AIn1AzcA5pL/pElkH8mLZsjgnIvVcggnFRmEI9
jL5UU8q8cQLGhLc0eRCKj0mVTzwXRufLpks5rWdIJqVyPyF1K+pfEnH24LfMo2VX
ErTOnqLw8jxy8LI70D9kU4SdHsFqVWI7aipgIxj2pfmBHBFVO95OX79T7H38i72q
gGk7nr4+OtCxbKMHpk+4ps4Rx0fc/yiLieEeOUZNSOTzmi1bQgThu5hcRTk7Mbr0
ZVEOIfFI9LebulczbW+EIR9FaYLfTo8UqkahFrr80u8AlrduU47GW4+ym9kA+HoO
tIHaf/00PG8AhAYdS9A1X7ySwj7Tpcn5CORKCbj6ZE+1cyJv92q/mW2cHHFs5KXa
BvZM5KxNlrhlPJM0PlHNnbVYjSBPk9zb6xPUdFPmBxwS9bW3LJVLXWbC5Pv8807/
rXD7i1wxsGtQ27JF/Kgkr9FxWo7QLVEErSpqybjMQb3+zOctTw2rW4zz77SBbIHK
G2iDr9pwV6pzxES5T7SmdoIZneHZ6318pnNbRBWlW1HByZzvtceq+ED8lqcuw9Uz
4awrQ+QMnkC28WdDwgu6Mm5Tb4df7tuPzqv7CLMBQXt0acP7b22h44Bsf9W4KPg8
xguoRm9+o8vr+Sj9gxGHV+EXAmIx5c99r6b1+Vg9BANyEWCGM6AT2b9R6MOPtxg4
/U+BHS8ONI39ZjnQ68gh2XKJJsxnJsfMkOXe6gKOm010z/WBfNLPtqGeBoVAqo1H
fTigpnCAZTtxFpZ+Irq9FmoYB/ztDsbxcQe3g23mgF9K0BHRYuxF1jQHXURTsn1i
dnntTtU3z1Ku5rWRqD8cZ4pTd8tqxR4Sxfd4vOWredK9/aNsDGufoI3l5rKZRa5u
sM4R9p5AvF0RuS1IDPFCasLymkUFQTuG1tJWTB4nLgjJNQb/FiZlYLhN/x88cPVR
ywqqk9gRZT/o3kfMQsLAFk7Hhrf9LIaxNvg/5JM/EWj1myKwCKuM9+wxW6Vfbbbe
hPymMq1mwhUYUeNsWldYorYvEHTyEgZClRKxEZbOXy4zCfyvrQyy3DWqtrRxrQqo
u8turVHd6PysiNykapE9NTmkQqcyxpRZoDij4UyWjouD61qP+rD7/jyaMFL3eyqU
QTG3odz2vkhHq3mIFiljRWACFP9YzQ7LzfvQrtLxSH813lTpssoXEmDFj3f3+Wd4
XASX4rAvR5BfruJ9EwQ2igTrh7xkTCXbhrzYjnyxhmQwwinK9b6uWpluCXpt3wQd
61r6g8HdVQ2JK9begSMbF5kKOOXQYdPpLzUqPCQgqe1+eJ2ss5iJ2J+Xt+bxxhsO
PfRAtII0ChqHe01IsiE9dVp3ZeOf+SSIkfy3f2tk4rfQyvVfr+AY0HNqyGCx294D
voOGEaqrAa/Zh6GgtfCSuUf5gahu3ZUeKBZ09CMelQBBlpzIzh7fXHE57LOkcJF3
tEe4MXfWH6/+KNguhWS2+3Z0OdhfGJiKxDgJEJX691T+yb69Yok9bp7TyiLsJht+
Tm7/gax8egdlSsDdn6ZuS8Y1RCkynmzkmkxgbj1OIHitKRFTtU+QmcneFyb+YsbM
mX19BW02tRueu9UyOJqmgFrk0F9KMh2PPbTT32NcFOCC5OhkWvruY0u5CpNtM95r
eTmuqxRTjHPynx4Zv3D3K58aoReL1p7jZ2eMY+T8wVj1r3wOjOO5LRfr1k7RZKl/
tcGXTwRAxzdsD1KVahHpQkErHSDfSJTrDcWSARCtxMzKVCocmSk91na4wjd1w3Fc
oDUEFS2AI622aWndELdytBUwzQjXyjtGTbYszPPgoU37rG9zwHibgXW8+vCIzwUX
H6fmRTsyVnlbl0JstyKNNri39fMhKMX28ysxGtoFlfAsnTE/VjTy8yMKi9+7i5PG
SstM+l1KueiAztoGKB2cnw2fxVnM1e9ff1dzGODXhSZlqU+yeqAr/CgqLPv3tj+d
tAO1Q2j+VOR0iLA7xrKSl9zHVXOGi1T+61Q5zjo7gyJ5InbTz2wxTwzSLtQXYEa1
Kmo6hhsjRqfXDts+d4dJ/YjKOAkEAvUoRJHL42HqNUS9mRGjPG8SZ0cyOJ7sqMWL

`pragma protect end_protected
