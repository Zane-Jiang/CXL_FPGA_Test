// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
THuUImyjwm1DDFfl38jWHfe8ffdDiAuTTSczLKbydLEENJ2xgdPqlgMwTWMa
hAGr8iEIgZaNxIOeJyQEh5fwag0b1E5UhnZGANWZ6L0AACau/YgE5OEPHfef
asw690KUwNH7KVtnt+WCTsZ6uwVMmoCBmd6NLCrFrz08A7ZM+ZnKcbECmZqS
WBdN9/HjvHEpm72nfbAIlmMURs5XMWlVQqv2GrHP5iJ8/jo8ZunsxzFma61c
cfUT6H5ALSwIklcdp7HLAjiNdghYx+105yMGmQgF7O//gypYUT1UZ/d8udaF
bS1HReynQQ3UfgNY8jSbQteifUCxb0ztfdap8I/WJg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lziag3yWnZtUlLm5u3Lhj8e2jsDZwUQEjM7YNFhw1jZ9+DaMau45Y7Uj8fK/
MzH2wXHY4SFAQop9IpLIGlOI/VXlWCDL0q9FTE7iUjDLLbx6cbQh1Taj/YMc
75QZIYBzyu1MyvpVu0O9quGrrKAh/3GVvo0/tOkItssEr0QHtKgNqVOz9UOB
cdjUiIhPVLOs1FfTcJm0adFgX3aGt0j598pf1TTwwX5QdrO2zA0jGKAkdqWG
wYArAGyL6NJQeYTncAS4foe6zOtsYFdSPKieBOTHJgoc8DAgTATr0XgcTK7U
gUpGlim93coKTu3VTD/c/TxbhJoQQo9eveWu+P8N1A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UL0m6E7bpdVs6BDTNmaoNw7KyNG64sy4C/Wt2uDtWld+Krfliu2HOZTxc7bI
LsLfDECp+7ND47Hf7sPxyptMdXPHVgWsH5Otni6qySmurGbLlKb7+g/i5aBM
r15tpa7bIglVMlAZZ5wBJC6O0raPzmZdVhNxWUH1MCbJ57YMTPVzAZE6ATrT
Pm9vvdm6+WULBYUzgjGGsfRDtwt0HckFwfo43DbDqrLstN3lfOKzSIr12diU
ceBFpcnjI3NTmMOJPL//d9VYOlYbCQTvUQ0c0OUT+0xWiPDXev/4HnWmQqeG
BLAzdPB1j6z16YdYQcMvDAc1xP+23F8PxMlCc/ax1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qD8c/JPA0MTi8TSodhU6wymUE1etUcPiO7YIsU7KtSviJiPDHcoIqbghF1DR
usYB7u+7WuqS0ING1DRG+Jo866qj3FmGWZVSEUmbvIrWL6jh/KRGY912OFkW
1CooUMbSoRLJG2vRRExcXje8TyxVUM9ynxu+/DxYIEjUow+kmHY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FZTBVapC6rgIsxOv0J/06ETNlBKodmpJtka43vaz99o9oZnmoqbxTpR5rdqB
rUr3lT3Qao2CBTnJBlD4C/63927iPkF0L7R7ztnXVa7GNP/ybr9o7c5iGMvV
7EPQy+MsPA8U/JNnaoxwDmPjzqJBmkwyhKL7ZYsaO0inJ2pBCG8vSHcqpSxR
sTjNi08oemkwQqtYyUD1IfLiFrics34mVgbwoF1SM9dPylhn0P5+ii1yhs0D
PaMSRj0Mvff1azJr2S3BeVFD1B9pTF/mDYTPJGu9Np+v56xBSV4YZvlQzvXI
rvJqVcbun2To6GKa2e3xz+ol54OtRoSrELW8fp3ilTUSjQExfLGca5eVeT4E
c3Jw14+OBVrNWzqXg0tbahHlc+8FQXkEXE1FJIld3JzY1lfpVRwCVHpsoy+U
8mLlGcTAFElwYGW2T9QhevbkCtIeyGCCcAot00Icc3DnuT+hwYZIfJBUO1Of
em/ga0CTq0hyPSHpsQKWmPbIsGTK2Lv6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kCW7dgYWvDUcEUI0rqP5yDc74l/oFV87eUKMSt+KjzKR13+I7lXEjAFjlmcB
IJwPjlM7ApFe3ibTvG1yRyv3+6/2/d+BjwM0Of+6VWdEdSWgmKIY0sZ0Ri6F
ANkbF0luuNaVW+lWQvqCsmMI0BYXXM4yIGnGIMVO+VsdV9Y97Gg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Z4G+n5/gP5T+0MLNiZQZyHJxBGsDApT2pdZbC96vQX5Iw64CNDlTbKGDjlMr
BdA6JFtygwYif910ggokTyLji2rETlOcFslBgtGQ5lRwp7Szm4Wi+Dr34HsP
I2zBKoj2K+u3dbp9kItex1RBSJD9XxcoSbntWSzDbx6SdnD6Q6g=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2519424)
`pragma protect data_block
/i1aeMGQ8oFuolv1qHtPd5MkJVk1n3ZumnjWTxg12GR+55DWuWyiHrlHdnDk
5FBlMbOn7fFr+XFXPDYhDcwOfQ6q2jyeZSXVcHKc5l9qU0Hcvws3R4fQTL5j
LDtbxfdgvdqg5jmwv+pDFaodqL0ywqtz2Cvx8PItClmR18BoEbNoKE35sY7n
THZipA8vADt5V1WGDIbyw7O/lAGgM5MtBWCk2ElX6ApcWZ3ruuefgJwUstUm
PPjJ0TPFSujIzXVay6MaBjAvwChAjhM1bXJimN0iu0GrnPgRDxC6ALgCq5dI
rEJbPGn+wS7gg6aNk7J3+ctZvFI5ESGyYb5qa/aN5PF+KJ3iw1wB8gwYJ4aN
jPTLPvobL4Uk8gC8S1XFqbjQNgtbzMF+6kzPKLTnuKF6e8Kbw84x6/fL+DTK
WNUc0XjbyVB4TJSdvzndJTcWUjhrndfiwAXNvQnw7OHSs40Bkg88JBPkzW9V
X92SSScwmC5RM+RTy70yVWysW1Qe/xB5daXwxET4MB3SQyCaZqIYCpvzVh8b
smDrGyvSDoEdKwFuaeZKiJXUbvE7fF/OdyPxp+diT0HHMCwAYdVyc1+WSt5b
QJdDJPZEvBAeMghuopd/1MCpWepXyKcb/DwNVLmOaA1INy3JcBlt47uIh2td
w7tZcr9eSbcnqt9Zgxi7qyN7w8NWC1zAX2yIIngwLSkICE9jYz9nrkctc4uk
Ys0Io1UZOCu584Fi+2ulAk79k88H+abyi7oQ5BxbSwAXitFlnckIbm0k+Gtp
riEI+t2BK6zpPS7Pq3YAXJvo+T2uagSkTqyfKXhl+DJZwv7pqgrSZloR1FCc
eShh0o87UnM1LhIZBVlmQVPM024wqZ5R7XeZbCRniUtZV6dOs9hZbPgoR0mX
I7iP1GZhEyJFAPYGyJgtCRS9ww7FtQJWXr1++Ex+koyX6j5SHehzQpm5pCaO
ncGHP/aLZKE0ZYGi+b3h/zDWqJjYOttfRrftLhabE370Wh/+ADaUY9cNvbyG
H7NVytfBMxABlfmvvH2SHExslW/9FGpjmWsFCjfjEfsMtvbBbHv2rlsk5anI
Pte7OPtBND+jzUFhoUhHOatZXEogafls8gAYhkstDqzW4yOY1zCxCVWp001/
7NcuboxKuvIwrXXiD8r6ehJ21oT4zJpc05baTk85GYfmQsXoNu1KioASn29H
tyHNtiYpoLyWyu9qHCU7K0ImW8TyWXlVKz94Fjl3HghfcaKMWaAB5aFi3CpS
zSh8/rSEHJxCyDi8g+Qx/Yks4QSPqd2x8ArTkC7Ou4gtBv7NU5wvDItRAm1A
WTWSlFgUzeFAruFyF8fz3sOSWns0xZ62JVWEaGHcPlDZlUfa/Gy9k+T/LZ2x
QsWl7bnUUx37933WPcOuOruvvAYd52PSpyGRIuYgvVrD6bNvlfOzpSblnZsN
m5NXhfe6KW9QrJHpJ+7DkedvMPzpFimrMUoVZtKt+u6w1aI/WNRZbtGUfWV5
IA78leDyJApiAwGY0yYfnK0HDmJYlporaHiABoLlnehq4u9+1O6DlltVyD0r
nN6rwF1eQDgopf2SUFHuoHBf047cTUnZvjYsZUS6Uj4FcKeED/oBeKNACuxx
eiWT0iu/iIDfH4+cMHQYrHKCHeV3IFHkWBOgBMZ1yTk9/1vf+knPgultwovZ
5xt9K0eDWzNxppNmR39u9wpfYC2F+RwwqDMgPOdx3hgWwwxhj+QUlIfhN8xf
k+s3Z1t37HrsTXROf/8J+leUVKSGMgHyhSTIWRus4UgXRn9d9MoNDD7a5TMJ
iobOV6RuwXddcno7y0XUvz/abfnMF0JbrXtGvpd9ND4VS1oGb0DuglsrEto7
reNIXS5aiOsu28TivnX8Z4ApfRIhxSePcChmMlg4E+Mumbdg0rHprTbkpQ02
2bsInQtWOSLRm+4d/GJ+YOS/vvNAjYVg4Exsgny7F9c1W2RRHlMiX6Ozd/y7
3Uy7lUH9QAfKQnovuxyaf8wX/A3CusZUXJQ+OC37J/Wqrz9Jwe8SHslbzRp1
kK3U8Zoh1eqAV68lomfbZ2nsbXF8Nnykn3TYzlK5qnCStBC8pknBePsUS7TH
aYdfReDq6l+JRqwXftVqm1If4/MuXW+nkU4OMGBQxo5Uubgh8XneGig7qcrH
/+hPMt2xkdhUOllmLmqgVuMXZ+UdYccPGFf5KHY51BV+3nxOWYZaSKwaIQ4t
hkniOylgsRkMGp53Tli1gTUCtN9Xex9uA7af7Ebh82YWuxSvmwxgk6hjJg/C
43Hv52XtHAqLBI2d4dCsz/t6KOnhQfbJ6/CkRKgOCCXXc521bOoBXur/THne
nwl4qI6o3SgrkJmspTba5VG2K65CiSXRoS3rcteJNUIVfGDaLLAR82UBOBxf
njg1eJr1WN1VpUAk/7YRI88XYkOTWWyORdcGfAKL8iFQXFRBraR0NkKvucXu
PwSFjzZUx/uVb2auWqU46OGT/rSkSOlmzG0fp7Mzv6rsHcoFAyYWDifzesZ/
glxYoHWeexRyUoUki1aSd3yRbcKWWViOLz8iD2qyuBsFl+yHNdYzVekxZq0l
BMYInR7MVrhJFpjq1ymaqCFoB1VBm+06tno8hiLSEucuwUvqZ52G/fI75Oo/
CjxC7D45ScNgOdt4LaNlC4cT0l0DZ81ZYHI/g3RVCW3btQ3wQtJGLm3eaN4B
FvqGvQx3jiNsVOcgrG4kqtaEys25g+Q101JF6baRrFHVI6R+dqUztN/fkPzq
FjJxwxThBnpjBgjlFAS680Aftz5pj9Oaq6MHaYL174WL1sL3mZTNBheG2VS7
yhLFULmzAcwkQX8Or+LnSbzCd/Y/zfmeLU/OIzMVfDiHem8NlWwPeLXVhuee
HvCWFY0QsTc+lL5DUTAtKLnlm+kibbFt7cwO7J/rMY0ej8ez7imZYG/VHBLQ
kIVWh8IjOdTdRCRoatr398+WzZmcYOjSjJt/ZAJFg+Y4ZZ7FcZ6IRaaZ0gRf
7EbYqeoEU+B/1hrcox/DZFANVMAGoz0DhJk9fPJ9ZgNdmBqzDFRwRKYLkTGQ
CAh/W/1hPLrHKmH2bD7T6TLMi/LSV/tKYBCuIppPIJUaOBIOaal/5CLAk7VU
6vRqplPe94l1aYUqHOzkr3jfqirNRm/azm8iMDyjqk1u+/UeVwnijsJToBRo
/5NyhMB75uwcNvYNjx6wns77G2Z/hyMgnn024ksLWmBuGuiEryTj7qxJXiGs
8E6D3gT9xfR84vuQfobirQkKLmJ3b88nHzvH+DFNRNBaUsxXoJ/BysNW88Bf
jCfZO1XM1LmRn4vV4UM+CwbZeuxPb5HTdXx1bBivRDgiaHypZgFGrYuq1JhT
LC799aYV4/KnXpUplNxmcKsm9ICTIMSxB7ta/ZrI+3MmdXIAucfxlAlZoy0L
8zK2mOWDvSfkAIEgtniTetm/B32uVSmMKY9hjDw7omzy+WyA4XbPZcYE6r/Q
P+0etAEHUabyZsc6cQzp0NX2cTZWKFlGn3H/FTEm/w8wPiOwj6RMt4D1WsZg
vN+wHu3fZclWJGsFaa0n6e19bc6iNk6tsYKWXquo4gAPkTa7Wl07pduVuSeK
4bjmwE2yEcrFi7ITJAQWt9/4T7Vr+6qdYiIY4YPH3A83NEpUWFb0dmXGfyjc
LjmmVXoITjLoqpFMRsAkNzG18OI7x34FkAtovp4P9FPI7yXRdGkaACvAEzXk
Gupesqnf6au9nGvaAjTWlyohbt/s8oDGbOZk5m7ja+4O4N3uPwu3a5F9yEA/
t2kppR6NunOA5pJwRHq4hybGozHD12l57HSHVrPem1VYTse9Thgppqv25mpT
dYiRAkvv12+62ENl7fJxStGyb8wEoWNe3YNSsOXnPG0x3cU977dwMUbtJPEI
37MNP+s5zFMCv3wqnyMpUwrl+cvD5uSnQ+GYcjnCWFnnNmYnpjlTzCOaKpPh
N9BB6BUAsYgBPDEnfpBxdjBdQDLBEo8z3W8Jxcx9rk3799mYlxjsn8DF+EQd
Sr9RfcWYXdhSTpw1Tus2nSojj/BaE6lG7HL5QtkVdu30ayLHsFSERk9e+OJU
Gkg01Xb5l08cNkrCqjhw6y0zFmE+zq9bmAlvKljBIySc94jMbGMDOsjmzabf
5JOkaDMslvpprRx8gn3lDFJaLXuCOoAxhaJDRzpGcxSeMdaT2nwemaUZLibJ
d27jAkdPqkHpvPr3gXwpytOrYnRcmcgAuWxFVE1whsDEs+bniBiDxAT58udX
FPdVG1fX6FBDhf5Rt/y5eMC/NU4HirD5wTaftrCD+vmpFQzaUz41l76qoqz6
R+cW3AiDQ3kOCvlgYy5G/dsKLhXqP7fJD7vymg3QSZ9djVX+bu0z7Hh42de7
cIaKu0P4PGAXZN9hPZbgmd5I5LGzWqpRXZj8p+J6M/PyxpjRmP6HImkUd70j
r6CHBom0NhzVAcNCgd6ywl8qJ7HCOzKmfVrwzn4djUIJnNSYb7lk0cLcXc61
EkHfbjFdpuObFC1ATKqHyfbNPgTgELrE+CV0YEED9eZQjOSeORaizr9JpFf2
rPDFXdJu99mzY1MmC3fjM0xZ2Ef5EgUoEBvzh9Z8dh+iK2ndwjHSpi6+2NZr
0SAO+7orDvnhF9RahpCPlxkz3/bQCDJxVWpZT5b/hk+6tCK9GUe1TeRYH/HP
aulPlijcj+zVSOv6Fu0FasdXGgrTU/0yYTwlazvz1Wp/W5B7cRMmdCn4hoJL
8rHtuKZNgJZus/2FukeKlE36zGxmTHfrWlaR5bg87P0BUbgpxAn807aCsplx
EUHhqpOIIgxUc47ARXutVgqFiuJvz9qe52BYR96RAzoY5HRtSPLEyR7n3KdX
aevsQo5BsPLG77aYghlKzyhVt1/Ky7qumaRfJUvIO2Gj3joj5iufOEHHVpn0
akpPPuOnsuIQ5dFSY3Oh3r3Xm4y0vHmaHwoo42wRd+CuvLOx5qurmwoa/qNX
XCr3wfsFfTBJ/2DD7SFTeFvXbcjfE8DP7DClGwKlO6bNE7yf5hh0NfjBW72u
jNIF4feLJzGuywmFuk8fnz9pvOg+7kQZ86UWw/6zkYE/xRKUV9+wvJIaAlun
5EOn4izy4Xi44VfsoziFGmd6/e5P8ly+P5kqL9on1+ul5eVn/JxHp77NOdnZ
J8V3toRvSFMo2BYlhzdqLeEoh7TeFKmBYwIOOaNiMptGpIOW6aFm11p8Ur6G
8RkrA3kJTkvfw9Yx+C131SFIv3l5Sp2jOIiGYVbptLaGkodVyk0ilgS4vjyh
tIrHPr5a8kAb70KuL5dr2Sk9ehBUyudaGZusZne+CUIlPgZrBK5lr+FSCgpv
bJasmyMT8DdN1QsyVUgNk+BApu5ptZCvZrQrk9hkOo1S46I4ZHasIGZLMC3z
Xuco21IGAykd1uqY1/jT5g32UZ/Lxbf1GH0pEnLjvAvON9ixkQvHlQXz0xd5
mMV4ahtWIMHVm2XGvAgRH/eCcRCnK1F5hbR+/OZZwBA5emVW+Lc+C9A2jGHT
L5nCqdGWZBcp881MgEP9K071hxM6WpaXJj9ZlXthYgGeJ7l7tecZotDt/ThG
0AjSd8RRdLL7O5C/UhvuaOG1oQnVSIp9+mvrv+fUdU4qk2n/wWXHCWk8WTKU
pCi0y7IIlHFSz0fQUNIdLeyd6pWVqNwDRcQXd56xyeeuigOp2gcbud4kjDL8
3/dtZPWjHbgU2cnDThUYwMvxpl1x8SM6TqjnmOd33if0BKvl5K8p3whV6jdW
DuqXebc7mu88S40QBnAUw8RJRb1u7P3776PnkRyGsezLfr1SvAMXk3HAM+r0
iqTO9f96TeJ2bnp3wnPKzEuzw5BnLQRmy+bQ6eRIw7Z+ix0/UA33bECGcawo
BaR9gKBFDL+kEwfunSSV0obhsoogicqT91sdmsvP8q27QMzE1/nlwPNA+pkb
9pQg++Qj6BI0qE3L/1mKphiUSXP2YWi0B3yeQQ5ThjbEWNu2XTYVNzQ9xFlh
hgUoa2pYB1XTv46pntMNEWkGk9RbEq+tt+u4zdtLPmv6aov1NZ7V8XOAAvfv
4BxytVBZEO+ZfxYcuCDv3A7KfPbjkhoTg9GiGwa6bbuceQkKChq1NL+6mSFO
rKXWIzkB1g2kGgqMSIMMMd9UHjo3eddYiv/37zRFVPMXUDG5Fp3pSFEC5SaR
YCLm7knTl034GJXMUrJqzWz31QfofSTrTaIJp4C+ZF+zamCW/DqOzYzS+D2k
QeH/LX185ZNzfddLDhA37tbrzbbBPUZ1keV4NZMR5SUTyIXNTf7XuaI0byUl
rbaMPwxHbS7U1b7LHFqTeVKI6Rz7Goq5YsBhBExAJP61YQrnw1Chkx/xJ4Ok
9zIVSyhqP0q2EBt63qfj+2bzf5jr/LW/lPn4Uip9eOohDDYTR5W5W0/WAGTA
sKrT3I/wPp2edRVnG+Sf7s3SCS9SXFgiXxkUsv0g6UXY415vtocCGTABhFq3
ajcV5vuxNA0+ymWrJ0kYVpn4mh2I/9A+FD7vK8u1WJdaAGVTVihLetCu+hC8
4+PyGbbh+rW+TKMxkFWqXSfPSv3PMhAnSGFjKuwLFezCo8yuh/W22uutBEFU
1vj2UKCWWk8jsYgNxUIEvKvliUwWGE75IKdqRr2px6j6SFiBxCLbUUsELo/J
uoAtRoQWLhO/Dr9J49sU9MwWM81Z3kgn5dI/Dgm1sXKDzt/yCNOETfFGTLH5
BY8L/BcONJZbFBD2galegxgkbApvDjiyO/h3lP4pb9/WQCTBNsYhlhKVC2yo
NygoGWnD2UhKpF51zd5QTK4DB8UMaHxiXKZXtyX6IPdpWw/q88gCgTudCEPA
knxDxr4GQGgb5MOEoRsGpONOEGyc6n9bPNPBwaKa6o5KJ5fzASBf9RsKWYCg
gDuJzu5O7m8JeRyfeM4Qju3hBY4xwqxx4ezdALrGHZrQw+IHVbIQCU+M8LKm
Fd9UQMKTzuVYIcJJ62+0f62mLKmonAbyDIRjsjQcd/nCQ3ILchJ7wRl1hHoA
4eAazdTGZ9zFhlABUi7HLDndVBI/SvsxcC07Th2kvVPGigK63E5Q0NZ7/fYF
KpJccH+Rpjywn35ChPBa5zzN0mLyRCdCrE+pgz2B8NhGF6Mf5Y7YL312CL0G
kDWacpckXG588Cg81kN3AJUEmtXSveAgUSjS5ktGWcMBEQBUM01wIxuojPZb
jvXFZ0yoxUNqlK84d/ozusqP4yobiDp1jYYCYhjiKPeLN76NDuCsT3NHmWxc
TT8/eqBeYwsrNwIDA1OD4ZTgXlzX7MkGbTGD7y68OHXcdfH0JUyndh/IgHec
QHAJjPeBUuym4tO5MhRcbfXJWK2BCI+O+/Y5aYa/LWPahj0D9q1i/zY6vL2/
h7xkQeJJNT9rLm6AJF/+0PhevBr4d4i5ZMztmljuCJmtnvUJ7MwC8joHcnk0
yt7CW/Dn0UxSbCshhxCXPqi+23g0lNPSQw2pAxAeH9QhJMkkZUq3b83AYbFY
GfwFTqdYrtvZTvivmrxpadqwSlF2X8POzxwX/gBKD7wgO4DSRHWTGeWBvJ2m
ykdZCdHZIQQSHL2zdWagTEAO88tZQV/xM+tjpsYPha+P7eEJI677dD09CFcz
cUzzkhKN4coEHvAD/S0vLeN+tyxMmRY6nrEPJD0gks621UiJX6VSEIdDLyUZ
rK2dPAhN9iTraYKNijXydvIhglt6GcRZxvJMB19x80zqhppg0lihZXs4C2KI
boDPY7Zu+LJlU6q73xXisngA6hQng442pJrvGNGFD8H4tr98BNKiFCmg34Fz
YsPm8/ZnEIEnscdgWNVhLKX8Ogfu6eAR0dmuV0bfBC+v3Ak8Grss6uudrb49
N9my9iTplFwRFATaDhbQOvuIekModx6DKyQT8FGRsPJqqX17h2DiQVrnmeFq
65fYzTRjYq3cZ3CfIrmislZ8Xxu2wbDqVFrlaMqCZXocCwoNYq2Go0eFvPUT
YrLj/qxj4fUlGbhUeAeZrR1LPzZyi7HyJ7UtD1aSBkCen/9rUfeIrtjtdD3H
CvwqIX3qkRhwLjBxesCIJM9OSt2ZEol1Ql+10IQczvgtgcFhMseQfa0camrb
qxT7p6tKine4GesqXP/3Y4Ce+dDdN5ibLzmMhyHACSlGSZwxj+dDAfO/T3vW
xCqD4pXdvf6tyxFEMKkd91Elqqvmv0E8lcah98HTDzK/lSG7RxztMmw2Il5k
auF0RhGvCX5nOHYguyUYfGu0nRvpH2jC6SBUe+cZ6Ol9O3ZgImE1mtBs04ps
I9SJLaszDtpOqinbMNkP0t3cvYmU2gBgGSI9wGnRKnduhqLR9iD/nWN+bpI2
RPQIav5ZZkEvuHlRw9G+tSKSUHxUwVYZZtiMglxu6u4WbWF9HkcKXU6ttnSn
FwrsDlca2BHqdjMwvyJ/W26yu9YHmiv9D7J5uLdVQmlxB56V7qeBGxLeusXL
rEf6d9l4OpA+2kbTIDQbeIZf2AOWpxennhsBotNbwaercns/mpmKVBYqTl3Z
BCxPETarGi0iqIZ232AyVdjv8lNgplrjS1p/cb38NjdFhAR7XuV5ahXTElIZ
UbAf7wnBi3EUz+HuRvl2gM07/Nlzu3qpOOb2OP51nPvmwJueJDJN0mkmhTnp
8eaWHYC0WZO3EqjFrp7m7knTDd7Cb3NSjv1wWrBwC/Oa7f0xtWL/MSyiUkeV
Lr+yLDuw+99KWVmgi0tfXBJ9NXe8Lrmbyzou6ICbIg5DpdfFJ6bc6jUr03k9
8elIp0ZDEblHObozOSTN0eYL31LJVEGVYCpgWjJ21oRXLzqcBx5fAQrJaD74
TUxP+h2exR1NM4QuXcXUGHVq3f8k0eGZeZhX2scHNUDGauNoR7dbYpul+Kxk
lx5F+tjLMigGsarUZvVwOvpIspa84WnmLkgpP30GgQCLW1CQwycbcjLrkmrM
Eex8YP/kh6VbFHNe2oDK5EJm+Yz1rfE2DVLgu5GYqkUL42geQ+9OSoaohV3X
uxZbBPhdorfwLEB5U2sAajiKR+qbhbSuNzGN4eILbCOSBZ6fLFEKQWFLUvi3
HXwMaXpU4wyWWuy0eFsvd4ym8kzv8/4z9wxoEbDNTnp5Ksxnvv1tgWm57yP5
0I1nfXxEUjdGs18KS3JfMlXqk6xxPGQi6S9WYiL+5tnbrYreCrqWm+b4CYuf
ZJo74czNqpUIeIhClzqaeAo39SK/Dac+UxgFN37byj91vCzj9ek8FBRQXG/N
XGx5XjGuXHRaQK6a8yz8pbdookRE0Tl3+DkG+qcqOxNbIZxKtl8fQAb7HMaI
Fa0p1GVPIsXWPCkl+tHlPRUlvqQFbmKIfmSRCp4eZ5Waaj8T2fCvwe22NV9c
NfIJE56CFfwWCG0FSqCd7wsZwrgKEO0OtekneBm/legPx+gY1A8Iv7I5nuV/
0w+G/8SHCo7bezejWGA1EgUC4o2WUs1Xi9ZvafjsfpL+xAyhGoeoWfgWZeNx
+0oOd/bvlnwAHdK7v6qe0IKqn1NODUoGlk9xsD3xdg8zrLbkdyTzIhzWlTDE
cRUOozZ7pkH4vTdtMscCar7F5V36gnW5WHXLthH2c5SeTSrHgVqevpB+OKTj
HMmjMEZvtbcMeUKvcmZQqXiEYy7O1UjpIwONt3eddcW976ZORW8UU8/oQB0C
PyATl8LV46Kx/Ot0GxEv47N4Zf4Aak5GCES+Yrjaj7zAtqoimyBmRFzHQOY4
ggGLmN5Cdov4fPOYPFEmxPgR7x3HnrQB+sGx1sIlwlkFyxjV5wf4tFhTK3gt
19647wZvWfXDgw9qksewZSrl/0nbyfTIUZ+dWooU7oOY8uqREIxoG6aEyE3J
SrgoR/NwGNe3Ge66r3KHohBLIT5UFaMnLtxEnGdQ4oKudxN70YuWgTbcvBl/
k+Ulz/grsUxgia7/VIDOZuMhhoo+ztD7Vur+b2wXoXRgIrqOrVQDGpGH5jqk
2wr2KQhzgWWXpzo/G9fXJXFSCNOpH9aQ1T+KN3X6gDxXv4UbpHaDVgs0svks
PsF0Jhf7JsQoo2g52pYumlUHGUT/OoLLJNLVfb1MikFzHl44RUxkTeF2z57n
ohUR8utUVPJPYCUnsBU+EvJSWWiIqxiwWDQ08H/tbB7oE9OkrnjBvdgOH1aW
cOvUNtreJQCdZ4OvwJNUeU/e64hWKjT6unAOl/wVl+Z9OjfQSrufjF28JpEz
P8MpgEOm+K4ZETxBZmHs+gQpvBA/u+U5wCdsDy+bkw5p5chCDLeG/CHmtwOP
DhF6mFZuk6TeEQs7VMpwTcO26CKsd2h87JiPfelaiHlxI6M7DdafcUh33ec3
0gMuxyly5TyRc+S2cw25WJb9HYoA4y+j3z2Kh6pKU3b9Yd1sqi0wR1JdlRZZ
uZ7T8vTzz4FmePcPHlihhSeAdm2tydGmu5LEQ+NOKHzGIfPi0YklWN5up1zN
L1QOvNTEVLrR8/Djhlr4s8/rSHtKzYDclmIOUE3v8z5u0wy4wM0XrlOccJ5B
qfFvXGrsytgNopHYOA+mDzJdhVbFWxCwTU8VgKnyqV8i7GaI4xsRZGSRt2uH
bj5SxrJy7Tglb0Awvhoc7QRrXgD9k11YDM/I+wR9pXObhkRepYgkO5RovS2J
lNFLNs+qtzgMnqQyoaT8Fc1EFbsXucZ278H7bIYREszHDqaS+LNFfHYSmaff
NDydwAJcFC4DSboILttDda0SBMx3MuIzVvGWIfvge50kY6DZY6o6/uEDmpLT
u4gTgTD+1eubDBfPSTsdILeWUGsDtYaMuf7wTiq0BGp5E1cnLCVDzMVPF0Kf
EyvQozwFmlJ9bZphImL+ZiK0vLKOsMpzxpGQHEMDYmxnJdstoUBaB22iiHsW
sC/3KzaFQhulTgNt+19olxaVzA+aXtJAzhbfKHd2MpfLfqGyiZO//z+lcfj2
vBlxyQ5mOlY0UgTzKaKuv2kcWCagHrbyRAZIwJB9k3qKeC4RLXTGI5CrlTG+
WSqlXcH4Z3FH2u55yC/bWg29JlEjcEi7rfJ8Lx2pkU77tBWLqlNlPd0MXDew
xdI0zJSBNC1NcYyzpKCFAVY6Vt4MBHEn8cXHh+lzgsuW2j9TkQAO3KASansW
zixsh7xDAh2P7L02BZifuDb/9Ip2Eotfbja9C4YKF8QwCOREUT9DY2OPRikm
xVV/dhhGAO3ngFbsKRdqakJztm/KLPIAHOc6OOiauEk6SV3CLjOGqZ/Wyii1
2gd45Ik61bSFH1pet2XavIhf9vAPICB3e/LvtODyeajPTy331mRMcPqK/HC/
DxbfhMvS7RVzKlldgqvMg9M1WgI54qa0cKdpkyYx1TiXSTBAET9YxTpiu6qF
EZKHtXeKrcou7h/bhaqxEraM1848x9RDlw3xE+jJgTcg/h2lh/4/1b8WKe3p
qIeBzHaWOItcZPrxZvtXaOmO+gO3b7MY9qTDOeLAdnQwJdpFy6koF21+8+Gy
HBprHWPi6rZF2YTbb3P3tnQLFHzp1jtFjVIo+p5xsZJTU+SdYKqhsqZNuyYU
O7r6t38dCu7G2HxTefTNXcd6k7ngw55JCzYgmagbvu1gdkm0O/fGdY/glLcq
y7035h39PmkQP1AMNmtBsO/TerNL7tS6/CpB+NNjNEza1+BPlZJm6B7hnQ0B
yOFY9ShcY4R+feff97LTP1XG8t082fOl1OnobfMsaX9aJb6jDE8u2z9Rl6Zr
7/XMiRlI0FHjxek61V2FNc+3GW1BBfgnAcI7npB0UX7WrwyjmlS3aKHvbfKM
kqZPnHdMRNaFfJy5BqoSiJpQcDQy9WwighoFFFPXXuOarcw45PmliSDNwmLk
x21R7WtUz1pM9qYKmSI5IPr05nHQtOZYw9kQXSlIwjE2Bvhn+9vaZlseuYDf
QZdsekct7NtW6CSIw3KDERQWrwhuF6THKz4ytZ8D3/fmfb+24K+hG4WpsAe2
MUwEidhnwDun28vt2mBYqR+7Av2OZA6h2gbfiohLIIqejySao/uN9TaPoUAa
9b1OLMgL77WWMWUo9B3dP8bVfqkceqm8Cxr9r+EBCrPWjYnfKJwd0JV+3SOI
45a13ypJeQGdE5WFiwVVdhtE0pzk2Vr2EJVU61q3lGTzx+syuzj7LdNDOpR/
7iYTMAWLEvrYchj3rTlEImKqN2sBbRxSH9DMAmBjvYlhCsG8cnLGZFLRFjAF
Bgwa99HKyWats5y/p0OAi3vdEyREZ8MQ38AJZVbvli/2x5o4Ztc9zYePvoOO
IJ79PSY3i+iHi4/ig7hQHmSOnMHUuACoyclT/72GTD5AkOMRbBT3cSGJXVJ1
OQRwpa+PDiSIAS1ZAtZcI+qL5b3pggSGRAWLU84h/5OnWc0lzYcajq9sm/ah
qkFnyVArpAKahjwrT7Fr9HML0rmXmtsAjt8VKxYinfM3xp4NOugSXTUV5P+r
C0aAjRh5N/iAy1SeaWA9qud5rZ0E7y8kn5hc1faecARzDK4KMCvRB/q2rFoK
lmcS8IGssLfiYQkUIP15HYugPg7DpiS/hTdF5ypJGLbIs/jXqgsS+yRapRux
fbLt+q4nFjDd2ipfgg1/0YadSXJKNMRMWn3OmbI820mgOCEp0NlpUNTWcxSi
o4hs245l01npW+wsrJvwJTWmpZo1vzDcfHmopuiaqY2RDaam8lFRBu7YkN1b
kvb9AelG/u46SPTakxqEsGMfzGfprAYM7SH5Ni9LKoqvMlLAmA/mnko4l2qk
F1XtJDHpV0uQ0mAcZlPEBRKGUalTD60X4pg3OPURXQOR3nCEeEZlfsnov542
1OIFtPpCoebzpq8g21RFQMWacYtSSsA4Y2EinVu9Cv7fv+UimhbcTzcXFW+8
dH2TL71e6X5vTA4/u0uIc24/0Ky1mW8NP0llEZzKoK8hhOS0A/bT9DUp5qzT
pwcujhlFLKItXnYyK1O+y6h8Dz0l28TqYNdk66t7udbnWJHQGG1KW2iTS0iP
ffOnpVo+xOHUf3XmlcUJBwpJgcdQN3rmsbvP67p7W8heLxJgRgx33T+znl5I
hOYygomciepXifCde/iog607QovJTWrEeNdEGmXbp0QLy3H70jF/OPYuI5Dv
Rd3sDI9l5+ez/m1vlDASMCjz2b7F03Sqdpx0Oqy2HLlZPI54Fy7Tb1EhTBLZ
ktShLORjKEd1X20vOPGLNUWJ3PQOfHU/sFRU73VgJ6Z2vXrVHEE8f7t6K3no
wbZnm2xSCrZMCC19QZDef86ZDp3hjULQTrhyos2pgBnC46SBfLnukb1WjPu0
AdCuQMWdSAcuCF1wgJdUEE5L8080h/OuTcaEqy2hrZLWb9J0vp8TJ4LbVq6X
vFULr17QK6qDD1jSCBmQTqz+oE6vh6h4c7XKKMw2Pf0kKrN+T0fZ+ZnhQaRP
8Dh5S8xsH2/b3H/sApHY444BrzPmTtmovb3IxZjyshzBa8sYIYauYZFppDnC
fNprdO3MO6ujFzyvPCVjfIF7DmKxF4UISC3FNBZJZIR9C7XWPOFYMJ2SC0wh
YtDnVyzwa6eyZhJHEX00nEjq9afgIG5D2VXNhwAUkKxsI3P7ngxoEsr+m4Rg
o6WpPLm1bd1Nr+giatrJGkXRI8y4cHSPioIL48HF9Xr1Ov3KJVVnqLyaIxrx
0oaNX95y/gV6hiKeVgQL/CaDwJtG4a21lXa6TY/lS9vjAw8gy4PpFz6hKzHf
kATCexeimQuFKBaVUi3FlazZ5Y80yrhjpyrqWEJv/H53Vo0sWavWNJ9qhbkU
NGcaXRJ/3KQ1BPLUYWZyM0VkioT010RWU1b1Ox0ongSvaV4Hlrq1PULESGE6
CgE+mG1VX7vdwmu4+4PHVuVoNBftCzKsnhkS2SK/zPlnHVyhb7HwXNr7ZN9/
GFqjI0e9SZT7mrLSL5vi2JY3qEyuJe8S2424NXfmAQnB3C/b6aW7DlEX7GXX
kB0ZbRb4yHZSLbUls8hyiJRg0G8iSqaG7cbQW6p9NUanSUyMjJDvKYkmdYEH
/2FFZkCfXGtolHbNO9B2UNAmsTog9pkoryXIexHkXCcHMFgCxEa+46N+X/3Y
Ui/5T5dEqEFd4XgkwluyICLEK8j2S6b2dPw49xKobTRFrAgSITAWX07ojnhH
CoF7nbk+vKOOwMxsOrBks9mdcv6P5bELVt9u1hiTSG+rCkebuBGprk9NLcYy
EbYYa1N8gJUch3w54yheS9cipYtumuxzxsMnjjguvLnAv1Ax1FxHjxBn9L2D
4nKhc4+R0z9XL3gV3SC99Eg0voRN2X4NClQzdUAccEL8TUdgJ5moTJ3rTP3w
hSNqLZz/h0EGHVpqABjkzRMyoDHDE42ioS3aS4HEmVoKiUELO9USaIr+BD8X
R/XordLaLIZpRt7xZTmNKPgMel2dyQw229A1mTcHXNOi6kFSGBa9V6oyckgf
L3TEfzupPQmjnWFBNNB7+a0aVZiERFRZXBb/QJls/A4zQYRYN5lXRH6D9iG8
F/89X34yWDeIY5QCgkOvr8wat0T7nTuxMfTpHigTDvoaCmnpEp6Z5UeJEdnU
b04wz6sUF/wqswiDQvaTMI5s3nbQ4oliU1nH1bMIA418EuDk7HWFEMlUWIAb
dUHcC4RG+fNsMfqImMXJdpWzhF3KSsOAXm3zxxtRju/50AhrkjOm5DdzMaa5
SO+dv+iAAX9NMZzu18MfBpvA+APVW/g0FKx2YCMVLTQEkTnptZlgZN4eiolN
2HQZjEFjDv/Ch9rGJAOedtjQeJNufUtQTTu/Ia88b8svnQ2Zbs37PVcbwY5i
0vt4loLmszwJQ6w6GffTfxemf9pDnqP3P/GU3zs0Vj9lIXrRtOPwF2q1wppz
yNn3y48Je9MWNCqAe+fO2728to4APx1ofelaLfF+aDTBzsNPRupila/KmMV0
Jo4YllhTzi4RxAqPM6ZFzILxekFktBabOvMG9UEo12LtG3og7pDLnDvCqwP5
wfT7uvRnx86qjpW2w1CIQ1UMh0agqIelnJ1bnLnhk+nQLtoeHm/1Yo5q2Hk7
REz6Qalhir0F03h9UjR3k0QaovzQOsblbLiNBb4Sh02d7OA5I1VuVasw8fKo
AjYocItffE2ciIizcm2G5PTtEy0QdT1W1XWYeqAaxF2k/xNpXQ8pUzLziSEY
2aC2EDIen55w3IyRAKIsOCEsscSJz87TC++7+CapDmnUciSCxcLYo5hck1V3
x7nwGtbm7xda2U7eg5X1TNgr5QwpUAYn+QFdSZrFRo3jsU78kZ0xe7SEaLAd
H7jU1RFJ5qPfsqHkm1/sNoft71hfXE20mQpNJp6lNbf9MvMVzyPwhmdLWkaN
SznIccixfFMCl62NZbdIaTKcgD8kNyKkgGb7rmYCWv8e0xBaGCqVoxvbIO8C
x66N6GrcfgnC+iLYyAN36UEPvbdPH1/ZqpSAzt2d89YY9SMBUZx4+ZhsrR+Y
1r/YkAMff3irjVrO22+gHRCwvofU/v5kSSj8rSvBDprwOkc76RaJNYTY4FRg
PYDUvtmgekJJc7Oaa/5DOZ37gtYOtkFLnLiIp/mqkCgS5GFfJK1gYJv+P7AU
1DsLhAyJZSCzt0E+ENljnk764c9IWcJ6NuuYwUQ80ScmKvQVcHEYf23pXW/V
g4eq3t0rf52i7Zt7iwFufTXye04HxXE2Bkd4IkVYLQSA1HleD9uuPJXNcB+7
DqvKWKreZjK+d5DjZW10cfv6M5nzBTYkK+vWnLpTup4h9mKBwHVIiKD3Nhx2
JpE8pfqMbNRuIPjru/2yMVoAyLCw3KNB9ncEwhvi1Z1PF6sMD2R0rPnKgdY2
TsVdyMGz5UITpL0CJOr46R1WxpKiCgsARmG08nzeZWgksobkMKG3biQoOREj
xhTTnqRkbmAXPai0NxsVhoQtSjFLwn/krsN6LDE5eTq9AuKBAJMNmOkRbZu2
nNUExrNhZ9sxhCisL9E3a8RAoIewVoyCG9GY8ZWXf7R0pHfQ3SXrwnGQERFG
FMSJ93dpN1rpaqPoOmGgXco4m/mAMUBclARsrHIB2lPdax69LJe0kERQA/IZ
Mj/ChURdNbYL0Wnvxb2JoK+bBcx7Lz9/7Ovkxuy6WN2R3JYi3yxldkoRVqKF
+FgUxCfIOQ4JkoRNb4goKLBIVxw8HVc8tcNSshgvjj/kSCNFUtleHmIMizek
EojO/8ETecYHPdPxkRvhByqkqsRUpVHWUDU15cJJcPbtV/h6ytK6XTeuhFhH
j2ljLHaCEtPPagAdtSwdZgk4m/Ph0ae5xBW22iGFY1facdDXrGrwnO5I8b0J
+i87OCJrVftTQeCnLlE2nIa6aOY4tcFCoP+6pSTj/g2ZgHLcgj2bvZeZyOxT
J/Bt1qd43OVX3V8WxXP9hWQJuJT4W7lGdwQJCBx78VdcvGHvtLEdLa+N/17h
jRi/eDw35zd0VttBCuw4wq02R2It/U1cIrPC68zfX3SeJDuxHg5kDFcQRf7I
sUYh8N853zuSM4RmjrVZHhVUmd1y9QSfiohvK2LLg3ZtoBkBy9LUjYyZIv3Y
hQMOGb68RnCugmeViXyEuvF4dD0glU2tEj8qVnLEI6ElTwHefAJ/SQ9g2KkY
jrfpePlNedZQd0D+cHYThr1oa9E3h2TJ4N2WWNw/ReZeRK1IqnZAMxXzo03/
ONYy5cUjdEX8bAmDpYdo5gmsFkn0tZJnHk4adiTO6BS1BPLToK3uxKufXlRg
Zm6v2nagr92I2650pJXzynsyOvUlRVkXhphtkCQQEQ7NMOQxclwePfBP7kX9
6rn+E/aNZHTFadjK95i31KoSg6+rsxDO57mtQDO7SSRHI1Ch3DrxN7dvSyaT
7CEwfanaHUSD1IU6LQe4HsVuFf0EDdeeSA6s6/EV/JIsNW8k6gXvZHuWILUA
UtCz7oEGmuo1cYH+8IQS1dvHYIzeWbXKHa8pKVLtEGzL+u/kH9rVmfcqoDCk
giGN/Hp4rWm2sC9SMbPPrbGheNkgjY/VxyXPlO/X2AwEpvahGpMpVt6/blpH
1ZUu95lbB5Lhg53r9F6xeOpgE6vJHxQ9+5QXUDHeYG6Niw6AUWKYuOI7xBR9
I9vll1wj/8jpZedX81xk/8g9ug8C7Jh/FiU3bTnNlEKcvkTq1YoH3T8iQ7u9
YAQida9K/BfgsaCINfpLqTQioclrCC4R7oZraL+6kA/0PJwNz7oZpiy5vEgL
Tngti+7mC2F0hZyAcgs3eTHwsu/Hh3+E9SGemn3ZrMVb+zQkYHSAQnFypBPQ
wIrglo2yj9LUyAZq0z4sVXOZolJTJDKW7/N03AwOumDVurS8B42p4P1NrKFd
6sLQxqDedZPjVQTFKQ2+6qnNl7+j+Q8egRXIDgwwRYj1nRenEnbJMFC6FfF2
ucqnzNhMHGZXbdhb6/Idp9a0Kfbxav7IO/At/7uoz467MYhgDL6tA5BXbclq
JhM5BU+ySItM58flsLsStCp82mSoVH57WZIMgv9HoQn+PNSNApbl+E2sPCfc
P+hQ0ft9UxgVJ2g4STB1pwp9CGDGWi/XmkCh2CROttCDIuYdQMig2DBZ8W1b
zQJGGG5oxSiCOvkg8AGg9Ce39X7fLbBr8mk2n6JkyRpmfZSMIic44nIW8/6R
IqrNwmEADBAfmutp27qnE5Nk761wfndJUMsirUxFtYThY4LjZcv2QisbZ2cC
NO/5/Iqf7e3NhLE4JlE7isjzzKNz+dS0U+UdSsNT1971zW2xUCWVnASAgDFl
Z4+6NMfp954Qn8wM22n9FlPJudbgxdX1RQzfWBkCqG4QUz4mnH1j9GI7O4B4
W1OY+N2XR2uYXZ9yVGLGJwAuJ/myLia/3xzeMQ2UxiRshaBjcSMTzZ7zPqSl
6slKWuyBx5Jk0unfsvJj6GSmBAKhHLh18NP0jblQIRPaeDHTg2nqXlu0NIQH
Fn3+tJ0zLVAUn6Lufc1G4wdM64NjP6VK4NXOAOsn8d54tAjqnkJRXdkLBRc/
Dt5re3xn5YoK+6rcvAlFzv9zxAfG5hL2J+p/D+VW0b3MYbXhdP72qDHNZtYL
Uvc07kui+Nnck4YZgM8MRZvgJDp6cyGFrkgdnRdMPeTNR01mNrAYjq0eSRVr
qj8cCI2v5Dk9Cma63ZvXfDBd6PZYTYFbjIAA3GfoTxtBat54O2m7hjvYtVPu
1KQ6dkhnLCcBs12mZgHUXYdvYbUH5vVr5ikt8QoP50QQEUxiIucK7SOv+8l+
vueAlaC7a5KI0/CmFEcYDw+6vImJusDSjfZ9ytGbA5oX6aFwbUnN+DbPAu6R
no5MoAGya0+w7G118uGxOT+aWMP2XmJlTc94bhiAdg8ld+22k7b5x3aFyZyf
mi9BWJq7zc7kp4KXJ6u4r/Ic9W3k/I5LwJxZG/C/B/rxI1go6hWl79KHc2La
q0/uKL25yQyP/7EnbPOoAHrwJJE+mx0qVILNvR/ADY+2PWuSoS8ekIczcT2B
Ql74nFkywHaM99xQ1vgH3xfYOKVtUxhLroNTupOxEqKoqW6tHmTI1H7vgeNz
31ffQ7YJuoGBHZTyijlN1+TLs//aXsVrxZTNXSrb38pGce8Ls78gduW/Zdj2
TJrehGzPTq5zUUTo70qap3nFKd3V2SOkUB0DE/FGgOCqnPwBG0VHZOJ0f1Zn
vDAvdSVOqjFPDAL6UZ/jMx4K3A7gIVZ7bHwf4mw6X2JCo+CT28yGLTpahxff
hk1wA3SS1Qmwl/bUz/R5uND9e8OsQ7xpxjVIhoVKfkO9txV32Dd32jF2cFqc
CyBC/PIX+Ib1rmT9kez+UjtmYXE7CtrtGYJ0KAL2mCQrj2jcM+aWh3wcJd7b
cxKTvBHlUx9k94Z1G8a0c4dbwAt+pbv7HhMf/SHmpWlfk0ORMYUmn2gqNdCB
hfn0TqxfN2gW+viMnzq7FPUeFUDd2BPebifnsigLLCYEcpvjjfOaT/ii4h9U
jJ/m7GgNm6uO4WMKExYQh2gQWAVWr02PiDr4DJiqC6iDSkuLcxWXpiNO+QW3
CAgp1U07UAJOZs4DSPlUqfgF0JK0DH4XAJv+Cfuq+sF3WT6vwUFI7nuqVaE3
YvD3SoCm+7B3ni9zWKSsyLXIcfet6DZnzPGRmTwb3QhY1Ie6rMAMP7zeU+ug
1UqPjC6jhvoa9TLpXTT6tGBlkoR/mzLUbWFYD2gMiAMsp+V/QSF3WnGmxk8l
z0RgwIuK1KzlFI2DZ2HnJX+FiWr0oDlCULankWMA2k7/zbPP3P2ES9dhPIKm
ApbOUE7D+bwcBiqx+5CGbcwH1bKglOV4hxGNDQCrZQNYeUWa0tQ9qdLVEXl9
76zghB1OJkY7AuxprDy38FTtEhHraoZgEUaDr1p5uto1EVdG25AG/Om8cTAP
O7I5XvSaVH+aGM931R+9So8oK8oZFCPebqVF7B4kzN4PzsnDs9CKEbDWko9S
RjCSubiuf1E0YSIJTUuTwvwwJgmR2FS+9KCVHU1tNQMdr+1XowBuY2Hu+z9R
pTbF3UMvF5czkRIf8QckoFLgJu7ieXSckCUeZzhA74hlxyzebW7ljAlvzE05
WrUt8+D8QyTe1ah+MvCQKR8gR4GwMSwQpZfNFzWoAoMjJ8i2LkGvdL3gZqRN
k3mPS6XdbmM/xt7eeJrC5bIPaI4V/k82DGgOO3D0+QLAwMQGJxZCGZ1CkA/V
wM/0UEGCClqIyJTqkboERqJNIjnmO8HyJeYxrtD2MISItZlf+lwOLVwAs6wm
wnW+i+g3CAVtadgRtUz1i5LGg5z4lC08b57NXuN2earFKVcrc1b+dsBmrIr9
b5HO+eHk5Soouw+75bb5msJpfgDY3Q85PFoQe5WYLghnSEDKBBIqABo6rXpC
0l1M4YFKDU1ZFgAZ/+dtBL838o9R69FXU2DwH5LcrwnyI6hap2/9D5WhdmlX
2FpS7fKxGGfUMjAX145P3RhElfP4BblE0ED++3QQNAS9g+hKv5eEGoznkZx5
v8Eoe4ZVyxVuQSHgIs+Y6oZnJeG5XGx91q0DpMiRFpsrJvzmN579zHVmoOQ5
WEhFZLtf+X9SF+kfdxifLm/Gj2oSEcD3K6iaRcvxOjESIhFd5kj95iA8740N
eAlQGeJAMHhB/AhjwwzX3hy1U+jGRQPCntP2EqDhdlcALykFdjkxYvopl2yC
ODZkEf1MemuwntO5CfNXuHRwaBAQtEnOebWRTtuHRF271HPlM73ReGvhq4JP
4G670aopYltlaNrzBeAWRR1UK0Lv5xjmXlX2a6CX7UfpWJ+CzqwpgiuGsVq1
iwR8wGR/vr8sB8NrPi7Slj0semwWeSqhbfgq8Ma5YFSq8vvH2wkNTgflCa+B
K8XbrfaJKjteA0Wddmo7shBh6Krmb8AMqsp2iqNWhkm+4009R0R7sFGxM8X6
B4pLixhZmcDRC5Vg9DHCd7rOkMvu66OqBybrAjMG9s7Pk1/jwB9fjx5WcZ1W
V3jaIYarfRdmxDTflkweG81OZv5PR0J08+5J5inwXyL2a5PYyEmgrnPtQfeI
iFd4CMDPbeAckgpZscdF48TZBVTpOIdKKxDaOfGgQnU9glGs24GA4BKgJ0bW
0n2bi1iP2+dpqlds6X1IZGytto+zRYce72i/wg73kNGtwJAQe2eaVlsrt1wV
8OIuCmBIYZm0+ZpQmcPAfEq4P0G9EgERvx2Y3hfiYjmyQ96O+AeqRWSUYu5F
edGijIuG2KHFimNLzMUHQ0tx2Ulh0ceXknRgmtd0hq8U23A5nDLWRM+tOAhm
oNbZq8opUzhSwfyAgwBu+jH7shPg+VDBTuTykyzXB0+IcSr9KIrp/TrlSVLY
tscbeAAq0BztBG7dM26cUE6XAexP0PWFwXCGpxKPhQ/9TRyiELYv80iW6zrO
9QyEEw/YaVEvNv7fUwMfFEXlcEGWHXh/GESzt0bqqJHLEakZGiph66LFN5Wg
b1sYb/Ve8zOya1C7ws0//oObW+n7r8lRxubU5JBH0Jx+t0ycX3o6kqIvjOH8
Az7aornNghD1vRwH5SEKs/YpvlxUpLsIwcULBgCjkx+ALG3u+pM0CQLlhrYG
UWJbpJ2/CTTeQdwxJrEa9QhiPntJYFYaM8JbfC60/FARuzu/lJ9/W91v4cjI
RJ3lA13M76YiFeIJV8CK/CZPGuxAOeiE8d0/J8wn9cgUmij3jP2OxHoEy6ls
7cDcd3jZCcKB/9bX18tTJ2zpT/bSbOUI+iUJjuRxvQQKDLmARo1o6FL7SB94
afzEsbK7DnuoeTNpUMBHoiHO19dD6zjVzUXXZiPx/wVS8+uc0Z0Cw0imxdDb
i2tv42+JMtPiWKasjSvKrVfF+N9YK3l6G1+UPm1OsVn0TWhw7+lBDQA1YOeT
DC+d4K7sM0HyojfDWfaDP3S6KeorzqAGPuw6vQIla9GiP/xIoBU2/fyJYARz
fMCgI0DuQYfLTD/qkM4FimHjz6jZe8qkqx0nMQMsZn5SMt5jzVTWZ9cFr5Fe
hCDOsl8laSV0gQUCnj7YLP/ZqnpNbROuqnULWzuFRTLxBe1hE8jAbl12xgbc
3MWoROcDR+JP3hBhh4X2C6SUO4v9qGs2by0Yk39/JZ8wzmnQKt3LD0r4FkvN
njQ4RqoCehteejj8friZfSc6jz+1tV8NFec3uCPBdb8gTxSV2M8jhYQnuQVs
Td2RxpIfPLslv7tOkh5OP4XSjI7xUdAZ+DxULtTnpDconRt2wGaozb1RBRvJ
YJQJolNL30w+1NKUINX7CuSzCduNVZbScGQsgQd0bZEvo3n4/r8Q7t0y87Wm
EF+uTvJaQGPBNverARgBeZdwMqeOVZ5RNy8RIr2qY1XOcIGkruKBdpeGFFEn
7RpD21wvq0COWOhLywA8zuWWB6++UlTVCcR488eplnoKNSTWjvlq6butTf9V
mIAREk2mw7JLgylEuZfs1YQHyWjPYj+4/sJFacmEk7JXQTH3Kjv61LkNo5TL
9+0i/ZZaC4Air7K8N8JjIwBch5h0bz6lvWRTVAJSuJkQJIo03X9yVW/0+O+b
MRicyw8HB2DreBKeid1T9xnkTsfp9qoNnDLxOWOE9/J3eg5N2ALS6/YYyt3M
YmfZ+/nCAewipfOPEPUHEAXz9Itp8TanwDqprs3xQE4g/fnX/cyHNN3wLu4G
9/uPOuY/rKlKosH+lDqJKjM7MtGkrCeqnkd4Wh9iZBOz/wBcLNiznf/dS4Y8
+1GG8RyV9OtExvRAVHG4O904spvMYXEQqM02TLajgxy8kFEuIRnL+8pD5DeK
mjGeh7v3lkoPSuyOSPVXwhNqGfZmhsDM7Wa2GAhFSOoIVQfSKy33zWuLbOQ3
tiSoUiPkWBp0UTv5BJrB3izwWxyFVnppQxo6+1MxuBGnNKBQO1eGPJ95ctAn
nqI7k8QgHcNusqQfPF/xHZRv0MQJ76kX3AukzHRpMpnraXzxE8qI42CYk9u9
MpXIuvQQXBbyTA9sq06LVn+VprWU0G2yOJTlFnhpep4imoeUB1J+b9AmMhDm
IZzQa6HOQwycIZokTL8jPcQyyGWOM28Oxjs9qql4huXG+auPwlkTbShmTggQ
8GXu0x1MabAUXuxJbS89ERDSJJjbiidZnvCdAqukoyEVxsBuy/Si1xQk2/Hs
kLbji1lEpsHq+bpERQQMbYFJ1GljixtFimG+fEwabp1JEVWCWJGsLO+4Oh05
4Ei9Ftp//kb2eqfWcpQA53xUbvvSo9SArQLV96lYXw03/LXc/oAJCAiQE0ch
6YybY1ue/BvReQmypbWjZjUSJfAG6HUCLWo57XLZxd3Oev8e0CrFnb41+zUb
vWM85cWW5PPAo3ZyvF91RrD8P+GuBsOUEauHnDUi2dusbm8qOhD7LIlKw95r
BOVdgJQARx6AZpgophIbWVbL/rUiavLtSN8As72kiPv93CoQc82nH0W08l4M
Fo9oVfqMFGNrXGtNw7dpYc+kvzkd3mFuJwFPiryjB/rNGvv2k94FGlrgaas8
SdVDml0WvTM84iC9SYYTDx6zc8nY3yHBZ7QaYuu+7OkNfQwN4LKrVOKJBmLv
1oc+1K9GmPidzsRHddEnkSTFpdkygBFycohOGB2PeWHgs883oHwxVqorJagv
WU5hpkZ7pdTNv5zmt4wthUxWAjdsMYW7e3rxMgZ1SkCE84SlbMr1UI0cQc7s
mHi8/JL7Zk2PL34VXQffb88gXZXPg+m50Krbt7kWxbbBvo2lnbOIZsTs7d/7
D/w9mbHQTmbZp0Cs4ZsQ4mZ8ZnDO9Z6guqBf93Z1aYvMRZIAXpOwc4rQURB9
gmYig1jN/6CgOXif3l6muW/WcHagv8wW4BE4TAGC+gBibj6iM7IOnHClPuAQ
70u4g53tv7do8qQUYuCJ3b9I4hctGr3rkLcOUzjW5VKOwUEsg7/AD3aEH0FW
cvjsb947m28hlcID0xTEXljqwcENC8et+EPNqPHQoTBbJ1iWawMw4iA1kx7k
GNLrul6X0ixpY4nwHY3jpZ2OrdBL0eSm+qfWFQ6BKss5QuRi8pHAuJhG4+Jh
fzfDRUgeTgBJ/agD5wauuu4VBPggJlFleNzBF0WQU2Oilm7kNECusqE4ZGX0
+EvTn9n+vW+BzyvaC4366KuTMnHZZRfo6WtZBteFXhF/tv9CxBjiQQSI/+B/
OCwOcMUBZuclA15ozVh0NkH+SKjh7BkMiTuuFsdkgtclblDVxqTqYLQiZ8xx
kyxAZmwy7QZoYXVZksDYHNKhHkVPcx8xjDoM2h7aUe6t0EbtlyJ0iGGC1pwK
7wJyoTldCVz055/Wm25Ym7bngI9nNaQrSBQusgzbPnnouIHHyU4hfo44A8wx
Io5D6RwlIQFEKG0vNRYCnZA5u3GGUMeAfuo7oe4m6V1vmId0LEerYHMNLuoG
ScIJdX9lZLuPGBc9CqJUm8i553YDdUfgRBw5aHjlA7N5eiaH3e8QEyZ3V3NG
aqzctPRJgOuXeAjpUkS11owoMnFsb8b6UxkxBpp9DcPrq5CB25fAuMlNe/AC
NFIipzbkbUgAG5UdyBjfPUcgtV9T91lWujqqk/Yu2ChecaXrbvz9kxxfzYIm
qrdNxfDwB8ieERZHf368ng7FIR/7Xqs/7DBzvM6aCro6BLOA1e/ZFaH8whme
9KZlQt6g5rLpu+Hu8xEg+TE0pUIrZ4TXXrSIBRic/n1GmSMVTbhctXNVgelg
SyhKDbOmtAw7ABu12L8L7xGBebTrglZwlc+d8iIoyfmfd3gHBV5pLArSgt4I
xDL+FQmcL51eP4FHrg4QQDj9B4IZ/jLKAZpqOn1KZbDm91wX532qV17sROuK
pl3enonObS02AwIFKBF/LBCNRF2ligYf65AlPuoUYZDRxdGCeilOdk2VQJkh
y98SZNKVKR+LWUNlHEQIScpewMziats8uwDue0eN2t9Hiew0RbUsjMJYj2T6
O7r06ygeTYWQ5cCSF7Ld8/na/mho28IKDabgmK9DRxX55sNwiVSdkrhR2z+O
ipcGgN8h8FVzn7xLYfsXlj4ZAxd8LowYZM7jrOnUSKFXJCNxt5nQfaZqcVGz
PM3/Bztv8Hyr0GpeO3EfvWja2JulqRSG6umyzGNfYwk1HXooRiI6CPInjXB4
21arTq6yA+jy/3hfCSyMYBLW0X7PgN1oYNYkIYLrg7ZCu4XAlRjYq1QFYfKX
R7M973Z1eqsCN88L6lJF92J6M287RDFJTWaJ3Rce6IY6pHZ6x6Pat5YaPQp+
y86B5bWlgEr2T5xaAaz9fvWRFujbaNl5AtIwGsSc8DfYipcOl5kJnfeakmeH
drnhFdsdk9q9wf4ME9GCqindQwnayaauKe42qApSCeUmO9dS3IQ1aebbYCVD
rGrLSd2ZNtcUlUBpFYZGTZ80RlVikGe/tNFdy3Jw7Fa2RMtj7scx94B4vrme
sfzN4i0bBwZqqYQ+oHTQ8fOF7DYFfh0lXlrfC1vSu7SF8HK/HlFIgWdjRQn/
RQDR2nZNiCjvPO8+K8VISEMmvLTpqQ7weM7GOj7s5XKSxAM6mu6CwCRQY8Ps
kiRa7DKr/ZiGuDrASKa6LC9oksuoFEq1jj7yp6qNUj1q8v18Oimlr8pIVWVB
kuJMT8hY32ahcfPC/FFeeYjN3vsOvcttwj2eYxtUwXo3wV/3sBF6MyN5AqdX
OCv2UjVt0n9FQZ0FmjFAXMceGnmJV8ALpd9lB06hdcyP5FyJaPyqB8iLidbo
Dc7ce9JMG6JdCTYc15JwRbAIqjtb2jzdWypY8QXn+KGKCY8HXdHsMDXpgRGm
yTphwAXH442OX6DuPHyZscHdJRUzwKdJz9wXbMLSrDLuwqUAxiL6sBl6Hz6b
hcWoNGWMaGjfl/mpZYfNuNxFLHffapXFui0UqMDYEyiE4ByazDM4Qz2s5a1D
7i23mB8O+0YNeL7beZy/qMDyxXCL8hq5teAmFXFtZqbLXJhCkVLU3lNZP/2R
o86mVbyD7eXNSTG2IOF2cV+gvwJwfZQlTAaIIIS7giNUXnFI1cVZwJ9fin1x
M1RivB4/scxGQn7fsHu3jiFCTq8jIlrkEPM8MIIhDnIPPx8KPAPUIWVyXdCF
2MB7PpIsYoaz63+N9FVPwNR7Cp6wJMaKs8+rIhAR59tecpoLs9ooRlB12wT1
KEX6Oj8DRa06LbO+BpoVoPbLrcNvsM8Wn0b6FRmP+zwYV+OkDVjfxz8vsG9g
Xl5yd8GOdOSTUjeved9pJF/NAz++oCEftiFUQ5kUPeGRW0F6zpX/XTV7n2fX
Cai3puRWNYjOKnEMbBlWK7uov6ZEWsowO+LKIsqPL6T48cARC3gBLf5b0J+z
rUJTdsZutwVlCZk8DLAepqLGRxgu8L9/SM+cVlDuEP44fFHyDNIV2FcL667Z
GG8qkrVFpirajO0Is3eJ+aAwT/GLAyAPbJyTVFU+KCkEMRbelHFpVnwpwWd5
ttG6Ute+Q5Pda7i69J5cFuk8ltgLVXbnJSAiygAxt5+41p7WTX7AxYrot6IB
l6kQunJMg439AOfh/0tXt4zuEfHNogkEIEfXSpRphzDOO9OtFbaT3lRwSiov
SeDCyxCWqBy14g55p+vY8xlyXe09AM9MKFgdn1C14coaGrJCczaOPRgs6hA0
B4v5R1LwcTJ7djDW031t2AWmaf7Yd6Z7XPf5na/9vb2OMs6ibTKB4qIJjjnS
AFQYq0LtIDjeXntLSDFDa0pxm1RqfKlKhIP12lyuBSliaXnZNBQPD9SFNEec
/7mJpvyaQBe3zVeifdfLzI4Dq7ZQHmnh1DnKtLGIvnflcRBpkIiBUeh88q9Q
bta5sSyw6M5bnQdpo5tFrEU4ENUB+ByrMZujAWLsZf89YJgwSae1AYweR3T1
eBGmC/CCp1/aLyXmHoNRUsl0hQo9VQK8cjsPzoYyls+W850/YFCVdWzGQmfk
WAxEhlPXOoIwG+7yk/CfGO7qeUjdSSIWJMRJA26RPX943A85PeRuvwdyuNut
4eTUsxRQfpQJmiYv3MiEVt72ChvnJXBn03Zy1ss5+dQp9sLQLc79hrPKVt+b
YVp/4lElCjBvkJTaDBpryt3eXFQt9f96NrYrOhftUY5aHDHgG32xU0Df9I4E
nl8H03wl5HRjm/PSuCpYmyGbjr7f+pprluUXdIhuJtfbS6RKxA6RoNB0N0fK
z1lKgvP5VFfLrpvJavCdAyWKTM2SFGlCQe+NMFObazW78CLow41UcOnkVSQ1
ar5CoE8NZVEOH9ULEpIpgu8yl1CvJpMzTuNzhetJS1PFKDMwDOZ6sy3UKArv
KZG+YYyZurJ6F7zr4QPtd56Wm/JajgkxTpb88vTwqov3ugocKlo18fvKJjCl
gbzFYWyQUpclaBKvRfWapeG+4Z9zUwkVX94+L752UHt71AhSxdNQ3BQJXZya
7zzV7rFuZAY1aHQgrbb3f4a6ot2byj1zpqBFYqiHCcdcLUS3mItKPp0jw7m3
sXTIgA+mlIalDyKCDQhj4S6PEMEbT7mIxGsiJaH7FeXK11DPn1q9bIPX9YZz
8lu4OE8/eyUUdGk8LC5AYh/niQH0biEMPh/VipI2VxUl66+keshxOMToBAUU
WkzH6swkXQ/Ul5k/gJWvzGxdsZq3XjzxQSAo1qbGcGbDTOL+LxSmG34FYsp3
XoVxDGz/2HfYlWCyT7tR6QySsVPgZ9ylj//MnbwjhoRgAEqypYFUQeO//StQ
iEpi7SYhRUQI+9XJbpRtwa/yP78tCF5w5iYkjYs0VhAd6bhuGwioI+6YRJHR
LAVrwSQ15XZhMcMgzZKXAFIEN8Ji9Jo1P00HyiOmlf5A5jHsGd1X8W5OBpiu
loNa7b0SAF6o/VUMajIEZNGhL2NwrxDrlyng3gYa+2+/ieFLdC99I6meIOoL
QGk594xQkeZdpM4z9SCj7rLGxd5u0oFNOw16odKOnNaVuQ8pCW4zcMeNK5w8
pfWUI2jgQxvbFTzCdYoR+BH8PC5CvFyn26ShB53Ky9wI0EcSrQ4K8AHMjSf+
1jw89JHCRRegQTxBF10Qzc4IUXaOSaDJLj1yxnv3vWCV2jurycJLDVwgYait
6/KTf6WQ2UC/ViP2KNzzEZGR3dfVRTKMe6NXUGtVthixr5WVpR8dqf23/C3E
ZpVFnl7icaxJz7PsV0N6YROT1/zVjGbTPGyuYTO1pXPApEFjW37/xu2bY9ai
uHYoWzHSqQRcD7wAKExsUrG3d8XKvSNuB+ik/g7/QANJaWdlCG+kOEbnmsyt
qhTuaItaT02q1T8MItdhGizGJNAjgcKLFAtd9Jft1n0Tbsl+A6kt1ckhmU3r
0CKVyv2RX0trhaaI7ZpNfc31/H/oy4Cr93GO9OHS25JTvTavuh2sFyc7j9P8
zfyOSZqyEUf6BwxKfuWl26tLWZ6kUiREqXZ3RHAlPDdXTxkFFeBqgz6amGSI
YdGeEwmX1ceWwOcaWEjRmT/3tMr5/Lt1sRf+r8hrCDv4YRWOpjvkZj1U7NA8
W6lXQgEhlhyP+17E9boa0E4BACAeVxAtqizU70imSUOQ99ZndcrKgCt+pjd0
Y6LOsFEWAiwqomkbDU50gPrnwiuzbskuWVRpLg65s6WFDTsrwHNtVjtOpDfc
0TaMofOhoqXiYRHmj9cajCjnmx5YtaEyvvsMzuCbt8ItEJuXBT6wix5r1kpo
y3+vvPBdtFqs0c5UFYwOTPcXBMPkYZgry24xJ8NnNuR+/Tf0jN7WIuqgB4EF
nJCRz1J74Xd7R6r0ak/j/InAdO0CEA1Lqv1Fjx3ICMdZiBOI8HfAtemfnqIa
IpRHcjKY9WqUzeEl1rXeqiQMI3BercWbIwRwtFH+eDY9mHBhQZ0DCUSPpRuw
2td3aSn1pNRRehDKkM9GSw/7HIJVYYbQTO7COYThm5E79/MEkBH1cKlZoa72
3qJhgfhPNXYjIfi/5Z8n09edzUdIKgGpBFrc6joJtCIYuet8QRzzGlL+O3Rd
bIjPVsbrGzc2hsUiNCjuDvqA1fmeCbNiv9a6rylTY8pzlcA5m3ePnX0V7P98
9etYTOTu77wenIjl5vnNni+1RNrqQJv3X7sMiY/iGPFwbwLwaB6GwMERftoe
DG40GuOz9IKrONUlm5oqA6oDHtsgJE4yl2VPVWNBeWVx5VQcNBefCHAvsdiy
a4N4sPIHQ2sGelalcCCklyHOkRKOkr35H849Gp8+ScutpDrDpeTzIO3jgh0D
ggw8JDyMNvE3TsX90NRC71FtBoijs1wAE0653UOymLyt5T9kyo2WTyOPrldc
dxUOebkiyU7rAkty/EbhRFIf43NUNFi30nZ2su/quYLb3k2HMZIT068jVpRQ
pDju1RFODD7epgk6YOWvAXTBHXcZOsjF+MgIh9QwOv752gwVGy9yD63ibVov
dPUIk5triymjsOHioHh9Zdf5+cC9sGQM2EHEOaOdTAkQrz8ffKJRFTuoEjpT
XNqMlv3pg2ALJREJ4+OAoi1a5UzE5pBA1a+CNMpC3IbguPF52Xzy3zoxdpPn
tOKZ+heq6qn+p6DsIn9MTRnyO/PwP4YMdCf1+Yj8PXdGMjOT/3nx3dunmsHe
QhkMORJmo5ShH/TdLaCftk5asn4OdHZI8jza7sFaD+G0P8NJAjXAL8R+dciE
P9x5Mp2HNB6Ku1obAAPGrG3LrqQpRwHv7euSS69rR8mL5TO27oQyXLZjOQbX
angTRw9vumxhFg5YIpUAN1dWj4sfoSRlDHDC6RfmZ2knBXTqk4iIiBL8LOjJ
zKvUBg760hfPvV0W7K9OQX5VnI3H6+CjUM0KAZxEX/SPSjjVHYQ6fNW5DjOO
DrN+3UxoQQG4+5AthTYkIdAG1S1UNtWAACKDiG15+VRLBSte71UN+iX0amQX
4wgXCqEqjl+MCf6jXOK+0qqbKAMCNjyNJfemHRHrKhKfBSuGgAfVzETFGPmS
cyO2f4+w+PlqQPepYLsAGD5skOyQIcfs6ov74Gmi+6cHR+IoUX9JjMOMe0wU
r/A6wLtpGUckl72sX5Sv6CQ9C/6XnMCip+97HY2ovMrSrj+r4BY4t0IoY4ON
tekmWjbViEDP2PN0h9vkNS2k5awLDrBlUCesSxMsmGZJH4vDfAN2tiIjRs5U
GcRCC/h8ZH4uG7eSC9xEe+esMi6ZLphZLWhQtxZEtCYPCCE6oA6rA8RonUsT
v4B7bPZ+jxoKu1jD8WsxBd/JszGQLL0V7HSTyzL0VRj8U7bxZ1CuQNA6ohx6
gOvGjx75l6KGzxbHKiIR9C8jej+A/o/lWpqjo7K4HTsJnnf/9MS9yHOrMEqG
oQ+gDIPcQhqne4cP97OycQXs5hz9+7seD0mNTZ0Olhapn6ipQA1rt9LCH325
CU58iauxz95eKnbfZmiSA8AXq+/OFkzUimDDDT+HPYQdZrsrghVhcbb3l69w
y6gVeUH8IGdFdL793qYrO61b82Tl51erRtEXUDcRotmhFXaDv/gcJ2Wr3276
33OQa0YqRWSX/DrNZSFX15VB0Y5DgcdEmerFzGD3cOyvPNt5Zf5bLGpDDHgr
mmczDlYL1aoz0I4ZpfBfMTUYaH056RM1aIb7vUCVcY2V3xEIF6SFL7m5/9en
kYsmEM7nqMUrwwwZUYhDOXgN3BQrus//i0J6Ph0YEmu12/KhlV6eQIJJyuh4
osPpAHwZSooE1UaCRTyuDPdFpuSrVvD+nQ1djNPUIMpoaXF+o45qS/ebfZJ2
X6+i6j2wd4I7yQgt718y8Ob8JXskZjLml07l7ggFbgVhkM7QreCFaq090+SQ
zXiewT6hpz+RAUkyxQVN1+sxg6i8CisLDgTiVJiwFYqeG5dEfmK71h6B3DRo
KnQ45T6cj1XRTy0YUWDXvaxKG49VZb0zg6QD+aWa0RMr9+RHkBjIkAwZckLA
ldxB/5FO++uU70F8sSx6jgzG/gmV535w46xUWglaeiRSNiPccLPD2RAfMJUE
vOKA9utfJmW9o5QvBVy1QxGFHGxKdP02ICS0uc5ry/bdGr2n9jGuP+P0DQeH
C6VOUmVby+iGiAf8//512IPOSq8bwmjCp8V2r8ZkRCzbFIHSDXftLf3RSkzR
VLKR/YBY+puOkXDdYEB893mqNrm01KxVq+zceejqUOoYpwpRdhI8kV/+0JC4
0TbMGgHFBqmiSguOuL/wfccZiXLyM2TpboD0701uEa93TYEqR6vb5t/v9I5R
n1ukxTGcUGCN8TN1f+Puo6vIcu/SWjOsvt2Q/uDjJd9z0+NoZ495v94PsUNl
G/C0V1swkewEeB7uH5LIt7MUkYEKYaeiUT8Qc4nbnU58ELoBpSHCzLLYOUhU
uW7p9I+Um4rho/5fctGObxBo7ibvwNdYQSs3jRKFBZ/XihpQ5q8fKneb5Rzi
oHcXPaf6ieD+YJoouUDjdrnguKh7FSTT9CGGXZveQhUAb4xvUKDhm4Btm24J
rgxcCs3/uWedsD7Gx9WSBAfffwH4MwZeCHrXHrFTbZQLWdYVhZNh3sKFwS9p
pKjalC0Lu68isiYf/NHn044r0Np8aWZc2uRSc7TsFjXuxJDM9BxtXRy9Zm+Q
PdCo6QqR8T6cVMrO7Jha/lJn5nQr8VzEV1lJinmI/hwgPAfKF3472y7nDLb1
x6RMktc6jOhvxUl4KHYXQrXOJNGsLsFssTWtgTvwXH7QBIrzidKK2lDd5Xmi
EocaavwsBUwjJm9f8caqCcfcQJOEbXA/R9o6vHn8ZWgyPwm5GS+/iL6YekvQ
1pUzvt6ZRyNbi2B3Bg1z4j/dNl9uBxNbU7EHIH6X5pe2O2uJmBKmZc/kkc0K
41t2sHtdj6NmijBWk9BPE3d4uuAHrKoUEb4ZV5z6nzrjz6RV39QC0X+mEUX8
N5QPg1+e8UVO//1wF6wFTfR9krFS/+BPAeBPuNfYf+9TDGbAwZG2cwUqJLPm
dBGoY2SRAjECxVH+ifktFEuqm1Uc++pT+JvrQOQJQM87s6bWJAuUQ32shzfd
BSp/zN6QfgKZphm5EJ087ntoMSC+jB2pyihsMXcDm4gcnaM34I+Dd6X8Fb3e
gyuPc8yKtH8TQ6cgD5FVuXWK5hibvIShIfkGAWF/bafIxvXeF0nGX6f4q53b
2++VHIEzu1J7Kqq/wRzp8nyDGFOj4XHJY9S8sCAxD95HpRK8eN5ZskPsvkjg
5iTdHlETqBkY8mKGM/xJhSDZEEpB+ngy9K6cyid2C2qT10oQeiidJQM3rJ33
O1dqhWfWI8TlE7Uc3yqDGmIQBs8az+Ncnc9psxKXdHN6O2z4nulG66ERnpdJ
qsGD8O1JeAlwyaf3i4Wo3X0dWuaIYTdS5scCbxGRfSCJtDsOeMR/xL3mAH9V
ZUq/ykae1boFO7+mGMH0iLM432/q3aJvzBpZ+dsku+ji+0Vf/uCdfojL8khR
jLGH8P8nD0c9Bj3NsPRSss42ncr3S5Fx0U6pVuektIVNEKZhWmjYHjYJsF8Z
lp2Y1nvc/59xbq43n2dQm/WB3wLEQ0BAkkfue7eYTkb/bbj5SRcqv57+Yc2H
6hPVzDAcg5tLC3pms1cwFIWXZXSR6gy2bH/DkLmiZToGql8GMsdX7fsK1l+X
1+jqU3sn7e02rffDSnf5HyZ9c9yf7O0cNBT43qwbt6KgossffUmaEnUcoyqQ
Np5QGlagyCY0cDy7RJvcJO2pzEZs+cqCNChLH9RVYB5eQqv7x4gsZwM2vfAx
f1s1piYYpkbjDBQvBiJcM93jQbe9XKX77bSKtEsRYc6YOjo6JHq10AkTpK9a
mxyldpZu6fV75VgqCzuVyYup+GHgLDGC5Yh4T9mx0tY3ePC1lqvm8F+9gj8j
HtAficAQjJ+lkM4+BXmZMSZX3YAhoYdyKrDpenXg2kn3RGV00F80fqpjB3MM
d3WzagXpcio5SBsL1GDyfRbX0fUBk/CFTqk9qnx4kStejqaIE4yEgnw81yxz
OEUM7fcZ4/iVUvej8uw2adPzmFSXoCPdSeiDa1242TYUPNNEGEuMeGSy8Vtn
mKnrLQXG/DdNgTrLB20oGVNFlYRWZvauZV3RSyypliIY5MbcJ5nOaVCcYIHB
5JTCL6wm8fGMM6H5lH+pJf80lBV8InCQgo/fOmxw0pTQR7zjAd1O8F2/Rznk
RpRqc8vVCKTlocuSN3KLsZdYhpUEvnfUJVA6Bm1/39HQvdZKdrL63dIPkL5y
lcV6jOleYlGcoyJjzVSalDiD3sYcvZ+HC8RgQjmQhAJMP5I4Mwz5YJDkNCJC
WagLsLWf9bLLJby0dHeWrD6xKXbXeKjTGla4ICvdVGxdOug0z23WnQezR4an
U25ob68CI54SrdzM/I/LEGCMIBZ7EylMkUVZG05Bc/1WLUFCY3rFEL109hYU
ILMQ3E5z1wp8lMvLaGOijZDuipA2oEKUDmwDu2SkBV6PTf1jxWS/0JbSDO6q
IGFbRLML5LkHC1Zhu++pffHppjf+4wYoA1IMXD0S7ZQqo6UpIi6e6SQVZqF0
hYz2zsAeLKTmXzMdKXQx/3mqdl2GE7CWs5gRp2e8ohyMJ6Q4oamCYgcTeIUa
Uabnr1+a1JikWRBzQtbsOYXJ93G9KZrx9BPIB9O1yVVNFQgLCBDH3/5u8R7c
N7Jhbc+yXteUvjuse2rvVqfh//MhG7cR9rjYY15JjL8iXf9jXVog1oY6QrpQ
7Hs73nK3VUoivXkq1TFV/GBczS8TeeOpu4Gd0tffSUQrMIEKi0em7MexRylF
Y94ld6TcAYr8Qse9GW3CtQewqBbFFvIiJzAHnDED00PAc0hgsYTioZ9r7Z7z
1VOKjYPLuEb8L4dYLfSFqSJwfe54XdjOfGNViHZVlsVu7OEaDWWtewX34Ak0
QWnRLG7ID3dQfFAX3czsuLy8sOjCKTXasLVPoav0Mn0SXM+yJoxJmaBRpHJ8
PM8E1mDWAsVu5aWcCdWdFFjcoqluFkSCMyUTvbb8NBaQ7YZRrAZ5fM/URg5Z
b3Eso1GQ8evCxH+NTXBiIyUQ7y5Llgskp2szAYsODRFudjWVKyML6qeHzVk7
L/bG8TGPQD8S9RII+NprLE84C4UMRPNgjXNIN86DokXI62INn1+ckJuXzfvj
/tTYUVYxVOGr2s9iXAUm1M7fInloZRLKS/WdmOJKDcJ8gML3rRiM/b0zyAtn
ABVQJgRuEY5uNW3f/EKQ+X5CBYp0A9jUEBIKuwbGHhnV/Vm1jYIR2my8xLzG
M3u6ju6IaCkJyO9/ojtq1suYHeeueJb2KLbg0i2lhKIVvw3J97zvAJh3nPuC
FRLpT4F1IFj5u39DBbB3NWn3juejsJ/1hdzfYYyjLban+648pgZrKnqtljhj
t3UZhHAgGqiMbVCkSMonR6l1l3V0RGVt30KAgshB/Qg65XnPX3d8x8DmDDpn
T3ZpcXyGGra8Xx1gFl9g2iOcxVn/g/xAVfAZs8XW1G3N4BJf1N4+kd5QZTVU
Z9mOe4/DuWv5As3ltbNH6Kr23+5w6gNa8J+7sIw4Hj2BUgpAp9JSq+t1KL3m
lnwqMa9ORoLmOaFRfCnn6aVwVAaTlWMoohJgR4LLeloJah0GsxD1QlDQbv5f
gY9YqkQErnWuPVyrdl4pRVL8mfCI+vfw0XBb0wc/0dLwey76jD6L7k2ak8yb
rsIEBquyVrAzIk7Sf6r5B9dkNxYpD3nctNEYLalawj6O972Bc717XDyew8V5
fp9zw5OquGkTwU3P+RaVXqxFn+53ff7xVl24uXx65ranZcf8UxSqhoh0ESs8
FIhy9WikZPJIYGHVzK9QSStjusgcDtrYRqiVYfh8mTfcIGdiW0tdRHmHVXXO
ZsCeCsUmlCJ1P7R/NfaqYVRh694tge12aCJYDJFRjD/CtU/XvUUI1y1n/51B
AJkhrITCYutM4MEM/wVpUV+RcpCpEUNz34Mg1mI2e1XtkmcaqY0xXMSX/QIH
2BO79Lpa4TjfOEdZClaGLE87VyRMuM3q8IviGt1aU0e+gEAdpzNGQlfqqQY+
YcYi6JLBlYRv8N9Ge1kAv4uQB91Jcae1RC3hUS+JeWY3griWTPcS6mjyA4ST
rCHJl6h77wwvzHlG5zmgy0aMUd8QropvdAzCAhVxJe9MPgkHzjXhp3VCTF84
1AaE0Dyd9mfK7Cd/zwaGmgsugcpH9sIsooTLQqYV7TloW/tmT2hcN05y5u8T
Qx+ij9uZjX9mrCFtx9nEceexorVv4wz6WqeEIwTWl5r1+nCE1WUyctRNucyg
qkLOF3DnXagjyeuZLUKabMyVS7hQwrIjkXlh4lS6kNZ05EgVyeWnybY6me6Q
PKHoxM9NZTaY3pQpAt+Ztlufq1uSiqcmiyJR8RpWkF9w+wonKfGjoG4/LZb1
2T5cZWp5bG3KetEAxIEQwbHYAL1gSC5+mOT9OC/XdI/dd87lsyOPMpjs156m
AAfjsDBbjnFPYB61jaIq51SgHDi0bxgN0DgWwpceot3S8uLd42mHfBpt9fAn
R8EopeesrBWH0xNJw8DZBht5xZkeszY9gSmkS90GmRonD/tMy7TrwjDRTbUK
Uv00POYHa1WhzyeFjBaODRFkL1q/f6ghU+3qCuDWTUF0Dp+wHVfPU1JudsO/
TSu4KTjJKtfKI+n3KLKXSKt/0QZWWw3Kn6d3n44vLYTrbeTHGJBv56072CwE
xiy3eUJBtQXkNrAV03Qh5PYRFKLoKLYl+lq7/aQh+1U2nI48iPVUIHH1v/xR
DdAsAuxG/znomIBROmD2wkOYnMC0zArp8NPgQNEZhNbYceYw5ygCzkp+lVIy
4bQN0+D/G9g096i7nrQtyuORYM2TTASxGurjEVEwYquUOIOiELkJHyvRi+zP
rTNVSHujdutPfHSopeMLoLLFN1Eb06U1ISWF86MFux7P7jjjku+2/gePMmee
tj1C4JjwaBxpr7t2o87i9V0TU9tQNkQLkjnBpohOEUb9DyTYQJCh/EQQ3laZ
vaG1QBfZqtlfHhyxVZwKmYk3AhBW0V+GA0ylvohYv5j+fSGui/u4p4KIU9y6
2SCV+5EXpXwTXxRn79tRFSHYmwUDokrGoW4yBpTC1lB/Pe5M80Xggb0pRx5u
rZ2PLsuPL/tnnwkRr0Rx2RSGVCPBE67Afnz0BSmHy+kWDuf9APDe2PuXHvrH
Q37zh6LiWZsX33iSbnP7zr9UDmQpXzNMp2i87Bi00k4ZzCv6vnaR34ykCXTl
6RDKUeHLMI5VlBbSGA8irDy9xrTAc8Oo5tvAA0p7WVI7KJ3m6rN06bP6lvvC
ZIacDGx4/lbfWQFeINH9XNBXTHmG1K8vRFvXWWB4GnuVSkqP0apzAmuXnv0A
GBX35szToZcZ68QXvYdqbeJ9NBiY6hwsui8kNllXFdPYVG78LqfpSw0U5c9D
XPWWZX/70+hNJlQySKhxiIC08latXHn0yY18SjA+smPENObgPmLyZffCNCzZ
5zY4wmfoWHJ7O9YTyyZoFucocGZkaHqYcrJXgdEUm2ve+xoCMH55rP7t6AIV
hEVOkW+PXvH0TRi3fl2bBNs4ZydpShCyUq+ptnAj/rRDXE2ppFgMWEB368fT
9BqZTr+MXzQbUhxvQyjmw6ZsKUFQ6+GkOSKH3siTQWvsHi+FtmiUVtI/MxWp
V3ib9jEbrxgzmSvff3w8oZ7r7t9kGGynRJ5JVIc50wXsHhkchcMlUmDkB/Jz
MvhIr3CdsPlY+FEaFdQa6CB8rbR1VKMFKGmsznwURO+i2dMugwsIdBcezdKQ
HO+8KQwlTmf2/S1bYurg1jiL/O+AVxlJjoegtQ0LaHJk6Fhme6eLAOTIdXNF
RUTEHJ/rrkiwIKjpZrCoGgAb91yBWMx+/ZShWP0k7QSQAeJ4qDzyZp7ZQoDh
jz5Gily2gv+5F/50lptb+oDGYBHUpp45yHBc1xecqRFy0sBPxKHjbLj9i0B9
u32dRuir3JWk98lfgsAGoewp7gjFpfuw3DSeHV//bvQVF6RJUa6tuZRQmYx3
3ogEMZ95D2kU3ClKbG0qkKuZScHNEJ5mhaoVht1ejOuNRbCnpqYXqk94IptT
UsOzjW+/yvuqA0slDDUhGuPYV0vldIasMBlTyZoj99IEYmiGowmhh4mghMg3
mMQCOeLtng6ZqsauRy8y2QWG62gDRiKzzAghtFWHvrBYtflO21hxj/tGjsM1
oAQtdlkHff/nzpMSSMaaijSz96pfWIz21wt++ICxraKblTeQY1d1Yxn8MZR9
n5enLS8ScXGDrfFSIJUV4uyVstr+lS7xgdnJGnOcJKRy+j32KZaiCP6dr5Eg
riJG6/gyMJyOZFZgfn7IzdRnr0QK3G7BU3zdCOuPK9nv/RezkcDMnDWwGrZJ
S4fAVjUsQnZw+0bgtQaA74ASgRmcaQh9Y0isUlSb5y4Po0g10aYPchYR6mlD
kjeE8Es82VihzY/wZsyzJ+BvNgE6wjrZpeNAT0dQLBE4nE5Ts5XznEOaI8Vc
NgnDYhIbxI7lNg0jaGdYNVRGquOQm+5+QbzFafG76dmPTpFBFf5Gb8Ak9SuH
WlfEkcJLW9KfOm2e8133239efpn7vs/JQ1XXYW6wdSDIkLGC3Pyp9aTjWcxO
CaVZVMrMJO5ATDH6GcGbNSNuTTJaLKLObMled6F+EfsTdoMRiWlk0nM0GfjY
gYTVf6aCmwNl1ssrDfm2auzBLamPaOah48meoXMX8SeEIXu9v/emGjUhPYs2
LLV5ycS7296M/v6X+f2BOQCDXlciaKMMbbU7d4KCeZHgcddSDAtuyP3PqdVE
PPl/XtCum/4hBCGvCweGS8qS9DTy6DluvyPILd6LauDVZh/8KrBLYddq8ZEn
nhjkC4YWsOpyVxsZNA+JMri6R9sjU3m+k4kq7dgQ9ko3GENVV6rmwYtwZ/cS
mfgzqF66bi4xuH6cqHqSuhzRndLae/98Ft186miGgZLeEmPf71bfcrTcCuSN
1AfatIsiIZ7XQKpYhNaGhLkgSIgrWrMl8GcEACqguLSvc6UYAr6XoxWEnMou
0fFGwvi2iYrNmrcQJ4lMjdr555ErJX78gHS8rYB5d+/eoQ6/gUt09BoJFcEm
xiS86jeXIGp6ZQMOY9EwOHPYabshStmAUiForKoPBhR/1E4w1T0NCA26NK5b
pddyaGITD398KyXvtn66+TEkIU7PbyDAaZa5lua0zujkB4PsY4pl1PwQTPOn
/610eW6GOp6U5rzF//XFxSK84Mf4DXwNoN4fe+tV3er+5HdvcCh+Ctw6++Ax
TYsOY97qpFZOaQJ7tykTAK81c7AnahFEjH/Lb7ryfgvGgbydboMcIcL2Mztv
l+mrMKRrHG53d9sCmpw8AmIzmbl9X2rMxcz2eNyRcK0dxOnkfsODczoBuFIa
m6GQa6ZyVt1u3xjYAgR+kiY5f2+10gkAJH2p3Gf7jD87/UdGaj3vV02o9f3J
1TzIlPqZws4pjej2NgfkI7p89gmV4Qi1l2hpwKkn1k3NILfgROT5VeegvCC2
6Tr3WFX2Qm2FOzjTVeq4s0Ga+8rHNu9rppQBiOp2Oq4QeskeZbqpdxusCf+R
ZF9/Ie43T9v03L1AkjOzbALiOl/tnPiKBzHyf0H2KKoFoduvfZ2yLBKY+Ipj
SFyxOjwciYbaDAqeHTmcYcZEIhxp6A+Sm+wTc5QlmBk/3NlTTwiq/Rb1A3aX
mf82nSqZP38byogpL6R+62T5IPFmAhGme1HDjbmkt+2GOia2+gBV9ZBmCfdw
k3vLeGnMf+SgaSKqOHjZYXKXoKBm33rFh4pNXOrNO9W9kV9770B0upNeIEv+
ZO34zy5pCloSVpZrwdNpESgghMfz2O3S+EG+ETcXwe0TeDgE9lqW3sgnz8kQ
mg2e/jPuEx4ewq0kHPbFP85SF8tLRrsEiHnnA/Sf1tdhc8r9yPSpqH0BjrLB
shtJGzun/N7k9rhRfkI6H2vk283ups+vuqvep4BBFVQD7DNHwV5uAQ3UqDLd
8xWimyLf/nr1CpBSUOJ+PxNdO2+MOkLpuXzsrQ7E3WjA3o3FEqWXuTYuXDMe
s/qvj9bUE0JYYPyARPDorrTsr0iXqdU5yLYQVKKxP4H/GngrfEXeIMLhyPEG
tJp1oFvWSuRjquikSqIFOAuFomWSPRgvjldS3YL0N9CU03THnW96lZZ/jPBq
W0rPeiTujQ0prSGsE3OkgtwVTBwIQtteePHz5ALKAWijl9nsJ+l2+jdJfvgT
uZK7591YzDczV36H3uvAbSSszSX2U48vpV/KX7AKYjfFJNfZ0t5HtV2TfNj8
ZfOri831L3B3N5/4SRXQ4GDSTZQNStsRoe34R+xTl7lt3HVKwg/goi/bWKiA
vNdZnj1kbvOe8FsUhHLHnYXD5HC6oISiFqnh2AkuzgD6YlpPkcWYgf3Nq/1L
qaXnXDF0DqMFZ5vGBuY5UAefSJ1ubOKUxnaHZ5YK+HVo0gXADyQ4Ti8TP1ik
LIui0EyChdRIHohmQbX5EhIgrwRhLEYb3mWOb6i8qGiwzWQnVV8rJbc9P6Pz
y1T8HQVeS2gq9yLn006DncAFCZzLy6d6uaI0ijS/BO9+2W9WI/1PuZYZ0JDl
816NDVteEvWxISww5CPaHkvqD4i0My0oLbHqoIWaHG/pmV64BryzkQHtHDsK
uu/k5umUxSXejBKOaGWhUx5euUzoM6rQNHNyzAHlap3eV5bqgAvEySn3etis
r/5QaCZYNszNfPmh3X/PIcMlIK1KLrthEemdmM05m9omUaT6zfscT4xZp05Z
EiSxB1wENicdjWPh32awuMEbzr8aomzGY5OhWpS+43AJtIy7zLW7tOE4ApoU
1NwpYh0sD6C/qrMFnqtM1IiNuDZU5DQcy0thuAGe4WAyFYbRLOOVz7H1Ctw8
p2oQjsRcL6fDI/qQ9/9WTO1yinOaRfaHaUyDEWPq/s74O/AprJ8N/96hnRd9
w5pxwmJRZIwdMDUQaqCD2NbNIMz9QM6SyxsIsoH7ts29jG0TTaioTOmNNu5A
ydjcsV+bN0+SG9dyGJgpb+7KaUQjSpWJGvxUmWDTTYeD5aZcQQnapDOorqt+
R38fXKFfoQG0wGl3VPdFU9zqxLTktlYW6twRfnrBrDN4NH5zJbzg/aXpMuQ5
Cti0XZUaQm+Ua+TGXqQqusN025/H53tZpKQAII4wH3QRKNFXdmv2KkgtQJbJ
dMjseDVWhnB3/ZIHpdDnmBiBpc2NchguMIqiERTrTXhuiKB5IMkqB3rzsKLb
v7185YDweQGfHL/pO7GemJfvGlLiwtwLW1x/mE2MnYAiTn6FTVZo2A/roSuf
Pch4RufFWMZRQUB6aSnVHcaO84JwJOcN6vlDpAPCa1ORjpmSfLEKC69p1Tkj
OLJXV1w/4i7UdYxUVyx9bm+o+fvIWvXjA2hsjEAwbUJx35+aencJsFV4LUus
CwBg8lnLn4cdzCLpp43Ii6DIwIKlUvViyVatG5EHU2MMfP9WSHINGoepKbNF
VBru1jcuM6IgMx1OCkHTu9yA0VI+bMqay4hExsqKvn/1e3e8v7BhfnsHTf0V
dBxAQr8v7LQr3Tj5Ak7/qJKDIlHAkUOs16nAxO8iFWrqh5KPTLB6Sh+ZtJ2J
U0QqThh+rJIPMPMrPMM9c7T2lLECkUyNdAIUZBGCITillJGBxSyEgm5aEVrF
fMEoycU/KsGcxi6pQVhRr0glLSj6oBg9jqPVRw2KwuHE0cSt/5zlHwcbNQvP
L1+YzF/YQUMqHmHVb9/xpNeXWB4SewrWdqNudrJcVy+NFpABHpBwgIKDUxjv
ORTTCbeZXZkyMVJfG6fDPA4GhAKSsHXN/GU7wjzWKiPLGsuzjP2hnuUnMFsR
2EYcYJz7I6jeC+bPC+dntVFN+9iD5mtIQed/aQwFPcOOOiG1I2ScaNx4M+kd
Xvt20IVNgCvQxSm2gnplLPzRgKlKrLOL07bL5u1I/qLalLtu563C11t2pQ1n
og/zxK6zqTgYmaGF0hKGQ2CuhlabnEsx33/CWj2JT5xBJ1N1rQQQso3YJxi/
IiVSlim+o/L2yJreLUFu70xOFhi5iO5bNTT57x3BfO03AWduOJPkIBygeY+H
BmNzlIJYVJbNV5fDinzj52VuZKIOQPFr/hS2zi8UbEY6GJ7BuroYwfxtuyW5
wVqp/KgIwlrGUDJGZt+MzzWa1OcH7dlogcpvq4/IMN4iNu6mVTmf2yXKXPkR
mmORhVy3EWxaOHPA/nX3TaABGzHW1rDJDC0kxTMNnSfzl7THzuxpL9LHOfFt
QKKWPJgNppRlyJxInSA1UdC3pBySuMRoc8DjkXLSgLavSYnoQCPQmljtIvv8
Rs/EEf66xXWBIHdGji69dSikE/yxR8NsUZMFrDG6Phd8S5sFhb1LaWbgQhZl
UoTuzIDWBPXYYq7iCGECaKvUnN9jO/2JPTT7j6idiqT0ux7jZH5DImXsxnRu
F2YgOVGpl/oc9w+JyjDT11NrOS8R7Lldkmh+DsTp+s6HW53pn2jhJlxa6eIO
VXXl4RV+stF0LRd5KZepzopRIfVx6p6nX/SgiimM24s7fWIhLmbGq0Ndblm9
Zd6aQ+CbeUSMDxiIXswI8diEB0a3NhBJOfBF1KjnYFyN4apsbjL24X4qHSbx
UssjHZUBqHEuuIZ/yTJQsrhWIyLZwek0pePo4kB3lyOenbfeMKb8tMzuuZns
0hVshnGVwl5tErF58jLQjDRPdK3dDTwpz7uWbGbnJD9wRv6dg0K9SEr09/CF
K1I752WPZamHspy0199VWT0w0xKA4Ga3MDSnUFTd5FZVfyIgaTT3/75QjHam
aehn3jIgooM2GX2Xo5qyfwaBFAPE3YV+baUsmaqtcp5ULa/32GNliouMZmwJ
xsMJjfucp+9435akcLHIaZllXtUtds9znfB9uzEsxopuKiCWnXJDv9JtXgTW
yFxA0zmr1PeZMcIPJDDzi9WtNljRUr92agX726nwGV/xHYLmsJ9UaNVQ+IZo
NZssBD4wYap2qtQa9BBIK2byFf+esHnp+B4MISPjmMkEmB2qeDL/dA+w/sN3
hLisIAzg45ZvjZk+UKGSYEF5Lae8kRXHx1ZGJCa9r1ACpF1lINgmJhA+6ttl
ADXYeF8JEz1NgoiJUT42JXTF5qeu7cpL637b3El85vxseL/kQjnr83cKvk5N
7DKiI2PkPRG0s1Ha9QL1aYI/12o8681A9xy6nxlOicTHW2uM0jslnkz198EG
luYjfkh6uRsFO+8ZT4HRArjvLk3xfgiX53ZrUF3YHumG9UIRrmka2H8LjIjP
cCUwg0WoSfEzE5+YfVom7GdxdskRLeQIm4Dq8xZWbH3WXK8lt6zgBvo2sDL+
+6LN9iF7Ai3qYyhCNIa6JNgPE6Py6rhI7/kPW9F5ff6OU0m+ipdHzYbCLPq1
3KgN8EsYptyPnLXKSULj2rOnO/+49wNvCnhHuAnshN3yDic628Byy9nwApq7
Q7btCDkntxG4ZErzoIK8jTqs6lmq/ib7UxcVWmGVB9frb91aBfGXX3XRpECU
IAXBWoocw8mVr9++SfT5UxMHajFLmPPFqri44MtzNQPJOJRX6ldfOJLubtxu
kdURIAv4ZHxcRV0v+hOLT3tPIiTt0mJzCitOSKSkVg6erQ+wOHKtrfH7JPtB
qBSTJJOXCaCngv+3YBlVZiFzxISly5UitW0MPj/sxbX36mfxI8nNsYSVC2QT
/a8yHSDH6iXastBt4xHlzqTAX0/J9Fq5LdKj0fFqDpZhF/a6Y3PnrJSU8gB1
fpXcLMfb4UzSM8ltorWFgzAYchO2fTG94410anNbLBzYTKTI4pzyfhRL9CDx
Lc5wldHUyl6tcodUn/jyGvtjgYP1aNijdRE6N27MuH1Zdv0Lhhd+6f7YIzzl
H9iJMrHOzxIHp15NmJLCGCQax5wMHxDGfMEFiKcU9qhqZUs36qy/sY1BIAce
YUDy0BLdLP/eC75EeUNMoInwfdf9eMhl7xLh5e+2wWEWx8jhMQV2lKCC9+ux
Grd+q0gGc1qixoV5Rtgm/jmthl6YkUd8Iq/su9TQOHEqCWzd8c0+gal5E+C7
v8A+QFjVGoPuXMQYUgNxyr7Sjef68n4z5UMNFFyghF+H95BR6F7HmwGEP4Bo
Iofnz68WPDBlWy9czGnmPQZSi8LTCQab2FukTNor3sGcQrS4/X8pOJZo5mk+
imAVVhFvzUY8D2tXJjiCY/YzHVA4aUEZ4ahRPG/mLpHDXYzKLen4+1PXp1hC
czlSlpn/u5tBIcq1cF4VlcQONPfely4ut65NUbuLKFT+lHGWr6KOmMUlYRwG
5j1uzQFCdHjHZOfRz+l3VBEimNnHd6lO0ywTjL0XrqeZii/olzsfFahKzzoq
Y7YJ/4XRT7xCiYMmcDAtCyhbYX6vi+h4zu/vuN5OSynG1yVhl3Qn6JqDLe8r
+rxdGzbx7+TkKL/2YCGgm6cxbjKFKdwfBC0XBB0yfCW0Xj/Pf8Bj/m+wufDs
o/v1ADFQN8YY6Erca8OJTd4L7McOBavY/YyEtoKuPtHsPOvXHgbrSkceiPKr
V280AMMS4WDJgrUkrQ5TLydy2rtgGu9L7pXgQLn1VK92Knd97Z83OM2JqYNu
rZ0oUoPL9FQKk4OHYpAv0Dyq6LVxNEvdPdwOvZ6z+P8YuVAGQYKRl5WqwClE
WSH5weZKtiGB/qhCa6stGUf34vfXmcEMYwm+0dr1cmLByrxqdW88usQPWVCT
UjHHHo8nRjGsQCM8DGjUGAk773imaSFeJWfRPhhQqtJJhIvHF3VjHA0eYxAb
FMwNXfl5weY4znYMzNrIZ4uswFIcYiwZEUTfUl0YnzU4usXuQyzCyJsx/wuD
qGzEINDNQxWWLVxYTaJLvqfOurOWt/gLNKkyXVOiy5H6ZyQzamP8Y5sK6WR/
Sy9TknyH4PiT4byPrR4lQ9sFXz9g64ooJ3Vco9IHecqnOGNQpc448BPhuNsZ
xSFKP5BMUETYclCBuR2GjG6ko3ICqy/yFshNLf/LnUYEGaoWi3yb7ksNUl8N
GvKbSS750mwbKhAADsifk0+s9RhjWmvEamVnkTn6EvyW5EAbz4wI6+OQdvhf
IpiFXRDL5G43c+jFQsYgC6B29N/Y14DOuX8IjNtbZzcg17cofh8V0cIaHEBs
wBFOCfuX+sJczHS7X8E6SOB0FBoJ/dAMl5Qz4UjerAIGozpYZ1OuBWVO5FZu
u0iGoyvhxEJcJ5rPOY63OOcgAJWIoyBfLB276vt22u1IuP0B17YB20P+HLUD
DewOHpT9vTd67bJMyqIyRu0Z0qcehvubuSCU2L0Qf1mQZtUmZDkyPr1uQVKW
pbnnf8gMURM8Pn4UWD6jBFjZF/6icDZG7DDbG099NjEw4l7HgTvV8hHtVtbj
kn/rkLdvPVJqOruHanU1PN+k2aNYyiB8qL7CWJnyVaiXScDRTLKzX566zTt6
DiNzV9kYQKBI9DdSP5qpnzryu2jWP8Gj5FJ5uu8cwnL6eqhm7QeJ0PorwUG6
ueerOP8ID3D3RIcluEBk9cc94DVw6n/5PgJ7kCD6ypkGUkx09lnCi0ilfpVU
GT0o081yGms6ET+QecnhVnL9dzpvepTkTEEnPyw9eqaCO3Z+XwqpCwTWo8BD
GiPIGXFKukJ0nbPstwcN85BQNBC7xhymQe6CDulwk+SrSZuZyYah8+hKWvf6
PLSa/0WYWKrvQA1azYg9zBod8oS5MMcRhZl0oszefgmAu+BUPYN/cxu05gtG
93N0fdZ5r12ysSiUVmL0ylmKmr94K1oUMc+w9GA9TeIiIiRGcK6q9Igyt1nd
1qxhCs9OpN0mnpjjUHBVW6OFvk5NQDPGghO/BfbNQf9cXexEMJM2J/nm9N2g
ENiubfe9J7j0LEGZRGECxe+hGatYzFA1PrV1v+u8piP9lqTxZtjZBlW44CKP
KNEOYDMkBfydtrm51onFRkG9/TOSrrtpsIG4qHpT/zUvaPuIoCvpDBgExJJU
6TxncLyKezU3MXWLPZMv+K6ivF2RhKIK6RsO2xeyuB5lrfHbkASq9m82/jW2
vX9mwgM4AO+3TY8i3l3xyEnpSt8IcYu1HH86y7HaelM0PzoakZ1Y5IPhL33p
Mh2mtplyPKr+zSTMnS31CVHEXvF69xDz6AKh9uxL+TK9jNYJ7o5mhwrLnmMf
d78nBAxqKn4rzTz5EL3O1igjOXKRwbTDG6SHWss5nsVVmmvJUvu/09usjDRQ
OR0cY2WWLhLDp4IRuqe5tmunsV7IRKBaXVoqwz1F6TDq1nPdSpyLjyYcimad
lyq5yWZlpPfmCbl6J8JlaYkk9cqf2LvaMVMFeqBEmShcfa0XLgJ0UHLboZG4
T2nW45tabAEsvxFLU/srDv+Og8JtD1vV5ZV6qmSBRRvfG+YnQzdWq8f5ep+F
lk2E67e+RxyXGiPwsfQ77CXHC3tXV5PURPC/i4OOilW++HOEHCQ3d9PdSW0n
E3jVn0/UJzY2gAzUdciDVj2MJ3KNaxe4stFYA9Jpm2jZZvJlKCqCYSejU6Hh
vpCto+0nMXyLr9ADrL+k/MiCut+l0IVp81GVNZvIAZUkrW5lmi2gksIxuwGa
RqBY76sPnas/serpkebBsaq5zJZOhy8VsWaRFyu5++xEOrfh+f/l7hzEb+ps
4sb7cwqY9dbVnR7izkzqxlzXLbPg9bDxa93tE2q2Cq2xNBeH/u8byuWGVVUL
Rp4+FEj/6sViM0ilBCVnoyODoxiK14L1OwtjBkxCerkybvDgZKYqifNQ5cz7
Zx2YI75qAejchEcH7J7Gsl4Z4rI94QnYOiAARmTkmozxw8y9gx3voXFsJobh
MqxOS75pS/ZckAqcd8XwfT+MwlbK6Cg0bhnOCanhicxwODv1oc98OEeyalJ/
y8+1MsxQciRXnBfjO3YGe6JWgFe1JOpzKY1kXtrtlxYRdRo+PD3Zs9vvC2OJ
mhojtkLUw7rL+9Pii068alB5BRrBJioOx/Uy47yJTAvB4kbxCiTIQCK3QFcs
nKmq92SGW/qioq6uBKAsYs89U8F/HnfQku8nIdIcI5cFpAC0m1lCqNsSx1Xg
fNyD3jygmwHUaikq1QzsouaLFFh//58SX0l0dgg2VmN6MA+mi5/NBB4GSdZ7
1qq+d9xOfvWKk4VCWovtzlqw0vbQnFhVdfDKhuRfX1n6kFxEuzDL8tIuwqQg
46TK6eR6JywMbxJi3MH8ShwSEI5HRyBqEuDB60Aiz9k2va/rlX6/a3kRBVAG
3faezNcIM0we1yt+eaIsXWxhIQDocaFIIy0Z3ob2DHy8mPgmT4rw+2tc6anL
a5Pw68GzCWDq4FiMEWcZu8P1cfJ4vdSC5OEzh8iSflSjAiwVvq9egUvxM7iS
ifRVhB9ZOSq7Xo7DOdlrNwt+izINwDyAEQbXvwvYNZQFjJPOSVSUKiplwWEl
z9kp6sYiBfPrboEwzn2GzlqFvI+Oxnuq0Ase2r1mZ/vYNouckP23SJXeaX5F
FaNwaMSDpVjdCtKXJfETttX973XpEZcfTGMHFDWMJe7GALbTIi80jZ4iS5d/
djul6QisKKeHxFP2PKVbtEHOmNYw0CnCqYWDELJOuAiNpkJv42aTyl4TuFyE
bo4DgVQZfovVKlvHolN29K3cPfWcoM91LOCin5sV/gL37NjyW5LiWTsh86WQ
qrAUaVIJvnj7d1sDHeCo76VhBwSuFWD33C+kX5VGJ2Bi1P2R6JqHWU1f3byk
K3WMfHswBr2f3LhnD/F7ZAnXJ5OisfccRuf70OqlM40bMzcJ29YGvOPB6JI2
uOQlSZqpUkoUS2hibbG3U8QyMxBPRixg8Pijm+gwnxyjaoAT8BXcK4XXzc6z
+LE7866eNJAMWvFH+LDom+e8jyyphkDRIMFmcX1ia+c1Btk4GpQVWkGYcD03
MSh85xN89XdXq7xoNlEn/0n4bX4PrFw4qSIgdV+AOYK88nlatWdJ0Rf2JKLA
978LNBMpN/hkHW4QU52kucaEtvSJUXhRREFs/j9QD7Ku2jHasFv2q6es+Ra8
kGmdgN3yBufFmxsSsjuB74MhvP8f1GeNwIiWgypCteKa6ykAs5jxfuVKkCbf
zmydElmnpHtqDzcxCdcmjFIKwUh2iit6ZrQw2z386QKctb5SOXbyF9iFQnz4
hiPjZxCAgRkJjqqQ1uNGudI11Res9azzFpJoTxW64PQhfIL6jUAjHci9uXxP
M2NwgnvNZ8FzslWfreANQlRAIoqY7xcXZFvIyO7g4gQGocYKQUz8zM4Wpi02
kks0D+SuRXelY0kZgdrIn1xCO9wTQyO0J+IeV0u7+TopZ0Ytm2hqpRu7ixmd
BMkjT0GrOoMx5MDJeZ+iK8LsK6tjfQLblNEjHPbSvhOF8V/hB4auD/Jh6tbC
l4ZhkdWNqGec4d6/9NL0/2CprO7hiMez4L/aStlia8+UMAa7TAB2+FrJ03hN
c2mS6ikyfD4oJdkqnVcT/+tmZsQHi/sxRMhrhTP8mBdoMnzVK/VSXG7jk6oJ
/SFaqfR4oCQG6Kp4v7J+bxr38wZqn6WUEquwB9F78Svtbbn+s5F/Dqrl/bGx
xFtSUkBIYzN6q4a4J/knf2qsskOOyhG9q47hX1BU1VNTdtH90UmgQdXnsFnm
rqA9rLLz7LQag8CClBpQgaBrKpiX3EIAFgLisxfyG738w/5vqLk0Fq4bYk85
nFYlebZ2fh3/G6nJbmBkc90pLCHShbfOoerXPIy647INsYs+8i80u61VE1cN
gxN0jqKVvHU0OyEkR4zihpDF+ykk2e0/gnkpgQhcBi+F0fMCKPjRMM3LhJLz
qoo6g9T5YK1gSbhUAMuMb9Cdo+Bi/JWQSjpG+dzFNl+Ntvt/MflzDlC+xYnr
bjH+LRRphrNu1S4TolO2vh/qzPwY3Gyw+GfJxCM7gYpUvP6c27inPcrKDTTW
BZfpm3Mebq1mKna1ruAZKA0DhBvauoFfG/+ZOaZnwtLf3NxQ6fkbAZeObzAQ
vxVxxWXy4AnxNAkDu6vgzyQXrYk06Rn20UTTPoQ/arSoM40oigLpMbSehxpJ
DpCPzyEMYFJGmYEBrJ3vtpq1AzwQ3AmcJMjJPjjcWmOYYX3ItO2cKuP1Ql6d
SZHMDt+Ug9/APfFv6pD+5EOwSJMjSbm6wQ539akin7IDCMLwSBWxVYBp2y4p
a/El4AUfWjPg17aAhD66lzVQNxnnTxHeeEzexXQXoDmogkmno4U+XM43CSVb
52XVOoJ0odrhaSnrgDZWWSUD7PKGMk9eud8DxDt9p1+PsoetVDVLncoqmz/c
nEcWNKCb/t1xiq8dqql/4R7MkmbrHrg8R9q6SXGeL9JTTqXRwJQ5b8rgpfUK
SNZWYQyRjcLCmk2SL9g6DNEy+VRSz43icryGeb5Np93NzS4foS3FaqlmqPRk
h4W7hHbU7lYfZvNDaBVgvh3U28T9xPmEm5LyrsngGQxez1Nr8oVaMKUZZWlf
ajXVa9/dKZhh8IYBssDS/DblkIPVdOZOSHSouB6n7TrdEGwINcpK6WXOWHBB
M1avBVxdLhm4/aHp1oU7Jnr+pFCacWL5txK5ld/W/Bb6/Nf9FoMkkI2wBWNp
9lhds+pHA3rKDbT7iz6Fqy9ptQBBA8aufDfJOEeYMnYsCszy30Mu1gBBN2l3
e7qHArWXoHQUHgSOJD+jOhn9h0ifmW4YcEeuPiHCa6aZFCqap7leVT17GZee
/xjV8i0HQYJJoViNmD6jVV5T0gqHmOrgP3cpMSgp/zLIJXiZvNSJFmsH4Acm
4+4dLW4fx5d1yu72FLx/dDgevejxNPRRrMo0Kds71zDCGu8mf31L4YGQSDcd
dBdoOx4Ygcpn6Z5sW2qStk0fZjGrc+Pki7tiMY373n9X2B4gvlSNDisZoBGN
Uwg4Lur8DtgM9RdDYUPbGPiC/79bt/L0iQXFzCCNGzup40Hsa4xlA6SXlCS+
6En5cWhhew1c0+WQJy4jr/qgwz7inazQKwGKswKNdMyYBHmVzLxjQpAFCxlY
QuknHR741suHIu4NGWrrjsw+7dVH85i/XugTrHYz8rDY8M3mOUD+7Xpy8cKs
9hsaHf6q+RXK8ZlR78+8kUR3I3FhWgUwWRcT67TQNqlcnvw7UwciR+fkie4U
gNCTaWv3Oxrcmn1h6xP6cofgjY0dvWqCK3gP4mToXDsD71jlWuOjM3rrVyjU
FpBiaHw97LHLj3S50lM61jyrae21XJyjGgRMPDr1npdCcgSU6VocGCYeEUb/
NhpSIjyZjaRVoX6YxGb+xdUrk/lKyZVpdSiyIIc9QBsxIDa7T1G7ah89bDMA
6zJ4ytI5CdMpFPejPLetJJnjO3n/pFK2wSIGXcOxrBtfiJ60HSQGDEoXABtH
Sa1uwsB62VAIT0MhCKGngpZkhx5ZWLSx9XGYQXUI80ntsnvZb+Rr1DE2vCK/
V/EWL5xpidbW13wxxewtaTBHypVk9xHqxYpz3/fFUKc3bGEDZQDu6SdpIUhk
QKOYrMq4UjPtn+Y8Bpt5Wdk8+KaBGQybjUwVBR4WCBEPJhmcb657nTiCTVvS
zmstLMmuh5WXtec/Gs3bD9PycdKS92/cnLeOa/kJP477AnZLB2GAOqo2tV/p
Jn4/l6cnPtXnr5lVt8eWjI9WQfZGUn+cY8CYTMt4Q1ELaDfUCSjmUOumKNlG
PeqxVXRNz7F0wuDQk4vCqn7Xv7TX8i7GFn68ZtJtzfJIYhW04/Fxpx7k8FbK
5S2FWpEasn4G0+TdyrQ5R14Bs1/UVSRAqEUGd7LTtbwdZ3BxIMA/IEmumlQf
1opakHj2+X3NDaqS51ddZCy/FDVNDgOe2MR+E7TV8AipIfJ8ryR6yKxJcERA
ekV0yQLDADy7F/4rEQwQqhfIplH45QRRhejR0raFJ2w1ADIEGJMTcNhQZNGt
aF49gq+fpNkD9PHHv8Dl2gYu4SV67RgaYnyL4iC/2dsWD4E+oXvaM+uED5cc
DWMtHdPhfQLx2r8DojRC6qws1Cf5XMS4pQBlyedApnDiqCxl8Sk2NEAWmkiP
o2OVXfhikAoezKjYIJF5PMsJ2zeOZO++Ne0tUhuPKgMIchCf2FBhFykbgUro
iEvJXmnabmWB+/Uvr8DbElL/9KAtfo4aN/w9lh8yxM+TYoxKGKmGSXsyYotP
F+V0t6zz5c8wl8bS541rK/F07e1qrzwFgOfVQiMhp/tZesqNuxCsDHqbWUOX
o493Z0VpIF39MZFaNyw4P6HmMeH8TSnxK0lx1KmHHXylwDCawUR1M84RIDX1
caY/Vnc8jGp8A3BQ3KUasfTZ8djTH7vm4NtdE0ty3gUKzb0cAGJK4V75RfQd
d8SdBOV4yG6dmhSIqmVB8BDtZM1/0D6I+fEEqJNATJtZFmm3xYP9Wow5sRtQ
b51xnPYtY+tTlLOKZa7THiTsd2E+Hn03nPeddZqzhCP6FySjHUsSZKAWQQy8
CIqBtidyjO8Z3proLhT274w7f1cQimWWuWrLa3+rpYsGFk2Sw8pVNuWebh2g
NHalT2jNmvRwtsSP5E37vT2LzhmKkfGV44UCAUYx4wNUMFnGodIUbZvKAqkF
Oh1xbGaizAk3cAlJeGoyD3SFxdmUlMdPB71WJC6IojIGAhg5ZWEvpJ9OKzyU
q3XPkVh+MCrGwso07/9YaCRMKH97ssYQKlYTPKBm7pVYkTVyN0F6lbuWhJ3H
7Gy8pCU2WomY5yGMSqOk6PESeJl/HPZHB4/j7W282wJ7HbQkcUWGmxRj+tHf
WPWuKpy8ovSKJ0EugNqzVDELfyuX14n4gS67ohbLAwQFwxSs2dqPdn368YKx
5pV+/BFWi68hD6TEp6w3shlAQroD2/kbk+zSQDWbau/V4oAQKOQIByVt90O2
eb9g3yOFQfo11QfFcEuff5AjgLa6auU8FGFRqPUcHhHcN+dLiUlwCO2psvNc
nMcJeSjKkugjjOA4QuXW5SWJMPpZ6E0bFlZrI5/71wGf/9/Lz1FC9XiSQIbm
rNNaqLJ2fLPVoQ95/L18xBWgSHu5Eg7YqOwtQ3noiljXQDkWhkkYczPPbzP9
2jtCNiD66StiCoAWu5Re9Vk3jL9NDgLLPWy4MS9V8widWiUfs+TsupI20BCb
EvHVwGyFEzVl0ygCBuPZ9Maxu3rQM9uhRVlgndFKurcvi4NlRmYW4Eec+0U1
Ht+wjcP9MsAY0GTfk6hD7cbDxl9hp6yWNs4HdKcYkHgukCn4c+9nbZprvKhM
HVHpyukaBtN6TLadepHEzo6674BOi8mMtHrd57JROFF6LZgtDpyRuFmekHiP
cxqPA3vJ64MbfD/HyKCk+ng/eHFwVgkgqA9Ya2+jPm277ziHYWrhe52xjaFz
dCH9OzgtCCwmxa5DMfB6t/XudGyGAQkHPr3Nw5xY/4M6SrZeTt52LTInrHAe
UrVnil2SlgG39V5vDVXYOjJF3ccm9lZppNI56RoipsfUDYDm3vFY3Hbxqxxv
7tHuXzDBM8jSzR8S10UaXYHrDkPdc4wXxQV40l5QVVitSNxalI5TUl2c0JEy
xpGXpg1HtbWdWLMfJYWUl6jVJ18mbDCEcbfyvs6u8wQntZYqWYiaiPKrdsEU
Idpi0I8cSLHkAzAqv6HA/O0Xvq4Le2aLswwZtYP3tMivxh/0oJm31wABeMLJ
+rJ062i+s3+z6jdxu+eqoTJnjheNKERbNWptskiM8maKwkk6KsKvoUqeWzkV
WkdSA+2B1dloFKk15VQ25Q+Q8dAGtyibl6lkFONudVi4562Mc0NRAyMmac6y
bNpTRmaAEPBUDqDOPvThX1GvbzgW7h5+KczaRRkJYh9KHgfeE6CGlIEp9Y3k
ojN8TkZVTNF+ssFw254wh54Lz8amn+JHbr2AEqtO/11wNP3Arbyul74i/Die
ZsogU5YwgnY2dcSATa25nh68COEwHgQiHYzaoHzc7G369khD6TvcDRaK2pMY
iCeM9i3VmKJ3nEcehmyjMxoVQac4TnKklN3H/kbv/g3gbddbCbREqno/sY+o
RXWa3cst/dpxEaG0ZCyIBpnb6ME2oP3aEjvyrBEuPv9H5inbOojaaSixLXG2
HXkIFh9jYNPs9G6p1Lr42p/1NGyD/t6eecNPPLNud/4rQm0bmH3tnP/lU3Bo
UY8Hq1UVKE2u3rZ2fnQhpUIXceotmMJe6HZ/esbFT9HDUF1drMlEia2H0H5P
5KQgn3/aFy6FQ57V7yr/ClU5HmsPwkAp1wW/XLoo5BSLQQpCLl9YQ4u1bia1
Nv5hFUi5FW4VdvhxhVoOUKK44suQsPctl36nc9dwuQNypfVwKxKN/+deTyqF
nqqflEKTZ9LTG9vU4RKImtp1DU+H6LH9xJezkHbAPrD41ER1WgE7YdwgX6AC
BelSO2GEMsBnJgfvPk2EEmI/9ygmy+ilj/NapT90Azfss0u0WPeCWK5ROS1I
4ZC/Ic+v61vGUfOa2Y6j2HOkTog4bzMdnJBaJte9v8RTRUy4xS2H73xysQNf
R70yVCtdcFcbWpqyYyJ+/P+zepth/A+AjxhedkWJIl3pEkXVp04hRpjMmWtX
S0VaEz501L47VEXPWW5Vkv3NJOkesrmZj8QItCdwgDzxY6QhdWLK4Svut0DY
Ul3iLlnsUdSpmyKR8vk4HUzD2GBX8EWAzWURyQ2kKj6IQ4wGBaMPW+SaLd8h
PWJdG72cR+AE0tNEaaf+MQUygQKUTxQM4e5U/qAd+JNhJyDjWDa1f0ZiXPdS
YUe/6KUnWLMWEWiz/yEPRCLJoyIRMMHNwhV1kmG7c4qMWOEuXCBKLl1FVUGX
FrNHfbKe4mKAsyI20NOrUVpTnEWvjgJkqzYKvhfydF+GLlzEuZipKNccYtMx
mQS9zM9PzX13AMUEDZY84bUveBQskixkWiiRBb6ZMkGghPrBApP43gtJhkGm
/DhuAuAiQG5RDUShoqsKxySvUp/eVmxhJxpVTeplXgQNRUhVxnuN+i08Sn3r
4p2dnDeePOAs19qQgJZH+ZrpO1uYGLdPLZy2zOg5KamH6eh0o8wjph2glT0g
aYAifUq7Db5HVb19cUr5zJ4n+eExyc79HgQrLQ06KiVsPmoeF13A1EZuGOAQ
nLoaFnVSxeK4GRxD94S436tWs5zMyKDf4p5UIGlg0oFagM/bGH+KzJ2BThCk
4oMGezOsKfRe19sXKrx+zzdjnSEg5m5Ek4TRSwEzkWbh0xYGDv87RvshPzEx
FckP07SGfbEQq4P1S7Hum46CdeUYQd4hCHr0heGnWkyc+K9vLQCgy0d9hPkl
F82pbHGfguKsQ1zl4ZyaBE8qm+Cocc5Z8S+jilLG8BraVAeWbsRdMBjBQwKU
VkdwxZrMNtz9eyQnGy+0PyUnGTyJsWMyH/GKx+Z4YyQpQeadwYZ7K6L/zmge
YBRzVDylTcFaeEmKW8QwGPU9fj2zZssmtrMbFpcpjrp2tfjF0+ds/ObU1gtW
fpA5YqrDN2DgOEwhYbeEaVB6f7kHpITNXmWsqHAmYXFTBqsJTkmcId3xY35I
m3okbC8MAScIZnnzljAnzMN5gUHEyY4mXzaub72gU1bu11MKTH4mU/9KWvRM
WE5nhe4CrdCYdBHa5YiCE5mY4+CCIa5w3zTU391btZj3S8iTnERkxd6AgTjx
ZS/l0S6lGUT1UwpQwoRb1mANJ/aiRgz3JwpCudpc8jOuEVJ1ThewbD8FiG9B
HQgTZqOyTcMm65/WpF/eAW825jHotMUhWk1svYXvcZVIGkfvOOsl3BtHwS+j
nY5Pvjub2wk9SXEHTM6xEvEhlQc2DtAR2n6Fj+wzWwNj/EORlqf2s2T804mT
mssfl4n3nsFGMA0Qy5KHHc4L2m2AjaQHf+YELIkcbBAwaxSp8IS7A/WyRrRB
QwAsOiBl7RGuNLDpu6/WhIooe2oIqo01dfkusk4Pl5aGP+s5dsIXg1uEK9DI
Dy57HKFdC+EVsz/5PTbYK9zANV76w4pzU5/mtmhBIKr6FN9T6zc243wu/3Yx
BQLkQ7QIVzh54NRhzPvikNBJY0G9M4zLEpRDpliy7A6I2gnc9NCPdWnE5m1w
1uKCMnlr8w5d7YjViUucNdfE0JdQhEhKCwj6+WHfHD0t2yk2nWhCRrBWLd3c
BxIdgL6uSW0FJ8kKzC6kWqS7F8vXl37Zdh1a6z47zpg3yGe2YpWnPcuJgoX0
Uasts9agQqz84CtTBLyPUHAJKP1/fPdFuSq4bxuxK+VFgzrEVpyy30gw4Ttk
ZnQM9ITgRvO0oQE7RUxMBvjilt1E1r3Y7jsOJd2K6C6YEFgLdJ6agccYV56J
LH9eGc/DSWUpzt8IKgebM0omrkycy2cDZ4QKG8aMFXx0NIHQgZqmYDPqgZut
Mwxz0DxfmpdV0kvUhXThdmBV3AL/WFGRJwLMZSVF/8mEOMfa9Srtz1AZ1AHw
2Vbasm9104L1fSVbxmFzuo8rBeUFx6ofjMEG8mUSOMKyYc2JE5UnI/s/7xen
p1v7zhscsRdWEubZKmO9ZENFp++G1BcH7duIhTJi4tDcZq826oVk9ktFkTYt
e7MehrujCHyKf1ZC69OgF0D/J+to2TJxuA4ycVgJL2pMgMcpHdSaknfpR2QC
+MnL/uIivc0gSqo6D8Ud+t2+nMbCMkn4WmKQDvatMqmH6t3XQnavWqAgtbFC
r88BKIPTtRKqu/1RK7aO46AotdvkgQrhWMJtOkYo7haXru8AMho1GjwG3RZ6
j4I/SIn0S0mPDu41Pq4tJ3j/6Flszfx0mhiCJg3tdiFdPqter4bbEaHhgjXb
T2rJZqjttq0qt1vCsZDBeympi9IRu+dMsjUADvztqHA3uYeuKn4eHsFu0G3g
YB2d/KMOgs8FKtV0cv78GUqaUTbhxd8d/C+z8yUrvHHNkL+vKs3JU1iRAWwv
emnSJfRMH2rAZN2yIRf67ldwtM75TAzaQffx5Aob0RsvElWMfxY7pVn5Fjls
2hzNDcN7CJYWPfTO0s0QpoepkPDfKe57KeIdKXhyEi1CcdYmWBLOL6nYpU4G
lPPbh2WwV1eqz8WqyFH35UBljt9+ArKwgPm50ds34Uq3Z19LjsEbVhknSJ8G
q+yfHe9JIng44Zc3kPbRSAWEPNF9lNFDOQH+MtE/ypuNsG0wWz/QXiOAQr7K
x/mDlMg2EC5pXa+ODJbpqKua35KubVsgLzPFD5Y8oG57GThLOIUzR/nixxEC
4H4MP+HLKbUoQbByM9urAGIhLHD9GRQ94QRNMkEQ77wJ70fMnj0k9m6YwrQw
Vy/Hfa+d67LEtO1buKCLg9AVOC5SBB0O6jy/UsruPeCTLptHBjhYrYVeotHW
7GOWok7Jnsnmuod4JNzhdwH98sfh3cpZVp5Nmvf6Ov8wml/Y1FB1BjI3GSuj
8n+NjRv0BwIm2yGK3qAZB1Msa5erx+7AgTlFQoI2s7mpy/PlRmfPcWm4m35r
/s1JkNP6yNH0AuSxcECV4LuJ+8cS5BZ95+ZlKdUy87VvhvqAcFMK9jXab150
IwQGRSUZuOCW+RZHCGzSKcYwm7cEChlrE9ohIDNUS6hi6bRWj32x7ewWaEWZ
YZNVzaYXhjA1V2M2OvhA2ND6Bq6eIHuVclrhWE3iWvIq2AkqBDCMgvM4xKC6
ibcyeWdYp/EpopAF9hJzz4hKZewmMH67KrmoGbzmwnt/MXaOJMgZmlrPZtr9
8rfVYTpenuP4QngwQKT8971w9ezf460CbKyp/kIGzA9d4b6pGZpzMIZmH67o
ldAc1J7EDapBQVCHRQM2tzrUFUDZBVcOghKxsWki4xpMJWli0la0S/fDIzJ0
mCMMV+PqXcYJsw6UgFQ5pWiJZMloZkWIMjKLYV11CJjEmOXiHfDolCqs4eqk
7bzPDzcjsuH0bSNBbFlQkvovfUMAMOAW7707ejyZxnOAAuRWilGKYKAPbPPk
7fK6oaj5TvsDJEnKyC/E15HxZQDQdYLVjOThVo19C7Lm73EDWxp6e3Us1R2C
hvNta5V7emfHCGfdx/RV/2sOs8rEprtcesbTgGz2u7GTmR//lKZNEdKF46Jn
EWPWZs6iBYFCV4XGBO1r3W8sWLBZ6JBvu8G9fVqQp8SqLra6Iu+x79dkbACg
yy2WnCEjnbyqE3KnxZJDEgKAlhYsQFRR5fYNp2RWugnpSwbg00PnfNp9dkb3
eRXPqxYwmBE8DQYxkWr/yAbc0quvaCgLgAr9pdlUjRWFPFRsoLKkKVlu0xpE
ViLhTSA9FvjB0/l2dGcxKSrKGYyEiVnf14hl5s2lcB+5RPEHZSkcsGnG1vQr
mnhcHdhR5tR0O7FwmLZN8t+CMEbcviuc7l4QLIc4MuHs+9TyJCA3lL7lV9Rh
nQ4wwA9E3h750WUv4U+YiYRwnMghqO2EOvJAHI3weTdl5psfGHgh2oXQs9XZ
B7dRB0+a7MhefhA1NtKMiFsA74dzEITRNMrm+I04+ouudWQlXGn1uw28J+ZM
5tbH4bVrVmIxlReM8Y/BaWZedPR8TFG7bhWw/8pWEmyPzxisrogrzBvt5esf
yzGuR9ztLlTygqxXt2PFYXGK67qv+n5GNcpsThbPyZlp/8uZ0wX45P+cKedG
UZn7j+CwsIfAn2xccqaf2zzciXO265I49d2yEiDeDGdH2QeuG08VTK577fLB
4S53th+JSxf4+kWwiWPJ/kBKoL8hhEwis+pPRf0XW6QI6WdbL5ecGxJAKjI6
3n/BW0mudgLi0T21EmSIORR8JjYtxsk4Zl5cAUzXjF+m/aeYOkoqAhC2LzjH
qPsdxBBfdk+OswNaSlrp9MxiYkK043wb7hLL++x393YOAG5U8k9MsQY4XKUI
X/ZZqMiFIsGfBrMfE4yLk9b7SwRv4O9UcEkLBU+JUnouuAcvVmz5IYnsrC3Z
fXFNAQ4kVllK6pLgWNw8ApUKic6Dt4d6M2sPrLWNsi9KU8Sp9yVCQv8H6kV2
h689b6KKCaaD1LibWkpt6esZ+dk1SUhbAkciWoO/Jv9pzkl9Y0sUyEqEY/9k
dT6jyvlhse2HGjh4tEcp+uplGJSbLreleXlHngdowj0bDIHU8Pqii5c31vnD
FhI32zI4IcsbU9yDoyQlnrZbakOuZ99/wFTSLLm8X+YQoxwkjVAKHYtCQt4+
Eyl1/zsIkOozwpft9Lgf+2xdrpkbeiy/WCqECkWEQwSzUzBa8VOEiUyHLKhE
lQrhmuS+8bR9M3yXzcoJX+xOXSr7X94ScKD5nb4o1km81Ae9VVM7ByhRmj5L
ehfzS7U3rHYxuEa+/0P8cHE16R5yVI9Db2wppuTjvbRqOvOFBzHnlv0zDITh
UDtjuoipDKWVunwOHC2BsCjUqe5XIINp3jMR6dXpjvpedT9TWQWZQBYF9XaG
cc1ozqByL64p1GZb6awX4xtYQod/phDMK3w9ZjB4lH/67devpc6uN4XcS5ny
G9coYqTVepFHsPv78vKgKfTI0ENulFkmcVTKHAmN0plJCTtuZdyw+dSZbWbW
lq6fP73bUXD2SdS3nhKY3cDBW8lV/lGVUhNWT6aO4Lmm5inWMJNuEsL+nMCq
SNpTX3doHmCN7iEztBues7GENJkCdlFTZKrTZYRqWg0s379mw7UdMl7CefTz
7gn14kPZGp3tkCpOIIryZmFuISV8epwWilR64WMsmXFORo+PC6x7+xddLKxG
FYOERZ1YzfEQKBLSt/D9rMHHEuLo0/Rd/PAMyuBqHmZWLpQ76tvirzce0OZQ
k29rpeL4q0bgmnebIKCsWU2aRi6axW20EJIIFs4q8olU/loGgFfhrViVS1pL
6q2SFK8lp4zzPBoDt8xdcOL1UQClu+ia5tNbpIR1bYGYbD/swPxsHV4Qz9Gy
RFjpPf2SSMuPXQbB3H619YAPtcJRhKFBNkGMARsACE3z9tj4XgIsNDe+gaA5
ElhtdKgv82B5gstkxesSn1IMVcWRoyKjOXByAz3e2U3v+3h35JyAiUpYK1cP
qnbb+w8+mRVxJYD4HzblA1rwNcz0XgZGgaw2DNVSztFujwYoO6bitdcOkYfD
bjpE6lxBV0k/DwL3gfwkin81jcaMxfYSIyto0K0eIZPJ1XtxKOFKaKoROnUq
AJX1RXPHRuLKfex113JiRlian//6gFLCJRSlgJDCIC01XP6/btnhi6P7RAAv
OSt41e8MbQaV52nwsqE3mbpvo/txWflsr7fS+u2qqtU8PBTIUtm5bI3RccEY
5RxyWCgX4YK/yBBcBZOYpIIuURnBHx2e7R9VpgX+L8PTvQH3ly2XQyZbGLP/
EB1dvEanHRN/Y6fbfzjtB00RU/QDnT1TuqaEB/5jZ6mEiP8feetF5v6gqyvJ
zX71NHISy0psc77peRIHnEi1xo7f5KePAhdzMhxu1eKun0D3eSHwZwtxv2vm
EixO0mRjtm7ANC5QDuv2NUmSWMGsEYLkjGj16TfBQc2Wkv9UZv2ro/8VoJVB
h07HeFy5nRGKJFoidmcpXAUFpGjTfj33oMjB42ghxlG3gn4YpwDzj66d00NJ
ZcrWERNVLmA3WqQSDmNang/ftLowHfpCePN+lFiKFTBXH0eVqaPLotxE36Ab
54Df6WxAYMiEO82pCEzYOcHhrR8O4CelBuSmOaPhDpXkSGtx5eny2quLqd/U
UB4NTmeO4arSOPYFF6w5o2StRS4plrDHLGdrJuBPSrtWOykWHoF/rqb1bMlC
MOVGTilPpM3URVzS4uIbPZegxNRw28XDY57oLqm0XUXxwvbw1rhDcb4/GAAo
13tOLRLSWWmkuyhkaSJOp4EE9GqgFGJUe3AiplCYVTVzuTIbev8uvTVZlyDq
And9nLEY0fiVzHsdAzQH+D9+FjXsz0M5IE8cPjyOq1W6TJGDPeml2ReUDj0s
XcX4owDXVgu6bbCDK7mRpJDflOpbukdyyz4vqblUhWFTkgzjFwEkRZoRS1Ao
DWI5aLgUaMowc/H4Wo7fEXvtkvtkbdvKDwpT6NCf05JhT1EBWEDdbvux+G+O
seBLedma7VVk5r3BmoWA1scVZiYSyScMK97wQHxKxd3BTXc348SljQ/fzLJ0
KaGEnYKozT23yabn5qbDvlhHFuvIIa0uZgPH7ip1Bu7FFjmLL0VVKTPitFRp
OdL2W7MHRa8jRXuUl03Oye/dYqOTQsL5y+M6AHy+WSFj2CsyK7b7GvDIO9dk
zcesToBcipHUSGTuiwH9L+/T0VKFqQ4Oq8VwbUOE8xe3ej7IEKUZxmOsx7dZ
t6oJ6GdHAcHX07ZEFVoSvvheai2f2Yag0ULHItCO01jnTpKKi7lIRxj1l1Wi
CUFH2tWcd9pgqolxLjgx4dkMBVFse2dG+gYyy234KfdNFUkomyDf73b3C0V/
vM/nz6ndxyXB0PeEDXIdbUtUhr7ljf/0r/LVF19zoLx/VBa9LEmfzVx2blYk
2WS/s/pn/1v1MNQX+xS/bT/E6ePFTrRdMT7qfRIZGxvqzV9JvXA6qaw9kv8T
ytJ+vYDxypzbkCb+oziQd/WnfdcZfwvfbYFIjZnvu+mpbss9XxZTOM9s4RUK
GE7IaEyU6pQrmKTcPGM2dmKq2f00V3C+7S9rBpYbi1ftlBoU87v7M9fkwzeA
Ubt/gQjVvcKT4UvHrkG8gyVqPyhNaISKWb9fmR54WeIqazWbVU9y9AQkEfG9
I96OovhATiscbvfDKAqjjm3g+cBGvLJe16n1krMZ3Ft1G6+3zU6Sc+JOq84w
VrHuxe3/0n+PdHd9mKP4Eo4++s8Mz8KlU8rColG61Sgbkv6qQKn2/AQAU4Ha
QO9BgSX105UhzIkV7AVnpkp6uWy9yoFfJoEMlwCWmDzEaAZ1gl9bIu82f+gk
Q9zS+mVuOBw+DhW3sSuyQZYS66tg9/4p80JZdquH/AhGvPXIK8spin11MVsZ
BNwXav8rsSAxrzxGSwS+BgMzXdi02MfBWwK8Da64iPnJJH+yIPSoxDhbzptM
r/yquFR0R1VL6KFA8P36wJZnGtv2rsM2oHMpYgFqOCfwzb5mnOIsDx9A+nZy
qxlK3w/5Jf5SzuvrLq8wToez9xpTeOhUc/PE7FOwuBZQ0Swwlb+5JEp/pupC
gpNM3iDR0ilj29i6Tx7SK3EmFWLMHSBBCWzV/+6ryv0LBWjMaINv6BuB0Fqs
aRobf7A+iiXP5Ti2arQFsZ1hLbWKfRHoEKrFaYN/Q0WHK7U974lOfDWi47Mp
18LvBFE9AZBALtwVvSZMijRsFRzdZRZfYWwWuomQcjOgS4eKvN8Lj5bWRYRm
EY6q34LB/Srg7riA0bmoBbZPTMJsS0ER8SBgrlpL+7iThFoWLEHJxO8TIwHi
7ayVTe4hQQrOD/iHcwzjvbTT5Rej7wXGvN7EkFhRRmX2pIoca/VS6SBg31WR
v83lDAtp5p+JnaujU9ZqYfn1CR8QEoLgav1+cUgDkz7udEhOHwuv1zHFpFIz
3HQbJFsWN2RCk9XpuGjA3vk+3E8ELSh/GUpsp83bNGELzoIIO/dKv6Me7eVd
jlEFEIaxahOl/FvnrcewBdfDAbStOUPi/pnWV+WcQYQDSzzYtRTL6MuClztp
JcEp5rozsbwWTj4YXLr9pNsxLth9+aMyrRIzkp+pFm/vjrM/39/CJyJ65P5l
LyPBhx4cL4O9zq0y/p58M+NaKgyVSz+C0c5JMgGQJhWU4biC0xNLU+Aq+mXd
RS3/9y7EVBsVYUluLJ6PXrP5Bhs6KZ8jDwyDAMh0D34zJErvSk0//BYqT6KB
ewdLr2ojyqLRFFC0tsK8EhyIh72qSWRNNGGrCXFixku6d6I2ZLS4Xa72t9iS
Zs9U2zxS7iqmbvpPleimd6DBw/6t+1s1KoNcbriPHgsKvNJIqFCNs/24Q4FW
SZ/P5hEN7frzF0S4lnteTIrdIPgyEeMrfjVUdGRfV1xVm+8XKNWu3ijVkJZ0
diQiDdLPcQ3b0vq5SjyQBI6HJWwNsV8xstahPwIuo5uEIvAZpisACRBYNnN9
fCmBE3o1A1TLXWYUXQI+GrRZKU5MYtJzbg9wm2/z2H7t/5wbY+nVabHU2kL9
t+NY/2dWBywJTpeQDpeKvlBF0Y8UFh5M5/ME4jnLGt5ghKulugmYijGiL1rt
LlJkGqRQH7mtYr4XYnKx6TNYB5NwCCsWGAavI6lmwPxjgrS30hkgh55wEk/L
Eo8hDMVBsHOH7VgFpRGL0yQL+lRepLu0nFqDK2lHhpGLwFUI+rpcPC025jwW
hzm15LIdyJZ15HFKd3ANCm3qE134W2Qv8lPZiHWmjy4fX2+9MbcgpB6iJMgd
/XrxLJzUyxy58Et1jdQLqLHidAabUL+fLn8VrLA3E9wuKPfkoKzIcVQkmRY3
XmqtCr4+JWCcKeLd/Gv+5Q0IPXLfLXjDQfEa5FauEYOTKNPTJn82a6ZU1s+7
Wt8D4shmbBsaZ6Kd99iMmlObYkii1Zww0ceDNwuVFrrE2EL/fVb2i4m62bCN
DGnYi1D5TUykP31bueUZ7xx2zBndF7bYh0bpLsKJwUI2iGqUGxC72vwRK2ZP
WZhWk1dcuD/8tPvFqPcNYVe7pKpUYhXj5SyKU4vtN0j/PFCZA6ZjmtlTzDSw
G3SLgzJfpP6T79DWZje+vGW+pB3OXny005HnOfQv6A03M/mv7vyw2NXSYxpM
Ki7Trh8UT6mTwTDpT7JRNBt9ByH5syDtCFsyarmsWFWBDB4BrX7OI74ESOt1
6KSsQtyvctis2EJYgEYfLk1OFU+3i9YfYRCCu3/+jXpuEMuXwhMMjFI+bXx1
jaBeUt5oOOMR3Wxjl3D8LFPjm2sjt4wJcClEyJtR2viVbioVrhjAAVY534xY
iIJ6mBlkBr0rip6WuBw1aaCaj375HqhAkyayHCTOmGTglJ0JasuHMWSMy4Ct
Y2p03TcseDE2MvbbDLr5ttMFGscZ0b4St9b0Dkj6+tje7wVsqWESWoAlwDkj
0dEpcxxGjzoK0/oHgF2QDzvx6GWyJtRPZJKYypfLASRHdAkKev40sO7fiSr/
w8zR5YR+5BbEZmPUOW+K8DEBhRt75tS+E1tnqwLmcKw37KYor2aC2A25xvkj
XW0SXvpen2qCG8yyCdUtIKoZ3nEmeQmnuH24uABqIQ0CHn7ahzbsSpezYIhb
XfpUAqmX7YiO3cjgbfHblrnhZjbjsI+ccoyUTT753chHLfEwNsj2RCIeuTQG
TbTudNapMQdoDEcI2uykM0i6yUvdfDp+HNDTfPMA62FfP0BIpT3H/nA4M4Ta
GNu1ilFTcRVm+DXNnH7t/jQV81JoC5FNTbNaEhutfqXlH6qL0QhJSmptDA+2
oOV3+Ack2+XkUh9xLb+ePtaeIhUhYwabQcDdv12/skwKE1T9laBy5eiTv73J
3fg2+goy+BhdpCpEGzzOrMZg62sQNtG05jCyTalbx4i/buNZY2qbPEmZ630I
huVt2xK5iIaQ1/1akhhlXykwPwI6GbiPl/DdMBTgnOD/hyRa4mybG4spId+o
ngi4Ddp8FhLVX3SQCnnoIyJ736sOwo2XxaPzDUseW/X/ROL0+j7wSCByqRHo
4b6mTknrlX9op0XdnwilvnnIMf5EZ47K80O6LlGkQYylXz+NdfMXHq0QBJgF
jo9H6EzdFnG8UDY7WYtxJrEXLInrkjoNkN/LSmPDPkm2BtI5b2qhiMKx0JAf
oAEddjDd0REj0PM/GhJxgS3/oIwREmVHqUPnUih2fU58wlJjCoJoFULzSIvO
vJqZd93l2W39gdS5pxaNykW8l54g2vkZCp8Yq1YyzTNmX1VSY2UMA96USrFo
HWH6GXshxgJZtvPoWQCBTCCKS+12dgitLnLxqkr6Qq2jzL++OQSh/FYYa92B
5rA5P+9lB2n17m7guVuhtV1ckODVTlE+tVVBA+cs+QhjCWt6Y8FTuPDqZZ9n
WtN0BKOFqK5sjPLyZWeY3hdi/itiURqrOnIfJlX5Im11SDNcem6nbxQU8/D5
laKz5lbO6Rbum5Yz/kl9W4nv/f2piK0XI4zIddyYOSpCoBzy/a9n+4g7ikYn
NSz769wUSdbkxMMGn5l0TtzYuUmuWHa8bCQv+ebCdl5+xRrU8Qa025VTsMJR
fbRRh6NoHK3c3Ykd94tUWIyqFLhjngZyDXHDW+prLiMOKs2Qm7B56gxmCVCV
dG35a+A0zMo/hDU/jOy/WPqPBBdZK8ZHRWM5/NR0fZ2XtnscQP9NuZUQLJMi
65RoB2NT2m/bAfOjwlGsgPu9L7NL+VD/UFKAJFWHzDDOFEVn3Tg1etxnf40c
7/sI7Ih0jypfOb13d3GDitqGZzKqTn5wXG9tM2V4ra8/48xGIEHjtQigR1DQ
8UVKt7Kd2OXMzcHwmyFeGAeoengQEF9DiTAaEB3UhODiAI9WNAlPpbOMM3Od
8/ZC+ykI8tX2pxp46tk13Rc+beg7kFHeMK2OpHfr//g6d4ra5aG6CY5JqFRY
Y8/TvmJggajBjq1R8G1K5p9EDOTPdmLlsTBtUDADunCRC1piLjtUduCvvXwT
UIEpgVm+Z4kQ12rpT+F53ftVSwzdNWIZpA3xKA7B3v8lD87S/2ztGibar/Tp
VLMrpcb68pmZZOsPB0uNeg0VyPKwOelNsCf2qHxhElaOLBrpfpPbpv2CeWjA
+EIzOA05QsxT9ChNkHBHfAfyWBpwfqKZVAXgy2UA7XhrEKwZLdKUYfg18Wc/
RozfbFPiGycDMQ8r4CEaD3GHcJ2nRk61SJ/J46AvRBDBA7VSx16ar6Lm+Pqr
E3ikBvxNraPYNvEGjkcb1NLN2kf7LTnBq6R/pLAC19hcU0JC/3Klmj1ALfuE
nM5KaTPtTDLuT5E4hQLKNE4p9dDdztjxgJHhlNE6Zmdv1canVnxYpuFQlIDW
DEuZTpuoTpna9zZhW7HK3sswvO+Rzk5RuTZPFU9ydGgatQrPDR//QeURO5Sf
9DiVFfbJ1OM0UHlnHi1ZdJT+H664Vg8ojimDLAha/rKDZhKM0IMG1TcVUMtA
/5IX8rTjPhBDbdYrwGSYokqQFw3ZJMPccG6wy5NIxHFy+x2oWui1hGsIkZrj
ZwPilvQKI9386EsaGI//T0HbVZ78QgA0nCb20ExdFEnlH4SWxU6EbVZ2jpEi
4LA20WXnkt3IdFXaoiVw6lHAL37OgOXi148eZLH0jzZBLgHYYoPKYP05tAsX
+iJksfMTJRJ4CD4BMYOaYEwwKnkraG9AFV+RufOMSiZBtoKlV9BbodcXSGrs
U0WNTm9GIkGe1LRWEc8y/g9J4TVA2x4nqjvdh5UdD1VXXn0Wcva+UXQAB0M6
/gb7I/ONPMD+1p+pTTLAd/uPYc8lJ2/YBEgQNPCRzSgJbOgB/WczJc7Ds7XW
yY/uLMejNhDTmaaNLcDtUN8Mjb8huPtipwU49gRFixz97vJUQpjF9lui9v3f
J4FDap3XD0J/0c/6bCU+JNLJxagYERrFXOlH21m9dmQHyl9VpzkOldl9c4Z9
x51KrBGQhFDB0jA4nl05NLJO7+XmscQWQIrFc5/Cvmdoogy1CmQ8cPD4YEG6
5GjIkfDKHo56K+hp07s2gI0VR3cKnzy0F/CS2IjGw0bO2EzYlInLGszK7E8H
lwDKHuWd5FpfCrgi+jJvgDCTIDCjKfgmeTks7ariO5+AdMk/1uBImtbb8gPf
IG+2Om6iR45SGm7Dp1pvfIGw5UdJOgayjyhBl1XV96mjniKVSd4/Fc6rpOni
1uuh5hD4lqA5ga6x+kdJL7uWH6vzBuA9bbwm/5e/CALd491Q7RISTo0GEewi
h97O9t/ZEP+hLmDbY5hfXlr04H4xdLLVi/of+J32agh61MdlgPn8m+EQ13pW
GI2a7Y0nWZonLOZMSlzqzzsOQEaQS8tY9uTn5MGiDkxxiiJQldNtSpDAMsYf
Lwm0BuaF1Jc41yu6jsnmvPO2RiMzTubTmtutXFj5QO9atm1ndYMevJojvWzI
ddxcp21RXmkUuOU8JSuXbjU4adIUoq7jfwFQ0Y6WTAfugfBkQWb+3W33w5YS
x/cVetYCSJ0qFJJZ7phO11AxTrXLfMd4q7j86hkbghzUHTKLzKgHCjR1SJTY
3YIhcRMGLugZC+FjffIFQi1SF6ztEHnbkMZvCF2UFZSmpOk2PKwhnAflZugV
n9SlFPD4Z7wxD++5L3y82tkShdPTIsnTXQDNQXQhyr0n6/T/mIxchwsO6HHd
ZfyNLGM24Eg/25vEOd0I2zOwykwjuG/w2Wt5O7gg5YrxdVjDa/hULdilaqa9
JR0ethh3j9UtIOVtFj64TiSNP/llPcSxl5BTQNlQpdooKnT107tcleIZG+Ww
JuhaOta+74VpxhEW97/pTQVDf5o0vnXQkobZoC7hZgm/8ijpT0TWer/zQmck
XV2ReT5HVnacxLtu4gX6iCEjWi/112eHZxnxWsbjim5pOGxm/kxTYuqSSidX
QmY3D6WhXRvAqDvkrsF7iJQ+DO2/zrTus1sDW7OjYbLxgzSlZWd7CiZaRFgZ
WD11XKKrRwb8spQCxou1ygwWEH5+LX+t9zRO9Z9n8HXpHAAuShGDAXtP8cLa
lLOL4JV3Ke8yBxSORRR8Rtd2oXL7T1NOJQsMw1jixwhpkLQJy5MQLI2liOjg
HjQSWdZ+qFtuJ33SnZDS/Z6+Rt9yPTAFudL4VeEiezVzz5t/MhNJLNrdZCkv
ppDpQJ6wsRWtpLs6W2jOh+SQgbhpz/0v4VB98JsPHDLvSrSyXWxyeIu4LcHI
DvipO5Hw1KVhW5lO6SBgIX4X7XkVs/SptPe+TLsothHZj1kB+E6R7VS9thJl
d5WXDtVeFpZtUrN8Q+FZjwOHsAN0AuY92G/tBrqSo5Jkab8e+umj8vURzQ4p
BnhNH2cNoJeXnm+aEyTOrL+v1Lnfg0rtw2R/cLiIp92BjR42TcMPJFsa8M8c
v5JqchvqA8xTMrlxcKLemYXNxccUUEkY1ppxYXxZ4wpEQ5lrc6G/+AS77i6B
8mUK+PTji4gDplRPN/Nr47SNFmwZk0S1kc6RLBp3mt4uBCmam83JN73pwNpd
rTjP95fWaJJ2nJZ0KwLX8RI+JVP4wTOr9IVtHPUeUMNMJBwk9/fzplA6Og+7
Lypln9KurqVuNYxDr6/qp80ONQsTNLFNCMjSSK+2xbhbWpec4ll6leo5J5uo
swABGJoT42Ntu+/LhTdxRWa3JAmR8InH9FeP+w+qFt7ctn7Q/3/NZ3hjr987
Kr06qBwH95yKR1knUCuiWTrvpeb6vujVsYjkPTvgKchVR6YDOjfusnRqrRe2
OvyWbTCB0YR+yPUGWnyE1tYnBRDwEP/4f2tiMiUtybgbrYx7vJdbBcDz7Nkl
2MbA96xikyXrfaey+OkaDqUl465cofHlhvYNcyfWTejRjcu+P2pLi1yCKLGN
XDEWYHeMQ+pbfZ6Us9wH5LhturRr8zWXl5yeTn4yzhPIc0aPgDTOWQqKvxG5
LNzwnHQxd9o4dPNLb2y6JshZEgrqQBWOghLIk2FO1QAx0chRQ5Y5+Ugg7jUL
IIvyy1lhuDvF7WKmibDr22iubkqE+X/kI+G9AqTSEceopGjYrUl9BqRnedUn
sAoxIOtRSTUKnmu3ojnar7kHeA6XA7yaxXoJpWLloEb4nHYSCmwWyImoCJqY
CK7eF1wakQTNGmsOKrvk42Gnk7iM/z+kmEL/rK2lVyVGEgBpKz7K3FcQHAk0
1BmElJetfpOevYiIxq01oPqBEHRes/frQeW/fMBGQ/Y1H7PBeDNdlbTZTBCt
2iQXDqmBHwHS95FKb+blGPe6UxULdUBrUW15xxqcuX408lYxJnY5irnXiNTn
UDSr5IFserwGixrW75LkpKFx9VbnivSihqvNpW/AjH1qv3yuScUQIMffcZSW
ruF5L8PpUCJeqEfndCdXqcheiw4szRFxfLHxU+wpSR/orSp5K7SdL/mcCAxN
PxWOTK2sH+y7S2pjD8NwiaxhiPYfb8rloZUlNwdGu5v3+jXA+SM5xs2veunu
UEaYdg97f+jxxrA2GAkskRbdb2dtzjlhPTwRVUBPwh9JoohdBp4vsEu7Ztlm
0vBFxF5q9Wc94jk1woBa+cb3qg6SYrgqRkstD2BN3TcWHVDXlxwJeL/J/gO6
DwLZSjuPi5gkGV1WJaZnYr/BMJj3UPPq/5hB9DjwOVJxae38tgwaLKRt3S+5
P24UoYk7di5PUPrVFdDpYMrP29NhlwJ61A4scxFFkxyRvLQxOXkxbUtjB0mV
hOmt4S/8PwFf3xiy50uzP2dVDEUijdc/mBF+gL3EeRBWTujL4qEWgAzxJnkJ
FkV39dEDtLvKwjqm0QZrTE2N5erbvJlTP21wpHa0rhSc97+GyX3MPLCAREoE
vjTrQ2cSecn7+64GIOJf0TLN+MboHw5boNdb7no0QIsnJc5C4YEsLadjw5Jt
0HDHHRmIutAAgdl3JZEqYr0hE4JxHQWSJfvVdN6H4NiBs/QRlLNoW814GsU+
tiBGNh6mZqfsUuRNxatm3oSwGM5nQbPdixcSOESrAXKduo4hd3drURmngfdw
c+s+Z9DpaU/6ZaJZF41wUdw2feImcjMtB7Z1+er/ULK0xxdqC+AYMbhJwllh
K0ztFIRSIBeOxsHVe7Ct95RUh+qfLCBb2bjo5T24R8CNJVC8Zm2/4tYrOc9y
WRYBZUw984Mjx5TWKXUW+KLkxJ/a7quB+w8YZrdkdZmUjaZ49QcDo1mDjp1e
l4gbtcqnJ0hJJ3MbSb4l3YxzaLHQAXRrlWOElJx3x2NjIB+zFXdFs5jRtdAT
YHKRVtVFtl7UjZ9OrEGwlNZ0gXjqVb6M8zSG4tGrqUtkGqbSa3qI0MI9cD9q
0B+95a9/t9v9BBn3RHmU1oNimeV6R1NR5RZcD6V9aSK+B/uQHCod4XvewSK0
SgJfSATfjEYjfWeMCpGT9TsxEVG6q0QEYQ+ChcbnC5qehMayPe7/OY+/M3xh
BGT74obPeZZHegWKV5yybsP2Gza2BCj7Ief5Ex1owG8g9Jndlc8IJaP6fzgI
EC0FZDoXesLT8/+KxNvJ9HCnkjAaMejvRW3ypaEUigFgS8qfbU3wcriTgc1f
5wGTtCEyBuh+cYlZ9HEQn8efseiTc0OTNK/di+M4R+9Pk/gcPlcuj75/xc6r
OZpJaskc2ThR+4bwwxJV7ud9HPKG9RCRgTh3dKVgTcsYyCQAlUraF+XdUTfy
KcdGpdxHwAy3+eQyChqOBDf+22YPNZIMvElBF+95O/6XUKR6F9Pl0jW2/z3S
ni+v/ygaMFqcWHBa4sIbrnavnPmDO+8jKy8+DswyOGZaLrZkuaBf/wG8lWny
N7G6yiz2g9ji7lic7xcNflQmc1XhAOmW/0mzEb19raDQNc0oEVKORxQ3x5x8
FuUHPwpnVxa85ifSUk/p+g3gQaQ0c2nIQMQa9/0W7tKKP1rMXDKOfSRFt7DD
lXioUbnQRubITK6huA57GnV29At5NXK5vWZhuGCRWDjb+bF40KHDeQQU2KnO
6IsZRTrVA3F2UWR2d/uKh5Lqxf5x+pOcHUagzDuccWVU6W6+UxJ1Orwy2Pt+
WDJdLujA3Jd5Mf7z3dbJYTBihjtAxcRwVRIa++iMZuTYVF1UtDzuMqxJp2hj
p/X5RunBcsoJj56ZC+OQl6B6BtBV5GZK0b/VoSQ42f0d9AsTiTfHtFKa1m15
z8HQflM8sxJ9mjZP0EWMUnfWKxw8zywTv10YCv6tNARbPF7EXk9BDG/PsKwT
+Spsd9YvNb+8ehZR/c9yHwdbBZsvoC1w2N3TwVpyEnftD7PNWQ00anSB62Jg
MVWmGgd5TRU41VCaeOwQ4Ssu38IUu1kmtnEzxVkpKZwVUfs1u2I0trvR3gea
yb6UwsYE1ptxBilnF4TjyQ4iqIFHbkTg72A0N3C7FwtLU39v3oWWXxNcCIc3
ZtZ1Zf3oatkJVA8UpRlVfUhgxU5WYksGKJfcJxF+FSHrPJNzUAL+q1Q0yNce
kEOe+QYTif12LA0ltca8vEWJTbauC9eo3IYRc6phbqI3KGvxucvD6/DlrX9m
hkITl6lRWsFnBr6SmRU8W8r0uXBPTr7u8wfEJPLklZ1eRcWJk345kfjawkKd
/UAh5fUrOPzpDUmcPueuMTCvlC0vmTtgBF2bHvCshyChCymR4lcpvomjvWOR
NIqhaaI9hPQQHdu+ipPujf5YLpqKBYfY0ozUW16mpmtYrO1XJVACF8KRT+1C
rKBfU/7cU3GTA5/NG8Mt4kGSS4e8Sf3+WyoiNwWIP9K5s4NkgkRK5R5ZYiJI
mW4Z2TvTdRR5remQ0oBzQzGbzp0RxOKFTBjhHdqaI9iNh4Dg3kQq+xQMCQK5
Q6qFusiAn5QYaTvMX2OsoX3IGGnhWUk9z9lsHZp/VdMru6zLzw5xfQW62l5W
PoSDIwcQ7gnCl1exCg3FNzBlUujF56U8c0sHCM6k4PZtQah98rLu3SjfCxvi
/nDJPOKlEMAt0Q4kUsLawRUqdQrZL/xzabaCca3Lg4as9M/He3A3oOS/+voo
kOkz12t4g1AI1Jjq6cr0U83IE9eBz/eckFhMS03KBO8JtZ6h/N78dcy0gaOL
750dTdryyXEwZ6rBb8txfkHaQio8+n6Anq6wLA50mDOwbtKPKQGZ7YjZ+SuP
VWkRGLwGZOx6SXKcZ9G6T1xZYtre9TW0WZhJ1Cs5DErzB8ClU1FzyC/eomuY
ZpdAhRjl1VwixzlmdDBMxUv1i30bnj6ztQM8LJrPBP4mJRmbvJOPqBKcJbUI
Y3uRU2aiSkijvgwe8vgxJYmXjHilrSHCVVQkixLf3bz4qLmuzcj3XQIYnmfD
T5wjFzUWdc+9LZ/osNsW2UsVJRWN/H3Jka8Kv7zbEsISNx8gvNw+7sqDi8ON
Y8G5PJI5intc8TTN+RTtdA45s9CW8X7bolZRoRQHQDE63QWZaFxbPIiZl7CH
u11JsQct9u5/XvYd/VIKBjicxMIHeahYXhDGGhj9D+m12KRrKBdyZk7OrDMp
+YdRDIvPHAyI1q3HBNMGvpEYaA130T3kYIMz9HLuuQHUY92j4ClZ2ZXZ17Nq
EKhyj8NnNyGZ8V9QfHfIYaBGu7IEnDub6Sp/qvBnnhlxFqhpT7JChXalrZCi
OweV1i4DP7vMZNgD4DkvpeDYwwAm9OBLsohdwrYEu9tzsIW3hibJYumN9AiS
Tly24TE4jTXNEdBaSY+yHzCqwZrYH+ybTn7RT0Z/jn4vIn8pSblGvITd7QIG
OKyvSzj2TTn4svjIjQWHBaxp1xiqRCu96zgncEHVFsQ1ijshy/B/ITOfhJhy
NgFUu93KGBvwZ5SjYy8F4wELmtrQvKhi6GRMRrHF27WgpJCBn7RgYPzLUEX/
YEttZwVyakWftGJ291rjIqhhFKpRj7MdXTfgORIc/irNlAx6Y6j6sh75T6et
EmNvxXOykYn3ix2LIkJVULG0PaM6/eoyvvA7OjWIEgJ2CJhO9qY4bzFv0/4m
fZS7glPCVjJI/it7FKnHPYnDjnw5VSmX+fggMygXgBFcA7//4OHCTeGMTdhT
fbz+G0bcKH1SxlZmP+mMKeNbqoWNWeuxTR/+udaHLeMqJQm/K/aIo6X00APq
uEd9q2Dwy6syH8d2LNTG1+4KmwWzEaQQyyoEfZw5Bb6AG0w3zFv62sOQBzwP
NTIMMt8pPSwCVhv1WxEb8zDnbw7NdjIXiNL8QPWVPR1+1k5n9/BVauqP8rEM
eiaTTEQ0OIzgKSbsh6GYjNCQB/KEg3XEGrOHONAMj1WIuS4cMOYPFcsnfEGv
7rejrKVhugV7EqqKAgXcbSqc3x460/vAVNBVQdNL8YND56pZk2oLBvr6GtbN
Aqw49k+EALA5oLl5xPh4xNYPN9gvYJLdlYn2lVImhLhtd36HCTxQAiBAmI43
gwYpLcGlbLJW3hna5pk27HZjrygy6oW+aZfmqmYeR/uhMPnv/UCFNwHKzs6h
mDTO+Ll0e+rFziZSlf8WvxiMRDckEktI63ZqG8im3RDs5qks5OjVSkVmp1wZ
XcDl8M+pMpDXDzOm3XY/toTBq5jRMStWFFmN3xDd2fbAyguEjwRoVOq3gpEH
iM+koHirVophc2KZM/ODECum1u1s4AuMFxzYh2D3EvmWjzB7vIL02Kk5XixU
HI39elXIp73l4tuQvsTxeu3iMVUg2f+uAnrKqHFATybCRJxL4MnmjTxeNFLl
PUrVFCvAATKRUeR+m5WnVPEEbh9x75i8xyMkJINJwDLn1KdQHoj2l9cEJNo7
VTQOCBWMzSI2iLJHZ4mmAhlovO4h2p2sWZTB9A1SIRCcG2rdJIoUBgxLuL1I
Vse5Fa6EggHJbjlVOn3h4ta05SxhHAiWOBT9yfEP+88N2yuY9n3B/wIoBta6
tf+eyXvbX/1OWFRxsMVTanFtWLaW3sTK0Vy2HxNOzD2BiNi9EGkN654knM1X
CrjQ3MTvXDD9fxrWNa5hzcaFJ4NetzbU49e/nYADbrNlAGarm4phzDf7iY2Y
8kMuDBf0l93V7CmAUZ0yyLVCTpRYhSkLNzCVa49Yv7geKuLmoob7dWYRUTri
3iIul86HrRuhcWPqzBgz+1zEsy0bcNc4H30mwYz+6s1ufcs7Vf7XAxlzumSM
bQuEShXDBInSGEMF8tQjEHZAAomJpPuqEU3Y4/Oe27OyYB9n3m6hH3NFo1et
uDSxQFQIl2nICDKqwoDKIwmZgEJZsbvhIXv0xuKrKIdeakUxUmSPsdhwIGET
SomHQU2zTUr2Ut864xZBjfwkAwSXrpVbDNyPTUNp8QU2f/AmpQ5kvtc+epZ5
K6aVwxgrUctyZ2DQ+o671DGTA4RI+odtTKxsn+4S55Ns/1cMNPch2BwJ8vUt
HUwqNHNj+jXhfY0aaETvOY9gCd2HugWUmkEmRs/B7bTi6K/P/bxj19RNM5hk
qNb/LCOei62NEVqUnXTEmjkIU2qiLMwg2xtqYHhmneZXNnNAVy6WttYhc/du
QQE2KJmerVyZp8s/aI52d+iMoz11seYQYvD/yOVNR1WO0Dyxp/sakvvjBsJe
JmHQsykNmjR9XrzMA6M/Q+Jcj4+I0K1Z9FflTf2MHrOEEIiEW0H2GERK1Ujs
c8bR0FSgGp9wQ12XoE53w6i01G6T2ajmeLivNOGJFaT4MS8JpspvhsSh2cto
1YHehgWEY+oh0nLIptzPiNqUekMlKwM+uvrwgfEnJp+MjygOc0LGwc08aaVK
OMrMw0HCVti8CMSUr7Ib5IakirCZDkPpj+A2npYfI+2qalw6IXiOaMkLBDe6
QHm5coOSUUYI4Cg8Mvkb/ojuWnFsRGuhu9o9/Kc+/WiGNKacA6hT1fVlcaXt
X+uF7M4fV5F9TCB5NINs4pbdSrNb6RzyC8qtu3V+EWPfQxl1PySlNCPVP4pu
0jawv05LKyQJ00dBH4kZLJF5a9PnKK5BdpEwY1Ci/OnnVi1zuH11rM0QZJVT
ndom8n3PJXAYdpieRrJzdKdApwMnfi4d/yBIqcNgBOzDivmv8IfI5AyOIBlA
afuny83EjyMcsmXsfyR6/KE3u+eHy4g6Dadvw9327XDiszWhTJs19kjJONWp
wK0rjcaKOlEnaOUAXcIB4yll0YWJz6oPG9s5u96FcCYIlxNYm+aKST2ZdVhI
MsH45SFW4iiqotCmZcjtkIa0XBRsgFtlUIzJIPWYQfGuR4xlrc5g4Q4aYlBx
hqI6a0iIPO0VSsp580+5BcyJI6NWZCbAOWlvBOu3AYeM0kLL/zjAhOb45gh8
j8+DWR1X07y8K+yY5/DTwoavJOcK7U76whJ8tEc3M++Bt8ykwzxNsXxC9JWv
etkQS58TibJ54XkqoXkz7pih85djjQilNwFz9KuaQGU4VzO9xrIYGEipP2e8
6CVDmV1qqN1bJeI9hfpvSwulIEMp8IGxFSnFTSTlDyGsf9XZit5uq6L/oIfO
G6ijeNIKHFosifzGXDOz6mNZ35NvHRc2j8ACxe6YCzoT2Lf3B5zl7g68jgoQ
t7ElfTy16yQqIxhsumHrCfoRqTmSJPofM/B+S1doyBr8X5JuR0fdomzJsBPK
9OSp0JMOH/slT+PAsOYvCZWhfxrKTs2KBoFFr9k9FWIvx2jOBKwnzmBskBN/
j3SWH1R2Lj0ZqnA9jzhv3Ms3OgRNOKoAHRpKuGqXSfkhqzhy+WtlKf5PeeKS
5OQxEIQW1fwMNH6vjQOpsXFQ3C48S3sfCUj5FLDMlTcEh6EHfeG6LuT9dUMU
4Uh0WG9+hp3C8ok3lqTDAZpEXQSm/Dl3MP0odlr9ZGq0qZHaS7yDvjYk/gnr
yREpb2twc0tnP2WhNZ24ShFFxHT9OnQ50wgzX1MGv85ZLl069OW8ZLUSXYGo
bJX7ZEe667dlFuQNQ5VrMpSghrgLGHQsngAyj4aCTSFgnu+K1FyvhXqs4ntg
XHCJf50MI58XHfi6Osd0yHQW68UIaKQtKxJ5Op4DqPJHuxjrjN1JKgZf53YC
otVrfJBHHzATnczQ9IR62UTJH2ktgZP3IWANP2qJB0Nbyl9zsa275k5O4hBF
Tr89sW1cJfxKRiHLl/9K91OV0yLQnxPLjYEwKekfGicIF27ZoPhYi4KzApF5
nw//x8GsWRFKevQnTQHDS6r7AMr3D68v1gPZYBRu8keFByyg5CdrhoDAt9kX
uZembfOpMlCzdzzQ4efqUst+2U7dFImXpU+Bll3TArWdcloPV0WszN+iZYiJ
xIyUU3Z35tH7FlnRnNuyDDg1vwqUlZvD7SbkUM+TO5Gi8afHvlPXWwKuFyk3
jb/g+Uyue+OINNNqzl5R+hsSnT5COPp7NowEdBPqDmr0x12atQ8pYk2V1HCB
0V5/NnlzNhIwxh6wMJhoi34YpqFnxHMxqY+4Xa73oIqrlPyD0rPgJCbMPNOq
M0iZFPeV8x2cfFlC+BSNJgY7evtnwqRHjkcHSjT8OPTnuOM6eSkk5652kXr7
ZiRl5UPzrSo89lhudRCDsivvKDaiWBm0bm5HSFrkspBfVMIFdwnEATdOiOJj
lXmOXAr6wopoeSCjyvR0pZtcfF3NEwg7hVyj+tTh+prGTHwoGGir7vqNunuO
LBGflIkyLxIa10/SLWF5rZbwjffSJiIh8Z5c6n1yiMLc42VTeMh378RtV1Ax
LP3n6CfJSRiOYieQS7X4fAikSNNeHOWh9U2Lg3qQ7XMsXR+nzObL3S7hbNJ7
+7VhYZfZMr976X1rhVK57ifOD3VUo7lKFr4yrvemukNW0m7SJO4LNTarbILT
9EhIKn6ZCJXTA+9UTBCMlgJjb0cVtZWuUP3eqtPw9ddh8jxbew5+/8xt+qUh
G85rkJEc/lEmq5UfmxfpcQ/3z7q0E4Yz8zpjcKH9rmuwXpb5db6j/lXqwyE4
RvdzC3kWR8QAAJapHbOWEwa9Y4WU2TTfOhDSnoZ7nFehW69ItlqAx8W+QnvM
tSN0T/S4LQRItTu565uQUD/5Kua4E6c6m/BvYERhSKrhdWu41rQ64w7Xe6Ew
AL1diMs6sXUHtXqqMN37PMnSiKgbuOAOjEszfHqaKN0FYMSCuDQjSnxjvjee
/2/sCVSbn/6JR7CIbl66rRCk/JqGvaU5tY3SrZYaQK3sa7ENijKDTII5Ef5o
q+XtC/2ZMcPYwNg3SvHt1WXvaRH0nMLcyBCVa2uwUNQ/KjUtRuaMs5egsgle
jK9P1S0M+wcPxjf34anMFwZ38gFT9VcOeYvYwWV68VLyAjm/3wnxHZYmse6o
eE3uFquiVFSqJqyytQAnPKuS6ML8ewg34/h3n0jkT28rhTilU+1x3J5eqhD5
yC3Ew6Ta9GyUCltfQ22P+yfdzU9wQksifTC2KYBSL8wCF31D3vzIqrUHzomD
mQIyjyaVwblk4HHcpvCzJ90T3PphxY0HEH1FwKJuKQT6GVF9HjpXbHB+TqiQ
BSoF07O2j5Z+uDae49jQctZLzTqY0Mf85HKhbYQKIi7ysyHXyB2Nvr18Ny8L
ull9mex/09HPTp4QZDUiZFshU73ofYKqQ8qCy2dnT2nWXnvlXBu31ZkC8VwG
n2i0junCzr0LOzWdeuZM0pyjolwidhyGiP4SRYWOgH40toq4pcceHO1EjbF2
6hsZ7kO1gkm62yIm2jO3wYyedkYd7F1TeByzv8WJHr0nQ5X5llMhLS5nAoqe
3oiDfyUohc4anw0supjyvPbYhMlS2uvf4GapCqBKOp9IM4qOmqJEcORbe0xr
19jai0NzBJhifK4FUKkFbwFw/ZjbwJjxwdWhyEETekbMibdmCcm8fMO9SN90
cHjY4clAjRJ4BB0iGCMR7sA0TziTq1+UHNBugGA8OFM+w1SSaW5xJV7fySrS
P5AXf90JY+EztlBQTvCulx0J4winklxdog4nicv6ODukgHkBkr8P2CgmMmup
nUW/13Ke7G/HMewHamsQlBo0m/wn//HVYxOxn90wRD+EKExRgL7tLSuR7ZgO
l+Zax3ymtc/BlZAakqTPP3neFTg7l2Me9lGXMRQ2dMNKd4VRYkLHdA53BxGV
7tdtLXv45aBrprL8PwK3aylHpTUiQVwnqeShHY849JzGiGa8uFAWIqfvbgme
FBeoE9hg+M91NyaAjG1i9s9xGN2GGR+iVc/SUsbPl1jIxeEffG5dIcHY9wAY
QjQ6Ui9HHrBgBbhLHOIFIndTGJ5kNt5j2K2qjJJb1iUlwRIyM5bujHDQaP35
lDyWYwuy3XRRvrvGhdIsletnb+YGTn3Itv/AlYQDYChdny4y45rIX6NVsjYN
prQ6PVag4eT5hNXwa58VBjtdT+8jRIguIsHwn009j1Aw1mOrFYhAHdTEMEmT
cs67V53hhZFUGCcyFXMDF0W1NernYSXdVKHICwyFkycBFD4n1AzluWFsCmp3
VzKyLELdyj7zI2BKEHyQ6SXo1Dsx+hcEGs4cpOaYikcAkVc433frJVLFWyhw
qaa0DdxF6Rr+qLDiHM7Upmy4dfK1u8LLZ4WQMTCmPmCuSmmjvnh8gUmVxKEX
XmdSnGSWcrj5Shiun+E5wL429W/9JmalKkZazqZlzj8rDVgk2mNHgvJm9Kbx
wDAhqRSCil1rGYNEESX9FPRVCb75kW6RpdMQ5z3DjIRgTwCjdXd6FKlLRCEP
mBpmTD1GlAtWKDPlspPUY21xzMr70R9e1m+StGCB7ilD5NYzAJ699pX22C1M
nuMcJn5Pt3O059Vfi+0RkLnXY8WkiCemZT8lq44spjddzHBfUPSj4McpcgB9
MxAVdTelUrcirnbeHOKxCeKOtEpvZKyW/gkPE81NFt0AHq8+hT+6dfIHYykQ
h5eDymcqaz7DwQ29m+ZsNrQYeLIyIwjb01VoVYAs12PYWfa53TldPInjNLWU
exZHxJ7+HusJbbmANIpcwnq5m9qifUNZsitS6xHIs0N7IC0YR37A28uwOB+k
oMPr/U3f2+CpDuvKLCrxORPEWwZcfoMM5y9BKz4kSscYcAaIs3BWuQvNgj0x
YkM1L0v5g0FoWhs2KWpP2BL/mu+PCpC6cXVoGGlK3N8+ZCOQeZtf3Ywd/7ed
eaBWu0Uz++QsBlwUXJw6jlOOT5M5F8/eaRIOhOaDYkDNdRm6boHtsTPXhii0
0S142NFjfFVua/emxA2SiWqkij7G2jyx6XrnTnviQJtcdAVkbqvzrDsu62Vx
/yFHpPW/n3af+8gLEbGvQixX5yG33kLiJpAriLqVjFqI9mkUVs0Rwo2+yRi1
5z23PRhzgQqfjacMGdVNctf1rNOk1LfVYYskwN/fP6Z4GaL8tSAQlrPIUoFQ
i8/5NC74VpvFHuJ09lUD/dOIBVWcGsitCg0RxqUziffTkxquUl6prJK2vNn8
2k72f7r277gfqrSyjXdikPiOfsmTCDajwaT3UrtefvUVf+0kq8DFofjAeZpc
TCejlG5EZUbpGUVianarAISQHmw4e+Lv2jA13+7yghfXqWtuVtpd+vwww6JD
cSTT8ts3CmoPEdDJM8BZW0S9nDGMGpqzhP0D8krsZvRI5p4EfN+wuJbVYDU8
5ipLNJxaWvjJbJ+wkmxnW4/Qtz1whmU0XYsFZAMFupP8+rGbwbjJsUwN2SUr
mgCvl4p3Fn6+E3h+NE+0otYjbxQ0zSbCt5yqLB2J0XneJlgLbr5j1F9XkIlm
/peraqrK6c7r4fMnsXWhav0UmcQZo7s+gdcw4fy1R7ihXYfjXZyWIm2syJ4z
Esjw4BhxZnC7m/DLdK9ximj6zjOZO8prAmoqz9Y6FfI6hyhnb2LN+dEHmuJX
A/43DRmfIOYFViU5cOrVQqqCEcbIL5eRxgqFKkV7Xk19fyVhH5zwLfLszuis
X+lluw1CCSOi9xsFfpCQN2Cbu+9lUSPUBMkrqz9wZqgD0FDE5+KRaPaN9+ec
15fiHX7o9+2pnFGcp5DwS+/m2xQHuQnVMSdCQP6qCLT7YTWC+ANs9qhwbqJm
suHvveHAlbDHhGJzzcRUi7eWaTQMAblXduYKVLtLM0n+PUlnlO67S/OuZ2Vx
NgkgFMKPVWibhbefXScKWsDq1vcwQAHjsv1u45enquOODg9De1LHyMmtK7K8
61ReNgPwFRijkGUPiaJkYSHGrpma7d+LrniM3HVglDfM4bVbMCfJEmmRuv0z
HRkMbooxwJfKCkcpQGrFvaF/GI+ZtfGovP4U2FYJ3IoG5/Hn6JpZvvPfzFir
nZQBTJIQJluWzWQt+1kbqyPUs2F2TZqZqYtmDUWEWAL/XPLeutwJomDfXKGb
8fgQnH/EyWDRAMpYQBsQZywMrgxxuBP7BfpjpX4xQppC8JaImRrlSUQ+2pYl
xlx7TQfPFNjPkjDuaV/yUMWmP2969MIWm0WNW5upBlJ3m6CRACK1gvAz4gKD
KJ60E24xgfYfulb/fCSJVQ4H7h+B6paDnTrdbuuQ2EGOsY0+r6EBhdCBR8d6
4WSFRmHiLA5Xv9eFYJyq1Qwngv4cilGfHlR2TMhCn03xCOoNcqsjos4kJNL0
lRRvUX7dy2AFi1nYl7YxMBCLUx/VUMdA0bdmUqA6ztb5yGBud1KMECYM60vM
XimDEf1h4btsZmhq3AMHX/QAX2AMThuUR5JvEddjMIz4bNgxh6DO0SCWacYw
wdW5EXYlZKaeNXXQ0DGa0G7fAI08yywyd+1PtqYLNDBTRKvzEUAzg/Hxhr6M
1oBOOdmrtaq7O83UBIFQXnr2fyMbOJNIsUV0xo8QlwKSQ/7maw876773k7QU
8JP00POxkCaA7B99BAkYPjS0Wz4RgegZ0Seax9pKYQJZPL/eG6f2Y0Gz9STc
8V2ipYHH+7218JLtaytccMxYlz/2HH7wmA1FGDDZhsw6g/78jUbrLbD0uGRZ
GguwKp/TAnic5rAVw6aZSUbPTIVx3CpyPq08DWS1MKDwa07KV6avG9o712NK
OKSl7puo/jfTddqUhmyt+LYSCJsdJWN8I8DTgltkhd2qfRnkfmGFDiq2gyxU
6FRHhPclhJ6Ad8uri3Xhit55SZA+Z7ZhX5LqshoWOVu/QX3Lt4Rjer0VN7b6
oU2gWUxPnmaYpyLpc4LrG9dNn0WtbVUnBQeqFz2Sg+0YfQk6HF2aom9zSiXc
/BJNJRLapgnASZQvABtPtEEO4Avjt8RRSWBGgQypOjT4WGfsi6nsBrrqjfKM
g2TgidRm62vFF89W8dAQa+Ht7nv+T9GJQrgM9Tn6lhbOgSVPVOH4Ekt2vzvg
P8aogvF8ndWtQLP0rlMltYOaN2oD5ndFHyQD9ect2unjLYULScVa47AR5jqr
gmcVvB0hgqedFvbcWLw+a7TpX6NidYHvQisrk1FX339Kue1vujhJKpT/dS6f
B/nOwt0l6nRap46n8vzLcoawKF9ZmGAM4nF8G3/thU5O9quR7an1mNk6xEcA
2sb5t3CYsK4rizuVbcPBqfXThRxiCvyasXdcoywLj0AYdsr6PWXkk71uCEXA
uthVBQFyp+z6pa5lahXXUiZtALpT88KjkZUhB3mqfWncuJAQoZr06WNIzzIc
HCousRtsXshiIBw+wRrBvyHMYrRRwIgAj055gjpiGxBDkCPzzfV7hlXYdVL6
t8yh99J32uWvLPWyWGl7uFVS75z6m0IjX8Pgdt1xi+7mdcZAp+1Y1MabEcbI
vtodMn4KzbrOzd9WcEhgIey7Pz+crpVaY+F75A7EgSJSKg/NRV4zcqa9LNta
47D8xVgEAmaQgFFngxNbkzehAqHCT6xIj22wTVp3W+J4DSeAgiNbsFfPnrVc
bFGfzAUemeHT3iIuvcNBxEMuln2aF3quYgBJ1OkUYOlBbLtIlyZ5/gcSJgfb
xV9FYdn0n8xqknMaTq1nr+cIYx0Tlkjey+3AjBDt6zAp3JeUwkRVPeBoxr5t
66hVdLt1vQ4UJK/cpzMAtSq78Tus/BJZYQ3jKiSRyG3BFhY3mSbVZqEKanpl
QTiPMd3xAf47QwowH5Bf//WCT0UbBOMsYcnD2yQEDy96wFsX2mbuFL1O0g8v
w4hnZlk9ITmLy85omsAq7E/PkrU+2Lw69mwaWR2slopVq38jzE6Uc17Kt9T9
b2v7qBmX5Zoq1tWJXCGJ/HdjG+b4P53EySCHOHms2w2ke1zpThzCN2C1Rs9a
z47wdZOIvNQA2jH4PWaDPYA+qznT1XWdjxE8S+UIAFmF76DD+O4/dtRK5omv
+R4WuZAmb4HQME9TMCe8xwojjSnQyG6bDjwsf+N7V2G2oLKtPiTU52nFr8nz
fQvQplUBbXKboaHfW580Bff6RuMXvUy5IuOT5Si4qroPO/3JFCy1Fj3RNnNP
l9v555kg2vWoFLF7YeNmPnlMiwezScFAS/0jwyzOyjn0zdUxjtuXcnjdSgVV
ME1MM0P5HZdYav0wgKiXnfa4BxT3pRwa3YFl3foBvAjZmRgU91YT3iBJv54o
J+OdWCI7kPE2mrvWm6FGyB8RXuBYlHvrhzesD1q/8JV2ud/CPkil8VMSoLAE
qV73qLLHPEyOcIO1FVx6qLHiNuWhVzDCttBRcLAdWHG77bDuqty6g9aloGRl
XBQC/g778LvlE6ufcD2eyPrM1bo4lsT6SZ9fs8aCHgmsK6HXE98O3wwu/J/M
4AIGnJODoJNARBbn7WN1PBxxZ4tBEJmdDnATuEJto4WfRSgRKIQU6DpvP4YI
c9RwnaUHaKdI3XdRf8VxEDfMCheXb7oMybXgwJ1dwMj/iBjD3kcR28itT/wU
VfSGdrwinPEyrPoVtIq5+6SN8nJzNDVjlsGPv6nR/qduXMEMR+DOPCrvieWH
SK44GIGHFA2j77lr8L0rqgXe0GF4DN/CnOKcLOejath4r3mW/Spd91ZIVZdI
iRS748GH2sseXuK8LXZr7FFLmUVTLwhQYn5PALoxRpkao6NMbmzl5FBJ8Jga
IwuVTc80skUqhU/l5NM2J+T/sv4ej1nPq21pjgnZqSiHun1PD6zK5j1+HvQ2
ThblcPMkvrH+gkpfO0MDxin8lwkLotePAYXMBsD45SCd/EPA36bsednU4u3s
kXYAyU12VgCa1+M51+iO2E81aAWU4VauDZCybXiKTehpz4KwkcXGajypoc1w
dir/xYoanQE72ot/KSdQ8/p4/8ErC1uWoil5g1mxtAHHzZ8G3/tHREmpapSK
pqWKk1No1IBgOrE5rGxV8fKxatb3PDuUAbCNPwadVbbY8IRvFAD2r4umLNns
oguGgUgWbAnlBBuelT7x4MU1+YVfTYtOHJopCKF4xkf/q825rn9CDBI5TtaP
Mke3N0R6NibVdXRXoHaxgx9Fa91qRIB9TTrnGdjRz9y2JHJeXWKH7CJq2JjR
wUxwVwMZlpV1pCBrHB2JynPlKm746tjLii1unltQ6fnlthmW0MbPsfMKzKc6
r9zjdagmf2NMsQ146zPqI/bwUerEwe+JKyx9IKew2f8ZKn+Kyd5daU3/N+WH
1TjjBpdE8sgWiN0Ik85l2To98j27CfjCIpBc55AZ5rRRfzhD8H1Bi5sbWVWJ
NwTH5GGFSLp1syLBTl0CHebShu+NTvwPvcXmjXuX6D4YeyywGoQBcG+gf14k
dDLHRCTmgXXi5FQlek9nCPtElyYNlg+PtwHNDkzgIUOyadx/+kIcZg8CLZcN
NiamRstOqKeo+vNuS86mOHJJhAFw/65PLkj4irX81eld2WqWcNw9pbW8hpMx
aXGvqYWjj4T0uakR5xqqMR7coznB3WYbZnmLJ3Gy0h29KdMW6GaaJcbw2QEV
czXRRZwSi0fBtoBRD/IgnBx+yMrJ8g9ZmsrSRobNo7z1h/KP7QRKHOoWjdB/
Q/shZv1Dir71wEHiY3hu1W0polEFPd/4VFvxkuHC17Y/SlAyLKLlRFhtPUNV
ltByrFj5VnhTIrq4Evb4K3gmppyd8J6QAOe/B8HtZDCt4yDgEAFrWEIvEhNB
uTiLH4XJCvkjbO/aKQsDl0iT3soh/5kCDGCAoy3Ek/QYHnciwOxn9yfmXLBD
A0zBkd2LZ0fH9Vv8eQPg0UOctoxsCNr7C9s/+bpzs7A/P97bn+q+s2pQC8BU
5elj+zX+y0ygwj+jMh01O5uaX7+CM2gOs0mkC/8QYpxnDtuAWNhs5nkNSRXn
24DvIaCOfBXCF45EnVUuWcEzME9nLA7tGMAoaYZSZ59TRNmldk9LoFYIvDZa
nDljupXdhxnA5zOEnMbf9Das/9rJ2og4AnoQ0RunPgJwbho4Vejh+U77nWuX
axC/31cO527Bi0c/UgvEvLKqnxGf31JCLxx3QtXR9Nr82noKqCSoKQiRFNyP
QvLsKOvENl2DD0/la8b21TzwdH8teOg2r8Q+pQrJDI1PiZqZmY4VPfAPwVhS
M4R0wTn/6iXGusMn3hNGfxbclqdVn9jE2suylupqo+oy8k1kD6aofYDCHNMS
Nq4tMEbSBf61I8aubXyh/jUAU4cMwdsRNawzSnKcwS40foIKxMV8gG72Eq46
d5mN814LilWvA5ycZSTD2eKkwrQ8FSoSMoD08LVUo81rA9lyJ63Mg+FBXEyb
lY543rEakCrezJ6ylTk5Xk2MeiuAkUKByYN0FEfv4lZGuEOinupqzCQg1pLj
gRtz31f+WS4DyPKkmJtmhjrx93hDeVqSguJ8zzHwIn26FiqV6pK59ALRgvHr
MpVBVIOYYM3Quq1qUGyVjxDdz1ks/mp7V98lQeUhH0NXWPz3pJLsMzXYlNiM
UWfQ9sUseOf90cGSdmpIGHxbOi/YpBiiZg6JRwLExMdq5vP+trmRsL5R/lUg
NhOFi1VTM2FHvP2/6OEKQsH0DFo1mEETNlEJUgbVYkao8ho1F+Jv7vtLCH2B
hFCGXSyh+cAnCE7vnsyIjxa0UnabUuIJLfAUG8+GFQIcMaPiedvEd1ijhBPU
9rfn5Rl+UQOqNUgU9Th6GNKFNVaoX8+4/zeGntLoIwZsvVgMbSQ0NUyleo1u
0bS9tX28mo9dYu568mmjr79e9t2P0ivUf8p9RXJXzKqok4ecvuTmiVVQ+H3t
8TVzrFDjK8rKJ9P/02mHrjS+Zl5Nvt5qm1AFMCZP50luW91/gLuZGZbQ6Xoh
ZC3DOJXw/QqOvwB59rmyBXRMpL3eFqyAlEaglvR9nt8rlB4H5cNCE0PTUjcr
nE1FIOngYZ7+iDTWHHgvKoQKz8R0vCC8HPOY5+/Tt2JVPP1NCKH900dGyiQM
i00fH1SwatONJgSdCicY+IOMAtBMruEpNnRqB5f3jllFpb8MUjq7J4ANBjRj
eY69vSX8ZjD3vaY0MAxCc0NRXP4xYqwMfxkkWLO1EZetnkavOvMt0lUV0Gi0
3tdH0HjO06ss6HjR3nPAG1DjmdORTb4CAZrX10o7kY0V0TfCNFXZIsx4T61n
p+BbbMyHPMCd0czyJdyWZBEs+Zz/gbI8G1iTrTYzp8adXWkamdjc/+cDng4z
f2nNsLKCiWyijp6t4/md5nB6HCkGzKWNf6ttoKIfKrIXnJpiwbWuiSpqqlX3
Fv2oZ3tpfKpincsektlU4LO/r911rIqLL7gpB2R8QbIT+6WBCNFk1xNh++65
5xl8o7NgvbFiN/S3OjZKA68+gthtaVoJzS7m1B7cSKqrpdryE+up2u/c+JwD
If3g0SNdFrAA2544cstnQ1SuNwBKy91l4Gsl2tritc4lDU+tRoWvCLgbjmw3
H9rFiHKBrQDgJ4/urtF84FzgxD6TJx1b2BK4J984XN2nVxBNdNi02hwNJhl+
L4pxItD/Bxcc5ankwVovhf3Kv/UcRY5zfXJDT10ucOwa5SVO0BDELHfd2j/Q
+DWbMbLazCEJWM/+3lMBRtMTlODBBlN1aHZ0Dj6y7fWUr2KmBaiB/EAehIDl
miTR44GbRW4hsBcByZ0iiTxnNRDlElUFoOxDt1vw1wFyNaJVTR+C+g/UvfDX
KSnhVp7ysLLWh9d/c9B/mp5ruRAVk3eltKj3Tfl4fui90VNyfD8RGWVQGKGI
N2S+tjO/VYedHCkfuTasZpUSeD4cX5ONSALwj47lAx15unvuYH0A+4lq3/dA
I5IK+fJz3aEggqGUKe7G1UaeM9qmkfZtOZKDEr6OM9VgmMBm2GdW1+xc/3PC
NS7Z/70eaWkBpP6vtjtJ0/IQmLKiBYJzbGYJ8i6UVSphs9VE9tOKVe18ZVmn
mpqC+6VrT8VjbfqKt73ctnEN062Bgvjo9DZGxDxmPySE1TuY6C3UF0X5+RUW
34JFAs/iwjqwJ13Xqz/ruNX7RVhy+mNunFNByi3ZaMDSgx1Go7w186SQaAud
GoWteBUqXJQwVSe2vOMWDkptNmAOuNnG9KO7YXW5rfrVOp7kgvMHso2If/OP
O8U4n8K1fEpAP6iARSmxNlwDKg3RAtw8yLCRyIRYUTcQpT5BmIawybQGQs0m
ju8D+tas9E8oqAf/+lMF9alefMJxIPYvRLRCIeCUYiiWZNQxQ3+O2OekGnG5
1mLt8DY0I1EK+Afmry84PEItvktGlAQLQUC9i5xlhE50FqDWph+ff3cLRAUJ
bvtYOybuZ1C+YDXcSWUO0hIv5IFFkYDqUvnvCR2WOapc6SPipVdoR904LT6G
wj0N+12zAwqap+pY6Nc6Ev2goLP3qlLgoBD/bHbYgNXfmvZO9tTWJd9T7Bdf
gjgjQeJQSzdbfcfAo7veue6z0s4hrRSfGYfsiF04NUj03qqmIRL2saSSJ7bk
l2bij8RDrt3v0cOzMU+RHa522K51GSV+K5ngcEKEfrCg8dK5/Goj7qtk5qqa
OhfipkTZ3kO/zZHCgeuPS40mPjCmcxvV1SNrMobUY0jFwSELd1NnueNQ9iJ0
uV8+2N7NOjs2gzKvLkIdEltTck5n54ZNoc6Sf3FGqwVkt9qhFGt8B0Yh/qqG
Qy3hLLGP3UTwHphJ+U0ttN1SrKzwG60nU244r7NdSmSp3d5vbY7PaBatmx2s
v9CXPoj5qaf2qmRIa59eYWYUAqEPByoxLRs+iIS6VEIZ+ocB4UwMHyZr8v/s
333Euu+DU5pgXnMvlP8TOPIsGGpegL3YvDXO/JwmxdtjOEmgMoAbssI7mIq/
SIppWsdNdfZdfWCf8VBq1DW0N4SAB8NWCG8wf9BYf28tAyl048WsWzCkwQ3l
KwmV+KBTPr/oug/gTVUKV6w7njZP5BoHNyFhDbytdRn2VEDe98ZXTw5lYSYC
9EXYdUEC51iKk6yAVVQrrCFB45NRxcmr43Repg9VT0/lo86ieKtRywGzXOe4
HaEmBaiy3ecvATFaScKyRbnSzjRKenPkRYyllrrAJBVD2jX2fS585DBgq9Ux
8h/UMpZYpsbLi7DL7INs1MzhTks7S6UTkLnG6HQpFlAUHG6mDhVJDZV1gUKL
EOCUAVldqmxB6tG3vpW7xd0UHXWEvni++GgKZdRn2PhshsNMmcP9KwSqpNW6
y+MFFTi9/O8lCIAPXYqRKaYFZnjeS+hLZ+ktLw4zMpO23jlIA8Gbiy+yhJVE
UA8MGCxQz4sAMf+Klb0Dj/hQw9cym+RdbozoOng1ryVs9nHOZKFPoTXljQYZ
lIpAsU27npGwXff4FRXmKq1VR+x57aR1soPFARopoLnLMZ9JGXW7z85k6TGW
oza1NE5mE/Yzk6m5Q3fF1648E0HrshlM7+9c7rp2J9MD6G1o7/a/6MpkupfQ
X/fC9PNOyK6CUtc9HF+y6zGA5FxPlm53/fFdY9Txo/2iDR64kVw5vtCWxJKD
LAmGcgOX53Dvd62yQYIlj6qa89SeYMfnshKy8YAFZhrNNx+u0DsZA0k/je/K
q04TwjzAam1K3sdrGG9IN4mOBZijUmwt3qpdkOkR+mTl8O6oroPmSEnPZ8SO
KpRBzM0CIf2n3G93E4+01yvAdYOeZPZjIiwwudVO+prLlhIs86Cqb090hJNI
3e5HcbI0ijF58nekByxYxwOB0s6U719dOXjiTGlKFq6NgbxtyyFolqP6hZC3
kz44ibLOBPltI5LEQ7+mg6LJpBMTEsshGY+g8/wlTgFPUoZirFWfSyuesD9n
d9vCKXW7qq396h93uBd6RmJB6P9B10NpWrwwucKfsTEBEEidM62fPlqfKGbR
vFuT4Gt1eXtna41PpoYyCnfgc+GdN1CMzZ9BwGGtPu6zLBsy9NX17985YX4e
pEtCuaB9v9YDRqO7oRCDZ5bPxZsu7LqBWZQ1MiFVdmESF2naUDbJhziQRgB6
bmeW9YxgYQnlzFZlILhcautTJM9J6clUkcGD6jxVYx9vAV8c9vTccb8eVb6w
sombgf10O5task19lIr/GMu5R4B7u79P6qVuiuSmwsfh8DheLi47gOPIU1n3
DW6gk8jwI43oiRloaKij0fOhiV97hMLQxJvnmlx66osWOvy9AH6oSU0jCwPm
V1t3wYEUsxjahIbBqefOv0Rb2U/N/sNyu1uZHoaCJ3A2HQCOQDqzxY4jC0xX
Ii+SudBmrR4dqY6EaKOFlot1471PLmgGcwGYf6OEfOR2ssvrlIZGVx3SLMpF
gz9HbztISzQ4BYC6w9SDsUWRtqgIpg3b4A7AtW5AS+zAMeNkEQnVaQia0yTt
rvWDR+rBRyzDzmE3SPm5GWtRLhTNFxvKWh5lzYz67K+FZoAECHgva6KG+Mgi
n5XGgWlQWX0NcvM1BwK84y7DMvofliJsfRcSnVClxFBWvxHybKhLJH9vIxBk
7QUJSIcxiJHkTzh/iW/kDr5rmEMiB5v1RdUkykQVL3FVbTQQuv+tjTmOMnoT
ftGF2kGKGt5idMceDsLegztcyp/VlalS95zAOV9bb6zg+YcjP4TIwxTmI5SS
GjySSqyXKEO2+wJ5iMd4xFQ9bl9U76yL9qtJlcRyq5oHi0Vuj0VF4ARbNx6j
grkHIa2jFJVr5iGH+RGCQwsYCUhu89OFvECUKSYWsKuGM8sW7jd0MMR5Td60
avCaHBpZR1eyUb985kQyEGpiEgsohmnMXsLzk+3CGcLJA4dFgTtrdUdwoQGv
KJg7fbxgkSK9jOgfWTflDKWqOU/x0do1gEtQ8EkKhHvdtMNrnAUg+hYvaJtl
TnIyJm11/nkJBiBe6uJPNZZ/2iPee485eG6ekIVL5u4Khz3Pb/to9m0+HI6x
HiT1RDSUNF2C9LiTY6fvye9JLQVlFdnFe3AFIwqn3LfyTZ8nvdpQsiaTRA/Y
sGwVfveQTWYxnnCDmNoOUVr1LBOB021+8GOqmxTQk5O62LIk9KUKV2v9SxNV
pGBzEJh1gub3tpqDVwtCRbPfrSCHLAOyg2xKEdk1pS76mIgpUR1P+3WknqUu
RESvn5SDQ82kH41ij++8+11IldivVj0yhvFDWKvdOT1CT2L4RgRv56p50cF2
eqEhL//N8hj12ny65IjkPNJGY6CtruU+3rEYw1pu8n6ex6D8abZBp1oyLM2w
1zv/xaYFIZ3097+utSIMDRC/oEX/C+kHas8YMaHKkgH7Vu+F8JTvu/C6IJRp
by0jEmqXhwV9zqxeXje1YTPVQ/sx7JcWkbiQMxE6AJs4SrwzbZ+e1ocsJLCE
8ASHAMXTgZheA7PVyzcwaSoGtqNpbV0jQL6LnaijUpAkcTnhHQX0VOYE/E73
fAW06zUh1TA9MOv48EG18R6CidoMwTCVsY/b1JRyjaT88JADB7KDxOmuJ6/d
uMVYuLUL7Ct4sivvm47gBbuSVRq/HdOMXS855vAx3Kcunk8U2M9tF7jnDFcs
nW6+AmCuKBH/WrKbJhMPR831pXwr+RZScfmK2xc9gm5bSZVxNoDaRFErwxD5
y762AdHljSrF+MKdSIIxSWWVI3kPL7omQ1ROFILbkXtSLmQHjMwBu+iGQkqR
uN7WeX0v9I6zHaA+EcfvByS/XoTLID1OFUsaRHy0QujBAlPH6z0cFonN3/Ml
TRDKfz9BbVXq88SIct0iFkoS+filvDFP6L0wVgAttJXZ08UeV+GKdrrBFvxh
7ZrYpY8IEteIsXxA/FGy8/DxB09i6zZKZ+ek102vCeR/lk5yQEbqz23Qy54g
xsilNPku7kxiTWvRUYkdAo4SWsRoBrVKW8zQqLSdlqY5AIkWbaZpuTHIkRB9
q/AIV8Gyfw9VsnUipF+6O3RriqKiuaB3tmHkjzqlkSDSWFw5rRQoDMOeHTJK
ULn0xis8Y8S3gz7lzmMYzf0uULaM4Qx4S1VGMyj2iyEspo1up9bzmu2tjcwE
ipHAwgeXsE1vCLknqn3rB7VulG469sRenWYlS0yLUFOHziWN9HLkOCDh41n5
NCOm2qZwCSqEWD/UDKwBSWe4r+UUIkUtK36NK3Rg/pwGMnsgfMT5YoZBfeer
oB12ICrAoWoHrlDhRrUsbIWbYJJs9B1oODGWhZmcV+/MHEF2VB9dlRtu3/xL
ybOxEi6G5MBXjTeLTpX39pBUkLax++0kzox991CZaU7gfuBJFfAZhPumx8cx
ujVTpMISRqm9Gu7Mj0QQIF1u3pkVa1uJjdMUax0NuSJKl/o/dIfjGkHNpyKz
HRAeAkF7o4BfJ3CszU8umYmDgjyoGTqYcLI8r7QFLZrB4sddlmMQNZ3OVcl2
WhYHuS5Qj7aNZefzWXKgZ/O1i3onapDGSwJtMIYFnVg56lVy4MbOMNmIcFxQ
/2gM34XRurtTBtT67XwG+4/1XtG+r5z+m0mfhQQE/jkWYqcUTB5n98IykpAt
jT8A+LGFMRHOWTEyyw8VMxfI+mdX+FFR5lH5md5vowuAwZ586gonEJPnyK7o
QBSlDDnFJaaX/x6Gw/BhF0ywxSoYDrJvaYl7Vcc2lx3umSfJlWxhsUuIuqjf
sQVtxvnKrZBbjVdPzRq04yG1YcazFWPwQ3uMfAcNjvi8Iq4VMcZkEp+XJNna
Hi0XoL8fTX+NzzMXtFmqeQNbSc/WD0G7k+AQtBupeD2cqKFujslyLbTl9tf6
hP958ppPndv4pkZyoC4tQkl1mnQT3Yir4Q7fURXgEWwmk+aquYmHbbkI/laX
a624XmYUfJrghtXCVi5NDVESeHUDQFZ6jJj2anGJuBfHcPvz1kmtPGefllKw
kXZOuImNRnAEEUI8XOi+tZsuB54Qac8ZNArUv1VYnELErs9IKn2b4dm+r0LZ
zPJN4lg77S21VAQYVESMahJ+HnBnhxfDDNnRnN8R9QHHLedDJNwd6zrDwlMe
IvticNvMtVCLNXrstKILD0ZNyyZfyb+a6WwkL8OO/hBRLHBBZ0A5uSo5L8ck
aiuIoGhYSNQMsNJoCb2e6ac3MC9dbETAm9y+BrJaw+e7LTHQoIthpfHLtAzL
FoBPqw6wehUv/7QH/AR32JVFvz/pqZfaoEShDJkh8E9pJOWa8EObIteuz7g9
Bdz9FtRnFJRYUdewZA4/0874ZFW6DsUhw+fk9T5LcYPH0tZ1Ej0sfu0+l/it
DsTwJo4gcLYvj46bJRF6csIIJAfLerZf3A/wqyenBp4hEAIbIB9T6pzOQtAl
JOJWrezoi9Ros4wIuSg4CP+Uklyl8plLRx74AdSK/VFWdR4o/KAglYiKF/s/
egKShLPd3t2xDAq+A4E9d2n+VgvYuCZJ4r+MhCBdcwkl+xQfFI7DIcGWSTrm
a6HCVu1D9t0A35X2oLowfOaWXcQaNfJQ2PTqPYQKlYM4XcJZaaUwKemFz7Fn
zXcUdN/9HJ7CSaaQi5p+pqgS9VsV1hRp/AtsNzwFD4+7orxihEbXsNZF60zS
YubXbmXOV4/S/FQ2+2qqfJu1CQPr7nn0+kidd/JbXasl7E7eqeItnG+bIZMI
als/9+1Yfevnht5S3osHTRXdDNxNRE8rzSCYFdV6zyvPTnFmGUNRKEZzst8B
/jwmJVAt4M81dJJPIbvptF+kVugak6myw2E34qFBkbyQrgJu3IOAxe+m6gXw
UmEO8NscKTkhIQbULHth3mVNmA7pe0cPacQPEuUDJrPwC7TSDm+IvOG7ttut
87kmv3tflMJFWzCWBQgfUc5uarcpgyr02x4ZpSWyN4GwmAtQy9EUvfrCuMQM
uLQrinFtjmVPGAKTG5Dua2vfXiW6pUvvaQwEkbOc+jEnDd9b+yXN5B5PCylg
i9DQV/dI2BD4Lf/7oimesVlEN/jh5pJjnOftJViifHnjkATFfX6p93+duPc7
rZTPkT42PhdE9JRP8IvahuOf7D/nibqvoMJ6qhjBV2k2mmy1Y1TzBIFsvRd8
jhRob5FYwl4A1L/NK8Y3rGY/ByLdu6kkAgLtDSuTn/b+2+srm0TkXk4B+aYa
6gDSM5I8Ycn1ZxY8MPTFOKrQT+5xz88xfqXvyAkrfihSUTsn+xYlHjQI3EMM
cOjMKkgZsmpdiSFWLeDhkU2MuG/oQzdIjPLTk9zYr44UPSrmDQg1gmmLbmBh
7x5fNJLt9g/EtwOcWvXgGbi3MGnvjJBU33hDGgiar2arvv8UaMzlvb4r8OYT
K6fVJ4bu+nmUBCZAhSFUtuRsIwJw1bZxVWf1kb4OKPYJMdbRYJN5jdA8MJMm
j4LHEgSKtCEoy5/XT35bic2md+JlgOmxQ1PaF1vY0QwpviJJTuBVPOpw8/2k
/BVaJC6gogEjzHGr4z66GszVf1nfby4kkNQyo130z3KW/XcC3Pd6cj7S454g
znCN2Ck+afCOK26LdWo926bRK7UJeSVzgzqRqJrv1i3fHl3aU/sPNv/4WJ59
tzlKGgZ5LBZJnvZy9IyMG2uSgDn0/MZ+Lupvjd59AcicHcBYgnJJy7kw0G7A
UhaEitWuSLoKHzDy4O17iGtd37YrrCSi297Q6gB6rhjg/zbDd/rgq+zFUrg4
3TJFbDiN61kTdOS5kD1/nu1LRghGIUJ2j9d6+M7Jr3pMUUoVye91QSbFSiKP
Sun3ds3PpuBeOM6fTuColW2+1QkQrWHzqYXLpvW3V0usOyfGyVKjUJrozPns
5CMYnATJD0ARQoeDdKiFbUSCtIbmLbFgVdjsAL6sTmYgKM6YxbKq88q01u2C
XhLm5e+CzU68vPqBGlebTtEF2y06jhywJdARcjWfnjNx7aDmk/YqvjxWYHqA
fNMASYxXE7jpYkBL5hImxNMIU/we/RTTYqgquebDsAX0MpG20gBmk+pw6hEj
JXEGH5v6ML65ek7YSRdgNEFfqpZXFKxQO40KpKs+7aDEzsDZSFLbnbV5RAxe
y6YxqbeMo9iZkFZDDut3owrI6daAAhb1lWl5MHPrF0h44YdZx0lcx9TRL/iQ
xIXyEoC4t+4K2qcLF+X0X5cxj14AkcOfbD0Gt56VEJypwkYhtewjnrFb6H2u
dCTZ5wI/JKLG3JVrUMzmoMofGKfAw9LeMgAzIKLWIOObchqgzrGLWdsP5hwY
hJwLJLyOl64tlCWRk6fVZKy6xULT2+F1eQXtSpCzSoDQWFCW1z2S7a3N7cnF
BD+vFCEzLLgvzmOvwiecpbYIhaUaq99YAVMyugauT03xcpkhyRm7VS7EPpll
YzqxSMZArwJg+iWKYOPPHICiRhOEKuwOEggEeGJzQy0kVdfWhj8uQxMUmA/e
i+kbp2LC9t4/AD64F6uzfOw+w6pTiUjgJNgaB3feGqIyhIWxLOyUThdzvJIM
ZcSTcmj7QVdkvswMRsyJfCMLVY2CJ5K4hXgVBCSjkhCxTZOZbgsc3HeqEkBE
MZpQtTjl5/SNiFVZaAS6Qmw/gXq6vV2KEONwSAviI5+tZ10nOTIsz+q6LBnD
fqCIKDvMqXpNA9NDYJfFLv0h5/6kEd68J7jSZPPw6nj5npKYiNbJ7ngn1Fkc
A+QF6pZUANq/bMmgdUYVsyIt1eS6HPO5STsN+t3apxRIIYMVEn1gzwtyvyu4
huWQxB4ghNCiEv6BzXI2/+qr7/3QAIEUk2iTLzNbrZAX8mK4EnrudJyePEd4
7B7daJVR1DOy2dDbr9qJePYasc3ubSh+rTJpbMhWcVI2LHpER1Wc1h69XXw9
6ehQ8ktQq+J+S4ZvwmQ5Plvqm94syC+kFHOdjYfHyjJTdor/VONCP2zHSOZ3
NXqh3vrb4Xt3sz1Y4tQtqZtmE96M1yRVsSvNgyiiAu4duuzQdKH5EDoOrfZZ
zfJIQGmswhZIg9vF+0eHlRsWFruYl+lXg0pYgYFEz636udpXEagnMcz729qx
M2+GNau4V/3XPYf4K1+jvtYEY8Vmhi8OrbdvHqkomt/Tdsz9FhJjJbCNu1j7
u5SHKp8ZSPOP+d6R2L7vuC5gEwtvM4A9AcgmfxKhiopGtqNrA5ZiYhq3ysa7
qCotWjD9NC3MRuVDFgFjJ5OmJ7B6OWH1yq2qFV8BKeGY5NObWb8kpjMXzyiv
kwPdrC3edpfwfhPumDGiJK4vutVd3riNiV5dsargvv+ylwD5NdjV77+IdSy2
cjXLA59x9Q2KkVAB8vGsbz7+RL65oyUTbP5DCe1AevEyOBu7m1dvDnw78X0i
ypTt2bghjRC5VC0EZSVPwUJ8/DcHo6Z/m7hD0C+x6ViQw2jOHM7eeWrs8x1l
8fjWcQpS8AZWAagkDYPKkEdsa2gTYjy5gFlu/+rxA4HV4mYpwwCj7hSGtspX
nuEQU2wmFMYQa6nGmMmjGdgzQb5asBoSlSljyyEcnN8NSYPHz/813LL5JeC6
3mp063ALlbxIoJAHi14Ju/T88fggOoUsjG3XKj7aYCXhvMesaPU6Bo/U7UO+
TAoE3QY13qlNzkOdG3ZaKTOLGR+ATssihzdDtzUUTIOv1seVTnkK3hZVTJSF
cU14uosycki0uBXQsqKrRBkGx88LGK9vCnmPidlFAmKMf2AS1hBupA3Mdtuh
u87Pt/EM5/cvqR2Pl19AHP3rI/Zmm9li0eSTqvr2tXnNBqo+eBZlCb/WfTze
KpHHI0jIeRNGOqOPYNVG2b+KE41KQ269B5IlURaMAUle9EkJaUbiUcM4dR46
guhfyAjsCBs5qiQihO+CuC1UdIBGnRAHAQbG/XjwIoHbhELmQSRRzGxPfopP
IXBPTdb0owBrOdvw40lKHA0LEiVAwj8XJXXSbVl/gerYvq5k/Jdpbmp3/9ZZ
/vQWNrgKVitIIKfwZiFlN97b10+1EjUs/kRJEkrpsjUL9r/c8s1YmjAKXqtN
MdmCFonxAdtnTQxSlUaafvPfJWhjxuLizmEREXVGjlhZExzJYFFmv0KZNtng
NIUYD99dB3w92O+ZXrGAVoj8MkrX/IjTpX1xktut0AXt3+vhXlPUbf3F/EPs
5SkP1vUXdCYLACZ1XCV2QFkiw91FvgC30lbZJD0dlQ5O/ORHHesUPWuqJkYL
hYiU1LhaqppyGJDKjIdXF7+SSQhtfR70FqjKNjsJTVLPdjp/V/E7C7gjJpA6
EYBKdlZVJA2Yi4fMmx/cq7RddwfPVVPAl3C+/ndbj9uCUZP/9+qiedcIbSZD
3mwOBBKg8rOnu8z+ybxpUpqhSBwv3PYTGSoe3RRVqNcW9nNia6kvEg72DfIR
R4cGVqwFzF7L92jqvf0+thqjYw8CYjZ3L6DZIQjAx1dODA1LE2Ey0u9xd9fx
p6H1h3Fn64AbiJEevc7aGEPUK1camNkYb1QNXbR97aC4HXXMcWagxSv1GPWA
4V6g453c1HgsIXXXsluuht3V+tcVFzbamXyolkZ2hhzILWW92PrgvLdIM3IZ
Ip8qjsTrfsQKAThFe8bb3Hflm15Zj+C04yoVHamnsB+YAXdbhQmaYoZlfuVy
nNOtaMussmjtNLpM738zjMp3WiRaZ1iFG0aQJkf7z6/Hs0IWL8cu8AdhXxR/
R0rKSadJ2CB/seW3YXagmE6uGF0rU4p1Zv7jp3FXQz8AOXowCF08azv+Q9uJ
WnlZwxEADVEKuv7JKNAEQLwVtqTP2kv1x4qjz16E7pAY+n9hDNtgMaCm3W1A
XDByDTRMDCSozPTSwHT05AG+Yx+6cWqrh6ujYCBIpz4YPJj4XizOhHK0YgRB
Mf/RfbRKDF4YvDVy+PNUKDN1lI74zAufC0Yu4vp9w88rx0g2oHEKSp/uZYWv
k91yuhwtxMMpCXtp3efHYsSHMm1S6BLpYKYSj0EZEBKZpYCUAwJfYcOwKdL4
ytWFYq1ieGibi41g+b734bwYUmHp32HPTMJcTNjHknCHtXQhPMi8JNAtX4xv
KsPoq7a+AcmqSIM8oLRXsr9uAzESIWP1PZ1jszhpCxX8CGmc1w0c2cNW6nju
fZZ4/M37eJlLNp2eVi3AtyRT2XU2bk9qG9MbNnIzXdPAGt/f2sMi2/d5Kr4+
Ii5XjO+PkbTMRRkcjnecv4esANLkti+sNMDBBu/aOEjIO/468HSpuLdZhe5T
Rct8eJ1enLqA5AOYYcrXUI3b2tBjgmdEjOiVxjg6pqS03VdVxNaljiIPlk3n
Ci3pQTR/MgEaSE2BwjwHr3k9Vf+px0xsvKaj68a8Ixdn5nzEBMoMnqmjk3JQ
/b4V0or0wfPx5Mt0sak91H0rUCVzoyxhh9+HcrS9CgGadC3ckh85rU9NJ8X4
AKHDnCECOpV5OOujBL5TJVOyas0fU+Le1WisVCmowZFoMCRLWcP1ESj0y80L
kyTjMVhfhbyceQIu6BUmWPfmBMKiWVMm95pNVghKIkUNuWb/yU4qG8EpxaNT
rlzvrx1qlbZM/bTIot3IpGfUzocV6/F72V+fXyfhl5GlkqQwggeF2IRF0R/3
jXJlNZxE8mg/80SYoQFKWRTjJW7a/CbKOd29cb6OP4oM+TBQxh35uNAxnzip
Gs+esiEqpopYo/VQmFRP6V5TmsgYJX6sbfSvt1u6ggrtJYs23UyvFDsE8jZn
1vdtz7XrCgffWvqyQT1NTgxFX09w55FFHOZgVlxKoEzDN1Vug+I3Ht/s0MYe
I+g/TIxR2AWgxXrg5sQVMdK63MANad964Gp257CXKnhh9+ADibyiWFRAg76p
SJtX6/bWpSJnqVA92sdSYFMSdei2L9N/MXTAX7x+t012Zc86XDRLLjgOBE94
5k9MqfhwoM27aCayXfGmDK7JD6OfihwJG7j6hY9+6lrvhYcds3B1BQf4C+Za
jRrcz8R/Zns+rst6BuBip+oNtTIOJBlui5y8vD50ViOXV0QFki/5Nnwpd3oC
mLHAxqAMcCW2TIzS2LUlwaDcE6iWGOLSKLOjgAXLqy8UJ6ZpFG8j4/MKSq0W
EK9ivFtVFHC4tKa6gbo2BNeJ7SENxoMsoJVfNR6nvPcbKE1TKohsKU//9k86
c5NQrGhFSi7NYsbrs0oYRILptwl4VgTOFq9qzs34V9r5QSjFFMQssH8lsOJd
pnzIYuDKcKW/jx8To0HoogcA6I/VPQRcVhnYKmGsrTIGI6oe0YyU01bOk/1P
+Da6KwcAEeYohqRwcnVaORBERZNPjEvTJZb+35oFHn48dVVVS6TUydL0Cvb4
WbabzgA5XBX9/0VYx+jFP4jOf2lJUOQ1X5oMqBPpA+oonoHKWoSBfnuRnoYH
uZA3IVCqiOSNnGGCoUQ3FvUKfkF70XhJRE11EjxSotVxwwnO2QOMJZQFyesk
9+YvY/p/YqLUElNfvMp4tEKpIpW6WCTySVw/vIEa2gl0ER2mkd88iL2BVpg2
9DTiy3y0WlU36a1bwVAQXICl0QB8iL8z8G6yubelzS1RmIPLYsNhS2/rsgSk
qkYsXFLacxyEkMX10NzC9DMB+JgZiPyJkHZS16fBxFAsI09vhGNzyH00Tnhr
e0VRo72FjfyBRDJ9rhLQMVX4Gce7OLRrgMLOW+vBtihtOqwSHEMBr0umHWcA
eGbfGHUGauo7DuQ9+z9hUAcQeIdzUcagQPaSPCHORcmlrWhmzss2IdKigvX+
AVq1zoHb262rjn63RjKZTfo1wqDMJBr7Ntp+97B1jcB9Ki5XyBD/7/EWpDii
3Xuq/uvyVo9Ivx9v7x/CQYl1U/w/yshgVx2lagWFfY4OxCjvXin675ZRtzSu
iednvcbX1gA7R4/c4U7fWw++zHVVYiRLuBBjl0bjUBsjDKGCoO0ZdPaU2XQC
hC9/BldyKSKpShFW3R+vAmt6Dfv7mxeZyZ8Acz3yCzp7ukUpKL/tJfpWw/Rd
gVwCoG5iOJnKivVgs534C/s8hfWkWkEc6DJ6eAUrAzudWZe4QeTQq70pKi2z
zOSyXvS88vuE0ERuePuLTqw+sxRwykNNy1Yz8tNclJkuDZCVcGXCwLvrUB46
mvFcumIl3edMIBvUmzM7b3FosS9v8tefrlLz6anKDcN6c2BmHAOM9gwzyK8U
9H3JCZDweUF2GZYJQbzX5dymrJUAPdRJl4MpQD5NYl5LYfOsX1BpB6lViIHQ
xpynduAiRM/MZOfoTnJmKTXHeF35KWsezH7BZmvBYiwmTSruKJjs3kAeiODZ
eVp4lriPusObOsjXMXto9HLMaS6UPuYPZVwrf7MjheS5GAZjnoVApUsSFJbu
YO0IoMoOM6v53Ag2FFLPY0VFt9q9LHnjZ6Fe+T3rdoBJJYvIU7vGWCUPyxZq
O73/GReKBLlrZYmZItftsekCD6GJWAxODzCiTVBO3zzd+lsyULB70OtNyNaH
8dSHnBexgxgIrWFxyAUfE7q9u40iPfKo1+Bsdy2HxaQmlw8XYT8ocinEPVg6
PGIPlzxpY7v7nOFeYKoZejWn88m/o+0H3XTCsBu+viqVdmQDlzXmw8VNj//M
HCmB3udzgG7lcrzjBWZTELicnE1uVWw2KLiE2tp6xaKUerOn05pMGbdQ0kW7
x3xHigAibQGK+mn6B68iJZecj0iIaMpAPkMqJZSaeH3tCka7RloRORLf+lkW
8BrmHnKUffNRFeXhYYL/aYgdIz8v0URVYsy+2KhfskT/HrjnbDCO1uUa+/Ys
XjMyXkUOHDMcZuuLmusOJlFrhgD9bci9ZprkVtatjLE3Ang2xB8WSxPy1YMv
HPqfkUADixGQj0YuDLAD6D3D6J9aDqUn9p9gcZ5vXEU0Ja+KQw0xlgu+D+sJ
ePxTateodOaJGuUQ3NjfRzz7PnVAikMzIlN9zDGp7ukwrrYop/5WTf2m0ezY
zk3FBsIqD8ZBXt8N7prhwAvC2KlxQvkhPMI7FMCLT+W27hAZC3uMJXf2IZub
mU3gCRcvz5E2ZVzJhJercp70vayhotG/XbgefdaRpS+RWKRwQeD5AyAUEINA
WCmF4xMmjB72CnSEuZA6UuVV02JEkm2+XvSqd012uZTMNgtTnZ6/t7CvCWnC
3Ex026AaS4z1Fog09ZNRDDcfJJ47WiH+aqZJRIX334GzO61G9A1bQQiHinSh
698oRu/igzSUdEperSJ/LJqHqQI58P7jJHGczf30UVYPibnk3e+HsvIAL2kh
EzAL6X+HARe/ZqpI55QYJzQsutJrYLkL97rytIMen+I4fdTt5ZmKl7OjE8E8
xKK1ZKPRTmI8NKrrgDbddYCBY3nWsu4sFt+ofNBffCcqXLRkuG/u9BFVguD8
okFMXQMU/mrLTigTbgsLt+Vwzu+lPgm8PaalvA2keKTnZkB0G48JBo/IapAF
0Tr5uP9HlmLZdHTM8Pkv3EUKwMYSWpnNRwc3p44qs3hyoYeQ7P8gTlOCGQHq
chSA47dGVw55zWQP3CQsJ5RmM1LpOhrXFIZ/LfwJMStJ9vLgqux7bto6lnCK
neNvMLrhNli/+PBoVTcYRqTsY+9dZC2LHLvinchH4TIrLBZnjrFJH86rtbu5
DvXqoH8sMcQ5vvyUTh4RZCmOubehNclXwUJxSQPozSGvviv//BcKlPLnEJlP
HVB1nvyvRaiWRTGYc06KfNt/E5UN6jLRVSWISXX+Y4NWvlOTTKntKb9So0z2
v4cKjK4SnzrHlEBDIIan2oiRd6X/1jK7qrN30C9x0oEQlyJ2tW5Px7nml6av
edgDrnaw0ZceAGmhjvMSos1lXmllZ3qULcifvsMvL2nGF16NG7lnDSDBylLx
wFWe8/uWfrCXTYnFLlx8w8icuGs2yUQ8uXnSsE/5s4tDhpjhvi64FCHROY3N
w/zYl3wLXKU5/PyRtcBzWrcoPWyYpNgl2wInl7D1OsCgydz4Tkq9ZUZfCqBu
K4jEDeh/BlOHcZgb0wE51je87WLuzTaady3PQblBZzVbd2Im62y5xD3c/CHj
vPxuTzHHe8hAUD/OrIzX1QmWCyF5aLP7MKE6C7XC4YDDJh2S5dhVf8xV3v8N
Dmiarh6j/S0iDzZNWVUjbcw2X39qCqIwTZ9nO4pFKp9GIHnqNOXcjHX6le36
MsgZobUUPEmX8JM9gNZ9Z1kscEc/uk36t5QMQ2LstZOBXkeiF+offLpj1MV/
l8DYFtttlVEaYlaMmIWlkqQ9kwCKV0rot7wpmtv3qZLwieqWRcxMHLJOdvC0
BP000fl0FOuPsDFfzrDPeKGoiPL5nnkFDNolQ8zjblXkIVEy5e7FDXBU8grb
ucwldAaFeUYEf3OORyBslTuVNr9jrGTAC+1p2URSIebVsS8BAYvJ0jls/pOq
lbZtKt/oorwrocqohqqgUeGF0ZiKpjWn9IlJTEMD7tJM92yNNz0I/XEOuAr7
UZbcnzmfxvSOuOhqfMg8xrh0bIaZJokKu9JveO3K8wUpdJF3fnwh65HnQkRD
yBfT+rShUGaFUdjOIBTnLQNzSuNhiVaUW4TgaFUWCgHjDG1uhQOUKaT+4TFw
wX8285HhDIY7b0PMvWhtN4UYeK0CBe9hFoo2RhHsML9Lan1Pdp8zKTp7Ek+Y
m3v2ZKp3a1EEeYASMFw7PUf+ioojc1RcIdmTuv61xLiu7+uPwuIIgRprkSu+
GFDtcF0tZC5bJ4yCF2Osb96Sd5Zn8xT6X0QPt5L4A19zNrcClYL7oRH2CjF5
br0pIExlHMBzA5igxO+6B5oVws6IkJGXzUzCerhScMxnhKE6Bu2iX8WIR0DX
UUUD/lQH56u82fCe4cUX+Pp6UDVSfyh7rJS4Dm7sMVL/nwJiVfJqhxpHsETl
1Itwe4yDFCpuMsz9qCM8Byb9begoEMqu3JaFN8tJudh98xYKdy6zlPd+fzsO
5tsdth3T/dDwtX2Dz8qlJD+p+XvXrtnLbPW7boIe/PrE2rXLuphPfaQWjQv/
zR8NNyGQ7lv0CrjgdO/7oeANfw77w86oQZiDqj3EVw6ZqoRYRNPcpFkm/Rff
5XwBXfQELqhhGwDWjD4AAI4WNuVA8/Y0AaXp6o/4/1x1f+t7Rjf5c0oWDkLP
vHaxIL9CRD52/bMt9sQLix/usUAyvlfbRi3534C6lQa0AaF1V5e2I18Gk11g
7yz6SJlSO8sWRjOoQIo1RvN68vFu5YE2vF75jkpraxbVf6FZEkmqGRb1OOKB
/ucj46nlYuxKXL9xMLsHy2W4eBf9OfVGP+0CdNbRzyPpzAB+0iaCLWCQc6rQ
qzkDIgaRbxvvpeYyVWBE/NrfiIwlIfrIHtX0GmX4l5lOoIJwl6kCaY67a8Dq
fTdbGMda09FhBrt6Vo99cBnTcPhvJFNhnMfGnW5+0Uj8pkcCNKj6KRFRn9CL
F0jEtwatldsA5/mXTJ6Y40j19droYl5wuny5t7T4c6Xi+ZObnzeqkx7UNya/
KIW1JygL9VZaCbvx6zY4TywrViKmMMtDgKQmexK+NK9MEDw/N2rYqjaeEx5v
GY4dN8/QTjCsPb+PBUHtFRjZkHEoOFiK6cjp526lU2cJ/LqBfDGGa3MoxzHO
hoVFBrUuiqegjZ++6U4pnsRuXtSHW/kzZn3Hk8spzS4k9j+cr20L3ymdpIBO
SXhwrsXrlKbWNVuAVKXHYhexKBZoz/tnoxKDCCamA6GbFmIU3k9SJejyvJOo
Hcf9Oh2k26X/N1S9OMeGhrIPTsyekhAneEeO9esVU9DXPIDRzo79rszOaIIm
mv2lpG48sS9R1M8mhQdD/s86xaeBac0gZIMZQyZJvw/RxfRHxHxCkYIrLT12
aTkEgOju4Gug8s6XLcI+wnLOWg/AaNbO/mRg2OyXkMfh3BaW20pm9aoAleHt
Isj4RMUD11QORPyJf+obno2nem0wcCpv7q2czqbsaYuoptP5ongqLUyjJb+7
Vg0mXNHsEfouDiMA5M4xf9KYrSAtg6bkqmqmQ+rP9O5OiYbKzLr40mKX+Uwv
yPdPtUseOMsZh7RXl9yOgze/W6QEgMVQfBQlaJSMgA3bMWlheHm07wNnmDiE
EMFzNhsKnd4ObkEa3Gbx/btqV3ZlauLJdUI8AmT5Vqu5I7u+fFnhkeCIe6sr
J1R4gUrJTs4Lf0iyPbgD59R30vdwBcwGjjeLpmrqzLUm01qc55cOjspgm4jv
hB8H4ZQRw+Wu46PL3bc4nKPZxA1Sy+T7LNwQK3osXGQP1Cu1ceShnjnl1OjC
Lk8AMMkfrTQbpqrR2vPA0yVtl31UtpUAQPCxR9wIt6PB6TeRCGPf19GvN62+
x9QJumaJvqF3zUbeR9CiF+yTC8ttpLlcJB1hCydhahKME1Aa7loWxNVBp4nE
mVKZzJuDv9LKhV+W8gwGDoFDlVoC18yosnqgP6UL6bZrOEtZQQi2LjHrwCng
JGbtHAAEF591UU0Wl6nrHy4FquLR0wCdQg74BPwRwW2gH66tnnZA3KFVC98L
F46zFewl8K8xJvOE/vXDi0TuUPyvN9pav7Vc0uBbdfVyZrExlqPJAgtPmZzM
1c+aaXnygDNNue3lvepVXWkoLCjQA72Wfhcd6aZagCsTv0D8ASAo6jYnUmVC
W6TJNd/fbCh12B0lD8NugAzLPDZyaygIghiLBsf7zD+R9zPTKBpArUToIrQP
iH6uFwkHjYQ2BYFdy6x43a2nPeMnn3dt9Yc0mXKoBiEzYHug/cf4g6ALUweM
ax4F1Br47iUjfwunTXNTZtsRJNb/sdXwLky9hIqaz03gmFtPOtzhFjogvtwJ
UOdDL6oQspZbJdd+Ucz8e83zAe6JBQl7M7w/nhxt5jmSXw/O5LgdtiA2Bild
ViZvBdlrjwyxPcJ+SZNpv/ytpMl+5DGH5DYC2OSgW2lPAFZkhfCB5bkX2gJH
Yz2axjRPe9ovT0owpi6IfvBL8IZnoVcRBGIwO3HIwJaffkiK0GkxtqZrwcQS
BwzYHS/jtlKBfUYHqAo9S6TchDdBvt3UzcweVwsI3oroo7GTDOsoy4ziq5Ga
ytVuq/6fI0T1ZCRSrMj551PzHZhbZI1csApM1jh4vhIdOw+V/Dv96VJNfbK6
/pwnpVcsTYY2cWnVp+6a48hT5ZBCeob3irNcFdtEzCH/+vszbj0wDs4x5BrQ
XnoiSgGU0sZPG/oxAwRH0H+fJ5Dp88xpQaBh3vaQI2vlYPJV1nvDE7tLaQk3
OVK15lDWr/ZpMjxlDBGCer2pW3r6Vcz62xboMobhWroXAT4J+XvNyzrcAHvP
2VC9AaPwdH2nwhJwvcZH9rd8bc0o+aLuek4FmTaufyhYyYVshagLTqAvKe8u
kEBTj/U/4eypWw31xSCvQM7NicDWH1i3dtRrTqFSJaPFdotvCKJJ8Vn9ebnS
D3iKN5PX2fmfFPqfgpuTkaW5P1RJawfpAm0sFKKwOqzIG0jB67SLBfAhpuBf
0tAa8nTAdowqxvpDrlGCgBxFZr0auk1FtutEjDhqLG7/QQ60rfG44ZfL3GMF
TzUd2zpFagxHk3X6TjddUzKCi32oDUcL5glBZ2QtlsNhb/RR4Iezi61BcsxE
VU7vPMkUiPHIbGSwyo/uF+DL3oB0PqtcpjIRKFaraK7WSNS+ihwi6UNPg/52
XOr0YFD8GU1yCc8gUfZOgD7Hc8/v8cwfFxoBbD5AfylbGjHIw2Pl8SMMmF8H
oT1f6Q188s//gWp/9S6lhv9CnURDgHdYLhCrjY9/sRnZCw2+Zt+aOH6YRi4/
746mvOH/m77398aUYHpTnKjQ2RtjTrbypcb7kO9TY73KpnzEGn5MFDoNrR2O
YyPhHWRCC5pSTXy9WuUbNjUqKslDkf31+pLJ3ypdk992SWkIWDCf8tLi7PXu
kKVvXVMEA/atYUhU0mnDO/Gt1nB3JNd7s7ReP3+DU7UupvCE/W6f3skNrpP0
dnaY7Vy7RWkym+9a5Wwtp6BJr7fGTR7bFUMgQ9ujANO6ND/uX4f/naFEmBON
dDczZiNu/k5NxOCzeUSfi+HQjP9Yhuklomo/8XY3ynAp9wVys8oNiIwIef72
Hurbk8JKQXKe0hkaHkK0q1JYzrUNHyxOdcKL7WYm3dVXrAKhrU40n/GnI0oM
HzbqRh/h4mIBlnrLP7+DxVJFTY3to3LR2A86tdAYc96lyJy71x6TMeCRYNmk
mgXXCteCRwEZGsx86kFvJqBl9SrU3SlaliCDg1XdpQOzxAy49c/zS2+HJv5I
0BgwiZV5h2vA4O5JbTqkn00afTUIGaxCXHn0srRv9m8Sk7YlrQmyHPIRsOGv
1NdPpihDNbPnuIy2mZkHHqIyWr3XmrNUNczg3F4lnWplxve52d3d/7oPj5n8
VKREBXD8LPpIb1syQT+Ip/CzZDqHdpTOggv1Dswur6x+2ggTFKnAcBnGAHKA
BuWLmiHnbWQUZiU3ztHeJFiD8F/7XTOTkIXVv3WneqTAZx757IhGq/ZOyXe2
gG3RaeFAzqmWHfNPd/BwsnMbGamCKV+vERQA/V0L+296ylTFcOajxw9KBP+S
BVcPygA+HiIcbwZa9XTDZiuOC77+nCsEVuAOA9wPdi0p6koqkij2OJyvKgzn
p31UlHlXoNS89TSWPHmIGtzeOnNSYDnKNMb+sXZuhXLUfEy4dupugYe0TGuM
Wdzulhxx094N5m28hNfs97kqT+Hg0VwIS5HbeTDTo39X1xw0plbKOtgymFWb
DKe/+fcpfVdIfUWfKRYeqxpxtoyU4CzysPCO2lyXbQvpPZJudF6q0wjKF7j9
M0eV8ZiafQkq9JDKu25RVQw30DFiMz2z01X0nu21ZYKJmrSYsgaS4kUrmtSJ
0zN/nO9JFEEjdxR/MkImstQGUlI+X9ZLd0YLFnAog190Gs+PPIFkuwtM2Uka
gZ+uo/G/yaWYlj65IvJTTbAXWa4KG5o+a6+DR8RrRF7QTbruJo+O0Vv2UE3F
vDkFDm1aW93FAQgLA+6rsfzz01Zju/716YLUEfCJaCDYWkw5JLU3aBh6CE3F
R/RWrga0zfGH0lAWHHGtsaelhBX99RugMWEz5+uccFZgkFOltchfDgThEUkT
rntZ4L101RX5iZAxLMBbAE0V2nKcmlGkYxUEynUt/nzXvzM9BA2LWYh3k27a
cOVNiubVH+KplmZs1dTJtR68CmeI26Dbolw5v/qlKMB1FhQdLxDRTHFCw8iH
aTuMAaU48260nhVhb0nLkVRz5hkAazfck5umq5cDcKjoYxBNLQEW+kLvic1k
WXaDZhJeiZGv1hicqPGnkt30GhMPS+Joza5VKd6p8H/ysJwPCzDG4j1Q5bQR
SAml+8BLKDrTLu70QZqUW9rGxma+uR8aw6SfnkvKFn/tv+Sg9I5VnO+hIUVO
vvFbHCAnETckYBqTbleaBwdu8pJSI3/sLuecP95f7HaetcbBiLzHHo4S6UN+
K315BHN32i9UXR7qYYXvFAbnnFHyH/ybPc9BQvp0VPXvpkOmZS/ugbeQIa6S
eRQATICcSOZs9sbe9kbQcFMIOrj10vNsStkliLEEdw854bs8tXts6oJfFkAZ
rfbtKz1CTTND7TPMXkpm5qNwYqDka9xTRanfNqF8Mc/BQMFo8P8XIX2rFTtv
JlhmpqAXGpQaCOOGzBY2n04eOwg2FeAAc74SXpKQjF0eRSLvTU6EtA751U04
5X3nvL9neWJoHfzAjuS41nShEnjmFkIKTzAIrwPlOuQgweLuWMhcJ9iLRajD
uxezwjoFj1UOUX0QX1RhdrMfKizyfDWt3qE8IDNpmQYq3mgmAkuUlH4iBwAG
r5mLpoGMyLcE/RQWscoAQUr591mSbOKaOjTDIyW2swmNKgUFFiLAMWUZ17yg
Qs8KLTM8HMA6O8NLEgsunzLOcpmXJPWujdAoBwHJDfWrRUcTS2Bf4EmAR1bp
SA1TLN+gAoK12n8Co4zgNKC1nbkx20fqcu9MDSrE0htCwGyHq05Dp+8v7vAT
bmc/rGR/UfNBiwR2B09OVcJ3U7bzwpXhuh4rwWLS+0qsjGYdnBzaGmySpK8h
ElY5lRwl+0S7vJ9UTBt7LUtpR0inZJw6JmwVPUCYR5NiImpmRFtSoDeeeOAM
54Io8wge5d3URpxo9trH6ut4l0CSIHPXGUMak6r70bV/CMZiwbSyF2Z6ZDJ5
uhm0EDAE6SiY758KWxeoI1jDgrR1y7hMgkCNzG2CyGYpBqD0bkQ9Xj3tbdYk
7ih+F0TQOuxO7/uQCLlmF3TfMZ0Fk7EbQlyUWPPgnZHeOzjL+052UTSKZdKh
LIsTekX9A0LMSBtkqHoB61nXpgRqcHEzrIktzWWp0FWU0z9XpF0lVz75wGtX
xSiC4qHHTBM/ZDXPAM1/Q8t5hTj8CDgZxDx9ePtPydmXcAI6hm4hnyqK2GzB
ZDnACERq5e36GJ32kNrTlZgwx2MHdHts7OPAfBn7jDhnRzjIx/xZ26EyavvG
10g2o7QT9N2kzGLt1bCCLCYpzg3P19Ulg2LzPkgSYfHJ9rBmGoXHCv8FAu+U
ItjgkRbJHvewvO4W6PFktdAOpNlBBosC7kMvg+NHfyGUSmtiFE00LznYO7EM
Bp/5qsTZdklv9cUTepCVNR/lHHMuiMU6rPGYj8ga5NUtedo41fYN5IyBXQcg
tXP48tj8PypWkXsLxiV296RJDkQgiLQaB/DLCvdTCYnE2fbDvM3MzyYCNXO7
X4pIgwdxhODoX4J0PHc0cKHdSeHnagRpVyd5o27qi5eFVZ4hsRWxKRnafOJZ
wwlZdCs/zU4SLCRDFXCv0vyyt8BOEgoSiEIwTiLTLZK9eTg+uo633s92bRZ8
68lAnj4qMR816p3/cnLcXMeK4bgkOl4HhCy4zQAI14B4c7xux3sHCIG/kl4b
XKArzw8/MQp0X2RaYY7agsHfg+lx3Q9eBQkeGdN3NuTY3WI+XGBja2NNyNar
UuPlKmc7B2a3CXbLuhUoZpLOgm8C5qr7gNSMubVxZquvgUEirPV87Evh9kn1
O0UEbG0CzCK5Y6P3MaBRzGmTGYNWV1MaV04pR7qrjKRRQmt6SVjIo6qqcxq9
u/FaxyUDNTBR3y+2vMait5UKk+h7XxSisbAN0fe4BJ2IhDwvilIpuDGkohO6
D/ok1qYet+z/F5Wb9fXwDWcmeRkK11zLZLyGW1005DuBlCgQz0pVv5klxHM8
xWt+SoXoz/+UiKyYk/NVGJ4Fl6QyrhDshOWM6S9vd4WpjMWOKpV2Ffn+mO4N
geL/ZjK9R3wyaOh3xHJU13eo2Y47n1eBISfc0JuH1W9YsBwLVT3XiXeka1oB
W9zWPcnuqxUAFi1gQqnW1ONKtPkdLKQpVCpQlhezt3lBtBBVdBCoUB4Z7BfR
YjIQAb0TMsICo8uXx0uVsaFAk1Ae7reYmMYzov2b72SWor8vm5q5c1XmCdhM
lRpdvFqAf/1wD+q9nuoy41kkmGqearamxIBt80YNbQC/GHxXqfG1lKgwq9/O
BqqWAPxPPVE31UxGZqsVDclEhedV0k2rSwaKlyA+aYRX2mLC+gl7czUdtOr5
+3TGYU6HITzCaBod9YSJJ27NcGHuSekdxcJfKfUjn31xhDlU38eBGPo6Pvzr
XDOTe089krfqFNwuGVAAelX24tYH1j+uAL7eNUS1uZ3NzV3nB3dwbIktbi6G
8BsEjz0UtmRLQSpNPGQ7qOxbFrNJUZEbrYMkAtc9inpChqffbpc6pByuEOIa
+JVTBXnBgBfvfJuVSoLoeukhQCIg3YjP9ujGjHEvyjFYbVsLbwv0Y6sl7fZc
rUu1H8vBgvmIh66K5unmYLotPRu5UaO8t5mf8yM+dMD0F3irW1Dy8911IQZv
Pg6sI/AF1bOg+Q8s49e4C3+lIEC7atEo2L0AfVci7kDnB2bJYaqJjb5q7E0B
k8auQYAHdUstmz3tBO04auztCdV8OkVJkv4ivBF93tgYgGp+WaBIBbXOFvY2
MvysVQ3Xi1I2d+CZb5jqNxiio9MUqEVWiDpABScWiwmNiJRyeS6JVESQzIfa
P/5LKp4qVspe2WPY4lIF9SS6dHUZ9dhBB+NeLYaRBzwR8BfpRmbZlvTfp897
gE8SP4tHCJAMNpVPENPmcPxKca8C0pX7OuUiIBWqs3VjUSS8mZBY3PSgTWQs
jw2Zq1SWFifR724QyS5z8mMK7RoS+UDFeFj6ep2qQl76lFuMPCHlq57dyJ5r
GIjgO15DUiLViT7eJi71NvNjSrOmxEfoN7W2fflV4Ybz6em8o1yYjEx1083H
LlzH1LQSkbNkErdEUziukDlpY0AQFhLga1hdrmmKg5kheDs3hdJ9ilsZeY4l
/3DKC3iHNYEsktsaOfTjg7EKxk4FZ5/wvvuxyELFEiF+qG9/HLuaRZ72q4V2
LZuC0vdicCl0APljextmf/aupb++YvxsZRODWNPyK4NfZfKveOVkqSHJFnk8
Abla9OMzDiEBKp8tC/qh5k0uOGJ6kZkrtC/ew8dNHaUig0KoRgxwTsCnWnJ7
qmUArSGQ9oZ62pQ+DktRSnU5MF8JHkvZd6oWvuDLJ1XaPTnT5jCLliE809YJ
SXc19cjGojRtIc880nTAQC4olieET4M3tFiRJDGvIDlyqwFRZRw/JquZfAgo
kYFEq4QOrU1QKsdV4Q1J0+iwlxTBtclm7mLqjac6SLYse4vyRDBEYljRuXD9
PgI7MCHwjtS+Hr53P008eryMrrvmmWvrf8tlzgvlkAuYIV7SciY5FwjIcCYL
a5ROw4G+WTCobD2uVaL7g0on+JDmIGT49dcbB8Tr9tWagMe8jynObr7hvYmJ
J7aKd17N1303q4MDNbwaaGw7pzp429UOvgYAlN2/CNRz+bHWTQnf/1KCZBt3
fL179gG2W60gFLn2yAy8L9v1tJ9k9ylX5Sbs0qTZ4nUrfqpEXg7V85hDX1Lu
yYz44SR4keLVN014BZoSGa1OMOdlKSsdrMIjpDTTd6UVF5m5BvhC05VzMTj0
Ik2GreE9jy/zF34H8tRAkX6iUOVHE76U83zrt+EQvNTl/qXiWeTacC+/gZEC
A3TI8tRYyKAXkc4RjvZ0Pla9dza0p0SoJdQNPeDPgOOSYWazj4A9Vm2BPUW/
0x++rHk4zOmLynlzHm7QBQY+KZBrzAlufwRgUqJ8wqXqu8Vi6qvW0xEg7eTU
Y+dnrPU826lGDlcaQuFquLnHr9uyj28n6kHpiUtp38/S2uD1KjXqV3mxsqCS
kGOZ3xfakVZ75vcnbrGlglj+f+ZdnXUPsd3wQBR2a107DgR8mT5E8hTKAhI0
f6WHWCsiVXH5tvk8D6dcpnnnd2NeXLT6anMlZUOid4WgzLQCBT+ZA1jV9jV3
N+Ch1DvZ+9HXFn8FvDgCjOForUqr0pZyYFV9gvClzf4iLtqnNQo/cJiCTa2N
+abAsF4fKbeygQ+hxpWULPuqWdpg89XpCwbp+h5bmOf2OM6KEQoVJwI/4Ptx
ZYlrtUbTYc7e38ZuN1lk9lLZ4K7znE+xoenTMqjNbjnJXG/cxeiNM8rppkiS
WIM/n9qK9vEXPzi37tOXmMGafSZRNYnYx5pyex8HxJkii/Qk7n+MQSYzrZbk
WkNm2V+FyKNj7cwMa1QAaeBv+3uAPZbkRUvORboZ1zyqGJ8j1jx9Tnj2EVjb
jwrACMcS2kXDaY5I7QvaUa83bmQ1p8pgUy66HJ/gD3fKi7u4YyYoNR+pn7OC
YwcQD1B802dBJxijXkuEjib+K6ZWQ8UkYG0IstAWcS4Pwpyg8SFU0xEBtl+h
uxxZHqDdGvVqwBl06ufpq1AkKMU5Kv+U8wZtv//eMqqC8Rml3uCFFZKJe/KA
WynEfMTehpqU4Q1ynOG5gbQ420QUZi/uTrgYUsszEHa5GInKcVl+dDB/lPxd
Hf8d2YfLBjJECjezTNR0HVfBttjUF38TS9DqLuFbgIGFR8Mq50R4XfHbQca7
Ta1n2qNn2UI4DfWpBMYmIgudbS/mkAO+eKsWxwXbWFCJovv1Tv3NGsmrm0qi
ecnMTbYtJ6ujirydFaFBVarAW9enRGVel6r/omKKIKDSQbHnrarFq+cIRfZ7
EZ+Lnmvc+FrHj7NjRyZQZvRZFTKpzmyYxh/itUrks0jV3w7z3V3mzgADGTpT
oGePBGXbm8FCMg/9UuOIo2PcChhMTDCiJBdqBcDM15DDRebX/u9YO4jL/uw/
bWMCTDS1oKtjUY0K5+Smu7yKqdIcdKqWAFjKN83gU++lwDDv7Rlq0UH89clt
0gJ3D/ZWS4U288p6gZTHPmN8v4h5qa7GONZMURdKbCg2A2PftIoLrdMJVI/I
usZsHdTkOcnDEAbRIz7D46t6qO8oY+olyNNInr8vmWg5Hr27D9XCqSHFZsPf
ZlpTrGgDNkQT13gnzJPI2facspB7ncsTdPg2LjM596DCgwPVKJtKPdQCvfP7
yfYSXEqjyfJzki4WCtDys+YVWGMuWOXjBIBFyfWABoEbkx3r5kWSFFe/GsY5
y+4uoFKtFeZzyYe8o8lVaHzxDQiOccZ4iWjaQDSPNizFUc4vgT+HBzmd9DkI
xMSpMGrRXAPtpR+OIy4j0V1LEEQ98QSIdpYm4Xc7e7eVT0P2NtkR0/JIT2Rb
GV7FGxI2qX5K4ZqAwlnHnb7OTs/g3x7t7OhoZ6Aw7JV7psrHmFy2XYrdbgbB
oicRIhYTXt1sDC2KlHeTVND+3Wj7TkMbGoe7VcaYrItl1H4Y1JIfKI+yM6ps
RipR14u+WwFlK4q8P0pGtLA5TxcnJ7ZRPMEk0F7w6P+mhu33+qLpc3aEUy3M
7/teGLBGg89Jm78HmNFvg8UdbtopIYJL4otKrqRvZxggRHOm6DC12wP9GlUX
UBy3ZSKY8wd6gPR5494YA8LgUithX3WlTfxevivYzzaDfCmUL105CkeUtbCA
7FFWbjhZ9vsHonSXgNI+XphBvXIMsMQTpulb9excRCFbMI4rKpEDD0XiJ6T3
rWP5MARSmubd6IDfwNMBOXPfVHT2Xo0ZhnaHPutCv5qdH9wdUprEE/X+89Rk
gF7XHH1jva5tchT9reulRLrw3MtZ3cCaNU97kgnE1VIcti1BeD4uczc/cTDB
g0rK6XFE1BgMPQXJm/dPUHA3jEKgRGiPp2P9ZnsNbIJWusRgozjzHX2zzDFW
bupBJvLN7K1PEjFeeuhqHkUCmI9gnX6NwGltrtKHAkfxtBQlLQTg0oT1G0Bc
PoyT/enG40KauXhe82mSwWMwhfDGeZEzyC2mk8ZflaIWXuznGyqjn7CbRunB
KR1v9cJZAX1jXF9vJ2piwxD3Q1tC58dbfW0evOsQvIrRhlF/G8WvHbDueI4x
m5ahvKc5hoYGxHWYJ865fK8IzwiuT/RFcTTxp4L1rMfCY3tTj9n3UdlWm9y/
zldR85p3EmJC2bxo4/FujndQiISyLwAO6OxLcBMZwGc6CZFD3ihYo5mAYlZt
poYABUBTcaa/GhnairW9cfvlYerPhHay6PFWhzXVyfVMEAifYB/cw4K87w4Z
B4hvXVzOC0JD5JJjtPLRt3xhgr/WnrAn2UADOBKVJwyWGHBDwO8zgrK6Ug6z
UQ/Y7MVboKyzuCSLy/vQy8b3CEvL8w1hms7bFXyEO8YGUZFjRa4UM8jKESC7
v+FQlibN+/eXByRAYgfoEDLDE/QlLTxjTHh11+oV6SQCZd+79ulX672a8p9D
relGy5beTX7zxYUMroty/wt2m/sst8xMDH8SwssbVCa4NJrIQxJdywpvUByP
VEzTx7Jp9NLwSrj0gPHmeWGBak9iZmyrsl9f/60PVWTnzRGVx0+DZWTb0cbN
dKsgY0gD9hpB6gj5Pd1yw+6qhqIiFYQRup8ffa/VdEv882ajFqvP3gYeKdbk
18zNV7KkApbj3T9uvJNOu0Dtf6BZ49SQgzChKO626sGYl/oACDzcwM12cV5b
0ta3cJDtpJqxJrHqYgsYq9Li/N/rdhuPBinlYnk8eJvY6UVYJIzdPedb1zfp
w9F+XLmP5tHVhAXbV920/o9Np7Z7j44CTWhcH7QPsmBxbfyvoULsNsuHkJGh
TKMycvSxOVnW3MHh5SnsWB5AyxWtseSWJ2KqMwly2gSDMYnnS/Nu07DHwVu/
sfrZCDCcf4bV5TiDQ9sIJQfAf57ifQsYpf+WSCBe4bOwJxUWPzkNZ5k+Z72j
xzO1ITCxVzXODTF/Y8ZReE/ZNNo3y/R9URK5esnwMZylQ9NAJZTq11EuIes/
2sRU5knorh59a5eksfKqwb0LU+toxGde7+MDxs18QOQPXxl3UuWWBljEqz0x
6skt4ftXZhS36FaJgRRqi9hQgVClBZ1l9Mco6s36xlO4rpp/yH6b/nVAfR26
QkM1NCm57EjRL4YHS7jdsbFbow2LyZrEEoImAJvGFxCs6vAhbGE4Thhzbkfs
wvLc+K5eK3LcXRkCSfsZv/V69IrDqAddSm1ROjXaMeGYwBTiJEpv36GPO37N
YD21HKQmcqTuu7se4SYQkp29CLlOdJP7Deo47Z8FS9II0kwShFTdO8h3NEYC
OV5uJvP0yna2wz+658cGhDFZVNJt0CwqJYOOdspNMD6P4sx8Vv1MQlyZHAjf
h7MrIqHeFcCZcxNxKhRUQmAN/5GGw6xKAqBXy2cg2mMfnkWk18TWXgtJa2PZ
Spoq5aULCq4LieU3tAuyjzPKKoSVhuCVruGnZPy2K6uOSNZsZqFAmZQdQHm8
pTXlR7nxcuyKyJZUOEDJr0uMxZWZGnlRjBi8J0M3sQJ2WD3NWOXz3IMifBJc
dY7UMyR/YfjuaRbErT3NvetG2sW52/PXDm3udYDJ2WQkZ5hyPqUS+G76m90d
FwKPF1PajNiFcdmGjKZr6Ba10z+NRdNYdlPgkzaeV88Qo+k3TxyHWqBXWY7P
cxCbLBCJm9bMaHzk5lgWrOfHrUWQILiLEJODWedtmOXbEyMXbMTT/8aP6afP
uF3QQDRlGyrK7YvSWDXYBW6DXBpxsN9vgkX4jyIIgwwJmCZaUkfCb0WDq25h
9DevzCEKpNaYMs5aMnDJoPAX8QoVsK25pYBug+Zt2C33GhIRuKyq06F/dBMJ
orcOPyrCZs+CKOnwOuKokN9+JZBoh25EkzYp+lu2Vbk60euc7+ZXUQtmnsk+
Kgvfldmu7c+jketh2OP3F3xZzgo1UYxN4N6aGeNvJGLYHtsjrJa5iGd3Fh1M
8VJuY8kPlt6CYaNq2m9xlQ+yLnSgOs/a71G71ZZ6VTzVC/StGZDeCHIQWLYO
R6B3V2hVEeNs3SvYbKMAUmiHgrATF6zAkyceblsigcDhLnBt3KifeKsVBRD+
YAQF8ek64k3QhlZQVQXfal2zu7MIfsTiTxxGjr//1RR2ij1tUpJTeYEv9/sU
86pEdmbnnT7QhIHBftPfe6ZtcJnlYPfZlCyzEcZiIW8oq5uS9p+mk1TvbqIm
qCDZ/t+BI/yt3WSOr4NtQoX1Hhj0aY43AVeP6MJWfClZojbW6Twt93kUYG94
Cki2j8/IFanZegb7KyBhfo7UO9qsccIi/FTJUlAQmcqCL1NaqxRA53NvPE1g
KVVLWPtiBpi45zNmWxLqs+LWr9GlBMQt+ajHaSO8DtqWLSckcbZYqDwm9P18
w0txTuYjE4VLGP/W+NHGRwHb7IdX/0az3sd3EOFTyZvwfa4r/rmqgkTY+wZq
Qq/meIYOwQtPEsoFz2vrS/WjBYJpUoItmvXgiKHMGJQTHtLe0HbMF/VwPWVI
xL52XRx7TsnKdOhI3+/UtHgClGJs0gZncATbMN0uHkCESpj9AGL4NseVxZti
TofVHCDve1+DgiMNLAErKJhQffLL9vsKlE1Jubf6NSG6mYZrqPztRRU/zV4W
0zOOxiBippnYIgTIwgZ6suc3+XY5uzwecm0c9nCoJUZxe2uo/NCTeEvUf8R1
ePFha1wAkobz74zmRaOGlL7ViSoWfLKlEE8JA0esOiePAprpA/UaKNiGTWjr
wsFIGLku9e1FoacUiZLaQxjr5J9cmP+hisQSuskl0UVkhrxmI8vHnM4iz4Pz
fhDnNyZBqdg/B+PoaSA4pp9lElV2T/ZUh1z3VBuN1e+pJOY+L8qqglsqU22G
zcTo5rNktd07G1sXnX7tDvaYrLK1IbW8w2XPKnrOEN5FOF19lkEzT1iwl/Ew
c6H/fEDzT4D2MpNviJ4CI9B2KwaBrIGCFk7HyHz3Zx2XXYiabU795HyYF1kD
3D7dkcuYf/PPtQkkgrH7ByKtsUxgtcAME7Zj9zsCj3KWI/dajwHYK7OE/T24
a0/cw7PPY96E2xfRJhZulCY+IraueLVR3onP4CeDjU+xUhXMY2KfhnP0ptJW
q9hyVXkqOpSUNKqB5DFa3zITOczasyyf5O7n/3kpuMPMxdH7kg3fTYTlmXzL
/f0nZStOTRH5Ej+xzBRXAkpVZhmzD5i9mISteqyEZdFohEBM9IKjZKCNxSl7
I+7oXpEmGox0UClQGb1dvjilmWyhqafTtUre+pQXOYHe6uAXf6jK0r89gkL3
0+1O7ZCX+1RkTfkF8BfILbualkQ6jGHm3d/QxefQPf86GvcV3rlkZAqQi+85
KDrDDxijRezmzh4GfNgu6x8MKZxat1FqVxkKc9qdpkr0GAtwFM6K+lChxgLv
dfvYPwMDqv/ZXeojy1+YAMvsBbYpIYwekvTONXZTvMpGRhTJfI8YlyExn1CI
hhR4emPcxAh2NdjOV03wCJ8/50W5FMgLsZRiUmlYD0KOS+953k0wxdTso25T
At2IwO2SPncRUw95XB+xFQfshq6l/Z4vr33l62n7Pp+gHY0OyvflFryex+f5
MwY3502SzaUzpiIWneEbkRtKuDBVDI6PV1Xp13gzpQ3s1u5JtUD+Wuu8hm4R
KOYgowewScsqBmCv4dU/ty3rctZwXMN463t88RBmE4MpZHOMW7bHN2uWtTZ1
mZzmqlIGc1Oxa6FFZtimruSb589i9A+HaklS/kFK+bgYLkYPgw9/BU9VS8bk
9hYPEfLiKPlagBTfNPcUZpC2tTl3bqm70ziUsYtq3BkI/20H4iluK46EIaBp
yPoDr5d/Znl/qXge1g6ppEFoaBOW42pggJ3IVNeVEhh8CiXTaiQV1YBt6O8N
mXcNOtwousKtmYoWK7DKATlkvUekJud3VsCoNuksKYCxj2Dzdx2xjI18ytBN
yis3Oh3khTlOo+sSrslaY/kLwK3OOQXMitfQT2L37caEH3sTwxcKkHHRjmLU
hT277sdH9A0T4XpR+qKoDRpQqmuRgttq0GGKpeB5s4EzLXbAy78Ml7pfM6qd
xfyOowE9n/AOsWWGMS64L17GAmTHBZVgczRcUhmL38kHXvwApnSeIPiMBBuX
XZ2nzOexUDP71fxymamGsluYZPhyzhmiPx99RBiqT4s/8rDE8Y4VSGRRUM+F
Wd6vD6DXaTWjq3xu9ezaENHJREEfyoVEKNjn84KvL5YcOSJuu+l3s4cdgSdL
WppmpJWEWrHKCgrfNN1TfRCDKKofABUoBK+tHv+6YXSZOWQeCH6cABsx1S20
OPMh/Fd6OGGRJMuyICfpgrwz2BOEcHy0QvbD/4whfyZXKDjpugTji16U2/GL
5B6QpAJCaYi63jrED5iaAHjQXgrVQ4EZkymrfSopWbW8R4m22cl7W8XCaxdX
Xt3f/D9/+q/oWODCWVR5jGUSn4OE5zMILj0cw+760YeVzvqad/VWW/asbK9I
NnhM2bhA0TdCcgf7VXwZ15uP+krOA9tQvz2yQh8K7yw1S4ymWN1NSpkmZi7w
iiqd9O6/bL9FG3+huPW0AOwSwiOJtJfRZnYbM8UGYN+z+CdfC8d1D16HQwu0
2FLxPZf/jCX0/sSaIqhe9I3pGj8pxhhwnO/FRUlVm8vcB6QODxgUoilBBJd4
lVyJdESOTPD4WxEXDnl0H+LPHBGVAH9gP10aBmY5i1sfSbIfuqepB6tDXrur
Fx39AxXWe1ic8Rpw5KvUWRJRAIuFCuBZ025yNBxwbfPQFWgSrzUySm/gNWmI
9z8DN2HeR0YV1ktbeZAviVtfowpiGMMtQ4HCwuKGdjB9S8AGF0zEq1EiElrt
VgjXcEy/JLh6dAnfo76egaY/0dJ6pY+VgcMxdPTGj/IIibJih8H26NT2lNNl
X0dCCwuR4rSDVENnfX3jCug0ouDEtHgSqgH06RBnGB4fn12uegsMB626KwJF
Al6YDqNbdUnM5/6fAbN0a412QfrBenlQFcNCh8xkCsHLLp8BNk3BEdVJfgWM
NBtfinl/BCCS1AkVmX8LJQNGUDQdC9MR33y6Knol1NhtlYy56lLHH4WECYJi
gIh2CRKe4B0ubr0Jt5ngc/t4toMVP50801ntm6tWcsLblvXGw392GoniWs23
4OFP5jDmubJ7t2d6zrMLr48jhOkVBPeDaFbmWkHEW3FrPwZuc8wBhwiZIPAr
KN0hpkJNzM4/6ZKiG/Pm7AaNnMWPZve99+Im0q53geoiDI78JhYg+EMLiBXf
EZQm2VxHGomhZ0fekAMBZ5eHqDAKfvXzSUAq+KVO46myeQ4T4lnJcCB7zzWh
nkaCu6Bof+QP1+iKopd8f24ylnhtTkDsDTXUobKM3C26P8hCA+/K42hAs0VV
g9sKboGYp1BO2vPlwuwQtHilc/IAnbFsBND4UyBVVVTc1m9ojRMmDhqUWLpv
X4gJlhqMNg4sTAp28S4MMHQAcoYoW3odbpY9XBoVgT7xydqVEvJnu6mMMMP1
S+IrvXmofJ3EXhBe7pNyWbfrpp8br/MLw9t3SV+tbZGoOrhWR2GIVABsMQ6w
cabgJud6+nTcbZ9p8XddssEhdWB18VCZ95dxQ5YCwjX5zgtPFxvaMUbRFFid
kt4w3B9ogRDUJQH2Sq2qYNuCTXZqVuZxn6wnOWWcMlm5Mfhx9hopI1gkHTVi
tMfTV8sgHJg7mpqtWNYlu83mAUm8utPAT9ztGbj5hx6M0fWw+XvrrE5Tljww
jycE8ebihAkTWjKlKPMqZ7M4wo6m7YZj+r+DdS4uwCIg6BHvyXCUTGHzYX5e
PFufkGduIgJ1bOQsINdSCm7acfkmnT3l9ehvsgLZwX8K1WkEY0sIu3NqOMxT
6kUtTIt44ARR1AYki0/bsp84Dr9VNNcqRPV+0SG+mySrpQ5v2sQsJNISM4zM
WMoyrC0gWsvkrCOue8nUc4G0W2zfy40xwbiFFd+Jl10jJ4rxn4GFsQuTkNFy
7yCfeqsayifWGtaFSFQX8jn6/pX1dFHUg5LVCf8zgX7Ms4YQG/uk7SBDLSuW
jhvlQytVXp3Xq8BB1j3vctZP+63RAnK3geaVmwTXGc3a1/4PgAh2bE7aJcAr
/jx/rJ1RcSyRBAlYccm6ZCIgSRiIjwBPiBrdMy5r+Jhd2ljr6nhAvMTAlaGW
YMQ0xVqRbGtqIgpJrOABEMQJ/zt0qVRsVlE+RLfJ/r/IgRb84C4BZZyHmdVC
OmY3EMHI5Ip9IwUgUIkID4EBJDTM73tiM1OqNMR8U2y6pgEznI1eyf/dzN6D
oBwUooD5x3RXPuq9536uF7py6Z75Ngb52B7FoHaLTP/H2noeCrwM6WcgkWdc
gHr1Lld+isnYovs25kRLCIXN4jUKeEwqMa+8ltCE1N9mQI/oSj9hqUTitB1k
r6lrhacinGrIH7CaoZHtoTZkePrVYRgt+koQeKGc4ctiwCeBsATQCrkB039X
vMJ25ityIL541OMQLXjWX9IzwAioIdU2to0L1n/Pfc3GU/NIijcQ4vS4rY29
koDfWRHnWHmFMlEku8p6OF4mMZY3c9wO72m86QfWC2p5zgNVem/nASUaUfQ3
ri4CXSe+ShDNcmVIA9y2hpsfhsEpTM5fNyG/HdF7pL9UHeUqXsBVc7LNX9N0
qRIqKn/PFhHRjJaQG+ozETu47m8i+RAS+4I8ijW5zvxdE0LwnybShTBE3unj
mSmgyRuFFnU7DL2oSkiEgmf5MGtKSpeEBaK4g8opg7mRVToQ9S+zuOAaRFBb
c982MKi4QZSQEklk9y1fIRwHcLNMmIuEe9IQvceWQhp8A7HJDCK5xsVfajr2
f2iuwWt2/3ouxzCM9TCdJazhempRhKsunctw/CF9CJwCrbes+Ddx6RLJrT/m
2WkVNY/i8EnU0t4Dxqc7Lydyz/yL/m8r+N6AqAhbWMBQozfsQpEZfMz6rQ+a
W+PpWspMlVT0k6JjuKR6RyOappH24hCJbZ4z7xGz7Cszu9vdc2lUxH31tcvS
thfAbhgQHwrqb0T6EpDGYqxVcCtIkPgri1379pM4+WapL2Xyyk5D4K1YH/eo
MFrlzzt8p1viXTwhZfiYWJls377keQbk4n+aTmE8B0iuXx2FaZgdAQPIDxyX
KEmp31NbwD4GpE/xwQ5VoEgL8zybm0Bbn7qURc2DZU8kdvZQZ8Qq2Br6jyp0
yEx7pCIGzNCnT64RpCrooM3tSq5sNYNkBZRaJ8IYIBBMIJbdyJ5KbjnEs703
9WUf47dTFgtrFxWRVbVpFB8XtQf0fK+RRHuJVmukIOl73NByoTVIrbhCN02I
DfiPSFolN8KUdbkljH5JfR5uQA6OjEAcH/4CoU/ee5TOR7eztfkBLTbWpJLi
gytemPPd8m7sNKyhCn7lxGhywdBInPrfIKcthJznKqW8VTlJ4q2cPUYak3yD
n2GtrFsD0HQPwiRjGNRN48E60WdyHFDY1tkDFIl3MUETW9Z73kAlsxUrR8HK
dfBXclCdKofY9Hq9hqVoYdO+ZNy1TKZsr2+tftzZJbncRxD2oM5ylJkoMqjs
LQe3XcLdKsPQX3ggADzo9BcDB0Z5tiag+MExPG5hiMQkx3SJtCZHplIYVeBl
TQs3tKKl9Cs9FGl9sw9DwJrjHykagA4exSMXxeoJwI4nZvwcihNM8NwKIWFf
B2QjX11jqnlEvU5cD32loF0+9impOT1TDdwkXb7Uvgo2Ot8GyXkmVX4ZYJHH
p41tCNYNJLs1XkA94a/e/yAh9059NRsXXX+s9h+3QBVxWw8+joQUocYCh99/
+W6QUv9+gOxyWrZ0Y0QVEzXYWmS7huRDN2tSP2lvI0ODUa6HlwLw93lGG9YW
azuFFgEhXzwUq4MBv2siOkHL0RAx82Kf6ApxjxiV1BWs4gOIlARlwINYRq+w
Vb94j6qASzVZmxfum5UEL0Hyh6x1SmOzjloca6DJbZ+RSEJj4O7R0kWnchn0
XYd9OzB/RERa0nGNYfHjYnVBzTP1zXCq5tRkYBplvqnEVELnx2KrY4/N70zF
f7RbnOpMQOisq97PSDk80a0ql7PM+bjbgYc6qJwxHdHBUBDNExt3slvRR8K6
AYr10ZE0Rcka7NQF9FlGfAdYBr5Ei5qj0K6BHn4i608qkgtJHNpVjLstwEMb
8bVCGmKfLLVYYvowz2zrAd6hBDgwnEfY3uw4a1yIDnx11byVncjHYVimvAoe
szg1P5vv/9PGcjny8HqQYB/dLLjWPk9QUJdZMhTuwXTzS/tEPbWSpChsz5HT
TXJSleeG7Zmq+wVNhtcflEd7CE7rw53Fjnt2U4q+e/sXGFh78fyPYMI3mM20
tzfThD0dYePXf9OdvIhF6XpzGDYrp6ppoASgTLQStsbuqjxtiEfPJuye7WqR
cVod4h7BkMPwmyDeBARmMxNyxY9vmKKd7MKvs+W9bM/wsQ0OijurUoySDlYp
dn3hZ/Dl6yOLmR2xOyNGoIsmH4t5WFGbMFMf9zM9Kkjw5pRFULgX28J2Zt4L
kYemBFpSwKbpgBRpWaFaMpFqiYwovljeZlmrby6yrOxlPpXtXrbtDd5U0T6N
gctJLidRnDYG1fR0B5sEmF9TQypT4rOzHc8OYyCy2N1KjU0RG13G2cWTLtJU
ifuDXfdabGJ/GIZ9TJHvHjDoOa9ejDw1PCXRBiLu7sLIKXGRgBT0654vkKpN
SCtB7luthbAhToa8y2T4GbCHHGmkEeOGU63UdC0Wkh3vZuvgbSP/iaU36B43
9zRnWOvF9TQ5Qe5Ps5HKGIJgfH+bCpmKljKREkMZNIzWr7ObBrJGXk8/U0N7
2yiP78IwaEeZaboghaoqmOH9hnCfTAjYAvq8ppiMhha/zufkudG2/nSRbaan
KHPS/1EoiXZmv5IRXR1psw4GS5ISZllwmXH3fsALbRUc+abTgqESfZo9JvnQ
TNF85+EHAt+zsljZrP64CS3G8OHOma53Xzf5ACOajmUATdF/zLrOtQ+SKin0
LNMCgewJtZxcU5rhxhQw4K9pEcKToq/fgNE/DUy5d0r1ySZIUbM9K8bacGQx
q4W2n5GpbeKdCVjngfSob6wnRGuu/tjn3Pv/dIiStcBRerbGgOjEn90fJLGR
pX1FV0AmVJkHzSmaWYIk9ArX8KZ8zY5aErODo8eIulEYPFBaDomeUtkvVQHY
GVBESkB6gkEjsQqq6AyiUqLrTobunIjzZ4CNpFU9IL/2LOzaw75HU+YqDMWn
Fcj8TC0fPK6R/zAovT8aEq8wXH6tWG6NlGicM4dV1ObRQ3JZOD7SVOr9J5T6
n8G9cX6y70bhZZ0dVrldyisnryI/O2o4otBIm7DShxbopyoSnDy9OVp6B9KE
FTyi7lfrVUKKNt2ZOidSydJvkxmjPMNN84MwM54KLBCXurXMagNaZH7HJL+Y
Il0vrT4wBw7aSweO/rv84bZvSHGscJNPUHIjvIfTh5hRGcnQBOUv0Dj/TgMk
zQLLvmD4Scl21kWPmTX18/gBXc7pIVuudCMSvvVdcgCXEIxHBSkDLo24I9yZ
8rA54VTtWsAzICMw9OTkTVRLyXF/4WNmFPQRlqvoy5kevG73n7cgFbZnKOcB
RDeh9/ggtOvchj8fSxocIVAe6TqlUAi0Gbpe2f1csaQ36MeLR+jF3JRbO1JJ
Gpc0Vi0/qBlg6d9RiUM5u8dugtFlx4oTPoQq7VzEvMT4oabCuORy9kkQsOkz
R0GLwCowPFNh+aUUXyz/L58r8K41Us8av/5Uc4WFn9vBWy8M4wdxlnWwnK58
Lhy14NlXROmseNAB1F/1z88ZypE7FoNrE8yr0o4UjtulNpuBzNXGty8Piigy
VWDTkWkFOt0bDi8yS0Vv05zA30sazIf0RgrbZ891vQkChlkDkMnZqGP2y8zY
U7L2X3ZuIW8H/RRnI5ClAt8RR9Lq4kt8RQ6Ii2HrqYScvshdDlIoQ8RoA+nE
eoRZNBGDBBUha/FO4HgzagdwAoDfm3PzQ4anWCaXNak4M6J4cYzfdAhLHgwk
yWvWdRKOoMbf+rvIP6RIRC+X8kWohkZXS2TATMn83TKIZfqIDxVfRCPD4HdF
p0ECn/Re5AZGZ7/pRCc9Glw5HdhjnG7DiiuAwkTlAgEW9kDb/Qbr+bcTvWii
zukE88NaaqFnmccswmRcJE/34d6Mfqa6S5NJkASeqOqlebcPQ2u1nEevbYW1
3rTTbQ0LVyCbmLL5vgB/okY89A5kHYFOqOy1kV4SfvmPZx736Ts3qFHSOOJO
ak9GX69Av4AtgavgvApky2MEq3FkCaaAfkjiyO5x5co4xXUESa21ZsnvMlIS
F5yickacPB1DOzDqhUZ9Tuxts2HWs1qennmCJtXNYTc80p804jLsNI0/yaFc
MpN/QtetOCH7+6MTYEGbFqwebGBuaAr9ZqZQJgSxRLnI4OjVhyNA86oyR+Fs
okOT98yZpQuX7csWHZW7JVcQ7P2xorNDOxonQyx9TgUscGXLmz/8nYq/i8fl
yRxvvUT3ldEYsj0Qd7KUwQ8VUgH5qFNaOUgvKyx3xJ4QjtFpV5u0qm0MoqRG
rlxKQ5+Mn3CuqtK8hgOnrbrJeUI1BD4awvBGQdxKsAchBtCPYoj7Rp+ADO0l
0Gpaa4Kdn991Css4xypCwcRW08c778aTfkewAkCkS86E9vIfAKfFfTFaHCkF
39t72V2dqd5INIIJbGWgoH7zQhTjZzmVkRCb+sQsQ9KxqxfWEbNavfN5O1JD
K1khHdsc96XnIcAsAyBDq75+T6HgmB9MlUzcPzOCrT7fNJ2LDgUQTG5WNYvm
d7XMViAuReZub8eD/4BVlrBPiqS7SgwWT7G094vOgUKiDNSyELQc13Du7NCo
Uj8UkAblCSTPMCaNk/yiomFLCqrv19mfSi2NXgKTjW+dtTSvDFTF46LrdaxF
MeEKTSINZIlLZeLlz/pyVuBaRXXrtgGz4mKezrRMyb6k9stsLlwyOPRVcdie
Xj61DxFze4Z1fMxRuUSlYrSbYvKRdOPJ+sgzXQUlyQh344/JRG4b/oSFBaIY
MqoRk8MO0Ztw7msfxXRTS+Cvsliy0ZUfbEYskA89b1iaCJk+YOSSFe1VdPLD
nsbOxEcL7JUUHquaz4ucY7HwbdMSWyVcDIm1DGwqvv7I2xhDoh8uIKGCSrfY
EPcmlQsum1fqO6Yr17Qz97sDyObdA/oiUzUWSOC/2RbfvwD2Et0jvlQXZgXD
RS6HHn1shKdDr13V6p5WCAQIMra0ANzYPQiGFIgLlmESTWeWzoWKV6D42Whl
mtA+N7aisRs3FYgc2VV8SFRHkfsFm1CM7m0WozVva1ZepVWU7J6cMRtTMY9W
CiXAyvhwYh3rvV6boWuopF1Ipqorn7EfU7LK4EuPNYnEkG4ngXtS6ynvnj9q
0D2OA6nH1ToFUJWDsWE6PMWrAwcT6T0QG4BCpOcpmQUl0C+gIYPvCRqwmQHH
z7pgefdSAUu/dj3jQm+Q8WdegKRL9s5f3QgYX1Yq3NKMZtWwDkEaeCG/Zba9
bSDZ+msCbayXJCMjYGW+l1ltB7Qt5hAkJ31jHUymho8J43cRs3c4UgXtUDex
t/ryCK1fDXzYkXIk8tBE3UNkXEPSwu9rdlOzIYW6mTocsaeRcM47kf7OVO1R
LIzCcXPdvnsVtb1cIjA/Ah0X+OzEXGP37YJoe96LPfPeJzxQoUHf7QAVyiRx
m/eyYnwf+4VbaM4wlr846J+n6lDPKNeVyd6M+BWe2yewEww9i5+qlQJkW4SD
PiJtK5O+mWhcyY+DLNTuQ3YV87n68sw7LOdQa4qbFrIHA/CHpkvpt8gd75YJ
399k3o4h7938g/c4cDWKbPdMyzWmvtYyjxyPIDWTe18IkT3QsdiqTmHqervu
NbcWCBbaEiHLSJVpFbqYV4hz8bkvJSG0Q+sU8ctEmUQeZbBF3hsRjkWN0LfT
oNlvq1HYGyTzBS0s7mw5LzJwc1IXpwpyC7J8n1RCpWX83yXVcHrYBmeCwK64
xM3a8O7VcY4105dJJQVO1PldtxQMqfh/p5Af/ioHoMbk2l5GxuIapsY8bufY
pyuZycJBZRDVXUwXckJgQaHl1DBtRfswv6uMBkF1nTG8rL/NKtxb/1bnyYp5
Hv6+9jtkNsD4OXiZUQb5mGYQnrIoKuOvysD94n3iXE5z2ejJHxCIrobYmYVl
nllLsMrR0QD6PQYbYW56AtB7lrjOPe8JJwO/N7yaWLN43DuIIYImnDUvMJQW
/Na7Vr6QACywEL3dNGzdmUQrjxxBcyC9ZvwFxxFGe2y2SpxnP2G0k/GYdDvt
DXJrSpvaykO0KF2rnCgx2GneEb0rQmU88H7PG27+GSiCKB7YWZBRT1jHP/31
CMZC2KvbJDj4Ftyd08aettLS2/1E1A4+ssP/NQSYuQjYM05IeXsFYmiZr51W
7sWYcof3hoRydTBxp5D13Hm9fFQtr8PQhH+cTPf+QHW6a4GSlkFmOFKWmDmk
tUq1fAXNLe8DdO8IXGQsinMaSx5Etiw2EUsvr8Ki6JkYasz5MatSqZzdt9ac
O97s+I85dNi85YRiUIuOgczHBrggsJESqlTxivK6gnJv4nVdANMIb4e9isfJ
7CglL4FmIPWkt7vQcvM/S9OwQY81ay+wmbCu+Jr+0TPNTgKbchN8/hyvcnx6
nJuIKzOKiI/JqEz71peqkssVeoS0NIjEF2oPRsWU5n4JRJTKLnioLRB91qFv
6NXAR3oYiK+cXyfkMM7Bz7AE/Dd3HdHrkOoIs0S/X+9i6Iob79GMrDVSdET6
mlOnFcUjCZmWKeJ8MMWeAoxMz8N7IT/Lq5N6rW7TRye5Vu6Yn8ZIgraC4CFe
R/9eSVmqxgXOMhaXuHJYdUcK51jtkWH5cUGtadwJv2nxXzs2ciiPpYAhbFIe
IE2DZDqk0DZDFStw5hfQd5f4g8Ag3Y3UgJlKymf+tFzEq29fD2iExlU0g6Go
ACrqGa53n/vsLQNcKef8BF5qr1ctbfNCKu0kfeZ2joGUz+WH9bzalmYvyEW0
VkGO7d0vNb6ptdZ8VMHB1Q5dX7Vu8/7/fksWrijMTlI71vij9wdaN7UP+kXP
SK5/O0GPXvrjgiqYlJIK8TvQPbderBb3fYAlCmSueju5cYHXuJX3Iv1WFORQ
oiRmaYGVlE2BQUOYXp7/m/MgIswlCaXE69DySw6khK1E0LIhtbB6CLi1/J+u
BAPYnmwS++yCG+ROFkCbq7ACvH+AGm5IQ5wgscTe+nkWf6MLplmVkXSWsgl3
YunEj27SEKXnVnSZPAnD4nefn/MuIxuIoaQtQzbOakWtyd75gHV2vATRy4Ie
83w4WkNNXJ9BPe1BgZ2cV8QoRxPgqKXyISLKUcq+bq4KbyM8VoqBnHitNvhw
2GZk3/O97wVCnea9fYJKdzHz3TNBDFE7YNYIrZ2PIK+Mfown4GW9OskktnGW
oPmrkEIXPXnZK/Zy/4sAybAk2m7uLoSXIWnw/HKquq77p30rzBw/08Uxy7cP
iwrIuvc/XYhagCYN297Un3dCOkENUe2sC+NpTzkFX42N6J1N6Xu6ddQ5vDxJ
UNVVIHtHtcI3SfBCITi07fkiOI6O5OUiZgVUE3ZCAbZI3fL7VbNDdOXjGl6N
b5n1t4B7zomkd2L0s7qMg/VU+3YcTjpXLCC87Wntsw5nKOO7+hlpb6y41gdN
mtHnwHGMz5Q1+v5aPMEu6zNRYGUb8N8ro3LL/Jq0Sd4BUS1UYDL3X0UIuqEs
pnB255DLLqWdq4IAX7QHCJjqNyuF1AAut33arPUXvPYFrMQABy7kMMjHalV8
MLFIwH8aKVZYcD8eETQ3RgdFusENFXwy49xLusvQPCqd6PQiXUqayubcYQaf
ClUUHrfs4LYjASTLXh+sY3H+mVS6NTiKXY7UiZsh4GlPT0FpmzKA03rE1Lgw
G3el5wacdrz8Ap4jUX9GRQ4KdNT9iEN1wZDnR2O0UrGXBp44+rUGOEiQxK6r
knwJgeecGMfI2iLSdWC2ktaqYbm6/BBbhXBNmbTiGTIObF2KdW8srkF1C7iD
q+3Y0dvP59g4SBdrzxpmbtl1D8J1zThM7dBZxrnJpXZaKr93BM0vX487k0FE
OcfbpEtZsQ5ldlraH+xYAhHtGGorum5y9+pLNLu/6CWjGCtuy7GHNqRbzIRo
o35AuPaKRRLpUdqPWnGIeeRu2swJi+MFqJJKM/5ooGSQs6pIgRCdUf9UAukb
CggNDkVdImu7yVQ7cmxlWpPd0sw1lIxGG+zxXPtCtbwnNk6WrEWWN9gprEP4
3l/Z0/KD2qFEMmiAVkefNtJimAMDM33W8d7fuQ3wYgz5bSDq53pB9QjfhqSm
A+6QJ4edFY/+Tr1P2YTIFa5iYDdZ2/tzWf3m8Ph8FrOL+aIdUCy5WeUoWes3
wB+BNSJxYtG4M3OFsy5WwafGld5zUL0Jcc4AmCji2VtoJL68aOp+QoLsV+dz
Hbayf9/7HuoOXBbuma9kD2fTIVRx0xcqGHDrlqUY+zguAFR71p1dluBnaaYQ
lesK7tKpQRyBgDs1aiiIPp97iQWpHTjXVJGsRTd8jo5V+X7RZBNW1b1Aa9Xy
pdfhj5RYTuRgv0MiocOZMmMhPoXQcRZSAXPOWK+r8BoAscNv6uo02UUSZ+VI
rGmJDGE6RvaXGBIKFpQC3ks0G00d3DTf6mpNc8lFvdevN9YYnUPKmSlZ7f+Z
px2Wi0LC0xuz7TH7WMoJ5I4HoAOJEspyu/rYgE6oEwQW8K3hr/nGzP95FZ8/
qaPigXgjdG6PzCe/86y9TFwBZr/vkmhtDJd9/ybNiUYZvDrFbH2ctxlmKIV/
n5gUuR+CFMvthmeu//d3tec6rADafZRJGp5Gn/LFsZh6OzioSSe4glcFB1QA
P8cLAw0vOYT374e+qlCjRR/+GbLEGz1/v/yGpfV+Vz6FNlsSCqfKKarhQqp3
Hz7C71CFIQlPiOHTNT/782GLG8pZ07mJVUs0HhCq1Kigjmx9A3Ua9wmtOlEB
cIAH8QAGl7K1qqRz2bSZ+BO/QW5l9rjWOiooK7o3RKVy/nE8SiWD8ZKpbKrI
vmKSbQ+y1NxxXcA5CHa26dp0q+a5sDjAwrz+49gvjFZaUT/Kh2n8mhCr9Llc
NAqkeZv1iaDX52KXFJaD7SJoTtk/W2mDy+49Wx8ydqbeuDoHo7nk54tp3XQD
oZvHMaxdivn8lXKwR11PMVO2IzOBGpCckwT2NCzBItk3RanW43Qd+UuwvLt5
tlK9Ha1+mAI2jMI0WQEDQppuF91Fg3dyPU9Q5R2mu1vKCa2401tQbcKPHdD0
wIW1+Qck5CKCpCXhPe8j8aDkzT2mNmYGxKp86CfQCNKmNEMpazB8ntF9BC5y
o2/xBMyqxVV/vq/nha+XstcXIWfN7PdKmri1UjjAzvLLYDVdfyFrbtsi4L9I
KGZZVLVISKIwT3af5omrSqSI72wrrsdNwj6Nuft/MQ/I7Ptdjovs4AtJ6/6b
EtVPHXYM+vtWxVHWPHx6erXyiKCls4QFiw8SREFNQvZOnpXXeQ0guc1Bf/Qn
x8ogdYWG1hyKkHvHMNUuImKplHZhyrxisLxV4DHnJCbHm6Rd++WHRxYGt/lX
6nSYvWulPFgY3/WfoCHRt61G5YuMiCwRYWNi2oa+uXCUEpywdRhgi0hq3okp
7SsKF+kEiWyEMn/qAW9QXS/d/NZXWPYka0QzXri/wlQfKz9Drv7HknBXjB/4
7rPGB4zdS9pocffRbnQwltzoq5EmBw4/NwAyyoYVPXzEgSnrkp14XKgMzT2U
8azA8sFuTf8j+BBDz6BKN9Afwb1YjB4C7nFdoGqpkrb6LPMSbHnlb5GQFyoB
pYo44x0xIbd13biuI43hcy+3eFgmkk+U/hu8nOnDnavNH2kFuc8s6UXb7D6e
DMzh5wYYS3SGg2OGqOzcfLwObRreW8x2zXE+2WDZSwunepqg0rZVH0KeCAg5
r3c9fZQOoyeGyxf42KUSSblWa6IZZDLRTaBcEZT28bj8KEypLgEiKQWjOdLm
y3G7KGABnWOU2I62Y8/d+iORtnqMBj9ER80upCXkZvx65OgoCgqoEy+kLbRY
Tm/4ypcAaqfxkdfHw9Xsc3Tmt6WFhgjC2DgpFDMT/Qd2ldWnNaz/K9D2q0tS
O/Imx5Sku+AGkypl8tESfkNVLT+igvepfy1SQrQeY2v/cn4vRhr8Hc/hp7W9
4RS5rmGb28TKpOmnOYDVP6KCM/YeJNMzxtccmZFqSCqqUkmr2wpE4gmRSM8F
mMdDDprGKgGO3bSP+b+9EELtAgkVFdO017uW4t1kKeZX52FagZKhTV0t69dn
No3+gKgANeYQ/+G9oSt2vf8xcE1X6NDtssXFMTeT2oCXsnEs7OF97joAx6EK
qHmtz44xzpTiomxF/rfpeFo3vX8tjmDM03KtpT4DDHUGvquSwVaUZq4abxGZ
p3gh9j/2dpdUKjF+WHOE6FM6rc94SdyOR00DY4nBIGFHtjrc6AHuoZ+Hsiwd
g74lOQXDrEt5KgLzKMC8ezgiKCaDwNv+Sbv67fRvBCsdnrUukQNJbBhsKEYo
WWMbEtR0byBjZf5poDxnMVPnHrghahws7DzzE8+9pSknKAXP4yLfTha9K9+u
Qn6m3hYl6J/H/WnJAYhaz/RdqdbxBjoZG7im85sjVzMbzzFMihQYnTkWJRuJ
izO4Mbg/3k1mPL1T0+1BbiRSdQyRIODFEeEQzSiu30is9TN3VJ+R0UbqXQv1
jfIP5oC9f/4yvESA/1jfV/DBaviqS6hak0NDfr+xqbY41l5y7B0spE8B6DT8
KMvbqQX9C9OmejOA97D4CTX6TODjvrwsVPOB3SJnOiE6k0oEQRol/MUW/3g8
7fA4J2hIpCEvnTVlezZ6ZjltVZMIoqfZDKMlNhJJWZ4q2WgHWMpZeS/iH/HB
GJi+s8+ULOJ9d2q2OImEI6jXdI42WtWm97/cxFSo6VVgQ5G8WUew/qY2UxQT
ggJ8T/2fZm35CfQ7RI/IOyttms0LMzyOLyEyUm1eI0tAm9rP103I2vpaMJO4
86C8+/ucelMoUdGzhWPr0nH0zfUffS+F3appfdYpJ3n1qwLpqpgtLOp46QyA
+ss+B6BcHeG1HAQEK4qcz7ksr7oM5EL6w5o5QDp4360a+vwW794rpWII9jgd
yczj+oXd0b5LORCsE2O4oT6ANvHJOjWZ3IYmTVtJnhptiQG+b/Zyp6iHnGX/
9MjwyGZEi31VpsyESy+486EcsUf3Ch5xGa52RtdHUrVlhH49KaBLa1+YS/G6
MvE4B6gzTWWKVAd6eF1J2hTs02o27M0655UVIoESw6VqRNM9FJ2NFhZ4U2nT
ojorRrUd1qtpoPabUHd5msrPPnDN7GLTH5afrq9mhFWjW234j2Hn/aFQ0Nds
KIZv8d9SphCgxwBHAI+xeGHrk2q/dXl6cr2lK8Zrk3RngP5icl+qDoQ0xdrR
zXbAGspXNYnNm32hZ8R+/UaTB57G/LdL0gStJIamEJp5F0iJvc0uLqy4HuZ7
4mbU3N/1BxIsukyuWgpg7EQQ02hyL0QCc3drNK7qUQDVjfr5+tl3ver/fiGK
IOKe11fzKaP3Y2xqv56IACcsncTX/sUBc551xzDyra46kyFUQuttr2mLX8Iz
qvDd06O1cEZwIekNRnq2L6/C7aCN6kZuFSy4G8z9xXZ/DQAHAQm8xUPCn/xb
ny261oKfwwgm6Bh0obTZXPL9Mgtx3l762Ff6AjAUjZ3dTHriF1KWtVF98jyG
Pqxj0vjkbZvq0F8NNc2S2qSl9KZcmaXUAMi36H8eit+FlrZPBQu8s/eXTKkV
nL4yQHOZ1XH4gaO+Qu0ZUbmaP7RAuKuTsi6qhOCOBgPUdBO0R7uzJIthb3H3
i2kpvi+LW/apAxgQmmBl2rvqp9bDLSDl0vpV60/6og2AtMgd1VnKST4KOgEt
Agc0QjeuBzJY5MiJ+fRiAvGz7CPrvN5I1KPSfULwWqe8JliFw6nAnCM/kLPb
2lzs6hOUuqeJ0fjNP/s+bwvqpt8v7bfG06/k0c46t8d4WEP/KqAATn9c9oMW
yyCWr1ZzNMNOgnBB9df20+g7s9HbI1Fl7cy+SHFd2QEMGWPCEDO8MxxsF19Q
4mvwuXVk2gimGOOEpwshcfOmMq34HVW33sUyhiDdcpfkPbAz28JVWowYarf3
gbemu/f5AY0QvX/i6N8/9euseRMUTzY5Rm1fqE238H8lbKwbwclT6Lu3bAP0
XU5DUZHZtlvKtTAXOwapC4OdX2r3pYuyzMLwyOIDZrxpDEFpDGXdAkUmTY7R
DRdGiAyy9PCUw1wKThy+P9EfgqlR8jZPLV0Zj6yt9reDryG1Oc/TKCN0ilix
Wor70EqILz3ybPBudJETG4vNhpc16CHqZHCjhH81j0JDIaE+1VtL66ui6LT8
0XjsqNcxLFkd4pkudjNMMdD1LcSobxMhV/Dgdc5rqHA+pFQdraOXNabfHTnC
+GZgJGG86E7FyPpWV2JB948jukB4DOrpy+ioHNSU+BMUhlGDGs+9vkNTs2NL
Yr+lkgZLsOAopZS8EsrMxI3rYX0BaKhFdN41hxHQJpG+69eypMX8Bx+NAkHY
IPHQfiqKIMmmRVET+o+2xsQKnUoyr7Fp0NV4ANfvc5dx1Tu7ywivZZCPyUqq
/t2pk/IItg89Nfm9jRFSKzzKqE9FIe6pG4h1domF30PHLaRf0yJi6Hh1MnP2
jDhMIt1E0OEft1YJDORVhFX2u/2lzRyzo+vDKeJtuq+vJCaw6IuV6oO8ggT8
FMUxn7QjWPTyVIwuLc9wQ1U77jk5JwGhjsj9f+hBSzkWzKrKF/F0B3OuCKNu
hfFfLbbL5wwsi0/BPpvmN20/ZF7/edOftQ7c/sFbthWrksfz+1A5wiUaWU1k
OknyOSq2W/1hfvwdlwKdBpFGpWxV3+tFxt1lgZAXazWG+2NhtV5NE2X0kZTP
iGt+xLwM0IL//DCG2oPpyHMNe29VHweczBuMJW75YrIzsw0+o5rVtkbpuFQD
HI2RVDKcj1IvOWAGXpG/OgZFH2YcWbaUEgxE2sZUaeOxggwjI7Ubxy5eBPWw
dVX34ppDD6N64mskyg248AYlm5OcNyc4mI746Ds3k6+LLLwmmREk3h+tQtlX
tdHmjVFMaynHEqtOf0fNkEBCLqRYkDeUc7RG05Q2D5W0Sz9TAD4tt5WrGNC5
C6cGvYd9tvd/rT1CVb04xWizOn4Qd5R8HENMsHbcecIqWo+L+giGDP3pXUJd
bVHlpY0mNv3RY8UMfzz6JK9S2Ut0amdPyyogesbYMNzkyQXotrWa+tW91Sae
T93dVkUL2bPzeERZGvbku5qTYVVOz9m3rvlMcbdlOcdkjk+04mcxz5db7nis
gXp9ebJ4BItfdDgj4Nv1KA+CRL7yP7sdsHRC7Q0q5S/ul5IhXjDStrzWwyF7
QxJQ76EqzxLtAc9+6JsTE5+O1jskB7e61gh9MRdg4hSZ9hg0lQR9b9h/EDFT
o4FKuBh0hXu9oG7KYoEoS9G/YaPr4Hb1FaOTCeKvo313mNUpp1Otvv7nx0CH
TrHFtHqC6sShRR6c3kna/1aTQaIz1JcoKunMTYCiuliOyWZG9/gw9cHzffP2
pH0BLIi3bDMhF3fcg179naDpdHL7Iua4VV51WZmJotUZi4GYU5OWdMHA0ndY
/yvPulIGFNx0ZIpB+HnpcNs4thjy+I/+bv8ngAOscprhVtFT7ybGKc2/aVZY
dJZuBcqxbj1/3K1mstkKcqTYVNsob3S+4e6R53psq8WaGr0w12GTUZy3KosL
8j01sJmCHybxWp/M1YGHIS5Q5YBfHuMZcSolRjKT+ZR/zKjhyx7joNGWqIpT
bfsWdrFVYcVc5RODbnOQsxeM0aV4n+TqZKgI5A2epJpNO+YTBI7CDjP6fpNn
6R1K98Scu+gCTW+pojF6exEpZzUXvC3arJCFQ7WbvwuFqqIY3sFSlOeLiqHi
YmLwvtIryMypkBBlGVL91fLbtW96K5WNDbz1oGAqtzVb+8X12YK9o98VFDmI
Txz9Ea+zqPrZI5n+OY7a95oix8O19HwDgdZD7t8kaGf5rK3y7F1jsXVNOI0l
EtPfOZ4kOYStesXJH/drnY8kiIQEdPP4+if2yi2Dm5eJa8LNsMwXo96QliAZ
LV7hBJriGLdorspIm+V+5v3C8jNvVxiDvgrBhnpVmWvoKYcOz9JQcasTUFx7
10xthQjDPf9kXPAWoh25ETLN3dKLjCcCj0ryss1lUCirymxxY3LPpkt9DGPb
y0SW/jvs6e1S9PPQpg3JtM+iqDfxKw+3JQuCsSntZbPopuFRf/vYqU9XOz9u
vcr47yG3XzE8HpqC8okfdjBimswB4MuBW5W8RRUwCmIRhvWhGwZs2i8g+vNw
uk96aW7BtGSmxftUV3620Sirp430lXq95IF7NcEfRE+WvZIo4/zXrHr5osTW
HZ7vzuuRfVrRZFOdIpv/kWBIuea/OU1z2fcj7M0YNrqII9d+YXt/IpNuzhfJ
KKLHQNfd4rkLqkSx6kQ8T5VV5akIx0Agojn8fVB6/rWv/Y79h38mUESl40wX
8IyDiiMdMDJoPAL2AXD/cmeGuPSp/MKP1g7a7YIC/UVo4DD7ZTzDpJCgJ6Tg
R/Ny/voo0SYGgjVFGAjxBbxbVBobB91nEmbQajIbcLaZF1z6w0fytg+GoF/x
7SoC62gchQKKXnjJ6VAfST8bcRX6QjdX+m6AUgxAIyWoMcjNgkGJHzO3Z4Ap
EtiHxJQCZwzwpLIQ5nurOSQIKd0ZPtFI2MQQZ4ZX2iXFw8pG5ukX10QLH0eG
TtWUJKniWOyLk2tjUooFUST1k5f/4JQlqW8rbndbvxZfzBRjdbG2z4Y4IzSH
3lDiXyNCA0yO55SfCyEtUfoLPPt0DrqKPnl8UmdwJjMoa5u23IW13gof1Vxp
YSQp0xHpH5itp9tuWIIYFvzex5znivc2wHXtK/kZCyHd+x/IRvvGm6jYnPU2
gvQ2PLra0oD5EbSack3wBF0QxC2WoW+6tG6e6/EWp6L+EKbjKB1aO4BEStH3
oRTFd8E1Q17y6KBh7//HxCXxgohPZE2L39/zmRB4MdVbQQtDVRkYUO0sCmuh
WjfRoV//CMaIHPCx50i4GF6YoPT0t7DgMRRCSpNy3LrxaZa//ZTXBBaohqZX
HUT03A/Jrcl4vSZl5jcFmVq+m8sg4GQXsTYaRzDrp9+N6oHvXuUqkaUfXwzD
oB4RTnERJkHj25o4lttsoWTtii7wrPrSnMau/1oWPiYlvqXGMK7FTFqlXrDy
+uOObEK8nCl0fASstuq9Wmw/l0fhlGqgxIA+wpyXdTfOppCD7jvgLVhwv5tJ
9Ckc6BNnk5HyQS+pPx5NZjLaWN/ogEpXWxIlSfiHZYQM8nm7LWu/GkpCyIl+
ckjYWl4aNe7+ufIXKkzEsLZNe/oebRqesSEK7nGJs5CNmFVF7kmZBAC2fvrK
ZVyARogNpL8UmjGtNyf/DUR1q595h7xGak2vLGSkzAK4Y33X6Pz6XxMtV8Cz
278whpRK4DJvU60X70UVh/600ZjwQ/iJMMJ2g2VwW68vAvqOkb/wuqPu/wDZ
htswkPUunVMKidcCkHhkG2QSDYZAmAsf679paGTC2Fa75SoYk8BH1zG6tXA2
AXV7ayU6/FNqs7AXepvL1MbD5DtIElV1Evvw9Y4p8CsPtGSB7yxRVDFmzsS8
SiMkKwY8ko91nDiE4tNeKV68wuJyNaNclPyv8EYeID14OqHVHzrAzQ5AkIRx
23ZT0wmwfM6dINKhDtfn0tNN+fYij40KQfwLLWggIpAzzScfNX0ok9tA99M0
fXTXr3NwqCgIPYkqN1968NIyNDksJD+e11Zf6HD9Kn34g1egyZfjisZn/lQa
8d/ngcBpz7nPndJKxyzFiKMzazRXR9/lWF+rrPGP6S60I6p5QcznA2vJwnN9
tPp0C+6l97Wo488pVHB58PoB/19XQAC0P6PtQRBmvJ1Ve/uCEjg742Z+235x
o4gMLhXXRdL+iVdbSEFfKdG3026v5LrRviHcJVbcV3s1039qif+pnkeZXenB
/Ix9dGke3xKiZRHlwYkGzM+b4Zghi5hF+ISEbQS6cTOVNt139GojpPJIL+bX
KSmuUWYwX+MrlmJpTD+cPlr1kfHgrQaG8kaZXpdtIC/fJS5hKpmoeCceW+Hj
1kOM/2bx1bfxwsPZM8KhMS03qK7E1ck9gpYAaDR+MOfJUBgv/Q3fSUCbpmzw
dqgvJfJhGFOgqVwSQx0L944Ft3GJZ/8QWdQGGMDdfokleUaM1StISHb/6uQh
cv4ErVJvM1BtccGfrQghkXSgdVxgxyVTlmkzMVLUEjz06D4SQabtDdE81kVk
P24uVTV00js7UZ9Djjsk+p+OVVVkzFIsKxMQKDKOwKqmaFlLN+Ysjrp1TRKK
OpXAGdAvAAagEZ8m3PiNro7SLKTiJykp9bK0bllTt6rsWNJ8JZ02IUH0oFfS
OIL04iNG0qPZoKQwxZeObzG4j3VvWDVxMrwtetvdIyjalHjf44+cPdFR8oQ1
IdRJeNqgZqmMBj13FUZiYdUwy03sJcuDArYqoK2ag1YuzROQaeaNFhGuqviq
jF2MrUviuD0SMnxxd+h+cW0Vr/StE1wxwkPOVSKOpbij58CmvSvtQ4A9/JxT
67I3E1DMdqBP39T0RfTHbxU126EgMsNY1oenc+YauxGlvM/09SdcskXCbU0y
paHkKDLN2chEkgjA98TqKp+zVxdse40d3hsmhT/XuFVp11X5hMfX9TRY4OnS
APcqErHHdzUyqIQ6c/lS2SfomwTFAyDY4vVhFNcYveXLvt7vfFakkWoqcsWS
2PiGgtzu7HrltmQsFBUndb014m4EiieCcAbB4ei343EHmK+1ZXfsFUkT3NY7
3KA+0YNYmPp7h2/r9jlVrGEjS2LBVBIQqilzmZejFnQ8Km2Cid0mCtTIXl59
eCjFku4tz0cHdqlEgtYcUx6bSaqZJ/ohmFtgPMpDhKYfgnDnkoOscZxdBPFW
pRtVFMSyruAiCJE5fNyb4bU/Alt/LOtTXBM1HEeEkqLvPNBtdy7NKVNGhOGQ
0uGjpVJbQlhXOEspl+92ZzcdlUeHkNea805UtjrLXnvHJSIBR0RQJxjgI0EG
d+o8aRHOHv+uIul0P/mzIWutIQFBy+veVfE9CrdthsKI0zbU6Ce6wxhzNANP
Hu+gh58i8e+TczUhIFJSIhhSB+UL893HhD9F8RzL30YYBzOYyBRGwh8wXzPo
7D8/XddLtACuGjKLZ6wu8vIVRr464gyqchOtzojvM85XundDAYbRZORTlfJp
N2TIOYHNkrbiDsErYjtElJiULQao9/03wj9G7h6CERoO/hvQnCsSloshKRzL
GyBXScQx5cBykTcm8Gz/GiLNfsEc/EfCb6DZVjY43aMTFWOT/TbqIgcdKxHC
zUSUbGDNpeN/mpabjwv/VNFbQvPlaNe8f1lmUQqc+yGMM/43XHGhJWBOJ097
xf0ILmqklBuhtwrFTA4DkHslvGHB/mHV9s/b4OFo4RwHjzRd0m53iZjPAhTI
lB9U0j2/ji5syyg+GsPVlT8uZ7qBZfK6PMnJX4yHtmTiIJc3uiK3j73nLqFa
ODNf44cmZz5xYRDj6K/F+epsQ0zpWxlutyZD3v1q0VyNzP6UaaLaqsM9jwx2
eTaIuvOorPEppSQuaxza8S1fYefYiQI4++5lwWEI9iyCW/+/EmAYj4EYUWXt
QB982CiKbrea6s742bgu6TNWqZfML/qlSTvFtD5sXGFgeQd5oOK2Pq3eO1GC
pH0Jk/nFgOP+iGtuyE6yUYisjsJUQIjdYGR2p4r5hp/Xq5HgrJb4KYOgYhqJ
zCpJku7HW/HI27z/dkp+9suysQv3T/cvza36/N+M2bB8dJBX/53ffcCZDk8s
n/OXSzxtasdLY2mkkKNrx1qEcyymOzeUWpwy8DIlDIxtoszf+WJ3sRBWdD/7
PzRQk1TukoDoKxb6UXAUdPc8ZU63baadfzglN+EVt3NtMvI7CI46IOLXaXdO
Qx6Pyny6DzZTaA2xK1wqhgp8t1LTg65JLjUVjMWpdc5cY9BQ+vKkB1g62P41
7Wqfx/8l5RqQxiIeX7i9vfv+wSrGWt6LRYsBosDhm978mMWcax6bVYbdpduF
KA2KQ0hYQ34dfN4BDP/SDRfAz6T3/pQS5wp5oidATvm/IlwctykVrRkBfcQ9
eXpk5RDEE7gb8fxoQ6yUMYrm5H9ymFZ4o1V+fCfrRJCz6N+HDqH+DrQ7iwyc
qkQPyaMfK4huZzy0jvJwZRzYNTzmui/i1gZqhkNrLAfCBeRNnrir9O+dmyb8
aOmFvYoF+jrVk0PJV276S843k5klpl+EQfwgnn1oKM2ldygrmAe79qsb7baH
2p49NcS/y9G3myuE4K0CkRB/pBBhbVPqicXlbZz526BLDb8Q/NhjLp1ei7zJ
vQ2dGw8lZadLrRX6rQNCtWsp3RbWb4UdMn8Td/GxHmPq++ww83YlWS0wGebl
YHyaEsjKoxhyZCB+iHthW+hqpnY22CYD4XOOuRHAAtl+KklukPu59wNUu4UQ
A9HjH132q/NV9LeK4KAS5ah6drD7oVl5yM4cmVQFNbtxqYphTAAAQhIcr8zy
C/IoFpxwJ6mJihMGZWs3EAyUvlrjxQW7KM53QtKr2gntf5z7mbiyBiwR3/1X
OWovg3nxAVd4BtVsfXkDPoWMVgv2eAbmimgoQsn4NymOMzhXoWX1eBnZAnw9
sZ1jqGVNwkavjtMmR0JlAE4ELUUJ7tPLsVHVbLjRSvRjuSTwCQjNKGsdJM3k
g6SNQKPM00TyDXG9ScEYHIEb0MrymumcDoQ21++6IwsLOO56A87juL6qW/5D
6uRzCPYvjjJiLH7zPLAfwzQv58QYIzjR5B/qD5Ua1XfsdMpFr8rnZESTqH1+
YfteHMPkiAu871xMJOsYmLrwVu9LcFAh0Klo6L80/sxqHNnSpGmtjOSwC/xx
9sXYtwBW5xrgHy+KI/OMtTDfFp48M/DpUVvVGb94MIkphuvJPPi76Qm74CVU
mfOlLXY/KF4hodg1CwXl7ydRz5y49y66X6iPA1v18iQHc0GP4lE6ZdyIR8Z3
FuTjYdcwg7IRmQn0tj0fUX/qI5zV9UK718VVOhVnWoY8NS70JG0x8eyomSgg
W3d6Afx9bfe53/4junWmXU3od8sNDB9VjCgg5xeq0iZJXf3+ll3kLSTgNQ4o
BSQcb69uxVl1Jyl/tzUKgEcdNW1llQaOXOWmSj5N34PvOPIUccxz9GaQI7cX
Vdju4OWuVVrFbmE2Pwo/IzO4YbP3l+l6dYgBplygQOXCStmTmYsFKQgOv5iz
Hqnidp4D4hBgEexs7thP9T6ebUfeaKVTEmEZZxWctcfIELoYA7tpAt8eiiFp
eb6OGiOQVN76jleL6nyNV76N/Yk8D3Q2+YhmUeM3YLnTpFMtxSzWGRRiW6aI
jV8UNnfBf+P6bfg5YtDeEtcUWtEBdrkNjNYU0ZCdD4OmerACyChAiLs82Q8X
bX4Fj4QFU3k/7JuGSBwhvv4QvOphj7L6X/xX/GqM6rO8f4kJDeXscpvvGBsY
QR0vMtAEd0toP9SrIOa9eztySsUOa4qmIV7PO3cNH54XVpDdOx3zd9FYd3Vt
FQCIS3Oh8JjRn87lo8wLw+Y9i25/jcFQRjdfSe5wc8uA4DMkmeFT5/5EKQAG
Zh/vw1dHXz2J2YgFudHU+HLnnfjkv3x6tPvgaskh14OXJ7VDlJLNDmoACn8+
DaRL2eXzuy2TBdR2T2W2IHLs2jBpR1mV9BfTwsbnRV0hdRddwLLkZdsALfof
tEbxXcPnYMP6QrHg50Ox+rydrk/JZIOYVYBWNcd0DFOdh5gfvtMjImztrprl
9HAUYji4C+3bXLU83+12jjV6ZHn+jmOVEICVm34RDBcEeNVPyZgDZld94FbT
92g6oMtt8Fl1gVH1f+HK+hvF3kky5EURUOpaaLiqBGgRYY/+FdwCkVr0g11G
PxpJNnUkHlgxo4GbXo05M5tkgyVBPRI0jLuiH5+WCaRSIKHxBFN2WsxoUXBD
NQby0YxAGkrwNRE+DNuyT6x+hSZpePn8PPZxw4iNLLayibK2iOTamRoiQgUh
k5TeiH3lt22cJENftB3ECtko2edJ1zl56LjGe0+dWRONH5R3yrtDxJfZ2J3q
kpK/KnxeWQauTecLyx6UvBfMELYeVaD2roc5ZOG+0Rp9FCvS7RNdXQxRwIbr
5F3KTNuD9A7UOiJBNjvZlsUHP76bLnIlOxsRfWNWB1TDVEBDtXGnibDPKRoE
+w/iAuYJVVpyWg+ZBt31ZNCkF5IufjFaGJ1XQhppOQCNiyOI0ADIoRWflPDR
Op4IYTEwray1rcEY+ntYRcYeNlhHHUHUFIzNaQB2Hb+sVgYk1+i43XDk8PpP
U4V3fgjGH0o0S3wC/pX7ote1NVMRQZWeiUc3C6IOArcsB+6ss3Lb3ESEQJ2i
MGqXWzyiZgbjXIzVsBCIx0z+L/8+F1Ub9BcmoWeHq6PiZzdX5htcotJ/Q9ov
XxVOZSrMLKp6+8U/QDMWBok/icnycZLmq0n6CIfHarIO3WyoYBn0XBqOxKVO
qjyvgHxtMW6FSiHs0dKkuIT4Ok98JGQ9pLFuSZ8UKNVatbK+4a+yYdh+QWo1
XHB3Nu8rV0oTkHwyXb1EEqEA77quTB1emsIurjBuJFeinvIAQNgtxwwNCo6F
sXLk2z0zlS6onKxOK4iZeP2oiEgie36CbQLvL+sRgIlc3OjKLHlaYFYhFs/G
H8nsoV627QQVTzTOv9XCy1iUyAoqodG/XqmIcgAAkTWgbQDkTV60OWG3pzna
ytdnJBAKx4irDnv3+OSv9LBORDdAZM4mIMJFQsgNyRyAIURgetC+fjPHDpO6
dXk90ob+VEiPEjzzfkPryPfiqEBvkkrBkS8nI158bdKKsedIWJE556UAJyci
9cdZOyPBa03kuZkRsnBraH/zO7lQ70D38wBeUn5FT+g++4W6KBkE6ANUMKDu
RyESK/RccVniVzsfhvAEpjcXSkPSyYHz1AnEMzIJhZlWWO7M0K9emI5iEoXN
FtBQfo7ShyO+Z31VPdxgf66AeBeS5MPntSsjq0HGHtWz3HBCzn99uybrSJji
FM5+7mQF2oE92kWvGhXjKGgIUHzUsg4uTtxvUbJs9LxfiygjWOMh6VJXp+et
5cu1Q0iiC20LkYjh3CAgJe6STI2PoUg2tfIXPHzQjFbcx6rg03wYG1xClMnh
ZeDVVCkfGEip7TlYwkPbTPNP7HIOK5mGRdTeON32pPF3/S44aVrZqxB5kTTp
i665nZuYFrwMOxhKJXpLPNBdmzgFkrv2BzfKL1T/6wkws6QXQ7Y53eHxpKMQ
TMIT3iYb0NPGak7tc1VsLAk5B8k1iS8aMM58J/DAeYRCgIjdp/NpyZkMDoGA
ev/3BRjEzh5sGlnGZKHbItQ32vPMnckEiXFc9HFK8LVzQA3Thn1gApsdc9go
FNzyT1JOiXbuEj//mqIRPJGqOPAZRhDsNrH8NGSs1LcKTKczFRN/TdGx4OCB
OvLqqEXlG33TG2y33M+5p4JzJ42GYqgtOaUmR0S73E0fSTDVyeIn0MnGuEBk
6hsIhvQNtvidWa8OLxCsHeI2A/JJ4hOhaR0+i66C0xoGQ+QOvl6zlST81kbe
Mxr0DQ/j3oeW/NmxvjR1BbA7Bx4fC/4V3wYBS18aFSelXNOvA8WOs0sVaQJe
vPTGAHpq/HxympUBgGcVkCiao6DptSNLDmG+f8iqQZfA5RVVSojwbAHHxY8Y
hMW+XqXJFc1Fx/TbKWW7jPY9sSV8KcCOUa+z4DkPkUg8HPiQAz0YbaiWk+OJ
BH7aB5fJSvx7NcCsz606dotyZfCfbR7TCLcIiUG91fyYU9MJ/6R+ueSLJswD
jVbleJTBBLGARsor8/Uf4Q4LCw2PYPYq86L/o53n0M5iVJyfil+DPViPJZYr
zS80I7LDXKsUgU1LWJ5s2UsraPWvM1WjX3WrbfC54bK54J3UdPYHcOhxNJ0q
1fRrWKuwY+MjsSEO/4xtsHhhe3pPdw5LofiADUaqHi62i4HDBkkDWdZiQoMV
pzSfIgyjaNKq9wAT4mvs9WU7GRqeVoAnhvj3oGTSg5aBiQOdFpHQ9l72hejd
V4oHyXjbQ8YAHEbrBvOodTXJ5GGJ3sf59K5oAIP8UbafNKuevAbaBok6H7Sa
SwvZh2GBjA1hNnbIqeolhR6A+JVw7x63s4ciH8EX4QGB1jlb3teJkqkPkUav
otpkqMd8urtHW4TAOQgmfEeOVlknfltoEKqifYHE76mnQvuuv+xuU3+PmkU4
7sP05BwWSrcutoL4R4DwdvTDfq/2sn3ib1PDYipAN7+SZd0Sk2sK9NF3dPIa
hYjNMeiaykIHsz7h7fv9te2m5dFEjdPacjs7i6BsRr8w8AOdxlotIgeVbzCA
CHFa3kB13qI+o5x1qXMEtLskPo7TYjsUgkz/ZvAlpvbzn6W7HX2qFJwfMYzj
RRunIb4j6RO4IjtW6DOjDYdguhiTK116Juvr/Q/Q8jWngZOeiV2Hua00nL48
Cf0Pca16mDLoRj/w6DfDApzegxLuuAkPDJFRVx7lZPzhkJ0mnLDIpEp3hrIb
mNMZ39yd+TjsCaSl7nY6DsJvlpHGx8EJLRz5CnuqfsD+wufr4lWs4Bm6znUw
jJyXk9SNFNsWZWw4CJK6N6VUoR6gulE2G0/TxK4LtFgUKV6b7CMKAjnLUVbx
X+ZQfoiD0gG0n3btzPssSHzDyA5EbZqUyEL4N6VZ1lpL5kKNhbBSKlNEfgMW
+ngKaGZFu8Ds9MoP7/WvSmz3qaQ7QilR7ALdgPzsMdXRw6L2mebSlJP9lZ9R
C5lIBiGBq2a7iVvTE901m8QVkvjjToEnuLZWi0eBlkX6iwN21MTIPzrJOfbm
QjITtr25Ostu/5dthk4XkrF9XfoZoprCWyK6OXGaVzcM5TmybkOzac4Xvjkn
cccYqvNkCkMnVlrRnytmCZ3HXzqWjRuuNM7CUUozyD8WnDJqwNS42YH4FsAk
QxGydG29AdTQaTj70rCXNBS0JV+zSD37zahw9UhN46VLCrAKhR88lNz2yv7/
4RHA6LmY2sHCiLIvNVT0ldsymUKS+4zkz3iFRCU6Xp3mokIoHetjzrSm73zi
p2fqnhnNE4LKX8yxS39wGsFU2ksusf1M/NMr6QRKqnW8z3mCUgXeOKp4Zoxp
yA/YzYrnBpSa/dVMjAkYbIgy0t51WmxvR/4nLecxMj5clbOc8jbgUyaZRqUZ
EWcXK+6o3+xnrYdDkBGluBwW1Ll8BYl8TldbRZzo9PkD6Yz7c+QhF/bMF9Fg
n3Fll+CTFZbr+fyvh+VhA1HLP8fEoN38Dgk8qwFj9zw6QFzaMbr3fkNeJDc6
Gxf4KbT9XOHTEIFJkZsdO7ywNgKOSw88jCItcMqS8/tidlCvWHB6H18wE1/d
OdnM80VA/Y3YEJ5h85sDdPeNmDJKC6xtqgc//f4ltm+MslM+bmQBGkuCtqyv
f7Yj7S2GUW9q/yR9/fn4RRtMLzYkTJ/TeuPTfujNxDTQoF4+AGLzcroXCfFu
TFwNFFOaRRETHoIBLdc8+FrKxYZ2uXfYwZxnxyfxb4ejUN2CkBYQw97gsBkF
CX5dP1yVCEvxDIF9S9T7H/gcj6C8GnSUIg6ACj0nP9WS15FDDbcYjHVCprgR
ywVvPJBTV/vGL5ESEEB3VYl94muidCdY2nbKtd+lJX4Ki6tAkUsrdsKb0TeH
vF67XPofuWpQytfSNH0Sr9avPpCKtfuE3297U9v3ecKD5T4Iy6Fqgm0zwCDA
Nbt5DxBTfxHV/1br1vxK1zpongB+6r02Dv8irqWziAJEvdGzOXpWp9sgiOG8
TEAu7/lcl1tjZvjAbCJfi1ZvykftlMh1BrZK8gojeAi3LbEkExtFem549BAp
8RtEA1Tdqj3ljMAn5aRXaaoqU5i3A9c7xu4ii7Lb+Tf/63KhRSTR8P76EaXR
gZhzj0l3aHMPZltSQPqIIIsAUW14+7t0FoGMeXaWDGESksTUBnvQo7iAxSfC
RbW4B6cFivnAxrCLI8GfZR+1Wktf6tbFeM2+KRX7q8ECBItezkBxdzGG6ih0
pnXzKzGPoNb6y36rZ+BMOVl00lhuwPrGihqvoW7eXWM2beJSWMXTR0d4M+T4
bNzyV24IffFsyJbSRmXA3vRvgBIAu0Oc+mzRi0+9TcwW4eSZ8ONu3fkmsp7I
1m5cIrpLCUQR5g6MNCvk0KgKx/xTuLiScYv6xIGsevarIw/g1tbJ3zriX8SI
P2cTm1925gyhXpfH1bFiXMEZyhuYvZdAKIBdlnwkgXn5cFv7MsFxwue5IHJD
pyzKZNU4Y5XlqspZ563uVUTZO1ms79/v6Gt10Ejqa6Gcx9qy6BJcpkLMC2Df
/10nL8mz9N7HY76i7xKkp/wiWW1NjmlcZMzc85FcCtK5Gp2NV7fbwZLPeDaU
8sHTQ71IaxWUptAcoSR4B0/4z8JEV+R61W+8hiJTr0IMyEKGNWA6NKYagrfV
oQAFkvH4RFs8g8GwaF5a5oFtPI0w+aHfDI7HtYjs/jeKcqsxFshrtv4fk/pH
UsvhFJZAMuugWg+umwUisW16Eb3z7eMap0zvtS38JYGnSnULMn84FjT0ZfQb
FAmr89JHPi0hhem8XImY3FnM/xgyXPavnxLvPzY2+fzgSK2MG0pI7BVVh8R7
q0p3B5HL/5xvHWvAk8McS/noRauf8/IC+CofbADIdACJlNCvJcD+6IfEiOvo
yidRLPomfgXleG9rURnKENYw8RGv4v09Rz5mZj+5hSA6NVvIzPcTjfDxUeQL
Ve+EENbT0Wg4pDGdgJl3sSb9cbWdhTs5o1Z2WxG9IcUFUsPaBL6zqJYf8kz7
1BtEFDESazzLxbwDbLq6q89/DPVBtUSWvyqzsJa0bWM0a0G5c2nrO8u18A/A
1jexHd+0oJ3JgoUi9nrGi3ysGW+l+UZ6GCfvXsge0HkRadChyfUpAUsUyaGV
sGjx41h7ZRpsKE/twXQ+ry6lDxfXzpw8xs7aq2BlakUiNLL+1H82Up3aN1DT
lDGMUqPgZyPo0Oz7zEN51LjLsnNzhFsViPTEWajHzz2RU33I8hTvYcUv6UrC
hAJoC1MB14s7xzKmGqcL9oy2yEtVe3u5WJGYCVrzBtyoW+sCQBRw0U+MyiCh
mbA4PZgSO5c7zH/sZYRb9XbE8kksg5TxJh7Ug6YbjgC2hVwuCfxtnB1F2KkO
Tx3L8EwWs3yqTVpt9l6Rw8qSQY6e455ivLOXczNFZQB43V34bo6viLXbHL96
AiqCwKbduMldAWLwmBV9eYWPtaFt0uuK6eZWLyI7haJQuhKuYe50Vgge3xMT
bY9bkPwrtZe1HqYl4Ye66nKEzUxCzrl1Xt7PdomxxAXz/HCJtSJEIuetkRlz
2Rbw0BwXzaXrX4GF8UPtkrD6YLfYsJ8fh08CLBBpnFuQfyhJCnFzqQjI1UWg
IZz4osHb+hcBJIFIDYBGCUULjgyrJZE/AipJvjXJw0ynq/ahv/bUmOjH+uWU
qTiCp06Vpmv5NoAtgrL+ju8NKUDh6/8KfTFzwHj0kczPngBTaImGt142O1Nb
Zn41dU0hYnlMWLFkBaCqRZ0BjZX0kYW2A34M6/KL6v0zpMRgdhwdASAQYA79
0Oz5wKIsw8trC0KiYDJIJg7zgzl/9evEXlkJ02ofF0DtM0k61p7KrJejBFiN
scT4bsSBwyC1UXk8p6slFw/TWbCYGnODQ8IMxLbOyD8kk77e9Un6KLkZLS/1
pbFe1Tz8oQo4/+YEOVOPyTvn0iCrJoWc6rbEiC9Hv7AW9cxHhqzr1ucxULNz
UyjqlVC84gFKtXUXac+fD3HgWGpWyufmef8JePDwjVinpAsFBEvWx7lPIpTx
ck+jBtUMRoXPtSNrykJP2nJz5/9oaW7uIQLTCRYy3zoby6XTN895Shfpehe1
IgYxJxHOAT5V+tdUr5yLZa+U0ekc1QE/BPP12z7wyibIdXMFrJ0B8zik7Pn5
TlnGanX09FOwem6bKNni3ilu/3pxVHlUTdfCszUaVpoq/rHtDKkgVeAW0GVg
V5QSYxKUCrkBXJMFfk4iH28IwralwJXriQu9trhbRw+bnTBT0Z/nUqsd28vQ
YoVdm86LKR4WWdR/p9TuD8qtNIhn/Faa7HHZ3D5Y/+a7SViCldB99D+yDk9H
5f8T7MEIXyhYA3bbKJFphbpuU3+R4w2lXb15eVjmQNHsmBw65BD5KqzQxlQ+
A7LA5T/coqOJyG8xNklrAqJPfpf35ZMhKOKtIEpgN51Hx+uc5W0uZo4byEPc
bgrFet2TGN9fa9O5u1biZ1h+6UyypedUAuqKIyHo5lD8X+7LCIOPu5B8NiFR
ff3vhVs0MCvPhfMMuuAq2Y4BaNdtUJ/L/5WwwyoVkRZIm6Cz4JJFOEsmohdT
z0zP1sK+mrCcpchjJyGpjionLxGso+Y909VjUXuEPgrzJUNdXXmg3Za0OR83
n1MojltZHHzDmOcDMFEUaV3hfEl776Z8dDl9GkXDxS9jEsLlv+wo0Yw3FfC5
OsJwj+1SmRB7UhEktZZlJQejKy60U82o72SmQsyh18KY6rhzkv89PaIGezdZ
94y2FB64WViijccdM6+DbYGgEGEDWda+TIQrT9aeeB8d3+W4LURHnmC5b9/F
F9LAskDJWopaI0JjJnHckrPLwtQsxozcHZ8WNF/nZjRQ2VoVaSEv4Z3enxqk
V+mIghZsxV1dmUlLbPIXZL6uHKk5D8Ss4I5HdEeplZGThw0YmEgIaKeVj2ph
8u58sC6GJ2WY/hD7/xyM7AxAnEtCZ3jvAmdH2wp8jVuM4B9yfGz+jsPRJwkg
H0j6g4nWLriQeX7v7Y+9IPx9dl4lnh4swbdOcR2DsLT9UeWBg4QvREYErf2B
P1fLiXTU7j/IFmWlhkBlYDbjOJjOxghibEsDKtM7kKdv/NZ8GcZ+UDhLbTnf
DATL8vW2xC7FHTK3BgQkGBlEpMUlSVGBWSGpHDMlV4cRoMKrWE44i2RTf2qV
FpFrEijBm94MWQJ8CazkemyUumD+ODGNYy+1JUa73ScfhC8omu5xwcs+xM8r
c2EFvgh7ckCHAciv4MTE79lM4kXcMMjt0A7klxDRDruIVTGDxfXK7VmdvRgU
0zszrJU5Fp+UEjL1JIwkZLS00eI9lleK3yb9/0JJzC992DHDpGA4bK6JjbwS
eLGcRSWYkei9zo6MgHhWihWF55N9pyfEVwjeRxoPgVxbLU/Ey6eUu/jWN81M
+uigazAXJjgrC9p9WM9QNulK2kjP9s5AW6zcEePkwi5yK/C8R7qA29tQOCEV
52aWUwtLE6ODqpToxdrSXMtRrZMh3TlQFf7jHPtfz3PCrFyhdDgJn+IWYI21
5xpiiEIzs0D9+Q+mz/tGgSwP6iUvWTU9J4XyQoQqgcZyZrZza279xA9T0nlw
zjicoAG+ocPEduAJdSiYILIiSn2LQnYnNtaZt5Do4OYLwRjfIokY52ELEFw0
+LvdJwDAZogdBloVz1cJL3ejjbNRzo3c3KUnw+E7USmAOc7mwtjcL0x09Gpg
H6bKy+rXwlzr64hu1Txh7q5F2aWzTN8e4W4uekMOubBvTIeNj+KDGa+lpGbP
LwtYbsPdUJqje+rJpVcGz5eBR+GmYcUOO5k0YVdotGGYE7HtnlnMyBTzJCRN
K0plC+sN0X65WI3mf6tw8XjTpocXFh5y093Y0gr/BggkDcPHuWiDUr1U+MIq
51zbKYcUBrD7VF7YgikCPWWfnrIBGPiELH9R8K5yYFXT1e/7CXVtZUgpZDjW
M7V79DIidcrqMHJCTAYL/NXxKLgpitidR7GMhvfR0AgCpcwjcPU2faLRwvQI
n1pV9okehdIxYHalCa3Ti/nuKO6ukKl9XJwcOBrQqMtd9jXekPmw7mGtkmSp
2NVAhEK3YRSPm2wcv4OtgFL5kdNhbYs5yeQFLcpHQLgiWcGhjxo6zN3AbvKU
wcTVimSZawEhqVyA1+z1oPyIn7m963/83hfiBR6u+madYhnr/OPEWfnSgFxH
uOpnHnVcVwoCR4Ll46PW9dgdIzGbPZDKAbd+/uhgPvf7L/CBBHDQe55ycpcI
TDc16keANFUDeeOoImcCvVCDdmGJMkY0EP3oz7NG3U2lxzNh+Hd7+2Yig3FS
X1sMDkkONIJsSVAMqtV2l2B4Bx4gxTVJBo38skbNne2ccQ43HQTPkQaZ+cxI
cCvFCKwF2knIiM6C9KZGTouraGTCffsB4FkuajZGWl7+LXuKqQNoTcDyWw9s
IYuAVNMsneca2cbxqPcrlpoecVjWWMXLK2UO2v+UvgXHUQRKUAVO7shFR8id
KB96Dfs6rUbmteRUp11TuPo78JQhPvGV6heVbEC824BrlXJWtAqnVpDGEM2U
n9k3NvmN18GgXMlWYWmq5k+dOIzCBCT5iej5XdOU6YpUmf+T0KJpW6DfrFU3
xirgrv/pH0lnMOq647C37tMWPVw8a+9Wq5lHpZkOF7ZisbJSisYQmcO0pANL
mvKxvf3T0zhbLzTzVoEilSwpLtflu0EDLE5UST+2bC5+K7EQXIaXXjR3y9lA
v606Bzta87tjsAu0Xq4Qq3PAXkBtr4yIYEF4NH2+d50nwvmvfT+QhbS7bd0N
NuSZmi55OF5UANXhtt7QyGkmFZggXGHUx2hhCLthH/yLsDYhMNmIqNub15x1
b/eYyD6xPAZA6rjku33LQF0hGGY+48Ut+Z3fKOgXgmEjDid6e4U/93vMJVIO
qvKvOAPyw6u+KAMVh9q1AZlX0+ZmwCQ+Rn2m2T5LNBnwgOTJUf9SGD7s0SvG
pQLCI1z9Rg+GlaLL1QNoEyGtXC4lbu4mzkrSEkMD40xPer9QiKH6jKggLhMx
9K34ozwSxqsp8L5QY2B4wZtKe+P0cctGxglM71d5z3ChLSCHtGDk4Kc/Et2u
l5+nZhm8o1Oc8Mb+LVARqrW3Q98TqKLTBTQBHZ6Pa+BrpvAFw0P5g16gsCb7
mBBvyhaoLk7v4c+Oh0F8Q5FTjh3foL8ElJZi9SmS9S0/au4x4NtMod1ky2k4
nJ9cG/G6ftMtcVnQUs0ka18FjRX0FdlO0W4cYyxkdESX0NZKvW0l+fgze4Zu
u1E67dtT4YFDhJUqB+HEuwuGau0IMj0R3PW0wPY8PPuUqM3qMBPKEb4YAKxc
Pz53P7g0Qoz6zXPcCI7SzsOl0fyFZ47CbF70HXzBZEfA5k6wSTBBUMF9JCmV
hYW2jUcNXMAYT/A8TFpxi7WIjnptCyOqEq4Y3d+wuk25TrwBCMsHSzudFr2t
bMe+gbumTKfkbbHHyN+flIGb8xvSpdyfX7lUcqN16ZX+wSwW1iwg3lXMcNVr
stYu994qYzwNXuzmdNjy41QMe0p8B7cbVvc+tvEtj2pAZq67mdHZiUt7i7WV
/5OSrZGeGd2kdylbfjGUir1aAcwQw38mUHb+QrHzCdlvLG4unEUy+iWK1dfT
v2wmtzZIAoJ41b6nz8cD6lgwv19EkK2S1rRxzrCxQS3awAwwpA5ym8DeAh9E
cKeByqPsRHIqf3ZoAi6RStLnBfvPp0MYYwkCUxLfG6vjvnQPxPb2cRokH5uK
wUXiyFADv23JoR9dGoBXuhASU/OMoIkIjtVuCkDcQS9p6O9AvCQahzDhodd9
TBG5RC0NXziugfi2eL3QC7an+sjXU8pzE9i0f79GSJYkHNJShXKM8Cki/B3p
2yJtrI06jw3ebbl53xF948OD8FUvl/Vbt51OAxGenvtK/2/yp8i0smb3pyF8
remEPCVIo2pFt9P4mpJ/Vg+szTFIH2vF/R/yye5iRTsR9xbcVnsp+ZrcC3hO
ioScoyILSAOYJXVie6dzgTgiK897UvP+1yAnfbFRg4xnj7rqlGlEMzFhY2VT
fe4rmXViEhbYM6e9f/dVpVa0kS614KyeRUyBQ/J0pMHlVg2Fe4ZrLAFcvtjY
Fic5B41ukdPW6DoVITbAFCX+9fQ/0Vq9iKV/bOXMzJyXeypvpSE0kblHV0sg
cd/kgZ/8hvDZ17QjepRxIIE9UOPhrG0uillhORt+pOiVSclbIuT97tk3p6dy
St3o5hHk/OrjDjkRq3r4iUAOisIftrftHs+QeIZNzr/OhE8ZnXP+VbckrgD+
JofWmyw3C00b4tpt8Uy4NgeG+6AGT/9gTCAmmjGpdLGGcc8+05T3r3MZGfEo
kgb8Fxo/XUbJH4TwyjoJhsPpq/yR3jqVdUz61yCw3xVvPnUH4pKrGfrWM8l3
T2tZoekDrZUQZwQVaA+0Ad0x4RjvFT3BCXXKCsToMDB4Q2ljBX5hTPXqmJG2
wYJpNMAuo37HPw4GORXoWNZ3VAm4gmYvpxdvwvEadGcPpYOQiK7iOWXG0dUJ
qB4AZPMIKRgcPThxHnllsz82ozonoJj7wDLzuAo4dMwNFNROiEXtHci8xyBH
U8gTYPmVNqc4JjQpKoZplavViia5Fofr0/K89BIsAyZCE8a4656Y0eKYeJ2C
aENl9bWMU/6W/kuThsmcjmyRByhusaMt7z4a8m++OZJBPClYTNtAseZwQwO2
6vtJ1Ih5ptz7uz41BJqWsaxfd9UCElffkpmt2a84XgGNE7zQjUZrfiZJK4KV
4JyeqkyspZJAXhsK8JHbuoDBigNXz49VxZafKzf1fFPTPuGouMPLeh/A+zqv
S5AUaNwiz93uvxq22j0i4xivjjEuKXYeHRGTZ+63mDebBq9mLAsb1QLVwCEV
y4luWancW6H+QbOewXQd5DnRUVsnJ45gufyBsZJaBZ/WfbnEDF+221Nxopn+
McecbdTpfTTE2XjYzMGqvsr6e9+2CsAGHKrLaSRnMQVfbmg98GfMeRtb5uLT
sSC1QV5+y86IJkH8etq9TiHRjWD/wz3OlFJ4NL1/mk9si6MDiKSf4kx/nt09
Mo4g/IiEpi2nM4OGxssEkOZpkScLVMX1kFSfxHkIl1UV2wzXjf0sAVKx4yc1
ZjhFkfak4+xl8L92C+++Cfh69bgaKSlP8R9ImQhvLeJ/vckZD/T7xvfs/SFc
ZYc6Mpele65oHH9vofkVc4mlA9KLsEcfGzgnTtKbEDDFqpUCVuJDdckdirH0
7HGYSnDZbQqgWfnQIVL9oxQUPWiizsiEbqtOzSYEdfg8nfbFceh4YtHVjA0p
fBmXtgAA734qh8dOm4oJtLMTfL6gUcJLTEVTZ/KjygX3nAWE+O9ENj/+mXXI
EziCZQHcfLTloaum/6lJoNhmP2gmiW/DLInwSKTOP8gmShM5TjJPmR01OCin
ZwepDOjYtcrvUaq1Vnu5zwGTAuZtZhlOTCc7FQ3Ufir6kv8OCQRjIBnNOI55
LgMtYeqDTDOgoyr5bxTNY3FwyAAIP0M/wR8tX0mM3XxImAkRjwxFdwZ5XtPX
KFiHYZiuQYmRhgHPQEzRFW91/R92Lu8ue1jjbgxvaxbCRrHFp+deZSHzf1m6
iAyB8togRSnMnRMRvRt5iCPlvrsYPepk17ssJ7y25JEoCbxOn58amj3ymMQI
X5FJAWo7hf1+4/JaFBNpH1uizVtLrYoZe2EMrfkx9hBRWF/Y6i0DqwrzLE/4
HurzMu/IWT5/WDVLjTFRqD0iP0S51KBKCZRY6ZTcKF7qoU8Jo1JarL5Li4uF
XlM3Kyw7DZsG+lWDnZdKG+mb5TsVsHRCc5pCVPUMOJNgyDbK8YXl0OxwMAXy
mmCemqiY6bZDDm1JMblQIYiOPjYewBgCNPu03YXXyqyLmOO6GFH/I6zgcRv9
cHqfoQHDtMMdvDP7PRNbPm/xukkoMoHdEOS6yg7QJAZnCHv1elCG1yHd/KQC
E/FwSzk+H0NL7RfKKPXjXqMc8QvIdI3v03QyO2m+9cc0hAFPDpoFb1fuIOCK
KGxPz3ujVy4Zgv8cgetQfo1MOlWahs0vq0pC1VbxCZC82HeXbqrdFZDm8DHx
8JAYqFudOie1jT3uEyZrrSyj+P5yBj7M1Xm5TrqOeWgBKn2Mqa2ic5WV1ORt
jFj8o4f4NHQJcOpboPmd0HTA9QoAGtQs1CZAFCBFreDa/YygGbk3CETPLWA8
5uYx9xTER78EvrE7SAzct1QO2mud5xTnMNdmR8gtCYIFc5iI8QSBn0PLEKab
oHeIhb2U4JCZFvDyeGH8pwQyawUfzs8ygVNZJbw223UPc4TJZxwpIGUZRjdm
ar0V05de1iS3zbKS/yo2iJJXxEt5Yk4UtDtuVG9SO3oxSj+tCAiI/SelyCsB
KTGatlwiXZdiWDCyVFLVT6ty72TlbAePXrMVeFzaW/IAJq8x+ZKb9deXFXFV
4cia2Vohz/cmUBwDa/5QEz7YYxewG5G2wpXY9MXsKa8XF/Wmc0/xKXzaeMNi
B9T63vXZBWG7CZz4ye2KZs64Z6sPYtKAJr55J4fwdQurUzH4+dwegP2s6may
Ua7fdIac1g+Ex4FoPj+uIdvgXdp6W10FsX0TCDTsXpRQyE+BfSBp8kqcN6Zc
LRNAiVZr8a6cqK81eOGBAB4/x4//d0NVExA0YMtAxKn6EocWuK8EBjawiC4K
An+RU/NmsoWdi/ex1dVj70+WPdBA/dWSTUZV1kXZWT9/c8nW/uduWScQAoiS
uTJzajE2BkT+A+8fEgVuQ4NN+juE9EQivJC383JJE6uwPHvEJjVKkDvI16mk
CqwXbndb2SCVAPwWrpi01r2Zs3gqAXUy+7E3yumJVDhs9JjD3LVprF2dY9C5
kcytccFH4mfV6oKIqyjwVaNNCbVoOe/SX+ZVHFobsdMNiV2ZEJpJXAj1agMy
76+yWaGcAngO2lMgWP710LCnCaox6i+C7t4a0+kLHMzBocdq6GfVJxgnS8dt
0j8hhYCOMh6hE81qFg1dnJUKzc63SH2f34pbOJJjnTM/GDbgE/yp2msbjGyC
9glo5HxpJ2UnvKKRSj4Jg5htYHnL0xg26jD/uuveUE4HVJ7SQaxSEMNUWJOd
Z6aYCmXCvUj89PkKmrwjoBB8/5C5E47XedmqxAzPkKZSha3rg5Yn2reYtwYm
ZOaiP3JoJNG6sS1j1GMeRNjP39s5f4NyRiBX8C4uU4tOSgLDtSyxMpPO2Ozf
7umGvXP57yWLQZzJ/do/1bQDO+y00Hp5Lj0d6R2A18Q7kLAUS0I8F/M7lDma
OjGNR2KBCuX/KTVUm47bLP4wvhvcNKSTktmrAumebFfUgxBq7L20Y+Q6/DGo
9Zau+LaE7/mZTYisshP8u943mpr9CEU6lVgo4aEP1iICp4GffFDumQenRAND
J71jnoa/M8MG6O17hQ1AKkYkr1Rhh0+TMgirm24KVU0iO605trqplGRemKIg
CA96exXfu0bhLyehCQkg/cn+9hXTXUTfmySIJ6lWSJ1PjRo42bdpX7/83TGu
oQNL7jbqkrTw6KPfFF7DxcSncMAMWpcnWuj3D7JjY6otZkUIlo/1FwMB4xPN
edm8x0YROZdt0iddwtsdAMjJORCeYNO2zG+yFtdXMTq92jH8goTh8T/Z8O3X
c2WvCXm8I9FVtDFb6chld7U0co1ffaqahmOcWK3tkLb/REU119QL0bCmUj1S
8wm9zz1ih85jUIyBf3WFQx6/xpt+ODOzX6KcZUiqw+fCdu+qoZ7aHEaopt+p
+Yav1O+kXI85tpWdGuuSYpiuKanyDS/9sAGOaRKEcczClW/8gJaaiTX5kbBm
wWj3TqjWExDsRedz09cj3w+ZBZiClbTx4eAtMBZXpcsfXmqDAnEAqKS9y8TJ
6RpHtBDDkhpXg/0BwL07F7j61OBLSU7/Ub2rzoEJuT8HkvMzpT84y+HhaSjo
PjbO75h0ioFRTngxK37jePNWtRlfn6YXWy31LLuZSssMnPTEe5w/wqfHrDnn
2do6yaHmGrlqKETVPJ8b7YRJ6iWeoKfxYZ8013FWvYrIPOQNoLsejPQ07TWq
ss8OqQJQT1Qvw0pS83GngetgE1DnuqAb5HqO6ZcZt5U5zw+nSrH3REpwlGQk
5kaedpnNZBf0MPMuML4CnqjGErLkkOWdxlb4muc9o93jEOTRRMmY1QBhO81x
C66Q/yRtMfZzxZbu4hcipilamIuUhMdp+89RZVbUrn4yD9bZRpetL98tlD82
tMNE+El+LRkOpg1NgaXc8MOseZNwBYKrGZ3PTc/dfDrgFIcvOQeAuRpS9fNa
L0RHRQAp9vbXu2FwlpjBxZ/1Eu346JGukHQqzjk1/RYcnKYxWjAZ7YiqXSo8
LPJ1w1F+Sq9/vhXEXrgceYP/HJLxVcYz3EB8mUy2aR/W772YsUjYpaj4eKe+
FPOtrvhGJUKS8n6mxRa80mKZNFOXrN97YXgePvbkiasHcKfkQ1hCxbfJ41Ee
fgaB8p1NRGVQ2Qymglgb7hAdOqC1ku2Jpf/QLfwiNseBtjQ/HaRLtD9mqSKk
tiHJlQhyvCk/JcYBb+pUaaPl+ImKu1tJkhuZf6L+pPBnm//vRgBy+tN0hDEs
69nd13MY9vR6BgKOKaDCnw19E3QjjGzXPg37ifEEQ6Q081LxUqrEd5RpZgcU
SdeM6eoYhxodsuGd+QV6+7nsVk+1d/FPdVVhM7rYPvMREEwwXtJ/pfMK+ao+
xje6O/HfFWU7HD7LHI54wc2i6uYhFiELLqraztFWujD2wpIg/lbQhsylMLIx
Kwgob77ODOPirQASzkytzAbEV3o4bYMZmCP7rBY50xecVPPBf8Ivnt1Yhf4m
BIumryyWadB/r9ghCrgsp/kARZoT91isvJOIL8ySyyCIdpEH5sX5NQr/3uBU
fOlW2ZeFbsQ/QMVHTVKOIvYiERqkrcl74kzUywmVmHzlRyVcj9BEqpsyXTL4
Ki34JyMO2CdfRxK1y349lGiHk2mr/UCy2V3RZ1+ctalWH328F3Ynzd3/LlMy
9u7stiX6ph4Y6MOnFbGKJQQqYs/BLQPLxVfFSz0F0xPQ3wxian6HedL4nBoD
kiYBFhMXVpgz4RgDOTnL3bO1ZS18OHo2Wmi3l14Vg1VdLJlBLTAdrE4FEtDW
YI0nOGa+hydwgWFoqFhieCJAt18nM852CZtchrzB1CSKIrrPCMSiPkQkgpCj
swdI4TZ6Sup4Ev/9YtGB89d5cgegWzd9A8zhODsYBJF9uOgeuRkptnhJ9fZ0
vFfHbaKFSC9SZid1XgaZAioAk+UPUdWsXWmzhJBEqKgFi31oDsib9BYPUoR8
KHnsRpXjfZ6SxxP7sebg9ufsyotQcfX4lENjD5yIfJWyJomh9ZJBnAw34PdB
2Oi9wWN8uFRSPKKlk2eEUDiRMIZW1IG80ESMWPj1xx1rtwGM1a4ezt8ntTi0
HLKzPdC3tzUD6P60aacOw+JT8F3eBXo2Y5R3aj4Fj6OUlCT8XjDP24DzD0zU
qogNA0qM9frcQC4pWNHcPiAywgzPY05Qnh1iGaqiH/Qig5+CKMZ+Y51WvbBH
F96CJ3fCl8SK+Mpf6Atu46scNufLfIYfohXEN28hCDBVjpF6dqAp7DLGEUlM
zx1NDCAFZwq0DQkQELv8Pm+HnzaTn8xfQMeQCqc5CmXWdxkNugEvZf3ywuIg
6BCfTA4olfWC80Z3PnaAS2KJECwHq+deZWYwCzV/ad3M1pBFqMa4VrkZQrQ0
8TNyy4YR9lVujI4bljXFvD7OBm3LHD5DgvIGxW2gqVVOrO7o1o2fcl9CJhG8
6uZBS2k/QBcNpLwpfbRjb78ePgLGtT3aYLdFJ4naJRTSeQEA++uODSbC5wdj
jd3UFdpoTLJHUXlYyT9nld4VMlJ1YDewzp0YrP+xRLajcn+go2qS1I2Hkcit
Rqsj6GFssicaukAlSC1nva4JE2LM2PA9m3DoVMyR1dHATxGeL3OGh5DjjJNg
YcgQsbRv7GniyyEVu9KeX3QbOIvH3OIBjn4Zbuf7Vp9AeSbSM5IAOLc3FmqE
7mJeO90ThOo1yKv0D5WwSTUaC5fMpwMHqlLfSji4/FOb97VLqGXSb3RyFApw
jL2DH0WEkee/PE6LoU1l4VN75Bnwvi96UkL9c2SZX39im6T0TzHtf5xRGW4C
cyIcOYfjYrAYose5J+L9TBFYULj9b3sXBtFa8FzopGJFauq7KDvBymLIvhy/
q4dT1D7AMSixb+843v/+Ulcnq6XqgJGA3rEtj/hApsh/PeN9FxAOqVP+5Ti1
5j7PG7buaEDUG4l+13/JRk8CWM+qZ3b9w0T8Cvo+Xo/fL/tPO+P4MigCXUBD
jyvInffeshoKcetYkBdHj592UP/QXcnIfaITRRX3VxbDGcutJ0jy/hmNfPNz
C+mtaeGIEP+MiS+aQPx/h6GAwj0U9gOALOqwoH1mRCGn4SsWQi1WDgdBdefY
aXaEnYqfzQsAmzM3fiCjvX4uy3+Nq6gxjhhxF0AMNTAb7dxwEL2/9ltD7xLl
OClTtXpvdrueKweTgALj9700Z4wXeJtMDnTgvSUvw7Y8eFO4Edq5eKA5A98S
ouhhaTvSSm/xC868eE9ibtJAoM6nQ+iP/7pycW9mjZsVZzjRWShd/TrJ+TuR
ivDpiK5cwtigkyxnHdkhJrpJN9vtmCsgLdUBiOI0E91+Ez2d/OIXi779kQWJ
EXgHZrYiDBhK91r45pq4If7+zpq/nhOPJjNNP1A1mAwwkvOquIGY4UmBTlwO
MsHpTlXoz5PIVEd6mBPrHd15CwFmzkwJHU63EtTioZGWqHU9GT/jrkDPfNGn
UvgYiZ8u44EyKZ8UvKPUnCRiK6cbPoNC3HYyzgo6bnVjMljfft9bqhpIvaHA
3ctJEDpHeim9kLJR+qJt/75ikT1DSzz8BWpKVLnZbL73DzUVbMR3UKejnr5Y
uyVUsdlwOwgzZBjcA2QCMbS+pi4Uc/E/RVSYm6/iFb6jp65ZJNxmwuI9jgUB
tVpsArCryT5jbpaPA3OCQIfTJ5us7nwg/guL5VbEl1lENF50si0yj32aJlm3
b/OQXDVebEz9oyjpY42DQHi/Keg9mPx05qLa3SxRDiTovreSipasgSUlM74f
C4oHJanE3xpgusoG/2qFecYRQGbbZqIoCOfPnXakJqELKY2oHDnsswffQOd6
Mwd3NmtNy6oTH/ogiTQDSKGrYepuq0k+bqL7tw6RwqkXco4yDjIPtKQpHtgV
TEXTAbljQbgIV8iRfPnwVQET1tm+2KalBIJqLcxHITOi8AEHITqcyDpmRnRX
VKiruPPU/LQop2aKX5h0GuY3a4KMV0rkTJXSLLo8yYNFbrnxZihPt2b/fxE4
kY58EES+GBoC2utu4ulaAAPZRoCICjRlQkLKIqd/bXh5LdA4VspRTeNmaYlj
/428oz28W8hFBHYBSab1gqFNIDO0SDg2SAnmXLB5IJPrCpJKTARYHVu7Y+yZ
GmB8gIVnn7ctj+Zr6nQIwi7q11HF8AJ+GoET81cKz0GTtK0i9s+JHNJzHIGu
iZIcZVlBQEdxJ4KsoMfu18n0cJbnhiPXRwbOg6YEda8z/xIy9UDoNasH6om+
Z9bqku4/yILYXbNElSzsLHG0LrS/mJDJrY/4XpWBSqBwz6V4g72NlESM/I6X
RL/oNC3y3Vr4l16cW2Jmiu+Vvn7iqpARAaVASVCiOm+ymPa4jMmuqRhV4a3C
VWNCR8PFmoP//Yqbo/niUJdJKGJRG3/mCZvlbF+Jv8OwZvCam3zoRCKAh61Q
xDTusQ1aBJxHDthhKFHe8bk7L8FrRRyw+QWh8xSrwbEIIE8W3gxnc2sl9xnk
kluuJJxsB/k8SQVmWsxoJjCSuQ5hwZ/U90X/FXaJJ070IHxoydTmIOVyR2YS
Hpkktd7pZp4evqhDSoU3b51H5Prp4nCnFfIbK0aGhJ8KEUUE0rOsR8ZZFEuK
nq+Zp0uNAQqTTgawgL+fGVEM8+zYSrfcOMAAThZjtO/hHBj34iv8t4tHxLJj
YMpWyP3wPCTvgjSdTpdBqDON138h/jxvbUe9M/mzDoS4QZ5Hml3ejXrFtPWv
/zMtAPweXPgLxkRF1mBUmAD3oZpu+mKixO5Qc2oX6dd9s0JXFOTBlGDD5EA+
+SM/YXeNxxknNixD3xrR/8PZJeKENoimUqvojNvH51lQlcC1i+Ck0jnDjnJq
oz0vzT7NAHvQc8BS88UShleSmxPLw6azdJdbkl8z8b7j71G72Fk5cnC78Fmb
dkmag6udICJBdn7/1OzEgpJIAtYL9xukW9xuTS2hon/sweEk0TZBJLnRgjAx
4Zp4pMD3aBUcQf0/8gCG1k6pntROeFNJ4sW97Euh0zw8WB6oJq4uEgz0BdxI
6wsOeYdmAwYja4qMbMHjHo01shVNQzvZF3yaskIBf366BW45ai8pXCh6axoI
vygsXtlWc7Za9LJrP7EGAcpUHXsml1mj4AAmrW7n17mKIlAViVZ53Z8YvZJQ
oeV+zLFF1obl87JIGRO2azO8b86U6S+turTCKIuV5Y+DUfbuJq+tAp17BBrH
eDTBlyHFjgBxc3oXZtuO7cM1UrxqrtuSvOLf/t/o2Km2aPhk3SLaj2ll+ZF2
vzBN4sHyEnXJuFctsQk29xYn4QFbLXru7A851DofcrRAbe59v1VjSv1r5xmj
pb//Z3tTnWEmyqQamTZoYnmMhOTTYj4mP2Ut0sd6AE8k6jb6Ln/3P34D5tR7
4+bKyZY1ncUpjzNOyKN+rXbkjHK24mkxOJWms4qKOFY3dI6k/qFZhO1E/50d
NEHb7AahTjeRq4r9zkNdv2r8bxKbI+z+HwbUDLOnFMqsWDKOGCOYhCgmsBTM
S6qCBSRapIg+V68h2EowfUu4ZWhXNPEANSH02vVbMxCtJcyjsussW11NjrrT
SllkCakebJb4ExmwbzHXtuR7TnUGd3UoPM/L1rPTqMWRNosgApdCeS8nvXfN
8zXakY7ZWxD5JQn0btFfV9pqwRyyGJ4d7DbVJohri3nWobIpE+UOiq4D8BGJ
/nBsSrSTmkYKu1cSj7aKe/qekbngzFwQyxte83jRLZ9kCFCA5IcJV2siY6kR
1ygbfDgg5yMQKs7BN/S9U5kFe7Y8mL7JzPYeiw3mekgW6MfmzWj4Z3sooV+T
Cu0CIxOTS8nDHGo8t5YPmvwzTOZcxrqlNUYtNRQu2VFOv3+48zsO7zNlneGB
Lirluy6EgTUQN/vP72wTBdLpwnuyFJWWMi9XdX01L7sToganD8R3ysv0XOvj
Z17aRysT0qTWFi7PzUZC8vrWIMX62jv6dV57qi5Cz4W7kLd+I3LJXT460AeT
+NrIjWc/J/irAioPIpZEy3gyFwVHepHCOxhKw/21+hyU5+l49Vcz9fM3Sm7w
YZT32Yk7UxRMVxIF5q6cZCK9hNOyylImj4ePWLRjRH12YrOOM10wYxQVebxs
FeoPUQ+AJwcVZatSzpBR6CAsZD3Q3y44LGWXxB8xQjkP+uJxdB/oBc4dICvK
lg8TANMa55MEDsTICx7y4UDkgPNK36oNZ7u+C2ZejBr1R/EpfPyPnZ/rbkbW
O6jn5/yY7pceYx28oIVv0d/6PM+7w5OY5qxaVz/tZDY/rIjDsp4xXG21AkWd
r3M5zYMPVvHn8yshS5pfsJyBWf5OXQHVXaJD96ti4VKp5OJgDPgzbXCDa/kM
k1ZWeeV9Ca/w49EigbtOycdPuPI3LWcxE3sMH6FzhLUCr6M9NQfyct6Y9gzj
PmTcFQucYAlVw6ibzhedR4/Z+uVtXKd1X6gwOGhUMJYYVQaKoIEGlZgeK6Pd
vXuPfpNCKE+xVLhgVBrHhJrKLYRIKIcc1FF5fLTMz54zSXw+ADVpp4C4gFX2
B9M2IL4sLXDtXuVxHWgAajUQhb8FTfypR/YkNqOJ8rkYIovPwK6ID5FO0DcC
zNI7SfENtbkeBrN5xHA0YzmtKLwaFtw2AwfgI1UNgcHK4sJHKADiHtfIBv5C
wzCpByG3d6HGcuuWhcNON9Vj8TE40vhkoEHN01cci/pRxJIJ8+GyS/y7RqYw
wodr8XtRvQZJWtvCumxFyp62+vgWyuudR/ZgSuzCEYwY/BLG21VVwIkU69p2
RYp3k1tcRerXwEhjSEMfH1ZvyLhICR+z2XrfH5Ph/x16sSDtNvBOSi9lMDDX
YVCV5REKz8Or9aNcOnLF6do+SElSOIEYgS2dBu8Ctcu1NCl8otif+7QlXMmw
dxho4phORBafTMIeSlPZgWjRsLfu9UqmO5QNbNQM/jhrgE3bg8RXwNVeJJmZ
FNoW55SAdbTEDFcdhoR71SCUv8AGAPYQ1LkNaJsC1pXpu0c5X63x79fHfTWx
HYw2xE3HgNPBKNH976c4BYwTkU8KTFfYW1jKB7FXpRuF4XSLYYoi2EZm8Wlu
1kbzpu8Odzjp9QF+e2FwWUl5gNS5m/HZgJDU8cJCkZqGgGbzEyekEg4PLYoJ
jk3yvMWd4jRZonBiNtqS/yKDWPANZNV3yA0e80DebP8SPLn0T9VWPVNfZ4pC
+ppyKJtRHFIzlLD5gSVEfptmwb30UO27F6CzvPGeOIHCagHKRi7WasJpRG2Y
RbJ8oW59nuts0BbeG94/zdXssSka2n8whpuRXVXPaMPQn0K3JGXnPmCw0gDI
YxctxlHjdb9tiDHYVZLV1w6cN+vmxwpGIlqttRSKRvL1X72trcU8eNyU7vUn
p4Oz+0R5hg4/XWue7au1zPWn58J8rpzqHdMUVCv+8ieZ2JfB6hex7T/JTzvA
92e54WsDoUmGq7uJHh0JK7z0YOMpYVCFwEnK1oVj6fKjOxeBgA5nd0bBaXIK
QEI2z5H6zGwSn2xdULIZGi834bqiMHxkbzl4KeGUBzMXqoa89CmryItm1hdV
etZIqDKsSiLHNThuLjwFwoTdtO7AjRhzXiJ8CnlQvA9GJ33WpnIBlsYxyqiZ
ymsmxivwta0btDomLov9pWa7sFjJYno/CN1FRbfn4qTokjbw9MPrnf/rTbo0
HSr176S3obsZuv7brk6+2Cu8H6ugPUmZEMKhJdJ5fhpZlX7DZj0I6AKkD+uR
Chpx2fO4gah4kI7MlZInDnMYc13NT1M5OomPFisCGRbk6Cup1Es3Q9ZbzqAk
etR5EDOuzuUAQOlq0qicovgBd/k5b+Qw6ZZ2jAL+RbVjtgg11m9uO3O2VkLe
s5R8PFC78R8xUYwqo0lwZpYjtuQs4WMgF4g9vWkRMAXu0c80Qdl5U9C/IQkk
6VttKY/syOtx9Uvc+sIjODWYRhWn453MkDJp6+SDpaKZovHcW7ElIS0x8/Rr
Yx+/N716QJ77ywtLJV5GGyHGyrPcDSNBgjMPwVtyNGZqF6NMi7KLgh0+yHdD
x0szr70ApAj+JYdG2gMx/YDvOM6y3Z680Njm3fUJAQxBWHxtcHho875YgBqy
SPAKGDGaBzmXqtRnrkvc89VmRQb5S1z3N8m/+M4AztbyAtrJoskzSwZYzayC
dfVKgxrdQPpKCpTsKPo4OKZICakWEGoEy+puXyGOGN+R6lIR0xUZ7bBFE0FP
fCLK3lxodAjIA4K73bBDuwKNXRQgt0mdibLn8ZatMbAa0Urg55+k2+I6Ocem
ACnVuwANs9OVacT2y8Hrlv8hDhuoCjFc80Ng+Euesns9tWsoz8IundC+lMnp
VG2GOyPVE2kFPaqjBMUW1aE5RuAhBv6wsq9DoeLsTAEsdHnet3E7f8H6JLVZ
D6ZzoIzGb4rIXBRVSlgZScG1Z1uLkiX4k5npbEYEXa0jmCW1LzqXeYXVPrNo
9r0zwN9zIguuH83+qtoZhvcrGBKVkSHp86Ak3Xbx/m2u/gjxbUOKvlFn+scd
a4CWwKqwuNaXbD3u1a+Qw8eTirujXBnnYEEX5lutVGVJBw5GxkCxYWbxcsEi
UewGIppURuDU0db0CXSr1y2FPianjOy/6b+EfNXw4CVHN3SFOVT13nhjrRFO
5UBPpAzIhYogfqGA52HO0GN0PQbeM7OLlIq4XzxbpUS15tZ08A5DbwVoJBac
LbC0aTHkzKyAUTMzE3g1E/3apPoZzJl+QvZU2UPt2XP4GmfEJbWbdwDi635V
zxfkBzSm1F3R00vC33QsENrGS6rAeD/CN8VFkvkzsXEYOuM6OnJxrtAnBO2P
04iPVxvWBgtRHkUpUL9o/BOiWaDwXe04f26jrQGwg/OYXkw6JjAzH59IN35m
2KCERa/IOChP2VBagL94qrZGpyJQJcXEzAnpMMatFPdmpZTmQX+zt49iSfqk
+piL/8XRP4Jk5iMZpJMHuAz7kBnKLo+AbxAfQYSt3BS2xm3ee85SDNQR0AIA
z+aZZ7o8pnkBvqP5rxor9EhQ8RrsuFJj6MCEIMbM6vvaqe0Ge0rAcnbNZWLg
8gJBfhJU9wuq34JlMOpl8eu7c4q1qnCBLa86Eswtkvrm3oU+KEIUjd0xa8jJ
LrZG4r5MgfQ3cmqFX1F+GFRq7w0kCibSCnzY8trhFDBQRz+vi6tnzzR/+SGE
NPdH+lGVF/dT8gVlzgKnI0XA4jT0gWKOAiRsrjxuHgKqlFL/XhbGUJ1MwrfR
j9sfE3GlDIwj7BVO82yREnsS7fywitLGIruoqu0jq4PZAfU1JmkraC4mb9VJ
m596wqIM1OHcdh/AX/y8WdBjxuJM7XiBmckB8DbhsxRsRtoYL0VXuhNnZhf0
pyzqDfi0GwylNRLnL9yYZcq3gq2DQ3/d1aO+jVW1xJUkfw6/NXN7BgW82E5X
P/x7rJnEwedUNmxrRXCafzOpTS8xkaLFoilrYvuMt/mFuEsLpevIPL0NJzt1
2ZPjQ/UnHyHXxQhDyeitTLT3IBjn07m6NoGm+bBqSok1X/rJCmsM5dsAJPCS
7ML2m+W7+dBhaVdAHko3iuIBXbCZtliPgenPnjGckznNRgMb6bCA00cz/olV
gJZXI7k81b6m7PwbfM/8moaimwwFvy50RU6FcAb9bhXzTU/dTSlmyoyM/BMI
EjaYdeoGX/lkGDEzGwgcrvL4bpExzyZVRiR/s35Di6f+xt2AOx+8Do2Jus+G
DDWpVmJzPwiaTBp8GzSKrtVcwMWFCfBk4PsVgTAAxVNX9UlgYXCVPVLe6dKp
VWSVka9Cks1ow9Y5QMy6zOkpuJlMih9oMkGNU69gQujqN2KpaQcWaUhBqS77
+w5Uoo4vCyYdfSeZQg9hwbYpN4pVnegxbIBs7vszJR2D2mh9SPD3zfJLDKG3
Yh2RKnpYNYbEoR67FJnWjdmN5an9kO2sa2AcmqnJhTPI3hMhgREBqdxjT0+2
h/xNrhTBHLYZboozvz98DrdzsBPaohA7zsI+aOaZLwLvlHqfXOQbdVADYrYo
6kNFt6f2u+Vy3l6ccytJlZlOXVasSakGkupP+KZ2TauYhK0rEuGcalz3IqRk
YBzeJyU/gPq/R7Ri92b1+Aot8A0nLJphkzWZsQKgHu0KGEuW0wQLx6fCeVGn
FJGTVAbdHUZ4xBOMUtjWHMXnUBs0DQTuMMM6gynzDgWQWD+/cGw+R5YkJISY
tw1x48qwnW9y4jxUon3GKvc7DVRSrEdfdxAe89BXTUzpvGn1wBBmY6kh33tr
6m8ttUmxpNNWQGgilQRFm74mhGD3wpmAeQPhHueTGL4q10GSnqbp/8bsGmMI
/thH2f750jjg8hqbU5qH0dRYjJjud9ydBS1H7VpInXiDin4V3lqzv79dHjfP
kjjoop1FMYGppIHGOwZyuADE6wfwmOuU1uMYSgyWknuiuzXu3nR2oh7uDw1u
aZ69Ay9JCiJMTmSiVJQAyLEiUmOcoveIKuG6dwWeirvwkp4UkMzqD055GEgS
GCwR6NKzTmeLj+ENFYrpon+9kiF9Pfkq/6w5FGiaGgJua4IaQabpp4Lx2Iee
O6xL6ME76tKLeGR/hjbk0TC4pv2nrkUt+hR9kRoMMFbXoRKUIMAPcVmTyNVq
SCVg2gznKn3oUiglF1v97L9KknapQUG7zUyK67m1mwrE0blGjuZ3mq/lK8Yg
k4GCu0Si7DqXGjeLHqArs/1pyKotNVSgX6HFWNtL8smPfBATT0z/g8AtHVz8
J6ZhXgDTnDChREdJJCrr56nkzemREEPtTchoVWbBdPQTUu2PKTPYWSX1CHp4
3bxPGc2UkLQFo1UFyi+DHr5dT5AMDaKe/BAwdB1MI2d7rOeAirK2nI5G6QAG
UfTa3JDXswfOhwsHXnX494VzmXYUGygzXeRMRvGmsvHBO2QCBlbzMZllMRxr
JOMJYk11G1Eqls+/M/8nFjczqJHrcBPD/w1G/D+k0WOPe1YUVxwwyfdbJreE
gr2rSxJhmw8NyXzYVz/vkm+kG1m3r/pEKBdDzhQ6dOjy0SBaedgkdpYEyLOc
JDQKYuoIIKOFlLHvQHtx2nhKG2W6h8nlFd5n2hl1AymP1skPTuJ/Hi76kFBE
LD3DPskd7o3uCsSrK8+XnsJCxu0p93mSspRp80LZtE+Q2FyElHDC5eOObFAF
VhzGkaV9r2d/M6odaD7grXf2S5Nqu9tDALWZ470Nb2ui/h5tnEpek/ZyJ8pf
tvJCoezE4RtJmkekutvgpnnIlLXd7lVg1iFV13nz7yoiHfA/6mHJIanoMCtj
HA6imxaHtTAWhPHcoUKA+IVkGW3ZpSbwBAPa+cNwwzTM99mUocMTxpGb4Pb7
EzqxSAofNR7rVjul6r6F4gxcxXQRpETAUKuQAlX3sHMYHuua7uDSI+7V27SJ
97Xl7aExRR+NrxWo2U6bSF96Ez/TIHAp2sqpVRyGfrPZDtruMbxL4ZHVuPj8
NSztKPOaKsSNM0kTEFiTMDmH6bb8CKp28yxV6dI+XwQJNGFIcPjGZ1TsOwtO
fvEmsrgsN2gvlFUUaHOlqt/nfnT1N5KxxjtZFMPefcBMmpjRnHAxVBAILun2
myiObATbx+MeSiWHiIZPe+cC59UByZpCYczAXtLxoFjKGxen50JrDc51cIyI
xIM5ch/1ts5E4OQj12O6tnpKnx+tCc0MfPu786zX9ulsfVrWUfwMJSio+j4I
j+TqAe7/NtGZ6+R6dZ+QBJyZpwxAIe10FZRArJhHtRv58oTpAvsgZ37xKmuf
YCQJrL5HsTWF0bTeoQMbJdwewfxpihgX6qjU7DjFC3UcDWmqPch7etf2VsLE
vD70TOUpkVukjiNMvuQGZ0X08E5Z1volKD35iw68MYnRBzozobPqw2NO3yOP
/zha364JLQylU4rj/gjwo3F0rf+KV+e2dy0/iraCXbp7/5f9BRQOvpwAcFhg
2tzOsQLoDJAHn7veNrl8JFW3aNG3nSij3SCwKhH5aghYDPl5QqiOMg1W8vaQ
rIWnEkWsYpfRRwbVUfGXJShxg1ur6Ypy658EjdsVpJMZDTiQg24og1j+x/9z
40WvT0hZ7KL3zgmZSDa6qaBRZiaOJ2NV3Nh0eD+V5WpjYa61tqF+lPVebg79
PfmAawMtm5nZxLnIzTT1PsJlu6vSGb/DtHK3eGfR7OcHDsF6yID1yR0yk9uW
+E7AqcPMEHyzDIcmKcODZgHn5k4RdLKI2QPaaQEFSxpsCO97cRU6Lx354d/b
I+h3Pn1Lk7FJ79XqnbbBosnkjvg4s9PXzv6AnpAAgcWrcsD6UqJzYFTlZic9
O+W/oJhr+WL2Dtq4xHG3GP3KqcmG2Sg4nFzBLlRzSYKeUNgn/ePlf7wjIN11
GPg5jd9ZErd7jeGUXNKhXR6UwFMab2xQIQT3GbD1wGZQEqdUSOTewfLrl9HB
W+1bvvNgUd/xlDu6bknEtZToSRDaBk8VhP4H5GWX5PMIItiIhNucTAUoZ8xE
Meh9cNXiZ0tIz4UzHdSOdDfuMjSxwcZZ15ODuMNz/yzHM026KmjAXGZ9Pt/9
eMiI2PyN5uhvtXgU+dm7iit00lb69rfe7cjOvboNbqOa3HS6xfpmHUlmE7wG
u0t52+RIYLxNo2ajkOCGOwN2V2sckYwnYxaR4E8uf1XFo5Ar10y42T6hSl5r
iNesaunBz5iRMAuYWtZfwHld8t8ntoV3ZGncqBzCEI0A1gvvtg7X1HdHLZlC
Tjq4WY5LUjby+FiChSQ538oZdwF2+8W+BRFBnPnGl27Aqis1qvVMazlTwj6+
ItpCSMfo7d/blzXWKEtTltcCuzNrRDYY5sfzkyPuuUoiZ79XI/dnT2DflZ/K
zvl0WHsDM6d6Hp2VKzGj4vs6NLfQ3ywt+G2cpqioQEJGKW8Mf+lI3MXSNZ68
9n9RrAsty70XApTC2AtLd3nJZvwhq+yX1qX3tT7st8E0Z6bdStT25kwvBoFU
bLY8cz+hFxJXJJMKdtaGgW0df316I7nuoX+yeVujF9TDOXaxCteiJqqL1/Jp
mLXn8ugnHG4aC/jt2f99gOaxNk3jA6pqxlqWw7TglkuhD8ylMN4D2sE7k5aw
eSc6EvLzp8zbnTAd69Lv52oBBkwzMUhbTJ8IJ4RKJ4ZcqkC2K2+q1Ytf/6YV
YyNSdcWR6pAVT2AMEOmgs+IOCtkJ1IhFyXAGaAUciUk7chPS2IBuIf3+R2Gw
burx6OXRYX6U8mpst99EjjlPgIb1dNgIYYbJjnlEl0w+hGQbWO5I6lFVQPkb
VN7BOhpyp/zSDK6Iw1aFyTGzI+igb1sZOMo9bWb+LYw4M+zrJK6QS78+wm/o
rFEWQm7Ey3enI4RD2cmrfOg8Fh/YIAh7VUeQ8mJ02T/fxXfdaKTsM2/6Y08b
w3e6dlvFyUCXjRGJSlY8M88ZDZ/QbNw7FQ1t5l8ww5Bndqb+wuCj0/sb9eLS
cSS26YlhAwoGJcnFPPoKB0SP0NTFVABpk6pR8e8IfLgy4hlkxjKlYBnbs2ae
eS2udr9awzxg3bqaFBR/8L6vjZzemLSOT4gL2dqE/GGbhTBV8dNsdxZGz+hQ
koorxerlMMlNXEUeFfnku4UiQi5AuWXd9i+JQEEVnHijVy8YorvLazcjvYC1
FDzlzKMS1Ll5AwDFTjB7RnOZ4Kl2UraRGDhmFoVujbCVTX3SVZxBIKQmyK1l
3ltn3ebIXk7V0jDdqUi80nn9F+WVspkU5xMTvuCofWIpRB+N99JXmo6F6u0h
wQn0reBPf2Kaiue7sZ3R4PJQLJPo/TNCsJnujWbTMk0MhiM0DTQ/qQyLboEn
ta/MTW73xM8rryVH2EwnD8L8J5blh+5dE1fBIgWhvfxl8ltZ3Zp2eHY2crxp
gMe7tLuaVIhmMYCD6b+Lo2/00BYN8PFIOeNM7yVM1IP5JV/SJFNCuSkFsnpw
YDI/BrNpkDKYuoQJPbZJq1ILfvyhFsPnL/Cykz/KRL+FCFgMo98DUpcACRrv
X/I2dY0Jl7XOaCzopQfozWoOFLNPemKuzrdQArBijFVO7fYY65SxGRbQFjfa
0ccCQji/TUJRu5yQe2hjc4HSJCV/qls9qADHhMa0jkMV25Lt/pXi3VPLrz2k
yCRWcrxSmfI15um4SUs2SWltUYSGiXTLaUAoMTRn/ci1b2yqPf8zki42/75m
2A++KLEnCtFfozz2zzR/bz15W5fQmVcIgXfVrIeQAJrQJ4l4Mi/qtSPsu6Bw
8/6vKrnbDOQDCU0zI8VsnNDylXQDH7yUle7EbcmCz9qQR4AXfg3dolmZxJ43
I7fg5LMUvN2DzCrt0X9TmsTUxvZbc1p0JlAhngW5HAMNzGWAauCD9948fPlu
MuKaYl8yke9J40qAxtYf5dWJi7iS8H7j6GFTMnDswoWqE2MqWhalWU4PH6St
y7ZV0B/qvGNeEbI/kRXV/O9GYBNPQp2gKB7sPYLCwJ8cTQ9CTuwyMKtXgY+b
YE0wWzBvkxgOB6AWdta98Z2YjqZXjiuADz26nPLv1IsRS1lykqIVwfHGhc4+
7RZn5NS6eFPCQ48Q6uBseDbUnkHnlHjmOWcWjm3Wvu18tF/WPDy2kIabIhuh
y7PQ9JmqLt7A0wrWxOV50JvuCSW8dVQJY4n5pQ9bOw5eObbN56n6gAjyMIox
yJTS+jwHWNs+4UqPH8hOrcan+UVEmZFSPIcg/UHRRrxbWChimWPvec0SoVkr
kU9PaFPZIwOprlaKYXd+czzrW3FDjEbd/JcRdCrH45Cpc366cVYRIM5bysz5
2D/fCgrF85oJq+afse1logR/7wuFj+qFkDTKbZTKvvsnzq/JX+1X9LKRsMmK
H630xvRhcCY2kp+StUpjgan7C5qN/vJYN459Izg74lrY4g5xN76hrsXqtKDZ
bZIwcBu0kEvL4iV6GpOd9kIB2DONv5N6DNNMdXTxwgFvXO3RsbPM2440SvUA
cvyVOORkK+Yzr9IL2sOPg5dtby6WL0esWydAWnBgKFZPlj21qI70V1L5zqe3
z7cB5R02pkglp8/4q5+2WydE1aYEsXakmClDuRJitGQyWGgCQSyHdUKrHamb
pJlJap07CsUY/FVq/3Qc/NPgJhR4bzgshuP59e6dyRFqhPcfqXGmCADagdED
cSRvriuJshZAOeaKuHFXoVZecSkut8ak5CyHtY7INlMzaG/K7k69Yy/x1VMS
1NMwIqZrgDVr1o8FmUSScrXQxYacXOIbgHSmf6AsCv2LgR/xsXbTfV7viFcz
0jz0jRVOon44AXILbMv9GCCWHrk32N+wLXNiasxPSxAwu83AyUFnoAd0B27b
42qE8OeueV06DRDcX17lR8yeWGTxY8WiwcXLYjcQw9JdzPzUvc3KkMPZR8ID
bmahf2v1mC2/RfJGAIi9H5hlM9c++xH4pvnzgn/h6c2x8f48FxVJAVDSukXO
e2IcnDAsX/pwqfHF4TBzKs3vVPcnmmU/mx9LRJW31mCmSPlZIISggNkowBZ/
r/aybRiUeJ2hich+CWIqUoLXD/9BFwoVnS1S7wk1eVxVcw6M5j6oKVmu+H90
JCUlLHEH+XTtIOBe5b9yxgyCwzZHklwSBWeqXISuCBHptnOWVvvbymbSXXjx
W6+8b3J2GmQ4Y5s9+QJ7nqrtHha7XbYatYxRxF5M4ToFTAqOJW0c/7s2Kl8f
qt8KK4Mns0a7xHoYq7OpSs044rfvwxEHHbgSxIA7IxqKLd7T3aYObQor8mwY
p8cV0Ovo9yfvknFZDTH7nssJuj4URkQnWfjBFW8gmu83mEa398SY8DJdgnFK
H96TzyEecgC8Q6+RD9u02JmerXxHUgKCRy2VQoGS9tzIC5Ug52U98WhC8NGQ
za/EwBDxwlQZLmRfoOeU67zwCeX5P72Nyf+R7Qno0Jfj8zDcDO6Ynb5AstkG
EDt1UvHhKvxLvrz+QCKZHsXyHkbeUB10mYKJcYWxNEQtFHEo/suV3EgpRDtl
zn4b8o80wBHlRV3vlRCeApvk7UH4A6UoPL7V2Wo2ekHG8AKc+6otG9s/Ltht
zk/oASn+J6jAPDR+gGrCWJLlWwJcP2qGZcFK9gbuojrzaqAhEzbcdQkIb16N
biKx6X0VP+oObasRuZmGcrhJyvLQWIlaj2kO6pdvBC1PdfNwZD6cIwhnr1vo
gWVpy1DM7v+W9IaurEKgHU+iR376ji+0rOthi3Ci9hWzdm42Gqyg0gWLSo77
cVXw9vew1k7YqjYBXz8e1JtCZnvuuE2WQIG3yCI/AmHR1p6/ruFC0yjD389e
UpFXSjzxm6j8yje8iDmsAUhKB7mt+HUwPCnfNxo39LsGn3s39KbUPFIRhN8K
dfsHHF05C6+G541idB3W7pr9qrF3qCFpsYpBRQckdS3gzmMV0oFg7AefntIe
KX7wh7X/oAgqLrRsXRfZ4hGH8kHkqV66+6U+wEFR3nXZm5hlL8hrOeZbfnOw
/mGUxy0kMgiDk2kWfQlhDBpcaNQwaH7UNFPq993FGLGP4Xvvt+QzeNXKQVeW
XZY6f/QEOTHOdzaPj5aVRPvxNzVbllz0WTmZlJgO/6LuM/N1IDps2Q6zMy05
e/zX7fN0dZDavX1oBayy12Lh9CBBXX0uz0aJdUAtyokpi8D2VuUwv0q4aNMb
0LD3NlgOGVwOzDis9XpaUR5i4PIQKbICDNcZmXVDsCr2t/b4OF2SLpq9xHfx
esXsyQjiHB0jmFfSUL6gsY0/aUrc6ZmFw9lkUY/r5ilmY1Bp75rnDRp5dIlw
VowOoVDWWOITrekvJx+CPI+mohI5tsQAPQD1AD0FD3ya37+0EXfX1jhd0c8O
UhNfWKKK9vK42YXFoEQRs53g915AvSnfylJUjS8fIg+IBbbXjZzZosFjePm0
3zIPxgVuyxWdv6lmT7mJw9nYQi8CB9f5dNnT/CwdTnGoM8ITG4Xv/X5fBXH8
xRhPCoHk20OakWyrgQInzQgmNZjHwbyM2zLEALpExsBxm5y4QjpcLdk5f7GE
c3I4DtK0AEOLk7wvhjTvaRUjRXK2S8ySJqk9g2uqMlrjB4ZmKrCgAWUrBSy6
jZhk5nv2eaqComVp8xWwgANw5Q2pzK5CK8NRw/ahlxED/lommQk5uy1V6Qnn
JGQosNz/b5oEOFhqIKQT98aAdSAMgpieggPAgSzZexmjYvptSuDGdeKxLiMt
JuAT6Jl5T55PA6otNyaiVLusan3oem3LVu/c3yrRqMjsHMvFmy/cEXnZI3B7
N1llqDXIhyp4qH7dwuTQjGDUJVOr/cd/TFtycl55AAPhug0TXE7XQYHrHbke
a+IRpqNF9aF04On2VYUE6PnNjgZILPpbDB+M0IbFWEgFJncJceGGlMtMiszh
EohX1fENU0tDpFAYhE8rVWFzo/VdyX8rCvqHk4EIuWlY32QYiHRVll8HTzAM
2DpKOTLsQY4XC5wZqc1kLEBfm9qXu9Arrcya3t6LNSql1L2TCVH9BRwtEsXq
CanEgMmWiEDVsVfcR2nutU14AGpETZgMuu4+cmBwPRHQY+O4erEDD0POUUpl
yQe2cDJ0ILGI3FNWqKxnymGAzM/8yp7T7CKMHzSHAP/cXdroROVHpx84hvfG
Y1icJYO1JxHsCOQVwKGj3wKrrzFUCwpqaH/EvdFg8OdKPI2cen1Z7iBVYFff
+mSRns6PvpWjevncAufc5xYlvReSVe469Jn0yIfsbxI6Nq5ZIfN1uwp51KEu
WUvjF7bRDKEH7gyPN7Jw/alR+qvmZO8IxNdhgZMv29crMmckU8ng+zu3re05
OS+6k5BGLtvm2D+kLT2MaxBBllSxooUAaiVXWM2zY89hSXUQLCzmPZFCDLp+
4gUcQgd3GMRBcpWeud0g8kxNATmhArZqNVOb60ej/Ekt6d7aVTqVOieNKSNH
FIFfTQ1oZ0NGTpS7V20/Fz8+KFei2D1olF8gRcSRHRFQQ6G1sqSdsaIZR5/b
J+EQKAVXqvviTa/M6Sm92/IXirTN8sN+a7J1xcIfSG/jbtYn66sg5Mg9ZjTB
0RhbIcs/Wtll6gnO94pgvmT4wgb2R1FzsesKc+ZK8aQ6DWPeRDg54yPjIxrZ
mfOYmer1Z4DT9i4j/PT7o2eiG1onU8dCe8Qkw9s3XmiRoG8Yl5eX4Lzq0+Zz
dhd1Xk6ihhTuHBAYyV+lYRdlxX43lh3LB0UU6E6rl0Gk0OQw9jTk2ih1rW5G
yd+tB9ubaUXKuEfcleyUD4Jv4UNatFA9zSO+egt12/p2s48GD7CrHcSx2xk9
JMX61EGN3wGcE8AKKqq6JCAJZ6071TtIMebeUp/GzFvYoNDlAnP7w88yGrX0
xA1lRXYUeHxrNDnrUeuhuOPE/w3NAVtRr5pzZ3y7E+oOsz69Z90LzY6N3RVu
yjZuRR9wDNlHbpU8fozUKcvrt3DDPor9HdmGgjKPT+IEWYzIuRcJGVg42EpV
8cbAhkh+J84l+ETrS8nUIgMrZelTVR1TWChNmtuEZq+EiT+NbWrhzAYMjTJs
tNoJt1hhP6kttNSc57iUUefxggksDKcOVsl2AAWunIYGTF8hRCZrJiLoLCK9
KWVWYd6dPTjcHZMNewVnjUT7fucgBffBC93R7c3X64rD6sH0rWUEas2mB/BL
wT5C1gr2SDWtERovZ+FuJS/0ql4Y4AaSvG2xhByLy1AQY/NSnuNDn1ulqwfO
i6I3RNpHaTGSXw73Kl7O0iTeAX61GbkKy196aCjKZ6TB4+rU8K/NYp07W9Ak
ByKWVT09Fi3fQXT6j7Sc/F51ntPL+NCZEo+Slfv+YnpinFWr2uImh8ua8y9j
xKnYcy5tvx2vbBMBpfTGSesi+5PUrU1uFcn5nZ+eZexFUOgzbj98UBoMGHlR
HF5arLh2CkAhCQ7uWDj4KcedxLxEwUFEKVgR2kaTaREC7KzI4JOsx1ZLIG8I
TAS/gnCrq7DISTzSO3MJhNs6bJ52IowDf58K2JGW6xy6OYtz+jsSBEHM2c2K
zVjmolPANmiLylBpwVMtTasQRlRLmWb3b6nf/E1ff134q0qlXVy6srJn5ntz
ivRbRp2maq71eTW9amzxBolooGUStev3Y8lvdV1JnMiOwhGpn/Mv8pU6j/Fo
c0loo+rPu3dAex/Q876op9OPwCFzbNghI/18XQyL8t84ZkdrNZC9lESpZT5y
mu1DXxcgx8CbGn9XU4NQtBbOAulNzI63LkeDYLBqpHK+QYy+QvyZng/2IR+z
5TyBlajVjHmhB4zVEvgnMrdNbkfZs7ELbXTzrPuyp8BLxlZaGXUafsje8nF8
Sm4y7b2eaGihTagyEiJSfOnh1+GDbaSjlXu7X/Vep4m3adus311tnOITuvTd
hjKxN72s6RQx799by37QNREwfH+4foMo/ZYWVkOG2AmLtL25ZAIepPq4AAri
Pw0bN8BkvM70PiB6+gTkv2EBTdoezGRWtqxD7+YbBNOt5l/PSj2GykT3atDD
VI+Vns48tIxCSvMc7nU1we5/QnQlmxZx//qjTl5+3lGV3sw37AY9++fLsKoU
4pvhkttPY2ZacnfuY38pnipq/SsptfZbpT48/PR4/cfWYJD/+lWh10o+c/uw
ih8sPJkrbEzIkxQZBk5ikzQceKz1zATHIgi1sFO4JK9lvljWh8XbhlH2jTMq
ooK1eIChIidFZ/26QV8LWuR86f40jVXgp5zKcfTjCrxMjiHaa9pGujSV1R+P
IyGb8CtXyPTW0X59WQtM4AK6lIrzFewSCc0Bz+d8tE3SbkIAzoKMhi9buOfn
DY5SRmUdCQc1TWYSq3PKQMbOrTMGPEGqikjFxD3IW24dYF3phK8qgarcG94m
t3HRPqjueqj1D0ovX2PUX/+OjKUNMmPJs/98mSB24TBWkmRaGm42NnQPmuIL
8IBNZTTmB6cAaH+osVWEEj3/LVcmH4Hnz20ybADBby5bB1PQlOs0WToDOxu9
9AVrZxDHTtBiM3q4AK6B2roGuaKgwnV2bz/9uMjS32RnQqyXvyk5RZuPry7w
Oa70ufEhQZtuPtSg0y064PKup6fAojfL4AMVtOtFK4YhQmWGKLVCpslxJCSu
xdQO+g/PwFYfpdgklUB/Kg665OO0Mk75e4yfDkxhG50QEjJP8v0zIUGDk/U/
ty8DbP0+6HCzpADxuu337qBAktxfsX/RUWW4PbJS7l0rg3p8SEJb0vBiamgC
Z7s5gwnJqEjtNIIWR1yiBH+GLdopiyhO4+lH80FYBv9TNpngRlqArnvtlFWq
CqnIIJ+WoQge+9wSJLkEASE1IvPC9WrX5Sz88l7GjKQyCcKta81CMdXT8bcm
0RmZNZnVH09yEpwu9y5M26MJBFcPe5UI2Pt6QFHz1VcENqLI5zh+u1sFUEe4
6eJtr2wzU2Wn3g7WbiV7eJum/R768deikWiez+gLxFcOAJPn5wLp9sWyv3rG
SNd7m79GGKfIXeEQi5X6sdcdgVMkD8XV4f9vyuoSofmhqLQUYr9BUBLBQVJL
fuhTMrCX8qjgStiybn5CeaJVms+XJUvwK2kUVHRa08A4qkROtsm1PzRcgkF8
pu9FDuKDeCfpzzjrX53Rim661Ney+6WQm4NTduAzDm/ZbCFOSbwJeK390NdY
zzt85CKrOdwxmEea9ucA95Wca4Wo/PAkSNHBQm7Uu51QnAbZbjTaOjskydCw
O/XlWbYIai3QewP4ZXzDoZoVi0qKU7s+65sGMbOhoHN03o6ioDFwR+MnZNyv
5Hveq7bI7iQgIK6x0nJzoOOPeEyXEI+UFnNBZKNth7FktfBtX3OA0VlTJV3e
iMRwxNGidZlJo9MjrhgWLcOniwmKGFlzv43cVBEG88HI+pMoSUfIik1tiLLr
Kl6+GiuJ9mDyYm2dey5PZOxeYnTS3U78q+M3vbZasICrv5Irw2RAiX1w3qTZ
3mFLFo85Vxyhzx17pFSKTxUym0tOuDQk2NeOdGXxuKJ20rTR+vf58RSgpA8w
ZM4eYeLo9hkcGgKjeCCTxOF81djf3PasCHTOjoC3ykWZ05OcHzn/uhAJhSkh
szBqb2YrLoZO9tZggDj80nhTX5bDK2bTHAuI1PAF3TXK+035YlOgqWrb8kVb
CZHwhfTXK6zlcvtLlVTL1QwmDSn908/ViM0eli4FzrApNBlxT1hCc+bbJRDd
0Bi2+J/JhQdLhPE1Ug4o/npfg0cI5mB3KY0n6EFOOaQK8J4fNa4I0XrlqA3B
ZxL+sMw0Z+l7AgccYD7p/Vsb0ncZOe7TKATaiP92WrD2QpSKdwmaBW97txmv
hmyqGZpd6e6n0HeaVqTAI87vI822ddeTqME5QH717wc5GehzqV+ZmJpnd8y6
eqcEbjkTCpJc3cH8GgqC1NPcJDS0DcFPB9atWBi6F7pU8SDA9ivgn+DchQdk
bNuWnp2GnBHXR5tDCaq6CxwWIVf8J1ZUQ4dl/6W6LjkKwcQjLBjyXf4X9Ihw
5GhJrobukzQLqmqjLEdIZLPVuUrtEiM80cPH7XeMG8Ll3USrlsZcPjOf+Jqn
0uodLtrq3Vnqj3/ti6QuXL/Mg5e58pFiQgQ5mo0aV/YZuIYPDLvz7U8w+zsk
wzBDFfr21eDlezX3SfKD5f3HXkSxVY45OgxHxQT33YARuHNx4Wm/BUJfYET5
BAN/C2bJe1lKxiuuk44Y0RBFlcSPRzCvCRwKfPIFl6oFxfSO+uHoBqokhKTR
Jue/wgS5hZfdwMpr5nDCuxwqcdBJDilr2pXJZuQqGtKedRmexz08RViJJeYc
pvBnvHAwUFQdUrsO/9SFz25nc1+VVWw0JxBYuaV+xGg544a3LhS8Y0pSAlAh
BbJE+OIhyjFCk+DbwJjjBrU13ZlovhZBgRZ96X01T2C67nlhoxOigNB3ULXe
di4lEfoHVihVKXCJgsSc5I78oXM6Vd4eIwvLi1OFyw46VMKZRmRv5Fap7Wcv
1mvHhrPoLYkoi8gYX7hKytFt1O656v42XaynxfMBgmTjMpPwBQE+rfZyoP9n
8sw/uiH9IQ3iVaNU8gbVnQoABjXc8jUl2zT//G0wzlB4fu4GC2WusQfsJslM
P9A7n2/VlgE/5lZBUQNJD16RAHe99C/kfRJytGnbMgR8O4goXztptH6KqXPF
BP5EmZ/oivJGfRTyAyf78PaI7rJpFjMBSpdtjzuZJLKHkW4SHTDyKDtvv8Ol
Zs06efFRJDjk3qgyxvcKTbGCYWSfBnIhYk+9YC2cOZV6D8jzwXW+IcRmTNqb
YAMxMhiWCVjeAdO9RaZ/sSEnOf0doaXBo6VbltxWJIkxUmT0Z5uZZID/RmKw
W4iiCZlLv+++vFDZcqV7b9bd2fB8EhLtjZNPjqgByxArSen7WwT3uKTieXYM
6/bvWLOyOmdPa0iBEmwf+LeV/glssJLBbUf6J6RrvGGygIQsG+e2rWGvy3iH
v4i6hzcvTPYBq7g7KqyfwAxtQWK9H0Z+hWRbuQoeG5AwP6jNHiCeOuYoBQdz
Vd87MMOCGWfew8VDtqse9sKRywTC43uIC4UdHXALDeuj3NEZP5M+hAKmNeaP
iSwctfpDwJ4pWLVVSe/qmizL06fjHPLd2AzzsUosXDfy/rWZcIJhVv7Dz7tN
u2YaCNlYhv7sNpIXrk4/6G2QX1hfcnd7eM0aDaZk3MFLid6Ys6UJAi5+rssa
iuElaSy/xnb+2xh11ww1T7N5uzFPEWxbh+ZtY7o7YVxexqDcZayS7NLY4woA
Drnid/eTuX2phTCd36Kk0kmg61Rbrw2MEnd2DA0/PaQLrXhsb7OSfgRYhNfP
10zId52JafvomWPUQnYq2snmmSB3imazunHNF1igOREIHeMoVyRXIgBhYoOk
OWTk6L6vXblhFozEmL2NKfE3qBwSD0hvndT9bplB3FpZ5uY7TDwL5WCln5Zh
0PJMhXV3z9lROFZ8JzOFcYC1QmeA3Ve6t1Kt5+g4leItQ2L5rrTGXGhJTxnG
fjkA1qkfwUN069dlbsBimMwfEb2Qwp1Erxlduf3EAYulDWHxMVlnZiDdVtMR
hKCRglODrX8+kzYGy0vrEOlfgrh9W5RqQhYlb4Vbo5aeHXJFYMRsueNb/1FP
4LoBhZ4OtBEkWO5Jbo3KDm0iC5LDIbahDnSs5DhLYxlKnFhlCPradsf/5eXM
qPxcc9ILY1r0oUWVNXf3v5G8K6/eCSwJgOOckLyMDOOq8Jsu7CvCBlEGSlTZ
LkchHY01poHU3xZ1XHmbdaNJfHIY3bJqZ1g3MFm/h87XkXGUT4IPCZl0TGeg
3/WuFXhVc+q3i5QX3o3hHAwaXf6w/6N43RD7rDDPwPNmpqJigdsRmBrc1X2j
9bVctmW+APp/wpB85axjdI88apGQhrjlYDUuJlIYSIDl15aSb+hU4i7qSCrK
ErwZRYQRjuoaSd1zUfgYRSrVgvaDvdiTD2PRRONA/KYvpjq4KfzhFJcH9UB2
8mqXSxWCmS5EFjh15Rz8+WiyPaWYxMUZv86cAvbyQT9kVf/HdZLaWMNYEBrs
2mcCMupeASxajPVJvM8ERvTqIEcOtRhXGYJImz1oXG5Yctx4ccl+PLS3JoIj
TDfg7EXxZLJfu+i1zgeEOQBgGWdI8SVAXXdV0kvOSVCZAqj6pBro9SfGSVm/
+eZQ27q/wkT7VWUTWT+1xRF0LqsvmYoJySetaDmJCt8eNZe6+OQWHAeHZPVu
I+9LOgjbgHxvwT4y8BUVAg54KtDCJ6WWe3UU9I1C6Ss3za+UCqnPjdIv+lzX
wpRQYoONAyXM+QL2RKohr29Z7Vli0G0Ypelc9y1cslMQrZCSJ2JhJWLy9llB
BHx11EcLZIJuISHhnW4CYRwk9x6u8MF9mYskr/vMG3xR1b9EiaGqvlEE1uW4
GVpDRH8lZ4OB9X59iVZj4Gc4MwiVfeB8e6rj0k5e3DEt9PdHJLrWiPOExVqE
E02DpVk+2BEHZY4S3WGY3dBh+O+1EnEsVqu9YKVBhTZIbJjRyekjBrTuGo0Z
wBIMYQrrkz1PIy04d5jZkoKt7PE2fSapvsQ3HZbqQpIAPkUT4B4ffTxs0+HO
c59DPoe/9fMa7cL4uGO4HoaNVON8c+jGrRhgDUtgQ4j5RIxBr0z1vr3RTTjV
7Efu5BXj04s7ermaA6EllDRUwjJu6slJsKyQ3XmZexr2A2uF08EENQi56I+D
wGPjJCLUuvMBDP2XcYTpRri7RgAM3qBVan4+kFeKbnQ0qh71MInz9S4+BnWs
QVpxl4gCrdIHhAJVIMHzBVga8W0rV31B5wM8qC2oz73inQpyuYDfim8H1SeN
qFm5hjl0Fga2copQjWEREMBBSPHmYmGI2MbQFirhv8umcTfmt+SALKEtthF9
T4G/OP3eofbLSABgvT62d3dOpFbam9Pf/6aJonK+AA8hHa+bmh8QLTrGX7bx
AHk3AlJkhT/tO8reDTtXmw+Gx/b6vb/oTHjC+2uS6NViit8lqCT8b9eaMOvA
THRtok41DioCyfVgxd4oyBQHLESahaZ44uwwrIC7DRM4wTGmVl9gcCyVZJ/T
TCjc959ifWjWdzy7H1euRTybx1cW+OOukIUW8CfLVYmdYfpzlIJkXJBhMcmw
CrFhsPAufxPgMsgoXU6Fos0QIvdJBmUB80BDdeEM+osvrBqxCtGy/5kr2qxP
ADyVssRYdHe0grPFdLzfpnZC2CIS7nvuJ5JeU5WWaMDSmLHUrhT/Gc596s4W
ONwoZvt28WDu0lF+sOX4WFKBAFisogMl3szbQagMWZ6V+Iz5mtGTPWxL6Vmg
Yi1w6zLftE0sOz4VHqE7F6wkd+lF4+1vJlKATRbcZmFnj8DQiZ7ysQuSqSls
lFej9G/jTiqXpMQxoMY+f+Bq0OOQSHCXHpft9AYD3lCz5iwZWk5eVUVK3xTV
lSw16W4PVrHFA5acfFVp0VCeUhDVTk/l0yyVHlyf/deVGQ39Dp83KAtbMqCE
y5xBguIUmINloPons3x9kNYZBBduZSOOXZKVjYWGH7/JafEqBC1iQu98asTb
D5jR/XQUGniB6jAtm4E+in4If/b1qMkGEFpiSaxggRi83j19bUHEir5VYVMD
VFoxuX45FhJ7t/DjFADkEoY++NKykJqWys0HJmgbBFns3Wg6RPHbmDy+ZGu2
CRA66sNIyTZMCd/G6zOJ0KygySAQEvhqr5Erjo4udY9obkTqAuXYh2o1paj0
c6dvp9sCpRNk8AHY5UqbVkG1tRctATm6jQFIdEi5uS+X0hG8cgk6KSc7iZKE
UqhZ28Irw0LHj5vvlNSZN9AsV3trMnu7BOGnXjqAM5SjsgAYOKVLLhtSa0M+
Jlb9txnJMTCAxMrSYaWYAZakD4563sc/4bJ45Z6u/Za+3d//kW60WIL0mmNX
0hgQSa+/HPcOKgwwt56cXBz71HLEozTYgLwLe1qOn8Z6M/34olHfurgTfepW
uccIVClOcibHenq6dBysHIfoCm7mm8xymZjgqdOWZjeEw5i52r3dIpxpbV2E
PVJMhDDlDl7pdFUMdwv59+qaQyCVOw+WfEHktxA2jqcpYrPZ1uW1seMQmPVU
ccNvrbOJsg5UrAyxP291brpUhRAci8c7c7bmr8LkBDYbO8sJJ3tcNohUu17y
Jg+verL2U9gKYD5fvBfm6j4fOzpWCm5NZetnxJKe+4NjLYur0ZqF1NHbTlJy
7/svAVZuGL+QObfzA4qwSRS1znhQ1SkkQSAtl6wyyAb0sAahELkFs6NNJAYs
5Y+20cxa4ew2ghpVnkbBk9yhadicbJuPfj3tPoKRPbmVA/XYHdhgR5J75e7T
Qv0euFqsJEBDuNx9tSbUJhuSORGzx4W8kN16vatpeCCw/ctnqjtTBqBkVNqw
ay1e/Zys+Uy7cLPyC1uftc9ASkmoHxtQoa9f65oyQsZ3Oj4FJL58JdkK3lRV
XPVqO9Xit5+4DA8RAoL4VKIkJ+UAcoOb2bbroLiD2DLPgQ/rJzmIefQtQYte
7ki2kR9urq0TfssXsGdJKyUHfxUKz/LbvfQOIO8h5R0drp0ErSR4OiNGtWj8
k3utMS22RzWOKISOobZXc99/vuT5R4ZqsdQ8NcoUVaYzV1MxgXrXBrulznqX
5EL0QIZoeI1GqlAq+W2uHCNjoO0Bn/u4VUdkVGQJLazijkuq30T/OfV6BMiR
hF+MPmuf/3HgpBHFtcUOOjnugfKG6WqKB5wh/LaLqQFAmnPZU/PW+mHdti9G
yge7vN79fJZHCPV0BnOZL2L9LO2Q6AdNBIMTCmXwjawaPbY+b5g4vi1XNIbD
XQOWy5xb8aeQ4pGhST1gH4BIhfsK624gZ6aHpfwGrDfX0PWtvxKgvMA2ljYA
svFO1454DMrO3ifSIXcqfG7ZxV2gUycJVm2y/BLOKRY9qBTmiyP4liOqaXxM
KqdKhRyrjMcfMM5jJ1yLJZw/5eME+nYCMUlsr452XsMpAxb7Y9CjOdry14bM
iFPpTdS7tQU3qYeuF9KWuv97t2nChc4XMBAJ8P3NGwnGwdPRTBoPHduCv4/Q
7gqCYeVJzMxFxdF4h1ZyVtm2jbrcL7uBD0R/qA9o8Fo8CTMjul+Oik6DXlEP
Zhio7meWdqqiBoZ1K6MmV6QUrIs6d2jkY1K1xnraJlbV8lW6wjZZvKlGkh2o
CZ5IBciqocywGn6gIOexcz/2njYCw4sr76plgJk91u+tNDJ3JRJNDLhMWcF2
b159zTS49yuGrSm0EX6g0jev7uyliNlazwp9lLk4hpH0/ovoafSCzqxfjVwC
DqwC6qR23AozwhMGeieQueaKevL1o5CNfIXrRgkyepDMa31goIowvNiE8mf0
UMBFVVi2niw8sf1OHTWkeVw5j/ko0f9zvLLFfg1nRQ2zVVuLgFNCW2w9JIox
ugTVSPJpKOr4NAEmB2fzJ8N2nss5trVk3d5RaswdCnMnlbA76G092lIs9rz6
tE/XTK72skdv8nJBpgvruQpAEVwLLEzxoF+cuJWaoXw51k050bobPvuYG519
duyNUwv4sFoe1AbHOCNOSwQiTptzhyCd/UUSmuxlwQ5ClfOWaOxgOmusHi+r
k0rDgeuVglxyAuVSJO+sYpf/mQDJxZgugyO8DBXhfzXPxnZbXzuc/YtrVV13
1SVsHi7xQGV8KMRFR+KgyPwZ+MUkfnqeTGyFoDGnOx47SEg9tWiQpUDNGsA0
RtK5tFjdJFFALGdT3yc+G5Q6AWJda4qPUqVMZ3Phny/1bNmK0+LxvnhQ4z8X
UlP0Fdqodc683MDK7PY/KrjAZu49lxYnixLcZjecllqa76IwhjYf5wNUnafk
3+po8TIleufaQb/pTY1OJU8bHGxBNvAyh77Z5dsOBZVeP2v4wmI5qU0F4vr5
LtzhfMXPGy51uutOxISwlKrek0R41K2M/P1A8VW/rvLOWvRvJ4sU1dYvlA67
zdqoeb3YIAkBnjzJx1txgxZdIEumE3X4Ubb+343slQlYYPGVrGSHYFj4cjoN
mMZQzO6DmJW1GGuhb2M5JDi6x8m3PFNQw/flTMTNTndt+KtK465QzwvnHui4
ZL3Qx+S/nqeSAISBz+H2mt/hpdBIvJ5UabY1n18bMGwgVcZMrQPsAnFVwHr9
l0xd4Aig92nWNN7Tdpr2FvpE1ZeqxWCF6qrhMCIdgPA30BN5PqwU1w5LG8J4
wwhf6QVwH81MUqOK4MTz0xiavTjX86Kh2BM4XmLr9IGxXexrtGdH3GBpRMaT
36BHvrLwGushFuZyhoMI+i2ervUMgO5UQGSfcp64GtpVQrCFbt6j2CT6KACG
5cfAVLoSycq8OEboh1KfPucxBE2aKxvCmyl9XJBSssEtKwAERhhHhPc0l39d
bGiXv0ackfZSlcVKqb4bIro4Vuf53s3I7In+YZlfnhB0pziT76Sxilh8jNHb
4QyyEvDKQARqLoicj6YpC/Qj5Dp51W0Kw0E/fJJvd3huyUWxqBSl+8/ueDOF
ieebx75STofmIl4Ojc3TgmDqGbtqWusrhzcepBGIHKe/xGkqRTmHWZk3DAvx
MqTikwPJh5puoY11mEllManYF6M3KLg3Zfw2JhqTwC8gy0eg4jjOWUgFNTY/
IxYZL0WOfAcyckQwh+1lvgMZ/e1XtdOz1F9OehZQ2XkxvRmqNGD6TrbzXwgP
0tqcBzraqm71hX8HE8gV+hVynJTiOKguTxe2ma1i3Fxkd11sDxYvoI+YTFJ0
WnJ0+m3v1rwAIpPx8HuvBYzC9sOf5AG/KqwkFZL9lTz6zyUrYOFL21OkzAnR
HYpxHIzEfHA5mnAP1MZ0v26UBVWe/2H66UxE9qoqoupLaLP26/UvX+bvyBx4
sUAJXD+RFrXDi2V/1tEeLw3kpegCkRS8b+j9mmraLWYHX2blQBPYSfayD56H
KMUrtj+tPOlspz36YtfQUiMU8vdZYuN6W8zjwC3tlvuaF+bHGHuQNzuAcLrc
5DtJipQAe/+uteDZjBBbJF06D/t+yJrZT+STTQzjxfPJKQL3KceATEjcoD0H
IcdN/B0e46JEZkbQkETIv16dA4qbvWG6FOogqmIP0jo4Bl1k/UpSd2CCpJ1H
gQOU67bHnKPI8fu3WL0FXVnxV+YnJtxcSwBthitmVDt3q4NORrXisIy1ugwJ
JQxavmAQqauhJC2ZpNRIn3R5K8P9UWQlxtUaZvrg+7wrDgzRLfGJmA0GIyIK
rg1Z7uhH5nawoWqOFsWI8yLrsZcBrZMZt2oMLLKWzKQsRdR2HCDtbzqtZwOI
HoJTL46MPM3tvnDsuj/gNzUW8kWnFJIVQPBl2iTJTbSzqSMmxgNGPQCVTOdB
+yYEsH+QmG5AwXVC1DmMet43Qq3jpSQjH3dMeg8id4keF4uwqexFSS3xs3dY
nzb6CmjKEcYWF+iaHi7JL702ad0sfP2WTba0NJZ6T2G6Gxc+kURcYoFDh9Ix
v6SJgxWXGi5bzLE4BRbk34c5ciqyDR7R+cyRFA//lFu28ynGQUY1ZXlY7mBs
Z9n8I9xa0sDzeaYlyRgHGYwzBFRqhIPI/igoX+qmu9yzeJYY7xkYYFTO+EGW
kTv0eMVabNtH1s/KGlW6QGVkSCmsyMbWK/fFe/kWzMPmO1DFr7/rDr1mPqt6
tkEJYqPL6Mwk4PqR9XdcCTBoqNdoNmlzdi+FT1wx2NXoLKFijOOAduYJIogH
TtMnOl1MNCp5HokhNjocng7bDMdKse14f4Jw2rvHlHHjXyGaDBRzXjsGfg1v
PYDcuMDt6cwzo0/YWDjqkhW1B+9sQElxR2RdN4+DlNCLQasOdJKsHzZ+xdEL
rhPRNj6JyzUgl0khKBJB69kDTiVMPOdm2KDId622SAPrx593j3V+zVYBVd/4
jS15/H3Lp2k1cDdfrJTltDiSP+b8ol+fqdCvUydqYYiBsjZJMt7dIyj0IAxm
jrvN/JimxVl/2WnLjaEAATG2ynlcRnyw5+gYJ8gRNFTUgdMz3wLotRTFXMMR
b5dw3fZOfOAAb3AbL2ug95K2BJj6G1c0/g6S3OPIqfTgIQbjboacVzrZ0JHX
HwOPWNUaQ2M15Uj0z46eg+IHVbm3uyy7MBJCRuwj/GQThXwzYAag3O4iYCSf
L1oIU6BT5n0P0xRuOaR3vUEVcAnnKYuC8iOYz/HidaOpl2AprWdtCH3XXsKu
Uw15rmkfnJD3Kiwn0kJe7HEfXn74+OHDD8gQmMeuuRKqxumolVrCgLZrh9Nd
qP4lVGlfax/b4kWHkRggpH2jQnABOuzm1B+7/gtuAXmKHiJ7PsmZ5EUK0clT
+t1JpI/KDXQ9c8wexHbc0FNx2mXAmQ9W4d0E3YMkY5gvz3GYjM4SKKnKs9W+
b2cfhvcxtkD6OapwzjUmEwdkWzVzzg1hI2GPFPv0FIlSN0I4OfO2/7eCKMa5
WJLMsgxAdwqsprApy8t5WmoXxkJ9fI/1U2hZdTHisqegcbfjoGx7biYnzAhC
dMwBCDyvDGKGT8hdeQPhM6NoUBtuawLsATNox3tf2bFbgeQFrcQCCb7iNahh
MKRXAwecK6rpEofeTD6jrhVP72g8YD4haC9tvS/mwErrxPr/ZcoLFKONtf7r
Wmr27cbJIuoNaC7ZuEVt9M9/lwyCI8Os19hLWYUYO4V2lCINSnmzTNqbiBpo
4JMHQNPsBnrU6//nZdj/qElK+LfY9e1NqQPO/06j9lZHq7QSfpO1yOXxEcS5
nrGu8sMIk9+wNxyHyN4KTMVxjR9W/GxgLI/wAiaVszLSHP5YcZR8ytiA/7CC
gfHztboWrESE87EiIDLt/HQvjtJvsf2diz4fM8BkeBTf1tFBFE2NFhtyYzCs
4ya6sAmEEhp1rw70Yf/NUdARgPn9u4/LlFA1eVvzygJrXsop8PcM+PfzpBpx
FHKq4laBcXRg7/B8mzrM7T3RYMOi2ENrcyboSj+258sYAECxAY/EDRUyXVc/
40+Nn274rSjRnfw5VZgnaXuxC5d2wJ/w8GEZapVlnkJjW+dBjrdAoyZtuf2D
Nx+wjr15Z8Cx6k9aLMZFu9auxN/0lyIv1iTsac/unV171k2ESdaD1LcRgzR8
VqeloUlGE+DKKVon+e42T88N10aU8vp0ZB89dsC1PxqOVybdJLztF+vD+jRB
2k3KRAlyyiU58DOp3QiaTWofAEZMDZPLMKPJIsdJjXlr5Hd4pUXpkd1HSoUv
TAzvBtO1pwBzbuqR6QcXfU4pLaeKn+kC2wzE+Nen9M0/2XNkTh4L3f7jmdoG
H0B/5zLKK4PLdvvJVSK8bPyKF2zA8MWpSg2VWqO4VmYpdeh0fhSB8e1lhwtb
c7PmqSd/wdohTXpmIf6p918wsYqR8GehbQaxpQVPZD360P4IXCNqRdRgrKdU
jjdlxI0ZizLbMDakRgpEgzo3iCqjV1co0jTgwkgRyQ+JYwGRlgi0v/sykJrC
UMoMJFIQV8UIbotO0znjAmf4lE8t53TDRD0Ytut9WK7Y8471i9s0isSbt3cc
QFyYKuUU4djUEbCZ25rPux8TD5fLRIPfR1KEbMCdg+XxFmBfDgCpCv7W1LQH
regdEv5DYmKng598sEvLrjPKJC43plLzFoP1cptUbxtmD2GOvIXPizmuUSVV
v43JZyqze2N3c3b6OQX94lZiXS8eNcd30c64MK3J5Y1x/OAC54CnoC2C6cP6
jsiSH/XOtDBP/VPW3g9OoL1OanjwhoRBlm98Sm02aOqqYjdp6bcHyrJpScQS
AqgOf3O71KgCzhS82fnZDyP2jaiqo6VB9DQgUPwupuVT2o2LW2K8vXUeky0H
hYuDrr8WCAGSiti8MXQs28lQ8EqvpnyabjEU09VcNpiQGMVB16WigY19djBy
NVop/3dQJg2MCyJT+52IU5yytf64DPE9EQ+DBXs2M5RCqNZj3Zp6wtKvvZ0U
vDA7Sdr4g3sHzw5cssGjGUL+BTno+EganMysVSZreEZyX2UrIi+3ex/bIDz2
bU2AHESO56d1MqFHWwyRZQ17aOgT78nNlDU9g0FxdPhQrKTK0cP8k4H/0ilF
O1PudSSlVbcCnG5bLz66NFPaShjowKdVHXHxG41ROmyKApLutU0Sm0YHxcaD
wq/yINF8UetZIhxCrn8e+Ni4Jp7CTNTRkyvtnfK53U2vIH1J2BIvsEY+tSNp
zN3T1BTqealTiSp0z6extUttyGQGXFWGBF2vpm8Ax9f1nSwpJVtWzZmJv5NX
MoeMs6HQjB7sPAPzLsvOyssyxAVcj7DYcL9lGhCiscEUoZPBzTvwIsWgNpKq
6KHbMJl6XDTGNQTx98q9+qxQZurwrsEU8JBZcQMWt1y/FOaJqGMEMchFQXkF
/KIOzYn4j9p1TA6HFtlfLb1rvcSQBzwHm/XSMojwarnUZSh8d+9tutrbLF3v
8mkFtX/ma7VRZnFD1TbO7cLQp3jNM6VMZFLjmQlRlLMJwnXr1rH1xw7PH3MC
z3Y7V6foWzguULDyXB0PgUhVYArWIVDSJzng4zyp9y1ZfkidchB4PESctusH
JQ7/d8MyiTeldVKPRsWP2WdKokzz1jqlScl/sRjDmYhn8HqkvlGmwt8sRkjZ
0JP4yYZ1/QbK7WWKUo3HLDkdId9Q8QqvbXCScbja9RaWfXp0n18WAn5K5FIg
yJr2ZUped9GRkmjzrPAaFmOeIXxFq77PHSgFfcuwSkrc+iOJQl/JbE7Ytf57
ikodLhAKcUTZvNHh+qh+rk6L85HR+M458CUJOFmZgGlbOHganpuwa0G84r2F
+SekBrItYTwcQtAWUtKm1hgwUV8aebmlwr+epz60h3rSfvwjGHyU/6/SM09W
5rLnJCwZ7q3ZYfZe5MoJmXgqXWmutlnI63wfkm7cwVmzq3TW7VOOVwTKJLgk
ts/iYd4FtVW3R3bqUmGd7OQVgf6YP9TLHFWLY3ha51XQZzXoYZwI2mj4jfDp
6eZOufDzJUE3pxfuN6/2qGTmrYsYWrlq+nAjFlVo5Gs9vi078wb8e+yqE2qO
nnwVBnjw/p7O7ejV1+amvdU42nQEKEgMM0e6CuNRsA0uUrTCcsgtmeLvc+8s
QVZ411mJtYLYi2Z91OqArguzFKliMFcdEZ7w1ohCr03x6GFARTfaOaOYjIVb
zQ8/t6ZbQ4tqY+AkrhRFcOiKecZ6Uz84i60LkvgxJRgFK5ozFPr/ltiqjjX9
BHmXEFQK6U6wnCmuMkXpoQhWDXh7Ip89z5Bh9Ho8aWMeqB2GBlMLLzZzVM1I
gclLeikOrTG2PCPOBRWyX3zywAAHc/n3g8HSyK1nT1MSH1MTB4VJFgMaaMjI
/JR/4QvEMKhn8D2QGzsJih2uyZUQQwJEWWA01WO/KHCpSSPUdKyrE0T89aiJ
aLftR1p+azZ8HSP6D+0pPee2BD3ncX8OoLW4vvxH1saHmsSxFVoqE8L2ArTA
jFMkEgVTdSbCekyqL0UabnLHEfyupezi/SOytyX1K6a5VGrEUahxqquePZs5
rnHMr8SFsfiLpzPF4RKbnKxPR2NaOXjFti3A2NTnflXMktj1VM45OlATUzjA
PJailtSrRJR8kZ+KXuOT0g4AT36SBQJSCZ43Mq2imrNKRMZIfqmTlUeJJ7N+
UWWvVWR06GDmcLmaFJSUQi3E5xwqQmxfy5T+5i5MjfkSDYe62PZCGdyJ49ZV
7VY9rcCPY3BkcO82FcRdbLdEGcmBVzOtXVGz0tYINjhKMajXi85aVHk170b5
DAD8Dzd4NrkfS/8ItP57u1rys8JFuM4TVgaqiNVOWAAGWXTbofv2OCtInZgu
4rXyjorqKe9Nwv7tJdYfOtzDrukE7+sYiSiKLeL0h7DT8ahwvkRjkceEF4oN
IcNIGNtEUc4Q14i7X4MAQVwoYAajbGgqKymNKSmkbRog65tu1YjZ6L+H2gJh
dc9pEDW71/aJQz4JkGqvIb9Q+IeqLF9aqP4s+agBviZKAxYYFwuRBiwGNQGp
DC0irO5NJ7azqhSjavxpk+7KgUhQ6ltwNETPRnjZBPZ18VsYWmCHaoN4doYx
XjlnlR9J/e0P3jk4QBudLl36wNyXDIGuc+3+jFjm3jtTDHlht6Ch3ayjt7ZJ
i2RVED3XXILGmPf/tvZN2QKNGncbcPKG+UesjM1EvJVyN9w6/PLZY9+BzyUy
/6ZD3MF/HnkTQamcraIMvkWLcjVWggpMW7xCOB2JtJt0NFxWGP63FJN8D7tP
p2fZevnrmcBdPpEQdoffZTv+NJeF9/EXIhRJfvzFhmsvtROV/CEfku4tbeF9
gOMarGCcNwQIkiYkw85K73iOrBtaPvmorl+1+goVUGO6oDyCsj1IM0Q4YcFT
GYnWff9Te7cVikDIMaKp7vkYw3hoUWN7V8+pIniCKzHMxMtLtNwT5GIpzil6
307nVrHIwgcgLFOvPCyWMDR6Vyqoy57MhuhghQC+lpb8+CXDykm1wkCqRFxA
tPcBAcfkFyM2eYIWtcy/7TjNssa+anUBPe1q/6geWX8l7xBnDsrkdIL+UqeB
7mKVCODdiMQe/yA0coU8WNc8Vdfwuq2a5e5+HQV7NxdmhqjWkagQL2HGyYx9
3HQJ+7GkWsxxZphrNKJtL8aSnrr8RfUHSbHtDBFOsQOv0Su2LOW253szkV5R
U8hqJ/IsZQjjKlFNbCcmVLP7IdprS4uPWG8n9fqObvW83ncUHwNPdmofmXd6
PfWZjTB1HE/M6lQDcQgQcbUFwYgALyZ9esOBd5dumgLf8fqFWDBtupioZ7BM
3xBwi+vvl9g1lDuXuB3AOMlp39RvVVAeFI6ybsP3J0K0qi/FiQyke5YOLvw3
MCrKz63S+gafb9S24g5bFoLfVEG/nC+R4shN1lcfuQz21sWUqq/PWjeul15f
Va2FO4PjFnMDfSkhWUDofK8d5Bt2cU9u5rpyFuSxD39WSCazxuNiN/ID5MjH
w+AdXmZBbHHkhUhvB8ohnDTGj8dYIhlcW/Srcw7YVU4fWGx6o8E5L5XdJ53w
Sv4lsN5xe2zM5QwJB5ruc0XNTZwnigIo5Kk4NnErhD9k2HMAYOhvBGrAyOVH
eRCex9YkfJyRcvfKJG/NKrMmVYB/bkbMXmhPinFDu/s1NEbaSfGame55Hf08
70ukNa1CZe05ZVNoWm52ZhvaJMbbOHAfrYQxo3Jlt11+TiUZnElngnxUDeu7
szpvzBc9udxj3Qi/CrK2MsEqMX1i8zDIFLMNEFviS+d39uwD+sSMcgMwtAxZ
d3IEybHRrp+hktsVQkqzmei4EqhXFp+HTe/lZDhKjtq0VT/QGgVhNGruiatW
gxdnn3DqJUMWzb51uEFYfAWHao8e8R1U0TGsyhqyKAtixbkM50g+glDa9zya
5Bo5xMCgrmll5p4HoTrw7lq2CKSIPoQrmu5PT84rSE0mI+B0dBZG0SxzNNWg
DjacQ+GgfRFQkdn+dxV780hGT4ajVb0EM/QBKT7n/6skjYz2yHFVcRDvR6vh
LooczEvYKS079FsKS0/kU/kKyU2PXX3sFYuhTqO9B3ROe9YxizyxrOGwy9v7
np8jPivWvokFzXleGUDfapAYOw1Wjsxh6QPNi4gUdAe/+aEA+uczjkXjJF3u
ZOcEDn714mSX1X6DqrhgCDNUgBtrfNRdYUFJoCHdWgfirL4hgLn8hZ4RVObR
grdfxKeS9ElsrjE25U1CO2grj5UjrG7LRwA7iFPA5p9xfDUz3F5pi7kRCzM+
bHdNVyegz5sgoPg3aWteBU/Jv2TCpw9FdC/e/HLFTG3YhdSQd7aoSdZyoWPP
6eqisPZQfYgZpEb+3sBBVmAB7bsC/SxJCZe5JFOl2uucGDXGNM6Muu61U68U
ZkG6L1R1JC1JYgDylyz2kswXcfr30g8pW891Ue5jUGyTtKkfzPeqpkMUvGaa
798zoSvapR+Mf80n3J0G2NKZFuZmb1HzA+bTv/oJj97nzNZ7DwcT5/kuKr9w
H5ILEDoHIIi5mKmmL3wZwgenNZGw8pdxLqIE6hdOkR/4TJZ3vQUqNIchfi6S
18YyumnJty6UOhXgsKAbUDwCwRZYS1uRq/13NzOoJIjHGLPDFi4RtdICwPQ7
eutFXG7EcQ+jbjzEUU4A8WCRd9xklhsrp8E7msIiPJcCl9SfFiIf1gOSjASa
TQsuej4bkEmH4IK9l55IPL5VaSXdPJF7H1dFE/OoO41qHxjL4mgNiYo1OyXO
2zleTM0khrIG8WHKpCjKBkI/e6z3SGbWJldBReCliRkrbAkAKkaZIms4SZ8Y
ctRYcCgy/tOivnjYi1Z3sttlqr2/LyyR+sBORFEmyxJxCYgWmJjBjmB6L2l0
/OnoHVD2r7rPj4elN9ieaHK4LvVdRSAYpfABEXGv6QWUOydatfvJcLBFjnPL
QL9ds4p/2bj1sKEZH1n6bL9U34qSmqM6Hsx6bHs9z8fObL/C796n98jbxcs0
iSXugIm5W9lejtT8WLOzNM9HcJH5kOZDp1k0SjdVpo+5X/FYytYCq7D0cdxk
i8Y9NVLTX1cGOWXge/0AUOgIe6d18EPBh2cN2H17Y2X1ZB6ezL5SV1eBacAB
9LvUZRVIEYmR4HJpppgm6Io7zU046iVJxaKUGP7d/mtROoR6L5IqdC5FHGl5
TT3RR6y8MlbNaQY0Cyatcl2TLARuUkapfXxu25TUP7Y4DExUUFqe2E5jIxxL
Z925jueUbQQruju/YimokQm3WQokkf3T41Ys2RuF3WlqZuIOP37felIn4/+C
UILCGNAbf8VFAmMtXSfOraO3RfvhZ2G3kIw7hLjrdtIiInpfHkbhWvY1xRUh
/TRbOuiCsUuvQcDHpRIzxIfYNa6mmVjX8F/OgipHFvRZ2WhtVAr+ymouqW8n
pUCKHTdGsRs+Eggw75vKi2FlaBgjdwCIz2JHJk9mFJ1CwaKkc2V76V3JnWiL
mTMEwTgPUNyW5XBk9msoseHX1wQp/Q978oV9wyW8MOvpBhj60+7KsOG614uc
ikh8FWGUOxMlY4iZT7kqD60L2nnPSKjOPswKgKAQIV3d09vBc8MhTS4RiBhU
Vq6Ml9bfhUg9XguHGg6fvMvMLIzKpglG7gWPo+kTWJGOprRbO251o7fv3Omu
RZpRhj5k3BOkKX0OW+sqBrn/nV4MwPxWKYbtGhGfz7uRlUP5qe4koqJB5UYf
c4Vd7EpD5WXGhglCl8uqRybaV01xnoVJdBVZ7qrMFrT8VPQiHfXQAS24RHnr
5HdH3926T2XL07LWMjerbeceJDv2Jg0T+muve9XGgO78nXBv5IQIKoQs83Td
/byYQwOBCMoHXoLRSCe8s9a3vHGqEEbbXs09/+9VyhzCOCo5m415M72UE16W
FAuzUWtxbJHZfaESD5/aJitnk1eLGxBRHaPWmT2QrzvzCP+1re2+I3dM9QG4
Mcgjk8O4c1ob59BbU1Zb0OcmCoZE0Lk7fp1Yen7d4+Vxh5dkT2hItpWBL31+
TtTjt4u2X6PibzDHEeFHvyq8wHuSfZwE5TvTZfDSYv0vcy16SVQ1f3QCAp0Y
OIyTJEKmrl+MgkrRlwoTkk3p9CC7CeXO3Ftr3Yp0RSVvYnDO20xsjIqeOMSE
I2nr1IQono9mAz+LrNuGPjENgcxz8QHtYsCjj58ELaAwv7RVLUIPEhBvs2eN
QFUv3mwj7m29rzYR9wJ1kR/ySvRUtUxTLSf2arZtmjPS79nLsqbDVLRCJTZS
aPLv4dTppA0Yq0HBVgioPnP8SMlmbcQqIQQxLJCKPFR6WwPo3M6t4hMPkWAm
57xnjZtUdfk6fWSXcjwlf4XPr0EyZiXZ/+4V8hRBlL0G2WWjEk59/+g6IJZ6
g4s383d95JDdg4bDNo/oIroLXTN58jqQliH50NK7cENKjKGW9KAQQlg0X6d2
3BEm5jFriA/zTRP80fV2HH2DddqqPZNTm4ejghsUxxtPG4xl61OJiSE/AexW
LZlB1dGgneSk2VzqS+pKZCB/pAoKjy8hulhdU14Wbs/HTVNMSGH/XdJgerGM
OcqboXP0Gwd5B6DZ7jn/zg60zZ16I1i/XU7ZKF+QULJaH4WBHjIU68CeGULQ
Q09GUE/vZJzghXubW9TtfMtVTWXrZokKJhQT9ls/wPRf6ogb3R7YjqKB4OdS
I4MtLX8osZ4YeIpuVKL6ObFOzcsxsKs/M4zH/9Xw4xScxR2g/MKn/J9rYKyt
xQYsZwRTrTbiUimsRTdb35+2pwNFFAMvvzCw2hSiM+zuzG7cKsex4tG+QBHj
gwg5uWE5+qdI7slQDqxTIRMbUnBUvJ8wRFBc5CTuX41IOlemkdefcoPIxvdF
3nVieVhuElfftQHnJtrgUBI17YapuEkPzPGpt8j17Opx36E0pV1A4B3gQQ3y
MPizjdJ50alMrro+c45esDHxuoFW1eWwTvaYVKVXEULSCV1mg6ohZpLHkNnr
u2e19huP0nriUwBvtA4fhca7svyfPTquZbAAgPJ3SHTZ119vXYqhaO/Y7vA5
PR/h1yycA57eVTBXsJ+DwXnm78bGnw2zuUpdkgd2niVPAIdYeJV1kUEK6d9G
gVXf+Jfwt83qklw/OlQTf4dJVG3+WpPJPR7i+ypBSt/BgbvBQUC7wDW8cR/3
Cn12YE3jxUeVunKIJprmktxfLqHsosRFB0Hc0O5933JZ3KFIeOEaRvpq80uE
fygoZrRPXn9D/EnsIIopYDTL6kzQjZsIRKQs+KDKhZnJc4378NZt+/sxv3YO
YmYLNqgwk9ZH2OHrR9LZ9z/od9PgUsCKJBZ9D/zYzdsTObPSgxbu1bZ2JpIC
wuu8dg7Ko5vfCncPiFaqKz7rhS03cbaeC/1MynrOPBQpOhn0lpDTAuLu5zc5
CsyTwY1hLDAEa+B9OkboJ8ZqgrK6lVKMAfHngiuyTkXw8GgF0KA8NagSBkXR
HesrauQw8EhjJl44y3WSESv0iAT2v/SnM/yQX+WlJ3FyQ/alCyOCNsCTRuSl
AmZx18OSz3KANCG+Q6KoVPCmJyLU7MtRLnX1eCO6VLyFsf2YbYt8IZDaN8FP
1WQTnaAS32/PrV+R3ApYJVITbCqYP1bvdNVsPrty3IH6gGoD2xs/6AaIdBfW
bXoaPz57X26LrZmegwoxym5SUX/UiBiJuGEYg0OrxBHSJaYUF+cocCWi1OGt
6ZFkwJAp65ufEHb8ZQzmnY9B9H64SRXBDu8jNmUWtlEMfljmqe8FlKcOnYlp
R3PW0JQDLu95OYUw1Y9QvSewUn/ltAZpEO1uFybfNrf6oG9tkD1nnq8w640A
ZTFkGUViW7AhqYLUfB28GPDVngdoXVCgilVOULjscZp4ePjtgvV8HMFE2VvM
wjjOdciQ6k3Ek+VeO9EKScM6E9/ZYzMTjvI4QXEwUnL4buHcoSPj0V/6S9Ro
1DNwgPBUjQ/rOu/dAvuj/8AVk7L65r2KA0ykHRY6wAOQew0KLDYGSJu381ff
SYDpAUA+qPNJRHSPu4Nng3m/CjSjN1Xsrf5lVcMWXcfXOWDOLzwUyv4O3Vjd
Mq70rgON0SZKbiSQQD0whGwhMMMqn013/55MWC2JorhF9DNfXgrpf3rjZiG8
/rT62Ze7FiEVD8ro3CADWV8RapVR5to2oM0Gj7biBH4l0EQiVumfNx8YlYZv
E67kW890oWU3uOylzHnSQMH4Y3M4jfOXePZIv31m+cP72l0ReGPb0TuqTyV1
xeHtSFG1i+ZoQNZQF+QyNLzqmuv2Fl6XqXpQmTBeBt1J69PjA4YV2k5pJYRW
sYsVSpi7chABtqQzrMP1oL5y3J4ThomCj0T4SU+DZh65Pa9yyWIFlE4egDiH
87YgMco7VeI09HrYkDSJjLDLxkXBalzHQQ5qvx/JYNHIC/QLphZPBJX4Roch
brFaLgTReFB2bwAetKYEFXXnWkdZzKNmo8DJfi4i9EvBQRy1WGqqxjtgsVRf
9i7aVOz4Gf3OrFEu6EgncTn/5QcBieKB2TM/yOCOm9KLZgcfNwhKqh14xDsV
hxjyhWqk2YWkqUSO6BesO0ht0+XrwtBXUPOpgJjWUjP2i5+BMWceD977oPoA
g4QAPUPWdn7HHyuDZVlGyLR2I1TRylvjFzEy5NWSlKPhnnRNocGyoy6j9qp1
HI1J/SQDmr+m/rdqvMYVT9e8/89dYmvLFqGrAkhqk6i4EGz5/qCzBovbOkNs
fJvZ22V7iYxAgizyu9jsaeBTQx2e5CftsythyEnDDh6cSy1qZG7Frce4VreX
69meXiLpVKRJRpggv7R8vBACaYyN5857f9fTgrEPuKDECXAV3VkDVVwLRrgJ
0hdbJW8gAVW3umX6lNFT33Hj2AbC5d8qhWsq6d7J9XkTUFNDrQ84TU4M+QqD
b4De90Sm/tFiPUCSV3uOr/dSCuBOHtleZuQk35HnFmlXotD0yytLduqRSAUl
VZQU008Rj7ONUoIiuVTybXB85CxdXzPayVPS+TG7Wo1nLVDX0s4ALn+nVQIo
e8xCna8ykND8pmYno02iA0SNSP0yeaZTMQy/bOVrkppfT3yPMPqNfxd9WzXq
/uMmSJ5GyNEq4JaO+5tXgYJASwzU1+6VVc6cxqomlqnt7YpPNI9tgzMApDhq
3ndb6o/AAi1/IA/Pru7UB+0oPYk89+qIz3OPoVCHU/kOkW+NdAqb+wU1VHT2
7Sb8AQ0J6jMfyoDazCW4lBHz4q++AEDmS3ql7TwQVvNRv8KdnvQrVF/j8ZMe
fYS6b4UKzAD2EDuo4gAKX+6DlLRVsbSGp5HY6BNCUGFxLORckLLri+4+ty7a
EIowTjWxU9CyQBv/YzU/atbEQWoXQMQjcl8/v1UAIJ1Fytw2fcUNkYiN2zmU
LioXuvaQXumWl96amJ810CgvaC97Na51cQF2/GYr/1XKvpwpzqUZ+Y6s/b/8
zLs5aBJ3lxWxWIQsJR+dvW1/KoKTJxjUKSRRUj2FWXhcfN7UNVdUAbpDzXzc
t7s1VssEuaxaM7xr2V3gk/HwKpc1YcUVxvk8P5pwur4yOHVatCdHQh14GDwP
OIdJvKyrvwDPOefnO5d7AgM/+FGSS7s1shIPaecw1wTxJ2YEkiegGPk4d2b/
5aC963U17Etrtznj/7VXiPTD/Z4SPJCeTjoXKkzUQQ5bBHR7uYk9UEbJQEKR
kMGeV9fvlRS+ga2UT/tGsrCwVNTRSTdxviToXfvb2VeyBkQc8gF/oQCPLA8k
WXMOQo5V2+9mjyq+TK5X8I/zlFk5p2Co2JBybvd+V2JR19brwgXs0Ivfvt2B
SCcOGoTiMUjZmK20xUSlO3+9CopUTFC02GtuBsb6axqEkTekh0Bm4LMmx5L+
VdFSNOuOD/no/LWgIQON1xIEseoCPBVCbn+LX6MHt3S2isC+7iSkkZRk3678
HsXZ9bF60kdP4ugYJyUIwoCSgcetp+2DESO2PqGOekethV7RRvH10vFZSYiP
8xeUBSDjWoQs1VF29mV6LjRNLHYWcrpShBZbVTgLjO9CwJCQWN2/rV6KBLkD
OvdgSc9XrPX9T/OAgMs0rr0oKnmd3IXmwEYogm8vVO6fQSjjsWxhWAy2VOmc
UvsQ5ABlDjSfSapY79YL0RoR72EUQEtmp8gkmcFSLm4zujmfA9LpsrrXtVgt
XC7W8QLxE24BNUT9oIekYQ/jMUGIcH1KV1uqdXlzIeuJwbr5GVUPDiHW9hYb
K/PRR3lHv6Qi1AuFQK0jgFs3uknP5sbhludkTDdUoBVyHp4XgxP8G0FPXjS6
VsWXBBaj832bmRS2D6q3M7ED8d3scYi0P2V0aMt+Dpxry8DD1fktpaIEVVWX
wbAu9VeOZmfByxPkAEu6pyV32wMfpr2mK/H+ksXDb2apYa9n3OC3fFmsimTw
+NX4ZWMFfHlIeiHjuJf4AVeUMD9/g0wg8vmU3xejkx6ZGgWY0co0yk+XA2rr
ecV2O3dubj74lTAz/eDXISDSPoK8cFAipt9+g83NPiL6128LaGwaqZw9KgEd
So3s7YjPDUTPwGrpXPJiTTwPAumSojSVSCXeeAfpNClUX9edZN6NwuwadtFo
ZmxjIk8S9PtQEN3KTamZKb63ZgRFZKuIdoreCDWXVwASKWKltxI9lEQAq1a3
6jevU4vVYdVrj7UsH1jZMpdpuY+71BxbApdRe8Z0cxCTSMe5B0izqFZgg+Xr
nL1iWrblTFdnvQS68RnMI2q9WPpbM4rXE8D6mvzqg9qTu2+o55fQmZ8gYIKe
lToS3mbQ6D4JPqPhDwuvmkzFVgmtSNa2H3lDkNSbqsS+DRJ2NZ7pYcCMpv61
h3yisWryPRxP6SJgXFQUWFQrdNikc/TbNlYkXv2fAve5SRRPsXwo5XKCgvB8
urV+Ct1giXYPe4QBYJwdc1vgvhVYm0skJuKO2XS7aKN2j+ztqxoxXGX+F/kM
e3eQf2Ak5OcIm56qHD5Z2+8qF8MBhxu3GxAkWjrEgYJVjkdu3N5oHOA2U2g9
FCXmNegr5DOyfrfxWEnmJYrqE50oVfZU6lacAm2jxHSx6xrdTkvZOGIKOV7l
ghcyTXElOcsThHSvSNItK9eovOvkXWd9aSxW0Th4eni3UttaRgPbo4rjIklL
yblyxD58NmFA1woiOe3e+PZW1LtaFupj/V9DTW8OGhMntAY+q4PPMukq/xzp
MqgwKleXUHK6aVn5R9m6rWflQV0syldLPIvra0MmOdJ4AjG0AEGiRpglgCVq
1TlyjjJu84K9Ymx0hAPPAq1T5NtJaSn+7xkGza2m8fY3ecDOsW0mMMnfJwNG
pGnaAgzsHuVxGqvCrg+2FdqCyK52kURUk7L0nPDO2va9PpD3Sc0DnlcYrf8/
yLMJNiNYOwrkD9YDtYG8txuGCJClys1R5ps916LIIthDB2guL2wbvWmiHWq2
lzsL5maA0fbhbZv/UOpoBUsReu8ky7s+zGRigHDGK2wPBHrA3P8o/2oJEpHx
VVoGnxLBGxP7JBI48shs2FFvWdoK2gT/goC/ccBV8f9PdLCAuyvd7pQ7A4cg
Slkr2zQmIQXaR8Qf8jEfBg+71onn6M1UeLOMXyuYjkwSHiQJfxNXr3ffvkJL
JOkCcdSHmxCVjTQ5XbKviZ59thCuzTwII+JUqinFPjywiMpKVDif0kdfxfY4
H+j1Vr45LPO1/jp3pT3eapRqrni22r5nGP/bR1o4n6jsbecGAuOerTGHCAb1
5IcPyxeomBPu6RZFO5T0qQ1r2oEOVx5VjRBiZKl/IxWADhho3WLRBsJB45dA
ALAkgklVPDl0ay/HoFb5xUyxYuxvMyz59LAfdUOrCKJeBwZnlfE6UEpBh1AU
/e1IDzgoZvzF1YkRarjaf+A2k3BnAtDmWF+d9oERZTZDK8Y3Txn1Yt+rfErK
4XmNwrULLiSVGmD2ka81lQYDoj4+q7+S3mg9qKWlFGkAdDZftcdr7/bUrXb9
P3MvNA3ScdFXAisOdtRGzqXaLh1o9b8IRZnM9bfuTTQHrPlLyQJVdyPt+z4o
dmbtEwaplJJXQqGzFlIlWm2FR1yQkcz8o1EsWw3ff/o0T9MHdyYUYZtX9iO0
jVJ6xdQaoiRuxfArSMQE/OstzJv/9YSkFKr878bU3VZsLqPVYvyGvCaaxPSC
/11HKfa0fbBO21Vd1Ssaa5HvUbY4UJdSgJZakWf5b8IZwhJ4Yuw20AcXymZ4
UBN6GUmVOKcpOB9DhUyY80jgbyqWXrwD7mnqLargVGIhTaHZeOKzgNtIQ1qC
2/KFSLGHOsYMGO4ldUKn9fSnwFEW6KnkJVAj6/KXEXymrY0WnshPhNOm6Yor
ZSNtYCHlFGOecxoPTwR9H0AYA5SZZUSGj0BxdVgrOH5TnotgEl83gMrUkJQg
tcwYFlsYcd9qxGGPgysbU4NwKXW2qwhxBDUs4qAWN7T8fB4B1Y82A+UkXiMa
cR1h40G5NAOHmUuzVR7rH+MgMKzzPHTWR6783n1PwZ82fMlUIgTwsPOcCl9R
LvXkhKsH2OdUBLUNTPCNrK7Y2ivdksIiNAqqzn+3JiJR5jfT34z7qKO1i6Xx
gNuxrOAbENBcKq+sK0hY04unwcXN/jhHW3Xv6OEkanj8zuSJZI6mlT8zqMRP
/QUuxIYTzFW2/ciF+Kr/Gwv5RrsJXjt3AEWGuvuIRxgAQzf9ArEfemKH+D4C
nTIWa7bS5kJumj8ZN2aHBOh+a4Cj/PLq1a9QNn3bTWLl+945Pz6gpLh+Kvfs
Wsvo+378zkjZYvCN/4or0+Mb+k2VT6g53T3bdaWQ/RZ4aGZvkAnNyklPy/hl
kvFb5ECQdQUH155na88Ff7qmOR8h3aDOMoqi/t62SkTHbBFe4e2NY4YOqfdm
ajgb6AWRL9lWsLzAnv4eKnL3mqhFPzaENXIBo5BAPCZO1cCSoUKNGACcJv07
Jp3/zQ7Xw2RlIZl6M79GEvA63A4qt4O5Xn1k4D8PlgD2Ddjx3G2SaqBkgP4H
rYibtc9XEX5U+5I/iLCD5CN3nT4PnDB7uGIAherLFqdabU+4h4NmWgg/+ZQT
0ZDH2G1BJrKKBf0IxbZ/496WlwVzpjIPFRt+VI2tvXgWedruuj8GfyF5gZR4
0xQfqoLZM/2n3QGr620u8yw0vILcRuGGUz+wzTd1nsfXdI02UBEImhzTogK5
Ni9BBUpYwUdQIsy586Q4gTVidX7tpJAkVJv0ECW9L4vMq9lbcU4ZjknYb3b1
xUSNYwxK8PmTkK26WazRlxTV1uG80TJGkBMwVsPJNZY+zziCVlIuw3TkEZg7
hyhGiExlAQZdvy8i5Zy47vjulKTXRJAjZHFX6ZWM/C2SmJxB1q/ASnjoDThp
A/3NVe6nJaKD4nJqARTUe+qjcYDnREP1u1eoOVlm0dfeiQGDFGSpMAbp5hmg
57b+ZaTCJM6DpC7QNq6Gkaf+3ChUAH9MncEurrc+qjIdEakC8Y56jTWL467W
PB5buw+JyUd/jAUh6Jnl57061BatBkiiZVEKkgn3QYOdzzqVBP5vYcVkeKHp
56FxfIbM9NUBxOfcZUXr63Mri/zvT7RI/QeqNpy6BYhRcoWK2ma/q+SU1w+o
jvd7O8QDs8bCSO9injxJo9eUXfHCk+M+ehw0VsTletsdQzg85mWG5IkOflhq
Be/aDkdfV7ZqCQoRlXJTDJUtcgP3CRJC0oddyY/6G5j8sQ5RZE/saqJ03P1G
DqYD8ANhayOu2SnnPBPbqWLEhtIIkEXTzCh0Mxg4AbeLCspSbmvuOkX/oNPs
hqJaARSHUkCsi8Yp0eAmkpfuw2C+I2evr4TqCOTcsn9/NKWsdx+CBwXzU93x
ZuQ96C1jk9ifPYYRX95m/a9mabUT4X9jxzoy7wkvpm4uJg0xjP0vhJ71vNfF
8PXoid9+uPX1YZjTGxvExfnyUsJ17z19LlVCw+aHKlv/ATMh7oEQzn4mjOJE
ymGQ2L1T/d5ozpUH6/nJ1YAvCz0sIswRodw2oR34oZAjU0NgMuW6Txge48Bk
GMcZfA98IFqLikat5151oBkDdjasfFZIEC45qkLed/4PiXUtIlY+bfr/9+MQ
7+9dApSUdzdBS0BXNkdOBGjwSl2y39T9ZQUocDNuGwz+kZ2gVTwo4scko92Q
pyAc9UiFoCNoHy6/6yAx5S/FyuT0VCUmyRyioyfbCIOx2OmYk+8vV7n1FlyY
JCQacRwqcPhlLuGJBX2UD1Ughlc6r8OPi+jkjKgJu3bRHxlNZurWpdRMAqQJ
Hr/FsrcjzZ5wO2Ljue8/2OsDKPbhV6MJ+n7oqdKU0h2nCKv5ic++f1GOy/Kb
nettCyDs3IVKq1vkmij1gfCIkInUJZa1YIunTPBtH1wDxZ7rqJ4TfYgZc4rx
B9LUUjLY2BTlBmktFRvc3Wxl5qZQZ09T9hgboHz76Z/faYXp5WIQPuflWIqx
FH8ifQgJ0rqUpwrMa5Jpck34lsZOVHVgc76wiGc166tdygxxDleeq/yx0TCZ
FcPDRhnpc4CKeiBIa9RgWH1dr44U3zDepPFZhVNNgG8G6/j/e1SwD58La6EX
y3VRuIz72vs0vqYGt/1D5ShZaCL5oKKPf3e75ECTVoBIOHZ5dkZhVWjYLawl
cSsiVkx1RfdRXjXohdS/a8S5lOaCEZt2knenaKQfBhaT6+rU2inB4inWuAr/
MlE/qePr5mvJ0cKglE01pJ/DzQdQRvasrpHiQg2/wu+Vh7T+y+WCmc+SbTSK
W5lxrbtWCBGCCBNfxWB/bU0gMp60sEfm67NDrjCLstxRdrff97vRwaDHyg/4
d0CgsKNzA3EJ8q7ih9WBV8hHRKFETjz5jQ0h1F0fxPJwioGspNIJMvOuRLfS
zXNnt6+W7f2i7CDjsOuRKdpNW46mWZXgQkamQe4xKYYHHN3LGXAwS00Qb2aB
Zh1JTF6GKsvWC268oFrhEl5IDSm2CHXH0YkuP7imd9hHNavB7i14W2gZ4xOP
pqFmGRXprmK9tv8+7Q906usGTvPFfddRc/E9ZovQrxe/JBcNcQ24AnvF1MzT
XAko+x20qadT5BpoaxnLJS8PAOFYKNm+HnWdAk/2rhDu0aY0h0DXKhHAXu8p
tW2kIg+SHKdN1w/iA7zyuhsfuTDHhzSy2fI9cn/G6waJNNEIvpWqTy++m2L3
cwJ3F+EdvtbsbelQhmSpVZ186avlfmqplz9vq39im+O4ek+0swd+U+RdQTPD
7G7ESZBwem81TX2Iw4ORuRFJS6O5nWmYP3zXWlsoPAH5J4BTOSr/ooz9nQag
eMcgVRlrzfLBdEw6bbkaU89wBlLi72NjhCWaaUO1GUfZHkhAJl3w1rVzDd9W
+aULpxOqJtRhulAAApfTvlyQunPtF2U0tnYY9yjdr3o7o0rXtiuCWaQbpsqj
j0WK9dIF2ffbHMAY2drqzq3lTyWklfZnDNSgLtnVyrSRdIXwJpMN0GYwK2ML
CFfz0bH0RH5Mv19UYEdgDOBlJCJBUcC6VnhTqZdURekCUgGICtNjbeLu46f3
fJeNqACQ4WL5VTIbCf+jyPrCedPP4lRjE91vbKKeqg0tmFERX26DfWigbNQz
xbSg7mek/VLZ0+I5Y0C/QPX7lU18BY6caHDS1dm04TThlesuOFMwYI8gAtpJ
dS2uZu/X1HaSWTFV6x0uKva8IiG81eITvZdzGMUj9xM4hZS2fyrP8SUku/yc
Qpd3njWsOfQpztBaFVGkq9/J/WaRBD6Xu/vuPiAJ3t8Bu5wpALJkXU7IsGX4
iGg02B7bczCVBqxDQgfbXcWtnK3Z2GILlbf1vqSbRZ9OjCCkRnAZMtQClr7Y
96S5aWkt2NgADMd+gbbsIoIQzAepezNe6VY45YXw6rzfgE51J5a0YQfA51GQ
HHtSYaXgnAzCwKD9yw5aWIm/VuR2EjR2Yz+nL/jAdp8hbtttnj+cZy1U4kjy
5QiBCasuou9wOr5ceSO7ONDWoJcxtR/jBkQ0URzU6QeynGU8GGWjjdTk0fS9
PL1Szx9b437+HwqTBFBdz0GLR5UkymQ0y0N4rhp5jdPh/3c6tKN8P5ijmyJq
ADx6P4K+ZWaJMmm/CvQBz/i07JW20sBhutSqM4CRs3YxzGJ5FiwIQcwA7ZgC
T2HNBzprUyt1IsYtIzybNg2P5eCOwiu/D1jgW9OC15IIK+Ecv1es30X8+3oY
L2duLRmW0b3nN0xHtipQvbBNQmfAApsdP1jCBn+ull1sNyibj7Gaf3w11xWF
ZdY+v6fAraUS69mndO+zBROMao27jUEIiFshe9l3Ym1KK9Wr2feaDEwz1mDh
kFmphz0Ua/0P8/+NkKTiBFP7db6cdIPUKLRbO1R+1X1h6c17TDJ42Y+or4iG
wguLdxH+85DHdwZPa8PjTQ4Xm37MRgdOakOf67JDb+bOz5DmLIXr0XIAMqSz
b0XucuWvTWrdhhWY+mgVdbXYcMMfQIH9sMbqMkQ+nYcyEPUL6YSukikTaS7i
OdFahrwrUomeEfy3wpfBaopO2tokc5j8pgHhx2KHzE+t8Nsm/ySg7PPNFaAk
MyumHDO3fgG+OasbXbKxkG4jhgGj7MdjuSK9Q5JhezQ0jt29oqWi82vfgAaT
K8AyEZaDuk72KQldMxxJ7krJjatQIdBU5860Mg4a/Tajvct7Y4o7pC7wWgDH
EhamY5Jx9feeIqlqWg0LefxyV9aw1A60p4Sz+KarGio/XkItas7zS7akHDlU
g74+FJjYWWgZ20thA3sxVTfGxRK7BkrKx3dh+mh4A5AYl/IIl77U24y8JrgN
0Fg/2sc7XG5z9xJcryd25dlrxTG+L/tiYW66ZtWw1FdTWNj+ZDCwoSj6YMEF
Uh1XkFQN9YFpI8IMRliHwb1AFq2McLnexW3GKiqzbuFlD1hUNbmdqv8JNJky
FnPQttxn0IOW3FQ4zgleHEbyobZN/DHyQxlvX2NdHXd7ZejsA5GNei8ty+HA
oQNvfZnkWUrfy9pCfKxW4vJfFhLvm9+qZYfDXHZQDlORbj3F2ewOn2irSUaR
r8YswSCF5XjGyOoyxiNPjq43BRdhvNU4zLnpSP5Hgz8P6t7h0nzOxBmVWESK
077TJFyl256e0osAeRIB5TVb2vAiYiS19rJqTtPvd6/FWlW2M57ETh0y3OyU
/QPMRWkh4dgI/ERpaQEtFZ9/RwY682hbfFSE7bH5isRC7MLFixWeK1LmIL+R
e4rfzIOaVsdadZLb0WKodfQTSFZZJ67Ps6eUdj2K2dvDShZlsAHbYE+skPxb
Pgoxr8hdGtaGKBOIB0fJR9lLieGZ3aBZy6dTagF+j2EUHqKyFKvnsG283bLL
kQCCXrJIiuMDJ9zdAHYYIeY68SzGx9kYACRl1XmgyJdUpelewsbOQi4K0kpz
mBkDkLUPhzf0Wee8WNkdb9VxvX8GCabYPDAcL7yut4XVLdq27yJXmW7FjdX5
BZcJipePMGxQmGdYIOLTQsy+otLVb2nfSYNXK4bZTnyVMpyTAPSdODg+Q6u6
8bDkC1+QUDT8F4QZPTEn4F5GOWxrsNJrIr/h/POHabix9GWUxjTUPNZR8xVc
ECdHZCfFT0SMzvEXKoHcDyN+9W0InoTyqo8VDv928raLIUmS0ikvUV7SyCqC
Y2cTTwQFqxGj0jFsgeV6zyWMAwZTOECaFKs0Qwfl/O82IGxWXn+7MIxv7ZMc
yGqetBpgQUrlPnHixgX+7sM8FxPnHPFKSbDuCHD6r6yPkHtyZqPSVor2hujs
rVyrHiihZf0fCkUlGAaNeBamw4hpQJoyqlWpKPX4pOZyJk9WJJPomzFjTv/O
MkXpjRHvGGSbAk6VkoIbMg6oEnNJbX6eJSKJFbrJgT728eguj/niILteDFDV
lVFWABbJgDQyFy6gTRgU3eqKEcA0K41frBNnQ7S2OJ7igLRbG1o13Gg9JYJr
nUBi8VMGuG4zldm19uo5knxL6g7AaRwhPfXYoyulCkxswpDeM1paAz95XD1F
DJhHUc8FvzhDLpQzypUCZdgkPqjpf1nD2QMiat61SHFxqarBuOBCST5QRGpJ
PWVV4qfIvMTSzOjyNBVHDlcRSuVDbmpS6wc1k6AnJoSrHyVGa+qKfvQLBFhu
OZn4nKO0MdVqAapXUrihelm/r7sccapa4Yti2sR8eejm8lTiydtQxuPDDpgO
iZSX6Taf6s2kwFk8cpWXX1+aM0DFQOyXen4W0EKfRChFjkOXo+b7GFws1OxD
shGbwxd8OwfGWHxbcMx0/FMhgbF7QgSo9zaaX9I2YRSt35kvVlo15L4XIfWC
0SYDpCi5WmZicn7KMP9taDZRjekduWRO7QW4kXia37T3NWeq2HZ45EhnQs02
kVAq8rx6Nx1E4fKl85IBduC24g8gj+rcoPaKxnApJmV0qrfvJvX/26l3rGO/
7Ldj9Gz4ptvfGBBHuI3UyttjiUDKC9iwoeSGkfKEycgB+YE8PHuJwVlZ0r9p
8sS39j6vS1rEgQRor02037FVx9HMG+gclGM/d8yNTAnjmJrh/CecXIk2Zc5g
nqxDfslh81OXZsUaEmgxnREypnSftxzkm6YraK5LnNESrxeaU7udAxwBeHY5
4vwVZWOQCDx1t9/wPifpvYmBE0JCzIhtu8avzNxGaJ16CJRtlH7mtcqBwlGr
q1iR+W4iL6v3I3oxWCTZbDn0W3yBIiyGHUG5Z/r2Yle+35KYtoYDGfgQa8Ok
XBLIfxm7E5XcBhYCjXqrrezUhlFSCoyIlz3/CwjEg+NzDIjg6qYlXiXXzYa0
VZnU9x+sUFYlmUaqhXPnPRQ3bWgKxmFzv9rSMbvvBYa7hXf8pGzB0WvRu785
OPWq4Kmb6oYJoVvQ5qx0yWX7vxvqZ7QzeYFtl2Z7gLjzn1Pn0NuIL0gDXLvt
nzYvbqZMwLUzfyi579XkrF6GbRO8cfaHzdss4Tqgelm7AxVbTi5JI/yOXm+z
ZTYDmIJ0uq8wHATSZN6lz872sb6rfGxPjUxvdTF9ML9yUKC8V0gwmZZjYv6f
irnNnJZH08SUhlW/S6axgsSMikAab7ko3iCXE3D10OkEYPdiqWxzt/3dxxSl
y9M9vHMWLAMqMq9t0EhbI/T1/APgqZoSmBrUu5/6ZNdCsqE9jD+O201BWYtE
xiySJKbFcGpVjog/svJaZhBOWnTyG5N3ArtMEEJzG3vCDV1ZGD2O1sOirA94
ysjPCmiU/jk8By1XopegH0BY7YgleXeG0MYxz0Urllq7YOGeUaX36MTpCOIK
1LS2c7xz2g4T+HLvktXcs/Og5wrk4WK9jPnaSm3A01TWJSY4mRSRaCbVHmds
Sfx0leKgjAdWcxHmMKWkNTllZW5tbTL9Zo1V/xa39k6KS51RW290nnDswjs1
j6uff9/G2IrEznzv50ygS0rIK0Qpdn8ZtJu11RRUMpUO2jta+nn+uhrcmGSQ
ApQdbINw2amt+1XgR1kMtSEqm3EX/lVuryuzrz0bU+xOogd+HIGYT7ijO73D
ibBXSEvomJDZxRLem/VJ59iLbasjnaGyZbX8JIpNfNvivm4Kzp/94Eh/quoJ
8ulFVv4na9Sp4PqAvMoqxTXd+Yz2HBLYBeU8aPUP2meGQ5nnHauO3+pE4iJG
/M+6JgDxIPXgEdxeRpnPBcJuJeiDGR7TpvSuupvg/0IR2WPTG7e0DzTANmrb
dGLsxCkPeCCI54CvMenc1pb/0/EJv0bAYLrGAZT2IeDiZHkKroF/Xmgdjynx
MpG6pkFFUeb80aLr+5nDGqmxu4tw8kZoA6ceC0zCO0Joa+aLzFjHFF3XSukI
QnBuNldSzOWNUQGsqHc2gCk5NW9lslWRofcg47ijzw9r7OpUXMfw5V5zmvtN
hEgQye/ynR87Ok8s07h+sW2aBBRoWXO+poRjmB15V7ffNEko9m5JwqZDuYOs
XhLbw3VEuasFHoWv8/KdGuiolKqiAAc4DOP8N34HBf9uA1+Kk0HtT7rj8uUs
nR77bGIFLrxdv4nMZhAGGGCDmBo8J2PhgizcdEwyAYCnG/LOLOGM2NxfIgUH
m6KFnK2JJ3cFbenf1kNo46Bgw+51Puu1MTlSRJeaxLLCcp4D8JkE92fbKF67
cKo8KK33/VptV1Fvf8K306P6x8YFtWKJCD5IhslDGN0XzF9wFHAeThVgr7Bu
5+cYEQzHp8DfMN22xohzX4NDNWIBT2i2flbv+lFqdhIlxOkmWvG65LWnImwt
8ubrgIfV8Vb5v16Je88gAaynYlxpKbTEGtIeJ7PJ3601/5spcJzQ1cyBJIQp
imrdlUCs57vBkldd5NnwUDTFiSMD2oReUT/6dy82xGoXI2NO2D43AEsxY7ph
XiXfeJD24qBMk5ZR7ULIvdqZ+4SoZj3RpE48Qi/PKtTFstzXeu9jaDVJgcGT
e+maH5P+iEo77A3ZiM0ruF7mvF8/Z9Z6xHo53locRYSmjvIYQUzSimQ5Gsnp
2zg/XRpGfOy7DX4Bb+D/9QsL0LgL2XccNiUwsMBsXm00msIDAWyXiLtRRo0i
OaG9t8d8mYR+fxoDx9JfIDC7g5qmtk/ZH4w2zEwGtJPJvSl54acyxmnHNSDC
V4bi66/OPKg/1I8vS5D4/B2hFa8NvcI8Ro9NpzbEaRDKgzzDWVcRLSItlbz2
Dp6EMltHgc+r68nFsIdjioVPBSXAri/CUp5PJR8wzga1zgmW6IBFZ8IEukk8
SXzb1uzWdZoQly07FaUiKBiz4YEIpltNFtOuz1r00Y4C3LbFWTtsi3Nnf/Pn
Y6Pcbvuda0670rw2XIdUMBpTnmnuk6QVMOOgjSKVqVBkB7tOHJGE185TmYSQ
bWT1WfslIeS8AFmCaeS2nrcF8OWPJlT1DcH6++4OAcIWR5YWV25Pf/MLAAuT
7z6zsriQxte3l6iC49+W7S25fv6+xK00apm960OoIy//Fdby/HRoRH5uUtjw
0vlS2KLgr76PhS9R4toQa5KguOVVvQLRJpiHd0WX8nMzqBFs/N5ifXmg/gE7
FMDeUCOAoErtDcm+te4OhBAAym1pFwcgRID2vCKHZKZaSwzCMW4XfVXDnjy+
fbBlg9O7tcV+gnJjbpzUv6xym2F28klHTPajQ3eSfPv7YLrofdA0u5SiXHjX
ziTgb1fWFNa/noEK16FC3JkjwsnPnRJ8LCsOi8fg76xxW6nqGLjOvrGGbdb3
rrZYATCojU2/7WJAor2TtdNJ1x/p2zS+iNtJEUO1TSAGh2yZLeHYaWE5WvO/
VVzh17k7yM0CBgPXlUpxl1IYxIOCZL/ioU99wT0PF0qo47hjt8ZKJWsFT/e1
cN7RMw8sbmhWLEl+3+XVvY6kzXK4pCFQ9R0MkJf+UXNlhkl/2hCuQalBP5XO
lkFwtVpuI/8x1nmReRsab5dPmv/ogJWHmrO0i2v+8Ur8xhgm8jYh+7fOaLkO
b1psHSDvXofcbjiNqNOFYab4vZiq5S8MTpqgvHztLUOmXBWpilrq5nIhd8wv
zFh/6L2jLooZA3w9NBxLvJP1IGtsr7lg7G7L1v/7vnRvLlGFP44MH1Clyc+k
uukN0FFLceofuknhgHl79G8/exhshEVHIAj8WB3pa9pm2jTCosLrSEHJIez6
M2Hfcr/iwgheOQpbnS1cPWSCmrrvw3Az4+Sp84dXf7kevVjYc9D1AO5Kuj2T
ZQAuTq2kOfC5Pqq5ObcKa4YTzqIhccEeg58nEcKL6g8yzE2rVujjsNjx5dFk
uYsmc5jQLnhxHQ+wF32Euh6z4jsctesehCQQyfyV3RAbUhecuGOgCsANThJD
xnvEX2mQHao/J7JRlPRQo9Dz7nblKh7Gt98Kd/OuEISkam5SyHcMSd4ClpNn
z4I5zcUYAb+osk6sYBkqXS09YIWcglTqti2G0Ar7BX/AU0aNf6Y0hvdS9qXV
t2su7RKmFSQUBLYklkvAzv4IxEtEHaHLTBXXzy7PO1YwACYT1bLA21T9aKIR
zvPH9/JMJAd84hfCTDbp/0irOrHwetYQuNKK3rdZhwKNEJTXf2cDlxo1RuWt
uPdC76U0UVQXP25xFkAmXs7tujn56btMSnAwxfBFTrIALPV778Cn8QJQHmPC
DCan2xDLPzEUErxNu/SxYZ61lw5gVzYl/0xdyJfkOu0ErHVs6KG0/GOxcty2
BTw40D2gikr2J9rFl8zlgDoNkKmXJ3AvqWk7xmPvNLWGhFSyeUXNVX9bFduG
bPnYVB67jWOpE3HHEDzS7+Gjdf34LO6gQBMQ03gojhgnvIRlWy2meQ79TxiP
UQTBnQJ3KOIWkGk0DpC9yLRBGI54GW5DwxNAUB/IF+TNvsivEL8mKWL3hA6i
/G87UKYgw0wCYGTLFZknAdhamEguRhoaoMC7GIHTOSCwi/r4AbLFID/hn1+E
nBlm1R3ZRxFiu/fK/Q+wbvVECffAFZB9XMlh1BSMYWHQdQ1SkFaBOO9mrzFt
27fs6niMs64gMBQvCMRu1ye/VELOMCmVlCQixVD8qlJOeBUawMbxDzK+1Snd
OtDIahewc9HYuepXdkBwcSPjH+rfJZHTkmlHTk7ZpVyAx8TvEZHafSiE9Qw5
C84qE4gNgGRXZCIjwsBP4srwGUf7sVXwUQDgR6O9taqe88QZB+HY6QYw5tFL
iyjk+JKUwfFe+R0Wsc+z7jgNyGxdwh6g4aq55of+CYidH/rAmRRdKT6OTeYM
5pXTGD3hvoLO/8/G6mvr8YJvC8oWDjx5Ll2UjrKrVtyKRMCI1PX7cdvRBvPZ
Fu7QuzC4MTb0LSUcX8fvXYUkDbmrR5t5gMGfoA582PV8J5d7tQZsYl3kjlBe
ZYMg3/OTxe4fyrWuT7Lo3kJOu1c+hdCRyunowbSmYSFLhUEfeFAFD4jjpiSd
7QZnN9f6OKCd+DFUsueztmhor7rKLu3YBB6liYYR16ovgQUr7fyCf4csuwM2
Hv8noWMDQwhUehKhpYte+qFioPKzwKHn5FczIaaQPiDU4IeapY6fSutgto4Y
dVVjrP6IoPcw+Emh/VCsjsCitoZyXxEaS6S0zAAjrAS8tJcHwbuJND9+GHKg
Cdxw4OByWXW46D8YQomCgI+yJefSpE0J3egsinzvGB338BQFpE5+kRIPqfsj
WAs7WuEvzdGbU1s9ppfWz8A3kC+x6SPbqS0IDSkhmxZKlK/gvWYa27CVCX9I
f3OkAUhETpOgrf3Tmv+ULL7TR3D+LKezZaZgIhVU8M6S0vuOxTECH9NOtfdR
TjF9mwYKaXGdAo8ex7y25CsYSbU5vzDGdV3DKyyi8pumU4Kd6eaMcuZhjzAa
58gxPWlGwq1Hw15w9z+mPCTYgISMxNtdStNb00pvAUPcUmAAuCIPs2bcDXVq
BtesS53O3GJb6A16e4rjz4SFnBgK4CXj/ZRJ1P5rjOh9t7WleOITXOP+qpIb
r9yusOPETSrCL+uSi7vCvItff7aM24EW1DNkaN3PQyh3BKFIf1IK9dQCIgVO
1+tc+y8vHEZP+wmT2wM0xFekWnU99PA9jd5ytVA/jLjut1EcCQBmEmY9CmSC
OMY8JuQZSSHERxGuyeUG0uziaYwj5mun3h86cQHxjW3fUhcZoqUY1jPrV6Zx
HG95wnPoYeaFckzVLUhuaT429oe6FLK+sQtm46YCQofC1gftzfD+tYWpdX2v
73wXO0mVUtR9h1WgwmJwLLT6fyCmpHThMT133QcZeleKfB7fQu3yeUfe1Rnz
btLWUeV0+uf7Yn7hDeMFTO+hUQA8dqkeYEYH+GtcwJGpFNToX06CfiTJbp8q
ybvRHnkrFeOt59RU0Kp4vCWa1fW1lXWUyiF1IREfQPA52/0OokyWobXJGs9D
uCHRJ07wz8lvGbpJwexPAC8vDjknUghr/f/6qm41YAMFjy7gaIhRQM4mN2d5
QsIAn8xsXlqOtlOz899lRCWd7Q5fqLGCBYZcxzsinKwOAdnAoxEJWGG1+kAD
7ePslB6i7YZpjAQ10ocRYwJYQf2jkDnih8HTqVaufMH3XZ6v/2XWwKRQ4bGq
0YYYNKpA7owF5rVhsLRVA+pIh/8p83vvZRV2yvvgZuZUB9SDKYKuf8l1i0c5
QYJduX7kaEyb4V1ZUyudq6u4qw5b4+y9Evg+FHJImZIvGovE+XoJVDJs5H6Y
UVA1Sy8YvxNYxy7C/T/RJjcjF2gdT6gyKrEoEcPk1+A2zVo8/YEB9hNopDPb
sNash+UvDEMJV6cl8AVIzePYnqaitWOKifwbJLUKyDSBvYXj2t2czHBFSIvG
vGl4zmS6BVzqOHPYLoVOeR6eVliJ7Sbbh2Jdju3Ts9ZIZeW02/gbNhpG75s/
mqPBSpL+OcInFt9DruF5Kyk6Nqw0PVCV3YGhmao2VwTo7QedWWQ/ZMdKcdSS
ddiVZQEQNtPm8B1fkdzK0ug3N5a4XSJtauo0MqAjkd/0KxjBHx68ngGENIBZ
OBnjxWJ09sH4mjQPQll/9lXU+UyUUPVXV5YVwkAYnEVTS9rtvP7NlyfbmrMU
LyBbo1c0NieWzgD2uSgFuCh/MUKgrHrNs/7H24rQe6cMUN/83ktA3aG5ztbE
UpdFI93SL8QnRiedEKjX/+PtSl8vz26sXjBNbOUAgRowC/NXiqKbbvrg00S5
RoIWczcbzA1tNiLvh7fxmgYS00cHNkN4qcA9Pv5bMUoKet14lsD7mUNVCyR7
fOZBskZgcOeOhTDsNZ5l/bfs0otM3Xss6aZTlaTKbI910V53sAs3lJ9q600I
TAkUEJp4B8EzZuOb1cWVMBScfboZMdI9GvYxIn+mSAKWz/2o+nrKPRoB8X8A
sfefFeQBTh6/BXjgUdTMZoAaYieM68WGXylc0fNQL4mOZgHYk1Gh/vI7w5Ay
S3BOIXbnNYH9QLg4T09v5VjTfHCdsyniFg88aG/QtjH2bd/usUbiZygpDtls
oJNw0BNCP8wDmRyKxGowzaICzN7/nwMDt0wzpat+VDSInChx88MChsStWRsv
G3ubNtmBke8MCm8joKGLfitJRYjebvSlnxjxhrQGkY1dDYPYjPbQBD6TByMZ
dQnEGNVjqo/FIUZpCjw0V5Oayz0V6+xtJ+FlipZtYLFfObdJTxvsng3553GM
52r5p3zCmnQfCpU79RmapNN7f06auI2y4V+gkcIJPw1uZFfHvqoYHHjVY6+I
AGrEd0xip54qRQMiU5r/Z97M+ZNh9wrBwxVkbZUQCvUqGe3Pc+PFEU0sUUE2
41e/d1yTz/QGXefhMWbI2FKYSRalxQIfdByOOp+whS6a1BHdZPCIhqpyJ8LY
yVGeqePeEr0U+rpPxTArMtUyfGrjDu7Lvc4UNROzjbiuQ/Mcv3UhqwPOivB/
baCTJ7RXffqlNjC1rn6Z4cAcwygUV53JhhNWqUv8tFPOqw931oHqL0fZouR6
7C7wpFBt+5yx4P50lgZ6BKzjxNCR3vjqJ54GbVn0iZAPs9wILV7HEwzJwzdE
vvbgs4K5U9TECkRyik52u9DPhBqLzjs94GqW7sXz20993Ic0S/EG0/vqjpfG
CMKAaaoL/P9JjB7OAZM1Neb3h7n4l5zvmjPm+WY8tiOk2+F4sXSZiycydMT6
NbHwc6ZfYc3xA6ft3Bb9BcAGr4um54+uCPartvVb3Vf64d+urJ73iMIblqGT
A62CYrkrLEhbhCxTAijSGfVDzu5oImsQRQsGXf4X2dlv0ggg1xKYTxiYskIq
tV/3jq0SNWQGD6zDgxQgZJpPDZ6sDkPcp/U0bb8pkLC82B31ga5CcNbNIhcy
oC/lh16hde9ZFurs0HB8g7pnom47dCO8Zj7kosFv2v3KnD0M2YRWrgq4qNIQ
umuupo/6QzzRs38FWAHknvHzGLDCWy2hugufdaQY3Yv/SWg4AXJBY5vNSaBQ
uk8PCFtskCl12tFMuvSU3/dBhjX+IVp8V1kxhcRhLUGSJSFw5zIUVOA0DD6Y
DqQRvm5T4AWLfaUwJDykXkT8b47+pQI3cNlgbQEXT08hy7eG17ppcGMRsgeR
OQ9XhWt/H3DbZT0LSoIGpQqZ2Ml4D0wIya4NBqBiAUAGo2QJid8YJ+lchWFe
h2rAPoqGwL7iA69Mra3n9IltxLBZKTO1pY+IHNxIXbnJH9Eg4CoIo7Bxo3Wp
Ab5pukjkj9GTpKJcTGcRIP/w+ndaEDdUIBtZH2zpyw1X1GDlNP3HPDXR+WjD
84ta/scIvVKLii8Hzg2rovGi70y6whIAFhRps9mUe7uPgshEy4M2CfkPm67A
t9yxXthj3uaGaqNhAbHPbcc1RfkJ3i0JKoJNT/CxQooGwKiaJv5GXBcaW8DN
tUzxDL7weklP+0a5SKz6u5myTXMGDJ+fzGWt8XzK/YK2hqFY56FHecyNkCrG
y4DuSIUUSA75ovvdbSgDxfFG0Czh8hAGEf3f/TBmsMT5IRC9f/DmrjoF4nxe
O+TEbWbvREoARPBNUTD4vYQwDFdSM0ZIYwFFzZSBykQguIhttpjoYCvPYLfv
mJNqY19ynI3jSQoI74DpQ3UCLxDy7uUvecT/ezu6Gwn+tqYSL2+xULtx9YNW
2lL8bbMVaQUbwtXa0b48P62HoSx+joB/UGRIyYXW7Cqf7pe8Dp3Abol9OS1q
lvjKFds8C/ugkZRoMl9cKVXIOyUIRJZVvYVmmh0LxmL7YOZDwYN8F8xL5oV6
WEvOwY0O4pCeTO7JRm36gBcpCYNNb6VnYlH6/rWZsJlHk0ulXt4Pr+zLNtB8
IZQ7Jza/aUfoCxqcpZ3jPYTPjsVO7t2Kvq70L0ypswVyTr6bMi6HSskvUSMV
d5P/Ptmde1vILq6RBAFn36a0jtAg8U5LX0/WrLObrc0LH6eDq3Ysg508rHDX
WGCTjtVyP5KU4x3q/FkjsL+0UxDPKUsk8xUyNJ/oUexWnwvsF9f8VraCEH7H
1xKlJRbG92B+h7+BYaqk4F4uKExAYcVCxlApgTpb7slsFc8flswYqOdlr3aw
RnJ9PgoqG6XJhyIkKpYBCcCCbKX4NTCnNPOqEiLPV+m9q1QWlVov1y1tfbf/
F4xa1eF1WAebSbRtwSU/fSI4Ux5QjUEFKxrVR2PlLXc/a8Fwe4twHqJkm/BN
rB5MPYbERlykpEGAuPVRN+wE7zX+soAcgtuj3NBhLETNq3Nsfpy2v8C9rNAB
wCgT00YWRf3hK5QkArcjVSN4Foak93yQCtybpgo+lyAo9H5aK78zNcgyIX2n
kxGv7wAu/5CJAGd0z6WqqHu8kpUTvVHbDga+dm9mGx6trmcZ0SXSGalvMNME
P0PLMArZQB4x0ulV5OR97HYx3MNWRW7oDf3yuKPuZQe7wIdtnSbLzHYYbno9
K2xJLvkv8DthXlFJE3WrAaEXf1IP07W3/875vuXPAA6ZpyTitA/UfIjSsQMH
1VPwMPw4QWSisv8SCjXVKt/MiCS469pr3nKuU26ZlCZE15FIf3mGYJ7Y4LuI
OMecoxRfghLTJkoG/8NX4zItEdupD1fFnf6zUqEgHqkxIVb1oDcThWiMzi/l
8TW17ijqCrtMUL0F8bOSuNc4MHiasoVvP+vdD0JHs+zMFpz/fudIDghS7geD
y4khG+LyGjNoKOi9D3+Px1WJkpPiFLTwz1M5oelP/dH21vpNi9zM0zuMAFDM
lWIYVFcjTMyTOmyPU3wZnmdYyfMuZdBvcVlWbaB3OtdWkNniFYJslUqGKWfp
bU9EotTtk0ngcDlT3ZX7qtfM5G66cmuYqUMPwhBKqEmGuuaeLHQAbxvfHXR8
n76+CwunnocpTuS8Jx4zB6/hXVk+X49UhkPebeT42IIxBM06bIFFGnaadcbj
NZ8A3C8C6vcGAEanbpGQBpfUcyYorJ0AsnlNCCeHysp1xda6vyd4m0Ehkn3p
coh4PwFX0D2Rb1MrnBP75S7D577LW1amHDfmQsU8UkugBjXAAwUBajonVAVD
9PR4HhkLDwsdQpCpUFklccrM7vnftYTlQGMbX4mak1tLPlZ2/jPR29ThDtKD
F4gCN4y+gNx6YatWOUcLq/C7Fb2UmYcpjEIzq7+IRVC58vzHQbpxHhlR6//u
b0ubYRnPdZTlRZgb001IGLAlE4L8Om2SbrDckLFsAUcK/jgWd1HbpVQ4q2oK
Bq4msihldHquTHHkt/Ir5uDg1LzNYK6dIc4LZLJU5KzzBMcRXfdMgXN6y1JE
nSdcXEIZS7e83pg3X2nAAGr2Xl+VMEoTVmzS5Pgqz86XCzOtQL6arNTicz9/
Yd3eRAQxV0DrDZ3MAPm3adDTDb448Du4AUNSso7A3hmd+6HmspRJD+CeKec8
2DM09Rl15SQP2SUnjSoJkYHGEVx6NVASTDCKypiVnJb6+M444Ahtdy3CrerR
ccEdo/1R1tY55n5mYsi1G6ATOhCW1+2kqjQHy14txrho8zAfEmxqAqTu0R3M
bAzQBewQ2HuTnHHHsoLW8jE0wSlvDA5qtVBAii+UX10mGqxFbbIQzovSqCNu
3VCBpdYFpElOKYKftg48hoA1iWd1fCJPGqX/Ln9iKaPvFZpUzmRbJYw0/uKz
BJLyEtbSzERV3E4XTaJ9QsGsNgCVXkGyzvmADQzOkvSGF7hNRF8JA6tVontH
STAxNa+4KOrbELkw0wIqCz5nMOQglBBgYvoYUaMTyTueArbwCaT0vKkXg0p1
bRoHutq44zWfqBbz/HwdCCZuE1J7UIpPczgEnwACIthzgHXB40NQOPuFl+2G
nsAGMMzyrpBiN8isOhCY+62SG1Lrj8QOO8ZN3sS/QnjRQA4PDPgj8GjfoYsf
kOOeEJWkTV4oVXUbj7NomhVdikcLDlWn3x865bkpdQrilz56sz+zU/ncwOgx
mGaVXe7N1fqIxQco46Kc5tq2YK3QT5x/nFFEluLSAOt0DWK+5vMM24IiAQ49
ryuZ+YgOrsYab4iF7hPNt0GouVG1sC/OCq4FSmwvjyEPfac4trxgBeKJzLKj
cwQ4aVnioqXKcByjnYnALpvXdBG1tTLCoArVIpzmv31Z5pEVlSq9KNk/4i6Z
xvmuR2GNNc24UX/2bAU7PvUv2kaiZvX7LpwUkFTWXMw2oKn9QNSyLPZJuRfc
MeqiKXEMF+h4CG4lNcZIf33ymu21a1mPeXtUtkvM/LX/YVWMgBGjLeCi/mKq
T0XJ866MHhy1UlvMXqiygUm2qUmrIo6VsNYgAXYeTwxH2wHqInMytG50qa0r
1EMafMTc8RI9X7nb9AEBeh/VsbuY3Jx9FWhd1PnShZbBiw2dnZNs7qOfv2d4
GT1UTk9shfDjAYWZQjok6sxhdtCsHJWQ51O/kLJhsmbETqdMWxTkV5GTfQ89
XaYXq4+h1eMai/wSSLDDPmssojChGpACKs6QMO045zQbuxuvQEG2xhIZ0cHB
3GssrzJhCdijhI6QdLfuAbNLV4UDjeZLar0QSgdxNOgIToOv+lH/jw838ksf
cgaS+b7E6e+9kMZDKWP9R9ms+cg5NYC4fVz+dV+eEJuJWblxbuIdaGuMTp3B
YmpQC4fM/x3tXSu65AwYUozCpr/PQIWhzhY8B3TbB3CbTjLs8QHwEnGDbO2L
LZb53iqSrF6hHQrk/hoU8dcs2cBLjky1CT4PwMUc6TK9CLCy2aZY/KFk/ZTN
lt8jNGMLW4JqihRV/UVZuh0DU4T0iS1GIP/nb3uvkOkU8IFV/k9wgeputRKH
EdMS4WbKJ65r3DWTehK6+1six4qIb6xR8mZYakKMhz4VOey5GuNuCplk1Wjd
CPnO46Hn98AZ4ZcspeALDN/FtRf9HhoDp9Pvj3J/J9PPhZPf0rYqfAR1qSpC
sJahC8FRE8DVeA90Ojo3En/SnuGf45aAGlP6SV67PevaUNroonzuo7oUmfzz
5+fx0yqIPmRMu3+nnLVVLD+Eheb0doMzASE3YnGi/rG01PY1r/3jfk4B8V6o
DfGiHQYdrm57oQpKkjbRtAScPWNf2BgO0IEBi/9G6BiAQJC1mLggcpar3VA+
2TvAkH6MYJdWWwzePlrmPcXgEGdejzJzJC0i7g931X5BEB83Bjm0/dFOv16K
jBb7s8VGBeY+hlc81SDK6ik1wcTJFOLFwPflxX1miPZWYFpuy2oj2uqI4lWQ
bFXffJZ0ZnskzfwXOtAOR/lymYE8CW848zJR7ge67jjT4v/SuGr+H2kWdqJS
udAxZnS9MXr7ttUehPC/HfVrcizRQtqtbBIeW0ayicBeHh1TTiDqpXhRpA+t
WK/vD8ErVPXi14UqmmmbtLjHLmeGeSms/ViiiHizqDg+b31VQtaEQGq6cRb7
+B2TXDb1SCpvBWQlD7FhvGoYtLByveQYIpN0S1D1sMJxHwxWw+pMCUmkL9rt
QZTurOwHFmZixnlBemdPmo4jMb8I8fFev43xhj3+NIAkabp/xkQsye2Hn/DA
HwY2on7h57kygFd+n15C9ovx379ELyd2DEfvs8Q4Jo9JajJIGLVUYhZnBvVl
hQWtw2wXSroG5PjR8y1xDsZnNmWaXR2DMIjusqaa/D1Say9KwA7cn1VnyKII
0WmfPW1SxyWpMACI+rU7HyyswWlMh+5v9XbmRqRleNHlYCRSvMnoTgiu2eyZ
PvfSDj0OodSvWMGkdXCNSU6HWc56bngTmKU4dK89//LbYc6c38pp7FNUq5oA
SJMGk+yWpZ3IxtY0e01YUj6b8JMsiLBOFxW1gRqLFVT7YdIZXVR9WQsOLLbz
s8+3mxIwGoFfHMH81D5UL9a5llWLDbPW61loDEucTDEwdbyknXMCr0yJ7Eyf
DbP6QGJDqZKoEgMFQrOLnvk7+j4OUHk440AdAwSLE8AYHsrS0zeS0PPRE7+G
fXEDInQxi8YQC4p2fQAmI0KA7wWs/tOP4/PPR0fRrsewsA02B6c22/wi7NkQ
fRpYThShSiGMmZSFRfA2G31WM8zzXtlZx7e7gaV+fE7Fd3rqNy6bPXjEnS1w
N78+42Mz3SMy0hz2CKO1pdTR6LoHVPxeHBTJkztltKAEYIH20eo5FzWT0z1+
1cAJoTDguiJuT1YzAKFyFOENqBE0pIOxy5mabu/j26d/ifdnGScpA6SWf23o
ma40zje0wBCXYisB32tlvw46xdNB5lGNYGaxHlLjmt431e7QfnMcr5kZCTSb
tUgeQ3B+wB4QXrOpruzJGiXNetRrlw0L7/Tz2t0zUK+hO5rEAjTQHsqMkEOF
A7L12/Y9ajGMFstiKbvOVX7aDXYMIfLbMVTHOC/UZCKchAGSJj6+0HAMoa3K
cLJnzm/iOBaXoMcDFFwdJ7tKiaaRTFJRBxhVTZ7d8bjRiMnnCIH2pFlVqHRe
wc/79PlCWLoSavqeZjgBhJCpzT1pJV4rrmr7SXyfKkZnVDe+a7YsIwQWntXd
/Pu0iB/E8wv8p6nJVguQvL/ndiFwSIHOm6gGkpk0d/g1rOONsBolg3qRC7GD
cvdMaa1Cgyy7yO2Jcpy2GKyxYwlgUZJe9YEruvs3sFi/7ZVnTP6U+u4koO6T
uiwtCu91Ei1lEwMFwA0WmafIy7EFaXnVadzWPDC7v3q6as4CafJB8FOMN9BX
ELBkz9O1u9+kNc9vCwAlnAJyxH7tBS5PO84c+qCLDhgW7K+fsbIYSJ/JPSTy
2bEiAADg6DnflzygAdKbykfR/IapKSLY7jkRFfMIg8JbjXJMn7FGoEWwV2QH
ttu+RxcJnnesy4iP1hfU0th9qqUntoZMvwHt2uOL6AtdTROkyCS0fxHPjnj0
pSKnnWVk9jE8l3EQ+k0guXfYPBybUPCPkV+vlIRrEjay7Cmi+B60X1I/nzlE
CaLMx8re/pSaRvDcmHfWzExsi9T3rl45LeaTfu/lz0fnw5NWHJEFckkQtdvK
wkt4SYi0lgcRN2So+FLNGJy6qFsK2AmvDT3nmuqqVru9JfaQbvayHReLI+0n
NPHuPG+IwGEN1fVfT+WN5fs+dHmnQG0743E7hPBznSu0bapqJO6IMsQ79pck
kRjfn9/kaH0mM8h6jGvknJ9SFMSvc6yRpw4aQ3hGqcAPw+KLLj3sevJLybBZ
+5y3RkzsKjbm2fuqN5zOJ7qacz3/MTjGzr7V/j6vyBSEwUT309og0Z4Iw6Bq
9fzblMZhZaheUTyv2fGjQXb6KdPLURVAsjlUPbVmupLtbOT/w4mwE+aY3qOX
ZmncmndWKQWAAuPmVa+hXHMN0GIP21yzw1jy0Vhdd0J1ZxDKGdt27Tw6siEr
mI72BcONToAx3X1AXSFxF4leeLUYyU8l2jUKOM6DFjteWF+wmiLJVpDcBlp6
4xK5zB+mFF+w091SbcPOh1jFeJPFIuDmwiU4syX5VBOPqHwTpiyG+8zU9xKW
Jz+YKnMyLz6/kOWh4CBlUx6zWBk1Mrf2wRnLYL0GCutd51bCGc7vBK1jhGy/
0dl7huq/vOmN54ea1pPhNWBoF7aR8uplwcKvjUPjbRV3ke8ls4muAJcUpODa
3UxqohSHndXmg/LOAtSPa9qD4sMh/t/UOIUlEQeL9WxPVCYdo1C8y8CVccpz
xdGaRLSVx8SCuY+cGqITB8eAoJYxz8YktRM0Nya9Nwe9nYfTo5nsv1MBLDoB
Se57oTUogwnT/tzPa2VCaHU58Q4rRh86RoZKva/0u8zEnuFC3h4TXs9RyOIF
zQkm4MccONp29FQEJR/LfidlfIobAVCyeBeZbSvgvRp3+286/2+u3vfodLX4
OOEhs+X5e3xvWaf2UZliwQqzFSmxlGMnXNh1aRVIrx/acHsrKl2ptebBbVc6
hdyFO8ic2F2v82pcEQ9WFgAKMfLVHsGWnzo58EUAMQKN9X9zAADC2hsQiF/Q
WQFyADfrMK2pyq/Ba6WBsUWJE1P7a1cSRlrA5+qOz/X9MW+tHK+rJKRriCk2
OVRWDB01L+7MTr9veUzzArX+Hvl33m+sE8L5JHqBG1K/3JRHYS5A+/pM4DfV
h50/LKiRmTstePM15ocDQi6rm/+7/+IcyJjuXifpWbmt5E2+gwH8ShChYpfg
0xwZaLEYpCQ20HLpQQEBrGKBtBwCexvemfAbbwmfjpgaebKm7kWBnAYsjtSJ
00uiRVw31rZXIOrkj88MEojD+tdgc9LrQt6QigPEwuwCaqw5GujXT1JudSYk
rOdzDU8UtrqA9ejK7sh8q9PliUAQe96weNoQoOTcOUacPd/1KDNtU3HiN5Ic
1C5OEkJozLlbsS3aFKB7KVc3HBEvrikXaPiVQkNhHdoTtXxmKb91biqMVjVR
9OHA3C/LDM2p2Yb00cNyXGn1vRP/FVsgeXVcqjPgwAyzdLcembs2ZBFSAXQI
Xu+J/eYmbi8R5cwrFqBHrZMbF3cmsasw91fOYMZ5qsTn0spr7RGyQ4016Dva
Fr+pObJ393MlPcJbYq8NTyLXo3cnZ4D9BIXNCdNHax9SHonSGDuwoznZdsD+
7hm4+TIXF5idxt8S8/jTDL9w6goZXVMPreMRfjJbwTHRpIOSrHC+52JEoXA8
OTtF/HXFpBCzJS7iMnp+LVudKHlKgK5PeVsSIqIHZRVPvE3ztPuEZeWB38es
N6T3nm/FQiHgkFSjEA8lQMC4CMuPNsz4/uvL015WZfzFnVRttXK33MPRrxR9
w0JrzyYqFIWt1yhfp3MsD0rufcE0pGliEhN/4JShEgbjvsQBr2JFu3HOKJsw
deHP+WPnFE61477Xj+epx7gX9Rv8vZfmw3Sg6ngh8NfENjJXkHkVw3ckOvOj
MNExWfiIOpNG5Go4TgM/8md/w8Guq2RMxt3ybZQjS7SSYv9SD2gWzJS22aZG
m/ZLbh6Gp8a+jSFpoRx3OerQ2NFtuZmSqQTkKEEIAdm5r/ChHy5afRQ8pVpq
Mz1dZL/dzvk22x4t7DJjb3pIG2gMaFuSRKQc1i+01d7caXlEUH1pH+muIILk
tkB3CgHRgL803TuOG+SW3fdY9xHRFAzNpuzkNNX/TGDZL27sUY7kT+7aLLFo
VE+vgPoMri3JwSv5LyHCSIDzB2alcdCuzYoYnksWexbAaXlgRZgsamuWjkkC
WLBDPSl8J3LubISb9L0LfB4IaTwMdyDyqeSQ7WwcjUwjDs1+M5Qcr5u07ik0
72G5O+TFNp7j5//UiOHr3mcn60b4qv4qsDm4Kuf0TG5fd/rznSPeRr73FyhN
hJXHuGYf33xCBlv1ry8VmM/eANbnHRh0HCH7Sk7I+6CA3HkLe3Nk7zi6S/qO
/N806ci4GWM0IWRZDqq1ZHQ1ALi9ippOeFsfMbHUikN8lqk0peZLlSKQNaRg
2h05Ydl5PJMv1aq8S1sSUarGG3Rr34HERo4DlrgpztM8vFemC8+epnL6Miuv
8omYYoHKqtmOEfehPAFveXqgLrSzzg0EdFjW046Zuet/Hp1AaBti2wkFYMg0
7eNaotBhAiIuP+Bu+YdA8Pomgk0UbhAGjFWydWWcUrAh1h0guL48eaxnqwMY
h8lYAZsKvLQWM6cANksm53QY2IGDy2Y6SuNB8slsb3cviXo7CMvV5ylE8fqL
MQjNYescuLb768wRYqAW5+rBaiu1ppGtDahYD823fSGaTwh2Yke9tyy3wAAK
saNji7OzmtQwvYwkEGyI1I6xjAcMdB8xrgflKhk4QDH8fIH3MiJo54EBUaK3
UOulFv0jvrlP1mcOb/Hxp9znjH/7F0D2q98J1J2H4lMEsRnDnPxL2Hw+c8LX
1TI+TaomB9TzN+IPGYgnmeH6PMQHUuLdB5GUS1ztOswRTYJUV/IBbBgH3i//
nyVGd8fq0yd0zpQy2++Q3FO9yQR6MMRckeXbAgBtyfO5TPpEQ/paoa/06dLC
A1iwAFUq3NqblOeKdA+NUobxtdsBz/Bb13HDZS28bTsGQieskp4z96vuFng4
5BCQ1aJdja9IWeXDZCzN62eBRLn6pl6oJAOaXjxXhyD2Lg5fqyw0cGQ3uLhS
w0iAiw4Ys4WQst8iE0yk6vowImN5fYNUFZ0ICoGeG7VYzAmhAfsVnpnppkZE
XN5wTrwt7bTQ/o1SKBqFcFRffiZuTxISRzh/XwiNOTEyyzyLe36tKCsJaB3w
PsHa07CgJLvZwuvgBgXzxZLKauAOq8EwOJ0RuS6zmysYKypsPV2/CSSsVX9m
8lacRbRdCK/AXbXuXYjDPa3anHxVpDbsFHgrUWwAzGxGJpod0iMlNmMNuBn+
kkwxs7Wj2CkkhWOxlNWBHojFw/WQcJgnNbI4IywbujB1U6UtJAgs0EzfLlUu
oJiwZjk2YagJwHAGi1KP9miTzhfxDa8dPmlkCEs12T5UTPMjbzC6sCY5X3Wo
jC6wyJl4aMHglxrziG1SHFN32/p3nZj75rqVTRMqKslZ+KpnH2H6WeGFYZHK
/bz0CYOjM6tbfoi7d9gAetNrVOIHTzPq6OMuX0TZwLpasbFUQD7zn6M+kks9
mKSWucisgH4D8mTmS4Q6iR8iBh984mvmnUoTguLJ46mOzcVTkF+w8HPA2hn9
ktEoogdiqBNKLOy7JPqLwlHiLVOwYoOTSUaHUqfszJ3CNlsOdX1NROgWdhb6
X5ABAL0dgaQCihUF62+SmAlHJC+NLNWNVV7nGNBLKddhD5OTw7EC1DpvIIjy
OK4sXwgr+WujS+Xmvn3yJBU8jDtYiETQfFXlU3xTljovvxrIab+h7D+w0Ulm
n25NsSdN/LHe2bI3TOCrmT22vDnm4W+v5wx2kpczj680kqpkClQS/79Ob/zL
kiDHsd6/RiNQmiu7bH5ASqVyIT6+DQ/hRoDtaEYFmMg/eNs8pH68RN/pzdy2
0EcPps2VWB1Xrb+mfxYMbI0KJuG6NhFUp/7TXCwTEEMGArhQSFEHlv2iIL6Q
pm+q9BiVRFl9dNgpETUwLh44lQ3W/LyeQ6IY2GZyPVHlI3F6Do+9DLYJzfFo
QQq7A43sIpKjhMzbI/0e0T1GDQU5KKz5o2eyuh0R3gMhkyj1+ZTty7EqxiWb
SiuWbGzQse7bzOWXLNE3E/vzD+FdPvB2hnTuTGu8oqhbQrjL7nu8ApYRQ4hY
kP/NtI5zzRffzu26FMS2tNYhZNMS1taO9z1VLxFTPw/OBT1hpiMF2o85w0wE
+S2LZ3eQjnbALOy8hsrQYesfRFruLeTjS73rdIFFuiebqHzNeRdHQ+QpJjF4
wZmlMWCUV2rvapDJ6dDQquSBQQ5vAKL1be8kCcIJt0isAMn/6J90tU7G4S25
TZgh5yPEBrTjgoG/7VZ/xXmImTVNg61qNf9KcT5ygdLR49R2IlRQYLNvYD9k
HcD+qO+R2o8wuW606AAXdkZl9YSEX6MdYmZ89jhdzTdvAshjClBxYg0GTyro
eolJ46RvUUjJNzRo02kdYrotF6BpgAvvdiD2fCj/0ETnHGoHBRW8atqbZ/a6
Gko1VA+gHEOkzrSV53jPG474bGIPV0I8bpftbwBURFdOvDIwezbeiNPKwvKe
H4LuEqdtFJ/I0YG4JZgxF8Vmtx4IJcdqjKskWcRDhdXJ1ak6OBb2l8JugEjF
IMiFBvkzzOP5/nJgLTuQbqZxaMESeNc6a3iUSqUnXNMp9DupBVrB0VsGUGYp
WHctafqJkdcToVJ0NK7UoBRRXPLl5NlwwJ+AJPPMlQ+BchpXKDGJA72dQST9
6DoOi0ico++iAr2cueidzHE8zHV7N6DkpEAR6b2g04HtR89CH0p40pD/E6aZ
91nDM1ddkPWBLifzoQdtD66OS3WLWLzRoxObPKQupiqL50YoHtY330Mh5+Pb
FkrW2+S2VXd6yDGR3WK8ml6uB8n1X4qEYS7ZYJNopVrMKa8iVwcdz0KirL+h
v/l+ZYOqIsFz+TyT6B+LTZrDWCQOPjKZrfDOrx4Vev9xiP+YEHFzpOXhUf+1
Sh3pY30em2cGpsclyBi3EF0zp6O+UsOR4xp2G/n1mAvH0eQxiARwm/iiLZda
W95W8yVz+nLisCac7TTR1l4a3SUu+yzTQkSmJ5vkAj5u6SNt3xQfE09gmTJZ
ulSJBlH4+pZE1z8qaJccGfmtKZaPuAlxDCz9vafn7KutGAHAEGDiZVkQluWt
1rPZjAeHOYRyqGak5EgqiTEYHGh7XWbC1BnlA3MWHluVo3XbWMGGNRQ+EVwZ
/YvBH2thxjprRAjBLztSreoTWOd+Ou0PDWrrQVYYK33p1IN/cE47DOqJzeij
mv3WGr+7f5/U+Edv6j/DPxTKzfzLDvL1jhBUb1SOPAKBmkH3imT+X6ZZzaot
E0+Xc5EmGjGz4kaladKwcY/CUP1aGo6801hHyGAgZVbmh0pOZLCyZQAcbBdX
CHJzPyMAXKuCYGIHrn8m6FNlSrh0E5TLkifUf8UO/lVwavmzouT5l56YCMK4
Qq276+fu8cQ5xF9LMw8VV0HP+fgqUlgRbdbk2YOhDVrngRPaGGEKB3HQfv9F
f5jDd2mgHiF6/2ZXKIqDZh7lt2oPqzWWe18aprY1pGBx0TWun78dPKC6I00s
KaBlAuo+gymS5Ie5NIOOd3/l70xHFBE1KHX0ekMynx3jjj/kV5J7Cs7PmrSk
iVT31QacGviHWNg575eS0lwOnu9pVbn6zOhADAyd6pQKDMboI4dDcdeJYx3h
lWL5FWJDKG7vmPSwy0NiqYrdujfM61X65gIwErrF9JXBabZE1GFCHyK+MXiK
GGkXT1DEpIPz/xU9el+PKyTYyRCwz9ZV1gr3frQEqO1Sv/Uwky29ixu51roK
OYLzPhRgEU/VG0cuXLd4GGMU0vRK9fyp4g8bMuSHC5qW61RQLG3YlvndwQ31
Y36+OmkW+9HMqdhn/iK616v7o1Ax7Dsn9uXrNcNUijGq+u1M9K6MmcY3KMh0
OALEzn9BwEHdFep293pQUfTpX+XuwIJTqhsm1RBHnP/ZZ9NJ8mr3oy5FKkyJ
Xq84chBCbhKbbwHA2+/c1dVF+vXx4djArQz1cQWUqd1L1Tw0a2gIWiefXAr/
uZEE3KtaRXsu/pWnSDs8yrdZKzso1bpyUhf4yszQeAPuuLXt+SghYTBSx4UC
Nc3tolhSmONnyGii8W/yFdtDqmfdxLf/CarRYPdmhg1q1GHUacY7ZJabMANc
rjENwGJJzpstmyGaXHWZyAoawX6Jx0WrFYX+bZIm0tc/PusFqSBt4mcqqRnb
2iM4TdeGuFtvl8JYd/3MkO5SyoTr9ScOOA9xgB3JFBEmTAUx8/SIsN2n5v0S
fzRAp0IAKXVe721STex0Ejg1xEZoQTnuQWSvm6rEhWMy+WT8F0zt69HbWWUM
jCBwx4EoDguebXvdLZCa5ej/EcTP6ExgbG4yMeJXO19JWwVb3CUraAX1oeMJ
bRTlF3ppDntHLGZk+xRWL2ZkEIasN2D/U+FanVaHAPzBvMp1L2BEb1H7TtfX
d8lReBz3H3fYd6miM0/ItUVVwGqHq0MUuOZQCSZ+QcWufdP1IVvizJv9thXL
RuhAvhfTgJbTgJAJT/mKVidtOC7Fr28xzN3WSYScAfQ/HMYe5iuabvpjsru8
MFSCBxDto9XcQwC8Huapatld+UnMrl59tOj2KbkJ56pP8I7nTdkgbn3cQJ8Z
gNY1SJBpo99D1YL9XtqRmyMfinfkbb2C86Pua2Sj0dPR5JIKffpsgN8zdL1h
RnAuK7j0S8zRqA/CBCZmDan5U8z5/F9yxg4kL4Q87V7UcZX3daCpYt0W83JD
N7/M8V26hCRL/OQjeAljzIL3MIu4QXc1N9saD+NwTunKrIPhdZtQ/8BfPUOf
pXBlyOXWX5CTCIfazteLkd40zHrq0iM+lnF+FJl8h+lH+UMmmNWLqBZaMWbb
6tHWyx2vqDvtNbj0uyhZ+XW/by4K4HTyDWCItvMKpZi4y2HHE28SawwuSTdq
U+FZSEjzLsJ3hePXNvAEqiDTwTg6IPXSJf0IZA7j6BjFKEM1e3Lm7diOwC8b
JFYgeQKJhwQ9pgjWdqTxQ1mdOUVerAbd0E9sAznp0XlIliV6tybc5P9Ry5E4
n2z+J3Eujav5trl/9X3KqOVcXCCslctJ09WUXj/CgI00GOKfkaMtcTbo+TiE
PDuLNUu+jcFk+ZwioDg6t8022yLAoRAPlLAXwWZBxX8vOKc6zQjCv94/gZcX
SLIbSE3aj070S8Lsmy65ASbH4kYPEw+36KT9NX/Ak4sz1xpREPPKpRVJwvUn
lomfsF0PnZk7qDMFd8itZ+pC5jmdJV26kEVsFxLq7sgZzVCmohJYEZPtm6IM
yNEyTygkvyY7HI/WKQWIb3mLouJgMk3PZJ69M2EBQ0IkX98/7NMx1sQznV6W
NQS7TAyl9mawfumItLt596SBXFSCmAQEC4o3SJvtFS/mZ7tP+ClpalEn8rMi
0KXdhuuUwEDdKpW6IvEBl5hx0gBHT6BeNzKgqAKtARRYxFhdXjQYAWe+Puup
euKMj/nZI6QsVLs23ti1J+/CZDYntYVZW0BZqx7ix/rpBB0dpHvZkyQ94gIc
kwbA4EeeWAuXqfkUdRHmd+2/EgMTZd2Vu1yplvPGaBpl4v51B/eA/6uQdV4G
cxaIAVQ7+OPN61Wvi4JWGmr4yLEfbAGE/XhpZjZO5uLNnlStPvIHC4Z5GZqz
0y3jnVFs9R/Ym1A4UGIcl1xRLFZE90ojmQ29SuRdpE3rOkMb23+wvkwRiplH
yiS/i85DI5039iTrOV6yPkLRI1Hi9wfYKK3LCEzEXTPMAwuF5D7naE3vewOp
wBCZEAvIyI5ZtmQ9tgllPMtX7goDTlSEUg9TuVSAQ10vz2ZepGB23/SUU44N
ydDGqGibtUsMbs3Kilcsd5nXeOz5jQEaJ5C0lm4LmZbrhBCAS/0y/9drXYCI
XhvxLFlJ714vPo9OPG/8dLfkQlH34WIdyZ+ceVsb+pnWGAgZjXShgwdg67jb
n2XkiWnUiZ0GEDxqhQoARF+5LkJPg8KH6Ya8Tbr7O4jt73+aJ7DBwSFVplj0
61bUWEtUopalzuF+av3DupZrpPL5tITpP+eaUeazFzTUIc+OEuh3+UnleXHa
UPg/OKsiDgePnvpnLfq0n8i2Khq6poExwvi7+daz5CQxYlqaU6MiNQnhseG6
9xyldOMfl40u3YHQXU2maFAmAO7Xkk5Nb1rpQWQxYSgapmV86RyQOx38sR52
AdfvzQgZ14rDQUbgEsIEWKsS8JgvZAWntUQriBdPI/U8/7tszgvaxRGQFY7e
UpBVDGnLTorzH/Hy+Lo3qcEVqa3TVfc42c8ByFElAAKC7p3+uz7sVpGEEhDr
DYLr5MFJQjI4SmnDlqp/A2m1+OKjinRaJz9hz6fiViUq3TF3OMzJPML1KmDN
7DHb7VCdEZAH0W9uaGDCZQUjtWBS5Yy2Xxrcs7KcZhcf0MT1MF7Kq8/o1N/Y
SMrAASaz7ncY9mTX2L7HUOyeDrCUCpP5XPpodNjWn9Ja/eJQZOek2koin+i5
Xid45RyJMDFzfqgiyBYZDQf4r6AWCmE0LF+554SHw7BA0wx6jNRMIzQXmWUu
wJfdPk2kKWGFLsSVVuWr7AfQaaWPDzqdX3HTfmNjDB/KgIp6Pl5WcCNtOjOP
h7zbmtrYtf4wGvA9PZSzVrbWf7/abezMqlfnIPFqf6hXFKDZ1u1DGhxrgtwB
C4KBDWF7p3MBbQkPuoy0FXWIWUyqTnv1NNYgrZer9B0aVDa1xutY4U2zw/Fy
mZKOnRUN+3MAClsAQ6xlwvk9qC/Qm004JdD5yC6mXTN3glE+jR+MS2xIEEp0
4K6xiAnce3SQu1FaY9FA/CzHs3jmOSy3gvch1y0qb5HvoG1bV5wUzBUqEPtx
tzfXjBUG2YyujgJqE4ogC+qZYvKQ/hGV/Wpvia3GNXuWf5CT52VdsGq1DlgW
MJuYZwqeQHESLr1/grM2p2P9wOV3ws+cAs3vmdrvxzzd44GeIrRtaO1zVYDj
s/6bNjZZXCux1tENjzq2aS+m+rDS/rTAoGtQxLdVIQClToN8V42a6M5mOT5X
rNtvBTR+jMUflSlmEkYS4trYh0QXeeFj5vwbZQ20DFFrYBXJKYxwgo/gGkj7
FkWp2WHZgrBlEKa/52ZZfYqD+wLXSALiLCbzAuInXBLu/PCdGXD89IkK8uCj
u9jr7Mj1DSq/MATV08vI/EEX1LwPMAq4TmK5BkCAI9Tq5aAyU/eSgIx79mmL
FeTsYQ/iT1HhfhTHtN/0VkofkUnoafeefxqCgWR4BO66vYuelMU7G0IZtqIw
2xf92UisRuEPQ/fl1O+F5uLuFoVpXJDsOJ5rGT0uuft0hsMP02Qzib6iP0Q5
sZhyYe3wolgDSRCvjcOqudRzbPQ50BSh2YzGYRRRkxA7b0wuNmIen0qs42rx
OwVBjeP4caJSOxggIEsfLHI3Viy9aSDvJXzlZtf66LirrTBR1RLJLwD744U5
sofEIjJ/6/tEUOq74+fYEn+bzf5TwCv7R4D7CGv6zc8BeYBCcFwCj77STVno
JL4uv0EEFZ5ujGwC6OyYxNBIZSVOPrWQOtEKiC6RcxjsWaru0s2ngD9shR0W
mUyRsGOotrXxKsNAOePZjUYfR2qLwbCTetNw6ToMtOkaGzlkxEHX1hxQqmBR
ehjHkVvm5xD0jiZx5AQnvb6coi9/tBhrhq3+XIukBzvXt5Fq12qk60jCBL8i
Nc9Ro15aw6wcSdQ/pmjJcFT2YeKbCzpgVAW9HLizluCkkmZ1mGAgD7nv78xM
/n5z8sFAkfk7/6VoA6GCRV5ZyB8bYpsG67M4Jhj0Og94ZE6c7k+ZaaK+aE1e
OPF13DTJB8CXQFQxSXvpxvkYQRpP8XkcvDcvET6EdMUmEMRSke5VzJB2x+Kn
y8enqI6873R/ys3qa81tWFkCaO/K3L0YRzYppMBiX+pYbimQPbcx+S/7QQgm
pev3Ez7eF4ZRVR5bm3KZubVEIroEQHpp2kkif8KuuQT6aN1/bySb9qy7Tg8d
NBcU+iQ4EeEBki4/WyvZZm+YpHmStkzAtFsCHdySWR9qWg0XnVdJ/8j77F27
4pCbl4djYdWyVMsOy05N+QvWj6Nz+V/Rp/cwLtAz3QRzIlmBG8KHjZTu3K8o
+HI0dFKgai/xUA4m1hVOCowlUGMz80f4IGbuqQZ5LijaBtFyCsjeTWY9DCNk
jMAIhCcuS0FVA8CnPug+YIWjXFOWzfTet1DW1yDYQ0ycCWP/giup06BapR9A
y1jMNXohUpz2Aw/lktBywhWAbNHDu0XI9fbfhehCnstjqtvqjuOs1E9wfioF
/mo5FTbJBPknOmgnCDtRyRY3MfS2wOKE7kyrm1mI2Lyj+szQnx/+g4c8KGc9
RUsrZF5ccgSsSDnHgMqMrXlCEzkmH0DaBOUvp4neWX4fQMgz3Ic98ePBKbTz
BCINfEV1iaAyC4H9b9q5xBLXj6DZ2O/3z6U0KgbLBRsttFQaYNzy2WYWEPjU
bzhSUjbcBASZC5zvqeexBw+oWLtvgCj/CGBp5/khTeqCPBeBN7s97I7aUoM1
145ERiY4+Lak8s7EyOSawA+zgl7b5QzYw+tp8OJpLaObcS7r7ZQ3axDzbKJk
gfsUuroBoucAo/N3hpKZB/ufA0JWwJGPPDSYt7d85HW3Mm/E0cNaaxcW3iaE
EJUKLd8choUU6uKCWkhRUDCHywEww/iH6e/dbp31p/N93AYaa6aNhj5ijj8Y
gdMRieYZ/DOHzDuu8vnpVoKj+J/YgCxqeIeL29RZoV3WDvnTW5DrdKZkNIXU
Z02ZmgiHCbHJ+UHwLEiXiWMZxHHkusrdx7JIwSM1pf7/LhTrtSLsBK7t6I3h
VrMxfrkINsNxsu+3G5BDTCOIUj9e3evHURYqHVrdseC2cS2sdtuMUg+UDqeh
kaqcAgCA4Ny9ZywgjAI3m8IcrR78fXBr44qlQDzLw2nBiE3m31eQ2bzkpm0+
OZZNpUTLT78IYpSsyhqI2Ksavy9Iau1x1gdmUTHgITZfo2kTuiben1rioAks
b5KmW65NTH5K80yeloMcwOTGZvC3lXY+0NO1UB+FPZvDeVjHVwycRNyFxpHH
r17hatNXNNQnrHe8+TOC9j8iUKOd4sHGyQzYjJG1ALgi4qUxHpxQMpLWBtfm
6b8YfXR2JpSuWfqCOZVl0jtkfiYik38Ww0u6XftQUDjLvLqlYxzlr7q2nFe3
qhJsg0cDR1C36ytTF2Kmw1ea/iUCwATrVR5B3rBnWFe/v8H2OnKRpm7e9XZ/
kwq1LXOZwcoa1gqdVPiAouDiDIZ6kfgtic81m7FHDtv90BNYdmOA49VIplwx
vISwGGtAT0sToVxoXevXQ30nTBU7PS055QcrQb52WugG6gk/5art+akMn340
KzoRNf1PAlt33R+NqDDBKLmWmXhf2zJTUH0ejz2WKT9WxYi3OQv2XVCFSTPP
CqeSJkQrUtGaCV94MEjJPizL2TUuvESx8lYz6i2HWnj1rLjfwhUPF0F3FtOV
0TB1TZgWvJldgURTc77w2xbV9t4TVoMweAn+2g6UzLbyrvbiXtaZM+eY8Jsq
Wz0IIrTDkVaQOUh7aeuvof8SFbwIMy2Dn/JXRHbteBIpHKXPsHNQRHjz0vn6
D6dqd2NIwpKp1F5zRisJiYHQ+ANyunabOha/e6bMvTic7aOb35HhE0exz4DW
lkiTwCuz8VWY4v10O68gT4mqRoSkZ7sKgUjZhIdgzmfbFcVNyAEWjBGt53Pj
SHMsVLjGqc7Eup6ZreFZyU1Mpwp8aPKzfHYKRw37tNPWK1Vr2edxigiQvfXF
hRu7FKZM60PuYh2G1XtfRxGZGO1l/1b7njtCALcl2Me02hacn19zAUrml856
duhuoh7z2XvOxtYHTCVcokCqfqnfW5wk6o5Xo+R7coX89U36vVR7YQ41xNBT
v7WUSL5BmFQ0Y9LUnOqQ32yLvSAzPfL2Tuq5VDRiivaDj7TUPdLjewC8E3xz
EcqrL7DVlkMIgP6vKg2EW4mEjGho0zARwl9AeP6lZs+IaW/7z6zaB5vIzTyJ
d1vwaCa4DiSn5VMb7dMilr1ZnA6NaIYyFvntX9M9rZ2btHFkdBa3pCHZyQtS
VjvaC5EGYU7b89oIOTEOi0ejWwHvpZh/3Lf4SUB1pZdZp70fMZdnBvVPJfEk
iYjjFGMGfeJEA26oYYBsetBvcfwzxSvBMaJaXIIXBbYFzIwfE76bHeFpG8B/
nqRcqc//ADXiWsY4Tj1MgJHxKeyQzOEHyqZMihtyPrHeHtRTmJcu/5bKnEC5
2+9AUl7+h43RuR6e530CSwsRTZhKN8ELai5oWm2qh0rf0ohpDzWv6HO5exY+
SDQwp5AkKOtI2rLxPCJUEIILsBUHyScR370l5uXCroXKcA1hSzHz0vHz6yhC
xNoJ9d+vI6IS2VhUq2bBBx3buF7oFMf8/stcNynXDWXL0Zu6zcLLDD9EB50d
37iHEgrFSOLWUVXnmqddLRFrWC6TZnj8NRBVAwc7D1dWEUg26kU6kJv+Lh3X
ZVeoVblbEhezFc8u3KLfuVZobuL2+6BOwl+CJTvcEMJ7a/v6I8frpqYnTy0c
WvchIWDVz3btE3b5J6b5YiN53ISc3WinnDs+Dg0vJ8SQFBnQP6O0SrT5uuJS
lEeKgx5n5PA872Oj+cruqyBWrsoRM9mxUf4Wr2QXvZ41UxLSj4QVYqyNfUip
RAU6kdGqBAzCAobZE86G/DJZdVUwBJmZ3WsaB6YAhWSlgKcPrJFhMGNy6y94
udxBWStAMXh1C+rr1nP1ze0tf43KDz83fONF40BnmsYWXKHDKEdur80X0hRb
Jgd7AI04pAaJaev4ffVH7Fkxy0+Ccg5pkb2cVvxEX3lEKAr+jVBL0WfKlhVS
W2kJN+35jK7Gtd34VeWhh0JnENkD1zQgv+jaMkwg/B5Yqk99pLqciXbt80PI
NgrmdVajfJkLMNDAoILZ/l4O0axpNpp7AOD3cAA8EEulmWGtjQ5Ku38pxF2a
2QfFhhx7kFLyJuIDV3sCZ3jj6hVt+o1IIT0AWoVk8j0CsB+cyNikBk2n6Cm1
fCFLJhaito2VmjBPBsp02lhPZQMw7HglXwPkg2SBb+B2yDo3IY5FZ1S8syHa
D4TkIzMt3P5J+boUf/bjPjT6jX/yVkVdJ2haHeBb/mX4L5sUhK7sdWeUGjs5
vLg4XQAQg8W+V/lRnLDGAi41sGbnMyusLO42KPw+9/8kTgnmEWJVAn3Ug71X
TLo+WMXxrag7Mr2T3haVjXiiOyfoX/mcz71TDlCmB2h8IgtzfH7t5RbZdO52
yNo9hWYoQnFYa5nmTYezWijsJh0gct/TsEvP0oxtEhxCbsa18ZLxz7zK75mG
q7p/Xnk2FxEFXF7U0YJVQ1x50Mw6rWA0qH5DLJO8I9/JCodVoBzO3/tGE5bu
3XXKTxu1jGuBMJLYcY/TaPBHJZRDoasVo4Jdq8kdYh3fSKeFisxBIri3Z+CN
BooS/Haq4UA0bGIrVDWiVqxKyjsx3AoVL8rlHhCRBuOWpHNm1QEAqfP623iR
U4A4t2ojQw0OZE34baGzaFXIPClqFAhcRXjsB522uKCLt8Zo7tW1Eu70AEGp
8R4KOW8JwJaxQwrCYlGfWDVeaONZQ+IOb7NJLlvmLDst1Mowi3FCZH0IzSlf
o9slpx2yc6yPOBQ1TAQbbqvWpM/zmtWqppEAggO2eCft4ZxOUkzICANEU2Uh
ioQbcHK7LZio1yyqKA2tzY7J92Wqsm9VOy/ONYPdrmHJtPursR9cR3ZIHgVH
g6C+1oSgtgZPT3ysapDLAOuv5BLbT2/nIibon1kIl7+DL74uAl46xGT5CCYF
+PvmGdp6IKb2fMsZTP+WZsNpMk6py5hrit1xtbE4JIPgkbhTfQ3/IeHv8rKz
vy/jQjs1JvlWmzxlPaPIOjInJDTcYFm3nieahsVlw67lMDeZxWIux/PoVDwE
lBm6WpdRvw0RIQfB9QHMp18FXy6yIec3W9PI/+I8cGTySUJpQdlOficePC/C
Q50r1LmjfosP3iAKTKI4HpWjvYQc2im/O4EEXB/P8A0cMdrXqOA4vFwxu67X
qX0/vJ8C9+Jpn8tiT8PnC4WxCX6wvSm6UZdT3Ia3EeiHvepL4WgjXVsXIMyY
hdx92IiXgYR87fvWrFYmGl4r6/Qa5dgZ4n42EY05nFrA6Bf3oLljTj9ZJ66Y
34Fa5akC9K7bjzNEcgdpKiIFou0tmVtNzqLGZ86VbogEDbIBhG7HI+BWFRF8
SsrO6Qu9+RZP0x+OGdKqwcCXWwL3jr+gZawvX/sD7tzK6oFT7i2YN9TJtabt
vUfiFMQSDeEU8/YnvYEZC5J7l6gjzUH9BfqKH2sWmBnVt6o01HH3ouFq5iQR
qwadiHfhLx8vclHIi3ZBOmsPFmQ4euV3jkO6F/SlTFkgNJrNfoI+/QSrRw9o
H8ebNRDMOOfkQjT4bafFKjs3rto854w/Eefy9oqZb3TUBAsrzXjEVS7JBwif
wut1janW6/V6++B4U+omxPWaT2BrQ/8pCnF16JI6D1oybFCfpC0ZWqUQmyo6
0pWNujt/uhvGLnoS0XSBK4qQihQeitOhtqGTlSvw0YOKZhasZGKVc6Rfdrd4
Ufy4nci/03AeRFYZVvTGVbJYF3XpEbfPSwNAFoiury/0uRdGyBrmTrdOAWqW
9n7C03b8r/Pv2WEfOH67zy0QJLyXNRhn2xz4HzkEwrY01bAiAE1iuytGyaiS
FvgSNIsUPjRLk8ZMNmZSpbZJ3BH14TbJ0w9qE8DjJt6/D4CZpoNr3Vn1mUcr
CIChoHGKf1P7tda755+/x0y6ln46njLEFFif69B8D8/oZ6Q4Jioq7afdnXOk
UZ6t5aH8PvJgmEodu0l0tKf0P82zhA8CmNstVwRQWuJH5bA28n6XqAy9tuEv
Yw/4Kf1UYoDBP0Ssy4ZfGx2xtXEf35tGd2gsjgmxZ7ZwBPcWL0RbO7uu1o3d
TqkpWLl1vn2zv6/XeW/wmXQUksj8zqhpkUtlfjVBHbp+YPwiGZ+CqMH3f7aC
Xz46tAhMv/K/IXb7B8MAezQ4vWStEOhmXqqxOa6VxkAng8dQGqQzzeCIbq40
PqNtF8MGV6PLlhe0Z4mNsYiTrpFLeItY94A3B5dERai16M/plrYmfm4KrwAm
iq3egGHbyusDGKxz+dZJjUbKge9ypvmKVYktUlaDgDD0y+Ry1qHjiESXdrpS
tQQwOWWfg+fG4KNruzZRJKrm8oxqfw/PNn6a8oOtgphaHUrZukq0Lxt05N1E
1EneA8HU+a9wGUHxWsyNvNHv4FFgNel5zQITGppgL6QCg4+USq88PkY8GFVI
rZ0avPEjUZH8mN1zNl55C7jlQw5qLDlHM4kIFsJyl7gZyYbQK2KiPQnwYjtJ
rbpz4TG0pCCA2IKjWJOlpsdl6sorjua7bIMUqDcFgY+t6GwgMcR6SZboQe/E
R7oJPWSO9a6CzWZ+u/ir7DaKhxA8WCZnZ2N4391g8DWHO99vcVncENCP0pJD
G6q9Rm1WdvY+1MIqxpLBc1YCWNZC42RUFQzTdiBSbdeqZJ6G5SgOnDgEHZKC
ZMlawuLCPSS5IGwTRC8o6BPrM+iYf36MDDEo8KNqJlIfUlOcvtAHapw7dI6K
bQo3oTD29qydsKdVRc2JBMOfOlJUwK7BkdZSgJp0kjpE4WMFPobOZRZH3e74
5yqSiUegqh6PPgfzC0TEP9zLVq/xeHUo1hrQeKI7tdxxB8hadeWw2tEoJ/V5
kOUnEEkzPgD4bAl9CMzz3j5FM+0oRZAxcFCTIeSzIPXFjk4Yy/rFuuN5ZGgE
1QvI2VV1g580vw+mVjDXx8ma5sc6IJqc0LdMGJPTJfoJluFjx/aLcM6VN+RA
YSKy/1dl88Oy/YkdE/yM0WrqiIQ2uUtDXcqlUHgXMcN4mhv3lAPoVvAEkhZh
JR5o2V+q1eochA16hPamhm5QrSRyGncm45TjAlE6HUabdVU5fNBwrRQ4fSUV
zJWac8v5j+RTypp6DudST57a0dAfnG4SLhVqbvWZ8quDrK5dnofC2rkJXxrr
cmiAeTzIC/7AHBRuMVGnZqiwkAnevUetEvByVtewKy+t1JqffzZCJui7BK2N
Ru/xIXea3Y7g9u/pixaHbeoovDDAHmC9hKrNkamJEltLgqltfcrdSczJ7aKL
56owAqTRierTCqTql0k0FD87Xki+ho33e3keinmKbDaTpkokZ8b0DL0yXn/Z
D+pS8mecAMhIgLAgrTEtMFfI3/l+dDBQpAbyv9eF9LBMG3Qqc8id+ZW9TEju
1Vz9rl9obLr1mfBrUSo+2hmKAMC9zeN+s7LCLyx1XV5sEmi4akdUZavLp+8c
psstRJpF63DM2iffqzMmdIxOGiI6Ryfp3CvNZDqjj442MrK5hJnaFUz/mlEs
ATzXEPJtMeTdX5GrMqE0OcugNALQPukkaciUVl+DXm8Lgi95GJtzulyxO+gd
Ps+J/kVxykQ06pZrlnz2bwdLu/l8mieFzF4GlCEILcXg/M5Quj/rv3kQKe7o
E04BSwcKT56fZArcKuPFswQ2VjzQne8e+fvrZyGdqW7MjidobvvNiaFKCoVB
J+iTrm3x9MvfqvmyEwb04pugozILdvnivketjWVqGRUcGTuVTp5hIDC9nd9M
eYCRBHDoUVNSxxU94wU+giHV6Xs/XUVnlf5WBlEQI2m8tP5+HfXqWsOlHak/
xjhMhW8yDwiX6FyQp0l857/3DMe/yYuWSLN1c65Q5z7VXRV0WP8fGHwXzRQp
XixH2ZmFbg2RxkuVuIAC6dyoyQVYdsTaC2QQ93dEwxZsAOE7EjulnkGrR+Om
UBlFRT0edkzelEv+eV3t5JpamtmyNsoCMF28m+KypcWD8teZt037obNnz37J
oyoad5BC+0tCHtMz2SvilyBxC5FMmf+v5a9rh5ewCocgtymFmrM/jPVTMshN
5Ea8erWZo4x8DtyMla+dXKsKz1L8X1n6qsDxJSAMR/qQKi3C0fysiA8b+m8l
mIh/e6dEF4NcQh34ZIb+H/D/1cqqJzzt7eTTIDtuaTjgS1eOh4CbTPaRLywI
tw8F9XLaQORLkaovNwKtwDA9cwvcbpq433eb9J0CY5cVY9tbf03AaizPqRWU
8yKFwzIMme0JkZBpbqmP7aXoMkAzrjkbJS64SYfLL3N18sBaScfBFVsKlAO7
pOEJduZDB511p7EQSckAnqwse8K18VPGZxQmkSu7i+aNeyTZFekIm9HtYDKO
kt4SvBSqOM5//txvo5pNsW3qdbsqOCe/rXMfx/xHEyPeRqVQSQ0K0Rm7cKnB
XU9fI75y4k2toD/8Fw5Wc2op7SVW6kgDUKXDYv+NTG4BmSMikMNCbEjTwlz/
jiYchbOAhTnqkjlYFioS770KaF/jbS3l5Grw+2wOC6o6cT7hBPw/tJSKgSR0
c18iYJ5XJIIqmuBrAUcuxNorp3wIrrSbsRMlOd+QyB6GbudT4Dl89cwynPa+
3DHO5yYf1yEjyMhfO0FYPYnbJea4ZM8Pch2nQJI9jTWoHKJ8a8mqS8DqyYOj
4OOnpaZVYH5opDc7n2epd906c8e0jUCb7l5k+lMV0S9i9+A8ejPxfLDfOf17
kgc1p4T/LQ2IE4YOl+hUHcdQI8FQa3ttmM/8eU2JpUIxMdvLAPTD0ksGXGCu
pJEOahWBLdG6sTyvj+hXzAI4JXvjYYJD9GhpNhbT/1Vrr1EQoYLQo4CMQl5Z
Tt2DcIygoTxEXOEfY2Wd6ISF8zfkBiJUPtvzasWr9fRxcaltG5NcI8DWKXEp
PPprmLAH5IeRTcysxaoZJ8WnChPicQfdb0JKvX+1r5gWAF02g15HOxOVfmRp
nt0MSKplOiyXUaqnzEaZO1eI90xmXNKOhDo5P5nQcXrIfQbA8jYvY2qZ6c99
e58+5JZihYHFvQlQmX85anw/nEUYFBC78FAAo4pBerEmTav5upjKqgJeXUQ2
BOFC0TBe76CmUqVRwFSs4PbQvWTwkzm5GJm53b3raNCrUaA/GJKrMAIJkbBG
7RhmG0XZ+PZpbo+lXtaN2zcNaq5BHSHW51hN4jemb9Jw6ijj4MP5DsB5knPH
8CzhkAVdGEqS7T1ouhqcsPzN4SELk7B4rzimGiCROzyIpyb4j6ioddK5oWq9
L9rdrevtaEc65u0HesV2jHQB6CEWlkMKppmlCeOLedbUo765EQiVdlIicdoX
NQ7jBydJ7QEuiY6mvoT8OYxIrA6Epc314kplasyuhSCL+MfCB8IB+ZckIIG0
7MZ27Ut7mSJG32PiY+21GkIr3OBHWpjTGH/INlkm/HmjwSICkNeyrwxT6Xvl
IPObghZuBhFk+CdTK3diN69/mt5pr912Q/yibQ8nvHXgAM1LiS+vp0nUJlyg
K87taVfh1/sAtN+7rl36z9jm6Qb6apfgOWhiFy8Q8WdAK5YEKw/dQ/eqaV4h
PwOMlg1Ny+2qFibEs3Pb5EgsL5cd/OicPVbhAPhqetBjpd8iTzneLw9Xp5UU
g5ep0mu3BGCGnLDNXeQ0qTUDOVEEXTNOQz2Em20poQagiWHLt1ukCq9L4ux6
B1L50MV1Fa4HD/2muoQHbA/4w626mz5PENscQo/mDG/IgGWrTVKV1Od37Sac
paWw4RiKwZoXusSyud/soS2OlAvDSRAkQWLE8RvadoG1WCbO5f1THqE137On
Mk0HPdiJGcoDRgjqUeQR1chH2A/QGg7JCLrNw7skEVlqAyhEOOhprwmMTKSx
8qsXhUrITM9ze+jttFgluOqt5N3lQJhnE80RKCnSTjH1O7liwTyvNnT3Yyl+
pQ92sanvUHkS4czFT9u0q29ddWyRKzf8T5LZt67ROPe0V621azJE2MQuLhCo
4ybZeYY5+1p6RxHmF6NTSxDWAhewt3MgNBzK2U/7bBiSbvuYZ2B4grL+c4Cy
c4oidPWtSR1MvKdq+D/iGCHCQdCgWKrpl5bGxbQIq35ZzVRMmxF4rCOlqEIW
Nl3ZDe8D485hOZcuVxVogQDRUDS/lSrDJOOSweAbC2HMTiJffmGexIG+Q2aw
M/x/fXPKpTYJcVQ6EXIIGfXjTnvoU3IpfxTBkfCUIuFUrvM7C+OvVSMtpwEI
ZkvIos43Iu2so2ATNG8WlV/+fubNY66QLOyDbgNbRUsc9/4NA3UjWbzlyOcI
Lf34v47tBqFkZsl0VYVaLAil6L9aeljkpHewkwEOeSTOrmquL+eXseFkFgbS
05uLgJwuulu1lB1FXU4d6+fRYrQs3J0FUBEM9lMbu+mcc6jkD567wKDUeZd4
Nb5RMqAZXrYVZ3fWeOmtsOzKAWzDGet59IgMU2T3i8POMJj3VF/NhaXA5z/1
kKHGnvI/5oqslLBNgNwyUBlSZX0XFCYIFM4/raMB5n/ueICS4t7GjwQGILoW
mAtlCWE/tVptZeVNyP1yz3zIE9VNLkjqaxTWQG7vvecW4ykcKkxnz2jMSkby
d5F569sGcgRQ6tWL0muLk5jP3Op9ypvdi9v+88EM9kenIqI6CDespEazs+SH
Hb6rH3uyoVJrjAqtS9y8n19dZeaNRXDsFkDnffpTRpMDcKsq83KBEM2stkii
KmDED+rOM5lk4ScY+UzwxCYKykc376CKbWxVIH4vcWf8Y5EVs5IRTqsOEldp
Zzd32z73IKOBeMop80adv/S6ez9u16DE0I5dv1a9z1JfNMWdndYqfTaAZ8+7
02jCPfFoZ7kvD7WZ8shEhAsZneWPx/P3jzwN6UBUuUa2ebbase7FW70gy8rD
jUbylDT3bGo72q8YvQNmEd2BQOiedPwn5p3htdJ/bHwlxZr/d9Tnb42tjnkM
p46y7WyO0Z2XUIDUiEHOX65dSGMJotGqTc5XVTE7uNxVzzGf1OCYu98mphsz
F5dQElrodSJrBQa+mvegnS5N1+sQT1dKIGnt58P2D72GuWWwOHyRQke/QP9j
aMfN/xL7I1noblfXDOD4P0ca6inFMCzHQji0K2ff0io+/JHd+dRuhe3X3XR8
Q8eZTvDLC/4fPE9sWNhqQDAXzPcfF5ugZ42+ArApwOi6MZdis3Lv2B55YGUw
gsJPn2Np74pc3WbjKa2ZJMvNFGfwD3IeujOjsda+8zRNdm/qs4u81kx8CFwJ
uf8CaAELB5iI93EUIIGB8N6ET/6GN/OS6cGz9JdHUjMNsRW2XNp+x9ad7YHi
UE/nxza0MM/BEdCQpKOf4FLKcI+/tET2JRY/JimHw18JH0ggdh/mvjj07x9G
QtAmIWEl2251msmNznyzdg58XO2KW1FDTTXP2pMfHn4Ue0/kZsg7TtfJchoN
XfMdqLx/saYjFA9ocWKOQMROCICXel8SlVbQ/ZUFii0TWEJN7q2mAVZfCMZr
mdM3QlEbuKtLvLX4DhZ7Vc+lRn69QZBexq3GNhU+mPnBB7vTLYzHYM1Fd6vl
t1mHRrHgOF+itL8iw+MzeNXL1OnzNohZ3XVpE127+tqAcFo+clF0UbP7ku/o
KGgEs2U833Kj3hjANc4jPzQHlA0ic41GC80aYlAkiZr4h3P/tt4KrSLFwEU5
fb2LdLi1yVcM1oVEYOsepjlseTu0l3Vd7bp7jTGNPjfXn09NLo7lFMmxKg/G
2VInbV0N7riSTsBPh0su54uhCkDrzHHFVmY4ccWIEdgSVt2Y8PrXW3yQ4uaF
qkhIKORAd0q78uuijVomW0sh1pZKUSU/g7ZccSm0BHDjMSMxqpsXQJdgSfCn
NGkcKjhQlS2f62eYHYeVasPAyWHaf5MV9rC3xMHRSv4OPV+NdfQIvtQBriC8
bZr9uacrY84RrmQMBhXR1J/2SVZlvlAvF1TkuBdweKbjRssXYio269I9F6FB
LIrkw67lxynmRc0RHV96Yxrt6dE7HfrxG2IBBQHlmC/jg5bd5fu9mS0MsHKo
YmbwgoYMnY9reg4mHGH7Jh3DlgOOk/xBYDEKXetGsvGrYG1RCXGUFdweTkX0
wbXgA7ToGpU5Pw8YcTgPLzxG7ZtFX26bBYasbgrxBzSHZH/CukowBoywAtqf
u641ky3YVe76rrvIQpcN6ULOq9WK0WTiEWqGCKYQyByNyxOkhtpKZahMefjD
BOHwFIbHaYpo5e8mIih9BMbaWFyvIgoC37+HlPQmkeHPwIvK26NBeYqNHSlB
bHOAgr/Tju20hKhFJ98/5/9nezGNe8EwM2LEnxU1Abn9QUtNdUukJtyECWiF
4KJmzPO+SU8m9s2HK1XUvukXIKkDWTLeikODZvzitxcxukboXdIsIYYRLSvq
5Zh5aTAqCa1Av7KsU3OrxQQdQumTmkYbmyd1cqNpFCFrRiLRCaP2z3jXoogV
6HVsGab/je3Ghx6Pxr1qs9CmMbSBeT5m6pAi2xO/ikm97BNKWX3BOiX7lw2V
Ri9CyBbmyItj/HKUB2JBAxWtWsT7DRlahDDZACxOrS5nYteACojZee0YBntY
vW76cdTOqXYSYVx2JfYkXhLluSKR/zGxlVPorgqiZY8jNXIt/mqcfxUhVb9f
PcBev/OD13y8Utq26bLO2prEldGagJ/n6UOJZOx/IVyq9w+dw2hDQeahHpQs
IYEpqS5uZwKpMZgwJKaNcuAlseI84TdmsIIzPlap7ZVqW9EzmAPS06AAkIrn
aMUSA87OKrurIrede9bprPs9Zew4nfxDObngofCKNB+1zsXZ3rEKUfNkUuUN
lhWFICQhmao18IB6qKtZPOPHXed47tZmcQm+wXA0sv2D1UnQy/RXw1OwCofL
OCIvPt0HgVklRPz7Jbf3WthvHB1qlW+fXd4L7Y6kYvIEdJVDMa4eQfdX2jCL
O3+DKv2Ids8QTlmvG0KPgV/JORz7MbZIST6i+L3r32KKCezI7Dc3QAVSsxoa
HHXg3Ecj6f8Z/AzCtSCtDAM7xBtWnCvlbi5NT3FBRrFeGa/ZOVums9k8Mpp+
CIKz0Tb1m4kEbmPZlqdEMQhLwpdJtDlUil2kQi4CGhx60nUwEIkrpP9ijf2i
vdlUM1NSIPhnFOKdavUsHYH3NeyT73tpoyGMXyR9abWAkVJUafmdOW6LEgXP
VqU8ScKRX6WZiS1ZCsUVL/Ok+GlP+zQ0gh2mnj4dy7Zka/mpTvZh7xSne4J7
FbbHAq6kAUyLcI5PCFfNQ0cwW5AHnZD5lkSYCNUtIPJzWt69p7v6KgrQyPz2
uiZQ4ApX4AkzrJQR9lBWVyvtmLvFe7ycPDryfgjq+P4HT035Zc8daWNAv1QG
HOmIRiwuIEGlS3XLL9SxPnQmtGbfM83lZNY2oazpfIFCfnIcf2F3kgFdNMAc
4xvZCJ6LL0ntUgxDguzyHw/02QqGS1590FXM7whjEXExRqW5zypR3/joL3Vp
yQfjDAXBMlgSUPDDY8pLZfoBZnyZEZtI9hgvReuGxBqG67+NHON6+RDuXFGi
ICsBDCwFvjDrz1kfKK1bI+ruPb578CUgnQ7/Z/JzenNc2Zl+8BIiDuy9lF0p
FAgh6NyKjk0VqRNjR5pZ3IvboR2XvnstP675sRTvmcpHU8I8ULuugeHrB6x1
g2mEQx/c5j58O/M41NKIIkTuKiIgDWhoDFwrnzk3c+R6OptCiD++ndfzO6ED
2IGuAoNu57X1hhGbv2LhtOmDznWeUInxge5tII3nPG/V4PU/zmwZfc42VZMc
kqka+WtKsPWHn9nMycOqFGKOAt2T4BnbC/BtxIYcXtjvbKyWglsP7izCGrHh
0DHC6ryhuYEdBo2B06rNRRQgOrxxMmJbB4kb94VAVxCkkUvHijjyJdbgaRUL
8tOero4709X+lo5khhYusAcSCwaZntqK9e2wqAkmiJZmYMy7e5uvReSnvpbT
RYp37HscNiMBDnO2hY6Iw25TfgJe7HUnvP2/8IopBfLaU9JRlNfeokRMgGXS
FkFvt5UED6jSAGv9XChJCIA9/j4gxMaB4OjkgFyO3bE14Vd9H7SDUHty8AyT
pE4HuvQfcWjAuFz8D93gxcteNBoH4UbqnLsa2bs5lg7P7fDfBv/Erjzv2U+2
MzK5qqarcUecI690OlctA5LVS0uTrZTRp7cXKEpqjxWMLJoE5JSgUi85Kxwf
06hylobdJECZ+Icrz622nKdZnSWpTF+SrKNp5ITV0bYfgbHssLp+ChMJDSgL
laGjuuKY2zn1536iCl1HY/lwDfxt+XSAFWoUreFl6PctllX7CqCQTe8BfaCV
5ypGfEdhzk3b/zM8WlDtnbElxXO6X9RTGLY6VUk+DnHE/qox/XGHJWfgjhZr
y85wlMbOAcanaEl7qm0PikpeLCvDpHcP+tQsMIvnSARHxhWJklUpDVNPS/Qp
N/RemBrGB2n+SDVFtplPJZxoXrr0cG/WYjLwZhnOSlgDpJHa8eXUWQtOTRjU
ng3nsUOJ9jlspUx27PHltQ5xfEg2IBXQlSGgnizSaQEaEaeJ9sfk4XNtC0ns
DJwgkCwpOEOw1rm8TozzyqQuozPGZk+vgZZpGDJhUh6N2J9P8UK4rCgC18rm
fgKIeQoV/cJIhxrTGY36hpGO4STpeNP1mb3BFT2ye2tikqfh+toq3v/Ai7SM
W/7GPotWmhTcqYiQIHEcKhH1V4ldknhp/g2zFMOi1k5DI9PsJs1mq1UIhozf
q1C0dTUZj3c8bohfB1H9F7PHRpyjvE7YjzNXAKajeB3JmstuD7vylgTQf7KJ
2Y5zdM8YQUgX9GavA2xh7NtHahZQBod3yQ9ZxOGMYFef2/lsiIi5arEKO64J
qtFYG82Idg8sIxmgH9HClCmC7ZAkGEcL+GF/d5rJHKi4+W8fYXLTypjvktOc
Z5yPftlH2UNEchYTm3tihlWbqNRcythklxrkP12/ULvgKO9vrMmAo4sF8jbR
LVdu740YxXMiWBXt0qyIAdwWy+dT7kIQ/kM5aZWfyOWj4D8kWt4IOL0WdGzU
bJVKw2zeABRY+RVQCIuVnrJ3gcJXCCCoGPRERtdgrC8N+uisgo8GwXySpdD3
kvwfxganL8+gK/G9B4UoMINjecoC06f72xKCLLwvko8uOdVpViDq5pn9OBe5
GmUC/02esHdobs0kLZJNY8J9/UuFDWisj/RFAKvJtH8MtqMLkRp0FZLnIQdd
ZqVqCcvitTbz/Wz2JQIjb0oZwri1BhvGZ6YtvubBxqLl5iCvaUj30PVvxELg
4Qxk85TER/oD0idsM2DNv4VN9j9bLhc9fCOTkr5H/QLYZwz/BOmJqUy+Doup
JuGKQdV4xhBEJSqUON8OvoehGnlhHszjl8rLbSJIpeVjQ14IyGJYIAtMVize
VoLIgoF70yREbW8lHTI3ckeFjA1kBtaevjqAlv5iNPYJzhXU0ykWEjabaR5R
4v4nClUVxcRbUNVbiLtEx0+Fru8VZeXiMyqBzB8i9tFAOIeexSZjz2ieNrty
Oh15SEzm7C6pEjpsebvArDQwJ5suCNu0msgbRbKiqngbI22g2ElU4jUvEtip
0nJehwHEyRC0J/zwu1Nv/L89oY9UK1F+o0H/NIZ16a8GknOU2nAPcChUubp+
d3DYS+gju7c/BBtutwoVACoQgJDbOGNTEKnZPB1xwINC0566VvKABCOTYjzz
tuEdYUCJGpLYshGWvAoe7qU6jPSruOCS5wAlVFe+mX0kuKrYaqveeihwE80X
QwiDIS0nvRIJBoNpE75bLKy9pqAfuQbBF2wtthcZfDJFoHTE/AcRtX8XL9PS
9z41M21/0uqPolD/sBdHO9KEffwuoUxAYbix1gTPKWFdUp2J1WbJEVTiVd5B
uDRmW5jUXVj1dtorGE78sCSa5XvaNd1mkRc5BEJgXtC+QldZ5JJOUlgZcoWT
fJ+kQ8OkM73CsBsfat0Ei4osUjo1m/MRCIaWVHn/qidRRDVESV0QXQW39PUU
aI2ZxEq80opsNGtdzdW1RQS9M+uUgk9QJgOy1PiB1V0V44yFdnUHoXaEPPi3
1xI1GXrMePr7Je2ucipNMD9X6JkiJez1u3/w9w0EtjhLAUdTxPgm9y2We8dg
X7wUIaA59DFs1/y9BSTXTjAoeFJs9/t6esaHRdw12DFloJQLSsSxVWu9+6Zk
4GdOyb+EK0vDu5OIhLx3hrNCmv5WDbCdI1fO/KbexVJeC9Nb8PqCJB98iX7g
AVwmH2rvWZH68HZw74D/IuE9vlSQgcNHwTNTRiJIx1xsW5hspShbs77gnYuv
Z6RdNTqVDogHwYur8XpmFWFEXcyCJc9H7mXCVv/eEeTgidem/C61n7R2DXWd
V67J7XQ1EE00300HuLlj9AEi3aQAQgY0ahKNL+4GQUbDV2F0yCnRjPAGXfHH
k5iAcL5kYfccd/jZrBJ18Pd7Apy4e9NYq/GG4/hyOvs0yQAWONP1H0cnT91o
yBJNqKjy05V45t5b00rpp5m93h55a/qDl7ze7uFSyMvOTfFfEzsbhKZcd36m
nnjM+iCbFn/g93MpNdPTcNfONTzRzIBNHxZ2lfve1UJYEy8awhdKq06Qtck/
BPuVfd3k/HwDGKNZ8662ofYbFQ60fpV/xI2lJJBKm4DSpDvd4uy8GiG1OMSj
gDZktBxhedPhTVZBbcoSrrHrjQh/SlVuyAPkAU9oqgRx8Nf2Q8y8NePU7fVJ
JAQ3fx6KYFzV2nW2QKvXi2c0+/lmCcBpQJA3mEXuwsgPL6VtOxzmlJ2aVRZX
dsOmPgfAqmitjZJfP5oMdwmEiXQ2EHW8daEk0MX9qSBY77V5e1zo2RdW93GM
8/ur3LwHWU+LIsPBU78mO4nXsxLkz7NKawgLMHQIhQ1liMtdYXKmHCMJNX+0
HBwTUwg14cs5EHgRMBz9Au9S3vqXYu7vPuUClnJHZV3RvxvxeXID8P6yO9w+
v4soHfT5Zs4hkM2UYLWluQqDzDbGFTEVF4fD24tUhpWPTbcUL6FUvE9+29Ef
MRbbaitwmhXqBgsDS60Q9qabe9ZFqQDIfkkYx5ZQqugUcnqGbohb+HKRABWE
Fy1gwNs4ZLxm6QiUf50Qrk1qVQKFxHQbODhNkYU/Mq8MdJAP9arssX4oNflq
eG0590UFHdpomRGZeSBFK/AooxMmIlxKD42eODXPgkiEUXdoUfz/C76VJsd0
M9/hcau8EwvKnO1FMJcaASGLQVbp6aNJLfHY9uWbcZQ/cDFdFM49eD+B8dCC
jhl8Ip+zhZqM2bzjRe+nrjAu+ZzOum7g3T809vpTH0GYYKB5nHJN1OP5CSW6
MtVu7V3/PEDo+6riH61jSFEq2hDVxC6gUatyCl9Pb+42XOpGRMnlc93p7xai
kLtgvLnnGY2mJlRk/1STVrgNpccnKEBSXkBII6bI55bXmQ8nudOgU8BO41+x
5z+CqiejT6LKz+g6mlUo9YTNgxZcwXIr7CuxTrtClqZ6YXnNuW79L46rcm+j
zhEJCA5Rhz9v3pUL/dwIjE94RuyuaJ8wBNE0Y7Su865nGMoUJU7020KFq15k
rZrduHIGuw+lOUpTeg0hMcSL6H660Y2U2T/CQ9+wvwfXfnNY3g3T06UNxOrI
2n58YrTt2tXK2dWGifBcb4M3Cmlo2BiyPqc6r4lURxVUn/GU48s6zj9bsr8b
TxzTmTiS09vWKxttiDiXBjsg6yDxim2Imyfkr8jjPKVkZAZVZi06BQwj7/lh
f036N/D9tFMzEZdRfGnMIhq5q+Z0pAw9yNAjN6jzfDuH05z4BxbvyXMTLdWU
NbGiG7vSXeJ28cUDulmUduXY6CM/xmnvJYW7hrGWJAgr3txtelDWxlyb9yfs
8NKR6PE66m926z7CjxbglCZclstT11fpIh6fltcVNf/SHTkLQMPIg5zwVbPY
4czhpwxUpQ3wOeDBi5CH4oSOk3EloHs0T5jSOTKyrl5ps64ltjXSbdQ3LxKK
wrHRvTfWvPHB0sCR4ZoQeJsNY925rUm9lTI6RVE8gob+P/Hk0QWk1jLI+6Wu
u2yRfwKzSfaFkHELDv3bu7D2V6zMzKD8u1Mcjs63hK/9mZY5ha8os2S6juH3
ygPD2pNZTHg9psb5sQ0phTTuO93h1/XH+sIOXJxrW9iGgBpjI6dFzTp484jI
kGP67z9SGisaWIqc0EW2aCukB85YaJHft1UQaoFHkEfphBBtYsHgUauPoyz5
lim+lF93NFQtEmmdRpnSrUAXl+ovR8Q7vi5dVA1Wp4DWmtfgqpwfWahZsK24
6WBj6DnbjlLCJDmlq0a9aB8IlV9DaX7LHukIkMCTlUX1r1U2kvIY8Z49ytmL
ks/5+GlKUBjHrVAyM8UGhYfDevrTW+ZA2Nma8ILW9sNVuo/N4EvULllJJzbo
DJZsFnqOlRcGyOeb2IwQ4oK7L7Orbl1zAv5x8bPnHlC3xHnc9FLr/O4r1sGb
znA2rFrgxiGsKY1rCDZdUurYB5wJH6a4fA0+ef9gMiNNKkKagJc8y8P5kJoN
MeT2VpvrGP21CW60EWPQvxz6sHp0tFSkPJqXZHTjUqq9dEwdWMC3eo8xeaQK
V0efhZa62oYtYWLy4r5v8LIvJcWYhcDqcggT7igur3qmbHvK/xSB8/6jmcfE
JlnYMnuqS9J+9AC91Xsn/Vfb5YbnPIcEYi3YFfQuV/+E3gbzNYBC7aeDabj2
DtEwP0JvkFd/y7CNmwGXkdbjo+m+5Nt9tQHcuewX2qntkB6TqAo8Wv8t2YE8
kNlq7ZBmZj83of7J6OVKId2xHxZBc79UDYtUEZWzer3gZMLGr64VcI32p3Q/
XBLRLMFO+Zz0swFl17no5IQJlEYeC4mAjxBUYS9ilwDovBA4nKD61SwkgJ7f
ap1DBWc76BU13EuzB9jFk9iO3gCnycwkkHI7UoraF/jENDBXA9F/KkTF8ar/
1pto4IIbbVXSzgALW14/GG9NYGMf/w4uRLlyUFAe5LkCFj1zgDlMDzuYJcDp
OKUyVUtsEcXWEjKx8NGITAgyhV9NgHFcKkn2fC52dGFPUn6mucBi5Xxu7jrh
rYwUoB7UYHSLI/B0knY2Xv956zdwOnYeOYoztmXDIiGioRkZcb7cm/pFylP4
vnDTTuRuT95lpG6qM3d6az1Q5oE0N1ERU0RFfB4s2JvkiJXkXJje6+P9i0I9
DH+9hMUmprmDYQTsLLJfHpn1Jo7ayCP699IJpGdecn5n1s3hBf70HmjAMXO6
aMLWzedW8IJ6ZdtwOw8WhwU+HKPw/wbv7BGP6/69DPPpvahnUdQt5l62M7F9
P2W7W1AiBq5XDt4QgbYzbrh0rPeBcJYknn4wzN9JNR5kdTjagncetaFUA7k6
Sxa8JSzFcehjuG8az85fk5vxds8eydJnmZcDHa8yY3PHIkXQ4HXy5OlHz9ET
c7Sd7bFw5PypanuDjSAFWXYp4k/QH+DBCnF/RV+6Z7saxDlvk9TLwfZg763x
2W5jI5Vu3U12tpBuJI+eM6B8jxw4pNjMX1Gxy37/tyUQ5fxHfUe1CoewYTfU
+2zGhr3rw/YUomeNdOWMu7TBvovQwU6jCMlz4+beofnwgTNZbOszn0x2YJr0
iEZzpoAbohNTiQ1noh3rZrjmkK3yJxeevQ8X02Yjgv2D0mBOUcHQ/xqL76NT
j7AdK8UU2vdFhUnOBGqqNaB5I/ozKufHniI6vRjUNZQAbVrmr88bbprstexc
kebiOfIvRoA6zh3NoJ8DmDnCZ4Hc7p3iGH1HmT+/DbIeEG8sUTxaV8hgZoOL
PxrquIles+Cp/FxTv1EfBdMjUSacJpAZu6dDAU28ys6rTfKLmgazjSZlSndq
0le/OsYsC3zKkpTTvSYnpCv6/uEQLCpJ1jJTMdq4MDAF0PJsk3H7hTVKuT/8
Ur6nn1YUHSwP/fE9XHBX5a9Cx/n6k1MF8as/JqLbN3nxEPs+JKwjOj0h5awd
c8I7nlxi4fky7Gn6lrZK8f7iLonApuqmAR9cAQzwQK/ITJB/+ZNzuX4APgDx
Lp0EbJm6R3j9nwgHSQND5YZD6ZSUDv6vjSpTGJ83NSR6svTrvO5zdIJusUO7
0aK3BAHPmEIHoDll72luP66EC3ygntS4jaKXyDK1MuJb+YdDT/9soNiSMe5p
0a4fuXxNbp/3E+aq7MsDdK+swyPYlQJ2uMUABS50fnhCQvPlidX1zGqmVubg
jm6sBzo76wSRAhL2yhZFYPSaSHhwNTOHZeDJUe4i28jG1C6O3qavOx18LpEP
vj18xjtJe+f9uvBb1fCO8RNlc7SAQbV4C+Fbe1dBRp6UNJTnycl8NXX1hBKg
kiAJsWNkcl44DeZxecBALNeib52fivjPv3Ke5insoinxYbPsLxodiSxcwO1h
KwRwmU6LqdIOW2rnoZDAUbLDOlF4GCA+oFL5Mq5IfpwrK6OHihB+5RgPFNfI
M1EoVv/mkANwRM3WyEbcQ2PoRZ958Ce6t7Nsg9UQxjZc7/HIjzHZGtlfr4BR
rqY8KrQJ9hSExW4aRtFVDWzD+59fgPFbccl84h0qgLtuzOndfnN2+OIXXqE+
sn6eJQoHwzD2hnC0CSvsXvcg9b6XoNhMTqWUDCuVtE1E6hG9DAmR+eaPvKTv
ca0hqkt5Pqo7cAQ4wU8xN9y7brXar53tajyZQ2zsfK+jDVzZePMr1G/MqQh0
mJha7ZjQWtxgpjruXRfOppvicBuCz2JOVnQKBC3w0bWJ5hU6I4SQ8KlvpZyM
AGLZh+cVXHWK0iNQHVXB3Uk5mxDu/fxecw8PZ1z0x4+HVoVCYqkJEhUFFtvN
2oX3lDUma0sRN7MFJgvN9Otjg0zMcEJhcsPy3L+0hpBszc28Ss5/xzQpK9ZG
tFQBMro0aQJ83d3j+kWI4ijScgb75GXmOAtw14EFB2NdAD6o8Uq+rLXjw9BQ
Pqhx5dLPS0u0ao/f52w6uz8vn8V/u07qfrE3lJTTXdEts7SNdF5qujhBHy9K
zBPmF2QkGkoXb+zFUFhL7nw97nTwd2J+zPtByCzLJCJ13P1LrIsY1VvOPl2S
mYR8MabC3Kv9RUy9+wpqcHYBxLM8NvdWqJUa0btIu6STOpfWB9WAHqveLL+V
NrRhkrGW0sq2QEg+UdogsTXtgUdLr0OghUi6vqBoJLgAG+hq22oh4VubbJnc
1gxKckOkuU1hdlkaEXiCP3Ey0OKDbW0igE79z6XLLdYVH3Cu/iti4oUf0ke0
ke8+D4a463hzNLOk63AI5yOG8Tt51BMITM2t2br56GpFGwpf5hr3wG4FOS0x
IZwCMNHunW1vmZKHfOJhZsj3l1P9d2XsAcVbxdPFMHqYDyQM/kE7bgzrtB6s
/mnUujXju8+WONidAKolqk3qCIzJwADtMV76QspCrnjbGuFMfpWXRfC0gW9Z
cEOuC6fKYlwQNYe0hd7w/Qj56ph8nsGN6oK5x/Z/sUpLoOuS1FZHUG2fA6jF
RoTCbi6uc6zg9au1P5opC/lwaPdaC/xICRvUroswHdGFIWRvLqLcYqARTD0o
CDkRtqsomZNg+pCzVI4FWlg701Q8x1p0vUIZ6wQjGJuHXOBttPl5uVNq00JQ
uZtXHwLUnQW9dHZLk4UPg2voG8HvVv8l3QfQZXlr5u0sws2gwnRWu+FBBQqv
bZV7pAv75LsgUqWxITE48ZIwZaelK1vGlrgCn9+DDLZQ9tTxo0CaeoSNZNi2
kL4/RgvTzrbhkUwyC9aQAHCVvgR1/7k18Qrr8HjMQ+eQY2dP/vTqcA2BLnRM
vbQNFDlHRef3I+5YfTYVdc/g9ulAk0mTK2cMZQdSTHIIBcPIfJuhh2FyNAcD
+ZerUsVkVK309IPXA2CtKnpnwXrAFDa6mwADtoxNoW8KJzt/3xkLtm+oRLGl
YhSe5uVWchn72HXeATaqs5AN0N8fCIfR6R11p4HPAXQEQo0+mKxiFb7hIPvD
CkLTfAaYPG7Hr8knN2XhazJ++dp5rRkHsdJlKvy+oXN3gnmtad7l9d+/Rdg/
7vfjovP92ZljCY9DDKVBasfgBbJLxdLMGOHa24UyS/i8/e14Hzl/PLs7TUOU
zG+MuALoGd2UMkijWdrrN4X0uDgU+BffX5y5w0RjCH0HVnAVVs9nu5EjaDO6
oJABRPpW2LZPa2niYXkAiYI+7lusryQn35rWo2frHeE8hjFMaL9qW94CFqrz
+NntXASP1xF7M/PqsyelFE/IXaHEyqPm6LzSS9T4R56cdIirzE7a4lEaSz5x
WXWVZE/T7/3Hb4zi4AbjdtmSqpQqJPPad8ch7/2Dhr9VGCArFG5t7f+w02ZH
w9JyE581Yn5vN8d6nbEw/IJoA6SR9nWIfdFjOhj8Fd6leMpCS/e1KC+CiikD
jQ8GCt3EuvcLrGOdtxLyUNMNt/CiHos0debmXTWC4kLjL8ifNQOYrAUNYBcD
qLWceYhn2WzGW3j1reG3AS9SkQutLj2SY2MCUqmM7Hb0LOR5ueWYxHT0wQAq
X83a5Myv73ddQ0TZg4UvkUoJxxY2xV1OPI1JTE528k6su4TIuVFot5I/VDFL
Gl4Mx86vGQ+XuSpFyMmP5MRAceVbE87C1koPKcceTOQaLcwH8gmZoueWqQu9
FDDqOnuArEeJUsVVe8tCCyicaMxhQ7NLIyfc6nRE7lz7+hdbcq6MvCJgrit9
YcOf/RUNivhd1YjtMF2XrllT/Qpirb9ktAIXEQIfclNbhAc2fmBdv8lMx79j
cou0oFGev3332JAjx/bRc5IlQIJ1esA46pTlUfAYhlQ4GYltpSYse03Hjyzc
0jk8p3P9Lt2Yrc2IT2sJrKHu8Db9Ys7+eVjxN8vtuj31ymbxgyBqUShEY+fQ
8R4uYxIN42RTKV4STj1/wlrWLQq2HPkUMlbfKEchojHdWRWZFEJeAZcejYAw
e8ITazNOO78NfRldX0ZIzxpRMFLWwrSftz8DKfa8FQuAlkyW0nNuoGsLgWCv
EtXs46Tm4v/4i5HypTfA8jHh3GLHp+E3QiUogkqNR/G0aWzcXqHEQtoGBFuo
6gR6qcXGKlavW/d4WzLgTRqM5BzULagIgutxSkySCXbzWTjtUaZPzruU4ojZ
fLqMOjhwLPRCcBkNkeLaGXIYahSOhEBixLtoNSTRvS/v4QwryXnmclMz+S9S
OAs/cBUPb9MwgTJvR+1zhJh0IjZXXlpGZN0iyjLMcmJzr9iMPkZP7x4GaSJm
QzOISeYsmJmH1aicPKX7TngDfBzep+cbxH96s2dFwWAj16Frjp0MtV2akfz7
amfr2DBtNb4SQjKD+vcA0fiOWmKq9ohUy53ET5XePNbJ7L95b6a650CpNtoR
p3Asbav3ixo9OTSWiEwJNnkN5xNWINtoARzSv1g72p2RLIWvpMWYkQTdQ2M1
HeMt3lnSL+kp7K0n7SSAPVe5tisVPMok1+DZCFPaDZBmF76KbZAjUhzb6RXZ
rzLAywayars01c5RwEm9vPap5ItYBUKESuIuMsteZziQKst49u6OWLZxz4k2
BQip47rnowvoL0ZhHbNMIhuE3uW9qctI978AoIro+b0LXBD4a1Kt2fY5SVv/
KXdpXn2R1kjQ9Ly1UdqcaxU31BvD8NromicMwQic4KnsbeEGg9X5tMSavA2g
WWMZ3euIVrmXj09I2EywErFzF42OCVCmsv4d/gh4kQW+6g6lCP9rtXK2vmq/
aDMqMGsOzwYbnTJSCeC8jcEti+59NQFv2PIcaikcxpvbG1KWhE1GU7HIrbXq
e/CwWT1u+XQPlI40i8nMfA2NDGfBjzSwV+7E1vbTkTuxRJYfz62FCscdnsKU
1Awoi6ZOp4iP9g9I7+mLf35449nx8+JU8A5hwOKhhE14+t+ePtdvZmBiXctX
Kvt9I6H/rA1ZLZmTupzuzhXEWX6Lz0jj3FtNXs5+ay5F3WXorqXf0xTKj6RK
YPMmmJ9P3O32J5p0+8beE0CIxGfWfqpGk4vjMjjNDu5y0q3J5uLqG3Hj3TBF
xk/WRul/EqSNBv8x77qxgphAr8E40hpkrMY9XGLSAQBT42CCN5YqVuXO2X8/
Z8npOyIQMrYoJK8wNz5XnJDKGh+EExHiELw33IjkZOTeC/uiFTMmwGOaEf5r
ycMlssgsGISKWO81GnynRmluOyXXHXSkOEDEaD3bd/1KTgTxJWsP6A+EfZKL
4bqECo8z+z8rOH+SkMgzRhQO8Xvz7xbIZL7/GSpjRJQdUjby02MvUEZSodVo
oCvtb/WtKRqhfECeGID1dP4TfXG+/4UehnZ67WPR2vnsUc17CtI5kyJZuQeh
EK8CTcCmOtWS99hNBe8jIGxKVu7ertM7D9J/uSkmS60QZoCNiZxm5LeZ1GUl
+UIVibVCKrq6YTqpk8LpE6Z0GNoeaRUu/RWtCDYWR58qwCKFEVhBinJWhHlf
txAtI2g5EP5RTrZRkw0XxcoGjUxCq7Soni8YFLjwZ98+oXF5zmcF7mGqhKPx
Qposs6RDNQyB119BfZGNpEt+Ib0W0h/iDNg72bgmk+G3XfZs6fz6a0jk8ORI
TD5mdiVLYUvz71xJBPCevBCb3HKPMmwhGalvfdZ2mimlkHG9eUSDNuXip/yH
nMkjuIIibdCLTtC8mVABN+6p8m1n5jXcUA9iBa5AF8nJl7ZrawwoGOID03EH
pnC+cGrZq+iMtI2T9HB8ZJdD1YQVtX45+CogDfL2DmHqnZIeebErEAG//eHF
ZcoZR02tlFlBctWMib+iHAS1pkHVFr/I6vwfjhMENWrnEDwPAC8VkCUqcuNT
jbuHQhgYSVw8wgjGVsPkTvFZvtCd9TU9Avj90GcA5m6JfQhPxy2Mj8hKo7fr
2f19mX8tpM+6HFOOHlEwNDgAQTW+ZJ1IZyaKgAb/OPVVEuBWgpmRo2fcTtoL
CSvrXfWFV6btp1oFL69ztt0/rOoabjJE7szS5uzNg7iLW7bncw1OzcV/SLQX
VMbdhCO9GGNK1WS5fQPNXeEkWMqiK21KDz3XiGoMCQsNnb20ZPcF+Fe7Ji3S
1BdVe9kx/to7wCvuzCkRjuk8nrvPWBhFTbmEIi/kvQdjhkipp0pk2Wow/nlH
XKa48irszsdcH7BA7mOo7owlo6O0wR9qu1/OjkuJrmDqb1wCtrHD2K6RnKaI
0HX/DWXL+ZIEB9bYifHbKuZiYvPWY06ZTR5ljv7Khi21TjSE8Fs6lyNTVthr
Ugt6oOmY+rE5RdYvuPzHB3Jlk/R6wt/6/GipwyGRhpGV8yzx+AOS75bGIoBa
u6dfd6APVRjOdPztWHi6W3ZQ/LBoReVOgOTgIRlED5m6Fd/9oVzokVwA7vq6
DcgdB2kzYKV0Fv7AU9kAMh2w55tCcF1t+KT9p5Nymh3VAY1Q+t/GyUI+Dpoz
raqXprZ5JANnH2gsWnW1dUX5Q3TksLg9VN0FRRc5226aqhTJ5XLPQ5uqNBrz
baOki5reTKvRNr8iOKzV+C+bVIPldtqNw1w4RAmW3lsPcvlaxtLAgQh03kSK
NAY6WAWPhpOoAKiGFWCMy/6oJVLj8ZTlJcZxnp+jNGYUeuyBg2IYq/VxXXxl
yhXRkfIR/uxBW6UImjTy4nUb3ppYReJDZpd3fQ8VqfMQ9U1aYMt+Rtq7S7ap
kr50HqTyJBVwsafeMtx5oXcnfy/Nc+jfjVDf8K0RklVM3oNa+KaGSj0g69sx
whepyx0Vf49Nfws6tzpYQnH5pCfFDM9BzqxLqlbhqK8HN2mHUWcAscquWi5x
IB2LBK0iOjPqawZgs9BDfibsCyM+R+N4QbP4mikL9gs8WBR65+qoXHf86IJo
SbYkVgtOiwxEUeXxtWdeeVqfF9mabH7vJtjWh4H014V8uk2mPMrLtph0B4h+
oKK3vYy7clK01shXJ3E7439wM6nuO0KjIHRxAURzGDZk/bQpbb06ddh0dyzU
jqZZNJXDnpvLNxqU9g7qs7r7eB2WeEFQO20K6x75oOXx0fDMYNtWK8GSWl6R
rvQ6xsjtL32RP8hdSYq/vomU4Nz0VBYuQSiJHELICaa8wUoVnuCTzC8wg54l
Y1urpG65FAfpC9bW3nKmiP+31GwT9CMGStV3dH0aTm1rb1Q7S72WetJUjPq4
fHhjzwro5fRbLpBDVLzugzsgolYZo6OkDZPiCUqkZireU8jGfBsIcx5gGa3u
h9yPxauGfOGaxXGKz2jzVRp5HTMJBpJ9Lr+bY8ftJnkOrKEUZWOT0Dj+vBse
qsjpEjKUHL362vclgKYcYfdZ3+LDwF+duUwbUfmqDG4BtFcvkk4Kt9q4yku/
BdS3/r3PPHQUAd+9PWRY6onwM+obqwxccLnQTMgUdPLuB1EVjMoTT+sd5mw9
wRIb4Mw8Ny1DdRl+B1kg64o7VqGGWTT6tKkwEIT0jc7opMwoMpZGDlcgWoP6
xrDK1om39gJ8Mwww6vG/NFnSG5MUmJBcKlq8g5YmafNHhCU0Ne0z7A6PxFub
VBtbrWlCPZUWJ8sYZTGE+b63ooNt7Sb43D7LSs1l8OuBU0NkxnCpk8bF8/Zc
hVPtv4tGbiSiA3JQ/D+/VsfKcmd8Y53BYBTpYNcQI7Oe7yyKif7r9sErjQ3N
lh7boH1pEbNJTirIxlcXnxHCc+gqZAOPqp75kMpJ1nYmYMbQd1UL3IXy5EMa
OouAFQZCWAcViT/7pPNtRrK2qJIQFY/eTFoj+hNA0ggEdNfwWEHgbwK3MS5d
01rm1RekTOD4Fbk4otI6AmegI0xNJJeUUR8yp8hisAP/oDAyxeuhSO2TvUwS
XCa10Qs21tuvwDEQz132/xcMjBUNqHdFj8C+Xpfdk+6OV5FPf5Hr2WlhGyC8
MlCB4KsDpVZl+KNduQf2UK/S6V/3+Bag/pCZkoqXrZandIJ4C90wXJkK+319
d2a1jRyRPzyrR339uUdsvguJyzth3nZEGV6FRoyJ5kpEB8FS+qrt2vo0edmL
PsEMihSv4xqkdxJ1PNrmYIS/6jJjBM4vSuk5oFeJf2df7JMYHmAVYJS3gJK2
a8EAvV3GYL2cSz13XnBkzk8GqAXajwq+ZolidvzzkMCf/MLKdgT6oaeY6w9Q
sxYlhjaOaG14jZjk3M/loplsP+A9z4tos3hKV9yMTIfsf8VZxgr//gNOJnKV
ZyPdkLDi96+60L8cnQK6XSuWvQLPtGiI2C0eXxkqCwH2/loIKbuW0U++g/GW
Mu9WzuJcka44YyXS5laouiH8J3+sc9ab7aRIHCymbYaAKezulrf+6UYWhj1j
MNI/tzaiV1vP3qNLOZ/2FhexygM3CBFg+tiC8nG7PNGIZBtgaTY8riiBXVh+
LASZjGZCL+lES6188qW/ytoy1GeTBM2UYLK0f7zf+MXF2AGw+WGOGgqatQwZ
pdkDp7DQXHAQx5BVmbBJOBInh3iiuUoCQWb/AphnPBMgBhRaMVNF2wPzFnsr
gSxzP/IjCrkTFTzr8BHJfthM3/pHbFEUfLT/umVmrfHzsB22xZqtZdCp8fjo
S+Sn6Olux6yRJFGLJkM9Ej8Lx2EuxqS7lOvtqWBLBNKeOZMo6FHovjpsNnut
kiWGB2F6KRzabGyUvz4S8WKfJlLjvZFghMai1ktoVYEL3rl2LA3rjD/ZaCQl
ed/8YgkjHixjgCmm580hGS13Qzq57OfiMlTX4wTrXbSaCEbgiekNGrZVb3pE
OkEf2jde8FLxP2S/9mX9KehZBT5VL8fStB5AYPDnsX64BjdfUdImgykuTvWK
1+arChul1OlSmxYLc6U/d4yFmQ1J0nXUnSX4P+VZgdvWqCCxvN6y7JFn8IV7
ssHLtQTnm2Hz0v0WbIG/odjW0ZTyWrZ035CC69lZaJLtN3qsAHS+eolPCnOk
pSkAedUtorxHSONgOzC9NZsoRqtnOdjlfyorouq/LJ8/V2KmF3iEc9l7Q75x
qGek7LHbuAhjSiFNkuZA+Lv6pnenDnjARA0vikvgSELAWJF2wp56cBlRyjrp
z7WCuUZPGE4xCXmXmJkjS5e2KCRDYTAUyZSaXmYVK8J20hRxNA3qIonLwJGv
4vzc+e8D81mpj34wMUb9BTZuzmsLEzPbTS1CsepU517WnwkQDmxPeX5KBMYB
CNTTvdQeJC8C9HtECM6Emf/0CvtgDFd5dwv9HMm4QSD0xlnu4ceqLzzDrTJT
zcrljGx90ecTlPqyKJPrIotLtoYnqIRvAkWVdGqPbnF3NcXhv+6mz6cnTxOs
VthG+hn79eQFDLKLc+/PkUevnnIT1DXDdFvFsWqy8UV8vTNAKQKmNZTEbncb
HpzsYJgqH/e/v5uCWCC9fneJ/8jNBZSxZYiTsRolFsiFHin4bnzoTXhkuLnB
WDbuA13VQne00dSXa83DcjuxhZTSMmWcTj04v5h3D3BygMP8BzCoW9Ikd4FC
BZRbenl6kahnyd3v4I0PiBk16ryE2Q4ORoiOw8zcVhNd64m9orisINC7Z3r9
Xzdbj6rCU/Th1Ktk5eUdFVC+AEFFVmEgsplYhIGd82y4VeMW+c4om7ElSKfV
MCdS5AwXRVL6IeNHn9pmdrteJBSM1Cb02bjnfO9lyKF+EcAtuMnSpsuxlVZf
h7Qvo6mZ9kg9L+A6sJJElUeNRT8aKrraOZb4Ik2ztO01t99EmzM0xlg0psYD
GtakKFEwOYbaMTnssZVQbNLQFgAETJr2BCxyucek2zKmRda/GNWO0dYVzSPk
4VyzAHxqqLenJDxD7EBuUYVfsyTLfoDw4xQ4aAtKs2vHIYfHbp/JUdOk7+78
AdoDyxJtYPHwKGfIG18kRWae5ooBQSUzogtV3Pze8SFVMfqWeXTHs8nzoPzH
bdbho5QYl+bcPV6ysQGYhgklKK9mSE5vi/ANvmQg+ibpT4YItaWJjpvHkOza
F+2VTakgZrFg4CqyHzcYkkSdGGFBk+sxK8G6zbBOY7SqMom+3xiSkooRIZ9j
CxLEckPl0EPNJEus/voNxZ1ZNZz0z6TtOvX/Me4JPdZx/lN+xJdUiYoBu/wl
5hlp22B97hAKmdaFlM1cEEUuQ/KdRztL2N0T2UrGNLWz8clTCtz5DkNTRDSq
+hOtYvuH4k/ZVIvIc6ssoxEL3eEGEeAdiBNdYm3vSl6p4BPJfjuw7ct0dId0
rwryHazJvoHbYb733GBzdo8Cd+vLi5EQQKnUMSDZly0iZd8cjoz1hBMvrpMs
4wFppOhnuISXFHD9TygAEbsAvUuBGtBk7a3CfDl3RBdUbVqwsILLiMHbq6RN
tTUJ+d4FQgI8T9/pbC5L1Pst6BB46GCiyfjRqQG/7BoYUhimuGa8Foru67+2
c6yyZaRZdTOIDvsGcfl/D6GmrCDmVEseP6aMOJHts55ImG/M83p2lwE5DwbU
zs9YvUEmfY3wfnGubTT2KIU4PwZpecO4d2oEh9uStniBbYtIhCVmYmLU7t2b
gBdJ31V/6YCOXhzqy4k0idQaacQkIGspR5L1SxqAIUz5YNH98CFS64WA4UDy
dAssc027+gUhsI0cvJKvpeDhVr5rp816UUWaSFEaRQLiqpvcMRRWMaJmY73H
xyKPv5fzz/jwp0CvcnlgU7NvXCM11Bpx2UG8wHo4iWIgzmthPgfmJ4od5arI
Um5WSH5u/vfarCRc/dshyOcK4cbo2cTQYgEYCYCH76w2GXYIY8vZA3H+sc2J
Al0qd2I9Gq1P7PLtYSrWwfmx4cQyZgiWm7WHzFSj8FcmKdOaCn9Bf5nYffcf
e57bosizGiyY6aZynxkQOAdTRgGl0gXVwINu7MBMCr2eB84h/u6zvuX4RPFt
rml8YsSUl/Nw1OBY+qsoNQmQLO5LFIxjetVosmfKEUAUDcn6a9Icig2nGJxZ
P5nD/R59tfD65gh+0Y4CaC+/XkrOUxEp6WIxVapF/XJqKt1YlWApM5X37TFp
RHlhm+yofXOnF+RMgjX4CuBfXeVrcHxI+354PUcTre37VqVbuaccxGsA4HpY
fzMhfmUDKKF6DEu0rorUFdUVe56/WT9psWJZhv47yM4UN85E845ORYhFmV9A
fh6jQqrtrSlhrBtlyeJzbT10cxY9BbpWBH6n8LN4HRJyhSNgbRXKy2L7Qx/P
tjPa8htsLFzOTW+G9qEnZTwDVNpBXueiZgz602hjN4FvPH4Fb8QRBz7Qmsow
Nk12qMx+tmtWIhIOVoonvjhQt7Y1LcWYdwHse/dqnOuwyx0rBL2jXGVbCuW3
pPGvEJGNd33BDZhYNkHvk79rQKA41YRh51/PeYNz6LUPHgH4hUk1aoVp3A6m
nfyjuTqAy0REuc8QnzGDYW3fxVq51bOiBgEwpdJXW19b55AmJq3pHMRmpx3+
R8Y2EpHymNRCYL2nqW5WUmNDbJjptxLgS+KAaOQpkXuatN5OTQzqIKlppPJq
/1eELdDo775qCNx7gW78wO5UsBeoXXUiHB1Y7jFmUaFmMe/JGQInRHh5yOme
MT/1QBUgoUv5JlsO4gZ5q9OOhXfEO+bQ2UNHbqL8qwN4EvwxpNX0p2I7ZYr6
5k72Oo9Cc/LMBhQPdRX/9fd6HlNx4ffAE4HTI/Chocw5cg6KecFXeO1UOcQo
hFYwQIxzriseQwfglYHCRMEZfp6MbSY6oqfgiZaR6P4baOceVvdnL7wKbv81
gS+apMDUnLMad9ZD9D3+wAwAOrEKAaBJZ4JcL4Pxla+uCCZOHWUR4+Nny0VQ
39f/IhHAOQ4Knih9v12aS6QbPJL0wDG8U8VjRLKSEw6VS0yzWa5V4QRRPWHQ
BZGY+91nbli1qowlTVYPMxFXo2enbHpMXysYA4RXYuxiP0ReJMwte1OPJtv0
NiAKwhnLsktav5xZupNtoDGbtmukLbPgYQA/dtbkVzGDYRq/U7txU4pzb3F+
nbmv7a9LNfWDa+ymVOVIs5mi63/xlSvkvWQeMQ7tMj4nPsXmaJflm5PFjbTF
OT+4Af/DiI8P0wWjAJxRAGD/FvlBKNJzSfC3HYGGHVTFLUQRbcPDbpctRk/P
DYPMALvACo5/o0w6SG5vB3IAHlKT7daLFHQzLk0xaO5RxRKk4iPaJUfRQV9c
b5hNUYs1g/jhPCDUgjB5n8Ngoe7mBNMneoJPCgwS8kf9n4IrK9RoV4vrMxNC
2m3zvAtiz0CY060GM9P0vLqLYFx6s8GFM9natglEsnLyj2Soty5VfU7F4Xyo
B/c8gajVc7LzCOcoWi7Td81FsUPnZk9CUL9f+uKQ3UexES7zQ6a1nBKLFXzo
iZNfsSMGn95jji6e4gne1fNjrLochufVWtvZ4+mj+4GwWzdFDS2VY7u5bXTs
Bs5R5BJpLpqpge+qNr3e0Gp0W07m8c5jMjPbWzWLFM6rCM2ZTtSE0JZ37HtP
NrNpfA/NqZHi5kLbOIpmEXQdTZbM2Mk3ZxWPYQJQPvs9m8byVggmjjogqZux
/WKRGWPKWCywwjLSqyK9+79NI0+rp9n+w4mt9NqGfN29SX/LOyzQhHk0Rc+h
Z8OGzbh7LgRSibXgMkquw+kk5UOVgACxekmXdEbCL8nLxM7S+a4YmfgcSvtd
35y3Jpqg4V5soTw/GcaPLILu1WbbhwZzlthoYhSsPzSi8mBilPdgkto5lJeb
fYFQZecVuzAMHpceiGdDyJk3l9OS/sSp2TdBh2Y6WiZ8Gj9fj8QssovbX17E
zXsLqw5m9sBXOKAPX1nrkrIEz9f0da2tUiDR823yuTk7hjJyZIc8c3ug8TA+
/lLPilTapZXIV/nOOKVBEj1CH+2ws3md+ZUWD2UVgL848pOcgUTgXdc94s/Z
aeWJ1nrmTVB1pIUbXEbuffk/9zJ5cgQ6g1ILcSZHMkuSpXpn9HMKrSXOmRTx
JRn08tAtXWe6W11pTWchPYD/OI1+aObeJzTafY6nDql1+MfU387hMBP4Ew3/
ySTDrOvrDHMQJ/+TLlVi3hrDXuwyyeoDDfUKqDgjxJb34Cdjv9ycxKeI4Owc
1962QcvAwO8tYSV1U63KYYJ7jr5YS5gOm7vlOd9cd9VNLNWU8QvgSmWe8oye
+Mg35F8BSnuOlaws4R1AjpfCUd7uSagEs/Br+Njw450EXHHhT5GJNWfN9vEF
8aetJYRek3/B6xIh159cn+s2snpFRutXLIWE+PoYeAfDMcVIFY25BFXmQWxj
MtnlhSaUY3Jki0L+t/YGPHlsvWqFw+HVksL2okcEphoRhmHQ1v7BU5XM6OnZ
Q87pdRUWdGsJqzRk02jGI1vA9UYckTlOurIUQ9byGdcMtdHd1EWNACfcYpWB
1f3+6z14NwZUDKFqfF3SZjH/Qyfnmr3rIBgO/nIKgdE+Uc6rWSug1ftZgxlF
Z3ur5wnbHh9ay/ikUz0z4TwvJiYUhknCoDbSfQ4a8CQZDpBLcowT03vUFV3d
UHfhbY21MdXNm0e/PAXkR+vEgu8QiBasBx2lrxAVZBF+TDpJ7lzXUeTyJk2i
05uagRphirVtR78Do5UV+jCTllUochDa8VWf55P2CiuJFZcWnFGVsZXe3UG6
iI6aCUoVEyffDOMMANYZQ156xfih8OllBDxgCzO6Cs6goCiVCxuYr/l3BCol
gIpq70JyXcYbVyjBMXvMSWDeq4v49NQLLCg7B2bFEeLReuBBGNE9HlfnapzM
0+z3s6O1XrAH4RHOD6NuZH38n8L3k4swRUQimH9u2+1TiLbfzs5Yu0xbIaiL
Fm7rGRcMZN7Bx3+r5kdoQJLq0ERlXRdW7l3j1y01hAWRFDTUxJWKgRE2LQIR
DbA6hlF6nMTDvEUf1FOoNY9tBcIggFViFVcNv7D/EDZsnbhz/2MY883mPI/v
Buzr7xzlTp3gRsDDIqtQ2EiD3G38Qf8Vy8c4wT1tbeWfY4bUDqPa8s3LL6+s
d2MrYnSG7sVhodiaxk8eI7L+J7y8qG3wkltIosGWI4X/4QM7BE4ljp0kWH/E
AWSiubrr3FSagA0ctue/J3yECrZdPKR4EPsTq9kMROfvaJmXhB6DzKvKL0wz
RQYWNMNDz0lW4TOXnrpVGZC6hPB0og10ll/ykO510Wur6/8Jlu7HLqDmMXDk
VedyRqDC7r6jPmRvQQxYN7OLifP+sn/+8LiDDLxEG6jzQeMAKHSXf2LPlGNQ
g1J+JdPGJSpX4P5mW5u1IBbjVVYX88U7jWnCsnT3md0cdQW1Y+vI/L1fCHoo
D6L3ihgu149pSFsuiiaAZjFSC6YI6NbGXkcnW0x+wQhXgAPf0y44U9NVdyyS
PPJdkjOz1TY+NxppK+7KAC5PrLJF2SZ0H4CchRgbcywP57wD/PRQYN8UYWGm
kbl99IAii7w5MrmlULA0SVp3rK6GE/53qQ2mGfkIseuhLdJ6UgtFAMcDx53b
9ZBRWzA7GLDwlyGEeyRAUHw3aQOtH9ASpHZ1C/VENdnP4iX07TRNexvbajLy
7+PCuVaFBD7Tw94mefYEDFqq+pZbsaww54zU/6nu3Yu9n27Fb0h1K5IUJmgK
VQV16FdxK7GKzzQTFVhKpmQXXQp6eWwEr+edVLaYq9396zVIvVEW23bei95B
s8VMOvdhNRMG/DCPo8EbiN6Og+TxAsOxyMhXlS26eBer1vJ87W8nstXtwDKB
yeP1/N+r0gN/fqKkNvte5GwJ959UytIZQLbeTgZj7YhdNX4yXYeb1zrvxM8L
7AK/R18/6HfpZmGmlwzhCU+xm3ku/bvqotZjVrgoKDh9BAxss6KLMg8uH+9e
mlYr3c6exCcYCFveRtBtNXswUPe623WxKh36WnaN9GC1/jAyxjN+rDKrenMe
8ZU/FDyDKsbe/f8bmWEwo0CghraGQbzHJ4A8cFGImpY1qiDFR1Acm3MXr8Oj
/USJJUK3MK2XgNpAhXlVvt24OufF+O8VoKlIZO0awp98pg7uycENXh0/OuGe
+68Ej9/VxBGrwmndcLrrR5E6cWALV4JgsQvkQS9U54x9kuc7n4TU5FDZji+v
UWXYAz9WFzgxGFCwUa3bZx0HLQhFyAeOhEJ/rihgJosjZbFnkR0yrxC6Fjco
b1s+i64Ao932YS3TejYyoT5z428B0RjwaCH0383KeDcZ9QjWslOQioBXjMKh
S3Hw01gsHJbjCD3LptkNgasfJMgxlvBQHepxrcrJaOQBuaIo+LBJTx8lowCK
f7/vpREFdAX+JKzrGdY5qjGd1XCZOVciGt/rnxiRCrbyhxmfMV9/hB8/Uxaw
CghHlxDmg/spypKHu7INYNmZ75091OoGRIC0cBeca+GZ5nE/XGfxiN4Evc8K
0L4e3L0WXaf2FD4vGHXFdVLx2YXCxepN4y62LC2171wkWNw5x3HtmVmQgHrx
Odw7vNW17dr9/Ftyl9vz/PliJRWUWIxQ8vp23pPatFR9n2fpne0VUuASu2f1
jBk/bLbKalWsY43hk52cHmodkheuxZmwZln6fBkbW7Ib8Y5s9DJYk0QVC+ZM
XaRFYJhBQtedlbh7T1BXbdn+ZJ1ZE7wSuxlAQPhIDnDThrJrG9BVVyHxnfxE
wyLFFzJW/zKTekk9DWJP3y/fxMCyxwGg/ssNsjD78Pbwzv/dF25qsohsoqPd
AZFiA5v/pf74cN/z5Sq5egZfjWCA1+IqiJ+Fgl1cLNcyq3rlBxWuW+Y5ks1H
kPq50PZyJAT6bWS3sCHknGtKg81Fck/2PWqWNAJqMAERlBExxbwNmBuKUKFp
xW63vIlZYcIHHfGBLUDEcW7U/M7AbBd9j5QyDwpc2Rt6U4aETRtjywST4Kwu
3vAYQARN0jFqO05vG1fGJQbvoY6hfdn8n5lkBMkwLIgFqnYT7zGigi1vz07Q
CxNfvP5KWpg2pSSLLD3CNib/lT8hnDM/JvxalOAySxTUXl4p3ofNKP3GaIdw
eufqp3vKnUZk/7RLxdpdMKtBV9/At1B1ew3KfVDpdRCH085vszdneDVwLPFd
WLOM6vfjbv/Ofoc+sh0qmILC27QaBm4za8oaTKjYCKo7CGfRc35SVW02zcIO
6yBQF4Uouc5g9wkRs7piPD250rpV2/PTsqB3/LXidT9oP0fioWJfT0d6Znkz
nEer72IMZwC/49m24a8DEc1Dx+2Zdy3JJdTv7qyMguGZZc8ljqKDlYUvkZF5
QFES0xLc6LfwRsMtTxhK81lsJzkyaX79A0Owawg9Xe4M9yP4MPg2CyQ0ktWJ
JH/iZfHQZx2WI6epY39NSlnMNpqILTK+H8NfFPnDocGK552+U6w/WiLUh3+Z
0ccSW3mdzNFCkGn98YVk0hnBIYrmoHOIGWpIhWQKdZeX2y33KwSKAIkT/AAN
Y5lHecEietJ6sPFACYX9x1ZTEEtfJbAd5NpEZPi+V4ozgPAOEi8778BuI760
mAGwOvRSv2znCvD+6ntk0IqsBEFnnyV6NdAgnphsx004rlsract6gxXRAdVG
jFoHUUFXPvuqTGH7dWrSlwkX99fc3R6XvoY/XRfLpGFqVF5b24nJin8GUPdD
JE0skP06Y/g+Acv3VpbF4ZazX8Bu8kgS5HeAJ2vYmSp4J//+mmZJrTMR+/Da
kuTww3+4Xg6ZOKxUBxltRn/GtXZjq0vsSNQ9ITKT2khffPZfWc/6B9V8ygBc
V22gHCLsBQfUBWSyGkF53zf4iJD3qLNYvfx62a2TesN97EPtEBTn7BMsV7nY
EPFiLBWPEH/8lD6f7hm/EhQkXqAmw1vAzWiz26wiJi0Y5sjUpE1LI2/qCYao
IeADsu/RCGa5NemjjlkQgWiFUK2EnxwhmufEjqY5uCHMx0H91H1clsACxber
6avQSyj5SGWBrLJ8GcsFR/MYpoEy6iLBFKVu2NsTMvG4xSncxYK04ppEbojZ
O2jhpoQH1OgFCXFR3+PllhYEWLVCBL49vE4vrxmAbwIjkntnLz2pil9Ak3Zm
wb4qxt0sn8dPKP2zM7N3t4JZ+RyXnKQL83T1IpG0xxUFprgiYcbP1hcytQL+
6lXFIpyVHeC1Wbg3fJQi+BrPDarOioq068t1+cMVw6zSsG1KteKOvqwxZIS+
w8kQKB/g5Rl0ytrIri7Y/9QAlXzEma7BejNmpA0N/8AIRX+QiDIMev3V4zWb
xTe9OKVyX+qjWtCD6IVtav5MpWt2CsEEADFa0G0ajC9f3oTcs7a84BBAG+Lp
Oo0YRtGBReGQI4hiWVFpjekqqfC85l0caj0Kgnse5nNMa1UJ62RHoDQhJSGj
6xvJS1rWbvkFGlKzUwfqAvyBjFL+ygvnGGLpMobbuA9Ts+7MiU/96xbiL5Th
jzs9DypUsifJ+57g22iutKfcWwBhUmZ6FjFZ0kH/x4gwYJx3ZEd6mWzdFbcj
YoqnJtUdWNRydp2Gq+lnhiTK9lr51ic8kBF5IsQ+1m03ka8utJQpUwWIvsE7
PbOSFwG3HdLeuAFfZEf+Cqx9fzVr0YTG4tYRrAqes/jXeRcfBZVTtiDJ1eTA
cyk44Yb0OFF9s+KSKTqjNLQD3cW0d0aPXKbNQwPFyDbQx9NYjtsg1F1/08h4
nO85J/mxTMWt1Ra83h8Kd69q5M4AJNy0zO0jE8S/XaoAVQi1K7JGuoAx4oh3
01scUvkUPFhZ8AjOscxnn1IVJX/XapqkORnOe9rZm95+0/CvB3A2NeCUkayX
5rI7hrOZ8S4QU00sWgiTHTZjQ1Ny11HiwdqBfuc9js1fyfUGODchQerHoLHD
pE7m18KzKTw/Dp3MdCU1cdSGmqIf7WwkjiER9zkVjZsn23Dhf0aVSXF9qxme
tNVhcCu2U3JPkybejrSBqazMoxqUpxIMYy8vFa/B9BY/abWMsNErm7i8Zlci
voTi9e0XVnklqVp+AA6JTja6LtsERSjgTqPgoqaz0R5Me8WXOaVmT2jqPV5v
aUs/gGSFO+NvqbnW5FJ0Q0rT77P+m8frHltYjHJenieh9+FRuLBnvOjluXBJ
LE4hPw+elLpdb1YCLBwfFYrS1inCtgfpbMVXf2kzccFPnhIhyuCCBorKSJOP
1LHEJBatwU7a0w2O8tCnBRlOGewA6z7dGjxvIt6dkVJpCiZPCOT4yIqWiEfo
Y5jPLizbxRRnaxXlPrP+LPhCcyPbQ5oL5RoN4aiPJ+eEMI0Lw0juu+7YMFWX
YgdAnPR8F17NzipFt7j+mDREwNpy5Fc1LJuXSR37UIkGoo4kQrOIU555ve6H
oHNYRe1V38ipnEkwZr+dSdz5dEbcnVGLgBWeSFMBK8D7bO2VKNspriaudo7R
ZN6oRJmcyDuVPb4g8/HfQlqdgPJzZIs5ewKZAHRqqNhuiUJ/OhCZ7BKvkwc+
0gihY4nNIKL9Dc9M0jLNv31uaGhqVhH355MxWVbA83etFTiXlJj149onDL1W
fE2W8++3GY3NuidHuuuslzfR6bbt7mRY9lwjWgji1gpXlxExI3e6nEKlihnk
VpyYHXD7fXv+R5N2hY/OyZ8U8SkXNdrjA7f69Mu0byddx8An8G7CsZX9DC76
YTh58pEGQ45EojhJl/LZY40L53r77NjeJDvVdWcMW6oGqO3/MRXB2U4cYIdc
J4PwphZ7Hba8E6m4At7PffFAwyLdTWnfdAjDCq27/ZBU9tBDGwdV7FQ7wxzS
jZz3+VTMkRot/y9+gsGdDKKpAVpCQ9hqK608VKdGHnVrPXyKEhnSOa78nkG+
8DLEyvJoJ2KzLr0jx5mvfRsEnNjZ6fOWT4IB3HVJ7HCoPHew8aZIvSHaQyD+
tQK3S323w8hhcbBDaLTIQ5ylPGWQo1tRL8nhPFkiuJHCgFR3xsSizjQ/mn4R
yiZs0M1lfetx807Y5vCTFib8uDjfJbhrcD76ouBlZYvbD5ADHF5NZ4sHyMyR
9bv5KpzUY17NK86Ti8hVy1DXs+tJY1Bfa+Ja7i14F08j87HE+V35NRNmy3nz
fG5uSYJnDtH0qPGVU1U2wkNgLyV89lljk8YMqIyrKliSjoYg+n5VupXWjx8f
q5wfghpbZAKWwA6wzxKfzodyxxDXFeK2WoVPFT44kdsqpYIufp3LZQDprS9T
vXnUoIdFD5mnWLhbBX/ntZU/Z72tPch1jygFwPPwU7NG9jKGo9yPbL3lQhJZ
ZMa6I8gBmlNMZHjQMDE17lRtn+LdkbZj/TN3KIySJploUJ1w01Aetx1dzBN1
F5zeqTpu0yXxcOs40HB+P+xJSSdoKDOAPvlKYp/6c/cb/VIaY0lHkqMdwF55
v/2Yh3GhVrLfUHrxPgB8CKPIeZ0IoGlzewi2c9+PfHgIEg6tqeJkeTrMmuzs
/rpsABsxjfdzxas8DrKQSnBKwUIMbQ8lX5hj98ScMuuEFzZeWdGeskudUghE
eu3Lkyms0rL5x7M/e3PUalACLpgYNvaktLoDFX2XP5TJCISMVpg8+Re1M9KI
I/zv0+jxLMJnCI6a7mKznQ2BR5thl09aji6k3Xu9SIgQLGO/gOJCqq60a/0C
8gQMaY5hifQ2b7ptqu6GKU2UmfxHHUFgSlEEFoHdBqMLiZrsFIIrHnVwV9TS
1J2oPt3G/UQQvwbvP3xTtu9jE2wfQjY3MTlnuKKiRxHtZ8AT883KiYYuG4/B
8mjlSnAI2qOENqeozQIJ8KnOJf8DY5NMTU5EFCZ7kwPyvNe9SyTmyVt65lsV
E9da6KPQtiI/rCzjwuUPyBmUQzLeIftncgw3In+dMUBWzZ1mjGG3HNOpT2q8
Q8SKZavA0e4E2tVBJCH1CSfktsi0bzdMbszgjEpArLOme3ZKM9GB33Gmhwqg
UeE/Qb+DHV70rI3s14ScA+PAN/0O8xFa1aHnaubQFNhQ1AdtXJx9PQ4iKaHn
9Wmc7pEsuombUPIHlUe5fX4n/g86rsR1sWXMaVLNn/F/knCJP8rN8AQugcxo
jXRjN8e3MQwhnndRO4GCMzpI/h4a1tcQENuri2VCXC8K+Pmd6h3cxlpunvmv
E2Ov5EnYF5iD3lvhMTyyqkJNOMiwzkYjurYqW3kfkqlDFMjIe6d/B+/+LNXU
qRD/6AQLvkcvGxTOgmjXlKndFjZIZmgXvDmIUldFudPqHqFrqnqhS1dSZH5x
Yprt8cuGh5s5HvlrFiZjI1gXkeCFyzvb3yDSGRPJ3g29Iu9V7lfl7+dXfrd9
veYBXiMiHhMZTEMPOKXL3mZf5NCzTDUpmy+hlhiUzj0lwXGgOK+I52d3sM/h
qgSPxoRnx6IAopHAiAl05UJfgLJuqoxsJKNfJaxp+ONgfxjMslcVvC53C7he
pSrZ3tUlcJB1nuBqe+zIeniAPXmbi6bdDsP2yE5Ge8GwkSEddvnCVjeLSdIL
rstmG1nN5BbJdao2hsb+R+uG8utOsPL168Ml9UOfaw8MKPA7OSrh2LHXVadH
TXxeaLo79QRZit9Q22DhQmaSpvt4txPQFCQOk1bPM3oN05kDtH+pWgQPVWYW
PJV4jqj4yzvbJlum7vKluhk4LF6BtLWs8ldfX/sELJJuXDCImFE7TWfjvJZk
vqCUAErSKS5lDAp+sXyA5zNNUsL+RTfUFl5ixpfFhV9cy9usdVgN35Y7lbVU
H4VBRdbU1xiYxW/tb2aQspgN4JbH4QVBrp/Hbf9p2clJeh4MBhZu+86gVoFo
bQ+W+wnYNFzxB0W7wO19d21y35TG0q5jGpE1QEtKoTS3KOfRon923G3NErUD
tsGcpE6PveRPM3sJsOfuwOw/CmLU8TUPgDD8s9ZKTSwzmznCZmk2DWA3kUyl
tE2a2tH7rkIv0wDkkaIewDjfiep+za4jMvkSBFsDIjEqiVtOF/nHq7kbgwix
zPt/vsgG/vNhFcdyPLjSMZ2gkfCIoL3WUSDPA6r99m3nhfVVH1DxknapOXWM
WfQ6kwoUCvgmgCcwTVubrecIopWGEsnjHEmF03zjqosmEfRurkfN/NviZWgj
gB633zYJecbzGdRlVg/njvCq7Xdpv7vaI513KSbtLN03SGFSLmuu7nEmj4bp
KVTeGGcOMv+GbGib4iMX4gEEiesnkoyLTrlRgLTNj0nd9ggVOh+9n+uKIqnY
QyAvzA//cPaTD7EpkgZwFk2awbItKhi9Q4ZR2dq+CVPTNYdSL3VZftAngUSe
1MzHdh6bgmVNlXiTWh49yA5LBWufR0DEK5jhN1U0AqgOFdjK+FtY3b251nfp
QaH05ov0B6MiKXwA2YYqI2x3xjw5pKLZSwaI2LvshcV4ZecvlKgLDBnTnC7L
w0Eo0grbT+7CXZjyrKMpAKNeDEeKiCdHMt2Whx/ENjOr0mJAGOP052SnheiE
5Zf2GaHj5Wjzq1UgPoSwjJy0w2ybNrx68ttp3AwIyFIg8rEq0eZBpmZ8sTMi
FrjWWebDEKRxkIzUFzMiTB5iRWelllp8pfnTIb9K/7DE9B64j7UxAbnip4Ce
Mn16NRVFYCnLzsneDw7HlkUKEyXE+J9lxvu3xLH2Zm6Ztnw9EecpKoKDPJ65
f7So/Dq8tofZJR0UmJxXHUCk2ELfNzHb5y3nB0+dUQHkiK/P8LQf1EJEqDCZ
uTuCraTxh4RVrJRdWSfChptwzzg08yfCw/iwSRwwgFFncGMl7SAGZk3BkAE+
iDfx1QhnX3ruMiwvTlBt1Ahg4GvlDo/AhgNCAGSDWKvHmWgkjgELVYLlrlsd
HxBkOSKDQdiDQbFN10j7NYYCB3MsfVyK4TwCT6eduEpHlewioPLRAFXJNB/T
AYTR7XR/XKfnfRE03cEaAw7w4xD/kQNONiRPsIMDJtmfcDlZ/G4ZOrdneEcY
31TdgPwpDqqahw8nj15jE+OIERL7w/RsCQL4u6gWK/YyOsmdS5wmUer/4da7
BYqxjrHP5Jbx4Mrbdr7Nk3zNXDBUfoaQBX9Dkqnc13/HIxLrWI6n20uZ+Bvr
NlUDF+St/6ChaioCDY61gtzXSc619BF7JPIu4kAyibNZTijtB3yAP+BGXev/
Ckc+TDYIPnPbPX59lQJ4AvPJkI9W5sQ4fIt9HW/LJUFQUjM4J/0dMefYdGQ7
E7OCmfbKH91vERNM+LUCU7YasTJSs6wzpFC3pAU68bMTm7tYZa/8Cnn+i/HD
k2TBTp7A6ewefg7hq+pHku6khoJ7GNIQWYvqcGbBdsAAypE9NNKScgewKWVT
FLJMfTr+GAPi7JbTu5bwZTIhZxgASTfKFFsWNJJInzgmMQcBlZkvz913YlhJ
+nFJLgKX3z0++RP+wry+INye9KOxzL6kLEL2KO51lne9zYmISpPO3j4XRA1w
sO7mTXTWLlmMPm85Yx71VcI0qhQQBoYxIO71adR2s4GLuTUrXaBX7x2kAAtz
gN3VBShKkktYQLXtbEKXleLlvNzcx/6ROBFG5CKLEbci4ARDZaADryV8qDwE
WzjOdd1203meL04KVtvT2sXmUbvVbCFhdI/fuMR2D3m27+MnUA6Q1jSfmcEP
iSmAFlhQP9ZPhc57hc49KRarn51wBZHCRaHXFQYNJGmINlUIz1xhTzdInV40
P60ypaG65bSfrQj8RIRGB8NdGSbtwkvUrKQ7sfhz4LB7HhM019qQdqdhMFk3
eytw8dLudBA6gEUx42mRjjjgkxbMoEbOJj9eG5d93kSVn4C1F9NRdydOSbOu
p7Joxx7StD02M3KHrmWNfTbA13C92x1OXQqJ1cxGefwt3uH+xZVqPPCmgYp3
9yhlKUn+pLjcKshc0KdH92vRXnHdtdHI+Zll80FdFBZpRDOPpB8j3peM498F
5psqUz8MPra3VYiwT1jJ7FnhukFi9iBT/rD+ErB1xvP8dAgkZiC+y9PVGNGq
JPUe2FfuaQMaNORBO2OuFRpaOQXa8KAjJ/cegDNs+1e4vvafFAyizWCzUgfr
kZvXfX5nzrqY8gra/7AizDtOlc2GNsrP+bJgOhjXY05HqfXME5VVph8vx1MC
3DS8Y4cSDfdzqgcgwFv1QgLa2Lc6SIL6V0Sfpj0vngHkNygXnZPGi48wdXri
szCk8sDafxiJ7kzCfCdQdPNcF7udltiHWZ94ESxAIMzi927vZLteunQnnnXP
GTeYCNXNkjkufqfEuxWUF8C/u6IILxqgu8EOp207zDogHLCSKP3wxx7Avcn7
tTz5MVAqaTZEImlHkEW3K+eRatGBeZVLc5m+RPb0K/x45IxuojAWLrvcPdJd
gt/jcE+gPhWSyQbU//2jMs2iCzhx3J+/1vse1lSShINqh74ATVxeWz6rj+n4
NGwIUxemyKpTNtghDbtpxCL9xbqaKOhFl78SFcYDTpGak8sRyGu8b4MJnU/x
FkK2/o8lYp0M7IlPlIDmkunRNOnOGFxmaTjVFY4unZ7lg50szhhYIE/gyRWD
cDmIMRkPdmqtl87IeErfB9pLnKComiTm/YOAQWomVCpIFCd3uhu5o74f51eC
+kGEDYIUQcRg9k1Ip1G+CnmVJVtjQ2il+oOdX923Hsfm2JyGVM87O7ArWUF5
6+xUJH0u6+8aJSuE84IIcm4YLUwcLu55P2xOEseV5Q63/P4WytcbWbmGZFLc
H/xofBawA2f0NVMnnxUXm7cGjkZhQg+TtKcUaPIgyvv3L+n0uq9Azqz4x8ZF
SMo8GfpwaBsHj9c+sEwmlF6SHV4a6V5gJiLrBUcHJYpNJb2aKgQ1YNmJtMQd
lb7gATPAczaR+0Bc41Fz4qZ8ohZtylxnUpyLFvRL5nI2SJNMNs5LysJW0UeA
qHxRYWgI6NbV3JVuZAxfaVIw7RNDyxeAo348JYo/0IRArR5UFuFAWxggZS1b
eRrFNqL+VIj050Sv9TXauUBTR66bbtWuex/2iSwfNHQSadQKMcR0Fr6zwrkF
SABJnSNM8cGEDC8ZSbDAiedwMvfY3+hVe9flEqM7Wy2bDLG2YZsCwPCNN3Xm
vWZzq5d2Dp2DxQpVEDS6buAMA3oy/LPhYswDsa/lDlMeUZt/aat0MCRTJ/K9
y5jf6ayT8iVgiAiAnOwaD7lZQVblz5631KuxX6m/OcgajOlTmkZFjK3zWO6C
j5LrHT5JmgW5q4qUBxwoFUQFbvJXRSbERd4BzZut3rzShSXw3P3q26BP81J/
WgCi/qGd+tpgkan4UC7RAKgLq/UPS3gbDW6C/7huIVEw1saqazU+A2v1pqyF
hH0omfle32rLC236i+N+w8qk5vOJul7Puocfs2AHnCK6EArVHVUXnvgv93pJ
10GX1xUpfSANygBxp35LF5kVgNm4ky7J5ZcayTjUr7gjGe0iZUDq5c5om1UE
34NjRhiddu4YntAkVJwxEK931llQ1Bj+ds21VcajC4wLTBqlAnj99qpuHKlB
VezHiFpk7g4OZifpwZJMRqb8Lash1dMXzqkcV46zJuqXlRchpbN48ADl+YWQ
YSotxMoDgaJSk4j/0wpC8fH/Jn4NxyWBrDVPjmMIrmGK+0K2M3UmFgSBir9v
CBDJLDp5h21NhZej1or8ilNJoU6XKLMVNgJ8EohjUBKES26iB1mFiWW5oKbx
AqL1wYz82pzle4qfMLsvSDYpFJuvziopFZ9Zkwrk12ia0vrMclJDg4Qj34E/
g1yV7owGwRNPHhtgQugWhZtJjUxFFPQiso/6jvAoR1oypmLYGT6jbJSJ5WsG
WbCrWoB9aBxqj/xb8gR2nkRxRaRn7l3GNruHS9FMDbLtsgcp1MhJv3KM4606
sWmAJSlosMkKH2PGbttrDjpCIVvSRhFW3srLJuefFaWxtyQRiZHcnsAbIBZD
xNPxwm+hPcKsVoSLXWLNXDRuffpTtKjZeM2ODmIoLHDxnala6/3umOx65jUc
Izg0dL8ncSjNyReqvKksN8dRkrhoG8/qomOc+W1xLIB4RGnaBAz9lrTQpRvB
D0pqzIB2X9tu2aO6ukpc1bixmqCt24GiH74mO0Yvmru+M/z2trGYZ+IXOqNz
4tes1CRmUIw2eqU+Ki+lzaCqns6TPT/ZbqkJyDtB9Mp+mEaV/01Y+1sN0RHO
8/Ks/ppYhevWetWV/JM3bFbbcaMAHrG91pkv7izoMR4rdPgS3jM63SDMtCCB
e0xSidNFDlBq3UYn4eYKemfzQvBsB5Hpgs0GIfTSkFx3Vx4gbG1++LEwJgLc
lar/SBrzfiKekxd23Q1P8fNrWBE4+gMwUS9px5xAaZFBaTJwg57yqF+6e21K
UqsJ5TbF6VhA/WSclAn+bGtMxAtuljGVKLRxehYJJCy/Je1CQV36pvEoYBSI
S5Pb4hNUzf4gR/IY9Zt9liTY/OxBlCeTBwOceV2b3G/vUC3C2ERelQgNqUoq
OvaApdfbNiV1P00ToGiX3QP8lS73+cKMbaenQRKhjR2a6H59wuz1sNHpZzwO
EJhmiDrc6DUuudx+kM51j3xJA7Xhc74VIjPXYx9Vq+G74Uubqf74H0LSCHjZ
AA6RKTGzIzQv+TZbZC/+R+n6auZaFs6gANYDVTKt6G5pW6zR3s7LHGpE6N/N
K/wJryHir2EfujMVt8wEfoxDDBJh+vSTrNySrzucN5CXJMs0AoSzRagxS8u6
F39Nehrk0iQoipjHkYZredh8Huhnnh8E/jdlIga6DW28vTSIChJMPGk+nrR5
IdgUxMRa0rfpKm7oQ1T/kJQ3qLbjVZL3NL4SrPqRcxLFFbzUQ2PJuLVQ1PVj
4ii5iXpcSzytDeUS6rh/18EBTKTg9QRi0J+oGpEkc8osyrNC5/zcUeuNekpR
1J7EPAKieoMWElW7ftgaTmakA3HtgHP0msMymrNlG4YFmTRbC2xq9KdT9ze8
r+5qJ1R+B4DAyssW95A7ijJzGBzHcIgTXfXpWA+CxRR5MQjw3Cn5cI2WFk5w
JxDM0jE8mT8AdKFOkKPgDMd227M5zqC82ZdjAdwJXrIq0yd/cS5m8dtvLjJM
KXqj4NeysAesVXYbfthJvQW7BI89xfXzIMKc2I7U5WZCNGL0/7OmACbPQm4b
VgJ3ycwzcFczVoHTmqrpGU2T+JYzZ28Avpiu62Jpu2RlN5M3R6V0a1AK31u+
z67RYTR7x8R6I2qd6/JJXvngCNMoy8/FSkCqhxi+3DtsgCwfcV+MK8Al8/Yh
FY+yRE32jHGk2j/00sR5Mk9Bxtxy5hCcsT6wZ+guXNW9VXQzyOPvtZ7woUIs
QiZEJfxpF6pdpQ6cbXrmi+fR8zQsYlQkbynN+ggUIqZoj4EXa7Yezu6ZVAem
aimnYoDB032FNuLC7ujtah5xojlaGXittfcAV1KR0MEHRS9e7pVVq7FCshV5
XD8UWJEqzxTawBd+Lyyu64rbVf5dPljACdv72v69zl0BTKC9leeQOeC093F/
J7mkIhW4qE6o0v8wK90SmFOdqGFBkT/wN/RIzRvCUcsikf2IR29BDVVGGxyV
pYpJemivbwuwiqydTlCn0nBYBgjaEKdjXEMzOiQTCXMxC/Oh9w8NqiMrk8xj
Jda3r6Syrc6y5jgvtAz4+0J/5E9oV7MXjV5mvpFKlwkVNSa1aCQkeMFOW4bW
+uTn1zuxsB8WHqkX6iyNfRhDcmMVLc2k85gt4gWe4+I1DnJ/Ptm+zkb8c5nD
ebuVvLTz7TSJllLvDLluvvbaUtY6/klVN6+T1prfbHMApIdxphDPuhmbSfYA
/NZxGzEQTgATaER/IsEwoM29LsC/7RL5B1I49ZozSt/I9FhJ0BqR2PwF+X2S
8uZui8cKR95GjzOICazSwt0N4s9GVT0dxwGHBmDZ8XDZWHx79Oify0nq/rUc
qZdAGx0z+SFA8KuOU9VzhIhZnC9RKIml3kKcyGBvCf4RJukTk8qPm/fTdLVt
g0L/DoZiTT8qXYtVONrXLowzxPwYse15XLMGmRCu31M5nufvLA/dnAtCSb8b
405bPSzMzSnZCImLrGMIBXF36i7d8k7Za5ZjAM00uR1p9wcGxksUgtHBFWry
i1by/M5V5uoRCmfeSBHSyVA3TzLipIsg4oJ4aM9Mj/sZk48WWil9ffdVRIp9
PDaXXEulryIh4yADUWVRUXve6eJbRVYokBKeBiQm0p4TAegmkP+t+fgZuNIn
zx29GyUnVhhO/zezWBEIEjlHV+EFQW3FaAms4MX6Nj1eql6KfP/p/5UQ8S52
4Xm4v1xuPmGYonfIsEsJoLpm5zm7kAeNxuWxM8WRPbVC4Cr8W6FlMZTYxX0I
EPlpZOGnY6qOqUhOUgwUZFp67LyaY6h4TTLczZCums+/uH7Sd7xZXum8BnHe
iXiMq7mRLdz5WHrg3mCtBuYBWX4Ur+kQ2QayoYgrzJf84OVV6/EN2J2xL2Mr
EJGhkzsnPJzCmXyJwXNU+VtBC2D5K9pS+dZR7+kZ1+K5aDJ4QWH75b+SZYrg
pIt4AwwX34byW/jRJ5tY2yndJUwohn26CFhxpCqZm+kI283S2udUjGObn/Bq
xPPy0vXWn2y8Yww++nWzOJRNkObQH7Iumb9SOqp560LLK1WmKjbFBtBEBf/G
keqLduws6g0i3wBpEWTp3gvIi3uetPCS4iTOVwsltt0FPQIG2otvTz36p6kr
2eIyatnnAPtooEf2EUkOmAvKme/KxaMKaihsV6zxcuceqmdYztu2wKgyDuY+
fIf5xhYW2OlM8EiIAfQzX8X68LYU+cxbj2Jaq+K3lXkGiiUur+2Egam09LGR
T8HihTiyOhhV+Ydjy/4VZoT/7C0OX9/PU6H+fDO+9NacnLdfYTptcYda3Mi1
A1K4qgIvvwRkzQzqB8+cYQkML4ekuiTrDxHojZ5szZo01SIq81hr0Ah6fFb5
nxM2lhRjJZ+/lxljBpkS32eGha6Z7DrR8AecEtgPiqo61FUtw2fF5iFI1mFH
jxcZpH6PyV70LMzIhamohFA/swYhLJ5P69DYGZ7INITC6/dDDDBT/daad0K3
VNsoH3PX5s5twmkdDW55RuxyU3+F2gKJbnMXCNzJ7kr2xXOEwA3hnrI795Br
ZCTJvDMqhbCFt8k54XN0dT7I7NOvc7QeMQ7b7mBkl4FBcDTRWZJ8KWEnkoQ4
ss4XQyZCVileKqlVRseRKXJ6ovWKIuqojHHbW1VPAAhGH8tWHk8PjSC/haKf
AgAfxNJPNwcOiNqBKRq6YJVZAOLPvqDyOVNfZs6PVO9f2eZifnuJ4LehIae5
fJenqg7b5NbHIsh+bvPQi0RdRMHRaR44IJ3vkYwt5ihfqwyTT3y/7tti+Xo2
JqESgwBvCcsHJwHBq9vFautGpbm4QtGkxtMmFwvXWJ4EaVyOJdMuad7Qy6kv
XwV0L/m07FSc+d4+zQnAYX2z3C+hkPjoKjxOh/q4ZrAdZX3LGmdv98PWhjrf
eOlpkF+eqLRaH4a3mGCRx4r4WdkMJljtyfo0S9ALKxHMEB+sT4jDOpUx+Z0P
KhCVoD5i2aefZ8a5s373bGe+CkRPZWPBSplqLpXnt5EmSEl1K6p37YdUXgLa
cjWiOZ5MivEDnYs8Lk8qIqMW7U+3F/79rd3lPOBtnAUK9W1PAo/v61IjXO4M
1rJje6xFbDqBklfySVKWbw1Jy4O165TiZ3+vf4CsanEddocgTgG3r6rGxbj/
Ql7c80A0z+dsqgCNBRKtyCzPXPaDqC98PVZPi2xkJwbdIvDySI72le03BVUE
bcCtogsaErOzT6Vwjh5j06gMcIZTofW07h5NoW3k6c4rxC87UAmznlr8G2V0
oarsI8I1cuf/3xEOy5g7WT526o9ESHKxkq8o1r+RlOw/ThpeaFNbyogjEubi
GYmq6WYIap6Sf6JkZdfgD9rbuwtLhMoc4BoMbw4nyhla2ORQptK+xqjqbPnm
SZid58I8HLZ4zGJP2DskSOL5bMTqhHu7HeaiE3SvcnHe9Yi09R0122vOACNo
9XZoRhw1yZ33UiEsxa1YqMilXVif3vLf+L3w9nymNrGwMhyqqSl7ybnp1Nto
XlSY3M1g/b10SxlM23WpMTR8IvRYX9ioAK55UdQocl/rYD6yprnzgidFdAbH
2b80x5jRq/7qNC8SsWcqSj/tsOiTtq4OQi5BnCDEl+fmM2KgqhKgZq3CKDOx
EEsSAkLspbJtFCMQT/0+6Kk07JeNAPu5SKD00s2mOwjSW0DTY1NZJ1JluoJ1
schm3bHhTgFhlQXIj2LyObpAnP98qd3N/3Ablr9eDtHwdle1jTw2vbYGq6/3
BBFGxnoAkGz0JX1iye9PoNDdoBEjkRAx7GkZE75bUVlCeXYgkWH1w0E8sNwp
T4ArhEZrMhC/0MVNruNoYLoyr6p1Rfm45N7NvYBLBys6NiLcCWqQoiRNJmrQ
J5Aku5m+cpoOUZWabERcSAM6svnSQ3ZtA0hJdM5CYv26dgwJfCo5FdpPg3hK
h3cX7Bw4ir7yM67JvTFJMp9mfiK8xiaSP8jl4uIXXJukSAJU5f/fL0eMLp/S
uPr9XaYaOPKeYZ7HQlloFIO2YX5c5/lGHBM5TOpWK/CN3lUdsDmN2Xda9dHC
cq7Hn+Y6/kreuiItxQ6KssxuwnKO4mzGOY95Lbxh4QNHcQXxCHnnGQ+9EQuw
JTe8bkgil+kdcyEC1e7dBjkA+VYa7OQlMhOrZUSPNEw69cxbXjasGBJEKw+r
BfrsIKoZVigY9I2CwPzBFsKuba0XsOB3vCU4JEXG2Re4ngla02wyT+kHVkLr
lZP6kxJoE6F0L38FZwYpoUpQwWQBPY5AeVtbebSVsjWkRUNyq409h+H3xpJj
UY1NYvFofD0E4cxPvNDC5fObZQ1COi9WgvoKcn88VyxhfZARYjsBtVNnYQo8
QqBpoNPLgE7G0zrOPEVIiIH6fEsTgM5lH+UuPQFg4iEOIMayubto4jawHpbE
SicO4o0IoY6nNjPwNMyg2OTKJnjleg6uCnFJDaD1ccqFrpChN8GTY7cjnHnf
90JLWG6322qYCOAM/TKohEy1ZMGjeW152po726MQ767kaC6BB6iSKe5B5uBP
++hLDkcrM+uLRwrQC5PlclhIcwuTtSXnaPKQa73oXrpsPuL8Suw+SbZ7WedR
xRcCDly4IQzjMvo0LE6VUokiFNq93SNz8fLdNZCv5R8GU95OnOHoyULZY1kt
Kfwklpes5uj9mqkH3K0vm0Uy3FKIEx2NK/oWFvPCdFeYhzpvrWW7cYnCX2Sx
vFuipxY9kPeMLo5Q5D3QDCel1ZzdcE6cFp/B3FLa9Cc45yroHl0oaDpqw5lJ
FkNiNrs1GYKcV57VEYE4FazGMVeC1ovVa0N4VdaERzNNijkOfogzleMHsszY
sopsBjdcTHocYXuzDub+C1RYBrvOV5PN4TKinHQSqFKj4JrHk6Nz+d+qT39n
X95RHKTzhO668S/4oEe/rM2KUJRnFOmw/Cq2KelcV8mIs6zkHvtRECVa4TWt
ViULBJ8naBfZjCJjY8IyK2FE9/Az6w1v+rBsuwfqyTQFJIzR3DEzro/7myIk
dOQ1S9ZdzlFwqjuZzi/CU72ZotgFgkxe6tZFBrjiCywJALAnAsX8DKo4f9rP
bNL81qKVPtOqU0reGv5WVnCntWlMGoIlsH7PZi/f69heQC2wJy9erunqq7Pg
ytPyjh3UWNBJs/dc+CinR7VLEqSA+c5UJEpQrQ4bDt1IioCw/3DrzkqmpmQO
NVrgh/borB8oKg8j5s1F3feg2922uJoUxDktrV1xWujGyfDBE2lVzAL90I6k
Rz+tW2+TH72iXEt4DzGweldkpiSm8pcfZvu5Mt4O8C51PgETG/qQdZjeqdhr
EoMnyNrT+e0t3P82I3iFToirjFTb08q+6zncfJk2ZL9qGL/kpTUlrfFNKBhz
b4Enx1Kw15/GIrPCeZ4i96urOVbl87Js8U5NKWp9vp5IeyoaK4l9FZ62gJSW
Qqyf2qpDESxkEwJhn7nj8ixwGnkpWXIpL/oltzjqLU3/MtM96Zlu4x9df72N
Ii5GUdD54OckHp4Z8ynmqNvoUVxsFuFFWM1tTCu/A5RWWpTUxIt5IXtd1zuw
56FtHuuaig1c6aypTg0iwyjxn8iq0Zz25XG2/TWw+vSm5/1SRz9sHD3xfMKa
wMXQiAVJHgA9HCdEhiOkovXjfzHNLJpezj/Hbyeem19iEJ2M1dLA/C1fqQo8
xXeKJeowmMbWCqIN4iT5+Ww7v3phosipNp9zpbMrXYJg4YkjlRYSlmtMaHY7
N43o+7kw4E+u736VfNm9qxcsuoqrTe4NJQw7yrBFBlyeY/mdRz5s6czc9mnA
RTvZugs2VdETx8ZpRAGJn7ES/o3WjScij4e2gn7WiD18SuahKGfJtad1hNHX
0lbE/kfzkkHHr6W6epzpgJ2I3jKSnFWHZ3slwXK7Bav16MeuVCMebSjnyDNb
vFwPzaWe3LMKsJF/38slhJMpA3GFUS8UglfwcI7rjw/ycsUkDQ41+URj3aNa
gSHZ3mrWOAdvurSXXsA3T/payoiNWApJ9AUa0HLNVw90B7/6jOBdc5PDM1jL
cp3EvE4ysVeEp7r0ff1noUhWhMf/xTL2sS8jo7ORtsuzA1OFe6wQ/3sHDqcE
ACxTKMdoUmKLrhUSuaefLiqvFl198SnjgTdvosHmbFbhy6Hhx1XefqCcfrih
24dFKXe9zdIwhhBr3+zfzkeDiMDiDu2NnQABHBTW+G6byYX+8iI2yp375g3T
I6o4/cEGj9d8rodFqmdUQYDIQ/bP5sgHHD2EYAhCnRtNV1hnIiHkD7kV1dhU
dUSk064Wzc7kV56AsuB+ANXytu0YS13Q1FjwfeipBHBMrksvCCaGSEG07cFR
WqjILzTIJpwntAhhtrEiPXy5YYfw939gNHWmj06uFfTWOMRJ5yB64VgT4GH1
oOp1Q8oUcBpXpVtIxlDswo5tfbMYaQlq6hKqZmXO8/bB3SO5kK5CZgcZnzhq
BqDt4/CC3himnzB//LIGg8Zj4MEjbBFusqxuBRGneHJAUPTjLogzLpizlQ9E
kfqvjLFhGt3JocdXLOFFtZ1L8Q2jdcaDYhkg0qPFqFGNXXZjYX7dq0SrjkQu
IaPOkv+uyidbZLcz64p9beRA8crYoZd/Bb9NBJRSebS0pmSN0Oc01NGfddc1
y1vgh0EShHDQa2e8SWHuZ3x/liwhG1POEATWCWE7SM1EybHbWNgjtCPocjeW
lcCjW7opqmzKuSIXsKb6thOUZWBsFGqQB9JxPniMLn3WsySE4nOGRFC9Z2ZN
o0dIj6ozYga2faFJbo0bbh5/oPYiIdUuaaEvUcVkVJXJC+UFdhgKdgU+1wXs
T4NAtTFGXaRRpkeZiZ1XwfQwmC1aWAycTwr02aYn8v4AUkImgdy4cAqo1bqK
yk4mB7NwjS5ZBvXBTYO7uJc4YvTCnkWIVt/8wF+RQ+2EFHesTSouGaHJHHxj
fEhS+BsQK7t6K4gyJWLYqhH5PsdgdqkE3c+Urfk3zHTanstW8SWk36vkGZWp
fDLUJJMRj5+i5ux2Zv4JMGW2JP5KuNwIFn9vSAGAC7z1SNyHhmY8C2uOt1bV
7T4S+0NM/Zd5K6EIb2Jirl0poq2KrsDsM11pC3uJeoq1l3eZIu2r68hbRtbK
UUBfRey8Bjlt0zloBbCDUR0cbuaJgUvIDQdpFY+nllR9wNx/DpIbDALKRPRH
ClozUJ322zZjwa+xmbXXKZ5reI1PXI4gB5HJDRJJn4Jhpd85KCJAzs3m+WWc
IV4fJItD0Fu0YgE5Ac49SgwnvakgtRZkJoJCGk523FQjFU0hsQVExT3hicWA
vAaHMzNr/9NepyOXguB+sMmWtgbB2W7g4l9w/ovPVfd1Uyx2qKt8dGuYtuwG
jjVDV/x/nIe+dbJmwzlFtB/iIN6344vr6l3B6TN/hTK1GZPxFB7bgJJvH26l
x4+9YRQ1zK/HnTTS2wx/XbqEmlMfz1thHWmhTyDNp/XN4gNxD8wGN++5hpRX
gHshl0pNAfI28qg/frrl/ReY0LZFa+GXaYbzZksmD2iZqrxR4qhMH7l+TOWg
uQFj+Phymiwn6xcBwCzPCxsOcto6mIc4nH53I24RLju2oz9tZmxFdR2ygj/z
dVE8iFqf2bMU0C3qhHCSc5vSILrAKtknsd8zjJ5/sIA46bGQPzpp53jBMFXC
bzvYCxCtC+H0ommpVo6TIlAYlyQ3FTggC3JoGxWoC7ZFo1DUyzFV6gYw213i
Xpo1sRxrz0vDGofne7at6KIQLaniZunBu+IzCB119C5dBXncA/uxpy7rAATA
/MyfzHd63/djAmiY3oagm6zGLzHk8siIpOf/zYdJGZ2rWeXVF68XV4RnQihN
DIC/2CdpNfQFLqa9wag7bGju98OYly/glcMyYRGpjdgW1nMZRu0AypPLvD72
yJfflk3hF/g6nNxA1GQvUdcNbBHrhy00JvGSTHX+U47eLkCOrrJ3n+VQKusc
SOzxRvAWXr+L7ds8P1qqWbrk7vaJ1fHQdSUIXLnZu4kJ3liTUysv4S9CkHWX
I9X8g4i3rT/VY+bq7OS7bfyqA79aGwf28kQnSck22v1rn7m2TH/2mJX9Mg/P
xe1RUOiDH/U+SK0ZeUV/ZN0ootg9pt5uPjHuenxzZI4QQT8zjsRxPpcsg3ap
A85EMidhhRA85Zr5RbYHp6gdRL+2Tz3r6YJGyzP8IgUcDnHlM7NAYbV7Q/kq
/lVu7weWmTT5huduA1lY8uo5Fb87FcxgZ/ltJyYOw5BFH6bvZ7XEurdd3wDe
NEqc/GsZLNi8z1PNFsnPSXssXhsIQgVhKaeJbpAsozJ2QQNDHTI57MvjWhyw
wMl02zJJRWKlN+Uv6e0XohorNGCEir/XKOLATSIVkwWPAZONaz8hbTphAaWX
qaxykab4FnrtMtCWz0jwI7Kvec+/lATSPyURubC6VUMfpdPlxOby6ugiSIcl
udIcMB423v928f4+jF2gVtK5RjlTKw14NlRMrm7FijXFySkqcwoDNRr6rkMI
vQk52TXvsM+TMDw01Z59xkZ7WdrjNueZsJRJYpzU3OvABZgGlvWTitp9S8IL
etWAjs2C6o6k3NrtdPO7rBNb9hau9tLYtf82dr4zHWvYloVXrhsStmuenfJl
QdnqGkcN+jK5q8kUPV6Q8Xl91VcG26Zw+qNyXttoILWYqc4m2iLs1aWgOKV6
tjk/a5feMmpT1UE5cBETua7D1zX3QggTwPhAHPUb8HrY/cTdFhbgbS17Nozs
DcDGtmOuvWca6vtm9t2lhj/I4uzxfjQ51FlPmNJhxSd+WYf/fpc8hPyvBEfn
cBTbuIOQ6bs2WVcCxyGNuArGIokgrFg4BCeZtLS2Zak4u/z00D7IRBcPc/P1
cOzNnlwj6LDrQMILH01GzcH+RxOYp2C2vzq9SLE/3nO/X2brdTFV8lJExeu9
2aptIqiYBP93ZnbFeDIU2kYMOV2G5Omqi0rPIyhrnajYLXCWd0yEZEPjJdFQ
bA1ejiWIrfmEQ5JhwUrZ8AufbJ/EiZ9pg7ZoTil2zSMuZYf1nlMTQPJNdJIR
zHKEbLzll9MkiaIhPXmvBGqKvYvqYKDr3ZNqE672+IAmZ2r5b/FuL3G+Ne23
nO+COOAgPO3wFQ1Duv06oYi9BeylzihgwA3gCt2UyW48s1+hmxmFs1gIYgAs
tgnkTj3zhg30+m38/gQuUGeBnbGAmvnxEZHvhAVno6zdMOn0+Q6k5FnGRnPy
4KAHSVNWD+pY9l6ISFa8Ex/qLKWHsaOTeW8pulO7835QT88bCiU72DyrMJi+
KfRxYE/T6IDUWpSXjyNlsBg3au/J6LclgbJtDrEckzJxc/ExPOslwKSF7LVZ
eI1BN8JgktJ0PHnZh1ZriGfIw0Duv898h0cpAKkfE/3XN0GScbFBWrAUx2fW
ADhXnkqq5HCB5vZIQNchyCvVptRGHML07EmNrRUdH8YS7qqaNhMtM5tXz8sn
iX4VnvhS6zUHHScOmOzd89GbBwE55b0mYo8VYmXPBU/oZ5afsa+pqDsvVUr/
dgCNqlT4BghlgtaUo8w/KCq4gH5O4N+1820EgIzV/DZOI4a3bylp5N0uh4zn
Z7gCuNhHRv+NJlmdSDt2+jEA9nEU3FKoeC+BCTaoxTtEajcko6/FcFsXjnm4
Y4p+BNoZ1A9EZuA4KG374msuE55EZ8khCEDmUd8PDT9bRzkWBXUfZreD6Gnv
7fRpVX33NkiCuI1m8bB5D5o2Y1axNyFTmFKmmiaTY757HuHV7fuOaPgVozIL
ISOgjobny5BeQ6blPczkvvD98YckWymsWiLXyh5RyaRoOZRXSQU6v6VpyYpK
cWUm9ELoQRoghhHs1m4fEZbYeRCOWeKYh/JXrI/l3SS8iBYYVuoAwiebJ/ps
HXPZ8fH6PNmAdpUanfUFWhQigksMSEhkuei5Y9xdFxvKa/V6pkJS9gskMvuB
WRlYaGyo7lkdGhexo9ZRh9E7SVgJyhCpP1GRhhVuVnQQuPpdrVB4QELmA810
YgbJJQclGstWjg4DjkXNdM338yN6uycO/umwlACRZhSpqkjN7ZSr4OCStsV2
z0e881gTbLQuIo718eR2s25JNc8oNk33oPojtyvvkuO96DmQSUTIMg5piZiV
yZJtuw9wgmCpVJEC2MtQtggvBhveOpw2gMpvaT5reIccLb5/tOa5R0uzinZb
TiL7sJE/raWxrN2NiqgT13IIUTshlCL8z6omySioGjY8NcyPJiQ5GpKMIPtQ
IjWxU9mLx8UPj/fuI95roUpUKYfHFOvanNY6Ieozs+N24TUKEMxF2XorUwFE
8rHXgKqwuIce/c+r6Anf0tvYvnKOQQ0ZvDZz5iceJ3cFMzMQXXUHrBVL5Heh
3PoWVghINIoLD3aOXfAuBMzrkYe7RjgMN6mekL/1pyw5CKbin2ahRtj/mJjs
Uu/JmGXUmejpeLOposY8odx/+e+6a/sPRujvj9U7y0G+xsJsUhkTD7+OmsU5
c4wi4l50Go1PIN93UShnOSmrKkoX+VAOOK3l2L22fWdSXhf0526m0linf+yz
E2vqXprlZcQzHVWoJxOKPCgGyA+OyNCvtvq0U3ZshbZvBezwZZ1rr+NNuU2M
Ba2Srn//97jznqcrKppeQ3r68r6YTYX4COPXCptgGlhmfhl3J3iHCfQN2qzh
knFORDzHnZDmyXrB1zDBYmq3XKe8/B4oheFWv+mPpwh4sd8WmcWMMOORb/2p
+4uptQc+mcRs+p8ovy4/0rH/K1fCtsmg38qc8Ea3ocE2xuribylxD85m9dDy
YUDOBNwTohNkqNMBX3qUiJZ3ILpM9bbu+eiemt8ouLpRks+BhM5KleIyyihB
Ld0Sdc5BA5v88U+fQh4D8KHWGcOJmXiJ98179r/S1wYdroi6far1HFmY/rZo
bfsjeJeVQkuD8KGO6kDWd15TAJFNaQLK8uu2mkSzZPQmZbp7lHEoV1FxHe1X
RI/dDjJ2Lxw5TCfnWQ5Z0P7gjeK5QR0Rzd3nJsq28D7/NHVdstB1FDXdUgE0
lkufkpjcMge74992C2KYvtrbkBIrd95eLRm0sAw3n3c4mTrexx3voS5Rf4rf
12OKILsK9afaQy0EsOxWZ03K8GpFd6nvspzeNNNaPUme595xcEnvacf+l6IX
7mQfY8WvSJlcx6MLHxbbdqxMwESk6Toc5wvCTmdjWygJD9vaKuNcNeBL24tH
WJmgA7mBsDPIKYTEwnhejcay0+v9vMIkQJSKd6v9az29gRt6HYBVJM8gSkWx
GrduaegXTGuu/qM3NKaqLubO1CYxwb5uZEjx5IBrc0iZ1KjPvXQxdOfr5Zyk
QJSJ1s9xejsp6J0Y1rhyHWOXzvK1+kv3ezoMOT44BZSEiPF/ystya/BbGvfv
FyjPzyrU8OcPhEBPYrYBLDZh1a2yxpOAQXEVcomTLNJpuxOYlFnkTxEHww8S
nhKZcrdmGvrQSCqUBFgiGLfiRhjTtYhacd8N+H9EVOXuw1R3mJEQKJwApYMQ
Fx0Rvbp7d4ljjlCrjNfkgZ3JeWLo3FYFsYAXa3Yqk/ONkO51Si40SXCzgGJv
sjw0ZiPoV6ufA7THZTTG4i6jNoVKEGZsnM6hV6XzEkQwKGdqXDsoW7l9rhmJ
IMZ61Zx8yarhiuXbQunQlRm1TP2FACUbcM2FOJ7QfJQDzG0zO9M8TxPVybbN
5eBIvRNGBVuvo6qE4PAKiMNxwRZLunORn2kuNAdJK273OgIW2uW2LX7avn8r
AWlhawM99lKLfkK9zijAQ4eOtM1MjkuQ5dXLWHIj5ztzeCuGH5Dc67r8Hffn
hnSZ+1pCULPATvrAAXX9nYhXFML4+Wr0ahpAWW1FIJWSayjPadswiVk4x7Q1
OVJ4NNIlM2Lbjutuh9c3SBs43LTGQx8N8RXG6qIiQ86M65Ihjn5K7ZwTTOnZ
KzsytmbkyQai71RBsDgVnVI4XSRwXbT9r4aZM9wYdWioluYlXKp1BDpI+ltV
iDFBt891qDuLK5ZFiOWdqTDm4eaQD+ejJQNEsY8fqwxttXJ2Ep9tV59RSJqF
zFZBfsVvUyaQtX9DVk9i1jc7DMEfRfxAxuhG5Htzsfh2/ukms5hiJkJjcf5r
KwiIt1DRki3ZmDupSVjnBXK8C13ujkD0c4mmzrBOdeCMk+7fYhJMZUiFJv9X
GpUIPPIBSEq5q/BFKwAOYGHm4Ai8D5UvE1PQN6mqsQzaE+PTNy/yoYny7bqK
STcp0RCXhTmhbEKuZBypfmMTPi2sZrEiApH9zFMCH3/dE4CxgOq7th1Efqkc
Dgh+8sy4Kt8mkR7pT/tZiv8JXM84cM3+noEHcmVST1fseEd5x5vVPjf5LOrR
/VslJ3Tp/FgGo6NC7B4GVZbbn4M6TPpnkoRaqosq1ZdXrAtQH87I7Fon70ZZ
tOX1cBOfyuYay2yWJ8NuLuyDjUKN8M/lZK4CHkNW1vUfji46EfEBkHPvmKtn
k6ZT8JIuII7SeZosLpxJYVznZkWiqeg8T0BT8dd9oBkP4bdNhJCK6xOQl/aN
3Db/5J1S9eoFfQh25j/HR+WyP6DRdhCERyoL2IYtSVCd74DeaVA4uklWpGsj
MPoktIxdxbRb1kn/kZOTDf/4w+vkBxoOhCOC3clU4MgtVsKE1xaxb1HqHJwI
4eA3GoVzhDeUfnSwtLfqngkGkUYKTcIynqo+/tPKxS5+KnLISwZJhRp5qRvB
GjdG4KC8P0nF4kSr2HFvFjpRg26Yj3aWV3mx5lYe44H5vevEoGwrowvyto1G
Uce68zXA/vpoZEdA2j9oSbKtVFbuhy/Yj2zpIv6hnFclTu+2qTO55uDKpnGz
lEGyL4YFyI7NlaE/iF9g1EF+GUE3Zi8gLclY6PeKQQ9B8UxNLlNqbxx7wkHA
nSqUWjc6Ww/fviVGKrTmRLYVtyAnmUfOiAXt9ZscwvtzNMRj/SYMa7c0oLpx
LwgFX6BcxM/LZN/7rm3fC9dB5KKwRWIoYWGc0MUXbl7nV9z0tmLSXt8WdsgC
rwp48DkJr/SPBLWAwzJ4yN55ERZqD8P5BbpYUiSZH05MX43S18W4O+VdthUU
B1FOicygre6BnF4NLQV7ND/MBiPasUux7PabEKSnWo7Q793+3jyL6lHDu1gi
kNpWzHeH9rAbjCDuSskZuMEnZM0uECp60DGDP4zveoso5Za3jQ1XFkL5a4cR
faR5WSMUzt/3OYetgZSBaANBwnye8FLmjouDjxfXoBMctohjOScJxkZeL+eM
gcUA0vbbGe47C+Wiorpw1fgyRbP/lLbQif4+T6de5rri1bhk2lz8rJRJAKna
OYtQzZ1f4X388vV8IwIftsfFJseZ08+Ftjy31kH/xAcxoLXZduq9znrhuKMR
wlRAzC4587qFmaHStDgrhjC3fqRmaiCDvGSVqpy6muX7n8K2hPye5QC7LwBi
Ny3e7RUH591UacxJvdMN+aCS78KpwSprYG1zmXIe49apy4zg47X/C61pP0v/
fAVehTeIhOXkDKt3W1WeI828fi0HXDhlvhALJwBIv0pqsq70TTqTJvS7uU1G
It08zbDZfhjcENUiOZRx9RZlOHaF1Dlr0EDKRQQSangZOEaj7+8DVeLgHFY+
cpBzv1eA1U+IxgxuoXXfNzVNMz1QFCuW47Ouwe1qpM4PkJspDNrs+BxN4U34
4paHXRGDoaE9cPysEFDHjin5cUaWoiVpik/n2cHCaCRcMfpUzaylWQdPtaXH
u+cRusmwbEEcfRjnwNUd5ryVinAZG+uSukN2K0F90TW5siWUzqfD1lEs/j0P
psdwx6z46NN5nWXkqJFYMr+0dUtTokpCKTDY+3S8NDv7MlBCH2+1oQCHXNBn
QQ36O3cIpeRMODxFFI21Tb8RzEJ7gwdSiiWUirARS2p9GZ/6j3XUxMHQDpCr
0HTfnC8bf6v8zvqeVrjardm4ROcjtwtUSWdbA9NlrUTumkNyqGM+YApxoyq/
lYtERA9H6wCi+4FM3ylyz8VHebL7clD0SqYKv3QuQUP0n2MQvWxmKBzyw6/m
7R7z0ImMomuG0OhYAXoGnvl5fleMmPqvooCa912UwcqTWiJXGHxlI4KmfZXr
aStSGG0r1C8odBz5/zefxIz9BTIPHhNfC6a22kr2T0CqMdkaxZrlFlGy1TLc
6TQfRD60hDDo8EVbXg+gOXXs0fqtrGwGN5QEm8ntA7/GebEf9FxQCguwecUs
frVUc2yaeJvKzwDZOyV1/oeIjQLA+nuqDog6CfEpuLxc5yV0zMzj4StJ+gMB
1K9e5LOQ3icOKcl3whDHsBMlbUKBVGFHtRjqd9k+bgzPd/oBvauFWifxmtLz
sFeyrOnK0tiqD6FwL+1dIDh7wEvKgOKmkW9qpm7YUi3RmZ8yXODeBeSZ96UJ
j+qM650LMClsaHzvXeNml7AtNufPJaHUhMXmMDirRMgVayW1tOsP8DzyARKf
eOWvuNBYgPqLs4nRxp6aOi9TgcQb4Q8ZaiDx2qCJwv2yM7b21jUedVbnNSVo
I2jA6ps8yvws6tfvHfUPfQD4iG8rvJqkeAI5IR3ZT7y/rT5/zz4kc1kNRVhH
HMU2JEbmJY8mvnb/OKrQaZAWYdzLI6PKzUygIzFO95/nRGhga0jKvDHBkYE1
i/Q9R9k7CPszuMgsOgxbu6UREzHOwLyw9b9/k1jA2vowrNOxce6g5626c480
l1rP1LlfQ1UA8eV1IZOqIG5mMwLPvBO9VNrhuKOkllPcZazqec2/KAVFbaTO
qBNgVuEXoWHqZ6p8GQ1OX8ZxaMG6hlIk5Z+uTYfkUst7oZBjwWp1AZicA5AS
dSxUWlriwqVyx/LixIcs7sSaARUjo4/qhQ5JkvY3PodBq1pjCPOhPCEZjsm4
GgRgO53DFZG65ufdnIEUgXKNsjIsgmwh7BxoeoXzrqT7jlEFlW/0rEuMS9W8
MRZCvhpAat8yec3eBaXdQKrLGJWXIL8T8iCDKgsTdVT3OM9JOrRD7t5G0oRO
sZdD6mflWM7ewlv+Qt+vZA1/HJE6UYno3jHXXeGvddBftqvUckvK+VBAOddQ
DKdqnVDBJU0n3WXr90QugfKluYbRGllu18Kg6WH1YH86vo8tIVwHN+MrbHF2
NnMxBm2i4oxJPhMIOzN0uTp5C2pJLctirbIcRmw5UjVn9GULwabn2UjBEGQr
BphI18XxHClGplQ6kMbNhvgPycWzraAiXrBnrpw4EUB45AlN41859zUs4Dxq
g72Mb8xXJIMjnk1vepjKQ76btOEOrL/cuHjerMrZ9AhKmMhFWyXy8ff1KoLl
sHVXZNKZf2aKxLFFxoR0rnsfMfOb1slcEAwYx0tsyDWfqJPSb0unJImC7gB7
nu4lZf8JpW9L8QwjGMAAer6kNkLivzIZB9F29dcdqC5dCUyqb2MvINqTzpPc
NuT+ajfFkhKmvpLaBnCMe/H51tnbyQsozdbiEPgvFM5s0FOHBO5ryX63Err+
+cGorSqa+VWQ5wWVuxUccE1u6dold4d5Gpu2cZlcVnGacP687lejAtgKlJzZ
BF5MWvPh6FFQhNYHMMmwxTOi6QFbDXj95jsd7F3/yoowVRYiNTGIu1PJQyQV
JklFep+c2mde/z3lQx1isk2x7Q5M50+tv3UQYKL+bGqfDK/XldFr61XRHmhk
e9z9TbDVucKJV6cWq79oHRhbDMm0W6jMKIrj/JmTKFGcBjdaYuAno0MUbcst
bCuJ7onHxS59YeqwqKgGhZHQksAI0WNVmz7ZWmFRhiZe2cJnOY5DhlzElbuL
6pUUkxx/mUNwRrEqxdyw+DcdZ0sdK3ZjCMZxTFeTZ0nZA1ELpmobHY7GIH9K
tfKZ7Yro9O1lM04tu2v1OHD2ywmPD6iTSjzMAXVf0T/WH5udUHMys//a3sKK
cpksIxuderXdMW7Xdz9pyUYG0v6FE1dIqeqgi/VOd/5qa5RCNlcQEJ3/8sFG
AdqCtv8l8OjTr9Nq/Y872qhyAc2lKlmnriGtnoX33rFdY4mlDFKwhscjbnfk
xQBLRWnNzu5yiBPTXDnVRO4OZ/2lHNqe4k/YOI5xBLGzU5Y2Wc3tIpvaOGh9
YMFDiDkrc/PwZnPEtZ/QL9LwifViqsktLOTAq0G3lgQ+/t9dpJyykUW0p0BX
vCzmx8MJo1cVWYKiVPJsUb0FZKSs/otcBDJN6k1YfhzAuzOaIOuYNKrwI+ph
6uwdtgQ9FRQA7CSXcv/15AqEtAg4rHy36JiXcWS5dPnZtHKEr9zfCEJb6BAC
QgC4LPa0ujBlAPhvYoIkkY8lwP6YJkiH7De/TL+4Lq9qPx3XOzLh3kjR/FY+
shtL3nbrEopf/MlKaIzx5ynEbg7Ag3lVUvBYRLNT6g3WIWDp3PQ+rCsf/D8a
M1WOvY24o5mNTRs8uX1k2AP8rpmdwt+y8LfJK4AY/l3RIL0pC6hzGqfuVDi9
KrSacelHQwjznTM76TTkOQ6suCxgGSavld1gL8nYI3wQM3gCJrBFNl1Xva3X
IPfRU2eNOqcEmNQxJ47RWRheisXer88jXKcgHTvF2y/4456Psh433ILWtcb1
j0Lt/BxH5QfvGdkhICQY5N5gD8xcpAONITivU5G8kfQVIP+46JasA42IyYWG
Me0xooKVYfosJ0ZymLT4wc7RXCNJKE9AehE7RzBBqBLFzRBmAtyAHlDnWxZ7
9qPit65nv074udt5f/eFEqID6++nIY82yN9wdPiBc0GJpHQInhca6zD7D07n
a2HfgbHamNcM6NRChfF/zj/QX0raKFieQGX4zedowHzpBYvEAwSjTo1yJknY
gbRNms7MFO/lXf/xWId2fotwD1uW0yi5kBYP1BgFfMzE6m6iFi1/fJ6Qxb06
2HxHRP0MCIWs/142GImNL+4mcRMRHl15Bj/HIdVFG8hEzmtUwSR06UpP62eX
/ck2Yj20nmu6NcXIiQ3CWfpD/NmqSnKVyZLWducoCij34ighcDQs/iVXgcsY
Udj7Bjxe0XMy5fm8SngKdDMrQTzoZb1YHJlEPpenK96aVQ+RjVYJOiyRRdEn
CrHGMEZBgCsN2VfXgZqhXNwhWi6bSAJ6c+iQ9LOM/L12ZpfYaoBRHZ/tfSky
7rjS5ZndhrWTzEsBgkw6Qi8VRBt3dg/IxZi/JVyPxdHU+6c1/nUs5fW5z/42
fdTKppoqr8JrNn7RurZikUOaWoEvaVt/AhetDc+Fx1qzAzhgCtKrid6+6epH
yo+JrRMg2kuVQJTQyYUMRlzKQBnzlBt/p+mDfVcI35vpBL9kXeBT2igxGmLK
fEofAGFZ51Ttrtd1ZSH0UkUJ7W9c44ul+1kd0kIBep8bj/blZaMN5AI5XIRA
U6rIaYf4m8dus2CtOu+alMK91iXGWpMXVeCP2ZCMGIcKiJOxtlzjotELUcZ4
nq93jt7ouWwjcYAz6gqe7x/m2wWFDJLrqqLrogPQ/eH1h/fC4h9dEC/UQJI5
PmDMDmkfH0I8r/d/wLlfcrPgO4gh6XNVN9Q0V0Kil7AABTzfNUDmK4bI1C9P
97mxSfME8jYoVsO4FxtnfZzvEjOBzfAuAgMf8/XmX5NxwhRN7oTVJ0jofup7
f0Ymkr9HzC0uupA+yx9egmaK6jONf7iMDppSc9yObCpyQlV+5otEvr5/bsul
MvGIvzn7Uok+8KaQIfcaNndkWnj/d1kii2p2OmXFC0kctwzZBvqPMQl5OZkC
bTuotRdJImPEBMUxblDES43Zx1IhopxNIyZ8cMK8QeArz7/UVGQrHFWg0Dzz
OkWt5iyHg5fIIABXRxTA8ySPkt1ww32CD6NW2CXu0W1eusAVw6yHMDkQu4jA
L01896Yu2Ec6m0dfaexY5oXpuQtHMN0FrYzMJ8pCbpAfXE+V/985Kq7JT/kp
ifwUANwpRErQJmO++ATCrv0QF5kGJZu4iCU0uLeLBUTT0wJ2DNl+lMum/OxA
EVCG0TTOBoxjeuPFKLTo9KfS2Un1V9uGyXTOAdAqk7mVF5IPLXT5KQQfjTTG
6FshJncbVofp1Pqa038lS0iO+BJmU4ckPAPuPJD2tX+PbVTEtSv282iJJC4m
OleEk39XHJdbul1UnQHlXpVfH08MlMzrD7HRl0TxMqUStmyNpbHNx9M1SkpB
YqFZALcXEIN70+5/hvGLo9ihCRgjDEBLhyu5j1IomEdBLZzMI9xB5PLIFUpg
FDxeNsvVe4trulVejJeYCn8vbDG/r77vd+AJ+g4UxWttrf/s/L9Y+K4kf4U9
oGnIUsogX7sP3gPX463qxxQgn0LJ+eVUtZCgK5FWs7DLQ1Z5VjXQL39wgcGC
znxMYMLcabDrctJFxxjU0z/wY0WxNItBgi9PXJdv2MB+uNmP4GobMnL9LnQo
AHGqkJd/C3TH4CbdGCjtc1ijVIdjJogb++7BfD7UGqtJdIZ3yTATZScpbLo+
FPnCumOUSGCOKS0LrlZ7pBRu5hTB6rp7cKeDos5sSD19d/YbhB0LpHJwDjiy
bQVX0CDmVWBsE5NT59ehgHU8StDJTslHjCEK80br847+IsqBkmEUzwqq5OUZ
UwWsqQ6JBWKYzwp2NpuvJP9SfcMRMs6OW/Zr1wHCcp2jOxwRTufyIy2zv5+z
J6HbdbR1HXkKXCeWBVvql+Ki+BCjlV/NEJDManKc8jMFki/0WqNwmMNUmfP5
m0Jhtnrb+VNQrzP1vMz6uK7sBQAlTIkqP07EObn6DBraSPThsrPD4vFLMOfo
dne5kFOPMI7ahz3YncIxaWpO0pculcjpUyDOxvb2cuAHCudOm0KDvgffRuBZ
sLGMEbZ2FaxP6szbfsVhirKn2xEjkj7lC7N04cmDWQy2rkY4IXjP/JHbUU8s
jKAMkG2piIZRRLvPYNYAeU8NnQIqsj3qnN5fqtKCJ++xdn/fOm6OYBXK1rDu
H/b9ivW3orKwkxN4qhao1X161YtfoFg4K5+PstO+IUG+Q64Eul+H77hx7vNp
fCzJG5jqJuJIkfi+sYcnPqXQJRvKw/SxC0rDM/Sa54jgu781XRoqmwtRDdah
g4WIGQAZQoTbHugGMxab0S8gvEHuwNA6hjwh5bkqwdKOd7ycmxr3keKwHCJ+
rlyvmtyzobVVxjVF7BNO/lSd1Q0KWc04TlGsJce2pxQaMmclXytVaz7gaZ4S
wy1v4P65t/KSIrBasa6uaWTIGuQ24hpHCag2vqcmIGG7Fd0QYZ1uVqOmYeSY
/ZkTASGBKqx3rpxolAKi54bB/ih7UJcYr+Ef2RcYLi3AXrbwGB06aB6Sxmya
3HZB5nhSGVSlRJ5A8VjrLcTac2SuBx8t9AtphdH7ZMX08L4kH/+BKPNBIGge
VHIIHkAn9hNxqQaxzVhOrccX1vlJrYpLlgpmDVZ1dKyXXIGwJ+J9P6iC8ngk
Sduu1XPXiYsly8hbWr3W1A+uNoS/Xa5jhEp6BooMxg6nHadct6/UQH9L7M2v
vvubrbh+VaIWPIfqy/gvVH8CwEu4QlWkw10JsvnS5fd9U9gL/2YLHtH3qRpJ
roeXikumF3P259yFusifUqh+XgaRGAVsEF+y/+AwagpgktmxtDXySOIfwYwq
d6z3ccVVVU44EWt6BWJVBQ2D032MIriINFPQBE+fO7wU4bnnHhMwz/AR76wg
QWYqCPc7rlMSotVDNarUAFiQvyaDQvbWLj0fY3rImEh88By+XSEFEV+3Af2e
p1S3M1BrxzWeicQPz+HSAxrfTKuzGS4NJTTMc8gFQ6yyVv/yGXUjkaFcNc+m
tBW2WzLTzHYpXxMfgKlgZMltb5E7sCKMUPzPK1YXtaT6RedBeJoxMOObBVNX
Ql0fJ0LU0+zj+bmYH2Ni6JpmhFsIo+1ZJgjACxr8sa8HA9ddes/PM0FHOZhl
gbgUk1WuJmHkDHTI5G3E7nDm6ycJ5eI6rZEzTIBe6Bas1L3X2FCja4fOGDSn
Bi6OUJbNXTxr91jQrxVGijSSUIIIAvuWK/oNamKpCHm9CKGVan+NP0kWSViQ
4jzOlKIonQRuy/N/rQAqBXHI9INVb1ROeUPRUeNip0iU6DSF7obUDh+ExhDe
0PYRwHEIuRV74mQWnheIV8keNgWGuYp9GIFibKb/SGYU8/P33kCuwc4slT5o
6dSslZRdOXPYrNkMYpt+x6fZMcTXIOdzbpLG/N3kbS0dgL9jS3eLcWoU9xib
wsL82fdviFoi0Y2VvqNTEk+89btAstyPz0ajYVmGUFUIOeC3zbypJiz/CNel
yASsZb8VLLLZZ+MWyu7Em2Ef3CJilQeHOzhmD3GgvlREZupP7MU/NFPiPq0l
DV9l+4V+VhiHKp+LPwrQCq4WBHe3gBYHIDGQ4rtw+HfBeyBc3qqPJtQoHODK
xm3lMJESE2IriMb5EWEkm/VFqWxcYX3Ntrx1oP9vhr7/GUlv/pMp8o/zh+JD
cF+Rg4Cp3yq9w3TsMNd8bdy7CvGjNwRkR08P/ZtvRxZ0VMIXHDXzFLe/zP1z
3w+UiyUfOJrZF0IB7CunIyEYUJxW5O7mOppvNAr+xFRvjcTba82sMVvckPwO
Q/I58HdW3/5P5/W43pMRPmfNbDhKbZXqvyLjxsUrTL+bk9Mie8D3KGOmng0Z
6a4MenTMhnf2dR2LQHPkxEvV8m/AIbAvVkNOTnvpHCDXNSk/ND8p3S+R5yVW
GblPvtpJH0Dcj7EKHvUsD8uK4af0ISItwxbSt8mP6P2G+5ZgWvnT8nx9wfSu
olTywSxsRnlWT5QkzDvTLdHRGhd71YdNADBoYTpUtKFjd7j8dBdM9z6aY2ST
BBhl2Oau0pFhMnGxYsXQcjHmFvPWGH4WMYG9R90t03an8ptpk1SPM/n4Re/l
NLsbbxIL35Ikotcdx/nT/8bVwM3M1TMgdYFz4V2T0arYpoh0tHmqsQq23j5a
iQ8T9iwWeQRYdkYyhyAgMdX+nfDVp27Fjkhb9qVVN7qjtTqFJEi590AgZ2o1
ctVjgNFE2AzyZtzSViclqXwc2S+KE09+XiHTxHUaDGPTdi5bfEagmdpeHyfS
puBlu/rNxEfPVsefJ9UC+Y77a8jLwCVIV8YcfmoTgwIZ66HVCWAGDpEzYDgz
iJ2tlEB2HLNMWqdmaOjQ4bfjm7H5KuCdwTdvm3VvLIAHB9noedp425mMeOFE
9FlExieWxxpQWpVDJ63wYYe6l1eRA7oRMP3sbG7syxzlJXKlwW8KtwDknXaC
iOkE39F0s0NCNulJ9lS+u+wm87gOE5Kno0h1NImk9g/uRQRLcrX/Yhg4dVdP
g4OWXELU45v9ejBZLiF6makNHDBH8K8LXpyXR7toWrxSph9Uajd67JW2LZ1R
GzoleYLyUiqi4k/mzMUkXNIc5jdJ0rbSmoya1ipNPTqT1SuPwUGMHclN384Y
HNWEvTLS5I8UoypqvsyPHoCfdgnhAWDY0/5fNmTYzkwJfnzpt0pU/g5E2d80
UiFHMIjXPcnfow5WUKTi/tnzvwvrM4xxcNy8yv37SEo//p8CMrwUtL3Fus3d
QeiJy26ACHbBG++YQITyf+Lf1uRrY0/E0p/V75BfRZMFqXj4YG6ZsuUt1t2a
QJqMuz/h0uRFuObPCOD2+YT7q+tgOvzz3O7LbtzuOVCTDPhd5jpjtvZgayQu
bCHz+BJGyrlUcQ7rcjaOsuTinROXExjE4HvBWCwUJG79NB5gu0H+/OVD36rw
jnAZ+SDG2lyiiqJdaxCHg6ImxD6ukTFgReWlYj/SnyZ8YpdtnyzGJ5noDSfM
BfrCcAtEcJrXICEIX22DkDgcBoRDkgXs9uC9mU3MzUwBOcXy0u2IcMXF3Num
X4D/w4RSk0PthcOP94ZYaAiyR3Z7kGOSDgb7S8HLMj/9yy0XiPJerQpXT64e
vPnXEd+OKLOLCkThlXLJNIGfExui3zyJkZy+71FD+KgEb1fEown6JqugcP0p
NQ0v1BqaUfWvGd3tYrEuoeU0vk0DeCons5ca+Bnl5LgR5jtBw7mCY1OBVMIa
4Msl+7KUcTWz1jDJF/tsUuYVDnUVM+J4W9iZp73kK4DPdv+D/FD672PcAKbK
fG7oKNtAu4WOW8ptQlrS+3NM68xJTvV0m3+OLEpN7Du+WYpVk9qh66p/X6aK
kxklWTEY0dSTVfvz4VBucSDmosKpsbH5KJKtXFNJAeq5XfC+IhmUGiiOQWwV
NnfD0nsZlLPJ+5iyIq7R8mdDofaDvIz3oRnetZmnv/HM7e9raAMolR57IcOw
coKqhCEhe7e6KobJBgQ3sas6jCgFzsaGXmQnWECjvM0eXl+BmXgvHuXafdcb
Px6JDs5je6rDza1Hw4lhgTrHTYCQq5ooFqzlwbiMtKH0ann3hQoauDBAZYvc
W4CBNOqfS3vjbM+N9g74bU3bkWS701fhMVdYSGR4S1cgZ2h6KelbBot/ByGc
Uldgmr8fiyvsWdrozBxRqSv6WhcPh+fqd8FRtatkv/sYPv/vwfnx0fV4qqLX
cUKN+460QJ+46z25zeT26Cpbd9gX2t/MB/5eYbBh91vjjHERFAzboTv9Lzny
iUT/CaMo0P4tnigkMuG4r8TA+9kcipMz4s7I8n/XKzV9iATNZkKBHGasToVD
rzr8lE0nQ7K+W98fE0IloJL/kZ0juuMYomOvihYNZKyhJINHW8GObIHlgpxf
Ensyocp/LN9ZSX9oP6/P+NBIwreXj3r+HaLm1Jsa4wgzVXrVDmlUKMsoMtTF
5oxt7U7nVE825tjwC2j0xNlS84zRAb7FR+UqN3dbPL5q0rB7KZ3x3YVHLwFc
HxIZabMNso3v/Ot8ecHMsP2K4OlvHnBuJz2lGsWzre50sKtNiqU/72vJH+Dv
KxG4HOxQ1kn/RgeDUsdB84sVxrFf5QiYzPkz+Ps/3CAgI6zLuHjktnrU/9HE
jtQHALK1f763EK8mo0xj/CKF0hiVheO4v4XbkOJXbdEOvxnSmM79jXaFQXOy
qHGDPskPtbigzEL5pBDJQR+bjuQTNaxA3e1cMRhGd3xEDxT9NOEz6musgb5K
JBXqPu+pTFkMkU32CpH+V6vKQRhssD9dGhU301u1VpRMiIV/jjoP3AWAeVkr
ewfO1f0ZlnkgUpNYahL+6CXXkLSrY+ULyyd+FL0XoBVPv3p6xA0TGxJQA6cx
Bz2W32IFEvH3LkhZAsrxj8zs8qtfHpXU6tQb/qJBlWM8IzBcg26jfJ0mZFNV
VO7MP/q3IeCy1l9QM820I57UefS4nJB3Ul4KgRaoP79hLaYdHVlRWjQ8psqS
Dtp0Dd+5ASdYdjd4ztnZONwelvjD7U7o+NOs0tE1mNTLRyXD23JYfzx1Zqi4
daiVJyQ/olfxc6CAvQoX1KJF/UfAJsdgnn/5vaOFXXnEbJ2yvH8x6jFArkLO
nKBDdg8/7WMu7qTjGeMIjjle8P5iWOTFAQc1JVfqOjzFD9STy3m+d/MI4PYZ
YUj+iP8OgTvm+cF3GGDgech12s1CC9SNyF9lyt9r4pbrneuPdLOiANap/o9f
vEuTZhF8cR0AXW1RwsHHY/ee2OQOtOtRb1L+wpM1ZN2hgwyGk6jxZI75H8aV
sPTLlA6P2r0YY+ntj7QLSX6IVdrX18ZTtF65A1ZuMBiefmmHDxcJ1aJYVXXa
87QRrGEeiYo5ZIftMDpU7YuEpzA4IVxjGxSE2e6OOfFgcqcpqGkDk6dR649a
D0Pnb/W66w/Kh1hhxEdtff2OLSO80b8EafzKCx5DpEEPMRJIt2O6kdGuPT6i
E5Vj8j3PmNF7nr2qDYSAxZVFzBELvWdna7wbTqPK5StnZEIhe4aoM2GRaSHg
fiElNMNypSiBuJYUP2QNPnBZh+UE5NmeNwjTH+dFV6YlA0REOmBRr4pPti09
zLFhzI28aGbPDTADTkHVUs34h/l6yVSQWOyrbgMn2WhT7oNTqoAH307UtW5y
E1fxDUQm3D6V5C9Ub6XFVLDOxIkvO6XKyeLBIX1aLLihhWFlctyYwKiEp2Kq
mz9HUU2xiASBv2mGcx4QSc1xJ/eLZVHUIvHkWpg2ruIba+PfikaYo6uwET11
3hHdcRLCnNnFTt654CBQ0pjlVmW/U8HMemhD5xlQYUEl7QOwcIoBg9LFGUOV
O/APOZZM1Mky6NoHG30UIZZQLU/2F80tVSxBKhMKsBLNbIp/D4GKNlF4fbzM
z/huqW5tvF2lr99z8w7VtSR+yZ5sEGhloADLXojeJdO82pJ2+69X9iOWog0E
v7O7KPZU0hahTgPIfRViN5HObjvz7R38/Ei3H9ATrazs1TAL3UrUaO+bARm0
AG2/m6fwLPU1ODvlOhKF6sarBEWyTuf+PcZmQNUGjH+iPheAbjPbZrpqasPI
JdvFTVPyasjSfPuretJ+ETFzbh0Wv4rfYscxIidm17ttkxSUKUhJrJzqIECS
R7YL8L49/Xpe8uJwwOGm2QEh2kfhosp9ZbHeVJ1BMzcLMG+ZDlzGQODHY5QJ
5Tz15c6VJ2GdKz81JDc8f+PE8V1jyFUFm584RuW+JFlUFJOSM98NQR6+S4ai
CwioWVNiRGuCrLNt5X+oo/nBmMPJkcsfvL02cchuTqXw1QmSpvpJho+E1Zh2
rPNgr1IMMtOc94P1zSm6BuLRt9Pd0K5vFeur/0I2Mv/sZCIRpGRVOnpLXGtV
q6YY8pdP9YxZ5bua2fQT0/pUOJiDZVm15doXs1mrM5YdJveKzvHa+GLj90oT
byXTMFRLqg+AkuAvk5N8U76KimWwiV9WgD7wclWbN/JFzOmadlcSODHsuNKb
d9wvWjuwSWVceDIQ8mmWNDXgFRAT04E5DkdAvLV6kz84Lqp/8WtP/qQO+EuU
6XEGwKRBlJhDB09qSa2LkssDuVFQpNDMOfuzsE0Opsp2caKu8UmoBnKQrTD3
beyM48TcWydn5/ztUgjvXVF0hZcEai13KZaxhkdnStdHjGxjzqe/aYa8c/P0
vNm23kEZQ8hmEJuc1UHe0LXmORiZCbpwD1A9epTGDFHyvkf9O7VoaMnV6hBr
R77nh+D4rSjdTNtsXc7R247RSLKQtBuspplzKSefqHK911rbfjnzxjjA9/jB
nBa1prsMPs0aHsaf5ipzYLyN+NZ1elefwsr/aQn5gTk++gaWsPTsq0Z82B8h
IZwseYmCnVttEDk6B232yKkKYOtBSw3bAd+aVlBy68JPTZA83JPXNhLlBRC5
NHA7Ud/9CBkrlAzhxItTfIE04VTOSPD2iCqWNbsDKF4NY1eBVnc6KdzNmyOv
qeq6ZOyYFwh7N8K+yT0gmNB4+1d1yBU+ASc4GSbjStwD6P0L6o9vbtabRUi8
HmDrOF4ghDU7geflg6Z6vQt+zaWJWnMtXrNNq90ugIMljSCpNgb3EEb9lfgQ
yJIT+upgNN20PdLqIZGSCRc+Lh5vKaKMyBGZ60PzgmrH/EBvx4bgRFUSA/zZ
7+nSsF0z18J7eJKdjBgcf1CZsiC1ozHdsHpz2lzljsGjGmNdEStTFWJ+txkd
8HMReGM3EppCcIUOcgzVoLrYKM4dNHb+D6d/IUAEDF46pBX/0pQwL71Y+/+n
s8B8na1QYHj5vDQCTi54IsoSBRUo/VgbDfHjBgF1jygxiWAsGIy0yafeSdZO
dw1DbnVQZXZ1VTqE5lw4ZhSGLREVj6EGMAAXRsp5CKRfUF4HRqwlF02qoFxb
IgYdk3S2BrZEMrqFCqu1MDJVFydt/DW8PT4bSsxVeajFLGYoSbSt7taowLei
lh9KGSMGXetFgqW2NuJmoWSa0Tb/SOVA/OIStGVN1G4Eg2Ty5HtDwQiR+0ws
tUxDX02My3NDpZSS5COD2GO2XyxwTX+e87BDwXTD8eimSvXC7RlSPREdV7CJ
GY8AJU1qGIBwzhinrjvaVzAN/iG8ROfQ82nIRru0TMdnylpWxLsWNmiIqPTq
icIdDnUupeJZG/6vi8lXKkP1EgXjjRq50/lEVeiL/MoYpo5UIibs/sk1ljtd
DZg3vuF7nhhb7vav5Fk1ncaZ8sBvb/B6683Yj1MKpa8ePE+Jforo4mQ+JlN8
y9rOG0ZffaY8UxKqP1ng6qMXNUJCovK8349bLphjvNuj6ValHA/b3B2XC91/
ofnV+2SHskH52kiElyWpwvOmuUOr/iU6bQVXCHh2p0tQ08E+MNvup5lxo8bB
QSnLbhci1merGbyYe4r2gs9C00ZYGYpOv1TUwJf1jsf8MjpyrxT+BALYQjpP
cPLcmRc+BPbGGUvBhwNQhF02i7YKYUkkKoPUIF4TrGC4gGJqDl9EVHL2YI9g
fy/uoGgvK4rXVE3Y/7rdaPP9u5m4OtXjAwdvfMzA7yKHZWxLIsFYd2lDCuu6
s1sr95e9r++Dkm+5gxSQdBJUKwaYbKwsUhjQadbitVJD9a88WzI/z2cAEhoN
Rqe3o+IdEJU4VUFUiZ6Y8Jv9twb6S+bYAqwUCXVDM4DBZZ9lPiubdSL34HLu
c7N2hZ76jGLzJfMz4PKwrEMyyK6k9ScskouzxPxj0wuzoBHMhPs+rX91wYlJ
SNxfCQqPjr0zWoLYiIgA1CTI4zT6qR2IoUWmwAmdvYzr+bsaiq7TeN8v3gpq
SZNicjub2AMgIBHrXkb5T3+ZYUb68V5QaaXCm4DeP9NvfZ8O/uBrJoDUMEkF
RWpRyvrlocb/m9nuwK2CtO1r5M9/FHqz1U0a4v7WLHacGFccrAdP6p22ZIF+
Bl03I+xFXsw3RyUWF9Ck00CDmGlh5PvCCn/Pz3OYYmo1WP7m9tJlbYoKr49c
OHWY0LfPpxVGwsGyF612Y6+didFZrTZMSPjjxUOEYitQxaoLVEriSblh3HF4
3pVE0i8cqGT/I6OT9FjOiln+twfD/1ry0hv4NbcRAYy2t7LaOKN5dj/KVyyg
4knKLnUYv/WLv5U5FlasmLudByLk3kQSwhoOm0+f6bP+Fq0YtVXCUDvqJ3Qo
U47TN27MEvRzm2m5lwxLyILUVxe2g1YIXBJQ1s38lJjjmfuCJNGIhzTINLHc
CQPepvxN5mjom3gTORc/K9C9ZmxxA9Q6Qh/m3GuA0ocfR6jYkvpF59rdglBK
cHkVpNHEvLWif8u7grR4LaI1CDWBPlT52xGrpLoqybDsEbYz8P1OLvZZHRuR
QwGfMa/CxHKcVA1RVwkT/O/qGKkKhDbhSw1rw76UnRxYBBzDRi2Svysh96dy
HRRu53DcJmM9s0vOh+Y/I5xMb/lCTzUJZKT6nJiU+CT/tTCBX8rqqMMzLjaM
xKXNS6ylJi+ZpUz4IepVRX+PkO/UfDLFgJkGAi6FJDIPczQ2qjo39WUb2F5X
VnZf/TZX1P7HMhI2wfMIsq3qjq/IXGao8+AovzKp3cgHio63NOXv5JoZ3VJq
beqxnHZmig2hM2GLN3fnXRACWNBqNnqwccHRVrEUWSEuU/KnNOhQaUG5D2MV
RmiDwTBJQfNnLzVfa2wPmW7P9rNHVRsDZb9SNG7Ge+Yk0v+M8IAYm07uIxZ5
xSzVAPjkKr0YiNA4PWOgvel3lE7+Gmgu4NF3UWv6pGipca9EVyqE10xwFpWx
F9Js9d+mc+Jjn2mVhLspygm8qdSodiu7USmQbJ8Omf5g8WzhUZBxrKRb99wf
ItYD9ypnwspfzwAj+HKxw21APrrUgV6N6G/HMd8YyLqERlitOOc56cg6ftu3
Gmk7gOhNbGlm+4YJSTLuxOw3kPCT7xU6jCT9YQue4Inv8WlOMasByYA5etAo
+V+AFOkYkWkbG3CRM69U8qdJZNBtSsTWerwySrWvjqHC1pG07meyx5N1GDv3
SNPxPh+74toR6BkxvDT7Pd+xiq3WLtvuHli2e4Giaqsmt0t5PFxuLV73R8W8
ZNpcVZXtUKl1yivYxfExaNUxCwXAL2LivjVP0AFXcXlMoOqps2Y/L4GUhyCx
8eHXhudfyiwUVkJ+E8xwI6zF7my/r/jOvNzmX9MzsTiNAkAZ43aaR7q58TyO
VY/z3Mk5JRaF9CE4I7yXGAjAzgMFhPLO34GRJO7bycCJeEEV/c7ij/OMOJnO
m3EQI67a5MFchU/9ltkM32W2qFTPQ3RV8l59rbdgfNJdTGolDf8V+unOLi4U
EqqwqLGGxza6xn3ncB8kvQ6CH0F5H9KwqujPEVQsuILGSlP83VOAf6ZP8/bP
ajDiL9eXuvSJXtjqCr4n/PFcwlDwEEM5RjG7hAsjRWJ9MnrEbDZLSekNs8MF
eEpcG938lJVY4tMkr2mylhclX5FIR/KDr2Qx095mf5mUBJPU75SYl5Ya3GN7
nTb7kEw9uaCE+ljXJW1bLTTnn9Lw9fXj3+Is5bca5Q5I0rRHxYYLzmkI2Upn
VSCVh6jVcFr2ceuid0bzfzhxifOznwuPRctiufaGUsWlsV3LEuVF6ji57j/f
BuXzfn5/AF58p3TbbPyjbEwQnRzIB73tGzxB7S0u0AsaIRECEUkAjg7q+ROd
eg+bAT/B30UkNv+5lEeXDkoLhf90KFLb3/D3yP3JnXUU8gtl+BVTQzn4SnvO
k2DnrT8OmzQyLcUPPtNOMnMejFPKKnLUeARWsE8HEu3GaeUZUvgsJ3m1irSf
Y0b0oSqo0sFmmtD8wYmuYv+d5yWIDRMk1aFfMeVy2NcauNffPQNAyuj7I2n0
MRLAoVh6Bs3/YyqGl0nyoKl6JE7/VoVG2Q0IiUcgfXNHW6kesdrCR0K/E+BR
mGBa6Qw3WPRbt2vCBmid+bk6AQMrVqDDQRdfGRPK5AybAlpsnMM/3YoG0NFI
m+S7X+eDaNvs+3vPmFnIEqNiT30qiyV+Qpx1F6NF1/dq53OveCTFOq0ngK3W
Ndbime7KWarEOUX23XKv1Fr/Wol35UvRMjsqqWxzom+P0qEr2s0VN9h2oXzk
qi2iWV5OZgzcQjIJmLTj08ucurQJTaRhvo+tOjin059HbFcvxgwypnRFtWR+
XjM4/Wk9oR+jo//SDWZilCMMchPH05Ckxc6Jao/pYEJ1uhK6T/F5o3IrNeQi
QI6RiDsQHFW4xPV9QZxQWfLKnHPUdP9xYzZE9VpivjLsdbyGBvmtABwKo8h5
fUxx6/GdClyarZq3N1eTbD0SVY67IGS8BRceNsyRtkkt6rrxxdLt7C/DgC6F
Jfw172fQn1t+uCPwcgWwiCOdiz6+BVYJ5Rj4fGq4b/sjqo3op6DmONLxh9Al
NHmxit1i7xNIhGKRYbGFGW29+obtZYnikToInZOHYJZpCKHfrZhIJ2Dc7DpJ
jrWoRADbex2RJlq88eAQqobBJ2vs241gvCoX6pNk+sOZ49oPElvS1zV6LO0C
958NWV6zqVA43Fnt1HZbtEl8QCz741kMVblOfG5cs0mLGLmBTlB8u/1dQPEm
8lfpX6APRHwIiWjTk8W0yccTJVBGddc5IzGySf9xa2uNkdWqYY82Z2Fl1zFS
3uP53p+hQpBByy/C45OGCAxy2yVDtcRFDJVamLCWXujdh2MFaSWFzZGWDyhx
+KHUprCRUodMNKQ18S8KHvfF2+KoMD4Kk3drjm6IdyvBSjpT/z94I7tL62o8
C5kXaryOqqHMT1Z8/UaTLDHo+Ou2jvO9VwLJHHheWtdU7VnbcakHBCjKrWPh
EsAK3b/6vA6P8+P+Y9odvLO17CmWue7mkdgg/o2u5o9YDap7xkCXdal57+57
9GIuhWZjkqf8arOO2pkbmfdCl9IPkHvHyrOVf0u42yYVFf9AW588h80EfSxT
/H4wRM3x+ksO/ijQviQRCTsbluELO6t0c/kO5M58Wpl/jv0j4EG0CpxsTjhD
gd+j79k2AZILq+lJOVnGzNO8E6y2YLtgtkAwsali3tFdoIOGILZAKSfNAIeE
AZmwT+k4EpJ5SxWuuM2wwjAbODlkE9Y4EuC4Gd9Y0qvOY2UUtWYHVLdEb0KM
Tt6qU45nCV8mg0IaeMCpPjamf9rsMl/Sk0iIEb1QWLBk2bSgrl1cqt0wntX5
IgHdjeCVI2Bbacm50kHx3ZoM5P7rtJZNFRNiVbjh7XSyZ/K4jc/yFNXBO4DH
6mPuhJHARkalmNaBCPAEG49A4ur5g8tpBpNKgIWixEbbbnkTq0SBnXBKVQU+
IUBxgz+Qlv4So16diJ6V+TX19+n47wnBVK+ywrIIEdZecMFe836vshj6+pKG
svf1c7kOIjthu1utZEvZ+L1acieXc+Qdf+SsiIDc2i4qR7gjGbm9YuAidN6y
1YBtyBYB7kQE+W2XqNYSxNw+D2vVNzkoYaS8wEAlEmTea2hVDggptUC3UiRG
mD84pEJ4xxEinX6XXHE3i1YHNB8+xW2IPIOUHmGZHerO/GImmeWBd0yVZbNv
Zsnj6w3t4sxd5OMT8eV9J1obizWTlx137NWNNHOeyGhccav6PL5C8CS68kyT
L4QW7fjxLewWCcq++mmqpZIpAoC2TR/sAfdFMMubUKZ+LWcWegXMQ/soIRdy
etg7TxUYFVfkuB/zbF2c+VyDR0uddhBfwadHr/0j1UWSzfH6WF46uJiSMpmp
3kX7iR1/KGmQRd+thMsqaZEXEXOQn0jhuhPf5R8rJ7bbJwzWvdnXiClPKlW9
AleaCP+MzSLNTXZfIptOPbAPwdxeqthMaHYovIEm/cEL2fUlN0n4ielAToOq
tMUTvmO55jx+pOClcx7ilH1F8B7TRrL61Q10NwS9SCj8QPYjoMt5gL9VnREv
wQc6+8TpSrXY00L3Qz+iWX4xAub/4zQp34GYFSkF4MKd/uagrZG3NDkPRYHt
ZUxNfTg+5VHidtwIozkIV+PSLrdbbQfiHFx/6rNVV9O3YqtkQlBkPbh8iKAY
aYUvabmzad4OisaQOMG9HDU6gjyNauBQDVP12s3VqKwYVwUGZPCdXXlZkUVf
3JAqxTfM9ELjHKlYK6YUDHoorWVM/9PXyhythiI89n1k8H8X+vok2fFCIZ5/
Qc9eCwutsD5cdfBI4hS1HMUW22m+g186t0V2AAEfjSAMzr1MNYxSutm6uTPO
Eb9ula5OEmuseHGqZhMz2lXD8DzlX440Uno6HUb9qgu0frBncAxnFGZFFEIB
H849psG39dphaK12tELAha+Apkx8Bs0P7er2zsIuAXaS0uGUxriJXTdDRux9
apGPJyVs2PD7dvaUsYfQOnDu0tLeo2t/obzspwAgd7WTfjwkD0O15jcZd0OU
0xpxomxS7Rs5oDMX6eQLyP9aPK6wwtO+CbVltkFahGX0g5Pq3cHVTCVEbLtx
ecZQncOQ5seev4kiXYeZie5FDir5iA3LW/Xs5THnjAK3CEdnHAEWBkQO+S56
BNZ2mZHAQwslAVIFC4XpbVU4ZagsdjAP/lPm6LAFBf0MGjjIBlk5oHrX1h3A
cqKNiIhD6dPhgUrM/SrMFKarwKTMyuTPLK7CziGCCIrvdZiZYjS7hiXBRT4n
H4r+VXwCDCnoyQufCoeiBF36gq0ZwhLCHt6VaMRlB+IanjT5Rjt5ebkwsBNR
VoybA7yE4aTua8G3uDlzNegMY+yOx5O7EEHdg1gp5bqBQ32l5Hm4y6PAFtjE
yQSP64mNn6UbeidLG6usyv6Pju4a9Jzv/kf3pxtTJLT92KfqeD7YGh/4IpTK
c9d/ZiGtHXHwGeKeN60QF5GuF8ygWmOu+hcDv6Hbd8ahCxJTyRQl1Xb6YPve
hUbcp3kZ77h5OZRJu6vkMNkrttZrSDcd3mE0CUNimkmBD48R8yuZZSHy2uRi
NrEwmjbQCIvgqelRWxE324yqlyPg+xLl2xjlrgW5FoHvq7Ux8fbaYCZr8k20
b5WG9I+U5fLvFNS23P8gjKOL5ex5hEy3gWlNl/xLsxK8C6BV+1BZZRz6l6wX
SdF7o+D0MA/1+d0x/pWAfl6lpiL0n7BfJKMkxoNcbiitdrX2Ww4qetzpzdcw
k768FmQ/P9tIBY9A1RRGlK5+dzchRWiPd3FyoxrogxraZ4B+cKpJpDXmAy7I
T8U5Gj9OiVqAC2n7ju1OEFbSTwqSSusYvFflsqIDfG3eTvVejehF7t5Xb7uW
hw1i40yCJKE4sRLRLpa622wKOtK4vERbT7zq1oPVZlHvTkzJb7wHEmuX3G0m
Qh+mzpJr+8qWA2ztBwgKHmR8nnNsg5SvBP5HQURIcxMFw7VAKy28y9bAW2pf
uh60A1pRqlhLNHltSSkrD5WAY2cqEPi8tfDOxkZ+scHrjaYJeOQYw+1x6YQk
DMMAX3lEEowwo63AUuOINdNquRmc6y8t/0R86Ti/gizx11jFol+mg6Pk9oOs
rAhuc7LAF89n8WxGA8Cs2goy0b1YUygVyBQYxo3szSSWtQGi63JdnanA2c46
PqxdwoNXpniNFtyONfeOEkP/iy/5RBgLLz8sJJCSxSa1vQHD5NO5pLXpyyBP
KMGkdQnE1HMsMIhv3csMv7L/p2e8Lv+15ufZWcyrWKb+6VLoCnrfwNzmV7eA
fce8KmXT0l/IKzkcWxdH4ctAg8L+j11JL7uomNa5zNTIGRqRG9uexWVjF8KP
hhXxW2+2ktZv1KnznAzo/G3qWdL2UlxCPQBqnkx+HtEn3PprsuFc3jXGP+Ph
dJcfaBP7zRLv9luaOmZwxRK3ussDXtEYV8bDSd/VQGnjcJqYePUoSGeGlMV3
EHhAUpfpjP/wzgZaXZsLTxy/LDK3TTeVbhwRFVlTRHK7THlniP05GeRUeuZx
qel/ekVLxb3Pyc91pAMbmbJe2kTCfe93L6DKZ5YSC2B2Zryq4LI+14LUnS2y
pJQj/rOHnbsXtWhiCZiR4E/qPBNWIucX4Pkb1qnWsOxacPRoUUeeDXdMdvpM
47cYnka3Lup25FQtlgOw9lEJvUUgl9S/LLSNxuYGErYq8Uz3wG27F91Na+ch
EVmS/fI9+EK1vx6m6snnc+hwdijB7Qt75bWls7RjTZZJAfx0WMZ6j/07Uo8u
zYwA31eIRJcQ50zfLBnWxfXjPquBSk3LVuEq0+R5uSYIYW3HU40eclEvyztx
Wkzaoki3DmFeKXC50Wums1jLEljzovTvPJhqGhoZktnN/WNXZ2MC6Tk1xQKl
ghyG75m06YfMCU/bz4ZOErMyJe65dpR5LwA+zVzdULAjwb3SWAPF8QSxiK4t
cPkS0kmEuhshBpAkGvqLIHRy1+Jg0mcCINale6Dh/fqayPwOTaurwCA6aNlC
Jk/7c7IJw2kDjc7jouL1SiO1hasnaD3jtBqS7+w9SJ1RllQPzi19tXG0Sx1x
z6ETfkjhV7UWzHhn1pIwkBJ5VuoVet1sTALER7QUr8xkvaQl44zYAFTfnyTk
oNS/Pil4vzP7BgoEE1M5cksRFGPU4S5aVA+J1NAb0XWdMXZ4JgpMRgSBcCaV
mFormHQd6RDYeCGqKrQaD+cWo1jJGeEJz4PVu92x5ahh2A/pUi8NufUK8m4Y
JAmFl2nRJFflfsUZarLlkfuGzyPxplUj+fR3RdnOyOpUe02BI8aFTER9rvtN
qd9ef4hbaQsckeIsis3gOpDLIFLz3YsRkkGTduqbmXL4dd/l8W3snK7TnO5P
U8neBQXjiwvAxGVFZ45tEzARCD3q4NMYlfnrgVl7gntSsOar0lAFRF/smVo2
XpRyAynqcQRSfauLsNj0Gjn5jg5G+RWrXzcvyePhNB5QgUaGa2f1l4nZiJt/
o59OaNnTulCYQsmCAS58FiJmi1gJexgnqbst7v10FnXU9DRcPsWD3HeP8qk4
gcAvvVzOEWDm2bBR/SR0sfnD/KB4JBKCXduEix3GEzp/qEu8cmaL1XZF8Gqo
TnPh+NGRukl2lzcfHjFGhCOU/BjzpqRTIlRNIe3IVDGYbECY7umcNCmYZUHO
sdonm4CfODVm1c/gBxtHuOfORkddCzDFEzx3wdD8fSKP2Chb7Ia8fQTTd7ZA
6KQuQNBNdE7mgu5VFuIkdOThy5ttQaazLnT0zqfj60x6Nz0EAh/8o/qhXI3r
MGqCqieHoq/0wZAh/jcPhLlKeE91qsP00Wg6rgdMEaE7PlMqhwqS9r9o/gat
ORv/xMRhut3C1V8wpfwz5Ef2dH0d7nOBjUpGIR6lgoNfb0PcvCle3kID5RBd
cptyszOBmtAF9COSt023fG/ljpv8L1HSpkW3mCFMMbyOWfNRqccR8N48BW3D
KCI0nzbwJcf0V16x1WTq8O0WijC8Vj+o/Lez7h8TtVy438nGQqJe7yE5lacD
RO3IXKstlL6eiw6Lf190hDue1/Caf6VB2Kho2IqSM80eEU/nwDfzMiR2zQ0k
NL174nPBQUp7luWUIjP03kya+X5BlwzskBxJFPqmcOukowACH/UE4Qa9tyra
gF8xmbK7jVNCGCy7znC6VCCD+lH8OvkfKGx+oRITA00V/4Bq2RFD8jKfBYDE
f1UGvTKPh63snIvqad9EG0QBslu5gOUUkqN3CKtJfRYs1w8TL+wUiTRAEqhI
Kger9w8toY/IutbEnTZRn+/IGKwFFiscGWhls2f7+eYQYKt79gcpUdBhsDt3
WczzGidSjc8sEz4NwY0Bpm5UJGBa6Zzw7N+1mv+OkOndt0h0fE+GwF0ggj0C
2aHf6vQgqmitlmMgPZcQdNMQ/scAo06OUdZAzAv+eEtN2HMTCWIovqVZDcKa
V7lgBJy00b3GOd62hB+FGNQTuWk7sBXNDOA2GCl/RiMtQY62insFIc+WpDZ4
ig9oBGR+ccGC7CbqUQZ3NabCDbm8+DB4DpwPjGRsp+hwzmYR9+PDtjZC1NIQ
l13BXcI8n0xYHll4Uf5mouDa6O0FxeIwnR+Jyc09caRrU2b3Ag0KiK+Xtau2
cbRY7yz3hatb7s9QXdUXYr0Z3SQTnKMwgw4ozw1DcDzLhMeq3Ps8KFAd0Hdu
Y++Yur8zqsdQ26PixyUlwkzkUzNgEmsQWsnOgAWXC079ZulI1euc/pqksHgt
ZVW+inyPj/hA7Ge5FEq9H38mMv7NLalkFFGJpLImm0ohV+rLURDQkreksbwl
GJCv587sCP/wNLhfHwZaG8BpIkCMBXemofMfDRyZU5BIgmcdBwb6KesnVND4
Jtto2Hg5ecQ/RQKk9bR9ZcEFVeaLBDSEoRmU4yjqwoFwjqBn/RgJYIcXzevu
ITYugEJFqr2njb/hYmkbgA+HPeL05rB+BdO0nxAG2mxGnlBTdhuVl6ARS+Pe
SEHBKdHhZn9uE29me9boANMTpKvKJs7tCn1LW/Oz5AVpPzhIXCwKdp5Qa/DE
H4ELy85s69qj+rE/2jxA7Z8mYytdJX7NmepGAqR6dLzPfFx7fHO/NT3EYcsN
kKZTFOPq5CwHkv3XC12s3mNJs0uxd4LWDyUGRJo4FJajiiyVJqv5epDuJGqT
q0+AwR7z/FjjbPwPltzegyr+RAoQXLdGRZj2+jCu0pwyFdgXx76zqIGrVfyl
A4Jpt0DLn0CbYkhDJnEhGxsBpeZPKsa3HdUsEg3w6Zx3uVftO2Vs1zIHnpAD
0OjID6w5GZzR+Np+PXR+3QMBzJP7qWJ5vtEIsh+xJranv0gUBZ8wKl5jKfm8
Jfyf/O2qQLfWewDFTfs80SNZcb+vgo9jZMhhuuvQ953pyQsQ842+FjNNCJjv
Zn2oDfAotyrlCnfWDDAPvw5+8sWaiQtIH177VEvXRipmYVJCrBjsx4sOKhcx
fXVGiCwnbdAQC9SdiTXYZTrp2D9cWCu37VLiG5piyq98TFlTaNCFAIEQq5BJ
gUZI2s4zPsS+9YErNHq82MI6fTDNWr3gfB8b0ArhpOu3FHQms+iRvMsAX3Bu
EGOOmSuxyibQli3owfiEl21HIkBo/5o07yj2r9h0AYH+SQ/mZja1pQJjweUu
tD30BO1UU9rOS9X2R0HhMgWjaK/RVRSjJGIdmr8uNHNKZ1+HoE16nZy2fq1r
216DlN3U31IEekHPG9///E3mZNa0R9QTKp8Q1Rj8cCruLpFa139eE29DfRUo
sIz73FVwaZMkKRWTSF8tKbwuREytl+i9dzIMZ/z5TAGCVrFke0WvwcLcN6Rj
FLlQpFW2ViEUc5E7e/12rlR1kL+6mhGnw6PTaoMmXZWYoD08PXCcsxK8FMkv
tsJ34DWxaExMO4woIjpkTSBvqCrAA2KCA7Y8QFdMn5OlvINM9ppiYxkQCRDx
g3NOrEOlCTRKflJvghRjOoG37u1MBosR5m2Uognl/trcFGKwgRLOE9GnpCWg
gxaHrbA7gi1OBvn9KI9ejR6rWkIJYxRu+5I6L4eNoZ2YjBwkFKQv/WSon64Z
rwoYg7VHdq18Qx07l4OQDbGODOeCdQviVT7xQk/aDTHY+B0VIsOR4K9CmW6G
Z/j+nbHBrWQxqzJbZlmeFljfJhU95xw1tj2VH9V8rCUEapK6rSYaJ2girVEv
jYU53KoFqKjp3kHxvMUMaxr7qKebhQrWGOgfz8rYup7NY7ZFxHKWPiT3INvi
3ku4NJA5N/9p59S6Jpj+gUEiqicNpSeJch+uUls0H+oyNX3UE6+wUMMqGQ4M
yFgiVwNXHYBi6oevRI7eXmJxIyA06WprvSNEzxXbaXnpY4JdDQLQGDb03Ex9
oxDD1mH7tpAL7Qms2vX4J99aOMF8zSq5sPSF8XycXhjBmWOis+RiyD78Qzxb
qhCyN/p6KkC1H6Yw7tfqmVsxwqqzW+mFQhkDQ6+rRTFh7df518aPivxEHbnk
Xq5mroljaZtjieX8nax2PuTKM7KPLKx5JKdnEwh7SAX2qX9hM40rLPsal3QX
3iLyS8T2AhSzQgf7Z9rqiZypK7Zbe/XHMBMcvGWN8+tZrlNbWE0sO6/nHpnE
CMVJ36ZOG0ZYPXAGNytB3xSdwY3eylr5qxPMxAulwKhNVb1xsZr3OQoFtdIj
xcN5TelpcPmKZb3kyNcjhkEVN6UUKpbDxZT7dazeXAlfd4AkA9j9+/IgX1KF
GwuUh2WlNV/RUIFhu4ePzfftHnL9ckOMlTivdpsfdbzGSZGj6QC1ArM6kao8
9GS4zhB8jp2NiorWLSWswsMLjHVDekscrPwZXDDfVvV4pZcZE6WzvDIOasjg
3TpWsgqMvirwlAfzltB/eBuV9sZ95TqzlGo2ZWZSWpyfJPXEHY5RM3nO4ppY
kH3XF+XI9caEpeEiM1Q75sggL8iABVateku5B23RvUcBF82JCETGF+fz1Wkq
hZVCghzC79pYyO2JVRu7t60xKjwZvD95ZVJdPRPRRiSoHngPsLwIh5PFwV8Q
w9daRlRGAghtPoQ6ff85/ASWIIbmkHnPdp3b2waFGI8EuQf5cOcDkAv5JJwn
H/XjgJ84EkJ1TLqWlMdYbKAOsr0lQ562rjJ643g45Q42z62MuNxRfT+KpQfa
WuoPP1heLZuP7R2abMsbAOAJ6Rss2i+Q+4Co+ExjMLmQblHw7bL3QTkohkZg
+2qZ4NbzUcy0FN3gcODc7PmoqmtkuEWE/yIR3mfy5ajZ/KokSQ7M+YNf94s8
uEfmJzaWlr6H8Z9H/tlZQXBr/+VNxprQCKNSgvFiiUj/eNeN3rG1n/xk8tWs
S0Z4DwXMbkMUdisWpbDWY4N7tLnrV0O6zrfhZoPiuNwoic+lwt5RL+vH1PBn
LzVw8S6Lv/FgF4ZpQdppZtP8C6IUxwZi7JS+HqSsRR0UXnVLQVZ3TyFBVoDe
owK66BkdN48U+BIkGmLuCSNB9Rwfy27rMhdPy+9OjT5rAdINkt0KEQ6Ctnl4
4M7+3ukQoY55KpJArvJ+VdgHMlIx2ZBN63EAQ+DM2MbsfTDEEcLDUw/5zg3F
WOWIqFKh/mB1qDlsMLo5MvLBkhz+scwLXW1v6icsczEgWwJm4TdCyYkz/C7c
VmpLKnWs5RxUzLpMBjajHYImlmZnFfqxjZUGzBibz++a0PF2Hy0A3u7RKdSv
+8Smhrs0a2jYNvSEA2bU8XLn8IdSfIkBsFoNWZlOnPBiSF18lxhSfWgivZ5U
TXb62dPkFQExrkO7bhYTmMxwqD/3b6o2rVCcrzLnDgY05f3pBHgLJPv4ZE2T
EgTlGznYjCxFJJcxv6Yc2AeKNF3OrNZQOV+T3kmtxUZ5WyxwaUPqhxXfz/Z5
nvhx8tvzAENY0eikrHhI16OJyfVXBIrIqRG/EA/+1UVKl5RdBXmx+/mO0hTY
KKIJPnf0L6+RPSyyN3GXiCImB6tJKPkvoo+c2DjckpZDWprpXf62SH3Kpknx
/gcI7yPQBJZsxVrxt36423MNYPjqYiYmyT3Nr6gyAznkdHmG/RN3NjYMrb1V
R9iNFYj2p3IZ1Fb4MTO9dE6PCCI8TvYsRALTm7q8saKOUldmALWwWbkR35lI
QjKm8AbSclEMSbj3YGmQ/MGszPFRo2caNB7sfujxCV/b57GmOGcDuMqxrFHL
2HwPt4TJoDTWLtgC3EuVf0bRhb7RlezqCt5clObk1V5VHHqSXb5Jfn3i64aN
rE4P6nW3KOeiDbC173kFFsfWVben+yEmlPLXTSGCxsMDOXy4Z6gR11PQjbVT
zDtZAyNjvMFUj4e5yzJcrsmlYXamJyC8jkyDZIChbA+CER6+QuvS6H8+99pX
8KJqqK+ZbVC5SmpBHchr4Zh15BG92ByHh2N0X+di3pRkWYUoLYGZmqi4kmWJ
XnYxPvj7MY0AXtr6zrHmTWojbHRrtxyPjjJhrjTsT5MRzdqmX0nrTl2oASeG
7q8PnhSOw3wfCnTUgfukzCIGBKUz2HBl1LfsqadiSoetNJmpwY8iSCQgzGAP
0kVmEp+RrRT3KZ2GXkvH2Jr6oDtr3xDP+l6GoSlEHrzNXU41oPd20lFR8md1
05AWOIuxqkfH5j/drIFDrQqNjECU56/0CbC9EdQnfcOPXsduvvYrMorkPQJ0
hUfVYmApbjOie6hxfFJpHpzHgtJoOVRtCUnV7wUOa3YrNrUhgyvn/V+vq97Z
LqBRS5vzHsNmkK5VrCku3uK9+tD3Gw6Cz5CkL/rLnCfuZodxWcQSu2c2NCgj
ZH9H76DKMv5RqgIDkeD00tE7W2y9RE6ATHB1dLwFIziLXsFTJTu02RfpjytH
OaIlpIYV9n5GqC4wcdT4mQvitFlEdcJScyS6yt+xYKeo2j+20R41rObOBd3G
evBzzueRtq3yN6+72zeUbHX4sJ3tqPu2sotVdJzu9bhEDlEjhXBKqCivCpHd
V7/EmMzg9dUSfs4W/znhItq3gUR6ofBxw8IHlX5RhFdqSMiOGF+BWdhSLCYl
Fout+xaVmvpuk5rAI6ZOBhZ7aB24CzgDgokY2ptxnjuSFK9UQmQ46v8BZIf2
gj4huIM0TgnMZvN8ZbRDwO3JzipmpMXYWvrXRhJLmANf4eYViy5+IjNePkNh
SYeu6qqOWWedmBo4RfyvHo8ZAD6kCrSuSk0RuCpUSK9ecf3iNU6hHuAYohsp
YAnBbvNydE2WIsa+Fxu8UCQfOA/rhRb/xJfnhRORfWF/2zBW80QYmuZTFQA5
oyWS5UJ4zndR3jOZxNAsmiRkWEYix06gYw45nmyFZ45oVxMzNKxTZk7Rh4gO
B5uKfERyyP8JZxio/SfuBliNEjLt0sE1M3yzKLhDrV2VJaDh3mGR7NUHlVbF
oM+t0EzVuz94EaMSCSiFoG6GwhVAYTbgqWf6vKiGE/plKsw+gYj2m1GuZF2E
inzHGHuceDVNg41DAqGjE+87NpkQroPBXiCCzDvfK+2LmTBklO/20TjgMPcK
0FtkDXv5OIUk9Ylsxohj7CU6FHlVawcM7S/Bn2kqGWtGPNpIAWjoGTGTQk6v
mjuT0oc6Pnwd0C2SmGS2bvMphfsDUg60yEAW6A5gMHGB2jOQcTaN9W3Cc/0x
Vn62qX7hNbR03WANmFGS+FsUVXiEZ4E+n1OBya8xKCmGmkwFn+8DPFwDMkDN
lZxKrTJfpkGzVYQRuDUQQDtMC5UXwHJPmNdRfiSVJr55hHZ9kOwwkVQ4S3k6
YiTbgrK2ZhqmR2OzE+3RhzeWawR/12joEI49PS/zhl7APe/ABdEKV0Cis9mS
Ve+xzM+/qFouA1uB2I91twzPZJN7ZjPf29GZ566MUorgWRMCG8rRZInwb7DF
/I38Z2DP7oa1XE4KlT562CgrG0/1IV+hfgmv+GlxOMcsPGxu8yikHBRwDOs5
dEPyT57bSFL9HEOXCjpj/hv0vcEV78N2LWWf7zXoa3oT/1swDJSKAsHaC4Gl
5+7pNTR4rpCqKObLszwYHTUPySfhLthF/B+FQsWPoNrMdg9xR+FWvZekmghH
JIDCA02cwi9NXb4cNHD49szhxuVhmRhG+Sy6hrrWjkHJyvW8ZNzx4DaWcLUo
F5AxEh2VRFtMZMaA7w7OKia/vQ3dzMxO1t2pAfg/CEwoTWrpWalzAhaEsKUs
Q1rGHCxvk3Db5xgyiIZfOWV2KaFo+EnxcOOElUSXDlA/aFq7Mq3lDDWksz0O
vBiRme/Bn+fMj1Y6cWOKqZYV7oyl2S/EHYPq5YCISP7efOkSMUMSPqwK8rYe
9JAV3G1uMTuvSnA0uHj4GQ35Bgo4gj4sAMHrW35nSPN0dKodP2OZ6c8+WvAu
cfRyCyhJt7H2KgIEMWX2FLDXaQ3ChliF7Hc6BAxn2KxDWfybqq44tlvj8AV8
X/Bg7HerNTp1mwwqLGx1F/dw0ssRK3HvKgRkgvuPDkNsyPUsnvSjtZv3yUdR
KObcaranNDNxfDfut/vb9Aya4S22x+v8JeZGFyiW1NmJGXYdoFUeha9Tgtoz
nY+sty9DEonD7XD6G7bP8FGNS3MA4sKsRGdKTQhJCNvlRprm9Q28mikWDN9J
hwDlyijFT0DRq9Bma6cmSxjIYdhJc18C2GZazt3b5QhiZ9Z+H3ADCPQFKYOm
pne6I8AlSH0Es4LsygLUDxzzhE1/XkmGyu8ApBpKju5AmdGo4rgFtUW8xUQV
/tcpIAvETfMTQ/c32V6iIKiIBC2mSM1SmQMUgxPHyq914z5v7+Ik7tCc8+Wp
QBn/RDt9TJSTOQ5z9vnMwKqDU1pza3p/jTU6YlwHfswG73rYf+YPmfx7zNW8
QEQrwjGnj6jWVMn+GYeB/DQHhOfsCJvZnGEJxZcGhMT/IEwZdqXW3V9WfjUY
+Gg1GtryVaxtuG0T4TCdj139l6r/ZCiLHdYY1AyKEDAegfhpBzBMCS/WMycp
QtV6JjzLSEoezjS9ShxWn87moNFU3MOdek+VQqpSFpWD5UlySsXwYQe5AK02
1Fmwsul84bVJry61AZEuOTHChCtvTP68yArzTcSlxJfd01aQ6GcK1RZ3DJAX
C5k1JtWne1bS650iuWvZE/NS5ZZKwc74cZR3gqYnggwtyAd8R7BUFwzigCBS
6+UQM8MlekcSBCdPuQUMF/JR3cWmdYlASr3QFGlBkbopx4vI4ZDW0ORmDfAf
PKcM3UcvdaHLUr//YXPD/HKnEgTYrhcwJpa/U1JcJRYCkx9Qo5+FjjvUn6A8
4dqH9WizlZt+SD5Jr/T06DaCNlFcgQjr3j083/l9vKj7n+hiT431HtpPjNLP
lpLYzDtO1wHTFA4W4PWeI3bYSpnpUkfJBMv6GI4kwehg0CxNdSW8ZfDNr1er
7MaI5LJG5v2817PdEmnIE4G4MrfNu+S+8R4E23F4symY3bm6GYDeG4ebQCex
wMPsZR8XaiYNM2HTtzGXC7uzS4ZE1nDTtBfNe7wSR9BjbAUeqE5UcLv/pcWL
5cerd2sfMVw/DTh1jU4G5epiWgP/2ijSg4UGKq9wJtHpP5f73Y6IRsr9bwCD
uggx8SO53TUDmv+PxAfGslexS5NTXCToQitYaIHQ1i3yfHPRsYHz5PXRHWVt
z64U2qUWXzwh4e0E/0Zynk4/shVjv97wlPMCn1tUrPYTNUwncoGB47aeEvbE
xKns3gMvfgBFla8HY0vHzxOIby/bm1gBBzaxR86ZMNNxL23RNeBDxRaDloB6
UdzRd+4co3KZ8cz190B/kt9Cg/EisN/OfXc7G8dBHFeC9jejy4Y5c6XZB7bJ
+aXkb0PLECkEF/8FsbDL7fctTCOVjdDiljuONfUE2qDSVX0bAj1PY/D31YMJ
rWVSOb6So/mhYoG8GdaOom4xdBzSbJ31QO24cTG4CCc5yHP+DEfuFJO2nOe0
P76VPvnf92CG4Ai7ZjQKuZ7/shMlko04duUGyRvdJl6hT3f5gkQz6SuxXPxE
H/yAimq7p97KDFI9k1VMy38E5kvVy5A+4qY1xrr9s7xMxVYxpERQKz/0fJ64
bfuTs5A4IeTpHdPnAbh/fiickMKl9sSzAtDgYwsurSgfrYzQMg62dU9P4zH3
RGHjS/snYah+kvSmWUla3QA52dc/NRW0u/mJ5m3Gbdzv/4aAbPbElsQolr8D
MH/PVD1bOz07h8lgkVSb/wUCj3LYJKVtxNQG/cKy2R6zLsOqtvtpm8F5B2md
0hb0YK5kVd5CU78kAhxvFLQah4Vryh0nI0FQALYbJQEU4pViUJJWU99tZKmX
YauJZWUX2KMLxNJbXqILw9Tjn7ZALFTWf96zDd9gJESpS+2SHvhx7jUPkoDM
E8iZyJvwsF6mgk3IsEL177JXCs6H/AF1THTHGPpOo8o4YIshgsb3ZqFdsRwX
hzfPxmvPZpqnn8uP5Y3A4pYfNRrlj9SNvelLPCPZrfHV4JhBnEa3IBipUDZE
TXtpTqbs5Mg/Y9GqBUme7iGffHWP3A6cMxVWi1mfZapRbPI1mBaUSwfauqEl
L10pCzLcWmJ0oBp5Vx5x+WDMW9aH24RQwsSnEPMFO2HkVeawAI88v+HSSLgb
tZoozgeMuVphOJH4r+tHIFwT/rW3fJDSKKLgWsf4ZkviDqZPgShfN2gAmkH9
Q5Vbk5rTc1ZFUL0cOi6Q5B9DyEWKwUdtq7oIrDD+eHgApaMbMxLCA6t3gqaY
QjeIrWk/hW5xy8acyfomSbU6rdkY8DNJ8scwSApO00+Ei4EhbopN5QGwUQ61
/KPV4kDptBZk602jlKjHGh9shs1INYbMd/LJhsUKsZFmO67xIcZS7bRk2ZnS
91xMM2ehToDh+S/X4GI1sD/lCabNTFPQCKtZqUNTpXUauVOlZsCZt1kVfKMf
EjUHbJns2aVKjhJ3mnsc8zqgzxS7Vf74EHefkhNBz/x4Neo8lvuvGoAjdqQi
uAQOIGvuiLvPJM2lO913OSvevmgSkpG7rDnUpyuresNoIk0SfMGJVz09Ye/T
EfrgHTTdJkxiOqBHmGk4XFvJFyhlmnw4Z3o9garSSUAlaVd1ICXldqPkssho
YUnExe/IocnX8yajTdUB37HoQ2iy7qcvPSvD5Ub/koO0uqS3zEW+o5XgHsXn
cqK+yXfKgqKyPjQ2BaHn8TMRnqqbeq7H8k+2VDxMwTruKVMt43exoqBt/Kuh
A4FkcN6x7MXfIvIM4WILzb0e6m0fh92smnJdpnFCdSUAB1OfaApvxuO9A66b
mjtK5qaWKGVSKcg8rsbZ3EXKpePP5kYjQ+B6lR1Hwg+0/ETAqu8p4oE4jjvQ
/x54qlNWwnUMdgGwix9hG0wtZF9wgGzNc42/bPZOV1P5Dj+F1WeNqK+kmc1Z
cQTCvzli7/z1iUCZA6AQnNhqMa/wvg3VQg59YdcFwFe14eH4zblSTPw1hbq9
Y/OO3sb3Z92u2PRdx8QI4Ev75vX8aToY369qmSn3uy4igooLk1eCatSVatCx
6WgfGqfAxFg53ygSr+giyeii+Yat5Gma+rAr74FnZ3cjVmKeYuDH7+W7q7V4
V47P3WyqQBfeBif1DgfmRLDsDivjPMHNzPY3sluZ3zqL40YKm7f0qL/RiSBP
bPiwIt2XV4bLTye0iLwjMKp08FPZGW9wgqBSDUGfsANF67xe7utLmC7326kN
pEq7jOCpdOBkRBm3hB8gjNdSbjpED3fnNK/79yZJM/fcS58Bn13WVHBLfbTy
dQeC6YFLlq+URDCZtxEERsp36QCJlj2NhEnn9O2PtegYQMxdI4MihJJISCbt
3Gfd56O3XV/wtP3wN+3jE9VzmNfIsWzyQXJdofZaZZ7zfwBnXVLSnVmkaggx
UKNibtkBhitFh05pVV0slPBSXSD2uoN+0oGPtJiIoLVlDCVNBzaJhccYAl/n
yBp6Ask3Z9eVDCYoTHW/KU0eKRw3F8iP93zws4DOdgUkBN2prjmOoCvcXNj/
shhyCWrNTnjRXODUgvMrgHZyoMpN2AemPy0A/oSFubtpul23Np05vl+WNz94
pKJfnxxoPAs8bBvcMl1L7pmTIOr9eZwBQnCRgo5tf1xj9y88dAvMvpAI3Mge
475iiiCKQGJm/m9tsDPy2887b1/6Cl2sCvY1lC0alU4lkhHZaX8M4iy89E2O
v0kB4ZBSm5qJvGoHud93m9L/7C2e4GFrOzVI5k+0wm0gksMcdGvHmLCzGQml
QUvbVjkVa+cqbjS42Yun29dXNig5Wm8WSFvzf4rzP/uX83Uox6RKSMC9im5b
6CMjBjuWsnc2AD6VkZtlUjMH7bnfIpciDoCoGZvZgDPJGSQh0wxkQyVyiE06
92cN2zdC4F4SepLRqKoEvfOLMMt7Lt8CxCe4qqA4PQ7bPocbCtLQC/39ZSpV
XfhlkxGq3nZIeMeHIw9Owt14SlgvT9zJqY1VTu8JcUt+B2955AstcU4ldrQE
OMMtCtY8oNJhQh7u2TgLNJvUwcNUVQMm/XeICBywqDk08tzI1KpTKUiAj1vw
iao+na0CoPSebGYktthe7c38R8kBCIUtai+TSZn+f2/aFdiBjZqDH5KHIxoQ
fVHD+HJ6odTqIjg/Pnz7q0s6ZAPLrwtGe61pF8SRLDfxYYQyjOdxdLGfgMmB
sTUa9L6avlq1Pxgh5SvbcqAH8+HYm6SKVuHiBG0NmZroda7sr6pRMN96/dfp
u0P4O73cBfmtGQrL5gPKtAKP5Q8evv9xTm5jEobG87VhlwjeE3zBCpUr8Jvi
fLih0Drk0sizgizDWqlCF5eVdKNO1f/s2pxlpkumb//+sYOdOHYIdOOl/tTH
BZwOhRIuA01tCXmrbktyFDu4MG50avoLrdv34rxFf+6T0R1dPJAA3Y5ruW8/
PLE8TJMrTfc5LCcVO/6h4uHpirLYqvMIgMfZegLA2zzw+CH9pnkFix58ZnF6
ghijUSmioy7y9pfiRmxU/yrSGfqf8JjovNEs7T0BUQ8cFPky4SSScOC5eRQu
0+pzqEksiSjCLKhM3JKqcnG1Hi592Bddpu0tDSz0f7UYX9AutqOHFRkFdELY
dEqfwhDhu7q2MM74ntCkMfqGGygNO/RORcIadnWYhKmJIbQHe3fuPdw1nDt+
7qnXidV6vak3YtQQN0tkUkIUQ6m7NW9q6lFqxdvHq/c6srUrV/iku9B1IpBh
oEpBSrWoAh6RtLn8uTCrlFGNvwMwpjBCp681QJiPJQzyln2Du77FpK8xD066
IQHTGUDTtCQKZsr4mqn6eBi9MMkrnAN7iISst2wPKygWy6ycej9AdCerrwFX
PV/U2Y1q34/Lk65GdsoSFepudH3viK7bf7bi4tRQ7d07UknW1Xf4TRdOL6iq
sgpd+IjovcsaxI/SirQ+9mqa6ZcJ5ncuFkk6JHMIsvP/SRMj+HhulGpZa3qc
/4KddGIOoGs4ze+KMBf+ZytrLHfNoUNWkbHCJqvVyZfzqY25cddWAg/TT2NR
m80linRiXmwm3km7CTEAq5ikxUuWkT8ZvGFE/KXH4rZRvhBQMpPWIjv2HZTB
2iX71Dt9jR5MQTqWcOjH+y5Vm0VaesT2trHXtJs/znrrlbSkV2w0CTQwIaQv
3f10zIf1m29WcU0T6gkTSi37A93FZQgXWD6LTCEeYc/oEBbm6r5+pzqo3qFb
dPbgU8UsFlm7/8AdNGDTshLKLBVCfNxuxIrsCrF3SKj+0NVbkGC6SibgC7gc
G69Lz60ivNbsvZGdXX0V+qirCibP7GYGMupalfyh/dqt+Fl8AxwxxfXL+6gR
AlesppFN/fsr/az9RPhoR+OuseASqY+Qf+F1wfT2gC72+Ktd4T4PDK8zC7Ez
qG5UQwDG6jcoW5a0hckDU7X9PIUTH2DSgtAw9WlH4WErq4qoPf+wrEdh3LGL
ffwfWG8Zq8SZHNVz4kSCyIfp13jNfC3YyLr0G5UgSyXToPbOh7dIiuTzphZh
nqEeHFyij6RzWpnIt0LHVffnsycbkkYh51GuYK4YUeTBzGfPKnIV0+3DTdIU
qSKyc7K1xpgIzBI1PImMd5GUP22z9RBU+uQ8MwBAghAiOBlTuTMXzsKlmqgD
t9XpoCKpP5V9Npvn8R0yKnvmrlwfHox9E9eF16pCOPznIdsxOY4XHD3SPy5d
ckCnC8Y+p3rUEKlPegY75cGRH7VN4Wa9FUgAJeXsTNUSPxEm/EvZbQTLAZvW
EYc0T4Zs9+tddWxBM7FY/ykXO1f4eMtQI3F5gChQOp1ex1Z6KqzDUWcsT7hm
acso8ieZVY1/R3EtEYvB4KbWo3fH1/YqXdgeMc9hkgy+E5+NleEWOkJQsS7a
HhfFOqHDacQeCoSvEXel5rkuP3Ssxll6E+/mtC6R+wGvQPvAaLIwD/Ar9p+C
Mf+t+UfsFdT+YBa86vGqlXdce0ehaSZIwgpuR6Sd4BNIER+jD7Npm4ZqWBBX
TnrWBVeGhOizdmzyWLvygHvt6VFL9Gf/DYX6UtK7H7SgDXkq95F3sKhGx7LY
Oihhp0Bs+/BPMtQXeiYwblAHOR1bl9bmzR1OGnHHH7eDPeo+a0KZm2DI1Q62
kbwwzm9nC3Lq532NwZalR1dUrOsN1AE/MIxlNYUUKA707cOi64OvWB1LORzy
OtOfotgWavo83BKysrZp1pCrSOUZ2jJzH4B36pDmheHRPpKnVpVyeR5hi7Dx
WaqiZf8DE2Ao9CbjS1TiVc6y5BCvlreSrEllF9jTCZrZ0Z3VNnDnmX5w22a4
snFG+WylfogOJrxzG/GbEdG0sB3mYqcICUa194DkjZXUCWjzg6dFFr3oTTOx
8wH4dBsZsJuaPMT0HR4ciOW8iRcxdGV23OIY0Rfa4s6wVoaudQdf5bvAqJXo
/wVE2oTCkn7XjeH/z+GY58EImXBWOMRM1ljsXRJMnkBiUHc4e6GYCfoWFUsc
GEWrw648ASa4S1RyszUT5oWFj3Z/IK9qRe5cUU6tD+/VKih2jzEabwqv2YxQ
pHgf5+0qZRmh1gWS/eBjh+dKVCiB2WvPBCjNcBVUOQOcKNY9Rggow3kkaSD2
kvtymmPwrg+I4i0KUN1NO1NuUyH9ZdZrpBiIg+0Y4qDotpLnCOz8zL6BzN7m
cWNjROyC1pPi0jopX5P7iWNDBItelwTAuKmJxucQChnmI0ChTrxmNTDg3IMd
gECwEoVKrASozki1jBYB+ZjKwv3bWEW/fSqRGeDSKSKDeLHGscYlOHxjHuNn
tkIq8m05Neq9+YRQhfL0sbLyrGOr1I4a23cHrZT1TXcbSvGoC72QB/XAFaCK
Q6kL65/W2FNWRhsC/MOEDj0kQkMzrII6vXpULCa7gNwx+Obe8PM/3kkPoXgW
eJoXfA/zAu3vmfybl8DXtLTfD+1e+mL5qkmgx2GGsdHjU7YyhLZI4Lbd6EfG
JO9K0mSCI71hB6gEK1c33wcMxcz6jeTFu17pIl5pZk1PJ6NdpcJ9racZykp+
b489C1o7Ry2IxyFfyNbYXFYOvlAtLu6zjJtNMaF/zQecZbjZHVywACS3ceqC
jN/QSHtlnHazfqdPPyIaljGRwyfNBg82SYjTY0pschR2BpHTvLGtlUnlZG24
MwofUWrDUnMO3HC7khA2HlSwMdMvsAgft5xxNpm3sJoCI7l9ZBTvp2iM+7hf
Vo/zQ9RAfJfOIzov8g7asoVX6it+CkAvlvJ7QVvTIvPqIBR/Nn1uxsevOcbF
JNTcldt8L+Vw4lPs4puUW38x/ht4tNY0NCme7OsEH88Fsm3qh2U2kPE3EDK8
rwwylxYf9W1kTzDF5TEat88rRjMdIqRoDlcK0CgVg0IMpHVXto3mMJpx/cY8
PvUpg5qpRJRsem7SxRk+mofIx0sNADderUjIKfpa6nwJ4TMJdGzI7yM8CbvW
fWDliuZsdBHAW6V/V9Vb+TJ5H/mujDW8rnlF02Kying7MZ4Qs84a1ecexh2q
sAf4klP/Fkn5KhkrOu5y84woKN0U4qGaWgSvK9kOCIV58l7EQ/SJN2RXRxGr
6rN+c7eKeoKfOWRkxQoaNb6ltL/AailHvd+VnZR5eE/LgIA0nUD3XQxE1KUP
oMg+0DRDRqmqeaJMTQCfM8c+drQzynNK1B78L8Qat792LAkrpBH5yxq5PNao
1FzOIzS2Cy8N1mHKhDJW74ssaSiKtiToo0aPCHHgMyuRiQ+3lp+ODYxAJlb7
RymZ4tlOMegvqbFiZmCMkm4J8ZAmuztF0LNdrUSCUD/9hXiBzxLCy4SLoo19
fRfv0xiRGF9IxlSnaC23btJgBZGzq4vXJLhjtRzxIqgYyUngWd2Pa1BTZpZc
3fOWzSUSy2SZzTprmxGTzqhEc1vKI8EQDB2FFaOdpXlRvT6breUdHgLEgqgN
NaJu9q9gE8OwvTqA/nLZNwAeCmR/wj76SWGBkpTHhQ/XFFplQ3v0fnc8EN9Z
bDLdMtbQCcuEQUoMIxDdVgn6Q13aO/USGGWQ9jLn7CadSP6n+1tDBqrCTgOP
i/7HPoqwc1DApDpu7IBo/53zb4STMUwjQNHJLbQ3X8akA0pEuUro+cY0lDC5
nc3fuxHK8Y5SerLYq4hL1AWiTF17YJUgbRQGKgFpVGFRpPXuRWS4TgpEM8t7
10Er1YFRHPJS5jB3K0VeSZQUcvlVJzn2DIu3tYugeKhl5Y+rkTlbH5De37/8
Q4gHpwJptlo/h8sKrFtb9hEUBqwFv+p+vKV7lHyjgMXXBYgf+nrS0bm0lpH3
5H2guLApfkO2CXzfINa7P+SnAoFhZ4qcm1/DRBZI4m75rxbqLePyLB3rP3Iz
H7A5wyEthIDWpQHOu1Oqjky+5FeGyDgvU/b+tAmxi/JfoHQK9Kw2VYY7KPwI
+Ce3saDS1XqMCAsbCcgqz9MpQJT8rGf1idcy7F9sY9xke1LvochcfeXgdntF
1DRzWaFNYCnu+G6id3cyzv+9h1dM5LXIGUaigsJJEiMJsH9X6Pa+9m1NsqJT
+6jn8tbpqni3ucVuEs9L7SaCJRxRUMbde2pcyugYo1cD6bJwndWfrxJFQioF
59iyS9EgTm2yfa3VC7plRHSkVpgukPh0Rx6ybWryLVUtZ5Guu6ymyDqzYYzB
2VJxdOzdBBkK07ImNAVXl1cqpIxoXk5mI13Cby/sUudzxcJ6MpVJCWcy5X9T
YmVmpIRB/thjRgCD5SD4B1unCOEu1O9YaYsgje3ePq2F0UlJfmV2aGiqdySa
V6yjzUbqgKzSt+kka3NU+dILBgckfYEwB7rKWFVe9F3Qnk6ic/QgoUMuF9Dj
2slxfxW5bOu73VA6Hgr00P8Ov1UylmXoXDDNPrajgHN5riF706DpKadffCb6
YOHRLTSXeoE6VsPZt3F2cKcT3hzXz7+wM9Ywkkta3GMrBTWGPRTR9kXyJ23w
igMFe6PQI5ykOmjDkYzFt9LJ8Cny44D2GQ5JHO9u8Nhdx0vGrkWG7Tw3w1Zf
ymBXXIamGArUSnLJW3Zgh7FKUhqIwEnHHhxoCjqWUrMGTp/3r4v+MP0+8o5H
HLwAq8rordaVJFSyBVOBC8MCDCax3lvj11km4gTFfSZKlNHoUtJfT5g+vbUR
k+I9tBQ2P/zgsXyaNlzgfy6p3XrtP0G3clpg0jUqwIkBLSM6u/xGKpnBEIzX
LSsiLIB8YSCXDYHcExc43RaLbfgSuoJm4qERdu7ygRg6XTzR9b/pM7+9+BNJ
1OUqb7+UcbQmcUKrb1t5CUXmQWYk5DnlycFBqyG9vMi5sJTyXIrFflR4hPH5
+Jsb3d8g5shokjwmvDspf0+5hP30xrQjJKDr8fkp74OmMq5qVIFHUBd8XszU
+gIPp0uwaytItbNVcd4FxOk9Pc751iUkIVIgtNoTIWTLeo3VXezvcFGnzaZn
pGOBQrCOSSfUQPNEzk2wlS5wwSvGVZznitF91mFWAJLuLV5hlezWoRygZjHf
fNABfz3bLBxrxTbR6hFpxNllfYU6dh5m8quchcBdguFCzBSNgnFvZOyaCoyH
1hYQQjAOTkSvOsL/yXkFwpHWMugML+HMrM+r1b+w9/wjYzAj5xVhy1t47ZnO
bhh5UoXRsdCVg7zyr3KlLrdFXO8AUXURD1JEV1wEynE68SgbPMLkFoqxc895
SMEZV/y12sSa+1iDjGeeKzte8ruoQhnt/OniA+PcPkbCQJUA87LKKrb+QPHb
/RkJqOe0Hs0Ik2ZlVHiV75RpR9Lekn5KBD0qjzg2Bn9T4dC4aM+AkdUTEi5K
uw0tJpUZo6cgu+Iexr0sSDrUwidVVJzNtkHjZ0H0QaoBJ5eYCsEsGXeyMIfj
cURfyQFDA1wqiIJX8I49tIJrH9Fkmt0p7oGyFIVvWwss4io54HN97cQvl/d0
64CcGHMVjgoPzXvhX1T2tbLFh/DdiF2ple975R/zHBA6T2kxFClXrKh7cstV
C/WTqaqe6rv6vGFCLwBjKC5nY/vjamGpeS8ZFQoORbqNC3SNamO/j46On6Tf
5Xye8/VJB+ShIR83acml0Z/I4lVhdJ0W4f790jINELiXWF6UjwY/qneFRYHu
0uMOw3h7FcHje4dE7Jx3VT/8V4oELLWobZArL1UWnMN5qxgpOFR95JxFJCkh
O91u4aT3uGNkEjyXsVqkF0N4T438Hk6fVkTxQyR+kN3mF3xofL7iBj8pkfd0
E8DCDacA1D7LsKJjDSM6DvWMVCv9DgVWI3gFF85lOZC4ukqEsK1Q0+HSUs5b
7WDqnjVve9OsgxiejQiD/gjUxAp3EPyy+umn9ZFt8GlMgXh1xikFBwfmYEer
voDeV9+j1fAAhEilyJ+afPJVJJRl2DiYDFudDxeWvdjX0ivHBjodwLJlma2G
xoXx3qxIwtveaYCagSC/9acQk8LTRIPZcJhHzJWi9R8XpCY4i4poq3lSEUwV
gx+aaiV7UmcWK6oA7MU0IQ9piEre2FmqT3VClUHKe4G+1ylWVqWtTtrwG815
6ADzX9KnC8PACppo0xie/PT4bUcwl3lD7R8wCewVub02UrPnySTxHpTCYu+T
u3TAxaUDwfdAjxT0F6WRM5qQxrUyYt5T6vo35qR0enoqkFDghBJYAglFALur
foz+BbsIJ6O/gCI/4ujwebw7VPnjm9Hy9G7x+EWj/ltGkyBpW1QU1gWilM63
i+Z6uSOd0mlsqMFs+BqTqj8ZXV3nBiIVE+HQF8ikOV62tK4VCA29OTSmXPl5
07eVKGsZJpZAn5sbr3xC2oGbi2s5vgraVYjJIWe+AXeUoGgg3cn++RAMcK5m
7NEaf+eAy2xVIoJ36A/cGl2yJw8A0rvQHbPvUUFWWWnZAkCx7vyJVEu+BFgp
J6tRLt1VhH+h9BTUmvl9S6Dvn+N7ckl0j6ad2Z5gbEC4PWeUbZQ0fAgmJOxY
juGR7Vt5oVn0ki9F4rDO0HKnQIAhd5rPLdvtSFT85g8B8ub7+XtIQHKexuRp
MsYqJLqyyiCtZolWWqWkHFbYRBB/1RWmeuE87V5k3S0cRJS3MDiHKPFFmBOv
hs0Uh1C4PTDAKMcYKfCKTMeTJPnQvMRVSrXY6N7n1zOLBkwY03Vg1W7FSTZx
/Ry0OuIcmO6XN6YevkKaJmXJMQC4ywwh9b7jUSsa08RiUaBB9X3qaqDld0Bj
694Xbx9XvR1FzAw/Lpz0Lv8f8ZuYolKT4oBVWX+i5D8J5RulSLG+XJCGk3/H
lh+4CeVCOSN2QG+L94DECj6shM8SUkz0iRU6bhvJ9aib7EiDgnAGhVVffiIO
LwDu44fd65b2hInTzr0dcZvIEiGEfOfvKoBvANefq8t/FZ80Y1LoLt3kIjzU
IFXxWEXjt8UUsbbBS+oHo9WWmYoLhGxCyTPAMWA1w/ewHR4JeOMc2tgwU6de
vLNqbnVaLZCwt7sbO/lutOJjalJKjNG9Cf3t004UpIGFc4BibpZ/7d8ukEzo
z/ekOKem4rkRER12AU6mSYuHXvMsek8SpnEPDLVoPFbSo2kWuHvq06Oyp3CG
az2ljvqeX5GNC+QF/p6afOoEhz3GplAK6uBYfQ+ITEs+iMum6m1uUcgDMiuc
5if3KCmUvkU+VBLbAQFut6zcl5cEIKV+W2sY8Os8SSkuTB5/4yGMzG4phe/b
XE7YA1bbXEDC9Tf+aHPzOQ7Z/oxCpr5lEbgl6N1YJ/xOt6jH3TrK1JV9GiBr
YN6I4V6GIwGFVORowvQ5cthXVeBjuDqkiFNg26xYFAa3ZaoJS6LbdE5BKccv
7WRg9aDGQkAHo+qMKcbztQQuH5xYgxh1JdCIO544EuD2Kkjfa9uI9y7UaTo4
6YcY4k2snuDj1pgt++B4t7WsLl+W9AohbNNIpazPHnF3X0CJQMfxMEwscKLX
JfbFGvr1Ab0IjTTThMKI+vWedJB72UzPHr2BVHGhop8lx2PkBhACTr+dmp/8
XmVVzZivcV9lKgCpaIyMH7EkT3NdAHNrfcGmnjXsI2vT658Ss8Gzr5aPgwZc
8ISjsiIvnGJ+ayDynKhq2EDM9NXS5NcWBIfLr+Hl5kbt0i9G0DS/Q7jDSrSO
LNCI0py709oqfKuqCBW+KF8bSO59VxXY6HOJ1WQO7aDESHsfUplPCxgibiPQ
iV0jFNIa+Y1K3CyjoVyrZOwOsrx8NFFSdSe/yQRlYjTqs/e3y/2tdG9ff9wC
x144Ofn3vFnRFNYZfO2IrA8HX8is3WXWESt7WjFilooAme5kJBVj2W+HomOL
QBtP7e13MVrNoaZTfPWlDzD/G9bJjVyu5hMuJDeUW0qHkKxaGJS/xbh6+CyP
cMiMp50uMC/Qe42ew5j2Al+UTqwnN5XRhQxEbKDglh4Y13Syw7WVFDknCcpU
NiMtXtvc8DwI95uvlQVeIy98ugy0ALArLr+RHQvMfSXugJyKGNzrMQaJwcjY
6YvohC/bH4vbJkgy5on+v5oWN86FcxYwAkZFFGIQm/Wb9asVuYf+GzeADtTg
BZDFuUe+/XC9cN40P5BOBa5ic+7RJP5rVe3NgSu9OElz7DUXimPPoaILGjit
X0NJ7FiNazb2uRGh6BN0YR9LA3gXKWr02p6hSQu+eha2RBBg6xdp42pjcn/g
QoLuC2cYzWmG+/X6AkCZye5Yf8J7hf7mxJLHPRxnT92dXa3OpaAJ2PVGC3ZO
MFXzrjExxsL7tUQ7pjuY3momOsHK19ypra76t4AfgC/9rZ+899JujwhcsPLs
0Gc2TiuVW5CVCF4xUHR7/2jgFNeTOyX0Xi0QV2OOUxlWQv6Q4DgbSyzIqe8h
Iurnia/90HC6wKolE9ORIBuHT5qGtm10/X2b9bVQU4pOpMoxli7amHOvChhr
AjiJwZGFldIa+aZKebGrUZVAzyVWPd751aNC6t8+GZw1F4flBSRX4o4w+/3n
5n6FUERcLzb7Y3rj+JQg5fjVfc8wQxsUTDp20j41gO1QWEzPvSADCzPvnXBg
CJCfRqo44AvOWN1NhlM1uUH8aS/A6tojLoMicetaxHZQUhpUIf0N5aWeJEbB
riaPETzPKlt4iW4FXYpASr6Hw67HrcGoOGCbBGyK+ph/T0zc8g1YOR+5r2IH
9lueKGLZbGY1GG8ayuQfbpBE4ORmw/ukdKuqnsw8Rjc/92Z8L0gWqmO3oe2Z
y4jzVIXVV7EZkq4cEIWxTmwFmSN8q77r9MH7IAvGFZbY3QJ7NXfoPfF2rzrq
nr8ytQlZxsp2KklVV2YQbP7DpFFgJWrClhqolxut9Zth9lBIPC/9zzLip+H/
lYW5qeN9TWS/3ScY7Hnr07Ls+216aPzXWvFMYCZp97kIRabiNdVb1YgBMCL9
ZckxXRzmCv9T0+kBFFcRlffHvhwz/IMJRqNdhbQQuEp0bR8AfdytycAk0psC
UFuGNoDuL0e+Nz/sblxtfpYsH2GypTSlygQD7I0jl6/k//K/uOJXRbHeC7KC
C8Jqeh9Oxkjnuu1AhmixUauZA5m/Kru8oyvUPB640U3S0fUxApKm9Uv5SWvc
HBcIyhyXaqPqdrx4oU+Zz4EBFHfReGxdZdjb82t016NnXEXCptimY51D8iis
f1jlUtkguAFKDzypErH75Iny9TRWlKo6+6gMtOTYS8tbXTWc+XNI7LJ6Jx0z
MBGyna72xTpQLoelcy2D4W/Jh/DvUae9KZrFNytpzwrev1LwSENlZLFQqpLv
7Gh2lc29LsVfdpG6r6GgQGd3CCun5A2oO6YWITqY+xhsmgwwkh7lpQy9FCnr
AYevIN8UbNMESELPmZKvShYnFaWZAcHuH8V235MvyZtAGO0XjWEouEaaWl8T
kcYYs8A5fdxLPe8IXFnCalxr3nxneJGyLRsTMjA92dEXG1cjDxLwfMAfpMdx
Ikm9cZnpJGtU7aajKYyKz3LWD9hX6191tYYPksVqygCTHQTrDU/9WRZ5SPNN
rzZmHDXN8UwJmSDsLga/4phaTUYt9kba0IhtOPEZe6gqyNdcf1eca+/S8e+L
Tg25FrCWe0X11mH2iWFl45PwrOten9sTJGIMxqxIEIw+LRR9Wm9TOi/j2KzS
K4g17KZCDz1yGEtLw2HvVSWzjw6zL4SAXty0dzx9XhxjzgJKcKHM++NcFeDl
8vyzMp/gebXrpdN4RtC6fdVPWaydDTwaWlWm0pdh0RH9izGRMGama78Zl8Fb
bI0tzJYF7PfsUOAD3apC9zhmFBhkSgHDhuVPJYzNbbyu2p2l6jtTZtmboBV4
gmejeT09VTPJwlkaWCw9sng8d18GzQEHNtXEnwP1k/LA7VdnvqHKYJ2BomdF
9+DzFAmmymb/+u5QWZlpulFNPjJZZzX6epESmjmhJcOh/u+GZkykGtD3jOoE
01HzQhZjDizs685EXy8tRvb6ot4jBDASQb8mJHT9s4sRPwZOO70csFCcpgMZ
T+EsVLp2sdcxOQp4Zj9inSmMIEvzk9pZe5/HdbD0UTLbE7WI4gYObDEI2mcU
f0XyKAMg9Wcdlzm941HDjcpXoWUMauZsOnsXoUAoUPqW4BoMA8gCaaq2pCnP
M8FfIW8O3ds849Tq8fKosv3pPyt4HCXJpmtXgayNNS9iZorwtd47TkbygWTi
gHcxPljX0WIZlzI2PAypUhLVv26Lg+FdQKs82pyQh3YnsNOmvoXCtJSmdKRD
Rsm4fFu4T1t6Lvvgf2iK8mRtMfWiDz6RB7cvzqtih4W2wbvfA9Ot6rVt+1jy
u5K8TRWIHjH3QnVf6lH/OGX9WF4vkLSRssHrIuzBA8MmrcK0+Vqso+uBH9p1
Wfh4ijIM/74cOhByNrJVLCw6GXjH8JSDRNEw5a2drErdaQKLZ9I6P80eDNnt
7yZs2sQ0kI6WTLfKlhYzu1ZX3avBWNLlRNdfGaPs0aokMrbUXTbAmnphZhJ3
BwQiS5OWfRzKU+snZep4+30a/f4h4nWdcgPc6Na2x7zn8xT/pMzIYRPOsEPQ
U059QqFwczqB3W/4vK3S+R1Rx/zijTO0upJdpcUFGA7VxHqy4oQzephQVYDc
dWbhkvD6S95Pecty+Ky1x/Fra/oEr4EC7/thjp8zCoqfv8HqpSkynlGDbnK7
mNus/EFsDwVeCcCl96tiLRBrsIOp7eFTm/K+LpQswVY69pxOeYh+FOFqJ/Tm
R+JOgDmxqFNb0RhCjaVvoM9DQU77cWucThPEVnu0ymhlclTBgiCuW51WO4r2
7Autw9ovaI2lC1vuG3JUpcnd8dYxjhbVA8WTdfNA4inWqltFsC5U3eoN5ShM
hT1kM9CpLfHSRx7rPuJ/4P92pVL6LCswDJBvEhBvU8jwMimeWUzu4hvhQ/Wb
n6a3ceMjKR7X9D/1yaatbfjfrelGLR8Fb0f8a2ysR1SDv5W+ABsY36yVx4ZM
+vc4EApE7JIBdl4jmizasmYTrOE+VZwGyl4wwMjd97OLt21aytYgZ8jEsX27
6NkdeKafelvj/haXrZTcr0NFmbzOU46ATIpC6JxfG4ZTiZAZcEYvz39Eb7UM
I0nMsILox+dj0HG4gN7+D4MpiBeEJcNlEkUIU31r4zng2X2u5H4w0/6xWejL
BqgbBDBfnXZkt43WRF+YpWSWy2al4i1BGNCvRnzpFZCChm+szULK08qReqE1
kDji+ZAQX6XtXymZC6A2ZnIR81vitnHqa/UuUsmZNGzbdNPDYQ2NSWQfgimU
bb3oNHiXa4MUecwPVqpOjVl9beLikxrHU7PrIn6AVFuIxvBAkH90thySS2ZB
Hk5QSJr8rQ5ryVGIamCn8fdjMOYEPA1SIoAka+yJX7mH1a0T3MZZBW1J7zMi
MfEWKPgtP1MxM2QlTbuQMTUeCKUAYVFQdlAINEZTXWMrEtyupZj9sQIlN3oR
hTeTa49xoYEYIAQr3RvdSpyqPSBUgVHP7eW+ZFP2PYu2d1SzYG4NLQgslOlP
+NAv42kAppjrT7FWypD6UYuV59MbEvdLy4cKE/vgawMT36Cpoe6zSHOUcvb8
89JDopeRTGJr4w+5G3vpLA+wLRbOoHrtVHxkrzJUmefUNpkQfgHZfC9sSHQ6
+H4yo8XwKKht+RZbE0oPPqpyKqFYlXC+E7TUo+LNTDiqWUKfJWwYQcq3t6o9
yslKL5nFIisDx0abqIsrjOOC0P3ha0ddH0pEe2UKM7tiBtJzJu05CBMAt7Lw
28Z/2iIXp7M+XLh5zQow1LVgkBpNMVucNIZkHHj3WbeoNeugTt7fLwzORoS7
rvJlYTJGzPi86+S90p9NLnlq88XmjBtY4fZJ6GsuMO7612NU7njNOldkruSS
fGnKzYoIWPGhUjnBGLptVZRie5gGT1IpH+r8zHykroaklfD8kgMBooejG1pX
UhM6T2eoN/yMFTIjJiWtFBiTtKWn/st2dLaq3dyPAx4M9deX+VZbz6xyBxT5
dJHgUMv/4NXuNIFoB/gtsv2TS2LpA7OZfTZYvgyWsOXzJN2+DIb0QTn+7x7A
lQi7ql2GR2EhBqlryFqmBOwWBJWB2p+j24aB+vIQgTZYZT3JuX8BioTzuhzY
EB8LUcQ+g0VtIQBQTkpDMlST+g/itJ2wxw+WUbk/9RZy8aePt5hRau2mXOg8
fXydR9c628wfT21P+ZQRK1wpDU7pA1L4d8AAwqgNHLf1gU5vsl8dp571lP0b
KStuEHLwZ2/bYsZ/VF//i4OEvdDuf1rxwI3zf7WTd/xdo8kVAh3F6DjQtiqv
SbefuOqb0SUtOl8RfG8K1Sbnex3r8+DX1b2t5gvTM4EmqlrfxG2nx8xU9LoJ
kje1p1PjM5QSg9RBlvcAs2ASerrDCW8bK9JchcJPZUH4pnZ5m7UF1g7489Pp
k1d/2sZ1+GjR2uomM+3IdjLEYkmZ6zP7kaXfQLG7JPSw/HUIe+XxvLwaU2MN
gXRuArTu9iwWMGDmCOjIAhnarRABi5aHfVJnpxfFk2Xm00dNU4VufdZZsSJt
dVcabrwXkgMJz8gyXaUqndwlDg8CFQJVBDo9ovX0SW+kf8KrLynCBSkq7Jmd
BEYICdXA3x2uxvwjYIU+UmFdQuuTu0jSsxM2P1j0DajSOGxSzvJd3StbNP5C
5MMseQ/1mWRTR3TzP5lhTUN+isd2lROPqkyg3IRbx8aPjKKYzGA9suoXQUfP
XVXdH/36G3gdYtLXqx126Ib5vxqhwQG5gjjUI4D3CzLWJekVh8Gms+adH6OP
MW5HEOk11sf/GYnkVApG2uM4nr+vOJQLuZvNcqAUsaHNEQo+JsJh0sHmmC8I
ZgYbqF8/0uDCcyFCQEByuas1GeIkut0gOAgxGYsz6pXTa0duvsRZ8yEuh7fN
G7SFY8SrCc7d3Mw83MkcIVu4UAsB1UE+RNfEthAdiMwVk3LTDDyBT9nu4lZq
N4SjAJ3p0XuhINeR7SoEfjypnpjQB18vKhKrkExpqQ99Y6qpra03UN9eAxBv
8dAOE53Yx2V7X2jdxhM9AodSSxa1PQfvWR45i0A8Wj1wPADLI6rVCDth6rKL
FdzihDBBOhTRlRq2FeaEAk8Eruf8RThqhBHWdwFOuysl76/jHFEWbxULb391
hPx9s6SA7r4VTZmYcHFcmwbyckCGYiqd83Vnopb9JyBxq6hkvANP+y01qUbn
QPDUZhItiABpVMJH71lBoeYR5tIrB+tDBY7eb2Rk26IfspGXRLHFV+2irQxr
aZCBjRI4JBuXwvdrDQ/+ArutVTJXZoKCzbN7ExJ2VN69sCu+GjFYGuQcljV9
YPfQBa70kS0kESaq7KpUPhS0VinF1CxZ/QAaJ2OhzOiH0OIdz3phPN58QfSl
x5BvZtPP8er9MgGYI/2b+De5uINwMXtQs2bIA4j2uHimELlNbanqUzEB27iT
a9f8gk78h1tgWSEVj06zjUpa8/ndf4xfBjfwzKZhSiBU58pIwv49434ktdcb
fPgmR2t4hlAj+H4bxEsT2DfShEF4Bkk7jdVUJYXvnOlySvVWT5hQZPOHpb9S
YTPsDb7G6bXP2iQyVuDlLcHsgNg9f6dGKoeFhBrl1jYzIflwRZL1HOJaC4Dt
0J47nn8eIfaJMW0Pyjq8llRf+93Eg9U/92uPxP2pqOvHsSCo21MEq3Iodo4C
4grgUPg0w6cZt5XlfIXMRla1MFy49s51jOnio9K2rNl9Gpwyfm0A2vA7GyBY
dr5UYCdkY4LKOFiEQH9ZQ3wOGwUmqKHFXsEb3/jNYLYV4t+AHk7avwo20Nv7
tYkX1PxX4CHmEBXfNT3LeBUqPFah7O+OhmPcziWTbjDCxyojbjNGbcUqmD8L
t2+EveA4ty1vWZHJsvOKQh9neVhPu0dgWdhuqbMbgKAZneX6U1OJmjkrBdSb
zyXKet4B+0muL0eFep1VQCJSmnXMd+HIgB/NrOgqj1xHjP1XY8lMglAxK5A8
kc9H93ru2/PhgBV+IezTKgfChWjQz+tAPBRqTKvuXxBPdoiqKs6LvdRLzkc+
iOSyAOCVX3V32jnxARK5362AjgR5HXxiidcCDhJD7Hjkiyj+kt3jtoYM9YYx
BFCAO86vmEAzSlpw0GKwHoHbZX5Ws3oMlXMqyHc5Slr6NFlaQDWbNFq3hy85
abmQVucfGVvkpPD9aimmdKIyYDO7b2TrZy/BAX5XS3RXUU07bbhc5l8Fqdox
Rs9KHMOYbzRLO7Jbww3lTYG7i1Gnt/67R5XSR+y7/5aBJEfelPU4kd4QLRqG
bsJh5sIcaxthF8z91tH0e7oEdumR4MrMeGbiYtGdiyEo1EZDiihDmlrRjbjP
PFZoP30REjtzBzUSpk/Jf2wd/ik3oC2Ja7HnL9MNeTjqfx1vT3DUcLBto/U3
k7GrzWsOLSqQCezE1G/iX2yWcTWO2w0mVCzX4N3GJQEW0DywMy4YTi/2bZYN
uyqkwZGrpgkAk/JQ7sAIC3wxLQ4ZIfM45XSRRqmTC+6hUHulfjJOSV8GvZlj
0As+hR50wvLTOOOdo5p7qd6HHZ3qthcdqd24nqEHgzy0pev/5JqjqUDWGiyo
UotTDXHuSrWNBvqzM2Kj/jIPlbLqS9D3rrNZLiPSXF4fIzpyM5qUVLY9wqrI
q5pD2pRToRxiF1gvg0An9g+yRWDzOXH6sXsW2dOnauca4aj6WFlOTspOfEHw
goYNfJonW2N4W5zw3tq5RDpiiGduwPMfEsiDy9NfuA4xTh5xe8B1mCnjgbGa
p7VjU4stVSdZwPmgOA0vIzPUxWDM7w9V+D1Ixbb8//mwwvTKMQ3WlbeVIuai
rMxfngoHdfGiOklz4d97YXU9EJAOnZpuUpMQfh27uXfA57aGFN4pS0eUQnis
lO1GxN9PfnjGYEBIXLfijwubceHASFnLspc0UvLMfG0EOMw6n//F5JxpMdVR
FE0EvVjs511KidYMxIZrW+Wu60FmlTwhW6GOO8x7Vil6QNV/3NIb23Acj3OE
1X9Vwo3zglBfxcrktPDoLXgT8rLtTjEvJ7MG+hw9dMmIlXMvNVUPHwp4Hfbi
UIwrvlR2y47KGgYBTyLULiAS1x7my0tOKI+bohinF9NS9oQ0NQ/QZTI7LJSK
fv501zOukq+phyyp0BuBvRJw8Da7WdoHrNCbxDnGKjwbCdZZqnwxtEatNAAc
0/D5m6S7EFzzyWVbBH4TgUIK3rKADEU9Nm6lYPF0HVRLOos7vl1QhivIeDkx
Eh8zLuNhRko2o+sU4qyL+TzbVjDOP+nxnNU8inxYSRH3kqkHLVqrUTcZpdx9
brRdZ3BoRCfhbg9fxZ7B/pvvcxbQ+18xzAaRCIhK1DEa29/6uhmtQdckJynC
5Qo22SYJInDiL7/oDeTFh5OykbscVtWFZXNQgamKLKNYyF0lDjAdcqWv/rPX
HwJBm3B58njgAmbDnJ5R3lLw/L82ULQIlLfmbq0jCMHAoFLBIQJJeeJp9pXd
8hM0+N7Wy5udA+1RaMrfvFyfIStl8dm2l0emOLRuMkmen6N+UEH8eyILwWKH
rKZ0mhI/Wg6uvv+HXhhppgwu1+/XTmHIfjGQ8I8cEDtdG7JnhR/hK0UIZXks
ZiJ1OxP+u/BNIhb5eKoAbZZv02OK/RN+MPeeYLUnvgc4FgLgEIWKl6ISBH2M
LaQOja3+cBR/3G2BtKcms9cSwzOF/3LLAhesuKMesynhPXitmEmYA4hHgFcP
M1+b/Fsd9gNdwxs4Hb9n9nUHGn2JU2lm8TH9uTou74C+nZWbq9x9cYnyFHCy
Zrg/FPcgmnaij3T+qlyah4iMY6cpusjvXTRMYcS9J01qxJYLjl5ZX7J4YmpS
MpFJb43MjjpHjsDvcBubDzLulsCecVq5K6mQnNOmGfm3qnbiEO5Kn5ifjil2
dlyEieprSl5HayQv4WDwLw1Au7E626IQnQgLukDN9++IoZyzQT7zOFgoBl+f
p72MrKtWMd1I9nnbBhrzoR96yLYhvloxTkBYSNbnpwDTtL/LgKh+s0hwZhII
MjCMcV8h9mENWOVuQ4HdLcXGIiaTHuYHgxDW0psip9+HTXJwfcX1NLN1prCT
Ynst6pJj5u/btD7oSPHgRevsopXy7Ubg4AmV/SxHweE1YWCzqyddfOPRAcVt
ONksdjlZyC3WUXHcBszjx1s7fDTbOc0mKnFXjF4jCOLyVpk/rxq2cCfrzT/h
bfcRH65NYrkyUmZfqWx76ML90RwDiVVFziXTQIbKW4E9jU83HGSWNc+q+Zm2
DtYnZQ9Cho/v1MzJnnYL3EZ5ISjsQcp5Z2ycVAKjnWJ0MHUapsonjQ4daR6d
xFeZAToGhK06HpfU9lUm9ITKIoRgyUMHYb+l7+CiNRU5Hmv2o8rdvWDaMF1g
9YtNcyzkmU6Eb2SoV7rEuNnloMN09UXT8Mpew/IxSPpnfQ8LJn8vN4db81Ou
GHZjMicHJSIzTytk6l7cuE/wLxpouAiyyt+xLEVEzBhX5B4DwW/qRGrOxYT0
/L+cRQIU6yihj/KtZ0MOVigJgo9gHXoeqi+JH/404VY8gY6CRZgxPXCnXggO
H4DQxqfYwXlRBRzXpVCea4xBK2zoaUM7val1CmWJ6gy5Z+y82lMKjn5JUuRV
ifTA7N5j5llvyWiQ4vJIQmoe+Ysr047QS67x4YWtNJMs1bWNDj94a4cUsorQ
ofM29G+p25zTme62dsNZ95PedlZUR8f4Y0BPFvXyTW4xBvMswVECn9Ru60Bu
zddKpfpzCFbGb9LAI/JHr63S5TD0F9+ZyiODtkcZR6NfduHrqSfnNP5PkcAw
QyAo9m2fc4r2cyKjflgY4a3/YXoLR6HzXALFcCqW1XjiZlMR4KH6ztvmLji+
kOfBR05dnbqRPsSoYD4LpH1rfTXGoRYnxXnhWzsuLs+98YuVSR2V0SFoADcm
PCeyOe6ccQ9HsAoUZaW9OtDO2+06Jfa30KdTOQZT8M+PkA6uPMTTefp/RxJ0
1kAoIg4oauqPBRZrqoSf/vfYA8Tc8+yB3AvSheybcBaeY5dnB9hF7F1iA/CT
QSSRAwbY4CafPnpJBzafBY8LOdbdY2S7lW/PsamsFvRl3lMBUB8vViMv3XNO
T7fLxjirgxU9FHKcuoZmYh5ocmwT1HPApXOXGp9GmBnNNRfTyUyr63o0edpB
bHy/K2fPhF60GKTpMxE81iEsuCslcPtrTRBePR2fyUAx22a0ysMC/AP/1tSX
9R5S6qHP/+wwg4tlJHTasi+KdMWCHetJqr8O4vaNItm522pE6MRWE20nmzl3
YiondDcL6qKF7Vb/DdRQ3RWzCYAk3VTRwqNafbOwLB5/WOWLj/HJUoslkz/G
wh1HHRC/F6BT2Qf4VG08VmCrCXRGD0KvuwyHIYtIly/U66MPoTeOioFKkzuS
6cJst3ONKfgQrNQgxVdeuc5+16k2/bJKcEouWJeQuNctXpP4+22ZreOdyEMx
Wll1SUrAnYo3uhwqL32Xpi5yArviKpms+YHCqzcLYpxLW53h4Vn28IaUAUGx
7BCbvrgslKFHw51uisEyEd51TdjGU+wEy4ofhHQmSx9FSoXyuBHv3vKLBz/H
NNkMB7r1mtFabNMOEE1vmZqVNm11KUjs3Hy0985L4Dlx+tPEmHv2tY6bjL1/
s1HZuF17iAnv5qihJYP7y7FyFSyZuKznuH1yHMZa97S5HoRJ7kJvF4jKAted
2kN56P25Hty9DQol/EBW98znfoOO8lBey4yoiIfnPsuisQzrnD88Ski0uU1x
6fNVpfjjADxhWcKEBsc7CTH22Yi3QshAmD3ry12t3buusjP1O/V4+0R8ZFbU
OnJ+osLClK7fdMx1nQcs9ebxABOiwkaqKRIg8DBS0pvUhDKmXOAY9mpd8pV/
xBcuORjg2EqDrjqN80UbYS9rdM32fvSP2ewy9vKOA1nLqZ/oT3HyMXFiAxb3
2pb3dnzH526+GTbMMRj43oPTWJkfma4JSVPeVUqs5Hzg6Z1NfnyFFFVW3oI/
fKayzToJm/Kzm/TIqhUxUcNjUXCI/pVt01RAR/YrV4jcQOJtV3Sin6UNfug5
kQz2xFajGkaesyxBNK+PtOfkb50JQoJDKuAfZgAp1ELK1jmK6smr6Dbpu2EK
aO6OcdVurfXnHYvapvKLf0AxvD+D6poRNn0N0Z49mSZEZpBmA/cn/wp6am1m
qtinPnPcr+VyWUnBGaTs6zEPERN1mO4M/9ITtTfFmCVpYopTUnynf1AeWU3/
mUDANAe7YXepMqHa6c9NjvnCizA4LTzz3FVWHvYNWWopBc2+tt2vzxzks2QN
md1Ob5N1EEu3fXpg8pJoui80O6C58q1J9HQ/fAo7wDUjSy9IZ8bJ83il9P8X
FdktbVmVCgytvFnM3HQUscNIf5CV1DrRM6b1uKwtFNl+dpOvkAQgVqA0wJez
tmzkAEVFOmncdojpxpSBOCC8WiO4YjmqU3BSBiY0SMCNkrXoWl9Qvs3k711D
fnFhIkLk3pJD9ARFxiiKf0EhrNVBeByxvL/JAbRiWIB7iaRPA8sc5xXBPyP/
Cvh/r0fycts/cVAcHYYevcRHbAg+IBJhYAvykSdb16EoeoLelyffNTNrD2D3
psOJimP7H52r53FWjG+Ga5jdN1WhcvK9qy31P2R4RumqsAd6HTlX0gCpPK/w
p8scjlqx1rxpZECfVFnC8c6stR9Jym0/0kk5DEcwRyHafWh+52SXzP6q/Obz
fePodnytdo/ji3ba4IvlYSB4lRITnQzeYP0qFXDkI1g4LMCWLMTVQur+WBVA
3wMSFJEKqrdKDchjGlVy75cNW7PYy6VsjQeSEc4pdw3rNUu0WmOsw1efP4uE
0mNA8fKz1fdKwghnBhdEM0CeLI8cw14Ajl7nQm22izJdhgxFJeEtXJlrUTIn
9YVrIF9UzF6Xcbl6Lz63R0kqm80wOvjfEe4jaGmd89GqJ+m7Bm++YeIcdVc6
Dh9JtMM8qwsk48YhkFXGCfUDEQGHaTN69GMY7l8yVZRNH9jPriLU96Dkpb6T
9d4xrT3u50h4HUbO1n2bu29Z46soE5JfBkzgbAvFJ/IzFSb06QebIN9qOIt3
/bo10q1sLaPnxg4bn6nXVy2qjEUp4zTMASP+gEjWLKx5TU1ZIFDif2MkYWHA
OrA/eBnbgt+vL0fCSBXime2bcbQDw7N87VPp+MHU6vrw8l8C3UZ8Ztn939qH
BEV90xGltO/DY5GCalhtiXJ8FMK6XL26WAvIG6EIk4TJOxJiKHW/r5RdEmov
H7bUxunyRlammCgwn+zcttAPUq9+wF/dL4kh/oUP4st5+ZGCLRrQyuDN7ecU
6R9o435u1ItDGqNVelrMAlN87z31JjJLp2lQUuHaWk26FPdXEl0H00qojl50
8/8n3pamvgWkzVtPdI1mKigrK1gFt5Pn4EF4E6JCB9D6CXoBRaRpT1dqtKMM
I2qXolOl9KkOyF4MnBC4avsxv/LEPVFqQYVIXnDofAf/DpBhYOWWv2ZYq+QX
6/5YxEfU3BLvSpp+Ig3IPW4x57Lk49rOvJQrQQIYlZ2V5LW2zzPng3aR3+8B
t14FYiH3meeorFlgRvTs0chv8psDxeNld5n2dL8Zkszy47fsOLUxCbWgzHBS
U6ps7CO6uBefr7oSCWNEzJaQKV+t0y0MtIXRviJc6aMk7JY6yIjHcG/FscUI
n6f29DJD+Bm3oCW7xu0cPiKo9J4bZfnD8wIRmWWaj9TpPtwswFe2E1/1ASGf
i8GHHpv4hh2Ulsan4rwJgqwj3uRT2mjiCxXXhZ+tTZf4z+cr2QTGwQh/vq0I
4wK/7eKC8TtyrYpIpK0DHVS322bVSsRN94oTN9Y8pK2n3AsYDePpKpYya2/U
Fj9iaVT7e4BQoEtKke8qPOLWIBBXcJBdNCq4tpwjR+h8J0dT60/YDZhtGBJ8
Tj9HMJIASN3WNhhxR9F7GKYjXi59kme/V0LJGuXGg45/sGKtnyaohHaY0m+n
Nabk4vxEGVIky1+epQjgVopo7FmwhOfB0IYbpcLhEVS2rAxH9n7CxqpmBqcD
T8LoiEQZmcKUvS0GM020AJjl8bSnmXGOqPD5Z9H4KpoClHvmjiHPQ2Nm7wSP
PJmkSo9XYYTw34FwEziZpLAm6OIkLOhSf+QZ6p1+fnDVK4YN0LYrwh0FjQ9y
0Y2XQvczppyCxkTV6QV/3B58+Q4W7c7rNF/l5Fq8upOTgfCuTzDBNTf0PdIe
LH3Wdd/TmZgGedKUyRRmv68QpFCyVK9rNoAXeYYnqmVKhvSZN0y2H0pk5FRA
Puzikq9JeZzvG9FLS3IJQwr/p/h4iVEXnvWg/YFG/4uWR/3Y3p0Ta4Qwpzd/
6tuxv/qjAXIc3dGRLcliUYzZGuKSUdViYJdNMUS2oVzCuyB6eA96fr1ckxA8
67uc9da1j0UKUtqlo/jwKDx0LaiEP8N62Owcz4qVOmkJwRJW7hwBo6OmPcs3
+rUmPz0VboSy4TUZxZ7yOeohaoF5daW4Q8oZu2D7O7vZq0RdDvpYKdezp0DK
h6UnAirlE/ZwRp/jfIARhIzGsnXsAXP8ECLtXdgrFgTcXWgXEVLm91U5c0F6
LmaalP3R3RvGfOnzfydZj8zTJqbbeL2SVuVJxNoLVHq35JQQEcVgV0Y4VZGx
WCWOkdhKg/NHAU1J6z3xdqzXwSJpGPJjwpQle3HcdamwxqZbXYTFYhZfRGiM
J11TUkPctw0tNsBXIwMCs0MI6uFRbglF+rdxcrVBp+lbLpPvsG13veXwopKL
/ODJPifJURkVwi+kg4AycGcFii4TmZMFbH1Nadnj+YA8o+zjHKQHPZfMoaAM
7mloshKryJ1cxGZ1wrmX6BPC8wrwA8iMUaxWb8Dv9ha7YES4D94vEAHgsTrA
lWQwM0PMzrVXMMCw9pRxC/hX+O/MLMQ8IvPp8g4PLVcmFZHPy5L0GBV1fKZw
Q+3lVqnx1uIs/+wU8OQjnNoiLtWKDk7CQf4mjk6xvOS46zm5mztO0OY6kD4o
D9N0sja9ar1joTtPPQPTvAd09n/qTOUD/uNRPnsGfZzglgHFbgEcQH0L2G8s
H2yEyo0ERCiaDIAx7u7iAUKics8c4oDfcHQDxLQ35qbTxH6XivmxSqb7XYQD
okedVX9AFYDLlnyvEIEW4HTYhFjE5R97mf6oB12lEFAPyHTwIXQZgDyeYKV8
uWzN/KgFBbnIvC1A3gCtYiFQWP6deG060Kd+lVDfXBIiI6Vxr/zPgXprBDTE
ALOkBUa3GMOqWdEzDEa9s5U1DTApeqALZdPMBAanR9vJwU+uDTPtjTWKzwXa
iIEUxBvU/gil9s0QY21X1n1WYLPQd1Af1puuH2CjLp29BDR7tGhzainN9NXd
maIX0tRUJZq+kcl9y7uBG4OxjduQpAt2Q/Pn66BV6RQyUIy+BJvGYYyLrzhz
Ypkp7ZvZiSEIG5EHqsXfD4ZzjcghoJfeMqm6HMHgGMEZR13lx0vv0WNGhGtv
y2r8wl5+Tx7jSCJFnAwniTL/ZLNYjZPEJRA7H39/HCs+za1uxQ6alRiiMruu
lu9oUdgkt2H4jH6yBgegMDzzWtC2GLbd5QWmtkFz63YB0Hbf5tWkg71+zJ7Y
mt0gA5H7ZW35xp25hQikHMKYJ1xgC5imIZ3eHNSO9d+kVDcrGpyocALjDZrr
z74UEPaRVb6OyKa6p0NqNpTZUNykQ3E+y+4uWI5vp+Y9SVD/ki44RS8ADPu4
v8D0cWDfsr7skJ1DIAwm86mwNKK88ZxqA3u4t1lqK1V8MLsQLIPWg/o50ASw
PhwClIqfYC2v/0F/QUZ7Nh91mdT8FXhGpw/o4gGYb3w0xp4HLBOiLOIGBWGu
Ma/8CGg95FN8IByboXlvUY899sH1yci/310wcBRzSQuvgvZwu1ypfRwP5H0/
aLT3iZLvZrLQ7oEpW2ZJ+QqS/enbp2Dx7qgQx/JC0SIW3IiMxPI5XS/BKWvj
5zOP+FCIEPtKs7u9evVsUPaFgZXJqO5g/I6rIv8EYQJBkVnXR0OtuYV/c20J
vhSuJvjUBQlUzPkKgdNj1KwdNtbDi7foSLhatt9d6zDmE1h0ImrDEwVAoePl
6KbjNKXlWUJassLszhigAWfqOPz0dd28DRkg+B8CpyzZ52bF2W1RUU4pRn8O
VzTZbrJbt7UEBOY0eIh6w6+hYFnc+rm9n3gBq6oKBCaU8H54NUowgaSdvr8z
7Ac/QOLkrW15tc8YMT+WvOAlrVffeJxWxELdzkws3hlMIYJjGbtcoPr56lcR
css7s3rkFiA9wE1BR0Njfx2mr0LonzMaHTTnJTfajXSijEG3n1wBSQrK4/aI
gly8H/MRebuN1K2+lk2VZp8dW1/fChCgqBn/upEmrHJK9u0vhrWiD8XsM4bU
LEl2s0tZhJr7aaomppjcdX83SlIOkbXknTUtZagFtUK9pdnc7JXAXljC+iJo
XVT3QBl9/NYyCYyWQz1ZqvCUwCnig9AAIE6fwLAZlHOJogdf7NnjlaBpIDYS
bdzUquEbQhj2SpmH4ppLfjaSmgF+7nBWd1Z6G3vfW+ZkAS0bsNZZH1G/QanB
BHIF70xaoreNubxG0mKXGSVMAznJ01bRO5vE5fZMdcV/5Rej6d9e6mjfgsGB
kFHDcQ5IzoeenLtg0SN6Bb53tC+Bort6xL4GEm6QrFy7fSgkylNv/4KCCzfW
Zqy888oG/0w97e2tUFiLMA59/eW8JdAs3Ch8znRiBhuG8AxpPR4c6fDUyScN
C6leTGRRQ/zarM20FnCUEh+fMevSvpmgI6YAYEeOTj2kPhvKpWh0dKiNyJSw
wxA9Q4JG1dlWyDvkxLo0R9uIkEf+4+j2WGqH8vAoHbM0/1RxQHDJV5ruWP2s
KCI/JCr0qhsrqihP4CsbiiR7ahYD6my6aZrfxnvl9U7O47TRupE83hbypXwT
6UVY3xsoVasBm9Xc4x4rSlYed2BFccD9VGMMThZJdRBbhv8VEsxX+PpyVdlT
GpkLo3QAKAv5c/PQur7mi6AcYHQFFMVSSz4sb7HYb7mPWPveuErwckInpG9U
PUXnNPSdDVVoFKtWUvCWQCChtOfatqO1xozP2b3f7qxb16f+GOt09nhqaNqk
yJs6kffY5W+b6mQW3/7+KDT6H/tFT9lj2ul18+vhXiU2AUkPvvzET9JsnOHg
V6zyoBCYRwPsZh7bDd1puKAUQuD9A85OmZwzTZCoFFNYzbBcCCIxBGCNGE5L
896av6jFjP9OJVq1vcjf6fSQB6W80XGG0iqd3Xrk8QY4G6n7JP9o+yaIYtU3
NMqe6M5xRrjGfH5fDFuDFNZdmbYXG8h2rJ3N82WBqj7OdgBv0C5euJU0IFr4
GFnbOpZnGpV6FA5vf0pyKNmxTBg2YcWI7FKaKp8ieo9SOSLmjRrUCSqvXMtW
Z1kfSFPtEOjFirrOvHpASjQBwY+KG1X0P1fa2RcU6b5aLJj8jjaHykf8SqZN
qULny2Pg+o5tY683q7L5rNXzRu7EhOkG56IAx/TRyKx18mAiqdNkdrzRl943
5dSNo9GjgYQYQyYfQH9pGDSU4lb+uJZ3C1taQHE/tIlb5IpYl/uKytOSR9yA
gRctATpG6e6fPymYF3l9UwO4njALsvSuhlY4+B67a5WBwLtQdiZTtsCKaSnM
vGkUp4ifrdLz1w349OIubAd+PmPTIfhbkPr6bBVQc7qjdNdt9wFYZLArEahd
nH5uPuS/MopNJxbiL0lnPM1mmigNwqx4hQ6k3kKkUCRhim+6H1L5CQe76jGR
yxOi9hDGdxa2TbZ7h5xyef2eoGMawrTrzm5wFo5KFsBKkiQTGgEfZG1GB5Cr
8ldMMvwnw1JV8ANI1HyVVKdsnYazHmeeOXmhCSPur7VTf15d30Dl3rOla5bx
fyhSg7lSCYmJeK0vfPcRbsuRlikIv+Im5V6d3GBp35LmnRf2Z/aRmPTkAJ1b
6fcO0booPYdGNcKp2ERu3NIpYwG5ExP4sid1S8J5XUg5Ty6rWGIt/pfq3z+e
Tp4Jyjskt0CaIHWkGm1lhrFYvBwN8cq4vQjeN874mPVdTteDeAnDHu5AMkDO
SQFSy9Ujhx0/hgjoh6legyYmZjxIPPGdYaF5MMTGmnTe0YMxEEcKnxXnQnsW
Z4Nr4akuGWHVN3wj5Qd32xuy1bxrqEWQcWHn2UttXw5eXias1CS3IUeElDuA
WzuywBCxhoYgujJV16EALy+gMjcXOA2pfZ3YXS9Ued3jTggeHSmGlg9UU8gJ
Tiax3xVwObz0faVBU0kE7ey5/px6pMQ/4MsWMghlIWfUZYGAGRlcqZyVT+lB
DwUISNOgZUCgxtt8tylFIEfcMYJALotVKNuuzSN/wuK0AWs6dWcdSw7tvdxp
3qIpI9TlzDB0OysSBMmAlY106RpCl6LDIYJHSH4HUMrwQZQJCEgCE8ksgH7E
KQYHjLS3bskb+B1NI40jwUgL6Oe9vkGP1RlZO23iRIrBWFn0F3Rs51gOWHzG
nw9s+tEK8vq37S33hZdbECBUILx8AHddpPMPKCrcX6yVzavf8WlGQt4N9vvg
HTPEjOGdvO9Su+QL5oCA/mmFGrLkVvyERwdiS7s6locS8QCgbyvbTqlnVavq
OwXRaRKefyHI9swb4xv/JzQpEjN70w2ZAAfkUpPrAZaXv1Gi7sF0d5Da+fsu
eTC7BwrkcF4IiRKGTyPg77EzsSAx6/OaNwDuKeEtrax3QGcBdcjCZZ3JWFGD
PKtlFYUcHQDOmj90IwPNEaykTfSFo8/SOBcmu+bYyEgHXdBAmVwLsihJIMp+
6osXKMVAdYx0Gu3HW+NOz4VQYUj9Qhu0qZVyIphbn2G3yRTLbQBT3YrKGZsu
72Sss8PV20f7eAGMi2bKkhqZTgFsfThATCa4Zy/0U1hcymyBcc9NVvOhqeAU
YiHaNEsTqjL0x+XzBGUhJWH3bhPNMR5nKiRE8pf8IGPS1+e/YZQEfBb/Bhdm
m0E24YnUJzW9vCgnHZUx9Zj8zy0Uz/tOF79IuYiB4RjnPK3yXesTur5eQaHN
JchVn72JU3x9Q9PKXxGNasbP6iZEKu3BRbZ93Yfbl5Dng2fzhU4f0ZV5G10Q
ETrPvIZPHdsW475g/6+NkhLJpp9c4oxW7vrXojfnDIVAmmDsfW3uoI1QMNmV
339H2qsBSTGuMOfh8KiG2vtTalSVJRa+dCS4ypggbFP7Y/AIME2n4hyEbkUf
X/Nh0B3JQVCjkV705eJ9hfqjwYRwotM361s7e5zvTn3CEC+pSv0HoNahmhGw
N+WRq17kJBx40ik4SrkSMgvwQkGhimseOuhYnQ845Ct1f10q/lVnd9gbvaWv
5JTszUv1nzFeLL3wvY6PcroensUNCWahCOt8+8Wm+q67Z4YLJwezf4lAVhbz
b6EswWXZxU+/p767Isq3yQ5mF0K1wj1DPzkQHTFmiuM93YFo23pUfUhWGiQv
6SxcYyZG8AzLkTk3QzVoGU/JrDW7CfykAX920gZr7O4ViG8CZ0qiQ5XXm59T
vhQm34+a5fC/VIspxWP3LYq/Osz82nWpCAPZ3asdki1WmGKHbUVq/A8/zTCH
9g8onPl+D1xGomvHGbb29eraHxt5dJDwodwnQEqvMDWmDYv6ljg7GUZNiizF
pfc/vs2xjmkKwXMIV3IIqxRnPmG7K/cfomLGlP0wA9rgFnSZemFWNNIkCWMD
frCMEakC3tpgf6YLVRHNmG03bfVngXIsVjgRLgzR4/tHcpE9fl2Gu73asdSu
r/GChR76aWgz6kZyZJCaf143N5HIVAs7BlqKRNuiuAuO8WdCndNxGBPBguII
Ae6xPeHd/HxaWs9mxndpGXzs0dBHLHEcmKbzbdXvovExmsjfic2k3Avfx498
uWd0VZn8H904m8v0/7io8g8Es8D4wAxppN2TUsfCGAknUKIwj9GPCbBZ3MXn
C6y9VbYCAnHaYPGyrpmOTIGjp9t7Hxhbj+7mRIL2MDBH2fqvgohDXa5EPhsv
o/Hd8H0OILWCBRBflN0lGxcmo+U/2PgrAh7cEGVQWBQgi41p0UUvi3/A7G2T
vTdpRedCxZGi0At0sbkfv4Fvo/7WqL0kVWwJWqCCDmZ0B5Sxsobfcz4928yv
qlFJVhodg77gjavwH6n2MVvGjyxPVvSY2QYrJObP0WvYh9Gia7z92F3ydBZf
eHXSf7y8Rp9bxSOdHF6zYPuxKLJRhbflJDZqeszBG8FJ4JVGS/l1dUB7KVZR
hyuQRrYike7RB1aIou5gde2ULejkrED0pWFWYkU0eFC0+AdkqKV6vhkst9ph
ZTJxLfS9YJblvBI1c6fQJv84RDFf5CaXptRR7ZFF0e7XjxYwiUivHxdbIBan
/a4+7FkN19EX7bY9QT3DmP+o5F0k5emttRITxqR+AYmPVt9uiYs9E06ASL+u
EJ6wG8fdMGfsb7co42qphTGaEsIdioCDNh1vlawXiBo6mo8i5nFm3WvFS14U
Myh/SJIg8301v6ny1pZI7cwpsCEkwxSAwBI3MPd4S7evT+dWAWFZvSrBH1J6
APOsByWA+H9K1Fz0NSLO1rzggv29E669DMfyAxIniOuSZYQNafVL3ZhF/Irw
S2jA8W7PUM+CzMYGa32M835AnfrqWihV5uMWZvOSLb0RvfvA5xkj6vEbi9uw
tT1/N9tsk25t/J3z7qumx5EEAFADQT9yHCEFPPokoA6s7rF0kepJCoWzi6sS
wH+jav5TZSCzV/IhCRyzxdim0stiO1So/3BE67Iuz8zG888lRBnUf9i3SWJc
VEwT6ggrAwrE8MRKbgwdunFw8XV5H906kDrZyxF62qGeRxRKBLw8yQ1d5m3e
kBm2PfBDw23KTKu4CIwl9oxf64P5jypXIPKOuOsLWNZV/d67WfEtMSlUVZQB
KOJLDF3R5uqGCslCezjgdT0GWCzhLPuX1XujdqDOfcaMRWY2Vz6G0DAwQpJB
ZOWs+3o9jTRLJxr/UaDLmW6ICGqGO8Lje4Gl+2g6/fzgjK4LwTvusMpdBsYW
FMnZocm2uXOAn2UQV2jG5/YAAmt9u858CypExrgB85yMT9+BjpEvwVfWI4pZ
HextK+o5041ubnfkNLHitFKNC1+xKqMtlA/6iVVdZAn/nfYSiodco+6SpMJR
tJyRg0uhs0LLxlOrequOPpqZtwQ9Fy+Zg3cV1eKxz0bUFXr2Q/D+ZihFr6Ib
EaoEFWgwvyIYxnuCY+QV0C2p2J30JNz77ntiEDovA6EtLcQv5fo6MO8ljC9x
wzzSmBRCdQBNQNgr9Hje4XtIGjblxHJ0Cixrk1+Mpih7L3RDx+NIHErz4gl7
ni5KtCvLLwdvWlfr3D0/JRw4quR247HCjZKA3UmjmSmI76gaNbeZDVlnlMI9
GvcG5owr5WHHipDzDCq6FF/DdeklhNcwAciEN0C4A6qF3hDxhGvVmjNoyRYm
ZWqROdNkZy7GiK65sFbw/sTq1oKUMqV9u8WT4QHJ0aPjR6szLkrJyhWXK9AC
hs5EiLfJjbIrz98LAaFq91AlM8t8wP0xleBkFMjx6TqmjI00o1Bm4feYBO0Q
ulmierzIMPag0Mi7U1Urvm1mIKhFCEHzXOQYRaeaGcQk0ZwmGQZ0LjxSH7HV
1g31/A4276erSNBGtrzDU5waPKXxRLVAVEaI24h+wgamyCrreYH4BU03TZRg
Qn8UQQjfeaoHLY6J0qMRpSWVbbqzba7nR2aYMvJSTYxs+lGQtk5Yqazu/uNm
y1kgQwWSOiECdwacMj6TVeAODn5jnnZavUfvMi3IVmLILz+5EOm6RLb0wt5V
Qwwd0zLrOwvCTFrSWIVVYQTampyhWrEAWEf/ItvuRX6bw41LUFVF9jXHqYz4
9kOJTEUELJWWIlITklFK0gCtL48jrHgpJ2wFpz4YE6IKBl99/A9PyR6sguiH
1Wr9tbmSji6jCGEYafBbYOBcoUzhbryZN5CcPZdha4XXw4Uz5Btl1EN8YRmA
C9Ryfh5AQvWVYWRG/LZztXPbrK5rbwahrHqxuqiz6Ot0DlIvQHZ+2jJjlUTQ
15N4M7M2quhwVvGz0UDAD+TAdHVKOqjBsuH5SjH9/GwgAxGBy4yoqmwHfWtn
L3xVjpuXpmbyfDy2Vuf3b+ntPeqJe5g7KQ3az4Y3TLtlScH3eL7IAlQ5wuux
vsHsNyrSSk5nnIljm8Od8nq8/V4DSsBTScZwQlk7uC7c4qd5DZi29TEya4AZ
+XRaNnXP1IZeTJafo2WcgBEoH6ZSQQPyPql6y54hb186Sd/GyxZCqQa9mE/j
ISxcNMuolNE/IIJyTjtErSf4lM1qeiXHyqYNQdbZvoLIZJtcb5l+8TPWT3NL
DHKpQWWsa4kly4MV03wjebKmbvoHYrFO852aCGhlt7vfuEsdwMiwuDt49r8l
l1UwfE8f4RAO0UIA1yHApGemLg3wbmS9SPnCqfs24K53MGvRYmB9Pj/1v9nf
OxN4qZgomyAC9QgBsrZYuTzu/EjgJwK2Dl/qQGFnp1HAcNDWTRRfQNP7PaPi
t1tUFY0IrpkAFKprdIpcCPJgNnwXRPP4ZUY4H2iiwCfC98q/apWre7WjY17W
04N9gbapoRnJW6Z9OW/ooeoQlKZXANocs/m+6PtYOCLi2P013UqsyevIiUlU
ojdzGNpKFNfGEfCdKGFQKjGCqIS7x/yoo7a2nzWlxm8XKBUF4Nul3cscI/KK
pD8JktVl3wsSIz14JsLkBWV4gfvU+0t1nAFYOffthUXiOR4IuEAsZbx6sBwl
eKUcEFyL9PmnSHLgK13ixkY/VTQsouMIA5jJulrzxcU3Hiioy0+w0ALABnPA
QTOgfqtvAFBVBCbWZYi68UFiLpWOz5lrMYhyf4VaaiGbqD6RYnvFdYfmDUAx
rhpNwT6grqOa+9QJwZjnEvSPH71eUheW2nZmvLJGKvlpiPuAwvTAf0wCrzTw
/I+AdxW1r1nqgQzlWAEU+OGXoTueyVnKpJrfkqjXbU39iiD7BoutcAky0t3O
73uvnUbBSDSTQ17dYODonUac5AnTGC4vc4EG0eCHIW120uLhhu+cjTJhJZqo
IQa/xt1mKlDALaUWrWTSZh5zVx0UdurQh32Cm3/yjXM36FX69F8md31tQ3L3
vZMH35yE5pKTf2yV9bhJwGr2Sq3HuuOz+NF+V+4uSQPSYU4TRbbEF8sukRZ3
aBT3XSmJHFwLSI4riSRPGOHkDem0upyf9F2LrubEp2HYfSs63cmlvU+utIw2
JMyMa6ERgL2IBUsPCDUSHLhIfp6Ewo1ft83vIUyJa0jhbicxNiA2Yc6rlInl
ZlCMjmX2Y2Qu0L+oFPlEb3A/JqyVj8PvwAUM62aB7Y3pqffpQ2jT5syKY4FX
ydKT9wdu+ap6MV42HJJuH1zTuSdABCYmW09NZXYGrqgUL67mQE7qSLUk4mCb
071IgzY5uPWPVoYSZFNyXaLRHKpfyxzQUsCP5hzQQoHd9tDKhujlgO08MvAw
MaR7UFrqVTNeON0z3Dd/dc6d4+cVpwkCysFzSBh6rwLFu9oAYVyFrDfg/X++
9cTfH6cLjnwV3S7b/pVJYXv1tzFMJHHZ4gV/l5QWRPfV/yezG36FgTPDSA3d
bJXfxwFkp7gby4/YHMl5iMrpNMXakaw6tMS/33lEyRCh00FhQPEAOkMwwszT
sKtR9mght67fNMypNrRSEuKPmh2Qyj0oyeXyk7o8Gfxn0vIgej/pOwyuJz30
GdFU3iqTsQ7SJK0gVWx96XlywpSTV/RN+iA6lsd8qw9Z0dH7H+WqPE3qAis2
VYaimqQJd7kWm7MbjLmSG+o4kZyp1h4Q6hQspBa65Tygtql19feGDsqTLnHz
t3LpI3BqfOOD3JG5auueUSdcH6NG+AvJITfxlEZ7pT9znHOwwPBGn+F5iktO
0zEbdFlSaCwTPrK0LdXIgSbajTAAygqBc/cbRUSLwJ0gOeeVffJDvkunWSL4
u2rp+7rN8gxsNTIBvNIMWvRe81bRa6D1SPGxnkjkr9NPbKdHkHefLdgj56I4
5/uLWIOu19Bdh3C+4v5hLYIseIyuyL4pl6/aFx+4VNlP+lhUmJFJZW6FLx3H
4j21pxZ7pNdTwIhj559ZRGuE3h4OsrNu+vLSkokb+8ZrLP0+FTDgreq0CyPG
5Pf1chaH49vAm6NUuLoQOIEHHS/kjsj7m6PErQxNWYbRqDUTNRz/QpJt/dQ9
AXic1G9HqdaMhiajTgAYgPT1PfO/XM2Ainke+EOsN+KMUJOudUDBF0GBKvn6
UkqFV+GfN8143zB7LuC6dJBj2i+HsT1sAGS6Iope69JQxLWl8U47OhzOfP15
YdZWZ8Ku4GtLZelSjx6cC/CZ48u+dTfxCmNGsPFvDoxvVUSUi9m0sICWUeps
DyGAy2o9U7j4vfXiKGIBSUY4InCQbyda4/EyyHuyU69pZSceW5Wv7XSBxEUK
AB9vJlDeGAw5ydXOfIoObPKy3M0S7qnNdIARv1pM/ygMu7GfdOUPYYraEyku
ZzvWd65nwgBIIzoy8D/Vgyb6bZFzqPdb7CPZdlYSnh/0d0spH6T1g4TrhQ4f
QZ9QC7rSIt2fAd7495HubHVfcxjsXJrKP/GCozf0n4AZFbaW+bI0tDmcFa8h
LTteRsymzL8WRI4QMAfij2z8J78akEGSy1WIIJiGvjE0MasszbB/coej5t91
eOqVV2xPAzfTscaM9dQ4Zf/hopC8t3i3gZdA3qT/ueDoXAQ1BYNltCKGLWX+
jDETE2L2xQOK0EDvXTcojOdXnViAKYwigVtVdbxDavXSFOCEun0vdShjfcVy
Mv+9k/xOOxedlEIl3e0ErkzFUR3KCLU3LzZBD7sQT1/8xAk4xcc5vbiTAMtu
Y4AKf7Lbc3CljNPG/wNepfDwsdKoHs2A4Mym3/4lqInRC6iTwGNoNr+u8tyB
j4rHvWrhrKBTyWIqA9K8AgYYEHCk3lDdS6xSSxFa5CdEJShfCKjfnfjbgwYh
h+Di3XssilG6GCIxYoGU8tJECXcWW6wWbpy33pV7bnkc/2Xw2zuBjRIJd/up
q8NPPuqOX3UR5srPJrRimGyV6IqND9C1aGJLNXJBkSOom2DKwWZHKcxjpLme
AYYl/y5ACKIln+pHTsa3vLEk0RJTa53DCBcvM0NWz3ZhH84mtEl/UQ78tAic
L+tNiJTCs47HNZWplqPOp/p4Zm8iI005W0SC3FLzTJ8oWa8VDUa5jTEFIYUW
XRcm8w8kS6XMEnt4Y95MDX/ZM7MfXixbzhPInKv80HWitMrXvuIJGHffNohJ
MEq6+Ks6JhayCdmzaTx2FT0nmLDGYxTsihA7v64S8brAWBs1vfkJq8wPORM/
CBTDf2DHmLeP5yM5Fnbs7yPe0v4mVuLrus+5FOl9Dwtsxvs+c91zxuGArQge
N+EE+2OCndSbdfUyllHaNq+aQkDb597z14Bj70rwVR1fRHlMwvO7dCJcJkjC
Gr+yH+64QAStaAdi5NbcrnwYYfBCdi7PJItwuONhWp3OrGutnSfYIai9LhIo
OLa3A7k7pK5QKyvrYTorrxkbxOI9KywGdhidSgm9Zqfdhpp9w6AHY/+cxgoC
Gv+qmFjPlJzc9B7FNOCTRaehiXPIxJsrKA0qixOJLB2S64NTArWApeNaAs0k
r8bJm/fdHYBf3YHbZ+i5FBd1yGOznpooM3VgVh/6M5tbReip5N4eUrZa7gNG
iswmQa4Tv2Dry497JnrmgyUCY8VJcQHJPfVU9JS75jF+T0XxAwnoStuI7FW3
dsHvkrtH8+qZVPyb8lT2bzFjHuMNfhRAwB/3O+U9+uNIHgcoDWYTZSoVnL8n
DJyGVHyRB7pz5uNjyipJ7iERBu717cliw6sOBsp82N0Cj0B47ZF9HDo9KzkC
rcpLsmBcTT4Jcq36qEIq2z0TLDcoaC+JpMlvuitNROghHptsVHMcAJqTg6Mb
c88U1ik7taRxtZo+hsun/ZlDsEQwLKbdjDhdIW5N4pzt/n4ZQQXbnJK8pURa
fpdR7zQS0u1XPlvB8yqaeA1WuaTeer+yLnumIM+XN7gfUufTe9r/f3PhNZh2
gQRJt7QhtUrkvVX7PEhYs/5zxIwmQnZKmuveSgdjvUAkdQQJZ6tyofD1HQwi
O9Hbs1AswuKoC4T/WQyp5dR16+FUdECU5l7ZFJZ6kJXx3NyzX8NSd0ZtcEKd
ouKFTza8G9AVNA9kT8UtUAPFi9+/H3bsMQSfp9/g0/Dim9k4JN9Qfe4HS1SZ
NJCqBLOXTZZCXoaNrtyvG4GKFr1so/G0NJbp0xpaxqpm0a/id7QbefVUS8Gs
KKIPYsdHk8hfcFaZbvOx89Il21WQmBVmLZTIwUSsmpZfQ5Fa9nNfJfIbk25W
4OG4g9Yqf7vAx4NNJ2W3Afe3whhRx3uxdzhX9I/90C/YJNf/rkduwBxeVubc
FKetO8+vY3mLKAFSRk1tJF8Ds9C/vt0dw9aqfRHQZQJ37/lXnvBAHU1Q485T
iZlqA+vi9ZeEXZ3q9hDege4icx3gWa9ZB5BxCZARXfiagY/aLw8ChKKdWJNg
+tRglWM2sAkpYOJK9cd5lxrc7lf3uXCBSCGIf409S1nPrf17NxG5xvd5RQ/O
1UNAqd358UxV0rcYkeQ8LKXStBlEXNoaARLzWZwuxV5emS5PdyXxBvIDIcda
2ET5W1xGycO0FD/pPQq3Fnukk//F0ZS6UYiM7a155/dPREZuF6XhBUJbKjsu
S34BBHrW1xGP3TDVT3xJxt0YxydhY5jcMG4TiuMhipRH1xGz+bQp7MRwgbGA
fBrC2dAezfHdEOEZp2naQuAYbKPuqnWzDIWyFC0puNReuoiMFTQ6yjBq8kb6
PeYVX2+WsSRnduABxdutInOz2oujrt58KBJQ/LQbh6TakSg2hOxa2xMkcvDU
heQsOnQX40D4aeilYUClYuPq0/GDVM9vdEpMk1Vh2B4OjiByPyfZiPe0mQzI
sWlALE32BHs/g1F+jqTOaxNuFp9yYMQ29wN8V+3lI91EGB5a3pb5M/WOyU6X
v2tqJYRpDUBxJ+Ye+1mWuMJPf33MiuiX5M/lWWNlbZEMZ66K5gXy1/lWvO7E
3L0vUPf+Xen3KUTuGm6tTueomYZ249W2eoBLTl3HbxEXWT6L9B9cvsYRmtks
3lMgE80szaMZ4Y3pzjljz+/vU7AwD39pZKhUEzVegdQUM4MlJg/L6TzbFnfe
2Dlgp3CEFVuTQ4nDATuOPDhJeMGVuFlPxQ/Rl2EVGySl2Ao+EdvwoI3bheS8
+PFFgPbf1OOtHsAH8MSr2w9anxDhPLmEPVnNh7svVMfd0NmcMXVZ+F7g8B1n
jt1JHo9G8VxX3kIzb2bw4nW3hOi3WyHBoJ1VDcf8EjsW9EjIqVl5XpfFvpRy
C9T4dLx9Bdbnc02HPrq7ijKO9M0lIewt8MYHjPYSAWEtj70B5vcHrkUUBwTj
uF2X2UMyPbX6l2OUKKHvkSM7fAlkpbcPR5Nd0oexxDWda1gTHLS6goDgP3E1
7iwTUqweq3bYfu4JMI+ziEK8HN1JRCHLMPpa5RT+587vjpVAacicYhRGH17w
vvrRueamLAbW/LKl+dTWz9jBGHL4CMT1BCEV3PlvnwIps2doo1QmPpD/K6q8
uFcd8XBN/beDDe0yIiG1u9C5LGHsrmhQqcWSFhyj54CtHo3TWxjTsU/aXsR4
AD9lQuW5uTBHQs4MZZY6Q1LZkIhfvLDsvNB3Nc1BcGMFVDM6DjmwziWnk20p
VjErgJCintVI1NDqiCghGblQxAeOWaRtn7LFgjU3OycbvxnGPVcfHiODjXs8
LdifthmwUN1B06E8cDDa6lFVuBpjmBNagIc4yI0wQkDKAbmBZ1VtNfd8UDL5
ErHBaCCZKccKPgIhfdIjs2ZziULtGYzMgM93h6BuhWZGYVRuzXAPUZAWjSZl
G528ucKOE+3MTpvkzembRxjZddHu2ux8DTcjBuKv9kU8yEqcNwFXGcQ1X24K
f6gtJ4KaWiw+r+Qd1TSOSiNgSJuUHzshVeeRTD8Ljhws75P8C9icOyvv2hjB
PlQSgr+gmZFUxyDYQVZXerwq5exGFldx1wiNUnMmVKUgrOZ4c5Je2l+ns+1l
/6tOWM8lIqHK+eSidcb3pWpWxNwnpEotUtio7R1FkCaNztnyl7A4DaW5pnTz
rOcsrQp0CRdDV7iqpI4tGp0r3/nAwXpSyT7flBwceM8ObPJg2FU6U6VSjJ9v
7vOlP6Ez5qCoIRu/l1tpYvECIFvDVGncdKIcw+WB4BpfOPpOmCnd2SoTVmy1
/RQIHTSw0n6jkJ+cyUDpSgx9MdXE+1LU9Pg/z7qFCQ0U8c0/4LeiZR0Xcejw
9rH2/6JZXcfFgYmBDCdqsjmhXqdcXa8maZ3w8QAGyI8a0MlqLWPwUZasQH/X
chd4Uj4aDob7og7iGbfX8aJOVZp/24NncX0eNxPfVkivPGqRNULX1KTDCZRN
wI9Z2OWcsJWrxnb3xQGN+V6RY+HpVPO5xznrpbpipRf5nvIIc/xn5C03Q/0B
LLEGRSfWpfbeODXV+6NiJvqZsAloa759nNi0XV8OOM4Y1t97UCda1O/+VWaB
ZGjfR9stRuYChS5a4DszBkXliCHsZCKjEW/24trqHrlsCj/n1gSuzBwFURaG
HpQeLwnPBlFnHYULF5lbGo7J8cZy5AzPRhNoc628Ia4z8v8sU4jDCK9+RWlP
/uwCx+wbs84QGbZpEWc3F6BoaJnDUcnW0WOOw/c6JzCIplJHXbrITIxEb4LZ
lx4FI4bO2aIB7AAqP/zjOf8CVWfem+/qV8+bDJCyUO20UlSqpLZmY1hYtnA+
VFkrwt0bu8ho8hmJYT9pmQEhxlk+MvNxOwFz49FFtDAbq3c1lFoIeFgmq8Pg
1YQkET+vRRY5pp6qEj+9Q+TXLwWt8XSVXfyY1IMp1w+1z5FjhwPWarMNeyiY
Cr1G+eKNHqDctE28wT+DV+SJdx13pP2id+FP/V9YSeFjmbR1jQ436tkb05/U
DPoYmD5McvnzdTN7zObV9vEK0Z8r6Z99Gxr0hp6LyBIfYuTL6y5xj/MGAz+T
egM9gBN/wXtrd+Ec+0AwtnYYOrbqenUdh1S7+YYRRCNlLsXoBW5nIJgNeaXx
uq5VyJz8ET4JGaVh1Bg4M45Cge0KySluqYEd1O+O/o7/eECdk09eYyS/IO+o
WT5qnQb8Rl6bnwrI4cBjeIiJcVnBTkE4tjc90PFmrsQFYI5RynPK3xt2P10a
M6Y8wnXlItdFD9p1mJAtO7b+bVUINGu0r90lm3zA4aUmY9IL4f2C6Be+Ms7S
0VX8FCw7/Gfs4KFnPQiJr4loFCx6d5j+pmrh5IYW7Ebtvo9YsrLQnAIHa6xd
HImohncLmBIEKAU2i9+LV+2qERZ7w0J5q51WXnrcMtDlxcIpEz9w1CSTqD3D
Q6IY/vtdBzPLaRiSXoIHI0snpjjAg0MH0kPsVQ8wfJDkCZKMe/UWLa03c94S
/j41JURB7Edi8v6ocJ1Kavg6lqdJUuTXRVLrFWdlVTK2iZLHhJyxEe2PZJVy
EmGC6hQjzwBucalpVC+ath9737Nszcbi7oUw+JbcKmfyqveBCwg50ZTTqO6y
Z5hYAN+dB18WubPO2J6bXnSSj0N5S7xBH7ttdz8zY/XrEQarhTDEOpLq5y76
J/0HF0bKexWA9ttk9/Hrt318i8Z1tECZPX5OvdFum42rvw5kHH8NenTspWjC
5tvUni6L3YtLUkrxNceXvmKXXYgJQY47xvKEr04tvjp1F9OpAetK3xO/15v+
vb3/9hhMfbeNUogJS59Ih1fIL+02ACJcTz0VgXjL/quByl1i/BbwoQHha45J
k4ArfUS3WscfLaKKkeGzvpsy6yVD+MQ1m8PCIAoKzUuSzpC9vFGgoGDib0bs
C4t7xHvE+qXHpCjsArrx8bMh212prlywckziJt/ekCN8VeRYVsZcaIIm06+G
bgOL/9PbeNOsyNheyqNKuwfQDNb+1o1K+2sc66x9ia6SBvUSzPuQSJgeuGUa
pIntL5bKmDi5aIrw/4/qP3MbLR6PYGoe7C/pNSY+s85FAw9trofsj7K5RG7Y
JpSFt43cDYm52LrI4U5Ixa8ig/zs1ythVZ0W/4iOl8IHizl+QR1feEuLnJKU
bTpdXVj2O717sJ47/dxOxFmN7EdXM7GhCoHGmyG28e8Iexita/oATWvf8tub
grjskHrdmZwefeOezd5dMfvUaRLvkADo5Z8reK+QNOdkp6r9CialO9HYxwox
39TEK/qQKVGx0yLaaZ59RdYdtAN8oW+pZevQWhzAXSQJAGTEtZ/XNzGJY7oh
rf+i4jyCR+78EoWK8yRDF13xcbc94Lhwl01Tla8zQsCZ/QBO30zRJhPviF+O
qB9f8lyzCZUSl36Vp3eEgwbpeEfrUg/dmEfPZmNVaAwgi39SqGO8EPDkKO+4
KY/JrOCp/oNnyEeDFlr6KJjP0gQzNyxJOGdudxeitQ6vR+UXV++9WuJBVMYj
D3jI2s1W1sX9fuMCW2O9VsRHHA//naXLavGrPdpV0ZzhRoMUc5MS44WesokM
lo59qkdf5eZcrEVX3AN9cpBjTUT8+cpJwjlLtRPKZYCySrtUUB8SyImc39ek
3HKacU2Sw0DFe2U9NcAHE0FFBiDM/FANyKWIp7BuMw40r20xfDaUDJpxpgoH
Q+QvUJJ3ytV3BvvdxS3CLTK2wEoOzovliShWCmUFFqiAa+mYETbXecbWao9b
tDlS2P506mYu6jxSkJZiOiLeHUE8uIx2oKWKWWNcY+fgj+5TgeB1OtGddw5j
FRc4V6s4QyDl5uGR45ukkRXMgKjEIcVjdoMbAPvvfikssBFZ+H09BBOvGzEL
m84BEVo/6JyI5J4HeO0AKCbkjqZtmBA2CtLfJWFjas3G1YmMcdUrATapF26Z
IrrHYp8ykxMU1k/pUxzh3EdqHOP26lAvoGTH0nXMM1K1bLz3962QC9+UOzLx
5FzXGJ1k+Jj0rK4c4+b8NWY/kLdbg1oQxsLXeVXzxzklpCcJiHEOIiT5sN+W
bnUA9Wmew3L84qklc1h8rGpZ8Ym86wZdwgu66bukuddMSN2lWlwDj2fl6pka
I4dDjhkKNUazxtCVXyxmKX/XpMAlt4KPG8DtRZ+QfVdLE830fGOqqPxDudU3
yDCiVFP7b5ZEjvq10sOYCWKXB4H3y27USU07OMdQftxhL/bd41pB4SzPng4Y
5VEhAYcKqp8uyvo3h5sYYEyWerpLJR9nGtRwjz7IuHECCx3Hnm/+146yIrxN
MsZQogodak1YfQPjww+hyOxk4ug1WPmr1hGHYQJlNcZnVgH2Kx1G1xtFH5WQ
0If5SeWurj2aJJDrIeeSUFfsOFfxKzkyhGIjGdqYTtiXH5IqmVndf34zTyuY
B/syWUsC63WcshEB4NshWMODS9yDOBfPlT3C6DVqWh6sfDRTLR64yAz2cJkt
UQ8oiSip7p6J32o/hwMS5URYT5g/O5/GziOz4OFCckLBtgyOTR1e9ZzzidRr
HelJbHbSqrjCQ8M5R2nb9yrev7EWz+itkrn8RJ8CkAHx7sRyhRo4NAA0nfp9
8NrMfkP+mb/8Cy6rL27WFthriwjIX+GvTM2WctGVUphgiT3PIZqMgs8Cctgq
mCNnullnoSgurlFejXjnOCtzU/RWmIOUHrK8hgEpxkRwfczeAdS7tXkW95Ji
VjHaPs7lIoWJTuTqeJH0F33/IdYN5eqChUDmFfXesCsWcRh09KBNvhWMFraY
QSA0GN6RMHdKUrFSp9VR17FnThejV9M59O1w3popL0Ldm/PwsvkXlvA+bwk/
ZyHNYVUdgVdn41W51dgs1fgNg0Ey7vn2vl33jtlFY/1CrpuZau/xkfX2Nw6+
K0YmKV39bLCbb77a9OrIrqGvy2o6IpcSYBRB08fAdZEjR+dH1QpyO5Wx0WEY
5H4P3zjYUgzk98DFFNGTDRiikxETn/Hvl9fXO242zUHuH+aQlg24oDTOAzlu
dMuqB2C1331Ihu4DL508UT0VKLSvrmqr/F2c4UgWqVfz14EqWnl0Na0NucK/
vwvL2IE4Hemo969osTsIWBkdn/eurdte4AmpWlLp/CWs/p1mWXXiZCBGeuUD
GNYvn/82Y/98MOvJeEkuPLYqPqztJ4NeBKXCpxJkOJQi+t97hNqQLmx8KXG9
HwrhPbAbVqxvYgSw7TOBTBEuW0bP/yxdxktk1uxAJRo6+Fmyqgm7yOo2Ffm6
7EsB9BNL4Pn15Q0w2+h+tILELwmiesfQYBpTC+c077NcEjKuq51Kj+CGKQML
1g2AANROv2beabInCZWUDhOextMxaIoL8oznYEYJ0KhTq07YbtKiHn/ZJKAC
nF22zSmDHC/TVEiLQREu/I/A7MT2g6/kTMZmpx1Bz3g6b70vkDBYZsZrKWEr
wmVbMLp1K+f3RDtWNQJv9DSOWteNWYNaR39KS2oCtVaRYxRotlVIHRPP0QH4
/3CHoHnyhaa/1NBL13CvbjlJWt6mKfOu44esMjEzOJNnmJ8OGV6ghmRuqmWX
IDLrco6RnmGG1s+e+zgAggNzjSB4BrqcjwSgWjjyBtKZ5cUe8hQXUo7zRO9p
QX4ZP0+FUySiD7O8yTZ/nR27hGXBjDl/EohfYMxL8PO3cxIdEX/zOTw+SAkV
CHBzH4oooWb8wvZ0IsRaZCObQ2jgXaHmttPvzee2zIDtj90KRNeAcdTGJ+xD
aqltySLFqITvkxUbH3sa12qRQ4ZCEZsWVKay9/UgxAAfvN4TxEwOfkawdBTz
LQIhpiqR+Ro8PhTsI/5p+JYAiZxh0J9uN1VES1WyiWmoDdXTrXR4OyBjbBJL
8CZ+QsES9K6jBH5oh+XoMQcLJwjfwRUV0h9BcdKXlij6F5n6gtuysFAeW6Hu
qr0fchXsaabdtMnT3mfrcOAA8lDOHTd4XBBe92trQyY09LT1Uh9jShD0a/AS
r0FymJzK7zdzE4t6Dh4lEHUFyY+i/jA2pREkEJAFDTiXxfkcva4UeDIkVF8t
AggZ3A9B3TkAiu41nWBeGLAnGv01GlVUV6FDkv0UlffQt2xEhcaTc2NBlBpD
AqV3bFHcQqdBSCPXR2HeyIhc1v9oaMkDLLEG42DKAyEmoCHRTbdSPhXXqz9O
cYp6ObgS5hDBanHHgBO6Kxn4TlZn2fprVYP9xN9CbMproCH8kC7JwxJRWywl
KaVnY/6heAmfbnIeRH6OD4TTInA29RNJnfNp0jmyprXxqlK+1241QNUIdKXv
L7ni0jpz7Ilk0bnqoHw74j1ov9gPfDh9cyB1Nb9XNV/B1uTb2ahMSSsFM+Qa
hxcDZeR4uO3hQUW/cAsgEGmB5LwreIWHW+XFt+MKhuySjZ76DKZCgeOgGWW9
RCBs4QrYVdNrT1gHVjXlrV4VFao9Md/fdkBeQWhrBjYPONwmVs9S1azMyWIY
TW9KWLHhaF2Hx9PDUEHJ20spAxdVZ4+h0ANteAFyJII8s7U+8KPELCsG7uDL
rEimCBeNTBXGEKGe8/5WH+yPhcX1ee6O9x4BKeOllWrhHWARMZjyu3cOtIhr
XIYbsp0aXFfHfQQqpMv5PnmRXb/HEG54xDk60uGVVC0Lyi5m0ryx29ifWH5Z
qNEBoKbGoXVfi000UjM2uoNSyMv5xw/Na5jrBV0VZMbX+uC1H1Nk7DEltuBI
ve2HfCATzFWjNfmsZmW2xL5T2Gd9g1r9fBoMbFHFHBuaPRdQa/vXNwfKwb+n
q3hGFlbeHcgvH9Gs7e0h+tfE60sRAqbM2tw+0eA1oHThGenCXKY4hzIrfnpk
pTYTQmrCLhHvxzZNjVchT8pPgvHmUwT9paEGB+/5DpAF4Eq43e5t5YXXuJk6
+kCJF1+u4kJ4A+y70X4FKMVotFt4tHz6cphO1eS5bAQRuDFmWq8KQ3SraPnU
JcO9qnsKkWXCfD+InQQPndD/B2asMq/JBfRPoD5cQ1QyGE3dmRvGkGLiDJWm
rU9Zo7rAvigVs+fGVEvJPqN5g8L5xtXtloh9nZAdz6XCEmeJw0zsqLxrVzSz
7dAC651iRvfWOBb8bObjhmS9rjAtqgaF+szW2vc66xciQCviY4dsyCPjSHoM
Xz91IEnU1OnEfsem1B6QqpoHegChYJX/07Npcn3Wh7UEWHkKyRegsVa1EkzL
4GntDbuTIDuMm62l53tKVdI8jrronV9wh2ewH2+kZfFbd8neRxjGU7HM7qFs
5nmov7gEVc3f1UUoSco1iUvQt/AEbGaq9Sb7FWKcXSjYni1Fmo+hJ0OcoU8L
euouTdK/Ul7kpt2qPGNDYExMES1ebsABZGpwG1sJg6eNI0QfDijYCgYw4PkI
1nn9QQ2FvDSU8uHFMNPeayLXNvwDSxbGCn4YtjpQoGw4oijJssFrAA2zFbgZ
RyfDF3MocLArHD9H4p883gyMyCFi3n1fY9sjHgZKD1CZsZjOAL1HkgzRiW2q
iTxBL03Z6px7Drkv04Gt5DMp5N9cTzDezLw6jtgHxBHjk396a9OpDLZ3cJqu
id9Io7hXGtmpGn41IZfzDgDCVUiLl1wXhuCPZWIMGbF88rJqLMBZcQaIkqw6
K1bRYSd2as2Q/6ec1VKTc+JDGz31aNLeb6/0jift7a7N7637nBSslhvqx3YH
wAEm+UieTfzOVDWc3J+XYYiA0snyV0NhcztwDVR9Z1KXPbBVKISlENioIZWG
0nIsefbNzvbCK1YJ7KEHGUl+pLGxQoAu/6KBqsoIwZQUcn7Rd1YhrQowIyZ1
JgSMI9JHiPZB/2bM46I1Zlq+BuBpSi8PlVmpjMDcu39/csodkF230DFoU32n
EBShhHMC0RJvNlk8D4MDtIF1d7PiGYEjtB1giQRu+Pw8vn4x0L67/OAviwO5
GyuShTIwlGGVIgl7CrrZqXHLjTQW9nzHnIjLjPETMF5jCQaPGk39ANwssLq0
OqKp59yWyF88n3Cgbs2y2XDq9SoL+zF3TE+9UXrvnuol0cvxuX89vzi02XSD
4pYPp4aVVj7qiDVYuiGbWPvUWchSkF3xjhuUqOCrsN4KPGNpE1RyCRoTO39d
Bz6cU07azrBY1+qRG00oZib7XOSPoAYBYKjsJ66Aqd+Gvv/XgerAmTP4fuTB
qBrp3yIlB2dbDhtZwpwaXsgsDkduk3LiNkOtv7KJzX8W682PPvrmkBOjuIHV
y6S1Oct84bLozfVE/czgPX4yrP+MTstU/oo3R1xHIw0d2/Ou7E7wIsriwFKv
UVx7jobaNi1lQz4zSNmiMLm+DqfHpuhu7PPdi0vu9Te+JfJSQqqqoJTMFm4R
FjvcO0zJ79iMTm7p3dVdKP2GRenn4qrk98nP6R5sxQn2PcLLJ267JQnJLeDA
Hi1YkCnvR++kQMFF4KMGz3uZ5G7bkVEMtnHa8Xb6SaWHDoJkIqAciX7V4eVh
JMox0bclMdzBpfcKTa24kDAbuw2wP/WILMBVfuoGovLkiXq+aMHE48wDQaDB
arlPtxCHcidM611HOHmexwXD0M724YHxUx0toOmFWLWzGhIeumWjE6lRa3j+
UaRiwj9Fh9vfl9N5BKbPObjQh6oaO7gFAwTrAqBhhLSsAb8fvFZzyE1hwPyD
yeYfpw3VIOYamKq8BHloZ9GFG7g9X7qlSx5Ek6xQbSbJoqTFe87nphen84E+
k6jHAgdMkU5xRPVjm8ZVmgteyWkQKiEfj130rEEOtxvJuk+eZNulYDcX7Bq7
vhwP1s8CwnUI1opN2Qrw4LidkHCw3xPtL4PBWUiUsyTPrA9AEQkI4QPWL6VP
puY0xECNHF8mYc0e/sNNMvUfag7Zwlbh1DlKMGjg8JB1Oax8fIJjMyg22ZLE
KtbqdooZZ63i6Ncsa3DbnAgKFbcSZ7KDyrMUY0lc8X+xCgFSvJSlLJSbKWQG
XDKQTUfqLp8e4Rx+Aig4hkeO3/ihHqRpRlcAoUqNfvxAlLdbsaGb9KpVJy8p
r9xYVbMZmQhB6YzF5hWXlw4RtMRq6pa7eQoo+vNjELqEMC8ZkSBOgTCo8ni7
3gTmeLbvEenv+ScIpZLVhqn/ydk1wwG14x8hMy8smcN7C79VLukLOwpPIHdL
Dtm9OSoAkqWpp6cAZeTBumqiDkpyMUh5xB9osRn/i8L5fdWiwpET6qIy/o57
NmDcjX/oYy0ymI+ytEXFyOC0nMh/4lcQNr7OdgQ6KJwsdY2YXaqIxLZY5xBm
U/MGok/Ww2WuMkQqBhxU7dZ+geNyWsmkxdpVwApDOwem+BjmmcCrsjXdZ6ei
/g7oHCsfBkz/qr0BrjWPRbNR/FgtnuvJqft1uVjsdLT3grJssdcw1sJJnorh
vPFec+9Z+a6i7rdXTYqr3f00Rzx1ZgMwM82G9UfsovdkfmT39xQtNoqAi499
xtXZpv6a8spcyiXD1A0FWTkSzKU3lOrbKjcA8lumV7jwrHwnXjI0vZPz0Lgt
y6qAIdODHOzW6ymFyo0TgghTJM7DYHWQWH95SHo82h4tVVCSqHttruyguRqv
Tc+6rLmmKUtJnEgeAXBG9eKrXl9dR20CqCOH5WEMPulwqlAu1QfNMKoGcIN/
Omba7/Z8vP0J7pqh8Qt8e6HvCSu43Ee9D9M4xs1Rq/10NTk/EnmAPJRgAAdi
+UErozSlAO0VeLanJi/+VBhmWZ70UQlEbW2czqxYlAHAB77ESpbDnlSXZZ/E
dMtDkqhvk4o1SWGbqSlLtxJrsi9UUwQp/14jH8OE1di/43GGZAvu08K0dFbd
NKz0SrB74KVTyPYvU+JHBRvcw+Ez5PC8Ma4+O9Ht+4SOoAprjkTYuP8/3LiO
r9O2LBcMPC79KOXZVVfrLOJWgi6l+XYkKn2hzSJnSXHQB6S1G/RfG/Z9jKV4
SJ4mnBXriXVLFMH6sx2p+V6vibva7zQlaLoEmx38CFnlkC5Nk4jSzrELY91v
S21KHMFA7bDgbFnHty+TjCQG3xVmGBGU/Lao7gHxbPAWj3ToVvQKGY68FMiz
S2BTTQXDaF/0pSSQ3UOlKnnm8rVXTRJbTljhFbQZJOixTvYI2fi9Pf88sufb
KjI1I0iBVTeWRxsRNspybckcpcpiD5mozE08mIYR4LvtSCTGnQujmrNMq6U9
sAMkkIf02aX8CgZ+1EWOMt1omYCPMpJ6Lphw+u4IcFRHY40c1ZW5Mv1mhaWu
Vl5+NhKqPvrf6MTRD6pYqoC9jcmtDxuEgtdpZYwGBSccPKjF2L/tamRSHDgZ
9R2FoWleHGNaAK1+tIfcs7BdGvrbWJNPDoRk0QlMJW6ScWl213XxOaW5WseF
ewLztQ6ayycRaa4l2gKti1k+0ujrIoW/shcvYPy097asv/DKViqHBUrn70w4
LNcboC6Am+WcaFstWGUqp17nMaKP94egb7zSo2+gkHv1lvOjOLWJ8BWn2p1a
ey8PJukhy+cEMJsS7iuWQ03iqqkDwmW51Sfh/G6Y9mFnuWrGsu5LykK/X6Kz
y4WoGX2gvxdEg2ofgJDthTz8lRYLfFzmWD248HWQs9IsFhG4yguoau3hAvcP
sDcgmK7r8S88STmo0v8qieN8FdMaLbqeKvZ2seuJ0hiBdOR7e190QILvBAjx
+AggJH6L8kYpkKX6yJmACtz68wPpNuaB6NsDm9akQ0m9Dccqtqct6ScVQkZ1
D5ue87+OsQ1IsVOEGWMhE8nR1ewlJ94RfsrJVQd3HPqBiz1x0io2MVdpW7sX
UKs2uZM17CXE9H+63wVgSAhDP0fkXJi9khQZ/TrjHjemw5sbtel/+mvwCjwp
G9314t8CTVv8WZioM5tDE8koqVS7abZOd7XX9CyLmFGiVYTq1qvKvLFJa8uU
5XWVW1Sc9kOD9C7lUKehSLrrpLkYjTwXZIHUurcFmsngZHAuujnpH5rl6W0Z
0eQbgAUFmBtGPc9pdxJi7IsHyyCnGrKpm1zZFxs1/9fQc/zb+qkLwv0ATqT9
mS+5SeLuXL6e0xy432MjLmWp6wHHEhLZJY7TrPzkjy07Q2P9HRkV1Lif6MqP
iIPFbaP+y2WHMIqoumTfyMjPGti4mHpImIIg5gnAQt35JrqQIQWIih1HvJ/S
mRqP0Q+PqdilMyMTmuucr9EpOlshSa6SKrjFUm1gJ9RGw6b3xjjegHxCtkPG
HrG7JjRXExtgOxxYXTMkDxsKkHsD9LdROZB0k2NfFmxx33bACrj8SeCIyO2R
vWuJGNxs6iCZomuWIa4WbE3d1qrvrpEtk+qa6JHbFwd3RZuIEQonNPDw6BPB
DxFRzNMDpLZmGLDoA46hXHLK+gJM3su2WEnGpssYvswzq7+MxMIJaSOlzHcC
TJXYcdXEDKnEoLwBfgcQARkV/cE7l8CbIdSzIYqodQhHA5zxEOgntR0qRc9+
m9rgm+fBXGp2+CcMzkK/DzYYbAkAWZTbKStT06DW6fYoj9LV2Ov9XyfZPN1n
7VKn6LSylTRVyNWUdWcghgp3JQm8x8lDcTTcMwCGTkLuderoipT78QPvHQqE
HvqYN6VMbu7rhPC9pjFDY9qZfzNbm23aYkbQ7wP2TfWai5pUWJyvq//wG0rh
GAIcA8/vfkOvZWeHvy0YFcGYycZh7FW9/r5BF2H2wjTpqt4SvDnC2tomkcSx
zIckWjqA+omL5dynht9ZR8BkeJq6aSXznYP7dgN/mQRij5Jn5n3d9BUEXdC9
mz2lTr2TD384YaPnuRJQHWBNgf4poQEN+RInlks+vUHIswHRxez4pCps937O
Py1yaigNTKVzK/aKY6IiyeNhzG1HDyWUvGAuvOILjDePss+H2GYe2U0eoYb4
031guEZkAt/+TmQzZCCrZOmOqrXKpyalc6m9pb4Hr0+QdYHVo6jAtDQD+0pw
YwTdsqjdY7n9Wl/z8pulWKh2uqUjdC7vBczVv0etOXhIMGd/lqQwf6j+bcUS
qikpYKYRx0k9Yi1SCb0svLWLQkY+znSw++wBhVqEjV3u5ow+kI3Byb3Bpsq1
+6IACZBqUUbYB0j3XSCjah86TpIci9AKk0zeS1FV7yjaDiNPz+ZAEJSa8vHk
k6Bdfikmx3nAmpRfg7RW5NzRRejDiEwwojUoSMphYY6FlNAFlBnUwTtKGmrm
Y+zHedHqhBfTvgXY+Pgq81D+Z6h7N0cMOf2EQIPbSm7ifMEiEAP3M59FSm1d
HhJqt6GQGRaWKAQtNebX/5/6U8HMgaCWfPWVsme+/TcGm9TX+fvy70O4T0Hd
BitLfgYpqzC/7Qt7mgVLRAPTaTkbci1p/C2q/FJ/65pIk+5DpOvq6eOQDqNL
SbXpnYElci00leBeZGp1/aOAPeiY6iqvDtUC5HB1bkYfu+DMswjMHcUHjEnX
uIzcnWBP/lt4D7wAzBP+rwg9U68d7L+ZWSKO3GZb/0OTduui1sFVHWGVLb11
oFknQJMIUdFJOVznJlSngSi3mNYeWnKQ1hl6Ofk+OlQjkmvYhANoKv/4MUxn
qee0/Z+wmjx6rPXVZg000L6cUIpP7cwazmjUwsX20BgsK+6LjZm3Wg9EAHOx
pzQKALeNx1RyGx1LdmAKUZxujS6Rve4Xk60LG9pe6ik9Tsg5cs8JvbI9m05l
yI2UMQk80jNgZc8cftE5UXAsPLCv+oMVz55PzHfNoCVDvIcAptgq9Vu6Q2Vo
N4SKM/7k18kgsVSg71m42FTS91OloO/jrP3UYJePyV9/d1cgoKZ4hfOwWMeh
92L5ngENsMuO41TTUpRM9JedlHdQ5Uwxa0mksqk7heS7X3iUnyqyGPff2Z+4
KGdXx58ZSPD6/dBq9ioF6B4P+bLeUQR/+jxUMbYLd1J2yToFl0BWbHJfr9Cx
GB4/u/0y5klPOd2hXzGB+U0sdI3py47IvxEmAy+bZmxgDgzkCw2POaYLxa70
WKibMtF+LFClnl0KR0796SRFEVwSxNg7JcQqy270AXQVW4PMIiZNdL1wou60
/FZKpCu2gk8sLnRw3mWrw70OxZz0NnETmnEHXuNAGIX1BKvod1XQJ2fUzwNf
znwOQD3srJLWTbuxrtzY5cA9SVjrZxFSzcnOJbF+kC8WXmBoiib2twBlSCvM
oA/1DZ8nJgGVzbayc+P3CoiNQh7+3g+LTsNR5qI7wNARpj75riHcGGNJURW7
8yzsDyxxJIsFtVW1G9FJcv5tbLAdVMk2O9SAvXohfTwXkrNvKcPxoXiEh2jc
yBfjVXF32XhWEQD7ssvIxEXaXFKL9QKhePWr2L9ThIIz5Hp7D2MrO5/ocsWy
VN5gzX8CzewchkR0m6a2YhToQMtBe+E7Hp/fDuPPPZcuL56DEYSGQVJAaEEo
jW0Nivu8PdB8ljHxQDEuCCgM/AXYfJ4Joiz2tDNQeIvX9kgoH9++JeWtzUdD
iG7Gcm76F73za6pAV65HNV1H3q+grIl8CBD1VzLtJZItffcnhog51L1cQ74I
Ye6rWdpuXE4Mi+H7T97wy3p4EUUnPMxjkVUfOq2IMKy1gFKVTYtsGFzVH5f4
dWtKQxP8cm5M1rDbbOoRRDFlNmCK24LJ8PpndQO8JUO90fx6KTP37eaC7RJB
yOT7DxnvCLmxIr0FuY2OpfV8BPckG/l+K2xdFdLYe/JSF4Vwgjfp2GECX5qM
xLUZa5Xon2047m7wlDv1UpU3dwvpcBAO+t41TWaIK/AmzyDOM5V+xE9CzH/7
wIcY05DJYPIF8yO10XVHdlzzIaxVnCtEEeACYgAK5jjJJ0s4kM0psDDWGTro
DJD+yh7O1d1Lj3TbgAax4dGWW+SJxc0Seeuy3GRByIJa3hskB54eOiRAMBF2
ibbtBVZBGC57EZDSfUdyn8870r8c0XPGiePelb87DWKMh4GWX82BvQswUX2G
wlbweBMXUY3thbQXAQhCQtWQ+TqinAhoJJjlorBTiWASd9DZplchiwz8YzKF
aiAyI77zF7kTXF8vYDuTLvLfJU4HMuaXvpuA4K3nnxGaXyoLjZ9J2nwAofzP
czU5EuZj9kiZAJxpUCDafYfC8h9YkYVz3MTMak4y2e1szg6wPDIcSEQTk5KI
TngXVuFA765kXQ5eyBPAPTT65riiUdBBk+nAXGWTISR2hI/CiN+iHAN2w1F0
MnDfJfKAnhZCU6E8Scg0EQdB7qwZeLxfOYjI3D24JT3kp11wG/jBUBBWEyGo
f7xdpE8NwqMRKt5JfdIEw3J6jmIOzYQfHRxVBORBF16ZYteBYTRIvxpCdd/j
HknW3Ne6DI7sp+XpkQhSFBDsYCZgeuxgBCWYKwFrrPHKu7CxD15gccFkRpFX
ZVAr5YpDkeFP7VIysEuOKsOZ+4fXJbTT+QlRco9Vg5zy7v2/if8HC/DtyjpQ
3d05CX2GqrvS67BTWn1fUb9hVth7m1SQdYmkeuM2P1xYZQmL3x3dbPHZSBoL
m+PSkQ7zxIMlnB3KhxjJFo+q/xQFMsSRuJxAkOoGXDpvmprDTYM4tI52aIwb
dNf0QcqSVIUTaymzNIuvItMovllNJ2og0eByPNVVybet4ZnVjIuCdNWfC9EW
voP4BL5Dh8mc4mAj0qUIxzt6W3+KfAOPKGT2vW1aGeu78LEYmiHcG8w/pQGI
xAvlseBQJwPKly2byPPbuxCsZgRBVnkDnx1zG1vZ3jw59bH5n9FdSqiPLhs6
fohKa63OTfWHoDIaHJWTDxlu0sDuAZK8jzIAxzffDlMXp2Tc95OAX4aVohAn
ax+1P2ZojtRDOxaY37Le2f9iVjMywpMQTEVYBY2gQhbNoTk5Z7H0Ofn+YE5+
T7LSQsnGaPpzgVSf8wjj6hiTCmsRoQ5QLkd0nhBaaf8oxFMlxK5anAXZVfaw
rrDGxJi9/0Uz7aeHtQ5geDQiOf3QWQre8I2zOtJ5rfRpcuuvpCVh9zgRa0rW
gV0elLVfwWJzBmTgdiLnYl7O2qp1dqE/38ZVw2t2kFXqz6cXMAJZjwyG2FWT
mAlW0nXLKpi/iydlMKa2hZoq2bawQH9+aDG4YtN/2dzanUM2iSyrKurWL6xc
4PuGy1KSD+BYLC8Cp6bUFY844KdefFQcRQxn70IhYtTQm8dZYera6SgQSg+f
m/RYpPSZffeLwQP0cqib7lt5pUmJ33D7acQs1hPjIrMUosJ39DQl0OEWC1Zr
eF2czO4SnUBdjnmxgshfzshcqoYGMLkvV//S/QcsRe05dDedIcWhY7d7KIRn
S0gOdSL1BtuPR/ez1y6zJVALMGVF9yZxf+rWyzzC5KZ1ZcoX9LefhDFutACW
7ZUFP8V/Qd7IHPfZcrC1XN72LIu9oa9jzzVoXy2nQfXqc0fVue6z39H1kRnm
vWQT2eEX/f1ffM5VnMdR3iZh2IGrI3hC24lxNQk3bTlTTvIs+jTE4uKX479F
k3Xm2camzTbI40VgDYJFa5fjgJSyMwRpk65RJvrt8LZPZZLuqSRGuYVnxOGq
eHKMSxdyb2nQmo/l995RLHkRsl0+4EzdZ9l9ntLjRuLk8k+r9JxVuGDCvt7s
FC0DdEFVWJK37LwlK2vTIgUbH4k+Hf/MXl0coH7pT4jl7/rZDHRZmW8E0Nfh
e44+y7bIH50gzi5jx76CmxD8p5uviD4ryza9g7vPBve12OaznrkVERoEJ7KM
VY2qogVGpxSZRHVNPmjV0dGo8NIJF4VKPi6RsyqQac8VNh2cs5970lToJRbh
gKEzt5L8yNfGBM86/BY6Z+2CVa1fzrCIrHCAkZG9EPScjH4zcaLNFeJGMm1B
gV5f1aspWo1vy3e6qvHAwckDCqHb/9AWgioNiN5Cv3WHfv8EtUuMe6eQXlIt
YX4ksfmXcwBCnCttMbXYea20zJsaYYp+kfrf8k8nXcKk5DrCxOVe8XWlC9gQ
ugoyAjDC0HKUVfN5BxtL6PSpUx5JIHEJ4VfOUAQerG6cyyyi24coSD2clw7Z
E2MhrxIHxgC5knDLiy07cHuQSUnqpAGNKrz9DQpT0zTyUlQ79u+LrfPPNw0l
vSa+m9nC+QUH11fwV12rV7zxNQvgsCvTlo+XNlCUdUJ9S7WyF9kNK6KSEWBu
fzGQJ5SYf8qVCNlxNodWCLpk08fO7uLjAxbc6iPKku+F7787TdCaPa74zftJ
QsXkte1ZgI35h8bc3GM3teXEkLBJH4/bXMG0hKupFK1IXBv0f6GwmYjZzWjt
46gVL2ahSQifyF0Uur3C/57brlVLVEfX8Kx9NQjJrVKKLMwb2RXhpMsg1VJH
Nr2P2XjvpwAcMTv+AOpD7CQkGbEAsh0CiGere6WaQBlA0RHfw3NHW4pZ3V1o
VX2Oauuqch9DqsU2fnDm3eH/yyOZIbuy0szJOcfF13smZESA05R5mc+bCwwO
Vb6aSb8pLcxk2seg6U0AmB+UVYZ1lsujpD/77KViFqMaFsxYHJaueaRavK+x
Jb1CL+pmHyBaZj+9+cRj456EoMODxIyqnHGx4LsaB7cDu4CT1QBIkP8o6nk1
q4iX/FaXqrZkPNzrWZlltGQrCts7As0ptPtJVIm0oCP4G4cQcX/RqJ+4xKaW
yCfsC5W6NKB7nTF1J1Bb7XmIM3k1YVEimZYqZklgscUYOBLclggZmTgD5Qqw
J39zwB9Pyg71aFNPKya/Qg9lY39y27RbQosEwfic02hDMk7ArI5Y6XLcy1cu
97aw/ePohWM3tCNYXoN5WlTtDO9jFgrrgsdQJpEIolGBrt5mMjxP0Pp/Akhi
Hxr6UJb+/2FDAaAflzK6Z1ya2g5vH5xAMrsBtmrHrlYyIYW9A8RSnGblSGf6
Ha8jtV51HRU3Bfnc0KkjC0FXrVgTXyLahgQCzHd/arMXtnsoOIb0YM2iE+aj
I2+izbTEZJCSL7kKjoe9wMRILHiK0/lXUJdNssxTh+K2u17YWgIHVDGkEZco
h8hx6GjouuE/CZvLq2RFn0ioU4IzITvgClpO0f6ICgo6LNKn7AigV7zV/3+k
R5GD5u9fuf0qH1wbl9ft9PjWX0+cWNxDigiF30PPHkp7EXt9z7btcpTo6dMd
EjFE0/46wL0A5Vu6RyOkPu/HLutFiL6/WlEH0D3CDE5KltCQLk9QE4qX03LK
didusHj3ooCeMmGHnpUtgvzehbMc0GtLwNk8GexBRaPry9i2siKf9Dp3CBL5
x35YbXV5Glc0Oie93clOB0uWxinI6FAY6/5HG7uajTdnwSj1XA2/eh+V5dVG
vuXJ5Zs20a2dUgKS2ROkJmNrgXjI/WazFFuFHxXNAdVEopikxRUGNn2ZTnBI
ZM37WX+DrBbAL6p+CwiAI+/nUXd6snobmHwZi/aT0lCx3RFGoR+YOG5MDSJZ
xqtrflfPcC2KOnigjGihJO3rc3hEUOGjQj6wsZTqYj1qXd0c0t0is1PAyllm
NqJQktEaVKUimjUkz3tHi61QXJXGCvfwsTPdlROVxYFM5slt3Fkcn9h5wtcl
U356NilHbpzNKCJlzfOBwMxAZMv88cX157LuQ2zQv10aFJqSkhcH3L2chKgK
U/QNWLQAEzMQaiV9/Ui8E6ZDwHSmknBZaqIpPR+M/P6IbmyP4AF1BFtG/rQ9
eSBdQ14aATb+MsV3aPbfXZR0VRkO1X438VUgyVGdcmQjoxPTHz26zHNV9BQz
BnhKkY19w4ZzwG8baM4qP0j9KzFBUU7OwHu2HKSMeK8h2/jH/tkYX7KAMWYi
A7vAn2K+/FQGoijQIqL6nJLZa8L9qoBzeYSSDp51ChRWYA5QbQGiYdj2y+eb
+9d5vW8N3eEbdnr/g7CVyUOULP2YVyQFL9izHjiGNiCVHttNMDz0T95KHk6c
/bqnj4I1Q4BqlMaMdini1bzgX8c0iwp5oT0+tvbBLwspDXhAf5MLbEDxGPAR
wnPrPFDRa1hnXYZr86LZbbxzR4JPsxRzhnAe7IZH2OssZGmJyRzW9FJYYQoe
8SwTHL70xg1FFbDa4v61DEz5yjddXMNOR+HHJNdQo9YebScZN3UjRxAMKWey
+ceur/C/JReoHcyqjAiVBGf1k7C51J6XgBGbEbIWGwe+iM7QNzWjGKsCk2xx
s4yiziI0L5L0yBijf2OGE+8RWQK1RPHhALDHNbvWDHkuZseiaPnVHJsJKdfm
/MSFDLh3A8wSibKtsUQdc37IlNa7j722QJ+jPKze5W7bE6DtqplVKr9jfbbH
q1PMmM7DmoX6jLA/B2niDeUa9Fp1ggeVx++Re+zrhJRaE40gYNDEHVKOrK8b
HzJK/HlSBENMQy8S/5zmxUf9I3OI64b4GHFkS1AGNJJc1cPjdYKPPvfioBV6
pczrSl1m97ciX4RsGhu8gf36sE9ZCo2XAcvBDHE0T47rTx7c0exRN8hUmTty
PJeOXHSM3iKCY+ClUo5IIkF9qd4Z7CxnHLbPqLTqp9Cz/AJZKAJINFsqtEvf
TguuUbzc5XnorX//VMl1LnYJn20Xg9TmhpEYhhltO+BrLAmZ5f+9uzurNyxH
IJJ8OKaKCnaDN+/qKLinUKC50rPvm6wPWmK3G0usXXu5vjKLoosACaIZMd0I
SVOoyWXCWe5gGpoe92VsE2Em1ZB6end80xucnO/V4M18DxjlL6RqUh82JmBf
NhFyHpaHZZSbecmks0kuXl70aKknEuSltmpskttfg9ewZ6gi68ha/HXCz2NA
8EAYL15hs/+nY0TyEZjyHgLl4hHKVBetDmFP+eTCco6v/bJyVOVo3Yde8xxO
a3adLl/Z6Phf2yB63BnPd4oZ1fEJV3WghuWnHHaS5hs2zzBxOFHfEJeJEtgS
96+CFJpY0hEwO7hU+2WBOjAHopmmkLsDnWw0kInLP5Vi3pe8KiLnGJI7RMh6
zLFke9l9jO72LTx1sljUpZdsdX3Q+FvkAJag/Nr18RROQAmtYtoOztwyPlkJ
hLOQ2IdFNVHQ6xRubRNs93vVggxbNZt4YJJIpHyjNFGVxCWbawqUKnleajwe
JXy6iCpEXXfPZrl//f5aQRECNK2e+5ewE1uoVR+9hCc1RK3e1LIibo8WWj/5
fp/elr+wKihcTK0iRHTXBIAWnr6tdi/2GMzWnc2GbRS1SEhcvauMrB6VBE9p
02rKPycGqFvvBYxbRaDZYVQ6eN8r+l3GGyuoOxkjIVtTjGz9jxn+VU0weDz1
dcKxRqDh85UHre9644QB3bICED8XmZczPidfhpMS4JIqW/JQ5Xe/+YEoHFQf
Q+zWl3163U0GgmylRKFzvMBMMl43qeUEMEoneThnVI7zIyaIl1r4EGvOo9AD
/Bt62uS2N2cFIdvBZOkgbVOg+B1ObACsmCd4CUBVX8BdtA0eQyNFyoqCxSXd
4oegdM04JYsU+BK80+oN2p8b6DK37MX/8qyM7XrKVNS/7Y58PN9kWsuZYCXr
x2wbGrbcrR3OgExom8Sz5i6Wa1yUGFuucyAxCs/b8bTcxO4XkNjIpoukvuaq
v5PQSH9YXnysixFiOC3fg8uxuSbuSkVpi/wb1ZpUPOMJ8QQtJnncaVEI7ARj
6wBoqDRiU7aXYfx2v2hQ4h4TBvHQH170B/5KtKuzcI656RksgNTvsamuY0LD
4w9Dw7Gz0K1Gtpj6UKzaePKwYNYsWNbKWQMTpH+qjCcRtf+gJaRyhyM2wJIc
fJqSvRedxWnCpClsQG8avKXPZRwQgrf2eT5EA4qxnvbDlzQNnK1EVVogFqqD
bDWVfHBDLa+gGnkkjgVUAMYvW5fuDhnF61VPidBXT9J1WXxm3ef5JtYcLqj+
3IcqKGYNsDsObng00+ZAJd9KkILIJrtrkaTYu4z5/qKnEq1F0c1lWl00a6UA
RPK1sQOIs7KmvHjOQMSjD6f6StFzcrMx4vDacjpdPWEFpfPYBDBtu6a427YJ
jO/klQTcXf5rxLixYECG1d9+LGHbq5TBEqRwuttVNdO2VGpQ001Tb9R59xsK
z6S0i0NkeH3H7uNyiEbMSsGMtVYt89jrfLl5r8Tht8GW8iU3y1ooWgCFEEw5
Q71QbMd8I+egtoaHZzEnzT5RRh1whSEVhMW6m+xiQa+fSLo2FwmraQF9Knzb
u1tDb985Ap0P04V4F+2gWqtHUJufJk6ZV95Ff5Zg1sivDG4+7uiVfBtPsJ6c
gDd9Yr+Smk4r3Je9ZbyHAmRl8e5SMxtBtwoLrOFpcBdwKBLxKEdcqe6pG6kE
Uud1pvv2jJoeePge8ir//CepYfwzUbEBqEpfhIJv56Q2i+KCzTOU76qWLZHm
87kjaVWwwhEVtvn+uo9EbPedVTmANTmuM10y05pauz+aiY3W+H9lVMxBo9Da
pO3HXpeMaqD3w6BDDvaqUXbZyYYAMh9yQG3TdMJ5GCwieF2pEB4B2P3PYEbs
fvNfbEobgfEEZ4FOEKzlS8IPvdr0bumFX6UDAU7U479dwy/tLD3TxEtN92NL
v8mCRWnZ5Yf7rB/U4u6CF9o+C2nxa49/u/kUb2j2MyohCWntoQm2zlDMLbFM
v1Dr6aSHKaDQA434AsoWavpYT9Y2jTdAlb88f1a4PPGCA+t4OGOIAxpK2D6J
d32VlLrVIRN3+J3j2xGIpCXe4CA630nGIRnV9VW+NF8g3RrHPxFs5s05Im1p
495MdyTA5J54OYqqDTPpRF3tx8A+pB+VW4xhQpNVKbFEIuOIkqoFbwdnS5zv
qJWNAaEXsgHj/Fk2eslwJb8fWmYpZo2sZLeP5gwOkIQ2znygXOlGf3pVwGlC
25zGOjIGO6BIzHbRHLVw76seh3IXaGGufitFOd7PjtIJT4iGW25G7oqhipwZ
Jrfox8vs+pysUZ/mAiVqEskRzsBon5JP8gTYRRX3dKvYHwRk42nx/lffNHMg
jijuWJO2goXXZYz+Q2l4q7VUuhT/Md1O32/HSWKGamzpV7pgsSGTzYLKVPNp
aTNHSh9pN+paI1ISw7L0Tw5smDQTlTCoHWJIWk2x1lETQ8OBIML/TgzgKJbH
fD5FjtnYOAhiH4sr8Jn/74S4f0qqKxAcjlGsI8GH6JAYfk5NTjZDdHC+cl0V
NbP7Fgx4j0QRSxZu8vdzrC3hYCm1d1Ic16t1kQXzVjYBCuuMXJ9+EcENGM6P
rf1yCNz2M77YBH06oE6yTemy8SkRNzCPeaKhwh6Q1AeocJrIG6JA7Y/l5GVH
OdCsBi7KKiqRLhAzIH/TSLo0iPqi3NO4vaVG9DsQTqnvtnwH6LZ+G6QKsg4x
QxSG8Ocn1fBImuOOvxo8gczy/h7zjHuj8IR0fDn5byuSBajHh8YtUTuN81iY
x/NQ4FipiLlKtzfaVRvMOu6Km2e6IQfjIZcUoNCDpKSHfPbbZUcWxkHqnnnv
nuNB/1OecGbW1daEGiyTbaB3I24lvbXHYks81eObNqWCDNqHdIRHZC3zV4Rw
KjFtUHK1yj/zeMOU+CGZMFD5tPgdL5Q8XvY4GWbLj8r5X5I5p5D+R4ANEkaa
0g/9V/+ZwXDldIY05dEhTahlqRg6ydAwbaucb6l6cl/uWOahRyAlystQlIU+
Mj3Ig7bAHV+FhoFSaIwre25zhq44YZ5aL4K+m7GqVXmOI/E23yVPaSLFYeRI
1R8xIRmZT+Pcs08c8CEzWsfZy+dJvv1V5Sma/eoxGOIyJYQxGDZe9jBS2Y2c
bVA26Qi6k0mSApsqZea5UvpKshkndQ3tCNlD5SBGfAtvogHDumR8vwDgn7Qe
g0Sc9u0gI9y9fCQ1Jpe26zZahaJFZZwwM9UDBCTYIlF0CBxo7WP7PEyA0MWJ
UzFrXMGhlMs+xy8kIq5bOwbrhb4Q6G+QsCxHxx8yXrxqH7TNpJXn4+du4+RP
ICTDjoFvSojHyWSPsgsz+m7GXxopLGSMTHMX6OpnoQNoKWoN2qQPVrEu1/xi
db7LFtq+Osbg/Gvsn9/398rzbIBkgJoPUlah7sj2Dz1HhrraJkqsIWNddKl0
SNh+ULVOYStEC2vWeckD+TdL82GuH+QEAMsp51oAt786Ck6MNB+NkTa//YxO
d4pz8HcjLGudEhalT+D8dgZclISW7L1UeRvQlxlLQS0ZxDFweZ9e3zAy5FEF
0cq3PygHr79YiMZsNboXfoO2nUkrp2i7B5k2/9R1fzCrsJsJlU99BTNFgIxu
pWP9qUxSt4ZfV5W0+vzFemgdIgXHwFLghbE5ODXEBASmNq5cqdiqgKGHKDC7
JnT0NZP2mEAzAsk4LXbJxs1GXXjT0rWmAsPHg9LIX4RoKstRxOXbd4dq283a
KHBP64m8tBunWX9zx5q+JLyhakyR9CviRpvr9BwCjMnCUQFMgzL3KisficIp
23Z2Bbxt489DzMYJxRzdYqbYW1AOacVcmkvisESKPpQYwS+D+DYBSwLxoCkP
auXhfZDVPFzYm2LSFTBn6raIH5cvTiOyXUm29Se//QubN+NgZqdyc+9O30jH
Ah2eshBhqa5XQrt+Jwp/g7I18thHHbHPBg91264dvSYTtTRE6pNrLrzWNmJB
DvYqFz01s/02bRHCczBJ7Pa+FvAq5Z8yHIshNfhO0z+84uFm2ynA4Uq9yqp/
snD55bsPZe4XYSy0Dbx05NRSFBWD8atnQZWvxqzluE/mr7CDUhHDMGc9M7IG
G1OrwmL731kY2cRMcN+6GTxx7ZWR7o830Iu9e/1caDPEgdYTzJ78MKARZ503
gKHNeGXU3w6s+kkwMMKD85Uj3NM4Inle7Hl3GEmAxovgNd92vTNqjpLEMnE1
D5YE6G25qPGbA0KYKl01d9Cyb/vOFrbIvMrLwzmnRzRhN6KOp0lamseu22i7
pQ7qQ+u7w5xgsTddtD8Ni/Yh2CeylwYtVjsX0OCMyytZtX+KtwKPKZ2xWFtj
9JMReVyLQvzu1Fg+Z/a14TtLlybPwrlySrm3RoEK7bujyjS9n/IZrvwv2ozu
mO48r7DF78CK3Cnqo6kbx1Ty60CHNhJGL8tlwR1bgCG+r29ITzdVFqnAxvNn
hr3INC37sqXicMIb/RwQ+b/VpQ/tqDBzu8uJcWPWx7Cg9xwpGUDH+6uLv/jH
Fao676JASgk2ysymeKmz2ySqf1EL6KnRtg1JfbtVlO7ndtMnmH1Wyy6VJR0L
wc0KH5rRiYOv+Sp5DrrTxwCIs7gNyeJLKEGFtQjIDVdHBFat8v26bUdEnnwO
UojYHeSWD88k3W1kRlb1CBSCPiEKppXxeDc467nK82OLLlDN/5FtAOgQqD3J
ZQssaBwncj08zhmykVBII4HP+fVwlH3Gw0sb93jGrMekkrDP2MVguGo28hB7
TRMrewbugA0/CHoicBzpPNk/NDC7kQV9IC4S4iafoyxn5yebD/hhtKbtemo4
qT7Dy/kqV9Qeq8kDSR+f88nOhhQckz4MGuqMvDvYxhf4Z8Dyj0QtIgvv8IsP
zWRm+DIPHvUUU0bYWJJvioF7rnJiKsKsjToVY3ky6s2d07z2nKkW/wmQDvBl
9eUI95CRYRgLO86cZosYlh9nLR7Qx9jgU4MAGyhEUzmSGTVP8rZ1Y3AUuEVA
D843AKMD1pC/SRcDtd/4c0OEwYYl2qu1k2lsm+LbmpbxNqMduNb33A3gN332
u7pewNLiPxK1rhx5nq86mhHlK5/+3LfIbW9Um07nVIoU8d6Kq9sd1VugYici
kyTgBzxfqoZ1vRAEEatOFnJk5sAKxR0La8xu7mkEEJnerkZ4Mxw9li5wKmzC
RadogZH3vlXSFc8CEfnh0ob+9oeiN6n9f+Mt4/ovNKoZZxnYwMQeCptyjRfn
VPWKTNs4PiRQ+t8PpgZ2kVeU4LndlkrAoUDKqgJw+ZBk226mR42oqypUCzDv
QxZ7vJdMIRg4FifXpQtVkeJo6hEPLvQSd4PYttYyDYikYzMENlGIBNeOYk3e
zacoPTkDdsq0iBR/Wm8DqpOmhsn/4FPQJUMShTfoSCd2CtweVboOA62MsYTq
UjUDOT8lyvw0qSbrdnDdtMjP61DrnvzbHLeVVRMYDNKkTaEpRNt0A7a8CVbT
EG1gDVQuD5CgDTJzYdzxnpNRvtW/wJoa/3wp8lwQgmF0WCpX/EXsINasb8Hz
FYoSUVsx8K6kJx4ohE736YNrfr3bA4CNaoGdPVfWjE+9Qn93qz4osukhERgK
6CPtdhVqRlc5tBz0F3Btmcw5whuAAWRnRdTyXydMb1ZKTi+ce2VGT9aCOkOs
ZGdv3nX1vQ2CT9+TbXOWF4QROZZzCq04/nDfU6TY2/kEu6bjQLs8NcD0m1vw
WVHpfRi6iRXoa/3sxH95QKdJQ34Zka481k0I/kaeM5G9X4bWsoQhhrlXh3xq
uJ05FlI65Sqi3jluozOFMeKjJcNkvd0HtSFtmLWGLDh5GEik7TkQ/yfymLyo
JaZIthC/j5faadyBay/Stj4Nf8hMDLOwuQCSdd3m9/kfJJ2qKx7u6uJNSEWz
dnUz+v1Mj9wVgW4aff/UTuFK34gDO51S9gNglMcGpk5hT6e5X2GfHLhr3jsY
fruTJRSmSXOVZusVq16vZ25Nm5QHDJtqUs7UEr2R13xI64oS6l7/07OC3MGS
bOYaOmEbVgun0xoEpCtIwbkxN/E6YyTG6lm9w1OyAW0EelcloHWTLrzgWcr2
i6umCHhGUL9dGrUdW/J7Z8X6nhJedvP1su7ncdAuuGCGr2oXe9XhEynRHDfN
LXW8OwVxvKtuXiP10F3zOLgATqriSWHEOYwFw6ScOIaSSGGO2V/r6sU6sFe7
RZDN7/P6/RbCedNTnE4foL7fvSAM7pxW2MDK8WWwcSWB2JuZPgR8RZD/pNJE
ghk90XhBLG31tKWJp+gTNmzbsvDF2zWAF3xKTdZA/7Z6WQkBh8+sLani+Iwg
HcVi8Xb0E/LpN0qo3HNdqKKGfveMfvd4KtpDpVjVSHj6sNh8Uo0jcIS3bTcj
Jt7ez5J2Sefyjt38OsIPLefMMsxFa48Q6crNKTH533csey2aCL8M+uHH0AhP
+9rBEZRq8MiVuP3hJrs8Z8io8XZDJAI3w71F4QscxACPQUoc0787N4m265P9
fXe2oZfT1vjWce9iBB77HVVpFd26YY8JCoDaRlpdQXnNoFphPtwLC/QcayR1
1ORMELmMS891QTCvU7bv/jYoZdtw0Zq1/8HTsusELVgjO90N/+H6iOvSHaaO
g0NuJsrqYUNXq3tx6Qe/gzTSEHp0MuN/Kv3AMjGaSC43l1rsHQixCajjrYML
BXvrKCo7fOmpu6y4C6teVqGoxmPWzmUBfVRDtARWqrepi5TswYMmTw1xrieR
NX15/+HgApJySIJ01FLtgMnNThLeO15AXuT2YdLU3sJi5UmuB/Kry09MTMop
4aDcZNXny3SEC6QKd0h9wEvA8I7jBEeQdSvvDsaMAO0j2+NzMrpqVRo967Te
qgmxma0pMqFMiRvEy0IZE16k4B/Y0AJFpQ7lWlPCPtBNyGm4ejYLY5Hi7cNT
c2FhhFZdKxtahn1EjWeRB2CvCRHUmWOH/Wxz0uEKkBPxyerL38fEItblOYQ8
MKCyEU/paKp1FrvRx5UDr5iX+LNqDnV76SCGB9qaZZh23xUmnCRkBM/W9wFl
Y3aFZ8VXN9Q+OviI+s6z5UyhYZ9vSIMqAwOvY13mXbkM8dbEruGa9NK3QGEy
nTRDWo+Xa7EoTNN/VMpvmeQS0xOXAgzZ2adNQ5vrJbayOJx2QPVy+MBK+Wk5
gnjyvJrtVqAG5X1qaVzzlWrJ9Kf++uFRZYKxIhLX+YXn8eZeZu6gOoeYNUd6
vPqivPrbC+vTkTM/SqpkhwCtCE8EaIPA39C7F+8Dw/wPx8RvVOl/Sahyf74L
SDWh9L0mWVk1iR1VEVrTR2OVa5ln73StpqMG6GNBmNHwYHiUi49vY4jTXyzT
xm5UY6g8ETQUrAzWAE584zhHtKeoCaPnczS7pf+5JgZvqDIMltNGk8PR+wT5
+nT/S6xcSK9CWkdd0aliNeqIgCb8L9UOaVrv87dOl9q1vfpYCnlhITMKiU5J
zO1RIq4JzjC1qREaOz4NzvntohuLEkBscxm0WzuwfcPf3Klj/CyTXzRJxP5p
uDHxqh2UWbN7L98Jvw2G1QS5VjnlOrZNr3D8nz6tbj6+NOUZ3ZCawcImM9wY
6MAAwsyhG22GpdYB3lNu5urmT8Qe34VBgA4NtWLbM3R8uIuIjcB23AvmFtIW
h6NmDifZD6SjGqB83jchX3Hgzteczy/DySALZjSRYHtG4y/uhSbFTX/osDP7
MHy8//mGffCvXyfzRggEZvt1yZZ7RtdnwXzanIdhpkLZNVwvbGm9UktKPz3F
oC6v24ejvTe/6itHdDl1mdzMVlB7xVNYrOnI7gmmfQcIuoDDHXxOH+ignlnT
MBRnJ2jlimDmqpwj1w02LkzjPnYgMrwpdz6inINWPoCutqAbE6TX26F+ZOvU
xF2q2ldHkn3wxaa5l4xKQIa1ajmSWIifECLIpye821GmJAIkLG93E6+qNeQG
i8nRpq/2i1USPTW3ABU+z1UYi1d4tLGoW0e6uGyd2VaEzOCV9XH7K5HbqREO
oRxv7uLOgUX7+c3liSqCPMPPpQXOub/R8D5I0h9x1ggf0OgWXoOcz9QabV0A
379Gh/d7mHvt9qqnsyDca6UegGgfuxWCzkCv1FIiV2Yirc7Psnpx76C+3wTn
uAT6pPA+rbcB8TrVKFJLKdusZLloySfPSKS3ScHosOCkcNh1hQ634V8Zop6D
Dx4FLj9DklS+UFRBn3iWIWU69dBsJ5DlHRtajvf88tfJjBgwTBDMGb0Uzkpw
rSvK+M8gpZviqQEGH/gaHk9wLDu8fIzPzoBFuF/8CXRREqX9GhI0miFPZvXs
MwZl0KH242shtrZOXo4MOZWyWxQ7HR8peqlcoeMoUlhgLBOswbMuTRDDK9Bh
vsibOUa1AbIy6MQqBeJJnRyjRZ2NEie0VcDnllhn3+UhdOxWjR8DlKPCuZ5C
TAdtc+wv+1PNAB5jxcsVXHwy03kCIaoTuj9sd4pENrbL/iRiN3rtU3jTN5oe
yvvEwFYY+vinZhMDoRdFjCN9CghfYnF6A7NSMR/GXjmxVlMf18e6WugPXYdA
9iwBUUUqVh/mTReFg5ZqMVq7vw+WPDWFVCXptKQgkU4Xhs/5pSkLXCg1rPDM
7G90R3NpeM2S1pZWzizuwVCLLLo4fFYMzV7hjO+Ry+YwmDPVjkU0782bOmY5
SL+CB2+orwJ4Om5kevrDojILox4w7/I+Lh2pyBFl05zwhWjbqjAdQCtaJ2zB
Ipj+8r94Zn7BSzXv81CmWPOyIE+pAI4v7aeTYGYOIc+XWP2/1N6KWZYf3ItV
0hKbo74nTDQFUv28bCt2PVglIMXpNshYM63EoQmBxjCWUxlkmPc0Xunx7Nu8
F+IZNXCZDWl2H9PCDRoa5wlNp+0/g3cSU4vi+usKDu8g9DAv9a9nbNEi9ekI
pEveuS/3MqbVc7osQ7Ai918fyqXvGxHJku+3wW18f+Yx8/KyQ4pgOuDbBMuK
hh/ZPULWLVyotBHeyxd4wmNZN41m8leLszpFLChP8w51WTSPvQdKNMKr/uSs
tLnGJoCvwXA3FOrtgXy2bphlY2oATO+aoenYwJoiz4SBPhwpBf+lC3b583WH
+JUeyrohVIEif0c6wkRF/HoK+cGhUVBdWpKCWtpXB35PnJRioA6VBA4O6qPx
v8GpM/+mnPFRNc4D1s4VoelyEBho1cITdrGJtJyEp0+friMKyeKRGKx2SkN+
Y/MsctG0eSlNmkr6sst8WfzghxO91GiIqzuS8r2IApXqIOgyiu+Wb8fnAMi3
YjEyeOTi9+75eEhmfoRdJ462tN5miiiUE0hEGP1C8mQmtBqC8wuUNmJL91sz
j1gVYSmyND+TAuBmVOD+5l8jJmNsJz7+iuSYGL5nK8kh4SyqkGDpAMvzZfPm
E62Pf51woScGGXTdsGu/n7ZSA0IYRpu0cI4QUT6k6PA7jwi+wjZOdpCqkFGm
EpRsbKcPJ8wR79dlk8KVgh0g2w2b3Xc9c3MSguCzdSQUpC26+fLgMGgmttFq
8tJXKoDVULcl76jlKowofq+YCrTgHuO1t8j0+jE2Jus9oboaJPfYh27oH5fb
k6DpTsJ/1r5LPVC6G+nby5lZlYCbjgg0PQ736LwxYzuXfIYG9n6jLz3PST94
6ZGzK9H/Z9KT7XBnAoujlh1Z0Ye4JxgX10Dsx/Jhco/XcwjSe/mNgpK6cria
2/pBZmjCTKi/rGLJGYTlOxZQPr+nd9o881COaG61KFk7pMe/bro4aVZbbFGz
5lCURiAlSQ3+/F0SExaA/kid7U/R+0i9L4X8Th1e9WGBk11N7D+fvsYjSemY
zoIaKWhAGg2Y2RJOSUPez5+OpiGXLkkOpSKVi0peIxkPCQqMn4s13Y1PEOTq
0KXRZpOQaid2T0t64CsOae9qII0UpVXfcVaqVTjMa5BxBHM4KQFj+3VVqGKz
hdIynKBgYeq0ENKAqhN31i4Uz3fMFybrqkI/owz3xADhWV/8HoIubdkyz8DY
Il7UkfNvSp7b2TKiggOu3t8vq7UbsL/l7kpL1531L94F+/6Tot6Clmh3w1yE
9vZdU+3kuQr/QqMhubGVR2i4MPcHt/DxbYea/yyWGVBWp0IE1tSRmRwBbIsi
iqiJK09OP+6ZS5Ia5z9UK75F1c9b3Lt0YhYZt7k+dO/2gymsJs5drLhfxO3v
ItY8fmP3NILv0HmRM/0sVAVoUoQ1ZI9wWe6N4B4BQHkTeQXiWjZ32PNiJqiH
y2kqoCAliUUsnv4+kL+cgDKGmWLfo1j4qUxUb2eY8cdx7o02CV8geY1f5vLN
ZHJovOlwUfWRAvj0If7/ap/GEKPR0BVN5mZjZzZbLZK/gOR13+pGFzdHKTar
CDTwdu3pjGTrn9qzHhUZ9ahiV+ICDtsWrTls2LQs3HyAAIfYwk3z/qWFzu36
GcnrGOuXcioTwKJv6LIIpVKHTFl5zB1MI5jWuV+WfyAaE9P7CVEqSSacxKmu
JGdm71Nq++SeZHqrW9IOkTaQ8Uf5wQ5GHWrz/ddmrefFMimFaS4lIk/2U9+C
3ZRas83lOm9V28hvsBct+tL/m19gGIIQIORu9UZWHQvcX9GBKZ5RgUgOgaPI
FrzmhlyzyCOyfVlC3na0p5fjksrRZTNdfU37jGVyxu3m0p9cdADfCyc+AIYu
UA/SN73xlXYSu8HwuQ4Pdwid/LcqPMA3g4gnnE+RffLXW1c+c3nBNNr06PKd
sPgH5l7XyM7CrxaYGyfWNi6Ry7HRvxHWmyrvooZBGbbpB8ddKiD6BZ5N04Fd
13wjJPEjIylsqBvANuZytlCcSKan7iS3F4A68/sFyOOu9zB78+TWW/8PN5gE
6k7LM4voRZf7xIRKF3ZlBsCZ1wzIAOAsM6Cio7g1l4V+LXiMW3RIMelIGevr
1M+lmzpOnkxa8yJKGBFbOChzw2RABLUK772NKVwKT0v/Q8CUuWhHoJsnOmWT
cw/xWtJFkhpQek4HHLZDUwtrdnITtLCIyKf00aOATRXlPvH5lTmTGnobxk6S
o/nS351sDot1z34yiHiOE6J8VJExsxMj58bfetgR1SDX+igL2q5Q0Dfa4R02
W8VIjW1LThK9dQs40fw/1UgJcWddILSrxMz/OGc78D63Q66s6RXwr8CYRde3
lkF8r5TQyoVh662VjiGJhuqHNPIg1RV3X+U1+nufjGpRIC51a2WJ0I4yGygi
7KUbWuIdmFEM7meEyF8qj74j1iVlCPSXu1qc+WSMAqT3YlR/ikWgWeXn6jBA
no2Cwpr2aVZ1Y5iZK4T4d6LLIOls0cdOAGIJ6opNx3Nk3XpTkj+ksu/bq1bj
Zv5JtG63F/D4Uehh2ZhR7heiYYSV9Q/s8tRCqBkz77bxFGMBa2wjCLWCR1Z0
AkwMzj16X+xGQGaqqtibKQ8zVKr6NilLFP8MSyhQGKGa7bOfr0XCeEUAuN0K
i/VO2vi3RGvPKr5D9x5LCvNLD83Z6AZm7PXBfFJN1/Ekug/b6F195biaC/Ly
gbyxZzuFgZYUkK8Saa9Q+U5WftH04BdSZ3MOqOmGEHBE0ktiD5LcTjiB92+t
yk7EEPalzAhOL/VKjB7FUhVtJGiZ9ibLFHiZBGSArgJT/Rcw7TE+azcJ71EZ
got+C11rQvojZl9NVaBuQy1Hv7noxyXsJFKwcNkBHIUdoFik5KnbUpSFmuBh
+uvAbj6ezPAsHEJERPFW/+Z0R1s5kmzijKSn3ci0HoKeB5vD3NPr6b3DnS9s
UfnqrwWla1JIssOzxjc1nGDJuLw7gXntqst9vi6RR4khQb7IFnWVT7HIff/X
RzTLbyleDo6comsriICqIpEn13VQAVzyIRezNytFDJz+406uwX6Olj7RmkEv
hYbzZ6MlWOEzcgsL9XwZ0P2CdOTul5ipxGOckoWQBd2j4JPKcQZ47DuoBFvs
05eM0bTFjUVwFnxyNcxo+xPWkwBB5KKnrQpL1XpGiARbZGd+lZdK13o7dYRY
Fuhbi5SnQZVvL7blfNnwEQcdQQzMKWb6VRTV+vD/Ia92F/ukr3MBmkX1Zqf2
DOk2pw0xVqELV9v36kizOJ8gh2N058EPxs+dRQa9NU16M8KB0/vpEpb0512f
puULItkI9e4nJpDWjo0pypLr6EWgdVQ82CxPBUP927CWfWQjtGEyBEkav9Q0
OoGX8kEzwThrfXyxxlszPb1gNW3kSipCshfZYBGf3nbOlg6WhpbqWAo7Mhrn
nTfuZaOU/gbXS32new+XTKf0xXMZlSV1yqqF0KnKhKlnUyOsXuJB9H1+28a3
iNEv6LSQ9y1N6RzfJ5y2GacrdjHJQTSHUo+L/g9qXVr5SPbAmgqLTGiNi+EK
21QBBvsW/cLou396Fp+w2s641mjCQt0qMhMT1uYxLvEKtKL9xRBoxKbL8pm/
vuOmilzi/+AqICc6GmImUOod/Urcz5w8NsxzJDmZvHtaCSOg6bhtg62HvYU3
JRqVoZl0n8Z/s1XI/1zcPFpWBmfJ4drOhuKA96Lk+iXdV3DS0f3wZRPVtNiD
dgTBam+ToKxnsEZrfPR85Ku3Znujlyd/Yzq0SAvW1WdTRfvtypCanrEB7ihK
RIaHdH2sL0SrANBy4unrbJ7ob8MVioAB6aPwmv8gDzrXU6jPXz4wHGriUG9J
oSEhuqqPtkdgP6jlbB0Qs8r76TmU67KfvaiZjayPkr+DDemCb6/l8G3NLLyB
wcAg7CwGIBFkgG4VkNKF4KDNNasRl6AfXD9/7Y8Hv3KS3CyzrQyJKZDZ7UnZ
85PwFUCCt1UDRu+4tSFefdLcEceyV4+8iWVvAaW+SAvjdnBTZUshVq7o/kGZ
1oVUXpWTZcndronMIpRyJQ0q2kCAlkRVWubKROGg/Z637c9oszM0ZnVNqXAW
ylZi8Le7yc2OSIRWP4xlJ10XaaQmFImMw1DVOgQxtIzaaIJltg2Ptiy9xrg0
pFcG5BXeMzZKALsNoiqrheX2seU1ohxwSAip5yJEC+ioEA1qtgNo0zi4PNxm
GsllABgysSkGv6ZAaW7NQ1TeYpxZGdlc1+41w5GMF86i80waOD6susb/Slpp
JPS3pUYOpU0vqdyXZWYCtVgCmU8NdeGzam3jUZV0w/TaFLUaFH6w0Em3gfu8
/xSDWjEtKVHi8LL6an3eybbWmaQNGe3PPjgi1NG+yRhJ1CxqEXWJ1cGtthGh
juMsVELkYZ4jsZp2y6Db658RxE2rscbyTDB8U9gvmpIhfEFWcF07CQVuH9fR
XRYA2SQFtYlPvHLgeKhisk+6M27oFgIjY2v06zT0WnJ6/I9L/En6XV69IJK+
7HjVSP8YwnKn0b9s7HDKj7VOzCpKdixpA/PAZYiYvi5mkXZTvPvO9UV1UN1H
im6d6FnZ59u/XTHIug8vDn+iM++cBHiZq3gl7je5e6KAvMmtmJ8BptiEiuS2
/QbUcI1L330efBfl4yytQ5wUss2qb+WyNlUf2+Cpwcy6K6rgzjJ3HAAgxQsn
uaUIkhhEMU6A0IwBKU9DHEhqO7Wgu5IYpe3FGx3MUnMajsG2SbXaDRjEXH39
ov3wBMeHw5xeAYNYB6DHR1cNclW6bVDwESHye854N7p2z3Vd69iXRfWaed0I
2N/uvKDSlXpwk5hIr2fdHj+ucMLsDbbcSSAeE62esQ9CgjYOCoTqgWS4NCmV
6h+PFWsax1sHYwzppxRMUDbbVBFfTbTr7zuqoKQMcRADc0o5HLNogzgRZJ8K
o7O9acNecrb2YB2dgmkBo+Ku5x2+9PP89DFhTd4w20BZaIdzaQmeb1+V8d49
RDfyGWZC0Oo8s4Z7fzAGU2jcdcDQj2zM6NgBrm02SphE/fg31Gp89m6WpHiF
lzmtE0JWxHT0ZBuLS5JCvJ7WwX9/ndTxaIoAKvB1Qx4QY7v5yak6cdmmq142
HDa6vkjyfMNEewBzZ24gI0hqXnH2MKIorhPZ8SgCOxXg55Wh97pxQDCRErit
PL7zNmjqINMajH91IhT8OF4TtP8kMnTKB03SRyyCFUHOkiG7CNwqWN2IRp6d
ojwF26tzw9HeCZwG6xtQIr9Zk9m/qIc/rCvk0v2mtGjcOa3QYJ3WVxw5iXtr
2BBzcPVZGmPWIf4k28dccNyLGBLKi6J7uLprCJ0Rt7epIYTlzm9opGLue5Ux
lIQtRQ9DxDUv/5Ttc/dsVkxH28R2m4FNCZq2/Rfh9ZZ5ADieD0GtbGuhrMC0
S3w+S1L/2Mn+6T2VnG234TcMjmCfl9Cl27wJni1h2Y6k5LNCc1/9VrWx+306
RIBGtaapEKgsn/D+haxgKTO5v8GfqRIrlgO4kh5jo8JAk9ShgqCqwSIGMK8W
/Jy+7P2KHkbH9kURJXgJKWUOQ0rPwsJvVrb8+O8r3uCGuWAN64Dfr4qgYVLH
wBBt9lShcPvBswI9INilwC0t/AehP3Al5A1CxXs0cbaJkv+IBNW+RXvovJs+
FRYz3fbReH+XG5c619EjmbhKPxcI64n0Z2hs6OrEo0szZHDZNI7VPyppzYW+
FTI4H6MwKXqFQZMQpNJUSEkYAYn+9qA6JMH1tkpU2WhNWiB9LZfOSk7zx27q
4Kg1osSLABqwQoASIt1M3rtGlJ2OncLaalnLslWYsRo9MoAg/zkJqNyXexF4
63Kx/7Aw6wRLHsGb2xcTQMBGhs+Ihb1qPJa1YiWJE+i8hvhWpmYTIlxKoHeb
XayfQcPLr98oyBfZrA+TKLizNYQsJhW0rN08BudhxjlvY5puYXYWc8R2+Ul7
Y/hS0qOCy5QiB0LagfgkIkromyWeCegxkGI0fIesMnIc9ja04rvMx0C0xfFM
+2VG1HWGMd38apjigQkmfHfTUh46rGyKd4D6APmwEvpV7j1MTTxl+52d9oCl
SSxA0GBuQrQ7bGQpmWWu8elu8l7ygiSCfzmmw1dzW9bsRNFdDk50vA187RGt
Oyebespzn0ZARx2DJajTEg7/j439uc1zM5o7GZLiqBu47Mj0wQYM61OJbNW7
8B3JBq/47XqE4ShjEjG6eb6uF+mbgPkitFpyB7Hmh940ZgKBnaqC1cZyq22b
ZSjNqwMqSGZHQ1KoBaSHa/NgJJP0/BqTJWkDCcxdWftLtstpmicxmgVMJE4P
YhxA3hUPq/5dpHuR+LQqZUeXgbXslnAYGZ4gD/t19NfiaOLsAk8C8mywjO1w
UHXmRWbBI/2RtDLDKxf1vd98nb0xVj0WHrgWpPp64EN2fNP5vZgqyfYs02v2
GV5EGxtYPraQ2OcmE+WzBnJ1yR4ayfg6G2KZQMRPQKDbM/WNKEjq3LMCx6tH
/lZSIrF2ybouqNzxtuTYCxPq5TF7IcbFE2AXgBekEPZD2GCbjn9GLhLqClRT
ESC+LuPWkYvvTk2lpfYMACYbJTgwkHnBULwtJtFOeW0JjOggYjDhxj4iLTaF
yCyqyFlTZ2HZOua9zOHB5Nk41onb9j3OzMereCG41o/NcvUc86WIS4s8ZNdR
CXEakds1kE8LvRIUPJclPxd+GwZ0+llBhrlwKW4vp0055XufP7Ze3vUB+5Sj
J1pfVJPz3NJMy/MClwC4FjNExhgCi0vgFalCqYWQ3Py50drSkpR9c3RFAZgR
XNBnglkUsOTqhQNt+N04rCFbmp2QYYnaJeY8u1XKqbAlEsErO7I6PAdKj88+
v/D7l4ozl/XsyB51B1m23YJVDOKe61qlVegNMlp5kIT3bg47TMYZW/zCNaRU
sjagSTKr6y56fJmRLZFyiGF6Ds7NHBc7OnGEWUDb6cBFBmu6lkD5Qugn2O3E
l2x34cM0+y8BNVGJ9+pYZWPPZ59pZq7ZdQ8JhlVztg/2Sq1+EwGxXpWJFqyJ
8/FEWTivTQlpjVbShQtlSU5TailfX3z88E56See9hXkyTcBI5uoEHnDV/LPO
StouDX1akXxb166R/zLTjAPYnOpP4sFgLBeglUvYyQivEZQm+lvw4Jgs/LTb
L9u3paH1pyXWtWYdBszdu3ykW7J2/rK0L44h1C5RBQ/ht+ry6fiOfbMRbH3z
HMCMmyyk+wmhgm2bo1v+AxhRFhh3hZw/6Qh6tPby5wg3fnvmgKl/8wErKCB3
9VBXJ63D01MQRJRznTYb+xvjVXlT3+vsuz88jD7l55mdl/UT3tttMIBwQMet
QshbOvOb1/a7B7bWrtGx/OyItJMRdcWtZ9g91r3ndDEHbyIF4izzqrQ/UiZ/
2FdBBvyYjuN/k3CnPnhh5qBp4dw7VgrcfrrDrg7sB/RqfAEpa1A/8A54R9eN
Ep+Notnm4wpoYNMIEgWxSXJG1CDTRptutEWFruCIjBfjW6CI0q6vIDLIZSBt
sdipRz3HK5PSJlF20lFk2OopGHlFGlhdPq6m7SUU4f3ucvnhP/orBssPCoRE
/07w55th9XKJJ/latRUrtU9BrZmWintPxeTCD6ykuLY5heoFgVztLZPg+XdX
lOJVyKXITPGxK11SyBkeSevZBw79/GkJRmV5d1CfTCozJw0AA9Dpiko/OrmO
f4Kg3MWM0nhWsLhkmigoB9mGfsWqsC58MH5FzuvB4X5v/luig/fY8PSWM3dL
S1E+yfWfHc9DbOyBb0aDaZhYkHqUz7r9LAFQFVc//tEEsUTUCZh37UghA6FW
laZkwcR2TnywmXjmaSvKvRB3IkbRsdVPNPO1OTeatOtjmjf7f5rpAXpXCg9n
F/P7KcRg2wLb5KLoTDlYF900aA0DE1F/jukZaivCAn7ovE0LVeeO6g8OEwLZ
ktUjvPmwsT04Qv+Zj8DLu2qBCfh59Nm5kGrI50MP8EcRQOHVug98v9HXRaN9
CT9OmhHT9d8vQU3IBSVG3ng5YRQiTM+jEqqgfg8FZ6UsyxWrfW1f/5QLvR4P
/aULvVhj6gkOJrW3+ZoVSfcw6Hr71B6ejjaLNcp3n8bvVa0q+j7INVhWwZt6
d15Ues+VisXHmQYAY+3Eaph1VOCnZ1rFZw+FKtBa4lGSAb2+cekHmyvf6BhV
F/xS1gCFbE1MagFwJX0ZnLDlIRKyutXp96yaq0srO/Re49ICcJCfZhf38PIx
XGvASGISvFBOODipV6tV/jS3XPKbVlvMjHObjRKvfoRhR0cnUgiBInAEplg9
ke+vRSuqh4fU+PNSMa8Wb3x7IzmhQLm1dcYmY5Z0g9N0pK891mwQIcfKGnV0
+Sv0xsMB9SX5ArjfHu9gP0MfQR9f6SbXOr0ybDX+hEtBSnzhpbOERPlq252J
o6P2yXkQ0naKAlllGRS+Oy6Zx9lOIBImxvL6Yfzdj6WEDu9B+AUyhzVyagAm
H1CtCyDwCuwAcDaeegxWeW8+q8+aMzH2bX2S7jRvi/CSEXAgvAHELaGzCchI
Wnn8HuXUON9OKNsCC6COvkrlu+zBTcJ8dVOErNm2AHrSaf/AxI/S7vaJnlMT
d0XFASuEKlBz+yftATsPlm1pfY/Y+djfjX+w/Z8mIB6mg+zpXw7AMvoBWrwS
OYIts6L0qXWC34rNYYXXo//edhbBwz6ExiDoZ4s9UtSVNn58L/R+4UstHs7G
T+mvkmdPVUinxfdEoTLnD9W+//QzkEGTVnQI8UNOh+rQwLencdmbfAj/zl5Q
y6OxJ9b0fjbRwpZdx/aJcx8I3J/Nmc37L7ykbOlQ1CVlr6mdW9actZSbNQ2L
AIdFWvemXXkHIGdA90xLEH8Wu0kACdc0yuzXqW+Z8/3UXFIfQBZzUooz2spA
uZ9NB143aqXZY203so/mv4lLs4CKxl/QUg2SnP4S5VhnAQ75QkO9Ak+s8Qzt
tIyIwQ447hy5dD85JfR1gA5v03XTSOZK0HkSESkWGKwRIYUl4gZqbjNRcm7u
gH7cu1Wc6P4JW3Ok2r+LHm08dLUkfZZ0U29iIsjSFvV8CIt23Zak9ZfishUZ
KudcxmBzjO94fOIUMU59vUpVK0le0KkvMPGMZXQ0pISdP3gVxHBnBf7WUEIh
H/N49bZPXpufp/hyu4Fv9WnAytys94E1t8BVdSvzxApSvs/T4u+zV+ncR95H
rqABDqmFVDTXahgVI/udpT5GxjPJHPbSpWfdaSCFePvopSDV7M5PqNvt4tFi
mb1oNcdJl8bKPTfmBuuZEm6oReb1HXciekU5PGXjR41A+WJpvy36yagDJrvn
ye9/7wTOcUDAlerhsSySEGGodXO3VaaQxSSi280f0wJfHmK3RlmAVBcngitp
WRSjD+TnA3SK9PlSFZOrrXJ44XtRrHEp12VFRaWt3HumHDlxZ/lyezyzCyjE
gNJW6d4Mn6vWCWwNLikDQVonOZq50oq/WRJ27G/5c03RGPZ2Zb/snkylSQ86
7vNB3Lw4iD7Uk4eqs184ZB6yE4ixLyGUZ3O+1qp+/D62ZLe9BglnWm7KpVrM
dq1hkZIBB+x1T31TUkJnA+D40LhlPuKgDClkIwzIMH6q8d8odCJ17yPLY7t0
S0KQ+HYlOo53XiqWTO7Zf4/HUwGwCxpd8S+TehQIZDiDZ1HIrCWoiBY68jKy
OjISlQIINq1otUVTap2XcLkuva+8gjQAL5bG2qeeS2EzELN6itNSblxSbqmQ
4GOktPMx4e4V9JAjIzSjqPvuIQuoHe8Sr5hFKyYkckZRkgzFHdoNf42l/kwf
IC44qq9DlXpjwDIFoQJ6qQbTt1EzAbG6TKReKtfh8ft6WVYeuyqQON1zWC76
TkvV5UgXMLvciOQtliOXcRPYLk2Lpv8GGLixxrAsvyJ1nPDewlLlW/Ib95ZT
21xxTPBAg8d/HnxIGNmf6vQE7ZBhXB3XSGKeua16kGtrD+SMBj8DB6E4j2j7
/20qFgT95xx+NnMy9Bpnh6RbCNZBE4vP2PVByPlDH0U03Lg//L+3sGH0JQp+
SqW6icZVrDH1lyNivk2lHmzPsXTqsQFF3X2YJjDBscyBcodfYN1sDd5MhkAI
soHuNTu+yWtPiRGEEtdPYJRJlhiku64uGp+OtP6AMkw+ZbQApzMBBEx1OilF
Vumbzx1VFWtCZYJRVXykstmo8zwfY6ohjMzbniWTgcAOFKwVWqLQAfr5XYWU
/IO8tkuxH0dx3zWSa9BuoFWNRuuOsvGJBuKNP/8kPGcathN1K3Q5k9JrTudR
Dy0mRasD+w9K+G4rIxD1ACURGzcfvN83WXfhtDfVro8UvPRBC1/PhNfImQhO
uzxoYB+UD3CbLFfRcZakVObsnZY/DI0rpDxJ3FEs0jfS33sCLMAFYNC4QNem
4P2o14+zhwIAFTskXERTxAYb+KOVeZyhdE3SmU6uulLn1H93+NoV9ZCJ6Jml
FiyM9sehH1gcuzW+Ns3TSa7VoomuBgiu5siza2NyC+foD/vrBbBddQEpVMOL
R53ybO0nS5Qv/IprBFvfCfSkkC29z1Yv0ayGjWAfLp9/b416PFQsl8I6xTwY
/DQ70Uyl7QV/rQbyvOgsZSR4iZK/vBbhv86KyZemh3kwBn10hRiNqgJCSUMg
xD0QZy0oegEHY3CCBp42sfDoCKR33g8SQVRgWDK14MY2BYcGA97v6lwA55M6
jjEO9MWSGIWvXmgf5CFCGEKielA1rtg2H59TvVGc4w0JArYXD1Gh+BDu2iG2
AFpX4/OoY9T2X3XVMi2/m0H1g8VO/IFRUDQlUcNhn1a/sg4+OWqME4JullQ0
QvWILVL3ydPEby8VYa0CsManN+oxObBnAfulQWTNj8ML4lvRsHQUc26hXWxB
EIiCpbryklgmt2xQk35DN7yDIUudbPQqLFYXRQXcSpBaBcDyQwwXM/D2YTE/
gCxchfcSe/kkxyh6yCYy7647q0rawWigMGfFxs2BSB4KOs23sVVf1M1sgj0V
SoV/IbM+H+MMdK3mN4ih4JRytF8za4NIaLMFaSHc7+uPCYF3umxpTZeCpQYp
po037NbEt0Ec4h6sl+W1Ak/gdwSY8uxz1jlH9OGBdBpa8VFgO4Ba33D1Fiaj
1k22TfarXgn4GwG03eEPYb+R1LQ51F6D9rPRHeA22Ww5uzgQ8NiWHVgfloez
MeViGYa575C4KtE27lnFDH3CjyG7YM8hUmKDy8dNITyULqn3y0Vn+3iu5Lqi
4T/fLUp9wqkQ5H7k1U5TfuxhA6E8OpO23j91kk5+lFoTsq05KT7lHYGHzvqJ
J+xpV//Rnj5VzSuTUD2/NI84EhmwXPneXGC7qXoDXsLCXy+2qFfCYc/WLXiK
9y6mbboIfwS9Li6BkHnW1Fv+8m006/W+V0F8+roWO2dDhSR74H00u0Ti1tV8
IN2hMBzxvNhCXBbhG1Iv5EQvhPIfh0JeyjMa0M4GkBLQQ/meAdX14fw4imT9
O4iBow1ONyNL19ZSk1xU6w9peIk8H+JQQ3LuZL96RfMmg0/P0lCL/gst0haR
7yGcqPRGZy9n0nBXYS5AnjdB8I29gTR1r/vgkFjuhQhlcDYZMOUN0/iSfOGb
iLdDju3brKuBbaHagiJDphVccE3zbeGazQ6ojquHKzjwtO9n90hm7g1L6iS2
I1XVundeEPGc8JOmIYVfUimgWr8KXl9Ybk++5vMrgbgULERgAe9TXTbwXSxz
1tL/uAjAFxV7tNJKmIUQjbpH75CYy0fq9t2tcFG1bZdJMoi1NR1MP/ogxMBv
19+vjMwikRW+E08fNRU7htjDwgqjwvGHgqRdcl5OQ2QQkNfuBXjRQXJfQIXo
3GfecC9zjDS589fO93rYflzNwbCHK5sDFFj2ackyMd+joHf56AuDiXO9Vevy
93pq8f4Ys9vkjq7Fs7qDJ3D/DKAGeyoJfM3PRfGlAK3mWev9r/l8J3h9VlG8
eC/1ZQhNmn7kHLecXzqQBmfmIRO56P1M4Q4zhjBcDpBdN1KCyQzsCzQSX3d9
NOxoRHCtv87gX3Y20MkeQ+reXwVTIhOJrs+Qh3C/VVglNHfF/Yj5CltQU7J2
nbR9LwPdF71Vu75+0y8H9tH2qRPF5w8Rox74J3owat6TRCfnn2NsTqjxQbxt
9TW6HQlM/L6cF7y6UY4CSR40/D5MBaxrkZ7Pems2Syjkh0101ERl1Icl3Tao
ZfPzOHAFSJNQxegtjL5TR2a7zS/MFTQErAPdhjOKtiL/qYc3VP2IXAOJLpb0
XfdiQRvOmhyHQa9Ivqt92KINsw0DQduhvOYtbRl46imn4Mb/bEMLf+b2mb1v
UHqdPl3F3d14fQTFM1yqo4+uLSZQ9jOyZ+NJEbI+ads8prLw4z0aJq+XR8l0
LxTMCWX8CPctFeFa1j62lTrNp3SYhdXKp0Pul8qGadQfD4j0KWBjayhKUVGg
AiLqmmqyE7eX/cYuWJbXQd47coW9TSAojfq46DK1eR24ERVOXf7sUTlfPEpn
Fc4YwMgaz6gdoTRUnMSVAGJ9ZBtMAQXeG2ybKv3HafAUwx0+XPkYdxDIGpw5
l/6jbmydNPA8JbopkykgCgmkzSupiplvEScvLk1hWZmUvT/jjrMz3npe1Qcz
KsuwbBh3qTs7JWkQQzpjQmrwc2EfRP5OFZQSWTUp/IO4W7zpEQCvpi7xPm6q
6X3y/EoCL/WY2oZ4ubn8tMxlbJowmsDn7Gtg4PTEMIYHx6mIftRxQmsvKIMr
2QO+bMn0BBECvzdWHX0wu9ehrRt6eNBuxoFcwyTopf3ly731gkp9MldrUab9
kbZf9BWrdbb0W/zuQw++IQCM/BZaaPWOwcXQ1taHnbwZ7OtxMLBhgs2GglMA
tkOShjuu+gNSl7olDAdayHUjR7COpDn1sI4f/xlNjQ53S2DUyYaNt8dtT1pt
iQH3GbHUQ7U4qdBCuL+vipJu5/Q/AMgaLS9xnb9/8V4kUUAKtGLTbjuW++M+
GJXZ8LluIA+7+C61TFH5vZRDMj4md7ltVZcYVSLM2DRzyew9sDARTtKpGLgG
kpCY/CeTkHoswVWh76mCVGtjBezbbLv35Z752QnHrVK/bt4tydHol8c8XVvv
IUr0yG6eSrUocBZVWRpskw1NHQPyvC53vui/ldmYscFeemm72nU65qZROGxs
VMurYOoK3g/k5dV4tYX19WbcgWq/CFx6fqXUXLMSbzTYK5avWFLTJphZxWXn
vjJnQRyx9iTcoLAZOvzorFI/YNud63MnVmG19lfV8onuvkuCSKJuBfGF+/KG
STfCBRsKN2PK4lnSov5lyToa7bizCv4lAIigZKLkjt9NLC7SH0BV9nIWgBBy
QY0sfC88Orsxvj/WOf2AEPfJ4/SxH/IQJwEaigNXaSu4az2VDVLH2JCi9eMm
+PghF0qkow/zp6U80Bmychk429fAJ0FmH8yDr8iB7dlK7WZfULcs76HzPYoY
akP9yOs7b4skWb9D16Vc7bBJqGesZNAn0timV8W3fqv1a6eSZLd64ETXWgvE
lPrxU3GQiRahRnfqa6S+A6CDDdtLm2nbvE/KqVwOtqlp8h+y/baaQOgfh9fT
3IlVb4lgZ2OfUqTF/Gh4+6ekpEiJ+56rOSgzHJWqZIm/39k5J0A1IEG++Xa7
wiDDOJx1fKno5S3XM2j2tEloNYUhrpOP7DFJrqfAkq654sPjvTpqXmXbT3bv
AJkRWwwx0it+01HrUkMSNAWlw3rJfm1AxV9+ctrkaYtcSzwESs3J/Rg7R/rt
L0q36qszLgD+6xoWcrALKu11qJNMulG4gRx12AmJwiOx0e5lL1ev28SqiaBf
pHSbIhybe1iXy/zrQca/IpXQk848cbOuflWbRqwTJ4JVcowkkhso+Osn38EC
niSELeVcrW0gTq1xKlYoxw9o9v5Wb+pwhx2T8AC/eAke2R9Mynnd5/RwBTV2
juF0kCGhrLlhYukCS2zGpwg/mzDIe5CSdY4j7r9ZUsuoq5x6OxoSHInqQEJ0
VOXNJzewLrLevYgWBt1OhCWPz0+TAZMk6Ds5X+XUqn4beSP/BQ/s1oV9JIxU
W8AY8r0ZP9SN7jqnv21czIIWF/p6srLMgXjYk8il1YopiYaFFl1xtw+bPA/A
c+JCqeTVecVVEDe/i+hbiYc+lHBIWKFQa9UWsaAd6BaMoJDyT+JnGL6slkml
hdoedJuuqFM+gP1pNm9J7eqvuEasRmhlJqmq6WQtTrBCFi6VfrA7GUTBTJwa
hkF8ooIf1Oz1sW6GBTpd6H+LE+q11HVAhgSfwYRwY6YKMBWfR+mlphC5QsVk
VRzNwunztG1uoSMjRuZrNnQdMJn4hJ/UwJYzUYMmu9koeMPFBXZoNgUxtCND
J+nxGn0t/ixdM5qB+03uMirndHhnqGr943l7ViqqwJBxpgBhJNy9n7iggh3d
hZPwfLU6J6gV+VbumXBWRIuO1ZxKHKlP8iE/smPgkvq1vkS0FmZt+PxXm9S/
qhKTg4olQsjEOosabbXhvTyHptrjpQ2l+N+Is0O4PT50Txeo/e+CF8r2biSP
gwOSBRBmOyKmXKsVEyTH2NLxfoehURT7rsl1QB9mMPQQT+Jq835dns2r3ydk
LpypkhTykOuEbczesAwhjIYBigxxt+onHwIYpnR+mzI/lxbphNJw+8azesM/
VU3aMWG3F39ynT9QEwmCE3s5oEyopBlfkaqK/S5wHiz/1320Hy/o0d+0nJLP
TpskwZGKrgeIekKXcABDuYcThSBLSXSBWG5rAUml1wo9KqePQjNEzncF64PP
lIIX65IvhSEYlla1zeGtUL0BZsgMFV2eLq8BTCi5I4i7U1aCvc5joyRRtDR+
R6kYQwhb8E9fHV/UZ1QsRNf1GXjBMtA4tp84WIm1eZklu9xgDdyR5gKz9ian
Y0lAMhYFz9c/4Flv/oTcd4LgABOuW7Kgal18venbL1fZds0E6K+UoOHdllp9
zG0YSCREIRf+IyS3HY9b8bJmj91CHrzBF7vXdx6mkXj6ZA7Oc8JLSUzM9/VH
/pxZrlJeUL17ZPIXLPx17hQMIDWWjOEJYVUDXOBbUDl0W3GQ2+k6ax7zR5fd
ekjZaNoGfXGr47ZYnYleLZjkWgBcfiQPXCYVsYidmo0ttML/0Ikq2ykFbKpH
deDeqm5kDIQdjrPQeNr84uGo3wTuKS1sb8po+U4uIZr8H4S7w030N/8GJ8+u
mZ8dLtzM7UQXV9n5qolNGiMQMmfBWkGAyVsIDbgIo+BCcKvMhHb+KB9HufMH
50kxNdB4O5I96l59cBw5slKnW+nJPvvzaaSqFToZHTJAR1XOddZssoN3FVij
KHh6xeimawEM3ZM4MPgawWXsAlFvo9z/fOlrPuDQvu1RfCPSn7Bc5vs2bR3P
JKtygX1Z/A58TJfDbqD8ZA7uMht1EeCYnmvIs1zT3qzBi8OpTLQiBAKKPF+O
NojBU5/WdR6UXgYfTCi26eYPdOg9MNNahXbxApCm2vJTnRNAIlqAPLsjE5ly
HK49f4Iv6zEwziLW4t1KQsitpdSewoxylbJ8O6LIMUw+STKgpVxes4n1ndNe
yTYaFMXmgqYELWrNdsM8Kv9XdVvm+UqpbGbi5UEe+jkDRKGSJ5d4fsByOeIY
V8OYnjgCKeBaF4uNZTHKzAD+cggqpYNgJljUJPxDN8syGSF/MCwoUhFZ0Tg4
oYoWQjxAVUj7jX3uoxIv48z7qrtCfl+uiX7ArkIuvB6kqpdZvra2tg1Bigm/
NiDmf3dXYfSdz9y+zk5bvISyuTPxg/j3WCiX2611QP4XWHRw2n4HbCd1d2hb
eCEw8objnDNDp+xz+HlfjbzOckEKwY6S7RVkhZJG6/WyZgqJ4I7CuHEAh2Qd
2PzR+MKFK849EqerR6naJwEkCJBok4w3hsQlzrB76arOmtDjYEPWUl7wxRY/
S1WY67v21UER7bfY78NGdVDyUdP8tb5+9ghrT9r+KKQPOWduBDNAymsN4FBS
32x4zDMxlGScd+VcfM3cxV7XoFoP4FmYtszDCrKtaDO+HfA19RlpgX13h9Vj
ffK2PGSoyX/p1Bsq/y5+YNTyP0ItEGpUVq3Xw6Na1UIb5/iU5VWRzhKPQ0sD
cJm/gWWtUqtwhkoI+CIuKBFG9KEdZ1JgD55nIl8LmB3Q1qH5e3DQNbkkH32w
sqqK4IpXO90PCOWx+Nx3Pt3sFJ6aVsaFPWA8/B7MqdHrC0mpSl88i/gbMuvO
IPSuiiZQdVMhPD/NHq7UK8Y4UKwRqlTJ1X6Z5P6b6eP2BtTSmc2A0e6zZLUA
1NhzsWdTrDx5hc9QD5yOMfpa00M/h5W0hE47O4h0Nwsx8ol4Ra+4D57Pfg+m
7GVLTrxWIzNhj2nFBv6v8Kd+7S34WVvx6/2me5rpnJDzwNGg1oR5JsPVj2Ox
eXdjdhFYwvcfVbcTzTlPqDyqsKFlCg+kPKxnBXsD9Gamid2+xbKi6eMUjdgA
quTv95GQY1Vr9FUqsJkEJftk/bmFQEttPuD47AETfkxF+O/NHglTBCCG7iOz
wXTglz3908uJtWRRYKv545oYxp2QLqAOQylzTdrIf85mko/wRl8GSSGYHrp0
DOYHTEjbnaT523dJQj28+p3g6DicTCExgYGDXVTsS0zeVBeHiJapQ6onME04
6Ld5peAUyD04q2JmdvjXDdJYiQBC/PyruC6flSXGPgWgz9wqO+30tkFXmTyz
ObnUvwcMR18KhkMBREsWAG9C/xMP4eOdEuejnendWOzPdUIKy38sg0jd6BzT
HFXVDfvj2G3uQDj/N0YdRzoYzVynPTBBx5WJspfMfZoPQeYy8otMcwxE6yqf
YLaabZy43/dtQuZuC6JH3WOy4RMS87fVgWuWdj/t/VJSHEUWcuVAZAdNxrJJ
JZJVZcYHot2fkxReW1kKvvr/imQ47Lw2ZwuXPyE/DZFxSNYUWC8SkqFvfaad
W5r4AB66s0JI6p9f84ibmtR2z2WWPTfwNyjsrljDgbHXGWKwN7Z7aVGnfbkS
M/FopYZIitqunqjHEvEY6IDFV/r2aHX57WEfuCKi632LT56GmOGSdt6v3Bt9
ANtt5hKgGwbU8DPbFmCkCoPh0Rf8q7qZivfx0FuLKqpnUNsaAlResL5pqGpJ
ZHtmu88fB3ktHvd8Te/++x4x+rzVmx23VkOeVpB7FE9ml2Ai/egG8++LFLq4
4EzB9gI3S5Jbcdp10d1YK77TA7FrTg8ezssMAAJIOxDoGNEI1aHwUDEyzfkF
VcY6NuV/dzt23K06AmVhThiKw4LNJ57RwO27D/hypniJy6TFRdQzlnvX98US
hhypGOoCqi4i3+Ns3MyJsE6M9OMBe7aGLRLia9rgcmTRAjVAckiamVGy4JGd
TlaCPQjYJS4L5k0b7O0RVii/SG4a8KrHdJZ+ZZf34eABZEV3wumMWZYdraGY
eKFoU8e/NOrpsl7vnJzeNIUND7Jn0wnsWYji4r8dRaFS4ySxZ9AQxR6+8ic6
t+7UZ8iV+mI6sqtP55n0wRAhMUA3HOdN3+0IzDFWWIQUms1hMcgAQTtEnZ8V
/ThUUw88X4k8dD9wRh/YI28nexff7P3dMTi3jF9UpLkr5OO+94LOuQ6NS/4Y
HtTCRSjBoTfMUJjDcxb46Kh+QxxQuexrJ4lD9QIVB9sbpDgEJKe+XHjBjdln
3tqWolUqVEmiZiY/FWkxISg8/OfJf5NZetcoaQNVsNl2bZ6HInizVoMIqEGc
cnVVV5zk6o/EBZBthc1LJuP++Wjg6foaisShFIu+joYkGATIHH2OhUlZp5us
wo4LrELDtJxCvx1nq2QdUdM6bDrgWLvHQabDyiN6Wso0blU/Wpx323iuoXov
PfBb5VyTvQFGMzJDza+dI/LwuK+7mcBoNg03pkBJleOIyZpvl0BpZL4/v0QY
EcMJbCFbabDXhOg+05Gc6gT7l0uD74kGzSdvkaN9ZMv8wFPaI6TiyaU/GuOB
KaDYY9y+DkEg6G9x34uZXohldbDJ91eWyee0xJ8yGPAnnPFYgbHMXQ/who+Y
EL0CA27TiCPArAr92O75fWzILBgDPSgaz8pne7iQSFcP2YeJdPqQAYvfMyVJ
/jR9rzsIAJsIp2AnjqVTaruYhkYhe366f0CpKwPUfEgcV2lkIQtm3jHIOrKl
t0uwt5/FkRuxxpcIdJkbUdBHnbni3V6KvVuJ6ZM3aZUefBCaVRBbSjwh4r2g
kNjRwfgD9gXyIL6eTNmDaUMxXsjIYFEhLHvwcFOeKuUtmOHEUMD7Z/lOIkVr
+gibN6YRknEjYX82M3z4VXBPsYT5h6/GhyZVnu3Tcwpm3+z674GwnyFj4eZP
TfMiVxEtAVFxd+tY7FjTSMeemzThpQn6wzJfQ9Gp4TlfhoeSNG0wRm2m/HUK
+8k4AI4x0b5YmTOlcgyq5gLRnEDhg3tJmxJcEgJdIE4WCl4LRnhMNYY3Zjqe
sgdG34y7iSSUt4oItcOeHa/qq3DdLOmqczEauBYN0+MdYLY8RndmBPUSDhZl
wcuovarUU38cd+TApoWxrPpJHH4kpSA2JmFWg4ph0X4TGQgeg/WuYZBcf5lb
KM0UUlAPQQjP3KePPq0m+0aSe7b7eOCRiZbYjzMza/HzhS9LuRKo4M10I6Af
G6Ey0FW3T1UymO/uB+Zlhy62RDJsMf9UTbtVNT+nP6Ba6neBlOWmAaz+1TZT
tjLr8eAfWR9ALdicxZKDwfLLKVxnEXuIO3RYgIyTG/rpONQ0BiFlIlCvP+vL
NlOZR4ySpvavi0ciOUcU2gTwGJsRBlWxwM3l8a6GXbWpOyOyGgP5uSUcD9L7
cLEFWDvFLizFvGZgyGjIDKHlb5yKiOwyYpSGScXwMO6L5E8iSU2GArFJnS7F
I+SJQl8UxwPKGrludelUVbR9/HV3EFfRpIgcLH0p4scyD3tYr70TSsNjwswz
nFqawXRSxfDcDuFkB14xh3vTH6USVbSeCOh4rlcDOJA2cMlErfl04RJzdBpX
4wzn1lEAgc8TOJZCWQO1GWwoWyc29U/RwVzxqbalxaMDIKP78XR43AtOEsWD
+0V1/NE7Yo25aieTTBf0E5rU70RPhvNPn6dTZWwj5567ua7gkTMGqmnkDMwn
0Qi22pzyM3D4TPJd/Rzcq+qrK/6GZsUzwVT18deWKEP2Wiyu00ELHytJtZ/W
7+RPpill4J4BpShaG0vqeIdt53WbcWaS2QcM8mHvVu2iYfqm7HLYPD3/TsA7
ciVeyfJQUbwiz+hkdJxhhVHw4TYBAodjnP8T2G/hfU4mHO9MrzZYMg0WCIY4
t0rkAxsXRlaQVO4KKMXJw51Mcz8GGoICPyNO4C6nacmAhpBd4dtPYY5VP0qa
wGMmVxy55rCGKJYZwTTk7KLdrblp57WlI0NzC+IxFLXUpRJ7toNY/eIIdfYe
lOvl2WodwYmQp7wc+11jP7MnOmeqsPJbSr6Y0ZxD4tnKCwq0JZGKVigteD4P
csUtKn4GVFXBnaihSaodrU4PBtyEWmxDCZhTyzHiTtRnZOu7gqbPHiJVz9af
LXS87dXh9pceqw9XCAmz0Rj90+Wq7bMt/08PVHwzQb3WFn1xa7KQ7i4iz2Vi
KrP7hX8yAg5epxW0keOPHdk7HWHbIN7DOvBKbazCdEBmPCfLx/EIHqg2zQ+b
9w6px90HjmQgXKcN9vlYDaAVsZRYuwtnD9I51quIV4GhK211TT6YAD2whq6f
o8q3xppc5LSA44Hk9wVVIfZgVp/4x5wmBQNiiAetcoPfETZeDy3MzSmKN++M
S1OWo/8ryoYOE2s97ycEC+8lS+q48yHemQm8LyqcWW2cMWXMAdknWzCsQDPN
LJmB5IGkniMwCvbYeMZ+QBqFvuy36IuvhC5JNsX4pzZyaU6Ny4sqmPPndpOw
JLu5jrn0fGscXjjn6x1UgzS9t6r0fcupn+jtUB78hOGmqP0nPGZNsqCLtnFy
zw95F0tuma3dc9whnFvZntxwk510eFkJ87Df3R1GCyWPmr5heZe3FVlyWSsD
FWkvi4Z4qPP9S0lXjPVJg4WhwcBXFRh/6p8sbYzofW6N4FT4hFXMY6B24ob+
sUxZN2zcqO4kPtoU8VlZICMdc9rZsnjVSxJqMCdZZ6utIAevTThn2H3fjKEU
hw86vjxLF4yjP21D7kfJDST01xiupVEpydFfDUhcaD4dGTTCPy9GdyjzJTUW
wMgzHsTnRgJFNdAHcPYXsmEVPSY18QjFG2iKsj+D6gAXj0cit7+e1HNRmsZb
eSV+wt0/GcCdu6XF1jQR1vR8BgtKCi+sOSkzxj9sQNK/zw9m680XAwO8rRhT
Kn1XeOGdSsYNqPOsktihiKCaS5ebi00BoMQIcT1K2mKubTy/oysAZuUBd51v
k7tfHP8nDSL1UIXKmiY5VWIe0zOkSlf9vSPYroIVAN48mXCyHAZNhruq3dsq
tXBWViNfPlUsx/nGCrdbFqLHvwYU3Kx8el/oXWURZ6r5RVrLnxqS1FoSAKc6
XnB+DWbvyUtfYkso8lIgWYw3dxV14X4NSMDeNoPEZR1W7FkNc7xxaES6lYsU
NbzCNPLSILzM4uLKlNYejT/oA9day/W4x3zJtfo13GcF72fSA3hIIQvSkvBy
QKi5qFNehTzMpKJLdyQ54MnPl4Ymse3kQh661t+4Fjg878ZOTuk/mPTL/f3h
dXs5NyaBXVzdRVCsuU6Y1d6h4Z9dGJruVGLXJxd+kqaiBfjCT3N3bUfayj3R
n2an/XXb9zF33XX7QIhBt3KhFGZ4Vu7cgd9XDhhuZ+76geRpFz5v1FHZ/LV8
1wlcvt0x06CqHRs2uNYTizSnirP0xQdVjuczofLijqdPV+1TjjzRgAVJgSgU
WNm0g9oOEwTlZFY8ZrQc/24aD24OSoI9U8YVgMatqzqlM7ZhEG8jyOFrcvK+
5tiCCuGK+H1C/+H7YbxFnv7xzBja9B8BFFloy80LgSWVdk5clFJVzE3+Zv0m
DVIX0AvhwDI5RuJwJM5Q4hX55Zdz0lMjvD3+DhW9X9ZQamVWIXnd9D7g0mLC
9w/Xc/oCHEXcksLPaNsGR3QguTTuD9QQY07wrB/t54uZhZtOwWc49drg1aBY
ToBLuKHuEbVl1Fl3N5qE5XzNO5KS/O0Esixe4IU6bJ2nQQT0VKGzzEeJmmpL
u2XQ7mRgWQYFcqktNchN+ripp4Z2lOE4ffIYlO+hV8waZTlYqVf2Bd2/Ws4D
/SvRzKhmq2ntizPd5LQ9ISNTXjOAflvSasjqJXWC/nTowFoPd6nsyIlr58mg
oEM3nFPbbC6UnfOrP0lkTtmnE1EZ1ZmramaXF26iyep82cUymK3qyryUYlkx
6Yf3zDYiLEWbs3rwkLkZ9+NMIVnGtoiwyy2sz+Wvwwmt4ai9lPDJcIWHhMtR
r62z4IHwmUFeTl19SCT7yAq/Be6h3GBrwXU84oHdH3U5a0ERX+98CMESiVcR
4Z8FbqhBiMbYjBBlfl1O0V43x9DDsXvNU2QIhUmikQf2jb9YOO3gEwiHIUs3
N/77eqycmIBVIRvm/QUUNsWKS4O1h12AF0HL4kgOPUiGAh24EUYTkO0T1pwD
cRnFJNK9+iDi1hnUucgqJ20/ev04z5K1frGqAw8FHuG/f1ZRKcUck3KE/AhV
+TP5JCLXbA5F+/do8LDVvSO0rZ656hNhyX8CL9lii1FpqZBrrXs/KC5llFa/
EYxoX0P7xC8xDT7FvDIrVX6OzLkpEjXeoE5m4wOV0gRrRWSZGZaOIDBnW8/u
tRzxNnBW51BfmdBzBOpppj7WFctHjzRfC5yzMpKaiY+38wIRbe0vJuA2i3R3
Y+cQHxDt38zSbjl8Dn70+tcgdnrZohuMAopinXDfAY5vSmZiB1AAnHsyx/au
zQAO9n6ek4E1Nd1TsIBzk1Bc74irx6MWvNgbtpqCf6aTbsAC3hpUpl9ydG04
X81FNe68dN9O3Z6rmBrGV/yth4vhIErNquNQrkywoDRHINdZHJwuxT4gd/lD
/CgNvJc1igIfiw6/bKrqC3ZiPM7UytwDN28Aj8NlDbBwzz5AtnzuSPVIZewc
3aebvtAR1On+QEZX7+nFRJ+VNJFOks9tx6XsJI87Ezqxy9TWTqyC1YatTM+K
+uA7FR1MX4wVU/1Qii91vTnqkU8WhHEHrNU7jWQCdU7cO0ql9SaK6b9xi0qL
Ygpp41llt35LNTsBA89IKOE+DjOJpBnHvJf3Il+7HUC12huGgE6s3OtAMVQh
V3/qrb4akT5PTuayZdXX2F1kAS4xo54shywxdxS7qUyNRMjmt6i7F+6RO6dr
p05Lw8kkMoTBJsQNLMy97C+A6OWG2nkIKbru6p9/R8x06yz6nMvVG/gZ+CMz
2ZRPAKhMD0Da8u/FOIzHR61805UD0nKgZcPkhqktw0sxlkRE4zSgIqbP4XBa
i0L3hZbV23Us7HBNPXPSqIafntE5xZZVq8LKNIzfygzoB05x8eLGoiX017VH
4DYKFK3eu2kARBheIhgg1QZfoN74V0e1OcFkn4NPQZe08+NMNf1IhhQ+6wni
CoVM3R/qpo1+9Drs181OmPPo06ZLQRCDaldyvoIwNPnWxVgGlOd10MaENQXs
7DUEfUTbyccMD4UPZosc3Ejv8bxa6HR5JkrWakJWb0FW+xs7XsZasA8iIkoI
MnBoM20msxwc1cFwzd3rUu3gBfuHHD8xyHe+a6MLiOWUyN8mpo5zZwIq/ikL
tMIpPwQLtQic1OQHF15IIP6Qq5XXHABgmwkkjf4sHD6DBT6YgpZ11js9iHn3
cHDUqMXuSYMGMENoJpxMY9GcRlJ1fi54csadvGckw6t67jvQNFOTz+rGmDqP
IjqqThruuS7bWwLOAGri/J7FC0xLZhtRBGcXZtxmGsymlIwWCulINIUDC4N/
RMDWWdePSu0rC6FDtF/LH8lT6gTHJGxyTBzl39IYG1u8kjJ/dHQbDMbHWlOC
JKdKKT6Ew7f6FsyjJ+WFczG/P4sVYFSfhfPqdJINxjz4JvxCg4jRg5Yzl/Ma
gPGdijwKee7uVBUkpTsYDerAFnf0rNReY+U81PrVBxYnx295kORhBZMsSEeG
TMFJWCJim29A0a9P+hP+sLhJyhRHTWO3dLQvl8jlMShun6UaEycs0hxwa174
PRWymCy42Lv+3lbrCoaQd2tgrpRz5r5/AZKSwt4Za1VPxqYBxVjDv4aO4t5h
uhrtGqTTwDJLAlcc2ez7+qzxYtu3s/E9j5q/Q6SoH1yfPYB2z1Owr0W+hufY
DDVEb53wY2y3or03jTiCa9MK1hYeGVp+pUQXN8apKog2h2Marcc4ed1EToUl
iU8w5hqKzMZIuUM0MDHcQpUDhYX9bkHbVuZlepnTrVsFuHnnsfg0lxSS92F4
eu1/A0pmYfPxNLCeXS1L0Gx4Rvi2ZiOCpTnT0XsGS3hDtqJaEvUltJjRW6pb
wIWpG/PdLwWdkl+H4L3hOpOSMhWaOEJkayEwrHr7GUDe4juP6BVrWcpXB7F+
fG6Mu1YY459KTlkzYGB/3Rd9k+iJ9lcg3/tRrj11dUjhrdyKKd7MckIW8VWo
DxL8EMPruSsenuUvmnMXPpL7/xPDB+eEjDuy/xftGV/Jdbx32Phhsa8+gY6w
PI8sHTHPYbZ6ayo5/dvWRcr8pPt2tRMKu/c2SudguYNeif8T+TAJQ0R+JquV
wpstYTiPMP2GuQ8hLQqijtg2u2ugQ9xz/3hO4CMeazMSBXNag/64z3jKJ/Ca
5A4YsJk7cZzRxILZKEF5kzEIO08W/V2eVJPBKM6LoqOzA9eNKcqbOjqjt12O
iAKKeS7YicP8KPsQqGfytF3tHY6KNjRbUFjL90vVoBOMR35dUYib+DwKQNef
0S4NfvcshADsd+VECcDQWSI0REV+ZvbaF0kHw6oYGUMuDRDiGrvNjIZ0tkEN
m6rLCi1WRSe4j3ohI5Lq80GypvrrTSXMcQXrS94e+eSu3ndg3C5C8pVlmB2m
tJzjpmurlIjbrHIeNhQ46SYplLH7LgTfQLr5PoH5SaOUmo7+b0N+qkh0gOw4
yhEFJ6wHiA4R/gp7kp41t1Eti+dTRS4xnTYHZqDbux8G1+uTzkdS27bhaYEF
QmVeifCqCPw1s3PiMADW8yCQwMRRmDWVqCQP4hCATTpIehLiehuFmoOqWMBJ
7S+eckpxc4/4spGs5eMaxUN8UImg9h8u4FkmkSL7Pcjm7X/VlAu0y+z4YPYC
xB/sWUr0GWGhfSkKhX5OvdN5k/TAm6M+gFxBTc4SwrbgT3/Y5RYNFgbqvjGc
+Gh6vQqYjSn1S1YFG77d0yr9Y1uT2t/n+QuAWGfUlFNcCdC6F7seqoe51On8
x2jGSn0wOgfPi34RRnIm1gZuZyft7uEwOrkEw4zc8i/qvLjtV6oA9lH+IunN
tFcJzYEXTFBKXYAD0g/Jwo3wwxWDbSnXhBh/KfGyhlt6gwcrfL/u2E0qel3c
wYcuiXGZ8jY6+y3M/NUGmWUVSSb+QW2BmJjaVCTsiJZ7BPRcXpY9qBaOsmrQ
xssdEaZQVf6fq1aw4Tjtia3PgBEJJOak3pt2Omu34gRwP8lk/cpEmHwVdZuc
DO67BI2m7G4CkcxUEwh5OnmYBOIuQodeatxdZqWKC+ZAEPeA2Th26u3UCngU
oVgkj13Y5nICjIBv/IQjzxvCmBBm7fOKJZKoUKDMZ1L1M82uEfBx5usU3gZ4
xbLAdV0xxehe1vHF1/Mrxs43ZKAKWspogbYqBCVD4UEvIvr8SFkB+vlxVFv1
KYsiBmxZRH65R0AQkqMwx0Ki8SNFngKQuSR8vD0vW2scWyDFN6qh1IrBmyb2
XuqDNW6JKKvBVlwr5u48l/QAYQ12smf9FKuXXKkiRgGRhUZrMa6+WMxZL9Gm
QUi784XXm1/Jw9o4jofB+NGzfin8NyCV2oB7rUuiFa7EUfo3p1flgep6qn7E
1b6WyKA7EkcSeOsoCuke9KJTtj2ZzRuMYZN3qjJbvlaneRhkKWNPd7TfwxrF
c2DUT7ib9Xpw8sDAiMXrwppvUIakfkTju7r67TYT10AOmckGVhCE+3oBGaPh
Th39l75aZBXdFbOc407/c5h4mw0PzXFdr+WjEyOlhyHyYziZZQTK0uEMzsGy
oCyzaDUjqbDS56sv8pXnRPOwEruqNTqToTxnxMjMZnqXs9KEAxjXGNncWuiu
K7Rrk4gCYiRkpxYq0dB/JOHI8H7wXuGXqewln802MhFOq61baxfBa3NOkL7e
Gal34X2o1aeHS3xcYGZvWzMtI5z3g9Fzk/yc3KrI7QyCsMLUZD7PE+nEeldt
S9ivP1vPjS2sWpbnu1NwVCa/+X3aAuFpd0GwmtXY7oF+vgT/74DwqKuakzy+
3d0ttn7ZsFlXM/rb1jAERkTicS7FFoPgwE5Ucq+mK4S/P+H7iDD4N25Xqq7X
X1BrwSk5QPY6Ux/Ubod1SuDjXZTDL9ikm0uqXPT9aZ+FXoPvJ51OmNSZDD5+
t96NNdB+xx9iHrXurUP4n5yc19Vzw1+RgZx0WyFkrK3Jtl/V+r/7oNaANguj
/2RundiTnnAPOBQnkWu7+CjsW9kyX04clqU9nR3bvIQwqXoa5O1KE6FlWk/j
XO8HJMFzv5INEdZuEjfHFSml2J7S0q6qcm0etn0DNgf6/89jg44Axntichc9
xAc3+C+3tv8T3wIzpjNZkS+DdwrWiRDQcPBzlNE1ntdKgVuNbMjHJ6hUtf5E
KiwoE/8m06euvHj1EkGJuIN5bTCGYZoHszNU3+bV+9eIhJVqPWWA/EiszRcB
OuRvr5o9en2uaJuGhB7+9Jr9+IKhTcBNNuo9UTu4UO9qkbQC59Oj43DQwB6m
mgD4gscqV/8Pj8ReNqOkNQjvi+wOzq/T8ViGFLF3T074mCmxYYwjCztnL6z6
X7K74GhyICGl8Y/sLU8xGYetlQNEgjqNHEnlNWSIb0WF4E8b1lMh7WH/nmQH
AIQSY0B2o/i2xkx/5Dqbi+InL4i3fR6g3Udt6EE4nh6Ha4awrGsD6mi3HvEw
/DBRBaykI0+FvUWk+0dEyufEl7eaftS8v208ln9CZZpqIWDa+yrBBBMV2TZi
7Y5BPK7/Q/lUjwJAwyD2zDgwMisDUoIZaLE5WLPFHVdwfB0gra2tle/Wz/I4
h8kvI7ovbBDgicUAv6gflhQOTCwk1vRPni5SrwMErHXsaPwWn5VX8YaeiWp4
qg1t5Pe0YAox815IwMVgleCTwRfmIeIdb68Esv2aixvToV5XFoNxpZB8bEqK
SPE+EhncXy4sWUikPtpMuT8n8rh366Igu6cV3hiPkzoZ1ILGdt49grRKZiCf
uXinMBfv8py3JeZoEYIgyGKuXsHezlmB0nQ2hwkfhr3zhhAh3kdAi12dplUb
hYcrKH5KoJbSP9XdcovkXmNMl+UG7hotoMH/ygZQ34sPdtrWifhqTxiCype/
XGb2nuiIYPKyr9UY6SIZlDq9buoyTRidwj3edtoyRzHTeoq2yGFUfHhINeLx
WtKN+JDaWcWrk+Q/BZAnKxWeJ/aHO37u2WhoDri3V8LIGHJNbxt51px0KZ62
mvNzoq+yse5opPZc8n1Sq1sUt5imvncN2GiTLgw4iHhmpDpPoy3B+z+l1T/n
SUIpWJaWf6YiHRkwG6lOQmN06scHXDSVQ181P1OqQ49Zlql3tiACjT02gp3N
oWqcY6xhRg+aJqI/EWxMyqcR6rgmQ+Iw44b64jkLXwgU493jmedmG6Ebcne4
AOoA7LzzvA0fnE1rtlpfF5O71q4+54lu7IEQjIFqsldooEwlBnLL2UjPZxm0
A77930acm5VrZVXZ4yFpc+Bq6aew1ELHI6T1p+Mht9omsgfnlUrxkzwgegYm
lKlYA+wRGEzArMnY4Ik3d2WVi5xrLP8t7W++CTJQvBUNt4Tng7VV5OkldCpI
ndkqcAbOeKUt5bAVxJIu/9PWcf36zqAfNV3btIW6S5r8Fvb3MutCV3BHg/Rw
avjmVaYPBoy3AnX6VShlpRWE4pJvVg7GCXzhUr3+NwnTZ4LjsWOR1RnxDx7M
TC4DeddS87rN0PG1zNkRJKFGqejyf5YeYLsXDb1s2RoqLYlmwXtkA64rytjt
Q6WIjMkF+eMyKBo9MFfqxS91CNnUjek8YXiRY2st7yapVAoK7kOqGxY7lO7V
5CZotOUCo5BnXKi/9lyn1RfajwvnMyLc+vI6eXpOcyCzljn9zua1xTAp8uTj
+BNcsXIj0dEYRqpUB/nL+tgWCGBhDvuX76ymsoCrR7OuOfdzjpa5cq60KpW7
/OnVNiXVFZ4vW+lRwEjJkoq9u81MA76kJ07TCfu2U33K8u9QRTUffZwduRCJ
UUJw5WL/9wJAFGeYAopJVzy2ZCK3MmSYd4l2F+NeFNv3wvB+yds750wKu1CN
JwpccLmf6pyb07eyIdp/nfpynRkUYU0Cb9eoQX/DVza9MHtNqQXChy27RBp8
1eBVCi0Rf1SNTETmSWNr710+sy9D32xSxiSVI4WFk/Wnw4VfqoN62JxZNno+
rQL3f/lLTF3DnWVlp5euiOqi3s7wmMHB7fFfnVRv+E49vjuhTMi1t5/V6tKr
mqr21dELMmCkz1HTyAXK7u1TnMt/l0msTM0eYagBiIKn1epQU6GS23pmGQF3
Rfe7Tv2aC6EzNv7CUYyFps8eyzSk7ZE/F6hHmXxrdbD/pU0YOYtP9BJMrZ/q
eA5Z1GTLzCv519p3p6WC2jqJBG58XxVxmbkUg/CQkA/fqxU/qBM+B4rVRFui
CKexLrKiyc07m1HaXBQgKd04otc5seZ7VwcDtT/YCxoWO6HG6jkfjt4zShKP
z7mnwsLpCKo+05S1Xhs6DFzOrMAscXuQE3lEJWP4IAtHN8ydkfbHuk3bsCjv
yilLHlaP/NimSIShDYx4VmyZJYaqwp+tobYwMogCLQCFgBX5tASivjKGvh1f
s0EiYrh7VDd8OCwciYd5YE9FvlTQUquvbqIXND5N+eS1n5nsiclB9MJYjx50
I4Fs9FKUNpdSnEd/VEi+/ijUUhW7zfZCVeiZJZbC8C5zLN1cSsqc8GfWLbuE
8JdnFaYIZQdqeypAJDw1TV0l5mFjxAOWF+AsfO8X9JCXjcHP1+5rAKpRT2zy
d6bNu/ohVpRuiIUbHq+wPQlz5NLc23r4wcSwWnMIytv7IpRdoIfICTselYRh
HBYFB2Cn3YXWyLv9OHLsOEwohzGlFfZQd9e3X1tTKn+WP426p4CwVAJ8Yo/c
VT4f6KajzSJH9TZbYTGV264qaFx0xqUd1ExEt0i0W2gHWlPIApApDWNQh6zr
PYDC9pu6crXxWb/y7d4bm6UHJjzEbNCx5XLA+o5iW9BKtBH/v6CbaDgenMy5
0rTxMMFbIpELwJ2WhPLRVihlhqatDrcaiugQ+lpMXf2YfwCAxMB1mUBCFIO6
85x1KSM07CxBUfkPK8ZbVbNGVnPJhpzKz0Q8nox8Xmiu/DO0I+/5fYSimqcf
TeMXZWLfMQX6j8KXvLWXxJxCSbkTEh7EdipTAzGumdmdgerfCuarIP+GR9FV
c7Hr3UeRgYO0rHYw5g6R6diV/THSErVUNYKNbsOW+MVqqIn2iX+NogRLSVyB
w+OIAaC46FTZlyuTasZjEIWr1nHMjtsLoxkDDqYGmhhG5pxbFVFVeaNfvZDO
a1WGrG50MB194imEWbPTk+QrrebjpTYwM9ZPLJy39xLox7+YHS8/hQC6FoL3
nzXq6/NxnUVs/UbACTuDMepEQf1z5TkXqfkOv2WePP3tAarDfuufrWyRBjIm
naXd5Hrr09nf4HXpH92KkOCu9UvPZ3ifL1bul7jxuezmbfYW4DVWYCjqeiun
u93V24E4ZaWlgNy/ayH8fExmSvo6EH/B89Ay3ODdSRpUuv5vGl1vWRERcema
ktFi8Y9PcJ7EI6B6F42zGeJsKmF2FMbIFM1DBAv+LGGr2HemOf/ZCtInUj+3
3ilcV+MzrAhQsU5dgLV/mhdFc756UBpi/0SRjytX9Hx8s9ah0odI0ATRAnPq
HBuAItecCCSexDY/0Q8sjNr7DlpP3qGjNnY30DXlPuLl7V5q+qeuVvwzNmVy
XEEzaBl6rZarKafTPlflRDUi38NZ9wqvW1tVteYFTpsVHPBxNfY6aQyRkuzI
TT8kAP3nVszRUmttdgJUubL0YqCas+LW5s0IJMAjCMQdklb8IXeO3JbIkhPK
CrQBk559qfkOEin/LDKT6elgQEYLVCEB9cvzRyoZPF6UDkJuIfJOw+44Dpp2
doVJqSyaQxEleF9qkdw7jqcT0/4jtQ9zR+1Hr8LSj8EKnpeZ91baFowDlpiI
c9q3gCJLpASO666ZFRVmDJo4Jd+QzutWFPFJMC+fk35jvt/l3ZL6SjigckO+
e//qkyDNIACJYAI3zLFlBM5CoFV6P6e5bWj/oMqRWYx9lIu+7Fof/bl/sSCd
4FQEZf98IXiPmFHuKTbwtgrLrtt9KzYP5PKv7oTWCAR9qfmcnTnn/6PtC/hn
6P+Cr9hvWMMU+Be8p9Bwi93npW3q0WwbD+iC3vOr5kWxKh2bTqAzmX45eVtJ
dQX731M2yKcrUBKNo+p6que2RXGRMtDse0OkBfyM1gaAXgz5A2NoqHM1AggR
9xogsuWGpCOtsF7GCg8ADKk7sTBkOFgAOXKrv36rCRQurJgRBziOmDhCMAyh
coNGVSOt8TROvSwJJQgAEJzmA5kQH2p6nkYW+QtbkDW1z7g7Jj1q67rF+CzU
vP4JR8wYcMePCJqnAiAiZwrnjemM2NWGN7M2EupOHGuanTQUcs4Jk0WBYiRw
WuJnC9e9aSaQwPZaZD7RKhlvF+LwMwOoikhcLH4JXN6vxbwYlxNeqZpe6N33
GtIPolhK/QiZw38GosqC0+60LqZbAtNc4tynZHfFq1HdT92fZPJMk2bHS6Ad
6MzKySeDrqO9Ell9lIloa9uRrq1KbnNlE+YryTWNoaob38wewg1cUKw6UdCl
l0KrWH5jGrLnZ9JMXjyDU9iRj4t3TbPChrtvSq7id25PsjJRM03VKvXD9iQK
cXJxz7P8MtFqxcsm/X60Gi09O5whJe0c+YqBfz7Qn+ejTyttmxb+vbzQo6ke
gJTgFNsZS89MoM/1AGIwDs+CL3qdy3TCjnd9OawYl61L+OU4flKzJMS7lor5
u4AikE9s6B5PUMPWPpqMBifbK1M9NdUiJkfTXwXDRwM+SVtouP8yOH85lurh
izwKwPkxQN/moWBexE0CmR4BnRLeIBVO4+RxSh8D9XiVaeWPkT4/Q/7SaEvL
SOxKN5K7PJXHKjmf+cOk7PVtnPBPvDMLCkaF4JgRmkLJHjI3K3mXrRpMlTAf
xwxvad0PfhxtoxEK7rQpkIVgeI9aUKF9a7dMhY4dT5HQVIEXpMf3ZwvhTdcb
lNzug8Sfdusp7imnrk+VZ+8G4BF8Vbblij7vrJ0P76ZXBU2Bz1/YDvvHFP0r
9E5xmTHShKTaArN6CCBC83VzRo0LTbq/RZbN9xCy4VJjMXKUhATRZXWIIlhH
M740/WbwzznHlzz5aIvDgoLGiDgQRHIVNLSlNcvQoSIdyc+OQ1pHC6Y81vix
MLlwCyMESu0HEqzK+0OYBtstkEd8FE2eloMUVtHLqUVgWkfvCDvOpVe5d7mV
RkgJxFW3XNSyzfloFQeWFS9tbpkuUrF80jgKJcp0LGsLjMzqfrnnKE6Hl+Zl
o4o5fjEV0dJ5Oen8Yg7WlO0rl/oT8CXOehHf9r9Rs8XJ7rJNUHUY94JiCZNH
6ogKbfxktGHUFn+iyApYlkTr2v2r1HFFWWY02eLkzw8/7XjSTqB2miJfZFcH
Rl31VmXUxAWM2ThYZl2XVz5khcbXzR0Smx3qughd8MhJOJl+dw6dC37VlErg
SODLOUbP8oc44kpS8uCjt9lRlTQ6z5wTYoRYl6ahLZNwd/SXMoydaJMAWGcC
qxSvImrW+Y+U/RfUfS+nJ7A2ObgKCHhtbi6NxFJvGn/LkZ9kf4jec5EWxUqG
viBNNtQ2Oeb8EhtiCyG4huRtJMLe/zxocUIcUpTI4LPq6Hd6htOsRpU7Wu0u
TJETvKZ9fwtItPAXkM3lC0k8Al3+QmeaUNsQAIFWoNe1FofLTII+hg+dGNlB
V5hRaHQ94hVKp3Y65AKBB+va6ZS3pH85/QFjWI/FXVHIPOYjkYjMk1TFPjYJ
BeLK494ISQlK6yOznWmtuA6lX0hU5FW1KlWAM9bdAq81Cu1jdiYBTTND65Sw
Bb8H8TaYatLgx79hm/T+EJAEDOgf6jivQRPCtJ8FOHgwGp+R78ZN8tUT/CA0
w26yyjSy6q3DY/Udvz11nlpwiXGG2xkoAT/UaHSmmuKp2LkAJTI9qRlOfWsU
UzEqo51uZeBvjepWf6ezSTi4oQ9pHar4ZZdCM7GQpp3g75qM1aX9fvVOVY1+
YRQ45EKrQzMyMGn5ubyll7KqQZkXisoB+MIdTMhoU7mAXGPNHm8LIoNm0fmA
HcUbvwFsbTW5ZO2J53YlaZmcJOO7EcRGea2KBzumQS0JLXt22xy/1NRupemq
Tptj9QcDycuxFa4t/xdDSs8Rb1wyJfvCbyenlaUC5Mojf8Gd8mfwvgJD8wLE
/nqFNQOyWHUTCe2SbtRW3/5hD+ds9OVd6Wgypn8sPgV0wbv5zyfZNQxx3qxz
OgymTUyMD0oc7aurJUzzFI1bIDvlUHDNX+3qK2ti1E/baZnJQgLVgMRpkqk5
xPm3jxiC404brS8B8vcEczPvBWILh74LsZPWGrLxDrkB/6sjuQvECyPFCut8
qdDppBFt7OmBOgEWj1WVZvPB2AQswJbUrT25bmklRa2MEmc3/wYOktai+bzg
S9AFpixLctZY9SwoLrcXWseKWIIr0wb8kdJeRcsIfoDnNFOuLEUvvwAqzb3r
gT/S7VcAQFhcKxFNIT/H/8WYq7hIduWiFan6WW2FXKto6ARdnQPzlGXSgk13
Wdewe8Q8tmz7w1ynh9neac3JACONIcpnnya7cmGP7kCVgEV8Gt26uxYEJwgE
429HliZEKtJESSaOge93FF8pUfCyTjv8cwyX7CcZZDiH7pxmXHMLPwRorBne
HXkdaCuV1A3whhAQfK7dXw9Kf+TEP8L+PyJm9Ax+RfFh9FeksEOyTtf5bjtp
a3JkaoSiJLwQgIF5347ynHa/eXnM9DV318lGmdTT48cb26BBhyeDq5cs6qFR
SLErUJkECgutVfVlteb9LPx80vpKUQ3Lg/Mo+fAOi1arV0HZ5VboRdi9NBdr
4JGNpxxuNLrIiskpNAfvmLDGOerwpWEHY/a2s4P+Dz42jaHGtvjCNkMY8FcV
K269Kb4P7gKYigmgTV9zkPfxwIn/ajhZdPrZrnbTZm9TxM2EZkS1e+TibtwW
iijk+wRo/5FrYUryO+ZQbSW/UtHX+CY25LADE6HJJTdaUE3PUAPwAvaRcn70
qlkyPHilkT4QFVSgMfwnYNTvn5PzRU8gxEIsCv7e1mzI3ZFeHEOXHlY1mNb9
CdhFgvblpsTSWDWTQx8p9aXa2GLsvPaj0tQWX/tD9yNfszZ1jt3gtQN6Ekq2
bUgrzNJB/0yib+gCsoUHFpWYtQMp6/ysCrw0h7mqsqoVWFe4pDI/TNl6u0sd
iMXqNpJcHQLDNeceRSfX+R2wOBAKS8mAh8IE8Ki+D2Ixz3Ft/iw/Btc1vle+
07UXx8BqjopMCSS46yonm/yybcCURR99dROvo9JwYBMwt+/htQrrIYxzvVef
qTeqajNTvR96FG7CFEKNbF6C29AsQClRjd26z5kbmztGSccbMerMXU7Yjbq/
X5sU2aSimMua9vTWI0ws0A5RtsUhp+pUZakecHpePlq7rU3FNWcTRCyOjsxM
itqSE+0eWTwfIoA/ryxpJgpt7owaRBnKpMMIgUuDW4OLNfpmve6X0BSSYEN6
wqm6q554wfAHQ6uWMhyNcXV17DvsGRGfyH6hs5SonBGjPW2DCT4wLhlPsvjK
/WQ0QGS0LxnmPMbcbGUX18yqCdD4Pk8xFLt/edxIS6bLe/NawId4lJMpmsOC
wK4ZV9XIXAjyTA4hWppCPUSSjkuKPtMtvfpSqMigLUqAfBtF+5A72VH3iZmG
HslJiAx+kDfi1dPb7w1FNMtBB5YuFOBxAEQJl2Zzi8loIVImF09COzco19EA
nT1qppheioAgfpm68WG/i7v2iH+eA257xCAXJHsAxlmWr4L5uF9pRCLR86hr
GAAFHMHvuwssfcpuPkBTPmheMRhgDHaXnKMAogsVv5hzQL1ybaNHQ56Xwii9
vBZt/pfAO2sSyDNKRuy9KrrA575wces/M7OwcS4BD5S/xn/i2PNAv2r1JIrx
KVkwDBueON40Pu32Jg58wyPYgQKkqLBQ3zQ4O/WJPYGt6cY9eAw/hNqZgwYM
KCvZsntCnGmtfcUTtkvFCY9mUxibo3GhMIB/jqF9CTG2lqPdvgimM2OCd7/J
dgEgmqAfBrY5i1ZDCW4dZ+R+Hv8MOqM9n1Pz7c7LLl0AuW6+6YHFhc6sT98A
JNXpXzzdhM7xp8QXwI9JH7XYxHb8L/uRR8CxlDZnAqE5rYCVtfbHfNZvmbV2
+ZYWkQu+7KzCissZr8tL5Ch5WMUBaOb3ONRa1Kqm00vPU/6rYPTwjPmkb959
ZjswRo6VKo//7wlxPVaDhGsQvr0bS9Hu2jB24h6WN226unZE2t0ixh9a4Qws
rZFrYE1NpI/YGhT3x5vVNDQkESh1sFQKjN32T3qRr1Kr6hpG6EEKbDie1zXN
ZGq/gBqKu8EkbdPCDCqMz/DjoAS9GmdibexgoJlp4XdvJHtG4b16z8scp/lS
UkH6wPAtjGZzcFZ6ORGgceTDeXrxezjsh4bHj/cwLVG7vNmzsZ64nLA05lyh
x+Msrcox5dQah6k/fHfnhZCMYJxphw3dyqAL7Wq9+nu3r/FGQncZmD4R4CSp
e5rMsp4EmsUKWBHGRBRDczKxfDtrtnfEYDeO8z6l+FGLS2IvfDYceZcyl7TY
RfJHGj86K5WPbrJy2cbE3N1bssInBpQ+2t77zsn9AStzRm/MbTe4GHK/fb/6
CBvicpS6j05OiubnQnkUfEDJug8CYQYNVZMkVaK9kkJOJ+ryeijsGWCMaDBx
87P5M9oaSU+JbqtUNajah2xTFX7Sody1zLYYLuLTF46r8Kp1Fo4lE6tXYeFY
LXTsdjgTtPGVqWW4IspM2Z10+rJWnQhxy6gktnMC0fTYdVOWP+bRl+uKMF2q
2nqbXPA1B9n4ZLi99bzcO8+EsSJnYislAe8vyFbenQ9M1bKVPWLT6HVvGh2K
DrErZ5s1MEcjxG/iaZRFEBU0LTzgvqbH1OrnrPm9XV03uMM4HMLtey80ZsPr
l5HIf1RiSQftrO+JKSzYRmsDedUhHwLW8cnaUinE7LkD1tiP/CJK08O02uwe
SZEiKneBxCbsosulum2e2HS0X4ug9s8eaL7FDrWO8tXGGQeOViaQK2akeBAl
uzckq6D21AmlkdQTUPkBP798qYoKSzu/5kggg43qE8AOBFzZshZpbIqdIZtS
oo1v/+zZk9ecaV3AlV8RsCXmrrSCy/J54UKRR/LhNZXIkNo9hfhBaL1xqwa4
ngsZZrXiAB1RyhCCuzYyRkBjXoKtJnFtioADITO55FriGbQ7mv7BfMEY2s7y
3JGmxdUGYKeFSt6s8olN2qgLAdILgNGvfbYSeh2VRWISMEGH0axFFuVLsiG4
ViH55jKCseCPFuDTT8TbhyQiRMlMeHjkLz9hBdoi/mO50zsPAiU5WitgTmZT
KUTgy1H4v66v/GCkBK30AlIS0+p44ZWPvMyZTNxLMfzHqxLtqQ2LpeYmYG9m
a0zz+3nd7vSN+yGZCNKBJzuNyOcuz/jXebj99dyviQBqBN3mkUPG3Itrbv1o
L8jCdcoOfNfuUW1wo93GcF2roakUMhV2xGgRWQcxOqRYDB0jy6q4qxjAaLuE
1zW7+JL0NtQcVPNYuApEWN+JqPYU6tnDca0L4cMZ2R3N1V1NqY9EBA2IZwtq
b7xadBBvOa6rp+wAU+IoENAksk+K7PIHLR+NVHgF6ap1SBFde3ysSklSstJ1
3WOT0FWANvqA1hVBw+y+dDsCcxunuhCTa7F/JHLJZLYzOgHIPwYTwIeOgG9p
0rFXCJseFEDK7MZ3t71sv9RFKQ9q83zeVPeeYQXI0yNdkctqlBrlqXROiLGa
/ntrjNwYXpK6IesjCbKeGy0rHIdn8AQzaJMQ5sUaxh34fPR2/HJnAjtGBhEW
cMNZRLJ1zPApcKbiL/1fVVrTb3YY/ahQT9BDqyF7bwDW7PpoVklgw60VYDEs
/Z3VWDioGMlsFPjZJzdhzlqaJ9xl7quQuQJ0So23lRxS4bwIrEM+icmTi14n
0ld4Uq8AqoJEY+vfufsx3wImwuVi7K+3gYxAzebRwY149okc6kbb9Y3JQhT6
qaixs6aIFLMZATdbwigCX4sc9oFQuuJcqTwdhd1pQ6LS/DVS8AutIVoRpjhx
gCpQNCbaQQuhhAm08tk3UKa3DQYknVtNBLqacXodJi9D5i2Bb20jQrJP7yk0
AZgVqvM/EYhC+UfJqQ9hmRCvr3HQjngt3oVBYRU7vreAkTeRRgvaGY5vH1t4
RmFPe3nWxriaUFOuc/hYxsMb/uMcSyeSaUbxfXuUjF/haGxo56lRNBdqlWOL
CMXsZ75op/Z6awAkQ2gNfKMwqx2Mg1inW76oezGDVfkSxXbwD9AkRG8gLTXr
yHzal/Z/ALDLkOlx7MstJ7ytDQQqVpK3/A7rzYQ6UeCA9C80P9LqB2fcHo0U
fy4vhLCzhDw9ofhH1ezWpSmqB0L8imek/8lc6bHmb5hDjnj4y52WfxIOcyvG
to9B8XkCOI0ty6ieIRD1TaGU1J1laq/pw6+0d3UgjG5yyKlDfgnRx8Kv5YNf
/yjP6euganaI3QGbjX/mSfw2KKoLCNGuLAre/x+3O/2UAN7WPHAfoFJkcY2F
cIFn/EPNMopdckK7DrmCl8BN/M1s4Iqn2Qmd/BJCztZ05XfnICcormBRwTG3
G6BTlf4OJleiBdFGs9jaOy0B7hVPcHJ/oJ0ynsPAbT3UVZ0p7Jme+e01bhd+
L0yNPMhPEhjP/GGdvKYUkAG2ag1L9eNb8kNt5EEt3kmPsPMb3xmOSXFtN24m
WG69RX6T7nfdYwTR049uQqSp0athg+TjSFpz2JX/Hhiu4yphLEy3km6Fs+aT
O9BOcuRDZABhrDfWRq1LddURL7UAGaFqDL/UppEHkOt8wTubMcMTC441Eguw
1UO9BLZgJFIYu08WMl2PZUD6HLZFL02rSS/EDirwlDkdyJaYDZiKkngzGmdK
LZIH7wCzKGVU94SKQOzoext95HqiWXgwMEuYnxrS78o7Q13fCphBJFGjwl8r
c4BOS87W7WBF8ptBX1251KoojuU2Txvu7xcOZXhb/C3fxCNQnLps8Se/y/ml
8D27Kq/RRaAocv3hLKO418ho3Z8N0IOLDjWjM4cnj2gReHMsk1JIVrc1/kKW
3q4QOG7FQsGLI0HAzPYCkylU/aek763h4WttCHmWpleXhn16mFCuhJmKX/d3
kmYArzdoZdUVb59w2dv6WlsHwbaK67nVesn1694XVb/S5a7yRafXNWl0md/a
Dfep2A089MCP83BzFQEhQcZFUQkotABY7Gx7THIdD+66eNqNu+RF7XrC7ZL7
trakw5YCZAqGGldZ83myIV+kBfnSMizUGYPlAq3SewCYKmHb+YjdOI3c5Q+f
CoWUFlTXZwx0ztBa5/pyOg05aLJwYmY+xQCSwpn2NLxLVCWcHjJ/zZ1KEHyL
jLv7X9Z/9Jie3EoR+bqKPStc73P/ePeXwUhMiJxSG0X8rpVk9ZFqO2/ovrod
ZbGgga5z0zG88dzPEbxVvdmix+JqabjqanKd0n8Y7nKGuQUg7eyGg1hM6v7M
h5bCwYbHGUuSVw5yP4M9UXmMGl9EaUSc12P9trqy2F0U+PdxZcVjJDXt863z
GOKK00cKLY3GCr4RGybVpPQ6upXwmozG0IRuy1ejIX2bfOq4TL/8oXyf1qSJ
biz8tPUXa37517gZu0lECWFk4gj6kNjVizfnMaNOvB7x1+5y1aiGuriuV+yE
PgiBN3t9vt8e44zcZE8jRtkfs95eL6ejaG3D88Wt/v8bpirmJtz9+WolDI12
UWdj6qpZK2MeSNOGYrBLtUqLfIii3OcqXHpqF1zJeC1cmOxssHv431LGyiOe
gggb6TSqd1W42eopsFN4ORUR7Bigaxt18ewUOtDPC/SoHZVPbsjGlAln6Q1N
AghoLAs2Kp9tXOuubWvuvE5Q4yEjvUZGrg1gbjqb+xXN6/vlUhS2o+431MJV
2/+zQZUeENzKu3/UeeByrHbcnfYRIN2uexH7VnWuw69iyh2Qq7YLE7RNg2R/
q8DknSbv8I/gooNdKIzj1VOyZjh3Tfz+MtzxxW17Ip7JAG2kOpd8j4qdRJGT
19LuzGZ6hwMU9PENel0HLVPOzfCU5R3HammvfHm7eXWaNwCz3f+GXqZqJvq1
MuY/zpOLcNLKZffjYZNmgVuK2U2jHwgcYwYIcJiYoqW+V1dT4xdnQbJ0EFyf
QkKSbK72vAVxg67Xv2zwk88G2DAUpmmysngP61UUsyYo8IjkKx29htQI168b
8AUuy8n3dt3745KnjrYdwvu2EZbpbs1OSeHNC5qwfgY0dkAc/elos+hzhlAH
GdHS9tSuZj7RDy1PUKkrSr1KhyNXTUejWETcSBb6OTn7HLXTfZb3Cm5VsDF1
mpeI3WsHnRmWsUADIGDJRVk/k26J4Jupimu5FDshmVMsFSTxmoC7iwXgJ9HA
euKbo7JkLgVratSVGK0dQJ52sNxJdF1oM3JliLtnRhYr+kVSjZUlUAjpLrRL
CCihcAPkebaowumht4m9FgTFW0n9E0XnrRN5uvgxJwwq6QIv+eHWoGZOuiam
n5jwrPok9xDThsWaCar2K7gEr2j4XAZ0CVsFXFATzMMOaOnmhzCwtxsqDWsG
5EdFO7s1/OMqWyKw0MrSZDIasY4wL7KmgI7lzV0tOg4lkMMP2+qHvefF+cMP
CFFANh8L9y32C0+pxgTY9UpLRBueSM5tjjdJk2+omSIqyIu3Iy2AcbrNv+9r
rbSNk/zCFoHkHvM4kY5pLN30S6DaZlcNo/BNchqlfZD+tEv3gyr94hVYJ4O2
RAs9junsa/umkC7tTUzugloW7PiX7p3/0ilUTk4OPkpAA6W7CwCm5B5rtKTL
iIB1BDhmMW7gS3tIccD3FOApBgke7zOPjnpBY3t0ArPXU01wAApknspU0C6e
Cl0mRTCEwVJwY+ykoXNwOzGogVDSLKmkjFrbxJCMi0OMqbPvUkCo73rlV7z2
y4U014sINcDxAEyqQizxFcMxgR4dV/42zldn3W6WFQeuIoguRCq2xV38hLbj
ZXeYahYnRQarxwgNdC32EL6CB872vVwva9fcjyI7tFHLuL+VfhMS3qEOKLKq
JRSt1/UntrHtJ/l9/yMrBXHj6xE+fUtV1LS+W8ZZpa1pecJ4FpK40Gjq/biV
7Dkd1PCUDLRj4xcrrvbad8RB+ZznStS571U8CrqmdvcZsaO1ucH06+n0szhh
qslXQOIa+MEvfOqxB8/IXM3pv4SanOyZEe71vWNVc46Qp5vC79W2XPG40C6+
o2xZzpklCTI0lgHlfQ4B9MUBT40vjkj71QmD8p/XViH7xNiuYaX298JMzdOj
hSJ32QZHQCZf7PLhaly3MVYsQfPU/sxs8T+Z2l4EqRRkvFa3VrAug1FP51zc
U2aqc6YW+iy+CjswuK9H4QKGkpcWG0g3TBZRW7DmqS56O5szUZUSbyi3q+qY
YS+1uc3vrLHfxujDuL749wNFRjQxkYCT87780LsAhKW5IpIPAEQtfSuf51rB
a75oYT6Ap5vWlCFRcX5DugjIUWJk32oKf1Q4rflg997j61Ttp7rL1RAI2D0V
Z2ufxWlbC21HvBNz8x20kn4N7Fsqdi+eet7oiKPgOsHrV3vC6HRq8sBgiFUc
Gih9VaoActFCNXXfnaJABTUeoGA4umF3lX1qFp8ShJuPs7j4+Hlp9KMdyEtN
Q8WN4lzn+2c6YLnNnD2BzgqDBJMXjs7vP6uwZU22/VJpFrV2j2mqEYN3xpEc
Nvy0kVowXv1wZVNOB7c1Aq99HSxDoXLlEDQL8gHusTTJYMjyA5+fAn26eGBS
NJPNljxXaWZZfBErNhSSbHeU4HN/O3CwHHGUtNc648d+C3fvI1qWXzshsp82
UUnKqXJtb/pZcHC1LcVhui2v6mCEAyBRsM3U5/+U+D0JE+O9IqWt2arQI2GH
LSzwyg2676/TYjztoCoh/lUgedXnxKiuNKuVYAtOzmxUCFIP2SE3Xw0UutXn
BPq9hMihbmVt9WhJcrP3cuQPQ1QZrfGxkoxNMFJaeFxPiLFwMjaaaXj0dVBc
VDEWaimLY/urEMWZshznUPWk/SIcMI7hJ84f+C7g0pas5cuky2hsp9n3gAFn
bDWcMgPWEWME+anfxAfw9l5doX2YxxnUGxjGOdrzuPcZNXgMoN6eu36f/Lst
7lmIThtHcY3oxwssT9xdBcHvT137RbNgi4Dre+xoDIVKYevvQU0KBk9wC5Um
vZZt3/NtOGLEcKr2EmvvprXW9mBzhweI6bpirlbAfT3Zf+3Lzl/PyxugxO5M
SchTcI5f3pOZr/2LbysZeU3rLXV2E0MzZB0+wul5P1Ws2z2PTrVoiXMB6pja
13PvYorUC5glZw8qfLfWagrpsmiAif1fHXLq0qfE96kbR0qDJ4BVLM0Z8wNX
u+Jj0GDuTe0+9QWjq+tGontSowPrwY7kEhmbTuMIfsXDYe4mra9sfP1szm13
FctwKm87AoHRigvGKiLtT+UeyWI8WVHuqV00K5rCMUFvC+MyuLxwSeLIFyRM
QNZoP56aiFLvH6FleidWc2AahM+YW/+Iplszmgf4gMWcsMT7v22Cw9tK+S0Z
4Id12feuaqG04ubdHdsKRDff/jV+qHKjzMnf0kLZimmW5buFhOIKCW/KvOob
+842dxepWsCIumJfW4XVLz0xeeNDa9e1nZh0SJ2rjyNMo+5AsZj4UMENSGYe
QjmAk2XO10PaNY9JX919zYUHB/yL6kWpdZb287YM9LboopQ6NJx0n34cTB7E
OCse08VyYbdUUZmX/BM426jFwd8mgVkPsnHaea9XgWSiQOldPZK3CtRey6MV
BIxc6wbxqqOVgqc5M7zsioM2z393vCNQE0KXa1bhXc0uODGa7vIHhEE1A95u
BDh3XSWKIaDr0NH+sI63eUAN6PT+W5YBvB9ShfaEyseERlXc4/C3M+XQOJDr
kdoKiWRdR2vSbNFI26jKtTCve0AuV2MsI1kMa8UQolVJayPfK35p6NVfBS98
BUsWq9eqsrtTZxYcC3FWdX9wmc/LP8oHSIgx3kVgXIGzBSImKiGsX2Zk3A9k
0CfcRJQAqjGxPG0Ww6Q1xOlo8hQx2MV6GYVtSDSrzcojm4NY+iLPkgRmnpoo
u4eT6QvKqHXGffgtFGSs/UZ6c/VBqMTQjeLFBL357UnNrqjbbdP+P5dVoa/f
wVl4ujEi7tHsanuT4V+MHdwVLRaghSb+IYkKvDjt6Q8hnU6VjghzsU1d6Ti3
MwVavaB7wuhyAuHkEf1gIls7nZKCcA2VsRhBEcZwwbGEhwousd+1xxkAuDra
/uVams75fr9ymu9rES/0m9jEeeRRLJJDCdaV7kzFLFnq+BVE6ZEG+/zay5Vz
XQI0vPsL56qpuDHek1p/jleLRGUjjmJXJAZ9Smmu1nnQhnntrKrafKIfy1qb
LirwQsFgRfiEprpp7hpmPq2+E9qacXME182JGdU9uhzVP2+TNPFPRRHtZj4d
OtvwyHUFv0SWSm+TU45sZ0xlpw3q7DSCg4UgN+VgrJplcFcZxr3Syuq5HTb+
O2MICGb0NBCovpiZQZy9JjUMVOUUgf4k10PzR6zLKzsE0vAW3PKGxThR0yPj
Z/FCImeVTBr75xMLUnSw69ZVRO6duE2MjRWbQlFVF2O3DsyDqHfYirJYQ1EF
21Qrzy9uiVubix/DHYY1gXxyDpiGCbXr1QDV4G3qCkxs1RWF82A1LcHLjCDJ
I16hB0mnCFnQkiYDo63x0KB+BKmdnpFGrH+bLKvFvzj0vlEErpWfB73fsU4G
Fn38YIAEarp/mJ0jCli1Bsvy/PmJoPlcPESkJtooswo+fLr867N4MHlDPdTZ
7P9VIWxHhe3P/Ta9eN9mw+wiqYRrFo/SOEBTaIjGDSj9pZCN7TFFEf+/FfRy
HEtvI3htb/v+xxPxHqg7iIM0oq7YRKqmPAx/Em7/oRC8c+bRlHTzURtpPxBA
1IN2M32+8GNy5JJsvKqMReyY5MOG023Z7LfB2fHziXkpQgIt6NK9jicYneIO
VMvGvfQMbZttZO5GTNWoAJXrSKMUgxNQja8TvVRCVdnL1BstTdD44q1iKYS7
2F1Vzn0DQ3lezhARCR3sp3Mp89GjETSuQPCuoaITckxEDZVsYT7ThTflHcKK
UUCZCUHSQz7HP+J4ubm+eWUfnJLJvRi9ua0uxmOOUCNNIBBr6SxWwwVA/iWR
kVnr3TvfPJkR7106RVWyrQn3ctGe4MBpMpu1ifC/XKlWQIh3IzYFbIKrh80B
4VBFS76jS2hJGhimhodx2uUhzdoaKLfXnayCfJglTzLmb8nZIhM0ZpmJFn69
9hmKWbzfWu+FCD69iEEF10nwNBAT1C194mncMYCutyt2ZkVaYiyP9Ft+fKfA
4lfActD/PiWYWFS0Pw86cAVK2SR6OVVuv1LeiIWAoIox8HKFvGxa22Z4La8D
gPDMVHLmqOdppdMh2mcFoUY3H9OtEGQ75kCF2gFoP11EYXzjGjEK12pzadbA
xsomVxQXa25Lqu8XR+U5zBHdIgzz7NtuVPn9hgHG+nf6tWN/b/idk6CJSTS/
S6tLH1wqljPpNveoyM+YN8BM5TCFwBWsg4JTXjdtT5+pM6lt2DVWi1JYgWbu
p/oL4/P9CaeFl56aJ98OIYbyRjxNyQsxrjW9LQJjN1d0xLjhLV+Vo6E1mei6
2u6AQvgKkt05JyHLh5ERlc8QSi2tPnZutUrZFXFqgUaI4dvBlRnoYbq+VUw3
Gtf2rz79+8Sn+bMS9FxYzzV8fFEhWHH83zPSVjGPQGUTohCh4fHmHEitA2NB
Y1tCz/VoKsk/fS7jmSai7s7c3X/zWy/msLApfTLWrrxAtpCvi9TVi4GV9Lmy
YOMYT9Evx7B4nVZVB4hQqxWWbcDeYPHvZ1dA+iMgEsYkumYOnoOtwBShm6ZM
TTM9mvR1inE94jK7dVFRiXDwMhsGOSHiJzwY66N+F7trbFqMXZ1SANJedLft
W9rnBySmks2iUobAFjb2gwR+mfBKSpzyM/OME4gpxlaaSC7aNG7XJcniXlpr
NnQENcKqR0/g6dL9UpBCThaMeOnOaRVeoZYYLNZrXqeL6jQRpBXsUF4e/WCe
Sc5aXKOazn3rkZvmGsB8EO4m8J1iiOn9j+cK1xPIGRv1HngHEl3dVz2cb9Yb
aeWVMPRvb66vih2eCMnEzuBDamJeCWL6Qp7ruDDHa05C2Nc5smvDAmBLN7YL
M2X9UeBG5nx65V8p07La6F9KZujdJH9ibGTrIr00rs6KANe02Hvp8FhreRZm
nGj46d5ub/Ko6WCzTYkVliByv5f15l/cuXFmLuLPkzXgnmo47A+4bmoeZeHM
TbzFjji3ONzsok7QolMi1PZCZuiLIbPz/4itYqIcG9GM2rXycXgPaS4Vqy0C
dy/qBQH7kEH9LuIUArPluEMnRRomcbCxDhLISGuKTvGC4m/BBjy2aE6b/H1n
I1bRUzSq/d+m0w4v9BeTLmB3cyUmy8ZBzqIRRvA4ofEBUuo4DZNbyvtC7jVB
vkGAO3RDdnz2565wIkUslRxGANQYB17MhpmLbA6U4NwJyhQb3fYoC8hVXBZe
V7bR7ZIfHZZzxdaRQ2IrIeGjqwILWSAJPCKZQeAXYUydf3foaQic5GTMFvUf
hXTYOfnvKwMilAG3mEwUC7eMLmUpEeb3r4e5yfakyYxovka9JE/tsNaw6uFE
J4jnvBw83kb1H9mOh07tZ3dtlisIP/jJJdJ2W5nd6AZFZrPmVz+04cEWxMPB
jTI7a50oFuDq29BtcTiwfF8ZxIAlyqs/U5pTT0Ae+XHpKfNGQAjOCJ0V/pLW
+9bxkqx8f/PwzJoWoXKbW8NDtMJHMPfUN3STW/l6Buf/HOAOjRJus+n10UBS
Zf5z9Kv2usNvPAnEiMqKUdnRAaJHA+ropwFH/7LFpsXoGxeYlkJhGh5iuezG
KnMo4LIZ/iRgtocyCnOzl6pt3bmXAm1aw2IajjSG7fE00QuNJZHHi9v2vxzf
vHtGQJSQOeOX+9hqULSFPimUXb5SUVrX9/SggaCYZWUE3w9EClFWjwyMZk+g
buFjFqm4DSyPjT0ImssOlnAnryXEhLB7EZQOQlorfKfsHrYpQbWsZrA2/IT7
YHz2jaE552O4qKk2CV9UwfCvoPxuTO2WFkr9ErwBhdI2Ci7NT9IYuVLoey4n
pigZc/FiEuiLbfwRW4+XqHZNn1bgi4YBQ9SDq5svJ7FasIirvwO6Wy5jBw2s
drTmqg5jOZCAEf8hehasEYigFJDpNMFQZR6ASBi7jTqgSxdMMvfnpCUdlmF0
VrsYrr9x1ORDs3nQr5tmXBaqqeYupjxuedJQS8G47HnVGTPZsIBZpcVxwmyQ
ZglFdcJDbN/MQXzOgFo0mpgGsHhBAxsHe41Lzu97VNOkoh3GmocYGubHFcmH
sIdFl6GmW2Bh1xxriaprt8nix3EoVFV7rNn/Ah317jmDwPUeUh5d1qXq8KKU
1nrHB2w81D0OxRn3rtUXugVZGNvdpCDXLK53MgUqUufxw+uN7da99hw7JgpI
m+OXIk2dA3KO5LzLvZBvWv5dE5zv33tS7Z+EUdObOCnAXmAJ8DsACtdfl88U
uxaorJU9myO26Tk0sR1gw5VdAOih9VHs/VdkuCairbSfHtjgg/rtZdeISINe
zHbymmLyPjxr3n7mxJy2tJh6mWRZ9LieTsy5T/FX+VJbbyzPnJ3a2G0aUK0j
iuXU98KkyHNm6vfFHmcvkib28BtETT3rr5v5WD7V7thp8UKQQ/14Jp+r4LBv
Q4bL83UPNAsq5fQXDzOwytUv+g3psWdnVm7qL+QHJlDWuMxrLXHjST1blleo
jSXIC2l4UYFACg7ucBeTnX5Y2H/7P5rvsS0vKd7RCRWQayJDBShLxhsUQ6QF
fAm3BZojNvs4119HWISFy+tQorc7WmXmhKdJPTLR3LPeKhPfSbVfq5xe/v1O
nd0HZ2lV0J70ZMeSemQhC+v1EAkxMTPu1Udrt8cX0Pp5Yn0miwgDErkxsFx1
FZfrDd3DJjd64CGedW+B9M1xNODvdmK+XvIJ2+ltu3yHAK7XUoox1bs14Rfm
yZb9yO6Q/4eEwuvnGXS0VvMB27Zp5LmdZKxSFzKo0hvwC0Sar7JOmcnf7H6B
VSLJiRZAsoClIahJDcYFjbcWizzRxvUBOZ+7HSjzovOD4zN8+xWm1ebuj7lG
zmeVpoJ3MRKK3lBTvl0cAsYBS/Tn/zMreCDGl8V4ztbeKc1iEMGo1AXfJxln
WXDZXEWEGcQaOQkSF/rS4Qm9dMA87DV1ZGthJTyO/0/q8fANaFLAXfvlBGe2
aFbq8bu4PquUG8OhwGYAy0qhobkZ7k/bddluDHamXCDs966aFsivsCjgjYt6
17cgtA2Ajx1UPUxb4rVFiKEWHDFZXADOk1rrg8W4zn9YciEnxKdivQCJYFMj
B94JDRjSeOfPS+hi15nJleXtiRWrotRIzM07FJe1DjiBcObWgseG42BC0JXA
d9xtQX0gXi4hazZKT7ZdHZMl5SQS7NquHzDILhjDPHq9YaHiremCOf3XdHhR
qw+rrbyDFrRixGv7P6Si/4pnv92ruXwI9OYOPJA1GCFBq3CzYU6VL+vXESvJ
r1gefliR/5EKIjoDeMlR/ZrHRw18ry6R29mL0TRK7L5vzmxHukiV1LPZJmHS
u99KGl6rK0mGJRp9pLk5+lxX20QfWOQjE17tVBQuoTeGQ/e0im9iwN430/Bb
2sMOPj+kfJmVIzP1Bjk6TZGyjnaaOsLn90ztznGQz/CxTMfid4hWEdATzgCY
SEs3OD7kOclUuK0Mq1Og04PgOrkvqCgR1+reXpOQDdRnFjObBJ/R2U7q8qLV
JfaIJmMNSbG0tbrAKR8mwqaGC/hOnr8wUa9uyoepM8i3DE1Owln1p8+9ZBOf
Eg9PAUEgHnEYmSXDSi680jjPnXKO4BesGtupzrBkTXMzgwtvQj5Ju6w9qG3J
rg7c3fSeVF5Hr79nkFXx+gPB+Ow0yXGV6muBc7lFYOIMm89EDdcpI4+KbeqP
pN5jGuQ62hvV1ciO4IXuvdWcpV3DEee26O+xQn16B9fUuhXTD9wdjxREmgt/
f1YzyhQ7nVQW2BIJiagDz1n5zYibCxl8NoO36Li+Zgfv01mX0STq5k4dnb4J
8Q9jR2iHO+nd8VziMvZNQicU3GB2vWPD1od1gzXmOdlDD63ONPwji+knMT/A
273WC10PECgkbjJQ2kVOk8a73y/MNAyUpYdUbbRx81wYjBo8zt9eLVU8rJ44
ku863DLNy4beyk05nZ9+Pshag+nZRbqcFKORhewv1U2h85HmJXLzpNMLxjhJ
w63s/hofrAt1oA7Ec0Z+64HdsiTrUzn4qsrVuyJNU2dRChUeoJ6qDRVymR6q
03+CK7AGhs2+ZeDejhUnGM4HCYt52qmjFCuRSHciiDRQE/dtq9NWhG1e1egh
27DwwXGZea67mnFumCXrdfOm7/h6/m03szHI7LS53VNVwbE011nt6Lr0A75t
xowG/FxlyyUfWAPHAqaoaAo3gm9A4OHEnUXZhSlO3KOnQeG/7kEy95o3lrHJ
Q4Vfb9J0mNGJ77/HeTw7+8S2/cnqtOSKroOobSPAu8AZ+GaXJZs781HOq4rf
vcGfef1CnJg35VcktnvN0wBvMyvAUGBgIfuA8uMk2PvJuoU07Rc71aHGfVXj
CxtY4GXv2Cqo1UKGPUBj5Uar0iKQckcSLiOp10hrCQQO7nGvNrU1x1cIS5Zy
ysGbhlFkMxCVYjvlz+rlNw98lMZ0jtdOgtnhO1XKPObwbVFFwxNeZNw1JCMy
62SqHnJKPFVO5Q3PLwavnCxxr8QAZH5A5UHpdM0tVErLZEk+9TIulkHU73Bx
on9Bw+H5PXDc1F8c/Ku487rn6CvlVLlx0OMauQBvznouRmG66W08wU/rNvWc
cDxwVuKTeCFJ1sd/sFcX4SFodVZbpjAigwv7VhKQYDTbcPwCpkbLkWqUzJV2
0cmUbgQ3nZ2xGy6sGj9eyrPeFRpgDsnLA6WTmFxs+LFcfjdOSt+tjDbj2Orj
iseNAy2ki5agYCov2BtUg6wPuky8BrD6x67W8sCNKQ2OmQeLz2np/vUfO3gM
cBmv0Tp1uKZwM/yEU/6vlTFcRJZpaowYVIUDMQFvXz9jmmCbft8Xu6gGWacb
O1w61jGNPfBs+C+hXhlrypgXWrU4bujHYL4R0Qjq8OpA11iey2cMhfenyTrx
FvWPkdL8C6pMg7HewVyf4CDG4DxGi8IQsliGsoLBQEPjughWhTaKtGO2PT3g
MdHKcX6oa4/mzxRv/EAuahCj4fJ70HO3bUadKrICYPUqN6JgPHLcyvPTUqY1
Ojb6POkg2X8Om1aLJ7a7KjSBzxp9medE1MMxPJxZRAD9Mrx/h0RNVhNUn6es
D9OipLs7gqxZOIO3ZfJbDXLWTdrjFWHb3NjVqYQQJqUBDJvi62JxGiF834Vp
GoGrJbjgHkfdSF1YVfJtnkddhPNS8jsmD1xyvD0pB2aY7JxgUtP7XI29qm/h
Wmo5OFgU2VK+SFneipPJvh6Q+K5bZNtAuSz8MboweQhOAClG57iO0qnZXVUT
oYxJIg2ahtIaJdIoLSvHbYUngXrO+uNTlPs6SbRad6dMtIvhYMtipTNDI/QA
sAxESau5e1Va6Fs7XU4Ua1VNJXpBs9T+ylCVDjpfzEqmTuP0zsBdzwUyE8L6
SlQxwP9aszfPsWCdoqIFV6odnywk3WznjkvLEKubMWCwYcz7AdSnXeAglnK6
LLveLcqq3Al+GhdIJEjRUfQHf8d8e9sHIkClJ3iqR73U9CUvPN0wEPvkk3iB
UYhVMLRBm3RWbq0cZU/nZ/QsPfAn/q0DxGX/2UV9Veeh4fNH1My/orZ0b12w
SB0Srrxsf1unX82V2gLqjEpU0G3eT3FQVhD8imDph3+MlXDo8saYuO2BvhQN
d7Le+3gVd7Gd78b7tSpv6ltjuqLbC9MUwYFjGVRVmJEbF/1xPlgYMGIffeQl
l4BEdfsW5ivrzUrOyg1BcuaXq/aqDO2IliWr0VFaA+Pmi7jnsZdJFt3HVcWj
eI8pwRgw3dgC7so7PYBOARJJFoK5UzPX3CrakI4MqfB3z2X4wEbi43SYhF2S
43w1DbuD+DIR/SGSyFk0Pf3MoSWi7LhliKTngfJ7B5IpqhU6dozMFx/qho/d
JR1SqzHrYP7x8dit7PkvkHSN9XXiV3P7HYWffzdrUqXAtrJ1lKyxQIC86qt7
Z5/yp6X7e1RCjS7nzABZKr6NM0gpU7M/u6xrbNifIHsoyWitdOqSIfc1bK9Q
r2nv0EsUEzZl/erEjrFdNkSZhATLbc+KYooVA6HPigjcviWh+ZU02hKA/Kzf
Zb8ux40Vrb94rXGsHX52UpJs8ftTfdhaCe9LnOORj1Rv+nPlllx7vWFvJ+J4
2G7L4KuxvgJbcVswQ+14E9BQGSRwUC95/+JzuumJXVPX0pH/JWUFEA6FqfsJ
W2nZKHdJBEmzHwbDvZ5LCrl2EE0seoz3SsWlMDJMGMzOJOi+4+WfcdIdiO3y
b0T3ffbbdCsyU62PcUCJurbJ4e0HbDYrZr08U/L+6WLrelZRjKHAkZALw9cG
+0Y52t1vR2rZ/1aytMcsz3pIReI1qmx4GtRhPPSRVt5OrNUR/8gak8zuHaeG
X8moTpgjt2InlWfvWw9tV+NhvZ8X32F1uKsE6OyrTBt3bEOF3xRDNAGUFk0C
6Pawu949iu6Rt6YJKztQzIiqbD3e1iY83kl8fGWZ9D66MBDXK7y4CmX+iYtt
iBafOPTp9KmmBIIXDs9XUfv6zb1nhYR+tMUTI8OotQ0j8Fis44/f5E9WKaRK
guDEe81jqB5h6Pk8q6Eh6vay0zNBZkj7YylNPCzCpmBcbeHWK1AzsBdmb9Tg
hisIw162sNrC9KkyMbmuHHkuBsNxqQXYXYIrnAWWTAXxlJFlzmKhgG2AGL6P
mZvi2m0T5LLlE7VSbOVUSGg142j/UvqnSmJIYhCiIHGkzNhK8ZAg+2E1osgm
f86OkmGyOK0+CG9JUvi1BJd6s8gCFnc4ZEC8KW5tIaXJgI7j6Hxfj3kvvPtK
gmtruAhsVTVIFg2PqUyq4zGy/MtIx+9KBb8tiX3jOdCt6Y1ag+x4eUefO8FQ
w6tbrr5bWIGVOq91vuhGsbo4kf+8dMgSOU7HoMkNyMPQJHV+Z7+ex+txxfzL
+clugJ7bO3SbHK8ePF51CBjLya08OA7G33PVKgcwxIZbLh3aYPN7fq7fBhCm
ZJSRKVASMlGs6ZWRXnZx6sPv7G5vURy3yoUCwx7ev3VnrtOW3WWRv6gsjny1
uQdqCapWPzD+Ad2i4r5A4q/BFPrCxIn7An80go0s+asWaFG7cq8jqzGlJk3g
/RxG6Ntg/CoQ39TsCIfgqD/k8rY38lTduBlUV1hzNB0IUh7yWG5ys5NOr9aM
9ZndDFVPLqHI0ynC/K0kR2s13IPVaPlo1mRpTMssEhg+DlZcllJ6q1FALLS4
aRhEh5bWsTdi02StO15KE5iUP+0hnpf73RLd+kuMYyk2Et1TVDs8bPqeDa1j
zdbX9AgWSOAcDPUV1yDnldzS43HX7P8g2194hz2LQEdKBWM9EzZNqH/xsMop
jfWvITQsGGD7zGaoPcvQmymoae5OizJOIeRzsCqa0OYbSnGC+o5pEHt4c+55
1XDL+1domor4iU34w07cRaeIDoM8Uiv21a6cCGjveaZAdRrZqDgVSfwFvEbS
a7xThapqirkEZ8D5Q3ohvqMRrCzVIgSYC7oYexMxxrZtAqTwww2PGiihJEEU
Q13BEXqfIwJgpP7C9l2c41tA8fOzpFhaK7PfwV1h8EGTXJoAM+E3bBZq7NBH
zeTMwNoFElZc9Z88uDf2sabIrdG3TvX9GXL3sURahWpHbgqCFTB6cRtrPX+H
ABJSz/U85yGHY4MILLfOwOuuafkxTdcxxLF76izamJ+izM8FnTWMPc/pIkwM
GSeewgyIKw4gK/Cnk5nkuB1+ChU06SQUCf7PHE8E4yRr5Z1RR0fkuFi5YJIJ
Q/kDsZCyyEtlWuXle9JXMhRdH0QxT/3flbHIVO/HC1LV90qzWhSKQwrh9lOT
MpspaPz+CyP0p6UeHfZ+rPIBdRqc+Iv4I4bmu3o/0nrypNHE0m1XXoIFnqkL
/P/03RkTX+yp6U0g7nL8/A0icCy6M4dQ05nbmp9ktEXjwFCoj/3MofPbZ4wg
YVgEIopPJSB2h8uZptTL5gz8FSqR8fGChXB6rGRcpMPQ9kTblp9Xj4K4aTus
yuKnuLmHQWDzhFO1ieNcPub8ZOixtFe/kMqo8r1MyTwu1FTcg+2Cu7A2Dv27
VjP9Zd+i4Zf+zPc/40PMifHPnz3THSxbsaYPLMt+GXGplDMcrKEkk63PnU/j
fIlb7EQYCsfR+4tpmknBpKqEmf7+ePzqQw/5n37HdyqsGihSkIkpBr5sjNge
2YcuqMy01b6u0miZ49V4K2IF4Er/fpwCj335YmLNQAAEkx+DfrR+thHJV69q
JDO/C0LVxxo4tNOKKhvUsfSiRzi9322bfgqhmva88ct/mXo1+sjv4eIH5yPc
38KNhJc7f1m/yQJANz6kVi2BXQ6A6H/GqWgK9HJBKlw2Q/WqlelC3wA75Tlg
mdWZsvhm7+O/+XSoVaes08pdMjHszWL/5YXhDHSM2b26raUT2nrznyYqWuGX
2BQXsAVImP5MgaFH4E1qJFstP++DelSRbK4BvaQT4k+gtG58jgmkj+nooLxb
LAfJAHbNmUSCiC/QBbSGsssJJkhOH1o6WPxL38ApQcxUbHVq0K2JQclp1YoW
yIbZyJWbKQR05dFcYz0E4exd4GYvBAUSZyehKhSHytFi4CmDjiuvFLf1kcBb
tyQNZlx1/JO5zGc67jfobumi/FAkyWQzpFwQcl+yLKfBE3Nr5r7qTuhwkrZd
RQPeVxC0KNZXoIzxoqUOFGTMl83q+5VdDnQO3b+mcpILdFk5xEGcIgJm2TMl
9QENzCygl3bf9uoxomwjC5O8MWlU3tCaC8c1nlT48DKPtSzNhW0vYqVpaNND
d6qaRVvLiHdOND2vJNtJRTk08ssvtD6LR71/NpzhpZQkOwjNMNdQ+UmKoKGZ
KreT+6I0w1EE2xx+mdbvTa1dBacZMvea3Ygi1kHSjRzHRZyM/O0OwxeNLmKx
CDeZAGoafpqjN7j4IdrkJTq+W3a/P61qEZr4Vot1KfG07bwFq6PzUTJK//1v
sGBtuZC2mQS27Zw7hW0bSOWKhHpamm+N5vvfueVY+3lSFsDFLf9FdX/l78Qp
q79+RxyocvKgUKTTWvJhwLm3Q2B0kOBSDRf08P7qNe2KR9ffmaB2qZsW9GGU
U4nsGYIqJK0hHkDcNOiWSOslci8ucknwwbSWL10Z4IkybVY5XwWFxdZrXC7P
WMMkpGsa2Sxb1mtepohrd4ZeIsf2sgq8t9OrE6uWCvCbv65ArhHSVoXpdqct
W4Hv165Klgu9Ed+Gcz/FDo8EsUIoIXCQwuytH3OWQBwZ8lEfZjQg78DCpDxQ
ZFdSOIVQHBF+WZD78kDg235wtcEBT4bUw6pEwNR9E6wFNqop2+4CzRZ+YDuC
MYrCtKi3MS2+7JAn5dmFy0jRwJtTFyA/A0QKr78oWLgSWvMYf85u5gCELg/t
205LKGVRqeAf288JrlTNboNDR7MVW5WcVhG13khYCoS1AJ+yW/dNzNHAKvsF
Tn4ZhDTf9YOy20rbATNEiJRubquBIsGn/bOsX3IxXRwpngcAUZvEfo6YDOfd
X4byVjv0gtyWkn6dJhgZ6wdOkSg6qFjLpG32SG1LN/ZnaQewNFA4uC41UjMT
156H/8xUg5mv+IG96205CLnHZMuZ0E70xU+nW5zxuoaz6LmTDJZhAF6hhqh5
MII2M8oe6UNPrOHHrsXoWAUwo19zQws6fGUj3urudiFM/jIcLfk3woX4wkN7
W/YpHJHaPY8RpSeU70pBKNw+906w1GsT3g064fAH2UFIXgvHj4PC/QoGw8oU
lu1+xfMSMgwksBRVg/yxPytTOnhqhUX1sDdY/KYiCorZYBeET6092iMB7AMm
pSq3Em+JaXZ6WCHRHvtypCh9Fj7iKodFousrVvZEhOoo2WBvi5+jY6YKnHxo
tEuEkjG4UiA6LtXpJ3svQOVQ85gJakmu4pwnD0015zfzKORyZqWGaBukByQT
TUo4wIdTMYcVeRGKU/4s86nX0tMPI8gRdlHr/Zrqc/4uR6F56PSpMZvwyk8H
+opvxwlr7BTHdaI3XWkLwPsOcye2FTlSP9HJLlLYAk0mxarQCiTNrLm0ODwx
EQrIxf78q4EaxJ6In0cXfS6fICqQTwBvOair5+HZl3iizz+fdL2vpEsXINpo
f254lNCHSO+Wqw4z+d0wUFuwTPWFAFGgWLOfF4bCkkAKU090QA9zcnL/F9Rz
OBGgtXbQTylvciGn+HApTs90Fo1LHPxk8VvcJ7yRE9IYn17X01JRWomLmaT4
+FOprPCINVpayrgfRubzD6CUz3BjbBGvtIIYTLcq+mZstSu+31NQKrU7lFmg
24hCSYs2mjIb7y2j1vSz0+f8TQrA6EDRK1FF31pECFnh8Qzm2+2/3sjSbng/
09S96WGA480/k/kcZehJbjUFICxoYoVJThaNZHHGAuZGNq6RbUP1fTDWkGuM
OwI31UwLgx6CNiw19sl1O8lvQGjRZHuqHH0f/tVb1WFIBRokLKAO0sHDPE3i
P7RsItqF7HosjeqFKTrV0T7mcHAGLZR50tXSCQfIvej47dATG/m8qHv5JM3U
38KnUBZXTwzsZJSD3upmLh9/oCDTdMGwbUaDL5VHiMx6kpIQHIZMzASfwOpb
cQfagZXOvepo5egbTZOU1fJWmeyagvb4ZCuSB+Hj4O6tH+7Tpsu5ABaiWMFc
Rn8TphFvljptVSpVQIhGLZ0+uahdc40wGpBsNAAITwaUhIARPgPafJbWe/H+
CGjeM5UeWXwLPlCu14+/ay3SVQVQBOElibZa9AgMWXCvJE6Hi2bhFDAj+Neg
ui9NRh9frU2yEoR1ly5ec/TEBUwTYA2wK3sElR+L5QbrFdt+7VXGyaXeaD4/
jt7zisByLhj1qXRqcDkZn3jLRH9ZF14ZRYZHNzEiTsF0vhNNiKypqd7kGNVB
ioNFbHTDq3R81DKImD7IFXcBfGRYk+6JaQSh2v8M+h3uaOKX99PDEGmWtDat
qSQNBKNrfGtkzZoARed6WTTwuLL2APb20Zzk4bvTKNc45C3HFNFud1d7o+LJ
WC6KJz+maVgxtshGgJ+rvkHbBchwLKLG31BeuETqRzK6EMs5EoA6a7ixVFgH
fNcTqXXK4eEu/5VtscNgPtJngMMztHvcGHFXSSWhMWb2V5AvjhSfGGC7uNit
dMK48JxueeHLF1ktK4KsLeEGnLv3La2VIywUNfjBzfcRZaNDkCHOW2abHY8w
aevqZ0DDYVJuzrqLMaSf8cHAgXGYYe4FYB01rnVgAnIim8ZdM5ZLKJ7YqHc2
j0ry9F4vzXY+U5494nK5TQq7M0JxDvZolt8VF9D6iJ5I/xmvgH4CDXzlqq9r
Cwvn7D+Ruz1RICwmjoGTO+OMjyBTwR142ZF1yKMD/92Ri9jXtTtW6kY6rplV
Gy4BoEqbC7LIsdu+RJl2M5o1kmINPak14K9pF58tK9m/dzHJv7yq5MStqryL
z+2QqJPzMPoOkWwk9ys8pe7DtyaCE/6H9zQ9tL1Mx16F2hsAeQ99izlDbJyK
GZ/JFHp8Nbwz0ppRnVBoHu16wjiQdXROobxYZil+o6n8V++iLxic+GpvbTWv
XE7qScIiNoH/RXDdDrks2LOml+xPlCJCEyh3unKvKxP9g2C7i11JgNg4G81Y
xziRFzQbKjMLQuEgtS24mA5ZAuy+UPb0lESSouNF19xtppEmsbd1oeCnWaj4
xAsAR1DWDJ1UzR57yjybrj3H/2njClWeRFLRz2U2TqU6s7Uj9wu8q6zdJhZO
2jiJ/1xOFrP/QYPBE0tr28Yno0eVExhxP7rjv9WFJdoJ1ZcYdP7xaaX3pToY
pyVHNyWpaAJn77SbNAGhj+uya/EqiYtSnE6BPDWqt2YPqKtXADJH5HeerLrS
OXZrEqeF+l1kTStk02WKyFKmJb8O+DkO2++xHejfRVAaSU9uWDFNfuFmvWKB
F5gIk7Ku89dfmSJFnHF5qvxNSSjoCOdDj0IiYYlxoWePCQZ6J/nj9sRItYJT
S9o3kYPFUXpJQCh24fEAX+QC8uSH9vZIsweEycR/KQP5C5qY2uFGGr82IRzi
W6Gkk4WziLtHEOerx4bf6hvEXuh/q7q9KERyqpdITWyq6xlyrvJgMHGs9dtk
ZRoFabpi1zx5QNcgqVF8x5ZmFEW7DkPRZw+pSMGwAxbpbU9Y3++grDSrvHJP
hJIzpStxGbDG+hJKoshfwkxV7gF8AsA5PuglGajzDuPYBFoqwz6osUGrsRwE
pyH51IcfTD1CVlXa3U6ALv+7w//j3IKkWTaa0dG5SXOszxgSk6z947KnyEM7
CmZy4OA/XZW2/K1GBYS9qCWarJGtmkoHECz8y3a3AJGn3FT6336w1+w4yVTD
IspqKkLXpfh/LZT/AFxG9ztZxYdb+oSZed3SEW78QbYIeLRCIBoEOf8wUBRN
I+76ufmO/51LqwIVxQLAR9fyxirIfGMi3L97EnGBPYHpw0r1vj5HF6PopE0e
bHY7yP47BOGHWZPpS4CeLT7EPf397O6pA0YlnkaKVJw9wFmmwsF2DsIV1dqT
1ZQqD5SufgwFbf287wUjMOjmalNpXFBQTU8aCiIhYXmXon8PcN4zj6IgQxd6
FVsM+7n+XA4tUvzYEtB3309HcqNKz/fQC3ajgSFX05P9l3AXIYQF/mdKblr1
7houls3B4fB+xk+GeY1gXeSnqQld7KzqH7pDScB+sHahbiPin0LtZNziSRbA
wwP5wdnMCddBykOjlBbJBYCeu1CxisLVjXHGdz5MNkGvGuOjRx0JOVWC0v3x
xWhdOsgvOzJH4LuANF8j00F9nd5d3h1IeLnXf06oFjsfS+8YOvThNyc4gHWC
MXWyCeuG22o3PRZxLq8jJnPP/b3eNZowoeUeGigETZJ87CXaeUE1aSWfBs/O
6SH+4ir9AzdYWGvjoeAEhqDEcuJQ512VF11nbDVqbVpry1WUflBbKDq3DJgX
Z5e4Ah3XBjcrRY/FawDJULNh3FOugcMaVhZDOvHoF2M4lorMPDs5qI5XUWMk
0yrn/yvi6t5ndkupZavUEijoE4/lz4/FmIi21WgxBZ8BjARMVN1JdHZQMXQR
DwQgSjdJa1dgHOVDS8Jy52tV3Uqx2CicKKrCA5VEVW9ZYaJylJomClH3RNXo
85QXzV/h9JA72eMmF3EYi3jjbTfiZnqGdJJDbEMuYvC26vYmQPvI++YQTMVH
iac6oSOW1kIm+QhKbjtrUStMYEsMH74ZmnC9NepaHb9RwHUUt5/qT0UnsRRj
JZPnXq/xtTYdXIjNFy4zmWMlOI/kKzrVF8Cu0jashCopghPakcfbOX8g8YlQ
/+t1PWouJvyW7FyGKGsvsJbBtVqRWJ4CuEjd8vHxlEEla64doqQG13hWnBaO
q7UWJ92p4sacSFph9EeZ/dp/aGn6tGn4BPtcVcc4faeJNMjU5RuBgzAixBSc
oF7Y7YY5jM4QTFPAIYVasaJba+i13r3xBcXYQNU2clK8FLEOegGdA2le7Prt
FgdRtrHgrxLe9hTBdJxhFP6lLcU/7J1YNjUReoqnknaTAFg76b7XWu8Wz5Jx
62krQs2SoGWRPUB7JtP7oVx9NN5NXbcl+wQ/ta/nkTaOL4GTLZFZZ8MJ+yoM
6DKh879MgkaGUqSBW5bNjI+NQBkzMlJKLcLVjQgMJuN0KrM89CsDnF9G+Ubz
CtZ/QxBS7cHUxmpOQ5lKE2VqOhbcoraA6UtYnwub2ybh9xYRRfokEiPV9mY0
OMBZvWHBFhEtV3/a1Clh2ex7W2/820BndWKKtOa4Z7i2pBWtRVLWo+WAJAiR
wEwaHaBaRfWK2JhCGgCIF6YBpYXsiKIjJPKLBH89m5bsjMKy8tYotyU0E4Vc
Nl3my/+5lD4dM6nDVq9OkJbKAgwX54iC7tP/7R55dcPKVz9BtYk5JsK2Zbox
QAOpxmyI/VNAZRwJJsVLoLogTZJRP8VTobhsxcaZXX3hlubxiX/nDGdwJcwz
YL6+SSgBP4QHlfgdxaN4RCFciyOONgOAHSYVDKcQszq4gMZP3j0EuGqdc92q
6EwXzw2KrM8PCa25j22eRnY7cRwr0Oe5wcYYOwf0srQmHtalYUQve1pQUw7g
/913aDZ/unA2QzZt4olqZ6BKVRwxKIk5HWygM6OvZH00d23UxmPzKbwfTPL0
M+nJZzEwQE3omLJIRmB+0kDz6W6bpe28N0RVM7Ntsts8cbO90NsjAJ2WVMuf
O10BBBfdAXjnPjEeXmkA5QktLKQDcBYqyJ5TibReNIRuEjhPqoqR5/fgcRtM
+fz8VElMYgDNJKzDmh22L4oTdyTe9cq0RtIP3D04I5sOGlh/MCCzwH1SxZ6r
SYU6oFJ2D45aUAc36gdyB1EUSoj1R62FFE1mY6Y0IBj7wzfOwGNX6V47+Dmz
j0Vipm4hEYpb+GWE7LBip+eC4S6oq5czyQKaa4dYd/dT6FTKKVdzpQqkJT71
ubvbvO7XhQJtqxJ44hLphqBtPzI3CtMgM4aH5QDIx8DxbsXo3wYGYTToGif8
dAucaU0iIeDjIFLDO1rIKr3eGvlZhRiIlFRyOrjOOrpl/xqihCQ4YCBWtVFC
paUjMad3nKELQrQhH20CNEj/6VSdZvDGr8QV6VJZdOchq9ItZhRDGEfpzpyy
C1tm2P253rBkrdwL+q+PF7iXPEj2QJNM6aYsz+uErMrmgPXlkd2SfgDtgkF9
I5YCu5VER76iTKIPJ7ICzCTxrGlMqnPVeD50RioEuGQMkC8RxUL2fSTrvAOM
1nQJ4u8VUGDNeWuLAf7EXhSsiVDIbiTVCXxNfUgz4QwJj4wUeBtIoKbd/xtJ
z1k+IWqQQpn6IUbJpWhVzqVikYkoCRPlu/C2laYO2LdqpGx11WxoBdZWTHCu
7x1WMKJfyrFWDlMn+K+emw4jgrcgfy+fB7JnSas1xBbOYEqu3WYJWHkj0oB1
KDRpWsSMrESrUZfIz4ED1df7uPiW6eD3fAun7qZ19588L8nK9ZJG7eDtfjBf
pIj+LsdLjtuR/c0AY1/Xw1LLvGx0r6tkiFTuWSGqZLfBj7noTNjdCC35c1VS
RJVKMFaQHwhC2cRAe3qe0T0Xm1SGUi6PVVdmdhJ1dA7V/RnXA7aRMa56InpK
4/Faj7HoBejaM63JhgPIyA9rj2ZHv6FjadQZOFwpoffNf/TekqKRpBxHosEZ
KYLPVMsjcAxw/LEHxjol6N2IKIFOfs2h3lzEwIBTVScbnkj1ebsV0rdviHmR
6Md+IyI74O0stJRXjlkRPFXNh/uDce7qinSWT85EEn38xixOEHh0x3PqklAl
Qj/2Pwv+o3Eks3c6QeytNUr6pfR/ppfmrsgCj9UtlY+GfImWodyst/iShQ86
/Wtnmd9wCKjegCb6VbwZmvYC7Aj3mO2f/sXg1mCaYPHEiz8/ER4Ge/5I+W/3
fDo1WdfFO9OoRxkGIHPy0nrhXmb4QvK7tR4oka0YosB1thlxgj4NkpCRv33i
bQjO9nMFZy9ZoIfHShEnj3XC8lZ76M0VJBRbopAB3v8tOmLMFmbzrbYZVDQu
MCEQ1CoroBwloITBlPk7In8aMxKN2yaD8HdVllIMp/suTYa8wq15tYjNRqbz
uk05MyRrSlMFWOsY3YW46msGPTRRi9lJoDiemJC8zKKb3UUG0OzOnQwpm7QC
QdhcZRK/Y1eGdHAU73KZzAyzo+suCi7RDPv6A/I+64WRzqLV2ioKfUJW7o7j
3PpT8VOjFKN/xmURE6iE0PLJXwirYGOqaqlN1hWwByWZIe9YuFYj8Uq6vBqu
Dtv/tBm7+5qXyW51xPwehFC182ZBnUnzz7K6RQMsIK+OwzJZGFUI53bqjgdk
QnUCwb+HM3JsSVn0WYSahXtVL5+I0oCiXy4zvMHjePZ9et+/d0cG1rnMyUAu
zekI/5jXDf4I11do5JwWfWxkahjWqkA7DKFLnq6QYX1p33UGreF12A+xztl6
fim+RMC3No85u2ybphnEy4aPBzusAJPLIgy2+oYeFYwan31KwgLEJgRdizcW
2ebro51tjlEEksmvYjgjSa8mUJNWj9FfudWrccPQ6/Hi3CvqYhH44ksA/knF
YpKtjk8Jpe+57j8CNmD7DbkDsvuIhyfeWRm86dfjQdRmEKHq4aKhotcDETMf
+qthj9A69P3UVcl4I8YPLHS2CPnUgIs4gNpuhIEfFbv0nfW2YdUPblGx/+Ap
a7WuftMKW5SS4icKpl6Olf8uNEttZdS/2Oi5V/gBu33T7T3VWx+A7jDt3Axi
RGN03pVRGTaI/rA2dZT0EbDEUOxiYbyDs2SZjlukCjflIfMqKJ39ls9kPuRU
f4+k6qJsmUIGJhQ+1WlKT9BSehSADH4Fbzh+AthFbJD+CqzgkbrG039CtL7v
PnsWPh8aaAc+xQ2yczDcL/sfxRNL8GZ1/bWHesPTO0aa6bYzo+23aRx8rwfm
4L3oW73+RVXCZFjOnPUABdJBuh56Wj1RGStk4KGtaGQj1FCfBRHrAQ4N9Tpo
MusuY6lkDLpto45WCy8DtslmOOtdjsLX2CE1BSBu06Zgqqc6SzV/NHEaDNac
uc4y4Xn74nw/2kyMk7UYLZ/EnSGaJSOemFSCqWYanQwaHMxZ6TMB/b94gJoY
NlPuMHF+p23tFDEk1D7BMXtBlv0HysKmMY2sfH3UiTFMrBWl0n870VbHvO3k
AxzcJyZTg7DI06YVI0pll8ty7osuW/kEajwHvGPBeIHFkASjxgZb1PvfRELE
WyxY4N/JCtAI/7ovfWmOpWnp4Y8y3+K0EIaP9SVVn46Lfs7EYZUpIH3ztuu1
HyxArf4x36yauZf29wBLZ1YTlun40iYMP9qFebc4IexFutE0HjA3px1p3Hxm
kG3kDZfvKTssw1J4xBn8hNaElzaL1LuFslLCHpnIAo4m5OjVul5GrovtPI34
IewBjcKOpJCMVND07BMxJClsiDOzjx14Rf/cu28LMT6tRS01pCYiTRquO+y4
5mp5PKdQX9bvEU3TpKjhTBt0i+5uPregavGGknFFt0zhyzm60RicsWwQRgKb
VnrpC7XI/gzQGpNRJBQo9m8gKuRYT5UNSxXuQeYIE69aejufWIDwb+C1wRrj
rKR/tGKb0Z4WYEaTc2HOtK8zXgviBZP6WxGkvIFEBHAUIhQ9I5W60SPpB3sr
pxGm/iuYrgWxThMM5wC257JoYpygeYFu0YGszlqzufCKSw4KQc83rRBaNytU
4wG2WIXxyR2BLwCcWXXlLZM18+uDzsDi73w13Uc/FIkOZEd3oP+CBjelcups
OFqXk/UNUdw9gcvveyHfO7aYmPHyzQMFhiCUrOrVD6R4Ir7L0hiTwlS14/Xh
ZvXJXFJ2W+2BCshRjyorcFjIFTaFmA7Gkfb5y9JeWS95Jyf4hBGWUQWK86RC
zHH8g2Tc5msUcfx8+xxnBTLsGaFqxvzQ/E975UaPXBO5FyOGn5P51M/s4R9f
PGAIOz1ZqSxnOr//idgVvYF1KBeAvrajZJzzcd9HTGc5qN1W30b6aq+rSmGl
r9S9hvJS8ux0qMZKxQdJY1JaPLvvJb9yWgWlS6wPP2AdWuekyybEaUSOgxiF
fljoDH+n9J7o0dbGnlWQrLdb+RGiGC22BBRw2Mtb3E/gquiYCVIBne0O2DCj
ipR+BLQV0JKmOAoqc31uu7idEkgvK3SUV7uVIvNh8CRGwcC6aGbxC+wrdqxw
0vm6fJ58rRH4iUdy3QayQc/2/7eJtdJ1QZJaVQOTHpe9CYjF/H1FA2IPJTX6
CgG30GaQRhSBvqrrhxpi5tHzklry0Pe8KEle6Vbq10mSgtUISQMIvxfBk40I
QeqGxke/Wir5IfaeTYb2knrFeW5IGXRiQxK0qtq4Ddqzt51dhyJG4p7b9mN8
wIu8/+gN56sOgW4q3l5fo0SSasS9xGZvcHeaZYDK8KG9eIjtsAoyhmMnt6he
f+OTxCtGrCrxq6QaQzzwuTL3GCpw7ggJSdXIbyY0r8x+gveZRR4Cm0kacRjG
qX7fW68jBu/gyRBjhPnUUJ7HJi9tnifNNmoWVyxW7gcoJAlEHP4SoWVR6tdv
AyAYcdjDkK2tMKAUlXtLmdUTJZeTIU+AkZfwjo2rs6UZ9m/cTdhzGTbbHQAv
FX7oEXEplQPlGbcD1clwcgQudMSWxtQz4y6tU49KkfRSrKzdAP+9M3StphNB
BceR4ndBgD7Vye/3g6wXwdP/ugy6A/6lZnMDndSaODzHmk4DyFjE715YjX9p
UfkwFaTHKaQ0gvZcrytLJbtsM2WPYt8EvAhdACx0FiIl0gPSkzNaLsl0AyJ/
Kvc5v17g2JkxcM+mVWcf+vitBkFREcTIFXEpW7nk/Dhjh6it1GKA1WY/vnXd
/+ay1bRvojnysSJdvDm70sTHhbt8tCb5cD3cx7rAec2M2itYFEMVW0E42u2+
Ch7p17YRzvmMxCS9y7DCDMky7CU630q0y4+ek6bQT/Omalh5k1nkQGTBB5Tl
yOG4mz4L0fceeZXrGthdt3VdfaQp7zfsVCedNwCxCg3LMOOf5v6pqVBzREXJ
mK5hViST5Rcq7IzHmlu0EE2bOAfhw8FayrhqtJLJ2SlDuylcqsbHHmowCzJS
7KWO1LLPiS1EOsK8WeFp8rjeAI17axx7Zi7TxuUFpnUbEAghlxolVJDAD678
9KJqXSaOMxnzsita5zdmE30Yv7/r1GrrWETE+729RFbnI+0UuNzLUWBOgdG/
9Ec5LhjGCMynBBK0dr29sn/dGOmJymQAPzmviehTWlwdY72YNOoM5QWiJMTw
Q79mlGoKKSxsUAv6p0h+mmshvjWX1gm1HxTVbgZnfLmqFzPgbW5qqKQtS0Jw
npcIsMLF7v7eMZOdXxQ6JmZ8/Zr+BhH0W8qFUmUAjpQXBsDXRO4b77io73dc
myJ+nznu/lVstPzFa5V5kdhcI6nm5OH5QgMrmm0jPqvf0mFk0fniBbPE4dIr
2CTUbjzbNoTNr9vxnFQ8GgeBfLKu3pYkE9HT43nm3AvIgAZ5u7jcxoMLXcac
XbcfXjchxT5LdpQoBbmWWI+f0y3O3wETltw3CxE/OvjxKKlzVjwmNLvcfSM5
4vl8FS6rydc20ZMNyYvh2r6NWpjWC0akOS+ehOtP1L8cA+bhIwsWJiJTrxt6
zlBTom618XBqkUW5555UwiAtgL1l821UVBlC691zDv0XrV1HV+aojKBmcdRW
QqA3yrZcIVBhTGRA3Dd63VJwUsoxkGvHxvsF3Fp0Vu01LrgynacrnPukdEX3
ZmuYHsZsKeoa9/6+p2wmXu4z4h0GWBKwPw27Az6wKU78ZY4kO64aqYrVo9/U
k2cbhF37pOtHNnNN6ZaInjtUbFSw0JnSoMTFNlB5YGQD07wdSeNA9F94a+GZ
rsik2wwF8+uagPKijsMkGQ4b7U/i4XicAjREO1VvBVlk3P2AGvg+uPqfJOBD
+ZQQaKqSvas0dRqhLuqA25goh2Rg0tUWS988lbSr8fA3NxWx1W8lW54kkJt6
dGOTkDvmFMQnaQFxNuPiEiOnssIzLT/9OsRYjVBoBynB7X6T8xse1Yjprzwf
56qmYuLd161GEPM9BMPfIENo8SWxXgioQwq3QK/Jbrcq9mo0SwAQPeu59MOp
dkbRwHm6K1+tewnsgQ+2uHfBB3fb/xvMuljXZLj0QwplzFhAOyOeOdwRCFcJ
p0LS8Kp6lw3f/aslKV37/yP3Xga5Z8h0eAuZktNIrpzfw0LgHxYJ39EEG0rz
JP6+sGnusqsLjCItobp4If1pCzFkBH7kO8gJJ0PNPY8eUFDLYyHPV4pmvGDp
ipm6sq/I0COV+X/uqKv3Oa7EG8EnrcU8rKVKf88l3SUntn5piBBDc7TDwZVW
YX++b67yCbgNEQYsvrQ2EVwAymzvzfwUrddKctPVFn+iEgN2c8usmeRBV2A0
IBvl2gcJtm7Fskg7TNxrQI09Snco7PdY2GdGIvpOp2LTmgeJ7MzwsVwBFcQY
yq32LJSWHJ94/BAzlvumyrGgMEIHNxk5KI+happQuGKS6EcDGOH6za72S9KQ
fb3ItOFQdh762zzFO11SE9suB2JNTM5uco2SLQSa0GgC+0RAPOt1LA4eGsoe
VhSoz93fI+NyOpUHohdO1IypW+s4jEO282VV760r7JEoEBYMaP6S5afyJE6S
OkR5CbUeyZ0ipUrQq/HjNpGpDL4HF8+T0kcvnKg6qst3S4TaPBZ0bovHKpG/
0vccRY1QsVVm0BtLeIXahPhFAhWX00FFSLqP05qbb5aYJSQz98jnUycRgJHZ
99t6GmZhUo0JdTVnXfTWYWe3pSrDr+sSp4CNR2/EDaOAUnkZ1hQJA4M3j5+2
m2/BHLsvY1LvAZY0d8bz2Pv29wX6s/xO5m+dQ9x8a3wHNg2T1t+87YAQuVbQ
k4RuNnDvIIS6WgOpwH5g7etPhWrFRidIi3moHwaVW2skYTLoWZ6FJek5Id2B
9uENFXB++8YYtjhO2wXXwymfxDgNW5k2f9CpWzZZYrrNLcXQrQbU3yG68YLQ
FMB7MBxe8CT7ChzA756dkeVuiIcvBvTP7pCP0ZJWrLvwx6X/BmjgjUg8jAQ4
1a2wernQO3qsVUsX2ZgHxKFYYbeAZIZL99o0CdN+w/CbI8qHMO6QxXJM/GOE
flwW0DRk+5im8Lo/Aui8Sl57m5CJINKP6wVSG68jZfboYTkfeWB6s8hf3G/r
gTXcrBtosa3YLfFQarAm3fvFiIrzPcF5qd8iDee/bQyD8SUZFTK+qXEPV2ZG
P4blxb+dXq2zDtGNTBfqAUBHoacyFqC/juPKPHDUE3/yAFhR7Hy+2KLpyn0j
7lBsSt1OHOY+90kyTbG3sfF1/Y3XRXSOf5hFbyfG87XPGCAzkPelXIAUjIjH
eWhuib0rHi25SBtPTXDFoiyiX2u8rdI88UWJSDD+Z2335X9VtRKtQ7eRdswg
b3whuaWZR0PhwJUMr0PeibJtenE62Muk/BTg1w0tBujpuSmB9+kmF7BP+YbL
gBrFKWMi4kdqPc7bIHE7ohSqDjqcKrYw1LNz2BwTwA3ocFK/kVN1w+r77BG9
rxiMBZJ4qBUygYv4fk6gJlF5gFgI7R11rcJ5tPmDHbv3keoPuGOmXm+ooMWM
eg4B7E69Gm8EJr4klhlhYd1KR7uig4dVoLZ2u5MRCDicTG5ry9An/DwKaa94
3+w6XWJ2Kz7/2H4iXNN/FYsVh8kl8D4ME2xYjzfYheTi3kfXaR8HIla4EUvJ
O7Prr3AoRWOMnqdVxarQHLs3fx6yvY4uQU4lA8LWLCsbBebVHwLqrkKSPiww
hjQonmFqH2nGjwR8JF2ipjYLGpuyUeiID9Pj8VhQvD8KUsAoXtEYfi2Wq18o
32dqK9mokV5HiruN1G9iJr5TXfRDpPuG8xW+UZ4rGpO73CJG66gpj48MRL4s
xIrWXkeuBmp4QSJmvR8Ewns56RHCpDUPH8MS2sKxYIA1OzbLVMazhPMTQSsV
IXCPMU6CE0kETUb7t43AiKwul5qvaSCCDdArKsHxiao4x3T+XOVr1lz4oeAi
29eHbedbIFm7+qy02BrNMMJQLC+VzxaUl3dQvaP4mqmJJqN7Vx2rxricp+XH
sL0P/l0T2yjpP4JzZx0mfdGuR5z6M+jctXH43xp+WthVPb2opLU3REAUm3Mf
XqOShBWtJPLYDM45SZ0sSaqIv0lzApVsZBZpwTyeSe4jtvjQcMASeJYN98Ts
id2nh5fiUDAdgP63EaMCB+NDy5xHEzDbe8GKMY/FLM6NPyIDGEm7eBuRDagA
fMDFu1POXLFbkqYYOniGFgWOe1PX3WmdXGu6tPACyeHgaztmxybHBSjUbsba
PxHPf4/s6cSsmYVmwN4ZgiMLCAAzDVWhnZp+pdtRs5/wqGAQFOANlpi17tG4
5N5OD12HYma5n9BcCLBjds8QUKYVDw3CTe+a/bKo3e1KQRwBozi7OH45tFJM
W0Pc1E5ndUA/x7yXoOBQF4K6xT5lDk7mAwESmOV1obFvDz50aOPCEupniFOM
y/zxFgwCZZxMfL/dIy8TmDcH+4+UNUgVqBIBwB9eA/9m4nV97PIkSs//+D19
i+Ly70UX/tEctymMymI1ZBi0PSCyt6dts3ro1UxGkjhkCI87vnoUfXTh28ei
IOd/cMKfoUGswbZsksCf5y8ciOfypnyFl/9l3tqPc+utt/VThovMtuWwEeCB
cyQMIl3u5yBvmaCUIESzYACRmy0UoB7OQHsRFgFfBiO4eg/2f2ZKa9kwwzCo
MEuS7jp/BA0ICO4HA35Oo/I0gmWB6KyPzbuhQlwVUbBOut7aST/g1GvLgg/W
oDlWhgacBGhl3Q7OVW6ICNMqXy0iSl3UhwJ0y65uwhz/k/YIV2OjNlPGhOJa
Mr8mG/h0xLq34wu5PskmaGBbRU4gy2Xfsfz5yT6L5cLUk/PRJeA6DBoKXiOn
FSH0rlUtVUF4Qno+IRLPTHlpVBR/tspqeR25J9KkXIlFCdcWPT0WpeLYBmbI
qeQBeKjrHjXbxH+UP3cp143XHTkEm4ZvR/kVdH3nHme1bPhjg/Qto+Y942L3
5wShFc8GfaDs/RAPEOQRHSNnVVAI6bFmTf2hfbQcYKblCgw0xZOeFGh0JCyj
3hv9L9Q0qVPkv0+0loiOcNzbkmf9O2Fqi/a6JdFm14E67WnYnTs2l74RAfSK
Cq/lxsiUbfDypjeRtI9/JG7XEg8cMbuernkNGMPOtAXOEI8JJ7UhfOqgSmzY
zpr2DVTmLl4xjRtzhE8P973+oR3ZyW+vz50iUM5v42VY22tMh1Yrajzjhlgr
zk2vDCuQx3vh4Stwam1h7bbjespc5zxPPvrDonBgO0ICepJVJ5cjISHOBRjp
rwyXGG7W7WrVbl+cfWwJcA5JMvch8MMMdn4/zx/Ym0eqCZm8Z2KYJ4128hJt
sJMgBXn3VSJl8PjbiqyxkdL81XC8MU8AubB94F7udOG01Q5YanPNrdo0YLR1
u5WqOfEIVw50AOcRI6ceCw5jpYy+KX5HrHscFGENaqDAWerZj2S10mQau6Tv
k22J6Hua0g6ajQvcKvtKn9tjal9fC0OmqzAam9M9+P8gWGuOZBA6Bz+qERcm
V9EeZtsvLF7Mp6uJJfNapmuzyr22w7KMpUaJcLO1ZP6JookZo7xKDx5y/O4e
iUPnggUQ54BHflI1FsMGMwRcCgrcnaIN8//uafly9KdEA77PsQXKYpXq3Um1
NA3QdSB8SB5TU7ok98avfSsYMutfJATvKZjCd5ml9iQhlhKaYEkp+V6e1nwJ
gIC5lor6haRlVzVhzyWDXA1BeIRjd0yWfUTndKH2zlOwDn3NN6stguHqEW20
1FnQgEPzPd/IUWffaN5RRbe7gyzUb7bVYAzDrv7Hrwayn0v+8haMuCnTdJNZ
SKvIPoLaLkmGo6+F4u8Z6VwjV3m9jEUDa+C3SaHEjB8HKD+XjwJZI9h7zTKw
tlNpOGyWWQ0LEWnJqOTk3YZVmMilt7F9ppkXDVawDEeIQPRI6hN4AxZCU6lf
FiMPWDep5rPGuA3745I23X4n4Et24wY/2/Zbl1vVD9NylRjfi++Sbf+jYCcz
ttRIvgGGsNg4N5QiqZ80s9wGZTXZSeJd8coUojHGOtHDqEwfV4huLqOJGn67
s/wileuo6hITsREyM/fVdtJSONSfCQTHWKNEur0Jrn7PKEEG54LbRFoX0ZWV
5pLednayjXKr6mlbhN2Lo/oliN4s/iXBEt+YDOaDIOVD6NiNbJEGhFbOWUuK
QzbOAvjusTBE3Y324MzCxB5JjgW4AADrlhXTL1kIYoEVyx5o5qjHbAqADQB3
ppi0bL3fUpErAbXrZCeqHCoZzF5e0KzkIr6PbAotxCww0YfgW35oRg+V5ugD
mOIQbQUB+u9poP+Wt0hexcnpMhfxtY3zyi+m0bM/PBXB9bS3vN6M6vOfqLJe
sKU9aq95e8393hikElQkKAWZc2erN1oOvtXJyG2wTnZbCwhoP75hmf9KN9kh
2XWAPwJaZI63u4rPlEfN2SkxGg4YBamGMpP4Zb4AcbHk8DNTYODzsCVCrZuZ
zWJwdkEyvQ0dl4nc+FbwhI3hFrik/EvxopdXhhaFPZ2rM+PN7hENiT5vol2g
W7aOYW0l1Vs9SBWShXbt32nqFvEcWUw2F9UDsvB9BWGyVggT+eRVrGMr45FU
YcdUk7BI0RHoA4CiVUJJnIst1LBsGhpXqCqUDfeiVpirSBMxz+5qED7+VsPU
bu59TIBOD9gzpmSVbth/LgJLqRNV9L05XHSHofKo3G4v9m89h7pAJLAJQp7f
gdzmp1M9L24JE/fNfVT1Cztg4bV/lBqb7qCtUmXEDNF7FrS3VbL81Mtoe8T9
ZC33ot7fbk9zHssuxMg681Vzwr/ZoQPF8kvFc+dG4jtCWqnV4bUPBBvImFTu
N5q7AYC1S450bvN2WUaalCI71E6bJVueyq1+CziLXKjgz3r3ZL7dLc8bNsdS
QawsKD00qD59dWt7QUdjPlnKv2b9I6fJvXQTgGLBJEsEwQ6/gtLXqE2GHvli
NHZMI0V5UsXiIci067uhvvce2zqlD7zEmV8WUk4WBvRcFqCv5fX2ityEI8CD
EKiQun6cCNZSiG06dYoYGVf1HZB+jzw+c7dqYzyxas0k1GLv53TZnkRhWQun
GFB0egpmHp2ki5k++SRR/pd0lNZsOwtZbsZzJPni5qtmF9U6o1FisG91f/Cv
x4T3UflKKG0Mx85GBCssklMi/aDXgpGPSU73UP8IkXHMGUkWW4FueKtf0wtF
3wpEi81OBSNKUe+REmdVtDoXiefkPA2tUlzO3KgIg1nHNaTzNl2sKl2WV8AN
fBb+l9JAX+2E1QCV3aDSYGqvwoo1ffz/mjhyZMokgnbVeWmiNA0iEuBA3Gaz
pnaO+zXu0Hixi4jydDxxwHLySDopcQPQUa0HZPo7Xr4hBfzcZcIAJp9RDGRq
NIth61447HPk3P7VC3SkKKkZCiqVSmorKydUyWhkmExPij9eb95VGcHJgmQ7
G0H7CUNHSdgxcqfBj0buq5PUdzAKFqMCh0MtUUaBGtTfuYEpQivX5QCyF/sw
QbIM7H5st41Pp/GXvB0k4C6Hletq2gyay/0hHFMBDeg9fPeON9JiwytAA2dw
XMf2RM7RW0Tmf0TS926O1l/iJZxPHq84xzhn6ah1nmdrsy07OvITAH1pnSlt
oDxIEXMq5Qul00QioDaokl/inx/Kv9rxje1qYq0Knsq0AIKMx9w2Dii/VuGj
nzajO5DP8QO6X8mXnzzxcBAF3iRFXg5cceNsGtzUZOWtBFdSI+imBgoDFWdm
IGhOhAIXTbp5zswmnv0kEdc/tbQ2eBzErVHLXYGvysWB5v5s0v6u5Y9RHC6H
X/6wjckrwH31UPacko10ZAI241IeCYGsskB9BBmloZiXcm+DwTeh6glBiQh0
elaIP83W/3dCe6dxh2BG6TZxkF0Hp5RqgM6spQkaaT77omzo0C9fihfcBmvU
odS9lSA3cpkppKCUhflmM+aGw12XggqrJPRBDTPsX/loDy4YIqU9XX8o/3vW
ugvdMjOUUzD5MZ6RDiBzmcNwIyGu7WsuYIJ3a2tJPTqBdPFXM//25Nh1gr0R
uEJ/rxv69wCUTiq+SFoNrbqTyuxfmLjmb1E5ZnjBKkomsXm8wSfQQjTksRC3
UBdO80Q8/PfaBVV3U3jvNoAQIxv7jxoSLNYGfzbRK3IYwB8tEiaUNE3DYryA
ofYfOc8LhFQ9CJ0LW290zZW4ljALvTLdKcS+Xo+xyP4cCZ8J8p75/b+biI5S
CxbJqOVy1K0vu1gpdOyi7qzuJiGeaARPVGAD5Qnj4aYbx93zq9yGWrPHrmPf
iiesy5Ap3WuL/j0zy215IvcRo9rponIC1TPq2BY40jd52CVoqJOaZZ8oHZVs
/hpN06aIcrVCXt3CulJjcaAv8Oyqxh/5wht9M1JjHT68v0ezpD1LTmRgssBH
qy2gVuuuosj4gziypJE1a6fnYKTctKNcSaAaVU5ERhbx6EMwoL17m17PTo/u
zI8tOiwrUNK74e8tx0R8tR3y5maSll965K96TChTvJDm7LuYyNvdNGeQ2Gjm
5vPo1QE0BDWDTBSLObSKuqbJ6E00VVv0XOpOVALGOFD4s9M85L/u2OUy6zHc
cuyn+2V/WshvoSPOUO6dIabCE+PZIV0gke8GodKGK7Vc/ZIuU/3+mmkNXBDy
d0C5kg3IsHGvMj2mIBCVXz0KMUEQzckYV55JPnBIyUEbLwf0A6SRih01s3lF
Q7xek7hK+ioODtUD2viOUTgIM6/Pu9pMMTS9DAFqGi9pNB560w1+mMIcBsCE
Tf+I8XGLcG7GGZOMLylM6CaUJ2FrXCaRZi0ZSSPXGHzu66AyyIk8FswiMesP
yDI0cetC/Si1o8nV23SO6O9JBTkwQNZEQ6IbvP7NVYG3ueKBDS3Nx5gHfd4l
x/dW2teDpiIKyMjqGh920ncx5CtLBoiVcvMh7l0pzC9z6ZwZJ+U/iBJlMd57
uctvzBtpw9XI4scPqjqg0eeNBknBllrc6j9mmkOtzuMJhU/+FwJ5m3PxetLX
BZnIa4X4JMLfOG3Vf0stj5auI1bmfItaA4mtjlQAG6H0detE1rX7L7tTDz+v
/yPrJtnO6sIk1KvUlFv1irPu5IrYrPNnDsKHcPtB8EAzjaenGi9leRdd6feY
mgWFWmalZ7BvffWVCiALcLwo/Mh5dn1jtpjzqTKP4BMIWudMrHkRhTICUkPu
grdHhgTx57gF4r/u3dn8L2Zo/VKNVcW3Me3nW00E+4mfVoJzntGb2JNB5ZVm
lQwFGtNKbncCh+D9dxLbvk9R3OdI0M9ayeJ3Xqg4mo5W1exFzHFrFYS8e6gy
0TgnMVlzL4GfDfQCrf9vdIS2+O3mxfUqz+UMbdfqa5RPsRClDo8AAoVI8KmP
B6bMV51SpqV70DT40DTBhBNgshJbt0lbSSLh3yUUAdb4dsEaYOrTTncWCvMw
SQB6dpqGz7tsFeBUT9G6cUe5RNGsA1RkgLO2mRaa3KLZO8v4N4d7aV7khA9m
aXdEV6ScRsplqtkIrAAZVI/ot75J3sfDuzziz+wZtkeruLwpZsbH5A2fsNdW
Opieueph3Sn3PxWVVX2eoiUyScqds0jyhtBVTB9zs6k08gZ+K2bizJeJn40n
+4nS4OunxGbsOAMD2hbBsQcuM4rcwnkhOROXLLoYiZMM7lTHybc/IZOl/Ujk
AKyJWuv/aYg1kXjIr7edcEyc7L+ZZnLE9ZxfNZ0xCauUAIQIIAemY1SbQ3y4
p2op2z+aScSuWYnTRLjplqNwxvXW++iRXJCSbu7Spy3W83kNsvxUbbFYKpwZ
+D0imkFO+7upSJEJPc17SdlsqDFmmmnBqIioY7P2FMC0zq5dBZ06Mlh/00P+
LFHn4gij1RRud0KsQL21q3bFOX2XdsSUsrfREtIJ7mqSYMH47pbZSCYjClPt
ol+JQ006qFcKinj1yuLAS4XARR/xGlBzwO5eCK+tC1JRlq9oVMU5lpTqJW8O
s9h4GbCz6u00fLeVAs9wj2rIiSkUe5Ib5zTOp6qtf/ykZeVJ/r6491XgoWNP
HmlmXJ47MPLDLg5JIT3oVR7qNVRvRQKt7jR6beidjrmg94sZ0GD401PLoa/G
ZGoSOG/H1LQjsQe4JY/0PHWA5KYw6mi5zhM3twfvdpbOF+S6dYoAdU/SKr/7
bbjGBIVpNPJLLOdvNX/6WqG4meJdJGr91yNbgWlv88IdbCDkdGD/aGywDDWM
1Mi97/eJv8udmBbS+JrLQES4szOgeTerfvZnLxLSx0K3+NBG/VeGdZSh8U4X
Yfm1oVvVW+Og59mx83TKyNEO4rzA6bLeVkKm4BgZuQJbGoOg2ea9X9rYcCmt
12oikmefAwmtIGwVuZVCCXIzgmcQ1l9rhYM/qKLNb78m85FQyoRlbxo09D7b
BoTaDRQ/vcWxJb9fl5csnX+2/BohlvjhTLT41BSpoWzFlPtWYc/4GFHPA9Hb
FzzQsdjqRuIUIgFRxZMgr+f415y4x1cQMDThq268LIu2fKVNoRk6Gbcw9y31
mbdQZoim50i4nmh5DC36yTGV/2ajzDhSVAyQVRMLBepfOcZ2/pWgMBw+jjY8
PDxmGtrdZF2eOciGABhcX5fmhlFrocT/dbS7TEXJlyh0NQCvTVq5FQD09hkB
fgaB4KdCREO7N/QeFcTDFv8oIb6pKrwG8zQippwIAQafGfmXuts8xpHQ19y2
6mJC/f4BabWDCoHspjl28RhAAWKPfYRfx0icAq75F8lhcMWQAV7sN91hMvbh
24vV5g/pFwiTcJQAmA+0kKEg1k0gWufJ5VD7tgjuTu0StI/J57Cy8ZSH7ey3
SCKr9P6mnGfAqkhracQYOPcJsp1TqfzoVjqgjuUsFqh/4G2RhJgOlMklLKIq
e5121B0oqbEY3ZGv9PbyVUzxkYN7xkmDcdnd8vwICoA46JK7xeZLIpEZ7sOG
oPUFxQj2pw6szLbZ8av/TJExmuKoY45TFV2y2u6N+xj2uwFZtIQFkQCJtVr+
++uDf29T0rPsVY9xYmtuRNAiaU/iGw6S7XeWn+Gxdpo3r1HgoRbbf3BOA/Un
zrNiBOzjo2Z1ZbLwPQvHD9IB6UMi8nXyKDQxfAgpSbW1t5yhPHUCUOsFSnwK
IQyxBh4BqtH1Z9+GRWgQXwiwI/XyBJpMpOsFgpKFXCVyvzEZRegoXGVYSQu5
e0Qd0d01/B2GN4D3VX/yz6U5zQTd5uRiqbQ7wfgbFAvYjj9t7Bw0uf724pDC
PCoft9xhz17MXgqLY73zhab2dQcnE4zJ01t3qOMAEWNdHqnaLs2AX3zJjP6J
iy3ZAfbTrMH5Y/xEt+f0FEcTg1U9Muoxs77j7/Qh9izME++c8gg/jLQNV+ON
dHw73iHyrHJeGBu7KDid5GN6J0MFmkwfKKtWvz3qHYMRnX80XtKpcTv1+jJs
ytNBTyWNDPywD5nvzq5OqGA1sIX8oCkVqziRnWYaSDWAWxSTPnhqRrxy9wVy
EIW0YLg0n4mlTzQ7XLnfnGbjL/ST3VP8OO4NsHVWJEmMF9GRH216l75H4Z0w
GLX+OghQAuD3PBCZwPQv5629u2Tr3r/X4hthLaQeH0qsseA6S1MyJik/4Yz1
LZTthIAerB0vhH3WIHwe7Ldksl/YuRz0JnMXMbdfl1U5zftElBIvgeomVUiO
jyn54fVaZYTN2oixPB8pyP2fq+leb2fS217qGdfaxdV0JdKdoNP9CszDI4aJ
OYVd5EM98vItaWz2Idudnnn4f9JNKPtiyo9ystPeDET2cVpHNVX91ee0qzFT
iTmnuhD5PuGORcUsKMRog4Hx9D2n00XWn8JBmPxRTvjw3ZEEOJBFGNh0gmIR
LJLNTd3xeGL69S9xhpZJVtGoN2RDDUOL/TyLr32uRRSrj2KFSO1ZmLfukyTZ
lXOdn3vMneAzqwLaHr1OluNUgy7nwjxuDcJ87FuSrcS7UJEmQWlpY3rGSvpB
EuGNtOLMkBAksyGtuxtPAsdcZI9qONSmKd9rC4//vWzJY0+YcxusGlBx2Y/G
7234kqoxC8O1EFzVcGsz5DEJ0OWG5VQ7kAFMaeDR5glCCKop4DS8azE/lerS
l2kzy2fdI+CqcTOfuUU/7gUtAMyoThSFItj2sUN8CP7vZdOBvvcVzX7AgDgl
1zSUgXcdUVCcTjgUfClwxcLk34UIzWNeBtbzQoLdI0AMrEi5dvLamEqZzpwz
PdRJBwB/QU3Ki1sHOqIZ/vakcgsmwvqMsaF1YdGtekT3Kj+bzIA3aR+IPrs5
aex7xLUvkc2JAxUbOc7R16YjCfNcN73UuV5o2+kazKs5EkJ+PunJ2DsV+Edr
6/st9U7Ffnucey+aTOslTmUDdAKV0x5HDJoryMwk4+4vhQXcvROzn2r2OsZn
Yyjx1cuGJBgp26ZaSbXzMg0hUqYw70djyOMhSBM1o/yTIUbmyctbLhT1NP1e
s3aXLOD3pqe70d1o+v6vJlqOwVU2stGeVcomSdRwF3QH9upWjPGjIr12t76O
ckEYeFVA/CQCUcCZjijFKAzgD1WTF2f8qxaVoswR+J7VAJCNrG2wrkNtZOda
psqnpJH6oYpW6iPrzxpbqkXLwXzR1Q0OkIw5r58eVeve4kwYriW2sWO0UsG3
x5fdxAFywODmjqedF49uLFZNANHivz6BAHk64yaJymCFEtjOJ36SM1S2eicA
lPDwkHTaF/6yIQNKE7x6G9xYEG4QJ5ywrHJlgNm9JTrTAcPh34euVUWIfxcF
LR3GYtxrzMiXBdwaDVgqtXaQRt98J9xR19+qI6V3BUPPx2XbSZN4jKeVtr8k
Q7Af/14YntJzaiQJC56biNJL02H/RWRCEC+aC6vdaazdzSqm61hLNLpSPSKe
A1INwK4rUWWcjKXNDzuGUhAb46UyiPaPZGn1LTWnzpG8q2Gak5jL7G7x1Cwe
DZHZNi32j/7cc4Owhjzpl4biTXV6y6Wbnl07J+4ikF/dyyw3gBp0Ir1TzzFJ
4HePmR6FvTU+kG9+iSUV8KwpZ9OPm91GrK6zcP6iyac7FJuVd6zW/uXbNnFG
t8HmSiRpm4ocxlDxMq0YWNikN7WHARaIwk4bsIkgmZl8giwphDuole58tRxM
dk9q7ql1HDduxYY5FfEmmel144YGBOaJJjOtN4MJhwIFP0MCvBYFYAvTX/1v
jXA/518EKNR0hqEzpe7O3dpUzKTOKHZ6xmC8Jyp0P7Wq6Dt7tR2oXTcKzarC
erJgXoBKsyfQLV3TjAvVNbDBKYN+1NjkoEg1qkTcmYaMd/WMpnfzhYexRlpF
mNk+hSNg2HRbfFnC5LGsjBLnkRXIvr1v4vIps7aLsVgYnOSPGfDuasSGYFgm
yntn/w0re52ABQgPcrJt/PFvQRd1wi0q5iGcJtUWeZiakcPQcr8t21JPWTSS
DwXNlJSHKg8dN+xkLuonU4lPNYZveEE9PQWB1wY+qtN5ohFFdtYqaLC3Uc4y
Skoj06sGSX1BpI0BSDhGuOB4YhQ7poBHjW7JPLsQdsD/sZDJ1CfCYelHF0Qv
nNGN0uku8lsApf9M3abrRGu4973DSOYM+DEjvRk8Owbztm3/6KUSNS9pV4k7
wnh0F5i6VMaOxssgZBSy5lyQJgZ/K690tjHNRNxTkjJRsPIppduMYrwXnxco
+kKNhU5FDpQ5OPA4C9iEgP0ijzVBDC6fzYDEWbXXEYsQlU5GExVI4kqkhwvu
rg8JEtLcBE5Q8uareK7tT4OwNtHbt9MxkHX/kd+5hpIfr25kQkvrt1NdKjrI
RnNfYvQWL5rc1veI+EntW6LMiAEdmxF51aZIQHQEtrD67LUprg8cPF1E3NHL
Q75L7T/WFCC6+ESO7Z2Xe9+G7Tl5HgaH09vxtZrEbDOs9ztOjH/SUbVKJN8t
VtJAqIxdigWCfAR2Scci0i3XAfRZjHm1Ay72ATU+GaCFcY9hLPpxSNHKmctN
NZydPcGpGv8Op5Uc1/EeB15cSV74w8zbnuPzBDVHD3g8ISVm8LVvOeomZT/I
4z+KnjCB2fieLccJjfbP29+6dHI0IfhT1ptLcjeEM5QENTqq7B2OjfDFv410
C97DyJ2w8r43aWcFGhnBLBvzWcqS+GLvruXC+mH+ZFWyxED9Z86XjrZafgVy
tpm9Ve4P3KeExzQ6aUO9u539maJLZtpRmXVZmClWsuE5gtr4iP5Hh4abrgOS
TZVYVZMlPDKRXTZzlKEfLEuE64Gh3zdKLUSJ0RLZZ7vhbYTomm+/J5gKcFj9
cwl0bW44vLcoVrWb5RubV2G6dG5JoZYQMey4GifXkPfaqh46IrJbPz60QZiV
AcYXgY3cM7JThqA6lBkCWfrLrdLuZG0oQIhP0wGQBJ88PgekUmtcKy9NbJqI
xCHQ47Zv2FIkuqbKIiYPG2NU99I19An8tljgpUc6nveZ+TUqViPXl96QsyD+
GuvF5jWU9xiNVl5Dq4zTDQnamyGjSziPqt+Mbjyrm5DPbNwBnY2sH+ZLvoIy
UKPMl5Rr/MekHMihlVaej3E0mI1FGbFxK0XhD8bmp9IfyJUO115/ZSNXmIZJ
PxUyiE4b82N1Ju/KQNbNrPso22Qnuu3wtM/6WDetAdsT17HGopI+0kKxMcmV
/L6xknH9isHqVzF79JPNNLoyaV4QV38ZVLYCiCXnZCFWD1APtLmZm0D0recC
WCyNzrEe5Db3j+g+XtOHoELdDO+dNe66R7ZqRit578YItiafkl7H7X3uAfBv
QD+kx0XqNJwZgDAiMPUx9qRpaRsUqkv6gI8SNfum9P2uLdBfvs6yfb5GTymO
gyHjoXSFCtVdp2mzbME0/t5OZEkSFMT6ysowKtjywwNLuu74oyK5AK2EGn6z
1SEVnm+GVmYY0t5DskoxKT0/R+s/lTinNHfo0fklF8t06qI+46SGibYe6eXE
rAHSQtnlE2cith+sYkoPuGbhiCBboqGJ5nD9v/UPy8HoBbg6F/G9GZaGXFOE
KzUpy4PDcCnF2o+/2b7/ENvvpwLWpzYrl0kEQdkgglOjrYw/1hgs5yhugn/x
7ur/oEvSAMURV/+OjxSQXTd29n3LrMpLTEi7SxhWZouc6JB2kQnNovgQFoPJ
HqMc9OoVdQAuzK/sQ9UnagYknNC9kikj+JPvhuMxNB+xK5w3FJLfHJ4OScp8
XZ2RGI+d9Tdr0Ze+478l8QPur9OSRUXntfovKoIYIF0LG2/8yqxZP4Bq+79U
R5pvuzNt2VxtiRB0jZDksqk/dDb7S1g1EVSZXFLkjU55nExq+ng2wXbFHjkx
Zen++l4hRChT7aKRtbrj2JAu8bOwQd8PxEF6Cdum/9lqW+iApW6sAW4tL1gE
5CzKEL28llsO9J4/NLnvlT7dxB31uObK9vKIsYpjeIdpK5LHWGDdP99j5uEx
9At2L0TKjHAjJ2I3r2tkxggSxRGn8h9wM9HmDl9iuVRd4uZsyXofh2nvKyzs
AlvQF+Hdpo8MqxpHpwXPunIp82lYQ+N7gr0EZUhihlgDZ5wsaewjOxII4tPL
GQ8w62NQmj0UqiE3bMVmuBjan8+IUczkYnqEQzzpMlbWm0lMIdVjp/oP31im
v4h9D0RnkhJ0Bg6DKTpbIoB78jnHvsl/ZIaU9kb6X7m9rubViHIjpjbcpo5K
mB5jbeiCh7YcYBliuaD4RkhyedDgwTFqzB5qnFavTJnNLIcEycdXe9nmoc4o
r6wClDbOJbITzEqHiFeWmt//kfA521t+pRV2GR1OlzVfecNCm+lbMdU+SLEm
vrCyGNvF3e2x1ugE/RKbxqY2uEGUMeaaH9vjHUJauZnQxnOFiLDrqdAhH1ro
LtlA6co/FNKpp5TvrlSfzBS/KYoF6RM1qFMvEeuUaVGB+DNsZhljSId6h+cL
qX+MC73hJ18KvxTKiSrblsRL4IOssGBMzQlGXiIv5GEHt60YMPV45fFGV/Zz
YovGyeLGywkKnMFz1fleqbOUiYh6QwM4kYexf6+5BC3ka6hjPp8kjcFpjdzT
wrtxNZ+zUj37iwUe7XK2pElwi5oNokdwLYHdNX4iHjIjvLGevXRWW235MZg6
3JEasHUDjrDZWDghU/Rwa8UWCc+bfGXGR1ncBhS49tscx8rihCDgQenwzSN+
Tx9yCyufKOPmLmjSVcA0vLLir0d1y7o7ODhFXIrpRhHZkHUHvWWWIiLk24IX
su/oiDAzBFt7tXxJaX3e25eLi/1l9tIcMi/j+CnmQq77wAr6KNoMfb1S8jgF
qro5Gf0k/NYkgwm79cHT0yuqTO8xXoWiiLBV0N8g9sF/TtTJG5FSq3ZmuBmd
fSLNlSd6/uTjKLF3T7lrSlbPqACjCSiBEJXOtaxsU1r7tGnycVu/0fbqP+4E
jM2eEQA+ssaA48fjr+VoOIcVv0FzeMDA3L5PP3ATI7uuRz1QXy/gH2gv05Pf
ZiCF2tVTMVK7iFORsym/a/8A/gYgp+/uK0BIqBeQrZwbKiamYvwaZ3ayEoFu
1eGKaEkhN/qx2dCmwzYfk9Fz+UO3CiH8u10Az4HQ5bnK4yQ3XvnqlNgcmfIZ
zn1WTZ86utjQUS5ns+b8CU15HIMgonjczEWGC2nAUsZ0yEmUZSeSIX2GQ2tT
OwSpq0F1sLcY0uYKZDxpeXgPpxVjoNZErdWl2+WLDxJmA7hxql1dEqY2S81Q
hCqtntTzRoIa2RZp/hyrJii++68DYstfRkDVF+TtNiU9P2duH7v/erVyCEKj
vdRmH/3LWsZEBqBlKV3lrj7cqattMo//FTqiLUz/WW4NH+AeXNtiEsX8b6EC
vFp/73GiuyxwJn2vcfHOF1iVBdUPiFxqJnZl+U4MDb67YCujovzSFgbSEDAd
tki9+8xrz4HdDdqZVIjj7ooxLoK5a1Wz/em9jC9d38vhEP10ANY70tY1Pl0c
eFmX7GH3l6b6L8xcs2hy30xvrPD1D3JFeq+OIQYpdutgq/J1aRZEO6kOAHI+
jKy+eBYg5cKVC+2zGJ2it4L/yUtrt3M7xIXZBmkq2rwt58sigQ6VmStGbUIV
YTIQnBwLK4JplDc0d8TVvzqAUbmo3yBgEo4e/x1b6eAZzkZ4wpR76HdUTuMP
KKPx1GH/ZZLLqS5L8+YdGlkDmX7NTBpDa4KnOvlZ1/ftWyLZ5Tiwb33NLCaS
cN64Bte9HE4ABB9yyHWlKPZ6P2+jAdj3UzetQ674pKmsqHXZmByqmuo0klYU
AXtIpczLDz/praFZyUMeN79pBkbAF63zo9QuE8bmjzIcVQZXy6Fu6cHjfP61
1koeuvJHzsyEQ7zwJnOzwzrsbtlIA+Chddeh7x7b7E2E4aovK1fLmPt1uY1q
ss1vyTTXAIpvq/By2E9SFizFGUqZMeR0Sp3p0N45pQphiWuiJUEc70iTlHf5
adsB1E5AqlcGD4wuu8iSe4+3hlHqzbD3z9QOOmEKikYGZNoOoQTxmckJKDVy
H/IHVeeKwC1FElEDHjIszAvCI9aPjAznUFgIEqZsbfkBYBqYHplx971GqpVR
MAOI4AEWkKwW66NcThEEHDa9Sd9D5+AjAqugB9O/5BoV/jzCG7qLbZAk7orJ
K2Mu2ZeEAohFkxC9CsFgVIQp5KUNf+VR5TYmwYHbZc/8YDKpslKy4TqPCdJT
t7Ck8cxL6P1wM/c9rwBt1iF2zeUUNEi96ZFAgbzV/VMTKYaTGUidD2e1k3OE
8+2QVpQyqluB4QYx79jRmSl6sHb6M1ZCqDcIQ7Ih+imb4qKJZD9Xhea9ZvOf
ePDxLaOOqg1wc00m6lswvcjvpHpCP2O7Ml/Lf0ZZ0Obh5BE++KU7+nxwVPC1
nY5yxoOf+qDoNg4CpMZ9fV2poG2Mp3IGpNtx/dzoebzSptl1JlM7crcKrXYo
9K029k4+lTQWxWRx71ZPf96Dtz8T08pa9E3b7uCAq/ry13cy2w0bKvf7JI+l
rz0ygIqA4HCI3X92g/AUCefMANhhVGz+o4unGnBuaFQKhUmHvbabE4TK6Gju
bCrdhpMc7MdtFx1h2SfMKxtFV+9nh+PV8lhA56rqFFgs+e0ySeGX8Lmeaji9
KZv/t7GbXbi/MS91aCLb9p8aDQ2ncYZ0Mk1vvinhM7ksOmJJfYlTwhTxAUGW
kg5TS+BeJBPLH1Y0yv9rZMKkg57sgf9Gc4UZjTKeKZiwR/htXW2FwuPbcz6k
76T6OXzugLV+HOmmNCYE6Li+GhnL0LiWyxRdxewA60ik+B7ZUDuBS9lHQhJs
8YKjVWntTLnq+D5stgR7ZxustDb/TK6x5243YtZmhlnJuXnkVKxRRmhlO1rQ
yyqdaqIrOCwy4BTnd4yiMBDFMz9iBrVmeQXyY5BEtJ1pmSIwYwjTST+nf57N
F8Qb2K48+3G1nYbIOQlPFW9ALk8yQTv+Bm9HIUrwspYzg0iqw7B6zE3SnnRj
Nz6acqa6/jrsVHZ80wLPz/cwmrhp0UKe6Jv6rj4RAbAxJW7EzWuIvHB4CvuJ
m2gQQr2ulxSWUm98aU+ti060L7Gh6iAn4fxK8RiPXDmGVu8sGEMhPO5/pVDg
WVYZSiqih0plNmSmxbqd/MoHjh70rfHTweD1JmvOdlKAm3R1yZZcRkpJlxU+
8RvxsBnrgHtIrqdfKCMrpny8fWxJkfTkSqSV23gPIGIeHz9oe0ul0fHbdXQF
zb97vAeMpO0COhbXuErFaMcYaDgwk8EI1wKL54vMcu+iKUFnSBLyQRo3dDMF
eI1T14M+euy1sm0GOwbUCabc33dTQ3mcy8UE9OksV1y4Ho9zCPVrjJ/lvq+a
tLf7BT4yAdPe7ayJSeACltIMepodur5+XkGzojK/tgv2Y08ilnLFi0lrsVtK
zgfeUymQE+9F7xsqlQGPNK/xmoxBg2hhW8r50KgcOg39iX4CMkeTypN4cZnM
OAsv9bdcfOdyGrm/tKTaak6sQPhFmsTdKaQNpTcqGisuQrFfriLzYW/q98uc
DZNugIaVwbVT/f8u22MvEAmPUGhy8Nc6wvAioM1NcZTeqcj2r9EkWbGqIwCE
rssDhEKthigHN74//TO9giK6PH6VTh+SDU/vl3itYJoZ7fbpFX1wO84rIvxt
L1J24550+oJcDaSKyfVKa1f9ozYaKpV/NurydJ5LJruTjkFvapsZOk0oGphV
1xytnwAGQyqh+pym1T+w7LGLxTqnLKrGvnaz/7tF7Ql5Q2rmbmuFoUjqGghc
ozUb9Oq2ozhpKw/2QCSXmJhgd18SGgzsFpKOE2E3eZenzHZt/KGxfMu5u8jh
o2/ubgpuo6WI14mkPCjBp/TVEBuO9MQncG9m7fpYejV5xGpNu5ZzqbrLbh7j
Q1pQyWA8i9jEEi0xzSs5DPnuFT6W+qqDYuix400OHLw08jy8L9+2EKPV9N8E
dwzl7yn+B/e7wD4gU0yjdO15fRXzl/CSur3ygTJtb3XPlnSC5aYi2m4vt0JF
1uPCrZhLJP+ShEBDizcoCIXnI5R8ZjFJFB+KGU5ybe0zEwTBWVFHoDbu0gNG
mgteJ1BhgXFzTchjNPceN6cqyaV6ZywLWfojY0PQjNV4Kxt7tP08uoahDx1s
vtGlstzelkE5I1qGz1e4y3O1OZSyKtxBp6D+GvHuc/TgmYFgsMtpa8znnH9+
aqAhbD2gloO05PvXvCiqePkpz4QgIdeTm+QiUGAm+aiByjkx/YotlKeE649Y
Te7P8u7EFaRQqAoUbNJxRechGmQxumpH0AchGDF7rJ6LyiQFO9qWxxYUJj+w
r9C54TXnfmvoMJOpGGAiXBIKTznBbphhty904+HbSrP2XIXZtMFmhpJEoHbZ
0KmuSwlKHQV1dr31WeoB6/29VcXUQnA2jTgzIQmNzAbkI3NjJZD+kQ43oOhW
pbxlOG/70B2u2WLgCeN5QQSKJ4X9uWMcY2u3VeV3p/J+fySazjDGbC8OUGfQ
AZcpkaT9RR4a9UEfxt++LhWKWavmXJnr8mco5OtjPyaw77GrLChH7gQZgIpF
CqbKvNyx/meeMli1jK3u5EftG3zZu8d2e0J5RBFF2BCfS7t/m56S2hkLhpm1
TWOc3QpdNIHWK7AZlDTTw6CEZ63dtlsuvol6K+rFR1lVfFXiCgIOZxTL4kEW
LUO1+KMqUaUgDmioG3DBrfXX5KY32shox3w5o9SKkKI/b9EcGZTfRUztEmNg
X6jEYoQl+udY4DSBUKJfm5GAOpWKzh3P9aAozbAmlwttb7gc7MYVcv/nQc07
Bq/U5l/8WuRW0AJ2EF2FIVIRCx+YTAO2iBluI0bPF7Mkg7TEyURF3FttpZNx
lvVaB1wBxaH1H4cMQNbTs1+8cmo0Otdw1ECQiyEzGGRIRzUO4Pr1K9yukSuh
rJV1MOYhYukjChfJMNyLwAdXf3wPx0lYuJGsz7M6UQu8W+KzUupaHv4eoobJ
Auy5MyS5/yct1LVMCwK8vYqa/mUeqeCOX9Ctk6UIOaC+AHYQaw25lOjFJYDc
D5Ns5X9OfiQ5zHRLQfbe2lAdJzzHplwxAggN0MQ2Ij1rmPRJ9vyfOEIQTfbM
iqdgOQhw2rYBQJ4BAeewBLVNH181sl2CKDRSYk+sbtH6f3KlkiyWgP+9UDk5
wf2n/a/T421yG/+FMzqb95apRCIiBNkT/aT0STDfzxTJCaEllqHPqGxcEOMh
lrs3NgfmncLld1oMxIHIZGSJF6gKu8tnade/45G5kyCBj6ncS2jzGFgIkUw/
rAHjksu0JjeGUQz75xZKVaQy1eopzBAoEJbDW+73ezdo50KeNr6wzsoK6cQr
RJSZvq+0PyTo0zzJB/1q/wemD3ghSApQi7EI4dUH77HbEd2O2CnlfYf0WwV5
bEW5uCt0QCwaHSczl10eMpmyA84i0eXZ/seUcgV8NNIlKJ+XotWpnxVQYnnY
/yM3655BTAdZaVQLHlNJQSBj3XgOf9S1UY3gYQeDu29kAAhTDGawkUIahY1G
WwKOgfZRvV4LEmaJ8wtlhw8Z1+xy0eIRR42LwcQs6VKh1Al12sESo3V8ojvY
ulfnXGA5WI1to2bIAlet/yAngJG8/aRyj7xYqZvY536s3YaOhBk9gUObrlCe
EgK/VpSTr93OYJsbzLgLZUUsnsrHgr7JHErlfyyjyKv80y+nLIQ5O1buTBJd
naiWEkP0fXuZgzYyhfy1lW8yDvoenU4NZ9SPHXQAWrtRkmLccj7rsLmmZ7E3
oEXr1e3Nw2AEgdmtdr6LzdhYFxqNGp1xj4zQy2ClfFa+GajXAZw+QtgKUo1x
PH374BHohzs8s+ocv/ynqEzxWShyReNfqQEJ/TenL9pglzK0wBs7i4eaMWyH
/cttl792GLH54HDw/ewdglAjzQubM2HqSJ6z+KOXDw67gMkedYklxN/QSSta
1wVb2yunuGb2ohMLQI7XhfAiPULhDSfvASU9qLmX3W7aKG7uJZKqnurpsvZL
6ZXdRmzJB2J76vTPrPib75VTlU/GqVI4kz6yCOAaxMltJZj5RarnZVUHaef/
cauj+T4zwAeWX5VpbUmPVK/3ipLROb/3S+jtQsQGPGCB5wcqEIu8oEkBR5Qm
1jsaVGHQwuHI3vc37V5LxEroSxN8C4JUKECOsj26lVSq9YuD285sNP44A84b
mfKO7WpBt3GMDxjXP2Amv/qAvB06nmdNOZFDiYe0jT+fI1Nnty8Iccjc19KD
Ja4coBPg2j2fY6Ka02Gi9GFayAq2FizYKf0Md03qmUm/1VKgCT7scnjO+5o+
zcth7sHdPvzlAzL+jQI+2lc+Gjjbn23Nz/O61YL7anLSlZmBhA9rf0MJNXxU
UeBS5eixE6ptZ1ZggZll/vPsw2Z6wrEvXZm1FEV412guyNbembRunzvd/X2j
b/KdLK2yM07rnAaZ8yN1eLbjuFLHJHTiA3WDfbtUg7BE9sx77+PhZo4UvTo2
rUIwpU00g4wqJFr2//WY9x4F0IIL2KDZpY7kx4I4RjBgLY6qF9Ume4rzhWo/
fGIt1NkKuMi+9diCHKSFZ8AAc01o7abvn8uXQGpymdO739V2WrkBjnUuq3VU
Mcye41ipQXsL0kv70XbWpKWHNTq4dxr41sfzV6rt2iG3lLHYmAt7lyaYjei6
wdC404giiyrNfir2UlDu312GZTJl/sSwMjzR6r+Jjstr8qWuU//IO+4svE1d
WyeWL/cV/C+QF1s+IbI4DGAOkAeb7xQ/DjElfSBgvQi0fyHi2FR6eQVx2gJQ
od6uvtoQCjGM5GytU6Vzm7fgt9q+YvsmqBF5NahcHNfc2HXLFCavwA/jvM7L
Jwo+iS9+qLBjU7a/Sk8uH1WQ83Kzh/lihTOkf8A+3Eou8F0t+dv6oq7RfpfC
kvIki53uYAkX/a5uRvkpTiyIdlPvu5NLbEd/I3jT1Eng/DWr0Wq5r1oMWC1K
FZVDVkYJB6/DtlE30BGeCNbXKhZ83pPgqYFstKoD7DZOFPl/8Ctmek0/wEvx
ZfVPk0GFXN5t/r12w8LBU6n+SuS004Wr57TNSw3hHhKaH9txTgVk0H5VsoSC
Kw/Q6PWDYg52mAA3E5R7feKEIm76eVBUDxhDjJbouiVcFqwwqwAYd5Rwd8w0
t4PYSiqC4d+idY6vf4lRDbfCRY7yxY7FClMbb1U7S1bLAUoN6zkLnWdWnKJs
HwArTQ1yZVC3qATZL2Y9+I0sIrPt+ohmZI8WmMcK2jPdbB8aHk3xuh924eeX
NM8Et/oE7EJLtQRUl3zUrVrC7Hb/VPZRIUP0HKHMqvDerUL/RPEyiB/LxgOu
dCYq00rio9F/GjIJKf4nhxJSieSaUXwPW0upXPeHBisSVyiWPaT4rJsLuxBp
fXOu73RirudB4Nn9hoKRK9o9R+f3X9bNSnKI/PpK8jP5Rh4iVS8NvGCu2dZd
1Dhw58aEGjbLMyhyeX7UQVQHzbGQHRZnT6IghQ6trEUQftcaRPMymsfYxCwy
h1nutxXhMC7oISMz0FHVFmJmWJTOjofBVvx+0A9IxOMlhe////+K+ItZ/gF5
593ihRtDKeN7IpHA/kXkZX8Zk2ae1MhBdTdBAKfsWgY8uoGagbyT3Dr6mgqN
RcUgdFtA9aaOfvekSIkL/j93KASorAf01pv1yTK42Sdzi1SUsQJcJKD9f9Bq
PXF5l2dM4eNeDqDcbC9qAvApX0VLgiCj4M0woCh5yjYXH1IswqE7ouulNumI
bqLVc6/SHALZjsK4QA1MAwWOmxije1HwGQsU+H8hNGQ4mpooSRcXu9zgxC2k
ITRcoCqISJXXiDlV6Dl+nKTD8B06va51KhntBItEezghqcoPxZmPqjjvEEVe
7nEjiadlu6qUEW+CBsex+YBmdLANUBIK6CdE7chl/PLQdBgTiYlWv4i7nCXl
8KYRWCP1AI+N1Y72WbYuI8gAff+3FPU3HYX6827YHCT2nYBP7vjT9DPTC0LA
qCKSJwGCZfu4k5XTl2eNHECQYBaQmlIdblNyxfLxJtizWRlOaApRfWUZdxF0
olOmxXmK1cmLSIVQhtgZU8pYcu29JOabIvx2wkCUgyy9Igyr6rY3dbz5eQiu
XdvGoNBrI/VZvyM3i1toz4jPYqnIJ9ccjDWuhxKGovcoytk8XM/Tfy1SbD8y
9DeDl+MXdDZ5m4slMwl81Dk73CrQ2QqwBhOjBp5IQTf7DxhAIwjSm9somfsn
kp3Vu16CaHgm6Sc+RPa7qyQAEgQ+MRFpj/VqDlUekPLzZRdqw8WZcglosQCH
i3qJzJId8uKN6onfFrviBIqCHZ3OAMMLxWs3+JrJdoBtaIPKDv0BMK9GPp1K
C6mX7Ak9Dd2KwzHMbJ/e4Qic6pOId3IjxOOs/FwpXHMAxkW55qdBpUI60c+e
a2l5Rjgn3Uzd7AMo6zAgQdKuyX2mYi7Zi8SiDrJE6XBQA++BGQDYd3umPeU2
ySHxGrzcQL4mdZ+EF140oC4uKKxK13/NuFNugnsnxBc1oPFePooZeJK0HLyA
7wr10wC3jcQE8w4UTxtVbydsHXa+jAobDxGNm9cs5d0qu0uC0yHK1OT0tD0t
ASoEq7k1SIueWltOokMChEBJmGjDser83+SPE92IhjGZt6gUJwebX56NoULj
TrOQG1pIWJTVdwedyzewVT9ScAvcuDCuowhD6h1Hw1cO5Wa76Tdod8VDj4ZA
N20zYm4cNvguDFtULwoYaLTK6QugObaAtyybX01W22qNut8nmdV1XZw37EeT
3xu0wXEjYD0Ijkz/ArMGpdOkjGKXuo4poY2l+8TeaC9S4jN6ijAko45gdCmt
8iKblOval5vJulyzP/FWRgWTl/K02Yz0xnuu2LIr5iLlf4DSEgbgRdk5aU1t
/1o4pVHhXL6SsmUUjeWm593JQRgx3hg1gC//pUn1wEMhyaLBkCBjWs3VE4hK
WtTJp2JNo7Onm+I9aW912wBRjW/ohSdki9tqPy8WIxdh4YSi9odSWSrK2Ws0
IhZarG0jyQFse0x7+tC4OSqQzb9X3R+KxdS9DX5tL1NZobukYXtdBM2GJVxc
dts6lEvBu9rPxiFaLzy8kPxZlYNU4ElGDNyBd1uBwDTcfWAKA3HXQWME3s9K
LYZCPjOfNbs18D+5895wPt/7hOZU/0jNK6LlQB8HamcyqAVtviLSr+O+peA0
HryA1af7AR5bE/98LsF0mOcnJKSLN8Apc/IHmFnnBqYQQ17cF0Kb83/M4+Uz
/C5Ch/4Rpfu5cqF7UOz19KWL2TqFgS2JzWTJIyvyVn/1HR2m/DoFP4CN2jVD
Ayi9Uk5hMuLyf5mbN/Vz+XfOt+RjZOdkjCZswv9a5a9QpeKRJtjezmQeKFnT
bXx/tH5FvE+Unw2ITWpWo/odFibNutjgBzVdgWm9IjRdDPgIKKuM1I/CW4g0
J+F8Fx5jwxh3N2rEyhZycAu10SXzOVUSIysDH2ftFcTzPO8Pfe+oeqDP15nv
HoJ9oQ5lwVmwWRkuXmehccMIuTzGBWpohLDbYVRhgPdnloW0ECCNYl5Xqgu4
r3XGE6VxceMlJ1R5LDNfz4maqkMVd++uwu0tO9pz8U5hhJGyHLjy79TlkWmr
vIfGmfsk32ca5tl1FspeTqkoPASWQQ884Zi2Lqab9awUKg4U0pNCs/H6es9F
0u3Wnio5XViE3HkV4r08N0KCQXMdeTaecds1dnbClgo4/7aXsUEmc3Jbl0Um
5rMF7jbDZQUpn0edFyLY1nVhJ4k7nN3xUfAzgs2S8my90szt/gvdZiHgla91
s5z9FdcRl0+zPPARwuQ3V3HHM/Jwyf5IHkAY1g10AStqRPPd6/qPw16Y5veC
SKH6R2Po6rox2q4/TzcaQr1De0JVhrV+RsnezOP/j+6xrGmIzjlShjtQri8E
+oJAqQJqIjBtvlpjfLzyLD/x7AVF1QoeXvkl1SvKCPxefe3Df6ygo/8HmqiI
vuIAFbA1wDlymQB2k1liCroo8To0O5i9nef6hYY3MmLpWYBbIHijfBThgeVF
mXe8MikRzLyuOZRH6FK2Jvo7MEbAwD2SIWebGmtiVeCFl3z5ozxLHCbHglKv
52/h2yUFkI84h9Gzrb+gTyoTS+6mFopE4shaTy9K0zgRo2GC16jnk9ZH64zR
OPzjgN8RDPKsewua/l9ZaeSs4IMAfoowhs5IuEYvPAlXhPsAkp2XjCYZuvQH
+QLowUFFNPKyuCI3tEfO8q+qdGqY1/8jX9bQx3rvl1uK3OaTDzHzziowchbT
kuIrZOzbbOj4GsiVejMevszDhQlzm79CsIHoPGQCv7tINW1NgG8sK4FCR4tr
qBiuvoJ+J/UqzMhiqdXDAgGFiXSDH85KX+yD8Xa0T5j3Yz931rH/tSNIPl4t
ujBOaE/RP3WGODhZBG8uOz7kVXiwHLUSje1O4KCay+NEI/8wt5BMKyoH2fZj
ktnybJZhsSbLRNedUDTaJijcke8cBKF8nzEI5AJd68bxKm+6jDkeJa/GDSCZ
edyT2D3J5UkN9cVdtrVH5ek8twzXVGfE28BRnLbpXCVkNoAMYDjmDiyHVE6+
dr3CX5+qxvsajSCMUZ9s+QEFQPuETcvJhqpKl6HvbWlntI/NMh+IuLH+2mY3
Z2lDIn4wNxeCrTkdrr4mlZH+xWLCceg4shPtZzNbdXH02k5gCrDspNDCJsfv
RyFHjZHygK7vnzv390j2zSeu6YHJ6YyI8UsGclQefvnVjDVB9YFhhlSqh4Zf
ylgwWzAsU8ldBACfVvcaQICnx4UElwL43up7Edn1nBcrOvMOeSwoosf8Z47I
9KPZ5hnTRXrUZBV7TXsXmGZIhVeS7J6aQcpqruDoyYuQHT0TY3c9LE1khTto
F2BebStEOEeh3sIdsGyn7LR5lqgBArhiuAWTSSeInTbuCxEYds1T84SZ/zFD
WJFkfLEluRX6V/x+0MJTxv46JHyhh1zqd0QipXTwfpWZOG/EQYYPdlqWH8nw
p6woQ/BqonrDOmYudi+QeaxGPXXaVkulxYdr2OaXs/dfoz4fp7V7lhTbvIXY
hZD0UKDTU5+olkOl6n01ESQG6J9/DbFlbw3y4Av7sjAtf6q8qD1OC73Jjib0
rXeMoxPmIA4L21iaHpxaaE+kBBIa8A5+J1q+NNjNHz7XkNeEGN+SgVForiTY
UkYXZ+lkPzv/eX/xVOG2GkxL+Z8N5yk+ftNTI8ALN5hwG3vEzBb7JRNRNewi
bc+UTp6Lk3IOxnb8xkTpSlB5Fiff5l6pKrpkMvK8v6z5RoFcnXvt8vJMyOVe
g4y2vEYEX0t/s3oiBNh23gt5t9IIC+/kbKWLd5rOd+AUDWwXI6zNu72b2fZ5
BWx+XgM5ESO1pek4e3n+sxUly4Czg9xfvf1f9qlj6Mjs1em0RAoLJvD0wEVQ
TGB5RL9YpqUISqAEnDmz9mRq8LdOOi8M40gefv+1gF82mm7+pguYPqA6m3I7
AItrRtIcsDIBrkPaT4DuR5gwqNzT5eBGi3r5627suckqxAZOH88IfrNe6dfW
d9h2qxzXrZlJbvxEhhhkBFLvgZ4NaTPqo+hsZxH1IAJvlR5Ig2fd3IQz8Nec
KzO+H0dL25QDTpyn2vW2RbABflKUABAOCJfEPhvWKr3wTKUIeEKjYHdJ+jkk
kJiTFjIUOutAucjWgdKOfjGQ2kyVPXuWq2F3fCtrMtyoYHSQrYCnrvLU+OYj
Ac/VMpIFcL/vGMP7IB3cUSHSEaLZSnWjLnrrxdgh2hvzkUCBM61C8bNZbtwW
XpfLT3BT1vO0BB0usU8nu08mEUzucUX2XP3xBdmwmDMUJ9v2QYzK1wzzTAYg
SoQW2D1oe8zVdsPbBNXDIPAYbpbPLTiLoTIDFh4T70mf7l44sRK5X2g/0XwH
Svz0oTho8Yuz0SoJvK0+h0NmnPqXJoWMDnReA/m4eDK+0L+gRBRb5xDXOK1d
YCpGJYeuJLRNAhqucYpTdvm2KbV+ES9m/6VmLkRUAsDX1M8piAhJJlkH/qnW
5nUdbUL28LuUfThFO8dcuARWeihTZpT/PM0rV40Uh2uRVxcPPzptQfpq08nv
OcyG3VHsrgblYsoZcA3/t7vA1NI9ajZfAgsEVnhirnv8HEPpenRWPNp+ShG4
A9sTa4jl8mv9ocJDO8rWwv9Dh3/vexw+8SlQ05co9IeK3RHU87bCkI2NpwFf
dDHok1smD8L/SdI1+Zv0WqKjytSlQoKoyMyILW9iIt4wyTWkOp4uZpwoFQ32
S1TGBxb4wGmZQt7y6dc3blOP+ZkzNQnibqPBYd8hE8k1JYyhF/AZVKpyCKN1
8rONwAQjUQyVFOLJP0ep08toyJirtNe97hiCBJtZTBAdLz3SiYZznGkP+sRg
Kvu/MjYFN8sVp/B9s7Mr7Fnn/PE5Au++g27nUUeBcg4hMq2XLxCh6cyUly/q
xcKBzmPsFRFhiSs28nIWj/jworgP1moiQ4vokQSm/1SO0OnGGkGbdOtmSXZ2
aPa4N9X9qnGnz6UAodElVuj7wzVRzqPQb75sf/03MeJ/z9VdMnIPiY4yFlET
5H8/g/fJH7BKM1tw7S0/JL+eV4thO7u7Vyepw+k9XfsUz48d8Q3f4Cs2t5qd
ZX0FRBMYZeIWarQvWWs/aVWSv3Fuk/ol59ggJo91H7Gr26CNhqcC2t7Q4UHU
weKUg0ijN/3zL3iOBIUNaQk66IXtoByeEvVXzxtdWD3EvtXg0SrilQ8drWmB
NzKnCyXG2aeVOfc2foOPBTfp7xg+t5kwjHhUEUMTQE5OpdmfQTpRPdfRKt/y
BE2hP9nZhHN+nFrLaidiCHhnDCXtjVY/buGShCRQ+scGHenb3EgrAW9SW2I5
DtjrC9QF1BGnPc6Ba5bbhjG4YuudDc6mLBPajtZ3SNi+uOl+UFRGtua61DBw
7BModF/3bZmq2WRFIw8PBmHFrlPjKrLPHzJSV1T5NWugrC1JxcSsQTiVbUjS
Lep8B5nFlweRVcdLBYpy6A27fWs8R3+AM568WPgh/Khii/Y7BkephCFxmESr
KwlzdZpJQqmgpB7EYsZeH8mL5luAtg4Yrl2wHY/1CDj74IvtV07q5PgTbCBd
n7Hd68CPQsxhgb5e0H5mA0gEsoL6gAwb+XsbEbmMTd37tXjvaUU4jkrTS4zD
xal3cwzyz0hB2/TEQnigodKwmtBScvL1O9b72tIhLFtrcGRUHrkaSNUBkGnw
Q7B4wljQkqfrpWYCuqcsMEQVnM+UOzyFPyaZeCOiIVCAsXpUhwTfgokD0sfU
MEzG2mey3TWC4sdKzb1akPOhqZILNaY9lyHTlVx1ICYb8q17InQxQJllsN5S
xGK+Sw9X3Kab+m+086piTHOSfeVQGYqpmnZp2iU0/U98r0Pnb+HJFQsY2v6A
+OQsTAqrN0ENV1kCzPxoPLdvRHqdfvGCb8eVw2HoEBQzJmjGr0QCxlkCpZ3a
QTlQlkDdPp+0iU8odBkT1Sx8XM7VVoymvZpnxFMNWxHr0JOq0xdJbuoYFeYy
l9V8GjPZcjP6lWXZpmS0mfJmp7LOcyWnGEdF3Z3zHau+LoVicUenBbSx7MMl
YeLHvCny0CnyajjJqxWkwoJ3SeGjsbw3/2vZCjxSA86LJC1TW6ouDABajaQG
BJyLW/j6x/znsbLeFDwz9/KxAdEd44MzMWWRWEFmVb2QRtwrTQ+u161qTstb
jeVwi7DfQ4JGxIGDm5MF0pDJ077I0IfaH/3suc75JkUAh3xzgFj5uJXRZSbu
Vl+sbUwLnmLW758OZ5GNNdbuP352AYZ9KH6oyvH1sTfFEwOdaFQFu+E88eLC
4Za9MHVrktt4e0DelRyOIIveluA2Fk+ObFDQ55sBmEvLzWwO9GnfD/28TpRh
YLnyIrtLIIT5FDeFtuLSFCOJG/YxD2oHqfoKUtCbq7yDNqtwJoOJ29TbiZV9
K0TAJtc/b2jXaAozFyOcAVhm843IwNpdgagd2C7i8FgQ1SYt4ROaHY1EqTbj
Ft+sfPCe0AonJ2Oqt4etSCoFcPHeyDfFMVHMxBWpiQxkOzNr6lR5SUgDi4P2
u61+EKzmPHW+i4wA1JRFLLL6RN6otCqRWmz4xaRdfhQ0dJlstb6uHvyN8izH
2pEYVV6Suw62ms4SDeT0pREdyDCI5ZhpgHcZvn8paRa+DnYfCoaFxmwiOmYd
arqeiXGOQBcV26qqeDhYLxgUa9DnJTEaq6Y947J+PQC5NSU4HumOJQGU6Na7
KvZpJbx5h/KaDPMnrPN3SEaYPMatRdqoDyztrrmGCOSXfTPJdnbLbZA0BWsC
HP/FFnrHCzjCQLT2DE5TnAyXwR0i8oi0+tIP8c2HufBZLgwcOaiTLsiwj1E9
Srg9WkyO6IuSPbJhkFX9vCgsdWi6Vrou2EoXJz4egHnCq7Th3r1RNeyR+mGS
TCsrKhAmFFKlc/ft/IREucYWQ3F0eZULNeeDhUh4DPrAxJAhLQac4NISRn/9
4xlztsYFDxISMYp8A0lhw5ih8NDp/3XyyCv6+YQBRxjIOpNByPpNasgIZJ7f
mNu/qsvJ0agIM2BeCVtVIAnjV4GC/zl5gUhXRcVYahRbbKc48G/A8rEwnGz5
KTSDDc91bCDTMCJu5K1KN2+sc33VFRgLWnurFD7MRs/3CDOxuGP7JrEOWxmw
gmr0kKg7Q+0qvAT5qu4gcAMY0LO/nQnCEsXcO9JKRb/5JUt6pmyRYNvscFgv
L28axmXoC9hZ3fqW0IPZn3LWUrkC1f8emwrEe03BJR96ROffsl0fsKzoPjNo
8g+RcuGU4kKs3+6PklG3DOZ4CDIiOL0WE8laId42iAENfF6gpRaw5IEljqd2
fijOi+GGm83Uiti3zQxV6q+u7oyN+SijxjDohNWrxFuPV9thNrWG1adEcNRw
mosu2O19AdvCVjrZ830UDJ4D9SaY79Ha6ifGZIdZzrOobnPlOyXJ6gKIWfM3
nPHuDspqS9zUOkIm/gJ3bKgv/Or5tu5Gcq0mQO8M6Hp2OB7DeeW8524P0MOn
YWzjD0m66BLUTtIP0lO6NrEMOFvqx2CxDBL+pKNihaIth8Z+B6aFC73wg6jO
a0mzy3vEK1zEcbLWJd48sM+u765kb+ofElOe/9EDFhrjhDNr0TwfIH8gO7Nv
dMbFoWkwl9SbUNla5WSo2hMIUrwNxIY7o1+RGiy09Eh4OGWXl/BlxmhcnbKO
MdMbg5Ov3Oeb6nbtYdRupbt6Mw98Pgl7/+Qg5q42B1ehnulVaaGawqJyq6YC
NZ4dVezaMsqaPQvH5xPiD5CV5KoUx8X35ZGy8+dXzkvlB3NEaIZyt0xsIJag
Xnr4FUD2ZagBTEupq4L9SnnElyNXZ4cM5AzPdm85POH9UVpED69Icm5zzCPH
FDAyTJ3r2ByPuXm//oRZqDZp58Dv0P6SDmbkmcmA9ZuCwR8KQ6fMIusxtlAp
CPALEjzLYNKNUVUsF81D9Ab+PKP5kVx8wLct/AdamWNndjb67IxgjrPe8tCI
MPBMR3f2cwIw0dZRwpg+/E+9oxVVElpjbfGqM17cg4YlLql/PeDZZz0phxUU
YMzKC+L4t/zmsOXM62pi14Bh19GAypol+JbTrEX/FJsLzyAnluU9/M2cPHk1
AQGWmY15lrIX6OYVJZoXBDs92DGayge2SWmsh2Ac9KF15SfzR4XUfXI5bFE/
5si4YdjUabCTn24WSjRFSrvdlvR9oCVa1XFcseukcaZw1YIf9J1wLSiO5dBI
jFQdalkYTPoNjbaXcihCwE6LMMcbziYOF2vZ5rliZWBlpiqS6oviT5a3Hs1b
1HvqQzcQqY9qa0TF5439RJHivWyIyRRA7P6jLBuf5kcil29YWI5N+PI6lRJ7
pBc3gAQ3QhFXcPILReBktBdRhwAJkPyQfdygYergmRYnSgsUV4lHy+0tg48P
sII9oVOVUlRY3F+RxDLgJLuSWso67A/DhIelbSaP9xk4NFfrlIBIX7qzOZsE
UCIbXtntycm3AELddvQad+F3/7fv3P78a+scrRWb96bGjDAkmmlPE/i/XF5u
w1VPYu5VlaHUaXjKIQoHPKBNz56r0xo7h5F2ARRp6ggObBdcP3yOP6VKfY4C
k4nuAYxbiuXhQ0ghrCybozhkyuM2AhOOcfmUF2WRmM0SAxQ43u2csBLPjV1e
fTjTsYAVni5y+M4DH4RsP1JOJRgoFh/YJqxqOIrhZhpfbYios093GHzbxUPm
0aocFHKNhBxkV1/GFS8n7Tmcq13fvl5VYGmpefwzNzGQ3fmpgzlfjSPOOfeN
7As5lFk5WoY9q0GXh3oMtXlrkLi81HG6vlw2fw9P61QvO9BuxqdgZmnPlgu4
6d0MipTlZ2CRTgE44M17W510VcxCfXmqrxKqspN8FfHQgDpHycsemgnKYs9P
5eSUDuEtJVn6ZJ90LtdutnIxMJq9orNz7MHMr6/jghcI0buERmCo8rI1w8NG
okltpRJJJA8eMB8siI2HPFXmFn3l0ybHXll/WuCRjANHNxjsdS2+/sIwc+1D
+uXuYe6ego0UOsvRN+J2bjb462P2jO3+Wzyou4YsiU9jT8Oyng9wta2rZGFB
O+RMhBL+hXaEjf/zGd3ttWda7c24I/LrblHbWEAvcBGiaZZtson8nxU+6/oP
xy2BQ/k7sVG09vvXoE6NHWoxmA3Q2PZNjGXRmLzcBFK2NZdgvtt7dBFhaARS
pzqhN52IKy6VUfvKSSaEjL1ToCoSayJozjmpTuHGBBs92Y2GIcpxDPaibR/3
oIhlgO4Iy9cumJU8qQ7HLj6dxK5p32nGNjDvF4DXjGQY54LOc2KJSdy3ENJH
9JZFCuK7B77AFAJbbV5LeGYmtfyMBXzKJRR7dcwfhQIbVuhvrRYCPThpssG3
eQkbZdlRhmmkZmefIwkpFHS1lVvloThHMIynrKhkIWZpyVPV4aJqb1SQ+QUo
u6KYPMSJtSa4wEfz4jfxS+nyCv9FbST2Zb2x2Y+BdBkJH4iPQ+miKb9WI7tq
szKWZRyEbOVU1PVEamscP0t3TfuokIfk52GEE4PqmMBN1S9ql352l00I50A4
o76yXGiu3+z3NMVFSxI9KDc5ljLOgz3yh2rUVRANONxgj5dub2PCMdzvTCgl
zR7k4re8tBWtWkD65pGUbXsEXIu910qEWbJ5UpBwoZbnFvpMg0lDOyUi1zN2
DjzXuTRF2630fULOThv4fSNQT5jAJKFrP6juKzR/mKiZjkc6ZVDBM/c22eOr
4I0xFJGDzH+lgl8ozVBHCOVEbe0QZ7KwA+8gjlPdu9jDXVJImwnJSe13Nywe
R8CMdbjNVeQF5YCY+X0amlnJYGFChMalUtXcQRnKgPMBbWoiErjvX05D3iCo
P6DDH+gq5ewHHV8FHqoZoQmUC8ceGlAWdBtQyNGVxuKqXlZemzhkLr65/FVg
fNyNvfTFIMkdUWB4sXtVI5iUMOkCuESw9lhoZIXAejcz/tSMAi3rtTHVq3CE
rOdjs5zKtnaFBmMOBCVonBcyY5yKjEsYtYTxPq6TrTrv1Ct0IygZhCohWynw
8cXlMAo+yHUXl+TqWuXwFH/forPnRNEkIfuJcmwq8LBqvo4OSgnuHIroGJlf
fsKD0ohtmhT1VUdftxRfC8CM5yfVehRdY4SzAvnRBbxj3YWz8gekJNYWp0OO
8LdnTZQ+7J/XDApVthwLrKC2dZP+3RFvcsVIXDn9bVNie/1jxYimF/GkAe27
V67uxjXqY9nLNCuNp2y9kU/e1nMkOLmkldfgLec9W0NNJ81fvG2Y9Q8qHFt6
ip0LwU2Dql6wk0ktUvuN9xOrJtkARXEnmcJTsRwGuYurkw+27S2WTatZtRup
NKeX7hwHgoYY75Vq189cSqQLIsEhLTB5MgEstiAxjS6LguQRHGsjLzFDMjmA
wJT5irzl8rYMCSGzTEU3iJionfXRGX7+jA1z+b+kgRGWwVhtGcJIMR/ohXq+
lsWqlwTiPDVOkEHz3aZsWB7fF3hHvJ5z5Lob42qyVjBBTPn+ZU+f56N47mO1
WA33J0NY6g4E05WER8jVhmgYe2bQbcwAj4QxvymJb6J9dFYBGLcT+AB73Yo2
DMjTCzBPPeiau+lJYFgCycYBqDXjfqkmE+xIjVtKkVC20ZU62g8Kv2ytPSb5
Rs8K/jeW7SIniVCu9JiqeMe4oGKn7vXXpZ2faUuU7xv44O7AXt3QCl3HhYqq
JfBWSM2qtQSzE/wdAPOmuqXTbSN8JzuMonap6jfjpjQgpOYLNURBQomUAkWX
sNcI5GxdtojKlC7aRhluqFF1DuKNl9fhKlSdmS0Efm8TYHi6ecb+tNeTwPC0
gMnmss72pyRrf7w0HHphVL9R7HOPztkiv5FgCdUERFtRUxmd84uoNM2rXocC
+3lwgN5sQ5VaJJJ+z6/sAEJk06eP4sFf1Sv0sN98jinYOtFFrIQ3wxZhz1CJ
CjtTGbyRl8J78JfOVc68N79ku/yqbKasIaEjsvGCvmSvwPPRgHALhqa4tmYT
LFbWG8dzacaC7brPiE0MJ9qk3Y1woeempE3FmyCL++e4Pxth2jmFCFO3btGm
odpQa/mkbVthBTzWB5PZ2vdQoPd9HajSmpBKi/akltPsLcAaf72opoq+UM6K
ThQO8pUJWpEPE87bYGu7/bRAyU+du4RTyS71QzDAf8v1UnFowEDddDpWau/r
x9f3/mlLcehO6NVMPy2bxzQcSQKvPFO9lx0XfGACFx3C0XC+T+v4O5q67VFv
nshA+frFGB1kTIeW2EFB95PcZLWV4bG2kYDZPAssTNU3AzPN0/ZcsYchJg1y
BR613jcfci3fvvv04fpztU747p1cY9X8fYR7oUcaeIgywiDJA16dIytsDabi
6y1FbMA0lNDCV46ub+TtdcuJP7CAabZLpaZeyeNJPnNCMcMzzG9wsuNarh8c
OmDvQoOuZ4XqnnD8lqr3VX+730iEs9TX8WOtqeNy+hLWXuBcIXr2B1RrHSM3
73l606CvbErn+2qoXXId6wG16xCovCl/t6PLQtLxz8frqlSMFsJbYLmKtVFA
zMuuvexklrGCYpEOHN9/SYnBs9E4yOL/bpB/NRKBtjJV+bMg73ccHI04Uqd1
6SLsCml/F3hkb8ztD62DiTovwvte7y490crX9C5ZjTSKmjIulo4C0oGepq8E
tp5E/xz4hCySOcf6/0TdpXVxxVPxHu6hit8Z98u94BeUmOcj0QMolObt3P+l
9Sj/E5hUWHAdXY5ZDhVrxU3c5Ph42Ot66fa2Xp6LQorF/qYwLOIAjZAdVWFZ
dWX2AeHGjQOijwnyeDrSlBURWWaFmC/zryzo6HDZg9IwXnfPTTJ1RosWkwrq
OWDzl/4Yd3EGmR0rdlRafmPogcwhwt27+vop5aUQ8lGVsgLtXGZR47wlUbpI
B8DKDLLXKWHRRd0iqwmWQ56s4h6sIbysv8wgNypvqXEylB3QYmzqMmR9+jQo
gPmSIIh7069K3Z9AnAXLS05ee7OWG151ttFvmMGUENxXEtztrasO6dTs+cmx
FzkL224vKt33tBVeeqYRNnSWOMQEUBu63SIG1UbXij1glvZ3nRklaKzJzELe
LNTk1DcpJ9tayFU8RbK04pzLg0UzQHIc0ovgsb3Yi51C0TL9RlHJitelPlDh
nXwRIvlB1fPGUrn7z893oGlRL8/3+GLJNWEK6bnE4sfhGuLsiu1Mab51J51T
IbyhfR5LF2ZfH8flPjDOXBpSfSFv9gDQWiBzjJwKORuT0YDNd9kEg2nAr62W
BSwoooMRw9LGV3fZM+OEIeF7t3tMYTOUZa6FEoZnH9DVO8si/o+xQ7u+lVLf
EGumc568/gO7A0DDl9k9bOI/MZbuT2+mNU5okC+7ZEeXUpjNQhAXsVwToEhL
ELzw8JI9CFpMSYYbW9R2mTMyl5Z9eYc0D2pr6Og8I9si/7nmKwtsixxI0Y49
jzgzyGSzmJ7PZOHju8gtEfm+Swlw1B1p8gRk71SsMRHOzCoq3U/iiArHjEPl
Z4JuK3cUAeyhAq9KGRDqWUs++xUueW+Rw9tyt+s1lwbjIc5fKM7guNwZ0roF
aqFzTWyWB0KOnrsWoA4kl0tuB/zv0PG6/mht9+VH8x1QSJDP41I8na0zAr5t
IVGPfFm+gg6BvV1RAst3PXKCWkT2+BSnBne2xT6AK9FFr9E3VJLiIL1hnmrn
th8Te7fJXiYITBwNY+j/b8LsT+bqEclCEqIAG3JAOA6NqdPzATinwqaRzurO
jYYKhYefZaw6GvM7sXzKsnger8RobQ7uWRasiBBEUpsLExFtt7lMPHgt919V
ZasBw0zOqda3Yx3poXqDWXkioLRmPfaxwvGPAyLYkUuhIROx5+nbNzu3PlHq
PpmGiDwIdLFYGpBtpYhOMkx6bQ0HbSBIIqhmq6emAaPaDgd9bHydBlynhNT8
LsIXRhsUAsfCup3QUcotywXnXt8DHLk6phywkeTd47OZKKiSJQVMTxVUHG8t
+RBEf7WfxRq9kGNYzHf6evKJjNKpVHw6SbefGcT54EqdfIzTIlvhYpqs1J3U
ZQpZufain3O9KkXBeAVzBM6SCT1yBYBeCiFsiUtou637zTPMY3lbt+yU/KXw
cQBa1b30GKpnETTsLyNOxAozBTdMBIZugWztkOWIy83Ib68zNsrdQ9ppysGg
bt0th6fx0AEg+xaAu2UUQoo735H6cVjf75xOB3PbsAp9pq7IyEd3mF+1S+/v
95ckIZHstywVmzJiTTK6Psceb058EXAFAKVqlHtCYt4OtVrIltPAh49md9E5
ryxJgGeakqei/GwUmL0ERZJdQIHSiGzt7bTgOqfL/kwzZ/a9w1q2HYWMXmsX
hsUqOk+nsLYuJpU3A/hhRZ3pbVGbx2xZjVn+ShcZ1GhedQNaR34PcKxuLb7A
ct5SSlmVjSrUZla4RePGlJ83Z71T0de7xmq60KkatlpCDuNwA05zN+0YuIMP
lZDQu9V7SvnL5vXhBZ3rpPbD2eFiP/Z0AGMREl7s/SV+KmPCexqqHF/nCZHQ
cD+E3mMy6Z42X1fVlbQPu1kqxj9FaADnMmG1CYzYZLbEBnojnBml58bnTjm0
oEJmL8xQb/gweqWHastO9bGGE/WyJedcXyym7ml3OpnDLszHwwW9euC/5nud
JTgvDCFw9M5XUew0DbOtxKaZlXmRlK90fEtTea/dgW5YAEMEKGlNkIk97Cz1
HSQxr3oepBXh9PSWH2nEUlrumWDOQtUon83TXmnuMeWbm/u+hvsNpmzgow2K
iSN4UXFmkAjL1qEgFYoZxLKC+gsjOHHgO1pctgPP4XMIRbwCAmNVauw0rhex
Wv/C0g9D/MSIJS6q8lubqBI5MQQqCrUTX2raFMLZUZeiBi2Ky8NV4zBdFCBE
MvKSyEi+eJMgMYLOteuUyV8fopqdOkCfcyGEWvRV/SF4PWMdEdLWv2izQkp+
lPPoCYrluU55kKgGNfZimQcyAnQDBtJ73pqxXpEz6m4lOfFdn7GKbvY1iVT9
UYitBe1ND5drjV/mrkzAtnKgeC5dlBD93KdFiiDLUGomBg3EBq7nZjVUXOqK
h3BEUPX2nwUHfzAXgzvRziCb+StQisD+bx+OSM1Mlgk6J6OzPQEpQ44gzcEF
OnwcAfzlfscK2v9FeirhkDor7+1NzcL5J3NmOfoRHhGSPPJFrqVLkL3D1uWc
9nGHcQ1pttJar2M0RQj+lCLfTLLWd1FmsEkOJQTl+hjnG6LVO5zlCEBauiHd
lEdWGEljRHINJvXGgqKGkOY3xGOlpqjDES+Vn5n8wnuTfK/ePBBmpDfGMWN9
nU43dfvmgK1j5JQdQzQXhrDO487YFSHl437scHRD9J48sBIr5j1MiS5+BEfg
UZqWI5aLV+wlCTCAvHNW1tH4pInihK7FHS2VdWzNWyNFeGSUMwI5YJwDYZ5I
F7uAoFXNTUGuCHiBSlwVSLwXx6a+Mg6ew0TdRhFoLmpM8mmIu/iA9StqRTiU
kxkVxTqpbaV8OphtRIZ7vXms2Bvhtvs8zG6I4bKfNV8ltNvkT9EP/ZvT4sRR
ajtOdDKAGF8WqZeop8qh1DtE/92lVmN9xUF9KiEHg0EGL0FLlpT7qdhnKUVb
g56/iU2w8XQw6OWgyiFeA8Q7eSnhUXxFeG4DNZeagyWuvzOQazipl9Crgx+c
JJkAykFDJ+w+x0KJIcR3vu6VOuySJyV8miMaF/HQCe5XfWTM99LdyW//LJM1
U2u7UfasFuowGCqjg4bmIKpprHXACSbDZcn1CDRXfzeckozKHfGd2jTBCue3
UbkOPUaTMT3HCDNioliUpAtIt5+0MlUWgNG/3mLgPWdOIaaXzc3g4FXTBzyx
aQrb6MJCWplhNe4bjX0DETZL1ZEEEiTLTe9jvH9kIEi5iNnHWY7CGB1djZXb
zF/MTR3CrW/3R6Ts5uBWiIr1F4uAWyOeZC1PYjQCyHg/Pa7/AfEpEV1z+m3h
ZDCrl55izEJ461rUrogslTm3CZ1vF8j9yvQrMfVy7uIYGop00c3SYCkLm1K9
452y7+mqjjj8FjiT58B///okFQgIGx3bb3hFX77hzhWU51yTFRdrplJEdUfr
3U+/386L9YtEWrCMUCJJ8dUwhUaTVneTNxleovBGApggxyEiBT+01iDJzxy4
H4Jo8CHzWe+UYkltlMmy3b3onJqGqn63O8je5iAhoPOwncJYTr3rUxpG+oLd
NdyDyGpmPLDharpyLGNkgKwQgi01WXmZafrLCf3YAryMlUAwlG+377trD0o9
OPCQEenxqkZCs56wlq4raH5rQ45zZBlkX8JbifCikUNVurh5LyrWnof3vCGf
LgaIGz+79C1JMLYfkL8H0Yi8auaQFRpr48zcsyBgpBHRylg9ZiXsx7Nl0dY6
SH5vyzhw30XfYdCfKe1l17KzYgksHlO1uiAuuGHXaprnVT6mvNnS6F/6XeXH
LqVgqsOfqvD+rKY2b1VtwAFUQ0iu12BG6aAvSgcRmS4XxkQtTC7lN0MI/ngI
1AtErq6KDcI1rD9Z5Vp4Dl6tWtiP50/MIKxcowniKE+E7J8P7V222VE0+hRt
JwhV9M+Ny+s+9JfRl2FA4+fZArmN9cNkwRgGnOPZIDfI+h+XPD2NH/2hcTUh
O0ek0kynYBG6Rti/XEnFVopObe8mmngV/QLh6hnbnpRaAuc4Dy86YCUg4ybx
uoICnhTngNmSo57sbn1uxWk0+6Fqq04JgONnk2fMCa4Zr+wVs05ipcUB8701
YeNUL5+cxBLhqQr+uSJuJySsrDz7gdzVZpA2xAELzhxC1R49sIOI0W4M1vbI
zPMDD91e/A6XvaOFrPgcB5TntjSCRqgpq4FG88GleFmOI2gsdpxByaJ5W7sS
Z1WuwbfGFGYHLEszDpP2lhdGMVNxPNFXQ4qPQJnWZrYbxG/V7OltrYO9JzRS
DQxoE2lFrdejJ3qW4Kqc4sP91y34t7fZcyhKZVkvV2t8OfGmr4osNIc+XFTt
BdFnPxHrwgHs43/Ghs20Z3CqG6NqTIrxNqAUQFAVrtOuR9y19KIQJ7S/Iv6x
72geyUXf9eM2Rm+nQlSmhEQnaYBzU2RNA9KJN1piavt/LlFX0LNm+ITwtL7L
NUVT4SvcMwxEKJ679IxCAjhPs+8fOVkHpBfZ0E4Mg3MUVl6jkQixPx7tuRh8
BwvO6A9a/wIeHc9myunhieInCqMM7DWZvz7lsAJYEarLiS5rsAKQV25iRiE4
zepkN6Vj+peZsCuR/HR0654tvIyU9gd9fIKAOce9Nh9M21BO5iaxYTOVCsJf
Kp3nltl1JDAKvYDjD0pl8mI0oanEvFk0b1Xu8Z/Q8860xqHHwLOeT6+cGwk7
rwXPihq3tVx+Ybc/JllGY1vSmDSuBCIOW5V1lEA/4VkCG4GQ5grmLJucETrs
zHAwuqg4lECr0Xm1ReDHSX12OHZrhv37291gtshWjEcvUm9qnpNrk1+YNAeQ
T7rH8gEZfvfUAava0J7VzjpA7IGkaYcfcQDqgJILJuB4ikFUmukq0ANXRw9r
6ExnKq+6js0xHWveMVmyt4HXQFmTx2O3yDR6Sf1lfRZwWJ4l8N/gUOnMHAHX
rfBy2ES3zum4obFLMhWU93JdCHfQcGlbfwM6vTlOz4dqZKj0DHCbNGtsujJQ
X/Xd0tULUbK+t2/46I2gA0IcXZzXV3voE3+NPhMvwviLexxqw3F5YSIjSIpf
VaN0woQee84+0h8ixHiwmqn8ffbPQtHUcQ/Ns4lzgoohVreop6KYt7c5dyK3
holQ4+UFcgfeR5vJrdM48wA4KdmFOJkPbUZpL2rgA0a54xOt8fST9vzQPOcE
uy9zgo6DT/UB4/0ygrO3zqmafsLo76VMG9qdnh8Z+V2wamb/9DZNqw/qH9pO
3EvCjrbX1ISYMLStn5ADZaJ5l0tS+QNl0BbqrTYsKZGxtk3Z5zKd0EDKV1lD
avftuHyIDuayMyoBeO3AwuhzBYGR8U/b3VzYfZCi8a+x4xgvrcElmfweTPYb
LRmeLWbK3Mg8wbuUqGgJtkG59Nl+MzCAdXqp0JQFvWLHFmmgQeGHoaG52nxe
QIibXaW0+TLwLBx5zmOUe2tIEKdVsR1Uzu7sX5bCL08RgdekkWUPzZXbjtFn
qI+4Kl0CE7jxYgXy/9FUuSi9wkypD6D76nlnAlltAH6yBsyiy9Xqjr+BvPEp
jXouw/a1WdU2ums6j4yOWOMph7Y38u9tuS1OoL+B+GiJX+h+n2j0xRkTq+fV
Ovk2/JV15QbojfgeCvVp0iShd0GaQP+L9Ejfdw+hDvGNqXLEyEboiCVGgQpZ
jrNZto1OnzEZfOD5+f0djWD0ZeEVVUmS7DqQJlaL/HqOi9qE0vpnDDRZ4hYt
3h6dAneuRJRS7e4Yp1T9rAuoJEuLkISebIKo55V1gy4Cntf/ZDXw/wdp4pHQ
bnV8YZUkZ8qR5/AftAqLjV0ODNPi+MCyokFPlp3YGUuK+M8mwEgKUkH/cjQZ
0XeKxZk9oEqh75Ge30RDYp5BOCXL6zOGZTMzfHsAGeqqgtOIXuVB+1MJy8U5
vDpxCxa3YCrNtczS58EhylCneIqTbWylARlh8BAKPXUp1Is3PfptSG76zbFg
pnLpW6RcBi3jYZuLrFv53mDd5lEqvUkbtzX/p3kXrPx0obDZQ3/kz/SwuoK1
9oaUIlZ9b6bpsGHNjN6id61bNVxab+IiUib6IyY27iX864iL2rZgw3Omlmhy
NFRshP56NaFUnykZNkyEEfNCBd5Vy2H5at1Y9eYym3KI2chgJttJbBCPFqbf
g/6eQpKhGTu7B2g42DsQCOl/qgk3lvJ3oqkTn9kJW93Fmb8nHIW2DVsL3V41
33oMNpntaOlSP+ASXcCjoDH2GOmwWa9FgP9O+hIQ7HOvHqcGT6/Lvcaz57db
yysizORefVDUx1KqzcDe6YM3iD+LgsvUILa09XqGUduE2LGdQI+lNHbU4wSd
ln3JI72ZUQK9etiZj04uYEYNTatd5kZuv+8krB9tZ1mx+rLskbRBMi3PY66V
3p7XXsPD9lzkueUOvF8IGzBn8xM7bkwTH0pmhDLcNE6laKEF21HnkNxuMhDa
vNnTmHA74hdpbKZhCELiNFRAfy06cdCkNLnRHqRCXPi5MTH6hpKPyIv3eDO0
yOGCokQJ32DltRf6HSdy+2yxK6ofpZmPUCKlKDKcyuy1dh1My4Yegv21bmzu
1Is9zRUerlQrs+ybFAeV7xasJ3BXqfRmv72Crm0fmNbUC0vIYBlEMCOqBsub
NrEX5wrSZNWS1ij+HTNuIrF3bP/O7e4tjJcLodGJ8rmVcDUEV++qm8Kwuf5+
W2g5+IjIoldUTGzSGST+wj9hu3oFwR9W3iqR/JtZzy50H7MKku8HOGX+EnDh
IXh6g3PafqnVLx9XNCGHHMVSlnadatha4Ozfl5/UmUxTlf/05lSVxl9NqrPD
4IS7ZQ1xlKdXOWeXVpxlNOR2XTm3OAalSB61tB93cZI1t1vij9WvureY/Ust
CERNL835dJQK0dc89iJ+LChCtCYE4tP/klGhgIQcYnQC/Z1GVmBLgAyT9p89
NAU9v4+QK3dmBxQ4x0WNKrq6yL4w+kq8XTuuf1u8YcYsTlysPlSsVFP8Fx2i
XKgGhkTQ1sHr4/8PwPtUfLxBOll3mQTaP8mpyzYg93iP3DSyR2SE8Lbl4AsK
cNIEOAibd9Dk6v87Ie0/aVTEQsZGY/0j4IVf9I/wuuNY/2Dz0Vi64d0GpMsl
7vDavhhJXjl4Q9LjcLp66wcSKA4IQ8DUpNy8N7C/4cIyKFH/0LNyzCo6ueJl
Ew/9aFFJohA1FXinfF1gLQsWRvnBJpLEuHN1jW/vh8iAZ+od/sKTchTxns2M
wNLMK4n8CF8TFV5Y+g/1u8d6bFHaCgJIm5hj11OjWX/CZ16PkAFDpiBtbCDv
5rVik7qYwIJH0634yOD+JkLQKZmItdWN7sJx/v6Z/LLSFrPhPlUWk8qZ/ZFf
eQdePXcJN8F7wFppmFHbi8oB7fmpePJVV7no/DeEO5ElgJAL1wPuICPQYq+s
80X/uVzW7ew/asopc7OlOemcPixAgegdqo3LSswlIx8ZxZFYYQen/DH0kOBI
zW1jp2E+nVuflNuq/zHZTn9Br9yDa352+FDlnO+luNLDWegN88kCVfBFVuR1
UyWdAR7wu5WyWbzRi+upokb3KJ24Q5nqZ+IuIaUQmR67vd5WflNIl3b6SDtd
rAUuCh5lVbXxW23dd5L51e21Fl23NW37t1bl9kXxrZsdVi1km6ooRxyvkQhp
bGGLkezjYUBfJKAeVYrRJhN085On0DdcR8DAbgluumLutHI0vnGQY2DAXRGN
InukgG/1Y80u4p4gQ2NBjCIz4bPUSuRybqtBnY6Pv5I+4cKdBUStFgSjqbll
dlro4HgZz8aK9VQ3s3DdrjcxMxh3pvTlq+uTtzqiHfVFVtu876Pe6OCJ6fPL
j5IYzRHLZJAitb8oy0MtVPDWeqyRHr05Guw5TgX5w5DO9N1UG6TT4lOOnL2U
RTkJ9/ZDt/cu2vr+HSxRwInHKVAzghfffuQ+ke5FUYYZ8WzTIFcJ5B9zBVRc
wuRAHJCtUNZX2sh0borF8xC3FJvSRmAfoIu//R8YbE2XRft+VYnO1RG2F0eT
avFpKhZhLgHnUboJGiBj+1o2zr7mvi22sWO+FUJrqWNdgoyFRS6gyT0MdYJb
LfaswjBzpbdz+GOOX26G8fGO33ErTjD2W8gpNh2qdAe0WYJXpF56NOlPx+tg
rpX6k9sWkomDQyvqbGgnlEJNnbrnP3qYM8CrMavIec6gYxp5ySyVTi+YEtwT
SxSAcdciR3aU0gsFdr24WtDGfqHRBNlntb49vgZ5gD+mCwfqbi5EG8Kai22v
QnaO6hm4XxmvrFRw7gRgbB7N/R3nf7CCnw2AbID+otBdGxf48CyuyLZ2x+yt
u8J1PWLASZjavPqTsTwpTetMIrOdzlymC0Z6/6FnC5x9ezUQhclqSqEJLcfC
rTFCBgKD9+2gL6peqY9xubHxrvvsdByfnucn2mxcjXqYoLmdARea66G7R3gG
0EsmsCF37FbP9iVLGJAz5oDp/tPTM8VgG/cJCoG7nBbtGZiy0I7pCj7wgl1P
iJeMcUs/JNmLe9WuWqF3uGmLyPJ3OMqKZzd/rp2JE3FS4OBzKvNzvd4WeLpm
QdKFFwRyn59lb9MNjvXpSj1QsJtDLjumba/fgtz2pmipxIJ2LEWqLd6a4F+u
e5H79cRI5RTFBr9Hwk9Q2kkzcrYDKVjpys5sHu0pVu9qijwrU1BoMltZsnTD
CrAGboBNd3yHi8wBHYg+y/S5kvUpGUigtfLa1e1CydV38XB9mhVA1wKk4CXg
x4dqB6fg7zcuM8ZqSKHl3CBVdq+SLw15Hz2mFI0OHChGvXC7W5olfwII+Bus
kYQuP9K/3VniVYfKvvovOJSko80DHZOXeV9JPOGSX1iuMPKLIFllRX9XXfnZ
9IkxxjkDZLxFFf+oqm0+qFsE9azIn/55pXmxFgC/DIhBDVvpbClQKsNrSM0A
8YZvzXvRa/OybM5+zD7HfsuVAVyy1qcEqvba4IR0S3sA+pcpk1lLeuoZBl55
RUMLYoxTSRBSZDWDjgUN2am6+Akev/Bbpu7SUMclihEEjByod0dJ3cMdgnaD
Pj31o+eHA0BMFVwnatrSXZ/+P5btB4/crTnjQitjrK+BSUJWQPmYfZyRlV6g
fe0Zx6YSPYf4IFiAnoDCWpJ5rUjYPlIcP2+l+xsiMuS1Ub4QWXMH2OHgWhH0
WQH2eEx7R0T2UmQm9zV4jb3HiO5QOr09xpj0ddoEmLge18rxQrq/RSrzAaA0
SnAiDAYP9V1ZWGI/5jfAf1S5KZ2ickkKhCcIO7Qr/zPwdZ4oMU9h3a6vdnTN
PmonHPcbJDH9arEKExGVMI+8VmeCguBh9Y10j2Tep27Vq1tFgZI+99C3SYu3
wY6NP29CLPVtRrKIMOZ5/2adIq1Pv+Awg7DU5rOCa5c4bWNqkcxXETDMXCXB
VBhW5QfJ1AEVqCK/j/JyfcprRiTWIje8Oo6/313MpCvshb49jPU6K4WTrwnj
TVcEWSD4ToHblV09IkChD3G89KB9F+eii4PG9TBuo/0SRuJJEiyIHvj4pCjM
rqSB+/Ubs6AVF2Jzjgb3bjLhjjMLxQHMVGC2gp1+xJWdk+V8SbPTCZkCHzpn
yFY/6tkZ7ea/y4nXep6FjvBN+wG8RdWqvsVREX2yKpPXS+/JrFsGJ4pgbdWk
yw6q00KQZSPXpt2/1tPqRx92a92Wijmx3hBjHT1XwOmLWj2TsGHb0hhDSoJ1
y0JF+UF9JudM9R+qRga5oVyhkxB8gxgbDGDHtbr0ccp8IUBtLIa4Zlrdu7yu
/SvhS5WsUNMJCeFqd0ZfUQNG4bBHDQXiNH0AlTTAUVXED9KH8ByhL0iShCPj
hXF64oQrTqaQ8Dgs6YSpjlNsDMj/ZYBAvFm5JZD9MxcWXFBdoii2sLjadBzd
Rn8/BMEsBFi3ukIHNKI81IYwsPwYFQjGca/9bZaSz49WpXDVYVW8X6Xbth7b
YePre/7MwzfyplcfL7VysJhGFUWVwTlws45fgvPbbQo4z61ro39aGUZa/Qhd
9PHueyClGI5SFY0leaztP8xCN3WqX/HDNQw81JU6itSFFT1lJkXCyTxTqYb5
QETYQNQiTlcRb0YqXsVFj1CqFYkf0y91Sjyny57UnBDd4gzrAZLJtP6WZRsu
5QCeF4ClQNNzD11rWSpgz2m1zRCymF0Bn7x4nZzHB8+rFxg4hNgpdn2O/+Fd
6CouaImz8+9IveMwBnpXxgmQyVERmAsSVdHD3W/EWxFd+huj8wPIOYkHBq+C
1cpZPZ4TVQ7QudwDnVFEpl+ziRpufZPD+Ri97y9Ts4tKn+fZt+CXrjafQ3bl
+QzqtsjVdSmJDbtLsuxmdypyUsN5MpDhga88rMSUF7qnupiVzmh/iIhj4aT6
JCSaAbYB+7utfkak7bYMHSMfUUBzyHJdbxcjizM+1LCLeH0n/mslvynyZ71C
v4E4spDvPPwojBlq3491ar/GRZdid1gbBC9gx4zmue1148e0K7b70teOg5zo
VEsrgCFGs6cT13WNclZolVJnsbdlRpx8DpBfBFuZUftywNZ0SHpwG3rn60Y5
woxqviRQyov03Pn6SrKrZhDfomI/m64YmZwm1qlW4QVQXTgNI+0c09l6/1du
uflCE5CV1gEKvjI+fFucwccgmSNVtN6+odFk4iwL3oNGcIv5fi+yaqheq/uX
hQ3ro1dy5NwtzW+tWkAwF/TVVg7CWejMRgS5/gyzRG1R9wga4EywdkoTgvWg
+3PFIkYy/jOjQxakvBpTu/z9en1/P9XC3EL/LzmfdKxBAkHjh56BL8kyEpgc
ERxZbz5XQfL6cDzekswzLuN0N4C5NAcK9lH0tHBOemdBysKUtf4KziSKSNRy
EuUGIss7qkIpvrfyW4PJC1oJRqju2KUqdQ3aiKofZ2J7acFXe76sWqjLfNaO
+R10UKq8nGXg5M2D7VCV8VAN6bHTKAdzcoIrlT4zFEsntT5K8wayf1Ie8/zW
e1T83FLq70hy9t38mYzDnvo6vK68nzC2ULSz8yGpix6FjEc0+e+NLAlpAz8w
Vm8U3UbRKmoU0MrkCUL7gW8W2pS0WaV9VM7cQpgRIBk8oJgcyUcxPEE/H7np
V0xdvZnqewMZA0lIIWTK2ZIwzDgyeXpRUaxC4eBBo4FkLIy93wB/lpzfUoFv
zSIjPHWjKiJBJX8gzkYIw7dI3y0727gUeSgY2pNQEllxelYZ9v/X/8AXLYrs
rERLfxzoaoxhe+0VsV1RoQxH4/ghWkjMjtZXJXvMNDlou7Cc8dCjv6v7gomk
rIGzY/XbEdiWQPp56yLvLmzvNrXp9TgL+PFRZ5pSxZdwv3SPpch647T4YIox
s4p/rVH1+u44q+3d0/7cL5RFmuwIvGy0h5J2TG/p43m3XC5+LoXGmERXgoWw
zXLmM/I+ShnywnbcsSLL1yTsp6Uuc1GpdaM9DhU4Y1fO4ZlSJ85UCbOIFDcK
R+rnQGnY/kqMHep08QScYwsZivZX42E7UE+e+irROCNBMP9WARV8bUqCe9Lw
0VKGoLWQOwJ821izy/qvwOZbCSoeUzovbbvvCcofAeoen1g/i94+1sMw2IHH
D8cDAMMhmjEWg5B4lCI38zH6/Njx3Ali3RM8LAwko7Tq4IdJxFbSL03BDMoi
VcG+B9laRKNsu+nEsjtJ7XB99qqVb6NqvWDDFQVEJRU0eDRlAIbXAo7OkDy+
Amc5jvsnAg8JKcBNlUEMnd5A/RT0ayoz4g/NzkQ3e98idhdC3OUdldiyByQD
G5SGfvfR0nYthacsTDRhxzMi3Pl6OboI99pr3Blh3Jypf1qzv/x2zoo1xBRl
+Z7dMdvVrcrjnp31Gygw6ERJx4NX1+ZFo4D2dKCCd2MU6pfXqWu9weux2mxA
bpTvFgt3oi+60D6txdnmbLz7n1aCLJyV6sKudvWmh72EogJp+3X8TLDSfiRV
s0B3fMlcQM7Eh6wOSRAQLT42YOQx+fnkqcXyHKnvwXmIYsZnkAnpUJOObJrD
a2UZl7o6DrmXLRw7uOVMzuVCRfQB3lDYUPnYB2AuewHwaucvbzr3wdKBlz8F
QNeWqXzQ5fuNyMUkmkz+AQguIxYEyeg2sw5YF1ooizhjbEFLJEv8Q8oeW2gG
BJsfPF27dgb9hChnCKlCm09P03/3pA6nVReCcckqc2OgDyqWp447+l/xhZig
OEFZlCzYG0Jm75q1ls4Bp+VRf1BaPqZS4rIDpZxzWBTOVW2KFP1RBacWMAcJ
A1OP4Tqt2LO+rIXgkgFspXTeMpzJF+2ZbFyYusyEHNqvJXtZxCsFio5tXxRC
KwFquS4MkvN4m3QP6Hs8JAnqvUMBO6ZyOIRgEswrN/w3Gbi07y+GBswk0iF3
POcJIFoo3k9LYodjEm8jKzsiacwrxXdfS+j96+8yW4VJ81r4gesidBx44Znw
dCEH/nhvSfkEETjKXBARH0gpj+Z7RAx+Zu1vG+orK4VDTAIZmJ6l3UYEnZD6
qx/FoQx3rcqSPDQ029tBahktu/p+JsvhaeNgbKb1C7vZ0BthcfDMAqyYOU0C
5uSTyIX2t2YosVuJhCZGXy8VZZMadiuAxNaUSUWsuKmRpZ9+oQQ/xg73WFPd
YwqsUiugk0b0zKaORfYXOBBe/BVq9xmgGeR2hDUFmTJtCp022t/Q/aMIeJ5K
t591aZ2A5XfGzUMwzqbmMf0Hio5egvFqpbdDGq3Wvjhelglf0GnrQus+GBlI
knXqHb70pqFGkAtoAB/xfZKU5JkukYzMtJiT9N3X0sNwBYVMSm2I4G7DXKx2
HhV4wFgJAo7r/DgOENgFMKCv8Bz+kl03pnYZRzQkBnkfn8F3wAJ5cXXEr0ru
RVxjFPxUApqvovcofQo3xWAyRTt6PUdrEKq+tVAAeWT4zo7vD+fn/mRxa3Kb
0COiXaaelzA0z7iEsZehVLRqCGjYshGSw9YM8thx9gfrn9ySS2PGsC3ls+KK
0FMlvSmVYxWxgN0NV/F2XntQPoLG0OhXykNdE5vuA0r9pv8L52fVllEkDLnZ
JQVm7n6PZw9S7wAmBPT4VSnS/WA72zdyUPsgvm85eMzqjDbzT3j0JBl758fA
w7EH9l/48A9BVxkLNPHFsdzyyObrQOjJXdQ89eDgGABWpkk0GyNDdPVcVzV6
dLfxglZ65YdT2xPpUN8ZIv3xy9VmgETVNNuBimXyiZZ1SrJWS/+J6dJ0Jw7P
eCVue6+4sZS+HdJNUXuvL2SbSkxBtN6N+oOh7tKujWNpVTYq1u9h0bAF9G23
spRkrNKxraDK3EOCytLj9MZrsqPS4JCCthEAvb+6F3MbN4o6GjX9G016LsTG
0gbQKfLe/mfePcfRTTzmeStKPtlJFJMcow8TnIE+KeSnmY9OWoC9QFr7KEPe
rG4jmNLb9UZPN95vPrIjmuu70eNQvn8RIeveA/AR8eis7nyyifFVgZLucW/z
hM1EmPl/Py65keoJcBhRyxlZYloB1dYeP9xvasQlLgMk82dhdTSiihopMDt8
MCCKz24/Zvovtg+/iWPFSZCl1UYP0sf6rnSguR27NM+7Tmatbko1KQW0WCkx
ooU7sAQ4QeAfSt7I9PRfxh0oTE0DM+7NoXd2Kq0od11vAvS5KIoCzpaRINO8
5TPbRNbTanXxzYwMFqTxfYSaCikpmlXnWUpxciKo9ZwZY8QIHjuFIXeG4O3z
35q5i//yetycWlvi0h3vWKz58YOiCO03iI+XOBKt5U6ylR1No1DrlJYdLzPm
+xaabxdsdMWv1LdLOMkpsmaoJH0yLut5+34+U0FJ4rpOizNT87GoXXe/IbL/
j1Q28PyrSG7NuWEtNSxB20aQBEi3SCBkCx/l+FUEAzIefMy/QBP9LiuEwqkE
1u2JF1AhwcvNLNYtOC5yRcu6omdCfwdzwLgcRt7QDTiTjWjlB2lwyi+LxITE
PK3yGLh8ELZJUkMcKSUbXEftoa2nCdf3CnuVOkltDs0yMWHbZTN/ARNkH2Ry
r6DECpW/ON63JdjXJq088ZV+A/qd8cT6lnSftCQEMa8YydsDgUhogxqYn2jf
Mrkxm2VeHYLwfnYDXOh8JrIqxL469gM7IAoO53odJ+8A5RmQ6PKm8Lk70rku
cPlIItkLPSySKYRPV/aGHods6Dnazpv0aF8fuU8qoKgt6vP/5boPLiJGp0KZ
KGnbxlRe5a63AHi1FNmiOde/7hKWQC0VfwCzod3hmaebhc+5LrOWK3JSSEzZ
2pHJKoNowT+jf8asqK1QyU1sdvwmtfL9tTBxMOgSqdPQDIkz/r/F1VNpmaLF
oUD/i7lvNF3eRLAYCybuHFNPk2aV3VIB7Zqr44LWCPhLMqUz7EtMQSsIQs9V
aHN8VoNH1sb/U39R7GQYAKOw3mtm/4nJWOVAeI5bEVNnE+eUrlqOetE9Fcjp
Z8hQ6z/xFNjh4XysRqaXCWoFCt4GxraIlc5yfQGejJEDSJI1J+Xj5cGUaISm
1yHgSDZFEBw3Qa+KgIvpKWxK1pahhVHLFBybSLnExnKbkSkez8QzgSoxX3Fd
89KZjl2gxOvtNna0cmVbT7MCbFIjQH9LKAjUJvgdRNFzNTd+e0vDKpgj7xdz
w0deCBV0B1Nj6/MFI9+gRB6cs1G2xrDdsk9vFSc+Sv+l3Ax3PGhKbQJSt6Q3
yWJmxp7aasEim00JqRjuWDpz+wqskBcPgdd+Ro1cZKETAd+QlM/Yz4w8a7/p
LIyi0CYTUxpDoLeYyT+nIGc/IwNuscy/4eS347GZHpiPdz16+SMNuC7xmcCx
QQlraoyDPj27XYB2GRcrs9q+FUwZkqUmY+12dYTj8QA2cLupKgCnzpl08dcy
g44HBITi0R8RIxop2n8+rU9O2uPstULdNAr0e46B6wuvWvwiLNIKiGzY+PjS
fMfEAw3gEBSsOn1Blzjb95E5Kg92MfgtYLmDlzGMtg+cYb3stV2FwJ7DxYBh
/fw3HRPw2U02PYXpA/y0mjWwPV5Jj4IpWuvV7rG9VVJq9EURqKujdhLi9x1Y
znEQVqdiULwgO75wTQZgIbVAdBi7+v/4vvqnglXkPnzhWdIJSni80/IUcI9F
pNylj+jdN4uoZPUBnUBtLPcK/SrBeOBVhXcK8FvQt5q/8jgwQ45v6ztcdTzU
jRjO4jZaUd7O7BUkAxIRW6XG0FR/Qy5RzwX6iRY65EkNjfyNqXP2WKaSih/X
qqZnLmVGiR0eElTxLenLru3aAl3z0eiNU9rgMsJhh3DHUzY1nUt1LkLduhKl
r7zgBWoXIiWEwuY3LV8jsD69BkPrLBvxiIH+a2ioFE7eITgZubAtwTdxkMdK
8RsGFUW5puDxu2k8U7CjzRZ9fka4JkyWp78QN0EJei2wQvfNulHTHIdc1gKu
AFo3mQs1HmJjn2zuQni1kJ6HpLVoJapyhlrD8z98ojOcyRhCR7M9CisXNJq4
h8HTAPaotwVgrsGm2caccdYXUjmRPgKOuRbzkXezDgBmHd+ooSAzDRpafuMm
Z8oMoNxc5phbNvamitcSCriKiDVXwPbyVHfu3Iizi3IrssujzcGKWg1AaENw
/gsQs4BY+1Yiz4ObfsAtqUUdUdna6g+RvJ6UFCVdEbv4SRx/CS4S2xljGhJz
fuOh3dSwrnlKHZikB7N3NmBl5GfJYl2wC6gRsE3SktDT+qUMLcmKuWc/94Oo
w6uEsRJNlTFAzSBIoXw8Exus1j4g8p+9nvFN3wtwOSp23caA2TknPbq4sjeq
nhlApJaFeWF7IFY/w0HJkOV2UcvNPmVug/W0AO5AC3PJxOmX3i75n6wiiRwt
RpowkMfM3kYAOSolG3AyHvqrFu3BFyYgFTfcAE9IGFFUhUIJzy6HzwWrX/AY
NsMiNA7ZTf8Nghwpg1nXK1wDgFVqY5Xsd+TGEbMVH+unx4SqspSKJttQ3kOZ
HvQMzL/lfIq2q9oEH2rAb2BqEjBAnKgnyNN4k2UMAhknod1JdA9rOfCMvwHX
tbW4x/x4FlakbrZHRxQRmsJ/gh5yUUWL1XwQhW2aiX953H0PGlpuCsW3nSsY
vwkzpCotzO9qVIEbwpAkrC4KeSBEJ7ll33q49XiIp9ZjQIVGZnn+0ctl7VVP
2y9dBA7j2IAvwo99SCWJDSQIKu54keNtNnYokVFe3fVMjMe/T7ONTQwk5DP4
XCX5VJdhoVVjyiVoZUT5z2jNXy58H9lIyeDEfUahgE17J88rm6alyARi6w5j
XXe9QjBUAfyyc36EVvIqUnO7vdqfO+VpeePvppqqavv3DnemcrKS7Y//fszO
3XmqVoBig0FV2fHamN6Sq8ZISRA+R3eCUk7Xt/nZfvv03exj/ARyAH165Ki2
b/yDkuMdJPSNTZP9WgEPtXva+w8RMdDHbqbQnQ+gFO+iTgKcnOEcBcme6tu5
CMflfYj/UWDMiJbiNZVqN6qciZydB00EP0mjldjfrqhKvi+RdVR8rOHuk3TL
f5+Y7NsGXNnRp4jD5z0iDIMM49cvzELGPGhaPWTM4PtsG6xbaxTBbliLPakv
Snnz0jr0GqJmU3xWNsH8GojH/p67jf4VipnBxEy5mHTiz07HU5y4Z5pcta21
AYS6/A0Y4/f/SVDEPmLYKYDF6oPPGA3JTp874qrYCv6aFDevNwGD2Gp+pdZo
Z2/sAIwddNMrxdG/a83q/H6qGGk4QeAihQk01ddD38sUEkUzNAaIH3vutSHu
BYMnqgCrUDCN811vWNlUdFrP6R+wjnXVUweC1fJNze6/MOfaknXZY9PAn6ex
3pehk5wFcNUqkO0bh2Cib3MZeGkvqSkPn/ETOw3z8dn5G0D7RWu7erMWcD1S
pfyVnwsKzBWXfM4hMq/Slz/RFgVI9ozWoKU+Ek18NZfDNaqD905LjFlGAQJS
p69QJWuRTONELBwKpYVRSzsG8Dwqiny9N4xgLrirkpLPp/+HFHXetA0Utx2v
WArKv4ZTezhOerU14dXctnwA6q3bS8rQhbt+lGzc5KhANOQ19SnhHR31DQt9
HdxuRL0ml0TF3PS6cUr2WlL6WUIiYJT6lrTNsa7GdRmA6DP2JfPLmHXaGC8q
5knOsxgaL8KN9E38AJUNtV7y07MxtGD8WKlbzBUDUFRLatKyyq2SS9JppH77
vi4ak/zwxTftWui8h2bj/dJQPb6XAXPo7eAE7MwWXFHLnw1GO/u47yAep07T
lC88vT+HHjVR+P+4NfVsXnjnoaoedyRUZEsQkv9Fo/VXdvn0053ynxlHeq3S
ZU9v3n7BfoeLAR9Z46DADRk14T+LX5xhlv3J+bqMX1eXv7sMSpJUUYPs+sdG
edatVnRgHBCSGXMcp2pL069B4JYfNeiyM2zJZDnPzIl5USJE1XAKyzNVGrqX
l6giT+JAoWXBBPmq5SkUDJl07IGrQ166wQ4388AhN0GZttWtR0+jURF4SxAR
zsmpPBi6y1GcoOe1194AIFsl3mMW/24/vY6bx5wIaUGKLjka+CySC+ea21tq
ZiIdoGSaPwYdbUIK1aygOAnRucY2cUYLFg1LSmce/b2170sETxqt7N19T5W2
/I/vxyLOz9NEqE2Gn7rv4ljamnqiTyvFmn68ILNOyInB3Nsx+tYUGH77Y8s9
ofdN7VJk0fkscvhZx3WzB1KfHOQqxJIXmqr9C2KTi9pfvByNUWTEFSL9md2O
sQsYhkN+5XUqpOdw8xBAwj1lVA7NPgpntFuO9wc4Awi6gbs0XaP4pfgoqHWg
oBfAVpiEsEcJI5Yj8K+VpAZXqr5aFZsB/+kWGKSWQjjAhpCm7k+B8XzHHnzj
ocpmO4YIpkG6i7H7AFY9DIQ6S1hCIJ02CoP2qSQgRuKb1dnh9BhSv2fHOlcL
e4OR4lZvYGmAhzD6uyAVDwPXRWgAlXxuCBuEibsNS/jrxYALbA/fF+5uFtvk
H2NpCuPvDuZZNMhulbUti9W0PUo4LJA7Wab4j+TYbS4iY6O9eYl+8o6EM8wB
ChF4OqvKS0Idk4tf+FNZKkw0n9v2izSiaT0BTiW+PlD3BmilWeP+ZtYFIWKs
kCDloL79RlaHoBFQo4uQa0uM08rHA1mRWaB8x9km9VT5Dr9iHSGhPa3ernWV
wLcq3S71sC5J/D1Po+Z+cgLioUjr579pGt8v7wcLb15MXM01xGoGHVPTfuW+
eqDrMtxDjIKqVmrTT83lszEOsDrfod0i1WHG41xtmKS7vMykb0fWzwqySvdz
to5F/HvAN4eQP0wh0C2FGaKL3iw7ml/bH1Fyc8JSaPNDRcfz9ZfKS78FgeLa
/f0HIrRkDyY41IUqnRLWKnJp7dUXhkLOVfENNnd1m63oHu0KnPbWbRFyuaUZ
jm7v8IlgLVkfff+wurFVVWrawF+PeWP5GpDiLvr52NZiAMvYt0VQQ3ZRajBc
5ah3/ABRCLGRFnP8WCuIwXeIcKInlRFEn9/ABk+fOSh75CMgfAp8RddCidbr
A427O3pPtA5ZVzfw3M3yFQAxGGireGKkCg+gqflsaedcJhSAtd2k0CKrsmCy
J9Dmug4hxx/mfnx421/5lco09Jg7Gqqi5sSMw8lSiJiPyBaoRxsTvYYVzR2V
YMsSEbg8xdQLJl7eGH6IZX3VbrNUaYqWXut8i8mu04zjtVaXyiIWYplJCr/f
dydHbD2nwbFzOoR+XHkL3gyHkxdbHm+NiX3GJrnIY+NY3BxTt72QNp2Uu/3K
us7jJyBg+AAONTaXO+AFDgCrITJvKM6d8B9cZRVxMZVway+Gzhft9InBeFH6
Oz9GXQu51GHf+QgA2Mv7v2Ek1DeA0gvNm2EBYIqdOcmpzLXkSEZ18Yd/qylY
8ePs/Nj+7U5dQwf0VkNfwZ2F/w4P6FpkOJLkm66FA5Tqf/1veRK3qSqMa4vl
2+QmFuxr/jxSd80taaYT1dBq71nLzTA11z5eM8VhtYHQiKSmdfGHHZZnl6E2
dxvBf/P3ZlYlkrrO22kCcRYoeaJRKNodadbNQ/FdD+eSVIBk5RPB2XoktX2o
rEY85j47W81HocTXuyI0dfykL8zxvUn6rCGNf1EZIiAjc3T6cew1xArZSfVM
cRGn+x+ktMjEuJL7cD4b2lWVUxtWNgxzWjUVy5CNWOTZ6jKXSkoQLblYCS/a
TNOyeiq3TJ6ESu5KXiazc6mpvqT2E1UMorJAoCD20UVYWL+kvYchRrMrF6HD
Dh0ljjXhAlXuWsaYc9jsbKXNpDDrk1ClZ6NB6FuPcKRPsP8Pr7GOMjaORYfw
Wu3v8R1kVmyzPma3IB9fCU2iRU75g98NnEYJn0SA21PYay3HJV2t5t5LxT7q
AoGj2bMjVAcno2TbxyWBlsMH+Tmo23O0FL//miN28UgmElZRM8TDCjQ2M+g3
Yy/WVo/viUt45JK7LfweRxJl6Uzv5PULazJkN1wGSOJdNwmgy/WAhoPiKc4k
DMqlX/A2nBfqmKqeCzC9Dum4SII0Pe9sEQKm/Qy8XlYW4DzfMPdrIrS+zBsq
zQ/6nGqHpFmcau48jEEyU6jVky8/oYO5hDhldjgDHlduEGjBgZQ+e8cgh5GH
6hkedZ5mOYUyJrhNPD9Xi+wyZl26fFlSwsmSEb/Dl7unOgDv5fkNDAvJGZFI
UI289knErtkQ90H7WsqhM1u5WOvtK5aAnlJ5yXdRkZuTYl3LEEwWbLvDjomR
g4Jo8YX/7ueW7ONOgXA42Wah8+yGySYwJjxcYlz40eU6efUQJXb+h2DxF/mS
lBQwLOg7DyjD8oQFDnEiEDX38kMYd1bLvgy7jBzXTLSyTlC6hbL/AH4CnmFS
nIj5kCFyqUn0f1JzSO3JXvRGIWfofDW1CBw1EslxBH+TRXLymGwacTB3wYLN
SPt5GkRl6sTpalyFEYogzciepGccXOkvH41lK6dabEXclYuaTZDb7lniGbHr
I7gfkuNWx4Ol1g2VQj9zdZIOfJmfg8t/eqDIsh423drPPR0P760W9CNqcjxx
SFpdqfamRGSE6u25xc7E/o3MnihiHncjd4JV2XWwLoDHYQGdxgEwPAQA4I9P
J8WVqakSQcTpcA6XUw7/NNjjiYJm/hq6DUUA0vbu5I7aBrOFoegpjVtl535k
L9YGu6xF5jGhUfivtKowtQ8TrTfM9mFxLxbTET3jicJPi8N5iLmzbHuPCXpp
y/m/lFeulVvJx0l46So0wCfSmPiGTVN4xVg1FSNtY6G6MNoScVaO+hIQbhup
PvGPK2GHs4wjuNcN7E+cuXsrgQgDMBuXUbMWhSbMcNGgtiDYLo+vv7Gx3GEf
3675OxVfg3KV6h6vbn1Hd7M5QCjNpaepCTGnHg5HqxaGP/UL4Awdwc2/D9ij
k9+pHOcdq0Vun5andHlke9Z1iH6h7FO7J5WoBT7gdIIM9NykOOjmfktTLVEb
9YmCezNZyTIdI3lJ0Y1fKM+xIxfX5gaKZTAkK+CsNNw3ezOywjDD7IXsLdow
MCxHjxDaPANcvftMFyVxbAB8IvyprwjwyDXrPa5FZLauqgb2ggPi5d3YesEY
/LgR2IfRwwR0PYs1tM5pChnU1SW2voQBy3EJtN4C2L01z6dWHoyYiDFifmYk
yBDEha8Nd2JycoBTqd22q/cFSAHZK7X9GxKRQBf5iUNohvHLTsCo87flqmXP
+yU3GgZajpGpAQqeqbdhPSd9y0rcejnbeU+z/75ixr06H5BNayq2xgejJmiF
OArRoXi5G5RhKeoE5gkc3cixvJP2LpHwXlagLcLHpw4Lc1N+vT6BW+6A/oLg
OvXtvHwyaQPJFJIuepbv9lSqMYTq0ZhTJHMQmSfA9LpwIh6svoVjnFSKylgm
yzNfxbGOGmWKWbhiNpnMFK3hxfbTELU2MTHPYul1Mf1cRgpx+baXIFkcoP3Z
VIH/zLZpiCFI6ykeL+vJo8lhe7gBZURuBXrxwE99B2w1UzvLPHhHtQc9Khma
BbuIrnce08LaIIDMNfJjplRFlAXroOy4YoswTRZZPDcNIEi6FEIFjQ1kthgn
79zCHf7GTNQ23JuRgNUX0yMh26eQ/Ai40+Wv/9+PTHSWCUfNLGLFB50fork9
ELqeWDi1AXhiNfZdv7ARZ2cUpBaH1yEJ4+SvzXP9cqkepua2EpsR6HJAxXgI
3MzeCb1bEYW1d48ohxDbfLP3p2DlsD5f8EOQztqi2tqBF8gdIPxeddTyHcLq
yGx6IeeXPKcFCxvZvvBlwHeUrn+65IPgzjhjDcBzhsm3XShL+rDUOoxzY5dy
7nkMxWZdCpiz5qxybpaDU/X0dNtjP/8ObDQSm9bYGteKnsSDs+dYQw8cCtT6
pvq5KvrFdbUin3/ZkJrLbp/5cWEDcVLeDyZeNG92Q3j9mNnAYQNe+E8+qcZ2
TNivblMnx3AJhmLrAJNS37BYkSMImZ9jk03gCF5ljfq3OdJ4uT8Y70sZ5vN9
uT0aAfo9C7OMXzDYDD4NMKNhUtSEK6yrOwUc50efdHA6gxLgK7EFc06iMQEe
9AhkZrN0RKDg5/3MqckmOB2Hyi0LO19eq0mL0g2fMsskYpr7uvQzCnC8h9/H
WV8DVY8o6dXje5m8EMXa5/JcYuAFK83/1JgpMNLrFVRx2Y2/DfrHSPZwDqoy
FB0nTufDHpTFAXci3mx03CHXYSPtYINVlTgQXdI7Vf1YTE6muOTljtCzdQoV
NdjsW9H/OK6SqWWw8t1COhHbThUeTQgxzuJhMY+KjCKHAfTfOyGKVUlfiK6x
Fu+7/XLR2vAcXMuOTUYStAef3EAvI3X4F+71/lb7jCSJL5HMjdWUa+L71jLg
R+8UbsaV2FFWsf3uoQ02mW/zEux4EdQ32H7vNV3Ttc4/yZY9StNPSI01l+I/
ctZOW6sSY5wUDHSVRs+xGOJwtxwSn62XjKHItaLsedBPjYalPpdgq9LJ9q9K
mRMnecpEgmuipE54rRbtKq9DRIGUq6hxbWdiyueDCif6r5DprTtAjowlJ7jB
hQz69UIH1lZ7NPsesmFHJMk+S+0ZIBeUUtroFLyJcg5F38nTS3sJ8UBOL8ym
bXBNFfh7ZMOML0owd8/4zrM8gSEMt4pvaoTwfNghwxo/WUc72DCaHaKYlisV
OlmbsNycM9qLHF5EHsuGe/41ID9DiOiPQlD9zT1E2UzJZ8Uca+oGMEyKex88
JkkiP32Mv365nujsVXI4Kxq1LzhupKVSFZ/aWPtiPh9CbvHN/L0UEKednFMe
DKVHK0HoZed+CGPoSnp6fJEeslyCV29W5zuO7KIMJvAtQM2Ar8TG5ZOebG7X
rs3dAzbhvCL9CLmyFSnmfhBqAhMK6ltd3CRC/5CzdF+bSC7vEjHm11VsEQhf
hTKsVVKmJzWqgf9E2R+cTA62BxOwzMqgwglMMMOAwnDbuSBBaqo7210rvquW
49VHri+ncbGnxQweCsZ5Q1BUxaCZfft2iXeuUSH5f9/TNBgYahNNIynW6Xjw
bgFARY+RZGx5YYEhXU5mKH+KXW+OjhZfQlyKy0EWyGHKDqddqQZRWIXsW/zQ
itsBxvX0OtndeUBJkfMTXN0gxMAGidfJcOpCQCetRtTHuoJqNIcn6Mzceblj
22x/2e6rO/OmwOFnnmsR81DGNPpdzOdV5MJatlG95DPtGAmgpdLWnjb8ncqQ
3ebo5x+u6VYPjrPwmnyVj6OLldKgLQhpz2d5e+gUXRKeUOreKJPoibLp5Tip
Mshevph3WWkJ9X+hryKc8Nvl1V2SaPXoA7zQdAFPiWZbylZor37fEVAplB6z
r7QbMmWD/kdNLaA/IrkoTHT3fzrp0pnbXLNi5HK1jkkd/YCXFN58b1x31sTa
sTy4O3pYAEQDeUVNcX50xP/YdyYfDR6H0e+LNMpBr8BqR2TFZeT8ee3R03mX
QHrg0QOPm+x9pPQV//tAT6DE2ZsAH8peol5j+l77x88cTsQBPXPntgUItcv1
HXyhmg9rsKQm8LTzbemWJZpIlE97+6hhrAPXy90H35bp1dkBl+C0zuoojahP
C2s31k+QeafpWgQPfeCDY/tXoHN5811AUPjaiAOdhmZ/lxk0beL/M3OVLCn5
GDXiEbf8RsCwKcmDAb6p1EpFMvK2XJIx90VpiA9b630fDP2Z9JB33L8HxZVt
zmTbpC2LbSVzFmf/+z+xpul4xcnZRwS4TzdW5VRDarL05SVM7yrlUVJ8O+Tc
DI0DzndaC5uNPbBabzV4VzIrJzy8oZc0lt+msbRZ/Fp01T4oh+lMR38WsiZn
9vLbRctWTz3uXMUbahQ9XIv27+9pM5ziM01UZ+kURQwFIBe759dl4zE0Gmhh
6TS5vs5rsg4bQe8fGa2dJOqLKLs8R+m0v6U9iLZGTliPQLTLiPSssOi8KDrC
qtHk2PBsXHRwN3Zp3IzMHP14rMcXm4AJDtFpcpBqYPj2uzLSqHyzY6Rpq2vp
UjExDHXjhsb3MF3HhPZb0aFEO5RnXkDUWMIjrz24JWg1FJuckf4m/tfBFO8R
VOHA1cTu+CJK0y9UtPNn2Ea83bZENqheSnu7smoUdT9gLWXdO2XLJybJXRsq
TGSa7AfPKnN5Z/vhtZXmUDaz5r3neRp4cOjHL1iRDBhhmbgtRe/j9E9V1qw8
BMV0rbSbx5jv652AyeUM3AP2YUjPttW3DA6d7a1yEHTqeN2qf8WSda1r4xpX
/8IK60D5O9cVAlr3iKiIpNis0HYJbdQzPnqpD7IXTlrn4kb66rDCq4b2cDDA
aytq1zEDufKHHvZx7g8hfqi917zQgrHMLJWAJfHIU5AFct1BIkjNK4JhY3LG
bl9ZPAcop6Brp8aDSvkvM12JnxwGvJwWYJMoYxAovWS3kH2ND0rygwwCoj8P
oc6vPTRbp9J67x20P7yDk9wYgkJamMsO0p6gA79YH3kr4RtwCEwN5mbbBRHX
gRxs2ZBNodayhA1sW25LZcj0nQ8IERxTltebHnc7q7z4l7Kj60jgAGg25/J4
Mc6/p4n18j/qt+2jWj3KEok75J5VNWW2LLzKfKrHSQQ2QYj4aim8cGR6hZrr
c0phRtlYf+pYPo9DHptzwFwp1m9CZzYnvq9enARFjF4VyoSRilUhqdnV2ay3
YGHr2xQRXwtmkMiSeBRYfivQ6NFVpsCy2zm2jeAuIIEUztn6TG+GhUyVqxVn
obXvaPHDC2+bmcpvSBdDnnVV99PymugUz9N9L32JG5S/jb4vk88NVIpYWRzJ
rVVYkNeYdHR4QGCvLL4C4DJp9YFi1Una5ffG18y3FNMUwSPpQC2mtoN3OnmE
rEVIGevtf90cxjBknuDNXK4QrywOKXgLGC5GwvtsPNFSDG9m0r3SE1Jihnvw
F/7MW2WKWjEzr/RDz9IgthK+kZoEySP8pAYfwpWfpGrMUtMmF6hMCsIYEoLn
gKl0xpfktn/4Q87lGzmFOzGuEltNPRHxUKctoUkc6OGC3FwwrORuKq0Poq5k
Cf64CXowj+f1Bva8JBt0FpUe+M1z11JVHbiEh9jFq5958N/Y9QlJE92FrsXe
XbIYeGWvNWSxxuh0gf0phNr5+FPe3odFva/9C139mJB5xkoq99ZiWtiLl3SQ
MPVDWHGEVYEvD6KulNuJ68pipB4EoBr1FIkHuEgUr+1Oh4AS3mFlVCowsqXP
/AeWseJ8wgsRMUdyYEhZ8zYnb9in5Q6LJ5L22qnxbDl5i8l11r11WUr10NYz
/nsAVZ6QXxpRyama/QvRLakq/xg9ElbgO1SFQJzJwYc6+HstzYLFFoC3KJPt
dXfsDICLDS04oAqRYXIglZvwBnPgeG+Q/8MktlIwt8XzJQDCbnwJpLsNsT6O
9vM2zkYZ6PWk270YJPZ5IyA9CayFrfl8Ync3uQt3RzXkx9qgNdCHSiqCn84a
xKMOv6YurB7LtLS2lQdzYYGdGWarxAmOmVRBMb/PXB7CU0I6LkjHFXb1SbAO
IkdKessLYpi47vAa5pX3XpHNZQIwk80MgWLKAq3I8Suqw58zMKa//Yy0TiHF
LKYI4CJZYElUgPsFJXHi2VNBplmJHQbdyoLe2toRFtJy/lNMRFcBye7wH+X4
32akdb1J8MLzUugkDO8Fnj2fc5HwZYDQx2erGmHSXjWjLN0utSt4dH7gZ1kd
4zeqREy5+yMBgPS1l8n7hDTmMj8/HEWnbF2nV4lRzJc9v6H9hiAvfmbdzYYf
lXv0tYuftSiqqK0R4prQB6tj3a6GMN5Oujjp15IYyWhff80M0rwAhG2MKvqm
NRzKO+JQDTWHK1C0ek3yGndqYfe2bwvd1/olWBE1qtaWyG9n0i0cQiIcwGiZ
1Pc4x3HF3xGDDzhcWTrKceUDnWZXXQqcdVDXyyheRVvXDd25lwiM9bLQ14sZ
1h8m6xKDsV9Mw9o3c1CO/1MKlJ4Pz3O2fO5eWN4yM9nf/jgXMyIttrVHnNJm
yOApbyB+eDgU7PKLWOwP77HIjUZDVVzwq3yqgrHnk2+vkUrMG+e9M9OJgfho
jX8VRfLXQ9Y3aTLF8MJYsZC1ydQ1UVOOa1aJBCgyahFNxg3I+S5pmxpqdA1Z
J9TPPhICHO6CjCnbJ2bYW7cSiTNbx/YfroniYQP3NNqQrG6jDBRBFCscT1dK
b8pgEEG7NoxxJ5iYqyC+mGizasZDU5O5IfVaVRi520pGrOQ9xbv72UOQ2P1p
ukR1hDKSy0CHBeIJqQdpTV8vFIH6kt2CKaohBGCLmoIFbc9fkN25Z096b1uK
pGbIsxLyN3vR80VgtSECcfPC5L+7qh23zXV90xjuctDXMQU7Umu6E8j8LSjp
9xrFzPcVyN08dKlWOpHMBZBTu9v4UlCzMQMT2jjSEOsSlyLIgctqOmheuRXH
uD6rm+njE5tl1S/nRjul6z/ezpZma2ROFkt4SE/W5fhomNrf9LmAKwliQEVe
kHqXyP+m1JmLQ1PjR+NALoNx59otxOXstMPZBUeinkfMvTHKWzGhIVSmHm//
eRvHE1kx0yAluRyLmQk5ZK6J7mhrzakrC8sUK0hGcmBf49OibwfO4F2t+wS6
y1BV3NYpeolUPp0hrfobWtkUYmbDk7RHNjd1h9bpBXvLBD2RUXnvS0FFOddC
RIE/ME8VHuAF6tq8KejOeBbU1cODvnjIDxyZvMABBH3seExBev5EEydB3R6+
Jpb79ib7hmMVltGQoTpaVSwHpDgv9q6zfA0IAZMu8IPahcU0DR7w6XVno7/Z
+tSGAPZVLEcgXtCAlW+rauaIRFi7ElgnKS4ML9ebRGrUNmJ/xTjZEJXBfcF2
kS9yhInVIcyrWAdOu9LFZWtkF6eWZKqFaXAN7OXoqnmGLu8tY6UMn5YIoIe9
j36Iuns7pZK7Iv78IgtP9d1ej01YwExxcl6Ief5rIZPgRldKqoa86zERQ0Xx
RltBS4DWSrilPpxms3VQg9UuuAID4yW1ywJcA/7ihkY1ZlDGfF+y34rzENS0
KMm/dCcj8ZcipxGw6nDX6dg+WPOpNIWIC+ugqBYJ4BJr+xX0Cuajets7Qv2k
YDZ1qKMLCMN9L+GRsMwTIo/4l6DA1P3q+xExOiykrOja+u6WbSkip+TY7vrd
ZVKYVQlp4pRM56mUr6HKXJ1Gd9xYMusMDJVcXyLve2L/xnMMzKr/ZkZPrTeC
61XaXnBiNlN/F14Llv+Yl7AfNAdf6A3pl2XoVjvB2lh43G8WcgcmLXeFIHxU
yMvvqiZWMLYMHWYjC9FvBsf90XmBEMYLdgnv3M3l0pJ9I6xJJ/j+8/cFPfM2
yODkxFZNFOOnQeCGvwYF5SPBDyMFY07wBj0ipVN4Jf33+gaerppwOEZtaVC2
TsS+SpxVvxK8rOcU9aOBaQ1tGy0mygxn72lv60LzKMdf8bPnHGTJttE3BaVE
c8AO/1TLxf1Lhxn7tPqykBPRvqG+NvwtJ1egtLSMgxkL+GSfP0MIxb4wccz5
nOynUXamAv/NABu0G5iXt/3QzfhSY2v5nPK7VdVicWcuJ/2/h6l/iTD+tasF
S+IUnEpbz1loY/M0IyOIcjb5ZJv+FKiVfGGznoUE44t6u1+wXM2E5XfKbqaM
eIhoQXreiK+J/Xzb1X07HgBxXbF9PODe5LxMruPYWRMMb2s1SgI4e+n5N1GZ
UwwUGLjd3LNrAcyqlEZUHnukGBvQmT/JF0nbFVSW2NZa0NuyWnwlrbRdovVY
G5UNIqgAwygspS2nllVjSL3EruVdy0dvLLozD+zLF2w9edO7TpKC6RYAGi/D
Zu7aKMBnddQu8ZD7SFdEc9a75ibLRgv+WYwYDQ0V6gwprPOXIjT9xUltu5KN
Md5Z0sL8yS45hE2oJ57GwiWxOQYQEwxtw6er0LMOqItoU9j39+E4yEwnqha1
SXjcuRO+VqCPzZxvDz9I9kqL0Ot0N3qtRv0Qt2y5Co92OMIt0OMCvYjiJxaF
6e8D4lSmeMwK8XPTLuvDiks6+izM71tmBikoExJLg0jmArAHnloH+s/edBTX
sTuaK29tmoTNPW50bnJ4a9GZFPn3iopcGXxi/FbfFcfkXwTHpunPWVyd2R3e
zC4AFy/Lg27HCq5ylfSWXsNH8krPBTEJKMGpSF9hSYtYY+nua7dzBDvtFYJU
wiJpxPNp7ztiN06C2a9NcLeDKqVXx3yKI3XHr8Ro2nENrkLQ/wgAmg+X3ucu
TisFqzSELFdSqq3dstH0UIbT7o9rafWB36PB2pdDm39KxLD8AKHHg4DlcOQy
YGfqdJRlYb+9BXprt783UHl4qbBQMAQARONkwrZa62pYJUnEt5AId1hKi4yS
QG9W2Phc7BVXpLV7ETqsyFMvr5Ns5GIm3l+d1dtZheHNeD/c44G2JN3eYw+p
KWymDEJDjOWuaDdNRiKrLWy1l1o0lzRUtaJxwTYYlzZ6MpM/acCblDuME+DF
j8dF5U/8qOaJRUwbRSfNOsH/hfOyeMseIssnjfMfAscSs1WhjFtby/xzIcx2
/+q6TMXW6btf7X0K6vacJ9C9AJ5tcPiHOijyfixPHPtVXzt8MdheWPLrcaF9
j0gtXYhXflecFXIz3SCQrmlpqrMrK2QKuc7LNZIjnIjZhDUKJ409y0GYTvrK
IqjMO+FAouFEQftGUsKmDZBmYwgzKBn13kyWv499BlCawBZplll+ea3pC7He
prkHFphFyrUpk0T7FG4aBfZU8hV1u+gVk26jY7QDjfg0oqIlOCTzDmIWVdfN
oLsGHA4bvyxu8Gr1zj0glp+HF4pRyovKFf9sJn2ih4CMTBgJpTIBeBA1DfvL
ujiou/QmQnrkDbTpkSAgHLYIRAl45jUZN6o82Oc2MxOr0sw/tR36PvemT1zp
tHlT6HoZMRKtjs9ZYh225chvcccSaWyMLjO09q6Yi4LUUb/b//LakmwGwBe7
tru1G7HNaNyDIU7KEZ16V4iwCYIL7OlTDMp2pzCwwD+6yo5zmKzSTKd7NHVb
kjRJJVHf3GFIGRtAyT6p4vh6my3yk2EmLhzB8cYQMn5ciA755caGdfzIhesy
lbHC81ZiSJ+W0ANbWZiZljxPvG/TX+BNYDw60KKzLpKTuHunn7rW04mIRMP6
gpUnLOKxV8/Lq+7fA2PazdnaiifPEV4qibWzk8xaGoqQhv93JKI077a8SMQz
M2MO3CO2izOO2ff+kFAte0yOVlGhlRxJ7jXGioMcbLI8EpxPU3M2uGxKFMIN
spYeGRzsUa+p1pELA1pxWtBFDDdGzmD9vi9BDehzDgibczSruupaGDoAECkm
dDbd0DsZZpJdNd+I5EFd43g/hrjj6bA0gIDCVSnrFWI7FOvGkt6/oUga6OoY
aPCjsycBr1sOrT0zOAChR2xm/sO3gxHqmCJDelDUdefRDr49BiaEV0zNA1Fi
Cd0uzu8+StmhLFmCF0bywyMdKPrgA6VNe5FXumygx8457YttZMk+ObX9KN8s
MY6eXqmUODMzxm0vYolVLeU0jjCCOpHT5CXj7y0J5HMNuej9Pj0B3aJf4asm
DP/cBbIbxQsUnCJl45Mdvw1BxOmzaMiaqShtsPlwRwgXpvb5bDaiGqOEfiHE
I3mtCE7opaEQ9Koz6wyTMvP2gGqKDCjtAnC8aExxb9vtPaG0F2QlNcXrWok/
dvqPE95brDMkrOYLE76RXjv+1uuZZrGVcqKtosUZboGsfjWVmjpExw0BmM6I
WzuyeN5Gm/K42bh4xjSaEtkMpWAA3VzHCMjG/07JfBnepv+5QLTRQ56NpH5k
ZzMus0g4HMcfhIEAc4nIBMCr2JlDBvAM9oSmU8yz4wjJgG+iYcZmqqoLVw9B
EOBvtF9UCDcvntaTArFwiWrfmayozZgDnWftgN98ToaUQCDNJ5CtAUgqw1OQ
/7oQikGtrl+sAGRvzsrJTxjk8GFGGv83y9KgP6RB5Fc/o8wCaMaeptGc8QNB
RI9jG9n8S6bbqOBtdUKHgfMn2PF5AsjG7R/N6YDXtZKb1pakzGLO0L/RAQkY
sxJhK7mYk+VAHOgULmRrxMliX3aSQdkaz/R/yb/VxSKzsusJoil+SfpPnvoi
zrYFhagUrWmn9OsDKkyiEHetAoUyojN0L2BfVQBYCH2ab2kCfO17kGcg++bV
ne6OnHnPUeeyU1dnGIyr1HDnGHzlfuLQwny1qZ7UpQ5/y134ku6ebEoJ3w6f
Hn8P+KFeZ39auEgmIxJrt/SmyscWFus0/6QcDDfJPSxUtFUU5CqrGn4Wp/j/
tkTc1eo40B7X+HEm08KwQgDf+CFOJPrn+wWNWFK3/jQw3J3R9LAuQ34JJXUI
i8jB1xDMIs+bXj5Mwcwzv5t65EkSsgUTvKQnG2x6R15JgS6Mer3e4N0knYNt
E66pE6v3bxFJikxl+ENEOIKm6nKGOBJ+2ixJ1FBa+dUH0KUQr6IFoDrhJz5c
visM/V6iiV3fsZkGhG+gyJgIFQ8EDYW2RLAB3UqpA+SHgJs6LVWVnoDXF1KN
zchnoDurLszArlRExLm2ziLxNH5zbIRHjTdeSRFxTiY1zGDh2tEpSqWGNbog
4ARPZ3uHo60huS/7bZBjCExN2sbnvb+u9ui8oRHYN4nT8U7ufkV8gYcJtFOl
Jpr+LCnsONs5feKIdhrmajbTaOTkoYgKTVip0eVTiiqqa1/RvBGZcw5w4AZE
Fv1xNynUTB2288z+/kjP8TWqHm9vB0on7yboghNDiZKogCSeQTFbZZ7r4ZPo
1NJxA5k1x4nlaINqaZxD4/bXIdT21CcE5ABXDIX1PJ3mqjoXoDBGRk8CQE4I
ouVxCP/D2qIUeWrgO0E2sj8yfc/Cf5ZyKVCjp8oOtk1DuaM1/FKpRDihRuOk
9FnkQhM5UjojUXqQXG98f9rgYOg3r9wqr09PG269FmE947co3QrBSc+dm2ci
L7kQxlsbozqDCDnYmC5PDJQVFydsryR9t5Dr55M6TDCs3FrC5K74ka1J6ixj
BRNhwJgDLwi39YPgJ/APi2l+vMckUGZvDXpj95gxauQtUoIhDYf+d59iHGT5
Nj2KnEdhPMUMhmMQV4xDGGZGfKAZO+IASbqBLbr/xGzVwJPYwqUBZ49z9YHl
7ZDfvF66SNJ/VJWmdpQAimsWH7hcUqYux9tVn8T3BozcPvVTysctwNxsIpDd
hoduxp4uamuYdlKLoEU5NDTiLRKuJdqJyEkFSc8J4WqlxUi8JbGoBCjF2Wpw
Zb2y+HuDJIktGwnVgKulqRF4ei/lL8y0DOkxA0b26SQprvCtCGHGo8JYhG2e
2AygJXouaLxBxdfpfz6CeU4bD9wDic+gCO11hHnEjTFsvs+k9xFyNR4lBj1i
SaQvoMpX5PMLf1HLvhsMjyPiumZYW2cyz1MOARfnisn4+8g7fZN5KJcxpPsu
WfBV2z89TZaMAYjmNFctcg7f+K5ohvWcZyIdPu1KxVVXgfjNmTwtphoJ/avy
EzPX75//GzGAXGxxaPj1DctPrqzwiMj/sOGpCq4GS0VgTRzlS/TypWsuTya6
EX8SHJvWkwz0fg+9Fzyf2MmJ6/HAQDxQccYlnAY/1aFfioX+eGTwM9pxrHtO
gIq6Gzn7m0LdqBp3T6Sr/0zcWyvV9NQry+ZfNkVFCsIiLHQEPiw5q6HPHNy2
YAbSGwn2Vp4ZvvU91XtjDDsBwYudI3dh1nwB5FuG4oj3WWZ5SN+479ETksJE
oEHdVJ0tVkufW2Q8ZR55Be6pEjFB5AF+/b9LjBvN/yyJn58gKrvfTE8DnZLW
8+usOQFQmOIEZu9GSoqNsDqI9tGMbn4irVdpZ2esQe6cr0TZyO0bKhafRlBl
vd+GxxMegZRzMWwRWpcPYNHocuDSX6C/O61rJtaV4E292RrhmdLQdRrEA5l9
ZMA2eG149niB63kGSxuILgba0LsvD6jU+wheNTl7EnkrxTbXIyHv6GJ/g3u2
LOFaPsA9/7TpDCyBQQnP00c8FW6+6rZK0hXXiTCpnIRa4xm15xYzj4kKD1Ov
j4RJy1RkVPO/qmMKIpOX7Czg9fe65x4lsA5QJ1ZO/XsUUOJhhh8XAVrnrdrD
ZuC/dDMsjUzq3uqaV3ct8tkSD1/D8zv2HuT0YsNXFZQDfeu0L935GZG77jcO
8YpCf0Puvu7L/kSGET/Go5qgLZL+USOsKN0LXIVaVvTG5ehr3+fz2VHFOu1J
ZFUiXPUUdXn/ZAAFAXDR+XM0itGhEpEiwKi895kAwY3twAGy92d3eZWHrlb+
dTNw5Oe6k172uE9Z8j+lWnwLyo9sz7AeAQzO0DWhmXsoL5qzqmARBRLo70pC
R/MjV+72RTcuY6q7iqtHI3UgCAij7zuAN8LOD1vUTnk7c+3POodMtVm1y47U
ynw5MoRpyYl1uoYpYUI9RWKs2TBx2KEK1xZg1KnvepvxEcvKXaaWP9Vo+4GJ
5+YtCDO4sTVIr+dujslSxomjPB64xX6rXcOPhJom4PcBtBHrozO1ik05QSLa
igXo7mknwVWILOcAbaIZSXf+kZ+EVUfClG+WnlXTxkW4Urgd2UuJzTh1pGSh
+/92dFgirZ+Z6+dU2AUCaTfhuj6mGKCkjwrCOOR2uFH1HPt6U2Bu8RDuhtKh
wI/KPHmANbiuQ6BZSpAqGr4j9lfI/f+vBbXrsTaYCHoPHFdZx93+G3+XCNT0
68orOY9wkAzw+xQ6JtObm9d0uJzh3oHg1Ospu3M6Jl8YLB7EFu37cy9oseg7
uXSSxLzHK2P5HXaC8DeiTDoWAeebUdEPMywHVoqr+oQg2SDnDu2JQ56lZYvG
DnHmB+lQ6cXFowLoxn/t6WK1UEjHfyEWyLA8eKEu5uc9KD2tAz4pv7uYGGeU
ehd9dP9KANtXitooQ7F+63KNQUKuSkzG69gZ0biFwrVOP1bgmtU78w3IOJ0p
n/CamPWBPPeWicazm2t50C2g8OYgIm74q2PdHRkpuUMwMrTEwrMP7ohHvMU/
8hdffBL22pCi2BjLZbaOxxinumO1k3tMC/ddVjwHtQjkeGNwCr+2h690/ou0
JeSntg0ME7thxXFCiqBjFxBD0q75vGXcQE1zhwv2FttMGOH0B5W2zmv13UJn
VDDznRkVpboz7vJ4IOSS9IhtTb8vvlhYQMkVP5KVU4zpg2c3gEBo4i8uECPz
S1lISSZqmyB1rrL9wq7btSmv/xkrcy2FXEjMVQo/DQUCRIDyUZj9Z1icm397
h8R90OWXviWEIW07UvpGwb5RWgFs6SX3VNtZllyvxM65JMBAYVh6NkQHBy9/
+3lLRv2XBFJs+onh5LwF5Rcne6KtlfCtLbidIFBNg5H6oRPlUnzIWTKUbf/E
26CTvNJO6+Ou6pcJLIn5K4ts+vBxxeLK7aTnoqqDreVLav5Y0DJnzJnSTqaY
rfAr4pHF9V8t/S0sFzyOcjBTg4Y8eBJU76F4+SAccjWa29NuPNrdgeiIk9FP
7PCh/hFl0wqd/aIDkBF1VMd2JCOjJ64gGIa5Z5JkVj3OXLWUQKWt6ldkYx18
OQRlaKcEqW3YX+zpb031edgkJ1D/By1SXSru3sooL87FY/TZEPVTuBSHzRcx
RnY9mo0EjZ1cCNW9jEvqd7NsdoQA4vXWQrYfsAXFhCEtz3EVKS0EGQMGtA6V
Fs+CQWosk04lyhmBEYICWElmJF500gHBZb6jho6/eCHozuLm06R9GFMpXHfM
8NyQU3CidIxWBVzTJ+WUi9uXaXOOfW2ayALd2Xed5blS7KAQy3gbWECXSYJn
PDmWlGkoRGGOuImV3s40ZXX2vdzntJ/xh6ZdB//bjCLjeOzJj395XHOQze4T
on6XofhORutw3YdRQGHfb+PloFdcn6ZiTzKp5R0Zl+0UJCB+D60fhcW0Hirh
YoK2CEE5tvT+A+cnqvx0UZ/BvhRuYa4Qnr3gS3FyUlqz+gdl/TTqqMg1P3ZW
rpxPwJXcGGTkkqOEOc9AnE7ThDRmerZPgr4yv8zt0XG8GWUXJpxa7J+wBXrL
/1RG3t4MnAq0eVt3afpqhdsDCcNyQeiobSM+xeCe2dWmGxruH8MFqVJp86IF
4UCSD3533nRi1zDUu3SEW0LHOZLQGWRathRcpicmernkMRnZHXwtz+KMKkez
3GWsD1clQ3DmcyLzTgKOCUJlfBdmvW2S4nLKtElkzNFC+ahXgOE6Gg3pvpmW
OLyjfs4qWNDA6OW3/HpC91+yisTG/3J/XnZ3PFQRPG/86CMZVbkcUIckQJN2
d7jHjA2P3utldF+LxIhosuBCq3Iwb0/is6u9rTZhXh1KhprGa/SYXKZTKhNR
J3zhACyf4PQTSccmXX3JAlajBuOO2NUkQTXceEyKl3wgyDPfxBvgZJxoYgVe
Z91Z91FpSvS5apxjvwzjn+OtUW+Vz2IGG5WW9oZbZm1qbRo0PTHq+YmSwVz8
5GWdhKlDTjoHHbZew4AJDmex2p2zv0ZWpfjH1k+cbKXJ7gt2Tuov0mBByWVx
TVQ4EcuZ3TQhA7uQx8Mot8beiI0lQK4U5va5t6zcBiueyZLnb6r5agtosMvF
kU/xbQMBwYJwDmSqaEcHUjdxPcyz5gcbDF3aIdG6iiF3LcjF6gGef+VOW9o0
jSMFyr0EdYGGTFsbWvsjSzl8ctdnf3ZYSHskyJXmjO1u2Gexd4SFstoGBa8C
tHZKRN2YkaENZpDPX5Gu0+lp0lHom7+KKXjSrMaa48C4Bv1xwUnW/c1J374w
D59p9IG+fdcvac0gERL4pJRSNjsnoDyiwJSb92/e6jUEsZ2fB/ihnI/69r0/
3ppVUxVCbTm7sluOBc72vNlXt1IQ8undndKvCFEUGvySTN7N6nRB7rkMjYlk
2OSN4U77GjGPpcu2H8Mgzxq5U1poCRfb9EPpZtFyqtd0HyLspfgQuJQT43dt
StIw/M0djkQ5invOksuo2MoBBULeLHYr5bhmaWxqHE2yN/P8EmIJL6lc3t1o
lDfFsUws8civ7HMVPrB1CWywGBLQQpiV663GHv/CQJR11djkL7SfctQyqQRv
tjWGduKMlzyXDTVtWZAQVW4ZMJeBS3mLyXg5klFsPzGCVM9Bklm4LH8aWIDV
5OhYNmfjs6wyKRnAReDaQ8XCRF3v2Q/UT8AK0qR42fINzTzEfdX/xgzfBjxS
XrnJrvMBEwOPcAeT+ijO0j+km7RteGEPP6CBzZsE3WuaX4LPlscL3gwk3EKp
OBcPRJeBQK25GsUAaKuWC7HjLauVqbtLfzG4rfBCR8d8s69QGVqbhfjXUazb
PUPHsofvERAj+/L76HJdgwL0/PCgFy4+gLl4J8tOr7ZrOkU8TRYKYWrTbwRX
309bJO38rNt9Ve4I4UAGm26KO3djC93C3lPBp0fWxfXFNYUjQ8A2CYiIpF+4
IB7Bj23WtBJpEcpUm9FwghdMBZ9S9dvB361qEwGq7xPEpxvoaNInYMVnBeCm
+LI/qARzVqZq5EsqgXDRK/LFpGpbeW10r2DlzoZchrgrEeUHHGsk6HCssK8S
H5s/DPOY8tmL7j1y486e8CazGGjhjUcETVrQQ5pLffEgxofniya4XHuRBLFC
q9IxCfyODAq9BTfPGxE45cAwdsWetbJXfJH0n4ZyOFREF9alkfDfwDRWRI2O
yPxQdk2SM1sCyHK1Ouk0ooLHQdbI/z1N9gtWPwIHp/JVlt+ZHDSWTnQlbbBw
7xrNRH1945D6A5vAHBZze7fVDt/a9P2L7evBs0jTGLjLYyE6mDonh19QOZcZ
YWaM+1yHjcdMJlNvTjSpDRyv1aDtYsTGGKTsD4icx8ZAxKJFlN9tv/yPxVyF
5jziGRMwgtS7sofOs3BIBwubvgohNvg97nyyj/mbcHkvK0UlbXh6WLRV9Gjg
77UB/1+yfi8e5FQhp3aR6OP9/SPWFOWLxlUA4zCSSg3ETC2UQxeJvNyIT2WF
Z8EtHoT+FFuvUEz/H+PhWcPSgSaqzt/Vm/Kokw52mIIA/qUyg9yBXGDRy7nY
rvms1a/BiVRJYLK6VSXzqsAvKFTq80MGxeMbtPknrCCg8e7sjHiK0T418H8b
OcM+3P49ld57lb8k2n8+yeoxrb0nZSrQl8mOMAJxVRqGt5zmDztwfUvpoNlC
IpIrFDc5Dembn4HCd5X2XKwj7mZMlBjI99e8VWKLx1WvH2kmAWFCD9u/qMJm
GkQWlEfWmZ5ic0HS/CAM688ZF65AVD6tC6tToDfmI18ArWdpZ+HMugzRUNNs
IQipLQw82wRgB/MJcZqdqlZYHzCb8UbBBiwOxOIabsPfGl2c61RR2UF8ujcL
q9ki2C3YdQUTa+U2rWwKOuI8x+WSm2x3FKRR5Yj/rl8ObNP6QShFRR6m2ohj
QSIul44FlTj5Iy4y1+QdiLs+E6oNDekVsb8YOVbdx64SAWtJbsX2ALxVALyB
Fxcb4N5iscoXS/cm+E/r7LbnkvjL8GpW4U9M388SmdA8cyakNHQB8dcj0OrI
v+eHxISst/QjoegshHvEA8KnKb8bRZoxA43JB09F66+owM0Rf+QuOngh9vzB
HYgYCCFEBJtyDHqt+K//cxq/hgFfxGa7tf6Bd7KZFGWfLJQ0oku67SeB4lsX
d3BasQu3CwA5+qnohZEEJJ4ZyRouUZVCtqpX+wxGVPpHVaX47FOOb5lmac+r
LCuD70QAImB68MaOXnbzta/xG5d+XQXalVo4IF00fUfrm2aqXa9tBflrjJY4
PKtXEjYz5BD35c1A9abX50JcRJENBpHpF0vt2J65lF+pO0Q5AJgKRLUw5mSR
LVpsE8CAkwkBksbpuybQ0YXLpBLuv6xe3C7cOQOeVOEyLOdrvzpVAqDzOeR0
XR4OTLsBUYkeTiDhj52TpnYjxxUMiC0/oqB6wXMHu4aDseKswSw+vbJTmsrT
r0QnRp379W6ovRCrTS3LwH8KOxeYdjG5e7xEr1NueZynsV98D5C1xxjuGog7
lctbMdSBuVRwssMn2VBbI686vvspovMe11bXtRuHabaIXzFBoKbRkwbLIqhk
Hv49dY4z6gl0Rz92opXcuDqiST5OdpgXA/NKY5zVrs3Bgu7mmQJO03wrwNDB
/8mYnUpZrEv/MQZFZhw5V8vdFvo492C9PI0gyYxjlj2FWyFy563dOJ7fm7N0
l/+X8rlcTSc6qgbFBQncVN3MZZrMr6I+416ARekFlSsvly8nSBo16l8HCVud
O1BXQ5FlqShcUBR82mevBuLR31QkXfAi2NjL+1b06fj2zt30JJ7y0yB00qgN
ki0bNVuEwrBU9BOqeHfzVb8yGFq6JeGIz/vJbaV0+BaO/qA6IpKEOgDf6GIW
y7xzet0GfXZbEaonlvD0spRnBifOTp5BrWFdDvrbHOR6XXjLyUxZZtNySgWJ
UaH5mJ7ps6gzQbsRI396nnaTlgHUEdUQeJ6wpK+TaueT1d6fndLsOABvSUo1
ONiNsd70zYC4AlQ5NBJt1g1tI0FErRkMcHMmxA7wvSLGQkjT24FTsUCWLBEg
AcLS0SLmXOMvzDaDHPlQqE+Vs6aaJuI4Qq/F5OhktDC4BFm+ZAsVbPaC/KF1
ciZ6xWl5FS6B+svLL/34kp0Y4wQ13bSzWJvWesNK0sJ6HCHhW0pXCmg8OaKF
H/vMg1jfceX8KKX/xN0wsPO7Yl8Vg2vRwYt5cSzzAA+OMfvGW9ARZCxJTirX
d2Od93onETaAerlIZIQ1cooRHLuTufEMYox6u26fI8CKPPZQn2dpPReuzVq3
j4n3xw2tRoN8kS/3E7Kp8Q+5CNZ0bGIKiU0Ivp1SWytpJcyNDWr/xE00wvqH
7852ncI+6mT2CgknVng5AANPSeT/smQpEpafplLVAr+Q+3NuV54ZhMGwgYbU
JrSCF1sSETCNQlPhJlnI+/zBiFk2IGbVPaXabola07lAiaD7QKS6QR8BdITP
QoWhkEMmqzbVzqodBxbCoJJSzJtLvceXIJNJSGV8tGkijVzYSqz5A1EA0SlF
Sy5EbVZk2jgOa0qJUb9y+RRP0Yy/iO9A+uMBLuQ91ZMc36j0XQJ4ZEcuNT6n
S0k5TG1Luy+X4seTScnzSpAaDeCGu7jEVE3VDftDyszfBAsl4fTw6sNdZKOT
gUJ1YWps65/eWHH1MOsd8mpOIEXUq68I/RZywvLws06xW/WBgjgyBbMZrBm1
HHTFFmo7p85W6ReIxsS8tx8nbVjoP6+OGmkj8bLxtVTrT0a8l7W03doKOhl6
zm9iHNSHytT7mVzVqtt5WqxEtlg9xcl2VIuDElX0ScK/0YYS98NTBXdLTqx+
NTs+D8zIhQpGpr8tryYCVIicZtRVDkW8GICIJNpAaUJLmdETn5kd1jsPS4yO
LnlmYh+03q4/pY95hOqadgfRzGgjWH2jaJMH4qnMWcHctFp1MPOrb2I0p4GS
Dtk2u6v5nSHI68nrNGkqscj35NTndQ2vkDSaolrcVmmraBpUpjklgsZp8olb
hjmSP4p+WRvKOM217bNHh6sJcysaR/tArVDTqOyf6qPFEgj2iU0HJg7YYc0Q
Ajk+IHuDm2hSGVC98/852MhhWiyScdnZZ1J0OE9fHdZy917sucmMR3mPYyzU
te6ow9AjAjN8onJo5VcvzHLoISk5ZNmMO1QQfCSJPtF9hhutUukUbxqIfTID
RELoUIVbpdtd5lKvd/k35k5mw6FvvCM4UIXT8Oz8keWwWnH58u6jvZ4/gTXA
DqeJ6+WHkRSlx06Mo/eBGpDeqRnYE8/0kHK2c0ALBPDvdRjd33hG2WvQXgWs
cZk+iuDPQ6x5uYNKbk9a22fe/D1WV8FlGG+AcIqxIxNJCXJGmz88fXadh1w2
lHYFVtHroR/Sb5OJEkLsufoogK9gMtMnZPWf4wYRZYiygW4dUZ2dPniiTasm
z45dfWJOlgADoTql/Oag+pRe+zDpOXm6UUDjhOgwUSwieWHZw8QEJN+/oVK8
MoJlelVoCdsTnw+TRfqU8y27+wbDVfwC1l2O46V4HBBef9sap9oJiMQS+84z
FvpHArGcBmhAfQwSSKvd91VFDePxO2G6K+4p2wvFtY1ldct5Mje9KH32Tie6
B0tJ/ke+lPK/RDqNjJ6HvbXCz4jAysU8lhsBEPgdHDqPmcAlDfaZdnYO7Pgd
rri3u/KMslO+5zjaQpzNWCteCO+TAK1k0v9kA+l3Ox2Fjql+vCvTo1MVgnc8
/zRAn49jwLldYmhgDflHvUKOVRbZJme4z2RT9n7Q210gNluEyV7CAGQEO2/w
Gzm3fqplQzjPrkZS2VA+jtu0zZNTQar6KoGFFGNrLPE5Jx1jWiFY2dz4494I
iUG+pf/O2YIqQ0RL1LbMBSs7nIlA6EhcEUplPiA0nc1Z+tMz3+K7b6IS5Fag
LOwJvOWp9hKpEbzFqtDxFi1PR+kKcmZWwaT13Ygvab3Derzd6tLqC4vHgxFa
a2GwOvWOfcAhYhvfle5b2BYKP0bmjUjxmnupwYp3ukuvk4B/9zFl6/gFks7m
ltHl5xwjdGMpKhf5Qjc7Xg4irR/jVZL9OhuzfhDBtOypqy503WTesPQRNFCQ
UDnkDfHCQoXCTYwX1dvai3vkuSRbPbHNt2lw1Exo9mt1U8afSIIOmucO2mQq
HYz97xsyfN7Uje7qOoah/lRoisIIFDaM0r0PG9zckaVqzQNb/mP5a3cjPRxq
9sp6EFUJfIEvZ88I9j+t6GahywJb+2PQ7PYrK3II1s26sp0CbWgtHw7+weqN
Z/+5dyRPVxV+L+hc6n89IMQryI58VB8iKJMVcCWG+4y37pdJkFlRb6ahJOp/
jVkCqSFvYwMR0Dx0e3U4bnk6FT6ktOPGju4VrVw/aU5vCVIC+bVGATTVYBPF
9dRl9t5ZtODzHztx8JxIqhkT023vhijWXXmR6JiPJVweGoVZOx7yiiVoladd
RBYsMWsnX0wvysNCm0Pzr/MttfSUM85+k0njL+VCpFufKmJ7JIISXIbSHYrG
qxdUiGA8r67cQsllHAY5wjb83KIw6+mGhmYIxcw3JJM6DqBXPdDywRrhS5xo
uG7vsXL0F5meqwDZ6ZXB7IZgzHZN4kdkvlb4/ZiXsniVfjkWgpgkuClhgt78
x9+JMdN0NsJWhOdpsMa1VgfJTdxEfWUf/hCWe7cW6kF1Dz0iJy2Z7/3NNVYN
xST23X2IWQdifegjS0pUNLskhzjUAIdBTbqBdILd3DmMKBi4yY9VXSWoBQhQ
kmXDIt3EKdyv8Z+AyzH2k+s6OwOvet0ULgPoTCEpYiOAzsV3vBsC3eHIXTJu
AkqI0noJ2o/gUGLOXXI+Q2P2CKvcC0dFRKjxXaoOdxcgg5Q+weRDowyJPIMn
4WgzTWNDpK+NVHveWjp7yMBLhqNv58q5ZYCs4MpTZWxYkDySZIbaNapMhaCp
p/qem7KfRZxlrvaiPnchpmKwOtGOsNJINMvyrDSqT+zD0OZJACHz/iMYGnIX
DJU68M09YR9KsQZNFyqj46qjKlJMMsh9g2KliIchIOKu1q4RFjaQyo1OV1dl
SEM/wfSdW0vpJ5ej59ml1o5SRj/wc6rkUT99rbNyHD2YXaQAVk3Mec7nY/dM
G5TNdJQDpvH+bEoGQtXEF3VvoIq6zgEsSPltsbx2KHCjzdzj+lbs1tE5tYYh
nAMu8YF2jNTU7Q6KzMBt7dAU2mgPHeG/ctW9i+czccZBVccW7NEc2H1esW+l
MTbK2jr74j/TqVMR7oxG2NDrlKfXvnragF71XrSLho9cx4AqhJlMiAIMpdFz
o7PQOfEtjCr7HVNVDZ6n/Uk3b9VOMidenIzdchzUTY+39+FkxkhH0O7gNLGl
IRCKoD0PAV1GoGCvRXNOZmRdXw9ExR2IU49Xh/wrdEXoIEoiIi4p0/yVH2XR
NVRDl5QhD18HOuDW8/Qmg8ZIhT/kNSBerVfUo9qldC3MWCkZWCCJx1OwY2ej
/dCgqiZYAS90F1cllnUlOwTLPUhlMF92GmWmGq8LhhgTMH1Pc/eKA+UfCO7S
JmI96nA2DN7zZweY6HIBcp/G1y8lHlaDmD9WoeuV5c4uLA8biIHx3y0pcR2H
CTalFNQMY452gS3egURHPQMM8wPsHf1/gvJP3sZRAzqWCpsxYN9p6tF+0FB0
5dvr3z3hURa1hDnNcB0SHZayFW9Iq04jMp5RzlAKowC3mgeV12XSQW3qLA/p
BkUd2fvuWkSfy8r0bbP2HXbOWHFqP+tz10Tm3AKQ7c4Wz07/r/kphvqp2+Tq
0sDAsVpGNFRtSPDzwCz6xdWGyQhuMpwHm+905Cz62nU1XZhsCedy7v43rpn0
jP0j6vvCzj0/L5tHJI8BrPPzWS37b8MBCok+Np/WVWGBpcWpsMuG8ty6uzpE
uh+BumSD2KIN17DGZxjcjPECyrCrGNN9unQWs61dej8ljKfK217GQCQF+xVN
WlouOUXyvu1kPaV1appxRyeZbiqQ7CXYcU4XkHVlFgLZqkoIKPQZMbNH5JhQ
+VnBo9Id5NYCBNxFFdvPs4HG73KKSxNLbE1ja7wG/sEbMQI/HkytKxG+pGQo
mRTe1AgeKjaTQGUvpwdMA/p5CxEC5yf5xVstWYtQpQKDO1Wdibty7L9iAxFA
3f05flR3rze8hT9lCCA6eXqNlYfRj2tkD5hp7VlqbqMmGTZXEDgWPLmYR7Tp
4jERqJcap/8nqAokB3WuX23f/pdH68lYiA2kzLk8xa9v2H9/6pfCObcGkqyE
Y4uf9SCKIiw33zHxyAyTWQNIvnIlkFvqoesLPtJ4+dOb6HOsJ4DHdiNAP+L/
rYYAO2egAhzLZWv+oVyNZhIxxVD0T5l3X8RBac+YjmjanwDNRjlHsfE0eFgq
uay6HAruAtrZFKjYjSXh+jxvxnurO17CQDc+0g0h7pDD4RvctttRNY4saGMz
XvcEgTvgmelSdKfFAQpSsnEopFvM4QIN8qCQu8DThlP1LTluDc163TXqNPIp
fmS7Hu2Y2K60N2pRvHKz7hnDgMiDbGLwvAkwqKS6r0m4YI4BaJKWPtFXeZtr
AJQ737PHsEoa3MS4Mzy1jDN9AAFySfhyku44g4/WOGI5tS5kPavtk6ngInMJ
Fhohxnwxl6ir3KBXzG9XEVIN1fv8XDN2CfZIVHxsgOOtv6BM0sl0n1imhJkr
0y1U9A+imtTJX+cJAD54onc6ikoDfuvXhhtUVfFLHK6YPpErEKWcbPqkE/sw
ieNGdf1cJxmfULq9E4dmaI5+rrMbDL4xv1Y9/n72tpKk9/Dewd9QGPkg/ATC
m2JAWCgI4gctpFQunR3r1BmLO6QJTb7FujcpX15MZFZEo7V2wcNi16SsG95n
+Cz5k6QaoWHC0428qLMjgEwAWmHgXBFS46rAb1MKxJ1CgyD/slgrzrR73gNe
q7zFgnXNn9T3FBeuNHo/vFzedR52PBHiF9NYi1CN9/1vKI1xSGpR/S+NBJtU
a82ewrqPv9lav0cyZSlmZLIGbAuIUjjsB1hFOmnOZkQfeScNiLe+Rmc6ll5z
+a8mZEr55Mecs0R0V47jezjyQLvcsurKsy3Pt0YEXy/CBuT/pHr1KlcSSSGd
BKFPLksHHgKOTmkP0VXG6ZlxLB7L7xWVfn6M2H9a2Ys4DIfiF/i7rOOZOMjN
JAwSgi+EXw8bFZ2ogggapPEJavTC3Nbt/MswXPx47h0PGX1VRkADFiq7/SyI
23KCXchMI7o9XvUcAZmXh62Pr/ISdYf16bom1R3X5WdrdDwhK3q/YdKQRENc
dFofERnNZbQNA+iVDAm5958kpr1EjOAFFr2YNqi7FbEIzgi1pcwNwVV+M/6R
jz16G4vf646Ip69WoZIGfNqAXJwWF1EmyvhoZabITvRPJaaVoDuQkC255gVY
3fyVIRxsKG1aD9QTlmCIOcqVysIFSYKTdaTmkX35+nw7jqrFHubG4ZjYSW4s
QLM//olw3TlQcU03LmfyT1v7YL3bSi8v3RJSwL9y1mOdcPgWzorO5yruRaLV
lEsykcNju/3FO5WVlH93EOo3fLSFbhlfrhHCYcnDZUquhG6UfMp4lLqEGIaJ
HBeSdu5XwOX2mq3paUzEyLJ4ING8LSP8wcxVQ9rYFIPpeXiPJqMijSzsj7hG
mh2UU7UK9jpXMfkTmfTa2KqKTGqjVwxfjGlFicsUrnBmlWiO4eRCQ5TuQnCT
D8SvvI3TptOjCfuJRYyuDizBn95x9k6xMgGo/XbzisMMy9OV9cJrMKzwY5rl
eNlbfqKljOYUt26C6sEpHZC7InUyyZNSZ9AB4HIDdTkh1UjAhyO7ABj56WEI
klCNspnvhPwgczVIgCNeCJO4yN/+yflqTvZSTM3j05+2kEdoJOewS2HFHIlh
uDHsTjVH1j00JiG2kJfYwbYeS+PtSQGcm4PPLLBzTHvvHfzxLTn3KRJFH6wY
vyoEkzW/iV4myKp5LzSfYlcl46O6NIgu/8xI6TnQoW8vnRfqa10RFCC7g9kX
K0CaQkokmHa9QPhChJskUH9rQL4/HpFqsQFTPihgC/71CwZQ9X4N+dAQfP6K
skCn0GO5ACnq+09uSkCBpLb7owcKarUPeSjwQywzhsNSHrH+zuwb4hNhkD4Z
Psg6pwaBIq8u/duQRzMQpf7Liwu0+9VWgV0WO8uzzaoMLAfq5bDlJqKmUg32
Vyfb2Q3pb+aJ5P7rGY7qh8WrnNv7P0DkMjRvRTgz5kxYdgks3RcG36d6poo6
wsqQgWwhcWWtl1dC8CzSh/XO80m1jE6LRihILNhbKIIJ9XGLYDV4KMeMNqvl
ZK6Ee6JPtMaT70/w2muAdHPm53+RhhZoWlRlNR+YWYRW112xroriZvBg+/rT
WyBjLxC8EKyKiZae/7sq5yM28yfeHtdbP781R4ftcc/J7fftGG0nP1uCV55y
eoUpRuvmyxuJe17u1whjDHWYAzsOzun9o+Zv1jy+7XNrfgbEqTWGAH9Zf/Uh
QHQzfrnkvCJxwq6qFCu0yDa29koJ40Vml8hUTR0XSmyCe/YbtBUee9QTQjtI
oY+fSPha01tygQFaKbVwG0sNrPi/PnXmt+NXi/mduv/1TWhpYrfvTvx0AgqR
/liF7BuiOju8h/1u9m2zcP7x3/6sYSQNIBcHneLg0Ehui0N9qh/09Uqslsnt
Ff02susGNwuyn/BBoPLgGTIVPveig0Xz9oO5TPwBOAFZzsjzx5yVtD1PECyF
DHuSYflrXO9bID+5W0AMVqhstIgIkct09qLqnRYxobhjxNRx33RTy+6zNHnu
NnPWP/RcxVxQAoG3ANyMpGLZKkwXGbF1sKFh+gNL03JtmiW97L78VmRWvwYd
Zc9r/eo3GPXXFDCvjbNMXra4gCkzBDvLWAo6ZlhcvNvUnooS0M1t9K3T1s5d
c7KpO8rJgcdPmcVnVs0b6FKPA2FzBsLNj61PKVQTsKt4/mUIwEQhtAvJAlM5
dASm0lGTSigW9Fbvpv6h4ED4AYzYyLvL5j6+7rBDSq0y/aCP6cgNuXRo2Jc9
8udOIcAEwGRj++u/UWjtGTEGKxkURH25DYflV8fAg5so6/8Pv6qJ1cONMqo8
b1QkuWqd9So1IQsSAwEYjDuhLX4mcdpR50+rYzWYiA5fg/3aC3scyJEnw3zs
Kl6s1vwb++cmcdSIIbLMJqfI4VX1Tpvv2qK8D1yYuSwjuPQXotPYnvc06V4T
+4daOZ/bBhUYzBkKZ3Oh4RtCHQ8kWU2guihv75s5yZfKSDhJFgDFuhKiT4bP
/dHyMYoe7TlnYmA/6pRs/7VFdO6OKlSkQ50bWy2/wQHnPFntAVyO0pCwbGrI
8C9ltypl8UeT6+rhPfy/nvM/4lh8CLrlrkxk4qOIoEbkaIYDve/z6HaCWeUn
k7mnjq39RfQ3g7Hx2stfUb4np/aUCg0M7I4QMaAUMAlwfW/RDCSnyECupxJr
GcaOZ5harApscSyABRmV5CIuFiFX0DkBAmvtXoy6Y1p/p3dYX4vdvaf2BGhC
qJVM6U5BADyiq3hKt2Lcfahl5gbAxZslyDrJadoHMHevYPIhkCqKwia9xMiR
5bDX26WOgI8G6YPZWceSQHrhcvl+n3ohhCgGRUQqx8hYhw+O8dp7s4rqUYLD
ujS77OHkDPbO651GxEGt+2W0YCmKjljdREuUmcKYTZQMmLKSL+IhWrNGVHXC
Ch0/FHXKS0IBtUV8Fsxx0znIP6Rwnbwqa3cVkzV5uo9CNbBu+NeHm2dhFucZ
BD6ZNgtbxqnstvAVMxFp67gfaJWuJpL9q/yAS7ExBNcjsHoSeCRaWc7i8p2V
iL2UsflF9SSLCSg0Bja65Rqb+T5ysYlyQ8j9yZ8byoIpr/TE+o9EzjC9rXPV
+owHg+umsxD3gISwuZSC5FLkpB+3XIFvnfNsgqu41uoEr/BBAaDiLVKLbMca
dOemGEypcuzhLPqkUZ9tCUqnutKXEt+ERfqmwOEx3QUEHn0lXPyb7/8B9xU8
0sziWBdrEvfrAFrg+GIP9x1+slkmKIDJ4+BOzQEfgEhL3W97iphT1rPAJ1H2
IVJ0wlJjGcr2A3uvQu3/w7IQvX0+lFqOEkxKn/MpAjFbT8/AGqsKstDDfWjT
3BzZ2yKus5dQhyko0uh+op8flOLPJ6foA5MmvUjHpar9h6hRmX4x5O4wO+JZ
q147sGYshRsI3wxFoq/0Ow80CpeKQVfGUY7zw9qJzvmqAKqpRBX0NDR9slYS
Q5sSEbl7RuKpNFKGIM+2MamS0eYIDGXdKg5NjbhHMlJ963vWL7wOjoKreGbQ
wM493t8N/b37io7zHttWKrQ8kfno5ZTPe91lrgdu+iHUICyQeo78gUuAamX+
2nS9jOtvMZfhlznaDFAWxzq1+7YncbL1xLkEkxxuOw9sg4XosKCyx4p0tUJO
5Rx85ZK+bOZAobl6oyMdZcKZaktPpf54qg5s+Mxp7Pf/+XiLOyUYpB/GmPAj
Q2blc3ePLUHXzY8EAAjpBng289RXpDFIBpELyQvk/qEUfTU93s5mCz9rIQuZ
t663O1U42NOtkEc6pOxvlDGnhl7Jju+U368c7kDvCsxdI8x845zlcn3JUo3i
stuifY53NKSt/aMsRhc7FraFRUVU05o5p7MAPLw+U8w2d5mL32io1G/QeK+u
CRZP6uAlS5WP5zoGwAD/nWCfDcEs19oFloq5D9gEdPdvDHE1LC49q8v7BvDq
vbEWGuBsV3rFrJYsqBub/p2i0Uzumx410jBy181dv0qGNyP74yeuG2FubbxL
o7+M/3greVL+endern+rgNJbVGAFKHWz67ZdwheKFug9Llh/NT2mppT/aeeC
UDj2JF4bCYrVz0X0LuzfPrvkqmLzObYdDa419DP0pHU/sp6rSpNbGirj3XQi
7wdYymt1jNhct/o4fTzbL2ApTqzUR/N/HlUyQPkC1RDYjhvXy95HIrzuIyjB
X+/pVVz6UXeuSKrtruykvdi0iautaqIYgR+XZ7B/mWtU9mvDGGXfDA2pkvYc
kHgVReC8/uVvJpo1bvLacnuOg26YptJnMVa2MoMZhz110t+c5hq0Hk7PpL+1
FjY4LWOpsaQ/uZ+DqodmKxP34Jya0l+myGQDzRjKt35wrJoOXFbO5YSaLtli
tiT/6aGbnhQtdw7PoRDNg3nSUjbZ8xvdNLyNK2toZn1aqnJ/9JymYza3bUFL
lXdEfoqMQph1MKRkFxYVdUVGAAYJM25pPZfqpsM//WT9LP6vNY1GUEI3LsXO
gUp9IEAeXJU7waDkVsmF4XUyRtYtm3quMzj9GlHWC43eJiaIyLPq46Y+Qv83
tekdkt7KiVQJO4l0lr/aJpyftfVXiZuI6S+CwjTDM166PzaZpHl0Wpv2mEcl
CWu8z+n2c4TWdlhOgK2VmLSdMgtzEEV4B1NuDbULlzVdEu5xZgEvo7uor2+1
++ac0+E/GHe7avRTFIcVlSOOJFmYrw62w0FrHjvfTnSNULSLeRZ9c943xS5Y
ahyZ3xtY+1juORmZvM/L/KbCMD6/qpDs9nuyPEtm4eRzYhzDRAgLgxuqzRvR
yks/JibPV203G/nP5/w6gffU1hFnDqYl/+aMQMEa3WhI+wUkw4xexH/GiN32
Yj4CIY8+9IEc+iCA2HzT9fvq1LRzL01f/fAB9VGlcf/S8Zrx4EQv44sAui8Z
M1sdDmP1u9WqxbynSDILShGgGrACzwZwvcNaR0oaPUC8oTaqoukfUKm9asQr
DhqJUdHkkuQ27vBqxyjfCprppQaqHC6MVtEN+QjijBaY2l6UUjRH46y/dfhS
n/x951XjUEeGLWywI+pjTYsjt9OKCrnUNsrHrQNYjuv8RAD4xepxkmB3w2wz
PKiv+C70QHT4wkd80ol7ZEen7QdjJsdsYPNsgyvQ7X8OW32nGs38nVTZuDSa
7NTiSSTmM0/kHFvkaOL2KPiRXiacoE7zYUcXQqgTrsFyMz0yHK112ALHq+03
LTV3EXwOnYDv/yi+zyUzXtOZeebj+BkcPLAuILF37AEIr/LCHRxy5B/h0aA2
JZBRT2z3+5Tr2tg3dpoLrgzJuE7LVhE9d6zB7f/sQak1g0quWKUJ3lYZUvsF
U1bAcNnwk3EYefeilGGIPMK5stYLtsc+sjbdXFHiAgekxXLLK2spjkhU9s5+
98S5SMcQ4QiTyjnVZspbErQnxQ000oxnmBefOKug3bc1VGvSAPLQdf1ZNgKq
BV2hOrZmP1aa/SwY8gpbPWbjjlyg9HvcbJlTiLwL3t0RWrN2Gsas5uH0SL3y
SnKoAIOU8X6d+JEjbtypQC4UMPQJOFrlbTK93PHOzXqFX2YvVNIMnx6sdDuM
iCCst5JbXa7nslu9dl5IxeqsyDHtzotp0oXrXe9Dn2Z5yskCSqtKv43BYKDW
72MNhGZ2hqUqZ8eR5z8Oo4t9uxDsp8yd7dCWBo7qd/rJhYVGVWT5j2U1bdRy
zzcjbkcc1jHpjEM/LH/z68NllxPEh3ynO9tGOSqYxALNzMnuAbj5QpCiSOft
4Q4HTk03ZAsweLI/fVL9gsQLlZwHeR3LfvrYBb7RsfRgyfJJKsCttJrdGsfZ
iINmG8HdpSNdeCD1Xord1uTso2rZezUWFwUasnQNEGCi61ylUJ2pONqNLTyZ
6IycKUJZA2J6GgMlglKaTyTQHXJj0t0yj0WRnJjOnpkqlFeKjA1Ew916/8aH
pOfHK2e/76rOh2NRMPlma2heYpGteCDFYETjeAErvYPH52+EAB4iknyjz7pB
7lYEdoO44hg7BI9j/vuxS/H1jPm0fGQlXKOMfJ+GPU3u+ESmyJZa5gysHrg0
0r7oUkghSFCUMzCfKdohn/w7/sqwZDeZqRFcHtYFFyff53Gus7GYMenUcUCv
PkKii8dwwZGjz/BJmtvSjcLg4QdDJPy50NmFR8X+Q4wVIwyp5guqttmNBfhc
zMx8YmMc0FdCDvId7S43Bv67pHX3ZkIOZKHWgxANOp2iYLQzRcORWCtt+vdA
e8Afh2mxgrJ2RQX4zS1hlhpQPjzekpcYbsn4Y5HlNodHlxK4XpG67k6eCbxe
I2CtSFhEQlhBrzv6ovoPXFSfYOz9Se0bbLgbn7AS/LYdmg7hW7Qe1Qp4LM9s
fGDpXjnbnb2l7/ApTu20MGES0Fdky/rRn5mX5K/5sjJJpGfKLFBvxQ3Ly6Sg
oj9jXu5xVHxMycWhaiW6ffLH0mvsU+vcyqwcOyO3kgrRSUxOxcD5itnEFRzw
/mcmrgUA5dB6XIDRTRnYupAQUjlUWMIAeJosd3r3MeW/PatNqONmDTqMvy6n
iEKtIgUhH2s/ekL3tfWrOQVEtGyvJnHm6EnKj9JUcGC3mGRKi68Pe54fjPxe
CKeG/0noGCqH/FVlSCB0bAKmtwRyxyIGRiGswK08Uhi9PjApvplYUsjSCuBm
SdjHraPmD76Pjy+oSEpjGsgNFeDT0zf6wNs330/qUgNTfRCSMbrEvCGTvwWk
q+NjQ2ymtPT51mawgRB6TqZBE1W/J5XAwUThzYYO9R/Nn5nhwsxRLesf3It0
tPe5nuZn+KIkUeZnsIRNnqLXGXtop1fRPEaV3n0HjVeMyZG/u9aG/AhicNBy
LkWcfoUyU2uri86scxClJQyT4UoYrDfPOeFy7u7tgvnI6QQ37T4CzCDdxvKo
pJIHM9AMe2/l60w/9+IvLFLcjMkgPkhAPpxXR5NhqlrehhhIAx3Wer4qSLdT
WfJ3XEy8CrW6vbwaIDjoyP98cfNpLnmP8Ph5MV1pLnTK/sTskUCRPhC4et21
cyC/usYwwxb3HOraFljC2PhgsZ6g0VhnhxDoFyWVAgZgFcKXjc5lvZ0hw/eS
alJchLU7NIwR6AZ85xweeXxGEDPqG68g8WNcuCN5oulBG9bYyIiyAYICrt1Y
MSGW5Z+OL8PPEeID2hdUAMXAp/zTuaXtLmJ82iIzJOfdsTAQiYs9ykDjbtba
R/UGsdoP0jI02qp6f3ZZwgrgH864ly5dE2s7MNdQ0xpxIUTPyAjd//9AjRz2
NLqh+rO3kKPvAmJ3XQoF4EDf1Kx2V08bFy4JckzGZ1SStP7dmFdxKqwAH0Ct
lLZ+Ehwqs1AY6T9GGJ2ycTfS8/tT5jmdjdmugI1uhmVNHVd0YLQrhx9GrStQ
rv6UkGO+ZD/o1LFELg9ENrNfSTaI4DpHaGcjSX54sdDZrOOONaSVu/Wf46Fu
HGdSwYj4tqWPBnZokEK9kO1eWdc7HnrG5X91BRalVaR9HBClhNkk6xxovRmH
61hKPNmh+XUxy1glDW6FA/+uW+iZNBG+5RtP60ECNZ3Y+ch7JSOwr0sK8H19
CAIOMA/2aj/WGfg5YQC1b0e5BGGGO3GWoHmPZS6g4znFoO07iQE36anIJhrS
r2DV9Jv8eLZz8caDHPa6Oq8eDiM3t4mDUy96JkfKa0UBTzFsdJ4mpKydeKOs
THy1XrrRdT7hUSYceGER7hAE8CemgS8OOGDlOtpcTu1iWsD5mYgsEVGbHXbh
x4PvCq+Rqr7S1eE+tDxY3roykU7pAOLZt4ndrkcaMlfSAx+V8CSBP59ucQGa
AOoZuFfikOERYfQHFs+IsjfNyL/fTOpZKuFJooAqBfV+JHITHMw/dv0PMn+r
ojtyitQHwBsj4LWb1+47jrFIVSf40EE7yJ0Iuueo1MbzB+xcjKpd1uSOpEIu
+Zp35UCVzEotw1ZGvld1d/1PoRsSDJgWrVKgQW6ocvjA4mWZkYPIaNvkr7jk
uy+9/XjYrzrBoTys/UE4O7lxqyzL9jrz99tX1iCcQJP/O6AWVmEWCrFFr1nr
qt7R4IqZP8E+AvmLwmfINfr7Riaf9jaEuoyd3vNWdvSQ1DVWJhquJteUyEr7
2V6kmlwWSJhWT3R3rQZ7uo411fdSQ7c5MW+cJLt6GHoCs+m3doRiNALYHu7s
5mVruJi2xjg1hBM+4qkKWrXA+HCFhnrF/79WkhHqWNcbQeMRfZeBRws4NjrP
ArdZTGhbxtmID4ahb8TwMowVDf2ak+t8obpURZORZN9GV6aJ/eoIHQad1LdE
jLRHEPqUoJIqpJx+dURMVS6KsF2sYr1hxwlAaIUF/vblWCoM/33qN6pdrzDI
eNuv/NNVNJpS0MPtP7bDSdp+xRrzhPhVfzJGtTrvf6DOxnLri2eBGmECAGH6
qFJrHyg2u2fe01bvFPvU2+l5SeQu3dslV5bGBFPT+hsUyCbCBi9twb9xefYg
AKbmmN9p0q22l3cEhUrONN2wEvkPUtfy4pRaePY/FAR/9jZDiYIHBEU9sFd5
41wiw/rlMXx7BLu5wBwvtHFjfwg+QDB0drch0WBgYWn+5DfIwo5CuZG5y/ya
aC7fuAmxDDzu4Ov7POECar34oJB8CSUzByBrNe08uWq5PF34z34FwQmOO1o6
h9Aat3PT0o5i1dEZQEQSoL9HHDZr5E40u3AcmjJGLaBx48CjhwKpblHCO5xC
fOjlpQ4jozEwSB5vmjRlA26YFHuKH+88SS+J2N1jV/X2NV2o1RpE8mPRv6tr
hflaHriGtMe5/loda9K3WOw+eJh04G3Cizc9TqG7uZonRRdXGZkd42tJehX9
bfEz3erwjSyzElZPKDvoSOdNS7nTdlDbcouVA3iNiXzlqs2oQJorzIXi2ukd
K8lZQr2C84tWF6rZMb14GJSlCbXLuJ1mFu4gR7iF+4H3y68FxX09Z4lKLDTS
qa6OXMuOvUHFk44LrYhiheqh/d9WDVoTg0F7Xh6+W4dAv+kjTMKgebt6y6Bo
lNOjs3/CwxGtlFImZwt7+6NOypMGtNXXVlJL3jMtUn2SSirY1RsLv298CKO9
NP4hJv5PfJZBryje+6tFr3DdU1bYZL/XagVakAOcDbfIM45YmO7cSDuMdxo9
GDbYIPCuHWBxLPkQxN11g4yCm9Wf5nHigiC0Lsuvn/LJHXjnP70uMSsTlF1U
iXcv/Po69JIgDiG2Sy3lspIdC3uaw48ObHsC/LcGvZpFNmvw1NRyVldXG+nT
DWxEl9N8UTjI1yetZU9nObRYG/CUw3evmwKsv3XoQCyyy6wZuoaNe3uUbJQz
X4591K64GY0D7ALpiFL9fru8E8KH3yV35Ku5WoJ7fkurKSVb08wp2EjJA4yZ
WIF6dhJGk8RC1v45koiibkJd4jzt/NvZ3Sb9zJ+a5aAqIuLgAHqE4CdK/JqC
ssfEKhDMWQgdFSCDiy/cxpLyaq7F3ilqFr/N0KXa0cTno1B95TZFPPZNNpfV
BqtGgJvrYYWm2tP+Oamzube8PWj3ajalT6xFJPItvW01MWQOYZCltFYqQlfS
ss8u0lKQIIPVnoNbXh+9DCK/p112X7SHloKYYBOVd1WzbMPSK4acAWZHFpd3
bboGvsoXU1Cpqc4VqaourNs0nG812dE9DXxO//xxUplDaaVpBIPXAcbilOk2
175J+Hh23F0wX3rbFCT9H2nBG1VBuUndfUI4OHoJqKuRhn2l5jPzNC30b+6k
1cP0wUg7DlDp+MsndhY7bIrqppc+fqoaYYpDvZGSag8OK4qVxdSKwLWISPgj
458WM2ZgwFdT4m2p9+LjZE4WdwUmxqQQOXqm27aETXMNJVtTmRz6jJJqHwNS
BpJSqp+ykRZAZu7pmEH9xrJLkIoJdQhxGLdSHWj9mvptUokKIuRK2lz0aPAL
sdWdApPPOB7UxN2YcumA0mUS4uHqA6sOyeIgLIOVubYXkLWYcMOqxXaiKdCz
acXEgKbJuoNcRn+pci7LaP/dt7Lef4rBzBrfYKgGz14mMffmNbMtrQvTuo+R
Me08A2Dw4arHRJ52F1kUZNBK0ZSmEnQ4OeJmYWbFCVr7Se5ay6XaHsMzsuLV
bMTTCoswk1sXBlRhZBrCoc7OsHq9YuMw73pYRnFlYkKGnIllcf+WeJFhYrSa
wA8hSy+D7XNslNHSEOs+S5s9yjiOXkgxurBHs7wanrFVpRZNJQnQylrE6k0a
x/33SUOPViVH+Y6ZQzkQq2WH7LpziZGjm7Fy/ZfjMeUVsNRfcYC39aD+HfA/
EWoPfcjmm9xpyakUmgAmJPHjCp1jJYx+o3HYzIP1B1jdHhBxpYvPpsDeDDiL
upNrzb7sLxhQTEyQJ2DuJzHteqNVLd2KP9NzvZlGExsLzXIr/3LtFHjNI/QM
3O00JLzEYi8+MCLWcz4oMgtnjslL1H1yoapbWdxZKxbXCEG49jDEMXld1s8p
yxfd5adMjy/MQRSwHs/jqvTxKKPPodKo+5Kb735Gz3TE96r/5cEN5d1PnUT2
IoT4UUc9Jxr+ZoPXt1U0kWXk/kBIppn+UDEFGz81gu5jN4wFlkIs2zilNQ7A
djGYWCvdWBTv0FyQYD45b6I9Z374rN3T1yCjzbdI0xU8OkJmVGBjAMbhj6a2
nvG8lPZB/HQfP9nYwlMseopflUvNBq4L2hcBPBfTVgHz5Q+l2yYTHGIyw4iV
hnQmOUEHqUH0hwgMEk4P3kWMK/EGf109H9J5HOXINeefXnhQf3W7NfvyNXzy
G0UG4BNze/D7Wjiv8K06fv4XuFmgAhT4qqvIKvD93yz2mKYt2a1gfPYSgpch
+dMm8QfQaWG9TGNKsKP47zAh5xuwImI0IOQK4vLmD65NGcvAQ9wfBsFp73p3
So17KxjAiY+ZVV5eIe58CGubaNLF6733LLAvdiqFZQgGgc/FCcryRTh6dfzc
loUS0HQbRj7khZMHYPV3663TaqL0Wodj4Yd1C9vV6G9bHb+2aAZedEaZE/Tp
v4ZiamkqVtLGBZaaBIENxOU4ayzuS0jJQEGPRh+mdD1LUvZmF3ctpJBbVxXE
2FQx5ShWcfBwj+z7MqXGPmKfhWJ0EtclZZkfgEJWb+aMOO6kGL9qgPaxGVks
h+KUkK/GOvRAW6GX/7pA3mfD/VO1HfG314mmOt8WQCAY004Wx4WdDtQ6G7Hv
93NdVGtf5ibsFoeTCsq42PZhEkZeHlo/fwFDd6Qz7nUqzFktI090lVbACSi5
taLPyDMTDpH+3Av5BvoulkHrTx3KPGDCHvZQX/cL/wbMPWe1iTTxMcXrTqXa
FiYaXUWZRv80Tn3e+sJM0zDGz3lwNaHJrXk5XmeYo6h8rSMxPyGE1TtNg4ny
0B2KWjEpk3hPlo/C+69MP1wxY7qiDxqMDw7iGwzt4nHBdV+cifOv5DuiTP2J
jiLuBk288uJfAc2TPcALEO2MC/hhWItzaOkVSjc3dUfWYVvz00+QvaPVvz6R
M3x5K6Bkj+PLWh5pLNGYUj2Jl071hAA/QrxYRs8vXgeCzliAChJBihoLFtUj
9l7WjdmiY0daUfDYfV2lTCiDv7d/QxXHiyTUMvYzPsRGKuW/eZwzuToz2zjr
aowXyK3QVKoIEcbH8eRJciQ4QhP7EWSlYChLNavVUV1EmR7dlLS70nFcj2UR
38wBSbnFyQ5d28saNb5kr216o7PI87ZSBNQgNf05Wkkkc4Eupwtj1GAs0kVd
y3oegdKe0CjlJ0Vp8Jc9wKNarhscMTceRhVI6vR0ejizG9HjiGK0QP0zuDQm
lzgfZ7Ye3JG872GIGIwftqqOuT+b0uRfXJzZBH3SoK8cHnUZ1YQeqa/pyJvL
grqKvry78Zl7vAD7qB3nW3zp1xCA6Q+tsugtMRljNZhmAxgE1dIpIf+bFef/
h3JGFzdePRkRteEaoNzyr19+cIMge2/kue9bLvv99pd+sGZapam2B8gBw5UW
mcDjDvjevHVHH3V3zd9S/PDxqvmcze5dMggyB0/pLZDnlhrax08QkbPRZ/f0
HTFNhehr0YFPkd2mlh+quuLw1i8sl10Cj6L5Co4pVG8dLs0jFQItU/UQWWIM
kzpfmGyjfzfiKERecvqer5sdblsPUuCsd3jgvt5vdKakeixKIBdG6P/2WEAp
9dHgbQ64h8Qbyb9XUOIXDb+H17aZAJpBmcLVxDqjBVlw96jC+X5JtMFAg8z/
ko8q58COjvU3Anf4o7cVYYZswDRA50mgc0GSKuWFJWtQA7DyOd5gpa9Skw2f
9e1D4gQWdLvxvuBEjAPmC2fs7ZcViNClfVopd+WeXaXMCgStas1CkqBfVIRL
OAU4A0jy8DxGjmcxOHQVE3VUI4cmtheqzFB6Bmc60lNPqDFzDilmQ/0f7k7K
nCDxvEvxUDuh2G8SW+VRE8Ng92vBqhugRiQj2NUrlYKF4PHgHpL0QO/0r4Ef
lv7QjsZtGtUpEwHLIwBn0UvUpzF3dqEUMfkSqmKWnO/hADokif51Ftw7tA+e
eEIv4QhKDXOYlyX60rJ2MpQobeyI+32YNAJSoZ49GqpOrTuHauGljL3kQm8a
dJCXfvwzHVbJHUPxQ8/oSlV8r4hT7j7n41IDtFadKmPitFiZG7wZ9cITmTmB
nCHIPkQHe2S/fjVdTOxi7rkXyp2iFU4wAifWg1uNhM3trMSHHF4lzClg2des
RK/mS05DdkfK2nqIm4aNCADd/LMje3lw6ne4e0jouyx+yI5rdHsT6KCflEqP
3PLuxczOK7cOPr7l95G76hHWpYbVFXjugqwdNtdK/e2qVuaJcUGs+oQXfLXR
vSsZ8bxSX8iNDzEXGakBTCR/IXZo6NXxyoHtazWbwMVs3fM8Ni74A1jssIgA
L5AGDTeQAoEcxThJ17lq9JV5tWK0yyW/d2CUB3uAdSNV5dSBWbUwgVmHNfSn
8YOA7ItBizBkapft3SCL0XvKoxlFvCz4oyHDLvbW8mCgu+qM/6zBXDTS8OOo
zgsbbEXsweVKlz7aJokxfmIOqLfEe35qrKFJ8sgd/fXnFPkHeWCLBDYcCdYy
gvLNASTWKeuncXXXICd55cz0gC+rot1FeK1FOtPyhON51/xOiacz1GMpOJJs
9UPsBDvTK55EjxkM/ioOEQGfOuiN/jfUQOnGGePVzfgt1cL5JKb8XyBjDN2o
E723vctLykHAMv2OD6edhjZVs0kwYLdjoshKewfr2w0rASOYZsUD8aukOY6f
IJwakSUfIzmLWlqJLhJjm8RKATS3YlKsszCCtBO1nJp/KXGE0iTsS7in5Y3G
MWfwu8aEp8bcFRfIxSOvJvzjh4c8MAWhb35rw2FDfN/oEL7I5dN8CfbrOSft
J4BY3G/wXaePslXjFxC+5oEqlI/YJC5cVhbpmG2Hq84GvTXySG22iqmFs9Bn
rFnJxf8CGTUOcYYdg96c6n5IYngW5yNqWVdawZmWAjk6Xa3Rc+MGotRrzOKH
yDqrMAWWm8jx1aEyQUAFsnUVaQi7KLeRVAbFeLpzlBRjfUHx033txVsQUZwh
pALe3txXnwuZNFINOnTUmlA5PzKcaz/yY5ayLPFV0rY7taN05IKCOVD+X6X4
wBnalwGrhTPGcY+aJdrqL74Q6ZW5x1ayBZNHARamoqGwznl0z2bmEKGCfZHZ
jb8mbVhPOqb6E4KUmPGfRMMkcPyBhkwjCfke9hPMotWEfC1S4K6GeaNUJfNS
HI0T4WJfr1YhgHA2TRX8MxhWq2i8q724C9Ic0t9BAYDYMOKeAfSNIb5lq35o
gBIvR2JnJZSN1zMNPCDNj6H4ENGfOaMy1aaWDzcDn5MNHZRM6B0s6hPxiND1
PR5aFHi4ru1v2iwD/rvfn42/JM75qxV6I5+5WmjFkVBUXXrVs2p9er0wsAuW
4bB/FD7O+Rt8efGksQdtlXEyUoyD6rlgtLsw9qIWq7pk4zjUJs68dAIDD6eB
8G92neafQ2nVTzuI6yP4jIFzpcmNyq+9UEEmBNQoO2X+WVnj9tCPk5wHFuZ0
ml+XQH8tBG/wc9Jg6Mr+FkteKYLJQ9NxQ5myNDHHmw+A46zuF7yDHlN8I8zp
CyXTkjpAArM2fm/2xhv6hXX9wdiJuAm6rhYWLv3ZJ30Xtafalt5H9DxX8fgM
raDk4+ffirTIyoVDrzXiyf4cm0JD6L+1MPPDQLJ8hA9TFw3kat8g0yGoApGR
URsbx0UUKGy7Cvk3VYVRICl4htKH3BgyvTnST+63DUxQECXK8G9pap/uxuw2
138FqreOqtzJrD/A4tmWqumDWiTQ1iwxYHmdUB63oR6x9o3iJPQQsXmxq5RW
ZCin5CD8Acaxb2O/5H0B23CojdGMt8H5T6oxBfOddSLcYi+V5wrYHP09F+FD
Ch7m07miXZ3Sq9XpnjYA8219j+bYD5if0l0+cIigTY+kov2zWsZPuy66swx5
ALdg6hvLpsVWGRk30gmXaxdKukhquNHhLfzuq6Ke8iUz1vWKN6/0b/GGmk4B
fERnJwg4uqvoW2abQSeSE77EIFU74zMkmMS6thgZdZwjL2G2bDm3GPVeAlcx
+EqVJQCIsKRkTO4vz66pSdaVE/xNB0Ozvhj5wFl+nXAFxK3cwNMXXpapJ3a+
dY03gjS8gZmTtSouS9e+xy+1zZzYkKdqT5gkJAVc8R3N/geFrZ8Qz/yVhgm0
/Abaai1+dauz6UqeEhlVM7cyYur35hwiQYVk7Lj0dbnVfhNoVJ+e+H3FLhZ3
lIs/UFkr6ut4efCf7Ol4U5/PpSBAwnO8YzX8cNRJGNhMh/fsE5yKnhIUpUBk
5QEc9AECYN+t2ShG+5ie/zhIr9M71uF4NeQ0FEPQjP0Zi27lzYwbjsojC60X
ToK5xw1Fh/+s963Fiv9Jab1hkgKIa21mDdP8N7UbLQmaYHnmroFEB4kwqia/
twRpu/Fp6HcmwFfK8XDzvZ+TYnJYOv0t2SWGHc3cbBlncycMZE4/pATkATBH
izQ2D58vickSu3cjG5sUbr3sopkxz6g3xtVCPSc+bZYzTbW5LEGBv64cKRk2
MipO4kANNc6OAbXokjvDNbB2FWLCVkxiMujnL19ggKwR9/5aO7SFYdl6KmPW
e8sN5yUAPlayptATf1vyXuXwyltUwCWkC0KUeWoZViI8RwoFsRX6xc3m7Tei
DidUFEdPSYu0VY3CyRgvhpJg43fNLDWx6ogK0kF2OjOTIdBVzorbqIGaU8Y5
LN+MEaIi7D8LGmre9eU9PDFFc3sk56pYIJ51SajOxRmN6dKraCt0g/rNRtQX
puzGfP4m1t2+18oLH3fT0u1ItoKa+BjHOULTMHtdtzGEmgZOT/AYv8niG9/L
I+9F6t9T9/8az2j3I5qMipLPs0yA0VpesNF3ROg2VaH3ubxxalLtIKb2dYaL
ahlMFoxRt9iY5F6mDzdb5CqPPqrKp1qCc3uyQmAobcJoRAkpsxDXUhaLkobM
CnBaIYD1s2d4C4Va8+h3modyPky7oatRyu1rxOKrzGcH2ZOXMCGpz1ZkppxT
1bksCmAlhf/fVI0YPrs204Fr1NjLPTlM8vVCzhTqyoZbdrhZrsQRvpM6XZQj
EflRrI/40kt/EJKqk0Od5j14I1D2YEe7mRkE0JYrS1UCtx5quEixkhIWUouW
pBbMKlqe/6hJnD5MivitzUj16Z88KsnNG7fdOK1irty3RuwUzggbFzzT1P0A
J4vAhPG6G8uoHU2DC6vxnatA0aJmc38BORJ3sCN9d3t+BBP1xlpl9Fd2yATX
7vhOIno10jHWESejfk74COONE4FBQPedRNSz5qGk14UXSvUQx5NOYcDGGA9p
ezliC663hOCECi1fVCkr/tbfLLLnEd8fXBnF+HUc9PqEx4v+DEfU/wd33Hfc
S86aXcUUcXhsTDdFU1E4/H+GcoJP6UZ5uJW0mC1oyK+Gfj0QZjqdr7xlAVTv
/R2U+e+2iRgnVp4Xda+nsd2TcK+i5Nr5a0pBnxDF+uK+FgBqurn3rMmo/G7H
vlE500CfupZFqwhXfvCi00XVI5NML+MSHf4152vSPpor20+9Y495WgIh+qKa
ygZN44YFmnRdAjzQ3gK9JhskkH1qVOL8PTSCmsiceOKaDFvX+4WLK5wkKdFW
5/FZrYnS0ZF6gx40xHaH5kHKL5J8Lm/1M14mKogox4c0NnRPPV0Ync7DqY5a
RoD4Qx3uXLpehmcjzeN2qOkGXI3AjaN7V0HAYWQuUms10e/c3h56OUOQFtnh
YEU074cMK/Ll1V6oW8cc+mIVUVXXb8ZRmLHVkx5BVLa6XzLDtYt9ERnoxnGb
PpOOGI7vRCM4Gsn+W01LzvD0LjTJkTwVFv6E1OVx9+lcrbRwI1Wlvc9VI/jW
ZzWfO++tlQRagKXtMxX/Dz5NFkICecne/1+HPpctLi7VVjBX2LxT3/VUNocR
02vEXjLtd0LOapKgFVq0wJFKF4ZcLAfom6YWIChaHFayBjTtuXN5nHE7dKMS
48ITcWqw/hK2xR0pMMpyQe6s9sQrqAzE2eIJQnctSCMb2nMJku8qU+v94rsM
V9Y48V/0VmJGMKQFTwNFy1EIbyLsqpuC5dn4qLVjsr6pyu86BSBrVO9bfd4C
Di1aoCy0V9L6eAynQxxAoZ0BcHwwMkJhPtNa1cp1MguwQHGM7Hgmr5UC1zdm
/LNPHYdRxzibtzS+ythca1N/1OFfRC4PG3G9Qcm/NXATB3XJQWl1VZ1yJIgc
01kiHIpBbDk8mpDNUYM0XUhksyxfev52vrzPmumsVrOAaf+mDyqAZnu8Aj5s
HhBkgz9vgDY+xinNbjQX/WfRT8ZsvZpNGe1OJOrgc4KjGK0tjxoajXDaJL3H
7wn0i1MRQoSF/R0dgKH8rjApWnwcQ4tqUlIMlAFVyKTxyPK7DCcwRcy3XobT
iQfig383tlxD3ah1IguskOsth326WKraYomCNhojdz9u55CU690LhNE8cGNe
Jn8+eTnuHMV21HGqi/uUudOqnN4JZFPiy9frA9BfD/A9//yi3Pkw6gCWvtmj
8G9efifeWVOfuLHjCN3MjaVMwf+/N/Ixem8S3jn2da2WuI546V4e/ON/Rxmi
1KVhKc33V8AbSBvlX2TpPQ7P1p9B7DZjvSCvVFTl7KtooBXJB7zxhQNAfqwr
k/mTLCGNFn1VeQTuM3KQjHdwIvBDFVAZ9TwWSsGsIoX/XDpjEmjRsmdpA2dA
XMBfEQDBOdrD/bbGQJ89xB6wF9uFJekZBCk0KK+AmPwdKcjZvzjUcjeWpMwU
i8xJwGLB+jcariIf+J6OHb3vmtVmq45MD4ZONgabYe8XVFuW/UPkteF+mDAX
fX0YAcZmoWqM53AySj0plYS5RakDgVBaFZYFJrCi59YVW9Mmdbf0N/ottKPA
d0mwgHxAKL2C3N/BinIQAMbyEiE/dnQpcWn4LAXujqFg7JEFxasclHKe8g91
9dRTf2tQev75mXp2Q/Zkii+Uu68j7O3jLqhvuOi9MzjGYGaDoxeJch1o2aw7
lrxsDXn5Emz/99uesvcn4u1t3CBl9KT6Lsi6Hm5ySZik7LqxMB8v923tLyza
YvNq/vzri4ck5pOK7yx2c86Uv9D5he9H7U1BUfZsjGzne/sO+/maKSlFe8/6
78z4HQNakLWAXwFx+QSLEXq49UUTE9Moh0TWsrrNYSURziVVrDqPGVnm5MAg
Wv2M8SWk4vc8/B+4JAPfxYgZRZNppvGnoSo9h785oMdYHgp1zmqeyZVrWcQf
S7GoVkpJV2uihC5xbuXYqGFgjV/07y8zLhu3w15gUBT5WPHOHCiEU7jdD+vm
KyXiEAdXGOPOf+hWULNKlzY76SooYsWbAskMlXgFx8AGCGqYDR4Ap919T2vl
DqkOHguJ1HzRKdBkkFpmQr/TkKhlM2s41GPyupZBsLubTHNr5GpiTTJIAlgv
Ua3a5FGp3DMhIUnwyoQIxjLAbkLnNngFiMtGQ1BQ8+sCGD4jgMerQmZ9E6VV
jzleRXYhd5EoWfbeUUg6+pvLEgeCet7VnfIutpuROXqrdA9EIE//4SiRtMiy
aaT1fwTU6at6trQvrH61UiUoDqcrMGNW7ZumEaGDicwdpSNOZYOuBbtscMVb
BHPcJB4i/C/s6WbDBe9GlN0VdiZGlKeHptOfeU4sXD8lzc3lvbed4kiOLwGo
9ZVNF81R18QOMsaCcP1m2atG3Ml3OPQcXFfayuurlr6c880CPhRyzxaOxDAd
HzScmTnJGtKr3hyQnUOuTH8fABpGJ17fAxmy4miUyQRtldH7iFB3UQaHeVYs
qCfBsb66VAenPxN6ugLgKRxB4QRJk1YpADGU8hH+/oAHqGPd/Lu0kyyWzq2+
ItCrLNXEDO2CZ5kJnz/XYyKoSPmf1N6vXtFXycPRPOU7/VzOG4PR5by2qf8L
+udcxM0H8NOpDUvwlxTnm9r71BvxZHhXNnusISJTDftrl4KNdLnUoVoH51oY
Cr5mIuoJHv7r4/rfYkPvQVlR849W44dBLXqMdmK8DsfPjtTCg7oxMqLNf04B
W2l3xFaELG62i/Mwar35ReM832vZtkto700teqClZ7OND4XwxK2dTHFD3uFZ
YaTeDuYhr9UgLaxB9sXPjIEpoZDMKnPb3Ex6/kK7nSU7cRfrVlvVU7NFJwV0
FXGVN1Rt2vyrf0tyCvYSl6s/cSvK73qJBjDfFX6z6Gs4rmcVnG6Icrc/htAw
5tqWXBbHPorQNn5/IrKagVhfekl44PbU5u27d68z89pNOgqkb1+79j+iFcjR
/dEj87gZhhZ/c39MoVheDpsI3Drd4SSzV39BJLePKYbg7asIcs1F5j4A2970
x7oPbpQoiuHHrP/7bwB7bYEggsfOhiVSNzRucL4CwnX7jGmnhi52b6/UhjVD
4UzMl83mPl0bVARuBOVc0MTq+YnpRrYuTzJuugeWh9qsYPKXhwajKqqfYaab
9rvI2IklvrrQEjVDDmUGwvdTOi+lYlCuYi/XlXbn0oiae9gRLaHiBpVYKW4U
Ou8EpWF2nT17NVsCvybbTe148mp7jS7wFK8zWv16t18+LAmNAixe+xInv4Ej
RXNpIdmQsDEYAqg2zbZUcb2TcicDemVDvcwpSrF4+tpqIHB3kefhj3o7MNjg
fWgeJ0FCjM+ipidu3FMCKm81TPgb6ppqdusRdgj6FnZV3hS9ttr+RjzNKkJm
sHu9YGYwoHevhSdFb1vWf+8umxub5IznohN4uSxmyU0mqPlZjgW2xJX3OYYW
jOMQ0CT7kpwzvRdpZ1f4/669GTTkrHxYdZvqBjPr81v/ZHy400Nv+XayMNP2
LXoy6W1JQFXcj2I1Jonvokh2HQUkD14anEVNGUAW7lz+wqED5yX+Qv9o6UI/
e7gNdxjkYj94Tzmpcl53OYmfSc684kuBmi0Lj/ZS5smAzR0+jxjVuJFNcWHH
IVcJ+DanY0zLoXp/07eZrPYrqR7SE942o9mNAp6dJNEPC7OxAUlBZeMjFBuF
Fa+ewdhSSaoSTPcDxe8eI/vF6Twp74OLiqHao03fl5Y9G7uThRdhmI+oh7wX
F3yPilqSYrs7vov4nG0F/whgpIZBeMapTLtRNOi+VZ4K+LL6QGPuE0RGQPA/
nokhutqzV76pqPIIDxsWvY9jWd8RS2oqVHBtn0uRAC5JuYz+VcMwT1qnolqo
0SGjveG7xf9sK46lceL8er04j500M/K5bjODwhtumkgKcy7ZDKWZscigjvdQ
8bS86aPnUCckZpaWbNqEEet+iuCVf3N1c9z0uJqpGFruOXfmm7tngmFenc6H
qc7n/rjEwPLGIam7oMr5reSrUueI5eX/etwOKKF/7JzGr/etLyVdcq10ckwk
VLcCiA50c5vWzxPSptLxq96YNz9MMi5RAvbjTj0X7QxnyVXzdV5tS9QMR9qV
hx8Bw9hKHsl9SQ3RyES25C2iDl9OasrtFIHq/bvEq6der2neyQRlht/+XrN1
6Tu/Z2Ft4qdzUF99kpWhQLAvrxCEIfENqAIaS1C9kGJp+/zs4Uu6OA0Ii4RG
BOdMT2uFzQ0ntXpur3xhFV3uHn9WRADjdBKPvYlJXFzi/oEU18o1BIibFwSS
43/1Oxe7QoLc0qBJCV5Sdg/6Aif/TqnwD2oHDng/F1oYKtGPzaeP791AkRXz
7+w/Pkzrp5ffvimEyX8auwpi0DvDQzZrSxrYOXiwTIBJgm3BKHl16WaERgep
4uLsdV7tQCzvUJ+bJ8Y+JUxGMJ6q8Px5/pPBTX9SPZj5iz1XPCIGJMXGXHT+
M8/Yv4w9QLES8+fJ6qegsJq7JqjWKTM2BugP+GVjA8mBL/cwQ9ueG7FjWn4L
i+7W5eyXjGI799MX9QOS4D4TGwOpaTi5qlbnc8JBR9fEwgy78uWY5t61kDFZ
QM9r8Lx+mdj+cee5p08g5bKuBUXO/xaCrfXMrAYVlDSrBC9fvxwx5ICjQF8T
dAvGt8+n5ySewJM85TWIbYhQDJHLF0Fsto5gVlz3kNdDDqGvkWir1VfRCyFb
oPY/ojjbHsm919KeyYJEE5fsBAe1CxIo1xC/ow9tkMBzTCVCM1OvFnk91ZZw
Nu6y362dmw1lLRGhBBoSrE+3CT4V5yms99eT3O5w0ebHNw34pkTCIZ28qPOJ
rNWXZE6/AlHT3L1f6HUvm+eMptyuvUSBae1Qt7bBMlOVbm+LJ/HxAXFCWbqo
ZeKnRlCSTiWDH0ulrkC+kyosBWdItmcap0VP0posKz+Yguid9XCcXK7Y718g
Voomin3tWeSHvnESKMiQXBVuFYKI4QaDo3Y3xPNg115XKDwTwNW/u3EZ0wTI
9EptehAnENKQdlPadgkwED4eGOs0u4lCiQ+PyazOJuoSahPVtK9rgZhTRAha
zzKXPeaiae49z4003dHPezrNiquKgwn1a858cmrRAtobQWah0+eRuMg3Mtgg
u+FaQmBPz2O2hEnfrXYSL3VYgfytoESeQ/6TT+SnAOaCMVW49bnKhpLHp8Ud
vcotJ9bbJEcoPACOakNXYwFKi0qzjSgfXe05wBC3wnPePVl7LSIZqAYMvZL4
7TdOtq3Mc0MQyzIo3B/G8tAyt9uFWR81UU1QIQXuNXAAvwfd21LP9dojySRp
560684a4SNKXzszvGTwBLyWh4KW6AH7RPUw6y55sCD3/r1KHeE+C32MiZ8Dz
Yl9Ow8d1rvTteIFmC4qQc55reBz74EWAl8bFuGzal2k07A8ZzwEAl6MMm+B+
/KKU0Ahzk6bScUVT01Lhxm0yY82NPE8ejIV8mK9eXbbFtuy0RSIPI/NyG2lQ
v6giFDdmjB3G2UHfBwgwPtZcPAdTMfGzeyX6RXX/J+Q/9NR3XJYDKy8LbOMl
mtWfwp86Xp/sBNvQ2ju7SLuI+5OkteHEni3ZqBYY+eJV5R+W0Dx2131tVd9w
MnAfzSRi4TlhWFPM9XFGWoI6elEG04X/RDmWs6ealdRMkhY+FKLPXDyBXvPm
ZXN3tSMYPamVfTg0xelYiBJbf/6lBHDAXyiMG+/Rvx1MWgeY/h2m8g3iflkc
4TGiPBPIZKK+nX8CdvOGb9aerkBq0nb4iOTUvES9dkyKJy2B+jiqwhnQ3plB
vi+UWfGNODbP4Znj2y+1f27cdIuTo4G3Wt8n9JZSCw68vHy5h6hdAZNi8j1m
S2VT7BVpCDHqLrN9GUAfx5nGb0Wyk171ImHsF1Rtq+oZm6MFzN5WfICLTx+o
8oGFNt4KtLAXe2mLSopz0LzF+BYsWclRAcvl3nWA2bPpeVToD8vZiY4ZY7Iz
vI8dGv6P8RS9OZi18Igun8R2jnL+Q8U8Oq+8vpoN9pdor6L2t3EsOvJ7mvyW
xQDf/W6KKc3zn6STuqnCwCZptkH0U6NzR9asGmxjwFm6mZvtpcAWfdl1sBRg
sWnG2QACmQGS+bo/O8+E278Ans1iHSTgT3ez/HQrY9OdOs/piVxu41jaNzQ8
CWqC3ikDgkRs5PP3c/VxU8pdftLf4+VevB6Ym4FraudXQJAsy68LU2TK6NL6
Y8aov/cL1IcDOcHCwZef4Thc0Nxp0gq1mY9bVVkKrgSXC0L1/aC0sK+U1m/R
g0teTvBhzeeq8XbbekaMR579zRSm3pS8sE+3gJwOXKiAsYniG3RwxXb0miP7
X26rITgkWNJbs+I/QKyTS9pE4zn/j0Cx9eTozLhy8qdDT3oXIYX8a1L34q67
JRyIJmKENqSd7mK/+lUIauJOlTM6ZpuLiANxeMan1RgnTqOvjsxxrK4s3D1T
wzYBCNBlFNMHMY4DB58LLzyJ28VbFsVu9lvdXCdg5jPo25HQ2clRxXYPVuqp
powHrTFl+R+9i3GMvBC5IaxiZrCRYDLcyj2cWlrZ+WMp1uNx7lhHFZaR+QFW
qS09K867qkeJdZ6dOanr9hgrmnkyPSASamVL3n10hUkDgkejpJCcH9aihPQT
ERoiC/1Hdlx8JOv8WvIWhRuPPk30QbXS0o4jhH2S4+Qz1fY/IaLtV8YCiPnr
TG3RToyWXsntfPHOB8h/KON/mEYHFatKc0dRB8KOrWoccMNnM1PAOh52kZ4s
1wtuP8H1Rxy9EGGdOq4m1qhk8sZyZKJCXyEd9AMMi+KEfetrDIpnHBsiWD30
mc+UVAsPw7EKmhaiKsYYLKAS0uuGyZofDcctqT+paD9ExuzRyV5O1exz5OwI
gMk/RW81jDQhYQvY6pScQ5cN088nZ2MEJM4d9iDQVpymHFoPrL5K7Nl/Q7Vz
BbeeSukX7TQ9NXkAylp17TM4cvUVH/+imUDAIVWy8x9irng8Gled8KopZVT/
xaCgsJbqknnEdQ1hUcteYS8HWen44pfYpLE+nKWh24KTOX7CepAPHsVy1AX+
walUlgqhjmcylfXVCOVRtbpw0xN5Z8dwJ8gNTH3lZbZ0sH+b53nOR53gE6pH
ER16kC0ikNzgI63o/mfkfp0l2AdakBlpfbYCg+oAUtqBZxC6Ev0mMfF3Uvea
6QJr4+n3Vt2kdfM4A9tlNzuSFmyTpvrAoi0jS0Ln06rwxJfnHNqVtyae/Yvp
4Tg4EPKVmFr3Zo2R6JDLmLUTeSJXR2bHaLzxkn8bQOVqVOwYcZpw5MJ0KLzz
qUh1DRfBZ0n6AJMhXRV1U+0sXMNzWSUkc8lM9ABvLghPzW5/ayDE06rO9Dpj
U4xNW1ItUqc54L5Gix5kYNPArRFyPvEjOcqNTzJMhDNwaMSiXM+TodoXBUD7
rraU+jXt+D/jKNDIWu2n2Gm4y1p0593LhC8GPoBPWve8ipZbTL92oi5Veqeu
+rSL2yXehspeiGQa+7i+rcRRRaVFGqH6bAiJw7jfEIb/vVXD4Mqxzwu8UcGj
HW8ce/8mGBk/Xo+aShp10zImTFysFAL0RMekWNx5SCSICCOkpRFhtH4RKND/
Oxe90WowlKyOWMeV3l8mpncpTqGlvtuZCA3Fx87F3eUyEvYMoqU1XY8gNBbT
Z5ggoD5g4p1Q8LbP0SeeOlCp+yBEK2IfHoeOTaVl5GojQ5e7797qorcwbYyt
KXWenKnh2OIMuPBN/IVaYmhZSrQXozGY8ePcWB9z5Pyk+avCRJlGB2a3n4P0
dldu9XGnv2asxwhUNWBKyAB7E7u7fnZyNRioTidXnn6/wAvG34Hila37wxK1
Y69Z42T01F4EwesqS0fbqnUIkdECJBTew71jnYGj0Pz/Znzr14ID7pf8Vhn6
lcOe38xl7Xq8Lg/dm+s6aS6JutlTrj6dSU5sjtVJDH2/qAlEob7rxub6tbMH
LPSH0kasVrKByyA07LhQLRS/8ou6ljIv8dQmR03O6eYYv/N6l1giA8D6mRYu
RoPh/V3Ob39dTXLXvxx+lsG1ehgNSnPzGM5SgECzqwM18TebkXbebdWf2v4F
5zwRzDSMKwvABK3S0eaxb9ovOxpR3FYswW5OsVJeK1wnepG3wcM+h0zDVaeq
DVorY8FaJlXHLP3NHCO5OBLq0Fn2CbAnG1BAMbpgodwyJ8S60hHbQoBLAlch
Zj2gw1PX96vnC/Ce/Hdlf4z4XXvAHX6uhgV7iFQxDXiLzVpJjf/OVhBdPhs9
CvOCLBbBlwbfKEIIWvjvDR4gC6U5NI0MRN2h1GNlkb5SgXKrkoVbdOmZGf5Y
KVM2zvH9KTxtH4Us0p6SLREif38yQPxS2ZazTKB0nqPJVW16wo3vvw4qkaBd
XSBG5Mn5tGs9TU0by1AqiqZMWVazI9Wy2DOw6SqldxUChvXNOZ4CboHfXDwI
4Hfl+YaTb7L+Pptk+fikyb+RPPa70fX1bcjLiC0fYL0bFfGNpDhdtntGAySF
UMscMSMJyeffUVRh6sgcpdKLE9b0Ft8Erp8b5BZH/Rodkj8MyO6Bs0EMmjRz
a75C24U1qB25nG41cu2N/1n/Yr6Tt52OhFVMgkuhBvq9mEp128FXK+Z+p7Ge
8rXmhzUp/XnXF64LDm4/lcyhmlI0YMvZ4/YMZERtmXcBfrcyWL+lA2LJhhlu
mZVW87MgI0/EcibEd+bLoKsY2LNhcBvWP+yF0rmGu0h+/+LiGEF/ReJTYfRF
nguqUIOBHo8ezHZyRZ8xvWHooNbDu/COMSaQiPAAS+y4QfYdWQaUtSht12fs
hzjbocIsP93uoIgJ8e6h2ts9eJEPcnrPDgODsWm6VYsadxrxRebG+sn/GpAV
OXwbl/8lIsh4QWAojFXVsgowoQ2TwkRkBRE6uqa6Tagi9eZQ9X1kA5TQVr3/
tbkSLyTOdGWtneJl4cCvHDWS2r+2F34AMTAxUWy//BwgQ+3fBcEeIwh+CiTg
eUEm9ImwhTkXd0ln/iNbFVkRl6LhgXQ5Fm/3EWYGs7weKAz+32hcOVHYTeaB
KhkJgjgT5eHoX2UO8nBhHHaF9UECoI06h/cm0GMezQJGMdfliUpSN7JOvg70
b2iDNSC4Njsn9EHdPVWe493n492usA6k3ASabAjgZdzlnRBzH+nFGiQCvvpz
6JffAbfBKH+hCGbWt8bQ7/+thTalPmSEqPtVWESgzGDvOxMehQF14bAn/kck
zNxheHUFATyxlCgi65MXluGQMuhLSUHMpGyxIDlD3FcynfbktUwYNkSPoBn+
MeMD20zWH6x1vZJ4Sy1HBW3wP0lsZqQDwB+tYP4kQV7mRxNJ0Bwy8Dz7fNcx
b/zx4Sk9EsEGZ2HdADGJzXryyh0komhYxappELClZtSQTDBqcSaixka1UpV8
Ilh4mYknLqqaHY7khfr4daAH1bKcxTqaxo9KxVSl7ZDehnYd1ue/Z/m/DxZV
aR5tyvQvVEjxL0suBlulnxaNYtV1uJNQcB8+tl/4ta9y91A2wvc6iVDceUN8
318xywfuORPYApzHumKbkfOJjcI+7ZZ5BNw2doc3PobrASdwEQLsKTjGDf1K
hwWyaXlwKeZRFiHCKGiRTZ78W0ynTdo2Oocnc4qtL/2z8bnwYVUR+KcIRwSz
N+arMJXzq79mrNWT411JHOfOiKgyxTeI+3DL6WOnijpBErRlUePWgsDxL8Zo
Zr71beWlXE3elGc+smPOTwBnBc5HK8UytCsIyEU0LKLXIhOc8IzII2RS1Vs/
EphEr/2mtABt3dggJg0ZgpKi/Qn63X+rGzeW2RMASPH0yKt+pvJiIFRSouvx
95a2SGRykB+fLVcOqiUKzkIiEmf2GwvvkgpIszS1XOywe8iG8I/gSiHFx1la
abqaQduhZLWbGSGh/eUpDrJN++J8MhrWZjLU6JYUPbhCLTbrq0NzitCA5bLt
x4Iq1aM0ND2o1psISAhTak6cNaBvqFX+p+N9HrhjtSXTXI21U41mp28bnLfG
kXT5U1fct+Lw35xIyWFSszKCxRUV0VweJFAuuc34KhKkaoTarlteqAPsnyZT
xOq7tzAVYicZoQo5HwM5fmFYRFa1hlvvtrSDBLJHft3Hw3cyWgEM125Ude30
TQraeE8s1Uf2ckgYuIwc9zJJO9GuBf6W0KF13KXOCZyIcuZ9iSXyGySj3JRI
VUWsIzkh8w1vJ8CGRh1YyD4GzXXovG9CmOKX7BstK3M1axLAYjxny9r4r39d
Y0c1qo3ao0tk5RidD1kP/c4LHjUOL6tNjvfKFfB1LcUnNmq0GHKIlJPmEyzi
97RgnPWditJIIxvSFZDX3axx9a56c/dwUJ7bKWZu8kY3LYO65BSf1uC4mP8z
3YKOeLNvz/Ur9mboEG7c04aeMkGGawCV091g9SI4L++Fzj59WLDCDxqIGpXb
YsQ9dacPLOQSFgKvIrSOaKoLRgETEZtEuj3G7W+TJI2iW/XL+jFHmJ3e1L4N
OQnOTNL35/GdMeLrkloJwF8rXOGRUDXJrkfDDKSuoW6dKaUm1V+YPD3Qj4MU
r75WYG/nWE6mfIYHQDY+iuRcOh82TD4qv7R1OmBvzS+sjVoKP8vFjMk6VmEh
Ww7Uh9z9dNKSuClzCZZaPmOFxjxyIwT3sb225U6211gn0gEj81AyRHJTZNLd
6p4vOTg3gfz8mk5gWSX8yx792sgRmKQTt/9HNtNzR4r/59v3r1/eTRRwSawF
l7Q9XcO4XAznFUoHW6wkPIG92xWBvC6+/zCJGKY5D3GiKSkKO3w+2B6OKz+r
wmaaWjPW06+60+yux37NvGMDSbcYlDsINsqYTVry1mL+KirDepVB4iEZnpfG
6t5bX3z3tSrHQJiG8UZgBT6sb3PES3jTo5lLY91DKF158plmUHXKDvJ4Br6U
G8M+2YpkRrQhnnTwdiCb5s1UQWbHWzTuCh6WlTE14HtvDBNbi+qjLhJZKYri
75IIfsZZSCuu+ECm/vYeL9j+9gxAxBkm8vog85MgZx1KHJ/Ne302HFPCUfpX
No0a0t7t9Df/EZATflDGLT25Wt9Qu/QhWeg/lXM75apZoP09K6TMJDrLV6Vq
SjdOPqCsv3a7YKlNZYSfq+CnBtI6qGPdmpaf4bpUsgeRB8gPeXZ48rERfaPv
dHel29MSnQkRglq3aKQUZH38UPFMk0tnzHglyxKOZc05878/K5UGUsvV7Wj7
ej5njmeOTsuYDXYu9Ay72DvsCGxb5yS252AlJ5xmSY3JvIMVpH3hW8NHq3bS
oMorrTmQQl+CwY8a82uBbRnMi6/FFH+HhLFR2VqpgV/MUrl0s0U0Ab82nNzN
xHQMg4cRySWh1c4tVvlfB+Oe9zEoVePx+hcc+uOe8p4cgRl+60VkljHDQ/RU
n0O7psYN2CKt9uWbR8SI72vALkJwvhWHRQRjhJFkD0C6dp/E279Gqqy6WC4x
JZumRMZTNQ8IPmTcZ/MIAo+GF6bR24SUtCWueiEgKLmzPgrCbYmJzZgr460i
78M1Ucw0isFWlFtQ3iFW6spdOISXtqUTuniEjfZsOMMjNrmiYZ7plP9BtqRd
3n0oyngKNElaDhCV4rW+u6K0RsWAyZZWSrdld3gmiagwCndE+IdrCRfRD23D
52lox3agLB8VR/fG3V+NFusd4yBL87dBS+SAjJ92WXfdSFuhhV11jiZDBgBx
pBlx8Vi/9tTwtnuPVW+voo3UaEm+td/gKBlIY3um9OnrwtsgLy8LLNwl2aCN
LPwy7cXLRbAAJsIB8ZDndGBmLr2c6xoVjpSC7QDPgJbIm9Yfh7bswQJfFB7N
k3FQNjHImThkIKj0T/WIb+ymARixgzAcJC9R94QlwUKgSpRmrbRsO2Gm5S6J
Jk88tX9NMOco2s4C7sWyx56JVzE/eMDWU3VJpTsOtV6ZjJDSf5AIq30lXLg9
nGllPHWlBTy2K394Cii5JuaZVcz0iiFGa0rC/v5UNtsWkAg0ownqK94Q+dDK
L9YIZpCuwOpMtWMihmTtQR8eg3dN1r0i+p921SgNsEualuRwbi8kOvrInLlO
5T8OhVEvDHgPWJ1MdtTiz+vHRPUeG2zS8jk2zH4KrBRuURgguQltJGFO/lNr
I1nEgaBKKB/4wd3PF3Y+aDiIWZOMvyuXXjj+Pm/LLPj2tEVYP5/M4MjXl5kr
71CAn9UQ/lrVGAkUAYWerq+kQGXy7+pxn2BLtHfX83QFXg5RYMo9vDYZWSt3
L3Aq8n8wavLmoEupVimoXyFbzaHqbN3pJmSwyHAZKkwIwcWOMacu5T5d0w4a
4bgtsTGLtoT/u6qrlCTqkSj+IajawcLo/kqUx+UJAweKdHz1SZPJMqQK2dV1
ngoLhTv90vDShUbsM1Vlul7iVml666bX+neVTG9mC/8eSaTWaNj91IJ2w5Y2
dEjuQQFHP45DKt1buX5Lj7MP1FUwsWZQd6hOacVT3N1/LliGhvpX/aKLCro2
E6cmCaRw0U+swLCV7tTZrGmVVPAZ1jiVvhkMohA6+no3llk8ODNRb4vceSzO
5JSWI9EZ5DJRTD1yZoVTYvG2GWAfj/LJt/BHc5I7V9yUdOpsL26B9vzDG8Io
cyu0lr+K6eKT/2Xh5nbYIJNqUetY2AgKJ2N623W+B23xrAeMCsROretSsWBl
bdeqP+jyFB3KQehvQ8XLJCHl8eg3iTalGa00SDizjtnjluPyIeq/eenaE5du
g6lWb/YamytshfQa84D7tflikF5PgVxOhICZRq/9Pw2nMlVXRTjTL3/NZDyv
QoN15XHGwVh5KIU3HuLs/JzVaDxLX43U3AqYAqEANj0zldVw9tly1bfaX6r7
Zq2BZNoCUWBg5haXlHahdx8zhmHTYvVyfri+XXl5Y/wA6N17y08EQkhWHCeY
zocu8/U02ISXkh5oL69TViyLwWEhdZzrle/ehMrf8Z4ehIsmQksf/RffRk62
ml+cGWaNFiWvhxEN0cVT+1AI6C9cRa74FvH6izI/lN+UlAyYa0sL/ZiGmk4b
R0UNPXPDsx/vhT18p1+4ToaC7xSxglMkcvc3lbdO4bFwcTNKSHEKzwlj0D8U
4b+IKHv/g+6RbdAK3ccVV2gZygQB+qWpbVX2VVMCuTM8O7HtHAwnKvQNu2dT
zkjidYGUp+BBeZ8a11bpCC1P5Hepf6NxlfAa1hzXGbTicHgfV9PHedD25wIq
WihIob1hPumbHTe0NG1xfw4mw6Kmi6e0t7lEO5pSZzEi1CMo6retF1LKZAWc
dXpvquzizjLiF2SBTeh/49MrBITVVlJl6+Di0e9lroNjjZ4NVWqb5dCnhgEN
XSH8Q+pCVZ4XtCP+hkKdj5FPfsG30ZPNTsiDjOmTlXjj5v0j/XYJHzoU1kHw
vdHN15SjhqdwR4zld00SCh0Ms8RUOe7MaQYHRW+71iaoQj4N/MYpZ17xGk8g
ufA1eyv/mRNXHN30uC56RhcGELvXP43jOynfLKxShmRnj9Eyjd9fE4aR7j6r
gD4RCiuz8FNkAF0FGLoPX6jyrJbXmAB+d2C5kr3DTkopSacnRNlSMNh3NvcL
cPxSCM4hOKyVCbqu80DWvqAioSbyV8jJMDXgCZF5qKSLTJH7mcsxyke7nmC1
KQ/5P7BdatMXto62/uFMhxdG6HVMadP7fzU425VrGMhJ24AZuBzfsqIuUVyr
gngJIXVCI/bzF/6PuC26RKmE4QQI0ai6uydwgwIXPfrkgAadZa8xkm6XRVHv
7m5Mm8BpLiOV9j4oSlPSXjaoDKOVoEmTqhZLL9r7JzwYespy6/ShdUcp0DIN
RihNipXyXhEdfp95SZJ3OpAvUv6whXLgUTMQdqNPljiPdDporypXIwbTyBxP
6Ho9TLrNtHa4127ckABzSrohpzeJTixffFJ3h7MtWuGhsl0vEBI/m8Og2voL
TLoCrJ8SNzugCFkfAmMGDNLCXgNIYqIB8SCX4vu7fOiFw2qIHK7k2B1GLVz7
aQZ8aCj/qD40yv7jyCjT/ykS03WC5AiSCsk+v6QOJiMyQfWi7Yruzdq6GGxe
BsnQVX1e+ym3ViMsnBn3QUiB3RUNwqfIaHVMtH+p40CiG2CyASmVLoS25QW0
o+hSH07FTi3NBw9IMVis2D5p79np5eoMw+6iOXRglbzi2+HXsc6f1HEC5ukU
SUjjuowt/v8wnXXA2Bh9Mtx5FWIPg9EEtvZRQ5R23Hj8mielbaknUdHNzbA6
vrYyqw0xSTOt19j6yMMBR5MaijIIcDLhp6sCYYvSVfjto5Nx78SqyWsjn/xy
KV7+qWljbMrzWTDk28OPxGVpUpmkY+FdsUXEPRqdhYVcTg44bHg6fKjNKJVN
z9vQQ2Q4yyHQUldkn20TL6K8a6R7WUuvYn3gkq4Ix/OWZhXobMXC4EMjO8PI
ik9RpmO2XZePBxOSWjgFya9Et64j+ZH0w23naKZhLi9W96thqlr0S+mR0SO4
t+AwvY/lyl37bMm5cuEsu1NM/kDNhFzZHoHdAudMCJfzOLVbuwm93dneUWQx
az753r8wtQv0Ug54HT83QFeRy0siYKhXB9zpKww9yZnL/QTaETm/kjw1E4GO
e4NBniAEC8LTJ8uUqOE1qC0YbCqpx/RcGrwNunvT8JB+wbEw+z7tI5orEct9
PhEEPGnOO+DZvY7ZsiKW2GzxQqbCV+TSKj6Gai0noNXz45cG44H5iDI2NJQ3
hOwDBYhBeSYN0VLscMJNdQudCIZZJBxmo+4lHgqKkSUPIBAAgjKHXwGrht64
pQDtlxQr+K/lDk2qYdt2YDE4FBCldXs8SSDWvQLIVg4jioAoydK8PyrCZciI
n8DYZXfM2omyZ3cn1eL9AXAaGIA8ZhM6MejnL7LktU0q3O6N0GeNNoJ0D1SL
3j4vug7VSH53oGISfX3RwgkwsMvSEuYCYXIk1EcKeUBdAL+cTv6bY3C2lsvG
pqpTVkdcMpyYdrk1HX30xEFjXi4k/wT2nSmAxrVaLWEa2rRxO6bTc4ruLQWL
kvXaUr5doR+NedMfX5Gi2aIMDUdiS2Q3PB3qUIm6Fk3OAlVQJX6Q0CGAsc3U
Ch/ZbHa7tV2IOubG/m3xqAIM/WVxN99/LJUIXhKdceovvi61IrrEk1el85v6
UyavJulnJjPc1yzwWn+5WqNqnwueExkJoc6HOUDCoOrzpxSAbSTdn7SH5Dpt
JdX0nQysJoFcf6B2thsYV6z2NqnlsDa0BIuOwy9kwEVHLOhEQIu+dVASV2Zg
dyyzT39pYOHdTjlJmKK5WQDfSnYCvO5cMqMLYF9dxkgvtZlkJ7H7QzZWVNyv
CY9eeNbxW1LaxZ53jvjnfj9NdHiHS/EHhRgg0Bx4D8K7O1ObZkuMivdUEcU2
/AErDC7CH6hf/aSjON+y6Apkc/n6sdcs6ievzDqgi0Pwi8fX3xKi9HFeeVQQ
rJNHhdvV1NnrtNaVzzAvcQREeuNH9aMTyJswRKc2fbUZbx6dMNvleoofcc31
eoTAJ9EiFBLrDRQCDUzC/ZlYfpssJzDk19L9aeppBDS0/B48Y8FlmQjbXOhd
pJHYjt7dahsO/JEIfhC5dwJ05beI5ypnvSKFVpcTIQvBB4JKgNb8NqCqYubT
tyleIJuCHrRU5aTFCwB1dA5385xPh+/WVRsp/p7Od+OdAKOwkbFLUtRyNGWn
HTWneQZva4HFqYfzbhDtG/Mm/fUtGg4o/He85k3BYT+L91xhkcX//bIftVOM
G6Vo3ZUWnFq6X9xH7BQlWk7yo2VHCsnlBVxpA5OpkeLR7zOTm18f2cfLzNiY
leGRarzmux0GjvHNl+a3a7yiX3CDlAPQVpiOxRl/ALILm+OEGPuTgvAKomuq
BPj5POv3/yjPrlpeiUuXu13oc2EMzjF/nh/VzGflh3OdahLv+b9odjSfN4GN
itwrmlrsI1KAhndi6tmf7iFrozaq9f2RDrpVuO+SdLZ3m+cl2Gg875uYjX37
Q7BbLboqTDLjTkNR9kmBS/vy/IN/lH9793bDogwx5SCeGZqeuP6HUuZI05RS
K0/oCSwa2WPe6SxkA5+llLXh5Ea2doDW8TwtpW1yCppzsokMolmLBPYKo9Pt
HEiHwqz26QGqlz2SXYxl/W3hRyK6JCnwWueEs7G7Pg7IUZaABDMvUuvSnElu
DzuNa2/Th7YyrkPw4RYoUmVkvlnzzKkdqqZF7ad+t80qnt3iNzlyfdSD25V3
Qkj3tNEMR7yYi4lepvY+7KVkNbZoqS1Vn6GxvmdwB3YEHh7lbkI/s2rqh2Sj
BjEmnx8Y/x6WmWCsGut3s4V6o/u5UV38AQayAti+zF0dJE3SfcgKEK9FYr3o
ZkATL8HkHlnWqBqenrsOrCGBastJvCGqCZ+dhYEAyIlMHrSTFxG75uHL72Ln
xlJdtx/bj68DUza5nOuacxDbdfnHIy9eDGAEiEWm6P7tqWlXM1pU/vSnofGc
9dInv5Pv9TTudockDRGxY6LGuA1nV5XJ6MDbj02ixfirr4J+9N4N5pv2X/b7
hYKBIhm01hyc0DFtMeOdS8dQCOD1Rgq/UnYnS+A6ePwHj6s8XAg1n2LKXRsG
hxjIYb/FOP40TCqQF2rkyxsf38arZsyr3wu76GT+MnqEUOH1HJAl2Vk6QA+q
4vsDJAPggmw/8VxWVXW6b0HIvdDNsTeFJ98VA9iA4tuKul3Hqp7qKJDhKk/c
JqNu1r6Waigy+EzhLuxegP5qi/IXtalxhlSRtK/JnUo1rf9c/rNCXkYZlzgH
JkSPUchd48iiyr2mDIeE3vrT7v4C2h6h3b/Jw+RP7JaUm2VrhC2zY31LTFtd
v41DYoCIX7oqk0/NwDXC+Sww1TRzy8bsCw6QXorGcUFfi2KAkuZ+p7HpOXT+
AP+UkOovo3wfh8g3O/I210vyUXvXZqbo7TzOwbRlTb+2KRDlt01IPqAnlDlx
oFH/yIFF0k3JVl6A5OtmtSzlmkmc0mrC+XvXkwWsuwgdPvpyRrjOy+Tjn3tm
b3iXwaN9BqhwB/AylsZ0xCYs3q3bEytSyty4Zs8qF3PX6PD1C7wSG3yRozJk
r3xqrEL9u1i8J/6yGutfhEmX2ipummGGeVoje4lY2SDeaXoBnkfScMOSkOfO
V1qkx4l7Vq7wttdtpjN4+h3JezadEtYkPlf1q2ZEuGwxYPbl9/TR880mGBw+
9/f9PCa7/5o4GZxreC+REVpXQh3f5zaQR8FYSMLuI3HUP3YSZe3/kFcJfjmG
LY10cMI0bfM1dwvHDF10lW6enAREwyLvLdEKzf3cjV7WE3klx2ueCh4/T0na
xcSbcy89PuZiYm3/xHARLL7Pg47idWcFDoeoPZ2e6o4a5lmdXYS2bx5K7nR1
XTykcjPnuv+dY+inJXS/FBgQo8r7LR77rNP+jaG0Ywjs4+H7Kb+vbLEwaRuf
ypFs5d7IZRuxyVBjYmKD4BLFdjKpPD37wjMD/uIcIOrqi/x8MBwoPlGpzGNE
ua0ENWOIOB9l6l3/ADFE/aAiaxmd7zoYSnWtBj/tMVWCLjfiaC7r3htON7K2
1I/LDxwzZ5rPz8Bk0XYCP8EunRSjr0MunGJaS7Dt68GXeDfx0pI0G6oVH9QI
GVvoxM4LwG+b6C5WF/YbvJ+TUFOlx3j1yV8cNvFaisSz4pZZnrIlGeqc6gG1
jmzPmpOISTI4FN+3mCRhdJXJjc5CJtM7Ww3+zNQ4JZeAKjy2CXFEAlYV3d7l
V60OWmVn+hFQQTiNLNtuSSu4TM2Ys1OXbG/OXGalqOPd/MPGm0KkIPPKx29y
qr9F5qEcs33GsS/Rb5k2irxX1isM2KS1CUl2gPJ8JqUMh5LXlWZRBXIaE4JJ
3L5y6Q0k2Z+EnY5zM33OST3gv1THi8WKAeZz99vnhCW8SrhdN4lq7X5oyFTQ
Q5Gn5AMuppEax9KYcPodsHZ4Z6U3iZaRdq1YCzz+QAS6pKtkAs/9MkbGIHY6
vlqOmcrJa3LxhSKG9CeDIij9OjBfyct05oLlutm4RG4LPzaDuv6gu3YUWViV
MxXRDdN5tbiV3kOKYw2OU8/1phIxGdZNk+L9L5oEGpXak4cSK5WWciRivc3z
CqP5Qh27GMvuN316y6ej87oAC0DjxVd3ax6ACb9abmAa7ysMefqjyeeyMqek
SPyVj+N3cek5g0NEyeyIGrSPFjKyaoWbvwMjbHyPekwIlVcYV+WlwCOYGV1a
NJ+FtIsBpTjywyyS9Ai5TUxfHQjcLkFq5TpEDfOmabvwkfgOAm9yZ+CtAZGD
W6BN/djbNSSKOxy70MiO2Y7Ao/jr86ZFclTHbWVAOzWnLmjWob3UN0x1bYnX
qbANLwFUCOQ3MQboxmYooMFMsVtCiqi+ShP1PiMtAl+grXZt7/H2vHg+TsLd
7m08VllSdGQbfPi7WrCWSnJro6TK0zyZv8dk2mJF6cX8xDxJ1Did0jpBI2q6
gfAQWZtC3sVCs8rcRjNlbyDFNGEL17ERwnub+xn2a8bAkMuDc5kafsjcK8eH
lSPI6dmSEIP6vpevAGmd/bAaVodq3Bc90g2QJBibo68QnDEM5Cf6uNBBvwP5
11fwahLLfIChr0F0x0MrvD3f3c95Z4xDo+v+qgxhf7+CltxvA33fw0ivBG4q
XtZF1+GYzeAfx/pXievc1/xpOwossD+JinB9+Iby1FcYenVej5HinTOdVVjH
hZoF27FD+x91Xuk2lAwK4nkjdK9MHjawhlvbM9bGZM0w1Jd4lwOA3/NFs4iz
DNuQ2BoeK7ICo0NTbCC90GqcXPNUQbuFROEGtY+oB4oB/zKYaV3fnl4/sOxV
0yCZN/2Z29xOTXMMIMbKws4rYrKZAd0Xk15I641ZC3OePOc0coJHy970B73u
vNLAC1qwha9QabijsFjzxsawANzI+8drDaEqe1nGn4VUJdXsesIkSm/R8/nR
EzdixaFvWOuvT+0UMBMc4x5s/vWkJQmNkZjseBFTnJR/SIRX3j6QwS2guh8J
UJ6abbEmfr0AIGJUHK/9esRbqLFvy6BkbOVAYlA4vAAvHQ3Bs8Mgr6Kc7zh1
OJ+EQlbwbLRO901C6C6qno3jCe08DuKec903poCH2/MRksLGZqDQiZFC2+pg
8KWlpvbr7z7uAXc+q2Nas00lf2/GBdFMBKznqhGRoqlnDS3qWR3uMorH+PEK
L8E+hKhkfDVEMykhUg123wK9enwG2ZfF84iuwNgbhaPumUz+6C2MR9gngwUv
AB7EdBcOq0uzKjCLY7BdW0FSwwsMYFi1mznH224hVrSBWd1K/s46q491gtfk
a4klXnPwe3bKkgUp0/jPnY3J3TNHtEgPXluX6FWIMPyrDG7JlvzlAOvCtZ6Q
Y8pskr25iUw2euJo9Hm4eOvbIzvrdrliUrOcKIH+svsiTz+0pWAHqvoxy5iN
gBaUhnZ1WQdeHwcaiZDUyxSGmZYow9L3smhcc/vj6Qhcl1brzdPTR/0Cteoi
iHiZglBRo9epVScLWvo+ZMwlrSg5rMtD3439amktUHhjoVFka7qGkNY0jFi5
BBD5Mr7yUo8hFMxu0LrSgruEDjGDcVGm39+9Asav4laSKgCKQEqBOgZjEN+R
YQw1det9qEryzKBkvTbN6E2leN4038ms5rPmv93GBXhMsVwfrzvFW226cN6B
H7E+V2B6ubV7lENu0LwTF63JKt8/EH1wV+uk7boTyA6Tcfc8Y/p8Hm8vfXlw
RLH2Y5i8lp9H9MqZv5lkSCz7iEe5Xs0MhuJBmpYfKlF9EQ9jXuC3caO0WCg4
izm0VO1J3Fe5P2FeqY3kO/sfLViHIa2kMyVrkarJmVeVluzNEpe2QAaLqbhx
49HQakX2Fv0JVmm0mCDKwUR0l0B9M/89oAPwQ5nEqsUGpJ7sJEdycU9cT7b7
/coQdUf6+CLyXCif5cwAP6p9pXMTTOBoSoJU0e6qy0K83lWqjDVe3SUjyLhp
38owpAHTqeVncfbK84k5et8cySpJBg4frCuL8sspnHgglalGb/CcmJU+gW7S
eCd6e8zTmetdquoeGS1wwxNZfqhM4MqAjJpjDCJyTlr3HY3Jj5U7BZeiCCQo
KFuEMQm3a/Vpc/llzDjemeQ6y1suOG9ZRTtBdcp4Lf07Ow98XN8eE9OKSA0R
KpFZZIita/VRGFoCFO05q3DYX8xEuFXwH9olb5YjHLmFj5ojLJNW8KEwc5Hd
uJiuTY4q3dawxH9QizUoyY8yMJOj3+zIQs7jtBEcOQpYgOvglrFUB/RQokDJ
hYzhpQ1XU1AbQqf1mN/Dv37uVnHZRG0TUXZF0fJ2Zr1qcj4Ba3tPStTu9sPp
I2As95+WvAAd/JEdJLX8Mf126g1TVTOm3P+ZM04lHxrssuwUH0WPYo2qpAkH
2HNNk9AtgQ+kSrFDfrtsLbfxyuAU4f8vfhzUaD5/9JYFvuxHnCeExWvaMtaH
pVoXh38gXY5A/C4SxBhAxDMLj8MjL3dOeyH3tgSbGZO0BOAE2JJsPEE202Z/
wA42VxkLNHx1sT9xxhCyWbO85M5FSll+2hpS04svfiscVlWGccskNcf9kqyz
onF0jgWqivLJCMUKJFrI80hxK/67Fp8O82KzfFKapR/jbTr4aP7XjKsjw/4R
L65bJeS1IXtyxQhK1pgwpSqx2Yg7pcwQVx+eBZX5axQ2p42PEcy2bSIwxyms
UKCTLFmjOwvTCOo6G7Fcl1dH+UQt6y2kz5lv0smS0mj2DfkYzrHda6k/IguX
f7NPAXZekidMCqTOi70OCxAPDHcTcZvMTctkp1CBaGq9oN9lWAG5YNaW5FtZ
i2sN+FCJv7oMuN6Nmmui75fvVUWDSI3xVQAa6pWsctz9vLcO9yAhoxx50sqw
ftsWjisqDZtrRtyeSz+F8kb+e2Q84MVgQrU6gSU82e2yNp/rOtRLD+/Iy5NR
l+IXLqtchl2WtQK4Md5229WlR0wJta+rSpFQ6LXjxxoNb3a4t/JQF5vwld/i
yDfeePfsVvlByjNkpnO3QANo/HOoiQ8xzgaaU3L1JidJrJOTEACNRc7mwn5e
+XJIn5AA1Fx6CY0PQQmSiNhY0Xw8iqCApjHeywKXL2di95mY/jDeP4saDLVZ
V+MZnqg9j9QLqbc6S/NUe87WIhRElWdN45O16G5DFY03CQFvOjGnYWVOpmg9
heMmm0s7upffn39FJ4QYl6ORn6146DPnTX0B9XmlMupMdhMXnPXA7RCTgS7D
YJaHKGCAwgrKd9nKdRfTdS5VKcgK7aedR2tWuN0L1UJd47St8fuql3obhRSB
Pfl2QbjNzbtXef5lllgLhTfaDRGmQzS5R14uu61wjcQ9QT/c0fOx8eCJYsBA
xXjVbac0L79EtH3jte4nXnNeSnf1sBrHRNyQ7aRWsWvaYqfqv7IEqSsvGU2/
kKqhOV7VZQ+8174pCV/7amrq/+4HsPac8iqVEz9UZIMwaiW/TfCKdcVY0yaW
Xw65B7Cjgq8/Wd6+TcKfz0J69bYQYry+NOyOyZmgAhLs5YI6Jwd/VZa0dQzA
R6ejKT4GcvBDu5VlffI27NIKkLv7XW2u1D6tMN+W6pJv6a+zgFMdeVkMZJ20
jnymQGJWCm7o2A1uXLr+ApaD3VE8ScH3PCxk1mrCT9QuFqVxTpMwmTIzjr5y
INXYnJPTs0WYFJmgNNGAoaBVMMyKMLsSQxk8ausawwh8V9RUo9QWKq3IsDbf
/0vluwTp4Yx1vmXHN6xLPmaCBoWupGwcd1BmwzExaFABJtJUJo56xOcKmnTv
mUFoDxCoCc/eB8A94hAuCp61NgdV9pLpCBRbRnHkZt/TfxrK+R0urjhUSAAI
PMqrqafGd2OCuAZff3ZyyepHe7zpIrl+Wl//4L0DWdGZYb3DaGT+zYc7+XrO
BCFCqVVnyKVIWDkKqAP4Q+3ZuopcwfzFyA8L8NPaxpusuliN84fvpuE1l6MZ
nrxDry4a4zxyHNUc1+NSe83VifwWE49D0MUaPDUuzuyOqAD435+oWk5SMFgH
QyHJXro1B/u+lveaV1+acHag3cKn3MsPOEUYnbwaRHDrk5hsz/I0s0jFCGR+
8e1QGo31DKvYTR3VK/edUm15M7e50IbSCgbrQZPk4qCtb/Dss7EV5Fy4fGZk
aj3sYjgxNRaxGlqsQZfv0sAt6gUq2z6MrBVOQIlLXz5y2FDiTWrrWP311kxy
3lsN/HgTTjgKt7O6fbNf6sR0CwCH2oOO1ErGwUNah3PHH8UJ0NcwNZe12j3D
wFmY+N636DYa4sVDRHZso8gIyT8aCyHg8Dbt9iaqpTnYrw9irjO1DU5G/3k4
7HM+/9pWahfVtoU4iSWJqEXKo9Vu0z/8d1BfQGpbJ9d8yjRMo+40MHBwd8eP
J0PJxx1Pjrt1knCrvLmx4/lmj5W8T0W9GD4HHB84hWfI9RitCM1fnJF9nO7L
frt2NJdr/Tss34KhTjtQ0jd4exvOJ8JC1O/hTN5VheWbGnIa77H8gi7uTcwR
UdtY+y0jpYrwXJteIVg/f9m17+npqC/lUik9HgIsrrBqB+F3/7VolHgCEcVz
dhnpTXc7bC35JTBXdrXt73ccFINDstIWci/AME9xXTxBddgcZDXXfPBH1w5z
KthIsMfNp5FvZ7NWcmOdyadXeTDfxdz+q9kes/en8GDIUfN4dncYGyqe0nEY
bNxXtbyAt/ksu/yxUJd+JVLS0W2Ilq8Ov2seMHWS9ibOJuxUfyJiO25epJ1m
lDHM6ddoCZdq1xkNK9+sQbbIwWGEX3HUt3VhaLE/MzWdPmStC0RL5oiMHNmm
QyJgLot8w5pQpKDyBoDiT8mb+fCVySuvkmDW0SyCHj+wY4shV7c/rApIs9Ij
3RM8gbNvksR5BLyglVj3/1yWIzP282N1XRU3dSXJu8IF7L/7fLi0LESSTqr3
sOxsPrC/CtpZe0NxGr7H1eg1TESxpE3FZcRAU+YfjpzAyKc9YuyzAIB04pjp
Czbu106bRge9oX3nOzoFcJpiAcyIQJeKbKIP5rlUqXI6gOYNJuamWvUc901d
GS4+Mwe7JebVa6gMBXX0r8WmRKzO0ouyRWGdgjT9Ls0GIHdwSRNmLrTpMqTV
VBMXfEDSmeNp65ZRtFPyJpZ2cBEiLN7niOcVi86MAWBf4gMGV1CKdq+1oBoG
txbh5202SWQZkp4qvoNrEi8XlnDc2Eae8SPRpALF64Vppg41N8+CpV9090b6
SOTwDQkM6h3OIbRpDLEme3Fk5l94+Gzf89+d4gHMcyI+Stk0EuAV0MvnBCdk
CQ55b5HZpDRYGgRwsUURlAaVg09EiFPe88RMY6i57rdyOR3nNLdiS5wT77eV
BB5nLh8pkl0UG5Guk0J4BR2VrnhZ3jpb70Q8gGbazOR2tALZgSa/bYLDJA2l
BkwKKWDDmD/hE3eavSXCFu8/EWG8NadU73dgZgnq0i8Tp6LB/HCQW6PEE2rC
oWkm5b0oB1PTXbEl1sXszOCYjVmoZtDpp6ynWD7DW/FxMOD52GWdGSmpsv/2
s5o5hwHvBpbybEJ6UgZfyO4Npxa0ONYmprlvh5W8iTUpqWbJ8o4Uu29EuhCs
0F52g6yD5Ozsdo1KX6DpOsn9CUZnEPvCveIKD3F5ZlkXrbqOcGlb3GbeYB1s
NQKwjW3nj+lNU1KqGNK2E3Hp6jABeyv07iluJL6ChKvh/t/THGLfiVmkKecJ
uDdErsG4UmzvVjEVh8Kbz92Td/Pc7TmHmaU7iF4MrJ9KkBABplqab1P31VIH
Hm0FlZ1Hb0mfq6PrFC/1Wl4PcO8ciLh/uHIDt5apUozzMHwLhyzP8OL65lmY
cn7R2Cbon2oY+kvRBBnfeGWgsnuDhde0p9XkoRLfh6fj+TADspFUOIP/mJy9
eAM7U08xP7kUNr6YDB4k0fXUbh34XwSrBG0vcer93WIGz+JPQp0DpZDKsMdU
LAaSC5yiTqPwUQYFvJy2+lpSs+JJZjen+mSxXse6YF/PLdiZzQw/5dyKcT3m
EsRW/nSXA0LB0BLS4sU8ifXqIeza0eYaDUMQ4SXv3o7kIlUCb8dWuBQsjG0G
MmGe3KZuM9DK8uMPHOm62/e7Ms0zlRkn+J544nz9N7JrI1AUsXPhEPsij19j
bzhpFKK3pGZdn07QIzZ9zQSIOsyOGmvRjnojT5COhwVM1nMcLqv61clBLyCo
prP+PDTpjBVewMWSBOiPDTxYP2hIPak9IS2gbLU4cZTr4U/zKy87mVAzRplK
IbXJQdX3FLiv/aOhSWL/dSg+V0Q9T6a+kpPQ2AvZ17oaXaOpF64qVFPJP8R4
32XpmY5DfclAPtRl7S2xg4oh1MEEPzHDFMT0mmjm729Cd2C3C/r3cj83/G8g
xby2Q/bRDDbRsbOFnP0qz6YJg0wZvnSXQUXefa6x74WRfmw1SS+F2EDtccAm
bFfUA1bwzP5Pmnq8Ob1sExtgJknvPJYSW23oBy/+Ba0I3v7Qaj0g1RNyj/dU
IvafwvRoXzvBbKO03ofUxWTmaV2QUkzFl+f71r9hVUPepi6AGg9Cn8yFpV52
cXSQ7CfVSuNFa3lZM9Y+kWEKLW3mKwbO2Vr14BUMeBhC8r2r+ApXhgY2wVPA
2nCl53jFN0drUbi1StwcMW114Rspz1rfN53b4rDIOcZ1Ctt9bEtfLcZaY1YD
pToHxpjOFTV7TrcR6LIe0eb3mKwQAlemrtE7TgWhjQ2q96P2PrDZDU2NNFKc
+C0bNhBax86IgJmRgZvCV08Prpt20kDVe1PAju2pbTCM0QggGHG7cHsptfEY
dVy3ISF+7d9TW/cBtImWKeBegGLNuNpmmJ0XuVkcClncHAcz11IdfY1heoER
0MLxYMgP+95B9/DwBtj07s0D2N0iVo61PyMUP2lRFFAR6Sex8ezq7juhi5+O
cUjPChaPn/TJGRCrzAoo/38axTk71gbn8m16NwiTJTYTWaoBafqBcRZnAa4/
5wX9w0pY7tbEiNus8O7N5/Q3WkETjgsiTU4e0/m/sfxszqIY0ybmTsvEIbMX
9ePHlDpkCTXuFeY/dseQArurwvB4Ei6Zup9D9Fi8+/lLlF35gWZPDuKIeQq9
jN4lW8PqptrSvkCizurfVT10zo99w/j0LL0YYu94ZeqQB0W11AsQY3B5R3tE
Ma08cTDYxr64Bi1/hDhfuKHoG38TgAzmtWCfc7c26qHtSHPvrz2ZEJ0lyIJT
xprRRJ9CxyVNw1FsmN27/UJ3YpDwFR/4i0TVmERYHy4PqaT81IYoDS88Tdwl
4ue57P6/heJfPrkfQOh03Vt5PNqRAPJK1+2J7B1sBfAaMdB3vevq/SVRtB0Q
Gqqsah+ngrTuRIjWhib2mlbPnMY+1OgSm87CEa26FaHf0K5ZUhb3joDwXvAU
4mBUO2QCGQS6AdLxm/RBWIaGguY6gOeIc0lbNa70EQmsXP4rd/LUtqfox944
56nHGTtr05/Nd66ZHYsXdesEiPzfqj5eRU3h9dJRmSVJyXVgEEmI7GloJh6Q
S6FTIkDVJ4QuIaLIhyfJOFouZBUK9pUvtWSp3byem7EjsIYwrjF82d9ISTLH
c+NL7PUyShMP2+p51YRfTTdSOsBsVlMTcrKhzqmfjSiTfVzWpEkslgFUd4Gb
qgtac2CWDbGaNJOwam67MHvnVhd+tly0+DYZQ7D39fsN1vDJiohbKQfbf3hL
v2NbjvXQpFBTVuY9WcD/3nJerEsiTGfCK1AsInax+7vWbjmZjjmj1hNPTLlp
/Cdzw0ASUCmO71SQaWQk0a+EYcCNXdXCHeIXhO4w5iXkNOHtlgxL/peqVuOk
THyBJnILzpqsmKj25VH6bcSGONHJy+RD60bVOXnfdl47aCpawcdSSyP7pu08
EbP44PVbFc2NV6PvmAxts3PUQgTX0sMDBQPWToLdm9yB/whnXoXJ1UM+Tsbz
w625Ckq6isdFSKykEZZp0ic/RN+UkQO5yhIKhdwbSMfSVtw2S7tp2kXR9unI
OGgwthlbDm3oKzfBsKIsoriY2Jw/kOYtiFQdpuusnc3mKy7VxMLArJroA/oy
dKmYLn0FWKdzSdl1wwCg3JPMJ9gbPnVJ31OaJPlz8UeOHpQHzJ47o1wxznpr
TVhO9nVE0xfyLdV/LSEDDWyhBFixWnS+ILXyEIwrS+NJdHbN7+od7STdKQ+0
we7pfTzY7UYVX6uc3pb5Kvecx90qCWBdFgK+jAHrnb2lTNCj89vC6JPYGlIn
hwH6mpRL1ZEa6sxAH1mBYYq22HmxWDkYzPh3M1vleVt0HETKIbZDVx2sGhnv
YTKtXBu7LG0Fi/Cy3aLAwRQa1IF91MC7/q0ixUjiMnCt9JFbeNcxdF4wm2OQ
rNczn30UhwJTljygOpfie+N4sxg+rIhoo4cdPDkkFn33E3t2VuawuZdP8HNN
MNp7yAPrt86S6EwDIZraRCKWqVXjhCMPJWKKghx8MhhpyA8hzk2eJmoXw7bi
kKXFTTAJfRCqKdFkoqZDErfxwQNIiE6ZSz5yMC+2FtnNgg8Ae0zQR9ulWxYG
/CK2UI91TevRvzY11QpLYjstqJ5pZ2YvPMP9LamlYXkY6nOJDrDSg13Kzd2D
ku4+rt7nHjtZE3KMhJ5TuvSBGK252YpMQvJ94UstG4o4X45PbNGsoNzKoRRT
vDNxnO/509raRn1iKX6swYJzvHYFnDx4nGxQku2wO6dDhApOe//9i0slAkM+
Q85jBrNeRsuP5/7Y6dN4iW129gkRGs6KvxnY0aQjU+H+EkNugCpwuI/RNxmv
NRSVMECyFHIIO11bYT5UWqtR5LlWUd1fLzwh8KPazn1k/FCLZ/esNtnl3szw
LbDQEUqAWGeg2aiTN4QN6xMrykC6AFiRAyY9HnerrKAwc7qDRvHMbyQIEYML
NJpv62664uqG2BJsjon1Ku0lLwRR4VZtHRr/0p3Q/6jEtqQ/pjm2XCbzB8af
yePBwJW/VVmQsv1sBcGca0BEJ/pXWITeFAZRN4z9ipR5atpsuSG0Pjc+1wk3
Z0df7IP2Lsz4i/WcyxXKkUFNUQTjAeGAgN3p+m2EOhRd8w5kFfOwWjo08sp+
try5ihwAFilEP+moX5wXOuBTzeoQUwJLh7CYnILm6cjxqir0PkbVoIwD97uc
KXI/PJYOduoFx5JEvzMwWyrSK1kAd7waeQdSYbH1Er5P1GMyqcblTxdUFJHn
WtLbxe2Qbk8lLbnpHNSa2oanfTmCS21z1oNQDgMMNk0rmDlHSg/zDJ7zMXS4
v4SK6MPznrhAviHz7SJ326TCFUKyDTqvk6KnEWFq7tBGZvab28JFrm/sjj41
rwwc2CbcpNSnRnyn8LVIOTo0uJhXzasLT82YDilTz0NHdxK9vpI+ow4Kg2GD
pkjGImm5GxhXa/13chDa4IMwZSJdTkg6latFoiKlvc1Y7c56SR1PU2mN1D5/
vNGUPMObE6a38xztaBuzKmc/mz9gMqeoO+Kn5Nr/Ksu/W2FJAM6mFwgghTzP
tHfQCSGgd//CVhj7afGh/yYSuOTY+BiL22ArNk4dctIpEgZOoUWKKj+Ycct2
jUsXqUmS744c1rQ+32ERXm9izsHfHGMl3ALeqZcBasTHeIBxCpyLOwUBb+We
IBiR3hGHexZDCAarEhVNJk7YYg+qbpk7490LDp3D7P0AG4nofPjqZMwqvLZY
sgs90g27wTwt41UKgvnkcTwC+Cmh9L0jhimKmSxQy7F2jl1fvW1LlW1hgTdr
4mZHeYkU0I2iakrbGQ4QmIzyrNNfhty9bsZ0edFPLi/aBWUkRqjpcamvDdfu
nhrL2rVYkBvkKmpXgy4H6QIhFj93r0A9k/5YfxqIFF1GJuCCgwpQooX5t1h0
fJ5/iUlrALrpyKK6+ugbZOim9uhsRIrjdQpaNIHUCozYofL5DIhSFXybf7HE
G9NQdq0I+KYA+hzUg8iOF+fCPlg79vRhegZ7EcT3oKpr+z9Ltb4WPkk6PbFi
TZAw2p7Xa19PHs9mc/ZIqj+xnBqDDY9yGhF07HWBAbe3GTDDd9BUzlvtneaF
jo87k+OsEoCFzYeCc3fI2DTCdmDgtHQP4+dzP39I90D6JFbTS8t5yR4PH04p
JuwKXbjzcd1/pZAK0yITJx4S5zNnA2AYyXglwYDsVPUoRnuPzDIqUgoqvk70
0Fx8LIzKMv35v6DiJSfCSP8dAVb7C7/EJls9DcBD1aRsHvFfYNj3+xtmKxlO
4nFqKa6BOKdPQ4ZUeQKEphALN0lwzhYBo9BLKeQ3C1F88GAAbWzn7gKMvzSa
DrCXDbNSem0z6bqIcUblaHi8U1VELrbENThASLIdvkCkhEqKOepUwqqtlP92
DDETzMFchsZ/zWY53tofp3KQDva2ihXJTnoLuRWHPaSTwzEQrh++Tw24H4WO
TvICcTuci4bj8rEB+xzFH0ywP7V0O50+VzYAdnHIFPJY8+CVaA6Drn7lOgZR
Hp3GURZclJ3gT8HbIa/GW8Hb9sBVU7yrsZz0d45HunLd+/Vm9aqwZQAI5dsP
3Wxgt1F8iI7xm7lw+HOpYwc7F7B58rEJYQceQecitiPW//6c6uKr+LmOWEec
w6dNoEGFDzfE0b8g0ctdUc0Sti3WQw/P3lRiRfzj2BlPVqY+xEitW6ol6YNe
dOmIwj2DsOhZjds22uFMZBnwszSYAkkP/hWjdpN5qGxJO3FIcAAjBtrmxbOL
I+ibydNU1ktqWYzhWNsZyvwShMBiKtShwrjTBsRjmevrzRtMr8I+umyyaPHF
+M2WMq9yBq02DdK58F6dosHw6Dw7gH3A87JIv5bWcEwqWKQqyggZfxuWgIzW
3firiSpkry2DYrr9sSpFnDoI0/GyAOpzbPETKnEj/ETeEA7tQXV0oK46gK++
IobeDYH2Q5XHzg9l1bmWCKVhaLd/fJY4kxHyurlnQ7Aov4CZ9AUPTN7aQIRi
7zz5OuWxZobMqDVtnU4sx0MUdw+7TP7Y2BLRCXR7uFJebyFglNA54+Aaw1jc
4iFTOgGOWZU3eENcoipPIi/NuZ/fOGs6LXjlYXU7zpXfb2YEVoOzMGItjp7E
Ji1YVFpHHqY8e5cpsFWXoMVQV++184kJ8Y03jdJLjpL0sOXxBE9NHQ05hZxE
Kxsru3wPn/F9tMKIKyqPFAJ7Y34B4xAsP3m9Xde4ZZ6Wqha+SYsboGHULPmw
2UjBYxVdrLmEcVBKdwwKahRm+smPwsYwrdFTzQhDxCrw+RGWGfaiKN4St1gT
koKfOQRDv71gi8YMXxBI1Hu/EbSFlIj7GyJZSRAScGWBmEZRsPMVHKXREbDX
1xDj0brEKOo65dQWuotz0T/Gpvjcmt+Oymazp5Rs1rX5fj2RI1qAvoImydo2
YWvzPPM+ddj/1lujtfiLULitd+vDFLDe65cTJW595GQqR1uTDyWeKqkHA3ZK
LjYFKtkALxf3tmVC90ObkwvYZRxMTUAbZ7IOPdrRDEWBibewTPZxazoOJi9U
nxVVwn91OObcEkXIFimKTcq+yXCGpLGsCcK1ZeQ3HI5cPr5faXRTB7q8QSiL
mRJayeO1Xs2tdjXwnAjKoQCxVAo/oN3P6cgBtCj/wvsgF2YIYn/0n5wx3thj
K25LlJ8iCE2n2cwY/J5TWF6DQGBSNInUVEDXQYBmLHDGnCi+a0cWfbu+S2VU
Bd8xSWXFkhsHgP3P7mQgAr/rNwUXgj6CCihGZrt68mIDs64GAH8kKZYtqnj3
SI0VQ/2KJEip+zrZaHplx6HTKD0BE+iZNOcQKiFcAmjrsJtsAWh9BsLfCmn4
Giqf4BA31mptbRrX4yBAB6hM0KfkTYr1Bj4hTka9XTAOoW8dgIbufLo7fGbd
R0/2Ex53gsuY+3b6bc+mZnh53pf7R8hGOkUNk1f/76RXvSUHge+GKzJZdZG0
GZe3kNX9TT2kd8At/quHRxYrlE1IFGTWhxebP0dZ5PSZnHiSbHnmOa4WLSeJ
/+iOtIC/tTmKPntPev34AMRfeHpkz0N79wAHezlOx+JiblvbbcwxfUNHJiZG
FKix0HD3B1CB3Evewc70MXMxefGEdbFG3KgT9EjtIVNAxwkaZ2C0a9veN8qE
a+pEpke4qikJz1EsU5ucEqe9q9YyqUASfxGmglrhhd2K8vYMWVZyPsiiqqEn
2VsHnsbWD3STnyGYuiT95nTe4oc7ReHFEQZb4axRdGYEHjhAmkhMIhIRgpSM
j6G97mJxo3ppS8R74Qrdnx9+wIBOqysxqEfSTv3x6LRvEUbr/dBukmw36kI9
gJUPM9gDGuzHGeox46MK5lHVwgkcX62ssebP4wp21ymaZFGxOMQTiGB5wfEj
g7KEKqFrRaTvSAlWleqyBA46SHwCZvHATj3XEdH6W8jaf6JNkw9VwRUe3Tlm
DtZ05Sj937CS55xVY20KsQxO2wBcbSDUao2Z3knByqlj+R6munpjS4qgqmE0
tKE21DwXM/nNC+jBCb772J277svZddCPoPGTwebOdI0nEbvJIVdb1hIppeEm
kRGX68zqNn6dU6sEOluucRuOi4j7EtNMwnHyDbcu07rqjOKkmUFvjhOTeeR4
0NvFh2G/caRFWC9TBSokQx+oFRuZp9KVCTedEkNC53FuTV/wW4cwMLrheb52
w5+FBEsVSAcGV0A3TTaGXFYKKKxLKHRvBj4Ha8SFlxIYIy1BUIHK65CDGNJt
YUwx0h5PUNk4XlhCryerjFQ8Hicon1zMaGAS3KDxi5sy5OCtzZAt49xuBygL
ThTO/hnByle8SlxohSV5hSVrNibD/xCajbULchMBSE5f93ibirYB0TjDEHyJ
Kk9dnU/H8n2Ze8rJut1vIUK15lY6tk8jmCXdQtE2BhkT8zhgHcjDPEufhpzV
ijTQwAYFIEMnOdyZBIHwsd1vbBIExP+KpLfrZTTD9nYZSs1JY2Xty4768Ea4
Piop9uUCbdF6hOjbpUSWuw4qA/JXF1XySA5xQBMzdcvO7X4Vs5izIM6gfIcL
oR4MJYeua3b3APbZ56J0VbwYCgWpGpbraKdoiKF9YqBNLAHlqmQyS602/Oee
wNokBwMlVZc2gsObb37vMucl0xI7JpIotbyBjeWDUT8kywJC1hII0MS7U8jx
GhtamlsZkYXRpDIho0sAy/X+c9GjwgZYCQVXZU8eemQM6uh+EuvsG+S3W+OS
iJFYc88baQZRtSADQrvd2Bue7eaE+Ff6VfvTqfWmpgvKh0To5wcCJh2xThp9
uoK1aeLMG/8NHTUKZ8pB9Y8ccHYOS7W6LWv3TXY/BgiljcXvQU65dtajRgZZ
KLB9Ncy3xX9LWyApdgQG6eGD6zF7QL5Hqz26QtW4rpNxbkRvyLwPpKBSio4p
XAfKPkX7MB8Ais06sj76fu1t2da+EAdlN8dOO+PAFWsJP/yFB9YnHPa8yX0E
/n3tJ0Vpj/FWLsvwFQ7ifk68tIKZJhJOzjJWAynGVeDOMOUjM8JOxIPhsx/u
Wuwinc0/EEmSYOL6Sk3G0L/4V+E00sOVoGuI1yI9hjEVJP4Px6+2r8H3lgfb
bHXbugPekQSyFLvr3k+rAnwxsw0XdzriBAn5oygTdTW2YBsuRL7uoYZ0QvYd
1UVQZcJdFQChqbaaeVryrw2psaZ0Fpjdt769LInphyTUMNzFTWKA6mFJr4R/
TtUMmrp/EWEQF2a9f0xpt4c/LodMGKzLVWJ/CPj6LGX+cnQqOeGQhZdArkZ4
YocEHyZgQwXKLJuMYhqD1ZwfBp8Qn+UXwRv0wtlbLRgaw3/DBEVOpoRgyLv7
+Js6q/blPV35LYTLRCnwI0cnb1nd50dTB9Rka4HfFqoDC6vU3bSwx0fe4vY7
yCZBJY+KFpY9+hGrXaF8NWVZiXGAugkn8SKaJLnviRETu/F+Ottj4bf6YI6A
HVxhb695eaWGy7HvlIPI4QqVReGRURY8PYFutJXDSH7uyoNW4lX/FMgf36ZW
PrisD7wcQp7JYF2/jmXpca92fg7KyRwDmc91p8Yd9jIayE6BPz8RAtLLUIma
vXV1fZT04AyrNIjw6bD5LWMK7PItb6wGKEgp8M8Ys43MWDMQRfwk7IpxEn+m
/kqHJkvCz3+uNKmnzF/iJmxrFbbpm6+bPnAf1GzJm6kq1OeAiQ45jgbHqeIt
u3rAoj1Ewm/34JWMs5iIab+vdhuOO06XNFtqxp2+1kia8nz3Rdp4Y6rwcbNz
nXqto/B7iDdDb+0B0Stfo0OSLwyXfyd5g6TsqLUTWOr6PQlUx18tF4p8b8r4
LtXowrQv6iRsGriTj5AR+TYQs2Y2UqzgtFI3oUc9stx73X9h7cHBu8++PmeP
RxmFNdzK+pkSmZxzh4q5n9uHxjZ5ZflErkS0sFCCWCGK2gqBaCq/4/Zi4J0J
n4ICiFZkz0xxBh1pbLTWAQmXGuflqte+wsQ/dC2W04l2bhkg6hnM0h77mo9e
KvHWOqVMoEWkp8GA6YVAWmxxQg0i9ohrSvfspzFUejQf2YcG2qYe0zSphbmR
+ovwCfqf2ko35VpFmbPGF/Y5BHDnugqdYjtAPo0f9hrxqrIqx9wYe8SBQlRe
L4KBSAgvyspboMcVQuBnMoozhDtF++6ohDBacxhqh3Y5mnTJ81jh7+H+gOJF
7kJKPGON6MWBV2/EDrB7JZfaAjVfhseVkj+Bw+bfo0oapRieZtwzIJE/4NH4
uZQ3f9kI8W6nRfqdZQZCG1oXSbYyEtS3KtjVrJrnuFLqYS08azbqGFz+mUJw
YQwaSn5jzHy6jzsWGn0TgRa2XEjMZ54RcZJ1sv9BRhSIXV3l/OmuKHU1UFA0
HZAwdWGRQ/hdiH7N+mStJRzsXuDLK9g5HOK71Ka6BSb69hbszHbWNg+3d2Vg
VBz4t1G8sWAt5mgG6fNHoTYmTgDhj4HVeA8bAW8w6QFABAcT4K6V6WT7FljR
vKGtlvpw2CA1hT7by9plQNqJYSL/1aX1KfK0DuiQ4Ye2VGnHleVhr7cUvNKz
7nzXvoP87sfzY5E5aqY08DCHbRC13wEvGPrM+aY/E7KJgmGKs3ICvzTvkGqV
bq9xTd4GOz1PCcNVjMl2RyJGMoiFak0W0kPpKUF8ZOa5IblXQQOKmv79ifuY
mEPZjP1G8FcFSI9VFDm9KhLAWORi4t/HK320rX5nu4+9qgxdGKuLCi7oRTtZ
d5lFrSzJRB+BJnwSVJhqX/h/adbXAIajeuY04Nzyd8SkVuH/z8xkHRejOoXN
dXzMV5kxwB5LDyKH3aCF7OFYYOoln66PS6t8L/W5EX1WnbMFQ/trtOIAAdv8
fjdNVVpmiL4uUJ2KW7Lp/iSGOHfsfiUGCSCGI/fV/6Lx3CuH0cwZKqUnJ/6p
hlEjy8125FaXeWqHxyAvQwAYoqBR8opS/R9LlZMXNz5U6MJTACt4QQXgKuKY
a5miJB1n0eptKk4u8THTGnchqG0UG/4WNHYLuz3DL8SeJY55uba12S68S9HL
ol7p+7vmW4Qc/F5enP98V40li0MI75f8NdoSH9PUiUOi+a5iOm1k5D1lUKCh
rhgFmp97or8zSKzIi/dgaw7K7U//91mpNFxM7ojsWMvgH+15lQ3bpE45vH3B
3KolQhNWS+WbLwY/kBCXwwP5Q/NOTRcLs4ZkEiQJ4yRL57AXxu0QHOHa51al
KznDkW6wZR0hqe+lR89AzotgHAB3hVgyNn6NCwdIUP/6ozuy8BBKAvBh2u+Y
z/iQ53OLNO8lmpJHS4euMNcGXHYInu8VjpX/aZUo+VjmG1FF8CKvdM0WpF1c
HKL0eu+r+QMkrnlj2qne60aPR/ssQU2hk98KZdE48WvMSw5QUWpSK/CjCVEV
XTtw6bGgQwg2+T2/bOlNQ29vU+LD2nZDHWnGNxiVdKWiiL5SLd41Va6geQji
qqkJmceq7cquLAR32xV6NFN3+r3Km2OCxJZH0BBsQS2OcXKS+2IhQ8jZA6Vv
8MFTIitgYwLeIbbPslb/gmcAPUlItsxBO6+/bZPMOsRWO6xcR3IlLpBoPbLs
zrt3MV8DdY+k7w57YKrQ7SzLQbNQ198PgTrI/QdWHp2QA7gJ4FJJYjUdXFSp
Clky+5n/uIeEYPUV6jq8unH9M7QgoZf6zRqB6Y87U8zGjRKYNLvAPaCGSOOK
7cg0JU4yd4cx/Q8jwaF5px8MKcjFOoJiHdDI2xbnvoRPkmNM8lz8HV1+J/Hh
Z0GDPh6pUeLBnBJZ1EhfoepLXF9skgRhucLGEY9mGIVt3wu1G/JetCio9wEW
Pv6BBtyMvfBiG506pHRBdj6BukurVI6FnL8Jf79KSsZXlkhj/RsmtwDxk5f6
6EPzLEYt6Y0fkdLa/fpl/jv1cGaJj2UPsD3lBnMrDkftefVuealft1jiU98S
6WKqKlZE6I6hM5TiJFgm84J4rFqmdur2mrMRfVgDVOwmxbFRjppXsnzQBUAE
qDGU1kSkRvoLzaxEBXKDC3/V570ORDs5tIUhMeSPyuFyyLIKWsmWgSX9jj3S
GhVNKoqdWYNho/xVQnXiKPEVMeEzL3gHY931ONwwqA0K9qWWLPWhrqX2CIh9
86jEjN7hGUM9XfxyWGheMCsajInUZ9bxcEbwn192bOlWAkmuEvIp1wcaLA0g
XCPcvq3EtNR2e3yDv+IVcLL7snFmm+vGmtP5LMXnQ/2TI+JYxbWOydcnZqSM
/1vWUfl+5uvHvIqALxfZZeNeF/vkN11QmvkNuuUi8EVsVN6IFytk0iybMUz6
pWB+pvfuczxCrwWAXWpnf+NE8J8oXPR/qpJbX9/VIDfTcqo4tsueUUmqjjXJ
ybAI53l27XGNS7f+aAo6htFR6tdn1kGhC0eu4myrzmN7fqwHn8j6egWkAxTA
SkynumlJJqHxlCteixxIimUmBeOmFij+sZT9u3gC0pqC38Nbg1o8J4bXeWwT
7P5urm6I2q8MNzeGsbu+iZLSgPvJQLPEKqES2mYjvJG/KL7WmdxxsMmU9r5r
ZPVgL7fT9OG0kSypZQhKF8r8RFWj+DtXMSyLjMLvvWKa5FFHS5l5TnghJwLZ
ISEeV4ZZGZnoYk5IMhtL1gON2BHy9EfXUdx73kZo2DWqoQXVM3WvLgutbizZ
NwWWmj8b6LbpCiTDlqbxNulRHLaGOnsBSZBk5rElTBN3FcJWLceiaLrq3W6z
y/fc9iUxvJjJ8m/8fINA8d6Dh8uegSNOiydbAfZNxIkVMDaC5q+8T9PcW+ef
zPLwd5rSmb8iziNhcV6URWN6covZCGiktIen/8gTVW4BxtrNdSzFwrydLCO4
smO5+aVi31tK352QcKK9XCCdTif+Vi1mebA3KQtvn8eLtLooAvnNCQFLsBqf
yMG0KqRpTBfCib12/3C7fdyOUt1AKLN9M6dgmr0VHm0KxyCRJQETq/2Jb2p6
NnCaaTnm4vFNQCqDK/BS2EQANJEni3bT0xuy+rlAORSL/0LcVj4mJlyL4Qdd
++DK9mxOxxsnfryaztsd1i6NBmEjuV34yjHouHNoCBBjcljoM8a9mqtUlNZd
9qfopfb22TbJKjq4kiE3AViYjmw8pwttwM96HiAS/KQFzHFfDrsg8XxoEZvS
dTpRyUiE7FJahZk/0w6e+tgberaM3EaT3K878nV4SpDodGBuNyDx94TkQW6M
8zxe9CmmomwUdvYMkhmuNezNdoz3pjdNriHDumjNBICeiiStjkzdOkiajaki
H/nyZ8a1HKszpMBelI7r8VpZ1TdIqwFdlY4cqlt/s6hGfxUJMaH1m7h1elbk
JeTpD5a23R7VVU0hWBLILtty4syUPIS+UXHKfZSYdECkFPcVYoAGeIzWYMFE
yHi0ycfSOacmguRAT9hfIzYylWJO5r+zQqRDSFO3axMk/JxlYkD8kPtLEGqx
XP5IiIN86+x3CNNR3R4CF1vI+rAze1InBppydDvGO9xoPve57OcucZA+l2BB
JocI5Ijqvr1eP+bbVr9Xvj1hUAIO+vRogfwAg88sjb/wycqX9KwA3Mdftixj
PEqEYTeuxKrGwQHbf4B8WWj+ZK1Kk6Iyk5nt/c/zczzrDhSf3k3cb4lyJ3Ef
rT5KHNq6a4j9DUc/wogORZQfxCPwi1gAVTD5E3cZOLM/PhV2MH204RyHJi6N
3KS2GdLOeAamIKevup7WqxBa03a7cc0j8+zfMTxdZkLxYCsOK/N6X0eSL7NY
Tjw+7DflzcXfVzMf1lrV8szHZr4kS+jmnAjyrDoZBj97izCpWhc+sMaE9tMY
ApSI+bzPrPFWcBpBvjvAnXvjD+wRLLdH5H9cNSIAZecVQSbyFVsTRBLky5Bf
9HjHEx66Y4uUSU0FQt7tVVGgOx99h1cRC76IhsjraEAF5ZChsEld5S8ndSzD
G3QQcq+enD5BK1mR563y2yMOpIKElO4LxdP+zcjGYfOfkVRJeyAUH+iWhjre
7pgKa8dRcfSXTJk2MJIfvnGtYCXOA8XF6YfOANB+GL0uszBXVX4vWa+tgFc/
AjCwRxThEZ9WFAJ82BPSvClXLpjp085IfMV9eh3j9W7SMnzeqRJ7j9aiwXKw
KaSpk5HXGUU8ikMslKlelOBKMbez33ilSMVq/wjQHiV00kW4R8yyLv90JMXj
PMOBI8GFXHT4/4NEaUNtwpgVU+8Tsv/Sq8Z8XsC3nhFn1QPyTpYb+iKxkOrN
VxioLBMUkzTA/ig7YoReB0XYRty5uIvkAJxGu8bqzFFAAp7mmO1XfcBF0HO7
bphyEZpfyt4CbcDdbRCWrCkIxcOOSoDbGDdscOLoQBTJKgnGvB+HOk5Wd8sM
u7b65RSIfEFVMfJMpxpRZQn/xFJM2PHXzQFX0Cwi4poYqlXRypDJRp+04fM/
55vQ4UaP3jmTPFnuJtu1a2mFMZ95nS5RDf26JXjx7F617Rua0C9zo3zFYYwg
UisIrqMvnIyqQn6IR91ufZRQqrKWOm3dru6ZQ/P9Tb2cAMogBAWkpV6WEfhd
gwiu856/7UL6rhNgMt4qKSfcOcdu00g0fXVSBkzv1g2py2eSFY+abmsws26q
ojDZv1Ird5PrW0KlagTlUlXM+SIg5C39gCTJfuTJWFQmjrSvzUVXC6eI3yrT
s83FIpeJFNtUhLWma6Mnhe4XmNNXOfqp/25KXs/9IJp4QiCJaq6XnVMzYqJU
zP7CjGSlEmvXLYCL15mME2rp/eqWrwkDpv4D7JkxXTmeHWIeE3qG+APxa3I0
GLY8ZNsbslVJ0jvc8bq0n9HWkSiF7QhSU8Qess5rMaljN1lXawVLlOnWvisL
FTms7X9uMYe3R/vziCw1M2wcNeq1dGEYwY41BhDHH+WC5LHL4C/xpWBugosL
gaqFfZHbrFuLGGGQVHGQ7+mqBvGulBv124cHt6cFc1f09iZcUMoyWkUU0gDE
eRf4a//YDU0vkcaPv5dXhoE/yoT7Ez4fTWJ8aeP60gmYkLsHtlOrE59xlZaR
SsGbCQkJfuhjQnqrjr5auCcMnG3ujYMDvDYF/SbYfPVKMGfmq3sPpxc2uS0J
UwQ5gLBlwT+oz+RuA4sSTFZNvY7tmOPuKJLzmPBhY0sOPM28qDStptrSVsrx
SbNsDpB319yE7nQuOivX3VBF/BjFjoouEC2ySfPey4AyV12bFBycmzcs/aSn
UxfxLB6khlR/uYpq2lt+tw22oadRwu5zrLl10XIZXaXu7QKjJs1idGgTIwU4
ttQQ3asvqxLjJi5VPSNx/wgwvVyKE1eeVWKfaJ7e/gDgXKPetGQf4ZN8u0od
OMKq9QAWi2MG66Pk1+q6bHTNSPrrl4A3fmXlHSAOe3iU+1Mi49RvryKKmut8
t7lV2MZftHL6Bi3mDRQDYaXX6L9hMalAn4sq4Mz0bkiLYD5iJjyqVkgAtgan
5MA/2VSFiGo+35hL+t3MbYkO7FNQlo7NgPUnO7Yl2n8dWIZfYvvKG7fcp29W
FGe8KhrDb86ZRWpPMKRC5kFEzE9194oYFwYFId0LzgYb66bEdPVyWaY/M4r+
r6xETI2SgvunpEUMUzpinXozxAWqeG/+irGClVhyn9ILJINN5i9EO1IAPC04
nqiX3SNaDwNUjOdNFc5XG7Kid6zYDVH0lrOs4Nebz9Uum/zP/jyiKriU7aQW
F+Ze8zErJpNr/1ux2X5luYV6W4utnpWDlqTJogpBRMYAfuh/SG/6ltndaVPW
2MQmV51jQbACwqophSRDDrCHZAZF00gTZDsN6i7PrQ/bawtdwQCOHopFhgvp
Ltre/vx0z4hgIHYVQ8dir0WHsrs6Z4mOuGeVF/2ZGzqhqVSdLjFH8YjNXOuZ
eeINnOKBKLNfGJdrIHJmQ8+tlQJwALIbQuNltfYAbpDkTZWJD5XBGkieeZ+1
HPTfd3ZdJctpOb4qJSxtoxUIJwWefxQjeg9XK7xooNounZNu/KOYEQLXNVNr
9iD6yDqiO/LRFp2pq1HqWqogFzANXWETWnPXtrcgoYIGwj5UahtXCvnn++iP
TBtg7GdwZjhET2qF7JdW6XgaJE4WZ5LlX8QFAFJskomV7tOm3OOK5vN7ysQS
s36E2JsxK8st9hHOCwOxY/2ee02yJaM9vsWwf2u5N9kHUTT+Mv8C5DGxUwXW
8WFhTDzu8lL7qcRNqrKHPpCIJ2ncgGmFII34GSwg0tkQfbOdHLkTqlTUftVI
uxox/Vs7YDb+u9HSkrlrJjawyM3BKcFmDQytvRNZCDgxDhhhmtSU7iQCcfbb
+K2yhDVf1pPy5fO8Yi85rLXntcTaH9F+LbaN7gY8dXI7DCGSwKI7WmkfXq7v
0S9XKKiSf7nZusNwDBOgWSmebas2aYLjnOTsbel3oPV1viv4jV7C/f77KucS
bfceBLzG4n7PH25CdReU4/Vww9A0qk+1NTSX9Is5Hy7Zy0qIDb/9LsxQIHF2
DW4bt18qpj7othe+JiVu0D8R8s41TfgRc3A4enCGrSYAmXJklF70/CYovCfp
NjZRbgr+sIyfceStR3vhljNj8KjnpY7WwBOOG3PTiCmDsD2F92XpH287JCNR
N+H/pRKC5InK8tikNCgF80vGiiyYwfUGZKH6Xgwrmz4pHRIPDMZyRUb176nj
RV/S4BXzwQWRQVm4baP7Sx0vh33X+WLu/eSnlE3HXGzxzjd4co1vCPhzpOj4
4+Z3pRZ9DOGQTmhmQyLbZMX41J1gwTdk8BncNOXxcH8RO/bj5cISqlObsLJ/
AmakXuDpKLrkFhHx2KviwRCCaA/vQJSrEGer3yYdu0ryaaqc756/zn4Klc45
c4LLsGAmgUbNZeRWUhKFnjB5BfgKbeNyiyaX+0ZkNC6EjkIhYBUwflu8vknP
yE/IdP7X4PocNnBARBJpaoq9VXxJCRHD/u9ABHS47aorDe0Z189/TaXYA8uy
lex2XSgljFlw5mq4KLy9lK7+iKSdmuVnyFCXAUO+evNX70qswvlp9a/DlF9y
gbOYzsaYywvDK2mfykfUsWV6D3w4Ork6wTbVVrfX58r+fLe19zj9mPJuMHMj
+XiCxesw/5p+hxqp0Y4KM0vjjOA7dkhFUeoyNI+PoimQe4X+SnmHkqG7nFWx
g1wIEpc4xQ0mTlrx5kvdroWMXbk8/kVk6cVsKkLwtCnGvXnwZIXa792zGF4Y
bAOyxUagx2uLs8MSWAtz4jbyJBI6qaarLKI6vWH2pQQi8gIUtJSpCWN/uUth
/0+zIitxZD/CC83x00aMuqAF+jp4v9D0srFUcKelNJIi8IJKM3TbKrSG1TCt
dNRyN4AoxEKpuHTd8OUfeOXX/lnVncraV87gV+5ejugNp8zOdIrJVqnzCR/0
sxzPbcod4lZvU6C025NYRfTtzIOAqaiN9UZfkifDo4fHKtl8mxsPtMtZVK63
T996qcwO4F466onzGBY75VYc0LV3K+fmqQuyATb+0Gg/i1iXBgakta5F+f14
grCyEy4f8PukrhR67k6upt6wm/0Hu4nmIcwGgXN62NvuLOwWX7PeUIS7YVph
Y7BRz+I8ZcmqTpVMRNYdSmukFWv9PDamaolYR3SJWJj9mVVDz/rV9+fX7iv1
pZtxi/5dvK0LUeavxH+dqcZX4P7io8WAE/QnIjdw4EByGj45bL0jLU+hjMgF
76qLcRrK6VpqBPhs0asj7M3nu3h2QZU71NooNu80bmjPH/KG06hJ25H35zZy
LxD3T3bAO2MVhvxzu1TlNXcIIynsqOkW1K5XZPPGUWdcF1gU0LL8s9wA3EZm
mXzvO/Yjq9Um2udvbmIt6D33OGfPcVxs+j/6oaTq5jZAyCkxsknobGti2VjI
3d/iDVBS3CXg3SOayvQ+4ZgsAVlaa41uDGR4YlKumXHEN/GUTo33vgRXgBjQ
XF4gJlkinh5kVy+6XFtVrQh3EA9nqNzEevg8LqOcZoL99/ngSFHnfl3orXsh
bdWzohipRzJcCSOXSOEBSDOLgCHFk084zMfn6zGbaUhK20FYux9T6ekkre5g
aaQQZ7LUuFtE7X9ky11isv6zjdLirAQG1aly0RpX6ssvT/Hjwql7DJGQBb/l
UbNG3JRH78LT60vSSfo/6sApiCBzFvOqViDqrwxo2TtN/QRSHmGJ7Ghy69Kr
dh9cNDP8K2YCL6Xvv88ZVCorFCzb7onOND6FTE7E+xdcJms09pYdTRa9zVAK
PP/h3Z9ZFBvOmh96Kqfi1NycjU5kGfhlRUKbUA6bTwK3NvYeYoH+FwKOrXrt
U+PgydXYOOsDrAemnGwxcB7A4dwhp/OkiiI8Itqs0tFjFQ12vE2kjMJS1wcD
ASMBC6A1IH+pzrxy2EG9PuYr9WfuBzsvbADRZXmBItQFc1YJy011pIYmaO+K
K7LBygJimDHy2fjf3AaPN/u73cA7mkJnbXMdp+itKeXM2H01tayj4tec4K25
kY8uzKL633c+NxkTYV9Jh+4k3BlqnijmxQK3KjNwsZoaM9p3KTCzTgMoLiTe
s3dYB97ikyRABLhdzmppTkukvWPQmYMNit8mtRd0zSR1QnFp+vn6dcCF3YOC
X4ZavkvJOFQFkoTWJs8WFXSj1GsK+S1scB4sDkDtiLj98T0njkn/3M/lRyU7
O/BCFyhHnDb4zStsdSTHwU4PlR6nkcjUS7PVQeE3oSelkpCPSKFFccQXrFAH
+qVvWsJ+hn6sLmJvSbw8gbELMqGQLc4/G4NDkga4JXzDL6WuyFSwIS6LgBur
T7leAWvpBxibDxKa6tg9lXJIIdeJ/djJHe47PoZX33d4ueDU0NlG3/7W8wjN
SsPT2nfsvab25j6H1gf5GR0U/Afrz3AkDh9dFWr6gPb9Wioo7dk4f4ZPgIWc
vz3rBUpVjtaaGD80hr9IdN3MHCrFQFl5M1CXhZiqwtuyFxRq+2StgO4Jteh/
9Yt3bZtdQrDiGFtIjisZNVcQv/umwG/w59KnY+1ySG8L4LGKLEs/ICBIcQxh
86ogF6JqQL+1pSqB2A85pLaqVB31tQ/MHF2RWQhPyBUJVxDFnDUqdpWQHeeK
is/h9ztioYv73FIyT2tmvxPM4ifjKjCFDv384LqsWiVSaWp0T2FmVfz7dSLn
1R+osBat1/HCPLX5JKwGH/Qq2QnNpFBZX1XFB5AlCcIKW3cLNbP+B1jvN+zj
++jfj4YqZmykd06OaDTsV/Hf06YqKk7XS2oXWVl+8UzSNuFYPu2kWB7voyzO
dac8POcJFgR6eeufh3+fxqu7PGEJqajkrhUMriSunGnW4dXUNSikwvl+svsB
rsFBDLIpInXFfOCgORfB0v83vX2qmVrBaWrNFvNTa7uX8sftglUdgmjOZpcP
nwgwDd0Sa+Z7AMPw+mok1msu7Fs+YHQNFLsuY4ay6X2OS75X7EVQne3g9RWe
6xT/ln0sT9YBGT1irj8Daa/9lnwQpLjOGHfNgttWBqqyjGFO/RITbZ1YfaV+
RdMeUhULYL1BgtdDZy17T/fyIJmQiohwS7CZlmwhrScRVza5rW3p7ytVJZTs
72KKVMQsd2qRNtt6zlxNPCCiVv2/AuaKclPFFoUGDrmDChSPU5DR+G0AVENU
8poIm0WT9U6bCiMaQmRVI8KAClpndPVC7eqp0AQBJZvBzmLdZu1gWFU+0w4r
RemHVYvecX5gxOLQZ0rJN7PZUx4YH4GtH1MEgKFXIMukXloDzT4616yNvabD
zh6LfElKile1miMnJRvj5QtgeMW71QeXwRBzPAAxwdF6LXirwXC9GPCxlU9D
+qCbU/FB4wQ2hx+idF1c9yyCHlcrQCm/laQQY9CG58XF5uLOwVo7q13PXZ1N
sVk6qQi1T2jWApfIGSEwXw56gl8TR8f+Sn579F5joSlJNVHRWnK0jEyhyxFd
NV/xU9Hpe2mWMowL0YkW3rjyGtKITZuEOfZ4THxQ04YBEclM9v3V/c/KCtHQ
lcR1tuX1DTI72YY5SqVu6Cw22P+696Vy3E3q+oaNa3jHMjCEfv6B9oFOGs8k
hIonVBUvq62qT4vl7Cs0v7XV6os7w9066TnHo46jJH5wieFe+FjcHAYOvmPb
LUo4jEDMJHJsTU1NAg0h0YbC5/E6Zcxi5n41eFvP5WhEIxyjDSLo9UipfwGH
080ky1rqqCHYaZehGny6Q9N4+HkAffwCFH1mlD+TFWxeelJBbQDda77opjaI
dS41Z8TZivFL8TcJZdsjpnddIVdUp4EFdVliv+jUI95rV1aUmzytAMIS3fDo
l28b/4GHexn06JqVk+foxpwNsKroPXD8/DifBzpMMJYRnQOFV2/YygVQjTIK
7Noh+XVDClvvpuY71xrP2Zcd1nm5HZvlGzM0HHdBiYAOrZkG27WKi8I4pK8Y
+qVhpYOjnanBwyL1Ze8FBuAmHift7ZB5ngo8i9hswp5J1zlIhFr0H8ZAcVZ7
iGHi2hhRGPHZh6FZoOkXL1E8yY7M0iQ223bCOFZQ6/BLaNcRvXfs9owHtPuD
vk79PZjYwc2W1mufBsn48N3NyuoSuXzZ5+UbsIuKmzPBRK+D7obsx9ctFiDB
1mRGpFitGJXB4f1DLPmSlujNbVlIPMTAjg5TYz8nxSWaP/zOky9pM000oKS0
d7xvHW45XNIBqg5slvvYytSbn8g7SvRx4jSgfILfcWB580qPCtoVk9gYF44t
XspzhTmrINS9cACk4dnXvwgcP7/oeLGfXyZH8qOgivjmPMgcC2L29APzP4df
x2sADX3/RCqWxXctnE45zDCs4Wd0bgcV69WjV0GYHpdx93m0Sj3Fzstpq6CE
rC1wurluWQ0H7lIf1NXLPq0UpNzIlS3RuRvEWMHStFJ44gqs0Pi2u3mH2iDD
pNKS5UXm9qXIgzBh8CwiYfA4nJ4I5vRC+/rMZAUxC72HNKju0LreabjSFcRc
OAVP5ZNY96EE/C3qzKqOr+W3KznN+T91ftzKat8g46atVSI3PDG8xeI8U/jw
xdpXyIioK+HbaRODgtHy89Q8Yd4LZcgQ2GDyJTDPlyrOZ+8q4/9XvrdeSOUB
c1T1R9GAerJVhf5mAHtNR1bjeQJKr4Pa938o37rSix4Xjv7ZnyBOhlU8bFuI
zNom4bThAqZxbWip5LrvUUXVkwtiMuHLU6J/sJwkE2sEVtWa0O82+govBvfj
1gzR3R/C5JTwEZ+MUWZY2Sq8VxpFCdKtL4ygDse0gLi2Lwgt7Os/EGfS9mAs
XFRVSyGddPUgy/A7cgXm81yytmK2oUcSdRX58TbA4zyDd1V/PSFiva/G//Dg
0BWj1XtqFX+pueWWuw9MjjGAHQBo33JLIjUUDf1xFADG1ArG+SOwP1WlIj22
wMGWXBEMpnGz1eIA9br1lV4hCvbUEyu/LKegZzT7kk8S6QxWcjz53TolhsaA
OEOhKaqN5s5KYgIDP+KgUw7SvJELPMk8+xbuJ15+Ut4NiDm2eXobbnmki9vU
W5eCXZ2UxIw0EJFAM1hk4nDJoGJZyYF27Nx44OA7h0nkVrdqk8uAC2+j8z03
B52jf2wCt0SK1SMTyQH0KcwvxUj+HjSTVcPn2NQd8Nllswz+rJltacoTnWwf
MrXZSreaxire80nE+L/XXBp+iYNf5FGVOLsTAQs0Tb3l2uPdQsepKS/xBvo2
IQRWmWJBvbR6VfJbQn28hjux2NnWvynGkh2Bqjg+miFEp1PnHYKcwNUy8+ey
Rc3X4f3MeF1xluHyQqmaUTS3ImIOv/ypxlmGdgLqoVLL5wz8cOPP0rQARD2R
jouLhSVKrs9CgI1c6EE78pUOHupLbGVzljkVOZdNBMbuaLktyhzBkysPTYu4
81+d0yq74c+fnbKkj8DiFARPHc4B/OphtzrHRgoBQEPhwBE8ZhnCwVdcM9r4
TsDpO7wxNteAmxQCyjiv7UhSYE7Io+7xYh923mQP5SJcTLUif5yRHLgswJ2f
CIhGtOC/wvDVdw9TSZHsbyNXVbBuGULI3RAUkXxvtxAhZuRkFNEL80bp9RKP
e7F6cjj9lXxBmkIR9smHT8R7j+dlk5p/dzTK8urahlHW4CQbNl5s9e0hieO4
8gqidtZQGO5e3OfOH5O2mdplg25emKmegMoSZTGCkhgmjUFweuitmW1HCNDx
uHaImEX5q5aHjJLlsX6JzggqMl02rbwpBRj3LMrU3PgIWkT9bQZ5Z33/JCnY
4r8OyYzRHs+Q3nOLjmldbhCn4xWE4bRtGL4tU4ld0BeBdx8ZBXalDwWi0GcV
jLLcQKZEs5JaOkEyI7den7TA88OPFcBBdKcsvIPI/KHbjAJbmEGQsAK8IWg3
nqglY6GiVTnUK6bF/2iT5IpPQLapBRPwvFxyq8Ui7AI64IMEjp4KjeDmX511
Qx7xZ9gu19MsdrwyLkh28ndcDttvCYdyTL+GGt2cdwfCoi0lXFOLmh+3O+4C
w6SbW8LfOjSdhJ2QBug1SDuChw1YlWc2IsoPpjqU5rvjfVX/dkckIfNIS7wK
i5cBl5EBJrHDZ9qawCRUx4P9T6xIcBATEhgEgCinEQYkkaRPfEKH+eilkSND
KNroW8MY1JxTHOMdHjpKytxA9fanYimpOOiIgU9V+iCyfgAnpSPsnJa5Cns6
6+73ecrG188sPTDx+52l3OLwIjt3JN+ChCdHBIY5K7NGIIo+2eMh4uuTau8k
MneTBE6iDKKLieTgBj6YYTQqTdBpfufYz2HD19r/JGOZWC7mdTW+OOE1cf/9
s50ZWLbrApHzO1yfHNHT+ejlxgSRwnbmiPVdAN4nJAu5y7Xk/rxDeayZQK9k
At/YyClZ7KW8o4xDdZqkocG5qksRUFJnXzHZxdqFHC+9T3VxhNze63l7antW
hZCec4kfCB535ZHjl3XTNzQyNJdAh9ldzFHurse/6VMp4O2B4hn3+bdu7xnS
w960/i8XSvp//kZ6GhO7HVwcZytE5AqI4wml9bftSnQmGb+hJ2Hko064b4hm
RGsHltZEnf1qsP/QfxLohcIbtZxUqXL5dr1WpL7IxUM8E5dKkqbyMItUiJxc
LcQBomR350jtRXEvv4G8geMFQ4ghpb1PpjM0HffHrbUB/p/OS+qceC4h4xa1
jN5YqI8obuZWKcxnZGFlfOXvI/DVUX9+WV5WfBpWkl4UDrPlTWEI2KHEBpX6
Qox+wEoLVibFmb74RBP62gepBuXCCmduZ/Jh6DRUNFhyEd/j+Pr4W55jm7QC
9Gyl4XXZ4mGhi7+gEem6aquF7+zkJPlvfOF+naTGCtEcI6zePCUQDKV2Vikd
GOlUrLFWreX/kRzyPlCfBtgzc1LHrZSVz9xsAVPRZn7QQQZdeZ32ffTKvleW
p2j06iRRqz1i+L6a3yAOrTCm4eyKTxLedojJkj+WNTz3X0zZGUehGWzw8LXY
ptPWqJNNAhJfq1T8XeSh2cnBkYm68BEGMKU9gn00jAPRukn2Q5vZ7Vy7CQky
K2i1cg6E1ZUXJaMaNENfMWgKfQ9w8QDnxW49ULEPRBt8Jnh1bNioeBmO5j8+
FOD2Zx3lOiQZ7l0f6CL6ZNxTvTadXXKX8kZXpgoA/aNynWXMEvg0mqeZHexE
bVCHXrkO4UIHBKBcra7kmSwa89iPzxFxkSVfbDZhw1zv2f64+77UeTHFFjVS
HqqdZNEer8ZKXJFAZlkhJkhiR0XrhQGWdOVBidSU1ikKiq8z6HLf3KGoQx5w
6oN5X7jZPVIhy6NG7i/ELzceF702adKhcva5rQSNN9Lqe2czcmgEpw9P+a38
aJ4znXm/dYkjQjlFjxlQue7mRYssItodCioxLSSd2R5Wijlo6xsgGM5Qf59Y
ACDr1N/lUSXuiL+aEQIMXky4HIrja195i8A5Ak+GFWwjX9cvdo3QbN4IfNc4
UvXUvHuzBrIMnIsif2zhxWd/rLYb2cmyShRvGuITLjEEpOeBKJW54G2Ffh/b
grPDpro3hwXA/6BCsATyzJh2o7mmXhzjlgbtqu7GGSWbxd8fCaQsd0rW0A15
6hcLO2ft0puzIwv56g9L9JBZUddcneMKSs4x713ZVdl0cFyg+9o1DaErU32I
4LuhGAJmb6K3jeug6irNDTHS3FNCS2b66mv0TKkG3uGrCE2+yKCgVuvoIZIp
fXWQJUd+eJ0NSfYzErn7NC1D0dgq9j6GMbFgLujsLImtPV1UN4hHJEsQNuA4
icZDQbBwfA9NypGABocRaAyxz33ow5jO0KHa+lyEysfhCyH/OKt9eHZ3G/n6
gFTl0zdL2OhWJLzCZBXaNR5LHrCJwbYmIqC3n9VKAIzDOa0Ap5S/QcPs7hWg
G/90zAT2Qu9nt4zeZhwhtG5u5xHqXv9Y/h9Lp9Ba8ov2gwxqSaXhbMvCXhpR
4SerF1yxtgGaFDMbUUo9B9efb2yPV0KB36/p4YSQeU1ZauGpW/MUFruk/f0s
7TUDiub3Uuwi9tWMLvE9wPf9ewLMoDe42cVbGMlxWpgpiZChr5uhFHx7Jt0Y
FmXqcj0pHY+cDaLiVRhjP3UM6ooNAC2CQW39hf/9pPD0BJl0kGu+ZINw8cNi
Ja+IObOOlvE4jzERYG0cA15KqvGY2rKB+PRGSAWftoiPO4VaCQi6ItmQahDO
O06wHtN/W1dcq7y+uqynKescyXzB2EiKu2OwZFp+H92JJSKkCeMhJIIALhH2
4kfIJigvUMkNdo/gYju1+bgWq6KXvA8mPTLqY9AKssEBs8+Ll1RosyoTE7M8
0uxaftaSrOXRmaSMFGy23pKsbRQKtPMyBJREb+RUIgD/8t+3cCQTcwZsxMdb
lLOybWBxiM0xpDRtaOV2ThDqhyDjh/jNfRw2p0WybF/GGBkMRaRZv01QoIwQ
bD145i78NB+MMM/J+XB2Mrt/317TIPwYZYrJIS84WsmRcUPL+ZMVFrFxLL2R
hKeHP4yTqzhgMkGPVHSaKuvENClxq6BTd2+bbhqfay10br7W/913rwBXGlTB
nQ3GcGlnB4Uc4iJaNz+RqkuLZhkj65MsTyLIlj8UIC2Y6LSkpp1dMZhN86kG
Q+j1nKyFveRtjg2DmeEiJWCOq/wJIsKQSfwGN+fJg+i9aK+1OnYum8/bMsAN
sjDkk3DtJoybG214nRrZGrHD5UKAnfnuYm50nyv0YzgWfJQT3hDwu8vNQ3IM
4VZK9n2DJV8mcaWXIjIp+DwrTR+N3qSipfFn5+gqqQKlEkOL9SiD6/Kiw0Yd
11qQrDQSD5LCEI7ONG0edmbH7Pa2YonqW8ODUezovsvSmJpiZMgIVXFt/wP2
SFUSeFHKF3/WzEhWll8F3hj7cR+/xNoA/mryb+ndmLkItjq3ctNmUjBRAPzG
Dy4/WWYDcQ4ch6bXRdnqT0B96PLvz8T4+dVkqe3FT5A6igIKeLjrznT51MpP
ZChXQTQmsAYjIYNyyDIc2875UkO7itvLupn52SkdjyCYblRoeuRyThaSbUX4
z7Xn2UZwYJVRt9vWlJXgKKieY5qntkZ78YcwD6yADeFyoB6dzFU0JnPq8nUg
5e5Hp94r1wrKITctCvwLLAua4rMyxn0/BRl7iCyzzaZ0NWzv+tBFQnP31tHA
XnYfKHUHVT96qfiiLyuX4jdQz5YhQuW17Ug8OkDXUyB5GxNfmhCbZMBTA+Ag
FWpk7ibX9YfxvstrDAQirR22xAJ0DD9j+r8eLAnIi0t+/pOMAkSacPMBx0E4
NwfLcfGJInKwhmc527xj4Zowkk0UW9oVOASk3MxR/1Ckhmsqq74vrUOjIQgn
jOeDBfxDwLgJHq0zWiG3TTP7CHyGqQ5pyAxCsaiCb73n9fLudL4Q3sPXyaDt
EfUYqXa3U9wtifkgDMgVuy0HXVCZpHRYfkeNAsZlO7IKGAZhT65jerA4sPKS
fck/lKxYRb25PTO3ebRxjvHYtWWGuh7r9flYq4Dol+qPvCWIaafozerjz41b
EGp0cugEZdFErhb5vyd6OSov1dQ6SphYsOYBXGDbxeQvv0ODrG/XswlyHOr3
2p7GTZrROd33EcrGpmK09kU+tq8TK9xK1VQuAZ20a7ZJQTUm6WXc13QxW1kV
K8jAni6UePcwIDpT83zaz+H1G7YuPpebqNb8ETKcJTH/xkkLy2k5CUn5HWgk
mPQjb+mlFhX+GSH6S9dTSdaEI4bmUMRdDbnaRcw/A5/HZksm8mTHNwD8yYAw
RlWpCVS4afYUdDY8mudXD559vARGsw0D1/QFJMBl5M9woEnsKsIfRTIiZm/S
3wdTFfKgzyWWVU7cPCxlgEAFzACf/pwRIpp6TwNHGuMFj1dDXQjbeJydIV2M
kSDm5zcmscdkdyGXDmKpR8huv3G3mQZnk/vju5EkB5HEt78IlZ5WZUuS2ttL
mTuursN8KmSi5UqOj7Il90qMUMbe5g3WpQjPTuIOmq8/MMkrt0AZN5a8AYRR
IMOmn8y+7jWsKe9Cj2dP3y1v9gaqKSDjdGY/qfymZ/hUXXM7BU8dOU0pe12B
4OSLl/PrcLTODOWDYz7ycZ5tGMauXmqFaGw04b/Z5DxXbZA6KFmve2kBpI0P
3KX3KeyFHbTYEtEzjgfkfz8TKfTY4kwVvhh6k/fZ8sq/a93BfDCKg38t0T7v
4isGDSU6yoqWiQyxTzB/G/KzDUOcB3426iLObhU8eIgjMFp7H1ftHuwB6cQs
3OGgyPAj+oJYOCqJ4KpcoMqmx/jdd4JA8RGRbVqBBVsMuWSY3U8jHBiDP5tN
p/tx3m0gqOZl+SjMjesl1pxeroyZya5PDVotAx9HJx0xwV2MY85lJgpCyeso
w+8zilZC849AF6s1ItWTxIq8rI2rQ/MuNGqraCPncpEXJNtgNK77LYmtHn9S
1XsURqzw5T52bJsutSywkJcxpbCA+oF7mYKdOcfJyKROg0JJKWQjU9Z4HcVL
OgFRjPAhNRtksTKl3g+b+fi2jpUhy2KMDGIp7odzsCBzlxUskXDvksuenwxo
uPTRvlSt+45H+OwtFfEV2xH3W13Lx97GHUCIyZRzJCn7AWXyp1sITg0qEXKi
4B3AENzkJhY0LQhZaJOciLutC0Ni5gUWgeqt7W4hjg7iJ2ZIVZ6e1Wpp6MHR
gKUIsgLfjsyFqRLtOCdxCZjYet/Gibmsjx1KKAAoeB0IE+q8Uy+9eJcdPbbJ
+C6L6tEhCHXvq4i1UQZt3EVWJ2oNEw6EKWi+k6wdanBJavVOgpo0xJTzixiR
zjelsKOPuuulIFWPtOBS884JOChBzmCtqGFiNYa8xODy8r6QT1epgulQC1B4
Kf1QvqXRVZQm2dV7JhsmqRbW3VIsSfXl4qdWcH7XSKM6d8i/he+nbfmC3rvG
euY1DuaLPDzjRx81mkKZYBWlTBj2+BiC5x9iKN432wELCGv9hx5FSiRpQ8vS
XGm7aXLw6oyoSWEXURU630aTs6jeEHyFyh5qs62d34kPUjU0Kx5HVx5uzycM
hvSiGMkfn8oRm9Ol6RXeNBv2nXZeVY9HTJlzjEqDEYseLSCVz689kA1ASrYA
LHtazKSJ+9AL8qb6hCGWm5S86yIyM0HT0ynQ/au546q2IV7FKSiVQMsS0og7
x9jvDPONDuNrKAy4Q2QXwebeTnvWykf6qaQMzeIBWC9lnBvd/xXySNn0V7VH
F5ttKvEChDyEVb05zFKHhX1Mgb0gl620K/9bCjXNWPW/39AQy2L9MoqGFwCx
UMLGO4EDHkebEJAtDZEQEiLpLCYyiHSs6dQMx7SN7OhHM1JLpOiBgQ69uh8V
NmpXAsYuqCDd5OVk6UCB9yHL4XePCBJt8EfUn9X9/eZNdxKg/OJJwprITpIm
B2aepxUu75MYaZz5YBYDt1m6tUw3EgSWiIf7JPaS1GLOHfBBXiK2kQ+ivBp0
FFjliv2SE/O4meNR4Q2STEk/lF+v2pTmIG3pQfTKoKYKXWvyvqeb4xJgr9oH
F6jILRxCZAdMUGWxMpGrv4wVFX55PkNnL/joOonM2NAVA99xU/Tu1z7N3cq+
hF4qf0OHJ7OamwUa8pwxmO4I7TBF5H1m4HhPALlrlOe4+UNXpRqwfmGhfqeL
ZjlSdqIOhbthNqpnR9ugbZGGrH+JLB0Tat47A81K+t0eBAhhylNj0EPnVSag
floX32SxUu2DzsfvC5xsbNmZO1HvC1TFi8DWMYf65FlE2Fj1DBspdvsscF0V
mAxIDsT2gAosdCAMUzX3rTtp2ilPUpazWnttNkL86P34w6tWycIa46i2FIqY
xVRxQMwwaPD3FhpYG9jBCgLByY3M+cCjCi2KDSjOMOqXZgN0BiJnXLmELaeu
rCRCi/a4V435WZxLw/l99BDxyGj2Oi1rVK4EMPm3Fy/iY6nDMLEZrrZKx1cw
dKyN1usXMMoVkZxLhUYSIftkXsNvrIfZlM/zHaB8dqmmZBwrSJOIL7cezQA3
WG+5Ekl+a2pSVYhR2Q9pJpAZzi1p+1cnIYcPKj3ruq1y+eRXN7a3JovkSLeN
WdxcH3SfxpjzlcvxO1ZEexC2Dr0tEOlx5F9dQcp4taxkEWAkLq6dY0djgm4X
B3DLK7zwBlV5AOypwkgvxHYSaKDbM1JlK+9V4USdRmhn/beUXbqmgofbicMi
UAgyxyCahKeuh8s783zK+9Q2zhWUxyjOduEKEcAEqAxAmqcTeMVDQpucGKP6
zsK86W5yGOdU/RdIfAYAVp0bM6a33dPaYkuhKKZh9coEIFcS94Q1q11DkxWz
I8vUf+Ct/aA2qgN5t+kb83TAv7F/WTHxXdCd4KjUZs4Ths4+2HaxpAipZF3r
TdtrQuR4s6bwjkSizfhBEZalZoXPMdXQMymmsohONU2U1lmwqEjEaf95GO5C
N9BDW+Z/vvRuXE4Y10+fs812tRMe3TWtX1pHNL/+0SyTcEoGLdX0svJjGVzb
WsAm3JpFP1NYkhP8A/UpQf83dfPLwwI6py/wClVerhyiUlBZuYn6EQfZTjzg
1ZYoyDIjzPwiWzlOaXi0zbMLo10wt7DN/KQIHoq/fI7GFoFVPp71lcUvRK5r
agDm5XSL8dAOL1d+panPkTXkjRrldbe91s299xA1ZynkjT3QXtaOwhK/GXvq
7xDf17HEfd+1xEiblUHojYHu6xtdzORCuJwbd/GLjKWm0jJApgKMGGkDQhm1
QnEQe6H3BKhe+8HOYfs/2peDgFIA+lmbKWQ9no6tfxR/kh60aUgA04jbUN8u
CdBROs3+DR7IU/8I+/SUeXLh26oDSaf2bBNSIhHKP5/LLowYzKU5+kNlrbjK
sLNr8zL/ZzjVlcd3vbNFcnpV8Ua8IkQcCQujB7Zh3i0finTm0AudD/DGox6+
M877MiKNPP9ibmI3eLdZE5pZa53cE3rjPVPjDffeABb94aBlAMWA/jxMJkGa
DYrdArNPl5Br6rRjjqS7f9QOAAeToCxwVnmENxnmqUG+ub2pSB/oIza0yoj2
/jaZXtOH+Qh1kcVC1k5/IuXJKTTQIa2Yif2wtFXf5ch3d9RSBqQcAeRA64pb
jrGkEF+gbXF8gc+RMwNFSdfrZrYlI8YW+dFp4RL21rwAWo1I1of0wZuop0gq
QUxrOz9CI2omgTT4NIEo0B0847I1Muzqceu7zEJhKlfzLj0mEVjx9n5Mjkbl
3cPwFAJj5DI2yVg1V8iynBEuJ/kcppvW6SHnCPw1LONnbQZM5rx70Cpq+qTG
TUnB2slsSiIpOeta7qCzpwhbUq4kgUoxd/Y0FVdJC9Fr0/cMNPfHkStPdtBi
iqNonCkTi+jsR3u3Fu1JZpMw1/dQHQw53sPCY8RDb50H7Vj9ciPUqNG6p70r
DVPL18F2Xyk0mIIwRM9V+Ym7dqCYhrVMfAEBA+XiO6aobSV5yRqp0xmMJWY4
QJKQNuI9nWn4nyfcXw/VyrLXrXKNxdheAcud+UjueYahuS5NiCO78VqBbf2t
+4LJTDT1fZp/0EjcpgMqcP54S2t2Rcb/xqdhUKyr+sYrSPR3MxyE6CequKoG
s+7qd1sEJVz5ECpnwy7SfT/b9xH715I3Hjmt2oiH7UwLeR2PjFpZdwXxPJMg
smltzKwpLQ+kXBJdznNPypS+7VkQdGw2Q4H91Barlq4z5TYd0FifDT0Uf23N
hd+8uFxpSaIXsnU5WuIIsSyUlFDDrS36NGykBOLw9qU8GFqpMEpY+HJbwALs
ScQQxOzvpJtskp2epicgC+xvECxv0IWHSW30kcDnCsK82v13cPyfUjF78ez9
09NpNEDycU4Rwlf/It7XwJeCvT8t2iHqNTK9/1t/MLOGp2Mm9mVc/+Wzn3C0
+eYxU1YflENLsJswx3O33LSWHVzqFwG44+DOpjfLX575ZKTRE73eHXy6RNsX
jy/4ugAp7c4+fgxM3E9iQcBf2OmsW7BHZX9/mRMQ6HGfi3cbvZ/zwNhF89uQ
d092ViY7DBhYk49bFLS/EgsMg76cpXUDAEhJIQspNOa5tLvXkr6U9Za3uX9k
v+ijzBL7cbOKBdUhhleBLKCUJ+E8YRTGuY9mHF/d7Cn1v9LvqtS1j28dTS/w
fx1xlY5a67hxFQHAH4AsYtGchp5NbJr2OfJvjtx2JpQoJz43Rq02U2/XNNTS
NtFAGjo5THo6hDYwX7V1UiSfrcN4uJ5zZZTuKU8ypaqryEzopiZTwWqPHuvX
wx/pPm6fAUVegQI/SQOb6kMO5DIPQq/YxxsWa07rI1kAwOj7Ci1WRabHLui5
lF1iHhY6f4FRnpj7x/nE1rAVlvhsYMqEiOzsq7Ub9MWtmfdBgZ/dN9Nw8/4K
EJm4Z4wPtaxosefoK4HedvF7Q6IVXX/tsUtCsjFgQhuGUTued7pIOLZEbNnd
5gCxWvNiGZmfW1r6//UOvRM91XxGkaWp1KXigjiWQuQtGEsxZDkM57HL4VaD
4WfBpsp/kSBsTqVWZiP3DrUQXJ5X44VGWPaLJoRxkYyfF2TcqdjBWVcuC7bC
nn79WBFMScCoiUzUj0e1aq5nSb2nvZjZbH0/NZqWj8J7niXy9gyl6BkWT1FW
wguNC8c3WfJHt9FKs9z6VehH2gP4iywuklp/PF+CgAq6YUFktNBDrz+vVyle
DNDiMo7vkiw3+nNFtAZcyKtKC4WHsGwLDCxj1rY5iOpiNameC2U/TsBl6TYv
Hxek97mlrYskTWSJFFOoiSkDhw20HnVrny6I3547osTXXoNG+srikFlbX4yv
aXGlWOnXPXnG6PUUWJRO7OscnfmEbx8EDdLD+bLnCl55slz08nHZed38/RNq
BHV7OfgbdiJqbqUQRu6WVpxWDhs5+tzNxs3+uNFaRJMSdjEURWSrypmo2ZvU
riN/dYs+tS1oBOxsMW1uyL1IjEexsZ1bFIcMrZz8sU5rXtIS6N268B1Sphuj
600ND1trgo2CFu3dvhECe8z0FNVktAIRDFMiuG9oNZxJC2VFX9gWIpAQH6vH
/ojVnjIm4XFxeeD6yq07R5B9/HR9DY/MYQjkUYTEhjDdK7A9GRZjiiKnyGYH
QEfOU1d6/AbdOz1WjLwCpoBiHIFcCl/VVm6ZeTyzJFdeZ+YeAmN1lZK58Fsj
pS5xhg6VyIRECPtV/Q7Aav9wxMuiaGwb8aII4AdzMSbM4hQHU/4Cn17dUgMy
laL3Z5Qh66gtYs7KUc7PLrLXWOXP14H+gmbbHVWjWo1l4vqs9V7RMJ1eYxl1
58Ne0DSzmyIgYValPSnTrPO7R1iijn7n1YJpiCbNq/hct5TBoLhphaF2TLjF
ZK3zyGXjh05ar8fGXJmbN+JL7drxZ8S+75Geejafi7ijR7MIKQcpNxSuzvGh
37x6W0RhJ5cHkF7BiGsISsEH/q7u1exnuHjcjuqqAxl/qao3+3QPB7BnnX1h
WJCB9kaQYIakzullHa7z3jNrZmqulAWKzbsTMPfeLqRGkZkg0oWyEXEAOeaT
jdJxMAiRZ9sJOdMHdnLB2SkEXX7/9Mbr32LrrQVDT1ZsLzamKrkwLATxbBEv
uNZ/25NiUd7TAChcM5BN8HxlUezd5Zb/ehHxqF/6hAwr6D/OF8oGCTjOtIdO
Aq/I3fuCxO/YNE+ghFBP2yhy4XxivW2+qJHlFLw8Dt/Vv4asrT/nRAwS4qRO
2diLtjF+1CdRQncbprSOA1dcnNioXdieXRaLggsZB1sLOfuESiBCapkxfLSC
6zxiwplvmeSBgE5xvV7tbcxbnesZNkPd2gT5cXAe4YTNGROoKiRXOM2DDaTL
FZDuFNlR3/7LxN7gxBprxRDLoZUFFbqtXzZRO7wAHdm9m662ZHEp4QVFR+KN
frY5ZvH1WBiBxTntkM0QwuEJK0lASSsuBJQkHVxAjozypChXvQwvROhG0rRr
UJCbp0BVm3ltGPrKHTCZXP1Lp54qXlle2/t3L4oOKsuFYVvWRgRI2A24g0vX
HYPbAw+bjEwXdTRt2E9septOgw5y+wUAUEm48cAI+bEALqxFwPtdLVKmXwZQ
VssibBR0tbC2gSmz3iJv3RZpcHtVG3720cRJi2XqobLoGQPCAsSfWtktmiBy
mIhdtbpRiLqsIbLcu2l/39oK/KtuT8A/PSTbNQnhgkKSZz0CkLWWu/x98EZJ
7A5qiMJeuOHvx/FivEPHDF7A1oRu/pUQGg6Y47mxHyQKHe1BTX4e1DrtY/ce
Ns80hZdEyWWdIN1zMmLdCgVlu0xvh7fBjMw2HapOuHA7As93hch4+xQi1S47
PeSTq6D4OYC1R6BqZiZEXAT8DDogYetNbwT2Vwypxcm4Rn730b623jOZpMmo
MG4flcH6iYOyZ/PmOh5dRWRjSMPLEAhtqa0Jwm+Osql78WXMUH/hW3rG3RF/
lFiBtuAJtir9oxHLrpxI1IyfvYouAf+ZeSsCDxovHEAUFqlUMoLtfhOdk+S7
yrWrYnbLmdgePXKAop7SQrnx/oYTUt8Cy8SuheNNOQvBlNJNOHdI5j/v5fYW
E97qwez2um0UEPDPHspwdUNbotBQ1iraTfjddhFjvfj/MVNghjUjZwwzOEMK
1tnhcbS4vIBwHRg9suGar3VuOl9fmr7hZhdvGlb9yFhrOVxp+aS+maG/pDZK
k8MsD7vsHSTO3dpb73aMYRDxbwUyBG6Y8TDQtmK6mhPKN2sQCvMgR0JT+6MU
RhaUyLfZP0D+me+xIdeUrEh7n5d8vSTGk5ti6iumVlAvH2uqZK/btkPxCRXj
zH/FimBqZ81YTXVX1/OSvQUVusgUiEtkKiJ1KRSLns2rYuH+d0BE1zwQ6vNH
HBFVjWxJFR6z2hwqmwUz5907J8354DvArDVmadjdrzXz80Wfz2cKYH1UiB4X
Mdsp0cuRvsz+5dV0WBNPO5JAoIizNGpH39SpQEWr71vlKXmOrYthvLTiGa+9
VPNer6YE7a4kRTv1RyftAZq52NGbZ3Dh+WI0b1QM5PvcDirRX8heBfCqbszF
hiPE5iHjal4LIaU2erZ6VHdAGk0mbrB0PQDBh42ql+Vr88R5mUwWPYhpJTxJ
GFenq3JuGfUDCNc2/yuyognkyD/MJVDxFVpjUFnvUo+rsbDfa+iTl+oq6Vka
WwobaDnuG4MvHL7FqFAbUfTEcT6/qzUh969xw+vstmcD+ps0LrzlBpxArV9J
iECRlrhLTj63gCM4Ef28tNJkhwR4EOBUx/07TL/XOnXDu/bEIxQpVNPYfFCH
LRk6eqVCj38ZMrKmkW+vTbKJ5Ulw6BQKUoSel68hk8r4HbqaylwPdhyrFIp7
Ohbl0eRs0x4GrCHPlnwlqDMX8HDi8nvsU8S7y1patYBeD65ZKiwjCBSRxSjr
mNuM21ZFgB2cWq5aR+ZtseEiv1gWflOQPa1ijXxEKnU4HGg4/nWgK7Y/G4uG
kaOYt5UVcztvqeKw5eFnq1BU1Ezdfu58C+gQGmVqUZRf3T7goasc64A/ut1J
lwXj0oKELnfxcKkrcRsjFMSuxD5w3eoiCWheeXjl0GMNm8cC2H/8jNsPAEnR
Rdj583ocrkDBjlXiqsaAellXsaUXSeE8ITqKecqYvu1EmHHLh9KfJWDgN8No
lSG9jqJRED3RPJWW37ByoyRoRNY+e44yFZD4p7lijqoXpXRd8WI0PvRsOjWy
5nH1J0m+DEO/QT55O2X3AMREP/zjji4DFrGjOL3ntHqMTNRLj7zik7yWQogb
9mFY956s4juBRx4/pOwOP2jUjt2QPPl9y89xtTs5Ac3wHnYLD3u3VUguI+iP
xZy1yt3Gp/ti7lxNPTubtlUgexVKuKT8f4jemnQPIhRkFQjuWlb0Jb0nu7Ys
a+Q9bli6u2POY62EdZwgiBHjg7PhsifBgg/SA5jCYLFEksCa2D3i+GkxXivO
qaoZYVGKPVKQRkdY2lepPVmgdGOQXV7RmgafDPR2BERUgR+YP+2XTlwIwBzw
eyARFHPT6F6Bdi7yUnSnMA9oiLVM6H97SMRX3tVfF3oNc0vADlMWYPpFTApE
aXMKuMDEMA7an7nUPJmkIT6O+k/9Nv6CzgusbEO4vWf2N/7G37/cEZqNQE7A
fqw8NC4wNHZV1KT8ieN6z1/5lY309ERJbiqXd2/a8/iyW4hIy28K7Q1StSTK
U+Prk3o/vXDZYd5v4Wo35PF4u4KznAdDlKVQ478flxorZn3p9sVBTbHKh7Ow
Dob19/Jyb79kZM/9JcbBIvhGI2y/MUUkYpeR+72zPWL+VdtOL1/zPkA7nvA9
sf6cOkI2aGz/4hdmog52zh4Gp2Z5aALIgqakTNEA9QW56U2AmNd/FoFCYmvV
dJDtlPORX3sE4vc7DilCMk/2eABygzTTelLVW+0waqJPss5uDPgn/WTakclB
nQWZbnn9bLuwoGln5nrtqjZPxspI9rSgruMbiHioCYuRiLpbP3x60c8l+Eya
uw/4aSbUm944AdCPsTGSYZKJGQE8Fa1lz73mSAOzmzK2kE6TlXF/pjvQGerK
mQLXTDGDHnd1/eU0Sufvkth7Ru3BJ/i2y2yY1YqdSs2UKGEj0JHYnVLlCe2L
9iLq37O79O2W6oMaOVrbSwcXJDAIGJl0KSlda94kjxUnSmyMxdvePjDAhr3a
WTdcfjsGcu1czA2jO5xFimUu7MHKucjJfKouNEgrjXEWhKbsepcsOQipw+pg
vjCAfNtfwE0wsdqz1DigzBF44A9HbY3jr1ejXcuEyUw0AEGQqFqYCRXdqDwg
ntHz44GGSj6mjeqsfJn46EtCcevCBn3gA4qsxj8RGstaTxo3jUttke7qTO43
HElnORHE+Sd39WOYab4ij8zM4mC0hkbYe48Lh2qoiPBt5SNYiSWAiEbLiimK
hjvzMCUEEvGnmvzjZNQHJhKzXm6hhPtIfP8s1fPlQn9kO8DCNQs8Xj8HUfYA
cktqmBryu+xqESv4yvLB36emMr2nGdOdzps7+Dmn0lcDYlSobcjYp0KqubTc
QzUt33c7gb9i/zQQEv7va5igmJH/CZLnn7TTlmJJ1rtTtk7JuJfI9fSqL+5x
PYwK/b3sQ/tVrk0qiGVvVPB6E/stSXBdHDiiQLSiyOm2x0DKL0vYG57L9ZzI
augm0oGxFJQuPK4okWc5oN0odspiLq827q+MlMaDpLj4aieYU8kK8/10jN0t
SmPeqfmTA5J6LEplpwNQ1iElH01GKpsQgEd5I1TY5U/UO7duO04qg771uCbB
Ri0+QyxeufZQXdYR2662s4vtsmN2mL/CPQudzcdURTgBtg27K1m8ycsjbsGP
ehsb+xwXjGuj2QvD11fGLDV0FLDvqi8QDFQs8giYbbk7NOsyvY1w+9qgT30i
KtjspajhAxvA3WljwO1U0h+HkbkMKH1nlv6MwjikVzDRpEp0eA3QFp+d8IK8
cTpSN/WHVQLhdthbXVua1u/96Rpp0Hl8f4eh9xua9EBZqUF5Kvv9RTrW3qTw
owewAou05RpK1YwBE9qJUgb8ldQNcNzGnbdJW7rxRORfBh9Wl082RBgrJU6T
k73kOfYTNr8yPdxpjgKzi6SoxsSijv5us6DoThJAmjq24anPCATbA51wvYu1
FDiGV/zFoRRhMNX0BkdIqwIrPZbAXDqoUVB1vCWWfyxWo3G1NaKKTfPWJPYB
wxS5ftihJVfzsMoyM0K4VEho1fq5qyu/mb8S3Kwr2k23IQSbSwUiw+FojkL6
Jg68TD8ZZ3R//22ae7F58y2Lq6NGIPPGLt8lEQ1rShNNs+0xrZ0UDsSkwkY2
CPwcwlgRR5Vw1tkdW9VzFrwcvCwQgwxJ2fWXfD3yR4L09x+uzXiV1y+AYnLA
5slTDHrZEN2Fs0LmiCGALhhpZBqR5JaD02zlcE/r5kk81ePLuAFzzseH3HVp
nDXOQySZq6v4iD66BDxnIgIkHSGEk4pKhay/2ws7Coj9sYWxf5AvzftmP7Wd
8ftXwQJCQfqN0hMyQS4ZBwS8Gwy5uDS47DKJX3BVg5LR9ziRcwelXdtFRksQ
aAr6AHhv6AcV5PRG+UBQxSkYj3zG6FpGb11aioo0Cj2GbepktrG6aWt101aO
KZN4FMaCVBb2VtmvndFlclfyYFbS09W4ZpVA+SQJYEfZ7q6VEHkE5kOhwPS4
1YnZULl0W++/PMUxwOTeOPtP09E0V5tRYoYSc0depcX6libkLFxXMFT2PSzJ
f56p9IphBIEfvwf88FIHoWtqpJmPubiuIISuWT9twQNKS4dVx/toribXDtUu
wwcmt0N/t+VhyemyNJYoDi/uhwl7WE7tgIKvEXO5s3n6P+qVONlJNiYWii1m
7iBZjsHkbSWVT1LFkGx7nuAi8e9KestDNTBEZsmCrsgQpiv/mk5N1f6+YZ2t
XEI0JvWZZQMr0uWO5JRk75J9kVFFa8+K4z6rTxbk/SWE5z3UIApgagdLRlTx
NE8LPN6FCBIfPLeLyF2SqvGFg5HNYorMCr/Qf+Tu0L3WjVngtKY4LMfg4s5t
6wlppEftrCH5F7jbI75fgidXvIEXSsD6MmM6X7xL1YYGCL1B3uQ//Xc+aWC2
s+p9EZwWwVH1R1vyC4ANFbUneivKbnJP1w0bK7YNsYf3yedWSLup74Rv/oyc
16/paflgLkWDSMuTBa+vDAdvrDlOh8tabbo1qknEhPKwfJcVa/F3i9tmPD0g
2CNBzETKSFPp5UcDekMv5ksgzRSiBszXv1dioDnugtDt/CZjr0c46O2BSwnC
Vrxf2fGJo3gPHcGq4bf+xAnzaqetqPCRmBlwgljZnrKQIiM8oLg8Dmu5eoto
Pu09GAMSWtRRdG/qefk4dN1/MgAUyFfjo5hfI1OCLxAVB7CS3AavjFFU2FSf
Eez8vhOgWkO5a6kfzvZIEUujGKdzT7eNpqssUX2L8h2fw8AvzG5fjp8H6Bys
El2dvPrmx/uMuFOkRD8/aDcTpDsPxX7S+sUfD2yeXtyF55V3Db/vK4nvQheP
uwiNMCJ7akkrqAc58FDWq+GK1y5R7EebFKl/TGxzhgyQgATqddnVHmI+TQpY
dNPueX+O13ZfjI07h1zK8wIUFh6hnpdlcaEiYGPLfdJl8Z1cDeB3yM57ToIx
B7vj053k1Z8gs5G2350Em0GonMIONuW5SmIlZSFMI0Fw8R7taHuBZP5guIWv
PbRCzZvbwquJjJbHKm1kFqC6i0TpN4Vm8pb3kn6PSkS9KdPuD0HOuCHo5xYV
VZYpVg+paHTPSj+79f9ODeNUflMqriuKUiB3EX91RYLzhWmE7UufofsS4TKd
p8d6SSmv5UgCfVGeqSf/8GZcKtckTe1seLW2Osx30UoeW1rzDU6o7GT/uPqu
miypvnCiqEWMxUV12VrSiOTlu7QsC3hcvzYreUmi3gdIowLhvtu9norjhuf3
qrF/Y08N485OlHYOZdlcefsf2hQWI2Hu3iEe6tUqV6tmlz4aEyU4OH1XWvIJ
uLiqT3M8UbO3xvhFmTq9b3B8rEvHitp/eBz0S2Ldh54fACK49J4Tl4SKT9GY
c6OP31TNSnLPk2iiDuKZ5u1bIsKlsgnsF2U5nnalWFh9/UDPbeoFiHp2c42n
oLpgErw0y0HBkV7heqiOI9kPwnGHRiP9ofSvH7gxo/3yGGrv20lXWEXm77ME
uLG08fzmb0zCHI08e2yMiU6zCjGYcTfbJ626jmYL3BDTfkZiLZyW+SznQcxU
d/Rx0L7bY9MDKtT14UwMnYm3NT7dKdCJAdPaEyXkFqkZLqYV/l7I2UaoRoBt
MPdw8ZrFHi17zg27/OL6Zb5oCuPXknJRXDBTM8XcNn5dvIrckcUXNE/Lx4Nz
qw1pjJ5WMK0ojW2nOw/BBN1z5scI15vafF9cRUgLwhqKYIIYll0fHY3PBtma
A47elcO8yXH+216gmOcpw/N5Rya0XBJPp6eLoVaE0wgfA7CHd4hITeX2LsiM
jv5TCg/ewIIS7sKRpqekYUGo/aempI98pYz+31wU/eOEC0gmPL+DQmeTvxkJ
hbHn5Ht6o+TMAjSvEWMAT5yF+Miy4y/1ihILcby643pr1lnZpO1IMjDPZ7fo
CX2DflBbi1XEy6jLY7KTQj5Hi5kkow/mrdriMXSsMhb9lMFebwy+7BNAGjtz
JapjrTO8nUQ/cwGdiVW5p1B1FZaT6wlFcpoxcm0xFwVv8yqBF4UpbsCHewPm
bM+gdYDOUbchB4QY01SVUzKH7wm5a/XwcuN0s8h0jNz3L/r+yqS1YUsJJAau
ma2MOnhWbHNLPANAAb3XtVZ652jq8iwdx42VRR9+s2pBpjDRVHzHDeUNgAtr
ZlcsM7+x4/uwfUED1ZhfphzodyldsU6yK21Y1cwuv7IQ98soRpSXtbHBgnfs
PFRRDoIDFswwL3ysscN2vuYvtsz7XlSerPEtpwaZy0ZzR/vQUbm8fPbquxMs
Vsi2LzGKfs5CMucPdwIjFS1raYI8KzFuoP2TTEmXAxah7x6HfJG5u4pAgAbP
HM7QcsSJVr9Xr+gQLmzkJhe+Nk+m8+ZPuVzkxipfjKLC7j6xEqriq0/KR9mV
nD0eGPE6vF0sJJ26BA+7kkJ51dwSEzDVHRUvE01gU3dkNHdVzm5KlCEs3til
TSPj1fADfZESidn0FwhhlT3rLJMDzThl0LYcJP67MTHDIumEN0USDuPp5RpB
FWV42329l9/hnsdIOQPbox6duRFHDWK5ZwCvIsUrrsq3UG5R83RUPWeRJwDP
01lJvS1g4FyITKtPsAFs0jBrekTxGkOq7v/QeYHnBzYacnVNlDKPrJdhFe11
lzaU2qLc9XZFWJSyFHcv+LbCRTHPayYzPeZ82lqScWyJPGgveiwfoOlebe1p
ZyBMwSsRYMoMxyTlxEfuoqPYX/tlUd8xS169ohMnNNiSPFAyqTIVIelbq6oH
WnkmlKm6wzTo8F9CH5i/gQkAP8POke7p6bDxex+Fa+xFBfxBmVXYfMTErdQX
i8+4UPa9cl00oDEUhcDahn9sXoNJGpSz+FlXtYbO466ZxC+PGeBKnWMzjoZF
5HlcQt260B51s0cZ7PslGIDK7HyrQAgzNWrlPmQSrzFEOuLSkYxTLm7uqKGH
RJRsu6VlLyn0ArOx3gj8YebIBRnSdqv1rW4zhUgbMPmqf3FubyameFNbJVRH
yUUFN0eL7tT3X8rFJOChS48urnwTHxrwu/4R+LgCCOy1WXcZCEOWkwa3cN8U
nuWjB26ViOzwRxIb3znL8rs42MON0b0pnplUJayTFD58nhXCI1MNXoe3ncqS
NIm2Pwt5mykAlx4LLNNCKk5KT2f7SDZ5NDbNDoct7pDa0z5nHfAx8KyGjVQz
iRk4+vB/L3ucxRQKA5N2pPuyHwfvfyfyq83BPqsqehcS7SN94MHKYGGL+hS/
baSE7K+i3NA33oGnJUIaX7pOeBghDER4Ster1rGKJQt/2pU1jrTZJUvmWdDg
vDaYp5KHy/EDfyKHV7cU4k8EVEGF7egclM66B5+ogp9LFTtWiHN5GHWiqNlQ
qbyg+W0rXTI2H3QVLjh1MuXkoPYaXbiza5x56CxdSIbro0op+XA1yQ3eMYO6
WSmr3N1eD5KzQPAJ8syhXon06/7+82Vz6WFddrH7MemJLSG+43m8bExb3lWe
bLnbBAp9Yvr+YDrEvHfEoBlLTEKQ2TeQcv7TNHMxu+d1F84jxAlZnwAJki7/
MX5iaF20nd2P+V6k1M9mF5JkT1LDblqG/gLRKtXxaYztXoOqw8Fm2uEr+vSO
xv7zHB7jPj82+/RMOLvyfVl3VXtsd0pDvirXvIJ+N1YI0xroyOne8RrvBL2J
xKCqZWmdNSChcG2GcpVIXNYzALXns1NalAD540e2KNPFTFI8Qy6t7zhFVXA6
rPLpIPCbyN6BrN0sRDEhP30qnSVup5Wcl3ZgB5i5aVXDexbU+XiwEtj1r6Ki
2mYcRfXPeoD0qr78F/JK/RQaoA5d5lk2f6zdYqf0fgCzYInyJL8cf5e8lo6H
M5LipgxmbXI8YaB8grbPCu8IJkAMVsnoyuX8hWQz8ys+vUSi60B/N0HZBFd+
QPCfGB0jsUiMOuYMoL85I7DvxXKG5ppSSqkV3tzNkFciQu6u+QuG6y3Dhwj7
s8W5/Svw0pahSkTJqKUv9xnCD4TEn0LsbKD+rvBn/DCjUxI6UXE8EmGqbe3F
zvOUsEyyR+orr8MtfA5sEaHAd53JersA8490arEkEzcX1qON70chjAecCLwY
gUk4nSNtYex0dbmqa/5dNoo6pVF+zZyxEfRr5GHs979aLi7MXSLA5RWHMlin
Uy1z+tcw99FiiMTpOCIdjljtJ0RUtcgGWfECedJCqdFVisxlNM7VSlOF+m4E
oFy2GUl2xL13ODL1iFWkmlgNr8g5aKz4+aiyxok/y+pwUailm7YQg8XjbNCU
hc6iHs0bpMjws6V8qrJOOV4fuyHL/uCjPwWigobfrAZJ5lLRlfhuVgpX+S3Y
l/H3QhcrBnPtzDkxOHVVTFckNRlDVryzE03Es8uva3UhcJURIu7WKP4n1Euy
mtmYUaES2ElJheHxPi8gc+OOqvEsDkD2QVNF5mzODEEVIYu/KYGHnBk+19iW
5nYk1wiB6+WEUSiKlyXTxbWZjbYMFEh67nG6iZ0IXllbPKBctwZbFbNZ1BM/
vYHIPc+QsoCeRiNsy5pdIkCr/a6qdpYC4Y/4/Fk9NFEHbHElaFjA6L9KqEwO
+ud1/srIxZSFsYo52a+7FgnGL4BgqdwDKK2tDwbJnR/4d/mX/c3QMctU3gMr
ghJQk48WzPVpHqynDNQe/UzngDVxeDQvG77mYqTucSOhyGtpTs2jM4RVXuaF
OMf4/ov83W53eXFNFRl5Z4a3TVWJSSLJXUbsVSm52ymxvheYPtoFpTJfAZeb
8DzS4J1LrAk0JiBb3HM2dhXx2K8Ps/0mRceHhld+V+GDz8x6Rm2lqiC89FKB
0Dcd51M/8O1swOX31uZ8UwgXzm/QrGS8z3XWFUPG1uAfmCr0Lz+/VoR+jV/c
7/abS9EDi/DeHiA1Em5+CC6St6+SHtxETin/M0jCf7JQzpwNJ9pb+UO+JBCD
Sb/tePsC3anQCvQuJn/8MbCpDFmTYzQT75OwF+GHaS9hWAaA0uOzqINKG9YV
pLM/WPHtdxqrO/suwAwr34UeFbjInXqNu3ydD3Cm7tvL+VjVLveRd7vYm5DT
H8m0cUV2uufpBphJoZ0z6qDZkLBPDyZ1RUDwlmmcD5+iPpjIPM75P05SBTnQ
8n6nZBzStg5yHsUNW0adOYHThXbhQWmd9DOP9N4WY36nBY0UQcMMCCW7SL8k
jqbfFCWoepUPIYtEdhIpo/8eCxVWcJtn/eqWx1IoZ73LIIS/3hRYqR/BG6Wk
ACbq3oPzKc00rpvyf1DDUDrM804zpChmy8hK46GzuVenjEBfUKg+3LZJMBp4
S90qNAG73LiyzIE1ZvHxgDUT1ANFC3tRdAoRJXjCLcTx3WylCNSDGfwQ4bI5
EfdZmR5GHRoTEKboeQLIi3ElcuIuS8oCVqQfdZIaFkDKL7YmZxAeOi3Ecz82
NT07bTjjTo+owij4bcrtzs7xHUAmW7pWd02XOBX1YWoIG/GJZU8yfzNdRjOr
5F0UJCA0deOE7Vmw3pTUS0bGjA5f9L3KGOtGf+CMXZxODH3DPdkD39Vxo0DH
O9iaGuMfUR2BXUadI5aVaJCSFIsMujlnJ9TY8U/eYw1hsMoVI5f4Mzk+kQ7X
MgQS7Eq4jdKA32t+HC6Bk+vigT4utqaNqA9EVGJGcLieJWrzyuJHdh2rM7dR
DNxxu+2KcPRU68cQG2pwmHdxlmx24Uct5AjTOSL8H/iiGbwL3FYNv+083YUL
VOcUBW6Ra4BRWK6L6anKgOTNgNcEbLJCf2kZewDGgFl4qZoZCcgjTX29tNFf
h6t7nRqcFWQdlhI6y0rJoHjLjQTWCkI5n75ke2Td6GPZBxQUBLX92+/qRcpw
MOf4L/1xPqu1p3AFm5k3OfawurfvTpyrbPbwpuyDlIb0C5Lqhzvxy737unNv
D3BgXTnv0LbKnvZeOPUbBT6rddo8cjSIwvN1ZFFhe6cc5SmcGg/PvyaKG5vA
b0fvhQQTbC73DehnnQHtrOoN98133CkSnB8itqcQuk6U6hoG2G8NzFHemS28
za0J0+R+XQr5mv4ri8TYQv7vXjnqGozgGQ0cy7XIsikgCd5dt/zRO6Vm3ywV
b/vAWmDEjjl38hkyDzBABXXCb93MnU0XimhGWn/20NSQZQgtIe9wxBvUifpw
vl+8sdB5kk2+ZFe+DDSOpB9dC5NSA1dnFVojTltczZNZOnvk0BMsFdk2qiPh
6wKxsQnfvc1xPyn8qU27vL8lpUmq8VfTnK4KDYcxMaST78DFb3PyNq8/8NN9
67qN3zJANVWydVUlWZUvcbVhEnC1ndMkFeaeZ/ufggO7WXOQ5DZs9striyN9
jF0Wa7ke4By+MmDpS+EFOITgLh8f4ox/mBy7/A8jAkDtbeRff3jZZh6mLdbW
HJ840RpPq8uQMcSjb6+YTyr69CqU5jCv0xxPRXkcZ95b4WQOtNr+hbjMlm3q
m/10+12T5O2hRpXCuAynkOZ+SBPE81Q0SZj6M6Sg4CQEdcVlto2sytQyGcwQ
ZwDcF5xBzB9atlU7L2ixup+lq84EzWDqADc3F1K/UWiTkAo3xh8Pf5HtGJOT
0ChA0Bf7MmxYD7WdmA/PWDHgEXCzcuVO6i9Vsl9styKKCE/kHCNRbBnC2CIr
+Dv5j3FJHNCTqUnZ+dE9b3oWmvBhbsmy5495/A/vhIecDBmrsg0pX/+BwWtt
vaJOgVnoQ8U0L6PeMNhF9Y+89iv26MdJQnzvsfY7qMfNPpbND9w+sle56eoY
yiz20+OXvTvxEYEeoqL0u0wTrFmNeXU+4DXqU6IcB8uYm4E/sf2xDXiMNpQv
POmefVq9/pOGTmzrjawUeyZjTVOr3ZqQjQLJEoOAYb2onvDlP6/a4ebNNOBk
6Pluj9p7LgGL3HAFCuaz2m3SEP+0WsTeNQRzCZ3dq1O6viStEJ8dwFDZJV8/
DaxsFpcagLgiFB9b4JPgXDU3qLfVoSaU4Z4Qw4hxqPYeyp0JNmHu/1Zwx/wm
XaBKvJ5NW6+Gb5AakUR22ADgU/OEVrSS1hZGcyQgMFOtRwpy1xFc/6d4Iran
5X7n+73R9Z2oc1CW9wVDzIBY8dt/UguYZXrC1lW7Q9U4NeFnlRmmEWZ43nl5
TBnrCOQ6IegtpBGydqyX9CY5Gyk7kJwkOQByK2+LQMehxGZkSIk3U6ieYf47
tnL7sFUXjc01CbEWf6k65G3cAOv5RQe9AAyGRiu1q70tRvCGvA4AKOWWdMhm
xrx8uGl7spUQZOLilm9H135z6ytafc9wiDji01YI9gYt4hgYxRRfs8/E+knn
hmmBYIhoy9OXIm8QYq2b8+PxWryDMJtjiPmahOdO8OIGuhud+hscHkv07uLl
k8k4zYii3+1StZ/OYcMoCMjOuSuxb3jgHLUtMERvOeTgpMBN5CBUXDe6Y1FC
zFQBOa+je0ylvnypGrRCe8zlyhRVom4EBm6l7QgOaIKHv6QQA89VhNJ2m4h9
c5UF6uuGknHzsd/S8GZJgpwoFh+QYEuhOCCkpsvgPoRvaL21XrAabJfntDNz
VMoHGWbjZco7PHuBvQtoIAZf/Mfka8f40i2DcP2reLxgYQ9eEtxM00hTd+vV
hOhiJMAo58HXq+pOZSxiEgkLK6ZuBjwkVqYJjcKPv0lMUo0310Hoae7/gDCr
qUsUc0QLXqS3syScYiF6G3wyPAod2+8quLcapTaReQIOKOCTgBkuYCYAeLrK
/BK3A65WM/oBkb2NOm5elBqkHYmQ1j1Tl92nnNt7zpFVyuDEIcoogiofruXm
oZB9XXed3Z6INW2u4syay2vFw1582hzR2N7UVhkFXQUSBQgNblaRZL91uecl
0wVxfXNwUsvfBl/pct9qdPvIE8msywti/6Ypuop3MhpSd6RXEm8w8fFF9oOl
OXFfSbwB0hrEfDJI2rYPJewUQ2ZUWlWEzReZQk+jlgHyLw9JIXZlf2nkjl8c
9wz/gKrcbKFpogM0ZTtGmLHxEnLza0HrcO7RWOigLLqmLn++iOy13i97d0Sv
bp5UN6X59jJ949bkm6JShYXiGsB3kT6Q4kus1Pk+BJaEogcRBaM6v219zkVx
TzNFkJycQv4xfcbuP/fI0aTa5eCjSB8Y85QMO/3TPTKV4HHDJaC81OjVan31
jU7XrhL6sLNQ5oEKtG7vI2dT9Ig+QQ9gNve7bym31+BsZj/jKCCo88I8Fn9+
w3l00b4rVFMqhZNOiGwppiX84ppgc9SbbGHGa+6gmZOrrhlh+vJPF8oQ6989
bZbTTGNtgOdDFAVuNSOU/JZ8pS4vJN8sUgnwWgupGHBwuq6QYjF56Sd8Kczj
9Z8cj3g7R3wJ6TrVBIuT+Ia0boMdIOWD80xrYQJjchdZy0K+sSLsQplDP7oj
FAqU5ggncQg0dowuopuz0X3isCdNm996GdoGRmSAEE910J8myZ7wCeCREOWA
PtjLeb3L4eUIuC6VCBrRReAllMy27i8KIllzxTK2OuhIo1+EksvoVxG6ntT/
mY5BVL8fjysEfmuDzMu5/duCz0fq9K9jDDjLSpJZcq/jPtivD83Fqf/AoqaJ
Rgw8tCDbKxBJZDXPHpkXjCTIT2sMjR24iJeIPrBOjfAcyhanJhsXY0HD6BD2
pFLHx62lpguwBaflJ55lZKbAUgUdo6dPl7DHispPcGaeVxB4LfyxMj18Z5GA
vyOQxsutZNX/fdkZf9TQqNVWGzgZzb2SsX0OaYZFBQ2YkJ6tSITivjqCNZ5p
2oWxwGtV6asu6ZZVYYAWosEJZ+kxwn/Ega/LZpzgRRZCjrDw2dWhNz9BgudT
Yt1N5anDNXUzIw2JBb+q1kwJ0uIllsPFvWwAZQu/HP62cPR0nccc+NpbC8y+
NQXKVlyym7SsKL9Ms6LUGASJ/FtdwB3lnNmbw2wULJBNnxVbBWyK8zuexQmQ
cvvfA4UnUqpq1dPqF7rT5kXDxhx2FtaXQtGY7QJCYMOKHakMINaUIZrzvfCv
CN1DXWjErN1pPgltZkS3xtpwyClhzN07SxDMux8IuX1Z0bQLs7nLCCJFBpnt
l0sFMyBXsKxuXCQVisTDf96KgbEBOpirNwUHOYch33Aj7vUgcbDS0cqQ/JpX
b91VeMHrSm7oP+7jOZChC1wwigsaBcqmzPQ3X2CEMEblqyfOVa5BQLDcG+0/
x/5FWSrHMm5OY0x/Dy3b9vQp84/W18VDo/uvHSMyUspymMx5R9Nv3mA8qwc9
7D+qti0MNOJ50p8vm5btWcN82YPUSQ1JK1+mfxPBu3TB1xXSA8xz6q5jcmm0
lFLK9tKb/zaARt2m6ydHipnJLLqfydTd2sR0+P7mvLvweCPpH8j3iib1hYLV
y/P+tuJBiX817pIQ5eGjjw3crLpW11lP2qNmRZG6BoKNlEdPm2dnGox7BRI1
/ALC8T1XUbb+8Rtso50Wc0EXqcOye3rg3BJkI8JTQCk/5+fbOVxZFNdLqw63
bS07l86My9DGALLTfyog74MF697mc7pPgzn63l3157Slxwt8WgrWl8oNN334
Pxb75X/EgMX1Zp7JSClSq3sRcEDyhGfXxYt/FUdxa8Qa+ZgYMVTZISWZ6bKd
LeMqOlS3ub9rZdMiP4JHHv89S7Vhil4TOrgORR/GvR9gROultZeCGcRsBJ09
ncv2JxT0G92qcqPhZmD6IJaO4Nf9cy4M2qvnNlKoE4O3T+t86KK8BX2RcSZx
RJjoSwDn+HxUiQubPfJyhMrlHig8s2DRnsgYnufIf3hQG/6S4DmA2ftRwEMl
7PvvtsuBazKhZ9psXU1+HftdMAS1wH4CexbGD6uTbrYpzCu9sfI7VmcoMoCN
aCFndwWVZpGGSvGHibjwIIEbj7cjBzdVNoIJdUJR5Ef5EEC+ySWkrupmklBE
Bm3ybjLRRpl6hgwS+ysM8xlUfMHdqFCM1OYBK6lthYps7eaZ+vfon85nir7W
i1eu0sTowNv5kS44rqmt+WupXqWfdXcLqEvJOv3xIdEce+A1mXdMCpjjn9e5
1ibFvtPMiUFG4AhhQ1rS73kCwAiamolUBE/epTrKjluuV7Zz6PXNprvHcyTd
K7EPUSwortZI/scDAoeH+cSmDGXnC5giq+IJyt6qgQuOlX9ihgTe7Yw2l9Jb
nj9sUEaYsgcdD1WiQ1a+NvXo8r9ztKvGM2ONBHxo20tgngzvEzvhD98p7dTi
fKLN3RbwHLII+N1Sby7x/NlquwXDmclIKBQUGMKCS59ZEEo+SUO8S4qfVgu9
cdJ1Hu//KPdNyBWgsj0qoT8n7psoY5+lIu78R9Qtndrw9p/h9b27xKJaF1r2
ijU69OJFVUjEpqD1i+Bmd0Ejo06Smj6Nbbrp3fMu7OtSVIaKoNm0DjeFv+ui
peoJcJKkGSW7+YssnyqpgWN6+EkBZItgxogegASHJGsYBA+rkMhRmQRShrAH
lD7DOoJUas8va8c04xVg3KWDVMNr3ooNtSXHb+a2qfE7AATe6ZtKfQDJKHjA
hAK4qOr/uUzGZtHXtzAwAUufKhNtcV3gQnM0aT628PNUl7lNLWJfiq7XhrRt
Gjm85BIVEm1E+Ljym71NqYKvu/DI3zC5kLOfUZkU10KdNbuIDG870lwuMLp6
CHAYaQkV7PS2co/UP7oyLdnhbxk4V7i4iLRtkAAeXfaJKbEeIWT5U79KnSNx
EKmlC/H2La2e02lECzpsL0iPTTfmMoPC2yx2k/HaysKbcmgbSk3bWiLcNieK
FbGRymaJ2+UtLUcycqtzvBK3+ZCMaID1azo3H9EeJxdrnuTHezCyvF1xslBR
PQGsc3YnpAO+1hsoRZ3cGj1CsjDG6TqVCMkSQoNpXITeJ0mDPMpXTPPf0i2R
RypTfyfHh7WCFC7OoTua5DDXhJ432V6SfdBu4E+9VYTVs3U5/l7F4cp1plQJ
RR5hJ7Ddy/9dA7RqOwN6E37m81Fau76PZ1EI8+KoKDjF3F9GsbHZefcepQ5U
HKxpuRYeq6h2rbyKpH+IwGzQ4SMlVU8RiLu1oHlrHNuKzpvEeERjOCiRqOiB
QIv3BkU8d+rRClDr3MTpPx9auqrSJwl3PvWdym26dcTwu5YDj0ZKNcKcrGWv
b93cx3WQkzjrfXa8d8fQ/QBj9ZCulszR3ETQsscYQ8B6adNSWNl2JXT81s29
7SC279w+IuU1S4DMgBBPYv11RBgWufz7TqNmV10wnitrjuKspdCnWta/o/od
Nfv6BFW4NQgkT8Ecwh6pCDN4rpR9QD178P/HJZczhg9FzBRSeOe2bsk0BUk9
poENARqZPzMTwWDGer5gdPEDo3jUOiosOXJmZE5D3zA6PAG0Rmp2XOeFqqHP
Hp6giTD3pBNTi5kofmSEvhF0tQqHmzZMgZeG023h2FPIqRaPsUHyuIj77oq5
lcVq1UgRe9gnTLoGdKNTRRW0MGBB/wnVYhGhc3W2Ubq4hv+HfrtDpfmWdHX3
LSzc5qcCgTJ1aoPgiquNjLMI9lQuMDmqh5pNhHLvFOFT4k9mh4jpdKK/ifI/
TQbdVdUXonhwJ/a7PFu1A+BI3foGXmKteLeuoc0gktQeAqGhFH76pv2vCZzU
dbVMvdD9n8lfSiCZfgZWVIslTqWSP4h6oTH9RrEyWcbPBfmEBAtEIqrgG56p
YMc81fJNwrzatBy2eQck9lkGMsULtdl8GkjlUwIsAeF/l07fjZFZBA6X/7qr
V2Lzm1K/dRCqLgD8wnJKG2kqDDcOtzwE/dHdZUBaoXCgdizFokqugt2kHlLQ
NltmwgN9r5mY2gWifzUXL6qSHmxHBprtk0jbP3Efmi2Sf8MWU0u7a7p6JzPd
dSljfKZ/GOCT+0iqXus30I6XZ7KSB2VQuJOak9cfgulYMOWL3bKgR2rLsS45
+iIuTRcgAIqasuzhlWB6r3nmTq/CZG69pYxtTFhl9tD3PqpQ+L/YyNBRPsrK
3GzsYl9w59tr4w0R2R02PoQcD+/GBPL98w6E1nWxVe5I07dxaAP/h84hD/I4
suHlhbKAVNBM9w8lmZgf6vy85VPTQMNAJrXZQrS82kNRtw6k8PM+RvypN1dX
l6kOPjzNn98fcQ6s/F+nBjD7fPWVIKP2/11SK20TrUYuaUFVtJ19O0xInLSS
P/E1sV+m8isNBgNCWtywubApVALaHxIXOTV4vGNJk3qh7Mh4Z2+Vv7b0CRqN
jw8uYpVY8MHxnaaR1y6Fbq3J7YQ79ZHTstKUzEWnnw2DEfYUwvVgRGpLmvSF
WgP4E7ba1F03L8j9n5/un5ofzTfpZKifop5Zmw8ay6npKP+HPxXsqEd6Vlth
VdeQsPERrWOTIq9IJ2VDImY9dgs+DJwcoCxfgoeJJYo5vq9dDvM9JM9QYqId
RRj8oGKeuWIrhWk/dyJu5k48EGgLkmgPf4yTURn36sdXMvuGrOKxGUiO5aqR
sFVMgFmHhKRSuSLR/lZfu9Bch3kdreJ5zvbKIvkIUKdvLNgSQlVqfsnqhN95
NoOzm9aztzHm9zPWwlM34WhlFN259N7TI2zfgLwI2AASMIwclWO6WtGlMjSe
ES0jgx2ELchTXLDQ6V4v3hXrqkJPKQyaQ6oz3jxCJFWCRKi/1G4VPXZ2gAGI
3rrdn5o4Rqd+GwPKoynALwvJ0EWSf1qLdxunsExORITw7hdFmHrZlxOCEYmK
DsoM75w6S16DdgS+AAlgLtW5/AnKp5LXrVHKB/OdI0VsWjpj69qGiYdiRxYT
QJj/OE64mVC6u+VnkbFAB4lH3Shzt8EA3/e1rkkJObwdMz78a93W6Hd2kTE2
3MrkrJ44wn0eEz0Vq/4Cd8VAp/8ErJjm/TlaOwupNf2bIU3LIcpiHHr12qtv
bTOi6GvlDqKw2HpgfgzDHG3SEzQU4r/MOHFNs0wSNyUZlsQeLuK+C3e9rUxA
lNyayevSSwZNuCWsZJhdk/QxrsAyO8aUJB9qX5c3GCoDcOZFZdUnFH4cFp+B
2mIUFkL/nZVLBnvioypjUfzGBLdiuU54Fvz1ZrVJxfv5Ez57I2OhWQNyRd7l
0h3A0N5adgVF2HGcFUf4Ywr60AGgLkS/vB2ti6si9Ow/WVH8wf5ruSUCr/M7
JQ5Fe0MDr5lzZxKB7kh6GsHOX098ZZf+HqEf26Mr6PK3GBtUcgiOVstHwuMu
A48mDHlGqY1LsIbFNlbFVoF9AwZnvCRFe9lKC9sFiSvXgjxM5p3P9SGKRaI4
ocMhe4Jm/Hy2kEtjFUUQiBCZAtcKe2nh9VLydFElKLMzEW94/VRkF77qQqLX
vNApgydFRGbRSPFhawMxu1sOIKfQAaLu7O6VyoSzvXE9z701EfDQ9PIW5MMq
6JXhwCOoMkVXPcYMA+ih07v7mHd8ZE6UnD9VBFCnJsBypaTllVoBL1SvGIJJ
bIRffkvbCTYdILLWvsWHZIs2ilBT3NBXpMlxNJk07H4cF56A2PJNosvkus8H
D0B4XDzjdCIlOhFUrpUdlrDn/N6qPrZZLlXwceJXWaB7Ko+lDSCKgoGF5dYv
7qcWG47r4EF5UZ170+v2BpTvCqbOoEDvawQXwJlfgFOP13E7s5gDQwVGadbG
BLjwtbeNZ5+sgl7EGRGl4A1r2L1qfv4wujbIv+SDWkihMI2Q6TWm0vts05Us
g3GXs23nHg4jxFD78OKcDTW/a7wkmnC9XEnioqf4RVRKbtutQ1A51yupl6Bf
AVC3ZObueKcZtTTpP55yg/epif/PEDCijaW1jp0ACmVVTai1wC6jinZpwqqI
+VjpPH3B3gvVJlr43mluU9Ry2Sb8IVX7bLys5Ns2aTyVz3DxvSscfpxZqUvY
+6PtCdNuwN6lfMrK9pp9bSujEDv1KQ4RXBahX/YKJr0gN4C6zDvtJX02O3/F
WwHoZMs8XZ0MyiFSUhetPR4F0vWFKyji5PYiJYvaow6Ng4AzgGg/lftBlcSS
myjYuMSRM4fd1uQyARMIKbaIHxV6zcwwN+VLrOioZuFqSKop3cXHbi7fLMXY
jzLfd38vSsbQvY93yWBJb5c9a/IlFkLnG9VPvaHSFSOieGxZauPH7HlhdnHj
ZbvViKAGhWypBFg6ot59hdj3Q1RROeqffcubfBFJ1Vla4qeNRBuzSir3U0eY
Qy/0GyKglggE+MH0tXfgh4/c+/kRYYH5qtnjjL/ap2EobwGyWIVIibH47QmD
3vCBLOhAlAp3UU9ceehVYkHOs1TxY027L/yc5TMzFLqbZaio1iKg+5AFIx+L
EVMvcnEmFtPcrdWDb+psHYfuFpxtYO0TDWT86vtdxE8BF0sG4jjWPFXL+ZO8
DfPnZ3sVWH08DJ1CXueNxAIkifmGmYWlDWw1TWq9p6bUKAzbkTwWOlBPBKjE
s2klP4ZRs4++tTS29c4WIvjjm175I1tkJyLtgwCd0MF5xHBVwe3F0z2N5tdc
WJ4C9tbGugt0U8pP7Vrj4bgxXT+EO4frdhDXqg4UDXHSfV13J5NPz8k1TT4g
EPnNyrIr4ItTl/7vaPsnoRzZ+efDjgTNqymElA9JDwS00SaUolibAdrRXd2K
Ho5kyq2visybRDWdXvnJdWgMWZ8GAc1dLZbtYsugeHeO7XID1ZkdufkFvvSM
TlZqVBRZH8FiMqKgCWqCNfQsbMmrzDiu+9ToxMom2dfAbnur6Vi/60MWi98S
Fhz1l7atI0x9J8Cyz9yRdf+LebKK9GuS8OBF+F7WjYkbeI2or3LdIheY4vI+
XAnYPMeX9ZTIQOsysZOwLS2jgGqLF1xKBKdVTfcJTmoqpYbgC3TuLDjCPrkF
quiYQAQR1iIN2+N6s4dgxS9sMC0b1Egx4RUAHVYf28GlmgVtIpc6SSMpF1qv
QVDn15NCftNNjOnuwEzPdHiiy/yKoBcU4F6ciGJJKcPLK5ele6upxv7QFfeM
YfMvprIsWBmJS2TteCFjViTgY7KPyHUT+1f5+D7mtt9fLvfonmCZH8MnpLMf
aevcEu7dFSyCX6rofSRfW1xXjwafclvqSEIHMEnmGQ86/P86km9lLDd26XXB
+B+WVjiKYzt2b9mVUBY+XwHIeNtuh+lNlwjvf7gBjSqKb5YSdeNfZlh+FxT1
y1+5oCvgdrherKAPvfoDyURsB6VvKVEDhQVxbJ9IacD0vWKCvj+GhbKq/HF0
EEDGafE0NboVT0wcuv9s/zcSq2V2oTQnpjzZuEBhlV6PeK+kUDguBlvK4guh
zv25m9uzuLMNsGB1ljoqMX9MyKCpS94LGYewWZtVrEqNcgynO04FIVxkFudu
d7ZjtshgrS2lHjfOawvpPFVqgYYTK37WdYoCK4AzlGV0bcXUYkS6Ja3BDKDl
y9MRKt9Td94H0hiCCW/WBU19w8b0QycshgVvGXvE64r7En7oLf3rlt4hq0cH
tJBr7gMkYcfsRvGLFDBOcLMiJzjdE7/EiYf9YLcsMIN0G8afXdCFn/s11zKY
3VLJnpiKIHGPuuShE5wNti2L8DKhTAiOXlsVbAgjZsDaQi0K3k0G1qbz5hLk
7YoVx6v3K6xwsOK7FlQDLilHD0lnqQ/f4S2n+j+XOTCRnXAOZH237LG0xYvi
1Z4L6iG5lGDRsosxX0DprOIKJBsFgNbNQIq13p53NC/T7/Gy6CQNXpsnCrR6
8Nfeg/AIqGu8AIiG49vendlXxbW933/u6OhOu/tIFnkPu2d2uZv0+CdNmo0l
id5gm6X5DAT5xKy8hXd7P61Ibcw0Ds5YbM/F97HO1dn4968FWqyK32DOFxZZ
z4FmpYH+IrQFjkRis05tH5iOU6mPPObOMT6tHf9BTiMGa3UYbbglT9HWGM+C
ax3nsgi4TGLJgdHgC4GgOEuRSrw5b8XGVE+cfvqWCiqbJMr9IXnoOoDqRKKZ
CxLxSAbcZ+EbrQ+3SxGvilOvga5I3Wjwg16ZRucH3btgJPKJqedp8DUUOTH+
jcc7I9y+6QL/LyALr9exocAfURrZb78UBY4USXD6nTOxw8ZzxZADDFbXUd22
5l+J3KAywm38wVJwnQ/iaf82jSBMy4ChkbIwDZDQbkIJBg1c6iqt0L7z8C5Q
lYmqOR8SrLDERAyGsu2tXk1vuzJygosHidv7mnhJC8q1GUAC4d+sCQ1yqoi0
jGgW0c4RrtlCbzlz7IGsqZvV6wvE0JEcH7kxndDow+UhAR8PlO24gAT/01H7
xhbhQuCzE+oaBnahFKLifOcABG2Ss57llTjbVRDKwXOAzceIrjteHs//iiKF
kJm8kv8SlrHym64hacXco0eDWJ3oIykMi9e675aIuP/t/seuhwxlIDFs9mqL
X8RmAGi5oHM65oYsQQZBIn+GcyZU/q+NeHi5laY8WUPDMytK6T/gPjI7Zc0j
VHkiyIZC28y8kyfXMoHfOobAwWUiV9V6XyffYab42GkSZ/jleRB0T4jKr3db
bDg6NxIaTc4qfvUDc9vgD3H9517T73NSMliKH3cqNKyduJ9feUfmXStnM1Ix
WbSa8BWSQCcrpRWCUNAGHB8Um4gqDNcUnkC88rO5K1XfDKsXEE+bvDWxkt3a
GF3222C0yBzSRujoejMsxbetj/Sa/3zPKc/srzeevMru/m0fGt/z1YIFpMk3
3wAVIYzHeohF1hemd6w1u1VICfSmhthDwKhESLe3R9mocCcIiW1pMcsXm7Qt
ktlDy6gpAUzkOIDJTtiXc+PRd58XYGMVXfGAf2QZMDSv+wAWM8uVys9UyVSY
dWDQKft+7Bd3A7B5rjG3f6GhUSA3+KaTorr5xmujPwBBsX+Ucv3MgcqhlSKI
GMHTAFLXLBudP+n1okOWpy4m1XQRZKxi+ayMuNb2xXwJ5EgxUs96GQ3PVbdo
bGv2QgCedKzM2m8X6k2N0hmibnwdMRlQ3yTBrsvzjeGC+X5GlcrU4NOPZUdj
Vk/YCc1W9hAThkBvnnGcyUd/r+/km+wHi6IxC2XbRpeI5kmNXXP75Yq6JaOB
C96Fbil5yqTu8/SZoyFnxfS7ubkY61dGmR8PkZrhy4gLLyvPnCU9JIXQLyWo
KibDZKHLz+eXiz0rUblwN0sM6l1liVYDqxyp8BJ9AdPNl7eJXT00DKodkM/F
VYDboPbmQYcB7dPOGJqHxbnsuUgYWuaGoj1qWiVvoxnKgahE//55Gbxe+S8b
nAomHHD/WLT3Co6/R87sLEDlHU34JaG6z5OluPkm9LZkR7wYG5AN7hDx2q6u
TZd2kGI3VM/w5vs4zi5Zr8KbPttvhSW7HK7jKdTNIBLAXDIZ/Fu8IDSBnKXD
7W64dCphzHj7tGorxQl5xRxuTXwucBzgURnH9oalzTXEa6BLO2+UsznCZ48K
0QtQ5Gh8LBd6m2KnEZVK+mBCrqdbIV4H8xsbeHfEn3bOOH27I4jIxHknt2dD
yXPS/SPHxWwWPurAp2TyrJmIMqplUZX1sYiVGBXwd9isRuDvr8lgZobHFoHj
QAoBmBUEbbTZq4XVYcRXgGxnTXgqP+sqsC+2m29BC4yC3Hr+Ipxd3whjaIc2
gqeKXIXRGUbZKiI42ArEdm6YSH3g5wjr5qFsJ7zhSsXg5Lz3ub4IxDua8Gje
SjsOSBfJO4Yt8AW7CZMPYMz1h5nLvTTNheuiXvcqcigiib6piaeKNAPmzUxD
xOOEAc0YdfbZrHWVrQQ2I1WscD2zk21WRS/Z7304jgo9kHn2n/ZCAvCaHzz2
VtLvh3QyNXLU/YxAYwyHKJQdB8c7+ZbQbcAQHwXHMhRvjo0YwOgwHMNBXTDU
73PUXJLxZSZTy+r27LhyEgd72dStsTadqP6EezS0r5zogDlUuWlI8UDteie1
tqeP7m8J029r1KrnTzkK9zxsoGzxV0xA40hKDfY+gCXJWdpkjLG+Egv+RlgQ
QhOb23QPBydiPhGD7tXMtVbbMbtcY2x7NPaltZTx73JQ2GqR/W+nqJKYkBlJ
8G2amGjvXE8hP0xx9GBs9Qd9n4saaXY4klyPbGmYzDaedCu6xFguEfNbGOwD
E8n7pSd2xkbu5m3AY6Wva3bzEx4+Y9r6cBSd3hDEdrgYu/PgWbs5bcs2onpN
NAkhQQosssNfqwOBz/lIfoIZ8VB77eoxvLEdpvLmW+S94NeRmVox8/65aVSv
nJMG79nEzZn8ytIEQKxEWw0yzpKcpR2jom3+/Ux5qjN4kuQiPVBn549yhLx1
C/XNEdCG6cp4LToDWgwA6hhqfOUJPZ3rGrzipdKB451MRihRhTTs/OJYrpb4
hzdnSbcLLQhEsQ67E1NlGsnlnq41+TZm646oVrfNaboOUiFgRJfFoUNSJKgG
sPMpNnUA4gN6+DCR9enG3y4tjIww3CdokVV4Ye0mSi9FW1t3zam9itpueVgr
mbSxjIIcmoCIME3hMsBTD+UEDF+ENRy2ZBH4eVoe4OKR8AGPsVWoGZOcFzwA
KNoo0tjeMkXqPjizfIkNmH8mbBg/byppGN2s1L1LRx4AED101HT01uLWaP7t
KaFUmUgA5LKXMauFmficWQfwGEiIM/ZiobBjPNJo7dj06ff+E1Xh7qrNCrre
v1HWPHWuWRLqDDz8B0fY7fyLp7SWbMDCyZfxlTACaApiDK+RJ52U8yt+Hik7
AvwFCMM5s1aeHCwu2fzOw66R0r3FLrnsUtcQo2ijwTE04k5Ao8CW9gSvKXbO
btR6jZ6TBHbuFygZYxgkhkZhVz9NWdJtPORJQ5PFyorvMp5XQq9824huiq/8
eLooCT+pQwQA5gs/TKRg7CsGR1DBtLvu6XIJII2zMh/JIxjBXnEua7nJsD4n
JHzAFg1X4kA144XKYF3+ExHOHlYmdoaMvN4I2QveEyTueckjK0jBr7RuLsxc
eN06jcaRuqNQ814YqoPMJIzTPYwH8X29hpVnl3CH8YEbEN1uYxGc4QmLUgu3
hhj90Mg+Jg5zkyi25MlGoVv4bxed6Re7yzQai72oKIeFNF1yE+0bhDBPLEe6
q+O0VwCmfkHOsZeNgVsx7/rT2M40EDd3deujtsyJ0y8xtvEM9gyajgJEERk6
qYUFRZxksBJ3aEP7EI6mPhLWsYWFGJY6ufGW23n2dYIdhjpSkG4pVQAtfJvl
pF11yAWT+Uo/8ONxPfGDDAePFVmgjZY78RDasMzYvuBLoZebPJPToHwmLex4
eQJYQ3oFtAGdBxiMBArU9z2kACfXrJaReDVg6JNDmz0nlN/ZTaIf+HnKz+AF
ejUfZY4jdi4idp04ZgyeJuxNSIVXj92WhBHDrV3G0ZhGuAJsn3m2BpAQ7bhV
afbRv/w4xli/KWj0SAd3R8+P3SdpwftG9EfM8JhVikv3jQAs6eFJgMWCOlLS
BgmDzDgzpGSZFfvaAjWMnm8VKhCTXpfuoQ2x6o03qzVuKoy/HjanqmihRUyX
bv9UttM/54Ae0ImgbMe8/piQa3v5U2gu/1tTfobH7hc36V2PTPvo/mvYIyFH
ST3n64LsjvQ8t1lph6t2cd7FATzyEde3gi70AJSWvS0mbrILNBNmemLbMLeE
xwYFUe6t1DrTqXIj9kzyGoiNxkCl+AwIDsvPaY9F39EVLl+Sf4P+iKhz/ii+
qIqVgTNLaT1FJ0Bn7e6lQ6ZU4wTdwtPiiOzV+WVzgemLOiUztt9Mot3vFwU/
eQbkEQ5Ow+HboHItROzolt/VElQGRrskbqD8A+XWw3z58ZmulhXILwAK3ovI
AjGejtKYEN0tfZPyJoyXIcRwwj3bucp1rdcKjDf2YQOePviakfmmTa9C5i8f
dfLQneOXKP6JXOQ1Ekp0OXwG2e4AZITwB7gi+9D5xaqsWZ0p9pRyvIQhzdaP
r2c36FMLJgCfpqJJedj8s/ZAWlgkYVgpN1i7674JveHBMWp6354YV1Zo+BVO
MEQyyElmJRVhq4xwbwRQQTPDU3WeAema95heedf0nIGZ85tBuBMc/4EcvNax
WxwWcaSAcz1DfEV8N0+DRle1kXhfH0EheZOoY5kqDvZlQW/CaREMFcQA98gX
HbkBZ6wH+o+FWXQ4Hfm6eZCqonQ1paLKupzDeaL2na58KU7LyKR8djrKSdIJ
IiP5upWjjLrL6uKu0/siTVsHxsrgdZuAaUDq7CEDZq3CeiITi0t3cvEx0m1k
lrAuYojaCOGe4zHxlKB6e22DrFbsgJkMdgmMd96bbfvxow46p1ZJYqvCC7ZN
5+KlqqL/aitMjTyhZzYZXa0s5GyjoGWLIisJwn7mnH/1ZiVhzIGGP59J0DWz
AFMy1bjc7MGTiEXdVAFqDf9Ryfo0cdODAv0LDMhuk0CreNHpCk0OEtdCQdsD
OpwiL+Pd4r63g48sHsQHsME2uhLuzrqNf7vh5rLqQdT9nROQ98kwgKsljD6z
t3GYwO91Kiek62p5blgp2MqvKhRTdrDlvdgvc9359Ot6LC5I726SM3jGTby9
rqDwr2SOcpKKj+ei5nt6k2YY9OdCw4/2kOaGYg3kN84iVtIyJM/hIf/y/eYO
eBO5fAC5sPdonZCLCB9oRaJoKnLEmDb8Uq5aBszGYHFnHbopoIIMyoyaxXbc
KBvl++VZQslxq72kSnPbPS5VlQ7wtpKDmuvTQECDlu2lgoZBV9w/WC0UwS6C
KtyFXVvr0yrOXkqJ562LswDGkAsAMBSDXQ4RdzBKU72NiHE0OeM3rC5OWTAP
hrQ2mFe8ClFnqYIHv1L9Re/MuNy9nj47ZZq+Q+qT8lhNORXsJfFg6zDis9Dv
DWVtFLKJlnUzo6VjRvLYHzfAe9m/MTkKjn3X0pH9G+ygXozZ0GL9jDOdRQcx
64eeSfiGtSbRPNVOSLsOAR6VvsLwbgJN27IMZT+ArpjEZtbWyVGU6Z48QLpl
Hl9r5Rkqwjmswoecez1GyXUj8e1aD4lSDDAm/qB86OzrhPtUYCl8Ya2gao6N
DOQReIjR1e4clNifnpCwTDbUBRz466yDRFDORZm5XUkJtVsSL/ngbxTiCLS+
TKEfx5gWzzsZpN5jtUHt4yr1jo8+3cCbchQ3xi3kn23hdULsR6h5BQfJkIzy
oXb2zGOmzzcMR0JwZr0OdTdNCJr8IBxYPfhFA1J57cBqByg3Jkw0QMxsAB0y
NeJPUA8MsoqtSxZgFk4qBnjH/dXN6uhBQhxB0X5xvtli1zLuAxRFr1l74+ls
OCyZc7l7NXFqx3FQrhEU/RRczzPGouRBkRj6msQj+e5TLXbMNlIZgluL6CBW
NyMiMwpqRBV4Tpqz79/rCe/K9jmyuE49lf9tCJzGeGMUK57fAfeoL7Pk2IPw
3OCjlElUV33XLkQ774BKuDALGO/+37zlozxRrcREdNZBhQ5VU9KeuxH9MjVO
UkZihFWTreCPHnxSIqK6vewPc+HebFmjqBw/FL1LaGVYl1+uKEBgUtWIYTNs
NIBN/hmJki0+5ma9xFM1YQMINCXEeKtD6wMyCEap3jAGj4UWBYPAU6hEHRGM
9mpyY5AOKYTLY14l/NiVAjH0zTO53s0pHHHaMTmKeSmDoZhVpsvxvYzz71En
DseFnQ8RDxZFPR0dskT4fexuT7KWgM04ix9LrWtGITnQDOYkmM5l71wsAv3d
g+4vX/WpEwM9VsNYPZAAesX88RIrG+ll2lZn8JLZQ2lt5bHLPZKcD152Yp9o
ObE8BWgOi8Db/O/jQaRbSC2lEa5bPi5LvBDx6sikL490XDUOVwzkzkWiyeAx
EN3KuWJx/A6WPOUTUnL9DWvwgJ8qs1GoZzHQtnjBzjd9nQbMrwzRp0IRvKX8
NG+cu2QIb1gYkH41H14kZva8+v9J2J8/ukQVeA+JH4aSybG1WpoGkBDw/gzX
6ul1lxBWlPsiogOhgqkJ9fEg1SPPNtsEbQgosLt05befqayJvF98BKMBbbeF
LFD2wLf9C0of+6SC1oX02+ND0V8f1FRutX3bHQspnVzXRUXUTRNjKxDHS6Rn
DOL0yxa3P1T4rNylKtZH/HI6ypX2xsJvGxf6U4p+cxXdzRVQ42X+2ctl30qz
jcIKHxppW3pwWn6vKDQcYFwrzXDPVEX3lPO0T/l8uOvcsb2P1fvJGuvyTsBE
MiVEegUfJ4BLxYNeB2LsISOXkWl81Hv+YR6rnqiR6iw+Q+jMwL6JyRIHHhsd
pDB/xcPAa+IkZdxT9pkNHuV6CHKtN6E5cvRc+oU5/BU20oXopFNAtxun8YWw
PddvOWBzmtEXoEgyKXSpy/5lmFNi6FqfEG0WFeALF8hZVQ2iMvrSJmWBkF68
ABeU6zXB0L0hXVhZMnP4QJBcRTXdb2fQerpqoBk5cesmvARa//Q5nsqAJBdX
FF6Yw3EKK7pd6l6AIZfwFJuBWCHPlWVycE7H7d8ZcQrV+v0MK92wWcQOzqo2
yFmlaC0qxXAeDpFRhjdpxFO66mLYT9iSK7b4KX1iTVNFFwugLSS7GOzj1bme
dkHBEhrK7YqbSDUuJ4+1CyIcMW9rnsl26pUaEXtS0ygZQSuW2UFWHOHaPfv0
pnQHQv8opCTHGuXcqztDMp3yfGFLSAUkxqZPvaAD9tE8r58fWcJlGQZXzbIm
Zy4wpnz9GfT12iFfonmLJMDw9Z/mNeLix6lfaqqMT15OFXl8ZegNK70DdEd2
tTv1IfQVMvOyPg8WdC3Zom+NPBrdtqL42KR2C0R+S+zclhaJDnaMW9rcsD0b
1cFfit74XDu9y3jYOh+RehkaItRPoUmTMzwNHTqPlhI/LJB+DIp5/hb088U0
01uJx5KUhNwkinNk4tUKhl+NOg2p0iVm8vRrBp5oDSIDo0spZWteccOawjPw
ABpI7g9j7du+QZeyDyrPzU7G/o/iZDyrrWzXZi5kznFY+d6m/NR6p/mPnW4B
Q6N5b6/P1i8TaK1kkX9Dfw4ZaPS8u3pDTt/11YKeMmuX5qP1RK8Z+z3DWHXR
DuW1JZznFuIhnnpqqUZde3uOoe3RYZ4M4JkqO1b3m518zXClDUm/xUvM3kM0
vNN2Hv9guItJdw5S1CVxKscnTnXVIUCYVhbfyroPdAWLYmCNY3FR+KTVJxNk
f20krDXGTEsxuTSSdzsdttWrceMT96BS2dsSiwaU6/o9rJ2WTiOI+xaoum7o
jkMZcbPg2u2Vflr6gEJDFcFCTVseXpJRcsq8kLzyGL8SY9Y30w6nLPNKV656
hGvqo4yiWv1IXQE29FxJ0gKVfhXwlLjv5P5h3Y2JwuH2lsQlMYI6g1ILLUbd
YvCMTyrjrcuQV7WtKgpNmKUGAVGvteVEBoNMiMnuwOIZLP9B0IpPg+/TnZR/
7wALALx/zNKkrciJvJ4EJ29M0U7WGnK42lCfcHzpcuwAvPN6TG8UIIsiYqZZ
qR1QsE5QIhWDyYJ5iNU8zJC3wd3yZnQNa9M6UduJJvJUHvMBucJVFc9ZsxPv
uWo0Tphm/qS0sy0rB8kQ5AHF4oBMcTIXA5pEAhZHqTx3kU85ivAoaLWmJEyQ
UX2efHfTlZV2m8XCItj2Iq4aGCqVqV9+/U4XSAmsJGpR6baVIvzw7ighWbpN
JW1vbLawSQqQzmK4OvmC4riCJ0GTXagR2WuEOrOqg2/qR/KW8LjcnDWwX3UO
nbMKLiqUTdjIjtbjhBrXwA1ItZzIEkHXQw16CcYjth4/xIJSj0gTPZC4JFx4
GbK9YI0LRdS7okn2UERkM22yZhUe6T3wdy+4LyauemkNfPZQnwSVE+EAkHHk
3TpYkJjpv+0E5rf+ZKmhVLuusXBVRnlfKIyF3dokjU5pPBGIxoLOtN8phF//
2f6nzlM1wI2fmNbxDvS+x2aNiLw5K1o55QjsYs/kvbmWpJxdUONyqsdqUHix
lsBHJS2L23iD/zhQ5KkmyKvKL8RdKx2smSiLM4BY34THxryKn0z/QQ4NWoxw
1nGsn2nxooBzyvKDlC8q1KXYSNn71FZ4qwkJBQimIw3yoEiYmzlzYM3cD99w
bWVyTRpAMGkUAuj41+usRu64eE+azXJ26EaOeWur6eNLoeMw4dy5zYDe8gGp
Mi06es9XqGZ0FH8OfBv1uAgjFGoUxnOWcOeBTLF3BrnQcYWuIVlBq8RRYhk7
tgeyZHGlAQSuG3uNYtRgOVSjr5HX/ARI70ND+8DJFBETxcs3xm5DKCYkQfQt
KJ2EdKiX9VnNCuEpmP+Nn2n+t/Iiy2RbYfAAHEf2hgZJ0mGnOd83Asa4I4kt
S6IbGjeH171GWij2jjeM8/lhawSZ9t2XDEpbvr+0CcsXXJf9nHP1+RjiDSNx
4rTFaT9JPzWIWUZmair+4IGBhflZ+KPy8ax9sy2AWiJK0Ec/bUEhObJecuyQ
+1keddVoUT32ZcXVMIs02yqmUkpXGos10saKu6nPOSPbr6pDC80Dwi2ZTxnE
8Kpf4Vzno2uxt030JUkgnysHZmq8hA9gjS3jV89CDEXaye6QaHXDQjVn60/Y
C66uM5ewSy6zizXXT8TFzqqqfoEB5IJoLsoL8siFbmdAkf16SpiUi42GQ/Dd
ivhmyf8b72dYoM0pxCyUYdchd5YJvm+7TND/e05CnKG8WnsnwAGPyk4EflNO
xw/MTxngQ36ajUNOu8Pfp+OVqgL0SPRXffNtd0FAEXoy5L0BiWTashWJG3Cr
LGxfowQBzqB3GkL4cryZIqCk+ORKv/svOFQnYN4Iw5Sq9nk3cYtEKwhciZM3
pPIsyef61Xfpz4M6EEyDzkPx6YxZJXLKOsfHLqvGjCHf7v3N/UyC7Fz5XTmn
nwZVuknCX38NwaYg9QG3zuHC4UKUG8b1IUkdqFHk6iPfuqtQCoQ0swVoJIaA
qLxLx3+EnL3oKv1LiprN1WemDWWtAi1PfU358NS9pfUeSeMBpeVoScrmv8WI
SIKnM8zTeLKQgQaUieKHAUrml1U1+TiuciG2kyocp5glGtEUapshxWifDV+c
RSwGbEIczQanNrb4gIoq0ZKidD9j8+gCkRpk+Bn82CroZ7yjfz66fxDxLxmP
oRKEzvpaqxxenSmS35WLL9WIjg1yk2vDv0Qw8+KKcbgBj9DFysLEWyzgIQV4
al2gLaYkmFQC1Exav9gFlEzV2ZiViSr4KB5035fm5shw74f2KgcQD1LZJ+fO
uAXDmzwqrYNeyanHminDyy17Aogr+NMrR35sRBQQDc3w7pTyZrhKI8odWXVx
lyBb64kSiu30BmsrlUtIC7UYKIU6ZNDm7Qq6B4CVh2fXMDpWdT3mtEVwZKOo
jS8hV9d1kzxMz5QdBXPXn7GMDqofDN3DngZ1cEDoGwhr2eQDaNkiIo3rBV1C
BK24SwUYYMBgChadVn16LaVZTcAnZO86t9z4eW7jblBHLGNfI31gkvc3Wgax
Yej66MLp/laQonYZGCG64OnHzRXAu3H5/bnzMVH7/gkO/FWVpkSDLquOs/Ts
a9rFme1SSWOKZbhqqYxzRh+yDjChTaFhvIEGjs7Izkd45GYdi2KBiGubQ2lb
xt/cjOsWyQX10kin8KkvDiYzuzEYGVGwpqoC6/p74EHXU3oLKRzmixl6HwkF
ulpwffaV/HBFVL3aF6/9x5zU16qgJ+Q1nCoYXyu0XtT9oSEpkXX6ZQH5Rd4b
NGzfJPXbi0Nyj2Uyu4g8teABMqVq0n0Xt8J+M4sY7t/8eY/4/66gpBjd0CKj
B6Le0QL9zfM9KTJC1D8Au8G+Ml0cav8M+AWnBa2BxhHVAYVektOQxsXlACoe
PeHxydIx44GEurMnCUk8oQjea/0LYhi9TXI/XTiYNt8ykUGtVDi1//eXqwGs
8I95IDDQlEFDcYKsQ3G1qRzKvcEoXI1BBGJtHHUbdiJ7Ld2iUtI67mOkHNgn
/WfyJaysUcMxonoSOIFVv66ZcDY/d7byQYXONwpS3597Mz+K5eDslYBHxUQh
E3nC7WzFKH4PoSPLqPw2m6gWdmvgrh2NgscNxG/SVccbLueDfc32bpW9WgfB
T0SHCrcXz5HamSYn4KoCjpM0K16APohFs/j0EE9PCtTkqH8UR+bAX+hoiiRk
7GIt0sYA86gWFJimdnzJymG5Q8lNl6xH63GuefeYUOyoHSBU6BsovymDtkqa
nG3ZVbQpvH05MfP/4ikx2Lx85lHRvSRrntZAWTsv7A9NJwzKZJV+ZHBiloQl
UZ89BOyxP1FoHuzE2iZY9AeFJWd4jm9K1hzeZx8N7ZVXJfhFTRGhCQQBVJaz
Zva68FqKND0Zhd5qN5j6I3Noet5XoyKqmOFotKDv4yxRBrovRTugynhaFjvr
uYkyy/U9yOxqJhaTeLmPDL8bTN8sgmk57I/hSMEDBXwbWnoetcFYPtAhUEpV
YbkVMPcyrHfaR840lSX8nGEBGjHL0+oCXpFr8Ap2c+U8xy2P2EfcjwS1qOVx
Dyh9Vf7xxlFeTN+ZsgcZkU9+BvfNLb0O56hibLxyEu9Fq/q/y5+nbURlCsCR
WKZTUMV9trdSdq0wBibUGIKxWpiIC2vtda8LXXQYr0gKzO89/V45WPrloHfg
mgSpQIk0t5861xO6rYlbPbIsopyblkl4MH5RWhDtgIzM0dPGgizRhW0DfE5Y
Pj9sSZ9TISWyAfKSo7VQGCcWiaOQfSpVktQqkAjWUsexFU+TjFZu0potBrMy
sF76Mzc2Blz/ATgBwVHE6cH+ZTEaFKXpyjIXcXMg6fcCzbzHaxv4qaWZUB1R
7scDLbCtp7m5OEEY6EQijPQfgK4zBsp3L697IuAvzYH41auMwyV7+t0HT300
vJTI68Duqr3E6sdOn+oWU8Xb95AtVrL+QcwKiFmPgB5DEhoZoh+03qx2Nzjo
avoalHb8kdzriZ0jwoid6OoclUHlzVzXCZk3h+QupZNaQNY/+lTRWMQ+ey47
HDtIZB39D6SwT5SP5K/StXp7qs/vt2tmigb4i2srog+6Fyr7czwQStoOc0/1
gb5zT5WNRF2poXEFg/ktIV9TYG3cTW9YHc2N9VUJdih6jkNAH1gXO3cFKyk1
GqCRqRrqLlG9AXNdIvBKZfHqYXnonkZBGuGlCA3XAgdSe3BBz7WYRWgMdZMb
gjgUd2wwQ2jMJbLCU3cSYq4a767etdWPA3ff0HJGBIaIxSNZC+c7iLJXOgOd
5xJOj/tZKH1OHjBO916QGIAM8hLjyy9kolAYyWwNpAJLeTRucg7LkamUQVVA
5vMbkVX5hoYlDdblvyGTJCeYVoBW6BzqF0LnPrlmThALokPuEILkrYizWFkV
BRaPJVJnoklzvFGjVKGPyK1LnfXyCbVYCdQknqUxc97+HS0huAajcxltO/By
E+7KLU68KSn0QoAMh9RA33czjhL7DBmjS9mWXgXA666T3Io+YiBUxhHrqv14
d0m+GNnXB+AC4YdCcxSlFeA00t71vht/wt2Jm+z0T6ZfsgBOgZuO9RPJdv2f
TsiiqOPL1psETnA7o+Er8NGbAjVO4SFTG6QuiaPjCiCX0FHuK14ncYSHGIjR
MbxjxQxMxra5jqWkqqXpuze4L+Iv/XBZFimsUSWgfSrOVfM6Qu3ngAp7m9Iw
MfQfLz3d5KV2yMB6+s0QT1otSeUj0CpqizDLazSNmcTiHTt17bt3paz9v7bu
9cN7vjPVfURATy719H3zP1hxSzMM8Wc2dT4mZQAogFPQwiqUb9spTj2oTW4+
FnqPC4XLUgFKe9O12W5sR9Vj9dALKdmE5NCJmAmoCZ3uHD3ChOyQBPFfbH+w
YGMcikAg3xnm2E2c8PI+0+tBMBOOOOfZvRXPedCvVtSQd8hovq3iwTSPEJxm
CabuJpaxdMqXi/KKmv31ZN8nBdxrjhD0ePBqNVbn932QUj/liFKv1Uxyx1o1
1YAqsze3eWMjE+/Ru/mTTQP0NVwKYm+z+ZcIRZX9wYjaCLh+rUHx5tcwUL2A
Fl8NTXVoQywK+jj9HylnMrC96NkZ/LTmkHBexEAqZK23Uxt3kQQos+sUMTPU
NLMODGXSN1y1To3tUUeSndTcJBA/KyEVM/nbD/ckjssU8OkZVcRw3bRYA0sX
ZUQ+FThFWk16dEPYoaBFBj/5sCNmp6DHoIqu790k2mtm1mF9TqfygxUVZwz4
WNWWYcz7o75TpOxrW9U3Y0SAGwXEcAO+14olblhxc2i92uZ0nesnJ4dWgWeh
g0BwcRS00LZ2oeCBtJmBtdkKn9NpkrN0o3+yGhh6+ysDekrcZHvYHnBc+OgI
pPODlNGsWCh2a3K8Tx6Vat57qKfcfX3zucNzINgD8B8Wxr7Og/920RMtHjLh
pd3045PHc3T3Y5O9GbtN1evPSblgX/sZyCQhssNjSBzuhQSnAn0luuH2v3+1
ZRsD2OIf/lcOL3ZWfms9NK0Zjz6ffbkswxZNTm2TW3pUfJ1dMwmP6H8FQhgn
mWRMlX7YVUlalY+NKjgvopelCQhE+zIEL57iY56g5GVkPxS/QJL6wOPTFi0r
hAzabIVmAVLmyFnyYa5Mk9rvzQ7lRgjrVUy6ZhGcGw0yl+vJXXagVB9ztVT5
uNQ4Ir+oc6ofSd6UIKR0XPsdKABkYXUYXyovgHB38l2fd9Qvfns5xVKzOwxQ
86JPd/oQnPaZrehJ0eQOyWPEmm2bxj2IUI3rDKf1e3jwv/8NdD2DEM4+iNBl
q0u5ECztvQj+QJ/j61Jiw9MUWsu2qP35R4SyuS7yeqoJpbRCU0D1WXheEnPF
af4a7IJWT22JnMKaKxb8a0629JUOnv3VlNt+MSPWjq6w8mJkMOV00EnHxKFz
5D8DAYPGHvGwzJt5m7sJj+EvKeIJHWS2wbGV2kJOjrmyqfeI/FhBGZVusZ+Y
z5CrrPFCdOcJLNLw2890JcF+k/Nwrmi4YUIvbL0Z3MdKgL593LF6kHsSzJNQ
O68qexd5rF/3m34LiOhTRhro6+3dRKULHr83AeSZ4Rp0pSt4pfNaM6Re9Kac
vxbJLgpnpQLMramija++7pOPbOk790XzdexZ2h+iawNUx5k+WTKShVXB7Muq
Ji0LwXzUzdtv6JRhOqRktmGuGbtpQT0AsbCbYrAg5B9v4+pmxoUx86SK6PvE
xcjgtJWSl/DKBVFrEwwIAc0vzIaonpGa2r4SpVSjjxl+wjRsS0S4GvGqFBNN
2eC2ZHhPE1X5Uk5XXi2Tndh6Ye+Yj2O+/JC5iKDtN2/U4cN4GXXkr1RwhGwk
JXWIAHdatYQ/l44espJ1RT1tFM4pcX1ncxpVbN1/wOyJw7dBDLHaAn8uGz9O
uPww7QEdKHxsl72jjg8MJMMGnmACl5P8nAnJ1vcKdKLBJgvh/pGhYhos6dLy
rTknrlzNKCSWHjGh335/DJAoTyMmYMJJCxCDTdHRx1bt/tuzivOHDCuEHthV
ubAItd5tE5qE7PHnlMiWCLsOZXNMBC5XSKC4WLYB9FOyJLdMwUbwwztmU4Yf
a1479M9sJf2NQU/Z0oe9B7NQfyCO14/aXZBq350tE2R2HcUe8Hi80xXghmw+
sZjwGRuUP0RypYaXE1dVz/D2X05fP52xRTAtsFy5A1wxtp5DIu39a4heqTI2
k3ZEoY1vB9EjfBWyuRWMEPw/l9i5/dg5yJ+PfDmFaQsaUnz8Jpz4E+E3wzwy
JKfWfuQHRROsjfk3r+0NVWwQGaCqHKyumkc08mrelEXmYdees6F1Wou4/gxa
PLVEsPpKMuf0Kv8rISateWs2gj4w0WM66dsZxc6N8VZMZD/HLj+rM/cI+8pI
GPKfblqgd92ztqgL2TDYMK2sVi0Ol+COIhTSXmSkMOCrqgX9zlOO5xiyNR77
YKWiMW2SqlRBq6dzGxPvzZGkSmzzK2x5e6RZwdREv1g7+2w285T8s+qnVs8W
nn9DAIyVDqXTfxb1KNdvOsloWlk4hvYYbU5sVV7AdeKoQ4s9RCzXP+IyVOlz
9sHxAObZV+cZn96cIOP76R5bbIMbMB95q6e4HclYRVlVJJRRZBUUd+/KmPmd
PWlMNpM5SD8jDxok3C+nEWBQXzpbEt35YZ6w886v6lN0AYzBDQHzM16xNPAo
bALw7MRTSZPhhOrz6HDS4w7D0x8OdWSglOZIMA0/fU9nvQ9iopjuHRvigXt1
4ei0WcEskR3e+/XTnN3VgwpcLRPPrME8y/gExlXMhXHne9Qk9aVS15JTOJQV
JulONbiN6g/XMSW6mi/uW8Leec9n+jDchbKEDZ5z6cgvWHSE/DSnkXdVBfeZ
QHx7i5caIdHIlYanwtOk/cTzppaipu1CkDDNX6vr4eaxXlnPfBAl7ViJyHKZ
FpIlAIjrgu2v+gHdqjJgTYtgN49iBEy7daO5h0/4XMxue51wMnbesnD18R5J
4T44u69O9O9dE7c0g+mYn68ltm6bNi6qhEnIKSWqp6gzAXxSMGmXhQ4wDNOf
p+i7rJsrH9azJWjdVhh/gdEgPHvs2h1GbcVhmLSymhH9Poz0K/30BTmJbMHa
pl64JAnKX841HJu+rks/l+EhgI7583rPaRgg9p3z0xaIYDaRiM0/4sj4fpcI
uY1ZeyqIRmidQoP0bK2GyuwDzrE55CPkxielIr+AeIrHiS9nK4b34t+h3X+L
Sh/29OEgkS50netmh+BnagzzM4TL0E+oQd8vN0vEcUW9rtYnvDRHk8k6j8aN
zhHo2GqynE5D9UfbqKP1GEoSF9SMAdC/ufrbC9+jpPCMCP9V2Cm68DGmbz4T
L7+mI0hNcX/kzxygLH6T82k//WEZlWJ4qq6JyOBs3BNuMWmLwxmYRiEwi5h3
uSZpIuhXdvLpTcfu1/aFJXy8u1UIMBmOBP6k8NHON6VTxy9P0EelUTKcCDSk
dxT9UelXAA5cD+VJEsQKoniH5ZfxMrYB+9/6ueP2oKJKWFjZyZQfIHyngp88
VdFPhXzCAUc9odr/fk4fzyzo/fJeGsLNTfGoW5HWjA8AzkSpWoWeBE0JOhSL
s2viXdpobJhOSrkhFX138CBMAzD4zTTjomhEa8dzXnWhVz7AmdvZfqlIMXeN
rIVGqUVBaIChY9TpX29MpbhzM9jkT1QlILkpPodmEj/GRHaAzPyOEBq4lspl
NCbLsw5M7sc9q6NoPFHURWrTs8MKarAB+DQbe1ZAv/4mgEvSV/kVH6P/saIB
s28Jp5v0LCf6kSlXLFnYtI3hK8NIro9C4MqBTcwk823Gl9OV9COzpYhIk6M9
s9/lqoq6f118+Cxh35KV3LAkh850LNYlkH8BfwvC4tVlTiW6CEXHCMZVxcPG
yaQb/uM1ILZ23K2GoMB2szQ8cii+3jLS/cm2VaiZw8I34mYML9nEu/3CuhYZ
dLS/+QjzigwyDVUmI3foc2hRp7+t9yGZn2LgZUAJkE0PDV+7IP97tG7sxa/S
fNOJ+O8MRpqCcEoEhxPwcOmK3336N/B3rs4S4tGWddMZQyZA8HoQDWZaoOW5
k9PJtSAEh5Y7RWqgHNp75BU63kgmeUMqgLbu4IgkONVwKPQzFz89rJoGB18p
oVXIq9wLT+lANEdfDigaOAQf9UEmExsD2tRsvJ7Adc4wTUHuvU2gEsHACpm9
zA7OeSJTzh9ckBymi4+RKqiAZeR6x1YxN2a/kjrl7Gag0bbscnQMFCJDx3n5
mld+ke/euVFC4OOQbWmiKsN3aM1vqD+YfXWwOJ1VMuegEmg14qwoogjhXV5j
8bOs7ke4ehkF086ps4i1qWlyb72rOfct611cEdTAi+LniPPUIcuz3owenXd3
+7W0XM7CeWYDI/jvKnCZlRFzjT9Y89lt0EEAfs6OfVxenGijJsz1VgKlQ/ec
Z/ypmIo9UZUCdphjF3zLtkjQ8wr218IU+YSUYzwbm3Ia1Nrfwi1TQ2WOY/ep
oYkMz5dKitB3yCnzCrdJwUpXygtnTeu3OpDtdS9R523H947VqhvMa7RhMgMm
dBWeW30X4yDdVQyF+23KrmFERJ9YITOvsgLVuVTcrqWZMerMHkZDMNz2FT8l
Mas7Wilk4YHde2PyfIr3uiTXGnass/W54z/ii8iwsdKYqPMWaaF67mk3VGOY
aJYGYEs4Dw5ySvqr95I66WhUOvkBfAmy5JpqD3MJplpZ03fS9rYMDpXNehLN
gXtu8udILiRxf+MipZkyrLa3mLDUWTVSYQOUD52UO4eCfs03u4FLxMDSlcec
3qHRpBn+0W4fp16vurB9ngo3qnlkXkbV3Qputo0wXexecMFjtntlEACaDSzQ
0lNcs0KBv0ZFE7V5mJ6yqmj7NPJhGhFPgH7hsxbXPSSr6IQSlF2KxPu7bFU+
+a5OQoQbFIXOpg6DxMec4zspZSDGRJdNncRgdIDs9/COfWgXzRpZ/10SDScH
SSSHx0XWUKD8k94hD5LLtVIUXprQ5Se88xgzr5QQEx4QGE6ppCVS4eB6xiHL
nWPa1aCRqkfj3AF1oWjNIkD4VZK2IodY1UWuinfuifbdu2XnDxIvnL5uTW87
UGtiAlQpJZ9hB4m6cAFbpcM/enTR0Tcsc/pJvLK+EV+LxHacpHMU/rRjjCan
Oo9WFvdnjXQm0VBAFEaNcVvMWcHAkf5hcFfFYxac5CJ6JbcPFZ7CtRroWOqe
KTnchzFNcT03/J7bmCJnnHWb4P+MOnyUochEjxpNb/qjAIAGoJ99sQSkXZWK
NwWQCEtBnGauAFcKMhrwPTBUg/8jrDUFL6bk7zis0jvBMpX/f2IEfVJD5zCD
lyoMU07G0vt0H3j16LVXA7FgMEVH5AX6hGMlT1xQH+vTCDkz6km+Q86Kf5K9
CuH+GMYEb+n26cUM5KvnC4KlMakRCXIMqtWTf21AsJzFE3x6sQ4WG3VFdXtp
C4CsyQ9yeFUpKNyceGFZw1V1zo8oG9ewIlDxHortWJg8N4OyMg61uyL95HNv
+wU+9PaCGFBWkipJKNYrr79fP+crZlfLuItzC4nyNDuFsnLaSgs23JqHzAA5
Uci8tHtN+3G5X+X4sPWAbz45QwED/9Ra5WJHfHGvvW/ixKZa6PaeCgdRA1vG
BgUjKIOnTQgC2+AXNjL9u938DaPbLHQ3WE9aGYmy2khcX2dvLCqiP+Ou1mOh
7Z0labE9vG+6P71Hdj9Gjkp+9WhgsnaFPPohAB/veO4N0Oc1wht2/wdcpqas
I+qZ8R8/fNugw2XYoywapyPDQ74lb+C07K2tSba6JFHeOBUxEt6mmI/leOiy
Hf5vYdCpknH53hwsAFnAur+t7+kCx3+WZrubbGhKRGs9XDhOjsbcaqtpd2L0
e/2FYPB849iwqHjFBmGOBy4VFJbJAgOu9y6Dqht2QSwTAhypwfKMJlnk/1Qk
ONTk6NK0NqccoC7RUpbIMA7TFGJfqiuiVRUwKMU8oxW8wG0HHJpsbnMWQNGW
ts9/UqeHWkXGoAnE7g6zjil75AdnPSldX7nHDY5vVIlZbhCqCJA1QQwlZBWv
YjIG+OKC0rX8Uml6baEuAbQKt3sbErpjddYe5SlNWTmLamH36M6xq2AZMqbD
kjL4TFYiLGO+SlRFym4K/+t3oORUnp2LtF9HPMhqUWz1HKsxnb4X/ej54UaD
C1E7MLP3mPStj0Rd6dYmB8pNB0Vy2ewqq4fyjvkIhCOQCo9maC3ENzAYkHCM
mEHpFbRT6cjhS7F/3ynaWEUuTcPSPwQB4Ol+k1VMcmJdKr1YX4ygjvI+1d2Q
a4DHnV8movhNXBAakelauyusDHNXwDIkqKbv6AFvUEvNC2efWTwj8NnlMUzV
cXb3tIq6mFvz8CCnFt9qJnyzfTV1kEu07ITvvQHuWnAjp9WUvn20fho23ImA
lqYZIvSIJfWPeo94OscKNjxZubqt6bYWGVIjSqOiNSvmHj+xyfwrCvbSw7Qa
OMkDOEGP/7ty7Ba51Vc7YFh93b/Num6SD2KUMyB5O8uNpNRABbKHWqzmh3Bz
Ou9axsMutt4NwVvEc0SURsuH7yON1aLui+0gcQTfdqc839A1O+9Js5hCsW0K
Q6giRISUQm5mom7CfFYLRrXq4fEUu8asJq09IeqzlyzuchdzDqpkX5c0IHh2
uoDu7tbtdkBIO/+j5B6rolSK4aR9CawFLX/mTvGiRuB3VceUIxlZXbiQ8R6G
7fLLWDXnwt0yUWbsJIfPg+gWOeymDbzP2J1RUgdP30HjJaZNrl3C2wszpzsP
MmyR4b16OPBaaelKyqJ1AHr6yEycRnwczWfXsMmPyoCfq+QCPMrPNGe1vSJg
sw8xyClI4L1Xr7wh9+l/4tpB/PkdGC+7OvRnoAxJ7Rd3PR4qvdtTQVtRUh9+
pPy3WdfY+vtkR++GxoZIally7aPgkhE+4ZOEtX3/W76JUdi53XgaOOJUCfLz
Nc4ez1ZQN/LWxezbRZtc9gKGRTb6cFdIc9TLOgbMVuLsUlSHw6Hfd0ymN0ky
EfD9NaGbzkk5R4EJ0R5Fz8QVki0Pwp1yx6XyX9ZtpGWUQzg+f+7In73Q/mFJ
q7Tl8fDPP7+HPxS77STfM3lLR+ckmffghmvdmjHGocKqVY7kFmqvYzC1/W0c
jmqzgTWIwWncObNjCwGb6CoM+AtyRAkOouzPZbJym0bXiI8xS+rxtwVvCtkW
GdEfWHkzG5gQymBluAlOmBvhoJFvRgNP9YgrLAvZA9HY4nJ48oeNHgJ88yEn
mGwCtYCR3l9ftph3uTVMFXtpibvoYcQnN8aWpjm+kF95BxxEbH8kFPNodBIr
KhRlQ0BEUWdZTxoAwImgKltXxlJcaCYfkJePAuSTvaz6Jwa+VQ9N6CoelWRx
GBXqDJLdR+aEEcrShSy8aZQG/cMp/ZOc7HPJm2+50DOR1vfvNrQzC6XsBGeW
RhWu4oPP6QoB9hi4bUaN1FdDbTyjCwbHioGojaFzGZMGpmAu/XmA8XHBl4y9
GgVVf0RQeyqeok/0Zvl5f5JEigPFiE8CfWo+YXMUMYXZ/p4fKe/3QK4DqGJg
0Mc1MAEB8ykZQqGblOdq60qcSN+p9j0rUVljWJs6j2gQXTgzEkgIIOcvlxEk
Xhpmt+VSuTVoO11Z8xp/ocRN2XZLq4GdJ/FljgHRwZAWEXlh6swl3F+EadJu
HJPRyJ7OZMkh0aKN/nj5Wy+G+xCPgosRW8o16OIaaq0C8SuKBxBg8T9WywNb
o17STO6Q+HMQDpKX9ASpZHyaJHjqdlfB3kBFqPZJDYCAKWV4pRGiL8y93sAr
zyRxzh+oJN4X8qOuPKmYrhR/RKekMsj4GA2mM3e4IoZhS9hBawBop29C0Fy3
iQdkdkPOUvhw2LQrK3MA9raddnR3HBV0DQI5Zf2QL+I0wM1VLS7LKI+wPq3E
F0xZQ0W/RUTiGzLrKK+Ns7pp9u0P55MTlvS7qRarUaoB7rRB37Bcga2jmoQp
0aII7PKqcwj2/GKXEItBTnnBMkcqAYp4shIfsOo26J3YNQa3kGFdb/fyn6sE
lM/t32ayINhOaYoe1IJ2+Y7/A2AxNBzXvci2qQWaBOuBxtf2DHuXyh5gaWuD
TzqksVdxaN9ow9yyH8ci4WGg1bA03W5jeQNzZ3zByUqz8gE09YneLGJzaAlp
LXohpcT88L2eYAymfWC2omw5GXTbFdYJt/kCyt588tFfV07k7SNlIeVcdmUe
hxoxhCSUPTdVaTlpU3mlTHHWiP2oq4X/Fet8iaJeAwgHBfhqtJfRlA7PzNxY
ysAPxHX6ehOU3K0tfMwq02dqjEBLJMz8aSrtz5Px40Kh/H2bZB3xUjn45TdX
2sN/uQmY6/b02TOpNVcAHoS/4G02imgCH0UHbjwQUSDLofXIQoBErVAEzktR
x4xpm/SmpGCJ3GhcWjscb+fgIwyVYMAnfJGgnQhvqLYM7LCNzoY9t0r/Ydw1
ikG3Kwer2SNiK72a6oA27QAUoXGL3YHq5fizliCV1FearNALm3wyORLNlAA9
LTEtzyXCVaCe/4qzf4AvgXAsnOyCXu4cwNN8tGLxI5g7K2ZO0EKm+LUsUpaW
iQjHBteYx3ruYW5YD1S/LLP4iof/Xs5IFqxye8C5hSCi1wA/8fx+KesLFs8q
pgcG9bGBLHx4yz3BVri/45ItiDlnkwoXqcIU6DTPxiN5Cu7RI/VXR6xSM2RH
tJr7KdPvlz5mmWf3PaYDBVX/fXW4wDD7bpm8lT3OmUB1tm8CQ7s/74ohOYiA
bDiTscTqB2gR97dBSZRMIll0NeLhQxDFfND6e6B7RWNnr2vyX0YAq75krFYT
faGz4Cwnust8h2p8oifoUq7ALPdtiHrgmSPB5QOrKNHSc+9jtl4rt3zqHMj0
b0gOHLfDwNCKSKYd0NOTnZoPuUxzKt+i6nJlc3Ofd4qHSDxh97Y3asesd/1s
RQOFLMJQqTDmDKs4usPKaZoBb2Tl8O40rUOgbHoAuPr4c0JCHkDn359SA2Az
oO3AsieIt92nhIOGUseUYsLSGsz2tOuTaQkNbFliqY0vrrQae0k/FQVHSVPK
WcTGL6HtF2pJC70L55mGuj55imlj/l4q745ekMeDcqtz0VZi7ww8TCct0aho
BJtHVwWN7W7CTv5QZO/hZBLZoq+/2vyRMrsjvCMhob3FxwL3BSs3m+UbKRoI
pio5tpGgj3uo8q7Zu1yoYbyCmGDFNfGKmq/Wtvdw1Fpax9CLpR9vi3/vrvEQ
ic5MUEodbco2uVQM1OtAR/UQoqnM56Q5hgIegX2Jur/FQRwqAETVr4yXF5UT
07r+2A0rbNuWKK8YlvDnBP8FpKFZAhqLvzf2vCysDt1jpEGtV+o6Vj4+sd8W
4p0TvfImcxugWNYIuJGY7Agd9OsCN2Hmc6+EAscdUpjqfv+anmzCvtHpuJqi
9CSz3zNFhV2NMonZtsJb0P1JJOwZte2iyxc0ort782VltZYArpDE6+6eSF+5
eZR4BA7Vrb2NyvjZ4/xaelPRAdw+Ts6/Ku9+Dokd266AFteKqUqDviBxWgv0
ro7RfNEy4SrKb6r71I6ONvH31gsNMqjcSfPy7oI4ZWz0jufOfZ8k71vToqYF
BNoBnme9hnchlI3Vzu+vkDA7BRzrF8SXj10WzFDOe0ShuMEk6oeXHwVsKe4c
9ABGu1O0K+fH9uWjBSJl2rzigOdpzZ0w4yJllZve3YFtxDjKqcx1wqJVLYNa
n4lr6dWohM2y4ni4PL1ngD3k6B5izMZwsD05ZmboEX4I2MkBNV19yw7Za32T
p8fJZ139reLdGxiLVtSjcpPonJH1y2fQDKJXzYgoBH4rUapBdtmnHh46aG74
QZcpe31QrgeAY0zLZL+ZIUF3jsLqVrzxw9TsreSKu31l5+X9u5RgoecZV5CT
cMtstzSUF7KJrxHemf1Y9Ikc90z1UTIyYtVNE/Gv9u1IFTqKKhG6/mRFRJMa
k2Rp0VzwPnYnibq5AD7Eev40Vfy61864SuhAV7qGUcf7ydF/Tnt4oE65WBb9
PvnFLpYV33cuwtCfWJ3duFCce8/0SE73AjaBIeE7bMFAs9NrEdeSmb41yfqz
wDbl+OKPDK1kxCHAgmKuaiN67bEAuVJXQ/sxaejm/7s3fN6c2ZTlXpLzz1MB
wpPbKJNpRkIQjzj/vV9piabelSlZPylpi6/x6L7J6OCj+eTQamTDY4D0Raop
5u5Sz/N6pVoQgsvLOozMRrXSqeoFTvYt+nRcGtufMfrLJ5VQm0AQKnZkLg9q
uJOk1jeLc/WxprUcMgbHeywOWP5GHVeZxZRymSq55oHsyOoRM/mYmxBq7aiZ
xrpvRw3Y1IieQduhjwmGdZFeDtOOOqqy9bXEHF+A3eeHBsNxUy9Sq4yF1hWq
JhS7ML+8YUKmCQYqPxS74bXOUcC8lw4yVmw7feABLnS6AsKDl17hN+PJhBAl
fXO0rIUC+3QM0RuZGrUADFt8jFd+/NclB+u440wn8ReRxvXqcl0/Zk1Z13vc
c3HFOFk/IXXRtIpfjxycXdDbSt8amH1Og+CvKegaClvpXJpFjk+7frNR6NI9
8CH+W4Bn70iMNUq6usHCMZZ6WtHnT0TJD51Y0Ppm1WvZBb0qzKfwI82Nzmb8
P6Q/1XegdQ1eTYkCrUGUkfm6Ik2oXcLpghB/EO47j+K5VlD6Bo8yf3q238fJ
Q5zXbSdhQKg2kgstn7DbhmjinzuzzfHdEBEMG3sp7QtHUFomwPtbV9hypJcY
kEeEgOHcT7LJusul/EyJHPD/MY5lzvZzAbAMeZeQVfviavN2qphYFvqoMFPE
MCJK6ZfRXD6LoNyuDINO8ugQBwFYDZEbZNH5rcvz17a3iF8Vg69VPkwnx136
dvnFSajZuvrcDi81fG4X5InNcstknA4xYE8f/DsTvQeY4jC08U8f5Sb6bKrC
INdcA7S0CbgdjcQxQgr85pVSyMp4//HPiO/QD0/KCAMT7CnFqqEoBm6vWQZu
XDfMxqd4eXbvS6TaK2+Uk05iaqihLzKqxDt90dx+JVN76xnYXj/v3YW9WLEq
Ogjd904KbjBZJFbgKGbA/fw4GruIcEU1PJBtt8dVc9RRJyUrSL911O1dEv9i
nCL83bPskl/nW7jg6yBwTHNphtLlihwKzz3AaQXzWBDaBrM19S3MyGNwkLmr
4WTYKeAHvjEJGAId66tR+XCC4flcHe5h3bMPGIxWeZ0FsIuabkJkDItoB5zF
sIKdKqu8gHFa9JCA1qOIs9SIG5OPDuuCwBROZarh0lLqbhiv/jtkuPwU6oCb
Dpnvwq+YqbjWHIRdegjNE80S/5B4ks+RVbUuGix9M91OSZ/gF8N0jnbfLndN
yPDqfRChyISJ2cEaLZWp54lhiqVk4OqG2r13kbOIThJ0/H3iFxot8v3zdx+G
9OVEzMD0jpAFgReqomO1ox7iWXnbJLPWrcAgK3KzrbHNDQQGNohrl0U8UIo3
IkF+/vTioxOoYZ/fgqEchRyP+3++5lA8UisHQ0+wvuNWkWNUbA96v7k1CFPM
zmHOZuLW7uplbzxmCGO+jX3V3AIuxhXGALKZfxFqYTRQUkjbhcBBpMt9cTgu
IQCNbpQgwL0j863Yuo0lM0mkysJXJRi1hIwSGlrR64IsVPi5vfDv4vI/jOLW
c3APg34IfTx+BjI/VOGAQd0xMNGW+5EnX39bWgSVm4hwuPBH+1cC0FhHp8xc
DtyG8gqFFjPgSTYAmRzAYX3bZtWsmqXBCiJPCECaoxEYhxctgw/nxy2mEB90
KvRYC1G9hUYCdNFBnt2woKWulMGs3lhDW1VuY5qGF8yvWVW1s8p0EC9/fFRo
CJkYumBgzy3FM9RekxAB5lsj9pfuM/HotembW2/NJ8UyoR/aLNZ+rYlJxPM/
CdtvCSlkp4cTb+vNSQH8O+y3c4nQc4bVbhQjWIAQOJPFvVmcpoi6szFTCCgy
iOFwVMh2iQPjcwyghNCIkLnP1ge8gPyb53Lu/MtfIhBo1OoRdlv12H0YgGTs
wVeDiyEjUQK/QJnswzeBIz+CFV1fpaWIbD08W6XpOeAbu7j+JDNukGAlcWDV
VJaCTx8BjhxrYbjNY1BvIM7TFs2gIlJp1Zd5Yh24VJVf4pulf2moVQfrNgwK
YTf0AZgLsDp6n5v6uq0InMLrKtZ6NOApMZzytCpw2gasZ6DtP0ctTET4Q15o
2eCHVbncYXPTpMeTReUdS0mmJeCvFWi0O/kYkmyhfqA3IU2kAlaYNB6dWbLt
gBVOfGoL4tjIkcQwgVqrES3JduoCxQ3Z8k3UhO86lHOJ8VoCLwA3rALwuklw
3vq4r5v6htKzVKEH6zp5+QaDcPW3N7PdvLsbnfcr1dIUJdkTzY5WhMRa0cog
OBKmNL1tpnA+mwIRJ9Ku5mXwVne0/3gS6fg74om8T+mNNJQS7SNSFu9ltmc0
lHbdoX6CdMe7FnS2DQ78QsUMdj2jIC12MyeJcBAVL5SSvc4+M+tnbiS4TszQ
08UKGYlywyPOXXDW8wVrXRUMNCQApYTKtWyv5YXBRGz1CMN2I03XxQpJ8Uj2
F3dGJ+/sOYVfNrDVV8xwW2boCUSwqsUtykhrB7Wp9t03+3jQQsQXltxFVOIR
6Cbsa7mAlldHtNv7PcAFwm6PwLAojLn2cM/NhXxM1If1vNDuYrt5B+dhvKGs
VfginA28pf9UDBIAIXOKwI6mPELVtTWQiBHmuPrfZV2GwFUDJ5dl6W5rnsv9
5kaqpgMx5pO0UI5gVg4QDM7I+/smKieFZbMtET7P+aTFu4N3bJLNmGa/eNiy
IvI1ygy64ufYdOQF9PvnmrXnq8iS0Lwi3xn+MfikUT1Rs/nVnmHqMKTsqQOs
3ozfCMEsU5gOENhCxbWpotTt+9wlpiORwf3ekL0qqHOtOkEfPSV5KqA24U+k
ZzJA/WKVv4tERqpKcSfe6f+jwwEwTHBXb/VPkyxzL8v4N6qBTSUWp/rqKaDa
eq5VpCJoPHeF5iPGkDwNpJNx4sjr04Qn4Zwo1/ku0KO7TALty4CA4vhtiBTH
uHoCCtgxbBAXkN2lvhzXAfGJwRznlJlZz8S9Cq6YDNi6EjTAMrbfG2rsIP9q
1vA/xK/ctT6RKOP7bXjnz3l/0DTPMzbVHyN2OdVOcZFRlu33Wpv/TBmqn5BU
MbT8Ac1otsOqAGh3gjyndOQf+quCXaKZa6EOEBMK585xbCPxOk3L2QvmNgpb
pJUdcbyWU8ObTQQMHT0G6DP08kX0G/Z/RSgj9c4PMwS1jL3OnrRhftzwQFfu
qu2BErKBiBKmszZIfZhU7HjSj8TOuJnW/BJ2wombRTQ2nExQtxUiosFQyxBd
7WQOrboexjGF14w8Cnm8JzXVWTtPzd725CpyMKE7NorulN9zVkjn+X97vSX/
1j3Q1HW2DGOY5y4aTacjyw/VXA7GuOLA1mxYTprfa4lkGPE3x1jBztzvw/o/
MEkJ24wjZL+PAgvub8pYKz5OsS9LqVNmMhAer5RcVBjV53uGZOONkOfOQSw3
dOONB1iWMb5uuS7VikwY7Cez8jpebvaztSqkbkg2n5bHKapsDcbVvarqH9NP
okuTwofi5ueE5sPLJVAn9Z7/nlAavet0+EaV96WrCfQknrZuASlqFbvwyfGL
4yIGtBPSgaTO2iA5xGgiPAa/bzogEfMP4XPghdLwl92GzKUuAKNFa+3W41Hj
YApXuhUuFTpL3WyIwD2Hic/L0F5jcw6Q1waQTebAQv6EsXpm4lYnG9qWnWfY
H0VXEY5swyiYHK85hSXPqNZlmBFOmAodEbEOhlhWdDkQPliJQ5Iv8eMg0Xs2
lMx1hPf8y3GAJoNQBL5EtjDs8VdQmCxaXj4KQTbbbrIqyzqWE78Fhw30XTwN
4SJfTsgYpahb1R0tN+wInoghKbNAsSygd3Z5UybR3HkQWXDz+nX4GXduFZLU
AYCEnV7xk9C6whdLsp0SSj1jXtOL8TWxsFhjY7RRCHFDhN3qpNJL5uoUDUDe
l9bcBD6erX39olBiGNrZ1XrHFTyhJtDsdvRHLEacOP+SOoTauorAxQznVCQr
uk50oQBu+tUNlPy3I0Nq0wkXhggNaZ9UBrCWP5gkReyTG+30Pt16TKC1zIEA
uIzdDq1q/gRmMNBW6DKlid9PwQP4D0fRhf56zDDGLq/580cp3+0TdIF+ZsAk
mZeJUSF8vmIKZUs8SVvnxYpyjCWdUdl5isYMzjcfzbPcMMtvw6Nd7Zkq/hRE
ugVnzRxJ9+KdWp/VsftxLu1g0Tul0GNnQsHchK2AvCGz4KB1pkGeBW4393Au
Z1S52OpGivJZL2gEeXGc+YyUrFHvIUdXCb+jObGM81KI5XUnuMhJsLtZj+Cl
TILmCQhANS+UBnalP3szQSO4jcCI8E16/UQ8iqymID10TzWdmctKjd9gnaWO
LvVcUsqozWXOorBHvbvKWpLSQJzpdPr4BK+LG+ezDQaaSZyO6zInm0vUHFTo
8IeT/o6ZyPq/DOX4KPDJ6HnubT0pFGDfgyL3vkcOTxJI842AYPNMmgOOiAkb
rwvXHX+8Ybm3oa0YS4IaBZOOMVQ3skc/foiVZ14yeev0KCYC5uuJoOAImoJT
AqnlEp1GvmFBmtJ6T+SH4UYAFb5v3PIN9SjqFNMbbZn45VVB7lnZfV/9VMBB
dbhDX1Zg1KiMHUS3KWC0v5/G2icE1DK7FqIRYqKeYSCYObPKqbwyT15xz+SK
Y3iMhUUfOnlMI3Z6mncgK+jVe5dpGo5BwvcFp2GHDhm2Kq5KZ86CHV/Pa/H8
maB1DOxDG/uAXnKR6mirno6oFNPWVWTZjswY5dfF3oE4kDQtbZgMTXo+NKE3
wNx1uLqyhROpD3w6MDfzPCXc4KB38+Vr9v0el8jRc/XY9WLhjJ12Wk4pEYFL
fDF7Hd+xVpUzCzam9yw8hpn3B9fUU3oHX0clTpJOetuICZJrgAOiCjBgEZLI
lRjK2kEJLb1IythG0qvOFkQziXLF0oxn/2Ziyvps+J9Z4e0A5lTRf5QDx2lf
UUM5/FcyMyGApzYSK2rmoGEf1tP0oJIdUNr1biZPQz208sViyusFFc7Qz3Y4
1zXBvKegjia7yzYgDdabPhYNyqqYCVu+cS1Ev9P4VZ5YQDy+09UzHFv1NTPt
QoMq/ahatMsoMgf9rWpmUsgFwOswHSRwNBMHO8GqucQLRGs8GvUvfwt/LDbH
yfLbSk26G5/vj7v5jnGRyD7+O4+fcH5S4SvAOeWJY1ple6gFzQ6dkC9kQJw5
sEKxolyi2QTV0T07WebDPmpEHygl+s/5IB4WZJg+RZrleNu+HVRDJ1ibhrEy
wFvivZvivdjPJ1/I9AhqOdbZ2JEdENmJg5WEFo41dwo4FsVASUMlQlneR/SK
/OirDCP8VT4P6HpxvLCHBXCl59oxem8zc0WdF+wxz6F7BuzRVBczt69xeHOp
YxMS5Nw1KTAZyRiIip4Yd0tJdHnRb+ua76m6R5aA4DJc6S7fUvxRAylpNF1I
k0q5HYVA02bNYoCdJtyHn9iXUJUCSyzX77Ghl4ng9IGzwdjZpcUvoZkeZJfc
ftJV0RBUcXAvvN/WxvsRJG/g6LcTZSvOm4cZOn70HdOR1Alm6wfRKCYg/Ddj
bYeuh9rAnJCY7bbd1kprj5IYiTDUQrX0+vQP5MUa8xY953LqXg2rIiLoicL7
5nPdjJeGz0IayNXvSDAsOg1Ds0jm7+RzYOLfJbf+8xdkdSZIoCnByI9CsRh/
MDiCd6pw5Boz0lmfOtkzB5RSJ9NtKaaWBzgC/CfMx/SGg2QkmeobflhNo+yg
S1QPwLEMiPKan8m2/6o0BGhZjRWnNAAYB7yml/13+6lOfQnZqZTZpJ5vy5gG
fQQXpGpY7q4bwwyG1bycodw1R9M4J6w//js9Ro0Oo5Jv++6qZzh1ysv5YBKj
H/oI3WtUx93aWuHdmL4tD2Ie7/JS/jRvrqXkMW/nsnoAqJPQfVz2zTtVbbBu
KMe4CXVLRiH6a3z6+5qOVxcKTzn7pnmomc96HtxAmBjDnGzTDdZRsxnyy3jv
af7Fu6kQCDb8RuGJ8PtYCr09ylOCn1KicIEvQecxftMZcNWJRhgafYPLBc/b
v8H34epaJaG2lp0vUmPB52YwLch8quER7vlizoxji+d9WQCW4BwTH6b+67yv
/erQFs1wwc71mklZdGnUi79RF3g3YJEuCVlTnbkxqFHw9ZaxU9qjfccsm7hb
Pn3XANFmYf5WYoDDHccMuFv6OriJK6t+xp1ir55zPZNS8CuCU8dgrKdCTul1
uhT/UgGeEx0jMZ0rbt08RWr//q5+tDhOx3vbVXTilzTdjqq5gFPpedVak1DP
IOVlr7ZTdp5ZdTRLeV4ee23nCCYx/ubT6TMsHI4dzlkLHSxR+INg7TSSkHmY
qKI51c9F8x4zZ0bk+EOuenHR2+a92Cp9kPZrMsStYCXjVPrNw9GakrnXRKMe
0eiTH3ARSZnIj5FQJxJ3FzDts9w0H0JlfwZiJGaHc5B94b5kCzo85L2n62q8
hT9kmujyeBAMgs+t+IHw99xiBjT7vGy9K0aqHg51uy2xkKP72tJxVXxshxTV
yr1fguL2LVMgK78xPj2r2Fls6njJ0+Ibc8xurQGJxyCEaXRp4iGqGb7YX7kO
+xLPqwJBAeTNE0SSb0Rk0N0ykF/RGHispOALGCGnqX4C9lCNPoS3vdiQ2Jbc
cNWRl0QLJ6HGgcNfEzDbsBag4Iq/Vi9r3p7ZgehfW/lx4qp6Pk2+KBogp0pH
TdeV4sWH9nPAdfjcYSGsj7wxQXW8GJGCNbphWUjokJjmK/ddoQyfwRtIsX81
+xPL0NfL6o1l6IUGft/iEeeiKm1Zq0iiSFJI9Y5WccTpr5iKjc2ty1HuA11X
N34zK8CqW/sAZEv2BgzT0jROS0JSegPPVlH/F1E+whk+qEPs/kZw4ybRZxPf
IuLMJpo0WznWmXMK0DkcFODa50CzBX4allh1owruS6XH3/VyrKueTq/2Vz+f
Kj9f+4ANt8dr5cl2dUuAlPe6X3LmXtzP0NaVQi3krOUr6GN3MyACM0WEaxxf
l/u1TZnxlunGPz0vloSqjmJH9qQ8+I3r1Fup+DbBPQj08N04e/uh+3qFozdN
i2f5JEKe3hGCuX4aGlMzpg+MzK7zev1JltEAWQvPcu+jKQh63i6XPvqm8J0f
GRY3sIlTJOPSUf004AISi/9EjPzgNPjwT0SohuDALhC260y4GKYi4Xqy4P8N
ZldcBEYqOa5RAP0x9zRokOMlYLgT6lIBmGlQfEEbZGARGzt/KOfFcgdpY+dy
rrJkvj/nwziqMSxMeG++7/zCgomNITOnTsZv/TU5/eX/MbTGy+OeexXVFIdB
SIvVDsO10qalX8iDuqWS4kgim0SW8vTZwlGYpipbNzplVOVtAPAzzPog7/xX
UQQJVsvWIVTyO3nnov8Wc8AtmvgaEWoxc+eYJ1RPwWCl9pZoidi8qhGoweMR
4oLpwsYkqIjJ0/dQmmqjGvbrI/b0Fx0HHKZwM3a7XsW3UsMLL1UFkRJOduv8
BqmZHeiC69EeK+P2Rl0FvNF0Xl3DwSu/nrUCbSUzDyDahYJdnhPdYTdYUKbb
yD5JnF0vWoSghCuh85MUczOb2a+bWm2pdknX9beL5vH2ndzsk5sUAOi+wPtW
M2fc05DHfTk/J+LMWsN0EDUk+mWkQdyXDCJM4cSqNILLQc4ov5OpQHHZeop+
rRG9/DAmOFYvwJy18akyUL7l42N8hecM4EhmG5a4xhId0q7D/uYiAVltB7qY
7amCMeUktMmvL/2M9uvwKDPJtieLz8tl/T17LP4WiyZIeCJtC6oBlVmlsq1v
Ljp7SkbRTMYTcxJWdguPJdC7bWCicPin55A5I9aN97W5v2kI6cgqykV+ghKM
cVBmQCfYcqCL7iqMQjel9FPBOlAr7C/07gDnJMaU46/ycnqMCHpiBozlE7pA
dpv7Mq0cSLWS6AInZxobxlOpEDQdzcj4Cvl46NPs1ddB8Dcjh6fWkAZ5ePJz
0kAMlyxmHak32fatpzPMvqfWSZg+gEujXNFcMv88p/NPBLGA+d59cvK1wYbY
l+fpqKiNiHVXvCsTUIUhswQV0KioqpyoELbq8PXsADuOObblPXPMryX5Elpr
UDb7uoqbV0guUlgBMR23/YzRvdFNJj43WuEcNDEgtqnciyRTgQf+IIN/gBOt
1EZ0mUqj6NMVPTv96qWVHs4NKeFF3+b59pEgz0MoyrKBW0KT9SrZXXbc4CUw
LlirUZ/aENRqrPwKbjrPGpOC4lC4J9SShtWrkP46RWoOX2TTp0KcOtb02MMV
N6teFt3eKsE8fOQWlOwbwvgMTMuEtADcA82afDz87optprmmUs7017E6ExWW
bae+G4OIK+H30Daz+Gf3IUQQnFp2lwPy+vxOJDF85SGAcP1wUF9rfe+qW+Vr
I2QPP66RnkLUhyPt8KgpaO+glR/ozZozdWkrwLBhH6GWkJPjHASyHojVW0UB
iJolg1wQMVdppCJDmpvPcc3xk4ianFFizsd6g9DFFGdpacvQcOJ3bkAeYZjv
TaIpaVq69DFquMJZypLEc5Kw0ZAgulr/lzOsAJ3REv7tlP5b+/bSa/D0A+QE
bCa2FdccF2hivzV9ym+/PmH/GfJiGnz3c0n39nWTsB2wSE9oDqI0GoRGtT2E
wIoX+4Y+b8TcoSKHG/bKU8YKROYG6fHMIzUz5yclKBcBJ4LkfVDuE6Qi+pLl
BE2pYq7XhgJLlMXrIF3G3+ldRgqz4u67cmNsH8ufvLmmT0BLnOeqbuln0Rws
0RoNJq/pCVtQRTIJtbNsAsJc04HZspgSCDyz5qxmoCc9wfwLf3IXNfjFmWt9
DzkSMxF0xopSay/x1T7TEBbIlv2RtKn/FxmFgJ6RFKxS5kZWmi5UX4qoa3WR
IkFY8BQRDzWI/dopSKAa56YU3u2dWgYbyRX8yD4d2Q3lcKHjtp1sQpX9b/6Z
74xLQln5OvUi5E5wMiYMVUiG0MuztQbIcOs8St3+n82MgsjXsmiVtYgqz4ec
dkzHQ3ZiAzkFUN/91lr8T7+bbxOwI5VKnmF9I3W0f011yViFe/JikPnbBtMn
6p3+FXAEfdA2hecUWR1scrgpqNVIf07372Mf3XmvjI+VOTDPZ/iV00Fw7zow
oahZ3NIE9ram/+WAdcVfYAoWdXy7TAMhkUW0oPJbRH26oCILy5ybIhJXzlhD
WY9E5l4kwSTv8zjKSrFxHkSjWGXQo/uPbM025mxenTMNppE2y0TJ+NfzWvj0
o8nhoaXCxTVRfMmzwWS+zph5yFgSd91tkMJBMHxBqDbbWiJVZjfUPEjSZw/6
fogGtzo8y3NuiaGvzmM12DM+Z6HKt0LDlxpS9lEi+L/GsNfr6dffPh3ETK/A
kWd3p6XQFyeGPUcmTS5uve+aU1KUZ2qrMiHSKxEGrKc7OSd1XPW/X3S4my0t
PBU/yjEd6oJmZHkZRoZkKNNFyQlaXeuT6MD+Hfc88K0x+FlC6cP/zA8dGeOH
WmpbSjGbpbvNhsoBznWRW28xmsRvm8B8WBsdKrn102kpn9YDykiR8m4Yl23c
XlsGxyrv4Cack68eFsifkp/MqSC5aDMetemZrCr9Y/TrpzfOYQBdu+Mm3cbA
cq0xoSS3nb/O5VfGW113l+OTgzpfrBlJvZOjzp3dR3Ig8Q/swHBmaWrW1+OQ
Ft3wsghqhqI+2G+mefm3XwQiyycLByj/ti1PIihrTJjph8wT5qt1lHjf087V
Qxrf29fW8Q6b+Dqkm4YQFGK9iU/un7+9oReM5x+QS3jypyBGJvU3nldfasa4
+o50JI0TOJZzK+JKdHjTJJJBpvhlruR34jT3wzHkfPobqmTd+96pEPZ6Td/N
1eokeDXUHHM+uqhTGej2m/l7zm+SFaFe1YMgYYvGAU5ncoyQWCj7gDqdVGAv
E/Eke1dljPIB04Tta2nAMeyBbQPXN1PPClrN/sJ0L+v0AdKxS2RJVEhpHLgF
dJR/IHDC1fiaRx46soHCqYB1Zi1LLPnrvQfUGltWlM+rUKa3gOPGHYvmoy3N
Oq/Ij4UfRE68MOCmgy313ru3e3qnuI1Rrn5/oQTYCoJYFf7hiHiCEraub6pz
SL3T8uRe6B7ECKJWUVuqAipDP4SAu2zaXYGSw6mZTV9NME3A74yP1Cn9nLOI
Otue7PBNoGtCocwsRygCegCPMHJdCZhoGXTkMreeob+NcTyUz5muJgl6ejRF
lgXCBaWE/iMnZInRhqtYIHWLfrUryHMvdxZieNoZKaBihCl7eaFJEXmd4ZpU
ztK1iLHeEqDak5zXAvvawRha77neiGeBFkoprMEAgPoOqnE3YcaDCjCUHvMd
GfE0FvSvb4MOMeR+R5mw+dvzCuEos2va4qEpoO5SGE8y/vYPegfANQiobnY7
Qw+04cnLcMrr+/UOKOb11GvRN5nMs5GIqpv6SDXfQ6EqTDaeoX1TWhdJmEuZ
nmkSrHaH3xtNHXTBxyFDZPxQja/0KIgm/dnl9DttTPyUuX7AEhIZO4u4027T
1282AAynU/OOFWB+5GcnynuQsY98WKgB9MDOP/495cWRFTe2gThoR8fVJKnC
hM5pcKoWzPIn0u9nUkyig8sO8v1LksmpWbKPdD9rqvfg7D0gKF6h1IhaS666
VoKya9ek/O+QCvIYLpd9kwkbKP4bj8k8vPSgMVX0r5+CeXLrmhvY3ATGZlCn
HHrtjDmTp2waGCGqfywRgCfsC9Rb7C1G0zBIit8mgTllcOd+H3M++4f1oATW
JWyKhTaiPh4D6wug4rP1YXMkjT1VxY2r1XjPUVcsngzn3MGjaASmiOK2XHaH
RJaV9pM+ss8UOLeWSGe3sQtFliqxd7HTPiPPLBs/dOWXgjfkwivnoLi+Epia
+7baF9zBXd/+u5C6DmqZfKzXv+gTMcg4yJmGnXN+prAbOicP+qYs441FqFP6
v2F/WC3740i9jc6RzadZ685OYy6FV0ariaUDoDN+xiBHIj11UFeuPjiOQfF6
G3YgyxiCvOF5VZGAWLCDPQPi9FFWOF2W0Q+eVnNGIX8CsQFut0B0seY/wSy6
QvLybfFOtKIBd/tLlXCkV0kN8FzJf6QRbQ5heBh9gp+b8dBNgTAI34LEF7F9
AA2/1F7RMwBD8fZ7MPv+LFnqNGLRywI/6vyynWeFhD8+0U7/Wp96Cez2yU5q
8PnHoVJIXQICrpZSX/S5JaMiQMTjOhlowWTWhNEf30/qOfFiXAEWhIHjuR8y
9pn9i7wEOY1kfFBz/AWT5XcONnYnZSKzoabbFH2vCrnoMA2WZGjnvKCPRKDH
fCj7tqHulUMeJ+LFcCHJFYdOvElltJatFPtuJQb8a2pnrX8608BlprhdM4Va
LzM35uACLHiEN7vgZpyvjnRo/6HeDy929JQfHqkpVc37s9n8hv4jXuD1E+3f
zY2GWdWa+OwVhR1eYENIjTo8+0ISX1mhHifP06rXcPbZ/u1ToMoookbsryPO
zc4ImohiWlJtj04z+u5S8A3PRChEiS7uN1W0t3blwbTT9TDEpqW07QavzUwN
1u02lpKVoFJ+3r4gYXuQCAsuyDz5KtF3uOqu3KUsYblkSwgdi1zGcx9OcBCZ
3QdtvM+1HmLGMY3rNnqRctJyIgckBNqeedQq+h713ikhBZKkXSlbc9xEVDsm
tyLupTusuV5wkxYqA/CH21MDGvTrxztjxgotfEFo/prEG1HFnTnKW1UQqn/Z
CBesBkja2l5KFi4NM/uLoNgLGRjg9tdd0MXN72FIjCDN1l2B9NgqN8afzyyo
PPP0Gx3MjxVV+07kQ7I+GnhVdrZOs5i3U6J31Yh9MajGJYSeo+VWHCqYl6jD
s14VdbPkl36EfEeNgH2HJRyjW1MFo/cz+fkrWMLhKBCpX/KNCFP55w283pqi
lzn90wij89+CtGuCIZbvODUYUYUsqY/N2RAX8moCBQ/dg1PHNu302y9/VVSK
C477aQDxt93n5Lul/lLBNU/o9Sb/Z9P+ocUzXb/QlUt3aJRpjq9A1tfEIJaA
IBzejlqnsXdiX7UTR4iCjaLi0evfdh1QFKJ7+1Ha5zj3WwAYokwFuoib1XcI
SMS4XUl1p01Pm8AbCMB3qbmq9HrTXPloMaECHCamLVJMFKJreB80BXjGRNei
E3HBrEtyRJUh8bB7fcbeSmxOl6GuK4VHI8LvFZHxDCMf9QSqgP22bJdUzuGq
Fa/4jCpfQm5MHCs/6cqYqbVRrMcCsK+zWSG5iiERZtwlfc/UHY90yVtSIphA
49fD5iHd0FzvXNQR2Oceqw9neDZ+S0n41863N/E5b7zQj5FicuFumk48ccJw
M5llTzhaG0S0idED1TjG48EDlyUJAvGtIAobCz5NYjy0WAM0VrfFLyFpR3pN
4eXv6/uAOg8t2dStrOX/rqMlTnOF42Oq3XcHKYDZ8Tme7oboDWZqIcMsieI7
Eq1pZs8Tx+NjRIXifFTEbX/fAQ7DJiAbHsSIxb53CBnacyrT2mRUCMT1wRyO
eTtuNRgriLVaJDcvWmQVIL/lJhBs/XBRkKcqo7SASdTM4KVi/HbFg07QBozp
7w0yYUup6bqS76TMkMNjWYIV3RL5gPQ2PXW8g0H2Enr0zfaXIZ+WGxy+3ui3
yuV3w8xnZJs9AzBPXr8543IoJp7r/ZXyQ8KR13tkIl2ACaicZDjTirtAbHr1
pWxu6OFunjoILevespXOyJKm+io+MDuIOCTkFHUzdeEzcPw5ybRSuBCPKdt9
25VlsynlgCoFO35Ny/rR0FVnXRuqtR6Soarorw949aCj3zT7YU1M0pO7WUvK
+Xmox/KYuNcKyANZ3QeL7tu72Leqj0Ks4aWCUOWW0kPUqyho9RW4d1kwfUDx
aXkp1wBqhtTZwBg9q3YBJqrLoKFw1ZkP5DBZ6YXutCvvFNA1rMh7LxZrM3BO
cM1NSIpACysSikBOd4gf8YgxVXholP7KNyUTuIT8/GzcMZ+2IuXnhdKpfz0p
6SIlb4XmJr2/dpBmHRk8UED5cTMS8CvIZMFTQPRjQShVxjMO33uBi898+u9l
LMrgO4eUWH3Vx6cusANeuCOpvRmKv7xNOgGI8EsyRRUdlMEwPY4gTQp+IlhQ
wNdkAExhEl/G8WahadsZzOmcOjd3SV75K+DI5ZP9E2Xl274vaI3ZV8C8HRDP
MPuyqlX1SxO3R6BqvnafC1LFOjzJVNgt1Cz/+zmNsWWuh0o+MzEOS15Rgv14
AuHOLLgHLkeOlj1e+B4SYmOOF7XcR46DLNR9MyPBGwFnGbP/5/dmGKfMqV0P
oR6l9SUjrd4j2gCQy9jIvLakMIqkKBSUvpqkvyA8aZ0uiekeB5E2ILznQRkP
EVUYq4SzUxB04foRf0LBP2fBAH5ihxWyhceffZMYIbvppaXrNY9xBqxZT+5G
5afOa6GMm3a2gCQfXBcH/J31b6tgr/IHzUd6CipcdHPZr/PNHh2srd/oBONk
2XkobEz3dl5otcdtO4RLFw7UzuNMlX9oFAg+RDseofxWUv+ILDbr/7ElSDQD
DHtXFzlwabv26J59zOWYlKPOBb3yKo2Pz3xB/XvNrsGoxL0tW6tycXkbSWhR
kAuDk0inCpqII2bdt68xROqGKEit4b3sA+0s0OiCk5Y0Par5GSVYVhqWyx67
/23xw0dFfpQlTadj/cnOkSxk2bm50uK1i11kRk/OaBKFRKbD3O3vTxpsDP4D
pUN04sqHBC6XmiVNvtDZUY8XpvbSxqKdIVwBqzQf31U9UuoK5FBwgBy6uf2N
z5keRQ1lwr3yBg8TikreVe8Sf3Kau7SBHvSskk+EvHGEDWhCbZBWvGuM5XSL
Vjzo8tHMe9kCo+SopTwFNpbMKZPAzkoJiixjY7YGXj68I23/d1cgBtMV+nGu
IOg9d8QkH3hErgz0FkQ+bkSI531tjgxYLpy5jpTmiUp2DrEw1YmSTzf6HeyT
iyztWRaFecorf41WWN3F3s2JfBHMYmyuZDKwNxL70z5QUysK2/hqObABd/Dy
YwwR9uvfYqqVJgg98aYqwxcDqXyqOraY1uGRpHJ2HBRyc7NpT469sFqZD7OV
vehnEz9U2wfICwO24d2tPDq6N49frwu/GfhIrkgdXMszc/g1dNtexyfjO16k
8MrAAP6hvX45ApVTu5htipLi76YdZtAkGDIJBIaXWCi8AsamYB2Eb4+DdG3A
PBNsyr7DdMcTWDkFGtvX6dTgHc4CgyWMpnNHEoxVTumMEvFEhp/KzJjRfmt7
wlAKG0t9Wx2RXkJZU3+nUNi2AQnsVS3p9gRSDrimE6KLKqxGaXZFj7lTcd3X
4my7Vdb8FA+HjzPowWqBGL252pNdTmYkhF+peYaBk5XFyX+IxKWk3+gHZ36e
9b5/7BQlELAO0OnRicrNEzqUmPmMWguJZx7uNxpRLaall8hGXt9Ae5H9fk1r
LME55jcH7RfngqnwgYWes8pIlnEu2qgutCdLC/gY5jxwN/GenFo8BlLLnH9b
c0ePrbuvVYC0fqv6bl4PDLK/Pv5pOYewc80BP+OK1kzjfp/2vs39OJs8ifYH
eYHB0SGtAEnwkv8F2M1uYEbzlc/4Ec7cVf2cea41Q9nDM0vw5k708a61DEZn
wJ7e5FrpXl1rmokjYfhCU8JFPp7Pk6ELF35wzdqQ3dr4zuuA56v44yMxxzGx
yDQdAN7viMwpL0pgAd+NOMHN1rQNBUVAxobt5JMBm4NPwhNGsP1kS9d9641p
HWvlKKDiGmEBCqt8Miz+HDWKvLn/LWm4g0ISqaH/TB4BeVLqWPk0e9h2FYpL
KjWi0xbsAUsBOe9On9LDhaz7d+816yPg41t5hUxvHQr3IeAFaDP6Cv1E6NR+
1jNmzjha0bNmIP84hqS4hXhSRJBpHcDs3o2cGCurkmcCvPlIPKvGy/XcVj7b
X3THkJXLtHAsFpypyAD+Pfb/jGjStaDz+EQSXOHbX5klvf4HRavQzV/sjhBJ
x7ID5CdvVSVJO5NrDBSFnzqJeS/+hryZbemeOT6RWzPRLfXsv6Bw1OugcQh2
VXrlIkA4EDIY1I93Z2Md3B/VAwZ6fFRbTMqES7odll7ZORVZ2G1HDTpWg51b
pyfEtEP04INobOu018kck66q/Fi3J2U8zZrr/38XU22DJjs9RwE7aIG0EkBR
tEKFF98eC/2O6nS9DffqxJzPhZ3a03cYMVZZtKvEb0/ZiS1BRyPL2/hT49fA
MBnf5pIT11JRoGmpvqtrkae7iP4asS6OHbwJp6OtKPCPFErS1A9n7E5eRj+Z
B3QU/Z7PHZoZLzdYZ0t2TY52VCqFnrAngvAiDnAQ+ubSJSu9GT1dqa7cUmwr
sJJiUXfsKfnAMhRufgB6X1iDuKW6jEzGQuZ6rbzjjXVoPuQD+P1vq+3SVyS6
i82pxh7OT26RUNwMz2Pxe5cB5iCJm5lfwXJEX9ZXiRYf4/jsD2WdizcPGZYw
Db8D1umRl+4aC206MezJn+Y8vJNVEg51H9uOVxvH/uXzt6Igu0yzNe5B0fGt
XhKuOeew07qOKI1AaJ/46VqGNODLg/iiBfu186I5DxgEERClBSYS5BLqg4fu
PWCWDJkcx/Dag5c7mSkgbRlrgYruEUP66mmK0NBE4SqaMn4LBW7eIk0CjFCA
ghHO+TwKesMTHN1vkHEsq1k2keS/Xlj9SAasC1zUsQNB272o/Okeoy8lQyuE
SImE3kCRNTtEH+uT8v4IvQ58FoM/1D82NYELPnluR17Ww+47RJBO5vflpbDg
w0tybKbNFl67/fjwtdsVm/dJTHmJzyA+7hC0XmEbVxHsXFciGbP0Fak79LM6
BYdlubqISdlJp+Ac4+cD2mgBTW/vcjnbUEl3D2I1EUo/6b5nkznYsLZcIQRD
dmaUXWmzVheTTR2FeoEldWAO/lc4ooN70aLAto1G8spzkUMR4BkXTR52fZMt
cCUd7KmDPvNbpgWeQ6/F8/w/1FduyQKV8EumF8JrBPD7lNJtSrg/bxIKa6Gg
5OHqb0D1KqmSpuPHKNdgPv6BVc5owG71Aa+i+5dmVRk1bYmak7g1hct/2sSG
OJttVXI9MYAuZ78keZIO0lRycxVmI39PCcb6jG7rgdGHudQM526p1uX0q8YB
gFcfZFlxP1LOSQSqa7ekRj5pJ+9xGo70SJFXYBAb5dm4pJ3kO8Awgb92AQ+z
8uN4UrtDas8lOxU1KgkJBkpuUQm+45QAupG4SigwroRRPqfiJFv/vhReUW/0
Z5EalGPXitkEPe5nG/thKRnK+P/uTvucq9FCAWxzs2dDieMTGCouLOAjV85A
E2iMIKAu6BUENLFTyfKwHjGCHGNrazr1x+a1WgZCC1ACEQk3gq3X2OdQfFjm
F9DTWW7otnZi416hltSOtd4vl9r0HkUOfeDFBmTNOSAbeR2N9v+rCBFiu4Ne
zLxWH0SeQ6teVDzkFS0a/7ODdl63X4XA3KLTeknFoENnGcw+sY3F5g0ERNNC
W0Jr0rHuElNDRNwP6Y2pP21byqXC61KFrfO5PnWF+CA7nKNb3wDjj3IWY8+Z
w/gEors7zpBChfB8G6aL35kiaU0YwccjEnbWcagTIoDFOvJgm3vaxr+wbZbV
CJt2WPosJWSrejY73dmBqRu3ztLocJztokwGQDzTPMsy3ODunTqv0S2kLHa3
jfni8x4C5dkfQ/MokKiD3xRX8rsD0OK/UtU8w+b1BlojqnZfKSU3NoAdYw1t
k+fLU9w6yi02nRr6h83/5dkFlC/Af62JNbgTNo2N/Om9aU+F8kIJkI4P5K8D
JrTdA79q89jJTQZ2P3Ntgfv5oNuhnpfOtA/Bl9Pzs5vmEZvQ207G4ZWaaO+w
SGTAQYrhhzLpDDwgktcieQNQbCZMwI7xquFalt5PZJjbYo3kQD2oPmWFnOTd
B3k8Dkb/PM1F+NNQIEyoX8auVWyTlPDNs0UWxEn8RSLOmV/h8lpeCduI1wia
aQpBkQxgt7VJw6o5hpIXXwsIflpYZrd+ZIzLt707NPA+RY/hOaxIM//F+sv0
ZEi2qbt9AQBKl5crb4mQh/pVyUwGPSRrYZztise5lxpZ32eNsW+hjYTMEDZ6
cFFIuy4HtEYlGwkj1qHirlP/lVBpPloIznUPPGe3oftGs/pWpKkk0KqgcnGz
D1EABkoC+wN9qtYGbXzTRhiTQ/9+smRh7EF7EuBpPz9jn3fSILIcVjL6D16W
BAuGhViahkONX/IOcmQLcesk9Qaa/OKFHTQlbmYOCsDfSrCoEpxAIazli9N2
yGxT3W+a6Etmb3mAuboHTwh++1UgA09fhlNHQANJx/97BYie9Fe6J6mpBS7W
wPJ26Nb41OXF2YW34UWvOl0LDyoikeECrdsHcbT76mr0yaTKMth1/z6zCRsO
SwEngtFGkM4YfWEX+U2FHtjDNlqb3SeEVbGseoCQAWVVsVAc/4Sh7A2VpUdh
oxUEt64K7Saia76osEIExfX4kFj/VRkev8cA2cGmsODNZO2u8uBrMsPo/ahH
xF01eE6d6F90FpvGHW0cEUa8PqtM8EjTEfZab0UC4vG/haZ7gQJ9uo8EekYv
9Itam6mVB1kONhh4U+5wH9okH1sZF0sI5o+SeYMuw2CRtW6fKLzwe7gax9si
T6iL1qkbbAKsNw7pULMxU7GHSngoxZYj3yXf2A+tGJs3TiQNAYUhg6AKykjV
qYZlAFjQhFnmbh6uDmCeBPSsr/dtT61CKht+7L2NNjnR601NhF6qiYPtToqW
AYrzwOm87aeqnfrS/ZkcYeSHL4ri2HJe63cd368kCnh1TBgDHbyARXmV9AHc
HKY+vfoNJA5g3EI/njdG8ClX23F1ROatT3nWriRp/sNUYMHGeG8qMsFIL5B/
jtmeL7RYLHliyMuBFZ9uig3ahQ4mC/WJvKE76u/Es5XGaR5XOb/z1ifxLjal
IeyOCw/MPy41hKTjCez+F8LjL5myTk9LsIywI73/TJKA5g7HsZVkmkDbPtYT
aECcyVYghfeFC3uxYs1Ujln+now7AaRbYO4TjQ5pfkC+Vof9kqMmRrk/gxYk
4p/Zn1v5LTe3Z7HYUZTOpNPmWTV4KdIunM0seQv+HvjGuT3jFr9o1lGyUb/i
J6OC6cVpZmq9wYCtsIJHOsE27rGdW4QuUJ79Ytqg/m2i3Ennduw7htdwxoJe
p8ShLyZGdEVfFOiq1YjVPY6166yR0Pn53HcOarRXAzyJekZg5a66TmULv6Mg
xOMqe/wAS53xuG9PWh6ib2Bnn+RnS2Ew2xRAf0SQXkyDdXTlNTWsR02Tov0y
2jPPf7Z2EVIbR3XSN1bobEgVUSy8F9t3X5YBrLVee3SvFXTK/MCem1HXabXb
xqVw7x7hpzOOUlXU2ztLCIGA6T1+oQ2AhSQ3wEyX0vXJojs6s38Q4uoFqJ9i
p5gkODtS6UXPEvL7q+wRqF44U0igsIzql/v20UHVZ1aEsjIWn/eTl36W6WMn
eR11Ur6dvkw/XM0XhJxyDbp2nhmkpDTIMbsGgU58VIa6GZD9jk9rx3CBVa/o
0KeNj0ebKesYa/ec59OGXIbxcCjpIsCSD/snVp5RnhuycR6wOajfcCrCCVhM
v+PCXdoO6R36SS4QvGTvKbTClYA5RnC+m5Zu8VU3wrYNhbVQ7zk5gv/rv4cO
OJpxDeqrAcOr+RSNWThAtzgUXeslKTTKUZFa5ec1WB7PRxKd+r5EP1vABqVs
gEaL5Susq3jyLcLcaiARE8BGPPk2xPRIHiKDcP0oGhls3z585wzHfWcIrqw7
UZhV72SCooGKtJj9OJjpJ3gX42h7wRUnPOPDZpwVe2feZZRMUnMQ6xMMlglJ
AwZcnx1u8BGllBeLVLj7Qi5z1FRXG8iVL2B95AibYERmiwliCaxy8ykmzHz/
IV4GxBfknYvFkIzxRjziHn81AfZL3PmTHwmzR9cKI7dzeRfqO9bJ+Z+WKBAm
bVQU49SlTREuQGHBGTDQuQkKifM7vM/HEB6XgVQoz3vHizZHZ6jWL8JdjQiV
1Z9D6LTH6j3GWKjNaKGYAvDHOQW0sQKlCZha8y8vszC1mYoYcxNTyhNhzabD
c9g263D+Mn/eVVdruprPikXKVb8Vi1+U+rcWqPf9rc7E22LFl3dvMdr48wvf
+NvTqaWxxsO2kY1SlWvX+f8/sWhm6hyct3iWasWpGBJ9aNLJdnmf0uU5V8oZ
p64qLLDArVu9ToDtPIS2AvcNltbzhRe9lG1JEoYFKmdvKmWSVrumRuoQZFBW
Q8NjKIf60iIqaYY11C3IDL3KzeEyLJ+6v2Ce8LPMQQZ8GM+z2ExtPSO8cmNs
SNe9Y/obzM3Wq/2gsezxxCI3p7vxXxbqPpBJR95e4zI06R2NxfcXG9pPZZ8a
V34eZ+Y8gTdlBGqeGUrCOmUn/kd4twgvnhY1wGsMu5YMml0M3LNHxet+xrlr
ERF8c5trBj6ySwQZ5YOwapOknycvbdGeJcfh/ACwuCpgpdfFpAdOCmAbYStb
VD9/wr6M26C0bBIseylQRasLdvS83KpfFaL50u4SJKagKO2DJl7Q3lR/sn7Z
P3DKxyPIxQjmqGPRM78Mo4w0uY4tVdmRG459UhAr0lnSFTrhSrTRPJTWCipL
0a55HaEq2AQkx60SIWyjnNHMc8BS85OYte7oy3woBSaMFLTSXNqRLODAFFF1
xCUAhZ2/igNL5XRrFCsWRG0QBpiviQmYAWte2S5muz9sLKhqAEMNAdnGc+Bv
FzoxhDgl3I5bBX4sAJVTnm3iGTXNwwmDFmp0mfnm3yro8NmtPknSoNn1wKvo
cBbA38CxF20TOUB4/RHtdtuPF/LNIr5zUyLasCI+Ul9dPd1podgZfwElWWgD
GwpdATRrV0h/Ka55n97tV4j2kXOQ0SkaUrjGHL5w/CdtSbBxhukPGFXajNQv
GMuzUBucQeyprjExVODDa9O6hFXSI5LwYw51N0TBkH1lcMhXf6W9eVTdjBLx
a+SENlU8Y0PxhQWee2S2CaXFDDFOahs6pxb5SQXKJz2DWdVEJHvi3vwZ073n
aJlIpOh2hnyXa0rhO3KpWM/WueJo4ElJJLfenPIvk7XM/dl1KpZHe7ESHniE
LLLA3symDoMb9NRdDY3yd6XgoMNDlKeWSgLZMggwFO7XdEKHe+4PY68Pd1T0
8yzjJD30uZSWz2PvT7OIJpK4wRtL60qUZjIBmwqhqCBdMB+nZoylHO9VhqKe
bYdImjcfAUZzuy9tSXFGt3kKSlbPjAFy30iimZTBRqFoAshczjTnffL4V94c
jGpMlNGICh7AcBSd7hQRDGxJr1KTe26IqMx95D1tX5VgWqnA0LRMhMRkoNZq
fJdD6Gcdi1cKHJZA3gNImYHH3OImKP0qDRAFl7gWlv1ujwzYxICy4GfVOOjc
CLtko5acu3wJds29rE7MXgY90nF42xlypUxLXGmplwBH3T+3NLZYiwuZrqKy
CiebSjegbv+8f35LSq8kiYYcuQFduSWwTiRHj73zSCPHZcx3ansBvI4MOyGk
xNLRFSJJ9g56aBKCuAgwsIbQ4Y3MhRkkCKawNB9dYJQXSz1IvbMSYmQoF/Ch
ghodacg7CMfYcRRGMoXjzgQbds0RX7WBrIFqsju0gHrg8bYRykqBZOxGL8p9
AY5WzgcRguSDO9F3dTpQQ5RfIJTrkd/r0Ib5ipRkkHBN4oA7R+ADX9yY3TsA
Xh4BEPunVuo+3LI1AqJzb1aCu4DFvTbe15ccLBRUjtmMHdiQsXFvmxgExzfW
GvdsU7odG7OoSvddR8wFM0UffLCglZkKweqqBOIC+P3SL6Kgg6dq0cdCe37E
5oP36SY3Y0ZocR9r1JqBcsj/2qjjtNhfQdKgAGFCTCqwgSDfW+6cWcEWpnmI
xxbr9VtKtCipOfeA65kZmeGCJXE+kPxpxiDxUGbAV4NjWZ0301p0OylqgbYP
YDp9EBlricDOkknVITbA+/K4ZfDZ+w6AycBAcgdLR1RAL91lGBCoORN0uZwe
E9gMNrOD/aJA7Kjk1NcJMWl0PbYtKIa0tlmkjQiwo9bKaEBc/QVy87xvGYn/
rzQFEKebg0+k5ZvQyXuwlOj4fyHYl80g/ilcdODBBOCj6tlOBRTlYNI4K4vu
LJPQUD52NRhVYrFdHCXRW+qTcnBfhtgVTgKMUksgYwR7EdnH/uaHL1OcPpo9
5PrL0Nfb3PBKWFHsSBfAvXguyAVhQLt+PcATdQS+dH6uP2KDxIV7B8rO3Er1
Ex+NyQ4STjx5W8Dn+06uU9yCx7Iy2nhBUix33Qh6rio6ShJaXCp7/JIe3x1V
76qM1H2vqX3uVUOvFrg/h7XNcBqKmUNNM8/3sJDgDID0E9sL1Ymm+4qME/JB
Py3EQvl8ufNrqErBb9cBwdtiNebK7sXsi/ygvAK0pq4EuWBHCQM8GIC5G6Cr
a4VjF/dVPNnOFDljb+LTIBdJa7kwquLt+eo0eclUyIhXRHZyKu/3hMWo4Tq0
bwk/jZ66RpI7k7eBDm8k8mushQRqIAaUGmGnkBoeOvqpQog1iEgnMBglb3jo
0ov89SLR7JaR/fSVw8vlGEvMI0MwPrZvnCujPG/Syw9bjNzVue7KgmbUyOfd
WZvCcRReFPTrIgZ7jRnZVamMpjdVKPd587nWnpOvWy2lUZ/R9qrajiBnJnhz
hRI+dZKhm2VeZotIATooGMYhioGAmQ3F/jbqruIvFf5GylKnYRSc0Sn4sNyn
UtGIR0qIcPIK65A/BI4UQASKj4xqBfiEvpdFMxPIEmTsFPNSfN3X94isDRaK
Qp0dBrZlZrCqetfAdFSH1QhzuWdaf72WoAtvonvIstXKu/w+7sAt66X2Q66M
TjAPkU2u9ZHkKTqfCiu5e3sE4B9EN3sBCPhlFnn2EJAVHLJCFV7mkpQpuJYw
nndvfSMuIi8yyC++X7q8AqZVRQSaXBWWUhYiHzxVKCsSnuMapY0p7EmRZiwY
w4jZi3Q5fhrc8+GNIiYNMpWK9DAOtdC1TQMn/ucDqlbGQJczJRMzTaWL072H
QATkkxiEyfy+qLUHt4jQkEJ6d01jf51N/H3/LzW4qJaTS5M6VL7Yfjm3VafT
A2fPUyfs0o10MYOys0UtEtMGmUAHM+v4eQ+n9wnc4DexUFd79ROE9xe2mAX+
kCb77ukUWzJv4sqx2zbBwCxV13Xo0voSTQ71ek+7vvjeH2mfYNpvCcteP3mu
FXsyC8xDy2BRG6jHbPkVTL1DXkiZnkXl/1M7fcwwiJ6pkVXjqsbWP70DYmPh
4Jw3XKXKyFXIwO0Nmy7fEgqtSBZGp7du5YPs+384VVMBdgo/f2XDlVARq3uV
Ye5Lo5vdnGKyhah2H//45TD3p8QQJ8feUwygGulVu7q3EbuO5hItMFlhvhzN
V3UvKSd+3GjxoU5pYSNCWwvo2JE/x9RMKDRkrsPBJ4/ihbkqAKUppM6hzIjH
ZmAoEYxpsI3bd5HGM1QU5fgLFJGJGS9UwCzN893hcBtdlywYidnfOxzTjAIt
w5ls9xfAlF0xOhxmpaSXjZT8IlNoafnAYyOvySsVrpX8OBZWcWNziY1r6Clh
7111YfuwYWPcPvk0aLf4uGViKQmfIO4W0RFghoeMS0F5BxqCT9X10gF7ROBB
Kc+O28rnObuL54k8Ys+0Ky1JGlkvtql3/N1wsN3+aGppWcd2XBRE2rtkk0Zg
Dj2nAIjef/YLstKiDlBI6OS4CyfIViBbtIKSYKeuqD7SR0jNvcNe5WY8GGyB
udupttn/GhS1OkUGHNHJeh17xgy4vN8p4/GFXDk9R2aXWYqzRDbVoiTFq7FE
bkEhFImJO59+948LCpncWxXvgKloKFBZ1mcKv+IfzD+LijZiYqtXIrIthmsY
UB0e32nMDDKgKHb3jV2YlyQK0JwPjd3+6vnKcOAicWV59ej9/TgcdeGBGUoz
ZLFSemwaGi8ZrxZCWNkqf1RNo1JW5a5//MGjia1rNMxlVliKyazbbM48NDcz
9E8rnKezAgcOnacCN4zQkH5MTLtS1GuPV6NIbjGgABZKHXyGXw/mlVGDPFZP
QRbBZ0q7SXPOgShZfmLJT5DjGtai+sECRWDdGwDUIwrD90jmCiTask62LnjI
o3MAYuu2CEW4mQQCqHUYbjwEYsFlvAsOp2Cn2Dn1+U5o6ertGIo55VLf8cms
Bn9UoPWIrSIqXBxnzZkw8X0fQdmBAoXxobsEKjMS2PH4tKIkKw81ontUM4fs
AcE/u25H/PsT8CBWGjGiyjxyF4q35OkgrkrH9KY1phZn0MDsFN6Rj2zihTHD
O3SKAzDQHCz9fvPv3OG++/VNCvb5t0re9S5gSK7AXbxcf79F2Q+REihuyd06
T8hCvLg1HBb4nkemEvRQx2A3xlUG1EfXtVNnbPFklcW42d9+PZyDvKQCW/Iq
mTL8qCW+Pm71XFVlTg7sXYPAO2sprYkUU7e19WmFQuN2dpdvykkOf19lOeJK
gmDDas9iAVklv9gLhY/l8Esl3hMn0ek4oUZUtJUEPGU5Jr9n+LVoB0mPwsXr
m8fUuDOFP+Q4l5aSawTFXEsrlS2vMTiTzzXQshk6T4c4falpT2NkQnDFeDS9
NJj2MbAdgqbL8UGNN2DCAoucFqQMZiMFBw/NfkFqKw17y/217hw7ofH+kb4a
1WX4JEVIrhv5UwTspNESa+5p8ruJc7NpGgMy2pmR8yuIghj1n0jxHCDL8DYl
AjrKX3IdwzrKnZ8mfjvYbcMvgRpQ2TKJEVy8pAHqCdAlSZJ5DAPp8zNZyFdg
5+IvHP3Mpw6qYDSkE6EoLUjnOnr1WzpPvKoeyFt02Rz2fa+kEvcKmTdG5OZi
UfFRorz1wy6tYEgtP42Tp4FO+AzPb3JxYW386c6dUlwu3g9VmAmKi7qyJ47T
CDtmpKCW39ERup3ViJncn60Bd0+x69gpNgimr123i1955PXh00fifL1HQjYl
KkTF3yNF0MeCQE8MLqTr0Atjb2gUNk0T7YN1a7dmmuOgQjwf+6EZcIrxYWjT
IBOJjnur/pWkjcG8Ps3Z5wBC8LCDFofnRYytUSQKwSHbRgqOADQsP7smjlsG
bYSHRgIgRv2HODgcUdMWWfHPxV3AbU4hn0WnF56RiYe49S1dzF7WJuDbZ3Mf
QwnyTqdntwsD41UMa2uGpucQiMqhR3i7hxqh6G/GjJYXE8PUpAkoZgz1XVQp
zQS4Mo6lReUP29mfuRgjjDGmEAEFxhpZ1XR3eR8Ua9muSNjO3byJ1WJRFdg7
MzSswHN0cKT9fDqz1I6AYZNGG0tQrTFl2G6ice8fsKIN7H4syllfVUJISXYe
nzZOv/Jw5Uxofl/X8JqxoTfPO2YMSXNgmLAYlUREvgapaLjAXOW7ZzgbcKnu
YIddE6cJ3U5Qlrak6xLTI5rZbSHYT3A9UgJTeV/DFgyCTGnunwpiTT0Mzs4Q
ywqffvDO4kKc4bCGAtDX5iAJmrJO+AmALf3LVNP2MMgvHXCn8rwBlvVMrvKj
l2tzDo3a/UEqvoXzD+xrUYcp+bWpIS/vSP9ZEefFCYmRWmx62I+i+m2VJ+og
vHNKJksi8rpJePXaFDoxyfI+wRyhx3jHhoEbac+fo04MfwZuxz7xIyMkmGBj
kvosrm3jBuDJB6WmupS/HcXgGTbzffh166NEZKRm5zDRIcnp6Qi6nx19b35C
YpLQNAqYettuq39FJYpUaTcK6fh5xq+UCc0wB6OWYZtk4wzteUImd62S8EBw
wtaNKCmEv0I3a76YrfoNMXKaV2ymrKfsA8UYKnItxpoHcVR2UCcfbCiCacNI
yqXb/aqkIjoZtFmsyinRdu1y6EbjCjWKKhw/Yd/aVqSXo2FBbvOcTXEuSowX
GlvUCHnc1FIYC2marN7YtZL4MQD0D4iAfmFBhHAFS2EMXp2e7Wbx75MsEpij
81ubfxq6ESltJ/DK/iNOenkUlArf0uDxyVHYl5qEvltVtsPA35c5gCaRXSI0
/wFPzNtCrJ6lUNOanrTFBLgQnVR+GVMr5eUT4H2/9Do8yltBnJVeCpGSupjN
pALJxNfgFD1WiDx+fXzbwAe+CimBMjVC06STOzzEwp9k57UeI7SBwi/t4HYN
TD1mI2gm+hGbxZ8ElqHaYB//1fdQlOlUjraZX9OVvvdn+4nU/XjJ7W6Z6n0B
tEY4TyVP+orPi//2HGxpMFzS7EBcgCxOvSzOQXHGl1vuv+b+Y4jLn1xnfFnr
PCpHZ9of7hGRhPiD7b9lNLtQP3jYt5BXCKvyIn7gH5+1KsM5RNtQz+ownTTB
S5ccjm/aX+GdY5UJs1Eum8h2uExVipIptT06aDDPT98uxJJ1WyQRvYVnDpL2
IIxToqCoLr125nULXJUDKlsEPLBHvfhI8UIvz0oJOqixqUKBnx3uw5ZbbIJW
HOSEXDT0durvjQObmMV8g799hTm5IpyXkniKyYtZlwPfVQXkT1oSWgdsb53m
RG8ceQOvsYBIsiUdIGzZLL1fXbmlRhpzt6Pd9FT92WI6H3S9Vd/q66KyIITc
/EABaNXX5CDjDA3ljQT7CZXqjYuyU47Stwa4GvSu+f7sXnn8qIeYW65fOavL
JajF7Nqosp55kZwMTe1YJS3w/U8JVaJVj5oObLLA1TtqvSIpsJ5Oye29qu+0
SO4LomsdrX8tgk5oXURVEFF04Jc7DXlJvMF98gzvlVR1tlKJzcbcvGcMdP2w
cmYnc8R2kTPbw6FFKwdK5t7bvUbqU7F9KlooihvvUuRZjKV2p0ri6aFYrPtS
KqG5V4cQbVnZVeI9BYLfr4PZ/Gb8QIZpc72Cg6bftyS360N02LaKFXGzfdAE
SQCsM9XMXFFvDtBzpIi4B3ryxucSErs/rqCEqqknWzMEZEWr9hTBzGL+1KAb
Rhc2vD0YakbHxKpilzYMVzl6FyTdHXgU1e0W9zYaOClGuZNE3U/viGRP+GT3
ZaTMmApWPGvsb+ijpt4wkEsvtSuw2gu9rhlUzHEOy4jX79aB8F/Xww+IJOO2
k4A4t/exoUVaa8qPKWj1HrrAMOluGpuIiNMKtjjcvUeNWviSNpnN5GqIDmff
8F3i3PFGikrm3svqa52zvjf+a9tQXdvm31E5GQa//Eygo7+O+ySV06R2HaKY
SW6JvZMNrZABmfizOIoVHFJM3dwBaDOJMBXJuYXkXINDLta6QeOjScc30HU7
CMAIY4Sj26N/MTtBY1Zp7G843ZAAwKICmFTiBeyWdPYkk5JbWJIKlNeuxYG9
h1nfmBlaJNBu52LMH4+9vSS0ZUJi+viVtAPlqZeED1yqezEhNJPa9d35jFua
EGUMu41WVHtTLBw8ZgXEig53fyas6B/B58rNGVu74vMc/L3luw7qidm2EnmK
9raWjOOzqwSd/BUlLQs3NxgpfCj0WeQr3Zq8Q/zq1YJRKbyriX83SWbXk9Il
/mk/98lidK5LOjjpvsnf6tg0twCRUL1iY41MS8YFpkrwMem4fmMzFeXnrhl8
KAJfUCxQujiiGEl/+3ruohWXBO9IOVpvPuV94OTrsoMfHQWCVqUvrXriMrTt
FrOcmrlhb2gSlWRygms2eA+D1XK0cVciYcXJ69Z9tOwGiB6TO0FL7yZXJ00D
0/N1+Iw+Z88TIQO+eku44+FVcLthy6+ZIqaqHBC2laXqJY/slne1dTtLZ2NL
0ertga7ibIqy9kaBUe7SvDriI4YvF+3mok1lC2S3lAo3KNqIruI2iKa+2O8n
tuS+XkwvMvao1A7ybzTbuJNREjbJ8DBkR38wjByxB7buFmcrmLSZSNBkBawX
mSuh51YYjEoQJaHMuWdo+0Ku3Rincg0cXEx53wmB+MMdPL72WmxphO/1vCt+
7CmeGZfeAIpAahcoaDz5G6AN1n3fcGjqGSQDsrcPJkT7y9REBWU97a7zP5Rb
gEowLaCP237+Wut+3ihoK3hXro9l0zkjROiqGeK4V03d11hUV2jS/oeGo8Ge
wun1cZW2NRVwN1fQZ6ZP+KkfG5Xn0E9H0St4TAf0TW6JhTtzYavyFdiaIzON
GeqpwHLTRpRrCq9LPKcHT+ozLOD7pQmJ+yV2urCw+vyliDu6kTtnBmRkrrwY
G9mndH1zw2kzfD0ojacPezIT7GdiNxbn/ZGkMYVBnRmn+lGyi7/WEKsUrbH0
/avmTcZS2rm2Qox47jAbeIPJPQzYN2PolZj6XCaBcnvB2zCbGkWWMayAGQde
qX9WtgzJMUNGIYf3vmptu5liPS8+sYP9JyGHoal+yvAt4koEf0vVFUl5tML6
UPuN7Ag6BKBb/nwxmH+OaucOtYVWd9HnVB4VBWhzx0TG/ZX4KiyZFUMkNPzg
+FwtEGk+oM3XwsB7wkJCzJosFvYz37LSz3Z/FXkOI8qWDA7NdyvuDcfAEjkH
kX2XIav3DtbvpjmXb7kB87SW7h0qkoV57INSHWDCvW+a0/3tyPbRHx7mEO60
UQO8uaRagEg4keMfxzGi0laiFlsyoJTdPhugBdAN0EFsrWrkoQtH6SwzuJcH
UmQKVEwTeKPc6fDtfSygB2Qahx0brY7ftQWohjXZtP2e+5kCs3eC+x0IY3vE
FaS2Pywq7cFqCcWujTQhYHXELUUn6AQi50UdHTlqhj1G1NI5gcCIV2CuARWy
AmRZoyWCWiIVzyXYMq8SmeAUrsDhQY5vsxKBfhNHNYke/TN++Uk7DY/Z8dn+
uq0npL9gAzB2eJBDW8oZ9FLELts0a6WIXnz15AKNFL0gQaKZA+SRXfMugK0Z
8Xp/ExFVLwIcTPQjhzIaoB+x/XTv+8cyoG3cYkyvuU1AnshfuSgp+Jbh8JfF
M6CUGzO9xn2cQiOQ/943cj3n3O+BZHkfbdms1oAFtvK6x0p6dHCpoiHhhDFf
sk+mbJdhW4l0Zs8ses3i+7r2gqcy0YcxZN1MEZ0TIOIqiaQERJOssNizoeUc
7da0fC49NHk0J47pEs6xU5WVwZ69S52MOmqEIJOGHw0k8eI18JWtHfUYI44K
Bw0fbcd3XnLayr8tO6trtgrdln/7ngb6eRq/xR6xQR7zPAoUyUHdIbuoU7ce
HivUZZLsXjqd8kVliim2+0ba5noTt9GHDqfWZOK8vdJfu5W30wm6iyeoi9Yn
q3sF9D1yYYCZEQoAnvybAIBqhFc3eZT1mVur4kRU4kdhNJIZv/FwwT/8U0/q
O7q+InlQMVUGVltNpsQAYdXqgY2/ao+JWP8yLv/JL8DIiQ2SxM7FFEN9svrz
RWJgld/ibuqNxWGCYenBkWV2FLHDyBDgoDnb++Gf7gAjBrDlYi/mGtjzX9D8
uZUT4JSDWEqy0+hSNxLy6zQb+RNBJmr6bICANHNXQh7ROtX5M+3UsuDR4a53
K0g7O33AFTwOPCYtIH5i95uLQBw/SB5KWT4z0/6n/93IBmoKYAYq3x8ruKIF
H5bdLponCdpu0EA+ys2ffXO7tEf3dClSo+Z1fKY5akHVrLHfViLkJMSC5oWI
MOf+Qcus+IKJ8LUtC5x1O0bVKcXL1+Pv4y67suxYi5jmeQ0Hgkas7R/0wjK1
wa8yev2NQzDAAUQ8lwtZRh8DguP9y1eM3yNN4me6NER+J3alTIimplKJ2Zfd
kwkm04f5DKvIa8tVXbEYVwn+2w7xsvzeveZJdrj/SLNRVsz5OthqQBjrwICG
5iR4zOajbvTxwy2P65AX/Y+EGhGVENciC+Jzsrf8944Yx8CNPUBd0xvTdit6
/afGtczTxELDT7rZmR5a82HUOL9Oww1EzMf6RLKBVibQX4k+P6YU3RNrS5TW
t5edu+jW67HEj2jMGfIfg2C5NGY3YN30bMvb1OT74MWJaUYYwQmMjg1327u5
zx9cgEdwue8kmJQBnolKrglXxS1orEqIy6bAMf1F75OOhkvUe69yY/YSNJce
a6i8FoOo/9lgkvfd6ZiGufDjtLRfG8ZQtz48lrUIEo6G7UL0puzwvOYvDpHU
Ll58AJmWf5Kf93261K8HPwWwuTk22Yl6EJuoGwj3F/wsdLviSHSZhN2XmBXM
htoTJz4lLk5EBqhU4VH6SsTtLWh7ZuN7urTD3TamzLBHpxIQFVsAILxrOCmP
HZ4q9r8u2E510rDt8v7ugTJ815RrraqQ3EyJ0yC9j8W/W1ZfKBo28n4K8DvT
r71vnHxOIEzM+x0dXT23AeNFb0LExSmu061YtA1tig0+t7X7nO26tEuzF4GI
Mem6vcttNRrW5SkGT+BAY4uCvmyGfqimDW6rjPBA+Cc7uVv/BoDi14NWS+6K
Nqh3s0OXdUsxYNOWHN2jemujJB4U9C3BM7kb9ACUo91/B5jFQJU1bGtEjC85
5FCO4D8rrgAQylmw4mpiO9oKp+EYJm7hxJ9XGwLznpksT1kLu0G85hGC0fXn
fCaJp+Jhc68qZgN+f3jLxAV+zesOzx6HAYENbJYrCBk85WWm1BpMbCgl6K9o
H8UAaT5RndOT2oL74UdoTUfxZs9XcybNqUzs2ivTZVAS9SWIVcCCwIfUCfro
P9DMKsu/c/cMrIPjlqG3EqBcIVvASBAvhiub9ivnLSBFZZ2yJbNV3Czh3a/v
yPlHir61l88KMM0Bc8eRjlwhP8IFBBsS5h0GuVgMwEb4aGnEAR67vR1q/CV0
AdbTTXPcel30Rn7HsE5OBSRn2F2/yJxXfzQcZO41vMH5FoEBDaVEJaxLSnpu
oR0MK/grpuGytk6wP5yUK/FxfkBhHpFlrz6LQQ1KnHE5E85NIoLvc/2EtSyg
Hgw8tTmmn1DVheTDvI0Zilc/uGsT5ocKgAzaralPXJmrgnjD9OtQWuKY7suJ
gLzwv3Mts/mKfxGnjAEtL3k5c1lo7/3kYw63Y+1yXJ5FjyEZDM/3ZUHTj5NU
daQsCRiLl9Wdjhg0Q1kqHZjRWy1XaflnIXfiKD+NCHEFUDJGt/2fkN3p15gM
ROu8N5dttwHUwd32zoDKd1pu88mCACGIeO0j6rgBbqhpEFQm+doFqzDlbscm
wIpq35DxqztjfkpvBUVrwhM9aiOCcZmVNfKkNqcxmEvhYEAn+fspC2gdM/E5
nishWVOjxRgvQWLqyp8JKvAyB9mgtAWWBXOfwFX3bTuq7NgG3/vlQVMu3Nx8
tTusDyMEo8H4xhDBNO6Q5jI40FigbmP4r4X5UMf7aXjfNrSchc1pNrziTRUz
hqMqeRNdt+7j/hROmTdVVzzsTLCb/DQESwomtkvClgQ836sZsq563D54ODRy
D/5TiAkP1hli84UmTejWgyqKzAs2WhNq/npFQhM8xFxbH9We98P6/ockt87J
ID9IptK3ZOBxbCOKGAe/Rvk6IoQhrrCSP2oNxlAdTrAN8IuEw3SNYE1haYC+
PRd2pzsyyxqCDCsjB5wLPdL4hLkre5mhMpOMfzLD3wcnIQt3ZfcF5pA4GMP6
j7C2T8pV18MkxvsFNYCMPXDRwkPCWFO/r7MdBNG1J/tM/HM1Kc5NBgEZjZap
VzeRk2fabCwW3ThR31difWsLqA5h0algQkEQItCDVjwDwzAFv0lenxsGWWE3
rFTl81UhSY8j56a1X5+mJXH7y/kjzthQ4ljw1fkxEOYd3wncHTOjnKhPjDde
FU/BtGmhHlgEHwd5qgCk09GZmSEVNxy+PrDn0mn9pfdvA5gQJR7QP9PLZulZ
FemnX5C65IsKD+6yZN1Pjnq0ZnKXGk0zNPmoXj69oRTo5FYbwYb5MeIiR72m
wrH/BVdC+W66D2DV9fEmcY473hK1VT62/i5mCAl4iPuCufqflszG/eAiEp6T
4w79rxXR5DEkTkhVyTL3aK8tlceolxNLj2HODVAzECyKJ7o+dE5WcDXsOlsV
hTE4nfw/C2Yczc4BxKOQOxdnwK7Vwy0IhoMXYeJq2tunvucDcCbB/wXWmhtV
Xh06BtKMks2EDZw97F+SJ+0wjHh7JrAZ05jr5C7XMV+SHm0tN6PFzYUhXG+Y
WYBgxGYrFa2f6v+1cUPzxZpUHsM+PZLBhWNpMCCCEcBAqgCQ4dGFtpJ3aHbC
kufCQuHeCz/oGqPQiUyQKdHUzoidPZUXthg3tGBdt1WiRXorekk+e2NpmtZx
EwpycmJ0ck33clDm+aydXlCcAqxx/mLMdIOfkzwWAzXlGk2SokJE7q9Bkg6K
mDeckAypSmTXnxERTQGIBnUKWMlKW/AXyVD5XviY/7ANaHYsmyOywmDLcF8P
+YXA3vPKGufb1c00o4UrgVU8uy3nBETwdBJMtRoTSmIjU5iN4zhF8OvIJcIi
R2NwyxP0uhdzK0aL8cSoiWl9v25+OHXFncuIZb05GEINg+JyidS0uAaKMQVz
EfKbMLITEZYMpVmITgTG+fmeM3ukhU/MoiGSTE9ANek0Wj3XFTN7O0Iiqnmt
1le4vjVdnSPv+lR1YH2a5Bdg97n0/FbZSstnMcFuksAMXTKyR7oHONgvruzu
zA9sykEGtpkVYo+WHzCs4CIum2uutj+10DNA1v2dj2E+2XD/6hPuG1Zre3Az
y5DNj/SCpIOGLvK30uxuVRV22mU+eqNkvKhcGIxlSxi0vXXg01aqJHNC5DJm
elb2pgPnQJVH7jXdvivM1eaypComB5hKH8GUInKcumi9Ub+JQdXDiPE/K5Z0
jDsUZlF4rJcTcTzOqeBlohmnkidxNZgeOoLXTKF7wab/sp5yHS7ZW+89oNdZ
/w3hZQRhLvqv30ZUbdjOPm7XE32ZTXKwiHN1M1nSSG8BFccfusbLQdI8zFon
3lbwEYHPlz1GAD/acjcHKNGMti+ZOp1dv5WKxF9XgM4vWvOMWC7otlg9yS8D
zPkj2Rtuh/if7sCwHK+2Y8pG01adKxWoKUW+q3/mcTKPI5JJ/smkXndaoYoZ
l8GqaqYvqDIGxL5nbmGW09Zke7XRbF9jiGChjFIIbqq5+egKuQ2KO4kDZ64T
p4n3M8ctNXl5snOqDfz7+HUxZyTuNS3dAb2HPE6VwxNKa0uganRXgb5RSlcX
x4LSZXTKmPSctS6d7ZB2DT9ojBb6FhXaHwCjLtHlm+tU10uair6Lw7EQTCh1
lJyN05UjtQHc4aqpb1IuRoA5vq+CB2XJ5tH8B9wCbpogaV3qD3/NXhJ7Sk92
7eQoExd6nVMMIFATg82DZP1zLEft8oRfYBZk0/qZHuLP2QUravS7YL2mSzIx
1KPP7kUr5OPCwA9tOZryH/ywk2AxRC3uLiBvqMb9TIgGb4xd7KMUB3WaiTy2
B1Ozu2KR4hepxWeviuK9epEmfG5th5pb1S16F1jI2Awu63OUYcNGM9rSlDqV
QhGiUWCpQdbaIu1mLPiCpbpEWnrZoM3mEunHq6CWqCVJcHH31SeomdcjGLvz
Lrg3HyT9Y0cAbGX/8kJonp5zaG0cHCb+PKr3cAkpc1/5cloDcx/1qsMGyFzm
MbDHejPUpLbjWo7VKyafOsAGWPDsL9fY53f3M0gkZfRqtpYVhNpIn1yAIXIC
QIV475IY0vhXJz22hPo3lhtFajTzfG4K74xuKqDZyo0Iuswa2Wj7TJuuv/wQ
SP5OjnO9kxkuu0Siun6YYBLw7YdslTreYZod6yUGlscQykVgTUuXFolAENsx
kYagNNn+BXKDQlaOe69KY7NQeWWf0vAV0dBi1u5cq+Axeo5QC9ZVM7HaOyiP
JIn3wyl9CvkFHvZehVfy3P0XH1llNZLV6GCTFHAgWJGM+9WImfS7WI0GCA1a
en0niyUARCjj+8kV52iCYJzQpSGcgFTeJEuqDrY9LRab6PjyHBs9YSjo2dOg
m6MqEjg3MtQyjJUxCfXzyyHQQp4S/95dJIVY12QtHvr0a5QZOdxheDnqe0rV
bfnCsbSKtWcn54/UbXYUrpxLbKBlUGgHwcxQwN/BpQQJsbZ4ZmOaobetD/yl
Z7wV5gTmtCJtul7lX4Bk4tfJdkt6RsMWUS1iwKxoxp2uwRY17HSzvCiu2UxK
dRpU/kTlJIKrSpmHqkEHfeCnoilWyzlSqGH8iaZAtnyAobR2txU4PfSSMhSA
lbw7ldsM4XxUAm8U9ZmoRoz2bGXOmnYT2mk20QuszI7yzQmfhbvBw9Jp1OtF
2M65jm3b1W7DOw5C3TNYHrO2cW4evwBfP/kV1yUd9xiYZx62GQTroaI2+Ag7
vdiR/LOfptJm0Yv2npqW9A0vzL5kS7ukzAVd+fDBRKfxuUicF+LjZT+DrJg5
Va79RnGVR7OTV59MSA5XcxT3qWhITatf+ipv1rvVL5QxYVDQqXxPGwG33C9o
I88WEsn+qgzIyLLwhshqVAwwpJFXeSJjtLv489HDsodVTzk30hZxlqM36bQN
W7B8VfaXVriwp18wULL/UYCTcevNO0BeLbS0276gTOei3OCZiI00nofAuyQJ
hIJf/M7m0kYOospLU5q5DSXGMewH925PHC0QigQkqb4Aigtsdy0NwhOCZXTv
L6kQobMcXsO3KOTVJUo7C4WgrdfkOHMh4oGf1LALiwSPuje0itmCYeCqwqRS
XOjGAfVAgt+7BVV+SNJrauNHe/3pQo+9m5e2VNNI1dLyTxUcXwXP8mXoXBuv
oL3qXzqytD3ufRmUIxR5cTGFC6oihDHuOjSy+cwpDHo+efENkVKGG9W1spja
yU0tF0YhHfNNdjHo+stPmAc/LCqmiqOOS/YzDN2YMvxEjseHlgk3Zzw0eWsr
BHFnqGXlV36pjN/KYEzfu5H+MSLgvE/icqJ3SPnyGObPu/8Ib7eWMBsrs85i
qyI4/vDMI3Y0JInqIKwx+pqXP43eBcj5Np5IQfLko6Axv2bhu+5x8OjP/MY3
/ATXJKqwTqI/fsZ+of5ik7MTfxX9pcM9OT6rmczprOsuySKD9cRMSsavhN/s
1T2+q8h7zL78um9MAB4fEQ0ksKfWjwSZBlekXXjCMTIPqv2JrqSLUIWhgzD5
efHOoTGPH+I94OX3XiD7k6FAA89Fu02Cnowg/Zo1O61k0/itFzEbdtxrzaKr
MFu4tLSyl86N9xP8nth8P2ppmxHhsY+6FamlhbhrqtorIRAWF8EqA6VN8nFC
Pmiu0USI5Sa/akRWtd1WpgYC3bja1FVJs0NYJtZWoP33p3ZLDOpdxc9uXyyi
dwnrzVPjIh5tBsWen4TDPICfPBxVtPk0llVWyurll5f8WVIsf3FvD2vMMLt7
hLT307LxCHg1dysECFw/DaVE++Da9tRjBZPJNMaUXZwgoTguxo87Xg9eLReN
+oSHF+wDzfTb+026XqGk4o109yd1UHbY89QrgPsVnCZ5U+Fpluy8uPqUDu2I
fXOfF3quk0+yR9RPBSIbSaRoxcLAXiL0dkfmKBc2JSVw0wd07PCXxg5HF4iX
gfEbrzc9tDZDHhExixcKFMbEXbgm1QI1JpmFOro3O1bBsg6WvK8hkSpL/IiN
LkRah1wykTalUU9s0yXfE2yGnp7JejEkb6f2QQHLvAZo373UE4wOwPK4bRlH
aST7b5z7BnQjIv/9oLxL4b9aUXRFps4B49rKp6DShCq/B9uLVuOi+Bj3pbwo
qJlXRroVKZYpRNGxSpOi60KPRHDbZGrxKgkp6UTXtpQEJdpV+QNBr3f0qW2O
5zdr4x/W4TLAzkEyA2xBVBKXBZufcmbXdQgm1l2i01IUWKKUwnFqnnrrLsu5
FDmRDEx4XqoiIE3mtVJgjNk/nZIKmI/LUBKorusbPyD9AWnBQnjZuoLvPXC0
tGZah4rAsdndEBzYzNpu1KAK/vBK+rDASa8eGhJOMnLbwOvZiMfGHf1Grto0
iY1tbvDSpBe4fNRPLN0htWjFTesRhvEwKM3Rnxa8cE4Q6OvRKoOqOkbJFDMB
PnO9gV+gQBP+STDkDIfPF8JMVsyCWKF7MIP1Ojc9I8oteszmjty8Cb+cICKx
7Wtbra4jscKghGJ1b9tZt5rSpH0CGCGGf3RTNY0yCn1up/ojFS535OBSQWY3
hlWKtd5IV/kZaDGntBppSCQCdHKF9vz2AOZv3mYPNinESa1cwRNveBWhfmgZ
P6udVcb6oTBEBdty1xosJ1fVku2UO9YRgtPlqv3T3wFLG7MPE8P1FO2FRmmt
z2Aq7cm+ZqtYZqjR3quxUARyA1xn95SCx7sS8jcyBEy/fwyaADetdDmqgECk
jaUZHQXexIhJQm32ThibcD8DbFBNdNklIjfo7d/if1idvnDnEGYiBOSLWLkJ
nC9W+86GCBN4YHlF36nnJDd0OqH87cxP4NASJr+LqB7b19gs/4G3GmmEPjvb
Xh1T79duvNt8OPCawScgI91YX91y5dC6wnRHI3cC8vX24hji3pOtnFxf6QBg
eETIX1afvMJaeLfW2s2sQl4Q6JAwhDjxGdexwT2xoD1nSgvMFP2fAm5jKTGs
hGkdgYuDIA2CD+Ido+WgW00mS9EZv/0shHIOedvXUhDPn0HlqRYa7VjX3SJz
ESJFRzoKhPbzSdxFvbPQPaPK2NYhVyfVCjSAN6TpAw1LqwqOUf1+qBOY3ygm
Nl+knly0qGqlAq/gfte1U0k1rjBlvR131Og9HRWP5zdDAlW5XrGYa+oriRAA
fH8Vi+TzqseT0g9WjCkUZZfW8wY6GBUD1AODeO4qR8aLRVsB8YJSvB3GRxkb
8N1gUF9Aaw9eJisNTf9Am3pF8zQDZ9PbHljSFXnXA2Vb6hGeoWFwkzVH7mEP
UnFyiletynZwR8nhIhpIZa3Rsl9xIe57Uq9PE86gE4A1/hbETB427f7yhlU/
woZaV7weARtjjS8Ap43WsC52ULxuaYw1ChpTi0JUH+zBKjaA0yNOrvkwGf7G
7FsZBg0zQyh/MzAT1pl/GYE5U07aLWThaiasheeiFJAb3AkdgbT+6YsVTgi8
9vQrSczFFJsPujmyvEQBPm6LbOEAGG/V8L7qr64IvhgCHmo6WjwFVU3SQTLm
45H2dzUn+2Bk278OGE7ZaBOIs5TEtvfq9mhshk/mYRYPyF+XupxApAeIJvPo
kl2rgHi04OE0GY3Nf0s/C0bj/15s7/owA7ZALKWbvyN9EoQf66M1wqyEwtdZ
ybD8Wp+gg8IRYvoZTtZpT2ExyfnIQhzWAXJExy/wxzt7R+2pyaIFQPLoL90e
cxtKqRMzbk19DAobWAsaiqP7wjkFEPUo4w7y1XA9yONAllt83khdwnBYoJgg
XSRmU0gVyXUfDP+e0GekXlQPcjy4O3MH9cDI4DAQyerwOmZOdvHDhoRdSfWB
2fi+91mOGTcxS7ZxTrQD1c1anCJnyz7YxJ8oRCCgvyEp13x+oEbtPDd0AwXP
h7Rn0eKUgBxCWCs6xnbn0dMJCh1SgW47qaQNDHmxNW/1xCH/eqQwNoBAaKYO
o062+vS473DiGO/lcXpwf29bQLk9rGo8nwMxKYwn0cGDR3/D0oyVYbZltZXf
cz1m+tscjq3oQh44hnOgWx0rBxaR/rikma0lhXGXDf7C+po1dkxd9ujgV7M7
+wF5JUGw+EcfUsg77XtEsyvM2/9MDLel332Wn28Bl1fqN73wBylxBoWEAuSn
8cj19Fbl3rqX3mWgnHEPgX7oig1b5aqjZxf+7LpI/6WohstfmsIb/4tpFh3o
YMnqvcTTT4lWFWCTvgoMXY9aWBhQWUNKdan2scorCUV1upaK166H5MigVgRY
9oOVjWbbGqVX+K47aoj4WzCFVY2Sdo5i7hp+eHPfXK0Q7rdJDAMuUn859V1J
fZYTjd18jXl1GFwsVB0Lq0YtC/u6epUua93SsfdUEzBNZV1IKqfQcTHfm3F2
DeYR18bEzLqFq16AiqDQJI1AAFBsfv8Gz2EdzP0NFTdPIeT1i8ZvFchZimwI
eaZyOk9JCfIDpwDQw+YzXZVMvfgWYyD6nGVBZjGyocyU9X0sUAmU38IqplrS
+hfnkeQtSORbTJ763jSxQZjh2j4WvOTFlck9nptOoJ8w2rhhgbjgjiuF5Sp6
tU9PTwBeJRbogiF3dO9GFng8ET7pJS9J/4jk5lV8Yri5DAUeN13mlX5rXTc+
qYeZEcV14rQ/WviLlnT1OWcNIMS+bWHaMd+b4RfuWt4D9QiTcVnFWiTibgMV
jFH3YQksq6Fobr7eDqKusEbMX2aPJjoG4oWZRAjooKPv469Z836FhV36kwnu
AYhKM4DDmPupQmJbYBZTR8R09lkuEeVCqFZNFWor33KIRkdHYP9Y1s+x0zYG
MBzFzR3elzRzqbfRfqIExHrs0LPxbYIpZsUkKXDd6xHWBWprvm8yW1+da1E4
OqI5rfBj0RbcUxYNMJ/xfChUu742nUo9zJyZf6xWXi3JnqPgoRfi0OfNdaJf
A+nNW8l9bFozjeFE1td8WjPdQvKYoC6xbG3l37d2jDPu5MqfObilYY4+gh7k
SVnpPrQSzSiSTq9DFKHERqWv53ozY4IOA9mvAtMYFD5dNskHhj8JWpqh0gul
xm7994rLeCv4oB191aDGiYa+0y6+blVv17WQslrTWcqayeJCl6cqvOiST4oo
+WrmM5zoQcLpfxdunbaWPiUtAFEZ0JHYFJ1k4Ozc3KNW+AB5X4GsDiQPGPvb
29y1c/kETPyicA2cpxUjihf+dtGU2MXzMPu1/LtFhz3CNFaQvT8KswuKnP6y
Hy5Cebo1/tccZS0Wd97Loo+M4CcKbpvr4iVCOvqBe2WtXToXvthX1vdAgWjV
IEdn/LYFJwfraya5quxAhjuJRTFaUGRnZ+mHlVdQ+cFnGmP2BUOKF4i+YRlL
oMDd4XI39iB3SX6JqjwVQPH50+D8/JYTripO+fRGREVoubwJph/5p1rRMBk1
Ztzl5LzUh4nAFuw3AOwKpCysjSc1xgdMm2zjAcut20jFNKFlf1gjyLsNlAYa
kPKBBffy5S6epbhOlK5WVN+wgHQJDSQfp33CHPgv45UHfdW/8a9/M5DoaAGY
4zG3reM+WZmI2UcY98KYXWekHHX7KC2I67c3840UPmTCQUvF3fFl9xioqAig
eJGe3j+9UHVLPVOOn6EZyEzHXK5Q0/X4veg1bJB5qgDl05Nz6I2wuK8E/RBo
YJnSqEb9msTkDClbeJi01f8dWFPKpDMBnxaLPjrv5UqMVMJ/NtQ6GjwxHIhp
V4SFbCNBdsTDqHINRUVCL0FVl82Sgs4+mj3io4Z9LhreDsQxyV9J9sCgLrRj
Qc23SnR7c9zc51a2eMhHCBC3Q9baQGJbr8NS1KtB6AiHtfeWRzsCNoG6vNaR
6W8kXND06q0nndzF9nxh0M2NGUEUNGr/rnNzZScyivaIFZvenEf6o2sSiOQE
x5e9h861bQZfkIjJudtJ4iH41HLKT/KJ8DP9yAfLgS1WC5MOMljpnWLzWnCN
HhVi5oZY1egFMNiranJDISMzATJKFmF/X/QddTmuzuJ9xXp4ErfCXabyFYri
NQX1xbFq5wn97DHOdF9+phYwQSwXL/JvLDUT7hOFU0sk/6qZWMu0+19SC2Kd
zDMfIYFc3FeQb5ghrMAu1sDNwJo4x0pGlUpLFqi8ZieaMAl3jWUoTmDl8S4P
HUU9CPrppE/GsZfej2IfoGIaB/jW8u44ouS1ni8PF7KHJABaFkJh6l0lHaYK
WcwyBZ7STaJqIz+bzlweBznrrC7zb6NxPsGQKfqmhDSNzmzIiqgSs3UK3c6z
HojR63A1AcQeui2NNYI7c3+Y5DX1j+sDrDMW4EtPLCqpyJC1+xsv+TPqy3dS
XfEwsdZKpNUJLXEEWkNL1PnjcaqI50blLEnTe/W28/YmDWNxCvQfkioJRAVM
eEiZVR7Wnh/1GuUG4NxFuMVfX/zFrzAKMBKBH8ucx43+eQN0RXudAYZbOn/L
yDfZWUI0VhdtdYIACTSRE8XDpnYk9MZW6nUJib9UEIBzkL3a2ZzFbtCl4D34
wMhbmBW+qSOd8tn+29w33/a/eyRxJ40ZSdpdVt8uttQAZSOh2n6OgX5lvWFf
YJjKJ4xf4nv8CDiGg7wfBHqeKnH7WDiHgHgosawpSA8BG+2Th4Uyocb+37q7
0BzTzYf8le3S2E90IPVshaZGpxDwwfJQF0TrcRNn1ypu/YgO2GqtFfjN08R4
HUHGqVjBSc25oddeMgpNSNfacund1nkoEYB5RX2A/nEY69YXiM7gn/7hBZh6
HSK8xnvZ8TSFkK3oF8Or5w0wSGRiB9aAzWRwt1a1BWPPiuOiF+bmP1Sr/Ts7
qqM4xW+Ox0D99Y+TY9B4RUYbOVfhWUrW9JjB0BSBQMnuEP9CAJLxF4FNQIQR
YA1oOI+aXjtkMZLt2KvFqWKo0femeWLOh59Ankb7FQaea98npsB5j8tPxhWD
EdIWNN/ohqXaRQBM8Tp+us0CPNU/VeDKVfwC722iIlrlqN0BzeuZZUimimkt
pAyffIwPmm5hq/1FQtA3AcNSuXPL2vCPgl4ICtZXrnR2U/Qef9lh+ryWhEBe
XpDIHl2inV5l00osRLCOJQENo9XhZfkwLwO2bpUuDr97u8MQlWiPxQj2bVQd
6/BRJYj6/A2V9xy4sAvpMsK2QcjM5/KCeW/iNxP0MZbhux8iD3pR0tItIM/0
7OmzoUL9cCpoeRmCSxN3zKBsov9unkTgYP8E5eq4iMXmE5+26FrVS5D9KAp5
QoX11M/hy3wOj0Y2pfN563wjGsmIveX9OAP+r+CikAZYHVNfG9jFuB6Q1Ue3
+Vy8KhgCGoqs0ArsrW2vHnJpayXxhSBsIXrz89zLqPl3m1KqSSgj6g/VnQ05
570MbLWDlXHF1q4iBF6WE5+im+lbe7fZgJNskQ4/QMeEczrbdXF3nYkXJIIE
BvQLsHbThNM9DNSe3LapV8w3OyXjzTvjXg7N4W4ziyjS5DsCmaDMQVngL6wr
5AjwpYP8V7pANVxHv0SCvtiTBQp9QM6rROMeyk93S3bhm+EYpo9MuABbaxNa
45/LjQ2NO16OTXXEJqZpdJfitLvp9MsRXdcRWD25dZ9Q+jBHJ/zGyo0kMd/M
ZZE55JzWOa26JYySN8Ex0Sjc1XE3YOX7Vz9mEETdM0l0h3cxFw3dz2S58aSJ
9Fgd6ABgc//xWsaj3EpP3fdodKMYzHSIt4iy93JC8zE8IhvBgJZAColPSwk7
RR9Y2zUWF5rxT1NaekHb+YvhI7Tvl2e5McSAUsz/xpGVy6p4o+K+se1Ekoi3
xUelcnWmyGlDRtEMTVWe82rCyMiM1JWlV9mBmF9iurF0soYoaw6bL6QLUKPZ
nJYFX7FgBv7AIPmdlx6ChM5Ch5mx1Ld83ZVlbCR/ZctpfY7ohWqkmJdDtZom
uYDiEvyYsSc06QYZ+laERV1jDTZLLguAW3x/Y+/xQEzLxRpY/XfPqljCa2/U
dvfQWHi/AtTeUzvKXY5IdBtARV1yf72HWny1SSwO8i/sePM6hyX+NdhiZW5z
5QWd/axYlb70EiO4uJtqvfk/mNdOvOaEcR88DuRYtnSMV2muoJRuI0kU6MOj
1g1ignHFhYiI0WeJE51IaCkdtDaYtlT6iwvxO4NRmAACd9n9CXwBwvTuvRIO
H2/1k7WJsjnW6FrNWGLLIo6nSIMJiy16WD8fW1f4JvzsP+ibCRB5Oj7t2QHB
LPKXBi8E7Jo76DLoO91wj5iyEyj9mH4OJKvRK/G4/P9wQnzGBOWfgjlB8xWq
ZQvs401zSDlFCYXlll+lY9IvjA2P6gVrpC7VjQ6ynK3RWLrVx+rJz7yM3II9
TO2k37U4PBZc6xba3PIs+KgAPoRIogzDrTEmKlCwoRG3As0WIiYWr1yc4QFq
uemWwRzPyxYnL8vXpYCvZv63giWc59Im5b++5uQMo+5q/4k4e+uYSV9TOTtv
VfMz6rXSUQQM9cGdKdCa9CFpp9pUqpu2LwDz6lZ5b1PLU+5r8I+2HPOAgbel
t0ouPRK6JUS7CHB0wYDlqmJPetb40CCoooneY7uw0VTj74pUUJMe7WgvJ3u3
VgQCu8RO77tMmEZDQ0IjsW6+uG4eWLpEy6rQEzKZh79bsYMMsPvc56iZrI+I
9aUCMCrFLs+zZzRXHd/vzj8H7sKwoBKN0Ic6/xwcjiYuBjwPJ+KvauOHZJ1o
6WGieiM/qmZrsavmdx7VIxI1WQ3nh20752jbLtv29wf/qyzJSD6J19lIf3la
lVj1KpzKBEANqDHCKwOK26SZr+tvRducziJV6s2637myTeDSy72lnNBswWEq
1abmx2X8W6w0MpDXY8rqHwLfnZ/fbim2dsK5uVj13wtfIo9Fg1JrGoWDks3d
l6BEqzQlDBGFS3IsgeAAdNWXGZprkdV9Fd4pRz/4yNa2nzCynYiTLLV+JBH5
N1HTNJOQhmIrNpNPc3x/8Wj23FUcGmP2VY5EFWrJXRPU1PFLP3FgU5Z8Wdlk
YgY82bRGCkbQ6lCpkvAxB9nMyqI53kxvvXWcB2Up3ETbVbOigSeCvPBMCBxI
drIZO4UgAVSk0gmAg2xN6whtvfeJmHs0P8GLv7d2fWJib9HoB90/j4fIFMLf
xKwsnsKNaDj/oiN0wDELSgt45gKeQAx3Typ3TOwP786J6DiEeXvkW4EyTs6v
PEvhNMXjPMsMUg7SvbqCEBMt7l+tZrrUSl2jLojNJajQWJ/o+BoXGMGep4+N
+EGggkXzCEabAVLVlPjwMm2Ew2DAi4c+n4AMA5obTbPzRqblHjcXRA6a/6Rw
LCIbDbeW6yeZErvCfJIH7BJupaRf0v+MLZXGE3KRW68D5lSoHloDNkshOdNB
CsGfFoQnHqv5DaKXJuNtPjF8qWxE9hDUDPvNHE3YL7sHrAIrxgts9bthAtZg
6Oq8sALQyafhroR6At2gcGGGCMQOKH+AHb/uu7LP8bcWbrws2GkRNUmizQGw
h81Gnc7LQrgbbKqwjC9xxNVepLokHzfhfNBge5FySZizBwM9wuurCD9rMEjl
pU6bwhiubp/mzkyLezeicQzO58NSX90uNnlW3pK0BSynU5sGpNvNSrwjCoje
zs1iM1aCom1MhEG7cQZpShl9eO2JwlglkGu0k5Ghn/8UQnnEg/2iODJpVAFv
zBIWbhipLIeDLIBEiUs+2R/v0NSOTGhYqTBWCclsZCwRw5cwUwkNoUwvznKd
AeBEhmmujlpIt5W33V/8QWadJq542Lpzbt+/VW48st+gG7gaTSPfF3Yh+V2a
hlQDCiRkzESlLY2h7G8OkhNZ/nrZAM1kPR+VMBJxBI9R65BLul0b27qe/Uj5
KSM47LuzcxpWZpe5bB93uUxnocy9ATsw8/at4c7DAVssNGz7fzVLBJUv8X64
CyngLkqIWD7XThwaGkFW30iM1HLMquI6X0bR1GVVMKshnFGSqkk1nphcVk6A
1//6q/D4COhA0udVKuP0LTUGfuJNIhGj5aqAOFHzQliJrloLM0KBbd1uIsJQ
Pj1OFDVZyiEc9ystRnMcqJeEpCzKoGbR+Xz34CjmrDhmYjtFNONjbQ4MpkBS
GTPRENoJQgl3BFIfsd0fyF4Mej/aOtKi8/HgunGs4j0WucIRzPUwHHKkZ8Ng
jS6yDIgKaFNjm3o8f9oeGn8e6ALJ1M8KiqJhyjQXefB79vJJbDC5k1DDy3YA
Yx4duFONmrw5yQMZaZqDnB4yytpDwW2s6FBMIZFjDPupL5l6r5kX/v0ETonD
vJ3bVObOFR8ksSJk5YqyTXnoASwg/TvKGdtUm+hPccedhVWkNPNV2W0Rg3sO
6ubTnz+J2KxYbsjEEYqpAWuaIz63yPEBjjO6V3im4fmu6ryRYSS3HSlgMRiU
iOdVF/nn1/5fr/q0uTU1EiYskr8VV2cEPtS9zMx0goXwViUntoUtQsjA4EZz
+y6i6/4Ym064szLMWaNht7psozUA3dbfFEwHgUAgn3MTPXCDkvc26N21KuA9
ytBF6FI/74OQEQjA1ROgXazmVFkRzLUqJD7flrycZbbLEXWEoHyThevjC1O1
J0ajkTHnNlTGEIdjr6cIgyMPoApJNgo+pKzj6cV/ErIXf1c0+Bo5R0grzKBf
TWa0l6sXlj7AeYscMMPT17L+oOJ0CmoeC0YocHO68duXrA4HjZfdpe1FrAM7
rR1m9HnqhV1G5dCDam6TZ34AR793KoFmdQjWU4PcbwCA/t3l5L17z9TZOLVA
nw8V7CBEEPY3voxLyKsfELtn6BS7A0sLimvODT321m97XEr2phgneA8f50ou
HO0fQMnzr3Ed24hM5/c/14u7Di+7vmIxS7kAfzdPcSFa++siNLKeCiO9W9Xm
4QLwRa3zQjK/1Cp1DYm8esUfMKioDowKkiGoWcXpgG1/1oV9jSVI8FPMrNyb
pMmne29to/BlZP18Z9enAWNYAc4XXilaVaKbnfCVLoFIkM70E173qAgQYTz3
2/ThLrQwJz/Ey+PQzRlv2LeIc80mWoeDoeiSaM81acIyxaDIRdmJj1ggHA8C
MMwkMdkTy6AKH5kf3yNIK7haHwEMTDQEA3JxPrV1OgbTVVif2pg6jYt8zQm7
icsVKaCpQzspOjTumfMY37MMzg4ROGWH9TKaasPCLxiqddrtbnkvTgOAMK6V
L6kRBnQ2Hdr0czq+JmBkDX5WOxgfvVW+//Jz71Qk4I5CmIyP5qpJ2Ps4HNdk
1OHegdtKn3h3dcedh9hIuqX/08gTQzj4jXGYg4LO7VMRusEM/C6WWhBRRmwY
4QaQAbtC8ruIHtESneJ/IY278SvpDYSy5Qk7SXdEaMP+barXJklBH9SHqGgd
IpSkXCr7drvTL387aLCo5Uk5uKVTuJ3OrnEbvEQKQ72r4RzmWPj8WSaw8TTP
Td6MqnqTMQq28TiX3GnrswK4K8wSY2v+QYT2yMT3vxwpHcnGVITnj/9zh8rs
VaxnQa5YGxqQ8J3XUwPgUPq7+2Hm8xc/oUSbT/xa3iH9fSM7crKPfV1TjpnY
nIPxskZAyM1zGcZ4sWhg1XPVQGJv3lChPc8MdJS5VhtoAgV2T7MysrvwmUYG
p9gAOTmqv2jf0WDxaTAqIqV+5WepTmgSEht6twrRZ+oPFsslMfj+/RRwSjLW
PVaad44U8hjZgduWt0YZxElWYLLxqF1dRsXEIWDX30rrqR90Aewm/kyUTBXZ
fvAGGMdZN/76DWIyKS+lErKAJTeqbYUnA9UAFGCTAG0SNh/YuPDyjLRjpVIJ
vbB+pCsfAGFZQt8yKznJvq/Jx2kHQpfW179evmmvKNl+isIZFeV5RKbTsAdU
y/wW3JqX8IyKfFw8cFgo6oCiVt1gsn7HWOZEVKMFEPjilzitNgdysTVDpdo+
FWdl69+zyTIPvPt3LTsPVOJJWj7j1+WjgfXf6//jpKZbe2VDBF/H8xcrO7PY
3vvkwcgh7FOkdDKH6HOPT0RNvGBgwRBy8CAZmC85/XwclUKjPXm3stwad+ey
Mss2jK6ZRMn+/DRlvA2ID80pcfUU5yiFJSIoga7yqOjtoaOTaTXAPgpFcYsD
g5daTOF1qIpHbcQJqyQXMFb0logaZuHEujdCHdSkwa9YrMQjaRmtcJecA8H5
cvVtnkei5gKfiXYMflQUjWyEkLSf2TIEO+oadTY8H8YHXY69I66S2o2P4Rmv
8FG1VeZujia6Nw10ixcSQwChx3GWuFNHI35fKfSVNfwxLvYW605Du0DaqclR
IaFHpRYXKa3zjNYVMMsztMY64XWjzKAbb34e/mPzdTF1HeYniZJouwtFa6OQ
Q2yy1851bBpTDwqsBz3xsjO9NyJU7RHKW3ugJXJd48Xf3pOruNzi4XOV5cb0
Sv4AzkASb/vzcNmr3bRNa2NArpNVo629i5tnUQPoxOVrp0pzgW48gEaLgY48
2cxTKSPlgcYFsg5udykqqTatAIbmu3pXeUPKE6vke2eB7KMuJnfXfCz28Xr2
JdDfvMZtO0Pzb2im+6NJhgXhxEaaKRDL7f5+TYYjsXnL/YA1reYlHvsdUEYJ
g0h4G8H0wJO0P7KyZNUA/nXFPs8xX4D1BtHr1tLc4r6SvbUSTEEPmbHNL/4n
p+RagZP5jgIiovXMyrhE86BK+wn6CZy2cUhkOAMEsMGXb87bho+NDGmU1UqO
y7eK75Pxgc/ShdA44L4f27gnam/vGhs01msMwAAvqgk8Ezk3EiTj/O9oc53I
bmZfLNAnd99GMpnD/ol+FpLSg2pr6xwJVDLbWwHuUnLoU7UUZxLSjwvloFOL
Oma1+z0nbivOxZMhNdr7V51zNNAyqwn0vLBaQ9knN+PuvQVHnVKtDNmfPB2n
kTk0GWA0HPRjceIT8JY3gmM1Z5MlUzJKegDhUo/F+MlPeGfwNLdmyfOXGfwJ
MLHblwRZ5lFOXNDMpD+aRGJbV15tH/H7xHkhc0mK9sCgZ1bX8dgUc9QG2tPj
kKCmys6gwfmOJCN4r+3PoU9680/5Sx6Wa8C7/2bVnt1IyQ9EUWux8UItS56u
pi1WsB2HVNzoLVmKhVIHxIbaQh3qy+5D4AN9/SkqvC9d5oekEOkYtPOZJwFn
7B+5ZcLpYKecmZTCWJt0DtJK+P2AB7jZ9uQJrHP9b79sFKZlJlc8MrK/cFGB
W8rJEJM8VdV5MY0vMPpwW/ow1n4ffuMFrEjp74ACWniReGugwSVcbGQTXpXB
VFno/F1/Z5NLgtZnpVshyeyUn+1JmxWtQEoalnNi1+hRGfa/VLhKBsBIkFh4
vG4BVCeYkpedhrk4uyaNSUY1upoMcgNp/JHtxNk5K88ejToJ0ahebXfSyNtn
1bZZH0Ih2qfdHTDR5v5gPAA5sn0OfVrkJI4UzHN68e6Ysx1ZR3w8JBAV+O0X
ydoqQcwvBTiOdf7WjJlzhXP4s+kMIHUJ676vZd7SxlW24/0LGOqmUTyoqSJj
y++p1BzYG5e1ww7vHW/6Hk1DhWCovoLFlEBcoDpDxT8mlc7QuDelp7n7TRHE
aI4B6BEZBnw329BXa7ibq06OsZQgbsTYqO4Xg/pfWharTj/E2P0RGvSiuOCR
eGNDvVItZ7czizgQOuLZq1T1r5QipIGUfqxki2pKjhJBnUOz9j2PZ6eCG+Tg
KA4m1sbpZKZwGvLumO/O6L03KOn/7VtgSseYt3q6Ok188LsMsiUtCfb2+HtZ
+wVIPGUdEB8T0ueXnO6GMwpAzozluZ+c2xOzh3PsFDuZzkaU2QLbl6ouzheK
tS/uFyqyZQrVi5fUjGLO7rj3l/ymANyeU+xOguJs2H6iWAxi/fXtl44jJKsm
eoS2m6e4M6U7aQrRxGBHZb4im1vKUKQCLqb/x2cgAPbLZSOwxlIzgw4rV7fH
+zDeF9kGWJWviRW0+l6F6ZinKu3x0i3airm1OzLejRYQr77uow36tQyY8rMP
Fr+iNi5CWMUcsSIqgSAewMGEIcpQPW83M/SPk7TmFM3+aKUq0sEGdqZ5mzyS
8NHO0uwlYzn/I1n0zzZe4qecpRO0RlyTvmmWgQmabJIYeLcndTuDw7zeA0Ol
oCgDHsPpBTBQzfIHXDTkTznIvY+/XKr9qIjLnix2goSUT+fI+XHMueTSeVMy
Vb1rWVzgVpW+ua6pilB1yrHt4s+lQgQEeYhGKhVm/P4BAoWv9xSq2dVIp2iS
L5Fvc273t0fymAbhaGSDFnxJGw6kC8ctKOO9FmsJGWIFa0yxtPTyklQg3q5X
mxiKFnEqWBzPjhw5dN6X/Hj6xCUc6KsfStdEDD7kOZ0EOwgmItpb5WGjNUbk
+lkzY4ErFRzTr6SyPhMa1BsidWwwcOPTVYyosq9+VBi62CJLvVuAf4YmzbVb
25Py8e4y+wSEaklnaux0awB4HGc4aQ2YlOj2rjMNaIpY6cmKB26qsde/b10G
oN2tWyS+2sntVJl1/GQ9SVYJdHkWhrTWzkVKEKvRA35Qi7nZ+ZRskoGrVKZV
O6Xmx0urE7ZJPTdmRsboMviItf9aGAWs3IYpB+X8ZSjQwQ960nZvc7o3h+Ub
p6AfBE2eDqUxf5TnwHIZSFw6R19UYfW3kLpJ8YyJrivNUKiwW5CDkvC3q1a3
IhiTQ8SiI0pnEFQiywXWxtLk8CO+C/79jriXP9QZKCNjGQayW6NwrzWv1Un1
cr20IFD2Cx1LyRFdtnjtmJZCADynI4145xE7W+R4/hBvYQ01EEyjpLiYUciM
bMEbGjX7gEVwsM0cqDsNv/oNydwpqoOrihL57pit/r9Lt7eZr0amMVxZSaaM
StBm5j4Fc3gQOFskdGkqSaVqBpIVCRmKn+XeLmXXcaC5QwLK38b1OJtkhQkn
6V8WhNJHdvIYTgY+sXlJjfY8BUG5bLOCkv5V0jt+g5QXFUnXUccWDYNLD04f
FbKZkEiqf/jqpJKghCmgz1oGQyo/1dK+9VqmiZZ615aoVFRyYbN74xH5sxC2
mXu76xB/B/lElElRDgVPaqtQkH7+MYsCddC3eOfkZdsSDFU6wikP58dNNEVf
M0RxDH7z2CnwdLSSOZIDh+k/kLeJQy3Dhkv9A6qVY6Hm+7abaqLtEMnmATcp
BokecyuIdGyeKWfQ8r6ZK2T15fkhaWT4VUAuysLd9AI39zfo/lyUskwPkhtx
oorHR3FexvIXri1GaFMKlBLb0m4E1CttG6cVo8qeQHnLDzYm3R030cZ0HRPb
X8BjgVo1jfguGrjjjsUMFNa1JucZKTOUeehAnyIUyq0n3FeQ4Pi9mE8Comgv
icu/NTCJxx6SFlCHFE/CR8TdnRtzIzAgTzTIPdC0djqtdzYKhDQLhsi2FOFu
rPwaLaoNxTGIKCB/974t4DMZbwQ09Ib/5oRfHmvH3P7VWzP5ZDSWSISqoafF
TH0wLDhtYxtZW0CeoSq6yzuVe22K2qZ0qRzQ3ZS6DMAvqcsqHb/UsZObMeuD
n3j1DFqPaOrjhHkbXUv9XIQu40yd2ByFd/AsmI87//4tahoNHIE8vadorAc5
4HiuReoKp0FpXXUnlEyFA8Cl80r7Xfkjd420E1g8JRDl5lQ3tP6gZH38NaoY
ehDXgEVCbgpnHs7vld0IJ3a0q1Y7uXMGF8wj8FpvQus9kJHvJkHlZ3mjBg2Q
bG7z0OmKUj0441huXUdNO88ifgwYueBtdZkxuNMchhLkTl9RUakebSZbwXZu
VZfD6jAga1rbJrXT1OWo28leKyThWXrHTMplTC74fGLFTg3Zxz/gKbwxKG0C
KDAuicvSUOmb5XecoGUZMcTAHvrRKn4SRwKc/VdhPTKRuzkXrpveUa3NQ1eS
NsF+e34d95hG+okiP+UncyTmiwVE2npVI6jl5pjRoHoH5We4bRvFJWjZDCUS
b/yuZLjvcuFC6N39CN42lsRnUDiZ1yoD8QOj5dGzaE+Cbdh5fXdbGYOEy4ZU
XzXfg/zAiYCC8YUm14WnqAOsRjKvQnNnFvK4bKcj8iLoJ2+7IVV3M1G4hZwL
rRn8SNs9RfJkkakAPbYrZQ7Ik3bnS/0MzFF7OVHSwUIz4wrFhAXf4HfiQFdz
e1qcehyGoe1cIGK3RE78eGmI0WO06s2Mi37K87J3UtrffqzCyZxjHLUQXd3c
oLrjH8aaRf9+7vuvvhMOsfvGX80ZZJhULtNGWnS3vbucJDJDlCdgqTYbX+K1
Kb4QtkoQ1bxseS08sWQRWi9DsTx87dcu33yqDfxyQ66j1pwcybARTULyjGHH
bIJZvFPPP2jhHL2o26fjRlc0H2OJT88QIA74qIEl1GGLVrLGaarUmVZoRnG4
vCuwgcES5+c5PXLPqcPFQwNcBB0z++8Lg4bNNX06/Z5G/MM9ei/GKQKiZhQp
sjZqrjwgR1SfuiERxfdtisRMmSALzsdaRJDkG4O/NwhrYl0twjFV/nZamo5c
lY9Jkhdej6nzDF8B0dZBSFHIW0k7ZMPeNUHKqULpcdZF4F2c1a64WsPVx5i+
5KBajNv2E1eTWepQHWPTH30BPg5R59Tbix/2j4Oh1FD1olCDmjWX/AUngfZQ
bfKPihoCNq8sXkVgChJ7hO7UuE7cXlKlpUjPOurZ9M/c7WfSOBpjuQtc74Kg
UW4FBMkbw0b2kodhL0HRNSqkJI1ivHCgjADX/Q+tSh4aLZiZNTykLhLlXIPw
rFX9EsJkyWFssMpuj1VBWJNmS1FTWNkvkKTyuhfzmyeJoU7lpXX92k2AOdda
nnHlvt6puOy92+j1urL5JR42oI1SclisWKbqrLFom6hHeBtEs+HOFCpBllja
J+C9W/y4ASgcH8sJAUWmYMbhN9PWRAQ4k5jd+pj9A+feY5T8uh3MsTjxt4KV
OcWg9zY8L5z+625QYpWnup5K2Bzjz8nBhtXRfOpbg4dwdWYMztdzE7vD3Q8s
M4+CL1lhDb+Q3OpMhRmqqe0PshYX3dIDNjwj6zvDYQdlk70ebBwi2Enj8kZd
OcmIvRyEAQHWnffRgC7DEDyv5h6CHwkNRn+rmM+Nt/RlX0wngZ4yfIy2BISV
FJv8kDDJ7LBvxirQtrvFKQcV5c6rCcrchQCIPqOom+fRCK61u0AJ+FNrQBke
F9ePeWLThF6YJjyQsKWhJRelEC5dWdy1YRMjwyjEsTuSb33Qjtl1os1y16UY
QWrgyzwJ5wFmlsHB2hTivCeAjCscTPZ2Rgxg/AedScyPteGSlyMAHJ48AKXH
/XDBBRgkVp29c2KTekCdZmegOWI2wD4j+1hXCfrDCE9tZ/UmEB3E//YC+ApC
lrGjQWk5K+hLfu1ANb7zMYeH+5dE8Tj5m8Bj/9I2Epy8HV6Xjh0vJXs+XOC+
DL0D/Ch1ae5axsFvcb6iJlplPWIygUvg47FuRxupljbF0to0tM7XcFEHqJfJ
Uuo7DjmhjZbAAp2qQNJ9AhGk5aGLvxLD3yinplz+A1gSWlq2rnqxkAGbYnwK
8Pi7T4wHTGjgF149XZdj5DohKVKgg+p2Q08gRktwC39698M/Z6bDx3SmCt+B
dTjybzjgUBBShFp7pFaVwJ3x6uUbUaDYyDNZdhvdppkK0ANAMNQRJl6Qttrd
4GedJLyp6mVchx6W3dpRhIHYt4fmYEjAR+XMDpnHdHzFvDQfjtmKCmPjNcXG
nQPYO5Cz/U6si/R8oeMS1rEMJUoYrRC69gZk12I57nISelzOUstPtSxnp3HW
09GgK31urvH2FlcWtmOr4z/EkU7+O8zcY/7+SfYTRUP0wWY6Vs51/oFIaUiG
r2Jrv1hYTWPm8tN/104ZdOCxGU9iPDpMyqf8uWXNw2hiHlhzEclDB0+MHP1Z
d6mld2dTjFWPMrhVIyU7mPUBaiyJ9sXDiswPlhXesPOZPfMyUADFb/B48aYp
F9inxuwbu/jGRXICfEpB7e4k0cq3B9fA+1ya1xem1Y+kDpSAq4DFv3hpr1u7
DRh6fTPXs0tDHoygC6OM35MZg5ehXm34UQmBQxhp6Q/W0PasNSKcy/FOf2rx
sAWkg3+q59XCGgps9V54mVS1q/UcMnbBo6lG8akx+Tn+i8XPVaNNe5kt9Y1R
Zqg53fb6Bk/9ScEgLX6C8e9gTDVV01+8rukmTQ8IIg5U1sii8Xozc5JIjJn5
ZApiCrKwP6MsN9GwH1Om7PMzVzfe6hwFEDFcs2ng15QKflgWnC+80KfMdf9U
ji4lK+SyGUqCJaFxvpYOxDkOpouIt1aFfM+4zN2OOD1I61tmOZmkoVP2p5Ot
qI70IzJYCDpjC/fd771HT0LPXe6uTJR0KgBk63+fhVpJ5TVR+oWkQWwCnaeB
Y5Vrz2H8k9bbJ9q+9+HNFk22+qLVgvgdXcZxGls1ybSjRPcGM8kJ1gCRBl0b
JGzMWsSalfv4/4W/+BwdLfGXVNdj58SVhBz4rJKc6pV8gdw6pb3iHQPhJLJS
/sFpCdcWLEsY7wyywFkMjD9wv5Cy9qVpQ+T3lztz1XMPoFxNwIZNvVbeE+IG
CI9a+wxY6+tkRpzpJ+nsHch9QsV8isByHYFvhoOHwlSTcd9O5e/b+tAJuReB
y0aIJ5oXI8hQkMMX/4XGC8GVHG5q/7ZPatxt5qmKAxUsbOeQ32sBoTx53Bqn
AR62H0C9OmatacqKQTlb63lJlWDTzfEGsD5MSLG4exHC+u33SbEhDnG3Q+Yx
9WJMtM9xBCI2+7DFCHftGGxhix15/YCLy04i5y11YBEJu/7ty5FoodBJRXYW
sKusZnJFeKVGPA4E3UvlIoM+seT0TWAZpmWI0gXi31Pn9qGKq4/3PqEyKUt2
YWL+tjziqnXd74liRe8yC98QTSYLAqZtyG6J5U6/Vc/QiPGnhV4524lCZTay
5JfUpBhDaiZJw7yrC5T7xuvizkrTxRxOtXiIKy4sV6AmDahzqzPWRosJwZYK
rKVZmUS6YkZFMDjE9cCXV4h/8UWff/UZVuuoyCg33QZGMh4K8kq91C1q0MXZ
JZ/zaTx/K5zHticFVm81xq3OowFsCdv8dewcEt7FhHFFHdFGF2dT6e/N8lpM
WhxUcaVQPdXrBb/rpRWjuUpmwFHnw09CNwxu/hqSV1dTsj8vZuRfd/jk/gqM
vT30O0r0Ic8xZV3Kla/KULZ5AlrVPqBQDUP2fNKcRklQXsfVi2vi/RoKndd4
TptVZL0Pc3uIjJlQlh7wpaiDFX52IMiwNfqDWID8jsRe4ZsHrSUwvxwn9eDD
+NTqIV1sDuJUewkhoYTeQL0hwXzFvKgWqdxwabN0pwrfYyk4DcmMvkBPJp18
SEzI8Kg2EOhNYZokE96lgi5yxH6Hk+1etvUgtPXW3AeQAVObDDat8khef9YN
j8f7/6MbohofYclbKyhzJqtE6D/GWYznET0inWBfie8/Ugw/DW/rPD8/f0nc
R77FLDtzLT5g7fFovNyF15XfMqC/RxAyTpldU4FsBglcflnE/MEud/ZkNT0R
uhsU17H9U2FvX0Wn424Ks/QC8pRXRUThue/NlHu5NS/FiA3UMR9E4WILMTtw
/2pzSE9IzUTmsEkgaIKEVStgaCrc/ZHZs0pG0jvZU6FA1XzR7EjgMG5lxxiY
cyj4csyQtX5sEqprGZizcR7PHDwqQvjs8wMBNxcx7v0nlDaMhHNgVQMV1+KS
uuDlq1bNJ6TU4Qyn2HJYDvaMBZwatRyNqx5fpzNxeBcgP3XJc0MufNPFLSJL
vAqGJllO3RjpFKeV+kUW18KELpsI2T7jnhK5/16eAlgOzKMvVURl26Q/wrmL
+gjzbNKiUBL3ltYu2HzvWdtAie24vF2tsAINrkV7k2v1VKit1nC3ZHMOttEL
aHNo+sixvZmpJohNZARuUMBp/0zWCjmZARk+lEs2gtw9yeNBEogHTMg4p3M0
FfBd4WD13+CAh/NXjYOQgCEkj86QwH8ceMI4eUCVJKAnUegu00kg7TePrT53
N1Y58ZTcviTe/1R4k28W2D0EH0Q0YXPwA3FjKhNC9+3AhcfqxPbODOvMKlQ/
TykAwHAgwzV0zSMTV85R3WPsmXMfeDUewT0wTAPY9MYhuZOvYb1SGnum1Pro
vNYlbu3yqNp6Uu+SG90OmfRSZrQL1R2Pz7lkvs7+PSahY+ZUWv9TvqmqFTEg
WBmBHkmjNaJOSqSlm6ICKBPS/lzfpiKUj3mleGG1EgzEp71uBEQUcw63NXJv
5fNzHDCIMvmwz/exObT66mdV6N6Fr7r25a95Exwz6WN2G5FZ/vv0OK8pF30z
oHdwvmLR5mQZKCdSVydpH7eazo4WxofJcex/DiiHkCKkNIN5lEjTghqM13TD
rgXo5WVLtVR77qmjsKXM/4Z/0ZpJR9fdR50fNEYZ1b6A9BW0+mpxJMLdHWT4
gJXAPGKNHYS4BeSBp/lehPRWZnIbegFHajuu38O5IFfZmZsrPKutI1l91ZP5
6YWCSvj48Th2PbUX+XEjS01Fy9x/q9RBQURWWtqc0RdUlvjjgO8OhmnJ0Gul
f9GXQw9eceZ0sJB+ZJWsKHnmyW0oGrlpmeZ9kmx7mV2CWgV0S9Eg5jTNTYD3
EGNNE+9IZKIN7QLKpBOQnXnkeZbzN5fbVRJfFpC0gbWU1Fd4FKum/PP3wInd
OqpfBZXsIZP2bTJPuQvaMTASlhA8Q+799DLtoN+MNq6yN7qn3XQsKryu4lSw
YXqcF0XGj0caF4wBDZ6gVHttSnUPjuXR1qFmgpRG9ii6MIgXOCQ6BzFtYewW
oBA8+IToDv9B1SuJr4Hwi1TTXwlPqJia0rt2AWYRZB+hURgp0smKxf0X7Rav
mg2eh+AXOU+7Tejcmj//mcPBIERxgzqixk12bjwvV+Sca2jhBXkdVFxHVU+F
OAaqHz3+TBitDIHxs9lZ1oXEux/5nJJpjh6aq+GvbALQxvC1/7FEwtzNSrFw
jkLOiM3HKhDRKRfr06YtKwCBgeLyPPraH/EzQ5ee5ul6ZnX6Fa5k4lfX0ImQ
2o8cEKIpOdo1Iqrg4QJZ5SJ2tTk6zWknMPRvl2AAbEgmqptrBS2dIn9LzktN
Pn0RoESUk4EwLfWB8OlSzP1tshQoUQlisBAfFGPo0oPytl8S5bhPIJG748b7
MVV7cZaeuSSL93SAbh46/tgGeZWxBh/riE570xv7XOMJQzc3MQwGoBjEk2N1
ynwgwCq6h9nUJhh6Vo2OONKI27IzZdhQAThvako+bBia0HZIS07JHuJsztwM
hlpg3Hx6hnuio7ylwFDp6QNd+aMr6DnPHdaNklQ25nUl/2VcOPJICsn6YhBm
UccTHAOfrYRCaK6FyEUy/s0eiNfDkbUFZz9HxDYzU/I6dqEIzVdj3RUHf/tw
FGFVvSmbB5JqmmT2n7rceqtH7PUEFiPEUK4QOYdq4DtmX6Wfx/Cbg1+tl4j1
DfYAHbZePZek6jvp2i1ZfVwgY+BrX9ZKXBoBcyimnV95VVur1L8M/vRvE32f
/0H5obn8001AFR+YZlUI/y8Rcu6YiicdTioS+VRSY6MpbKmqWPGvTkTBfUKm
6SoT1wXjhn6MdDW/TUTTTMRllMA5X54CLb+4YBSV4aeoQuNsJRgjbGKzhF36
2dYn1PmAYhV/5BTTIuM/JdLkBMo6pwbEwkKnT8+62bvTbyTafQap8BHrskCw
vkGNxLYCmpBaOtAiY1/LhUJP8O883w3OI9uTJap/h764lscFsnF+pjLYPgXK
pyv/ocYLTv96K0uuMLv0gPHrBjgahAHXd2wPnR9naJyaXnXkn+ta2PAOZs3R
WmGMLnNiUdcm7fUNywYCC5ZXNpx+iBo7kLT/a5loCO/dLx93VqCqpzPyxWz1
UDUH95KZUy3ImDEs6qhh79GtqfFARATNmsooZzmzuTqPIZwcxrMJoJCWg2Yh
JIx9lTQ89O2sLhUOQN8ry79b96A4QIzZ5Iq1K8fgf8urcNpIyAtbsNSyEDM2
VoDCE60/RFPJgt1isyuQchbWaBdRVG78KEWLWE7brhyQtFRmR0I3+vuUOBXn
IhHfiXR5usEXiqsCz1V6Ga/fndSj1U03LMxegYNUa+yCeLf0ux3ym3++CQAA
LnU5E94qPNom0p4b/MCsggx+Z2EgzWkK01xoCmDDQQPbo2W6wJf9CDafNi0s
IS6Qo8TWdQkguhcbaXUZ/IrBooMdvMqvnFSIUi6QOzZCxO7v2xmtWJKfn5WD
66q4LtaL3wWLc/9GOsIUtcnvwZtbRY8tVas4Q6Ad42S5yoXZ9G91XY/VK8yF
0H7dLnemWq0GjZGcBvy2AYYwtuDeB2tyhasdDb3za52yXQNFRJ0a75W6FWqW
4V5AfIKVRi2bYdvve17y+U6swMrpTPtCfgKIi6tfXd62tuet+fjYJPZoc2OM
i/n0Tif14hhRdpwrQt1rxl8tKmVLey5y7PDdib3XYKMnu9CLy39eKyuh1fuD
ddTqeYvgWyGw+pLiUx5AkjGWB1ifNAr8qIqWpMR8dd21b9EAxmkHEwNDkSRQ
mCyr+9XJiYcZ9sE3awRCfhniHWqHvfIW/WqzJwktTzS4LMz8BviKmsOQlWEJ
60lFxISXBfoJsHv/DhZbz8kun58Zr6uYHAVs/R1ornC4ffeqCRsL3FH8OITB
PKGQfFnKX4tKCIXUKxYgax1iqdSJqCdnsmyn7iB+zG1OeB6LZrOrDwtWJwYL
0pwZIscX9H0kGTDkl7E41+TiQ2AaVPqhyhSfXhU7cFmqqaeilHVaE30yA6Jl
+wR0bT+43SqMuL1MSf8fEf3fldC6K/yPQUdQ6Lsl0XouB1nfaOWuOtw4E05j
0sKddDKLJBqcEOdGkex2leM49Xz546gLSVz+GYFR0l3wfVGCAA9kDRsnb10s
qYK1wqeM+bbSlZLh96Zi2cn5gfwMPr5OO1Z4ZwoUDo7rIunf/F5sBm1G/i7q
GyIOpcX0V+vBOzCDSCXTA6B31Vhg6iyk2+nY6pyisJThGK7w0KP3/7STPNg7
LoO0zjb3EUDQA9cH0K0Dzb0ow0hMGOI/8mFAeIcKO2wJucrzKvHeLmSm/yA2
YAvsp42LuO0UWvFHixA3etbdDTX1zIrogc5KzHTfIXbunH0hzXxZ7tbXzNF8
gezsC9dMfS5g7vzvyPoZrtgBjKjESp4hORbgTWySuKPlZ9Nafwyp2yvOzqc8
exZfEmGfaH7NA6YP5g3qSLKsTCptU/x0DVYi+TeQKRJLAmTH3W3YGUhDUmO7
Gb7yoDafUveLxUolhguW1UjLVCehi+HXLS4tn2QgUpjyBDyCt5PeMA7t+szc
3qpTOAfihHW28umi+VCE8OTQ64tFYaXXlKtu6uDkb+iQk80MPEQgkjtO63t2
QU9CNWEHS0fgy6eMH7aLZlT4B08c/0JFWhCpcykv57HIbMrTGCiTRplCcUNW
6t/r02hvCO9+gvgNhK8AC3gdJ7Zvxjw7eiC5ZrlKZu+wHYtA1/vI9Amu61B7
oGI+VrZDLyISIRvj31zzuovN0vv4pymFIWQhwAmV7O8V2Idp2FpaBr7JMoK7
uuZbp+4E/UOkYDCnyKMXhInf+liadWcZIqjIX/w/wCfbBEpKWGX2eIKsD8mu
kgzp0pJ4VBSCWdnpg5ufVA1MqoZ/W7RejkIFN8C13cbnnyfvHzVUrHVoycz8
T5P2yMBLLADqjUIww2NXBOuzhkzpioedOg1XD6aybCCKd34fD5m/Zi3YSwSl
1nhcYJApPoEuKWivwKFQAhs/ahXyfQvywyJwPjlOYR2F0zAWd1lAROO2bKLL
KG/vTZf8XGsH2nJdc2BXrTfIqxM5hE0ZZguPHJSn4CBqEO5TFnx1oZOckW1S
W4Hdh5D6e+KmjF0kIZL/k4xLsl4NrAOC/kz1g1H7Y6v0Y9jIyL1ZqAF16kdR
Zqy1VPbBpRB8RMkSMPnfmqb8MNRhZFhBys2xs0enwLs/PFwLpCYZDDLpF9h4
5BMDAK5XBhSjemgWtxHF5uZBBdncEeiJb1seApZqbTv7HEhjO0vEwsyhGW1Z
05OlGWroYB7wjjCNJiyQg5iBtl08PVsU7J6Lz8nEDWM/rs1xMFUdLEk9f78Y
+G2ZoTQ4lBgA8Re2dRghe5DRiDsKFDd71IKn9m8Q04TjbzBvgfGTeHkkROKt
LqXi0ScJgXcrFIDQDylxjhJrq49U714ydc5S1VOcQAnHChcmCebwVHxdQVes
NhIcQ1eqHn1evgEiFhjFRee8UjhjU0r9hLJhBasighlJMEJhTlicUHu/YA01
ObEjm7WkiSkl2Fr06UpWY5F2vw4JQIznOx2hZYwIjGcc1iXIHTKqfJd9jxX4
Oi7e9WLJ/EJGq4ICxMqXgQYYeEop/KTtaJIdCGbZNJh+TljAPDWxtRnWcwbj
/ICk4vrAMZmWsoaAQ2bYwVMcjtud2SKNqK9w6GGsOaQr+DFWPh9XgQ128mvA
ayrpr2tOT/pQsGHECT8vDfzbEiebY9XhmE/QjpY+wS7OFtOdahInJeJgAYlL
hb4z3wODJLiRYjx48PX1DvhWSK2bOP4FIV/l5FiAnfT3zGhGuin0GiL+wsjb
7QHjk6fKRyyMAFWrI1dFG+2sWQbUpqAE/ZChiis1uflP+1fbcl0WJBzIoLOy
/pgJIibJ1PRE17323Z5IJJb3tAuyhCukJyqfu2hqIfGZbCLDlETsCN5xa1qT
O1m76noGe0y4zAGITBaXRjr2wwGQ/bxXXLDHVXBs4ONuajYnlJoKzgxVHbwL
rCPbqsm5gN5wj1FIOgYXJ0b6i2ptsEWNTbhpbMNtgieCu7DGBoVaSQNdjUmu
O4v0N649GfwDLdn8s9afN4g26G5pr4jKRnnlvJ6L+KCnzie9eZ141HY8t0vk
OD69PiJNlChdAL5Vv6UHOaofxoMlBegv36mHr5RB8ZcDfwBvOWAGG/jJaTBD
wCYeFRSfXRi+Z9do0tlF2IoXyaGMezaEGVC0u5diEQ/5wLVzwg6XahdAMwXr
lABFfCgV/uz43wRbx3DRaLW7e32Sf7hhp5pa0egpwQLSSLpLF1/J3fGpmy50
rASP7y3rHO5Jj+WtKbI2rkOpKW5Fjmig2W5aMwyIoRUy9AEOjkQy5lJqE2uc
LbB2g7iI4ag+DKu+I4ZuKevsLyAPx62ZMYs0PSwPTD+kBMwAqqpikI6QCPyX
/REJayE4UWdx8XiVCEqva492YCArMRpMIDcyFjMBzm/Z3S4XU0sDtx/ysHmY
zTIeRbLKh9U4AyYiwMuYrQ2HuUYM9dPq/OxVTKGkgaPo0IvP3KoU3FjbPTR1
iJyA27D2gIqfpcl3GcU4iuo2cMKjuRE6ir66IWFeZbX0O26pDPh9p+RB7eNY
wylU57068fE8eHv5McN45ngFwvac8Fb9SGuf7P0iIwrscTE0WT+R6h4JJrm+
rwJqjYicGt+4uXjzIdGX/z3SDoJmq2kTV/YvPqZGlYU+rwX5OdQx2Hqr94PW
VyIery8+tbBhR5MCJ+ESyH1MW6lKoZcBfIIavoXVUlntmfrey9CuYJnFy2xI
U7fdkwr7X/kTSWyaqQ87s/eoSzdwV2Si5wH+97+2LxR1entepFkq/eF1ch3r
g9R2IHnS9XGHDsZ6v1nk8c/Q25prfFXsQenGmyaAi025v+ESzEgoAM1ml8CA
K2ZbSUPrEJnNvWNpk1MRTT2Ac2YZZjMA6DWEgKRBN2bTvUiD78IB6V5liM7q
7Meaha0sJa+Se4NiI2QxNLqpu6lQOYF1JxknXdSaoXtL2aUKkj++EaEpQaev
MGx3JmrHf1WEJ1VC57v/RoYU2EyKdWRbc+HE003lMoe8xpYcuuRsMOSIAYhX
H5eFRATV4vHFEnbFABidImScRincdbFUFHxThn7M7L3yjdeDNnOWSZIsD9U2
lBsNB8dkOBRDX2lofdOM8cD/ptLKw924qOqUljagf6i1iANE2meyB38CNDtt
YIXnlwWm1eveA7PitAFRlug/HDH3lC0RmnECnUSuLYxSKVPt3TXsyQaEJtBb
r1K9g4HQqmj99uWpRrSlH685mPu4dEtWHGPWHLhAS6Kq1qeW/jrcCkmKKnPP
Z9yHd5MpsZNmplpkOOP8pPf5BGrWajmzI1rsr58c20ra5ooAt+dgXw7KuQdp
5Za7Mrq6QNdJR5/xxeBBsHktxI1i6WfBvo/+6hJd6LnFnmp1OhGg4TdyJb6x
l8/7iguLPoiql5VWziq1DS+5I0n1qxmLTCmn3fhTLKy7RDG9SQakNuhixRtm
ykm9ZpoC4J/+eitJFJ+TaVJrIqUFET7F4aLtznoalymlcY47TvjTXClv0A3y
HuBssgzrtQzv3oWKb4WXaVX9MQvzeRmH0tRyDlGJsL+8TV3nOBnNQrslJpat
z0tYx2wVU9/SyU61jDlRmx/zMhhE1xzSEcq3E/I6EN0Dk5JaIugR7WasamNT
zNcejSmqbB6sH1VTAEnW8gRNsxNjYPG09zAMmsOFVuro62kmoIh7QpXWKAmR
uC+PZCACiKWAgn8nHo6MXZz1JgofGu94MJRW35yFA7ESo50WhokrJf9e8F/h
bzeXetRlFv0+MsB84ecZ0J+BJIRDNTFNocVC0xepCfAL2W+AwZZmKrhcP30g
u3HFWYUARQndX3eK0NzOHPIzfjKouSQFK8iW1i9cjsNT6afU6I9UUq/Y2e8h
l+fcF9RZFnIUZhIwUGC6nWULh+1pJQszo3K0lxLx/sdSl82KtewUk/WfkDBo
GRGEK2Nts5JlQyYch2J0gO+kP13cwzMm5fjbZXs93g4oVNKFPrjWdlpL99ke
DjXZt/yoSzPS71JYfmkARJ82UxznU5ul+2Wh+tseXspOB5edlHLyWJLWKz/h
bM7BaLvfyn0tN7MfftZ7fm9cdM7GNtoUN/b1kb4xgV2Wnw4AKKw324bGTItH
ztF7QHhH3ycrFqyaZKC+voluu2gkRMWQTs1CYX7+4jmEuzUWRmehOxgqZOWe
Rgw7OjH9d+/+zuw2NwKJHj6Fd3mItcZaDeatb/090ygask8RNAH35C5gkvOk
YgdiUl8tcnXXQ4wsMIN/Q1faEuS5hQ+hZDnm0SHcvHgLPJJ7tf9UbfPyVqj6
witCrQyHSzaPwElBJ91/g6XTzupC0zzPHASvTFog92NDdY4h4xvs4NB0yWa0
r4BAIEUhxt+enyDmyyqDJ/lAUUkA4Uw3kVE+K5gSAcduVMRle8aaFzwKRyhv
s+wTgg36+EdfK5/nMXFbcRsFdLyFNti7Row969UbvQgKswBcHBDV96XatnIh
amzJ5QC2KeoPIcje8LvnpURSH8Ep8vPo4Qi5Mv7ws5l2qSCKRPhAa6QsgnV7
7bR/Vv+hMnYOBkCYJXJKyYwpoDXKPzygL9sMbvmiRf1sICcc9sAkiotRMkzL
5F0plXFabY4yakjfTeroMduwHFdSsp9ADoK0nH33tAg/VGYlWD94/12Oxkvw
rZzLfVLevU1UqBSo1Ka7z2rXkF//jNTWwiG+6jBctvnRu6AnSmvbZgZHFhY7
bGiCs3OmMR8SznSbBJjYJ/xZ9YLRtY6gEJCvIplI3+8kZCJ8I531N9s2Q+7R
XGX22uI9D+orjP0iGJpt2jutFDf90MCNG2uBzAePAcoWfmhQ96Ihud+PW7bW
IjYSBuCPD22Lmvimisc6UNRM5giLi9p6hD/92BYsGGCy47zUR+5UGl9hrTS8
3A/EdNpRUY2xuxGcqZLDIOBGf27BkKvWwyheoxr89VaWFCHkbcG93LFmxobA
2UW5nbAaiolDzislGZWPoi1WhjiAJhLS7pIMrl5GzJeUaUxHRDG0T4qU+ws+
ukW7sF3iMVX+8ci1zagxen3nPp1UTowJqmzmkUzgLnqhmTscbhZnu3HD5q8r
LtaXIOtrX+NKHhqi38sRxRUYahJfAlZwtcgPJ/PJXPtuEqOEk4f3RR4kBdmi
9QLJ39rrkjMYSBTgOZlxbgj3Suu1rv7GHVdHGo8r41MLCvQ2siqdeaz7LTnh
Sam6gj/dliKQQi0Y1AiPN1WRjdG9ffcbyUxCAr3MsUJGaSQ7Cc3bauOfEF6G
B9Pu/PHnOVtf2vyt2xIXE3AOmroHlwJqtJDg2yqR2hHVW03PR4xo/LspHt2x
VwERej6zdrOGECAM8quTv2DlxaOk9zqDZ4txddnbZRPEGNX4md7eKuT6lH2z
EwJhXQ2Mr0VoDBx7K9wy+pOIL0ktUTnsZoGCw5cXVCEsw/e3qAtIFNkmDi8Z
lkCzYLevMjgoqgLwFtPaGR83BJXYUFJx+MDx74safgpSzNaTKa54Dl+5RGse
ogyJYXmo7JS2Q08h7dRRknQbWD+xV6IUdRS/41/fMZ/lfnoCzVxv1knhFHHw
aH3id7C7+EqHpEl5L3/e5DyS2Ty4vSTXbesppXp7ozeDO0vjc4R0ZOxVcmXP
IJNunLvlUaMXkvI5GWBUz5HHudlkaXMNaF+C/TC1wZCzt3+IVfOJ1FPjZRxB
WeiYK9YxB4xHjSscjGU0S70Kn74bxWfEv2azYpF/IvwJBQII1x9MINGKsPrg
4es0YsdK3po03OadJXGF2+YXG7lx9aLRJ2WZ6AOqO0fky16YyjpGEthid1+/
OZiWX1PsY7lbihZICVQ+opKbD6e/U4WNFpDTs5O4LJ5fU0Bm5gEg8oCc5Z/v
C8pzYs9EBpMalvrEDtdAGrTKrfeUPy+e0Jqo4LvM9zVp1JXsbQE+GCiaHFQ0
vSHhWFb7ehBHyZ1Ew/jt+IvzYOefCVi8rkpH8zHwr2tiVT8y766vGb+xYatQ
he/7UH3HjJD60JDGqae8rwTZX1D+H6zcxz9Lt9NeI1kgL7ZF2JyZJHR9gC6k
+eOt/dYGhq7jW81/zrEAGS4Xr5/fp3eU8Mwv1XpIj7JoW17chfjywqQSfM1r
yE8lSfnSwCdPQnZj1i7N8RHugkUERFEdRaW5NXh8drX4GyE9rRC7sF5vY8DZ
VfRSd7b/Pwju4jrqZP29/h8G/p7gQd768pZ9NA+yw9Ve6mEy+BBIDKAlC+ze
kBx2M+cCR5Cm0f+gy5Jc74oYAhWLsZopBnko7kv1/p6rIDi3pCzJpdf7qbXX
9OwqJJjojAVCw2ISRs8R9yX6OhE5oTH/Fs8SjBYHiWzi35N1MIaCUWxY5yCU
yU//tW/370eByKrqYYrdBcMXeH5md0rSKjm9h3J1DsbFt9OVuXsRtFGWz2LY
R9C4OyapWT5T/AJ+9kAdxfimWlLh+cWosCqmFjKLteKuC/bcHowuhisybgaA
dbTyVa+62Qxj0nhqXUzepvlFZk1IVSOUKsehCb1yRwz9xAvmrSSWqE35nbcw
zk4+bFpuNOFGI1ktX4jN1wuA/+FnteiA/WWkKdpLOidXkt+nuPHcoaXykOVe
y6Ffhj5URqZBTr0e/TlP0IRxAdg392Qzt++5ps3ZvQV2pqlRATzCDhWw3DdI
bbNhrMLD/9eSopnUORl8KVicU0FK6D4DyKnIClModU86KQykTyUTC9pb85+j
CKr1xBwVBCteSVFtJjqmZ2xTrx7+7VyRxtWFI14ohCPykP+e5XmDaosEIKG7
dvIX9ph4Z0pulATb/Y9Oxz7oTGB00w7+Rd+sWR7zPO/wl/Tgl0jAu6b7T7I4
Ilq7CX7uGgE78CgvwzrPSSrq+3pxOQZc89e2ChT4TBel7r/+pcfvo7Ckm8Sw
LdFeFq39W+rS+QJAm+NTDXFKM+CzkOsRHVHamLq/zOv5gZ3V0CfHMG2m4R7A
1im91AeEPPYD+tFyA4ysXM/U2JUIWrYQfaLfvf6uJrKPOYwYkFUFwLw9i2BK
IVkDxfLCfleHXdcb78ynSOahK2aGBB7iC61SsU++jeWywyikqGWDHTcnqujh
oKcbVqT+eR6CxmiExhUe/Yp2PmhPs37KfQ2sko19BSsgz5V7pfiKHCpqmfOP
tNIvebsBqoKXy9HCJCywWEHAEH6O947+nFJsDAp6LWraGEVQ8f3W8pzf5G1x
XI8RL5Ov5Em0U/rLgtFmhGAJJsIyvDhjbyxsdEACC4fJ8VhpAvFUGp+Jz1BJ
rMeItykG3MdmzyHcNm3QkW5vj1h7thXcHyTKm/k00xdKfI65By/d7xbw2qI+
CXQNf8YEZLVaYVMwyQ4bhzVQBJe/kvCsa073GA6V2GxfJ093Tknt/Y5AQTCK
g55pDQRiKzMG+0GR/KdIA2Q7KtiGlv44KNxMvJKPDjG9XXNCk1mZq6AJgOT2
8toZ5gQU/LRLAw9BDeu3Y2UCKglyGFqiBVL887No0yFlavj0tPEZorXyQKVi
y8+m/QH67vtYNuU65EXDOiodKR1wwjstpFDkoN0FXg2cK4AU9YL21/Wqerk3
msLBeBWnq+K3/hbsyT/cu2fNZfUEOR73I54t7uNMzOVtRPb3avPJqrlgzFQx
dVLIEUHcfRXTrJoakMXAVfLTHC72BivRkDItj8vbPt48UXAGOANnHyrF8rDH
f5h7fdZnmoDkO1NkdKMykb3WEH84zbu3bU2Q1Q/F2nlwFfSC1mh0zAdGYIFr
X0WVyYQ7JsWs+x+/I7658zEYNd6l2XPYJSj88Sh/pgxXFPJrBpXmtg1ba05c
dpHnmBicTLTr+OWObVXwbJrd2si57C4T8qZE7+TEHpSAsCn6nngxca1/SVpS
5sWqakZnjTVE7Gb7lV6Ccp2/1kdJeVVYS9TowI0L/OeF3ySCdiGqvCj7YrXr
UksQIDO7WanU3Lhln4U1IhvlIb9rLoTJnNxP/Ktxa1CWRk855a1L/ZFT4+YN
1T6IAqbLSNm3afzpt3vyVp//WzSslP1fr1k9NIWu442B/XKDK+bVs4z96yxj
I/3r4ByvGAj3wu8RfJHyXdAApl6XcMl3G5t5Gll9bdmz06Oq47VmxxOXrK4L
IqPsmBIYVWW+oHcz7ToGDBOtZr52BPk8PhSY4FT3EXobl0RD3IjyTtMNLqlF
lAxumsKS/SHcbX7X1TzPvLryC1BCAnjRjExNSqphlmgdp18rK0qwuyUIkcda
8MzR0naYvkZ1vGGqzOl7gjw+IJFI8R6jfSJ+5frCt/ZlFOLK3z7hS/nP/rNw
0NffhiTLaqIFU9x7tj9ChXIiuJmsFLG+llQ9O8HHBalFyDVfachB+Jkz5FNo
3EXiqgsfJK9NL+WlupJGGRvhIpZ1ps6T1TEyFVY2EWmbIqrz4OvxE1M5hKq8
8wfVe3XnQKH+dX1qD438H/z3zWIyKPEP+ms6uUdBqo5fibmLy3e9mLU4uX7Z
MHjDFdC0HRWIBIyoTptALPIihvUKfcAvfutu/Aw6GlR1QPZJ6H68Jvo4zuUk
qrDhgV4cCqOfepY/nX7/GLXkQVEVM/rmL5mK60UKck7pYrpdReDDvfCaP74b
5ord3YDbN9LqoEDucwQKQK7NF5mSo42uyHzDnyUJRrxx2LRSb1KEkwGunrOc
GK4SQZwhdPi5C8LYUhXau+fsFuVGXzxnUl14HrbcNjm2M5stQkrJLtgWfZfk
bhRokXuPTowANgk4vDtZuMlBHVH7YFs3kjNIm4aW1QQVCviwt53zM0yJtLg5
VOeV9FMnBw6HskR6A6TdhDbMVuPNW404OZIwbB9/XGqj2GhebyBPgjJLnU06
YO3vEAhtxJEkm+Cgq/eU8j7GpiYcrZIxiT67yOcVGaknZ1Z+C8T6cUF8ws3b
yBZg4PAcAUlkNrBJ93LalbGK+DN6T5uvCPDNGR4i6zm82c5ofkIE3NV+Meqr
8BcbLmD2sZMH4bAkqB5tDG9+vHOmrLpIHVMiBC2uVUccuQUANDHYcBfVpOXh
u+IMA3OoNx5LYXBB96IZqT3TwwRombMaP5dWBsngeY2Fbx4wJSrLR5AzKQnL
rru6EjCLFlgrY9To1LfJyW/77sXzPo/jL07YG5OjaiGo9/O1oUPJ1yWwpQ7n
FZj0xFkwvN6yRoXbfmJwdiyN7vV4J78VWgdIMzQlfS92A5rAl+T0MTE5evnr
368hf9LsqzH2DtDSgRax9CXR2J1BaMhM4didoADPWHcF1hzoBn1fF0W01bRy
UFyVxknqfTUIGZc9rTCu92NGlgtkdGmzuvOSvzfm4MpubCp8rxvZ7Fhr7ooR
wsStsEgkZ4nC7QKnXFLfSsluaQ7dOQQTvvbJ4HnYpST3+5FhUpLVzpkIPG+4
XtDS3G5gLmtbozB/E9UNMNdU1qYQxDJTr9YntjPE2Zp9z7DAfwls2Bpikd8C
E/nw9aKPT9e2dV7ftLxY4f6DF9/AnupPXw3ix00KamUFpCsdWnZuQ3s5SoNG
fqUofXXeaRz3qBhTje3iRfCozBDSnPp+NgL+iTs8kG2HV+Iyolfzir9tzWdI
zZ4ZpgKRQVqbj42PfXPMZHoicbzdiywt8EhblFrLpJb7+ibrnnBAcfk+H0+Q
hMi4mRXIOUexedYSFmBT2B+lrjjQBOBDPJrll6Op5WD8u5SF1JLIQASgaQrh
UrcfnvPkZeBYajlUi3FrDGWHeDbgqmqk2Vjo+7O3Wrt46LH03XhM4b0W4giD
7epGSUvkWAfmr8t77ayn2hnOrUafpgKgCdTT4sIghSHBft8eU+R2fMoaeZZM
6KbaVe5/A7rqTDQ7LV2HaQCOEAyn5mIjQ1u8aTONiDNhH3LDi508NMIpGxJX
f2MLeACgP9kRy6ku5Bxh2YAciAIJ4A33I5OTfHBbKeeZD4MKb2hNk4Gds7MB
rSl1QlSUPZ1nsUDdrkdGgCYnDl5arAwCY2en0hpl/HI54/5ZaOaaRLtvhPqI
PJR9WbyViFUm+DD4CqPPEWn1hDKMMV512Ug/MoEZq6yLXHGqFbZNtLfQQxXx
7LDelu7kPRNRgIM6jeh7tVqy1S0UwkqYn6D46bTpQJ4Rrm30zIVZFCLouvWH
Km1eiDEUkbYzwnGIvM9knRowZDYuB1mAjxqKXTpktu0PeUI1N5NqUq9dwVkb
+DBvsoQLa4ulXBCdwwtycyeMsdTj53z3IjX/UweEbmi7czaBsz6y1LLecFe5
4SC0tYUtQAVPoc2SJxAXVKLZXIS0Wx+N8s9ieLYfvEj1kRi3A+nCeTImexy8
u/S5Liz3QevztKrgQbLmYtdFNdXBOgDXBvmBQBHP1/dj1xpA/Q2UtWebtc9U
4xZQgYV/7vv6xo8tQ0rXjr5DGVG0uuemMHdbKJi+AjZOQyqEUWaoZkbp50+5
8HRzMigKrWIrXwgqQuGsFF2muSlUKZOb8XBzo/yr3kNnZ2WSmaf+UJNW5wU8
Sfm4P68N2Qbxmv05RzrFU7wMlG9cdZVLZwTjQfFPGSMBrbpHtHxic/z/anBS
1z58wdbLoM8EO0j3WPz3msrwyByI8a43u4RVL2+1SoxDri+4XkpnuHoTC5dQ
ySgRsbpNIJa4o7WdGGQqYMsjDQHwgAyklWM1OhORYFF4kFjYlRSWz7SG5PIB
/N/lK1qDGxU2MCiPSEhoec4u09XskSa9gYq0ebX45NdhJ8BSsFB9l4tpfpWJ
jmrMBRw7m88u0v83RgBD+hjGvZqK3/QV+4qawTymT3605wTZEq3OC9SehGBS
KYyLSnobx0AybZmEjlJU/zLobEcrrhI69CMa6/v3aS//JjMiRMZyMPACt+jt
KuDj7WOLp/diJhkqbtzQVfVJnZYAJZsVe8IQxxCu1R3HUWOcMhUrPIyPHc+w
kdYCMslEfbFj9EbsrVp6flPQH8ozpj7x8XTqupj4DVYzuAHV8y3sILwlI6X0
4Aglrzv2/Nvk3Wqwg5lLRgua6udqer2ejPGAICXPvDKx2MAF4JY+WEDJoOb3
BuiHAQMGgLPDj3g6qbJE6QVH6OnCxRai37f59iWfeY5l75TjVkZVn0LgwWNf
rmF+p7pbQ2gkSSLZ1IxVx/n+xc7mNJtYnKjz5LRQKKFj4o/gqiqFg9xWmKsv
yyNN9uea/GsSlAP3/EV2uawFoedY8GWbGAvJPnzsvDiXWVbViKrY5k51THb0
+47uZegnogOWEOh6AzFOF2kaox6oFH9Y57vgE5HPn8XkS5GLno1RJrjmmG3R
6OVKOj7ZSTMyUnWW6xZlUKf2p+C329RDcGShZWH5N9Y9OHf7RfWnd1wz0vAB
MN/LHnnL7zzGuZwHxhLc7wgRejZhRKyV0YMp0xE73sFbh4HT+Zgnr4n5fyQP
OdGPG1XsG76gY/9ca/5eCXS1Ak/ASK4bt78MpZqGRpg/P3ci341+UEDaZWLz
09R497jeMxuHq2P+ybtTtNPdvXZWrUIhgEUURvk+KfukMhfKwPml2FCce+7/
V1nICRnow5QhK2fbYEHLRXV3HXhcY+3UsyPiVzXXALIwvX26A/yKzhV6uxPn
nbMdj4du5YWj7bjz8MPXktDF0Qqn6DQOYseh1D6/is2GdSsZRc30fCNV2ENS
34YO/iM0lj4x9LvVtC+8045snsAeJEcwnmlFbaQipLmNhsKgBwqx/LIy905T
Q+NHPkW01tJTJnpdMrCxvRjCHLwKYvBrH63sbmonr/n4RBf32+FJA3vnAUnt
LwrvLgy0ZoScZ3RZysG8p3qjI6NAY+ZhoeKXcoVXEuiwY5lsPY5IVafkmpju
OLCS1tePO32a3vsTiNOsQZDOsLLFvAPQFzR84CUqXGl79WEhOVun+r9xGhKl
ULg/WySNeOFD1uP9qEo7vAIR57d0/qnqtx3TfN5kqba7vL7ElqG0nBSHK7Yo
GNOd/djFcCfQss2j90GmJoEtJoNIMSUV3LWm/rj6Adla1ZNuC4M1KnrzIQKm
3GKxV3wvY8C974ZxafbCXHaBLtU9F6GW2MRX+PzrjxV7lAQ45uF4np6uhCAM
P+Cz8G/YQAvXpj5gwejINxTATDMUJCFlQxuhYNpljGI523Nsne9qBkhahGAX
RX5+bVNeA8WZX0eKqTK/ANagEf54uEfd/l13OqkRGLt/KiPh9NsLX9zwxzcw
Bf+1zLtswpOB42mOMbo/wrkZsLKf2lpTn5yJrST3hAC7YLbuEl4b/53aze8l
4Mt4scgxuZ0q/inkFM5RBvfbaa+3eDWxsEMk4gIU8aNogIM14wr2mlb7s8dd
NHTSLV/CXIhf/EV8SkFaZUzO5KC1hl5o6tOV+4ACTvzmyOKf6H3jzIg/q4gq
57Ghzk/fXTsnU47xfCIlFjjmg9HqzFtjV4+YO47Ke28RPBFyRrhuLxLO+U+g
kJJ4jv3xtubda9euW+4PZDpw+30zuCevkQ2zmDO1J7w98XrQwG2XSDkRU/gG
RIZvfjkz1CKeobcLg97+P3eJyJbCg/uS1lZ6noPMMsl8mr05GxESpwZ0wshJ
bWJzO3awGGXIp5seGTWLiTRM7+rHye6sfAD7OGqtkF6ZPtE+/VEa8kuYByNU
s+QPTt8/s2A7mSNl7ARa9A11M4L5ZBEsRaKkElRsslLPJVPHMiOlxFZHZtXO
yNsk63Pq84gIMcAAjTWauceYeuYYu742Kp5hLZhPczdhmrjKd9of6MqSnVm6
7MDi29UTayuJEhTD2+9KvhjtGnl9Yh55jMAzBuzFaSbTSeZb2DcTCV7IuKUW
sEsENG4NIHPSwYPeCKh7YFIOlG7MzA7/bgjNLO92y7afEwgFvZ2ki3UaSFxj
xZcGmfLVnOdIZ8Cagrkt5ftMqlJkYHhL7EmYLwP620UdYQcBzvrktl9WsaSr
XmQqB+FRfhYz/ZkZ9tqd0q9s+iUPLSlcpYyZfg4knw3fEiQ4qv9Mgl9otv0F
ZYJycLBDMnSD4dL8w25Kj5Gbok/3gK3AI/LeYMMUiji5FXIIEO2BlbhsTo6L
1c2klti5gGLYFNvxCSMl65GC1jC2hET52q3m6MimiWVtaV7JiKsh79uOYDPE
hTarJk6VrCD0u9EFKR5PibdYKbWw8TS7SsOoglAR1W5U8z7f7jEcmr/voIlN
YYccdraoHA/iME15ROTcmvz3/ZALMa8/jk2SmnC+vQ6I/LobeVdWonpuor1u
GO0+COEdrFxO8VlS7dPE8Ro7leowB1chBhySVuwt6LTmZWCUEl4IzG4aKHqz
yyMO5l15Q/nZC2EmRM2xCtoDHuxBVwvA1+p/SU2YWBp9fGwRwwwIDI+NhQPf
Q/zx5EZDYtRXmiXG2bc7o2g2c36MyOEAYzw7g2XF2DQqKyup6rvzsbSC42HB
m2p5d604Z4yJuooivRnfvOyD1A+3vxUUNeAEmxSq18RpOKifBegWB2krq1mj
QSl8/dSQd/36hyL2rxvferzZkmdu4fYdVDsm/RYsJIRzuATJiam5j5fn/0mx
U59OLJtu7Xk0ir9GDIZs5YFkJfPOW1A5Dqc0tgWaOCDkL7pG1t/bVPH2+VP/
REuxWlY0ajOc7zmpwhKySYjcx/MDD4vg7OdvVVNlZV8RKVQB0kEVpf3a4xH6
qEdtyLL1II8/1+OKmSVcRLoUW8fcwS+xGW1SVpxfeB0elvr0LCkKjVVa4q0Q
x1IV2HvtF5WQj8bxJ+BfKs+HeB0g/VQkwH6B1hWWRf08qrqg13TWB4CCjpt2
/7LmQKkev1ZjMKQmdeLbptv8ZrIeX71eF85NYeIvYV34WX6f4nsSMVrp2tRg
jENjvStWBF2uUfs57UYkoGbVxMCkTB/guVVXOTEZP2GcyZQgcGTByTYxueEO
Ebw5T+m5Wp+i2crBn7/cl/sXloW0HITz+Mziz9l0mq9QkFM34cOmYYnYc5yl
BROCsBK3sfV55yJ9b6/LyPdCHDVRelauM3I4gJ6IalIOOvPLJqoWcl/Bf/DC
/9n2IDntC/q4xiOJklRGvG+zHe0mbtLZNOdoTliKunpYM7w0FWmsAAz1S9L2
ggshoj9hWIcbuRpppXin3If2SSrOBpske8QkgKZRse4GH9WA563Q1j8gyQpm
39PdzFzkWpayYYjOzpTjZ9/yOWjm7JBLHvchWUyZR4npBmT7xjFzB/4HVobU
L0MywX4QlLre5IG687eQbvJjBP4jM8VV7EaRRUoGRa2yqd3voKYWD7QpzNEn
Kl6vyURt8DXXVxYcOOhMdENt/jrwP7C1dWAvIHxNih3fCySeOBVR+DDaPg07
EGsHZWmG2e9REhqY4OkZd13BXfhdQmaZwo+E2wouYuKLkZ50joWXRGorWq0G
yqBrkjfdI5+ISUybjFOg0O0i4wfGqokOTq3ZRGxYhsziSqLLwgjSILZ3QaBI
bXQIwKdFsusTdpUj5aVhKQYxH3KMzvdOw2SLlZztHXN7G691qrFaY7vlrDfT
qL4K7oiQFZyNnpb+a0KXDBG2wG8rdqnU4UxAcoBHRXkpptna/E+nxReOy50U
oJfDzreJ4UhGiNj6ZysxQaZspxH+VEnlwxvKSF0mzENQycVkwMaCLM2vqu0Z
Ez6pUp24JZUr7P7ROwVDA5czJVrbCvXCJTiTOS7ASXZycd0WhY9CumkD3mT/
xPpeFCEbGvCgA8OSLhrlVHKT7XBgFSF7GC4r6u21nlNj9pqFq75/+DL+59x0
LoK+EQyTPFE9kLSbAIAB6wfxtb+kcFna4jeW2T8EgmfOPqYBKeFE0tBS6R0I
GOGty+i99rRuyznsBPzwL/vYlZMVXMVoPWjNCaYnS6uLXCvb3uBcOzPyKitT
5jONxzqKDS1FTLrLYCugsCdzMMz9Ed+wyUdZG0HTtY2Z6GWnmhejYBnLmbXv
eE0ARJdWRkzEaadOYObAIJqceM72nOLNTp4dmoVVzg8z8t7bCA8s9r/b+ntb
Hsnuw3YxY6MTrEAIwQYmQEU1fiXde+L6rIK5qv1gJ0hxxMeoEHtw1mDcCZkL
lvTlFVgFlF79sB9tXaMkyiLkXAG/fJuCuETafuqrMD8Y8ezaVs/oxz67IMQ/
bzwm6S3VFn6yl0+TT5MrxbqWoV5iOo3pqQ8i37lKW2TCmyZdZN1eWAv4UJuX
bUBHSShuYxTWJJWx7plrBi9Q8xoAk6wD3n44yKJlqSgcVx7a4R4AijAWJ073
3bYuYUmZxkAN+DrVy0u3X/o9fiZ1ixsQjddCxxidXiUILzeuO4qw+U4JJKvC
cNo9Qufa94FAQV9Y4/PWUHYBwqkStzXBp6/sDkEh4c8gzZOajsR1jQz4ATsI
ld9GCuruFpfciGy77jgdkuLyeN2a5cU87m717/ZD/58FKbzwfiBrQ4B7w5JR
h/29rLVM9f7vjHq5CpXXJTQTtoN2AOKSLxYCuxSJk4fBDjtQXTSnrJmRJLX/
NwWzKSGPFbvSmTaMn84d5UnJt/fMMSGrgNQ6KgNbcNag25kzcx3Zdk1l/QtZ
AFIuC05UB66kdzAgaxdEZuA38wIv6hNTFN7mnkNYrhUBG6vXBiTMaMB+k+Hu
Gf6k1h/FXVeCp9RSOdZHbWgV6udAtKonWKznEYaJ6a+6DT22mFizgm9/bKY3
O5CUaTa7BQvUEeBLzeaoy+ai9aJM9kyNl5R4C15x5OM1yiOEPJM8yFg3HLf1
w2TxIlClsj+VVuKINIYLY24aWXcZjxldx5BT14wQsxihwlTUGxIz+xJtmDKr
wK4+w9CQRCVuel0OH+2DUpIkIZtJox9YHe7OF6Av1QHcuGMVKXMToerKuVR8
MSqY0wBiPa2vpQMvYL7mC0r74WysUeDJ7gt0h4gPTGBlym9nrVuhMT4LhOgv
eWnG0gaCZrqVnagQEE5RHs2NbTX3PYOWEGOX1ejgkMUl/a9dUyYQSAHUAJ2/
DmdjXIaTOUBz0YtBHe860K+qjriaIzHVeoqdLCaH5MCfEU7JZ46Zu7ZKdsTf
CwopZzGhuDl7SI+TaPct5Er0ZHjJ5HkWxB9gdqCkSCQ6kp4m9jvq3VKgRASM
L+Urky14bSct9VQEA7u4VSaryRGBGeZLZWRDBkLvdcXK+vvYbVcDK1ONzUvR
vPiDoJH2u8kIYD+XMAMaz3KPzqo4F3SV/P6ysnFesOd9PBtdyblj1LG9eds/
BlOUd6Qpb7m6XwSByein6l1mQT+ozPdTzjSt7blrTHD0JsrZJqm9pCCIdPIH
Sm8WEEfZcYP4qKNDKnRPW+p53DQ8lCTLRfd1wV5YP7puFfSXhYqIUosLaGNW
Xe8d4DIv3CxYRKgfffpNZL/Yoc8WOxv2QpRjzraIO29ryIEb0RzzxK06Apnw
WQ/fFGtWetoj53UGQJP5E462KGnFjrhzzF2mWctbAMdr/ATlp2u3BCc+8TFT
ubqoXl41P0Vzxggk5yuuVrtHPdCPVX354SpVRi63XYPGSpzPzz0UviMiNHv/
j02M3Mg16ahhTHgDeekz39LuJ8vSeJWdVE47LhRNaTt3OZDjT44+2FTICMdy
hbQU/XfdwhViWy/7MQPZJIWhC7FXhcDKm1psmWhULsjz6giAKZQNvmr5zEjf
lXeeBtx/6J3WI9yhzH2oLOPuQT1ifvHLAVooC0NFR0qhzYOMSqHQgdlBM3vA
PC78r9WydI53+b1vJ07vN/Fx2DGxZxjcWxcIAne/7IB50jjUnx3b29uZKwRD
m33qlwK2hOxCYxwPlPLTaCto94XsqOTYNcUh/m53bqSQ/uwdtfR+6r/iaWY8
84PuPiOurFl3MDa2QvujT9+dAJNtM+FMHjFzFSnRWK9F+MpgwUMzlq8BvuBk
m7rcfMWNJnfU0zAr8125xe9vBU00YDVzKI9XsnQv0I6rmS2gbSKQgUxds9vZ
P+hH/nYAJTAm4Ua7ades/KWHLEJh/Su5Pdv97yxxBu78U0G9qOO8ljDeFzJZ
pmHVm1avk2GKaodSwbd76/qeEC2J6i5qa6VSxwKykG4V/VQT1eMevfz3Fpv1
H8CgLadW5q90AgvO8MXb6mDIKhUuFZZlRG8ozdyDpY6Qe2gVeHb90J5cdey/
H2Li3vjMlv5e2TsD4LgSG1/JSn3wsfGKLeLrOVAIgu4BVPjclKt/DxBNapdy
louUTXYYbYnHZyKuvFCwiSLeUxZLjTqR6K+7QmSBGuW/BtSaR55yDit+jpby
093WCWYZ3MHHdjPgDmpj3fHVjnAJWq0BLlxSDQ71Du3HdrTOhjzXy54L/mum
ccyu0MMyfj9fY4ibLCW0YV5YAKgq0BaCBXWr/6tl/rtAEbTk83DLl5FIBbY2
6kJPWBGvWGOSPi9iHJh4crL2j+kGQVqudSxpyfx/OfIJvE0qgUhYpHRCJE8m
awLlSIMmEIBWym1bFYChWNAXgEnuW0UVJ4VYlTKkokADRzCuVUTQ2TGv84hA
yaqM9A8ZNmNQg0dmMw5LbaPaQct5WMo49yZjYHCdrJB7O851gs7NLYX9RW+a
WT6r5i9uVk8uOj4UoN+k1VMpOn74tSAZdQtEZpa1F7ZtOKDK0uPEh+lQ0YTN
mk00v2OiBmPjuuBmzqFhDcDx+4YsBbG/S8rPWRNfsUu2maygbIJOITSZC55V
x9v8bQsBfACVGlXVuJqkQ0dt1dDmSAX80ChSy9vD4h29l7MdshOq5luU86El
Mkl7S/TyxBz15KCB1csryejnC5/zOM5GEs86Sihb5sItp0i1hXrzfPlQy8sc
+FF0DspObtXjTOHY72M1oyD3W2MSsnfN97UOQAQ93YhEJ7sY55XhicIym8dW
HM25ZwBxPWay1hc6PTDG/BGzV6ymqEovp1+eFgB54zXGpkvoxn1tM146w/GN
QiyNW0BjryC7bB8h1suj98UyXkX2Bx9z9xYgP5OZz2SF6mlAy2lSl6AI9gak
0leaYp2rlm9MumDFsJtjQUP+3y7zHE6jPwvqI4vggQzU/vSbN8clKPDs2EMN
IKudN1MUPajojE4KmC1zYt2DNlbWsF4c8hKN38K1oAVuHYZ2KuuJ+8POzJmT
KsxLiEiR5ZF4VOhYEje1M73gGhPygoZGt8FFuQ7cvAZ7ps+IHot7gVgoTzXW
wf5XVspbA5xShqu5x62jCk5kF71j9XIh6AHq/NgrG3ioOCgz80wCGm4QgvcS
hlBPo64E6gHwGRpZEdHg4C+EV3cxo2omFvEwpWatsqP1xj960VXpZIgGDyiB
WmaqLDCEKOZYZxK7z2AYKURx7LgaLZ4XxlenJhoLZxaheM7zXsjs5cwj0q6C
2Q/hX7e5ICdk1MmmwdNvj/7lxkS9hRpgMk29z+xtfQL9+/m87hEw9vSRAqvq
vxJ59Tni+QKEOUsRo1GaEiqpnxUU1GfdgUJf5b1u95KgD0+G8DXG+Xz7JyqP
yXq88eAI6gQaNwFSRDqdfHTeWGLFeOwTFdJSzEQNi+Og5CSgiMga8DdEg5iG
gK9AREELrZWyMueT3aQlblD7isynoO3dSHGQsSDGIYe15CTIz8b6p5aQwP1H
XxYWX1utB2sXjNsW4ywSyHj65HltkLmYEZj0HumlThQTnNHZF4T5dBv2MgvM
kZj9ohtSepg9OUVeaymcXhqO34xtZvEx332APFrAcQcPSKLJfCljViRBrMt4
cX9TFl0HFzprlSauTjISvGSzxgh1CdhVFqiOuGYY08IykKZV1U24ALYBfXsl
FNpECOuiih8d04H737Q7awaFXgMyeX8z+vyYm1aLToFJpLeCSAUwkwmyZE+G
BbQAkIHSOJGN2FURLcXAJ7y23VGI1tvaLCnrqtxmAfjOrRn5YF/xTRUSVK6H
DEX5J5paSXMbKrcmwepsYKyzUeuXHVERb7gR+TpdktFaYm+1hrvjekli5B1a
fVv7FlpSjoTQ/1c0VZulYNFuAi+6AlU6KT6z6hlPsQlFzsAhkxm7/htgaMzF
LVUeQ5Zs90OR7eD/3kqIjb0C+YncWtobmIHf+VcrUHso9L3JAezP1kYYAsR/
CxSLK21bWdG1/kgetnvFc7pjG9/xEpRL5t0N3byK39tCki+Cqf4X7djO2Bvb
SryJtTKW+yGIEQMBReYxMaGdP5NiQYuZ6E40YyOfl6nZ+8gbPsJaadIO0tIK
FV5Ginlcp2lagWtk0DBgmJJ9auM2X47THS2o0q9/HeIgwkocTHzfmP2yVlQa
7ZfccojfsBzlUVhG20kccI6cmCq2ZuJr2CyHu/XK89Arc+TbUbfkM1zE+9I5
Axq29SasKB+xoiKMffIA0pw//SALK3i62GE0JRy1PLodD0ROWKe+zvpohthw
yQGZG9MCt+ptD0BStINS9+j0mwo8YZ5GNf1Z2vF4SQuouRvSxueogmT1HaxO
zatHOSLENOa2CNh0eDOEILF3NZV4LMRmE1OH1dLUuSeEwXWoZlf+6NC0dZdi
iB45dTSn7aCYeqzGnOqR/r7XgQ7+MblMDzqb4fyidBQBjocR+ky1FULFvRkG
0lAUi6bIwU9n5Z6EpijBaLQhc17O+EhJayJKcGKdyHoPFC9gFp/nbqyUe5+n
xZCEP0m/6bWGpUjMWmyxig0KMRIA+pxcBGArDbYFIOgAuT9fpdHcGZXz01IE
0vhxPoly/uL6NF7+HSQ5tGkt3zUMIKjyq83Xp5Hu/MwK/7mOBEww8EIB3RlA
0Mi92MhZjX6dIHLMV0V3NhJPmRBa3xVBcdqyb43FxlLd1h0GsWmsI1RjHEc5
I4RckpmweUofBMZVIPKoOgCejAf2nCJtR2Oi2q76BspFERvZ762bLhOwl9EZ
c1tb7i7QQfNaj+9aaBFni2roBc7cUCo7evMGjNU9KjViY4nyBQFK+BUSFwPe
ZqEOlO+prKcXCUzAUJFCMEYkIgpiEvaIkmhe03J5DuD0597I7nqVxs6LkR0w
jwMNH+zUwLyuXXIk3dQqV0aKIBepCiCYM2Cy9F82QaDhUg8CskwYn/C9FM8H
MsnkzrxCgWWkJordM2dZq6AKYFjoioLa1xXxhkbWdrKCIvUzLPvO7GXsdU75
Nsj2TPZifDUM7uvT0U1VJ5q2pHDBKBCyO2RHl9aR8RLoBMUANWAM0qXLuTdb
PYt5MYJzQkv3LltXPrKbApLKTvY8eS+xdyTPhay/x+mXcybpN71AfGKXAP9M
1ekDIQzSrK1l0cVvF/RYWAZJl5TINnt/FiOU0WDdsJkssn5Y1noLktsMdTuC
jQkYT+oiNUgI2jVYUPsWB0URTlEHrD8X48RSF9QwLezx838hjySJ85Gx0Z2t
zZ+HQCGKE7ciU2XRqq2LXYhUyQf2HEWmNtx732E1dBs3a/0WwGuFxNLy5F7Y
zVtV8sDVK/thAhhzIwUNwQPfiPA0iQ3X6WzuyIqwGt5XtaD/SmEOaHKZs8n7
KhntaM6+8Mi4zFTOHnReCDXKU6YH9eGItezYfGwenhUJGyRDudobd3Wyfkde
ix3qYvzE/qU4VHWCtsLaoPLwQLrhvU/0dmAuOmSpeZz5bjUIu1qv5TOdegAu
73SWMlrN189HD2FobaUywW6+BuxjpKoVx+YzKcEXpWk0+yjWsicqKjlB4STM
r5ZXYA29uqIiREgnBuTtSUpRpKy0feEvf8bR9+Cf3oFcNRF7rFIhqmYClKgt
59iB5uhRNJdWIO6Jo9Szrg+WR94L/t8U9RUdM6jBJHnMorrjQzs7M6KF4sef
u7IQA6BKIhoQtsfoj/KfLFjjxZebC4UcegV0rpXZ5zYu3Zx2tyuv80Z080LO
3K+h/rSyvHdN9k6ACj8/NL34fv5Da3JMcdrhD+g6tsGs9b34LByWFRYXL2fW
HVzCYMtfxBiN4T2nDFvM4Azs6YSl5VcpjP86UAzfMCYVo2cU4VtFobE9YZV9
z2FnBwLxn+4oVlbTLJ7lcMZCSWyzLq/meeAKqM27shs0b7ZnzYYqNDEqtFWK
YcH9XulDYxQZPfsADseRCiiAO7zUP5kqMeHQfp43KE4qqU3xuNHKqII7S7ce
BS+GCr/c/ewtKHU3i+go6gmGKTevaN0B4T1jon+vgrWxTubeEh3SymsU14Y8
zUzx3N3v2WBiYD3WLD2nolEo6B+p0TwMyLy/xm70zB1+p6fq5Uo94gPPUuQz
mBctz/cRcszUyCbLYyVEl9CFnLRTnvsTV7ZasedvA5Aop1CoyZA/KbRwV0VH
8d4UklS4p6xiTDBKZQhQYbKkqU5aXLfDYUVdH5NviYWjqJnEKoqcaWc5Rq1F
0krwHlYsvarGlmFLrvMOSD3ofU8AsJNs4JJ+UWlh4jSOZKgvYclFDmfY6vD0
xMXwGRFiy8Jszj9LwJ/Q2faytoLvu54pNaQ1k302YtGJRy0GxSZAQ0yAWrI8
MimBTOZRsbIBfhxdmVZWqMQbZa7sS0tfu/Wacvs81rcYKH/J5ve+jl7jR0QW
yAFg99Min1pof5GwtjMNRiWj91aMN5TsYq4UhdvCakeeIGsAQ6HB3n7xKD0Q
b7VYA5Hgqxzqx0ZJ3Nk6IqSDZB0NDDTZ1P2pGclqpyCN30HlyJYo9/W0CrA6
hSCBQSSsKD+sPwoj2NUSIcQKKLrvVkFb+BSBUMLBOcJLPmtqdKLJMs/C5CBc
mfsNFHcVDAJqJGRAwK+tr1OJiF7ipZuQggMweenPzPYRtkLMcOtKfNVvv8BL
S1y2Sq7yh8mqdZzwmj5GXYpGEOONTDt3sGTAh/cq4ppeRfhtAtfw7CQrx6J8
rAGm4x4D4g7GCW5wWIDih1OLJtr90YrFM5G2FlAtd6JlB4JXmOU91HE/L4pc
oQ+RXpri1fUIXVjdwf5A/PLwssZcBJOywC1R0fsI7GjjSCLv25a+6sHpnfhK
HJPCZ4KXQQCbdvMXB8uCr/EAR8ULRkyWq4QVKtwssxXCqIwFVm42qQOauNp3
arWXi26608FRdwhq68BOQhJpsIL2MqChnh2TDtGNxDzTjPV5VZxM1MOtl4MU
hsiu3ELIdILuoaBtcCQVElTj1rdWuV2sSRKg4IMXA+2t4Ui7/a6AoJZZWHx2
Jw8Oan5BmWqFrC7PqSmVs87KOyXxquCAKJ3OPnc8eYJZIgsbGdlY8RZT4EWw
D7eu+3VfxKrg9np4+eVmRLvx+YqdoRmvBh22MmsW0v3wSlKJvpXaDfxZOXsI
wxwQCzIXQ7NXnqK4kwwzSKEfcJfp4YbdawdGj3V1nDDpgnz5ZsFIhNgQM3qM
KryR8LuK9LRFE4orN7PnGA3Dzo/Bl64IGKlcJgATKeC3Eykis+gCN3tZWK1Y
cwWHuZuZiLYik2VT/X6ZFhJhFhE0o/hUYBEx6q2e9+Epi5I9eZwjM2Efk1Zc
aTQoHnmnAwsqC0a25yRnw7GGfUUsFVBFDVKPdWeQJL0SzFKLHwKQmWjGGoPZ
Dg1b0uVG6Yrd+AETYM2RuU6nJndWrAOZ5gZ03+Sgv5E8bTe+lAbJijSR9aEp
58VUA44O22IwXlaAPSsFvG6t9JKl/ULfoVz8384BskjtHk2ytxq8U816HIfs
tjtpioCg/axjtVbH0TzSNUxFKC2NsWIPWHz0vL1ktC45uNHjWnb9lmdRyg+v
DtLfYVs0LiiWwuAhM77lKtFTpZkCpKK1eciLqbiQ2hhFB7nHNAyQw/MiHRGn
Tt0PVQsPrpC70gjbx4zlt0i8RpWgem9X65TzHa3ftsS0LAetgXwwz5E3UL5+
jSDeUCBXvmyqLQrvd0W1tOqlPQizupuMmz6jdVFjIUFeANcW+xh9PCQ0Qgl7
pHblXRgZP5e/Eugbc4BefIQAokaAh4Y/lO984tGEolOqIYG1Ei8AsVbg23PD
GWtJ0kgj5YnfTzTkHyJG0L+VpE/2rMfj2hD7djlyeNUJFIr2axneZ5ZdijHB
qFfEg6wfoJRKovXdzx4xg5ed9PYieVZYy8WnHkWE143HdZnUeefONd/ewABm
3yc5kxFFEcFVkhQwsqsbHWvUZNlAoB9SPTt4NziDTVYZzbIA/huvAhTovAqX
Y/9Xpv07fizaBxFYx8qWeD2UQIVltJKxRSz650nKgAjdZ2wS5FUreHMJPKSf
rdRl3l//JmkomIYrs+3knP/IsSsD/swZvYFcIUEHSo9+IPiZTURmzHYkB9mU
u8B9NHHldAJVeerWuQNdCYSr/OsRYF9SGGlwPFFvKIXeMPGAKUjxxb+eSMAU
r41nzPX3FMXx+ILStb5pTKdJK4fdBifi007VYX/nuHj4KNJ+GwQ9y0L6VMR7
3iJB29WRk6cZSYyjY8BNb+979Id/pit5whb1Cj3iRXT0ri/K9TP/MEGFZWQL
zsWlCUvVXxu9I/DDucky0SoG/Of4PTXYFxT53ktF53ws+lT9BSgpyR62iRGO
aiDP/M0Xt+inzuVEg+1Ets7g4QPH7dRoKWziRQEWsjkzIG5RzzBrjyYKQx7h
lxgdO8aD3xMIUAioZ1FxPr/SuodvGspZBMj7US8kQ1e6zaIsSq2P4MRGc73A
0QEKHkK7SewTDTRFudsdNt4gIfbJ3weUchxF84IcJx9PT3f/isFdWNP66Kbj
GiEG3QCMYlR5sAuQiRI2NokHE4S2Tfu+L4XGLQzGzZYc5woYxB0oM5o6oLt/
tszdQA6JW4GDjYyj9DRYaN4WmVxCtPpUAb79U7UB2deUMBvZODWjD9+F0YNT
mU9AGkun7r9EzkJn5QpedxtHPEMTmU8M/5EbCptA6ix6fpZC7/kQXv4gqm0b
D0QYSq0r5/vuII25SjagvbPyHpw7S5dWcRQPQSGQ2jLjZZHu2TTmedjt63H7
Sd66AqzZyGAuLVPXAsH3G/x3+pRfe6r/WqaezCcjjv2HaE3Xi4hRaE74jDBd
XCoGnaUuYYcGHXjoo/sLSy/ig1AHjfqGfQmWeHWN7vXN7m8eC83KPuQtKBQm
qzVP0ZX5YXAg8VATCfzo72zDbiLA6R5RtHVim3jARUmNXgRM71Q/SBMyUxme
Q1lABP7oHehUhOrOJvZlfoOCPKgVBZMzlVUPHj0oKXbCVI6D+e0djyLTI2N7
KrBGpq8MX0ZlR8KKHS1NkqotCwC8moyRlIA/fF5s2Nrc1yPmPREqqVFkKHGW
J11geeR4aeemIQxs5GZSQUT+Fsb2aOxTzhdVVt8IgUOpanwlejWi0wWC1Eau
C8KQsflIQ/hRlCTo2bTXHEe7snx62LxP9WciyG27purD+CmQH5eSeDF+C3iD
FrmpvFOrwPvlixg/lhVGelozwsJlvUEQlL70h6vUjyCrEsp98IPj8sKp5dL/
VC/pJ3U9jksobkK1buNUW4y0efKby7LtNuFWefpNxyckoo8TA/bdSSVWpNxl
S3x74scOdd5bTwIrA+4NyhFrb6KiUGVDNwxFOAomaPY9Vfd2+/476LSHwgSA
3tUzqNO2edNJiVFRUCFBcoIXDpofWvUZy9VkTd/ZbK6Xyx65q1EdyVc3bSa7
2pDN5dMFeVc0Luwhzbh/xdKRC2G3qqS6TJh2TjLThSlccZAy0Ch7orPL+IwZ
z1NU5oCiR84lN4JBccE3AFsg+Bj7+FX2R5gFeQzpW9lYYiKJ9koYzbmLT+fe
8RpEsH2dp6pIYtBC/IJ2x53Oh8AuRQcln4+W1sFfX72PzcEThLRItZ+EBRyc
WKjbKHncNJ9NmSEA4om3br3ckicl03sqJvPjHDpSrBI8V6Z5hEJYZSfhytWa
bwHCWT9q2d+xjMV2friiSQiUWaz2BPiXR72uGlLc1aRWm88ci7KpvwqCsURU
4X5sZYL5sbFShlfBED1E4CdtOESqcCYaTDedBr4QhfrJfIcAoC6SyVwwUtrm
k2kPq7sUbHbps2u77sH0YRPoepkq5pm2qmTdFjFfpWycK+I12IwCDcz0fDmL
B7hcz+LgAohHGjsj1FkuaT1BrHtp8mzAOrPlFrz0uzCCclASp59U5H81gdwF
NCDlmtGn4AvqDKzf+LrQV4i0VRshbboq1Z4lwV1niRFk0oLqACW2KUFhMF0l
v0QK7zTBHCR2IwczLrYtxCI93ltAUtE2WpVeoJ3v8HcU5WY3lFb6krgZlKrj
Ne2aj+0C4NGyfZR+bmVKb5/UCQRojobVuLxtuDrJ6KI3tRU0R+EhQu7TusnU
d89NozMTX7X0CNqCtCjmHFyVTHmftNUgKeu9WULOxLjkDJKALZXFvB3E6fk7
LXg9fgurz+f/iuBZg337Ql+3Mdczovr17djx56eZIzCJO28afHa45Y337UQO
9T3HRUmI+SBAIx4MEQhmIgyqy+hqt31SsDHdmGa/aofdw66fGVBFcFr4dyzX
g80vqdI1fid6Gu9eeWOzBL0OBZ8p7kLACpU1qb7uWmOJZKiibGlPQTrpTt2p
E6PBvjB+HgYdOUyjjsQMvoY/gbW7gb3iBbYhl4dmlU3CIwH/AKoW5uxjX4r1
+GmSMDyf49PeHBZdAvRQ3MBgCvIW6pUn/+e0+v6ZsUSu8P2deiOxa2Vp/yPC
KjiMARRb0g3cM2KKhayjuQB8X8oe4W8oSvXokcyJ06tp53gQo+LZtZjugJ3l
HWVb4mXbGyLg8N+PZviMPrcTI9VZkjvm8y3RrFZL8/phopZ8j4VE3ZI3uDlh
J7GW6aHf7QeYddgtgIwi36JIxqn9tXDu532ccoOydkqMw2+31SdZgD/XkjxK
6b4R7d2IhFeM/Sl+zlPGGx8bWcxbx+qg36EDcwgxHqclZZmwkyClyBTxxDM9
OTME6UGPz7P9COEGHwl9/HI5kfZDqS+yhVI9CwywG6nOxDfZTyfPPcL+gyuX
KAA+rlps9X63b1mmx9iZi2aGssTbj5RMGlatXNc+D/Uk6TQCYuB7kM7G8o/f
IirU1yGLuWf/uV7Nzh1MCaNIOY7J2xYVe8Tc19mZH046QwpQPuPi8CBWUOwZ
g3uKn7gDiF7qvVJi/JzVn+4+Iie5+iWbVvFo/M72vj1qdvTqS+txREzhYYVk
vrsZXV0L1luqWkRL2ZrxxHZTqyW4fyLjRLCTquAkkUuOTo9hDaQ9ktX2mD8k
khEBhGezt9dHi5fvcZYeWRF7iDuqwv+Qr7lRgPaIAmVBJtC6oCunQLHrL4vE
ZeiKF0ZETciRPKW9dNLbb4c8P1wcpuOlpVe7FsQzZbyUN0USw9BSlsckowRk
JQzqHltxTjhRDAnolAwIAzy4GIPjcvIf36lCbU8F56RKzOdrh+m5lGgnHd6c
EXbWo4APPVrsbLw+J07pjxo0IqonHhpBabUa2JKvw5AJFdlFaClnaVuOhI62
va7w53hn7Gn5kSohy8Rz7LbfZXdUlnXK+rmDOwBqrEaS22+k6ZbasVbzk82d
OppN1Sf7G9TqZBkeByS1xulHlw1mF9A/asXyM8xze4rW2eFj9D2FedaCD46H
tvnBj8z9QerXeRQ7vFCRFUVKo/6XUGyK11a7eQnaDJocvaDCCt/4RphbMN9R
xHsBKt8hrgKmKRsH2uSsqCVJAnl+256ZTE6h0sKIPVNxshVPWG9RsD/wfXsr
Vn9USbvYKY3fhddFNU+brNUkIdh4W0MRbM0CLkFWJ2BDjQqpb72D23/5nm2f
TWmdcOacYyRnRJ7KNck74+M0Dz/ZreAuWNltYsDmU7Ox6nRF/BpC/MHMSl3F
E3ymgMIkpDpv0TqC4gcYzHIQYFBB93WEy5YrHsP6CClk1vqR8JL9aYNFkNnF
5EbTKjXS67qGOq/2EoArFcCwlpeEIFNbuA1Ol2zDHpsSs84jTGp+z1iFzM/b
UKo1NzQhunpynY+LzycspfQJNcBDn+pwFyTzmHcuB6qmHPfsQ0+33llBC5zF
btf51ogjZz1ycPcqaY4AJkuTcT1gJRPFqDD3zIxE5TIkuaBU239/DwDe4IeH
NQwgrrqLts4+m1FpUXS1YE5Im5ldst3PBHm09Y0LN0XyxX8mVDiLHxUINLtP
TEgA1UqO+cqqDV4Lo/PMKHwA9du+5ppB/Wp9W7qjNkEaQ/FBldGgWj+eHf+9
qugeKQIy+ecFtYUnl8JeopF5HCfV0FZ7djQHHtZkT53uYfLO0fTHYG1R61g2
zkIysQbRViv4u98Baq+JZq38u+fjngsAnhxkxPmCWvEu9K0M6ulXEh1AnAdK
5FFKY7NXBHigGX6Mt+Rj8/9Glsgq9pfqZYEA5y2pSpaI7lGIXy+E5IkGN9fR
mPjwo/2vfICVjll1V15eVjaTzpoRb909nabTwXibE2OY1vzQH610dC00L9oO
FAx1sT1CYMuwbM02fZl69oMl4W8yHYDAiyw7U5MWRT8cAq0YvT9zloj8ArXa
9uN4I/Z3jIjFi+2960E+Cen36M8NWmkybZ/cx6894+yNz/a2u7pGDMvQ6sDE
Kto2QwgnlkUC8a5/vp95FjMS7CFW2tyrRaC9IMB7NmxqgRPw7GkPz2ER5ITF
J2XndONeKKlYCmUhVzHPpQDGlNj4eni4t9qF58QwCWX9brFvhZlvBsUCjUSC
ds+8lADc49XkZVC9hlawFx1F6QkQIJByfuGc7HULS3ZBxm4GqO3wckz7I5EM
Bkn3eWkHe8LcXCQR1XNfY5xdyQWo1+R6pAcD/LdvFhKXmO1lcmEhFOTXgeoM
oHrx3zxFgtNwsEfIe8+lMqnAvrtexQZJCdiAR31Yr8BQSqxqrWwiVGrFhO72
w0P2qfKCHTR4hUHwqYlgl3nJdqzifG4WS5napQLY0ijvku+qcFTtdHJ0ojRH
YqOTBQ2h3PB1Sjl1T6tgNTfP8rHts+ntfDsFlN0PeGTwKDoky75QcARbBULt
9JrPzCgXvIaMpFGc3+QhhR5vXsFFe3BCaWHIgOvvAjJx9kRWOJkTvMOrMGTJ
PgLZOoFV50mOrP8Er2SSSLHUklcEh5EQCKev8rBzUSDQhaJpPq1Yf4Y+ywOB
roOU9OI3cxpnfxnTkSiMvlLH3BUyTX/pLHj1FwLfIakUgv3aBAIerc4wAOJC
YxE81rWOfyHyxPW7OoW82kZGG65thEPqByHI2EJxnR0AMyp5HDroxeKyl8my
Asn/85sull7hFjiSCZu6lJopvQhIQ9+Pq7YKuKjT33JqK6BgaQf02cSBf+Ao
V3dw35bXWX4uSJ4RYtJ0lyWFbzb5ZBSpNee70n7e7EDvIcyCsO7gUD4HuzUu
EYj2JaHmy3kapEYOV5jx6rTj9QSMZym0RjjzmKUZop3CaQS8tW8c3DD/CDqV
QaYoHt9scbWN4bTZPnfIg6MdyfdHyjgzSDN+844U+UbCUhe7SnpY20skzXdx
mnsLVNMoyeP6v/IdHYbwzilHlpqOLkYWmIk0NDrN4hapXQs8ToNfJ0EjXDkL
RhDAlqAsd7lzOH7ZbFTs3zFmJqrL5iZeK9tvt5O8rfjFAJtwsfJrF8gZgqTJ
aPjZYnhcu3Vl6TI3O+UvwjtJnoFW1AgmIZAAlxIOIEtXhTuBxHQ5y4uhZ1qg
W5LP5WcUogpo06Yf+sIBWGnMBPknzV5vkD/xyt08xAuQ0Pptyi+pPN5CG//k
gJmEewCTN7lOYTHPTqFXp02x03zA2uMkgKZmiBSPzUc/n//MeVBmSnJJ9HZA
unVzXaV9GRwERSwhlPihCp5vaBbFi1hl/xxttnCH9hrXqvmiLeBYW1L997vG
eAOxB7QK439phO/JVdLQkRz7vrPuDmWut69VqKL7S9WWNBIud9sYum9P38Gc
kPW2soJfASl7IwPz2VSR7bZb4Sssj7kBlAbl+GeMX/ySZumpNqCMYHeDtwg2
iPuCDmqZ9at/S8rR83EI/+bMoYD7RrQO9I1qakkoxfCXBv6wcOGA80yrgYnZ
yUIMtRzohh5NfqaLxlJMXix7yTu055jDLM2Dx8i5H3xX6IT/DWqQ4pJ51ALF
XLWtswxQydQpzm3qdvrDPI+s/u8ykaxAOdoqyy29lU5vIS5JjuXKa8iBt6RT
5Ms4oxsMlsJ28dj05M7EcO737jgxHFyvx5LgX6Ot91O8hQmIPNadxoTt16Bf
2ODDyjDQOU6GRDLxVwKB+ihMNkxQD833QRZ8jrR2I8ua96qJ2fiJXj0E4qHr
EnRW7X9j7iyelbGF1x7o9XuK6BdMGN6VnhV83LhlZxGksR8/At7mclfMAeHl
EkHsmxarKOz1EfPATXjdYHLFh4ePpSORPil9k98wn9+tZhpWVOj1VJUSnDfK
t/TgZ+0fWbFThUBWht9UUT1ng5zyKtmjh1ndwNqnN3h4JmfZU2bLORR65s7R
R//ow4Y3MyiMCL2AY4uOKq2bjFJKQv3V0uIbN+Cnyg64k4osZyEYPbn0xXai
8hiJgfo+aYNA4r7Mm+iCWsOBbrxDjf0++t5RZbjRaFh95zx/pAPUyGDef11J
thT7f7sw7lzOmhfIXtZusMBCvC8fcQpsstEamW3SJ+tYOm/3HldseXAMmFn1
a/BAJNd9TrDhVFDmyVq/+PbZmK18Y2m4v0L6FE18fnVxcshGZ+vH1PYNkCiy
IoCgufcstyUoXn61QnKI4HR+1rUvd9e/cd3DnWNRkGelHquI2yNn1afixo8x
EPygleGfMK2dPKzfLV7aYAqrYkjrKG3eSPOCxteiKVKvP/wQvAC/tQDGl92w
oxB+p2IMpHSmOehevPBI5r6KLnfMgJVxTwm2bSMUqQv6nOAovrTT/RLxF15G
oQnYkOjvgYPF2BAvlrrzypoFlrjG7jZcXwJLWqe3KTrCVxbV95c15SwVD4Kx
994jSPYe0SixaeyszuThd9AutyUl/ytnWeW1t+rb9N9/bP4E17b9cSGbx1ai
Oo1mMfT8Bg5XrPPfT0u4vvWK5JjTihjztbdt4gf8+R/vm+zJ142+h+dh8h6Y
s+7uVDs5/3bQNdFBs/I7QVEn4zEoxHy4MetzGzQkSZtFuuI+c4frJ8yK20Xk
Lk7xgHCK7iVC/UwjTwfgkOO/QTrE+z/Ye6Emnfcw/LaMiY68FC5/esNQXkss
ipds+BnoJ1mAsMXYOBKKDhInmW0DWwiu2WBgbAGxUGsFdGfQhlJpUCqgeXB7
KFiESK0sBLk0RCzFuxIu4ZVWri4opdICktiyUaFD6rUJQrL0Ab4eO40Rqnrh
Wo64hR6E8aqpQQFpmG0u1T7jH7FuUIY/yarv17mf3gFi1hZFXKBvpcQtrRfv
Fd4IbfkFKIepy1/7Us/JWHXa7oBJS1lm+83nwMR5iYS8e/z3aIIryTvtvR1d
jCJ9K+9t3mAe/ociUE//O/3bWnXX9c3ecxZkBCL/em8lSaKHr6Q4uX65Qvor
LHnzDDl5DJEVO9VY/4vTFlP4Py1LRPsdozfGe6CEjvjToQ4bwXiB947hgPC8
kWMFaKM/dAmOTttq29NfeHyn/yEze4ush9h1WFW9+g8ePEQbNOoTtOgboLcj
GD/ssQcq6n+fBFhvp7PjzIPv9PxuUYKtQB7dskhXxe7mLLV0f0/xP1SBAoJr
4OgCrKV62Jcvm5bkGsOODjsPLnRaHWh/zsROrnZpYvn58S4+5cJJPTok/T5V
yaQivn8gfCjxEEn7j/+5Px3CVZCpO7/ctS1dT+lIO3O3s7ab88rGEOVucah1
jwGkI+frwMOUwdOWPBbMEA8p1Aun04+c1WocrLXNp3jReUMZnBH8MrOTiKMT
C73sIoW8AQ53A2wJWDBE7IeDfLzjkoIGkxCSIfcJ9NFvxE9clFYaoj2915aY
b/JbnwSQv9Jfcz3uf5w4TlRhPZmcHakmEkw+WGNI/x92rDsfsWZB/pSt1Awi
e+YRswdqI2mVv/tvuo8K+vU0ye0WyB5/DEtkH8SiX647k1n0Y9+4fbYRnURP
vdWtO0y/G+meWXHcF5VEyEG4Qg4qU5nay+TJzzskTIiMDLbJvCZgNHzE0KIb
HKCQglEqzuJh88fMQ2NrEyX3TdsCDbOr+D1MiuGPggdoUf5jII+cLy/MpEFy
PPD+/kQN52+DfPWjHNm3XC2JCFSo5FvOh5IGo/KrQy5ZBoYWf9lyiUeCMbO0
S4dSZDnAY8JqXimHbYlK5Ug4Clhwa61YxMY5dGKjA06Q5SEQs8laasjeVeYV
OX8lT120oUAqD+EeSmL5O0UjQzhEKdGP1FBmFCK9LdAGo+m5xzFPMHvmcyo7
z1GcEO6EGUsGow1+zyZPkDplhAA1PNhIZSnHZb69yYm6brFBPNwgoQkwQPkX
+01IhrTRtTPRWzjaWsPmOg42bOzSx6sVigsSnKSvwDr71lRl7cLq7IqeyCu8
SNYkm1KeP8kpmwhMY0/K8yt+cV4JMqtCW7vmV/8KkPjArJhHz1XDU7eC4Ayt
QLvEfZ9KHVwsITiOMn/uhrhFjIfw0s2qktee7zUmCpW0BT71SD0F5Hn5dp9/
KgCF/VyT9X+Zmfx9cULLScdmx4FwOK85FMCoDTQSPQ70vvMlJcawWpmbX2HA
FJqJO39Q8aL6PoCGMhLkfhVK7yN7ZHHE3bCZbvTuQpC8svgXud5NhTDJX3wH
4i3cigzSfXgfdBWjanYH2Yzict3K6tbvtmL/xaXCiZc2hAFc9CmxHaF6eJaR
vg+D8YpKirzKj2GP26K/TDCR+D2zJyP0gIn0eehKHnvsh/dl43iD61o0kVfM
/BvaTrGAibDC2M25J7Zjxrer3D/MFDXP0CRNFuK6cqxEQdKuVAas5c3ZjCK0
AWmEEb1g+1MhrUEC9rbTW+chgsjLdfg/XRx6GPa9Y36h0a7BRcnswGfcSXqb
2K4UwPTUqRqPjxleH+v+WxfbN7KiK8/ydzfQMXRxv9Nie6Tb6SR5sOTRSnvn
XqmeuyOjdkIHlPJ/3qPlwWbj9FLFTE0O/uRWBsRe6v9T8S+Nr6zw1oGBWqBo
GQBoW5ekMEU0bvTu2oN1nqzG5+KMvvRxplU6TFPKI4ZiSfsZXIHOq42J5005
/D6992Z9V7fHDB5icJw59rEA/dSbKWubWpDt0IEKpxSNUjvNz3DTs5ZgGyHR
wKgRpkZHkoZle0UoyFASVFLR4dBw/F6JGs9szed5DTuEMXDh/vrJErhmb6KB
8+LTlSiBwV/eycQWxQPj1GqvNhm2VrnU6ESUguCbe1i2K+OsJQwOoU/ID0W2
6+AYdHUyI70E6HcPddBScru4PBKSjNsZ55H3hkJjpWH2XzEPsiavXHiTxxae
0AZqELtfEMlw+un1RPbs0KMMDA8z90VGynZ6WfAPBNWkeRb+IhtKJuMF+G1+
vUWd7FgJuM9i/Mc7nmGV0ehke+ef/0ZWAWU3SWUKnSB5/ZOgLPdrq7oUzOND
FnnoCV1F1TlfS45N556klx3RuH1O4Th0xQEEmKJkBfX71SobUiFxDOzwalSn
lXD6vPgwSlXp1jz4g7ypxM+6DiSeFYNDqCoDjahzRUBUKb6jTPMYzkW+8hkO
6Hff8eYkKvDsvp8p+ergWQV4EU/I22XqSujhNns7EitoZU8J6DA9s6fF1Rdw
LaFLa3QvtdQ/M5FkyeuvyCXu+BsKburmGxkoKgqBwfHUG8JeR6m64Oi1cI6W
5wcac8h6LPK1l4IRhX9hePXlnRBOb9UFwCCn4yGHsdJwkAdeHOZl+cDgnOE5
+yBoB8vcYaCIweLyEpm3JZskjrFQm7iPWAYiHuGyCB2KrNdu8xVS1xYC+1xr
sCoPl62h9WsXrCxsomtUTR0pykS1HiB3MTe43da6QckEHqi2bYHovK852RaW
zs3tdIF8QNKqu9+H18FO/e1/Hg8Y5/ajJdygVBLtEg41B1hDufFbxlsQp5EX
HTYCTYP8t77gKqfOBmTNmlXyLJdi/Z+mrTsRnHmpJio+sjqctYygxwlOkxr4
rVlcO/nll5dMMxudWoonxV0i42+0GDGAqcpvDt+KcdVwRF9wj2UkRDsQAG2I
5d5hrJduiHa2X39MspEiwUcTTqm3MgB10I/BY4qBQxp4e9NLK2g9oAa4HXkb
kRp6qVyl/qayFiJTGctopDVcc/wvkWY06JComomDlqMSYCePc5rr4gS3UcTi
icz1RF1zMVoS06AdpAMWVXYV0T5lBdYIBU/XVVdX8TjDMOgf2DAXiMuw37tT
Ws3cOA4SJiDjVwslquZ4DYUwQo5yQsTBNE4xQEV1YSDCcVYCZ9/ByNG/8bwr
ffasMVFdiZgGLPC0ah5lYKDNvTEuW74dV09ulbMYm16CCSgit3xOqpm5MJ9F
y3sHUImuL0Abwav0VQf19fohCdcEV86joIkCYT97w6z3gZVHxI5oUm09N8LD
LGw3j1eb3/Yu5Djyd53aIt+OgZ0FuefLqovauCrF0iC22DzJ+G66Ahc0mkYU
YBAQGhQx9bSQBDnzsDupYfCbh+7jf8DijZafbgc1I9dM9bExV83NnfMSsTJd
VIvOoQhTfXD9DwYUT9FSp6hEfxQnwfkRPwuGUwr79uxGMyc0zd9sZmWwp2kD
QaO4G3z5p8qMhqVo0WCiOAAZa5dralzDgeSKmwdyR7t/PbBpgHVoKvUD9UDl
A2ZKKhTD5I4O6mGBsuv7K0AGstJ3ltgO97nQc0n6pnZEH8MTBXhwdatJrS0O
iC1Eih3l+cGjERSnLeJn+ciYehCyQMzj4tld8YPer9h4nSQjQdUxrEwupsRR
/DZ12h5dWo6kldDP4VeyjAkk6iB7BSvVw3NW2oczj5TYakwE6jsprDbvAyuO
sseL1kTMsIf/6djSF3OERZdc4kX/GcCmTB5a/iKWSUy1pzPPCSQv+f943g3A
qMEy2BUiXAGLBLl7dvRetc3hISzk3FqD6U4qsftlEUekzprpuuHh+wIgCnJY
ybAWYrpJwfZYrPBiuKCFEGI32688aN+JHcNdOXWIpvYfEuU33HTgSYiAPLIH
SiVHJyj2JGpni24NkjLGiR4sgZauRlYQDY8BUztnOaJMPOn/MWQcnewBBAQc
W+a9PixUrcYuWLNc7C4NCenVZFBovuiber+HU5FvxWU1Ujhzwd9a39pA7xM8
rWvwf3t4Ng63g390OQoL5Pl66GCJzcsLgVGXkasuhMw2FnaU0p7Nnbtk4pZ6
8O20C8zF13QAFf9pdt7UXgLNsAGLOpL9JsWIq0xUQQGugBPV2HEfCyDbRLt+
C51aoH3i23Am3KAofUErr/bgCpg2hIuXEHZXdHRpuPdL3IiTbCQle5R9ynRl
Od3u+7xpLXWN5ueFht1oco0vsjvt+5Ym4S/y8EkW1ECexf0rH/zPOu5j8Amy
4u7U2hhGd6cMpfGB54pBzxxFIu4KrV+Gyl7dxL0outq4Ae8Tr5DVTrKRnAd8
6twoQ8CgFtTWLTwZG9vwk+lW5nL3a87tk3aFwVtHTBDOWjvl1SH/Di3wJVrm
xoJLO14q7Te7RoxtUSdj55zM8/idh8J3W2XQK6p4pxGm7CLF7W+ZAFW/Brb6
8tymKlCiJNvQ8B6zbsqZQHzIxqU1JiUE9ETJymQXz21bk/815qf2hqQSvKOM
KCznfz8N0G2iFIuGS8HyNb5X5aJT2+8J12a5uEvzSftbvMwNfXmkMV9pDwW0
A3LKqkubg8sD0joHgmFH7nb2vOPrHC2FxfmFDf2NoyE17NHpT/r4BNJblJx+
oVCfil3DpekC77KtfDT36X2ZnJB5n7zchYaoShtvIC+DkanxN6ARO/Zk+XSZ
ew0TFvclJCdhAQv6xi9dNo24KKvSINqOt4J3NBy0vqSybHsf6/223M85coTV
bWyXeyjmA3XgqYR5uNfsU1NCPP7i+oOsccbUu2OG1KeFo7Ym1A7PFRH3HwZw
EPbHPz8XnxUi5Brx34+5Bm2l+jGIRq3nBdBa4nCO+5wSvR/HRlI/Wb94D5lX
2KbbVrV9kS8HpTEjsVszDwmhiM6YGfumT/m1xDqu0ghrtHGT856Ylpc2AQrd
dhYb/sMUxq1lEgavoIqQuxxAlqPT/knOEdUgvEYI3OERAAL27/eX+VfFbias
3CjanmCsjHG7txgAleAhJ+xhqqE6r46tWQaL1e26Ki7CC6NTeLAq/RsI+s7o
QFSVWL7Lp0yIOdb/oYGiptJxFup1n7STy6vWB3AfDZguRThKiy44serg6Qfl
Y6Qu94oGVfhQ/Z2dKtQxoW7RVKRtYKhZVSej55Sbi60xK3x+orUvVvDzCj3w
2Z+ErDIAY1JhJZwXOz1qQZ1uAcOvitvawf4c/8847cV3D7z8/1+ftke7+y1H
eHSbbrq5ojHh6kCNIyM4kiSP4RnMCxlvKJwhB6+Ju7cpRWaVJIMUKGT4erFH
GzjFikVnDUFsJCbUMrZy8FvaGV2Q4KTrYN9Og5+38BndjWbNIXgp2l15s5b1
n/4/9eCT6BnBd2WS+DXQKcX6IjUfYlJ9/7t16bzk9uXAduZYCGo2E5ih+klB
wHI/eOo0Nm72fn8/CxAgtNtaIJLMZpcmQA3Ok60d6K4nHS3zXHIOBoe03GZx
BlqzT4HV1WgJdk8n1CEDxX0llNcPqLeLbLzHzJCUlrYnBL91QrPuPJbd/e75
A5OtZyckLxcQfa4gfZrMc8nFOf33aTzs9D/9qumyWKjhFc+q+PhsEjmXgnXx
L8Ha4rrNa97RtCWbcxuNYKNpHisymLeHOiO7iYc47aLmLj0kxoHksYnH5kyl
/l3HFe20hJCkXo16dGeSceuhBF8FoWk2aDHyhqWGHseOqJ5XgI/nphM3EMzK
2OZev1ehhjHNOu3vnxEq0/KlLJmLDd0D3/Ym+6dnmjeh9wvz9dsmHJsQTcvb
MuTar9rV7a8GjIeWepk+qbJPv6AUgCtJfoqwLB+I6IFG81+zxXXVQ4S78Tgl
jrVDkQ+mN271NMZG0tNsYceLxFUSUSwPnfkX+FW0vBJMHUQTBKcOUd+Lu9Wz
QLeAhjrAoNRSLSUQli9AB369TrvStFeW3zPbhG94X0hZzVZ9DvlrJcPuX2Y+
ImCDCPKVCjus3Y8mciQNCp4SfR9mJ3GfBWAfBJ8GuOm1JmajjBfoI4v6/Wqi
5Q8nv8dz8ssB3yxiY9Y5e7xxVtsg2ZDCttpaii43+4gr+8258f0PDKWl3oGr
Slvbiyahtp+uGUSUBJKJpLJ8swPhupR7UeRVvaoapjJVDGw/S2v7LRgV1tzn
vP4SzWk9wl1GvJO9i33dKe+Po1FJkxNrYqJPIOK94D9YzvZi9rfkAZEM7PGe
Y/hs5E+5QibqduynJIaXjRxWTjJFzJ8wpDF0UiLGNn3sEo1WcfRKBBAFRNUu
gJpgCaWAz9U5ZpxcYjVJ8cwSupmgQQcBiOgDAD1E0lVYj1owlLdPOHds9WMW
L2qqvnmeLwE3GUqb70U3EQM0Z3FEUa9T4H8bW23TdKpkpODLyJFqXr71+vYX
XGJXOdXM3dlvzA1yO9TA5P7EBroSNBTQ+GgP6q0k+smEx0vOvTw/6Ftj/w86
UIee5t5283+x+baTGAoV0nVl7iVrAZJFWVs0n0qHguf+cPdRZHXwzy8FSOZP
fnoIw8pnSJcvWh6ZRX4mnHMCC6EGUzq0hvJtYzsbRy6U1xm5Wa3pditE30ij
FWxnxjXOD5DQ9mBld8WdwAlslRFA9DRKHRUyD0nHhZebbu83VGFNQ2Ez7s5D
GSSfqmjYO/JZx0UEwxGWYmOraE8JjXtjraW8aj3hvxMjWb0mPKAAjj/+ED5V
wvSz9EKIAot/JWk1LnRdqBITi6Oh7OVQQXGNYJ0r3QEWBqo5KG/CM7LL83AU
5yU94UOFOkdmJDnizipNPEZb7ZBq2q2wWpLejTlXsr0SLJpSikh4TXxbpS0F
hdCcfmtE9k12USDlCyCuAXy8qVaGdDnyUj5OP4ti7IDMQIVwDBsN4bFMDiG1
jxCBWd/bd5+2J39hysfwuQcXLIODwvFJCtqOzFiGfsO19P66Pljb1syhSZ8Z
+Y+e5swc/N2YuYxZCWJpGwsOr9KbJ3lPNICAfZVcmYjc6Mea/5mxcV3bmxxB
z0oQd4CSetC1cvNOTQuqlaZdv/U1Jh9hM4xKAYlraou5jjD2kerlGQWncx0t
CtbdIx/L2YAufecGqmicRiI6CC9vHSlPizEFgU8PHtyh/3sb+kGsJOTIe3Vl
P0kfB2GsOTD1XQHPJeCfhtZw1YeGz7IghOnBMtdfTUS75JbYlKI3j08iUgQ6
d28QKiEvRdqHxJQO5P9hSQzXH4poxa4SUismXVGciWhLd7RPQGMlxAeAY8xn
BHnLGbaxxJabyXzNEyCcBd8trHxD86IuFNPgtOlWw7bmAQtDA2A4qZulB7Cp
UC1h3uiB3qSwKc92KKddrhqPywZ1bPsQp1zXl0IsQVySYy5qQEvMQ/ZECEzm
+A3z8Hc9dxUQUJG2D2PlmSfrMMrAUWT2IPqyqvuaWsyIpTkv0zlJlX6Lw5xz
xSnTMDjY6EKl8Lpk91I2ifI90N+RM2F+fJj2SRprgI/a/Nf5jV1btp/J5O+s
LAhtVmC70Zf6r18TpQ1/YwCh0tKf5yuzpxdFZyWbZHsxtZ5AHYahAvJq/Z/h
WXtAaGfph63hy0IWobU4BF4t+eOqM1K65uWip52IdP4U6r2tFTEBfLrHczUp
yeE1Bjzoq0ypiH9oxtFKlzWRoudg+9b0SHQmSb400Nzib/qt7KqweqaOZ+VF
cqlFQHjR0JX/RoEbg2QD1LuFZeP9ftzg7zzIW4bOSDDnv8ORQFlkSCsUOkvR
lkeQxql0BEYnESuDm/iYvxfZIRPjpllW+b9w99ZJ682kfTsrl6bqJSOv3y39
QeBfNXpWrnfV2p94jrBee1C/gnwYdtI6jI0i5vJyiytBL+K77KYeLkvb6t/m
2CfPQof70SZE0kd+FESBeleFt4Nr5d9SjzM1oEvLlsUTiVHvmw7U5JFLc6pl
KpliTGQAJ7Vc+V3TIVD1Xsh5eb4pj9jSu3ogfSZ7QT8pJwoC702BG0u91MFF
RIo5MDbpBc7bw46fMLs/IotNkkLLzk/Ckhrr08/wsfRM5v7oKOT+TeOG2FFB
31g/NK9zIcCTkCwQQo5fwIt+odA9T1aKycRaR6Inob8XDclZT/ndDmBCyAkl
BdBY15tGujc2DHJEaN6Y15yYBBH51ofvtSUCDqe0qUO9/o+cSZ6M7Is6B85x
y6YFkCUPhJgelaK2CleVyGzDB2D3qx8j5lu04uRqFbwqDgSa3M+ykJsNiwfm
beNGbhM1uje0knDoaQrvP90uVVm//CXuI0Yylp8iPWPDyGH/UQFpM4FmvrKE
Ka83XKLm5Hrlshnl+cbox8SBtfGVifiuUdO0U3kP9MAz49CjqyGZau4fzhNq
64mBsXtggCyQwGvm2LhQzvN63J1aNTdh3AjAwjI0OMQYhoPzJTqlq5X6iCN1
ki9qD3j3OCCYig1MIyWwkKg4CEURuft2iNzDDVswIrBo56uEyf1t/Olpfsyy
+7C/3sAtCqx3giPuibCkK0Xko8nd3fdABUpaiZmyucZYrAx/rSermNswcNwA
aC0eYe6s/xJwOQjlM7jWHCXzrr5811dK1Gith3a9g4cpiM4rATYvZsGaWVSj
p50OP3UaMAY5x2aVd3wMZ6pkGbw2aFPyeQjB87hpt2/3tLYvwTJFQnGG81bn
SMu3bb4wwugxOrjDhhXgyZsbz5U8iu3gdigaPw0TxP3l1DdGrtRURO7TJf8h
qu+eOixNpRCF8rGv8bda5aDUVxiP4wzV6ogm5IberNBZ28fwUns4yL3+35Fb
QOPxy4PNxANCpHGc0iO3YfW9q3jLAUrB0SVdUE1l3xd0EsHuc7+wGdRjDZtu
3rCkPJq27zz8NR2yAM/RyIEh9QQvRGfqIRKnRkfA8QZ7MHteSYp+WfhFcLoh
dcrOzBCg4xtro5PF6n3SNXwqzkIsZ1VJmR/qJ1YRGpf9Gp04VreyjGmeEQz5
oczqxxiNgHbUGK0Msoh43WFsaTTeQXxT4Cc6/IbitcyXDoN6DmmQxvxQaF6g
vQjJEi9lFAkdLo/qjdH4fqgfEN/apgOlb78H1XqiI1U8woav4KRCqfaQcTz9
aJch8hwEreyp7CP/M+FjIvbXfXjP6unSiN5B3cOS92+0K2VrgE/Un3cMZh+l
mw3q7Jg5gRjSOIGBVkLaRWitZ0xjZaQnZavNJLhOg7dCLSoADlSHl+ve2Ozj
q7Q1da+q4kYjQRw5UgoWRCECqxeEgjzBS+HkX7WsfSvyFX4eGoTM5YW6PX6V
eQ8Sekx8gspbiYA/zPyjpTzRxxYlSHVismtEKn0goIpqZUgF4wVOhJxNY1Pk
wkxqci6X3F8L7s50sM1NGyslJapLEZk8TcCMlzbhrFGrPQqpAVaAZBX7N4z5
roic3LcFZF2d/v8FPhAdpTI3jBRkjq4MEUdkanyi6WY28sjeagt+KzdjUiL7
u5aY3TRy//Pr1+8MCAsUBdbtTDM68o5qJ7zU6XRcF1gjcQ0+LCR8Pt5aACng
Ex/XZEpuF3tPxsCPpDBWpE11SoK7oHLaxx3SL4Y/GJtIM1qVP9bsAGs9+lEx
/HQvtfMItumBKHXlos7AfdW7f8m1H6Q04f6Ru5zPpZpdco1jULWpneJ0OQfZ
Ej5OCTKwzrhYaZW7AciBI9TJgRR0hrNtN1/EYVFYwlQQJazvSIkt9hO7nN52
MXbPbhL8xQMf2SaFY8XTzrYeGKiKav+VAO7d1j/YPfiejyTzfVsavMeXi16/
YcV49bazdWUodtu6QqnGzw9ruQJwOKyQOgynK9On44gi+UYJhMMtojZ/sw15
/GXRTwNyXGb+9bM7LrAIOpY6oFRvQmBG3qvE0tvC7cZQYHmjXvmEvTAqoCfO
+8ErEqmxYYv/kUc4a+q+pxWxy0offKedkisyxhk5oiP4T32fMciC7D85s54o
T99KeqwEYY6/qSPx4crjr+SeZEL5nvQ7f0vTUqlhh12Svyuh3YgEr+wFJ3hn
0R44roatSE8chn+SBpvrX/TbGDoIqTjkpR+OB7alJXL1H3rYHpHT0rUNOAF5
kGq85cxbTYnB2sRuZIhDEnFNljx1YFy2db7l9+/xLVcDtoGsHqKgKns9UYT2
3/C53mvQ8bngTQxoSkyRuCRnbxJS9I7Ji5NaM4zGKMvAFAxDlYMF/WsypcvQ
LUqnWpWz9CPVqgzRb8j5aMKdhpQ7PTBmSmA+uCLSv3VK9SMpmarta4o9e014
DAh8tI8W07c2VWiT14pIqqGnREQ6XwDoH4QN5RzArRaPLErPm7anrsbgY3Wu
Xb76jvnagsV3X/FcK4SOm9EnX7BpLvhYh6KnG2vFtoF4BPYlu2a/KeqNvM/X
A2bytRlzpT1oeFeoinzjs5nxNAmSNIho4K7QVYzqykCTFSP2zEstYJltmSW/
ARByDE/UXMZsaX+NWQTCJ4MvaxaCKBrWtwHq8QztfwL9YWGuSyiBBTKjo4ro
hPQWyI2qKOeZIONkorltqZv8hSFUcWINlfojWHMnEVUAEGUgCpYplib9D0CG
cLN+FaZOG5hu+btJrrrWESfxaomKfrn6lOQyWCghZ1xnS4BzHQbrjMvz7Ykh
GzdabJmc6htdxCu38izi4+wy6I0Lho9rEqrXWFe3UyLv26qOJ66HOTm3ARs4
XN5bYG2npIlqWAnS85RNHXVn3afN7UPxaH18uLs6L7nqrs3rDK8Yt2+KTAZy
kV2N23Vk5LVIItNSzV45127ccpQJSX48tBTTksK18d2EaUr2rZF/5uTXW4rd
1ETMsYhetslY5mL3tK+vgpab1HmneadhtodBnD/EF7bEfqKizChZrw/OZRey
I3hNlpN981Manvzqbx9HP0iba5VOInYwaJjw+jcPUMJ1ZBAQSAe7lPW0I11J
j9Z5KTJJdM1URm20T4ehrCMqrou2YOZKJlwaykitLVs+eadtDXkMNhKFhObY
nkgb7bBmQoT5nyuDrS+aOhz5vJWgy7jOtozvZQU58KKO3uRY9/jLkKfnuHwt
Eds7x+acTbZEqcZQ31MR+/HEIa/5JOyfSXX1z3IrAfA6HgtiNjd4IQFdO6CS
D0kUrkYFU89StfASeA8RGIUETLDum171VLdGKBmo2JPob4qDgZohBQXeKxAy
QolvrQ2w7ezQIl5KEchJt+nAcUKTnIZ7xWEfw3++t3/S0iOiMARD72b8fmTw
VdiKNry10jnNzkJqMudRL05fYMSRh8JRuDXQ2VI9UB8Ms2WTtjT7MrLSNECQ
PfidvoGPp4gLX8+2lc3wNOthCHKXf8lWMYCfcDCoZDrH/f5np+fefCYTNpRj
KDcHW81gyZ+/HbF3gjNcHMNcTRL4nUnpoNrHrRV8+YNtJMdygRAZjJFz7zDY
Q7aLlIhBc6UHCUFnVVYAUj+1jqAiTlcIOOhSuzRxh+b5Cnz0icts/d77zvKW
/UHzU4v4ZEblMjHWDk2OSMIoY3Ejzs0a1sQqxXGGJz46PMZtnVfcUN70enUO
pz2oD/+8DjBaGC3WwcjOBMIgCGltQLGkSSID8cNCjMstxuik85zHRbPzVwX5
6fd02w80TTx1W5fulc0YSDj309l+0Se5dGXWJ8OL4f6oJSrfGIjfJeonBSM1
jNL//yAqnLBQTaeu8MVCF/68GOfS1oKpsEgVniM9RfV5OWhU1TKm3SdK5p+u
fVmBejCchzCVlw4AcRLNrRmTSLlhVwF68nvy5i0jqfvHgpotr17svUWzESl9
qbAd1cpLm3gKhnbRSk411KC79PrkilJ9M1zUyu5qPhyNlDXZi059x8wN+jSu
GbCGQCw28OyLKJQfaaruwsl3exhUb+zSoSla/bZl8L/C7PZ54C4KaG4/tmqA
VfN6HUZ7cdmSgwQfBPLXehOBOgGCjHI8EkXodvrmkpOdElJI2eWC3DzfBZ1i
qkGE2iU9kjqjJbAsOW4mekYS86OgCbkTYh/Dm1/v4zuuNQCYvYSH5W427gW2
MnyqwfL1ldKyU2+ENmOVOxf7i9NoJwFY7Wd39xiC8JzpILA+ZZ6q7lJ1/4zq
J6cc5t9d8E+da8SgBBikHkAxuMc80dbw+UaGa+E9ANt/RO1ncI5KGjYQRkLz
6ryptOQx/2mVdK0iPT+tqbjmLvYezyHDL5N8WyLR2RYsAULHz5r/+HsWa8ZG
/8W5N86SR856vnnbaW7ndQVn3eCQSo+foKIwfiogO5kevNXBtRZQio7l5wAU
xrOc/HNinQVH4GL+D5ks2N+ISH6HRDsVmST7oj0FZunuIptI1thk2tXOz8cq
v/fV7x4U158hcbyhl6/wAds+0lTSTlTqhANqajArV8zoGf4gnPgWem93Q7iW
ZcS3RCo4BuAobGsUQ6wvCTfqhfOIgsUk7qy5oZKp6/Vj2YYiHcGldpRPAepA
K8VYe+25JwG+l2ft+UiNhKmw4UWMDe8jYFsIvZC2Lv928oqRe2mIT59UOL98
Y6uXctzc6SO/vW1TkF9Xgxmbn1gmmQks38za3MK3fHIOiM2fHqBiRAdK5Fdl
81XAz1dsKzcgQd9e04qeFsSU9czj2OT1ak3c6jPtimDKv8ah71QARBVpxwZP
Tlf0D5U9wIs5K941HcEhM31adcWgCIvqZSbrfueCc352UggXjPvRptEEnE6I
80hUfiipD0v4L/v69SWk3BRKcRSPNY2sL/ILisXJLQOgiBlj+FsUQObw4iUj
me2iPRz3vZM/zZdLNU1wf1HUR9fxJ8UgqBb3Ck4L7y3KQFKkZUaH7HK6wjwV
tw2zOA3Z6n/OzhVFe/1ZKP+q6vWe/yy4+rsu1YKu0FjD/1hNDkeprKZkMlC5
jPXnXYkRoBQ9h7OjRyg6zwKgcdg4n1CelJQ/i0BpWeEL3NOvZNzKu8SmnK68
Wt5LVcktcimFfoIKssyfrXiLIsGwpLBwWr3D1KdRrTFhjF8R/t1eoFrKkktu
Cw03JcPbqsjExcn3pf5f48qQgzvX7YsCstVvLQ/AeUcX/waaaRB8A0b0mvNe
meFh8lQb/fzRNbI5QHZK5to/d9SsLZp5Dzsa7feBiRvr06Y1ase/3U6jDo2S
/SaobEd2R8WpXXhz3czshEfWpsoYFK6jF95UTMZhgPVWxwNtkQ2ynq8vvhEq
ZZe1nUQ1vnAGFv/iFsT6xVVHbKo1AycUaTbrmYHZKrPZ7VKJZA5+oa3QOGIX
toX8eILDJiZAhye01tToYIAzIRB25MhNQTd9wqiOJk9vMkCIp5GNnauzhbYi
9Uxi8o1iOhoGp9vdeR9LOu0qM3uNpYYOO7GKnUY7QEYp5gBtzRO8GexfUomm
G7qZwRf3sL1/Qy++pYZnGzva2VPZfGxKXhFCWZMgCtCvjytPmbMuq9nrrv5P
7m7LxrU5lB/FD4tddQ2O0BTdwyml7aE977bbPZMTRtGj+hNUxrJBsAXgXn3f
zdHXSccrqnhxBObd7VIKUA4388RiBN51JlWGubbDxt8nHNkOx5GOSffouTf7
Pbk1HL3MtH+CZBMl/FDgE6tvc59v3a+jvWczVvigjE0GeE0kPaK4JowYLaxm
Lpi47iTuDGVt/B0X4JSJX6W0muK8SUeIjU0ma97Ar8nQw5wDcfAvM8AaZ2pD
cY5ifzvcQHzp6h/L7NaH/ZudylekkJmYhdAE/Z4DtrQRWi4+cM8eQymeAXVY
aFiCcd/oFbsYnFuCMejpEmTBh1Xn4A1Ivl7k4QqUhJwkxa8D2zpO9cX4xZpx
wOyek/Y6JoBPrsAwJGVSNFGo5vttmkxTONldBapeIhC9NHwGER8eibDLPqnQ
jzff94WzoQoQDx1wS4ui3Diwl4wYGTMSLK9oOXIf+vxWH/G9M1JtJz1YyxGh
Zw6/I3JMuYfQaj6L7AE8vB53EdYJrV9rDF6DVVIz/n1/16+9lGWCR892fZ6m
cd327szEXR2T/WbSDYFcLmBu2/xqCrIZbqJYGwimN5YxMud5oAVtOrdlHVJ9
x8QoqMqsrQfbmMDsk/2+v8Jt1PSl81PR+EtUHZ9TaTnNKlOWYY1xLPa6HUzD
DRFXSPU44ggS2yfqo4krDFdclPh9Aa1/Oejko4G6NGixAygWKofVpn4FcLwP
HHApoprve3thFscy9vwsrhMVodd2ik0sQefj39tAFHscWVNpMmWSwaMV0xQ7
XMxnVL4cUKLzrhSiWnf1Zz078yP5DI/ui/e58oWlPkLdQxqDPHyY3o+3PZBA
siaxfoml5ysICCAksVJj82P0tDNRWTmVVm22XA2L6L1reiL2XWiM/XnPBRwk
fS7/+kYIq1G5G2miAf5Ewp/NTxiT8qADkWdBj86uHfOhmZowWI3ZVrOl/U61
f6MmhXQX9f+8FMiH102q9qNNbRK8bFVP7wiuQA6AKlQuzyJko/nJPpjBiY1x
/gG/5d80rTrxN9Pd1l7BwXK8S3aGoldXV4+t1rA8V0EgHZgtyH2OPfZZLxme
e9KWr95s20r1X/j/x02amnRO+2YbIRtd33A0dV6hovyplVkgC1MAeVkDDKZK
a3kJpBaYOmA60k1J//dQwcGA28bxs+u5+k46uX0zHgKcmcZkyaZcqqwJgecZ
BVjIG68DiZkkqP6CIo5lFhWo/4V/VGddeCiJUxkZokqWthNX0QAPvG0sTTau
rUzJSOFqp5ViZAGAT2LeyqppPIbwT+Z1Y2jnZGRsfr6lSdsG9PxUI1U5LSrp
8XMjybt4g8cc4rU33G7HVpzvTc5jEmJb4Lsk2AJW9g+L/1WQ1B9QmETFRotI
Kri/qfJDv9XxP3k3BfX9co7iG2mNHmVaPutunGN6VigcFXqpOhUtvHOUsiO0
dZ8kaW7kUQW5kdHrzXV/9DY/EV50JjYrBnZWSY7clOKA3B58tKjknjhbmqvm
C+gy8sYmM6foWgiMHFw3z571KAT/086aS8Lf6t3v0w++gKyNeYlfoStqvofa
l86obwgeZ4KJUAq1mSn9W8EZcvtitZVP6vO8y3InOMgxEof+qmkkHdyxaXUU
mJBIpTk710HwmFw2OVY5XzzlHyQsYWjUUWj48P8y+CSubmxgrTz719NOrw66
lPMfuGP7MD/nqhAFrw9AgLs02a37or55BQ9HpusqkAWhu79dC9Dx/WxrReB/
EHy/HiCcvRJuElK9T2bbWookr7oC/L8HHIIx7UbPmVoTea9Sg71LJ7qB+SOd
fOydn0aOLdgk7m9rto2/uoVG3W29PerK5ysjwt+9mNGET8+/sb14X3uQ0LUU
FJSzBpYifXgIQ1C4od/RdDok48Ulf34UAArMVAQHI1dptf1ntasYfwPA4YwK
ymquinX1jDuSgeA5Oxou/srLpcVVh2AhcWrKyx1sggAVrVgYWnZduSgcuYWQ
YRTw5ky/hp/4/w2OSYN3vAMRdA5jeiZyborq83ORwpTpsimM8oDXTdwJgFmK
RB2yp8evPeD8a90yqZK/D1Ycdo8nlXVSMohmckFPavNsH77KI+9MEKDcya73
qh7Dlaa+eOITiGz0YWpVIyD8zObgq8zQMJsVoxPEPykSXZTCuyTxiYsfUQXB
UX+Rny2wSwJGGXDoncEl20iU8foYCfF4954htDf0d99He9o2XxIbIH+xyFmT
i+0BIpizqYM9t3fo57oVlvdG1i7piHBMswLiaZGDzBCLnxwaYy0StC4WZ2Zw
km7ZToVNQPorW+rnTPgEwxnxmPf6/LpnuEe2EK0XWLllLNJOnU8pmmeTtGIu
ulaPphNlYt2dUY05sLNThT/5Ix8RJVwk/z39Hwvt5H06q+mKXDnRb1yJvApc
ex9urISopojBARs8/z/AwczsheqkpSMkkvVOfcyr0xSL7MQmX8Cu51K2R1e7
u8LGzTgB1CVm26oZkmo4NHJNMNlE3LJbI6OepaATVY3SixtcGFdGsTM9zB6y
6kpmKEloOJJZyhHK+8b8NMzvSYAfDv3gZiqaa3tZcJ4B9TLW5AcoKj19V2v6
JWqOaZtu+TbL82BWpxrcrTZx5ABoY/YXGSri7wV8wAUgh3giefBVNMMdmjfh
MmTuQ8SnRYkCT9PlrK1rbtDARGTrctGQvsTuhu7lFNYAiPefWxJBIiyfT9PS
1yrrcNhEm2mryYX+mxa8VPiOZhJNZZV78syzKba7Jeqb3a6/KlMKJWS0hYyu
qEwrZ42viDlwQ9fXnmNCNUN0D6IpQDPAUpeEd3SK0z8FgLag2dpzn8FbrWhK
SaOwoGmvq5Mx2XdXSULozIS804yp/5lg6omKFyJQt3XUKZYi7b0wKAIoNyrT
LoB2Ep/VAkgEgu8p6S9CQPhyvtayDQ2grnuop8vMAt1DbYAPkUPuyZc742HA
f3vjbVneVDMRXMI5Zq1USjQQavIBWHP0JFDHJIdujSbrobji+qBI+iG+lHRG
Yf3gksFbFypDqd2JU+9Xc8XzgWWBn2dJd0wRzmgCVrxAVI0NyMT9aUf31srC
DU/UlLKNzOdnStV6dBJn19GEzRAXVZgeB0JkfKcxbAGFEP80E0+QSDvepEQz
pz4WCnjMg79GGD5rRCOCivpuNnGJ7xz8d+drTTXEu91SBh6exoWzG8DjbZQZ
cTJZgQlmFNE49iWmiSrb2nSZUu925LkWdS30B5FQnbERxs7kP1dGidr4bRU+
wUitt+Hr4vZ5jBKv0u1qpzhqS4iz6ee9xS/8z/HKuCyUW++lhilwRXdcNaq8
ur/gJQlCbKnrlm2tmQVzawOhoxB9Q7rxzPoDMAk3mikPDKQfWvfkHh3FWf8E
B0WSMrjLM49NGOLmOGLfKqQysQl5PjNLkJpeDAQP9p/ByNjM/25WushNS5L7
FBh0uVssd8mWPsZhVWCk2l/MtW+0h/2WBk7MGIabbsnCwtZOGLyXEh8jPu/G
OcwJIibM6CH9dOZWcmugAMfVIGLB0pgz04lo0lRrk0rcPAhoqLFGik8Ugtmh
I2GPuyUKviMoDluV3dttrrgFO7vt3UdJgEiYG+uXoDla+0eh4509FUayJ2B0
NVrbhEreWztKUt/mdNHeylGY2ixWsCFEN6WS/2JfHDkWZl2JV4IBSQYzz2P5
vCVzM7AfoeKiNTedejG2qKq5qyPAD9cvL80a2MMHtrSXtuyi57Xs66fyUJTU
wZQJfJW+MOwuW8SADAB+K1w1n96KDQkBbxu2Zd2sRvfLl9YiywSf7PP9N00+
FRxo04YOyvlDPsfyZZQ9Hy+IQMKiZCwHRjujZnSjcsT59vz/ThGI0+mKhPZQ
hqDIxzfi46HIbV0CHiC3Zxcziyb4pbwwZXDxhDe+K0q9JFkFNhysOpRFqLE5
2QL/DFf4XAjmGjmpfvz18KhZK9deknuOD5NyRSpfdvxxJEB3lp4s6hjMTHrZ
73pDQbpi8ROZGZL7Qo6AV1cWY/AxgaYM9vPAjIzisNz1bpDHwV3l0YMHV2uP
Wz/MXMzbx8CW6YqhURSDYdFYcrqB4zlOJpKElsWHsz6HdUxkaW8NjRPJQKC4
xEtqwOezvetoKkf8knZwlbZMsuIN6iHDYZWOvblY4b8ctVNo6RHGVgU5HbLv
XR3MN8jVw0v8s54uzOFkVUq6bik5z4gikAIMGl7NrCeDK22ViqojHAwkh7K3
ebkpB61xwA65F0qjXtChDxASXi5hUeLfAYyyx6A1138rt9wJDOF2HEGnqf2S
w1VULuT8VKjUUotTkBW8us0jFqPhGD1QfuCtJHzCbn85hKPKOrFYzMkHVPPc
3Fnj6c5Zk63HH1uDt92SoeS0TZmV4gm89hM+SSE7bW4TvOOzrmNF7kK/znrn
trx/gNXye/oZ6LHQPgpx++TAbGVPEqzWeUTOmlABj1GJIg9OlUXkq/VFc2l/
dtvpal1ayn1BAL0RdSYHMDMtUIN3uSzvOBW8AMts3QCYWOGzksBjPHI0Co05
BaycYIyXoe+VDZ9sKK3GP1+7VetemD4s0gQZ0n5OwRqJNobVzh+lH7GZ5iel
WU3Cjz63D3YqVSBX9LI5x2DqlWCy93yArIQWvzPqmv/x1bC3Iuox8RrTm102
X11uSGSZ9ya73In7WOa1EjeZGIUzuhA0JWS4sxADmpDympGjbd1BRaRShTuC
cWHgK2CzEWv3xi56w7WXKV0vRtfu2MYYlfWtA9ZLMSHeLQZ+ZmjwyYjz6kcy
8Zinh0xU6VkXS0W4QUNzg3hEKB4ZoguIROKo/bsYH1M0QrI8JjcWODQqvUtL
otNYtu+YTk2WfTnGqd7PqFCTG7BVbCHq2P+22n08yPYSexbR665OQssrOhjQ
yg+0a14OOuPQSu2vKVvT3cGpD7/MqtJbc1NXxd0h31hIKWqxo6fK29zMHwP1
JgS9Hb7Di9lEoAWdTKQjPxmBWV1kCFD8W5CIWqIJaTdoXUaBpfKFz7hj0Np1
9ZgkO1zJsgZTVRGxS3XCq5lZ+piMf0pGD7/drY7+uFyN2fU9v0kkyz5kToSv
sOHyHbCN6DdecYhMV70EaJpPuQtAQtsImoe9yHsaydBZP/yy0SFWlcXZGWL+
hWXSYdfPUslYlCMeRiTgXGh+lThE9RzN+Vbo5SCqQORQn7Mq4+9wxtAAXj69
gr37Km/P1FeGOq4sduvZksMq1nWKKaCZZ30sJPZAaOD6fn39ro/pPJNK/gKY
L3tPlAi92TXA9TIEK9M2T5p4rcQ+hlPHK8nMnHUBAp6vf3prqyLj5HzrNcR2
RU8LpGUv4jtNmQwZwdhXNqwV4NiVVP14SQfJIg+roEIPtZu7hpODNrjMchXv
BmXfN/7IIhcM+7S5fAb5jYLNUD9/ZxYzu7O0BizhO/ReHD+ymolPLRnoaOXh
gT99Vo7Dmgin8gsPXVJs8jqMZrfpf41BWyP494PyRtBgX6fhSZMUtAo7GW0n
1ZpmnxFfwDKuRtNAbY6GIXtydLm2x9IhX9NJ/rOKsBNu5tjMX2BCtpXn5Y9B
yqsc73mBHH5ojXQ7VDDRFT4Cpd58YtksWGLBEfi0YGgatTImew5M24RSIl3P
bJxO8OoVYKpHI7Mxcua5wz65g6xrDDYzDNPqut/rLqikS9r+WKJ7NF5BMf9s
/RUAVGmVTBYhPNfTq8MOFoiAihdu+P9rzQpvhVQeF6OcEXipz4LwoqYYu99H
lyhdwngwJciJIvdU4tNsXbrhkQ35QA7bjobnpOfrdEjiyeF9rIHBjBKQG5yl
fEHxNj1hEoZ3qHOw4ZTi3kelcVCBsB5zecqom5aPlKBP7zHvUAGBvlfIS4nv
dTN80H7zXBZQrvlPEsewqFAHJ73asIXfyiU+4JNhYhrewQNm3t+Uo8WzeDCQ
i4rozxpAQnPqFczeo12IFi4lDCoRexFwTj34DjuoilF8Q5lUe7VfNwneEPRH
HjzEz+bvrHiTfqyigKZ2Sst9iMcne5GG9Lcg91Z0EHifmiT0Zo6ponR1UXVF
jeSpXyDX8lFw+HZHcLwJtFiuPKYXCisKCYOYg43EwvoQLXmKo79/iPXvXn0E
7Zr9ctummqpndXahIjaPqmUQLTMxaGeVkK/mHn9EbDhorX+rFGE0xQ7DRDGu
b2J7g+cJ1aGCczuqMWssrE1dcb/3AnMuvRJvacBvR+S0Z9ICMrT2szCOF8af
yXLtsrzqmuDJWvaYuaffwRr7T3jOhuBaD0kvXhkXNcx0FcAbqlGpfBu0UFns
cf40p6CrQcUVQFPTgn+0AT+zMvoK7ZWC4yqLPIw+P4v5pm+ZgMQxBY7rAIMP
t5b/Gev3UUhftar4Go6CTztLpc3S6t3gjI7kXxMxn/3g99G4yllvzEDqbqco
DZ+QAezflfViJzrP97e6ayQmbjqUjDwp3PhtsYkDI/sd5zgSdCyNSxDTk7dY
6DXdjX9F64Q8Y/KAlVSkKfdFS1qQwpife/BzHmyiwnFqeaffOTvpnHjWyjuF
SximoAl4I7YVku0EKC8oSOXzvQ9w9ZVtsq7yhkQe+RU7FShLahi0sn4h8oJI
ohVxOCyPdoowkWYrR1dXy26nd2rXUUGZ1WNb2Doljb8T6F/nHKwN5+8739eP
4gGMWV3XZXvFlzQJYTwn6tStamsuf31nopxcPs70xdjf/5r63uNWFm+zF8SE
HVVmjTKXxIwF5844DSj2Iwcz5JBrOPD+T2VVo3+W+YR5eAW59ykqk7ijDRXY
sR6qwSEQG9xH29nt73ORGLT1Fl/R3EyxBiUjXg91qCPfA0QE7n1eOE7rhuyz
qCIKcOhHyeF80ESViy8uQt3r45rOfdDPKnaNB2aSyQSbgTwOCRqfdLDNl9Pv
EH2v1hJgOpIiEl4WFtWrAQ5PxjPRdYAOKwS5P+Fda/Zwzy3hIQqOSJWxYl66
ino4QYgsJU+CILbErDtw6egfGiz9bJAoVoiBBWmHmtzF/yStUJp0zehajyIP
GUMm3LczINma9QcOtI1LHGlq7QxgmK05sS34JqitRAASBdgqURyU3iTcENFK
4rGORcWAU+tyOpKecNLzqG4bstiPeJP6xNVPCIu48vZTV0M5urJJVLsndtOF
wJOnWb7Yb+FfSuDXIDkqDcNVOhwvkA/evMkBHXAmPH5vJabNoEpSskaRekK5
ZueuD/op9HBSCxkHkQTKmkRQmrl4za6mBmgHpl6TqBeuSclvP5EVggjARDVt
quRQ5koPZNB4J1dWSAdP1NKw9lKkO0Ub4jAn4utsP49V5YKXYdVNfeUzz6N9
kPfUmq90AGwfPpgW9iKAYP7k471gKOM7oz2XLZqZW9k/5GyAy/DjwPl0rmsi
Tn4qqFsJaPXChWqPl3zatK8jigW0dOcssV4VCVm2KkZqfaE+i1WH8GuEtvuS
fJfZfRjTd8LTmf8hdQnK3KlD165OrzNDbMtGHyitetbCYOEfRouGFrB+jtTl
s9Z+1qYvk0Ii2B1aZCGMGpK7+WQjDRAUHEDsadO8r7THlr7X87MsebMHktdq
FB8dSDEnUrWLWP7m988DELiWx0LKxRbgYPEt7+xKr8TifvgWUDw9liZMW3oS
oj/fxbXpo9VHJ2nEq+wJomoES9aKp2d64ixL2IvL7bQZb31hKDI+e5jMBPcj
a3lw0tOGhnYqBjwhhe1K4WZ8QRonpwnxyW9w7xYJpouaZ43uSxnJBswMqgcp
mruwT6J8i/f/lx0/DZP8v0NNjtPp0VK9JHME+IESu4fzjL/w2dAudSTJt+ip
nAXNfd2dx9u2wFmsoCBiFq3mJmFD+uKEq32htbpydJkr2qnYOziIGRioHUOQ
mTrpHrafJ0/H6PoVXKkrYkuCUeip16b8TvP5kIP9xaF3+0mzrXWgYTEwOz3Y
Swq23Z6szKuRMgR6OILojhRpBvjXaA+uk+xkA9TuN0Lc+IWZAR2Yx2ExPRAE
2EvOfONA+cKwFrTWj1QDXDyC7f4Arl4KKDe8/+e+hImIQAMh0gdIYyWTkeOn
Rg+1txDCI6Lf7dlX2Hfr/YBbzOM8z3lC/ngT2gprXNHlZqxms3AWL7ZN5UpA
fQtuIXgYnvLt+GoVIXUG6mg0LVktWOm3juWtO7pX0wGnH9nGUqL30kRQybsl
1TYtI/LDgLaceJvP9DZoe/AnZH06URnQ6z40dOkEUXCdmXK/5Z2nRF22G768
WxSWTiqtRnKbIcCbTMBEMkLIhHtEhqFOweSzuVC3GEW1kH/1+gQoTVz+CsG8
5nQH+sfTQh/gzwuhRwJ4WnEBDNwg/ohwZNhwugXIvMnPQI/33XrKShDzqH3r
P7Od0rEzKJmn09mau/8IrhSJgutj3Xd6Cu0xTXRhwvIjqbzN874kiFGEjsHx
/oiXcEeiS3hNFCHTKEzRlvQnR+X1Fcw6PwITQlzfGb7wn1q3kBv7yu4knGkn
2HEH9qLbRdU7yioLqpbkS/xsQyv5ay+k4e93xAuauwFcLimmI2Egz0ipmXNg
7BstLeMhAYoZqE8bbYGU2xOW6wTZ+s3njvR+5iQMKrSoWY3FNeEMwfI6rqmC
zGCzhirRUdIxaRT2bBmadThRm5mMjG32EM5tDy/0UWu/0UkbF4piQCCosMwi
09ZMCa9pMEM3ghF9riwjpIoW1pfY/n10YDCRWTgTNzxtPfMObPUcwNE2Hj30
EGi5d9/6NZ7BuxXw0fYTCjmqKEn4bU4Dt6iO4XdZV/XCFkC7/GaljwoQ1wf6
dWoj0GHByqhIeUnyACT3WD1iwj43H75egy+7XM0p9B+1N6kaaxsFqoB0NX0z
oVODmcd3cnDFX316PfS3PWGPp8ewM/ZBHuL2OJ4eXafGLhFaN7EqRJMPwhLi
cdmm54teQYXujSu5b02/lSHmqDBZc28f+qSRXYIRfQlnMffc8T5/FuOvX2Av
MGOvZu0+seBKLW09QX5BMimd8Wln8Nj9LgJwGbYlQBDR788HO7ShQmyPTd5D
lz3Csp25hWg1sUm4upD+GxB2tEVxSCmVhp6olXUnzQCGHWrGjv+I4fZfMVKj
yBzdSGh5/hpzBwZF3zG5ghWNHde1rLk7xa1ShbNDRzVMTKsi0020OqLIlHMP
gfVVuyGAo8J2uCGdeQDN2dEkUHLwegF76iHAMElYjks849hk9RVDpeWmAlLj
YNGBqys8wnL618QxLv3lA5IvjP11+qI2fVQ0eUQFFv3CdnY/EnJnrzgqlLJo
HOdp6zjhaUF/9oC4VJOxxCjrunBxXnIn/YxHc20+borywCz52+aKd6bcHkRX
J7nPOQu0sXvJaCa8UNMx7CylcI0ARKDu1FCXhjkLwY8JCzzx+hfNRJU8SbMc
PSmqMj9pzPLETEvzDPsDVFSLpWKwwuo+NcKs1kjvQg1LSqJvZwBHyAWmUmg/
1gViDBP6liKPGoDcAbfEBv458bXv0W5LuEokx7BkUWV4/aln9r77IH6UgZYS
Qxr7o6dQW+9i534h8OqjB6jtyPHPRnIUDQ51+yTvzlf+yX0owCp3tzbegtLl
ZMyFfiEBWsT1bddJeeYQflGEM5IyZQOLil07QlX7MJi9x9wQbd02b8ScAvt8
zkKKHcefE+S+VLGRy7nPYioVroYTEosBIlcOML6aAt13V2qkVmYHtJSLZNAm
fkcFFzhrrmgZHMduS6k+8Eq2U8Cv6/GmSgJa6ehyaiS6ytLuKkjGiKUrxk6V
gRRYREH+ZVn2wrosi56lS66HoivKdJXmzQLpdoTiVQv2e5WuWig+Xofje2Ew
mwNKLDZ+36C500cfGUdjgPZdrmV5XbY4fJQQmn/9h71xkvdeteeKLCuwU4qr
hLpVOtgE9i/FxBzKCfPxTZrcLGLzJDvLC5iHPPZZkXu5LUH2aMr6f8l4Bh/f
L8Tn/of6rnetoSpeQzfpm5BsNq8sSxd2nHSq8lAmqHroLXeCErMPd0q8EHf6
0XgtcQKt2O5Meox5gjYCqZzpWpviNXxXwAWkXG3VpNljww6A5l1K8ZCAqOTy
o5KBoUemM7QaYqi9bL+3P2dRMiVRHO7uc+I4/XArgbWMsY9GJWCtykSZ+rW0
/sh90Pld9yvdUkWmMUxwSPA9XQ7qo4ooh+afcMMjos32Csi9jLebtke1i0Z6
AITmFkJ0c5Kej5ecJhR9oSKfK8Uc8ls9oheWnL+NaEPLnZPeHWzCVSWI4wgn
6eelinUQgofNUmX1J0z4a7J+8oMcTijnq36FllYEPj/4QNlDTXgEAMtRqxtI
gpZGqsrQTpJ+gDmhLhS46oEQcLXhY+/Q7kgVD3iY4bUHfpx+n1xiCg/bemVA
p9aOy6Fcjewrwu2xEYOMqsIQIGM5zaGm48TEV37QUaDZjNLIlheh7Um/Bz+o
qv+XHjtsWtdMjpmJEMLJHKKj5h3FMAVb4fThJ3luQZD0tK15TB1N7qcesjmh
oP0w6lBpf/QF7/ODwnP4rfAyxGibjlpob/BnW7jyzewNvlPyhWFWCExdiox/
QpWDjUJpueIIOMvOTfcNQHlJWoW7KWSCip34GMc/PyVG0z5iEaefrqhJduCi
1bQWGCE9Od1F//Bz0JP5HmlCfEzKQSSbaTyapUW45oCWZXNwBRdPhL93g6He
yN8WF+s2yY+9P3SSYGH8ddj9FERf/154sqYzHW45yqWha50az9a0iuuCJ92C
xYnt6kcHQ7IxQfBs/7jYl5GxU9DioJOsQ1V5Tb1tCc5iIPRYhtDUcWwuCJqB
uTxehiKLajoPAASBwBvrEHSmAYHIhkrXhZOMelr0VETtQbwNWij9RLA8aPlV
8kWuZ1qsQUIKCGwfqF6lSsy/Lv/nLKUcyLjcsw7qEqWWcDuvZ1Ur2b14wPPz
RvyVPiP5Q8/Q30aGLo+duK6wVkizEzVwvnQlZJ4ao8yoZSw7W37oA8gPAL3u
utAiNZ8JSgF60Bo+OEfMpWgLqnIxbyXjwo+KQ2g9YrMXvP+/T+ffMcuLeMao
AgWCrehj5htoRy1ty7guZ7WszgmUvfw3JzqEpup54syZAx0oR8eXu6A4asLf
+E3u6/2epKnWG5KGAb9+mSkih/+BTVBa9AHNuA6hCRh3e1FolYcCVierawgl
nOT69oRBu6JlxM45BIsu+Y4rNEylhGpn43tf1GXAcyAHDzgxEdRYDSDuoBcj
NVLYKjh36mUCQ0knrdYJka3hOBjNopXIxEk/JQ+k4VBRWOPNtXCnNduMtssn
t9nFoZgs2dH+CB/1pBBsDV6Xmn/xKOcuQ7H8Don4pJPszN3DuuphmTUnldHy
8b4RpJF8HYtLaYU8b34+yKAqjjZegwGePH2X3vOG67tkPN5Qci2O61zoNKaK
CNQrMeBKDhmjsMJN5L6X81M+osKdLKRojn98MZIiHu7zElwo+rdVTBpGBsN1
mCtYtrvB/hMgguaC66TCTHXueWn3ul2Lw6r2dYmALoZwfLq6MjxF77ixjyzc
mAn7HQIf6Kebmp8CsTnb2kgvREyDL2B9+3S4/pfHsWnRxmG+r+TizKVWEZPP
L0VUihqZERPrdwyAo7K3T6ZzmNgf4RFkz3x9GB9/0gEDqiBRjP1ZiCIvknyC
4ZcEuRxFzxw8gks2d0AlArmY8fblJy3QKdsWoELO7ICaDMXiFr3tMzSb6tj3
CgWadJVFkD+uG6HjsJkRqxXezFc8dR95U4mO0OIi0jKocLakcVQj9x4VNGfF
9GqKWLkxj8xsF7Vme6nW2TR2d5/JJ6O2E0OOWcL1khVctRKG3hwlIrrvM9OX
dyq+ECbjWolWmypuy6yakGFquwYLUc3tqLzQgg+Ux1JxsxJ6HEP/LgzeLA54
zX09LaBKI53wTRIyAsJDq2QiwKCIQoS9eiMvEu4+CezPF5nN90BIG+flpVEk
DFO8zVxJusx+4nVfQoU/JuP/M5VEteo7N5amYojMn8c2dmfGs6FXlwZ6SZNC
rNJ8BiUOH4by92oRO9soo2+QG0tihIlJ6+RlEcieJqwltKyflOrQ8CYeqyw7
elownCq3l1WREk/v4BxZzyq4ifPt/9zlb8Xdm5+xnq+QpslLXZLpdCi58Jw5
DlJQ3IFRf4yVGNhuHO5V3QJZwwWHbfBHx7d1nnXralLPtdr1HmdmVU0Z6kOL
ZdmjFCYDecrQVHsLrk+1Fd7cYu60yP8joBzDhP5rECmoizBmVoXUTnwRT7Qy
OZJvox7tbt1tEreqHzXBzXyZhb97zmD2nmo8VzD5qU3OI9tvBdw5LHo4b3tq
MfVIOLYGbCt7LoN1Oc8s3OYZcHtA5AwVH+k80dI/JdZaNlLRP4e3SIr2lH31
iKdCFR9Ybu6sqwNT4wEW4AxL9yRZlSAnn6RtZLqoARWzrWqmLGt8zP57OETJ
/sOnuN9vmxds7xVLwvAa9l6LPKocbWQuczVjDyQRSqvExrqWVdLkg4c9RrIT
DQFvvV01/bnoI9a24VFRZFuDbcl3u1nw4TX2vwzuOEdl2pcFwH3FI6jlUNPO
0gQQrILnh7Bt4bGMzn0vCJxyENRnKPl9JYB/4SxiSmT7XfO/JbbBmPhZNOdc
Az6AWh8mwgU4aE8ejhWGbWBLXQ5Xoq9lKOz8PetN2FEcOojHDiYWBnsOlj8L
r9JaKt2FOOj+qcENwsyEcH7qBYfZuQDAozxs4AHQdH1B8FUePF9XWk5nF/u6
m3bEo1rWASctdX288dRNHHpo62w49FTPa3XqxeVyp8cwHwJ6bJg7bddbg2UQ
9sVFLN1d9mmAU5+RBPJ7nhiNABEzdFcW8KiCIXaCobUI7tzLQ3igDm0IddBe
Jd3Ev52hC0NPTzYon9PIzMrKWte8G5xjgSAj6mHi5TGtCLwPmQ7Knmq5ANBe
Cz4ORZMkunAX+wXnB4us9T3H9kLZ4vlnGySn8jPXc9ZNzigMaeyyjgkoXgrz
afswyUucVRDTIWXpx+JkP3/A0KrkPdAb4HPjKxsVFZ05YibITZjxGaOnK1t+
yiN2T3F9q0eoa5G0eteuCsOavkI/Q9r4fLg0yeW9bFPIh0tu1XekbpWm4AnO
bRB9F3YkRZLYJrO5E/C1jqXjeKPu3rBpKn9QIPpE5ujfj+xqy84dN/iAhxOt
XRCOSyfi93XDrDjeLqgVGVks3m3EWolQDp56M3XRtvz6grDYKKE4Xa54KO7L
lgDvlnnIt9IhAmDnQS2fH2bYb7dUMza7s/RyQMYFPM/o5VTAJvimzX7A7G4S
IXSLoi3Yc4QDkLM6AQ50pqTDn+KcuNzqvWkzS8/UOmxGxPl5P3JD/zrLXAM/
nKyIURF+r59StIBx1uNi671KnPxgFRnhpHkJvnh4OBg5D6QFGOWyv4JhjHHG
H9kyxk3PJVKfq9RDj4jw9LyyYmla/fZT6xB6zdSl32dOinr/1/PEsq8xMu7w
QFNDtfe0MDy57cDkc1fsOmrsow1zKhB+b3UOS63/LcPSkVCOyNwQsNF3LutG
qam+4M1wVaEilE9JJIUqiFM26t6zIWneZda9DR/Tgu8Nk7+PhGNfmXgh4Cz5
7Ss3uBibuVEO4pr9fCe7nk9fUJd24wyNGdEbworr/dhOlcBMuV0qzJ/3wSuS
DZ0/TfDdDaQbu3LxWoTsJNVOEpr2CY5E/+LVhjPfC4eYWfnEayQbXh8NASDV
uijcN/4g2YlOrqP7Bf0dRIVgSon2eOXaxLznFUaQooyCdzxmQsa/ivNNaGEr
eTdvkI/dNPwxuYVmBmlp0TDhETIbtGZiQODACPoh9z3ntpwxmT4UpDGCvAOF
Qd5dz3ek11ApdJhk5gztLTnV7qA12qYrAqbL2Nb8T8TEXncYsbzuPf4sBY4x
dECEv0FJnh/hgYOP2vo4skJGwCpPJXbb+AUqFLEkUMkI65EOd5yrJU7S2g9x
3BaN+w6CpTnxa5dFvbJ/7X15IGWpE/baC5K442kzMsjRhqpumCh7NHZrdkf6
ToSGSQI9saBJlzq7ieCV3k+FiWUXg6WE9QHlkLKMUBXijeq4VUyKIbM+aEgd
0SRuBYPr5y1HotR6xC/talpnzu7UeTMjrF4zAQvrkuJySxI1ElV01mwmek1o
09TsscWpnPFJBWaT8Er+t8NJoz0TpMFD5N64QMsqwwWdTSC6uD1RMqN9qwmy
190Qs9mZnQKb4hk1LPx9bExbq2rYIay/CWqf5ghvv/SYVFq67Z4ivDzG6xno
VY/D+dvY9rWGVT1MfKWXduf/ToOAZ3pD5zYnm2RcOQ41/AFbprXvQuZCPHxX
60LBaOsdbJhWHv/2Uz8AKogPBAmQoWTe/46OPUQdCzdASZl0RIloiZnOmLp9
f9dq83eRC4imDKFNVeGQWeB/Ahpd8VrUmnQUtwDYzIeGMOluIMYFG0ErY2W+
5pmoTrj3wdKuzRigewd/I8iDex8xSetIkzal8y9nccVPOjgIN0mRsEPpoWMh
uEb8NQw5/hZh7CwO5/zoTTc1tr0rZwVtBtcWXQOzd4+UEDdgOOcQJhkWuJWh
fkCEp/XUBW0EOAENL7AZHJBTQ4kC4iF8CzsPZN9uL6dRAKCfmEdWBoyJSl6L
xJCecsOGJgeT3PxkhG7wFetkEjuaZiUNGoHWgLlcRIqXlYUH8rhNYdczmgxx
PHXiSBSXsPMyBzVRf854lgDLwGeA9pu2ZYKz3+8DEl7vRudE6ysJEsC4DCv5
8osBM3z6L/z+mvpYQR2pZC/lUMrCmit8xK25MUuaqo3zSsT38sI9bLngR0C6
lDOuhN31/bMsE9n6dnqxnE0XowrTE57T8uA6jLazLpqaxjjqlhYuhGucbmiR
Oku+sa5SGgiQ/MPNYOejnUfbttRuPSp7Ocz8baf8nEhog3iXIfishvqp/fdJ
LiXG4SXjaq/5OWe/OgBm1oq38b97CS+dtWjf6qO8EU9F+RWyMg6PYvbfd8JI
eDNgbodYAjz/KxRjMZyIWOl6LasT/Z02/d0KyyIFVWDcG0u+09m17HirwIEY
FNlJ+8TvwkyC98drFixdoJznt1TfVKUiB49ezHD8d99exuL5yE/yIjz1oZ01
dzkOjxBlRVTIE8NgQJLl+cfKd044ImbIk7c8MT8yyOTHqjWMLPRYHW8ob5/A
mR/boq0ZwSbrFvBB4m3gwa4yydvp88hP6v37+WV61/UI8zDbWQaO3EAvpvq9
zc8LxvwATiGorPojjJTVDTlUVv4v2oObHgvfGqu8E4twYYdca+Z/l2Vn6QKY
NFTpol9+zYC4G8nN/3j/k2sKEQIITSmcM+4wCrUsE5MQ3ZZN1i92R8U/xxRc
peuo+Q5O7v16t9CIFaiH4MFjGLss7WeclCxA3uN704DbRWljKL7Y3EyUMaq7
5VUtU7ceTxPgjpbyMjp6GlQNYiaOukWFtOdeN5JFBUhd+cPs1HWa4J0j2djU
2rgZ66XMbiLKEbsF+2gXr33wxZM8CHGSuCatG460GyiPTuopQE3ZO8qcTYkX
QZdEQ7dSb+wFjPet+tMiksO/HV525GljMmT9ZyC5/Sq6oDV1l27rH/SXR98E
RiIQwU9pHcgcwD2Buewzg+UUmivNzaVXhCk0vZxG6l3dMdQbiApAwy0szoMu
HWW2+pg6jYcew25dLE9CoHE2wqhh5dMcwNK10uQIIJ/gfO1SUe/z6/pglPr2
10saCDKizhGK0eDsnjulq7pAfXXjLMT5Cg4XIjIFiTjThk6AqFB9dLFK7V4n
z5fxpi/6p2WIB8mgNN5fPA6eSNM2qDCJod963NTqdHZrtAlHBs/Ewwg+lsLE
Calwr3OOu23MC+BSoICsrF05D0+xHwGEW5r6oEvjzxmKS85uNnYAiFCDzLBR
Nx7rx6vsN0cX+j8gjnGLaM5pkkDFOLRPERNYxIEvP76SAvBz6VWFZ4SkGqMZ
5TrgVbkvmV3JWO5PGMBgsyZ5WW4vpgnX+e8bOwQqdw5rEwlBcGLR+dJYW5b2
yhhR8zMvpaPjD4HhAI2ywUwhijT7/I4vQC4ueSUdmZ1ArnlAud3ogtBADTsF
b/PSVLDTbyQ3zrd3QwY0ghBmZa2hMJzzjHl5mGI6bjFdV/yCStMmTyqQpGRS
CrF5dtjhwRm1V7YzQAjPtWCLwUmLlGJ4rP4jDE4gsLMKQgcYXNBrtHwrXZXR
5MDgYNp5mkDX6FfHaPMWa/yyc4y91pWjfIJoaYBTNML9gNYBGHviu+nUHi9s
NJTN9HF6H3T/Fvi6coeOOimcdzXqFgyAW/w3bg1U9/g4ulACDPbtJIH5YbGO
cR8zQ7VwMHFbB+SIFiGB3CnoVbQBUIkZ/8CsMYK2MsG5rS2m4rEubybYud/H
jqVR9XtnX56TIEpzk3AidPJ455NK+wZt/GblVT5l4jqb/FCqy4tPbSBWr2kh
AwkL0tMoSCP28Wi+dSO1OInLoPTRHmZhxDNAU3hgIdO2sLPpeZ1zckky/GXf
iv64b2mSRuX2S8yOH7j85HD9hCiQH2wJQQX8+rIJ1vx1G4m2zXd53hwt6G8G
8FeGR9S22Ic0CWUVxrXmCYFPtZqn437FeCLxP2LFkyXAe/8vVT0C+E9WonW8
yNPQoJbuaxrPNZj+xb0JU6Ktab0vXGHk3V3uqEjvBnXhOQQ2TuFSyp05pnTV
CTLMyYaw4g0a1TsQT5D7jADbYdnhlmyBBTjvXvapNGnmI6w+TpaNuaDkpUrc
CLsr4Xiw1rZ9Ui3j0oAXDwNHqfVWEXFhbljR51rDfg2i3fL57FXkW7fKiY6r
ekgyN5p2YEA9TM6DL9l++FfbXlBeRASe6p7NjDyPnHxFNU0t2I8nxpnGGm33
kXLNnepY1ynSCrBM6ee6L6+1Ar6JCZHdxNjgC+IvfsGZBz8+P0bYJix0b5DB
dYw1hGnOIDZgVrupSyHg0PmfhRVcQ2PzepLww0GbvpIkEMMThXsEE3dIoamJ
XzQMHEUjlR0KhSmvB6skNEMEx4y+FxbDVUfgN979hGPxfErZHXu54rnjniVl
qsgIMVoAvcpRbMqTECe0OeAMwHTLTK28UYbVlEB3iWe8G1W3BAu0AhA7/RMy
Lv3b5v688iK8wDGrNx8qb6NZtHPHCPCv1urX/agGFsaqK7jWetTCaX9nKTdF
gEEzi/g2HQgsVt6M7op6sbepyq6yBB19ZL4GAzWot4hDEwX3Bbxok3yoGphq
Dv8wkUJc6RiCPK+BwcP869QU1daD36xS0rLEEvKcFAvcx9SiMoerKMH1xv9R
Omrh6AnlwpTn2dkH6FUb5MuSk8dkRSaQ/RQ6Y0uVZR/Ww9Je3p9JuqAVZyF8
fKwilB51x2xesKVP+EjrGHh7fk1VYhECraN5szKP/L8BGu5r+ZInLHfTVjjC
rk8RJrcoFw2mfZx2CsVSblOV+Hu4cFCB19z5/w7jDa6pKGqO+DjN0hTjKdFV
1sDkTn9/3lOtQsSrW4IsBOPzunEDcAe5qQlfolJbACbVpqZ7etgAFxbMM3VI
YGDvSC6Yy0Y43/A5tSdHVK7JtJ0Qn7WGbi5KQydNV0cDlIeAGtnueh51zE3y
yu/eGa8EJvIi0drOUWxZcT1SLVDglFYihBZQgK2AgMEAaYeFka9Qpqwxllva
vJID1pkdJ+KSlFR4fOvoTzv9ROdETiBLN0ZDM+2s6yZxly1fcglUixFIBpI3
pHfYpHxoOMLrJmkhQKZtj1YR/s0Q9r6cae4nCUVY9ZGnJ9wvyIXmom2e/KGJ
Oli2u9zeBdPrQ83gQC8FRCGdMvdtNV+eMJLCj7wTzSKaqxF4rWbJtPrbyCdp
CpBSSSGgeI2DVQE0acs7BHI6sSGbI7Xr3b5+ycfNV/a4ffyL1VoFEnMEaHoO
V5ySBhm3+2k2y2W3IWE9ibqTDzzW0OhFBkBbs0IPjzT6xO37YEZGGjyKLH2A
QIN5rYgOCs9Z4b0HMGKAxWwVkVEGW0hfoDt6TGVUs98Vudw+FKFDGYdp0K/s
fhztdbM157abPdbxyd3aNtzwz/GOzL8sq421xkiDmmi7RmzGjuBDCsCK6Muu
aoavU7r6nIugqfd6la4LJtXhj9Sbj0vVAEjq/oJgUB8PbtBDyAU5M3r48Bgn
4oh4MBHDtvM/3jZLC0ijh6W5ujnB0NpHcyFcjzipdZAX411fZP6/PvUmTWz/
EewY9slI/jl7B63u9Vh2ICGWqfrR0GejlTiuh68MfbZyG7uSXdsvcpPx/BxS
I455klkBTRNawVXEzAsTUyW8TkwyxkKKbdFwmo9E40SImW8XRJT1xqn4R/z2
qagPyKV1YWpxBVh5ZEVmQPuBnmmHTOayYx3Ry3XW0ww+Bq1vvp422EDg8QLu
4bMOM/csCLvNlhFOJsLeNiIcdqJCVbqDNrd8qAaXCI6FI7KuIjXoTddmiYmO
og5PZrgaly4SzzerHbtKYEle30cauVzQ0sj/BNMOkCc4SST/F/uYHTAcv2bu
irDiCwaq3V0egJdeyxyMhZKkVJGfjW4YtMH2vcBaS85lJgpNsMHOagKCpe5X
c4MO8ghQCEXK4ZEmuxIe91bRbAVoVqFOgZQCZkK8/iPtSTYNQVlIJinsDk1q
58t+JG5+h1JZaA9ILXnOt8yMpS+8Rzlnxu7V/+eNJqbTodHU1Q1rWRGTSwCi
FbrVIF7jIN8LyvseDU4Y7b3KSO0mHOuFSowyLg3oxn8f9GvSQPB1KvicJP1w
Q0xq1EPSBw1AkHtiBgdk9ZDTEdD2BFba4jkMS7rksh2Q86gVf5fQsQFLW22e
8IO2y7cxUzkfqRO8djLNZIX84gRFmg/mqzmd7N8PCKw50r/98BRHeUMJXSm6
By6YKgtGlJ01LPQSCrKtVsfbMlghe5himAKmJJ7tKNpfGFnDb0bb+esBZJZX
ZCEOD0stXo4FeKYDNt8otVEHW8oc+eoza0MauB9vxAv2iqLoDMPLKGKwbuc+
UHF1nD6EduUbtVNh+atPS1d6QHLlRhPckaYO0cjb5KEkJx5aR2INEa8gXEnr
V8ttNhrJ/HdRT+UAtkRkkryvc5Y9a4ibSY1twg8qyVixhpoafY8hKmbBxvpB
eLLJjvNHs/MMS2I0vvWdVPZjUQ2h1MYOW8z+liVPTABBAsQSe9FTqBvdoqC+
ru0KqDietczGy5QMOp5+lRlx8ImE/Y1LVgfIww5rbaUpO8rpJ+ywpoPf2gfp
Beo9O3ZSfSnc/EdYHUtmNpTjqoAgmB/n6YKOxYVsL0HoFk0LqbhKGS+oLysg
u4v68webLWSTqlioDBosGIJevA+Z1Mg9gRddNssUYBG1j/F8UgXVVkIANQ08
HWGWV6txoyuidDVXbCGUAHfZeqf+gybGaSkihqdbmH/YPOS4Vc+1jJgAPRFZ
HujvluZ0cvUq/B+vF6lQ95AmRwIYPKPSPYeFbezf5OZ7SEn3IDpEr7/wHd5T
4iGa7EbWSB4jWwaDy1CmJfIRe5mdL7YN0nR2SSFd3zFMMScWEUIg2lQQwomr
X5CFjkzL/obo7f0cdMwrmgXiJ+dktASk1EPHmTAgu7h5i+dw2dTBcGwze7pv
2wtAgAi0RLqc7ToCY0QNerfiWTQb8OF5YNGTl5YJ2pqzf9nMCulQ62FLa88g
xBrg16SXtYI5xfFS0UgBF03T/9Jix0jJqtkpDtpneviatKlyzoiGNWuMG/hF
fDXT1j9+HISgC3EGujb+uH9O0U6WMqAj/lRX8CekysA5XZKcMw7u9dP1osDK
Mh670SgPyUzs0i5clAJNnhremm8cW6DoG+R7/PGm5lKkQxNDfRfhFBo3CJ8E
aycmurxVk3B6cdOhC4M14yIXl1C9Z0h9H2GZh64v58Upj8gLxOM0AA1wRdUr
wpmW+UV7b/fX40QTWwpqoO3P20rivTkF4JWVmkJAvH/q0HGyp6YfksoaIrVB
8GS+cp3MS3mUT4OLqHdVUAr//sKUKCw6adl+8jg1JgnY8mvsi1OU2Wp+Zwrb
FGDn/EEUd/lrM87f7EeKRsNIUMvnKakNbE58eIdi4CWZXc2KwCZU0MfRMNXE
ecT/EKyFqVbM6UmbB5oruzqrfxQSreHT80OhQKS88zFeGeMkWKKPyR9Gzhpb
KWSX+JLz4mLs58rkgPfxCJYUHm2YpXMuiR/Dvntw8FBWiXNJwxe0hmFAvo2P
PImA/+/6YjFSmcf+hi2KQMONYJ9NdXpgpsyP8hSTJUT5PwYUFtWgYr7QB+V0
qA4y1rndN3mQ8GkUq8mj/9kCs/5tYh94AuS+E3cdsKRU/r9oRUvoZSTEFoVp
P0fN2G6RacqMkNGHTu4BDt/3bSyCIRQKzsU1tBFXXSZfZhdz8p7Up0i4Y88N
LW3cHb1vPYbArbnKy3nkGHw/HLY40lpjOP7q03QRQP5PokaJllx+BzneQ8T7
MOZikkUqQTKLXuWle6Pd2QshVE1xi/YcsrTU0mbte5pauE/GQJFRAjlgYga1
X52tBz1eu+kVQvzupVEEwQ0Obilv1+bLf4NxP4pE3vHq7J3sMp0ZQ1Mlkfmb
iWG/aS/AGtWIaS+6PmGrje9hETIjQA2HDOMcDdULPNIUCUfLL+hMdgXrdf8i
Atc3hDCMGmGf8vzgV0qi/Z3OKJMmQLC+YyGFFSuxXaVxBztfkItSeCOi3BhF
nDCa1aDdYn5D5Nj/1dD5xxr+MYYkgTjKdcVfpdddk0F+OSinzafvB11jmT0M
GU4pKIefv/M+FGOc0KP5QpCDyRPXy7NdDcR0n3rHH2DA4nmuL/OZ2KCmVc2d
r57CS/jNM9Js5dl3fJJtHT1sDXGU+P7IsfiFlkIk4sXz83vnASxkmrbb0Zrc
40e18+M062ODVXT947lfPlw+NvERRLDhdccrm7dJz11sETjbvKjTSlk3Jhmg
v7T0XrBmovRgUN7LxbQzSePTAIm0Qc3H717RtjoQeh25PzT78YwPLJaKyxV3
15U6bcnOYyBd9Jn4Pv1wLWov5jNLSGxn0fzT2Q7CYLQc/1EmwgBofs9Xzees
1LxCZZvthWSXPeY46DKEBVRx+ljXCIdR5idSf1m8WkGi95AMW69tuxX+QlWb
8tskFoj7+5mQ04mxbYcK+XGwPVIqWsroD1iwziyfmg8zULrbNS+cMYjOGolA
xbDNEJnx8xVrtrmzu4bNMcC3NNGoy5hJVDi+bR9Hrwuzk6UF12zqS4Jdy7A9
il6mKbOrsDyGCn6K3SyfnJtTH+il6RD5mviJllnoIW/CmR4h1U+wi7PJHI26
3UCXn4SorSzyt69VPf+4baMa750ONk2cUj8XuMaLvmtlrOMLGjoIVn7EPKOy
DL1cZ5i2Az8M0jivQRyC57G3ZiQpIVKYkwn7ooQa7FFL0BCGwjp9UnwmzAcQ
kqzi93IszotpPmOduDPGnp34jwLTcigjRnPChTbF8miG7usOU/CV9YdjamZe
0sOpveCK8hdAHpTYgvmEm7aDd5ysgHwtdOtCCG4WbuT7sTVNzhMipX9mP0K5
txzd2yDeAQXNlYE7h2aLPI/8AwTCOkxRnTck0rc7oKQXFye8GGZBJmWpvw/r
FYF9JElnnyh6WhcAbg+f6U5ffzz3lgg6xHSwrB/AW7xfLpkSn+KTuZk4YSlh
0wHYO873dkIFohyAPU1BOtu53QJT2m2Rdf4NhKFEoTk4bN9qq70QR2PH0yk3
mXNoLNKLtWolSZfCsBnaS0YoAql97IKsPq/UrxUeSXWp2v/BTbpJjv7DP/0l
18zulgb0SwuOzeTnwuPQ3EeW1+45glyVPN8if7La9JSEhZ+veBiXoQ79Pzxi
N3wbnrQi8ELgPoa/9MILEU6wpwFLkGVJsSUp1b9E/ocJ/MFVK7GdHT3eapOi
IefyIxXrwt5O6Rubt8LgTttBI8jcjzrb3kgNNQ9+T9aQTHVsn+c8Dcs1rQ0S
JLfQhFyQzTiORpzlKeJexmKKUjyNKutglxBjevRSJzbb3Et7NsMDPlE/kgh9
ViIo3YHcHKSaiEEjOzrpvegp+NsWSZ93+CjUvGWACeYuMxeT4CqyqAu0AyDb
OmBkFgLKO5L5+bCPNEoL+esJCzpFxlYrUFWXDrrTA5fV4JSMyq3LlBrHMNDw
n8ttl0PQxQxy75QjtmihmVCrBjS7dqdS3OjMMXdvQQUTL5Uh8YKe6fzW28TE
FjpqACWQs0xBR7BGj6S5cRlh4hnoVBTb10HXN1yrkQIob4f3v0jv9j91gcpz
axItqLLj4NDyWDeHVJEpxPtjaBRkn2oodkotVzjRsHcJO/MgyXqItLHcfwua
XkGmpHBrj8ZNP6h8R2I89luouizU8z1jYhVGqJoKUpllx5MrgpPHdVAHkNxK
jUE5e0Z1Jqlsz48FwELBeNkRuYrDpU6hF8Q70mvkM+/v/w+u+LDn0GYPWhcI
M4Dd0dPaI0Lm/6X7OenjDn6RFRV9oKSRxJfFH0oF5h1+GojqYs2iL/PwVN9j
xCWiO4as5NVltbP7VM7hhZ/VlNelGdZKVb+l/PMTs9sIdZoGnTECFRkcAi/C
98RaG579KZYnlUOmjG5P+UAzUD/aMeBMbrGS8kQJWtMxK0sh+NgGuMsDFBjP
bjVS3/uJD0742SbgRKvvAhiPHp4Mnh4mTMqVZyKvQjs52xHvYgUUuGIKl3vu
Wr0uDEci4AfUypIFhXKWoAe/DD+E6RDaZi+OL01jPqqxoAvpuh6ieb1d2H/o
OuqcbfqmXh9g2BRlfvfOYfNay422WNd12LB7vjUzupIokF5rRm33/vtZsc9h
LHr8K2xiDER8yeDBtQ7Kx2hqoOTNgU9V1PNl5YkCQUj6B4bF/XOthHH0ougk
VjY6oHxU7Du2vl6MfphrZTWuejLdU2g70G+WPtQsUxlU1c4Sjw61M64bbVq1
a3nIRpr57vEmuEb0M8RrLPywTvbZpRYuecLpsY6iUv1BF3iHktXbyzG1w64E
5J+YcEZsfQXjMuP1GbRF8fmZyfSdxDJgik1Vcprsi5lqGdRnxL1FJGaKGv9e
+APxxaLJK/AsGwXDWoyJTp5GLnJzh3YssxcqYGGl/f/ovtvHfGb1iTcHqVi1
97lW13LIutacED7CXwkcHBJUpfmpAm2vl+uV9uVx/c5dbs/GvtaiQvYYPoQK
4Hex6DxNz779bqHMvNiuKIjVhe0GrPsCLTH9cSGnxd8WYfvqwj0x3vLk7JV9
E93P6RkR8/A/BF7wdiULDYW41FA4D8RoI5Q3Px2P+UQYvBBtLEKsw6bdVONc
XFBfiQ21c99Z3gMHpRTsX9qi01DTpvLXhKXyjc7oDkfuBrEvI78bG6AoeTcK
kUeXvTxj3WAM1oZLJAQzxyCI4DZyuukIc7TyH3J7zuYEz3tY32+RCtYsKb4q
d+cLmrrSGcdrqG/88SWge1asFs48c7AzoHIFx+L3lD64i3SqgmXCGMcX/sA5
f/bX8Cp3NQzl0XUsteZ+wjRxXubOMGVKVMHMt7uf7Oy7NWNQNAzLk+7uNX3a
msM/Xmr2o1w4qvlcAmM4hOKaYj5Q22ugiyqI7L3AKUdpS2zSP1ahCXAwwfVp
rVgtgu0dwi2j2IaMQWi9mjn9tPbAr8opT5hEIDAVTXdsno2mkddAcmDfsENR
7gkJWI6dh1xOVwkxIDqt5Rv3873zSZmek+XTLL9E0AAqIRV1NiLrIpCJxk0V
esB0/0Zt+HKhcM3PbYe0VkNQuEJ450+1YjBSU4bki1qOhPcoNvgKCwVGVIiO
BXX24SYqJ4VreQKTX6XKF4DO7L12k4QywJLRLEddv+wyDD07XFn/LgXOzoe0
l1RDnKU3u6BXjdVWSBPAy1LughZEA93mMZqbrq+BS7hx2ZoDI8ukj77LqQYN
SX0hObBZ9Q0zgYZf2rRyd2rhtDPsQbKyriZ5+gjEdfT4pUvpYGxdtv4LZ6PT
qgPBicmeEdVI0rzp96OWZfYuWxdRgtoEqaLG+F92frDBHCfJp52/FGa+GGgI
TP07tkqiSuOdgzgJ3nGDIhywRKwyG9PYbMeQYliC0yLglb8DdP7+1uTlxZai
FKB17tbGzEX7LLAZLg86GhMDFdXqSRwmckdXbuckhETIgYOINNG1ZfsP4woY
lzxuTo2lDkSVMlSIh8pPPmq3L3FDPnstgRurh6pLoab3aW/Opx81tVcYM25X
P0tGr/fKxDJkrSiHHe+94i5KhgVA43jn/yP9Twy6kBR57jnBV7OsHHVJwYo2
E6Q32qwTb4G/2bGxCAgDutCSzn0lmtIfSyAlEoltvKerT3pCKO2ZAiLUA8N5
BfLNRgMbj5RtS+f7rrB3OZ6d8p1qKw0OqEYBpAggzwlClEN8SxoHQtzEvWDC
j/OV/01ifK7KYg0eFYfUyK8tMCpyFg5dx78GL6EKWBBU9BoWQaw9qP9SLbNN
9Q6jguwv3E9by/j4MN5Kh0YV2ZXN+w3vuw23ZBme9rikx8qajcOdABWMzGX4
IKvKwmbgP/4oKdbgJ50BpsRmjVTt9pUg+xMxkkJzwIVZaV/iS9Qx4ji09qGI
jywRVvq4v+kQpUNQLBywPoakjIK0q3qr7DXF0CmIr1afPBFRlAEt+HA8Hxnn
x1l5Bp5uhE2u0stQh+NUqvNnQuOuJOJH3QxJ3s9BgnnNHLMZSZQ6tZH8rytI
6U/rE0jhFReVCT6ma1hpyK1XAXupKmmjU2gFsycbcgr4D4UVR5JHDIXtJXHm
SBq/ZLy3QaPNiUnNQS5u8nA2NBk35RSz1lP9XFxi6jq5nKZkzruGl49+hWNW
GRY9zrlGjAc/VmsT65Bgut7rGyjRS151bkPrbiYA7JJV9iJhuiVVTREHj/ib
REp4+AgFLilgMugnuzh3vPUXoyFF0FVNSKpfdmBmhPvs/Y0TDrieIycUChUe
uXFlgRHV5V15F9KiAENznb4a5DoPsSsDNHPThWyLEIRLfLjp1heu5XL7HvMC
QW9+xIDbl0TonSCKpSR2lSCUr1rKwqFaPPRlZxUAinm7fiz/BocNsBEdxgtv
ZIC/jmUCrWNdXJ4xpdf11j6F9XgXYHEc+OtgTmZ5fcX9JHA7iJhe2haov2Hz
ujDqx1w7RS7zW7vJAFv/UG1NPkun9TZpFy/WfAG7av5xxGK91BKsMtJOLG8D
GUUo6YNTsNKzprP+h9c9aj3I+MqICP5LdrJ9i9jhcQCk9asU9he5rnP8xTew
l0av3tPeoInER3gFbBVSkOpIAoRSHTcDpze4O1wn0vqm6rzahdlyiAz3viUs
+aNHQGrWWOPmq+mZPiuvZx9I5kXpxlBxqTDY+FmLlTglwE43liKY7ybYUnOS
Otb00b7dgzLxLQ2Rt5EN++6ochDA29KDOJoP06OjoyBsdsHK/Z3ZqwRsAw1c
m5AyGCdX1LLfK5hNO35XoBAU2aD5yhTuhIdaI2OyUUYpJiNBnwoUxT+wKqCj
Qu/MkgXqsn6tx6YguByvtlw63ky0FV+YjeZuLu80RFjSrM22Qn4nY4jaW+H5
oMEmdvkAwHKeyPSMCranb/5UF+dqhYMFiHyN1mjM8rq5j6NneiwUUXKhs3Wg
0h72qxwRda4GfCsFRkPSFyy2yHvUENLB+wgQjhuHhIbc2v9jkQjLpBHBMMKL
eqNVb1JhkZS1oYr1HDlhwyGQW9cSmcgyKt68ODGvPrmFnrn9lT742jQlhjsI
AurdQ6/XWrI5tM2KrslN0KDg7OgjmB1midCdod0aUGLxnqxkM5cjui5QxO0N
54jjm0ejqAnnJbPTO9V9Y8rhJVIwN1XyhQpAONFzEHfS4PvO1nWdMuTfBwW+
03YhZAyYePWafrddVpF4fPP7ADmFQ93CQ9IbMqp1k/uMwU013jtsrY1lV0hf
EUZr+Vd+9/cUV+f7gMO+vceOnHc4NitQpvqBca7Y0hEEbveMR+vEdZPfM2br
EWkZirkLnNiqMZKyfmL9NRbVncbsKEuvGASRzqc4qay6wpd7HNFkbsYA8Q0q
/n0mc8vtYzFn5U4HzjGi5LxPJIESFyIL4PVXYL4SoF88mfpWN/zHxTjr33cm
qPGPyDYfg5I6wOb+IAA0lPLikwuDdE1Do9ZPzKEFCqwDT1Xe4bqUeD8GVTqN
VsNNGyN76mCYEoGBXOC+J78866SisdKAB50CTBxnYs6iCw6zoyjdmvuC1foV
tBQjm1NMpLHUYjBGtRpYKvqmyQO3Qu/zl9H3IpG6TQOgpa/KfJxcw2E0UPSf
M+ybP9IJJbWU+4UG+SvpoN84ETsMhDWi9V73rOAx3gTxRJRiYBSMkGqwpFj5
8hYsExQsUhnBdgufRkSEFqKpbTYF7gGBKISO5aEeZYjoB7asfT6PYcBoA/0u
uPdTs0lbq2Tl7Hxt5fILNLuDicjYCzs7SSfB+Ycy6CLFdEfMBY3yCPrf78il
o+3nI5k/BmgL+WpvrCh6D73h0ekLVwKmkFAsvk/oIOF7Y/RX+5yG8iM7gKUK
xVeBtxXwkdwWH/R62X4F9/ucWIn5kfHj9j46SDSBLpjhE3aKmebAYRy/5c8H
hJBIG9HOfHhJeFyjajxIUByCWxq5t7PW4Pt7XSX2kRsv8IHV3fhZvz6scDr3
zLEWiKXXJbGLpn8tIUf7Y1BpAfzt+pwAuUGm5DLfCdf9JGZZ6vBy0XflHSmN
w2+hUeqxoN0QZwmT2zNjB8PXGOz8+E0W+OuuK8p0I6qamfbsuDi8iwfmLjfE
PccTszhVvX7pyL0ydQsi2sRVhFfL4TtQv6k8IA6KIq+glvHAbNZ3VvMQr0v6
T0LFP3Gbv6QeJRp54EMfkjBmbd7+T4Qpr8n4Wt3e2f1eYHorREy0RaTfwSzH
qnTht8dQOHDkzyR008/NlmegQaJHSUy2eX+6w7sezZFvHW/ppFJ8ksMZKker
6n7xJixThRP2DYNX27kPzFPHTnjWzmGSDZW6A2Fm4XT1OJ2HHw8XG5KDAMB4
vfEXVuQdFp3l73EAKvgPpp5RGIYDw+wKRP4nrUI/bmfQcyddIuK2jkV1MXRi
rH0SvFAZQknOOkIVtidR8wUomCmfNFne5CgR6nkOirvI8mKWsLmslmNVXbld
74aPjFVi9DzcBj/0rLFIL2reW4bmHZ3I/ujqefCJUP1hzK5I3zI1828SrqJU
t4KTvzMKcg/7VSPQ71oUvb5K0iBaxJINtMyxHqbviOtibq5Vcrk4MNi1tD2G
NhN4V3r6gCyPIVpZqGHk2BOn7Lg/V4IFex4WUVx1nqpe4UrcGZEaEQ6jIq7J
lYMm4+6u95IsR71ZIyOZAVwNf8WT4nDwdsh0XY4p8DbgAF9RuD6dUGFX2ErI
YkyFsrWqZTVUjiaKBpbiJAdD8LhdEGOSirCAi8Gf2bHlyLBCvOIQu08cEFB3
UFf2a9EdjPaIWDWbiuv661nUvdeyjl1NpZpeHMOuhvuXxhG2z9qXX3+kv7WA
uifnVPfnqkw9GUVBUbrn2VbU2oCkcY2ouHPBwDXkBMnew9sYAFQ2OacFyNsC
5NZ3t4ZchI/HXOSosKf49DL/NC3l0ky5FYOcWurM1DtTb5UAgxu13uCka0p3
up7Y7neGGjdQpyLosvcgs4udFOXRoArIVGyif7ylZ9nbf1PkF3TD0xL6wmoP
0LWogFITMil0TCxKrCvzVKrD/+oFysXgq0+R14i/Un1r3CsAnS3Fzjrd4edf
fwiE41ViNO+bqxN2F5d2F3qXUupLBK3Bl54dxfYjc9G5alv5GOqBPYgI7oVV
bgY+BSQJS5uEeFaRpq7C47F8YsL+z07xoJjcB/k2DL9PRG2v4xYltnC9IMI2
XLkl1HSBsRvp4ejfw5LUKwG1yIcgWHpBc6v4eAVy/Zir9EpMTzkfsNNGkT2Y
mPQMSsEkBiEcDDAThZLtVekmYtDwwUV+W/P4rI07sJUpzYNG8aidUJQzNkYv
8KZF9WXgf2vWQXA6Sg+VwWbSEIKVUUBFgNwaUnY9vivP0ry82DN7S7Xi/Rc2
csKLvZh+kmHeFGHJI3yiACcGBFuVt8mDUr8ni5XIgB5IgnnWHf7GdErAOf1/
XA3usSrapzLQ7tSxrdmVEZADf6t/2Y49UEj+W19B58pOkE/KRx4kt0xVZrkC
TuLuCYcLEpLLx2nWDSSVHHVK7a1uTYzrxTVh71VwaFWSvkt/1XLSbwIE3c95
+LgCWNXvlEr4xS2kD0246psYr+secWph+25lMNAMCQTr+FT8ljveggwVK2Vf
40kS6dGy6jiESB9f1BRs0n7pnr1fTWnR9m9RqlngmYs3YMUN+WXNnqsbpdp5
ZvnHzt5F0F+RAy3+JN+WnlQ5NzahmwaW2hTgmrJyP/C1GfNd6LF0A0NefWJR
flep6vF77oUh3BpNT8Tx/tflKiSE249TgNbCm7yARpT8RnholsFf4ut44VXw
/fba4GtzSpkyu/FWif61uQes06gJ76KMj1KmWYU7kcFdroLO+b6rpUkr/cHH
8gV5Fl9N2uW97AyakNJ16iUYMkRM/r0jRPTurBZbVL+v9vbVooPL3AyKyK/h
Utg9idVUaeIiF4rORrQbCLo83ll02L+CAbyxguqYJHJSZ2E5JFdAHLbUpWiQ
XU5d7pajcLlCxpXRhOqWZ7dyx2yx+RrYO17xmNnzfrq8ztesb6upnKYbMCn6
0gpgqeIMw8Snja8RjZh9hDu6F0AmQMIvMuQ0RRERXa7w8dLSTJJGharqSmbF
T3vajreXAvL1QxdZar+V52Yto1NX9NH5kqKyEHC6sW/1hMtwSYhtLfvUkurW
CpuveD7w+9IpGiwYydMrDoItLaWa2mz34DlyBE97WTSxk4mRAs/MwWaz6eK/
KKbQ5gWjNLHNqtqNrtCH6km/RjM+o2W/Tgk2BtmesoFa3uO/To26UikCXOuR
9VbCxxxqXyfQulSvbn6ipx8y59CmQV/IHFE6YXC9U1gs4acLX91/m2MjkFgj
VF324HACDiSxNlF9iQnKz5l6ser5Gm+smCxbJ52yJa0vNij0gpccZXmb4LOl
jaZXrmd5CjC3dF++JPSiMWFNawoi5sDh9YFCQQi9ssWps5+cqEUdmkOdhnZ4
L2o1RIz+aBv94MU52/DlM7jj3XxamPXSQL2RJBi/UzE9Z5cyDT3GezE1Whtw
YGLjTkHIWAo1936FLgBLTHnIs0Ex8enwDiQSxPGwN70ZXvJ5HdwdSJqTfr1K
vI6NjZaYB79NWVLkifWMbmewyqQErX85x+JO5XVYvuSmf9OeqxMl4sc0TYzy
uAQWRxq1nUZsWc0crTNjkJytuby5TfKhfPiy41gcPHWE5ZmxozvHPGOxBHDQ
005KbWRAlOtJ8MXGnV6RPRFPL+Vu83eftjaRbvmYVjZyJiW1OMqufWawRQ8t
3eGO40ys89u2ZY+cB5J/oHK2kgi/qIzcmalm1MrG796sXLwqJQg+DCQgzcI+
rKzbN8ynX2LgNUNuCCA+VO2y8rT2bivPFuTmdScC4A8+ABWx50pJKMP+WY+j
7TxEeueq2dCV9XBVxFmetWXtMLyMgAHwgqOcej3xrD0UuF1SJS0HWKsL7OsQ
ymrYOmVOhj+pDhaAzcP8Otr2t3qxjqOOHnx0sONH6D93+dyxeEvNFh7/iKBQ
FXvKnnLRf5ACPFnz7+L2TATtpKdKh5Ds5nw5KNFdSGJRFGUH+0NeVD1x8C16
Xl+F5CTgv4JJ3fYUlQTgU+6l9DZnhqiflKzyyzfi2IKzjNZ8kRL9l/n1GpBY
ozkn5+vUHHbKOHEPz1QfPQoRDkMB6kO37mYxns2zieSrESLcp+AKgVWYfYy7
0219ba9PJAXDNv40oqGCQxxLs6eBgmmgklU5fIEeZftHG+wRx/CUMWfdlmDM
oAhm8g/SQSp9MVkhWZMNol5gLI9/1dEc2o3Q3D+SW+ZGPg0ziejtgFzrnMPd
8W8GwVuWPunBjwD5SF/bj9kegV6e3YAZtfRGbqGbCqjgmPZm9ufGhhbBVFXF
Oqv06ObCMVrmNjDg3B0Lo7n+x8PEB6dIMpVLpJH8Fihs6ZHuPavN96vQXvVF
LrLs1V1JFjzapa7SqikekYrO6xzmtXX9w8k5BAk+kev5hoYfyvSrA8U2mJpS
K+j66LS3NY9qmutllql448B9B/wvHFI/XWEffZw5V4UudYScIcpdEibuZz1g
R0TLHoW3Pn+8iIh389VC6+Z7/cPVHJQRAdOMXALJeoCC9A6W14mWMn3+1tZ1
2jVkUPQdbRfXGIha7WO/FT++Z0E11NxuUYOwP4o1hrqmO8N/f09gD7MaRMDN
640U9RYTk+r3DkKa4qsRQZRX74h5GVZUDlUWPDcOxtqqh/fBEefwUQkuJ9cF
53EW8//v0iMyGEiKJfl8QNQ7T54BjTKFX3UFfXNleC0RznSxoKrC1wPFKgVG
DwUD/hdUQlHa3Hq41aoYfDo0DFiReX+UXFDF7vStjDQ6M6YI4IaikSBL3UYc
u9/SfoQpBOqRllGuaYLB8cziFO7PGTfDxMBn1OAv2H1WUeF/SdESDnuCLqiu
fWkdKwLyvAGE4c5thu0Yf8RGwhYtFGZFGoYtHSstK/WqaLQ/rXB9mkWtdeGC
PYZPB9FLYkvdh7KWXIQcXNeRr2Zwh3CcAJM41OL5jB4eiaHZPCWNOkFBoD2y
qDCT3k7Zl2Sr3M1FOeDGCvEOG1rUMOF9TpYgvSJ+lXi717kMC6GBy+OEnop3
3IttLyWyayQiX+JUx+dqsbyX4teAd1o9GB4gbWOP4Bc+gwRgigba+Yyk99I0
+lhrNCJo9SsB2Sxe+O6Lx97Fw6YNQG6fzRv1vdz0H8cKimkzUry3VZ1+lNbA
B1+3FNyC20eDuZ23he6jN+Ww7llLFSzH0cYHxPSn9LpD+Xv+l7OzZ0N6AsC0
EOrrkPrUcyml2Ps2htyzqKVxqwYz/zcSp4k8hwttI/Vmmhd7VJRUrKEkBule
OST31vpqQkAMauzMMvnoPIph/PRXBBr4FVrP5WKxmTqp107X2CzUZ2G/SR96
y1+AB8uD8xVzskc4czR4uLWCP7apIF2e+M2MZS4gDZpCIqFkLrzvzSvv0Tgc
s2u3KfEe94Tmu7sO7F/2UuDrea/vkl9P5jCB425s+APOySXUzH+NefnYeRwH
s3Nj0nSGDI1UveA8qYcTyCAOJGk8jkhpbkLG1r5RmWvkHjW3wv82brwyHOYY
ej+v4gVmgZ3+Zw2ctSNPjyyacpJ9ewLGwMeE5kaRgEDFpiA55o3DLfxF+IJb
Mhb+dVdYWSprGh7pVeOmpbPz29Zx98lv4uYYdSagvj6HHWwODqGbGrvyNoFw
ZVD2FeV5qADXuO1JXr2rd7SOCNUsR6lOpru7dHpJsPjstJFYjqhW3H6WGGR1
xVqlVuJ/yYLyQuvB/76GYjYP3Sx6y24AQ/ERVl9Lx5kugslttSKh3F6lY0qY
L6RVzr3If+1a1xGZxap3mNbZ6cXsahcQVtbM1rpWNDl6Znk+GeJeeKNqTWtz
GKu2PlIE6jWZFESvoAG3Bx2ghCoOniToUCykhOQx6n8r/+WZmCdx8dtYEk+P
upHtmElCEp6dTdrOZQkgbSdrkIuwb5hWtYOLejsibpfD49kZ7es41rcTd3Sq
Dzcqf60466+QmmxLEFEWDRr/1sZ+VtpO1C1XP0eDIdUUvOBGeYwdRi5NiC+s
ZJTwQn2xcYkdVJW4xHvpWSeB92IsaMhpG2A05/a8k6oqpCzrCFvKPIl22MuI
NQBZxQvY9nfcQwtLSa/OQvtK6X96jYtXZBlc18QExz55mtjKgv1h1243Fr1u
xEGus8f7lxPlmNf3WnYkfZQlKehQjhNDjGBhSWgs3DY23FJ671zyWWDhQtMX
l2iN6dFV6nTsaXQmFsiB89Ixmi4sLLGIYJWFKTgzBKOLSfstDryY5vUP6VHM
eos1cYhsa4e2nF0c3bhl9uJMyU/lvlJ0EbisO19zr7DZ6Oatc0HkHGXVNjI4
Jgmp7OFyb1YGtLVQBnRJ53rmu7Q7T9r3W4Ce7cu6SqyNyPJCWW8eAqIxNWGA
4H8rijMQeaHDbwGrG0mZgC4DMnh7gE86xRhWikRRKUAx9IQ0MVAA22qr2cUJ
clH359XqIU8HtfNfFSrdl3fMWyRrjF3FwhJJOu5FfuugJrOyikHxM78ky5Bj
Ee5R82x+WeJ1dzxIApObfql/6R82gG3o52b+SrOUkKdrr6JfmTaQ9FfDyVu9
BdR+O4MgQd3QbuEUpj0TLYJ5kUGqpwoTooc5MackYsGPsRhKbm2d+csfMOvm
3/XhsE35bjR5btRwUtLNiWReMXiVT1YVy+2YbA/B/yNxPYDb0yDnW59owo85
h/2E7iU+KGcwA3DnuX6crL6fLpbGxLcBN+r9NxxsMMWISjd3Rbzf5MjaPXoV
1gBqjIV1AwVjX0SvazhcJY1rPO/Z2MdAzIUR1qOGNf5Aqb3AO5hItpE+/2D3
7mq7OLiPvdAF6eJKEuiK3N6sJe+bkk78Oi32wovmUztTn4KSkVLAUBiNIHhR
HCW1msIdTkY8y4C7Rd51SZSzPQwt+K1/CQ60YE5yTODdQmhP5q2HqGVJE4Ab
8lW54jy43zUMR9i5bPEpJm0jKmgtkAdCqaYocyy+0N9srLd0C+Bhlym6qvrv
p3ec2lwYzDxnYqY9Vo8HhMncx+VKBxsRAIj8Pk/ssqGb/BZwAVNzN5cN1lG7
BBmrBeKvtocW6pIP5ZUNqbEFP7WwazgS1Vq8voKPnJSesTns+/UWi+t4TUTV
lbuQ7hiSRpUNIYLQHdcuCcPiPjsyiJuvl9ltgbs+iApN45i4Gd4Y2G5adz5P
BdGvE/nx0Lc4ABfyWPJ8U/Zki00fD8newiu8Q2NZz46J8S5TB/cKWJmR4WIB
YEefXET0STULQJOqeIqgequcaOcX7jRKOPcLSlnHzvr41iRzTvht8rTISGUi
Uo6LYBEzeaIQfMjLINZ3A1qZ10AhtDpRVEBMe6TL2Ulu9w8qk9KtBuZHRgqX
J41JLF4I5SpE7i51sBAfZVFgk24f01z1j5YVce2OAc0hb+OCDHVGoJ4rfm6T
TJAZIJX6XoxiqqW1/lvucumCofFNVXTaPEyhbBohUmEMogfWDYDqhkwNRXUu
S6VT1bTSRO5iqqklQBbVeUlYHHuCvO1n1eeLuGDA5otZGXnZcOA7bE5teqVE
8Od7CdNxVQGrJkGijUJjn7VfSXk2xJ/hGoMFltUxYCB0QN7txi+fv1LeiLld
i9J9TQXbp4Y3SSRZ9GHtoemecRu+MgLFqHztBxC38bjttp+Pu+rI9hgixBSC
BVh5XX1Y7eq2NgbtYlS7Jos1BaJ8xrpBr9gRYAWzdA2+vfWWmdaUcU3PA7/A
oCSZYFyc7uU5BHpgUJANW+7a3/xHW9+VuHX4Mmdu87iFsDyzX10Gjy6B5LZt
cRIgkOBEk+B7OiPJZZ8f7X+FFfEL7S8+DTiuLeyCgSX2LKHGD5UO9y2Xq1kc
rzPNgdKHkqJ78wzcNfJjzE2TH3KkkQmg2f8JWIOKF7VRqqAxB2esTOptJqoK
LZit4gvvhrrizhyviZvfLrJ4kLJttV+cS1++QMR4xny6PQAG9yi69scHk0jx
4IFille78FH3W4mbx+l41SBbSaTJc7IWpcj2wYMIIdEMwnlv1rL3bwB4C4nS
j0T5LBOxmEX+GdkoxkV4OoCX1/EIrFj9veghkxM17WP+Pu7XxamtaZUBFKGk
W5q9UkQUecN+/l90+y/tYLgLSr37UbLa/r2dgf4Fx/UdSe0eZcysZzWU8sIY
3Mwdvq9wJ//XDDQ8acsXWdVQnti/3ogOElqJeHa45j2+1QvTI3BnC98L6Chw
/2bRAwLaV/AS52RLotisQJfyNsx5GUeHgdZAN4Hn8eh5Q+qNy2Nq/O9neP2R
qtZndYue2WCTA0opKc63P9oP5UyQpWWYFuSzLC/cF7QiyxBSumJUgM3m/d/c
UQ8zGsxqJV0SEx6uAl3fleISTrnhmi7N/8sJxbAOxI/SJZ/Q8w7ftEKJcvAl
nswtjhHY1SwIzkGA7uwXAwC+U/a5OrAAX6q2jSsG/uKRJyyhITI5hMXhrJhn
i6QGn+gpz1U3j775ty89H5pIR04ezKX2T2mbcnvm4zjkq5mSqcrKrhFpvd3p
/7MTYOwKqqFS4RIqcjD+h3JU1cfzY6/RD4+xYOpMZVhnJJVx8LlN5FqXBVYx
qvzE1FDitz1D10RuBGYF3SOjbQFqhGyxvgnDFywfhJ0pIR4iOnGNd66GZ2Qn
XRFUBXnUBCVbSZ60/VHAqgwuH+OTPRXFHaBUNUXfse8lVVUMd/LX2qG7Hvkn
bLRTaDT9yNIAvD2z2f4qUrQdohbgfXPY6G9RjgUS7pjmB+WhZLLI3/s2kCil
R5hcu4BXgATYfpX1i8gv+F+OVoJO2ZosrF2iBcbMyI6ocrzVXviaU7Q+d+5j
vzzrPAMVuvxTRTL0WuZ+VvxZex96V5tESZlKHAU7HE1eb77eE3305MvS3yY5
gSJ3KAad83zzoaHufp6fgBydrd9fefTMbaqnEURRVutezr/3QcMSG/tsAXwa
YRAfVi8XuK3a3rW3yGeEjPEKKcwd3Uuoq5T6LBPOHSx1kqqcdcqoSNr1mCDy
czK7W8bVl01H9MRzfRuMRJ001xhGxej3MJmzrfd0q+jykv9ZXfMgDqmK9zhk
LVQl0fbWwxcqPfbaEAyYfHe2E6KffyogqFaM4iTGd5t1v+4Tf9KrYXqteV9z
Rxga1kEyGxTPBDCihtGgbqoGKd4bztDbTLOU0PQmM/3aSyTYSJ8vaEQcrg32
rjorKksv77bruqXt3RKeuZA8GrQu8DaYWEgpAa7RijLSD+MkSMmkrjTXOu9X
lGEcBae2R/gOE8vrf6pP6sfvfELccWvYhqfZaNT3T+kQS6IuvMq8k1wGJEcj
8k27KJbZ7fQz7XemRNZ9zFWwb6+By6PBHjr0aW3VUdDQnIgJPvx4/UVmjR61
wHoqZcA5SKGrTCwzqMJm2HEIH+sI04/S/v5QczrdWl14XGtIYJlGqS0yzwTh
Ju2YbgW6j3pg71OX/0elBUAZuCnQRez5ZqcimVD+8iFkGHxYNStRpWBWwlTi
MwXhNt28C9dfjNTPuClm9uXqv+Oi5c6BntwIOQGFRCA7157xOnILC4vAaoWW
7ED+din79wCO+0mHv4w0LKNidj/6w3iuSyeyP9MheQDe5s7BCtW1b8utqZxa
FFvmll8w3j9J2mhUuSRT0qR+mPFZ8tyeb6CzkQW35zM7LdymS/Yqw+EEcNz/
lD7d37WZuc78bxYlg6SAfqy66/Q68ihgxZ7GsUngRuQ4qrH2u5pCv5x3o75d
nWLElXCdF7Atw2N2MC7cm+5UNcoRp/M+WVm8c3RhnKLWiUVKda3MWwHzPgG5
zPTR39VfaBRjdb0gLUPEooLiedQ2eao+CUDWQFQ/l4VfBjUu/UfA7MQ7lkbK
Lg3LzH3vylvfWy0xwitBHqjOBm9WnNyAdV9TiKbewZiARKbLzy9a9n+ka8th
WURhScid0VYLIS0cO6jUoznOLnCoDcIKsOxc7RuDtzKmoYimXXvqYzzKL9k6
ui7ZOkW6YYf/+HIHn3Zo2yj5MPUTe4HP5lxViHlkmqca2/+PerUUhP33MVpV
Ts7Iw76d5RGIurBan8OanJJefNFS5KizooQvvb3cJ4fXkBOa8oefFXQgo4UD
lqJHDYi89ot5U8NSWyC42esBVueIea4vUjuZQwIIl36Y/UZeNlyaDthljTcO
qOjQoObkkMkv6MyOkczfJgUx/MDB5CpvvgUzpVuL2Af3hCUVoK8UJ6Ko0dzR
rkzAcIr4fobmMnXDvUBNR3hDs5ewsqlVoo17DHVp1j/Tuu4gpocBoL/Es3go
WGjC2Bl4SWwGAEE4Wb3FL27G9PXHb1Qh2YeeJvVQ058ciKEvLZXtQgwveiuj
s74xZx1Pmi+/P4fgwKJKdfY9Ea7YqSEhFgThhpRQj1Zc6J0wa7oiGVBaYNRR
5lpX+cT5a5sqhAQw5KN7yGKQLuzqflorXr380fv8uMPd5vCODNsr8aV8js7R
9nISR9zE9RdXMczvd4fFhD5+HAn1ygpYv1rWWbNngbXZ9fChSatNxLUBuhQl
Raoe7hlnijJo/XrUKQzc2arXZXD41H+f7QMMWfeCTKvlBvJnL90DZFW3N4YC
AnQa1Y7cxAElPp1HzcekMT8tuQuSwM0ejmic3cLzQ8g+lUKj+sMeIVlcN/NG
kzAwRTPaCz3LPsicOdEGZipHvJRjBQTR9mAfYMK45QFWXJLUUclbPQfrgJwh
7cE/Bl2TmqD45Utrw60eidvh8I0doBRc/JcDVRW90Z5rOgN1jPs7aklVb3F7
UNexvrCAoV2emABoneo7y9ncG/CoQlgV3qe5+1EyNcKy8Wi35g0yzi29fDH+
5h0Rc3mHcowFNQUlS06MHNOJ3N/MHlYSY57fppH1IHsm/m/273fZUvTyryMv
U3pjSHt0KAGP9u+4QWEWgLHh4mVXtVSMqf1siA7zEJyDyrYNjrU0tiq1XqaR
GXOyYE8xTfIOkvulKIMWnArCgWsEK291PdpR0zrhBGeDI4N0WYRL+kg19TfS
PvCTRDcSlv2i7nysjSZs+wYsyB8wOmKclMfVOtEuScISMgQ9Mn+RQ9vXAsqx
o8SvI9oHjilg5obzc85sFS3q48pMMZkeXLN8sxIzO/YzYS/ny9abbrXZOQg1
PpPPQS/WHlSwAT8ubSqiJZmCMmZryCIUJgun+fHVvUkQTNzgtSQQTSCJsT/Z
TrQH66xy3kLAqb3WnO0JJsttg8FAdPugv9nVP/CEyMwctUZqKR1vsXnlw41I
b9q4tWNXJRd5zjc1FSXON9dGYQVmPmIuHdKizffaCeaj2PVQ3OcNHhtlEgNz
VTPJrt3GpBEOoiuEOCAqfmkFJNMGumPAiEDDc2KYiczAMGTGTBANfYL3VY6q
Ux1nO9/qzKRf+7un1ax7/9xF+T1C9zlaLs3TzKLLxyV94lRvBU3Fs7cN4fPR
Rz2J/r6zH8uyk6yv3LJsQtZT3Q2hvy8iBWhLE0spRxMI4qxZelg8sTJz6wvX
ypoLkETGy3MlVx7NUQyaPzqdZcFEJBF4WCizG9pWDXqY//qFsJ99ku4uRxSG
7zucySeJ3hNBI2N7uxYl1rXUXPTwN6Q28LeNrb0jxgJprS3y5gj/g6guyC12
eVeneRUlZIZxQxJ7/q9VM9J+q79YiwC8d0T6eo+GyRh7PApyNE209wzqStOh
5ijuS1fvtV4xsSBnz1oGtmlBgJVASfcIScPK6dCQMTUfCQ5p3Rxob6YzDEbE
YhmxqqpVUhjJ3Sav7LClwEXJENTc4ord1x3eA0urTz9Q2Z2ojzeSgsTdON8U
Kfvph2LLzYlVfEU4AUSnf0mHoZr4lVA2aMI4l2IJDoXkhig8ldxJWUAJDjls
XQHUvaHFcbKPySfXQ3r4ykr5csmzwp89HHx3LknZLhkLsmB8C/VMckD4LCsu
Hr6dT2mWaRlayiKsupyJ6nRZTSuLhja/m78nZDTcW2oymhklBS7P1irYgEHk
rLvc5Y8423ur9gqSewdsAB/9ewAMutS55+/CqgOQneUcjxb9jAUdTdUxdgxc
B2Aaa4wKKwgFoJqLyH100C+rspbI5iwir8R2idcuGu6UtPxGnBat1KYMbpIP
4n3AdK5irz57gGsruD4bMwjdT7RFMEtxMWVgEQz2BC7D3oyat8Z86izcIodb
Jr85lC56+34Q9BaP64EbDizdQnmdC8Q4Xr/Mw+mDySRsIdLmcFjuKGKMHwmR
JR7eYcTnWru+XvkPiCPRUm1Z66yrcFsCPP3r6rw5m0bpEIJW0kLJP7B7N5SK
czBaMjhQnrNNI4VmMmzFu+HoMaz00A22GvUmR4IvgMLQZe2iXk+zt1thKNQ4
ua5HWOjrfqu/Pzf8DCz5H9JonoqGFUEWhlYFDBAFdBaKscTEOROXS9CAFgkC
S5VyPVZ7Lbw8idCYth9A00BbDek1NS11HpIXlOuzffhqqM6+p7CceNkV/oua
DC6O/IuysKsDj+wbIN4xvyXmZ7+Hekg80nQ3MH5DRN4ETcoocDALC6MgJNEY
2YX+9oij3zAIRJs7M0IGsqY0Wi3d0cLFRgBeG/bcpZLHBCpCpC670sSf9ey1
b1rMH03fGWfRGfiSeSyVfTFPApNRG0S892Ov7+jx0zqAR6XZG/+zeUCWTaO7
QnMaIA3MKh/K5NAfleQ6J11+suxLf6X9qZYTYrPaL1Rv6XRkJ0F/hqKu0CwM
eD06xEWiEUM2fvMpxveKclselbSN/RZPLJWbkODAwJ41hT975KHS1rYdWrXv
uemrOwOerxu5ujuimx8pQ8QHXC2ha7Tv1CzOWJLmUlkH9wHuQVLXItkW+vpc
lUvGIM8qUVc2goTgDkyozvcWiwXK8vRUiR8uyfBshWWJhansGzJrO9ghIRaM
Bx+7OHTlupIWLxxVcwST5NG5o5EaER/AnQZK4wKoqMBZf8+SkPB9UCbnlyQ4
92vWA9WUQbcSXanIhdPMFgXG6zY8qAXyBDGR3sSe9EXrmzUivkOoVBQbJaHa
EERztNaHd7JZmumLIRffQPQWYvV4t2xPc5jFdbWgOUgi/iroqU0I+O93ghW5
FvgaZWmh+yNus72332Wy3WZZgQ6Lbcu6gW9iNWQeNjvvBjvEBmnaqEp2STqy
rM2P7Rbm9+fGgLUsWQ3c3I3neqDsFfsukXojxd3c8uMFMpLDOIDywoG1SBAb
/vwBmdtnosiGBHKfF31weKxGFX0qwmHJPbCcQdCwf26icEzFaBDV6fug2+Bt
oy6Yenex63bGYgNH1MRgmjUEGKJW21wPKgIfeLyLzkxI8C3RyjMVVMcd6GVU
XNmkU/CAMfAsYCdztNe6K3yKFNvdSMlJi15bvF9u3SX5yu7ITRORpImnwexc
9k32D7wcGvxzhv3OyLFoNkM90ojgS1nfpLNfTrZGXzB/P6dWHosrYp8mAB0/
d2ZGtgIQlyv+IA5RwDNMOkuCZdxatzkZerRgV256Je9tunzn6nNCTC1SsQyN
r3WDy5h/Z2LT/7ulN8TGgFXIikbbkvkE/7NwwV8kIIGdZagEGewC97M8sNmn
EIArhd5HrHL1bms6bkNYUUMtSDJdlt40xl5qO6EVSEnl4pbrzSbSAJ8gey3d
rFv15vT3UCFf9CbY8btcBNS4yb8qw/B/5ecC3uH/XEtiFr20dVkagLMmN4cT
uHpo3bLk1CaTi/FWF+OqQICZvk45XwrkEoeuY5y0ebaqb7qblseWylLRE7wx
gR8pbswrn6+R0NDRRo5bdrisJ5hsOKiMnw0C7y+usjQ3tZVsy8ITsoD4zm/b
iqIcPKq10ETf/yS032xyUpdNesMidBCP2bYHhubuo+wcP7BrwDBhVRiTknDg
g0OaKxZzmZqswL8mQicagWqKrbktfmLEQbmVJxdE0F1BUEJQ40e4jp2rVBxV
xfrZOqwwdSpQ7gBG6MW7xYolrEgZBLc3hD3fgSgaybNVYFdRXdnchzjXdL1b
CZeyIrEqwZ2YqjAb/ZPMV1lGoCkJlIeyMRCJDH9yR1r9OJkQBzyDzraWdsPu
tJ06UTAsywYA0PFVFtRiFnJD54ddnkjjR7JLRrUN4mfNnml3aq9K8zyrcaUS
OX5l/dKvnLbTLVfJwkKmbRg/JQJmI/NImzKdC8BKcvFx8ebRF7n3NVKiyv6r
oWgu7rigke32k8hWn/dsSjEsvOx2xBg8P+bC3ecZYFbaahgRQ0Sy493XBPlv
g9oIcbGWnhnXuBgQMhCWSTlj3ZEiifS2M9zM+O4tierqOlUkM7Uyka3PhjSn
JciFuiwaoaQX22H58fc4F68iB76yu9ZI34vJMthH5CJpT1usM1LTb/AdFrIZ
Ovndvi+GDcH5K64VdBgT32HnFgjLccxjI2dW8XacjuFJ49jTRBuAj6+Nf1IM
SvcbyZgh+GsvKQvuoqxM53HWDHamp7yWZLlbWa11inppzQJ7CSAZqI90r6kC
/j79pZyWOLL1KUf/tmj7DlLikGyZp/2KDOc9mQvL/weUR8tfEf2Tp3K5mDYC
PEuHhZ0lHvBGyBQm+5YI6EYJ2OrBFo3p+qbIZ5IUpMdnIkAgya0RxcrN3upD
VyhY/jxZtptX4P6KVZ6XRwDWQhwd4mpt9fCmkC5NYpyA5R+Fm+r9QlPb/IGh
jlA0hVvL4bvJ5dbsSlrclCwb9mOcyqhE+XDfUYMbpO7jzgPdFOc4/w/lOCpm
+bi/Kop/v3N07g/K0d2H/oUflQ7S9PDTkvC6zpJyCSv/GqQH9sj7BZoDHpxm
lvrIJ2IcbUU6hsvaXMUnphPIAcwPmu9K0yLka7xEyKRkwY9XAcyEktygN5aa
wHzVDui4oVgozaWtN30F17fW7KjSklyrLJKY4xf31BZVSCWaPfxGso1FnEk+
vQfZTWqv2xfW0Bt0InfGcQXffWFmI1S4Kw6OyptbSYGs5gXku72lVQCF/lky
jDOXSVLBxaIm6CQsYsttyYN98uPHJ3MKmCv/Ru+BxgJs2Qp7vnk2PsBWjRwH
JrZfEJ5rgCy14XpD2Ov6eKkTCJpfGWmB31NUKFOV/26yM4x069z1ZRoxZAve
XCYFp0O6aoW60CWRa3FAm1wMtXUpQe+rySl5vhVEmX11qWG3SZlPHrIMFstT
kR5ztS2CzMTGE4bOBsUc0l+6zfwZjUvw//nJrNE5XdV73B/SFshDB8bYxusd
Pk8r0URnbUJvlBjJ4tva5Ou3bRTTQMzFfyAICslOa+gth0EVVmYMtNAA8e8+
2Ci/Ep8QqoRHSCyqRNr06jt/xDLZxyYZ6BrLeKfQIsC+r6eqyyYIYOtrKwkU
Hsq9rhwF8DtRgRoCXTdpoGf5n+LaOAGKskgh+sVUzoF3hp6fiHPNSQ/5VwcU
vNcSkE3IGxU8X76KelLOaP+doP/L5mX7f7dKe0FcemfhxTPYhMW38B8rMSmd
ANSBvf9XKxZJyzdH+sirttpTY3hCMbFor71DMDGnm37gBoePXXSS5mwVO/8p
ONw25Jk2ViDcwCpcY4oT9QFKzgzIQh+ij1AG3Q2wJ5MUX+6rt7BHs0nfSWL6
KEzAVc+cXYh31F0gcSPGEURn1iKoXCXC6AkhC1mBsTrbuyWaKTI5nRG1zZmW
ut8bTBnkfuLd3kaz98YPbdUF/evLv2egYiATyYydmHHpTaHMBlqJ3AJRiKFh
596paOXPzkGWQ01uxUEW2Xt6Ia6mkCYoVOFlbnW3EbdpuGN+mgLzjVybuadi
1kuPeB8xkBFR6kyRRy3dp43tR3J7z0AmQZAif4l0M7Jh1L9jXFF3JNf7llf1
F0TSnVBXIjBeBuObHG0xhTgYfxqzjOKTT9QVVLYmt1MstOhq9GqQtdBRN5vp
Cx/z29eIS50hVyneMcv18zjZeTX67vKC6+dhOhFhS24pLWNdjO6HNBy8WxEE
3jK3eLKGxaB2Ggd7zCUquwO87O6wh86PXpItxm/l0CzL26QGdu/AjOzOEDgb
FVswfbp6wQTfORqQs4UBoZg2ofuV2I6WSKnU0zfjfuiOXuJIOu9TNE5Tqn4h
YHWVMES5zK8JS73y+gCOjaWaJmQri+tgfjcQPwiFHrIK/iy77WTY4qWi6XdS
6MzQ/ZkDJ7wVxxWufWfca2U5fj1h3KhtAmX8fNSdDpqvPaUrvNUmPXpqOa91
RBxWH1cJJicOm9P2JIV9VCo1pvUDj2SgFTfw2WGXtybw7EwR2CkvaIjm7tml
wN8TXZ5XqQBndP/56m/f74twYvXMk4C0nD7QRN4fi96vBuJh4jHxOLiQpLhv
WFQutMctno/HSZSJzK9xzt/2bNPy4PrUgKnU79Bu1aVajJCZQsuOFk5iYSEr
c/4NvrAtJOIB5fJZCeYiffWX+TL/OlItzIT9AWiRbGPX5DEAHWX/h42U0D8D
WlU9gjEphSA/jPM4XAB3i0cPUy1Rb3ohKrSUL+dwHZ3kHV4lZc6ccNfnwUqb
5zrCDfxrhD1MA+7iwAAoXQZNp6yREPstDNtZBlmm1TzxV5rKRxdwmIpGEu7F
Naw0h574+fK21NQP83STWZbdzqi8F1fBQ/2A+1a5BsL9MwTE9mD/d4pwoAbm
6liy7GAIIU3c4OyFAfF1/7A3JeJsQWCG3d4Ieh7fHMXYz1AjEV/349WOMrF/
C9IuX6c3Mq+YlctKu4QQJVq0vY+9XWIN5QTpAdKkpdAZ8fzbKwrD4CNY2BWx
hiybwK8YNO8iCPfJCNRfNvvpdq4Sr5bR99wSUjLA5ua5WdtsjfqFAG6RXNXS
WFBHsSAzcdbLizGy+bgS8evc6n2Yk/hZdjH7/uh7Hpiswyv8VZecmKVF8Bf/
J83+D0ZfVxH6AGXbmAab7I02beA63GnNq6zuF/IkosuaEzDQKuveCNkYj6t7
FcIFR6JFxFQrGanxo3pTDAYudBPlkhnCWNGwkBqXCgOM4Z3xZf/uNcwY394l
McNBDbqET0SQwDI7+pc+TDzxKjf8RrT0+CDUnWUPEvRL9eLepMeuaFkcFEkr
Kf7DKg7bV7dA/ss6cg+y0lEeqNM5VidpQ5RhuUwz2SV0qvTOGsBcDncbfSDk
u6OPuEdA6vhGUMUACZHaT5ENnA4FNfvrHXPNX+6upe+kfnQ94uOlehohgq0u
FwyGo/WFooNvSXN6vPmNj0GtpAvdsxcft2bnmnUsqYRKmd0onS2PAMODIRXB
zwoziebVB8pt3ZCcKFSV3+atNQSlvsDlUV9fBnD2ESaOqAeXi5Cx7awbj54L
I/dRqHHMNQGB4XMd8AVlJCvUbM82Nsf5FOcFKpXF8IGnQB8WHVxdxA/AfCuW
nBwffk11oe7yMXK7ECOSjykvRIoPeyBnfTstaw+fD9YUNijFjfGLkFWIoAtd
nUqxg/2U9OsKrzfPfzBImbFhx0nPOF/dA7gpyydJqnkmSCtLWK6+yXYFV+nq
l7yzxS97j0z5KEjVzgGIn3WIezL+UjWb3VzzcahwUVAuub5X4ob2TETSdMv3
ygO8o4YsIjm8x7j15TdmGWNhWH8T2k7DbQyeek32p6dzQbKayqgQeBjP4wqE
8tSOGXObEGOiLAVZhzoPkHl8aBj/7PCAQQBu9pqSI6gUZR09CA08xvVZpybW
9LYdZ17U6TtZ809pEsQ09sFyOpyv/rjz6CuSavuC/4ZY/JAjfcMJewrCORDC
cX2t5lcuy9+AMO9T52OnCHOilxzjzCgUoFfMrGIaEQXwUIiSSNE/goJJixeq
v3f5tnk8Vy8vFnufs7SxAPzJPs0iDazXT03na3vdHdozAxX5hi3dCmJOabk/
Ct38h7wwMqF5wp/6480XTPK7/6l0mLjD01XP8k07NAOC9oy9KRgu4R4ArAJ4
bwyv3iaUvmUAWlvhRiFTf3kNs5P2B4Df3LeCeodm9YxNQRoGuNIh4InVrtF2
+CLaQKxC32mZEIMFxDiAWTCFqNOuHsCsnU2dgVcpwRw4WwyKqbpxOV1BkWyS
Q5hAVXXhQAFXCmOYO+0QacKN5Tq9YTKdLsqc99SyzjsiT87eB6N80YidokrC
56mPJOOfPRdOctLDDPt60/pf3cCELmrfNo+kgjQpWNm36zcKBbSYvGN7PpM7
aHJ5T5Aj8SVdx9oRNhFBk1VNAQ+7ydTEGmxMT4rH+nrZZozh2of1xmQXibsz
pxDcHpKj/M5nMf90rMF1TpRlrPYXbDlFH23caZ3Eznr8gaeTZteAQ+XDdUKA
zDR4lGIHxgbrrDffDNlEfpadmXhu8MMEIceI9SokSq42hDj4I4np4BkB8d1T
It++GS+JGA4gMTOgtKtiHluJEjevBzcDklYyHdil4nJDTq92kBOFLZbZ6VLc
AwyR1Rcxiv4fDnFK5lP5OT4wx/qfQxWt6wcEZWJh9S07N+WOs6l484wHX1mp
w9LxuoRyNBGE5xNkGXA1Pt8UG/qlmQfSlGzUGqXsh68IFTW4uSAfOesuh/m0
LO8XCb5F6fJ3QhB8HFrGqP5PWb6G4wqQ+kvOvm70ikGzOdxy+o4jbkGkumD7
51sBJdX2kioPmYDOy+ylQd+x1VOX4HCV5ZkyZbwyikk3kkKr5hBIIJXM3nGH
lkMwT2vGdG+U078srim7M/cl+3wLK85Fhe2NPqDJR0IoNhf4jUdLWEiV+ln2
UBpEmbD7IaN21b330QGZVfWEAIjmvzcBlTYJzcUIv7YraDFHU16do0ZVX/0g
/Vy9a79KAxgmka2Vk8Y0PBlXtLU9JK7W41SLxBwDrYt3xWVFW/M1JcmIfqTB
HXaBQMm/zLCbVgCntec9lCFg1GF+CH1mcPWzGuUj5Rnp1HwHFwqjUWfTfW+z
L7Ev4fyBYB7OZBWDURTH0GqS+Ytc0k+9f0FakKytXUK76HjHE9/VeWPJFv43
SMUpNYH4HarWKB1dmUp6Yj11/jdz/Q8Z2CFsprVZW6kU1KQoa7AQ0bz4JCGQ
hF64eCG++hkinKnlthrK4J3A/pY9G/T+ei4wD5QRujZmBuDd5C0w1NJT+1MF
M7Lq/Qjl91g/+sPYXA3HSD/ZOdkMMNwOAEbuzivmQz23bV6UoJk32nu+Ay9G
8GviMjJxd/3cM1wKYSxKUtoSm+dvK37MkDq6dL1C7xeqzMqS+HMKVwlYF8/2
Peu+Lcs4ZlGEw/uUqguMxdL8zC7YRYFue05ToXqbFL80vkUpgdyb2Z98U7fI
nAqzr+sQa28fnXkmPYWUBGyl0cZBSMBy/HZJXWd/HVNKaByxFKoYZIymYCuZ
zs0SXHqsJnPIPoshz4jyz7rg0sw4oZK6CKNZjbKXcJyEQVGE1hv/lSyqxWL8
lZma0WLgC28Ktr17dLbmois0UrnavndeLp4eOVedg0xFIUb3dlCKVUz11KRv
uPjc5EXgmgXVct/kU5urW69Dsszs2bg0XktCsXoOF15cMgeWjUmE/i0ifWHy
LTGykUfN20lKCfIroOQ1T52OxR2Z8n7vVWbxacB3PrCaOM1mHiC0gG66hR3p
N/JzdfSWDXsCt8DDNu6Ix69B72mLfLALGSs1ApfiZeKXmHIKud4k1qTdaXBg
zc9oU9px1Z/u2y9OEhe3xE3PpzZocaEFArK+B1XWPTsNP3RRlbP3LZ2iLgsX
TzMoZVE9US2Rzpfh1KCZEQdIkGP8jQnL2YLurxbsBVrTUza3RYPGpGjg8xX/
4MxUKcr99GMlmkn1RGirE2d0rrjeQUWLmxCiPwrzs2gcxrPZTIZe9PJjrm8U
ZRH+8RU1mmvJjlH6ekSCvajIknRrQ3fO6U3RONGLb+q8Ej44tkWC8eY2vBaR
/1fRVHtoTxoNjr+D0ncEt6LIodDR/a+YaNikh71d0+hHZU7LeCQxhNOhcbGV
LOB3qN3wmd2t+Pk1YASqG+8KB9cBXzV5a2JZ16fu5eJCSQ4z3ARp5KY2RREe
fo9w6M5DeDtFJbjVzgfsVsSdFCEznit1N82JwvmtVx5u38pXzPps6m4twlKq
8MquvmlYqWM4a0MUwZ7Xg6xVqR4TA+Qqy/JHed20IPTJTGbKjs4GGr6QLPrT
Gj1A7CPxQQtz0eXQ9vYbnczm6wJCg+MOOuI91eAYF+b/BvGOiYTGHRePfFuX
ywkxhyW96sfepJ5t0K2C1sTHqfZ0p+Q0asy2F0u6rqmsj7LMMl3W0axlqNjH
N3k02DWh50WrYPJqYWSYyJjN4O83ovGc3XYOOy65KRYAUtUL2JAuQe6u2Vde
cbiqRmhfcn2k6HG+d0wEPmCqPdGssoyTYf7Z30/ZgzKYhs8OTuDNXrFvlq5F
lxfNDzDUL2fK5+x4Mc8Ec0HTZ4cPJzilH5JTwsLN4UK3hG2h2+ZbZF4yqDEA
IBh4goQ7s84kS4BH3e3MA6N7ZHGAlJmj7UpaI8stb5cr39gfuP4YbG4tEw1B
lWLYYswBhKDOkAFhtaEDFap2UZOHgxuN/WsPBnsn5Rksmvvvl4KVdykMnCJI
8hgcLDAQnxJvNERfLC2vZ5vMg/s5mnuOXj1OOUHlr18fz4czLSkBhw68AFaM
tZKQ1mbs3jXNytsAbTnql9ZYGnqYvtjJ6H6MZ3PbQSbrthudKzstqPkf9K6B
vCts8/P5IsGe5sgT/ta0MNX1CktjwV3vM93lnU80x8f9omq9TkDK3nmJqf39
RLbCautWVJXZBrwb/PTBKOL1aB58uw3dLwWE0ornqAwiYR1Z9h+hcxO46vIF
jLF67wAARRe6H4GjqmieA0kkI6IELmUR39WP3PtUVxGxM/8r26Jbbv5tuRfN
fxHmGBP3k/5QgN8gGMWan7z1lmGwW0/vIcorGoVlQjx8ecjYyxX/BFZKSltp
euJd3bVMXAhaICTxbf0jvlw5YmJOJqT83OPBe+Zsx6gKISs6DjF48fMOQb0e
gG+8kQ1vfyJFCOs9khWsBUoInzvTfpQdCy1Ja+XZnPUY6MZ+RS1HjxqQPRs/
OzTEOspHElXmMz3GKdBtQf8CoPGVxNnYUeBdB1J8RvFsZVjZh6T1QlpftYGe
2fErp0Bn/UfnlEjAINbyUi87lsCbuoHQDhJ11LkBvhBjtvfeG5RXVlSCfG/Z
eEnNCKGTj62JY5pA0sXC7bTyKjr0GFPRkEYO1nsOEyGbKJV8uV/aS48XVw3E
omZ3ky1I+p8Mu75eiKjBFnb9JTY1eLUL6PryBIFAWyXWWSdvuWsn+9rCX5L3
pj404ioIAOTu16efl27jfxeZdfupwZJ/brb/D+NXwzAVOejDRqIBAAOCeMLN
YObIS5ALJBn0/op1PhSi4YaMGzFG4vGfNUYW6jhKJULmF3kgU+/sMKkiEV+D
fEcIeUEz75BfXCECX4tyZFdN5uZaeh51rJU4GYRj3SRxY0qtAsiSL3y+aPBK
W2ECduSXo6ioeNHQWST2ivOYPYKXue7eyuZQf96uzoJIMrsWpLlN9AnWW6yH
EQljz2YD2Gc/XUc+yCehHOGM/8PlQfXryWOP+QvhNLa5f6aiZVygLe9myeOO
8TzBD87sULJzWjunzGkf8hKgA5obB0ARaKctSSyHYJ6RUmUCdgG8PYEIVv61
7ySFApV+KitWQBZoO9p/F7bjCxmDqOr73IzjteEtM6aUbX9o1mEeY0Cupb6w
Fibp+15OER0ZHZJ/3GWXGIGzIPVmdi6fbcz5RA9LlEEsyG1+Whltqxe9ARQQ
9pDxD6mPuoj56U4QsdALUSQ3sSybkgQ7405oBlWC1meDht1zYKCb8px3yWIx
7oSYj2Sli2W6lQJSb/p65o4OV8GTSszgJJMy0aLCIh+LWvQ8/4gphu8fnr1a
iuwq0q2CVRhwBYj/bBxvqRJZ0BlE3p2G9QaxEpRQf37pxxFKvnyUkOgn3Yug
7YtorVuuVD7CiXyoz1oHVC8UKvAuhwVwlZG7VF7gUu8aCLF14vJ9Pmt86nUQ
oPbEUSgXhEZOwixvDnLiA5psrxAjaWVPCU6yGFf+EktmBrXL1VskwzWh0uW1
LPFiK3Cb5nRqP+IqbQEb6vqkBZBW3oQn/7+HGoYW4K6pfdpceR5oxzhnhIav
EhVx5MRYNmaVf1/zJz/zJz1gmqG04oOmKhZnMzxnYtCKy8aDKLuPaUc+XfI/
yMsnyFgKBm5D6sZe9uqu3cIHNwiDNA6wuLL5ucM+SCv+0zLbS7NNsK8iUfVK
/zUwXZkV0ArCC6PmMTAy1VcLx54bkyuoTzyksdaBx9c8Vio6wIfne/rDkpFl
QKyXXrS9YK8urRZXyAvDGn5rF0CBVLPfQap2kxfsk21AVE07zhckc727ptQn
Nh35J0X5TborCt2yVM+T4BAFIHBhPZb+2WhjtJCGU0IQ6Ij61rnWRv4GEBng
4qi5DI6bdTkbf1AV6w5STiHXEsqB63tviq2sBaybestWk7zoLnsV0R/lFoVt
xDqqAB3MH5BKhUNFe4Fv2DVXlO2lH7YWyv0eCtiScvc9n5lcWKVKylB2Rzdb
aakBfO9iafgxaonyNJ35sVc9MbmBEsFJEmwtwxXpO0RbUK77Ma4X5SJZz7n8
xu6DfBgPO/6dwN+CdJEzOoaH9NQuf9ivPyMCzoAMSUgF+ZsIZohr6A8ccJK8
cKtlt0BYxusDiX06Hhc3d2wh79fyVzln9zHl5GDSyLfRZoxXoCO3EwrlWu8q
1ymC4cFyfzGDsyUlr5a92SkPK4aaMJ0usojHfbJM3K8S8p5RqEcKCVd3ohQb
nujguOez+oi2zjyEhoMIJARW1QKOXTSYh1B1qP864uJtfz0a+gcM4zpG9AyG
bBRUjl9qOKwGDTBAT1G2o/bYZ2q0ZsapMY4iVebdvu0u6QUA28uS612EWBQ1
D+Z/GrT2knLm6uGQAm4h1MCO1RUYbCPG8qoS9AaZBYhmAm1worqbfRbQ9SZj
45VBbW1pL/DrPrryTacwr6oS2Of8L95X5jR0RzchhB4bkB10QhWKGKF6Bd3+
624QF94ePwnQAyJ8SrG6/YvhQCHH+Ycn5NxD2iultZroACsl7Hh3v//Jf/ZQ
MaOTfEn1RyYc+3jslL75BnVk9MV0h61WoGEQS8PekdvvDE/fvkjMS57vWUIU
PbLjxQWZQmFXByHyM8rFGGqG5gxCrghhI9SSlQt83FJj79PzRoGkeHbVcQEo
d5gZg8TLGPmSc55FC+XBB/9Cpf60tD+Uqy8a/nS3JhI5eykEKOU97dDAhzS8
BRf+o+gS1uukf/4ggMVaQ4Vhc8XTvUfmgn9v845jnY3iuvhD1XDaohoe2rus
pV9nlybz/IuSaw+FHDSiWl1mz7/9Am9jGogX9gvk1U+I4QNiiR84uQmPhzlJ
jPp4f6/QVYfWtYqPyToYB0Uorv8AtqM7NbOoek0YECksxggHoIWqx3LnI4Lc
rX7oiUIjnKG11ipsBuHKCljgkPSI/NAGwKFr6PNwBx/dkO5gBzAgsFIbQnQO
ZqiGyX4m1vwcO5i+Mqfx+5njihFViQD9FQ14U7t+bHyglIfMzQSd2ad+okp2
uSzhPTiJ0+VGTJt4E52x+zhfUQB52cGhI48+AjlA2iGJgpIfk13oRYnESZiZ
EIYI17oKiuRl/kNV8+HT9fdCSEiDLDlH92Ox8YmDQDJKNmPGSRt4I3Pc10a5
M35vzjLDGFiDVEZeoNJXi6wnGrXlNCb4BFpiXBZDvLTqmYdQVXXRAyiirYYV
6EH9AchQN2CIzUaIrSUWxC1Y8JCv0qEfWV7cnG44aLFAaGpdLH1y4jbKXb2I
QLdEmNrIlpgyx1/g7qyYs8zMdhcAQDrDiP5hOt8pvtoO3gdny52bkjbjgXcR
wtGgEox9ajfGicCXpOn0rftzfS3OpAWyuPu3T+u4LPN0zARaKWo5XyY4OqID
jMvpMB4AP74h3l12+N1dw9KekaGkcxqFNb3CzJ+3ektL/3XIWcBzKbD59SWN
+3k9aU/tekHKn3OULvPmE0sLN5Rpr0THY5eQEIEXjQdMICpmM2XJIt10h5Vy
50QmOblbRucorJ7yeXpyD+IP8Gxe3oPq22a7vMh7UWlNTs038YyPF26fvuur
o6RKvnQEMUebyr+Jyu0paeQaj1RcuVASgssBYEbnM5xdMudL/JEH56/K8ygW
aywYTLvRVYo26FfpUDXmawic8fl+TkAII7MLXnvFSrhcG1xO7pu4AJLbNhy8
m5LRcPk0Mh83AisxnVToBedvRyhBdIox0N8diIxQpPhFnVA7Z+GxWjKpPBxr
cr96/Wpiqn764EFO1yU1ZPp643lC0aH4E7ubRdYEmULOkc4Alk3SbW5fCbaO
EEIimZFWOkLf3sVjGIHzgsAMw+g6BdyZqT5xGBhxeFX/m4y/DW4vqY0wYQBa
C2/gaphXGAfZ76swdICp/wLwLxbml8zf8A1acSWziAkestiH0badMoyNz/ev
J0KbfPLmFVDkKDhieVoGp42vR5+z/R4dYy+19y2FIF8xxJNykGz4DS2YfEZu
+0vr9iaDLXoaxBfQ7SO39KgeIkRbWMOqMZ76u+OvdaH1KQZVtzgLL06Lme/5
OYO5Htburx5lpmcghkibA2H83q3pHxHWNO4uJ56Wy9t42r4tQmhNYGh4xAL/
trcf5gPLYv7TAorOODg7sBNOy/pNYd7IqiCa0omui5n9nNZY6bCEOJCHkao7
34FmH+w9JMhzHvHdK/W1EvOMDwI6+95XpCqFQ6tY4/M2Br9Ydy+POimto5hx
ttLpcpkP6xLkD37jI3jIcW7J7AU5mwyMBU7j21ytsEMAvLwElps5rNPelFdR
4MkAyR0PW4Z5TfAxol5whxIPG8CkDAFZCmKjREDhdL2K24MFZIu55h0MHSrd
N2FJWqnW4ZxRF+PEFboIoSzIJc2CTvOhyfNDoCn5Z9cj7UAkWxb8P2o8vgJB
jxBIN9nfxPQ5k2g7TU6BV5r8Yv3UvbDQ+23XF+c08soUfoG3H77foCV9zUpT
DovAeB5vqDPb/zX54NNktLMGAvOIITldPSYLXO5Xab0SQ+6QotFb1xDOu2YC
OgY2CXHBRPZgdEbLNpdwXP69LIWp1cmyr7ZIZpVN068OVgmANeFUB/wxzujR
BewyBvTL5aPCcwzgoDLlomXNsYXxnEUnIYUUIhhBFpNLQI580TAqd+DbntWy
uF7a8laTFgDIy2JqzDl6d0daVM4fwgK8C0GXMqR4a20vIPk9Y56EmRLWj6R4
r+nFodZIzJ/jGN5Mh1dhMeYzKsJESPhC12QbdMRJVETBzR82Jdkj+BUntNWB
R/+bupgv76j+14LlhrsVXCCQoOYC8mSXGjCq4TJ3A8VMpPiAd6Ya+N9wT8m9
sbI8oMRlTDzI9BI5WU7K9dw//jI/Uj4fAyOk4H7nrlKO8fSKpe4PqCfTWtec
SM1uV2pPx08EBBiAIMCmj/bmEZeB/x23X6m3lYbeG/eqbJPiCEa8uLeLCotc
8p2/Uyt1k8aefssdCrOmi619orR0c0Z5PhpibB5V0Bp56S6LHGg46Pq9C/9X
gp0IST9gDom0S+cLO0fTMJg8UEZ47TD+5dnCEijhw+9hDNI3+EyUi8cwf/1r
x+blHZdGfiFcy4ibCE4GSjBwqTtEcT5qyrx/pnL7X9RQrwXPK9Y23yj7/RIr
JB5+M65pRVm9B2ZIHXNRv7Z0ESxEyS9wJVw6cdda2geEBVaMyLhJ56qDbtPf
B2IQVRyd0yT+91maU8yNoS/NGq5qr4WGQtKQaTARSRvg9WNdaSG8sns8FqBB
+IqYdHkYOQ/w5tauQf1Dixd1JMjAe1yoYwNkFrJLcDzv28IClIIm92kGKiNz
7V1DV3lpBzBJzp0Zv1rV56QDDs/WcOlilxBZeuiykBMEVnbvUYF/cyPhtmDF
T56zIsyAPg8fnzACQtmdCKm95Hj8d+kb6WsT1t918S09BArfumRJcTwMTDUm
ClUHdb96raITiNUrOfnHrAliRZCiD6GGFFe8wxKmBUTzaxL/yB3VGROjXQpn
esH6MPmLooIMMK7Easm/X3O6faT//ZVM51n3wyDaWZWvPHRVEZQrET24hbFG
RH9vximgb1lqZewBu6TvqgbkZiud0KjNS/Gl3Q6AQ0gRsVbJvw++XcLekUCV
nNUQcl3YVqSr8Mn7d0aRAj2gLJJ1WXo+9n7s4Cm2SME2pO9j22jxemHAhYTv
6q3jvRfZfDD+ngrgRV9lf3QlTQXtZtYX36bdyvLg8Ea9f6HlhEHIge/NVNQL
p6IiMrN04t1O2luN6i0iy1HorfDn3iNDI/YRBsg4fCSQ/KssRDMVGeiCVyn+
U0/bRS+ji+1RMwHLLsI21YLCRlMcgn7LQ98Nl67mp01gwbNYcxolxgnTRHU8
XJxJnZaDkryfHf9HFI56ILfnTjLMSZdMAJwS5K84tVAzJQWlXk/r/F+QiFE4
Dv1mgGNq9EuboPwcxjMaiqFJo55+OS1RwUnS1xJRhu82ud1z6aEPlMMY6eOk
GXEUpL1gJo0YWxlzxAGAQrCmWxMA9jmfqUCpt7oT7e7xFluSCJAx8Q2N0inw
f7aj6oBJ6KWn/FooU5Uc1c8tZxhBVxSvmJO/bUSnsHdnJK17Q0M+I6VPRPTL
I/711F1EZheHhs7EVw4xs3vQuygY2qJVe9JKfkfSp1FgOv+a0mpBpteJCXqh
iyaOKM8MPUw6YyB4HKvqYliQWSguhtqesLy37rdrQpO5pKhh55wR9e82kFqW
4fEbWY2Izcc5LUZ3C1/d6O95TCBdi5xSIUI7rNXbGR3l5KUtoxYKAeaPeELp
M/mWv8RyswIGBP9NHypOoDCXRTkSJcH7J2od2QMY37nRKeTpZWfyeEwb3NT1
XYP9+ZdD0BEhVYDgSVBNJAJ6vBUP7m7lPfEW5ER/fDGZEj/XmO3ydKyu+ZMD
p6fhRQG+7rqNa3NqdXumsyfurG6XZGjpIfoPFTOQUNF+sWp46aOxVHJotmyr
ATfvMnCvLF2X0pZguBJjX5VXO5uB+4C3izGfyDSv+lBB9KAZEfo4STAQzcwy
6LazD9S0k/ZdyNwq1nuCPJBYAIkEw/Szm/GjfD4JcC3CLEQoOpMMoCkKhEkd
YV3B23VJkkxEgjSedqJqLioOq+HI+CV3GUVMRRW2NcFRnB5hSE/aK7XWhpSn
cxEZl6muuoQtiXEd6A9FBhgviEAzPyAhGl6yB868joYnwa0rCIJmvSh/Cai9
FKZyHyfjtiA/T7e22MRyKQhj+8iR48wS36vFJioIQTCPgEIfdb8ZNSepU/Ia
gk2Q7tNq4JSAM5hlHFggo8zTlLoz4Tt0JQaQWqSsnstGTqtRGzA0acQfCN2e
e/JXmvek6nVdX5UMlbK7+ajGvyDjzPaKEdtvAHLp+JZPUSODxlwV9nipIToc
LY8b0z1CiEtReFXDtjUU8Zk8WUcrec2K9o4TLt9gbJUGyBIaTM/yD80nC/6+
VPRXxxTOBAgQaqDmywUOPsVrhdsA+xWH5ar4GvcoX21UF+7O0K8PthuIdWqF
7B4ku99omxoIvqbMmJgED7Enuh5GIzYlvDBTbPJaIchKtZiJqN3QNbhSD0Ix
lV3GIgRlPnsi+0zQL5c6pjEBAcH9YupS6SYcgxN+l9iBZuzRBet7sf2ER+Wu
xhqZAVtj5fkMSYNM2i+t5QgEyHUDoG8UcGhvDSkBR0S7AvR9AL0TRINA8WEf
IBntapCvMlLomHI6FaWdoi0e0KdQD0ct66nGx/exUhLSioFi8d07JagGwJOL
4dbYu42hXhemz/hsyJNJ6SMo9Il3R/J9GglF3jMVAXOgakdb5qF91kGtWFdt
F2kmcUPsia7WbDhvxVPTFUZKXPEfAnxZsvsXv5X4Q7yCqW20G0aH4fDcXt33
0GCHjqgQc1J3wdSgnd6ShzWCdkp/oFLHC6erQCfnhd1yqQH44dKAfT5odkEb
eQnUnZqsZodKPHcYF8pEexqasf1UBlNazAZlt6UPmLQocOS9XMJoBJq0YJAb
kEBVcR4bA6Eieu7tSFRC981ZP6PmhrCgg7psg2+PqkAkbI7FgUiQ5queppum
IdFtLO3iewgmjkcuSL40LnsrBXIW5qF9r8XI6rDlfmRNDhbrgyQwNC6CTQ+Q
NPXjXFJI5wt2MrLzQXf/zvT8c1Wq4m1r+pfEzpLyHq/Uv0qmdMlmCWKbd2F+
l3fGymnUrOF5NUjBCe8tRNLSLABNv0ExunSYz6hYG1gCnqYsFMoBi7RXIEw5
NnZ5+ncMuIw0SXuCi++6tspJ9Xe7F0tgPKl+RKmSULf8UewRi3hZbkYaeniU
xMfj/E5hOFICTvG5u3+nBpCQ/S2UJrbn84jeO7AOcZrB+bQRfxstMahHzZ2K
Wtf/986tMBd9aIxTMFKyvYVPbaUYw6Msm8taJLMpwZsjs1c/Yx/tyPwpB6sz
DWNoRCw/J7yoaTbnVgCglp3zikFj7HYK+bF+yNwpXkDtX3doUhA4/JRZ1pLK
+ZNeolRQqdAr800os2O/jKLOHoxm7Ett1UjVRCYp8PtMX4qqptxEv8UiFNHF
pMK9hZeHezrk22nrhf9b97OGUQ05ZzbaOrXuHYqOPz8qYElr6b7zI7VvEL1Q
QjDqopi/wOONH2vda8HlQ0rGBbaXOGETjcX2ncK+onkON0BAyD3IxPJXVYeb
yZft3wtslRwccnE0SwE7503roCwvmrItypZR+LeI86IZeO+gdoOk0VOiPYbG
WRAE9cf1FincpaQuOsNU4OVoBPX6SQcw92R3mA56+dkfUREkHsbc3EXzbcZZ
7KRrX7uEGAIjxMCgcKI+lmFCybB31V+KEIXH90wcjBqzjtWthMgw7/1nk21a
PNEm1ntu2yaebzCyE5YU2h8JJ4P78dKMTF6OOD5DMHmM8wNwBEkM5r1ZyGES
cCq0koi44diIyR7tLwioeUbkuGtZSd/i78wMa6Hl3E84Bt3D+fyvP9rJnV5t
j54/qB+083HPtGvuqyuH7ydom9GlNGcHyFU6akV0igZk2MQhDdPSTUhF/FfU
Y8XRlneiDzEeaqbfvcCLB5jH6Gs/gJSG2+PHFhltF4xGLCMhA6wNLsqyoF7s
zeyGG6Nc9D09jC4RTjdGyUzGmZKLaY2JyRes44OOCtMgmUFqg0XJ62P4MkVu
weDYtkwWYF5mrBtrEMrhC2CiuIWWCtuFv1F4XTViezXpxn3eXWwpGj5jXL/C
h9YaGaCWc4htEI6Ldh6OM80yKkGhq8MzImm0XebDbm14AXaTnlxODmHg55au
NuGvDGUn3bbBk+gE4eORJazwylnJNUnK3vg1av/EHTSWQBJtPJUs0tIg6MRI
LrcNyTkjWinuB4hYQ5uqfrWT3LhDBlcqU1J3aqirDuyM8cCWuNy7Alv5CUaA
vZmCN2XQ8zWgp15QB5Q6hbnQdqF8m6i7dYkBDQogx8sARqWFOJ1KyOsrpHuN
4NTJZHC6uZXjj1c/v6zrUkRZy9E64eAw7lja+F/8NZCaQjyKwC5CZ496fi5O
/42XXERTsrTI47L9DDJn0xL9uV61e/L51jrgHKK7sveUAnjU74DPLtuANSMc
RTaeVUYhlKDQ6hUD0LkYj09N1478sXDMTM71UC4KJV5sTiC6yFbGhxSUxDV6
Hbp1eN0iTAgsBRDM0kBL0vy2UswPp+uc5KWQ0urF1L0xKxsd1BJk5G6UDmPN
HjxpeTveuePzI2c7FWiJxUq+ya9KKScF6CE9jvgT/y9z2LCU9/j8twSVBTcq
eGnWMt0Nj7L/3s0mLg8w/sI2T4XQHJRqWyaEhYyJwzLSYr2u//w0gzQtAckm
+IvZvbhj66h0md/QfhHOjKbFo+nSwWV0w26kxZyvRUUAhuGy52OTvuHSprv7
ky/NuY6hRabkucTZSbHGKUFtCvqz/jDqtlEbtTI8Ro0jS+LNn80rx2M/6cOn
3OTzD9ZWjGA2kD9MuZgztK3t/+6fBNKc86yXXOx22BavOQieOmMVmIx13yvU
+gw4Hfiyhcw7Z3ct6vdf785n+UYct/l7Kv69Zc5VSmit+BNzj/uRY0et8Hbt
M4JIe3YW8my5qq6IHPWEVVNcPlY+0CgjbyVMqjRJ4U+40iq0F/hSJFOgz+S7
hPy65OU/9aj9o1B9m5sVRM8HX0Tz0kBsUylU0tH4cP4R4gaZsGiR7GGvpMsG
H5MUAu/lAZVhOdbaWoQNBvYtUsrnuM8ypjic857DXrMpn5UasSwmXwxpe9DO
2EP/pUnHOIW9Flop+fsVg4S5H6aYFHBvnqPylBtfg/Z1YxOY/4UX/cjqmgLD
MMd6AZwU8AEb0QRpnuxBo1SOIeGhSefrcUF5m1C4DbBXORgnrWwVLr35J+We
bcoSzarlSW0l4xSc2YaJZGaBooiXU4mOHz4726gOQAx2KKrUHkOi97P6KZvF
0MAESdccNJcmOX2A9emwkBWawn+liWtv8lO2A9dXkQRZrC5Cagc9WEw4b0U9
Uuf5u/NIcKKz5v6DoYW+LHwBkdDG//0J0y2eHrghHZDjY8zRUv738maZZVFm
tBAnhjkgstyT5olHPnNWMl3wmtV8G9ozhBDtnJocaq9Izj9szeHbUqPJwT83
djEUKV29hK87pdw/VHJzk376peIMN5HdLjpvbeWDfu1MJTOHQJYqjApmdy2V
z3XTzWtWCDye08IN7FTazyNNL6D9xJefjATXUUoUftTQv3E2bk7NltT2Zf4h
X+K62PKfJensfuYAFQsxchrqdeOaNwWigIeZiPVzhQ5bWuU+RSycdewNMFyz
m8bMRdMZaStI8Itb/4KYoFIiSKITEfRqg1dbD+BiLGLQkGtTuFYMqWICcQ+2
CFJ5d4FKMwuSYAJYedeOq/CDceEdtex++YDLACrD4IC7nRZEa6F1PKskpsQV
Xe9BeJLIvT8XC6u67o1T8IMIzaxqxXL6XrIoigXcnSDc2vKoZwkkGCsi0BfC
c/7BMSXRZpdXbf40Ybh0rnfKXNFDUVTB4qyxMvq5//F+zk/jRoAPnYD3dTv9
X9KeHL9tGruHjNxbNg53lyKADRoJrBC40VKG3aH/YRsyxy1ALEUROdo7hP2b
TE0VqfMwvYcxmIeLFZcDjhrqX47RZ0JoE7n0uydDy5BHzgTlOujuyJGGhrm7
W/1bwOZ6Jz701iEZGZS1nLs5ulEL5Rk+ou0NSM43joew9uhKe5yhUqpk4bfl
B71kkyBlqPrrlhnCNOK4whTM62xv00kVRPAh+J5H4QeMPZ90V/ZJ4IuiqSgA
rtjjUlHezbIvH6BUhMxL8ZG2yTs2TCmDeDdiOsxU/FmFG0YePxCCk7290tXC
DfemRxnkOwmNxt4hkGE22X7s2RclEjzJ8fVnqJepKQebM/Fu2Tz6zfxgQJEV
7Y0oisDrMclK0CDxPysh4/Q5CF7dlikG+hdvplBgPr2P3POcGvxoYCpXZkAD
wFZFTR7vgmWyRRaaIk67hSOe4OM1wId/7eJisctaAiZoEn8+692cM00/ayUv
9V6y2Q+jnrTfJFAf15ieXfC/x6KmyG9GRd6fHEqQ4PSX0gqx5rEhn7ZX38yt
5JGidkojfQm83LEtbPWFbL96JreLjRFksXnzXy53H9jNbQ6nNIwSr2V1vKBF
F44RvGTk7MMRGlxL2ykMmBUo5mekqjBPypex8hEAHs3V+eJ98trKweoUpKN8
FL/YfN4wMXZk3DALfyp/v4U9tAxNeLGdziWo4Zajsje1R96Motgsql0FtawA
qXJh2oeRie7sNQf3K8TWXe2oysu4mmZSdj/DR74aNTnTUwbb5h9BlktHNb+v
X/7EznWG6WdXrm3eIybVhTh6gYdelYLLa5H5mHqpeD9MiMJ3JnYq7MdL8Ouh
lHmAOB2IOq5JM0msn4GwQ76vnor670GgVkAPujqMX1OufBd5wndqrdyLVZ95
9Vop/2d46NYQAhjfHddFPmyII2nyOZui3StEM8vJGuDwFfAJkU0U93PDU07h
2SMPnjH2+YTeF8rOqHunUiI8J5yfLDaygkMTga2VL106FjVPvd5HtOTawXLi
aRhKPrubIJ7UqQuJ/Nwe6MaKlMDuK9Vl1WUi4XrX0ysh9fjZFSNOTUddIiBp
QXdftMR75pXz/Ax9yjnQNMGqFOV3wH2OubLY90osCj9grA2t3h0PZjiePXRu
LHHTMKWA5FYUyuhICPrntJqc+4EMWZshmRKATiJ3aFtZw/wS4RqXU0ktp5FA
DA8fxkZGQsKOMQ2rurH54Pt38uPCdOCBieZ/hmk+aYLb6csVZe0goU60x0bh
mi/eMmRTA0arJqkg7qSGVC6VRLxgWs1j0oc692Rr8oaib3KUfoEapn4IrdKm
y4mbGh9ie2IGLx3GtFCwqjfiqxpYL8DA08MhdJlbE4DC26YdzfOPgyQqy7fK
s4Y4EfaAuFqUVlCfFQLJRUYAhnn5pZzWHSGbstNqd6SDGc1MsMvuAdYtYvnC
Xv6eGqi1hwVSeKphCrmEjptjmN2EFZDR8NC0lRub4g4YdszvXYRU2FQTTKy1
x7c61WUC1OtqI6vDiNARywjV2gpGCn4IqbPxwKpaSNWLvXkO6HjDRUcLYmfc
eNmyuTUWKqsjIp4B91It/qRlDnshyBMjhD0Xkw7rPuHycd9Ynee+BMTx4wvK
auebjUH74FVAhGDN4Mgmz9PcHxRwDzfj4xoWIRct7btDXqbWMX058V2hV6ws
pOSjwE5vzws4PMKnnVglWrSa7rUc4fR7OdxRsC3JtOSsX46COdoKevGFId1u
a52aeKJPm09jJLkzznjgczeLvmW65JCIUlhUHnXxpv3n2tXXhZEx00MAYrm1
wlBPXPWwiaCR5j8zJLoDHWMBR0PGiOuIGwtbmgb7Wp+Sqs/Xm7RaTnVRtd1c
IDixCB9KyzL1iDQh1J/1GCM0FSM+lVDQkhkk+yPcUpgNX6wn/lnELBqztPrf
vvR2s1bcWCap58t38eCAzrGEglfEzzC1UEMiD/doTq45WB1knwDHSUMMaCZN
fQ3LjpJdXTekI4CXIq8lRGxHyT1fqGaLszHRahz2tbMvnEy+fwWPXGxusVSS
5BaehE0gkA0xDbKF68pJqzjv/woKpHO0jn65H16j6/WW2CJZmehK3v3oDZBO
AwysWwWlBUYgUVNqSBNElFjsw1yXqSIx0ylka2DkvKzGbB3eKH6qfftSq3vq
ZA4hzSHxrsART4Z+88rrM2LM3/TKpiOLr1pGbDLmXu8Qur2/6kZlkITD3V7x
iJcbiF46cOHZFM2Z2njd1qlLK3j/Fy1tfE843WlB7ihOuNar9MhEDCTrtt9Y
Iatuk1Lx7w5UcdF1c+CfiRgGviHY6JUYoMLrq6aQrsjqdJyDHugUF7TUs0HP
uwYtGr4HUItAL4HSAK1RDUggYNJBMahK9b6Eql1Al4NOArFj6QERpUod5b7O
b2ltDUFlVJsmpJspxY2RIHdNTqT1Aa0TbFFI9IBSGrbImOmQ7ntInMUTh8wb
yuZHVIk2mw1oJFQLP/WhxpiqJAYHT7E47MKbwWcAIaPIcWK9FnJX6IlGWK43
+dV27mJONTXOFX7SffFDcbXsmKt0CXIhntuv+xKNIRWZZsY71xElop1zPRZd
B3ZJGYlMNHvqQKPdzgWoKcjRaFB4U/g02oCB7k5j93ZWaaBzgo8htpGi2YHO
UlojViIyyPLtRGDxQqygSCZB/fUTrxvj/72mHbMuNwQiPjQqQHx/f/6lUe4R
eHyBLygTRBe4JioCIz9R18wRrcaJePYfvyM7GD3TUY3yHu/19yLY0JfBbUQ3
97B6OfiT0KQb9xJXgQigveY+6KKefB7VMnYjm2FzHZtaSV4f3+Tw1b+nIAuP
BleYkWcFvqXHsEEyTrgt20SmZkCwphffN/0ecYZ77Hs7wEZnsCvOCDCENdtj
CiEqE3PfsQuJH7/XAAtvtAWWgD4TWHn1wVOmisZUvCdqk8gCdw36dq1/f09c
2eV3IcLnigXjQ+wRk/gTclOpVcTVib5qFPS0L1AVv18p2uhh73lY1iO0pcXc
4GoOnxADnD01YtqJA4Wxl/Ka++ukydx7QO4N9d49P26qRDG8tuJLbZtqh4q2
SokFjcKxL5W4M08PKz4/2Y+vmdsn3jcXzxChqM5JYB4BeAIP/jgLnaqrN3nb
GPcX3ykkqb/x/a1Mot3QeFL3dzkQzb9Uc8FovZwCKLTKb/ASqKQDcmaXFc9Y
UNumVMe9BOJJ5vv+jnRM+QwhgGVS2hh8Z5Tk20UaWpnJ3dq2jzHdtSTJ2hkK
3q9zbJKEt4p3VswSgmcSz6TlgdVKdlTPMf59rFreaa+9D447fnpEVVXHpq6F
UmnI55iJnhDbJ2wQJ9CnkpJ8az/XHAuSJ1SGt+5XMGCPJ8/+2Uc216LRkq3L
Tt37S5LCGekKYCwzYGPMpBiIxCLY5CUwX+aCgocycQSpQ1aUtZSv6BVhe0GM
ba8sMAsrqv89IZvz2Uy/arkY1uxJdcbkuyMZhR14Ztqg1vnyceNnxUIYW3bg
weP21SzdLFndQ7E2vpNfSkfG5RiAZRlBTwBtouwmUDmZgQqetS+hZX3nx6mF
g72PFeEnuT01jYKesb8J1JuBQCA3hFYC6dR559V6jt3qNZn55vefSQFPM4o1
ECobtNzNIly7jdrNyh3kO9zXNjWeIEYzURYhWQYxKiDomspxd1ZmIsr1AvoG
FV9IjJc2BekRAOh7J3ivP8BwEsx6poM8rQz/dHcQDVhv9n0Sz2riEsQ271vu
/6KzcSz/0207BKubQJfaT+bs8nLLRA0449PCn3YKKTXnLfqZdq81gO0jgjr3
/tPOgvthI5vqhYjXl6y60fJHvl36hvf/2Y89xCBcPm7JJB4kIjHl03KNmtNL
dEtML9v0G+12EgBjhKh4WZo7kwgaHgh6ywFyRuyB0PIVQrAp/Kajbxr7qBG7
qMCGp36s6btyAr5FGHSCyZf5j7HEjRmRWeRPckh/gX8WB5hSfxwXQrWyn9IZ
2j2D2wfzUL3n1X8A2rRSk2QvHykNqmrAjSmPFdRzxadKYtM9c/eJ6fqcyxm6
MlGtUSfmWhAFxz3QpsGwlZyp9+COg/AC+nLaJKp7RzyxwoiPfj5fyXgEiTWP
0V64TStjUofAib+JNDkBYgsDuQdv4apDKFRr87+4WUED887gLpGqc+lUSRc4
TGDarJ6J4TzbfD5aP4zM92ilAr3oiWngyb/XT40QVg7mI+I4Ke6MMqUpJ/e1
NDt0MuffKq/p4nWlNPO2rps9576q60s5qmPzwztb7b5GpCCjN+oF0nJr3uTn
Sjoxc6hFCMyW/kqghBHplw+kBy6IdlGArG9CBC1Jkp/J7EjkEsq9ae1cgcQj
/DlPgC0xzj1BctM9uGY5dK1K4XiZdhQGOBZZpycNoc6NZdfnqnRcoHh/JEps
QZCCKhlQs+F8Qlo3CDIzoAhrjJpVj7QdQVs++LdqGU1Z/BSrx/EK7u5Rg0U7
chexaESqk8Mhdj9l6T7SjClPhQt1mjdbf9K2wqRf/J3OWWwGHCzuxSFum0BA
0nD8Q38OyeGvHWXk6UWDGKgHA9dPI9QayVG3YQ+y038LatJt0sU0sIyoshCI
1PVV2Y6zN6pQFhtSghmhhOImJtwXIRGodf9H0v8DcQMt66AkOEuDt8LwGBvQ
mJtm7LWr0WcyRRAuttMvAPKFKo8kRQd1hFqwWq1q/VMt1opPBrynYisVs64T
L+Q7b60fOF0K9+7VQj1iptiG0PXYjLNIw5BF0QjULt/BA2NT8/4AbXADw+Vm
k71IwEJ9MEM8cxeXiDMDPM9w/wk2zz7pQo3PXZtL22/6h+By7BLz10hQwYx4
EK+cpNKKra5oN/b0PbYy4CKP7nYLGflb8pUxj/gKErYGAesIrcQLt0BHnIwY
MH1fmDcBrivXQJGCWURD1YYanF6pAEn1HbaflnOvmCWyQ5LzqfgZJsrJ0IRY
MP9sz2XaWOKG34MesyGm8pYbrx9waAAzDGx7QK1jRaL1xWi7FjScgCg4zSql
2BkN6k4gWP0scEuUi/vIsPCrIk38aN8x/V1xvOcIhj4qAFG3hHmNE864nRik
hNihej/L/I2Z3/j5veLbtpjh0s/ZN5+6U7uW8eq6Qt4o98kjUIkZAOG6xuTX
Svs2Yohh2NrhuQoCBvCqaMd8ldeN84EYD61ACl4tTnwXqKc4q4WkAnUy0HyZ
GWzZ1f5pGQUjUQZBbU/Fd6A8EYOF7L6v03yESM0iRDFn1f+UpX6qF452x5Fx
ivU3jdKFE7aO4L1XmGY9Fz57iUAg20pd5amPYV/2S6knFi79pGiEnMeJcHM1
ht4iXocK116rGwgz1CJROM42YV90iCnAFp9pU7VhafOUdet4kKPM4xLPGQVS
ycdNPm05R+79b4UIu0e78TNjS97MgCg7ERf1MiKautKoJYmrYnfTu1X2ow+k
2OCTAxidrVfebnp9MFPObirUjvsHV9nyss8WHPbcvHTgmynSVT4GjhqczxRS
b8qS6RrMreZqm++aTEu3riODobV3bjFKLkOJreJBzJ1rJbjqUJ+2HYiLS99r
GhrGGYf9To8Ju4k3GPLtJTD43s3wfgAN0bNO8jjfS1ZCWatGs0YLRQ7zbJAO
aXHzGr17RZGJIHrS/Fmo9/nfrs8GEl6I2GCDSaIY+UAKIdNLXFkkSE+oqVsy
CNoTNCrNdKDR6g8BZuR8t3mxSfValQ3+Kv/gJL7J16L3UHn7//6JFx3+JVmA
l3jeGePGTJOyLDj3uiueH0zzvKlx6nApuFKg5KKUKPQiXXm7Y/U3kp1bGQR/
2zcFijboUuN/2eq/0DVINxkqpaE8g/SVc4+MhCAB6VE+zU33LZY4aRpv6eU3
EhzsYgxTvOvimxtGaMk07TaJKdFW/tqZp3EbwOBBdjtq7zizx+trbFO0uE6C
oroHMSt3VvHponuDz8sVSRzbiumLstMCd1T7Ad2s+7M/DNd/4EDcFOYqJLfh
FjTREH8zrwo0lKthTWZNt5MAfSyD4dGYZ0zkyV0VXzlUh51AQ1FF/yqGtrsu
XgfOpJOgQD4I+/Viz65x/nHRt2sIKF6XMGfDPjgpDhP+fF0RTuxOJGLnAjfA
SqSeZvgyUNU+fZp/ig1HrG7LK0243lVDz9enipjq43qW1z5XzvgDpWmDjMUZ
UhzpIzboAtq9d8lZZJ7u352+N+P9bNTNJiEcpftBd71EUdc0sQ2PgPFDyEgO
rZsT4qOr1NvBajRpeE8OZ/+a5q17yY3SVx0M0aL6ltuGGJ+njCtlUwAqp5MO
WhTyRA4ORubtQ+IYtRA3EJ7n0553/h+Ti0paom1XxuBQOn5PxspHYb0+GSNv
7pr4kvWKLeWPTdDlFeTaLSaCR2gjdArpGeyWhBEfn/ltZJ4ZludDtqZ4nMJR
tDSPRY5TfKc9P0sKCh/iLzHa8kk8H7jJMnz7mBOGseEImKMe61w5KJAvV11Z
DcjVYbi4u//drWMZlZkQGkU3q3/av3T+VzexBuNKcsUkA/VAintOvphBdhYs
+ZJ9w+d7oEd0dl3LSHP7g/FkDJtIwJLvUTZQSHbh3Ox9r/FRsZnUOnQUboMh
t4FMNIGtgn/kj6EajMwL9JljWh15NP1TOG/pgxa5j5Tmw+9bJ+L6Jb5KCtVf
30C9GAtRo6NtotVy6oWXAJhsmCs20SoYtjRPHrksieOoB23t52UIoMutbzvv
djQTIv0xqHDk5OBGB4Cb+HE/YwA5MQzP9kaTa1NBGXtM2ZvL3tD1dPHbEgRr
LW8+96cNRVjX6a1F8RXcE94Y5UsL2Bb5S2WRjlxRyC1ajnKzgRkQzNWXq+Xq
qzNuaA+StX+VeWUfBZyGUmPjh+y09na7jEt/snemQYNxX9vnz0XRaRC6dHY0
mgQSxv42o9K3wQLw1yjBM2keCtYLZQHmQZzoh5oNfhZRwoV+vFuQjV4QKfH7
YshjWhbNkw6T7GJX4IZTK0pGzePR/BibPiCc/oSRV5RwiK8LFPj2E70A4KbM
ZfefvbxbqScS5pqQ8zMxYXR7BFrfUqxuwdIme2Wt1ysoFc0/SuRP830Azm2+
9Yec0NilUfaZxycyUvvbs6WQD/Nivcpb8seRdSns+rie+0VVYparAuPSmC0D
G0v+WPJaEMjYdIZ2PywHpUwd6IVbjzBuuLjC8qlXST9FCy8KRgGoyM0kXk9T
p51eQY64aKnBWTNWDYK+JgZ/DNJQNCi4CFxxjkes+04r+rQdyTmgWR7XFYaG
QPLBQRUZMj4mX4mqsXMl1a1hToPLkw5JLwTRlonCuNbzF+L++CSCFmzKsCf0
btNWirVeyvMIuJSKnN/wdKbPwKe+1vdWFnR4ilt2BZHQEvzTngQbUJxU0kZs
tSOw0Cd6SKl5bWpfWCG28iPo7/6J0rn2f2JZT8jHkjCx4ZD/EbP3b3640XLf
Et2HSO4QyFXHnNcCvuuv+aU1JTfTYKtpW40ffxFc27dne+3Imz2u3wIpq0dx
fPznvKNzylFrzzFAQXQ3B60vt+v76BzHX+pXkPL+D7Ro1826FA0ycc7BbFNJ
tuI0uRfrmchSEriSkNTOyOMOgSHr1+yQ+e/xWBMCXg6iiCWCB8uzfPawytzX
p+iR8voy3lSsL7MKyGssYqhEGGCNEGOxIcpXIXneeZBf5fn5d/SQmBzm0pcO
WkniOE9cRtDc5ki3JrAo8XdmoMVRpC5xbtwFfAG2AUER369syb5LXvnaZV1v
a9q/uvGMqlap0suEiCK7v/BX+Nzipq0H0RoMX82AFjjtxAg6LZU2uPnIeUQF
8iSvL70epZGqzKkj5gZ5jKnh1lOv1+YFVF+Ad6w74DYY81zOglUv+t24oK+4
8NxvYZt4K+diCTteDMqJWHBlvQAoGtYVPKKE2XIgkCdjcrhZO4kb0bEC4rra
blvmS92OQh6gIxgRA3j7DObqmxBJAfUT7A6H4b8dj4lKiJamSYu5lK4XQvFr
Lpxo8zHE+RvAn/yr4b96QZJ8yJ7qo0kC+hrNG+1AlqUpikA7TM1pFc4YV3Cc
u6vGCMFDagSdHFrhy5Js+4tnWKB9ERIS6UaGrsfj/fzEfDQXQ+XQdBcjWkHz
9Sm0uJJO3g3lBuJHTuntuBcQYdanweCukcG6he6MDBnlOeXKal/OVLFZC2W4
3uNiCnzVinJBHthYi5VHTXkyn4TpVn0NhPUooQ7N6GeAR3UWONpPgGZXjl4S
L8NLXPBveQbO0zuBETV3zbNAvIW0oRkVYpuzkJxYTfCLyNj1O9g1SbiheMeb
K7rhbp0eU0g1dZFOTyN+nmCfIRdITyGwQu9nXuhqW+MiW3DIeF1th3FlFiE+
ciykH6bPRSyzu9A9JUvnPAnutUtCWQAMEedreGZCiKTPBfD2nYXr0tHO6oQg
8JIJm3PBqeufKka3mlegwCl/QuWm4Mz1pZbGKtbligMq4dwfAprAD7AX/Mzu
A2tY9jWdOg2/aOeDkHCW7nKBBm2AwREaXLo0HIblekefcOmFHF0vtuzd5ZkX
qnh9BdjkFmcf5VGpxED7LmvtIYo27nXixua7m2E1fiNP9+vxVkO7KogbjEs0
pKsEtC2CQLZ2uDjlYLJGxk2M1qe8HBZ9AaH2DQWZGgdphqusXO7E/FmcZOQU
29kN4VWfBtZMzT1ifPb3pMNHnNMfbRsZ1dV0YaV6H+7MlFR4+KLc04RxGMMN
vinvog+UI9u/lxu/86nU32a2S/UBpguaplg0biGAHGrWfXX7dCBuHY1CQZ0E
FJMoR1vnVxz5lJHuHTSuH95XnsvAW7pXv0AdQx8pD5461JUkRLcefcPR1VPa
e1iAeg0QaZdiNg6Sq9C65giJz4a659no4N0abwwf8YGki0G4MojTlVaEW0Vs
XH16eHPF1aPNxcY9gOcDiKkU/0iJyJtY6mLfgWXW+mbDUue4ry1tbNLTMCFF
b7oGpoZMFLV7WSatpTYmq2/y3zZqbxE4MKCOvgx1sIl1ZFbbdwaCh9WKHvIz
zZHkZ/WETq3K3VZhLkHUvpc6rgxhFAiS+gEI5Eg1xYJreKZLE53oxF3p8yZa
2Z5HSrzRjCdWk2QkkGPqAcL2p5xkxwMGU/iE+bZbIiL9pxSZCuBGdfEePiTF
xRAc11L2gBEJhhGwRR8cySP/xblUKnmIUKwJ6sUx/bZ9lEwG912TRTTzHgbn
4m2anJ8fT241fsGP5Wu1A/vnFMJSaRLZDjeig0qKTC4Z8canbpGsipk55bPP
TFoo6eDRZc4fyp8QlEg5s6JafY/Z1eOT7ngzJUkMkq5rETcwsgtWTcR5WF7n
VH0eUi0muOa1hBQ1p8GWm3sIX3rO2k0M9fO3klMEigeC9IWHBTGW5r4WXxJ/
xzI2pQ15JIZig2QmqTnm9nH5tjotwjUabRF4ab2yTl79uCyGGNlmy2jeejkz
gESNcDCKZiyE8SEgdOrUKPkplKiZkwwAeOikUn1doBeaKfhjp+pL3vidtMuO
MDnJ8LWSrKL17SScCvextfqsrHOubyPB+7XYrv5WpIEqOgqpI/Z6x4YBAwu1
QzVI4po7jxY9EBX0DDKOB32cnKR9JOLlXWcmS8pzULPslqZniyCY4NnDbC2O
42LlNGlcN84EOMA2Z1bOMD0boe6SHp+TieRAvApYCy4qFYxeKY5S556EsotE
Br5W+IPZ5t08YYPosBgSxF35d4g1gl9QO47R/kYIzQYnDUf/GQVj43tqM6qs
RY1/MT6hcW4bdWmSgqIBCqcmUwjFFB8P/M8RPK7DYDcQ6YbnG4a78pNigcR5
39TOdIrnYRX4th9tscXEjvO5DcsiQn6CAFmjtAbzUpd5TK42fKtiYeeYEnpZ
ZPWehz7o8TE79wbYV6fliwvLJF62QDmDP1rdgu4gGdbJxbrlwOmsotEjvGxB
AHlt2S46dbiTpRuR9SMBUmrnXYX+sZMLVxdMjYoNXwowv0Zb4JhP1JSxgkH3
Tv2VJYeT0319s7qXj54nxM8X91Wm26pxeQgVMvX3ivFOjp7pysGlyU+PUuky
IA7ZHphqndTw3UnhB3SVBje4F8PRhbe+9HsHvBoXXuA6owAm0Zv62eSd/A3t
FpXsNMQEtYjO5M7DLX+YI+0N0mVrw5misBcWKUcsTewpdjBsvAmXX0gAqDug
YKiElSMfPzBtOwv3bXSkM9K8LUwbX9hKgS8kWtrn5RViXwzl61nGKB4w4cvr
M2xi7/cR/RDDV94DuGIh22TbyKiCghtYsJONIpY0D036gtdDs4VdvNdsKPvD
15wmGr5ObsYltmX+MZaZ2hCK20C3P+D1uwi+mEVmO5YIS8QzPdfIKzbUbeOD
6CNpPeCA8SiEr7KiT4SfAtyEpGr4qBYbsOZjY0AS7aCWRrwSK/yOwKKB4LnW
cRdMt9chSHj6gcuQqkuLTACh4imHxGLm/BwWJ+uJ7nD5wkZXLua8k/Bwo/xJ
J/ZJs5jx67pPQfewLYW06SFC9/JG8Fp0UaHExupoeCUnaDHUrtDtvlLjf7Av
lvhP8gabpYDF79AfadnouaXp0M8CVQixa4l4GXiNGwnJumH9fLl85Cui0QLx
R8F2CP6G+VorUOuKJsPVrmoCYwCNYoz6332Sj0/QcWaDJGyEIdWt6/Hj4F+k
FmoiUTLTcLy2DLRts/iNwJLYEdDPgnhqUUcftxgL3wfAmxOL8hYP6Wd0TM3x
x3LyXstAcTbDD1GtHMZl1vBWYTIHV+mbVUaWPYuVJUYLUGQ6LTqvvxCrBuPL
bRMIGt5P2iKvFBAi76sEiKJR6UnWUuNHCXNbXr33P2OMVR5pG7wcc2ZUUrOH
HgopTBZGCxiFoQn7eQZkb+ycI3YYb96m8fi2MVc69ggNjsP/nA89tymd5ca6
ik37fwYU72EORG9elz79OKY7lZG2HEDNo6lFUrBVZNZLLAO1HWq0D849ForE
wIMlACgJnegN2oinLgI1zhrRmaclHQ7OsnGHZPdh3lsxWAOwy/i218smisco
07ENo9ouRMrW9HZ/fp2pUaePvM+mSrPVtTlgKIzzbnAFn2cJZFXZi8MDrbIy
6Q3pJemNB7w+2vLHZgE/xtXL9tesxYFRFXSpTa8oNEqwS7IUwXgC90MEFaKP
c4SfU9Ls9InDfnfOcztJxbm2eB/1uvVOSGHW8XsedKT9um7dkeL5mo+A9ttb
hjZWnSRPujGUmQ6h9yZTZhIH5novf33SqFDzXy7SfBj4i3dSyovMlKu1weaa
yl8g9FpDFUfbEdd1ZZHebu2NOQT8I30Tl6GqeOKwoveXozxnbo5QiJIyTwWH
ULY4s3Iug03C4CaSu7CTQN2g1xq3jcQ7r2ZQTJBJvRR0ySlOupskxfB/M0ez
WK6ljsWw+ck5SbVVLPiq7JNwNFEn3urgszQ5MhChkCaEWehV4eKMF8n780JC
x6VzWsoOsY29yHeAjNzftaWzfy3bpWGk3IxRs0K9nE0l8nnSM0SEbNtDiUfD
mtplwzcDlwoSuF2kBVoqO9O9NPQolPatXVo6xteIhQ+pafNtLN+cf8sVnQZG
NlY3wmmXycIERuiLO7782y81DFm89QGXDC63NYIYD+dX7zQVxoGuUTYJ7BHo
XQ5/2F3cVU+drFa5PD9utmPcc+XcO0r1lecKtmRPdYByorFQID7c7y7JzFRi
cHGkDFdHeZlYbLngRazui0ti3xZ2RY7bqXiXH4IGCc3CrBvkn4kPgHY7js7m
sJByM4mHVlhZY4dB72zOA9ERJIJqLhvzWJvfyXHWDN/JyJOaGPFAfJ819AGh
+ieNrrK3/ZBbU5DAKaQjwrzkFqqLCaiHe+cQ777Slk6S7HnHw7N1damET/dl
q+BWKWUni3OW5LKvajqzWQxD5S0UzfH1x5gFVmhS3LT/gfQ73Q/1GnOH7cIV
IjgayXeOu/rb4o/E8BmZvOWoEvUrP+eTUbGEwR7xuSKf7owzJR5qFjvQXgVF
hT10pto09rBXZanOUUhzji15Avq4x1p0B7McJop6P68A9l3ieydmEMuvCtx/
P6RXPe2GQqN4rZufJVrteNvi1GmH4nGY0BYyZ45qBtshLEpZ7bU90Vca6fKo
NNn0mI/vOjzOY1R34JgF8eoF6Zt9Nv3ZYKRDgjFahoiQHWuBZaff0EFUJ6b/
s8jImOJVhG/Cvq4kJjNRF3LdaN+iYFHqCl0HJ+gdLiOQMK/Bw4Ialaytjtmq
pDgle5JmpXcaPpsEX4o2k2EXUnqdA3In8a0V9FV9S6J59bxsi1yJn2uyiAZf
A/DB8R17lIm1pDXGEbYsZT3s1lYEGGwKz0A+CL3zI3Nm8zTeevXMU+z+cqBM
SQuExe4MG3WeYKPcBqRcxuoTEPmEcoRQeeOIwWn7rb/7TyQU5cA4/hsfUjWP
j+wkgUUaOKCbh3kgpYagJ2gyLfN2Up/EzM83Xs59jkC9a5zZsDMnp+IOTpDj
EMUC1znPmkYoETmNtW6dI1SJ0fDqeiTQ0po6X6yM1roQ4TdCjhta0+QqN2qR
1aGBjU5/yz8OIfF8vS+fI2l8qYKeon58aKNXZ2PUfJmCPWJVYyx7Al3pnePc
iQQ+uME8sMgYHsVbCu1anv4hfrprGlOtYNaKlZmUlNLYuDKotV7ub5edLKJe
recsVFSldeCcBtjPIleNB5qCIA7LY5hjnLY1LybaL10Hoq9RUC+97PzDsvY/
WnjbuJOleoqS42mJoGirVo+cST3+m+jiWsPtK4H9K64YrFmHtdmsVmV29pMT
VlGvddmOdxu/y7AFN8PzjYeqZ/+kWp8Emv6NrNGSnftKDKrTWTMTia7brLHO
ZcH/hWI8qRb3M2aKqtOI89bATiZZzP/ytkVmiTNg0jGkayihJDFt+xnPCGwX
yMvR9KSyxjLrbAPD4DURGoTzCn6HCZvD8PZjgY1TBini9F6lIEuP0DC0XlOM
diUGj2uaAbQNH8DXYbRJ84qtq1e82Hyz6vK2zXBH7W73nK0Hsjp1uF5GxxXn
gWi9bRdrBNgD3hnY/wGLvZyIimfUJHMOf9SVPa+Ep0BEudjlVMR7fyNF26+M
kYoF8mW+oTOQCkL+OmUxBf9vkxccFmXxCxEa8cPxDF14NdM8kq3ZydTI0FTe
6BU3MUrTJcPeP0LLnlcqBL0fP4Hfyi3dSqElxkgQuRIP3H4VJG/8yhjug7+R
EJVisxI6dcr59U6RrqaW5ShAR5jKWYK8kD51YzC5wIqxl4xr5Qg/tm0ph7nU
yIKTPfDVQXxSmuc8P2rswlO55LcP6V1zPU4HEd/4+u6+HRUdJJPSiL0lwNhg
X4mjih5lPZx6OcUajN6ZVAYRhzvyTB37XBZRMVThnLPa+PFDBfASxINZlHyS
VD+FPUpH/4ql1Ahof6SQkwd1Vw1V+3Xig/+Edrorskyh1p5HiXPePJk7wTMG
pnygixjneaf3OMP4M/WVwBxqGQSxVA/VPLc2lpLBYZSxtHwTWEJd80aUS3f6
QNV1JBSGGlDh3TuuWy9oxB+vQ3Xig1pWVMxvavKBAFif0W4YikijmSbxJ6JL
KZynpr6aN30zx5EZNAXpXvJ8LoWq8Ir1b5uSAejbMF3gPrduq37RJY+Do3kW
cpVpWNpNits3oBx5LQ3VfndhkhROGPcWQLBsQch0cO9ET3MQ4IICLN3xNlYL
d/7jTSC25gciXcYY4hhLSOskpSt21cFph0LDOvn0HDemLAA0L54UEknShR8B
Uv+k29Wvzvq4ZcqQY/3YGPfAoM2f5IXfLuMyfndZVOubjvi5zrlHuSz5ehj6
tb9AqSD3eeY/DTD8Twrkoh/3dxCAFvRE+nNpHDUShQB//s/JaGXWstqJUaaZ
IFYW1zQkJM6+kTGazWiio2Nljifh+DHULZOi+Zx1iKjjrKlBsDqVyWseNSGx
Y6w7ckKVQ3b1QhFeCLd6SIXQIBe55TB9gJ9caxgQ7+XP14+EJnx1xZ+dDOn0
F0bqRtAVVCBTKyu3APWHhpoXvWMzWO8VOg9VMKUANBVaV2ehSycCqVDJ8+9z
jEDTAAD614v9+jcvKF3yOkE0T+lnjlAhKyyE3Wco0SycMJJ7n69dx10QVGt/
uN4iGriDsi7ZXX0jJt6Dv/4KNsQhpKip4xCRBdXlbjZbJQF/ONvpoP/3NpyI
2a7ZqeCunwIi+aeDQsbrxbSfYxLnyttuvlyI+UO4KawEh7Mam1tUH1ULxo1V
brm5JmkboBxf03zBUxMTtzVwBFzwuOHYxgK3jU1VVUf5z6AVJRcRAfmVZrNN
lgVsV0tgf70Gvd+dbnxplAFrn60Xt1Cxqzkf8NqJmI7KtW9uU1nFo91isUX7
XRQsZpQWHBrNJF7p9cNZXMR7roQXSdQxbBfugs7AfzMtysnbM9mxGE/IX1+0
Udz1zWeX2NDnVqEvDMdw4IWSH6kfYNSoQGMGkdpaQr4PFfcuCvL4ABK5xc8O
8OI+GihH4Sb9Q85JvnfW59706gky3NsDwJOa6PiC/5B8fT20MpkUlBv4vYGC
1sOca9cSEr5jhpQSRvjXI1h/R9WdhFJi4NbYkBHOqF3Cbceo9IlTvEquhAaD
mzXc+ossyMlhh7GeCeQXRIbgZb9DH8WbTl2xaW/wCaraO1e2SFykMioVEjK0
G4nfmDkPfsdh2/wCV0JuzfRe2f88haNV7PSLie0JioRqISDER55fB17bJW1z
R17Q+vNWN/bwjiIlbJ7iKRCvuCJhtE3ZVKxSHtorab5Oam3d8CeHVk61iaS+
+cJ+xtoHQZfK1qzYr5UeuL/SN9s7rUEkXeQeIWIBNVmG3vlRWshb5e6GJDEt
/YmEs2IfahKOr9LizVsPNCx+q+cxIhIpVTD4/Q/aY1yj5wc2lke+8/ba3F6N
jGTFDKfrpG2wCIYhfHaLd3fKCqKCdbu9PDzuBXTUO+jgwmxGhGN9RAVZfP92
XWrnXEkv4CTSMArtvs1b+sKqmYawp75WHTXcso3LoNSawKf0VsLYiVjbxvFW
ged74R+0jM9HvwTCUws8VsLDtrkiKytIbNjXMYeWZLSkgMjsK1642Qma362H
UGb4O1az5xlk30BYDYR5d2FGax8vl6gqLLTBeQmtT4rR7nMDtxDyfnnPM/f0
vKXi/R4+Eg7eIxsMRbvs40MlYUHxvv7URTZdCvm5zoVhqxzXEOQIUrZP6Lh3
7uKfOy0TOXrY586UxPsdF/WkdN4crC1wIPDB2O+nAHip5wKSMYbBy3tToxgQ
+mydMEEyxif0iz1GzaXvWOuFp+pfVV5m2ABYIJ9/OMJIX89uPamwb7EbjE0K
tl8PSQKCB3dW/Sze6nvKQvc2fnIIvURBut8xOq57V+d45yE3JAZkdy+uljXD
Jz3HcxXC7CWCvq45cVtX1t9sUoItVfPVn5vzv+n+z6xCEyPrY1o4NTtlLBmd
9tXmujrprt83B2KVjXaSv1gg3X5aeiDM9qDduk7jzVP4yGG4nTRV6MqgPKGI
gpvGqQ4bN95GoQ3n/HOaalitGJ5ylgnTZZPYE4lFfEBgbBIXHBxeRmcZUb1k
GZSgucNfiscMT6eK17WUHKeFrgY9w5gvqKmnflW657ZHvWVzNHMic0AwZHa3
NwxUvZDHS9mnh4dbLi7we3k6Ft4tsT7h30AEl/lqoSCtItZZ4uuRsJCbO0k4
rCbnuzAe2VSc1G3Q6trqRB/qO+CWNQpZ9+yOX+7pPJSzK7EUsYonR7aL/jBY
WbeHFE86vLAkOtYAyulRRfkC7lQHbMsyKyw5hp7RJ9cx9wogrE8smgWA7Vvm
DsJeMCmpZXaAeKGzEFRAKglkp24Daf39DDgosPL8Iq2NdZvJuRPohsVdh0fs
1cqj8V6Uv2oxtgKYL0xQp4Q/0v6pVmLm/Wj4H3ryt1dwsO05t4imL+rRLaHh
0ZJmG6jMNGWbsPIE+pmO7uJePGQn13/P1YQ1D2ozQO9O2PnZ5J7vMoom9zEV
foV+MQ8ST+I40nw8gCEE05zw18t+EYykwmKpdTUT15c5M/Tb2j+so3LQltht
FrNA+Mos+Qq5OF51RW5ANSQfrZI9h+vvJ5ndCqmpU+4naa8DqZkNnukCOK7x
9v/OqktkUeuRHhcXYtFKvvThUpJU8hImoRjMEfwKXmvNhKc62utx0K/AEqOF
K3Ul7kppeKaVZjzaUH+NPKJd+uodXhGohLJHJwvUbZGbi/qDf6ru0GP+xW7T
p0ulZB0/M/D8/xN/TQSd+48HSVRVt180cTCSZ/7KlGGmGAISKeYK7r0Yml+H
2f8WYqmWl2CDRWBapOevjKEdLamoO8jWTMuWohz0cID/FrdjKyemjYVUnh9a
Rc300By3hmQT6QURY6bbWSFcg99QPQteaeyleJgbM3rYLIFVDUM5yxfTWp4s
M/ezHrZgMZ5msezsQ+C9/ZFbiMa9rh4d2DfquXzsYbS721mflBYKb2cGxtay
bQVD0epgBJuLyBK7ycfViWD3Zu2Hpz5QGAgJs5+b5e/KUKU9uByduRTc5vhG
1pVRqu6Ei44MFX+hjZZ9ruzjAmQlvvMBRMgv4QX1JlON2O2fCkJQa6/iUU7A
b5LOSIKtPbx4ME9PE+NP49sGsZM0+D4HXf/EXnRAjHRvhbAihetnrT0sYy8K
c3hHD3DgpiW9b1nje0ISavsq8NtAYtBps583KLvH+YHSkmAatqSbaqbVwkEV
OCFd/J1/cPt7qNZO7hou2XdimUBjUzQ7mLt+eCcfZ5zOlJrDI2Y6Kqg3IvrO
CwqvhNDRP/ylQEPFrKR5y6+QuMpzw7wV1K7wwHAgvj0mAsPYlQqOAt/lI5LR
2pRtiUXutc+fIRsIsJb/8NflkjzB2mFWTsLHb8Fk3Hs9tXPgX1XMtMkwksU3
Y3SiQ2d2pGtC46wkclFauRf7fRkXc9tm7I9VYcuw/AaFO6XA+1wSFvyxXLxa
ZVCcoBwCi4P+G4CGVpYqP2Zj+XZB3UuS2em2DPGfatb36Py2fpVGl3eXWUV2
qJi6FSxafounTPqlE58KFaF6wy30MGs8MJ9ocOzR5iPrML7TS7zEOJ/PCCFc
s7Xkoj2ws/4t3VOlgZoyaK7BgwvOm9k0D080JrHe2v5cK2cSfK9N6AnzVFqJ
BSXN8wYS3FqljuLsf76cNmT0LYOqa0q1U0DNXmlDVL7fZbVUUaoaBDSCk2yi
w+3qvZFdzyoH/PInuvNxPKzKe65sGbL905cjXd2A6OVcnsHeELcZ6Nahe3OW
SBGccRwycpmsAwBVODngf5+tJe/CXjFGhJwmYnIPyalkunqNA9tCCavelm/j
JKSWmh6I7/15eKuPBqey+XDHJv43jgyYXtmBz5ykx7LAanUaQ+jDVDgG8P2T
/V1wwVb5XLX3bGURbu8mykm9Vs1psFFwVCwHVazFcJM3DET5gYkLJNL4nfOc
K0zseZuBN2GDxZ0abAxfacV5ay4PtZQMhlBg34kv4nfloeXVsqTpeOHwFDpe
1R3PYK3sBp9Kc+fcTNn21X32CyfUdeWdgFQdScUP9gRX6w06q7QYFn4SaPyc
DmjaYpjSQkE+OoJOBqMwTnzWR9pNM8vNIYBZzIaRimOqPBjLvrjIb2Mo8Kxa
pUOD/+AH56+vy411l7bdJ9xXfbIT7Kd53x+ixad1ixmkXsVhTp8lnaJXkKPU
tkHIX2heh/YDaC+ujX4JRi5wCmgKyyp6HLpog7z8SuanY7shXY4QtVBUo2Kd
ZK8v2fUvX7doGHIaRsz1AMfr5Jg/0vfwKekJKooL6BPJyDComCbw0c5KbOQS
gwCzsnuolyFN1P6dfpAUAc1oH/7zxj1hS5CzLZLyTvVtwVv8/FQrmTXtqK4m
QOUf3gq9OARCznto4W0V04HENCqjsxCc7og7KwmJQ+c+ZSPT7xTLErPp/9vL
MTqpPSMmM2Z+lh8zgYk40GlHVRUdzZR4oteLiAn0BoAujtVksNzoJ+QGJ7X3
iUdA1GyR6VU/fiymop5p0oKtZhajDX2eWYb+xRhMrwZbHdSZuTuXgpx8qxZu
44PuyahHAqeOW5qwbcZ8oLU341aYhHZOnoYGIYl2isBSpEml3uTElgITrpig
o10aFjgDLsu3Up41nf88rVhxacl7ZzdfMxszU7Lr/VBZXbOZWDFWDjLUiuXO
CC+0M6ThT18WSFvU/rkogsatQ/u3UcpwuNKGGl0Pkd/tux4bD93gl4xFXMTT
GxrQkTNmuwgv2+GMi8+ccX455r5uo+CdY9mt4c4fPuI4hYC3EPJ+PAp1cJqm
z/RTxjqXq+SFvm6ERoNtIu4pSG9Mvro56MM7veCTuvyVWv4Ohwx3sfc4jOTs
zhJm1qHXNFfWxiXFwzyioYsfxa6iMHKybtQ1Ej8eBvkuhyhOo0LXlceBo4Q2
kc4e9cjRebiB+2fBHisG01i0/V8sMuFJbVVTUcGLhZbNCEduEaIAAwo4/iB5
EoRMe00Trr/JJ8yhAxNB8SGRyB2Ij8VzqxEEMYGg3XySAVpW30bqAjyMJJtJ
kJbc/pLEAj2RUg32XYI+kGUxPhgJJoEP/tucXgg04iMmtFmW9Wh3qfnfpiwS
QnjReyHEmh/2BeeBtYHwaxdpwk4G7P42KnEVaGY9g/LUpyPD+0sHX7Wb10Qo
BDAyCiKAcvqmcsqfv3Y5ZGGtC5UVeB6Nu/d7VgyZB+HikWH/hjVg8PmhR0eV
9r0mUCMDb5r5+X8TOnd07yP1nmGPL7UupjrGM5+GhTw9sClYNxfpmOBdePve
00MJOoJJNZqiwB5+gL1fCXiv3G7kGNS4E4g53A213PX+ZKnlgLsTYhgMoyCQ
y/cm5ocEKWXCbrNgxhFKOI/DSCiy8U7osZg5nOtrq+qRiHET4VyS4Cw3ejPk
6K6ZX7kwW9UiMifSykOQUCq+A7Ncdk9XNSvP4A6y7++eM+thRg6hV5CeD1zN
XuPqJ/EfqttuHaPD2LKrZmXWL1ph7+YC3pN29OqH8S76TgVC1Dz7m4Ywb3rS
uneXDSA0lvxUBTcBIeFhfw/3coWHlMmn/+06+ls4J2PpH+6JdoGr4p+5Pe2r
b2Eoo0ZMv2ksmSrPdARD45+ak4lYKzyqwqwod9kJDNTusEWNc47r/+ijp6Dg
4stXoJ+qpmAVCgImPnBImDZJcddRBnYpo95+1vjHW9URooKxI706iVmLrw4t
/y+lZSr3BcFdmzwKQAjR5G5EC+EyieTo8eWZMP6wPsV9ja4zEo9eDDfmfsc+
QPFGap028xPdSM1scxRP35of587Q/79BF5qjQJUX4gicqZBo7VD4HceXvGb2
55YQ8JRXgk4bIshJiH9l7Ntb32yjh5I+51nPEWqDtGhQBW6iXQRYItkhDDk7
2mZUmS5ZflSmHb+yKfneEi6fNheC8NdDpZzvrB7cwy3EKB8mHLuIpjRNAEw5
Au+EnG2cV5dhoj3BddDOaz4e2XLUQTaFjQQhWOqV1KQ8X0uapd3WZnZd2Svd
wKYejG0CzaQu1ii7eUDZAAUwOgal7NWlJRVPxXae+OXe9c7duHh19jz/H08O
gQTmD0uOfpXH5o/YbIguLgCXrW1Q3yoUqKPiRdL3jxJQ9xA5SHK9MzzmVAS5
WmVd+DmYNQ434nyLEULN3nJCL2tzyC+7utCckYLLGp2//XzoBBL9kXdncfGv
dVtTg1VRYaWYny5M4R3h+8Lu0PMszL2OO5C6uxbSfA0VQb2OFcYBQIOVENzt
gmFDn3+2lknqPRF6faK2+0/bzUdZfGQ+E1U9PJa49SO3Xtv7e6z4DvYxWDVO
tn5Y9TToDNFFJ39/TDX4cO/Nu15bBjHcYrJbjc5QhsIU16ws5YzgbcHw2ifm
bYrRVdy786RVWD1cBRJ8Ql53l4yef3mY9y++5gUcUwdAEtqsM4jKw0n5l2av
k7dWPet/C8zydyE8OGyATfiwimK+nu+qYhu1Js0H4uYrlJIauLw5jXrmaoBC
MEjuvffoayccdnnlxv+pNWhlzu7aqrlppA7Q2mVtLkZTgTKk6S6YGcWIRAv1
/ZlsNm8KmH9Yil8HKfmP+NcTtpB26I7XaEMN5Ya+W2HK4vZNqCskT5Cp9tb3
QxEoNNvDfRfgd2Q/vAFy0Yqvlj6LVBHjv6TOwc+Mrn48ABJonuZKIdGo09uV
KIsid7yh1HmQerAL3dB5n3Ng+FCn9XTjDWSSEdMs/N/HVjhLKX2e+kRw3CJm
/IMVyBMeHaNqYSRk/UMNt67vDOzRlIipTCVefAlz/gfHYUR0/Xc4FJN/ESCK
WsZWXuOIAP1ksC3bbMHWlH8mem+zX5WHEjBHWabjSbnJPdwComZMK3tqlOf2
SdNA0ZNTGtZv7CYYZbkr64q8U5DD69YYlFgxo7XKulZMmeJrreeF/8M1yhqA
EIISzLOnuWRyYQvEM2gO+ueZ/4ckyuJZxm+wiuZNulYy1ZFmjmT0WrkhljNj
hbalHENgaaYX0V+EQ5fBZ3aWiQgZfBtAeVfgJVUIAsIxVOpxQ5EShcYly2n0
s9WfLczSiFoSwFjKwPWQuP9YG5/sMrJJFKfLxMDlnuZuvrOjdES2RfeX+aTH
KSV2bs0JYbp19LnvHa+lKSp+JFldJmkRHcBr4/u2JTGc5VQ9Rx0lCuysX3un
f8hhgSB74+CafdNSa5J3rmqaQhLiOD2rCiBNHG3JHFRfYvTLYSOUMCmWU5Gi
R8y9g2M2wT73VKcaQr1RmBvfCKkfDieCDWy9neeBHEVGVm3HkaYPwol1P8tF
MkvLlNuTqc6OJoF43qu9O4s1D1rQuTJO6rKs7+3KiajxJFdoJ2Wdp/TyxR38
Yh/yIwwpcsm7LHQFS0Df/tsALV8vivXFLi3pEVRiUWaOES/ieCzSu4zlbABh
Nx5yxWKQealgTuzXlHkgbX4qhlFw8A78ocUm4NwrBAe6LtTHnO3DtA+6mhKJ
wFOEbeVuwEXgYvauUhkJwP23Bi+pVI7n0Q0hVQ7VCwKA+NQUOfnofBbOXvEv
bDqDL9lWd4Iy7pZIdOckv0tm67mXcOJEmiqL3mPcgYHoDy3gkE1+7qB77/Q+
QFA43orTMxrq8sBoE2Fhvot+K1UBikjrv2Bl25UnlGJ2vvbODlrJ99zGUfqM
doyLq/dLcizNyXahAZGXADPkEAT9rLd4dhEgjypEMJJGmo3rfRBQ/2APPllb
J/+vNUR8pM/Lp7jPv7DJ72j6EhS4FxunB//Jg7l2K6feEL/0KKUHo3hqDLJa
olVnnjvom2jsjkw+1g6Dd+MLjlDL5mPUJ0v6D6BpkBDqgZAMrvvzftLGMEzg
Me2Yry2z0DF+X/n2Eup4iLUSSeFcqWm1dR127zn99cpfX/2TGyxL/FTaPHH7
ziHnNgcefTOjKScPwGRxpPoh3Ex0cGuuNH/+47U1MpHFPJsvrEsnSmRwCm6N
safo+NG5phGC5I/+bXqB21ZUtYIeDb1zdbebVz9ADHO2VtySkp0s9XW2NRoS
lHHrErDUcSEB1A89znHJPga4q+xAJCu0U/E1KtRa8bbD6JugkspuYJ7GIbC+
jEz5r98vKMpUg9MoNmTy5qbHIt71ViOmmkImqtl73f2v6LnZl6ScrjDgfJSh
QyVx/1fnm9cVnGXSq9Vx9XLZYfXAa/AK9eMsVeF2E7LxRJv4j/aSmqlUe6gG
HWjrDfVDy3+zgYsRBz+1q7+7YwuBSvEEKqV0kxwRpSrlhQEG3M4E2I+YYZQA
oHIXICmIipa9py1Q4lZiouTy8lCX8yw5fKkCBa3leZjiXbf9XWBpvY2rsijP
V7FmwQc5m8VcsYy0HUxAzbCZg7C+JtFr7zMqrP3zAOctnRCdLaefnnPwe+dZ
jpwi7yAOKCQXpyDUdpZ68SQwhvtkrTtD0d1p1HkmfLqeloeCAIsz4LS3+4Zt
vxh46JjCnqlTkdZ7HLcOQ+ySmL8wIExluVnA+fqVLHhNcz84x/zvsAhDEjdN
kYL9WTDYCFEPh6+x84SSuMr8VI5HjPU2u/zLn0gZLdV/PJe7oRdS/t5B6HH0
9XV7mP+ZEX368s+byktJUfAjITAI30Y2tX59QcEirayS0hqbqSqXZBbauMR6
qG/iK/zhSAipHENuAHM2SmI+D+T7kohdKS5JsbpihTgdrELl+BS+QPWdSzKJ
CrQ2YaNBMw3BRrMwhfP33whpBDBz7IpXe8zRHYcxE1Va1IG0zekNgL2Ywk8F
52eGaJfvbixT6hYZLB9GfTLl0YIoev+7MrZb58az+MR8R1E7T/ceb87ywt2w
M4k9di+m6rdLfLklGhI+Q0raTnB+d6z4tukpwzU4kVmGua7vsYFZ5yvEyFog
FWr7Nyb1x9bEzOCGasfvgsKxUsGVDX6j/hLijacZ3BQn4HA+CF1DE8iA/eIv
ovvHc9a8qdJP/utk3s9JgEOuseiGwADhkYHdz/gu0YsqMZph8WITBb4CfysW
sPoM7yRPjgbVIrrUZhB+yajcTUxIBuEv74I5Lf8DqHhjIh27flXEmwbP45C+
rXhXM9eo8ECrfmIj7tD9bbUgB+xCD6ObB+/NAwnQXfvdkh7xJfbce0cIfvCu
yfqQhB6RKG2SHyO+sljVt/qFtUXU7WPvmzHvcVeVCOuvkhnySbbk/k6D5/DP
8jJFm2oShL9j5k6Lz/3haspW65bt6mGZRY4lUlS44Ir3M92oqXvgtyvGpT8W
nB+PeaUPRLesqVF7loOz0O4uTAtKYyO2qD+0AhxT6lGQYEB6KN0fWHvHDOuP
pYRD1d9/c+6BaDXbdH6jKFkuTYOj+fBl7b0d0lek9h3XGFJw8yoBjziSQZzy
64FMe849ecQCIgA/Fj316dr/2rvB2b3TxrpvTU+tt6aKB1/hv/wkcBXWtxKc
ptZANwGhIT3Axacjy819AxB+/4pmFYH5QyVxNKPHsYZwi9a3tLA8etAw9H8C
M+VYyg340pkWC1cKip7ixfWclP5M9Yisku3jTPmS61QxZlYIDU9GoXFNgxKW
BUffhV64NrB9O2MVAwtph0CWODjx3i7qoyvQhdNtO8lp/pWJeZwH53m3RZeu
kPFZLgljXdc75nLl0XeIJKakomXeeBTGZ9tVss1T/kHjnOKyOWTXYsmyAJp6
zBUNu5vJcoFupHJ2AAiHCiq3+U28+34txkdA9Gf2Bne6qMITNQ/hlSvTVaNl
fVnlqSHCt/KbzjEvBjk/wS/7i9s+8fkQmytH07GA/mWYGTOOpwF5VQr/Gi4I
BJYzaevJWOqpSwVX/REnv4kwgYRPtzMZKmJkivRqFULRLN32cgoKcf2Znu1g
npF13/cHCrzy7P/JCAXFI6DLFwQTJehm57tBBAwesx0TQik6P7lNhRH0pxzH
6qH22WlzL15Tm3dHSQJbPCDSin59jFeZGRxiFGumpOrjE2a8zSZB3CxqiSCG
dcq7ys1LqhrZ+Oz2MF4I5mK5uTq8OaTcqAAIs+MMfXHJmMrX+KwFmYpgEfCc
aVylNP/ZKY8zxFPI4LDvNOwYAwHd4FixTH/0JqLCbdZVY8Z2y2HgJLQHQqtl
j1o6/L8o11O/Qb+gVXDOfg7AcE01wjvCaWtFJagmxCu9ev/kwMy9U29omRC9
hy6gePF4I+RLVoWsVdrvxxlM2HbF5oil1R7evBbRxsNwwx3lamU5Fqq5ksN9
Y3kvLylqdoqcH/lDk4m82aOWrBj+K+OFhJURqwrBFzzs/mOvhVdrSIqyhuSf
i45Yc0gcNw17FrRxd+adiRY7QVHKSi+nV6ejjbb5az5HoLOZqqUeWP2+v+0B
d3oZ+hmAEfprG/UogmJ+GXaQRqd0NdG7NUGzgw70VYJYdr8IinNEJsF0UNWT
0mixan1mieMucPGYuQTlVMMkzOitySR+H6bL9aibJAoEl5AHX38kL7dycniE
rkzCr4rBHs+sI477p/pckv3tgUiO/Pt1kvM3U54bxmRWWU/vPBzQdq5szdQv
ilcq01hhtA7I3v9WFiwLcGZ2ofte9Kido7XQ6YbqI7p/2ye9Z1B3ok5gdIqS
tiHH4A1k0BV/1QW2qGtFuZotxS+i5x7xYQExzGR4LfXXkrFO1is54uH3f0p8
oJusczHDKFPhPhuHAX+Lp508P6TJ2v9on4rTFW5Np++cGHRpfUFwVTIpstIg
as9pWoAl93AzYRWCm9yioFHMN04Vunqk5TVQDMsaLS3MaOVwrhnFBvyjNkAm
uJoFz8dXluiHYDqaGI8PlXWsmuxO06sAmivF0h7THGNCfPGCg4MsQejx/vKr
Orw6wgYu8r7A+5O7kqINZOCQV6KWw9kAF3ib7tJeVGQwvobT2+Rj/k9e10fq
ka25k95VbOgGr/6gsdwfqtKm0h39xayvHJ7HKdMvH0HKic5V9sHmz5+H8tBj
i1jWZ2jW9tuQR0Cn2bFC1G/qBpQs2cmd2K78dJoAWivFJMX/oc5ISSfzuTTy
2DxQhj0HdDGgENzzE2nuRyiqld4iRgyqK+7xezdO4WbWllVSpei+1VNHDz2e
lhXaMaEDiBiin1Q8ONpKGuUU3AHMNEliM9FiYsnRakPDFlaGExO6P2rwXmNT
yK1Cp1gvadLbzMRfx5zyY6MzXaF6pEtB+nDzMcO7JERb/gGEUdNME552jLBJ
qslk/P5FJn+jpssjvtYstuScgE806PHjorjNB+mZxBePNvfTqROPPO70m1hp
vza9ywGTl1VALKaG8NTGapazJxLAQP8tRMMeHKs57idPptn8pOYmlgqeO6oM
aZ2hIxKAGsfnZMACrvqoyxL820eFMFHXkQnXl+mmG2GDeb+98xTPUYEEz7i7
5nscdXpcaNny+hx9ViaZyL8D2YLV3NopuVyuNsjscJwl+HiBhD3rnAHdkdDH
hsIPx53lHWynoqGSfokFZ6Y0JUeGM76bdgi5EgUKO5edbKxQweYXdqX/VirJ
8CqgytElUforiW78J/x5rlIf3zCnyyB9VKqYMNV6QR7WRZM4ZUygJVxhxe2W
264iXMlwE1D4Oo+dsjms4cI4EvAYam6fW4z/vcUGhzdJ9Ymi7oUw+/D0mrS/
UHD1wCCD+i9d+zOzEs+QMqfTVtgBvq1pQ+IUV6xjhZj17DST7/QztMATLfS8
qbLnE/dGyOzgEXbxhak7OCGvE16nhrCA7Ixh5pFjfFEKN29a2PtWu/ffz8D0
EMVYUe3EbpMzkU2jqXFtP4BB07WidHHne5uiLR9sM/W47tZBeK41QC33B78A
D6V7qrGwqUmJezti8oG49Pyh+sU69GShCRi6owvcmOs1B5x2ZGrtp5nKB8TP
hnZ/b+lfTp33QG/IrDX84VvedczSyWxSR7aAO21V9OtAF0Z/Vy/j6xIULC/x
JsRGDBc6Xm9Y5JSnSVcAL+9VRti6wwvXU99xg4H/4hAAEW5peNrqf95O3g+4
Vn1fcim0QvIEHIY9N6gyFDnBaYHEPctHyhM5faBQqGZsIRP09S6go+APNQ+5
hwxE1oP2XsAZKk7teK5lHxLS5AweIFzzKk9Ud+98OjmMpFvJD2QQurFZeVkK
C1CrN7JDTKN9WBWlDoxgsjIh6e71TscFV3f8DrHJmK+W95pZWAvUtkCN5q3Q
VhsFqrp8HUy3jEv8+03QR9E3CQnPdkmdqv8DK1nOeXLMULWiesxRdSgSoO+U
tk7GV/x+pnWW268JZy6E5dZkxYry6JFsD3FYdwCypBDdKoSRsaj5IJLr5idT
IzBmYp2Za2YggLG3SnjyJ1WHSXk8Xg9+d48/xmIdxBwx1MfrTjL19XCR9ihn
+SmvAnWoiEiJYSd3a1xsGPNypNoLEyeuMyxCfA+dx2gkgbMoPoHHg5MrKtc+
TSUn5Rs5pG4VmefVw3VZJDfAakN1ZAwF5brtpqV6BleC/xhRoUT010OcVLUh
Oql31Zni1j/3dzAzxrMEthY6ZQCvaNS5p1IMwkf71V1sA8tR+MvakeKX4bhx
4jD2RNvsG+XIQ4uKv6ilJkoMdDiBi4f/LUKYkBzB1ZTNb269PEgN1G06ikBl
eS4Pf86EwlNQOUNRNj9NnQ4zM5Q9Zjo1QySv0f0ZYkAsVGuqijT+WK5lPwbb
o9izsIHUZSGagt+6cnVgv0aUG85/bpyT1j7uFlQj3cvKzcdIlCpqLF1fWDBL
PRctZdXlLIu46OMs07G7M9Z4usU+lnooSojmgLYL8KUy/lk+wJaJo26u60e7
i8L/x5JpsPx261uuDLzS/5+XKzOx9KUPZ3D7FoG+37oHmUW3AftWqAXE0tkn
JGBtwxIPHHgOOVchT8vX5DKI6KGa8fAzvLcPflI2aLaM3kSrN+Tkudw/ooM8
m6RlXfPNMu9rFx+XvIeOCO5iT6yMSTdCFv48BUcSgJCf6XSIZq06NzV16h08
mkBL8ZWKXLilKpbxIGFVbS0R1DmOSUYAr9gxMvdMU/GYo/H9gKnAPGMLAq/s
LRht+IYWqRYK2FKbykNDX6wbLroYc4ouP+LlsoK8wcdIGM+xTRpRKVez+ZFm
NUfs8kTPU13FX9Z5ExcvYI0EMFkhB+9Altatcn4bvUy4D0+wn8Efde2YPiSs
F56/E90q/Ol5w3P73oq14RfQdYROPrn2v+jw5q1v9k24rZYLRNSH8OVqtHQ7
45ZgXZnTqbebw97nNPYIZdxMsc/1Ok75qfvo+l7qMjW/JBoul6NWxJMbYIWB
AknRunlsm+XmK2lrv08Apspk2saPQFC9zNqNv0zD2HsI2I6y6xa5VORxZiZz
hFrRz+d9rqTLkysEf9veL9uJscc9ry0uyZmtl8EdhRmVRGFZozB4Vi1wUBgg
UPyFUv0gMkCTcdm6U2O4NKBRGal0PBQgz6Tif7X5lrkWjqaLmKjpr3laeALO
AZwYc2aAv8Ic1XLJeUps7tbc5eraZkKEcE3azZy6nwgN/oGaTJ2DWF/NUr1z
PMN6Y1MlnOdfKNI7zrMORGGMRGZqW6xVSzslgpB9Dx0xnLRRyxDN6CwOml6H
shrJFX6Rz8fNopBTiXQkpLHbzHiOihdccyYRqe0yOt7x88NJKFFVgsNQ2MXx
JZG2aQy1ayB2C0hQrT6IOGhqsZfx/MKpgO8MVZO6dOBQZewPLdd6NcvuaVoj
ubr75CJ95abteW5+9QsTdHgEZjbVPPCZ9yLki3V+gPQdtV/iKtcvjV+kZKlL
OkqRjFKGi2gI9zsQ/WiPsRUexyH6zVo4HaTWKqwrI8vTbEt5py513ebRC3eb
1f0k6Tkne+73LEHxiV8Keg6h4bsuv5nBbpiR0Q6k7/lgnnfdiF/WY8g0W1p6
B+um6OMwIgVkUicD9InHNjLa1jFKriVn5pTCOCKLRg59qFYLNsQVV9lzVUCS
A56Lrh+pqSRAEDcOquV1OvHj2KQllxXxNgwCg0EphWCOtJFgPAST+Iv3nR+z
HObFfNVfK2v2uQovvpBDP2Korw4fzFO2cIpIzlGmiEofecOzG8JpnQPDpTUt
DN2sja3xk0pMJjlxKhoGS+RtAROILOokQmiM9C73qSqlQ9UmykBF6SzXLw0B
GfXjz1fswCabUx5XTxVobhaw3Z+brfMvEJlvsBth8GBKAXz6U6c1vkYmkeMQ
7pvXAsPiIlhBaBieTe6SS071OSlxAmzbFehp/HXPipUaXcl4W9d8c6rM0uN9
6p4ZjV1I0tW9mYcOuE5pP8jv3zXUF/enwFwl/I8RyEICNKDBYwsZ2MYnAs0v
oqww41T0Y4DZE9nobt7C/qX2AJjGwOKuKuAJO8J5hxL6iInaJicAcH7NSFh9
IpI8j4urwTXfSLJIeQbUtat0JIj59nKs37bJL5FBBLUrrjQVKUsb/uFbYZh1
5AmPeBm09qGiI7mJAyy05XV6iD4FsrL4vTBwRkQBnzjkomHkTlZhiqQQLU5g
20Yv2c4EOX12/QyyNZ88AqniRTUZWb/vBeXCThhfs1Et67bA/nZh0zjT+sW7
FQwZzjUTuNTRFdVOx+FJXPIf0rsj7Dzgk8w/q171rUrSxd2opGQk411/Y+n7
nsP3bqOMnYyfS9ocwkOTzmfUWhr9CHtA3MQk1eyJtVDz7t2qAGLSR8jKwCCv
ltQGS3W/AyVW0wSUoiRzY8fxhmnHZdBGoZWAQAkWuyz49ikFqstaEJXzJLV6
tz6i5YGlaRolnKZYLxriHpYf1qC1FbFM7n+qyC/826hx0h7rQdHxRNKKSz8T
9A2tYNgq0sODQiokrVWd7Cgf+TovFdgKM7q6IYBQNj03KxieyYbQrFy462IZ
iDV3M8fNphORbgjml3lVdtQ+tA7b0ndxUuvP3wE5A1/Oh4vRdDv1vH2bzVnV
z6GTkyeqoVYgWvQhyVkJdRUUey9pyXyAA0Dh5voG7nbd7G6ZSE5ZB50a+3mM
apPHvGzawC0rrtF/mFded7BrW3uf9hSoj/b9dMumZi5nh+pfZC6JJKzEkIsn
Feb0ZXRSqJ2S2UuEIeNhtNwsw9AipaXy0Qlyjz/VPFE8448C46HHc/6hk6z5
j6x/lvu4Cz1R+42hK10V2tmLup7lnjZwpwsdE5x1Pptd39U2ofdjsiJTo9dE
knZa1EbHn1z6OcMh3R/dBeLhVX/kg9Y0ybcFR4pqREl+LmSqs8XShdA5QzUi
ucT+dNBJNuW782qbER5sUEKNtalmk5E4q8Z4ARGvP8q2gHz9P39P3mrUb0lI
LQZ3Iuc+/mgTyWMK/D5y+JZeC9ijpwPZxDgjws7phzcX5FBMJes/PnzVXUox
hh8V2b+9dcIL+7fUY/0+QcJ0dj9Iekt0CFk07pYnG8H9MsYfNU6PBIOKaM1A
DRrmRcCf9fl16KTrtbnqXRU8xu9kVU+0+D+DH97rKIIt5mAb05Z68cQifrYR
Lsisn8pfLYKmw6ucHf9ZxumS6IU9TLEIe7Pl9Iid/Xu+xHTGFK/F0Xj7Lmn1
vUlyfKHTpva47L8xc7ccm1TrAmYfq92Nmafk6kcJM5nZWmYjgLRC6FzQ+XZ7
gtnmd5ml2wnUxPhgj36kxx5dsH4mniIs6qnPmGJjzDHSE5KBolWapPE9V5jg
kEC3Pst3bO47hkmpCXxyPrl/woGqC+DQXvffNDiNCbnUACg3MHhs7UxhI9J4
8NTjIablDslYNHhvBFloT5Eq0jZ6Jk/MkBSYgHQDb1bwMCGZymkpo8kKIEKL
8rseOmhhFo4Pz1seg52AZCvEorOzxrJjng0YUyPGspNCBwGq0FPqPFs3wBO8
iYsd+seRuOOu6HrXJQMcAPR0ub4JEpcgtzgU+yKzr6E3TIFGYouoxMlxcM9X
s77DE7vw7qM40weG6IKHeQ/6jgj0/P6VxcWhCvlSsT1HMHDQcE1KXx8H6Xug
v2QcqtcTSPVV46bPfRT/RJHr7HGI1gK0LpAWtiImd8UQ3uJgYpqBk6x6boBn
V1zYPduWYUDLgiViVMdLQ8R5vldwnQ58dL7tHRK8SWVWnJyDtsJgD4VbA0ro
XePGj6VfwaujDKcIptjZ4aRsBKVKRe4a5jCg9HGP1CfuQG4xpS0QrfNRZ0uF
okoId/htRIAFZUmCMPBRbKX1nskoi/NGytkp3PFSWUHWuIaQkY1BJoJM8uYD
FEb7QYtYHZ0NLJhOa2BizOfHxf5XXOYsNLnwKOcsFKj5N+qUN3rY7ErBxWJv
y+hVK67t87B67ySbrIUbZHZVnKRZz7V5AlXb6zPxM/f/SnV4WGAc2W3SnlQ/
tRO29eFNTv1tfR3LF8heq9ZhDrqFy7j7I23cWnToHjqVhdui1ab+nV0xGC5E
Eg0XMaOFJHehuvQJSX7mBURgQtFarHChK/XtQ9xj+EwQuywHHgwRfj1QFI3c
8nyVEcks+QEEMvv+kzs0VooknKv10pOtFni9tliRdYcDKJm+1nO0oCZBToA4
wQawWEDUvrkmitJ/zHt7jkzFSCOe+AIIs6HTEhHL3sPPznQrt4Xbl6T+x38R
WPYfHVT5oT2SU6icYLP5oBCnlrd7x1jMBvDDEtzdSYhJ4PdIARXhU3ZOqCZu
L7NBLjAZR4Xb3N1BJJIENUJWlc6eZf99cgZRQZViy5TYJDdz3+b1cAsTYj5f
b7lbwsIQKjHSZa1BPWBAckY5P957VXjOKD9aqdNc9Z6MQf7nAzLh02A5kqsz
xxgtHf9p9T2eZ6Ch8XhlHPoA8trPCgoyKXgaFGrMPXhBqYj18+I8300IkKZz
6YOqmrypyqNdllkLdJBNLuTqUzbk4ErPC3u7Eobq+f/R9UTs1WAL5Wu/KmyG
LSEbhpzKua0irIFDLpryOqADF7BTUt8fxFXkB6qSB84KhaJFdolw1Tvljeda
b8vLFoK6kQ+myeN3Ab2jJIulvFRBCPp6C8tOA4R7wTPCLcv8pro344DFL4AA
E7BrOIi4OxO2W6zZJNacYUqObUFjzA6f9x41K0sYCvTevfnt0grQPoLXmTHt
UeVeAXEqsF1FmV+XTXalwF3jQJa9Gb5wnoOQlYVJtUV4lczl6xkC6q2LgV9A
5XPHInJCKFZJ4W6ooz3CZux1368H8l9D5pmWSiN3w6mDmpDG7wGwk5ai217Z
3X3oSY6XLzlaRMijn0nlLs2HY6FbDyC5U6pE1h8JKOo3gk464iEclvtVG/VO
KDtKD4GJyaw3UM0982dBtmMLzAeuD3poojM+ZZD13Y+fwWyUxJc2P7Uv8GUG
tSBVCsy/7ykdlrVvJtbGFA6xzXs1VrB/gB420kIHAsG5SrVaxF+tx6lay//M
o66wXVg2pUEc3oZyf/Bz0LdxAFs59b+A9xOXuRgIaC9+MkMRJyvZnxx1w25K
i5G46e9bnDsXf/hA40/p5pnQRQiKFu33J4ojHpXhOHTWlQxgu5ASm25B1Tzm
8p8PFHwOSuHqpBjtNJofplGo1c5CNiPapM6G8SFwBb23Qjpw7cBfdSemhf38
bfVayMeF9hostMJZmfqKPWBtpJa6IP2krCl997wHeOKB1jJDYU8iyDlH4w+a
XPI+ViApYGREGVS1yTthbuUMqn7s72kB9vLrrPxDuzvidto1CfBGLdIVy3iv
EkqW6r4Mi3q8nSFKOAXuE8qm9NqfiDXt6TiEgNJDvsX6MdZp+LMbOQ0CyHl0
diz3AbCtgNVffmUPoj4Fo1H8q7de5Xf5o1+s3BzS7wyY7ATZx3cjVY3sNZMB
uifVukLxt/hXnoq/veffhfWyMJ1C8EgcmRA7nn1NM/3H28JkTr9WYR0tBK7w
xFUkziphrVyRu0+4I1AFSVR79RDIqZe5Z+sEtaq5VDIzNLxDzhkG5Pm4yNME
7za3r4YWYquv/Fq2gibNQb0JOPRr8sb8P/jSzDcxForiUeiHYzO8SiI5p6Wg
3kkNl0GYGCiqLo/yaFugqS7tipqcHnB7FAvqaWxO9wWq1xD8VZmV63jxVqs8
IqUxcP294D5B9i8POdOtYe3HdjiPwrwz84GaQ9/hNoe8+828FTduu6holRDR
HjWkEGO4Xq2uVLmfB0VfjqoYwqdCcQaWZLuqWVwvV2X4ZIvYErPB3Pu2Ss9f
Z2ZLwKZ2GGFdcpj5FZ6phYz+gaGQ9ZvT/Ua/VEQBfqy0awOOPPfAz1zSmnGL
BSa7pN17YlqR2ASZZQsFRUY2Z8Q+K+CdYghmoRmBx/mow+WS/A1KjTYLKEfC
kRlJPTStuPhVD26prT1Iz56vHjRUCahKTkiYS6t1ETNRiEM3fa56QRcNW5b2
jrPSNSsk+ycS7oEJB8ri6NkafXZKKqDVsv+0moTkcyHOjZMfKsOZqco1Bde8
65fe2Kcd7/97Y60/OzYCzPvoIOokWmh/tkjpD53DBRwiRPa1SL4eeRioT/ql
ENsBWRwJKUjN+7sUdCD2aN2QS795pT/mJGXfdgiBohEh7I3zVXHlyFmNMzLK
waG+UoSOmOK/8SI5ohDIec+EnZ2IKXPfMNFTL/zQJrn9rwWnJxew79HFZvdf
AswQe2AO5pb7++jbJ2HX6eMYAdrsv3a4JKCnkRV7HKGeK+VXkMRFVAVfUavv
6dpts7ZsOcFhj8GSbh4Mj6o63iUUY5ek+/MGynhdHBK+CbN540PwAJ/o4uej
CBr1sZ0VtfEIm1jCQO9mf6veZwNibWP98MxNo6l5GO/PKdlFSHk0dzufGvZe
670DfY/OZ2Z/byC2zH72bf/kwLqIPySvUxooM12NWLojPE1VJM3hP9I7RMVJ
vcKNbgdTV82PF5Fg0emImje6IEuvu0t/5Bw+W8CUQhMYG7Nyeq3pNLU/W04P
hzgbH9Jn+z1Tatu5dCJMaP8CZ27an1JQcozLgcMGOEI13RKT8RaX38ATRqx7
3Wh3wMM5O3Wz35RKkWLVVJxp078WkgnDHAktB6kFn7IzOmh0uO8i0WwZaNgM
nSEGkBtqyEV4YlIfrQV9ZJT3XrPKLUhzdFJVs2bsETX8EnFgB8IWVLZYnTbC
KGhcvebbYQcSRq3r1AmoSSKi74Q5aUPnumWwjcmqr9CCdBcZaYTxOe682AEn
Drj5hw0gNR8cGsIsCw9mAT0x0aRK+LxDf4fsS+nLBGquTl8sZY9rE/H3lnvs
4Y5+ZhsPrZap2CXyknKOrgri9gjOYSGMm/mPR8jkez0jLwTCBOmtfQ6TYnTU
9XhthtDPnNm5hoPYiILBambbux/Z7IgM1HTV762oc/udO1bb6zfEUpfLA6Gg
OOGhNj96n3edzMrIvEbsQyJMdJu543NlLs5peZfHDIsI24vUFlgrC0EN2pk1
VQhZTLzCI7axyVJLm1Qo4orTG5uyZhnUxUICAD0UKKvJyuB4KtLtWMIbVmb3
Yxm4aeMiYpNP5OueQ2gba8ezUr0PfRu+I7ga+OAejctCJg+ok0tzmOddLfXO
li/yItMqoaNHfpU3ybJkn9dG/ANduDSyXwVf/N/IAnpvKkmFz687NGnsoKgp
bL9nmYsMhajdXdisKlwcVvbk+DPAaR1TGYbaOndNkPLi1udqh08sQF/9Pdyj
dJX7BWUUUQplVqhGhrKI3loTSoM+XeHprepSr/8mAPV0c6jEU5hPC0GSit1z
O6RAqam2IfvfUGU0w0Zt/NLo8jebzUQdYT1hjKuMFCJz7G+eN1QlqRtzobbE
tWcji6g8aCCnQ12UXxDg8cD5K8+ksenahuV0XWwnkDMvfTlzmVQlK8CG8n92
Iz+5iRiGcM+Oa0eT63zNiAtF99UnjAo7YPSS5cy8nfi0uM6ypucsECcciy/z
4pcLYnN8QmwfIl9GI1qA+0a/N2ciZxAiX2zMZnCZkyMis+FdHuSzJdz/BYPy
hQGmUA25wiPOsWbb9IqUEPs2L7BjHYg5IG+/PitGCKCF3mkFHv85yf5Dh0Ve
1NGYIm8+I7AZrT+nFvYTOgCUFC/SklteXF61hhT9wGWmjctlg8xD0CBg64tk
SHjOcxdVmNeamomD5MV9cAsiBj2xH5OOnaIvDTPDPkwhJkzoXWW48Hil3rSF
bvZpe3Z5MDeHwN3njpZO7KTAS4jM84g/u/hEoIJQtrYq81EIXdUS3Ui7V49X
Ok5++s+eztEfFDyFGSiJjB6azGQt3C9Y6A+FY8t/y3NIJvr8GBIdZhZ8mijF
itvlvUHCqLiunfNe48zVvIqcSVrdNphCMuFeS3BsBdVe1NjuAEQo8OHpZPW1
lo1nPyrCMx6o3p9mj/ichJnd74oKL3vl+r4qDxaixoyY7imX5sENtbpYKUxM
Gk0dGq9uVrcDL0ZDPERE28kKDv87fI99l09fTmjyiZ84lbXqwTSBatvvSVgI
VbQpJdTxkISUUEbc53a8JGFqMgpNIr+fa9Ut/biCD+N4wu7ewgziPvGYHmyW
GQPjvDc21RwkV859ZkUbvLK5kmoqTLKaOdaaZasivTq9rBcQ3OFtQ47FN9De
byU7PERwjLVPdm7JY7xfI5ovSBF7h/i549tH1Ht2T0SSqOPu/vQO/Wl7Ezld
70yW/JSpGB0SZ34dnN56PjyCAFN9wcpSIyOupcEoW9d2Uy6F78nQT39t/YD3
JGo8atN1JvhCnCvjmQtwvFy6HsHgp/vqrh52/0SxJfMCNabOl58jHI80IWP4
K7/R9gfFA3EWJGL84SKTCq3m0We/mm1jbX3PtOe+Ax665vlDaIeEt8ge3klx
4Y/OXiBjsZ0OuBHqfvLsIuAlVocCa+8ebWEu37X/lfJ1/1Z1G6zdAbdND8Rs
b/IxXTKGkXsWqIdk1eqI/vOTvjVvI6YTMnnr58k7SERxcqWD6LQ7juggfuZQ
fTsDzgEVEcMZKr/iKY7ndgkLnJXQpO/jal3/eZMO+PbjZP1toc/vAQi96/2h
SIqNGFx1AHMubGB+ukza9QcSCihuWearRRCfvpVyv4c1f3uUIf6NxX2LKq1m
YRZXVDSggeidJgOHAYwgwkvOU82ERJdbrR4o9GMC3F4Q0mOYbQ0yGt7ZqS8i
PK0Z0j6abgpKJEaAkVhc2zo+RpOEOFNaPHjw4T/AabbIGy0uCJ00lCkM9jCR
gKW92qEU+onubrIybauPRHjP0Gb49Gj6INxslriplihw0b0ERrGN217Gzxgp
uzckad9ddvOlGL6gmGcf8Awm8fR3KAT/NVQvb2h4EybTMa9kGhhXR+npPvq9
Fyp+/NTtWo1SKWUf2UfPuVtUorjHFay7XrdIsv+UlgNvd79oC+9bh6VnYFd3
yglHtTTpk91n4pRvCmZ2/CirTtty/EqqOE6tmOFv4pfYLPEIghHkS6C9TjjM
0UQUVenjJ/Z96m8HjxGQSoJ1O3qB88jKttT9aJlD4kjpg6CjA3DgaYw+aOly
VI7JjxP9goL3WO4a3bIiei/DvrIbuEzHFcBH5191PTgyI3IpAPIY9Gchparm
3FG8aGeLLczGlrG/1nhtjSBPY/C3WvyoFkyYSTW0WfVOQby+Km1JkezkpYBn
xagzCQiftFzGYqhZvgniKHn4+rM+/ogvuIK3M3594/AM4GQyAmIljwXdom3Y
7wCfHt3IXPyv5Ui0EbsW4NlH3wgeJyLOyOnGMCGxC1uRVAW0d94IMyyVUkJ6
X5i4Xm1nbefa2CBUTjUgEx2Yi77Fh9aNLoxSW5GN16QFUcNcVTgDV+/7r4w6
0jW8gZeEvr+XJELYEHwhNlq5r7ehHchqpoGWp6XuGYD9bgAd1ilz6lKzXVWq
un1vcsGeTJ44YO1YfgIrih1DjE6BI7PXCbhyqXrhkqfJqiZ8AH7YNVyd48fx
hP45OEzUMG0thAVdueSKTvXAG7JcPjVbkLVAW1zyVljcbAnvsCMdqFcasWjk
SKInY9gTUVw5fY/nCxP6t/TrCqJHr7gR+cEHaksi+NC4dkrFEyvzneMmz7qf
z5UUWBK6pX3Rs9U2UT4xERVpUX1nK6r9hn8lIu5EagEl8ttu09hIMGRngZCI
02X82xdSzqFo7lS/+DZRZ3N3Gfi1HZzcZOlq24o0APAGZ0gnt6+knUiPsZ0z
1wGMV2vjyUs2yRCcpNVCIdoNpuBSfh+Y9FDfIuIrABPhDWjYOjUzDbV4wZ5t
tK46Us5Ons1ycVuByGaVm8RRcsKM/T2IsXqSl/TyWtBMkb9jtyKBc8bJTc89
PQ6r6dJeXeX3cF5vtZnRUQV40stPnFV0nIhhdDeVfIoYr2/m7MaIKJYRm+L8
jLaptE2f4PIlyQ2a81Guir0VWxLP4p79s6ifreWoceedZEBusaWhahn4IzLl
PT2tmNPUFStP/GA0QMprdhMPHEmAhlvgdD8PTntaXy/2cltvVuHX0okEXZIo
/8mzgvIH73c3KrJceJemaQgUEmEBQQHVjaMCR9LAlxroUjUaWUv1EFrp1yTq
1Cpf4GjZ8rODTAeNh0ZC//Z3/aLZVIRLq0g6nnVnOzzq16zz2QZlfctuhSOg
xQ6A3qBiD9acZoReIFbY4riI+O2HvhHHbGK8tvItq9vgWFzedDU+GwPkOXJb
runa+zz3NWr5mYkfuyDwsj4UR3CNMWHXMNuHfd22L8UOsfhKvKJZ3GknPPlO
+nUjb5/gRlSusMYyGPdyT/e3GGGiW9/WMkm8kgvataoWv6fh/iXq2cx1TZ7M
ILoMeFVI7XyWtLitsjbOEkDUGBZiaJOECHJQin96GzI14qomfsCoARyHJqvR
oCtSUAWtBgTISdsSBheL8WEd01EhDCVYlg+xf4KLIyWbGIy/n6DXDcjKNwr/
dNYk0loE6vuGxyQ1tYbtpMuoeNG7F+1AfIsaC4PdquznfGC7beVNQ68CRpX1
bx9WXk6+BGfca+dWAmEpmp2A1ajn2PAfy9iwYBR610WY4FK1ZEILG3ZM05jC
WuI9v0i6Ra4dEpDMV9EgEL3e5jmhA3eMXXqClKMGuHbila+RBWBOu9SATMQ2
eJgw3SbtjKbrpFn4Fza3sxR3fIJ3IaH/xazvFJGbBHd2Y/gDAiXXJTZWpwru
7Fe0HREfjTxKHHKjjb0odcaHIwFAnXDDybuZcIaz50zYASCfM56f+7QQt5gH
lLhQkyYn7lOV+xkNykA38yA+9lQe6KrnU5CmDsX6zpqLZH4CpOFaYsO/PQ4V
fz1wua714Bss+bHrM+FRUQIEmV296qaPcZccXUlHSwuseyjArEvMp4TDQoc8
hDf4gs+dbE1qVul3I3XdfTdmxirR94DaKMQyiJaWJj2uTiJIebE835E5RR4p
Ceoz+LSv0yHej17s3e1cfq5FgyZjiY1BOPwUCQht5CcYh14Q/XPcIRHmkOQ+
Tk623JcVVWjJCflvBaucjT/IJ3WewXC5UhOs6WKe7x42L/hPVaTUec5UtO8N
FeCm05kT8eIkae5YGf8I4kaWi2YTQikvX7kWoD6Bwg4q9uHeGT/EsmPff4TH
i3RJcLHtsIl7jA3jtW3/IyWHKY+xysHf4rdRhmctJBOSpeq35b+6wf416S0i
MuYH6d48HXDL7mJBPgGvk9okri8KtfxNQeX/jJrPU7abg/eTF6VG9tLCgUha
ZpqjOVauGdPj2u/PHJ3P5HRUM7U7HX4LhFxNrWR6j8/Nc+FdYVQDRxZT/Lsr
mlO4T9iT+ACBKc7YbnSLp7jYxdgm8sTX/MufWgxBXH+8y1VweYmht0rDwLCE
YGdEOfS0UaNrRjlaEf+yYHyPTGwq50PMa62WT0CkHNkgJ9o6ALKfWmRtCeJn
lsijH8FKdminsRQ/K+XRklajC9wjfafFoeDzierZEBJIVMfJlHtlktaA4btJ
ED61RjrB2Y+nDesIdwo3+5R8501O3F/BO6ubWaXy39JkUTDM9s0PZyn+7EN4
HYaqNrZEBH/gq8a3kYe2jx2fG76WAlnP7AtMI9guBn9qwz/8xQ+fgXOILROC
FJZcNHOM5GjxvJRkEzDyiEzIVtRPOAWJX1qirWXN1ql8tHjr0+He1S0eS1UP
SBvosx97NEVog8t5oq8HQCI80abLqNIuUHZ4Jvfc+inu0ba5fZofNc1L9I61
tD/Ul4XbzKk7Msp8eCPYDj0rpO4lBgZRLGuT0eReU+etC6xsUzKvmKht8HQL
Du/TkGKh23VzsF/8UUUYQgmxsXq/IZyL0/pWQudol/3t7plprrCf9B+s+pcf
g1mWhXDgig6SKoLhEIPVPuxkfaSsBB2FsM1++zzVl9tajbcOnlcHqGQ6ci0y
7TpxT/juDLTAiQL5mQpZSAZh8HIz9G9orraacCrNJ5uEA3NW7p5fCUBzZvwr
CiqAf6L2qMHBn+e00ReLD+m3Pm/G95idIHOWslJahynJqElh6rCPZE84adJ6
mlvr7bi/FSBK4k3G+1MdzGRfQEjwFMyIOzHB+Xae8bZLx9+P8086WJKRRH36
+n0oGLlccIjFNqxdwvZ09RLUJnBgM+qUPj0u2EfttFW3GG62Vr9CKRd0cAok
Tqq5PK+SCaxYvdEM4suGZCQhYO6oVjijKZR+V9iDnx3j4yyo+NVU3O3gbXLS
jAfCH9RPQc/SemtNdAPnlzA7xkf4JRCygYW0UAolBC5kUWFMtGs4shcvfAUu
yfqhlJJg5KX3Z0+5cs1f+z4vIizunF2MvmuE/XfUl8so4lh3tFCHMUsmnpWy
GXmk0x68oy+InEIsv3u1aCjdo560oNWK/gV1YOudwgEQvCMEB8+xoYOLZbxL
fpr+M5UvtXYyjVSPXAQIMzrzdol3NQ9TcPBs5BVkmStlWNhYDiOtCjTFz3aw
DhSIvcBvj7SusyQaPVBEcI6IOPJQBmwmZ1wgZR14ERwz4Ut4vS/RxcCwjLxl
+QYtoSr7VPWNmzIm3HznRBFDBjQA09qt//oBSV57h8U+bgPNmx/BrcV36wuD
0KvqgR7b7Q3JhYrrXOhCAYqnbV8kXp8dbqBzcAY0RmweQPtXFUixQbKj+dnQ
hJ47n5rKvVeFLrIkoGPus+tkvQMRDYxKgdX8E8jdvQ/M3YW/18dYnoCgWCjk
hpFNgiOP/kGhgu58Om8pq5YvFoIaEM4vMoOEPF9/lAa7B4j98OLewSi8QOCj
D4Ok9YTmsdrzDvhsgqK+ZdYxD9iSDgP43VUzM/s3rJNq22TcAP+zFuP6UoMk
Gz5HApY0/2870QWoz0wsc7c/RAwzp7FtkVpW4Pemix4G9b6ArX3pobcvzIOv
3Age/9JU6kgVqZEyt1KgnPobZnOf9/6OHu1tl7gPDfFWny+VDRKa/pOvWBnd
3JWtw4I8AoaREpTCZiYg2rtLxeWHfHlb7eykE6WPPATFvibQi0NI9tuQwaA8
Mr4U/r5wQMIKlznet4wcnOvT9GoLjFTtXu41Ym4GR80rmaMLMSsqqApEWKOl
hvvPQwr78PygHKy0iOuBZ+jR3+9VRMXj1JmkcIi4rspC+ns9FXM8IIPUt/yp
NAN/fJqot/8RYunrFFbRkD0sUOlkxQgFCoFz/nwsgq2isDy57ioX/HpGmIS1
BGGN6qVmaU9UX1XfWjIhowOPT08PI26jB6bLmGzMOV9ptsIj0q/jxRW78Wt/
6Kj9HV9nys+/mtegE27HS72viuQq5nVR/ZHSVa6/rE8xl52pj3fEdcIQD0LX
vDL0tQKG1xUsj/pqWEFfRsacVqWm/SyBt9c2JpIfhlTiae7C++eGzvCjTVm/
r+vZyT1NJYWJsqhYvwCEBEMa25+0LS+zSP76fOXTB0CHRXWylPo71V1eom2x
0D2dqd3gpF6TLuriUi9avcfmJoK1h+1NHMVdv3QVx5gnxnOAMBGRAF0C1gvj
68xBomP/m6L6saxQO781VWY1GiQzZCM7eH5n4j4s6lHJheNtpB6t0bIa+Cr0
0cKhR2yuYp68FXfOE1AK5garyK1e15ansZUJUczF/U8xZvYl4wAXimVu7Yel
HwTUOBWRGUkcOsoiiPgTo2WGpPuP2IwkM8IAnc49oLajM1UUCE922Fx8qf6F
65CDRwaPBblfSuxzTH4fbfzXwc5WdP6NN/X41s2uJcraoVjoZJeMfTXwXDRd
pZHDIq3rYLIGgBSuFS/P0TK5/Ml1w/wjcADm94MtvuZgCIBT/4mH7QTM4RGW
Qb8Yjt83hGJBnXGy90CXwSVXibTQyp8WQud3T2ju+w97iH6RPkSQlxruLZtB
MLd+P2cCYUk3h9eb+TUY0Okm4un2aFJ8Av+2HjXk/qnZPQaDn9LTYZ9+p+B2
Or9KMdYm6Htq/+Li2OMyAtpcSs9kNVk8DU9lnvlDSLTjAOUOBjjzngzJpkUb
GOB434DrhDG5t02LYCQSOsJtiMHGt3/ZFCMfOk0Jny6ckz0BlA0FB5ioASjZ
zbyftvUQkrd03h+1CUFLKz5X5vauJpc0tK4yBeO9zteUsU2/hz8rdW5VGsdU
viiq3jM15ruuiQkwu1NAREtuEk6xGknbfBiOSuByo/tvt90BMPkQ39C7RuP+
f+5StsRMK1qWAyxrEd90nt3OZ3tGdPKUbJhGOPYmxd5AHPfxCjRtj+3NBmqk
aE4IJy+COuHxd7vSLhKLWJSFna+wfQ9r4REPXJws3oYiK6DpLyIySxiT5sAb
W2/LKwVYRn211uQmv3LFl5oYOtsO73dj2buaTi3b09ipDryhhLJ1A34Ixa5S
lfIwaqIOAtnSA7YZFB5cxxICqGEh8skIVpIsAvpTmfEOX1VWhxQizkWTLMeD
Pzzl0C1aoIKTM9u7lrVyBlJ4+ykcwiMdbJInRCl0g6f/9cW1NfgeIQQyYRQI
d2kzHN0qnM901kt764IJ9RrH31/XfHfG2dJTSR1LItU6CmxLvCurflN5gY9f
+hUK8MLJ3JQJAe8UGoF6Yu3ThewGdoyqZ29RJlVZluY0QSTjHi1DFk87iw4F
VW4Bu5ai5NnFZjGUiH/dSHa0XbF4BJtB8JUBigEo3ZaQR4ouF+YPKLVSa/G2
zu/Q5y25xMdCHkw+PDxyYnUTS1EhVr4sTWP4ll6PwtGBPri/ItNARSZN0P8I
gaMG7qKIjpy5Y8ZqcvG8e9p8wh0nK9/QzAoJGdVU9o7cgJdnUWiCrI32Kewr
jZ7Wm18iHAsUQ3wETy7uHFUZnR9Ee4FSixY20MDO0cv7hwCQ15YBj6VVQaLK
2SS3A65IAwzpEVMqcGYaQMlaFwCF01dhQudBt4qI9Xpyu4mTo742pVVhZYO7
/wSW4/4O8iH16D/WpEIDZRThfmnvli3EuWdqrMmODIxgGhvwc7QOmgtQTw+J
rOwqjXvxl4XCdgt5yyxpHUdjzLINIy839hhOc5cv9zkXwvD7gc8T1OCBr4al
rYVVZ1uY4oY5bcKj+w2Q836bDwL4NS1cl7oL19LeMnUXmQlFH5V6PnJh+ify
gzXgbiTq9Js1WSfAfqfkCALshp0cmy8ZcPj6Vw+DqRjHZ6Vr2fDaHWVZsc0j
acxiWZohq0tfwwyvdYYUbkXrDw1f7HRoMOm9YPt3o9HXofqfYDpHrzX4dPfi
PEeMcqnppv7ND1bpVdm6HixxI/ihAcVpwSfnxxmZu6a7MpzbEthEojT/6jAU
VnfsbVg+SU5Dg1XyLEzbOriIDA7GGsvGVSmz2Wnw/IdcZKSBVCF0uiRhImni
tHNTEcVl3d8FDlAq8QZOTlm092mguTmwgqm35MomOwc+BdxHsMYibDQHAhEN
cwEWAtZzl3yiT+UoAotMDjER+t1zbhVQ0BNFQBodmGl7uIbmhajT0tepedq2
jh8g2gEyDyKE/JBPZqWoQQjL3jZ1R4h1f/9yfBcevlfcXEebGJZCsqm58Fei
Rn9Sv9SP7IbH59ko+ttUtRPgjH0HSP8fh/LRWVOshuZAcwyPzc5hcyYzHJ4W
3Dqts1ERAuwPU27mG/xQ/GvRdLrATuySk6g2QwZAjIDO7UE4VdNrpeZhm4Y5
7a25eN4Tn1kxDf80Dw9DFoi2rrUpmXWmjZWju8NRQMIKESgVGGD9w/T7Lk26
Q+32+VJ/AszS39B5u9Ydf8ge/0JRqf+n2qlLk0a5XRvG5dpQzVJW7t9M2STj
TWGEIjhEqJuxbjiMc7rl5Ac4Q1eD2svt0uKfKgGHqfmA/Yis5+tdHHqOD0kj
n3Bc0TdAFN4jWXIEaiyzGh9VSlAqhpanGqtlORz3Jrx0bVhdiE3/DTZp1JrC
Qfhh9wyKdSt22CHWRlMWBZ1ADuuA1BrOze3JEKaPqt0vRPQ7QgKNAYUF5/xI
bgnVVQCFVoAtVbWFcpX1VswwaUJv1leL4LriqQbxmtFDfvGvOKf1zwrx2JIL
lMdGI/Zn4Z2uL9LBiaQheSTrSX1Y+mdGZKVBe9S0gREBzTbWMuGyd6OMFBGt
cUacEQd2v6tWql7ZVRiOn8QMyQCTOkKYdgmfKVDhEcINpR9jDYrEp3gU4+IF
F483GLKZaQDJqpOG4hDJYI/4CBxE8IRy87TwZJnZLH/fOdrGuu7BYKnfq7Sz
5zKStWmtbSi4gbGygistn2vo/BDti4KGuM9Fvz/Y7vZ4vCQ2M7dFhjQivp1x
wFCIMlk1eavDTlbxaswfvW6kSzO7Am4at3LAuiPMYlDxknCpLW/M7ykyZguV
8CWWWFJ3C/LhIcm72obT2wrx2UeftPMW6+kPGPyK12jgd6OFn1smd88M/2CK
4KTon/6slFkQhPq1HYbfdxYff4MvxH0PL0aaA4xV9jZTRKoCA+6MZZGVlzA6
3CE0CLsl0Q13ZvQpeSZ0X1Hrs8DST0OnajvNDsI5feiwNer9Kvspy7UUMdK0
jNBz/jYl31k3PlvDZTBSVgML1dsrm5HZaeVcArrWOrstxBnykq0CnE3CPsxO
b+rK0z9FSoYtEEH2fXSniuN01C2QMfFdm0Q1nQIUBFrhXIIQ4QCDEKdp9wSv
URUYNX6Tfbm7/EMwcHsW7d0Nsd2dauwPSTarAL3ruDH4xtTExAor1flj7FYu
/eVNi7xi8dCwstreRnU3ylzyyJ8rKTv32Dbo3kjF9sC/885Iq6MOO1WyEgZP
2tBbZlb1IFH44jTjZyCtEuEqiAYMdSE1u0kjrbjZEvKFn0VV6alzCyWNZnU9
qeSDiLCuZ4LBIp/YhnAiJDzGzYrLSahI8rrMbCDUuXiUrCVXdkIkwdWGd8+M
oYPnFqdMQoxj0SKWEST1aHhm9eO0m1t2KofAoOUguwRGqdCax+YynT1dTAWX
3/krv1MXAvXqBR01AN0ceWUc+TWOVIPkzwu8luf4sVk0hQyQPLxA/VdZesgY
30Gta8b9Z4m+nxFAHmU76rvi7txsjiTDhqse8UC3A3wXE69P3VCoHG3txjrd
mww1qLUmHoZstkbOHONgzeFwbTw4GrqDv1wxB9c5uLke1AQaG3CsTb1GTG8a
BR9UjZ88EsPgmJPMSJOOuCQSOs3Ag8VvSYXbU+SW07CzFwfU/skUIo/oa8ny
Kl8zO26sMbI6qjc/vDj7qKbWcpdWK6251U8QP3/ejjbntJ1AO5MeXVDqzMOe
dg+UBESlOjF6FrA+vSBwm3tldb0BG9eY4sad2LdNXog5UaOAZf7lpW3zpU6q
MErNUetguqxpTJABJDjNZmqd1CSpiiPyKaa3AUg2GteAuWs6RnkceMMBrJVJ
jTwPR+46o2vVcE0RO4uawFV0dtdcGZu/UnHvMu8TlLg7qjUggq7Xm0MSNGJa
C6yhYXrI34+DrnJfGenV7h21ll0VV23z1KUUy9miziy1pVWsHrVSZDaDtpOW
0kvztj/eleK1HraIGooiFCzdE/PaACmg2SOCBkrZ3zlYKp7FxoQi2J+45AGu
Mw4W0wiAjlAguB7SJ356w96rDuqZCjRFqfjrMB1uB/LERSndFO6EPC5bDvN0
fTV8yKVvNu+EMcz7Lwu0glnQ/eG8kIVcYbaII/0RWHiHP327p0Qu61uJVT9U
+/tFaQ3Y/2mM0OCCiEe1hXtZL4L8EfjFLkz1PYChXjswSnhg1ngNrXB/UqqC
zTTRxs7UyssVTdTl/fOjU5hGllMQ70QJuVIVhPguji6u0UpMGDbUwa7iqYwz
er5sGY5nvRcOa6YfYbEFm5wNAFismDEuSn7XL0VU4+EFVmB4uPcpESeDJynI
TUf6EDT7xdOs7D/dYd3sW3g4VWVIGIjcR8X6Hn4rl4DJJUzBbuT85u2N1bKg
rGYFaMp3NxQgMNFaEeq8EBwYmTP/Z+EjHyQqBPtXP1z/cfxqU1ACw27+qRuW
hQIcfQ39GcVxrc1IuaPz9UdxNe1/A+D7xLEwiW9TTAbCyqO4qK9yP7nV3nJu
5b9+mQmRolhJdEzAwTEP/X7rV3NcLthQGG/u+R5BnyPYyDsnSo4TCr6xXRNm
ojJ0o3fnH2FLtSkgUdqtMMO7tsJeILHx1anozWPFZ1TVeG6NJim+s7rKyUnq
XCYs7QEf5U1/IabheqcGe6gcL7E9Ce3wzNPLAHZ0CBqaMAvtcbDDhov7th9n
rv9/GOlAWRg9gP7PpdsPojLNFWCMKyH1zwFxaJ8F+PxCRkXFMaTQw9ifsmXI
kdrlp3CY5+fZfU1lNETgAtousTGeUFk4xO9Q6thszDs+3X8Q31TYq15sVX+1
MtfVjNG4469gLHYlWOefkpahOMPqBCoSbjVQiWgGNFJ8vjcMKIIUlNSOKA3i
STtYBv+ErWkCsCUG5GOn7zVyV8G4zWNYBweqBxKW7T7y7SMGOJdoiXCn9Wmm
tD5yooZfOLXTgtKjhTpIhL6O79IU4+eBc/VkhRLnYGC0i8QhSvde4qe+Jdjm
yBwBEHT5ee0SUILBoQVMbEOR0IgRziBoKRTNtyfU3jtuMNk34NzsWIAMvxj4
ovHqKamM1ZfGMEs/p7iTrX5nNrJhpcbvYY5OfQMY/AMdLxC89TJYZvkA4Gbq
mrcUi6G6Q6TtS8hN6RhOJ7X4Bnazu5vPo0hE+wQpjZc6x41rQxTFTwqosNP0
13J0kb+7rvqt14AcanVUcUGLshrx++TaGYxB/wmP91vXKAFVlZhoJRVL76Zq
hDqA3PdFxwgmZZFgX2RjoMd/Nb6IWMGkQNPWVFZQcSq0KCqM/bM5s+6oeP+h
vpWLbaaIIaMzvstlStVUDdeO+eEX3Rwg3FbF1C32NA70Ctre5Ll87xt6UXr3
4lib6dJValJN+/uTtHFcZQ3xRdYib3xsixcZuvYQorKlRcC/bcz9YH8V0HhU
BdgcdCgU8u7aqYyNgd5M6XAabN3q74aj+x9F9NvnZ3Ulkh/cciwZmob8N68d
M5w2eKB3F4WivxR/yLoZNhU3XSdCOQ2sSNi3SoPQ/kH5DWuG5l1vGWztyCJH
nQJhTCATanYLIaTh0tYqBKsazMq7YynBDdTFqIalIz1wv4ByaNZtl0GhE577
MVd0j6wyRZA6atqFhPKFsPm2M1lmF3qCg2R3RvSX7N8jaslsz4fLNSD+Ecsv
9fr8HNJmV2Z0C8BsbSDMlZi0MrTMFpf/+SI6IFDa8gZubmNyV568mPCqHzl3
Lk/p91L9J1CMC+9XNnfHkdF8FEfWWgAyvwVgeLM8WmX8tAdCbvV363ERSxth
ed0V9WXV/mo6ohvLRn2rKCnlATZeCAtqXABt1hhUPL56kC+hVjX4bji8DCnr
EzbtjMcmRqBOiOHlSzEWbWhTzhOpVJEpn5S9nhenVXtQy6VdBw8YfrajMqdM
2LJFxQPIkkXANlCo4fZJ/UcqjzAcp6pi3S1F11xcOe8JpXZvLIAWNLti4mxn
AMj1vaTvO16CJGs759ctvieweeWyLH1sALiExw3BrQnFBIlJy16jlnbqH65r
eMbwV8XXTkj4Gdo790d7EYLZN5n1+EQqbbX0VOtXB+I/Vx7aKE0Os+sQqpnP
jcPCrD2+Vxl/KrffLXLvmBndD9n9GMszyD5+D0MPda2CnLLwTaiyudTFTCmR
3hQizjHFD5lmYMKBt7W/r8lVmo41gomaQQ5b91kQu3/DcRz/p0n/TYi5Mde+
fis0zCBepKex4yiqkmNCsp3JhOugCQoJMp5/xjKc32N9O6Y70eZYtQLRCuO8
Zdw09OdADeUUijzv1ne2tjVFxdeibSg3utRsnVdJfvr0KgiBto8lZAKr8iJD
cCKNa1b8Jln/+mObGX1IA9H52ZSbVbLlILEBl5ew1ngwv8YMVJsos17uBGPu
ZlFexAzeuefGA7rGUEJvkuBUsBub82MfxXw3MGCKp95xbKB/R/cJvV7PE3OV
YlHdMVgf5MR86sJ4yp7vp5tPLvhyLMtSKsV4sehkO4xBJ5TiIOLbjG6fd83T
AD4mAM8vIqOW5B6YaIOPBStiMEJDXqokzvGHcJ5dt4UNfPjwWKg6wK6LBZhp
lEmScNzILU6q24+jDnuJfY1yZJ1ptAZe22IvH6fYaBbvTUzQQUigpR2Dm3G9
ovuOKZ2Qq6DTSVhH8Z5rHYuAgMgI1sPyc1+/oTGE3tAH2ICWcDmPXi6QWiou
eSiF4xX8TA9lil0E8XNhI826o60kp+5MgR/g8E7fALBGO1Xs8CovClP5MPhI
eZgCNXEAZwRxHdq6jX2h419QxqfSjcgj/U2K2yjuPx1ZwMS49EUU5tYOGk+2
VUq/rKRLssFb8a7TL/ZMjOFDa2IW3AjdjcUn/JS+9S2DhcFThfLYgKB589/t
o0fPIzUkCtTGafrkDVdNbK/QLzqifTqkKKQK+oFNphVO5+X6a9u6F5d5NTdm
EXC7Fv5pAsl5Yk59IAmMFZ7RKJ+SaTEVhc3zdYz8k9FCvu060JNe93ctFDrH
2dCQZDLhMdW9G9NY+CQoS59ZO7Wp8YKDdiGD+kigHj5aO5aXyfqHcp2N+9bZ
cW3zBUmaNjuLxmX6KDyCckRY4OBDbJt+Lz6M+j5nImp+DeA3qQhLD9X+x/qf
q/6U38St9kWSLbTQEJ15ILb7ckA7lmO/OhKiUtqm55JXsV+AHqPqIVnS2+SZ
774+yoyV+IPSyVxmE18lnZQ0HCrGmQUlYGKQKmJPFiSkXmE+TktpRj/jOXeN
9cm7wNLinaU1TiDTxDjopEI2fws6a0kBdXa0VUKZWihY4Qt8C81WXRy5Vpjs
gL1rfHgobG6ZUginYR4tIpQmxaC9ztM/sXyk/1j35+7FNgyYPylVaYBFRnyx
83pjgfDcgEJk+EPMhi2Bn1gENB8HaFvPg1UA0gp9z4DG1+E1Dt3wJA2pO70x
Y2UL1E7C/M6sH8P3VL6kTZPN8i3TiQAcEwcFnS77Vp4pzP3gL71JxlgO8onL
YbFj+wYNGXefoi4qOJGxKVAZN01oKlE+moNM6MHmnRN2Q9rOXCnA/lek7UYR
axM2ejJxzErWoOq4TosiZbA5KmxisIjaSXDWcDJtHZ5lQOnptloqSlzesh3F
Sg4SwwdrAn6YlD9hKcIeMRNB5hbLr4+RcjYqHFtP2RHkp3gTmC1IT9N6MzfX
G42UxNZctHV9sEVEH1DleFKDXFon5P/9OKM+Fd6dqexwstFfEEKd22WvPic0
1uvk/t8PCzRw8V0R1z1jgmZ9FZ0Z5pDPRCcSrzsfgou+fOSyTMzKrSQQSgz8
n92sxR20x+kQf0q+RQKvuMMrgqSZcBZ2HESUqccxZcplzYmwZcZOvQCBslnC
r2Lx2BHdxepwY+X1WuB+bSNwNwLr7s9I+WI2gjsybdsriKYZZmS0Xb3lEQT7
9cP5ngSV7dzLuMju5CecYeNvzzV5OumfBD3MnQMEPOumNu6GDbue3Xxl0O+A
JlRC+uxrqG30W3RiYPb3ChdK9IDPh2XfsAvsFZkY61V6FGJfczEJuz7Fv7Rq
i0p3vgGXbRJ3mdBKxQsbhVJbYmZVdMiIjHBG6iMKeyhGUrvyEJDSPNinVvDK
UGSM8t5kds9pFjJfgyLzeXlTFNJGCfCFAKlPIqHLWghQ7+Fh02YdHjp6kPqi
n5lakaJGOe83iT9ld0rXRrxUQrVUVGO0tC2ZzHu8BBSIcK7TZBg3s5JXJZVt
pl+DmWqKpce+OKTIW6FZ/Asp2P1t6lwmnjsrK7ZklruiZi6bDYDrcfNuMwax
sFk0qh35UMsG4fZVYPLmy7t92xU0PRNnLrmYrlLivDkyTK1PJAfR6LR+87uv
uUwLLC6o4KBLK7kbntxvXkA+LksHckoK0zSZW0gJ427Uayc36RN3GytKI5de
E/0ExsIh/LyW/+6Q4qJAqTILtQWfc5jzEfzfV2xtzRaMtZu+G3vazgS16A0F
MwN7JRwkues63hdgbcgNOr2Jd84nF+cKDPUbwtxEpKXnRWDjdUrDyKKK8wNk
VHgQxWeKO7N3Ng5KIgJhPRPlLqArysf7ff9bhdio1O8bD7/g5i/OuoPhQz7M
rFbGhMuJIEdKq9GHr5DlgQ3lxwC0f5fuA9g78ENf6osIkIWq5Mt7Z7Cw4F9q
NqXwpI4uJ8MZ5bkt1thUwIwHJFR4CBi2LMOzpXDDtblm26W/jyt/QB5S+sap
pMEdFWzQTBkmeRBzyRbir9aj+i9X9mwjLGEnu0qa/AJci8Cnye0qqdI6Jpke
fQQSfaLLzPvqq7MSIQ92VjEYcssl0nplu6lzii4V8RbSsfnznXN40L7NjIk4
1yKtD50q9sIrzGJLZ4m+GdQITKc3LOwEaqQGaYQcqxfaN1kHUQ+lnS7qHD1n
TLklCnbspHFsJ+5OBJ5tvHsSTgStdrqLf6M4TWXP9egDWvBIKwa+l7P9pLlk
z2HqHKkX5PmXf4SY+Qi51Rr7pKN8eJ08KiPFMLdaLDA593UFCxU2uW/ZM+vO
vzlNRYgplDYkjuoHxZLygaBW2BosJ6ZtYRwS2NklU5EyhPUXn1BaifUUI2ay
9qZP86KVQ8kDMvramC8w3QllcUtXp+BViSsEKv+h3N0Blllfzufuva0Zz9qD
dOwzJGlOxg7zL5xWtzn4UGGO3JASeH5izg9kMLy/zK9ucX4F111wSINDO8LN
4hR+JSqmpIt/Uql41hd63yY/yOfKABw/QH+ogZIC9ZvtlVgD0mwMir5crnvU
YOUUxlcF1i34+iuz6oul9xUPQ1Ybq1QrBPrGkqm27mKpHn7XoNoBgPOPWNoD
8WJya9gHlcd6UGgvvIRkxkgCqWawHEj79PHyYOWPbppIV+Jro0SbyloKMjCn
M71zH63CHnJxD0Cj4pokinthjmtJ6ltHc6IFdD7aWO7qJOiTr8/LgDFOdFr4
VPxH5H1ncDVaxDTiGIVtReHGwC4l3VR4Y/SgLpQkdqRWoRsDlShF1ZTF8vz6
zjRdRoNHYcJ8quG2B8lyZVuKwxdE5NMZl390lDPT5T2LFqY7oLh6YuU2tWeE
B/nzyWCmSswacRUTYhlt/BTBa8M+wu046fln1KEmeZuZZQylINfPPoq0MwUO
smEKJH952i8Kop18Gk09RPci3AdqXCImhWQ12bhP0F/A7Nu0xU0lGtcmutEi
8DnkDTDlr6x7wwCNP82eloCfV1yS0ty+hQZ6cpExZVzmkOVO07oUYdkcbVAq
PRWZX5UwmFt/4Qcr16mIRRxQpaEWviCmSODwAFzdF4zsgmAd7dytUSud7+2R
wNW3eYfEgp0OvkSa5B9DPjs63dTkVPVwKKsDgbklDYfn0HoneGZiFWhD70Pa
etwoELrmcy2AQWB7D4JrVMRXEzDQ+ji7dSCoT25xVacHhiFn2mksoXME0YYw
0tiyKXYkdPmLrWncRauU8or00vj9enNjU40BD2eL1ZA99QlDwnKy21qBw5mC
LEof9Y9UK89RIpzk87TovKVfDeC/dy2zNtTu7G5X7q8LWLR41zTdHf7M4bye
vxkfyUxp1DydB3/a++QB2HRgGdNplogzSoq1r9i4EaLp6h8lm11VwnqXGe1s
BvheZLC/5TGqb5ZEymv0n3QIhq/tfmJWoa97aeenP1QgcJ9oDeZx0W/ERlov
me0erXT/GEOYowHe7KuTdwVI90dUwN8/iv3t9XsbIC9XggThVFb4TB3SR+Fe
OvCjqnjl6Pwo3xRPgKfpPVntweg8c5VsG+3qcwRGzFZ4c/SrV8Gad2rRfgDQ
Hx3ooV0pP6QubevS4i/T/CjtYL3pG+74ye3GjprSWXsTQZmmmi0ZjsdeQMgl
5mZxyNtk8KhG6lBwUQLTao3SkpirmeuuoDUet9/BS536GfvymylsrfuCEZxf
OuhNOkOww8l5cVmu+eFkJ5BnQkR6fo3VY4QOhDxbFNuy9FGRopQnQ1YHv2yO
hH7vkATRPmCCKKW6e1MV6oNotGZHmzjUNMbWC4kq2u/rgQe4wTQmg2CWRXfX
IhRaTeQr+l6IncbmMkbHx9IBFJWOjmgN+5yDv18BiwPfqa2sCvBBKI+0mkcD
ffGeKvixrQ31KsmsIP4CQTNPjD4ndDmKMeYK+iV/AA0DfBCL1XkODA8n2ZuW
h70DPM3VSzsHb+gF8h6bRgB+0+oOwHuR/OY1zPOJh//MqYQbvcd76WhNLpUe
UlQtjzc0QrDO9fZ9GLuoubmYVK2lm6N+K9tUsoJ06OTFv71NVmr0W8qZbGEd
g6MoLvW1Lf0esqx/z3hUeRj99S0IiO9zuArKGwqRap1gBJNK4MpL7JBh+wa/
tWB1uBh4GcM09BSJyi2H3xAqhuIotvwMzsN13fhzlGvtCJsX9J5clzc6gj+b
/1ghaSYdAOe87Gftu/lWDweknnKPNFaSDCY+NZu55QPP+7LS0xESwuvIMcVS
bgcePJZG11Ft3gMHjDzpjZJLocos1yYetEAKTZiGReU9SpuaukleiV9fK/wW
rTTmj6sz78a1hFjOu0DnDpLWIvv6t4vLlO3cewa6YrUwyWbE5iX+245S9E+Z
oOIlGSdkq59CyoBPUsEX/uU279bG+X0Cy7nlEIroPrJ/pB+GytzQIZySWBJO
eKucVCUQrYx/wc++HecK45c8zKt5l36CqTnnV+9R5MfxNxAw7yOBNSoK2OrC
+v1HZ6DCedBejV1c1Au7vzIspEKDtYR/kopb8GRWGzPnHkJtn3ihgv3kL168
Ztzgx5vMdyief2GxpzopjUb/7kqH89enRY8xowSa6EO4DNACnkn2/5M/qCJA
+9Aow9rtvK65vTkzJiZHG37OBfIQNFJxeiGOlAHBlBQsEbJpZPp6nbgq8PY8
3cGtmPHvDCRqM8lVmOLyFLtoUEyTJ9ktd03MbKLoUBWb6NBedcbRxIpDnWpt
LlnwLZdZ4zQvxj3r1esy9eEZx3A/x4LgYwfU6v34SxSaJ/uYV8hGZiUr0T1C
V6L6ecDLgNOQ9CC8uiJZdn03lI1aIxQ1z29yDcvxACjs2goONmHTwDErTFVL
tvuM2JPtUezXMpw8fJPbUiMFblm/bV7Kv2YGehqKHmFBzPahXmueCn89Vduy
luvg3aR6dXxELFd8l4bWyaw2yfI5AkP8qp3vy5jysfiDg9S4KoDeNVWD9HJz
xwuzy5TL0NULuDXRVmiYArtEl0UxHyRGy4mX+1GLSQjbwsyVcNBIPCL+NkNl
AdVbv/7cvBcW3mibYqeD41PZRial5rzJjtgMR0s+fMvPP4jd9hrP0UMzsoaW
Z56FMTtN+rVM58E8Smiz8aOiTW+YCubrRSKvDievp02NERf1omnuQlCddm1y
UUQuk+GqzLqYX0GYMHw2bQDEek8Vgh717/85nf0Y8/bSMzVR/Utwbpwn7azS
FhsRFF+ZH2uJV0jefulr8w0m64Sbd/qjnmWtkL38xqS+tRmRmTlSp9ofzY3c
OxNVwbHwQ6bNefCr3AQxyBvi5nECBxlP8GjMb7fUiIke3moPrSbqwOFIWeTj
ZcZOXKsODlymb51qyYCGDKVb3DKS/d3SlTET2y4huks9YwBTqSN0tmSDrsQA
GMkT1a8tvJJ2WOiW2UafDGxy7ar9kPMPgKRLIzcjTEoqjhA9SJIed//WXrRo
hr6nXWlfVl/9HCyoFzeqaCeeTBA3i9Pj0s0WNAfDnK1Vj64Tmy9TrxIAUCsK
CQC45+O8aSs/wcUGvafnkJyp3KNInyqI+uM2ON+sMjqvoHjkszDFc60eigeV
nIdd2D7h7jQS71kFzOvoW8ONGnniQoOYX4um4Sc2ZQVAPxnObCfMXebRCPJD
M18duoMcb0rQe+DesJKpg/bS3NogEqbofGGHBS9bGTbX3A6Dgv8dNSk3IrF2
vT+dmBYF/d9DxlxAtZTw6vre8g0rd3YBCfedbsgRCPlRcWaR8rsBP/oB93Sc
bg6oVCmQ9UejUru52zgNuTb3e8bYVB+bX/hICJ6ZtkdQ0xb6ZbBma3PbWuYd
mPvlpdlqRRM4wMfaYoONsGYsNZVRhVa1Fx5iV7KQAzS7NxGWo2UO+PjT0xxz
XKBu3YDA9Jv/Vo33y25XqglEzfjDcsIRRA4XnG3Vip/58pCgrF578LYKcUWD
QReBWvkw9bnobm9v2S2PdP0XBmqqwQdRyH+/lLmyV/vywhdqFJfMXHU/9KbN
7EHAYs7VVl1MyyjAXbEWoZ+6c3xX5LdnECXopt+/GQlGTRn8JOqWurbz2Aqy
B0QA/qVngg2vmqodhy0GCJZEwtxROHqjRBWkivvJR7Ubfmv+i8oEenwJygsC
nOoF+MoHGlkgEqTVO/c8hr+brlsjzF0bFRK7twHyJMHaFey5KOa8Ulehhzhe
OY25nfu5ses3UllNTOEpNh1UVNYl7v8Zx5zmdIoZPWsoJQcLvehtPohLrC4O
r5G8giZzPuj4acjPMNxzds896drEa/NUzKh+VKUdG+3/rA5ukBvGhkW/dT80
mLLfCT2uHK7awQGoFF+GJmV15VEdz8sor60JDqCkNu72ufNjdPMML7qeHmrD
b2GDO/4BMuiOG/HsmFEX5rKdqCynIjXyfzyV3H42/nsGFJIfLwdTd8jcBKOi
CZYUhqBS2rqRxatbiO6hmpJz70yrnCBzNJLd+lSnZeEefdmLKskvqN7PHQXP
c+rB+ShXoCH24ZVHJOUKR+2GRL5pwAo262E+bBE/vTb6LcKVpfXVY1yez7YK
rsLaLPmzm/sLCFdilP0Z2uljRFbTU/PKmKZzscXSppfrAcxiU+de/G7VciBC
Iy4UdAn8egFLqDYMP/1sjvojOg0PiR91SKiSZ4QTVE+xe7kMgoRW9MAe5MpK
a0EdfHuIiQEOlOYPqQLMaL6y2qdehe8lSn+N2O2eCaOa7oyeED12RL7q9jTs
LorC8acxZ2Vf/+l1Kqvbfh32ilLoZJLOuDQEaOIyjwR4178+2cruHnhIt4EX
MMIoO9CvLNEi9m6eenHae7r6khWku5cqBFhUTUutQAlPOWKvXu14ZWIZmAZF
op7XdWbeuLLchMSDUPzxtpG8iwBKB8ff/zXCuOXvYplqMV0PkXXYBP1tRUC0
wyxZmCY357Mxb3VA1FNyUwhcLBLuS6tduenYP1a17P5L2hHInuTUN7GpsTF4
ZqC76LmWAvSDIR+1BUdtq29C7KocbA8b9tbx7QhQVRCiyAV0XgF6woxCvRJH
tSxd8Bb1gpVLoOKwXUINtTM5K7LrT9o+K2tOwu4Q1zy40ulx6OAe7tD6a/Eq
VNE3o1o3+7/QYjA+I3Oxfz+6N/PxfiirRM7j1R7BpVgQowrvIpxB8lzQWXkm
29oohrEJEtsIXTTXqEjdy1x7iIc71g9O2tC+UL/sXYubfOqixQWZTcJRIBd8
yug6A3Emmg7LoqgBv+qsNVyhQBqlaa1bgC99vcrB0sj8QjtRRqvq/U2IURvS
y2CejB4zTtizeHhmkzOLi21j8V34qO/btPsunXmRZdrfNQ8KavVujwi8aHQ5
kEM2I1mI0Eq2KXKjOcdbTK3GKQhdOHMpmztm8JaT2b7UX2V0s4lWzEsSscth
2dPqxs8ADanAUjamH1P7Ep+h/zx63G5jkcjs0yLMTlmx85bWCQPfz/c5phWt
zJCC3oqtIcPgK8+WuHa41qUxTEY33PbxV2XvM6GmR6+Jlu5lnyg7q054rYbR
GNcUuZ0fMGi7Il2vBYukFjg9f8cBDtrvhp/WnSvWUlpcQVJNsiE0Qosh47Nu
+DTJUKP4Wr//lVTt/N00qsB6jRBiqwTR/p4hej7PcFK6DwvIAQQGPvUdZ6T7
EuBHHpRT0iB6SKu3NoGjmZCZ3lws91TztZKUTwPEuW9T/+b62SHY2lIG1pYI
29mJdwlfLeyKP/8koeOGat0quwfRS6tMukES/5XPOQonwFjMRprezxDGiJRo
FT4eLyDZZxB0WxyTGYI3WVjlGY5aZfXxo0SvCTr6WraSNezu8Mcqjd6a+TLD
l4kCPW81Uq0VMNOM/iHvC4W4XWv8NonONaaiXS1SiuNGAVtRVaVCqTp5oCYs
lTBR7bdZLG50pN5CqPRk0OW1I95hG+pr1lebfyYUSjRiDtw+CaHGwhBw/uxz
gnX3GaGOBwNEBKZibghTQ8DLKjlq4Npb90bE5cDAaSVLCBF1XLjq1Ga1WOMQ
71gN6pNh1Bf1sdpw88lvIc5ZXaZ0do94EWSaWkN2NJM9mGXxmi2/9euloCDu
ZPhzfrgmgkvc5VqvjWHK0tjPoDBRrjG7xnWXJJWQ23rjjbIH8jvz5l4YWTCQ
UvY8TVEjjKd+PywBWz01Mwf7tpbv2PLNntQxglR6nKMvuUsiA9+AmNxYGEom
vs/jgymJ9jpQA6/UD4nms8dVB3hjbaW9TahiMA7Ls3DREeut5VRszSitIAMA
PGcqSF1yFNSkDC6WF0mwWoxrxDXYgr50akUafxXBN+kS6pXQUetw3tfyHao1
T/67oNnc97cLisN9hlMJqCHqUYRo0Ji+KduTVDeP1ySR+88rHLzXsEtG/fCN
YYHy0fOojvi/CblAHlcArlJtel4dibwVkzEv3rKSGLx7gTpcfNc1PHPPg1SW
z1tQlr0E/Dcdr4iB6+m819pL0DefVrZXc//idVwsjwBW7LPOMmcM2DyyxOWl
9Cd2qUfqZrtWhS88Qkl0+wI3Ne1yIvW6F4LFR/L4IWbhWXuviXbevL2OyWb2
qTrCGSpNLbwP0rdZMC6UwK4PUYgHSMkUlNu36LEjKwmpfMNGx7D3SwuAoljs
cHLlKewYez2ZV6mXnRYF4MFNiVCub6ifgN80uV+xbgARGYqN/F9KvNaYUTYA
7JOxoXJbSz28mMCVT2D6WTJnzci2uhRXK5EWUMYmZJ5rDxR+sYNJcqUhGNkK
8QJXwJn6rGAxV4XmUMztaEJhP49K5Rw+zdDE+hYO3sjBQMZ0LxEowXHy3cMa
VkcZGTnp7CeHeTDiCJLNHHj/JW/WV4+w8YKSHqSi5rOkEuYlN2IfkL9izOcm
vyqjnWuSGoqINvAX1X9Qun8yfA3Dg1apMRxFMRUioQ6ImvYTYHQ450L7IEcS
8Zdz82ED6oWOn6NYNPprqlJFKo7u23NaGssBYA12pikHV2iAshc5ScG7KGGg
2FfdAPR31k9tNxq+NTA+klIkm9V6LCKxxf55RRR+1WUQdDqagY1XIzPUXbzk
ahpUquV/rADticcACLKiD7lSu6+7g2fhX9xCP9nvkLVwiDvAjINeDINrTN9V
g5MTh+s36NGPurMAgAUiWq/LZsHTiHZujEfqxCUfz3DJcZMKJNAsFUm4T36N
LzkvvUWSoQ5DfiQEZMo7Kr1hZXjWEG+87i5oxzlCY23Dll2V1fv4HDadUhdD
mf6oNUtEDG8XLqxao2ma8JyUSkKhK5B/qO9ngBw9m93P/KvuvUP+aMMA01m4
QKUm90aEdCrZi9/64BUUNgmj/sf2SNnHo7LbIQX/NRJpAzoyVHeiXsTrxesT
1FLU3NTth/hC5IuUS5Sdpt16en3pU8nnO09+JPWXrUa116KNxcmukCWwpCwC
5bo/RK2jeQqnS3ESaAGcaGiYzuKuJcJ2ymrvCn4ba6IrNzIwC7WAakY6p8vd
nDZskPFsOuLZY4POBQp5a+FZCdEWLJevkvJUCy6VRG59rBJGnplP60XxgrOH
N7iHtr7a4hs+u5gMH0YyO7a3vxSUucEm+RhDtmQ4s3hKsdjDEkgbS4iRKGmM
GbrywrzGvhFIoRVn6+j+sdRDdhYyifwgdBkt5GlsTeEMbVBY7cDu6F+H4Ksz
JcypZmcyNUlZy0PZuk/Pb67O9q3DZoymqnqDm1UfrFos/dq7DU+nwuj3LbCm
zbWRIbzOQUAHb7L6YVsBdrWQjfVg/CBw0SMifr62BA+hVSUei4aRMriBnKA2
dCaom6TB/nGoC9CkIw7sD4+PN/PfUUtAsJzL7OBLHYm1YwLKIeBxmX4KBJOe
T7yi7r3hfgMU0ddQVhtZMhRpxctRLesFcpnEvEHa4DH9Q7SxCEwSe4iZ4efA
NPPSyICUV1rPKfy/dNPNQ68nu2+dMTbB6JKHMWO/lOj2zhKnVm24UxrU+Ebk
Oz7PhNZ/EtRhTtbLFlw35SePZYiC5jTUs3gh3oVMixVo5CNaQ3yIr1EDfB2V
tEIBO8AvdFUL3E8dPpeBLqY3v3yD9CNUy6yASSW45471q6myfnEUXpE3++av
BqTn6zeErgz31KFO4epD6FjbETjqAyLfnG0sKiAtG3P5tNXLPD3p4/4MH5DN
VAmCePjdg8/f/DfbUccz/52TOT0KTcFE/M7I6n0sxQnyDM/b8rwpO5AZyrIZ
bOJHRpHRghD2zW7uL7fOYEz7kmHfknKC94NgmKjBnh0fS1zRtNvc3UYAzHqv
P18nTKj0zUkNhG6NNhUgXqpZ0eaB7yoVND/YT1T7hp2RrpY6sfyzF6wVPk1r
/rpfzQoV1bLtpITYHqdFyyiFhxmAGoSRNx5gSESe6/I/oKnjWRynhuRAdWWg
UNCm5IMeAoDO7cBo7SznvBWcPOZF3dTFbAUSXIjW+NmfB572cqL2dNUtfup0
meepFv1Dfa7aU/oHpiKSC1XREXrNGyGd8wZUpg6p8rfE6qH+KE4bAE1vDVia
EatbrqT47Mf6xhU8MrHi4o/gndl6lf1bFNPco+UOdHHcZ6E8J75v/OA/0x63
YxY7vUYrlEgRgWJOREH8s7/wu2YczvxjFfFvtE4UONZFRZDKJF0zuvCD7yC/
FgKVNWwuU9XMj8XMUKGMa9V6I2BpSaAdtIiA1+RIDCL5H+lg2mXJ6d3bP8ES
h+brkX/CJ3HqwaAjQYz/yWwrJMt7/qpA7AMa6NV7FuVkeoY8QspcZxEppWhW
wFKk969ucnogbyRkutfz0QfTNncNQV1u+VwGF7mhO7tImZnBDQgmEyixZM3U
6yThdbxrVkSIYpJZwDIqCs3SZCNc1RL6cGDTEKMNudI1l5AmNhQORNiccqDY
zJQw2P+GmGUh6AyqNZ5FOIyO0fh4Avzmh2TpsNKsCayjmgSy38/OFAwENtMM
/bZXkDNkFaoPryfu1zXA+MFE6mgp/8wtmTDxPt5wtpMNQSHi/tMe/o1mxtlZ
VZHO8GviFjYJeWTUWu/XsELdhPd3cjy8YTzhCJAR/9NCfhd+K1BYQx/GCyno
NJtnTn+A0poEosSIlrAJ7OhXY+2RTW4qeqIqiT5Dzr4RxMFnXyrUC+a6f1UV
EtjBPE148OGf7mc8y6CPRhVzUI4jOfskFFcNwBbnoBqAd9DGHeYzWuTO/PwI
SR4v+YqOVHSbR1yNGJlXH31VV+pN6RpKRM09IqDMY/EkOGJl0Mfg0n1g7RIy
x6DDP6q4nYEc0ZiiAUi4e7f4B0WolEMVpmYKauQiuIwQ1JeO6+DlaAn2OKtG
wdVAiv0L0fYymqx+uqExqOhz0Ok7Wp+feddbFFrW8BSvbP9GUK058ZBmLxNg
l2jPSrr8rsmRJiQts/fq4i9akvWA0lDw+lMAY1sp0Ox2S5wbLugL420HrZRu
Ws1rPdirJxoBh6Rn6Hq2Oz6bPjip1PIYwwieCAAmyuljnSN1P40d4eLLXWYk
ZkGGewS4hSJCrjiJL6Z1aGm3WRmvAJjlJIU1Vy31WdPozRo2vkglZCknsEEs
DlkAvVYMJu8Hk92reF+LZPonjjvUIc799kK5j50U+U0qtLZNSbqOpSsvU866
AhRWb2UfMnS5tfZQlY7T4GfCWFeVudW5NxzLsMVlRXj+EFp34XcYawPJarce
piC0wuNdTxaFny6fhWGNOCR/yftoXPtRiYw05C+AZuksJX99Xqs19DZVDoBH
x/aDZbVz/Q7gvLO+fWCfkcXGHcP/mJJ8vw71WLRxfBkrtAOlHMd71g8qmgpb
2KTZk11oDINngI5EFX08YOmE2hHzngfhhWjrx29b9TaiMg/TZtom0nLtwP3/
u1jNd+WayZDeo3v23wa6CAa/Y0mZSBjaKDffckg75iuRoKqS6Il9YdlZNLWy
ca7BitMTTDMH1AWa3B2iRCxnCh75/WINOJDSJcQLquENsxHqocxSjaTITWxY
823aRpp/nK0MjPmMag02n8mw/VimPy2QOiKKmjStObrCS2prWuRsIgCCvzHp
8UKUPy7knaCKIcJvLIH+M+1MrbcQWptH/jhbXu+Dl7S+CEDHg0cG9lxIO0uo
VbkBgx5HxGXLs4WNapasDANY0PUwA8kVfY3DkXSMYQ0g5MtVO9SgQnAcCivs
VD5tgSWLn2FklG7E+bQiBGNKuD6M+xOVcTceMW1NVZjLsHVymCbhddKp+ZBS
6BNwAg8A2kLpYIGHvnxkUCA57LJdXcmYCev3uvawwQSjm84bcMNcgePu1q5f
5ScVpdTGesz+6O/g8tBO7fTzpLA5lHinwW4iHPrmAsGpaBof8chJNuLNItm/
CyYdpWSrAc642mlDHixPZeS8hYJM0XYdEVAJhrM2znmUFW5m6LnzxK9ONMbZ
0OF2Dnq8u5uZp648T5Oi0zpookX6hvdlyZ+D+56yN2W/y75M1JeehaFs7Pvf
H+DRx6I7KuwltljW9ScPPaDmmoUMabM0/8WgtB54eDka/lUWeG3/KjQRU8BP
KPCauFYYT5VoB5OslSoC8391z63WXKelwioMoJbs+zRl20hWYhx+QNZlXl7O
VPdNBbInbZUabNixGNtGnttm4ihNWLm8YOl8O7zOk8V6vJOhqiboBFWRzkk9
m4o/CfhVXyMjmnZb5q5yWHSy+sKplm2bi4so42YNoOP/cxP30gOn/3imet0l
qiiqGQwcE2jMRUuT9oVX3MYCZdr3gi/2j0IkOTOMOED+1FJ0XoVqtgoAZAOJ
qphSZF/19X6YROIp437O+Tftt03qTE+bNjNX9H3TdUu5HcyfI0X/Y8iPjNUu
/yl94mXi41Z3fuMhyrdj+ElgYbKbmJl+OMJKHUzflxdVBAhzF00dNoFWyPQ3
LaxBKFzeK9gPsR6e6FoSM1DDcKmZXPvzZhFKqB2lYknwAFYnsOOsE4qPvnl7
YEAn1Rea8obK8NWot0U9fj7A/7UkYtXdDnQ5fc/ZFXbYr0ierbY0diFY66XU
WqfOM9s10eEvGXTe2W92MLiMzUKhtQ+kMLyx7YQB9KvvRp2+6RCY9BTy97ta
4BJrK4o1PofJCzydNgAkXQWpVwfQ/6jk/292pqyTs4J9A1ktn4ZAl0xU/h/v
83tvvpEo4jDr1DhdYeoSlr/GRvy7wLKBQ+QGqN3L65ZVNQ6HqP3rF1BeOWPM
wb9PTRKHwBQbeYWYgRzzxPoQsGPglyZzfogFQTrPnv5eU1vK3Bqv+W91HHbM
ok4w4UILVAb9zBL16ee+Niqggm+zqli76WhgbAL7sQp8aeiD0azL2PxNgDhx
BOIVT1bg2g7FTvsjCrH45+vGtVKGYhCdRXN+sSZMUeIvWZv/8/iHqm7Enw/y
XCQ9OnHmEP93ZMfXmFsJPtABHkdeDz2bvJVvDIzKmFBg1Y1Yc0hR1q3hskpo
CVqFxH7XMlM/Q72pWmtptQ+tfiflvQQ0v6I1CVSuUGEOHOre5ynk2SuOVRhv
sQ8IAQHgqZDuZBWyWEzp/B/J8z4FqSZd/m2sZCvw4KTHTJNoeVOKXU6xWyxb
mT/ipE+rSE4fJcrjiV5Md9xyMXVnCKv13+gp6oaclYq3Mh4ziu/F0P+kgwWe
VVd5U8E85U7eFSIW383w+agNg/4MfSDvLqmamCSPxkWP43ratdgGB7KTuMvN
L7tnUT7ih4T6TlA1NNxmo1Cs/liQMPUSWoFL8IXxRTd0df4gFeMFKFic8l8J
MF0BWX51ZFTLqEgEwA1KzRoRa1t4EmX7g/WRjtJPglQmnE6L1fvyLxrbn8Yp
Qbm0BWJ9fNxVSr7SkYxpvQ6AiEnIzgcND/CuMafs1MX8PaE3gnwQzRGYyTRS
JWonxLCN/p5EUYsUw39Xp/gmOMq2qH+4fAwrdkAIKWTRzIIypY3zl7NHFgKl
HiKh6/zp75A4fsDjkLEhnRcfclgQC0Zjl+HsET10TrWAgjsvi8Kbt5jNd9Cc
SDT5fGzUzcU5763Uqb+fhTbEbsUgPATQX9hEtxdkV2CIDrLftOJrSEp/dODd
JqUFph3Kw3d3eEBJH9lV1F0iVAX85btzeEXc3nsLTobG078I0fVIBRf4rra5
cQmVVeEng7kBpnjgts38O+4D9LvFSzY35G3/r6RfngOjDlwJZ4OG0ESuMzoc
QVp9NLmW9CX3kXXtCdDTK0gKCBAMqY5i2y/vVDk+8JdD7kSxZNtzyTU6mKPZ
WffhIConi/VX67ta/Exx3kWelLh3HtSlI8PcZmPblhw66r4Rm74DSz8fA8hO
mFqZ9CBSpB1x6P75KUsBngsON0z/r3lvbKT4lBbHdeHyOnIx1hP7XCrAESos
7a6//UA906/EcuwoSiDaXHJKjLZ3mcsLNNqP/z1TpB7HLbmcslj97BBzrI9R
R0ujGTaAXubdyBzaYMLupDDqaPWDQLSOalSNuBencE/xxGhOlSll2bNYzpPc
cYt2U2gAexY+L1daQOGS7IcD4fj1JgJmYo2HOIlAqqxxfO7BSR3Gj4YvECze
MXgKT5bZ+T5RJL9JcfThOKUjOYw4Cxu+tIMOHq1tzq5pzVItx7hsf2H/K/GK
CIub2bQRZLyps03qAGw7eB0qRc/WrsnoNPn2Jzpgb5IQDjrqtDYMQ+m2z9Id
dKxxWvSAzz1qgEIUfFXYXSLX7woEU/9r1NbqkV/NeY9XkkY3Reesc5hfdeEw
Los0NM/AbEXBVM4sm0yQwUzJt7rA3Ma/TNWedfTqT97+f/ket8bnihOh1Byb
dmntpko7GYkcXVpXCA3TNtLh+2reF1MXob3eKkhMqiG4eQypwDiwsB4aAv7J
S4Br89q8QVIX/8cEluN0XZ43TuHLsO44OlPMlUpFFcqKVI64cisuszbk6RbL
DMIRYJGTHQVhvy+UsJOsdwfEni4DmgwOQUJRJQPS/D6Fp29uhVN+kLRw7vcO
QV1NETJlwj9TtJGruRcYchb4plXcUFiMhWNNPCgBvzbnsD8QFH4EC+qgBOYM
7nCMinhpXv8+yOgkIBxV5HdlXAXTQ+Ng2banGzNdbgsO/+v9ayfUJP0iWe18
9PkLRpLcC+xzpjcn4LkA/FVB395RnaQTq7u7VeMA/MyD5cFMlrM/PPY5ydkB
GtPQa+P51ags1TrFfZCdj0KLuviSGkZSjF9KKsxrYTT686DcFcM3dff/PyGD
MDbfpc0qYmeOpxvxrGFtCWdNBXDzJPbqhsii8uSu7nyqerAUW8czXOopeWBH
ZcXFYWzZd0Cj3U55uJ+5hDHH3xJsKaC/0Lrdpq7wTfwIQNliy6h55yrxWNKP
mCsUoEyWWfn5K86Im2nJWN0AoILqlQQ0nJeji4FZ2xdDj5vNm1168WiIZqi6
2l5YUomCmjreq9clxWg48mYkh+ToQxnkVsNzFJpMl6JlMsi9766MUwBYTMu4
cK+19ffdAAb7cH8SVfSFGpOEjR8oqDqwDIhHIsVAzHol2CATlrLWCJWmGzNW
urMqISODJop3Ik+4uQ+bDTAvOlSdvLhYnDBZftMab+Q7BiJBmRmkMoHVQR8y
OfIjcdTRRcTYb0FWVB+uErCZ39psrHeYi80WY+Ta3sMyqmlA8sNcSeN9JWmY
+RGabccHaQly5ncuOwC9YyEsW4w9rBnngYMmDIe9V0mtaliDrYhzlvCpzAWv
ruUhCjWZkw7RbpbjggqzT6gntJJpkUrRN2+n6WWXI+p4GPL5JVBiXbF5O9wC
PKQFmUAFNLVgsKO2veq2JyRq84P7jSoiig5G2TpYWR9/r3+tZ52Xl6Z0BFsD
hEfohqdpUv8o2n3lTimol3Ql2ezZJkKEAhVT3Yu9rDykw4OXREHVexoo2HMh
uQMd+A7lNlw4XSrfDLZx22meII0sew1FZM7flw5Is8pR+flfMaE2eRAkrC6P
/NaxZVbWOQwyLRzkDfLXpw2R3OAoveW6RiAeRI5V7qUVgRGSRZaM+1bHiegm
AML5Y6CX0zoxfTF9AGR0XdT5iwrmVRz9eCDTeIp153ZsJ25djWWoK1AZxmE/
9mLQMw2BMcP6HoSIlY9L8DLSKyDmG0mWQ6yF1RrvjnoLIRDc1pUyYzw0N0tp
bLT9jmMYnq3mo4KTWOT2RHB0JLo5t6ty1fjAw525stBiOwPSHy7U/Ir+tZBP
z+ibyFzEY4PxgmR2CKB7rXSGPDfDOgey2l7MERNQ/PoBZXBdHODBxxBrCO32
6xmtq/cH+GR1JlpU79VLjX42ciXCQ+JNW816G9RZA6wPxPO8fTNrZewIoDRs
oUZRvfHZrndMkxrJ6BOx7Vv0EMBbLPIrKQ43OiPJHk1vHTt0QSnqqPsB3bCU
CZ8+V9AsELAAnD2Bw5NVHNOYwbKs3ElRe71AJB9llchr2ys1CkZRz2j0xByX
/t+92QXGLcUplroZskZ2KphdTpeD7kesUK3hQhU9VM51BKLlW2QndFdpWaJE
OzmgSZZGGh3QtQ9yBqe9sjP4gNm4OY8SDqLdUL0oFuhNnmlpSVZ5t04x4A0/
US629xlCC0AQOJK/3ti76gCdS4up4VAOEA0mhIjGjpHSPhWsb5Xf7JCCYG2j
fahaYhVQU2toDcFI1kBIcKc/ZINghwg37KhVp1UNj4LSIEEoNfPQfuRTYi7n
1UW640AP0cN87wE+eYmTFhYXW0B++gJgViEdPEcqff1eWLP05ky7D6mqq7MZ
w/YzsdCW8x1HJs+yPM4GTJPt81aQTgSYlEJi1cSF1AgVt4RCd1Bi3Vya/2ey
Z3/c74peeLTV1qdFcpg1VeXQu4fcaVHZIOnZHWA+g7jgNDj6YRVL7LKgTpCw
q6Ert7gbmzfVf9+Cbz2e5xAhPOoDgzQL8vFY20fw8ug0teJ1n5TBOIcs5i9T
cTsCNg6w1k/0S2cJ9QonH+VZq0mtYXtHQwPgsrmZZeTffXCDRgFAIZCWVQTT
i+TnqoIDx6xDW/c/aELvu1/NcfrlkrS98jHkpiR22yO0HCWBmqUHEL4d5Pg4
NcEsPnj7M7ti8S2kUyW5Vu5bp8BAqt6f99B5LAzbOgePErWK9AFlR5sB4xsU
rKwqIXW9Yc6sqy5C7AwvrIHYEuOghJZyw0AF87hG9HUYbW4dvmWaCRZvoeof
O3Sp65kZkBh31adN8ik+9gMRmPd3fsrQqJWdSEnP12/kKywON9QX+SXFRu4v
+feU0Z0dcLeD1wGLO14cSujbIjPaYVKaa023PSdTjy6aijCPUpUQ8zWThTLM
7eZzwrQM1USwbsxemOs5qPQ/a1pRnVVVybljvxQzDDG4ahf7ufUhCYppGtbJ
8gKLFrPZQoVmoIXeiDgq9ZKP0cHXeqDbkjWwH38E+Hp9CghJjVR5lkTky9fW
pXIYyZ7Pxlv8Ru5x8XSsraa0F4c6YcgTvZ3nsPipzyskDljbCtoILQU7sWfT
/fgY5zPRMkJsVag7veZqoFuNTUUe03ez9gZR/ofNKlQE8Z21gIIlY36K6mZu
3G2NXQGPlWlLlQebCBb9HyYxp2wmYsmvLyM/0kSstcCbZtWn25ScIxsiRbTD
UwAjUXmxmo8MqPC66JUMvWXD265QnYFPDe/SoemutSsR5r9CR3JkCY8Icsw0
FxUzTNIFRKublkAg3WfIpc/cK4DagGQ7JEEx96j5QjtkhGJTdG57wK7KTF2S
B014Pt1lzID7xod830GA9fziGCGYScwW+rpN0Htjk9niagUWHMcrpfgedhnY
hqfphG0lPSSAGMTU3EHBFqYMPEhhsFCga0f53FXmBk6fbEg/KN9cwRAr+avu
3+vvjHwr13zt8VB4yRnW8ig8SQBkwIoxRH7brpKv8duwkoG9GoqA0bP3HhOj
ZHPHmlBKdmdkKYRvj7ddw2C+rKuHa1mYDgTG+aO6mqJvCk1j6WKIauHyoEla
DHnv+s6GEiY4oHmnFkg8foCgGDSOG1lZuLgimcfnTs5nKtunZw1rysiuImw1
3njyzyuDRVyHwZEqhPbkJ4NLOgku9kOb24PVLOdvxjZOa0XO7HCkdseJrx3B
PpvqmQUY1O4l+h1Zif19R/JMp4UamhQfpQ+Nim3NrtNxGFuAIlOVOuO9S82b
N1nF1ZXZNE0ASZMrghOjTsgxlNNtmJuGHito+uXOrd+uEY0k/RZIAgXKqt8c
M09NHEI2GRd4abIRHHWl2DfYw1HulKZcv+OOQMA08riMcGvM1JIoAF7ULT19
zlamEpql+ieH+c3SvkjUOngrsyDKr4BmN8h6p51+ob9ZQce/q/g/zAHSWxnK
PZohfomHDuucZZPpzLkuMspLxePZtYra8Gj6T/6StypgeUs82kgVnwdb63pj
18Le/e1RQXVd81SNSSYkrCdPMAlH/atVhwXI8O2X8o+oCGbNlGPjmaPzP2Dh
/V2HRMLxaBKAFSFdtCnPEDRElFSMDpCI6nVq60vNS+hVXukD3IZhJEY4tGsY
/IPRpRxesFgKnQAbXmtEs3yoix3t0CAL3PLLLj+jYT28Jw8oz1XTYiaws98U
MeXV494yWxNxyYMu56j/gBvecxYjC7DApRfS47dpl2hzkLemvANaWih6nc6w
RVPWUC5r2Mekbs9uUStsDqqiWEHjAPK7Xk6DFKnPycVgpcCBM2ZW0+I55/qi
7bbhwokV615jXE59tDvo61RahSiDaAtW2+Uo/BOAD3Esxy5WH4eo8mGX4pfk
fFaBu2PjwWyKabogeHDS7LSxjqN2MXUgthubdEKXp2biu7Y23Q21/8ZDSXyI
rlH4/+bxINGRRq/kZ5C9++TXbKmij63un593jT9o2vx1UCJTZs1DJACGYi/P
ZPji7o5XYm210i7y/l1dYJpSy1msnzNTcYwJOHFOUQfd9/m21KRRnHBO+QBp
eD8HlHToeGI0yFWkhKKciCws56xFF5RMvneeBWwfK+i9399J4IEh7cV6siPZ
Z8rOwGAOCU4KfvqNAMUqxmIWK007rWCrTYxt2cCcndbuJ12wc2f6gBJaOsGi
pZKK1C/eUvxsn9RWk0EL8vC5WC1m9ZHxfX2uNeJYRTcEYV8hg+OIUHGvAdQJ
eB93lJYxjYL5bfxQ1ES6gMtv7rKuhub20GQs3LXUy3VcpKtkoKHs/fjlj9j8
iHSzfbyf3U5D1u4K7SaJhQK24ai16fVfI5HHcCiK7OPD8AG/7HG9InBHjbOL
sEKBPUc2qVyCNGrukS+T8WGFAVyBre1/GlCRFRFnhdWW8iJXt2DbUv46BXrP
jZJsnjS5gouVolci0CM/pJnlKXRnqj1Jhud1pjBUkoaNWe+GOc0KQd8hZPuD
R8zJTO/4qZ+O+45cRLIlCN7FEQ37nzBSoPpUMpKRCFWkJ30fQnq6s+i+DvSh
sVIH4MQGnEHnslcem6cFlpqiwtLrZ61KX/AbEwOcwvQuGVdVAKSPGl/u3wRs
1cWuokfnY+F54W+TockT/Icl7iJ4JnWA3vmKTaOAAispj3EyYa9zAEzofe2p
7z01a0txI0reoB2L1HMyhCv+A4KlTO/dmQLfLUkiVWPRijIPhn5ulT6XXujg
Rc6UzkPDWBWW+CHSJHvvF1AAseMiutae3UFz005p/xUiP1xu50QdBCZOrLFy
63kvVPFmKNliTxmCF4n2m4FL5hYcZY1gbD9YWNfyVl3aFxNU0yG9HQrS1rtV
u/Bu9gkW5vocY6frKbdVN9EKHOSBCKIMmyNnGdBqxK+sCc4SU1XsH/C8RMFG
WINQejC8TgnQyhmfG6q5Mb1NdssqNTlrsjBtCVRERzL0kuDjfeMRnnnhYo/f
h58RG6P+ZNyx4vxvYApKYuweJE8K15FgxeX4Uf1NH0Y5hOAvHD+1sUKnIrT1
5Qy3zq39acZzk7AgDpBNodUad7gJv4v70uZDhu8zZuvx8DDdJvZyNOUVjkRo
VUn08La8hWIaWn1wA1KCZTITwWieciXzn6Xk/HbJx10HXiSMIXlgQFOOfSEc
mKTCuY3l1sGtJX/0x0AljOa4cVdaAw40f5u30qqTFSFkFuWWnD2YHq1A06B/
XmCTydGWR2TnduWQIj7GRqusQJ8BbWCfYcVBkupUBxWoEhtawr6Jf9Gn5Pl1
UXlTtYW+I+Ouji68+oHru++kKlcCBzfvsmQ61A6xNz0rjzhll8mZDBMoCaIs
VH/eGWaFJRI6RLjnDG66kqOMxWgPWwM5yZcyVgYQnGMy5Cru8A4/VV2pcDwq
tP9OeZLuGZ/9DPJtLYKy4yNA5qeYj8JY5djbINn8Rxt04awA8+FSgJF1Ei5z
qzGWNQTCVZ1fMCCT6B3ePIVjJ6b7HnjpFQXA1GPPCjI50sHQhonUzPs23KFW
SDJ6SnxrZnNvstgXdLyaRYBTDxXyR6MU3xx2uLRfLxUVtoi24RYrkHKqvIXy
jtAKP48F1j2i4PSIjeox6AhytHhmrJcwgELJmUkb9d3RtQLkbh0YPldeasR5
XKbtyetzy97n+F6LycGWTyPKIZ+dfrLr+gL52GAUfS6gO5pNKHhGB+/QaEsF
lAoyTufYGYTzhg93kTl6FXBEPVmYETBi/ePaR88tJVxow3E27Q6PE4MBUtyx
2/hkSibdrIoQkYJ2aqVIDWkLtn/zKkbyHKNZpeQcKL7eLyXb+h1Yff/QwWza
UXoqQlGy5nj8IIDVHiqDRcJnYB8VdK5CIm9qsAtHQjJ4xnE9O5qTSfd0p6yk
vz5461E5kbJzTEVqN2NuUCDX+xx0LC05OOHrkIGweT0HsnNCepx8gT8uiaf1
xSWpypLgBuiPiP0tOJhrmlnDC9J9gn6uN7XPU0Ebe3YhuIa5Z/Zpsom9g9Yh
xijFST+zjR5n/o+dE0arhiI43jU+oLTEiHBYayKxfN2wyGGvAleoWOFIDKvA
+U+0hyyl++Df5m5fj5ERpDhRqDNOwSFwn2gWN/zS/tgWqLD0lIleNScI1qxp
0FRq9jx96lT4+j7YC7nS5tY8EjkN9FbTHtzBARLO88O163CwA8HJtRPGWo+y
AlfD+U7G05aA/3JtB6hBy/4zvFKTbx1NCKpBfjFX5DFlQqBlW71FNCK0mqbT
O+eLUkaRXWQJJm736wXb9AXoKa3YL1srb2oMUqk+m2sL0tELis1RxXOBrxMt
OBDEl6CqEJmh+NjEmsEqfrNHeuGMpyirLQ4pbXUwvJTbWalMRoUylZkYn3Hb
Hi9uAXF1HvKWCGAKoMRamg5jDEhxlYWgZtBuv648ccve/qEpFB2Io9rRQNZG
WatvTsV+Ss2nbuooz9erHvJRCr+IsLNEB1reZs1vLt+ebFYFkJTGUuF609Y1
uVGp3mXC5O+a5f/qgYx8m0wE0lsgecmbo7uRvfSgPGpAca6FQuoK2c12hN9W
MSbmwRNsp9U3y9XpOg9nHUZFPrCRBuP7HR53Zsih/xcaP4/VcX0Mg7vaT9gw
JdAfyuyW2sG3vbs4Hx130/puEWrT+2tEXkGBjmZwbhaJF5Vtg4kmcBJxUZG0
aQnS9XHCpwPkXR0M4UiU9MdyBrE0SA5inNcvi/RhB5re/nIIbFeK6INE8AIU
oVTN0BlYve+2SlAvO1jzQpzEM46pdX6o5L9vPmhBAMVqKAIWyvCuFnqoSTk2
dTXiqwdjq+p5YSJor0+RAafg2kfLZUT3YZLi+1yGZDK3XtHhxiTtTcKtfZRL
dSlHnltLOIrR/re3LXwcgUpZ1HLkISlDhZ1e6ySn6PhHy3sElCR5b4m3KEcg
WxovP0zGOAPWNJbujGKH4n9IoqomD4V9DIQkystYXD01ThNFYo0OJPKpITMR
bLfoswRiPBFNHg/LL7moE6SkCky8j7n9FlYtUDys9JuJxjfwj0cV+LTW/LQt
nJEce2r8kWAfxnulxZrlQx569XkanWJJ7gZ/Xtn1ZRXwqxG/rWRXGj+71xSp
vYtpQ0HvReXy5HusPxlz57afG949a7wbUyw28pr9xxYAtQqH5Tn/4yAoPDw7
bgOic2NWiaXN61YdD95F2/wE4uKiUVDqz9kg+EVRM5EunWkImjSGgff+God5
HoBxn6VedSHOwW0+/XXVuuitF/QGebnlh2TlnQxTQQO5pQlfiIg5RevRPb/u
95kK04C70vqK3/tt+03HBaELv1bhFFhOLJNqJxqBBr0R53eloTzjUA+QoLeM
SAo11zNVlbD65n6dxKBscMHf92+O/UKoVSVXlhADiEBJoggsbLobgHIYggTJ
Jy9cPzu5a5wLKEhCdYEgJCx+kF+EvpSlS4wWjq0AzAZKoExGCQatKfGyh53g
jWWpZKVBYUJq5mYibVFM3sjIjWMwWuTq2J5FjqGS8zM6gzIcYNyLYnLUd5tL
031DCy/NB4DQMIf8NfSZDf69id/Qud8PUaXaBo/AdWw0GqRMljOZ9e9aem0h
GiOzcDzJAphwrXG43N8t2bgntk/zunTopvgqDlpeUOe2fFVGz16EToXduoxk
ChEyqplBOKv0LcH/hHOzgZblBtsJ+K5ets+a9UqcErpWNontqO9VW4ucDxV8
uFsEO2eAqoHqlYXg9lXNRADngxlOPRBwdlwI4tGUY52i2cQ7RdLzMXhoXdpj
iE237NQOrsL0kaek+z/xY6u3hjNK1CrtsUELv0HaMC4xpDNCFABDl+I0VHV8
isDJbInNa0KsroCcOOn4e2M7zR9yheAaniD+Tpg4pY+Ein06Kwg8MS4fveAo
q9pv2GSGhIEYmLJRdwyPb6VpqqWSiXIRGuaat8w5/euWeV+qfGZku+lmCwc9
KVJeiX2dzb/U2G5akfF32SRUU8bpvMMlCQp5CYfiFVRAQwINFkjxS4qV+NwV
JAbdxWlaWJLlWimy69uKROTCcO8ikCjTZERBrwOxwYVnj1K7GnWOrR9s30HS
qljgXNq+lXQfzB00inpB1YPNM+bh2rGCNuqkarzA1DU4BG7GaQdsQdYRWaoe
3E8McNU1Dn0KUahtCbntjm2DKJUWxytpecJ4o+qFI3Tbd7uEru5LcOmdj8v3
rlZeDoG+SRE/OVSJaAU2+v7Z552C0/75nj8Pi42C/3ngksSdN3yhYbdSB/fe
aeYnBwer2nKP+mU+PKKwydc1nU9mqIAQk+d5z6aKYDa4WGvCL3xOjBExha0p
ETzbxTYNz5KEJJx+aK3IEXG4vl07Y3pzuQlE7PlgsTxwpIQI4hRDMNKTdy/c
Uwpetgv8UhxN+JyQtYZ8FrK/ghwXC6gwzKEBGQD14Kw8x5kcSq2UN6cmzsyT
XLrrgdtHxqPjmcvDPmbuBt+PkRCSUoa6dHk8mIyJcaVHYBv4mmFJpWZxQi39
PuzZk/7itSwgIXQjo1xofV8lBJ9EbLT2q+Tyd+5LnwXwm0UU3DanmcXE2R5Z
FeticpvWoZTFgLuw77Ue3jvlJ18Enl7xXbG6dlh+uTUkiczRm3PhwwAlSnFd
s23GsCd7islQ0VOspuwdwF2ezlf1C+1MxjcYCSC5Rr0Aevz1mzvmBGdaEZFa
IuAoEa+HEPOjmoyvbjyA41HUCRwjvUbyvkLX8GAraE9rArmMxnkd6nta2MFo
VZyHCVllcPoctIFZRuWBX+xw6YgCuaem9GqYumP2CtibL/1zO112oL4ZPHUu
B58ivl4UxzO8Qap6tJdqNCLAChx+FckvNJ27qPwwY8tnZ0/PwEaY1XpKMRsA
8bpCf6kLjV3QgvRu6MxdTB4ZnoQ/607/Xl0mD84O3idi3ZFyTDir64lcoJvS
4mgZNHpiPPQ3wrsL/dFaT+oj8/LvzaOTNWKTUEfkmur6EwIx/1chkzRi3F0D
z1J81ibsRjqxXmZ0gEOxj7gsIQzCcCfUUfJ2C3AlynaQw2gY6kr7Nu8vcscV
CGoMNJA8wYLpgOOTMAQw+XGQe+j0Eh3Yiy6YY5f/D0vMwM+L9CTvO0Sv89Ur
h+axgahdXr4YTMFcWY9K1Ky0D8O+mU4G5Zrfyy0d+Bdw24sAADdN+NFtcTZ1
Lp5ur8cM4Hkk0q4kdR5oS8iLbC2dl4S0YFWfHvZ1m1EqY3Q1QMmzqG+F+JIF
FcWVwJR14+n8mro1VSSVkijKuc1IKQW+1nKO2R/5pTutK7dCiYtrsD+j7AMb
6E3CC2IHIdDxczfyNjn9YAo4gT62h2/EXLkY9aBOWKzQWCiuu0hpQBhp3glI
ce4S0y4yxBWviRIqhTYPnc6yI+B001oNAl4Kb5TcK9ZqGduD+Cx6UTUmIA9X
XD9O9/lXsln25Ykx4TXkcVmW6rZvRBz2CH48w+P+eb2UolgW9TOXZmJwxyHY
0+X/sk/QvY1gKJx5pTVNYagqP3H+qRrFLKW0oCQOQnRWbjCxFVqTleeG8CCu
Tbw70/qTuHppYOauojURazqDdWTqIa2HQku6mO1BfQA8U5MTzrR3fc+kUaGX
oxmTYCFu3ijz1/EcvFQFL3+GlV1+1yBhcY17/BDeDKW9Aqij4FqTINqxbu+h
CMjtOjqdiTt67wxuyljzUHbN87R7K4TGhaSauMyYdbJWunLrwKtxYLEhzNPI
qdqMYNt/zWTrx48ffGScm8U6WMsh+XGOfrkZWOdJVyvJGB4GfRkmaDWNTJQK
/M/5JktvjLF84BDN7NuCG7TV9HDRt7or57w2FodI9ZnIVDxwzn0hKBmOlD8/
ZNybkG8p3QPx8HYVdxaFVHdqdfCd7wl/fg4gDa8WxhTwlvvpUDGzIUNPpzKH
L8YhC2h/+uhH9xtXuWVRvY6RB4guEpQL+k1bCpRgnor33PqyR3OistCopncT
U5WiBixHcupirwsMx6QLyVQVQfr47ohkCM9I+qPQSmvOOe236NXCFpoNAO02
B+u9ahYuqpvnVd3fmJ9Pli6CmP1Zz3SJ1SWLHvVDyXNd+NG73dU4xWHE1eX6
lJ3Ndng9munSnyD/CUO2jJAtMa4vLs2ncA++GM8RYgE7EsyUAiLBNST87Yu8
Z5HWrPWlUENWlO+mds2IiNElxOSB+Sb5YQlWuN3HjaP4GrseM+i/fEcI2l7A
dyHdnINl1+VyWOmgX7/4m5w60iQbESy2ysIuf7ka9XGgw4iOI1T3+0sEHTmv
uj5YrIQkJodCpljaN8pYn5ckoQneJsobNZdoj5t3OlnDo4eX4wwq5ZvqwUV2
ksgr/5TGKVF78OPga3ZJlOTZMQn/aRvNM5yDkkntD31UbYegxr8Vjuzt4qju
V2peYDZ9XUU02IpEYHeGKhalFfOjsX/yF9GOAHFSIfn6vj7Y9NIyufFNHnpm
XgHAq93CENEM1ju5F7MS3ceWnSJjF2zRVEIduNRnb+ujKYB9JuWxUyxFOrOA
/LXbFq41TKH47Sq3j1JmVFTR1cBak6Y+wkvCJ2qdv2abSeQgo+bZi5nfS89Y
lTaZrDC6z9bbHkcnMjI/2WqeLzE5P51RwxGcgGRM5IXvuvxncsqLlNjC5BWS
gTh3RVl1p9OeppLwYYImRW1EOmjU9trzKOOE/ZOkjyfdcBoAf3rzlv0zN9wv
mednhMc47Z43w0uqSluvSf6/j4UwyWXFzv7zFOxfRFnZtXY85yKs8tDI1qn/
H/eAQIpTxJZ4uF7jpCBVcHF3+6cfgTui+DbCq9YrgQigyu0xNffBGbzaG97d
jGRTwzXPDNLbr7HkBjt9jx8rxLjbKr8kGCZeULtUXwDoRSPuPPBV7I2ENejK
Rh3QMrThc6TNXH1XZ0vmiZEeRBImghY0MRkD5asLv2RhD1lao+ESEd6w8DWA
ATnFPLslJv6cdOPxvaNvcdqVARhfczqT3x7fTv3cYYoyFjGaqRN/iCaFRWHy
7naO53CO4u0OVyzr7ZldPWz4+0wBE0rdhlJE267P1nNgNhrMeBVHVrHq34mF
SlT3beO896XtOhlCucBlwhET99lmF6N1EeeeMM+JUEztHhV+ud4s0/eNgrf2
/SWXt9WLbbaKs5qPBeb+97HneU4fihErL8ChyD/O3AvKxutI/nuYdnI/5DKg
meyw8wEDTopIl9IZX6pjdpAaVTR6uF1Y/k5jVJjZN1T6+WWWU+eMbHDzVqSN
vNc5QSI3Magcfkd602+PSpYynqyB049Q9DmGLF0SjGsHA0QWbrDrDUeqf3uP
6Qxs9e1v3yMhKUlTmP8vGRwXznP99pNSF5cEb/6anuzoZc0y2gEP0r9rVUom
fQFO8+yKARMZpzD19XPb8e2VfYYSwYI89+g5ee6WkD9eTu2RXsPuFKCDbj/o
MRz3rLxjDyTiI7sLWoT4wMC/hh0Fxf/xiztUTa0fCNFEgRZzqbc8Ku4kOIYL
Mok29/O1Ugf6vr3pIi+iq/dcdtyMFHH8pnC2gfM3cywJ35g+Z4pW07ao2CrN
R8Bbi7RTqDcMfvKWZH5oFyKqpy5IpuWDbkFFdzOqFc2agR07yo49cOg6WqVS
fhVmiMEqqenTDCBn+FJVMJcsljA9Yn/D0q9chn69Vlg5ibqt1Sgi1XzphjoX
fD0aj9qzag0Fg5+peZJNa36MGH7X/Lx1xXiTIB0xhSMvxJ2KtxCNMCgKB67Y
bJOu3PlZi2lLr/uYU1OjpVU7ySaIU3KitCyHbV/4EiTCT/rH1sz0HH6n0tW/
UC46if2Rl9X3idk624X0RzXf7hKozQcA0Jnve8X1BpX/ojjNuQ0eWv0X2AOw
c0mEICh/6EsfGHeITFeSa9C9F8cIyDC3F4gV/HFpD9G8sr8kaXF3G7Qg2co7
McPLmsubZUFx+YzJuIIUt325g8tMrsbEREoh/OQsSWqhFJFR0mugNXOh1LX4
BsagrewSsOo+zPXrFncxVYKprU0r3cMU/wWc4QfLQWyvLpu/2lDP0Y1/nu9d
E5W5vI8mbpZPw8G4+0p7FacO7KMdVKd5Y48VLqtdtK7iCxmB/8z2sSpM7VKz
v4MXSo7MRJ7Cx8JFwnttuRB9Y2Ln3+9s5KKbmrYl7uYX31eKFldhEg/eRjm5
DSh0O6LZ4D63OiHVxdd58WPS7bZ0v6xCkNwjc/wUZjJgEfIeL1iseL5AykkK
tGBa8qXCqjniJs5Ot9RCgwWGjPDnppBGOpVh16x7mIvPRjXLPn8VXenDFDKr
+aVz7g5hSsFU3WKxdug0O6aEMdeONSjayTipDcO1brn2m8feUI9YprreeDft
B3/8w9qwpJiL3LuEKcWP7SYZxeGXtN1c1MQxgoGrqmuRWhN+WTrpGddpWQvF
sEEot7cvEKmctRL7lg7hfmmSLudnPabz6E6CjFI06feO/iIo1MvLMUciV5G3
qDFkjheRSsKD1J7ExatkW3PBUvaUvqkbrTJmMo2PcEsa2SBWh2kORVFaWyp5
AcPt+LjF3C4izQ8jFmazO/vzwCACoSDKa9uYz1BGb+vmKScrAo3c44qNzl13
7l07vXrITS+zWXaYDjNCRK5Vb/EiAiMi5r1jHzxRdDild5a7J7xjVA3CZ3E+
oYNRqI6LI8x/fbN//MDxv7C3R/ZMjJqpmgSQ+rhmd6fm6n77gFM//6wuBg9d
eslpbRVtLcCt4bneW2X70sZFLISyCuQTUOrIQQ3nZ0fXthQ6HxEF1L/QnMmX
yrxvrlIYs/CEKm5iI9Zwpz2imy6dTSzQisOmU/kte6Cjdb09l/5EEOggoH23
NvtLdxrgtwpeNPoRbJxQlKocwRQN9S8VZFwDySt09B/zxt5CXCTPmHAAadP4
wjcPz9HmgBVLo3RrPhXtutFpQonSR4iMnxQr5twp4mRRyfoxMe2+Mosw7yLV
pLF6EloY/j02Oh+RYUtoniQOIATNE4Ej01cwGClQiLDa4VVPQpdHJIH8Nocb
B8R2hIfyYb+ErbKSUFO53TC5Lpst9ZHkpbKaHs35LuhfsZzjkqkdpjQ3H1iA
/KA5OiUhbM0phbhXG8hduN9NQeeQv1hmolX/+hINzHRCNPK+ZcAuDpNwjk9m
9ZG4uhXMlO4QK/VJQXLFo/FibqV/5nAprPNTO8n8SjUFzJD0IBHr97frLNlz
pirdaNmAQw0LBqzCQS34eWKCrLePPAHTcRNlROXAe4q+M1yNn0SvWmuNAIct
o0603VlwAR23NPLfkayB7cUS0G9T9ZS2juUkWcW8h0EV1uzPK2Svjx+OThax
CdgvWQJzM8s6CqiPkVWiBf+h3zQD5i91s8xAM/1tCe6e8T0Qs5xZyKlcYcmw
tWJ/eddkW7zE5bSxrMserJVQtLJgAcqlgTlGbOuqeyMvtPtq3usERDzWEt9Q
4xF6bdEI/peO0Hb/onA+Gp0uWlJPjOBBFJgml7McsdEFQEMj684HudggdSUi
URcTBoc/MMv+130I+8CA6qYQB6YV2kxPuct6PP0XL+qiQvW5xOJY216ay1W0
DYDYYmHENU+QtORJkofn9Fu9bw5GIG6ZwYtyqgcc68FPP839AgOX9hat+fpb
PqybIAZtZwoD3LAizMLhQryRjcVHHpOjspXbVwbWsYW7YZNMG4Zu1b1L0L77
UjJkAAPbsG83CSzCaodl0I/jOZxWIKsf+l+OulsNGSomkCEypSrt5q6BKRz+
g2SYZy5Pn2tYsOfpV6PlTQz8W9+qFptuDl3MK6yNBoAPXh+s46RbgzavWPXW
Q8ThhwGwqa/5qLwCck+gY+YBteig83pMcYph9hQV1yaCUV5wYXJq4FsZN3f7
Bvg/l1JEB5IMVWHZQlxpLbWpuEBPS8NxxYo++Fmt64J7SWeqoI+b0WOi5P+J
rg8GUUt8SAtCFNTW8tdgwSl0yC+2pP2obrwbjyKUUxK2lq2C9DnaQ7bFef5C
oUy/zOje/pf4J+atta4RJbd99LJX4UjKq7Tcpx6qY9ovJgObbSvzm/CQ77fk
nSvZ43w3H6EnA1bv96Poied4T6UclEB4tJO188U+8dUQCztNGYtRxPt5dx7s
z/LhYHR0cBCtfEieaUxYzZW5Pm7YAmhjmwRx+aaYrmO22+1RAijMZ8JoFFBb
AKDrrKWEQlpzKNepDWvc3Pp6Hh2C9gs5/ngz9F3o6il3toB+mu83+A48Lrns
07pWqpp3FHiD7qj7Xv5mZFj/QcczFvN5eIDEbomQn/xoamgsd/rnh3tJSz6s
vJ64uyKW9B4NIfXU1j3oXV9tzzjBTZf7vk7IK7j3LxT5YiSUuh5OsF0ZlhS4
CsuDh6fIzOywgFxwwn0rYYjebxHQB8bpHT+LULCdfvy1tpXefWvOp3pW+MXf
ilE+5iavLkC+HrUwD0tokh8tymIIlkcrdeokVVrsl+xjVeLkeKE0zsLNn5HG
loVti8BDFdEfBwipkrf4BIFXmUkTjVgDnPvaiZ+AwPmLWJvxF0aYR5eohfop
dSFKmx2K/DxAalWv9TwmRhfdNscIvX+dC/8Tj3MCWAULdZXydqj9Y+xCZhkh
x6KyXGIpwzMUlAglQNNb7bFm5AU4XxFuw3ReUJXVwxAbO5vR+jcN2FHaS93S
JHecdNfTNt9XmUCawvzFiL6EIybawNRtCZGJGO1CJ86OoiRjaJiLzolLhRdc
ppi8E2T8BLNl2zH1p0KUF4o/cp0/NSZJGvp9b4M9pyuU+LcTrvR8OPJ6Q98A
8+5QOVfMMR31R4ep/yoK2ektfGZ/eb4KuPmQ5jEceQxbNcvayDX2GXnFdYLN
xd13vPttzYufa+XWP7m0OeTh+e8Yst8ZDwrDiCqVZlRy/+Jxs5S7VnlBS7Zv
zOvLz3gYLHQbXoJ2SewvNhwWFmcKP7ik+evmIBEwTO8lJ8OAZDrP7z9Jsl5A
KvDqV1YkfYrs3P0L7cuBXwi5r2Iht8euDSGdrMj0n1/zeL4mGtmybCrg1SuO
p8LXetp6000PZ0ymg5qP2j56Osiq7BlAp2btU653wiyyaxK0PnA2h8Lyr4iz
efd4JMaNB7xLeFN1cJcCDREo/7ZAlTuft6YPylPLW8ojbk6cV4f+bcbvRMTs
nOSzl5UhItgqoh8nQClUJPQg2kI5WiiNLPupZMnyOSXttmMHn9LYdQmiTfOF
R2QNger5LFeoJ9fMIBOFUGWz++fnZbj4SUk52P6DQRuMiy+NCYthoG0Nr7tf
0lZHmZ2c+27jciOQeuG1bSKFTtxrj1LYeEnJmTpvm/8hJExQNay7UbqKnMs+
uXPT6h4W1QGwT1cSwC6Irh3Wg+GzCbjlwmx6l6kQ3XTtIFOwunTKg8oqhgg3
xU0DBQwZsLl747sIubp0x1/QskjgrgCWILsg/tu9wOCnWgskhpZmbRAPSuTv
hNSkfyRV9gbxlf1IFXtxBfTAL7Imdgv8E9GS5pUpymRcz1JjIiA6+0u+g2vU
LkQp7gLNoqXrK4bLloqT/Bub+6kb8FctFDOOemWl7JbHIj2CpqkhNSqerx6h
kmHTKVtir2oH+MoqQORcdC2Cm91OpHLUMJwWoXRIsY6a1hJwaIl+RzEW9wi9
I96cT1iMvPmmwqbOYM19wZOmXo+W4VI5gOMKHFRGtGvNfbx1Bzidpm2wOfE8
/5vVxix4KVkyrgaMkBfiy/vK1xnjaXzh1+lLoqm65zjkaVex8P0O0ckRHo9T
QD4dF3SGs/D6iB2z+xzfINqrpiYyC12Eu6YkpR4GgdBzEi2rO+92igjka7od
guWALndEqtXESiAh68DRFPTFRG6Fd2ya8+r1z8k7ME2XOy9CZdwqbl5A1ifz
OCpxJ2mfWGN3D3LR4gLdrlhYa6K0+ApBapymDmEdAnOHv/0o5FGvsTZysT33
56zAr9uODGhYHxT23xIYyoJLx7zRuzcv5u8SnjjPHIi8aH6R1Obb78hLGLcj
lnxt2zg0V5nCcInupwoT4vRqq1XAWuk/csYOjgIiwomp3WC3NIQrc95uXuWn
e3itBrefcUi1gUJ/sYrg4zUcxFsgz/DI90MFVcL2g7Cq0bB9Cz/kBaN1meg2
Mo17glvpCh98GFJEXNlaNNGEZ/V4df4c2Y/JRNRxYdNQA4RgMy0GvyOmpd7e
t9eK456AYZB15ORXHVdAMmfEpATIuegjEfRiw3SUUa/MpJXVYl7cevikekBw
SYmnz6ORJKsT2HzdeG8CXc05VZ2t+Y6B+2iDLwAaPJ8M31xb63gdF/HIZRhZ
tQjQZ/DzpaXQUDZ2XMvHqYNv21XTo/2BLhcuvIav1WqjVzj6nU5wzsH3zXR4
n+tt7IEc9jj0RNu9XeyCcGnCPOnEqnXiBg0hq24LiCSvuJx11mrljTG1hosG
MavchJyFil4g2HpXjnG1dg0Hil3GSeO7uK4JV5V0XRlaINcA5ZYnZvdgeS9O
ClqUvRezh8fDOTjMRNuQBMDqcuR3kVEWLGPYD+E0gvaDiQ/fiMyNQK4Q83hX
B8N3NBQCvVFXppFhJaTjV8fi1/F4lc4RNHnvRI5y1kDu1Hhu0IfP3TCRn+Ef
lT97ucmkv4GC11ynwRN3MzRMPpOYk/I37REuKM1N5mk5+pE1w548xUIY/KNo
XOcl7rz2GzEG1g7wllNGYmtu7cVLBD28smtzD+KD/XQ9FWHpwGwvN9B46k8Z
gx7/tvWeR2FnogTEXqODCQD3x2Q2IszHr5psJJ5Q34eJqt8hkCVRW5+NSN1t
3hGwv9eEKdiHiyZp5eMNZnxe2TspxPVGrNJamJ/lsr15mc4YPAkVP7kLB3Xi
+XgLpx6a/FLPDcRuO1TsCLZhAyNATTZh73WhGwjPRTcb1L4YC5P9alraYEnN
lRUx9XznDBBapYrNMM19SWdDHNYhOBS1Nfv2nDUBzOHfxbafUOTAb8XCFSC3
mdY7CIIPU0WYyDA6fKw6WKP40/boIcOh1oZZNNFUqFLb7MDwhq9IL/bYkpn/
f1x/aLb56PdTfL7PcolAhr856TUNJgVMIlaZy0vdGnKN/NX9XnS5OSwh9UuW
uqUhkvByiekktLw8bKXJy6txZrc29wPJXdANPa0qAbnBfAIa/L1NzjsfltgW
TbhMZfydQdbWsLQGULbVLMk53N/+XaUops/C9NKb30Nuca0lhoT7Kdn7VjWg
yDQbdJTrPLlPvfxhDtTT7kM6BjgCE2ZvhapSYNUgMzW2H8OHkOrGTv1WufSk
VMosJUcE0vm8cQL52q0PIK9x3HtmG++d8UXOfe+5z+EMoz6CA7ucm+bRBQOt
gp3HDTuiHY5L/kmRHtJcFS3tVzwtRw710wbqMQP4vQ51wZxV6sorJTPpWBgE
XeusAWr+EiYKvhnFNNKsiHPxaX3sflhAp//XgSp/oBDeCghYIM4ZNwVW+vWr
zCQC5PW1nsdkJFTu0I2Km+IHe0yUyonv84u9Wh15VPh1SLzSIrNVvo8I+DXk
6MlSTJ4QGV0lspDfMvgAdnsk1z9biQzTq/2ydG4czbvBrR4ofrHEn6W/fvvT
sFApFQm1jNq05lBgKGWdx+uAFU90YRXjUMF3qrl4OoiWKWPpruJRaQjACu3O
3jpAm8OGSCMM9Jqw2gYRq1Xv4tZ1eBhis4YFGG9rXBOkFLxr4/N+OgxFfCUb
xCw7+GQwF6lfglc1Y4aukbUkxlNWAD4u4EjGvGTNnbr1uDHcQRUVYnsr8c4s
DLTSIWNtSQeMPuVvph+9NgJCisA8lJBinbpBWYtwk4zaLtyup2ZZMczCk7lq
f0gd0b6m0d7us6k+05UF5Dw4wSi/Jvxm+GR+8Ba0X1T254TFJIMtqhyG5XLu
ScXAVvD1Dw6haVMJr+8y6uwab/lXMaYjyNxOasH9vn0xZthdVXKTifcett4h
2p+CAfabos1kgL995xyTQKjJw3nLdnRIsP/R3nq9MZeFfUoUMGkyJft7QBg+
pL00wuuYNxefpjTNYjNx4LwQ1vfE1GbaRwqLan7YtFLotICcrKnHANHR5XDT
wYGMLmCLM/Xm3PVHa/GJgcY7/uaaLKwTcBEWARksM2U8bqRZVaX8TfWBs1D/
dTZWSaJSFvNaJwr9styyea2R5s6CJY9D6Bcaw0Hbh0jZW+E+QB51EruouXGE
BMrEgQjTTonZGLxjxHYUpQPDrJH3FgFIproGUiUC0Z13s1jEBJSM+8H130Lc
uhza1HJ+WeRcaJcInDS7H/268GrGDuiOHaqFV9gdTvSv4M+TFxK7GfeNy/gx
25M47isiGZHGVZeJ5DRMccDDQT9oH3D1YNjhNuTox7xZmOys6GoXk+1+9bS2
x6PvEm8M/jDaRVpJy6sb91orueG2H2zeWFpLHiw2VpfIE0yiXMLY41zjtFEK
+7+pOx2hEYa79S8zCTTuKkO7zsLnIchTie2bSTPSEUvIk/ql6aIBeGg0w066
GV/TS4KZeT9ti22fYrCPx04TVOx3cdLJqGFRtI0tO+TE3qB31FQmvZ1neYlg
ES4710Nwuy7ErTOOfG1/y8JpRhPG+Sk1iQweY9Phjl5HGKIig1vcB9micglW
ufPa5eEa6vxToJrMJwf7tY+rG2t3KFk8IomyumtunnOqYQ0m93U9MKLwG+8q
1JUYCFpXDXTPW32ZFWfsDnvTM3o6bbNgNKSjHJOUqAYVqbM0CdcBTs+KYCtT
9yq0Jua/P4+AkrfQA+BMw63lbfYw0bBzEJFGj+Y1kGPrRBV7N7aAT2AgYwPw
wXlsOlXWTorBp9iUj4pJSwc84pjwhS//zriVnATwdznjNtmMmriLQu3hCOvr
Fn4KXSrITSnD47qy1xvcJB37ndJ5jILp9iQ9SQBzlrdPqU/I81ycmuw63f2H
k2z4Gc9q9UUZucTLn+yb0oDA6iDlobN5x4uNX9G0lWW+RcOB0b77XsokOlds
i5NVyZlZsHwO/6Vpp5OFXwwfwLzJDE0alRlQZCAheZihB8ec25CbLCWhMyvP
Z0suhy/XaegDL1+fOM5p0z4b7GQ1V457Au3YlZXD91kofEWjCiMm0Qdgq/VD
ZqEAVnFztEb9hmLs+VF1CSvQDcv1b1DCeXZKlMQ1Sn18xGZLVKZWB5gc5sHd
LWu2ZAM7saD5kJMO1fb1O7PghhPTywnYsI7xb10jqKpc6IxmiVfhAbZErHjQ
Mepl+WbajlL2sfg0kVp/47d1LVOCP5IBArV+1FAQ7K/IHU0Y2ReNGcVB5LbW
u/jaDf9PHyIQzXNLAjBf9RuF4pqXCS6PCdcE6fArS/YgH/98GQPJNa93rZoI
LArRnnbyXf52w/6kuRJqBpv5QvgngdPfc033xeOrSN6pPj8E9HLUeC7cmhs2
G7i6KaeRC/4YqDc856uyVuW6Ukqauum497zwj5x0kUiOfEC43CVaKHl/DYUI
0+MnuktBRE8xmA3/pokjQJxzpsX2AUt4a1oaZWJ8o78IC+taksbF+Kr3B5C7
DHbYUEfBERaCZ/J8ohdht0B911E4FYpyznZ9gbpj23YBuAOiUbUCQv/OxjmZ
7NjdCeQoyPP+MKBnodMCqraE7jWdk+daz0gCOTvHfnDlhwyJGRj3Ye9BV9Fi
aVmZviHC51l4+yivHs1Aj7Y9Z469C2fYfgNjAHpnWcIi8Qspy6i3xpUyTngR
ToHDIJpAppingoOy7szEAzXpOfhmyFtsqIcyd/1cS2EinKNpF6BNSsP/ePeB
Yj0zdOwaAYZT7CIMOQShtHg/byijVOkZWGqSWzXqtnKLKMt+y4lufHfbDe6I
sFn0om9YaHbvbRYpWTKGCuHY4kZLN0oDkXw3HVzisplFY6BaNLw1dPWv86MA
ZFsIcRJtFCSH1v1umY7ZmNJdAC9PbSdVbcA8/inZWyTZdA8VmleJK9brCqyV
PsrgHYt2iY6u5SIu6VcFaC/yTOQbjT4rUrhLLEl3pjPgAqLWvcaVW+L+gFwP
V13LwrIf6oDcCHF8LisVeBjBbWJ0VhUQ3crSDV+EfGsDh072Rro8K77SQcA4
vVqZf8KjdKC0Jx+uLlN6jAw3B46G2B9zChBuZArXi/pHKxYt+WYIED1ofQNU
cTQt7xq7IRq8U7Alms7zO15bW3ICyImfS1owaPfj+0uwqP/mxOyj8YnvnJBN
V3W2SJ2KYbYz7dyFvruFeT8SFa6fMyg1LI0xPZOotJKpXW5ZsquXalpFtvOh
v/ppdv2PnmACqHFEx990D7VbRzFxTucocfYGDeI6jwdCuYnNotQoEgJe9T0L
Sh2UhBnfs9ZXQ1PTOu269p4BfukGrTR0k0V8jK71YMOiRK3z/rp8GfbB3JYp
h3Qu4RQi4arzdeQXMtZnnqFaR+uMAgrD5tJi8YATC8e05Z12SYePtpTREnIC
nHzsOQATCsckCxNCuwYtcRDhg7iioBKZ8cON2V6XZ+PLT4NIO8UNiyXVq1bu
yB/PsrNWl1wifDUx66A6EXNnLoNDGd3OgVPkQovMdK1hAXSgOA5XGS3loi8b
ClgWerW2jigKaggBqMCXLnZIXrs/skQNCI9OKIXTl1TyAWXfQbd4yOAJYMqO
dFbkQbg4cyWt6QsI6whR1dr7/sMXal1C2vRWHvTSIvAvBw6l7Ywk719/yX/g
hHEaKicp3uSeKDvLFYFpckOrt9S81rXe7wRKp3sMcJIIHFCepn2sN3hhEvg9
uqMFEXXKu+Q9MKxdZUf3sZnRDRZ4pmi1RVllsPNC+N6XkF/iHOEnWJ4R3hOB
fccPHFc/By8enO79WnT7St4UR3ME/wqzlCRI9B2DVbyGyUHiVn4Dy8Q13rPe
yDj8H0u2TF7hCoqhYPRD9xSTAvM5cvbfrcep8zRiRqd26K7Q0otZdo7JNIZP
vjhtjdP7GnXHN6I9auQozFFUkTTx5Pj6RZmJxlKqu4qfjaTRNU73Ne2QjY+p
nQQuMhRsyVGU3LH9GuhoiVwPB2CjDPSjtZE2CB8uSR9KoshZsW3Rc/BeAD7d
SgWmSw77ac4yWhpWS83kFAYIdkriJV5X1UcBdCGH1dkQ+y5ceYTiJP3c/ngM
4f0XqwBBQOg6DM78jR7y2OjtxsYect+LznARnQD1eeI1ZKUppETS56H35zcX
8SvW/eAARX/YaLIauNwQ2W4eNQYRGxfkdLgTqH4WfZGapAFQkpUeb9N9SHhr
uL0ZX7fs4ip/wMggf3UgQtuLh7NyRyQoGRHLfp/VXQX1cCrV1HrWi13LO5dG
MSwXvbgnoUHpgYQiv0lmvdehExeWde22WKm3WShHDA77nsjjq5+5TiOmuQEC
wQTu/oL+L2o3vYIDH3GCboMn8DNU87P/pYNWzlGvTKL5BDuv/5TTtnNlxNsd
m2018qubXTHLyACT79BRZG3aGj1vboYJLZNoN9HWuvARRRrm147bWUZ2Fq1p
jJqXL1rpkJ40mIb9c8CcT7MdVdPzeJx1EEQbyLjZtxRfGC3u4f4nflY6db/W
Pr8F5erniLayL7LvImx6yHEpVUizV5StdVWNpAqDzU94GKZJCnWUk7sPMbdv
5hz+O/PXS5fwIsVB2thXe4sV3UIQZsTyJvLYl86fdx0Rm5pTMQiHpqlrcD1c
5YyP1UkWkox1uBrTGna8HCULF0OLN35EVARw7+9wz1QLaiTA863YV254q3As
TMizkelhiLPwX11p342NyRwkWbELIl/Tl1RE94P7SiMywMoT3NbDDRZm/Gpy
O0O8SA2PjmjPI43o617UQYcNt9DrZ8A8YChOxRA/MvNIZQlBSmMaIp6gTXSb
asVmb2/cXEBSJT+M9NfhyzVVB0w/and/gAt19BG6AgmbFD3svRyMqEO6MFam
nYQ69p6yfSiRyLm66PHBBkOugN3WAjRPI5wQsBecYC0QUCKxxE06Ib1QQVEq
Q2GXQvf7H9OR6BQNT+2R0WWT0wJhD8S5yswVsxfgBde4/4Aqle+Vgg/7z62R
cTy9YRn8ebOe/ELeMMzspVJVJ6KIOPFf74lgUlFD4f8tuuCEKN/NXTUKrGvS
8mWV0MDZ7u1ieMkP4S92oRR0x6n4s5CGpsj+8rqJemjXfpIlqBlFdQ+KKq0h
lbgSH7larqPjKsCDTq9CUzhIl1vqrkyLdi9MpgypXahX1A31k9mS2a5jYBx4
qR3SiM/m6e6VlcbYiD7ytvlncjEhN/vcoqDWu+0M9x5K/RyS6n0ZWKCxn68w
SRFduxB1wiWvhn7OrVqdOLvjn9oZTM8i8nt7OYhqMgdjcFKiVoAAQqm+P4A8
bVNUF4Uzt69qebRu1KKkT1jKHRee+em7r4kW+rRYJ2i5xycxwFlmjh3h1p3B
v2eRf3qU6eJslgzG81MEYkS1y3ZxqM+x7xdSzv5QNQmryvEzR7hHRDk8Tucl
OvDhl6o0DFGv+ie3mOAzesJRKxCTMwg37/lg2tsfdQkBQs5A8vMAp/ufHKo6
yp/PbS3L7uuAXVNedqYPxLgt1XNGkbG96lR2P91oAqV3Nr44WDQay3ch6Znp
8xzeUEhaV0iid/YnBHmpr/vHvVJlZtm2+tx+vNf4eS9qWOvzHPsizdq9lsea
w+82xTgplR9ZlyUb/3mvsoMt3p2a6b8Tkf06MgzvFMfIdJw6cQURg46I08es
pyiOXBo9suEz5EA1EjbEjO1qjIEDEUcfxsrY2Unmkx8ugInxGVNVnjzQFhCo
DiamDyqR7B+EKre41FncoidHAiK/f8y3AOzRA9Z3ZDXvYtQOKBY/o1HIfIZP
sN3Kka5UTRVkhBYJMvnw1EOntH/XP3+pgTq57o5MhAdF0JUxbnaE2HTv+d6X
nu6I12jOWHDrf/FWOSAFAMOmkhHoPxRkfmKlgoqwRAQ9G3mT2zsB2WEXlHO9
pVTipkdEx38I45l2YSz9mpADC/GU57OS0pLsP7CI2ChwgFbdmk1d+ujIfeRw
mcsuntdr0i2Ypix3h/jVmxg/h8ctgVMWQ2W4fCSvQdPfgr5mXVyAc3/tG7hc
OWR4CWUGeEpcbsndnFubLV0srgqGT9eduwCznkPoncE6byx+aNSJlBZX2Y2S
lq5meE6trOwLc5rguZy7+IzDShaoC9yUkAFQ4eq12bfG/VmiSZvBWRmy/dNn
e8Z+FG2rIIjituU14yqLeGUyWPe50y61rYFUp2TZW67I3pHtd7bB2zMGQ3W/
5h71D5TjdF3JOo2bHW+WhQU3Q8MSGFJaZK+qzS1vmdIP5gbwEZ0/Me1TdbDj
bK/ARwCj0j5ChKLps6opGOEmR5vo2Bf/m2lSKA9lh8gYXZ3z4D6AgaRSgtSG
yMn96rRfHzKLomNWFylKejwH0naLS6izgaQiheTiqIhjmli+v4SVwdn2IDZD
a9cVKY7bI8v2CcUin1GsVuzrV8uW4NxtJbZ5+vGL9epCrXrHE5ewmAI27/9p
vtXZVFqiX8B1n9IU7p+EPm6DFBmroOqNlkevdj6L92gjZl0dq9jnyvlKxqVV
3bNU2W1rttfAG5EkOgFRBf2HfpfEwrVG22Qz6/Dfj97cR0ZqChoGP4g2vXn+
GWbSDkph7yZ2LLbIlJSaAIS82CAcTs+bQb1kpS7UN4/sRaJk0ZKWlXgBcvr/
WgrfLQuqRdttxAHa3ub3Hn6iX6yusOQcHxb2M6NYckmeCvzxBOPwEsC4zlFm
ZQfa5N4E7DYlZqLlUs2LZLOpalMftY2MUPl+eTspO4TGvKAUncijCX6QMziq
jdw2bEnfk1OT/6zj7L1frAi0RMGWgxpRMTaffLxEEC9YAKsCG/MXZmNzDZ3R
1vteA7dEZrmITFe+iyGyHtd7RUvp1ia0XgEVSi4Wl9HQMyW8ZawsaQ0JGum1
xsFUdXHyB5a6RnpV5Z/VIrmbrHa3EPrglmcqTSEaT3ITe0cReLIjG/0cYhxS
yaKcMgv6KhJBssKvVk+IhDacNuZ2NxITb3/E20lmM5zGaYxXN2jLNmvVMesc
nIvZB2G9VpmqHspod9RHAvFZBwZkgxchypWpwaCBsngcKVk7ivglr+dsbPn0
BUrlg5IwEpl+U0efHT/vOJsypZrI9sXSw5thAwUX6dRakmi1AF2cV4qbIBSg
ekTEglRExx1biOd+qKR0bPSrPO5H+Lm0Uctxu/9qyUyBaBeTE8ojZzTPVAxN
PcGPNBbqyYAv01yq7Dq2BwlP3IEWts6nJKF4YHRHA+jsnOEHNi3O6rk07XH4
HSx2895Qj3cEWzpWJcrG/TcqXEpcLm/xwX8j19Oe6OT39MdibCbbDOsjPhi5
caXFJ+rot2ERwy1l99y2opFSm+fdmzQHUGlys6PnXjKyUkXqYrhA5dbXaXGk
jhaZ7THDYWKxQ2DZ/oIjGk3iD6FbwUVa2ZMVpeLAGfU7gWYo8/Pfsx4dR2ss
KV1bxkaHIZrsrkOStr/PSmz4QUjV/Kki3X8s1SK0NVVS4R27KlNOu+DOPbZl
itgLOEy0D0K028KvMsBYO++DSxELQA+E7Nc5G3+4FcryFfa0hbNhdlOXB8gC
c1iRKQnID2Tf4Dhd3MYjFQHKr/zZfea0MGDpo6zU11z3/+No6xy5J6gL5vAa
PNUFZvdAJCTVBqsdS9zhYnkPw8dmn5YUTdetkRc2Kd2RHJkChAnQw58CUDBY
6yAALQ4dI5A8POre2DsGUmKgdfSNlFRfv9LsQumzBRo7uMM8W0RHHpiV0xgy
bLH2R2l5StY9aMWCsQN3Asv/50nceguqiqpTA2y679mohM5Yh0PvH0XVD0tA
scAT+PDHNgzq5Q5dwj0Qrjk98n/MVuW8E5yiBDFdREZVAI4NFjI/HX+uld2H
ZChBtcAs7j7421VjpWju3j8ODao/rpa/1VcHellEbDqZ8sILtwevUF/nHqE6
qYqiuVxAZ7K5Xs/5S6YP19/MpTHOd26e2tFXZWRpzHHr56Zgt9StWqSipfG0
3W2pCvAiAHQT/XrhDRUr6sdw4QqE8k6eyOYXU+VlK15MfCgFnFWsi8J3m6m1
/sjQEsUt6nBhS6M4tKvHLGNB4OQ0n99nSbwn+C7CN438dVPyibzGrPd6+iiz
elwl/mOb5vNEKN+WiCfAaaAixaNWj7CJ7lDQkatJjHimJHkNCkd5B5B1ZZZ4
l/3ydHa89kfr86hg1yPNrm28sksKJHhVoSWTT86gvdm+Q/RsWbjOTjhfLVo/
Hr+AXhGstW2+LcjYHs9ejHct7uP+5tRxwZAB2zdplsBtay/ClBNBUqNyE9Sk
zhf1pBLOEthKD3B9gq7q0HmrnTw/4JaHeIu8UIhaw0iWTORFYufE3hLTg7ps
o3YG/okCEu+h7V3LwdikZ4SUiTKKHtSKV577C+4CpVte9gzIi5TZCPtTicPG
maHgigoOJl0tJPCALh1qzemvg536sQo7edr2+Bv5EgD+elqPjJ9FO26KzP9P
cZjKvIcom+8dDSLn2y6FfzueVqt+Oq3VsPDXOZbaFL0uC3Ew8b6KCOgfXLNM
trWNVuVdeFpLGJ3CJIpF71BEUvdsHcNSdCkBUSfRJO6Zq+rMW5/HIpDvHo0V
QHFzQI3p+EZBS5ADxFN+WJqRJ3J8M5MAzLeh2epF/RmO6CgfYD1Cer32lfGT
vjZkTy+twABJj5vwhD1hwq5lA+5qkv6lr28KBHWo6ftUr/+0VhSiU8QWTQdz
4Iv5X/ymqGFlycpdGS5vy+jFbgoLaym3dTTnsVnz/+hcLnbRLf/i03Rfu5hI
gE8soHpCLHXHac8mfNb+pw6M6uOYuODNOAntrlAjosFGQfU8Idl8KhemFtML
wFLbDygDA8gZOo6oLLOF8EIuKkPtFpZCNBnjSIfwffnl8TzB5zrLZZYw2rNz
khERy1TKQphKMOFL48BHh4NUuSKsSgr7etyIyRoHKRq2aITRJiKxTEjDAvGf
tVYhCpAiwJtYhgr8DTaXJ4Cv9b0BWWpmNa0UdQLsNP7U7Zm2FpHrLNKvdlSw
+BcGhkQQZSxsdgRi2vkwo1ggT+S9yg2ozU1VPSrkQxMpJa7LwO5bfFV2Bn53
C8/tIBQ1dhRnvdy5BGdAbZs5I3DO3NZ19axP4enE8RWautRJtqgtXfv//xBp
ZC9mliQqjpMQSyiDs04+nyOmuHTA78r0/SfrdG6uvIZ+8pbqZ/uvChlyCcM/
3lhSua9kYz0LITVT/zN1+0NOf6B+IaKJG50o107RPELfUF1RGqx+KNELYcBE
nOikxzahAH2MlNt81h5gdBZdtk64P3s+r2MkU+45yivjuXeLpi/AnMs9rquW
aNou4XhWG2tF9tBiaxzlfwNzf0ScqE4MorL9Pxz9T6tGoh7hPo/5ZdzKOXJK
nXUaMeM1BQKvXUDEHOxkhLYaQlCSnJSyvBg/Lhrh8DWn/ehMWUQ4JhaLf+El
b6T2DtNRTVPQU4KpMWbTfQimbZQp6R0biSAZ72YRoTBJXjACZXUd2/Wsmv/1
+c3LKDHfyGwaaPK/t3UrJHG/CTfR0bX37XmDwapiPE1tb+i0rHNVlvIM8epU
7A/qJn4axHhDgJc5KJCaVTzDkBZC3s5573yJw2evY2YLMhZR2BX4eNUgGivc
kmV19EDgfxegG967Owzl6ZQDWWPvSfomHjY4F/zWwYDjASmsO97ACIv9vhw0
C6+C2hriCHXZTc1QAyivmNxYqiU5ua6Sm+VgzpFWwBOKHicoOwD+kxWs3olW
WnSHCMZEPZXZ4f/IZf1aByKml5gC9+l8jxNx0tKcguGTxCiVb1BLNDBqdDdb
6Y1YBj2VV3uNID3fmx56wtrNC5fgiRBfLoufKPOcmDAJTtq8MPUvk1q2DwTt
679Uy/b6/0N8SO9PUK0U5yGA72QivMj4o0XHwM9CozkOY254pOSJz/jgCHjG
sYrpJ5diBK4wnfvDmOdl9ms++Lj7b8z5z1j+lzff6BMuWMGF1tFoCNB3ia4Z
NZZEGWbWvqQubOnHC8AVQ93w7OTcARYuzD67NIXynO2bCBiFYknx6xThTTri
Kl314Jlnw5EhgrGqvtqwTALTPLmFpVWBtOHEAsZh03fc8YtF55tkiYEwsIuq
0w6w0MR0VH3hq09LEq8j35AHqR2f5t7CxgsLgadc7Ui9iVov03wtO08/iT8A
nGG5wnjoB1tCRlJa9arIkBSxMctYOc9PBMp0sJiqDcSzTIG5wJE0ldxEtbCl
dZbre1l+wS1dquW8BMqWNRXdFzT0NL+ubJY+q4qlWIewr55JBFZjUYkwk7fC
9aFz0ZYdOdUdizezerluh3u4v75DlnIQcK5kudA6clwMtZMAE1RDgXC+/4gC
VYMDc/mZjRFE8mCpoeBLuhifxg4rBsK7KEMSvp9D85ueFFDAnK6RAqknLyGM
J6Wi4oJlDHfSFyKUmoLk941KmHcJqAzYVmsAer8WWDyAmX9wMsxlnnvQj4o+
u9+6r8iA6mtk52zFxLV3bGvWpsfZWMYdtonPs0ncPxWP080OzLy3NX35ZzU7
GsdvxKtQHYHsJF/G34ZwLnVm5rQgymGsp34krldUjdeXUPtlshAIBqp48tJo
bYOQ0UX2lHDI/q7Wm2b0djLp701nYrH0QwVWOy2FybSKaFmc3rp+MDUADhYI
BJbPOdzdH1FlUa1QsER/qdYK+riCNUIyWes0paLboIebypuV2u6Dy5+WBgp9
f6eUMa+MsDshNgPbjugyE3qR37/AgyGr4aEhPl3YcBKYnQBNT8OD63UuqsTa
4Gk2yYsEVvE/boYRFgY4qNz1YRMQEGnQQY0VQ2dE8Dt2/RNT13oiatHoqeyR
H08visp73rsv1s1afR6cf93bZtgDZbH1jlru5TTpRv7GD1t5ZVdb9/xdR88l
PYZCwBwLFwlLcl9msFwOaSF4ht6MzQ+qnTx+M68fsnKtclViFSTF1PXtv/RP
6hr+oNzvcloiW6I8M8LJfP4NMe7uociEfx1a/ovA61F0uyUqEGCFW1sVNGYk
YXusHrA6lufsxFxRsBTDdIYZRYdUnlKPkmL138vmdvLNBtLyztH2FuR7uai2
KrlMokRb+IOGMi8aCqyiVL28WYSxRXMwpHDqYc+EUJwwYVRMlg2ucxyq7zbQ
kep1IOq89VH8ARY3tBHQniLz/AqjqFKgGfCWLihmP2kJgQQCvQ/LSkLeWDat
dguZmu+5CdC7PXzwHu1yOjM7rykDMqK8CjLFb+d8B+zfMvtUPAnqSL3E3ZrQ
Q6paiX4ooYQgZbH5uf82kJB65MYuZ2eOWna6DBrjHHkH2/gr5BdzPG1wBA51
yoDfBsYbdSycEZ3i5w+b++zv1lSGvHAS2MSIyjdnNDTZ2D3Pto30hZsiaeN+
gwqznBQjAvrm5JDPjPOTQOxKTaEtXBx24yCfxrCv5dkP4TrIPr6xAtsdyL96
RnCZ9v/y69zFtLp7up69l7jdA04Yrw1xeKc+Qj8ruCxQmXOzwCeF+dy3qDDO
5sJ2oLG3gwdXdTsToNWJH8azIwK3c4+Tn5fyOplPcSOp6rB0rtRBVhstctA2
3FHk/hlISmnekvViftbDTFgjVLiYV6R46N92tGmRk/ZXQBe0eg5mFuaB0uIg
AIc1Dh4OZB62Jlx4kNiPDI77ilmKU589G98EuAwsI/Tdi7TKi0q39Tf0ULmZ
4xGmBuiIGjU7DlLYUWW8eHuXQoN+BbXo7KA8UqlaMlGwwPmU3LOxA7s+Med3
KveWygy5o88XURCKftzxFa8W3Rb+QYrQp18aWb25iigJXBjlh+HPfr0qdaHr
JKiNtowIiWGl4IZyykv/T9SNR31kYtNrRBgjZsNdWrG+Vbuokis2WynmowsH
cbyRGGUIJO6sDf2sviUUSgkdZAyeJZOQ5cfWoVN7WV4u61UmHbaXQyNHIi06
Amtw65+hNTN4igahiqrUu2eHMNGto6Z96/rrTA99koHihN1Q30NcIDsQyiXF
l4VU4B1ClbcGlpeLOuUaWeGAV2BDKk9T0Sx6uvJTgsTt8NWHHa79PCDqDCKM
ewa2iykIjAeQPVqeJZY7HP+xt7FJHPf6GwYH4FQNbDevUJHfNpqyFeAhj+BE
qd9IopdLE+kb45PbfbJ5QKUt7WxRdvmXXHBr+ROh0E+mAa98ZN/U38LSesOe
vqnVjUQ3YXOs14oXhEAOOlac7jXBPN7Czs31XrvZjmG519huNddliH0qZfJ0
63+11GafxGBOEH8/7AcjlGrUEEfmJv3UbMN6vbWjaqt5+1moOzIiospW9qh5
HOPatzyHR7cRsceZpYh3p0I9yDxMJL7gYOJZnRNb/orv2xPbhf4Aa/f4euwG
t+T9G8SNOTF9eSyxoxHOdeJZUYPYMHuejWVUH7IL8se204FJWipBl3f/TSrt
TUnwMXH1LcPIo/OM/jDbz1FOQHTCtgLtgPvothYxQCZx2eYLBSsVUOqhpFmm
aKKTcKlKbRKqR6rOsg3IKpwW5PlBgwp65iBvtylCmderkKwphwxU+wSUg+Ea
PKTCKMHaJmAHXHLYsuG/ANBX15hYnjr+U9GR57R8tDm4bqt0GpUyg3PwDDMO
Vdkcv9roFlj2ILiiGnj4JeqRCRqGZXdxsmcH6M1mgvV2LmZvvI3W+62YQ0dz
X6fBvxQcxZkn2aNBpJEXg6JaU0FRlBL2DbEUYhFWHiCb/nlLvMqK1TAo6gKS
ROffXjIaV4CmvOXfkYaBexNEDRdnF4UFiBIAxWlk/K22UiBeXNUCLoOccjdF
bwFbY3O7OmM3YjP2FNYGQplpcvBIXIhQ5tNtcyKkZVEUbChpEOwr4ZwI0s9Y
4vJvY9b16HRlC2KJ8iUDQXZ4t/VXLDW2ASQTtK1mXnRG7k8aZ56ffLQsHPW+
SsV8F+vxbRuU7VWsIBmBxj7iMQst/7IfbJLXdTVV073x0lnWSaNQU7UQhbD8
KaqkFliKw4/kukBGGadTwOE9i53Ca3Ys04lxnit8H2RPFVY67KkBiRkVdRWz
w21km9kLYKxC1IJB160n4+S3sLUxJQVfHFUqZ53rg8vAOIamIidbixcXw5Fm
RKMsvb2vvyhNWwSfQtJNUlJwZsf3aZB7lJk52BsOrg5P8GUHJg2C1CcqUgob
BePmmxyB4hLqoOekqaaFNQX8AyT6hqSnttInq4l+IYSFSWxHhYZq+RE5ODVV
ptVf+/GSMdZ5u8xgzpON7SxdI4lz7LVptVSQTqFhdY1+caPIQGp+3/UoqzM3
AfV9YIWJco3Ml8rphdlfaC85T1n+iF2JG8qqkpwP0WzLe1lau/NjgZUu0+z1
O9nt2nH+8f5P3niC67Hbxdn1k+BIucME6HCmnz9QFfrePZ44H2ZD/6R8c/6J
43APSbxC9PLy2mwVawU7bMwdLXInL61xrI90o+heN4jn2BCZc8kpvgpuCIem
efxjQlIK8p4f1NfNmubtv3OIJBM5wEzLY/tGe7I/0pnXZsrXiW19edbqpL8y
AHl9OjVkSPPK+3jx+CCyq4QS98Bix/rlf8YlXN4IgojyomgIWEYiOxzVuZhG
TbHDdBOJAfjeoda77OtM5terIIhO7D1YE+E7Y/o0jQdCXKOJA2OMhvt+KQ1C
BlrDVmlNjWSp4rg79DZA2ccdPym8gDG9C6K459gyCVMxtfcL6DvU9YPk7q6y
xONgGZCvloqmcrrnSwhAEBlKPL/KcRVr2mqG+RRC8r6mGaiWuNvmvpIhCodm
hgymdfN3k/CmCnWHrrxAfy6v3d13pUIF36uo9rc7Cdq4y7WzHP6VBNH0LgQf
b4FC8k4h+ndgQNbzxf5pYhKEsWCydpFkus8IU0mFwvmrIj2gV9dofpYgMHyd
qhUFD4BQ17v5fjKaq5fNMX7+1zilaYcQL3hzcV/+/pTQV57Johp4PvYK2mLp
hpNXvhoXFDbUKKsrHnO3vh56npnz10CRvQl218y58K7/FyVRh5ARBgGNv7nC
pHlz1iKjk8zrMX9j6g+X/2BaoZU/JrPz0/bs/TG2lwoMDjYF7zA172iufsRe
PZL21c9U+jqhqQNUAOEKcVJEHBXIeainKEcufah2Cib+UZqJ69Fsrha5hgwR
QE7e0LPxbMzSj+XE8iwJ/G+pYeQSKolfav0wnu8ppSrR1fP+evH9h7QyE9PQ
qi1vnAM3bCeVLj5EUGReyu0WaUWukNbSWH4nK9wXSpUcT6t+Zeda1wjgjNLw
adSbiRQpC27XDkn4GZ9RoIRCGO1Jo3J8zMKwzN681PsogJMFba9hG9Lg/apf
38dNR55iw/2D5dHIPh6kitfxBQKAWSgTmmcixhkuhPhxSsupNDp+ZCQ3lOpx
UiEd2si+trk2xTcNmtdrRgvlBp6BDi3pTW6wnu2L4+yjSgBefB8eMbHXL3uf
psH65L7qYwK5VOkQOpX7oMRJas1HK3/qFkMOiq+/FaX0sAIFuiykifoTde50
q+StxjFdfnYMwR0VMjAFj0VN5CooeWEnIGMt+mivJEd+vSIqbkDzWMwxxJSI
3lpFyowH3p2SsIPIEN5o2q599Z/U3x0LNEExIeYoQcBsyF772wLkHcI/xZXu
lhJkuKxjVPDYtBUGnq2f8bH2Bjwmdo1Du3JiaNQEwvIDS7RS2yGZOZhFSHsc
54oLtEw5FnExRraixNobi6EWfuClnVzSxBtcNb7l8gEdmipCcqx4EVjlfrfD
tV1228q5pAI2y2DEaP/fcG3SqiVkmaKz/Ax1A5mRmzyDJpd5acEcoCs0aTrq
19DiaI8X9c1Cz0kPFXkQG6S87dUjy/moJqc/31+U4WlTkigtvZ1o2R5ry+0c
25f7BIxifV8S02/GKKZo5AbWhl5nQDWo3G321Oo25Z3qXR09oAJzbFvUIESs
9g/2/iWq6cj6eAjnO5Is9dZPzEESv2kk3B/n1+63Nzuo+2evGe3SLgpHgdp5
XLtXauK7tgz6nfdwBmjhf+by4lBSg0QvQc8qZmb3Lzo4O1eTHFp8/hB/WyFK
+dBNQBoQd+6d6W8GUhpA7kHzDOEOD6IImcCX/W3O3LjHeNLpoM/HmluaySiO
1OMdiwiAoRfbgQQ1ijQJ8eWFd2sIuf0j7JNTcErBU2cPpZKBwQFvK2G8fSu+
RVnPQdj6p86IPnEg6vrEDj9P5isZd7kSdkzrlduJki3Kkm0NV8+tg+k8t2eT
wCuLbpWS0HBzP3p6I1wSnAfaxI0nzoO9RkAshIbGZTXNIghkiczUI4e5kbxI
GdO+vV7kyygCRobridg37uBmqcqYacdb1dlk9+3aZVGV2Gqq66zddRDILTfk
X/QOEe4tPwM9fRK+KM+yNFg7G0Ff6dC/n2vaIYIYeyHBRceFllsjAtwEyO8a
9r6PiZa0XgTGgnr7JyGMAmGCb3jJalrtFevhoOAiY5Sm6jAMbxuG+JZWIwSF
e3MuLq5QcWx/sDepyAaTYAkwjzG8Wtn+o99CBf21aVGz+y7gWlO0mtdnKNzD
Bw3wRx1B9k0cuLOvvfvqasXmBvUVDlUnDTZQPIQyGMlPyFvC1QZ4l9vhSVfp
HztfS6X0IHeRzCgiTbmF3mxx/7RyKXzcjrj6GWxH+R2QevXUWzHTX4mFZL8O
yqlEcrVEWmO9Hmylsc6+AgqXmtAceR4nrpB5rS5FmaXOXnQuDqrop+WukH0g
6QHCqv3m+dAQB08JaMEux8eYKxccO85CvllXaiCniJ3+B0lDRYZSICXu40Ng
lXY8h3XKLgVny+spDIBfNsJplpkio4DVNpP+5j2xzbPJe9WMWJywQepCjsHj
/Nl2AMhniQo07JmSQ4H5G3ChMPyc+isuIZZQDvFRBodL9nO6wMk4hiul5HaA
ghwU2GtUnFloWDCf7scvw9tSPtaZsONbGt5lw2FkMHyZ+7pK69GzdgBAfOVq
oo/ysT946KeE0J+a/ht/ZaaiwAPbjjMAugdSzFZTd+HXxAeyPvNr11lUmOWa
6tXipxzJO3lMJsZ0khcbJ0zCMWXjjUY8APjyRZ0cdh2AHsyJMqbiytRTKT5u
eoKCGyH6+V2x5RWcn4oN493vPtuItrQDeGhIorpDPteT0S5GdIavVoWFQH8Z
jgoMlb8AuZE/mOIC0EuFe4mbvE5sMI581LbtVQMblGdxyjLISfJimJa2Vuks
w1cgCOcL7zjX/VcBohEe14rkqQ8ciKY/up8TtAaaZVb2UON/Ff5zktTf0RR+
rHmwMa67jjSYvRKNJMGFS/3JQuF4Kv05ui1+Z12GbZQRIn7jR7cmmBB3f0lG
E6AjRTJzoCRA4a6mGs4cX4phNgyvGJH1rjI8URvO1xWLxOuY08OnYMDq+w2Z
zjAzhXgXxfUegRIxBVFcQ51tDaPDaQpHri+qTfGWTKNfrOAHhehntOoJEF7c
x8l0w6FF3ion6/C6c6rohNwV2b4Euiu+eB6vWLPUkUxPphAQrPd6Y0Fq1AnC
chlBYUI8qGqtsq4U9T8aU6p5g5SwuDHYSssIztM75hOdZeiVuV49e/EgINnX
POG29nKw7UXB3bCtMRRvn5LqBiwNvKhuGCIXWy7eMWJywrSv+phPaakBFnVK
Ys4IWUvhfcKGa+iHbwgsTKyDhYwrIuB/rKtaQate7iGGkZF7S/D156LK2dYA
rdtcf/zs8tbWLgi61/beDpTBxdMnCp3/zMQDcuiydvOqDmnkhFkOvDZJKcts
8FiWYgZ4IYmlz/Ocfe4fwv8y7yVmidjHMAViN53doaaOgReuxDVdMittj2bp
ddrbywsTNkRRp0qE0qdTmOMytfyJw+JKAxxACN6pgj9ki8jrtLTqZyNwdCsf
W59mS68TBY6/0/JykpX3s25sEYBDHSok5R2SLPwfPpm8HpDtsYlr8SNoFW5c
i0Xe+vhVfmH1uX+A73VAtt80DrGNb4QtaXRQ1JueLifGIUb+MYj7TzNXIOr/
Jbs41LrBG8TkgKA7FCpSLr7/TzCmg1ViGgb3X1RFgOFWffFE9oBczs8uGXTE
y9jCicje66UoIZWCaSs6oECjxvVoZBQpzt43vCXPQjekdbM7ozbOrN4FQWTs
mYtcjswjnhPdgHpxPfJjiy/CJhE/7uf0OwGnviti/X5nCk+GhMVlXae3nxcp
/PHu8sDjDX8E8IyqVtX/COIkvVrTa5qrWUvISB0a6D8q3sCMb30sM8ToWzCH
IEzVkt28/jNuJkogrnJZGx1fQNgyE7pspppvpYQsoG4uouRopT7WiAUebj/p
tVBx1SCsV5z6rJDBW7RjLq8+p/xQ4KJLy8lcc07vfbkF5t8Y3t1n0pVJkkPc
l4P4HlcmCD+xvfAp889HJq0LXC9pkxEiQGdcNg//MuE+eOgbDv7ciiMU/C2d
CHS4uFVXdYd9Zqbu3eiatdpCvGkyjZStbLXMFhmpiq4uv7tu89YVNh1ZXOyo
fGO846QQ19jisir0dadIrSK81qWO8LXlk6JrViZMi8mIxDUxN59VJUmbNiTe
gbgi3/iRf8vV8CAXltInGsAI3jYCLCtFyud+GAv3nnJKDOoytIK5s3TcrP3w
Q8jvjj9RHlTQtKcK26eug4Dopi7lkUO37jz6OFGUckBRdJ05Y+IE3TgJgjTr
L8LMmQbN7l9bqf9PgcVM/70hL9jjK7+ujWfjveHJ8lbdIQqr+ULwwSUF0Wm0
R+HaqXNWiIn3LSgnGs/C8s1ydLAygA6Ozq6ZjFQeoSi66IZr2YVVsdOGtb5t
Nuq44SCM7ptUZUMGNoL6LwXta6MdCGtvnjDyTOiQCDe/MVGk237NueT2ALUl
1yVGPFk/QTqAz8UytZiTnmUcMRTbdU3WYSCl3B8iOFbpdcDrtQ2XTC6kq3z6
PBRIixRjoPHr/m2gfj9TnIcuaUGn3fM/BZKvjG6R3SVyZLL+hLHteeDrMS54
NpFXXac2qXobU0qF5IEvqr7TfASunTljDjRacdM0dLyHMHyK+17cvLq+2zxk
zJ0DprjdhdsSmV7HZxm+073yQyt6JUQ89OB+YaLgHmX/D2Bhev7WkiM495ow
LXg/7rsTMAhyy5jD9cTiZ7DC40OTox9DbobDHlD2/J0HG8jKPwDG6xzV0xvw
vBzwOQAVdKGSty/mhLiPmWOrhnoUW1A/JQFGVeSsDZB+nYgsWyonEXJL8OAT
N1r1r38mC5QGyUcTcQXjX7WJQwAtbPyraB8LS8sHwa4G3SHYAqChjBAAsjhP
0oWJMy4sX2cda2e4iH1n2eAttFei3ldtmcemcZc9/myjKktqEDy+8ytdGZJk
YMXEEphfBVMTjZRi9HvH6W07PvHpi+MYOMrS7YCbhMZJ/TYdoNiPhJUrfUQH
oz8LAB4EpKftuXos/xb99KyE+XeBaEZQpA9QJ82LjfoGaXS2/PkOWicOMnJf
K2xa1s5EnKAcNhNntf42/2jam0ICbiWb0+Cjo9diNuJ3m1O/3Ha0Aqa6Qxp8
tH8TuY3Psnoc+mPZyirrLlRpl29q3ARuNnT6ix3/xXPWGgt9lxG/L5LV5mfg
1pbKQHSjpTplX2+/MhkJldeCFilVAQ8nqBsG6rw3/qlaPSDf+bW5sDtmgbau
2PLlS7l4ifcqjUAqlXoCMpqbGWdCpuEUtpMOJSyEjFCK1Rg5PxcGpYhpwQIU
p3gH/ogxZEUH7XKG94zeK9yM+CVWaqghG8fgyzbBIh5l0Quu8/R30n0n7XxU
83s6/vmJEcghSd6kxvcwP6YUVKdHGCD3gUjkIqAOH/U9egzd7o6nLyeQhyXA
K5y2w2gmzvoGPD7QNuhmRtcXH/tB8JOMJxEArswKXdU99Nn/walNsvcG+YeU
T2RFOF1W2Y+U574dY8JH09C+EzWlIANSB3vMIdpBdKQOkGpNGxRFR3mBoXDF
PkI4hbJkMjjv7+1H6oXikM4/7qgU9K2Ltxymf5wV9kQUzhlojaGevLPU0q8p
7dnOgr5eltKG8RdFcCRt/+/Gtv5iNgl23mZOTzhnr2E8/Dy5jWZnV/HyFKYl
aI+PPs9dHqcizZALtB4QOSApCdU0ROUWkd7LRBEgEQb03W/pYkdt0LaTKYmC
LTwhA7grlpUTH3ovJv4uF7VhHMbJaNDOUFDR9l234WHVZ0mKrHEcJFJur3zd
VVAgTjq2Ac/B/NG+Ns1K/17xah1L2oBGESExJKWGyDHreETKlL/J7c1dILOG
krvV5cSWHk3ewK5UXIusH9rkeVTvVIjnBd0ygpRRxvCSbafd+N7h8cKuVbrD
+0/6YWMUP3xjJAedocii9U0ieOvosN91C6IV4uxmcHZBLPYxat6K6lbExMVy
HQNOnLPSZrrjGl0ixA8tUR/MG5J+XEi5ilr6h7fmR4deln8Ip4HmXK1dnbFo
CIvuoPbUSwMgYTY1QrZWlr2l36MfPJBEpGAnPL0q50aI2mGLLaysY5I52N5d
Sb62J4aBoPFkovMr2dftsoUwD3rTWkWdYvrrrK862UYuJJhGNNkTjPtFPush
TEr8jpVCGM+Kt3y/aDK0Ry4lewUKrHp9MjwOXyn5fUBM0UC6aSX/VMYXT+rD
Zpoh9QuuLR23UUj2NGhNe0Iu/1k0nRXTSAI5zQ20tfzoMDx24B50KTIkOrIt
Fd+cbfQSFkmAYq3DFTdnPp7Yznu+RRbTQ09K3OXC0874GTsFrXiAda6qlbCO
njIeMRvx/34KM/AWDAfyksk3oeOR9EllTksc8frKlzENJPP7vZSf7v2pM3sI
vPE8L2rkmpAAt6Qi4yxo47BSSTPKE5tf2MsVXPEbPR0IBDxfQVIVG3a5/qoc
6fjuVIJdDvpjcFQ5/Q4preWIRcIA6XrdMeQr+6s8IjHL98hOe8BDOfULgXmY
XgunNWaTpiBigiHjnRmacADOqn4G9lqCcYrNxloRhX4GhKJxIaNs+FPNEzlJ
zVirvyWtm7RJsyweec+7W9NlLoL9TL2zLDxG9pTv83x2SvVynVX1Sq+6xDk5
KjsZ2zHaQKfMcidkoEmF2uKwE7L5cogvreQPiSCYb+QsWlFMCN5rgiPGaB0R
iP7k9+aXFs01L/Oj4WXEvX1bFUfG11PTzeYFOSb9yYKBy9NC8hq8aOqATLT2
/1FLM+8CC5+RFZyvxGgMxJc0OAVFaZyjeOajeAfQ9svvu5kOpPpVKpFTLYgR
xbNllP6Y8GcwoT+q4rLDdrtb8yGF/bMQCfy2LeWrwkoghEEEdQL4Gk2/RkUR
q2d/QK0sb7uVEL28nviU68m+RTF5Cx59w1uMIExqaEfyXX+gMIfStxX2LP6B
6yPRe9b4FAyAyJJDvROYiXbWjekK8RGMsTr+5s3mqGgxMBSJ/b7Oss5UQzFX
awEKUJkcTuZ6Z7eUe2xF54bdLGAV60EMhibN65NWMt/urKeADQeG3iekc8Qt
hUWL1N64x3PAtD0ILzirz8VLMGiDClFQ0G+nUjVNebm8astHWEbSzttqa1m9
PnmpXrlwhyOqMK7UkQJlo35oTwBtbhPtzUgaNJuGN9BX80daF50d1JwEcQDF
5rUdb0NY3Mj8ARWtXxDs3zzSP3ehKjJ/1Uu2Oc3LSY/7eAcwDeTHRYTS8RBv
8YMGsCJ5RrgSNOb+BrNPR8K+nSF02C2aXK71ncNa3wXiS3RbomxIN9EKJrB7
RC09tNJIkBlOxWaFSsseIfH7HYFeRxk2h+a2CKUwz0UdA0V6amTDifXGJQus
0auVE0K65YJ0NGnNWPsfDOAslMzVUJW1cM8Sq/jJ9H95ihM83q6FA/EKc/8O
CfZMXaHjdZ3Bw1hSssD3ygOwfRFlN/UsgymOrWHj2L8DKUcP6Fh5HwFxFCve
dMzvoiw+7szt3jRQ6LAX7Lg7GvggUTdvq9XWFWIofHSfiMISDS+Zau/IJJdL
s1a5LI9zwN4A//962ie1W4BJ6UfvHcLQ9DTFl+EzcSC+4jmSf89mJP8E0xQC
yee5kAQnFycqBvAHEufX2PvrgBgWOzIlY0O9z9rs4lrCNP53ZkbHPRCSOqCU
uD6u/E22Pj89jwiUx0sUYLuBI4jXH4v9bJYX/EfmLs8QPo528/YuVMERbPJ7
COyaXBkBJx4L+uYYgMGRL3E9SCOMgXviyHQndrk1S3OYxx7L5h//UE45FR/A
NOUoRupvAkcCSJEFQz74sL1miD+6y3Gt+QTUM9JZVvMSQaIUf53GyPzThJ+1
y0x7KWMDoC4yFRAf8+odbM3MGnd1bHAuYYeoor9MAOt7dJEEM+W98U6mJ4YX
hgXUBPKgaKwc2i/tRnYlrfbFqbmHDp1qYBm7qB066cAdQWpeJk+/8P6jKx6U
YDD+dapzNB1/AsEo1hKGwWyQEM8O2cULl2d4/7fYHOQ+FBXPOqojiWY6lLX/
1Wwo54jBb++AuN5ZSNWZaaYK/EjauhdG/S8oyjGuwomjc0mSMXXcKLdJYkfB
eCzvm0z5vt3ZHWdM5QvCzoT8mnl8Is/Wdj65DNi3YvbmGP5MEXDQ+J6jUTeT
MtoBp7FRYsIYoFGnqZkMOZtTFHEzPUu7TtFUc60QEeY+Cst3unELEWF1F7jH
MBbSf5Vmi8uXBP5n62D0SkGFJopAhobS8PpHKloXW4AohkFsUgkIk9KZwEk5
kn8hSM48ytPNT9NGvYcZESb7XYGpTM4+NHUhZDUGu1HCxVwyME1E/8thr1xZ
0uJ15+o6tqdojH3I47vWNi3Jl1ORTOYKUgb2n83eUrnlyJ8I2vZxLsubzLyy
JbfGcO7a+HhNJ87PlHg/16Jqq3CHXvcZmGb5YiuBmSg0CdRm/iGGHJ7TOQMT
WiY7rLhfAWwG3vTMmUk4sHCY+7/z+uEshgi2Lyvry+pSTLWUYrG8rYB2LIT2
EiuQVW1PGlgEC5GqNSEynYgJCWuwnbric8ayfbGatuaTOM+a+R+4z9hVQVTV
qz4w9Iqh0FOxGXf5VUi1CC0EHYuco2/jEE2y6AGiVK5Kt9m1DRCqpDh5pVb1
Kc/DwkuMbwikWpqwpForpLsVkxcJCFhd1YTU3gYoFuSh8MxnuKKZ02SfDdVa
YgPEidM9UbndT7vWerxEjN85q4JDBxmy1XF1cOjZME14vd2EkcALoWH204HN
ir3iMGnHeG2xeZcNp3uTrrFgpqk9FLgq31xO8zsIWRW+L/taDeZWgcnuAFmq
GJFKkcE8w9gsWrqq/g7R/RylJ+CfzZiImnCZZniF1SJEAfbHzFV5LJepIE1e
ANvBP5AGom2kD0D3ejA8AyW4PlAZ/W+4efZ0wFhUfy/WxVQechuYLYCMaBh7
9hz6NOSdH9zzQdWd3OFE5wRLz3ctqpU7NSYMDauNioN2bXHFMTecgcjTM7ZQ
qYtwcVYoVjLQ3LkytJ1t3O7/ncP8e3EP6IG1Ze5vrH3nNB1yPj4to4cIW2ms
c4qPZ1onbHSRf1iqpsbn5P1c+M15ZXL3OX+86I2JQov2Nws6vweeJLWS5JIa
P0JJVOHdEyMrGHIrgS4K/lNxrKcp60g8ugL9kSzzHTP5IFYhnIwzrgXj7c9J
zRBIe28Z362WjEeeki2bUJxYAhV/MobkBl5BRTzPra1nPKXx/kqTMfHmMd72
M7QElEITa7MbgM7dLMkWSdrkyyrn7CEiVZFRxInmNi04DIo6GKzcUh0XXVBg
UQGJp9hTzqX8zlfuUyVLx/rywxN4eymW3u3Bh6Qcalpalb6QnudJ05j3dTM7
B8RQ0i3kz6DB8qc7a5024mOYLKPllFA2p2VbGKJkgQwVjZLvseipFs7tc2PX
BTySMSzDF52bZJhg+X0K1RdezSKXZklmgo13sPJkHGO+lWjop/Zjlt4drN03
ajtdjGrakNjbGOJbccZ40dn4SjgZ3AYBQKkYJu3mo9qmZcuTYGmeHtOyCrb0
lZ25l2LlQvCsK89+5FANcafyLxyIufAnOBdMGcro9kaGiKTyukcKNgQEtn/5
ALRY5twvo5M5YHzqu9qgZmCd4EYjZh7RgGfIsCUrePJwwRidc44Jvw1RAMvb
DLsHcuf0tJ3hRIAsPdMdavL//2yy9iBuJd3E27Vi6Oj97NVgFGyHft7SoEKu
YrvsoK5OMq2DyTRrcnOPAg+vWH5nUighN3IyhBafQKpQP8CiV7qqaT/FP6YY
/LS3cS/eUxlDT/dmfPj0PhvzPY1AKQtxWJlWRfo99SKi1DbjVHvFHDjwZSIu
qnIvjRGJbnjcjkvNQcASr9DTRdU/mtVoDnykNsGfZMVaHfEVuCmY1XkZjuc0
nNq7+4yuF6uSFf3XAVYVzN2nOhe0i9eq5z50i+aHmtWI11SdmvACDiTYgdNz
tUlDP44znxHVerCRgrNejv0hKAHMgG1LIHQaSafmAXxBDWhQILpOZZ/7Rw1Y
xkgEi61A+uAJDy4WHFikZF2GfEjo9kfL/Q00qGK/al4UYZOdxZCl2Dp7nOcL
9YjjTPbVoEhmnYDrJ2HBp7JeD/iTlq3Jshkt7DVglQw0Qt7Z6oWpWZxfO6x+
4szueaITU4YmxKtm99AI0rGpk6JPvqgm4GgIDNAeqTMjovDl0NA07OiVq0gz
tDzhh1K3FJh7N2uKvoy8ZyToemMTEgm4af/N4wjJPOwRRLbDTsPZqhS0kRXq
85gopCNMOHKIXcWuWXFDtNHPmBPN/wNeRvGVaA0YetlBw77RBm6bqmn4bPDO
P+YuhC/1r2g6vkCTPudxTEKBu8JB623odPpl4nS9hBp5943GK+7JU3Ip2076
GSEPMqNtrtpHL8ihU6rnNsefEvRBV3xV+bqJcOBaQo+eLOp0v8EG6TTxZuSw
qcf9ctiBGjmIadSYiEUUoU1rRkfBsOHOwk6s46jnO5CxBZUAIIMd9lzOrWsi
0tYYU/6tcyy2DI+bmYrJi5f0B41w1m4I/6ioS2rdlNUFNv9wDYmFW1C2vqzL
jEbtRHqIqJcOmbQzMMQoQpXOQIEW3TWiD5X2UsIjGnacjWX5f5NJGC9A0oEw
BEAsUselR8myR1O40YHDbitGbSQJoQjW6rPvjOgLx6jojCiUWVk+vn6kSBMx
iblPDFNgL4Ev/YksMg9OB19lYsFiEJutjWzJRaUO1bLRm+Vv5rg//6a6Ld3d
7/dbBzJTDwoTSpeuTdymdQCUCoBAlVKPpcGkj0XTOB5ZUVsrfWPriG4kJX2A
3P4Sq1KSXTCj0VQMVTe/VZ629zRde3wg28NBaHdvcuV2Hzb4TPUv66RObMOJ
vZAygXZ97f1Zq67pIHVMKLk7Ac+Qd7xxEFjRP9GHWaPE4Zcfpove+gzJotk4
mGXVKmjKsauyILeI1EeSGD8PprYDRo+LqF9lYDHzGnUk6DlpI3IQ6cfxWA5x
KcA2Ud2vU4DMPJno4RL9lD/aeAba5G1j0kwP0BH2/plStrFgdU8iv/oc8jZx
BdCC6iuGaV3c3Ad0lU9/9uUZAEsK4uqGwcHA92aAKDdZWxEBTqfnVUgGmwen
PdydftceM1S+mrswhB695+89ZASS+yCYaaM1UIHAuniHBkspKiBsTRs3/9zz
o0Yw9kkquyPtTgTo17LN6FZP/v5qyH6d+uyIzcZ1GqcB+7rki8sgc4paTqNO
5Vm8MSPWwzpW1fWnD//sNC2ixlrVwapdIYiEww4B+YVwCHG+kdI5PiJHXt5G
K8/MyoJkzhbUCt8E6V9bDYMyDLOPAIbZ6GELHrwU64GRl6SyRuec/IPP+B8Q
eNmFD3CWVoUFSHm5I6GykWliBUKgM+dmTKAHEtxQkPZXZZjAnO1llTq8xpJ+
xrN+lloqt4Qya2V+PKsilTNqZ1L1UvhRMyxVs7d+51wHwuUOXhm90lyrwEb3
1VX1llBfGNWubLD3VOoexDVPitzb0sQ7FH/5SWTilZJascW52rzmiMN/NZIH
7DejWeUnQFOTJrYBE3Ih8LlU/oNN+zCEVtH65kuM5aGYue8AfQEsPA2B6lTt
DvoBEV8eqZqbibe0yd1Kjj8UlqT9u9F5FHrFoUjGeVjBoPZ8OEdFrsa0v/5z
qYUapNrYzHOPo9aaNczK/rbr4Rfws5H9AD/7whx/IGMwpKoLUJqY9O26Q3AE
d5XDv8zwQkt/hOsRD1vmE5A/gypOWg9pXHVRb2C+3UUAnKGFUUTg+JaeS9bP
nvJyAuqiaHe6sxdythd53p8Nh065VbtpbH2y6u+4zo8cTJjhMR3D2QJr+r2i
3/oHLnkqMR1bM+2qxbaCNJgwP+M9MHAe6uIE1f+Kve2wPhwwIi3t10DnYNrf
m8VtDZJ946nyCd5BO5Z92hf1K7FeaIyOmO+ENY2pOH7WzAAwm5Vi5QJco/0X
UWm/McmLzeB4agkrdwGCkC8JgGqXUE5G5N8twR/xXnxzyUqWeZLksxpy5zjl
jabVgYLnmocib2RepiDV4dhDosJ8nMDkswKatPnaKVpBcZvmRPQkPaUqfeWy
auk6sGLWbsAMVBwmcb3Z1UQM7VZUY7jF1FFnWkqw/J4DkaaKWf5GeNJ4Uxo5
PVJwV9pLFPpu/YmUM3VWMsIaS1io7Fxvom8yC0yr2/sJvm9PI8zQbx/1yPBM
2P/YITeHc3PoIaPH7vXGI6a1v/cX9YZUgmYlOgQYmyyXPpsedeueEeBTvGr1
sQWU5jUYAeU95rfhFfsMoUqFlGQtZlCDm+bZjRzKUKT3qT9XLtNnkTQTMyo2
8Z3lmBTGJ7PlbLlLeFoJj7ExVDR0hr+K5Ml8iKMbtcGGht1iQQEReJo5i8AE
8AmYN2R0csR8SbzdeKtS3uVEgRA2J2Cz3QaKKMh+HsqdVFANi5xlWQ+IJpWo
EWzCPbSP1d9tfJMJ3sCTZMkKGZ+L7jCdLqC7Vy+TjxkzDSeHmQYy+xM9T4lA
Htl9jteNyCyWhUVTo4oX0IR7cAP6c/atzGPAUn+6QIyIiIWeo8fjYlQVxiI6
sMyMc86TfFQ5BRl3uwobqu9b3SavoeQHgh5/fy/KkDFnpFl4IDLot523dFqI
wDGkyKRGrW+JwQChsDjukaRnFuWf/6mo07xzGjDoemwAuR7YuRmDFWWxwv9y
rer86/FUhaxPHGwmjIr0bf4So3rydQ2vxjH7VIkjuj2dFgqrKxgcoZhl2b6q
FFeCnvNYHtzsvElnpIEmkdbv5LRyx/+ci5X2Nqcs0hz/nEySsob6Ab9Hfwjy
Dk1D2pPjRUJq5GBmgZGj+rNxMVkAzXi3tpqsLrRhO4K0WygMlou0s/9L8XG+
meRPmp71t58yFLqjnqCAFTUnp909l/FKRTmEGyqCnBnAYEaF5QnEmN/y4msw
uWerGXrUoleti//9oeRqNnPxEY2cNbNAF2l62ElULe998dXICYAX4BUay/1T
r8fM6DFwAn6umvC6qQpYOWUfmK+bpgj7IgdAPE4JB70yhgcHiRzKDd46+Cx6
kmIBrFcW3uCXH4No+9g+ekKHR977C3n+kN6gKxkUa3g9XDiDGA7fdPXksKiB
7f21Du7UJiAwNCtJvvuxekMYGpDDB0DOJ0HJ9eBaQkiC3NTukAiLZmIcUJo9
FqiFSVcIgEM7KaUbSn4RXxfYUD1qk11e553Kb3NVzOsrDmFp9f8oicfu3cyh
unpArjW7lCyJdjBl5aXX4+nhKAeNMsb2gKeiggNv1/2gFvsZGRF2dq7hHrFb
y1XZ7CBZXV9hxbtLcWj0j5qIqeduA8z8OoOVBylKXl1AVI+BzITPkzWoxW7+
vnVnaVn+IssAGfdeXwr0YZJqS8XCN59iBh+OgGXWPzeDGho/nb4a7ObRJpAg
VqQPy+vRj9k1EVdzLVwTexaZft3UIoPlpC+5Fl5+Nf3QMgZYyqQxrDKD+SO5
qp/jj1P2ERLKDlv+uAT+NRLG933xvHmagY9+CRK4K2NO5b2iSC5NUQShlyxG
qn6rdy2/BoAZELKlUN+dLgQfgPelC3LPIMoJFyTAp3VibPM/ayMiEb+fsWVg
DksMi+wTk9lsWkdIq5mvj4zkF4ueZMNwEMRc5S12FTaVSSrH4Xv4ZzHp/WO0
K8YbcQbUCqzrSzZPoQ+mDwFSYh3IJ2TaALh2g7jYXhUi8eyusx2ksCbxXKu8
Sh97sghNEq4lH7wi0kshkIGKLlQCfttkZaSgXV0NpRO+pwOQtPtJdK3UaLoz
15cjDzUMUhGCvlZEF2R0edrunekZQd8LozBtfAXFA+N4GkoN6SfVQcYhqSK/
+xRwhEvgDFR39dPtJt0QfKlOaICKlSE7cVZ1QewIPHQd5ZbzlU33Wbq7XSmf
cevoJGNGgNc5hLUuemS8u1hLJ4FdQQ6tHNzU9iRoftKXfUfurGH0OOQns7Vr
EWaJvzJpuPwfFdbdA7pFTrJtF3pTRHnYzqhzudSvAgm6B+cDT/4JBj+wMpHB
Cwi/wB93Pgg7wn+J86FStIkTMwqjW6F3jtyulqocvucUj9/O7T4WICFHxUGc
d1BesVs8Di0giL9Yb/148gz+CEvgTyShV8Klr7k8OQAe70TUlLfHCffQEWL0
EaFl8k4S8okK/ysYdyDHPl3cd6sNKAfuXgaB3QX3hyk+RXh3OlpIAFFbuQED
6kONXnziSYvx2tkPW/Gk20yiDEHd5y42VZh5EWdnM33r37WVRaGKO9FTieG5
vdiSoG1RNwScSvEbRUU79jM3IGELr/yCmrTRGmO3rf29swGOWyFxnvuU2M+t
nH+FgBbdtK8gI1/gJ70UnQbXwmB69IJ36L302BlOxYPaHLSuLP1KBBkTiQY7
XnwC3pij3Reizj2zKe3A7kQqCsfwZRdn2JTDqlLvcp8ib7ZWZtjx4FQvcMVY
FSIxqULSwAE2c9OMPfLQ50vITYYw/1UmYOdpDbmq+dEzq2KRPXJQIM/q0r/+
LEEdgoV88D6mFxIeVm7fI1bS18UYZKk3We1RmJdQzi0/ySU75kuax7CqZ8A/
4mjHMTsW5kP2Vu5cQkEBSskz/zIQdbyDm6Ot81pMOIiTcX2JB7reKnV1l/N1
gQJbodIW1pVSmLZ2VDtVn7yjrXSOBB5JxGDU+li8o0jnVyjg6dnakosnBZgn
f863sQEo9cDfYW8M+rDpt3+pjpfujZ//yY3/Q7ut13jWoxvNEcepXw1oy7VD
lVmwE1K4QUzpj7T0kTGdfL0HFxSLI1XonVThU7jgAbfHup8Wo89cnrkxowVM
RGwjjdUI4+fXzNYtRcKvB5qWWPMd68rEyoeiWrErjDNTsTibFX5Uqk+i3Tg8
hD7ws1vrY/5m1TJ+dh2946h4XKdCrVFz1Olox56Q0dmr4MCcx5HjALZ3EGTV
S4/fdJHb2egUL1gi+CBrcrnfgHNCAEm6j7tIQX9ChPdEtjF+DzXDqZPaviGH
/rltZxN004hubPldqW6HNgyAAZfE+HH2UIoZeeQVezZBcAOawugfwxL8zHFn
j2MIk4G379i6C/vt4GXiiiVBrDCG8ob5jaZnAMB4z7aPbrsusvpnF/RE5ZhN
E6LAtHLUpdvIGj4ZMHs1Veo2JWC7S+I3o56L8FTxEMokQettVECGxj+Gr7U9
zPhHu3u7kN7xDOj6ivJ7xZ6iVZpwQA3+E+RUTDtuHZzVm3gs1Yq5iivQm+dz
MVLfL5ACqACc1oXdA4JPWFikURLKebWKaEeMLKY34wH5wj83bl1gVaipvAqY
1QO2w0/CB6Z4u65yfVHteYSMIJOTX6/BnmEUQj+Dg18Pscf8Lr8Zl8uBJgEZ
z6BkPRlHa7uNWAVqpglycGOo/0pJqweoC4f3aJufmATpO2MBJd+QzCkOZrN+
VVR+dRnqtDw2GKHRLjetBOFr1f3uliQnM4MfBI0prW2U9rUH7Z2cgYwslKlW
0D87XFi1NKwYgaWctJfeSnckeT8DVVtGMQLeNrVy4xOtsjeaK7stqYCGreQ1
XEWj/ShaIa8LLjs+PCZ+o7MjxM7SAudN7yri5w756s277IDogN3Mn/PLKpaf
FVk7/28XM/nLrMDmyD55VaoZsxkjt146PwNcnP6PT1PdgDgBIj13GOzeL9kR
HZUM/A3IESGbTGDw90TN++g10BZNRh5DoMuqdd+wHD5aVi1DdyNgU6Nue5B0
sJtEVsLg8HJgoWc+cqi22H+PmEO7SdAP9o0pwhcyl+1rBc/AzH3I8uP27FMi
yAp+hvyW/SmER6EkYlt55CY+PLOBbxf/psUQIgJh9qMHpirDJNtRIwLu8hL/
+gzbQMIzA2vw7F8M1ZXpBBU2hzTsEc6I6zDE98axclkMaGPSGQTDBiqIzn4a
IvXh96JwBtmDBBLdUmoNeGtbX9N1MTB+MCzWMEt3fW6q05traGV/SXST//Q4
HaZIvGQ23jJTAS/6BGv4Qeth2HihtnHiwlaHVjGkVo21Xg5fVIc8nX/pj6V0
SXATBZ+SX7C24oWaFYmBQKqfNiIx8eVtbuPA/rktTdHpAFkqqjrlvmbxg7YF
jtuIhvoKLWOfQtnIObI+Qy9xG6WbJ694pq/oKgxgAbO7OmFHqVfEKFfsEX6O
LuYiGJr+VVNQ6QF9wY3kDXrFU7J/rHKM33IUAUUDxtMkTdKV5TISyim+va9z
rdXQYzrQixrM9M4kPD5BauF5haRPv93eV9VpSOs0cPpzEKDY1uN+ylmyWO9N
+OabpR636zLrhrVfWT7Tof2y3vwIWwArMB2Tp12EY8XyRnD9Nry/AQkIVThs
wtDvVLNhWXfu2oWzxC//pD5tMK5NA97dRJnW0don5okbG4Cvh4udzho+KUBz
A4poe69v2cdgAmPQmRQKqj3UT0dXa/beaySPsaMSKt9bAhiiPrvjZMn+acd8
zWm7dgviZ/Srgho43ytUtwKygHKWxCxmn4el+A6CP434ASZzCKQ8xBeT9U3J
0cXHejr13S/uUOFL3FmDDYPkkAsHk02nzZKk+y4Wy1qqIeUrf4uxidV1ohQL
o2q/5Fv0uLP/5muRWq1BvgBC3Jmz1KFdQTKd52HJRpP7peHBvWOUCdmPTbZS
zmOThVxOC+xWJ4TN/Qliyl2LvT5Fdk8zknBFWxf+WGwFEh3rCxwRG+EQT7+/
7X3nIiHxKL1VgZsAr8jsvcaYYFIT4wSMPBpywjp/MVkBqh5ut7QOuEgZQeXJ
8ZY8ko9subVprJFGQVfnbK3eL/wmIUhk5exu+3iQV8N/+e3dSlkYG+fkmk4Y
NgaBzs1557zSVwa6hH8oSQxCaAoTT6+jrQN5g7dIMjUWxaFJ6prak4xL5drd
7IC3rUn2NuOmv5B+5c8qmVCSa8I+/zmtErrwoUT1GlTwOfVEmaDnnR5B2tnQ
h1eSug+SNrN9y9cSeut2Db3ohNpOuTWTqTXw4mu3VoewMH8VY0HnyXONiMcW
5xgD6EOmF56sc7wxRBqPXLXUNp9G5U4PlSq7GIch3SzsHKjG2Zr9YfKkwWqJ
uGD4bF0lB94cB78x68pfd7QtEskOO1hdz8IEwwrFVR4kMkzkQ65etPFU9Fga
valjFrfZCu3GSOKAv//W1cyJU3/H62O/SVb4nw/OWz0xlHoTq5YmSFnjjlNl
Y1KC/8GbtIL9f+ls7wg90onZQCgPX3jUHv4yQg/FMqxK8Wvaxx8YVQs7kc4B
y7uh3TiBLLs6KziYOyzZYaT9D58j/NWcq3aVxoO0djdsZ67rA+tl9M5mWNZw
BA5j1iwHVHc1rS/CbWMNFFfCqlcmq35zVOF2CO6TZ/IgAiX9xbCMRdCg00O4
9CfhW2XYVeS9/GAHpmw2WQtTjc8JLpO3dMJPdgv702+ogx+HKSu/qEvAkEA8
OtVfnlGlYuOTiAWS3M229lfMTXph5d8Ssry3pQ9MFCAhxAo7m+WZ2HPVwJbg
EuRPu9Nhh/VutX7CNR37LR7ED2+DbLlR25thc6VrhLZy+8v+Y5aEdN6rHndV
4QtLs9qhLzVYnlyOHJw4ohHGZbFfcQQ0qWo8oPRy7nCqdSmu5/mHO+rjBhFy
4d2mmFNE7NvQ/6dDeKo3rZwbvha/wEEIyk4qHFmBdCsKuawyAKQyGvB667h7
C8EUsrYkOJDR0AFmS5mQ5TytdtgYbKGMcriiW4eJQoplns047uj2LWoIByio
AGDLCGZlRfceaiUmSn4+fhiPLpyqtwWjnP9SYtwg9elkDwKHJYvC4N8myVUl
6iDOt+G1n9faa9wcEFbz6IScQPU47uFtXuh/kKOVbdkh03y9aRUZuV5CA/OX
eBlmdXlZotUWbi27leygCHbvFqpD97wN5y6+J3hY5B8gf0sz+gqKwLbj9GTE
sg9lbKy4aNSv4BGUNxHetyDYbvdP1Cf9QR12zr41nWvLegC1gNO0sV6oO40i
r0KxXu69k90wF2PvHWFsBUZQzf2ACELIbXkwERZfLPV3VN/bqI8ubkU2m8OL
z/qA+YUncLjbCSUUHGHqoaDEXSTTtCXHnpediIFYpshGnW3TAQx/SxjSoLk8
1jXsqQWMkq7hDF2C3d82juCZemT/xGBWpGqWe7QPhsbePQ4HwEOLB2gD+3fJ
Dxp++B5lp7JPACOtzu1lzFQcskfZkOORNequFg1kvl7vsbpcvhqt69Iznqdr
2eqU1fGSNvaszxHwFtr9minFr1IQtWCQuCT5aFZx9hPvzOL7XMFrAwKWQxKn
A0BHApYCxVgEigkSjgR5MXFTURORFvZvEka+8CMKfZzS4VV0s/liQ716+B0u
7Gd+EA8qb7vH5ff8F3RPw3J9xvGnenT0jUZjoFEwTrO89Dt47H70f4up+RUu
ig06XfLdXAbNe6+qMYX0jedrqpdELPCxG15fSjfKif46uZ38Lco7+9tKqyHp
kMiRSevyEjXxwX46MGYfzUdhwuRQmnWFhBXfmGcLY8m6IIkvbRgOww8Lclyf
sMwQp+DP2YzfnGqv5GkWoRqcdVE7wrsXfQI3uciaSYMRcEtPr08V2Vlwa7w0
PS3byFF672qKGNZhOEYpmjtawZRzOcetmJNozoRBmmWxuS1hbkl7JfCMh2Im
/oZ80OMJPA9lJaWMIfVwiTLvNtqPewBieVrFobRdVOIpzWvCbwksF/WHz4g4
bIbQNzgaMmJ2YXdxkRzMfxHeYC4GXUwzcb+2k9w6pbhLJrdggab0hvL96gy0
gbJzBzTXOYARqEsXYRjYrSLH4bk0AwIIWjSP1tT2mGAWRwNphNFkK79kqeUq
0Nk4z0i049yJfLeo3L5AlTLmWmbkV7EAM+ordPehzFRtI3Bw8LkFPj8n3H30
GKpWebnDiFpfHzum5Veqn+vVIyNNub1u30AJFflmtE5b0Y1so0nhalgf0FxW
ybdF9fhjDEQ4YXdjpCXtAsTghu5CAN9lxH9LHaB3B8HTb1kEhRu0ky298FsI
qAMeKAWvY3FrXpuG1fSZYEm5V2/BsRc7Zmzh56JP13WxWIJNDJS2x8PuAyxI
K7xqgTxCNjtiT9wfMcFIEqJOXtNzmCmW61w9X99sckcvvxJ1zvWyfVhzqK78
xqkFOaEsI9XNHoLCUyo7Y/0WRPRYKAsZIRXfnqhKKexDP4oFr0YpqmmGHUfq
kc+43ui5Xds/ytQVftsWTTX1E8IXfkSYyxmDvLUk7xiODo6L8hSzPsbR89rY
1B09wfV7L+7GfNprUrXFlfeJ+uTNCfU1KXsqKYypufEOM+R92KmE6eGpzQNy
MczqYIvtDU1bwAGK9Fb2/fLucuewMySxN83uAKXY9n9F+fWyHvoG+m+XbVPp
HFdPsbL8Y7wdIUp9u8ckIFNXJoPTJxuNSoSxoi1sN1lzEpDJJvGXaFpiM1y/
ngtPxwsSLVlm2ISJ1GOLxPnGX6tm9nY7XIps4JibpP9LF4aZdteGTy+HH4bz
idP5980Dv9Mw/sDSeiGCGwuqaiDfyWV/Lrj59BUxBJa6JeZUerZyCWFDECQG
kEYcEQ1Igx+o7ZBNp9IRk+d/34Dw1WCIXO7m+O8PTeCrlC/xG4zBIqMVP545
EbyLyh/2Po21L0ayXrsMFUatUv6HDSbM+/haLB6eRRZJ2brsbAcQUQYal00A
CdekM732M8DZVSvxd4Bz1FGkSRY7iavfPyAP7ycHH6oS1obBZsMjkW2ZBUcf
of6dLGSoIhYbzkch6a1kVYTIxIS5gr/1RcJ7P77sMsmnAQhlFF9s9lEEyAC6
3gqzybk2AGac79q8tAc0Ij8+8/LxWB0PDEC28c6T7t3tDbzk3qaa4eEc5MX1
HRU4QVFsgvDF0rFfe9NVkJ8MOfE4ATnshN4vO3lq0dVUgFy5keYkWJ3w4kIB
CdaqnGJtmTcWhRZDL7yBL1rwJu9fiwZAOocy51JSzSGIJipCI8y8NRZ2TWSh
yPLlVznJOxvQVzdMcziQyBdoJtoc7y8QytMtC1EsaDwVHH3jnA0MrKFxwFo8
KK/IiF2kkWwixpI60SQ3D8VQQXnr31Ewi6g5Wb2TD0OtHTI+qAjCmb5Fy/xQ
6wOUTggH6J8Hxcj2lYyheM35NPdH9abP1njyb2T5+wRI5vEPxXu03/n0E18E
zwaJY/k25aZpC5WQN1s5CT3I93W6VTULRTAwIvu0AeNodMvUxF5si33qPjMx
9MZ9jXX9CA0KMPRClo3VIKsQS+4VJcs91FUnY+k5rfsINgfFqllp93k1Iir3
yTfBvJ4Db7Ym8DqXPFuzfk9SmLQToe5AKQC3MocPmQjYbCuXjBkgTN86ViEq
wP4c90Cb/TilSaWzdpcXNGdKLaB45me34d4sk9tkgcfSghqEiu4bRTGNkIUW
R0l+PdTnr8tuQv48V7Ept2slpU+FfWR+GhzRyRsOVEET0oHL3GpogUzfcRuo
HQCReE/BSdeuSvDuWXqAz5ma0PugGrb3HoIC/3PfcYgUy4DjIvvq52QDj0Tn
6zWVbH/OGE4twWNg6QfEJmzEB7PRMVB8XIYAVYAblrsLiyl4TPFEU9PMdAeR
FqUE3E7JFtNzn0aTWTPg4tkeR80YkBIfmWv3aglva3qKZwfUEijE6OYs8oPT
oh3TCJ1SCIFUZNhEp8XAoYsud2Ki4kAy2eJ3IW+bfsrRMFyerVJ4GClG441f
6AwCaN9G+fLSCu1wwv+k2gRyy9seapFLuA95WMrSRzNIkMyjMNGPH+L6ifEz
ed4Y41bXek/UI7ce2g+ud1ioEf4ls8ch1cIwKKIA80CJDwbo0P6hlwRvddq2
g/IZl/uvDrGv8k790hHp868PDVgl5GhCy3UEcO4agJlYkejurHQWJh87ecIu
uc8aPsNlGsP0JN0PgoGi/U4Q4oQDRAvUvpOpSVsLzOMU8QhHVR+fS49pcvB4
YXSlRh/E3R9kfBAeYw1Jt7M0Yxo6hICPRHcyGwQ3c41Se7oQDIAxUB5gPxW0
uA5OVxbPw9qRxjRh4nFlMAVcjQKfZ4goWC6Z/DaFaSC62X0i2j7Usnd1ER1a
9SOyTwbqsygrw+0bz9icp+k0cevHBPzoA5tqQN8ZO5xlSuyRcUFyW5tT9KXj
3UHT5wDe3CnLNHNltkJUhlF/jKERC+evQYOKcElqIid+IsW97xpxT2Ar9BxY
9Xf4E7Fxbi/R/vUTByGXrNkiWZ/M9ILnuFioOa7N9m5PTY+zz1JOaRImpwAc
FR94lgVuM/7nc6iHVIWCZMJWlOsdtxixQBQQm2BKx4T3YNecG6V8k5LIY3FH
i5o1DsgHyNUvZaxwKi6Cr6nmE19LcuVSchM7Fz601rWdCszc+p8bZ6mc4fyM
57oOFWw+mn7PtAFIJBWosvdt/+t7W+pJZeBXPHW6kTV/STxtFG11XXJrZRQm
rz31UkRRaE5w0+9yzVdtFjneL0Goc8VTS/RtepAdUBL60xeHz4YCqcj8wVDW
+ZOiqRU8NyH+XtAtzHdl8LEz9pDAYKxFcbHex9lz5nPHFqrz8koII3qXDDtR
Nhbi31c8f0zz4GbSftELPyZOKX6EH2eDKR1F2brxBkgKw4pp0vh4GvIcNr45
G5z66WXyDGyRQjsGh6uBUbO6K5lKsGQCRcBCparkR4lY86fIRhnSP3TeyMTx
PQaTtQ1i7NoIoZMZCuOvesjZRCRb4abrSKMsNhgGjtP4GlP2+rM//0+RILBE
RseuWELOrZ6OrBFacao2n3dagdKQLVQd7oZT/4FM5eb8fI4QuBD/GAOooTw0
aF13Kece+6OmKxl3jiUpUS4oJzzQTJVsKU23c+Yw3vVFIi2Z5mlux3Bouo3W
WVDVDGul1WqnwmcmtDiHsGO7wag2iMclFwOoP4YAGWGGF3SUo1Ijhq2KnpI0
UiMQUHNCpsvYRpoMk3QIEvbYik9RhBHZjy6g3Q2vAM8Eu+OnOhO7uX+WNKW3
WjsNpu656o1P9HM8qY56H8ngu0lz65bMmdvXs9LTfARSJ5IE6ym1yZ0VBm4F
Y2WcS+E0OJaDZzP91Z+dE5SOBUZAU3hh/AvNYgISljWGe4j0fT3Iu5oTTxGk
SYtCe2uI4oBHIOD5QBj64uj3iQc0/Pmwy3wR402JyY5ootkle0b4cnB1wdYv
8fM3HRk4wpbyAWG8dB3PRdRsRY9QqStFX+TtOe9ehzyxE9INWZFTpMhyfbvs
3XdMxpLw/+A9tKx9MX3IMGql9EezmJyvrE6G5VHp9L/QZs9nCh/A9BkKGXCG
K7dvfmOqXTLWxvkZUL6MPURJkv5qsv+DKO5rOhisHnCXY4gP6d9OXwY9/sKr
0ShNfyNd10hf84TotNMDwgn0bQ1ku7Df4Pf9VgEDQf5c7vDv68r/Bc6OLxpR
Xz6cHzMvhhS3LzE3wRnUZgcn+RxtV12Ykm77OKjtFIY0aI9w1sULnIqAz1gK
7SHVOlwRRHSdyFV47epjbJvZOZyx8mOsIV4mPfFOtyzBtpJIVm8cG6YXJ2CI
8RUB6VWMc/XzEKykX0JIQVU0h4C4448TT5yj9GFRWFCjeSr0fpHQyBMhwh2D
7H9Qbx3/fdaUEhS5+PizC+6iVNWlW01Wwz3V9T+q4mYxqRiXzm+EY0LEZnet
Ga5WJH50ZW+knDOxqGYqmO8kHA53RgUBL0O0TxNEHtRd4v5NQ0mYB0hEeEz4
dlwSDWCdTA3mUxkHBJCUBxrkMDo8WIhw3vySuvRwXtwh5IPuislsL5FJr2lq
iWbNTgslpdsdRU48Zp6gc/jgHOf0CCUHidE6hrDjBMYVF4UyxV8wiuFyhBON
W0lgHzmMv4bp14HFSRyDxgeW77k3ihw1A8DuaIyGBaa3BUKKmwN136A/Vev4
QSY+LynwGE65Xo9G8DKSv84je85C1CabPGMi1RLYr0PDwfwcDxn7AC9LPFEZ
ybQ1xrkhqGy1KE+OC/ZH2V1qmJeFH7HmrG6kY6gIKcvlzYsM7S94qgU1nA8G
vM7umQUj7dw1OLyjtoiUpt9C3qpY99LLJviICLUL8MbwX+lSSDOQqz4r5YvC
C/xM2Dg//hGrVrT0mkaEZ9R/Oa87Xw6yLtKMxY93sd5w7DDaLuKQ1fzxWhNz
EYv455ZlVdAULCw8i4PpIzc0EHXIij4yuW5LNjoCa8Xn1vVGpU6oFWPl/+h/
Y4fyOLOgTu4pxe87AKpVbpf+5R0BX8oFwJcwjMcw3Avmh8ln2QmZsqf/70JV
PUZwAyPLrJYw3As210ptRie+fgmo7WzLDeLxuPRKWQJLGZkLjbg6ewN0MP2m
0JaBqufd3AZRkX4UsyVSAuRstB7Rl3xx6agVQIz0GqT5jQxOFD0uVdAIym0y
8qwndAe4tEdCmS7TjFvTbA8ZYTyXmQSetHI0f2IgwWfNlRXkwR+xQXmYJ28r
uuZZ2JMyYDAm7ZdNWX2HbWzP4SLnIpeu0OCNSQBc9xcRa3JV32r2gTblk4/y
dg+CcoQ6yjzduU/fu21xUk83W2+x8Wn5fqnj6QqHZryEqkhYJC7QomnHiKSa
NBDc9aDdiPbdIisTYis2JAf4Swm8lfzyifg6rRksJohzuYLwPddv1vqvWboA
B+4RFO9HgDW1klpuHFPVewNhGhsXxhSpLMFLsto/QxlvLrCtThFi2tUrZ1/j
jON4o5QRoglwOs/IozGHiCfDgCXdbqe1O7CYPKtNISskSXa4m95Tu5Wws6nJ
4vzxJGuIu46ehci+PzzPMD07fJ3UgwRA7bOGTj16ApWT5xKba4VKxUxzrMYJ
llgppIzUyXSjXXxfAhCmj35A/jIm6aB0QyUSGnsb2DVEjJRTEolX4Gu9hRqK
35Fi4nU7lb4ZebrHPLPK2xvkGyXHlFjEqEOBtC8Gw7xOS7RhzihdgNpVnoRC
LI+VdcF42mkCCTuCyN5ozqRmgtW9R92eJBvGGbN05Lm04H3odgabDaDeTK+C
WErubS74a2GGS+x2dBjuaOQRtkmkkRjF9MuDTGtKwLuSAFtcBMyiRZ2sYT0P
jnDvLqKqoqLqACHRJhuztTWj2+7k7oOIodg8jeh5x0NRDsDQlzAVyO2+LJ07
pgbe9JXvr0X1N6QpMBDqmhxD27wVWDryM4VXQXpi+gc+VgvhT+uWejYajxMs
eEKpKSJr+euiSFAt/adKFBV1sjt6oGoRCnKb/sryXU81adXk4VjBwSQvn2DJ
M91ACGW0+jwGTWuPr8xwHHeIU0ahULtkROPBql5rkZoYNjaFYTi2D0J0+aWU
C8Dwy7lB6TQVQf3PVksk/Yd/HsyvUOV7h/YP4m6r3FAV7WWvRAnnXtwmg4KO
TLQtUSsuhHL+Qmt93umiNj5F0hugQrXOh5NyZut2NtRUuWQ7unMEnSCdJhhq
N/HwwWj6JF8HjwP+rdbGMxtX3kGoCHxgEDy7kjGm+VzrmiFHZoMz0STuoPTJ
P+jE6hbmFLx4AdSFkTuMOh5SuhV3bJKJVMmoiZ7B72Be+YwVsRIZG3YMxaxp
QVnL4bwCUBBngIvE2E9iGQbf1/LZBq+oqGbst1vHM7oHLOUBtruL11eI2MzN
AfNBdr99FXmKGSoKSAoXe4Z/aCHzbDl9EVEXmGxJ+F+i45RMJ3FyKxGSnoQF
7gRCFgIsyws4qmxS8CwCqnN/x1Z0G5uv2pIKB76CcFaR43Ywus478xwW9cRu
MqsIuO+2j0KkN2xqfwRoHvCi2hypFvzQdJisHtJeX+PjzMF1i6Q1CTBfr3wY
VDLYk4PK8ANwjGiHuoF9EHF4RNk9ZVRbDrDg0vzSgEccdgyO0p4r3I12nDti
xFoatKkRw0RMXxaUw8nMpxcQ42q1lB4JAZemMBiilizTRtlEOSRhTjz79qzq
zsLg3bGvJRtXMvB8aRQ4aEQKumax5FAavErmjv6a0oGl39ZPajjnzfN72FAu
TMosocIbVYvZXODjGha9r1KRvWhLqYjPaj2GrJNoFWwjQL34wpRx/Ng7tCxJ
WamCkRHGavocJfjdAwSnvgp5fYpK3ONG5LeUNPsWtDHLLvoMFdU0ENCPzaJn
Z3So4+2CYCTuwdYdoq7J4hpVBB8MnMrtCje/rUJYcyBcU7eMZjFTihlAVbO3
eSsG2P9oXJOnIzRfVsm5dinXxmQHWZ2+62lo38Z4mvlGY9EYL5OAH/AEwKiY
0AO5WQq3JwcumkLErl5oGYTC/OPEL1C4smK0VgecBdTunlEKJ1kc6QAYt8wD
EcrPEDBzKMffaoNdPCyrSI5jjuRbzVLlwhrvNV/PTPFF7ywt2fwVTkkSHrKS
cu3U0dgvwQBTSlHqDgZ8B/KkB0r1OqWAgfUhwlpy3VtgVpAZ1IL9tTtfPdHp
Twc+0CcAgddVCgXVZ1NU4Pt5O9XjcGv/1xSwP4gx6Rdj1ZnZx6C0L9wLpVOX
HO82TbUtSVvI4o/jSSvI2hVqhZM5YOoxOr8V5UKTb4vP2Mwlp8PfZ/8GBydF
xg6CdPgaRR76/waeCqHA2HtBUwUhCoR34d2hH67ezvRfSczGjGGBRVxVd86d
TFt+ocvFNWh8Slt7OxewBnnCHZzvn9G0ZycUlzgAOHXKgmwOLuyoRqG0dsdp
hKEU7KQFfPmpy6+9naFLopIPvCfWcq4uGHr3ePqQzlV0VlBsFYPpZA2ZPjkg
c3Aib4UwnMw6spJjRH2o04S4378nCvrB6FKUrijBJvIoQT1bLts1FlA/wM8o
/0ZzblksSWmWPJNzTzz+i5VHBtbzOyUqc/ZeuNc7xJUSIemsay6HZzgM/ggQ
V74aJTetQLMwdQO+mtrcRMKVUoATmAmhR4ijTCMvaEt1aiENVbZ3rsJNXWlD
zkUxSmmw1Ju9nqefkMBcRUwi4bWB620uGFHE31d3bS/sM7rdZJ1anyrAF/9l
k3nLA3skoe9/BThHSi66ruHRcItHDJwbLBkKQpQV9JrPhNonKe6IsBXCMOVU
JXMiV1h7tMPl4Bmz7sRj5stVjvlZ1AVDOznpy3lkX+qd24PmO1p2CHELfHat
80Yebl+zNsMRifW8IocC6fSlZorD038Bg33jpsNx79/uQUn7fva+RCye5Z/L
NOUzVWDPCFg4aXceGurMiaox6V4rB70GHx/We/uVFxSX0Aex29wF2kuICXEQ
9b7o3Wr6Q6lbJ8Rkd1f9dNVfwFZkM7JFTCoQgstCCuCfDNTiluKJqVpiqqJ7
xUJo6VshLhZ5VQ75P74H41t15I/y+E789XuNhvk3oqDRUZ+Xt7SrWpggvXua
LqG8nsQPEPYpqMZ0uy9oCfr6ha84P/4BP9jy5gm7s+y6pasdk2fHbH7DrGm2
rb/qRffgJ++MpIm8cjHu/Jiw/gbZwRBJFb6gquE+QDQp4AnRCLFjrfi0sNos
af8yD69ezNYIBObGN5ns0v774dPqXXGWRG6vm1M+oYzD3oi5Dc5ZamsNM7y8
8hiRYIySXsdxT7xupqC0icv0tU9lRv4DcQHMiP6xFBRvaC8+UxuBXhaAORCA
CJKRomEd+sF6coav+VWm80fvJKWsX0+6yIKGlDxVe9LZUnq6XGqNstY903ce
/umvBf9tBiARzybMl1CppgV5D98b6qG79knp734FT7D74o8yjsAeQe4XBhm/
QC7QiPN+H2lu9ofuFMbE2pju+rkYsMCzO/jiDwFm41DeMpv0b39hh0Wqt/m8
wQNgrBMXW2fpRnqFUDU3WKxbW+4QzHf2Idfoid+74b1ZE0yKFBNnCHjBOjbn
TbEsyuJFLs6Lo22S2SBZiWzc9Le2HTfazDgK4KPflZd/XjUnNvQqmqDeX6Wi
qqi5QVjjg4j9Tec1DLaqUx+bzZnblTbQuoL1Vnk80pn2rDxCnEofKxWiDuo/
YIIf1+iA4NwMQCMvG6+nUBVe1CwdEwgQ6qvzXfVT7WUt7gAp74vf+NUQr2Wd
9MDClcWQDCOD6Kzqf/l3IkcY8T0PmlQPG97uvA0A/TRA+zJFWkea6Nj4Gx7a
4Sr1UMIS28z9/ffq6X/7cuqlWRcSJWh3Mrs4v6Rlw+ZhKGqRbXoAuUsNeN/C
Nzpf/hL5xl5X9f6OI661ChpubV25H4fr7nD9YSCd76IWnQ6QAR9ellVAH/XF
/bs/9tQAgPcH6kzYMRP4pTVSJ7Udpl5m0IEhayaKW1eeZPOLrtcniD/Ge07+
UrIkhboFhMx8rwP+wWHx66rKpg1qcqi4vB88+Zbr2I02VQw+RmcC8FBVhzlU
W8DOFOJfx6FlMNkbOqu1WmRHA6D6ZFAiPJJjPjVMs1PBWtWLGMHFgGn5XnLe
aQ0R20I9hmugE9VxOJ8f12GJZMbXW1SbOSaHa8zE8Hk8BTWaVRytZafKnjTg
X8Rid+fEawf5ykz+bkhpSemhxHmoJmU5iVCvTBn93EvBcwEOTB76x60RhRBh
GytIhV9DY2J+SKAmzKluNlW7qy/C2bBfex4D36NWFKnIDbeGPIuI8jyDxFCn
OyNXSCHix14BvbTAYhLNy6YZJ0RWLpA9WgYjQjRQX+3kTpS3IfNh6Fw5UoLk
jVSkXsw6Q2fqIDqigGjKPGwExpCGkqmfR94CeUdLIAkijuzYl3stFuhtsz1F
iZX+N1iQUd+0Mw+8CNCTr9YkoYuXcpa2HhUnFRzfyUKSMLHqCDyYeQD1Nyf/
SPGMI/k4xQeDSr2Pb3Eb3SIvefrsx1PI+p+bims39F7zCxSMX5iaNwAKy8oQ
Zgx65t8P5OxPqkJCTNJNF+2zaRs4c2uZLyUKNZ2lBK8NBZePXmVNLhcd7wm1
mSrdrA5sLCxahrld/AMJn9neIq4Tkcq81zSbvlxI3CzaxxgYBAYEYRbnFWfQ
0fXgX70SBR77Ry8xJJuhGGg3n7DHc1yadn7ht2ClpEof7Szq/58YEd9WaFxL
uInvILlPv9RMslIMwtb3TYjJT9+H4mMzbOL5b1uX2IVBaWtWSOOc3tlVNzpG
fIBO99Wisa/e1AV9pZlKJ2t7LjeVhqly+NBzGuZTn2fCF8g4ZjlUlivCq6C7
8lXuq8Oe7dfQnFn0tv0aIlwe7yIYqW6MwgCIYjF2onzqWYJ5B+vV05Kfd8xg
+8BZbNLLnb1+3uvG/8kdD3YrBkNZ2ZIGJsJCasj68RF1V8WLTZFgGBiv5089
Z3zfMo5i7Y+qUyWxeefisz/Un2Tqwn7ViVV2V25dE8aLTj32QoJmy7xkCbPU
tlHC0XbYQF+qm4WBLxAy9eORhRZDrlbChoMP+ZsZJG0RowIt58B3vpzSFNfG
NVECkX9pgIoBZnJ8etEJmNhjxafk/145/lYySbhbsoSwcBPy7dbGH4JvoHH1
JReoFuL7ClnNPNzrrDfHo1+f5Moa7IRD0yGfVC87I6cSpypPqw1Q11kCvL0o
813RGI5MyB62QexO5xyHMlVCGsRu1EQamVgrnEv0b7VfzYOIwLnwDEQPEi+l
1oJtvsnWI759jpwx45H3C7Rrr6llyoxRqeujxFwWnKuq8tK4U8i+uIgb2r1/
l1Vb+ack7PRK5DIXgdPbjyvAXxVXurMYPH1+uXIyei4+sMF7hXsSuxMJuKvA
R8oYnH6ir0X88hKSmfSQ8XLxXvH73RABvuDlDoPRHkXpaOC8yDw7h51EjoQB
NoVqMNjNITHxlx0JjyXGMBVJXon84C6Vw/OCmstJ6JSPBtUJ1qH8NLO6kyY2
E7fSN5XJURLGVdLAT900mnocSglOIQIK1IAvxbY9Rt+FE8HuJxpYtw/6/o82
4nMK7VQq4p5z8z5OX3nbx7U3p8BCuDwUiiyIR/BAIRamKfQ1FYDt5Oi7rEyZ
i9kN/QrqexqhNnI2OPCylXgPM1Qj9WJD8AxOvMJv3lOocWsx+0JOcPmWZ/nl
h6U5dfrDCUjmSc0/jA9cqnLMy0zCyi++/gAL9l9nEB6fxpQ1sZFITcnFKJCB
VUL5trKgL5IeP1uN7Jil4Jh+F9qFCjfA32BVQTJ0N6aHHjbOOD0PJeppr+6X
erVgM69aGpFS+rTO4FLYpJ4SglzxT9HpyYRTnkqWEoKTAinwcFSVNXWXk+j4
lKqPe9+XUy8oQ5Re+2KLxiOwr42vw/lfL+jisKPUnGC2717YcyewitbGH6zo
9TZedXO64HDxY7NuG5nEj3vbgMjotC9C5RAyGDk610ngACiO2onF7SZ5VxTo
XVbx0LFSXIiKRWLA64qz6YOUXyV+ZyQAQvPxLxghkP59myS/iovxmTItdt6l
k8SCl8CBvbp+2+Ty+9NtX2TaCk+KXir8P4t9n/6Uf+MPWPuFsAoPlxM4uEOr
XMDEiTjuKUt7ToRYpn65TF+kuZi/78BDVRj11HdwTh5a7r8EBwRy3bW8+9SN
A9GtUr/Kjr09Jfl1Z+Hh2AZ0Pd9IaqL1M4piM6bsbjsNRr/acNwVD/b6S3Bc
hDfSxF1e4LkfS2FmE792SCFpN8zvOt2dxBrlkvbnoQIe8rsdkUTqBbBezA7a
vyATwcW8ZlLfu3CojrGogt+aLoypvha9sFayghEl9G6lvGFKC0Bolm5buA0o
RFSt0/tFI8bSNGIrKv8gdrNBkSxghRtFp6+Hq0PnHeh103Ea6Iirgf14U/GH
7ua9+vXtUnB7pjOnDdjov/Zwg5PC5dp2Erz0dJcT1cAoHqvX/1l54GYKZTGc
O8W8pqE7uASwAk4adJ3bmN+aE3gcWA24kJceQje+ZKf3tl4/FUaVGWpIjxRd
f4OlE3miZzyxFGf9BnEpXIQD+28HS4KDrlXuicQrpecQcizM/LZa/f8Yssry
aaBHYPaI0Q1/e5Id9XQVw1L2xg0z9PRuweFnTOI8f/de/9Tz5foph2Vb3n3J
oO0S98l0h+c7WadBeo+ADY3pai1Io7siiUq/UCM/22VVrFl4EfqJR1N24AQQ
tffA2UJ12SnWqRwq2WrokRIiVdF9AlcacBAMto7fDQq5g0OygqTcuafHftAF
p9rkZN9x0FcZQnA0C3lgtKa58J5yUHJStT0DPf8m8AhdfxdFetIf/O9lVqyf
Pz0Moo0fiHc06zXXoxBpNwAX+LlRlcAjKXn3l8B9dvmAt3eZ9QruR+Wf4xfv
PCWZNMEp8uPg7GepP7nFhTV6/QIpBeUwwavsao7bgpoj1t4pdokl2BCMoqKn
mtmtr7+lhGsgMtw+80g44fpslffGxm3R1YVLZA/eqOU9eNL7EaV6UNO4gAVY
ZtPkDSovurJ7RSXBQFEWY7Z629UAO3zP81JUnmQjY6D7kUdv8nLKjStEBp68
OXJ2aHAh7FmiCGRNCirx/20H82BoIXhsxTwKUj+Nz8PdiPK24cmXNR1+mypO
Pn4bNEasRgep9wpoonqnNllUwuUbjexfti6Dl7Lrl6iCaBomfunN97WU7FRc
1L0YtomuyyaBc8Q8WVDBR4e9e88ONUOtPGHf46czEU7tKreevkMxqAHg/6gk
UbPvP/cjMdjFbEOr9UPReHbDa1R0yHV7q0/yhT3CYY9RH/ar8y3BqG2EgoJZ
g2DLfxVMoSeY6Z2QQtAFCTws4ZeYhwdUEDtdt5BoBA+p3iVoE/EA0susXTYa
vVrQtm/Vk6r4aHLRdLs4dymAMVUDaGzhZPlaBkUiuhGVTmQPdxsyG1jtTZIe
UUbIQ+e+JsvotQDlmU05Tfeb93HXaM9x0/1LLeekbr6sLZKH955dRyqGIRgZ
zj0VK6lQsRuuyAqvK3YmdlwIRlxrr2R1fmwwgrIRANTpf/KDMEz0GREAGimO
ImIngDlnAOrVupx6iVdbdg6hL9wgYfBQSo+GJGjHwoOQLfJtbibCyoIcxsjz
EQR/gFwpRs1dNGQKSVpWiEEGmcnHW4iP5IDaS8SE6P+x/CtdxoAeg/RDFy7e
8TMfwGb6JYGY8BnkLJMTVwtM7sxqZ5MVXp4M/8TUlrqTbC5nm6OGoaYsyr62
ZioOd4wjGtX6C2E9Y6DdnxLq1G7vuMRJIJO1q2UdBT6F6GgzRkrFMIHU21Y8
7VzRjBWQXYEMwwo1u1H8ftjgTc4TOpsUxj/Vd5hwi9D7SFY9i/YKzmgfZoCy
OfemAxLEE92ghMeOuK9JG/2VQJqR56+yjxld1mcX7g1BbvjqpwYDVagohbFV
mbe4Sb5cf5VExakuH+WZCFr+5dgPsMYj5hgMy8gkQU4M5U1SX3vGXVEJRUWh
7RnWYthvr103LyEg2Y6jImzPGm7g1iOrRZBvkXmZC+m6LY4WqV6Z6toTyWLw
kr+RupWXymEnjvmYrnbIndbRGZXqb0SD3MTMCV9f6KoMArgn0c0zw9dYGtWA
xUKjUX/3n8zOTrm7lSn1+lOauwhr7AQAebrbmxxZlIuLedWOQYakyREnL2Rd
daGSRAoMbrCtsW0hLc9w7C1a6Td+HrQzwho7Z9TCgztaB2iNs3SrzuiQUboX
5FeKdCGZ0q65re12hYaFFI94ZFcLZz2wmQ8GGLnyDmTSt2iXPiA8z8CB+9Xh
0oktZpZ7GC5ci2vEb5wnekKiwmzLdPRC6V/SOHItE7CTEqvOBRUBslcq7heZ
RBUb+6bcP2IHNAqqj44tBrj0ca82hT7xS9sh6tFUTo1+rL4ovHietEiImfmQ
Na9xS+SqkSJIEwWO05Ha5PnIGN5n528H3MwevETGMZsTAaMwmfxj/6UrbB6q
cOEaWSJ3hyfCdGEpNjesgso61MYkPn0k9SgqD+ybep0wpe/odxAr/Em8CIxU
irTzBvkeuuszpO3Mx5zCnvNMJ0lYkfA/pl7OpA5pTZ2tFNLMEFjKP5hJdwnV
IZcmtPnE6HCvY377XOdtwFSdIS7z/Bto5wyWe10i3JzAON7/sbGi+B9rN/4X
YyVNSVmAdmIz6XkCgJSGWuUkD0bnBFLoXAOvv404lJo3AAbp+V2iJ/Ci03oi
OuO/k2QCqQ8ixb2HuaTU2wmVElhViveo/xXcK8ONxPC40+EkCP+kvWAnWFUv
ylgBWka/t0XdKTCrKPDOXgJ0eKqJKcW0LdJSsZ1/2sqHi16iovaH91txuLca
UZKbMEa0K23JCzRkC+l0Ss3MJ81+mQM94Vk/3SpOucKH4leku/ne9DIPWLj5
me99KooCZXzaGgBgDdySHqlh6jCo1xEOdHV1w/S2zC1/+jX3M6YDjUPoIJeq
MnBl9PJCnmWQeIyQ0DWq1rftgaWeR0ogIRm3vFDOJTOnKyvtIAUYa8NrNrFJ
Nq60qo7CBXsxiIp4qMbF6qOtjcGQvLfBo4SJqw0O+nJ8RhkqHccMnMKL2Lg3
gdjnHF9x+u9ycaGvvtxzX4KPEbmDPRUWDV2czC6Va8mIbrVNY8mZ751dP1Vs
lIv7wlPfWo1jbNJkl/9q1qNodNxCnHMiyoZNJAtYCNoT2M8iLY79Njof1Cde
i0P+0X65G4CBvnBAIO0a3j+7qVa/OfUPwoROny9u/GLDNFzNAcuvUtBsZv2y
7KmqbpoqY8308Dz9GPAeIpagiQ8sX0B/tW0WUBuJQMxJnc4hAi/BAmJi5tkW
FnD9dQ0DNtNKx1u7Roia16EQLHTLn3PRca5J80Af+pT5ExwP8gRleGJMvgWm
HCCOdhnfJkGApoycVvGUXh5/tZEd7rlT0Icro7i+4/gM2gBZZIvr5LHDL/q/
rfffrxGUIZZgYKlpdh0Yw4LQrcOuUjgux4F+lX5OlWMsPpYy7rd3NaZNYrBH
bnUnTdqqDeKBKhsNeNTY1zF86uA7KcjnnKkZCyX3TQbR/jTbpK0X5h09GXhz
qAa8umm5+jJPEwfYbiA/ikIqHDPqzZ1jwU1ZkJRT4kst33k/LeG8ouGe8PEB
uBTq3xrsrxF502Z4LZ7o/EYGwXwZ4LW6GA6wMQxtDtHGIxxcgjd4SM+R7m5k
58U8f12GT70JWzD0wQqyattRazJ5n2/PY/vkbh4d6/lyyvGVTgQhSkXfG382
qFs6SHREsI5qlHL2GecVaKCtjqborxn41XnYubA5cQIUPHVhYiCDgMoIZxe0
qvAIn8D/OZRmVExRU139yxHoDJpbjWZkCGYSnp7Y6vQG8arbgx6BUB+v0gq9
+MtxV3JHrBbcn3h0BmPTUiZvNxaWHCziJqVGmAr0icZNd5v0jCHM8ORS/3qG
MfWprZ+V29Jy8JDfub2izZrpaO+1H7a43Dfn3jGUefa6r5Vol7+tWLTL6tmC
ffr4L3QBUsi0U1O9Wdrrrsd0lwqDeiBi/wu8Ji0leqsKCAPKqv1uwgmMc170
/JaQKEG7JrBPhhDI+5JdRH8Kr5yjr6AGX5VG1/HR05pq2W5UDDLj7Vtm1Olz
w00or/8Q08P8vB1KS90zZDszHOvuKzKLiD/8ed55YkUE4uQ3ySotyn3AmHkD
1ZwQKyPegcHOe3Wd6gY/bDRUr7ne55bV0CbAlmd8YpHYfzgattolxivCADXw
QZRGSnOgcNWgESVjq/BeoG9wjbOETXK7Z2l7waInfaBjEp6Qlg+zRHZ+eoHj
l5DcS6Nu4BRBcTdkRXfYTmrjI28vxoAt08Oy0dv0f5FuYNNl3aZspa7RJqz0
10m6SN+cCZrMXdYqPaGWX4OXDIrni6M+oCk3CvKrcuVCM86Ww6LCmuYYmKtq
8HXh8vcA5i5h+bcvF9qiQ/HyDDyWnNKACUS1nvV8v4AJnnIdH9MaYHQFKQNi
hTG8cWs0mi2CfeBBXTOWTz7b7GwqnPNLVE0isWHOR8Xa0d/pKQ42thbC7nAs
gEyUyxuASxBdfOpxyjbiajXyHVoZylfUTzF6MBDvC7/G9OzmM2njy37GoB9X
RYrzCtqedDgZl1U9oilAkuJRjLsyrbdnE4OvbPDfd18UxORclMH1ZSq06oJ6
zPzxA4gZKAKYYQZyIgr+xFNBkfMC1LZ8ScPZi2zIaY6hsmeFRwTGGwJyIIzx
tTp4+Mix6ITOh7qPdsM4RwY/YvL46hc/nWvctadpOuUvToSfcY+Ci8weitCX
R+9p1xdME1RsNtzPdsNHgHxt2mdcGiRljYPDyZMSU4jPZgX9jIkBfetj+3EQ
HQH6SWPmmeVjLLDUFnuyiMcZSM0CyKfpR/jyZQRH2isvYZ5PbZtg2eczrbRw
tiHp692VgEiF4XHBdTdTBFb6YqnlbXrol9O5g3aT47ieLZTxGZkFspuECyfR
Xr6YIsox0pyzm7hYVdCCVuilSTM8N3JNOTrLMsBmFnzpa2UFktItpSlaoo9l
+J/fuImVs8KUlyiijV4D1rB1gLm2Sd1CZw77Nc9WcxxXg7mzKR1ugxi3u5ef
PYVfMNtWt6vj7CZNHyukeVm02OPcUMhqweP/pZLO9zsKHwMKfTrrqlGQTriL
cFQWA8SBgAOaY0iTComhRw84Wa4DXW4kntHIVgIWSgPJZ2muS33E7taJONqG
Ktfy8eVGA3nPUm5J9+nWU8FmxNEYIKNCudticoZiNQwEkcTkdXWUuu3/u/VD
Z+qt+mNUwLDdlSd4K/eE81QvlUusjFXqRxuska4cNtjkP6RlHo0K7VP3Xgn7
2S4rjlo4oO6sOv6DiToLawhP7FhGzvV87UijAT/3QP6Of2YJV5S64OxzdbTQ
MWRGh4g22GUQtYMtDon8Ebc0tzdv2i1iD1V0z51T2N/LqDrpFthugWgNPFOX
Ak42tWL57wsKC5sjXG0yFKrec2/1vvPXPWNFzWlfRIzu38UULyZuitd7QulX
kZ7Q/O0NXzYKflyhIcxh+6MEWiqC8gj1nZvBk2/znK0f465jzk/+8kH+Kwee
3jM/i3pR6sBhFTop6BSCaqfCcEpBwBu7KYKCYpbm+fN8HU0kJ5KJogPjcFq/
Z8VWYRr//ZIgrUh67iqE+sUvRnN3H1MkremwB5SId/xQ6wm8uFofascad0Vf
U+SvFc2oE723NaGCTiV6Rmv85ZRmEDp0Ywx8ofEn3K8oHDXzPven/tknIcF8
1o23W+OlW2V4bbnj2LnYSQFxspd5LFIzikqvJ3dCg86vkt4wk3el355bEbDz
XaURNWjsiC4ncmLq39rnTP/BNN73Q1opXaXxUdqJ3F2Qrdy3bwSskTkjmq8D
VY0/olAH/buoiPa3QPc7EL9hH19mKpoK2tyUHZkZl7a87+nJ8blQsVmRvDru
3jUVqe8SNqZbafuDmn4tMF1vakR4LvVkckadBTLsSp9i8kbNh3zqThDWKkZP
gJqq8U8+D3K8TL6Og5lkWrzJdy02BDNCOUw9mLGCgt8JG3g9xXdylkWuoP6n
HvRfOfcyfmz5WL0lm8l0N39WckTVGQSJ+O8kGUQORWNhaOrGpN3ld/+aJHbu
tcqWM5+sJCRjTr6J1Vojd81k1/XWVAZgQcVN4b9UQe5535PLyXiVsl46us3K
UisACaMR99W+kH/j8duRQ+mGo8Ws/ii4mt32mlFyuOtbtEg5FbYFKMyKz5CQ
xXZcPDc97RpXfGa1/82QWowC+HNJuK9dLfYZdMYiEoMSIVFFeTHb8oCdvOWr
V8Yo2oze8HaySh6wpsCV0Ig+8Wd2qB8XARJjNIpqGiLgMmzkFggVpAlINOcE
Oue2/6+xh8x1WaN/332z+kEHNx9ih1Jfjp+5+rF6JXhhjQjWC/2W+9jwcKcx
JuCXkFw3yNIWnK9MTc8j1iInV916P52hqCg7TnPbS336SReGUi2E/NfRI64F
S2rHas/go009XvcSW945cpKtUchJ9OvJ69sTSAfwXSk+UBk2U7xKzRu+5hMP
UwU2ZMsFRyJUnGAbkT0QEbO+Dmb4VGubSeheB+07grXLAb7VOm6qxokwm4mu
m/iLPsgySLD761UKVV8P388B0oeIlHq4o3V5fuvpvpUYQtGkiK3gFx/2ePyS
nQqb4qr6rXAwQJhFHLSBIPsIQ8WwxM1yvbipapT8m5m9CORLQFQTARc42reA
d3KOpc2htuUr6bvybmyxCzF271+LbltW8vG0feS91Mxlc7gvSawndt4+T3Lg
V6NsbNz1O9B1uC5vUEzwwFeQi51UMyD0suXJmrmf9VNxs8LplZjR7qF+Pu8f
8KUaEvtr3874RUe08qwFabsap1g/gVXoSxa6I2vSXmhhoPStgCBUX16qw43d
kg/J2G5Judlh38LLpe8P+VDx9VAUdboCYUv1M5z/U6I8iHgO5YGjpkpo0TrL
ywQpQ7qESU/cFhuL5EfsCB6YddXlmIq04VRgz1fBpCKs3j5G5xGgn/htzhzG
5yEQ+5ouN+CM50zKCGkYIUjoE+MjEHDIjhY84R3l5OseNVPchAPZ7mc1/uN3
nla7m4SvuDDhtUl2KpqPtG/alLIP0HOqLZSIoeAgaflfoE3JMOs0EQ8Z6DmQ
FgZRuMPcd5kWd9Wpx9FwgHyfYUHy1NFCpbOkgTlcwPyOGIj6wNDRrEs/Kzwe
eqhjXdqHsXsXyc9TO/a5jhc1EU+Q6MhFWWs5KZGc+vwOhu3V9qK4jguLw5VZ
SE8xjFnUA/6VsY7048z8Dr/KtnExSsC1JVaL9lFkcZZhaj4uz1SVN6E8ilsl
Cv2DPJwYbIGqXwRM5X900UZSU6ciIT7R7QPkaNyMYsV+8Jafeuo177VV1SHZ
0zx9weAjkdRBYB1rPfS9zqF7l1B9UdOqrAdjrtpJBGPrW4WQ4CGZhnnafJP0
RvVcAqf4r6Y43KG5ymj7CfyTEKP4YvwQekDXGznj6BXN0G0mU9KKiW0Ndv95
fKES2NvDp35XNDVOuV07A+wzae+PjTYGzQ7j1lRkmeSgAA4MyR3L61yWxSVA
ctPCXbvNc33Lhp7YMyIs8bsK6sX0yE8IBpnhVM75b2b9s4QMxWCcervS1uvT
eAPuZsM+uCo4kmv7OhGwT3lhAMkZorGt1SEBeAtqc4L2TCx84Adihj6xhE3a
aVPJV6Tdxr2LOpc36u9TAhQ4iayI5l/4qBhYaIbvBwyvtrfcPT2JiP9JRb8c
mRXFnz+OiMBYUTCDVAhai3hsYfX/CeFz1a+3fRFrl+eYlFZFFirb7ZJ/FmaK
puuicsXDVjPRxwGneoEZGnCQyNc1s91Jq83vJIPfQ8WpxJpjxZD1T3hMVBoc
HiPJnWpOA4T1o9ctZWgOM4orcnPkMw3DgQuHTKR+FayySJ5B+rUWBsgDIQLb
nl5ivmlsxwhI+cQ3MmoN5IwTCN/fLRHZJkxny/x4QjK4IYn9V/PoGEVVfeTb
/e8A4kBC/dw2/Luys4xTXet67u5lLSdZjFKFo2Al52rCBk1VX5qzECwHI541
wlzRTa/U40wCkcOW2uhf5UDS06TPVDlGE2MLEOllb/2XhooHaBDOS4blVKtn
RqHL03OZs+f6mgGkM1nOdRbP8rm96DObBW6U2u+GR/TOcKbpa4TsBS+qH5hL
8idKWRK5qLctfka3w98ZU6yPThi9kORNj/VuChljenxrLaNhi0s0OjkD7aYn
QiC3amdeefD9rj1B6acPuOER7ta1FtDpMHUPSUXC4qgjGRXoecDrgr2tiVPr
w+ZU7W1wBAsukgZ+LQ+V3vPYzKOgO/Wg4ulAziq4HVyTq+TIRP/dVQRr6lzk
65xycN94v9cXhro9+imqG4pV9/TtdM9nsNqqAgTWe7WQJyaSq+3SoWd136lL
PEGzYn2NhAIu5sli8CUvGK1D7D1t+8k+Z/igkDA+3SPaMPQhRr9Faq00gYIG
30mgERSuF0FxV1GHg3wULbcUo7jg5IX9UXb7fgQ/CyXDLaWR2i+6I9+FJe0c
LlDm8ScKdgJG9uTKxnEEEQ+SNWCkNRL2qYOUOmX0dm4lNvn2yOpnVFhxErkX
1kppV4d6LW5W1uXNfpLj80de6ueAxvfZKQ0WRpADR3fj+yltMCwsLMu+JPTA
eSOfHueoIpQXoaO9nV0n9lrfVDj8NCt70St8tH5ctxvY78/L/MYR9YB+bzcG
49FLzMAQd4UzLzhZq7LP3PWS39UCjL2vURxiLpCSshZGDFIYIp0MkGNR026k
+KY3r0CxBAF8KHvVs6C84VMfHfGqPJmTY8Q4Jh3smG5PItHSZ3TJBbVuee9s
gDUGyrqr+RaOjSOBO0/iP/DqBtGMXsRJEdD5Kpz/07kQ3tEH4tGEwcc1ADL8
EMLGV5ngaIdVklmYGpWbn1QlrBjAkA9v/jVGH3y4VYn34QPKhwBJf+8Ih8Ig
nLkWdT5MfADADSCnRLuMZAf0MunD2p0h5UFQrojK6SG0v+Rke/NIVNyxiPaQ
+rq6N3Ndzp0IAUj5LbpPLvSAIfZSgeJR0I5IZDjyRV9rahdFpNJ8CHTP8Q99
1BNUEl5kpICWsbLW+ITToXzVWhuQ+GmCXLETowpB/K6aSytCDvD6daZemCCX
oLsDi8+HS8TMIb8kagkCql99Zxa2NbxK1jjiZ+i+ZRImGIJlOuVuS9stPB+5
0seKqhH2i9hM96oLSbPL6NLlTpYXhQFmwM99zncJvB8S0soW8kmc8ihVcQGc
a0k4D9ZNk31uyRBJYqTTaih0dlPqy01h64LCPJyYRuXp1llyIIc1XTdutsTa
6ftFgyid6/EXH94/xy5QSUepXr6AGNmpRQnD8gW9mbEks32+JFzmgKWa5IKR
iMpr1Uq0iD78q1rDhhFj4DYgYzqxPOk6G787kQq5RQplk8nF0jFp7TDUwEkY
0qrdcRMPpMI+9MZ32xuD3uIAQN97AGJ81uM4YTobPhqq9+fM8tabPIjzJm/S
HtfDS4mun8l15wA1019ah5lFgArg/4ieDV7seEzLTwy/hx2of1xFEgAN5a4s
/Msdf8EaXKR1w2ire761pDM2RtgJNiu4cSWioHuhHz8v/pcS0IDcCg3qW2hH
NDY5cTsWocB9WZ4BQnSeTEkOcPUJoJ1xzpyExOfmUi5sliV1cVlOYuMlUm9a
tzUgxhNwzYiSgFy5zv5ljMhi4Z4lGVgNqntXReoKXbFdbQPqYamn3D9XsXh5
x2WX6IsuPN0uBBKZe21aGpNqM9MTAy95o0ZuQTPOb1K1Rum4+OO+pfdT4Lgn
xQcNIydnS1md80d4jpkE+aThpRUCh/sywsDSAwSUiUlUVXqw5RJ7a90d5hDP
iv5KiYmkFkxF+ivhl6u6v4cXeCxl/z+7wSIBK/a97wnKugGo+inUkYnvTYht
3nHVMEPVbb284OR3gFZOzswdPGSBIDRLHq6VNGYqjzsoSjxs5vyqQzGY0b+4
/m9WIIHozNeuCpmB35xbq+AnZ4Th70ikU7uVH9fHZCodpPZ2Qzaf+3KtFyag
e9mkVy00SFhdQfLOyiuVV5x1XEZb9SRE3KwPo2ap/7vpA4OYMy3GaCm9qNs9
vZu03jkOaXeb+0J3ML5F4clf2Vd6emuW4aONVm7oYppCRBeoUwbKU+Df3uSF
yQOGWSxJZUvVU4j2Zrc8FGTKUq0sWDm6CzHIYJkS8to4xbwJlIZTUY/PYOoo
JYmGXWYgs/XvWZQ6yOQBFkgZoAfi4fSL7pM1IKcZfRuGOHBlpqX5+KZL+3o0
7W1qJU4jLyZ2aFzkUfs4n2+LcwkcPh7uOmVZX2CtLtf5xUMCtlfrDeZO1iQo
uRSYlCIRcT2wqRTrcGP+84Nn/uDzTwMBmE3z4JkotqCgiG+EAic6I8rqPiWZ
346AyNMsipIfhWIq2Yj1fQJsntbrMkDWkqevhB+QfVzuLlqKkUem1LD4buEy
lPRhuEbIjCySa6zEczvb+f2zP/rEmqTrhQamzy455rJJ2ZvKf97Z8A2PDb4F
MMdekbjg7PVmQagqCf/VlizjGeP2BKuwzB1aezFQslNIrkomBkkX4l9Q52wC
p71jTTiyiMZU/rubxK5Hj9XZyAn68Xz17YnAP/8YbiDoLBAGntayzBVlVZoL
DmxL/fMTcSGMeFchmzno9d5Usd55QWw0y2qf8jU8KuZNKwgGsEO7MyxYQmTr
hE32RJCW6ag5rOaJOE88IBYq/t58zU4gXQU7y+WZpwlqdFTxv1ka3ldqoSEN
eVlhtCVEXpWN+L2YB1erMKcIU5SCbjLYylr6dTlqoqZtF/h5ZlwgqM4PyIV6
WzpaOqA7netbT5QhGl5AnRd6Fbnfs1GYpX564TQ2dG9GFDfaPDdj6fwh1mJD
R9bBvb2p3W2HdvercPzHlG3C3ZIqwqiVA6cZoEa/M9zT7rqysCv5Cp88vNlN
4I8HMRr59oRAW+5t9hbjeouZ3bW2CuUrIMTioEKYSMVU4tITcCF5JCsGfwoo
c9Fq/aSZiyuSSkklQJGeymRxFgHw7L6gyKZqk7GfMGchP4x6iaAm/gA0kDTj
sNGrA8vyaK6JxBQ+D7fDPO0BHzRnF6jlneB4rV+kasUWtMhWf1gGvdig9WbF
n4233v912xKrbZ5g9vV8FpxOa7Dbnjv58GD2NRiyLFjpc3vT4Mv0sBR8xNm1
YQ4DJHh+5T9m3NVyDjKkmJhdm8+PMUOJjBEt4/TGfYBvBGKZaZKPBtJcebMt
BsTz7hWjUxm2UJjt5Rbw3jiejoJnD44S5h0/nn3z3oe7RPlz3ZUuzpkRJDG8
oIrGrWJc65GguZhR2xh42maBft82GsfN4JcWsj9fLb+IV8HT823EWmH2zfvp
Jv3B50cZmJaCMB9joP3zshReVr4KrtQ+RJ+pVi1MmnDXeoAvGwUqc/dkWs1u
jv0rBivZJ8+geolvBzyczAJIJl3Gyc2qUzy1Hlp9y9ZHfCoLRPhOOBFksneH
d+czGTPf6zbykZrtLwLjxRgL5tuwDWq6yUgY16jsEj5385Aj+WhgH0PV8UnJ
UE6tLOgoD4m05JUAlLPCZdD1vLyuTd35TDA9iqJ1sSEHL26KON4HRJcqwPs0
r6blWWD5hiYtAF1rxjd48Z5222caImoVc24MGHpAoi8gzJ9iuKsaj9hgGgnw
NhbOKqOlD0OxBpYCQe1mPr5klD5lVcYmCVC7vinFiXcZ//fQvaQ0B71dhJad
KnVn+p4IJahTSbiL9Px1CvMloeKIEQtL31du7IlF/jYPoIVHonrHKJ+mzfHF
4285QutUHmxz1uCQfNB/CRRNs5i3uWbW+wjj9Wl5fjTug4Y3rI2siObfYNQ9
PeS+b9PD5Hz0NwGsvkqRqEPfUtQIBOBkzDQeScdlkt3pQfKPw73Fg64KRo4m
r5UdH1J4NhxY08btQaMTG4CjxIPkEBFhpQk0//5mI9xD7GHmX9GQiwyHEhwp
HH8zBYJeoblobUv7cwWeyPKchAP9ZxZ0bAHZE1MyYomZg5LkMHvQha8Q9d2J
SkvX2fJXJC9sWYiFIySAiHixIJJc6W4jAhJRTKGw8jrF28ixhRTdMPwPDViy
yf4zLQSWsn21xP/HDGR4nUnCU5KskZoBl+PbfM+bUgeBmxfhG64szCyIiAkT
LRWkeeOISINOWrgUyclGmoidF13T3MUPWH2Iog/6JcRm6GHX/9ZDB7+6Ke83
IMXCgf6fX/Bxh0A6OxShexDOEw+tsmIozHd0b9GTsZQgPl8SQ9BDeUdWlHSC
jU0RC9KW6DkQ9sx1ZQWq1XfntUd8lTaUC2MzwHR2cLrEtZEr1Bh5lzl8jLgN
eBPvDxLU3WTPzZcrj6H7p9zzRzFJRkVu8gelo9hJvB3fT+OC2BRG8WUszFZ/
6jl9GSbL1OpHSIETE4GrRVK5KgIGBYpM9lC0by4t7YD/JEQwN93f5ie67jS6
BuLuky7bPyu/LXDaac3iGf2hmdwGE7G0w3tSzrJHedu4ObdoSq0s4QldXNd1
lZdIjMJpaFS5ukQWCk7x4dc1U4lmK+hnKYqr3de56bQ5rqOvMlEKllDbmD1O
2lLQ90hnNWTW3Nv7KoUgynlUo3MKzOnej3GeJxBstVqQFklCyMAkr3oQOQnV
EOpGe/gBigkER+w43Q+svHSj1SEPVHaF7NWXP7bMjnh8tOT1td5VXOnElqLi
SDWkAjvMHI3POc6wZhv/LCnIFAIlk4lRswd8InJitt+nBP64Iq3pyJvsoHXl
wOJLSgNZZufATCRGJ+4Na4WeQzN7kzPoqj+Pkbrz0USo0nrQ2HTSafFfMEqu
tljOVwgPlml41m8wihcxf5n9ER2mPyrwqgVzyLRlJ2oi1x/0Vyt6DVcIMP8C
yBrhL8NZ0sJvgvcO5KkjUvPsrgoX05diL+XwqC+6+GHVOM/peqZ/6/3Dyizu
AVK/CiBFBY35sCRZmWaR5iePwmTeZEC+J+5eO98L56mtbnRV+bNlyhrNlkN1
FMquOOCGJVqXKMi14y3oMz0XqrTizNvhY0h4/4kfAKcsSJ/vSKvzU5c43RnG
sbF50/69Fsl6lE5VvMUpIdxmMhAJRtxmt3snZN/2tYSkN2ARStnH0rGu5PX2
6PsOFplPdZj8iJj2a2+3jAO260t99bqM8eKGZF87AsdFiS4LkSLOnpLx13ko
dRVlK2IZBp3NlBS6yCgo57Pi9DCz8o+E1iEmQkeIGFXQ+ZnNMpuQ7WjZUJjJ
h9SZ01uYWS9+OfuNLp7DYenX2E3YmeNK4vroI4R08ZzdntwY0yit6gLJhlen
CObbFlj2jwzKh/BN8M0YBMc+ptA4tCG5hbBYb86d3e3t7WdwcnDhCLlJiScB
Ds6wtSUUXzdzTyyJ2K/NXmBw5r3T+Fp8+vY3ZqGWw8mHFegMZr8uG12/vfNZ
M4sOFKFt7H8Y6HP9PwtI0sZ3GeylZpWaHm4DEM/Ov2ZgyzbiPynYS4bs1oKs
p/qStYwvoxv82a3ldA7UQeH5f8/EmpGyLVKf5p+2zmuue0+KoYtxRiORN+18
xxZX37LJbHXKvC62QMiDVKSQE/u0tEAEtYkkjf1VMuGIFq9rDfFPjhVqNpvN
J9SAJXDIIwjRahcF+PTzJuTe2DzfneMNVKPo3ILxPb5uNqRWhlpHNHhvyHkQ
gRgl2a9VAw/fw5ji716bxHmwNp4aKJkq1dxtQmV+RSCjz4OBftTovmsuQ9OU
1Ag53oVZ/wBIqX1k0snQbi690TzqYswkZJVmouxL/ZfLCy/aK4N8ReHuFe0T
5hftUFWR4Lp1lXobsT7f//2c0sBWIgwjbUy8PNs+XvgOarkD+z4fHoIqB3c7
i8bxBe6bztaKPlphadVmsIkjSamzuwr5iBICq3bnguAMItFhwt+yGUaafEVy
ZpSpw6ShiYuy6/BP5YrxDPxyNvvtBYR4y4OWA/wCKTgzba4HxnPgeH46l/iR
wfGv8BjDpsDPb6S7nRfloGuw+m01tJ5nlt3qoD7b9oEEW85uY/y884KIAwna
DyUVcWScwIkDbHWnGPZ69KjOakfozZami1Dv8SHHUslQjDKo1TyHyBGU424c
Femeoo0oud39J2mRP0XJWkVotN4QIXFUgA2J/DqneTOU2uqXwW+Emg7v0eOC
84TSjZ2iCYU86kWbucywstn4IIBeeTrZHRI0cliZlNi1Lc8iT9+hWA+m5ECA
cloUerEmEVPBCAKNq7RSyTMTIV5QbksuwExvSdgrDy0h01a7hbMglcVU54pt
hFTn7/ZykjdVBGDevRgvdCGwgT1xZLuz1P4GkBm91S67qv5uK2rin6rlQCHj
qa+HKXft1n08nAnEONxDCNHAv8DJeLbFgYdVTVH5/02XTh6jQ38yYJLYrBkH
yPgCVho1OFFai9FrTxbQTVNaiPD+TYQLeWrv4xU3xQDKe/7JrNasYQfOGKhx
bNsJS4I9M3y8luQCpt/PCrMXfve3LNGVJ09dn4VSAgAdm5K+CW2R8L85oZqi
c67b1OzrE2fN3NVY7iDGyTh0PHCNPFOEslwFgY6ZHL+iOgu3PGNk1kjWOy38
tEWKl7y8hSwrQXd/gApNumjtqdbsIcZpgRuXjRq+R4/RgvjyjktVfoHAwnLG
EBd0nzNpJmAx0bKh6NempajpcMF2UD3KG/jEKHneisdwHK9tgSRJBmSTuoGY
Din0U3BldVTkblpamWk3uIbRpdNCSXM12fj0m+OefL4XrLier9kDWfcB1QIA
uiTMFc2bYpLTgn6G2PpsHCo+s+NIy22VOkkUBmnMTjGYP2pmwXm+Hst3fIwO
a4O4wWfZO6qQFxzirbDKuSEfChecsqPvVb02QU/8VWDd3dDnRcQiG8ZzaB+O
3fx5bhV/eXCBXHbAVRjl91fA8XOXZyk6cjkOwkolvTbO7BDKBlqaWH7c+PV6
uKAEj3HVwIWzt60KOZI/WfAvfrfPKSa8enevvqyqJMV+73/tVVCLBdnR4/IW
5Rrmz3nDB8uOP0H/DUdQlXaBHmJv2nJCSCSJuh6QE5ljwYEl0p3eqZqoJuh1
S2GXwkAIOEu3GS/BJ4/tvrAKbyd4BndmEtn7P47hxcwLM5Dyv6bEtFc4yIJ1
MMCyG+Q2YQiPML8aDqV2QNnQelnFJ+x6wGKz/j6DlenI/3NHHTh92Bhf6muj
lKJeAwRYX36px12FMBnIuJ9Dhw0cOMPbMfQk+U33uFC83PRWTfa2D8Q5NZ+G
BfLfMJfHfvRSrRLEf0CZSFDXsDG1sjELDCptM+pj28f+SqYtafOTfmOggY2l
sHYLfnhtSS7ezdn/ngSnr7DRrAzwBBDNQW76we2aUZIat2mbRk+I5FsZa8kH
gvpPx2yBSpIZS/JkL3i/i0PGXX+xGmayGSXzBGjciN9Y/Ma1qlyGGEkMX9C1
VnLYwzYEVwo3txr9xAAPIbQdz1HDmp23wDz6JpXtn1E+xKyrZFHJf3tIvdmD
XY0aNRbRZlchR/dfqS4w6JBcqFOzmom4j7VfyIW1zJD+uCxVhzHEP++79gGY
0wNi8hEHxIb2kkatJzI2fkEaJfhvFL1LesHQE4BLPA/pwVq8+3W5R6iNSVdG
UkGaBybGbB8ed7v4ItVtYBydOvaJ7O0dvxwoW1WS1v7R6ZgpUZpqE1E/UlM+
kXKCG8HiOd29r56EexYss0fyp+KL9E3/ZUBKhdJbzhQRfcVsehAu+6IYIsjc
xMPPFSAULwkAXhU3LMM0BgsOjXQjoGpPD8qWleTEyOL1CBu+1zPy3j4aKFsl
e6jr7+PCEgERv7c+HvIfPQ+NpECAMJbynQqskfWiGAT5VdOSFyY4QqRBTn4J
g1X1ZWGTVzrdB19KJNRp3+lHKR5xQw9uvqMLco7hObSaHTXShPt31rprBIAj
YUV1H0x4r235P/yIfq4rmGIPSN50ONuKv6ZikVZOOoK2JLJbaO79O5eVIrTG
JYC0NmQUonFQnSkALA5Rn8Y9KyIv33xt+hZuSgF2N7XZc/ulwieL1Nd8W37x
3TUyuftuVFYy5HRh5yO6sasIZwQ4WzJVEp+tzp61Xg9gTjtd+yYFbM0VBta+
ZY74MXxMIq6AXXlSe+ZLIAiUH433uYWRaFSKzXqUs/mPiVS7HFDGVxMUrhi8
auyrpDL15ROgZ0wWTH7Lp/eKQS8WdUeGbF/GL7Y55cBP2Qh+130a3t0HK+fv
8unlDSg7p4YLsa/I07UYWhFwupNz4du/g8ajZ7Qx7Dvf2RxDFmbGJVN5gcYF
Bj9yRSnYzxfs9JcWIoiNrOMYQo/D6oBCANAxXX0TzeyoiNsHLgzD5GlAY9Om
2cQ4OB4pRlp7gsttuKttRlJ02B0EE8YmZahAGby0S8jMblN4e/0DNNLDPU1N
5/PZFoTN1ToRvZpPnHxS8JPgkTrWjg0ntV2v7AqZpxzferfZyk5An501OfCl
NRTDkuKNkz6gsGN3mKh2QKFSRa7IdHjpslWtc+ShvfwMBZIylGVWTA00JRSk
fdhFzKmNzVkzxp1jNWdaLIzNjGtMDQjkj+MJKUWCTrt/yiYWXtw41XWp45/y
bPmqOnkRngpHtbl9Nt7ie/zzBjOWVKmaVczVlT/3xMmdsHVCDClfAKnOefgn
3NoVl1UFZ7z1uan9PSuLHw6sQlKYz9rmkFkqQ1Q5EvXmrkTrWzw491ZX7j1S
AN3GD4wjEP3gBVzUe8Cf7ZxLP6Fm83/EfNveev0HKfHWMbjxMwvT1LrigjF+
lZDWFHBGXTdCt21uzdv/Vd4LYg+W5wVmdKbvTdJxUwDUhcLslGX4lznhKsob
GmFbklAd9ORHUL2MxqIo3R+ReNIQ89+XczVSqiD1C5XJ34ImOsDX+BzmSgom
0+7dZaRvt5Ttw5oH4A/oDnPovou47d1pqyu8CD4K+b79WHqSnlRDKVg+rrXD
9LTwosSQAPZqUKg174GUAndvct3ZGRkjiMKz2RvCKahyjy/4kYzlu+8I0Cmf
R3B6yzf8L1siRNh52gs10xDJvseVe4KpHt90qJ2n7ntHOrVKMFciAWRe9u59
KgjCEiQZZashzbbGVNLs4khPbOjQFOyJI8ppMatp9Xv8paRkes9mjUqPbwAM
Hb7IylTX06CumrHybYgEmjawJH967/594OUy4xIGQtuEKot5RZqDWydYrytU
Icy+GQ1llaDnIhSuJ/zWoHC207TFe++kOiyQ3znDn/aoKJOwEz4mx8A1uQG5
bxBSghZ7dCxyjJAG6YFSFbQUwQ6zZ8fFPXrGhyo+VF4XdRw1kDzxnLRDUWr4
djjSkSI3yKYrh0shA9tLTlCDz8tVECQ3oRGme7BEZOxr7Cx3MG+11mcB4Hsz
vyPwc2zeJdYdRxcObMYMJRSawzIw9xLlv8J+f2UtPXxpRyr4+VIyk+nrWn5Y
fH/P9ixKxznAE57qBqZGAG1LiRCnwXpn13QwM+UXlhCyyo0qjxRCujvXIO0z
7OK0Qyv2rBQCf2CPNiEfVPGKl30aHXz1Vp9QrewFQiuqDoehkUmsoo3B3eUb
WXmM2elrETMaMgwL7+Be+E8EOjONTuXFswR9+quAyHWgNd0cpcAdUZOZz5sM
KMjpvtB5Ufr4chIQtjpHj5kuCZdBIPQ4Z55F0vMwhgjXV+5JPVy+JMdmWxNA
szTKklVVRUf92aWw/UMxO+tJZAn4oYaO4JL++ogZU+eb4/o8Cq6+BQwGM6h8
1qdgNQZ44bhBaQF8B+D4n+NZ1WdfJh4sE0wic8kLaCa678pZwFldhd8le2H6
exObeo9cBVDymO/+UOPAQB4U2KQtlSvkq6q3Uh704jQn2dE/Vr5VXnPvQfeK
kc5sas4Un9uQn3wBbSkwJQnIIwpMzWtFyYsQ/s/6xpg9ze53w5H6fKLKrzuN
WnIIFoHpY2v2YRUFnFU6fT92ZYV6jJr2C3iMFdAoFhUpLRW5jj7KsCPhC+R4
o53hrk/m9DCcp0YRKAi9dVPFRnMYcHmZ69J04MFoIHDqwLck4DRqZp4ZaCeh
8wY55+iK7f4IfOO6U4Yh6MW/Thb2F088tuppzv2P9ZKZ3z/p/nb4NwEHU0XL
lsWjxwbPKrtoSlyM7Kv7VDBz9EtA6jG2chZglCleEmLcecLRuYQ3wRnC/z2d
rMB/sFB8zZ3MEc+85xsyeFAn574Np8+BRkyqxQyH2xaoraXSRYnnG5SgBx6y
vSEntgBoFOXB39/05CPXWPjIipXz8pms8eH833os0rWGFf7YTjQ9m4qxNqbq
Hpz9460f3xTqzF85NqSxFSiRzi3rxxcbqiWBAHOj8elR0aPnxnKzcL0wBuGZ
DxDPPmZ0R94EIgJxiTG3nE/ep1YpRwDDAvJHPINB6rb56jgpl5lPFktoaXSM
uJ6gQ4Ja/TOtecoKtSrpod1EraVs+1Ogyig3sDzhPz2hUFlFfgGkSk83zct7
pQPwEtOFk1ujI1wkYsrTCI+3I2vhja3944nG3VxIPJUhvNHJGf8cMfVw476y
6hoQN/TCj38kpqT8/lz4BKu8G0q/higdvGwF2Nwru+8LvxGOOaRcXbTDoBBp
sIyjpEBo9L1J1VBki5UqC0HD/ObHiO/DCfv0XRHOvhzUveVyazLsvjw5nwOo
sLA157KeAsDkoz+RFZI9WCwgz/rAQ7qIf3RTWp2oZI5iHtT4tUipUrU7COWw
QooDgbZdCZC6Bxl1WxkZ1HK9rgek1jaJkD+zTkf7idoCYapRczxt6zqIyYdI
oJvp98oqRpNngPTfFEGbJF/R0jKEeR4MLMuFAwxCShDnhCjWxcEsNTIHV0Y5
VV8rnT+nqiLZrKj7HHd9wojRFhqbgWZA/GS3JwjeK9bQ+dI6yNe2DaFolXck
ItZPDebQAwFyEKNobRupZJ1fzFgUyDStU/oSM2Pubwqv9GmAfy8C/9L4O7dr
ReParYuOteszDuSaC73thowD0H4pvpYHE7fWNq4CtXor7LTJv4Yn6gLBYtMq
hfj5NqlBSl3n6u5b6Fdj6BO7VMPR90iu/71pqfadcPn0txZPjrCpdg3NFNkV
srNph5nltMYA3Oclu6eFgY4ijEqjTlFQVB2IRUJVrzyZHNontYxdACIcMre+
YjHCVDbIvwNSl4aqpl5dfs0iPgxvipxoAQ8AaeAkapIZkKyL32noUXyBJJNQ
y+uWqvDE8TOolj30/louBHluohlGueQGjSIULxMGFFGU9LhulMYp6pFWm3Fa
lItK7XymKgyoSm+lN2bOC32gNhsIK09k+rEMsZ3q2Lve7BkkotXxbLn5gvIz
L3ome7/kw9V7F/PDVZO/YX3Gv0xmjbWjZEQYZ1cqzptDHk3jObn1EBpjVNj8
PLsCEHMIsw+uUBshiO2frgr0DF0QT+X2YCqiqT3J7G7q6BK77SSSuFDM4/p+
UygUOLxfr1+n1gFoBxFKG9fFoh8WRhHgMo3D3rIf+6fXeEC4KmmVjU+jcE/T
W4qMXXnZShIaA5Xck8qwBurOhgWDsjxah56WhzMuzkneYsTb7Gsgqsev8/DL
TgnOjjXoZYX6K9NXWaFIp3NMgxgp0cQ5OjmDZJFDXNPanpisR2ofeV0ai6cs
7BPbKThpWU9b6Fw06co93Dq5zHPqvzyiIookKGZA3fJb8ztqIGVSmyaE3Vkq
W1zy7QlwiXUr0R+ufOyZW0iC2HIAsmFihO37hMzcYefJaztsJrYWRjCaE7j/
QYotJoqBcMHgU3IK/w10JBT4BvUgcL7BXOOSvCcDgvpm98MlVzGj7tlOWU9C
lLKb+D/xHIyLabURWA4aRZ9fZwzaxfNnMfYW4taYLPs6WdqxsITtV6uAg4/U
2RuyfJiZg2u9iKGp8mut7y8kUBxEh88MBjEkAgbdbCF6ljIWJLeMVqhdwHdm
bVZiM3oXykiVWgS/t31VQqV526rKqZ+jpk1zKouxXQ6MIJtGGAGlXp9IMZmb
GoY2hP1/4RubPEAO6353pjMv51F5WQg66BrfKPAWI10llQEOYgSfe04C4q4K
IiyAt5HqHKY6OIx6G+R6UkbtrPwDBtq4LAyeQ+28HEi6Q0jHdHnTAlTsDbxL
p7Xq8ae9qxdyLNylCQDHS+XuvzYKfxPLW8x4yn8a4MxabiXefLkX7Zo6N8a1
tJMslE8Uaiee99ogSgOnwpNyuzcsjfu72Kp7qLR13RngvJiWDuhpuES9oq3G
LyxdHmDaslJKiHj2K2np2bfwiP9Xfrinf0RLeTHttBwCv3aksxuT+s35UhPR
RIpN+KApMr4yV3QQ4YZc9Lfn8yD6X03Ot+qm5TfXrWXaD5FCGR5sbILkrsQ1
CHrwlu6C+TQ0ZlKb38qjS+jhjRFvEqMV6lYs+8bjaVRwihQU71ZumM+niIGJ
tJy0hGdgcO6fM4mQkRTdaqC4MIe/Iibh41EV8daQ0KI/IJw4w7ij6rMwNRPs
EDx/c7MsFCBk8OheeCb8vEGAs8h0nOAQjpndWIrPLEZNpyvup1MDeZ0IaoG4
5mee5M3Y8rLH3fCBgK5G/1tJiAOrua1HkW5ykm7J+lHnE/XwZ8T52sCNSOpw
c8BKxgzKzzlONC2X8PFgsJ92/5pQi+V2Oa54CnQgkjlIyVDUsCmE7eUkUPyX
m+qsdUj3HChnBVUuKnllz8lu8lDzjJeC348Vt5bCYsGf8VOtL5zNJSYp/uFB
eMQwR7eUP/2x02vaUbl6eowo0MNifgvdlvBJpekwnIjvC1lud9ADjydI0wPK
Onu3BrF+aM0HdQYSJwUoEnKLHnSvDvm0xiRy0w4qNDK97e14Zl19tmINOUr5
DUDoqWBPH+SDQCmUQ4xsPQ5c6lpsV7AnPH2v/Ux8D4XLAICGBcKLX2nww8zZ
vxCuipe1iKH4oW1Svkf2eT3SDeZ2JfbacG+edmpWKERWfTsit2sJlVzCkiBd
j9XCWwX+MTmFYQnAlXTPRbv2eGJGS1Pbw45gWeALmZbTk4JDsaXT8lwl7ADe
8aUJBDOxGu9xiT6e5mqzNXOoTsap/FZDKGILdNPdpdgM5KrQ5yyNNb445g+3
N14nON3mHu+VIAxo71jx+5sP1znGCOE5qYrcSbLjalfvlWMsuU1FMSaEroCR
jaHFp7GahWzBrambDVYNbdce47YgNnym7oF2MH/D4VoWgGToL3b7re9oIWiF
lY+K56/TV1XzOs9axXlp30q1WwuT8NluounTLAzVo/ruNPjm0aCWCbafHs3J
j1IUiCLsUpAEsb0cWuMnEiyjDYEFEK1oENIHHtgjQxCikGLwFNyYL9Zg8ibe
LzQQME3es8oxjTJARy/8prk5jwP7qff6AznJb2qMIswlPALxymBr1LzTqP/u
gRQYkLydb+j33v60Ma3Lb4BX+KSRqUE+igqLTN1sFJ6Ibs9UrcpY/2FRUM9d
HBKctIgWIoPj1+L7nlgwgunjsdWJrDznC3IK7JzgrUDUc+fULg2fy4yRwF9B
c/lXXlEyUXY8C79PUvMnxM3y+EOfNxqcJe4rUYYE5mRQnrpWR40K4cUfioqO
Iiv3POV/hyLPe5QpuuycMlcbcGJvFOatN0ZeFnA8cQ38rAWFhlTu+fR2TfQi
tY+oVh3SdkDNugz5mBNHzyvzN8t280LJ3EO+Ld1OqVgwtHEURRc0dY1ou5Rb
ZscRfJdyI4NZJiinOa3V/VwO8v3/UX/4wUWsRIEmEoSY/+G2YaezvdxK1Wh0
BBoDztk3D3sbXvMF8jvpnhmqDlglpc8468c8afAmaeYm+zPbjHq4FczAFRlz
Bv59aVW7puNZb4Yh/s577k9V+0ucCINdG6GA4Smhs/AnqzKduSLuTaHUT85w
NFTkSj82+wmyxKca4oesA0MguroESm5XPH2NHrxG6avkLB0YPgYx2VpPY9KR
3d0NeDK4PQ54wl4KpGtBRtLYrpMtHpyA0DLqgfk8RgTNmaCJVN6/SEweDO88
m5NSCQtshY8eClLrEvS9+d7BrpEDq6BrcEexXivgQS5KahyEhMZkYIntXrEx
Mody3wFKoRNgz0vzxZxxAt5IVLWl97Y+o3A71/2RVaCW1kZOTxDDeAqpt4nG
Yt/vwePXIKRYWOPwpi2Jsfcrb+sXhplli/NCyHAYvoj5kBk4ZrHVQzN+HmCl
NVx9EF58aiPSpeDmX+YLeDyJBn3f2h+MatOFQO4l6Ar3MXuib7gH/sbNLiAm
OxbuyzqdoxbXgafVr6KQV+21HcKBFSYUVjg85gq+q4Z89s7gBNf8bfjVKPyt
8boTC1qBzSCKN2PqxGKqB+aJohvqUC420lhHfrd7vu/LSHku1QctZIWyjt0u
omZPH0+6lfKp0ZBV8O6YAW3h+vTthaR5XCaM+XqA41pLZ3b9mnC8vJuqp+eF
caca7EFMYWw8ybDEgbmJvClR4J0i0MUD15VwedDBaA1AvXIfREl/sWYrsdVj
f1NnKPtRdT7UFMecql8UbiDAKrIvr2Unz6JFM5uuRDsmUyfVBGh4lPUQgb2H
/glFR2DtDrEkPtcv/FnwYHkRGRSgk2NCJtC+gPUjta00sM83iwDQ6UF0TxlH
hrV4w5IuzLkQqGAWAaXHpD5TUV/vYdffVJPakPTurblf2rCGsH4Awz/zzQGB
dWme/MmqrnYUahlO+878/iPje4EJJ3rB8SIP4AFClsxkskKp46+fePYxIp4F
MMnrXu1QYKTv1Uti1+1V9CCqDJnRYav1zwMJMhFhRlFabJy4DL6zkizXLSHM
uFloX0yBtshOEDNsXpEdWGwh/w6bYX4ezLxpD2CM+Ck9NJH1Qxk5Kre/GxBZ
8h11JCd/e3441dYWS+JS5tjKV4DvvrewL8DNL/AWrJDfLpL5UJ37/IhNUItL
TjqFSUbOvmT0jWkQhPOE69MKymFQwc+umGfyi9OtkXzb8RTfM48d8yGjwxb3
V1qZYs1gOhk/G1/JnGFMLofpTHFHGt7CYigPyNZCHWPW5mUxtkZP9nIJhfe3
hS2NRq5/jmPOWOR04Vk9/aeDTYFfqhymO3PdK67dq9+U+Q1bcyRi5ohQh1BX
LpobTcSE0ScHfiznaJPfvXFfnMjRXnybKgYrUoiVKIKhzs40mis57Z3d6Hk8
vanaFvRwYtmagXbZPw8rnIl7GE2BfedqsMrQcKHItIVxZzgusVVeb2OsJ6tq
kB9Qy3C8KsB/kfVkSmaU43X46HcqTwyD6ZHkVEQUY1qgBAa2TzgNtz+aRWDE
+tiL/j7H9X9FxcrfvwGifUNIf7BXyGWSsJjths9u9lj0Piq3npYXL8hIrLMQ
/AM8zTVLPr1/WPMLynMLnq9LZF9Ldn9F+iOlyFxNDgytVHinGo/5cWr1g5GW
iFgqkpDUy4U++yFguoZ9V7aVx3E6QF17Qu0ESAIZ+XAtzqFUtF1xf/frrM36
VDbrzw6Vc9nO5/40PUyUaU3GbLM22wJQgzS2nA50ewLWGZgaaK3Hg+LuMX8l
PDVbJF3GueAvsVEmaKOSCQOKZEiQCjqbwCfX/EG7zXIclGTrgKUFd51knaVX
heINBtqihtVx8M7KBJo+jX1CkCPm0gO0uW8jYSStG3GNkYRd8xMinFgy8Ihu
fp7DF+6NWfQYZikN9RwwlmJ6sHRlrz9uiVUcrTYMBFWxc8bh0GsbmuKC9pOJ
FS+zj9LtNgp4u+twtS8+vTaln+rizUaFMM6CeEICMmKstfJ/0ks1jfFpftEp
Dnz3CfL9lPKnTaijH7JS0hv65Rba0QD0CLigCFmJQusMVQvql/1+O3cz1dlM
MvQfusUfcaZCzw9nKkJe8+OuT7kbhSJHvbSLtkMZaze5cTBaxsuWmEOp+7Rb
05FhmWnvy0Eq7eO1jEHPQ1UMCZ0VSVLFBXJDU5V/FcxwdaRhdRadU0Kb3+bl
/cO19FeXJPfu3VlxMRTlC7IRv9c1QBqbrKx0+GjjIx21QF+DJmhqAuGBB2pa
LZBQcQp730T47CbBhOFbSr2A6PzEKcguRmztF6fEWhdLMfNleRM/GRaK3oh/
FlTLZn2yNaB1nwre0NhR+dLhDs8L2xJVGZn8no4ZPBy5RzFuVbpS3B9HT6SI
5oSg8xl0smjybszH2RZIzw3TbXrpQfOBiMOYkqa2DCZnbvBWvC7KHpJX92iU
Uhv7nWKoaWGoKuc/cDSx1u2NzWC1mTtEf9TUjR4aMZAHjQ3+aPZjHJxd5HOO
zzyjQl0LHmxaaWGumqCFCXeZO4HtZZaerXOcrAnySd7pu8iemnhaMCRK6GoY
ykkYR5mMhT54YuaL3paBj/7NCq+0bkDKxJtPIKtiqMfGDv26QpJ0XQY93q5/
M+a1i58H9FohBdzVWEarHMGBqxvFz9UDsBMZjOYQuNFidFC6NJpHlIr7eIqV
TkLc/v565p2oQ6AjTP5EDNyPZq5X2jIcJpcOdrUUnaoEnfCFb7xq+A8RrYFg
03emClJpFU6OexAb2Bp5y1l3noy9+gAqPJNyvx5Td2w3NNH+BYqwRHXqaXq3
HLSW6E6GEFc9v7ceSAA2IG9+h0paphmPVaYsBVlNcPbUxhNsF+OaoinOEV5R
h76ikJ2+J70hetXPc9udQCpMEq8QjPjsj5XBTkmQENkCWRErtuL6xoP6BqEy
7PojZXsZtQp+r2Uzf8kKy5gNCiMszTQHL8J6ZzyRPyF7tkH6fw7Pvht6XHLl
He1QXaPR4GvELsRaGRuJYcHMMx0fxqMGCyKplef5KLeXsSOm9WbuZHuEE9Li
GT+he1RluivlDm6YfeZJT57Z+RVbGfAt9GUOaQSlqhXs9POGDaBi5Y5iUnvO
tR2Kpshm1E3ZEkd+lUW+O/rJ0F05IFgd5fs1XqVGOaZorCdl7oABOa5EMGOV
h8q+d+1tZg0hqkvR4E/t3b3o1oU+FA9QaGik6IG2VynfXrKZPr8Y+BQbqDKZ
Eh9/74ISa7vGbb3pPPkuezay8YQmzuk19tUBELRF738tesCH5IimSEDn+YTX
mfrcEDaOlKTlSCFy1DM59afYU/xqbXOU7bbCz20JoZ6ltTpqsUT1i5LQB5jf
+wMg4740G2v/QFlLOLBw5VK/9YgoSOmTvtC4gnFbDPkr0meLW/ns/4NVX7eK
xeXeCOKXNw06RSb3H8KYuqOvezoY1bkCHyzsoR9pj/bZ1GZODU0p53VTRfGT
PrELAKEeFaahZjXHfp7eDBZirKRLAhDwXxZQMFCL9x5n3kZY2Msk4ow1Tbn9
AeY8pb4cBZIllyNMUo9jR1eSux3hTzH0izgREqjlvznn+0HLvgUfRP98BwZa
8TuqvcMMn3ODDNWf1iGXEUMXlYLAb6LcO6cw0kHGyeWdONlzlu6vKPtfZ+yp
g4SMzd8HBNje62zoNTWhxvAUIaUmRHLqPLBsT+0/88NShRLzCFnblwmhu1VL
vf/aiHaWwyCjdEoxBsrL8bTllx8cASPJETZS45OzRyULis+VBROvRDLlsDGk
PYXVWBbLTJgw8YuDGQS77J3GDD8E0XBNVFmHOGUFPRx7h+6eHjPGEazaxbeY
vatEuyi4/qkSROHN4MPf3/fJwRyx+g87m0TBklaKDjrKvbmVZEW7oLNdr8+M
+/V6pDzXvENr4kEGOoUnFEF2+Wcs9qSLZfnUSc8ydnC4aBBM2cfXPlLjZP9v
8/dZNxa9nhFk6oTfytoHWRS3TicPjvl5imd67LDKdTcNFx27nGTw1n5f0nR/
PhZVl3mmn+YKs8wQwQ80nmooT+pvAK2dsCt+oux1r0cO94pB+akQM7T9XKzQ
Gi/Dzq9/q1oMHfPivs0l+HOZVg91FYu/P48XwPrYIP2q+0v1wmi4+PFosHsw
S3GunSFjH97oPyBFsbrbzx/GcEw3mYnSXDxtl/MA+UoLUtybxsAM7IU6QARH
A/pqeJ5x0JO1StNKbiKZpnrwm70UqXB0PaF2HyfgkNXbBsZtzzQFxRm12Ih1
/jbaYiKMZxkdTfzv8RZ3G8+qFJ0Ol1jOTVYqCnHoabCNGueWvkzl1EcTcEuM
4lngsl6cpR13gdrRm+MIVz1qnJqkE3F5NRRAsXMsNczaPIC+6xShxbLN+8Ac
Pi874I2CE0njC+DpNEPihlMlPaIMb01J5OVdD7LZYuqdfqCXj9QeGspPJOqv
y7JTWsy8upTWq+ZfK8cpSBkyMpa1ghd5LYI2hoNjCkcvXJOxPjyeo4MoJJAI
xlZ0w/pwlZN9Klb0/uDmO9D6gOF8VI0kBU2PiTfMeZpWb1XOaTOFbvuzmjGt
eaPbvelyaz4pkQ0hBUD+vKAI6Dh4uIvNVGZBX2pRdYFdJKOke537EHHmE8bT
tw0wcLJDdbxRWwdUoORheOQhO0nFtrpjzVW/O61FCr7wYZQ4ZeAMDMPNqaP9
PD+/BFeSovCdz1ZKHhBbfk7zCtA7ciedcG6zY2RkbRUaHtA0azfbTS6J8IoI
wq3pzaz7XVyCVQ1OGDMXR+ajojTbgw3DlX0QogRUP0k1UzPwLkTv8YCwqSVc
maGrea7HD2Fe7DnIHCgvBVtCdXA9umL9VxLOP79tD9UFZ9nkj4VfJwDywyfD
SJbVbFkEnZwpHRhadGd9QtYNo5nt6ajfOB0SYwl+LbqojLcQem7HmAk2JMVP
4nhv94IDwwZrhw8pGih0Eo0fEHaRqkeRfy+GYi6gKCsxBZgvkYXuPdLMNa04
6x/0EB8gUEdmwSNJnuIJ3kjdUStIuFbCVk4rawKGr3Q9eDx46uCashhv9YrG
KurGrab0L9W/DoQZ/rIwe1WhL1U3HjNoQXzD0/UuEXSUmKNxAz2+vA/XGCHC
F1XX9idPOFDwCHuGRzlXqDKjP/4/qNAPMMlk6DsOb4EVgotlQyHeRWzeCK89
IA4P0KW7984dlh12T4XOznZaswo+oicmV8S86qHznDARDUdOA2Ys6pjVHNe4
mlpJQwJAi8VYspFSL4LKNaSVcV5XNyMb5hbuKWQ4tq73E4uVMFFDQPKE+X29
f6eAMNLHckuMEV6P4xvPVfLl+QPi+y/mAjzb4yNFf7nb1guyTJtM02FEAiBs
FMjpG0Sm9Moo3rLC7Qg+fTtF1F1aBhd2PwcdsPMSg48r5Xbnu/9j06GovDDo
gcPUGlMvszg8ucgG8SbqICARlT1z3S8FsEVIPGP85XLK9z0zs8C9rCa4Nwer
IMi5bSrq/Q8rB5WkuA6SRr5/EIZ+GcK8k8/1wjsbopsulj4CK82qA1B6lqVp
alSPBDljjzQuedyTgwBd9tlp+Jm8Je68P0FeYcLQ2ClvSQqpaJ85fn/AwoOw
Ob0i38AM+Vx3wOr8Moi9Py/2LSC1obcVls/eSniy27hlnuf1DjhZUuyQk+Q7
9dN+t82BgixkZntG72XzgKgyeZ6kE3p68gW3n6LX+07RoeBhh8F3JrX5UjKS
CXW7W1PgZQf+6JhPTpBiQb7i5IYDGUx1ZBloV5c14LEigXSq9V2aDBkNEPCh
v4SQeMM+GDUTtKPwhXK5pGKWudS/H3T883OFFK88qJp88Y0bDj3MgK1PgBhY
6ahujKQDR0dT86RuKPkIXSrI4cTGmXh7SovF5O40r3IVmzL5oZ5BlJgEuEGX
vXtBDFZEeQwxbnIAXe+8fbuBOQqb5n4wBLyIloPj4o6Rh8O8BKLK3qjJ67Ja
rjMCyrVliSU8JJE40RRrkJcnNHSuLdfXS9sGcO8vutTx10iXw0sEMJr8jSZb
drmIZzmHStj8mMZqeduK9rgDm/wqUmswELvfHpP/GQAPEQYV8wT4byXk+oKf
Gii0rhO8Zgf7J7OFaUDfUUNkcUMSzMVsv/AwoaFkGsTv3bz15un5V9B/wom+
TosXMMnMzOs3qcrvmtANXSbucbvxOF/0Y+sU/tF56wFph350hlViBFvWdxJw
zx1WJw0GXw0NT6dTtb3ZQvKJSeYt/O2Ffv+QuvkEnE7XjEzMUtvSS8oLfbXv
7dbtFK1B+CdMHiQ5adG2L0GVjyT97iRMS9WeGaMx5dHW7dVgk46YbDH1Yz96
KKvXR+AshYTt1/FVMMPl36sONA1biE7KaHdyuvc7BlTuTliTU/WZZoKGWLqz
iLSJLFy0K1vVKSH5VYWNq7li8tVxmv626XXbb6ElV5r1QYy1OfyMTpiKH3sc
AhkXfAyuRSTyVwdc6RaQZ6z41Cjs6rLLyONOSrBm9lxON+h8kD37HKcDY5wd
nkZQCOZL9jjpusFEEZp4w1UJsV/FqV3BYtD8dZ+xVCBKYnsQ7iRugVxEAz2H
KqB1RqW35CORBH129tW8ko8HxQVT+y6wM/KQsh7COo6rQdOInYXMjmlQ49P4
s7xuKdx/yjvZdNaZ6uBPBg38PS8pv0aMWEBpgMMS4GmrjuR6dNlTPWj5ccgZ
nqL9eZ3A2g9NtAQ7jj/BDVl0Zr7zqMvVQeHtej3MJZugRwhKvgq0NjKIdcoL
xy1IhA3woAX/m0WOClZmX9Cq9ddMGNouM9xKSyUL4mZ9ADGlbQSRCuqawsCP
8WX6es+fgqd94rO9F/BzJSLfd2AzriY5Ln6p2vrb16WWbfQm76idJP7/i9Jp
u9v5RByiZKZ/Wfp7nLfnCPvlS5GsMP4FESQ1h3TCxzp9nIXZc4//M99ozm1a
rHVbSWMXhz+G46vuwOJv5Kk55ip4hhyi7DQI3wmyWZ5C4PthGa2BBF/Fdxej
X43p9OL/L8lIS1vZRhw3gVZbja/Z+SfWe09zEkyKRHkhTbNxfDx05+fWJMa7
daH8QWWqUFYtle2zIyIzakeR8Vhj6k6VBLGgF6Gl/q6WY7CbP4QKyrgf0YKY
gXoab87Y5ZBjSsRXnB7NwVM/vOwibyBdHWrgSP0m7NH+qXcskd9Nm2aj7jFb
WfQrFmkxyI3lYDGYclJiK2ybmH7Ly0ucHwoXasbkeVr05xebGoRfasjBfeiP
+kxBqJUsTu2VdhmIx1fKgoXLRGrtSHLF26LCNSmv1zzRJdAhM4VX3U/pFKWn
/ZWuU6lFf9F7RpODIHdrNlDGgOwK9gnN6GDpo2niptESRItSeRVv0o3grRzd
oSLU+w8aXZStIL6EyusBc2mI462+XxRsS8bbMjT6ZYKLK/OQ2POlAg/d1ox0
dvYCUlGg1xmeR+DufETxSkZL9KiI4IibIAB4JGHlGMvOBRC5tnO3tkPszs0O
oCTU4/mazwbOw5735YtUA7WHyuo53BSLZR6kM0nKghvZfHrxUMhPwIs10dXq
D2AfichTov1WHl5xDNqXDNp66WXjN2Iy7goEs3kcfw9E5TVJnSTxfBKXhZ4D
e2qa/qL39mCR05Ucy3nJoz5RfgnqGuoweKa+DnRhq1/yjb2eMAc75AZqdeHQ
NknRSj9RbuvWGIKpMbe0mcrgP4kEHVgmNNwczkgJZd07V6Uq90QGgJO1V9nt
wPjcOsM5s06SO7kA8lf5663twNDJQ9qhin13UqkkQuGCFlDB8Tv9jlbn4bQR
gskevOePEWU7qSYRgCdEvYwBNWfU3kMmL8eJ6yInZayE8MDi311NPpO3nKTS
aDPwdDEq4d7he4Azod+AWFAJnX/ZRXt/syD3Bqxkxu89cVxKg97IEE6DYRCF
cVdmrDRWLQdWwTNYgsK7VsH7SEX4pm8jgBVLOTl31H74aLqjqKYe0uaf2SZZ
To9h8NCr4QIOBF4gapWLrnVxXowu+OCwPjwA6QUFFjJpwJKCMiDOF1+cY6L1
8b43rgHIK2QJ9AeBOU4wjgY+wg3xG3N+DBUq19q9F2QyEAiuZdKOsMH650rR
iK6WEbiUIAUBE5Zh1CvqRAVRefK8VP0Lb2FttoGoZZNPTasYRLBHWFSjJJ0F
x/0A8iFbpwEHjdC1HWbh3AL+w66whrs5YRzppn66vMwdcr9BaH+NOh+044MQ
+56mIIpvjgTg9+MV6vdA5r/RAMYFDEdjxB35IAP9JvL7ttD+7Ml5oyErwtpy
GaTswHxIW7oDGF8qhFvVqzqh5LF5iOET/K+Lk53SIEXs6JbMGm/IoIYxRnjH
7Qs15RJ/Uc00kfgp+ol49uvVbrSuDpJtfB5zTYG2CdXYLop1Cs7kGlBVHo0W
GwI2R9YYvwv2JgunT06QjbnG5fdpIjBLuBs/v8+p9Qfzfx/kB/lkZoQNCS2a
JDL8dI68boXJRqnRiwJCsDPAperj128zUT2yu0yPDdV5ZIe+8jlSoYVywNUb
PF85xPcX4cmQTqZiCiiX1ULda/OCRmo/bwT5G5QTe6umQivO0BF9zp0uQZQk
Bbv72SmQLVFkVNeQBcVIG/wQ/w2KrqVM2RyhdoC7zjQy9s1juuzzUGzATxEP
hRr4lxlSqBQ4qBYpgQEYZIj8qapV4mwbUN40DyZsUm5WCEp5R8dfaopHd92H
iZmBS3KhziB1JyFjST+eQ/o8Y9l8sCzC0b0nMny3+T5TbEtWdvZ/S2/fJ5TJ
4iZJKGINIV5HjV0e0veCqkeuD7LkeVeYIoAgC+fIjVNrhq4m9yWCC8keRZ6g
Ta/S8IcESUWrF2wg1HlHvL79jFbBtvmmkVdEkuj6pqgyKYHD1kkehy0AeORh
Yvdy7dM0hrqlOD6dQcDpi+T/bFwISEJGWvi024MojrA2Mkbtt016hUoyElZ6
F0BBVCkJBJzSLD4ZuzS8A8CdTpJdxl4ZS2j7ydL26lUXs8hGDgz3JObmqYsR
n3nfFXzz13mJd+xyN1IIRPIL6KjvMeTsPPZqj9m8auFqYY5HRMIxOZxsFxpc
TxMGmL1lHSp7nU9/IHeT0Qc6QokwjQtf+FchQVgjmH+xVjL9/8DzpG9KqBhO
oxSn4Mf0ewWLc6hHDTH28cJUvCxJmcUoedwyzVP7e6Y62Uu3LvDplPOpmSJP
C/uM7t5UAbX+OHzoXG2W1oUFponhGXhD6CrPwRYMESJDIzoYTQYaKjnOIG3V
DB5O4Bx9Uyr/8hU/dsnoNMSlvbb+p/a0SwW+v41khCVvGI3xgOchgrBdAIZM
/AB8UDGWo5yndwcHJ1ZLuQPXSN8WaDtc44W60UqW4IFhr9ZDofdSnlnH0CBM
NenMzONSTUJkN3bC1ktaT/nWzIvytaJS6QMSBVCqEob4mMzknAw6wgrXXofW
bHu4qffyRiqeVzG/ncIekTKwF6rzVU2HrnKeM0cPPHps3KXFLQW6nmoUD582
9hDfLb8UBHkdAJMCkXaeOsexqhrjrLuBpj34YVzAtb/jOmLvU/IRMLIWTX/O
VXnLHs81HcsuPeOFlr1MV+3z5a+gqz5qojydkKF8M3yvPYtKBUgqgsFjgNhc
0rQ5Wc7MDJEW5ZsBTlRFDm2jCndewL8V1fi7gFHcHEcnoGV/AooIpG9GveLj
/OMKEEcCJHujOmRCHXtuUpWfwI/eoevtyCCVzsV/a55yCVOB3Pwh1HL4EyFl
kS5J5sTQn/5u2FMYOjw6VUxlY0+kxkvzLD6d3lwHQiqeJE3cR/p2Fw3IW5Jo
2ORp8vSehX7n2hgqqGSYkgeiw9v6uWd28DD5MH1F70Er9VKxj6Pwhlxt+iv6
ZlPVzQOmD4kTTv8xxtNE/xA5vQPIdS1Pqco1q51gclZ4Qra+Up/bvZE4kCa/
SLSoxJz9EWMZF5B7n3IVApMo6novGlcy6sUs8w5LkfxCrJ1b/m9X4vaV35JE
7QZiIWajGbqZaZOd9WH1qGwszVuBm7YATu1YJeI2Iky6ooIiCx2iWfvX8wTD
d1i5OrJPrewG1Xq/D7noAoQRnyuRhu9YRPuCTYbJ/dbL1HSczXjFXOoJjQBP
S5hvSyQ1CvIssTMdzkbopIu2+ivkEFZqyl+lH2vf+J/3Q/Ugg6wjRzFVCcfY
xVnYKk5xD8Phy4Xa56SrcoZT2IsKoa0pUWWPkUr/kR7lZRMoj6USHFVQ84Zt
D61lAPrxrw2NF09eb9rj3U4LY/CVzkAEVag1QLohC5WY4ByWNkIaohI1pGrE
YBMdLRgKNYID+5LwrtQ7VRp/SBVcD/PmXEJwVRiz9EgA2rsQ8DN9I3xBsVMz
No1//nw6IbCcjrf8dLYR9qHcBI1tVFKJkEu6DE9kfz9iI7x7X+bO/BhfCQMz
rP0rgEnm8gIAOuA9kh3KuR//quE33XlPj8DlHcXdDGzxjFvv+tB5/e0VzYPm
s6F7BpTJRSsZlW/DWFt7RKOyQ/iSfkytqC+0v6C+i3uVpKzaafJphqCMHW+x
yHeF60paoTi/Dd0e5Xit3veXXShgBZHuMqDKpSZ8oAMc4lRblEKccu0GGVNy
HXj8fiBSih3VEXfj1fMH2dnXY/1npMDY9Dnjx23gEgJA91dUcGen2cIndeUV
0rGjNTvQSd4U/cBAnzWoQXUp/GeMeawIzKSTVM/Zo0K4yRlfaCVHzlXqDZp0
iUGgMl5JzkMtrmJ3IDXxLp65PimiEcYXgUydEZhll15yam4uP4q+U37oJTXG
1MKnCX3Iu7+Z/lCNFJ+V5enQ3d3/szbfXdLQ6aSlTU+EU0/eDOvn572UHoqN
qZrGZZxhVowC6k8AlY2RAlNOndvJLY44D4gf/EEZbmGuEXaKlsiW+t0JNStb
XQ0ct3f35yUhJ30ngUmUVRhXE5Ty4EvW61ACEKZ+d06NVBFuJBUln1MeJKO5
NqtWOeOlUCHucWbp4F5VMa4tc49BH4BZ+Btwj+p458+65KLrErtvmFBlIZ7p
opgPYV0Blu8ZBdOapsYAaQHWWc/PjFspVUMhPmc14/g1iRABQtaefwmEJ7r9
l/kCgyyQgvUTIgyTjPR5naFIiLFC+bXSeqhuOQsHcR4bqPmxbTLYWUjrFpOR
Reg/MmRa80ONk92wMz6HkvlWISibtWMtHSVytukakHnyAOsKPj5i1zwf1M2Q
1GUKFkR+dSJ5HN6ZyflHy2xDvTXTe7dduUXneCVWWau51P799Xh/koPcerjM
NAVn875BrkoY+WU2XPh3K5n9V8oCZd8KLw+YW1USfy95aotp3UrZHSCy0+Bf
hnZk4fUopyQfJQtFQ3lDs53pTzKHodfU+WPBd8ZQYsDAgfIh7SrMUX+ygWDY
4y6GlI7aIywmse0Qy6KahfK88b+RSFOh627HiNKfI9UoVs34B1//zag78cQr
uvpTWntEDWZeBy4kIDsTGmi7Zp49nGro3WuX0vPVDovpbbuxQRnT3f3aOd4k
98SNzy7dXhSk+pg/ex+9ldumnkL7xNh0IyM7JQ5bRAg1KZc8OgrrqD+ZIpp6
p/JIfg+C6iI/heLhV9o549p1y8YEl7dE8ZlOtNQxkjCDArTVa2HyOwWQ7edx
ebaQq7g3wJMOeL3Yqp6kMhaKUPt/imwqLmIQSu+e+t1bVf0Jx3Oo/BAwDsqz
y6/CLNtbtJLeQJn03HbHYNtoduAOT5l1NLZ3vnSR+ZSBsVL5UiHo2q3mJOOb
D543RffnFfBLVwM+iRyHvt4iUAJFaR+ErAn1ei4S+TV0ElQDw1R1TReLzo9m
yokJjSKdi26RVaDzBK2//CC2Kzw+jtI4RYRgjdf7EY+gff7PzLMZGBWfouRE
/tm0JilX5DMB8WR1aR6n6O/tN4OQT3DpnGS0K5SVCs6lF2TlCdU7TMbEu9fp
PvYtUV+7XWxdggbjH3oQ7kunELG2OcQzEupnn3ilGbXwhViIPLIhL+CwQ+Ap
Finz/9YwH/goiIdt/c1PgRC1xOXqSLGBcBSvq2IiMZN5cSXlolyNGW3/y6HB
LFo6CNOIpFD/5YkOQZBay1Cri08FMSX2BwsTWs1cHMJxV1OcIgIr5RzD876N
W+bYNB22uR+W6JCR3Ka6KXx4LKXwSa8QkEuNLF0DPlX3Hn3SuvoI5UtGr0JC
hf7QM9vKmZnlJjoexqoFjq1ifkEC324PwvFspbpPBgFnZcesQsP/KAj7aNfe
UEOI55g9AghEwXZfAQRQ426mJ6kydG8Bqh6BP40G5xlu8dV2P6GutDYyn9tV
K87x2O26m0WRhc+phviYi9Aq1i+OrTmkiAJKh6oyOCnXI1f1lyySEsIRZysj
EswD+0x/mW8b7CIi4CCws5ZApdpVHUXmb48uATfWANSkCdqrvoc2uf8hK3hP
ZNW0FUxv9ppLpzhSBCmUaOL83ExSN7kLC1Crq2/FGCwGch7niAWfcgvkuC9c
daJLYluHhG9ctEe9i7KxLheqrvgy5ktYYlAoj7l8PNT3ObkhkdIzZFPYfmtK
VyJdp5Uk/n5wPYfTSOOv6SGidAcTWbtRxtQ0JufgWxIzqH1pLyX4V3pBj1Du
/2/3Y3ODhtLZTZeernW7YMSwgKscfsbQQfXaSnfWGOgreUsMigLK7orAoR8f
DQ2VYpvIWIBaBbZYlYCjKWqh6K92RZ10sbZ4bUlp7AE5PGZI+7dB8Mjgm7Z3
zRfZqSwiyg9T1a8rAWzUoqirCWccQ6SrYECfXoHKhJ6XhaxWf0ezIlHYrdI9
jj6TT3mqIKKD8VAnZRsZLSsWk6vCP5XgXsB1PBm/nbY3wr1vri+ba2mUrB/Q
zui1NMmOnP6J2aJyvLvXpnz7q0Fd5Zz7NPaWW2LHCwHFXdmIlA78CkvZMxrb
NSZaeIrLbKXWVHWUlt2/GPcuf3msx7655z3Q+JS7ItPmRzYnn3fF2ABsZgjd
vdMdq7GqLmbZpBPaYPcIp3BBZ5+ZvxvDOv4o/FUh6c5acTas1AheriTBqyGV
1amG2BfTXwxSF2B3/E18TJp3ZlpPooyGvXB5uSYul910mHuo57koE8ubuorZ
TW6KX3fbna31T5h7N7L3j8swiz07tIpVct/jwfl+kS3C3edUZDAtsQoErTo8
chUHyUEIDSjv6C77eke3os0Bq1/ejh5KW2Lg6fDAYs9Ov5uA5HKjffmOWfSG
8h5+Ym7hOIzmO8ivFjbphRQ9klOMfuBZoscBi90CxZiq20ykk9/yXdkCJmfi
UuMp0G7iwZc9S9E6RqYDMQ40ZYGYujMmKC/WnjgIPC3Wo/XLyD76O0pEKYj6
CzpYXDee6nGzECCOwwosG2H1Rqm5Y11mvg4+N1gv1Qszd3+Jt8Y7GGbtdn9M
1Oy7IXDPNdu42WaEQ8HcfaUYbee+VPds7Tzf8BvAx6xaUunBui2g7GmQAqRX
58fGspah796S8rqODIqOsTd0KxNR0ui8BbIMlw5H+TzhzDMyO0D9aJcz2BTc
3XbAQ7jJ/kt3lVZ3fJfJ1Qpd/aDtpUCvitZlr3GyNY1sMyeTcAfya0NjseiU
3lnmD9bm93fSyRrMknupSiugWJEJpj4ITFr1S5QMtBJ0czxHwTFYUTkwuKYd
FQg0OQHFAqPAVXRs4GgZh68/1eiHkoQF6nLWIaAdCZmgpnKxpMTJZ+hsjDeM
C9goLdKMP00+JsPtO+uPgfqZu77NEfUrkPRXz6PBE6Peiozy56jPyKFo9iVu
I6D0Uf7+8LB+Wga7ByS2pdavxndOxxtT1TU7mGVZGuUwPVuy9urD1lxkjBWr
kGpS4hYB+LjJ32osqz/cMQKAERnY7nx3LPIwIGc/fQNF4Yera5A0h9Swt+Ur
EavQl9gMtUpugr3Qst/qaAu5SCC4hl9x7UHrAQ/hfQWOXXAjHme9VuzcBHTs
BPNWQ826EviBR8NWMq6T4QvFwmIwpVj3NIkrGZcDsVFQtKWDqVHa+F1Ff5Qq
xifXlzlT+n3mlGOR9Kad+axMf62m9rklXgFMZhvCfij7DnaqmmW1jlKfg6pP
wi5ZhdLf1NJCN7RSZQIaxRAfSJZhOuGtV3QOc/q5XCFYGEwYzlwhPOE7ZH/t
0mCVokKlrypQ9XqkBTVIfghyy8RMxUrciP2hot+LlAYoWs7YO6DoU5r9DWOq
bMvCismNf5oGKJaXEFTxDBTLJb0CJqICft4HRdtqyg3kArHd6juNluA45SFO
fZk6ahQbo4jM7a3drEeLx+UyRTXrg0AG2CGdDmgP+ldjH8CkQm2oHOVYbTTx
yWU2C+ZqBRXc9hzjfD6wi1X/1uSaU4m/F3IfXIjAHDljDCGe6L9Mo974w7UW
N5wEKhNakgunyjVS3UNuedVzaIfSJ/aWDvvrByQeSowEHrO85AKmc5RKPHgY
p/wLd7kN1KPGUCr8SmoKYq7DNqwlOMg79Zt7hJ0RTXXQkJKmZSBra4ZSl4KZ
3ga4OPVJ/fmlp/EWdYEHPp9qi4AVdcX38nSRxWBIsmpYC4IG2CuFyIuhYCaq
D5tb8Cs0f+ixXo18XpkA5Q+8SNuZvSBRiacHsNAA4PUeV9Dsc3KqgHg3LSZK
vRBgp79khRqu3PPCmvMLGdPdlVC7wqIMc8TCrjQy84ORv9ewxh4AMwQxEuJl
wNgcidJ7xWR4hdDo8kSLtiTsS0XBCqbAFoMyqcUqHhed7vbQ+BU52dQx1rjv
9DaDA+AMTxJajmmiPl8wV4rYwWC9p29DVHyJZ5oIm8gwtKr8jDkJclpqY/ZK
VWTN04TDsT2EflgRfcPYisZdVpkScwsDrdLuuecraoLh9+CutFMj3jIZXKKR
25l5SPeQlCBTcG0fHxnqx37MtAlRKY4Ei4pg4RjuMVVh7sXgV01NZLjxr7up
TDsTGU5QoDNvS79z645crR9arKJB6l4HXrrQN67xmmg3pNlsv1jeFGiflI2F
lyF7o+HXh1rZ+glBIiRJDj+A2rEblaPOTd8aaYlGZxGKUxILSsllG84BND4s
21f2N1dITVBOFKTIXHGqyLovB26C7mg+9vwfH7489qdI4Yzjk/CaTzhdnfst
/VEh8eRoo36aNu56XuPK04QYQ+WhJzNL3K+yyi5mOcMag3+FwNuQfrOP9FlN
/F8ZXJHLiEuK5rV9iYQO7ZoYrplXt2Rw4VzDIx4xb8t6lQkmHVmFJ7nWDJ68
SAES8yJUfo0ZVuIJ8wgas1v5UsW0o+3d8kKBuEWsc28m2lfUcR2ScPWgoqOh
GPIWsxYk60WLACs/3aX1lpVXZ0mY/8H8Vc2ce/JnSW8nvbr491yghPybeuxI
PN0kcIrctC8Bae7K2zelwaxEJT2zuBSQ9BnyBm2q5AnCFWtSSsPWRkzcIeEr
jxzIPWaatwKS5DoYiakqKykX2D++ZufAzMGfsOZ2KSpN/NBZqJu4N1BZpp1W
DEPzWoAIje+pFKpCYNFwHXnF4uv4zhTwQtyWOiEwj/DafsHzIEgU0z4/37Sd
hViywxNvgA8JSrAStTt8pnNmAOhyB5qEyykGqMTMnnKsjuV9J+IqgiqDAxD2
6Jt76NoR2+x7GJ/GDplesKHp0d14vjhVrUKxRSh9f2BGpLcLxom/eF+hAL3m
AgbLYm0B7AsWqEe+PJDHNmgzwpGn9RzFH1cuBwzu5Mg8d9s1nAykgyny+764
6J0kw7kd5MkxeRVzVfO+HEt6zkjQBhOuz1tw4KkiEK9JAzH/Metxb/AH1Dws
ZPITjCwXaQH2w4MT5BZWc9T8yDVDH+qs3+zgSSfWXvij0xHiojJ8k0uKMxAZ
//dFu9pz4Frfykzr28WTHUg5YHcBcWQfrcoSG/N3JVgYO7K3EwpAp8SK9qiS
e8Vg8Exldwbp5w/Nay/2JWqFN7xv9VlUL3gpcy/PU7iJXPMYGMzIJQXvP8l0
YWBnETPH7pMhy+UFZAgKCmER5JTYiD+OOWsfHZOU8g5eoqp98yjqKQ09HUGc
DLvjTYIzKntFmvqts8lInc1z44yx9UAhhsfGeXWUgpPp1IgeOUkPkhjVXcCL
Xkcq8KNQW+Pdsx4xns/YD3xXfNmxog2MRjRXUEL39BbCoLkFnEl/ZqQkn6ZG
ldKZ5QpcQQrHoz3M0PwIwvZ8lcnD1dz/gTYg9OEmEMkj7OgUgjvBlW5GAJna
RcaAR+9sbqsUFBj9CSKgxUNaZ4/oSZJSvl3LMGv1o/tZ5yb63g/RQIAliUZg
AaLDTxXatD3pWVsNrNDSqpd1smvsM9pK3v4oI51f7kCZmFlc5RR+6Ah6AQ2+
BNyTqoh2526SH6iscJ/ZXUEoNevpRc1DkqWJbJxkfbvMXWDSMmxrEu0KkS7o
9BDnls+cAIhQKKfVt0ozpp0bsEpdfA17tsV6zDFtgRurNxjdu6VR94rT7JfJ
d0Pv+btBe1dnOGZs+pYsu+kXQ/OMN5i0UJlB04++Oh0C1MZ6n22CtoymJeyT
jiH6wseZvAMMQaCUtkYuQUApFX57/JLTGmcFea06dXVSiQvNA1DJJIt6S1WD
D/otkg6OnPy+yhTf6yPJKoMYlbXiCfND/uRtv/CDmX6FDNr7Vr7eRjn6VpGx
h+eP6+JY/qg7n10Z+XespYwGNPUAx+GONR+xDKgl8Fmq0eA56/+jvIFKyI7v
TvkmyhRTA4SbSBOpfoVGwORRSdkFq0UyEwenRPruC3+ClQ+9DYHDa9oylZFN
5tnPBWIypK57+4t/I1VbI2aap+Ja5kNGeJx/qEILav+LUj4EAoJv1x/rLG25
CkdQvyKtxa+dBX6U2GS55sftjSOHgFhIfb+Cuqi6pYk/cA5C7G61McRbcKo2
BtcHgbfWBQJMAZZlkvlTgyEx5gVkk3a1Hr7yqVrwdyqegcEKzgHaNbRx9NGl
+15mUU5s1FZkHIm45aS07nSV+zuVEcFOgvb4em3iOPL7R8+lwCgv/RsE/GXK
DiQxKE8Sj1ve+Dfmg80aUug4dunY4B1j7xwgkf4Ieyh8cDmsS+5/UKiLdDNw
U/da+ky7d0E//fXkaQhTQRutdgEMu3Vd6PfmDcquabpiZjZ+JMYczwgq2r96
nCTSo094B9kiWqFooqWMCOrCgPFVUUH8tsVRAa8jiHP5nJAhrsqZfasTjNkh
sjxUY3//FzuULMYf09w9qsFhlRn6bj72Ne4VDDvIWAtpQaAc/32CB+dU8lT+
r2RZsRlhokJZhxUHurqLCh+j80CaaLbNgatcmPHN1e+AY6QEuLWiBRYfVT5x
1R0fUZDjk4xIuxQwHZm32wAQBetUU1HcBONv0yIeiSMLyMTey0zRLepFduI2
Ko/fjbx19L3OKNRBEv/gT+5p7n4ljR/JzghjT+1KGd4W1o/rvafNuBv4F0wZ
kTBG+t+fQw+FEFXRyN53QAs+R/+2TIFZFyWsE8yvv1KRgQ3ZD4TZPDIeyuVb
j6zQlyQVnIEwpTv7hYmGpWEW6CE5FEz4C7lvBrL0TzaEnOMNUqlq1852WmFN
WwfpRsC8u6eiJNMLUSF3lqYqduYuqnbJxaQgh3KPAwHvH8YCd968z53Ppadz
mXqZFnMaJuxQzToAJDQzxeF0d41mc2L4SAhW8UIZAaxU1tYP0DGSheZIQK3Y
jLH5yTWlc6FwArUZV8yZWUrP+vxIQ8TtHIBg77EkQdGOYfMJrLd0jaehgmT3
B9AF0b41OSHIwHWKxa+LSkX4+exDCY5oHCmFuyeWcdV5+jTpoaf9MqL9rDal
F3MCzvomA1/dh1W4CP5mFwz1Yfo28luji+nfglIo2/X1P8/wpOJIc6h0W0BF
KLYEt8to2CpcEiGpy1wIUeaPfSRW7HcjrDmDjqf9BIr8m1UiaotOYHW2j5on
i2ZsyGN9gwla7j2F02lG0RC/M2cdWhkUkSWXPTWE7JcNx9Tap7zxOtl1PZWK
RS2QZVdQbtjzefdI9ls2wYwAIr5yAAdGWefmDp9SvQ16ClVCBOai/d2V/FS3
qs/lmLPIeFeLukfh2OU0w2tTtHnV23d/pANJLg5QuEtQ49DlR/dwe7RDI1kd
XNV1CERJRICrL0h6HCximR/C0h8liZFdsUsJe+DT5hioaLDGvu1kIpVr9Wu+
heN4xnGnbBk/bmmF8tzTMYgbX0NUp97cJHlzb6ZqHBgWQa8FV5FovCkZTrDD
elIDXe2ylLVkk4TBp+FvRG7ITyYtbSY6g96EyU40xrAhPGl6jWD9yR7jCivN
iKmLeI0F8O2ffFM0HDtul5zsD8+SXFjeZ4VRjAJzevjTQnwKPx3u3J9eV78X
KUZQ3AsrG0IDnDMdtZkl1Iy1u20/tys9nNCxlwqjn2iJt7XhLdHmV5OnErnM
c3hDDx9xmvqcP59mjT6O6+wY90BTRk9vN6b2zu53tHLsus1ED1+TTHXa/ntP
dzo6pvoZIrCAH5Rnab0ACNJUIqxGNMUlxEaQImf2YM77OGu03QlkNsbGNvRY
WsIT+hf5LYgrpHZJsX3nP33fZbmfr4b419ag/hbm3MOabFflzIuQW7zgRcj/
8gk64EcfmmdnmraauNmNMjtTwG8Vp8XdGjovNIDgNIsMtQzJ8drKGBxmFtl2
PhS+S1TAWp1uhAIeomcYE6XGWzJy/IGYQlLblBmUuXCf2RHbCUu2grLBFbdi
QvHWKf3k22XHkMg8Ot34EBUYtEK21trieEhpBaGFb1p4e/T1p6YmcCHPfC9G
G2vOPh+2sJupekPFFmTTAORCBiB5tg5z+3kVjgygsFQkVMtAuixSnqkcRPZV
Jv97kgEsenJ+7C7lKnN+ongr3waH8TerwwDTU9Ku67mfeg9HIu6/yH7LmLuS
HF5cPszCoNUD289PdlBksf78NH+XbHEbbajDBOuMV739Qp3nLRhGOQ4YSuvX
tMiLL+BCNhL4RGRK9tr2/ZNN3RPNIcZEQMnEloy+7rJDb078TRJ+yHiWHCEy
3mybMgZdkR1vMF6n84gH77ZeraVHRmZpo8QexVEhM6KXWg/cfFN+9LIyMV6o
U9ts3nemYmWsFT0p0SssmrDwdtMOgBH70buQFVLasxI3YF8CDDTng/hwD41w
J1nBZr+zfJCGXvL35U0o2SOIEGTh/kTUwQwp5WMVnJNvNX3U5zmeVUw/GH65
Q9yvZWeIuGVRJy8LdbySkJ+A1Nuq2NW5zSvSPR81OKKCx2uKilWSxc6lXqf2
usZmiFxknrKRPsf3fVXZQUewBJEbIOsAg4z0ABbziMKa50y0f6pwh7Z2lDFz
QTJDUV7YZ/0gqS2123FfrcCs+48Jw9PxV6an8ZzJpCyHUEvwOM9Un4o0pqIn
dEHOxtYY3eTok48F4ONTEW7NCBIiXpNTb2cbomjGwOIhSA+2Ayp2p+KylJa8
KK5hV9m4iW7JKY/r/jNzLdljx1bfeAsLbJ+CgCvpRCQEKwkWfzgp3ipvXC4q
dz78+T/NkpvkDHN+e/JR4ZwaPvTgIy3pER9pRIK/0bDhdCF/VgF+pMGVwUhK
yrYWrcBuZPF6HQB9V8uccFG4YwvU+Eea5Zujbs5DxAAfI1DSwpSgH+lEfuVD
wjgaZeOgOd165wsMeiCJNLKWHlU1tTPo0OGbOl1I3jShC52GD6TyHfdtU0NF
zHrQOBmFtmdOf+36Jjh4emLAnRfsjaXiM/AVQZN3BZx7ZpAWcmjB1n95ILVu
KAlldjCOdLJD8fsqBfQXwr4OPv0XW7uXiuAEtH6pZkpCYsKpfOiltqPSZvFE
3rihdyKuNPvgQXGxP7uLXTabcpYxMbSFcDpJwtRgsFFbhf1yQfRcYWoSlolf
SN8kh6haeqO1vdcD+kCtRKrNGafcSwlQ7srPRdLntHsR8jaCJd66V2KAq8We
Ul5VRSv5becbiON/UQ330a4JaOeI/NifVCtmv+G12MO/xeoqwBEQm1e6OCUg
fOIWNYddxB8ReF0TAfVqIkUjCHHtouUE8lfk4XGSsIY+YbZ1GQSo9oNDwFHb
/RTfxlJsAW0bUErhDpQH5xYltCqOtfazKWw1hR8KGfsNYOGWuJgb3+Kgit2L
I54pXr+wHme5VdG/ljpLkfeIAiTrnEoFbei+z/Y4olrn/A/c1ERWcKy+Szq1
m72byozF4FyWWIaXppGy4gZvf+iARznFN7SDqc0UxUs/3ucLmUCJ90qUn+zY
8K7x/YgPDmjtGxiDNEZY778ziAzpnMjVf1LBrPKFg/9Yvk12P5vQ//DvrYLz
/isdjO+JhkXOsth3yLZgs8jJcSqXLLWAwU3aQ35VqFG1oydF6G4mG64Gfqdk
Qma4AjS+lacWK9RyJAjLnWWDE6wptXCzH/fJaAphvIvPPS85JINBTGoHrQLy
Idxgb8qYNGko9oZQvKg1siDdCizGdoNslUspvYlS6WuLLu+rvxZTXEi9TfPA
GRXK3CczlIHvrUhUdPoSXLC66Zcf1d1/l4j7bcPHHIBucIizpVVAqSc3GyUc
ZoZA2AJ865c5Jsp1WrDe5nhdLyCBhT+aIx0jyQJjFOMCuy6sdzcAG4vBIg6i
QMtJaSkj1kLgBjJ4UTBOAth7fXGKmsvCkQ8jUJAN8qHdDwryYT/3ZJmkyjK9
rP7MUUUT9FFMjMIb+uRO1EPr3PwUE3x7WAzCeS75J19WzUEh36vBhIeyfV/Y
Zbn+sCs8xFolb8p+qPx4K/mmzdL94RQjwGRIoCGmET7+7PbePxGxcadNVL74
0bOHYM+02SIkPb0b1fw/e1cyCYYF8pk8KqaUqUMBIxW6g1MCf3ua6ey7Mk60
AQ/3O1Nmg6l3vkRhgqOZpl3v8awdbKMHwLCVUTpJRmKasqKvvcxwC8XRuXwX
mXg64F6rAQW+/Ez6BuXt15enzM7rgP8sOkp10wceVrWS+gepHfECVTH2HS4G
5rZbWB6tGp7JLIf6RaHDgzHQeoqP0egnZU3KQduVu3M5GSzLqsW0IpqxA1Bg
1FcTbLDTcDxyvKzuxJTLHaMQkSk+MIB13qjjgQtkeuiJUBToDFebOuGHo0QC
sKQFhFa0FYDJufvHkQ0AR/TbshRDKr9DYLgBL3Z+3Pxl9bZeYTuC0PXZOV1a
131qEEUBE7jCkIFUdIwsJiHO8QLAPr3H5ph4GjPe7Ad5GD9JFUHMESJOZvvr
LoEtkUbkQ8BdVI/Px0deT5d26kQmxRjUpmHvTCrBFh+tNzK3zxjtfc7Tkys1
GiJsAWwOOdnT6dAQSRlMZGsTK9rZf4E0qiS9YnLX0mdDez67iqu8hrkbkWYV
kc/Tt04mtwui6CmZKn4f2ZjLwJQ4KJUcStQxAwaPCir06DeYqn4CtTBaerfM
H42o1uVkqbg0JCCthbjJUievuLEmvMq6zJWTdBnEszlTFFhUPYZ+Sttc56A5
UJUj2s13A9x+mmyCA9YHN8Fp86EAuwiS6iXb3Rl32jDZfcq2KZXwGBMrMHz0
agMWfi5Bz4LaVSBJF8rxtsZAR5IJJ23DjxdyiOpnNUnItDGpVhec4CyyQ60d
Mi7J0dpRDwJY7TbnL7fj7xrwf90SwYEDPdi1/1AN4n+0B7N0UUVCix257zhL
wdov4xaLX7KLqPX4V8lzyU6IXqAjfwnCuYUfzFkveLrZV2L2hQWz6acxxH5C
EwkAmpQsJsdUrbJMc/jgNJsora8tQgoHLr8wSfp/n114993/bZnyP9WbrIqF
Q1Hf21fXKt945FtFGVgxqH5yXUO8XfzaCa7gdfCSbVw5liwU2+Kf0KainTEl
QeqgUW16nj6ztsrKnrtRTxPo8V582bbLumYt2ZEEGKWJ7xPM+B7FUoqHv9eY
3kSAvs+lmfnsfFG73CoTuzqJtJEsEoawlSvI/hKJXhrd5lMv2lGAOn94wpFc
AfYd94kxFgAWeRNxwdGEu1U2thKQavSyIzBxC3PCG2XvCthUWN/JrMktgEY3
bUJug02kokUHIO4b7X82NI3M3QEdhK1nmxAligHv7PZHEyDres8Fhv2UfmAU
iM/WCaVtEuvRWHXRkPGb1L3/rlAwq6LYlturLaVE+CK55F8hCSjDCuKyMnkA
noy7SEwTcu+2iKoMYZl1g60tAE5N6z9z9j6+d20wVuFPXDws1KW61pmKD/Pr
lZF3ZSgwOFLOj0SI2+qKyv9tMD3ynItBSLloObvvstdw8O4UF1rKI+HI6aQ9
dcBefsyYH/r7VCsxLw2ngNUQUsEgP27CX1pF/55glM05YYV9JPyTR2tGqzVM
0GW+7EwxZBvig6cuLiy84Xtf0+yaaG8sO02R72MOdF+2wV/C/c72J0Klo3qZ
6Kyu4O8sAo55oq5p5xPVDHNs4Nwc0vsggPtKTRCELp6OEh8JoZmN2aR/fvTn
UZeLkA/muBU+YOQlS7Xf/KMMJqGO5DrKkBGBDEMc9fEitTnlLTH4iK/AagwE
U8GbgHSZx6HE2+MEexfGyZm6z24zRms3j+qOJOTgXfdrPio613t+yJe+XcmG
xJVrsgWChgQfx00EdS5/ImD3L50x+0MBbWM5nzGphZ6JtXJUfm2Mxqy/UljU
4fkv8EJShWr3WTeWiWqvQ2tPPY8p+9GWbh7f5Z4zDdwCPH3lqa0hikUjTAzN
hpSYs0e+QOTzaIjPk9OAjYOFVr3b+Rneyw5jzgJNkXQB+ZzvMy+RO2afgcbI
zMLGttnFPnhuCsnxNuof0Kh6eYFhRU8VRz2Fk8rfMTLRwFvDsB3JveMdpUkW
zdmEiwWtlzGTzx+93F1xX0Zc4ZeEfuoA44mFyJpK2iOG80jL+uvRC8EEhyF1
+idYftRHmlfVxf6BZYp2kvN58D3uHYfXB4ABkYvbneIN4cnwzXXdCcFNM2Km
5v9j9Utkf2HrrpTgMZRQSMLBzJwW0iMMjPujWlcVccsIq1LpYAOFwP2+q4jW
LRh5lSzYrRfOyberdzzKWJ+cDnvf/OdDXTkIJAwCBqGC3OUasxrY0y3ehAdH
Te2TE/YOTU7KnEBzuFwqf/o1w9tdjvcK+c1wfqvYxZky7xCgSmxhctnzhWaM
IkWKSfZlwODIhCkXBhUuCAA2DfUuoOoTmN3XRg0rIu+65R1WKvD8yDAHNE9h
1QhP5GPUqiMqNq/bcl8hEUbyzCDTkYiBc3Hnj2nQ6fGafzhDP/iM1qeFaBFI
TEJ9o/nwyzFBRCz/dkDJCL19KL61FjZnRqUoKelKFzujdEcSM301imOGQo6I
GZ/lSfw/3PCI99j0hAUFwp/C1GBu0hoM8sVfGlb+TiyBSaQEjWh0k44WDEgH
fFoxdnNTBMYBDY/71Qp7pRucTrXQPmAiUQdo9pu1zS7hFbTmT1Ho5zdy2Ef7
SeclHlPpbIXLnhSwLNIvLS73cl8RNJLWWpa+3U9OIh44+8kgBC9SMCHKBmKK
DLN0A75WamsOCtHpo60SqhZdbZFkPCOUuOPzEF2zxh5j22fLT0ePcKtkwFsi
VAntpzI7s5bjOBHf9fmwKRSvIZ7JcxXVLOcBXbJ2PnLTill+Ot1scJjhGIHW
n+1xiZ8NHMFXS4IXK5ER+7eomL/5pUHvp4XET7O35Lu9db7m9nTiZhGL+ebU
ApwnqsC+1JiwGYCjrsQS+Gg2kdIe/SkjHam9nocv7geVGpWLtiEhcfS0cOd+
yPAM2bEZZSB9UVTkpERWSWFR5tzbM/5SQaF1h2LjxsmJFmufOyUam/PT/mio
EP5OIiCIF69fAaeUuN7c9x1Spm3QhKk7oC64eojMTZfuzr6j97xKi5XqpC3n
5GFnS9p/T+YXJxM2Idbk82KEyXBKyb23OETPG262L9ccd0HdT1o397DfpGOn
2EefVSVcLNAlZp2XQD90gk9POwJydze/YCvlokPb1kaJusW69ipJa7ijagPa
ewdRRe+ni1WNUFejE8io2ER6blErjz24/CUA+/lCGNAU413ZHJ9yKL0W8jJl
yPSZoV908tTqzB36NlfmsK1j7wmS9xIzj1d10+Tb99r6fSTd5ZPcHuf/SWdK
2gHvjY+YKzES2WhmQ93CMdOzRoa7/0gD9k44ASoiqO59TfJtsej5F1l7djGy
WObzP45aMam6UI9UbE8x3H05cRSVR2wS/zo7kuIu4Aqao76LBL0ScXH7qsTv
AT03tv1NVb9BjRjQrnbc6F1YSqQSv7pyqDql544LKpx/ozziDnTqexiMmP2F
97ry7VDXiRs+Ow4IUCqaV4CkDNuk3r6JJotMUwXNLc0/iTojL0VgcAG4vNlb
dptK04k1ibvrnOAj1fEIuMrYi4XntK6ldeZSKEmIuHLyXjJ4YRRjdaFyLjhI
YcSgnWMXJ3NlVKnirY8T9HvKeGJbfwSenSPgPPFGgZCu+drWohsNqFwdSWWR
Yos/5GAD+Ys6dAbFl1Iq24ya/XxvUAkKtg0W6sqi5TnfRWE2AarnkKT2RNdw
puyg7aCDnkJz1TOBc+3fE3twTjuxSLlLToKW12HwlCpKNXPNBQL38cVwImXk
om4eVnp1HwIFlCqwmT1/IwW3l9hoahi5eXPYfnFJRgcuZqn9Xls/wGhsAav0
NqbliUvzwZtdzwz/t5kr8a12YxPM3QgN/g5f+F2VJPa++9vgDgwBiso9JybB
QuDbJDQL0SDToWvzXlBF9ceh7EWZXsJTlIr7cZnGPgRrg0vQSm5wgDZx73yX
xIBtzTu02CPGT2k63NOjPdlChvxCylcrt1MF9L0WeZDaOm95i7ZuBwYqVVux
PlyNqupjNco98vFH0jrL+EXFSfxqNtD8z9aJkDQJ1aCpmiR1SOJxIYKLszSO
iF3Pr0NDA8XPdKAGkjVBKH8zlrEv9A228HU1HjmtGadJIq2368oZO7pNUIqz
htQ4x+6NzXUAHKaFobJ6Tml4kSeBi6QgN+Z6+bFewqlDJ6WScyujBVsSCi4Y
minNjor47aMaYCRpwmPsF+4aiE4OcNXgfoczpQ4kDQwpGG5u3HdLOpnSYt1U
SLqm3XtYp2Ejr4YUp1+5cUnGrDBwkeVRl9+BPQ4tNtEN+hAY/Wv30T/wp/22
NY/h3WWS7zIPkMTuOq5/kw/6zeb9fxryWsWkNm2jF7MLk9z3zpZ9qh5qbhJa
QC7xwM4Yq/C/SVLW3y3PykWuq2rwiaSSVaDOe4/IqmynbExHraIG1lJrVIZI
+rEl/9Mj4cgBMb5XdZ8MrwkJMmW6bn0oy6gVU2e0lh60rnYevnVJDsubpfml
PeD85zWczG4Kaxi2ytGEps6yRvMBMPNzB0PbPI1qW9JlGM2IK9CbIVL1VwJb
rlUUKv04jhYCmtEVhs3+W2mQA7ouA/EORXIKGloc/H/f3YQpdx4NTN0MS2DW
4wk0Le5a1wgG1LHvKwGP1w9z7GAwhKkabPpAsxQWSXzdbuLbltLm+1RHkzl+
GL6We+JVbx7lC+v5UAwG8TS01vNSYxyS0LpALdSXGAia9wS6O+2H5vD8/yAV
cBMfMhWUqZ1OJl4+Z6oyhbfqZM254fQ+OBpR/6/7eKUEI52zz68dBznkVGpF
tXA9cgZ2YyC3KZlQ5CxkxFMOd6kvhpEGhtJ3BSrwcf+rACs59ZfuTLgj+2nO
QJhsrb5SM6h4k6La+2k6GgFcOnIjq/U8yXkq8aGlbS3fbgHn+o49yVTFz42G
rjzWouRzSNMY/20OMaILzRf8rziqSaeyz8SRbfLvFm2qmixsZ3MwBEMR+Mk3
gRqJwDsSbpmkOcAb2eBQh3faTkiID1WXRE3L2jUaHieFObRpNVaXrSk/WKyD
8AvEMYQhQS52imedc9iQQoGFZlll93pQJ2ynHg7AvCJjhYxIT/EfDiii3qdp
gE3Xp4ojg8J8Ignt0CkIUKgVLEJfuiugrZ/3N8PfwPLmJgcg4qeTy6Z7e82b
OdWsYSUJ9HcD6yO6u6xZ+0TM3GPOXOcSchGb1+IrN2Tpqr1NPKT2TKMBe6nH
koRW9CL+xSt0W9xA2NxzDqkPrqklCcHi6LFKnKKNvSXh/wkDsVpzrjYFBvtQ
7GPYB2hNcJK9A/my1TKumiSl7d3aaLGuyj4Ht8yD9j1I13N8fgiFNOzMWkhx
qtluV53ztOj18lZrLhD2H3hii9EgzaRoBDUlhXJB4vfe2AoDs01UofXZPesu
kMWikD2uIQ5cFTa9xILywtrt+SIJbEyW2WK64Icrp8f+eFmMfSGBGk20/h0b
ldKgJyIQ7h/cwHT9QOleeOUViG2hNsIp3BhDS8pCXohXLIvyUkBTBcPlY6ts
KfKaqpDuW+FtrfGXbUDnt1+yxpj6wp0Z/PC9WHRdn54wPi/DdxZVZFzdeuNb
losrLaU+PEQRexXrX6rrs3fBvcU5NAiS+8nDgsraS2QwLQFtoTwW0Sd+ovL7
46KgTM/YkQGZ5ItwCw75ky42Z+uFC00LXSxGYzQtzqtcxxwHbi0WEtU5efNC
jGcCqWU4KGxw7hYf+BW1whfMHJklIL5jBe/PSIJX6PMOsgrhyLyZrkKpMwCC
UdQYALVuof35QOyl93tDouCWFy3IrcVRvCaZ4XtjMVmn6KRfYqcplADlY/pi
N5o/L/akdFzOn3UDVtjzRHFlMGkNg0Bx/1G5l5WegZP6/srg03Vyq0eMmnsU
8OuLuGTu1duKZidZpC1yyrypjFT2ByBrqkT8ZxTesJgDKlFPfoMEY33zxVUf
V272xo8uGgJmRPUrSVjqIdsqwXW+MgxvU0HJwLmaU32bhnsZILzlH8v0MWQf
w0ERz0H0QEG5zsN8oDqCVPxouqKP+Kymi2Fz+E1umFi+TL1xGaWidJiDSZWN
uENtFL2IDnG/CXAtTjQGmDzP/6hif+OF9+MMHfcEeukcsFJZKW80H7odmADe
AQpOe7nUuHerSArUvPRTc1ACQACQfbtRQdcQ4VPae32h0q9hwQ977SsKg7JI
Pj+tm4XXapsczWgRRNl+GaidJajqMhD02n4yf7I2SAG981Xa+6iGOMvDJ4Fr
K9f2/pLakHFaoVMcREju9/LbMgPkD08v8JfCZ1NsWmwe9FxCUJkSaGyREdoc
wUO7xMMsErTDHoJL9lxjiKHgIjeWsK5eKoNGscGPe6TdNAopuid35SGVOn2q
lwcK3M6e0G2ElAlTVmSxJpIvRFq1fx+xNPqD0DmWdXmXV01i6LcxtcjvVb2s
quv478y10dx9I2t8iWB7VN+nppKAbzXeSMAqJKVrRvYzQRvVIZHU051iV51v
VIwOcPCikxDfXSSFgXl7fGEA+bZBaAjnWrQC8p20UjeBe7EYLanZyK2kYfTT
t25hNGFfEV4cejhwCwm4UQVS2IuD9uVvDBy+jBDsJzFn09rnPrCBNmk6jUr7
3eXyCaC4cxr2YshEMyLUH41satqbXLeGFPUSWe6MUaBkP80ahNmON1XP5522
GNaq73AtzNDXnJR6uT1gk8z/zqSzN76VVFsNVihAmPcTfBe7SNpOltIbj/s9
AloLSS02bbm8CsS+OQGH/9mpqJBD7FJtXZq1hJEPqPG3B2fWxzRD+aGKccYo
xLr+xgWrQ9q202S8TXvmMTAnRBhr0+pfBoN3equdWVFuU0DkVsrcsva4upBh
RILH5UBPt1GAQA1WyAQ5TTGtV4n/NKOzszn39mAgWViBQ5oJWJ6VVuVAFhHb
rxFH/Cx5wSdlJpwNjoGD4SAev2GCgoUZO3w/mEPZ/zNKYkNxCbgfk++nVK91
vxf45N2h9P/ezRShO1DDopFc/QuT1Kzd/NkHLfAnZdiiEyBB4NsUcKj61Fi3
uvOphmJxo1BIt/Gi/XUDWADhtdXteSVCHlfE/8QTTQTpz5yLcv3qRNRSOgcB
M2Ezf2H/oA3Cw8+BkiaYkkwAej8EqU8/3MEzxSzWN5FCjDsfaORKwfO1Bo1a
gXoTuyGAA1H1tNNbZoInI0EhJAO7JG85iA1j/Mr38S8I5NMCsD2H5IhMhvFe
XkBw+3LZHqQVEMm6SrJHS5PNBbajdZvYgkT/E21TmzYRPpNshoRkkTZ6NGls
EJPZ13CDXaJEDEhxlHBdYuuXteFH/0A3CSMMSJ5NrnAMMOHYAiJYw3vbzm8h
F6J6Z5ixdmf+bkWuQRmJScV7qo/+a+30mPxpwAbJ+ww7FX35Yaimarv0jccs
8beN1nHhhBIqa3aFSVozVF5WACohFuWxAv/9VsyRqDDTI35xB/Suim/phMrL
+7UBBslqegWjbLquRulOJEnvq8gUGSqNqB7MVK73isrm43ac0GqvGsmNWy8j
tQkcYibjVQj5vgCXOqxY55O6LqF6uzBT4umGkVLMU2ViJbGN1JC8Q/7WtAyf
ad/PYHV8Lv9AjLlygopAENXU+ysYD5bffPE1NgDgamHcbtIZdIKLaWcBK5mW
6BeoBaGQlAOvyBMnxVt1wIr//p/avpt/69/lmiuTH0ItGfCCO4/MlVuThde2
xkk4LAHbAUg0y4THuKapimDOEUjuu+nDcXy+hQsmxIpORgTx8pIMdtuJpJba
Eqc/WLuW7SHvfLBVgN4dR5olLevZ9uLvoxd7vwDTgb8/Z2exTD38Sq1cxF6X
LhXBxJj3xjnaznGxbWvn+LoQUCu+QTWyx0GKXYr3wGeZk5baeqEslt6gqQs+
/5bLY/J704/CjA1ix0Uz5vmuGoQQREi2efFLc9Xh4Lvtyef+rXEdqq4msAjy
pvk7v2wz5WkAnSB3JwSI0Oo3/odCf/DX+LVe/lt5OsA4xa1VUbIU54ImDPct
+vZRFuyZQ3AudLkaZWL4jjTtWZmnbOIm0Hj9blQcz3ByE5uoAWUC3JjRUFI/
YbttEhkK1c95eHSSJhDVrSi4xyxzlPiH7/oGnELIX5ucMOwxvtDGq4p5gwZd
uXLDtA7dDvn4uBM4G4t1fWfyKWyWlZA0vXi4ZjEqybXSGWfTdGZG0VCyinDQ
Ad4fh92/pVzzXrI9hVkCf2PWzKkQrdGckzUY7+RpbZvhfEFuLOw59yoajXCP
acvt0N3BZkaDxRuIPX1FZ0i0h1E+FtwLrXH3okUvU+9AKrJQxLKTspr19SP1
plV+E9HJhR6crHSWh5tWwhOSlbKl/WV4R6hOHPv9rSFsWWM1uTodt5RAt/Re
Uo+aG8rla2jTk+hxQYJhwKDjgIFk57O2si1d1Cjx+sL+EuO2pD6v5AecOOeG
AW8jeAxRZsTeccO1cNePrsl0446iHsfCLzfYZMyuguSAsJbqib/5vJTQEyyJ
sidvpnSUpHeuG6o7MA5R2EiOx49nUCyuy89x2hyhbd/XbQhGs/aJd9qPTh9H
DED50ls2DBe6xGmU20GBNAY9uHRJn63yawLSOr5OXhYu68Trvnx3BcY193Ar
uiamDpTavmZZs8wIarMCH+PVmr9MLPYdeujxNDQcDSqgynBVfb/U2Ti2qMnu
cyq4Muyodq0qE+vMEoPrgox5OmLqZPg0qfWEklWfW/exaeGQMaM8FkR24Yyd
LnHYNcTw73hRG3Ci9NLFftAtEYHd/UoOSjz7Te28HHAlNJ+VEdoyD3fDP4gk
2mAQTinffXNueZmvS0+VU9OBljBGOLPupO2fXJHKGSXvFzUsCfi8sMs6pdJc
WvG8nC/8r1KE/3thnpTdAhe56ilhxfliqIpzykP/gBNMWX2R7YJ2fpzc9bV2
46YZzk4piRpWwokK4DrgecvyB9Y8vQxXdgj6zBRXVhOzpc7Ti1cqUjyz4JQg
iNxl9YFXgzI4R8IjjI8nzVcTueAVSK3/gGPnz0jZNxNxDFI/U9d57yi0dGqM
sTstjJNvgQ6TLPSbw0DtU883jGj8tEH8tEpJwYc6fIFnqSXLbB9hzy6X8pAJ
vylCau+5PfEtwKAc9Q48Y4E/edHIWKc6poxmA9AmcS/gXPYmYMmqrR+wnKji
WjmgEluxYtqeQDCg8KmuadVeDnFLB8NhhFu0PtHn53QYz17W0XRkQTsy/Lo7
bnvOrG6/XON5azywuN+RAHvZAqb8aV0k+LxNDMJgDUYjdZ5kWohxfC6kY+KQ
wPtihtteWyJBlgrZHiBlwfr+B9S0j3iYjVWyee56Pi6DOSmZTi4nZNPbU4q9
Qce3xwj5AzFXWlGcsk8U/5yNhiOhlC3516QNkrS8JHhZIfZ36o6LUtdd5piR
btLN3OrseaGXlcPCR8DvgGCGXGIT2lznQMTALRUpAVZZvQp0jO7T4YLd98cs
9LpKnIahI74vrweXvtmxogmVqLweh+Ds22PXrb25M9DIkhM+VhG+wKWGv9Ui
FMNOSeH6QKjJYrWc/CNXFDNFQnE6UTE6PDEw62tF56qvrUnbHuHUJ/+mPk5M
wQO/26vpQM7F09egYVbItT+GHxu+vjSxDYwaK/0mLOzBH676390gPyfi3HfX
3nOwe1yjjxFyaML0WZzycyb1wQjeH8K5mGMvQc/4Jcj9nb53dJNeF+ugzbfU
kjVlROhL8kTGAiGq42g2dyf4MoRsutTc7hQXI5Zv0XZFBEyM7FA+f3wMywm3
aDhE4s9x68FAjdN+CYKfNerjnQhkNAg3J1JwOJ/i/0Y7sBrHPD+LJ5RPvPqo
pd34s59jxFBaWbWYxbBo6dVsV+nhnPPM7M/EYo3C1Fp9ZBKTCPVMrNOk8d1g
Z8ve+3XVOhJA2BKriZt28lFBv058ipB8QyT5w4e0RFYYbKPNeqLZf6fTNP4R
qb884eHUOSD1Wbt8uCMMGWdx39GrjZoxIYJk+VeC543SkqSqSN7NEKSDVPL6
G+5JtXAgfymHD1CYFZmfhgiIUcAnd7IqAYwfoJQjlyyweVDiUGFVklISRqdK
jD81rlm/PJMC0m6LYeSwBlaboZPPJ6YlnUd5HaL+//+ma02lNS0c8sxDwyEq
JDfPx/AYtLEc1d0Kr4AODkfHCvuEyHUCsD6OZAHzCdp2tJay8gqPcejQ2uxk
BehojIzVdEPPS9v+l38IPhbyYFiTCxMHqHKWq+zCNWd15pODk5iWzuKbUzMg
zVLh34dyYTIkmmbDB9mWvsFE7mRoSxlpZYDpSI5JW/f7R5QWxbCaWu/7nGas
4kfxcaF317/6/GoaHxOOWIrYz+XuKHJVhWSGmsuXXX9y6gpUPlG6pySusQbO
ZifG0MnCUzElwA4f4/msqaSKwqsCotR97PwUnWoW0zpLcsfCnpyj5MPdSWOc
QTux5iRZu0IiQ5TjwM0ajlt6hL2ElKIS9CMbHJ+5ssfuveLzp6Ai9wRccFbd
AzLLN7jG965xS4NkwLc5UVjChQoITtrfF74MdS6OQ9HEUXhuwluHYLLFIOhY
nd3MDvFw6WZjjE1hPE0IoWKegZTXp//AuXLWPpN8FU5CB7buseUghdiNe/7l
Kd8g3vnyrdU20z6GEB06OmFwhQyU7KGiJjbPnrJUiyYlav8/kLkUebgWWeiu
rQFeH/6fd2YmQJ4XboYd0f2vr3MidAAG0ghpBcyRC23/Rm1hSEJ4xkHe27CU
kwo6KgRLDlKEQDRm8PDricxoFHexsnRsjVSKUZBnzirbi7rxUDoYJKNnKvwX
BBBDVhDHLRne21pmCo2vEUknAMTGhLqhGviEQSHEZ+M6I37xbO4P/uoUL0h6
c1s8X3Eeg3DoEzs4t5HIPN7ttqGRTfrmqjWl5tGNBbSXdqvHPbvgMViMoQDW
GJrqfAIG8NtnNcp886sLlMJiEjCkHLgJqkx/QfJ4x/by6ADId+nOIS70Vvd9
UIVXpwJ6chCYqMoKfBWOQE30w8n354Y3wJmr/DRJ0XFwhut7Ma2KBVdWL1a4
PPeLsi6QZyVBab6yWR7Qrwma2FBi13klilbwnYowodFksTKWMqNUckBLib+p
hcY7kjkgGUejJWTbOzeVobtApWpfn9BFpkiH6c9RPv4K1P7FmG6bHMeFpNRh
j7cW0a+2+jL5Rk3vif5jR3ULeTVJlDRaA+Jw8lZYNcJ5bnDNzJnhS7SX3j8M
9z4pQXJHXL9TuFcwPVK7XfNmm5z4dFj278KKjK/oOaleJg+Ad/o7mVJbkjPZ
mQKWBN6scVvwuUjHh7pETYwIrPpN+nYtKJdc/cwQ4MotUgrGt+Jnf2hQYl72
Pne1xAg/91lLwLCbN6a3ddWwI8jqQWwlVh5P+PsSnjr6q6pBjMwyB1MTnckQ
8A6FdY8e5g2O7A/ZEqw3BKSqcdA3Z0uX4gnzwvcelB6D/g1IHh5NkYIubWce
SQxxHFbOrW1Uva/q8YONRmkd7Py1d46r0ZD41peW7mEF9Peon6LEOdSNOZke
X3MdkZJZL8jJlTsg8G9/6hS6r2OsUepz7DWCXXnMj7Fln+VibkCutZ0v3iHK
xAu/mJ3dnj8UeTZ6Rybull8D919q8MWlYFlc6pMhYwH3/yb/4sJ6F8TlJ9TX
coesUEmZbAApyGwOIBEaH5e2ddbtTIC9p7IKkKDs2BiLRXBSJE0Tea0ZDdy9
oEQ2Vr+nSXXFqZVojfTlm2fQ0FfSp2c0HUHVxqm/TSD3q1H2zF5dVr+1Y7L2
aiZM9jFl2NmKJ2Z9ywrO5n01AYj4If7pmPWHPImznl0vPLS1i0JXxpolP4aV
gviT20pt6TlX8C8tEgJB/72VjV6KgzbkbE5l53C8Q6sI1xGGrgulb70mbHc+
RrG0rU0q4kn8RP/QPKAYDCGsOG02eoLbumzaJ4u/KJMKespCoMc9aYM5z9JB
ILN+H1HhS0sKHDqGwvRZgf7oREshSbq1td5QF6G4TcY0NZdMzxwtVTz+Im2X
/rNNS4PmT6wjRAUkyGp/NdzU/oKaiuE8adeus/9pDIAM/6uWDspUFFSwcQTg
3BHAdruR2qr1ctVKRAV6mF7hB13CrVn/Ca7EV6BBL+3csTaZM1LpIu7hOVdr
/3CsWNKNg8R/x/f21q16JwwLw0F/xgqFxPDShnr/rm+obVW7rHnFFMNUueK6
2DkQgVNjyxaYA4GZdsr4a7AYxkL2lq9UIu5RoCJg+vkaWY6eryzPZoJLn0jn
fuog3Z6c6InA1Smr5AulhHD9jMh7F71I6Zw3yTShUDLPBbF9JeGHHijl2Qnu
jBz7nO2zslwWptlQkbr9FwHtt/Si0J9+aXIopswz/5lXBL+tKGenEC7xkDF6
7KeleydzURUK7wolLl1mp665rGAJiOhGZgLbi9sNEF+ffkhGLQNrS0PjcGAu
IxRTUYEshYFRg8+Y4DraYQZKhlglJv0aBL5bbEskxl7bkp/4LOSlx0JOQvQz
09/dlok68lzSuzbGOhdTs3bR92uuTrviD7uxXnkWdpI32ECzLy3tJzje3fka
7YZ7bZbjKgqtS8auS3KVSEih/U5xyXpSmVQz9W/J7ABTU0ddw4Dhdg6ZiILH
T5PY19r3Md9hEq6pI3S/pm1SPsIDTgJEzqktA0Wc/J246vEkxRHsZpJUZXeb
CpN9IJkGTE4KGnYPBiJJypi/swdVLa2/oMoRSejR8762h7MbXgQw2TFlP8AT
QxtJnS+6tq5C4D0KH+jxmmBSptFsyL2BKQt7lq9I77o07a+NJx7/WQRsokxz
LDgiKVNzhZlUwirtoMSaRayvF+O9kCDfNHqQ36h0mcc+GGu/Zg7iQGcB37X9
vMD7SKPs7fRvJa7PkB3yKp7IfcSA5wcv8TCxPHjt1aha+KXSxb7iaIgWP8Ld
lCWx8Fazvh3O7PKsvgvBmW4RnCjjJsTclYGBVcawJt2arw7z0jIZnIUB4zJ+
VdoAMU9dwB8qIZT0rloHQyIINKVRzyJDVYaikOjDpnNLxTUghK0U7bQ/m6WA
JiCZBfa5axQFxNuUs5u6Vuca+cp0UFkNya2edyz1n5zXTzvGqcu7351i1ENF
lpzdkqCb9qFI36Mwwl0OqrqyZL4DulWp2amsvQHv65PdweU9bzLuD1s6sTFr
+u6vHDLMM0kWoKcODScJOagQ1d0snplojBhlkEEDdVkLPJCj4QidAk5nbwyZ
4NKwQdXK59zCr8282bp9E7f0jwy2rHWi7iCM0u8C0X16vwkMqpGgJUOdrLzq
+jgH8XGEFd4NGEkq/zQyen+0VVO+3/ogl6J/FMAtgkYtGA3er0wI/VXk8Krb
ly2hOxJKSe2k/Hq5W7ISf3SXzBpRTPJQi4vzreCzIWW7hDf04quC+QoFi+/z
uHLxlEjTiDH7tuq90+trOwlgC2Kx9QFvaIUNhHt5M1gEmsY8kIFKs7hO4kdg
IHqziH9MXWJCNaRemlex1s7lo6/UYM65V2t8aWyI2E4BNXsGCs4c33RovGMp
6zr7vrjbNGnEvOJ1wqHBz2StMcng3yA4hxjFddzzW0zycgyFtoNzWcd03QaN
UzVCufvdWmQtjeWJxsDroXBO9k4acH1oBCn5im+NUJ2Nc06d784mWtR3HcBt
LQpqRo614JbAEszQJFSoTIIgGG++iWzILz8UsLUf+hT011h3uW3j9sWh1p7L
tIjZTSwuO4mqyZ4200zoooUYqnuv1yL1KElqVQjlTaXiLGsJkNqM6YCXO82X
s4toI03Z/vnJ8kgpLNPJ+56bSVc1MLDibUbeVmqcQSLCkK80mb9v75e38mt7
OES0K0M2uin1U3Nl2bAsu4D4tiCXn95J359L/8vSPjMZx4u+v+84+Krl4WGN
BhTeIuBsKQWzJG3SATxn2YU3iaC85ydi4HQy5nW6nwXQNCE8gWuOMP4KRuzT
niSO3KOJf9va3vQHxDMNWEDPMX8tieLmHGFKB3P20sWROaMkKEcs2+gjHOjc
RJesmr5tuxgZ4fLpNQHyrlhHhUL0tLune1Dq87ZaItv0/6XLzafT1XJEUpCP
D9XYnA6hzOCv4WTc4tzFLaHOahJMlRHFQylJe2JPMaRvxEyMOENES6VNkH3D
dotiyDzZkZr4fylRpV0uhIWV/9DAwMvy1Ouqvf1ccjxtRL/Gh+HW2amzkZ1l
48XwwNoZPUsm7VL7aztsCdzhGveliUB715VmOq9cG4FkAaqvzvMpgkk9m0JL
PO2P9uhEkrJVhX9yjanl3nR4PXyX95gd/YXxRMQ4MSMWvJMtvi3OkWx8HoVp
/1ibQNWJClMAA4PJbYL7dshzZRw0GuVnMeHI/haLHgitwn62H3vN3yilCQDK
cZp5w4yC/1Vq7CxfLOuN6VSEtw+EKgSka1ht8YLt45yCq+5boA9dnKWW6BbQ
IZjhzI3o6YGf0wqKkNF9X1OghdwPRQR+P/AT+KAEhQ46Zcn/OoB+icW9bd7W
yTupPPYJikR1WVXB+unqsx3PTut/HrA1nMXR0c3IEwspqrhAlxnox7ticzxO
8nNdefza9nQnfL1Wxng/Ebk2/JDZuTe/cbPkSOCMnCWZM3fiwJLtQVY90YCd
Wr94NQgG8RPrq1GSqQnCs0h0s46FCCRF81W2jgqs7izyBvXNsC7TtQHdjpG2
qi8gfHMZo6TCe/eitSrdYLRfbC/oY7ClT0su9BYdps9HFfEWzcZBb0JrTRZC
mzAEG4HQrQm9K0wtd7zAQ79j1kqZGrmEgKRno/TPasaKunoJMNMnNMsGL+Az
o4fh16YXa0wlIjhQqgPDtle9fxrZxMpDZbmtTAr+P5yvZoFqLnyh1GKKZEZe
7fK6p5gq8F9mNZ4Je7tUyNNP19yugMZfP+PPKHdm2UHJgTl4YvmVkacbcysL
XJoOqZxJ+rtdsCv76IW+ybGDUs5y38V1f1dfbP04WTsKcjYaNAOCPhOKJ3Wk
sYKHq8N/nVNgxOxdk+y/OfikT6U55uN4tqK/B/QUg33qOVTdecIgcxTZazhr
v6v0Gd3Pq3Oa6txpZJqdaEHu7HwgydRdn6t1rG81kyr3Uy9Ff4RSlZW7PEgY
bUQlssZ7c743DQAOe8sm69Hl1ZFqb9ARZ+E8pc+jybk3K3aiG8CwXcVjZltJ
ZLBk3M+UMm+7IRHzFMLHS94Ex8IoC6H99NQieGVy1AlLDwLZnReX86KPyNNv
X10n4IiAep31vmNzuYQE6paYE50WbXJYz4ec2pD9qyL3eYiBNxAcwgetMWmo
HbA/ypd20sPtHn3WhoX7k0nb72n3Em6F5uKVhbNB5NWlHlRwu7udcYKV+aUy
YXvkjJIS0FCB8JrvR+uuC0WLk8OnRlxWF3IJ3OrmoKlGPlFFZykQc0pV4CQA
AAMPua9gTjDfW4CyWKXsdMnf/ZkjuVk+nOQtdXw53iAUWlCwUyTd9QsRwM8S
uiPp8u4kF5sMWiRutOArd8hceov8KKjTP/HRHH5A8tVyAMabfz6udmE++eFf
mMFB/dJ42vWonbn8klLwzXvnnCB4zxg/fiaJkP01V8NsxhzDJWCeywrVI7XH
xQiCukRpiwv7/Qdp0SuDFeqX6EO0HPn4w6Wv5uFhooX1eRhq+h91CMGBHuFy
4Zf5Vx29fTd9RZrOiyym4sJ58AjBHouORFnZ6gIjZnINgSPft4XYqWgi3ooQ
wJrG+zrDsnusZ7lsMtl4mFcES/SoCkDDmLWomu5EBecfbmpBH9Do/zv/9WG7
BQUvitTpJyGjsQLSxn+JaTUxFYNuPpC7KGAG29ljWU9yaNxrWbzppi82s0ck
Jl6M6e4UuQMMf/O9K0s73fpZsWfthZpZe+y/CutNiUmdw68/uTAuhoXvtQ7K
xl5cgSdSAFVXTGmoLtUGD6whbq6S4W+bvuDcudcLgbmZhBd53/6BKY93gXPi
t/0hZoqqO3sCm4WynA2wG1285ylNVcb7WS1ToKJh6KYXKFG7Tt2SK9yGJAWv
qmHzGBiEv5pX9Gc5IsTd1FUyPuOwclb9Fs1cT0p7LIw5HvnlXJ1oDYUrSGlC
Y6weAbBiqBqgH2V95WIye2RwKJa83+FUTFXX0EJXc+9bVAAgiFXqNb13y7tG
hKsKL93VBnjzB1V92cpSOlm+IqnYX/sngdi6AOz8h/iHZBmvv8tAWsB7yzpH
BnoWjVyz1fmOZ2HO79v03vhV4cyOC8wxlrgHZhJZf/BlyYdJilnBwAy8t7mG
N5aSJSyIWK82RHVLoB7wPPjzqppDE1LLtZfKwy3pc2IW8BMGSeMcuJhoZvmB
i9aw2e5ZJvI2F0E5H9txoiqM7hhQSXYEYS0UoxnFjJVDjj+I+guUsO/qr0dc
gCHBUyfhKyGHMbAF6hdrgTyBoKt8z37a1zAV9N0j3QiRZucAY0wQd52Tn65b
3ZLXQK+f9ru2TW0ziZ9fvg2xJ9rsdPhNzRuXMSs/jt2zaM6JxJiH9n015JQH
DT8xgV5e45MzCLS0mSGguz2q055Mks3SAhEekHh6sjhJz/VqQcLNZ74io5Hz
DWs8bFTlm5At7rph92cesYpN3tcxnfO7AHcARveoHihpNVF5nDbSuCinczRl
d35XvO/ywTw9XOB+i4fnsxOt3fsj9wPR9nOZkoNqWaUPzSgaK+TfnoAOtZzf
avmAdvgdITG+p1N6xJCrVX5CDqu0t5eDxDhhseaQdSrmEJtromLiuTc/L5ve
n6z/jMdY4XwrEO07Fz+Q+6iP42YO5LnkF5ESgcVShiwDy8v6WXjsDX3w9h72
kxT4pXvhWzphUY58HLDDlcYVWKBEhxkDQ/LVE+w7gZUA+DUpf91wJmfpuy3j
RC1TO84O39A9Mre/hG6Qsc8HKoIui8CkEfjhTLvHVOZn1C5qQosC7ZNhHI5G
K08vEwkvaUx2yRYYd+svvpIxuCeF74pZxu0T3lsH8MfCnYkRzrbNyZ8elDI5
C6Zw/rAd+7uVpS7uafBHHwhlViD5VGaifjtra5OVbSVdul32s8W3SmMogKS+
XzCHtfaXh+AvyLnaVAS7rauzdligQ38S6m6/YptQKAp5OJGqODijUPLHtwOH
6rNZQNQdUvGAP7w2o9prbnuRkH4rgRzB8WwX85ozW6IVq7aOA7mVlnBxUZDN
LIz0+FsmtCNDpsPbwSMHddxQ1whoEnfEliQYfRbqu1Nkyimr7HpldckR0PyH
JUSHYiNEvclqGPjel0NvlKMsKE5YnCz2ruCT9EtaB+aoXo/EFvTkidrCOUNd
fJ/1M3Bev6DgnuiOcdqozW4xWkdgGCnR0sbskgYyUI4nbjb6k0jEZmLNL9w8
wtnHVSAGKAn8uEa3IsyP/wyJbRoYk277j79FqoPX7d0zolMJxY3uEvkUdlaf
eWLSC6/KNt0DoZChwL7qWorLKVa7nk3xG8wyzEavA6F917zOYgmo75N87Tpz
8vXbK6fFeZfhc2q5WZYDIwT6abz2CC5cIX2ZSIoBwVsr4ZQw5TjCsJFioqlT
hDjn7kwFV6yUqYKG/8n7Ryh0SuUic1VZjrEW+DBVEpiUZVw6aeSZXaoxINAa
PAgDgnrtiDy5qTSD12JQLyZ7vZPyV3NyuO2J+tnHYF9vS/j7eF6kuw0ldxck
LJU8Z7o8huHvwh8ko+Uuo3tiDIZsQXEkQmIHip77TEVGa5Dmaxo9cPgEnTWT
2qbFkXtX/umXiMSWEhwDx3XVx3E5QzQbJfitRnqwxaC9zTUSRGqxHjbP41Cy
wa02/MiSrAKAIzkjkujhlD9OqEawkJgkw0ap1uWLgF7Sf9ycq8Kl+3nkrX5d
38rhzq+uH1Taj75CYmZ7pfRbpBoZ5EM4AZpmNaaI4MnNHHRAdVQhcKHD+BIg
+dRzTZ/GdwCHFf3c0WpFPU3T21dxxkl2mbQLxBzYaEtipimdPxeFes9Nb27a
M2ARFPo7oa1wGUvqjhWO4F9oKpgLiF6cx7Ly6Ke+vbwSWdbBFSDyR87Jiwqw
X1GPb87y0racQCN1VsPEozFOIADcpprIVboepTIxiJIOqDlVRgoCxzyOVXB5
dIaCMtv++E0643Pkcm/tZeZ0pv09sXxEGy/By4goUdufBB0ARW4li90KUN/i
TcvtL2JRbBFP6VrgGzufq1j1bNfYySA8PJA6rlhIviTKzI6fX24jeS3dK1mm
vUcZt6Z5OVYaZhRS0vVst78lAquqq6YYYo+GATzvXMtRVtXyR4xI/qffy+Xc
oSv0b3V88li5c9RDQySxP5RFZjWnpCP6RWDiEKSIz+pWYq+bv+qqmVrc+j0Y
jRhej5OIpXSBE77hmen3ognHx0iKCJb+kJMWBWQdKzgyZVzOobh/i/8wlVXR
uqCbvUG+4NK5dGqsQCdFb8DO9/+6TBpBGYtgZYDK+t4VLHPtproFKPI8NHOB
H9pVWN+NJVYrSjMzd3xpl+YVeSSp8FocJU47huPw3tJ7sPrbjcJoZQsqebt5
W7ewJlkZxZwLOaQ+q5YvIa/OfdkBs7lCoF58fV6poDTU5po4NEMWMcaflMU8
v02uWl7XjgPFK7fQLgW2eOj01KSkR+g8xT1kP1kEdifMHOedAGMULJjaCueL
BJOZF9EgdUeuqOQ/tBUokedrj/OI5tGf4iyur13f9lKFyUajtqKtfdWi5wnV
luI/p5q9tNr12QxhBDFx4DowxevU8dpSZ0b6g2bzRd00CQ11ykNyol+Fn1LG
1Oq8ljlOHe1SQBtZzuHeN6yKUP8hunScIIH3s4mMvKOT888N5dw0o2IdnUV4
1XtAqrw0bJfKauwBsJZ30dFm4LZtNu0KYsOQJuYYQDIQ1PceS02PfZ6EGPIM
0o7BghGl7agWAiKtc/cTZcaJePaCcy0XQRsQL7/lqI6pA2LDSVPhZYoU3f0s
ZVU+RgYRgDePczkCfN8cPwd8zT4SbEX5WOcN37zzFyp3WfiHn+UsHkbO2w6K
qvtHlJzVjmiudFej1C1vpBokQkGSvv/q8fDJhnU1BNTUdeAsm7X/Owl02LXC
gmr0i35npkrrOUQVHc2YvzS8neBK/grL28D9+Zn3VlhecjiqwH/fuS+O3zAn
SqbNt16YszaRmEMpi8YEYgmFlBrI7KtgDHPE3U+y3EB+p+1U51dK7BJmoHU+
xt9YSQLT7DAa5H+2PNr/L/nJ+ueQNcLRfdKaxYoTe7e+mePAjL//8YNA/npI
fHO4AVdJ+lxOI3C9MbiSLL1XnTyjQAfAafW7WpQmIxmi/brzDMHoVzqYP8+A
LhhkDY893Yy/58wxMOSBcL9p1wLJODcg+NA6u3w1M6BBAm1PlVvIUMwghcYv
R6HONwEcDgxiWI0Nug/GtzWjSJ00CVQoyRPFYdw7LoTs1O+HbV+1vLN3uYRH
VJiYTj1I0W+pHKFvzGUdT0Fo72ZlXEimZSPmVGRTdlx+JrhasCbt6eR7I3za
VpiP24Ds2kcMczekBwfklQX0GKiDNU8dKq3iEP9k414Pwnd/zD9NzYg4n7SK
tLsc+BetRTqIg68LaBqjA49bJI20iEoAO5ztwwPrZTrqdVpVRpXnqds/tLv7
nE2UOLz2tP510p00yQhwXm7URIXogvm35zpwNu8RWxi8QVtZA4xh/SKoKOw9
TrvGcbKo9gmGZ2yaT1CCYOsc6ej1xUupo/Gwi/EFxxPi35GAhwgt+zPr2LtZ
EiLgfhn3ex/Walx3OHtAz/WITluzuutPSqaPF9TTxUL7vNmTQgCbPOtGksNT
7MywN+rc6ajIu3feWd2sP7hlk8InfLMVeCv0txeZ08tT9ydezSh/mX37iPld
OQletEKfzUigaqxycI8KVe/A/8hlhUrpszo6/8dqbS6xMSDWGHxnE3+0sZB7
nsv0KvReJ/v0aSYZhH9rleu+xdGc0k1L1flqEUsLJflCn5GkB65glItTB6GC
Aar/80wIYg26RnJEQOrMGWH0NgdjE3bhZJ3QeKp1rr/l+kNecnySAe5SHqxc
3BbiPy7V80UZK7jzMiaOl2DbEzw4R7yxYFLFyHoDZr/B+R+fj97nFmYrAd2R
1c0y4y0bp8dtmHlaxX4YT3mxtLxjoxgJwjf3EMB0M88FDB0yPR/zKZHEXP8z
k8UQxh8lMkTWTZT1N9+/qoz2gnbYLObWMYHDNK4rB7BgYWSH8XoW784y3AWy
Z0SrdI8iHixyJIgZo12OSWvM+YI4IGeyhIDLkJK739umqPLJ3oWp+NrjdKsg
ejasEBiW5Ge+akU+7Hq03ltkJV6RQPUKyqFht3cRNHu2C3pEYBwHn9t8yQPS
NFJPZzs//v83tRvhEVHYyOlypiHxH2ftXEhKgwDDaxJSK3ZwqhKpOmaqgR2f
tKgoAnmSPb7/5NDPyegAs7vNNOm8E1qUeMlAiDWsktGgD178v4dsM5RRm/md
TXEphJtYxcqYlcsChvUxbi1h+8LuB7GJpQ5YqWqNVR3UNKPT+iOhRQDRV9rC
v0rxd2FM9endQkYoeh62W3UvWYyTjDiATxH6gYnTapzgR+UuSyHV/T1YcnHD
Q5VxmVdGvu57J3K468prCvJurYMSUxzUzc8Uq10DGHyYAwy/xhHT3GOuVNvx
ZpzR1RK1xGFLYbSsrhd1QxRkMDeae1pR+QUj/4hi9voFZ0z2S0t5IuLEjwjM
WoapGtwTOMFuX9C9Oo2C/cugRTiWpXL+D3G2okONK0FHI2KVYGUQvV1YWk3p
ayzX2fxQ+i+r8iPXWyAC3E+nQHEDo5zQAWHRfBbsvYTUZb7qufjnYM362LGs
5odpJBeBKL5lW9LgYCQx8P538+hedK5zjPevdRF6FaDjUpZ9aUo7aRbvVPEC
CGnXYPs3F8TM9595ZpJVwVR6bOptbB9pTK/lUefdBSQE58SUzbH5p3APVkG8
M3CBx61Ba+F+924qAnqOF0y1krMBX98ZkxZOTK0oPJc2/cmkMm+sFLrOF/jd
10t8Sa7rlUg4DM7mZHOKDW3Rv8lsb9k8sLdWBJml1IR8LPNvRUTX+lcKXB6S
OhBPgE3BOQ9hiLmCDRJFrPD0NbKYGfZGQDGyqsmzCdteM44q4LahT+aO4eTX
WNxqzy+07GfG1MTmXawLKT6BJcTGqnSmhNkoPQZTvP0Y4XBwtKwNC9eqISZW
HA+fOnM3XZFarg4gw6p47ho1LzoacIg3n4ObVDR0YfCzy7qpOaWfMMYIhB/7
Dy353ScnetFVqMI0lkRRX8o8V8s1Hi5HNRBq8DI+AszF+IfZiO922dEmVkb/
oLErs6PVDgbtAWKX7akE8cHmljwwu8bnv+ldDJxpOmg879xr+LYgzKu5AlTk
eEzl266v8/Dd1kb/mxtlsv6KmlLZ0w3v5fgvnZQIiNeo5O3wW5zm2Puw1gvD
YigBpOIPB8JVxvLWrLinY714ZXYAXMClSLCh7dRjzYZVTD38IJddWunLz4O3
7cXXQ64R02XI2DrvbTdTY7uFqm2ytJRMZQG6rKpQOVl6mfE+DXm90cx7w0DU
uEtVTLG5J9/t7OkC1w0tKnr8d9P6gOz0eHrMN+Njz9M3cbcCUSxFXP4eS6JD
Dd2wtUAxDYLg6cCEUVgjDG0a4OtLMsMnSeNqkltOlXOcXNtNYiDp6jWV08gI
foXNuuUBT7RGkg0Dp4GZMsAfO1H4MW59RcH5TAlFHqO9a8h7v932T2xKEICY
eF9TNeW65w40DfLsd7AixzlecweAhHK+8uAoaTx2li0p3Dt4u+HUmPAYHCKJ
4/ZiOCrTTAezp0LHMDzkNrhawdql+nmAU4vDOgYZlUxCOKlYNvFbZF77Mvx8
gRXY/hGwFGbT5Kjk59Tpkg4JNp5SbHHHQkCEMkFCbxWdZcUsxscJ4W8vkUe1
Ivdehx8z2OpNhpR3PQ/i2KubU2jIT396MAzlycraT7kSbS/iR5f0X+y2pmZk
wrRzCkc/eS3Fck/0nN95UxXjlbo4ntkdCbATfaXB3f1tcV3UMbwq/3Z2ff5T
BXCVbo22tGDdyE3AYptI/19UHkyl6E9J16nSY/RcvtBcQHGTrOK/cnFgpQNs
KYpTXvUF08pOwDuCTmjCr/haJaONS8N9B+gd4jhMSY1NDp40kT18NpAj3yMX
YKIp1JnJh6xAXeBCOReuUes1Zw+dtjUvs2UwZ3jBCuRZIa4v4r12RS/Xy1RS
GwxthFmlA9ZMdhuBdSdV1lNDhdO/XBv3OiQC4OBk4Mz7nwdRinYzPZ9PPrBt
UkelB67xJe6tjGxJymkGTDwRw1j26elnXbxFwSUdTY0tzotkEid/62q+pUdO
92wdiVDTUYoWcfumd/me2ILNSKp8SZkqx9JdCXum3IEet8vfvPZQBUGXtnpE
0BmE5ZkTe8dB08rAouAxVHuih0G7264h6D2UhuYCyVgL5hLWIzKqmuI6o4lz
x42p/FRAeXMua6QJ6Pf1Pb7XVpkB8bHbHz7nP0fdVw1u6oG5jCBEJJ91osfd
S6QYvWcNnaMT9X4lmAdZj/u6oPPhlcgdww51UiSPW3q2q+7uPqNQbhB0vU8N
nKJLxzXjYXlZ+dndH87eLdAD+IfeZNxaur8K25eyDRB2gli3oRZypV6E6izJ
AavQrVJrNpyaPh0qv02wqqADWYGl5o1HBMqU0jQonm7Iu318W6zW68cIz3x+
B0ZKizGpZFRMJ7uIl5FLa9qGl7UBZL+O0RTtsxfVy0wUoLqU/FSb/BiAKD04
XKkxnIT20uPOlOZiP5MoxBINSDrKNRepheppJHxzz5uEtUpEZsf7Y/bvlj5I
/FCAhe3hvzb4IwRf8TjFsu2l0LjM8p8RiXCdhzt7eATCDN9Ei3YnmcKumYc2
k/F0+0O48SFgPJuJ6PUriRKgmDr80YRz9fNPLbmA5bBHST6D3uTbP1OCoswS
PcZ00xzPGl1p1yIiMtRkD52tanMqqmclWaK5g6OUwAv1Rz1wilWcoO6Zubjs
av0A7BvIsJkV0ahGU+4p3teKf+dFAa4yKLl+1zoFfWvdIU3m1gEBoru76RoZ
jEZk5Nv/SIeyxKRvxbF7FRzfjf0Nj9vtdry3UsV6a2RhoBWTcHd4BRso5n9B
RUM5msBMTydbjWWBFJVPl7dUsu+OyFmq91icpYPE6HNK1gNd2UgqTUlXwvTK
3o0nbw+HQ8gmDkIBMF9+JmMXnZ7kpY7IaFJFffT+RcYMJYX4tJfgeflIluA7
r61ak/Wc4l6AOKD/q8lcM0EmP6LW5pxGxYxFexdFfctZgoK+AqQ4hfq0dtv7
G+1bYDEamAhFD5XIcDh4Qgx6dTAPTRJKkxIBfmK/BkJf7yipdXtjhFlNdWGj
g3mfbVz0qD8ZkoSItV29l91MTInUHEhGtlpc5XZujuPRQElqZhSsHv0G2cZx
1oNzK/uw2HgZCXvgNnzW581RAhaKMzoKc0sxQPjZLKMDF2YTyqYe+7xceK+o
ut9UwJDVZnwG1zuOG/reJkj65rXAfGqYI7w+j7mtzmyS7QT2av3DuooS4s3t
PVFTTD5LMFTV46l2aXX7IoJuJH4bcNoCWzXJxNxABP9WPpL2Acx8JZaSxYDg
eyuyRN/NHD6mwBRe2WJSZH1bbNHaNozgV1WY3mWTjcswZkRs2ydCD4PbQbmT
l7eW+2jceYTfTIxdZ1X5EvIDw8MjQGmyB/JGpe1mXYjj1YC1QN2GOay8WrFb
mpvgpiKZoqzkfxN4qIiFeN+0fUj+RRv07SgGAhxanD6twqxfCA3ZITfjHvmQ
qbI3AlHJ3GiLbL77Nk2pEzP7ySUAAbgh+fow0mgH5wg7PoJjFSpg+LbilmPw
Mk7jpiU9ahoFLOjyyIkLqzXO87kFX1s6vI1fsQPNwrJiD/HSCIzwpTnj2V3D
Z/sRjmr8cT5ciM7p8BqfD0d/zF8UfDN1huYblW6f3VzGzRMplNzN5yBo69jk
ue/4Hzb9K1/A7f9L6UgYPQDypKV+Q1jyCa4mn5TpLQy9HjdSUsDC5MZIc9ND
eMP1vyZX6HDmohNIGSqaefRELgjciaiA1J5krcNV6QPP+9RsOfxjcFasatMp
rnhiodaihMNdHBdpehfAxC7Ttm8+YnlXOr7yIbNBNXXrQStvDFTTMQcbPOAi
kVCGyk/eb4lgljGOmuxhn2oZIvSh2BsdH+JUGpNJ+KvspXOPigvmf6zPWtRi
1pxNWDAqBpFoPgvqFZG9UODZ2xMWvQoNfK4o/jzP7PWJ5nhNFrc6IUhgdUDT
vq0tb98OmBBFGoNGdbZgHDWQqIwS3PRgpjhpN1hpWfkf2eXgMEeyaHcNr60Z
3oVcb6raToLGHhpN0+9kH5jYBAEVLSim5Z50jdVPuQ18ttRDSpjwdcYkhcUw
dmIsWBSVkgWMhrvCiYy4uOMeO6sFsHbxw90EjFfgS/5M58ErG6DZqea6qFp/
pRvqKiGHv7KGlblmaC9O56ljlvgNjB14AzUF9JIAnSSa8a9vy0EWnRGd+Wfo
F2AtF9Lryk9PpJ5qPrQTQaNPnZujDmpBdZKHAnPGtJb7pDt3CoTUjC06KKHj
o9poqml2k4FjWks9F5NwWEY+9EFF3rdo8A2S6CCavcIf2bpVof96epvDF1lI
oaa41nXWqXpF+JHEXRA9SAk8jmjP8w6FhxHXmtipUuuG4G4g3faIoIW/y0fo
qFw5WBlgP+y5BcCJRtLQdUmVtSoIw+5VDHdWIqUZPILxrBWN+EXRsB1K8kTq
R9pqtgz4ORHttHboz8alrqvSW209AqbpHrXga45QckZloYfV7t0+O6PDtMqk
uDR1bNupkS9E0w0T8z9QPGvZSWOPI5D5IFXyd8nkLyFZK8ZcicwTCtVmZJIj
IqZETKlMg1200PVItqE08Z87aVqTIitBVNBhm1MlmB/ad3s4XYMXwGUmm7KF
qqmMGysP5TBC7TgSh9Rqo4VhImUDrL39oDloSTjE+XuzAZQvq8O2BSRsGrTl
5Aat2BiQsHkR9Ckg/UNEczvtS5smNedAZVjg9baJIOgNkHzrrjuik5N2Ld/6
dU7s6sbOGry1ggqiUU5p3nSKetMOz0CGS3Uzy64MVQkC/DQewlWIPTUdK7Ic
u0xan60lSXP4XbMF7nzx5TDFwb5O3B7IwboByihZoqbk7EaZDrIUw3a6f/wl
XyTQAmnmrvSCH7Bouuz6tAHxND+angU/mWzewA4OWxTcsu5CI9R71s9Fqe66
ENxarg7H5B9jb4SKwpVqVZohJt6bjBzt+X1RBo3hgbiEt1Epugpwq/c+67tl
jI1vNPytHZc51cimhiMvdqeNU7h62Uk9nQPv+hItJgh1/vMb4Z6bHSuGKLH9
yaw3adxZnmQvL0St0abnX6+Rv/t3zyDyT1INJeIEBenzJM/H+63vmyWQAaqs
faHKCDCBUEdPX7mM1oSlt5U/+QoW04pJRQ+VbpHTo6YiRVzvejrjiS9u9PvP
exs2evF+pIJvwnmpaiQh9Nf7xfgAh2d99rwXtAeF5Fh25AHieVHQVyAnVfis
NixDaliVSr50YXllCYEdYSfunr+ma6vZ5I8m5rI92U+GdsHZ4wsCk2Fyx1bN
vxBgxleh5oBtBeJDYVoKJmA/J3/4iiOhefsY9HU/Zo+N9X/wZN1wCzCfWTdf
q1dqsut+bIJH7lq18LMUyRqRISosiqeUxTNoF6N0ihVmnEtJcS4JHGgO92Vk
I0SjihT6F74fO/1CKZgZPSrdYU392aG/fp5AlZH5JpaG7m/yHOMVIAT04Fer
ItQpo/DkT+KFcs1XM+zl7CnfaOJz7FYxp+FS8EqWyhYnkCPIu30j1V8Che7m
zq8w9shNI2JG5sHmIxr+crOwREJk8srxmzDEWAGb1VwTuZoK21ms24FyetQH
AI2t0Fvb0A/z0e8fBYEBZcPnY4ZNeKXSE4aPDJqYdpbQiJLRW6EtTfuT8xiN
nLHkXMDY+6Ll8LhuKKSRFnOeeLuB0UyHzLWxuiOyOvJPEwjTkBkaTUUlW1pD
87brqt+VPe3jEZQqMaxApa9r1ELYMXldWY0iL/Q0gUYuB4KmiHteozk851st
kp85ZpZhs2CfVQGegeA+NQcL6KsKDeUuQK2CkKptFnbVYvQ7b0wvKshgzfw8
kaVOAQ8A31WzmWHyYoD3uSFB41v2xOputIf8Q5vkTjNqdKm04JsOe23K/pSA
+Ux7Em+qRsCVHqfOMWwEIRLgicfq65W6zYUzRyhBENr3rnPIjmQTSuQD+FgI
WnJZYz2v8sIiwHXKi1dUUJMSUgg27WNefEhz+BV0qRRgEev2uqu/x36jq0vb
ot6ydsl8yzXwIG3kUTJP44+4qA6C/f5uLh8nv9fB+1QOujv1vUnRWyaXotvF
4Rqz2qu0UEV+HLs0hdPUmRnoKHcqw/DX4ocP2pCsSfO3MhD4l23U3L1dkkja
bh71tD5Vx+T4h1J18Lr5XjPigCtcO5yTWZv0Z0e+myfEeXMv/3tXYDvgdqmC
4pBbdGjb3HuDNxlrO+3l/UQgKGfmtODl4CPTePUzCsTZQrO3xQA2FPShcnZw
KGp2Axm70zHslsVMnx8EA/yupO9Y6PoacLtsz0gwEhB/JHRzat1HwoRawx6p
DgDLsTAiSoyZ18I725UQWPs7bS/8QYhg6fYQwWmOc7jS46E8LnWQFF6rtugg
5HlcSN4gqLTDs8fxO/7eKaOBLAdSRctc2HtHTNeKuz3qwN9DnF0GPSI3T/YK
+2jmn6r1KPLTeQzLOqs3d8HkAfoybXJJVDru8AipezQvjK4QYzCwRan2xDDx
jEtX0BDxYoKfpeGoHlZnPNQkyIGot/H6nnY4irm9mh19gCkcABfnt1LqcKI0
OF1zKQShj3L8uPuczLB7Hhv4mDuhf62tAejGfw0TFkm5DpvS1J+6uHT5VcMC
9x+xPg5tT7a5G3Pgg47Nupx+67ccgAtuJbLKEC8HS9hYN+ECaTneG9GWJDt6
2FhCsiV8WqRX0BTBstzlo+4jxbpna51qxjlHvawEozodvzM7cDsmn/FBaRY1
ee2kx/bBqOzrGpv0pBqTzut9a5sfhTbzPn1IH4Gcti+xQhyqkp4HDj+B/wc+
zZ3auMrd8C4KsrAxDDE3gOosbNeQ2T7Pvp2hEHs6GSkX6z2XZF1DDibNKv5M
0VcOkP5D0hBEKXhavoZfzUdm5eqG0npyn82U7yb5J4a5iTwehWlCEtaLZt2F
cf5X5tDY2VMA+0j0DYZgN2AzqWgDw92vvni6OoNO3VIdBJheEuC+a5QofFth
Aedi2YF0T9Ds0varBdn8TXJKFipTwUUnmjCme3fTdBti1lYbeOZHqdEeKeiO
nSg5PZIbHbfgl3MFLDHUzCcFlyWxNxg9tEKB//4LoMtnQUKesvLGpD9AA3Pm
dpDfa0V1Bgq/MoeQf4MtAAfkvDlyuiupQQK+t7Z9VIJun6xeipeQd7TDrUI6
siP6fXMYzCvEOoTtvEB437BthLsjyMunG1kckhnbCm2wsWJvQRZaAf/x0NIe
jlyPfGeZpgWkqPrxaObAaiGtFp0LuSg6I/su1vqgwFbjF1LLm5D6pdgzbxCy
QTQpMb9iYpBdJ8P2Djn7HT9qSb4hmXeP4S+bgVAVcvfprL+bKU/Pk7Ntmm0M
HW5Z4Gve4n4AMSkX37Z7HzzIyJbS61AfOwWFir2BOWWAkyN0WFUhDRhJWFiU
eaSaqFEixHI9qEcKDTQBtOjBUHZvBo83nXBQ9wNjWlMTYEWV7wDGfSutz3Oj
SA4yedFXUk8eSSoXOiLlbYbxgVzDmAEh2xsmYG6QrgRCaz+2BrlI/KS4hBV7
RGqvWMctcEl5l/7hhGpzJFCCB4JbmDQaPDkAzQSYMy7jo6FqfD4l2ks6vUuw
/HKtOo7RcEsUm71UL+aEuAE1eHVr+8UmpYeds+5LNT9arX9/alekPwATSPZv
w71YKfx5uJwJnSjVQ+TepGCf3I4hsHkcHaOkfolsyF9ZF3oaMXXd/CBayJ0e
2Wy2YByf+XAxQRT8GlXuvqnEchugcbTTAl+kz2xsSZg0lBfk2S9dhPgWupYE
rPc+aUMSeuol41s6LbntYLq2H9Kxxb6gpIMTuH8Q/KL6w6MdZia+9+AxTWir
7klmtL9P8S2oBC+wRJOhgAFAureSChoEmEbdClqWr4N+oize6rGbuyUk7Sb7
UtqP6ugFQ32g0m3YkOIqMmkRwEZJKuAOUY4AOAu3PbkctsDie9SMX9WoHkwS
D6Pp54ZBWK5ciKhNIZqlVCcSzBrlfhtn/1LtkQobXKKAya0loj5obRGMVXBc
K38tweXBt4wNUuYmNm3mGwg2usI6EDyzwYkdna94cSeNvAaeL0H3Gihjc9wa
r42zqHt+NG7qQG5KjJ8qO4fQ6+h/yNoMy3ZH7M0F7u/tG9gI+kAyhRceBHt/
C4i5pkmkmBkEkMbL8QwKuRskg5Gwg2EOfulZqq84ANwG2/WYQiJOcMIXyu4b
+L3rlUX6qtdm9rFWygmeEcFsbA7uHTuh5L4s5zoiU/kYBb5GTJp5FRjtNBDa
KB4JL5dWlGVHmndzbqlppl+CRsX1i4PWO6aKT2PJxfWtXy1/qQW/538jwINY
wuXFJbwpghPZ5Fs0iPt0XWPtYWBoFp7TZqEFB4KhryXjOYmswtgyp8Sfv5md
2/f+NCe3+gsHp1yRwPWR/3mJwZIteDB7GjRitiJpaT/u/OadQebNNRtVz6th
wjRfidiwKCTicQJAQ0PqnJ04d7jEsqhg79Gs70ILCHJzL2xniQhNIMO6dSg4
+QYqR7aEyLU6N+4bpyLRy7eBXISxa96Dygq7gneijyNZA5iXQ9QI9FLayMSd
1snPvmaJXsyg0P/7+GrIhjMGC8xE33ndvt8BsK5ifYDJlSXXceWq9NGck4Kn
WELOsl2cFCdXJjbJLIrztSM9sd4MlGODOvJ3dZDlJmXxYTMaIRgUkvOTNXVb
//CQl6pudKFSn7Lp7qVNxJE+dvWvZnF1t7QVCobSZCZxbdadb22Xo/+NM2Dy
Jr0DcI3+/OQ5njhBHJlDsE6MOpYQLLOQHgDRJBzvdAijZ3nKuyr6LAn5SBOA
DUH9gauUp5V3671i+LxQGNNIb382D+wipBc+40haJbz+lEWLYi3pxb5bDL7Z
ELwrZHeiyiu9dfl684oZevHoYWUCIsIg3yBhhnLb314TuzZd2k729hJK3kCh
W4hhrXDgV6fKinj6ckrbqix9GuXcvEA+n5fvzZh1mV3yfufxjZD27X1g9Zql
Pow+5Ti3FBfVju/x7yrV03Aygmqju3EknuMNhPf+sUMpRUyyozl9K5ZS692o
txQpmAd/OBhV9YWsvSauA1+3eyqhS2bRHLR1hoIkDV1qj/yR9RoEgl1ZcYbT
Wj1uSNO5+Y5mN7JLpNhvJufWimGkDJ0/7qj1TVusl4dXihtVz9+beBiBOQ16
WLV4xVCcQVZqqWv7b45MoOSTAWJGXI3YDKNLY3Z28nnfepMboTGql+yMHBNc
oBIkeu7njQoU5CmaqC2qsJRLRZ8LQoJYn8qIHLZzGMQHsTBU4foPLBQCAS9u
tgHhvbp0cLuBdSPRMBSZQLnFbMc3/XfbfDYGFuCxdRE9Ha1WunU7vUL+6WB2
4A0LLZI1jwgXwmnwfwtCgYtvQ48rBJsH4DjBzHrMGBoU41F2/m8D7JmZIM2Z
2rvpBdJL6+p5D5K2d3aLhzVn+dbEI89/LWAKTX04y9Rb3THUUkI6MxTpMuW9
2tas8FgDzoqKKoS9/2VexZCLDCRv+M6xpJJ/g6hb2YcUVZlk0uWy+Czw3fgN
aPa88ev4FM18a5jgmH44QJdjYUZgv/fnQyrX/IB9qsxBUqxkS1hOKpO6DNid
Cu53sbEQuT/ZkPsW1hsAq/0b/dNTqPkpW2KsC7CI2UTYDt2gvZGzTVsR2zzE
BTjbh9AdbmX+ZlMCSzXw/BC4GBEghUuViJcLkerHKMh7RLG1tbTmOaQKspvv
V8zzzz/bI6g/xEhbO7/kpf4uY02kVbKUokGO0FTHZGaa8v5usLp9zvcIA7+d
xqW9S8zJ+inN0zyYuCUB3TOWXby4Isb+VmzJ4zndVrxbUlU+daEucYEF+HPO
Z0PhcLzbYr/98FUWdctfEkU2UxlQXRqJTa5XdAasMTQ4Zlj80u8y8JqvRFBy
XYNuolul2pYghQdYXQ5w2PvNCJCgPHt1ti7S2tooGKmd6dMZ46Vb+TCBx1Ye
PudiIKRBi7IYNP8xUYSguAsZgwkY+3wG1Q/RT5J9L/sVRtN9XHIIfUE9tI36
2Gp7uZgZAMWt6CCtCFe68Ook3+In6ypFuuUzsFHDtwTlGqEZcxc0/pJimbYp
4yWKFmXtr2vkdDgnYNuBqFCJ6csgT79zZTohX5Jm5Zyu86rbT006PrfXkqFd
Tp5c//edMWNBGbVGoimc3cdkwufRKft8K+oPdjOBt7Yon0DBNBYjbnbAaGs7
p4WeAOCYePnzRwXKuEL6i2KigH3i6kBO9Ao9PcDWD8wm2FQbLvCbMpWcJ0vh
wr3Wrg1T/ppRHo/zPrOX+XDqW2MXdTpcK5KfVk2hpn5uK7ONfbsrbYhssmmn
vKt/Ei7K+bsr+D7xtVoMr51LLPQOd/TGupdSz0UkIDoOCjgszo8GdS1LQqqV
9wJ8/s5yAO2kFdxxj3/gQmthS1gVl9xKKvL+Zy387b3FxgVWDe1QcaSfxcC/
4IDF7bdGjbY5AqgIcP7zm24tod+oXeZypwsvZ9+s7oXZeguRrc81dmD+mUOG
ImPt95STwhsAyqNQB48osC/ZDfbxP6CgrZRaKJAbY2dEPbW5kuixbcv39q4B
npKZ/Gb1Hq7HbZ0qFxm+3xzI4xGDtZkMW1hCpLSHjz3dC9wbu8DLXI1i5jO6
YldlbWhE82K4E3tatrJKFb9hB4l+QCA46Z054SJF74ah7nycyRcwSDhpUTeo
9LLurc/XNzC+4xGZzbhXlgIWLgGM6D4SPO6HUSvB9hfk6XQFdbiosykEMPXX
mJXzHdK63t/FC8VE2nV51K2o9bLM1NcqHhdIneuUnr7rxFzKns3UPv/lD8xE
iobK0sthf+Kr3L93SOwxLeC+SxqfY0CVcdCzvVWesXFF3medZRArxlBZ2isj
5I8GPmR8uqjyOp6zSf9zyrDejXb3l9nwKVeXEDwbLHc/LtfoMs5VIwJIzAwZ
D4KHE2AvrHMbarfXtCdAotOeniFRa+2NRuk8X9CwNnMHwSJc8+ESIqodAMBv
GjLJM9PrJ8o1Kz52Bkg0sRmGzW89RXM6oQAwr2ERWh6CuwVUIZx+rHaCCh82
ezed4EPaaBZV8gBj7QaJNx+YdPWbfuGj4suI8Fx/kHkEfbOEOLXpAqc/I8jn
W7muwv3KfaJUNK0BrPrxOhDZlC7cKnQgXckUOdhEunMovrpGkaWseDB9Vr2g
Q/eOGtuRBJrIgtV3FBPS/vMhp7UjjezxpWgddCxUQzHEmqA5j5Uql5PFm9ND
qVG5w3v0ApcoEGkWC2jIXlexEE19Zeit366AI6nPVsbIK8iCKswwrMIWB0JK
5CtOuL7QUgyDMudaQ5q6o5kLqjP2O5ObggI9VfJO3K459Qg/9U1eqmpZFdMJ
vmJqIOWt55Nvn4Xgl/CrzfkdqplmFsyvC4KxkWRSU0Zt3GkdQfXIV/157meh
q0LypaqY62xXL54LxRU3krAfl/To32tHRvqyuvHi8JyF+JSNF1Nqta6DoJgL
ojNyxJwEyjyYB/WPuqh/aJg5vRfXrUNPgmaW3/b1fpnJiJAGtPW20MGApvqY
sbp9g1NM/aPXgJPJ40HD7BHdt66cPWaK8zr6kyvHn2tKKhVHzNEoAMxFU83f
ABdaZh9WErn55EziGjrkD8zNBYMckorR+jz/ABzW1N+itlaKZIbJXwSx0WMe
3cQOD9AxAmqr1AoKWdUT5dKKnqlvYL+pIsyYFnMN/SaozhN1i+Byt+MDkzBZ
Fb4as6Bjg3s6Z+Sb0M94DrEfkg3uC7N7q+CeGOh+iTLcUyIfTt9nlVDl0g6C
SIW2i/BqNikyOqYYcIs5RNiGfxeslEyDUXGNAitev7dJrlGeWhZ1m27yODmX
FQqFTbomxvJb307ZDYwbjvJ5k4d00XROnRzH3C4OeL2fJ5nV+xpb0D7vK8Tu
iKeTW+ALYTB7EopfrP/uQ9Fq7nEITIpKCl6FlCOfqt9QC0xG9PbJDOClvEfz
GqFB4aVwJwv9BpZRWlzyrzPh4CvaRsLTqZZ6V6bFUjW9uYuTrAYagDE5Cpxl
PfO8zJye1x2EvQ2jhYsr8wFoKIxHY9PiGVvQAh35zPV4Wjvq/lzO+hM8tCYN
U8CXJv6ro/jIjF6jGYzM0hKOLm0tYvG/o1iq7w14QfeIX9kGo2F+kuL00Nna
Yp++NGFATfHc8WPPhTLLQAelDr3hn4IBTNVP/t1zy83rNzxTPIQNf8SSR21g
XQbBTrWkegTE8Os/t5dmKCm4irTMQViTop/qsKVYJgANI3B+b8Yas4SpLCwC
R/E4fPawrdcxEPDG9ktVD23E5r+8UKZ3bC95wbEI0r5msad7STKrWmwzStkN
eZkRJKlycfqY7DZms3TmgaZVGkMH4x/ghLJ/l8CfPNNA8q2HbUIdVkwDQ5PE
cSBkAa3r+J/UaBWNXYOccW2IE3hTu5NNvSodGX8czBAeWHUlyjinLlO9PE2+
Y/uAeKelT3qTDJy05G3qExF0ppqAFFIc8oJBFaKQLN31Y0RK9knvkoIfNK0A
WJGOc0cn4bz2qqWrZSPMVUifZFbZRawhgKFt5bVwPR1gXVHjR//1PpGjoZIw
wF9vCcm6tulJLVn+eOdxjKvY3Asbe2dmjAy9oYTP958IOpFUz6tME+LiJYYv
vWNGj5aMFholSDGd/vVC2FRFXsTXnn5kZtqqqTWhBumxV/UxRhmnbShRhgIc
YjUsEWCGWeE+1ictj/huaep4C80huuq5pNWv6ZHg7wwsiQ2tsEAfqIHIjnRX
kr+XXK6LD2NGOBBSDkes2rD7mRvmIFAVXE55/16krl0kHe35MRenyZWCcRx+
XwZUm1k6gsQoKEIIm1OIjJdEdcRv1WiZaCn5PwOBXNu71vlxQJvERE2KdQLo
B9nLDOvSa43B8fSo3Y3aH5+N+Ns6fTrGydb1CP9Ypv06+tESQkfSPjnT7t+i
BvYmnJ3vvE/GSxhqrHTwxFj0jcvb9NABbL7ZM2G71p48HOGhoKMGPH6YqjjC
XVwGZ1A7hhKGvVjbLEObW0fJYzMg5cl9q9N1bXpWIj/SvOnUy05aoqRsqAnD
m0cIdYfNoujlpOGcOw8zZPtSsB4QawK3nmfQs3YfNoV/us4IQi/uQrKLBEd+
VK/0r+pSqZNnjqunwv4ltn5v+xjAfARWF6u63x7mUroahu3bQfQzRDVXKoM0
IM/L0UN128LDvP3FVhnJMyZ86uVQ87FUdS4bO8A24Xxvxa8RTi9O2qU32mva
UgFsVH+PSWDhW01BdRbn9pOfErItE6eManf6I+k4P0Noum3goLw7NmVYxBV8
T0BeNpuzR+T2pRfFIcDx1xcRBarI+Q+JMqpTLmZ5Fg0ukO0Q4RmDaRQRb01w
kkTlgyeeHV0a5vb2SnT61iqqW+Gq5Ae31y9QEy+kPpHlsMNEyP+Ys0Dn7kMs
jbkz6iOvEyXq41dcbnQWK19Eda/02SZlAHPOypva4a+4doJ/X5/Ev3C/pE8g
TMtuXq2ik27uT/AZ1rUv8jJjrZNnpoDd3YsVJ4u3LX95D7goDOpTsLbK7zAW
bVO1QIEJQ+27Y1Fl7ZJYN0ApV2TaejsqyQ9/CA16zYOs3b5NuAjSMFV+PLZF
3H7UuerSQgIMDmzN/OETCuY+H5zIDdGxp/cq2Yzn33Jm/HRBxAhdO5+FtSfz
Tr8rirbCeTtg/7aVvIjqmZP5pqnQmT0MRGYtWJqotsFEpxCD3BUHjWf+OS0R
agPYxH5d/AinuXZOZ5aZ6dHmbOwKa/KsLY9DGZmAbEpgjtBqXL/vBCQ6dVX7
xXFhWzM09P0Kkeh3UAmXQBkqFoqXB0d/TvQ9IhePKbtPn0yfTwRR7Kh0jyUs
lCQeR154nb/TU+UHgma0T6HncCm/gjZm3z/Jb++k6ajEPDgZwnoEr9O6jsj5
bJSJCn9x5rjV47OzvT1Hb3FJR/VvQaBDBPXp/wR7uKRfYKlgXcFe9UgPHq5N
wuEsyfmN0wye/17zCJYGImGfEvMxQWjEpeHZiej43zYon6ikJwRxuVlDpdKw
cmjEX+Umf5Mm9aOoW682l4Qi5hPJdWvR8SXQ7D6gwxhn1XF2Y9bIVzlW8i40
QaMWpokRu5amtVKTM2HnleCHKtziTRaNghbJ0bG+r1wepxxA+MSzjRu18W7O
TfgsuvLuH32NBl8IYozatZC7w3/VvzKSOqmQ+zdPpyPcoMpn8iFMa7YiKR/e
E/tCvUu+4PcieHcVEAkR7lDl0MHYjEOO6zhRL5qI7TTpXTZr7azmrpQFR/oY
31+xk+MF7SN1dUl1sCu2o+gpDRL4j/5cOj16xXX2sfGWVJd8Cnx7xiew1e5y
9yEYYsS7OF1tCwvPNoiBXElYKjepwjE4SkmONHf0pZ0Zcna2ky9e4CVaSwNt
7d9OACmYEZqJAwlCBwA3/X4LluoMekLIfa3JvSD4yewjLqzQICFlIcvwkKLL
a2XJ1B69Rsdy1zY5lvok9otNI5wBNG1TdHl/UlykPEsmoVAzLpluc5afJQ2J
y0Ogs0ecHWP///oxlPR6ZCdzyquWxv3SV0btE+XPVw1OHbyTcqIscz7CQ6Ex
kT7ilxGyTKL0Oi6diG7IWn+3tt13zh8z24Qc0XLu5aNTpEBm3QuqiUvVEMJE
YemRHdLeYDAp6RCzKyEsHedJIjS4IXsEVYpJ8LI7Lz06Mw/3cExgT1C3rt8c
dK65AGJDx/6FnTovH4Qbwi7Dg6K3DJVUVWvEszPmwnxfuWcKPyxDoe3yNKMj
ho/OvBedOSysK9SCwLXAwSn7iSD991CsOxqg26+IwllOsI6T5fZcfM0l7RDy
kKBqr0gisyAaBnmFZkJIIr8TihrAglLcssxhfJgu1ilCXjb94EXMtmDtBZyj
hZKxZT4Tp/ZYHNaBNDB8Hcc1ImHzpuzodwInhSdz/fBJwvoQzREkLKWR3AAw
U50ykBmnrIflcMBCKPm3N5+nsmS4NVIhGHE/4wFxqil2zxf+tqlYDaCyOpoa
Pz38dxzxdVzIEj09a0+SrlCN2WGPuYubFZCuyuaSG4bCVr5dZWhH38v5QWlp
eKYPCgjtIs9O6zXZKsudDYE08S3eyI4eFInnvdMgIChot1+Hzwz3NUZEMmVp
zJ4qfHEk0kxugwViJy2aTY/oK/wJM0nNdKt6njze0A8LzsFK5s2ktosWNEt1
u8jLhLU6ic4+H2RUVCoIqrtjqaoaH4m97JkvLz5qMEKQm7Ua7EGe5bpJAdmu
6fLFIGjw5AHlr8PFbkDZeLp4ixxk0KptdPR1h9angq7CzY9l5C2YftPOtfvi
jVm7yb2AYlde1FLfd9MXF0kVXvPL/N3rpCxMO/ujZD3Mhq5fpggTXo7W1DRT
C00hMz1Wn9gXsQAeLqTdXyilHGJ5gfMKVY2QVOV41bLwKseHV1ee6A7q0ntg
0vHg2vYD2PguZ2ibQHai5yZuRPhhY99fqGb0V3KPnl/fi2qBvWB3y65tOK9Q
ZFGFYnbXzRfMh+RLdQqa4hL1REHYenrbkNmu6UPnJVDwPNOIxMtz4gCN3na9
eEclf+db1w3BaKqiHWCsxr5YW9eIGeBG4wcXrpJSL0+Aa/GqTauqCONNiYNK
gW6jfDqiII6a+yveIxst/M8wpkwUOG81CBVey4Zl0JTp44JFMg1ovF60rbDC
gBYoedyFi4ofc8HoGbeVrzLlBSjHOOvoTz0RxSUI/qDwM3hFC9eMi1O31Rsf
rj9WdQCaE3obWmUGN1HJ1GjzMtS6tqZ3NcqvniinmTeI+eVbeUsK9o4NDmsh
eWY/HbzCxkCBZxiYNsZmmUT4P2UoNXQdi44uT/9xZfbhRLzJKQNvIW+TzzbN
vjPNGBR0ixuUaumxT2ChquzHuP0SSWJKIorD0W8TGnw3ltJcTvHyABTTDuT7
HMuL7du6D3LSO6FRa3Dhtxz/HVOlwEhGRsF4X2UEEn7BQu48F3QgM1QD+NLd
Uhyi40e28LkjBZUB+3t7xOlnIYdDFDsixW4G/e1Czdt4VFTUBmhQ7+LWSzuL
tpiEDPHuesHagmuv2YwRORlPJLWxpU420yAE7XmVc1EUuL8pBMuc3Rim4Sqe
GPISyr9stTgcn/u0/bjG0nV89LejbPJOWvowKKmq6HLsp8keG6IY8wNSwsLp
OewOjhCWWlapRwypwNvpJ6xZiJY5brS0mrdjuTavUOjml4sfMmcjZgOrOGSg
jQMnebJvbnHTAVbcMd0W7k5GbbmLGXxpKjE5wLXayMgidL+oQGx3+9cHYhM+
SRaJbyEke/pyercdBjQ/V5ezLSDNg2NJg0cCjMMpP2pF7q/lPdnlk6ettWxw
KbOXI+yoxl9lJi9zbfJBP3JzbBIfQB4nqDdrSN8Y4npxtws6gkGd8AloZiJg
qkOwdQWnv4Q0AzuUSaVYXbGFYMRVaYQAwgND+hDTcGTnZ2kjIL1ZByDQokKm
Q43ojFT5OUBHk0c9EX5tJy3p4d2DkAnasV8bPIgpHRQLQdWPl/92mgsrj1yf
3ba5NTRgRzdag3Q1dbXynyibyye7Kjyzgv1zM1cdMZkRpwXsd5KaxyE3So6j
+X7HWGbeKyHwLkRzS+571o3MEqlZG0UVIyk8VUx16JeXryoSvXAZ3Yp9uav2
zguW35BzVt5CLJBQdIOiwNE/bNQLUAmKCAeyJJmkxPL8gTwZeEb9HuKJBcRB
cO9n6cb+kDBEHOhZHd+p3qDu3KOEVAO+812gmT2gNhPUzWkXyWw95WMP5gNZ
lN2cYQQfI/hmuCnWi9dZiX5dzaHWl4cy/zYVQx0GQMJyti1+ZqyTPljqrkIf
GvipEz9cN+VwVGZC61l7wEvUrgsJqC5omfDadt7ZXj2Urt6rXCKQWWGZosAB
rPl4UH6awaslwLe60hxUGlZ/zbxMNk3ZBZeKtNTaez2Os31xbkAVSG6uFn5T
FZR9yX5CmohHyToTD6ixhSWTeJdKJnA6EcJvgOefE+UbNYWplN1dNK4Ff2f5
7HtCIGysN84FwOdRJfaWCFYGB81ZqsCaVvLWFd/FMlvDyOALm8OhfUSL3eRe
XxYdj0HQc+Os6WvqV27wMGfRd3cFMYcRjsGbCpZlAcq3jy5jKI4cftsFdWh2
SrsBRJB7C0Y4brDUziEohFUvRC0pfdC5bwq2EPr0UUlpUTTsdGGFmwQaLFg+
UoTeL24MeDIHFhqra+t9sbyWG5kTCYX6LsMBl58HKTryXcX5lG/COG0T4jW1
E1IjlhlStQXV9xX1mOICjMh46JZQnB3AmZxC/+T9D3BylljOGrwJgXZP2BhV
9iVv4uJm/GnE0VPRb2iEYth572lMe+vQIQQxwTB4CCSXy68j/x2F6PmMAX+e
ibkngrsuFx433r6MpSHnqaNiDSNFTiNBsHiOUcUNWqdKfqwUdtKyW77tyEOS
YRIGAKVVFIA+g5n7rqBejHDMGkvsSFSiCQCKyu2vpWIJIK092Vfth5+T4WsU
3wUOaXXrIQ1JkL2pp+xOAkMYLzi6TauoLSDUmkPtY+E1g4bpOj3EVUGK3g0q
8IGZ5XPOAAIhPROr1vg1kpD2kK0POi1lL+c/n7EZD/R3STpYn1RGwVmaj4QB
n4aT3UFZ+5gPQLsEtuOvqMv4cC5WEtaiHlIWmRMDFLfqMKCoalM9iJWP0e6b
MAc86Qs0XVLb1ZM0so0CLjIP/iJ/uN6gvXiMPlcN6IElcXG0fPVGg7GeRHop
xTHHzSVLnkhICTOgNI7PS2pp6XzgvUsQj3iSDCJgofTlcAIxsQBVkvNTOfg8
24YSJ3blfWDbI4BUlMBGcG6QL59hf0arpEuMToM08oJ7aikslP68t3Cg+2BB
zfoUG4ZdWfs55ds62UKDxGVytFITTwkG/pOfi4kBIxypZeneg3wW2NfQ1gsW
yTWWyDRp3xt2Yg44yhq1M8BIDX56PZuIZEbHH8rDaAFfeUGvo4f8WZH+c5/l
nZid5X/UWwIJ/hHr6W1Lzn91s/AutndK8B/+gAyNl652AfbUjjvcRBrqRw1k
ZDkmBrCRSh5A0mTWljsKcV0mWsIfrSbmDm2LgXygyWJOkYwumYMEEbQUE5zV
/41vyIcXnX+g7n7RKEkrb6hD3Qta7SY1KZccy9S2SnBVP9mJKe9QJv0pCGyk
p9962UORAIWP9nh0b1F0JPpWSZp17nZs6s6/Vaf4Y3LgKKyeNCR5m+aH1slv
uV4Yp0Mih3GqoUwZNs8zaOb9KQn5IzkGRW4yn0VmY8vnGtF2zbmfS/VCJZEw
OiJCy77ckz8V873rI8yYhcnBrTS/Tz44zl3U1YFUDUJ/w35H6bZRd4BIcDUS
0SisATDoX6aP5W3ONIbjFr7lYSbcCa3d4Fnd1zKlcXnYMB8Ta+nfHSkJjeRG
o/QTMuPJ9A9V9sl8XKE9WXPZrx6YO3451EPFMdU5ccYSo6yFQGehZcoQr+Ga
oX1puM7amuFePvm9FqawzmjacnsIuKPWqu1MtpAaWS6upWX/LJVtvnByEyXm
bbQRiPt7yitw/xokhV/WoWlEsGJNjO/2zBDv8mR8uSAW4wjRAhgjXuZf9CSc
+6dY46na0erjnzswWT+NGeMwxMoTjPC/VDrpGBMk1UsJ260nepRcMHCpYfaI
LJyxI+AMKinwpVLtpp6qDxHbPsFYqsf3uLVPI7mxYlDs6Ool3tJRXANIjlyd
b7BqLSyTIUkSZUMNNqqv8crEa9CywtgfjOCKaQSolyn1Gx9YNBzP00eySYRx
NRAsSntktqcXRI3hhcpAqJzFo5BYJ4GsUGKyMObHd3Jk8NRoddqOCuEW9JRP
gBnPTb6Z+Pwkm2yITORnMQvS4xoLCF1/0xGJNjpXrXyVO/UdpX1uEmOPE+6z
uqRPpmTFKq7NsrqDTWJeSaiZUjaRu6TfQVWL6uReFA/V3RBxQlGF2fJQ5cYr
hnbYKAXu3NU9bDJyUk3gni1V3DDLtMUAB3N8l4ZjAqYvtZJ9rZywYXA+phdO
H00lj/9U4/RtDPP9pcgSUZndIf1WTNSfqOYlrve/lQfrLf5XLonSow3EUWqK
Mln7XJYYba5oGjd8imGZ1eQ6C25FU7OFZM31tPvPG1ZL3kEUqh6b7cCFsIGh
QUdO20+TB1c433LWBN8pQd1G2Wu6eO0G7DzBc/N2E9WjN8GsPTc0j/tLEq//
8BwtVPZXqkt8GidAjiD9iRDiArByUUutlSl8G/KYdIoZs0VNx+o5nPVkV8wu
YY6mXf+mKIYSw4OQajUWw6t5+YYU6ZNGxFGN2yAcAZeR+A201NkoLopJ4qJ0
+x+lH8N6L3VU0DmJpT6xeqf95p1GgCRpOnd8zLeBcVv5sfUvAJSxkSlYCOda
sp6/fhLOyq4Ag1FaTt7yEZBPHWdhVToGzLn/IxBD6h9wsNYg98XK5xDxrgfA
tQOr4nD2a1+jXNQG5fto+PvtIMCYCUGXFZE7jEXmXjs3ZOXOztKR99rP6vVx
ucxfrpzYGt5+pzpUrT8kYBhn6zTZE6CFKH/RvDRoCkdXnAQz4qgA4xUnxtlf
nsi0/RyRQsFC4Cq4xFYp3nacyA/IGbmBihV9NjClluW2oDxsNrSFw+pnBCsd
znlbyguBhgRQVnFkK1bihCVKud0fAtZcPBE3OcU5yEydMzyH9wuJZdmv3KIk
7vrB1Sliy9hNM4sL9+q9Ysoz3EsaK3Rh7NCUFatanf7TD08mYwwfmd/QBdlH
FjTqi0QlyDdABxRy3q+QWU1onG5/eBb5S7sg/RSz9ky5h6AK6N24/js/9r+T
qWCy8NNtGiU03S6LwF4wpFvcAYhpUDp8pvoWaztgUASu91OCemAB08rADBI0
WAypHB+m+DmFkDOA3666v4bcz12x75yiEcYPf/B2dVKUKN1vTgUt7NI66WYd
7/8DY5vQlz/oopPsWb5xlSJXK0TVPUCDg/3O5auro6Juw4UPuFNyxrFt4yDY
wUSdqhg2Btwno7wb/wqBrTvKxQwsfuDy54iQVrnbarU3NexlGFppoVz5bQT3
Ngp/Xc4wOoe26v2Tvg9OLgem94MVVzr2OcFe8bP8rVkWA2meSyZtPRqK847N
lfWECKiKv40lh3GzcM58P3VPZ+raaQmOdLCarr2W4zdG5DeiWtWNHlFVd+Is
QLs5HnBqAgqHx80htzPQHKnvOLkFiVDpO6ucXSq7dKFwQ/X5rNoJKsH2rKeF
zHcs22cxMaT5wUC6BVqz5aI8gKD/vmCMaUIb76g6JYs87C9DpiY011mq/NlI
Zlq8hFRXPhIq7TuT6GYExJ+Coc/iIdHTHFVo3QCC5X5px7b+KRiIbYam8YzV
jVzjTSFwE9m8WHksv73jbXnhdUM/7XlAESQMpyAf3j37Z6CL2XdWbscjj/Yx
Z7Dr7vQjsHjO9jQ86RnMk9GO+hBQQTTY7Nu/goBdqUQRC9VyhIYsyNqk89f5
DNQjSqNYChRUe/HT+fB8wWk14QLcPmSFfXJ1PG8ShbY+NWBIWYK1y9AfUs/E
ySIdVRumfmRtNEsmqvI7dsLO6JB5FF3Zn7GhvXblm5v5E0v+iq9QOIfhW5o2
qbfgPkJeZP46GGny35WT/G2MdYql+muFVHLwiG182Zx4UGLns3b4DoihiRtM
iHuKeyF862OP69MrmQ3WOJdkF2Et/B8GR1HWK9eVcYSnuDtuk7r4lpAQf60o
Dax+CyAhtdhWGzop/lk+V9MT5VMrU1PwyATiFg17KRGG9Ai4e79d1wZtbhKG
/T/E0DK0gZo9H7YQV+X2Ljx6jPkVDCP+kmZtvgH7c2mvT7RDNbnUScqGwYGJ
fy3ffx3pcsrunOw5urm40Myr6wrOz42iIAJmA5TpuMC8p/JYYTnfUjVbX7bS
pu8s5sgoxboGVdT3YyMsbfcepu0o73LLiQctkfAHClrGb5TvZu4J2wlMWgBb
wVD/TcO3JHibyYdCsV8wymRf57YZ3ETrfUiRrhJqI+w6nhtfYrSb9ZB6UkKN
W4M1Q53wFf2KbrC0inBhP/WCWONRM9DnvW5wHrq+o7/9/kBwRSvvTYW8fWMe
IEdfxMpGhe3hYPZPUBTy47S+AJ0MAOVCN2LIM+iSYvOqQ0gsya3+MavkkewA
iltlTu3eEbPrung/bdJnNo+235bw8yCvrHVwA5gP4cw2V0NC/0TmEP8PeyHS
onI89/FaNwtzLRB7K2CIpRC/bHhXWUIWypPkpl3+EHXctBOyRdO9rbuGpYSQ
L7HQzxAFFUgsndBG061qpqMZuq4JvawRmxtIb6ns0YbtUB6DBgIqzqMOty9N
C3LsAzIaXwl1wAvWrhrJJBPES1q99FnQtAY5CZuYZOO67Vc5dHNj6sOZKYTV
0mjOHib4NA8JLF/sFoC1QBBvOMysyQX7MmznhrHy5j0M4djYKhcU9TEFtGRJ
jL35ahhYBoHjdDXSKBguTbuxo2lMrDXUSgu1hJ4w02vpZrpq5dv1Uexv1FL3
28xXuVMQbgZFL9LXVp76QAiBczThS9pGKg5SqNNobldv/wm+SR4rYLpNpYaP
pHiXbO0IZ4z3d8jG6NR+2VOMbzx2fxhEXQ/O2uoOZGH3kj6EfPRnKgJnF2+f
I2ovJu1y8iTFkU/r+l45TtSQ1F0uBLNuNf381N7cxR4smI6M5+3XnRlj7ESg
NYXNU3jvBiKOmqg9kZt0bt9upOIK7W6GdhED9fQjjUfQHRjICRC+61NepRmf
LOsCL9gNIPX1vV3Y/jF7cJeEdbQ5/w+ALqnJOtH0wtUtmcOdKq1EkD2TT3p4
L1bynCV8fCcewnq8sKnFCXpB8vsQEcgPZaQ8r8tD/vuu1wueJ6GelE5un3uh
2QSP7HtEbYjmX3pZSb1iDT5N8Vm+64oOLmQFmZlKMcNk57EIaMVCLspL4AVQ
GFEQ1+bg1VQ7EwJrrBCQd2gDzkQsokMzSczziRxS3qYBk7Unvvqv+FOzYwcQ
gtsL/29lEdZOOTlU7NPQm6JzD394KUxwshlq+29tWuswBkSTSv6jCDdIKNam
UXbD5ayq5elGJETOZzkHDEhYh2NbIdZ4ldfHU1c5oi1Wgbe68y8RgWBJmzvT
nY9llisjzP+paHq0KaCCIviGf/IqNtPZKcvOSbtL5GqmhFzzIb2WXFvGsZJ9
xmuKl1XvMD4fFt6/ZLb2+g0uug/N4ND6gq1F91ttWLkB2TIpikX0+oyqMr3Y
BQ8ZQOrH3ALm+Y2CZYzoGFVDADIUV2GjhCUKJ9DJDHwLxrMo4/dVj6OA0b9N
SB+90bepLXaKsETJiDDvvYi3lfYi0u9TsafPkpv1qD0dyj0n5OiYEF4+aEMQ
sK7bJKqPs7Uv5OtVuvxQb+sPQ62HBW+HJpHIVwzQo7qDdmunR8m58gzKUoLW
fTOCTvK6z5ZmoSwXXdw8s7qgK70UXAoMyvqIk2BORSNWffpnGUxkegno9+BD
6hF9s/Z2VjaYx7nSy8uCr62kbTIrg2brdAxJ2sa0w0XLupMnh/aQrW+QbE+A
67t1+d8p6TfpVKWrLwoKAh7Uxz9+pujSS0Nv/g+6IjKHbz1A5OUyNEfdNyCv
LtXzu8JsTmQgx2c+/X+gTu2zt/nYrMzjWz7YtyYC8d4Q3B1AwLF1uMszdjCE
apXgyJk/aoM2HtWLmkjlAI0jpRH65p945xPkxE06Rw/QV2rNqDHwspQrp1SF
c2krSZh6kOCDDknn2IjMQpbMexYOtzzaf0iuSGAM8u6Pg3YPccWBTTH6HOb6
SyVHtN4WmPre/Fs+8oaD7j5HjXSCF6gTDzeI0DpeYciGMDwaUqqYl7NQ422y
C2GSvHXUsvIw7RP2Le4gxCM6mXsNy97E8A3Imd0p4gsObbow2o0DV8NjVWqd
1QZbWPnh+ae1X+PIlsITUFFRP5hP2AJjyNpETQ/28x6xXVOZxCXzMoObqxYf
GQqK4gU8vtNhTqk7UVP5D91G7tgeT3RAYMK9NDKrTbKBH34LXRCDheB9+fai
GV9X8UJzGAodYqbuCFkV4CMrITBhBEl0nqdCK2m4KYzA7N6vBlEv/uc70Et4
m58UuLRA1Bp3FzcS5hVS7p3LeqBhZRVrxCW87pvHvaqfyw3EeXl5KOdP6NEK
Icja7iQn6WWrBtMi9tgQZxlg5UUPllfANxyI67cnUE3LPYxSU9ncvzq0La15
UcO5xcmNreO5/wzDuOIgyvRFF4vBMbfG+H9Busp+QG23snaIRZN/1hz75pW0
vi6+bOei0YJ16Lj8mB9fQ5fTkptTYTVFH753pYlDTWZI4CdjOScxBLLuERsa
EbY4D44eOH2Z2PVh0ROBJadLXmEVeAghcT06fhMDA7m9HMPz5y/bGfPIbR+v
X7NBFNIAkI04BR0pdc/xm7BS3rx8dWn2QHkXTnpqSEcRe/o0WwEfCXMtYUYY
8xz+cIkDMEd/lX8irOsRFbG31kj8W1yntkjSuHjQkO7EXlywUco873SDOEk3
MilLPhxEO600nw1h294FoXt4ZAzokT3NCAKnCdt0UbCRoqPpTIjgfhqs0PLr
obn8suIh7FFTkVcBVwl5tiWELOpRX902U4f+1tI1KcotBKbtXXg0HGQeYdXh
zBcsJkYfI8sk/4Gcj50LEM0ij8FgF81ttU4++KW/qe6/w07lW1ZMBIjMf/JF
U9yYVj26vhbQ8EuptBlpy+yFh36gilxABqHntJdlGxSPk3Ny7oWWCT3ZFHBO
M2b2mUTRDJqlbBTaWDU55F2oXjm4KajxFq1/5C78wGw17/mWoWoQNZWV/mdi
yLn1Tepc99qHNuYDhuHng7G46gGMRijhnggfRYUKhVv3CIurFXimT+Ezj0eW
dzR6OvxAeI8SQmIGqGej0KodSdxbQyyse7qQdxd55EHN6YsXHDWNkXRET4vr
WEkq3SulP6ggstAE2ys0hqY/vqtrq/kuerdu6ZHOgqB9ig/YcnbDso7jhwL7
QdRWyAcUh+qC62tqQR9R75bSFpZ2NKCV3fx/b/QmPcmFF9Fic41oiRO5c5ZL
f6qkpYCE6s10z8Oeo5P2QX+2gTEhkuNhKKiW8UP3j5rC4ZJYREWYLOKuBiOC
+ezTjEps62e4AAwASkoNjmhR65WXraFHlGToerToB9GZfOrJ9cMRzTeDSqVl
RGG1CHPe6UsbGs/TbFvAf9YfLoo8UQ/o4Ya9Uyj4G5BEANUGNfTU5wP20mOa
LCpTKQaX8boIDGtYsBe1hMDONiy/CJSpDh7UPJSbSHdzSYN+BNLZVLLrAGu/
qq3XxLSsB9twGDSl/dUHJdqz8C/CyRsa7GREWS0tML34q+QqY2DuiPAgk6M4
zcIm11f1+3deC9HILxLerX4Niw1FoakZA/NnmFI5EF04b9przODfox1o6S9i
Zqqlq1n5VvN3b8hEMmolLSuupWtFiVY6CEtI5gvi8sFKCYtSlVc2kqoa7thr
YP5k32cCo+/WMpBicgbmZFygqDm96+HvA5OECPKPDIrkgSmOofB7frC1IVjD
6jK9Bi36dow0Dz8s0MPKlzvbvkBEdvaunoeUbLZeeopFLecoIhBBno6t4Abw
wJF1aKdhGRbdgXEhusHafmJBS/ExnBiQbU7LNosoGwMDONqWLFUeZw4hJGqe
CtiaTsJ48dLxCYPVmFxpQdcnwV9Sf9+dL/9YahoSL/9f4IyHQCcyGvzbgVNQ
8r8R+lQ73P5UBWD/fVMQvp1s6pcWh3qs2UhKkW1VZXTiBOW14TBnm8/TXgh0
WFceFZF3ZGBMcoFHTiAvUN/BerNehELI7zJacVBaQRzj92bd85PLSK4St3kE
1klPXxZcFTWFhyRbZxJDVF3KmQI1ICwzUDk2peRPUg2t2QEoWQqxwJG4PKs2
qVuL5Lk7O6e0J9JTFpvF+ERT+bwmKlHpqmHzkqMmks6GtRWCoZK7oJStihIz
O85wFul5lfxdCAxM67DzbNbCg5gk0oN9qmnOIKA/Sv4xzieMPIGnQZCdpPTQ
d2ML12F+ZV6XvjfM3hQVQVnZ0xgH7maoYqBlyV6OTzMIfX9jQ0DfiBC9vEcV
a+iXU7pD1SvS8hpvaZH2yKaEA0nUpI1QNa0iWV1e1NBXfiu69McGrJIZBfTl
yaVhzcNf9UdI0aRYuRumrfNwvbkqhZJv16i8gqcBNeRrp6Hfou9aZQpPjixT
5zTtgHUUbxyt1zy7/mEW6hQdvmyTEMwrGec9+ypv/Lvav2TXKDDNpzbBhGG8
CiI75RuUccMsJrV4N9ucC1hbYAL+2YRosDzvILxvdiihW7Sgkd3RwmeRcu7i
vx6TeybqLXlW9gMUdc/x9OJkOOuIdgzzRQwTE8jmpD/c6+lyNtvs5BJNUFdc
mJargs/i5ntZBqmR6OXTJpOgJ+BBBbr/rsMYJcSKMMZkg1g3JNxK16zrAvPy
WiSc/r3AxgrAXBvwPBybiTugXb6gQre2QX+Izu+BLfproR0vd+Wz3zPynpFD
5pxqLUTAljPO1YukRwnUJFPlMRtYaY4qGIM0GHWSnCNZlf3WhLlvOeKymGLb
U3ybRf3ykMf4C1vPKdmwVXhePRK7JMmAz25Lv2TcWfuBQo2pei4ZN7vN1vpL
4HIIe9lxnm7jeGggVdDpGcCOxQ30l3Nwg17xKEGZuSy50Qm/Khz+BBAZIQuI
/QaC1s292hKd3vTXUolO0shOw7oxR1mTNc4fwxYHebof+g1PU5SHDY97lvX0
VTifS8xPcYpxNW54Ag9iC+pvN4HL+l0XwCQahM6F03IjHVceJ/oaqFnRjMdR
nAcQZA5lYiheTZ3NEFeCxSthDi6U7xk/qvAxyapXP19a20MapTIt7HZS1Z4d
3W1wVnBVe46zyeZC/fzihfAjonNRq49z/ZbQ054D9X2bg27TrZGtdN/5qBpu
6ryeu+iSnyG/oyEbKgVKbMItN356p4/4OR8GHtRl6fSOqPx/GDyPgBTOIjsp
ZOZxjuIzj5l3B0N2aJKBgyFgR9afm03hoO4qtpdPbaUCs9V7Ui8/4vlAWfu7
aOPuuzCBmVGSnC4Rnx6Crd2zOO4xM2bLAx6MH66LM8hyUYgWlDK0He3xbMxb
8GUV57rhVnqKJmMcnHvdrz2BS2yZb5N/ojH2qQrRbBQtyM6NI9RHod6Ix98y
mGo3IvwIJ1VvMM0hBm5tE9F37dTjUPSad6Rnb3a2fQvTVaKbEty8vhX9wU93
YeVslmx8DG+NTOTLkCjgRsfxx2r/6uu2YI6LwTa62+Pt/IqCT2VRjgwUVqfq
czyX1xjWf42iwSvjAv7fa5BvCA+NkxqIHp0WfnSZtcxkJGwgbAvgfeAVKieY
jpnDxESZ3VQ/u2M8hEFitRNvLyzdsQSYdht4TvDYJQU0FM/XdML+Cj+qZG+p
BD1FgOKzmkQghRp52WW0ZhOq1+XLKMEvMFF4jgz+UryJK8tj+X+hwiPOkj3O
caovN6ZqOKzHhPw8/lylskjVq1uvN+1Y6gNMUxtgdHwUQXTvfv6iWLmXnWo3
2UVtoFYLKI3bSGgt1p1rzM7H0Hu4dsOO/etjx7I7htoIBrEu6qBaZH76xsjI
znKXALNuG2za2YbORPv8BQAYhu4HJh4uiRicP2F9BMwcVxBbq2bwVVW9kbYq
bcYAyeWSdMXwx2HG1TS+VZpXhTIFbr1U9Y/AAkqZhuH1KzEyKZVVjEoSzO7e
1aF4xK8HoQY8ar68RxkRrGw46sK+gRsYGW317d8iEUH9zQ7fpW4wINFQV40I
BjQO+8D9u34EAMl1ZpaTRldGZaWpw0xcfMGR2B0zt+n0bk30RCTmy2t57oEN
X6prAl2z6f5zxWOniGwUfYCHdOPFgCiTmLkla6hml/6egEAbCtJspkU2QaUv
UMiaT6b8P30CTF5bkspG/ykDwMyUkpfVm8jFw7qJieHQdq+yBIhRac5s5/rM
MhazqS8Nr1Q/Kwk+qTtYDMz63iYBHziLOJjeaIA7FQBxX2QHSjan50AVPaTU
BKSgC1vGp6l2gHWFAdBlUO8hb6T805AzdZu6HR3Mjva30KMiQwexLlfZfvqz
Z4DUn8Vy8SX0aqZVfDRI2ikRPo0CgMoYOx/XqTlWjpvtLCsXRxGwZaU1fS2q
Wu56yKdxW+1HqEoI/gu14ojK+mHr624bp9IBGEViZbwvh+U9Nw8+9ejqRepm
3WBjGL+tz2ZJ6FiCiYgVaLZuIA9ESkZq6XToBzFdiVxCgyomFB74b8q/339z
D7QE1yzFUoo0yYP2VjJAyIevPZXo4C7hPpyA4pLI9Yvn/TwSBkQM4XAeZCnr
5zkHCTxRNxIaWUOzgWMrgdcTjmo4PLOktESvcMAiJX1fZ2WMGpu6UeSIVUW0
olUcvGfAJQELR3kY6vObdL4EJPPf+058g2r4fylgXiyRYM41RZu9ucBjOt+N
hmjNyY0yHvuhyVfmmPtaSGuTXkoFBBhGr3aHWA4wnwFWbIHL5O+gmu+rpU5/
e/vvmflXBE3mS8CsZ2yhsM8yzwO1GBr0tAjs5NqthtG5+bsnxgmlvFBNT1ql
U56wh7/dW4BAS3ICZneugb4L8pUYO1IALIeMPV5YiYo4ly/cQT4pGg0ooH1O
grCq4EJdgoKyxmVFF2LLMcbFELXSiN7JYWoqBUh4vuv2OlIzSUUWiTSytEWs
n45Ha3MsWWIbuPDdt0av5zoOCr2bhOAmeYh1VdpBASyiKVcYR0tZdoC+IjRT
++/2DwXInZnZYOTmeA4JjfS/ajCfmcV6eyrAdp58TL3eh/XSn/PIs+S/OaAX
Cv5yPnzuZ5/+5LbRz4WxYw7McNEop23D9GrQ2ZSvRrB2gyp5TBDCHG/3VcM2
cDtfc3KMKa+aq5kcu3M89A0uvN80WfkAQmxn5HOwu8dvvID6btE29duNdwc6
Mcmg121RTL1sQyilIlB/t/pqfePwq46+1QBjryF7wnlfF+qluSWa3LKbdg5n
/8gLk8BXYp8CfmJIsbjzYrde4PqST6KtkrVFQyN1eChEI1QOxmFsj0mN5CuD
NVj+5qGI7RFNLjxm8euUDrQyDj9l+5p3H4czoaHNCniInM9jqS+PJrv5mZ0C
kogjdkcwLpfmfchvG+zAX3dl0cNpYFLeQg2KgGnGqU6lTHL0ha2Yz+6KK2Ur
M0raVlfHklhM/72Nr/4kNsmu4RFSDYdPp++TDueLYadFArRFEPf96hPCD26t
ZaRnWyEQB8nrqVVFD/4DIl0kK414AgtaKmsfV27DDirt68qXKtbbVdjJJsGS
W4Hq3sImcPC5zhLFAEYOwtolxdwMjzSy/TvVI87Z/nh9K0sB/wWezTNOm7Ln
vPi/1ssdj4NroH2nTjPrzyAeqnEwauzE2EJ2CUcZLcHXCocfbR4dOfLnB5nf
mJ3lP150loetkDEMIgvYL9F0GjzzcwiyZzWGOMA8q+ShOgb3Q6sNQYqC8iJh
0M7UuwWuZePyeUvUVxJ049842+UeqITr8/ABHYB9wQYNzbagXDKi48m0805M
ARJgVwuRecubPs5oBphZJtt4GZaXOuxkZyw0ClOLob0ecafEKQZ+pwtYl9/4
DUHF7e1JKX3xQ+3P84QXKJqzPrjzDnj5bV7/xLm+w0JaKv1pHfXie3RkLYVY
l1AMlisMhxrPDE0kxS3T+hVVgnyELCOrB2Vu0ajRt/zhK4DbLeQGeT3Qsce5
rt4CeUre1XbjdNrFXUB/jJnWL9BI4jkRJeYcG1h/65i522hRPIFv6EyAevKL
02DcmwV0JjQQqla+UhdQGZpfezyPSifOsOLvM6YqwvlNmf9ruNX2nfQC62CY
45won+QjES/xrFLAe8AY+8Nntgfi2cjkkZXjdv7SvRBGL31KHW0WqOya4Vy0
ZAAMbuGJZFa7Ch+dUZJA0BS23ForFook+VHM/Fqj7DSYpeS88qriVgkBEqos
JPJ3dvOeIOX8YpckeGO86PJIyHHqWTX5yvzwq3Sx/KBx3LViFHviBZJWs1nQ
rxrfa2Pu1dHOa1pyo9AMYaQhsJcz6QXLgvvo7xkZAYxZ/ChpYtxn0WNDpGBv
yPtV6eW7COV1S+2y64VVOyI27/lBmGirLA2KbDIVVWDjWoIAELBkv0IziCQX
EOfroLl6hr43yshrQHpTvmnYJ6XMyMiVh5O5F0Sz6pncNK+xYFXtax2rafBE
niabcPkn8GZkIgJJxp7+K4UInJynHopNOMGZrPlNH/PF4vQLz0ZMJXwfXgHs
iTV+eTDgC44rCAqQR1rxhd46FvI5OI6yVPsiT9Am2mCcJabH1nweKO/7TYt4
FybNA6XWZufi4ZQr733IRUx0AsjzHyNOEiDnEWc/7FwMouzyUR/CuyBkNB50
PaPUj205KpbQCQq3PQeC1LfqE2n+DxXIZyD9q4CMJlM2HaNGlbPNop2fcB6y
ApqKo8x5YK1FvBCofji9GYAQennGxIuGvLjFzR9d/PEstgg2AvwA7nVKBc6j
4ped1HIlEhTqYrRzddxzXdNfKp6251k1v6qziDpo0WvcnQQYz7YmC6QcUPqv
mU+CSgkp6M/kwODNycm7zrkp8QLRwzlZiF4AunGuMAd0bzq8uO1ZGj148Cm4
SQ8XqeeSUpzMmbXPvIL7RePvqiCrINFDuukCKabBPQ1Mbnsnr0I0j5f5p70c
xJRQNRSYB3HndLrUQIwcFiQAdkYXtFUUgum2d2SZrUHLa8jbt0Lyg9TtKUxE
08TZnXDBzYpJp5U9k+JSMQOE5yxcYkCLZtI4gC7p+T8VzLLdbuOKHYHwbiUt
l/6w3sIc9j/uD5H5tilVImH4Rrx+p/Y5ctlXiy9V/85dC1FpwxNVRjlHjjl2
FAC0szJSnkVkQD8mWycSQ5y1ERrWWbCa73066unEVNDwbxVj2mssT2PmXeCz
1r4BU6YspNU+NwelwohtoiTJ7MhMwIw2yQjs+BU7bxpuUOuggxqn9mrC74rK
u4ILUoR2Ha6njUjwBFmuXZ/ej8xAbmcsDhLywWiVLDj4hpdmGWpBXaYRKFgp
99ECuvhz4EGoiXHJaIiwWRI3+2I64a0UfPek31hYteDP6b7lPs1Q3juwvMKg
jdDF3pUdbcV0NZR8/JOJ2AwOr2uPHmnKhvAHugq6Iy0DjpCL7gRa3pYHOBzv
Y3WCB2l4Pcd8TMek9s/W1of6nbN9jb4LEjVP8W1Ok1cFZiXdYwSYGphglCMm
NhunpxnsYQPaUL4LmZJ6tvchY31Nxfh4NVv91rJ8x5IDawsQSxw//JPziVZF
GW8K2nRME5YvfFztNA/pFytqMsqEYsvycsTbUhR/R/GlJXppXaNwvOGhPdOj
y07ApDZBkUefh7YBjp4UpgbK0up2vSPSldkT93J6uqMsKmIKjJEParkRJD6+
N+KeIpfwiad8uayhVksUlhQq+eFS2JEgHQgswB1eyhZl4v8tVyH2heVfSstW
7P8vE/ahHrCRvRwWYPttfJ/RSXenwqyup4nBkBGG2C+ZElyw68P2zJp5I6N+
dZ23e8mk99RgrrQ815a3fXlMdOBXFT7Udj2ijFyv6cFA8MOfkUf7NBSoL30I
w0D9nWautp1SnxQe37AKq86Nw2y0Q9gFhFgfpqlNnavLESr7dDccHXNZQVZC
jhEhrxIoPqe1BXlOp57a1EmgyqTST9EJj6AXoaMn1Scauqg0e++io427rXjY
HRML/+/e0tt0RCw/rA+uUuNo9jepXXawuy4kmDySI3nLUBBvRJfM1jvz15CY
Tjp0JbloE24fMXxbQNsSxQUOsCK6Qr6SspgTkt/83v+KzF/Hg9UFl65aB0ex
t0JuCa7opYzglEy0PzqSDy9jmEg35H1zP/ni1VeNsDkxNo5T+Lnkww9VuVQs
xOumgboKmvtAjTzuSA26Wj9xRdpuR8sd91SUP86iXmsR/y0WYouEX8kpqvPp
dtapdel5MJ+60bLDZBaLz5/T6S3QQIVZgtnnJ5gZYHwKUd3ary1RSYS1jN8b
sNODdk9FjI6Vm2vpGCUp+9S2s57QXAIMv2y245LLMeu87EkmkmTky37mIxMb
29GX+f7EPksC0loi77GNIRP0xg+673DCmbflBulJWybGJASfygqXtVQ64tNN
OVth37bu+gueZ3e36/MYpm+mReULoz6IwSai48zqfXIsaOsBp0OORCqedydV
Zdq9cOz37LzaqvU0hQK2bt+McpgKxWlZaB3sCiDVlb9oFZazrQ/EcmQ+a/+W
t9Yx4NK6jpUfScrPVVFtuCODWetEv/R1PLRd92C+DO8pdz3/INzrlm8skJHo
KVb60B6FiklNZDRQmrBhzSFR6QMMTRToXGltN8dBHgl/d/w3Ch4vb9R7ctCv
CIAOgOXY7LGXNzAmn+xxT9fwKPy4DjSS47tp6nbPyd0FD/WG95mybhQBHT7m
xG96KBqlD3LF4RhB+elh3y4htpFLZUiK6Qh1rnIWQEuQPMbxccHay/58Yoa8
PuSLScc7zxNYg8CgmK8xUJwPCcN/Yn/ckcjl3dZNMheUfsFkg42iyAMDNVg6
lI+vnIs08XIWso2vRlF2zcsNSOxnxKPDEIpsNawBLAT8JEUrwy2+OYAIThcd
LxDxMWK4VFU/GBkSSQaee9tegpE51qKJlb4YIae3X0irWKNKArKwB3zNuN2K
U+h5NLASIUzUZrHmWy1x30wGnyFpU5aNDcE4G3VlPOxXxlvDdXXJaFPYxN2v
w4fZHdyNXx3xF4xtqPjuYKHp+orkuTWo2Vo4ZPKISG7j+Bxe+x1/aG8JCMcw
iEgPTVh3IZ5r3bATqRD2MR5dYtgRAlqmbom3NBs/yjl4ga2b/OoDj5vEv28m
tX5lv7kfI70SD/2sXMUwLkdN9qGm+fBxjcgmyXZGoI3BuXnpH2sJlNzQwwMR
X/fxV5uPRJlTWl+cR0WT+Oin1IVsmYGB8DXG9GZBPdgJfkkSIoJuKROWjTGQ
a6oNC5XUkoscGoGoqObYavbe9fzCO1U9ZYtUV7x7tCMZbJD3DNMB4oq04t8o
X/vUIAn8yHc/YUiJt7BOJI4MZGpm3NKO7p3Ai7Dm6gxQHA4siOurHCaYsc1d
EU7nkAdqjUADAyUTJ3j3p9LxgPAqpvYT7RYDVaZYh83k8RlX54ysV23TBxh+
mLgpf7zk5LVoXH7YZw39hWhvmqG7kcRpi6hK2J8CHmavouBq1pLYBkHCnT42
DvkkbqDJH1sA3Ss2boZQBXU0mEjHlPU9gpPiFvMVV4x3I8dXrYEKmRf88WEy
oxnoKoxWYTLlwXdatjB2by8WugqF+E1BS8GzqJf5S3aWBqzuwmyDes8cI2OH
wgvo85HPOn0u+eX1nhk8dI24YxDHgljw4Y4bk2yw7vzJNLkeReqJxeDImdfo
kwE3mS9E3O1nnKvPzuNDqM3a6kmE0FhSIPdyYVoICsJuGU9e7Ro8nqhaMY8W
m5GeT+NtqJ2XuKTpFqKkS9coh0h6+yTUyCdF9UkRQF3gyNtaO+udIREaamTR
/n2LfqC/lO4jRIEhNQ5Jk0V9lSZnBnJ2nLBWAUPlWjUnJ+J6NvGiMg57CLJZ
80hHzNVo1thsnPAEXAZYuDP3EbZEzBtCIJcsGkxpsVuQV4BSEDBab+M4Q2yv
UtF+oYCOX2ZHb4hdmOBGhj41anzKpM5UmGQ46MxYcmxnWrjd97ITJb5W0Fme
2Y8NE1++W8W2VOS/Mh7ZWKMOe1YlkzsM4EQ1SWEQwVYPvGdgWTGLfkj+WA9w
kHgdMBl6z9MHlsVvPTJU81GX7x/wcWKH9xIPaJQjAJRqFlEZuWbd8C2WXqwW
MkIYaUaNFxCDbHzBlCbZ+rScr5kSysQql1EIOz13+WW3zsdmUNg2WRSPdBCk
wLQtzPfWvH9tXynUe9PZHFMvaJyvYZFxPY7GmtDhU9WtL7nJ0Nhl2yYO+uf+
Xb7GdKwaZDEmD+5oireM8QE1aNbIryJicOoNVeotssBg+R2P69uzxwDB0HcA
1NxT2spLPK2nwuIqJ7lgVPw3CsPExPx7TwEGUKvMevn8ffqBmRZgyQRjt+Sp
ntMKVFNYmVnIBUL12qE+F9VLu0WNHR4C/8cAJKsAKaNny+A2idvgHsUmUCUq
FPklLMjSx2r+MDvYxoab3pFKVij62Mmtm5RS28yf5+vdtrrFZxf3fSrYhE7o
rUCdDuon6+BIz8hawPZdCbQ9q72REpbr889HXEiD78pTfSJWvN2/A8RjAjPM
HYbRkyUXHcJWmcLWgDvbbU/YepIS8ZG/cqAlO+mqxSSC1/LQDWX2A0XtQ9Ov
WXQeMLcDacTEzzCX0yhhKcDBZayAog74mtwv3s1fP0+zHPCHi444NZr/UJhM
XEl0XGvFCWE0trPawUOmjHQil46PIQFSJT3JPr6WFbEZE/a6IE83ZltuWQa9
uJempcZoDFvKavRoqgvEjN08I7adkUu7orGkOSSKaYkW5axlYym/oPkBUZYd
dTNDl9qWbI0f8BgrM5sjt6slinWCXr7FJT0nxQx9oPtbXBi+MsmWvXir7vO3
2WBBMOwtDTqtzHUtJim01fmO1ROFQnkht9dTsgSQb7cAGbmr53NMynrTgKNj
83KSREWrhKHPX3DjpFwhQJnZZuknDAc4X56FUItpzWSOdHIPPWlHcWQBzCiu
BnCfPDz2r+PUjOH1IUzq49EGu6ojJoV4BaK9isXd1eWNGOY+xKMOfyuPGax9
Odg21VEqjHJzflpr0JGMImSfjfKLnF6WD5GFs58OeoKRIZ2d+U5hqoCsAjPn
pT76GnAORVyVPebaC7rQMI798VQn3EWuUrmsNZ7dvTZymaTGEmfy4YakFQL9
zxyPNVe3N09tR4dvUFQ7i0OERhhUpsm28x1H7+mVpyBT489h8ih2k+spoBHl
TAZ3EmQAWk2Di0NJTg1meoGPbFcLEvu+lrd2FUdpLI1lYA5VKDMfEBsrw/jY
X1KFSU78BBb2ONTnzvXtxp+XMbWJwxg4ZFQ/QJlChCrnQddb3ubrOWSUZapO
FmqXLG3PIa8WN74J+/hfmc7xvK9ZqAViEK0PuMbXCg/MJ0r5uno8UVvgJnR1
ioihmfdH6FXhcihtRNXWDtUOGHGW7eWisp6kSso9PlpnEtp4g8TaT0E3GPJN
3f7ZHykkA17bawsFuTU58CRk8Ny77tQALtsBIK3K+ZFcPcpxAJroYTuJ/pOT
ufnluSRgrlTaLjPhFWYKEkBGV/2PZpNHF/F6CtD3L+UAK0d6iogb2gIxD8ee
WQNCzGcsrakdA5AjK3PdMii/cvZPb7nSOwNOncbily8EpDsorle5wJ/hwI4K
+KYAriU5hk/c2WYqvfpKXnNdLRjBKeAD0Tm2qQrkGEphnAj6ShamQD3LMk/H
J3KEtzqwDN+A0rGowjPuqDsp9bBJ3wjS7IPnGmDGAhSwvZdffzDO66aZt4DE
7xE+ZseWfwHTZZsrKODne85iWmZqOA56KFojxD9+oSOyW3PFWtTrW4dQWW75
fkfwdvQtpsPsTupxIzJUnjbP0WCxhVgW/fFv1De+VuP9gmzQFXLM22KNsVgX
lyHdWD2o47ldTWzMIvp6jjZVL6LE/2D1roORTis4jMjUTQ6byzY2RWJ3KFnl
+pz4N5sbFqJ1JKnOys3ELB75hhckim9AXI2YmkyVXdASWSUmzUbceluQdWT2
lyjqcs6yHKULenXSmss/P5m2xbgb8yppdiIUs6TMkxHt8MOMth3HupLcQygH
aOqUCIZ+frZua7H+2jfyz3N/Kqor3RpJuvLZAK3tCIsN50cfnkFws5AlpY7Z
89Nr7jo8GsHICRv4tVJ8xarvkkDnW1i4lEBhlZmZFJpLwFUH6mifpDJNmpxm
jj6bsxkNd6CAFGsTbOxP6lyJgAwpJ+I/VGYuWCi+REek5T/+Kav+h796iP8l
n1NRHSCxzIf+xSEJogwCPQ8XAtprU/4d3LAs/QRyB3ZLZGNQ+bzdveBnuyaO
YGYz+dfWxW6eA51JGwdyYbkIKICx0phpaSUah9VimyInwgCvAWn83DKEXgp7
YhaSgLuERnliqFmOFBZxBAWYynfulk2BGbPLsJY05a2nfxg14yL8WLTXHS8R
WgFtvn3A7xB2/5O14Pw8g/dwV654GzSr+TNwVJb/DGu4Lsjsca3BVp3jt/Cf
Vij6ge3RoS7gZkSgCVu0ebhY9KgAZ/4wEHWx1pZxg9PMN/PyYDp1BXaFjoF2
JIGT2iWpjwd2AHUzjvReyQ+pSZqSxlzVuyEobXPdutlZKVsKBVuPCZ5C2OVZ
EudMGgIqo1HY5sEmzjJkAve8hessCHv8609kE7G1WOEomFYgy1PTqKGXzxLX
agVhKw+XWBxWMZkdrp4DIxFGoIOVjYL358OjrfWo29seBUJ+1tN15CDJHO8/
lm6RZXBhh8lZxq3joy2/IybKTCsrUsJsFBM7dtzrvmLzSszh/O68H0alDKpx
FJXkYkH8VtHoX86ZhsoMAhJ7SgXVrA1GrsYLWzVlnsrlLrbUwhiEriI7I8Zb
sJt6In91SeFPDDhGHbIWlOvJ21Wb8eGk1iyVUtnZ8zpyyYxBUxKC6oMsh+uu
cLzzuCE3SqSUKxk5LegQZ6MebSzFkoflBHFE8hId7UjaqfQIA5DEmKRmjJpw
I0t3iQpKlKHUDGtS+4ZBwEtOGAwxks/CTZkkwzuERiO8tOYq4z03pXjD27yC
ieXPtAwx8Xp7lpJQP9IP0P5nuqpjltbgZK6e5IakvTj1WPqjL9gAaMoY3OJo
6EU0P70OxyLlgIhbm0yP03Ir7QLAtY5AQs3lP4ZDleMECdPwlCwxlk16T9+e
m3qG5Rth5sPCZXIJfhnH5wj2u9l69jTY8Kc4q7v0rmMe5Bl2Yzn6JmiSi+fX
PXxAdTJSpW+4rzROBklTM1UQG5AfaH21AsIQJyHoIC1Q9AJ/ziKyUviq7T7g
jW3zruCMNPGln969zwUOf/3Pbj2zg/dx/dGQrNlEAzH6NUsEZbxLTjf8ZUxN
R1QGkSStfUfPfHdUzMXMhVcnw/sT87i0Y+vvLEg6NAQAzv6La6d56ZvfAoIK
zlR7GD7Q+gbZlW2TTG+LuBGPN7def8FlLZdTYB4AH/0qYUooYC0O+iPA2k0/
zaoYq5UjOyC/J12eQcEGAanGy8Uj3udV/nU7QKzQKk0kNaQkjWpCpozuuqQu
bdOhRcAyypklXLU29Ij9pxCI7N8uu9yrBpbfKfoByh7Dee/qmhGTk4YlMrRv
1p2gMTODCLxKEk7MJrG8cGX2RcMfU5EBpAO5EJpKJH366sLDwV2pZKY22fCQ
TAlOXQSir/OUo4Aa3IOL9ffDlSvK6/XwzSgw2Cj5Eq03vGXdEN5t2QIb+B3I
hbbCY3u3dh0PGpKgoo+1D2N6O5TZJ8cZafZ9amTK5WQcalWvE+SIGh5gCaAn
kOp4DQAWdtLSk8BJE+IXUiw3/ug8FN/ohRBHTUTFMXH8offEh/pq9ZvBeqGR
aiLBDGVJ4hrBA4GkMwwPotbikA6MBtm4cRYwGFHI4afLtf03hhu74izT7l/+
vFUuyU6td8zhNb6jR05nUR25xx7jfJjeNTWKMdEJ82OAx0D/ChQ9yh+RId33
REszX7FSE0JHT9sMeQw2qPb/2W3rA/BswEVze7yT91gE8TZpQ3D3jURrxUl/
KV3PQ/vC1zrx+3XyumcdnqezyyZSxg+qyeiO0h7CQ2YPUbMVqhh2zH+Sp1zX
xSBhMFK2XjG4k014ReulNZh73fUK5vfTJBh02wR0YVT5kAfJxQ/eFuFflmy1
QfkZEeE38oiqy6r5gCuiKH6MRTGMo+MXUuzw8VqCcSsLAt9LDCUCF9DlLeQJ
gZJprnYsXjDBjYodlfUEL1t4G4xLRylhXACJoR59U290kCrRJ8jmgbG9SYjP
ZSLot50BxYs5Pwb7C2fCfCZ9twB2CrUgEXKxMs7mUoshiKGnqbn4VNjBK7+1
8Bl5bdD/qAo8BCyCDtSCWtd0xT14ZXgzghr71ZT6xCTtj9BzomqbOVrTle6A
aRawfU2aYss4wcrvhrVDpHQtvtfZUKJIUAjpBSS/xcZzyPElnLL/YOW/SMeB
v8nXBWQE6JfeUdO/1RNrqxAv/vEAjuVcjo76Hb5AjZAbbAwIqUdytcoVN/Vz
DWMhjAxZVNZIm4LFxVjJJipoj/6ZWutJ5atWY+mJXgRNzcz/ZfO5m7JwilIK
3fhZTKKpb7jm4Fu8axaUHoFuAagGcFjrYqvcBxEEz4wwrTCB2DfEhTTLl6+p
0QZSwf+8xY4a0lq7zK/M2SOsLxtTWR9K+bL6LkLcaOOUAbv5xGnkWmS0VcsP
9toubL/EcrIrmHQYjXooqmLjph9GQVz4jZby6GXwN6jz6hLUAzjIUDRg2YvE
gQxDsso8IoalG4HhwR3nazi2k1rV17wgr1KifQmFK90EuJl6INDFMczj3wd+
HfaY81bSN2JqKP+AV+GMUXp9hPH3sc+LTzGDg/W01/zvqGRtznK7Sh7JdYA/
R7330cAyhF1a3GoLhxhHn1W9p3IIST+SiLEBTl3q4dSfTZmzKG4QtkVwB80d
4Fkz7IEom5TdQOuvthbtl/R4+KJIQLK1vulSGAHwGa/K7pGVwOtWIxCj5O8R
S+9Rj/+i2rjXQkDpmJefZGd2M6ISpHpPUUyY7Bvwu8I3s/kO3XGHWJrYknuS
Qfc0DJKvfB9CqzwVAlWLDjjpraxG711WFwIWFClcuzI+c2VLuCoUPSy2tUAb
FIa45KrjtqVfQ5q7XPXAHyAuBMPpEUCVrsKpTnzSHhbkYeVO0XjYw/gwJJ4I
sE4716CFM4yZzn26hIYK9fuCqI8sRIvO1Q35OJGUE77yeExd5CNlchQ+9G5V
PrAQyaa0BSOWPNDgangTOz6FIVKCBaLqztxwENLDgvV9zDvrNsSZP83MKYAK
JMhv4xBu3mjWPHXhTqBFzzs7ptP9uNut3O4N7sZyzz88HVOCQiZJ+lAF/OPh
MoPNbTCbtVG7jitEOVtbY9ht67KlhrvcmzHbTtWUnHshf5sKAHWfVPIysVAm
g9/58R68oHJPTA2aqzLf82lpyJMh8ijywiyErQ6HwdaiidSW6fdnuO+Q1P/S
HlkgsSaUyF30VPmg3WP17VhFAlOvdReQT76ULEgNk8bpZYToHpi51tgpUuLS
PMV1xMW3jKMHQzR7p1YTnCJE+6ca4yYDz+6oL6RRyBxHkW9q43oruw1QrWGr
OLAT1BAeUS1SjUxAZKpP/HVvTauwYFauuzyy4aQN1zun/p8ROyqe4dp7J4yL
MgGvppFXqIzOxX1c5g3JLDMJIW/HeOfAbBCIC5Vtxc1NY7uCXJi6bczTe9Nc
+skO+IyCWRcPFTWGIeAFR33z7572sIXcrz739iO03NjqiyYBKXPgpwu7GAiQ
Y4Y1a+Ek9EI4c4uXkYaxjyN29hLqEL+LxeSJcfrDxK4sMe7Rmss44MlmWPYR
1e8t+cMNmA/90gLK68pMj/yNG3pWJBdCbOEj5WZrXQfpYgjUzgaumw6OYI8z
LsJnpCVoU63dAjG0g4SSUzbEcIEQnK1fo2QeS38FFXhmzedt+9i0US+/4dOb
rXPgdtHmggxdHWMklmwtqcmUyYlfJlihhl8PmD5KSHFOCQdULdsFKmY+PPEw
zkXYq5ycn2h5V0tl2UA9sqpXHHcsrDw8HjOtIe+k4teeWus1JafVTcJsP7KA
vB7eYP/TXOG9wOH5e80GGbZaxEKjvhQjae3x60KG/Aj22P/T+NEsW2ze2NMy
sonEmshh+QGMA1vzcintHzT8Z9fn1Hcc8CA+n8Mr8FLzSakbVHHxTTKpN3Ql
qfHRQ211XWyCmLK0gItDfvtUytnU/GA/eoAkqjPVuimdhjlCPi4n/RUE6HDu
0ouq5m1v522eXR7RMRMmiTZkC5x59XZNXbom2imn+TTOG8J7uArQBhHBj9bm
2GAm4J0vvwVeLmqsK84tNjTEbdsj9KhTdzqpLTPllVknBBMCqP5wHAJ1xiBJ
/aF5nfzLm3XP/NXT0XMn5k8t7hMvyRGvjDX3WydCgbp0KexVdic7Y2hr7QF/
A7YKZgFWXRZRbW1NmD6pkVUxzecC25Tw6JviR8ttbTiZic5a5QOXsh6tU6HQ
ROjrgdpbivZT9s8pawIr2qA1cpRmYSaQMNwp8t45dfWB0Nl9jHvc1DK7X56P
ypl7Tqg2wh/gGqtfZldeb3pHQ9xUJYn+o1TSfAmTfVoWOVPqtY/GQHREm3lA
LExwVn7KbxPYxaJy8m+OUtGCFFB/LhbITSVjSRyUnEFVMcq0gYFGUpO4lmnK
EsS2fOFe95ROnU4SwYtAgPaw3SGI8oY5echzfAKZCXEyxwvoJehSWy/esfOE
OyXf94mOGjQsYaDPkTpiyHlHwWxFeJzSGKugcgN0n+PIU6DA2ARVvzAC0Oca
oHkwTQDO15O3n0gmvUX9LyDvJbVWSsAh/6OHaS4CpXb2MUwVy375LTJoyTb9
lkBJYK0mA8heNelK3ZIml7WvFlLE8BVpOcJSf5j3XTmq4tjcHbhQ5zDwla9h
RQkZmqakpBFUvcOdwQz051q/NmQaGnKBvlHAStxkWxq+yDC1rO1j4V+BFAUT
o7fVqB697rXD89+ynirfcVS/wi1C6K6MUUhXkYLfn44Div8UskWIX7ebZ0tO
b0byToxFSpRUF6vJyrpHVYjxhpSoGbYB+k8q5xBMvbIaurC1tIPXmtz5JKY1
po6JRhBdPP0lpUGyeOOA/z1geAsm+Go5kkkYjMO/fC5OdcnSYIyve/is3BuG
Tt76/mjNINzunzy29FrKonI0tYbQ9fk5Di8ETO3Jq+06YAIA+xS6mIquxU5o
oPmNU8WGSvdLSKIq2Nq1rz0BoeSgNJKWbu05DIOar8/o29zVoubozSYsavvo
Q51gdb5dyL5r/OsgG1nb/Qt7D5KL8fTPoDoluMghdCYvlaA0nV3HS59tKdnN
49KsKqjWBFpcxUs11Si92X1CJV+GwTq7Kkp6SfPEJJ5DNsfh+1HjAzalMXzF
EP4zTKCz7DdQct9yF8AfvaEpqTtFr4BCTnigkNbyWviMuuwoEzF+1OvsJPQn
vOO0Dn3zq15TiTlbbVFZpg8qn4YJqT0ethSdV4nbRYR20XnHzMdCAxyV6W1N
pOr4MLxbGCBkBsj47ozDV4b6sYeN/Yljsasr5PfWJfA7cJBW28KZdiQufhcB
pA6EiflfAePfReYabXC74h4jRVn6/87C8cZeIFt22wfU6vUbtqVwRD1ditIF
HxqYM8hQh+Bdny4CMK6SSxWfAXLGK+F5ZbfqZ3U0vh414/JXTfHl2uyMGaPg
vXs4Dp6JDCrGrRopQ/+bJRtRPDmZ98cu/IrgyM83EE2g6r+3g1F81tVC2XjK
olzt2Nq0DQBs9+ezz+q+aQU76bde15d7yFCCYKWywmagKQkfJczQZD8+UErl
zKTtirYEOs34WH/hBdFnaSKrgT6flpSlc1CNKDm6PSEa6DJaZfGPZWR5jvEB
7yAa8zRn56MOQvfIGDYGWdRFn3cbYIWX+0uHLeKct0gOY9GzoNP8KdP4xUd6
JCD3cn2cKzwc2uqGvtcAmf2BYbBnW5CA9ER1/IP9jvGClNQSbjNFqfHe9urT
Fb08xjSaKYg8izKAOwNrihK0lSe7bViLxP1xEUznLdwhx9+sctxX865G0UhL
XAzaqRp/csGPU5Og43WzXSSA2zvdRV6Z/12cO0kjaGAdOg0gDwDSIdf4V+1k
+X1gPQ+8YrClHsFM48xduULE5zm97q31ZqIR/aKinB/DjbO1r/Lrct9+Nk25
RpwLZmPAeLsDchyvFHcrUYAWDsI2Uum+TDYvsyQ1yJ4ChtE7ORWPM/pOI4Kp
cbBS42TmqOuaa5InjUdFCmpRiRx+dXHrAL73JRQXhBtcU3UojnQuHaV/JD64
UFFToXOrFBMmYvA6RJexvykdYhSW0Gvw/ndEBaQ3KZJfcX9olz3QBhftsk9u
oLJPrhRuDBZWiELqJIbBenQ32bMxtl04oVe2UIJlyI3ZHYTAK1CbdQofyPx+
ePbJAsE7p3MXwat8oYT96q1FCDGZXp5U6i+Dq/ZZYVblKYnDEzWia7PxSufU
O5RCIigHd/oQqiSxd14SwDJpjCNnyEi6I46E/2JfVHNPH22RKgdi6CmmcfvE
b1FmFDBx/wUSYxid1Sxx+JOhK4zTucthofCB49BvNYaAv8Pe0kFF1bDv+TQ9
kI0pNKu0hzM/weNQpirsarroF53P9p7FRS2uSOBNlSwe/XyLbMtCgggTg0lw
5TpRz20ZLaCYHNG7JtN1TTVNWWGKmricvbr2sfdLqE6uEz5BZ07ydRylRpzG
LpefN15aOQ0oYL/t0qMDhpqeC6UKocFXux/N0otyRNRbo/IzDw6Lyj6vnxbb
PwuO8M/yTXbPrhdsGYoHVjbYItko4dUTb58V7kYdqFH9uNPtFmlPRQsvHBSM
gFeqnrpSSYXDvPNMhEQ/l63fROm/tSeoZTNuMtpsuURbURoERS3mvgIWcw9I
BQDc7nHPknWogy0eYv0OiaA8ztR3bS+GuNBpHra6MTua5M2TedQnkErUBb0z
sNhJIrXzvfjP1vbPZ8kDzpIPinpqWnc+EM/PdupPkeEIGY3Qleqwxn/+UV42
j2Ik/FHISTqW7EWximC0V3QoW7oHrj5rMpDR3z3IfTb/++QZlZxWHoDJAPHx
3r4CSfHXgB2t5SN3Ue7KDSAGEHMwlknYU1V/tcK3pgGY+6hMtom0stDjOiRD
y0wWq0WuX4xSlHSMxWSTOU5anzVd+iy7ePr9486g+d8tM+zeri7O1D1p/c7h
T/3nw56iuDXfGZjwLsnr2nDFwwmDLorGtXIKNWQHofYV+CvQniCN1YTQAbf4
xn/0poblwZmhjws0HnvJip7M77ELV2RQTBcggMw8pA7bltEoPxOWnBCQKYbv
9pqTBoTcjo5zqQoun1Bp5h02+8xBx+hsPbYNqAJBfhBRQphS+YJObTTYtW7C
AMzOLLvJbQPgA1oPI2kvGmauD14Vv2DQUe5xJElHHLyqNraLHMReqb5teLqQ
v4Vp0sqHVVGT119xGFbPAOGX94G9Ar8a8Ja44rDiZdLpqXsdnlJgszvqGXHg
WUMXP3hOEA8WVAD2qmhdxwrtaD40TV0gBkLCa2FsUgrj67U+tEMrAgpLBJq7
VdvRMklrZu/8lHvOePfkw9/IH2+1Mj3CB6Q7XyAYozIKf7dtuuquYDCc0CsL
f+Sl5DGBAj02h6KTNMDo9R8J7CZNUSbt/LaYwkaW4J9lEPMXgo214RlLZs7L
TWUQIwMgs1oLNto2dVrbAL8nX8TSkKywvN3eFQFcOYm+OyKizsVYOD7vCxMM
thHvSrrFT2pE6PmBhyhN+QnY39faY15wbCn6Y+H+vJcnuuL6/E25Tz6+QtSc
T2WZ9bsv/XAbFO+3hkWYAcn0WDzD02YrnWOnJKPOx94CmTIIME38mrrxaPiT
ozwJz2Z7qYqlX+kFFYOt0rPv1lK3ow6d4u+gYiHdC5ouZiDVPJfqJR1kf/O6
/cNWL3xWpcNuNCQduMuuJuRbu4mdipQRluhYnPCK6oEHue0lNwt7oW5HPI5W
2Kf0voUGz5FTP54Q8ZZt7cZuMCDmvpAQnPX6omoTBCmp+8vcj4bu9lw8Ltah
E7cfIHgZRw3eS0lhvBcz6k8qQYQDwJR8NvD6osy9dGa1hpG9gtwrw0w4DgUs
yk8QZSnqR1uuEcnUNPdJmwVH67tdicWWUAbORph52fH9DOAf8r/GzMLOTe32
qmxJFI47RV794qdZga+W+86zkAAkl3DdaGWFicDIn4yg+UN7Kqu3Eg81ZqyR
LIqTXAhUgf0GcJ0FH1WAEr1Imop1Htwr5x+rPCqJjFzjGRnbH8A5koJbrENb
WM1VCbXMZzByOYzZG/KOoLV+F1aEl7+ZbbDgvH5rVkGmp65Y8H7FrfUhcY1K
VntzvXk76lQj9GqU+dtr1y+WfL6w3KKcwX214FQvABjifnEX6jbcXilmfNXw
gVl4hFd48NHy9iunWIAsvcw2wZiMh4jE++XSVtIBo8TG0t7diLDhUSt0BDe2
vZrW3C6CywMHdez7RtgpSchSg62F/H7yyE3LUeJO0n6NQKMD+lRlCfRW+xtT
vIS8kSEwYSyUBrqUfbovxEKG02mcPx2J5qCGbDMW0Xc3iIAJZIEKaTTjRDMM
qmoFQ0mCX5VqlXnQ2QBS+8vvq0drDHvprZzyUCMl4wAnDCcw1kUfJZ6GPfX+
45XVeZHkJwiKOfcaflbzY745/5yZguFDqSgWR1SvfM354DU7POmgNPxv8wDj
UV+lSB0Wg+w6tGu4FGNIaseW8T8fqCdRm0yk9b8Igf3faj6fT5kIhrnv/dRV
zwqapGQeQ7TTRIHecxt1sWFYDrdcdioVcjEzreu6GkvDWVFsfgfKmUzIkDdS
SekI5bCsWwdlt07NB2hEKKLJ6Y/h3LbHUpBj4d3QWAJEkwVNKnv1E6Ya5Roi
naJs7TJGHVqLcfvLMzDphjiX58uPBBBsyvgK1elKPnRuET933Bs6eSjuc7iB
47ST+OVrUWZTv4iBLTi9sO3EkZ5KrDiKyhdIMaH3CvghaMiMI1xJUvy+XI4w
MLt60HVoIaERSIgDtFBS3bLltSitzGlA3IJeqfUz6e0qlmoBsbHI414DlPNr
iAM91FkGePMbeLtkR/Gq3WXQB1JOpJeoVULjdpo2mBoG/XcwHBXCe33eqhaN
KMshpavpIfu0/iua+/Pucg62K6Yp/U3jlmpoPUAz0sdpfLQmHDUvJhnif4i1
3LiGTvi0qquNuS45RKR9eaQt4BBRYB8bTV7XP3O/D7WgsJifHp0RROgqazlQ
LeiKVYjmD3/sHeYK0bhPV3K/3NchwNyf8YTbNoj5nNx0/YiZEuovCjqkMBDM
LGTQ06s4S21LEFeOj4QY8key7xlO8PjebUydblHPO7MVZq7krwlFT5vXpLd0
hmBg9mDjnuPb0cfJjIg/nj/TEyLCzWsZ74RnerIPYVhS3Sn+CkGxNAW/Lh+U
kE3b685SOJNItfio1MakuRQ7AidOm0CipSIuyCrhAqbrF6rkcf3xc/4nj7tA
uvuQUbQ0VPZnDwD3kRzUNOIDtQTWS8e5msbRq5aOLUTeNuJpHoXDTRZtJlzJ
nItt353OgAW+h7xrukUVOS/uv7VglIdK8EGD/2zfG99gxwt5RDKqbK26BbA8
N9nCtX+Iqc/LKYcwtXQJzrvGswhS1IPupp/LIyAKJ/w/FL/TkoGRC+mpfp3d
dwKwfEVlcPPE6wvz3RybCqWokCHV/5vvdvHe15d05063txdhKP8Uyrl4lHpS
6f5m5XUe6M4wBgCtegVn4z/5DsJ0Ra/oeiUzf1zQXwLVZoLVzc4dWtTDpgha
o0S8P8m651yIaMc6JfqAHkOVrz04Q32KZ8/HdFXIXlRonZbmuPhEGRdDhNNZ
+KC3hYSRH9ww89C6HZTZJ7XjirEKOKonz2pqY7TuZcJ1TQpu0WBhY5WnC5nY
xbtdnC8ogEavkF3Sk0Hk9C86A1lF4RkDlVDup38s1MmR1RG8mYt51nP6SvDl
6JiekexCNwfV0azTDn9Lg3O8/Rzjro/4ErsDBsh6dX8czBdowEWNQVBjP2Yt
pXb3mDhrozmp2EKRertRwrqt7fIvLtXdGO48mJhJSz00jUGLrDKeTnW1qpl2
APDr86Uy4xkkhz5E7R9J3W68RqFlDWiXzL60+oabctRbd0oLWelhSjSZQg2o
4P/XC7rrT5K3ze1AV3VtqpNq+irswksu9NUu8dwSV2noL1Sd5lvGN92lKPmV
JRSYnEZYcFIfn2ELXBaS9GG/35wzy2ePAd0CrrBP5s+QXJU5Jo6bR/268r5k
GEiuA2K0jz9JOQtFZy1EZsKpxA34FFmLWBgGQTZ4nMR8QABsJvWT4CYUvWY7
H5MkEJ2N4Xrh2B/+7y0LiakGvehpkPUQ37BiDH4m0p0Tij9CcXzw0ObZ/aaJ
a/yRA059AJuC5h3m49umEGDDq57xFnCEI9VaVPmSmphAo0StmYWLdroub4Cf
YJ29+QgoCc+gGtXf3gVajC2yCHqNB0XSebW2NCY0mvWN8es3Sc3615+JTg5Q
0GjHXwEKgQGhpLB3v1tmtw+oMdJjlcSa/4OJNvLxUux8VYiLCCKI8wtZndt+
//CJVlEYo4cGxia9FRutM0UdIIRkgPXGb4/MohxXWZFAAdd+1UHdkLreMdaI
J1AyAbOXEevZBdAwPzFyyzBCiqM1qgf9NWB2F4Zdg6zPJ8VBkUHK215zeEmb
WBpeK7MBLD7RBWBlyN9hJ3XxSAJgm8hv/g96T/3fn2v3qhgwI7jb7UhCoGPI
vKqQ+pes+63x9dv3C3FhfWl6LySPGO3xefgRN0InY1WAUc3D5C8KYP49yaSJ
XB2Zh76rY3qRfvsmgZTbfDlazwRavWRY9tFmIQz+YQVQJKIl4oh6EsY6MuJZ
eFJyrSXcTPFD7aUHjMB5UKhfRPUavXiLD3bnL2ZXDIwHU8+0Vp+uwRywJ/7V
h264qXHQrufZVr25+ivLEu4OalOSWzR5Wfpl/IpXfu8fyJh+TKRfvRbamYhW
Q4nz8y+6JDdzl6HqIlR1KqY0LqDPbMn7c+TiAZH3AZbnOUUFQSermS6exi9/
KMvfXkp7Bz2uCvO0isMkeMQO5jhPO+2gsuvC3MTNj3m3BjuZde8n6ES/WME2
vACPH5ZrACD8ZI+9uBd/Pak6wWKKOreG+xZtKjRr+MHE8lQpfuG1IS0XZRIm
/5k0rU703uB0p2JecZyb3Czgy8zy36pWdXVcsDXSsNidx/rd416hMwmAeydB
Xihvz+vF/F5uDzCiU5ewMyiEjD+eQwJDZCCVht/wKJ6CwqvRD0+6iIw7MG5/
I8debu8oAuWH2hhdvY8xVlI2g6sPdhyT3aEIEreOVfLlnkh361T3itVO5EES
CqFI6qib6RVdAk2p2H6wXtkluLtJkFA3ForjT26Z3yA02dNCSpTHfMVl3cph
yc4zymYEXGNOVZQAnji9940r+kceqafNTgBqmARPMncO6M1jwM84YBNDTTjU
TkpvNKgrwffa6jyJrHlQ6CW5npWPGduXy9a4CfbOgJz7r80qrmAwXQL2uFTI
YAZF8TayTLoY1nBj30RpOdKUOWaIX+RFvSCTLpoMUZuJvHRx0Hu32jIACH5T
jOIqaRuAr7hw+OVqC4C9d09d5SRR/FHw3hnlf5BFwFjFgU0O60fL6NcOzzQp
DkGMBjGh9mXiQRXpaf1+UiIEuWha8wF2ENrtbrHM7dyY2XeDm9v0ZYN2YAed
XQp7ndxHzt+X0B/89HfUAuYijjQNcicQRqVOo7A6xit46ZdjKIX4HXytp+Q5
cVGkTVQkURjr6kMFjIaBwjteu1ApZ+eJjsNtdZJ8vCQ0Jbs6Fx2bfeaIcgBF
FsKWW+xE1+3lf+5T14HvpwIUGRRPUd1PPLDjcshZ/vDMdmWV4Q8NAu/aBE1r
P8mII4EsbFBwLVKIaw8dAQAYeJ4Yhl9rDuPAdh0YX4/vNP7F8AEng0AIuCwz
+AeVuCoVT+FzKsdrb3bbKUWjn4YS4/rhFLXnSZ0k9M1hOsRqNXobFRkZlyWC
uHyx1AZb/NwUd9+gdtcgmPIOHOL/QM0jkJk/Cq4Y/jZRc4Awu3iv9H1V//M3
9pnfHzfbd+aiWRIDBObGVRuirImdwbqJSxcPMM94YJboePJh57sn4HdPPck3
yyVMbzx9iDXwbiwbvebBtKdiBVVc4fJJQIpEoAg6XcePqLsiDv1oIEGHun7x
tW7GLms/d5TN7MqzRQEoTg2KO4KIxeSqtYfV6Vt+0kuHwB9xTCdLaHVQNz9Y
OYA2zsN3M3KWmoMlpqA1C1lQU+lS93hwy6/KYdcltJXQfo/7Bz0mr7So1c5o
zxCdCVSqG04uR/7sC9+/mkB3BVIe4H09n8+SEFNsjF4oRZM6q02caVRcXpV3
sQS2IfZQnkogh8wu/hIc95tO8W3TVu5GbcPQeVJHlhNBeqd+TqZgvmMHOhia
lsNzTjoNtuzSTzjw8/GfiUO4F7jjZbaTrG3SswI9S8c0uJyu3XoFtia+AdF0
MmCFMFKpO47AN/4Q4UKywb1ZDdMYz14jBK91JDvcax0kGpFOc+NRRV6szNXp
NDIET19oYCYp+4iB3Dgj1F9qpTCwnQ8y7BmYrbBHqwU71HolfyzRsjpeg/bu
lvgE1Ow5YsUefKfgAmrobCtKp+yVxLbwve8LLICsMx/16JxVVwrruV5JzhW+
IHsQj0pjkh5lWlZZjGOJsM0fZPXvQcwI0LFKVEamAeAzJtbnViNVehyBVfNc
ZIBIIT66Cs7jzqXkeYuJuXnK928NLPB+ib4VMI8/z2MmmaNibtt+yh5GD9xc
ivK2vO+a4hRANXLqw2LoUV4I6Ur3K9cV/bAM5i5kROo06Kmv5dbFMPekaXTU
ULvk9eflr+X0IF2rfTVQo3tthOdTH5gAdC+K0n8sothf+o0X+PeXhj2LHMfd
SYoH0//8GFVrwHP2wKKj5XZyrzfQsNzbDVGjUmuP5+3hOcQg6f538+iG5S4k
1jd0f97gurPSD0p8dmEiRalu5gfqyKg3ZwN270xBFcbfGwr/YuDOAbi42vwO
MLGkbY/ZkwkZqkAr9TVkIhi3Col1Ehe7sEliFEgemldpMMu61vpnFIpeiJvc
M7deJR92n2h57ENkK25hC2yoEkjBmq+UlDHa9rCOh1MuPBe4dgAWbIfNX8Z4
G+/O7j2T2blUW9QhpjDFn1qJbwtZStGUkgQnVSj4STxAEyF//qrHTdwIHg2g
LePq6XXOAYrcMzdFYU6EN83AtmGOcxDuVN7+COoajYW9RCyQ/LV/tOOlDA2h
wgLaCNYPUrHYgfUrATi881FAUwJpbx4fuJPbNZgIr0ltKpMpbnXRVYSLmlVN
TnAP2nnA0G+xOC1CaJ+8c1Be1eHntOoZ/VYzLdsHKv6H50bPgVxmHMVPQPKa
RGrvWPW22TqRaXfv+mP9pCJYqZGTxVYefro9iDxYs6gqXEFERC5CLd31En55
wYmsX1AshrOcDjLsfYbkDXhKhXoxbA5JtyYCovnX7S4yOLtEME8NMnueGhdd
DF8io4lhAQ6h8zV28CyFMlPaZrgma+mJ20G42ESapCZs0DVMaCRROCRswF+R
MrFSOqq4upDQ1FzSy/81YNRsM3R3sOOJ6BJa8BWfRcG3wF/6z8w3ABZ9tPCN
+ii8rN+c8Oa84kusACLRgC5V6YnzrQMGJu28N/xCktDLwIGdF1ejZhXiwmod
WbEgXHPZZQco3AGqOf3b9KX5abUpJsCYMNS050ZBI9DsNEaoe0XVBlKXwaS4
jRvPOf1PDS1SjnCrllS1/Ax8DhF5ekYyjTcVA7DFtRsXIvXXwGsn6wLNtvo8
+QHNs/czcA3KwnY6c6J67bPHIm9TT/7Ia3UT8fWx2J9uOTsVEkTqsbNL1R/u
8rSCmGh+pLpzI1ktpGeqxre3i0rUaivT/pov7Q7kYQGNK7/6iuz7R7B/GVeR
ZZoZL9njsSuFaaTZj0IivY6jA/dt8eV3cvzMVBcK+9e96lyMV2sOQrLa577L
sDjoEG6enpybQt80TCt7gcEWJ4OqIDMszz9rMcL7rCmRpn2odPt1ivFio6//
SdrPhrrvND/vrPHgnAsPnf5bqr0B7UOepjHn/gyj0EJCUIphPNPsHRT7Y25x
kaxqNCLehlJVPNyBXtitkK2K/dIqIu5jtQsNG6On2lmoKDR2NVIsyKsuFAug
yYjF+8zMhlJJNtYnx9/m0EAOSZLmIdPsFZwbD4bx8PBf3kjJnF6OyFgj9lEf
WIUFge6mqjDrpTycWrqG2z99YNSYUoPa/xrYatIzrA7RBJJdD+oJAA2MLQxe
5ha4g2mtIrbIPODRF/yB3ytvSenKdZoNcW+RHN3had62OvtldBz1UemjBm7H
T00v+bVLG22U1Pw3bsqz/yZY/yZcdN1gbdrsrnLdM9OHku0jSf/R6B7JrARe
uouo7/jB9TSshwQq9ZEcQreU/KPxlsAcvzy8rGXsvbqqjs5J4t9ARlj1N0Xk
Kaz6oxVr+LejTLZaTgRlzLQuJUNQOqAgZSwmzc41j1kDXn6P4nae/BKFLsSt
cLfjmEhlFyk+7Ens/0X3WOklgaJcMXodoibpOE1Q+0LT+wQjiXkyxLnMBcTg
TQWrcOW0WDszlfO5gpH8GarfuAgcz8TStUDVbRBsLopoevO66wjgVYK7FrM2
cA/6CFdfT9rvJdvPHYzhN5pZ7rWaxBrPggQTC39ONuM/jrwSdeispP3/+4qh
LT8DElVX3PferIWGkw3osAEsMiaBlDZhEHrrQfO2GWqfwpunnCYcVgTrrMHc
+qN1HdzhCprXgCKBU6GX5kWd1TK3IlrSRb0pXDacekGtaCIC0D0ScVtoGJNK
pTmiZ64+QVILMq9fXmXe2ECH1wJCG8uH5QRGuH37jMjgUSz8LGv9NPfTY0Fx
NKLh2hzQrb7jNnbjD68iJDBVvXHTXr6OR+GNDWnsA59oXGjMOxWp9eQ16yqN
eqq77ecPcJNMdCKiNBDLi1cHv3SAsL59gWWoo/UDupdZUtvmOVysQVWPcBow
61K3ce2n6KcmjrrdsOBdRZlBjCzJyFzURPgaFvU60RSixJZ5UNC9tXB/9tT/
0QHW9SupNktp0j42TR2/fnRtMfVx+0Hsx/9jFbI7XVZ/r+X8i5XDNLrCTet4
sOoUlIC6h42BaFx4nYzYQpQZqvBGS8TOinC6gj9euvdA9bR3Qeqvn4WUADR0
7gpbNmc2UdeHgcLFuaaievxYPoppFBNEOtbJwZJIdU/W/0AMsNWiJ8mN6x1H
JjvaQ4Io9XBns5J9YHCZyjuIPsvI20xzI1BFJx0wXh4/IYklbMstG/q/9pw6
xSbVTIWUqbzYbRi071RTmJK8W79yVbmIBrBrMCR4PqeoJN0dsUyFr+5YK9V2
ed1f6SYj2F77xpcky1RjqkmV+/Zv1mwq92478tGonr0L7Md98XXJ3xMIlaES
fh3Mf+iMStebIA7exU41WoBj2gKnNGKqRS6J01jRJhbOr40L/FToAR3qV5Sj
sOa5VFwM0X6t1EedW2aAj0k/ShXlwMqw2wCSLIs2nxfoMZJyLgIQdZNxlq03
FrrpWYzIZ11xjMLZkPC1qBYps7LEsPdRvaMkgAlgtyN2WdTEzM5sN8yUn8II
/gpP2glXwaPqg5uGT2BloQu2F8iBEHhq4wyltTyrYfvkABopRRZcKPjzl1T/
7QcZ+RQPzr0uLWAcwTLmRQgb6bUhaWjh4Vhx0k4YGfqqTS+gv0P0IttJPPGR
/G4YkYHrp/v70IGvLVBEDIWZ6a/CqF4uNYruIYdsg4p7zNBXdKEQAaYGqjis
/d95oclBTTbJDvD/t1tD03M/VuloC+NQpD+33L2djaTOdbBU8bVkxKQcR73e
KmUrdn3sdSkHigOQMK7ben5hUscyOl9sDorWLhU4oHBK0pmB6/gvTBMfo9wx
MEMflwWTTwHiUfuQ5vRFfgnmuKGWp+0H/M4Wa0FH8p5P7NOxwY+WqTegJ/wb
p8ZzGvXAnHSYYtasBTEBF92g4mHMUJSaTYp3k3Ca0Tc3A5WNOrsHykfbgz+w
5X/YVywrhxz1i0SCW24QNx747aS5CwoAPHp6+QyTJ455Vugj0vyVicot+huq
MTIT1vOCxTeRr/zVs9rUp4+uSispSyWg4JBGOHYSlHLV++EFKuGWsSOphgCr
WHWR6+jG6fb7g2KxtdgyMypSXES0mmWCX7WZb3ICmSzdquwAe3YwwBy4Dnbm
ySMT+2aojD6ka7Gz59EnLFfieUoGLckLuFIwe0vBj8YQIBDF1lz2PG9MDAcO
myVM/YjERTs9axaiL7n/xNR/bXU4ILtei3hpBieXDuWMpLztvpe9YuPEiD7x
t30A+RZaI80VTMVyrnKkt+a1XPF2pJ9zIORpZKCv0VhXF+T7VWXLhcQgA56U
MbED19dxiCQf0euYxYYue2YAL+PsQQKi+KyZdkkgu7Qeu6E4UOGI39gY9NXG
pl/lmr/fjhYduxA1msg12xJ2Voe89mZwl0ArSwFCUttawK4SwxQNuknfEXsW
7ZqaFuZMwoU2dW+wsZRsrJZPWS5lne9m1hOSgz4unJ9tWezDtvwCVcsf2v+s
VyZHqadaK14QJpl1TjNmzxuYy1BMWUoWUFaABhIqADdntg3DbcCkRHV04jrQ
H1qnDZ3nV4QGLDrk6+hyj4DSVn9QrPm3x2GC84PgsBLZtkNhGiTXAXzifsWl
FKRUsoPjQhWeT4/vyLhSbXuQVZpkrdL2rmUuh5v2z9EjmK2oj+R/iTIEOIXI
Q41tFdnf//Z/9t2RwG4iln+kYniwJKL5AjFc/144YD2SNyXFXHEggGbBV0e6
Wl6EhBNi5xDAvMx0lmBLf/wGmLzrDzgQFiH5F96Lm7BT8UxmiefUjF92UZcS
dwgG/0/1eUqI60HTZHf6+MehuIgv3szsFlUK2DJoDSZDBvCX706hXwrs0IWJ
5HkXkuBuElWV6bjh2DG30UtX46kv1FCkvRFjstzG0LV7QHzKGYw7ypsChp8d
OsgIB2U6tLjHliW+3es0RVvlOgAvLh+LcdQXTR2LFOKo9FFb/i5tZ5DqGWy6
6oOzIu/GBG127vcBv3m3MFcBWlDkuLPvzDi4LenWe0F6uXLF7f9kHKWOkhBV
VF9/10HCfJanSQmxtH1phINYw32dH5Fr1ZNlb8GSoJcnej+IqZgjoRKNym3w
AQiNrEGKS87P318nQStID0W/1hU4Zl27Hp1lMi/xP1M+W1EydpDx7k+HFAHD
cNfWeKzAsyO4zEWEoM/k3jXMFk9d4xFXKiyjMzV6yIMhwwFH8y6N6RqaH14N
sUa36j0AL7WlOdfUcqZM+EclghTsurxlhqFtcAKKtlVOiabNGEzmoGtAHHyG
8gUc77QZqIeX31w9693H+udaj0W+zAWaPlqJsPvuoHSZfB8/RxMLJq5UQn1/
AMso6w6z3ey6k9Bhb1rlfxJG6L8E0Bdnbanz2p0UgJb8QdZ369EBJHY/YBuh
LiZL0xoenHp0h63PM1hqjBleea1+Ys05nJ7VK2jrWdL2VNyBVBRmurNcexXR
auv6EJ+xU8pEH4aRPs03XgUC3clo6nHz1Rg5yvtf3D44jNgHl9C49HpJDB3f
gN6x7q2Xu1v/gEkA8Qf6O/WSnrfkjcXaZBG5u9ja1M2Lx0Vefcd910OfVm7b
1YdMVhxI3arnfIFb1+V3T956mM7tRht+z3ioRRPpLqONSnNDW6Ugnfbst+GU
jsGRMlXoSPEDjqGKF4rznsJBJ/9W2gud0r7MboGipdB47Pq4QMu/rL3mjkz6
0xlZyd0fkdd+olkNng5IIFO3YPRB+f+ZXddJfB8Xujru/UDUXC+H5kKPsHWU
83lk2BEjQWC5sGsxplpUhGLNd4fTTp+7XlaHjBHxavdqrQzrrvr2RFmCq8/u
8c74BM4fpj/QlargUjs+4KDy2RBbDhsOLh/SDjE0hI1RW3Ztt6YZkWvUJfc/
gBif2zidMb5ZeSyn87S3aMZQtdLM45sj41lhZ8qoxQGLMryhJTfJxO/eHKAN
NFOGNAV1psc3dS4eXq1NKq5xniD0yJ0eeRAOWbz7ZGBZM0oLR/XwjECVhs+r
IktU+eRd2zeQp3vMwkejYD7ZGwe444MWY8lKvJf+xx6bOF686aLMYkGKTn7o
BWG45zbhsB2edzX49pTe5Nr547YWaqkbQEUR8m0NN99/GOuohlyXi0NkwLNY
bj3mYJzmNI4GssHDuMB79D0ztPDJsUKgo62vvC8ULMHvWhvHPJ+nob0jle15
+MA3o2F6S2lN1Lta5LbGBhM8NXjZhZ7k4y6IVTD0huh6SPBTIOuZi3d20YAV
WgW9dMhx89YTiNx8fz8wnGGG5JGpgKK3Xvu4U/mQCf+7Hjm+X9011ifu/9Mx
E4/KpyPvMpchM1IGyER2U8hjrfZZhoMIy3ugQHs91iF5aOjg8GVTIjzOqvTD
Uojtx8p+y3jIpCRfjGTBQ6Hog7ki2zrbgyjJQtYmtdSzsW5a0CcVe3GChPHL
LWYC3xuYD01JHkr1TnMXUafpNnxgzJxasfuD9y/vWkCvGB/wktGfPm+SYgQW
Mbxx+iPgd1F4iF/dtPEdnmQiPq1XX5ANBRdLZycFPb2MTuqA5D0JcCCo/jkT
pTpM8tdx1Zc8137zQL6dVpBbTP/W3DzGKACT0LGJJpaXSBVg7vwbdBzcLU3i
JJKuMqQl0pUDlt65uQ6PRYM35bOgFQ3/IlI90lpnlWakwAx8Towr9hm0zuaD
Acpoq5V2asHLCG/rF6TFPhfSCEPSxp1IQdyUZdmPIATjmotH5czTyGQV4hoU
f+W2pq/6adtvLJ8XjOcC08XKnt6AwkH+GLhUyLtoEv80VIIbbvknuE8cwMiW
I+JlSlr00PsoeLUG1H6k2vVyj3xviH3Fxook8On+eFqYSLwX0bsn6Q11THkc
m3dZDxHQoA/pzcSHFlhjNsZ3riUjCBNY/Em+3U/fYQuzTEFBXt4erljNilO+
JqqNxvs1C+9HbgQuzeaTRbZCSnycWLO1Y0Za73pOyGCz1MuWFK4Ct5xxbEPa
vKpSaKfJKgxj4KRKHX5/wWOUGE+NfpgHgrZCz3FmrRz1gKXqYXtqvRxg/XDr
0bojc8dY48lrTeeV0MEr6S+naLz+Nwn2EQHjvEHUTdeSMWH51MWBqx9sz2PL
FjYFUC0wcMNgtsX1ZHlciGTvgUQaPdxzlsZzHLzXF0G9O+WfTyXQur2lkqob
85vV0so/y93aXYpAEdvIXHKDda3orwN8NnAfFcX1KVClL8YaNAmzoRb0fhj9
1+cDgRnuaoSa0CrTWUEWATp/T/wgBZrKAzMftjC+c+m/WgwjAjx0ZE6TswSU
u6k/OZGp6KoIIVyUbaBO34cnWIvtPgum5jyM0793rIwlnJ+L7P3d4lun93lq
gT9nzn/mwHBHyHO5vOmznrOhBQSUhueRTCCxkbkXYjGyUHyq9Hi3aVJJOjbx
Vommil7mM8OU5gArI6QCN+jIRsF5oL7iXLzHVelCTSoC0UB9HlbH7pHxpJYI
Z9T6F+HGJw2ijkaJMQOhYVnzGGY3Znq7jNvINCOP0WTEb07GE2Lmb1ZOg2BW
83eVZejeeHHNqTHbxR8s7b2XrteSdjuauS7vqzBj+Rp7Lw6doLpSSz8YB8Yj
QDaI7RUjbZif528re5lKNpLnlr4Up9kC5ZZf6qnrdACwUEHgeqCVpIXQBd1M
vH2QogmKhKz6Zm1MplcHoY3vX7Xtbbbqm25to6T1rgimkCy5fHEdFDV6Inp5
P0yGfpLi98logXF8pCMLnttpucLoHA42bNIeb9knK2oaJDdHPqyHLcOqybOi
dzJd2gJHutlbwJqPtHTEdVX1IY++2F1ffROaIMb023Tj2gvgd1W8rSSpm09Q
1iyoXZ8//vBAybndUg52JvMs49vLDq7L6CoQm3yacENseJTBVtwySi2FU6DX
Tbv5izcHVGA7dVRgOkklcXqUwHz+4m+xFsJ5C1RJKRrZjRnEB3yk4jaQ4XTo
s/Y3BlhxviyaQaKtjdFQ6M2E15WsSD2xcOB1Jmr4t7va+20uTRbeEhh9t0Pb
MiYQ6fF6howdPOFAumA9SAD29ZTJD0dU+G3YUN0gke9A5vDgFVHyelnBGe2K
QjdRDL5UmKuD5dBZ64KppCpO3B1YwHBKsYbU3pY3rH2cpUeACQolNRywg/q7
gG6OUf1uTds4cprVsECldIUaTju0h4lSMTKGzAbmq2a3o4uQVd/Xn0K+TSra
BfBYHBQ3Z1sFteXOW3zIwtq8eIFyWO4NZgPd3lPwl2CtlyI5Q4zVftNdZh8c
4KpD1RBNBDJEQZmE5WujHlw3Ucwc3ypVEZvattqG7+yq54B7NLbSXAbJI7QJ
b/nc+ffkg9I4XJqMq7Pr/gOekgV+AeulRGXMHLKYgB6qx92R8THAVVFVp4Zm
P6gvU7bPfJO+XyhRzm3M+gPI1mk9PTBl4WiHZg/s5IrAJpomKm6H4bHCOVrs
V69XbwWMSsfo5mEi+zhEB1at2xMp40gBmBPcfNvy2RuHlvl2V1ZaN/cfdQEd
ZyxfjZ4sCiIBv+i4N3dnZD69S3oSGmSNPMraA/pRtTlyrZMfnNJmpFKZI0F5
p1Tj06Hn38dEkhA4EQTorzt96iz8ANPo/aK2v0A42Fc4Ry3hCJ6aNm0z8va0
DFp3tBcxlojn4vjvO/AhWw5U+N8NZttYHHYm1WPVQdWP2PyiSLLKUS9WYkII
2iBpn9uoAFY9boIjpYe9mwmSePk5hukP+jDzYi2uc/gPBX3CcXH3AIXKbgop
VbWOsyZEVwnAfs5FnM1QXV+lZ777roj5awLre5mSpVTOGd/oohetM9HTFbVi
clAbeUFJNPIqPd4EaFz3s+OuknyZOPQ024pqLWG6LN2GjL6fLzHarku3J+6A
lJ+hgf0vzH6NXBG/647sKujjxi0j7gRfqtLIgISWznUc5v6HrDrhaLSnatO8
s9/qPg2GG6LqVhjftbawNgAZjiLV7nq4Oupj6I1Xq2GdtGY2F6mB6lMmUyp6
Zev1QCOE+Ll7MBi3qCS5KfsPFIZ3mg8wIq9MgG14AnTIIIu40gsdxN0jUN5y
S/ds1/vy6CScHOxlsXTISlunOo+9gdwbL0lNmH9Fdo/ptyVAvTD4CZ1/+2wg
YSV8TuhLgzDTKJAaAeh03WZyi6QFdxRoTYVvf3JrdNKyYsp8BrE64OYi+Oc3
OsnPts2/I0JLnexPyHGKVjJR8oEPJqdbv8qQiG36VcNzaRaa/YCLNy+vrNg1
qsQg9gqHTz0ZkFFTjuxCqbi7kF+4Pi9qPZ5nGpolLDxQow48CPGtTiOEfP9s
LlBnDPSxCAmTcyuuOwFCwZs5KYPV5N1UkA+lX4dgWVJmBPC68NuO+QxvvI6+
s0dUU+TSY2Pk0L1OXNOai3cMp/VLGWWdzqI/PhlxlCnfzQlLGP5W7nFbkyZB
KjWmV3yzC4A7Bm5xjnGt5SjV4J1qhuXR2RWkKkr4pcdQWkkwoG//b+8B/lub
Zr3ewMuvQybMHxCwYSYPZedA41p6+0saI0K+eSzAUpbEkfCOTfW7/4+uzK6s
KRq1a0IGvwsDIPGvcR3FA8D5oGC7c2QzkxcHUWilmhUamGP0C3lGuiKCy4j0
zeSZKu+A2pfcGobfdMmiAboZqgbQ8vm/UIVs/hnj/DK5t7Pw9wylHDBnbWS+
Vd0ndPHvP8zJzWI1QeqtMimroQkQHZDABpe/5MzE2mKl33Y5PxRABFoJMhk/
TKW/FuKHGz5hbauDjPogX9V1X3N4dzGmothew/52pmUCxA1X7w0nnzSIy5v8
Y2tWa4GZEAko73hU5DUHOuMl+FJ6usRuGM6jxZf6UfviUWzkYOT+/7wng+Bd
b34MhTEoBUzVP9oO1YrY1O4aCZnt75fiPd2HKNJyAI+QObHYBl/mUUcQBs9Y
dEATvnhcM3syOw4Zha1jWtRINfqTKpn0YYs0Z59jxrI9HBiwIISCvqgicStV
QUL29gQfMnwjIAMCa1gzjsHGgI1y3G0aS7EVoiwfyUX1P3e/NSPnpj15mCVi
6HJWfcfm+15JbVWPv4cGXoUv7sGb9amIV5slqUpMIVv7PjLH1PVe8xI85PuQ
hG4XFKvpgu718TWL+WX3V0uUpndFAN976HIhq4uy/jUpU/bARIa4s5B7yZYI
ankJuUtLjHGtp8v1EUmQGTXwf2m3cgqiZ8lQzcXDYl+E+Tx1jt6UbCU918M0
7WKax41kQ+UU6Riw5US0rZMqnAj79UXOlnbipEMwh++qBpXuOMzWX8+Brfm8
dZ8njQXdMLbkk2KVnEvBNnZRnGb5uEjPsM9QXO3RtB8BErMe9lhPRBtwBJAH
s7/adrcV2kR0mWAkaLG/ujMHD7HrMM4jxuX9pZQoJDeFh4+Z7nf0xUosjBE2
yJKJ+MqK+7PZPu9EQbg+dAIApVrbEPzpXlSxu6b/KE9qdQOmhMfrg0vjt7fO
G+ZoeVDRmjoB2a9tSv0whP2NPcCW8l0skhABY9WxhJ8PmuB67IoqO7J5i4Xz
qKSuzj78eHs8bp7XN3hVhjZ6OXCM9rm5nrNTddETODuWgipSWb551NT/qhWp
Clu2Mfdb0SlnkKNxASNuel2eFTchahqcypMA4sX0L+POTYuIl107YhG+K2z+
PurKa3sn6f/3ubWiA5k2J+9EJXE0ofeKX0A2WnB1g4V29o21KtRwVm+QUOZF
CqmtHe2FGqn7ujSsX9ITH3G521HBp+9owP2aTfKPltTXwSV7RA6D19p/d4Q+
maWbS9oBcrcrb2tRGDJuLzYs60PmIvKbBoLHv9MyCYzW6nMnStlpDOj0Br71
LSl7tOZgbBA7x9s6R1udWv/L+PGADU4fgaLq+P6R054fsZsUkfcTj4w5+iZ4
a9pz+hO9hTj2N0IyARjdme3/NWMF3M9dp+Y7V0sDrW2FsCO6c74kjCxkXsiY
wsmBgFFqmmvxLFEeq1rC3+TdtlE0e6w8/sVGEkT7RBzy+d3zvl8yHprBpTu4
YF1cmOcaR1NPEKEn66LCQKKVY/9k+LwgKh0Rafo0/IyinIBEszPhCDK/I7DV
WWrHYxkg9rURS+lISsECqOi9w+dg8s0DNC0KKs+bUA7CsmeAG4KsewdgnMxI
UWAStcgqx3Lg+/2QAok+AcXplohx2YD5wRdn0qvPUU9kXOtdj373NLec8VUB
vEZNritXFEFpE4Jbxxbrhxt0iR9/yRryPf+fpHVejJAsJefhtecRwSyH3Zul
GRNNldCPNRuLFwzTPvd6LMqrVB488t/Pvm3OuMFWA4+q4WXQgvfXKWEi1ZuR
BvcAR3I7YyvdC+GK5Kt/xsCi2gNbJJBbeJnVzh+17VQgDmmR1putmkUDF3dn
UAPhqfsrJr5dimbypLjvXNKqgD5ywN/wZ4SDnwpHt4Qc+ptIWUQDsRnkFyK4
Z57A17vryiOh/o+q5SFMjXkABWWOMspMF22ZJeKpPJFRMMH2HZqy0JpKwniM
HD4/ZMzcNTdlak14FLQaOSBDV4GzRhcp0OLv/1i+3Z1zscd3I/FSpGANoLJa
qZEEER6cj7h9uEImJxih1u+tK8Znrn6N4ldlNBFs4GoWftRGau9YT9Q5tDrn
uOzvxHXEEuMvVT2x3AqJrImeqvY6qm7MP2ei45Iob2KO8CMYaVgQnQYoSvv4
6J4oWf21iCSOffI4qeFyfenzhzZuNzg85RiGFYB8NpHqjvZVaTvzbm6n749k
2k6Xa+vg3BLAUraG2RAAqnZMy7OLVvP+uQY0aM49V42+CV8nW9Q46ASYFBtZ
6FBMK9rReQYAojjpM8HNS5FfR/5vWTkQ6qkxpzjDW8QUSzacgl9ZBFS34Uk0
QLt1Rew9c4YfVipgXxQFUFl0dduVf23Vn3Sc5EUA1FXlW9F49UnxoQZd6Ylp
aQgo6C+jvw5aeG/msyIdxEafERbeLIpGNB806VZfENLAveeLP0OlBMBNjCcI
BzVNEN7AYqzNm0GPAMdaMP1qAgerCvt8ZVMop8A/phc7Sxs8T0ksYCiMwd5G
hzlGY96cl+vOkPb/5zUA1/DisixZWvS0SBuk3U00Mc9ml5ZtQndQtrFuGw/w
Aio7IuWWJ3RkdiRr39yJoeFFSrFkg4jMzF77g++0BUdjJLqZ2qEZoywAUfmT
f74OkmgdaxbEucBFMILK1/G02RzkjeZwWi/goXc51rFEGGYDEpPC26Dv1lbl
WILMgfaGOxHpPALSytWgranQbBKZ9LRcu1IMpreQ6QPSUp1VFaR+RvhLSZVx
0r3Bm7oiDqL/HKWpB5rGbucC8djQdmdrqRtdR7/KKIeDqupcjoc2Yl0j44xf
Z94XUt2wDnWlXrXey0R/WOc7Kg1WRIkgaPpHpxDZX7RI+ywDXCJTSlqbC9Ny
fsJrI955TLi3MXGMgj476AwucurhPuC7DelwHwRkIkzqDoqb4AOoUA4i5Ew8
rBkiebgqbj+D9WFrjai5xzUSXqFEHwbJqLjBKv0rZ+KJVAGmwlQVdw4AlGy+
5YkCOgoIO9hze/ff8D7f1LAlT4Cw3GHces9Df1hQiYDVIgmtN1L4/VkHhGm/
+jEh/3UYC1qCFN1C9DWIb8XPHG7mq/yNoNcUhTMIfi9i58KLFtcLvfjPgo5t
kuaaxTZZBg3J3rDswbRba+f2mytN/aALHJNa1DVwbJxUAsE32bhW9YojPC8M
RZluv6eHIrRqFYaMXySq98SgT162FpIU+iG2oyR12dB7H55veH+mBLeZ4IxY
OcfoVqsJk2auUC8RzHZYX5efVA+Hjf/mUWITvsQkkIXqiA92FARr2I5dV1lO
X7og1diON5D9qIV1A86N4gdTWl/Q0VqerP5if2JTXQ9dc7mlniXSn1y45D66
Eo+Tppyh3K1xrBhhO/5LMpUqAv4rZH3cE0ytnq/PzDRO+ReR0JJrzt5tMcEI
ObjCC+7ygFjKE3eVeGhjQz3AII865bQY9qpo8FXVe4iETE/PoYSma5bDdHLk
+7yg1fq9GxzYgtWX9oI1BWJqoW0x3INGdGSo05cA0x9IWSCAEz5yKftN5SLk
r4NbMLDhG13KVPwq7O3Xj3SBlLEBH3dQZk+bjgZONrIywOZaEbhi5sW1Bujq
IuF3Ny7NUbnOloCaHFkX0WCnVJYLmGSvEYnHQamrrB86bnxhQxNS5dPUhtmn
R6+3Rs5P14E4A11hfs7og7slxc43yMmH3x5/N2CcnmCRMbmNueJUfPjRie5I
k5YDXA09wsT3vi/iFKVp1IEqM7nbD6I2MCwKHQFVLPqA+9xp1U6Q7biqCJFZ
eUsSFHbw4wipjg6k4wzymCenqrEj3CIx0p+A98fOt3ya72+iWeQVv0diCp5E
UE9PNrVbjUleDBrhDNDEvKKDUtmVSHlAY27idwIFphKf6E8+0gQTGbqav2il
Nkcv7vQJGy4VWFN50BqOJfkVIWTgIdiQPBsOPJgIyc1vImh8neeT3AZeYvHL
1fzSQs6AhFOXpRMwG9LB2ovLboK17JOEkelb5cdsz7P2q7lN/+Xa9aQTbWu7
rhiDT7BaGmEKK74eUrsFP1zCFJjBLsuACY9z9xj2B5VrQ8ng3+KJ8ZwCofjC
pRbyu1+pP+2RHQLpTEC83IwMy6OkExwUycTRYgE7SK5BLXfu7WOyt5wSwtB5
xHyycn3Ki+Gmj9qheB9/4tVb7bp92nr/MWDX73llluQxE5436h5ni8pW8g+6
R/0meO14xOuVz/1ysV1+lX9ApPE8mKIROfXH1LZ6Jv0F+nbxE2siHsCteHkU
2Kk/+A19YSrqoWm9iX/B6NalVII0jioLeU/Otomc5PEjG7Yl9uUIsBJcos1w
rN13rthCSSmoYGWER1Foxv94+PpKo3GrujzJaZ3BEHHTnSz02BaW/fuDI4Wp
mj2cjlbhAKt6EN/3kOTjRzX/tzICHdvXXiBUUlq9lbZoFJtIAUUEEXVQvM0K
5uHp4b8sWMuqR8Tb0kQnGAFlKJvP3PKr8CE0JIAsaPiXzkFfa15T8PC4wbKV
n32tUelKerHDl0e8xpkppaSDGvk/vaq/BLDNiaRbvhxMwbLYxW9K0b5rmR40
VDfcay+zN0v0yNnOaCgRvG9yXalVNcS432FZ8/Ff1xr4kr9xCod5I+X7d0mR
EDu5dfDROF3hI8qOOTnp4Zv4xyj+qflsQgQbHlYhj/arBSC6dASqY0Rkh8b3
kqJvSYkR00PYhvu4oW3+mL3uVA33Teo4+5F44n13/R/7c/9ePqAKa4wiTyvv
ZxyyKm088wlYIvT1xeQajtOJNKty+uA/b14Z9CXZPHsFWmL01RUp87oDF8Gk
cjNEeDag6s4UzS7GyrSson9/lOYtz+uNJPegW0BWO8xq2nwcwLBb4uNqpDYJ
fsiWHXF39lQr0qpapK7h5+8ODVC9U1bIybqYaQslZ8MWqZEM89pEthHYUT1U
yyKFCdy4SN2qActay/YSGVLuqYHijDKIpLHUp+cZGtpovD2AZdkg5nMQZFp2
wPUEjZsYtZ+x4w7Qq57aQioiSVDWOJBv1jenuwao3PPM4SL+BBE2+fqbwQHX
1L6vSwTbp5gORBly3k89/1v6SJysW99fbPEBT5R+9dPYNJWYSVFChHuH8UlP
hFOZs4LAqlZJUPdofqDmLkE9srpweI3F9CComEXI8ezvijANpfmze+WU+TGL
iLC9mJzIbQJmJ4ouZYENUPCVAncevVogugrKN0siLU9t8Hlh5BCnTKMtv5qT
t0BYP9JGYpBXGe1D7aETeVQDCqX2W78OQ979uesu6cgTFswvSSWwd+Eb6J08
jQ5lyXIXRM/90f2h5b9oR9bnXvkQNFIHuVyHcmdkaSE18SHg1uma0wKyfx74
QHXLp0o0te0co31qCZ0OlMA5RU3K9XM8n/+fl+RsgldWrznBb0G3fZ+AR83s
Phw8OIRrvTU3Sl6lPuNr16AYIcoOd9LdHXQJqIQDUzfIT4YP903Z4TGk8l+K
JhYOqOlp+l16G6kpIMCQDPUTiFu1Nyd1PVik5oKRqsoFLkJQhr3rbpyriIlU
51X2OAh15T4NJgpYtUKsGKymudttiHeMR6eK0LfQbXJGRD08EO7liX1u6OTG
aa4QldtyduiqfAZIi1gtVzT/Uh6rhyDoMVhVtnJsBWp9ReOXxeOdgzgAn9zE
4BgMfe7a7TCd6kxClYJRn6qv85KSaYzgkxi7wrhmeShFTQTYU1pLQk8cr8fT
lQxPzxdpZUNgRojLtjy0ap6df4rJSKAXM6kd6YBtgpS07fjjlE7K2gELYMcc
mrDOJDE7BOMdP2jM/q2brB0DQ+5nFEaR6kO/AN0t/l+uDSPBhwHLS9h4z9/e
qQLAToXIducFlTAcx+ufW+5GwvwHS8MWm80i567sLmC19uLnIQmTPzIZAFd7
l71+WG46NjU6XTO+4OuLR0cZXWKjNLcIg04WAgkcAMSuaoFXq7Ssni4s7UzX
wDReocn6OnnqWI25x09yngb44Zvgtirxc8lXgJ0yyGRmXYGu0o/i/ygWiYWk
LX7zfpPC5/I2YBLzra/BV2rg5tW5O+B8Zt2dL3BGutguXFb4gUMgybuxB2jb
BqH3nOjnQN8ProKJQCEWrTzbN3vQjDVzHZVO09JBqpQK1inEnQ3DfsU69CMV
hCFFEVnNexyLNHRuhqOiVTugd56OzqUxZGdnc5m0NTwq1ayQ4/Lc3PFYMVW2
26ZiizL5Boa2Q/oAi0iK914P8Azt7uvkq1ycBKc20zJ8xwaeYR/JmK3nGXm8
vucgZzuHkJubEaLWUXEJ8jtIlCjiyNi+u3ZjUwCd1dcymH4c6SPJhJ20iB5i
AhXCYQBWap0xWgEv1FPm7to178qRCdm9ZATAy4B9k/wYHBzGWfDXi0mYz+Go
svdh4oEfleFLf5UmEc56obxCDJo0hmQOEwcN0mAY1TPOMf0pNNDZRsgtstOf
rj1e9MdMJl+GndE8Rsyr02ab6E7B3E8NnG4qHcrZKSXLuBCoriAY9Tbd7m8Q
qUYGWwWnPUJMcRVGHI1EzN7YhEPkPCXWP0Z2vtZl/mCwVcJi03jMCyarRZAB
KFGOfpzCGUQpFtBDdHEPy9jhlVzaKaKP6h/BFzSYoWn0ffrh/QpBtE8AoDGP
uDKw2Ob3NQfoBEC3S5Cfo7aFyL3WXSPfdbohFzWG8oMHS5rtBrAx7GUQoXHI
BqYd8yCFQiCNkJQnbrZ0uA++IuEcb7IpTIUZcj3rgAw9kSt9MIeZJzb5Biss
I8XP2tfYnVq0JJBNtIE1qmbTUSww+QzXV0VxNcapd5QvIrttHFgkPJ5+cPLe
V+df/nJmVfPeI1Ybj7arJO/ha76SNNKiHocm16f3Fmmo6us27TbEAKZqGnY/
NUPa56ObsA6ddj6FWglwWgRV6mWWNvuJ3aqDFs5pNSnqDPTg1Dxx9c4YiIUy
sVVd0oNHYM04cttXydZT5e59OSbQqWE9LAkvo0yIKwdDXNCqyya7L7lNWDgg
4/b2NdrJNkxtbidNbEkQcZgDJczaHOm17I4vwcNXuu+b6QkLzh0Af+fJH6rG
DT8NSY8BJfmOrJoj8WiHoFl39Bv3NpZquavIBxps1XuaKf3aBa0ekLqCdZRh
25TfBAPWfP1qmDYKF46GbdGA6tNdkNhejhpfgc/iaMSKpsjvZ/2ddssvD5VD
OeuBywL+Noya4AP9i4J6McN15tQ2ul6APO4RDOZB8UY/hDvzet/evbsOHN1v
d8DaAP+aIpE97VbvlPQVlgyR3gqEjkPa4q7uUPFm9LmbpqGK3MlZYPYl31Px
rloroeorbolP9SxHJxtzo1xoTtKy15M8WDBbgOmsw34KFWvFnEIP3GSfCyx5
nc4oNVmX8MHxNNUVj6SH2ozk+SCTnfsqpHDF99gkZ0vBbBqBEPpF72v0y7IO
3lwDojg+4g7I86HhzFgJyKty7ptTChxZC3JzsbC+FiNp/Fv4GlkyZfDKK6Qq
QKAQh0Sc7caf4cHSeunkpjG0ksazfP9+pl7RKY2yZyqeDC+ISohYukbZEMw+
MAnRfHhc88QEC+YMxBTTqwjirgHEOhIvltUelmvsvwa9fytBS7nKF2FghHc8
4hZlkJAIA5BPs8tqLKLpGCGLfhaG8b+t5EAY416G4xZ97fEyMV5aCHxO17Cq
2GVqrD8enUNJQUW4PpX2N8Gs6/WTzB1WUU5DtLuiTnO8hL2hgNzQJKYlIEL8
jpm55bbllhSwjcjvNltRNoAOBOOFyBN2Rz/0p0iWroU5kz1AFhron6MjeF8V
1Zi2MNu3spVSG1/9kvbkgsJaLQcvaujzi7qTP492rgkVPdDJRNpjO0w+CiX6
VS5UpTGFLQFXsokYxC2nFTFoOvKr+aqvnYomOGR188tUdxabIKsfH84jvBTF
qLArkUrX3QvauFhcTrCvae9/Du3rLPfCzbI/fPKX3dB8z8jKB6H1aaYLebcp
eLsnqqZm1iYbnLT3ljzPi40eN2lQEe7Q1MO3/cMOK65e86+BBPw4uNfh/I27
DKEC0CLGKq8hLBHo2yQWDA4hBDfQWveM3l2ZYDaa45U1PfUmweixpDkDHm0c
p8ZXciw/gPlXK3qsPJaU1M/1sM6plYZjRKOgbsCMKC4fpNh0ttoratYriRES
PRERaRqSvJxmqFaim+h1MjOVJ55Cz2kG0SpBS5taq1GPKMwV8uFLjkTjgzgX
Sxkc0zU3XN8vmA2snWVx2AFmXgU9I9zIesmLEN1wyBUO44M/lsWBtc6fPanY
ubA7FSczrD17Hail0lTQZTuFTZC82ivcgMi9rMS4u9N3l+wIxFYWwg6ncUde
uoLMufCbG0WG8kTEUJKDshzrvqucFhwSFiUjMTQkVrOuQ1Oh+cVncwrK6qw9
Z0eS0ybRX2E6ejzcrpexXGwr2ikXSKLsMvZUtCS2fus6c3q1c1mB2QJhyVLQ
nmUgVQW8QfnehtP022uP/uR0t/vSP076KaV2NKQQraO3OGhTKGyWgpicFWQy
gPBsQBg1cv4LA9qAryEf2hIDtait94O4iv4SzSerX7WE/9ph4+b8/u5M3dGa
DAB2YSHty27+YXiWEJ7V8abHYTOmjhC+qVvy1Dzt1P+CZKE/FGpWpo85W0gB
ofJW6/icONBoJE5UMvmc1Qy9Yy/qXp5bj4Ipkaq7k1DWaH7STL9c6m+UGVKD
kweafD387xMELnYVVxTe6NgBGuw6sardAhSgd+XahsaimgLtErFKdI6qHkvR
oNqFKLDAnghiDsa+Qs0kQBFu0lE7chK7LIK7HX4tHtClumV6CPxmIMW0sXKg
kR/ouOmZe1d4X63TYAWeP1L6g3GjRsfJ/oxogxfOpCo+2nl4rgGzIrSa+RWe
q6wM+uat5yXBWh3HiCeqd6egdxB0YrmqECbIByocE1KOBijGljkc7q7+TukK
E5NkB5xJbNP4AnoWXQEsYOxWB+1dBzvnfxSsR80b1sIHQnu10fulTJiao7mr
bhU/eMbTbj3PgiNBAC740vHGdGbmsu4z+Mbq4jBqyFfLmLpx5ajSQ5DJproh
viQejBl5XyF1Xzqmqz6oKTlfOYzxy8PYv7W/xbOaj66bxzhMNAOwKl0nVTC9
yzaZZHEEjnwAZam6vl1QOCGwDvHCSFvR7x4euZxPgzIhPRfH7FR6vCM5wiNS
lXnSZ85tLdBfmy0y+w735fUL4/pkkZu59/r4oqk2GE+swEyXOuXIsYpVRge/
nD2fOXfUsk/jUxlJ7Auf1bpiTcSLoxh1apVbvCcgW+c05GoATrhwyNUipdMf
p8PbRaZvAQfrFcEvWt7LPdqOVraZgrYyPvjHtK+P9XTinz++ThBEXHt78Zhi
jvVvjuehabZtX4VxuLGNbYKdLBbT9AB10C1ZdCIrgiZRAbILWD7o+D8wVNju
Zo0YP/3TjG1ahln4uBIHkIJgO3LKnrrUnv6fypuz+McEN+I7bxq1BKQNlH6j
ouzEx5hRYhON4Txy4ZXMkUT1YK7mRug67nNg9tw99sj3sDzS7OVGtHXdoyGs
ZsW3FK/LaqzCVjChTqvkNr7rZ3awI1L9ksPf1Ah9IM5O0ZR/E588cygvHczG
y1JX3frpPHwby/0cppMPT38S9wZhmckZ1lAVO6c9xC4Ms/bK9u6+irXhIsyE
R9j/DWh2COG1sOJ+PyiuD6+DTf/jTzOhqnegiNSHmVR2N3pym8xwhUN1bzqR
QTo832FBChThk3cDdEr4ObqTdnHBl8ztFjW5FeKYTHRyk+antzXjb2w02jYy
jk7FKJzKsmMX9B2ZrI6BKsecELX6sJxEVIX3ap6yu3hhSNjkXpzuc5yg8CSl
JfvL8jW/mpx3OWXvm8DfPpnyLvjcfAHllN4M3dXyldCfaVxXHdiN9gvZ1rN6
4b99lc/bMSljFDLvT+taEZK7zUpKMena72qFVT909xu3MDQP7xg2IuiAR77u
MaVQxbN+I+WINDX4jBpfx+v0YR83i2s0BDjQwvVaV+ceUt6D0Falg+qa+zkY
8WQscOWTLMyoe6psfXf7Zg0GLaZxJNLr4JgGb+3RoR7HpQjmmsh0W7+qAnt5
W03ZJtFTbyo0I254JeCUWet/yk5ICNlzvYB33JgeIZ8yL/o8meFpYSs+g5DQ
515w7uonuiIamFcooqh9zEvDVmrjks3kojurPHfGebaMPSYR4D2r58PynCJF
hf7sp8Dz2meCPDA33KYofM0V5ba5tnugOyj73GGlmUsEkgXWHTkjgdpIPukn
jSUE8adEshl7adH3ptkGb1R1Og1iHpDa5bF6eAGop2VWJiaPTNId640SSV/u
ZUmgsUGXBjfkWJ/d1v1/DEoZBCdEBY3DkyYREzvNX1oBcVHDQzTMq5us2Q/c
D1boEIDxLkAuSifF4SCdMusb2FwJiOH+JXX4btGB+dGWPYX9wZs012q0UBdM
biwyN4YWyNsdYX+EVIfcmVoBt1Sff0f2eqpKEZQhOXNSV56sM7NQebDPkjbN
35WvWmVcetKpnY2yY9V3OvOt4QVC0RF8ZFLV6o9/6ild+8B8jr7XsJiAIYVl
f77LZhgPNNaOvfOekyjogq7+NKXWvJABg7r5i32AP7Jk48NUeUh16N7PBWOJ
p6Pa7XkEe3452Tbu5LwHqrsOWtT/474d3CuHjkptuGiFyVoWZePmkLiYc9la
ihgkub5gd5bNGDCGK76n7qbs/itOmxCZ59cwtywPbl96PFvBaNOWhgRcRAMd
QGu5QDUM5ez0+ZHEEgadjRa9EK5xHh9ZPHhmXpb2MEL4TivNyy+/cxxqw9+u
kThzVQA6d5e+Wlkb5epTwKX7tfAQNaKGmgFQDA1rO0xfJWKSdRzP2Zf7fBUx
9GEt5rZaLYz4apZMm34imF4DK64yg4YDO3ZNxAVNxUS5lIlEoyuggBhM1vC5
U22+E58n6PXhADyO5S4hLzEOoz9Dmu5zyMCZos7xrxPghEtxnPemItLB3PHZ
dC5wZjWEkpJcTp231QXlDtjOCXTqRvD0JVxV583GcMV3+bDIEnEsiCVGgQwW
R2VB81N+EYPAXCV5utWESGHm9F4gRCaOghdFCU7GKXPTIsEZTbfdb+16YES6
hRscHljId9Ju9tI+sQfTxe5qNkuDsl+X2DdFk0q6bJSZyXE4dpPr6j0E0fEk
Jp1hkgmeoo5kDYvka27DSZNKF5/lJfKrrHYE2E/gvJN1Geq9vQBd4bZE2ETR
5UYdom8KLxzbtpi2ZPfu9rHiIFGIqnzmP8cyn3yRF6hJoK+kWhIr7nu8rz1c
5dp2/BLmb93fJcI9h0QjejEoqIw/5z8D2r9mY69FB+hy7i526QzItGchTppo
Qzhaew10NhWHTilpGRFE/uTKw+ZgBrEAVvWLnWgkHq5ZKpf3mFg/fOYCF0oH
2OwAhq5Oyai152eqipOXH9z5fG0hfTnSre9MwYpwIMZpy+3RTwesHuNttCoW
6+9xq2iyfc+aib/in1M73Ws1/runK2iVp42QieYDNXyUao33s1Uw9qCkAxS0
2VhJualqF6y4IZ7W9e+wQdXG03hweCml1KVAqVvYohuocWrOyImavPUImq84
zMpLiiYoUKIPmTOeTxDH+VdD0Dhiqalto3u/zQ2JpM5T4C2l6dJrXH2+RgAJ
QMeIqf9Q+K9PHj91O+9lq1aryk0ZP7RnCW9b2vP97bmoBzFtYqAPQYKsTMLZ
5ZCeOrVcAaT4zJjdzF7AjF3ZE+b9URcwZ5p3ZApSZNqiIwqhrOM//98tmAAt
Z54mAUggSiJzsa1IlphJk37Y7yJl1HiWLhCZdyK8S+YiHOk78o6pdpSWk07o
f2fVsaTcASQboqYZKiIh9jeq9PTQ1ZafL0sgJILgIhsU3zy8ybXWnddgf6sZ
q9zRT90L13gJ6VAzqqN3UtRko0YLmNNE2gYy/UbaxOeV/m5U8GLvHdNfWCq7
s96CRM+FNeXPTzKBtHkRbjr4xsuzuz1dev8sxkhSRMFyOxYGPxaIxwg1H+Ep
1LoL7/pJncI+bbNkp79mcG1wzK61T5QQcKHTloo/UxSHuiXKp5vaOVe53jZq
AbnCRV0sd/p0J1DeGqNGzzCwdcsFa01O5ys18yLkU++cB4PHvOePbvo1vOHL
+kLsz71z7vnnksYDMcp+bKdLAKa4czuBc/3DVh7aUZ6PDCm1hum6SNkyLNjD
ITq5S7Ut62elzNgDFXVcrQNu9SPXBciGlskQ/oeQx0/VxpO9ar/InfTzmQxS
OGfS5BpwMr6wJ7/w1vvZ9XnN9DjJkPMOtyH5Sai38NXpyeiXYxeChZ8likPV
sVNevCUZ7zfNqp4TU6QXokvcVqjwdKR4BTsLAz2tV7aBt4x55fWgHtCrDokQ
mZs3Lp5+pWhkyNm8G/InlA+BDH2uqRwWPtGiqOQJXnYAcOzAIMtqTOpQQIxA
aWEwlaorcR1zb//Ceqd8eTEe3pHi1uaZbVXU6BfEnRJMhqtwQQl+QSCn5ndI
7hs8yresqXu0Iq1tQf0AJDoIMOkpTYm4gLZJUJM+3IG4A/jZmstbimXn4YBM
6IXjdzXG6/AQEDi66d64q4RvfTri6/KKs2qmc6UDIqUqddLFejUYCoE/t2JX
w76Ih1UAg4d0nQjzXnNGeuQbbETvwosvObO4uRa+WUgL5MkMR8dGNxsxOffB
1GFcBCrYzCcKMoGBj79v9FAAIsbL95NCf6iRlzBXZro2FXFakvyVSs2tKFmc
lEkECeL+rPMO+eBSXElkVi1hrTcz9z7bYaW/OcvSDN3ZutHIbqFdE6GyNWGC
+nySwcjrxlHeeC2TQXkL2pig2Ysxbdr88fLw9M8UUN0eYTc5Wwr5RpCz2jyg
HB5Meo7Tmy4R1s5L+xr2Wf31a/Y6S+Y547TfwPfVly/cnxF6EQdK1Vmz3awW
tHz/YtmIDvQ7T+7CDIkHq0Bp6r0quHOHRaqcUSdGtnHPdkAvQZqroPQBA3/O
ozzwixYxs9jKIk+TfVCPdn+WfTOFjjDNV+CogAF3xNp4vm4ah4xOjZA0jRQI
ew9pHQlwIKtgJaGsP07rUCmlAH37zPUCkDQJ3Og6ISSkMNbGd87ImZfWAtMH
7CJc1TU32M54AHtgrQxHS07ni1kqbV/N+WJYAwoRhiOnOfUy8m9imwfKQ3rs
/At4BHPK1sW2UtnGU7xeRIQVH/JxHBnWDcdVLDf8LNR5GEt/fr1Iq6jvrrkV
K0lws9Z+ntVDxFV6kSuvyF3LzZbr6DCXjgwehmseahRkmXQ783OLrTzzlMKh
O1A4mlgSOwHdL2LvtJJH1uFihwObAcYlbV6rdO07+XwPwGQzyb6EA+EVexeh
4s8Z6Y5WHlnbtOIJe8gdUxMnf/ZiVyXoU4cCHvQ9EePbDPyNi+RU7eWBGqrH
BM8RUB1N/GtIYkBOG+RWfLAuiTYPTCcnr1bvFZQlUNXrodBB4nqosbvokihO
W2woKOQ+U6d0Vv4EYavWsLabclcXB/yTEzcFDGrWOrba6nG6grKNf6B6qCUi
FfSNRucjD439bboVbfy/TRLYmGPvN+9i033FCbxYO3da1qphcThXgSuqyYpm
tpI3hvRuM+Npl7aV018eUIP6+ziPBBlBkmmBFTR2Tn+fd2qB1vM1fktErO0u
b0u68ExJY0e8uDizVn4L8G2MdxezmJuJ36IvyBmlwi8GSfkb72kvBQ/PaVvz
+S5XtkCmrjqoipCGKGVg1yPdfccwsrQp1zNRIaAYRLRSvEEsMUXlvtYsirtN
YeOTuv/hCHzmG76rfE3U4t8NoGtwjtinUCFSVAs61iJeYXsE3FIVY9vxeaTm
1Ttt+QaQyjrBtuQLJLHGzgMeHn7ZT11Lpfr4pMkMIeTPnZrDYuNFXSpv/q/c
Lzto4jDx8V3JbVCaJAnlyQyViqEYxqmyhlaUrhSiz6zG6hl0YRhnsKwKQUA9
6iNjYKQwUsK4n6x7kfon0E8KGd2bK3ckGs6SwcEETQBRC7CHBFDgCijnI9WC
EO+Cm0bYkMS+AeoS65eovPQtOU6sRxk+Ql6SXJh7UvK5WpoFYYc+gf4qaQRG
ZRlM0/4IGNPiJcJYX772BP4ovahK4KbPdu46B5KI9MP/3s6arokGj2kmfqn6
HheeACD+DZfftTD8iKVEJdSB3hAkTBmq5+By+ooPEGw7vBGC/eZIW1Xq6pye
4VdHLD+kH1VrsJYtjZEyu1+VcMdyOiJV8Bte+OkJM/mzvXTFzbIDgVuAOETB
i5OKYmPdHjal8jdIVvKNGoFj+zyvPNkNW3mWJFlCk8BSdUmm2AUFkISCXBKC
1XCqCKlvyH1I7CsUxyWS585ZMKrDLaxy9A7QTTs09kZgAnl0qVyFav6LOei4
oGCX8HhtpZ56YPFgVZxZh3F4PX+RCCbH7OOIpJTB1iQdfj56ddsV+uVZ4Amc
QjxVnKB0TykfiAEj90dxmIOnlkSqirir6/tqeiSIs0dF37Ir3xCx+RDAZ5pr
yXiwxPioHp0ITgkJvpGsLpg80o93K6K4RyUZA8RhC0HsMxFcQvmMAUwUGycA
U8mWSxZv/FPSQ8xMw1k2IXed4xYUYStHRpzRf6kQog+xuMqhkfxanscSLuxC
OZYw147HcOCgLkwI4YyTdFyrPnyIjF4mcSjIj+n+9N0abZigdghWCxuKrjAM
7qCtuJAuHomlwpoPWLAayEj4xWoPI7S1L3QoTnr5ukouXDI1wrd7xizB+dfs
9xbehFPrKQm+qnBeAUihXZluM0UANBJZ1cz8dIAYL0jam1m3Ez828ResfCk7
tWmBlGdsBBcocmVFfMJFCXW+NUR6oB02HoWssVmeooIenZ99F7ZOKeT9LC+Q
5OhBlmpjYqfckGexKNhaOaQ+Z3XX8Kt+xwq9sPNO/7ho0at0NdRcLQ2rnc3c
I7Bf7TQ1g7kGHz8Xu2GBiD6zudPgjiKXTQDTBRmjvddCurlAaRmVF8mP8Qs2
6EEiNrUbeZ5z45nso+/DZbZoNlRGCyyGPCQF5F9HjLa+HWCi6rS6OQSfqxOd
ma0k1VqrXC6hJKsVSJoeRT4Akoe2aLV6UiC4qXTRY5ui0oLVKwuQvSVX79wv
Jx8N0aV+9DXXh03urj/klCcWKVXzubf5BZq7tTq65H2KhBNS5TNW0nRyOnvF
H/Xa02elrOnUoqcD8W37zJ8FQmzi14rD4f6N7JJavc5t8AXjR+hLCMlubAVA
hedKtC1wiWlD9UY4pdbkNk0oR4kwrgypf0OyU21T7utbjOPy8M+0HwdOTt9I
dPoJ1kuWsHvwqxwpk9O0FFeq7Ng0ai5s/SMZ730VSn/LHOphA/HljcPmnpjo
Hh3fN7zmIcLe41kWBhbGEmHuDgo1ciNESf6PDSUNMZ5M6MzIS1HLwsR4LwSk
BjZ+cOzfCNVlxS34z2vgxOlkEqatG8Fd8FkowoBqbTe4ZBt0OU77Q05RDWLJ
nu98KaHMT+GlxBGbH6dSN0uvm0WX5rTAvc8lYgL3WFTTF3yUN3RVJqAsKPyn
MnKXAiqMz17tbqwfX7VcdlehSyaz6pWLEBTu2UO4gUYCyCpRZYudP50cWRsR
I3DXdLfm/7oIeo3FIubthY0NX2JXLigyCAfQwMrALBzxr4jHU/BKP4V+GJOm
jif2CL/YcXcybcVgYdApC+45erVARB95qq1pO0J1m0+deIOwXCrn+nUlkAhx
ikV8jryQy3x2ReqrV5GRtjS3RbL7tlNEZoxSJ01RsyrmkYtuo3DsZihfof5Y
sljSfdHiaWDU80GFODRvZABaPxGt9ZBciLZnYOWGXbvRRHGVPVZ8l/gcWgHd
wnNo4y0VltPT/K74hcaH6W3D4YQQQO27ZRVKRR/TJqPgGjHlQHwPK4YPwDUJ
mv/V+yF7+/35ey8tqjB5QgGemRHmMwhZijnXn6P/4+erM97aITiQcA9qvcHK
hA/KfJM9W3Clt8CfWKfbE+mjoNAJ5S2Fw2yMf5BCMEkU6NYHmlrOGD25kf3C
G0szpl9exfN02KwCtMEj1n7SgUO5y0LMuQ1k9YQyPD4lsR4qRAHK/4QHQTjg
/+VhgM72cplTRwnJuI+mfWGujV1TJPLODAfw/HavnVrKA4MLsxAE4xG20NBu
A+o4t2f/V8YphlKdvia0L51S1vUMtGP5sgdVeszG/Wx2yqYxw7k+JYnkJcbB
gJeSyr/w3fjGqNqPDWFe20cooLgeLVFMtyIhPdlbxnnJgSh/RCT9PZu0xX3C
qqEd6+nSOWd9E5iJ3l3U+O/y587T/U/hNFwaW9u5ocNDGJWDcT+heBtg/Bwg
kQZDz/ZAGYvDcp09oeRGfTKFA/obfOUOy5MPaUJoW/6xfi5jx/a3BmGeZacH
HBCMVkYkp4gfS9l70hHRJHyzuofKwcv7j4VoIJo8h9LmiFoEGZrpftEOHs1Q
qbDZ27QNdzlltXtz0eGrtvweSxyqaxirtDm/vLjHZEkZLJDf3vIwKIRcWgX7
W2TCYQXXdNMWRlLZ0oPt+gX3RFw2ZeftCtN8b68cP4lUtmVhxBCRpcTYzbvN
C1F0q5QeMWHYmVd5LryOKG7Jkv4mP82um8HY5c9Lr6uh8ciQ6rjegNp41o69
qFnPBKi88WAcDPH2kDfn+I1OXkp6BkwrxkD8vVPjlduclAJR2QIgdedHoilk
GLfRQ0DIP+ilaxtU0VpT5n1o2cdPGdUp9kw/MD//W2+czQ35/c/sGmGXRpeS
s082AlHPzG5HYrJaEC7xvylvcnAWVXnhlWJlJoiRsVqJFWjLmPSnH/kS5isN
Rz2gbsnS9fIfCGC6usDTF+gILWAtYE9HwdeizfCl3lmlhPlpYvQZmdMlyrwd
WMsFcVHysAkmMNC77zov06+H4SLn+4Y2CZJxepMUyVwZ/K8Fiu/epj/EN0YK
uqL2TV0Ir2csvALTGHE1JK1CK9VYww13QU7L7E0HbGnAVrFZzZoDgD0E2CLy
E1VFFRmNo4XfDT4Pzz16lfWMALHThmPCkTXrbzEqXAk4sGXwhNlUVnagSQGh
iBYDmsNRdPREFVHL/4ECTvaIRTRblg+0VhGYeB9vxrvMcQ26NKgCdxHv9lr0
ouWmxJpMKWJs3lmGQMaZjGccKTYWebkXucK8WjZCgT9LEEvgsa7WvolQ0J7t
KTRcs6zzqGfErkqFcR7Ky9vl+7Z6nKRr8rpWkAEEbBUheO4PAEtBzsjxVFiQ
chpIOk2laOQHqBJHLd5yVeqb5gY6uDzHURDHyouoi3ko0xuopFdSFKvSTchn
hmV86v4XdnF+ZAa/DEuVTenF1lCRaZjCakHsLptYepY5mTHI9turZ5hoZS+o
fu8G6/EvTU5dkzIj8CXheeXvvH1kOcFAMNaLAB2TFGzDSFLod2MKlgIqy8sz
t6Rsgw3qhbMsLrXr+jhFgpgSVvFjyg8unkoMDY1pn6isN7BcraWj2AjIQ7J7
fVwZue0eM7RsVukSMj+PWjhUh6c/iV97oGL6KNscGi7H3dTRnnm4c2jwHueb
rz5XSM8JWCRPlwex8tu8NFnVRSZ3y8E+WAI8EOq16PO9HixF0vV0FDZFnqNV
6NkFd6BPscqGFLL5KAfkXuRzTYavBsMDAWvIMja+F+d4LCBTsSJVzlLDvUzm
ojgU91WhTNo5pArJcxrPkrxpSLOvrjIvb94x9Cp6Mg6GVxU/v6C0WColdumy
GQuJM8PurzaDaEa0bTBvln4HXZea6TS+tkeh42BDtztpuf7m/LBIOpzsloe3
0kAiD740L5xPTv2rS/F6/Uezl04k5LXA3864JEzJhDo3eombfI/Zhe1ydfwn
00agFZMY8pVW9E1uSbjqVCnvTG9UYxLVd5eFZcelYybYO05CFf1xM+5IJ979
isRLaNeokTJJ8SytTTcbtjX4UkEN14EouJnbk8lfzBTWUSJTV6Lg2EJqqeNt
NZ52aW7sXuweO+enN54YUcuNQbjjw6yK7sBZgKZiKlj3nRgmQGRq7KNVCH0K
Ub/gvx1GL3RIfR6inipRzhJMVaWvLZ8Gj9RbejDw+RJVVJU4EIGnR1QicM8e
dIS8Q3V6g025K6DsPK/DFdspbZCvYx7+OOK4V9A1QPqIhaUC0B0k8JfFATmn
Agm378VXSnOq8CYxR7JDMRmo6bP9QGOVOg8ddASoR2rSWd3FNoKgx+GL1AIn
4+AkWPNDaeBPW8L6vzJ5UUBuUWcqEajzuHH3gjpF9LsIp7M5Wp5dtzYWcYt/
/PFcL3QoQG3n10hP0zkuaDiZgYZyXEm3VzAIVIuit28UJYlkZOYIESWPe5v+
5L05YcvJv5df7sT4ZiwwTZvcVlbDSx8msv8W7+TmCgGBrA0wDseqsaTLicSG
pEtqv0A9Mkl8RMG3LyqMOAWjHCkCRAwQNBwOGgX6KZWoCxOHhXOO2m8TK7vQ
ErwUB+P10G64T6YhO8tPJz4vOQr1yPl0qEQnUMIT0FUkl4H8ofMhl6Sd5IDL
WQuRPuzeNe2QTOEwbaUcgO2RFLOcqRwnQpkBH6npouUW5cLE94gf5LYxHye1
gXwiaQEfTP0Umuj5ntxTXamuGFLzf0hv0Ysd4016y9T91Ui7Yaz50qOpu/tN
b9uBelztZ8EfJY8WGbRQxQkkuDzu61Z/9OajOJSPu+uvycqm4gQwVzYwMSdV
+OIV+JGdMGa/95H1y435xOA2X9JdKDgLzDJhxNd5KQCyWZx8eUaIWj+Sw1uQ
XAKr4+I31t8EBnI757yeBlmse79yCdNbFrn9h5K9LOqAsljGsrYyB2FeiqTx
5zOxQ5kKc97Y9QUSMRCBGdeSws2hxK6dLI03pSXUycGSteBhkw5sHpGght18
V1fOyXk1knQY5XTk14JIL0nLiZa2nfy1K+kvDBrqrb0vJukSA7p9LPRIFicM
HBeDmbBazKMycxAkK9dzJ+NPvPsKHjOmg+LCKgfs5kIAYl4CTrHp1rFwj6sE
kerKvAimzGgB44lE5jEEspij3PNtEiXinl9U7E5k5bwvlGaLCU0qMHMWn1vW
tDFTmcXngmA8g/HuyD4yChWkgO4BAkPOkPTEd9C3VFfHbZBOJKdmsDDXNl5R
79HFujomMUX/hqF95fTAd+djhx4gbKzJRDWCjauV15TGW1BfqekbHavnY+vq
KgSngncDha7UFzIxBrA8ab+ihn4L1tNpSwkl+j6lyT9iXB4KJf5wShR0HkNh
sbzgYx2wgm4+fH9xXF7HmfXdy4bsox8LDEAuVcsgxxfhyZTGOMtM6bQ86zIC
dsVdSDKQFT2wOIA7cmFPO5mJvNdX8BcaWAV2btyzohtSMYndGyRBaMhqi+L3
LenA/db5LXDI70P4M6v+4AE1zcz3tTQYPsYMOxpRB2rKSFwRBzmxJSUYMVAC
U+zCpKSEw/JL0NANsmkM6FevPCqRagmBkI3tTxNpJ8U7MaHZjufk5TQDncWM
W+VDy4sgwdpn1QEfDCuGUypfwvsNAzdYS76aWyTjxXIjqGj322ZKVoG6pIy2
UeXUm5pzqr3fb0ULkXlNnLhX1+REpdqe9M8YKIiO5OmIDYZ6YhgSIRStIRaF
QblC9LXiR5GgUyaek7iBCPWGe+7nlC8CXVNrebL5z3n92gCHd1SzrIX9VXON
H7vjKQrGhkZr4NweVo8arUZ50djnAW3gTJq0JZpj+BD/aKb8fzR/1zAB8SPs
i0YMomcA6tdb57Y4r5oPHTRe/kGia7n+VqAIzkIW8QayrN4CxSNi4Mi3L5o2
nzL6nC+nxklJjGPtdjDvvIW11x9Y/Ci1Etc3Dbtqdf62XzG0y9bFLMCCU6NY
t9jeMmHsiAOiQx4pH8/k3A+Tosy+IVYWzbQy84cfIHY/+l40U+qlv0ErNw9m
MGRY0Mw34rDHuc2Pf6ySpGsy7jKkYhLcq6y8I2NxKWc9oHGIzbo5h+T8xmmC
YETJlHuJ6iUVA7n4bUHsOEIhq8l4tgWmfK0d+ugl7sm7NmInXM3VeeCRSF6y
ZKnPbEOno6ZJxiDJm9gLp7zeW6+PAN3hA40v24GLLcFJeWhO9sKmAFSZRnK7
5FiRQOgtA3/hnHRU2kCOseM+20VbIuaBC9h/xgUCG+62sXds3i373RW2nJuK
jFBi/6hKUEIIcJGuf+JwL/H6/duEj90B8d3Vtf8Xp97gD5IRrOQ/PTPnYUsY
pK+Ai0T8ZNrdgZ2Fo5BEkCXjMIhUOMYnl/grr7ldCZkkJmtTZ+nsBcbt7m2A
vHtmjucNKZWcIkP4zE1cYMbqYqc9kGIomWtuppiVw1M4uT2KRxtv5eOn3poh
rVEroWMVLXUWG5ElBCp7Y0P5WMRfU4imyl7yMLTypRQPEbWppHeBZ7PC5WhT
kH4idZa+jLE/ff5WLKK0KgxiQLWzvfKsJE7BLXdM0CFvQI4b56JokgRpCD8I
m7LFXPutllKR1GeiHdrhRS5K1RDLaAis/cOoJjwiygpvQ/WI23hd57iq1VDS
8tPsCzVXbXhm9x4bNVdKaNsSfJVJ5TsU5kk7Fvem3u1V9SxeEXPSbcLnrnXj
bVlx1gfuPSV1Uf0tflTGL/FIv2A2IFnLPHX2PRs7wCSB8KWDfdRRQwlB2dOY
mRSfQlSznXTjmgWRFdPLg5iNYFaI7CqC9AfRYknUFm66MrWnfKwYOoyJLBBT
6vRqTX84FvLOFMuRRkkoXlfTUZ+lXmrhp1asTjx5EYtU22Lgoe0/VfXOcdkm
WA9hHB6qBD3frFNJN6viuyWra/I10LAgn9RZL+k12+WIYgBtzarZmmW3bjgQ
z5fRzibY/5pTPNf8qc9lm9TBdX4wb2AqwHBghBnfS9eiW25UGUZy+BKw/rr7
h2WeLbfwNMrziz8zIPQT23vZ5JCWletTh6ZLYOUPcqXbvf0RU0loOddtx9we
QIRlOhbO8dZzcyg8Yiky6RXlh8EcTvisWsrVOHmlwRZmCy/8uxZjX57zw834
ySwFxv9PT1cl8sZL1U+Lr22MCyiO7gtcaERWCUhDTD9tO+xEW9gSTtdyYaPJ
ulAI6JIdJk0DM1cAQKXsxe2ND8ejVuoz9K4BJ+1OPvtZnm7DRIcqmJPj6IpL
UqP8P3zmhhlEzlpx/UCxb4k3LiHZ1Q5TtPcerDDLI75cvn0CFQShy795v3Ro
wslGcGSlNPo7C5TngGg/0R5OlsAhUpTubKWcRAJeds66yPe12QbDVl4Tn6iA
TDHAXLmTCO2iCeEEW+Upp/KXR783xgvU1fc3q0wQ6muHPMqzg771RSCs4Utt
20xwPR74TygFV5KHoTk75K4sP/o5kHmSrcv+uMheF6F/ObkmnKf8sYTB17Pb
tW1A5In1bxhzZIJw5X+JZsI04U1MQs/nDyoKwLLHTZ2lLZ5bpJkmEq5Jo7rC
FpsoBPK4NChXbKl9vDeJSDezin6NjFx+R6LoZKb179srL4OwyingIbvLn/UO
cWUnLWuA8Y6zIPgnTpRO5IvFHEAVsJkokOcFk7QGmGmIbfA1ELCSvvNiqVOh
4uJs66fQjDsGtMgahu8i0dERIShieVwWiggKggIAUmBgnKKDcCJHkuwJzWce
lJnojTpOe+BeUtLPPPWVq5IDpmo1tVHCNCLIsClVI9qwInaDXfLue6iOtT5s
ow3ICcHjRD0tO0RRkKg1UaTRLvRoAJW72aOTiqgxqvlgs0SEdCSb14ZNyl2f
ZHQoDET8q3IjNRWhmd23qVSje4BRYqBdU+SngdOBvTRX9Zq+gcVZYcg7lOSv
kSWaqP531uBdL12wNSImPqaBtAZCIwQPtZRA26dUc0qYXFdxoBsvdrs99lLs
t80f9apHgS5j/tOwHfw5ItWCqR2wB8E9NVS4sK0GcvH4E8oInZFLqnn0XCTV
FQqtYrqYKG6lK3Tb9M4tTvp94xFZP32ZE/I96XbRnE30Y2SLBxqVOWcWvs0z
OlyTjL+amEBca5FsLYDb7yaikX06S52IAIKgI7dSLS/Hf6xagXKiwJ1BC6xt
rMtrLQbq+oAVJPscaDfR4CE+VTzG7mt0Zu+TQzqDM6Jy2i1wGFsoAN6QpqPq
k0QPWWgv3JSNyA1cEy4rULUuKgHep1tnSK/5ZNKHJrszR/wlBYvpmMHWB1sI
qLRfdocoZmyAjnmjkQnEUmBekIgdu+XH0EQWnfa+IwNW69M8vKYEP0MFlpx0
7KmetZHYNqJ5oQRZQLsvyDtuCx7btvZmkkOkZrc+Le+8iSEnDHtDrjZADAjh
6/JdLi0L3uXb/GLHuk7i0HjdupwIHNg1uFPFOiGJFyvw/CQvY7JfL3CvnPOx
KOSDywlxMihM802kc2jp9aShcZRm4QZy9fF4ZHkv+Xm539NH55xkJmvIlNiu
rTY7VbNLwpgYLMG8Y3YSCVpBs9HCeF6D2CG2+2jycjCPeK8ZZgKk7lD+EP+W
twimW721d3zoz7Y4b1VMiLCrqolwfxAtTpepagtWRe9o0pnEMmKiHyoYFKav
di+pQab9y+Pk7VgelF0DLIcMQZPxqbXJdKceMQj3/x0NigZiB614x3vnLYw7
WcPYt5iuhs9xFQx7dNFVkcHMjUuDvNdR/taNi6SHS8JFsUS2iMKBE2YltX/w
i0CPhiAagHvO2NlulFlpuTDAFW+Mwan4K/7HRNqN1mIeK0Sx/QPTI+bNdjC0
Qf9zua5QoYG/keQsh+YDeBMfbc3LeoaUj4DGNERt0qIaW8KHxo3+S7k8fLIL
XGrZdPO0z8h5ETTWJBjYXZJa/PLe7thJJ11LqUNiuy5jzOQW1jyirxdh1dll
Uc8ovC3gJ+TSvuFmnwKPxORLWICPr+wP9jJsFqjjEo/hyCDD4LWcLx4zN+Vj
Y285yPM51pRcGYap4lsNMYNxccgZgtZcKfS5p5gq/lMg3F/YkkP4t1UE5AiT
vem9NGXm+AxSfdBvJlPlU/YISgipwDBU/bdK3N5++JXUEtrPUVuUj4ywWbBd
lahh26+x5BqAinVvDlCde/pKYkftUti1bC24mqF0kHPTb6h/2t2BXD/F3eAb
5Jh+Zm4y9ulMAtQOgSaoS/AIUt3uKZAhleNwAjpLWc5JrST6mVYBGm/5lh5a
asqxHiFGLvnpkAgmZ973cVo9dZHNMkfncB2GXke6Vd9Tb4EnsnscnEP4j167
kc1PVyCMU5SdtgOhmN34St21IeAJJR1PvFDufE+HWROFwM3EmS63Bvc77LoO
A70VUI7aOtTb6QchZh97xDtx+qaFQUQ5QF2SW24Sxc+zAGOJ87Ug+a8dCoAe
OS2oeQUaDsIthlh4AZ635/DQUzeK+tHoOvnMvaDNvxSWabmAQHV6/mu60FEQ
mSpxD0H2PYvVK+QzhMDaNB9E7oPDqqs15GWXiLv0C8djSrk/Xuh+rPwUHdJj
6W0hXoI4kezCTgbrdkOEmxwoRtJSGHoXRXSsupL9xq9YDtjF1e7TA6iic4vZ
AaQqAVwPWpgelRmJHKfeOPc0JE30WM9u56b6hV4x39n+XbF46OZj1ijMm36a
UqD2oUiMj0QUbQv+BoCK6c+2u3IO6ux09vI+En3Y84udNvzeQlQYdR8AoYGm
QNsHG1EQm65m5ZMPnjTKBML2262SKInfV2wdn13hDgTW1f9bAmECZNvXaCiW
1KXDbwZM5GxXUlUoRI40W6m89OYK/1Gjpap3PNukvX6cuQNGnCHEdugvCltE
jYdOLma6CV6qlLWYamkRfg0bPB5it528JV4olz9ZrGZ/YoBGGTj8a+xcMCb2
fhR4/Xi97HLIHS4OPhsoyh1wd5KQqEMyE/3tr6aLztvnSWpOAbzqpiaylxB0
Ar8saICQxtBO8z/AVV+MBf5IYsg9WOXXFP7JI6824Kf5qrWfU7ozLbFjYrMj
RgnyFjEqw0e5dnGUl7JrxegLTrTy6+NRO72sfvy6erwoGJH0Hs/XywKj2dpr
GsPFz1zJtVZxHSy1pzeBF4jyvZFCpJVg8JWi3KbZF9AGPRn7TsE1SYBvm72m
SnZfE7mUkpaEv48wrL/PZVt5hwO+a+qaOGfAQoedURESDpTd1Nx8ofvDU0fM
Dp8+0UCzGKF1KFgRWQdnoDAnYH2RMUNzppMCnWLgsmOriCNcedjdoAZFzXw2
GEoXiD8IZv8U/YlYvBz61IfctK0IM8SbvfNwYeJH5emdruqnVz0IlMnavms+
R7u5op9DfLvu+tfgl6osT9wKpaDXuMqT2cILXScKM6Zq2Im00afv2C5vtQHd
FTxYAA36eNSywOShn2idhsWosU33egS451K3Eh9ia4riib70U84pJnGG3cht
dCyRd19716A1HG0sDwoHn2tJv3rGkGj4fsSj2fqOginRWNTp6sZ2Hj5Sn3WJ
yqR4gpKR6PUTzgvPkB9rwnicOc+pP7vd238JJ7AlWz15ivKwPtQpYxTQPMmM
Tq4ZBBWJagA7GMoGv+Ded3Za9FbT/szugV6XaGfx6NNzjGUqVADu736mO/Ni
eCi2ojEute51eee5AYc+QUqbhWIpEdhYu+XIgShj7dzGPJ+HvbKvEXQdA3Ke
sssCBIV5cC92x1FP/95se1HEy5739XdAB5kAgrkb58FVjyoXH2kvh1yzJ9Yx
7HxGv0sA9UpsHXGQmo+UrYpXad8DDPpBaB+zfy+9hPQ6SszLX475abann1fa
E5wI2Y5wsgnCBhiEautzQtl2VPBZluau5ehnoje7FrDod+cm1pkjsjM5SgAi
EWE9cyKNMu3ZKbN5FnTOPmdJOQk9CJCp2We5R0y+m8cEHSe9Muz+WuaHtunR
rYIyIxYzhM+8ExEj79y7WjmnD5G1VGhWP8lSOVnvDmMQmZ4wUNLdeWfkxc5b
c87Zy/W0VMhc25K2EmTVPQdAmlAQgD2WXpBFzWXojgXJaF5TruliUleRMLEJ
8fDBTTVeoydc0tuJrTLHzioa+DK0oUgzjztO6OSrHf67rb7SXMkNZ1qw1Ak9
xkRtNr1SSQo3d3NSoszXjvh8YwwfLA6F2fB5WTv1LQZRkKNtyG0mlRnxZHAS
ZXfRmRsdeL1/YeUyop8MQUaseU06CA6/sswOCvM2IOE4Z1xY2XxcQZq6bzLz
j3jOw0pwC0FRY61TNJyTXWMNzRE50R+jahZRxMVpWAcRwxcv/ERx/o5B7MzF
sAoNiqKgXhWBgr5785kVtGwbDkmwKqUg5ShHk6/FWkJfKvfdSg5TNxj3HOxo
QynG+nwQvE8DYGl7SMlrm1f+RSweRla8KognECiTJ+GtUkkuxxJ3OQm9HG5E
GnFBEIGRubm02HtgLudXkIItarZIWFCOtZfnyyexZmX9Y1b6Rz9G1uJXgQDz
FQ0mZj+H4ZkDV+zHGCyBuHSKbby+RiHobrdHTlETcEM9g29Y7DneHwQoQa3l
aENFxpUW/EVsSVUbD57+4pVZBThaMhHu+ECMmY961FPIf2mHRL104Rcvhgof
XRJH/qzr9YdmsRVZmTZ0o1/af1e4DNnhen/5CfOseCWk2+cc1BMpHuM5OloV
Emram6MYXJHdkoxRQQNwL6P5UJJabGv3/X6ED2kLArsrqnZlI/Nu3Oe+2GVx
Q4/9D92pLkfJaO8S0VfJ9pBbD+q0Rh502Lgv0juZhZMeDSgMRKghuXaMMkjZ
U7IITUp5zkTwIoP0VzSR+v2R2bh+ww82ZD0oW4WluhTFX90ULF70j+Rrhzkk
a7giw+qofGqdHswWAiar6PuRBUdNIdWYuxLZsderlxkeFdTxW7DaIow8zhSL
WH/4BEHtSz4iwFvPhFPSU7SK1egEJeE1mshZG7NRZP0Puhmx+DmWtveeKIJv
7sD+3u1ZHKn9D4bX2R9D01yLZ9+tbu6vzhQu/ZZswWT8elM5Qb/Wp3bMUtzr
rHO6odSE8JwUS6Ib72A/B5CFPYmA3iAC8Yt1R/E/IDmvu4HqI4wst4xR+DtG
AfwRQ0RUXnVbzmLRyEe2EBEk50DY9nmLxCBguMS2OIu6eeDiTPX8NozOf0vd
QlWCkHllnvrr0hfswlSbmE5oRWs8Fj43Ziv2QdlPi1+HYCuDrEGivdI3+3wl
8dzpxZG6qyYnaJip5JR6pvQtztZb9mte1ShmG1rl5m+eLE0bd0cs8XxgKfnf
lHvz/IGnSrbFU3snPIv2fsCf4EIfDc8CLXOb/IOkeLV5sZqsLB5dSTNw41Iy
rumj1M/OMj9oII/tSQCEqYxLWXNeyDTJV58ph1KZ9tJEfxb2TTXHkwqkyo47
0hly+x0OiWBIj0bM2zZV1ki7HUPPX8dY8ry/ZuhvkwLeJlRhCeUy/MmdGvLu
in7ctCMoXMBQGE4PsdPsxg/8arud/60K6/TZTozDrS8knsuGXT/oBWL8WaOg
Rlm39BVUTPH5aVbgaFY/BTzLPPLhY3+SC5UZ28OwVdaSnjjECV1T1fOsKdq2
SvzghZVqTuvSrtfQLnkOvJVmEgXbxaIXNncFWMFoSecSiZqwf2bNo83A7RDo
kKlXD96/O6Ie3n6UIZydFBDzz2dZqM+LO2y0tfzXcSe1e37JLV+lx1XmGaFr
HqBUtJoOCivazwld5dqM4RBS0Y0Mw7PsUwZQsaR9tK0kAYookG67S2IW/4at
KvSvw3kTlrP/LZnZrPP2Wfh605pb6FhHuas4yLJ2lvl1yzU13dx9abShr8PA
QUfzk5gD4duQQP55L1Fde5CN5LIcEbNiWcw/nBckKk/gA6S45Rxy2e/DuJJV
1GluaPtz+t5iucuaysTQGnaM2qv4qwwmtT2oz+niuQZjnJayi1J+GRx0HlT8
qKUIhArit1V1lyjseyaLiMQpx/8xXaHsszA4gd1y6zVoT96VgecsQBZFupOh
f5T7NUhTMA1w9XL7/KqHgs/XZZGj7aC6wTFyyVLB23TLKseUa26PRxnRtI9F
RCqAeR/xXgGYWh+T2crrYmFs/Num89ZqkG1kK4CmC0Po7mJwc+5OLI5yInDM
46MRMpvwtK5z0u9pllMcP/vSby9eetl6CjO9mjOEMRvwzqVPHGmjwKxE0/eH
aQDoZjZQtAT5nD3MTZjTMtxcVEV+uEb57cU5WH1uvmlXkc/WpSlcST0gQ91D
BxE/Fnt8VpTBGKe2dBZaiivFotZAvY0zu5/CjNMPF5sjfH+9S6NBhoK43jl6
kIh4UPTWIhvzKXNUd4556sU8KlChHIeNuvk6+tSq+0yXANhrMef97RH8V3qQ
sT8ikAgHh0q2Gx8UMFCLg/R2VspTSmJ1cDJ7sf4geKyhQJnOHkL5QqpZRAha
QaCQ4ns3/ZhICaAevXz8pDq+y4fleVV0KLafsnNMlkz/i0zW+57nfoFTOt80
IP/XYl6Qupgy67Fpt5+tqx+3L7JOO0FCGQzS22hmeHvjZqHlIiIQylVFpPQa
kWYbVmrWm1P+UU5m+CZa57uGaVwMw6p6copjKojW3mpOvBNKQe0c58fqaX2/
YiAdJL9E3ckd/Op0LeKA5yV8ChRMQJ7ivO+F4eYfsyWzcz2cYNgJDaloocyx
ma/YWD3Xp+G6xZHGsmkm+BXH6kAUD38qtKotdOAXiglJG+jSbS19+oeFX4zi
Ea2zIFcq3b4ds48EmQYXvjIF8CMFf7Bv/1jIz1q/zD/9FKNYnX501wAttKk/
CHBVSMeO1njbBpBETAAtNZV3FGcZU+/cZV4aTLsOwKVQEV/W2MZ4OSUOMEui
Rej7QkXhDhAfSGf2/7bCFljGc8Oc46pwJuT6HQeUHTGUJ+XgKO6Gagtm/Lit
X8r/uvjR7CSMy+P3Ccj4RciLsTmRyjh58b2/ah+DDN41gYYe/7w3yior7p7t
RaTLaj9/4oGl0EgqRarzHQSVHfm+CaDElOuf4ZQqCR+QUrNLP64Pp2vmzC88
SO4z8K1XHcRiO691U7wcnxT0d2dT8R7hmS2y+fd9i/ZpwuPsSVHgY9TG2l7N
c94UwQZuDhMMjZIoMtX/49pRNB/c/90kykUHZuOvx0H6rjcUYoEOa1aZyxQ9
OeQl4Z3BgoC/Bq0Wn/FbnuxnrqGlUczOrQ/LZLiH8kHoVBPVPOqWvmQAI1ek
B8mRXFmkVdJQaj6C8jvAo7mc2ybUE3/4rn9Yr8Htsa8N97abMBDIvMl1ljNm
haDgIJ1AvEKJHKYXDn9beUYQqcI5En71G5QRuZQ4cG7bItB9vDFQV3QBV9ob
poOGWo/ErjkqRZJcOB6sU77CaT4yW5yQ+g4bwH029p3iXzn57hQn6DL7Gvql
t/d3VGfDe3cTMMbxlNyTZJhFMDhycgGy+jnZH3JAjx1awcASQaiolj1JWTPc
YvYLxnVbtMO6EnMqw1tZRTDCA8wYBqN5sIt7MeZB6m9qeGVoCI9Uw+S7lzVS
3uNawe5yk+uGJZzJ6lDbRXAseoFzKasPJYl4GA8RkOCPNOfzWKnuqkCBSzIz
aZl3ZOrAlJ1enEkpY1yFnfZjtehTZ8MFwYx+HoYySzrVTh5nMbY3XpKVSxGw
2aoe1fOsZt6efTuzDGo3n3DJwBMrFLPqKHyZESVNcLXCsM2EVF1KyT9AzLHU
YPa+oXWnHNPGR1oXIGVyf375O6cbxDJtBr3xl9LeWEPkdHi1Ewtv2RZrF6kU
+jPhz6rR+AcZCU86CexOOHsVDQxhLdf0QMWrZwj6dueEE8eitH7Vq/jXTNOJ
2vwL5uVBivJweYCjBm/l1MZO87VhsWv2Otv09vN0f0l7/KvsyazY/uTTLIbn
QLM0ZDye3mcKdFuq/knrB7dC7M6P3At4QYtxTEEyMg1yr9KfdF8NN6D8H//S
oAdRdddmV2IAyUfg28g7253YFrGogMyk4d9NoXN7OBtfZ5h5MSSJWvs/YaNL
cS/GKwIuOEqbRrNpVKRgBgKhFLgtx0IjcZ1rV14YMdL7d9s+PFHSgXGuxAfe
IC1/wlOQg8WdS4nMkfPkeAXt9h5uzT2JwGGtG/j03Z5ZjpaBk8ljmpa2frNW
h9tjHYb+NLHB1Ey/PUntufgF4xclpodrcK8Ud3f1oiDYkNZ9mvzj5Kx95r2b
RyvC3e1AP1XyvXS9ifWZu2a+hwUj2XAgKf14ZFNjeK9YV+CxEiSFB5na4Q/b
TmwFnvFQZrj5bv0YDxy/aXZVljXdB9exkAM4uTHsMvqJorff044niLOnMsAM
lCkpKjW+QX3LpJ3Qg0eSC6Vr1myHT/vWvp2NCyQaYCQf81xMofr9SG+j700c
O9Bnxkhs9SE+Mw4dNmrCTxQhDTuA2ZQLRCQ8Ha9Vd6qwzmbcPNonDHjBHfYr
xcEdxUJ63Sihr29KxRFduUV9/0jctZP+bcFPwzzuxvZV8cg2IN7nsiDXDiGj
NnjmV6rINUewJUOIfkut19+ZbAf0bwVhvV17qs8DUVwpp6Nv4s1fuU6vhszk
b78o7Vz4xJxVo/YddBiHys+4Z9E3DKy8sBX+ATRp/HQlfTKmoZi7UOqSiNUC
j2QV+xLVZ7NPtdZwK3nJqfiNkjw7P3LnzCviJ812HMCQTyr18G6yL2tIPqa5
QkRyY/ZuQUqyL1oKnnOpKBHO8XuByWIwzmZLJn+bONv3Bd6++Z7E94C2VggY
5JQtWUa08NsS/yQSXOebzWar6OtYPSM35E0iq+F/l94v2MBM6uTiH5VyJaM8
9WcoOI1fWSNwDu3ibjL0bGBWN35ijc8jGUkR20W/staGgvsfdyb3WKRhVWai
X+5gtjeLzk8kHSEMDtCyXRbOKAHLNvFVYGP/FsVwkcn4mmFkCYfA3vvwj1X6
amPR1m3/6TtqsnGKo4HWlhlExmhFmAYmE3IeVd4MRD8tZCnTFM+1JwsagbLx
MoSgAlBFuKVOFxjc7uW+n93X8kIXBbhUEIvbCpfo9AfJWqfPs93wbZE8Odaj
zUxQa8yCJy1s45o9Rc5HRZd01z00wqSP1bTowXKxCrcdeDVNxMpFV5g5DJah
rZd7uDbcAVU3oAhxvUJoPDFnUocS+jn08nLzkRFUJMKqoNBYku+E8fNJrjMf
VWl5rxFWAWVZrR+kFJc3jYME5dLgHBsOUrqUlTZUFB1VhI6VgRO0vHeVBk2+
6gWq9M7TaqnUUGMFb7bEpwIhsexuUaO+Vki5cibke5u6nKm9xTkbgqhjId0+
+nvp4pjO/90afjrG07eIgzb66IhaK8CBKmG/7Of8Yu4KN6QqVHHnV4u979wZ
D7KxE/SLdZM4lgNRr6okFv4yYwKerHcBaD4srF/TafzkxXYJlz21UUjhoPBy
r6aIaB0k/l195pBwt7ADpF942TKv0GxXBQGRF4mwXLiDPpGJ49wTwDej4OSr
0gZ5biBkgcw1mtDjkTRESypM9S4v0e2DGUoJwKT2IgUrfnn8eaOFHtT6UgTq
emptDJLJZ/9hBSmEvE4hfp15EhvdzDq2c1tEj6Xy7IDs+MY0ubiExDfxfN/E
CgA7Mb3ZaTJh/nFSAtcjJOHcvromlCfDE/v6WPTpS/SXm4rkluz9GNPdKiVJ
CoCM6qQqh8nhZ+4i2QTUK0eWlUkwcDJb4MK5Z7T2mgxVHcPDlUM62VvcgI63
BxJav1loI8XQhK/ACL3dQuzjMS8wdV+Tr+M9rNeL0w29mnXJSeFlp40QztST
U8kCdvZlQ8TXUOtVU+nlwL1+aHPjsRvqgqe5OBMb4VLna4xSIwZjsmzdBZa/
74q1l1LpTs9rnqfP4TzIaa1wfDaFUQR4B0OR5Y9Kq16dleQ7xPKI4qKImMuM
geCE21sytx/mqO6mWMf62BrroBj1G8wVbP6tB5rXXyPWTTzCHS7hOU+RdDV1
vX9zmiDXi6UQ9SgURXLIgBvTCcJGeSa7+1+h4zOxdx38kNKyKxVoo/jkXAOC
yIvX9z7h9hNOxKa/MziyQVNAVRHtZnH0OvnE0phFqVNZPyF9ARXksvJpr9Ks
UezPXEHzDQCjB4rvTHyGgZmioZD8H03ryM26Rlcjp1jIHQWNlJsDdPv6bhPw
AS1Bfq3VuYWJSw1Q1qfnGla7MrGqxf7F/+PgvbUIeI+P71bGeT964RX4nzLb
g4HHpLwqz6K36zy7zn1RaZ2+TjlYLYPtQ3D5P640u2WfO7/Q86hDk6s/sCT5
gL45JqsTDamAKWJn8cmV8MUAt05fin6jxq4TNdMi1WT9xZhOvEnpjgHfAm0c
ImbEDLnwMadoNSQbvXXyV2t/eQMcULVB7NDue+3LwOnpLWqWxJEdYlXoDK3Y
Aw1IDNYZ0wtdh7KfT89Tlfmqvo3E/7CKlX71mmrSUhSq14nqYDdBP+e3alv2
h/mTm61WeRzCEthF8dQ5UEax7pfynComzfLej/j2nzMNTlJ5SEebO1Yvt98y
5d41WM2mwAgiI/lgrYA+OTmYMXj8P/42bw+RStDTR27oW2XzYuLvu2AfUG3o
lHVvE06ZkRhw8P+Hag4VTEx3+M1MCyMzWgpjgwr4yTVwHPWKtQrjt+1eM9WT
rhNSRi2PM5Z6mCGOagtsVufw0COmOHm4bN6K/RpE0DkjrKlPrgIFyfmojIPp
0Yx++zqMdoa197TV0aUbbgerSXyJrSc5OLJ9j5ZRWpkkJvnGWEyT9iluy/J5
5K+hSYiOgdO4KPyBQ1rUbYCKl+IKCNcPTGT/xBKZw67VJ7bT15f/PgaP8L74
PeA8gpXlVounfbKwCWU7jmFIwziAhUJxqi+2/VgdDNwATyISvt38/AofQDMO
6025EZUPVGgF+1szyHU4b4UlYrAe/XQDd2FOnD2xhSGPMQqYPx6H2RVtTjwK
0cmssyeAeebQBGJMyDEPNvS9IB0lUHaFRkHN9SbTmrGsfkLz0rrSaIKGUl8+
UMqgGVTsrze2LQmxDd0IG9Cf0x2UgghamniYGEQBfPkj0KRHm9JUbQALxhv6
oOaml1FYGpyZEJdHVME6K5MX0U241cftZzVVYdiMufBdR/TxlLVd9Rts39iD
tnCfacTPWbOt6sZgAgxpXOBBr8TwuuRtJ3+SNedBjnNpSy8xpYSD8LNaKsuD
osmA+5KPrZThnPkhaaPo9PFzq0LJsPhh9hW2rL+u48LXoPkjkvBVuQq4bSA1
7qkaTusF05aCl9RNU+haj0it6Apuy1X7qgYDiyzfsQEKJVhoAzA+wC5el5cN
8kFT0Dc0kP4IjS5X5mYpNxXG3/QZIu5cTC4BrnaXQPdBIUyoy1UdXRDcM6oM
YlAwNYcuS+qxRigXmZvnehyirChhi79LKQoaADjKRta+sWfI+XKZIu8ZGcBq
Ig7xmps4vUUfVrEl6AB+4Vy7elKcC7d3PZtpxZnp7eO8aIz9FQU/ZeWOeYyO
TtLcmS3vpLLRJ/Os4RiuUfuf/iEIqOZZtw6V+wvt7sP0soy1+dcdexl8tnBl
cgyqz1HiVFuJI+7CTWVV9r5imUWnml7m0KbVlxo7/JVl79F7clr1mh9OtFnZ
/aYlvA4CK0ItymrmClOCEwwBKa913PbRP+MIRlcqyYHpaRFrXxWczgO2O6oK
SbB4FXAd8rofAhqFQ5Y7V3wfsA927gOgQ576dPsx4GFqQknEmuRRh22oRIrF
qOX32PXJ7VvpcBxOJG20zYWrpfOTj3TGDRQ9ugSjtjdU+3gE8WrpefJWctUS
GGeCYL2IWSx8KHNftj/wZ9yhfMTj4rrx/RtAwc9SwhGcuq2DNZB1Xky2Jgfp
ox4Ctrz/OqdvqOnbHd7nc1n/qn8hRexFvcH+r+JA6zxaB2UeJQxI3E0jPs0d
3Rx7PoYZ0QBESK9QkLyoEdhxpj9G95HKHNyv38cXineAg9qaZ0EmhFpy8k96
/Q3SIrAcgLMuzpPORaKNyVu4AE/Ed8RF/am4IHAqfgyRDkfz74LW0719YGYs
g5nps62zXjLumP06FeUonaTXpWIQJVKRMnmOz+VIgTU6EInCa08DD99KHOhd
ENcIkMGaSGvNgyjtUIIMDkR34OTTGaxXfQFpq1Vx2fmOICiQyn1wjmNFXQRe
jgQxOtHh+YKdZwm6wOHsGjjx28rX8gLrQf6uvf8RMdBOABY9roQyElD0Px/s
Ynt5qn6kPXrN56Cq1PWFuj5TqprRLk8N7QniHxjLNFV51ruk776Ec7Tb6I0G
eGYF+eA9mdPoXBY9Wp2pJqfcBL0ghEpzNUia54quHE32PqU4dcrG+yz5p0rt
DCuEt9AyvydDXlLaNFN45FDTeASjsyDHLjpnWukMiCw11ovj0IvXrPuSbn3t
Cak1j9yhbcAGMyUcg0kpEsqH/BLdZBgdo6O736/sr6bEwsdArDk9DSRgQVMT
LwyEVTtaMaX/pPvNgPnsJ3RZcjTwbzmO+bByTUn1fgwmsoeaLEO7qr7iQNnw
6+Rt5jBkQ5Uo3U8pLnJY7wOsSR3cuLrcewZ2uXbXcCmLBqFlQZzoQ5LuOqPd
rvEhd7z/X4hMqF7ALWqS+DxPmopRQkTtr134ahefXG0se8DOlNRJb6yXe8L3
LFADT1qGO5KbGfi7RMrjLO9fjJZfxPRz9WzsaLUXBu7QeFHyemAb7BWwNIN5
zUySB7WdV5Am/HMQoL4jQopcJHywHFtLFmX19D0e7x0EBi18pznmKNGX8KsO
weNPcJvPyxASgdJWJJS/YJaUOHcQa9qpZbVqDS12vDwzUckj38qujt9OD3B2
3/+yOmYEwKhC6gVj8rMHQWQeXR0vJAzu87QCWy6rwLdvEiHpakvHcSe0b1FS
wioQ5Mq64+eOOpj/bSg++2z51wYFJNoz++KMO8c7CFQLYftvwl2gfo3uzv9v
tmyC5bifHbRmM5UfjN7fGXOlN2fQtWj27kG9j+CzmybbPa9qnroSI3bUOWpu
7UhyCvFi84kUzKW+X95MZM577nZuserLVYGEr1wS7QFwVgGZDVk4kQ0rvMew
VRccV/qSN8bDDuy77eiyPyh6FKkZhsoWhbCR1q9iiF5xSqlzYTL9/3pByJWk
rLi909RmI4FTSOwC6Eg9K33YkFb9v0mAiAhzGJA/ezrl3FFQG0BSCjz7Ymln
xSvz/SQaySUQU+RpmWM9fr2bv5DTC2BcDUZu7LbAWGjnS8Xo+eJPueZoXmkW
fO2sOx/HhhmZYWh4hIdVuSKrTHN3SaZ3ud71SB/gg+dG++BFX8AyP50UJeNo
+v/k3RxfiegH6+0h8JRSCBc37ueisQtb/Yz8mqKgmeBB49oclVWWb9rROhKO
T2O6T/utxf3iKjgdGJooaSY7c64bGiQRQFD/CwcmWZLlTr/quPmkpzH3TbMz
BjCTZO30gbK01+o8qd63TRT9IxmUKNaBGqmmnT08NSu1USJ47/4eQ9Qr+gF0
aTYE3eF/Oj9ASx29XbCrPiceYJrbXEdX1wdcu5K0WWsVigWo55Kc1HM5osf3
IpiZJJWn+3XbEaJd/0O+JB5XDlIj6EX1T0h9Azwhj6DzD5WfDggE98JfU5wj
FGaCPAncNdmcZQUFh+uQm1sw6jV4uJGxJdIlI4UXKK0+NbHzn6xcoEbOQFlg
O42PErIAa3x47MyHlyRVf0MZeDNUyGlSkgKPDyZ7bcDMbGlYuse7tW5o42z4
sw23/v3j5nJXoPBoW9Ie09eqbyruT1kE6NsldwvpdPG1MYDhcHeVdrUPCUlU
OkjUmcIqGLNG0Sv5NLQ/iZXrMzKQWC+OSlkzB8HWHhFbZvEZV1blIAkn1dRi
mAj13a9UvKIhPI4vODw5L2P4qHzpNFRM7ShCwcH20wcSV4yUz7UzGKdpUSLu
Crw9zkeJJQbbqjBtnKgU8glDPVWl5QeXygT7YhLlaMF/6PhARAJDsDIBrw9Y
3lhCnclFhEiPK7XQ5Xr0PFjygaRHnuL9Imf16/9GDAPCupTkrpHq7GVXbOgw
LKtzNIHAqm69V3jplUixJm4jp+/dbUCmlV1n1BR0NrzcPYGuPoSa4E4gnx5u
/1HpyyUqbfc5MF7srkpex4o4PSaab2CQ35opwRHucr21owEDOA9fgr5VCgP7
69u51g1f1snllnRjWmu5u4xRJUe8Tyx86VIzmxT+Dd9Ln5SImWoVivoXWN3h
Nxt2K3RdZD7nKywdEOAWGhILLJ413ADdTrjRNCytlDMXZbCAE3wsoi6XwBQZ
+iceutmS3hvYsEruBET3p/0cNpHzHV67AOsEd2NsQn2KoHOOTuHEMY6GdvxX
7soyqU96AJ1NmYpvWvW9hhVWQuqgh076rzG6HVUsoWExB60iLzoLIWWXCxUZ
rssdyVib8iUFU9PuIaJCVhsdQs0Nh0aKWqfjmYQjMuTUxlFPymqgljZID4XI
fY2niDARNHelMjD6l4ow5qIQo6Vth4S94Z9RQyU5hG99rQfeuBphWv5+Vyhd
AyGjowBzsV6B8+t77HzjhPtqFTYaEKRAFFv+BVOkKGdmgMY6uGjQVSwF/HJF
+FK6iM+yUYke2CitsCqqBB36y7iZAdudF7Zh7TxPdO/cH0GhBhnC+zaM8iEO
kqKd1hweQK3RsdbyKMI2k/Br5oDBqPsK/d7Lpi0QyMsW6Aeq9aXs8VGX8B60
gg1+HnU6Zq8jjHzn+tLvDOlDpO02XSceII6fD428bC9V2q01DFBR0esUzWKj
nGE8tq38vhU+S4nN5jAbh3pN1L3fH2h5uThyyO86R9trouRHY4UIvbHTpQ/p
KUK/y1LbuKxd895lmCd2h4SAd1HrsUQGGEdH/2vk/m5XelO35ZRkyCJsZ9Tp
L05DBZSsQShKE359cl9u7qnpzfPbLBe1qFBePi5moP89UmL4XBEvVFSzM+8d
0JrYiv0QLMhFdjxpzzCZI86PQUWdP3/wedI3ZkvzXwfpWffnIQcJESe05RPW
g1Ej2Rd7dq3gRb7hIH3RQkNO/wlPBiKJEeqSRJmqYCZW8YauUIuksnEWlPSQ
8DwgKiSbRVjY/twD9NljOB8M+uHIeK3ERM5TjUkJ7yJMnyhTCCuB/bz8rIJ7
ZQzaDmKzpOyHbMG68Ws5/gHZuUTYEeMtvMiBaClUe/+iOPJxS+TRRpJx3idY
fY/RG1AsoXEsLYWViftEJoltmwV5E5pmOTmWnKmfvvCd8Zf8n4QaDXYEt1Bl
CpQq02fnCYVksRszBGW3x/oZ9nHi3vJCLwjGcF9cu+oOuF/luA7DZtM14W/r
/UtldmIrDJQg3l9VxhcYBtzgLO+iJRlZDdiSUJRMhRdWVQJqBz+r5VLWZHdp
OQmJ+NyM3XxwnayjGYsYK8t0bEx2jOTgVdXn6iMAd6eSLgr4lyyp9ELcLA7h
nSTCnXHsMgana3bDHETnv9MOtYH2eO3YeYz9f93z1qSAGPVuWgBpVOsPCqwp
xDKuwtrdACkXH+AtKYRslD4aolCdHKi/bums/w8Zxku+DZVty3FezZZGnXPI
owuh+F1Xu34ai8F/xtKZeehVMVzsQeoe4+flIBDUaEHJPXe+KUMjxYvX4n7P
PZwu49gpILl2FlhGitmfgly3bqWY3tv8+jF0XTIiDxq43slLjPt5vs5+nnSp
qXyQ/1Kwm68D9NSahDbJpCX/ZwhFxMxMqsuATkA7AjVK6Ot50IefQ4fBM1Ip
bHLq8h0ettrR42SL7xkjkC9p6v/XVPi/hCuQ/kBOMtf8ZSg8+zlyMB4jsWFA
/uIU26XgMFi4Uy5auoQORWAOyiiqeICgHN+GUSfQX6uY6qQgrjauReJEtW/a
FtFHRPNJYY4SD9o0WFWjidvPBmN8an9mz4I81S2kVlHhYLN0BdDzyqnJ/A4M
7vUkV1/rjzJy4J2VIis4uSMAEPOVtm23JbovL9QSL9NBefXynLXFlDUsoGi8
M9nhWOMZl7cVRev+PFD4WTHKcHjTh6JdNJixNZ1MDusl+57uWn6EvIMf7oyD
H6yTSTBQCTlgvfL1NjwpmrxmnzsRVDk+kNizJoAgJn7GasyRdnEdIkYmYaCv
tkZWQyR7qjnR5RlYbRV7tsNr2ZDwRqcP/MaZI5H/YO8hTOb6fY9grtL01SjP
+8pBavS+kWdEyAf9vdwc7gD6T9Ir+2KZ8r60WVbimyBX6RZLNOPjgJ0rET05
PZCn3Q97HBaY5S0HJ5tpBkuRFIZxZblZsPC61+zcrdzdLlGv3MrEAmLyHlH0
nzxJdJ+NUQ7NHJA+wn1z7h9Na9UQ4wJdfMWKqDY23zjOmGuBjSpyTiPfAWU9
SEtu0FZztR/rnZZ49QEbGrFin3wJFLvo2tZL2Vn6+H4dLz8AmWbgi6oGIZWj
Ji24jobvnCp5Rl6PGckfr78ZClX8y8jg/38FLKiR5yohy7D4KM2FWz1R/pyV
5LPAkEB8JOdYyLSEZIq81KSOwEtffnXxrG+MCp0GI2Sr9XgkG77AFJXFN0mQ
ey3bszOE5ZvsWUUsFPbM/Zsru8g7E9c2zq3EYbyG77RCXCo55FZm+AVEf7Sy
Y5zOf0NhJIC0+Qm34A3u2oaGxVLl0tITQnQeThno3x1/YmGop2tB4jgJC6z/
MdWglD0Xs6onXbDBeTDIqLqPxYWYoAjHv1ex0guyulBut1IkXsI5yxRBTX0H
iUXXs5FEIl7amjawucm0W1G/bLoPchfRid+aa2e57iTFZBYPRs+K4DchoCMu
y7+qqevUUzccd28QXdJsFCrDQvjpTUSQPSaDCi6Xxjp+VvQFZIIX4H1d+XKM
6a13VAgNMKvK4pjmfP14GzAYM6lkgYKDfs4yNVlsbHd3Uxu/l9O35lZPaLsm
YXAoaHGJAbYDB1p1b6ZhYPFKS0ZRN0ZMxHE8jTLZ1kpwUsM0JgryXBHPyBXq
SA+sOF5SK2X+wSZUNv11TP0TRK1NN/dFO0jyLVxNiYajKOKZgLr2Skwsj7Jg
2HUGwwWnJi4h9RY1u2U4wYR59XXRjgMz9nUFxsKagpPcKGusdR0vbSIbKbM4
YDd8vXHx8aL0dYHEp9BkSUJtu/IUpkvUv3RvQENgoiZeJZshEY6HbluswmXw
k0xf6MQ9UCXj0NovGjzhoBnv8/w+L67v8+CbOdyya3DVTX8PxBuYSRFh6DUo
fyYGqPauaNYi738NtZVDtGVoYf4ArydYXtdTrcfT5R3pETzNhoNqP2ARrt8U
3FCzRo4iskMxV35UXWiUFi2y3Yl9eLVBlnhlbc7tEJfjLizi48tWLUYHt+ja
AV0ZW01O1Ftxa2WXbzHDEkIhgPpCtxSITDEAENgMHbASL0qacHXSEpUUARyH
qjKaLubLRJHFl3Dpsu9Z53VZGPJ+nlY9WAnsU/HOhAQdRf6ptGK/tUMu03U4
OUt+b+V95Go6kpRIyKJndPosWNFbl5nZ6WVNu5I5hAr6O/q7jkV7pUIJiUkp
fSTfBpNeSiYwECMeVQonNvR9+bxuI73f0+GqeZfyoT1/WOKtEItieo6BdTPI
rzSk7TdCkXj986w/7Xywrt5vggpyM+yQLR6BtZaDqSisCa0ZfOL/95QIC45H
IMpM8vjwlM0HvVhGpmNGDgMrFMLXOsyRBaXU2D+t47dRwOU0KYpIYusJdPOk
HGByhdZvwQjmyCCrbzQuRkxTV+JE7VzFPMJyHyZMuPGDzHStVNJEaVVG93Pw
AxiwM5oH5wZVyYlZKhNoYAYFDZFN6mIpwvTcT0SEVZZxrKXstRnBt8xUJE0e
Bn8swkdpJpmP05VFuwEsn6cOgwhtkOa9WTWNzofXoxFMBP//QoWeNVrhcTwk
2Ui6vOBfyQCPl9OqT/sGuaIroAj5vgslhLyTRdYonshKpeTt1dp5NsZyzjzK
iJ6sw/dkJTrGsGf+0JEXFu4K8AiCgCP44eHN6xUvC02z232gRTsUa+OGfyU7
7MYoPWxyDhkxuOTP539WVGnEAOpQUNzqtSfjcfxtIY4KKDHx0n+ez3xuX42o
sY0DPJRCVdUVq0gnHEqUB4RL3c0xY1WMwioeL/EFAOjR/7Sc/QYnnNI6AOKJ
qWJfqBN9T+TtlVpKbEi8QgJzDpypsmkDFf7LEuY72UcwmlSTQKlPqccfZqT2
dUEv4cLmrwKvKCoWZpAU9GnW5gdP2JMbj944ZJEAqrxcio6uHUNqiLWg/hK6
1Q5uuRq5eQF6rjz4mgqkHflED2Rdqf5XcOvOjWi/ORanIwJThflj6XJVlJUf
Ib9aw1v0ZES9uRXI7BgVJVMqRy2ZP+E38evB7RuHIv7a4bS6JEZ24PCOBUvo
UG4tvLBjyV7FjXd3qJp2AEqLk9x79GRNmSjTcR7UFLr2ZwOuk4NBETPJolEq
MwLhy812Le10JYus744M5aQLiu8G1GrQYss6Nha8kwOlBvisUWCbZilZYBQs
kTkhuzEK9z8ERBGMFyeHOZJJhgcSZy1Q1igYd13NFZ++ocw399c6m79Qevg7
nAxeVRprfuAeOusWqKnulwIOonYZZP+eDi67iZ3pMj+sBlpkHwE4gLJdoj20
O5eN3529iZOuL7tYeVo+/Ay8bH/GnPkQf3EqTs+/RM7vGBmKlzXRu2pqHBPJ
sYZkcdEhhCDmfETZ1xJC6aRmNvjpz5JtvaIkeMg/fd/aFK//9ZjF2QQ47uZy
ElWzHkPEM6MkGL8dp7CBujB4hGgmjsrL+3ps9gSo+NsFnfCv4dz9Zbo4R3Eg
Vw7i5xuOLGpx6KPJLQvSduggqtxGuJpT0DiQ7pZWgT95CqKkeW9x/kbipJ+V
2nX68PeSDqRgHatyjVdUs4jA0gol28NxQict2B9kdZHmgT1bh8aIYYOe9mtI
lLhA87gPRkIY3ufqo7fnKfF15JuoRWXSkuPknyZ7JG8Oj3fV54ICHbt8HF95
d+qH+f92b9SHUV+szsBMOybByWqq64PLKvEOgUyYB4mv6014Dr+Ht3Gj9EJD
Z5se31yhw2Z+befflSIinaoPAYE+7UyNYOsxCW65D3hiIacAW9R85V+018Qa
biQTRUW2OvZ6bHJcarpM0sqsv9ERFjimxJX/yg1wzs0+DMJ5KaDdBrLzhJBA
fnRpuFZlkg/WESY9DtOZTafjcOSeFXY6mxnppQpYQPkgr6CaryyM03E6EDdD
uDK3gtSy5jI3Cf7STtrmGHxX9P1i9Z6LWagqZSEc+mQsqakwM7Hj9P/2QcOp
PxM+SscVq9mP1S5iPMOpir2TVK2G2xZnwL2t/PrZdgV7VDl3USHCm/I726uH
4TNpnorqWyWibCbksS1AQvIVo/QRFt6gnUa6OkwJdJO9l3ltq/5rxS3qyjT/
QhydDTMBLvReMNsAckvagew7fpxp6BlMlFCAKntORI7DzLUhcQRgMM5GjbP7
E04v7Nam4+GXn+79HyiMpmlK4ws2GP6yGpvswgI3s8IrshvpSTqZNZOfdfO+
biOjSQEKIjBPhygbDq7FeRpKKw83fe86UfPMLkiEa1+fNprnZ8CUsPRcfdil
LdEGsCz9DKSanUNvtb6/yj5BzRhbss6s9h7O+56DmtAE7yj+eyjvG8vAEgTg
QLdO0Dt3nZYRGwsQFifv1j0ppm7BNiFJiDUBpZ5jh6q4TOMVA7OnelGZh64O
/8fxevr262n1OYg2a/CiQwbytbAnymeRDfJiVBMjHscK5EdSwkzyDS6qI41K
KGPnhRqGWjWqSxTUcvNr9UWZlKURliOue1BcgddxrnkTHz8mTnwwBWa4J1H3
LpNsDMunS3/oE9y1cQMw8PFCY2L8M4BmIK/DDePy7FBitsJLavasH45VnKbX
Wy4ArJWiHIfx6jigNfTHHBNZSfd/JP4RqGkFc9pXXQ6LyRlnluao8Lme53LR
kuLDg43Akr9zKZeXPRxH6sJOjPhsdyJnL0j6/GppFIylFaJyduDJbLJvBHch
PtMAHLVV+yfyqZ2ojZzX/B4xtMN7gHdlQUCCJz+2+gAyiaMEhRpTxOvRM3S8
fefk4GDN9n4u25ipv30IkFBB6ou5sIEdmCDOdh64OnQbPNH1Bw4TIuFDkjvD
o4uZNxGWMqjjX/m12lofX7wYQ7+3uB9U8XfaI4/NOvROTH/Jxyh2VwyrFtCT
3D2kGh+nZkqmYgyuRWddw0GnPoaaPxbRwkqJA3J4Lk8jbcAEKsGLVNd+Z5on
YP3BVwM9HR70M+6e8iZYaLV2b7WvS9UF0PeMo0bEvlCModwHw+Fp9rRYusJ3
SdUQCQ2hhfhZexOcGFZbTZGjsAUrdurEhBkEA5aClxbU7xGF9iF2xeV7SbyC
pwGLhsJ7yTDczHJvG7U++Ftcu8p6qD1TyvS0r3aHnBXppGJCxYwJoS9xH/3T
Y1/W0Wq7VuU/JfaKvoyMhbuxEc+pu0V8qCobn8ZXWZnC9YXwm1Tm1e7p6sUD
0wnRfdUicNgtv813yPyxn+ryK0GrO3bZ906eMBJ+knXofrAKNxzNlsmv8AZ+
dMLkyUFw4R6n0KYShlT0w+4wOl6l7dSe/XfjRpKixrskeGMqL5HfHD6sL61n
D69E4MJQfIk1YFa5p0XtyM613o8W7XK7u1592X15m3YjKsTiH1Dk/7KnPvz6
B70QMvqxaDa7enQPs9KEac/WrEgw+JWawLAAbHE9EkVbtawv7ORcUKX9SVpu
7V6Vd6NGdR2REELyzu2aB3Lq4jdkR5GAWX73GvJCqb6gipmF7oF5cpsORoBo
KZxPmxjkUOk6w0z6SoONr/4O0v2XctG8amEr6FoNWdVqavNabAo3jEmVjK1X
f1Q/XJg4H1bwe9OdgprK5o/EdMnsCa1yqFPHXMY2bEGw76+ACBIWX4e8ffOs
tLgTK3JdvCGEgI8pvFlOs38uTkfmcGqupRKkUBiGQOGliQuBjqgfcai9YcjE
nEQ7PNDFCmzJql5b0xzyGC2jLc2krLjwqHjHuhiShDGWKMLG9709iWzHHSuq
Zd87G2WKHV0eUdasyZMIkT0kCeBLJiBxPFi1kYlMp7VMf7qeOAphMwbRI0vP
p4QcArhjJE8uGt1oEM3hHkmUjJG+4GWcnG7xZ4GdKocPBw7OHha8n/xqb2Eo
1BCe2mIXj9VVPtMQEoiAMS3Vcdh4SB6+VGAtijgNvO7vOkUpg4XHP/k0MCNG
X9oD1PgpZMLRStqCF89tTnsMZzHGMJOf9NuStgJ4tCSW7WFx/26X//QVtoa7
wVmRYFpxcpOY7CCmHvI5AkKLyz4AJtKQ1hD4MFwMSi7dra8tkhfPKFUugHe0
twKpooXWFWZ0hc7c23CyP84KTiW6hPsNTqvs5Pwtr8ORnrcoKo+YdtTbitF9
yJun/XWwg6d54sEIg/g/XR047qa37xOAC8yr/mnR3ml04dq21s+HTZXTYz94
p5Rk53+mHqukLD33E/Zi4arRCFcWS22RJm59/yTZHMEkLFZi/wg0/OlUFt8b
MelnxQ4zrpe+JneDs2QG3QtONheKoGhpJaiOPX9F5Qfmi4iPDF8AOp7j9nSh
7mZ35/qtloLrLqVynRRIg+ozqz3DK62GdkY7yWZ7Qx4BWStoMsjLymN2zfDb
Q8fO1y5CGCQFp9Ze0nhq3TDSKh3BeYPiIQqK0DiGFoQz9u3Kk6TTCUv4ez14
U2deddmqqLvWnGSdFEfhVzsxr0yPJvJt+VldjHzjZRI8ZrSCrsnKdzf260Lu
Keb1QiijquPWavIUP5tB4noXq81AXbFlDs30mPaiHdFJtNBTNEppcAJl5DKK
db5q3unzbEnoNwX79z8uFnWWe4yFDYjAfQcmTINWazrnkNlq9xlHN+NGm8Xj
Xxhw4TzDqr2QHDrHNDd58fz/4qT79d66QesYspIYMrN69ubJKq0RQE67erxG
Y4CeMRgqbifKowUssH8f5R08aiCWAIiifvPaincN3q0NZdnSJrqVRCTu/KPu
JHUdDQi9BHh+Tchvg4AEtsYbpaOyHygTPlDX6Emza0igwQmDLkc1DeLEvPFU
1VkHk/2kyR3m50yLVMzsBFo6RTxz5UC1YMcnJm4UZGEt1d+lZmsMMfrHKMFh
rbWSVw9jLDS3ivpFjhvEXln4qBsAVNC1CBqESwNdPyErxulFYx+yU/1sEBlt
QnUs88GcM9vNfzD8W5QgNj93eNo+dolRQ6aP16mBhKAmXVVT3vbhN8Ee0vvK
gQM2KuAEiy/Mfdwl5r1oabFjCOfyYYqhK1KgPMQY6dsO3pJHHi+xnzy55d8t
QxWa5ztrE9KehD9v18dQrhBIKDpgF22MbDi9vWQS3ukMnlf04g+ezMXQ5NNU
pbtLVAYpyb6x3562Hcf+lntXOS1kjIjRoc+DJ3CiQR5N7MJL97ThP3BaV69u
gJcz7LFo1qL1Pl/TbjbIB1mMmOGcR3qrX1elCwIKdlXPhfRtsF+Ev5y9LC9C
Jz8atQTA41NoOAlbK8Rr0YssiiW4LgmSLkEAflxTadkKqs5piTV3F+nAl7Iw
RbeMomwVes9Jns3VGPOdGZ1kFtIGXa9DGS9UjycYGVQlklYm1jqlYtY4ylpw
3aCLPOQe2ju5ezfvsdkbffQqF8n4nDnw3YTfKbU/LxMKf9QGheyy5lRjBkk4
q9ymg/R5h10XRJ/l4AIMZvBmkEnw81c3r3+V3eV/B8s+FIiiSr/Cpe8h/GVl
pnjRy+fm2opbq3IqlnbaxXLDvALeDJHIX8+11yaIAE7f7qDwrrcWbVoH1fiw
LNQvOv4cwr4NxcfZodpPHOvMjrmAWx6inAmmAUEojMOkWPtxWyL0Widr8bje
OfEOhBg+jXChgMUnbnsO1CdlgsxmCsd5HfZI91XYjaV/sRFjuW/91vzCp7YH
CFaR6jzZLi6UBrNaRJgVcvQaYqr27O/RbZKc0EEouP3mtuD+pAkZIbjofd9m
AsjkslogRBDsfeNbojovrye6arAZTqBlGxcXUX1xjA2umRwLHTiyzo/J/2vo
rmqU/d675VqImjZzbPSNTGQK/Xc0B6V2NaTm96UHSMGRSUmNV+OJVaX2TVj6
qrlMg1+UuzQ1v2rRGs40kEpf8D9RCEm0gyYV7PnXlZLdSHojuNDT0cl2dHik
htnpixd9tx15Gls0iTj2mAqQ2ND2+g1lzPbVPKWueQBiMdezNwffCpmE3/oa
I8wKCTsFcwKAsRNO8aM/O8lyjKI6/MSBXPB5H3/+9inRdKpemuWDHNnu49gp
5fPwA0m9l1IS67rytQkXT4V/FqjriifCb2iMdPuZwxL1QdAJ0eOK9oadToJI
/CbnUDnWQ7Uh9mf3ua4MT2zW/HdnsDJUWMA+I43m0owV3M6mWcmDvLSzYonD
UwgqZYMTvAsMj6EankK487QQh0uoUsvey+VmRPIKjADnOIp0Oi1mNoR6EM3T
StHdSDYmrjDIy6+Ik8aTxvqbDVzfXqFQMaxYgc4vT0Yfq+0eNOVHjkOAMmXn
EiD71TfiVIPQ9dHM6QYjOjf7nQ6lZjztpfu/IWFhDpb6a7u6mdMhZ6Sw6Kku
pPN9azh65Ww3jA1CquwtYOoT+prnKMhPxAT//3KxfzI/6BI+aMaVt1zU4uFu
werFeESck6Kp//Ailu90GKMPTkqM5XueBHplgISRuX5bdKK5FSRg+TSyRMXT
mjWLG1VAdaZfyL2oHGKh8uL59mn4xx9DPda9zWKE1FzMU+tDE0ORcoZ5RWXV
nMYjO/2fPVbv9PCimLoyJc1JzstoTCNvFS2UqqwW5kCA9+XeynOWqMlX8s8a
x1+psAEDDSImnEIAoHCuhmOPIPPEuJ1xlvSFclfYwxa0kSJsltWDmiAqPAQJ
5j5hb1VVUDJ+dxQ4RkA7GgDEui9duLx1GPbqtzX6ryZwHob25HzwAmasK6/y
yU5+canGH0pMn+d036/ryd+TXuwHw23C9uQyxqSgxPN5Xdav3axrvVC+I/t4
2na6OMbXRp7hVM9GcFBzuw15RHIxrHX9L52RuTGDtAOhjt4edHytCydS+MoX
bNP0N3kLjYosUAy75ersWWALkM8gV/tNuwZTJ2q0rZHx/B6E9Qu+28/gIuHz
Oh7BKONzclOahj6PVKaaYSAeYNCabobNU/BQJUNRxdJnj10ibqYd4HefYu4/
3E9I9t+NcOiWcvHJa0KQsFUVw104DBuzmuuufBsXTHHkyM1XUqDtYI3uyRWc
3Ca+21Av9ETuu9u6jnk7YL+SfyFPZbgZ3Wg6Xup3QpB1JrDy2n2nwZpGKbnf
VlP+8cFEhGHJb3VpgPeY87BpO0KYDE9Esdz+wyWB0ntrLX3xaGHDBKaxpXsz
zQUkegUNu/S/R66ydtPxHs7qJpe8DP4d3AmjPNJfgowhgOd68ivAF0emWtRb
P2v4Ie20DwJ0TbOiQdebJhUeyjqlJEAsY0gnsGYorvUcJJexwxxancmHpqPl
qrHjiu9HsXHqOiWd4aSNAuDoMmEEEvJTqGsnlK+lMGmsK35Xgdt1+egkHdA9
96VHOCoQHxdVVngm7AokDEsYrLfn1aMPuA25cItxu1NL9z/Alt076zhV3fvl
mvWP89lwbQ/0THIvOYTAqfbUvl7zeMyIf67IIgihJEEiu/FjAk7WSBRKiYpd
GWaPBVWstyAuc9HfQeyvqNF7G9MEli85TRq00CyeOggo76aoRaiVameDw3aL
pPPjiU/RQeZkz4fSgWFy6hm06+mvKPa2QoVqhuz8tkqdRSLIEZt6ZZA18jWW
ZFSlzzT7WUdkZhGYIrqGQzhKfDRbhpncjla043ultvRgRrDxmWFsQMcnK2Zj
vkuweUE61Lytg0ArzVoe9x+S0eXI6pyltVFH8Ly8MqWdc58dscd83NOR+HJb
UwG594HcEsMQIbfndEQtjaAiOUwDjPNqO8hCaQ4ryUcyK893fq9jRIvd42iK
5vxb/18HhA2bZK3h2h1qwPFsIY/CNxOXgfDqpeHXdUPKVc5Wow5i5iis4pmJ
NcoG0dRVu/Ma8lSU+gSzsYrsUxJhFNCR0Vx+/iwo4TPSUheqFJ1s6J7esguy
A48+wxx+0UXhMQk5uOfQuhX4zGiAJEXuKh7noNdON0mo2jMuAtUdzp/6EP1y
JEpe4wh9V2u9CfWHDKcDkkQePyt4cu+iuFGwWqwuXy8iTPLoGRL4cLCmcrRj
m493AaRh0jEufbfpY44WhMsS0q6ZUHrc7U5MklMJQJf0rq/jwn+Ft2k5cZ+0
X5Ogymiw+khYegjDIRUGHPLUG0n+GSa6Pw0705hPtq9evzzFYL3MD3WloQHl
PtNZHhF3yk7rbc3505NYV1dHANlEAtV7PVfpybjbZcZ2E6dhE8QQ7VeZiCFK
SeY8cZHzYar4nMYeZSTi/0De68HMXs1J8OsiiP0fC+HmHluZbC/pu/7YGAKH
nz8J+N/IPWxpuyPBgK3Pi48w4TpRcuwCT3A8LUcwov6PqaIf7iPsd8tW2tVx
vVP6Jhb3UyJohlss07k4CufnX39pLOCQ7PMcbmgMG2vmyKEZeC4WYk8YXId+
a0iACRfFo4VlWj3+YAep3Vy9iTW45oq73vN25nWQhIwVBs24yvhod34/QdQq
do8IqzkI6XCOkbGhg/5cz1/lWU6hr99aWbXsvtOPNqZpSqov09+GzG77gvq8
jPoVQFmMsDkIPJcsp89W6gS3bTMYrHQ1NCgy2LuRw5KdacV7CMZcgOVUt/9u
dT7MvF7ogBArVE9xCCFmFKCmjzK4BiC3IvPEsi2YEC3TTJ2Y9GGeLcV36Vb2
09wyRu1WbiTDalri28NvJTglToKTW9YWVEhXkOOSL6wOwMSp5D24BTm5SI0J
/MjGU/2Ce5lJXIXnsI6fllU2ql7IcVn+0qfcUpvj/Re0Jb8Pv6GOIWLVLVx2
qetFS33TZq+Ob0ucbVnUVz+hEUTO6rhuEnEWt+h6PElB6l+Psz//D4wJJBkX
8j/7eN4TJ/g/REeKVAGYmX7Fxt1PAaIPc1Z+xWD5crybmPzQwZ4iDaDGUXcX
/gJb6KHGq+ITTDrA/vTWem59veeSmbLgpLAdkZIf6j7PZEdSk1mB+1q/iUJW
5e/Cr1zdRONXDqeWwTXG/7bUFJR76kYD5vG0jBAZ7l7ZaNp8HCNkxwG0AAg8
sD7u2TaVwHZ4Mvxqzm0pbZCjQX3SHyTKO3Of3zK2wO01aUoCFEATku1i5GA1
Lp/zmxqr4vqxhNjN1R4ln7FYn1RVWKRwFZiGMHaQjQ3558mauw9jPihRr5ey
OVRjzQo3NZ77LwSDFqA7C2dWaUjIPWHGcWY/CW0MPLaSq7D0KjwOdpOs8HuJ
79pQXjVZABRmSrePU0tKTz8vX0TyNHGnzjFbXm2sz69URCrhdqjLSCbH6W8w
UWLy2I94vB460rV51Pfvkvi1U2GFIkq9ittk4IOyr4NwLO+x2N2UM1PxIVYw
usYVL/3hiuic1/u8HI0Dy4fHTimxQdfc0Qkf0AbDIL4QtItZeCXLX5SLyoAZ
ht+mOcFLhgxmk2hBOsjvKQbmzY2n7C/NVRWb9OUK8nUAx0cV9gJcD01YSjWS
AkBhPdxj4HMfP6gRAKVxG4GvAzjqzizW7OVApvOodnHJNm1cBBronqSBZojT
r6vsI3EKTkLTtEl+kTZ1J73YhKEg0+Em+xpwJAFsvUH4wqyJ0DQMeJxkyVAH
icE9Sfb3maDKpusf+hQofnntvN2Cz95HLn0KI4sM50aRG2EEIaqiRwUD0yco
BKkwKtHPsMVbKDfm05AojhQwfEVjtbbUKqM5FYm9+3PvVcH3qFyuKtm3opMd
iAyq5jmcngmn++hWN+4F3slzZnXI4rS/0R7KdnPHTO4FzQeNW/GdhiI8+2U/
YiZmc1NIF9bAYVvtpzpFKZ9ciC0w4XJxi6KuD+OEA1ZOQ5NgQntkc0EQeZxN
a+iofLKN+w8WQUdnj0SKGgkaB2YZg+DANYpeFWsH+Qh7RAUD6Z95hLS3S0V6
QCatYvZ0gq+oAklpYMK44gjTbERd3l3VijbIp2qu4QHhbzqaxyZs/tGu9N7W
O4fnwRgjB7ri2cau3ooUTbRSMkIB3GiegHBhOtAzrBdUEE4lwhoggE7wfMkg
bRzH/Bo3SPHAK9UOEyKW9HrdGmVSITeIgWc/YE2Zra6mJootJrXuM2qU3ydf
+BO54XEsXzXNcRYAoy4ZHso1+td5XPU+X6fJawtXw/LC8pmSszgeIgfyU7cY
PgzVdmzClp//XGYE+DyeFABSNfhGY1F018tHSRZv2MpWgH5ngJ6X+LUqGrqO
zvpLZM8NG+BUaDWS86QG0J6r4ZVMbyqLobHzER0j2/aeWIR/PaOXNLXKw8er
5glumXSZZnqTk1h+I3ik9udorvSaBe8kTjxynWm/ISlK3aG66UBgOahCu5pH
l+dYNvdyaTNzK8ZsU3/EZweRLE2dwSuJQAlxVSPJIUrnfkjhEj/ZKbiKldFb
sWpL+/AR9yhFICexrd0I/y91iQGGIhTULKuGPZF5/V7VLarVhWAaxCZF68TB
8/mvtxnxq3V0yw/G6OsjSSLKsSRsmVzbUrdMT1JohNdID4ViB65HcKY8PnYb
+dtBJXhBELt4UaRDRr5MRgFHIF9SAA6HUsp9tCTMhFACPPMB2NYIB6DDIONd
yjo7Ivi8EesWfDxLxL1HLU9QUaDGhTkgx0FJdo+HYXIirmrBauCkQpBu7agR
0RjGeAjtSXriv03AW8uUajOvJsuDFnxD0HlBjvF99s0/+n5Rb3NeuZ3F/pa6
3GPDtFWDI1B0rYRj8JyPfgXbz4uj2wzwZasxoJmB2AfCEWLDjGtF0J/JU5If
vTQWCfPMEuUEL3y9OvwWj02lwFk2qF/2zSNCquwMReDSc/OaOaxLKP7KankY
/LpKYrizXughcnXUbROrpvEuUdfinGiGHtriwXOtJiqEqJQkE2WY7/y24Ks0
nn5dEQ+j9S1rhFWaRblLbLivFQ2O9F6RxgbXUN0oRRwLqTBf4R+B9EN0LkE/
TvzKontGzeS58Dqs21eG7NbIaXPbtLiTIZLea7dOQN7jKHmogKVbXSsBf0nW
Z6VqS/JFvMip4+BHKf+VLVp5SHG4K9TGJa+zE4WQ7h0dPjokrtdmLgZ6PTsc
EZq9KJWpYiBlZ5cmC5ZdBYG9q79xd9W6qYQIPiJSMISvQlI3DBsft5L6jo6k
h2d0dwd4v7Lg45eL2fdgB1NJRsupx60L9MVPEepbr8a8fyDRdj4RdnTO5Qc+
/II/1m6RiV9eGHWsPp+qotPRjeSGkyXgRVcS1A/r+lZ8d9hgtfsKK96xutpu
LGrp/WeqeQ3f0QqqJvOuEiG9qdBotn1Cv2suNqBgq35pdXT92sZZSP1CsH4I
9ixHq45+uNN8orGyH1vtY3mLzU8Ziq2ajy+rTpj9Vah2kC1JDxfvaKlocX9E
ukhm5V6dV1xzXHWazk3VepR+uh5iAuBK/HFjxURYrT3UfCM3f3qZ4KnkvaDU
K0g+6++u1Lyuz23WDjyn6OLKtmM3z8C3Or1q4PCjnek4NPwZk1NN9SHttnrU
/FoPXqZse7wFR3JTbKQUSC8GM5jjeDlWvTDkfoQzeu050f6QE6c4gbP0+zAO
SdMNGse0i9evZTf8n80bbYKbxDbXf2LVLnQW8wG6n2wyKbgwGA1Tl29mzUem
JN22eTIlldePmhBwoiTjw+pVURxjq3mqFkzcCH22WL/Zy14p/hdg3OUCZ1Gy
PwTmdJfSr2/rM674A2q5jLjH49R+mDXyX/JUm9jARumI28F0pwgkJgUg4qLR
E+3aQ8p1/ZprMGt9NwiUY/ZW/zJuZ22ZrS3UYClbfYLRgsOS+IHBkHftrqgv
kuC0OfRH3THDKJw4VewNYleHXRJE6dTmwVIHz5TRud7AmeKRwGVczf18ZRXz
4XDmJJnOeerCKJEKk3M9gWg57dhmznu64rke+668pAUXTudMHiteZ4cjYH86
I1aao6agzN+Ft7sbzV8D4Rkq/ZnHnJe/OAtv9/yT4vq3QgP2/mICnaVObLhN
tw7W2jlo367P1Nn+zrL1WhriYHffHL1ZZO0kXhkNHKhDpyMlrO0a3yeK9QaK
/7o/fEtz1KxE2kWbxkxfhg++zJdVxaik1FU/JGLnjx5NliXksSNsrs5Hkbhg
zMRsOwG3y33bkhvClHBND3DTq9QTFpPFt+fdOkP/FhVpr21rlrrt40jIROrc
z4g6HOtkrybJp0KwhXhhsmkjyWC3BpElQNzDaiIGYEa84VuPGsgWfwgqsSUh
i1tzpCIsJGDhBIAM9aDV9fBBShTG/Y/Fn/U7oLhzlKicsi2Or6Sclx2zCo9u
Lw9LEm3hx6eDddXCh6Gv7Ia39lWViZl2NLRy6odYnO1f8p3+haLiqbnJJ/P0
tUP0hvwTmrY597GXCI1YkPfgr6Qvv4kMLg8j172fL8eROHGGI+jG2uvaKydL
LMLlytEuChM4UEY2LJT9WRrgdMGESxmChEdYXviuS/9yLRwwKBD++5XM+DD6
/bqGJsfge9QHXiwB2T7jm3zm12b5BK1qHtLqlrGerZOmcYoRH62QkmhMuUV6
Yfjd2Af1Ktpu05fUPgSrYfvyvSPXjCSvIzHmS6Nr3vYfoVXdDdfR+LqUDNOW
6oWnTHhJG8IpA0qkmX8AR5PgZ9aHVn0ghEf1uFuAaWtxmLYzDGKDSWKrX8Kk
zS6SyS+yWvcabUhs8ffclMB9hAfTDxrfIrhQTKFJqCdaHlQx8N2eYIwFN3I6
O4QnTj/JY1mMqMCAwX88ZeautUpBAhhyTd/+AqmtLz3nyEh7qMGnyCXc3Dbm
a6EkzC16wYfpq9oHUwkGIjjmqNkfJzOQDkOC/JU7lTnAS4hbH1MJ6wEi+zhX
3e8aTJ4G7qmZYD4Nm3kSAqyIhxk3QKEqyq0yS4Bj17d2Avi2utnW6IWPPYlx
ai0MGBSOBkF+4NsiAxjyhKvFy/03l9IgzbqGno5HCq5nyJlsJrLXRmy2IH4s
UWHvJ78cyUaEXRJA1E1pzzI/NKgxUutAVHGqjf+WixYAHM5XYKEpiSSJIOL1
YdEUQB/vu6oVw/f6Vz2zhIbuRmydUNBkQs+QvjiHXJd/PFq/s4yzqYCd7che
n1bNcQLsVy6BnSyeEGrSU+DKpY9cerQ/6K29E0zl0inVhzaW2Z5EwoRUavjO
bEUWhux9O9EllnjyElinOE9b0QNKTueaNYACNjkHoDY27ib9dJn6IE+HBJXl
DZW5nqHiNvEjqSRw8bVp16vUEXNhZqmP6vNfiWF7c8TlR/nepxkMPZ+HXGbb
EFbK/C+b23q6Q3wMCuJfBe4jauwti1gPeyEqPUvkdPM+0geJaLwFcnuygIao
LjuNzizdzntmr4e4LswMiDnU3Jms8T0F8s+MpgbbabYr8c7pBZ4yNHR2jSsk
wrboPSEewBL3suCtzVARNiBDBOMXK/acOEG/sWQUBWUqgf0oNws84ideEnlI
l1X1TBl/gAnwnbRTThG5506kqk0KR3TtbT1uomC2OdIP1Ui0Xy8i4iX8p98H
iVKffgwo+EU49FQMpcTc9s2yMe+j4VgSwpFNxt0ItGjIcnL1VgpsZcTanqqz
CS8HJ+fM7cuO0vt0TvBqHQLOSCZ4RoZ9zEFtWVLXO2WuA7QZsZTgJOuvbl62
FqMQm81e9R5zyqZJYa0slvDMCHiTnAxHAT1qsK1zaGAkyyAIGlbd/PSQD5Re
gU8kxG8AZYU8bMcmB8NlXNOG8SAZ59R/bsT9pyn5q25Ai3XAUfueBbLT2hTt
YikXqNODq/A+ze6xbY+z+DzAl6cOTDs7PzNY+l6NjZe7N4aicBIk8mRuNfvv
sGvOwl0x/C5YCJ2MXhznypNSZ2BEJso1H9zkXCRSEtpYtPHNyCbq0Mvfrks0
efjypHUtCz/eILRyC5mjPvIchPnlJBJB7ybWM2DaOG0MnC1Vta9z1pcYpqLa
bXrbbGscdw0JBmuqvLOQcikov7Xz7oEIbtdsrCuR0nO+ezg1fToakfD3RHhq
xXTqoKjxEEER5GkamgBXNao96X0K8gVAkXgXvWsg2BeeCiyF37NxKQ5NrAH3
CvEvFlOxwsBrDYDbzwwfiowpVj04S5LkyJH5Wx8FqTf8KOAjVfULWUkoFbKS
AdpXNYEIJeDq5UDo1NturPkhlK72RnjA8IvD6N4fRxz81bw1+16V0iW77YUh
nwNzoBQ+M4jUCehI83/Tawojf1goeXrfuTLWYaKiguiHLuvNWPRv3WuaXCTM
mVBeQKDe7Xhv4yuDqA7GUph68sHPRnKzJHqZhCbyLYIdNGgIPssW9WVYx3MO
XWtrdPEJotvRBDqxIlHOeNJQGXh82XmN0dgaB90UQZwdD4ldv5OM+Em8MdUX
6NCgE8NKa/SSLwyJpuBPtG59F55St7yUQNrqzW2/KCHmKaVqnn1muw7zH4WZ
9UeFXllXdNL2nHBKKfp51RMJhkPmGy7MuOXJp+PQa3M1QYOVEIhLgomk9SHK
euHwaqWmgCDmQ5CxCPB4DQvXYBs3OsmJZMAhqzKra53T7yqRwM3EXzHJBBmk
x7COduXcmyL02ssgFjLaVeiIY4C3THgmiM0CcG2UW++bz7bhqYx5BQtJEj3a
O/Y+P8Anakh/ALDt4o3MF32FqamcsaCLAryt2EFCD2TZ0OrYF6nSCzT2ThI7
c3H4TNK1Rekrd5freaxEOAy4RDc87Fg+qpsD4bwkAeXSB51+2+zf7VZyT2+u
H2g+L9P5oCXLZhURzTDLYhH7epx/aeqpONzD8XoXzvRgDh7wbqJfKqjrB0wd
DV+zZFIFUk2gdEpC9e0KT1IUvF4NtZR0JQ+wOWKZ2ewBuR70eda5oDPjZS8X
+J7SKIJRxW+gCWM+bnUdcgLSq+QU09JyFI9BQMi1XO12B+IZxtbw8n8WEKzp
D5nf0P7tgQvtadX+yCEGV4GMzT3UJbgs+FMuHYEzwcTzzm9rr+VpVUl7mLgB
8SAGnkzCqqpv2n/u+l4ZRjuheSsJxSD2NZAZUcieXr6xnEGwNhbxw/v8lWQi
AWqPPCKp1tnOZ5VbMf0trV3NUdVMRcYcDNTZjd2j343jahvKDxNOuaMcUiP6
pKoot8LMCBYMBsNPevb9CFsPQiY18WgjNjd9SHnzAX6Grqa8eJU+jj7fpDmi
nGSzQ+HHONoo5ExYLPnioQHU8mBGSoEydjFqU0MHNQ0hdSK0JaFp/mlWuLi3
UDTK5Wn+D9DXk0ZBoEtA7CLv1OdwLU9JYnIaa37kx9+KCZUvowQmWotXmSp9
ylHBiQ+VlIFEvEHUoMMp0pwh3e6Lzl7n9BBlfuJqNie8i1zxD6VHV/JvJZXs
Qn+etkLxK/mec/kpNCRLK3Xgqvq+pf6JVGobNCZuQ+U+vkI/olGpHYeBNsHi
mvuR96VaX2/0kH107aKBgTXJqD/STzMDZH7HO18zsqrtcK/30pVM1Vg35t3U
kDQDr9ZYOGZR1sSFmDI7QXz8OlmYIFFsMaV2YVOCLF8nbDwnbL/iCKcqoDIu
mSu5onNHg4w7YWW47yQJgVhmTDsiytgjTWlHQ74O74/nVkacUK0/1GNRHW10
FjLW6BLHH/97unxBTmYCHz806cjJ7nQ/TKYT2IFMmnyNfkebtk9z8uo2vKJa
culo7MzzyP7irbxxT3DYe8VAsoNXj3tW3aUL/CzXxdXcLAiquIRM8asBrem4
uU1jjPQFDlfVttmE3jWlZdAky8v4OaNqyqcVTVLyDj17mM98v5etk50WOawg
SiVRZH6oZdo3SYoj6/52oNc8Klhee7X7byGVfnJOR4I4BM5oO1US4PoZKUbX
z7e+nSU6H66wY340jr1BGInkYOAzDvpUrv3UTHskb4kKhpVkQOOiP8M4cpyH
2XTzlQgsrBeh/E8GBhxAQF9aL4vJh0Jf1D/9xGwVX8GRj87qV3yLWVEIrW3G
UgPMAqdk7JEMc8Jh3GzL3op0EJCw4GWLUWEQQsXwvZdmO9aIMBADr43szypc
p7facXUAhEvPw5PNhBDcXyu3vayb5l62OlPxJlZ5woq6r+f6ByCvd6isEYZ3
giJ3zo+e5qtnnhxVXT9zlzxMtk4oT6P3MoKC4AeaaJBoK/MvudAgSYV7gZHz
2GAcmakjhTQbycHYsxETpCAiBiq8XWTC4vnDX1uWvLU0idGGPToD3qLKDRR0
ZhrLGLG2MSfy3cHMTtI4LAygsWoaLdXu7gP2R7mS/t7uKVWFgq8bM4Xjof8J
JSxR6HpjMp2i96JOuJRIRvJmihSrnWeDfe8hk4IlSMBX1pwjDMJC40woCbxp
Nps50IdiHM2enDG4UEmwQL2s2CgtzNoUANP7ffBi5uAeg5v3hYcdxRrCmret
9YA88COZWc8oA76HKLvw7OV+tVjy0MyeTYZQAD+ylYpWDx2HVAXOACCs0P3z
YciVPACQHi/RJxnJT8lHioJUeHcQDuACrBdICFCTFk+6KBexIz14eeZOJBtL
TunSxQbQs/WYqS3et8MACiIVolwnLy1sTv0MvVyhbAu/PBQuUwpngVgPmzKf
txPvgCD5ZHkmfMLA8Shlvl1aRouQxRAjVyLFSB74IkPG23jJjnQ1+xS19Ylv
ikzY1MtmdglrvNLMUteZAl36MwSMsVWvDd8DP5uI0UE0sfHEg8ykAobBe4zw
v7+GDplUOPm3HO8vuSqsGfToeMra75DsP5fVb9iebqeHXpya4+9pz6Hdy9Cj
J0MsbR7OPSjDuQl2XXTGble6AFTP6NckMNOo1EDRwt27yhRGGp7EzXmNFPGo
Rs6MmimhDuzGiUwQcmNCJ15X9csamp47m3RfBNaqNCPnK92AHYwX6rrEj0Pj
8a6BBSXQ8cYn2sHeMr4BXIa4jPbB56PkLOlONHu+m9p63jOdvVDD7eCPs7lF
ZsUN6n8zO4oag9jX0QkEQSJBF6Q51MYVX73C979O9kX+vw7GbgaH9yU7szbL
sqUEftDL9V8JMaGsiUgIamnKxLJWBmhUBI50E64bwOEMCg5yqt8mU5DcFm/O
O8sByvGetanqyiRtJt6+/dfQHah9+7y0TzB55yeihLnvuKROG++Xhm7GOh2Y
U1vG5TA09MeDR6ckrMh9gBm6fwBJe4z6FI3lovy0yjZ5FcEf1x9v/tHxzB1t
9ymf62vhUdEVagGFmHOqiOl/W4lP4BSvS2tyA87L4+SDxfH2bNQT52XkpVe9
DlNqVEYMsAoHUCHv/7sNLmVZs4FoKMfsKk+r/JYPkdOPZ5y/Uz5G3rBAzS7H
WHsX/aEjDvSbAl2qHBIE8+NiafUda/PdRY+dSdxV32rs+ldqdhUWI2G4j1ph
Yen2hgaXQBn54EFXsL0KuV8GnCnJQ73/CQ5pBGmdmoiRkWwoBcDnSZ0z1A3M
CbHHNYWdkIqSNXHi40y3MGT2u0NHsBYCKJqWeFOnB/mxla3IizSo3i0waaFu
D9iZaoWralcdl1aRAM+M7vD4bQFdxzPyXzqlqdSCK2ONsj9qJjLHYCwWP+Qj
Ji0o/ToopthekcqA6JFRKeLj7BM9QNLPcusK4l+6updVRJYXEKQajlXSjh4U
WiS04m+uTNGki+Fu4wq7gM0v1ipuESTX9uaTYN5LWISBSCtJXxWhY+xx776+
Po08o1eJnpSrX79ylGKhjEXTzZF5NCXpafHpVAIvVSLPpaYvJLQy3ZAjT+id
OfVCWdLsHJKiHF7jv0aCx/LIh7fZfp1hSXOlEoCsiXy5oLOkAZ8WcmK9SMDx
yhUsIWS4rloLTQ8ac6wqd2Y6L3S5ZsL0w1+5ecaOHpg8d+kU4vpw0jSUSrjv
z/2BMG6ksLML/DC8cgOZyfTWRytrL4FR5iagxJ1NdQHp1Lhs9SY7vdhtZHyi
XVcQecwszTraiMZQtppSIEbGMTfxas00lIENqCpNPkcw4ia6VePZ9mI0sCor
XPMoa8m0sp7kCobpZRHQqKpmaBb6dm7Ur2cLmedzu60na8Dfpng9Fv1LwVtd
C9EYiPp/hHLARnEUa6g1qyqpcv+ONPRDUlIdJ/MdN5en+ZsGtU6The0ZFAkq
LMObZrGKtiRrp65M6Bbv6DH7gFIsRD6VHJxLZEdIVz29YIrhBkJX7UI3AMi7
Y8ftU9OD6MmyrZ0+hgWRD0jD2MVDGHzJw1rKjyHdLWrlX70G5HIRwsWzKxwX
Q79e45z5URG0qqO/lRUyCUzr3OApYH5MKbF9JVlOVuTqAfwvSoXPJ6du0Ia+
bP5xh+zWBCM4lBI6GtJ5z8NzF4e9zpUjOV4as22dhTnSClMAcGJHucq2zCp/
kCGdDZCXW/7SmdABTUwxQ8BxkEB1wvXDqAVMUj76DMSfefffA66HJC2fW5fQ
MLVRID6Y43bsm2/qJD80xrSqiXR0BR04N9KuDbJnaOfo/wGuBjDwtqHw1Qq3
tZBGJDTgMoye1XYDy9L2AbaL21q5A0W9qrk/++plkSlgF6yQLnQ/eZ8Vgaej
vpsDkirkZFCQXynTKA8+IBRDnItnVCeaiDr17yLPqTnKGvBJl9qaBrv4LoR6
2ZGJPIYlbCn5CT57KlmRvsu+8pxsJlVrsUf6A4SJjPelRVGa8Stroax2ifsN
s86DKIoMh8cJFY7qYS/Om3aEgh0gtsgsqsLaEkwdEjJ/OZX/OKbGwqFq28UC
dxL3+FUfna6x2C5Xq1YMElr6NIGBb3e56y305SXNo1BW9tCRYQplr1uvwr/A
MWnKqG7G9+k1ZyGuK05hEyjO/tUaGZ2w6SB2cLCdgvFsceI9fOiid8gcouAi
77i1p5FR4M/z3sG04REWQTJNHU3I0/CPPNRufWCltFJZaSEJy94DU0FJPgV7
XkykhP5btdt4aX3eCBuZJbpMDg7gz3toJiGidgKa3aIlea2YR6+E3ejSv7WP
rDiErXwP0VAs5Oah/NnzZUK3N0OV5ZMJkNq4j25BXj/vwJ/vZVMzbYLYCTDA
CY8yJeAPsMVMcOr8KLf1xrpV8D4C2q0asj7cQeFk6P/7tX8j4UePSPOArbY2
cS67nyCpp/+yHRgI/DUtkXJjNY66SY81TkeMwpyRPJP25vxSh94JtT/RgQ33
CmThTjj2IlrtEOUD9cFPAHGDthnWch9BjbzO1hhz4n/ttYyLMnS/d7qt34H+
cwDyDsAbtOoePcG6VhVcwWc53KqVB9aimQRZUIBzUd0jA7rTJtUYu49po7K8
DKiwTvPgCeNWVaLFpL0cUQVNjZEN+kAcAw33nv9auzNze0C4aNvPdHUB7dxM
uJq6EIWZudyRxI2fj6OsV4eJqKRQvdB44mfs5LgKK8KlKwJUAAMgc/Tq/Gbt
MD4PjjqjZpRUJG/CH2hof68Wc9Ay0EDyWcsaLVBGq8O4JFwyGRu1cCtttrdC
e6behxdpshjDozK5GvM2FcCDtJNesbYvi2BBTNmo/Vjq7YnFvtXlI6SXMug3
23Pc+lpr1q7/N3p571Oj/mEOEMA0+GUd8k111jf4a+hU0mseT5d45uB6LotI
MVTsWmQusV2Bsa6kyUyCMLlWiij0d/jPc0prfw5pou839IimyLTX5dVoYUlP
Ydhnaix33YEueappKFlzK7FLF0IfJmIYB/KflT/2WIk7kQRh6nHuZ9Bik3TV
FBNVP51G8DuF19VBUMkN6rz9ct+UsNx7YAVnEqroGLwmlWG9Yfj8rql93/Yl
85B2M54ysFiKDFTaD/uuR15RQVxci154LFaFzliB0y2D8txJN86wRpW7uNIO
Sfw/9GU2HyLnkKjZVGkVjhRfT2izR++SxPK2rUjn2eYHRFERGRUtXSxnXU/E
siiMPndtab0gHRogVFlpCrYQmE4A2l52Ms6O9n60hhSFiHM7Ka6LrFV2pwoT
IDuv42ITNog5y5nZMJUHWkppHuBzchizltzZITzMnUHRCw10sSwqwEaFtrmY
n2TTA2sJJm64rs2CeJWTmK+q5PLwmVNLgaA/hG/s6zEp9cm0/8KN4k9JpGFX
NXBbndIF+kjTUf0tyUmKs4Fr+zLir3sS4MZ8Gz6HbNqqomiblzPi8jP6Vpib
SFo93vfk1CdcljIEQp0Us/hYcSqjzT5VsneIU25aVYXkTcZp2qinrLsfgCyS
GFX3D7AVbtRaLAb0/0PB5V8uJ6/sj11Y/Ao7onkf8UkOMWJjebY9CRl+BgnH
xx7FjapgUDJJcz9MpTy+GlbT3pk8MKgtGixx7aSR/pMmAj13b7XV6kEiwmwi
zxSSq6urV003bLBpq7sV1sCNeUq3o6Z31Rk2RK9CgaE6YmMQgaKJ7RgClSym
IW+NxZq5DrHJ4quMQMCEUZITp4Dz1M3J6XexMzLA1c/0kXoM2vX8B3AyY8aS
n8iRtYO3Po+pLi9OGYRrN0X+nZj0ml94/iW8NMjJfi7ISyCnSnXNHGGPOsRD
ofRCl+pJEs3EVrgYkq3e7ckA/6QQLTRRDqyNvx720U5+pjyoPfZfdwES5rZk
t+z/dHB4M78nPtEgX3i6zJ5hIGd8p9/HD69edIj8oKapR3ODGe1/QP8byW2M
I41D0youkVPSot4RRzpzT0Etvy9MCnCRpGA11g4Tp85L4Fh8/UQ9sgWxTEZ4
O/lC6SYDV3dfpNDZ1Mv8Ge9uSVXQGlzXj3ZdUibrNT1HyFSTKVPXfNc6VeHt
PJ0ylBUs2vU4FDWQO1QjmNdvO7G8MBYPdhUjc31LbTgOGoIXcyZO2lNDYgho
56enuK88T+MdxVtYoBsHW6kCUqFCNY//mTuXdopLuLPIZx0nb0g2uBtVjCEE
gB00ZrDZ5gc4AWMX1NgummIPRkhQj/uFEy5UBpFmgleb1zV9aK64Y7hG2yZz
G/PpiUJZmrW9Ygvp/DTEnwBI26Mh+5lah+gXvyWi2ffZeIRq0D4TPaf4aFOm
xouSsFdzp0gOWNKU9tX+Bglp5YKkhD6PXTHCOiQrGabmW2mEdH4W7EpiTkKi
pimR/oIQUnWPU/CXcf6klP0c4ibVtxDDnqj7pd8ZoIDo6nyRKTykaZHXGWiV
AumGynOiLwaqHYJjDjafSdDjfL4owVA7egcOxB4vy/GK3rQcuZi3o4WkuzmJ
r5B1apIcD2GVmTpFRqb0JbpFMDweFwSV90ChClSLk2etaUUCB23ZZ8mMbDZq
MHuGxPstQu+007xFhL5u1fCaE1GHmlPEPpRJTygJSYldXrQkIIdS7A4fcEzr
cefiupf7ALDHbMtjiA2jjUoY8JAv82RT39t6N7wssNO1VrxVdjI52o0Yy3OF
H+/u9x7MtoRu09/P/1qruslVGvhuEyZc7UE0UATB0l/5ttge/8ezzl2e+9BX
RcwunyYlOintXC3qz6++ubxaZoGV+xC1A0bWKvgiNJI8J02jK0rrAq/6kg+W
l0n0YAUi22gufwfnPFfmjzIGa5jIB0hzCLxkjnXbSuPlXeVVC7j8oYI/ez6U
BNcjQHKXPE4a3qp2icb5FNe+npIFLnOPu8JAL8cT30tQT/MzsxdUGITVhucB
90CFSh6JZnXbelhoxHRcLH51x/Ah7k1qDDompNHaxwtyxv2XeW8vbnLOUvx+
Fll8A2MoK+i5vhFsw5WlWN5vp52qqObkncwGAK/1no2nR06VSshC+Is6IdZO
v7MW61o3ZEIdKXJqNC3A674X9b8qOklvbBs18k5W5/wI8ZAq9qmcZkWaioPr
9NRxVaaoofg/YRmRcU4rIer1+Mgd5f6+e6R3rmDMHXjHPeripoPwKZTIuJjf
5jctMgHBFaVIqtBptsuS5d3d3xj3P4FkMEKy/VhAs4JfdMwpT8xuPR3HLZPE
9jpRYck32V1dbkY3zFOqo5pb2FO2OgzhnJTJz21tL4GP75dADtpo+GGQAHUQ
PYg0tj63yQX2zP8d4CV6a2m4z1VQ96jghOh3w9s28MWc+u3US3MAgT3JHado
VBIma3ig77SdjqzW1pH69Y1qrtYPfw4uj+V7YOAKDvKdB6o2X9oMmJMQw7U/
/G6wP2fbhQeI9/Ts5MgB1X1iL9BsGRCn9hEcz72ZdiAV/g/EOvIFCyWlDZCh
hsuKQwKlYmTc/8KXLx5F0OUt8xE+Ciq3MlkgxBPl5s41IPaTjd1lArMfL6/o
j8UXBOQLfQncPgsF7tTcVQgM8Pn40gI54xbaV11qDjYG/IzFCgixRyBOzIGS
Pi0VkK6wmBBf9Fq8AioFiIx6aUPOt/IwmfMmyvXB6LzqTTC1eT4ZJIokdqvF
NN8MMXCK8RvwzMT3VONUbYlxPKNKvuIhxQHqsXmd2u0pkKkGdm1eUO+GGyM7
KdyZGX9EPRtSTrs9tig1+NtGLvErRcvdJjpXUaqcjsesKaLba4J3wJRoT6Ly
aUJciq0fiY6ii0fJLENhiH+o3B1Qo8E1BSyBn35oFh2mLX590z0b568p4dTY
XNiQw+/VxJPjA1yCqHp3D8Ud60qw3CQOQnum/5lR4NT0AAOEPUJoshmRuKr6
J9y2q6nW3MFZ6B+jkgRdMKCRpnMhFA8D56Hymio2o9KN8HsUQO448tgIJ9Ip
5CVzYjdsSMF8gibiJdTp4dxejOtst5ZWuQ+8Lo09UGUHMJkIcE2LykV8wwkc
lxgKZev6C18E5xjw+zLFwnwxDeqogm96CtyOupqdURJEauntWgIzU+Twz4ai
kUVWfiyTt0TrPAblUAYztfwio8piKcwCCIv1RepV8vwlX4n88QDorjkLWauH
iidFWdeem27kxJlnPKQCegdNcK8gM2KP44ZaPMAasWYu5Ap9352vGYb2eOcS
nYfxktlP/yUwvwC0F4uk/jfzlsePzlWtknfFnAeeDgtwO2xwz73ZCJfZEQFs
nfAOSH2ZP4CeFGuX/W8H0mO86wFTwUXoQWFGKaNZTE7TFwXoYyhUilmocoix
FnO9RN4UFAZ1y0EuDngXHJs1UJ3wiot56sEQDLid0gqVjIC2VdzM/bIojcED
blY221hQ7gZcQjsXVrrHKz66kJ/N7MD+NPo9lVngCMRR9g7l2c7dIi/WSw5X
25J76mFCC6W6OFMKu0z5SmzZzd+/HmHPeYO2BpyUZRjRYarDSH5JPgwiakx7
A47rM6/DWP51tJ+zCOLBqRuuNPmhCBxRvjBiZSWF1vCy1morPaAkEuyps67f
03maA2UtPkDilhfqRVoziVVWnLisjz94hTLSvxMGdSkx9uB0H0EWJOgRR5I0
B8JSTScRqOYR3Q1YxConhaBKxq/RHrHS79yCA0eraedu71MF20yL31tRwZ73
hHzx8FH5dP6UjVb9fu5W2CrUyVL4uQI9oej/GdlidfC5fxrhF3BZFsxsz1Xy
yYXi3wYpdN2HeQWo4+t1st8nhcc6NGEbYNHkgGG/8Nr3jwEJhqLrUZ1SKhyG
HFh6V6IzUo4fhd62jbFuvPnRxCwJ0tsxahN+q/IoTivHHVGMbI0iFl79wpX3
SsMFsHSeizqz2MZiI8FrO7dXOGhPQ91wuBJ4uQxsG+OHoF7iKi2PH1yOSq3o
qxSxBNDI7sEKx87s6hGqpHuoVyoYh8HJwKutm+4xofcmljoCmukAmX26C5GX
d0VDmuMIDXNur9Nlf8LjlqcQFjVhP24ow0MRNHhfaXd9sLC3PU+wpPvp3xmR
8HBFA0IxjPbsb3T3ts4L+xgKj6STphZ0I5d58L2URDPsKclZJtY9Oj50LEQy
RmCtcYC5hb7Y9RpD1zJ1Yc0zBJ2ve4qUuzkxyK+PErKHygauz+N8uZH9dat0
YHFT+TO5c995umLt2xBfpbxD/sW3p7ytJ/brIBBrpw/a+qEUzKQlUiDiHAp1
a1nCyvEJysFtnbKEJvQqg3pGN/iE1nyCPj88+lRzQcOVOOvB7D5Oy5CvFonY
dNwHpO6pXxc2nEswg1P9Lo6H6AWRiGcx34UtLRY6A04xGKIBcdjAk/ROHojL
Ah1LEWc1BhgCu1MTYrEzi8V45oYY3Zak9xQ3OV4/xNsIlnIRlmuupi2jt7YE
eBFcQrMxp+8HkUJVld4EAjKrKsupWqjVh4XEkdoarz0bVzFLnHMJpWshCirQ
X4/gQT4E+9NQ+pLQ/o4ydyKBz9Q29XyT2b98ta53Q/NZ9Y3i0/5jg0WX7XKX
V2opc4CZGnnA6ERy0FDt2Pt1Fq9ozrq1GB0OLtV1kuKjP58od1RYvnzEWRcY
3LWqvT746+v+ZA2tLkKMFaie/PdxkzOfL8gODhY1fvgpcd/UuH4psjM7B+rA
RvHjI3fX4h2XzvQZrinivxPWW2TTmmmtneh0YO/fXYOXZid1A7W7qRSQyamw
dLeWdYFqenhQec/pSMmZeGe+Uu4mULLMm52RcmcQ2TnJWh1Zwk14zDv6Y9C4
VBuBRy5Q7aiqqwWe6rRsZgjK7EF39hc9Bm96BA+/hNrH/ULeOPtEVR7JopKq
By7Bp4jyTSYF/4NemvN1sy7jZCdVzjDczjAwOQeZIUWoTBIuG8+Jc+EV6X3t
TGGPfskwl2bH6o+VzfiE7JQFnBOkWLt4OyPiM25zfO6/hZIk13hj7LADMk5l
iCL6YKKgjC60DlvEhqJI37rEoMFAGAiJtJEL41x5Kc/HNka/leTh5XIPGLwY
xhIW/O9rudPPIjxFiVPnuC1VYhLSrsC2l9sDV/2aIEltY+EUkdV/rETtvXxU
6dbUVwXHwDmKZjnKaaPvLFReVCvjjcb234YDozVc/g2u7mn0lj4ueX2HQnL5
L8oy0aoSpKzJW9+ehLU6SYUTkG50cc3QVpExNTWAIwbgChf1FFtNIJu9l6PU
S38NfwjhFexhzrNI2wdNAqXz2Cpjc4ckocX7HYpAFkfBgAkpppVFHN/W16Bo
TBp0m8DMBWgW2AGjGbh2UX8qBM1FlnPLny42FppazhweO67P6KHvzKmEhUzz
+Sd5MUFOWw3XZypluuPGY+wU+1MlKZXXM6L79rhBH2D8jhBh6Bbqi3z/XOdA
RF9Ks6g02kN8PWMf4wMdfMGXlV25dQif+xXP18jvPVondvhWcK4HBKdVJ4SI
n2d0RLFglmcenBBlIom9/QCgCW9tFOU0j5bef9xl0DpyxPGELW2FPgZCVWJ8
ffGf32L16hE0UtF7YJFELgc7STjK24xfNyJQEfiwZ9aUhocetnAv9LuBtR63
4/7cH++hZ9rw+cL7rkDbGzMm3eJLGdmCSiFqmOoNHM333Na2yyaS0kldvUSX
VB1xb/TXNoJFV1MBY62l4i5tQlDNB/7k7hTz8Ai+nE0eL1nKLadpBHoWzstk
ecGljQS6EkCO5+JMzFcSL32TUZ4X3gXLHRyHMelM7zwZEIKLpoiOWJsz6rxU
Bgs/TyQGIfTzOcEFaHvpXqvfElYj7YN8tihIQKT/Gfd07JzMRbnz9GF9o/nS
/DXLdieCN7aq7gv8vNGaWLvGiRh4/tuRBeBKaUAAVyasBB0THGXKpUX00S45
GHhTETHwTvEYZgX8ncLOvpv1R5okemZ1mrDGZr6PTi71CX/c9V55Xqp+c2fE
4QQS/731EFcQAeLZ9JtLv6rITFF5WdsjLyoWi6JjhPfmzhuQPINwJZscp7Ev
TvzK09pzxM8Poc+/c6S1ksOtkFYr05VN/Dovdg6+a1m9b5m+2BvTDSH25efR
OkCRE79DyRLG8J8WCH/WsU41Lg4ZnDRuKVjfM7rABGQDXEr4Mn9LDaEoShK/
2JsazaC9RdBbbIL2ajD+WuVUonIGgTeDQGlmHxsgFU7lIp0gv8KkkxoQiZIZ
rFX5ZWOZcOR2+gKan6oxFpGdlVvp2dstF1M18mzQLvbzjGX2LLZjSq618kgl
lZQ+KfbAdRk1UJFZjXsjSsm+Zi6xAJURqJPBOcim0uu8K7OykjUgDIGIzQ/E
kIS9+W5n8MJ5GpcV+fcAsyAhEPxecBxLGBQ2qR6nVWfo0oiBasrUWivkvaSS
l0n4ET+VV+JotEGuPPf4ojNutXI5qAe3zSu4NgqqlCY4cl0wbwj1ccA4mGsP
2ixyPnzcZCidV+ZsldQuwHqBlJi1uSCqi8iSM0JLd48UYZxc3Okv0Ymq9Y4d
JCPV3/YF3UW6Ji0NxINwZHascGKI7KgDutMx8wO1/BLqdKp4iCYJR6VXFe7N
2nvYXjdFtrGep2/F+6y0XQmxx+EvxXNMKxIdn+/FKrSmIDBd3kBzbTIupmo6
TXEKIsdBqv370vyqAccAbICGIA05sIo0I/AZr+3I6x6Z73bbYNHbnktaDz+l
U8IGZcM8LY57XskuFtmdfgx1YjCUQyl4Bre3JpOF0+8BRofLeoRO70puLOB/
3hBgqvnoBvQ1H2KFYkebHNnQyAJg51Hdj3T2k0g6uQfD5mffoQasuuiU5Iz0
t/t2dInkQezbzw13N9Qp/3PGBojV2ylx7caNvbetR7mDul0xboQFIRIZyfnc
Hb8TGcPmpbhi4n7MAjQfaYYZF0Ockna/QKq7WALPm+DLNQcYaKRDVKhMiMIA
ONCZMnrAEEV+5Q1CuJE1Me09nEn/uhkk6XrrWblW76F1+NLM0YwwsH3fY/OH
X7Y5hzCxnobg5pE7h1AN2y4CTcXxA1dX+vMZI3+YL2al2w8aP9bQEfvTxriq
B5qSct6762Z2MqJbSP1JYtHZ/uN58XWpCHu0/TRtO0llVcDcMYcpPJLomm0s
+u6OxZ8rUVSj/VKh2Ems0OQ6kwqyK02Lq1Hq1kQAODVJ6hnYEDGD7urgw6mY
wmpEiG/5OURjeGNp23yJUNijeXVPc6/J3r76eQci3Q4sLE8cSJnw1gLwMR/x
gxzFBUPsWzTM3H+tCpPFR9UXilgFu7EaDNK5H7YCf9sG580VYR9JCwXS8lVK
5Vr29UO+/UT2dccFVU239BA0WzzARN6wVnA+X5kvOW6sJgZoIE90iJzh6OZ1
Ffds5O1EzQuApOwdYlD7e0P+QaxOLBfFWtvb0sgEAVi73EBWkWdod0LyTXs4
rWOAJGejqxBhLiIP4XOiGBxKn8vE8+wvPo7i5PESlin1rw6Ju1pBvOFdfKog
bOeHoHXCtWI3/t4sYk4qTV6f7Mkq9ewr0VbQOpi+ig8Q/JsqrfrSHUfE0Gg6
GTvjK/4ac9TVtXKv5fILbwyD2pmbkwpGcaXoiidrEqwFOnlVmJRDQsJd5Vyz
GSsT1A7yPFwMjDJbVUGiX2MqAMqJuLF4szqbyp1Z25TzYe3dVOufZRgKCnbq
bkyvErQGaLA368MYMyrkIggmtZP0jqiY2gNSlR8u7FVc6i0FZZu887LYpARh
NiGwcyQsEDBp077699UewwlEVRSB1csnML7n5xBTo0MK0uKHKH3vAVeAK823
nb7t4W5prg/IKd/84dsnQ/JDdREgtIHa/ydgIHwOtoVnBn4ET0GbkPxzj06w
6u+tqTP/qEY16WZcojSv/1V8o6+j1n5RF1v6cX14ct4uKyMo7lpVdYym7nVx
8mngzhtXNY6Iyg7QnQE21CSu0h9LbY+D6MoPFaopHh+XAnhhaBQkOpOYI8Mj
zplyllxV9hwC1Il+Medml/tC1LglP7Nmx0Ui96gnDjyDkjLHx0CVqbCzve9u
gBvjLegVB8bhlYtFhDka/KC0fT9ZkcIoXykv/rtaYY9K3ffDNbASPHU1gPTV
e7dw/544NAJLUdwBZuOB63FgWh4M4EBo4ohrAAFhO2HZ8OnH0fQlQ9A86YEi
7SKKUOlftVxH7E0Lzs8LmU0Z4vgNlFTuTZlv2vf80hMipEU/bb/AZb9aXnHa
gznKKKOBmqSblVpwZND6Uf4njuDcZqmpBmT82ocDZZsKndVpNeoLgX3oo1Oo
r0G6dTbRNK7bec0pbKCCEIx84QDJej+goM4hiirqcfA5kQysUFGiT0FEEm3w
7bhsvkGORSDpJ4szKMt/iNpCzuHVNVkIwq1cMJ5YlnRlFwRwYAHeelBieBBF
1MphHUH50+EBkx4dHy9HjSMh3Uw72AELcUXR27+ojX9z6HTCL4RGf66VEEIp
SLNb/S/3y6gAreff1NXK6YVGzw3Swh7VjajVNCzQDuwrgn0lwHtPqJeYNsSK
6WqlSD+gdjtpkuyVO4iPcly++zyOp0f6hnG5RznoJRgPwCCfeL0xKa0UPM56
BbgwLHMyTLm6InuWU5m/ckamiUzCLBL7bIMVGV1B0YFigTUeic6TUfbh28GD
LigHeIC7xLuJOezUEXImyd7Fsj9iXj8CMCDIslDjUP4Nuqf31DRYDtQCE/1S
p8FePN3filz5oUDxAPX6RvaNC5JtzGe7/NaCImwiaA1LMRoa1gya0tun6PQq
AVGC1Vkwj2y4g3ypExuXuEQMpvjGcblT/8NXnRw/Q1qi6H6b9PPAx1Y9QkhM
TNQndTPKvzsdpKTZZJKl4wCL88QZcnnJXnZ+86d6wzvzy2YJBXlDM4K7wH7/
3Dnch4thIGCAzJrYKrVEijmA3BlqGTdjTsGGFxRrcUFijexbJZYo1NxpCwi0
l1Mtt/kM72acdUB5uuucvBCe+bR9XKV0/wqPC3sRsHsNpHuttKustIgUZ3Vi
eLPhx1QIz3KShGlH5rNx2QupiBfzE12hH0rBT8uQV9FFW+jj4StzNDIacHZE
JIGDAcrQIgkpHhaE4Udx4LQrQYdzZhmaB0lHc9yZfA+KgDTw2P88Y/qgXf0T
gxl6zBsZuFJoO8TGHMu5SbvMydOYeYgsxBJT9Y+tGOwdR3PZJHBMoFW/qPiw
HtCh2iyusoWo5dH+HcPSfxsMjbDfss/8OjNh7KxZ1Az+R4S2zsdQuGmvR6y8
ppYDy1Ob1Yaog00Q01N5QAelMItYoPI8VI/YybUQgKa1kCn9Nfu6HetJs9LZ
PzHwCuZn1Yaq+rycpi9nFRkad6xCsfNQH9qIxWwC/GTgKh8TK1QskUbOKuUe
SRjzuSqCa5264JCdlYJXkY/3hcvOTdHTD9FLG47KiuANKndTIwh+aTVLQgmh
RMSZXa7qa7+1BeFA/5FhyiVjP5ZrjM0NCHa8xOryjEVmASJMDBvanEb35Ik1
NS+UohjO0OS6K1lZ7dG0Hj3/muzmsi3qRlx7CgEpaC6iSShpXKbqyrGv4aGI
0okk8acW+37NvoeoOX68fVLQKKark9qV1+/mhAgk8N6RVqUjuEfVaQNK6ano
jJfMatIHdR1ilttXmvzPrO4R2QiwdXvdtK2TVRDB2kB06I1S3V2Ev3OXabGC
1HBOXOHYJSndANwK6I19M8ycCLOvB+3i1NjkhOu/GzMe0JOwa+GQwmUKKbP+
b6VNHaOTYSWEcC6JCwIVAqYVlpWsQ/GzzDjTNFSwVAgIcL1uLk0nZg6t16su
fUiRSyjjA5PIn6riOaUh5cSy4DJ4pP1KFB5k6va01Oti8wyTH3WauPSGfnb3
HuYAJBK1BEXIEjWEMZT2GXxeqZNUGHUD0AFgatzGWGNNAgphwJ09+akmgfCi
7zbXC6c0dpmuxfGNnvWVhk0b/gxnFw8RvOLvaFNSSSL1cZQiWwRgQHWt3RMB
eRwPmWJ2CcaW7KgCFh20hMDnNTdS6XOaWeuvohAVjvyT5Fkg/Zd+COGGF8qc
09qZ/en379U7956rJCusSa0NvmbHjj8Bjz/CqhFwf/2jlKwUuma1awoRry6+
3ziS7JPIBjrSc++7p8yLsO/y1ZYZjnwQc94fz6yFxDZ6tomS6TbxnLxWE0vw
9n2MUhgybyrdBDJ9ymZtPSxbNdMQIkjFnbEZ79PWnooL9bEXKDJ4YpOdGrLk
MgpZ+cxrxCl4j5LkJOuI8ftNUw3cpRRNJgsMsBUk9nqfDfsqG4PtKkTByY16
/UXvMaS+4qG/4xsCFxx68apID1JrTS7Fdf56Xu2DJH9XWydbIIl3BGOsiyTH
UrHJxEvnGBDJEeyrctBXbqo42Q7TrB9zaT9xlST01Pm3M6RbZL17ItWbQuVU
MWLZwZc8AWjJauK6t4vBSVj9KagpE24zoAe0g7VeixQOriayoqevraiMbBku
pqoucb32iwFBANUYZoAKKj46gfqxeNpd1pqF8fN/+HK2Ta0rCGwkVlXTtZbd
9EX44BXAnFCsZJPQekBwnphTKvY4C7+sI2Ejh95O5dIUz7fIiFU3L4Eh3q62
N799ZUOJrGaYjGuQjp7ob8PkX9JGCIr9ewqgZF+uWNrfmPlkY3W32W9ZHYFs
vhdraTvwpnLQHlNRUYmwlPHN/E7ivw3mlRAaFM8CKvxyElfMSidNMBUmZq3q
ILLWU3L4Ho6e1JRr3RuhIXzmbp95lLAs+YESm6tlVbgvKNfHGr8TqMhDaGn2
8/ACa3T1F1BliBk9jhgu/0axTIy4LqJ6xihzwKkDnQ9TetnYBQ67Xq2T1/+W
gm5zRCTJlBNeWfKfdeVus+ZH7ZqpxYnnKhoqBlKIGIDyfrzooWu3YwIz9yl0
wCJ05Fu/TNoQ2BAmMHm1075OKvNHXisI5Mtq72vHFijSV5Rw4CGr5WdOo7Zy
LMaggRQsfY1VtDFIbjEYXMjD/4DmOjHh4vOmGQha0G+bQ9NMK+aBxemF0/oa
2lx09TXIWbaPqKXsZS7SqUU2pGnSzCmCqvaj2hqk19nymE6rwDOnfaVm8ckw
w1jU4nQPexjbX6wdRY6fuIcpy+RgUuhe2Oeuay7pOXpMnDG6No8cw6nRvuWi
s9wQLy0UoTqHbzVputdTfaIRw3KrqOqYlzW7L1MluPBvHisrVC0CrRjrZzyd
RVgVXsah43bxCS+JYzhsc2H2RvSfdHQ7yeRWcMVS8v3DCG/7Q4FXHsdbg3PV
Muojkg5zSqv4RqYccBbhyYBg1OOmIeVxM18shlBB/C4TOGc9+rFx1yhbGf2W
nhOBN5yfIk5tidJz24X6jL7BDbUXg//H2AGm6M6j8+toN5rd2Dr3zJj6JrH2
XDgsrOnDHpinjXEWh64PsFUTgWTLEEsSs8ofX2lzfN8KN0Xc4l3Sc+83TEi3
IxK6ql+Ax4ZGa1ZziUMtjfSfEyEZ5nrfaVd9n97e2FeQbKPO1ii+9cqsgyOO
6Vg17NGVJ5/v3kz5Mmtifew2khMSF4SmXPhgMxXforRz5BP0Se6H11Y4yMke
EBFWEWMQr0avmlzepJi0zXXcRapRcF/m/u6Va/gmuNWXtzISI5FIapSjoQTU
HP/ML8mk5nkOkQxZ7mm6GNphJAdma9+N0GQYrK6wPYWwuDVzGjzCi9Sebyvv
yCHnRcyw/VD5ks1yeBLCrvOB9weK1lPOY2FYLZaNEPKUG1Pf05yGDkj+e2Rb
QNXj/+pIwfDoDhhDGPQOBmOLoUK6aew8SJjzfqcDvKZCfYMJP4HEj65Sfbbf
tcB7qDCg2TmtBGlq1XtC5TbQ+pYhTH62rOZxUj1fnY1+4Hosklfeb8K7Lw6E
soElqUZt4SfBYmMKRKv2p7obWIZcrBK7v3MBu7h7gaPF7MHhmOxSjo7WTu0I
ic/PJSW2mV+K8IKbf2QUt7IzNwAzBAMnwWI5HKBLXoWrBRJkcJUVqlOO6/zt
DXqpumiz5QvSV2trZCuE94CrPfeqi4Ds5HLl5keAf86F2gkIC3Jxd6kb9WjJ
hnO6QqRKZKvkpX4OMva2CJ/NRZ1cErvDClmCI1UtqQVwROFXuzzqQdscnIoB
ZP4Pl1s6q3BB1M1O24Af1ATI2Ml/7pVDwUR9xGVXld4iZ81HK1/Rtb+YBWO1
mT3xmP0L7/0ROhq3a0DJc3I2YcAy8T7wweJ2yGwVYt/Ao24mf+QpgBq3MC45
9zR0rQD4cA+uJZCpSU6pHvCs/gA8WgmYXqejBT4dY/xjsKzQdeM8OQwLpp8J
hutOPZLNTkHhCKK6xEJHzGcq3lgPWv4WJ1hv8pIML03emTKdx4vluynoiaLV
VTRp6NXo7hi0WG3rB/migczavf49akqz/LnGT2G4feAvpkaJg8eu9tO/norr
m+cIPW9nFRGg9nA1Wr/szG/o3EmlqFaO8zRY1gVwHlbFxU2Ck9p7mQb39gZ/
jxouRMebypJNF4JjNPbsPFshUJYXjUCakuJO54bJqn91a/pD+IZhejOU2L6e
uxh2l7QPiKErLLo3QQVGohKju3ePm37ad0oSHffeKUEURUaLUwLKrp06jcGJ
Mg2uyYL8l3RRwJaTgS30lySu+aEd/Z7DYA/Vm3u3eAeM0EqFudNJg9HA3Acz
nBBjztrwYSmcDqE2me8bKTSk3zIXqwfSOZVwZpzTDHwoefs6D76E24Lzclvg
VbnYchHF0iGtuBF8aG3lkZF6OEbeILnCPHeyxdb0E1P6d3wDmgj6Fyes8sX8
5huj5WEbPUjc3RPkuskPjFc1dKtxGMSlrWy/NtiCz6IIj62ZnkpSCSTb4czl
IuJhysuTDAGf6+cYy/yM8/OqJjSoUounOXYLhjUS2yNupakgfHlbh2kzvNm4
HfKbC7Lqxq9MLPKpbDRtp4YbPVa6oNRQJA/mw14KLtgnil2K9Ir1Bz3n2njQ
ckn6T19LVPQsC0IOmWVwa25L66JzHdq+bETd58sIj2susS8j8DMqhd0m7WYl
0gu0EW8V7WFObuTP3gnpe22aygrjahsTU5B0M0LZbSgCw8UJhMmsfs14Gcn2
HBy6bejvInL8Mr0B4W5AZ3BrLW5HbBiaMN1cfTjMrSHmIU2A5APFg3PXt+8B
rFgdfUleynWO2oIZWO6KTr1//Ij9QxQ13+53HrQLor65m1+8m1NBkaBS1n9a
rG/AyLbxIfmt7TaUCMdZvbHxXMswk+TLnpzfgT6goDkMg8SJAoAIu2fGTrmW
AsCzvPheQB+WD9IsgsiTg/BSim5CTQm3JRd4YdzUsoG4Io4IyymY1EaC1xM7
oQPy3YH323WNyslJRLcuipau4wV6/aNY/XURIgQAPrUbt9vdUekUyOqeENRJ
9viEI8JskwuVLGwxNrAH/YXDT6Heu+86mpVSeOUGz4/toE1nkYLP6VC9VqfB
AMeTpEQab5I+xLgh0v7BDwFuiGU+JmQW+xpjwvcIdeVQvqjw2iaEuCwopKqe
ca73mXZOt+WkQPM28/3fR8NBz2QI45ndorOSukl4cPhtBZ1+Fdx1rMTsVpNQ
8ts+zn+xgSf1O8sEaJOOn/jUQ+u4flvtTr1rBR0j6e/jhhr6A1PgA/fAOYMl
kV9PCd5QricSiA+k61KfUNVbUTZwzVz70mWvx8+IrzlMnorkHmaa4q8UUsFj
+nK944SUMYRHy+Y9qs0M7X3jG70iuEkcv9B3WD2j3N/43ZdS5dGGrhZQnZ1J
42jrV14ssO6t6VF8MTJg5BNsuiApQVjWnSza66WizzpEm5rWiBioC3LdkzZi
9K4PDNg+FKQyljgsLjIPrvOtvtfGq6MzflmGax5Dn8GX+XIAvBTtY6juhqPX
Eg53iuMWXLBaFQnG2+2TNDPMyyRPazrrjGe97VXv235CND2YouBTnxLVNA45
nCj4WpFbkr5wGry9nkPhvR2WRgv6wV6qI0HNuqiFxFfWXWfhyUcq72xXfe7q
qnUOfUdyGITXqnpH6k93001im70W/czpdmDtnjuifN3wlZqHkgIjyOzptUGr
5bi7S160L15TH3t6T/Lrjo/+Kx9MB7O4REuXekft/LzkZuAxT/07Ij0k1jgR
QX2V7ZFHQ+fR8OPg3ip6CP7hwX3wKrzelnKecUgtZEfj4xApD9LjCVzRan5r
1QXnveaL6TeBp0TEyg9KI4BhpqASD2R9hw1/P2R81FyQ7T5+OhPTszMWO0AF
3bnEv2ffLEn9RcC+UQcw1zCusIbQ5v4lLmz+l4ctxDclYzeu4Egv66RJ8v9r
UpSo/XMacIhD1qydXuaN24/6ByE6OnuYk3NQSdltUk1Wd85VPKlVsfnAcevt
9jRzu4+8p5LrGjLHpi4SO0x/sgFq4vVrr0ek6vW7HlzhACPN3nYrou76HMzk
S3rAdSn+UuFzij9Z6aa7PDBmKaLpQivrFI6cSIbVfxTi+agdHsDlKfTdvSXu
mURwlE4otwYiqFHQOmvNtKdzJtfB5hqtxTnA+G1Ttb2JfiBrMlYjaxYwc35o
dCydTrBvwTDuHOfBmdC3tIHAZ3rYTEc3QysBhkairqrtLwCzyWUeuZxki8jG
RtgPRlvCa/c0Fe2MAP1cKyJJQWwvBkZiPX/gRxc3GXXXexq2MsAZY3me/ZyL
Ghlg1B1vFywjdthUXx+GXQSBKo0dktKk3p6etY7l6ojOW2vNdwjkI8YMlzlg
LSdyspHBTAVvSfR3VCuz672NEzBXQhSoAa6p1K5ro7Dg7yoNBfQ8CYS1TZlY
lQ/OZZa41Y6IQbIjoP/RrJurxpl5CbcCmSzCXiABwKSyO43TKDuT+LjU3QJM
FJq2nOTduODXVFQNevHijJRJRmQZQiytE3vxcBAi2tBvJtHl+ME8SwkU6BPl
q9K1sZJUOAiS2Mk5dl9AE4vVfxAH6Z4eHet9OLpZqkrH5vxfitxY+LkIyTDT
cFdtT//YNyxZVv8Rd58qvFmgJcZP0efeCgsS2tJETb8QL2BOgtRnS71xMLTt
vgUq/U1KKfdM2J+DGGRgPDVDb8Xh8Qyh+S8PCzT/X1jX7eFIjHAjj8IVmC3K
LsKWex9PuEqQc4plG0NEnz6eNmBvxJoIiB9ELLa3bbroSklZW/swcToiY+Nl
YpOT8+UuJ5FGOUAzO3lgxlbxSuYJXfVs3quIMfT7e7xnS3vVsWGC6Tpu9HE7
qMhzjdSnBy/XoPVqth/hJSCCt5bpNoyjpYu9EpEYz0KZIuZyM8JtXLTAf1jC
2R1/vxUuroKTb8EHe/GBkZshzaG5YuH1gq4h9bQUcyjSFBLjLHPSHT6snSJF
KRbBcEqswtXYkeAo1ytjag9GDpgObsDrcBTE72RrvXJX2K4dkfs9U/1Qe+yD
Xp/dUyQq6l6m/kqqbZR7VUBBDXCLQsHgM2GmEajdVj/q59lfg8LrnRlFbqaJ
I+ZkBi+gzSoJWvvxLgNSYwrihSoUWfHkPQQV7V2Drqp0D2nIS9giJkZX6N4/
9K9Giw61snp93SdQiZzpJusHl5FGwsqOhKtbxjSfVPakNGfLW3UJjWon0g45
fm6lbxP6SPeOMiW2TORDu8yPYFBZPS2CsK2Vc8R+4/BLUvMTNsNHvpJUMHLO
5Iwtme/Jq8bH8au3VpIVF4CqHw3SHjLOS62yZiRU+XO2v0vm+peOhAm2aDPR
AQ/bEf+o5vT6+hQYz/3a0j5+EhdVrXFY5lnlbRZHztGKf+R6lroTv6V+Fugm
5a1jC9s92J3c53uSfpj7n1OUPIXcJBJmKiq1mIYU1NUqjz2uCN57TN94YWsx
aEyfA2QyecLgg5nED4V3Hi0jlkHxomeVj1tOicjqbHSduZOe4t32AQJGrbX6
AbiWuRgE+XP2EhFk92uViuWrH+V2BspVEni3QmQvdsUZYbhPjrQqMorEUrQl
BONam+Tkse5nARRbYDQJ5U1LviBhjf7+b9sM2P5THNSEfgQODt3iS2vIukgF
1YHpZQNY9iqBw3BUhmxfsZ9k10csb9U73U0ofx265bWAJEhnry6Xd8fh8G73
6kqwrYjszJQ6Wk5Yam4gJizTNf0FPxRSV7Aq9APEZnec8O48SHIpTSqX3z1b
virk7zi6jyjqeObTtPEMdCW/X1Px3TTcJwiVCLJZMT20uOyBehALZvOdR9mJ
Zn4F9G3WqbokcREh4TvOjihjcO2Ak5YnpggsucBU9Ti3rwSWFOUnr71PcZMN
nA8L8euVjlUG0zRuNil9iw+QBEJFFb3sWC27g3vpClt67drM/Oz8fuuJJhMw
35CMhCVlcKCTFfsTJJOnbaRg/QkYGCuF0/xDCNO2jOSRjlZDJI2eNKTD2YCm
6ZSdEl3HylpHkJp6vWI/VbQDXURLVyX5bGvQ6oiv+21Fi3Lu8r+hzqJ+0ag2
HpnvpIf5ohWOibTGu2vmqntGb4XFXGahU31Q9yRNSE/cnf9ViRL7i7e7eVlX
ZLP2LoLc3ZTb1yepz9VVa4EZg0MNAD40QUv//rjuYgHxM2z+GFVyp61fBwjK
6sntiPQXnd9V8sHbiYsjvPO31rppWBGBv6uKaSko+MiRlBgVcC3kQFQnz/K9
Q3lwC/17tPzGBz+e+f/KYniqcSOZcdTx40i9o50+oGpUJvT97Sswp/YsAxIv
9XUAdfC+BlOWxSixQqJp6x10BmbzoWfheIbLQ8hqxUEE5LDl+3aY1I+8GTF9
G08GwlZdRBAbZxNCG9bofItZdLJ4bsRirmE/oeIc3bhigD/uaCJgCa4GzCtb
8y/gbUE3no6iBbpTkPgexn9yGBJ8ihyQRhJxAPSEfM2hqswnsPkZ5PRS+nO0
bCHf9aHYEiNDewCGB6oo50lyJeNxBVb7876iYHvzFI+5tRQnZw6U5GqhFtwb
zw+UduYT/kLPiKXcOCCf1pjU59S211pso2y1zuWdadzzi/4B81Qre50ZlQDT
8FVI3utTebTCVdxackMqh4uBOy+FhWs62SDJWUYUnwaDW5Nzq54paHGuYFqf
1Iqloo0WaCa+kquH9pXQC3Vk8vMP8ENNzcj2LfpuBuep1EVg7wB8MF6c6f0Y
e0/G8sILA5nf/8ZU0GTj9nR10ltynmS7y1cMRRziGiUYiDWg7uNRrEZKNaaE
Msxs/WdkFoO+HKuR8yWriFahjFfeWdAHQ5k8gztocI9Q662Zduyqq5u1EfGm
RImsEBq/x/2BgtVHNC5TQUR016MHmBjj/SxiXTXgDwHHL/eiNs1S7R5M8qO4
V0JxJJXmz5z0PnwWEwwKfTd/Vc7Q5DaONPzKk4CIUmu5W27R6lm0jQiu9LIh
QTS6thVwue7YgM2c2GlS3v1yZJEHt7zywHDW/cYCWoIkCyGaefEKAwDhs4FD
FoNg73EgmcqIi6894ET7uq4/7d1+Nnz0075yApxzXOlcqMGxhcwl4kIJlBdq
d8LE+2cf2WnvluwE+f9IEUZaWO6a7+x3ntazd+Bb8EAK5cSq8AeByKyUXbos
nIn2CdfW4iywWdaelYzq1EThJiId0E79wVY5GSCqPZJs/eUJiM/K7Peih4Ta
JhFxGZEgy4Rk4hcrIC46ox9jjlCAbHakORO7+uJ8nDvNAFv1WPmgfBGyBG19
kHb2FGKXN68QDq3YPaFPsyp5CwVZKfAWwNETp0ohzu6WBQbbvOCsQfI/KYyQ
Drj2nJGWnD4ndR+hUGr8FA1jrGKthYqK7E+uUrsa+bwhofxvovR+DJAUSgWD
/zEccV/i89+QwxG2mKqVwz6MyKX/+iXgveR5cMqL6W0ydtXafI2dO+3cqhAY
Gdkpd+bikoRnYA1Oe92/PG4Oi7yVT9mymjXVLb+Ctc6zYyVs/3FtCTa3S6y4
h32X/Czjh91gUBNKqcegKWVtFVv39oilvNSb1wKGaW+hgiSHBB0hEQ+jka3f
w4x97pF9tHQU6ALZHg+b92e7ZLuD+tBsOXsxSohkjpqDmLmHdgh/pUcXbwar
QxUwGtcTu5TQuFVpW06HnVI+zAcGafN4YZXyxo9YBMPt+qTHr6YPEhSZLUkJ
vPchbBzVmGEnt3ag4bgt4Wh+ni85yaAtXzSmApEOOQZg3ms4druYRgCXlojT
//TV+uR+onECVRrHapF4hal0SElImcYnuo7gaCP0SPgoCNkIrp5rKjibQT+F
TphULe3NqzOGx/IySoQ8TEZaB26xYoMxIBFA4YIdXTH+AxsGfm3+c4BMLqrV
wzXraa1Z5y1iZ3QMpSZATvYnrM7RjZAyg0WslWJURbZd6S7MjN9B74glyK1W
W4jiVzEGfPwW5AZhT/wuwFd7UA7tH8rT8uqFl2ugqwJEq/t5oIjwYMHFC3Nq
IR1GJVloO0mywyj0W8ITqUMjhSxubtp0P+p4syd5TTW92eOfKSo6fUi6RCJ2
XPgYC+JNGuUAPsuoN63tePjRdIYLmcv0UnKFBYEUir0+gqwWcZP27/lxQvXa
0cCusgT0vEG3WO2HdJqEH9PebdTmvaHy8YhnB9ZYi/9D4mJDfawDytwsejty
l5ObmK/T/Zx/oVMZqQ9ZjsvQZftD6pZ7CUQjkgECTmzrvWsFraks84UxELZ5
5kCV6kyb4PAMYP+n8leIJx5Nqr4LSd6WLGITmfnp/a3D83/vfaKNreQKtr3g
2GZFwk4y00G+ETvA9/NO4wcBV2WIMb6dEW1z7X9JbDIPNy718Atd+bY8bfp6
NqLVjBsfxyLhVwpVYBJ6JDjyZfcfznER1hvdRUWp/bfaDZdQmTyKmjZxWGek
G8jm6Ev5nmGCr1hLl/neEDCYuGgmIg88qu4MOhVspIp/ar6f4j7jQ/P2Nku0
dsc+3hThf514h8iVTpVC7jRMkCrQDIgqA4P7llhlXmNlZgW6S8p2m7QpMi49
JA4RglOo0q761Ao5FVWgCnVLZLwhrCgDYk2E2jokrK8pviaEBm5sBs/YyhAn
7QAg1vAREHRFaO5vhzSTEzbSxy1I2UnHFnDrXcr0cMk+7xCkQJTNUnBKxs3N
fTGfmmg4ECZmL42yXfPgHhXG3Gr69WO6EvAG0vagqCOY0QlHJXLb3phuSFTf
AHCrVIlqyYjkU13IEPkRErS1h2uIK08GKkTNFOYR7o3edsMCQULG44tr2eOy
lmii9AfCksrilWvcUfGfEe/XsQcCWr2/4u7HsHcZt3tmBENjxxpEJIbMb0zs
/v1zpa9yPgNeBWQaL0E6iJUR74vvF4NjQzrJRXyzzbVvy8EUUnGwQD9XNhQh
1NkrxDVskPkDrpYyzeKVH4+wOrRl19xTNVpUdVm1Kn4yWNnMDFDprWBUofwc
ajf/UbczdUpHzMKGuc/5au+0db4SBnN1bTMZyR9is5TtunKM78C/KUkcEDgQ
0AYiQhOW+S0vvMQ73c0m4NP6kGHGa4FSc3+HptGvb+8pBw7mZkwoq7sW6IxH
e2tRM9/RI8fEyLPiPCtP8V5S04P+6PdVArgGFt5SIATXCv3rhhR7VSvvQ4HW
vFFYYvkaO8093+h5z0Ix+Gq5kauJY/hEFOtGV6LMr1IXTFLdgHm4mVXUM+gr
wf4lf2HVPmqc5aQnqEChUbA6RUZktUgvxSKP+MxWKP59ybukMIqL7Pa7pYM4
9kQHc8CNWXbHrTIo9kGiRYmtl8ciV1oPqqjmRGG/HMnEaIA9erB5m3WyDKYe
GPLSlgRW8+8xCn8cqOWE/0bnhEYAtNk1sqVW8B+9THAChBqDHTOYBU9xUZL8
XAuLTp5sDQLhwYGP4gp+UTzhDX/0WMZD2htZFa1xgP4eydd2AYj0AkFNL08d
yB2IdZx+KhVAcnIJb553uY2vxk09WRmCMYgK4uDSrjIlbeMqSEKE2OeQD/xI
32npXsQq5fLUElm4F85ffezs2yCutrCXLb3aTouMule8tef5JJVS5zOpv4DY
zoplcoKEMimu7K44zEsT2Xd4ukDVn3C7C8MkwxOofnr74Q2jVHlwRvYIwtKX
qMf+AUSVO2xLeuc4/NOCqmUU0/ciqk+LsBOvLGIWSRDdTeP6rpyaxbEXwumM
bJZQNDLKK04JfM/IQCCyIcQb1X+jfgJ3rA3vOwjMSmVWXPqQIZM71KQc1V3g
Xi1sAJor5iS/odoEKJeW+GC2ilT1e34+bBUYjWTcQkxIH3N5m+nu90Squ4II
ASGiYNkhp4rFzpuY5YSy64iCXXdjf37NRKonjXmPY62yP3gtJybVGPdBqUKe
SkwcD6Bi+ARzIUdvHJDRYTUGVykgmGiR42g8ykwS7loL4ey8Fev8jov88K9o
bKZeK4dgS8ZsasiPTRdAdYVSCV4ssYqkXkU2OvlaR0hQrV7hpLQdpVpeX7cN
XZLqz2u0cGwcT7zAYoO1oS1ykvAhPqj/DCeQaWAhupuMIuFRKFpTnaYb5JTd
RIqj46DPbr+KRMzYSE+7S3PTgPyO5rxgX/YMoajTMvJeuCC1gl3C9Q9ofAau
nJ0BunQRleVx7irY9+d1LvLyCnCGHXgBRqnHD7d6ccPr9SBVxHoOKifs6lV9
x8p6ELj5ILia8/QW+hT3Vq0phZeVTwYF82iNwKN+drY4FRLP7rO38Wdli8rm
67+WyBcPgyT73ESs7LKDq0cvHO59baM3L/Aqu+SEY4PTGmmEANe48WA9i+Cw
e7AIX0cJG3MtVx6buNAwesMrqIul8rg7eVGPEDE++6e4m2kqc255BX2bgknM
XTQMEI2VSLFkiQdAng9HdftomUWz5UJ67osIWG3t0CCOJ8ggivrR+sFJCHEj
2GZJziQIpRPBdj/9bI4iciniS5ZLGjCHL92lm5fAg++J+1fIhhGdy+60uGhV
DZyoF3QKDsaxKcjrgX+bbnifpOmnRxM4yZBzJD5rRaBD4xtohJQmd+ZlHDsS
ft6CfYnx9+10WBGkisGIRRugThgZOuLR2tW9bAoVW8FnYmL53Ek6DcJLmY+3
6qOKEuZLIkf7cboSrapEPWJ+e6zf6qAxXPgXNKSISV1xDYVUB8iHcmBl5uBJ
rBXE9OVO8ItUuOO5gLaZPYaetSxt+0jznjmrpJBQ5WZCQfD6rDuHf0Iw3LE4
3r1cVTD1KT3DpGOkfsLcGAl9HgMDz93tpXNPsd+yy+ZIvlDYCJ2/AJOkW3/q
PaOYvIDL0ryEizDhjAovDgPtPdojDmTiqtjUEkH3At3o/0epKuZIRPIQOcsE
y8cVjlzURywOfks+/W39Pmz6v+q1W9L0HHiJYmlwTSpAJFUE8Y4xp9WlXQEj
eUz0/D+QQUO5WlNG7Jq9jNERSdhfsKT/rINlAp9WVWWI/DN1lU1sougVzmwN
n3pd+HckbmHkuAloovdnllpnV9M2SliSNRr28f9wf2jC9yV1o62YECVjGXvA
XNKOjO5I2gwlW4yJZCll5UdKH7G2TOui2qILhzbmJBCAmdNboh6ayL07CB9d
npTJTtfbR1ml97Keivq4pgU+CVXY70u3Gde41tNO4WULl1bLi4xFrjRna4tm
01Y4dPwGbSRsX0YmqnWgZuqluBaiWeuyZIX3WTRCzlu4NejJdo92/iXN/tDN
Ezaktqed2BA/kY/v5F/XOW3eYxwZcukn+IpjbpgZGAZK4ux7GB/0TGumju39
oT1ToA3iCedaY+YCrgGVN833f8HUNwe+Xm3ESjIPqKI+gBV5yt/QAsbKdjwo
rgBGHAEIJeOAg5jlAj3v7YmK3ZI44ht7oHfxsouS2uHpPT5EjDmE+N0b2ivu
b9UHh1DwpVULW/k47kn+Chrk7iGP05e3n1CytRQ1pTs6bS9bNv+yAwdD3/21
Eyqui38iJXvoekY7tIQu7qusVcIxpmh9wOfIk6gfTtsgwIJPlenuNnzbjFm5
OEQrksTM7bc6Pq1seD6ApEyZhZBYBbGRZtfKiXvGdL1wqAJVFRCA5r+x8wSp
w4y4a9NJ5asbgJJouVKgEe89WkUfbrKGLpFL+JfuhLnjJ/b3FINdAGxVWmul
TzpKT3Z0xEpqpdH/pz8vm/ekPBeh/P5GZF8aMtH9WhFudzdNlTeQ4xtpRRg+
sSuavuwYfEGfSin6YaUTLxpbm6Mh2s596i2i23u4QVZ957nZvICaSMs40OMt
O3RA2KrHfE2g9xm5K3Xi1wFE3lI/4VRiYQEwITQubJ7s48ycQO3AJHKce4pF
q1Wq9rLoppj8MveV25OmJEgCouJG9StxdnQTi+7iPlwgN3LUtqk0fC4EsW2/
COZUebw38fWcihApnz+Ikc/48fmBzpElHTfenfOkS+BmFchbqLIA1eRSIwig
Yc/1UFTz/CJcdqes0vtUnceNDugKcWU0scpmOqAfdETvRLOFta+xwPt+WYW1
5CsMjOCklruFPKdsq6kf6rLZF6zag0iMcb8q8xVizgChHczPhD9CMuJcULP3
O+MuGM5V2apzfC26ZvyrdRxt6WjHkylY1lk0mPzKKqXaSV2rHPTVzIi2g9Mb
J4OfYx406cePDchsIVG8VzqzBkNE+O8Pb75f5D8Hb/Zsdk8ivPbhDSZQAPsf
QvymvDu+95JBWhFVhihaKVcWlBcgUl88hxdwQPWUljpckMwnmBCyxgJE99Fh
enmsuf3Z93LgiZzrzHNTrBJL13xtFyVnOHcsj6VBmBmT9c94Gpdk3OWGRXZx
9BQl6hRFOOBd3wrz9xRtgOIke0M1IaA49PYjxHsBo5G31pFr20eyzZ2vS48g
x2d8QUYX652rFAPmCW+s2EerDW0H+VvyWnKpObpOWTgXKzIusUsl7pV2LnsI
cOjquqyyxWT/e9t4DKkDBMGVmEZ1P7wN/Zvu8Nu1Tr6bf4f6SaybFx0vJ472
kGjj4lDSAg8boMbLRRFKOQ8x643sEgafeTQBrA2fdrKAwqmS+Y6fh/AqERli
zI6E8SBdVWil7HGXrUxHKHgC5WLNb0WmreIPpQBvrj6vyBBNX91Jh8t9goPo
DkuuHwhJwle77e711kPr78RtZzs2KhfMBTKTyN9G838WpLAPL30+NQAzHP+k
IrlUdy3LEitrzlKNgzb4LDa1dbq10xVwnjAlLBMGg6RzPenhh0UQhSsPSd5N
u+mHTTjKIXRZYQ2qwgxcyTT7sKbH0oI4ogyGk2/RwVSJ8kNfWxjQU/wnpgha
aHdmoQFNLYOuV527344bOp2LHHhHTCEqygcj5y9mZx9lwdW8tDyLaQ9ckncl
yhha1/x8q/GvYaiI/J49u/hp32vLEKLoTZ+y2dfGgug9J5YqLFJRd/H24Gqo
GSQkRjHPdalgpjDFsan8pFXl0IQok0XvXiKsGdUbOKnfk30C+Wlg+CpEesdX
Vb2NuFQx8YUNxo3ScSHCLx9UcUIzILcOpCxB9laQlrwbYUWXdns+kJNq4byn
Dth58SQXWl+5Je2z/lf1GFUl9rAXbaeoqmYCTYWhEsLsHNLCRhwXrls2ZRR5
LOZFiqUw2EFpxbBFVnkii9OQjkzYSwPTnMljn46O7rdwRzlIDwKgMyTJ6yc2
8GLt0hsGJl1pUvEwQsEXPCgZIB7AUrBOxrAYoFbft3Lz256fmoa85l3iS4ba
iIa+Nnq5WHwXrbnpqYs1MaA4Gm2getbv0MtDl0qdSbyT+R26YZsow0Rbw9t9
roDvoyRZ+qfr/CA/HRQCrUfmJfrxOlweUVX3Y2Ey0VEL2HKQjBpSHN2dSXP9
tWz8U63iM6sOwSSdiGMxrkE7IeZXTWDmNl6rEUCBEeLdiKJ/PCL95sl552ZC
vLBCiYPW8HWRhGyJ9jyZHokXOIf4R8UY6dwxZ4GiZgvagmBr+IgyvxxaJCgA
Tw1ZAxoFdkdkhsiX2U2ULmIdWWdcFQXYzhy5sx6p/CnHCC+FqiEDEWbtHACR
e5NVjhNlcYnSF2RnNe32mTQ7Vko6muzBRuCwblbGUMEwmgXPB6lVoeuLIdn1
+6FCrS4trOQQoJqnIBWw9gUd1WZ3a+tlyaNybTc6YMxSOCpUDz7yQRfE73Wf
x+um+5log71PMS0gu/0VabY6l/yBUsiSlGXFv0SiDeN/HfR/fgGYEmPOT2Ul
QsjH1lQeL9fjeWxg4fCg2Np2FKKDOGWjsNZ0X2B3nfSkstqWQMdLivRXQQUY
tTAYOOsc2Hx9PtmU29rubvkQcILYouSiIjSARNrmdA2B+lJERfaclc58lmBz
3SrENSdtFB8k/53j3/3iFgOqhU8yFiDvzqoJjxmkmheb/xsKVqwpe4xEZ0B+
yIrPtiPmaR7b1S1HXA2H+4gglrifpXvshONFFZQIsXH8bwiog1uvPAGPyniH
m7XA2w6ywH82siTVSAa7rJfDCpugZTGVXYWXzIaiTg2mt+4Hjl1nO4tenLYj
MJLWX0pW4lkkpQ3Txu/XqlQGf1E1mJQWoWOA5ionE/Fz2HOHPjQmYxthLDmj
osBlauVKvQSecKyqIdg/90ScVQHYEOY06UGmDzUwbGZ/Cgmu+L/1wWY/WCsg
3YiNs7ueGPhXYKuvjzu/VYFV2HaGMYqZJOXZYfJSywn4oE001rZpcZ/DEQA6
DS5tHsmuSemlueu7lHfF24sd3FFXPNC/OonKx0rGkMn5kqoQQ2GQKlUvRJba
AckAlGUr8TyS4io5hlq3QaGlThl3UKApl1fiEFyHlQXTr0B2fR933JNXER4e
2DKPMVFoMQUrTROiMg2OE+gUL58apHifDczkEWMf4NnCl5UawNNcNXAaANRS
llOt/+lby+pm+YQRC8dnLYwAem90IomBq8EPlTXWR6aoACBOdtLsyIUi1Y2H
2QVFY40YIQ6dHZeBrjmD2nJJVjidZw9d1SlQ/r/9BjH/J8hwerfWpprOUD5I
oOKI44HGs2Thy4rj5wfUsmwwdPMPozmUJeK1tdvtBVckgVnknP/TnJx+QD5a
dhVy3iCvvAxaBMvFX97AjkFbxpWcY2ehTk1uVdaNctomZr7DOq0r/+0F5de3
fH7tdG0FsEID9E8HqRdURNYB85escxHo/LJhbJsk15TrNxJEkXaNibbtk2Kd
Lp+KKpuhNYfNxbDqDInq1rc9iZzGCzc/ua+AdxJqzAdhpoPfTO4lDKEoz7dm
KAT167TS6Wo11z/V0v6YuLE4aANJ3eeqmONrvj0FjgqKE2afyxrQ20j3zgVk
gFmTleX9uS9Tbwvgx9I5nPc4fjDZNV2zqz2YBjg5NsXN37jWQNmSDVJPvNTZ
xfDyx0gEG9bfnT4go3TzS6MVRWT+62C1hsAc2ovR1f8XaPciNj5lKaI42ysS
9fdK9JlRdHpnth6/0qwcpTKvYUFZXddCynlYkZQmINJ0ywjUgp3nzbMOBuvQ
Ho2HBsawVX2C7mu2vCMSlx6WjPgTTMLJSyy8uT50yeNMkNzg9vMM7ROdqSbd
PG6atCPzKN9jPuEHZjeMhm0NiezhXYyepgLRPJBoU80wrQkKdGGCujOWhY77
AphJL0Km7NSO0vL1q8yW6EgmoF07CgMMcfPnfGI28jUn6Uap6Gc1WgR8CNDI
1MedloAXEG8MS6olJ9Dc7dD8aLjLOoa+2JxB1gjLCYRted0pjU1wtjohAeSO
ukYm1Zcdcv9mBIaNt6ResqosMqnVpGeTtJVIWR/2bgm7kOu3m7Icxz15IOiw
7WPr4RGkUJ2sSTySScZDZO/hv/R8QoDsHoA+iA8Rwaa4i1B3ocLgNJt3sLNw
07PGeU1mcEso6nLgpNjOgdQI8SmtZDA5PdXPonTPsGK09tAekWv4PYNC10XV
/RGyYdU3voHqLYsyQknmxPzB6wdBpCp8oj20RvAz0N484sLb7AWOEF+PPkA9
yx8LmtzTAsUMke2jc9St1l1KuMvdKT/kYOKSAONkz92BhAPdFgv9i9NJnhvn
vIpqMipayPCfGujmnfF2bbgWfYxLlbj8QJLtoZpza0/hoqASv1GwNrGmhdYU
XnjETJa8xgNVqfIc77RprkgThxztKwUziuhA0ddMCH2fSyHw5UJEGLZgVOs4
9DHBdWvuGw5MTg1lfXcTdZ5CTXi11UWQIYaLzABlMeBCZ8dqyyUXwKc9N4/n
kyy9Ll6mURpmV0u5UUjyyZ9GpEB5ncotJ1wjEUH0lRCe2lLHy/QjxX9NuRTL
bYPt31FdstVcUCUyOKjwYXZi5d4Y98EBY3RLVrYiTMLz8yH4ug5x7ocH8TeP
0rvDfvPJ60uuSsp3DRYlxTiiag5ntHKBMq56WvTdgyXdIW6nBm6RhqVNzPO4
HLS6O0iZW204Ljc0pUOJEgzx3CNyoFx258dqXillmtaP9ozCSihW/5yWoC6R
yrGsQNHLzs+RNfVGisj2ypfotWfyO0kxrd9rFZcoDeLsKJz6VyDNy1U8SDMB
HCZZL5YtZxXwuQayG9rfq9MekZYF7J+F0TaShu960qviFWUTHfZGsrNdyuF6
5Amhs/m9TPNjEQlnfAzscxgF1FERKtEQiymamj1/ISZMRuXn3/GL6rBdb4TE
OSteR5dvOqosH6n/uYazxKFgd4rtUwSRDhNaGo4GnlvVgdjR0YEd9IGscpzt
W+F/Ti9mYS5F29pVpG3YDKuPi5tv71EPOYj8sPobHaL/kmgSzgKx1JLEiK1L
/xQiTybTQf/5teHc6ziS48s353hcAnBDtlKYN4Hpc+KSK99IwyQtcZg118hR
BQ2TX8lC4NWQkGOieSIBWmMjY2uBODkPrx4Y2scKzLwFADsE317W99NFNCSw
8ZQVtGNJgY1hbDXJYuAuHXX0Gt1RWoPdmXvVreRF+mkijrtV+jcdjY3wjb72
ZG3jltmRJEsrbBqqXxOdwv4WhyRtf4FCLOPZ4hu5Qvb2QM0yccHHQ9a32IMO
Py2YkgDxio2tQ0nzD3qBfz3KYy8Y8B3bZN6khVrSegByc9tOZ6/nRbOmecRQ
rCfEaqSaSjSx1EtkgD2KJxNhapH5m9s5SQTC8bZ3Rcyy8IkNHQi1UWbtZ8sn
peThAKSRA++YCtanPUdX4nkaQ5SJn17+N3+IDFkMfoJIwUKZxRT2G2RxCNIi
kwAkV5iVf2g90T/jrO0bbOxOiu50F4yS4bjfNV3VBYIAQf5NUY6P9tnpREn9
jWNpFhgsvHABmDJRtc70u01auU5UkLXUEcgNgkVvO8atnaYCCUYLsMsOxn0J
iyhxu7wEYzHnNOUFrBlMA5G/2VZzroCyAfeWIaQJRmRMNDtAtn+5JXGsQNp6
/nWRhq5hxL6lYqku2oBVWaT1FRp2U42FdgYx4q8MBn8Ci9cjWE1JgJUoKEAh
jQJb9w0s1hr/MTNUIohGSZDB0kT9hWFBmY6FjOqsRs+3pQnnY0fJOHD0wp80
pH/1SLn+lWUk+mYDIu4TKzvfLIXmIClUgH+eDUBsA6l6F1E7CiyPDb0tQ8qp
l3WhPPs4D3jQt7lBuu1N/6HbwdKaR+hwhINrAl/eM/bjECLRjWAkmBJgaUIi
c8az7hl42bZpjvE6JvlG22vc8R+FqgnZcXTq9b6UIW0Qbb2svLc/Y+JrwFyl
ocOLF2OvonT3ak2FBDQHbBEvKzQ3QcuNVrlQOMgUONhMifiN9FxBG+3ElrPF
zpqOQzv6IXeAtfHb1jevMS6gKbvahXax6tQ1wYOn23nQ9/5VJ6y+9OAF0gEn
xJ6B36pe7nZURzIR7o0/19d9GVtIJxtrBy62B9prTK6UxfCZmwOxNZV5ip8A
hJhRNT7nSzo0FRjCPceCSrZ2KL9ANj7g1n3uKa3ksZSJbdFUVt3+Nk3tP9qS
XZknkNHqUpKYyHET2hI6B2z0B3Z16gqoTqybnSk+lq95HtLuvaHvr60k+zRo
tintmHJyOBi4GQtPcfDtmDwIqDqPBYML2ej/NOZ0i3aqUz4HalOhWGm/sxmo
grsDnn9e/2eZpj4euydzq5CCLqdMyTs6br0+AZnk8NiVty7FX4dN6FbnrHKj
yZmBcICHfY5Pp3L0qYRO1wAcaOfVILAvJEsUUxmBBJW52jdA8exYQOgGegB9
RKvjOFIQGDN70xQnWZ8b4ua8xNxEzflWBqDSFL0do/l8rhbbPoeo7VG/TQcd
yKpX1mo14FvwsCj5Lgqb6XzehDyVP7P8n5dkZ+4Vd0RbOZ8pHiqGtNhFIjPE
Il3Ls7YieyFiBuF1WPGy1jTsaHh6+VFbLwoZKtBiZZXslqCXf8cjfYWHBUcf
h06nWW2VG1WJEIFFdXcBUmoXKCOsRY0id3j/EmUfKHPenXEhUoU2tKtDVVCd
5pMefBdUyU6ujvk3Aq6MnS5oJwpYhsYlHSzidsjVNHZknP/uikir25Zf9jl2
9snfMR+2YMS/+jf9XXF0cLf6xhnsyUHtJrIqrolcc2PvlpFctDlUuRU7elsO
7AK08A7pYAh/xeBjuq3xyRbm4OK9R08je8eRkwyhOcwBH0r9fDzbHfsbMj0I
FGODCP7wWY+xnVr2mt2+xuj+a0o6/Ju/jDYuExIFZKYwSOgGsxwC+mu/1jRd
pz9e3TkPlJT21efXfo8zwEMj2ICWp7X3dqkzAATJf0S0zxyYQtVnT3DEjO/U
9M1x18KC2L3qcwyg6ytMJvnauqpXBqVNxYcgRLfffVk+WebJQXVSml2cCBK9
FNDEyQhmBODoTqFUEZVjvLhvXhawaTzPM3awA8pO2VzDjE6+Smh2uZ6FIssq
wKjd7HJddIstka5VtGNGjCx4KgW7ZvOkBl8MjXagKQEB7QrpBApcqNFU9V9M
sSOF9KG9wvxoSjozcHDrvfJf5KKLNQacfoBHRqmYINFEx+XfpQWSd5PIzCz4
Rrn4l3sJPhKsWNPWgB3Id5U0jZ2BrXv4llo6t6BM42BxNsnQYON7PRF9yV0h
RXVv0swTnw7mKKwj8tH/gJsiTHGMpZ1JuOjrqw0OjH6rqLIlSyntZZhBCrAX
B0SX8ikJ6j58LYWJBQlDFqYj6AZVkO612G6hYFYJO11area7IkQsDUjpGYWS
w5AygIdwEfHzPpu/Lh8dJaPXP7NLyUscSIh28UIlQcM5R48LZurWWh6pPwA1
dHIASb4NEt1VxDiai87gT0wwleK/w3K5VA4jjhGAVXosOgxUaRsVeSr3hZ5Y
KxrSdZ+cEHaHpqnWzAU7Z0hKC8cdmbkMh7gWkq8UtbpnevmBwhTldcxKupMu
vWSZMvJ21y5FkoC2Xu2uJtH+mP5iuNP9sooPUpwJslQ+gsFeTarA+ivpe8sm
7EuLY8+7sseXdsClx+Fkdqhvwbqsuk5thYrtXMeUqA1zCFBWvyamLIbk8dIE
vx2tMyn1aTWQJBAOo2GCyTE+bhWNy80O+ZM99kVoqU55+5yjDwsjA6px0dI6
rGoVO80EkzAHgbRIiFOKGct5aCM+d8ltbVQrIF/TlhETPjqQRGKqdCaKn2Pk
AoBHUaG8+NfpK2tWgHqn9LzDMw5gh+Xo2XeSBV4+pG+UY1MV1LflPYxi89nN
ZcG1zY85BcvgsKCSFinvPU39EjaUF8JnyGX/N7Ptms/iYcM9s5LRDBG9Vk39
bwsjxbHDHw3ElrtysmE52LKc4VEbuAUt6Fr493ecyc3E9NkqjfKxHAfe2srU
LAQQlNYQL2wQ5mMQ+AChk8pXA2RGbuDyshVNCtNvgtuFLbgB5tige/NsZunY
U6nFvzqJ0GMXfsoRC6qjluh5Wnvx+EzrY4u9o3M617hQyFGZWBXAN11E3TK2
wHT37nmb+8D86eutUI5Mb3LQr2io03Z6OMHVpLd+lCgf8A5yla4fFMpEMckf
9Dl5fknpkyrijzUjk59EZ0HKr8sWRvwVsFVDeHbs0mH5FfmjHa4OZXr9TdKB
yzZwzIAZbijVMYLDFLcEwRtgbIcoQIkd66X5gOAtG6BPLxAtqBNYZKLRU7CL
RBQO+ZHV7fr9VaxbCQDoQnFVErkBii1AeeVIubZyLLsqHiwgeOg20+cPQTjC
k7G0GHSgLh4ZjAHoHeyqjeZ1L1bQy+TUJAN32pjZ2SycrQ2BEz7o0HJaQF2E
ciXvVrt8KuhSqNxbMZ9mUvQpWG56mnO6F/yDqk3Wr8ZmOy1S8MI0jMtcm175
dN+6QTMmG7DAW2sv0IzmCraLa0wiS55Su1iaf1lUXgLG/fFQkvMTVkqZ98+a
Ei2PmZkanC5F+LxZTFELNstOv+UhU2ld5HXzSI1Czro3a34CEiEznK9UrV+F
tkWU5/KMukjp8tfzODsZAfDxbx3KKPvYJb+tgsQgUHnpwPfMKLXlxhU4WbjB
GVt4yuaTW3Ei/OJZbGTw2RQrrT7uhzJr8SUGlvVs8OwuSw7u16vfzFpcccYv
whkTS819PAUeGrvP0oFYFMul7tHL7k70yy++02GpkHmh05a0rpVX9dxYHe4N
KK8g+zuWtu0lwkNxwTZPpswWsrR5CDfol9xsWlqzFMfKxS6yBKENgyF+NnQm
uQzPsBSZ50VBofITHZPI+cfONJ5+aUXQtiz37/gy5F4To02BkS5wKFM7Y4vZ
1R+V3aErjVBcnMJ5Wtt48l1+EuYWHPIJ9xgT12hHgGT/KThi/ZSemqwf1hpW
7Qj8/W93jDqJjwTT7LpOV7HNhM9RnbUCU5z/Xtb9hoGWL7y25olh49BF5vuT
qvH36yr2PIYoARzsbxOECOws7SxA/71ttSaag68SUxhPspcskPAmZJbqTm4f
abn3dVce128mRIWnz19IaCAkGOlREilkh56AisJEN2YNoqK909MaIvxUr1xt
w5qXobRd4G5zFX+o00sBY0811MLJ5ENu9qDJqM1SprLi0TqaSqhgso7GsS39
NkLxN4UMc/QpcdbFYcBYJxewQ+LAN+h+1yu1oAisn7K661vkN29kzrQ4sjM2
NiuNjtJ8D9zSrpJ4g0hprysUxgXF9CDmvzqrYIkTSWhJD1NHG0Gw0566G4Oo
jGjaX5ja2m15aCe8t3/EjSy0V33s/nbcBy14NDkM+pXhGbwNRLREIiLkWKf0
PNpQczKlI6OF9fAzYs+cJOFpfMrDDsfKAOW7MVeUHYvnTv1HNd6mdOuqZkny
jseFRseyaWVVlz0LykdF4ZZs96/kR5ZvyMHtRfmBcgX8FBS35lbMGWQBB9Lr
8CFH+0cvJfR4R7oeYjh7TuFdqcYUnHes4bgsbzVrt0vPC8EwFSufIpwHjzMC
BJ2fdYwjXnCilN/MOBHGOJbc/RcxeaJlEs5J/fOI1ii7tISQEVCgKX5b4DoC
rGOSrRP6VzuJB8MmSJ01DhF/wbtZUNMTcHFpKw0uT/pFJusrU9BQ7EDJ074V
f2dyz7O623mmCSoBbicXfPbrJL4jaHKdiSC2u7gzk8BLPF9kIjfu+tvpX2F9
7z4GiMdAKawnm++nsrPt+8nkmky5zApy9wQnFtlTcoaqd0tAdibHjPjlr7C5
dHpI3xV2U1yqP0QbwBYNLFAuuXjwdQWuZrqtNbjSRx8OQLHxCTmWbnAbLZdJ
sdkzQ+ZgcKimfrQ+nA0JFAH8/JK01gr9XQRKclu4JA3FJqoQcBYLpC05PjUM
R7w0EiRNTMb9iZHdgXKFz7/Mby8hvE62NOKtSDJeQ3yDXqK6OlvMUSvomQsj
PQiCQOJndzok7vyEjVC/th5CIqllukk7TbZuu9LIpf7qbqWzx231LO0G+RrD
C3Qyh74XDOUgNDZEzxot1BB4ua6mwtie0yzob10sxm3dLMee+Aui6zFBUgtF
G/SV+2V7A0zo1g4YKW/Bv0VBq//hziHZzzlooStQzSbtouIjqUer+qGjw17P
qMfzUHHNuLUEh6BLkBIf0tcZCinFAI1OO404DNTzBZPa4mq7Sg6Xhuh5AnB+
zKRnwM2x1v7qHzEg6h2ckLXV1uU5c83302qXKyCmDa3oZQE6OMshtSjVvBPN
Dh1DkWm3167tqECWdmNWtEvmomZ5XcrR/hoasNPgZI+RhdxCZIoaDH+/yzAs
5+5WA5hXhdr6UZOnoHVCu8G87k9in/C8LoQphq1HI1EGaSBw10GQVZBXApIk
kAlkbtO3EPo4iVM7Cv9PTVafJGuDSWW9cVm3TPgETTzyIgsB1hTCXG3E/G5E
vsANDm/AqnbMuWPk+GSQ5Qc7OS1H7m3Ijzo2eF1U5pyYhKxA0bt7HiURnbjr
tvAds0LyfztOHVL8vxzC+gNvYZvRxOm5EOh2vQwgoVxvqh47qeuttezNDAzv
bcZwj27Ym8Ok1/iZ7fydw7khrDtNVVig/HZMWRaMHWkmAZniFpuBDWRwRZZl
MUZs80/yx6TTHtQeX4/m63UwvJvDV+cGbMsTJWsXCZ0vSXZSx3CtQKsvQU8N
GLz+3m+SJ+cZ+u9T8+1NwQ8vHZZANN18yI83uJP38G8j8sBHMGybJX2iG0pQ
x1uMq2Ei4Odkf2s87ubk5ec4gzqpAqqzMWmj7dHvH8l+XB2BNVGDyYVfnG/w
s+hX0e/DlEM7DbOSpt9H6w9lmlu9d38wWi+8MOux18+055hkHIz3R4gQ30RX
ZUzor+OpDolu0FCjh4CcWsoJkTYiDs1Dx9RhuSfKQZ/ELqOEx2gVQEpnaY9S
c9IoO8dgOy4wyEJbow1Yl0lcfiQ/7Q2x6iCQwYKuXd6lvHL07doKcAeGgcHS
gCmVq7OvYYWorJhzdb1MUmgqdt15UeFXvnU4tbd7tMFHtuUPNO1mszV4R0sK
QKyygEovkSrsx1l37PhqlOBPCW4RTIhzYJYAlUd9mGdCOzli1mpT0SybGRjl
qBiLGKhmp57nfrvg2wFrt8GRZJc4mx+LcagwErdfGx6jKTveCmy6zmWhoW0+
vksqa1iN+z57PiMCmlgTxKTJAJ52vk3Cx3KjLkrBmeirlFyUY6Q2rXMfCJWR
0cZKZd1uHN63tThBc7FVzn1FTPBHNbMGzNDkErZlcr1IVd/dixBcpv3hUC7b
cmnuKrpvRUzoidvl8aGzvsEqnt+d5D8mVdq9msuDlrZSV6JtFiwvYW9ivLkH
IkP7m3hHqA36ynk4Qfy6yXrdUBa95smoTdRgERR1tdfArhtNKJL9x4U8g++I
TpN020A6qbpSpZj0rFtKlbBpDlAVZW91jsiTeQ5fDEXO0e1j9GhgBCzAqEM9
JAWN4MtuxvF98ZY97ZviWnLXVtj7eBmsl/fcZYbvZy3oBhD2KeuIRP+G0et6
Z+hahTW8+pFhPn+sGh8Ue2afCGiTMaBwtjsCdD3vAAfahyKOak+uANTkVgNx
KS5+FPZXRaD1jxdNN91RCrMHW0ygcifCLWq43eN/pXtb3vQM6KhOJKVZ77ZC
tQqTrEBvKzgWcDDRcSlOwhD44Ypo16IiOrARkv1sXu3ZQHMNytEGjVS81bW+
uNo8+nW8C7iSahf+QPYxbmI5e397s0om5Aktr56pY/4RCEzKkRBESTwan+jj
aPCTaaBenAfviKRV+DP1S/dEbcYoab9nuRgv0ch+5FRa1lA1WAv02oenhvmY
h86LJM7BdUWufNku6ZNQVdVTdwMXk6zGckydAI2HyDMRXZ8jbK9lQtaOBhOf
SzgVdS3Bv01HmVl0P3iWBzoIGKdEpXCOeSccrP+xTQRnFBCgA9B067cPsY51
gIcHHwmSdKqgp8nz+yxviiOV41d9CovrrPVKXaX28AfzZdm9FElZsxPiK0d1
mNb8cp2WFzVxsRcdFnx+Vph5MuKfhHWcajBy7h7RQXFrM7gJ52IN3DdaIYgm
rQ6WRLYXftj2Crbsj/CIwxGKRWjmNR1DSovdzON3z1h3QzGtK7hoxgr1IcgC
U23Cb5AF/rX8ydQW0CtsTTZWWLCZRq29AYt3rgTH90AIVdIwyBfBf0QRrPDf
JaV4Vet9+bAAF7zxIPZ3TZMOc6mXgEoa+7PoWnp7W0GQ9U0qA3pfM6QKe5vQ
I66HPs5gOil9RYI6GIy0trnwXxSlo4qAFiKVSsoIpJurZ6iGRN4DyHYs1Fgv
9FIkPohr55d9wn+WnFt8/1uAnjpkWgMyTv9Cn6Vme6Z03y3boj7UMdsl9Ecv
8dx+Jv6EALey5DuseHM2gauRWcWJF32GZR485U7cMmTnMDsqnUOhGJmlpYd0
lpFNVDCbLetljl1gjV36dvWofCK9Q1hcNehPxV4iPjUHW4zN+eF5/vJIc4wD
D9RYCYoH7tFIzP0ekP9PKLYhOIqPs1GVY2LMkg8UrA+l9UZRcjTZvsC0/N7g
NKb0R0DMlF6l7v+WdizhAyVrRzOaSB+Qp3rWlkzTKvo506GkbiAb/jxmojQY
eXzxMzEKcaVw0P3j6evwSLPl4tqyMW/YoMbS3zQ0LlJTF8+FTF6swTCKjPqC
FGC2d2p2PBj6pJpRpo0asvHi5HrEv/EMgi6PUceH30B3ueNMtXab7fWNdq/r
TnXHABL9IBiu3YWgJQR7qMxSpRrLe3mJ1glcqXoZPqU6iik5EAO6tAeUol1F
njs8U378jTpsLxCyXQYICuaousy6SK2FM8QaTfR+n1m3xdDON3YxYwb7z5My
yyCwrVZw1+NL34kIuigaIeut+zd9M0WRUze1nBxDzRDrVJNVwMsCoLkLu0qy
bYwwUvHptOuDoBUCyPxWCZV/bKL6ADRKgvAgtYPmDdVm6pFITYVT1D2zwsri
ryb/4MhxBHrrUJHic8Okg0EWO+s1BbmdKaIoUwDWLULDCbI7J5fh3yuzPogF
pgsP34aEetIku43Ug8yxhpyISvs6hmXXsAO6UxZC8iRfQK3erGmUm6atyHdT
IaNGsBmfxulEa9pRVNPaVTCYbjGVlg+nXl8z6I28btefwDBhuGWZFo4Iy/Co
IBDhPaQaHh9qx99oFAh0UOlnv9aJRXh1R5iZiQIZp6wg+3jb7K3bfXGFVYTZ
Ama2Qo20jfFri+Pnrs3xZd+6YDdtnpHeE0XTbHZE56c/ENF3DLiwLlprPI3A
juBVsKhVBa6otGkYp3lgsUX20YjKfC9EA6dHkKg0t6fNF35WLpIVj9lIVJg3
4tqIiPIRmYMOYJ2xTUyfoqTrYbD7SEJfGENW7neV7xM9cXcuLKfggwjhxlpi
uJhQXCB/XLw9kkigSxL1+b/KD+9elNJeHxDoXDyhd0SGzUzYGBBxY2R2zLqo
JmWVW6NLktiD13liodDhTuKK1ozf31x/dNtV1ljiom8IyIlnxhwMJfpBuLVD
5Q8yW1iHpZlpl+81HffFkOM2LoFwCpNKQnN/QuQHOR2EoVLIWDXgYF61YWSs
Sl+4eYjrzNhZY32g6tACODnBfpzm+L4e0ZO/DH5+UBNFr0tYwcZGXUfb+8qn
f1k2Vc59MwCPCFo1QpPDeSiOamzZF/wXdJ/jb7iCGFOQUydZONFTmy2wSxWb
hNYrbUDVCgvZntAHOLTGHPoca/a/y585k5HoGlo4mAn+AnH8sWBf87dWIqlX
TvYXCQ18+BpK0MFJ70+gT7drPeE2+V925s6JlC8U4FE51zDzQ8bQxKsSTAhg
Bkryc7C6C3QISrZGWH3Mx22gUekEdSPfz5IvAaEekMG8IpoXukqsk0KJFMkX
wAfxoc/zVmtTYw4o61fcKx+9cow4pIeF5cfvTBixOFfGKHtvfvtNn7x7sFCS
yRcEWKxSdYrGV8V9608ykqBnv6R40rIeEWGQIFhu0A2Rg/ik5cmUDNONwaxi
2i4niZ1wS3371RVVlcQjRXIK+IvQhEEmfkR0ruhWP0BiPdXqwPvxxklCS2Mp
gtmll1nPkLy558un2l6zZpQNn6zEz3tR0KltYFo4BRdRfCPkqOlA1R63vy1G
HQ4J4SGnfbIWMrDYVdPE6gHDZgxtDmnDOskF9UCNRGQRE95tGb9r1hTAtDMT
yT4nxMPPWchJJpRvhqY8WyI+6pPNAEJnRGh0+pjRlYqv0pxuGYQmqitiScGn
hDfWuau3cHT6HLSmvrJfseGzV5tR0qvAx/rcGfX0kDNBucjAVUqnzHJJSsID
ib7GwTENUAz5LRya8sj3QaluAI6A80zIhc7sKWn9OIV4kYyQH94niw0qJq1W
wXYTQtw8iVMk0+CrhVTvax0h8j9yfxhNPoQaFyT6JtvR1um0oAdjCpSHR9up
wYpCAcEKIQBUmN9YUoyAhUNb/OPspANGOwGg9cLHVgIIVXiH6Bq50zF3Drsi
Z62lAPC4Ng3qnFAeUZSks9ll7Artgu6R96qrgft321b6jJHUynLjt/N94DEt
S7iD26kSZeD4m9hqg7OU3HasLmb3HFcpqNxVTuv8eaHo3u7M5JsnFraJoalt
cLephwvdVH6IJsMrb8aCUi7jIB6kVYSfg58yKHsBQtJOpu/9f+/uR7xrGQwx
H2eNDPJIzH9xp9U4z1Hl9E9/hfaJ3DQNb89k6s2rqzGoVarItE4rv99yX23o
v5LjIFv5pIncFujZYfm2jmhlpr6AivpY9YGaAxKSqzjWtPvMdaWMH3ByNJDG
dKVppZSwiv7HzLihKdzqPNh61TL0hed/u8AOgnjlJBgmMu3F8YfeSIapj+PV
3qNBTLv2DTtwkQu0t6thOArCAZJ4wTBdBKAxC7LBugSDUi0fWTVFF77JMLW9
Xwz9+/LDxla98zcvoNlQusy2CF3gQUJZ/HxweH3djcwzCo0bJxOaFNULgp3T
UwSMeoMq8wF/dHO3srkQ7gFPMdY3/uUotOLuH87YrfsmXs9Bjhnt5ucJAE0Y
iKXBmXRDAyocpk4ZXewpw8wPdL7wNiS+Ci87u/s2dtzibbFJrAS4xFlL9HNT
tYO3od1L27F3hKdtX0DP46QVrqV/0xi8vQoe7ZK61MXf3ipmeHJ9xXxAed+K
1kQ4EaUcV4iTRJtZVJco7Lv4bt3YlCllBWhB5yXSeZOr67NxQE5X759GPad3
a4Kn36IrRypL5yRUOQE1uzGL8Em8s4AZR/srfNqTwDJsRbc2Xiby38dFNNMk
H5+PYk8zEBBxpgcdRrqHfWfZTSfLVx5EcI92dOr4Xme4BB76Mdl9bFo+/hKE
YYk8vnvpRTcVbWWgKjDXEThW+iJg5pI6O8Alebz1lgtxRGYTJbju+D3COEI5
/FnpAtaEPxYPBMPYZj8LKzq494qH86RqS00ftt2okIhfaDW3giBYGJiwe4EG
JE3ptavpdWQ6C++hTG6dlDOEYHynVujk/i7qVEw0CyNglLOfGcHKItkSn8zq
cdY6VOc/FeU60JL2oYp3Wj9BS5WY7/2Ag94aJS7/u57Ifm30hbTXvKedQfwv
D/Qr2YYC307XG0MFrk5lZ7csGRFwJZpLxLhv6iAudaZPo56FxwgvwxWt8h9u
R64m3/iWXxguglwSI74lO3KF/eF554aqslmtvw96XstFAu2MlCWi6WSCd5AF
INHhIp8oIVbiwwQbGbEunyjQVUlCuRiXomb4WqKeXwSlhKyabA30fxnFs2BA
fOqXUMUdB+jkIv8tn8v70cnCqnobrwO8mYGlN5IDvePqODstzfTup/Mt82HC
zAM1rm4bfpyLGRA2Yi27KGTxlB9s5Hd+owgx/JATWfvkXxmLyFzf5k2MY3tH
RdE+3Lcrr0I+vRTf4YGd/vEP208CCsGK8t5TKO3t+K9wtfDHlfCW04p6mTno
eCqCg7FFkBDnrBuuYsNdJNTNqkGWjTVB5nAuHI8/hibHPWloNkUUcLQXjZ2l
3yq04UDC/sqkyFaFQwNPwvLlr7+VLOOxP9PuHGgKPUJqRlMyqjDCofhfMesp
ZunPFiPC/4XNXFscWeLVxtkF9Zh9Hjz7tIaTUpaw8kgVwBdCw6pIahZSG8Dl
Z3fzTH9dyAV+J2qheNGbNDPBvifK0j84FTm+4m07dGWRL+VN/db87y5habLY
oS5t9NMPRfUimBFCdMtv8Kg8Tz54yvf4dSCHt3oL9cM4BCMaaHOibCsWJww3
RXWPhQexkCyRK9+5ANv0cJnJJ897Zv1ML2UYlvd6KwixJV2CzBOoKoJRMGTD
b+ZXigRdwCzHdG/MmhzXiL9zn6AnbeUMcKzrjhgf3vlLvcG77mJnM2/bSeKU
gwIAJAyMydsk8cMDhkMSoXk12QHNAdhRqQScl+n6n4Qq0yZazxoQnDkvg2/k
p0AYmmn+KkdSa+fBsNbCO8w0awA+dUhi9Q9eShgSKJBIGVK9nkZZXbOwK1Lk
lROcDjf4nfjD7Nqksem1h4ZzHcWe0EDpyGRAKi2iAdU5tL/cNuw3u/RPrhm0
o/BzPcU75SASTxWFd1IRBb3yiVA+jRr2onrinwQFgVvywD6OmyOS+fmnLoBp
xIG459I6Igc8CF9C4vOjDbHK7v8IymlfgTnXosGMyaJnwO5ezg7Qk67HZkIg
bWc6wPmOjdEpjKOxtNIHidncxTeZv19vHD3i46xFwpkxkC+olJ08758WYPFp
G6iKvoZrPVoVNPAm3jrWRkZfSxX9jpYyKleJDEa4hl4j2T21pJeQX2QweKTr
vVk6VHv3f/IUo/nF7FG4F+Ni1z8afAsOHv94nUFwBlMHbnrw9eKXS6JR+gjW
VArrK583rMS9ttN0ocY1xV6i2bXLU9qXWJu7Ivjn97ymNGQXW6y3kaEqvzSi
LSNo19eEufD+eK79/TEObJJuG6hosEq4TwKBpXRM1A8zpyee5WXbTINNlXct
i1C4/Y+rRc/lvMcXwxzvk+esVd70N4ySa2aQn9iEOQDvRHMqwoyzVHyCJp74
HDGlX6OW6KiIk3A/gFzKdU83E/BjdSrycB4+M/xAjPgO4Z55ssGDszdWZSeC
FatLCNubruBs8vVoBg0JQ6FpW3xOVmd+ewtEVH+qLjmkXbXSsbEIQXnd1xN9
mbSHjmFM771Goodir46EbWL5QL+EpLyWANcD5xxM8xIKpdqMu+lCk3Lp0vPU
A/QegyacLrxPuSxDyNuBye824uf7tQsd0sOTj4GE4azdsS+TMdmvAhXyc7RP
IHSyPh9Fx6wgCQQjtLBJhXETimra7nY3a4d2F/ZZYXpqNFk6OOYmQfU6/uQz
TvqMZsN66xrBCVZoy25ux5kwWRFQFqnHOY6VJrNlgbbpSGYqIL8L2eXlQUbx
Bo/cn7kBsn5VY57kxITc55/vHnbEeOxsqioYKyt0fDL/yZa1sfcOT/0vlDti
RiDq+ParzzyeIqL30LChgT5XfMapidU66yg3BeC4CS2EaqU5BDWyrWixEhQ6
t1A/HFF4BhG5rUuKF2HLlMmhE83GU2+5OH63v9eSKTeoA38m3grQnf4wI6oc
KnUlJH4tz9YTygiDChxNUlVGGpEMMG6ZTOgloO9NvEZDgDaZkZG1eIXj1lsE
l1IjRxlX+xrpddnoK7j851ErRgStNUyGZRX53XiOgAezhDGJ4NHHxvQ7xx0R
OQiV1XlGBYfbv2gBo4CaFLYrZ0MX/n3AhZ0jtQYOylEH8VK6ABReFCzhL1Sl
hEYyEfzy6C9ZSQzCHsJ1Y2MmGe2VCJSFest27qm1uW03RfEelLxcCHw8YnrN
y333gcI3NClzhXg9XWUPt0nVLFEcJkh2QC6pnQXjeW3cVu6/h0QO5d1qFPEk
L3opEqWXPF7sYr7DhqqcaycjS78phcVhyfWouuSIIYJN3FrZYzXdvJSsTIJM
DFdO4n3LHrtNw3+OPWTm5ZHOjruv/+llWub91VUX/vCojn88H/ipXe7DsXl+
uMMJrOHt2Kp3900V0cybh2t6aJGYiYx2kPdf6kj+bY91upA7q+O/4BviLpfB
Mo3HpwnqkAigKXiTrGcyQGmHD9cIkzmiaHTjqE7Q98dJi7ynBKHXhY7Xyzdx
l+UKa1W4/n+I+2bYT4WYUm1Ook2Zgzj9NtvfMs5F64qIuEj0edbj+Xv5WiOC
aPg9J9arNgL4jb9VndMfHi771EKfJCgWdWTnluv9wIE2MZtmKOsWvtXhZ0iJ
JYu7pmYAu6L6/Ad3m7M+T6kNHwsQtuCskFZgMGu7/k/Jv2BC6a1rFuXhLDQP
SEFHxgWyT8kahCQ57ZxNzp9JbicbMu/laAhhEG13p0wBkqsL3xujzfOOkLU0
Ge2aRoqwB8L5ph94gAZSsBcloHhUCwhE4/NpY9R7jMFKNvUMixWDsUhtDE9U
v41C9StsrbRrKWLk/Ygm/2TjzsXL92tNV29hQCugsaxNydq0AsJjuIPIgFPZ
bJRnr0W58Zg1UnMr5cpzUQXMFAkN5VIAJi7VOqgYrLwsoCIHqMmuCo/tFU15
UOv/KIAd7fFmVEbzqFLCBxY0wojO6qyk9gw4dzU1ISzP8SKvSBr8QkkU/01H
dWteWsVCj/nutei/Fh14f4QLNLADNb3CUZDuLGAQyrLqeBcmWNvcjglpGgVk
HH8UdWacfpmSJL4/SUg2u6QEysPq3faKI0AcW80zIJNYbaQ1BG2rm/1x4tvj
ygL1J3nb+HB529Rz9Dv1S6oOCQUyfFYearVfFwIUT4Fjyy8uF8K2rN2vrA2s
OIK1iu8tqlq9lmlGPHvdhVhdsxfbb8PqyV3kL+iTHFwaTZtdTPljV+3R5fir
8XS5z92EBD4b79U7Djh/7/nI11UlPl9PVofKEIeQmxTgowcWJgST7tm3/LnR
bA14Pz4gqKJAzCrnirnkRCVohNzkZIhdtp3WQ9P7GMjGHk5e5jNQcNOhGIcc
Z67Iw0w4nFbXYnzppB2/X7lPOXnHIxJemYhsZGaEwa6WFo+xq0heUFf2zwbq
tvl6umPCpaBMmbHcXAcQ/SOgEyk3yBdQNrjGRG/wop+HnxSxiThX1wRznrqm
uaPZuOFtRLADKqLU9Ux0d93RPrdHuFnXUBbrRYoZU2wWHgxHiVkfXrzDZm+1
b/gdnZ5YG+j9UrMBapLsRwaRSmY+prlZ8gy2JzahNL0Wt4Fg0/xL3B5ocdQi
HxzNH8TecbhYW8wcmo2yR+Nf9I44PkfjxBX0Y8s67Zp6H2A7mtg8EgPL2Nkj
ANfpaLs27XOc9BfcNtneRz/pfkdwa/O2QPCn/RRnReUlcgHbVhGd40Vd3Csp
FN+W2yg54DMfl+nGG7cSEx2dOnbTO/aENjOgX1njp5tpG1KGMl9ru7hdscHn
CIf1YMZA1p5WKWyWjR/fOFMz7exrA703ZB21AnGVkNsuGtusxnCmGW+I4EU0
jBNsjzvJdY63dY83tIYDBWzYoC3hx3S6k0/IrbCwdcr9QIK2HTbvAPqgBuwl
usA6oHHe5IfJqxyq2rRQZDYzlvqkPd7RKnjStob0t21RoO/XzF4zooy+6CGh
c2PnJOThvsPnma9Ljug236PiWzcZpZC1R2+c5ERSaAixj4mOAAo3JJJIPR7a
Wjc9NnHOQ1taDHbzaWDo+xnG6IBM4+3BeeHjba8g/vj/6NrEltbAb08DcSbL
b423Omnb1PyC2X6YD15B/WYhoUjo0G1n5ZHN95QKls3jgR5UkPT/FS7dLf5j
RsJAQRfHIPmM20eC+6QEarLXu5pHdui4VLjMZKyrbrN6qTc1r6p5R6Yokn6g
Q5TfFLzex1fU/iDM/b2wI9kTiDF74itQCCIFcuabdi8tAXyJmtCztkjw9R1H
A9zD9pfMNA6Ex5qyKMExHpKPTXWoYp+K8uziNm3NXcDJdWBakignONORLwXe
xSYuUp2923n6B8ukzgiF+RobZzMItnfmJJHVCsBAQgcLxxfMJddksmIcFlJZ
SN3VfIQfOPX45ocsvrA4yH3MhQ4G2KBD3ftXX82hXQ1h8U4IZHAXaCBNxcDW
NUhWSN86BVHplJOuE9yilgyhnqmFbT7mPzY03248hh72e2oEZzqTaG4SjtjO
zh2DJZr5OFGjeEePmwwTKCw/eIGYBCtTFiUHMXnDqIsKm4p4vVhJfgL0U9iM
UIx7Gyazur3aodjOeCK1fzXb6OyZBpk0Qoudlrh5EdJpfusS0857u5NLzuQg
iZnH+B4KfVtMI6+OjetkVqX6dWmiPNGyN2VYLzeY+3UZaHYQzzJVK1YuZ98T
36ggaApks/ch8Ujq9IG4WNZGaLyYXFfyd7lffXmWRta3sX48iJhqBPxP6RNo
3IbBHapiQBLEqO4cJ3MnY0j0CzVJd0IiDS83kFa4pCAR3Lzyla16WPbDJg4T
JiHa1wwLKTNSkqR4HfqijJRBMgUus4tWUkxiNHgulZE/QjcO0iPLbhrL74S2
VCRATuBg9VLMdL0QMB7SCgpd6h1finxm4OIjD/vA+ikhQ3Fn0lj8rZB4/6uB
RDcCpaG7ARkwCcqqkc+s23q1Gmb69ugQcsDmjMRS32x4BzMJCsaccZK+I0i2
lBorkxgbLJ8+AGq1B7yOC78sAxc9AZpFKHP7XkGoBYdT3821jQHtgpF31SSf
KCYvuBgc1v0BNp4T7hamdA2xt/W5reCW8+nF3nGFB46RMuHyiC2p0M5LBAki
Q+eFXT38eZv/iUKO8ew6gmjBPg0/5KVq01QmLR/mj1+/YuFvPQH4ol6lgxS0
yxmfDRahZjtYFCoAQ1f56IxWJ3Vkvc0XV2RByGnS3IPGQ3yObMGaN/kUWMIL
86R0s9seHM5a88GTeRxsPiOuH6F6HC8nwPM8zGTc5RprK3U7bxAEvcjLYYvF
6xqEeBA5d/H+GNiuwtYabovI09SnDtAHiow+kmFm7QaxTOIDmteJjI3saFZJ
SKzhZvXsn8QOiDYWZHXnN0ayr6v6r+59NQCsSCSPdEumoS+8fnx4kJRDF7XN
6BMKiTa0GoDTxn64YHhq1OAWhm4EZqvT44Hgz4a19ZYDglVvR2J/Vwj+s8uZ
DOoO9qkkFEK6HDaG9A51NOs+gki+nJjYX3swl6Sl8R07RL3uwnXbzHP75Ggk
EUbC4Eo0Rd6am09CbtRRq6xpTCqEJqk1qPTnV51KJ/fFWko4+eJkG0XQ746J
3r/wURKi2golIDwqzvivznOblnvKJMbF+gV1v6m1id0uXGRXTBd3Bl4dJ62U
aYku1OohYVyiuKENHUqVITEFQUDQISKkPsj84bIvW2OqT2aaH3gf8T91yxEF
ZtAbmdcWfg4bBMw/PoVqnjkB16D7M31vZ7M3VEisOr0Hho7b0Cf50WrtPiMj
op998TMqDUl7bOwDFK0V7YseUZ1WA5C5lMo2Jksvy28QmYx8Y6Hzjm3VqNdH
8DW4hsUFiPocnrGpGYMHotMsCfsnsaDTcadkN8Hi/GgHOIAxMOnAUxNhc5Tr
Vz82N6A7UQaQ/bYxbCnkB28vDXuzJJAnU8xM74VNt0zvt1jWf4fOpbwQoovD
6xq1n8uRaMHmSLuuiFjeABh7rEQmd7iepTQqfSAydhdmQGzDKapiWaGxcukx
H5DnuAV86vH8hwS300Xz9hRO8mcig6Z5B8LXXt1XTJiNobHvA36q1mNep0Cd
EggOQ0HTXRCNtcbBaLLrupHQfkgBTwFGsuTG1K3IxGiRlsE7tUtVZbeyAJvB
GEBJTHDGKJoF3yOIoMXdx6YTg1m5hXpRGoYIy4WReEqP3t2TNyosP/ECi3iv
4ZWquVd+gn/L3EIaSFaEwHmNe3BKQOTLBjdZkhYkWMra0zYvHVAkHrzdRAeV
ClUCXgVIOvSPlxLCOYWIFBF2byKUb3P+R/PjKA+x97Rr6nFhBSceDETagCF4
Xlw7afmP9rq3mbnA3zNZ591InYv/F/gFBAV86Lpd0ZasA9iHTtgoRtNVC4Q2
M3DB4flNZ8Q9ttIMYGVuKIENGxdTmDS23vT5Q+zz0n77asNO5QSHs007yzHk
KKCZSNYYG6IN8WbxLtuJqw4chgK1+nUnViVXyl3YSicxxvQSsMdInvYxnXH7
vHP2HcI51TL7t8afqQFTT9ckkwHrXQFmWYJIWrfH5c8tYsfCZ/k/AoKLbIZx
WFSm8tumk04qEmCoKQ3vjhCc28ISEgu7fUrLF93pfGQvHJ93Ll6MyRHA2NnA
9asATpnJPfCPnnCfbodKsd3V8T1hVb9xg8V58AaPxZ60N/cPU4sd2AJdURqD
FOFMifPq8CkyMO2U/l6v7Q35Uw4NgxMp9FyPwgva13Ye++uMPxDccyIfDj9f
ibZ4XWMwym5ZfF31IsYa1vl54Z2BHR6Aif24sU1nPb3bJeCBLH5VNQSV+KR6
R8NqN7AYZKTIGdeH2+K/g1uRy0eeylbkRYxa4uS7n+zTU5+p/gLAmNLJxBtO
V6g+kxiTs459Nz6XHx7mi84CCpRIoAwBQSwMh+zTuJuEPWnMPoqoLRGIt/AD
T7fP820e3oPdi0ckq2BRSqUqo242f7uXbiA5oHSGYe3kELk7m446Kpr/11pS
NnHSRleKe17HwreboMPcIEpwONNBc1g/DvnIK4BsKGjUfpxiuzgg8ydpHClD
P+yUKJ1UJcNuAIZhaIG+dZrug0ZIB6LJWmQfVhboPfd+LJHdVffoe9Yz3YGg
ZmoXG2giUnh0JSooPFAq4Ut5ZcWg0CPNkgqoyyx8R6po1v3cwrTODboLZ12U
GgHDgHhZUisr6a2r5gW1jIjY5oFX2GAlIWhKc15LN5Mv2FWwLAi4gmFDAkWg
FbX5J3zwQG3CK7VbgpEyP++bCuVwBrmqrABq9FjRps5ekcZ9lkLdH/tSiYwa
3kbE23P+CkDtpb4Onkx/tBurfcWB6FKRsLG4lO3wL42fom36mVNflN+W/b/X
aStCw+hrA3jA6uMdj3K2D27LJg9NHiFcrXLY5W/A4s3gFOxhdtoOGlClripd
fjk5qHtBGMR1o6LWGFUJLgvdsWOv6apYNPOyZZsE5Nu1HdQDkp1yI/mA6OsX
uGBRBfAHzAb6aYnTAZABckoMnbn/QxvGf+Q7GPWCfyGDbVGcKZsDyLzoSQ7D
3nHpL/ApLZZ+OJ+tc+tOUQpWnTI1yIjDkVmghJYPWUQzL7ECdqrpvLhcOXyJ
c5qwZw4JzjTeGL5rIIYGLbpLtaWqa9I0Jn4r9Qi7wbRmXgX5wDfC/BrjG3BR
uhTOv7eCMeF1pknOoymPpMAh09H8KJSNghbimIa1/jmtTaVM67o+K2kLCANZ
6aTu/TdCQHwmFgFWWx/6WyYAqPriEJQgwxqy+Yom2ZfatRZkmLEoGmZLEZgh
Ms3+8G1CznyYmeGcGlYTOuP1PD2Kx/pLy8J9MMBlyudfcBPXL/Zo7czVsrzL
3eIaIXHzQpBELR0u3gcCZL3pBOjMn0a7w9o0iHhRVjs/ABstNJwzOXik1QSq
0mxtUdzK+hOr++b2aZZDvWArYJr+X+4tpCwkBbaRBQvFdoJk37+7nHYmxt9P
7UJqVm9xfnWX2HmJBOQMX9jW3sXkQt6DCLjI6iB5VDTv4NxZBRg0yQLj8vhT
esZECfs0qsVJBpDJ043VI49AJLYaD4mjF6qhZnhVDTJ6J5T8BOHx3ehUmj8V
QUL6xAwwG9JTlYwpb5MXr16bDgyVRBBBCktHZTbUjEkORTWFT5XqlUiQTVv0
Saum3d9IUYZ+qpuqiN0T/gJyXrwcDKm/UQNoW8inYM+CSOyJztAJNFmYA5vV
W63amurM1+z/NK8+iXGIE5JgNt8otsww/Q9rQBKGQj45ACG4HXqCe4SDgz37
tbRuilsAc6l7toZrYiO87ndtZdx4HD9UROW6X9zDJQgK3+bXEP/XVbxdpxJP
cyUjNbU81aGDbG++uGVEhMx0ZTpPfx+0+Vg0hqOC/G0IlMpb+ZnmjL4a5UMc
O+2SYGoJeG+bd8tuBY91YDdTUWUrLNcqEcuJe/a//oXF93NHR1SXq+QDglQy
skKClwyDuDBhxuObaEnKAhUvpKINIInK3RGzKyrhqYHw/kL8eA20gJaJ9bkX
POHvYALHY20S+kXm7aQ++6HLwdlM9rWkYiqaB8tJb7f4ilBN05olfxotxS5w
xOmZZKTLlwg62IbpMiDGlLhGzuebdlg5LR4eClcu/52g/MRrYqD+be//nBZx
V1NS1m0hU65RnUbI9K4fdHAJK4TvIgoBsX0wZNaytFpxlZG96BRZoj3btZWm
7vCkD90LAG48rcd3dSjcB7Gvl3khRuX41Nvu4HnJ/AlRf+gkqNBcki1lKm4q
Fgrq7mhDSRLCtw2QLmZwNinOdLDQUt3/ym8cYyZKCkMPFtQsxfxV+h/Don00
UoKqGyCfslDt9zngP7zLL0ZApx+NsEnnAH3LCdsDk2H4LIH3gRbP5ps3rDbK
S+xFKeHFXm6hjg7veQbOXb4NnY2VBsM8alczN/D40q/gGA81QZj7aD9t7OY6
mvOhjp2QQIYmBX6P4G4xTQ9Spf8oNc5TBLLTQEYY/S7VwfqSjtZLmYaj4RTc
zqt2Jdwnh7lus0FWGiR7hvu9bYINB+ZWpZbAqdfqFrg6sfZg5RP06ga0GDAc
EcG02SpIJDWn9pG2KlN2n4S38kAH6jfZcmY0+Tax1BIHJJTnr6uK9NRMLGfc
YCSS0J/F5zFvqB3WCVPYdiTQ40binWzSFLxn/GWjL7GI3yIrBFTJHmJVCNy+
10neJN8/NxpuHmQKdeaESQpJpPZns5X5xkz8ScsZy9dpDOWcjwprpQ3WwuG3
3sDTKAfK1fUnOpSXy8Tj3u9alQ62JGDRU077iewfsvu8JuZcdO0C6NaZq2KO
9XNl5rvOWzuKBbVISYhfay/0C1SDSLUPwMEkDaeqIxc2iWm6NeUUVEYSNhM4
2GbJfZVMB3gmEB/IDGU0MFF15amGUYZNjkrQI+f9Ugz/d1qY4TiXQKph0ath
0WH0qwtt8aANRlMFrrRel+7MO169+WByd320PihsozZFocLJMq2jXhbW08JS
RVIIfESiHwuGwGyK7XijQswXyhExmhK8l9FrchV4XAG9OzJaxLS7I05odh8V
8A/30RKoFOnHkclUoBR3tA2dX+rcUSYpxd/3QSqjpa6q9TDGTX7kH4AKl5fv
cUGkDwDeRCn5n7qzt7HnnSBLQh6XCLcWq1kDaRdq0Ql64Cy97NIgqb1PeIMt
8OyRPA67mRfymHiCqDcpuUY1fAl2GjQaxTbmtJQgvokEaeWeiZNOMvwv4gU9
6Lre336KU+VVtT/w4EeUbS3XmzUlrKmlIflHwyM8xlD3YHQGboPW6HK3lUNu
vm0kr9rvovp/h22/K6P+woGSXtY5XTjEGv0wyHE09RSEfsTB5FOxnPtI7cUm
OpTm1DDuiPNgl9LXGhrsRkJQMVrKxsiBbXSeONZDDjSvsLpzPTDpSbIY/+1s
Y5rIAsROG43zlRvXze51tHUOTpTJg93rBBYl70a+5wUusqA7Ibqfqi8rdwUA
6OYc/hO3y7W+cv0XFUrEZ592SpqixCXoDWzVO3ul6Y2007O5WKLOw/XJNqIc
PNuoLKMeK6sEad0irmuZJbo9NSI3VSG6ElscjWGvriahHu8C0Fmrg6xzh6dO
y9FJh4ZLgV9kdHrvZTyB4+0QWqyUH/nFexrP6TOa1ccCVEhZSbb8rQBQMPzE
Lc6IYo2ldgZQTd5T3Jn6bYkaw34rikL6PxYIUXjFKtwtRWmtgO3geW5u6Dpn
7XU+YBAVCYmiu8uffcXaWqG/cVZYoSVlhEt7HkoW1YxlyrpxRSvaIxcUmTMu
v7fYZb4aRENHoYqZUWFCfP5Q/q5jbO/bRDlY/ILFIYHXzdU7gQjNeKB7PVyX
eJPo/5Su7K+0AR0yZxwK3Vnf2+wZTuyp+5jjeOBdJAkyXoyjjqnbOLJgQHpn
UA4y6sVVh4zuOo/OKqCpNYItFHBogZkL9W3obME6ZOYr6BsZ2oI/1ctSJo4Q
52fibeP7aMI7IrI9+NN4ycp4B5MRBsMGXcydj5FeLgwlnLKOl1KpMq7sW/N3
kTvlzaLAF+j3NwPnLzOF+J5S5dWYlAJWeGPaDR/Laxzvusmr2yy4aAiA3MWF
80ZwBTNGLkJwzQaL3uBjKpaKSzKBi53j8Y78bzG24tMVYJGjT69w0hur4lXl
aL24hjOSgkpI5rWy69/hx5CNbHJADHcQZHKUchtDK3UpiCX46cbYf05Q7Dry
Zim6QWHPPAC1UxUnSuYdZ9IcO++H1ZpzTCF7xMYShAurrZXhxZ8MzvpZeWZb
spZ57HsqF2Qd4clTTng8X5O61+j72OTlfuQmg/OrfoyAy/6brO08yUUm3A0T
1fEue4iYiIE1JR4REvLxsnYNjNCKLE1NQq9xqzDOAbvs8WcqSki2sxJByDn9
kCNHna/1v/TQqyuWKLR0WIVVrKtj8sGdGvhs0CCamOuIXn81L0WJf8BNveVb
H00YV4Ozmh2hVQQnbrFoGGcHFlXlVXmPH05nwmhZ4xJrnBCZkWwfHLWdDaWc
bFKy8pqp13SjEl2saG5dAHen2IDAIHx/sdfozyCd3D2fwnPXgD9HIGIdAx83
TrD2qPoNtXbuSAvu75UQtktbGolIHPSxCCnH6wPfiNay648i19mnRaenTyhA
Ro2STCkT4YGASaKwsHImbWmTghU9VN9T75JkYkl3PJnW2uS9oSCfskZwHxvE
5D1QWJuRsDtxeEKJf5rxWe5Kj+MUylgD3JnUcyYeoqpxF7v+oue/fFk3DL+Q
wDwNYL2MDNTrL90SsT/V8bi3IrA9fYjebdUW65kRUsaGjYvrYr6PQZOYgSbU
Hv4xS+UIpOa92bJzwa+xZBiztrxYkKlGgMuUikhnN0DjKXpcGI5n8TMHyFMj
AMVlD5MloBMFyBZRREdwYOeNI7Skq0t8kWJfLCP2n2nNJY63qSQ2r5R9i1gE
vm9roTjvZOh9SihCnjebtGnGLqM2jRqBrlKaQF4gFH6DBpHxXu03ZsqyQLN2
e8+VPyDPm8ihgEq59kwr0thyPRKcmTux2ARDB+xHWdt9c3c0JqbUtAzpKjBq
88/EsjuPnY0Z3MiSPEb2YjpBYrLUQ5jsfbX0ZHM6N0mh3rmzjR+MTmmPeCwQ
PxYBtm3COdOp5vue/U+7nrPR+MOccft2/awlej7a47FIppL5hPErqQvlgKYj
3Apyw2OVktvaUXcwFLg2rIeR1+p6JAy5C3ZmAdxAoc/SI7CxOQrvY+4srK6B
Z0QISxBSB0Z5J8DFzDBM5tmd0ka2gP7fRCCueEuL3VO7v1jmRyNSasJW18vJ
tEshiNeQMe5mBAH1qWIX7PanXfKbdrWVF1UAUoQ4g4oPS0H97r6orKPlJIvB
zz8B07jZmYcmnbEy/mYN1ZNDXzYbYgSssymZ9AXOnH83ZJozDOpNNEWov9sh
rhv2JqAeMXEsTQ1XISzfaJk1T5cE5GlfnCgP60R7oYfzkBZ/k0nRsyydX8rR
gxlbtsntyLR1wQOY4dO9cMNGKg/HqpztGc+YlOqnsxRMIw2tcjDgDsp+giKZ
puIcY/uh7QEBh3NMOBmrnE3gP9ewg50Zjkhp+4z7mb8JVoWYIBZUIb5bczjg
Sy8EnEF3Hrpk0OSzyJAt2o1PRCLtzniGFaQ1M2aSdQ9mZIw4tsOBH4z493Yk
FVlIxb+/hZOEjcP4f2fJw3fGer1MRV4NHaU0w1bJ30hGhXhAXlylWSB97JgB
SdWHdjA9aBLwRHiL/9/BO+VGYszOChXNxev/lGnD32vcPG+hIPFJUL9ZiyHw
fzASF8wUnV1mFXIzzHE6/zbooDprLsE/7AlXrVNK51Ew7es4mJhWfBbSAdoT
PqfInGzdKwjzpUsxNpcACx2GuNb5M+XPdh5lhzfvDc005V516OubW6cEe+8D
oMir2K7ULfcWimzXna5SMzFN1ljfAQcdsvG9vxPsTL9kNSshXrHh53MjMafD
BXKbZuN3YA1/Ztww9AahwZ5sV/0wl7X0W4F36E6PCvDYF/yLgOx0ksE3X63s
Meqo8Sno1Q78eVi9wTG2FlKGtd/+l1WocWwNTNa1R0siSY28D4puCHkH/Tss
EuvFbj2iVRD7vi5CuBHEBRVSX9/UEXFaa13ghQ8S1UpGt6uB93/qTWjgSkbH
9TFt1Y2uKOwzLn2X5ACdlyMb+2bGgqKfK2/hE93UnpsGlDVyPs8L7Q2aIXXR
6xsVg9emWvmYqHKqY2VAUiFaKZtTqdInrZunwBnBmlaaXZ+ZOK51B1SStL3l
8leRfbqeCpYUKqWp26Gkx2puHnOgsejaApa0IukOhMDKXU7Sf6YOOIAiIcme
4Eb1zDeRzw9LLpLk73X0G3jQuLtNMjKOKxm4X7g7q/F70k1Zs651WSxXTJAE
Ldq7GR/icdkyP5v3T+XitXaSGT/H4SuiA4a9Rqz2/SXZYi28noE7Wvv7p9QH
YAB9R12AUyzTdte+53zzfjBN9/qCayQGXkDi76PXJ/Gl0WXjrEpOy8LL8wOx
KmPPSB1oPpphydzIjnX+h4sLetXsrRFo2QYyYOAkZWrjAnD1lNfPdlBaQaXs
zBdTuUextF608QBXKVJVDArYDqa/4R18rWM3XLyQv8qzgAmT8zMe/Ns1fDX7
T4E/oB2gsd0kDN+kCm0MJ+G8d3rtobY0jUxJOO4F6Ns8HfQKhAUZS1nJ6uw/
gPLqq69VJ+gJ/FYgj6Ev/9pUzztMZh0rUwQ8h9YyLkjZA+9CUMPsfBmvOpYL
sVQDh8wNXdnxoGymxSqCffoxDTPMDu5x2Usfv/W8uy2rViMAfKzkuQTxjKs3
Z6uDj1LRUUqTSoj1q9GGMYRTCrZTFp8/HsZ8H+3O9LHxVRFNF223oktf+0rZ
ArA7deJ9bJlSc1w1C+36BUNaqH5jWmgAHpnH0YU5nmaDWyd4VEwW6qzWkCXV
L3qaHRnj7L/kmOX0//IIi4nHkaKDbFW+65negssCClpwVWaX/bTvtVYiA48z
Y4/hufHB0oeWz6Gv4N7XAjlXsVnxHjbi9jZmPaI76WYo7cD+/PUwF0diR2YJ
nb52CXf5sSRnnQz3O3paqulCHry46WPAQyHh5O39Dt3Kcg3+jivHAddQyn/6
iHs1E2P3SO3qNA+LRHYA5fpSeMbPxIsb5JEJNxrcQmNUAPmca5dPCIRShOTP
dbR/EykIamX9jBovSuzjVw0ybAH4hp8VzZP9+A5ghrDo/kYYWVoAAnJ7Xhc/
nqjDiZxcTQtcnExwhQWtjNDH7ojkWb1E9wvSRIGFkIZhUlC9EsFRRWBOZmld
IL6JrahDHyU1K/tYMnv+BAg84L/ctcK70sni6dQyqd7/aeRJKJPg3zlQzD81
8diRSmh9rhFk00njWRIxaSS5N8PpWauBNKrtsohzk8EeYmpcmd7AijncJxaG
XmUQR5DpDIpJxlpqISWXX5Vet6XpvUMHLS6e2+bSxVcsSnHz7uPNiTp48wRz
MTOO1WnNOKH5tIjN/D3JKPOcpeEw8lBdDmhI4amlx1DS9Vyg8F7jCvJsrhRd
0Lb7tDiRsrQlSeFWp/fu/Lk1hP7t7PG5ReDNN7xPgKugdAYjQ9Fm7WtRd5rr
MRs1Id1SeWS5hg5MF6cu+tDe1UOd6G0jfMp5sNedjNpj2UX24BDOvooStKz2
aAsvCs/KQ3wB+OkdpYyUtZF3mbfrF95I2jHH5Cq986xBhzx7c/o7AAcIfw4g
NE2o+Y7t81Z15vb5V63cNHA0F9fZPGpqV2kcFoWFCqg3RElabwZR1T0vbl8j
5aZW18g+mhEXFYtGwFCLsih1oeP1yqxI7Dv1NwQGr5zqnnKXG31BbBRnJepx
kMTuzsTSsyZbzijzY+uoeD0OfNaC9gvmY30HzMOYAW9x/l17lYF+9chgXGE2
2I96orVfIQbFWfAi4rp3bst3KOqlCxoR0X729YNXTBn21ePMO4HJ7nR85iPC
8+uZoBQuPeBtPvI6EqmXY7MJ1dfbXI1GZfb7PshiHmpTiH1SE6fbAdNSANye
xR5zMxCzi0w9ijsOUPZVpBwmyD026pA9bz9d6/6caZPtMHL7mExtaqtOR825
L2mGNmvFPhrErWUW9HA9E5TrHK4vrZ4MQX/sbfyIH6ZJE8+99zkUQo8Y2JGK
c+ZOThjSwYHXE1JaOucG6s+WVEjt8udiWumoCcoEDWaJPASUiT9WiIfaXFZ4
O0fOEA5wJZpAsJcSVL2kB50DMYWMVEhKNwxvESgVffpROGkZzt96R0Ss8txA
40vadZk5BUNCnD6e/tisiL9FhrKYZV+Qgt7WkJkUHsZd1VOEz91ME2JpdTeP
SMwiAYagPTysdLQRGX3XQ5o2hbXDLhuCf0OAoFea4iJXQvRgBUTbMjsWTBxH
qV2k+5yBAlKf1fOb2oO6AZihZBMVqQ51m8T00jjxjPXo0Z/4PLyeSoN2mA2A
5OcuCN5m7LBL2hGHrzkUMm9z4QfTtmarlrdS3bYgMlxlrbZPOOrN5+j3+DZm
gMNLkGpy4sA2zcXN+/ahuUI9XpjpP//SgyAkYCBpZ+7mtLJr6yc0hqoX4QCU
/I4yBNf/kRjBMpSfeZr115eXUpL+bY0avd+/51x/ibtOzxNQZ2eKcVHkxl0i
kSsEspei/6CTth6gj3vyaXDINNE8gfBpuLS3gfNIVbdYYKY5Dm5ndOG0kEB5
0GQM/WKpEsbDp0QhUTikf5dCuBtrtNTcT3IjcIL5mhPrP0veeAWIUcROHrAA
VMcrZTvFo8LtSrimPq2/b/k8KAHLFtYvSQHgIE0Q0fwhFS2sdkU9XvCUkJ0a
y8e+1pGmX9D48kzjS9LBo4PvHhGP8ED3enMhjZJE4EMTSsD0RKK9hE+LbYqe
ly7d9WtsbB5ONjQsrY98LFGhIozbfRwoTeXCWZjcn+PcSYz8VAb+BotlUz9H
ZFk6KsHMlZMf1dgX8HPAf1fxY3q34v+4OFZYg1hN5K6JAC3fowBDbhFl3Hi2
aGzvbcONtQZMAyyp2f66hyvPELx4fM76Inreleny4v6t7FtRhB1XDvtxDeIR
PfsRxnlfLq4MRTHH1BRYMWg7AE0Gge4YIqG1pwtLoA2OUucd8b5Hm+qyfQEQ
nc5jW6n+yID+uPb0PQ/z58jVT8RrdQWctEQLR7q67BEcZPzfj6+KkepPBwe2
1y6XXvqQa65PQUbT1nKPzABfSNt5T/Ln1+BJPXagItoF0PlL0rrroT8jfZyx
GTRF4HxTaVowIyLECHBBtbYSCQ06ZS8q9/qEDOW3siOP4pDgnp0/Oj7Way4U
xLuHWfe7yBaE5byiVROMOptxiJnRS/lHSBmfLGVSnx4q89A/NVgGvny3JAOg
com2Umr5wVqYM5ojrmhL+ohZ1DoqtVtA2wVbtpziwmxM4BMH980fm1cuJdBg
9zHqS2XgXSkdqp1hPk7ogE+ZoUBy04U1NhDmy7FB383epkAzy+hU5ShurN/P
VH9zkGdDLrxHI9GLfp+qPBWaEnNw8opJFSyegaKkkkwgVoj9wCpFbiIx7tWj
Nw/DQ5emF/4bs36q8ZfSogkb/ErQxJHK0mysqoLIEFcEj365TRyAuThuwvdv
7phIf8zPeacnHWj6PFlUUaGpj3+ld8wSFH4FoeF5XwPZC3Z505XrhPkqR27V
9sFWVzpb1RCz/walOC6tkrwW7GgIKRbsVCK4lUWSg6Y8tDxIPtHBTAkbDygr
m22qveHNcyLDkyh9Fck3r61yIY2m2I+BygIWk06ZjTNqFV5ylHYREv5CY062
Ivb69X7LaY5H2oWAlF6H4lNpJjuMkbiEPZvWBCb4yxzkLWJIBZlsM6OoTDM7
nlLrfgQWJkqjIf3LKV8JemNQIP4HT/mZLIPmsQUyxdVjxgrCUhmvP04bj3Zf
5opQO1RZNY0+Ibp/ZxKIMqzFgIOx+uDHmLG9bqvdhuyl8NUDPgFqUHeFMsZy
/+5VgjyFdeaQmRnf0mLvoEooIbF3ZR+gqnnklGqP+LHXxGlNXdodK/TIQ9h4
Dkqi0dXtaBoGIrotQTp6tj/YM9QYcLL1k2J+FmrAIiJTqBOGcjeecqSDOZjM
WO/mKdEL2zqqrVymLEFTm043qJvIhtvCfDrEJgJlDDngYLGZAC15pwC/hXtq
WXqnRfSanmIyxxel7CzL/NU29NRcAfAlFkI09zukOlSffrGS8CT/tf2xWooA
AUMUkro8awcNbASWqZ502vthU7Pnw9lOCwyh2ZudXHdbNqRj45pEmn/Lkrhy
U6la28dGsHjSAsuHmDN4d7RYKklB5q9Q8gQr4a/aRuOLZTgTLz4lZ+QmY7gm
RZBCpscQ71GnM9Lg8EsPuiyZUch5EMbdUbNX7SHAaLURuCBzhSJKJgQPHWGz
gOyEf/tR6Rj0Ld6USyG6lfarr/01qSnyPV1A80mzzjvQmGWoFdPzloG9GzdX
ZbX0tVOPvgtBLgoVs0tS7/5+/qUohNqLohGdZuJ+Ko4Ww2PXrcJQju/CanEC
1OS3+SJ8u4Q4elaKoGjaF44dv+pZYh0mE2agwk91mN3MDVKlMEM3b7aaH5uu
lBuVQ9j5+uxV7ihmx5H443nAlSsWtu4+Dl04YcuZVpvPnA+UhKNgqGzon2rB
eqMFnutb4qANrntMOBVdCWd3U+Jx0fW1lKcdEGNt4fhRuzo1oJa2qKccm8P8
nLYyBHyPt593045wkqrNbBZBJgSj6vLlO78ZLCNMd8hJoaOupgzbEhcNm19W
Y46q/heINJ2thiQyH+ewAP70G93LPHseQfkP4gEOsOYXdJQXZCPA45iDMvH3
Vs3IF3hsadJwn7zy2FMQEZNVojwXtV6uhCSJPPeJuom3CUB4ckxIV2bNwCC1
0BjrumqbewB5x1NnO0gEELDr91ouEFBbo5sx3RyDdFcO5m42kEN83YMvnL2X
+reoCJi0bygmqhBFZiCpt9dSQayufjI8RgureDaq5Oqykc75CYiQSx2ArYNw
9JtoB1xYr7i+EXIH0mDbudH7h/ZGOX5b880ABppcaXx6BmFqTOX2dBojY402
15/TwXxgNFIels0Qc0b17ybPyrG4dylJ4CtDLh3Se4thFOHpVvwx5vfVl/ZP
kgbuw3uWx8b4xK3lkccpadueJYR1x6TM2FhivGALSttr+a5MDcDRhZSiHJPg
SxtgARxr2DEgnaKkGMUjY3YSdh5gBB5+Q4wLA6JYawKYjsDUUP7NOydEb3q1
flyglpxSB/m12JNT69hLg72kdjrIGr1R8H9WA+B8cZw3Cb5JoMeJeaLVaGTc
GFv8GKX/mn2DYnI3c2vmPFTkkD3Eem8clBeWcLJK4B8EvGW0goC1zG7NTdEx
L4tI6XVpUSparus1BQfCi7f8MGYxhsRJNK9dspyaFHEZVQEqNhaVMVHnM2eu
U7869vCSEUyjB/F7wYbheuiGrfkq37rLTkzFThuD8P+T4bXTsrVTBTkGYEb/
tIdSjTNf9ANkTN8WxpXTy6PQSjxVvQ4TF/q9dFc1eYziN06SLFSfdq7NPMUU
cjaLwKmXXh/KuRUS7WUAC8kmsn4XJ3VYR6w9nPMi9UVs5uV1jQNvbmfry4to
hywX6MhhbkBP8E+Lv1OMp1y7h1IXDf9dwMcxj8GIOdFaJzDAf+a8BuIQ3AuX
gjFBhfwyPDEuGY8Km+ZMz5ji3mUzG/y39SsB2gmZA33rX32rKytwfK6dI38a
/slQ/enrBVsCHWRpUvaAsEoVbT0srP1SXi5BvPOvLCauT07A6U/hb/NTyejn
1WvTwMJroO+ucYnIv0SpaGyRlK/b1x0nX3Ppeo1QvKGguQ+OukcOmSpxyVnv
PD6eo/NgfPABhk405TTWc30obiJH2N10NjkVoAf3XfDgCk5ZCVJeilFJrv5a
P9dbbceeVox7woC5GX5Cu4+Bfh4Ut6YyXsMjZ++q1Fb5TiILFQ53bY+D7hyK
pnj5l+1YG9uwMW7D2fJ3M8zN20llcaZlreAt8/f4hoCySbkKombQ1ACgmR+z
ws68Pmg6mdeF+3kCKJkwaLF8UWMssUOfrh9hIGOLKhGCrsj875+Lvxpn8A23
Ffv7lLI8EsuakKl2xJJdXZ/aWFC2ZEMtdKvQDmwlyQts6MRqiX1wjIUGLIeO
c8bqjXVZOo8Ha4QOiMqNgFvo7chE1pC0uRpmL2SjhD5TEo+r1e9MDCRXKCv6
QUd1sDBn8tDMQt/p3ETYCT+HnIfEfLhio3OUYcLsg7YUI/Itb+93Azfw3MLW
MXAUhyJMhOkehfCSesgrg8p0PD9kr8vRF334kbUC1zeCJtlvMyJfx4mO3kIg
g0NmChIMFKEM5p/y3IOVxnllS7XnAeXfro6zlNgf3Ivh9CI0WCvtXVxSCcBn
4ThbE+X7sFA752KQd4G4Ku359t8DnEgdZrEZcbQNpXpx/i2WTYZ8oGIq1ppE
D9g2+oaxvWMTeFd0WWB3T9ug7pzHVAbbBjwSl/YSWBEyMMAOOG+mU6cySDaP
DhJoEa7WTPCYJy6vFudSyf5VCoPtbTmGfBifI7xofgM7szfDsCVEbxz4O6GZ
A/uLQHf4CRfHWh6C0rrydb12gWjM23KPODhzVKbT+/MlPsvl/hlgTPXen9ql
CrqTIAHl7hETurfrR35dqPY1mrRpSw3FJyLIX9/8J49B2bfQsuPyaGSjIbdX
TnkopMrf6+mKp3yA+z5hBegquOw/G8WWwhoS/RJ+KMajlrg8XdeWeS9mRu6f
gL/IzdQlCGjWZzuPzdPDOzNQI68vEyn9R207etWIyCiWmJMPJ1IvqaRPR+3q
esYELj0ARouMMptwQYu16DpQnYbV93Fr4/YvdWaNndDjp+DP+ttbKNb6cHpr
nbZ+F2fBhnSQgg7wFWbLdmKIfrcGBQhYs3qP7wCzgEUcbL+8lrDrYSpNcLvy
vfCUPF8hQsP1SwQzCznUiHVI1Y9dGnpvgfSEIr9lCizt3gkD7FPZ+h25TxYQ
EraEiCCZTD/A+dZSfGWk8t8ZfS+YwlXF929Ap/GD4fCQcRDQ+Si4PiWWXF7T
OVMliX4HFu2no3iIwEy+rcrCyIPUYNqsWVI7K5Rd8VeBf11qywvskkulSHkQ
IemWTethVLw8FUWaAHJrub4wWWHI0eaS+gGnscmlJoUzQQJ63Yr8NLR/vmf5
RzeWPjNWj9r4PYC7zUKYOd84/4Nm1eEMnq2EHz62ByNM/0aKPPuqKI4RJje8
Q8U1kKr2bLPzPAxZlzmz/ngPKlwUBtmyM1X7I3y2f5L+m6n1qJG4Mbq8ETiK
8ZBic8KS1Ka95LS2OpcjYKC+/R8RsXamE1yM/pmRbE+B6YFRbKGNORjkCscE
QsZAT07xauRTtADuWwM/pIGO8bE1F4YjWlrya/rFH1oFUb8aGGPsS4gTSc1f
5V5l5/41lz6B8rybwM42mcBz1sLkpMlp3g6xpTery+POqpipneiQ4hIHUxZt
uHnNfrfEqyCYgpH0d617S+OfUyR26WWO2hn9eafO1MYoibE421lydZ9QBOXp
YMf01au+ef3tCAIEDexBclu5yivjSxb4dsX//MwydFrh7BZmOpUS2W/QG7OC
wNTqCm9UwzhSNS13egs2JfQzB3SzL4/itVhg7FIM12Y5oKIvZw8fFFfaXHOy
M4ZL/h7//yPt6BoKPdY5e9sW0/N6QvvdrNo7Wk6TiVzCYut0YqPg2BkXcEpB
AC8sK9ar6enqpO7cWeQOX7hr8T+iVQU9hByloT50JCBB90ZndCgoti8KU+BS
tY4wXADkYJDQ7FEFE1S9KYHrwMznB3KVFIqswxQIWuyoojBZukc2ZEmEp8b9
GQ0Cmz4bB6oseVxm6tdvgsHWYKdKVMvRb49aUDJ5jxoJ+k8JMK0gr1G7emj7
qoTrJTwk5azNijr1zxGDaP/XkX2xAzt/43gTtPNgEvTCwYHbg7sGXX00+gW/
KERgYG8DFeYCaoL/a6LyFxt/DNa45J9LJpoqCcQUXiguBRRfebArtdFSh8sp
CQEfr3l36JlV9XulYJvozLl2WsT8reDXb6NnEeOUQwZ4zZk+zDSr+sFjKRaR
vYz5kJAMnh8d15qWG9vUkcgoq3zn3dAA/fxKO4TdfBs1eoMyg2HI6BqSFRYo
2DcxsrcHYGVYJJVDVUHYzIaDJKuK6PhLt1GNYT2RwNxVUqncv124oIWvVqmG
XWFN+yrdOxMF+WUcFZhlDovsg06kvngeMNyG2i1Fqv/KIho14yTk/GRq6qbz
s9o5QvqSsPoZwYDFDTj57MMb2DlK3CBEWwFX7b5W4QpLe5/UriekaTPZL7eI
n04obRENJJuKTqbqcCpROIzrZ/K79HYsm0xSHLyzaDH3LqXJIIYoZQPTZbl8
7N+Ya+GwIIgeKPXwWOOkuBWk50HR+wZivIBZnniEHK3az6wmf9/G/VCZpyF/
Sg22DSz9AVlDIeIuKSGUUipwalXlKkYL7sqDjdBSS+53YcsJIggsiufSJj8c
NfcRvL1WsiD8R4fSqfNFStlzZ9RAQDGVxkDQy+cf5m0dqRzAf6bHyKwGC4oj
ht5hZuVO2XXY6Gspl212wpgJ4CbYv+LiTNZlyrtcRzUsHHBTSt4/Bzuy0n+B
BHdVOCiZ75nbBtnadmE9V9K0JldJEBXRfCeQ3Op2RZoHws3gup2w4hTl4Pqq
ym50wTjzPXFuOY2YvZk+B7XqTbvo5pVK9imcxqgtpXXYlJ/d3pN4+nMfx+DX
spFmnf0J01wKbSMXZurEj7ykdvTMYuvtRcCuVikb2YHYHefwrmuJPxKqEd8c
yHMYiLuhryTj6JzJ7zAslsyH2IVH8cz40E2ZcgeaVfQBqQnpNQ9t81cclwvJ
pwkDaM+QcSw3zfT4r0ARd/JjK34rCeVvQz1FXPxF5deQ+xc4NlY0lzpHUR/m
6bx/6UrTb0frt79cRpYxBxObT08TRyenhxL0CZ0q07cgckr0k65omeaGx8uw
btqnJjeCiguJ8a5yumTWWpiHvyOyL7BDdIgGroi6ANFg87sHXXO4kOYASoof
XsEevyJfkqwJeZaraUKuMZizk5Pwr+iPh3xlk+Mlox7oVBKny3CONh0t6iY5
pV9XprlT9fTozyBu6eVqnJECA8faC1j+R1/Aa82/cFLjhVGYaTFTqhtjD8LS
3InzqtSuJ5sDX1ZjNuuZH40WC+inv0BST8g5x9t42aQUIQ5rgVju4W+P7MFR
JXT4T8Cv9LNfI3lMHZYqYT8xaFp5KDQBebzr2cgpDqrIQ673vHGa2+lEATZV
hxr5m98cdPIhiAKPtzXviRYfQKFVSHl0EXvn67iv0P+J4wrTOWLby0jLrx/G
YNijL4kh7gRQMZkt88xeqZhD0ZLV/vpt0pEIbvZ9dBcgQ32MQOL/nIQMc/Vf
VsAmCj4npIMLnqL6EVXXnTKShMj+2uHimRjxxShxM58WGyLMcgiI7Z6U2ZvI
DRtffK8oZmsYM5vqnPpvEd/M6yyzQ0FD1+bz0BrMLpiKZGDnhDKYZxXroFLC
6sjANamGQEwqCHuU1cHKoDhntsFfZy4thh9QUD7vSaDEt4k86HCtJdY7361u
Rmz5I/imgheLAW73x5SjXK9gfC/HxsW8PEuGf+TvJZlVGw0uxlLzYG4JvsIs
RLMJTSkmhxocjuAbjVSODl33ZSRdwNvZUFR7HgYOk4KbmqyAQ8NWVTeOeuTZ
zIO+6wcW/YCmDUGv2de0THxfhbBCeJYGeh44QD3OTQI1HJtSqTcSl1phI9vg
qlCFy3zYTTkS3Poz4k2AyTfrjKXDX1wDOSyQwPYcXl/viL15yCRdvoqGZVaM
9SDEhpkU0JKL0SleGV9P/Nz71RhgCq4pMjaVYctyJNvBjsXIhOmr+fpcshfR
Ym/5RnSTjGAdYehkwmB6NeOi8wuVePvUDLOmvE/x15jYHPMlSQa4+3ob4qJ4
ULAiMamTBepakjMFHtX9k9RGEPzgj8SH5cUV9gGzkGaiKqSt9/M8bKszWeac
NSKuiexKfBZ4sLVCpQXK3Wb+aOrlL5g1ijxVqy9Lzz8ewd21hbJufpyQk3Rz
D+ESfGmXz4I6tLsJ1vZEYdURwoOgPrfw/KxU7KwScmQzr3v1GhFAFg/0b14i
38sF2GuLHmdfmstszIFK2IIa3R6I4Ww7V9IFzs8ao8xym/BjQOLmkpBUxhiN
8Bmkg+gy0RLEWlwsMGfvLKzGw/zA8OO3342IST7S0oFn9J42OeWdg1zcILp9
0YtlnOBuuMa3NwFxDRcLt54LgJ2GQAXuY2SujGbJeCD4qIYRM3wwuwRKNlZN
hiiWVcX+wUuMpXf7C4OqkggWieTBXbYVr1hpq+ewGPiZMdT1LiwMCJdTr3Nu
fAOaxzSyLmMQNXbru60QGJCKd9OpBB3BOH5LNCSFLjw5sD4XwHLtYMWTJ7K+
sEFaP413bVn2hX44rHsVHVfM2fnlQpqxLseGTRXMyqlgYcfrjsBaGBDY8ZK+
BMS+uBrtwVgFo1jsxZ/4VvuUSGMKpAJUcOozuhFBzpSodf4sNNGxAZjYubRD
fAAw4WGCn2aPyY+QU0VhrfA2vBswEs5OAQ4fL8yX/DZJUj4U94WpZtmKHTZ/
ybRU9fRYcNmL6ey7lHHpZhbBIlV4DDcnTATNxNp1eHOhpTe48a1o+HmuFhWK
gIKMqJhKRpkDUpbcfrOY/5VVSNx0XW0qLOyHjyfCPyCeWX44tosm/MWspjUF
6WuldIYIRyOoBoMjwTT/i5+hJosdchPATEvNrz/eEsh2V+UfSzlbzxPFIhPt
pTTuym9u7vOWGPANL+Q61PfU6Gxdf2DAr9f8WCZrpdLP4CIv/16xwBX/4eLW
Gn5zqaJ9BUNGJwc2dgoKnjCG8xDrEHaDsZzpDwYd6j2c1fmUrU0moDHqormc
Hag+fnQTPel5TYZf/nd3V8Na4KfHw/j2TRzoS+D0XzwzQWQ0kodzmrs1XjmR
Yb5e5RGUOH9BUytdDmRALG7K1cw1DnvIGxQjgw8oc5lSJxzszD5Iw4/8SykV
jfHU1ngaDxnPUaUUjPIKjwzNgYneH0xy1l1U9kh7JdyzIQV8SC9PAorREx2I
nXgptHHA9AYqo2LtWXkfMVLmTnFS8FY6KClfsYchKfP2bykdKcxwYMj0963V
WpJqHcmF37GoHpGLtJ4fMfTkVfVtdG4NMQG55zB/i8quw+eZGX4VdmaAZu21
T0TG9ZUiQq/9mdvD6ahpSjW019MjQZhRWGgZ331luxgFOYE1wHXVddGPY6HZ
gv3JiPEfSHmF/epve5gP/O6OKrX7Adm8gprCZg9Q15Af4seJ6GqZyIyc+8k0
SKXA1lurgptR1vsxcu9jS68JfrUQSO99y8Oo44uNZeyBIsUkX0DuE6yCjnMp
f0uQ1dffbtQnWiKB8fAiyf1MkYQMfvvkTjV26j1axuIw1Taz7Cj4yPf2x5/i
fnK6SpJPpmtpf2mzGimGzjtlbd6w4Yfn5jK5Op8m1zJHG4/pkL7v+IASO6Yz
/zEmXCs0y5BalQ8Y36top+slQ1Hrf8+rxTV6qyM329t72g9R7JHZTjENonV4
mBF4irUC+lHOwK7dvxAClBaBdzvsLuLHkD66rpA2ZGi4JqINWa8JJ24wdLl9
qcy+LzpgDPB4DoEkFVeU7F8F4/oPh4y0Ltr7scyajTCIUybaOAoLQPNdNS1o
12AgA83VqDMQstEoILk1KJjbDl5uehW0J6b869NifWpYM9eZdvqb/VItxKfA
Y7MUum4HMa+CsIL/IsFCgPAupj6jfqQNEghOI6WyFODSRYcP109J3F/xcOEn
ATSavudWQ0NIZNUaFIt6mcYaneeY7cn/WIQZcyC8mTqyopMSqAHHqyG+e+NU
IQNgukcxWyJgu1Pr1PUcV4Jm0wsBTkUam0J62mziHXrMsfk29Q0wXuTDs8vZ
Lx1pc8LTYnfhYHh6HZZ/Slq7jCeh/8fUeqMfMsmddYUAIBFXPpSCIGcnuNSf
nEqjOUoWyLYjfBW0Lz/razoKYf4bvmwMQw61kjyQjm9W5Ou9ouiS6IYXyROK
AAHxgghU82WwOH5pRUUVjLt6WFASqB/eNs9UawB/BXJnH1s8YfaY5IJlm30M
akzMIMWXpI4aPTu8KTRGOWilr40GnS6K4htFSZewMW6fhMsKKp/2xxZHxDD9
TVJusl+dQ7MszCWZGr6JpQTEDoD/KuvEWBtyPsa27sooWHifsRjOGV65796X
q2+KpR6O6BWgolxwWQ98Rh7yCkiWNwu8jU0+1zALFyz2Y8ppzayuR0w0a9Mc
7a80c6U8xWWnwL1fvRiL7xIjhnTHOCkpQh5b9QH/cqjvVGXbyKIv8tDqbVod
3n+3oU81UD+m2bepOjTAUkXcfjyjEwBBAxb+GbIMrt2YpMzvhgCpHtFQL6Ws
jXXFk/n76pPQv9OZvX+4nwesDi3NF4i8I9zf1tZ/4ALRwi4AJ2VyLnQajKyM
/FeZQkpKB0Qmj2FGr75z6ni4AUK22VkrOxmLCv+FW9dxpAehyWZR276AL9gd
N4u5ICV7hdYhZoQz4FqNeTg5IRe1pp5CUn28V8imGQQQby82fWP47CsvWG1z
dXgnJeoOcnbV0BLlWRVw7Jm5RtDk/rgsagOBrMz9zzOSYVt3CxVpQqwizm9V
Ber//RYlk+fk1z8rMWiXFyRTG9/94SkYYNbx1eco89MwYvPsfl0K2AyOEEYN
wSl8X7th3A8Ih9XT261pY/3B4trafQa9U8oTW6u/2ErWWVnfhUFJg8gb5xq6
ArvHud4O8wEWtMlb1ycGGbiQl5bavPppzemc4p7lL5mo8KfYRPcsr6A3U3Sv
Rx4NcfcjUJZDNZJkCmXxbVSjpFll9zvSoiui+c5XRHFIfzNswNZD3GVo2H7D
Kb4KM3mjGJif21c6oJCV3P9tSmLxDfyhHmcDHtTWwkyFKM2+8pKAF/pWKOTu
N0G4jD9tzXeaJJ1rXtPnT+2ypSzd8+YO9KgWQnmfQBh+r9d+doTtPuOAWYBc
jyXkWtUNGYawzJIquL4z4uq6G4787+LosR+z5YfaCSPyNV/gQd+nbjZwh9Q6
BxZBVu3YER2MFhD6Pxd2Np9mFxT+Yuz7lHkJL3E9qLz/45dLl0qzlg3goKqY
4fMByXZwGMUWAPw0ERbDb8rSLHTccjw61qTwC82bo8JAAR2GKMApq8cKplzI
pvhCKjeN1g3u49Zjn2Y60OHtZaxUwglJwiVi5UznfCqWIv7zzkWIpSfEFeAg
iliLpk+QB808hHJ8IS0AUoUjN8VDurI6AkK22OK/d/vuehWx7ADuyKL/wjUW
iXGtbq5UoHtvJ/S7RmNjJhfqnEcs1NVBvRe/M4DBZbIdtqKanj4v85PIjtxi
YuKPG+uzxspI2Reo9uEMuw/iDO5+lRcJAvYKkaAC9eWx1Hcf1qMkP/n3gJ3b
vPO4WMKGB23rrx8dKKsM6GieYxdPPjMmCULLUSBkFLr2AFC2HKeKLw/52nl6
frbyS4kIWz3nj+oF6wDb7Y/RRVwSMsrI+wymbwEWGKPzOPfkG+SZLWJzqd7v
H9vtGfPjMUlR7u6tH8p8sSbIDxEyJW5j06NhuwkXigpS8C/BiB0JJE6AENmH
x5TTHM4dLjqqSclIBoidZIUwPM7844T+wOccVnUJl5NpWlBO60B+93A1E3iP
VPCHJnCb4lFZujU0nK4Gfzid+3rLyXwp8rpXs33dlrYm6u+KsJ19CAfYMoGP
GodjetqLGoCJY0RO4ePinGxTK7Um/cj8ApYBWkankzjMDq0CAfi/1AlsILXm
GIjmy6SqN8ZA6lUOeLb+fX/wzwA8H7ES7tTBzFBLrsSntdPBjwqCoTbQgtNY
d2au9oAZEk+COui1yh4I125vH8uWFPtD2biHBlExqC2OHIQlaqat481iVi1o
YcihTdVVMU+7RooGv/dKv8mro10LuoYtIUF6uHil7ltTKl2+Npa78Sg3n3NA
ErQIl79KC4WNQMAnYBDO13AQmQBy3evSe1CVTiqRm4qlFshfuodP1bbu/Lsk
bUzIiMNrLOHEGWmUQnCeC8sJ63C2LW6DiS9eqsWuBMKKZIv2B1hsv6DtPfGo
GXSiHSpBHTd1VhGFsmIHwjLKGbkJqaJuYTu9J1M0alaoL5IGhlbybeTDOk7y
1yc1LhXwXnOJ/E+ceWqyIFhUNhbuCSLdWssZ+RpstfC0DMFJsewg2QyxaWdV
j1qrXppSuiRuHD6OU/Wim6x8QIjNDzD34S/E4o29sjLOsCR8gFNoVRfSeFDn
Nn/9KF9BywiwIV0Zmfzvph6oy+vDUpkZQq9kLMygA4PzIRoo18Py7M/Dj8Cv
BeLxXpIDt2qKt/bzLH6CU6cdQHrDGdCtpKR6d4dABFjChI6JyqMJY9Bxp/Ct
bMKZPY+SbGhILpJuO1fxcKCV3CNDCWaNNnI3m1TJAfI673aoGRPltME481WG
d0gG25eBfZJqGtTtl2RxPR2WVLNFlyWjFNq8m7bQ4XUoeR8gbw4QMc2L/f1n
kv2G1ODfrVxau1lBhTvNA1/AGqmDIZYe3ICyAg23drl/YSR2Z+Kh8DQRT6FX
aalpNchUXeyba1LxtqjANq2lO+crk0bDyqVVp1oHcDdxbbRW+UoWnvzRMsJP
/rRYg/0OXSFx/r3OUGEWHZcgNmzmLnJhVVfpiJ32xuou+zICMXwgozwGX1xG
XrUp2NFht5+W7emIPW4PqJ677OQRLmlpccxoOUNxyz7c+S0GL+lblxe7u+Jf
HxWRLNesQzlKRjnpcPdy0BbPwHQT9pWsxIUT40dj/+voUp1Tj+NTWadAFwJx
YC9NgDZX7u6fUpzugAd6NQFWT+Eo8cRzLw610VuXw0GS1DVWmBVX9qv6EYPV
7xCtJwgAcdyTYXoCfR3t41MLGOGVk4/+TUwT1vJ/JCfhEg6tfL4ru0vuNoKR
ikqcPx1LKBdTX8B/xK9UO69JSiOjCetky5g89AdzbUqpvmSV68h7VSQJ+2S3
4os1mppER5+GXrYl/jPqUz7lGMnHFUQiDc/HZjb+RLZ1HkfSHt2zKFAob3G+
KgmTBcrfHjXjrVFHH6OE0gK5tg8cxGiyb3VWp3CPuvfaWQfGNnHaX1kqo67/
rSaHZAr5L5knfFka9EJfxC9dYg5hR/B1WmPqcBJXfVFDoN/FthdJIcXNwO60
7cGCa52FSHK9RzLcllt6RiCi35lhdMMS29eh1gGwXWPIpUCOQcUe37lkMOkh
SyJsaeds+g4hYy/WwwXLKA1/sjq+qqu5Ux5OqMGOREHl05JKh2GxO6E/KzWK
ibjpf0t60kgP3EfRE9CuMFZCmB6Nss3hiRnS4FBcGf8JIjx4WTIHfRmDj47W
k41z2fCPOUkEGGJRCrYz7/FObcfIWtOa9VaS+alKW1F7hgHsrZLbKxrcFgZw
a7iBUC+hysWEUCfbNhJmFyVTyTQOtYSalB4HHljHxuLJ0S8n9E9ruoOvIulg
BSyL81ApRUn+aIdWL2C+Vuq+N5h1cLxu4P8vAr4mxqJzWTvSlRhi1RVbu8OH
68BDiR5+LpFJ5yMciixrj1D60wSlZE+KjBxjk2ORxgBiS5w/hfH1PDhhltBJ
JcctafwfIZo0f9HunBE4DS31kuUUeqHCluSNr+BgILnDcXuU3Z7xZrsg+Ghr
t3AZnfzvJJq8yLTBbM+BoY7viorm1IvkmMEN6URT+NaCm20CYg3KLoZRyysM
sOdOOVdDVFFlVp+Cax6cdw0J0A1Wvva4WnN7xmO3NBsGMiQw7nwhRHsb5qpL
ZziJq4+QPcksosqnbQdWgWQUsms5SOfNyabuUbMUvUdjABm7jBpK+Rrvom3V
g9mOL7dEIa35ZwYbhmct75xC9XMJo42V4NxYyu8lMMCKnqWEhPm7cJR7tz5M
vd7o9rVlzMwZIoiq1tqGtU/mwWVhxvXZR8DkyMFMPDBlUkNoS19IObPsWBsg
tfx9WMnxDyNrZr3zdp/PmwcSFoJZPGCOlIJ9hL3Z/vA/TUIucm+zU46IlygD
tN8KIlkmI7vjw0ukR1ymsvcN4Bi9NgzLJeY3vlocigtNryrIXWdVaUKGHyMw
l84uTeQs9gcYrMZMxWI+vMJijKhl7voOctuqIuDk/Qv32yJzoRvHmZDNqi3S
rv91UHj5JF9MYoxbe44MHgfz3fD1wRyAkABBXqQL73moUKEBHQv7AGdARAsj
+g40S2nDfS/npNm+TMEBQ+uMUx/D88+h7AAOOn9Kc/eKoDZP0n0Cprp+iAfu
zgeB2MSPmRlk/SrIfjAg+zQIAUUY07/uw9dlDRH0AAjMcj3SopcymOd5OTLM
CHXF30pDxD4UN/fWbuUEMv5zTUTiHgkxO9R3ZaViwGzBAXURd8bL9hgNNiPl
AV2t9vJBRtJkEo40FymYR4IcgeTWtwweO5H44v2uSHWFATzD9lekBBRe5B5d
nI47mybTY1RamhL2Cqvu7v407SruXqhP9273DD/0AYWcV1qOKHE1IHUAF42f
1BZ/fj3hDt7GXDgD1N8xlSw4glP2d/lg/rHYCZiW9Op7qNsEhbUeljc4lxtN
9E3gTpyskPDQBwlZSgmv7nM7g/W1UWsqefMEXnecccCm8yAP5w+Nxv3hPrjh
Z1F4hNCE0W7R+BiXCE3dNMAnHfHzG9Ou5DdgChHb/9Lv8k1nJPAsv8dzPUtO
P7w04BMkeE6g9UmcDGL3TDGmyoX7oyTt2Y/2VWw7Tl2k1c0UnAej51wz+NyP
2EMs7kZgYDh/Jk29ZBYEnYhDqMYG+O3oLuaLnDXleTQQ0UFrAPre71oYi/+a
KZTepbTAMUBqIyIc9+rVOiF1zTI/5G/9ja/XdpGoA2ll2zAcUuJy8hb5FpVT
YXQCostdFzNAef98ilO7SsDlxoCFliCu88FHVTT8YOL2RUwBtqS1HB5Rb04X
nNRD1GGxrKpLm5uj4E18pDcVA+uLh68XYEgA5cSkMLtbOk8cGDoQGHvfS2jf
h9i7klQcRuTAzGtWr8X2dJkP23ekVdfzUB+WaQNzJ4dIfS80Qz4xQ9tykgnY
qkHhaEG931+v42pgIwMuDgg7pF84KYFkF6SvqBeIW3QijSNDbje/bDCKL++m
BUZD8krOgOOnl2g3yriEygSvQx57j9jVrjbvHAwkLeOlCTiQ7fGHmq5tPt30
3jp52L4TWGcFhA0kJlfby7IpjoVTHHIMn7KV5ae469j2sdK5M5liF+ENa1MA
YFO5dYsXAmmB4FSzqYIQ3XNTEo/JdWRooTMCqq0zZxo7uedK/JRRWAGA3rDC
bqJ6sjh2BajNYaJjIh3WVt8cuFh6+3Dsq/S/P2sXS/PzYxY/cjrq3ZYxjwd7
xpuPxVYaPKq7SrK8/vTCGBNa4YEYN2tPs/Hb+jcHL199hW+dFzMpGES1QptB
1UCsPdsZra/6BwvEcebaGpfHBtqScNCqyHQYuvThWGoEtElLt4QtkM+8eDCQ
mNZJlZuNbBAJVExrLlhO4jtic1u5EfJ9ZqOEWfqqQLuJy0zmGYgEBxZYZH7a
ntErLENe/8fx6OgX5Qw+956inPjqYhHRwFWhX0qZc3ygotq3btgYJKIqSvIr
+r+TKQocrWiTCCFc2lmmW6Qg6i91qyyvgZ4I/uEE1NmLv3B4pMuVuwqJ3MX8
oLCH/kMl2OfBCwGbjRhuSFhVhKDHgKLERgHv6RUxEKTRUcM2KvrxHE+TpGex
lXab+oIuXWe6QIxZvqwXDxn1nBx2nNYxspQF4kh29M5J47FaJZkPZztGUkmX
bea6RtxtOVXWd3sZ9EJlUs38ouMQSTLS/8RNQ105O/aKe9txRiq6y2MUKEyV
o6iEhgT6gOf8YybX78qcvPcgfBP5baUaox5CqvW4gHm9TDeGm+ca4bWKx1wI
LCazIrw96pTO6C2hKtVekK5WemSzls3Z1NAai423BaRs39/zwg4b4Sm6+Y1P
2NqmrARkoZVgFIxFfwxXFM1D5cXFYKooVl4tx5lom5OOEhhTTHkg5nG7MVf7
4V0FztAp+/gwUDhyfAVHWC9Fn52ljXFLo9kIa5lNQMWcuO6p1aNrvi+vDBFz
yZJzaUWWKfHE+TbVr7nQuApMCvaWY7xalzQaRs8LwxdIW/Qdyz5uLjJ4M3lb
gI92oYEobTZgMlN3KjDrk61DvbiQIm+rd05m/K4HINlimNu9vYuGHgGVE2I8
fINB0w1pUPtNVcrL+rSUQLS5eXTnZJiuouivCmnJ47wIBfHeqa3YcGw4M2Wp
0GRzlBoYw1alkO+nnWdYqYfvVpw+d0uAcXNcJVgpyKsZSPT/xteZ5aZ26Syy
gOt2iUDrV0ib6m2ZvGXNuRZ4CZkfb4giGL2ho+PullJ0+mHo/xqob55cEjLv
EQx2JvmuingJx6uttJeAGcudWsHuyBtvFrfnWkZ5KQ1Un1jm+/AUAUuzNlU6
effZu+c780RCma/G1tGoDFeSIfCUblq7/ftM17tM0OhZAlgjwhr49nSUESAh
H0d9dtb6TLdrcKsxLBOd7OvltIDzZy6Zy7HovA/eTxm+r2h+wgxC32WnsVog
8sHwi0b+MpLwheHUcI/4xnSd9oE66p5O3umvdKOra4cUo/K31hiVXO7lMhDY
sZ9u7oi/ntua9Lxcgt7P9bbjrPB/YWKgpHpgaJWVJbdA3y1+lfgozVgY9Em6
C0mtQHnqjRH4tXyje2m7Q3ZBuhmW3LT5o2F33ayjeLi215S47DvcX8r8rTev
jJ81F5NjArDcEZwHYSxymBIFgF7vIBcC7n8vcvhusRNuRHR9qzRhM2X61n4r
vT3v5vNeStWdmUwEW9QErJPE8Wr82p26nCvRZMPx1gAUNRcH/UTR/Q/1hiO4
o5Nf6cd+VyyQmTkTvQf91jJiQQjS9LLsHqCCroyU2gd9IhmclR22YwzUrZhJ
wQycCT5ofovzaNPS+71z7kDNGAMUUnLp8CkG293yEkCp5p3BssCjCs3F01Uh
D8MywRjkO1WLn13NqQ/3BpFUfbHqea/X8NyBgMNai1TqPjJRwC5PZkXXgVF/
y5g0/WIEWAoxgI7LMm9SPpPPpR4pUKd5Sw/CHQQlT3IQHCNmX4Otn9muqMoL
mK64wdDxq0wZicsaB1b01TDRfGncXSMMZLuJltQFNbO6b3rdNyFVHM9CQERp
5FH0A0DWkKxxdMg1Ur+CI28nEzqRRrxCy3k2+iT+wVGvT1q3VaDcJLDqWxF+
TfxN6h1eKNMJAwDubebW0ZrbVP+c+IS7FMqFtqDEV1bb3k3Qx2T5oi7PHwan
v+LQik5ogDCB7B/B0nHIkV+LAwwB97qKbP++Zfv7eo8AbbuVY1yuDFbG+/b6
Nyvc2uDfE0y5O+jZwc1sIU21cPLVHxpXwiseQjKcDrJa+kJThU9H6YwcYqbe
3XqnVVE8LJuo0cLbsjzshRmMcdvDPTICyQ4JEcl6BVL1K2U+HbLV12mHxvEW
ezxBI4HpDB2gI1o2IfCPmEhkNcsaUrwwThVJNW3yR0odzRF7jnqFTiwYQRPD
OHNa5hhHJZHKwOoKgktUsYdJsRbjBg6GgVQnPSWeGLmyPiTGGemuHN90t1w0
Hk8TDc3IcoIHJy0MOPwANguPdSgSiswb1M+1AlU0JCcb8E7NarvG0ipQKKMm
MBn3GIGwNgjUJOS99bq7cRduKybkV1asEjdOxJhqFSkHdWtahHPgjL4D1gFF
9vr/VxE9HY9J/hSb73YLYjxSWpjmm0OLo3URvfqNC7DLRq/fRwjUtFf4R4xv
4Zrd714Bm8JWL64f5D2w2UCfTYIcV4u2p1sNJ3kgTZU+19i+zl+orkz//aOU
ouHEnkPqJ9ZkW3P9k/j2TxOgSf8C4qnM2SKJitpzOW1Bk15hMhZ7NKvKy6yQ
Gqw7ARGyRmxukn9suIweSRkHPYKWQLnrJDE2mVbpz9dpoSouY+g+8nAoH9cN
jknoHtfkQOskI+krfBE1rVpx03ohYg0B1AWlidiqSp1eIYGtllvxA+F5m0Cb
+QS4FlMHXBx8EopTSdNqo+HTNph2jsR4htG2k/Du4iFiQw8ZHYOAd2R/FUCr
MNCR7P9HwZJdWBuB9dWTZO7U+rrA7KqksKyksaQfrsl6TefIcxZ7tipwj0iJ
2BdtXJNzaZ278YVkdiW25arAD3fWZLbIrmNqFvBNLOwUDiLT9dGKgcZi9BSy
vKGX24nb3byX1VCOGMbaqlHasPv+gwWUzA2PXXhCTkZTr1cYuegWPjAZbWm9
9xMOzK049qbaDtnPoJMaiN2pExMkox6igBAxwItSkpffXP/PcJ/yXcytPQ6X
OSBpXXix6SUIn6JJKggk7UvLcG4x3IthUIiZW3mwmI9TBedXldhgjOnOhi7B
pTmsAzeY7C7QopfCYoOJ2Wv8YaIouBByWOur3RWHRsu0VqoLNutcMt0H6HGG
HI90nosI00iBHZCqDzm9q2GpcZLAFGC55D4gT/e16bIuhF/M51l1BpS8JXSG
eMz34Ogwnz3Hzpkcys4iWVvPdDeCuGbs6lFZ0tpvZ91iDwfdFD0JreZ42+8t
AJkcfr2pv2jlednRQDE/T2le93DlLviVqQUuJ8X6zZfWO5dkWQrt6N3UlB+6
WfzPbppByhS2XVdhColRwq8Q9H0YyD+RVioRamtspPocJNGomQHNqMiMfDKS
xj0ZAsIKmx2TIL2J0CKW42H9JE7XKcsPFuf/FRUhFLZ5bLRirXBmE2y00yb+
BB9bRYNwkDz9epg9JymehknjKIEGxZx097EM2FKTaZ9h21EBjWUetVzSiuLE
+U2XAZSgCukEBG7X2UDsFbSPmnM8AXCzdI3EPNgNZBm6p/RYzVBf3mcYuVx8
GlibHDV7TVCAhH95vI+ECMKhutYdy6G17U/vo/VULkTRBvlfcC8JPOlGLC/j
tQJbJh+fAoMg0WxoPGfNIfYANF0RtukS6XbNKuLM2hcxDjsCrb2ue+UpLDdR
wDZAFAbAtnH/Js6F2zs+TvGeN3R4kWa2gLALKLv23Nmz3oEffpZ3aIbqRUdC
xB/4I3DOyCB4zy5uRseHorx897gJ6Y7RW3kUS5cPI/gYvbaR99F7tynpyZ2R
fCjUPEp/cAop/bXpB6BKl3hF7Fv2vr2eUz9Y+/NPKe/fP7+6NO5aXE32fs4m
xrvkm4WE2cpB6YB5d4vNPTbccwwq/F5eakL4GOHaaP11f9y9VSeCHuLMKLnR
a8uWnW6wsFayV5WsZztPP5xxFZzktkBsJ+daFGAOaSxZL8maMVDNXPofehrG
apvFyuLKAMJxOPznO6cO5JbmUcHiHItY3r+PRGOngZmiZjlGmNrzYYO9UUOe
6HLx4MaB6XKo3p2EHmogw99q66GlKHel/sN10escM0Mw+GL+g36+y1eyTsrF
zakann4oAvU2fUOdZcrP9+DUH1+PkMgdLLUQFjwVe1Q9J46+VqU/f+Ur0a9i
QkgMJBVn1eJW5/lLK7v0q49CtRrx0nmlS52cx+Cj+D70iJeUXjz0Fb1FR56a
9tfMUeFWTTbEkzuszEnYI6tKvxyWIH9xhNc/5HhreNhYpE7lbuM4aK78i6Oa
/Q2wclHLnLhbypAYgGfeeNjFZDrpyOvbEzvsJ5DB5pzJB3axnIe1jSLHAgVE
gl43g4qZuWaaRmZH/m/CkLW5Rq0fKUdfCuhGKZYttMC+RiuZCi5omQHt77HE
Pb7uSRD0moNBkiL677CiuleUPHoQfs9fm25CntQZRgJ9FmywaXisVT2bsCwZ
K0THAJL/NvvqrbbH5BPbfcx2+UvQGMg/2Vla098fyviFMxMKEhm495+By5ay
Ew+CnhFYH8mGAHYtsEFSAbEweDPbsI1Vr908tkQ9I7eoCScREFbiPrJZZNEW
EYXibJ3MpuYB8XJAdhVR6CMGcd/SFUh9KQAY9kddGW+TaIayGwuNyCxh/2Kx
/OrTEhJRQ2LjpVgdTSvoBblGA4VxOqOwVdLIrYySYU/SG6sYq60yWmcmQoh0
GkcN4vU662pm3cdPeoIKcsrTaAhrCGspkFVjOHQkNzWX1v2BzlK1ehyaIYLq
I+NVaYX563O896d0w1ZUFDOisZA1G/zo42Apf8rL5WyUsSQKIyOEcEILGl1I
+e8q8zM5FKNAC6m5V/U+6tFaxWdZEek7MDahc+rayY4m/QLjfG4UxyAAFEw1
oxPhOhb0nx/FcOivR48aUmYPuR708MfRy3BFQ4WPfgSTKw4WkxKB7BknipjJ
Y9QS9BSoMoUKnhz9o5hYmcDUsmu2cipuKyZgF7jXmTBcRFnm8DuJjhEdFJEi
OxUvL3uZdqE2MULz8JdyT6LXl7pA7JGyrnlDyeAWlL0UQd1j0+cgdgwVm7L9
snE4fy78MSEO4HlviS60f7amaLuM1Wq+R9d4/b4B4iDNU0r8LDH71mNe4/IU
Qc6/0TY47kXnl23n7558pZR5P2GJX7xn5LzzlAYRW3oGdsiUaBXAmkxRZtGO
XUrGSncawXTMXXzO2ECLuPbRrusFoW+Lr+QdTBLaRl8G+Ai6yoxCtg7Jr++4
NLxrXdVE4IVJd98PO1z1BWmuIEX8Laakfo/3qXGWlFdbhK2SHDgcEIBf5cxs
M8slTN6b290jRoTi0XrOb31dmiXkr+HOpBsTBLwTLVlA/WrtC6iX6ulJ+Dr8
7jHS/KdYVf5dd8jy6p5m3BlpFTeO3oxTKOcHgWZq3sP9lTVCm1dSIQnTksqp
9Zvx33c5fHBwboaLHmn+vOLRwNjugFPtVUg+yE2QG1K9+02nDxfmLHCU55Kb
GfeuQ1VrnE7r5DgVQq9in/mmSQvIbv3gWFiASAO0PKo/TdSv3HTs96wF4/2N
FeKAUch26RjAFphErxLpf7u4ZU+uRZA/bB7uTFP+egqGRJtnpZeYX3pQYuw1
eT5jrrm29XObFZd9dpOe73meOq6N9/3as4mCRVMhxcT1mCamBaFJdIVLq+9c
N3BpwkC0NZxX5CIu2wencgqdk40uYfMvnvl6dw8CBMCGz1kKWg8buVNGjINw
3tCEMCY/16w/nXPIyGM71j7rT383Q0dGhTECnckfu3f/BPVpzWq1NJ53AYor
Hn5QDa2y/h6D88EOgfi/IBim0xUFWCRMWsjwtYw9f8zW8PRzJObZh1V/CmAo
qCXkeYNu/zuFDwhz9xtFBn1Rc5aZfj8wdLL6LNTwSwMl0wU+V075NTD2EUK/
ivZx5inMVPnBfxnQPLchJqCWYGw3DpQZjW0LCdGOYEve2vKr2Fn9fXWSsAOH
8RxRbsWVgx/1B2ssYuK/Bq2xw8CDD9JSDo8XMoXVcP16JdeDXBdqT6+BvMIS
x7DyvB4Iwg+De3R6h7DaQ5Yq0zI0/BQlFT6E7I+soVj4icMiE2xrolxwFgNa
rcDNx8In6pg48l4e6jbmWr9G4jGpLQwYF0EPYKAkU7AXb9Ct71+4zaDMt3mz
y5ETGovJs2hzAtpUcWX0rY/l+E2YJpIqHrnM52zHcxCJ+VJRX/k9IjTlbNn7
daavoAJfBFFFvSNqY1tyjvFP6es7OyCh0x/Lbu792lq65tz6cYG8SgP46GmR
THPkUd/KM6hvSWnuw6lGzf0u97rT7DG5Ka7pJto6BZ8J0y3B2QYd+gW4q+61
gWDXyXqSp99LaS7jIqQHCFZ5Kf3QVoDOeJPRiMI8bczNI5ccz3eUTXNtpskJ
mDHDazr+R9eoc91hioVSKeBL6yZdvaRtnbDI/AMtSzk7MOu4IiqJ6XnUXwC0
EaUB96EQmAciPoki0bDPuDNyFtHSiAKMm5e0tACxpuWXjeHm1LaxMn4WU3zp
T3ANmghH9tgtLf9KHRJjOP4M3JN6VI+bu6lUN+IurK7Nz9JYP39zHPduGrWx
cmOAc/FCkUJUr2ne7x94F2pG4qeY9/Eyg+1OM1IpEpf1+de/1qnILCsUh/By
peZ1kDfsRZSeDCY7CVfPnREp2Px0rBz2euJTPTb3AmgLSEdCqFq4ACAgEtOp
FdUvh7afiF0RuyugdsgNhM6ZbnkhP+PJdau5WuyOzCJaRWjAcqbbsM8ekXPq
3dRqvQUzT43oBOYahgzEt7txqAzcvDiykoPfQK+2MLGZ0NR1MAx3J03shYoh
OnL1AW72aRVBDKUEHnRPzghCELwrDh+ZLDm+NtHZayWRD7f9Cf/531nb1e80
GckS1iYu1gMsC++bqmZ3v5qmKFTsIzjTd1JrhMsT7AuLmEpd72l4bcAhpXVG
uBWgx27m6o+mzadmp08ccCQzl3SRTMdkl9r0zkh9cJqee8KCA5CutvXuGiD/
sV8IodlRIBA9AoGIBb7rGhivf3j8jEDgvqx2KT9y/20Dih6TNlMNnrOyZR+J
qxbAssaNWJ5fnhCEL+CuvDWJ8l3G1K+t2LuuWRH2z/BS+MCbTpKnHvurz6QK
ThkAcOdPbcldv1w8N5XG0zNRl8bmKmPaoitZ+VGiLST3xCaVOSN951kivJOS
XPgqtUitRdapqXD82jAXhh6jY8E3EbNCLGJFXP1E9eHhhtUMHZw0KhF8EISh
mzsqPt6XcJS6YPBTmU+ioc1iLFtTWqNQhfkwHGU83hz62EgjedQ1SLC4zDTO
sVbkAL9A5N2GMtp1qtFh469rXCyfApoSd4pkqTyHk/WZL8lgtLze3ShcTT2W
BZ4zEbw0u1uiajz20nhC0jA+4qvnFBUEd2DdNMMSq0q1ntQ2U7aNR1bgVEyG
ncwnM5FQlJo4MCZ5B0tK7T2yOJ2j9/OxbtIjKG7NywrTnlq1AsZFOdJzE2+Z
9ACkOV5rSPjhZlwqvVLxgg7a2KqePPa6TONpGbDI48TO3LPffiDL/0orwueO
MHg7v1ZyahRkg8ZyTwGICeVtxjzvq8XAlC6Y6noj7s9PZ7Z+AfmiDDLJ3rXK
2AbArKgi+PgJHCbY8/std+z6KF30VIUDKkMQisV0GJ66B6/Qoj7ZEXFyQ4Tt
71O9tgIShjkfLqJv6h/dD4kjAfbV28vxAM+8w5NlaPz1Gd/o6gcaVOBd2EgO
fY+jOhYw+yxSRkjZoO5u609BfsWTpdsUjIFQxMy1n8T78DKYkrBpUW0lyeNr
UBvwgGWE7mfYvbeJwHuzeRJfbnaWbJpzXWqKbeqdrX/f9F/touIGFpKyzEBY
Rz5V3r3Ux3Ac/37OPGHYtBo5HVJ0CohhL1h0tbT9vAIYY0b/lK2mbA4fPQ7v
CYhKvtxzJHb6UKYWZEMT21N6f0tIrSCr5pf8Dn9j2DCfIWLyHlsNsGUd41Mi
HMmECJQe0fcfeWvQ3MQ34GPw31DHF2aktzyWszmDtw41qz2opPQ5HcejR5X/
vQxnrpWVJvTlGpKKTi8kzEvMKezzxJwVsG1OAtdWtvMI8PMKAeKwTjZx/82J
Q3/SOkjSADbTNJwYEISx/tP/ZF48/RI7EGyFOebX8V+zb7QRwABU0SA2daZD
3Og17KQLQuj4kK87n5hsNlml/P0cgoGe69kdKY7h20cuFoOccfEqJx/8UfM+
AUqsTxKbXo8Uvw1ZuXO+7hfNopyHIL/Szrj38eanqnHEOoa+FyygAKqRnmn3
aZD/ETOBfk2AdLAUNDtTJ/gbjlbZWZI134PcMY3QGiVj3DlEmZrHLYVn/8n8
fImh9mFRCAm3O876Kl36h4Kbn9LNHlL1+090xIOZP7+IVwWqZoNZP0xeflcO
e3GNUFRga7boh7LOltsAnm6zYyQkYiFkKQv2gcevxHj6GcuVYnlyFCPX3jFb
h0v6mYbe7I9pIswS9+Lw9pZYpOjMwliZAyHhBjXYIi0Ud46A/K1N+vGEv1Vi
0/GgRTWqag9VOA4FEp27LjSEWYk2sSAjpHeelBelgT1DhWzeqXUdcPrPRkqp
B4QwsDqdSnWrZexviESrlL6RJSbHDmCVoH51wlELI0KjusDamwLL+823mv5v
qksImgUSZH8WnQHrEMaPJN8F4drmzWsQ3Z+103188IwX9wnuefrNSZhQeL31
JWcrz7h+S/ql8y7SxOh4+GGOZhjWHk55jLVXm8DdtaEYda3IGRUQsLT0BwqF
duBt5yX3rtoDnuo7EpjWTeoyhxB+FRDuOt/y/TYJzhMmZOhM2ycaIFQbyZnA
DJk4CQsvaUl473oRzPJ+0aL1NOx10e8PZ9sb1NjlotJWb/5wgP4CPkvwNlHV
YEtcliaSj67W7hFn9yBkMnArPr/bpJ8P6cltX+EFCkMgPDb96eXN5R1u4Z7D
Dk6KtGcZgxrTJgANgIevrPnQG6qlyLYvgLhE7EAfcL1/d5pN1rIXjui2lO6m
CdLzk8LHxN83VNl4cGVxl8UpVdn+vCtgvm//HM4N9mn7i9RrAVhCJI0YVfTm
hcjbiGJOp9cMkC3CYcYpSHwgE7jrCKbvRG8zXfBtFg8eQGzwKmykMAK7+UqN
/kPv/L4iW+1KNwjv35sJMbzcru2l57ov6UmyaD5OZd+cgTHPAyIHu/zeqBmX
KIAacm8ksUQrePxyiraY957iu2SgyPnVH2Ks3UMWY9djOd9dgHiWVRS8Aeix
EAMBCZCpS/Ot7Vku1hKg754Y3xqgYbvm47WkdJkYWJYduSXUWpIOcxqzpNcW
sR04dAHB5W+3lRMw1MoOJMbuM3lK6gvbFGnoUv1Q8/o9uf/uAQFl8BbbNYEy
bXADwSBMU/mNQDcdySP0EJWlbWYADHiPFCnG1eNLgOVd5a6hBqmG7YHeJvZl
JKBarLHqG+yhUoFXMNiTS/+rS6dvzY8GtW8pA2iZWELNFQl+mA2e8z4Lb9AW
5ULuU0ujtvSsptZgfJVZIX8TZVqQt7gX8bG546FdZ0GjP3BoM9djRxhXKfII
IkpLx4mPQ9kqE5bIHJPQ2epQcWj+n05bgHVmE26gXU7zxK1S18kWHdo5lYJo
1ld0KQYVTWGUE6Ww+VuUAybljghATQdAe81VYu0NpX3EViI4Um5aRnjCnwZ7
8ziM4hWt1pWs0igILg+kWflUIVrV0LHRtfOBRlrjFGsDS0DWVE71toU0+Pxg
Mc883XZrZH6guLp0FXlUkM8TwUN/TwV2+GoZaIDe8wEe7L6ZrSkhCMHgqPeO
mT78G6a+J3jzRPy8OTk2HGQ4EzgSk+XtHQp9ayObHA4l3W59FrBWFVclP2Re
iKYToC1sA9fK51zfPz1Y3YkHO9zHGaEgx91VyXQpLTYZN+IoqHGC5h913Xz9
Mv7tuvQTjmEX5K22V4E9OGegDpehr3yv7L9LG35QjW6XYzbdG/Vpc+InX7HE
BahyFbHEQqxoBT/l6mKrTxEmMwKlhGVN+nTzlfHNQh4LY0Xt8Cd0FW+LVirC
/YMH38Rc/2wEp23kUtJ+dSkeFcRbLe9nY5bzMgbKft4hQw2GMfGtwxU+vgRD
5w/A5GSfpdVbnn09F/iMjvUuRzUpjYfSBqp5FBeShXOUndRhZAvEjHvOT66R
gE/Meld6AmRchSmVMU4TAliJZdcCljk2wn/qcra1c+wsLn6pdKp6kXmoXuPh
h1AwUbS0fcanWqmhtJ0HoWcLpog/zNYPxHNU6cCAqVU4O6j4UiavnwOMeNcK
ra2Ml2ulDa8pGvg4mNuF9t//N016hpYoAZFFX6GBKGlVOpuOyY2I2Af4EyU6
Kag8negrQR4f+zBJigvFCoU6G53c0RMAVHQhBJrnFbEVUE+445IqXB5l+zZe
x815tzaubpsFiJfVNCdsNYmwXBjWbHcXyi5J4MXZLmEfcyFxdOOv66xAx7QB
40rPrjtcjY7zs6ldnP6Y1Rbk5DlD3vTN6lewuqc+2r/Dz5kuVv4aLqj2yzMn
uESYDmvP2/nga8s2ToO06SetYsZIQTm9ZtA2b0c3kWowNd9YXE/osLK+fsJp
IKe1A4+rNErTFlbaTDO1KrPpH+SkcX3/5ESdh71Q99/tECXm9+9DzSgumbTj
dEfjQTugqtK416OYg3Pf5QC5ok0oIJ2HSSoV8hf9kUox4lGeYY0QEZngyuXL
Q5kyMdMdLvYBm5FC+OJ+YQGUUlZt9uzF0bb9bZy9QcOo7dfemPktpTpMZN1r
/dAz/EMLKeNipg/HgRliMdU4XGgAhhwJpr8NEL1GIFCmV+hwe/JOiDL7IKH+
il7Lo6KIV37fP6VgvGkUX38waGSDM//i/a+vJBFs6DcTfpnrcAvv8BYkOpjs
Gk0NjRoiPCtMFrp2YyDXW+XP/Wgc+eU6Pk8DqdywxiGi3MBsR8LAO7tOG8Uq
Zzi1M2u/0sjhTakzGq1FvbNszaLPDPOXwgPskTVGA9GcjR06tc/rxAS6KD2S
JEli15jRHYRMyVr4dG3sZk6Aqup44zplxZ0BwfypwwP7mDSZeTD6TcBeoOyD
vVHbvtodh64SqmKkrOnrtY0Ltg5+Nsmq4zKHAHh2WoOaCwlkHbNm9kwFVED2
ZT7jCBtUZ9Xa9T05+ZG7azHCHqMQmNWecfiwP2DV76p+CaR6b55DogwiXlKL
PKJFbuLbAJDMJoFOV6wTY9Pt/FNHhulzcvy6JyB19ad+EGreWt+Ws2TE6M4e
jEzUZLnbs34c9U1JJB8ElbDoZ4wCLKw4yWTfMI8zdxTQ3NVHklKS53xjKYQk
Kbs+DrsQmy7x0S+vlJ6FSwVEaq37kJDSxPeMg3cmvxnsD2PhWw49TMM/YpQo
LH8ubAHfyuo9XYahpc/0JI1hVEXVdNHFUG9KMphZYGBC+OZ+z78uWqsm2ymH
NNS7aknih26eaeF9xpMj75jiK19kCH6quflaaiqsP5J4dtV0amg/W5DCe/s2
ucv9bObLheQIZNthRlZCtEU1gZDNPcWRJGSCWd8mF7eecpxMVAcaR4pnjN2L
5wtaqUdzllgleMh6RJM7LzUGG+VTuPtyo4Scs1vxikozmBCG7cFDsHivF0Ts
QNOdz0kx9g0vb+OHnxXdck7A6OthQYIG/dCbtQhmGDSQXiokyA04wL+s6e7j
VnXXzSkQEm+KXXIMqXRYYDDDrV7yNkhebgZw4qhJg9zO7/vt6xrg71TRxPQo
r7PisGYkBPVIrm8+x6/amHI5YLSmPCfr2OqC+f0lfFNJc8O1cQcHnXFUxPnh
dzAlJEFPog++WUBBgGq/Zoqo5j4mQu8VPkkdegLgj9EkvNw7KOCIuF9sTAnP
Al9H8US7ZDxuzZaF7pV9wAFJrf2khWvcw9DqQqfRWXKbqg7Z5kuAgv/ovAeb
zrdHl3/Ge2/a0zf5bn6/7cb5YmoezrtxV78EyuuqGRevCapCg/GMcUxhctUC
qX9KL2GvEqqZy2MGMeUDBBk05EOM8BK0oHTeGG0NkroXu93NAJOurDus621u
cQXjr+hSxFNZzOVdzrp21h4+Bnj3WDB/eaQ/Rz8w7ySqdUwSjO5dDn3kV53X
MzsUalypmyxFZ8eQ+TtqJAYJt0qKfSPWrb8EeDSMNfXjydFdY77QNCNo3b5k
W3kQgeqaBgsVW+qdv8oOhF/MfDOd+jLfS8rqUCYZcXeKUYDk538t/FQlIW9n
XvF2y/LgSKinvcSEFA/9tsDwl1mNAoja95cCG/+3c35+anLc5PaPIv96SYgu
u1qyFn0DYPMnIrHM+rbWZ8YZNAiDs8WY0M1fOpLRicttiUiwnqCMs2ebw897
rPQGBcP0+2857JGffAha5GhOyLIGIVd+R/Hch7mmK1QxfFLhYYConmNPalYd
bGZ636nlKFpKjGHA7b3ewkv2phFF9YTLKqdcFODDPjWUCOLpsveaKgOPlC9t
b91Iq+hjEhhyUM7yvKpd/Whh74xj2jQuV6M+3yr1K3Me4N45qMbPkHY9C+Zw
U/PRHKmkMmQoxWVx+puTtyBpauWK0OblB1wlKsWEL1l/jm3o8k7GlpV4T2Dd
17a2amwIQqJbYNmRLyTOegX0fmdfGsdGJU1vRFucHqduzV5lFmvPS8Rzls99
mHzDSC511Qmq+ziiHSvyS53wWxLmaO3hSR4dH3a4YFIJfeciqG7xqzdCxT8s
zC5mGUuVl5wSc7HGtn4vmIHzQ+Ls363Zap0wfbegW+QslRnBbrHixofwm7F8
vWzu275MOiqUOYMVVPLy3e6Fe37HqDMwvoEE4kr8VV04RpqVtfZUBLYKTMvB
6+hbdzT50mFVchUl7KigeAuqSHRM8RmBFPU9tyBGrdzGAiR5H+RwsGgKjqEX
fFxKGKUvDfpUJAkkjTazUGEgT9eW4RVtqQUm95WdPJaqpasEmSgB9e5tUjww
n1Kd8phWYgfGFye4MjL4FfVDNihrgNFyfxXGtc50jc6pKwR28zkZazJGLAhO
zTimGXfbubAGHitoiOjunX5rkUwaV2A5XX+XeTpoIGoJQ4p/TOMIVMUUXmR1
I5K8TczfkE0q4xM5Gq1q/H441FxFj2yfFdpN0kb/zHmZstItKn8z/Vwtpm7p
EeC/sOdo4zDdPtLTcrDz6kAUIFDv/fMxfmZs6FM6XHIkFQ46B1okBlbaSmV+
ZO7SBNxk24nQOPwTEGKrhMZZAqMkDwXA5tNfvNCMO237j3d44oEc7i1uz+9C
ejyEpcMunAvFWINSP64QB3+J+1Du7nMB0eD9ZkH4noId6C2jqaFsWBYiG6bQ
WYsWQKjFJofoqsZ8YagldoYt1A4ugb5sh2nempiyOi1CVP6iFU82ircbYQY3
E5BCMb/cHq2q3681qBw+Ubd/Fe6Y/0wq+L1NOpQcRY07noSjn/59DJ25ur3d
uBZjAUtkVoD2aS0Po4jZIjbepVkAnINKjafKObx9m2YwE/zzD5M6xaLmm2GY
uMhiWsCkL5qZW4+G0Isp+IQ+pMh05ZRDLP9UylZWsg/OABRjJjgpCVBbNuIb
LTQxZGoo1l0z9oHUTmESkBorV8E481xmlET1hMFjTb9wOp2mDvQ196rXIlkM
Hxlwtl/3cln2eDWFTdHqxPxkFem/iNICY6LpZuVyGrEkrOmrQjqGSf1ItdEY
aUOtcYyYDg9E/wGT4H0TFPWYskIOKI2sNbFKKYRxHloh+PdYH2sDvuhppSW6
5+NBAP5xQ74md3IdhkIgcgooglOqn6NkI8vunZTI+yxRQLQVKOmD1+xd91IC
5BAKDu4j/z48uHHHymqw+JMRrZW58ZROM/TL8V9oU7jV5UJT+3OaQSMiix0/
fAsXOwqqEPBD+bHd2AfjumQui4zOYNYDWscTpbshwmao/w5dBNe8zbddvVi4
IrWn9LxwFDg3ihUO1kXNSIn3xLTLSdWl4UM/Z7W/qjsEZt8vESZR9+o+EJEQ
qZFOHNxmnPDJJ5O14ZrzFtA+J2ndDJ1bSttC6+YrMoU5hHDK7n3GSyPGajKl
TN5h4gYrG4Xyg0EfvUiTJ3L5rYQ/MZPS9gk/UDFwXwY8ksuGeDSh7tcjcL1s
240gGhUIf5cpkcVF9ayj6CXfXMqoP1Nk5RSwu7S95e4K2RR6yxdljDh3IfrY
8i//J7YJlUYAwMwdrMBVOXzdeuno/5K9hkfHI4t3VWg+TcgzZGMKPoI/0M9P
3LN2iSk/Rv+REKP2EW08yUM24wqmCcCSJ4MFjuX9ZEMMOE22NoBbteRUYe7u
hXwZgtge8RnrRDcgwUj1jNqFvmBjOCR2gTO1FyuNS4f4Q7uSzpQkEejNvUy4
0Dia5hmdnVcMkthMVK9WeBUE6pSUrpLIvohlLEWLw5lT0GjMK5EN+w9k6Ek/
nfuoMPARjzPafE3H2DJ/nabYUsQsDH5WoOGzyd/jxa2JAkApwHdSvEO0CelY
GEj6EO/cKaD0W8SIh5uTscZnt/xMoSqbKwTHkR5Hp+/L+kEz9KKw7dEqIK3d
UuzXmmU8L8iGkQKUrU/LZku0YLt5ob1FrvgW/dqiR1RsDpCf9gducDcKk5Ne
HBgl851gsp9+UI1NE40Osm7+gpmBhgFos1wicoUfKtYE4e/EhIubhr9GMccP
8iRBYzaVAbdiT59DdoANuWSNruYS83tEvA0LI7Yt/tgG4xqChSoqmN5s/S4M
nkVryRc93j3J56upbK6ensoRBCcpvzePl90u8oOTPw7U/O5abDgf3/CfQw2O
A7zNYS+4v2USZLFYOrVxiUE1srnYrwFbYZq3HZNp9/ujxoCxcB2LRHVABNdU
VFw0v43A1B1yLlVh4OaA3pqbHjheIWfr+629jDGE4FLQKJe5ZNhoRPdV3NV7
Ji3ovjQLtT8xBYM/pzKS0NIMLEXp+gqhdSQcsnDrtI4rqhSnyyUUceYGRpmR
BfxbhBlEC6GIu8n+um0MJ+TAnlKIIBJpbgw9RJadzFvZ6HZ1a+KnXMPmffSQ
bYsaIE+E0iHggW9UqfBRbwm0kKmgIjZAXj6XFeCSaULS728eKTtOObfhR1To
HNqqU7Gg62603KYWX3IM+cb4wHsEb3IQ5njqdS6Z5M2Q/BOxexPm2KM7LAm0
XiEUeB7lReFSyyWRDA9kmiZK+7algni9p7Qs3gBtu0Hg4SxW//KSt6tK1ThM
ow+PKUvDJhTG34zSLr+cjpZLYeYH+GO3hEserK6yBRQ+0Q/VnBEYFHBGX3+3
2+rH2hT0dD/1ZOjEKslI1CTldzQ3uBCoCV+S/+Uwq4s2HaTXLsTTFs1xXNnP
jq7M3NEjf6nftJizuUL5MFo2c50NNYDPrPSe7vvdyNdAFKvIt0TcbazroeYf
m3bvPFLUpj+ZoPZlfC1tl1YpfayLLuHETSwarIunbwqNYzJ/pkDksHqgGHws
ka1O9IE1NKXlQwbcVFOufQz+by5l20zVj/zSY3zoHlm/fYWqfpAkr2RiNKTk
VUUvggaFup/5kUDEusBfxcm46QV1P4wiQD8PCAlJlBGK8Sq51K/9hBhccdDk
JqhARKE+djwEsqmlBYMBC3nIehjJroK8GiFigfhnU2EWRU4hz8ioXmdyp/07
Jch+hKVQar65W6EmlyOiyQkNaK5IR6ap7RtVbANx/LXN2uIYYxq+pioqvd/v
qPHHnpw3b0oRyjRKH0VkWUQsr+/jr8D91/3I/IcyrWPp6C4yY2g8u3DSvlnK
NJ3/wKrRFw2GgHa6ytCMgQw4hvahoVKGhKtdAavqFJ5O7UvvbWTqp+z+BpHI
2alJpwA1oe62ai86EH04kKUdDrbBG1ldlcq1n2zc0/C1+8l0lAfkAWwK0/U5
fqDA5EyDY/Ps4XasgjTiqIZOVfUlr9qISkDlyvlAF0ZzZ65D0nZjP6wFrrYZ
3P+qnK0toh2Adaum/yUD0fdrgX97e2ATALgPIregliLPVmHS6WxZNPzcn2EE
4bWues9oiHuEzt+y73QYEZ2oNWzwF3T+GbHSG2Ngt7H/Y5qXyx7S8taJ+q5E
T/o91iydBYXtaPXDqKANXc9u0XCjNf6cTwlxKC76yPzpbJ2SqKpzYFtqO0KS
I2BGUdObUaj+4+X9mB4PMXUUe9FqtfsMtStQx9f9eN2JmPeEEnxX20uzuvOv
TllJPZ2ts5SipURc0jonZjyTqO/mfsqd9gAKoPyp7MRwoCNFrm1MZTdLlcJ8
Yfyt5e9qYEYzmj4NRVMooww1onEnG2DOYDOIie+8IZoiLlj4VJuld9xfvwQn
neWeRUClU7Kpyqu7yr7uGVcqne2KX9M3nUlVRlVAmmcsK9zWBbfVUsspAYGj
nZzK9jO/iFyenkFybwlG/GixOqCO69A+DPc3zcPA3BJ4AWzHxluu3JwdOO2C
IK3KX69VYdpMzItoKCXQ/QBKqjH9wqj1pLZLA2HNINSrEdD6TXBLuYT6jvBs
8jKIlni0A99yY8Qsmu1pcOVYunT3BB6w2s0vk4nHD8njS2QaQbpIS8xbt4Fa
nAlTkmfsG+kkLH/C9haSyurJKaa3MeWw9k3Fb4NBNn8dr/dbzaI4XPDqsPl1
QDLjAlQsiqd5ZzOZ/V47s73db2c0akrS3McV3v3dwckgFAVSRhMtnYn9IEIL
57gGVvAh+0ByQE56roRL8LlaAgJm/9a77AgxQyOpm86cvwWatP1HCCHqzHnR
IB3u61R0Egg1/DCZEvX1mrvwJHmwsEUl+pvsDRnOsNFQGxJpdaX3UMGHTOAN
dpPHuEtcegUA/MSOkY30xQo2alei8mP8H50TSu3G6ewq2c3X94DN+PiTMTz3
LKIQidOnLh4u6eTRG8/SCFybYYAA/BzditaDoxEcM2gHKhDWN8HSYBmVz8VQ
7DtY2NygJzLF9ySkkAybvbTI3xr4TAgD3JNwRwB/LQ+7nsvL6qS+0wJWQZlX
IqDuG1imlVjOCFUQNG/1BtLxrnvvRmQzGq/SENiIUrNXNHE16sAk8hPRy4RF
eTmDEyBGgsUCct9FWwI65QPJB/i3qus+3b/+Y/DDGtVbuTO/RL4g4Sp/W7BR
OFvrn7RURakbrwlsGZsroPeWO7oScZwoB0XEa7mosh/t1AD8uUiVChL8TGZ9
nKkPLDtLiK3/hC0SipGQFno6mDPw3QYjiUmeRBfnkWCAARnhoKMmrx/ECQMK
gIGEVt+JRuELQBgQ2GtyE3q3GksJwPWEAMO4bUujC4XLInTaM44BFnjG/S7y
DpsGAbs88hugOOVnI5oSw1Yy/XoWTMpRZOxCHstf6JK5C3VYQs8ooscWIdHC
ilvFngJXFVe7nPQKGzxOYyDY+UBsbt4+Ys7dj4LD9MUZ4TW/2nl3y46oPr+0
z/iVpC+H5yso7p76d0tPnkFhAiln7J+iA3kMc1h9kz7jgcHQ0bTU0XRpOl+7
eEhRTMxUQrK4SNHtN/SifZddpadkeCywucn/Cw9QZvLuJja6iixS7VtftI+5
BCToz6SW1vgS+eO1OSeBgFWjt0fp3a03cifVfWEjSa7ESLZPbiGYBt+C1P0p
4ixLXx07TBlBRCIDH7pEV/pO/KdcqMRVPdo0NOm7vmmpSaZ8qLk1uDOe2wJl
SPTiA4HF2PG1ItbvzuNORU2Ms6sQoeXin5KsfXX9iv4cyCYN1ChRxg8RAxMX
CXCA5fBUW0hsTQ95ht+prafntQwOr/n2rdYPEUKyhXAf/kAtFZF7V/M/OSbp
67OuB5Fl1bpM2ynNUlvsVYRUo98vLrLpDnB74rrFU0hhSfxk9I3aWEcoCl4E
L21FAAIaEnZbIwqKQ7wMk2ZjKkyC3vSiswV/R0uth7C/AKgW1iaxVIIOlRQ+
GOSg2GnM9sz8mWrfBCs4YJ0c0YApr3nQLE0dlKpUfdXWscGclAZCM5Xhwysu
BbGvD3hJUZVtdi77z6xdr8cTJKVwSIdYD0pV/YB8GZbHBzx9IOllAq2g08s7
0Qdh1NM0PDsJhjcFHyzlqwIIty+kM8WdpoZjjjHXqsMqsvZTZdEWcs4hOe1Y
s9QNMZ1tc4GR8S80k0wbyE3AUqxJChwq/DmOuIcWQaSPxEo7mzRMDVDyKGlE
rmk/hqZkEdx5RoF9uji4UDMzJVAG8dLC/jogZvu77baff4vae53l0XsP2ayD
J43TePqCk5zYyt7lDA3iVgMDLoCljpSZJfNRd0/NKbVKyNXOfpu5K0p1/1FB
TmbO+UfZcRfuH5P0v2dODRbaWFPaA6UyohEuwmimmc1szei6DUSZ0mSkR4qM
xaDP/zxh/QeD79B6NRJkG/gYGkRE8kuxA3YfqxFRAI+QiTkgU4/E5au73591
zlJ1S7ZssWCAzmsBALd8J8aj87iTffQBvTeqSMb0CXNmuGaVoO1hzzl1I631
OCmoKi7JFdvS+w2ndaVVV6CwOm0FMAi0FTkrKBSEnkpvZEkgE2p97LakatcL
xjTGUF69SeoCnnLDfhFf57uA6bp8fjkgSwQou85w7lPOQYMLOIRZBIe2zJuo
BuAQRFZcTmXBRYBl5a6MIpT1zZZ60JP3sQvdGSKW2yncKuhNXMGECObHl1m0
+CNfUp4Bra4chtsYExaZSlv6/Rw3zB++ECe9d2Pu9u/RDuPlwKTHBClwoqZE
cwFSJoLXcUrNkBzOjJHv9vFVFn3mu9VPbM+TrWfWKf0dtjSJB/BhEnutEfZ1
48ntsRXhpXxEmvr0/65eRz+b8K5OYSk3BRX93NjyIvzrPbJ+Z+tuXQxB9Ejd
uLc7CoEO4GHAuiagBFsr5tnN3TtsDXsJf5OjJt5CD9oJo4BXPHnE0ugu+eK3
V7oFpP3K+uSU19Zg7wGYSVBx7nIxoIYgarbGQM/7QkBXWwauINnFi3Zy6nOb
iYU6Zxoz6i/UFgGIFkN5N8qVT/YB5VFnQN2f9yFIpTPDsAtJWHL451QqNh35
I66MDJRw18YPvmH8/s8rPH2/QrrcSHxM6YhcQD4jKcw/56WovOrhzTgtIhy3
u9wbJIcnTdkGVZRYraXdJN1PRqIkOsSbcB4fu0n1saDIH+8jUTaUhIMQ6Lki
eCEh7P3weZ+YaZUG+TjBunuDwGK5n/aaZnQ2CBaZm4DmccDeS+rN2VSEWEAO
4K2YUgdRZHN5mdS4HYQDkHJo3EJezEyhSSusWT45uUxUcyVGdAbX4ez4wxmt
bnbW0RPO7GvtXnb2WU8d3OrZHfAVHXxVVm87FryJs4AA1Ym1WkXpjwAnGRCE
bDdAX4LVfutlWwP5pgqmh6x50N1NbFH0BIa9C93kqIrEOfFR6b0b+uesV9Ry
QtnsuqV0ORygXRUOYv6e9Sq9eEjUm9Rdf/8bzfHB7AFa0nBdRiRv4+qwqQVB
5GMKAmVhwO5BNROZ1fyVJMlUIq8O1rM7QRtNF/SgjJ6Xr9MjeHssBUdx5UcH
jeTz6mhIL/OIMfX5ajEr9up8qaOV87h3V06JC2oS7kwDG6FOtiAqizJQMTzh
bx8my0IrmmM6kBb3zd7tmuYN36qsjwSZcq1T/bOKbTTr71wK5y2GH52wbOwu
I1R41KjhJNqjwp21ScjUepxRoP68SHfV+K+Gh0hifX8HDNN2bV/gbhdo0tIT
6GJGHaoksUM+qMDJge71DwFv7I/V7LxdBCtZOexytE3JqSgXWYor4h0eZrpY
J4irZZCNBochAiOV7FNaARDSdm32Jwvxs38MT3jqyJRapSZjzeIrRsny9fbu
jBI9On9NwZiKjuJkO702+NdW+ov6O0U4yLIKF3mDJ7Gg22Zi+rcmMhE7GG+W
9Fb3T6OC9IdzTYkqia5j1s9BMyrd8sCnI1H2jpZrxxkYt7OhUmVy2CXwBix7
/TObJ9xCjc1xxLZLz38E2aD8yHyCdoUaIBaaYqFfzGbzuqCP9Wd62ozmlh0E
44qs1MWd400d/XJb4KVgWjgqQznucvWVtv8orGPre6A6BgfxxQb/67kVkS1d
JL+Cv05Q8HQhrMRKM5PoxAxiPSpOV+tUZDXpogByeEcg8nCMYiD9y11u92QQ
IBMcyGdq8dYwInmXSn7iQvDR15CMG24r40sOYlBjQAzeCPxV8dwUVMO2EREL
Po8+SUB8x8K/Bx+1+oCQF/M/NgMzW886VBptJKLR3VV0oPCX96Y/HejdD+vG
6Ke1kUL8EouEsF1Ig4KIjSMDERPzoper4Y5QU9j2Whtx1EefComPRKAAK/eJ
GdknuDVcRfa4oncJ8seBEPRh6zWrO31aaBXmrmdpbLFH4f+A8h4Bg7GYrlVb
jmwA2/NuzxO1pFHMSDluUdaYRFwje51YSzFwTE4nqmtplGw1vEcMUXQtjLyX
Yq6HgkqQkUSA2et5sH8C6hitxtCZWKf+yYOZ0Su+8mepzTrZlk3QfTpMVuew
V/60DnL9HykQ+gGd2XQjfb+u0uVV9BT5HdD98w15V0Tx9MBXpHO6xakpQlvJ
K2a/4GEdr3U9dERV7qP+zbvvUO/j2//mTyZRPkLzzDh28vvrcerZ7ZC/AKBL
YA54asdSv6R2A5G+OM4bY54yaR+sC4abwg97k3B/93agCFRl+gJPBxiOKFMp
HWmKNcfTXthgDb6eOytC+aeAxnw6Bd0Un2vLPUxNfmT01vsTkPL9eIFofCpH
XB/JzV6QdssJ6b+z3bgJ02ekeJTTMjljhg4t4BK/UtTSLYqpo9fMakjUaWrH
ZJ8v6uyTp1P+/leTmnD9VEgrl+cn/x4GMBsQK1f+/kDriSH0vvZdaoRA31Cj
l4fF19vJQgGxGg+cGXNw86aQKiiptwqhqNJzLyGOL5yUaQrOhmZT7+HBcvCM
k/uokuqOa/SwdJQhy5qkc5mIh91vEtsAdDbWCydOWKg/z7XSfkWSSuVGjbxH
V/Rx4/960b2Hq0GF6hx/94QGC87v4EEIHWV3zZg8SHladbAtxCAzhynT43IX
aLuJj03zdWe5mGMpn4d6WPRfRm6htm8pucTJ89uFMmhWVZRjDy5RIrQjcvGr
9R2lDdcxnkvil6jiJGKUtzGRk1pzqxMjf7QDLH4ex+i6bPsaDIZ0peLHeIkD
HAE7BGO31IqC0cBSbUDH37PffH/dJqp1ymZXSthqFouSZbxWEBnUFsBfVOVQ
yAlzpdPC5+xrM9BuWU1bws4YbrXYfI2Zs6DM7e2+TjTUalp2gtk/DFSYdUyi
E4fomNfhJJlRfqrIRKX66tH+WgYqJfa1A75NFlXRgaGPwxrdeB/LHj3VFU9a
iYRh/6Wg9xDBDncp7IrXYhDKeDBIxp+3F4CN41uHsDzvL5XfPZpqNS4O33wz
w1M3Ljq2E6AfBLPS6DPQhro0JTrR/2GpGskQW6mWwHO1qSMknFlJ9VNQmkUH
+YT4lKxs5qTNa53TRguVIj+qp3dPkl+Frlh1QNWpkHe28O3W3aHQrvifD3LX
6UUhHDLk/yMa+3bfsYbIUGQqoI9BuWq4JO04Yw7LOgpBqtCaswcS7l6uQBIo
rVhTS82h2tClNcOyP9xJyEJnxaYgsuoS57Y4FLFeyeSljQybH7ap1Zuv7+QQ
Jb3XQKQXMyGmnODoxENVyGAughfKBcIhvDRnWV7G7ZhH6LFyiwObwgJBwVYo
hXYYELgPz0TD1Zc+oyO8VK7KVd1UUC340zq04qFlIaFMvelFGGQGmhFKNx6l
ZGpfj6k8bsydDJ9SXpIiNAsWWuPOE/jq2S6AwnVc2ShGeP65h5vcVac8qlr/
6tk+03bBkv6cq7oGKdI1Xahyzc7K5xI9Rocw46Hi83OvFgm42sH3aI8eHxbn
FO1dsQ+19kUz3tkaz2ytRxv0skSPX11x9ju89xs7fgZNyhwvqxHYtSIUizcw
XI3XnO9EUZIbmxlcHkUC1+Uc6LgPe/Th4DGO0C9ly3xfjegx6Vnl0X4gRQnQ
Ltm5ZDT82/t2ZF8jfOYdqI79m07XrUixjlR5TBRVPVDfxxSO7ea5vuhPAqlU
p5y2Q0nKf7ZZFpVA12FcfDh47G31B2JM0N+AEB6i3fa7BHBihPmtX0SMrhVE
VMAJAz6j/VNRcpVMeWUHuLbE9C3t1Bn8p0vriglmzRuOOGvCo2kysQ40l5jm
FnvnBoO86q4L8QiMgg3hphok24jWa6evdGTNHIiNAeYH6VXtgq0vOMSZaM8f
qTnAovuHThrc+JP7pT/lQa1LHnNEcTnvxrwW6qVQvuWWZpG3UM/HkjAw+YPE
jwd0crLQxgNGG1XwwtpjvJTX8ZZTtAXwyFhbz1GJ0QQPcVjG8j1UPpWrMjV3
e0yxmxHUNRekCXrs+1kt7gJ/YPYo7B+hKKtV6uZW57Vs/3aAOI0qPoXmKNGH
b9OJ59yJQ4K4vx7Pa4sqZ47Ck2/LhTj8blgWojHIcP6jY/l5BtKf/sOeB7s9
+1fy8pUjRYJNUh+u7CRhn3CnkQuvrBgDHcj9EMDAMLJaJd7e0uJz68RC/f4n
kc8sSb7I/bWCyXylJ1im4UqMS8TXlDvOx1ULjp/CGXZmmsKLN+JmOR+irkIh
wl/1h+2WOYdd0sIXSbHkhLSBed9/wAtRku6+sHnZI7j08GEp2It0JO5/Jm9i
xpY2RXimCAWQqLPyiMIXvEqXQQk1OLS56vBLJp9H23MKLJNBqT7Jb9jO/s45
f+mco5C1d6MilnLeLjk6x6jOGT+GJtpTMSKnIqAKveF+0p3RvSsyOazpYYVo
TktjYW0/pCCFimfmEwdGacBLDZusWXYr0nf1a7F5LGxJkFhteRr0YXzO3ww/
nfmVrQYj+ea3+nFzME6SVpFXJAjpiT4M69rjuV7A6rUEj70B5sFHAWa6XLqk
ZRxl36xDaWLc1CCciOv1E/FvMKH6oh9Hy4ZG91j4juAhRiEOEl9Od5CxDJmK
TSMjBfyQf9jIdzxQhsUemaAt+4kqokFpXLHEyTJOENSigft5F6gCaOHRxvm+
XvLvhMp0v12kuUTgY4KLSmtAxA/ZoM8ARX9QBSiOYhPvfrGuh4a6LYJl67Be
Ps9Pl+8fbR/Lq66JGpYQvbUIO0betDCot5mnk4ifmAR3fzDxIX3Cm0Fvo9gi
nWVow6MPdOkF4Usa5wJ9HQks6V2zrWxxj0z0ChD6R0aww/dP4XbrHuAANGt5
E8Yg8JJ2XbeGtpD+4jqBDznwECEoGj4pn8xKLZ1pfqA4SF+Bxn4OTC/q627t
DkKMbldiU9GSST2bUZjxi5tYg1kkm1mpgUjFK7gt9VOk8tqhjJujkyXRGFDT
TeaDi5K0rHm7KuD7pIoq7juF0iHTlI/61wbTXh61c467Vq14Lwra9CN+zFzt
nvEAC+PMBI/GERdGonrK4xj4HY8lDad3FCDwmDMVkfXCYQ9rBqU2fgU5a3I+
s+8056BZy1HCaIawWQqToyLlsZfT+OCKkfTZ5bEz2gtloZ/5HAqc+OHAySGj
N7VUN+bhMH9jWIJ2I7QVFrx2WUCTsw5uLIURiNhQucPjj1g5AqZtYN9xAZx5
3o+sMi/XeECxJ3INicdJUEx+rFIrx4tXUux1EpHlhvIcvlERWCG1sUQ607L2
m9SRZUGNUizS8R3QuPOCp4T/vg+emLr2f3RZtzCGYZgIPV2RP9V7c5YNLqgn
HE5Favb0K4Lgx+8x3SVR/3pmPqX3ocK0RStFl7O4Nd2+svop8KkK7jYRyfF1
BgabGMqJEGsfnQ9ghNJNAcg+rOrUXymEt/as0y5TBpma9h22t51oWFvVRXsu
Wm79HN4AU4ky1EKxTSLqE7ag6Zr3kR7g8DDxlbwY7hV1ojFuk5UjCLML4YJE
W+yDauN7w8d5kbb8zeDwXC49MyFVxoQPJwaMeWVabEGiFvb7wa1HSBGIQWNL
rU/0VvBnbXSI2O/pI+xKJN8Xo0NlA8PRrKldppokG82xX0BCKIcuQVjk3jBQ
Q1SjdInH70V0ceFu+a9hi4cTo3nT1nFwz5Gr7nCQ5bw3cHvmJB+52UCIpMPf
19l2/fzAB8XmoslX1P52TtbDweA/iP0wxsg+cnegS/f2LOC8a3yiqd58SKx/
mJqydRBzv1WChsyLZJnzyXKRPZurRk1kFuAl83ujs1jBMGSwW+R22kxiJqhI
pCdMZNMGlshxKBDOH575ODRu3bLt2Sn8rfAzmoyLbDzNO2C1P1UkSt9B22Uf
+k/GoUtGSiRgqod8uSCvxsJ+bM8RJuv8Z1BhjBbXsCGEACDZEb/9DLCAsEnz
UXHTgqsO9z+PglcjGYjJkfc/YkFsrGQD6dXSAL6aGc5cfHTDZvPsW6zdrZgb
hMjkbSv/FJW44KPxq15eb/bDYhALOloN6JaWrYGFnnSxl0evgwdrY68q05hX
GQ1M6dJFHutwNhjm0hx7g2feHDYzJaQ7lDP76Jjbqfkwi7PhwFwGzjZlhWTz
8F1ZF/sh9Sc6UpEwfeI4PgLEpx3RC0knT0pv75YbV48WZykwKk/txteKKVtx
fuEArrEk10UPVGXYY5gFjcTqClig2+2sqVXLfUavWKj9ZbEpEcJXvDchxvjV
+fV79SbS5FEJMGFHYHDgvDC6+3ivC6GEHQbsLv1DFdcpq6uQeaKdK4CWYoR0
xParMjyR9d37n9A+PQG+PzBK0rQV/ma9RF1rxCKJn8I9F6nryt0RRWDsOemN
jBHbXK+yvlYkaBEsy2OeGH2ExXNFCWK3nH2OVnnJU5q3DVoK/UC6nhITVWNe
PnRCk34JTmh9pigzFkbCcsgQmT7efdqf+2XTgIMJRW7A+EFhH9sZDY1LJqbM
uir0tmOEo0i8jXw2vXUx9YhWVdrjd9qxTuEZqDJHd+TzpCSSwTplN9B5RKSA
dW3OlxuZlIdZJ1SF5CDWD0WzE6/odWupjGkZUFvNXdAVEm+kiNSi/wcwJtiH
MU5KoKVge6CHqtE6k7WsakD9MM9PjKV/+8f5U2cp0Qgv9l54JJs+qzobPKOt
nP0O8MNLzJFbjFdjwOpqUbdQfCGOsjEDALLJDR7zTOD6qQS0MV+wB4WmUjcN
mR4832tWqKsnhbc4oTFlXOzHHtYkkpZtwUR7xQICHNIMl+sAfdyl5/8sj30O
cihuc2WqpvhRSmO/MQeWGQ9PlUFb+O+eR/OE19/kiGfBqRL16N3ZZvHnQePy
BXL3z/RwCYsJo7cpkpZWNtQBXTJtJIpbuobz1z2W3DrB1hSxNkrNkrQu+DNj
UmYU3j+tg3jNPbGm0DzhJX2UM0MwKvdt7VIpKuixlB5X/zCTzMwOHHVMQ5J1
ry1nRTpVmMPiQD66oqK0wLEowdS6B4UfgQ/BJPrCSf8qPiEh9NcHRvW1LjUN
8GbDcom8NwFQLTVpp0qwTzY/EdAuiXj/pefz/gcHMr0ui7vl/N3prepUsdAJ
yXdAgUfh6veUrlai/3H2KzdLXiCMJeT4H3TPKOfZk527t/YLK4M+0kU1z8BV
REeASEonSOHBmJt7Pvq26d6VqiuFZkmbV4ALs1CKWcHWNispdzqb8LSCE9rt
toZgtgh74pwz5sCS/9lRaWaCrKAIKbtPkABIDRm2+iLcm5ERUQpwwLKaeLFl
Tg1RRqiFyUl6NEWTGR5RfXIBP+dvmWtJW+cYWFzkgVYL6AIIAMavOSZBnLUM
5IWgoUNy81aaFFp9OwbBnVELDrcASt7JXLnN0hgc0qkw/s7x3CDooau9Ex/5
9elqOzVAgHalLaFRuGTFVmUl81twWdmVwA8I+jy7sKaQBk0+DK6ltEEClrqT
w2dnl7TVh7OHwkuEkFautKEquN9XUNh2nvnZWM6cqW3TZamR87NJsqQT8IRq
BUiOMuW9mLJCoac7K5K88h+Qj3F3tyUVfiqj9o4OcQprkcH6g+b7tilefsq4
pQrpzk/GYtIvoGln+wqndgmKYx5h3wknCZMZwM0fe5XW0qRL8b4z9qCxMfy1
T9FuMCU29IdpcGBuVHhEJPr95T42zOVFgYp14RxT/VtvhWoxMm0Iia1gUvmi
B9e+cKjw2ZCnCcCYvd3J0HKa94YNKotGFgK9kZls87zhTIyo43EfQi8ZaNt6
vdZqXXy7nq+ImBLWYdpmoxM2AI0zuHPPmWLN0X2cRqUwqYpMGb5Sf3GPvHEt
iTYWtfkiYE5ISlJZvDwERPj0+tACGdM/YdAD3Z5PxgTI8F8scc5lSuwO3rD/
pzm32gwg7Csih5p1+khaqiXFWI8UKs+24SkFQXY2odzotdTut7jiwwedHe0p
XcCjUh/i6Gem6UdvL61D5w200G+R1C4PPA5cqhEiolRshxNtuwJCikaOM+lM
/cij/nVm9KsPWdh6+kXFa3wQYqgy/U0hx0shQTvXkKyiCk1Kx0mXvmdf9SxH
d0+lrSDS2OAtg6CuCKRxLBgqcg0MJ7j0D5s4Rj1TGrUagLkW8PAdpVnC0X0u
bOvgaW083PlnS072Y2VzUMKOIwLHiNQGE9ce+4o4LVxhokZMMBKQ1pj+ryyF
iHeJYiBa9RvwoQ/m3hVengiX9xYiD+WgcoWEiVmxDr3lSCEl6oThUSCOQoUr
TeutrkywMogSUPKPP1zDTF1wO4fzWpTU7ASQ6ZMgWolCVy2uO/OBJeVixgOB
yMmhtTAfK3SL+S+WzRD7gRBNlASod2ag73boxB+mI71ytNX05oaZHPc9Qrro
oPXgyQhJntmGefXlamreH8/QrLz8nQznOImwOXah8ZerZLrFFdznHVD2AS1Y
vtKqUXpa3QakJEniqYomuSVVi8n/bkhzAvr1Tjrjw6XPsTV2NOD8V2nIafqp
A+jwf/6jB4reAAeBOTfang17qoDRX6iPZwByNbIVgiAOPi0uaZq3QANo/VVJ
03X9wxktUB0ELck0uTIsbxv3z7nEZXvxe5cGTzwnIsEywFgPx61OotyRdIjt
hdNiK+KQfuyxg+OMTMRoq6RyQEmtq44uojb1r4PZIZEXsFV86me1zPjNQ002
HY/nR5323sVbNQbVsV+Hu7VFbe0Q+h2o4ncmFDi7ziaaZvvqrLSh7oby0hVC
JmfoqCRaRG2hXFnTShkIu7wbFrzZe6j1NtFPt3SbdR3wU4Dcobe7okrSNuhR
Ty5/XncxBj/Ho3MnAkbT3sQOflG6PHszxC4APZ8UMd4qAxJ8wfrfka+3kVf7
0CPsc+urYlquSaO6qxuRjuB76wxQe92qcLRbbZUkAKTV8ZSsuyUkFvOSN4AT
o7d2tze0YFfxVQboKauoqQplGSEXIvLMQuI5DWRS/SPB9b80lbW9PORQfX1E
jZxJLHYx3vUhHgGiVv4R81Srpe2qHT0FuXN3UgpemCp5SYSnVremnjHpxsiv
gBDLGVd+oBmtoNqMXcwoYSJ1DqIz3hIJ2wh9h6M+n2LhVV3s7y1zGYKKLtcI
vCJJovoe8qtimoWVQALP8Yqfh8y1G4hQS0Ga+PZTdmSKZRhAluZdlNvA6FGX
uLBDLVgJ92atKX3nnWO9IXyUYSMbrTonpAW7MAat22j9S2ci4ZeSoZOqxf8P
s0oqYau59ulNEJ8zskLwNf1kS2hW8+E1qoQBBK1O+tDqz7ZRZM6aJ5ZdmpiM
0pRqt9K7FQXosHfPGD7x2BEqrSQEth78g6n/YNB3adPktD9kE18v+C8jnnMy
xzyCrx8aWsPvJW/yrUvteyb6yzUPkMvHAsrpMg2WaUpzPFpkos7IG9yWA87J
vzQk7AlQ9P6dICEo5OuQ2rqa3GLjrC34eOoispLqEsQoGBD3h+l4A6dph2JQ
Vy+qiHqymls0IDEmD0RM9hw/hooqSfUpzwZk/jZGXu2gfOvnDI5GpHBdMoj8
kiLA7emaEpySCl87MaCl+LVlTSvZWsFxb5lwLOR7Ht9Qt9Ux3liETUiEudXV
AGBZhIucw0u971B4xMphNcIUnAu5hGT/OVhEXpCedWRv/fxnQQwh713PyWw2
1GX2wzHcIiwRFqNO3SGAkV71hn1+MFIrBlJRSlg6Gf9ZanYQPEfgFKPIC2BD
M1l8SNL4HyzDdO8pg+68HaXAFLho+hHPFHyUnduMdHBFOa56IWjLqOSmEqcu
nbHBuM/bZpImwRSeCoVe4QNoYYendwipj487Y9Mj/Bthc6MHrGuA0xH09i1E
LWR83fu8Jcx8dUXfXBH7gYUntIULxb86E80nO83fsNigWfagLtFLo+QbFL45
j9SSaHy4j5QyXv+X2NVbkqQlk0gMkBq/LTpVvT+h7odJc/grQ1x4DKOR3fw9
BZaaKlTyPOg7BNqVlt+H2E+qVakoo6TNmGHRRXJzN6qDmzMB3dfMxj8fZEds
KnEX7LsOz9+FU1asDiiy06tB0hKsHDwfJWxp3ebuFnrsh8apuBHXumoqPfWz
HLUETtimPoNyO3HmYVv9If3VkhfJ5SILT2vNAm/+meZDzLbQE7iTJK+U1+Vz
sKySY3KxXN1do+5EKxVIJDuzXBcDFZctiocxNGBvzK67Vcn72CMhkk86MzX0
3h97tKzzGtb1IcfncgERQynKB0jwtPg/W9AggslZTQpVS6XY1uJXohElDEkg
zGtXxClBVmfMfcsh2lrQO9POGI/oGNGmRxJ0c20EEJ/xdctCwYNcHV7zpF7e
y7Qfy8SlyupZLYY5Fb3ccRkv9m3IeHkQin/dsjRDSOFh4G7iCjS109NIGKC2
30/LgmYM3yTExX9Tye4GBiILFX1utU8Zk/aHCq1BIDie3965vYzS6P9fbhWe
o/xVERQW9NfRtcRatSSi6yV6ugjjT3UqOhadE/z23EZtuws6nfohti8jSs4w
ewhOyilsyXce/glxclq8zhFOzXlMlYPFYRTymVx7wr0EZ7G8H8W8hwu8hZTH
/eAEIo9+H1QB/8vyU4+e57Jml7gCvlQXj+z85Mp1ZAmQJ1vY1MPP1uLlqd66
2z2dwUfmRCfk4bCibRY3PW5AZELHYqS7IYiv8GtZrt4pCkQytYkN08Dja6wQ
Rg8M50u9CvBIDRkdhAmhs97H/2yWmbzBc+Cd3AzQNHfHmhwryxtOP7KgF9R7
0psiuuHIkwEhzC0DfFDl6ww0dMD+vF1qTwCV3448ITrxguvbmZckvcLKua2+
kXlobP7WFvCWyUL1rP6qnydNqjYqGzzhU516ndSLPph7kmMMmXw5kM0EKQQ9
RDSNnoFQHoorUe/mXXTwmZR3LhwKHquotvuvSZ+rE2D0dgk1geYzC7ycRD8V
jkUDIDgvr27S9BkMDCORC5U2s1S69oBIw/zofUqQTsHxOMXIf2BFKsps3oh+
bEgwEIdrGs75DlCAcwiGV8qfcnPEAu/e1EdxB76aYArsWsvwpiUeIce2JeL0
7rLf5aqd10JTTrgetsRgFdjt1Ax6khyWbKAv3gLFwXmGMN4iMjshPW0/gUxZ
dovUXB+0BtDXqwCRlhZqbeT0tLxW2H+FjxTpQyWi3e5aihoPrOVm76AuL+6S
vRCGeaDBPC6w+6SjjH3YyNThpsNfPoTxLJtWkekdJmKjYYO2INaAITT/2pLi
K1vxSKxmEX2ktrm3Jy0cGrZfhdPl+SdpL2ly5I7xmq9926cqT6EDAsKkMBN+
KSjy8OHZulnAJIpy+EzpY3zb31yyegcLUsFxbwG9QN/gC96pPLMXqzgiugxD
b5nyfEojRcx0oC3t6aEeOTsI8NQhA9iMCdHF2Sr8Y4kx+ts3oMw40z0dRM0x
DTcC1UOGA5oXP/fMpziYKOLu0YB0Yh824yqND/uZkIeiIXvwAwlRDCDyV1rt
LYoTIjo5VfPMPKQMcWJrh69rveMXA/jVItqiI30Y6bzrxyQk28BD3pbjKt3F
ZlRIoNyHc/Bmx2rUHyxIJwKk8NY4S/Stj/JRAZexU1t+lLRneryoBtaKOc7i
HJWSFapehvUd8xBaVdKcoU2aIspAktwUi5IKIlxpHZ7MBEIJNNvgmNC5PdCa
EiF+qRlXqxo8OP97wI3K58E0CGZ8eyZQIYQ6ivi9ROOlHylR9z//jJivuUFr
deSpT18u21ypIGM4j1TSqiWW41IMbRCzlMoNwujqQBYJwvRKc1kTxnSwOBAI
E3prrc6HzDkeYXq7/cm54uTYj3dWDCi96weCYoAgd4GNf/hHg9XlWBfWCGAC
Ju2OJm5xFpMwTJD2c6+y4u8AUw3M0RU+WdhWOZ5VJIsmLK/SKBaefo+enDlO
2gmFwjc0nkrBSSr63AF+S8aR9V2kBfoPbWuEqrcXIOwxWGDXe9P3WUd5UJtf
M3AMhYhM1U/uKElVB3WbmimXHQER9Ffd5DE71lYqEMVpD3tn6AWCsMZGMLnb
0m0tBNuMqtwjWi9P+bm2/mZws93Cg7h86UOZg92MYBAj6AEc98h5aa+yQlUx
9ACzaoMq0IA7oOk2PMZdwtWvFa4wFYvjnZRTZAhlucQA7VDMbnQAQljpLbcK
KASDnsXQz+yn7TSECzRqi2H3CrR49WV+4NrUstDpxo22/C1t1A2geA+kBU8m
N6YWWqgIOQBFV8TyNhb/MsOfCrY/jEYpr4hs5qUDYSvs5pLTmP3bpRyh62jc
I3uSxFaQu9xEguAqOeriEUkjb0NdgHVTpQDfhURsTmMreLuse0y/L6obFT/s
MqLvd81dGlwvr9PcWnCrJTxJgUYuL9eeAEkHs6ctDHUUx/4KjmUMJuvdjWs2
4mYiWpbmS1VkNQAPXmo6OthsK7+r2Dyod13zwC9DkWT2uH8RPM3kDDAibkGB
heX5+K+duCBI8WLwtt+0Ckzy72UXaSVLJk5nHWsRUXzNEPH5r/zzuzOtwdcO
5YHzC702oAN7RnOKtVpfHzNIYyrXmnfk4mJeAgBcPxHM5nqr2NEy87bGIxT/
q8ULL1OxRQZLwy9Z9ZXaOlNe/XSOi+TUUWjKDIttUznmqYYHrHmdM7XY1o2f
roASSmXO5jXaCtxwDxmCXRdIHh82/h+uuz7IN02vkJovXtIWUdKEayg1MFNo
pLbfaSPv4Q6Pp0+f0ds6ptkUXPHazxFR7aIu9DlfXUNPaCLsQTNxVNe+940i
st2I4Bl6fVeBTrlezrxFGrwxvsgB5tgdjw24Jey9dtOhijSG7WjXfr8HnBGc
eftSVta1VidtbKzi+cml7Qr4CzAqVJ6uPy4WUF5IQHf1LybQO3y8B7/GX55E
+bFw4HGS2BcPx8Eeo/pui0gDPsyVjFriqqSzrpYGSD8eFfvI32tR++aXjdCB
ET6qJMnChgEi25FiI4/e6eyEXmLSlKbQLD5IZKtOSZ1O8X24UcfpNuXf15tT
NdpwNnpxI7yA8M0iSaADGR5TbR2eGQ/ynF8eUQLYH8JcIZtREMXfEfBh/r8F
idBMFOkcLaOnITdQesZcL64Fx+6bELYJtIcjZ0fWtu7Xbc6hm9MIYv+YfrJq
ecPd/xZnkT77GH4EM6EDv8XxYmTbLK6KZvt6Mr4/yMO4nx+NZvwInOQE55tc
Ehb3QlNLEuTPcy75+sVLuCwK9iDCTqFR5DTV1Y28ppawrh+RajFbvdZgZemJ
dDSdWneBLUBFCnPejoaOaiqSRzxnff7CCTMIQyBb2hju2z5bE/mLWfo0fblY
L1mlHsPVveE91evl6LyNmvuVMYWz0n2RJSTGx1XYFMYvDm9gXVB457kDAZYD
H2p8UcK291U6evQuw+LRb3CK/fW381LoK1Ixg2zRy5Qlywtnb2bVdVXZij0r
VnceyCTnUMIP+IMj5bXTTQI8YWRbOCx5NxnipXSkVr1CIGdYq55lBGurSBiC
15E+x6Ury+pakvkv6Y99rKAiEFN+IX9upO2avtuj1HLF6CvJSU90/H6A6d1z
K3xjTK0GsePuxJ/edt2oIwvaHpap1jsmVMORQ8EOkdFq8tRF2gdQ9Vk6fYa7
LzteHkEnn0sVEXeVf1toCIhQxaVtDUWPMjSuqiIcMTa+DLYkDGEqGFg92fLn
erDzf+TKYjWzAzLwqKZRBKCGC4UxNJMfU31c2d0BPXuc9Vr5wGzuYb70amu0
VrJoQXX9Zj+nxZD7rS4r/nqn0M4qh9PS2cnp2ODsjNpV5K2+l6sOxnYJHsC5
5h07KipN7xxnZuIhP9QQCYHWN3LEVnTuAtju8zKRoBNxoKpzSvGxbYiIKvO4
+Yi03JHd2Q3l8/VoQxE1EkVUx5mRjyG2YwlK0YWs/OYIgv++f8HlPPy/uN6t
8R7K+BaTkYP7yKRxwIE1Q1GEXgf4h4s9X8aRuwY4NVq6CamRvZJLNVuHd1La
sXYLK/VzDDeWaFlif/5XlRJC3m+iMjIYNjSgxUK9pCVrr9BGmUteXMvHHtVV
F+fO6h9E1CX9nyp1LAJD7/NDTx4nTezhozDWKf0FOaFJmxXEO2m4F+i6NPW1
gFAOR8Du7c5LbTsXkT683CGJmBPVbGT+CceWsBozwW9XbV6UhSdxD6/B70kn
+NgnA15oNfqtU4L1WVQ5Qvk8KYinbF1hSJNro1Z2eLarsVmG5kj5LgJYI1yB
HaYy5z+NIpcu5lx86Jw5v2aa+wz8U1lcvinJJaRMGZ8jG/WFqc3J/xzSAvUJ
Sw++0a/3m+Aq8ueSvcW5h7QB6alfSMHz7ZK6ClpvAlKdXduvCxtfHyYCZYgd
eZt12QjPl5n8+HWvDcvdVqvuaGWbs+d4b9UUQksdOCHHYh2gkb7O1cTgATDt
IvNdM8d2U9gZFRLrHwdMoxVzUiBIrmHqqnGIyto2/vcn2HuEHjo57ToPzrj5
AJAO8Wum5HjWx2gYKVI1xR7gz31GgPoJrrjnqXJ7CysQAc6R/dc9lZuvhEzB
5bxwmgb18NdsOfGPME6guhkvCiompQjaQHRo8VuOdI8WVdn5cBW8jhoP9j1h
qV5wG6EKhkZFbA/Sy3E1sAq9Fsyb2nTROxTMM4TBsy1s17lEM6nkri4fzp+t
ej/1LotOtvAfJoWzip3WHDTBJMCOJBQb/uX3oE9Tck3D00xTEfy/kxHmjdg+
PLU4rs+zhnYfMvXwusUkwBgpzffkW8RK42Th5d30fGe3rJJ5GQvMutU3ROHq
WQSj7urfj+9hXRQfaO9/WzcO1/pO/dJXMHFH9imjqVlixXkXyRgIF3f5l4eP
aQEsOyf3c3H9iG9BRoS7iLxQF66d1oQW2i17uF9aMKuhQRFvf4S4VT3+jOKR
Dp62NYN+Ilr8vTenMtXN9w1n0dETBTJxVP+nvdVl2Kjrl2lTB0VwYWN4BTWH
wuudCeVrO7W7lCfPEPOqWFQBnA6plH8ljaV5UfuRPDbK81xJyl4hZKapOfSM
6QQY3guNdz33MjwQ/IK115PiNPhD9Icv4a+uuw5MF+diyFJSQ075cgHgfy+y
hOkF5AOmpgnPU2xs1jBzEl0hfJAF5t1dBwfoqjpkLSc05zKAR8LH0vXws1gS
ZXUDp3WzA3w1h3N+jNhICPOyvk0SEN/VOEfFgBciNBK85k6Wp/68VGMcBmli
k49cX/3RSOaoJorLia0uKOFefKiKUff2EgQ+ZH2dc2wdfaT6N8lxiEs+UxPW
GZsFOpMRj6AV7rmX81IVHx0T4BPTCn499zU1RoP8kW4ZQkOvHMWzqEGwGUm/
a1wtjqYsFqc5AnYY39ls9fP7H2RbNdXQxpt1wNvDgQQ918NUewfFOfEC4tis
hk5z0jVVsN8A8I1+vkJ5csn+BmcY8R9OWlX9jQXf6FVkVZBZRThR3Szp5ul/
1Lj4LHAnLJUt5bpMl6gB22ki0Vy/+F1rEJsnH9Pi/EoMerAi7ktCM4zU7Drl
1JzTXZ9Fpyn7fbL4qtl9XlKxQQtvaS0FHlWLNGvCOFHIxl37pYXhrMQemBsn
YHR2gpDCQUXNpDyZKClQySyRUruho9PErodbEgYSte/x0G4Oavzwqai0htnf
XJymx3fyvSrVz77isvyv/Z7XifaEsiTyMf4EKAviobK99xjEk9xivT9GBbeT
Sw3v2pGeMwrBP8q8bGeITKYEeQsuWW1J1wxBEJqyyL5L8UQhZWzNjRiVxUM3
TgfyBH0tRlxdhIot4jLECZymxAONc+SfWuvOo5p6N2Vn6sxYVR6YHDwsn9TB
BK2dKLJZnRzuzPmejIxLSyGtbJnVxTQHdt5fowEvBn54JikYIkde8etVdCN6
sdO0jWs4xt9zsf5F8ZxcVTaDc1GHc1Vk5L1S+rAkMuzaQeTA/UczqF7GpLlY
Te4k7hWnFJiLoUFz12U/wunmvQieFif8Xc/xZnDbpNCpZVCEbGHgaHPOVLOg
C5/+xUW7Jjtgo4O5U7Rp24cYEQlu3Z4Q1BLzyyW1e2VUmf/4Qpti1f1O1E+v
ZM7HVG5oMwu2wTqR2ppsUh67nF+9aIvgQrUj4ovcZBhWFj6+pcG7J2WNHw21
37WCXGQ1Ld6vbt0YJqkQNmGt3e72FC+TVZGaQVWPmdJvKWByznO9dUnsvJSW
4kVsOB+NQhG4H76q+fj63ZnGo9BNvyyAsaMLOK2mFHN9QrQ86N/r69UDHK6j
1r3enlKXHKwhHROoioFi734ktDzAo7e5higR5DATDgPmSyNWEnqumauR2gu1
LSzNmEF1549I9OAWuyiDVUgvr7HEawm7gZ4kM4X0cpfap4by4Pe2NfWqXLwC
ER5gDdLO8MlMS3Vk+BZsQzCw+wU4y9t9UyEOshXIyy9f6R4qnLckhKHTzgQo
qo3FOmzSNc4i45hjtPc5y5VCjVmtxuclfwpvS5qaJcmxv3Zuc+Ok1YITOlIg
FazXxahm4OWnm4OWToanvLN4MvcoYtoLL0Hzp/btqkZynhDdN3Cf9XChjb3Y
zPdzr6AWhANJqvm0vVcNKXyi+ZHqTArBq+zrdkBYpLkeC0KwT8BdyfCWSdBc
UMWPCio9JP+81cihabQmTmjv1JyB7YNGXbx08KTUSgssIBvWGhKC9K2T/k3G
+SWmCWuUT/jgM5sj89jNUz0cSaMQI15e8E8OEibXh4ihFHDYO/9+FivBbbuc
CW4mZ7X3o0dMqkzlhyOLp8kV8Y30Q9zk4mNI8+vMJJpx8KAex7DKqc3GQXL3
TCeuAdZW4/uQkXzoUH/eTgZa6Dnb/tsGt5+Sd0LLtN7N60iZQS7ISgck/a8G
GPHFUvb/g6PA1WmMHju7Kwiz119MAnqBCT1KOXzdyrNw8GDgrcgm/rYLXah0
xacDiq0uqnDKlNWU+RjoOllge/YSZx42WzeLshtAZmePCTqzs3SBIUwnPhcI
NLC+JEuWK5WSz1EjrfnOaee7ExfGP4AM1h0MJQhXSgK63a57LmcZ90Omwbo3
mZjE1y7tJtc+DQHuTyRwi0JXWrc/7srNwrQ4DDROWan8kSbJgBp42CTiJna/
NMImtCTh02GEqQo+1cyRY1xp0j5NDVcrjH7n1sCWQtrliDo/G0144XMbxaQa
d3VNukatp1k3qn4D1XTPIOeLGsSsSha7YW0b0FDSUIHW+E+9P5ixRKaAacJz
y9nX8zm6jIHyhDyk7I9ZbnkFYRY5Inz4qKyTI2dkeTUuQgghqRokHo9/DZYk
xtOcdkJT0L3NL8Mr4lEDZhsSbfufHR+XZPdTpSHnxXKtWBZeTXadf4ZLdTfS
4QuLATf6Bjis0EyX6+iRHGUPuT9kLMPH4PnDWAPbV7v1d2Ch07Y/jfB7Jgw4
Cl7sGCdvXER7s4f/aCS0VaYV40w0WpiBH5FolHLaSgGmd2wI9SvfTd5+50p1
X0Jqujnxl002WFBXmRbUwLbJK/474HCIxAd2SgXROs6yFHost2pRTxp2Wija
CFDQwzsx469lsLJ7zYs4t0OoeArFYjzJ02aC+eEY4C/L4F8u5ROryrRP3BT6
yOjCh3rTezYT4Gdw/dJutZytBDbtLKFK8SHtbfly3Fwd27rjGmRIrHt4Y97W
apIz8Mcxk7M0DnnBb06u7g45/SbzTzsAQ1B2KyEcHH9RuUf31MAp6LAI8p5D
rS20TXcbzfzen3Hl7mI+g/FkG5jyDXQ0SHJbaZxqLoSCCMZPNAC7JBVfH6Vb
MPISdpCAqcbmzfDtMS39shca87hopfukpk5NOBDUKl0HP79IGxYb/MdbtnOP
s8Ml8cORk+N/KMMR7caDiS69EA4NVQG/nke2JZxj9emxKNmcEAc1a5P5KG+H
w9ly74Yr9RVPppK6t4fSe+gT4By9/EiyxzM7TONIQTBfaRH0KebK7HgwB/wU
hR4vyD91f/xx+eBhvB11a2rNgARQaCL38PTPvSO5N0tSx9W/4lfa4cAswOyo
LlSZhwmR0+VU+AtDcw7Q18iojatRdyhcR4ucZ7jtVh+zHJ81Ej4pLTjarYIV
7wY147log7yB2tfOC6rxXTmFnyV5SvCM4zdLVrY3Cw0ZnEA3Rz+5sndCI3iu
zrLcSZBXt7fDzuzVXgmRkOAqiIzC3w34PMduBipMZnlBsIhHUYNoc/rrc80I
xNVk4EC8hAbPsEYEh/XDUeo07d5lhjSvcXwuKjF+o2UKb+MBODDb4AUWKCiX
Q6LPzQkyYFa4wAh5DdMfzhtqG1dKDrr2bKRdgrFizUhg2CysBFDh7Fe45vNs
cEJPZB1sj+eJYVfK1zOBjq+L/33bzboBwWqWZ2QHmEt6AZ47d1AiTOEJTAwP
WmZYbHCO3826aaFc0Q8Y5+devrpkEmlT/Q4x5+CtvVmjpba5yWY3KYGQoYii
HSE8NggouWfBMJEi+981u3pichAa1rTqL576uHQu5Zk0IJ9HKqEQkFZzIoH2
bL0+e2Q9XajtMRIOhuF0KaJeBhJE+32F15Gs8DkG6jBGIwci0bhIzMpSiRst
KeUZXuWtZ94t6lijI/GWZOV3RHF62P1L6m1ApqIBtAF/tj6cHSzn2++ogf0O
p7ukaicwzXr7NryDQ2fl8hTCduXdq0v6RwD113I+LFVeDpoS0lysuosX2tZy
4QRXGBZvqrxII1tHUfY5Gnx0s2wK3kxZ5GytX9N0A3UaFwEvse0vNaXBgrGx
fGr/Yct/7ixaBT2FDrXb/oQI1kEC+UCvtnHtu9DCeueBv8h56UqfeyVmq61U
K3u8VGqjdUi5vn6HZeb0hgZD2lVo6WahyRgKM9fKI/hUQ11/51xTowSVFdeC
ngagsWDU0hCuvZOdJhHk3SgHc9smIkl5jYaLN/5+m8XBcmK4JlYL8z9wDpPq
j3CkiFx8G+z0OTNIwic5+rN6tkZ4GvkvuMW+Af+lZRFbNS1X2h5pgjFh4EAb
5HRwnJN2n27LQ9hVWG7yk+rUWeph7alLzBI+B0ILO4x8Cr1wB21mPf0Rt21Y
blXG4eNFTAJYEp+eEXwd2yd3WosfJF13Diy1OgK447gkafmw4h7Ep6Fxpa4p
1UNGuSR3L7lLikeNf0+gclkeHHkxIiG/VG/SHls6ioNGNoe7k1i7urJ5QB3Q
0KNFMo95LOMd0gnQVhrMRkXG9gqnZVvmKfb/i0fVBYHNz4Jy0/bPrNcHlInj
J/WAKvNuuuqcBwMxnbl5bYDbK2H/3hLuHzY5/bmG7DqIrTJ9IQkzmu3U3nDK
xIDNMlUoPr1fyCiQ+IeVXA3yuD9Q9vmD2q9uaavbHIBf2cwsh89wmgLtSQOM
t8yVS5eonUFsgqEZwBIv+XM00zNmBXr7koUDmnfZkIhi8Hwj15qsGb0h4RLJ
1pSNGtUhm0Mr0+PZfc8ydYJGnZRpgMUyMsI3y5du2nskZwY9Pn0CbspGo/up
oz4jpapnMxBwwCmscfx8Nswwf+cArys5kDAlSP5VV1XtLOownKqact6xMau7
GEZPiEORL6hEm8Njg8M7bQWA2Hooz1z6LUEy6Nw1aG1I36e6aXtJ34Fw2ZbT
wEgSfCKbU0BLo3VQRiKFwHSZGITLjRkb7FlBprUEvTsB++vbqeAHeisasPXH
nPbO/SD8x+LCAcKSuk6t3alWAviHNQOrnmEaoL7t269lpqggRKqakttyVPUG
+LpiFV28ECXf1Q+Y0FLb3UwIXr4U9TY+Cdb9A24h4aEwKY6LC8u9X1Hqz2Yv
heSf3pcfO9d1vOKaD5o5MYezh0hUjvGdnTp+WTeevUcgJtPJhN6TlQ4xxa1i
+BO4pbKIuSZfMhJExkj3cw55LgYNH6zzMdE6Vs9+w3HgwcE/UOlq+TnNbCCf
1rY20fzbCavpnFdBfyo2AOIJPnWyxF7GASpNbMVPusa097I1vHSwKaK8HNi5
62SSvQaZomJbfVptb+doLN/DfQFDLfFMJZZ9L1AQmcftG8H4bZ2rymNTHfVD
M75R6fOM3wlDftMLFNZin3/Z6xECZRsSb6TQ7C/GD6a6khZ6KcxL3HwVpQ1o
PEcMlU2s6BTNXP0K2fpDiQQRuDxejcvNu9aXOgJv76LaHQOWkaTZ54Grf+9a
1BYsyFgbPq6PC5VeuNqKclkkLgaKrkhbPAWz1uQYvbc8e+RdpfSQGYLBVcL+
ujEMh0krh16xWTjI6RNaUHzeTPyrBvrY03QYeR5mIOu/2tN7zE79z4pXFaPP
sxMdAz/iuX7Uq6M6r7dQpBKqzomqfrn1IbX3lmeotMfihfcsXQvhfdzIxWZj
+zTQSPevt7x6OUwnxj+YWW+VysPpcIePwlAnQWu/V6FYzdrJx9ESdFQY7xLF
MdeWNOS/B/bEHCBmhNJSIh8HxtPXuY/9lgKDQk0fdbbSP8NxQcOflUPZQfwL
h9a9lGL8LK3cYyKHJdWFFT+Fvwtayx10KkbFYhJizAEeKgXT8QGOU0NgrMqo
dIXkaOUmdmtEydxMmkffNFcIMH7kg1uPiun+YvTDW1OyrY/HYSaY8E/MbaEz
zDeLjgYWo1FjPg8TLDzE0QmYlekytc1XMW3wpZcZbEZ27Ts95F9okk2UUQAy
6Iuv+rhNGw1x8LsXACAJtXfu+de1XtKrO8KSlHQrkIeLF64VREpLbsUEXCa8
kp3S29BMW9/8VmrN0I+WTq9nh82y/MPBUxZRSdp0S8+hceAaf0n+Do+iNPnB
u++K6RIZWVkLEByJZVO8S/WQkItJc7G74ILlkm1wyj+TBzVrnPVq8BukwaTn
DXaV2dRTw0+zqo4eaFQ64xkUcHSQ+c1+Oe8y2EcvqgNMf8TgNb3iOomoUkdf
kVu+vM8I9v5Ghxv6dVjL8hznRlFBdksjNIrnGagG/QdqXCqDLrgawTPzPHAH
XHBv4PFPwb0tqPYTH69p6ytBYuHMKhUG9WDZsQvqKiHwQUhboifzQAyLb+sr
eTlAIutds5lAzxHlNpriZjSEzE4AW0dOMRyNTz3OY68pGLsQTnXgGHHVV5LL
qMG7oH79TxXGmLD+eOXbShpcbPyfR2swEmYaaDrmHwMXdSztvTIpd/Ueo7W4
v1JhygeMOZ05wO8tuPaLt8V82NSKOLS9RQ+MAvIUP7Xr04UP7Q3pMaEm9zvL
oCu/epgonY2LmarJJ/V8jwmIVELyySGqqJqvoqG8xci0XWut03Yr9eB+bvOH
t7iHB3Y9yDT32SGC7hukV4fRk0JUmhi+RNTnrGL+dDcVqqXMhwkHAWoSqOVu
JnNAbdAIh0YyVUbUHrXrydjHTMm6aFmteDIJiNffSdHR3ZGk7JUu8O8owT5z
d3+aNzRMGVcLpJio/+COW7I9AFRessU1co13D/IaLhq9b5Q5F9UT7AN1w5Am
FqZOucrgq28Aa4hLuMDU+8QicBJ5HHjXzEvca6z1CX+ejk1Wiv4s+ONJ82LS
4s9TOe3BIm/YOzvkrSatOri48Z0syqkJNsrIrGr38WP0Xj5AxjYNtIEGFkv3
F+Vmyw6VJwoS9wsqlk/B2yvhQy4wL2wFrFKaxsMf5oM6Px98A097/1cjOJGK
yGKuLASDJuqFsPY6pMPAxHoQ/kCEszVRSV+Ju6PGIzzUVGdTfUDkTqYFDFhI
74aYxgXFkuk4pigSffY5mdjVBKVHvURmk+RHs/bau0RIqZ4ClwTCuq2yQQ/l
mq0QwtkrCCMlKsloqCnGW2HiBKmICU/VkeAn/F8OeVuA2VGe4Rv9iPBdC/JP
pnFQsGpK1ZILEyW2ddwSiBpDNfQIZEpxGYSYA2Ajw9z21LtyhEWkbbVu1kYI
djUZ14XK5qraWDIMEaxOwr3tDthj9MoFfh3QZqHn7jn3dkUsZCZvsPU3f3SM
s2P5YzwZW1fMwyF+fCvZhi962CWikk583NELjyagATTIO9qd3xZNPGhs9MJe
F0Zft7i7h7xUu3AOS3ouBb5gHPRsckEebkpCzou0UusixXC91n6KKPQfTKI4
ZJE9XfRexN1ZGu1pM6/hbvD2Dsj2vOhDaqvYbqMi+YEDMGxJ11V4HEF3THaR
7E8uFKb09pzOAKL27crkuQ7TLj5ffb792ZGaK0H66HDgJawy164CbdH/gzxf
kP4+L0VhBMkErH/gl+5rp/moQbd0s2gU9Skvpa6Dg5b4DEUXy2ypyUxZMdef
mBYF6TcNp6G/ifcAKyfJk5lbF7EO27RwPKpuLPZBDgeJ2dzI0Iz+HUseSIUk
P6yFoktvaMo+mGVFZli4JtkLHNJjHRFXNJYRaZSAhFo7jAEkpUxPLSV8vpHm
qxzwFvoCJJPkZvHwDai2FgBUBEYI4uhQepRjanFdEGx1IM/aW4kzHk3RBtNl
9d1YiRLmxdKGoLosav1XsFaoWgHTLRtuTc5PAUtDQhJ+7gkxkOnHvPp9mL7O
nMmQcdY87JsgAl5NxdB6RI3fPPN6+JWMOKltqUR94nKevHGbh7712o3mVee1
6/BfVyGpzs+vjE9EAZi66Pvn8ckuUk/BhPHxjzJs1orUD4v4u33yMeYHqNg0
ODgLfkoRZDsltAjmuRBMVxTkEF3jvwNL2EYIooFX7CmSsHQC9Q5+wXA8z8Q/
QqjmvlfD6/5W9FBP6GufnjSgsgZFgEGnR1O0l67lcvsUuowtGFAiL8ud77eQ
fW4u3YaaUz60nbKi5jK5SPpvK3SggWwmpS5K46gRVFMO/Tq8wU/vQbDFAqWH
oV/Jqvq+n2ymILdWa2f692p0TIVXa1zmM+SmzNziWMfap79zhMldbhHWattH
VZxaCnpl4ugdU3dvZt3q0+NEy7+SrdEiXeqQaMejTGTHt5RSGuU3ro+DpLYF
qyht5CVz+6DZkoLTE+dTVEUM0/fUan2wznlsbuUjmkG86ar2bxN2BrcQWVOP
6qilweeE0wflU06pp7FkmtLvQv+5DwkMtPjLXK2TQ60UKaMYK/d2FTdyokEq
XFQO1OKhM6g6B4Jn/og1/Q+a7vvacERIFPyOIoewtyRoxhbqOYEWYnoULMlU
o/JwsYvwBZ2hVh2UuxbXPH7QuEGLWK2dWjMN0B2HA5YgTw3gBZfBreTb1lsD
HbTCbCnFw08uAykFhRQiB4wC0IQLMghdnZkbswT3YwxE+k60sR1lv0aBaqAJ
y/IcAlT4I/9CWgA21FJLxbxo1IJjeSzMUTdaVwELt8sCif7aZTIE+aUP7ws6
XYgW4J1HUQbYQ/9PhBNzqxtd+blbAajxLh4E7wuSLk9gqIq0n7bxLRavrRUr
nB3PJBl+1AFYR1Uo9jQuWWACHfmSTLnb0obmqGPgLvnwwRuVsqkJzDbgWft3
iDseRe41JzolxHe6IhPgS9vmbQlgpWhVnOBmCRCvQ9L/i6eQYOTroj9ryxHN
wDkIXEPDAQKglwO9iuKdXSi+jNYJ62dzRmSi7a/r9+sl5PCNa/MkFSHYgNKO
Dj/wMLBXFveoavigd7coBHf+fRXE64ytWMoOTg0o2X60NRsnxQrlFzLtZTFH
NbLKLEXumCLMl+kmqqlJc1oZ2D6vCAR0cPtqDpc5ZtPBN6AqVl+wxAI7V28s
XVXre9l80M3RTQsmNbWxM3FXU+tVXgBiGBgDamNYhyvi4dZhSN9hvcfRfoRs
pk3JLEZhYdzP01sd8m29DbYvQC9cJSXKFZA4+bdm9nAQf8zzZbAoHi5zsxvG
urnWVnAB68mWFR6WKPuphy4EI42JGtomGWus/7kI7S+pbeoCWYFhESV9URNe
8JkMOzoOktei9rL9rDBOVRIS2KGLTRaMEBjrgLUQ0RMtUGV1A//njzRpYTGP
qSo28u3F06QhylSI4e/Sp8d1RGyz9kPvxbYPNTNLqC+CumfYQ90nI9JoZ7fC
uENCcdg8R9Sn36ip/HKa5F9pd00SjaB0bKZnOfeBnfyYdhkxYiNh0xSroFoJ
U/y9FVrDHsJnC/uF5wywrwzIKnDGRErBxh5XNjYVUJZjexcXGco0xxVmaLyV
QLbjzpYNrxrS7reUGHZvaEf7RW5zSasGPgiLTMA8em0NB1KBbFYeTLZ4zVdm
dz8TeydDUlazszhbxAFPRgNn0hEjiPAt7WywYahtCkHOS15zxPJeeekTPWfO
zHJLESOZvfOWjKmcRs+YzJZafbvzdIFH+gU4NnJBFTD+AjhuNdclG6Ib8JYw
F40P9YJi/JUdwmwkq9TI7aWQAHL2ZWRbdGEr7bRH9MfRfE2bC+OkmBshEelv
z8iRz2Js5eMgM1wXAxINab2JqCqneCiFa5cyzwxWtSd0U9cSnp3+sn6RvTbp
vIxLjzRj8Ga/httI7uiYD5mnT8NFyWi0I2JnXVQDCOkC8eHmSFw0/aM3EN0w
k8XqpfPwuz+SKOSCZ92xVMmr6OKtZka4iAcK2pYAsCNSU84LRxHEl2ovF/m0
DlhTL9V6GsoppFiy24uOY9quAG+TU5Piisk55vYNhlZul7dO4rQrqUkjOTol
+8kZFlYnoIqbLhzbDnh5B+syQW8pChBcBlWfx7wwctSaPRklitjQr5ND3u8V
gC9XJ9QkL8Q3Dq5EwPQSIY/3fiaK7+G8SlnRZPQMIGlzdihbdcT6Srbw4c0o
bLUXoxarPjNeoPgvzDx8ckY9KeLZIRZUrC52ROyuWStniRiKRO4ZBXnX69Z4
TkhhwrcxxTTYvZ5EO6i+3Q4K4HXDZ6zpnUgB2VfvO/xTDb/8UeNkfexP3p/y
eWqQc8D+hG/NXf6bvI9JlicqvjpzRI3aqZN9QhzAb0uhGSAqJjPnVzY+PZNB
z+ilzvIF8Ksn3H6eh6MdARw7E1RIoUKi+Pbd7G50BNfbPdnK9wgmQuiilabP
H6hFJ3WKf90cvBUxersloXRdedTtnCSEaUz4SBD16AuUPnExQeJOl78SCqdx
LtGZFCkT2QmZXgqQIyOD4iiuG5j9ntJ3vUIQHAf/V0E6g6H6sSQ4zM77YedV
3yMRqJTI1DsKOSCDo9KW8C7u62GeL2QIT+Vrxft5mQRu+bogDLYB83Ki4ONB
9wv3D9sIw6mcR+t6JSKmjzJv/u86rvm3AydBxji7pdu8LJA9RQZQhRm71KWt
OsZZHGrcfco4lGSNDKq4ttlfvQGnZHUo9wzygAuwtP82p3DvJCov7+hqrZ5q
pG0dVzYFMufA7zoLC3+0zwT14fMvx+4vkMekT312qQ/SyMOx86qsA4vbzkzk
YaYIkjFJXudON63xaO1RW1PgULly4UFZzVwQqhPKQFDqcyUtuggyzM2a6jSv
ZbJQJAZNF6+9VLNf/wKXUgemB9xivDL8dOrgZmV1dTzulv70l87SaO2oGRTR
N4CMpibdO/dPT61HRpxrtZA7GzmTB0RNtmYrlt4Vrl+bjgh4RuG4toP+Gy1q
BUhpf3MVUhurdP+lmni5HV/s68ALFoYMq44h5U+aeSEo2n097s14taW6f/Ey
y1w6tEh+2hee3GImOt2/e29R2jxnuyI5sUZC/8nRJR0VHTVFH8McjGj4RVUQ
WsdgiPtLzzgIsqxrak9yQVcTphUB8nAycFNrz/1Ob/qhzS/bGgXySKra/b1V
OwJJ9K11tcVXnM4rGbQxlyuYp+Fexg5bZFhCNrNj3Ypa3zPLpkR2DOF4BYdT
uQK7DgEdeleSLrNyy8gglpvL2pPIWsb0hJhkO6DIy6W8plr1qZs71j5GQ3Bq
EIZyqw4X+riBMPopBUzCjpus+SeoX8tdBATPwpdofaa/hx3YwwzvC+4kz4SS
Q9vRjqC0TdLtyqLGhptfoWmOBsCCEcWEAOZAO6jK/Vq2KXk0sBK6HhevEiEX
uTxy6MePEUhEUsfK2go5bH2cjmMzCMNTVb1myfJh6NPOIBOftF0ue38lRTgn
UX8j7DFKWQIcPrfIVWoSemLPGTxq4/gfNHA4f2BzLl4LQ1N2uyUriSw1Dhif
fCylaaapKdmMKa2iJEW19t2BQY3lJyBHPqo1Cr3t5Bnn1ns5IPmJX9ri/l+6
ONcXWuzBJD3WKh6BeskFCaKAWqtBiJRE0aaWqQJ+WWFI6mC7iasePsBaQ6Bx
M6/4uDxpHvcyv5MBRGD77uoDfO139DLpmLeK3oyfcIftxlNXk5J2efqog5ta
hVl26g7As5Kv+J257QOqraItS7bGDXMzJCYTo3930GzyGYknfB36qq6aImPF
z2nDsLZMq26lk9MYRHaFNnZzm9eg0vbp8DRqcyJSCyeh7FtyHN9XIwZ+BzmX
8QyrtaaksCvZkg39TnzKLRMA703SdVpsX97oxa4Mdt86CSisMRQeV+8eX1aR
Ucr5PWP1QLP/mm1clmPdq9GjvopatE8WR3I0tpnreCQbCPZ9d06h4alw9JLJ
/9yryVQnS6Wg74mf2Mch7wdTfV1NgMpH6MITQ9ehZE7rLefQUvgd2zPzSwWi
8W5c/MovWK4RjLl58TWScpyUqyPXJkPj/FKMrMlzjqe+eb1sqiDbLjPO0Sql
tjV3ZkElhjWNVj2UXitBVApAtA8R8zrwkoxGu5XkomVGpMiGb1fUubU7VZLJ
8wC5fi2GkQMlI8DbvtgWGCb7hRwZuSFLRTP+zzulK7MolTE9AFMXSCySWlwi
1CJA8XXWZAfu3bXA0iVY2ua1B/pYQvP2Jfgv71ABhS7JlhclnoCENjvYNEfe
aouIHHfhbUr5GRY7IFJaZKYwmyIWqEecEuAo6NXicDJyFanb1gDyLqnMTugg
uaweycUj3ub6bIUo76h6LWTbv60aP2bmxb21YtZkFjtxJRsXResskoKhLtpC
s/jVT5Y1i/NTwtedImTUnr5mD+klqn9jb+cEG4O+3F0w8flq+gpz38RRTcmX
qXKuVUO73FfB2BiGgZG0dSO+TJ2fGdLrN/2vAXt+nCm9STpQawuV4HhvCB50
oHQcIwmQY27NWrH3g0omvG66XCQ3U3Eb6J+UjuJO4zSgoHVAtuuBqkNvd7uR
CxjBzjfNxVXv6/MeYwNNTUk5py8vSAo4iZqR5hNVXZ9Xt+GYRjRioyihgssJ
IT4eyol9U/5lyDu57hoYy3rXZxSul3dZK1ZhTh5Mxc7ZEfg102Dd3u6M6bJY
5ZG2giibtjPAqO6uWNS0jMNVe/kL0QyFjgsoTm/0IbhW5sUGcXg5B2D0aDxz
6u0VC+UKfuBDl/yvOdsc/8IN+bEeDvhaqyoB4pVeG3BHSGJwDxYcNO25UDYH
nUH9IOOElgmw8LasiyCpriJJnHB2go2IWKv1zL4xHdWnxIchhRfQnJqHLPFC
a6eqI/uwEgrt9S12xobWAHMD4o9ZPAFEGDkriswyhz/xwqOGXTpNeznpbkHH
qHZxMafNqrtz8WVH+jFOpRvV6q7iZEYqY6ZrOy9qyPPu+5tgj/C+lOLV2syV
7qJpNwpsN0uC8rzAP6C+EPQS4LK6McVKmdMGYpvKzlJdzxEkGjoBVdhJrYvT
HAC3+x6scaeZRgeD3tT89N8k/4sIY4egBtV3wpR2fRL2YY47GBzntf4HNTz6
PcHj8xZuJoyYiAsrNi/SuYWp8/3QKUwQD4gkoJmqrBcln0kZNPosbshUgC06
y6D7wt5fESxRuzccg3n6RQibgb2ye97hRT7319PGuEDjNR8xFDLzt0qpTSxz
GQ4CS3jWjo3YJzi5xD0vvZ4bTvplWFXH6WLwXCDLKeFwWUfJRp6v1zMJLONn
CZloDMXSuGFdDF7rDVMYjJDb6abJyQjxe9rqA0r5nuu/4yKkoYRxGXOd+q/T
DZ59YtEz2W3lYlyobYjFbdEyYy+jIrY3MiUEYV8UwvqTkmsJerwcruWbG3mP
IGKyU/yHCcMuwaoaWK9qj8D0a+IBitkAez2e+4RwlGNMdUzCVYDrzYI5eyXP
7oF1xI8XyA80wUjxCFcE6MIP3VsjGOWNJEBJ9RGZfb6GPDHQDeS4cJnq83ys
gGTzFFE1Kv27o5tG3WvTx6i48qTkAIN8WGGrULt0gSdvNWK/1LBvSVi1uBDt
xijnUXp0aY0vprR1ZWwZ1SfZA/4j05rYmwlkfvt9DrvNQ/Cnw1D1RySqOiv/
DPrOiVE1p3l7T0o6jjDj5FUiDTsbC4dsCIfstAoEcC09Z2falqZVrYT4ybFf
Ep9ZJlKgk/xCVEwTaB/2jokf6MrQU9iQU3NqDW5xMLEL7a4MklN3amRHX8Lr
S/QAl6jtzkt2igBKPGP0aJfSZBzNwNv3pcLJILopgkgd46t7Wh3WhLWQeMDI
TRw7Yb3KsL94CV+ksxCMr9WdMRU1T7Skm9b8xg9w7QAciRxzoPgSjhfwZ3eo
DLmnek1NmBlsUwLicSl3kFodRBBdUa88BayhyyhL+XmmFlYKjVL+B6NknG+r
RrvV3nBALmTEmWpylSe+HKoIBy0ex0cdksxjqa++WAUPN/Sof4qArZOahZRO
1gC3P70r+0KGEXwg6QyLe791x8c/GBZpXQDwZcrVblvuZRfZb5KCdfYf0l20
N/RcEVDaV0tJwHrWfXEl2xOyHG9hcgAhqQ9Acblcg5aGrRniNPheKQzrgY73
7orvoXxt+Cn82gnLbb09WvbETRuXdopmTnOp0aOzYt4IOHWUQpoSz5YKu+Yr
M1ksAkqIHuZfoJMgGTltFu+nY7QgFz0oagYTVJALaVk0LhVjZBW8gu/0A+el
oq9SqlL/h7TX6J2sDtC2ovGmO1eeVtxWTnqpz3xYDVggQgHwt+wUWiSOpfKP
gdW6UMWlwoUbHjsqblTFo3B+cYxm4T2EN3v3y2F8FvGWihWhM13oqBZFfLR3
QlQqL2o3MY8WqjG/Z3LIeQguPaJvs/FMoKABjFm6ev9Sla2IYngi4I6pHUiK
ipdGPZNarSdrI1HMOD8hnZgXx/ofUoqi9EfrYQyd7P57O8V5j56HwmsQY44Y
Lo8Nqp4jSP2YVekZExwkeGdPQGTC/O/azJSnU8vcbrMXCi1Rw8NQ4zYh2ST0
Sd/Q8oALhUAgwvZpy7wQxst1nIxYL8E93zsBVWcf0jFf+l1KW2PbamGqFB5i
/FfupdCV3YWRddQTZN7qo7MFWGUkhl8SuByTHR+CO6Uym0w9TtF6U22tcIEf
Cac8px7+alkdfuIKWbzdTto+vtRNLjq43Qnw7wNOfxYx0nDg+Uz1e+x7qJuK
+QKatmkjS0nPnz4VUpUb252PxB1nqumYVcZCDdRjWkT+iDSFrOKBlxtxX2hY
NJ8Vxg+wqGzhonGlbwt6yYS6cBacSedxhslrGlaMLgCVrJKhMEE9UOfLhQlu
kU5BF6M2AgOlayVxATvnrrmqIR3x13VaDJyabiXA8rt9AT6jp2EYSOwhVhj/
8IWjyEIz5wi5RMjkiBNhqsmjpHTSzHeEflWTLB4UiANtU0lWuJ0CGDuWO43p
Wf+a6qRJlh0hbHJix5k2wbsrr5ToJI7RPHICmga2HGMNLDoqyMaxJ8Eu8SCi
NfuSeWuKqzab4CtEOAnvAKnl6hcNgzsEgakxRxTZSi4Su0BPIKwidIJ+HuyT
DpjR7ahs2n1j3KsE6gaFe0pbwdTqyOvpQtM+/8zj2S+kyRqo7D8rFWjVrkCN
0MDINra4waH2XnbFGBwHK4o3KL9gFzcINBYPOb5L2tKvGgxQo9tCf4NfuM0A
KQm34QpOFfJPzuDGEErNEGdiOFKVRxfkWdRZQIQY2tWfIuMN+ffgW818fOy5
oiZP0QYCnfCVjcIx86h9shgtFhjneVy+81/QgkdczEwVEYy/UJ1ntnBaXg8J
BPw4wx6fvT8Rm6Ilw/fkqNvp0n/JLRC+TpadheZZWXJsWOo64TYcEfZdvqdw
CQbpuHIky0izpq6AHbZ3+LbK0NoM6RcKfAn6bDKrUvjhoRu7UHfII486N0AZ
9nhuKCCh74DyGTiIMnUqfrJT79J8KgqqEMM3d9bpGjDRVx9V6WJ70cCoSmDc
Rcm8hAuopHv8VM/vQsFzSwcL6m9bx5JPsGjSlHHcdQCNHxyIlRQP0snpn+cr
3SugZ2+/ZaQGn1J5cgG5c3BLggOC3WmbFFC1vJIKCFMbt+LDoXtk/qLQwyh+
tKGjmJFqFHZ7Jej56dobxQhad0cxo3nd16xZKAo0kI20t7fUyQCDLOZYK9fF
OqMkQ+qwKrlI01RQ2GsG1NcBejrAv68B4AGsu8MDl4XKVH2kcQUr7+g9V5Lf
uBv7u8nDMYqRbWIivRJikIUT2n3udJ46qfStQ+Z0AyfCeYY/VcN7BuiiFmBv
HIcwFDoYuIdm7zKGs6Bfvm88IKrrTFzO25YA2SRyhMxAVJCr57Mr69I2YPCb
5geDegl/WqCwI3nsxyZMY3rH0j0CJ3Mm0rMMwkkml370j+nlvJSzUy8vxHd8
lwm1xYy0RwkoTxFEgVTYrUW7UG6wHjgqiZ6mup4pK59Wi/OPSJnXQPvvnOy0
Zz3PisHCu+/Zfw3hV0VKDg+eK9fDGzZtlbA/wB7HbOknucTTGsVBNN4dre/o
qpvoOJ5g7C+1R8/7MAkUOtf5u8/5iR4z16j+LeRM9z8xIP6iuo1d8HUhJs41
B64eqKzzgEALmA9YKudd6LmK0QQ2Aq9eDBG5NMkn2+0dIqa6pkUpN7s/R/eE
S2uBWPJX0Lp/x8Sw5yJ4t9NqtJAPFlkF7pe32lIDYgsgycC2kAsxCJNcDSvM
xUM9boJkzt2+AtRWlUZfgLNyhnk1WZmJU97zvEQ6kaPnIeWB1Pj32FUy7v7K
ET717Ls7i85FGYFLOaO89H+LMuIFjzy5m+XbPKpk7kvVQDOwa+AxxLRyER8U
RdFwt//uOgt/+z1bHoQRA1eagIstVYGjsJUiJn4mixW+3szeQUwF59V4qzER
O9yAKalZqdq7DgH8QkDGKX3hwyEH/1tfVn0o+jbSf4OyT+jJt5jz5FT5icVE
HGC0GLq045XY01jI901/KrjlfT0oF62Nd7LPrmgU+LltushlWYi1gRGyBg1V
jZHippJ3rmwW7slBKR8xyYUfsd93qcJ26tnCVdvKDFe5NKkWUJCuBp5nic6y
SRXdJmdH9oc9t8yL/AOhlKIFO1yMe7CQfXT0WiPRHFSAgqwyUDV9Klk5WK8n
qFoq58OokobG50N8QzT3pfiwICYMcX0E6ZBiz6EG8ypIsf9+ba6LgzcY9Wec
uHHxNWc/46WLQlUOQI1/p6YknYKhpvAWeNukTbqZq/QsdLiazGeYJhjunWWl
DG1RMrMPpmgi1LTOtgZSThESfbgzYQxAGlcehfWpbscl+i5uCvPl5GPBEZB8
mh9dg9u095W05r+CBHy3GdtNmxtI6JmO4CZ/8MECsGFOsJZKiC7ruPuM+q5w
OnrNGLdA2kHGP9UbIVdUICoGHc3AvxuD5wVSDXnw30NGn+pQ3VCUqcaIMHh9
qflZVox/LiNmXhs81u+DbxYqSKVBYjifS0RkYSIiHJjZ+Xw1aEI+Qy97zTNg
zQ/2bz13kFe8CyjqKmNjDvprJ4w1tZOUeQ/R2Rl2RPk5zRzeYtK5P77kFzaJ
kuGEH2SyDZgUCvP79ruVLqqtp4KbufTtrvpbllcCw/6EWMimlE9zI3HHnKuP
6HDFfrCtKeBudouNUPjYOCAQSxWWm3HXexrhKjB53IS8dj8lmUseOR6ubWQX
8s6EvbN7GwNWv/X5mGeRc91DTrHF83dmvBHzREUyLhJAwwjfPJhff+V652G9
eYcUHPnPbIWssY6j/ZfuGuGBmvvbOVSv2ewKypfc1UvrbhlPiTpmhNChVdw0
T8boFtUmvrPnx8I6OaPKMrzc8Bu1rMcb0VZpXd6NxAoDk7endp2E+eH+jTTj
6qc5C+/+AUEhbFLKSRegg50w/Uml9bqGnedn/sNkAbAgbyf79i+c7/HgPnBR
rnyOAomswFQESZIjIK2nqjGFkv+HpwO/qBt2YQd/47K6ffb8X64v29Av59xN
dsWPIJ299ZPG/aX4q4w5jZT+QIr8xYkg9GD60tRFGhknxDGWRdcn3Zyr+ljY
bVWLdJoUmFpadETUVlUr9+6cAsZ9FvkK/pHXZZZ32AwYC5dgw8Z7ZMkuWJuq
54uyA4PLDVkOMX/tXbW/6rzcDsniWf88rVKdpMaxUHVNH0YfdQGBPyE6IFqI
+WqnJM7cZy1H2997ShLCivtsX3Xll5jn+laawpZzzHCTyl+6p53NELzhbLVp
RbjNBaP+a5qRRruIBg42f6BGWNJwbmYFNikNucnauDe0ZDDLFxyoKYaP8guV
kzckYuyJFZ3DJkQGrZsx1+JIo1ho7ofbmivXWefyJVJ3KGRuYEQyXA00rReX
v1uTOwtLx2Wmzl6e4hBbkO35K2/okGb9NyEnOgJ/I9eg4oqKCZmUdnLLMVJh
hJYp4HMQT7Sx+vtNpsxRX6F8V22cINU4IJJWaGc0c+ky/logxNBCBff7WHQ8
AhHrY4qi1aimOWIHqG2UQSmdtAiOYPFy2ZuLV/SFW/r7K9emRllB4nJ2jpLf
Ty16OF2y/S3+gcvxAQE5qIzK/LB0exh6BLr1dSQFCMfi6gW+w8rewGBrirrV
Na2GzQbVq19tzjQWz7VF/mq2TLNRx12bP+0iY6OVOyCYDhjPN34jHH/fqkn6
Np2Te2va/SHlXVDzXc+Q6LMZINpPfFmzA2W3gEYH5tjlf7ZOYHD7z1Ist8Tj
Kii42XG4w71272j0YRcFEgFAFglaq+i100FBaq55Rv+SL4EB7oQ+5gLHjQOX
JXXz0lGdXr4fnXD47p3NIcHTw+JRykGN1xC7lFAtCM6TKh3SYCM2tHJcaqtd
iZJqtZFBrAqplhMQlDcknmhxhIJavDuGqsu1+hIihTfe59kjtuVlIAMGUZvx
7A7rTKIiKcy3h3IN3EGuZod19J4DZ+J0c2fWYN5MbexWy0Debfzh4Q3ZhDj4
QP99KWpq8eJZ2PXSDkjjuF839a/Er+iMsxy84GtYyz9PZA2JXY4G9/YtM37N
fNTJQeXMAdGqsvM2lzNNanpZJco/dyQj0dGPLshBoU9SeLwayVwRCMMPLQxs
6pHi+daGfG1p2GXDbaOua+GR9a3rPkYetxHCF3M8f983fYE+UyG0gkMYHtVn
KQ+TWNU7xWsKI8xNFP0BJR7ZVzv85UiHJh7aR6oDxIVKI0dyYrAtqDmHrZQ8
Ju/SfimcFfxbloCSMMW7hAexsVcM/BWin+kUAI7t2lEc3ak86zHmmceg997q
T2Q7iGX6DLRz1jax/FFejWWdIZflV7m5bzVWXRvUFZR4Kh/3QnFbc/7Q+VK9
abFELrrSQ5ln2EjwAW8dlIFi10eMvCWYHi0Xr4+5A8IwPoaSqGQT43c5eSvM
2bQM9BpTdtpAXY2TzEXzGFtNQ9HL12ihGkQAh2g71VI6SmYnIOMyxrkRNb9h
h9QGPVwgaRJrDYxObhPqXkDkxYk+tsN7YDxOAL2k8scSy5qa4cgeTpENjMkg
gottUnrD1yHr2WlH77YIUGFNBUBKN5n+dDkiQq3Alo1rcUo8DvQz1+DuHSfv
Ukhk9ICMpYRE9VaG/Ek2QS9KtMRYGrALUIVRtB3RvMKA8KnvHgQXrWNxAz6f
avpYCXVNW8cPc6lwHQVjmAHXVg8IrkyiGet6yziFTnP5sxRqo/1Btf/F4eb/
vBOP+u8qRTOlVbTchMvcVT/byOTs9zGt3gLi+jT4g954X71P/QA1lt+yIiKo
+zm6fAAaZR8V2Jyb1luTD4c+lVBLwC0Yy486H+QVZ9LNX6sdpJhmyt8saQPP
Hezh+BMAKWkG/2hZsizDziTKxCpArGX1ZKB1Rb6tsrJ2AwTsysZfMHXKGN1f
673LErXCbkFUDBkA15W7I5CuvS34IKbbfzzzVckCnFsM66cQ43jdRlsN/1L+
t1JDBVXt3UKsOh1yQ7T6JTaDpZO0sIHL1LDj+NQai4QjdC95KGyJadiAZZFn
QDB6KnSV4Leb93tckaQpwQBI1DJFqXLLy6BpI0Ab38AtmxI0MMfgASei5DP5
jZY9F/Q+wp2e6Q6YhjOCNe+rem4d98YkhxdeccTsxUIKsVgF7jLlblCHNzI5
MwfvTl3TW72fatL+msxhdYXnj26U0k4PyCpELNyk1ouWgXt9adpVSuGeY7s8
F26TrSMS/sqSt/Z0ZsO8PnCn8EMtg7XUhx8GRdHz1jSfw6hT6ehMPJmtkC7a
JQ47q9TsFbaPUV1U2kr2eMej2FUY+cpgJeH2qV/AEGrOTjuvNNj2hUluEQt8
iZEZ2PfbPhVN3jPVe/v/W72JVr0w060IoxGvyKSe4xHz3ExfM7M+xcQ2miEp
SSAfR8UKvuIwCF9ZrFYHbT2uGs+7e1NRUZSA1jepXON8h4yvigNFWNDrgzVn
R+rt7UWJ4mDmBJS4Zz775nqClFEKYj2reIV+6z4RBe1AtSTxjmQjOEk2AmE8
TZntqhmQpV6oGWRe5gshh5r7VMFqRfubGqK0PhuV9d9yU8pbrAPDPSAKn8UI
DNxU8dKvTS2rWdcw6bvf1WlCdzJymjMrGQLdRu/icgshx6cJFuv3K74Ijbwx
TekVnTyiyWvzcy55yMITl8Gk3q+YZFpojKPHlcxc2s8bJnwqtkWMyPD1qfWI
Ff+IhlUVYmD0OQTSzeRs+W9FaAAeIepS6TCIynUI1zq6mH8oOTni38By9ObH
UVNdBjIH90A+ZS8VanaIVCQKCLpNAHLlVYA0IPGP/SpeTZRwd/NoHZLpbFYE
/RFqMzTNEF62S0E65blhZ9NocWVsER8tovkk0DH49EYYPHMxX6mcssrWc1cj
SoeFYGwCK8RjKaExq7W9vjBIbsi4zSTToRfBhVF79+lg91pcQuLmgjNClzeB
TLs+n1tiUhFJU0T4XswSsi3w7sIBBf+W3m1i9PVXcFb7cFZcWMWZlNeP3kv/
Dkq147Y+/T/SKzbeIZAOikHiUS786BGmeiw4mKFuoa8OQXGqxoaWODoFGtk6
EQxMzo2VvsGq002jBlTfBsf9SJHrRUojQrzIp+TlNoRBkM0KWHEt3v0AvMmT
0EIg5GTR2c7+n1PFx+lckBl1VkWEfMUkMQe5LE9cf9Z2mwe5KbJvlwBiy89J
XpyRhzidn1AZAiW+ejgbNrMbJw9xSqpcmfYnLU06kKHyDgoroRTHbjIo1BMp
i6RqEoXmHXl5gNiVqrButcXy4pcivNzsB7QTVtpa/1FLfGWsHxOJKZ77GwZR
P8yYxHjE9xMABjnSjKu+ObFzlS7foxqL/KgGhPrG3X1AqbBjFoZP3xa2vLIg
6xmSHCHn2pz2RCbAq7exVbdX8p8cc3l0MKT3O61oanu8cE3lnOUkKtx4SbOY
+EFXOK16TuWsgMPj+R/8iBqV7dYIWreeUOMptJ2YxoccdGIxnbQQUtQGzeNM
GxDoC2ekXA9FMS5bGox6QDxYuhCwZ2pPSqXTq36CMVCEq/6sY44IivS/3K0v
+lzZvnW75VlekK20N2jVhlyXIebg4H2fXSnZkDOm0meKyHuw/XBXIzGIuE1e
ybVfJ48tQGUgJjJ/hTJCgWBTXLg6F4QC4SxZ12tsw6nylPGuW2FSieGZPcFf
d/5hSo//58af1ADP/my8aJ97ymZa/DXKHudFkcxzcTaLsHMS7k4Z3CnI5C1X
f1+p+GjuhOPiAwR64X9HCFb0znsX7EZaJR0bOY3IOusTIMjBfBGlums3gGBX
kZv2qPADYx+j5O92jEd1aPCKtlbFqBGX6dQQtdon0uYn00pgALHxEbL/8spI
ck00+TsimiALTqawGRAEXwNCjAAa3HNrEeNiBPwB/KD9Dn7GCOCOGKvd/gPV
PvfxdEQ7pyn3UEMTmtNMirZkaXahLOeLY8fPoNtHBpKzPL+vw/xgYx5yl4iq
TdG630583f61/L4QIwG6di/elMSijmbrcUpp0hHYSc/dtHY36G8UwJMXTYUY
Dw8BQDiQlSEfgCTwiCUWycMg2tIJQamcVuvVSg7RFvAczaKN7oezX4ShHKWL
RBOlarAH/oV1Dlicpz64q22DM8N+ZRD/wNRTeXkCbqDQAsmzzPrL5S8Piq7p
Py9B2nKNfglS7XDQuxLzV2AZTljxV5qdO6xSmmk0VvXoCdiqzMSg8i3RQr3h
qo/3pvXtMNAWaUH32/bDisgZbTQetBHStr6LUXBYIAARiZ31aFtNvyZbZClD
Ys1biA7B0H2lK1rXZg3Sr0zElT61Dat5fMCRkDxCo2yW7YUGW461LZ4kGVGn
VEkCKLVJqJP3NoGXdV2gM2XdYmPi3eCDCCiBuOU6In6kuG2/IZ3rlnk/IpVn
6czhl62c2rCbquxxwUZ2G8HM72Vy6cV0/idZUHFxGYGGDQEozu5LJy6qH3Io
pN30gs62mkgYl1piehldKgrpjWD9uKXngIC613jMu9QbZHFQwcR69J0yNMDA
5xU/C5VZkBGplTZeMdIXLMWyqqoPD72ioROQPPQHFm/IYjTkBidUA+Zdk4f/
wdk4k9+s/XOVy+c5u3rJw4HbQvnOzSUkYT1IySQoED/05FZvSR1RZG16XZzw
f0MTfaRdNPhEMUup2/83zN1N5MdoMPj2N/buFT2YcWpqOhJO94siRZ4h8Olv
HJS79puvykv6l74qKo9K74MMWEdjqUghP//3jJDg5L9Twmt3tOlxBkCUU5P4
lzo0m6WWJQzmC5qFm7G1+YRZ297pSkjo4L7LdU8LxqtFmIY+9cPkukH3O03L
tT0x/AU02kxFt2/Ajs93hfGPJYsuVnCzcYXqJYea7mecO2tIDQOaIdwZlDLm
56bJ3qaUTseBeKPp8eDiCP0fCHrrTXz9FJqToQRzEHiUG/8Du2tfrncN5esy
x/PVYng5soVRy1ep03enB1ujHBJ8eyQ7vkWTPzRxSWbmGGGf4u7MHGoUd5/F
xlUubs2ZNKzJqjwukdkAk+oEk4UGUkm5NjaqXaH+NJgxVAH4/a1fYt2JZRm7
MyZlBXDGAzf1e1eHKLZnPeajtUlPR+ib6A+PqyfnIxnQKyjQXfoGnrf8AHV1
RlpqLpXCX7m1fCDo9Y6greMN0EDvb/feJwot+Lo5EHe7vtJs1FqwFgX4NL7V
wEfUg9JfL3Zhyt5ZZHpsEsXSSYas/T9ZScjWU30bIikKZ3nvY5YnCMuO8U54
DtssN+IC5mrhUP25bbp289zsG6kPr7nj5JbfiNGYSLfQS0/8p+c7uS+Wqw94
vjPct4ZNKsR1e82O6eG0uhpU7oEJbUZ4hFe1OH64wXgufM++4Fjuqv4h5O8x
tJlI0XIafLcz2XNBkaLI+RwhM7bJkvGuwTk4TRh6sFBpEDKTQ6JPgJBw1seA
2peAU9aabvMSg1V8GKYgYGPVO/jtdEKYjmhaHV5cV+IOvRfMrJ16pL4IdJqC
ultrVOCEefepDuJtgR7SOmNlVUXv7MdoMqiEl98/BLCu0UjvNvgDkuWyfykD
U56L4cUs1sFt2/b1wK7vVm2Nd8jD+YbnfqF3EKHSX09qhsg/uwwHTefV0A31
zukBEH0Nn487rSo29I8KPjuoWdeBUTa8y1xOvoRHYUfe467FVZ49wuN3dHn6
gxAgX+xx4e3bBZ7q3A2jqmiE9/oOek3U7mjRvU68JzRixW7TeoCLS9amTuoQ
6xxKjcvBqk2GkOFB3qAmqLbyljInKsgx0djgJlvJ6Thb/nOSA09ld68WVvQ4
+PLlvgfNcAtT2/Pg4SqyThcyxRAE5sXtkCXMDtTAhqspH6RbFpv28MJP3mhe
b8h95pwvjvOR8bh1aVDcTwyyCTqaSJJYJ7Kfj+HKFIvmQfKXKkdywDy63rgb
fBAb+iG4hAHJJ8CBLSLZmvwdMi+xzyWt8GGyz8GIWuLZCbjXR0ra04wwnNQo
eYwGMz/dXiJckb/trzNN0MlUBZzgE5Y9PndXUpqg/jkT3XLwuR5g2vLYvYzF
f5EyqmZyX6sk9F73HkVHHn7mHR659MRC4Z4Y4k2Ppg3LCFgDbvfd4o6ItTZn
mqBwX06rzIMIbSp1yb88wye+B3JkkGl3Nxtmx+sftI5i/u8ruevWCghVBkVC
qK0AELhpAsIur8aHFgqwPhm4g+eiLaCp6Jr9bfSzIIGHYEjKUYg8BhI0KP/o
c1wPZexWcA2LBXK3Jwg/+dQaq5oKxJp7WO3DbGhx17G4eQfK4dSwNMZH0Zv4
sQdLNPAUqUEeURsyO5ej4E5H6VR9PrIHsmylX6SfZ/Ej+Ll9i+pA4fsAgGmH
L4CTh4i/GfZHobd4y822zKUhhkB2K4dFlICNaqUmvTkGAPS0or7wZWldKgc1
sNlQCiauSQ4OAwyp1qQaPv0kLZlVRKEAwxLkvNZek895u2+4Yg8lCwa2p0SG
H8edJTs0MXqhbfiZxUatqHgRKtD4cptfhCIseOjMLdxaGoBwWhh0OjG71uBG
bQDLZeS7lfAug9kl5pbQVGQV7Sk5bap2c7uTWyFOZOrjrrzA0VwdxxAuv/w8
gjTfgifJZYA68JdjixSqAY+tHnWI/FGrOHJMTJMGmMqe3UserVFFUheyDguO
ajKJUFBEsNr20+UqU77tHBNgWk8n3C/VNj+yIMdmTmW2bk5dywNbkT+gr5WJ
maMAUueq9p+xRMMjo+6YUg5pbJqdEHVPIloRzrwQFC5UjhNl2eSCQB8f0+al
VNVaAXtPIWBe6kIEI/hDB8h/G9hO7Tstw6uuPNG/z8UN4SPXzyjAhZ0D5AYj
RTqhe98WImxKhYVQDIMfH14mn+/MsaaMhK0c63KWk9qX7qumQMictiGHvMLd
Z2hv4NFxtYhaFcMKN0jWAHf28LfsLWWUYiSLzi0fJjsLebvLJtZCX5kvGP+I
OU3R1ctDB2djEOejsaqbgCKy2AbCxXoq4vGNdqzMc6jYgFVdW6grz9bFJIRB
kc823ld0Lm5HRb5mD28q5jDr+zwy3JIoZmUf/O0bS4j0xkqmX7CtmvfnFcEs
lh69mzPm0jvM+V0M2332mbiADZwQF+OxkBNf3+TulWPbLKWH3z2xlBjIaT4W
dTXylJ/AKOlzOZHhJw0291gD7rluz7dTVv6/c2EN3yTuPBEg9BpZa0vfyFUq
0TSQ6qGGQRN+WPT0q789I6R7gGxe4O/Tljri2MpmVgXNLimaApyrq3k2Z19I
eJPsqUGcfzh+wZHMsLcn+Vz4r0vlhmkTFiM1esUdKUfZ/wq7SHpoVnLElIll
v1MOuA9mprog27zwruwkUtp9f76X7is7dUUmuErjFBVePY5BaMlyB7XECSEb
EuXygoI0mkw/n+rFOpPMYKSNT1jFErV0BBXQjAwY/Vu1hxA/V4wEApUw/TNR
R/QHlOOyNXzwO5bnqn47ifKVgLzK/7k+g2U6nvyj4Gbp4DwFpnePG7lqQ8OO
nfGrw0fZHAwrPHaSJOnlXkIF9gi2pX/uKCsju8lk0CMV3PyemONbqvJRWbWx
ESQ8aHBYUoFiqnaqQZbnIxHdh6AJ/6NRg8laCmHwgM6LHDu6lL6y1wHoT3va
qkP+Hvp9DCx2tmFaQghOez5CL59SRlcQukUydH/ySFhBUg3jFZubi2ibEeqi
Hens9J7S5j/Gkur4XNHOVMg5BEyaJVlJqup5vqTi359YmU11RjvNMjKpJlrp
dZ2fFHmzYo5aHMaI3olpoKpubZ33ECmAwZ2fvwzCS9sC9NiGEUE+dSydcJxn
SEzCYVqtoZWxxOzxq88pk3iyRgQTGlSwWpLLHLLP9hOxSR35YRRDOsuXloti
fuXeo/rUSnAftU2ts94YxNk6nA0okAZ8j1Mc9aCa4S9RWrGpNuxINv+b4Upx
jTBxG9258TAzoG71QmuKEMuJ2Lem0EdoO1ILmfHv5naV5+qfVQKUT/f5+Era
wSriQxiDQaVCwV3h4wtgRkBxzw6C9oAKlNxAR6yiSLiUZy0cUVpB88//odhq
ff09ePU47GhiPcIfs829tnPiTNcCUf6dafw7eqluVFykKC+Jy1hbz3dv8hjl
HQ5N5CcI5zJc7m0M8eIsA7WGIePbCJO7q1YISfecqKFCSC6rs47MnUq18UIx
MHknWz1ob4GvtRPbO7BRkHuA5PEL+VfnHjaT12Bvp63gx+9vsE9FrS7bxHWu
hk8MQGhH+fwNyBhPMnRZLzmJdzug3DgYL63XegQIbM73GRTWPbp7FLSiYcSo
R+XVxon7Q1xnzOnzi76+pRSReUsnrFy0ihZid0VMjkgO9JAJURZNPqiEI98P
GN+jRd+TKY3qExZQg5r0y4jCMYGhAWvUlbLrZpXmbWdcvSX8E5sxXKFalzfc
7ytjtY6eJrYhdNU+04grHajoOlQafBxdwbAC1GR+15WgLix9tJjwuTca1hGS
emks/dEXgDyCcW01WWaS4Kxl4Gm3DbF9WchUBIaDCrkQmXtC06MgOt/gckQi
ACmZn8GZhtCzwisC1wuhRMXaF3xG+/WpeM6w7/3LFfL0elyd1KLKV1uq1BnI
FJRksc9NJQL1ocnaVzXvyqoUD8PREvLYOLO+HuzeQnaKUYr8CqQm0ueP4R3K
az9h85bRYivW8Am9+qjlj/WTp+cypQHMvMyuyrhlX2oMOeygk2q2fEku1wTu
dklaqh49FNGmJoNOEUd3K21NyT6YvW8wTFjCc736p2/BuicfzH8nzWtdimwD
s1SMjKh1vLfeNRi+TSe+CR4Tesu2F0tXnEX1DdCJtjbfPapWZs//9NAHKBBN
HaqkDSTEONBcUFeomOUT0S9nfzJ2a0K9YGu4WZRtwtLdIssIlC2NPRnyOH/M
LY4RuRCtFfYNVYTF4umVHayCRLkazWkZ//qlexUbn4zwMAJxuadWsC2mvLVE
14/ZCpNQbt0wEyYgpdWXtTwwc/KdMwmDcyZ+DpiuwuoDboAmMr3sUkWciCdu
/hB/vGPCkf4GZ92Rc+OL+RWzWF1Nl8vGZ1WPxXZRDRpL1OHPLDmE17ROTKBP
iotGGZj4UKhqrvNHnvSlddOsKg4DxtsH9RsOq3kPWN/N68vhmiTlz35DKidt
WG1koc/6uo/akOZcNa6qPlUN7VJ69N9wAuL2r3mXd10Fe8meOi8lDyRkEbTk
6YasC3Ku8Hni+U5xU2CsYw/TyzGf7nR5m7UCm152h6ni9+HhE+cwTdlxNIZJ
uhFFE42UPCb3NrBG2yMfLhLjHVbRYky6UL8vrsLx2KTdWf5KBoSj+EUDqiZ6
eH3JXXMhgj0PEWBFKqlW4sp8GWsSMX4e8kcWHR6GHdywFv1i+6LZwjQLE53q
CPTMYmzW5U67snrggx4qr7RlZlhIGAOWpopv+zPh1dltYb1LvoKEkiTRKtBw
xVokGmdEexSKd6JghAjRwN4eaT3EkSEpIlu/ZDKe60vDEvXrPiMtk9HmtmUu
msUpV66HHD8juIjvmyTnX/lAXJgRXzSpiKfYTBkRKlLeSkeuSeheJmE9mQBt
BjYjnYKKdFmcN4K7Lgm7tftSVsGuuANbUWFIabyW+l+HuHG3DFKg9noRGj04
jefBRrGVlQ02T/JTwNBwSySWqXjSpedxqaH1xlV9W56TJLKAtP0iFSoV9zmR
grCw5hjkVcG9ZtO/aPTjVALEmZY4Id6ABLezqlMtPjknl87OzLDEzdeWx0kA
9y6Wuy4+Wpy8+QJTcwkV0is863/p+qoy+l2YZyybEoLvcbHff/WMulOBgpda
DaxTySAoOG1O7hOzux/mK8BRJt4nnBJOgvr1DYqLfaas66cBsikCaG5tNYDc
CBXfGEABbWaSXXNc2SuO9y9g2T4NbYjMUCwnYdv09yuMT9qzEVUKl359ffS8
QucLRBXKH3eBmC5KKUBjP3FDCYVoTSjNxqWTxSuIvpTgVZd7yOo27/MG8TAo
sGIaevJ3qSQe+UOIZVcdTet706Up4m7RYFR9B3rVrCqqsPytypZTXf5wnMhN
RgC+4kjdHYSLyMfiNzVtZ0Ig5sz8eDbWUaJirwNy58RbMZJZcjuQW3deRTCN
ZMRzCUpO32Yj4SDAX5Xom5fiDaxujEKbZA1FRbM87wlBc+aBGt2f9l8DVOne
1eTRJ1JMv/tIzHBtg7lU+bFnJQ+J9+BdkFCk+rxq6r2D5hT6rQmj+KurBlS/
YzOo6GVtDxM/SI1VEcHH0zuJoih95/wHgCRnjq45nNb7RxuJEqLY79jGsRIt
lrUVMRNg4z3LqJobLbU44qeEh/nK722x/v5Uek10mw8uHVguKk2DcT58SgOj
OmTidCOliAKiFumHqdDs/4k2zG87JaiHQh7zoCUBFnPwdFF0E9lvrCt7E+cE
4UhvtDP+s6haTinpUcAHFGnmpgyJuVRc7CToXHlbPvfTSS9M/KgdIvpeKezF
r70LeAz5tjCzfkpgFbBQCalrK3iVw+FNRfh3hHT/7I9kEVQdO1LbGiGdEjap
uJWb5xqnoxw4K+JMWEmbbmcucYUSGAg5Gs4tFTF3eoDsTmYyw7mMAvA4hALT
A0bwo0r1UsGwvhyp7FvFBzZ02bvgmAoJSlnZ9KDw7lMDicE928IQukJ4mcM6
hcS+7WcNSlJ1xtilm/ZyOP6OyHbyIPqhw1rhSdO8SteRAg1xPgqplwvWb6B+
vAKKXIZ0Aa6R7Hj1LRcrk73TMc0qCQXb7AxRd6ObzW9TQyh3KXSt46nXJkCh
uq0L1q0SHhlmX2R3gc8/Hec7iW9oPMq4TpyF6duCg9qJzqs97Z1aYZU49rHc
qgOfDyi9NH0QGZ15M4Cl9YFpm0WnTGR6AbhIQ1jfSumoh8mZkoxl8k3zdChj
foOm0BV9DBdAyWrWaeZKup5CjVgEh1Vxo3B7YFBWXMYZD1kYjAFyXGeSD8XU
U48jyfYNVgojhFSpgm1FbtLOxCJqvb8DU9JayZkDIKepJYQtfvGEVfLC/YSK
0UKMYdvS7INjXQ7PMwWPOZq0wUrmMJTz+jc4l3+/249GYPF8Pn2HAVeQ9x+l
sXc9sZr55N7TFquVQh5x93Ldy+aUQ+ADPUo29VR8bq6fSQtQxfgHEukgvENu
yOiehtjjnh05SyPJU7DE1nlWyj4MPT31CcAcRkjyvUuHN0vKRdRfeGBLERru
Mw+MF2TQ3oKQXQLDxQYKjxfyOCc6cRSwyYe3sw4aYOBCrvFMrnojajwbeh9e
9blNB+uJiUlXBwYX+zE5J8TALHb2cXbMh+39r9sSfHo1bpnNHvTFwlAw+6Q2
19OVKZyYMHofQFVQRV2hvs6B2pV0hvsdXnTQP+nHHcDNl2TMGMNrMFL9o/Qo
GmSXpVMdee1zP17Zc3if0kr6+sKpnGh1GvYanX/CbpF3DRPkjFIEeMGhs8wk
yL3hgj6zwoyaDUZ9sZC7aIdyG7P6ZvIVcX7DarL2/o2T/xe+hdYQyQ5HciLy
qJ+6iWa1svrFccC0+pQ8CQlWM0K++URUw745JSLcJl2oeFd+muCFki7z/zk9
WS77cWgwEhVITFbO9DdMXhATfXLZ4+10jMpVgYNij8ePmv5L072hgj9iYJbV
KKfJPzcf8lK06o7f29DW7mRpOkMOasu2RBxQL/duuOcgd/AavZKDGtFPSvQC
vhZ8Gl0oc8+tyWSgUlzPi3rc92YoJFdRyoPp7Kls0zM8yA/2egBDGclRMgrj
gzPZaY7jGrJA36hQgcKkMEJy3nH8u0tHWk9cG9HcO2sBmbwK4jr0z8WT0udz
FtqjNkC4kDS1ubgwYPaPRR0zSYZ0VbkarIh2eXVAoORP5S3XTgQFK3R7Z8Br
mb4EgrBrhqFjdG6xIvo5BB02qHvZBLh9ljmY7ZOo6VISS4nH3Z1XfAn/F5Kp
fWI+D8Uq7ZUFOcnfzeTA6vwCtD98/gh6fYnkDopzDipmHfQFB2OMtgK5mA95
aZFLXxhLtf83wWcdWaBRprZQjLDcbW6Tnoq6Fyk2QqRu/f0wSy/XNg7oHBWa
8lp5mgXpXWZ0cEmEhE0in4XqO0pcrLPkhOOkEC5iJIJeojPmIvPRaskolvSP
GB7dHJD0CDaD0R5huRAhG+KHRSgZFQ7XDDzaIhXU68yfzshQ1zchdVtot1uu
TSLWjdjy4/I3alKHcJHNFOfbnuf/VADU18DONxEMNAkORHzCOFBT6AdQXHIF
PX1R+RNk4QA/KH6hCjWlJVN+bV9aiEd+W17SDHQitYSBnJDX7NTqDWLDSRdh
mI7d0czLz3k8rytiUeC0BD6h44F2vdFpVVU7TT77N2v2sKofczUyak7uUyyt
Mvv2rR5zm3uotIOhEs8BMdxObUgenVJye87zzQeUxdN3n23FdlCDh6m8Fzi0
ICcLlHHBBM+OcQ8Uydbzg97YtXTzqvxMt8O8U0y8fizDD4joJ7Co+jrYAs3x
pasumDVDepC0O69Zn5vCqsGPsLGrnYiqnWs+c/YLZqz0ttuPAhc3USBSntyl
HBv5R6p6Ce6PRDY3+/iP3nISLC42+m5AYrkM483QuNUfi6YU6SETfkhMjYoG
+TQZVjPfU6t/yCNQLnArFi3Tr13jvfKYH1DGOVXB1EEKQ1NFExQknD+PI0jO
fUZGvRfbMO461umbf1P9pcdEhw6fPkpAcns0uC1f93e1ipA58gKAkcbpnmmK
Dw1iQF8MBo+hDJHo1+Yiduk9Ow9m+CyLxJ1NF/Ds1h4YNamPmWWnN4eyfaFm
uHMvc8pedQ1HyGxLU9c5w3MO5cSPm5Dfmx+G7FItnju/8jpxCCJ39W8+WNwU
O4iN+LwbZI84HVN/oRIb47w476PbSzuDuBJ0EYqVeTE0dmdQzwLOux7D6T+o
kd0gMU6kYqjBM3axIfll4sOKO1HMC5gIV0m8ytp69SgB8A0X31PidOPG8yMV
OS9mFDh0AHdCUaPb7f+LmBOFMoU7R6iBl+87AlyUZRXCyaeAwXrIhjNhXoW9
rFaecWT62hX8B8/vZFXv1pvxy6+znTCxBnJ/jdQY1+y726XdbxdS88TxPA4H
bXHmjfT2w6X0NAolys3RZMnMOzRm/HytQjsa/5qDwScKF2vUbNX5bvcscRJZ
BoAsKEGfkqvAdQ98ofu6Wn/KvlyoB9j4dyxeSAiBtZnxX4ou5orf6wSgFjWO
vKY3swtZESHtZsNggDtMFkfoPU/rXEj+CbF0Wa7d1QAdUpQk+r1tGc34NC7Q
+66J6Mp917PPaE1eY5otfbU/F2izUAuqTX3uQZN6cn0ARjkK8r9BEFAuKnb3
Kj1gHhLYMOWyWzsM8bYAUSqcZfLG9iBF+bm/tbDeC9KxhG8jvDBUglYpPpup
BK0DwqSzueXukFJaMpuR/+MXIBrC3eGmR7BKBCf/cLubBR6VoLqI4tFbUiIx
MFJYrtoDSMrhtNpVLMMAat86niiCdS4X27GA1plX+tLrP/BajKJ6gXtlct4r
7EmL+4X87yeBIIlPsYgl0CJfTacyRy9rY7+Z0c0nG7Bql0DNcFlxn4jnaQwc
I9Nju7a6zdKEiBIQGK+1xbni9uBYsyGxSv4zFRyz7kfSeIB3K9fkB2mwySou
Sh3tdn60dfkRSYR72DBeg192UVtEGHz21AUa8cZA3oqSrVo8i/tghgr0Urdj
2bpkcE7YMEmJchAMqr2Kefyedgojg9vynoqXGX6IMO1JJ0KL5VIxmyNNbDGH
VxZ4k0GfrVsdnIuIM/QUdxpbFx6WXGVcX5RR+vSNyfExDeDe0g4K8jf++Hol
4MpIX5LoXdmMv4JVEnrO3AKgxqatnaZf/PXFBb8mw6t1cOkbPgCs+YtU9UjM
cbqMrWA+slLIW6Go2PwfrlfwZ9vUOVO02CruPvcQrjckQy/kJYFBFYQXJAU4
ALnYusTwu3+uch13Zgg7vXyblOXIeB0QRENmulod5rxPQkpjss2X9jeZomh3
pCVW91/Y2ZFXsCqrNKvaTiQIw9NznkZuv2c1mA+5JhgvUuHREnft2rSgI/xH
NVca3w3QP9ygRmWXYt1GtkQHQocSwq7JJGjK8i1540WfyOoOawNDI5AGLoU8
Jw69i+UE0gWCLrLq2A3hUqvWrPe+zMCUIjmnw9lEiqMo/fpJqy+U0Ej3ebYO
VlZEMjM8irqy4xY42V2Holw5s8/hUT7aVmivZGGVFlsh+/+SjUwmx83BD5K6
5UDnYRGS4g9ZLPduFuN61R+rO0HLbUGJBwfnXSrCO/u6dvwWVp9uLTAIbUQp
BQBsVZ54OGup9sL5TL+vAUn3g7U64oDfRhtSeFxUu/g9uDJBGnjUZTxZqCXc
scfluqJE7GOQ1wdP3cSeRNGi9eF7jNiVGRhRQKjxLRcOpjvqozIxTVyM0uJp
I3vKN+2jmn+bM2qSlSz4h5wOz26yKvl9fRMmPYyzbRtbUJvx3AOu8GlubYLJ
xC5P7vbjzAYY3Y42Uv+yqNH2A2iYcPHjqWmAH6KV4p/8o097reBSlrdJxqJM
WX4ZaynvUvVMfM4it8+NCUJdR9tOzQvqdu7D9PAhbgXpiYjoxLxhunHHCnUO
Y2upot6vplKJdYl1jefhPIP/5FKrMZ6zXyCzx/xbcTqWIsLEM/efq8T7/7l6
SRuY/GsKqWV+cJYTVO+cy/VRHuuyESrbOwxuyaCYPh4wa4+mAvqq5j0XDxlG
KLQ6UGowvBfJ47PrrelvHu5HqB7S3Xuyz9FrPHHDLDG294I7VlPADBJZgpUv
qGu+XcwRoyNYNYkQfbEt/iJNOXSeV4cLmQHdUz5b+/GUpw4Hx2CgaXCmwmwd
lLV6aCWuXd0f+i9puYhiZ4jUUn3oPLGdCCpXh4IQjQVoEaY4qaZ32FNySqGR
NDEZRswam12OaBlTaHzB8VU7ZbXWvJCUNftHsw9vjOQDpDR4+VvuF/e2fyEe
SbBZqyg+WeSeFWBxvSyf3XOCQJZDvip9VAvU3+QBLpZxARKAZhzEB4vz5E+p
8YPf7PNpSCtMgedPenJukJdKwh7gS3EhEDuF7cprqASbKXsgcaZU3ts9NNDx
aEaWyoWDEiiRC/53z3fRBHhIyJESj2BcnDfyMR3QOc+y7AJhszWglFmPr7ze
N77lp50O3DYLKHOTWGEPTnjjSfzkbYG99/1S5lgGUGwoY/QJbaD50XfMbUO4
43qmMDztLsniPbMoFwphmfKQhpuIUV9FTjaRVftCjgeK9pyFeU+y9uQYafSL
/sFA3N9jFjvmlX7bvYaoPUSDrx4i1Oa/+tKdoOA+SL5EpoBKsp9nmNP7znNl
xX4m6/hiisO2dQbEIb3TlenO5mdpEYfQbdDxHW+XtteBEWQ9whLQ6DAtYaPH
rF8dmT59JDSJwlP+iz2mVWl45Icxv1a5qpekctrDLlavCpPZ/x9XceBKm5hu
Wu9ub7KQrEtsHUM2l/KF2df9LqiQXrgttmWOpUKTczytB3D2OBhd9F+EH2If
wy8DvhhgVJikrUaNzZmaRXrm5DVSv4gG3FSLQRDPV4oPyBDJ7F9lF4GF6rFi
BLPgFNh9QLDbA/3WRpAJK/3YwBnj2FoMF/n0SsILUaeh7UPvLwQ9fbR3IWFE
y1jExINfejktc0B8dxjOUwZFOj29QQeQRR3DbpAJqt167ZBdXAoZ80abghkT
f6ryHNDBBmE1kYU+Rhulq0lRtJnRyIJ56R5ESAonhsXE3a7Akgx4GKiRdSzi
MAisK+8bkj0K619Dbv1yOUR1NRLT7JtBM0fPIYoqNy4JPoBIYt1XHVOZzSv6
RtCxqM4LrB7L2c38n53vZtBlu6rNygjvkYjr9xB4XVnX89XNANUqmhxFykty
g7JZKJ5y/4GBpYaq4X1OlARuIU2dppGsa1vJPxiZte3G8rKfYQNOZYtnixVl
Ie0CsXZTIvHeFFMMGcsp4J7N/mZZrVkwU/qKI+KYqNGMZ1QETisOeAMFiMVN
90f+O/8k8IVIsSgVI0rsITpO2GnNfm2P8R9aaff+J8OKlYsQ5UWR7t5+hfEO
/r++8r7AIcQ0muVSDcShRBVI4cMZUlwmv42/Pn/Ijzia0P3SSZ8QqtUcBydb
ofsb4PwiVvuM+jlnGLUTaxw4iHbixqTR5/4thY2PxGGAew0R49AyGs0qEZih
s27nyGRpKPHPLReGcEI0toHaGEMuqqvwj2YSo5CqRmS2jVmzfz4pYOH70pf5
9PMBLY1remgZi8iHmzFEYQeoKj/sBtoFQKS0FmpISjjwkKiQzAbbw5l6VqEo
h/Wh1QJP0mIhPXhfQbPd1FeWHPnno5luqv2gjTHn47GY18LNTFgmoA1isEfp
L6+bXC10BWaStbGbq0KbY6Y9HchMf9G1YKZ1iWJDezoGh7PgR6aPK54OvOPj
SDOi3IbRdG940X7W9HnhEnzUWGy4y+yhuncCo6dDsjqJr3F5IQjI8Nw++wkP
NBcF8HZxXFwajLpqoI75hSUkry0ACSu2ZSfx20Cd3OH+yDagY5ZVPaJe1cxJ
5yZ+sth6myBHEJ8y3H3iVe6BdCBvzkJyPgO8DZZcpgUviM2r0UUPRHX6Gvkc
Ny3DYFwY31eS32VDCUD7CZuJGDKA697w5Dpep+9B4oQTXyHA2SV3xUkuZwW/
/sbG8cbfxwEcaHufyFRTs5REjG8EmNTzvi0WNPYthcYssgWDK32P0lT6QR6f
oXVrOJYIih8zr1yt6+UiVZo4iAbRQiqiNbcyMCD20qjJF8qrkN2R03lAlMkw
7V/2ctEwXFGFzt93Mh+G+r1HogIjv6nluCwQP2z95G1pMurqL03q6tEcbPAO
xUdoQWl2ne20Hy3213DOceXMfolldCtmqUWFeTtsSRvIyFp+kU26qDqpSuvN
svogR2e+Zy9mQt3x7aTVrV5Zp/mNS1sJ5aB9iGbdokPI9wBMJGEm58SA1QDr
kk5FdG2is0eULb8ZcawZ4Ov8NU70ou3ODkql1iKc8MptDy14UzKhMysauJ0D
V/hhFpreVRVUDTw+ILexDWwi42iOjkg+0y1eXc50jRRmaHgCIV6uSLNnSmXN
JjCEk/+0NzSw5hPmQNHOO9PkPo5e998HnvOrxcBeiItECtHWDESPCB2gYSRi
5A37xIX6Cwa+hGbZwqv0NLQzNpIey91P/AgceVSTdFvSoZv4iR9b6rEqCo+x
Vr66utSZC6dNSUwsS+FVCYlBTyWrwWHjw0WpwkMtr7DU79vtuRCMb3sXms+I
m3DtfrnyUHlutX/0W41vnOcCkHpYo8MDpAdCdJgCxNtMDesRLUQcqkoCWRLP
mu04htYpeOy4H84iSLbO0dILL93bTarVm/zjL9F2MOfKZlVf21z7gnOL/tVw
GlXCdmXcu6FGl8U+kUsLJWK5iuIVTcJE8y+VqtqOghKwaGJuPLDq4WmsgMOj
HdBYxo/ITdR3NNIaeApy2cXtbnE/OU+rZDJlJUOJDgn5jWlMenwig9Mroyc1
t26gD+Ajc7vtLVg+rhmM1UJvK1q4nXWIpB047kqZUcgu5dYGFixIAYfWeQgo
K2ozdM5BzekbFkGh21WDi4oqBoBBpIIuZirtTps/MPhyjR4Fh4KWIPCXL+A5
tip2QSKSHh/QMPKo39Klz8ySjnrLMaE95GAnct9b4lDFJ0SX39xOtXpU+10c
PblDRJzWqOKyeQp9ALBDoFle7NH2aveV2+1OpyjG0nCMcYZ2FjTgLTyAMHiz
Qdx1VGtP0Ep6EbPMjzUlwTKBQ3b2NQhxlstV1EN1q2YJBtDkbkSbV3jDjIGM
NWr5/OuD/3RvKWp3lhLT1RW1WLT4oZcgtiyf3RE3kKTJleh9w4GJymcx+ZwU
aZza2+M1ndLEnGgdpofy+0LvbSMBIkRum7Yg/DQvu0i+sefzDQFgokw9D/ru
zhzyx1gCcu8Pm5mqSAySJ8vc17huELekooW/5nTsjFGrYOTh9fAR2ehrW05X
JhbLday7MUEZgsSc3gsvPn71KTAI7Z8z1Nfy7YZYL2poJbWSphMUFqYkA9yE
2JjqUkqeuamxl3fk/TP7yJprg00m2c6dvPQIWu6DfMAELy5WLZblqV56pb85
4mjGVwJWspsCaXSXJll/9jP8e2wUkHt5Tfexejl7moVXFjneUR1ke3mwQ3yI
ptrZrAfVnJkLjx4bbW9vjCOHzMM4IsHyIAT7d475YSiHm5EOoqfuwbb5EObG
SlYiA9KEJxqC+qYD+4aU1Kz7Ep1qkwKv6uz5o8X1+36XoFyaVCD59DIIZVIZ
qwbf0PCuiq0VP3yMClcookp00DaHQlnZDdGks/+iWMvM0MGb+FWgAep9HHyh
SExQiP6mfRYKvyAdCe2K2PM+LepGlycLL9jCYPMzI/vQTn+ZWafTypOFXLyD
rfsOR4dOC7OZNRMy3COkF1eE929wuGRRBGX4dQtlzQ9/IpFblYrQbHZ/kWWa
YiENnTrFhtT3EfrkEEVrrrOWSEPowG/4GwuUOYmGyBD16dxNOhPaN03hNYpq
p/ywFmu6s6wikoktel3oECQbGoWW/OeRhuN+iUqy2v48jKm3aQFkXq9mpS81
YQrxzgH+c6Eu1keCXlDm0IRxuQgPf01SZ0nMC2Osw+4fLl67exr8elZQG1hi
IKmnTFGKDr1SgVLGC2Od4k3Yj0dOpfxujpKAs3lrBFGgDG7gWwS3W4K2Z60W
7fwEGdvql8RLQMzTx8mOAi4LDXSzwIAyEy7jB4sW+cDY5KHXhuN+yhm7cXyv
CdLJ/OgcMkgi2A0HExJ1Ij7uTwfAXZKefVZsyY02Alcq1M7Bw3N5URQQLLsu
uvHdrpEuKXrmMWodinxrABfF//VTfHFMxHiSLGY280kOr3nEdu/DOUijsw5x
QafgQN7FKnEeB83U4VIqFLeXo6wQTyRGRY9HBSC1MV05oq5ScNDgShOTgw9i
IxPGs6v/dBzo2UkfkJuq1g2mC++fVAmGeltB6mwXES/xT7AzFWqa8SGWAxGE
lsEAeVMMXAmjBl3oQ4qLMW+m3i4/U9EScVo5eCRD26HuP1Yg7D3wPaCRca2J
ddZuZPBAQU0NYD73F+rmjzVgQelJ3pnm5IvJGgCVEyw9x0hhLKpKRBfZw5tz
+Q6SJb0U1Y7QfCLkvBrHx3hrcO7G2/edHn6Nmi1zCfPEk20wBT5NYFl55HX6
lhsMIYTFxX+QKW4ErUKhJ5ysjB50PXriOKZ3/V3jGPiZFlDXfCu/IPRjgTkS
+/XdIoWDEYtEOb9XvmmrtEOF3aPpUKl9zx9hN3dPYOCOthu/kBWbmuQVEpbr
GD12HXRKRxALqCEDplOvFz6yi/4bjwpZpqDtmdSOLABN9CiLjDbD5ZcyHcXI
T0bxU3xs8y3p21HwHjcechdT1Vm79l7E4GgLQhHc8bu3Hi7POW0PdcwOgRsL
7+TgxILkjF2x3uqMVqxN/rhek0g5iwypdj+tGmJHyZU2fDtY9fovAHd0eRIa
pf329jSGjpySAHlfjbP0sHeSUl2JP5CWSmo54I9DWfiel/w2I6z2Xdc1IQjV
Xcu/Ui+IYkSFaRrwaxzonBL0c9Qk247j4tiQT4fbLzcJmyRjsL/NQNIPLq6z
hYkNiJWPhR1trGjYMx0QCw3/Eps83Zpto+frXpDg9xySArAjhnd8XCveDwpT
Vg2HTIz79UDbR+Bn7GQqwN1a8qe1mMZ++UHPr9IgxKl1ROZTjaWZdNiiU/td
lp7/ZGBUTx3Q1NEpSMkpstj0n0LvveGwM6E2jCfWAvC8vH9XkAAy3K0ZcM1A
S6JZ5vgorl3Kf5EA65N/zQzjbnyQBmWRf7r6JJ6sHhDMtzTNT5NL2fRFQ3w9
lIg6t8t3i8bOCpBohD/NK54sKyVhmu2gsht7dUyjeTmT1mEGkHfNdl5wb+mR
tMQ4vZg1+649qsC0wkka6kw0PAlofd+dBMT9KgtsUzAw/6hSLk0wAVSbDL1t
1oW4QSzBENuXXSyueLTSa3xSoh4Sdd4nzR+TpOBQqvKlKrQ+p7B1faapqr7O
jE/RGMzaDmRROiUmnejlN28RfybYdIaNCVqYKEIooa0xYKPifZm0PPvRFriC
+hlB2rC48fLrEMlg690qbyTr2s5pDFOvxq6t0uoqlt4mbOSeo+dtlEjGc7Qk
gVtvaetwhfzUA9Y4gKOzMPVDh4NukyI1gvPa5T5iy7aOxZ8k/I2nlZW63IRj
zgVce4BttZz+wizhdz5LVUdmEOYD/QVuO8zaG5HQc0Lf1j8SCr4T7a/+JpOJ
8ff/ujtd8w+Xo32aJdZWBxzPeBtgnAJMdwLqGImHAKVaFJyJwVPZrO5tNthg
1QJLyd+O8bGDfytn8rerxk1JPLbmPGXTictEmTSyxeKWe6/0zMKD+oxVVWn2
DThoWK5QAjsUWnABF7WxFeLKgSHhcMlCE48yDfQjSSC9w8YqOSSNg7puQGty
3BIyjmQI0lpTznz6GI0c6U0gUnlcdkPlcKiAd3nEjOBbLNXMRL3ygRXilDZl
g8foWxnYfzpQwy9c0Dk8xAeUpv/vEHwEC61GX8LSOHOjaHXDYWdqVcXy3TYA
TADQj9azGeVCGf4AKRodJxrBXNYZpyPSerVKxVS+nbaG6SSF7U98V5fzfpio
NKWPEZgrHSXcMTCnMfkPZqF0WN9IkjGsah+rjg/Ec159kp3DIg4cyLPARdCx
wSZbVfJnhirpcHE+CFoL1na0J0QT5phiGIj3oV+zJoQSuQuNXi62S+fXGGyb
80Cbgcj8E7PumRRaiCUhtad7ma7uPDgsKw0pBV9xto+3OSkToE6/sZtUbe+F
coETHZvZCrgrz0v3tlUcw7TTaOmDVXoO8pAR7pV32NU5m/CQi/Hf0ObMxqGi
sRh+CdJ/ryCd4Nh2Y/VPmNU3pOhmDgMa3xr2CCm86+2RZjPVtdzFGtJowTOG
SPdi9OdBBxPDSxnsIr8kN4U0oy/MXbdjyWzngOshvnrWQICrIi1UpIsB+4Fe
s/EnlFlDUq3T8IpsxuMHcOSU776Y7Yk8Se8QxPmjmCbYsdrBvpkslgsj3R+M
6vdxuIvm/wTO2X3DQY6PZErM8j2EHVSibky1X9dYb4hsT/72dQDJXiyWFGGs
7Ia2X6MXC4jyGAsacHpQy+H8mBN7eRememYjxO9my3Wlf3t391ZKEyHlZsZg
ooddUZ9KglDc4Hq1AuwFZWi6YvuKDrUyhzkSIxTNz/MIXvNY//xLE+H09lRv
GmUumnAgBduOvvJ071UCWpOvP0BCZTDurth1Sd/Z8JEcJYBSarQidwitVI8f
MrLNeouTexvs+qmSu4Nc8LKHmMZIRT/5NCVg4Qe9+0Y/VNUyfYr+Y4T9KU1w
OvTWn/plFNzv+XLt1ttAFOqPutTs0hgiq4ZVqul1XVKHOskHKXxWvSHl9ui0
QbXYezhie5wALVZqzq7h570JYUNBsKCY5ZIOxQ+mLzctpAfAUycqjAjZ8FEx
j5J46JcZdQgiUAN7+C3dcvhJ/rqaWHFCIzdN6755g/rLFwK2XqFSWnnvHZdN
JRRifE0aPHyY4DZmKzunoFtWtupm1oxO0IOiUpd/TcTt/FIW5l9HJdS+o/N+
pDrlzwnREMwQ1xFTYVLEsxGuL80ETkgwBDFdlmFe5H0xhxCNRvmANC7saj8S
GxC5QIfOB52ejlm1/ViPKlyxwfnf1ZoN3hT5lZIV6S+XOb70A9JMHmVvswVA
gG3g+69lelbI9KBu4nlUybmovVML5n4ZqW76izvXl3pMLYxGUgm+1zok0ekB
ssNVdNxnUBfApH7nZ/HbTaquKlmIPITthB8mu8KZY1usCte07Lewg104nawa
+jgGfokDMVaI0AU/R9CK1WHP+BQirbOE1lgVGIkkEC6Kz3MlFTafNhogzJgP
rITJ8efaR4WHgJ3SXxmtwZ6+Mon4OjieD5A0pnSbao0CVH3tUxwAcnefFHUN
9P+wowiAaNtwMQlZYdieauPA/CSekSr6lkABXwL/PpJhoAXjTucyA3Xt6X95
Rr7jysXIg9i5/WFjMUSJ8+RCwViqDMPlxjJWq/RXxWQHVaOAoiHmNNiJTLHX
P64GCJ5dFbOVDVcNSjrxLHRaOAZMEoGimZ2aUMQfIdQsZsS3dUQay3kZ7sKq
dCNA+ModRzfdGpBhtepcjtnef/aXaXrLEzM8JKOy7gmbh77I9ES62znDcu7v
WxL9cOwn7ER8CkvqAofqwn7nX3DkObotstK6iconqL0m7yK2JWXl5/KHoVXm
ZYbPBfm6k7YbasysrtClXMpiSQ+/1wWnjoyKRmvraj5FMPdjTvNok9FsmriT
39rc0JVs3pA9SAgjYkrpBykul3RyaNlsdnZmCsVTuFiPRdL1yVCoM9ySCXaw
YTWild06y68IcFN+1NrIqV9Q71OitQD8h+wV138DgVh8/n1EntVI4Ux5o1GS
U4m6rQZZBALdYPpRjpJs06GPUq1urtFi/vYcZY8Qhr63N0I+gaFpaLaB3D++
YLM//7D1UCpO02N8RtoLmqVL6XrZT20XN/Ozk769lfzdM8WULPnQlqdRwwzi
J76PshbBfZZmZoOPmeONKF3AdYLTmsRy47/nxv9yYej8TqCMgkbstAM4dclu
sfWOGoB4nex1+/9/aZfEA0EWbL8YK7n4pKnuRpt45GOL824pYdV4Eq8WIVzM
deSri1q9QuSExt/l+1Ow+0Dk8XZVZzr4tIs4WvdZktfNkYvjWPH2gskhvHeA
sctensahiYp0Q/oKBzTveCU/N8S5XEY4xkTWwHRM25oAHOCZDPBuLLzVvI5X
b2wybx6ylmAAhfPgBGzzH8B100ig3F9fzzmm2Cwl9q8FM5RyQtoOYxqAnS8v
Lkonm3axuMlLh4BeL3gSVc7lAHiQDiVMUfnJYdvsKGNu1jOyT3748Qnp1Kvb
eXLmarwEboTTBePQ2gxYMTrHfh88MSpTedk5jQLlQrjSizcsa6gRP+ZbbVHi
qJIe7EdntJitCgnZoLw16otJzGuF7oONjunlyFCfduhN/GlCqyU+1sSxw2GO
IqkqmkUyOncN9tBo8cdsmTQ/SUUJ06HrvmPR+TJp4HRdCHLcZ+tcVzW3IKcr
ofWkvPLKjbhg3aCYoJqDAldJelu2CzPWPoJi4/JMqsOlB6uJmMU8shINEU1K
n8wskzT6sKBkIisVGK2vXm20RYwQqMkqel9Z3xWbWe9lhAwCzglT1VfQ65IH
lkDv5np68GNa9HO2H4EP3uj0dR+hEmt78xN6Awy8QjHPiVk3AWibDIAczYzm
y8JQMrz8qtgfHaiQTbvdDNGUJe7plUt0kf9N2E/QIUETajjsOI0Zj55JBl5a
zf7IYDLrc8Pl3fsc/Eg/tfQ8u/lTCtCIna87YNTMciymu6e7x/ORZtAKfTGi
3rPNiO0lR7oKHAgExPiAprue+qwsSDtNL87Y/A2YioaVm+TE8vPXJ5maoYI2
FiUuiVgHBGnahEo+fO0g30eKsNDQuNg/jqik2TmQPoWBHurB6mx/p/y2tsSn
JhRVWYZucIXW6YWaQJkuWYmyxSWB9mlWdFelNHG1OzVWp9CMmSfCWgPsC+q/
5gAGbWceWVUjH0yWyTDm2dTfVP7nTFqYxiAnOXddNyjStoruxVFK5u4kqWQG
CFKGXrIcDoz+yfcVL2zt4aFlLHbNQcO1+TEy3h+vkdwxELb+SRBCZuPm2Zo+
fY/a/15OHZvcF8iK9FnASjR4nKaHP0IEgBH8cJvdjcXK7fW9umb7TJhFe6wg
0LS6KFhXpOfz4qOwBpVJRZu3noDe8m2bq0qj/6IfUskdS3CkkVEJjDGiJ3FA
mmbg9ydPUDy5YAqTnOeVTQM1uu8DKQiz9Vv16/2ddGnmVfYuOAGetXsYotKW
VJaqvsVYZzo3hLAICfzdvDmB998/0hSy0t8r31EqdxddYjNsPh+WCMT1oVS5
AzthKd/jUp19/+4AAlvudPEFYfvNFMrEllChZogEtKHxBdyLE1zSNjPN01sv
WCnud8CyKj/ovf4vFrUGdBQJr9lbNQ6X4/+MIvFPDPeyOvzYXsu56ipc03uT
P3u1DQMCtNIEcM2ZUf8HMgj/f4oiZQ8sBQ3jpBvbVoiySk2gZooZrFOYfDcA
YO3yDuidbYEInk/yOenRnVKoITdBwsOATXNaqjLQ60hAZwK2CoxGEg3LBIuh
etZNwtaO/Ze4YXBKXg1yNrPimFXOfg01RyWHnYWWEAivT4iO+C5UfIIsbL4z
wIQxkC/0t2iwOsuzOM80G58DMVLVa3FsYdo4q2fVX47i/8hNsQVRSmaX02JB
dKaNNL6+ge8/z6C+xP3Xb2ZjSbbcJJr392EEvW3c/TG2TFGGK0XkcL6lQfVM
z+/t7NE+2DGC2Qh9F7P/vXzI6jLqO0D3QIDdAbq6ioGF9idMbxvynUr1evxt
jsx1Y6OR0MBDfDKxBzZlWnGMgYydqer9mXWpn/3D38Mj1Fiax5REp8+MMdFU
fho7gNo//WQAzA3L9qIoixrHt5BTedfrHEqkDi3VpaOJLfAr+tEsJX5HocNv
n6P5l+Ikv4IsmC7iOobCRT5dI9NXV32MhP4/dP/srxcU61sQ6kMgm/X7e6Bq
M2anjIGwfESeePTodifTS6Xox5L+vQLKZcA4ru+KEVoPh/YQ7qBVhEgZrrPE
DBahoPDEeVDd5uibBN11xVbQljDaxcPid9FJexWjawHguDN4dNw1oTUmAg9Q
CEbqSVHmEZUve+jo6umDxKMvct0CoyNEKu1RC7NBVM+j3Ez3LSNWReSN7N7v
ywTMd5zyQ3RMmw2kV6wZDMfpV2da8DFmTHxpT4ULs7fHAj1nvBT+fdt0mRB+
WHtMg/PvmmJj5WeOS51I2xIPwucLSdAsEQF8tvmA8/gzk/fD7kjnzRg4+zgu
1J9xT4ThiDBk8rpfkD8HfZfgGYcFw6RimmQmmZfTXiw/mekpIYkb+o2vMvku
30YuFBjVNodehKITtmynx6e6pw0OuNOil1yo6MjNdZdGCDqEG1DDUWunz7d+
R2egiCT3cy2hV7rTbWeLUi5osnhvhJ7/L+T6joXysDR3IBAee8+Nb590IRcZ
Opn2VDrMlr85d48H2F89/1bhAhtqDwAYjQSX0zh5n4pKF7TV6sxRO93xBkWS
7vY6GfXb5gzOMRENz/kXD8Ol1riyox0P3Ca/OSVzQznz4SCo/D7ZoMXHW5SB
D+NbBzw8cSqEvR+tjINiNj0UUUj9gTURKWRhlR9lk55xKy7PceNKncNoLfqt
jRwBqMwSRlWN+9r1bYTVZw1v3NkOlFvsXZnwTlBjOgURKhTSy2tGSUmx3boL
CnoR5MS5u5XhmbiFLkt3Oni2kiTTmDbDBiKlZhWlcBhFJPRCdi8HzVFd6o6R
PA6HkPEnxnR0tEwy5n/U009anjtSc8XmNoq2uuN9BtFDE/lRq0r/mMHuIWr6
vxvyk/App62Ghorvu5vRjqnS5m8+bPFb3SUe+Z9iRK82RGSazH4eWjrksuHp
OZidde0O/ADX5IqdbvZUXyV+r3k2+Dnyv+cH38qkZVMPiUCoj2I7aBaA+lmX
4HEhJ11+PKXEbxd19alxUmJ8VU/mEO6Cj50pLOORT4xM4IqKQDhzlx4lIrx+
Uel8SAIUqKnjLvxGnT9JyyoX44nURr763LoGHGGvMYnJjE04x2r/5aAnyPfn
d31aMrKwJ9Ic7LhFaSFw0E9/COPXir2w+AZ0yddXmtOSVsBOCmQDThKEHEeu
WUnzQ24CIe5255wIE1ObtGYwZJ9j3C2BS4n9yvs3h3QjIb3dv2wckeVGAmBW
Lw4srcgLcoaQLAOzhxsMVB5XEeW3eS6qFQ5rzJw7g6WxTCArHYLvYlQR4Zx5
uDxQYTKc6an7QE6ejzdz+x1AOI+ygm+Y2Ch7HUqe0l7r3POlNyNb9CvFQRzd
hRymb7lig0rg3mLcMa8XcHgLbWx+/SLO6khmdgmL2n+FGklgP7ukZENzCdLb
ML+C5+LThZgxACd3woEEPhje8zHWYGnu/ihDbbvVI444wuWbU3hheWheuNic
k+cqLvDq6Mb1iPkqOfDw7SJXD8mZYK9EBkc+xvPjb7g3mIS8LEyEGskmRQt5
bBcy5aU6n4aKLAOYqR0U0bFd+dVekppwOrqHWX1b+b6ZWAUWaIxWqClLu9c9
ZJ2/Y2h++bUdb0Yu/OOv8ulUnu8eFmTiVLxQB6hzSNc/WsJN+wRbrxTgJ+t3
jnezCN1CcWPKUaNOwdnu6xQEPDSp6J9Lf19Q6XF95sYAZZWHKEFSgA8MVReq
Bk3L9dRDar64ja/JbaTn4YQjobsLavF+HoHlHDJwp4vpAUujC3/kwv4Szp7Z
JMCXNY/ImKi1j5Nd66Wr1UqqcQhcl4QEH+0fAoXAGSdufam+wuBV0CJpSaMV
8vAF3KS/WwHtdVEYnfiKlP2AR+IGL/TTNABqKKD60mDmw8Q57UXnbxw/DSgk
X/n/+sQzXpVsiYbsD0Ns7SuPW4DK3v844yVMJF91TQPaVSh0l3c056AXwPHS
eilK2ozyLj2gIz9WEbfKto4f6FGcGxZ7bpjl6pHkbwxN0MwY1jarjaSRu6+f
c7oef41EdAyn7Uo4J1KJaQVn8FgPMVOCMklt0px1n0DBvysL6fmPdjLuWWk/
6tn12eEpbyFcFmb6qbvNBcTIR/SmwR9dyOghsHs89l0Ot5e2K1n+e5EJIucp
837mFS9L1DhDDhsKo4ViYKNmpjFGaEQdTd2Fv6m7vVUpMF/v0UZ6uYqqQraU
NbsGibUU7IxgESW3tu9sYCp6NQ2zI22o0Ib3ggo2uXKib90z68Tkhd6ax5xT
qkE3sKN41pK9u0ioChTG/kIGj74cavhMr35nvnVU/mz55WibrPsEuGocH6F9
YNlzhykZ15ItQB5slA1JqZNFApvc7iYe+DHUFjKzUEa78L4kxnxYAAYXNGdl
I6FMvNrW0yuHZk1SR/Rtcv3gtsqLNciGf5S1D7+8BdhJYPdS3pBTgW8rVYWJ
yX0gxB13WVlx/QLvRPL8hJUfXnOW7qo/48fTspLi7H4NVAYgxa6niFDRw/bj
nTpNo8fTZ6Y1wxmEE4kf823+GWnzqJhBDF7DFk7HJfFf5GpUTPnfDZRY+nxg
xn73sxuvIXbNWNiaax68PY3jN8fdYAYcL1kesGAV0BannzzoHxHQdvaCxLH+
K5x7wH4/pMfA27dPkm25dggO/dSjBMUyVNfDmgHgGC1nZkdS/p5aGojaI5zK
/eSY1Po0RfOI4qM2rCkbSSAZuefJegO8OG7MN9loBeo6YdTF2QY7gYPfjUJy
rGlhVCR2OVqFfpjm9WvRQKMH6X64ubalZCjLpbubW9vA5wjj4WT2s0j5lRZI
+FVRDw/Ur8pK0zdydZbnSjV/Yap0R7r/OjZGLxYX8LMjcCznXEGsD3Flzb+L
Zx2XsxzXMrKGcZeC2SLOYzYNTd+j1EV9ZAmwEr4+hmlLWDNjw8ePfeQDd3Sp
fzOxqZbs/VabbJ3nJllFuv9VMYo/bLm0b5rpRZap/Md8VcZ1LJG2LP7yuRWv
kCQT/k5yzjLh1JFkJWPVtpL54Ou5WgI/fqJdq9dyXgET/YK/V4dm1RiRENms
94UrNrFL7v70VJ3zWZg4GCjOj3z8Ssqe4JvjOS2RBnTF9kUfZr/R/f+/3Dpx
2o9zaDU5JganHOz4KG9vsIuSXi3UQMViSJ5wBOC7wbTLMqvUWQeworXhtS1e
Ty10ST99gDwFJGF86Id/BGiPnqTldLfFYQkvypzQjFEm/HaokC+JfqYlLjFj
PoCmDXrNyPoiBi46gHQ5eNqwpxp5ofsAG18mpq+h4BVwxc9vzOgP8lQ8j9bO
V4d2VIn8mJPOkXApGXgzDjOUFH/s+FNLFAk5ZwKiIuu081aTvehK1m/ZhJ7W
ahbW+8YGpTynKCBXchckTNGp6N2Hc47t8jeJceJNZbzYDe2JbY68By8TA7+Q
Pz/X446tJMzCsSJTwqsXVuZgV9vA4dd4d4WCXZ2YSY2boiJ3dkD5oywPrduS
0brFmlSe+EeFUKv/db2NmHbzEWHvMKfNNj+2NUrrf6De7W82yhOmP5wIF8b5
UPoTecYOjV6WuHqg/A5Iy9RrulplvuVqFMLPw7SC8Ci7s7m9xANPPKwde3n9
wFYHiz9wNe87q27LRjrb7/IxB+0shNJtVGFfL1qX54lK+NeYDfv5kObIbOQd
E6epvnEXDgYOPFMsKZSNQReAfGtdreQ7tusjQXmVoRAuS30+VC9KIwyYB1/l
Nzj63xg7lAmv2DzvP/P7A+cpPwMfJ+ZiMq3kPzcYPKS9aakoKqz3dDrzxu3n
h6ATteeJfVkzo4Jh3RZLtZ+zgE2XcxgV6LntRz7m9/9hpa1Br/h7JcXKRiXW
cIHfun/LKmIoUkV0kCVVKRpoqcsBtt58MH+wKnaQEdNLxSHK+fcZS7ACYPpK
t2klTTrD04/3goCNIopNhnWgIvY9U89Fcq6D4njUpEKIN+ZvR5jVbRaa0fCS
Ldv/U3ewNHui2ELwhB8tUK1pI+F/5lDzFX5SZLenaJ+umu6DxEXqVHkmIypN
Flh1xWuamNN8pXEOyC4tIgkAY9YnEbjG5u6RChU3fi4IuT3pvahdXFr4TA5v
JeKtEqj3Jx8YJ92+wtMYk9+dDN3nbCJGSArzqVSep0coUklmW7kGY1VPn8Qp
MrZDJaMpT/GdUBwAxTlqwNTxLNjT+izZ57q1RJEvNOeLOHs/zQroPw3P93NO
H6OchX0+X6jsjGjaq7WHw+59OX3TfoVTsNxJhsQoyG5I+M16G/YStnmTUvbL
FMBj0asFaroLpw8kXT/dmiyakhKnOSCxjV5XahpgSmSIivh6Su9O/I9+nCj2
ifXj0VbUB9/KPb33ixPJT1uUH/0NtGhufViftN0+H3Hs57hVKzOjxTcHKHXi
vfmoUA9ZCa0halRHFw9FSNAcJ1fnTReCV/WAhecnPQTLNVHRXtuPoMUJt26m
otciTdN8oiYWNcau/gHq9FfVb01sAg3KTDRq6Iv/jJl1I3TSjQhiZ+ahGGSj
uUaJr3n2ZuEdMw46vtCaJpEJzUEGroUkJ9pcynhAB1W94LcIZtJTqIQe4JHu
lg3hSbgEAaFkLff7OS/1YaDwCkyudiOwijZFXkVdMmIuPz4aHxiLgmlGfJjN
6FFuqiHjk/oE8DrsUsNzzKJcuVHXKqfVAEmnkZHOR+P7FJ1nn0H9Cs9Q6Pbi
qeiimg2X/LIafS9ydw1ILyiaECVkzoCxKEy7dl/kPBoqhIc965I0b4PVxv+b
94Jp2FTmvPplK2x3HfXGNJNozV30aBSufESTmOteybUwABvltuei1KUwgMpi
amgD4Rb2sT8nwX/eMgU0tIevB3g87Gno2qwKVgSeIwf4gdOLqZjpBPQ2f/mJ
XE1gCyWB/1X0zdiQ3FlkfHi8g9aaBkEotlIgj8QBR2qb2VA0MKEeeSyFalQa
uw6SLpWk0168nWoNoINl0NkeIup20kKAfdq1dXJJuzUhXsGu0NvnO1D3shLw
28+ul9A8AQP3EnbMcdbBkgADehc1nOJn9vGrNWyf90XHUcp0Mrf5shY6Qv5i
Wa3DKrN6zDbYcUwRyrbbcgjO/R8BbxQjg4XnGaUCadLQrywsHfwMZG6ALPHA
XN7NeLqHWHR5XEL4HpCPPUpbR5c6RGrI5C5Wchxtiu6GTUIBE6HnqOeh6fv2
o3cmDf8hyTc5jQeABkRps1JHxq6ELc2A981ErOTZiCREubDl75DFEP4EncWG
PfVKL7QUN+sF8F5hv1OeXg1YzW9MgZMbLRHYsN+55F5rULOrAxRGyC/LgliY
V1H/2CfgAtHEW0DCD+/JBG2rKjHOw+4tjHVIes7hXHvDCBbEXbucabmEnuVD
TPW6XbfPnyczWYTan6pxj2DoA6qq4F+DsPhXrnR0RSsHYpR0bG0UDAGcGz/b
Mpg/0KW0KyPEakYHTODIeUOCPlCstJrbR8Ke7+CdYaUOLh2Ul17YYyI5A7Ta
uUzuTep5G6MqbSIpbLFXKV7AjLdgdY9tVhdb15I1x4t4vjHbMVATt34ClO2o
gsMchBX3q+7PO2u5nu+gKzCSr4auDlF8lWk9XpnR3KJD5WJXL8Tj/d+e4hvZ
SuHyzqjf9CZKtdZBFJG+FLhALFw+hYB3hL8VVTG4YxH48H8UC3+s/DRefW50
4LRfFHmUEmVHWeuhQ7lnQ+EkwVXfWurG4eMRky/Vw6SGlzBdp75J3qt1xOJz
XKvlq/k2m4ixusO+IKR8KKfnbCyCJuMnjbSlTjBUTh4UqtQu5i6QrIGqVYH/
21MQhS9cEEViGrLHb7n/L9IjhhHRyj/kPfKOiXxv2YioZVH1Ip//iOO9ZgTD
J23TrwRrDRZbGQhHcPPY9aW3V+Bc49WFMUPmh4r9ylam/Wc/03XyFbhfjp43
gVAF4HL4l0J26ZFLiMwwDh+Y5IbKFZaQG0KIKypC5ypEsRTGBZ5b+kHb2Pjv
A5wGnp/boa6on3oMEZcpi8MxaVanQv+kjMEDV5rGqBxs1TQvav8yZ8rK40sv
NVIVU9Zvr8eQSpG7y/uX2lwGaxykTryZg55NbuT6RxwuCvZp2ayIy3uR/of6
03JrCtxRH0Z9q4X6DJy90HlLykJjPonWLtCUJhMGCRfnS3ZPQceMDkVXwOn4
QWoyWJCwZgT9ruJL4h+QOaOlWRf4vdGYdEe+7HSVou6uNYn9LdNQZBIfJjyj
OIhnP6jA9L3sVmLnEB6mHS8P2OV4EvVyXIyQblIxnubPwcYi5JGpOGJ4XK9+
x1iiGYss2t6+pHp8NYoLAjuXtlfNt0CkxWqS7i7w4mCntp15kgGI/JBHsZoS
jfCwEuYv5/4QnKcgCSW+c8Fco73UZQmFKqKLQfuLe4L5Hw10a44rlKloc6yw
Y3ifYw7qisXFGlBuV0Eo7rHFtM5OC8M7hhqSZte68V6kBAe/rPtAmuSqelvO
4j2abwAcRtt8N4BT3kQna3iQQbS1mojz963QQgl4BrHb/4jDd2WhjooZvw34
A2nMJ3QwFzqIYJG3lo96jv1XFrQmTS5VtgKXlLoCX3wp447Ej2yr5x4uuEXR
h8mBnuIRBn9RnJ1XuFgQeaZ/nkqHvNv5Bbe8+gNCB185R4zPgiivON6+iK+2
Q51Q7nF/an0xpgPgQSl6grIoMfsxpFNNf+YkhZjIZumkBZFz+oc/oUXOUHpD
NhEAgcHAuhheqe4DYb62BawpwFG30rL+NL2guVFyD0TjH2RYv2/EGiZcl1+f
zql8n0UPtbjkmaYXe5lzrJCHthSuCzHuoXG8obrHc/sZGAbFUCbjOlrTfDcn
qVt/+iVg1aCO+tq/UcXoIrh2vmkhYZy52ZnmKyfVgbovdj7cG6SEMyRHLciC
P+pCDKmZ3f4+YCC5nF9kGCjSq/jkdHx0DzRN/ZaRzFLU1PtVKI9W5OsArYlT
8+UNVPWo3f/KiWs22LS5O0mHXwRydh/dvXNLsEeykBPX0rRIAasEzT4TmAnD
2v7S8nsoAHGIt9MfefOLIKRx09eFiBTJQ3W7iM2Kxzeqcf8FiQ55ATJxBN81
qogelKoynMdJVscTQuQcLMe5Qmsj4ZkllkKXNyuPxM+JyBYwYIV38Jd6PQik
RzJe/oOIiFs4H/rWPfA/L9MV9eiYhGEIuUoPuQHG0SwnJWt9Gc4RJn0WfNa+
goAQo4L5fsmHOtoBX7JU2PMRrfBe6SXrpFEiZohUMAfyB5fzysJN8UsScZvF
/QNvIEBosS/pRpnJuy5n4BZBYAowvb7X2yZVj+2VFd1dCTTFx11lm8cC90oC
i01dBg4r+lsLp4jD+xw0iCGr8SEotDEojt1SUN/VFCtRa/sylgGhIfAbIGTG
5z+G+meiH5a5rNfDfLPoPNU106nRsDM8ckQvN84YS7+YzhwpdxaVnC+kWH0m
HSx13LNfMNFwJV2SbQbTMNWEI6PBQXZov9ki9wQzHH0OmCtjVGnLz65Y0ZeK
2q2+HVFZ+pVaHBqw6R2/prSpLIO7NwwLM/iCOxRQF+hkeGu+Zx48T0xpxyTu
1ML04FBFd2kk0uEJqDsYhdscL3Ov8g+3KyieghHUJIFw0W4fUnPbWfPW8AKM
WsNcmPjwnXYiHXSYCzNS5TLElLeeqw2bvjWSX7cI/kAHdGPpEldOe0usG0T/
iqcQF8yjYYW6P/x3/y2g8y1UDNUmg2r/81Qa4dc4U+T6Ox+J5ze5r43sHLX1
3EjbyG0QRue9pT8vQQaF4CgZCHvTdd+v2pGyHF5YYHcgzKklUpUgA+knVpSo
zp3uIlRYNZX2eRR9Apr/VdW3cH8OTEjIQLnRdl1fiWZBqQQ5k/dGTePZzHfG
yXhMlRSRy6vNNl6PPwkOoS5D6oUY4gZBMEzu+XYxespWQiSzgS18vx5dXTFM
BkaGWvFaeQiTJFBfubUJks4O8aTJnC2voy2tWcYbTvulBTjPHuhwKSYdT7bV
f9LaGisRY4A7DnHYzYguozh3h81RS0qX8UNcjetMQNkBt1xnGNwBKhVjiL7P
2da7FJ1joIVDV89ysGr6sFP0sLL0iXSU0KPgV09A+BnpONiLg84j/ikHff2l
02mZTMRibICkpQoxGiGnVKI5lFVBbfko+J8kc/VQwS+vSNGf7zwJRKIH/FvX
bF2NDGrWsOtembegpQf1I0kb+Su6tucX2Xskl83DYcO13QNCjHx1lsLGw3og
Uk7ZC4VqAqtNgIL7V+IFT4VcN06Phxhrvq96fWQZ49U3qQnGjLOYfdB6ghpY
yOar/MyvuVPOpzSz45Bb0Woewy+ZbApjpRxLNSsi55TTPoN/qSZuNU/Z4PLR
EM658nveGVwYEiMc3DdPCzE5Wnph6pdr5jJ8XXa32f9DEgARqcSqKykN482i
zDH6t7pIaLZJeDvjkvKS/fiyxAvAjEqhFRdAN0N5CCcjhvJR07wAsOctRnK0
wZLdN4fV2Rac0JulhGvCr94e0K7UDkQJqmkhWUx/23o890ffxTEDnLhDZHEx
6lWLk7sQJHvD8emoD/ugUI4YK80yPoYRfGC6MxUn3gT+jXsT+d4k1YbqvrvZ
GQbUgOptYgOXUSfX/3z1n/PQQi64K8wFJrrTHgtaHK1Ckx+8fd71ItAMYDOq
k8+uwjGTuogt2vAeBoD7HNY9WBU+DOA1Eo5G8OIB2QvwLl35RN+V5pGj/gv8
LysDTCjLMwOr/glcv+WA28bfqcSaoBh9ghCEENYgQdd98zAWPOjT3tlNu7Yi
D3TXjJMoouJq03PCZtzCJOjS3mXnF2A+wqUn5TFhrMFe11d2fkrdNYEj++Ot
lyy3vMOkTvUZJLmlqLxr5Vi3Dbpit35fx7mcePzIUcv0Qj49r8ezzjgK1Zeh
WEzLSyRYmonA/ZriDBvgeG02tt/lT6g6MdGqk6x4dRIlRhE1zrrKInAH+ogN
Uvgd0y1RZDttZB+mInokarmYQIoEnTUx4Th2kexwN/+SQa1GSagOE/682vEV
FJR6WNw0i70+ntDIA2YxLUSEUoYvwO6ZcY6GYV53VgrfyR0ZcJOoLa75cZfb
H/v+EfabC6rATJjGsp+UMQpnbXg6H5GwYS/+SjyG4eFrpUwmV1+EEW7bn1W5
CGzeGMu52eC2/y5Y1VHl79JnXqBELvaENIhFS0xF+b9hL8sqD5DKI+ofH0Tq
QTqMINFKmcR15LP/a97qfuDY2CigY75KsoPuEXrf9X8nkcxLlD188kBNowYK
7TyNaiQbWCQRxBAbW/nsr1sKDuC2YkADrGo6AIYGTsUDt9KPenAhBIwM6eKq
M+BbYOEBVEF4YU08B89io/npMTrpL6iRGUuHzTb2PK2EaK/+q8joxWETwXLA
JMx2BU6X0mn3wCMTQBKaVu0Cqe8mEB8PwHVxusCnoZ9BifVP/cywbKaK8wp+
Z5uuwMM/IDZ92fPOrV/BCBGLc5UTxwKNZO30Yg6Y8FkdwO4PLuQNU4qyb2el
+nuLtjG2ut1uYBZDt8jLIUu4FBFMb2ZUz3g19MlKoWCEkBmTLxhoad7uMwB+
JmVhqVhFJ5T15yDUaa6mEsfD0O4mUi803kg6j0L64PMYb+J/4TZE8OVP9ise
9m7ejc/aekfNt1KhY5Hu4TLPxjIC3L7JsNTuTUjTZ5Xfw/ltCH3kRyIaWChh
msOqelJ8Zju5l+eqkbKg+hToFDVqgEYbByMj/UQfmmJXQ31rygk3l0zcfGj/
WQrdee37kL4GnXI4ZEmQEI/9bflogvB2fsKcKNFvUpB8TlBsOgJH5HneouAq
V6Ocq0ksBYV0fkifl9VWiOM21ynLAweiHi6psc8Pft5mQikCHIZauvYUapps
eB3onvLgCXKCLsN4vliQHP39srbod+mCNx/lmFayk0AKyTJiGtvLfoiwCKyX
WhEnDEghB925yRaRZFDPbTq0Mx+PFwUCuCsNW2fX4G4JzFi9I4BwG5WfT7j1
6xCtVuSpI+9oZH6Z7T5SQuYTS7ULfsLlLP48u5Jt30JQS3j1MLm3kWT+g3gi
CPD+dWOEZR2aAKpByGTftaqWELBCu6D9YDZW1GVsNAV7+opcmx728yKbOYCK
HQ8Cm4vjupoBeIJBz2GjLj+qqMSVAlKJnuKOCYRDxSrDfHJHXp18Oq3JNajD
hd3zNQ1iB/JBphjBw92/DLnZORkAdz6Hrh9LkDGnrk7eAeRgmtBA2r5TXJc8
/KidJHb+GpvaUSJZcE3gu3MMGyGgSfD/L/dZAgI/tLK/8k0s2kVDC3P2T2O6
ug/QXpWHLCuW5GTZLW/VIUZ28at6WILUMQ44Y6AEvsouw0VjLCxD+F6D6W1G
ucc6McGRdr0DGW+WZjvrojpXnDhKsY+vgFAYUqeXKY9h7tGj6ig3GW8cWMxB
QloeMaU9RumA7ZOxAEJJe5vujIErGLGdeNJI9S2nJUM/24r9t5DDArbjwgao
etdJh85mBSg9veHvrfXC8dVCIJHXPDmZh49vttxQBXEGI5yAKSpPxJmWUEOA
k7xBV0UlIwBeeYrx5kzJoQNjgARb3jFUi+gQNuPNyNUBfMxbN/xJicaOZ9By
cPbiaPUNF4b7sEygpTZGIdDytrUEHgzARN+mJU2UXWEeWAYeguLvabMR3CqW
n/vbyl8Cdf9Ba3c9zXmO67qKqbY/YnSC4a/VbkJt++1fDMGpIMOczsHg7pJT
JTCeI/omnAJPiJNewkiWmNMm4PchocAZRf1SyDu9zvHP8AWVFvCWqAUNsnhG
t+bjZrkoxKz+purfepIy7De5FuvXMgoEf/nhxquOeFvJ4bSUWVT2LXiZlYcu
X5ibou0nkWOdPddo9l+8UZjs3U56PQ8Cjzd/I8kfqptJvnzmn3Jdmf7tpfjY
bC/F1P4s8B9NVAFuYlPRcb27RthGOHtzQJi9suzq5iaYwbMAOptjCBI20g8z
USB4LeFnF7d2cCxPWgMcUEA7Oydh9qxSBV7UrTFk6+8/EOB2pjQCA04QRyyG
lfSJ0giKzFCGwBFxG3t27QReHkV5+iPNUpggW8hVcQ1kQ5nPm2cAVkYXB0tj
lVetTpseQJDkw0sWSL3ddbSgL+wiWpgMRTLlq4KnmLBMjr4FGrApLzFNpPhb
jbrkr7skKPGt330GpjNJICklduDSss2eAiPbNPXv+vH7NUjdTxyLfKpSfXke
3Yw9UiPFWFQZqN1V1EbDNIjCjCEZ6CC8zW1cSiUcdYkXY4kFzDzLoFzOOxCA
2qRNmYu3KDSv+ahZsGPufVH9aZyyHJKSI9ndOLAyDkaNvov5LkJYRgPllKbm
jzn6QfA76bhebSDUDGLr7YI/mrIbbzkn1UFxq1/vWrSwsQ5Kf+6HTmlSjvCD
EQJ+PpkrvWY9aU+u0RwH1jemkWhI8VKjhlhAOMsPFLhcfrdcybWdeNOzZK6C
pza/TSXRS4rKM8X+CFEZwIiRdBlRq6+thfuFH1l1maYUmASjDP1J8IfnM7dE
SDkferWLos2ca0PaOYaSKXkTSksq/lWN7P8TnfwXEo95t6XS6YFik5qZDPRe
SVHtob48y/3CP80VAVnuGgmWpCCqtquBxm+DMCOasqmQMm+dtasSpn+6wG8k
1+dDTeze9WwbSlCrXb+FN3gclcNvSZ7CB5rmiOHPeRkAa84oKb2qVG+ygic2
Z1e2MGwSubjhl3gjf/vqeqC2UAKAq6M/cxG+C0cdFuo10r22AxLsXbLQNZk9
vn3FiNxkSaPwfd1eF2mryJQVn0gQCpiPA8WkiXmB4Z9PO6T7NIGxauYb85Rf
dqM93pGRQaGqXN0xepNg5qqUX4yvolI9bEY0Q3VMnQsRHn0+T/fErb0+5YKw
4V2uuHEWmm+QIkTARBqmbaOsHfGab3Iq5lsqZDPzNUSn+chSrgUcYJpw5KMG
UiZaxJUW/j0bFTWNVhngjQPbmdW7AsYfch8tR2xKEspLwKf7kvA32IqBfN1Z
I0E4QjDfoU1LzxxX8omh7nnGd0bQRAlf9Ebj+oGS5F6AbxVgIC2pM1QTLn0k
95TLM/MEX86roLs1E0clkYLo+1+y5LX4Nax5DzqERzwettym8PJ3Wf9Cn5T6
GePBBRtQRRpaszWpBOHyB1fyitvcXD0q+lw4Azf336Wj/WhRZLmuoWfduoVt
ejqIgRyaKpeDt4ZNNBIp+3w2XK2xCnrBL8OBrPOJ+31XVgarPIXydx/JYfJZ
p7OoWgYXDQI3wjjscqJaPq1IuXkFZ+ZN4ENCGer8oDgxLEqRK4vX7tETnzZ/
xUiMtzP+LiYpnBXCw7AnqWXDIaE123o5AdRCXlx4JzJPjEF1aqAOyZY8zsaB
oFX/Hvbu4hbKH6FWA4r71KIv8gQZQ+4tn7se66/lcnQVWZ9OzDhM7WE8Onpn
QLsHeSNAAd381wH5UZbr1jKxy4Ec32hN0xjYjZhYVnQc65RyjvYMiJMSEy2o
UgHWIRqniidsCca9Zvdvp3oTb0giunFNwrI34c4S+Ihk//AEyYftLpOaKmM0
nU8HmZVchq7R6xz5mjOW9gUuKuOYhR2xEcMYQG0g2p2M/eYYQb5HSLqU/SST
1f/VW10+5YX23XtjX7R+tm4pyMSBzR+OQ5tDg9ch2B2Y/otfW/TplCs/esz7
l5yVz1F3PD/ynVmBbNeLe6t8kmaAhdGD5qfNVQfBZjydyCN3KMmb/TiwHsyE
sDi5LKpKunuTtkCFCPY8Z58iIcteLGmUu5K/ciFq06B7RxauR8KIkgTyME7D
1EQwmte3pnxsUB7gGpPU18OIYSA1GH0XHb4fWwshHm5HGaHFwSCUfvxP6v2l
H/YKTI5yHm6u+0LlOEhzhv5XBiu7KO0ZZnIVCxvpqnd/P0y6UUglA2v8jEbp
PO6/L1OBI/BD8qGgkzqMvTjama7M/Vf5KkHkCMIBJ7zaNDQCX+En25HZHy0f
zYmEUhbg92iLoojnGqqrw4fnxFShhFVR+CWCSIQ3BlpE2WkOs8BhRt23DcEs
VJ3f0e1O6aUmdKXzk8rIybs8xoJN5OLGD7z/mp8C+eNx+73QHpP4hPgEKR6M
MTSfHVlS6gOq8ZmSE1MDJMQ40tc993XscRVIQmFFokEohHKWdYMLFer1h9wr
7lMXFECdAd7Rc9WDU4NmtQy8eNtUc/cgi0SQ0E7stx+Yaq7jJzS4Xzydp5Q5
8ojQyTp4bDt3GAXg16G15/aKbjeeLMEYt8V4yysu+eBHtf3vmSV09cFdY04a
ME8cAUtazyv74V0YoW1Nc+R57SRS7wNMZiiYFtcQE+Vxai2yg7YHvleVM/32
VgEmiGT8Cbgi2s8jKU85OiJyf9NhKviy8Be0HMGFnXPSEEE7KQqadgfF8gP1
i5Icu/pOE9lN2qHOQ5tNThJaOHirStKcD2nA5n7UBf+AGsGCWjKjJuglu23L
tA25DR/OymV+7CVRCzDIg9gJHIQPTDfYGHhdfag9oslwFr2hX68JcQLfdvVV
v7ov+/mc51F5hjK0sQ7ImxAcweeKnUD/ToMGI0Jex7ytByHCrNDspP6l4KhL
vrJaHN5mD40BKhiPgDXJuoZwTKrHhvRghivISCWN20uEjlblpS69jqo2uiys
zzO/zG7Ax0egFo9r2RB8scaXYEIYaCPFoevcV3eBcwI64Geuc7Va7yc617ai
sods2PTW/qDd6Q4ub0yo0arS+3sPIT3STlrUW1TQg61YvA5pBvBjSuYGjAfR
gvImMBYOPrjtEvYzRn5BwzFOd6BKxE8Nl42O7bcgAjLHMS9ccziGm8ynpT27
vubDF8fMhnP0e74fjqe6u6wBZ9o0EW3xFJ4SAyJ8CGbXsOJoAslBpkRFAR7C
HYqj8whYnb+wHEcedZM6e4uUFlPstSDLPgFtg2AzDC8DgDparZINBDrsC2lm
NoG47z4Hhb7OIrQL1PmN8+4yBF7S8d7wL/0RrUrEoC4jxhZVgWDfrvd+aUp6
A0qM0SN5AGFxutV7XgZBddUmRfa0EYmpnrRyKEPBXFwfuLAtuA0kPrbY7m7A
tcRyKRbViaMZHKNk2R0xlIWypWtWc7ahmpIvvBqi/tKKwnTRqbyHbjWr99V8
B50nKo+OeWyzpWKuWqEn64hxOEp0yqubXX9jbHz7h+0duWONOKSlkyGGESyx
Ca4YTkI2lFL02A3tN01kgjwdebeCw5sApMrHPJ2lZwY+g5xM1UFg3HRxXtyK
MRR/cTrgN5Xr4KVKVss5JKzap3VTqSnGahSNffisgJdPCpqIW8CH3icC1bgP
kRRWbWSnnlaXgst4vlQvl42tMEIJiYknArjozrCXBkzIIUYUckXr3QUT3Bp/
WMn3kuUFLVtGPjQ8MaEJkgWaz+bZHC0zQynWPJYWgW8aXKNd1fL0xKgoBHhD
vixwT7PZNohf8dkzr0uYSTIFPYhZcygr9ksCcvSfrWAmSV9vO1a8S2MDYX8H
Fikcu5xhdmEdS9/Fkz6mAajSVHl33HhcDpAQzqX8GLOpOvuFBpzhZoksjXJp
mVpO40gRfYJkitiQGDWHE2/j0Cviz3YuYXRYlLmOIo0aQtLiX6Ds440RT1Me
hKcbos4wLLKoOBPbYQ9GmAAkDBMmEVn7KaQ1QgYZTzer48fPCIkLWwo422LD
c8+s+zuOA2ST+WdkFehUhACHeLY5ZYU32WsLCyYLJInNNlneAzjXsFMwmRqP
79453PNkZVcrC5yGl7w+Cctjy8f96qmrRfjN69piuxF1oHT9w4JTB0erdF3t
V+5RiCwqnMxGeyJ311r72VxsaJer7TpUPrvltCL10zlTNTgtv/xMdUCeymzt
mXTzJ6gun8djuRf9Z2G/qRrUL1Sn6MeUwjRdgZhaaStZxEp65k1GAr+vFzJn
OEP5Fogv4odfQEyPwxrWMWFWxH7FBoVgcr+5N3fdpuOLCnK6uSilP1VEPXR/
DsZAl4n98mY8b2OKQuI/8dVzp2dIB0xzwltFZSB0a8RE+G4dqYt9xFqKEyBQ
U4m/stebuDxbOQAJbZ0Brke+4gDujL4XFppY4KS7rHkw4kdgP3CL00inFykS
SEOoBoEKX8jg1ckKPO/XW350lZYupuParivMwjs2aG8KzL3e1+4dwsx12MQT
2U0fmMDh8NWOmu/RXkrwV2qvF1HDsMwIqheNiqYRz6UZmhKQyAspx5oI0OyU
tVyuEDW0l5cFBfRVYXUAyYeIIlUJLifV+QytaSQqWcshb7/N7dgzQZxx7xWG
HzpK/ZVWuXiwO/AAUnlPknMmnQhND/qMarpuFCf44V0Od+/ZJonbgl4pJ9KR
2oc3xrNpy4TYiEt5hvvSlwnliJoM2M3BXbhQxkBmRoCjGQiG/dyfuORH8Z/L
zSv0ouxjiUcn3F3jqe9mNIHfISVxI031mD+pA3vEPI2YGVc4+kzXQ1Qn5j9d
LxbpdLgVKC0E4oGkH8BxF3GRkuLnlktSf+YzEFC9FTnfwiXYBaFqJzaXfjaN
qyWhbD5pZeHlRgBWdq0T9A5byCNnsvtaBuUZubyNLFIezi6a9xomU9UD2lom
eYgSM+SHSQAPbpCe2ZB+ulqYu8phiuzY2OH4xtKAkrljseq2VzU8mGMFLXc/
zaYgCiEaDMoTKQcGAKVyXkXwdHeLOPgBY4GXE8u9ho5ywHnVA6qL1bVy+73a
BB0wpbjjK08NueQ5FabV+QQUn+7uRq0nNAIo+LFhyHobgNfVRT/UaWeUZ7XI
o0rRibzXOOEozxjU5Hb6CC9pbiUT9M6Ol+BubF6B8i0Uaokg/CneanvFpFp/
qpOkN/FsxO5U6VK0yVklRdf33MgE8XBuvLw7mKGrsJIPCEb6RBLua17E5/QY
lIgmTv3jeeD/jg9UEBP1g1BHbJOif6KSLu321U2zOOS6vxVFaWsEpIzxL6sT
0ieptpuj/8hdcC1HBdHBXmJ/6S/Ot5guYU9l3BxzMPYu+LKAShCR2ouqaTTR
VV+blaZ25us8CYmG3Bi7gZR6W4SkNxiuO4Tta87olCSW0+O4APNj61yj5iWP
ke2O6rxc9UDY3u81ZeVHx0OBWy/2FDmyjdaJN8Xex7+MNcpHBdVlQqVMqJg9
bcCpu/MbXgX18keFH6KLWRqv98Vagmk3O9DIQi8Y7G1w4oicp7cUvsing2YN
lMaXdIYLu6qcT0Je4Bbr9h8JtdL9t1QDcUvHXNOII8fllUVe2aFiDYcxqGwi
cDvJpytYGkzt4aQlyvlnTMCJI2YKph+EGL98aZLVagKSgE6+w+64wbx4Tfi1
pUuhUhgCzS5nLbSJpI3J5TlkaB7EGxhg1pO7ISFpH1Nz5Bh7MmE9iVXCwlTj
lRBzL5owSSj2lFNV1s5skbX7dL89+boY0XVKSW1KHgH/o0kaXg492KOlkglD
YFMIOnS4fIspNGh9riBN9jXHj3ZrrL7yjvemn45ijUuoR8rEt7aAJ3fVwPr6
6jCFCU6va0iC7s0b3HCHxQTkiqa8UeH/rHvDzK42VFZqKbqS9g9HQdev6J4+
QCxfCD8ecUYEA3oB8M65eWYKe1i6kh5vhTTapcDWjd3lHZ5yxAV7lZv+VpYs
ANdXJ+o8tE7cR/B4vwypv06WdkRqenzhvW2qFu5n9JU1tIZU5lEiupDknLS7
YG8sSadourSgxulNiS6XHdYNS4uZh6K2srX0BFGh7t34dtZWiSXkxry3q1yp
+2UnGaI6KfnD9nBvzKswR7EkZFWveA06F46KSYvMXuKU82CYtiBVKU26gBbF
bwzTxxUoWjlUn4HYoM4kyLMxrEl//t3Bmfwn47ZqRC4Z0lhtVxPvb+vGd5ry
qdxSC00z5TjJ+XxHx5+TqFKwDxcR8zYNFfk5elLPS3bRopWdvklSw7lJWrh8
ImE2pUnLQ1xAu/yVKieurWo8V3XqXc4w9Qkg2+A7xHTIKy4IRa9i2pzWMLyV
/hO9hEFaXIf68fVNaHxIelb5Kwz25IP0ZT+Fh1vG3mC/qB8V2eSxo6uz1xDD
Y3c4rDW9hONH1pKqVCEYNf6nWn/MrwLqo/5ZdixM0lDwF/vcbfbwNMkOf5Z9
qA2Cbz8DuhH8WYIFzu0C6/YUpi1sq8YDWPTNdAcQdGN5bzmuM3OtpTZ5ZnRs
KwY008qD6Rny8tPRAu95UYEzwrpXnVfPLVbgnWGLAT0HTlMqDTqe80lNRGz+
wax9xP4IPmvRy2fCRj9L0mAOdwk17QkPQGpUZfsBtBBBwTvfmS1N4lLJX8TQ
cxF6eBn6dHaJ1AxhexlDwD7INS87s3+nqSzbewugfH34lg7wq7UzvVapt1Ft
lMz8/8xW9sZ+wc/hr3255GQ/dKAl9x4aI/IYg0d4vhhLlJ2ZcOd9cReoV4IB
5Kw1KthtOn+9LpaD6YzLILjziZGr1d3bOCvif4RXkZhWcjLTVlnDZpQDO1n+
RNzCgGKLmt6xAUg3ecRAiYC/4QFaZX9zEyRKa03O2dW/Le39Zw4TYWfqHRAd
YuUYvJDdmhXcpkwwDfn+CAGmB7tKkcvyx+RN2eWVmOki1k32oeGSsF7fb1cV
NQAyPkEimlOY2tFbrmyz73KUIcDcCIokRD/WisnjEOQ22CXIRGocdHVaL6Ml
8CQ5uD1MBLa5s+0cNhRbzsZv8YngUIYCubQ1hZtukKpMHFyPRaRzmMNAy1sL
aWDL/oeq2O4RvTK90uk4Z2GPHakHDB1SrUoPBBWON8yzOToB8IL9L3dAY10i
zL5xjwY8j+nfCL57kRbIfuXFfeWAILQnlHF2wUrv9cNTWr71p3Q+9UrpBAdw
aU8oGBAm4OkS1Ny34Qfdlyi213yfsHVx6U4oSA8OXX6q6BULj0Ry3GX/omA6
GqtZGMn+VJnmKBlo0MFvkLVYNB3nXyJgW8ZM2SbRcofOMxipAUAc6a7s9It6
R1Ho7ldcAX0LppmeKIGYyCZdLpN4s/8UG7dbCI4J7ORYy10tulP8IAERJ8yG
AT+LRMXTOBOIte/M4uvj8/8TJdAuh2D3BWJ8Pa7WadRMnZLUxn70tjjzgSRn
2tM+CGNhwduoDVMLFDEORAGmZFrB0Y6myEa9LzCdP0EHXRoZ1K4lnWxY1zsM
LNAKtKiEXBblh5hiwodnoJji0lk+GDe5ESzbk9iQau7kflAswugaQGevNSUP
aKH8PE4cViUh+zAkJM4IxisN95/uOHQlNSHHi/iN8bTTKINPgj8Ejj5C2WRQ
mvPVjdFMsnzqFC/sCZni3KTXQPwQrusaGpkjVV56HyVXBcKyTfAYsz3k1RDz
W+YjgfYZ+JQU+0nZSF/lSguAy6isIoMy6swi9ddC7/26xkaHheThDj8YAf9s
fi9nUZXUdbDK3WeO5nDkzL3+nn+YvixxX/XC4RZkl5M5B8/g2ZohjqEM7K0k
KokR267tc/MTXP12JB4NxuHABOCSr5rWV1TzgLvCBZBn+uk4HEW2R5uIS0Li
Q8M1/z7P4dpZahSJ125EJKRqjM12BXWlfJwYa16R8NktRenm+YsOoBZTZBXf
R8n6QAlbL46DC8Izh5jOpSPlWWcwQQ0IRw5xbGGEqODtXvvjJXg8ujdYlTAl
IyloX3tNlxOT0MnE3VXjCWgVMHUaX4UbFEU+55tI+a7353JT21jwvTE2W4gh
te0l1+CXnob6RHd/dDgGod+wot9RO4Uf6KVbNl9Lcgm+1YTXwTWqdPvsZQ9f
fSVaipo+YSCryu4fV+CEY9uqIrKDqiX46zXb9vVt2sMu8ASclOjGlrqwst+q
JCCQEBweZbihonTakR7ss9E6ZVeJqqwWH8M7wfIubffCLicsyh5U3qXyhje4
c3OzBd0hToyXP4KlCW1TeyUBYiOaqqL7dWeKcRkg/YqCPSvVnODyvbZM+I8e
Yzi7gFe7sSRK/MWHyiFybjo3zmqH0WCJ9/zbQylE2vOvVUtLX6kqJGaRASjB
mcenEqloy5i0zyz7C1t1meK3Ho4RrWibvASy/krmbW80FrLDegpmPsMZZ1N7
uErUKJ1+VK/u3bAzGATP0pBYXaUyZ+Kbqk6BIES36Tli9MBXMx8RVuVD8rel
AT4lcb6DGbTD+C3y9a0EJYeVH5/TcxrHzV5RThP/S5lVtVvT1uG47gypQqIR
VpJvn6KqoUkB0gpGyxZE3iuKqgSGkcvQ0Vnf39orXzzBPzcTh7uLBA3t84pL
PWLuHXK62jL0ZGZnrtr3r3i8EdN2g7UAcjGIMM/OLDXQCx3+TcU52sQRpv2s
1HwLZW3HAq2hezTNvT73PJVZ+84j47/k8Otveq+LFo/9ALkbJCmOzKpkwDxU
lLv9kI85QJntiTRXzbzyPcLVBnm4CIzlB1nXu0V5/nBdMCJEr2MOFdmIfXNV
NDLuUyXEjxxMbrS6hzFKVRRVcBayfMJoIAX+ByUY+wZRyvr3q0v8Q3lJklpI
v7wiJe89HQjwm7oz1Jtz96v/U+GMShV1TtkRjHGddn6qtOKFe6c3KoMwMY17
OZeYL0h+lnjzLYgVdpov2xuldgPSj1xogUlFkF+X37JjRP1z1FGJKBeUPUfs
3V27FcuRz3AxZccjK+0LDjFXGGoU66bLb2kvGuMNqoGZA6l9xM7QAQ/NNLTu
qLZEsyhmtFZW29dqPoJySJkFzvuPIXuZARu72WWrzlRlQ7HBUpOqJ4ZDaKpO
Myu5ufWP6t4TikEn1mWBMd2BUGelXfrCSx6SmxkmLAXxHcVUkqsCoKwEhUBc
BBC2d+oYHwOtxunidXtdDNYDsUDcQFEQEiMZjigR5Q43gKB9Wd+GwWTV5LLt
lqLZR1Fu2lutr8IDTHw3F+1NQd+WOF0PI0Ve+Qc/khRqkqhfhzEicLjiVsoC
P+OiB0iXaUwuf7knU6XSTPw31DmjsI4Za1Nw6v7elSdEVP36xvMfV+usGyfz
btm4QYB1jF+Gx3M5W022zgpPZy+sWYUoHte7b6udt6NfmZSxIftiOe24aQOc
+bzy7mmD2MdYdjydkX6wymEn/fbuZbogTd2PEuj8Pjajtad68KviGP9p+5sq
7N3c2IyHPTP9dsjZ7Lj81eu+dMjkrKPaF1xcUKFKhp45PahMcw1J8KNioEWE
cVfDrl882CpnoRqC7p4XpP/5RP9+ISfeGdTNyBFsHWryDLBpxaRLx/aAmR5a
/wZKHDgpWTMPb4Gd/e/PTRuBXXSmb43xODM3OtDLWkv/XN14kmV+KYIyHLSf
H1RNa5+zOb86WDJKel/52dA2BU9vtv3e34y6XkDfJ/pybkJAJXCd3I4Qnoi+
es0hsP27CfgSdKNZH2tEd28FMYOhfmcuRcVVq4v69FRfMSLOIrk8xuMqwZ9D
ZbchkEODNLnBoSINq6pVckEGXBakhDEa7piILjbY1rq+r3152Ut5SAQTJPom
d+FzItAef0eW2J70dXK1R9eMaKZduaYKmMyV0Av7+sB+dDhT1+R3XKP5rsSu
8DCcr0OV+feeRxT4nMYlw6xODU5v7NEb0Cky/lcSSDcNIMvuKy42i4KzLu14
7u197pLN5u1hXyTn8AMwRg8vAXIfK07DmFwtPL91J/QFlLbk+UXOdQuAoZF1
y3kgv8XSnjnquDBBHbhePwJ62vVmXUWLdrM4kxAFXOPUO3U4XzcAqosr9lPv
zqHZcIwf6emOfkpRFE1Co9lScrS9WBGO9YF7OEK0EOOQhwfRBZqPmfuN8jXx
ZUy/s1re0KhkewuKO7Xx/w/pCufunBLPGoL3oxK27VkTI9uvMZfwe5M77uQ9
zsxcaJYK9CLVn2Wf6i++esakDLwoxugJEythJ+3tPOgwYGKkkeQYTc0i+Alg
9he3tvwJwcN2ShxlWhbhNdht6jH5+GbLGAyDpzTujxUaI1ciIVSJc0VDKN+d
wm8z2jQAdo8N7snkAqBV01zq1RqreE5pu/9OX1iNDqk/RyOSwMc8s74VAsj6
+lUGT03IULKUeQ/U5mBUqO7X0SU76RyH04wPYKLAzNQ3qRS9lOQ40o8JMN5j
1MvxQhIY/cPfQ4so1FcHZ4o2i+rNwV3yuG2Q/TIwNKThTYvlpoFwM2wKnLB/
N+HrY1Id76ObHravVEKknRjeKz7MkIF74vS37s5+u6oXCHq8PTCHA0G3Wrv7
HvuW8dUD0n7xoBKE9Ay+6m1+WEtZnQlLTjqQCJOSn3H2l/FCZvKJSIwh5vgl
r0tUvE6tnQEmFgOOXozORy4jWw2wfcUtMfirJxuYVSdUl0ZYg7td6lgEPhfp
kT+AD+ll8tvDkTp6WZXD9VpDjzQRnGqBUJfl4tlq8EACI59fPFOH5T2xWH01
+ox6ZPY7GA3rPdEjph2N3IbzW6reJTtp5HdDRH66EU/C/OEyI/9JHwi3WY8h
NEaAbSMQX5olk3/uTCyezuypZlr+Wqoni+2A6mriAqmNqul0K3l7JhvJCvS3
mmufrlsq7eVT11BQpBodKsJAzmVD8Qkgqo7YfCSBQ5mphGugNDcRlGQH0bIo
SIn/EnY7MuJe+AsQ2Q4Ysummg4RFKovSsLf+B/o6etTXA9jb7TmiYPnUm1SW
nC3VCWS74D7A2kC8nDIHmPjzMT+nZTHL0k+XK9/z+q0Ep2Xuz7TAQR/ucaEz
OYtxDEPPPRvufo2W0Eiq3MijfG7Wig4mkVaAtHk7a+R1Bc+xIWm6HA1DMJTM
1SpmXIYeIXDdFBfX9NxXGDlPqk+TqYa79L69X4LmRhVCfWUayBb3nAqkK9yi
XIE/egTj9RC34oPsu2fdQeGqB95CfIWn//Igu4C9m86Lk259nNl8Z1IBvA50
NtY8gCfFu57h5apdCYMkD8BG9hQzA1uc9gqBF+742/73dieU3MiN1GOvLxwi
1p/LgGWYDISCqHkHUOt+ad2PTTLKD6MhNHwcDshe/Lv7nNcb10DpISzvjM9M
eZmIbGW0t5xLQAUQv0/Kbq0/xCD71FtWjEniCWZuxJHdE0w2KfAPXhS8wquI
A69SCqRPeVsS8Yk3Tq3IiQN38SK6tXnqnto7CyNLvNT+q/u4MPsxp3YEPcdy
0eLT++8BuCgnMyfeQr1doHOnS/UKWHArpBFnsIq4WlpQnyKGctgLa6JbWzrk
K8yeQ/YGeTCXysazr5uH2NVsQVMGRNzgHsazYq7fVyMiEzoPCc7hPh/T/Ht0
SLv5Sg7cxGqd262axiQLaCX1RDGk7LtYaDGxmY+HtCN+523NWjOAsUVm/XeU
4DPNSgE3zQce7/UP3+aQb2acgofOtonaMC7FZmPYhTVjqsnS69LdUQPN83qp
pTNFnoR1GoYS4/zSmewyBpNJgECE88wwrAH+ov6XRicQDttbkf7Z8ZCzMtnQ
wsTxUJLSsXa1rd01YTwLeZuFlXXq3cl9cUZTbBuv55FS7Tl98qXfUrf6saqR
bjHklNJqfXlDANvH4yRwpyIVeY+TCuaZaJX4bHjS4uv/WTjs6E/gJ8wYmutE
BdwezYMxAtTzQzlxq0LOZKqlZ46BrcnMC2EUdCF7R5922z+UuncqJmzdVFMU
f4iWQOi4VSsKMBj7NFRDVuZEz9aPyyPj8An31arJyfEm9k2Cw0lBoerXyqib
3PidwKmGc7srriOJuYkabLQZAAN2I3RRKMzg4cSJ4O+Glr4X9F0e17LCLfep
RFYdhI+ZO0f0LcBN7kF73YfzxXcig16l1xTX6ZugqD4Qxq4YoCIJjyyEWqcv
u7bNsaSBJF/07S2ZheVX3VhsFfMDQOVETfamdt3MXAWpy7pvF0PPYyPjjbFf
D3DQRHHIaa6u6LQ+tVIBmw2xSkQzwVIUiJfEPrimTEGJeLggEKgGuJeupvSH
iEkU6jKB6h0qe0DGv74BbyEFQSvH3BSdtwUdlwf3i85NXb4PyniwDQ1psrL2
XmRo4kyO8Do71pI+286UsK29qF1gqBdxTe4lM44rcan0DgcZJ76S3nvWh98o
LY7kusAw5Dl0WNp7ZrLo3TGFbOb6R874qzyski7ljJxcs64jw7WCRE5cudmD
sg3ZSQG7KUVKvqC+0qoW4mbJkgW4fDIcvTD6l5k/koP6rX1GoyJv0VFwtfpZ
TH8qFjW/pWM+vwE6s/CxtsL/fE5Ycih5EqGo2Xp3SuxbVbz7HSGojApBgEdr
ySn7lYhcGmBGs1wTYlk0PzsFvJvNFtXxQwwGCC2SH8uKvpRwjklhUvcmxR9R
3xOGgO2CH3bhXQiMwCs0qDPXzvSiEUrLaZSIE0Po5OjQ1o1byv7L5lDUkhuR
ybCz4LoxupQZoWvb4t4cAoeIj+pa2+cyFjb7LalZlDOdAD3N8Fz6ECJ/BHjn
KKAl/Z0gorbzY52MHcnnVXEHWes2jQb6OFWbKEZiXbdILRh0KAyyIrvcZPqf
roMvkwLU2H8dCw83BqMDQF4CTDuaL5XW5VEFiZKXpr0X/LnRFCuW66XR/CRw
K33HQg57mzjD1T6dMwHLKGvxUWQAvXOQ80wz8mgqAexOYgFdTr5PY93VRTQS
j4TeBQfxui9ZCpmfW+WoUGew+wThltPc15+gFAfDdeb94movCvDsWAsexsS1
z2zO4Ar5zWrbU1kA3XZqrWEsVaOKCb326m3Xc19yB1JsSuRxGWeDq82gMEyl
TCYu4dXO1GPGcq7NFx3b3WDxrp2/67CuKLN0Iod2XSK0ukkk0tobLUKr7JoN
AtUYrWISG9mWAuYVb8HKLvRsDnjFux4pvKCiTW6OGfig5pMXXRR3DZQkk0ho
Ci+64i+UwOM7yVEX3ICeX+vlHI7tTKFi9vLnxUqv30jQWC/ygFPD637UimzL
czQI0GbRdJX1WL2s0gByxWicYbDLKhiaQCLCZK7NdrwvdmtcZoJzD3GzkdnB
8nCR3YlFMjjq8/o4kSTm6AG6++fIuYX77XW0nnago4XKJN4azAeTncp7/AUB
FC9t/NLHZtUZUwSuU9QIvPEer64CG7eLjhYPCU6a4MSgVrfit7UttU6RFKnK
BQL3333rIiPZc1Unz2ScCkdoD94PVy0GqZmqOblHkymo324zqOO/cATQxC1l
qLvYgGiGzoFUjYiBOCQX7cwJ5e6XioftGPOC6UbBDQ5cYpFbH1lT5+eajBSW
WKe3RrXQEHdotoo6INwEhrWbeXXus8cc3/UzJolQTiionBT8aB2ccN7G2IiT
UVScd5KAcG2sH+RoYt6h9KGgJEtaBU8H/6+IazCr58m8c4DbzVffDQt09kll
2fGaJb0/p92b4q/gYCXWtsfPe97oHnE10uMeY03C7GFJP+gzJPQd/+nJ0AFl
pUhJvjt2eMnzuIfTmYACjDLR+EhMYwecAl1+EVWlG2ui8tmELxSaxLdiT+Bb
aYOIx/8p3/MT/slpfylGjdSEn5IVXM21E7Rd/p5wW/dgOcExGJ8vKu1imHhc
1ly8JRh28bKzD09E9W2gig2/ELnCCfwYDUHHByN1NFR5NdMN3J3pfepi+y/+
cWyIMoljm4A+eWrXjZisXjDivtnI8CL49Nez/VVy8uJqahulq5WPY5q/fqYa
t0mu1UMw8nsZOgOYJeKCYsG+8233h1og+rVaL+mmSVTV5GU5YOG7SOK/gVIt
oHYf0QW61GZnNdHs665sJk+ROHlJ7XxL73TlIOy1mCWj7gkI7LZ93UMq8eNA
nqKoMNAy98eOIng8oUSJg6y+tcvFoEc7jpHzuEys3/XdaWMpgTV2xDw4n45e
XZhdI7dSa7AdGHIi/mrawkqsMZIfYtyg/XztLyAh8MNe0psmaE4l4dG4v+iB
Kkq7MNA8zUkiiByaEhYLKcg4qmNpNYKYcrJzCPS67CeSVQ9jqVNLDRAQ87+8
/+qXDesnTnWo9tkKOV9T8Qsji2IyPftF5spI8xORc5eq9zkmejayxyQU5Cch
FhyEUOV4lz4wfzBjaIcc83up7Q5RBVIcAWlqIvkXQyLXFoHBlGPKZmwSQI5Z
rGrjSulf2QzWQWTdo0cSdeoaMFAnC33/MqQzuCbcRYURkfZTYRTLX/yluN1b
8rOE75Q3hc0ueGtuDVIMVfpFZgvJAnHqtpVXiicDWiEvTo1BFOjMgGl3ggrH
1If6JGH9k/T22N6AavW3WLdNlEeEkBY9hF94Ct4HXsz2RSK6TNUQ/wQqWHtz
j1MYFpg2idcA7BqGJ0lRqWz7hbLvY2jhzdAzrewF3x9O0WtmizAKv/ZN5LO7
qILT3CP1iOkjdz6uAjHikb7v4FA4TtyF3nUM/++SbkJHYizOqCHcInrGoGux
zLBeBBeHjGciuLM+NldL8eAHM5j8AdLoi3q/Zo48r/E9t6VVsta4ezLH6nHx
TyvsbqiYKyW6Zv2BUQjWFrjR8YxCaoawuVGBTW+hZ03gTQjhc0zbbLsD/eb8
KoSeBnvAwl5Yl9sAdFQ6jMubs/NKCZR1ppBRVsa2v52lPIeXDCVvXAwhjoDw
RYjem4GcDReKmveDQljd0I5TcPKlB76bcHD4mWP6pQ6UmOaY3LL4Amft5T4a
VyHRutFSRGK+/AyWM+g4HUnqg+qqeXEbwudzDUJyVMsKf7eU2aEmmdkSI/01
bIP/Ag8300k2Y196qInF1jvT8F5gAI94mYz8/Qf0RNs2QpqX95jUiGuIsfve
iQekLlwTWgwavBF0bmEf2s15yle5Tz5ZPltRZP0KkX5aNsZvG6ckVcF00dMv
saxERmLeX/B2YQ+U6EcCL0JU/e2JRIuuFYbNGwyuwOMQmw/fNqV90AIbSpbW
h+/5LKwdgSy+DaImvasl5yxUtZQs4l4bd95+5z6Dq+GPx5gvBnS0ASeMz5K6
QjPJWs7jq1mdqfJIP96BjxoM4IdWl5LNobHEKFgvag+Leq8bJJsK2e2Znj4T
BAXzT/HE85EePw/32oH+2kRD1+3QWoruCY9xJ1ZBmLvPwFvX+31HaRVfKxmP
vVMMgr9Y4edJHn8+E/ZWQMTSGmuhn8IHQLYhAmLrjVg1MwgHPnUpwKyvcLiR
teooqlgDlcx06ZBRZirwdRRUvaMcI9gV9S/gtTzrwMnSplkKjN1GCFMbzeLn
8sTpTK8LB98borR9Q7ok+miSbeKH+SU7k2wadkFqRd4eTmoqFLGXg0vCIm6B
RZDw9GMeZpqiNS69sGrvLU1y0GUsdOnD4RgXu32no+yj4kzUBthQs8ufDcTM
SSqdXCpzjoA7lMj2aC6TR5fj6kQ8YV57ExcWU8yiJaf6nPHTDYLNbJiZMr/u
GDAoMherYDaPPSdGditX/uqwQ3ukNaIzRyvuvYngzY8u6CkXG6Jz3f83SD+N
dL6YyPfEVmU9CxH17JfLOfoFljkOHtnqEBnaBfoLwPqOLqt/A2uDRCiaxzns
hxs+4f0K6VWGH1lnNbt7ontOLBDDOvJnOBai/+aVFsRWw95ZUMEE+z7TbgZW
5lEGjVZDNV0XWSkOItNRABtJO4/l/drNKdCWRibUUab21BsRKR7aV5o5gqHy
h7rnYxQ3dedNvxRvo58gWvMObLL9qaH2h+10S66bzENtCavo4zf2GYoeWPkL
LsWEGvuh+k9Hbi/CLkHNRn5peYsgT8HpV8flHBEEUmoyM/88hCWDcUp/3/kN
U6M/HbBb5h2Z3r9tO+BSeZeP3IF6LTQ5rFlQLrE/o4SmOwnY+A+ngBFhrDq3
sMe/1ZjW53LJHXPraqmp4dtcfRyty7rRB2wfHhSK4pgsVFGv4wxbWDffzkDZ
ddUKjgSef+d5aiXkB9uo9H+YsYGr7Al54P9XKb8iF+fBePoNDBbzYEUkH/Ia
s6PGrhCaq2QOSwbvXZNnWSd3wl2bq81JVykpAI4UMBeGnma1x5x3P0vbX9YG
rfMppRPk4e101LxvL48edCmFgf5XUq/c32uOu16ky9Hubg3sUDQzR7LEjte1
7ZjVq0mtFPeLNKlf6HFA8XC9u7Lgkhv2T5RLVXvbVNaZ049+KvQMtEc/EHfc
cmiLeXkEFb7SEiyfgtY1xvbf5VvQ35ORHSLBElidI+5i5hnbNz/ipxWog5kK
RQX+y5DQMi6XnhQDKzOZ3vq34oYugTexTIHIptG9ysjNXuGNT99VJJJG5JW+
6H+4j2FTMGdNfamFndV4hnxgvtubaqyBE51a2HP++efyOzAeW3215uoVFBT5
ZJuPwC2GaPCgCd74DStxug3hXxb3eMRXauiuzzOPlxlEkYyHSAekkecHNPRj
KCMTY9/SaHzIeG4DqfNJGhg7mlZIovhz9S+F1AYylcOyA7vLdxLmOoC0rspB
XMkVLI7SsOb8RF56p3RVKDJnb1uT/ZSMXQwM+2gu4g4k20UWPJHW3ka3Zwc5
We9bQ2hZMX/DsKXE5h4KKxnpB+w6Qy2wfSqFh3QYb81gLtp6x2Ompn9prOdh
PtqxDwdBvMICFmzOeqMTeMxfLMcmgZOsecXg/j7Z4IdHkWCNGEa3ZEARG/lY
op5PiqJeU4Ytop5R+i8QJI+WBxb9y6ZWdCbtkHmKJZ/HmkkvASnc+zcbCQ8+
p8AfMemLYaNX4P9V2ewH3/58PWHXKRCnhujOXmlTDHJ1vnkubAmT4AYLAN1l
Wek6ZzwzbYLIo2/mwt57Q9VWEvUkBdOhh0K+Av0Y/gBSyoXW2MM0KwodF5+p
4M+nUwp6qcLQM/uYZvjrd3By0DzLsmuiXOLXglcomy+yZnaGFmeJ5+BOAXfT
uXqJpT4qR1mmOfBg5eUDdS+/GSlK8oAiUDddamE1qkQe7tWnO4ooDJhw+s0t
duVX3VwtJWgbMWN9B0o1CAvRAJ42i1YbQAkcoNW4T4e7vrJM5hDIRB9hEkHg
MbOqKQbFcFW0UFeeCYvXC4L7o70X05rr5g2epHtd9cuWv/f4ScDcgvu+6jFV
kH8jjNGTQzizpOFwS0NUBE18JXi5UT/A0THVhwm2Z3ne5uWINcfHrekxC28m
ibQFLKlhkTLJU0M90X47zS2Z8O6/fMfSH6jCfkZsculMCMv6uOx5Ig+5uSPQ
b51rNzt0loyQEAckBCl64erPy4BHWLB0bWIGWixvwsvXz8bRbB4Hnjru1rO4
JQdns2HCB2IqqiJApGCoXTDs72Lh1x1KfFbzFuXbV9B3og5LzrF/uMjnl3dO
qkxdh2g2h+tDf4qbyrJyYRWJBj01L04puYrJ7lo3EtMRr4cPWy43cztoMMXE
mBXWS4VFYSox8kC/ZFN7y2qgi368T2fkQf2f9YOoB5LIg1/U7C2earH2wz6r
ir9kAPFJL6mQXFkD8nsJxyIdpwUmTYFxA1gQkziHpHlwnC/aAazEFfJFPHj9
fZe7HuP/7wLCpuoeQPnfZu1MlB2/suxQxAf7BWAaIc+ghYE5h/l9TFlxKUiz
n3UOTMhrjCkFklrj2Qp/p72q/EMb47JBI62M0WwWWzoO5Dq+T6C/rWP6lV3H
fFhBk4EEE39Fan72/bZ2adWPFIKDTgX8DDNatA3NNIsYZTB2rQudy40B3Rd/
3biVRlIm4/fry2nnyBR5UgaYV4sdEJwtEJ2+HX2kPoSSd/azVsy542SXgJP/
gvEgZMMb5ZooAPMKMi63ywUKbmSOMEPHho8U/D0mDJ9sxI2HZiw4Gn7Qp19l
z3mDMz14ou/qDmYtQo1UjPVnuTdIg3m7lCtxBfmO0ZGvaagqNBjb3B4tOewa
7O9+qcxy6ykk24+5fjxKE8BSYWv01K9kNedXuB2mYAri49qTj16L+Ha7F6B/
k79fXKMXcAE6q7PIBAxFyt9aHI265kGg4UzWzH+mnRiJI8Hf6FkdwK4732hk
+8hkN5AYtqaAz+gWf4SFGsJ4dmeI7htCn5oV5QVAQMnY6MJDzOfoCbTcXoWq
BlEfYln+rVbaHy8vhLCUuZ2Gfe58YzR/rczBVRVT0gMifRxrWfPMky7uqZPF
WpPDj44fJipjrUkonzlrDSRB3oe9ETiMva8raksLoLewP2H/uK0QjAgihVii
e0RBpftBqPuOfUrXDc/7DhPsaIURrX4TBvHXd7NeGUymnHvO67aKiHXa12mN
B1XQitTWaF40DzoMv9r6sAyXuAHtiv+evv2XFrcH0kA6PrhTFBJtIDNBhpRo
lxIDKBzBD7rVwnr1qJDv5rulEbcbvOulHriIC5rmnRo10lR9ilSnmWJZFX7x
+714/6hQQH7jjXUFc2ewCzRRF5Dtehg9njPlS0Ddsn+tJb1f9JsTn8OIbdmL
7nAj7nDmdK5/Shre9fw4vwxhsR2PsfolGVdsSV18oYI7WHW2KXzPpOGk+1M/
x75XdpbU56KsfnaVEciVtkqhJZiTLMmW5HBhhIs39qdXusCX+KfBEosa/Eh8
2gmpTKqwpMuDUEYHJyPGkUj9ip1Xgk1vK/BEZdxJg8hw7IgUA0UKCZx+Vr55
SvnkdPw4w1GsSdhCeYjGRRJbY2byz595HLEEnEtPGHLJ8w0L4zZPND/wvzMX
j6wd2xl2qkD5xxfKaq23L4S2Xg3RiZJaW+wxG8pdpqO3obLBSvIjxSAmA8ri
Gx7avzz2wJZCOk3R4Ble4WgAFQx63RcPT2o9vOCoWisQwIzxUD6rhOmLHqCv
tYxMSbz28UhXe8oCud7RLDx7gTepM4/eMPzmiWaCXk3tORgw2cpZCWLxk2PX
jv/omSwy+uPkWlyb7ky30LvgYujDSMkwz68y3X0aKKOHTHeusX1LGulkEwVq
mX7q7nQVyUhCRz2WHCWP5CVVFBlcUkiVDfKoyK8341HMgvGLxqyBwRJPCNgq
aOfCg+i4LjGajUVtasiXR6f731in+ukyxhVXCqAZYzVJlzddFgLjzQ5bRtPv
O/lCJr0ADWMgF69ZZV9inTtvOYgGBzrEm2MbJdX62TV5uo8qpq0yjIUfA1n+
my9Ov3Bz1mPCr92pcIh1uIIu5TVfmwqFV9rxdgLgrUJej+uzKEsBAHOy1TL/
Nu1u4UVTmVpi1W8jPL5jdsDbqYt7FvuxyIlpXQawcF59T95B2+EzlDX7qqsO
n/DIIDDYNs7kAHMqyoZ5fa4s1hw57Cqa5u1QN+XRNGng6M6JpiC2na161ATg
d/GYMRfQPgUhONKgj4B6D4xlyAwIlduIagJnkpYxlNZAE+rM797PhCjTaABl
adfsN/bhZ+td5l/7zQHKNNvyG9RTrzRnMlultu6ayG8bt1jcrTAiqiSuA+CP
UDsh5kG8GcKqe3LbqgqncLUojZf+0IwnfwvB29NoYBdNQ1tYys6J5H5ToImU
u63mG9Zl1biQDjZkQ/wjuci7kBCtv8YImIsUls192Fyt3Ncl8Bt9J1ixNzE2
qC8GUUJrFJq2XTIP5ymZsZNIyMYH0Gmdv42CfCODbA36Cf14qFIOgkxa7Kqs
PIFaeaVHFE1US6/GfqQhukRb0jdSU1P8SPFU/wXG+y8LaUi6/pyRA6Z1Tmhr
AOnyZt8iha1S6N1nDo+F5OkgrBvPR62AIaP11E56MX8uSbE1mFTLKNmYuIXi
hMrq0uuv29oUlbYgoxt0WKGmn5LoYvNGAiugdlDoBuRDDZk9GCbu4rFhEil9
ZAVtRJbtQ8kosbsTi++UMKdCWAZ/CxZvq+mMsZ8WCSYwM1CrkD51Mqr3e30j
v3GG4W8UyH684P0gCFga1TqFmo89pm09rm62wEx2Odw+r41nX24WOK/9AqAw
M+pwq2lhFOOEEaRORGXzxOEscA41YlZa1oAAk4/KJK/n/UDDEAr+63BYj11b
cBGL8M8Z5HsU2T7SKw0VHhHjJvNgNknqbT6DJsgPqz3rV51P/zTWAICIk+zB
H5zhSPkQLkwe1I/4X2Icta0g0SDDQgBupJ18EcR+RSHibqqNB+ZY9nLOI7fR
6ojpigB2v64DxEWUlWFKVhse2f/ttg656Cs0zHJWZhiMjqRgvLUjanWPtkSp
jgm153UYzvzziYcrmrMB7c/VQ9pQSF29S8STvXG9m9a2KyofBAu98F1toERb
Ih8O8QD96BVlRWFTeb5SedGEUWBGVJIKRSEI1T7AnweYdaa6pBqgoNHcu/LY
RHCPTnz4rFiDpeZ/FrnGo2yM8LJBJmePPOL8CDtMzvrsYOc42ybVoW8Yr1U5
1nW3zcojplDTt7IWjgcRSjhTPZhehexV/3nfwPD+U/q+jdmjNiTKFpugk3mI
iqnFQIOC+gHSJLE277jV7fgUsno4IFqZLUc2n/R/xcqCwOQcWR0t+JWSLttx
3z4HfQFqnmmHn8Fbvc4CA1sgsoIuc5MBaLhkk1lWTddRkwdnM7CGMZaxCrwx
CXmLcZbCBM5Ym/d4nPsAw3MXvirdUQEjnHq4RUBclNmEpHB0W1vrWcIf2Dlp
lTM/MxbE5bVU71XsnwcuLV1Pa5seY0sZ2sKSCoqusGIRqBrshLoxiNPRXIZP
H1jeskBiUerBXfOnnj79EEvtKuPdNqoBnX6DIQpf2GQpLpG/q0mRyi3Vhdmr
OvlktExRgdMtKSPn9G2kybZVqR9j4tYmDuhuiGb6I1MKwVLF7xVBIj/UndXt
OG510u1IxWMTelshLC4jC2VK2IKsB+Afn6TcmaMEOKPuzeJ6O7sfRH+qG9ix
6VP5gVaydxFHOpnTRzuDnI7vCThKH+BDa4PZIQxD7JFuvYw5iy+L2ffj56Pu
UzaO+emsgxY7+btNnUQM8CoWY5j5ZZmlaC3fAikjEFWFeQ4tdZ1cnlcHphBn
zERDm0TCZF3O+pg8MOmD7Y5jfG/KaL0i/rOcs8u+2pUDhf6RBvgaMxf0m+xj
Iuig4QbJxXelxApnINW9XYlkztMkDkQYXsqepQJ2WQvkAl/LafkWM1viX+mN
U2hk7ObpJZaSKdKUWXvPx2Nn9U8niMgF+0amI7pbgAGTthv2yMJZjcRk2zU3
NCB2qusgzAVrqQMmxtSoh+CI4MJgfYVcApv8dhhhQOdNNU+AZd2uYb4clk8L
oS4OxhpMpEXzovt4IjWFGboZxABbGtD6oqG669amsaEVzYpXXQpEsu8FEY8Q
4Ha7Chku9AzP0Lf9FmCSOkryfd7ZvIYKkq3YG9W24x3JyB6njfso5SmEmP6p
W6dElGi+ha9W0z0p4M+IOENA0802msoaTenQbepUIkVsly0VTi7wSoBfTpVG
49o8rV7f4B5V1YvKARzmmtjM4QM3Y3SXkwCkqOzMN57YKXmHSXLeAEEH8wPf
V3jvUFOppbJgXclbcterkUfE0x2+kde6HgvXinR2I/uWd339iFK/dTA471hE
+saFBm7Y/JNyHIjrUZ1tQPxEQvJqFHw8bMVCRJBUu5Hcol32XaW6rCuDAPwv
hY8ri3JCAvirPmukTg5jmmUc9IowaacZNUj14oRyk0JI4G0yF2MOkd9NlV59
adf69m1SM/nyCpkBSFw4YpnsRBeRiNkAy5wLKl/rD4x97skKyj+uBIBPz1Nj
4IaPYVVCRLqmE9VK01rFal1kpdLI3WCbtwsjZdKcsAH1d6jF/qNDYJvVy6M7
FJMWbnCIe6Q8KTEXoeeZpCI9ksiiXe5vXV9w9EUi/q9lUeNMgEnxuXSGqsOY
/tFKyNxUYsyMiqFCTCLhxDr0WDgBuLihiYNe9pDjpJTCmyII42zmd0oVsS+q
UTn/8y2VAu0zofQGarUciz/79MElMFhqP1LLWQ3Yywa+8wKtkAanTsFzIR8Y
8vs30GApn+QXJrm9cMKIC4PcwdKw8RrIbQSLlI9qASkprOyBKxO4hlPsiToa
0DWo+0jOo8R5GlMaM4WMHQkrix2t/yUTUKLxYSTB1pYIoPm2hcRplXrAdg8W
a1pM7vDHlv1hXUlFLR/tYCAuvuRPxEDT3KwTqIDIRa+xLNVZEa8XzFKfAHLX
LzG+J8ZkZMv0JY+hnCIBlwq+oocqxadoAEucALRMwJbsYT3lc7Y6e9e+VuED
feLF1Q/o/oBP4YLUgJOXM/zpV+3GdJpveu+wQzhXXyijmTB4jGIErvRE0OxC
WalbPES7FlND1CMIP00qCjP9l7jRMpD106ktVi95hZxYcdIyMYWZosmdYnGh
f22N5b9dBm0wM9SIb3R3XmWFXtNkHeYaDKXuRjqOv0ISZjj+6/gT0xuxXYdQ
vJEz19uowUk7NYcG/IUAr99OA+j08YytIA3Xc5h+h35hioo4wB7bqjuq55t7
k8DROp1Ba+RkVltaV6U9PCgrTgQxuybnG/6x4wz+Fiuoxwli6sMsoEg8/imd
QHpe21nh5bV4XCnNJoA3CguC6NTV5i/P4vyjFN6YYxKqVvZKOAnu+ISYYrJ/
fhuMTIyUMRwlqVVezm6No/vMIxQu68aQhDwb136bp75OenqP79nJP9iTOwg7
NeW0W253Imeb+qmwI4awECg/yIH7UXTwQyFeHkA/UYQabHQP6+bRQO4JFGvH
LcAr8aN+xN8I13FbDCvO9TRLOu4zpyi2gD4GXCFbykSyYIuanf7nijneGVMA
X5XvehF/WKOuL9cw8oBN7IAl0EaQhdI7qyZxechioRTctdfqoG2P8NJU0Ci7
ShJW0wWZPnJBFTw1pQrdFGjDUuD/KtF0kQU+Y0igTszcV0g7/SrmA4TJ3pJM
T3OBf3Nkfa3X/dLOVvuXCp/PtZdSUVB6lazm81+544GHu5RAOqosdWAGOYh/
JQxEaw49V3eQBlLTNqDK4aGRdJgnSzK82g66SCm+ICjhelM4XfwvhgdFdYG4
4KyBd7q8Ffzn1zU0Y+s8UbzrJxLEF2dGoOYpFwPiKBDEZqEWG0K+mtLr8Raz
FXT0/XFrvwQ9G/R0M72Cj6q3a/z6Ab3JMCHQFziUaKtsvauSW8sDPDBm+ymT
I+/wlVAjJPahB/nWYwiiGvzRbUM3hGZ0X9S5lz3ndWdQJAY9e+aPh9bT+dxR
KFuW1326Zp9CVETLUeSrGb1qeXQ3cMDkhcTiFb5HvWbe7V2lR2h8novTp4vx
pGHSDoOBshA9ALdGNqmzQsBHv5eRRpZfodZfgmm6sPdf9UB3mHM7tk7J+d+K
0r29r9lwJMToi539tDYtx+vgvLcJlC1gaV4kn8y44B8PJqDTQsVvnk0g3OmZ
C2fsW0GHCDry/46Skb+1KSk5EDMXU3/WajdWAN4GiD7BXUDMcEe5NiIku9x8
iwil4VZuopmer8BRBExuMbnw92SqyN4/GYT+gjzmaIwGQGIkhrWL8ng/wy+6
Ct4dU1uT+j18cj/io3XUr4O9XyVxpIu4xG8TmdLHf98e54WJ0UlK9vOMSFI6
XnBtaC6wdC9T1BHc3Wzcaq1Xz1NH4Uzri5VLFaG0RvyLF8/EPMZledRJjeEr
IqzxFWYDgcUUlrMII6zVc9gR4QjTAVtIEUXpVZWRqGz7JfWEvOEoVUBmfKVh
Mk+I3A7mfMUFogWYO7qRXMGSoI0kLdZtdstHklqBRXrBOtjUPDDwr8/0BH4h
O/+7xW7Zw7EezHY0FZAwkJ9VuHy6CPUtPsa8Si/4oQNQfXgdpbomqetknxEj
gc2L2/xKrwzPmePw/WInzI36yt2gbcXFawH+N0pNqtNVJX3l8f/re6XBdH1Q
283kodM5csQfDQmOgYaI53w9jkvFNfPQXPqZzfhkXd5mhmh1oEvhAwMmsHBD
4emHx5QXbZi1QCSF0i5QQzPyd4WFmzBn/7L53vkfs/SwTW7iAgrfM0P03jtu
5br+33I7IPzAJ2LWsvsLRSu3jCI5ukWp24cmpSDFZZDwbTeiUueergciUM9S
TWGgDpN1P53yc+Lj/4xoKVS7/RnhSOO4GiJICN4T1VWoER8C5LQyyaV4Qwg2
xZVnoGB/aKwsvzqeG46M6Ci9FUmavIMKLbmrRhNMCNUMSiGEH/wW9sJB7BEG
EDcEOCc2uijhSOOBOeUAKRPJ+7igCXfabBOR/sEbf+WQh4o3CHqd5URmHiVi
FBppPYHwBNvIa4iGARCOj3ZiKM7fNMu+z3s4iueLP7/sEMsClOqVn5aQ9X9J
ar+WtrbPAYOSicp2Cp7yEhLziyVaSFdEt56OFgPdq1GmTP+UgbuDf0U22Ask
oCiUwCFWjUYUnAR/GKvK7HD5OgvCSaJh+XkP01OBVZFnWF5xv4XSMStpPqe9
IlpJnvqe3W5kO7mENKyI8dij61uqrC1lHl6f7t53UC+Th6PrUn6IWCPgJP2w
8G+s7rD2h0e9eUwgnE+rq+XU0tJtiV4q1GFQIxxIp4/Qu6grlBZ/61MldxCw
aq00vmUBQIWpx/p4OdFWO1PVxk5guIspBso4NnUuXjPQZYaTeWfjjkeTNgvh
znGERa+bx9qwk0nSiXCramVTDZTe+zM56+MjsGpyjUDO6NTP9vCGFGfbFoCP
b/BqjoAw1f+KCs1Srjb4NKb9Z8FLAeJMmgjYDR2/fARWVe3EL065ckr3DTql
KAvpnwW9FdhOR2abEp4kmH11dUXuHaEHQbh9rGGoibwEONwBbD85IgjQqSRr
XijQ+zxOjYHxjXwOJQ+9yPfWS9HJH8+FNtynj6p0ORZd74D8GS3p7RNH8rRE
p9ENfgKeMuyaBTiV/kCWmxjv34Hpb9Wz43bbZHMIWZsi+930H3gNit0Fd/fw
12Ctjl1kU3BfrNUKb/kUxR6uXnwDyWlKu1xgIac4VvroRjvn2sHqZGZsD6rq
sjGfzRYNxONsTSc0DXd7cq79B1H6za72sj4ovIWNsGP4fVatpCMiexFqKYyd
OvKW2bpPWyPi8ee8GhDvEu8f+Iz1+31AnGCNAeQW2txxqsD8bo1OrJLt9CmK
rag3DPX8JJPjvUO1c0/qYhm9/rF7CItMBxj/jUpW3Hmtk5duE6dsiP+6TroW
XwMEvAmRukmCJqlqDcjR3L+jsb2UFtLkOFKE8wgS/zpnPeGHeYcnEg58VXWr
s77j3PAnzQ58xJTxW20uM6kTCdKaTv7CQxKnK0y9KSSagRVzoTMXWrraJCg3
EMCf7Lk2E4QuH9MBPHtiCFLlkyOVrrHZ9YnTL7sdE9h7wqyIRYkbkBR+gJss
4HANlEi4QDAXlW/FOjazO7thd42L84fva3swTeQK63heENnDh6d329AHNH4s
gB0+yupIZGznh5p1Tc06sLnF8ooGuaAOW4mEYWjC4KcAgW1ix6Run4TIhXHL
SW8FzRpD4BE+6wneY4hzi05X+xbNdcAKt6Vkq5YLl+Q2NQ9+lsge+pezOow5
JJ0RU4we1qMf3QIyTu9qyaAYwtCoUQs1U3lTxOTXpFKcFKO6CEwbRo1DOCPW
AneVWArP2jqLx37gxPbFyJgfH8cqEaLb/rFEKlVYqjdccSMlbXtzHo0F81YJ
1UQwE4eekUIMgReyz0YMhf6nGWFmrr5emiNXflDn3g45EoO8iZQ96Ji+1mS/
DaoWLhBvgkuBSLunwogeJYCYA7o4g3KcOoAIcACxK4kTn33fwcyfNLLO6yhZ
txQuaCuyuDSMvIDlSzguITCmz3cGmbOdgFfSzR6QvWvSQ5jKq5ACJtsQ9hSi
NQa45M3iSS1ElDoIfiggawSLnEoWsjlV8aFM7K6EpsGShr1x21HHP4iWSvn+
YCx68FzRqFHDNQWQfbN+tsFO78ArQZTqvoLZ589wq8mGQTX1VzVL+j/InCPY
cwvU3m/yLR5XnPJhKQsbtCFLw2UtKshlUpEAEUd9Ui6mTs5iSTe0UrCK+k/K
zzyaFoqHHJCEO7jpxdA/jdXZmYL5XtY/Ztbzl4k8J/kK41Uq1B7Rwt9bBoVe
gvrk2mA+6TQoy+dIaltcp9s+XssvmG5S98m228I2nhCqs3uWOERiUE/xnT5m
AwWrOBFgEis3dUyWMsI6581IAxS57fSDN+99KhQShay2zruzNFHIKqBfcOQH
08lW/KXEVdIGMhVUshJgDgaK+4sUQ6sByRJaVWC64RABP5lSvVsk298wSwQj
98PBwoNtps5iPbeqioPnxZAbHj5wYEC4wmRtZmpeiyGlTO0U+FPyJs7u3dX6
3Ld/ECXvq2kiSZ5PHgS9enMu+UurD3lCjyKa+g5K0j3MNudmEZt56PWvKeoW
983LF8DLV81rYhMBRGcKO1F6uqV3QsCku2hjCctJ0zgaAO7Mzs4aSttcTK1/
bPZHl7WsHkn+LvwpYeMydg59VbCjg+frB1QyFWsbKgU0S5ai4uf2GpnWQPnC
zSNRe0KGELPIRNeTYJ1k6kNBXK1wEkTcJEmIaIn6C3C9XNlnQHj768LsTahq
pY0SgjeS++8d+LUy9nyJFB5Z9mKd02noHfW7pEAcY40XthiI2AvRQiLFAKdL
JRzStgOUY2BcStlVRXqgEzhoXDl2cmuesjHWjzNjcxQ2EGcUQCazPBjNm7YF
6hsklG1fGI/HxgUTVRPeMv/qQ+ZVuYhBeo8DibNH2L9wVLXcAkcfRUwuYVFY
N8TAhWb5WKNR7jOQg2cxE6zgibNeHv/E51jwZn53ATnUioikWYylEsGz42+t
zJluDcRiWY2k706c4+4FIUEbQtwhHZQjeWfvrt1PQC8L743GOBlvlFY75kIr
7jUENH6x+jI/X/wLXbH4GV6GHiMvjYzm2U7xYk6JMxRIYeSZW8BzvnZFuFFK
fGJtCV5V7D6QUS7oAH4aYATBzQ/7tydXHLOyNzXQmUxKAJTZHlGWkHZMWEdh
u1n8kctUj8awdUbT1oMH/pp8pKrAnjVnktrtPJpjgJjYC1Eo8rBR05LEyr7I
oVoSdNSRnDPpcPWtWZUtOT0/Kr2+IwdV9jTqK05XIkpC3AV09oq3t2klJdYY
y52c9y5YT/UC1ATJHwdESm5QRu91nua601yraFOfCVJxJWAKEHrIEgL8lItY
91fCv3n2IPRvwqQmYIMQCM9/khRGFWyYKwvWDwIHVTF4ekRRkseunLlqvO7q
qRZlJDHqYuXN9Nav+wwGw1jTDyIs5YxvHRtm+JS/oF/Fqrl3D9/SLGMeUI31
iC6sgB0p40ZX/RqGFvgeLJLI6nsl/VJvNRNxHIOg4D7lG+PFK20xwYFsUhh+
YWZyKhLem5EE9HLQK0NqafFasvkceBtEdbFj4CAFLA2m8Tlhp0RBD9M/E9fy
bkihDg9lIZuncXyb7OO6jFmENWeXSoUqgT2nuiHgJQvxvN8QxZIBXj59VAsU
MOoLbK/5sBXW47Gt5UtFyo6Ol+tXAAIM/gGbniX9R75QmhsgsuEKeEix+Ick
Q4y7tVoghx1wi9EXV9CtOABjOx6zTrLZr+yDb3mpud+XphYiAzBIxyxEI8gr
SxIHH7HHaVm1x38fMWHHFqgsgJ9ISys4oV2dMk+bd6xzi03h2O/f522dBf2X
mYC/9DA+6vbV3VPHKlRmSZJrs2oWrRIwpIjqiFHGYlfiWFoR6odQt1tyV9Ib
lTfDalrj7TqEuNh4KHTO7CyRmE4irUJfrlcsOoUEOVnbuQIwrxUWwtRTecZ3
vKLA429jQ1VZKzQNi4m4svn02lH1LXYPfER9oiAAQM2Q7Agj0K9o6sjuCERo
BtHYJ9fUQUxoFFTnvjgVMbbG1dHL7cn003nrGcrFiC3OqOqDUoRVtrPVuTOp
A6n4Hr0T1/4ksfMr8JqLUb+rkA0PsKTT849DPmdRXtly0+10KoGAYSOTqTKS
XEusbO0sfDhnO1CoBK91XsOEkZr7occ1ACLrOSK7PzJ/Z4VkOxLwEOYV56yX
WvSfihk2uVD1QhEKA/FRnhBOvNjY1FrbLuawJkdrIidujlh0VM0Lg+ohoMMq
pboc4I5dXSWgmn2ENdtq2TJKfso+gElxSoWJ5E8qf6OvIlJwpdunFsBnDNTX
juLGqb21yXozre9coianKqPaaPLLARz4J60Vs30uTew4fjYdaKh8Pb7ZsO3c
j3nzMAMsjB3o5I3oxUV3brmqqspijjakxo3ftASLiu8wmf+YddMgOKV2M+UY
6SGrL9vS3ql10jJnSsq1WBpmR58wAt6XO8ZcpmN5DbJD3jIhfPGI0898Db4n
0Tu2wq/zSD/AufKwqJfSSkxrKF4vOHnrW7cySbBWp10VrhvkXALtTebhS6Sw
4iWf0zhTRy8ky5m3OfXpB4tGHEL7XYajdTMwuOXVqFsfQv3zX002zvxD2knZ
T7GPjDEITJcHpioh8z6LaRMM2plDTEq0NxqfOQpythpXe241SEvPhX8fZ17o
4OEYLk7ubAJjGwc8EITeSOjYgpCkJasVd9dVetBMEet2JnBULqYCDn0pRpQD
sWKzfNt9PTbWtd3E9sOSewngUMm1SoxqKsXNLSQPa1CmQMeR7MFT1PFM61rH
/82L0NJzTkHFcSj3bZBdNEBCt40mrTriLdMBvFknhg1/383FQlDnnoWmU1nE
jwJBtIPa9GI7so6Q7KhsygfJMbTpxgNWx0P1yZEhtJR73XqsJBjtqXV6W33K
UsgZLd2lmXHRcX/FisfO+/xZ/5ffCY0iUNx49Vu1h+lhYF7sI1nXO+UFQ19P
3fSF/u8lsy8WhGblKBOtBAomdJlHGWyeWwu/VZQwv6QeIjLOJN7X89JXnjxy
zY/Y+AXiPZj4H6gk/QG74T4+ZH7yfmVCtQUaKkPsaCAwmX+zo2A5CpV8d+Ux
01Q9LYp5ebfkslgOYHX+kZX8tXT177r4KMFLC0X7im3A1iXwT3z4qz11FIFg
y+TF1+KPKRZ10LMalieGU3IKB+Nh9auCboAZp4FNrAXcp2m4pwUzSHihSN7C
4VibXRJ7y2vGQB4NsKI0BF2rg2qgvo/KQYHDcZcubxiXJkau0umcr/gmn9hS
L9uO7X6nGb6GD+e7X75Vh5wVbAXdbd+KPo7j+MZM1HG+upzZdArTneu9gdFM
EUurWqDFYAS7Y/twEHdwUYoygZj9bC3qKJR81yGBbyZl1tYPut7IStPHcx1a
DQ9H8qTXRFhl43TOlWpWMplNLOkurPLAAny0Xsml5Jl1rB50TFqWS0tU2+I5
KKS/gFhuxazjm0JxIT7onrtcupcRQHWMwfggwmEkPQ+dKlbxEtfmMnfcWZxE
kPcWM6zZ1AQw2AKgfKiXkRONd/HkiCQ6V+ywaqFSEc3YOVkys2VMMfA0geeR
ydeC7bxX/R6CBtFOwWbbHzKr/bpnbX76PGFAclDIB7BYaadHIr+1yzosbp6j
US20mOBT+PYefEFpJXZ6GLyWQfQaE8mQdAdD/42vJhvfCi3eVr1DgVrkxbuW
0fT+FHNeumXJ1rBqJhupAIBJFynH8j1hEaWstiHVC3PEXVfP+AFRNLhlqgHu
k5tmdl7ep9sO17/6JdbfR2Es5BowNJr/a1ptwAyS4F0GU8ggynmUFb5Qv9Bk
imyFcRyhydXrJ87EcI+TD0sU388ZsN6oR162SLupKvlnGCqoBs/zSW7Tr7NM
tLznqCM2ees1/NH2+5nlQ5qHiidzz82yh2WOxZ69BKzdcyqZ0TxH9qdrmatO
FtOxVTBKydQMuFDyF+E/w23CpkyA2L8pa0FRnlciWvJHa8+Ykad34aTMlnn5
CldrnBJzy2Y6GA6vH20NHobkhEVLbvIpaMurNM7U7ZaWJ+E3OpZMyFKGulRx
XhLSY1z71WR0KpxlXwi52GqwI3PQ9tjTXxnExnX4Suwahpz2cS5SEuSkkO90
OKCIpW5x90v7so2weZu25E90mVgBxqnFZzFIszwM32DyXc1UblYYXnANA37e
UqdBpxvDA1HBByWViBEYV2gsqvt8YkcbpjDtZd2O2nfgE84Uz/VqPXHEfF0i
AeuVcN4XfX+G2EjQzSgs3bxFXCXknD0koiVUh+DUeEx8T/vvedM+Jx1s8Upy
yKmBdFroaGQ6IepS0Y6+asARCwcDBej7xH9eMJTO1fsqUTUiLc5NL5xisunO
RQFu0x1+daffpi+jzCRuPx5zSmKG/AnxZWt57lgoHVQA9uCQuL+9yMn30FfR
D/6XmqSXO9KFP+IT5YcBbf/7CaHcbhu7x6HIz+pUedgu0Bdzh0gpKjlGYroO
49mm9u5C19HPI4RDfzp/lb4BAlJNjYLLbfFO0N4QZBuf3IFjhYFK+Z0ULnpn
DdWx7seHGdIQ49FUv0Yh/G+lo6cBRHgyQzj2AQZar12Tn+q2GKsrxiq3X8Cz
dHJKNIBOkMV0Q8yjQJK4mETHvLM4j0W4caVCsPzET1dMyYo6V/DQdjr99Ft2
8cdkHElRJpjGUplOL3EVyHE/g63qvDm0ApSvAzO12r2h6ZHaVC7yin9arCAd
1tNMBZ0fpLDyxcMv5HrfXNRhLnFEm2tQkZQfFQbPD4QxNiOOHaBik8cX2PHu
bL3xjtsMjRT3XCXru4yEB8/EnEIB6/lmV45lvxUX5qEw4PAAzl7WZ86lS3vd
l7KVD7gXNux1h+umk3iR3Glk0HzamH5oxvcr4E7rZ/VRk3WN7G4L6A/ZnLLZ
7wZl2Gz0hPGejuA1I9TbyvcfyKG23F8HcUDH2N3ADQYSBtV0rUe02hEGoU3S
mbfmZ1at6lgb4GV9h+dVW/Gz6wQXg4DZeloNg/bbR21x7fezRwQlRgLc6Wn5
07wSFpE11hPWiMP0CmvtPJhF10FyizrV6Ek7+o033XV6YQVK100fdVx2t4VM
NCLHx/KGz8jPjsfk6Sfo/LO8HWRb6I7HPQHILD3nzurIGER/TrFoZaG1VkU7
IrCifzh+GCVqXMTExAMseokILTrBWUbOVE+WBV5u8PMuD8IbSvwiBIjKz7wK
QSPfSAQzd6J1mEIW4328BekIPqEdPZJCuXPlk4MaKsI39xG989lYqN6UF0Ne
uj3br8C6ipWx6Mpr7tJyPlPHQsa3ynIQD/d7LOUQrfAIS/s5lI0CX/neJI82
ZkabWOEHZxeu1mroH0aeRtcBHGGYPPafrZoz0KgZUS2xBpRD2mJVCROcXxej
f87rlTiyU/ExIuvECzu/mNJoXXYL8LhjXbB5FUzpmmmT5nSdQ45tw1vuAHQT
CSqNzr+kul0fDh4TyNC65aCRazUnCAX7RPgUUfv2VyrcygIiGA7tb+d0sefr
9Gzr/LsiEB8ZwsD574hym/smYSVail7GTPhqTJtGtHZCJFif1IipPUoNhxqR
NzRl9EHmCmuOh41/xOjGM3mH88zc+HCqeZ1SlUCo1hNzY717DmOpKHK13D7l
TvHExjAChJlOW3JgGxsOKk5RR0PVjBp7kbjTIIgim+i6noQ8DgRyAtuwroHb
H/l9+bNU0VpkmANJNX5hnaCU2A8Y96d4pAY5VLNHpsT4kRomtP8pyQvKNncm
/RmzhmHgkMBxCjTlNjNO8zkoFylOLQBmz20stxYcpPqoDG62d1FhUD2uM4Zf
Ii3uE4vBiY0wuVjYKjzLePvHy1devubuKu37CIJeJOwp6uiSSSZ6NWCB6y8U
z94Ejg9I5F5aWW2IUHmyXtCr05iZO0Lu4jMImYT7SG9n+0oIx291yiZzyAcc
QpTNPCz+OUnC+UhFC17djbMsRjsSaaiRDrr8Zaz4Y1LsdcTWdpfO27Ls3zYE
DW0nNrWBvHKsRKSGnj7SUnNin9Mf0NoH+Fofv9WycM65mNqVqTKHlRLXV17N
JTiEQ65QFK5AyC9Gn7B6655mCQYP/l6nl9/k3YDZuVWqsnjZlgDF8NKHs/f8
UDC+aOK8g8clTrBVuuur1RvA5jzunZoPWIM8obQP7RO3kbOWTiy/nOiWfq8G
3GE12dIDS9jWisazISWWM/VA4x3qzJIrgnuAn9Ws7fybHL4/1D299PBEfKW5
dytr3zuvhY9de8Pc/Owj/iti+I8N2XGZ1Nc8AIeUQQB8bZNqVq2uWa8FhzFj
FNIxRCZIzG6tB6VZ9HqVy5hXK4QuTOZBSJK8EOX3nhUqP/BBKTUp2Dyr5NxP
R3eU0oYzp4HOqK9DYS400IexcLGo/bpTe3HtDa1U74jbM1PnTSh7WE/Ew+0L
/gYAJ9n7bYXWhmWMyzkYRRZ09F1d/PqtQL4uVzX7AwPuzfilGoJKixnVniOb
awdxsw7EubYHt83CkGacCgSbmw2zqgjmie+C98Ly+EwFYZDqVKf7aIl3YFrL
fvOqOiXRdwnZI6R+ITiF94qhlQRco9BJMUOOOsi8wuxjstbK+ZiC8HaDozvp
WNqPgm5TJtiESMlQ4cjMNMXJGDM8+Yi6i5Hgmi05bKCAtiWEk9CbBCw/iweB
BkRXmqG3RxDIT7wWBaJmiHoGl5edJmaORV4r6xqf5xM4XLY2C/yaZqb/mFxi
W8pqeRH5CkRsojdgy/8PqJR0nhhEHyjm0masEBuEgNVmFbXJpVu0ii6xYESd
z1J+7zfFbOGIMVmRLjoUgfSrzbL7c8H+OEw/aSqOJHeLFNR3K71vYnU6fR19
Dk54r+SjfkN49Ew+NDnwtLjzpoEgl7BF1QpGGlRl0kLrSjoxoiVrDwIuHcY8
uR+nXQ/7ngD3gveK1atSxZ+If/UF1WXCjNiIyk8+50VoaUd9XhEfq+9Dp8uP
tfAXfcq/9OE3wUDpHXHNEgBmQcXY8TYw+1MfK0MmG4YirPtTo8FHxaDzT95a
g2i2XazDv01l6eZw98D4ROuuf9CrRqbT029kfzQrvBDWzZ4Mr/GpvmcJUKaI
lQYcVWG4X4+ewr57ji/QYYiLVvzNKOKyuoGK+IV5bBYjuhXaPlr7HICgxg31
8soHVYo60tFY391PgyNQOP4yw4DPeyB2F8ySniMPsasOjBJkN+NEcxPvL2Jx
zBU3/vIQ0APVt9ADcU4yI0qTs+nY2QWchsIje3XsYMi29o1y53KILMhXy4EO
LDFAZidPjQ9+1kLhrz1YI5CRYD3oHrNs8RZlfTKHuX5QKeJfLgalQ5UMd9aw
FD2gnW66a45gI38CGt52KcMYDdFIE234wpsgHaqJs7mBd7nFlXVir4vT+IQ4
xtVQn/gZeyCzZ+tZEEtI0dnYRNq7bOGFR4jRkt7bCf563MutV8gSD1s+hLlT
YdI6eEqD+uR4sE+XFAQfnAn82J3q7Uhnh9eKO8yOrvB6CGCK/AUT/tz7AnLr
a7W5w8TZiZUkFu9LhwOJ7+aLQPXwd8elpAxdpw6OV2EXLvFR3uz6ZsS63/zj
mmE3M8nMcd5vBiwuc91GzTUxxYx1sYVYU/LzsCCcfOeV787mlAiwJW+MhVG/
k53m6IhSW6fe5fup/EFU3iA2SdH+UHJzpjxjKp1G0DTK82tZ3TaOXOV+A7IE
/lzXaCHvPCYmCOpxphWiUjI4muQzjt5ZY1e+Bt1q4C+aUnQwJGB4Vhjgzsxe
LskH0Sw51q4JEhlpXTbaAWkLCXJsHkNb6HoyD5vawZb0yL6HftQbQAC8lmzQ
UiE59fOPt4xW6bvTE5fmhk+GLak3W7EzKzJe81VQRuSZdC9KgdcF5o56PJpr
QJk3H2dAqeFw6hqf0CJ+8KY5J4vJ8wJ7CrnBcmXFKgP9ar6d3g4os/GzzpPS
Mu/Wfl/7ya/aCy23cuZ2ViHZpg0aSaPRlxBpZaLOHFNyVsuizWkbYMtH0G53
TVcjFL5n/BY983jZ0XrunYzqrRasKnX11WQduR1ApoMRoKitizC39z1Rheme
jg2iqxNjArsLLpJWwMGvRaKsBI3LMHTwqW8CJ6qOG12EPT0b9tr+WCmv56vA
Fk79OmK8zuO/grpEbPLh8BWuyPaUPIp7LEgt+I8J2jqjVIW/MfrS6X/IybnY
g9CTJ7hLuFajkYzO0whbOBCB+b94ewsk/TDsQouvxoHNbfS7fa1w95FeAcU0
olaUdROzaOObCh6VSWlBGvbJr49ndqZD4GoelCK372/dSVtayCIM/p29Xujg
FTXz9SuhYvZhx5lIKuFH74nOvIGCdNpbGWZ0vWZM2iMPxVwAKIDxGOH2ckrh
39C4TE7q+wwnXgYVOeiXGCTicR4bViWpsjVuAgvJH9jj7KOLvfthewhyBk/a
C1rlUTIcNVWp4pDhzVlfJ6SCNAqRAwWO2Tt/YvgjmQwouT+j0ifgqJiMV525
V72O4Fz6dsUF1vaQ8MguGI3FJYu6vnu6gEb3fs+ZVEne0tOq8URaFAU5fAiB
bfOzJkLVos18AHF9Vw4HSdH2KTI3zo1SJesp8Qg8Mq2XsRd682qeqRjr7Q4/
m3l5ApxiJjKY6ojGzKfzFkC0CDwEO5/qgFPr+2kpdg3P5rDgsdr/V44m6wmi
8I/4VBQJKkQKKEH//tkcm3qBSlLmSzSedSA04/hXTnkXCaU25dwaQ0bSfSx4
XPnBPWePco3kfenkvqYjPwUWAhEl8W0WP6dTXQ7SEm2FNTcq9wxQbp5+78w/
/kJu1vsLxRoUPBtDsB94xmhjzjpyo9E7iiceelhtX3NNLT7OSS+Jt6I8JoUr
7SAHeP0eD3FojB79CVJ2NEBSaX8/Yl401v6X8QHh1nksQdhwHTaa4J2flISY
5mGhAHz9CPF7DUiqB9gvREu08BWzb+14Lh9nG4g0daMG2Ge8ecrGJ715OPyL
mnrcyAHMRhE5s4XHZ2TYgf1Onz2RFKpzrSjZIlF3NuJ2agDg8e2X/OHxDtJA
7GT7WlUTeUvAMHYSZq4oCJM0Qxb+ELBZKsF04W0FjFoEtzB6g8MBKiZ8pUmu
xuSkMCdKH9N0PigmYhynfKHL40Kk+tww6DuEgZ6aSb5zX+7E3jyXyFpVgIqp
AM6WZU197uMDYH95lm8Ca6K0lLaZi+Qbrz8ZgjF1GvoK89G8HhN5r0kIJErO
18Dv7GPiaSz5LUPXSo81sx4qa0E4aB9yqqCkzymMyHrjlIJ+WCpcw+P0SXAh
kPwmoqtOR1s2oD5PFQyY4spYfLynBOiHnrXSD/rQlbyiEUxztmeadHpAbQyl
3raLFFT5jVGmbS/+y32ZxNk4uozfLghFoyZfsm5suHnDhmLcFf/O+7e/RfyU
L8GLwdwIJmRSYEolbkW4UCjxkDPO0eDIVlzzW/iYee2EZ+niiyENJHv6vEkw
1chb1OQvYj8btZdv8pbo16G2Bokx9TAIzt6btak0aFsAHYf0jCpK4mhct31I
YAt/j0zliBb067fvKrjFacutuoUYOzpr4iyF4UcKrzULd5H19TAfTZFLlFCW
a3uBkszqu/CGkWlLsP6IdZosoSD1wx1/BLcxty2jjav8pSk3cvbyBD0/kgIs
3XXvSVb2kxi0VWc+t6AXPbFIn2+kYWugCgmsmnsLE5hrc9Yy4ZWhHirTt13o
G8Tb1Y9cKmjC8rBDfHhn1D7GtFFzSxtTQ+svdB9JhTVhEPLoRLNvQMnHrUvP
EhUouEpNP6x8RZoFHuOKf1Fui6D8aObRekuq9JEzZZxwNCwUgVULdj0R253K
+yxveCJ1LxHSAuj2Zum8OG+F4TF7773lXfy9LZA263UjfRaqUbkxcH9MaBNS
KNQv7BKCg5DRMMCRcGDzsXsyltvXt2LTtIOqiVL6km0awzXSA54/3RirDp7W
I15jPkV8wiFAAkmd4P9E6JeNdHKWgE1g84U+24Zcf+rWM11hbzfxOVaSrmkt
1bCJhUbqmPQRG8u0qlR5u2+/Yc5YA0Siqp5D7r6mrB7b59atOPoE9aDIjyrV
elaS76OCo+t89R1Dm+PIsT/+6gV05/5sW8tBOJEyO8JY3GeBGLu6++Bkg2TI
b/+wHqTPHyGdomZ38VPRVp/TRgwywuXEPIFShvnKgsw9f26QLGOV43ZUbWYK
8cEg023c4AEjLtLfw0vrt+e5uf4s7so+gcZd9iTsP2+RBhoSQJ231hg1QS0t
evODzvGaWYHRZGg+/7c40QFHl+kn/CMwMGNPsSelGJ5eVj+Qw2m+Ep5CtZ0u
mmbhQKEHBn9vRfe9QVDXuX2RZeE0RjUGF9ORBm16DKQVceI8t8SYP6uY3nqG
vN3P6MvpeLFk//6cXngpz+CPBooWxuK/oZBjcn3wY3z0XkSTGKeId1iufkHt
9B5eKHYE3X4iqXwbRusqMXslEWDtskoi3ld19PQcxAt3+zkqmnpo5dFI97YH
DZpfLwmbO+A5ktmnvAV7N32z4JgO5+YLcfI6E2dMirhwCzRkGnerV4b8kzuP
vMWFvS0WiF6GtIlOyfiGd9l88QgiqCcE95eiz6Scdm3W5WgfcArpzjJgq9N9
Eh0maYejF1oO7zjVhzeWsSFyPJIeDhi5jDw/fUDj7wHBHIhi1jjiZl45kPf9
ziA88cxStlCI/NvaR39SqG3nYwz28UQ37qxloMgcVX3+O9NmilhHlSZqf3gu
JVXcituLgr+Hergog3096A327WmzE+z7LogKbZDuU/0WyxNUAorO2AjsZlMu
Krmrzu5TLlJ+RfRDh0CmMd7Y0M0TjI1OoHvXm4mFD2Jd5KCMaHekM9QuNhBa
7WT9DSTadRWTzB6Yi6dpTSlu6vPoG2t+6/7wSLg4hN0397WTBw4Fh1eqzlsk
jvptlxQFjqakM7MqS7X8L9MhzYQhXC4oKrdBhI3UjDdtPxw88RjOE4B4MBYC
bNAPez+ktquo5qxHX+VemWpxFsT+pU4tsvkK4FBBXMi/UA3UrN4F71RYeX4V
cewCsIuOQeewLJ4jHM+58sVSZw4PvW98Zo+K6q3LRmd2Gbd+sffr5xoiuFGH
O7gWc10MsR4eaWQjwJ5vMIgmu2NAoqqRP3jXa5Gxs9RV8L2wESvlmlFYz2bf
vKpG6qxvf+z3GqlPhR/JR/4WX8yZryJrIBjmPsWU/BGLVZ5LDqIv4gEp1MZX
0aIkoCjkzDFHAtHTFdtEV074DYg3KrE0+V5knDfkhiae5EyCO2xqLftjztk4
o2rzPXlRwlycpsK3j77nD0uVi/7T4E/hRmC8oJL08oGskXaS/sBYN1QNm0q6
k/GjELAAtRLAfW8k0VDYxoRsHEQXHb12eWEU/isy+QgxxBLTrz0LzaBcTw5/
5gT59MAqMvcDU++Q/VwUcSyUG9Tck2C7qyFMfPHIEfAeCB8SiIuCqP6yKuGB
YklEFr6JFa4IEgp3hPxYlqQ5ocOrAE555+tvTk9FGg3ih25OSsuyUGFqUmTu
eLxn5rGDsZcgq2ipJo9TWnjs4ktQsbS+YBT8Z9KN7a6Ms11T4Tfb/njFs1Xc
Fl99awva2zO89vMOZGMJjTeNKMrmvf/G79YAPquxOGZMNXQ/yA81FfugyoDt
HIbPKeP7rmEbhMtTXSy7UTFJLP5i6ja+nnav3SkcuTjotiSl7yY/HGJv9i3/
GhqlQ879WPO3wC2mb8FrZta3ftO9TkMS/zvhfZAXzEUQXozoEfg3zlM3ZeGu
JVKiWpYNST4298lxXtZzximcAFN2vT63Eg+CMFttXHDHQIl09DU/VBOlQslr
zL4YZftfa6+8ssFZcUv2/bJPPO5uVfk73tmItaUszavV2J0zC94RJK3lcdmN
LMoDxpxvMCeL5RmGxEsTHss8Ahvt12SM/O279xu/3ctQi2qXHA4Pi0yx4973
o5ycdoWkHbsTXVwuFsDbGLmX5l70LICgfCYgCJr6p/qwCeYRog9bm2D3BTn1
15BcUb664/ebbAatwt2WY78Ib90RdwwRyOOVQZm2D6zL89MW0X27RLd/xrTo
/gcUfF8YoU+61zrwNAPT+gjH6JNgM0bNxoLSvKky7upOXnBi0y1z5YtUQ9io
/+ppXFdPIZhT6rgyuEWF6Nv4FaN79PbRuyq8b78dzFBVDxdNvdsHe3sQqe19
J4iAxRk1cka26UCp8RE2Ao8GcR6KLvjzZOKKI7OU44Z77A8yjsXvVGCduWgC
/U4IjYWEV8+2+gMmTGbynCohw0TpqZEIPXsfqfhnfOySoap1ecgAY9WKKS0z
waVoyFS58O6JNkkJEeQCbFbClVXeuDCSbHlhyoXGuT2bQsSg2P7Qzdf29hpr
65ZDqDFvR34sayWEW2uNy5j2WfWorC0jsYAvpx2OPS17Exm6ZmFjJ71EQcvk
VtCzBHymo8UYRrmW/OEERUqicmJOYMmT+SYmg4yX3HvH4d4e/7BzBbIQHLsw
ixtlToFLwZalcLVivFLsn9l8QwD79vmr8l60CKS7tgK8Ny6s3J+x0fe4Fe3E
uDOSijcpj/W7xgmxoT7V7kp80RtWzfJRp49cNmuRMuou9TLfEVD0EvHlSIgj
IzhZWVQnrfup6cUoEyTqqxwW8YhGshZLFzsjdRS2F/UL/L0YgZOxHMHCKHrp
+Z2CUaKdfisPAb1wUMuVfhAJHH6wuwSjKvxnBxwnvS8wmd12utosiiyQcydN
4I60ukuqNrgdllYGbx2DPGXVcn8Y+chDP6DsMIxTkwT9YYawPrlLMlJTklEc
IqEhDRm03fAxxrQuUeGCQZlvhbsqtfeZ2P4O0QRqfDfKCnTR6fAFp0wf/vhU
M57/gXfm8U3jCMuUbZzbLRqMCwW4wtl3uMxemI/0oeHAE4OTbQSB5tbMv2mj
Nm2Iozn6Wvjrywoeng1NVWQc1zMp+jddOaMoRbnZEm4e85V739jW/4CBTgHe
Rx0jfSXR9CKp5LQJnxr16qNlKoRTya1CNquZEMtOdjwvFwBTVWb1GhqQcRw6
qEDvUKqznBKo9JzPvDdxGhnaoN8uzhZqVb0QOmXto1QglmGeemVFEAJdWoaI
WFUwHLx5aBI1z+wjOTOe8czq8vdV0k5cwbBGCruRrkb5ZAToXO16RhJxzAX9
lsyUa2FFIrnKs4fVeM9fwfB+My9jTIhtyh/Tdf3P5K6L7ctISAcWmbmuR0Z8
u2WdNez8VSCWvcwaHYWFcaFfOVUsfZhRVwKhcDk4n5Y/wHDIv3eocoq2S69o
f3OelGPXcjs8SiLmyKyJgZLFY1F91oVacjFsGIzcX0T4b6NwUUn+CuCnaJ++
39892YBNJOkl9GZuuV9Dak/2iKKJbozo4V89QbqhvvWFET1Qe83ZwhwxEVr+
1xmB8+5C2WmmXGYjTQh/jBZUx66W++pQCbadDOswAU/VRGQzAIEribmGHLON
1Zs1lW4dyIYSWAIORH/u+bqCxON18gNwGFpfG/bxMqXTPDIfry9TeznStwCl
l02IdUCiAMyZ2GrOW9etvertlWS691XAVuyqVIEYBdFRVMg2zpBPHV0Et0oy
eeNZRWY6YcjtKdZNXteoGZeOacgwDULq7I89mMy7yP4AfhbBiJKiwNwuY9LR
jwTIURNU4q1ictr2rplfqf/Ujje/j3//8W8n5B0Ru5Hk8d+gsU4rbeKLrQ9J
/GTwfUZpeIfeVYha3l9UGT/TzjDIz/34ehefoqcx6KwWhjqE5IX24toAlIca
s74D7loo4n/9tyX+Roal3WlZEuO6ryAZMgN2kwXOnqCI+IjGZ9nsnt/CYhnG
APideEcSDJ8XLvXGCUM2Jgu6uqSsWZHLB2QXvazFDv12Hx0+2OoVJ9WhStk/
I4lq8d0ntsrLgN03vifrbizIO5zL7kYbTmSodu9de/tpgjyljr6C4wR6BMWr
3jY9fOpsGZvZBqevLqRPevW93hHdO5eq2Zc817Vn+Gww2p/LTupvEjLy4Ow0
O7ZiNy34L2rPk84ONfgvZAmeH1hzUjfBc2QgComxfjAWEvDD3jVlhT305Maa
4NFDk5nZBviYPblI4xjOErvb09ROMfuixiR3dyliOJQJlqQ2M89HfVk29Jrs
Y5xxkZz/RcjiGX/6AesvFNkO8g/RVifPCqRj+gk4Rdts45WTgUX84wHgPqqZ
5ygGZdwUMXVmbDKJTNgy0o256abgnED4W9x5bB+zm/joHjNJxJDs1IIMc8kl
hcprlG8X2jBNoemSyNhsZorv3+KXaDTcLW7O2qOoMmdH6Vr9RP8mpG/m980Z
HxYWGMiIBHDs7uwzrZzaLzzRaYo8WPVt2bi1r/uykdKEN5RjBZS77kW2F//U
wTbwYHQ26zc6Jsgm5aEYI8VMH0JSxPitvv8eDGgrBsaOHLJ2P+LjSZLBT/xa
5lTKIw6MeHiP4Ma1k+ELV0NnNu1ZyZHEitLuOwG/XGYcO/G/6tIAwllAsbXV
06vW8HyDHwohTkAQn76eEJ1VJ/Ffp/mbpWYhz2pIYuAV0JAF7eZwhXKrXS9f
NhPZtIBDu4dJ4F8wM2qqSGFJ+RfjgGmi1z0VTQ9y8yiYB45CzVp1rFPg6Ynw
CDhjpM3+61I8w39QnXAYyQjJmXx9jSIXLwVSeYl7tlF7XaM1Qs+G45+H8n65
HFpYDXEpFodHV9vl9vd3i0GF3vlXrCTLxT6/ZLCKU8Nk5zuH+PjWh4NdW0SA
J24iZYppk2pZFoN/NY2BUXjNjpjC0D/F3UVHR4EkOg0LnxvpIecMrHW8Iime
A8vwkrkDygCgkG5Pi/GtPOj0IR7xgAOw62AzJWLYo+lxL/b8pjkXihDg83pY
sysToekIk/sJg9AjlaKA23jciinF1WaG3jUFwGtnr9SzUVQQ67Tdh5pVOrlr
/bMaQa2T3VBq0zDQZyOAGcPQlLEYDpz1BGZRmg3x0D7ytmzM5yWPncYNarNm
o8+z5C1Q3muQwhIu2ugr8wrg98SrprX9ePPI7KReXQnw/HBtAkV9KXZivfTF
VqU+1qvfJrNNE0F3As5x7EXnszfU9YnlVNdFg/I/Wpi7X2wjIbcDMII3woFJ
yvMNwHFXxbi4XbKf1qYmXwM5AWiWsTYU838SG7hZFtLPzl76l20fJ5kHp9EE
FwJ9jQSMmgzOUnpY5lhC55YUzIETVWEPEgLP//jI0ntfYYBERovcokczbbvQ
MtFTKfVUxLvrNzXc1Qkpe0CjvkEX9Mxsn4ZFWTFTIS5IXYwgd5ToOeFBTf78
E33Dlv5UU8quX+NpvQEUUCP+TdDeRgb4fqr0WeGkqM1sKzABdvJ21+pyTYhg
6B6xXmlpQy7ZOsQeqEj8s6Lr+j3e2XvYXs1ftod1ZYE/V6GoNNO11QxxExzM
jTTWHpQAKQKeWoF7tLZ31w5N5277CRPrWJTNf20yGo+XsuN8JyKZIJ4H6p6Z
3gXsMyGfTXjb2k5H+r3Fsdzs8qhXTPy+esMNRHMtIYW6iUZq3jWM/mURjgyV
/H5T46HL9I8rgICZbKh674t0Ps7IWhi/EswdSyFayfwAaxaDScAJp4H7mdvi
tA1Dx+8jZCeVOk7k1Yp9vDKjvAm+QK2M0P2HPwq3/DMOlUVb1WxjrYwaLguX
S3/8MZNEYZTsIJwXSU2yud/q0O3SF0BPzyqd5xZt1Fa/sWmR+FvOzdHx2Lzj
SVz70ZjJpIP7K2lZoH5GqC6q4Mg93USJTNPqoNO0HDWlwDsiSMmuiJhqrWlf
UR4vvp/7uKh0C7y0Jvi1TE6FkbTbnPoi9CaNGXjwLjY+r00a8d37SAs9D00k
P/poeXzfSswZIjFCjpCHzfmzsBjsDvcjOUoMa1xgShvhkgODPK/cUnUu2xRD
IyPBa6GcctSN1UUQ1nPAi8BAcRp14ruo5KxppGZt4PMIrfbqvdUWgLL20Vdv
5fwrGEsaSbHWf0vM0SwCJyVp/+uRPoRrQvVyy3Q7H/yiPykrhsycHlJlnLaH
ATg+tMOR6beDGwU39idc6DslfOsyZc/tsFweTvAWtBfEj/B+LyGVkic4AgPM
b+0wcs7Dc6OgXMg29ZKO7KKz7nkD1S5A/E36yPPh51QPI3gGtbV4itrf+ck6
bVEf4F0hFF9m+Ce2QJbPWmxF6Ta0P/J/6YaBy/3O+EXyUOesXwnsdhu0Nxg8
IHVgP6EoT2Qm/ap8DT4NSX9n6hfNwj+gab+J/iCjCbbNJkFR1/cU1lxCaHEb
yLbhmlA7SACiK2a1Aukksvl3H6hXTubg+rjmQ5CAv+6UiI1SkO0tH+uQOysH
StG31v6ixUuFYcIyraDaFhrbCi949mxDPiY0YSxEWYi+v52oKM7IKrMeAU1B
oOnW6Yv2s4hwYcWKs5IEDwgfQ32W6Pset8UsJX5hZPK9tuPtHF+e2lS98kUU
10RdWOidArKBLu5iZfKqk8TRda6/1wKNxGl2/1vu+iS6Dzi4V11Y2xJZX3uE
BV9owuHPXl+0+fcmKZSJF7r0N4Dr4GdcB/0Fcn/qyzLWuisrv2Pbs8YkOicH
D3LZZf+vE5N5wUvIwGiA/gZzBg/GTYLAlBYWRGq8RPSrnk71RauEu5Vh89OL
d6FP5yrWpScGCN8dESfuufalTx++IpGp4zgaXJa3sm1pdEoMl4P3hVo9CYBE
iGmJl5Ycg0JFiTtZHU1w1oF9lM6I0F70m5dKScIvItJCrG2+qnY6bzTLcvK9
C6PuD9agQ3kqIWqPkCouUsQiR05qg2ltMN6wD1ji1ahRuH549Mvxt4apx0Ke
4yTAXxJPY+xjehsEEqgOnb+96svSJsUf/ZQTAeGrinDVIAhf2wDDz1aBDBh1
MMPTC0uiQzCdi7AI9kz/Tld98TarSO2TgYAy6OH/gQtjWRr+PhcRdzoG+V/f
R7XizQQ2ipC4WPMCUTUXLEsjLXa8Ek0OVhcUPp07Q1UExvfI/AQsaatNwE52
W9mgsnIhxHJuszlTqa98cknlpPhEbG+ZyHPL7mlL3iKq9TcPI70P6/eREwyC
W5VWqcfTwiEn4cPT0c0eYUM090jl+oBXNQyvHgIIr0ZgxNEKlkgXb+2yOPtr
k0zuaLP8hJCL8igUo897LopYmSlski1tSfPDiYRk3huELR0ojEYVaeWX2+3Q
3pohztRahzThNZ7ZPM1mqtr9OTwkOJPYUL0NNzEDA46/pDvgGWzl/v+jk/JF
sS7EBeQfDPjd11F1qSGIFtnkB6zkagdJTCoIlv0RAjVC64DXRfTpn+o5Qwky
d02gGpLVqAmgwS99I17ZdmUdj0I0z5YuCme938w62jZmYFMnO/MLZKGJFh1l
Hx2VP+HTL/l4M4bfzxkxmmWLFUnikPDEE2EUPUbl7TRmmueS5Daf/XX/mdli
gHhkJsFoR135dNbC/M4zLo4D0BusKl2Ci+jAczkxqyqQD7TSFb1Vi2H6u6ry
E3Rlgth7CoK/841K0iqbT1fGC7isN10pZqbLu5mNlYq+FWtMoljUouGljRNi
cBpaYeA86Z+Jul5UuW0Oo5xReGXlTD2HIuwweUgjSVWR7QD8Gv3P28+OjDgk
amhe4jzIRwt4ylV7hwvyu4oJ31awdJtJOV+ul4L7jmZZF+JUTJVIaFBP2kdM
Qo1U9RmOPlh7v9PUw1bO3cYuRFD7oXnZSJxGgfR0RzhoAwIgDSYsrcOFI+ZY
sqfV4gu/8AGO4nsOxqvP5CsI3tzFhzEOPTbgjVgba9YIQyTb1iO2C8g3HVbW
WzLNaEkrjpmvqggmecv0l9zUokPF7/iSW430YPxsf1gbPmQwwxvCx0OvZwEH
B+OinFKRtC2TLQ5uMmSoB8rZsIdUsbyJutYd9PkzW2cJ1D5Z1b8z9t36BFhc
TVIfLJWw2RFQ+JyUm0V4GNwsq0SeBFClDoYaSJxGlI67KarSD+Ca0FWOPy9c
RNcFIS3iVO6UOoqapw79mgPTXVUyVqEPov9rWoprmJSzBtlye2Yw+KwoT7ne
PcqmEgazA97jQbPlq9FmRU5e9LMDBOVBdJ+FlPSkRuNBABjIn5xH2VTgaKkE
WNYdZdjXoVSDHhghAYU6AlCPRoPM8DeKlyyrkQLlnp7nV9QUaS4y3BLvtHmO
W3sH6god0iooSfJpUzER4FU81ANslkPUkXL5YOHxhzYcYiiwwHtqX1F8C9QP
rAL4TOk/xhuVQtCxLonrALVEGGONLooHvG5hcahpDqIbQmKTR8Quw5nYg5lD
SAwRW2pc6/2GBfxoWHqw513NWvUjCYqCj+Vv2uUSixrc6Vr82YaPU009kbp7
682G3sW7zXU1EZeNYw0F484L2l1XiYFD7VOhzI+aZqra5ij1yIlxu1sK7xD1
izGSSP68kcnAPVbr8+bmyjCxqofKwe/JjS+f/zy096oXL+PFCDPAIkZILsjM
N7+zpsnl3hujfD8vCWAa/CoDeOO/t7456cEuJKnOf0rbIjgdXAC05JoW7kNk
5rvmPe3+7SlVdX1W4BPHbgX3qvxW9+dEaJ3wu1OusAh0JnsMITIPLKbIYznY
RzDgTXo2ZFyz+ry1RdxS49FfdZflewt9nTG2NPyty277yghigzeyRySQTWHm
v+X93q31fzwbJ6iWCDqx+dOmkBSE31JYL59L7+m2cvqbWo08apNo788lK28a
jYD0+o5VpNP0870lQehuDeGBA3/q5EvW9nFSbnfDdcxrQgUfyYYKiQ5/1pnP
wCZwu/MJnw0noyZA8fc/TkXBEkjYJ7RAcr0Hk2VE+qgdoJbNqKcUE8RvGMN3
CtVLEg2Jv2CjRranrQoDG/qLuRHNrBxTW4tWdGY4DxQlzw87babDOdyRM29R
ISu+EFXt6N+jDgcWG1sqqn5qAWf2N7nsTOQ7trlhCxcTnDAYXWGs/ZgWXdip
7+VerP1nVejL7v5MsXP1tmm5u8IR5UXI6LvOmzlKh7/kLgxbhxue8Z8gyWkR
Ta8HqHN0KIf4aznknQRdqFxVFj13jSzT1ZMWG37l35Oz//xjuTjePDBnIwuF
QbEbyts+0IvO9rzs4/toxW0W/ndyeym7RPJ3SBI14nX4kEArlGBD95c/Vvm6
yoEJ6uOpan8HGmYGS74DfqBFR3JA4HfyAawecMXFEv8hrzT1OSo6YoHnmTUp
jb7Wbot/wTZD8Sn+G5+oXYCpNDurXpV35H6soonPGXOhxq1jZ5jI5EvJAiy1
6RXUNRGdtmrns6oYBVEQ0+rFx9zRVM5fJxeHP6hZ5I/7EMud6HAxfkBN2JRN
3riTz6QiMMwKLo67pQCQUpehOXr32nAerGERB/HtTwIVVzQblfkrrD5NRmqL
K3J5mgwJ1GYw2geVPMeNnh8oc688qHTxq34PQ58DSLW5e2PhGc3n0hMG1sl0
lftl6rfm9o2QVqDlJWaE8yDffX10YxycuI+FSL33b4rA9nFBbAB1XZzuIxx8
qCfcLR1y5wIamItsrdiV670Rb+XsOxGLpYqOFB4vhYBpwxT3/IhNQebiIO4n
00Eb65iQH1RVmGLCbgrhWufGWEynHrZjUsFPvKxtpVHrKEmlJnGq1RkcU6lp
WHs0Zr9xJcAjsQLPRH+VGcA7FXMj2oA2wIz7IvHst8OxN1btrKcHof8ZrCpv
Ra7qTv+30b6PALu1OP1KzhvHZX31S0YwERrgwTwCbVDI28XdEsRAiIbROgof
GOiL1NqY5W2a5qRXoBr/U9uAlI6sjZWjudQ2TYEWwH7Qb9vf+GZbTmbLiUxr
F4AtvfSqsouTNkkn92eL6MikNh/E1V87NaJ0OpiQDlGHb9PKz+0LdSCxLgAe
HNfHtqAcmAz/MuHY4vlDG8gHeGpvXz1uZ3Jzyl6tAUS5D5MRe1kv6wQZ01xD
LsZIjZ9xMb5UNFATwqg04iHayHRXXL2j1FPf5PaH6TA9NWw0En4YqjEu7nbr
BGZdKnlHNXKBIbwaT4xxHEt+4w42ETZt7xX8Z8ZPm9Nc2xdyPzF5IAKh6DM6
rJxezAw3lMC/7IpZdtXknGSKSTEJbCjbYruJP5FFQDzU+MkcofiBuvIyuFQP
dDPlkHMzts43FA0pQBSPQTEhrzqFh1TMjoNgtqC4ywvTxXMGcI0yaHE8+arV
lr8J0/VgAfAT/meDxBIb2CsX8P0LVq5PH5Uxeeq7Vmi8H3Sz1htQoWAX8iMX
/nGD24GijM9obkP8GSBHZ4lWSU3dDYuIsPRwCzF5NFD61HiHCjKS7UEex/gY
4cXTzWdTHvC7w2P62ldQngVTNUYaSQiYMX+gziBH0dvJuOOAB8AFIiJFOzRl
zCpQYGLedBI1VtAc1Sc+zR6PHlYwhIlaoAWqaZyu/Tfwtd+iVFCK9YQ3vMxE
JJjiXXYKKtGsIuoqpQVpc1TWyJpPEivXbLjD2ahd2v9p+BfCsdT8zbYWSN4A
yn5drzxJtML42UNxp49wu4+4ctf7D5ozXM9YY3B4FXz9vHpDH/pgpbdqLM7n
zhPeLi5twNVPabYIsjwUgs5Mut5K4WKWXlHlFHU8S2fLlmXSioeYT4gecimU
85bDnqbndrDD6jQNn/SvkmqBCG4X/hzTpNyqU1XlNUAQuA+/drgziss6GQN4
vBku7lx0w+phhMIo9ncdDhq5IjEW9rAxT0axkBsr7qifegkcidGJxOoXzgAk
Lz63AC+cJZ2k4eNVkGpgy+wZqkjLxndYVUkDf32QdiUyIsx+ENb8RnWxcVB9
PZZ782jd3g8biPCA0Qo3oB/LXMGAffpZ1/wo7xBx6Wb5wYyTJKdIGGXCUGaT
MgshcFs2sTA28GKYwhqi1qHjHXVvDUpC0ZWRrDzgM2Ye/hAPvxp3J/MQkrgm
2rvuB5iGkZo+h221nAIFQwYba1YyU7EahTABhVvbeYfZ64ljg3/sL4IvJEqP
8HLJ3BEjy9L13+yg5ipJs8FsinczlVdRO6lx5wLkRo0kFjmIkPwHDmkgn5Dj
q0lgJzSR3uqaJuS+jpoRSSi4vjM/5ZKopUdDPMPnDnSpCPARxWl1D30WoDqj
YN+icUYp6P7w4c7772WcBNeHcCC4yzUSrbuix0SIiIgihRkNhJwTK7Xp6rWm
1ChkjZqj9XgsGMbY6pZaH4CCzKL2vtZQYW2NFkkGJB+wmO5YPfkmc4+wtba0
3X1ZD+rJPGklzIVHMWGa1mh+CMjmhAAmVk1nafzGCg4MWU6+FifCEZnsn+z8
mBG257OrnLzSfsffUNIxYreiQjgCzRu2HrGSJ0pi1B2BM5L7eoHnB5I9CsHN
SkVB6dIgD92gtrWSxhVmR6jCSyMj45LLmJhmZZOfD8kY536Gk5Jx6qD6qJ4B
49c6SzzcSENIc5YNr/6l2MabyroG3BnmN00agnAsrM0NaHkszuuZNapY6seN
52ZsAL+2ukK2ZiW0QxkKwzWimRbjHknpMVyCoYtdXiqxPzfqkN+h43tFA2U5
0e4ktq1kyX5HaH373OGUgMGOC/5Ji5MWWQ65SEtA7w08KqFNxaMLCrRfsPj8
P3bRXyylhPgnQ164HhBq7CPYFqUQ37e1x1YdAj2R23BD5uYS3jKzScD5SLsl
44DC6X836FuO9fc/1zRuU+5fyz8yWHusbLWyGBGlcT4y1ILerJn9VD67kE81
a82C6bn0HNy4qbyU/UcpgENMBWng613hcKzlBrSWpu69DrUM8XQRKCYd9Yao
y7kJtMCAvGKHIhaEiRqhFzbdbGG1wUbrmTcW0sBIxUMPTmPSjcIfCiUuFB1z
t1WmZo9rVIhq5E8lB2lL6Y8N/4FOdYpMZP5ND87I8hResQeCM+1vfs654W2O
VNtXP6GZppgbCOzooojSCaBTP6b9CA0sQ/utSm0ds3a+BaCBXMgJukODrnvR
23PsZGUnsMUjx7tbUJRvJuvYFUjuVmHIEFGXD10a0oC1ykxUmLJkBC0El8dI
JwgrU2jqVBN1S7LJCyZEZ7k6sObnQhVG2zJqmXVf7zPUjmxzmXIdtRPDadXc
ImyDwV5BEsN9FtiTA+KvofnBVGZUK8/vVQVvC2oftU/uY3PQaxn1gTsYnEu9
u1WGUyju0TNuPKgvI8uwWCFomJVNqt5JqeFn5ltjNZTMo8KoIMwFCFdNNG+R
qADLE1BZ77uHJGPNLr/uBBPbnjGPU8bBN7QPV7XQZ33xL+sMWUUe/PtWIxMr
rCQXL4Xu0bW8N/39spfwlkvHhtgE9Y7/eOsIjldAl3qrQ3xRWf2VDYX3Nn3i
WpfB46+pDP4mDuFP7w1zq1NZYYUMqQfPjqifJQhrZv04sdt0CrFS6KuB6Mb5
fPobXOpvD443HsmtqYEMjCkLcltHlGU+TCpm9P6f4N3RXCIJdE/wTIu0lhjH
3oQBHiokJ1qzZ2v/bl9Sl6d8z5s5e0voWCazVuJ1WOdbWjda+fophq0WgCM1
h6sHJr7Wfhw/WJWtslM4IYUqnPUdxTYJ1BpPj46i6BwVz/NEzYI3zyP5qxMF
pm+vseAnD2GFfsET2vDlVt+oP8UysAGdSsyJwVodgiGqQz9+HHFrIKDuTeUh
1gwJvD5rtvlpZ1vy5erSFINVxU/PxJzzfuaBdiLesKKOrpyxa9fSJ7kJr3il
+C5vFBUZUO7FP0uy/H/sLsLK8jv8hWg5VtKvdPSnkAE/GBwr0dvmtji5fimx
6PCjDEfcOovD1v3dca8UxTWIvaUJ4/AzKnmK9W4SEUZM3W5IA9PCw1QEthZY
5sjLXui6OuyxMQUsbhEXeh0+lDg2bdZmvV5JvxdBUgfdsl4JswhW3mRewnjF
kMjPvZMiK6Q5l7j6z9i9fyowF8pHSUS2ZHzEThxRF35x66TvWXP5mwL0JQEg
7zdmId77G7PYDogd87eEOL30eREgU0WwmljYSlsQORP2xVR1NoGw4Vli+FIO
EHhtBnOEyom1BiwNmcPwumIOdLUpuXfw9jVpvR13gUCNvZvbyZOL64u3SR18
bNGKyARygnrQLh9x+IeQloZDHYYbI/MsW8Gz85t8SnAtoXE/cpy7DPmgRxv1
cKNVL20yw/zAVdNwYWbCU951+NrNZZG37bDmhLqp/QeI1yxWvDwNvH00dN/P
LCGrT4vZKplJk9VyQGzu4yzt+CRl3mDfEQ+1VlbkC8wcJmgZTD1PXYitsuEq
5gVTwJR3v+cxZyxu35BH8NizJs5+n9UuFZotI6lYjOwOVB1Cu8/gR00CbcK0
rz55cIzqADCa6iro5gbL2J4guDm7AH+P60+Bwbe+qAinsHb3f5PqJZFlJ0ZK
QOYawJNcQ5yFWI/ZVDwcEZ3TMBfFUiZgo3utsQbPxrkwbRCu2oslD5kmyyjd
KRJkwMNUQm+ZozcLIUqRL1aN4Ix+iwTvhnbK8xkFdsQMKL8LKwcGACj2h8Th
WqTGasCr7vE/rfpgpWKC8MKuKBgcBclJcLUUxsacLDmvBMCQPW4+tmEAtdkt
BI9Pzh4MlbjZDq4i6Xmv7/zp9Aev0GnfpNJ6/Z/Qnw96S4ChVjAOyDQjZYeA
BH1qhANZizEzOBUrHNftYmVrz3L5XBNo74z5DgOeQQVxZTkc9jC/JW+6NW+R
DdWrfX//+zG8vVEIP6xyucFt5LUBYvLK57I2JMd79x8LDWqcolQ3NTPyeZLj
yUCg8SmOm/eeaTBsgK2hpUd7O2H6zI+V4DeSW9rO5wKHIljwb0c03mEm5b1X
NZqoQAsf6S70UQ2g6jxVg+3b1ljsXEIhTbDZCL3wO+dO5kzb5EnKHtInCp5K
SfH8/RM5j1SZyTWAXgQ9rcIRbkm47z/G6fUVNg00lNc/bQxeP8nbaIzh/K90
94DOocFyMDVcbhyxRmN3kUdfkqm2JMrAVuh5RIf/MjqP9SUQOj+eQ6fcEaX1
sxKyOUxXhrRCFJKPbbSSWlcsuFtRPyZgs2SmXKHi5Y3/M9qwBauzTnO4DA8N
BhuMdzOzpnYsEqldRnmTO0+d55vPvJhtCVCmKJF9wa+8hoqRDEfDA3QJ3MaM
mJ/denyUOZebyTfvjYkL+KcG0zgrq7UvXp5y7KSApkj4NthHNu3kOJ7sT0Iu
o4xKNExBmehQBZz6QPLCf/bdUKWwExw4bcnAAiTctZp4ZPpVanZN8DKCedJs
OFpJg2+B3pId+bVn/ya060jTZNNNT7OjyHMw+IkyZC9Q/tzn3TV2sGLn4XMu
IIBD4ahu9gsiyAU54iiocDMPu+5ey9hmbUwl0NZugSvU5kmpq/sMTKkeGfkB
N9syoAo1osp+S4MT59K1DI4VmOraM4pA3B9ZVKdv5ksciTk4oeTaMDhYuP5r
F+XkhVVf0LQ+ppg7xVrW8nD3dPD/HyXHWtKn+teC2EWYDjh70revrN+DxZV+
+Kxl03Pr96SQ7MMwy/WZCXJEd4Ok9NZ4mho7do+Y8RpJs/APWXSfqFq+RijW
4s/zYKEEhf0mCAi9PV+qSiMCiARm/KuIsz2fF1vTHU2LyhsYfv/SWIEeA12Q
wS4Va78sN3i4POoH0T20VguTB+5lv2C+VfcL2P/hFiheYQCW4nYsFH8WM8Pd
OPv/Y9Cb1DmCcOmuIP9jCe7wyntd0XIo1gUt1yHAjXZMq9BHmT4jvrbdzJEr
sgn4CDVsx+BCgcwcro0LqHp162RmhnKjbb36Wty/rKzayrVDJf5nwfC8Cfuz
qff+Q9D/YeJteJqVHZzAVEAatGgY8rIzXsNEZ9ddd1rdX5iGywMl+M3fUU3J
L1YDqBMYNB6wV1C4kWbvSIR4+ocNm7sdJlF3x+hWDiqMMG5FApgZwVXHuDGx
wbjLoonkVODpY3NKdcFp6lMTCAFYDuRNH4YrmWKcE1xku5sSdNWWMphmQuGH
mlqD9nD6iMr5OQeIsxST2AngKVCrqIHW1DzkKQio2VybCsGT9SMCKxMtpM5k
ivkSGXyqNXRsyY5uyjnFeGyltBEUOS+wmHbTOe/qdnpJLB9FgcGbidtwvTIo
4sPHXA8kuNQFEhVGey3O/bhk4PNhbhAS6pk7qDcGwMQv3gdZ5Oq2XICbDN5t
nuTyBcIM/D8CwWZNsSm6w2nfTVCJ4mM/8n9h4NvAflHqyNsnfEdiCThKUihF
aOissWVzY4hu8/t7orU/kzsREqh6kjlRCmFT01nIG6cel2AHMbk8Cy6PBxI4
RxQ76CxhSBSkNiJMlf+fv/QGgLWX4JNW5kFXb5vuL+bfOJtzcfZ1qaEgIL1X
D6QKIR7ubNnYzYrufbIaw8H3nFT4WLbKFktq9ZlV2b4pWPbE1oRX1b7bDpIG
a7ODLPOYFDtcXB43GgQWi5L3lrWBaeyhopmOnGTHhHMBsSxMRaHZv7yxWjzz
2kxe72OC41rO71BTsodpO2TTFcXwL/lbo55fmskGoNDA2gZK8K6n8NqdgQQu
WYqfrgtYldxNcoLzLln/KDo71BGkXBKbFRxFiyLk6byDWj01pljfxVk/Zk04
QVOqLnuw7anXZcCTqUZFsgtLIMai6vfwqcd2TGPoNloRMxAzfu7OTNNKHCni
oE6btk0YRunQSqeMWg6RKRP2QPb9gYnJ2aK92hM6x1AFcqylGULMHPEgZbEb
bf+hfPqIf/1GvyCnhwBNNSO/gq8kcGdsA9m0u9Ha40Lvbvy2BGy2stFpooFt
tudmClNnb4lMUR4Ze8E9YYEdEqDUD6VD9VCC4NqvmFBJveX7h3Nk6Stv1gCj
S4GDJHEip2ketMTcLhw0LoUSfxjiAgzUp8lVfyXw5WBrhVA652IUcDCQuOzP
KPJUKW69OjhJhR1cRUVqJuN+PbCwkyFcQG3nnokZyo349eDZ4l12iDwPGh2p
P3bRhrDpf3S6POdHktDNfYa3INIJ10SPRINOWmJKJMWK4NJf5BVd17HaOfNv
V8aULHmHnJmXOqz8netc0L1VY1GdtWPN5RgO2jKUr9BgzcrBVoA6wtGXIsBH
7B0Nrp3cELQOyUk8XKmLiNyV0YT07O90y0B8DLe9aucyRHmqbm+1JMXKCxvL
pEj+qqZWvZwBaQogwPNhQSrh1Wg53GZFZifNl+kMsdKyaREgDX2LJJJqMuPT
QEY8FJTwQhnamL2eN55JnH6SzeicZ/t866Ph36tsKpbQxOYbdTZd3Nss6Ay/
zdEOkSC/0PpzpCTggQc0ouZaECe/+biJDCyBIPpKctU1hc3TJ2McnoCI5vvV
e3UBBqDSPi0j0xVKaoeqrz5DvAPWisjdOH97RBgxem0XAnDaF7DdI6/4noD6
M9vj3ey0LdDh7n3JgSUcoFWx2i6f0Tm4j2ky1OGyhblO6KnS6q0x8SXWwlWt
fYTXBvgcrtjYPL+wiSlGGKxtCi4v5ovn2aSSahUEXtf2UKWL1B7NcNEMi2kX
qi6bOIQuWHUpSrRCxt6aTOKQd9Vvz6fT/6qBDjUQ6j7zgl8LY8S0T82uUXEd
CNSTRe5SaPwynsjUHkr+aXUgJ6Eh3b51nCPkqFEvvSkM9VRrQRXfxuqR495Q
YQSsimnoOvRcUKRstBQQR0x9HJicdwEPL5pxIxuSjdgM/xbu60usavHmXlUY
yG84BTnIRcjAQ1MeZc9EoSs3jhfNPzZAU5rPhEhWruImgfueysc9EdGn3ONv
+//lqRxk4pFjEiHdLwmiy4mbH6Q31JXYdT+TTCdz6zJ9rGRGQvvBaAqyk1LW
YX/g0VhUqRhvTPNbjhxt5sANn0lCCLnAPUBGDS3Trijjy9ScqY5Hxq9zZZQ2
Mi+3FOoLjcr8lHNA+zYWFBp0WDboc/I/DHSx7AinPNvs+RAkD/VHhrNn3/7c
fOhlG9ZNFj5BLtXnampgy7zTYtQnjpYNUXglGjF8K8JmJgyq4arwz0Js+DrU
zJNYE7R32UwFE5SeoZ6d+pOec70uplW/wzDtrVqPCsjmor2ETYIzjzHH++nM
L8mrMaF3/KuMEJXaHRc/DJDMMM/VPxdkbpVgY+OoYYFI3i4Qb39UlzrVQnHh
xPOvFydG9lG3fj7fzSWtFdYYJHR89IPmgwQFKbqBFV0uE46yhCyN6b+Tx9ZG
vekMqyuDjZFW1K/IV3PmxEDNPA4xoMHbCu7zRxghpgNgoHJPcpBvMO8uRChD
GnPdcSXrCXmGTBXLWNHval/7NYV5LBUjV4Vx6TmJr9B4OIGsSzdboxeESb6j
0csQvtORaWbdkgQbun6D+Hwnlae+u4JQGGQAubSPq94XEkC/0D+Mj5Ab7y5n
sEbbKxtGd2q8mM7oBcLs+N4jePcfItRaiVE+upbER7BeK06Ds9J7f4KpuDUh
SUO97m4+xZYTdOtTcRsfW/r3Q4c0J1AgefGxXv1cBZV2otsaXEwRYnep12H0
KtFI3mBmbu2vZWi9tFOPEqMZn57zNOyya8SY2vheWza7TM6ZNcwqyE/VlPS5
tmvllAFpm4R4EzstOloQ8F7GVfk1DjEiv2XkU1T2vqpm96Eaz6TRiLYCAdjX
QFdJ2HLQgWyTXAmcfAF9MGpcIqgkN1pQg73tYWXTDCB2qT11aRx2rN7Rx80j
IQ7frNugdFIjYF+5+U4DskRolaO87Qgm7BsSJGYXTQJmp+pJyRfqsU7De9nh
pHpkHq6utLUDK0DrE3gYBYFB7xhO2+8bGxzv+iQBQTODYHwuAGSFKQGSBNTp
hgYprcGhuxYPLwiWsEcdmInInXALeSR8B6EEjhP1O5C4OYEQAi3effD+HlZa
yXt1mpudKjS1ynuD+NqmGHouD0OxIe7PkCd5IYDkV3nHv9YzQY61fmVuDm7Z
R1QlfYm0rnjbkGRevYuookFxIkveMM18MmDWOKYmX+qIxKP20qMc61OvYoTr
qGH9A10vZ1jbar49w8claYXsC9tJubdk+9FdTfVnJMPWXpxaefwhlqQws7hG
Mh6XIbxuTRfQ3xdn5HWjpzxBObF8/I1PXMCmXhOBoLl3NjhPvXvHj2O2jThZ
fpuEELQd7jf22AeU4kx1MLSEM6uDjtMK2owiIop9ZHleFIjHkRfsPfMyMWHb
0aAq/Xxq58MBdXlYrAPU6zOPdFJbEEGpoCwHEFFNOIcOI9/64gYhk3qVZynP
QDSKrAevaE7g+BaZU9h8B61EZisDzwDoQrDS7YbNbYOPrbwjBFxXPULPu0g+
bmIzx3LPnEjZRy8Faz25Sug3EvFjfinwG+S+C/FKyXCohfJz6Om9tyzoeyLU
QbNsTJjg3+3Sxbk1X+SAbYOvunVJ4EXMfO0tbyxS2rWP1Pi8TNof80n13l6b
CKbkWAHjyNFGnMrzG1IzXQATxp1qE7aVDkuSR8AQdsbQUuv8LFIj/lwuM8SV
dh6gWWCjJVVqlJk2dlykejM3shmc15xLwaKqfyPN+5kzExDbioOQVqcjJPc7
pm8fzBvYQLioRIP/ZumRgLe/TRQReZLFXs2PxovxG/Kudg0fvxp7wn3n2ubS
PUkPZgxrbomoPe8qrKuDMtSrogRTRJbC/b58HvT8DxHFvv4BjqKNJ94D6Onw
hcaPtNxLxaWzjyMgU5Ziu92VZabp6PYIZ4yuaEy7gk2XDmbsc4/62gvBON3i
GG6WJq8gwuRJu/jEWv920rURznEgHPk69DFqZ18gWFNlfHuvM0/Q3SASWHp9
DZewX/9MPq1UIi6fQu13uMkDIq0b1gxa+OUkI6obSPpsn0PlnEwehTorjJ4F
UL/zRvhBgHxVBFae3tgeIc7Qrpen1rXsD7xzF80f77L3wqmhFdEGl6pJzFel
OREfKJZgXrjOuaDM4ARjylYAfae1yCJbBjJ2f9+RMmvmCQg9sU6D+TQpy3Gz
xm7fCDbuRM7G82ptX9ubgAff2kHEBIe1y9pT84oAzDjzJCryDT3QBOuQxVdf
hBYU1ajC70wDHiIOVtsij93nJII5lAk1x8Xdg4pZGyjbx1HN0qxMCXuv9Ibw
6Aw9YAOTU7L9ZY3dfTBFDuwpuwiRspHhV6LdgvhctzcrFxqr41DoNzBPhOIF
nQIX73rCca/T66YRp7YbtnEglWfhixwfn2WKrR/Zjq6xvSvDsuoz7uN7M8j3
ghLSSW6y+6p/C9hDfMhNojxE6gfFImYGdz2sivIsk+F9CfR9XEOCY1W7fh77
1HuzXoUH5sieasaUNiQpmuNQ9q32o/gAFRVUi1dz0FO2UvdBmVI0LwD7L9vm
jE6APqjOFUylz1yxjKGUgtyOJ5680jzs3OqfMytDFxXhYgjeY4LW5V8aD9Pa
Ki/S0uIUUjJfhFNCYWSDOCGezG3wBzwM8F/EJETGzH7UC1gm8zj517WBmU8U
qXlX97rCW08z4hCJF4pc4+iuBHxRij1yee8pTzntz09TqywLEcHT2v/1/hhd
wGlGRQYB7JYbtByyOw/uSAoPfnhA5R+pPARnfPmqOWLTflONo8qlFUiaWatp
pFgWXxLAo74Z2l64KiJb9PO49vowwcLIkcysTKEI0vEubroQoa024o7Gsc4S
duVpTPjxCWw4v7YfZEgupK4isuawJTVdKeutZGu810yOXNCobzaVSpW8/al+
q5YY6pQIbnAOqF2FR/ghYhr0i0Jg+okki25SDCpPnIakTdo/IdWe4bt3W/Cd
xcFGjruBHAd+7vdR7fqN3FBtNOKzXdXDIkaAKuK5g19+g0UQHJOBoYa/UUGP
vF4e74XsAUnA6v0S5gEva19KaUivk7GWxTkykRxn9pJQB/0UgmX/rlRD8h3H
Cco5X03+2FORVHF52aaEz5e3ReIpAE7XsYjT++UBKjLexC24UrrTxsXffusY
pPQH24WYp6n/nB66z3BGkALHhowykRFepCqNtMA69nNAE+tOQkdevd2jj4ir
kbb8WHFxPLC9QuoufEVg2go9m4EZJ6+l8dDlBHi6kjcDrx4Ik9yNWQV6dJFk
Uu2BwsPl8xnzjG5XxxyHOQAsRXEXpvyW4FGLWEKPZUarzr4oZoqWXqy/IZqg
O1ygcb442kx9HvmI1VggjtL0yPP8p4/tzlnTuZRWwjFbb5GOflbHYe+PX5cb
rEvdEcsxZtsqJ1D16l2FhH3qCjsytw96Fp3bCHAQnTIlg9RpsloS5T3zPkaA
/whYYptExJjLnBWwID1rTm42Fm8urQfdXuVANBjzRd/gVgV99wXUGQZY0/cP
cG0mvvuwyj6ecViXjIOw4iDX7yZND5iJpv/FoKqwlMUau08swqV0Ah+lT17N
NXmqy+7wYYm4CpUksH0NwIGoYcLzzqLZUOe0mcxalNZJB+pX6IT8BI+l3cgD
fKd2/MQSRQRX/d8Tu26B6ydgA2WgVFjA3CpiRhEIVPpFUroaxl8IvD5tsrWE
SZxpqp96/NH5Xzz1ljs9PucvO/EqYcrMZofRp8Z5SSGoYpKrElymgraDybED
YGjAtHdEzYEI/DlEhAXmaz3XhLuIt5RSYJICeMyZqZUVKsV75I750hTOYZzA
rTg9CKA6wP68QNYRwPzn+9AqarmE3K+GbFemGyX3vNdzX5bjMf5SNn38wTO3
NDUAkmtwOtQffP4jO/rWHO1dpicHZEPJtdiKhEnYnueYxmr1rY9/jNd7bPA5
N1qGvza4aJslsVxJ9v1fsRLtrj+NBXdzkJjewrh0QRuKEqLC27WllovsWK0E
nZc+L0TP/l0gZbRQ15TAtXTpyLUh07+kqs4jdFI+CmDwa6xx7++91N7j/EHA
1eDNrF7X7F27taiU9wxnp/MlQfrUY3xkoZ3nlckL4hko+3z7sGvfA3l7iq/Z
/eWGFrGeuKvoIrup6mZ+Dlx5D79wYT03VXxVUqkJt0YdnL6rgqdo/tk89eUQ
XryMufjATCbzBgYzZ4JrLLOsNedRSanPM4Jyr3X/sAE/h5cIpQKtbYrU6vwt
5ZUcyFml7hlxRofme2k7XtNQ7U0t7HGBP8rK2Op+SlkfHrap3uUoYb5ujns2
UIGi0T0pzLbWtJ4RhmjYQhh/ubQekpYsyG7iiksuAIJRjMYzOu5Oy92vxv3k
Vhn+wCQbV7DLpKvA9GeaEgjZHMQ7UrxeDRVWmy7rsy44Ajke3oJFGMSG3aVq
jYEfH0wWUcMmoDRr/WA0BRvCaD97U592C+cT1hF3oXYh6CpcnI8auPGr8XHu
1LyMCcdN2QCS8ARIQLDKL1NybBp9cEEh/I/Tq6P6GoGprMv70FwAxvH8Katc
7vHjaRk2x0g/xGWD8gxR+ZWayJhIROjQXDz2Sm3GCi6dopibG5Z3nFanqltF
XQ2M0A18YpAg8n4eqMaUbliiTdV7deu0IXI3iRswGwb+KqxaZ3xt5ER6wTnp
NsWfF8se0cjAAbKOiwZJaLtlWaHq9pUMbDIvF7puyu3D1iCNtsdW8zfI3aqU
z4ezYASiFg/fnS5odsbJDwSVhBozq3y7HbTvogoUz4ubADOjet5NxfPs8Y5Q
bhqGXMGpHK5Q34mDRgyB6THnf8L6V8DOWvaLhfM3a/xx1entgFKP9ZWe22z/
tJG0Nf8qvqHyKLJF4U0RxBDRU0bf1btTTqXumQ4GX2ocuCoZACsEaWuiwDRp
FqTNgeA0FilH0dJHOwsPR5+aXjdHFxCvKYsph0j5B1Xm676wEqttJfVHNNHd
zyMGlBz8XlCCWZClFA+qoukfUQ0vU0syqLcuZw7iJfB+rVpfUmawYje1N3m5
MGgdtXtvyl8XoJY8B4Fumb4AzBXKnV576aG0A5AANToDtmPEfbXIooWNq1sS
LctD55RZcA4qmy7Bj73rdRfYPC5dfrmJMNjL1rouhTmwXB49Ywdhu1jybUm2
yrxPw3DhRdBkzdmBBNR1/qtGO9m558GaC4n+7LGUQoyLPBIdlHgGCYiEL2Sd
1wNT0RqYiKlW3vi+vxTPbOaSE2TQ5urYtJ6JfWozSebK6yj5529/EC49npUw
3RFVNAjXbA9HtMlrcCK/U0Sr0fu6Twy/gUrw82nX8brxWyre5GEzfbCfuLAU
qDP0gGjyUep6sZJWfTuPMp8b59tgNRWBo5hcNcTTpTc1kSMOQj4SF/7U/F4Q
ip0ovd6PBkFLYjNBQiuYNhDPmZRBItOwNK/1jYB2vucqGYwsSrlA0sOohNDn
vGOB2admcldpRBcQFaNEFBZqzYie43J/Vd4BdoxVNnbNgR0WCo8XfdYD+q2g
YEpEyNFTdjjz0JZt7JS3a1gCF99nDS96MuvOoDM6Bmx9LTNnsZKDMVPWfHyd
5aZjfS9inaV24aPnIpPPgDJBo6Maua5Nzb+O8diDG5aOcIfWFlll7s/RfHBj
32M0jKgJcSUxrBvITwxuf1z8SCqYCVb1QhSGsiPmLxAMmpYFM7ulaSnQTwNj
uShqcSXyAEAvQYlrad/mgFKVzlGHLfJPcntrH2xFLE/GJdEIMWqz02OPrX8R
7Ozd6GfkaXjewAkyFYAB9UzsFiSQVNapClRiN9Y8PMBm3Hp3CLsT9+2BVx8+
q8GxTy0QrlWzNyYRoPtN3eHuZfNkKyGW4f/iEpzEE2K7ijoEolsBYzrPxjZl
gk3O++kpMBTfrisDQR201uSs9k8Xp+/raFjd/sekCnuFYiKQjDIt1NjIMypj
58ghwyFTBRGTwUNlL35r5KZahI2fXV5a6/5RfEOS73x4dnvZY+NsDak7U+TH
oU79L30m6IW/QJgIVTFKoZ7hTHsyUuRhQ8P14CUqMfh4xWByJ7zKxlSU8M5r
7AaOMe4uOyMvRcqc0jUOAiHDgza42tvAHKDgHTObAL1mtsbqLeTx/7wrf1hN
3QQtwQBoOtB5Zw6+2w/0xU5DeAR0XKzfRUgJakAwUvH+moDkHi+o2T8335Y/
jICh3oLxI3qTMpyQ9BqfZNge4KYogLSO6Q6sr4gkNTyDBeORgKKN3RSjDDQ+
OAV6E85gSWR4/rCCbzM05bay0b/kVVyVa5KGMjZZg/5o9u65Y7cXwCZFKjUA
R9eh99T3zeqRiuupZ8VHj1dlyuLk6+dHsKM9zi1nkC3gpOoa3j56eeWq+IGs
SKuez/4Ua/hcgH9oWVGPOf79vKO5jETM4UDdRFigqq5X9q1ksfOaqnKAw7Fa
6Zxw2GHm/tfg2GOYA4r3Mho0Q0BiXyXFmjfgFKUe5huqN0d98ujcReTperr2
k/l5wYUpjpS5FTTwWQENQEB8zH4/uGWA7xLMA3iUugRsUQU2rWp8G85tLhCH
DkZjRs0dK6gcdlUY0C6nBOgEnkZ5SfxP1+sRvShiWVS2bqSMtfcbcfCg9oin
Eakmlz3n5kqsOd8r/l4a8mZq0EPCNNFerq/4Lul24kkkaYQW7PHVtBPpfygX
USGUGK5o0genLQHlS+MXQmzO2XyeGt5KMyx2ShhUQvpZcdeUd2XDynfu08nr
mxJMokOQzgGz7VOTsovdkAEinFLinSaB/4qOC8G6UtIW4aYmC9KMwBxiS/eZ
evhzNLe77vOemZu/z+XBvmpOwfVegECr1FCyiBWKzTIclg/uwGqnrM/joNWR
96BGeXgD/Hzm2aqF4z/QV6Y04pck8ySpSYxZcDLVMAMSPGQAIQXubupzBBz6
YWJutTGMxLYv7uSJNyeDTn4JuZJuXWXmP/NvAwUkba9ArYuwnEKiwL8QJeDi
g59yT5gxgZi9eic39RCskZfP3tJfcUdA+7S9iiiciNRpLewJRaeEPa1iEMF5
N8N0qRfxOAb1kY4HpjG56Zqwg9P33vCQ7ceFt9TOmI+J1mU0NLKUs4UcFp5Y
SojX3EHHFf5f4dSiw3c5xn8pC0nHRLYZ9pTemTKMU/bvMJhJl+E2YWbYog82
qx/EPXwfxMINPxRMuN2Tbvsrajd8jUIJNd5XKHGKSQkBMidN2mgvmAImE8zV
atZa7cFvehgJKc/rraxPl27diQ0D9ZXAsNrkPbQY2qrxm5p/0IE5GHT1TmOi
5gMfBwd//dy/Dc9gDYu4AZT/Zye0J7hk5IiJROWRUMkCxO7FiZemDQlSNS1U
TaRMjI92BfxCdDKDekvI2VStqzdWqDvWJJzPL8gwrjgSmUihEBWBjBimz72d
ZXWvNM6senNms8HM2tQajbD8ea664eyfkofaeGD2lfWzZBfC26Rgr46W9haF
eEqyfDlAQZ+6X4SPSCrE6njwq2Lm1gM6DjUgT08nMi56DXJK4uL0HR/lrfQx
wqAyuHVBEkAtVSXsezYnK3NfR90KnkqF8pRbheT9sGHwVsLB3ZBHwGtPHnC4
2ZF/1AypYfkLnw48O2+zreSDIFO4a/J6vBeyXuEWnDjWnxJ6CZvEGTPFyiWd
ZYmgX/0HtDVwf93pDMkP+eqFCWRRipwjpuymQTDFGz3A3went3jkNX0wbxZd
mPUYAibFp+AqTJf52jahSXylAX2nSWV9PjPTocvHnDPsLhgXXj3fiv6M1ics
GSo5QK4c6Jv2ZFmOejOzJZerNypW+DXVy5xD8oBDbHHJWmlhKfcSjGdrnSa7
Jcq6TVnSExHQgxnfJum4lHOwvPIKoyZEcTF6HtH8D2/pfTt4PsEMCr9reHYu
7j+xlgvpoG8wSSgfJ7QT1zdvF1AhCdGKnYvaIWDysu0IDB59FB8y1ojyeFm8
mP6GmMdReqFIpe8Ki4OL+YkA9Hzknw7pfudpP6OC/PoSp6VlbbbtC6dnmnRX
c+jR8h9M0ffiNJc8xlqIUu5fF/vkOaMPNroH1MBFm5RaIOxd2rJEsiIn9Ny8
LWI2WhCp4H61S5tbZUK1Y3LI5vDKknWMhTNey78nwNrQnF/57Yz+Bg2F/ZXz
Dukl0Y/0E61tlWPg+b9w+b8+pNzMR/NEvyxCTB9t6Rhp1i6aCs3tIboQXTW+
Uo68IyGcGWa41MTtsH0tAWa1E9rtCBubVCCnFFwCy1uevNDMQ8gq7dIE01ng
az6/Cf3zwsfGiYh6N7BonDJWG2FWONL56QoJcwdBPhLtKe6SvXalwbMAzPcY
CzrBz7LsiiEp6yl6+WcETgiPGfJNXH5rfbF/rPHzNg8goRsap8gw2424/W1X
BIYy6lH3kaYDlbSJdhg4q7rDj+NQ8nO156PKb+3rsGNeTSv4+uEez5FNT+pC
zNrU1dIqmjypVV5o8c0AC53kQmJy1wAveyaACJ25ii8yReKtS+/0wEy4O+1M
8GLUs1HGdFB6uHOuCbaqUoGSFf6EtWzA/HAC0XUZD2Tlan1neS4bhdr+KXcC
qmi0XRJyyb1vSB0UZG6QwubLr21xvsKMW8Zgdi3Gv/kFfzHYzB0ajDbyIdhK
2WARPB2n5U2yMF1tV4XwQeSkrKeOWOSzMqbwahWZ3GRYOEjYxb6QMUS+lh1K
g4dA7iKNsYjU/4W2Ry5nS6ucmcuZd2SMr3hEFklcM8fUeGanLO36mlA73jJ5
fP/ETA045LfRVp1ZekZI58Sf7Ot1Pg/GDz1JPFrMEQr2K6t9OeOQMj6vwzaw
mS5JilkdRRY71lADKy6a0uNuk3yrq8DGfLBZfn4Cpn8mWqpB1nJqH7b2M/lL
/S5EF+ZoFZCjJVgUyPiHNb3j/vjBEFhoXbn6HJygpRkv+FnhksVkNaElGLL/
5eJvQPZXKWNWlo9UOBX1Y/eNCP/5jHKtvmk+yvwUwYwNTssMO1dlotTV+fWc
fRqWpK8whBnEwF4TIbsfp+aSYVKZpQ5LCYU0ls2vwlKlqPCzmT/wVds+bH6U
8dva3940vl1I8RsWCv0W4wJLIudInD56WBodsauRlsU6lXAXdqkqi3YgV3rl
hhYA3JPOGYODkjRG+pSL+XEu7T00JLQhZ4w+c9LNH1ykhz7sCGG9rfM6UW8A
p83JDCgqQ8ET0JgeqoaGSnvdVlt7pvOWW8ir5kwnuIFF1CU/buluHaYTVQ0Z
i9EJA9EOQ26L4DPLmqyI7SMWWJnmyFwRoGuVTjChP0vbQPG9z03Ba644bXop
J10k5dNd8vEXFIAyjs0x6q+lFfErtxW8wmFUa9Pal9ayBorBcZFUCWUmrwds
Zoh0NYhvbk+31vW5aB/EhSxNF2N4XwWK9eddauC5/Z8uJCLczxxVD5IyLD5F
J13qbRTQtSBaypBtv89CdHgKdHIxjVcJqYaFPzHS2STFC+tKXdP2434eObDH
ZAn/M0OI3MJKZemTHM3hLjCYsf+bNeI1gW+Ays6Rrpe/W0uGpVWH4wo2890K
eOqfjEu2YbHj3ZGy1vPv3YXO5DT+deWLmLQ2NxxalYP8SlAJQho+YJ2CXB1/
v4QLV2FHqBZKlr3tWm7Z0vTKs3RJyueWNyWvGNNZqgAXodlA1G7uPV7CaA78
L0J7lReL8H/dDbujw6vQn6+apgrChYmBe/Ljc/kDVJZ6ISLXAsBku+/LzWY6
4bUbM5k3qntEWgy6rSyNtgIPqiC4z1JqC5DOwhelUR6dQshgHQgLdGy4qNNY
AlTsxDlGS4g1RqCAupoReQpcx7WPR0q26yE8AhhJB4QDwNoENP0LmX0nhLUq
OPRfZGj5rHk5f6jbbie7GD2RczQ7jG8GobTSRu1d9vFLD8d1o5TsaESEUkH8
NMzx3RItRQolTll5Z9CBu9/8XS6+OEeu0XCob6NWv0SrmHyIXW+Th+DWPfPD
2WMV9fRJ6HRvSpxIBiFTm8CWBZ7+DVQ0gB6Px8gqXYPAa6SwnwOJfLneM/xS
iM76XyhfKVI9cgw+0BBQBIuJnYoQv4szRigYAfFb5q5nHVI4X8CFymmqgSq3
2TaYJ4h2OmFfegRclqUKKw0Hlw5NRGb1IsRhUWEDZg3VQT8/dGUCaQqmU915
OkfYb5x3bNagnWVEc496bYeyxDmLLjZUQZbyE90NlUH+hy2g8D95EYFn1uUq
WzNjFTuOX16c3mH8GGXEVhKQNjUx2i2rdCVe3Ceg+xZUN79rHvXoIb1Pa4Q+
fvYrlRSXAU6IDxBl779W3tNPrkXNBgEoJU4+AumnjbKl5WhkQZ1OW83nIDCr
8h4uUQEIZzbKrFdCR1YWQD1krSkfCOEXhRPWSnWk5QKAyKNq1THVmpKM/jEG
d3TdG7uj7g+Dv56WtTfvMNWQ9xymH+GJG4D+koqLVEfWeLCQiShtPdfF3895
gfg4+Alt2JoM6bHYwaKjjLYI7CHtm4eZqq4s43/URbCM2+C9T/xFRVTZSAsT
7xU0JTUHCHCy/Fw7zYtDZFlnfFboJuRVlJE6fw5c4fhqaJFsAYiqVNp0fOyC
pc9ZoDqph57m8R8W7uwT4rOVhhH4J2XylNmDg6m3cDRFeIddKizWBRf7/Gtz
1v+p8f99Nt54rZ0Yhq3j4MsMw/nOgUrMW4aSXXVtOcGGdLaYSdU3XmdPu6KR
SnIhpT/lwmKwJBwXA05+FhTF5IG9Zzor7KJbF/TUUoUe1FHkbPDTF1hYB08y
oeoJhq3sNdXKtT5kgNFZWLZe53RIpohpSQDdn3CTS+QA/XdppZGDJdlEHIue
ZC/f2+UHPEwew3Ys3hSs+3nvGxGQ3HotyUJ/yZP4UGtEsQ1GPmi24tMBv5ac
RR8fBqo/9uUcu4JpQxnM0VuoHOgX48IPexnmNu28nlwQdgDQqGDUs52z/SMo
FCS2Z1MZQKPGbz4CmUVOkhIfxrtrP7dAPuo66sP0cFiUmE5KyYEHY9ROOpVF
kn98HvljO2/xuqKFgojy57OYZ0cYh4cRQwytFmEA/7OzVkICraDsaRfNiFl4
cO8vc6i790xtMLE/Y0Ru7TKeB7gQ8zsAblANwQz4tEovkRsc2qUt3A3FmFKf
rSt7orCcIFRL2n2PufyeWWsckuzJlegC/nnvIDzTxF585G0xqwTmnx5zXfnr
RDKe5n3cCPFe7bmavAaU8c0DFiwy+0Esoyoxsxz/vBPbKv9Y7C2FX8NTbDnR
dzM041k9bHZSebXO3R56E4MYrYztw8xGKijU2dNQcpTMbpgbZwZAzCs+ZSfV
tI7WSfU8iesDsbgjAdGntVRnhtl4jwvSSbgNVNMdxYj7n1w7HdFXkQGEYQkA
p8yMX77BoB2gMOXvqp6Ri/ZzxwWLC1r6oyWeGllo2Jr5KR+ZonFApz+Dgivr
Hk3NqHF2+BIkz8TgK9xVBAg8viV7O8pMANQFqHRrIv8P8ExV0qHz3HjMbvsH
ftBk2jQMJL3PVvIGo+PqHAYmZKEi8Bxf0D1m5+3O6VhQS72ghwuqLhDeve71
uNWC4CSoUhi77IOJBMsnhqSEAa9zfjDrEHnOFMWKjKiFsQ0QhldBTmrgrCKM
RJHa2mwBTAahGNFhhpFG77q+wTpmWAT4IQ4H5+zlCSiBOtcF+cEOawA002VS
vmzn0XAMIojPdGFjHxv/YXNDCVxDeUrV3j/TnCzpubvMdy8ufUKMET44KBii
q8uUKTSkR4Z06YutW01r/z1UNn1H8xitFk6tHMyNmRihHWr7OZsx0+RkbWgy
TfspmUQJ+FXOkkyyLFVsCJPk2p0yD+eHC7MXcFoZCpVEzjnc+/WYdUEfp8TD
QvfZPrkpR2TPA+WKrMMZGvx9h+++3E2JWQ2D/Z3JkESn5PdM3Xu0fSl6fmg5
kgxSCa6Kzu0bvtBlG6KOVjc1kQQ4ovHaqSLtcmr1g3XIE/gp65tvHJwqKm3o
By32xjBvOog7e8Z9RSMPKuYYBHtAD0L7mp7rBvUB/fw1dPyQFv9f8yk0rwYp
z0wBOINMqq8x0OlL8+c1ZSIKQohPpwbiN9dcf7ij+pGfW0HKH3mqHtVOTRrR
rZNYl/ua9ATHF2K9XWQwwxpBO67py6Sv1M1wLoh522nCDVOTI44/QE7xrbTv
H8pCMcN3FzW2uvKxYDKZkE1H1IaFdtZI0T9LsuhYW3GUe/btVEFRAzG+CBva
BaqIJ0JKUxFFcIlbgFPh7RszVg1WO0U1bYIc2sGcr8cQ2T+M0JJbXB0Su8u+
nJltbx4dZuXZ3mfwPLytBP7GM4maSR/KvPx9BeKukS8lmqvWqIZAYYWrlqIj
SYTvxzuml7vDJhI2jDuh42IFpnDwzTuweyFrttLHclmqnK58kQb3bjQ4EmkU
FArtOt3dWZoRAW88RNj7C9kv+Di6vfYqVpLY1NibE03BWtOjXYXTs6v4BBrw
EGTqPc711S5QLtroJQZzLgh9+HgHMxTDQl/FHoHmBh86kZU2h6apCfyBAExo
3MQjnBmH2Vg05yQdeO2DdGVXI12naJiG1uL3swuQAeEQPy0ij7ilGIgOyFvf
zHjMXJK2LQi9C43qcGa1sJCOuP9VJmBuop2O3PRSqQ9CTJqMp6Wua9MO/fXl
jr9eJiisBFuFK/fFKkMMi4HVFYXr4E8z7xgM77cWg1JYC88iwwpiufJnT+FH
GtlRu0KjJuXwhRZq1YXm70GZgg8Rsj0XIk1t0pEqsk99FRURdCdvkMCa8FR0
u2sPr/fXW0sjudx1V8N76Zlcb1BngbPUFsEBguAz9KqlkSW/xlWz0anZL9oA
w21JctLO1uEjvArB80+3cefllhd+MGhLb3TKIBNFd+4qUfKY/07Y2XkwYaCr
jWrdPTiMFhJHBu3Xg6hW4iMH0Qwvy7lPS7VMk8b47evcfLvNsmrr36tSL7ft
C1s2OLaQAegvWeIDQyT3GzE0/g4+0JaD8PVfdC0BGuo/WlQuxBzCyCJdL6Cz
0chUNfcIsRQC6gkkJ1bXhSSEFoFqKP0zUsIU12XqMOtHoDLy8arq71v9lJ04
dA5Vmq362Y6T+SRtlhIXdZjYKC8SLBzx1OglbxTyN982FRD+LAXrS08EqeAN
r/hV5SkAo8BIMzj+n5W6/6mxT9TV9JqOYL4itEoI71O8xcoBBxYutIUv9ERG
2vkKK4iDrBB2zgccM+rMX6XCaMrrlx+LCxEHtk/uqkeQ5kNulrxkdP/5cApb
WyrW/xazw2mKSoI2aDaCm6voMh4EIkYEQW/mtrT8MKRPXmSG6knEvd5rCtC1
WOUVLeGoKupFJ8AVZxF/bDjj8vcMDMvaL7CPvs2FtLASDf+kGJcGNLIGF1Zj
UbBjrh0GBznosnbO8I9ALU0kk3MWJAfn3fOvWPI0JD3qjCwo5twaZOxIfQj1
ZNg6KNcX44hEB2IfrHxzMiDnPW2kmsZcTMmocyr2Ch0YJNeH6sEYYL0mX9Q4
O6gItfmRxFe+NTvBho+/cE6dnh6cSIXG8v4K4Z6eL6rWvQ56SWvEBQ9SAl8x
DxXIr23yMGuhT7gmaF3Mjq8Y0jBAO9/O98h0a9pfyDckjkG8jnYMN+gg6eWR
b8vYDvFeyIJQlBD/1aR82uPyDnLdcNSQzntYByxz2/sqh5wdh5wTUi7MQhDE
gPy7tu17PXf2QQ3O0tVt46qAAIcEMyuKJEDAmQMW4hq8M2ewg/tbUR1s/l6w
qkhEsECfASkjsHXOH96RUoyBklOxxFq1JFEMFE2iEKUcgal5So4jd/HUQnzT
4RXpEw1ieO1kqxx+qV4jq8Tp8HT2RuQTtGbyS1wBVOTJ7yCAHqaxgH/IznpM
ZksdZeLj4FTTpuMlyRfyyOmTL0O19EPF1qk2knIUYsxDd7vee61nwjB+TfUF
AO5weCI7UQbYd7b1LRV8riBfrcGpkZHPsako0LEowlUso00CZmQu89CHbLW5
rC2QsOwad/LPzH+E7t+ptbi0WuxlyjY+3DrPRdjH1xCQTHEoo3WxAQJVChK/
+tc/txPAWXeW1TLzzNomQmB1w3CglUIT4FnW8leOR6YVh0aJEqjoUj++Ciu/
nOU3oIuWX/5AOJuirldwc51Uyc6HCRCUyiNCY2FJGy6Q8AkT8AyLb2o+fpEi
quT/1hbSpsEu3FiGUg9xUqgnAcAAI1vAcxvirCUhON8gG40n/ds7TDPm/Z9f
aCnau1dWNSecuJidd5O80auvc7fCEnMeUMlzS6A8wgDuQUKQXC4/5Vi1ynkE
urBVLkLb2o0V4rsmyNulni5vLrCTNvZaFomNQuSjbvlGFYzeNLQoF6RB1ZBR
VYLBfeGpcYfSM6iI95Uce2RxaCD2gry3iXlMq/IMX1Z+XL4Pe+wK6wEUV9tR
u0dZGc3yURdzPGKGDwts4P5xcl1k5Gir2/kTpJr/N2CYVSS7fun0m8leNxqc
s2lHfyaVVCwxAEgTxvK9kbv+hNDvGMzFNKg3B21Z5yFlmShjBUCLEwn9tIFk
MvPhOW6CnqW8QXhlZJ8UXDs3qlNG7/dkLS8myEpUCf+gpiCGro2jWPcTwWc9
WogT4QM1RSeJpMqALQzld0z032BVVn1QA7seNAVp3yEJW3A1FiR1FbJGemkI
OD5LLhB47kKsTPuhfduVeR1JHdhtTcZNOlJpIwqPjQbq2scyiWZCECgCtLhm
fABhY54cq+BgRLwuRcCIhZhCALHCnb/Cbzn25W9UHvxGAZerf0a9qLcB8pgf
FH8d5SPDgKHPa0HXyKNiL9SXCs4/YPnfnGKIdeClbFoPBmSwQ0tVO5SqHQJh
N+VUpWjHaDLSp09VZxUWCJYP2E4xsF1u9nxoPubrZ2Y0hQDDlLdXckA6kRzs
Uxlv24Lkbh6lNgQ1A0K77GX9GTJWAp4G0hUt9onQOILCRqjm96ytCAVEIg21
c132o9NKq6jBBnZr2HkYVLmDRmitzTUw4szOqdIvhyI8iQK2tqPpC43SDlMS
9cVJtyjIoX6X9YHLtTQJdvv3I3icuN3MortiZeUNgj8+r+91TCp3bvF3oPur
cQD2fNpUjoyR7o9tItZ6KnOvlnhnci8wZnYusPAFdlE9DEtgSdXgbFHKqn5K
qg76KATKuZlUtwg6N95VjgWC/bCw22y4LA4rnpjkvQ/5IISuE6i546rf6lEr
Xj8IcfqTpd3znhvE9SnsMnp/ELGTYV33QyozJ6P3BNo+0hgjSyXyP29XId5v
G03AeLJ6vC/1E4S1ftKyFeHcNMCqmscbVoDgBUaAy4zkyt2nHHriPh7bc9JU
x7ktNg89/CLoLVttlVklosOtpJLHLM1dHjToXV+sVaUzvCNBzBS6crd52lNg
3jL9M/pMX05vhIyi9aE2Axh/PNNZDzDEgZWSD0oiaJwPPXszu3J4OUez0sfQ
7QZ9YHZA1Ndb4Wmm6nQBlYUHSeeQHB64Ons8IYf7NSSz72sg1z2JBtxa+azx
qzI9UbmtDth/lvRZMsJKeG7G4xkddSBVUZLSIsrZcjytsMnlNpEMnbKc401w
Wy1Mk/rL89M/yAJQukQUNQmwoCmRMPMNHv2soU3Ry95km7pOUcaT163pAolb
6IpQdp4yfgPBNYZk2adOovqdwEQjbjGrSgc9dYW7/37tx+Zns8RW8Rm6eHHQ
tR3ADLzezgtzW7ouv8TyG+Ew2M3jPOQGiBD4L8nCwXzGd1lAwR1+fhHtwox3
5/h4yoUARqaaB80kn6QtJEcLxyiMfDB5vj01IttIpctCkAlrJzfUvo9wCCLD
Rdlxd2N9LbQnnK0n5BYKTcoeLkxwFerKeWXicWYxohd5I0sVbjXZS8T0n9Ay
tLLvBqFIRHW1mz89rMwOAGntB6wzlcxjrxNGoXUg1dkn406bhzVu+ymjOrTm
d2PGfL6J+RD4ta8d4S8evkHxlzqyX4ny64O8XK2gr6UXD66pMNmPbU63ENKL
g0Ihc1mBzbaiTFYYzFLg7tsg4SvroLD4+cHYYmvTZXsR8PtGjove6s0VmDwq
in0SInYe4Y2u6TtakSBlh/CqleZtyQdaitdSM7dxKFayS2i7XmWiLqvfQsq2
VicqXZ5BdaFe5lRhBhQ7r4RU8F6fnLFlbxZ3L0G8gmqO3Hnc9z99WrgJydub
WGO0jkOycQMdIhsWW/yd/jMwp6UTTg4h50gyMLFXZNbFEe+c8ECz8DQ2VaM3
xE35slNJZnu9p2njL0XTAGAESjBJ+xkoZQ4Mx6mwXRHJcDM87lTle3wk//T7
asaJYFdklCEcKtQ7SF2XcWD1y9en/hp7oH4z3lm86f64X2yNRjbWQTGt96Xd
xN3CPhMURsh/IGvJZ6f/7qiXb2ceqPo+iLHys6hAFuRmLVG8qxoO75Z2Y4dA
nceMSleeHJN/OBPGq6LGqD5SwFEctl0wiQcxHIkfxxPz0zqbRTDge+9toD2U
BsrgpnO2vTAf623ALVzpAmqpwPJ0BHS1sv6Bvq3Tgk/eTboKzsa4rdRYwC4k
Xs2AWYHtwcdYRANayAH1mCqqGANiLE6cma1lBcPHqx4VGkFDuO5AGn8BcHe5
I/KBO6VFxbmLcSs4jSXTHWmNqHyPaFIBpatWjROLnw9SEFeqMthCHMz5Z8EU
wsbdrCpCUx5DDyPxLMBrhcqzUY+twmRkylHsQHZwZ8btSFd70B5rB3fDivmt
TDVldi9/MTdvYl7HdzO8CdJcyEzZg15wawdUBKUcPl7bgA4wb/yq/FloG/je
bNx8wyOs8NO/zrfJbA3EZ8jb33KGZahvsYL34/xEa8alZc1cvi6Ye9JPIBmR
vIVkxnmY3hn3eWmM8nSJadWgkMuPx+0EzaeowYDWCN3lLa4u6kwVIe/UuL10
3PzTtZ+kA7k7Ptnrnj1y2POPQ6qWqBqHEC/F7kaCwqBfuWGRvyGvRwOQ1+XA
WfgLVbLNZ6Oh4BwTVEmnQuwt1Tq9wVJUXSk32dCR8S/15RNX42LW02WtS5b7
jJljsJW0QCS1C5VWVTU2s4kDzX3L7UhEouTamFJfltd/OXsNrxqF1X1lO1td
xr5yH9zvqskKgz97RJmTsVQWA/wbTmIoZ9EzW8HC+EpdYK6pCVBaV8ley/MS
XXqGtvHE3lV8q386BRVhdhDAH4roOV1w8wH6vI03TCN8GUjSRYp/s2NmHay3
HrUYAQDxDRmbREj5nMHXAhRgt8O1O4JPjaGh/+c5A3JB8r/ftTNcOTG8JVmf
1RC/Hl1WvMieSB/JLc0Qvv3WMKmpa63kx/VCWW9+OIY/zi/H2uipllUFhA6l
JtOzlH1WBaG29g5JRfYRaWCpn7PH15+YjdZenLJzbt5ihCje0NH6zlFm6BOx
XenQKndqgmq8Z47esVv3LWPRMALLVPX6CwgZutivy2Ud0OD/3QqRcm/pUFWO
phpoBK77JdYLxdE0tiady2g+KF7SqtQBTLNT6hZWy6EGfXgT7QOtJtKjGzMg
crDLk157Ftkk0vjbn6FP/I4bXxVF+W4drEEdr/nwbs1lKFAOnkU+xHrP8sfJ
8mFFeTBRAfir4JeGFc/YQTQO96dtJ3G0pnWYiKz/5M8tUMEjalH2J62QFb/6
Jpy13y81TCAT1aFjzzqUy/9nU59ionu/5cyHcEcyX1CeXHbnxTJ8HDAOsyeF
BPSbqg/OQqY0+uWvkq5vRo7NLo3ZNUxGYsmMiXEaYTTgIN6klrgwXi8httWu
YKAh+gJyoxJEBVP2VzvPe/ec5YCVR+eVbqUuO1W5zdsW4rziF1b/vMszyVII
IFaX1hv+G7dvfM8hcPu/pFxHavVVrlCxLk6VQj/5iN3FMOOwVQdTTEpk9WCq
lRERcwFT9NKsor8occwq7R3rwTPI12bHiF9u/ETnPRdnDo3KdSZMWPLBIx7Z
CeQqEwRP0G6THMvCE+gUodq8bH3i55VSNMo+kmfFTiPjGjDF6vTdOWq9MWmF
IYmLf5nTi2eG0ZTo1EPoN776Dx8VRFatvrArn2u5ehfqu15gznP3XyW1d4yj
/T6N2S2IMPRL6qJ81U4rSPtfwS6dmfCr7pewDMd9OTuqHs0L2+1y8XijTSIb
zasgCPhM31E2ERWUCSGYEX77/LSDmSO5jO2U3kiYCKzehr/7+276n5Gc2z8b
U2t3u6u4lLt+Gg871LvccgqpZL0LsE0UWeuz4RGIgaKDD/fbPb62OLoNkiDc
iF3vH1VEGFN21PtRzlJ6OldD8pxjhlL+pJXxHkyYimFJmrnrLtrpKubKXue1
J/FHVvTG7tDdvG3YXkkLX6FbpmmP3p8e3viW7K2vsI6pSWw9gKEq2aVNG+L9
8EQ9/OFELtejpppMIsIJNZJhsrjrl/51UP7PQQt2urloDwPQADmiTlFCGSwb
DrCXAVm67mGZ1QvSzqxSy2aKNsRqMDlNXbTME/+WZ38RBJPH2oiv7IAt1P6g
vLuRh0q9eOF48r73WiLjNITxz3GuoWngjPVMwXpo9Voj88V+xgJFrrHg2yXl
dO92tOCvhsX8DO/qvT1Rg63UIKD8k0H5hERYCOHp4jgDj77TE6Zv9mPvi34P
sN1Vpwd+dFJgwx0fgahoM8Ykidae1CmJI4sEaGKBIg9BXGsP9Hw7orflLmrH
LVNfzGc7r+33wz/SBHt0ssmVui8HTFL0vcnzF6VzaWNFgeoMs8F13VHI/9SI
fsucY2f8uPmRPb7GWy7OWJSZCEoH8rLI0a3h/xs4Ph4K1iIa7NeDCiM7ATDd
hxEfzkNnb5TK/JubKIcOCkhGBs2mDzJhcx68rWYFrurx9y7rQSMHZFbMWpNn
KE9znpDnn2Qbp467FFEQf1im5CwSThtyp5hVvkGf+MEhj56se4Wb/FiKj3zw
jTsSK9xUDoADzY0IGmo+B6X9bLghEBkYQcWeetJoWQnFTfOkpnBCWp/6hR3A
gB4EPg1k+uKF9S4AdtDIWLb9keCPbwdErPUjcek4hsuyMfwIWyhm8RFu5H1K
TOYkHYHcjjawIObfAmVJrUZlj9JQ+poyW3qBBs105rvf+x8o4mRD6rBQYlsM
D27XAL4Lvn9TXy1m/Tf0haTrd+qS+3sURGKW+BzP45ghz8gYiEBNNLxNznyj
KpOqMAv1miypqflEn4l+Q3fu97U0SRiQhvdpZ74LgmP8H1nzIaMgr3OIg+Na
CaxGIH6LBj4C0AjPbc+WBm+klVDIxa4hCv9bfK1JzPXVgtJD/J9w0n/wayNy
3K+qmxE8SV/m3n9FXtw13g/14/Rx21KsGSxzH0w01OZiO0YaSLPe5zWAgDVh
2V3Viu7R1jgqOIiRx5UVqzDSQ4Tde2h3E79Ou09qOtjCyCqKer0BdacpGBpz
BOfXWnC/9OJbWy7NzvRU1zCZ9IBbCKxzx8R+/RUrKHci0REWIwsoaVfEim6c
fij9jAkyA8koN5O/38zQ6SZywaMg7KaMimDTahfD5qTj20SXdYKNWB1P0Gte
V60EDGR9ORp9LdAqiTW7eF7CNudtg/LDkrU3IFBNtHbHH9Cyr1rFJlMigXef
Vofb2aOYCQbsM9IF0jjDUKY+OHY85ad1TaH6mC5vu0fWSqX83F2qPsSprX3W
BEjEHfWkG73Xdp5kxCCUz0zBu6fvifs0zn7vBlwvJ+RrsNlH49CemmrgikVs
zW8NzqrQlGFrd0BKRlRBQY8Ke5pnjdhcw7Ik7UiMq2Of4E3IE+H1QxlWd/Fm
CYIqiobU6pGWa/qyOU3MPZJd292MVsTsAgSXgjAIz7HoIL2fGrtgBNhz3vXG
vcmkRGoxz6ufdmvtlGD/sLxZusg1q/36FuMNIRmaHyYN9LFzaYxKIcMszfPa
SX52nl+ycYZs9EIUsIZjK43QtR+zJSp+UVGmfV/DlQJqZsC6JY828rmi1q8F
3HSbzu1CoMVXF8TQoxApQ8JII5809ia6iqSgr2tAE5ltpOvrlV4mIgib6elY
2JJvycX9YwUGyk+L6Ze4PNYZ7KvU+rrZJZSeDHgaxJzMbRkLNE4lR6qUz8PU
wULVOcE/GMaCLLhpogRfsOV6fMP1nQV9KCO7ARAjeZnNoc36ecBhR4iGOpUq
KImvZaZxT/PpM+f0y0tRjFo7CAqxKjYelqQoSnE5oHogDm5WvN2/uTzxqojt
15hdRKoLSi8awzySUOVdAFvlBaGBJ6f6IR0oNSFJDBIQDyNry0YUl5xtaR8Y
0HtTdMxz7SDDyuPIsPpbeGkLktFxhylQxiUpqAMJ6RyOO7wNqmsFJItF8Bm9
zzlkDHM9UMptFiYWpgjXoIJ+XXW/HAqbxfKQVnvJ44sI+2/9QRYk2cKRGN0j
gdDvK2JLi2BXgBa+F0dQrQU6VMRr3cxwomFowdvNsiT5eUcfIjKLGElEo13k
RLMZ88vfK1RSCzjzxQAL2NDjYNsNeahmwTRxajom7i+U7dO2nHKRrSSV+0KN
wGLxOML7/JeP9N8G/bEYO8thrQljyOJ0866qPJIyO46Gaa/dTIm1i2sywcHk
cilbPDNE18S33PrcRb4l3GakEoaz8vXyHChjyMKF+aaHkPT4AFP7hw0jLJ7D
QpZncKlbAEP/RIyZAnCQPp5jQYEJ/x8SUe3dsPMUMoukf3XrlW+kCBoUv5Zt
Zip0PMgFoTWm9pokgg2V4j7vm1biNA6vVmf4Tj4jpCZOJn0KX8W7aQwle6er
gj7WDtKt8u09NTRBhtEgSWLwKJJuRMzlS13yZmvkfVAxvA0c8/LJLXfADP+E
UCMopYi75AxacsSFc2p8jsV3kPH9wMLjNWFBLfPMBPDgaV4w6gED63r9zBu8
uaaPAI10JEkpMGhopZbEwmfQ+lZbLt/Ujj64bogYMtUp31tkyEtvKj7PRmZs
ihs1NtDgnsjoPERm+mH5jLqAe+PNJiZn+1mVR/Dp/evzjcaLanFTGr4Aah0u
I/D/FICGUWHcOLBJJ0ni5c8xIiJsq0ZF5iK4STom15co50iBzEKWlawpfhDs
ESS//K5fnh7LJebNj/KBEtIfnTucYxIDhw1gE2TBlAxdL5NTGkTeHjpJsWz+
Ua6+buS10eRyVPMxg9LCkRSdS+hJr6zDAa36MMKGOxFO2pMe8MUwExMhHgO+
ylQHxsemsjw1j4A9/3dQ3Y+tPSQcshAlw4oCfXHhDquxMlJDBO+Q6zchR6tg
hnGLBl2lqDokFLDgi7THZwdw36bZNz2jZR8kEYbl+7ZNKl1WVFfRy5v3k1Vo
3/sBLNozbkXTGMarjL4slLl/UFqYengu3G3A9A7uBxSzEmPmCVINSTNCRFdN
AqcS6bvDzsdmsXNG0d/EnoFn9txa14m+/lkPiD9O8teVGlVz7N+QAVz35UAz
QwMxGKcAnZdSPCzTmJJEP11FbuSaldLVV6PEXfhtCcfo4hZtpAAZYdRRuKMQ
plIN7ybX0/oAnM8QNRI+glNXH0h8ds9rFLqSFyHgNoA2NgsHA7LbqlR9nMQ9
qpxm5z8+6bOGqZg+6dNp81ZA5itoOaRG4IgGMYT7SvjQbpCbLFmQkpntiwli
FMuQEwoQiA1GR1chw4BVCBmx2zmN3ScE3BrrOSnKbwc1nHCRvfc2H+8rKW/k
iz1Jz6PdAoAgTVmMoxQWdvzYryxRFkkMslfHcVZ5DenswFrc5eWkT8uT+TGT
aKPhb9lOyYYt70FEZ3ocBLBJL/R5zA60qdkPSATLwBCDklnKBikmrLIOj2ud
jdSkAr7p1jeRCtzH3RRleQ++dW4YOk13BgneRpQmzvo+rY6STeXnV6zkbSCU
lcc4Z6tIc/xBePwq/6wiYKvnvG/HL16VI3pSo+/ylwA78s+X0JPHm2zDwG6f
nkcnT+7V7k4gd59fA0XdZTkj0vwooBOEtPdAUTN9raQP2yIKSUq7OEtj38mj
4uZwESEN9F8g72f0lyKVsjs1pDK2uyMvL1vC+0a+WpCkAeng0BuX/y0HTRk9
CZGDDVM6WgD6irHcEQnTN1b6JrjBFcybKTKCCndymQ05/rkLijXQ7si4ZZwW
uOHehxKjJ0XqHc4GSaE6s0Cr68cPtn4W3nRXkVPxqFwEY+0B/+g0Gg05R88/
He1NtkaYd33UUPKSaQ5Ubts02+7Ee+/IAnPxxLVg6imOA9UHr1Y5xhCxI3Wq
O4AuqZOKaATKCTpgAuK8ERBCxdmA0bBzfm4lTkMlc1yCCfnu/VksK0XQ/Q8f
rCzAVy5lePPcDlL6QFrvNDXxzUM6uuiuNbRlPPig1G6USc4gTOxZlWt+Ubq4
YbmfIQRHNo1si3xrKiKQNz6js5ohcAjA2LG2IHOWYgp8JdtZjZtcxvsHxQhc
jabkRj9h4fIJs5bpn0MCpVvyt1StsxyAHL3eV25X4KQY9BwL8Cdo/H7GUrhz
MHN6Sa5YUOjGko20RcXrPMmrpjLKE8c3YLfgLEHXREXIoUiHsChu1/6hJ78u
rS5v/OzeprTWOgPVMPV/EzR4WfHwvV0d7ZlG38UafLQdiOd1GQTEIOY5u1En
uNqQibEY0y+xFdCGAtOlxumQwPUoDXhBOJ4XeTKglJiS7Ottg0RrWgWUEj8h
16AUIsHK6UZRHgCBizVSbIP296L6sJ9TTVSg0Dw1C9Uh75/NG5LpGmkiHM08
312uppKel5U4rODGGRlHR/lD4VuVfEqs3/Y2j9/pC8eAyyHByFgxTb5Q4aaY
EqBpIZU2HtBud/Qtss4FVSfIA9ODoUoWVEhDML5YWCDez+K4bPCjZvCAz6c1
SkGhVgS/Lx7NBMO3xB99NnJwfBXahswvNICEw5TMV2y0lubwYAgosW5PkkR6
7pTYkc3BDiUYwiEJaPV7AOUlEyD9P/JFIx3Tvzgud+ezGEMlklqpy+1wFDQB
RBEr3OjY2wFrTCL+X7TfkDAcpWL06tAd9jWX3+iyCYKcCJKbsLz1xtW9BfOd
vPnrSMlxw+wVcaADfINJq9GoqNcc+3nZEoaidLU8fIAiJXiNsiIdJUnnKZM0
cg2Hy8IydBXGaEqnEGKxDsNsDd7dZD39Xsqg9NtGu3Ve4dnEan7c51Rfc0Mf
fAJWtw0kdLtt0DXMnODudnSQ7GJRoSweJAiKPDPtaidxexq0HBcb1kNvzrJi
K/vz8Te1d0nD8uxT5XwgAh/fNHVicJT1EvP2EPES5c9hNMUrG9jcj/pr0HQ5
s8cTeDTl91JE3cp+NemQgKsjoq1Ryx+ajS33gycWBWsXdXHbb5Yl1W5s/PZY
ds6FwAqm+3ixn2/h/YF/Gsyter4FkROHRdFRQce863f6mxtrK0UhwytaM1h9
hTFWBFGt+qZQKwZ6VOMidKRXcvuG4WiBfJ+CM/FFAR9jyh5XrH5tlHOMg/QS
pasY408t6WTyPwrtoSQDSW+NLXyhdwGtPLfPg1BZ+1NeHN6N0G/V3CKtHTWd
5ozmFOqqP2nCpwYyKNld0yNdIjlSKvxPt91EXeW2FZwtMfms4POWEApwSzZJ
fXo5Re0EHwCeO1GCuXjh1++UOAUfmkb9t1tg5cIVASsCsrBIbZM2sqfcIhUP
SsSUghuG7899JmR5dDEhQ30TpqSknNXKZK+yZUoCASCDBTkPiVOystWUgRjw
LaBAxZcp8wu1GMBfEAWhT9eRikzyc2Oa1ZwZQQo4hZ3m0AX+ehlAXaudCBcb
r8qsQTlVcEeJ4HSkJC+FykPRRR4nNTmtqVbLMaq+XkxmatOMqQ6ePq3Bgne7
u7lTOXOL3VzsM09xEmxG+58rnY/Vxeq2DF63U70qnhBiAl92Ac+lJ8kj/NnK
gOwLspdW4XawWpbSzQ4ppiaNim5hnjqeYsBOxZBxoFI64h+2f/42RN4V+POm
ghORKwepGMZgpFR9emlGSygnx05qyGiBcIOSjcoiOut9Hqtb+UBi/OsnK57v
URxAhkFr/O7meo0AWLdA1Rvdh9WkQt+prJRY2BAxwzngdxAN6ByP+4cLEBef
GaCYZhzSp5Bro5s2QFlpMuqGMfjSgS82R1zq/r69qp54kPkoqVglRb97k5KO
ZxqnzMjQsjVl0xKDsuxCbA6OwFDEXYptQ2XhuR3tzbwtfTk8VWbP9oh2MuvP
9RJtmCj3mYLfZZdex6etDhuKYJu67HYsVrAB7iKkYwH9wBBUqP77qyWQ33qw
vkPt8mbBy77Qr8LP4ez0es68RlW3dMSaPj7sFf5kmkLoo0pHSV5bT9E3x76H
FCJCt+1rJssmjwA+WoDVP7N5qr0YkWVXCpsi7ZC3tsHw68vdtFloGF08l4Gr
66Mzl7b/wwwRYo+3MIXSPJuTiQCFUEoequD/4cpUWdstFmXQzYgXJNz5K787
acgmORzg5S7atSHEBbutUSjmUzhaZKomOMH76vnSakKLdpXJsneGkvt8umGT
hOrCIHYmIJ52Ago+ggZY8+Worujb3xsnrEjKrUF3YjCbP4cr/JpjZRiOyXpu
wMR2fDnHJMSFAPQlEG3os3wpa/YyRByhcT6ygjqbImr51YidOoKCVE2hlKNk
VVfVhEIv0sXnaHYy3ZzDY4j1D9jaY8+BZ301YrdQVZ7/gMQYdNoIpr4xv1mf
u23FlGE4zjpcSm+9TkQouXmmPK8vCB5VUSMDfnxGOQP2vtrzzk828JhlbFL4
8lEmSEMQ5ATCG7mR6QPP2NXsVkd6bk5heTIxqQY8OQknw7JO/OjJowCGWmIC
Aw/cdB6eQNvXms7fTttItpsugGJbbXQNk1YH5EUsrY4p0Wz8aPnGlj0oUS+9
pSMidcN32LQ0cb3o0v4ssfLFQwvzIqrMmmpEMt1A0ezaSkxV1KQjZ3zr40u7
labTeWO+zu7DgUq3TgiWeS5LIWlGX/Og30evT3FwJd+lintD4npTklUYga4X
cVNcjlSqoLGYOYfI5cCrBP2z2RpOEC2YwWmC7HbdxF9AvMH6KYXo01LBV3DR
6sALYSp8Nixrj44kzXzIrCjelHKPZ8uz2BT86Hi5oCIjaSgTt2Ye4G+brpHB
Hq6QY2PrriRsRRij9AcYzaMX73oARRwPBy5m10WLtuwdxqfnZ6B4jmkslKJa
eUE/V/G0LIFm7fUvm1xjW7UciC0RmBveWlWbh/4LelbibiHJ97Ci4mSRLhBG
ShA1M1loCDbx7lUEn+itT090a2V6AIAMOWU72SFgmXUhS9d8eBazSTB58n7U
Mi6q88MPMn0OvEs4QMpLfRoDVRnG1lPWz08ILgrze9hPeyNSp5mJeZLRYPZ6
Ztj8UvWlrqYkwEVBY5KpRwN4ekW3YVpjpCq/GUp4V8IIgZNDVh0pfs2hEtFu
2HpihYdVuSy6Kp79cbMoAGYDW4I32vvkXNFS8LXW51TnXLJodAjS852AerAr
0JeM6tSTGUu0njHVkMR4g/um0NZCrhU+jwksf3VtbEqw40sDd+0i2+0DKyrH
8GSW2EKFS3qzlpMAs6bMpSr7KEhezUBW4SAFOfuOe40RMeoll2HXOeUeWxBU
IJyN0aQeW47tZXoJvuc3jDU88CCN4BBXbggxwavP6GiSHU4EkWccm80wB9SM
4LcC+kezlYwlSrgtSWpmiaIQCZR6K9ePKeoDoo/9A2iQKfqGO1Zk0kUtzEx3
XYWxofvryfEU8fBr5LYorMG/zH4BjcP5EPM7DFzyQL1OXinPID7Izcns8UnU
k1oebpFABLGzDQpyuIatnBoD8udYaLOMQpbTqn+xWj7Z7AuCjvQoBGrEfffj
LQWE7il/SK02jkU2hFhDDNYW3swdHDTwHLhBWDj3n4hZMOo9IJ5W0cMj4n5U
aPGbCHmZA12XeutUi3pn08DaxCbKsrllP4mucSRUQw8Dn3+mdRd1ika58Kto
uhu/TM9X8qvv2tzmozPqrM0SsaLu1NQHgpeG6E712swXvmzDmUsqgjeSB6lk
bjZiYGBtDHyidTg9gK3wIGUPskjx+vSjru/iyfI7n6dryCqoUAlA75bsX7XW
AnOvy4U3uz8b2VUqgIa/TRCrRC68HkiP6sR8BGkOWtw8x9htm1XhCuTv90Ag
tZUOPvolm1ow0b2HIYnvBAXYyGPsahirZOh6vSz4SMSyYCRz1RapECR8seW/
XCmxB/XmWg2XNXKoH3cYvgrz+IJ98GMJSE49ezoWXPAqouTJ1xPqGxCoQjj8
LOEKebRjyhcNZHRsj8oZVGskAfpzcDEZH+aWZl9umbVMCyvDtva8/PdbaNCK
MMmf5m+K0a4mtD/8PI7tW+tRUrCI22X88fwThkNZtVKmw9fbKCpMhRjlWIuG
AgkcCBf3a0PDws8w1xQU5okCBS1jkKEKmWgcG18qPIEByRaQ24Mm2vPDO9LE
aMeGxgRTieTr6McaWvrX0fKdvqzH5ogCgEV8NmrSK6UbOJxOvxqzj79mBINh
OkDJNLt8RTbG/H9xE8gh3APBt4D+F5AfnobL1ElZZVwg8VoSO0oVanMsHP27
e5kR5GOORxNj8PKy+zZ6imb2bSWDWkYmM1Hf9JLsYaIB07KNvX7A3CPzeX2y
ZGEqHUExfxaLdizvURRsdQQdpbZ3pLt7pW18BBMkMXPOTVvNP8clyJsgNM23
oGWq1S5DzY4NKx5LtaBPhiIhypKkmOUhWzXfXPdvF/QkD8XcoihcLxvgaIA4
QK3aj4q9BV1YO4NMV2xm3b3FqqWaaefNPbQRzSCHTHVGRx1RpRPhzRo0aq3n
sx+TTXOSFMEh21ogiGgW9veDuXk1Ftxi1isfxA3E5WVw6zrbl9Cq+4goxrF3
xjLN4eLSugnekULdiJCj3Cct2q4z7wvyKg75MHpOIuVRPFtvo7Jv0jzdx70h
PoWkkfXLXNA1QfFMGBCaqup38gxTeRGTMGdMJxwPi2BH/NZDzRf5oEUJKr7J
sNEnyLrAJgwcn9sxUAI+kQ8KzU4Xdkwedq1/6p1YeU1Qa/QAkEafQtH+MjyP
j+P8deiQNFzA7r+APGYyci/vFcltHuWAHzI9+hoIbs3Zzj0WLeZzMfJe40L4
1J/J7jtrPittCsdmx6Jv+pLhw1DyScHFXcuulWVCyFZPx7iUOeceRAAgknnb
GSA1sCUr4obdLeNpD9yrrgPnhO0mHRdkAEl6pkJ6eBaWSnQheEioG/oYaZZZ
SVKfqwrZlXEoBmA1eSuzSa8dBuV9YxfqqK40naTx6x22sHngcuOZ4sWRyXfD
BZ9RF2LYlrqqmnnaGUAGfM9CEUeP9j2PK7Kz3AxV/ZGzcWsbxEMRcbXQYlDW
MMOstbilSNxXSMVYWozhF36F9XoEI9MI6hmG6qPR9FOUP5ZA8IY6arHFjzBj
S4GoJ1u7I8WoGMybwQqaAGJLaaRGLsVdQgFk0JFfCFOd7IyJhtOywnR2awNW
wgdvXkYQmDo5D793MU42xPFdT3M2OnqdvrSRlzkowXHfbt5GoWLtQ5HF+gss
dQajOiN8L48Z0pA3u1hsI65bubBw+U4J3lWR3j/V8Jz42NQ0nJQBQGAEf5rg
XG45VvdpPKPOg0YzFTesrsY4wR4tArjmC5ULllrMw7S0e4h1EiFbC6WB0I1F
pMTdzFMS7+9sCrG96azTt5uyyFqZ/Vf5rLlkCyPgHrmbqp9IXcHE2X1rwz0T
WEu62nZmB3I2HPH2Lr1Kv9OUa64hEdVG3FVhi1dw5Z/U1MAr4TDr5IVUM1wE
7SDYFf3lth/tGkwULxdd920QapGkH6+b1iJkexr3haxW3zMWpESG8ieVOyHs
ouOyP8ZtGWIe75fGYZ+4coQ3gsqlrUbre59U3TAQgGzv1Yp6ayhyUsYiXlgy
Ys63+VSlYR9Ea+SpKrCTJEmo806wqZbbqYkcqJdI8yYZgDlz0Mlp14AmOdDI
ky6ZOimi8Gek8Pp/4w6EcCe8ZS3J64kfxhffArhuAHx/u4PDKCgv9LMydRZz
b/UKVolRiLqxV1uIZFox0rGarwOUyYtRffXoBnSA1tZjR6aF2iaZZi6yMr35
zfgVJrIBItGDob0bEmsMExLVXgGEXPrdvJ3Z7SkG3CnADV2zLlhQFMBzJLgW
czm6QX2qRJ1uk4BLvg8PnSEvMNOpRY/mXWx/shNQXVJ6rQ/v6ILxN5sTLbbH
EslseInYPNvVzvWtLdxRs0TtgKKNy/pv6Q64Q7VOCU0bcNfi/pOLP+XOckYg
fj64j0qz4PTtmoHAEFlv4vuhVETWDU2LRsyNPZmlmj4ela2Z14KWS+/grnX/
n2WwXt9nbetyMfvTAq9RP/SV0keBdadnw9gBnJhN9r0ApYh8qtL6VybvUdT9
UIRbHnY4ovNN+ipbdcvNslIMIOq0IU9R1Rf8eaW0kzjabZF+fK4F3RkcP9l8
5KLQGYljCXqjOCC6kAU/h1YgPb03oXxIuXjBmsYtoOkSvUkC97oyP7KVvbD5
Wq/enhGBr7Bnp3ZnOjCwJA5wEcFPx2jNO+HanAV8F+TyA4MQOPn4MficvCJx
13SdUohix6spNhFSltWcMx8G0FK4EW7ksYB4h0kfRo/YMIHcNelBTWK8DAzC
nYdC2yVebhtxGcy047AHTQdkI6TlALXvaVx5mzRimRg2jYdhW/cvdKpcopNd
H+od46Ul0M4YWbtuVm9eBIeJ3qm0UuDIN/N3FJ7lPqgcOXWZCT/dC+hL7vjl
k2/vxA1lwP16mS3fqfhhj5hHR27Qaqf6DPD24tu7+D6PM2tI+jMZX/Dz6yux
SENfiVabUgHGcjFlyvrdG5iHiP2U8EDzG2ueAhNBVJPYQm/DL/sFKGx8aBS0
gkXLzVWb3Xr4mkbJiQl0xtFJmyuU2/KDOAuuUMicwXYkanl6sukpm+n1d+O/
d4jyfevO1rc3fFB7J+ZkYdpLAaB2BzaqmTti7vjrabKvbXhkv6uAIuoNsSDe
eA2RqTj5IpiBJTBV2IOSjU9LnS+suGPpbXKDPpjGZc6SU1193PGdw6yG1tNx
VAdbZGE2fPSR5hAScjDU94LlJepDRWgAmgqLI69eGmQVDkrWH+eSUcYvn1/A
Su9qjMKShFX51Hip2wySxlCryyAxaBBmTQxQLuB8HOGEdrz8p8Z4wVopvw5D
pDilMoPzFkIk7ldwBJObvc2JwhCLT0OMHQDTCmZEptW6Umk5H6kyeHVk6oPf
QkCwZKhFelYf+qo/zyIvw4juylG8DzlY0NWkcicTg3e+Q5KDju03MftJ6ATZ
u0oiXKHaXZ9XWcoN5DPkE+4ZI6SkMK7xX7l3D+G8GgE96lFIS/yXiM4o0JYX
JYQ4NwRZm41ixZuDYD4ikmSzazHNeLUtE5kZLPt1aoNdkwnQ2YRXfXV0+O79
rsgbW1D7skD6qVQtpZLryNQL8jLycXcqTxIXavPu10zimYuH20kZM7nXtO6v
xpyOcWWA3j8oGUapyFbpreomS0Mk3tWflI1WrDoN8z4fBnHRKwnV+PtsvvPN
EQb2ULWE7u0JmnlXdwfSGI1bsGd5r08xt8G9LBS2gCQlMZmt+bLpeKqn1tOM
WvW/KFfkk2ecrK/TnjWbozeV3xDyHiCEJaje45ON9JU1GyPGyFnJ1cjL5Vmd
+jwECUcOgGNKW9RRHgTdPQ1u9+QIcZdpvIDMM7hnBaFL2Uwumtub6/kzoNVL
E1PpQXPl6oTZUMNT5p1ydK9/ZLFYpX1Y8gYo2yB4UNnCNkhVg7BkeffnaCpk
+HqTmy7HklPLczHK97HKTooWM6bGGriB5Gzh8GN3E8+5Yrng+h6RIjdNuerO
GuOtEBOb0umvb2g5k3x3qQEhdPw9TpWotArimZU/kZAsaGBQzxiCph4y6cay
Nec7ibKI2mA1sK1phL5+6uPkJXIUV5GOyZXavbH8LwHB8xZQXpAp75SpETTb
VnuJiFOuogkAmqZ+eh2/622iJ3xWwrVjy7GmInf3XiowA3Uf4hWxYel6nR6k
u3LJPcLzYA6WHFk4KuyrmRg+1124ieIfjP2EpEi05b6u7JnuVjpiOWyMpw0r
dt+d0WaOch//RUpj23fyuGWBSVFz2vwR8460m1BCPiXKxq4zxZOc+oK6PfsU
BcJd6PEAxpjgNJN/WJxeTET8bjHC6zj4PuHEk5AokBLrXSoVbQurY6p2kBMx
X3AfpPseToBQHxi/8y2886uNsM3aUEhItWek7vurs96ChoP1rROIfkYG73fh
kIcCgZPoWUH3+i9MXV+53JzUlT0n3PR3zZWWUAhHf34jNto4WEeY8WJEragO
+SqJlIaLGpyFpUxHQjiZVwvDA8crzt+TgFVXhF+0OtihJFS9wjFFBDiFefFl
1HRcm8Dzm3UgrCtWCoPin8Yih3/qb3oG6uM7gZhma9Rb7kvqqxI3aSWZMg8W
pKopR0DkOjqPwZLE7zbm4TEaesghEZzNJv3QlXXVsDMqihm5yfElqJFO7572
rQWGWSzCGH4i9HiE1Db6W+J7U6RzeyNjIy4cCOfwYG4maaBf/R+KLjm67fU2
Yx0b/k5X9HfVxkY6y+B5xq8V3WZth6QHuqKi+1QUHoThj7/J828WBAB9kBOH
V5PyD+sGmAT5Jgr5NKS69OY/Ky3ZQWX8f1N3wiAe4tuCOsdbMMYAuuXxPJ33
K9IX7aC2nLVj4/HHx/lnzTtyDN+I6sS0tXc0I7mdsCGvC0CK44FAdx0Jl2aZ
ypVfA7Gy3oLr7d261tfHHLGLlA6xgRbf+amUtJf8amsWTTzOePf2NCCLeJ9n
lOb1EtUwYlFz38kUMbn8dYcTXc+PiKk1f0tDYjMGTFi6wv+CZSejNMZUxBtE
c/cMPoijTvTCcuIEnd/A+1iTSENrz3xxu15YiD02On7IBc1Ul7GocRmQCScq
D412u4jzRCbJgytrkBuIO86OG0HlkLWBqTKAdom69MMjSIZi+vebTmjC8Owh
VSlqcDLLn2eQZogxmtvy+B7EO9idVdeLwuvUuhl++8qmrmBy9gkZ0cCoRUw8
4in4HwSSIF1yByWBm4u+CUbh7XXMG46VMov2QXozuSD3T8ilxgvkVVfn7Q1z
TCDVpp/K4Uz9tsX4n2vFWHG1STRM0oR/muC2jYvLJ+0e0LSg5FdO1M4HsYqP
vUWVmh4HprIeVdex9io5wPfYUEsgdbiIntLB4RZbtBdye60MNEnJ4r6S8xg4
jvwdAC54tTIxVVhnFMgSl+WomM9dmG/IQOHXy8pZgzarUB0WTTIBqHoH5HYD
rbesvLWAV4cx+V/qxvQ2T+zyyPFJjCJIiRklAdjJghzD3fY6bJUP9vpqCTEK
bkjlV/Z2LjRo2TSb/GCjP9Yzh6uAlTVdj1jzYm8tIONwq/d7jgkELsIcHdGG
rWQn0nO46OSMIr0WqEYm1B5rJ8peY6vYv0xTkBPWqFgW6QZwbqQVyL1ZGGGA
LkfMjM+9SORrIH2F+GwIvG203hL+3iRJQZNVDT7RQr20+IW160kCvptgwFPQ
57B9YrqbK+IksbbQ2IWzjbXicozRJpK96nrR1QA6Bx2OniT5R+P3lw6xwKWB
XNxm8zjBN3Qb/qNdkoRCAF/8W1u8RrwFE+T4Uvs5hs813GncHwlnSP68BkFa
k7TNkMmgTpoYZULuAOanYMtQb+Gpy7Uy181Umf5KCvElILndjqA/Cz6YtrkQ
QYFAMX7l1PqRmhUp1epFLIja+IkY4Uz1V3uSEaIRo0qntS1JqBcRrPbtMRk6
Q5GtZhQU9cWuvppn/lRVszCv/lC7d2ZONuG5z57e4edcqR6md/K8tZKbKPJG
ZkWZ8oyepbpn+qX74zh2HWbm3+86WkJBPbXvDHmKvk0f7l2kC43JlmgVk+C7
lH+aPn4FUj5PG9pWB2/xVGjuVJH/2AwrbmpLjyO7epNiGE6T9XRH5+t+Uy0w
BC6avhL03dImsPcFCotNxdMiTw+9bUm6jPbWJGsltRbX+bvQHA+iOTTbNMlr
rJS6i/wzxZVoV8TxFnudKv4vSFliDupY0TuxS8m6/S/jSQfjoUQlUq8rp6BR
V5pWq/9pVarZjZipL7oX/ZBaXqTepYwq6vKdb3SKYlPdyoqbIGcesaRLbxR+
TCPP4gr+Ve7EqaeBnM9IFKRFwrRlLhyBKNJwTPr6MvPDT95xzAIkLcM9j2Tu
Fa8FcgtAwuVMzE5jRZBST+bV/JKlQljvczR4OAbSwWHcYaPk+atu1+pHEDRV
wTgT/vVT9RMpY81uiMhZkz59NuaBfufxIyMsVAzXvHnDe3LUaIXLdXz95si7
C05iXwZsP4VbpmOszTa8Cxa0awo0rMFZ5yJvdzHxZ77MhmJsmmD7mDnOIW8W
xCAqb3Pq7ZhyWKp9ZP3d80rL/sVLq5by/9t+Amin3XMpnO9APKsD3a3lpEJd
8SlxyQ77N7l9SOU1As9tcDD6WNd5VGIMylPRgXJnfXQuD0G3f5UWDzZuvIf7
dV7zUK5W1KtIYsk9D2su59nI5C0GD0p6P+GwY6u/nLkOew3IAHH2UevqFHuf
Awx08gQhM5b2vlJoCPYyOTRXKJsujduPcZbLUk8A6vcfClaz6UffNtDtkydH
v5f24a8UgBX+nn9nBGkCo1EKdBglKd2PpDEaX6xcoFFHUk9qyhbvcLZPEHoO
EVHK1h2o8yciODGnZWG1X3YavQJ1J2qDU3JsB5LEqoHhUNZKh1gFnIgRoyoI
1MxLNF5TCKtEHpVF2vJ3wpm/vc2ayT/LkFDygDKo7dUsRB/CXuBR+WYH0R/R
CcKcDd8Rop2PhjsNvXigsPVr0gmJa/jfe+V31GuTkiIpZupp/ViTSsOPUl8g
FW9HvGz/9gYvQc8j5JoBP1BewiZ1N2HVYAE6pCpJfUgrj/ycyOefOJRe4hVo
xuauJ7F7bKYEm9ifkkf8hEOVisrTEkzNzSdLcd1MhSgOq3F1jEd4Z12jXuGi
6JdSeo6p1KDTNDPzee/5GDyFUFPbQSrxu35ZAIeGoyf6ZglR5HJZgxua4k6S
BiKL0ZLwVY1SLxfKB/nhSNjekdgIyOgBoL/POQ/dprsPDVt6VkJqAFAQuAU2
+9aFdJAkDnxf0JCtnuqZJTXAWvkpO3LrxaDi8SABNLj0GhdXDNTocldxHT+n
KbZ+phN2thH7xZZdS6JSx4NAzg/1eUpdY3OB+0l5jxMd7JfdUe0nyNTp9903
D5UMmCnMYASjG3ke9sQeE27D7v29zhBvwZDTk4rgdAep2br4GFtiIxEv8Zeb
O2Pe0QjoaOxj9QwvEyvDNgEGjS1cL1PfaQtBQ1acKX+EvSuMSpiXqmIT/agP
X5fdCgVoJrCY1XKWsPw4lauC4JFUz+kkX4M57AU6r+TQ2CV8UM3VpHb/YwP2
sjXxlcgsnKX05e2x76ISGPOkWVMith3J6MMTRI/76pBCxTMkOKgKt3A0411b
94CQyMuV0LPWIBc8hTTju+Ni78tUCuKiV1NauqONGxMTjU5jkeVf8oWiWYZ3
XadRPPqRTAa6e2OIgS/UbMxW2rz/rTvkO1qVVeQqqee8sU+IVAVT/mho38v/
/buGF3T8wxT/IzqoYxqDVAF9HL1M1H1fJG8r1ici3BtDFNts95CBAVb8opP9
eWVLFoxnauizVlkeNPeNBtd0ZvhgKuE2VTJjvw/uxPb8KMjGfmUoYcCoK46Z
XCFnnWV5wVTv0hhHkQTgC08cFuAKQYGF6fTGJnf/jWFEasl3wC1VJsAYf+1S
HrJZZT26qBXypGXdlwdx8pUlqz37sztYarAjVLtITB1bhZKC8NY9A9VkIVrG
cLMZ/rejTUzkeKzQWSWaZ8c5qO5B0CLzyZRFA42jQXBLkfeYHu8A8XY2EyeM
qABrTSoxctQsEsGDJ2ATJ9vQnAymHQ7HijEH2DlOUe0z605ykYyM1wGbFW5N
BZsJXQmOtN0olyBCy2xTjVXjf/XivddYPu1dkaidHnTq2IZxrD9VNckQJncv
gx+YMGcFwOWUI6DtXmEOP45Hk3O9lvwHVoI5Qh45QZQJ1mLBjTeAGHxKGOSa
0opwu55ZCD+vTg1zZ98YeNEF2Dnyo1UWb1Zn6h81vVfqR6ZCbdmLBIMtpdmC
VdvZ6oYqccTI1V7AsyswQJtYEkdRhCMQBBgPsVrKkjj6I7LB63P/qGQ0DtLh
XYYYYYj+yaqXOB1QH8ouwm7w27wKyAVRDLL1JHHWjL1wBKL3fhO32pmMjjVb
LdK5wqHadRIPDDMyo/VU7EntrlNSYViZjosOdIAOkL1DoSqdj/Q4B5WaL3Il
nytl88eVWwSLwTQL/Yd8g7+10UEM1EYt5PPEFMMfseOFb0uWe1zH122X7ceK
w3IohbAm0EOe6cRKXNasa4qMkF7/Eg7wJeChiu6Cg/FRq3SzBXwC5yyMA8vK
O6YLaRTEt6sprzdVCyUnBXwzcWtye7LLCG3xzg7o+fbqC2WRow1xUdlYrNuI
/NLouMzbKHAZ618deerFCbeKywsDt/ny88g36a13stTNmOr+SoLzR03z3ZNC
5+MSEFWBOCDH+EF+EbrZUXurynQazs3A6FMxl0d0RgQI7ASo1cQPSYYOtI8t
R6kAezcxq124/NxuwN1dG08HMxc7K7yjZY50k0I9t9s3AKER9cnwI0FJSxo2
z45iXy24Qths+6DsIuxjLBxs0rv2GwFgnPk27/5vOggd0mw+JauHwJFeTaHJ
IPUWTFrqa4YccScphzIw0netoMHLnq6/bpXDm5WYcJXOFEnXMbrK52P7oGWq
YduRYfqzf0KS4yMaTab38wpSMvfRcc3l61e/FCcWj8gPFwQenA9Ot/flV95+
gye5iR68Uh1ZX+DnK6arfzr33yJqHrYMLdeSV4jKG0gEesbjKM85MZTo1vdc
xus3G6Ywtyp7zp0/Yg6kCmUIi4577bUZIyOm4UPC3LcBBf/6YQ72sURh2Uoc
0687Fv1ddeH9/IlgRbMSK5cpKm62taqpZjlWTjMyo6PRriAoqVmlb+Xdq49q
9tj50XjRKezJKNWnUjRaGG95JNLdTxxCV6cNfhPHmfdKYsHig/Rd/aOONfpQ
TqvWtiTSqHBeUxBnaVAtQwqgCQD5i0BeP+0/7/f4Jf41XsQvaC5CDQFF1oYG
qJ0CCeT5vZtUWu+b1598uEoosY9qgFlomlIzYn3kVvXjIVvWRZOgu1mQmqJs
KLhCpRnhvq2ElJDkkCOhniueSjYoRe9S8zvEAtp0iMGmg15rHSXsFhPmv+M6
RjiO+sVJsKHt4tGgRCn0sfpQa5hJ/itE9m9T2f9muInth77XOxqnxLwE3fEU
RfsSHmkJiyTSvi/gfJOWebZBCPQwhXEU6styaC4xDdAkP2MZOd7goew9TWhL
9S9+vyvqRwcL2SdO/ohMzjjdI61wBNEu1+2R6AHUklmhpSkfybn1Xi+pApGc
tpSrWJBoOHI7mc1KKkelzjH5iazUAnnmTvJZ5z7ceDz7uWfsS9WMBaPlXOpK
l935ag7aLr/My737JYOUSLZqZVHQPn++UfxcjBA4/yXEtO2/M5cDBzuFhfK5
vVyHWtGrpjUQyosVKrI3UYxG4tqvkn4/qth/SBsbQFT07mmFoVdNwUQQEDh8
3CqOKCNMCdTyX8D571BxH2avfBWAVcxXkN+lOU0jnqSGGjMKCl1Pg7okuHlr
F/Y7eCRlX6Ls4yyrmLy6eSfT832dqpG93/kr70MSBKZOKVkgINOWFB4I8ukC
SAByeNbwgyvLjbdPKAPR5JY4fFNa3bev8HFSMyz+dxM4fMjivm/Y8wCHK0hT
tsSFx82kIDRKr/qg3REmcdRsEK0LzBzngLq8YGMDFvLonr56AJJEgzHDZ4Zf
D4Em1cuJ+2nOX/sQJKjo9AXfqAs2gJZXC8cztVTs1VZkmyND6neCFMqRRXL0
E85iCR2BxnRxNDMDiCRMIwSNHSvBFXYMtnNnIfB+1MO12cNrkgzyfdiDCT5t
nTRgqGr2z1D9z8dO3VmoSO7tDf6jCcjK8jU9y2iRZxpmx097hxgdzG1OlnT1
8AN+/SUT/WiXHm94JOpG1P/ASs9H1LZLa1MWFkQ37nprczuz5r4hqbrcJwbr
ZVx2VOJNScpkjQWWhQMmrImTof9x3K/Zys90ESMb4oAhMN7i5uJyFxXOHVJF
jd2olzhxnELuqYNEpfCdFbS4+bcZl2evMnbL0lOQyV+OpMiC6ZSN23hyfzok
3fdAd1R8SeF3Ex63HjOUQSIG5UwuxiN0/vTxpFjXRuXxIVgj9CXugSLk2ca5
ncUeX/xgQrK6278SJTAoRfqAdWfNOxuDR4g+/lJlC7MuhDZWLxITsQLE9U7z
Leo9DONshRHMI50gl3DdjjBgFPxNvgIwvjWtz2xcUFdTgD7bIJmyeYg8QfOd
uCgCHZh7ytpDw5vTzTdsGYCRdxpkKz4Er/FlgeSs8y2WunS5i+ulwjd1bRoH
aS6OvCbN42b6Zi38mstdx4eVdZmx6SUdgl6ontOVAyOHj9y33FQryX/OkbKj
Km2RixLxHFzi+XHPslbAeISzD1nE1YjqlxQWh5l2f6rc1nomghkgqsS0oszl
PnlZCL7IZo5zwc239PmyjhhbDWDJRCvJ/qPEIkzVyqIjVuj3w8E6IuH6G68c
wkPpW0pU/aY8u6zdpZxnH3lfnXiAOzqa7EcD6+MR4VdFjuRY3wIU/5hTBb3t
vgL1kSxu6G1V/cTpyDQzgJBqmWpoT0QP+xP3+3taMS1wQVQpas0mFPLTEGwt
DLKCScC6XepU850fyE+GmSvKSjNFrHu0/QtXLHRzA2KlvhZIIfhkqvsq+8Zj
GOHhilxbvhGUQygSbHu+lLsBoFLeVIX+k4YIYLvIifXW9CvsE0c6Xs2NoJ9b
98tKiFljvAG3s9QqZhcayp4jLDN0Nth+6Y9BMyXVYTRRDy/pSpDWA5+G86TO
cL+KN6pC7rMxPA3SeYM57Kym0920N8NfrXF8vnBpYgYd+RhBK6sZ8pTqM+Ip
KpeLjIFKF9FEMxf+95/tLSbFPpJbyg3zslsLS+UcWT5t3a/KEe6VGpqk/3TE
dVzDz/tD2dxfjyJzgLeDIw1xX57h9oylIAPo3SAVvZ3lMjidk1M3NxJyNU+z
3qnK3/EaZ6YpkH84rwZfuwBCXBekGPfuGy/dO1ZfY+Pqc8Ar0ql/97uPlmQJ
DyXhhKqTqUmfsH7FG5UhvoJUaFYV70SQ9HcgXFwEKGlpc087DKZONUYFr5Tk
uvoskPPVFupe5Y4VBoCWEey28EGHpOXLuCNTYFiZaA6FFZVWMI/06AohTdy4
sbxRB6JjF9cTIow9BMBXtLkjF8YP1GZVhspaY4325/aeiykJ3NEqaEdLt5sc
WpuS/QNCexPzd+44bzxcupM9up1mylYR2t1jADKr6DdUuokUBDloqThRBewK
28FbXWBoeC67nV//iefvjHp0BmmjafXo1lBGm9sxomLAExdsuT9014j/Cfb9
NTHzrZy64X2RTBoqznUSdoTUZzrmtoL0a4xzmEMRdzwvlrEw3g1etzVCmXAQ
9emHaScqRUsEaM4UwpAl++lCgIXQt/zyfn5s6Ix7jsYriziO5iyXDOwKknqy
wDRNHIXjnNg8Emjv+zhJyoIpUJsH2aX+TFDvIsurGWae33nuh5hNl3lE2dm7
HvJnOJ1yusRqYbvCBeduTaXn0gzQgsHNFD2rCh+Q/nKlVgn4BFW7ZUxp0J24
stv3yxUjgZaWbYts7RjqbopK4uToa0VG/OK4F2F4CiIEba/lFN63bXSw1ndc
f8tGNNiVTOiq2bY+s1E8PjKhuYGrgAzWW5QQMLax3YEfrNdEMpOIHGEHj7VC
WdbXbTEkAfcrA5rK5U4wc2YsdQl5TsrAD306Q5Dm8myJGLD84pPa6rK91ZoJ
9LSlGohlR8FK1TsibrdKxSPonh98MH49J5YhPwbmKm8s5yM9KMLwgoF9W3ji
FsW+ToTFqbO+FHiClRYcij6lO6hxx+PExtjpj0XjLyt50hx4fs5jNuJq5g8Y
4CSz0EQ7hZ66xCSBfdLhpjmY+eBULNLR2F7vQsN9gNmRgsGdxGzbKnmNA/eK
ygncgrCnUnh6H8XSMOWZ42D0u+/A7h0LTq9yw+YKkcptrXVC5pp5PMuP1jDb
T0++AUbnxdpvcFrgHUvtIIuthyjC3gFO/Ud7Sf9vn9FHCkzxE4fJBfDOve8y
j6a4dhPM2O5neVibAh0svvnJDFRWnGFFmNgTlztE+36B24NXOstabcEEHx9r
w+uD9cxaIblBdFnXfR2OUduxJGsAzBFHIbmxXMFdBeKuwuYifbddhCHrk6SZ
F83bg9TLjW1mUnZ0se8hnR1qsfYxP7APp4jTGlsCDRTu0/4GQf3DmlCwH0Et
+DXuP/7Hwlxp1FFFjLhWAFhPxo0WqpjFUnReEA/VXgSZxagLZISt9qtnOnlj
S/ccBVxho46vAickhBwAZf1dp7R5jnQsu4kUXyTN1jkOmEiDBj0X+DPo1PIr
/1TC1+JxuiEDneOfL7cdvMmv+BK2j3aoCRT7ZoMmJNLA9vIVQ/1yYNg0ZnpV
Tb21cQj55gWsBD1M8F6/n2AbQsfr0Ag6PXnKhiLrFxtVnju/qelsNQPJMEJe
IbYbSgH0HU6N/gpd7yvBAJ+vh6m2k3fFfK6dlololumPoKhHgdJmlygmYDMM
4SreuyO3+wIw0Z/F/e084o/KYneYLipg5kSW5WmGU6Ajdrn+wOA7oM9mOv39
nxsVLa4jjBFOCyr2RWf+kXghu0hkxW2eR1YvEoA7W9dHR/wdxfqfiLL7u9n/
4FSc7qjzWkMpZxLpkhPGgqop22KIRQpMMtXATvH9sIH0pOZcL+FJBry2CZdQ
IrIUFEy9tnAStrCstm++11A/25mgfwQa1POSgeUNQlqzPjCX3JxJX6xAvd6W
9PPScuMjkkI3aqgopTPext9ksyiuE9bJVK2KQ3y1j4BFUtpS5qJtMHiQq3Xu
gVzx0/syVdHeus8LMLEF+PG9Vy+CwMA6wLL1WIVCdE33bFbZoNN5njlysBLU
uAmJMGWWNZXHlJVtxu/CkfwZlOrtxssWXA5JXyzaCAYzqtHgO8HK9U/3FVag
69MvhXPlZ7XRfsiX0xTMbgJ2vKgcAvHHN1mKbrFbm0XKhER5tdOkKgFr0zXT
A7+UHAoA4wYzHre+VW09zajEc9Gc/Jexinnzo2X0qlpmMCFxGlHmZn3LTAVe
p9mjH2n1xN7a9jMNtJA2/74XRKQAcURsfJEGFHnEjRC2yGaj+/FXfzw4TbUh
14ZLEB7IKSLVQVY+H2LMzjb8JNzcjmyd2zieAEauLvhBCNw6dx8kIV2p93o0
3tkyzMHF7m01Uc4eNk0lrfQWLnwn7/Ny3r/cckUOzZ+2uZp4Y9enyHuvcaMa
lCN+x4O93D+iwJhPyeT7rCG+l1dXSSJqDJNwIEAlpxgvChS1dpe5sQA/+kJ8
IQVA+CSUPsYrOetbGvaRKAL/dEDbx9q8bOz3lQRUCrdyvZm1lRozeAgfhdsH
+rG6dplhoUPNiVoUiPsX2F0rxaIp98j9KAVbVMbaoOrYufL2hlA2+mV8rHpp
RvbocO+25s8wSJNUulj1Wt9GdMDsJ5lsp9X9GxnEa2Mcz65BoInJkLTcMmvQ
4Sob4BfxE1t3VVpTYH2Y7omIwzKnJ4FYdwH62rjad7nAgg95MPUhfCBmxoiA
/IWf3eSi0Cu6I0MOj9T25PdSh3Y3nMlU0Xa2MxeCLPFgfyeK6k/yY7As5U0w
QIJpzMVaAeGc/SG6aSN2/1fxaD2Mec6D7OYTv7zhMglDpUejtzqsWONmUJ/O
OqGaYJmKUNEp0xlNb/mVgM2GQWA96odTg1XJInXnACGH+7bA1WGVSIxRxt1n
SzMPl/u66FjakcU/1VaTHAQvmfCsVvTPH1z7UrMUjhYWsXQdmO2WFslZggcd
8r3cb+4Uoq+HMQB+bbINPfHJYkZ9KEUt5j2ISm+7tLK+BD5BfnP4mKOlrTx/
PfM5IO+u2h02BepRakeJ7dlRznhxrc4smfnewbaIKIClkIwm+jmPKA2k50kg
8cZV/rC3pYtv6RdCs92zE19aJJScIX+b7P12ofDRbEbPaOivnnYqaUj4ho5+
w/Yv3ai0LmJ6AhM6dmCTebYRwtdkwDae2weLRgaHHjnj9GTEu8e4ARiuVNbJ
t5wDIQvrSKbT1Ch79WlE8O7QeDdh8+Rh3fc+uaYmb9VdyB0BFR058tAIqI36
C9K3IcuP25Y+TaByKZn0KjQi+LR51KaD5b1J4VLLH2uhEPqLDUSs8sdip4IH
nDebw8+oJ0y7uEgcAO5eWuHqbu5ZBuCl+Mwkr/QOkNKk4qF8EkGb91gPPYB0
0iU/lQeHDKTdbL/37/AHrs950PylXy17yohr9Q6PM6KS1AWZIYtvQXb/RGYt
25KjjMVvQ8lIjQbqD5eqHJIw6RIyxI4Sx4NK43fGD34damfYvWXDKBsSLoff
WnjNAik4ntsooBRGpYzMz+q4qGmMDxLgfAo41LlCaTYAoNTt2Q7xON1oWBEw
uMFrB5KlwExv2Mmwt06ZtqgCj1ucENP5wxe51mHY327IozcXlmCMDqUWYuXO
dbQ9jfmQyf3YYoZJxh+Ktb8hbKIH+WRVyDWaIOnPUMSQg2GNS7ovLt4+AYh+
MtClz5Z39DiLAqZJyPAwJRWZtiGnvs1NO68CXjNFNe2pPPJZI2xIVnBqz5qZ
GfBA7I+uUsHcZFv0FrUxd+CgLUeuAmlvGei/qkucZDLKqb8WZafq8xuZkbMo
etX52JYKRTwzL3kRYXy4VuQBzme150Z9XPvpSrYo6+E/Rtm29pNJG4BRo5vc
31mq+aR08wtRIAiWz2y6s59hlGtBwWdO8xzgf6A9PySM7UtkSosCjX2RRg4f
fyHTrxkddjBuLhUhOKpawvEDTe7FEikQ43vTNhOh+h5naBbTVWd6QeoKzBQD
qfwwfmYoS0wvC1Hp6dHGiT4CDrPJnFQGknhWBbdYibrhhvdKGhxnR3mnAKiE
8hRsgQlNJ3ymNs1nLg1z0WmXfiO5X1133rOQcqrVemyzZIkzEKHWDsV2Xtd+
DEKEboZn3X3xpptad1o6OGJ5vKFYHkCiTziWBNg2RqupOJFwtVS7uRFqb3E/
gXwQ5zOb3JEB+EG7tMZIx4fIy6qNkwmm2jbr1ZJBTd3O6FZ27JgMY1OdlWsN
cal9k0tZY5xw205/+GfkdDsfeCtjUnG7TFPQQPS/2ytOUZCNCsAHT9DyNRwo
bUL4edvVI9Zu27vXHPWOsdjqgw0o1ctA3FOz5bSFp7kbzIDWajCbSna3N8pB
DH+zpoZ9Qdt7sW4staAFssaRbpvmWMp5zO3GyXx4lZ7//VmWzpQkD699qrFs
D/QjEsl62YPyof2cz0giH2c6hhLbUGtQlFu9XHnU46K4cvoXNWz/eJiB+85W
+SND2zTGIoZ8yISpq0gePUeMdEUn7PZZdlofDnv3yFjcN0VWt1c3594t7Ctn
rnZ7TJZhx91l1YUbPPzXd6Qlax4nBGDmXrXMC0T9LdoIyxWzx7dl2Gj/ofeT
9H96yRwvg0oRah3jFzOPdWsY27Dy8cEtOr/53szf/4TAVwOWB3EBeCGUqOmG
73UP9oqPYq5WTnarQwyh/UZvHh8TfPz7S3Xj9LFpppylhWvuRtKy+HL9hdCf
zMU+qc2deesfH/G7onNkA+qG9vxYHTjlVXi9rsCkGKFgAv1aQa34hZEyP2zI
2f/pYql2LF5xw0XLtldFe4SqexBU1IFBKOCtTKB5sWjomeunTzcM0v6X4F56
0+DX0rk4gW2621BFTb5zBwx/fRpSwoG4OdsHBF3X6mVnu3VpZy/DJutqgp2l
JeK4vIRyl5zhPEHQ/VSVM3/8xKHsIpJy/W0oN02jNfNqyDbgXJGBjwW6kUsw
gtsUh98rfYmm3QZLoVnaRLnxuGQHb331S41RLOLBqlEYtM3pZ87b6EV5b9wi
GCTZrCK4uXsyCSlkZPLwZuztxtOHNV7Bj/NvS+qCGtFoKCigk8B6x6f5tbt4
X17Mj2EMthf6nTfWolsOEH8MkHYB3HYDZLPKkpWHwCrHvC/fh2ZEPa2EgGiK
e/5rV9MMu1wWlbX2rUWkenSlxMBf9z8f7AWvMPn9F9+FDav9tFBk+wm8ENgk
JR36I35Q9A6XZ3gww73Tzw01SUcDbUU/aoYvuQ0H7EFigIcBAGl118sYhHv8
BtbAh9kuSMeAiXozOz7sRmzPTYBnRragJ9y3bdwPQ1aQjQ8RpG47yIqvSqDl
lzHv9jZOFtyWV7o05xsc1GYz3CD6iqJEtKsI5obWfIYbsf/yxytiCpghpIky
/gGxPCdVNq+jgGrXRyjd4wqQQK2MJvR01jQTu8AvVAWs2XM967xhh3g2jNk+
SKvSgSYp2PIIcAh5RqV00F9z6qYZ9z+EYNpWushWHWRtiDM/y3qsF6PlmADe
opzu/m81Q050LLsapDKIifHFkCD8Fu+kSrxaszKlePmAAzjMv7lw4uzA2ugF
kWpzLgYjsGhbUCU96oQZ67YobIbjvTAAUj0Wxy88JlX6wmlGfmgDGb9UM8nX
+nheUGoQdvErcm0U+akB0bxpVSljrOEl9eI8iXpPWjWh3WGnicpQUx+2zJTX
fZDF5nEi3CXeOrZbZHI3Q/3oRexM+oS5kS17MJnM4bMhSUeGlG7+DhmU6pXF
ATaohy5AIU5jIfdWx3wZqFnU7oxJYagkhY8XHvYI07dYREmZm2nMDkXNhSwO
JMn8qHXBZXGI4be88dZL0wZFRDwktiHf0EwxPmr+1ktxTMIajvgGZFQHVu+1
1r3kAifAnIOQuXYKbnEmUSUs9VAbUpk3tNqvkVCcd7fSRvDiF2CWQoftx11o
jbwPESYTFGZ+2Xrl0mmfWhvQPidnj+DXQdhMct63FYafjIcHPJwTVjBRdr79
PdD82evNM08NJtOVrZ/CpFIO4BryGJBIe5bq/0FxkHyiKbRWdTlslJqfB8GK
76AwpHbywyM8wzDhkT3rDRSPbCzxOmLAfDYwTDjg+Y8VPX/X8m5y0VybEeZV
wjY9PE0VeLAP+T+ALiY+wz/BOhr/1uQCrlXzIPELWCyDxjt/saGuX0oKTOCp
T+TsZjZdnYU6LUIBOuDdzHewSekNBwnlep7RLjZVaM5dvvisBFt/dIA/HrST
2Sh303vZ+eMmu/2sN1Ui94XZT/Yfl7sq2zuDZ83EbVshqL6BGqi2ik4gxjCQ
9bYzAilSOve6VJ3JTmrVnexcq5BeZ3UV/4inIlQpJTlfzeu2Jq+8RiHQbkOt
11HOAjLqqPegYzG6kbSsGIRNhjZRvTx7uRZQA1sKDlVg/lMSz6NJEjlGDaCm
oeJHNL86AodWsPFO7CTScj8lSJ5OI+N7ZDsOJBSnV4cey5/8j6ds+wMpsEYT
7F3iIB9gu+u6BEzBkvK+vuqJOXtcMb8hPm/Y1t4EuoL6IFPOTkZKS8UtYXhp
5bEwZ5dkqWlJjhwi3F5TN0x78G9pjJ1ecwhclF0z62R3jGmoLkmQqXG6JHa+
vH1ajNOkByswCA+mQJyBptTh4BnqFI2YZsW3LA+Xhzxi73yeFRxLhesJ+Po9
3S1SyKaEeDXr3YXzhfVZcP4b9+/YS3ZvJyI359GT00Z/23eYGw34bEeh5ZFC
7nVX67cTNipVcWh4W1RXcF08nEqutrg30eaAXm33f/NR+B5ureUk9/0qa1Vb
SGdd3py+M2fnrhnqJ+dXUhOFVLtQ3YuMibm+NLMsposK+88vGM356Q0XYXwc
hn1i0g7EU9s34HEb4vJK8NZo6fs6evYt3OkM6hz0T7bH7SIjZO7zKMSbmM/0
ks0ue+te6of8MrcM2zEWTr9BJLq+JPdw5mgMTyavhdZ55Q1GpUuw7dR/uiOU
AsUPFciU6OTTyEI6HI/S0PWRdnLxiEzhPRT+KRq9KpxPj0VC6VdKkAh0SSD0
pc4aMgA71dKNowVOJF+fCvS3uda3M0Z1DBz3hbjnePLvrWxPaTjr+7vFUfX7
9t8HIm+NM2wH3CKaGYyejnS7yQ+SKNZUdTlkZJc7lgPaFim6TcVTh+PMyptY
lI7wklLBfZT+nq2JR3r2ulZlT2Pj9jc08u6KIUE8gnlXxsV+FwdCPvuZdMyx
ctIR2nFzKDIAGLSrN0NClpiMcBSqDXVLwSMj+E4SbjP4eYReIHkVGxNdN8Wh
fHW/knGerM+Z3Lj+LOdAEYh4pXeZFL4O/iEmMKHZbHCU/1AcTMoMH2RAWldJ
hNdchYThngJxWUW90fbmG00xCjMzBfmCMynx82/Z+SZXEH02Ze9/zMK7+F6b
Co9TaNeTGJvuk6sAi8UYYEP0bsAt+MU7eQx6Y3RlbB3leMwM4BL65clMzkKa
pf0ibVGaoSaXNpswGvp9UaydgLghJ/paC8f7bXoYZDM2t2TZ4FuV8cxF7vvK
eaJ5D0DadEAytlg8XalI23a3WaWlZK0O46ME1OEYdw7pGMLx7T1gb89Z0rpc
sK+aMtXArMV4oac/wFcnPRmTd5Gnou7sradZxl86jqQoglXmfRVnkPPZueW7
zt4o0F9Ec0GKNLmLST0cLzOxZGO8mO1EcQ1UQnCO9QIUeCkV6ht9PiqEpIUl
+fRKyPWUNV/FdT6wF+BvZu28R8t+Y0ESMQ/4NmmR7p2S53mQd+ReVcvjxhWy
L+6Frx1uB1pH9rdJc6JhlmTzKq1Jf7xeUq34ekEnpiH0wjbIKSo7zQSgrbNS
PrCf6we7t1+KDmUorSN1YuchPQF2WDvHrzAVQyEqlIL0n8LJutw5pZbubPUo
m/+OCD+FGTjgmY+xKFgOc+z1jKhXE3vYilZ36T1L1cNNiDEGQO5ecRxdvMlu
9EC3vuSwoPnnSau3Yt+sSHlqQ/keR40mrFq49Hc8tcSZtdOPSX1ChHVyBXww
3DUnIG+h7rwpRg3JNmuGL1cDSd8ZDkqu9o4aOvF8R7K0m+bJsFCt13uLn4Mo
HQxUDlA7HtH6R0K1lyc9gVGrs8WSJ+wipRsST1/iyTWN29WP7/YQS1HJxuIX
Nt5/MFTNpPMm4dDoHCSy0kCh72SHROEMRoi2A/fXWEFI5QgqqHix7TxCRbRA
n7vNx2pH1rAKJifn0xBvyqL7XgIXHMqlobD+vIvI3WLt4KMF0ajLadwmjgba
yDAgdPYMx30N3ouFzrd+iolQsxM8rgxTqVVyuJOo3J91Zv0djm7iQYmzpiT3
Hi6+L8xzwTmxryFgrQjnTzYj98yXe+p8ULMzMM7CwFufcla4C0NjgCOC3+Ny
JHhiW1ka3RQuJoNiVcklmczBMUm2M9SLGVeJX/91oFTgDCEry+KZocScN8IP
siTMGDKoVAJwyOa41PHu9yayhQbwJVbIhS/WdcVq3j6JaQwiDFaot2gZIchJ
YwZ1BlxKuMk9xYyRe6c4CRUqFD59lT232PT1jq4ZKV2FUdT81Wg/2gTCN2J7
/rnwNMczfDTdQIc6GHGj4G2XoXiqVsrY4oYAIAdv6MeyDQBezLBkvKoGocdH
vTyfzGFf5oGVfiAihZfdrm8JP4+IT+YF14oKAhC36Q9OzFp5ub9AfexuZxUQ
ZfbcsaAlvvXRqDM7gmuZoZltP7FgYr4OHYleSQzgN2lPijKUmqArNhTRKB/g
bfiipuESjC5e48A56cquL/L/JvJT6Su1ulNJrkrgrYF1qLFtapJRScBTd7u3
xbjoQxfj1FWrBJbbxG1IqvZIPrVBjqkJ5OzDjxsVMAu3qwGXUQ5aH3ODxGZq
dg6/RYNMs0Pxt7OaLRMcJPoDKZNWBrsFYx/iIa99uN8jiCM9AEqloBuyNWYM
t34dnZ4OjXq3gUOWLcrTp+T2U5HU7btqDmx+1iyj7pewtg7t77MT6fq79Pev
7m6G2nJBaWK9oyGrRdE4nH+yKLp0S5tZtqOHqiJK75EkSpC0OXW5ueh0lMX2
ACQcpuWoeoN1w/pKm4Q8ftP6oqmJ/BGOwPTp5ZYnuqxUZCQn+FziYCzuz6v3
UHfSRopSrhLGxXfSZ+ueaGuF02DKvIxDStbOD0bOXwUjwsBFTqjVEbPC9fum
ol7QpBdMki5oYxchNDeTSPDJOllN55PzA3c7AwuibBlh12UtEaRCZqyVXNXw
fFpfX0Vz03hvrKxjXa4YVV9vex67pvCvLrRQHZtLYT/XT775FeujbUrWFik+
9beSVN3qixWthmSI5touYmpRNE6sGXMTlgY5LjwvYFPeOXL3RoU2F7umLLGO
hz/AJ4DUiiWjzkfKOs1BoD1b+PrsRvhV3V2rbXyRY0Xv6KuEAUSi3cdwbLuy
WHDXuMaB+1fXZIpcQDQ8WGR5TXgnnGlpd3u+34Ynv/2TuyXDvX2O/QD37hSJ
XO8PdPOplrUmahBjfbm2kCo2lBC25EMWx+LP//SFDkcaObbTPjW5x4lZi+Sa
ziA3oYAz51wrFYVVvyrl1pfgTLzL32ex5FhgpgTACfbmbQTgDITWVJbllEtP
kHaf8caGCsu5Sq+ylJL9ZcKUdnqVDGT96Yfl4wQ0c8MX76yDWvVqR0Ntl4Ut
UN0Ht6IvUigs3/HrhmlML2fjEsemBw3c8xue+is7NLUmeEBckLEPLwAuFtlD
QwEuZXPCn2IBtyv2klpjlGsCtgmcY2DE9RUlgt/oMcElwb2fBZSn6NrWDuV/
iY+tbKjOuwcq2XLV+weC6SWJswcNRV2ViYl63p1v/gGQ8bdbG9S3HpQh/AMt
7lcWV7jQ0AauKkiXwTm4VvNNjrQ9yg81xUao4Z5/gazCS+ikMGgtiBUHa2BZ
cp+jWBmmGh9INul6JvlJG7BeRb+qUtmHhJ8pd640+uYbeoq15nvlkipiCtvd
2DmlDW5Xj+/vLDgKdeenFJXlAF/sp2wBPgSGOdAEBwE2gk4BuqEgyeVMEsvs
V/i0aSdbe/VNBJOZJ7rsqGOVLw6LbbOKFy4fyI+ooxzyUA+rgCZyQBWnJ4wD
KTJnKEaRtVGhUqLHIrPgCuYm7TOBwr3oZWw7X899qzVvz8KalLmlAdv1NHh9
EObcU94cfSpFBmLh/5hL+75iXBMP5AliEX08xh4UHbwGEYdyAp1iJdkdbhmZ
wA8VKvLHa/Z4jdn4IMw4loV6S5c/Hh+97CF7gvH6ahdLuLTaIp6/+I7OzUFF
Qgu0flLilJ/3eP7elOQeLwQzClYwQE4OGfLguLnIVMP40hzqlZl3RgYWQ/11
Kg7FJk+uAvk6bFXn+OkH+bTYrMkkNqNQL8PL3U/u8A3lYLrHWM2n3uPQq8/X
l8wY5I/ZWAKiu9MwlzLsJcZ1OgYYRJ4SQSQ8VnUR0MxatlMulzvkjJ0nFfNk
Ifa0EvAdLLDcbyycDdUf8OJZhy/oMjyXznBdEVLR0MQ78bQIK6x3Pon3dVef
8olbSc4T9relgyLvkxx1JlDHdgEZrt+kkmjN6eIk3eIs7wgKULPIKFNJ15q7
fPwkgGfq8EEYtR2o0qWqHIFyTQuqfxKWUQ2DvE5FjJjpccXf86r6wnzDB/Rh
MftnX60UAf5wo1QHLJ7dr10vwDU4gBYna06ipQv64xr5TQAXHTT1/Z/rv/Xx
yB1HS+cJlUU+nJDA0qgOnbLje4cJDzZ1FN7iOlZXgjnw852mnepMELFFmHWf
iKlMVK/y1ckr8vn8wQtR5dWyCZhf8PSQVr7CH2Q56S+BhFTa5r59Cb5JxOon
YEltKhzgLmiqmcaOeci9CCsCJRiQDpbYJC84VPSsGL26hfKPuNg0wRyZzD7q
pl4SLSHeCGdULC3tZlNg3K1roLA0hFOu4DfddOz7oMXoeWyXFjzSOZWWOrdK
JAoWAi50XdWNkMgE9B2MJmAimEWA9aVtJ9JYawKTa99RpOLKvinclkq0+V4Q
hPZqE77/Tj2/tOFfjVLEOi6qJsZmSNQZ3dCcN8MNSQW5NiDrY2id0Ts0rm7H
EPmdN/PdrXA2gWeH50LprvcX9kj1ZQ/AK3QzjCwPQ4NBSl9YHm83WG/TeVvE
y9QCL27fYqXNFN+tYahA6R58ep/HKu4bvMw69AGOmiHaddSV5UDlO9RvIcQF
MgVAdA9gDWe/urqY/0vhgPu5B2q5wbfQnT2z3N5d119NznGti7utCvLJNG0Q
S+9tFKE4y3Zr59ZLbvWyCfTPCJZ5nXu3LyGkivZ2b+kzmztwpMlE5JhqS+zQ
uMrABwuVE2C+ewMPKmPbvX/K6m22RgopjvDEmfWYzz24wzeRdX/mKughuhpB
lPn2uDb+n9XWOHsDK/Ge9FABMs277PytPj0PF02nY6wbBPznruzWTFvo1Mwk
K4Iub9Y3ku53uWXBE2S2nZjV7PW4pOdAGr0xqH7GXxYDvpSwopEQ4VUgLdV7
KSsgSZotbFonj1b59a/e0AwtKKobA7hrxmMl24syS+rrR3EYy189Z3ZFxpjY
tMvoeBiOCXiAr6gET9GwJwGR3Iy/8WuPWDXKGmRclUWxaQW9DkYL0oEfPvv2
6z/nSrJFdvopDqKEMbAvsuyqrH34QpWnPzsfQbINDo3NMG+269sVFV2SfXUO
1Db7NQFm5v3ZelmUAUi6dSRMV99w2hhg2Xmx8m0Z4rsNLnK8O+FS9+jz7hhd
16hfhNqxvCTK3B9n6dr9FY8pqo7Xp8avkucJD83b/3JSUrKU5m5lW3zhcVWo
Sq2RgsmODEFlZ2tVYGaEmvILChR641ttxgI9S1MVJiQ4o8xaDA0Fh+/JLqNK
ZwbNU9fEpxpid6nZqEtoupR6hWzEUjIras2w34bAB6Qj6Ox2blARLWaEs7cK
XWAfPRt9tyBEIkA+bOk2oFLpq8z3ynsoprby/bJPV7uMj/PrvH/+jxYt3lRT
X309+LtGDTopLIDUgnmOuhRQIvdoDIJItZ006oW+oqoZlq0CfXLm3cwEaEVD
Emg8fdGSKDdrT3sz4lXbTJbL5w3GnFAVDBuSQYtL/cxCdrzf2hbCcApUKzD7
SlF+6oAG1Z2+xnbkfqV+Ld/sYTl0hq8LmfhNVBFOSk/dCVgGaqGlut8Qr/ea
Luz9SkHpxP51hUtSZUKdAqlLhhg0PWtyjf4K1YGtHRTDxfJ5SKAfD5LDtdOj
OnZgIhmenWU+Fo39r+12poV9t7fztbhgAy63dGLb3mPNsGAvoiTq5+OkYwV/
QMktt/TSsdnDZFL4NaLyU/TVkqDd3C5huRffm73DzH6DlzID4Z6bOVj9khTa
/P8JJtT9SjzGCWnJ/jZHK0zU8eILp3TY71YokHEXUG7lovnRJoe2ylaUZtfF
Pmisz00OODyX9KHg3sAsmgk7roR7GRpFTJEUYJnFEsR7KoBBNKaLx5EnGcgv
efZeQLpfTX+BBKH2t/MP4fIjEJtTmXJ2FFDT1AQ1aFHwc8blL3ajjA6IpCIH
F0VIRBSGnS8kv2axX3Vlls3YvCj/40bo9CEiSgsxcqhsr86lAAO+b9jmBaBv
7NQiuRQdFjdCiJCjriWgf+1cMoTKxFTl8QyopOK1POVFsCAz6wxSOpftu5uv
Al1rbn5Hdtv7zy+0LvkZAaEzybBeUk9jB3S/bELTvG2wkorvwZrhetR5ji9b
AfmfKXvUTQ1e9OWM5pdk3E2ZWmZZuwt3aj5o8Es9HlkdET39aFqSoTLBImIS
nKIv+50udu61VshmIaZJX5Agr6Vals9TdBHkqAs7L/BwxorBhceMtPGHW7QR
9VjUegJkWuJz3eJjcos0mko9lgFZyOrRWaCu1YY3QmGsipNXkiVRUyObvnL1
cqUPIpX7sLcP1VRJ0DSRpkcXL798yx1uaHpFoFvHfwj7kXzTAhs1mo3ry7NL
Je7VI4q4wb+gYD3td7EJ/6GP56ETz7Hp3ym9wqySAjh/++r0KfYJS6Nbweoc
nldr+sCpy5dvwANg3sLfC8vff7j3qDdLiX38nwaiD26AW9fP1iGqVhqwMRFC
fxeIesltrx5h38vAOZRdFEociSEG7HDiNglHBH/CjT1ZpKUzC0PYy215SSkJ
gDFSVl4DyshL5Qzn16BnZJ0hefgILz93eCL00AwNI2Y/FNKYN9no9gKEVex6
hVZnBjxFe0t8V3OfU43oznlJlh9zAahwbnw+bYTGLSQN5h6UfigZ86snYKpo
pQtGFBzz8+cbgo9QPHj/qRfs8PhaeZ1bRyHP7cpHZhiZUAAivrZTmcAT8vFM
r6Le4F/Y9qX7SzszBs8by2LPvPAQmauNHCChZjoubvch7Qs7XRhqcPtulh75
biaVGJeKzFl7rLhV9STmFhSXZh8g7ouuWKje37j43lgp2vg5oymE48ICg5rx
76At7ZRzMUBYBw9y5g0vj+yYH4dYWPT4JeVAh430FuXoqXQIa4fmmirZWLab
Qg/UcfpX+1rC/JrWq0oplzhh5Qj0V7k1wVIIcrssb4leOF3Jc/1p24UAG2+4
p27V4jpArtWE3Y0zyykfohUXkyoGCW589IOg0MvNVbbghfkqz4HN/HXkuFHQ
Bn6ogW+JEkj2yIteBETz3OFmuyv/2TyaNMDl/qpseBZD2gfXk/gbWlt8NlnZ
SUubDj51yYNBnhp7ZxnXpsng6/4Yar+anBiY3VtWfKl5kmAHapGx6ZwMj2mS
F7FAb1iaewuup7AhYI9e/10wPbTUIRyyNScGZ4FLdrLYYOUMQ3A0Ksk2+IHT
Ojrpbk3cgbbtrMeVbEoZKAO1mXD/wEBpwUfk+PyaRsCvO9wqWln+8LzZcwXI
JMMDlqMYYKyQ+276FU7Ih7/AT3dl21xc0nAnWP244Nb0rFOHp9NfyoPTsodQ
+eadVeaMbTexT8x3h4AsvZ6Xhmj8HmNyZxxq60yyAm0/xg/DC09Z7LA4Z/+x
GeaQbMymxbtnbNEOg20ouBlZp/hPC+6n+yLANiCQBzCdJ9hPnmKhUbmL+r7E
FPTOcyR7fEv4bU++7sI/MW9e15n0qGUhiZDckwmtCVjttgfjbF0gBfXQeiQn
QKmc5LrM8zmdnd+9H2SmQYyLIz4qSmNLXDFCIabI4KtNkcQgf+lk5PZ2uJWL
ru7CUp8QyYRy5rvof8Fb8Gy5YPc5QKDZjW36b2kkxtXQKIfuTYsmzLblO+YO
Fd7/J7BdhtUv3/upoyrTcXO5rWm0e1sX1nVqv7q2dhwByo+hoNaRaEXjSZeW
+Hr+smgojorl2lQMyOgaSMyQYClEUDSUs7ORvainsLzBy/e/9V+oPf5KW8Z4
4WkAzy9bM6r/jiIKcn837RueM1k6V+WNupAXcBNGbhtJ0Er/XtnJEkcMzhf7
Fbfuvlq/eessyN7ZOP+AObpyrcm5mWhiZuYYhwTrq9748Mik7tmHwL7UfyXn
+OfaA/hNDF/6lkP2gj87I5e6/rHDaJdH0so8HiArQB/HqytLLMzO8aEOr+DZ
qAzjx7QljlWJS7Otx/IsvWjwAYaLErHwTTzpvoEpbLKUk4FEPM1Z2qAfKYiO
hS/YLJ2xL4a0NG4qMSziJC5+pRoUO2QO/DGTZqih2jGsMtFfQzzE23JcUVfq
WVwkYAujmNhmqOBHETI3X46dhORez31EtbkC1EN8Ao7N/fzKdlV5vldaoqlY
xB3vfOSpUvLL596+W/D78N13xKyjJe/VXxnAf1CXDRL1w6H2KeeOmlPF1ykF
yx0NW/3XxNZ9onyhs9yUnkBLXaXe/aHbkoIR2RuEZuPZGlJAfxkpR0gEICb9
qBn6AYDBqDowKZfpHxtXKHYDHUMnOwWh3liXMeJiqRhBPXtCeHhVeyCxLaEU
07FvZ3dC0D7PcI3QIHx35WdeRPibHQSpfTAEfRK7+KYtoiUm7kccu9Ay0s2R
qpAQDCTYo9T6oYI/u4b7AYUzc382EIaGamvjExT70/eZ+nh/+B9ybXQRCn/O
aHaCFLkb0CQhhuPZ3BPKeWRrNDcywCOO1lEYaMGlLj8CPC5RJkJzRz/Ph0IH
sZhJnaVGG2hTXWDUYxvzS9gK29LvT+esUO9QS2GX8OQkBHY9IOhWlCgHGtqe
QxaPfSkvMR3iv0DjT6JAGa7FGF7batFBUJJxQChZ1KtcpJsNq4m+TVyp5+CM
VewkOgkuarBr6Jn5d8DTj3dKYiTzcQ1MamuLWObHbFTUAh+OXRNN68Vnfp71
gGGwhbfrx5X5BW/iAo37u8lRA60Up9A3yDSeupdMpvpYG1NY3UsVm+ICkD8C
mi+GGWJJ0MCz6VckGtaW0AIwWr3nUI7jwamc+HnmxbRBnHWiU7XKIAVORzsv
nQxdjd/ykOpOf++Jl0CIG/teXt40OrHj7Wgw+eOLddsNeDQoR5Qp8a8fgNlv
LHYls/vgFDyAovz0E4YqZt+hoV0/Bex4yKrGtlBD3tKAGJ7CxAUN6EO0sTSv
MKJjBW8x3KhjZN8Hb2/C6Ec36PJrhtquHDqBhOghkC8K7Ozw2bI3Xx9VH4xR
Lj2gfgw3xcmOEdZ9DgDypy+/q0/YyaMgojp73/RKuVECbIm2oMjnKbvmwUvy
VdJ1XZBe/ddTQ4gw/d8eXYZ8ikg6spqQPfjc7Nh7jqo71CAnC1pGWepXSO3d
sUD+ylFS9S9bSHa7U/dQcAza07KArf7H69nZPK6gp9fnDruDaOiPIHjZWyVl
Oyat+yjmRhGVNfoD7nYXC9540rzw5ojzl/bTyPoKnI4OEVdRFRiLPX7TdIUP
oOCItXWafCj0rWmKb54iVQi91k4VyDx8Wzu/brO4FCWCMvHSiVqZ+ve9gDZ3
WhxeJLlgtqdBKMo5toHnnAGmMNfmLIpViuDcY7cAeu7GMYcjxKou1uQn7Hpr
rsZvaYb19i+zan6kFCBmQHyI16JQ3rnhATXC30jR/Yu1CVe+FL5m7/hH8vug
FbtB/SRAEGFWjAFUstWNj9vAmDBwxQmC0DdP37RzBYLBY4P3eeI2KqiY2LbN
gEs29ECjhKfYwFAeHFUF1K/7Dtay+BWVdpG6v12EzwVupBL/12Dg337xFd92
5o8W3IJzCPmvQ6px/YNRZUvYX1OVoGRUfCchXmGQWAiompvo/tmh/ZLyFFBI
FxZaUDcqeRbJO79E08nYm3TiH4PKy10j9UOqlSSBmGszMSC2SgxzhSV7Sg5J
vI3YnNj8COzn0F+vFval3QZue9w8BZZibNgocof1twLLgNhgJHLKWhga2TDu
+1YPBauSadVcE9gkE9Ato0BgGhHeF6OmZ2ACbYp7ut0WlMxTebzav2CpDX/o
CEhPJVmYc1u1PvICb2YyFAj/8PbBIHXQOafZEukaLCHcRTxKNhRosmXcq/gi
QBxx0wpip9DEhTTKFrAyLd7A7RVWFqtr8xBg7ygPs99cG/CC07iHTREVtaQr
O+gNMkH+ryGGyxeUNmRbaN9NrEwwZuI100UPIwkRDkUDOcpeh6kOhGun0dn1
35RsCC/96W0oYX402NqyulTlcRRTZY2WDkF+I6e1HDZnr37ulVqGDjRRaAbt
jW5hN0N30ywedcjWNsll2MVqY/Acvf5KpwpKAxDH9Er09o7gU2CekmhuEL9o
0EMA+z21jbkU8bzMjpr2wU+ceRuMUl+lOlGMz4JRM43mkbtJ/YWdNgB9PKnY
UMfJgDiPl5W8eLdYcDUiqWqWHEiyxSI31ZvnVmTsKafULdK9O3fcpseldQCr
ZrfZAHatSnGPPn7184XrkSixe0I9pxr+Ejb2U9P8AqRtRs1K01a6GPECpLCo
i0VMMM/KN4MOKfWFsazuSJERw2ZsGwht7iFo4VEXQRfJ1C0PADJmc6I1A9gd
wfpad2agZgdbkZ6oDs4PTGdNhRtYvfErmEpwyMQjG3lVo/qqaxP0RE7iVEvv
gkM7Cs2lMGvjDF7+2eeES3QGpJtFuQae636PanasWa1ht4dAFNSThewgFkUk
yxmQc6UKHhP/5BYsWfZFJvKJr+6QR4hBVIYscvbKXPPVTwN98Y5U2q44KEDv
c/RK0A/kohXfmghZPB0ydljcLe2sRgq3px33q3/OFcdXaFdVeOKHxTJAIiDd
OQ6sZpwfF8l9R0mD21E3xvAzm1C05UWu5lK2jVCZVdggwtBaj8XBOD5WuXY8
dz0ItrBxKEkRrJZh1vY3a1lmVbHDQPhKD7jxfqOVjy1y3M9B9K6dPgvwgEaY
WyBAjlFJM3tjmpVU2Bop1wCW/FutW1vST4t+990R5YpFzojmZcr13mbtClHY
p2Y87Bqt4uqM0mJewu3NZodVYSDfQ4L8KsfWHeH+tFI+BAZEAiWX/qgFWSbB
HLwXTvKKmOCksTCBr8XMM3Qt/R1dxj7X8JcMxHeru23zaObZr3OM7YGt7NnQ
SL0t5byWi+UNmjemfPedTSXTzUWam7405aDkbg+5eGmuksBKbEacaUUcuh/d
Ym2jkzRT0GjKcSdbfGjxDUYcCPoljWd9q+dvZHZqwIXN/qGRKyCW3Na6VERX
3uYrOVpRkaDFGcpRdDt7VjLCrc3MyBq/33dXPR3dDAsiNk3zYU1y8XjbUaj0
osfWSiSEd1KKtVisWuRSl16o2IJ+T1Dt6hcGklDhdbzc+5fKQ8HGl3O6L6iV
93Muw3iLWp+kwPfjEV5lBjXxdjbqaiGRKTBJb0PkaRYh20R1D1vSfqktca28
Lu780mvyPvCQkyiRK7Ubh+3OGXIOfe+WrTEGySKUNzS2AmzLYBtiURFrbKUV
E51fr2s201KwoxKH1VlHDKBNZz4cDj82DewC6sCfjJmd9Cr08Du/SUe7dpZQ
yhGZWvm+Td6PwRso/JlggqzWrp7sYlmQKUMVppTZDNjHNQl74YGYL/n/6crA
82UDD7I6qmiOmkeJD8Y/3QHsBSQXWDw+i+o9aOtdlWnMfMw0fzETu7bIRYV9
N9aDolJBivh1pv5YrmORgZunwolnpUAYmKqvzv0Sk9nZvGbnMb8UOKSs9K34
sn2mZrnE2Kbg9+wYO0D4+wdqBYHuvy8TOOety6AFKn1QedLEVWjFZQ7W+YB4
phiipX8jn9PDc+AyIUwnUi8/2mlYc+llrEP0QIN4TKts/NuehqDFsCcZ2D5w
mbIvV6hJMPV281HazouqLxMxivt4H8QtMavba69KZnV4cG7mS5JluiOTK3N2
Ucm72uke2OvgNdH6qs4EcxRSYC9ZZf6rNnlxj4vclL0Yhc0Sx4QeArWZAiHi
M86hzqlRPbD9Zqlvj7hz8dQVeGDiYICqLZezFLBtLt3BjFOWtw/uILZCqqg+
pRy8RoWyD6KxWmGd7caGE9+dS7JtKLGCXpjnUwqLfLAuUVVQ92GE762+Ypg4
cK2xPtuT1gTSwFQ7i3sdIXP062NtncDuVYrMB85hOY4wNxsE1y8yv+7PdQjT
Vv8GU+mZaf7yBldl/u1mdnhe/r07G7gQgVqB8AeUfplW6aRCW66+p4L1ecio
VyLrW/stLwlKgpuV4S7qvdQOBK1kuTr0L2tqL5kmKm3/aeMh7zygbbdZCa6G
3NrPRhM9GaGm7uZQUavXMa4ZqXNSHahGNRyqljWyFkKTu49LYUL6YGBOVORh
3a1umHu4iHHYfNur+GrjIw7kTtvm4Gs1T6d4V0pjlBXNV7RyImulA9tlsii9
F1HuEoXPSEheqsQLeN0RvyKyTWDacJ7br0gUi32vYsz2FNFwnVC1Rw+3fhEX
32mGaufUOHDQSiAEZgXfWWuij7UK62FLJNOSOpPVVV5dAJ9+DQMh44gw2hm5
5w7r78rdUiHT/+6FbYXpsJjcIVjO1352CQ5p+gpAr0ZcDOGJu+AMu/RXrTge
5/AsngrpngQhMHg5Q+DDAmNQWjscxs4P2jrdvRULeY4VmLidDVLApZm2GIUV
qn+ePALQYqLwBE/ypcS+BnfuF39XSy6dPTNbY0uJC6I2o+V5JgaDTf97bwum
znJWo0d0cRWi2XoSIXnGl9VEnxi36C3SDl+ND2e9tzhi2DyW202d3S2VPLvS
pMG0TYnQbAfeVMYGZw1swSNg/fw7DIjqNBvPC7XYPnhd5C1R7pkOViOrFMLi
aAT8IIDD7jgQAqmIk1bVtNPUlgq2giAc9Fsn4ea7KmugA4IPRXpCR0NIN9n4
LOnbJVlIZmAXuNdMQRTZnjaZBcAVrCFFgfrdI5UhD2zjZJDtgjOpjxRVGTTx
1Uo6I8qXOcfTk1FLOSkChgk4RQoAj7AQqT+wti236LXSBm1lnsxC/ZE2Eafj
3EUT+TSzuIimdz+aftjmcW4sbCd83LoK7S5xwoNJwUggApFA7dDDXpxDZ3YZ
Rz6U8lvO82SYb7SCRDweix/bgx/aS5OXrFVodGd08BI8+BZWXEn4TFuwbnOo
+kG8XxaqJQPftglcgB29Q9vBD574ctoqpTBIYMgjRGFbye87Z9DbtxyK4icT
nuNnTW+psotSvrPdTNE+Dy9EAnmB/r5YM6QwRl7sNJR76jqEYKbtRDxW29Cx
aznYC7MsIVL6bOVfqOT/jyzW8+2Ip86Cp39a69LCzqN/VT9lS3Z1WOkMdTvp
nohvBkqbzUV6twhMh4pwchEZhtfBRngJVzOEliky0jMHkgPc01OHL9bdQSfN
VS/fIjEHJbcw3uHqxtli3etr+YzSC1DL1BZuhnJY7mtSPlkc9bwW9WvZ+I5P
btXOGWFZm28eKv5ioaPT07hDXhzQuinPJUPql0gkF0rlGu1T+iMoPMhUr39D
TLjjGgDy9ogcRQwp+UZ+OpwFZ4BTGvRgPXxR8XE13fLYN7BPJyLpneJlwb3K
F5Do8Y+07ERvHo+LRGO2oYgeURW5J7IZEHK4TzPF2rd9ea1ynZBFRYcv8KXH
eGVN6rR0Beb2oJ/NUqb3f+19pw1WDs32DjWD80JadgxLOzAk7a52RiXS73II
mmzfNYamzKRWuzXOq1t8widtR5PNhF44d20g+XGp+PIVKB5uJwnxKxj4mw3T
C6WOHwLFSV3mKWkV6aTMKyB43k4VEND5h0D/IJ2TU+6KZaZlbQU+hOyuApBx
aaRGdjzLqBt6KBg4mGi27KVCKm/5xyS7z04lUJ/nizM/o1X0vp4rKeTx257+
5m9cmM/E5qGcdZOX17jWFNXSks85nmy6pTsSS2yEaa1/q2SeXuIeJWA8q1sP
nAWflS0n4M9lbOb+hUqkf/RzcfxSIDseYX6XL/a5hQ9Cr1FxHn/cxW8JGzBt
V5i/2aZpft+V5h98odW/9uHB6iRifILI/5cMeNL4gxW6dSY3949zMaxkDZ2r
6lwoLvRLu+bsGxE8N+9++s9e+UPD8lA6OIihfCrb+e2Y3A27MoLnD5iqH8hG
VMuh5lKpaj8eD3RyBngtW+TDJ7KgkJWR1v7CnTmmClivVtaNfebMypDZc2cD
WoqO08IEX81z1xC7SZEml5yEnMCCihh4peJM1XgR0m3/o53TzbvX2JRKwm7z
IrJD8rpPaxzu8G3q5UpFdDdalrAdCazz32nLKh4pPZV5LE/z6/mmXURHgNns
4SQDtpNEDKIMhB2klJZwPBXEnrirKGomeVkcKushN2lyiZkDK4nFyZ1O567T
qUQKeOWYz1w0ZtR/x58LsDWertDMetyCEekoTU0IztgXK3sBRdrfissu/WFq
v1N0xpZoa1P9w+os+g3MGdb7R615ItUYTXFaX7xg+kw3zGiVXlqf9AaAcAf4
odrOocWPESb2AbrYa/FiQfbfn0gLPj5icl9c5MneW2/78AX1JLVNgH4vY0vz
WbPoVRyrTFkv1O+y0qNWNsVNpSPLgMDNvIqKcwYsSG4BGQXKJlw3A7qlglBe
Y/6PdsQLoxDXV0zk6mGmR8Wfva7kVGoePjF3ShGFaI+6aZVmMICp4/RJ/LQT
2QAHIkYkxsvNM0jJCApp2MO0OHBwlty7VnHgIIimvMo87rrdvrvVUFGN+ARU
qyPkzjcFDxCnGVSFhXoJmnP2dBUfjmgOg5hoE0/W8ItmXkAlNLbuqtNl0dVX
l470Tw2sZJDRYduh2f4q18wBAETTBkVYPgxbh6ltoDJojndAvw9eNtgPvwn2
uQCRpi3ova/PfeY7DZcX9LBsSWr5bs9+SrfEXPhHTTk0ug/K0q26oT4CHmt1
CoSnnNxMFPd7OxxQTUCQm1TbWicH7VQmO+5gcP3H6koXGNJUcN32JOcGGu8I
hEXxJWhROacUH7QbIiFW6ADlVheOO8jx61euO9q+MEtzKbr7k1KLP1Bca891
H/COTRnkdo2dVAnaBlRPi4MrBccVzyNSWuWIK3bMlL9j8cIUSkgnpVXxx292
N3LKEXWdJ6jj1pxoiTUNk+6NJiWoZstdIJwc7aH5HE7ZiBT7qK74wahB+Nz6
A+R66JlFOQ8FK9T1GRGoExZBX7AOPkeLc3C4NFALFqIIVmxdsLJyi4YpSamY
HvuBr+Jld1aw2NE3Z+4ohgSPxIZqXxZW1EOSE5FEYmMSM6oPEXcL+9oCXyQu
2mtBoyP/cvMAtmeLOjxSWyMmuaY885xLlPPr1XqOmEg8bS7Gc08olmTidCL+
g77+1RM831fmkSqI4DJggwarX504FtFMXT2kHwfEDKQiHJjuRcEUeP10zAaM
VKJ78VFVRUJU8iOY4HaeBrkNCdyoOVZMcDgI8qY9Pz2qA6/nvgF0ts80N1TG
VZEtTeQJmNE0Ptgx+iU55QpfVI/LoNt8WWTMXHkQo9UME4lPI/h+/uDFxFTw
ucFrfGUj9RXfxY7B6jx7OVIFhJczLqj3J7CIG62slVKJ7SQ2JuafYUmlpDVZ
3nKb02MwAG7+q3nThM7bFE9L2Mr/zF3736oJbzFaqgTI/+/wvhGA7Fq4/0wK
iJ3i9IWNHP0S3rkoUvQkuzQ8InBJ83e5RXi3jNyP0yCAy/Xbag2OhoSBIfFS
XonIFcNM+voV9O7dGkKgrairDZqf4uTl/6MKHC8IuYZCizwMBBNsLfT3E6u6
sz29b3k4kT72cMeeNGeGmXJPn+IwtJDoN2V0E5C0kx0cTBBpVYKhblb481b4
tV8zNDfowxK822iXHQz9Htf0aPLsDdvacTHo8MHGEIIQgmwKomCCaN75UCHq
VXwukW+N2H0rM+MP2WwHy55F+vvHAiUOmzcZhc/F2Wuj/v5pwaPuT4cTaIzl
L81kZkRBMNk7S8g6YACU0H4J3vBozHPXyggMuaFjfNyAzbV0HTv3zZhiC9mJ
fBUJ6jADbMCq2KvcE7Q+3g4hhVj8eKHybwUeJ0ZJrwmV5XGrwGrJCi8x+k1/
WPYyIdVTMWn/xQ9gFTwj8zhFqVxV7gqyusrNPKLAkGvA2BLRE606k9GI7+hf
kqunmq1r3QmNCryHX0jSnLHXo2t2luVObOvvjhw4MkGcVSAW6j3nu0zvtOjd
Jwb+cpK1I/fHE5B7RuRzgnEz4sL9HlJGc14PI0RB1nEGnaC5bFcUXY8yi93W
l71koINnb4ik7sxEki8j4+hsVkWlOoSPABb0wlGD/+BSKZNBagxURS9B1+FG
8+uPGyr/riS99TOm0Bu1Bif8r/OALZ3HKdMQLJtjZRg9SD1e4ZvcOFymA3VQ
wph8PaLymqy67bcvJ8EkVhFT5Sqq0KbQZH/f68Fayr+omSiWyI+OWiSLPUoB
deWq2iHB6SJm63ZmsZwFIq7siEHnpzt50xlYCTzZ5bR0AxSvaxHpBgnAuPIP
tzjytit4FVq203jS9WhDKhHaYzmC0Ry0uZtDI3Pvd+v+pqSxjWRtIhMcCFVZ
yH16NYcptMCPLm/J61E0a74IMkPpRIXTU3FBE/PQsIGOAj4Z54Y+J5TkeHtr
XipWF0ZQL+5e+5Bew27pgYcGj5R4nK8ZaseQpOiaipNxEz/ylVOkm4HiLFF+
vSSLNQiufOS+gZQfQIMCl1Wpu543XX3gYSbuBfrGjuTw1DbTJn5YRRKnNZR1
YWmH3efcxK2sYBE9uOD/BBDTWhTLtAY12JPRY3eBreNq1JcdD5SAIw5hDF+i
a54PWzfY2vyzZgaOR1uht5ZIdeWG5cLknH8CxM9GhEkVxkR0kVZ5lWAdGujX
0Hq8PJ6kMXwWK5+qdxg7IoQtjzBNwoDVYdPcPbOe6lHTVdWJHXzQEEmT72vM
ouPwS/4EBgnbEZfJW66ov4iVp+FpB/fPSAY4Av0vxpaYVjJyJxRIcnf/nAec
jvheANj+OsiKwalox0MTntR6BeDa14OWXjPlM8io66gU+Npop+0G/8Pkwjes
Zf6aGTcogIpI6jxuPxv57im4qZQdncEkk2dpv0NB4ocKokkYiSaGVXYKpJgM
ohs3UztRzaESsZgO5efxSk+vnIf/pXyWpp91tHpnEGJIwIKSbmpbukESgbpE
Nc6ymU77EH/HzPznRse3X/ArLNUYNtvnIB2Y6moS0wJddKLVtNlczHcrZJt7
igO33vmODhSr5LmVr72bz6VS9KXVc5m2ZpgaC0Fze0JCdI4up4Mgb8+GcNBt
0S8aZfVemE4tRIH+Dvpo1zkCtgTo3lY8Gjad8rLgicRIS6lXTbBUXnKGuPhp
OWCtDQxkO130m3xK78QDj8hj7ClYI/jqxXO8JS/SlH6lIg2sBmbveDrMFDTB
ZiESAvytnxkHCbMwo8hoLF2AbIBeb6UhdW9pnNUMm78ihUuPd4ZSMkmg6wND
nWcXzJ5kUQF3Y/CEkYsPGP6Pq7CzNmg5dkyCBq4Zp2mfqqU9NH7ZtFtbucl/
tVGXmD762gOd8DAyCEiViYXgIukwvvyk217zSOnoBJk3ofbwruIAFf9tH4/g
MeWfWOs/1DbVpfVPVrGhYaIB8qoQso1Zl/pycbea0uldth3tgzmKbdqpZgIA
nAzpDAQ8M4IFHl9as0715kM/bvnaOQIhgBJ+X0upVuzdW3WmN21pc6B8JFZz
ckloU4L7StcY9xY3cN4tQuuv0NOfFmk8MY6UHmlzKcX+v1Uq2zt+Z75AMYDw
02JbOq2zUDv9/iJ/fgl9frVY4FnCqz+P199568pbUUGeSEqAxI9MlCjiOvMR
RdgStJfWbbrfqB7SQKD7+I7kvIj7SUPxKAfewMfhEm2k8xDajdFWpMJxOrmo
MmIia/CLnDssibLJM/rmGsdQK1jinEQEJrBJrPoQaLEY1nJrMmjKZ3Ivk5mD
D/IWwWqaQ8W8ruB2EhT4fqyfWIxuhylxTqAIID0UKVNzZKDePhtXo0Nnv+j3
s/8E23q2N6UA1HnVgJ8mcns3YlB3HZQDmryvFe1MSdHf/tj47mKGSbrK97pm
+/CDgcHh717hADlnlwWym4YTH6qTcbAuyQIbkIGn9jEG2HuJnfyMkukiSBr7
YAsxU2U1ZHSwtVp7xi3o15XX8m21kGkL0mfWx9WbcopgJDoOxibYiy1WRqJ9
470PykxOnibDrDwUbhH+TorgjvRLTLzisoiIqUuM8iHNtedi7QauMZd9qTvV
rQm/eQ6IDjwPXIXTEJJmcMcoNfHDIik3Myf6gXa5BsKiRvLaFLTVNZmqxJ9+
UPg1HsHkO1NnUAThdQhYPXe54MkAoYNJReFGMqFgdoQ4rsx1H4jY0RRZJARu
saJJJe2X/VDSKIJjz40i9SaUPzugN4wdK+LbG2yVegq/C5sdscfAwrK38nLC
ZMem6wg4RE/gw1Dj9Fy2m24Gp3XY48yCSb4pu5k/0G77J4/q+G3R1JVWM8Gq
nYlYdVP/2xYRgs16KeQCd1O502zGZqdT5nUxBEf+ELnTA26K6nvfbrnwLOqE
S5h3s0e79W+f0l+vsRwucCybN1J7EgnZIRrgDuOz/LeerhneCekVwTuv31ku
Wk/abIM5Fi0hVgtll+TgFMKpae31FKSEeS7P6Hd/pYt9Vv57aaS5gGsr/u6B
QXX9ZHhVHkmfe2wKJaRi5jyQkOkKWWVBl4hblAllVP4gqg7zzq40RNDia/LT
SgJHvBuGBPXG1+Ly5AkNAkRpROeGsri426dM/MpWndN59Yk6P07+EPT5iOh/
5ZwDag+vllFjw25TleqpxngVTVYcwxoRT+fFVj0ORVZM/XQHWppbkmSHCz7d
OcVtOa02p3Gt9BRKjSCO62se4sRIvZ0M/jA3+YVKrMVaH30VBADmgqmOzAIp
r+LLYK7+iC2861lncvVKf+1YOKsrqe+LlJ5HX5PL4a6CYNe38EZyPYUtHiMo
SLGCuXrS9HLVzqQnH2kkS4W4vcRjJg1Keqoh6OEJJCH96RPQq38VVh9k1yv4
MnkahhuYJmWZHWCf/p+9sHrexNQVf8Fzls7+nzvTAniGAkvRo+t/RWAvV9XC
gKNR8mixb64y+FQtzqA0YnD/7X+OF6fdBce66ie5I0NmW2PV7bytv6ujjpwh
dmfs4r5tu1Hds71NU8d65yDRt4de64Qt9/zw7JBAUimu8JgAVWqrq4QQdc7S
Z5J4W6PpKTiKEMYz6qyk5cZwGZ9HO4zzRZ7C8Vr6e96/oelqPJID5+GGbDLu
kccoF8d+2MFOBqsmEJAF61EoixmweSsSFVB8pOE3xX3FPBwU+8DjuCRvQj0J
M5ItGW32i4QKHm1MrLFkPFfIaXCsem/FBrDgzJ5hmha8mUoj0w/2m/zefr/s
ZLQkCpbEi2/02PzU7ydSJkOugNJh/9yxdvJ7aqGwP89/rVBMRMjXhfQD8cGV
iSqHQ54eTkxXhUkKzQ1jggtN9/H+SK6vCi0dXxNYm5Btsa3YBU4VnwQDAAWZ
h9B/5yVdGjOD/ES9/BBsVMU7D86a69tFCSv8apbHEN8nYhDMx4FVKr6L2BcN
xs9E4OPXwwVlphFPX9ap+6nfXbS51onyWB7zbKpnJviFcdHml/l1ma5wuWf7
rqFJ87VeCQ0O5dBLBIEl+ylxwlNycE2EG1igUSgQGogf/LFClCxoW7xJQ7Sz
WgpBoDP2vLF2i7RFQ9JSBkKu/8p2o4DRjHdK0Bm9GNpia/xLdG8ha6CnO/sP
b+asTb6lCayCz1Ls6n7VcI91dAK+90j8fYl8nugDQE15xcl7ylPfvq0b0PJl
2b7VSyz0MlwBJVK2mv7qppGE6uiA2Nyxdar7cR5RdqEZWdkLa7I6LtWrZU10
JErSKGhUFXTVu0cNy5RumvhDd/9Fwp6ZDRMeg/E+wPHv9U0PQlpXbr16/VYl
9SM23aWw5BLFfXkAtXvUsjbwsXLBoAdTAqHgSdoI6uHE3mnnaTcJy8qrwaIM
PCMkz1wRX/ejjeDJjLX4k44IUH+fhF9dPE85KJHKZBlXDlUZUEisu43BhDQJ
Bp8qTbJrnj2pZPcMmlZ4ZchF2mUvl83C/rJNprcuH6erPKv4O6DKqCs0RS4K
cWhLr2v488rCo4UrjUr5kYkTJllKzi6I2tEgwDhQQmQmjGC4cNRsJmdkw15a
ObvB4GPVFB/l8qE8V4OM5d2lHVgt05+e2Atx1Cvdivj+J0oe9SNJ1D7HJjdH
RAi2J1aUY+KUsNpkoXTQMRUA2kkyqUEXMLZzdghwp0PixwtEzgvvNlo082lY
2bTNSdk+XMuR7QXxrbEUwzNe3fCKkujU4DGOYA2TsuHn3SgN5srjmUyUklIS
zNvlLUjgx0Qe1VmpG2n/cRV47fMFJDSTe8KFPEtb4TafahHC8akXldAWPjeC
mjESoUwqA3Qdh3W//VJTvWkmuqCZoAWKz95donRD0yajYVAUARTTi0gTiOeT
ttu0s1A9ob56bWrjlaaAK9E8Ro66FmNNvepkyAAUonSfY/IhMOchnCbcaOAl
UghA3I8/1xrAm+de27TxzLvNrQ5SPZHdmZgk/RY5OufEHCXIbHVGoZMXJRmy
P0smLXEVjTSEkCO9YiQaPs2eeyM2mh1WAPr9qgeI2nzYvci21yrz93s88yBr
9/duKueL3c1QLaEzxpqb2cdjzMpvUeVL1g1iZxcoHbr9EqC6QZuWvcN+RmQw
rYcsODjzkwl6ZsPtYbpvgNq5oDdh5MqqZ6lZUnktJufjktbkcYwTxxCQtW5W
ciAfcLwOFowwsl6PoBUiOTJZschuuuCn6GMs0yl0R0BMh4nXgjIawsnHSd00
H4/J7n1GGFyOXx5gxxeIjenvRzzFOXOHZIJYoB6sL/i+phTzL1JEa8qjG5C5
nBO2scJwEMvBdf3196VjWwMkUafzhrMRo7ZR0JQHz6vW6BjmNJ8gjg2XC9Wd
c1F6c5NNubEHfSrzTHr7u8VTJBR6ValT2OnnMn+vStNF2JFNEPoberZOxEH3
O6LtcquY4Eb9WEhgo2ztWp8wIW1v30He4/L7LeVC+QXBH6+zqLahce2Zdd+F
h1pXuVWDLafFSTPk1aBIMmaoHfvsOfTDVpfHeZdf71/7vb4QxJzx0v3ys2id
yjtGSsLMspgtoWRGD3fH1nzYHU83eUhz2/lHOcLHkEAIeFvPl+2sJGcWe8uP
IvXtceBVFdfYOKB+0jDHMb677yFSMjgauqKpDzGoI2HPvDm0HRghWbgZOyXo
czgDzblBG3QTRtxFzTbu6XM0MwSckPAt2BxVl79bogB8ECxDBsCbRxdxVd3J
0s3IW+FMiG39eyRXa4oS0e4EXqMIUmDaJk+lqc8x/0NlD3m6AbDoLXWcSQXl
bMJSfgJUo5TDWvOpoLEwxX3EPTjn92sSlEGg4ZsfEwrMyzRjNqH52Utgjd/Z
DwOx8fhwXsGyhJvcg5rqhRsRDPq2/suNyyZ8YXClg9S9gZ3xpHgkmRToKsgP
lCAdAZK0CookHcQoO/jpuIkNKwE/yj9ZMNPVvszXKxkdc0+l/QxNJBhI3Gtt
WzBj9+dNjsPD+leQWT2oivJFiKqDj5547jD0l1UJP6I+NDlSdLyM272039nX
INVC7GhV4Q/CmFfC0a2iUerBNnfwlasWIgzEKEJ9rUApHDZ5ro5/kMBfPAkj
MUZyEtggQMTkIy+SWJO6QXaB+mFXDA1Fb191otCS+Ncf0ipu4R0p0bzs9NKf
xZatblke1gnR9uVE+dIdWmbT1H4vkSXETnSyC0bGh3BAwXlLVqqsqb8DBqp4
dT1O63qLqqGUqVcwVefZ/Qcd/sKK83soiFWI+Lm8GF7bTHTh8EuCF1iRZnPc
eVQCT8dUxTP84o+Gx5SnmM7Li7OyRf+laAPUr9tI2H2NavcHDcQZL3qDInE6
5xGqnLfBEGvJCzUcm59O722Uv/Hh1xRc2B+1hPNlHdmq9nGdaLel3N7irGQw
JwiXugh4p1tKvI8YDoYbZDz6v3Qdnt1Gv+aNmaAQgtw5UxEKt9ilE8W4cJMk
EOA1myCu0hjQbsTacCCc1yVRy12GMiuh3+3bZjAEYGTFgMFk+IFtXVkhn908
8yPmt4fkzOnCtafZrD5F+5TAmtW2m7I3bies9VarEJGsdhQAphRSwEA00SXe
JwKMgB/QVXcIEptT6kb5daEdy+KlQLb+F0hX4TVsI94pXjy/pGpOvc3PdGk9
3WQM0+WltkEmofgZkwMVe6OsDPXH9ks2ciahvHUViBt2ZGySIOtmj62cFrHn
NaIvELVdHNT/HzegRf6xTSv5l6wSFoLZwojiS5eRUnDgPDq882zgOVyQRMzj
TDFZklwp3FD/ajMhlk6T6M6ol0chFIbJPKsU8pktyK7P0t6VP87Wsz3Ss6zq
k3LwYZQkHsz1DJT+RdeeNFJei6BhyZuAYV5Fjr8BbKlpsCc11y+xddramh0N
YRWFnYTtqCfsEYEdDO5hkUfFR/PE4xXUJtPyKDditGTdWbUc6b+8bN7sG/gO
kGwqbC/y3ScVHw6yFhBjRohjdmMxCphOSEOu/WcsASU7lgDH1ownZJzdTRQ/
m13DMZ5fN3BUPu+jwKEO5R1QK+4EZCjADC9A5w38DLb/5ygvncD0z8s/1bWi
Wf6rqqASO70vU+g7mb4gK+0dNJbS9fGlaCls2XSNUzdsoZWa6EiVhdriUx4D
/VcMf9FSvmLUbL7RzcXUDdRtpsmvXFKAxZe21kfi/ENaEnaauCIdwzl+7CBb
kQqdGuSyNUYVFDKeZhYPwDWWg/jXBVGqOmcOFANlsR6JHsUa0bRVVv+Tr4I6
26SGH6Gxo66BLzlio8IlWip5vyogoUceZ/WGoMFjT+5XezZvUuIHeY5MSLRb
lK4bwbzgH7J/3aRFeP4rP3+zIE0a4SvOdQ6LbbfAeAsz+MU/2rySuZ12w482
Mau1ShV2ycDH1JYx4qRBcXlhJw3Dj/qkDmEzoHXtnbBImvTsL80fn0rMq1r1
kF5DXD6UVXU2LQQPbH6BQnCLDZZOfoREIbgtYYo788daqlY52Cu85EydHpQO
fBGmRZ4oobW8Ta5aAVD7yfTIX68V7gezuggi7dZ0YonarmWDeLJVJN5qHQSB
RBQfS5lPmlCW+D7p6g2FQErDe/wl7/g8HOq/NAcQZyD1QE7xDI1VWjuLMahU
yiQdnet42FxKotKu04emN6DchiwDwa33b7u+o8fGu/1g1JDDthBq6suOA/hS
XuCaWMIQ2UOtj2GempasTdRYDGxXDccxZ0qFb/nsm6r+aAFTd7BLDnaY/5w5
VM1pWL8cwaEpTdzp9YoSEL+Fl07Q4m/D79WjfoxfMjEaoWvCkSDmmvWgWBR+
IDms+izJcRkdgl31sptxVyRZMCjCKlsbKxx/gwP1NkKjMpnPsWIgh24oHcRC
+NDRxjoYK9Wzo+i29UxwG4RQFfjw5iHWvrwBOTwaD8ohsEM25BhUA7igK0Gk
1b2LyBJU2QBNOeXNt6Hwo1kRo+B2u4cs2Q68QQrojggMJi9E99/wAipJv0T9
YF7xrqHA80Fyd8iAc0DWglLut1qPB40i13obZQ+vYRZ2meF6KZtUq+1YVo78
JVVyFLxnbRuQQZe+Vqe+Vx6daFDoBnOY8lZVZCJzQZTXXUukRY8NZhMejqTx
xaZAV2ZcfMC/0UH8PrLii2x5EsKsN9sOQOTcbo66aTJw/Py9art5Rpl28rSz
tfCyNh7rvVKBDji3dsjqS7Yr10lG/mo0WEru+xl/NCF3kX16+QLiyMiHyUqm
u/gf6g6n7bhkqw+Sj8LsnHxrG1DHdkKBPX8QyWgah9fly4w62VotlQWjWdzO
9BsixmetWtVzLq0IbuyPAaAaY+NVNcxTgo3kdLCKNCMh90Kl2Ou7nj3K54Qw
pUSkPzFupJkIwKKLLcvFfOtJVAfE3CnYskBWkNwU9g4rhYRJ9w4mMU3InWC6
wtbN7Ytg6s4kb5tUjEIZgiqxiDFT3qK74sftkI8kdd9f4SbBxJ83LrLlpvhJ
hg5AMdtupqKRzi9gN+VhGbRzNaSGrmd3bq16DV6tDwj/tLYCiLhksv04joJ1
ifHZlV+BPW+065+Zv2+6Dn+KN2lGFBpKJhfZa6cA7hdzcyoPozEvOlZAKYFZ
3eAiePSjjDSajXjGIvDvzFT3sjr9aovvNq0kly30FuuNTOrnsI6w/VXxbnFb
w/xNq7P8M0nFJvHLFMCsBW3UMLR5oIx9QymgUiFBeU6g5BzmxlZpsZpUQ3Sy
1mln/PQ2rYa8atvoCIjT/j3UAtopACNq/r5bQqVdfxxEOVVGqAaBcDxeX+wd
FYPuvqBwYXrlvezVROAiuPtAsh9syAPKextz/YlJkhJcCax68syjGFL49VhK
z54DAwRbo0ZUQfGRp2l0NXOmbfAHNsvtc17phR0xbSXw2GCB7MlLqsXMpIRU
1OZHegsiYHpZzpwXj0LcOLAR02padcxx7Zqov4A5sC/uHAPl+evc5wP31baY
oPmELJUcx5dulEf3Y8gTIOedB2SfSmAVaAt7nTPATsiyKQ84Aeqyg7yd/Efb
WmuK6whpCI3PUzsmVLk+Z2n4UKMs7ksjVWptSi094m2rYGOIGG1GX14cEed3
M0ElbooYCB19Aa1jZUmhunH97dtXsQsdsRxJAHn5DNzs2DSDH2SyoPbyDnSD
DMw/o0M5wi+xLhugRpcjuFzwkvzgtPFuMq8hws9FfeJGv07pkmjiqudJq1ZM
bCmrM6gCZDBTuQRdJ4kwVyf660rZdbrp6pjJtIiD+PRuisVCRQcCBaGwDpQE
WPeJcUqe0x/URY/JZHtpGtR757j28agMQVSrXgg6BRg79+OlEMzQS9/9GTiL
7MPr5MeN0yJhR/rUTTKecbYQzMRhU5EGIue7l+AvzwMkCwfdTZr3G8KHhNhU
3PiQbl2nx/rMqpMtZIA2vWnFvxG7Ch5R1W/gRBIxX4yG4g8zXwiPjtICPOo+
NQlE87MrzTMqHWXFSnyhnTRr4UWp/wMy4fKGecTZiELUG46X5S8DU+caUAz6
U7WvD5hVPWtRwJoO10Xe2K7Ew3V0Ul8NX5VUp5OuwZJIsEfDzaCIBry3D2ka
qYj6L9ckcUGdkbdGv+yNjXMat98a9R8ujALrrvmAKAgJyJ30n1Vi5qmmQ/xa
PGi5+2dUCNk1uSBbRrSKqmz/gTJnrZkEb3IBr98H9XVMLIllU80vtiZQBeok
Uk7DTCCLFcWn9fQtP4c7pb+GuqlORLFzsv7q9LDxdwNGds+IF5nunsPTuliQ
oTMPSKHLpKys3qQkWUS65kME6enX/mqhHOu0GUxc0xwDqUWsGnWJWHMVTjyb
5QJvEfB0rEJHMxFviafRI7C8Da+qCsPaCYCHHG+o6vKwparpBmI7Y+Ui4hLG
GQSnmjJ28DoOW3AEgKsmGj/DizbUopmtpJEBG2WUF1vmnkseRGwW1uCPV+RJ
FLe4FszehdlLUJbVdTFpr+CIobr8ABmT3pq8u3mnLS+c5iyshsmOOvLifUKh
x0Kl9nWfXZZWVaFLGLc6n+RVoFmB1fqqriaDR0gI6L05OC+P/uxMlUHwUM8u
9j6yldgt+kIPhhjpvMZknQZ7GisM/tf+tJZICQckkxdLN52ApbFsmjW3AGD9
TR/eVBxOABwc2vpIMoqN53n1q5fkne3kW9t4TbXNlJHR3QST9I4cXPnATihl
w59v9BT2fbdoAfAuHTsEcK5Df8fPEft67AwbLt/ZQDEHEKfPL4vykrgqV+8k
WIKXdlNBYmeqNozZRCv8NS7Pw2urYB64afB1luy46QZ0Yvv0UNJOZsX3Ae6E
5HE+X/tKy2geV7RbRGCGeCkRKsB/7eXi3GHI4raAeuAsDrnEa1poda6xYFiV
cdzmK/ndwWNdAXS/2/6SRxs9EC6uMw/vrGN29KfEX4uPhyK/tHQOoZ66vq1Z
kBwdmTasliCZm0/cfMT5yqzPhUz6YeNssFTri0iy/2JfvEfuZmzzZ1UxbyiD
g+u+5ulFb2n369tTFeN/hu6A61RFOqy1wlKgBqBTv9vDscZe/pwxZB0JcooK
hzOfXsdSRpLroGxTy13b3Up70fg+46jWBmfkJKTIr+vf5VD9SuGL4kkCwvuu
GGxaWdQT301n+QnlyGEFV9IpKVjCcTE0lDFIWOzPMzOPvY1VV79RfB8i2ire
+YfPehF6h0LDmuw8Chiri/RIdxPATtXeC01/YFZ/y642AmJmchpki6jsOr4o
KAymcCbuQq+A9ScyRVfOpeu1dc1fWAs5M0TD5TEd9/oflpU0UN2hKIKTu/qX
lthitFK7cQeSd6KHWmLN3ustIyEC6I/G32X4n91+6ynVJCRWjnvdu6QQk5EY
KLG+jNBmElJraNf9fdeFvYy1yxN0xgMQuVrUXSogM2XabAZxGeMWvwinJ/gG
USW4q3bFTVIm+lhRjrd0StO47d0yJ38KD3FiTej/cJiG/ybOBgxLvldGybmk
gB2zSZ0/IxK7pKVo9piNYxYbd79+1mTEolu93VjSIY70rYU7Mb59wNJdDoXj
F7FlE3CloaGqCWScSeT67eNnoPdD/YMKVMGH3CmZnrqW1cGTBUiVF9JKKiW2
qNhmqw1Tx0A9qeL16ySiW8byVFh8d9WnzxBMYT8RnZ08Q12u3R/dkNDUqSlf
fxoQI+mhs3lnqVxfksphdAbb+p3tmqcsS7sFhZN7PiYojY4YjMB+yj97cwgT
MzNkXdcPcHtS1iE0DRWXY3QH/mHKlSDHneyJy+xsdzcf63qf2RMUN0Pqwi7w
9/367fQTKOQnLlW2sV4PlxBwwTPWIAvR6BKNUTDIIk1IX+R7Fdu8Xz8Sw85s
qpsGo9QUod32PfdLg6Lwx7B+Ndaam2oNiI8kwx6J0+SPe6Q+7QuMRCMuRvPf
pEK1e4Y08D8DfwLAgO6suhYah1MBxLS3es8/70uNiFgtpyqdUEEa5CtZBqpJ
MxOKIaH78wymXqUPrfEC6Ld1Y9yOeXZPRXLbz3pDROmFr6/BusIChBxPxhw/
864ZKmlZhsIGOmGIw9tN3DpQmfGXRhhsX0PmfEI23BDmSA/dbp1cw0XLiVmQ
ie2o/rHLrfPGuGB8aKAJVcENPk3PLyejnRMAsEg72eyyDrTgJRnkFUrCO2LS
S6/gbdyGQJhJFKqX8YlBLDzyJSsGrgiw+kIRhmLvr6IPEkPw0DA3tXOqVdD2
Nd9zH0tvAKhnOX7OEjYe+f2iHeafWc/Ka6KU+Lp38xOZE1T0cFXjV6bnn3/x
29Kf3hCyp4f695N/TLry20afZAKhjsbgY7WEs7YIeG9IaXoNaTa+vPw/10dh
twLmCD6ZBH7BoF29eYpi8BAkr4/eNK5JjWA7br8HNW3/KmsVIQ8AVHG/QJs6
tMP7ffcG9igXjtZbIDHXS/lMoUAuKN0lrJfMH0e58/PrbXl6pKTkEdVV34xV
VKnGnz7xwgol7sugxXz2MmhOn92lTSOz+Q4LTE5qq8y07YVnUkNv5dwBs28D
Oo5nuyXQZCEvwZ6AYKDDX3YA/6B3rFsh0foHRkcd/9Fwj7i+KNCWeFd+OxRZ
bMZjYAHyleXeHJuyicTJUE7C8UCVxWp4PgMFhPUXT0RTPQl241oHFfwX/jGs
Hm/UZYrHj70nnTFDjCswPr8JNQqKiR50+I1gxcm3WWehd+sAKp8DynpSln+V
CzakbBz9G1mYfSy3Y3Q+GrlJl1BvRx0vzuVz8BgMZCiY2PBC/DqIIQRRIFEW
q1IIt7mczKuw6bKIe4EuU9Pmj0yGU88fHomRxFD6gY2D88er593eo19bjtRj
GKmc7p1IiClhazGj91ZD5ttMsk9Vzl5oXsVA/QHhlWgPxzrc3Plkz/YDdN7R
x+QkTDHch5DwyPlW/Ah+zG2ubBwwegiAZxMbzGdqLwRDv5F8Dno4jMkmXKy7
6tJNSglZGgp4EUpNCVlgv5hOOmOvbvFAS74+JnDKYatqpaPM72nk261oJ4Lj
utd4NA5WVe3a3jHnjHZ8QFbqrF9Ano2mZbIp5pGiGPM5EPcTM3SsUQWijnRj
0gg4UVuk01ZZRDYjb3/ZkKpMJzvZZ7YsW82oBhGIWsDrZr0r4zuD4TeGfVUe
ndsFLbCHuM0v1t+6dAwXdkJ7tB4OCF3S5ENho4x0FRdqrgBY/o2xNovIlzjU
OY9epS3EwojiLmditEIuaxT11tyXydcFI4uYgSnwOvR8RGByCVNwIqOwTN0C
2uY0AAW6/OwTwVceuwfujv2/kKprBlUFLG/QeNq64OPHVUQhEtj+Mx3M2CPz
gTvtkSAhizOJd4q369uEN4aKR2LhjZ1xd2FUOgO0FqH9f6dO5xjbPrDkL4an
Xx4nglD9PI06J1/y7+p8TJaUHsIsqdnshc2D/9YOJoIaK31gBSWJTi15W974
YoZd40AP7Om2ZH089Vp9lAEY/fjJRlVasqNBMELlPcGJq0NrHcCQsx/1RElu
iRr4aRV3xQoZXTKJ868FUrz4ysQmim8hLMCKY40ti0MOZcMOwGbGam24Ze5I
fzbdiSgGbmzTLW4u8bWqOkpYwY3royZlIt9Qq84vxu2jiqMQ9/ww6WdKwMI/
RkR+N0ANPM+O1eqzzba9SMuQY/sokwtIDGGMF7VNsn8lwF1Vf8OYPd36vhI7
fKhlEQBb+ILjRu5YCkSLFEaVXW5etT+6VdkjJTX3RIb9SkRDigfv4m0Ce/Ef
fOQvukYimuQttsIszzC/6eFk8BGZ1J4w3JevMp02dfyCKZhjs9cW8maAR80E
Em4Zzg/TnDiFZDN8BOxU/hdKTykX+SvI0iWJDWkhbBiW6CvHWGcwGjcsP9u1
oYMEbdFH3mmlbx2Z9IKOXajATmlmwGdTPhVh+yXCkiqUnE90bUV7Rkcyywox
s0PH5YMdrogGtFXdL99JGtXVUiHmLKSmVyb7XdFmJwzZv7QI4MNRTx94xQt8
+nGsZ7HZ80HBsNUhVpCasnmFNfBx+9ofyUKvJ1MetShd/6Rw0/1XlZF1/uV5
cLGHAQF6h9ebqFQOr5surbdeHrkruXT1KOvecfs7dkND1NLs4W/j6X+smjwN
aY3cU7tLDIN6RlEYPuNp0toGK0r7A9wZCBH+5HrKWSJ/bzS8LGsmHitQ9hJ6
/fCIv/rFGE9+AD3SsINbIisMDve3gVspWvyvkLXTGzWWu7g5mvYmtSQtx9CW
miF9dCfyqnQpzzl2VU7znOEfJyHV37vWIWjoJqDc/iPIePLIAqMPNcYIyU/h
GdZlWKNbCZl7PMBm+aWIqMjBXSR3Mqg6zYTbRrSARmYCeaJMNnjhjaFN7e/V
Dv0w1Qu+lIAcOm/YwM9YlyJrdee+wXKw7r4IxDokZ9qxcRoNOAsGcXdlnkmJ
8/mV+ovLi6QUKaGGfvDzK58CNfR2aUsRz4EwwWLBYBAAymcz/EoPP0wLK2vE
qrltcWJ8ZSzt8YN5Uja6XKDQ0rHwRDS/SxWKwwNu8IkPqBLjcCNYa/7ZEb+/
2zBtFxfJb0N2PO4xvh0t50qep4U3jKAIQNAyKZvTgKq+MrztlugXqoKo+yQv
4zqfE1ww3DlTcUBtfgd33M5fLrptOF9Iqz6s2ZsS3cnoB5qKlNGfKj2i3LWD
b+R+nKkyG+7n2GEvbkoBEKzPFr1kx35hD4UiWkx5xNoQ+SbbFHkYN5wHvmVc
9PwHDMksQHO7Ehg/Elo1z2NIaLh56JGHew955YqmVw5GX8CIIAhSAlmYtWP2
7uQzSRCodAc3rWKs4Wxpj6El4VH3WiG+6dBvrlG8baHIigDKme/+VX1CKjQr
vstZiwBz9kouK38aWAXaUyzADr9VQHPdh28wVW6knhcFvQpSgwKzr2C3ekUF
cCd1f0hm4WeY1GmASC8gAu01QXIUmHRptvI6yhdy4PEoB5JbtJbzAXmuglo9
/8m3ARiS5Kj4QQLTw8vbwlMSsSPiG9cHBBVyG95agACkPpepSNEQ/fCaS2SB
/5YkAg/jlJfpnvuh4ssIuMvxsJsoftWzdX3o3EBDaZW46MO90er6O2QNxgPj
h/HVsPhtNw3gvbPzdZ0Ns1W9YQYMTl5zsgs5i8Amj8HtttVNgJ3F1X5H4v+d
8sMeCTkuWcOvBCMfAmAMBe5by+WuC5aAhtj+8R2aCR9VpgWzzTyojMCADk3i
1UmbhXHPCvyG0f99xsZiTbNy5+l+ZGpCStO8YdQJc+ZxwqHZgq1sghPeijBi
+VhVoyMhtsKS3XsDsakptO/2O1Fr9cSOfR2lOLB2qe+J97CmUcSeNv2HJXiY
mwSsVp929WJphXNZC/cm/wxQMf7d6RMMjhDroWZyLlaMSC0GZTrA3TcfjaKU
S02hP48SfueycW+hffY3Hh4+b8Vutj6UfF6s1lpMItOshjOZ/5F1A09aE4Xe
g3Z7KwaNhXF8YRjSem+FPXCuSE4jh2WXkAh6KsYR7FdaldBFAwz5VFlDwTZ2
ahJ2pYxNVa7jTB+YjW0YUd2d7dX57hHaHRkI6uUVpDRoFZN7wDOySZAMZa0H
rwZ55VbCsVJk5N3JYJj9dxrE3aCQZB0qMOkf2MRsWd4tr08O3hYjLNdDc9Bx
8ivJK4cs8vcbnM9AWuwy4s3emQ0u+bTsbotTyGWAgstcTse6DWUbOvUmxGup
YRwNiOkjR+kwXqFt9VPhhpGDL5st4L694rgyPiyqtDpYjnSraCkpmuk2EkeO
q5+gLYfr/VZk2x+lVtEu5gEpEh2TEZKT0HXNPSbt0o69kfXz1iLdAQrmJSw4
vyFZIGq2dNfaU8uMJWpw2t896QvcXD/daYZhnaa0d5OmKXwPZzMxmxqWogfx
kNkxsM+Aug9ZKw1NpK0rrwAxDSnpoqKCEg7LI1FgJV1+A8XpFxlmD2swfAL0
jmMWSC/a7aMlm5Q7/Bfu8/X0yk+qMEFmPuBKtUVL6l77Z5z0yRjznSh12Xtz
5oTa0gZ1Wc9z0mKOmgBUk01whql9AXOpfZpUZFBO5osmysjlBHa2VWKbqiBI
W9zF85HCnQIkA05Of4VT7F2lp0haS7DEyHlOsJYOPkCB4h2s3BEl1OLmNdZX
zQdMRxEm59q7t57iWcqbCvQH6PKKM4YCqqwH9EcxhXzwqDY2ehUI6p/9uxW2
tQOaubmpwaf5m6lkPIjQWCtmriQwsH87k/ooIlcutswpsG9mQsFIhc/PLnnS
E7nJ/YpnzMjFFXBHebVz1VP4oaisNZ2IA9eJlLKM9+eHVpbmJ2HF/T0juPNU
5x55itldX+deybdGjX49NroJgqNeKBetDTPeGTzNlrGSs5is9DakOtsEpBKL
shy2avO8jNkbKKACk9s/dfDiew29yjpwMLcjGrDLq/SWZDdfUx6KfMVTD2Kf
drisY9oy7JXk8i85n8KZRmtE+MjbTpR06gTUMRy9yaGMmT6t9fFvJgjofZrF
Yo0KL65h91N4FXZxFKum4sBj6gc9sZSPQo/q/WHkmrhxSgJQCTa3GBUzpQcD
g4agYhpbrPV+cBi05z2Qdv7VEhnD/ofogzYAOldZCyv1gMbHGF8CQHNaIL5o
rM6F0LbBz+VOXura4q/jidEBjv4oSY1bv94q42WsrPy3SJaHmupNHfcKCErE
SaGoFfBYWvwnUyg3XbAsqnednlX/naSyXDn4yQxjU4qk/rxMe/QKTTAFRV/Q
PUtdF2trpR+h02KxZP2dbeqMdtJ/SSDtoRBEqlgrfkQ4S2NjKDniONxBt8JY
KtToVl2OBR3D5aXj0lCa+4Ayk1VYJ1NKP5U5CpBjfYDWPg8ruBoWKSs2Weyy
wFOaCHhmM8r4mIj5ZlWSP7Z+HiiHAMqk+hYkhfCVqkzB8YoyVw/K/hbSqT5F
jWYGoWQq07FVcTzzv6hGCf57WUMGeO19pdYE/i5oXncu+tIWr5L2aS2yZpo8
vVmPA4e5VNZ8L7imlt1W0IODou/cGmfC3d443okfMO+Kmob8IWSzivAkPPoL
HXnBV0Gfk6nysJTcNC2B5OOKPyb/18I6SUoUIW0snKVgGpEZeKSeJ9R7oilD
r9MKJKZj9fUQujNT6531AWSbuNOsAYn9ehUQS1PG8iDf8r9SsiPrbAi9LHzT
WZ4bBc8rk430UgfLk2yqRYDYJUBj8lLTIwDvRsiaRQ8TYou6MkXcmY3UlXfp
wx9YvK6+k5M7cFI0Kmx83clhmy5Nnybl9ecRoa0+KBSUGkPI81SRJQWjdZGg
TGbCCDRfcU22/qfcOdb+ksmL6Uj0rUmsqtoCIkYNYafBvM+yTySnusKx3MMa
oOMPoneZ3L1PqTHHDHjMEkgVRlEkG/s7rgBs3vZ/mEIuHAVRUjd1GiUnsOrE
eHkMIzblyK+u+P146/icuYrGRHwZsmnpeEIual6FaZkvKdFPslDQ7zkXY/pN
E4Zw9J6w5QL68jM6cwwewG8QZfpNcg3mdruzZMCdKkJZxePo+GTJpv7K76By
wlo4d/PzIsCQYsbDNrVffj+sw3inG7WHiXB37nV8tu96gdXw499WVKWUQgsG
oohzKQgUtrsd3fW3de16EHDDWLed2T+pYf3bTBBxDWVmsTYSasNy10h29tRW
YRC4gNbqGRhIy+xMwnAmvO7xQHnp+omIZjnTTK5VSOL9y6gwo4kRTorKq7Ul
7xUZ29cF2vkCa6C/2kWtk+1tDQWaqtnSzXu/uIUT39gM89q0Ave62+gGIOCM
L47vghJNaWX1wLAK+W4e6yJEz2aB6RcdFTefz2wkzgtn6Qc6r2TAT0tR3e6Q
qsTDZXdhUBlwOctet6Sj8r+RaJqI2xR1aK9LoK37EgX6oxLdvsuo1Z2FLVs8
mFO7mcKJIVj+WOOA+YD4qCs3Xvv+opUiIIY7IN8TngSbHdfWWMugBc9Wn3IT
5STJUQo7idsXMdVL4T9Brr2c3cTmHmL1Fdm1eDtsgMNgxOTE6ATXpxXx9pUC
LsFIK06mBmfG2boBwGnJnqIRmY6RPeq0Mgi2TxBddjPxNFCu+HqY6t9c7lOm
HH5Ur9wFAvvlJWhsCg2jg+Y/cnSctXwzYJz+4hqiU/+2+N+H9sSSyB5zobvu
QSFtrsQaANfS1Ss8wCRKsfFMwO4KlAKeF1XxX9fdOK5s0jJV60TNwpspnzyU
U415DOc5b/0DXvwVHY0EiH28SXDOtiCWrzdRXLhOQ+unWwF+tJiYC+yijvWY
4Ys8aJYBkjIdVnZrN+jGCRoJ/H2VRUFLu0mDYF9XZf51UFPbhcSOWj9oSuuU
+tkID40tVI2y1NGGk6AbhpeoI1Vone4br+/E2pXRBXgWxSW1KWSRGhfYohBW
Ny4gnbjaIXID//GS1u6BuqrLLBhKewM6mI5qK7rrpKKe1JsKv/S8zakz7sAw
v8IjTrfb1CByyZMvezcaZiuqISlKwNGc6WRYGIzEBLhxWjRsAxvFFkpv7jpK
aZFaTFEcLDGR5hAgKbh/KJdspBgiRBAaMwlZ62UaS0zHYNrkRYJXzAuMxOAk
Oiu9sFNI3mAYe5zZO+IbEtRU5lEeQ0HJySBmsGnzj+gogS1KjPwZebUbsSQn
3ec0YmiDZmLM/JHLCRDTkgBgjdIBX5wEEmKtWbIdjZmMmK3E6RjlF7YVTzzb
QdKE4hfP5wIbj1fwdYmPJfH5twE5sbJ3tU0rEF3b5Gh4Ryhwa0fq1U8h7xuH
oEN+THxPG5xjITJFsVZE4q6wpv71UX4Ji3MoY412z8X+sbqFAhR24saf/OWi
9cCHsUls1vPMwmYOhNEoH5ndNB2dtpUI/yGKVaySeE3cSkN4qzc36g1ENJge
pGlK5q0UERMFkR0MvgyCaPqIbNvHQRnIpsFksu3yHD8NzrRXcUfLy1L+Ke3Y
kpyxosIqL0h7tV70qVe9xIbM8DRqBH3PNSW4J9RbMlB5uszne5tkvXp8qU3T
jAwx881Si3Hi71ts9cAw41/UMipWqz31A2jxxkBbsZ4r5toP2KP/ZZk54YST
/bozYC+FVaj1q5+JpqCWcmVEDKZVWmNwOt8S+qHCsFmiB8oq6QRIajW2R4NR
gp38cZ5ZpQt6oRs3VHbddYsLpYVlj/dWLMlVih3CBJnfPUNK0TiMQrBQUb9b
OdB39ffU9KUhaykZpdslG+wv9hpA5+ZssixPoMQsXWDvbptr1NcNTcGA6IB7
Z/Q2UFFPKLYVLtVPAY8NEuGWoyykbR/SZyYH2yLmcMs1IHhjywTYm1rXYmme
EIfLhEiUebbZ7rkAnN614zhe5dELQRNQ60Vp/tIZdM54aY3X4/peMy31mL0O
Xa+COPC9YVQjUbfP1bBxp5/IXRbJkjrzbp0fTKqAw1AA0dq2i29O99dXH1eM
u6K/h1KpyBGtH/aMbsur81yBr/ZtDLVMv25CRmXlkveTz38k57lTRBT/YQmW
yZ1f/XK7It1LOB624mKO+bB03WNJppTEiu7mPmRYaVERbGyaskmSqG2f6Dwx
9C6Ihyj/fAT660udlO3kBqI43aSGvRQOmU6PfBVqip7fU5lPk14RUJ7hZsOE
nUxUu3q1BI4rK/SwRh/7UYyYDCDi9/qDmJhhYE2buE3Hf7JOEeXzdK0zeKi9
wS5dhMNtoDkZaX5buxW/I0hsyYneJZBZ0yI7Cmks6YcgRkb/2Omi1qcx4QmD
3xMLggrbDdjlQkb8r3OdTpFIM5UTxkzEDhMYHH6gefpm2O7PKc4MPew59TLF
0NqkShMH+D5aDoAWAZemXpCqOOwcFpyo7kYq95++FqgnbXdk2ZUa6IOaYa8u
0sjy0chCZ8VcGu3n7fR0frsl5XSA5NAgDSNjwO4Cl5/fqD1j2GT69VpY3Xsu
wjDU6CWRS52A+DjUZucw3kU9BCfcmjSkJgfdALPxgGxo5sfGs7rm0aI5Navk
gVZBf+u4DQy32cGJgyjesjqAge+8Nn8gF7JUf+fx5vs0j4PXnnGLhNpj/LNl
RnGfAczvxFaOp6zo+B2VLML7Gi2+UmwZwtOMqxpQ8awIwFNEEuVxb2eDTRMv
cQGnu4+KGh6Apekqvd6zl68PP8jPGgb8/NL4QeQxY6YPuHcjfBjICVbq2q3g
VRzLNdhItvi1vO3g2PEyQHPsQLNGx5rvncJo12wyR2PivrHqV6+4YPSEGE4D
AyGeNUACckDcizeXepk4YLM1FPonnAUUWgYjg9awur4gU9VtApxrNCbeLD+A
agAIyCAqZgTNdVm/qpd7Mvwsd+aAbcK5LxPJm6uj3F/KeE8lJZdmEtZUj2Tg
U1HKqEl8A8mhSNulLhsJAdkwWzvfdV2ouESL1eTPo06qcvRy+DSuaQ5u4PRV
oxd/z5ESBiiBZE2+SwXbv9UPzx2RlIDC3GSvfG/auVsXW7b0U+ILOuppRFDv
YT3LNxVhawH+ReK8UFUUOwf2DuZgebsjLCfKbG4VsvC+aIagPI76BF2EvKzU
bmc+c4N8+ulGI39HF+5Tl93uBI8Ejl7f+Ef5evW64bzE/WMYTYTHWClSBiGE
UMgQJw0gepPO69fPHtpMWJArdHs05zTPkjsHIN3HdhvKdcjynxnhsw+w2INv
r2OJ7lJhD/fraS0DuZH6KggTVfy5IljC+BLjLAk+anbui46gusLI2H2n/kH0
UaOGxTUb/zTX9f2f5u7Zh8PvHKptZIzp6nc5lsE4InW3ec1id/1gqrdcS0hU
08ztrwyhvHk5T9+Nq5e9ROcmd3lB1HuRS+ZJJIPZGAcZkJ9SoE5wzeaYPnIF
HfUeNr+ajxT7rTlXIiMoRqqtwBNDWebZQb8jVEeMcxvNsgPSwYAFIdzse+uX
mMssi3vdwAQp2lujxpvFiTTQ7IBqF9Q9Lj0fHJUyUiGgd+ufXVy8FNUoX922
Ey+CnuB+1pOBlGPXK/4blOfOjcpxQ0IvyICivySHD7SLlHFUGHSFcqVz18u4
gSFN/Lqd6hQ6ViaepWkIzUh2M5V1A3pkzHcqloqlBzXB5Lv+888kiXy2vFfv
iSSEvgv/lEGqhXVuw1flLV8oOFvZvGkeuBAn3lnkD2zLucFc7SUp7kmRaHrj
lZDEtJl2goh0xL0NgYbCuuDiUPmM/zrMW/MxMIxn+NnvaQHtwe6END1daKBs
C8iA5IfDoQZ+bImtT11oZusoCXfewum6uclYNpvM+w1piebFrM6Sa1mjvwV7
R5wA/E0gXJJma/91nUwPktAfEc+MvK2PRU7+y504Fhv/t7FAPcvaXcFW9Vbh
RExABW8hJlfY7Z9BWXksyaE+AN8cFkTKgLCa15m8ERTmaE0k59ByqssXSNh7
FPxZuliMuiV2ejpTGX0hMMQvTyiN+YsRl/zgV15IsjNNvlrINVNmnImwRJtW
MSqWbvTzcMnH3h/p0mreiFJwHcX8Xb+NTcdAZlF2RzwvS1OBmjJ4stQzxsYK
GYFu36Y/qlU9rcab40YgvoAQ5ZRSisetijSJO8UEjXHRmSQGw9V6MhwAG9C/
xdcxAf2+aNPJPT+2yFzwJ28moly+bLH5SN9/M5jZll88Su3f2/HOwbVnZeBa
sQHb1fvLjmfKkjt3FSWn77KNOcA7LpAlcL+tG0l41Vu80wbH1nYWe+IJJIOi
GSEAbw+p7pANqX7bXuCzjnOun/x7VxM5URaNeMZ6wSBHblY6a9ZCvAVJvSz+
TwUafpH6eDm2Zruo+TnUN6AP1SvYaFCzOY8rexM3gl6MmYdcMzNX2/T+Esr3
fl4udOcoPCOSU7Ko07HhzPILwN0n7T0QEAJEMuxSGgcylx75SkLXvPi2NnBc
+jWy+pbjeySyGV6+JLfz1hkaJuPsv3/SV16eoKbXQamXEuGNL2f8qKBeNWFd
9iz+Wvp2+TkU58gkdNBBGWx96Fnaf3+y2wqgTAEgMj6qqcnfCe4ZaKU6BUWJ
Oy+9sHLMbN/5m8GsKvq5bmphTJ0CsG11vjE5TpUVNdg62cJuDPcsOSy33b1Q
lH1TCCJmcSuuN+wayTKyofRyKN7YikSCEmrZJUan1Pp+yBCIU++wXUCuD47W
D57ZDuhO1rAX7Hdo8xt5a1MH5pfh3DB0uHshqYTH4bUQ/CwbRCtw2WBG8Jmc
Bomt+grlE7AiTwwf80/dP93/EEGPbt5QObFKpFkVQG8hjqPklZGW8FjGFNHi
zI6Co4lLdEmbcjvl+tvf/vfUwojxygaNyfgRG8MGq6VLfb0CPui64G/f1hIU
OkHHiv/OvH06N325fC3vOtzfNS3U5YxKtjIlrKbc2/4qHqTe7vPXyssO5Zgn
oo3YCtJ7qOn63lfG+kI2acu8d1KN7ELbzkljJD4cN1uoCpAWS2SDMqj4/1LA
S3f6yQpVzE2yk0hT8oy0Q7CMGmSPp2bV7bgytEGG+RuBCfjIwTWPFHEu4WBw
DJmgvYDDseBgXLmv0APHLGrHKAWOfIdJ8e/oHfd8KEYu8mlK7qpGUOBD9UJ1
z1/1lmcZRKhdhMLJZucd87/++UhWAwG/48nWW7DWiQvSB9bGO5xW8TpyNYQQ
9Bk/u3mVoU/AoX+2/aiFIs/yzTQ4/WIz+Of6UVazJ3R6KQKJee04tOpQOkE+
Y/cjvkRrqxlsBcte6YeMwnVB/53eo0pkEVFvhIcNjs6yG+DTt4hy5WxbNOSz
z0AOnGLNLfWDGEI0w/8VKf2R0YDjqQP5EungZ206r59qrVMYIQdwCGI4nRcf
ISGmk2PCHmXZownwRIlMfg7brQ/O+Kohm76ajIWwub4ExxCGJ+6GXNDWVb9r
9jwbsO5L0FX4L2wx56ySGePlNa7JFE5p+4e+k5kCrpRk4V9T6u4ny+9F1Ash
g+6xx8ikSjpPrMz+lZ+nw/IKBioGhicH8enNNcd1fX3naUxQBdKfDVxQypQV
pTE36qCG1+8hOomj6SBdBHFXimIP0iK2/NOMeovJi6dKar+ySHaGLfXJodKA
wVLU5CP9wDBdf9LurFqhTU93sKLFOEOVLimGy19CAbG47IVSuStLR723OxbM
VVpIGeoQeqNhcdAu7I7qAW+ZtQgtw5BYfvA2KFIx9Ce1uLHnlgfRTJrkzLq6
aCquusJvQ66R+x2eO7/SRku5rwjAED3iGcpnknkQV0f3KNrtwaYmK1oEyZHT
L6/D0D/3Ex6/V+oB9p9FfFuiHzYiYVTn4gyZG0FarPoEYCsnZc38JpG182us
BYNtCblYz8mjRZaWhas4aAZmPfdArg6d6GTxa5n0RA83xk24fOD0fR4NY34m
uqFeRj8VOhFsWdbWVocKgofb8VGnzs0IkTn/DKT/Yy/Afd3hVRPL4vXLxQEV
rRze4rtALIkGLqAY/s+XPz6s/yQBCv/Suh3sy8ZhbvVu89thmg0zsOlLoArj
2gEi0Ikgk6QB5sxeFgjxDGwHTOKGvUwUS8ODmUAWuiih4FFSdxBWwnVEoAW0
zizchCjfW7grre6SaXFNfQArpmR/hOQvo1CXmyWzweCidJ/a8zJaDjLUySDT
gvDY71DILYS0aopILfmwjXyGyLFAxYDD8qq3bRyDgH0CFXqH0fiYZhLSt7JN
Cj8t2Cv+BV/RGDodUuWCyiklhgyhm09870Xa7nEcm6ujSG4WIA229ejJ5tyD
KDzVqWwBYjHJ8jSTyL+Xo5RrKoca7+fOLLTMiX/7y4UMivPN9BCIFkrrkHYE
7LerqNwSU/gHH6wQgAhQUANi1xrvpOwaepqp5YhLtpiDkL4Lwmiz/qNTnd9Z
I2WD1dyy+Z4rfiophnyG+zV1DZG3QXNtULfE9X13IUeCNDI+hZwJEgQMMHUa
r5ybmEehk/DPaQS1WKqsw48xgibwpLLxz6bKXpLUUVPV2PjOlT4slp+ZqINK
qpDYlhkcDg6ddVfOk0Rey3DxtzKKowIXMG6wkPaqbZklpNeQNcfwi6Vv33DD
IBv6V3JXzSu0zDHyOsPafztrOxeotdUPlBIAWrOQNSugxBuUkhWGkO+pGDw6
7sUW5c5d9W3PYJKdp4Ix8xqqo2yINrK3bbjdtBJtcMGRvwgOegMwN7CNGhgr
PgcTVBgEivmoxED0hxSyDZlT5ZdyfVGIA7/Unt/cOxI1eSnHi7JJ4txcP22t
8500t1heDHvMkq3xdLupu2kqI267WByn2cewy2AC1S86wiEA1OVkHnHXrkMJ
vX2tu3e6YzpE5EYol1bS2scsH1nZ3EKnEuJvT1Ll4mHoB2u+b8QlNUeK+JI/
ULn61qIZFMNJQd8992mcCmTpz+1rVEtQ9P1caJ3VDbDNTz9QanepdZX6Fh8E
KDBt8ZzyUacBogS2OuCxHjv/NMpx0bIIeGT5wKFhoRA5bZl+8mkRwjM4yboO
OxjTRQql36S0cYf3a9pWD9OpKWH6X1yMix9O3VVilPLRsGbvz0Ysb7GBeIs1
UywIosyAWvRQ6+f5ENU0MkrDEv5b8ar8CKLGhutK1QDSf5DVYSkb0ySMSdZr
3FGbT403121jLyZxYC90/4JU9DMrAjOjlX/23FK/vNi1XQuKurbh8WHxs6/K
oXwbmY0hkJkaC3Xcsv6f1CtYXnBM7gVEUb6TAoUZ6vY22uLbfbHO39BsZHYG
KH7yoTn1DpgzksLzdgf4qd3ij/U9IdrzZDCfrK/Le6B9cmlj9jpb5greyg6M
GTJTUOCrson/Bg9mWpj0bYwlDbGhugQRIZV7hpGIVLaZfu6lPLtddCDKpU4S
mtHCLpr6q1hANsEUdspsy2N0oGLz5sBJJfa8RxGO6sq1myL31eytRVmR2gNh
oqIxx+2yGRYL0Y10ndHwX64uGE9NxDsFRjWNK2ArSR0xk/u7b+0o1J8yWBpD
pIugbtxDNLf0Kx0v+DKahBvJJRRbkPkBMKjfLvtW0QcqCnYQyXMBd0FVRDzW
LpMipmHCdNHg4xrp/PozfuxR5vq54gqLroEO3y19YFek5YcWXuBd/IAzVWHT
tb3fEdYOFuXG4o42rdEDFQxW7frMwzvidg7FbQrDUyL6Ichq/3Y0UpJpA3QQ
6mSkEzRXZZOqYF0z+YGQ0p3gOIOlRaNJdvtIdd4bLsvdOjvQAL5Cy+s7s5rX
5xp09kKuZvA16+0pZr8ctpKXd0JbJ0N+nX0s1ElV7zwtu0uaRNs9M2WLWr0z
Q8j2G7mxs1U01pQr9ZpSXZA0Be2sdEOILn8UbcT1mEHHfQ0NtUW0MU1gKcy5
Ipnqvl6RTv9JQlvi5g8gl0xsqj/1w6Eo6qaSpldSP3rmkKj/T8LfSZBUai5j
wUBejrWMFIFHtOtuQQYEY7nF6JJ1NnigSJ4kHc1UZ3TBOkgdTBAAZNCixJOq
RiEnulh18CDYgqTfzWcPC4thsIr1yWXuGSiKM/oK1Fio9vE5V1hU5sDMZGa6
vRMJUyBS5/Zqjcvg+Qw3LJ5Rnr2/Cn6YrZzngu62S8LKcWutJHbweSIlkzI/
lw3UqCIw2mYuuKt5hWLP07EvFvx5D4EHW4YHcvXtmIibyGwQPZPThAxUU4PJ
E7n+Vnh+u5trEDXiSpEq04pkyZQeuDNugMe3x5eK2dMt3hNR9+24f/dMjz2z
uY4GVbA+A1emtRacylg9ztLOyQTj5wXP4jybg/gOTjDhvt6sg8ZFXFePJDgs
uIUbeoOrOfIgq//wo7dt0R+Y0YU7/R2i2mz9xzGAZijKKlB35sfFrCjgWHQL
61GTXhR6p4NZTRvp0jKgEzpffwMMHTcJPzyEZXfIKX6ZNC82oH5QmoQcyiHS
C5+EGH5eGjyv8ClfqTolUkLWqx0Hxoyh7jWCK9Fvpp3dnPzCAqSUvg0PraX3
Ge3RpINUIEUolhUVGxJbalAiKRl9efzYJkE0iSQA8wbUstw7fjq9P5U9fsUc
XN1wiYASJ5LIM3cK7fOv1KTpZvcwp0ZTt3Gh+SOmFGocvGehgmsK02a/pl3s
r/ff4/Jz3mncCIkh96qvzTperYR+eUb6x28OxQVScdT4fh2UGX1X6XjsabfM
fEjqfgd3DGNbeG50ppGl38drmi4oGyz2nMQpmIWKDW5mLXFbkQDdZgrhNGQL
X/WYCU6szIf0ID8Ff6zioSsMYpxQBUsunnUDdPQhyXNqVMD4G/yJBL35DPO9
G/hXqAXJQwXWNBD55hHCVnalT9/ZHos1Ri7BP6WWiHhrP/dGeJU/YCyyIyGP
45hEqjmZmeB48shQxTZHCmcROqES3Haw1gZ27/8JWeHwyumD78Uzrq7ebRPf
kiMdxlarnBpjZwC/fUiHS4W9Zrh3rM+3ziC9Jvjnl9VnB+s7a83lBzq+0QmQ
tN3V4BXR8V6NrkfH+BuP90VwU3bbneQpQTsqp9pQXiKKszZ0nKS2HUcJUOj9
yHt0NBcWamXr9rBf+gVn9KkZQfNJs6Ya+d1eg4qQADm9zRWvdJ4NpFowywUE
tjrlS7yGc7+mGpDkGCvTvTMPf8MSr1coqGm8+OVQo1v1EQqwU6nwQTGw5ECQ
vzMDQPugdg05yP0200pwoEm0SSV9JxqX7la25PM0390esQJA7vm44Qqq8Qke
PsFAs2ZydoZxOJ+IddK8Hm2o2OWcUes1Y/hVNUXzGc1NowJ7x8CQUqvGc0wz
ItdstUlTMOq0wubq8HUfLS9TVxivbDXt4OsmRkJXfoCU2oCjF0XIWo+V66R5
7LTpq1mPra3SH8EIhMroXV+ui8zOc6eoUA0MAZSLettZFEYGkTb/ZE0HcSJr
S6Ke/uVNXauiXI485dY5wnveAXUiKQ4FB4IjhQw8g1wAv2x1vyKirJqyXONk
FHCYAaGoph3tsEUwf9Sb8dYxv51e9r8MHvCgWH6q4pTHvSEHB95jzzpIIj2u
jlDwD/axZuKqgAr4Apf3Hf4Tk8q/6AUfqv1nKXYGsH6Hx77QxksmzeqDx7Yw
ijj0gxl2f3Y10MocF/LFViSNGgR/y1PIkPg1Ms7mav5BZWXBq4TXVtr+iXac
1o2CPxAgPI8ZdR8noDcl1iGq00WKsZZsfy0d67f2Q1ovuBwHpaunM7P8lDFp
nXo7uT1xlxCNPaw6zW9+c7FE/+ArKPrUYczAPylWiiVdV5Xh0XkWW5i9ZeMN
Z3EU8DnnqVGCgVJ929EF8wcf5cmoeU9lGhsPwiAKJ9hT1dFQk13pWdI8Bb8a
OTLzQ/dFZd5nrcjz0PNW4B57MTwuqEIoHM5jp6Fc2Iw9HoYTcRvoLqLVT0X4
gGd3/6OCXrwieVx+Bxd/G+hDRCJZzLdGtqP+ApdqECmsjpqy7r4kWKcaderE
+hDTpGgi0B67SLsUhbNkIkOYea706wlv+Nkipmaszn9sIW8T2ZDs0+CGSXMT
QZsDSm+MWqQcIrzGrBa92KOUfJuSaR4/W3bryhJ9mCJgVBa5NB1PFbGgKp2e
iOnEuOE2YDCBQoggd15cIExu8pyMPl20fzJgleu0VhXBxeQ8vr+HbZ6f+RIZ
aVy1qfGOgQ9k5qq3fdV6HQz/91UHhU41B+aMQtq4XswTruilggigSd31bAw8
2+NinS64cvAkX17AgmO5lgeF4moVT9MRnERYbwpLriC218a7O+AZHA8aamyO
buzCbiTLvrOIRKG+X413mU6ftmiUBEaMcvjyEIe6v1lAWIiyy3bf9PNpinpK
FKlCwEa982QgQBeFkKuc47QDrDp54EhZdDGT7jM76kAS+k+wv5W7xtHbp9Ez
XuQ396M4JrbeUGMW8BLlWlxjwnNSFwxeMc4NtX4o9T5T8R/U0buDJQpC8xkT
aaH8zKgJqU0tsNdHQ0Ce8Fp750BU8oPYTy8hWcKto6A3c50OFdH9EsSbyyAU
ToAZ1ticp0LM7s9T1Diwui11OFoQyXqEpE7G+zSUyhh2qsf1+BZwpyZVsjkC
i282XrqN21XvR+fq1qccewsQY9ug3vA5G5illQr7Mtdz2G1k0B6HnpSAQGul
vcoJShGHOTScygWzDxw9Ir4bhLVO1ztPBUUQiGCK6YaEyYCiMCMkEUt23Zvj
Fd+Y9VlEuaM4in3iGlc0zDoDj8r2VdueIjXyZjkaHnZAc/tuATi6tEqTvLYz
8x02szWXfJud6QfPj16RFAAZIUDKQvls5VfAEHjyR3wH56azQ6zlTCtexI+X
2MTxPDN/ShyFj4QVFpGK93XxzL7sCNTVpOy4hbUj1F0apwsuZ/tvbm13jd7D
pRB+DR8fcaGHsbtJ/cuecHBhZkfbDKgOKY4vb7qkyrzQ+i4QfJNqI43hPn8f
hWdOH9jm2lh/C3QxzlhCZNZF0vp/O3stVB637kYdPUbnrmLR+nZ9L7RGLccS
DKbE07pTd3g4VHNii/vRnhUNDOx+mQDylUNuQPJc5yXHfGcJnDCSdZxtd0mr
EQIaD5z5n0lLUegWqL1rsY1ONL4QOTMO0brsCSj4CXWg5uFF7zqEGjZzBr6y
hFWnpHOpdRYBQ1uyoQOmEFZEZmiQ4F35QmyLcOKw0KHCMy5rHJfbWprElW2I
0hivH7YQ5wI8w0GLWtAPtg22ZiZ7dzdvacq8EqC42xI+gcEa2hFLHOC5TpyL
nVN+D58miWRzwVZGEszag6JjJ42K3AhosQ8lhEX0CN4ZOIxMrjp/eflY+qOe
nPbJupLBnrggZsN/kgHvTrwsEdfXa5LQnbI9rTu6O6P77YkWzR/m5b2LuOeW
Z01sCLlEk+6c7ik8VuSG8V+RO4VncTVBiA/MK0jEPv1t1VLLKdZlTj6O+3i9
R6U6p8KJ6LUROowfGbIGbdoCJkdtST9kTomJe7NDxvzjoBbAO8ezk+/dvn1V
aKU7/7zRwAvsSN37SWPuhkZ/avMSHBu17OFLxdpXi39VUGfRZChaW5Qb0UFS
mnR+2EDpuJEM1sAtkr04lLsIqZ1Qv3d7VpxJlfak7Qv+M4kBKm2LjKqKtFT9
5q3OP0l1YKxaY/vbjtuUsyvDwsU2PsGpV/ejgsMe5/P9cluq6UlCkBLVkvRC
GBc/TRMMTjDuyTg6DrMOnHpFCptGgRNVKiuQU9Yr17dBtL01/czMHKBMhoA6
ekeDK46aWAGiTSEoP2Za6ohYA4yYGGPCGfQhyoh4hoAF8Vc3T/CBBfHC8rVI
pGKmhjkgbuLLMKaYzATZsx/q4UWZKe4q1LXS1EtVE0Nv3CX0fjq65uS4U9TD
G03gBFAC9lFqtbJzT9zTgMyldG4VS1/5xDBvTsZPV8LObp0MNIYHULE7FUWK
3g/UTi9Y6vYIJ6JvgpBP8m5LroeQ8atgKEw2V140D2M/xlBfMZZfBMmhq0Wx
NclLGAo5W9rDQnkTO7UvF23ETE1z6drENtA1K8Dx4w+dmt+i2vl8XYtAk88j
54dIoIgLyl/4R7z8WfcIVN4BNbLNFHGUl6KzUOYWv+3Vb0TAZa9jM/FuCp+m
qSlrJR0NJO5g2kJjN3KyMu1flbzVs5Qm2RNzlomFbIJ2czQ/I1/Ybv9Sp47Y
T3Xpr3OAJBsrlNYUtHDFbOPrrUHndJCUZyF5pDe8bBzxLCfiKZa1Vq0LbLzO
TDDheSD4gHOThcv77tmHG89EC0PebwY7+oC3YMJeVVZXghxrDW60XXc2Q8Kg
Llt66oTgQ6efgunAvFrc6CpGsCvBVYF6Zl1ZbyOWqnBKWI/+IpR5RiXBPQ9a
VKWagLg2saPrR5fNM/vIyt4EmrOWmwOsC1jbBNck7qujaNYfhCtcozx+kk9P
cTF9jJLQzzSNZ7gx7nCJ2j74k9MagqEo5mnri3s9iZx2gZS/z/MmWNYy4vQc
jDJ2V1TwCnYzk8u/RW0mhOEVEHyhhZQ8xKncFStXPbFOGJJQGg3IhIT7OfeK
h3Gse6gsPpa3dP4xDUr89zR2WB5+nM8aLCnNfPTntbjcJTd4Ja82OQ8Za1aP
DYaEsgL4wsbJfFFdaZ1tFNIZKfKqUGL2JgxV4Xl9p6luWFM2U0Cvfyi1Hikh
HQhbljvKLF7ExJBQcsXiBoKwxU9MuB1l4klsfRMmlqMcsjGyrYKsqC/fCVqd
yrS+8sCeIPHptA/APpLo1f0DwqsoJh725dBarlCyjbG7L+qnDKj+4qgtM7PT
NaHWfZHh0Rf9euyy8LUduMZ3R3id99kiFVQcptHxy9RBCYzPVIiJvfvengEH
WQRGe11x9UhHV99xmmtujlE1Nin5MzGPXoy14nKJnDPLYiVDDA5qC0CejoyI
Co6kI72MkPpEhf4rhZOXd5C9kC5RhZBr7vUSckyS47i+kwS6kFIrlHMDcnGE
OB0uTGOGGck35IH5QDy5ZBXj/VQHNgICT76SVRNjl2klBy4nY4dvgoRWUg2p
ndMDBkyjNO2pIg9cDfMhayAIWQ5VtrnHm9orQL65P6EVT2vz+5Eror7v2h7P
nc5GsfVO5RrHRompRRpj+rsvDf8c0cOUQFx28gCxuTQ3Yt0XxdrQa4UR8ZZe
36xWSEoKijYT6whodsRL0EU/WBldn71KjDenvNBMmvTgxN9uhJxF/E+RGWo7
7pIm9YKO0Be3xoynZ8ueVqb7KjhjvSH1w41UZ4gzweWh9S5Nb3JY7Xnh9KxX
LN3E0ig7561qFU4LDwQXtc1hn33Ko/bLdP3hsE9DKliJMbyLFwThngdopPWW
D5rD27QjmS0hMDAbA+rQ0OCJAfMJjAZWzgWDu9fjBOBQUjYOAknl/Bx9GRfS
cDcYqqCfD+lQ+QL3VWdkuhg0WxxerWyUuzexQZ83fd8JR/W4g2uw+s2ofPeG
T/D7eTBMutpCabtN/2V09nG099xWE6dCku2SKJCJahivW32/vj/GxFuH/NOd
nq/EjJZUtEtknkeIqwanDiLGdYiiuXqU1PqLyd+f4ChJ4IB1Ck9LlVzA/sX7
tMVd7RyLcsagafhFG/O3aK6g4hv4L5omGj7uBu0BZLSlUwdV2q1FF7N7R4Eo
NqWxBxTF6MBr4kFcimxrBfa6FDEb5yRlcHTvSPSspw6wUP3aikOGdBwf4hOQ
I9hYedSaYJFfq+u1OwpQKBFbumek5hDTx4Vvv2bg7uYmoDQzFKgARKQZNOUg
veRhw9y7eaOkDpkKEZ6NRMd+EuoxMtXLWqivkifDhjasHsPAGlG3wlfnF9ji
UyNwcSNib+AfmfXiHKeI626jVQLPGpxAbkIQD1ZQVX/J0kzlKydjO0QzqLYg
abrOle68Zu+4pPyHdw92Xb+TIPjIbtj7soBgi/b9IjNQQXIyv1Q1Se+Oiqdl
IWZ4JlxCmKE74iFQbFRZ7TKE4EMx4q9y0Aj7VbzToJgdYHQi2l61xsgTd1Ys
V6wfu97BuDGKU8YdAERpVvNTAiWtYHqnQFmPscIqGe0aTB9478tbCOt89rhb
6X1ZRUkxZW5dgyLzRme1toPK8SeWMv1AxyOtvq64FjDQvDhASPZnguYWhkvV
beaQDMDxLFnugtUJnDhfUEm2yYhTmeRSRjUwKINb79Ki7WZy9N0cM+fymJKE
9H/mhFx9rZj+nGBv7fkb2Tmoq42r0CgeIcbzBWPHyz2E479ceT6qMDvwIuhO
Tq637EFc5dIKlc5oiagF3Y8j2lD2bm6h6mzoomBk56uBXiEq38xrA2ioe5K4
AACi0xfEE12vmtqbT78EULFUzMZ+GI8nFwpoxe1055ooU1ng5n/pNQbOCDu7
hOJCjlr2bSJF+bDW5BvGtv7SrUakyo4aAHJdH/mmlxeMWg+04N+jKo7NBg5f
dJfNoto34imojXyfcpq6dhJgpJwM52a367VAm/x2G2vWLuk1Fnrq9X/Ev7O5
IHjfvaf3ixon7nX79ovFGq1Fs+IoBQBiAnM+uorYt5SMEnWi7HYpKlQh43w6
VBcM5ql1D0hLoMVuo0H0priRr9vTb7p8fgx9FS4TDQKOYNHzywtmd4Nd/09Q
coB2bxtY1MDPwfHerw8I52hNxWq1Xu1oLrCDB3JpSVbEvKs5sOiuwEvD6BT/
8chUYLhEr558JlN6KXFNOu5h7X63+6eNWEaJq0GlnYYxiCe1M/IX0VuREVT1
YHbEAoktzXivrL7BaIxS1CYKQo7jnq7jDUWY2G2H9NUkR8AKrqWGsmb78p6p
ZvdCaCIYmmCKJMHk4jhdG+3JFeOgNv1R7gv/0xccR//b8L1KxFsyZmsaJVEZ
uCKNOCvfsNerT7p/BhgeV+m9Hemv93NQbHU7eDQBhGdYGbvFnpl7VZTfUZrL
/PK2u5IwVGZI2xVOtF4+LfWBYRiGequ0PjC+MjCQxFzKMoQ/yHfuSlFAk9+e
XAMWijNfRQXc/YcL0PD2N27tYxaYrykm1mcZ+1ezvJ8q8wz9/24ltcDlWlKN
EBQNi9MQYW3Ig1nhrBGSyaK8n3aE96MCbwdb12nJ4R3yUXbzeQ61/X7tHoMz
/uZ0jR8Qa5esbjrAZ70+2663x5nSEcoBIPhvZ7Z+qur021MVzs2LrhWdD+hJ
w9MBel6cj5eLG0NO80PY6Q528+xWODQjpaO9H8mY8q9YzFHhmYoDFu8U9Ln+
RFZnu7avwG8V3IafKuQDPqzINwbiwmsT9Ya4BAjOjmFNk4w0oXcMnt1V9jmy
MfHCqaFpbPoWr3ENnbuhL0inb9Td2YY4ef9CNEG0u/FAGtV5zpS3CQbikCJa
LbrNTaRKCeualk60IUzNQF8UzShIG5//4rm/PHsVjJqdgZX2SD/N7Fbo33I6
4KFE7rCVvz4fXXagx/Pb8TQFKqD9XiV9GX7NJ4GwuFfs24S1Oq/EYHKZRwrN
N0NXOgAOCeJuUjRnwTQ6F68n7WrtHr40pdkwAaKvk7p2KOX7kJS/5tpp9m8p
nQCbAbaC0SPYTdYCWYyDGL51X+QkEdFuT2/6vXuIgtPMAp6PX9Wgmi3+UFaK
t5l2o8k95Y/SNSyWy/LYxUBeKB+C9hKED7kovGDTVbtRCBsuKRwfYbs5EFAj
xGb2jYVoTT6rI7uG5JJxGjySTQSOFSdiV6iEA27+N/ylY56qN42bMqeEJEvx
GfKjh+Jl5/PD8VQtkHqivsfrSGGSP1M51cVNZP4K8+5ZCFP0ZztJEl4ukgYf
GAWPebXN4vreKfL6jF72+6kK6ZDtMotLRVZQ/u3jsHPndy8UQ0kEXr6RodfR
BkfQJkdCH1DBjpAacL/KnkqdjV/oz3z9hHIbF8FnrhRQVmtqGThDC6/bHCXk
cCXXi2OYb2NNs7185NfR13WDLldD5sKO2DlXjX8TzpYeB57k7D4vzOqpIpyS
m2izmZswy+iN2myCYfuLtNXA5JCCaTMlU6+BRO2oc8l+Ch1elR75ubpFvVWt
Smt5SYWFcKc6LfhgkgyHWf8YgF/+odcj8OLr5G+zdlUEuagDwcInKW7N6XIF
3yteWsUkbY87Izywp45scsMMTNLJt0guYHFF3JxVobZgOEUjWv/CQZf2yqBL
aWAjkRsi3Qi5nupzjNOaCxxVJnU4U3JUKxKAuPY4xk9D8I72oeDxHdSz7TAv
KegId00upmKM8UZIAibgTfLXKZmoxUK4UiWgG6NvAO4c+CltTeNhMovzjkF3
ckw+HEW+xUeACjtUNhlz0+pPJTe+QXg8A8KiOjuDV9Sez/9qAJerxc2RPW9N
EJ7t0+9r2JW6BYm9NcNrsKwM162I6o9Hm04p0ZTsycSX4JE0KL+G0Uuo3IfG
wtsP6Vvf0aw9qOSlCCV+4CZzgr6MJcKmL3It3f+Gdw44BrRRr9TzvuZrNvF2
2hCUmDMzJviEzOJUJwC+Cyro6TpOaLLFsILLzzYAJuOAJFgMhDGVkCRXB8kn
xxAx65rUr2ldR/vIpp4FJwsRCfp+p3ErntMjR6TighNC7ZHvYVu+Twp/V7Gw
Bph0ZS3K/qNFgi2xqeC6ZTrAPm+Dzu6uSK2o+DsX4lPHs0IJ2XscWgCsAVke
CrOwmVSm4EQdwNQMp+gSYonD/rRTt6A7iTW+3H0PMSDPexpd/gbF96gAQ7Lo
DCLmYcTQ+k4tRWDJM3m69RT8N6xXFRLNNM8Gw2LdbW+hrupJpzn65jalvZ/E
m8/4koNOg1i6VWb31snmjckn+5ikiRvItjBC2mhPHAAf0QRr0DwlpmB8ebEN
9MUt+jRyPU/vSthZX+rZeALZuYe4K44fnP0leGDYgaV3yM0d+BxiYXCPaY2+
g12UQp242nFcjsVLwRJYJ4hWpeqy2O6yusuYL0DvpAoEk4Wn2jxTs/Ijke8Q
K+w26a1Q5QuMHDAozVpkDaCwMoWrzgKZLTODsbXaUUgD9OwdUdkcHHTMKWUa
DHOmhrh2qZIn6mjLGMMEw0g3WZswiraDU9fmFFRms6hy87BjHxtkh+EPxezt
gyMO4H5SnJ5z6KhTB9uCyQr4PeOTE6pxC6k4qUsN5a/UoSGQiXUjmeViHq6V
80AzLMy3xXW1AZTtd10vsunf5dWegckxlFDEMIEG9WZo4eTlRCQn/7l7NMsK
qmPdG4uehYrVJpZzKJt8OYB5RBut233CZTHFqq2bBSYchQibrHi1yiiM/qLt
FUdh+ovJc+qTO6vcKDp2hx+ytPL3yrZFKaKTBih1UX1AEHjdXZMPfaOhyDbu
K55mQoYTdwYpz+7Q13NwtTguq7VsVJICjY4s2YMf6lxV98OK/591fTShwo3L
UsJM3C9gQWFHBc+I/NmG04t80uyk93xkURvA1F63MdFG3TJvhg4PX+twtZJd
sq+qfAmd2ClfSgcW5UGTblYWWbG3YNlMnDjWTenEJnzIHrl6Y/gOX4/9+oKg
sz18kJ4H65l9+7CnoLBiaEO4WRpEtbNmjWOeAPtM829+PPldO9eLMJlyv9JZ
3kd/PUne5u8ScuYMQxOV2xF+p4Ie/kzOZRQE9quOsyNTMSXFWTRsvC68g0/N
YiAbZKKF1aj3EmtfFLpcmITTj1jil4PdplQXz1+Jf5KyEfaYF/PLyPsuhqyB
nq9D3fyvbB8m6VU/VN24THxPngEZJdqfO96CpkeWOWb9ptBIRN1U+RXmxRvW
+ccoOkMC8XmyuPe7l3Z+C9uqusQMhVHKp/zHLCdtaMLlAngBk29QxEFbvSIl
5s7IaTcXd6TPlQwdJfqLyN6/StgHLGTgtqJcrk+VBnVT9KeK71iaNOBR/PZl
zAtB/RZUlPz5bXGtD4sSDhuku6EiGo4ptcQUFs68kKgXxae1HKsqBcH+lWtH
V394zGOVbFOnmv/6p9jTcoF+Fcxq6WFqI3sF1p612vIdAUThqIr964RSpIuN
1PkVTUYltrkyufX+njDGsgPXrP4NYEDwy0+jAsX4GkXnuhaTCHsK/VQq5Ntr
vlT73DiOkElAbxznuXaZH9d2ZT9amzdqClogiuuO3qRW6Sm2NWWuY14sEUfa
LD5PXepQE+sUG8Q+RFKHAMY0pAk1TeTbjjLpmzhz36DzaEijp7Icsj8ulg7M
hsjtcnGuGXRJWE9zstzsa9CL4pBqGOhbIqafmKgwFCKJg0Di4kBmHDrB3rF8
V+iNJdRUY2QtbN0UwdVg8Vmjtq0J+kOEFjDFRA6Q5e8UsriImSLKVVVQL7Yl
kPK0iv/qpgyRXnDBSmE7S1q0PeHm/uM4jrDcVo+KO3o5mj6D0eiNTmCksyTf
M7xjePtETaKmvQPA5xJTBl/h9rZGCyeREPjShj0NzVjMC28DfawqyhTlLG8L
42/odWuI/Wpb1Le6rQcljehM1yDZxG9Azif5SL29QyQtknuYLtDMEvJffePA
Kfp+9SnK6UD7rmB8whVvdZfyyeJ+8zrM3FSu8m25vEPTdONtdAQ+LKks6CBm
+8rfcq4NK1QhIqWQEL7uzalpcgicoYJT0OBFrQliV7vctjQbM3YTaBFW84UD
vkpPuVy0ghOQImcDNO9tszwSFZGztt9ZJoDYROEQ7zczz8kWadycG92ddWBa
kdX7WVdZYAy4mCTl5CCREAFXbTkVEb92wP7OagZd4d5K26uORTzP55r6qTvO
e4AOGwt+fBkzuJZIsdxCkUtmPuVxXYR+Mr20eGMoVQJFdY8vsliMQyaVBV1V
XED7UFXGObvB8htTZ/I2pvcM0nJ5Mu558fu51v2U55u/jdhp+CxeUS/3n0Hq
JFP0GBB/MbRDk9ClkQP048UyB2Jy8it56+bOrNHOTuVDj9sApvY933PeEvog
w5dUq6YI6HrrKXXR9I557IBeO6Ae1UukLQSEVsvI7QNrZhB0/CFbrrmFHjuO
xw8FSmvgMs11xVuCi5kTQkIw1sdT2a94cRPCcKlU2SDw90lGNNK4TKgA9BBB
6DAA5jLq6w12i5g0U2pmtnYBwGI74zoNEw2A2tL1BfBS8f9usbz5lsa78zpR
FfPMSiEXHNLWwPB0CweECJbw0BoIox6eP1RbWe/E24wEFrNXrDRQSZSJzWdv
F2sD3NvDEoTZAoQMu8/NtkTG2Q9gZCCWOJJoKSnLI9FOBnm8x81KIgBJbZ7U
/SXwNXNvXEzjC2MRR7Z1sUr0QPTebRdCKeFjTTUhIPDoacb2AULOaPnN9Zbd
F23+g8o/o59+XGTDS4HqQpAflV2bB91OHjr1ygXMmUR1INNYh8i4OxEgGuJL
pzbckav7eY1SbSyK8AGODFvdEmPHhWh7CvxxSyA9JypAUDW2mM9bO2e/RjJe
GRT7KRL3+4PpP7w+oC++k0yVYFDqNtGD+jKLx/lqq8Wdo1Bon4TG1xsRIlGq
qEq3Xkizq3xDxlfg+2R3E2aFgSuxz5weojmP5IEvkWO0iDKCT5aXPqE9AZYq
YMh5VtCdVmJRVqLHvNEZ5sysuf9ScJI0/GvGdExQdedHyqOrl5e3ifwkBk5h
s7/+o+2M1URetP7Du72QwajPdaBu96vGcyq4hSPqzBRKWgUs2V9MMu39AAxM
TCpBCaQR9A4HNrax3qF5fvG3nz2qvkid2AySXifUx5a26BYqIyVE6Zv+B6iC
YMLju9FUmsQPjKJlU1Drkf8jf6vehGh2yWuJKrbnp/tkW+DTd4YqNOyMUrk7
5zj8CJuonq3N7r4Z4ceolew/fF9kynmHDbkoXMwjbPIhoPE+NX9v3cbBWNgr
qAFO+WFSROOOL4XXto4HEtjOK7nJYXDvNLhmcG1AZ80iMp4BZM/cGMLUin2R
U5ngrk6Kgv82oUWkI+flbySAoN3M5Zc21ruMSZPAoo9Fj0eHzUdNekVYSVVX
WeZmzr+6VHvyw/aYkON6FMK7+9v9j9k6zXrLZ4+gF4hskYSy7LaZ1Gms0x0q
rypP86b5cidef+T6whXqNi5UG925H64ud0zRVUeB9wLTkMeRRr67wgyLHOnu
EWMQK0KOM1y85PLqVFUClNsTPkSbDBWD6phlGjr1GrNadr0a80fnIKx9osgr
craqdiNBHwvvIHl1vHsnE9SsnMZl7PWHeUxtDkgSySJek8C9ste06dkQB4hj
9PtT7gmBAWixgZ8os1O/79MZCNwwjjnpEBWFaOgAr8Y7uw/AJwEPrilfdOYQ
3PaBIm8aSpGdS2eOZuJVLHp9a+YKom1+lezV9UPaS82ZSZaNIDufwkqFnG/c
uJaEf1qgHEsMaHRnEqJA8R71r9YDtNGtI8YE3o5ULL79IydUeT7nW9DVQUeH
yieLnm9NdthecQVi4Vp5IAietGf1IdZ7jyLSljnKH3pHoJNfMqVpeEKS5f1o
A9n4sxbpU5WcbpA3z7H/hY34VlXvfDf3ebHFkLWVehryd+ImBOsweBKFnLK7
92zqlg9Mk55F8KpoDVYZ7P4+e1VoM1INLvzftKEUOOGtHIw2tsxqLgV11JkK
omRUBHNqEkGqyJc/4c0XEpZZnk2fRgre19jC/50FoOeQUFsTbR1SWB3LWhXT
xDCoCDXTNybZw9OjKpYOVtIhVvIGQO481UbBrLqEtsKCR6NMOMzkJD13JCvu
y3LWuRglAEG3OH+NSGygi8wAYYbJcnm+/9MD+wHS/PFTt0cl3k3MiUcO8eNN
jykPuMICwANjhrnYxIM/ky/RfXme2RN090DNZjhZ2XOl3iuLoqty8eZakjDN
scBMxl09X+kBdiEZ5itHggvK8wQhAWR5JQQvo7tks1Ta5V+cVUDqSBqAyhM+
JBHxwMgXaTqvVTjsvncgKSblz4LKi48P1txr4mdBJ9ZcvnQTakYK3oNTNnl+
52D6Ku0wZGNYkKj0/MpjW3T8qqzfLaz0nzk1jGP6SKQglS9vN6L/Dtr5+Y8k
rqmW8Yv+5zsMgrnuEgSVpXGRUGa7E+sxrpbBIUJS1D4ycYxEFNq+Jmx1IVd+
XPk7RvcxaF0CtoqmJ4QI5a/nVhHrA6xuJ9RTNH/q7iikJwvwRmd1bbrITOsI
sY9/rvTMnmm+xUKYrbG6f7Jsrcss2w4EiGCo0ThyGKvI9nVikms04A14226a
NHmN9pZ85dYPgNbuG9tbeN57XrCaJUuJ/iltj5/EbHfDe8v9gniwgsiaMpdH
p1uef8ZP+Oy4Te6Mn4H39GZMNqo193LJJa3w2QWwviI30ZbPGchoXoQ0tEi4
yTmhQLlsKCCpa2jeNPL8X67d8Kg7CpkQhxmlrHUhk4gl194bKuY196yvCVFI
lON1HQnEHL7S99jxFZ0qUlDAE3wdn+TB77EuvW35IDnAITIwfVnCARwck895
F7ChXLyoAlaP0L0u2bcRFly9eOtSoyPIFK+4+9fXFbzX11g/7Uk7zo4JW6zw
0sTweMuVJSnSAKsS9OjUt9k/2j2ZyV7ZGBuvVZIMTy1mgbYDY6hPe1IVWCd+
ZeH7UumegXMjrJp1Y2jgXMOY2tK5NIVZaQZRVsJ31p4Vpo9+smszQ9mkCXR5
TZyeeTdbbyzZq/r68FlMLmYEuP3gu7gHsOpkgV6U5HljoUYkhoEpiOMHeNlI
MbxWPIW7r2PiCLZjbDtpctZdVoE/5yN3olxfUQeYZIeuRl2Dr+QjYkAHve0u
i7q6YLaidj1MV8pcB9cEAMwMgRZsHKfvrb9cnC4TSbisLXwXFxPoEZo4OK8E
aPkwEIeBBWWD6OfX6sdBT8G2e3MQgalBEYTBBbp0qebt6y+3ZOrCQWDa166s
BGWmEL5XV9sGexrCvTDR5LPUTHn1tuF6lVBLHhBXVlm60QYx5vIE51zLoEtu
21mk+Ag2UQCjlGQEvdLzId9LolzN9d1mhcYR/tpzopFwQNR0Gj5PzVy75k1F
7gqQZFMLjMhKoKqiSplyc/ZhI43McuEaQtYl8FkBg6A0LZFyDiAp2ib2f8bC
N0dpGx27bn7Gqrx4ni4y4b2faXSIU5M/Ng25TkAstN5UUMdzd0KTa0mV5KK+
jenZW4f8CkO+juLO8uMo8A1XAJSnX8lIizXMpRAKa47z9Io1Mefo10WX+DXL
W3Eu5dwE/3hKbyFrI2dWDIOs/qhyaXmG6Ie9ArQhFT7hqaTTpSqPbCIa8uNs
cEx67mpG8NVetOBC7+BUZ9ewADWJRgj+wOQ62y5ZsjcyTO/nuX/kGgFiVbd4
GJXhQW+wF6wabH1Aeq9z3qAq7NeStQ3tBdxbmiQHczp7NgPtsnuwI8Da8jBF
Ez8MDHehwxbXWsAXvNgjvh4xhr6OR2LneAn7sjN2kea1FgpZJ7UoaOdzOnoL
X+JtnaYkkw2P9HXkBUsLzdoMJEDgEoBa61d0lIXLq6vOHS3kNAtYFs+0phay
pDvwZyi+D6W1rrA2mD43JspwDTwi7y8V1xWYWv7mZwnQe9BEPx9kE6Bj4Le/
zUT9xbzJ5LTx2VXxxLohntk4F1JvV/ETdEKvqJLWL0WPVE03+pfcNx6Htn5o
A1bp1hLKNw1nrH8uP+xq9/OOQvAJmfEBwT6Iq5X4hPzAi0fE3pOwvytKjQeu
irem6S+9QgQlsY8+D/a2OZ6iFShcZvaVls5IFNhZAKE7CVePpms3ERGwEj2a
zsQkanK5DovIOiEdzC9DqlVIek3gf571Ee0Y17wEtkOP/7UXfzlvk87ayFq/
pnrHv/eywcxrJc63NFV5iOE3/hb4kfgv5AGBbHHLYWQD6rm5K0SchNh6nv9h
0QihrJoT1DznVmpNot9TqicI1iExxB+ZRyuN1Vc/P1edSee594cco4girnmS
Gzq4SVhNvS01VSHMZWbmBeNxqy8mSyNHAP9LnpnjYpqR1coyhFlGhKcTX5+u
NBlNBOGEk+MRCt4u9Pf+MV4sqiJJ1zW199aNmgHchjXliKiArrMfX9JGls6I
FtfysTezgGtzNAMzJhTvwq1JPd5fIIQ9LMNAg6TZM404XG+kzQyEf1QnNcJN
q9jqBRSvxEpdIQDr3kO+yoBH7C1VJlHp0qLamdvZLPUdVTc/d4QlSy/Ipmk+
HCSm+LwQ14x/3XChxrAr/2ZFbleuayEgFUPRYWPmsLenBd3k0R8kHeHGjcIK
v7+HaqZZtPpAEd1aHxiTvPUlMyaJpkTq0B+gHYYvOxO4BcgXcLLHVOyVs70t
xcoDYmUiZM/WBSRkSn26+AsKhl/ZGF+fN1CpqcSa3c8kRJEuIX+SwXdqVPrs
ROF/QPQVFLs19PwPhQ2DA6XHLnxPl6c8PIedowAssYMQqkakfUqUJaCyhX6b
uZinXkRBxDxQtM0fhXUwZ9EvRkfLq4ZMozPLKvVRiEf7AD8f5vN47ggP8B2b
psvb5yzOWr24InWIgOTzC6hn9mcQXeeBH1YjyMMe4etw/dyT73ftyOPJE9tC
bWbU02pgyqSijIJzIliPjrtyxKoICmS+adKcyA6BSw2Rk+yJ4pmAbnnUDAux
BCpVoszju2jN51wlVLzTi27YUAHXYIS5uFg1y7+yDaH7URHEdPIaaARWWXXa
M+M9OEElfRm26W1hdl8JphWsGsgaX61mVthio6mrL/2JuKfwGdzPJVQZphR5
9ubSYxN9e9lFtPbY+74xGSw+hVCoZ43sSGhF8Is4Y+ouNeYftGwZxKKrsAgy
s9MZ572YUpiNuqhCaCSJ1Ai6VJdi+2qK5CQ8fuWDsOIAOA2h2titGm9En6/J
yS5YfKLxCE8CW1OggkfGvBNOLClESgz4CHxPWwfvSAQ6E1kotjkJIb7Bf2d7
m2S32t60LniYHf53uk5F2HYZ6NX83LpbjF9ktFGIYC6x1tDuBLWmO+KwAWI5
GUjxIiZkr0p5We6qKv0h4g+nVcMYRgsu7XsGScBLXT5qg3EO85KHrw66dJGP
spAIrfgnPvC4c9l4J1tor3hWeGE+X1FgOCSh113ZnzdFNWIoDjXbqhH5hIQg
CEOJRxMxu2jHya7KIpnscBi7ZD4mzWpYh98Dg0w5tOdSKe8yMbHPxCGI5H4m
D7fXClV2CcRLiLasBzLewERx/EaRhYq1ERjg9EINnV//pfVU6jMHcBoslsi8
+7H1Wruzlc58iltLRkKnuYkO1EDFAfIzeWRZsGndK9W/OObA59awT234vREc
9r2a9H+owRrN6Se4EivLceFStJewO2LRgQR6U9AbESrTauLLlw63siJX+Xfd
pilycROgLS+fCU7Vy6npfJd8WQLIEll4ctgY82YIc7eltWc1diKlOghKjTVa
IMb/m2Xhx5HOHYHbqCe/luViPCdNpcDLJ0RI0VLmHXDVVkmFpGQT28KkN3tW
jVhPmdxXeSurWpb2LrhB9Q33SHbgBpOqCDgtaD9I0O2Y6jIXI7O1m1uRZCLc
GXCzo39o2fuJ0aEDy+hH3lMIYZ9LQB5B2JT5S7fFx1/6ZMnsQ8qYCyjfIWxM
69giMXmwTo+t0TyL31AQEX39xmXk4jJNDvwSn1F3sNogZ2qXXKSbbrZh5EsG
Xb18E64pnhdazUKu9VETSPdP14YmgrTIdRdS4PqPJHteH/QLFhJzsQZJ9xX/
pQniI13/MisXnLWFX53w6T/2ibm3kaMiZ8R1OAJ4J4v7kJ0lWnf3nBDbqBs1
3XZkR5OLf1toFvi9NCUeVVID7d3fzOAHhmnsVIMmX30PEFe8psGMgEzNddms
2zgeMh8Dp/ve5JYJtRdK6huweibYnIJO6T3foTUBMoStD9NKXucL0AJdSd7S
Go8qls8+0vjI7NrKAmfOJZpis9zVFLdZP0SbbUuFgvYJPlU7twWC4NT3xFQD
nR/HWdwyiaswfRd3KwqLeXn/YS6A7RrsoyObeLmh6xgXOUR8UyT9qB0rNklE
D+CqnVr88YlOlpOgMt6lTbEeB8N+wTWS8Dz/AhpIKAtp9WyXD8aEgoPfdphg
ZQ0abxgJ3L/PQvy1QqzSounji9N05fot/AGl/kmEIOlPaYVysw3WSsNcBOcP
wVmhp+Sgd2elQWvWYKQx3fuwcMbWmXdXW2AU3FwQR9QBycSsdDNdvWvHiBTf
lPs7o+7g9bvUjKZFQ50tFrxuMvu8pnHbGdwQlEXU+3d5Je4OEEpHp20TlBJK
LwbIBcHM927ricEnD/5Sw0ANzTF1ELf5DODSrrUDp0PKguhH0wSCZgJDXJzi
Rv6vTFDBoS048TZA2oVeiBlneNneQMuCMfsf+bowfno4uPawbAd2TkBmFw7k
TahA1F+ukdBDBVk+RCmAE6dmgPl4nUxMZN0IOWCFT3dMC+XNTt7YSXw9ltBH
WMlvEsqp3cd3sHJzsG5ViHkLTg5eqAYPKDJF8v2OaPFZtsl9G6NW6WlcXUzn
PFqa1taJ9tw6rjDdL9/ExJKqiywmcqpRCDLvdBg9uH9rsep2aeotObMzoT9y
OfHr2lP4Hbm3wlBneaTqdlSmUIjCUyZ4p4ZAudfNP0NE8/Xj1eKh8MYBGUXl
/nA5vgMyGDBwO2skMoJsXKY3jY+EkfehiHlYReZgipp4yP1AQcyVFvYPLEBZ
6qur5fOsSBnkhUQCzkDKb6HwJd3Er/xgsi4le2LWcqxsmwrXMYR1J5vjbKoY
ozQO/rLg4Dt7qaH5YwFjFHL1zCXxDU9SsjHGz5NsCl/ROw9zI4mxwhrMJoil
eJzwJgiL7Fah8ABSmKNaWvyLRHbZAyZ2nhrn6qddu0hAmwCLm1Q87DgsWhMm
fqDFAWg/v+jmptCC2KrqF+UXAlz+Ampudo9BbqJ7GvCyUsQWufVoXmTn48eI
Yxhxz8gIZkOKlzapWNwQNLbv/1Z0PEGjzAX/vGmqYx5mXTnRqQuByOW+vsKz
6h+PAAm0CwNYYWQ/9xIYToDGTi6rwF0SbPuSbJLymMao1PwbjoJ5GN2oveP1
zA8a7t66blV/FyALpNns5xLqPLb4pnb42XdFb3PdKxYSGcDmziFrmzlg5eoT
d2n4UIe8aGoCPNm8wuoAsvOUSoImjQDG/uHkWMR+RuuH00i9udNkAxtEH0Kn
lVJRkpNKBeVECsVCX0ti+CA2gg/ie3oR1tgOb4K8xVsd+UafIVBU4esxvx6m
hXQHLj+3NENYi+XnRhsF0UpvSGSCF5BpqlRLeeIc+lUm8bg5k1RpApzpgFH8
a9/W5RuQfQwOOODuMjEUmzhZwb1sq9xIVHLVZELz89oT1hNTluFTgsX8VWg0
ZPRfuvxTBdpkMcAWIzZJKBdDHPvN2LbfKEB74d0lYCmZHEgrE/XK2fWRLS+5
a5nIJM8OSnTnlx/egNAIkIiJ2G+UhuVe09gOp7ZKdgGoW0InMxIDSHu016pE
uGWcz/shRiHduDrbgqJTTZXELV0yRRePCK6XEKDCWG8MQQy7Gv29U6bCc+jE
nAUX6jlA8/C/L97m0EksdXTq3RzYedKZv/1cd9al6iMNR4/9SZ7ljUGofGvd
aqYK/l4xEhgvRRMQIrcOxqj3Jp16RCZwW9lTM99T3lFOWnt1q9gPo0jNU1Ag
GSt5OQv88aV/8ChMnj5GxpqvufwVIzBaI7p07lo6j28iOMPeaRvVOXcShQXU
8G9eNaJwBMgc1YBShWjlnvpaKuUSNG08JjY+lVR50zYXVOum5wogNfe8jFzX
UxPrU5onXCKCEMAZV7mokUfRPQpVzvzIKGMSNsJ4w95P0h/KFj9lDIdOkqXN
Vo5bl9Eqf5gcjE9VQDVzrIFbtAewEo9RJv6Mp2KxBNNIzIXD+j6v68V5zoTd
aiTYiBrXTTrUYRaS2I13roN93j/AdQEiwScj7X9Y6pU/LfmajSOBs0SmH/q8
xTxU5Rrv1hfw5z0UnjVbqk75ZHygJSnyIl/s9vRLsk2m0y+8s4eImNA+7qlc
3wvGdSEt3r973TQARZG+qXN9WcGtQbn4o8bKOnJw/4xXb0WZzIm6ISCADYPW
WZinJCruYpY1HrouCz63IV7JuxPpufrf6Vmbxn2/A7tntI2aR825FqCjGgMx
e9Ri54paaEkrXfh6qFLPNeBfgKV7uiiIzFrIYhpV15wZvVmbrXzQA76rSPFd
PEvKz7+3bF2HiKLAzqhefYUJ1610rFhntFZbCAm8xyLWzpmQkVxFesUrIC3b
krW3AQ64Un+CX5s918U3FLbxxBHwH3caLNG0F5FRE2EaSTcBEQhzt8g/DIzc
/HOF/Mt0KA6zfwfL8A2w6Veh9rQbrAOATouHQFCbnNS07HV799AJOUfwQYaQ
xPe0w/pU4xVFJTiCiEQ+U/yuUR8MNh7y6oXbcS9fHI8JptwrCiJj3y06ZWxa
Zxv5ABQAClMMFj8nlZdcRcSDQqAtKFFIv1UOoliOYNWpGzL9uaf68uADBhAx
awi8WC3CyGQ/6jbDQC7lz6Uxxfa5VKflfxkv1JkMo1w+khdb7NKd4tnMWgVB
FQ2yvZgo6poBmqC0TSGTbyKJ/gaw47hPlgQR4YRyGLoAykuHz2qpDDRM3OO7
7qhoYuPJQtEs0gsRhE6hRW2uN0AOfszcpd7dtCZ7T3+Tv+TLkbP83CMvGgxq
13EhG2sAHabNg3dU+vkT22tX4/Qgbr3EjICRqmVZUytBgdcoogQBpYnN7qAx
M6L47qFkqyaim4sTYrFg8O8GYVpXAvq9RR8ABDEAEVN9vfFhrxRLDrOnKBTG
C3aZdvA5Z+nD+MHwSm4O8hupzLu4N9KqHrqiJx9Bae0TqJEB3mcaR8OLjxYR
RyjK6UuTpvV3ei392LiS1X0zo0af6Rg1wdMwslRbHchI1sX39EDx2A7SEwX9
BCsduLn6oXdDxhddEhh0Mprp5w+lgd+wV0Pe0r8d/thIRuYrsF0kKjGlOIlR
vt8/xaqcrmDx/TJbUpWZn5NkNxBvlSKiJJQJk+HEmEOIkq0Cha5dXJq3CTjT
SK6GpvSHUX9Agcmm/YKazVDFiWpQqJ071KGNHpadf6jxWC7MQUxlNKzskQnz
cs4msgVdwdUX8/4cJdBs1sMOpmuA9ngF6MG3m9yvexDcJa3eArZBHZAHfIuc
1afyNTEHmZYuRdsa3nRj0Qu4fFGgXJL6k1STZJSMgzJMuwIZIMU3sH+LGtAC
3fBOXsl6zkdbbYPFAshQ6PqqW4y+sWj8+Z934LIJLswCwi48Db3DNJDKAswL
pFKOcmBcJts2wiRBUIHA22Obbeo3NBUrbwrK2tRA9WcmJO+ur71B/HsTCql5
sMuVYjX0ZioAoSkdA3vsovRVqWk0pT4jxHhNeh+UqgezmSJ57SWnHg/q68h7
E+gMCMGbrb64mjZlRViXHadrFsGbSoq4rNwarhgRVfKO1F6VJUkF7bcz3bcq
YvvlC0+Ds73Qif+7E3owoN9a6ECv7dWGjwTkPkRzYbUfM9xmM5MnHZ5aS7IA
KpQtFv2NXUNJyYpOk+DhGQq455G2jwPOK0YLUZ7vlOMfCq9H/Pvm0pYsrwH3
p+tebfVIaVt/ofrSZUBEqL/G3/JQJBj50YY4WNDaClmumz1E9A2UdaUroPXt
A63rIbH/wLhH0ELoE6HoCQBv6slLd5wrUUL6+K7OSzK7kImB+Gkb1fTAW0ZX
IbLbEPsI0AUcBUGPZBKWck6RQbpTdx4+NnevmHbRNf+GvQDSWCgwVZczZ6vw
RN02rmNug98vpajL0/DHRLvh6J1PV6FKyE1gCmBBuj9Z8OTPD7b4d0vh6js/
vMwGQYo2p6nIBGD4k7T+AcuKnK5DZhYchgzeUbq8ZKDpH0/DIakOKAKz1SvX
PBiPWOSuuquZwjq/OZ4z0sDsUhifjgsJLRtclBn5BPZGXgOW+P+MC8lv7ziw
p8zpu+nIvyJViHa/LWWopwz7Uy/THUgZBwiSJkQQPDZj8HacVHokhnsRsvIC
xhE0X5Y/UNH/dW50xXIkOp4pV4g2LWIBJBdLWXR8KIQjQ/1RnqbprlemysnX
fN8bVja/Y/51kUdRykqHi3mrYw7Wc4s9swhS/MVp7odAoIT+eJXTKJUybnvX
q9y9z1E33krcZYXeoCAKTdNOxmUUoBUiuyeXR7IXQ/2fmJSMQ2TVnHQiJOIl
1PcKi9qer34tNMxIYaDnk2iHmifShE3X/x8fcLUDYYJci00SBKj1nPlDr0WL
gjHxo6r4TBtLTpIwdUuJHYdxui3blhpW2c00hClZLDtZvitZtn9lcv2vG61l
y7Gi8jG86Z4qFMR5JLU4i0LZb7sJj0nbyh1dil6v/SVreuzcL8GWA8fZE2ws
c9R82gHw9I4uzBhr/fQewm9J/HLSzLnTTceB25qYJTrZbpmgFAXAV/2jJfqW
C7odhxQtsrVHdzNjIZ+JJ3DslERyM1oI/aJLUJLRnifmMQ/jsnkH1h1Lfg94
uBGb7jOk0X1/9RPosvRQNpK7e68gJrnYSs6l2HGNUTSJ+m+F217sbNe7hag4
KP0RfuKrIwjhHfGkYPWBcxmYU3+wnwCTJGNwSnzexrTKJet3HM9AzUT1qYy6
WE1EON2FJGXdhQtcXc1CyrF3S8b/3SOYeE0/eaexjYIgt2gZ3KF8gUtONUlI
ZMogvgiQITED1o8PrNYVY5MRu0D2xlozk63U5L4vmA7LbCUOnwHK3QEDS+kk
QOQZqKqVVMyQdeAE3fInXAoq/aV2ifvJGxhaXt1yFiide6beqw95YYbpTMCR
13lOUlAcZ1GnEe+dleU0EZ8/+H1fMqnWlxdqOKf1ab08Y1E/hNHXE3pIfddx
Y9ucgDPhIIgefEWJdJXRq8V1P8SynJLxn4D/3d1nsgPY2pyA46s094X1xAFI
syv1/7UkUUAEZ28xrlkZ1Lq6Q09WzgCFKiaeJ+Jl3E6cBigL9fkQiQH4eYto
KzEv2/8Wqny2F5Baz779JEMGI3NWL5mWsBxPFbkOLYViw5eJK99kd/ljvp/J
tmPQSaY4EY2FCRC7tjNU/MWplizzHrpRYaDXL5tUqBFfT3+nKl5ltGRBHk3r
8ZUJpfO0UgtFsLENCSbs9BfO7ELvxxga3JCH2c7CJA7SOlp/SSpa2OaZXXHR
4oGIJny+SDArAarSgVhvgAPdO7Hk0KSE5FqA//J3lpuGUd3dHu9EAnlHO5o3
aEVH9yapQCwF3cFH25jVxSajP+wYdZ2mPKrNgpzJyYiOlkKq32fqW7QERhGX
9AXBpr0LDBIboWqgvviBXmP+rgXjaEXK9AgVoPbKPx/KDCbcssfxDZlmks6C
qOuIXNq5r6NaAS1LNfY3nUUaKAwSu4cJKX0mwCGMtnpELd5AvrGQJgmKHLqU
8HhqNGfjGVqzpwDCcE069BOYkYV6i43RWOtW2e/Q/MPrit+BSC3oXrgK1prs
xZpE811JhaWHPid55c7GBT8u7nc4YkzKTQ7Z0CW7DBQYMc1Dha04SK635ZBC
T7JSFYG/X0LS6RzrxDN0dffhCAmfCT7lAWn2/2S8NRH8Oeq0wcu4PgyqdmQ2
psql6htw8GSh+voc1g43CTLG/lYxIeO+4tSlxM3BOKvXnns4eMebNwzgbyb7
CWYGjwWQSOOdX7mJu8eLBthj2S2UWZFBFVX6J3bUAUpzZtgqPYlTyH4vO2eQ
yiDJtM8ZYhdzKVeDcjl9T6q+RYq5N7gJxjOYoJtSi42Z23NTVVaWFJezXaLx
dSu2PClhqFIMRHrbX7MK7R11ho8PuqmoaiNSvZRBm12KBLBvTkFhCZzwKDWA
Sh7JTU5ed/ea37BDGxFVE+q8SU2u37RmBHzi6s1px0eHeheF2X7UbyEdCu9n
kcP5K5LJORdzDz2eAj8s3XBk5pEPmvZnle8PmA32S0Q2RUj+Kb59jK8LjOH9
0iY844dN4h5Ht6mJLA6umJL4MCC8xirEYQsezqi+vRLuRXXE1TYKeu1EbX8u
ZD9NWvbryr/OOHirxZNDzgfDvjtjqfl6ZDt+eGqLamLxycj7yVenHAiRRgt0
6Vw5/Iqq5Km1eX+oB9UD11NmnVx5bBDV5Z9yKUY4AqcPjhxpJgaYQOFR0Eju
Os4P8jgXaFHkaC5t7KLR1KV5WbCLtYvFxsbGTZgWCFiEDhcvvWHca/I3eH/j
e8WEPAtC5aZKQ3lMTvC/jHkWkQiMUjOJlfZCf16yKabi72FDHuxjifNzCBJ2
gVY3FQCOcSu0Stvq8njClZjBfwYWvi5N9/93OpwLEwgcF3JUNMvSPmlYBIN/
U+PWw6R6S4xZLfcDJNtvA3mqpdhe2Nq2lxPM/mCrnuxeS8u7OaojLJ+cYtid
T9teUumdZEtSQLQF2yzS16emibwLreD1ePK9ZIxp/cQ1nygRyFs+iBYrjJT5
Lqudv172j7966cjQJ3ainjxyN5Tnw1hBX3qFfwZlI3W5HSVGvp+C6uY18Ccl
VhdIt3QAByuFAezebTGO0F26HjDQrpSXfrLFAb16V7j2C0Q3UQygWi6D8efz
NkDsivIbpQZNhk7s3ZqZ1LCr1VPKCDrQLLZa3VIww9Mw5lYeHxVYXIUrIItd
SmsAoI8wBhGLCCIjsa3JwuOkQn3PhPZ0762Kdetr6obragE3P+NCOCQOnsoQ
fYu22iUXU8+m5iJ729nT5w8goQmK5lolF/OQ/4TXl4jE4Na7ZPymOphzNxhu
gve+ou1qOR5vxDfdE2uSpf3c4PUAe+CePhu6TXgT3OHhEUH7XZQNFy+1Kndt
Mc7Z1sdoQ5vzs15dkpPvqcIEGfOcEZMqpo/AQAtzz5AieU3KvOo9K5loxHA0
z9i1WJ4dECaa3NpkspIlNU914HvPfD+LDI6aTDXlKfiHIxpAKsl7kCrYoado
2WyBHimmqJPjwc2klC+T6braqSsCOo0enmVSV6NV+LjdXfE0sPujtQksZP1Z
uIsV5fE+2T1MYIcWFbXVGv5qWHff60dVAO8kSwXw816rtSf78ju8IiGnElpR
DU+a9uN0c/a57rIXogLrPb1nfqrycbqaKss11S6CMiw0ljFMSWO9rz1PMQe2
jZb+lT7QTUlOwny9wH+Moa7QFI9HOPXOGXPAoqX1RdyzDwMlLmb4rW5bztEB
sNrnqlClsa1QvU1xjFcnzHPbk4reiYmte0JtaqAFnN5VV54wiuL073i3MX7w
5k2mWAV/gC/Htu0nD7wwudfm+XqaOsZ89DAqXLaDnrgBDTWVU3UCJ0vlIL6V
E8VUPA5S9oe0IdBm1x5JAGuUXg/kFYiSDra/QjiQpkIYa0XKJ+hyJUfJdPtJ
uTtjDGihbNJ0Rm94gM/AzDnk0rjRMXX/GbBkD9gbIa7uLTbSwKLqw09qRdpG
8416uY7brWtppgHQwQ3E743qYztgX281wlKe7iwJr6vHnmQFnUv5HN1LzRe1
8GnCug+VVVq3R3dPmx9YQQ/Qi5ledZnk+mFecvITwH5q2cIf2u4ZcxR6s2A3
hsxevcngjZdIt2gYufP/x+6XDiDngGLUiBDbG0dZ2BHWR6g8tv0vJoeMMOzY
5VayrCxXBOHgEIUeaaaDHdD/jxNwni450uoubPnmn5gHX6BIpx7RLNYLMTtR
tHRO0piAVMpMq78uJBefV0+UAq5l5NMWy/L5QyO/U//vA3ra7BHT3zqrduT4
GdK9Od5Nmu5n5icf7zUgP1VWy4oOP0MYpBAWaNHTdD/JXUEw0Q1jRF3XA5Jk
y2KkYo+ynAS43oCT+xO6jLdGViUxrW1BFEKKu0FB5NM76jWKETfKX2QhMlZK
mY7EnArSIHEs4om69U6YpPR0pMMwVKaarqc3DOmorSLp0NG7g0X3iqsI+tDI
uwp5QBV3J2nhWkCW2RDydlz/G1zteE3g3MPrvPVOcHDB16xeGbHPiOv5zTWi
K0aVl3WowW5SHfwCy8gkhhqRP3Q/UePnYXTWYWqvvPaw8rMhnTBe7TT4yJcr
BZOc80+JUGWm9LKb4aNYTQhPa+Y+tYlFsyKP1zwDr7e1nl7Yye7tdP7yKudE
gDuUZr48R9TT+qk/A2MQ7ARSyAxGzS6BBNY4LdWMynfXhheuMvuFQ4W+DuBr
yId9Rz97uH2gtgU2NIzI8dH8TohGD27ZXKqgN1ii6ICtJycl1XORkbQQiJwN
VhF5EBLLiaS28XNTlByXYHHbtX95kM0GGkeoHHKz0jIBiwtlRiw1MWI4HC8R
+WmdhmJQJxy/nVd5Ns2pAH2gVgrhizw7tIBoS9qBlD8p+xlk3NsoXO24wrEQ
fIx+CgxZF2TkT4HilkOAfxPaQUnmDPuOI+FkJlCve8raVHXcXN+ZEt49n/RU
22qCuXlgpa2X5gMvMXJlpo8+cLsuc1ut2WAChaAAro9UD1LcnU0UjjC1ccH+
pa7DZR8oZTXF74/uplO1KJp77nHc2yNQvENQSBlcBzHMbiKfywTebNnEoiW1
fiKN4am4wmcFDVHB0eiHPBTIV3317oKjm6+IYcqyR6/Ghy17HSg+iBxVH2rx
7Hd0hkQlQh+luIj6rXYo7xA8PHFnUHY/oTQY5uEB4kI0pbdF+unAkL8yFZ1A
C6rgp9FyMnbf6b8VTa0R7lKqJsmlerTstmBch8wlfK2NZH8HEdixjYX+D6UG
lxoyFTzryTzsq6ZiIlaAgtk/tGMnHOIPB5q6ff966qWqu1mLR1rUTlzK31Ii
SWmEFatifGUyUiaASSzFR6RifOxp2FfgOEQNTCMGeML1VirKHqUpwl1LzaEy
SBSzABAdzSjCcGeN/4b+Zm+vCitIm3GnuUm+mYeP3M+wXVhSL+a3CJQSOufZ
gfIL11f1NQX1xWiWFPd99Hp+h7kmmQTHM7FAd/V21BQ2um4OK1zWRSTHifuD
9cuGrcSuBtL4MHIdL9/Gt5pfToN0MECo+JaI8DefrZF2CL/VVUdpDSD1qPyE
7rB8imH+6igsKWiy7Acw1TDulXtN2N9nEU27Wa03vNHD2qUCN2LI5NHXb98U
UHiijauSapJdjvOJjKwqsz8VbYFKDSpERzDVzcF+ju6DgQkiKs2imqA/vjHs
vwaCUnIjh5zhroKdWZN3BDalfn6ATou7OovC2JXsUDjUXocN6Pqt1AgogAGh
fZ8WYIhmaspE1unBljdyiJaJ7WUtYW4CLgTNogyStYyalgYK0iDsPDq1Z0tN
ZXQyMGkl2afC6yKNXFZPIXZ5vJ9XhyF7lA2AFId1AMpAAs+KbJMSqNZLxoj1
vz9c2A/sNlEv1GLKylRnS422eWB2MqeOKw1Uqbz4td3G4+ilcxmSW/8Tr+Pl
EClsLxuv4Kz/X169Umc2pTRbaOwW4NTw0IGMlXsxmQSuymwccvB/GoHF1baI
6GpZqAvJb2NnWCdgii2uoQ+H1F4jtBYPNBUsufH6nw53Zo+M0Qxtn361jC7s
dFKiyvGBghkFTW3jGiIwYViYgtqkAbxP/DmS9xBBBp0ewb/5P3l1yF2BM6NW
3+yO7PUfaYbWy3KloTr1zVHX3V7yyqWavwwBz34oR2R2igsyY44I0GU25YBs
jdJ71N/PjTPURppWfc8NsyOEYEV7A41D/WJt7pFcEGIonmgUZRRjAk+IY9xd
qOy/LKswsXmkP/aB72yx3OlQwjeQQfXTp2Wykbm884rA7pyu4zlnHn6NjhBX
tuUblNOEA7g2k9WJKrbyPMkypUz5Op1j63QmXLxSpwlZ9ZhnOex9qbw9HZIj
ubhGrMjTlWaGu0ZnZ2r9n2HECBg0k49AtEEGbLNBS/2m6J1Qq5JN3FBwE1TZ
plH/38AfJkMBoOU3QiniwDD9hLhEXxWbXRd87Z6I/BcQPcQKHXkDYWCdtMqz
eOHITyfpTBHebzEZ53ygCzyUoVpASz3rbhcfq6ZUtVkFJyy+vWIZXGVbdXZf
pXPQ3ME6DgQsEOO1/yfpwAOYr0xm6IUjYWMXkdrK+/7vTR4pHts1/eSzEspk
HcqdE+tV7fwFzXqoPezcj1Sk+PBQnjsLzJZIGJ5kKP3buE4mdz0jKUp4zwWo
/GCg+MR+xiJaplyevwkONgnkCYcEtXXvXsHSACTOVak0kfYrixZ0GMBEzRjn
3f2Y8B/9MYo+2GI/tfYEBywd0BK+znGRxMVzyzGUdgqj9STcQt/N4mqbZARH
AQVZ51RvXInIcvHlT7W9v5fQDFSRpODMLLt9M6fcVMNTnRk8MrQXBNoWef3a
tZHwC/2uAe1f6Bn/IWB3AnVQhLMUVpy2Sx11j9pxzDno9DUzX19VV+KaIUq9
ddyTDgfCvSjoC2ifKT2md7Tw1r2L4fJk4xY4Of74GmCgbaGH9MBmZ7auH18L
n6GrZSHFObQqQA/uHPDm5uDXmyrhh2gL7kicOb06zNyYCpruAsP6CASo3+Rs
pqqut7Mkf8fLeKbAphDCHFIaYHc2yJzjrkLLtTG1auMmlSpy3PjKCBhaIMys
akqUqrBquDlD/r/OwRAEMqNz/zHtO3QeK5E5zLyc4n7uYfQBGBsghdzq3MOO
Gdjvoe7Rc03hnOnt8Bdpon/Y7584sKQVSJzTThaTql3Enx9p7rUjF4Agarub
gi6Ne1sTMiOS3szdM6yMUOvRg1wBH7hO2Kkxixkz/0T4EGxM+CvAk80w6OQ8
+l/5bM5K4fzA8Si7OH2kGtcj0sUx8iK88IyIST91ToQBrvSJPRk5cJRftM5Z
Zt0XjA2KKuJmfYtR0Cckf2BtFRkAP6rhhT+peTE3xL8ozdGMamskHZ59k80m
5nL6wYGlt+4PVu9NEK0rAO52RAAY5l0PvkbYcOEt/Szl+6hMturVphVIQ/FU
ff+sTxCTBimaP+75vvYRja6AFm71QVKfRDnu1Bno7vHZUqHc6FKVJcEy9nK4
212MtVTkWB7AsTGlu5S3VC61Lzg/NA3DybfNnkZY3r4cOLgdWi+R1G8i9fd/
o7S5LkDElA3LAqTGKWisq7DrKD5LvTkIQJ0cEDxq46yz//9gA+Y6UFJwWS17
SHW5KZ/t1vmkB4t0PBOX14qiz6H8zIH3tjmCMHziAlfUU2lPl6nh50UHy5EH
kma4uDakFv1jz/KdRfaqzC1PWkr0inbE9fLt6w1tVGCL1gcBSBX9zCnQxYIP
XPUoptab7xS89BFjdmF6Wy4OhKaNtEAUGT2SXQwCY+tNN8MLl4dOUJCHSTB/
zs0NaunCpB0LWvqZa7L4gihhJDxUpCNp+Cp9mvpq9TGRsBrmyQfXIcCklZu3
uKpo6/4bEfKLYI6j3Z3TmA7MzRSRx/MC7ZGXhxdkthiSSV91NdHE1EumEqxo
aJvVk2QDnmzqdYsVp31BytLsrrqhSKC7Ute4CMbH+FOyadY2FtI1VdEFK2nV
UL/nXHu9Y3F5HTcx1zVW6rhGmlII0XH5Y1WelO8Gs6c1Tu89IVo7936qoPnu
VheUiVegNohvIgeHqk2e/1A3Nac1EmmvUvvP/Uc5qieqfatmAlwya9FBs6wm
5BpO1OB2mUsaGGR9B8otynGDbbMhCh69HS22RX093dyHqA7ElBpUZcY0IMrI
qOw/faYMcrmCoDIcYgCPdnOZgIzGAASVPpNkY1q49tt1PaSRlxUHCK2n3782
EZwqgSL5RQQ9XvnSUNdKsorhT9bBY1ZqxP0PDkO9XCaTABi0vBCQ8JGq0ePV
pAqtlEfU3wyEeIy6cD4LRxA+QliXz/InjpHx2FsSkKVH8JXl8gN4V2BqkV9x
Hbj5pA8Th9/dOZxbOd1hQiNwS9Ply/b+xD0dJDvgmYbIUFVuHsHYg4IfBT7O
ooI/TfFyZlDpOjcqTDxzSkQUT5VA7BxTHlh/I6GvejLZi/+HpjTzX2+M4UTv
vk5W6KtLA4/5iOO6eriUl7wymAzHMobPImjUpLqtYnew0weUVKcHj0aTR+ra
fXJYtoS+Z5sMvffLITRlLiQyZXwh1gc7E85em0iTZ/yUO4YfHWxWH+1csm9M
pwmGJzsuJF/Jkdys5T1L36XvQg3Q4CmVb1IurjS9Oz6Ggbzk6ME0IqlEv5Ir
TvrImP+jpnVEYwol0vqQc+Fjh1v+zPuyngPfMv+ScDkfq6PExyVSKhqt5tSe
7l8mGI2yrXEW5jQCbcUIJdqSO5Gjo18JZnGmgM478T5riLp1NVoRuZ013Xe9
92SX+M5XvlAcQ3GydyEk6sQEOtxbgT0NS1cUOEGSNWNV0WtABo17Csj36/c/
FgAalLdPgdsC6geuEp9ElFirHTGtTuFNRGYuQw+bvjEFrd6pTlSiSv5V1nij
4Lah8SfB7g/5CsBneogtEOv1DGzA57P4YKNo4GrItluz6NkDed9v6A1SCHId
ueB2En8VpDye8vYrgcCmDvJtTTkO67R+iFffl8Z/BnkANk8FgN4v7XqI/XPH
js8Wovf6OaTzKTSQcfaJKYFDEuoRlCkVuVExEfUPOWpJPdU65DjgGpxWNMta
PYGAEtHMLu9C9CssX5nbauPdhm5/xYgOGGks68zfwBEDq0cG4vjReuzkqPAZ
ziSFVO09DzeNbR6lJ/C8lTAF0HrbfoNEL/I9TNWLw24TpfN3XI2PnhvTWh7L
P/qv7w8zt58Fsueu78S9rKZuSvHAUfzMwtY1QO41EAib1sUDeL24ly/I/Syh
kvkld9pLVaXs4t9dxJaMuKXwJfbOQXjGSRy4Z4dV3YMsXOWanJKpHzs/nie6
gu4NbZ6gLjaDQiaNqPvQvGzPRdCZJIW5cnL1HhUaX2Lx3NpMBG9qYolhQ7ME
zH6dgO6RNuCEYplEgZ5JDFjPbCt+AiqwvxiRewsCqW0PjWqFeXDWer45LXYG
gdvn+GXQr4VkUVQS5QGib416KrR4y7p3LfGjr6VhMX2tz7CEcjjwRKlvRgkg
47NYLL9o8PvIKYRkDUP+UWGkm4bUtQc/BB23xbFe5BIHUVqEpH92peBtO47P
XszF80EWKp6VK41l8KMVFRDJ353D277NKdTLZ0TVe8VhTfYJjhwYY344WHmv
RPSs3n7kzk6DaTXp3g/6kYSGyraVFo5CKr7VR5XV52isqSJUMmWxrqatyi1D
rQg7GNjyf9360TNMRBGzuCMSK3dhBpRaQgsikYMTdSSgCZ/v3XtHiHZj+3M1
CGzSDYJ2zFJYMYCY6WLkovr4DQBp1rcNPGsM9bQe1nxnbzAZI7fDGkO2x9m2
Bb/wx/LNDWoJnwsjSOaw1QmSOvZ3jUPE20hmYgoWSXuGhOMt+sNQ4gFZRwEb
PeHVUZQy0YvnuMuakxfLgnpErHpsui7hE6sO8zDQ3spY9Zb60BWjmuO2bkIz
GSVfM15VfuYX3MTRf7f3qK11QeaArlEUGvtCHglY+rLkWels26D/5ToJ7DnW
R+4okAO7l5HjTsMygelWNqLGWEl9vqL5nx1UZmEHVcPYdki7LlfeWtCoNovO
h3H7Jd7TKFyEjAO2930/+vizdtbKn8fBOE/pKmRPv42+cwbMWAyCIPTXJkrq
CHmfucyuv8g8AZA8C7+1MtJrYHzHe0CBafnxqssFoNnlGZNDBhVaBsaAGGXq
l/v4fomJc7uBHV4Ph9fxAa4cO9jl4JNxuwVDd/edrMB8Ae+T9bBWzF5sn568
ReEFNS92sXISU3CZKuaKPGhA3Otq51ORGY6TAIp+wz0zeVFx6hPPezCjybQ0
JQJHkcrSzFqEcpI0SETT3uj3cKodvpL/3LFKqiSgnCFOYMns7G/C+tR9EvvV
/YncacJmg4HWeZ9LTJRv0PnQh/Tyi+7CtLjVJxUgaRkZR+V1EaJ7ViV96AXg
4zhxZq1IIrbRCpaHDoiJeZfvxj5g7hdjvHt5ytrtLjAVL8x1fFllxdsL6aY5
QsF1bdbI2L0nGbYW7QIm1FU2Io+R/dgbtb0nG6oM+prbCOVgsxTwgM9tIogt
EmSY7xXbdYJ9UnZAf/armdLzCjPYo/wlSo9ftr1MWzwM5FKa5oxkyUepnub3
QdNEfgh54fa7F/t7/DfhppWQYxfGtoGXBqev58dA7n6fM0MTlEDUw6p0JaB7
tGmOnpNsZH9oGKOKfdPxgcfoihmZlj85R4RyMVc3oXcr30V8h2z56Hup+hi/
yxjdra9664S45LNF8hqMY/4KDym36zZSlYwUAVfavq0iJ3rheDSq7XIPHWft
35/vFeVZCYSj6koSD0dFiMUOzMNWScseg21PGH4qFEdveVJG5irWDESb7Osj
OBGUTiOkCBV1/tR6UbQqF0dp9LCj646T3QoFDKJvwPpxelKBQVLPVH+naw3f
itHEHShABU3XLvpeyGYEBcABCQPY3FhykbMArSv7NoiQgMmYVH4ZigT2LCzf
WTeVmQrlSQCtMl7Pi4mcMBoNAwLG/tUgZ7bgSji8qwS1rb+lmKn1tQQtnLW7
gVrYDcPSzIs1FtwRxozyA1yamH1KlZAZ97tAdDjUj6bzrKJqBY55XECf1SD4
V5/y1+uxNVeeNrz9qn4qtFakiBJ1XskxzBGVvJzRw1XQG1pFCQzSb4p5fryj
2FKKui2yxoOIT6RhnR+7zuEcAXq8tA6ihcuxbNBN0TjCbqXSSkAppg4rK74N
3y/e0evyITQ6vlVIZuQBchEyJr+dYI40U4sSD6EZZwDKgZcE/8BYVS7dMAu/
LBZRouSUcRQ7esurPDyrAKsn2dOU+YmvaG5xEkigZKqGSvWauMNGI3IeH/uI
XjVrWaExsWEVYhjPy1AMzlCtQlp5F/J0aXhuBJOiiz3zSNWVJhJHwL6yiW68
auje2usPDjZwHV1GNWNhWq+Zce1Sa5dOyN0gGn4ml4PtZJ123ZHmkjhdTH0k
ja6A7vv/a/J4gc4TaoXXNSY77bgCdkZ/kUf84bzgfXDY3lINKpdKbZa/VKA/
51Q5rJdQIVdvvDLG2BuGlH1gblQbG8TynOg9VXIQnuTJvMj1DbuGaVEw1bh5
j+MD3X9lhKQHP/2Hng//7wncQQh6B6ROPEhF2sCruwPXC+PxYMc6lpXoCcRq
lE55TzTgqM+cAf4wG8ljcWMIBVOnbzDm4PaIQfFBUWpaE0Yrqn+ROgPiTDBT
JcfSZXoKyo1L/1KQS1fo3Wt9Djwri/mUGlmP0/uXxv2l/oxe+rcpqtMT4Z8Q
4ps+k+umyeAG3l8hfrtT4pDEdD4HY6YAbSslPuF1Y7sGatXHIY+EliTRayYl
EUZ98OXAVpMfOr3IAtRuVb2Ya4lZsq99lfA0Up3Fveqwm+ZT4JOQ9/ELoFdB
GVmiIA3sc1afkG9tKP5k441PdNsmnubSZfViPy1zGS7BktA0HKw4yK922U3r
1+S9V4r//CageDWbM4zvpbOB3dF5/ShQwwcooPKyHYDYv+1lzVlMWZIaLFnM
onlxWcPrEQcelK84nWDWaKIJjfHKtjaTJpQUSlueMt5n9uIFJJpL0hnFFp10
gv9KrxiKtsfx0S5ykQTFzVHEf7CBBdPNjnpCy4Acr+liUDEZYyiIZGm1nnIo
yJKIXy+0sQvpAMw7EtaEsXXP2Ewd0Q31UM3M9urv/sCBIZqdOiEj5Hx9+jh3
cv/Lk0IC5faMLGHZCzqO+OJESiZ/HCANUe21wiicMZFFvZbSdr12/8dBzY5B
UJTG5WzQHZGvHi0IsGhSyEsVS+pG4tdRzuYsL2RPb2hHOrB8WJtzCraklp6o
D0t7cZSDW6QjpTH6yBGFzNOsPnfq5mh+K4vQqGlvp9MA8sj7r7yVkN8jLub/
vEVU8M/PEksBwELDUFkePhgoUqiQRtrC497BDNog++whtZk1meKbIswqgddq
0GgDW650tPjxhvrPSA6U1a4SI2aLGsrs1k7WdgiDFwmhZtCGZq5nVFoBAmdW
JGqkzg4bKYuI6d4vIDnHLoRJFaUZbj9RvN23AXrP5yMmj7Ac4Tcw52NJLELN
y7saPxkAnSDLSsQtmE3z0XAY/fD1KW0sSBd+jVcKjbWFWINnElwRtKXFhEpZ
euYHegonBMKlJ3Why256vajCBicb77Fi+9loF3OO9FT6PC66RBq6fajlxVKx
DqsV4ZfSF02o6X3d32mcXnjvoQMsmp0svQO1T+gXBtVCDbLEJYU9OmHzxNgv
ZPYXHlnC1bvi0DR3nuKwJWedugka1qQo5H7BTTCJ7WOlCyp4Fm99eiwMQI2B
PFk19atigcDG+zvgtISLZcR8kSFwtYdFSPWnv+rmFzEsBF0fdiHDsrYD+ieE
YoOZB1AKg33+MOc1YVw2L7eh8cvNisKXJIZUP554UdMyj5EYUUbZcR2mXVmH
ZEZHHxRqe262hmt/Ql3VkOlF5xhG1u/ZuPgfqFcGWRfuFORdiz86MUthHLCs
TxKtv83wXQGdBDjGK1radNeI6Zr4qu1hnaSXV3Rb8npiZ7DFvJSkhiU3V99F
0nwQ2B4Fx3JF+fG63TKQ6syASG0gw/2jAGH46kNqiZ+3TyEV2ExBIc+3zBtw
E/5nuK37jZ99QKBFDmJRqUE1Wzt0PUeZXXrvV0jtZ2VlDpqPHUwvVSYFxQ8a
m2+XrRB4EmhhsvRBxyaTa60Twh8gT/gWvUx5YhKeDDSs/OYUoRqdZlSPRHp0
vd60mW0D1zEUKBumRERZIC8VytRwMTpqCfM0vvynC1RPrsikM4qggOTviihN
88rw0tOHoBaw9jT3WkqoyE6yMHtYi5q+ummO9wPH0wfKXqHSwXGF8oQHtmMx
KCty/L0jHgQX0dduy2uUk+KUEki19d4cQaNO86vdafOR0C0daRrmDOGEZhUO
ps2/JnK6CH0rFVh+1rgvqKNnfKc6paN+eGc/z5fEjZ6O0CPVt/PilnJEOH0g
Ck5L3hxSIe57AlTbxQeRU3w7uO9E2dogPdzumr2rk2rW3t6VpIl5Mt7QIed9
WTrMPJ0GmRzWo4nNfI8/8gIAwmNcZNGoDn4zJLWQo7yFqn5KFtUmfZRJOrxg
zhelB9v8rKpH3ho17B9VsjBPJRXing3nOj6RAtqtLwNgJv5bC7fRZQA1mEA5
ebGqFSu2eLsAzqESu1Ib88jxruVZ7z/PbSTN8ftTZqP/pxBxgb02uvZNKnot
UXhV0xZEs22ir8n74rQMbQF1umDcXUOuNQ5GrZXs9aywktvey1tA/xLwJ590
h0qIBl0+QKh2H6tYX61Kad+9FW+lqe/F5w9JFfPLUGHC83JgdseqXDQiA1Qu
RwgVBe+wD/zNdFG+LlcSUs8fdilDvmw5E7PEpLYHLXYU6KJ8RO0AXzzz82JE
fRueGzD/APz1Hk3Odi1F5nQJtYXPkaQYRRvdOWTiU1PnPjZoQF8Lz79G56Zh
9ZkvOOcbL30q/28osqP7yZelOpYObUOVFMbgV5oxFCEsYpdpKYOqidifsXJ2
oczy2D5Xl5kh8lFkxl9oHxkKcEAeJGpWBddV83y7IhGJqfUoS1ftDD1foWmM
m/4xPJsipKxtFmWS3mYrncAOocuuuS2RXgJ5mPjCAHUjj+vyp/wp+i3bI5Db
yQcZm00dbQP2rAoMm4Is1r33VGXSMk431ldvhylIc+sfU+68nh7j6AZxo273
gY8XHkwGKGHNCxyGlrVQkZxbEXsP2fIMUucv17WRpfKn6EFHzsPi7j/X8+Qf
op5h5Kkk5bRscdgr/zZzvag3ewvPoOp/T0c6Tv8faJ6gDKU5eiVbu2uWXOWT
vQaSWMB0okajGH31C3aY5uQtd57/M6ScK71g5yPPikD10JSoiRbbPgq/zHLe
K873orlswUkXGDbO678hwrUlX6MXAhu6cuhoCvh6yGbu6toyC2uOA3jgkq4u
Xl3IC/af/z8rfuBMRhZG+706YIsRdPP15t8tZw4skrw9GUhf6mC9FKZyXfvB
nA017xpgWgjA773i3toui2au/AGsWYHmEA4IXOEHjJ/3Xty4IdnjE024noKw
tWIlI1gCyBhdj7Je+qAlD4Ka9Z0c6zxN7zBO9jPCNgPH3/G4qiu3MisvCdh1
+8Gtk78OpkEmRUjHjeMxOzR0eDlBkA89arxJHeviM6/z7ltHaTEvc5kgjahM
oO1FPtig/iB5A3UuhJYcFXKjtHzbM7vymhDQQU3pgC7E1SzFF1wia+ZX2HGG
n9NbuncOjpC6FZHWqSlT0DvXHqg7/s3U2LkEDwlTT8ivYguDfKv/k0DV+WgN
sde3O/QexhZ+WUBjKDEqbO1JggZ6Ir+j0yUHN5Q+l79M9sPTpo392r7T93vf
Ohvv4wS5nyn4nHCF6NFxZdR6OjkDJIbBLtadEpxeH40HVySWtTkdDoEXMDxW
sJcp6kvuAkMJRjskXf52mn8VEk8Q6j/hZJ2dSG+pXoY8e18sYxXadhFGPdib
dCq+WZlPL6JonwTzUkXAUXeBbfqVFUO8EwnZdQIWZe2DqMP6EC1tvOWprrcJ
xAsPDxtOaTgtNtgyRrHYl2Ayy8DuuEkGUHq7t4GduSGkS+lzAQqglqP3B18H
fDMD/reoRPay3ghzwgNqOD7Y9T7qDexvo6MKfxmsZEV2tDMIA9rqGfm3z3tY
kZlwHl74zGPLe8pdZiZt+0j7UE9Bk8PEj3mOyssz1AL8q7GkhnRXB/MnQmrz
o7Aruw7pzava+WwDEj+9QcynjAr0xcVmnRBmG1B7aZtXAZ4kwBFBJNF1NpCD
N/jgVujcuxfxCrk0wCVVfXHgGGu9xN0NFQ31gBl3TYD4I8QqUYbjdOVWvtpg
LMSa5ZXKHsPp4+/36mDBwH+bYWQhfF//eby4GxkbnrecvdPduNkb3ylHg0LN
dBfx/4km48Ba5gUdfTGW54wl2UNKiwjgBHbhNtGbj+D4nt12ifjBL9eIJxfu
ytWDcG0Cn4g2YiH9dte4BB0DKL9JodJbpzC465KvvIDdLE9q3E8m8qikfC0t
Mbndwc3ujwr1DHKdpR9HsXdiqwtEM8vZi7acYENl8ZiQyEskRxLEm3VmmA2h
Uzhrl/fIPUSnoeI94cG9Rcq60W2vAK3Vst75C5xcOKeDGisr6sc1nxJzVsX7
VbYD1H6sRUk6LUoAjHERmzCr9Chyt55iE/6GIOCI2hT5A0ubMaDKgw+yOqZC
4qANuTB3fUqdS8VrLCiDI7fNSWMi2ZUF+vC4JGpEmrWwtxuLT7QsZt7hQhBJ
9kPOCTRg2wqQxJvqdsEKj+fSmjkqN4NYxMG5edEGmcHQhzcYdCmZFjJqL+o0
UHC4eaaHJfXGOzwgdS/whiD25aE6yLZ7fp6ucLp4xuHpedWsNXaVW+7STUJ0
YD5Jz11Yb/vAMDpCfvT7EqWb8VGiw+/2OEav46k5Z22K9Fp14hh6YBgw8x3a
Ka7IWWZ+QHZYqA5bwkGDarF5sbiMm6a12dCJbFm+ixKP0olSJGgvfzeF+VNA
7C7vrD1kAP5gYY0ILMBHqupcgsolDprPSIlizTHKOrA7ukLs4nx8EUEQk6ZT
+hEsusvQfhXMZcohRBDQTbWv0gU0MnWwBmuiiJP8hP+6QA0HnAz7DiI0Xr+L
iihHsPWbvJ+wWXW0xr0cItaHh855B+aWNTlWjvnYoLM5Z9WYDfjquWJEQ0LK
sNgDnciEi+FQibt92UgXcIP6Gywroz1ZRgQz3Q23vOfrjYylvc+4SjVnyJwl
z9ag2kSrJ5p86shHUrxN4zKkjKIEsQLHmMbfeSZVRhjjHD8kwDvxjDVbgvGn
4uo38RK0YHtt6MFXKPuH+4yOhTos4yG2LG+9rTjAxlSBhCU8cHe06Xnn7aBU
7qYpBN3vR/mhoQmFDo+MRDFxaTsyljaWTbnbl91826w4SyHGcxDmkiauzX0K
7hZPnDav4qoQle2XILpNrnccJfBxSzquk9WtQsdw/fJ6wP7Z+4BLFndc+X7U
0LXAqqp/wlt8Z63ZKGUfLsH0QB2/EdcMj4z2+inPySNPBG9fSPTT4WzHaIH3
nUtaLEj5q6vyOxSOpCzDW10iFPczOo1idOYXmybZLqV3H+OMctyh7LT40BS/
ct90cOhimwC0DCUITTzOR692dwXb0/mPDkimJTFnaJy2y+5ZJgPcJoNT2GTG
FofBxFSej5xijToBIW+ZzYKZXpsqbT7ruM6TBFFp/g+TuLsfj7tE13o5afKn
Fx2g6Q6N7w8sq1qM61fPptdgZsLIwVyoBej961cE1eRRWAJO9n1mEvVP/JO5
2vbukitCtBStsEFoYbnyR31zzkQBru+iTp0NcXXT5UwVU0UTH9Z9KUTCRJje
NadnJ1LEJ4rLa7kai8tz9HbUgNYx4aZPx0FnChMdV/K7cmbN5MhTgcLff/ZY
VIyGkQZAlL63w3lsj+4K0yOQ9cXOTqLHpziN5jnP+35HyQXemnH5chLzXz6L
W9rSO3PkIf2TiLUTHpptMXiCgb0pFPyCiPhNpUOgz740h8ORLPbWv3G05kfZ
gxcidBOPYzZta/TclDZpEecOBNi48CT+bAKAw9mCQs/1nlJ6RjqHLiq6zDxA
hP+Gs2BaofJpP0iBMhLTG8LvDgosJ2nwbp8uhQ6btvcUil4Zu/SA3XYYJFUO
dHXo+sLgtin2A/fU55fxt1tCR5qhcbELMivyjHTyeOyqcETtILlRNkaWi7lR
2hrNHN64jzYd6QC+a9vQ1ddYfx6Ix2E2K0lMoE/nJthGaUjwBNiY9+p+4cB8
zLVYc6uRJY2Kl5Bsw/X7ESk1dwfmyPJQLQttT+GrWXBuo6IV+NzFHN+O10HM
vayEqoAqjAOqIkWW+8pzpHUNKKDjHFTDQIZb1Fb4Cam7CiGXEqMhwcZouHNh
jKhFGX7OwXRxkeX8eunpgP1L9fJgg5y2Bn1QSIVjlM9aodYB04dnhXilDO6Y
LNtTAuDEcZc33Hzfe7bwCKUHBwZF8lZgOMkn9hoQV4GZYDLFVCkRAevBcHLo
q1WuHg3VTJUGZwXtA+pxtHYWE/wPd6ck9BIsap7rdTQjinf8uztS3Xn8/B1b
w+JZF0BKA5W84/OP8q2ciL142cJ4C4SyGKX9BebleBs6R5tJqBWJ+7htvyW+
JlrjCPNfqpLJHahSWakq78QE0XOqVO++P8yiK7kOPa3LhoLoBQoeS/ZDRSPf
oSKTtwMCPFj7I7E7RwEwR/jBeexc0rIGiWo3WZ6QpRRmmmcUZVNaPWuOqrYz
XlfADV6wXOVNJag9K4LxSwUGCU7lPT9l7okM28ezJMHI1CHP+OPBvVZOrASb
W//Z23k0+DVgGoVkP6qt2PxAujfzXjX95dnrh5NcV/9/194sLCRuuobzKRwW
VyCrDrAfFnJ75hgBayPkWE0fj8NdwRQE59cPIElOXEla01VFeFVqLbjC5tTA
5sx4h3JOiJgrTRnhkneT+rFyd0Xz05E17wB/1pAHvX/qREnQczRSpoTaAmvH
FsHLMLq2D0UEjnH57+PyYtOe62XncRThs6Oiy1p5ef617iI1RK1RLCrQemtQ
KQi5Hu5KCuW98kMs0t/JyzMNl51nIKV65u5A7n6nqBfvh9BWyjqJjae/Cy/3
bq6dKOnukyL1hgmLrSiDuymxi0lYgl5tX+jwOLD0nrGMZJw1xO6GvUTxKQFu
XnnSiYwgNLQkf5KX/yCWDjWxkBLm0pTYdv9g3h3gXx6wXcARhvgcato7diaO
FhFkAGAD2nYlrd2WlJQXKHRv4+/K/laiHRu/FV11pONv12BpuFOUM7LgMrCW
/4GAKS1mqOla81PYgIhn7wSYPjegMCD9Q521gSDOELiU4D0tqbC9kIyjHymE
Ll5aR61DNwePMyisV76TtEtRPFYHdQufu5feGEwyD4paG9J2TI4wJbuphFao
yQN0pxfThvgXRg0HZqe1P6lPqoriKj5oyFnwzN2dVp+wMxUZhbsfUqROPm2y
VHb1APL7uW0NBfggzXW2sljkrs1VwrMVrcg1wVOQspgK/B5WR8qA42l1Yz3a
mi8Mj8tR8T8/y/oPvzQ+3L/POEKr4Tf53rzhIyX6JhfWl1YLXtbrqtLmJq7r
AGpWL+xzkB90cBfy3/0lssAH6ZpDdCZxTQCBrgjWGOuademhrmMPPHrUmgUB
Ehz4SWRemvXfRQ19kNKgANagZhFMJkkvdcZu/aLrcaMyIlABEYR0r7PhYt6A
0bWNkBz8bMN1dMs/Gq1ZDivqA3Mqd5wgtMIw4uafN1NXIyYE9sxMJHLR7doq
l3+SAVNGK9JJhj1kv9wsSL5YfQ4hl/ixrG1BnatyCTZOoUs6/T+iV0Nv3CGN
hPmcinDOhhYsOwwx5+Ul3Ah1IkP98EFJWnNbS2tEOaolrsP73cAc0k/CkqUl
wZQ1WZ1zRNjF3Kqop/sxZpCgUnQNTOzevq8srOxfrQ4eewHgPPvonCA1gfon
w1I2Qp2jRuY8ZzUBULE5zoP2ixzlNQ7bxFcrgA5XRcSywoCTegh/QVSdNjlT
A594NTrOk1dlR/c32pxgVudCh/b3ZHp64so/Qp27tpf+eVzyH3dfePCdrEMd
ny7zs4+LZotTxJgv73wYts32CON13Q2rluevo3WKR7fDSk0/9tyHRNw9FLVz
+77MgjIpBxAIu2Ud7s7i/0iG0ITyRSNm3JljreArAmnjSJeipFuerV2m4wdM
qvVj7xSD9AQNwQawGS9/xN5aeU+Y5+JAY6NpNhOKjcJKmErwWOlG/STaLrqw
XXz+3tpjBaE5IG9g7DUPqFjIwouuVUaVZLXGxMJfRLeCXKN4vjERm+YLSY4U
htBJ+XuqFXqMenMTRDpVMfOIrG1Wm1Blp80Gg4e23sUMwsEvCFCZeIqwybjb
i9K2oN6IcAdZzSg5BJFCHij0F4c1cd/5nx7M3LAvWBSZEKK81bvj5GU+csKE
lw5lVgWFjQ0nzwzu8VtLZ5zZGEEWHuV3o01Z8MPcTkMu/9fEz5CDKBmY1HOc
3gRcprmwJG5uowMj5XHuGG6tTHVe85hB8caOUj37eeIdNvb43tyR+Hv3nsxD
4S3kxX++lcAzO+QrpJApSG8q6dUKzbHXhfqN/4afWZ8B9azLLxGMlBhB7Mlm
XLDM/gVxaPiZ0rARD9IRdOau51u0MLQP9+qUTm2izC6CI21E/O4f6i+5ZfeJ
KQb7SBh3wCHKgQxvV4DpS7OlGdsbnUarzI2W2ucXFn9vV9JVOqdQJbOyOa3m
Acocuxzz6DXZN1O+FGfIm/qCIq0KKePiYv3J7RWZ7tQrt1YgyQr9wxo0adb9
8whTXESvA1+uy4YyvsecmZQFdhZGFE4ylVhM7Rc/uiPLthwrBstAgl02Tmlf
HjITrVzIlxiH97X+iH0o0nu1NMvo0i1fjYI3ck1YJZNMk+J/Hp2T3rJJYIZ+
K33Iyw3o9s/KS9tLUUfUInl2AxfDyhiI/LU4ynlE0kFff9sLz13+HCPykg2k
EdhNEoc/wHKM2qX1iOMt20rQuAjCQji/5oowcp9AOywtg6AZL7z1jGQGuKc2
q6fKct0p5V/Y4i/YbeMwZa1M3FM3wX8vdMffJc1H3FMwBbfOC1rNlHuZHjSV
gF77Kb+/bFV+jQ4aEG247IRby1ceBAnxmzX9l90XnLOy5YuWffvZ1Nwd2vut
m7dMAvrMoV/cO2X96dVPhsbaE1yHaSTiYH6w/TC9NecXdNe5Xn3f7oaLue5a
biqcGZhbfDDWWIaQ9dbiul//3MHLlOyfWXOkG1WFlvVsF47BeAxmss2pPxHq
drlEGYrwa1HqZpDWI1P+IzW5s9qPPQjts2NlJy5H2v6MpB3hcsdy0mK/Wi0q
vMiQkCDA9pa3C/K6DdVBBYn4/2FQXe7uhbzd8P62HSxhhCivpJH16X1A6Pk+
mcMHuCfzqfZyj617bijjKDBr/n22pzR1scjfr5is3ee/5YPL43ZsmlILpur5
1hptDRf1r4uDP3DvuHF8dKpiM/bVlXsHe2sustnoaA1NSJS+Mk/1vQrUTfBT
kCiA6PiCFl5IQwOM/IPHgeK55vbu4/Qy7UkmquzeCppHipcBwpsNph1Ylkna
oZuv31+kWhT9+AvrX8OLv+iDNm8VjFvkhZT/kG4TKZ4wKyErm6mrbKKCLDlG
SbKmO2piPCHd9E+rnbfwELgZi0nQkFxl3LdxXWsh7yGz1ohwJeWdYr4rQUGu
jvG0q6PYQL7cBUKnAPAmcalMEZoxMdlmynJpJ0tRZiYrW+Pm1uy2/oi0m5cf
80I/TBLj23kKFLQ2RtxDawpEJQcXFjrl1S6j6J3RGvxQHuep9XDF94kq/J8K
c1suMox0Q63HP9pFu4cmxF8UF/gRBnMkkEnb8Lodbw1RTOMASi8klQoPEuFO
IpuvP9ylm+jlQrz8Q9ZzIvPHo09LoeLhawiKIDQXr2x+FSH+4c62sWEcAzs1
RabKRJNDmWtVaINSRwYKd2We6UG1YxfxUHzxEfoD1iSwWZ9cCRKFiim0+dE0
+mDu0kZ4uvZncW4Hqi8ymtUCpcjcDZgBuCCBT8qGWl5uaICDHZ8hJgW4B9Wk
RhlOG9Hh7IyGbfGu8RdBeESz9IUpxtkgivLSLUrCbr/sv60G8p5JkEa2ET1R
EgWFjXZkfFBFUWzG6AqOm9Z0206Ze6C6WBQRmA4ozY+vJXYJ6yuJt8rHsav2
8QH0ozyR4MUBbi86CZ2/uvEkx2ll7VP7TW6H0Q4eiHuOA04r3CEXsOd+0unj
Hu6pgLcwVz4CwrGpumCfcqIUWgGDNSwf074j+OgIAOklCuIxZSGxjuxIgEHV
o0qK5WVx0ChKj5XAH+hI3toRMAiWvzBCAYjaFaI32QKo0rmUWlENvIpQIzbJ
QEeSt7h0v4WXovtDs6lQumE5kDXf4yKyv4ZHDJEPCW1T3sJroo57K/p1jwjw
TNu9JZALS5UTZdYhrhz96ufb4o0PSLt96uXKZsQ4EHGkmp/uOEoPetooyLgR
RFf7zpc0Tdzrb+g4mYoz/yPjkKHw+L7thDy1TLaeQiDfWZ56o5p3xwZN7yDx
2v/5Loo028P3QqTdjhyvAPETvE+KVUK8qwYaN25gAeOaWvg0DDb5rYmMZAed
M3Ft1jKz1w1L2A3st5yCVAAWsn7zyAlRHfWq8mWIVIJlrJPzv+jCNX64vx+V
USQ2pPAkMQj34fKC2NWNeQnivBti/T3IVwUlPAN46yvZlhbsfGvTcdlQwE+o
k6t/voElGNdmGHgiARMP7quMP3NsMYLiwnPeyLyzr3ZEppqSXb+c8QJQmQlW
32tUHlCY1f3h/WNOsUyR980YlTC5xhmVkgq8y/Tah3Y74+aqDalzGGq5rDzk
qYbHr77qHJhHmVFRcTlM0PSEDtIclQKPGUiPi/bw9Gx0T26N20OGI+feteWv
jpSC7JxeQs/QN0WZTuzCekHZeTzjinrp73LUdM6xaLv3xi119RwLJudoxAv2
P8JZbA1sFOO4HRyzRl8yBcWYMKjBIHh8EiLbMcEui8ZUBweM/4WoCJRDI2M1
AeMQ4TyPqvjDNgUUxmRewq1v8o2e04+/tOW6HSLXbl4G5ee9lMiVwQOQTg+9
2YABeOxSn4L+c8wLsFIKxaVHDI3AMdn5sfOskN3wHMgyGx3UZewtgPQv2uVv
kQfrqhXZS4jo8rpyCiuHcaP+47WRXxL5uoMgDLCYKyPUl8rfXe7AWPBNe8XO
sgESm7v/JdLwseYPT/5b77nsebsdXhCQ/2lAK9zTt6meaSgQHH0TNVuWRfda
+Cwrw3LVtjcxNpDSuEfXoZ2sKKIHCXzbWnp3ZI92IdBeiH35cUjukZ3/dp39
GY6VIfwrRJQQqPiWgKZvMKfIRMQlh99TU6LAIbnu22vRHCAqtKV+C8xGuGVC
vfrQ2zkjKu4Cq0XmpXOY1KHyWn5Ka/vY51nm94yqMEUvLzUNAAxnAevRLiFj
BtpeaNHdQ7DcJ4YOApvZc3j9oHR5pilxE72af5qB0uuEPY8Zb3OWbcPssmXz
7K7k8m0QoxTugTNkBU+CYMt1Qz79d2sfmpkkU0E7DGkU8UpyaArKcULTv/nw
hXwDpRmTea2ppVBII4H0Z0ezObyN7Fm3/g+9XnFH0O2dkEeQwa2Uv2+XxXu+
5muA7d01dS6f4MMQoxGJ+O2dEbnXbGhhTLb2LCRB3RmAKk9ACKm+ESvePPVv
RBbNFEqwhvJqm+bWz2/FGfQL6TojIvdt2x1ZwakDHESAkp8f/dAfw2AYZ0WC
PJ+ifNJDLC0nI+kQj3QI02VQo9b+Nz0THOb7MN4IWgUhCSq3IH+GJ91j4gGi
L5ftvfYGWCho5PUmOM3KCnKBReIHeii06AzVAireJAjT9wUmhsmohx42QxhP
Ok8qtjMFjtDRjLjCwa9kpC4aNZRcmsIdT9LW4bPA5OiiTSqKTNxqSlkjUQEe
RtVdRHWjOfiiLstbBdRDbCSRQCN1mN0semy6wY6DB6tknXpnPhqmmn4DERXb
yitaEf+ezDz67kVVSHy+qOVSi3f5FSli0u5xlfR531W2E3CpqrAA5+nPdGz7
erH+1qCRe9AM+kysYGtVLOXonLHXHrAhm3TJVJaIekgg4ADAPiYQIAzmsmAJ
1oN5vHnNflDoYS74G/P7SaL0wOQl1AcEBxGlwT2kRjV+HMZ4vh9etCHRVITb
smXmazuwY7WLbL2JFo+1Xo+xR5WB9YbajFq1ZFaf0fMropO3CFcQ8MqCus0B
Rijz8rh9/k6GNq+td7nq04xgUj4LNe5zaxpoTf2rLGLE+ZRWEil/ZzzYoIaS
mckFHVXliJB+eopC61Ku4cEVxYA3ydA8fXXhvNcTQloRw6XyLtaArlC87aL6
uqO2GnFY+KT9Kul0KAUaHDugCjGU9lpWwzzYYo1+ufmDQB/lnA3Ty3cob3cF
QQM8sKK6EW19jdPxtgk2FwrNUv0QncN6mDv4JSaNLj2fjJQYx2miBOtOfyMv
OuMO6gClg4lw6PXQ0t2Xcn5Eqzd7d66QT0eOCFKmVKTuh1+OLIvsZmkryklf
dgXf9OV2tcoyOHiwkSRkH8XYaGdB5yxFczWwlYJor0Tg3C3iAoqU+syvJmnt
TXRDTLC25m2h5D9ljx+eZG3jSL6H3QarZwvk95p9P4FHRTjuo1Mhuu7fDtY2
/3DPmG1jRTzphq4EYvuBZQNxALaVwBgMa7J0wDD7JFAwblxzw1J1CNNikZHr
JuZe+/rb8VhbBd5OFMR2h5+7i6dV/DztLBdKVx+wB7g97Te9X6cDDJa0RsuV
jIRw9tRrjedbST7iznQ4gxlCWzF5KGoz/9It6buU8hMpcZ6fACcENSzQLGVU
QuTtmr31j/0kePynL/Xly3BTI8dCvbUuHHo8NPx+drFQp/3s6rmMvGq6jDJc
RR6MCJDTjn0QUI03QnUA4tRYXupMk80XzYTi+BEG4RN1P9HZczRe2DVRJ4R1
w3jG1Y4KboqWfyT8M6SZPnvjCmv7Xiso3XeanY7LFFpQIawBTLSyVZDS5Q5N
azKTFAw9UV9MV5uFtDX+IPjFTmyhiwyRfEfP0XRrGFFzTfaVogELj5+1PSkM
RDC0wrtHFy9IXbmCVjB46XMg1mx0RSWykLbWA+uPmR6xyO80mdkF03Hfhj8f
stPuuQngRjDCbfmPrfiROs68UcEalN2H/SfOczRAyS5euTH5S2ltu789BIvf
NmD5Kxzh1SHe/DhpJb80sw0mEeTtoGjMNsmVchjITtrv4LyQ2xvGrGV0XbVa
tK9LGZleM57KbIv8P7pBSYqcN2XNTBPKCI5DrbDE+ZRWYYHEbK35HiUbL6Vi
wHs8X/yVz8EBm1k+QUKVVyCzjZyAAk9GF8UJw/bsIVCS5n5YJKXTXmDiipfh
hCb9eXQNm5N1O1J5VZJQasegp2v7KANeqfCIZOXIOhUCgbuDOw93mVR241FT
M/joePawDW4tZzyasV514CrVXve5BpRflE7I0HZh2yZieksgBHjfKpkNtfw2
qwXnXzsO6qOkOrMtze/CT2TfkwotV36+x/zGPy13lkrZr1JbZ2dfxkTfZpnX
0pDFdTQZ+EG9mkkY8ts/WVsWuox7d2llUpeCkUHoKnrXvnkP33byyXwppVp+
kkUhiVnfNjuLr9KOdw3kESKwr9oJdtnBCtJ3uLaB5XGI+pXdPhK2S/pRgHhb
gd7NXHLeqVQ59yzXUF44t4fpoz18HYSXKKK+49FbTPXYRZOmAfm/Wzr2i2yI
nFjZEspRAN9pmxWUzD5PyP9SI9KdRRYvdz0fpFJfXxyhuYWg6z+CWz+bHxmS
hUVC/m46ObZoPtT2+Jmpcky2abBu4mCSiT6iicD1b7wb453qtXK1PvoHQsZ0
SLqeZhjZmw2Bw4AXh+w7W3xPIrAT+Fvs7TGU24IjR6YvLR91CeJ5wubWb5DU
rSh/J46xuUs5UT/ZHEia2nhipq8lLbwVXVK2al41MvLUdN7yJqjij7PGL02l
fSYb7xy05ojP6WpwIPGfkzIOjCQnC37DfpZvXGQQ27/39jXIN+xRhQjuOxA1
xXPFfiPe22yS26OHm0XoFDhXE1TJGTru30TPr+yZdwoCIxzslNOkpLBx/Svu
nCh8Ln7Dw7Cd8MVPc6IKOKmWLjolLDLclIh0lg8efHSAVa5k8sxxmKGGJsLm
mlEkAQ29MWUYR5bXVaQCJCELHyqEhjPeqBB8nkxo4XqBXNO+KgJkYD4JtMaP
I+bsRHtYnI3kgvHMVplR+1vfS/XR6MbbKMvPjRNksrVF+eM/thBKu1WSCNlc
zZyP4je487FgeQhoEGDJA0yt4tdYYTf5RuT6TO1ufyHp/W0QK7bapufV5W6d
Aj8RlDFk9Eo4N98rajCKZmcRqkcu3m/7Ynoi6du7B6ME0Ig9/jWDkt/eh5Bl
6ezzglUCsyAbAU/rSissDsg0/8yWKFbZsnE7F7x3zcm90yl5k7KWhCENaV6m
K9t8sCw6POQrv/LhmzMU4LFa37a6ZcbfUsyiUZXk9B3ts+18regVcsM4TKce
R7jMrtmymBQ//5wUWmd/na9ev8wzQZwlCellLatQPyVWW+yqPoNNkAnCaqpe
6PTQIiuydJHx/25ScBO+YhNn6BG9jYgrU1OsG7OFEmz+PwJTT6vQGDMZszAK
WyxB0SAtgdaOo92LEmeJM2qw58XZtgffUfgqparE+CgbuixRfrn0VsAjj92+
ud+kNvTJ3FUJbuXgrezX7jSujEBPmLRbE6gYzCemp16lIBatX7YFI/w62jpI
bMb0HlLY17+AW35vpeMlPVGT8nZUJGI4WGwyoMI8WVRTY0CBvLmcXtLFASBN
EVuYEzhpPN5Tkss+coEv9UC97VIgfMPWVTNSd12rWffmix6RU7uiodh36xIz
WlEpSoXI4PwCGjpxGGADYu/mjk8Zs26/ukNDzT9yehmtigc9mSDQjACG50kF
jPmubLjXDfe8AsiDHmFn7y9nVOJkASsyMb1C6ox1ebRj4ZJiKk+uUbc1Bgv7
kKKb4LwnrloN/HBMQxEkUJohFEoVPzF2MTEUvQVna9xqZ7pShqOqCTCMzsgu
6DF+Q41ZLSksp4TbjqYP1UgHJYyETag9I43S+wD9OhfPTlQuZZ9v/Y1hy5yw
4XN1cao43bUNBSrSEAs0Lc4l81N7+Uat7mVMQRG3NHSBLo/KxcKkKPJg9Bbr
lMBKx1ZlJWY8MgMPtqGe6HZTOFXUIjGwNIPM2Nrraqrtz8vOlurKd60Wzohl
RUaGhYi8X/hVrcv+uvyBc+cYU4CFc9HlNab7vYt+wVaHmvshxCslkccrzX2/
VpvdeHBMZc79UQbyBz4kR6/g3EqRqNAMb34FYvRBouYkCMKyTrVMfT71rBqz
GNemjwBIbWjKmoWQG6IMUSOTBVRhmbwZAxe2Hc2pKt5oQh6+9URV8LZ+dSYw
5UQFYlS81Fam4tg1Vl877rIE6jf/JvWpbmHbgeQ56XFi9fUzAMwE0RhrbDJo
vXUv1bANkK7jOiUgHeanqqPKVbIl0jtNe6P8syw/QvazHh8FVOuufKRPJnHV
VaGHV+MdVt+QfgxS4PErEzvUlSb7CEEx8xTbkTo+KvQbcXsNG+/QZlbzx8t5
LlFJt6etK91ikLiFw6SIRcalIl9Hk2VJKYivQBDhJoQljrcc4hyD9xfXQYpw
YCLVj7XTXqQyH1pE0W6xgagJmyTldWADdom8n6aCq/DBdO/2nTfZByB/GpI0
iKaWAaEbq2o0Ch0Nf6eGYRDUNp8386Bt8ZRhDiqd9ZkH9MKHqXVhc1X6uEKd
A2PwdXBrc8pxqJ0+WHZ3IeH/8wJaQ0LvyYgHmHZhojNbM7czRKMXqEKJbFfd
nO7SXNz3WXSS7yVONSRxAipyysqlqr/V1+Bb5O/dNKYUTCc+wqwORkVSOLLH
d1ufvcsSSWQn0I/OeBnR6mdLBoFskjIfLmaeFfLDb7upLPcINY/ohzBsO8BO
dDQscw3Hsg6QjKLjPOCVS1Oi5/RmcEfecXrxvhVn6uwW55Eu8k8g9zQ02SUG
SOvj+rLDImRsEkO/8liKs0ChFSMMMAs6t5g7BiPmuXXstbDRiL+hwPgsPUHz
5cD1xMGbqVsC0cvKlhjuUCgtJoS5MIGNK9CLZn6xyCTpbABVmEN5mn7/+h8+
K8mHpJbKk2IxQrRtwauyQOUrc/MP5th83Ii6PahFv9PeQsx6lj3G6Ientz4T
Ryj1lHxyU+8xWf2VD07IKsbAanNQK8hHNPJvRKpKrP6DwSnIg8Oft6Fo02l6
KD2VR9Squ9LyXWMc8TIncQqV5FWAdFZK1H6hSSw41sS8OHFt5UkYdA7LHBbR
eIhld7jysNhsKJSFQSvwqiPLYaGzGc5XC49Nfb/LetDt/lnirwnNVwAkEcTa
tzQ4q1p1iWx4DjahxtyV5bmNtCOZA0JJzIj3uipq475iSYacDbx+diztZfyq
mt/+8LZfFQgDRxciCjPUPBRV6bS1iuHwoR5X/vaiFNBTpS9YxF4w+QoHrTGG
hpd5AgE9ErztpC2mWV/BLqvtcN+hXbJI3W/qqBZF6pl/2FwVQ30XN3qdUJEE
nnDNscoPPpx0MX9GRkCF09v91t08rAr27JlW/Bgn86PHGtcLrLrTtNslWjDM
bxVg0Nsow1nn8fp4Rk08lB3QEy7tnuB5qKL1ZcRfhvk1tWce6cMTDEJkQUuZ
XBkO6pA1wzbW5LtTTfZMyJzA3pBEv071fKHKIE+b8YTJLX6eXsmNu1oC/w2I
2oeYR3mMgd0OJhsTMfBsmkl8peo8j0+ZGcB6XDr/OD1FUpZniejLnWrS5OsM
OPL1UPQEEVOl4rLhQPQz/kAroIB9EQDVI/W0hq3jtbQ4dot8aAJegy7z/a7F
3A59HN/wq5l1x0ZEKBIkKsNIUPFhHIBLoVr6kr4RNn8C0Rb8tqiymLfDx7lm
BHx8NV6bcpc+MGzL5CWVCM+9nE/lNyUF7X5JSk3uWQVGy27+GsAIwuLRG4/J
PTFQ8MyGzl0o/cvc7yrPBOBuQWKGnMXVJ+tpcN8ip+7YLUTQiABL5fGLKQAz
sTMxu7P+xSrWMPnK68YdoTsCrPDJ4WiSscfqDP2Zq4TJOfUS+86DHDawS0HD
/vEM537KwHnd4ViiVRvvQ8F/LgB1Nt5ygwJChtZW7ozIAf4QP9BtnTm8S1dR
qzVZvtIpaE/md7uqo6TfeIDwDqQFlmT1pA6A7Np0bvigi/kL5x75QEA0OzFI
KEImQpm4ihBVfPcS8n7RT4ekCzpskIkH/G0wDOvl4rieRpXV2fViW2RkL4py
Tlf1aqvjSwMthVWqog408u5zygo8+5AHC4wDNDYRZVs3uQb1CcFXNManAC1H
sdwewrXngWIVOWRs0Mpm7NIrCB44wDsLubOc4TMu/brdqSl/qa2/lhE/9dwm
ttlrT68QZ6jeaUM1Plex03PRjQX9BeoOlacwYeXktirlgQjdE1+6SC3yo3nF
MoFnChFIAR2KISljqvbL9iTrlXh5nR5WC/82pXn+eNbLwiC8wjL+nPbzgTAL
XYB7FkECoq5QZgHXiGmycadI0ishYQNRqbPiYCGMxekLllny/vVVQR7jbBh/
3j59mJMZtm8LCWBKx3Hb14r+1cyxbjc4p0BfLHxp14MzepNLJaTG8MC11Pdq
mbcOOGbqQoXZyVKrHTv3vI2+R9rRg+SlySq0517eC5UZxr+XEYXHrA66RmKb
EEiv51xd0m5gBb0SyQv2ZWWCegTu0S3bZ1D1sBtOtJ6Uk622B0kskL0J9Buj
vjgndqpDG32Zyp4zYwS1ti9cJ9lcKBwMIP9ZZ9jL0OMTQWEI+Vx0sAll/Rih
FmG3/cMwLy6FYHjHPmtVYnHdS6kSOgt80WdGVaJg+cZrm/P0vkpWGoJEBccm
xxvdJWZDwXo9bWmBvLNeUWW5QfGQJfVBLz4RZx1lz+srjydS+wKCyMX6FIAl
y9pfMofvV2FJ0z/OtweRO/ZhqR+7mwKs7tYft9/LcN1zpli8j+ZkoJs5lVQO
yOrUMoT38P1NTSxoU2BvVkgf5VTZfu0K2+7UefGS1MDoZ0mKw8jIu2d4SYnR
4ODlNxyu5iqqZhoxguK88FBOts6QN6yHt7NsIbma5oharVTNkOEw5+1NhxJ9
ZEwyO+OWIMfjkOnUxmb1YtIiYKm3/JOafagComB2IX9372qXp79Z2hBFoiyE
BFJbMFXXznhTsFXLVw/5R+GDzj4eYQVQV3RrXHNzYjDxxKbzNqFKz8C6z2p9
9bm0MA1PdxYjU3td0CsmrEBQgx3G9liJfGH7AuZGFzysZwez8C/m9H/6KGgf
AVLE+t2s0Wg/OJMKl3Y3tN85nhycnKzTTV3JSBEcmL99P5AXXMHUpVccVSts
QWGwmpeHghHY5jmjBBcSs5fg4ZMzbIquYzG/r/INf0+L+UHQjPnFMEjb/qOZ
XFSWuGRS2jLGXqzagNNmimS+/0C4sKnNpFmpfOn3Cqe+mqpfRDi26aMtWs9L
yzF/zkwfxflgobCs/YTXWgAKKB3z2XlTBqxzfz0Mxb1+Ao4fZ2J7e1S9P/Cc
xe+ZtP7+uDHfiBQbiL2hoPR0zGVkGmmtk5sa9WVsGQe70/dhtTrQlo6vAwlp
YldCL+v6LpN37YTwvOJfcOI4y3Z5mtMRUDoDzAnWQiio4+gyhiquQrgUvtHz
FCDpwkx4PjY8o6c4Rsrin48C7ReXrMxuDmIUG4gISQA6P4EiAb77YuxqujYy
v8BiMz332uxst2NHVkV3Z/IjSLfkekUL2MqfyjSDTePcWcoBtV2kkAKF9Wgo
8dpI79ATrPHC1I2VyxCQ6R2r/xzoKzyV0Nn9EHIJKcrmUbAyWy3f5eaj8K3q
L1qJFZ93XLq476Kc2LDkAMsPttVUKLSTwAwSlt8bEl535NFw3DM6p563kl6f
oJ/GGNs5GOR5fax+/mghC2QpkfvLGpFljWvCs1it8bOK85HSFMjtNl71B1FE
8rTtWFgQPTHiZzn5Y2FsxhBppcAOuz2AfbR4As/neuT4Vb0cIhv9jeCxdWef
hQ1jlPlfnm4DhZzLTo/4RL2Lptr6e5egm/AdhSJIqRQwwHnGWM3VTINE4kYU
+wGrbh1+MXFww+yKESVyQqYEt4W2QPBk9Jt646JgFYgAtYVxJKoS3IkZjVow
krZjxODeIuY2nfOjwegHyDU/GhFM8Ggt9zEAxcUAtxU+KTg5ux1MHi0X//jN
flKYV0FfVD3uMd8kATGWrXFQkFQ91FaAbtPLdSk4Mo+5Hi/p0wN72C0+TybW
pBg8/4rBMbK9R2U1rGro3UZ7mBZnG5apRfTXGwKy4Bc3cJPWboxbpfRb5CHr
NziOsjuYCbriVBksWO8l6wY1QqE+q7/4rq1DHrafMtiHtvzer2lyw6FlRS7m
dP2X/hikedU7JDetjRAAfHigDThKopcg82wNUyKNEXa4i+kXcWgagFdOX4Tg
+5vAbnz3KDepKk+bzJcdLDK98p4nynWoKDCLUAnROVd4UfQfXm7QLrCWDf9J
om4Dmj1VusQDRZVQqzzwvIFlF2Rq5CHaKCsbre8yfwlbUnj+PT8KXsRSrbNK
cdTrjriLQpL1YAV9w3N4WwJQOdLgNutAPoCFPXc0PnOFYNzbT3iCmqdZwAV5
V12Q83Gav8N4Mah6KVG0ardbBHZWL5Hg5aJZlOJ02OF6onK6sEVxWGxi/OJY
uUvPcD6P7dAYP24tkzTCsYWTDOfSrLKNVSi19zIkG/t/Fxx0BZ/1HWMTPFgO
fUwrJ3mrkM5nBbLsZsthek6imS83B3G6nE1e3bRz6JucUDeGvWWjAt2mzZ0E
L/Ufer4fL7+imiF/bEjZseKaleBYMpX41XZnI7LQZnWumM9s37yGn7mbNJF5
Ouy/M6L2ogG1F/qgAoZMZT3ChwfD7vuiqAPYtD66Z/gf57ulJ2REfR3qHcSo
0SXDRlf3CJcorntpHxp7/SdeOzMZvSZZ4cmNvR3+ZjLYEY20XK9/D01sDzhc
VICObb2r3mDu9Td1W7C/C61Ysbul2fQxengvZMt6v63x2dzLSXchc7ChKeca
p/qMlzS3HdRzmGWIIcl3BIHeCGTC0HGJSVar2B+trofEMvNgsBLfFuUbR8Kx
2Duh+QWeEtOzVBBFKwQ95+NBP+rAtOn0Uamci6Wfh4e2J7+X3OA18MhvgJcD
XiKNw2K0VaQylfSqNUhwnQ3fhu8khejQTy9v8SwxSqYTi8nOfYKVTnbNZ4lI
NLJZeVA6c5AAH0EvFHkdW0ONhRFU84+XrLGcU8BU5OPW0tdP0tDuMmCmUIc+
2gGzzlLqyqt9TKD/UrFVlHQ3GfUlhSCyDhDTvIwUwKlWP5B+NXeaNbbC6SJl
dmKU4veGOf5E/Qw22Yav68BdaSTioTgtwkO/G+/3EGFt8gDuILlDfWLMVGZU
AuM7uh74rIl3elnUrLmDMB83yQb0/eVTVbqeGnXsCKnbStFwHsH6Zrrj5P5d
HJmwlKzrBora31kYopjk2z7x+SBFm87XPd7pZFaAWEPWhfRXXWt5zeJkxUwu
lrEh5Q9oBQ1J7OAHxYjkb3tVZbTWXBrpnO2UdcjntfP+9mWUDWkOE3+fOzR0
m+hxVMtwI18xDXq/5mhdzYaawnAOLeUfcYkK8vfQ305rnmWFC8ZiYVyPQAsY
3aNgNFoSML0WtXQTIWjNEovmuI8wAEbeVLUwcn3NYBlHj9/Hywt/fa5fyFrW
xX8shoqrJtf3nGIWxYAz+SY2ycK9XRXACBbsLniheoJRwnld3PX8pZERVdu3
dNOpZbBGX7ruvucN6mgjo1bbrHmruXD8sKvs5i+TOBdMhfakDgiXDStlVKLf
zPQjRHH59hKbV91oUdFsszoPw/Wn+7CHs5apspTbxmUPN4z13CqcOUV9FHCG
XShjH/e4SMLn+gEO2pQbGL+lMdozT7ASU+BlUVOEA+AxS2Xrz1X4FvCoJ0e7
PnKkpaI8G9PeoUAn28MOQxCBieUxBhUidJgvG1CavNGB6iZNN413UeXwDbUX
ba+ZEI6QMvMI9flpx7iG3YGDE4v7NPVlpka576TRgluHCjqKtSYeoQRsjELy
CqzhsakjSRWTiFDSxNZ1HHXysDsGQFajRiMJ5ROBbP2sLZyC+PjuAwXMoZVF
fQ3YKPdZQXLiZ4LAKsbFtpbVS5a2q9xWBU1xmF+VE81obdeyMNkcd5FxUQo5
teCDzu1ljLamzggr9UoRQ9STqz3KteU2YP6JiaUwUGddxRxxRdGjnDblhY/Q
7WXy6Q2a66LAySCSjV6k3uqfd70grIkWNjJdzZoqahb8/AGFvYJLf8bbLJyI
qsAKFNM6irxxprsy9CAU/YfoLodTCy+zpxY9FbHgsL+SyIqu6CYAFDAKVXa8
0mDPWBgH6c5Tb/lkPjP4bvoT+x2Ae8sHlaJUPDYBUPN2KQBFJopOelDXtjG6
p8N5Zq3toAt3jttrvCwbxhHNB5jLdHvKv6mZDCSrpqPKpIpWoGR7AO1TQgWz
+kxFF9GJ7mVc96vYbF8EWOFWfBVzXlAR+9S5dXB/AegEJ5ZMP60aVHg4YziB
oJWG0MzST7uhuKREowFdmFYLd/RDxkOa0uy+Tlg9lnj7A6J7fSYJZw0jFNkN
PjCUeBTkZKd8spdQXjJ3nEzOPZcdVrgmmtAxjhV5VGzyBLdpUHO2ySLMUCQR
f5hYlT2+tZ/mnp9/hQ152c1AT2I/22Cg/XV5F6rCGUKb1b0FwB1FW7xYeAL9
g0+kJ7Fowul6TP0toMH9wdD9XHWcvfwslZEvNSPMx1LVnNKNhNlEJ4z7ne/n
VmIzJQRkMRq3atJzabNGSgynpkYS9Tws+jEckEFXmjXfG441OTCT6oeKLO1f
vGsJ6ILr+l+BNLvzYacYbQFzu366u2ThE+m417OgkwxXXdtgCN9ezOQWn+Gy
fLlKJq1FAxpDOR9QLeMzi2+5wKTMaFSuhU4CZzheAUT0PGsZkQx3DvqO4ELd
iyT+Qe4b23TA1iBVOpo45eUZqLEATzYsHbbY49IoJum5Xd+5iXybSxy/8f3w
zQNwuac7hUl0JoMHlFYbsA4TzO6TeyjE9lxJXTJBUcTIc7RqCAUstm4KpNU9
1BLR2xRAVwRsYaPVAERjN3HFFgn4BZ2WYmQc3qwsyjn7ifUTt4Utb1ozTQuA
P0xOo89R2rrGW7k19vAEKRD+XEY0h/PgcsfmBJwZ8CkJAZtS6BQC556XvMW1
0iBaho9gOdY2Bw7gD+/d/HpXvi76V+pM8FvGMFBl6KfIG2qvJAUNea4Uo56D
fgfQOKOUFL7vtBBllAoCtJQT94azyeRAp1JoQHNeSdjneqoGt1TRqw4Rnw02
tAy7Qj7Et1KQpKZijr3JEyelis5H502rGeicXzMytrvfq0fBvsLhyWxlNB5i
PsD3voSu0r2/2rkth7DM4+kP4vs1xvFugpxaLzmyrA+5R2QqODb27JB7d6PZ
2YOeQbz1YTnEjRg1Xbsd+rMpFzQze4oDbJbdF6ddAGLafyI6mk5eWg8E4R2D
cjH+xVaDYfLGkv3sMD9rBKmrtFA+G9VFq1I0vO5fYobB6Mjsp7JSjlizCLlj
mp/5ZW4fwrk0w0wLD1n4FCrNxQX28tJB3jcz8tsMoa9Gf0Gn0pU/7NHcvNbj
ZgGuaMEf9YXbf+6B0gRZ6tJin5HiSToLwnaTT2jTxJSTrQXgQ0DiizLibagl
TbC/IJl2UznejGeLKefhRUcPPhQaiaUZX5QxmvSfa/1BdEazY1ANSdm3erma
w6CeXqC+/ebfQ01Rqy2s2V/ustIHBcwjUkvEQbxMT8WDUnuyokFjxawy1dwK
uzNld31yV5M7yn/NMoXp5l7u/kJw67a6m5sEwjiei176Rtslr3uHhM+mFZaF
vyFnfTIcwW8fVkmBMW9gPuDNSyiR0s2HXQt4k9pTa46f3Pvfmfkseow/JdEO
Wapdh6pH6N6XiyEnjntfOJq6DCxsKH1Gj5Gy2+DsRib4MazwincaRLAqVVj3
jz0mvCnGFeGeVKReK3Uwa+tjYSAYRTqaZZ/QRrvL/PiV9r4JtOJtXkYyL4lh
cpWIGt6ZBR0WVdrCuldIkzi48qYU3sG1uDfbhyXXrNsEM0K9/QjcypV3VZ8o
TUk/fsooFIUfc2TdlR5ZFzpgmR9qFn4/TOTtS9zqD07QIja7eb7W0JwudxSH
gofJWB4W85au9qPLCOoCY6wYQks4UbBsTnGp+ZYJHvTdyOApkZ1RpfLaeX9W
nFCw3RFQy2062DMz3keTPukl4eVigWvCPtKT2fr3omcufHwiQPSH7HIPxwPw
4u0ksnjnY95RlHnosUHFt0y1DiYNjaA6+eafh4w0P0Qg3AX3hFjrJ/c9JAVl
yyWrdSIo5pNMXzXM6TKII4eFFIZEpMAOPIQ7OXWW1n7dPEOq2xzineA1idSz
ViKgI8/wO09Cb7L3Igld7wlCqS+yGGIylxEpF9ouMrQzAlT963Kt1zDhYuTg
+0g+Hc1+TYUWFJKg5WqIkJZ9AxDhr0FlgOAEKqOR5BH4cXkWGH9w69UBDZFS
aEPvlsnOEO0ifYAHssKKPO3zcKqWekKnKZCfV7vfMTQNLxsFt2OSniNExHFn
jJZHed1pM9dxACSeDuWmRSOyQk/zuSuoe+lcUFAlG7YTVhYK4zMSpIoLI4UT
jGCwixmtlL/lHIUOrNoZnIe/DeQZ/PnIyndEvaX5VCXKsSYtQgU0SkQqhdeQ
PYu3yS7LXlT8Ii5f4U0zM8KkuufZEe7ZPP3MHTuGYiJSeTO8jMGje3yDENCX
YODBwgEmp1iUK9HEK9pnCKtLMczCoo3TUvQx/Gm+4DXDU1N5DA64HoIGqI3A
OpD5Yf1gkGn6YRzPKjrP2+IyCctIv4PMWV7OYUhjoOt8G9MeYk8KjHbIGy24
Fz1e94On5qGzGrZmaeE9oKfMq2KTo8O2oQd49QqUNXpcCHhmtqUuR8i91yrF
Bzm/Ppm5xX3rzx5s1bWFqfDp2c1LaziduGuBdbKaiyASOUZUW6wrnijQbOnt
8K9XTWDL7rp+BhmkRXAhovou1Pb6PHuRgxx/pvZoDUyGefRKRU1oCmwDQo4q
XX4qMCDDXevQ9xZkTnsTvBp33SUaG07deziV0cCP8yB/JCobbF3NchWmxZG6
sydjJ85W7sNA5e/iBDwJQOzXT1yYj8ePJiplforX7cfh7WUBDN1f3KLV39Nr
KDTTJgTqX4EtW83DsXxUPp2UIdXIPwn1tnnza5fTS6CWMlzcLwMIqIGegoEf
yPQSVa1dbQVKFNYuG2PaDckux646f2BXXGWmzuZZUlhbdrKS3jLWXa8Qa8Pu
ILmm+58tag0F0quu2MnN/vNlgPVY9f3e1SV4kZEXPIcmxheWjOYPHSClw97d
NiRJyjD6zeRImgVq74HHPYhjvR2bFQHMPHwrfKgBrTDRdfjwx4XmC2LIEJmL
4tzK1VZ6SVAtaFFvS8JOMxaKAkNKrmVDXocWBxnAMAEMmaKjgN0y4UYh9sxt
GLsSvrR8NkPoRaJSmufeiiSQa/ykusAiAGBj1Bo7tdaY5qlY4vHBdefKsDbl
WxLCjONrbr74WxP+QNS5mcTtH380Wr/fsXfkCnn9KVVRsfGw+51FvtF2SiRv
P1sBWqTjGY8xC64AoSdlk26ZYWLqKvIBMyxSC98I0ysC4XeSlR7nkAV7G6Qf
6w/zcO2j9Tpvty5D5OsE16nvkx1hjAsMXqKQCjDzFLuhqoWNZWCWtkhqFUf/
uoKAi3v4dNYM7MadmfTEoQvRzhpS+AhdrWG+AB18Y8iFp27ql9p6lG1UnQZM
by0nmHgZ5Qdr1iAn4QjXbsHURCCge09Ro3p5qbLpytwKLm7YgHvulrdrAExr
PZtqJI92XhB3LUJmUZxSj2ecDzY2u0BM3ZI/+dlOIdpWfCRogC1w2q5OX4NB
DjO44P2KJDOUgWb+3zCROUYYqP1ByXykh1pDWRy67X2nYyqlEbyO4XvwwrJT
t6o2dKFWTl3df0mjtRfpCX0Cb22GDZIL1FGHqZeD1rt4NlmtgpjOHGmsC38F
66QrgbrxAu38BEhqIxZ7SXwVk5XUMXqfhBY0ny5eUftlz5QTqwivtfqeKrWd
BSDLfkPA67gE+C04zPGbyF/12zpNxQsN16jRKVQKeBgOkY0UY9+FKP8f9nlg
MCHsgiv2bm2TGi5Ng6BKBdh+SckpJPdEX3C8T01YQGPcjVpIYC02BiVzONLq
wNRn7lDe+tOelBQqbct+0LhX4LKEGN0n+nOqe8qFkf4e7w8y2giIL10Ajpgl
LP5OFtazlNLQLkSLe6phbfx1jlaq+J3bQCEotsCULDgcSgOFGjTrB11YO/cd
yE99/m5RfvZ3GmGLpUMSiWJWi1WZ/bmg6QZrABa3bE9cwFiVHLFz32nmZAx5
2NTfWnpqO2gOd8LASnOAWneLaYywAQMNpN4T+h6X1yM4m6/CJUtqW2wUb4re
WMyFM+mphNVDVJwMbM8sp+xRCyTdEkJy5Y7Ja6q2xFzikZF9FHna9HyGPril
odftvPfie2aL+ErMmGUO1+1s4vBYNfKV/06uNgCTxeXbn1+Nqp/cf2dWpT4H
nYayNzK84z1TLr56PpRzPHfIKqM0I35POz33mJgFsywmFPfnC7Iq6ghoyke4
/YKVC53ZM+bl/wsIUvm0B105phvXXbjzEZWr2S/O79q4BBanKgzBAiaUeR8g
YtKUTnEzV1LxcwJ1Shn1C866mODN/swILybJPTxgvvzRtNVdNBwq2Y4HIFlj
jzM4affPsnuGo7EbgVqDqZ3MrVMC9fv/ScTVi3+kvQzW8bS++ndYx0F/DlvK
5+/ie0Rx4JMUZV3QFKvtywepRgW0AvaZ6b1+0mEdLiTIF2Df+dIxB4sxNILk
X/vWlcjiFCPp8fDyokaCwxELDRNTOxXAg1raAy3Qmwuc2USC1sOaMT4hg2pk
RuILy/Js/sTojTfdTk3Q9W8o6fFUvu2Rs+H0jRTSBcdRCZUnT4xefD9Iv84v
NV+hA9rA3m2uDeU7lKabaikvxN9VjwQUZ/GfWY6yAB/d9pl/Hu8M5j47q7gm
l0JUBpppwFUT3ZD0hz0JDm06jbBlqFX+6uElf4NSxqxBjHHccfxC4qwxeGZe
dDIfWAwmSsGsllXweov4j1SpxDjYjZS9G/WkjCveX4mTz6KzopbsHQcgqJn6
iUbst5xUYfM7ZqykXabfzLhKUR8cq5pLZPFJln9P5RUGxVRT0GTg71hNQnNL
nYK2DuL37G67I4duwWFGc8FqMb63x0rUow8QFRD3lHu1gBXqwgyzXAEKtCFI
2l2lfdC6yBLzm2XpSmwNv1ysf0Y6LhPsDwqap1ucAw5108/GjWyl69YVpyPq
MqyiV+qg8CjHKLfU8jdJc16KTR2ridPGBNQHU7w6oGA6ZzoL3DxypgcmT4pW
tsksvTfnN44BHzXOaTTWnva45FIJuUesiSG6ssR9VjTr5/TVcbaL71ZNLobg
eikSxKk3JMTBcUFL0mtPFQ+bp8qU2bPOZk9Y+8mx1aQfBVBO3UIaPqC1ov5e
jG62luVGW+8oF5g6io0Yz0BZxEMWy0K3c/4eYDLopg6daUknp4q3SmMWCC0K
8lfA/GhZnxIyYCsn0tt1FINv6MLFsSZ1Vddy+rYDv8a7q1uHm9AURls1uI23
9Nocth4v+HUUvqKmfpgMmeQ7rlP4Undy1pflEzV1xpA0ZwwA4RNfRifMqMHt
mDOL/x65v3xAWPo/CDolNlUNqC9B49NDzn6sBzD8KgNkFLqUkT8Se4mdRGnN
EosgJwgsgkprRHuLaFBqwBpJdBdXJdjuAudehf+2NxfkVjvb3Z6nqW7ENrJ5
RBVpUMStZ9hQ4cS1kJ7ddhKUuJxXD2iAGE8AeDiAscuz7Ysn0tg8oVLHp6BR
AY77yoHBaQX6pUvwIct9QI/onEbX2tZ1KauYsKOC2SBk+ZdBkR4SpVjm0oNR
HwOUEvSLBFRK7a5/vQKLggfYbl0BCSaTURrdoYQ83YUs6vaTsfqB2VfGALBv
ErdzlE5m8El+A8MPqMdShCgs0ghOJYX2epN6086H3SgoGEGFjX2ZJiMxsvOJ
fYLl4vfvlHaCCZQ3gWuOO1UJRuob0JS9G+p1MnBSgzBU1yYkKRkbae6IZex/
L6+Zi16qIhZhwe2T/2M1DURW/+yVrJQSYokDl1ddx/EaRpUi/VpIQforyMNJ
JpRYPDFD5boVnZBLDCjM8Rw+qVym9YR1ZsB5QWhgP5A4s2Bq+khbJyVc1DNi
QMN7mYaW9Zh7ls7wiwl9Yq/UwJhUMke79pQdTNE5QdLZPpYdMb3yAVKceWTo
Q1W9PitHHXVibWRgw/UyVfM/Gi9DUZx/vIrAq64j7kEpwkV7x30DehuYXIBL
zhOv4D1/rsaRSRMgRioihhCkv22Vk0YYdLnW99kdmeEX/7Urt1rnzeZ3Mot9
GEtI6/ragPkpk8Ww1kxilGyeK1lqcJji4W6sX13rsf+eweQ4yneHTFHEeXyK
vd3YuI2U08NhfKbAPsj5eF1oc094mSg+ANcu6/SVpCkzK5eZgitIOHKl5BLR
2BRFb+1TFTX79lg8XxsuLBHuyHCl2e44DBbJQ8TIRrfy3kxvMDxEnwsUVe7F
eOPqJWJABz0DgxzRQIeelNxj6/vhZy1BhGlNmjlVZ7hNDXqEnSo0GcfWvhFf
ANBs2TiHpddIrZX0wt4VN4E7Zn4qBk1oo+Bwjja8ZgtxM2TjDA1vxPCzSExC
MKFrX4YTYVVd7YQwtAYsFKLnRQ42WP+9K6xA24FhOcbP4WCT+mewJw8fQc9b
zNFXX5xza8ff8jmV2HjQrXJF0xeo4zQFOMW7RD5+rs4ClpV6gtlqUP6OZ9My
M6gTQYlYuKXN1hXsmtd4HLKl9Ce9444M/d0fHfRQLR6hCo59uCHfU6k8dCAH
82TqLGFU+yoaU36g42XtV7WtkVNKXOfZ/BeuiZQoAXQzGrmw5yCinTymTOn3
k5SXJkHoQD1cPyrfnMzRGmzG6VwkVQG6o/FRShdEncqtB259O5hDub6vRB/8
tFg/BA6OlcV8khWD7+5ZSGQeU8hmwoaVzDQxj1Q8XkHvmfYBBSKjHgrpW4YA
hFM6fMvuPe+K72/nnoVRZ+AMLmfDhpctxPHGgkbxGXtliYfGIIERHH7Q+W3j
KHiFoEsLcjEZeFCy200N21vaKApwbySVuDdOUCyK8C2LuMRvGyuMU5UnAhgi
LN793SXHhDAfmyJ01tbYhBhfimyYWpUy6MmU3jwlOk4KPGG2Gt7EjRhgDwAH
yVdjKWTRU9Lo43ByhZPV14DlDR7NFVuV97mUCkt6J5KNvKCzKp9hDNLhwP4n
4UBf/k0Bn2tPWH9JMdk3CYs3J4wb2EmyWPDaXe38WqUKhnQWE2t9mf3JxctL
/1+tehOZGeEAHrWstViaFW052W53JOJOBG3T9AmbahHYtfz0iZBwiFkjPXK9
RKzKQ+fKqgkE4zXebOM57ZVUt7+X7FI6sw4TXQpEtoXu6la6jH3okFUtxxlL
DEq/hQC8nIi1KHriLIjdJsapAgxryPNYMP35WzetMARcOES+oByaH9x5b6Cw
2fp1pRUJNoTKHBRoeJ7VRG0/AAY2jNZcrATcLWuK9XKoIUuCHbklj9z5oScC
lZUflAH7Yqhu1nlzvbmhcCoFLqH4iCTuY2KUbJZjudpg9Mp5+l6sMFIogMVV
LiBC9IONaI/GduAW5S8pw2AMczVWfZVGfqA+eLdAFfgOH8QkQjnLScm8QJHX
lpqGgtsUrSDRiDDjfQWXtNaJdhkPrivZgL2ivXyFhoZzHRuXQc7o4tBXm7Yh
KoSf59vdYxdf+e2xxV0LgGeFVT9jUCmnnCnaO3yevmj11sUKpFCehdsJV8X8
0byvRDYp6lB5scYh6t76WEMHe6juQ82g/2L+uDaX76znCjKALR2r6T3Ir47N
3PCAvW4P6nZMMXR1BPVtsLYQiPr5v7HKXNGWS7loUfCUkTT04o5gMqwuBYDn
0wM4m/KXaSAkD1IkBt2IZQEZ/O3yyNzeS7YZAAyEkfbaLhxj31MOPoFu9eYq
XlEsrDRusA+l5v7Z9HRH8rZZ2EitMrbVlUjATdWdKDbYPjMAMlqZB0qnoJ22
OyVrRjIYbNCwfy1j2Qw+fA9H6iAHIF9C8+lunUyO/rgMBXPRJcV/0iqcCkph
zvOJ+evmmPAmO9gedhvsJIfdTYhd4l42kG7CykmaB1fg+NblG9nVR/4S4f5x
cOlKA0lcV4/FJSIclVptr8ddEaMe62YlgURmzzvmP3f292wcFhy2meX5RCB+
uRG3XqjaSIDRLqPDBEu+x6lI3GCTwgBNw4sNbOqGz67Xi9MuhBFJgMrU79vr
kgsgBWSwMJhzg667eqnVuvE0gwcES2HHb/r1j/qZwFzonAwxDZbIE0WcrxbS
WtGBCe5LWg6DePxFC3eNftO/vCuqj7oP9Xyt8BykmXl9jeMXgOcxbPyoampr
IfgsCYtvhR7dp66tcKSc8ZsA7UZxwjP1ol+GJEJhC6SPUja79rc79C7l2Qc7
D0Ely+mAfMdEjMeFNkZCMGpyvi+JaknFuc07XQj9lqcBOuiIP5VrJ42MoZkH
UC72WxYyLPe2Ikd9nRGW26yXVeKHApOjmxZ/ndeGb3nBV71UzvMbm44d175t
Axrvwpo0hzlkQ/2SGCxyXC4kMTRQBIwnI4ovNbD4Sq9hUfu8h7sOAqZHFQvu
7Ji+ijB2lWnrtvSTuKBLHrC9GZUEo1QqY4nd0vCipeIfQrcSpoIlrHkBwIJe
KY9gfJYPLcRjQq6E5TKL7K7fmsq1Ix2oLdn1AMaceLpHIml++cBH6GVafbpa
sUF0lK7LVyNvCBjGwYHenUPN+6jZiK70RysN2plnYC10n6eSpjZe2xJaskM7
y98wByC1QfMEOrcNaXwu2L2sqEh4xAPoH02Dg1bb64HArFLZNMSadocyEZHT
k7mnAlWnYAXurwph11YRwIPL+iaCM83Hd734uTF/j+8yJ3OMSEiSUvSjQqQM
qGexeEnMe/xPDp3pBVs3MQrKmS78lQ1jOom014R3sv5sLqbxCyLPi+RIaX5z
w9Dw46AsBhmXxklaK06ZZxXS8VYMYtHsmCjIB2VXlHEwiUIclS5zb2UCKmOr
jCilukqe/Ht1ooIa9DgJnGRQKkRF2MRp0514yikDQmnw+ufEfgJuZCQW8uIK
2HSQu6AMr5cgEf321Qt29Z2h976w9f8DBbTc/C3calLkLuPQeuS9JE4kALnO
R3m9qnzVAPgN9hYrY5VR+7CPmk3K/DoSOWxXz+Qt0Bsp3QPUozIaNBg4cflF
wx8QR50PeOja/LjDEpbAjQ08IXTQNNgU9yGJpvIvKeAfFUxwytHja47zSGnH
KZ4ocbpIheVSQYmA/K7qDnKUoH2FGR9jdJLwQVb9zfJ5bM6l8Vgg5G0hlRPg
gMuDNqZHGWI9ZiUzLGAnHZi2IWKSyKzTRS5Fo6HvQEg5XED87vpBF7orWN4t
BJ2CozR3bklRr3cJaJsIge+CMiwgQ+fnEW3I9OaOsDZVSd8Ulc6OJsmuxmIl
YCf6lORZg4GAH8WHcj88vANeswr/ipaL+k9EVKrEr7UW8XljiAs7JpW7RE56
DQwK8dWC+b5wa3mt35akEHQFkY1K4PjgYVqGUJpx1kOzs6mjokl3XxsNVgpv
YdkqQztSYMwhpeGijwMYoJwCLRtpE0ww+pxpiantRHCItYXv555WG1nyehy6
TfycO3iWioNPtLePjRDn7xR/7mVBvWWP8+sY2QX4OBB3JdPOnFb2RVp+/Ad/
Kwdkr5yxpzkDcI644AbhNWW2umvE66ND3OMBh9BCz1D/SN5k2xnGQCJUzEN3
5CwjcvZmffX3v77zLd0IpRrgKiNN44alQD6TTlei3bBrSSeWMX5t0wXAeHYH
7WdqI52sEVjA3PSmLPBFh7FnY2HCGEqCSPhwUab9H0isiR2cIhm+g9czDSgA
xk6X0SUo+etoAjkd1R76OXsM4III7RolVObswbqsyY6CjLWTm5ga5PkJMY9i
c7R6bO0TyVmhypmUPEVelhw9LG3G8dK6yIwmgjTjM5VcWXPoJcgKeEq5Unig
vf1lU+0+sFPpXOoVbOFHLtkWunNLoIAEvo6YcHdoDO9b3Kg7SnB6eTP0kF5w
HmLYHAQWqAN/bQzsIQ3bo4ybCxrauXYu15IsXiInQIJDx1+VY9ImDCGT4pGK
sLkQ9d2K27QIUpe6S4AgIz4r3JVTmY7jL6jEcyRxy9XjyqmaZrfmEpDu6TW1
UAKXMHtQIqVx5YKEy2vL0CJ186GrsO+r/aVenBX8vDmYpWFlURsxNhErDFy4
1ihLoWVOTZtQgpwVc5iBJ1MtcG88NozPl03ZvUfiBmoCmpPmTWzVvczj4R+J
Ap2q7jutop6xl/Xaqf1zTScV3PGoM0sFEk1nH0h17RnG73imTs2NKpO8zjbr
u5MgFsYLSI5liZe5eJAz2HFsr2G945bYmprG8KIODWCjitYFHvQW5cHwJUgo
8p5c6kDcRXeAvU6t1Zj4nPFQyUsCkcZbm+2Q7CyTbs7+6V9up7+F8Wl/7bRL
QqC+vEf8I+35zbBH1DY3JapwEpBwY0cWP2iNVZDGLDtp4ZIwOLbSZ1qzQg7z
jy9va9crpbcbQBicYZeiShYbqKOeFXJvwbGLNmX83w6/RLC9tYSzvQDuEVyw
naaJ9gVyNlcT9He/fipXB+nlm0HG3DOykB2csNHjeR9QTI3esNm0Odfr2DVu
9fRwoD3DMlox73QVajXOd7UbbiSVm3l6gup3rZNmyqW6lusYRpXy3CGJpvIg
PrR/t22VuLUkM2TFtb8oye6A5gBIuyhsmdJMGH+W4uhTU1gJywdsiZ5tIDMU
rvdgAkzYoVzp9LL7tiYwXHevwQLxtoVlwFZN1agAnNWDYFq6H63Ti76Xow57
sL9t4Nq7w4qYvCvs9JA7sqqwJQEUTyJRCwlQuW+7ZzNBnR2BiNTuhd01E9iD
/J4U0ctF4KAJYUnaGWN42t2I0AAgZQ2nn/q4KOr1yQ5Cb4IxPMbtBBKzEjhY
94Y/KMLG0DoR6QGKK61/URECTZG4OX+SJtHW7U74hv7/bHb7OGx7p24zQfCO
fvfVBnyfG3F43NdZHlBGiMV6hm5zhQ0lTmooXTfEG14hpImzvTiP9AnN1CpE
Rt/jUNBCQd0cURdrMZNjU2obS0YRnry83bxOAO+wtZRpa0yZKlmrW2IKRQ3c
NblQboSnhNhbvK0ESl2KRFNfH3oPjF2eRLI0zlbbyvOZSuuxLET3i/EtG/qA
DpHnfA9+xIG4K9ZjsOuJs+XN8G65210/3sC54bZuDIDy4N2CprM95GNPymHs
QsG+XzXVnhQtY4XXCm4GlvM+sh9/rZP88BwKhc3lj+wP/CYfKJNGpWxpar6N
x9nAIhj9WZZ6t1tl/cQqEEyBVs/GH6BA+7b8ZwTeN5+RO43k/rPbc4RjkNJh
dfYpRgxLaJqrpfO4czWX4wr/kZVqMOxbCABKsr8j0+YwQO+JcFq8HVkJ3RiU
MwGzdrQdyCkhmMKGwhTkprecS+EMuG6EEUdMQzvUHdE0yqzLf3paYbMHgymt
hSkIqQCulwesxvsd6NKi3qw8WYgBrDk+1RDg7KEL0ylELMVlEaHHOvhrMYts
NRIEfgLkzNArhfX0RTMo5wQK+No1H3iq+8qAaL8xaXmecWSybM+x2PcTsNKy
YyGGNARs0P9kibJebVAXCAiDbGIt+o17ZOFCn7XFbICyzjKIBwxE5livNUFU
k+Cdb5h5kTw7uQ1sMHe86LatWIdxiZOrqx9z8cH81TrQEdCPusZDxzaGrzxY
fJaHrsZKB334SCs3iZSP3U0EBZwBP1PHZlM/4k3LD9yinSrxKPqHaaJRNQnD
LNoHNVN28ogGNprkBA6oRPrAqe9lS38f8w49P0C746weH0Ua2VpovpADk7Sa
jbcc8jo09EM6Np8lisHFKF/OPOkYUAeyCmg9MIE1c/52FGIp1/QrwfkOLO5M
9SMpcX2erlOZKr00jmH7ebsFXbdKZoRs06qbGzFaztLYN6IKPDYykd6MFXQa
W+gN0duuLiXTxYILTdhY2w2DkDoacd95d8aqcsrazOTiEsvu/nSGlVKtKAuv
lF6nMK9tQ6hab+I6x5DXv3o5QUcBHM5kFpYmII5LuuxvxI094P90EmWGx4nS
9MB6QRsCPBni2NGz4iM6KJOUybWrj7fvUC8AZkgHU4/6QjDHJx2II73A/wRC
7tSAuRIT7KSQKMpi2tA1x1Ivbr4TGgVQzGE2hPgrUOzGEOABYJIVu8mmGPuC
6m0a7pbXrEtj/9yIZ9L+hMM6U+QlT3swNdPe/D8teKyOWgD20zddq5lYeB+M
grpJRF/eRrXFJYjdXEgLgBnhVVkuW7U/OxQi92wMBFDjaW6lcjWxeq8ybCmt
8CrRanCZqqAXFM92rT5YC1CzWry1UXmrh3n9ICaFoCl2cdaemg1X8VC/geP5
6iGKVSHxB2Zsf6Gi6p7Xd2Xc6/+ZZuYyQxnws9vggipTN9rhAicgBJJ3covy
HKUa1uwkHn4wW2u7r7vKHE6FgdPP+XUzsWXC/paKsjDYMIrZkcx2bw2gttEB
VZ12dYH4t6iFN9HgNQde8gjTGlS5GyRHHd/0tyHElLZVZGWwFYnX8CtKmGII
gTi11bQcz046JzDq5gIWpWJ69cplrdrJLvLFIyWMn7NVEY1CW4++PbX0OF+f
kz69sp8gkBi3NcGurJXWLGv+JG63soNcC0cloa6AFfWgZgvL+UZrUpBZ6PvT
IgjlZHrzAPu2N/eNnV0V6EoBzId/wZoMhz4tjSjJWC3mexHTE7Y2MplG1Zo7
0nyIwVDLTnxqMMJPU9UMsSZ45kn+HloGzeF84dg6gfZ2NFslxTBOBncGU2Jv
0qffd2Yz4GhFZQRZ7TgW6xnV4mttc6YEpDW3ynPVDgZeUgl38D6c27NnoMds
LjVGl8kZ8IQTBqDbyLKXK7FuQ1q9GEshUdhq6cGOULMDMrU2GRyVSGsAHeW1
1UZEVn4asXfBCR8DoaMT/HfEdPI7OI9XMMTLGRVXHkRfGJHMNYDxQM0h9n3Q
tg3V5OoOg60iIAEND4QXVhNUkaOpO2bPgpDEmU7NrmAJlcTh79bq/8BJnIVp
uaJJHLihGyoS29a6bhfGon5P5R7x4zHN26D+sEmotCK+4U+X+PTh4MES49Np
tViVe9bO6viHeXLXov25XXSgRRni8bBrWeXnzOBSE98qG6huzJeHJMclUxxX
Y+fD+Qo6JhOOmT9wTh5cLr/te8d2gj4P0i4ueOrBfHhC3yuijOPOT2EwowoP
EhguD4jlc9lwL9CiSq8N60XMot5w6NBXj9v83r7/DWvdQ5dsyqnv/uDYuLYN
9xWBMSPIaM+SZusaugPEwNX2euJcVv/TJTGoCW47td54lJMlmtaEpv6eS0Rm
bGdCo1MMn9aD0wh9tCzsSsrSZGz8aD3YB5Hk2w4DcQAx14PX0QwpZstmwOHd
I2Pb9FBHI7BgWs5jnRhAmhMcZK0+Pp6R9p8EhwWg+4xL0cUdjBunpmr0r6Rd
+c9/1YkEiyopy6zfVQnqIF8YinDMGVIzkjw3fJxfXaXULln2TpqnVpSGHCSm
vg+0mwLYHvCRAjSvgp0gS/JjoxDm8fiKA4T4y9KeFOp+n2Hs81lSwMbNeQ1n
vDsbf0W+gCdldyYCQrMy3pCW+6ss59M9wT50Eg+ebrdgCZHWUpbuuyffCb2r
CLN3RonefQ8eKBSHAboWg9HetAJOuCWBWednFNkcENDduYWT+njasV4HpQp7
VHfODym7Uk8GXpjMc/zNyh5pQp+uspvTH/hftsAcAzC9v7o4Y/NI9KYBm6RY
z3FGFKsjOGrPQ7LzHl5ge22RvknHYYXvWo5hbotfotzjyWarYFN82An6ts75
NTtuYFgwuGGBp8EH+vL4/BJyRRaRhXLvo6RqSEmXq7zCsKqwlrmR8wdSFoPt
QznNmjGuoowWJfaTev4B63wcv1GjWnyu0yfFJ6gQ9Z5IwYUpqC6aTlliIl9E
FLBuoXwRJXlqCTmrY1/mpssXyhc1f7YrpPbuLq2obIDnPuEDRy1ugP+tj7n5
6N6SlqXJLrLhnjZN+NEZGep7NHZn6YmU6Bqo5I+atVnb933Wv6peE17ZW35u
JqFLR+dsocF1rBFjZv1CIzhqds0eWRmGuPNnjcBsCaPd3YADCKXvM4W7E/Z+
qu+fKopOzusuKOUlEV0qpRA/yxykfR92MOFsSVohquy8ICLtOch7dq3oBThR
MTT8dF3BA0eV0pfO9czIolaVdyEdgYc6mgWj9loaOva32ms7eVNC12eZMGIw
mXjeXs/6R2c8SMdTD0bWD8QTnBgcnLrU5S2GWOIZZOkWUs0TpbeJ5T70nRi3
8StidLa/QmrV28Jprc/vVGMnNj+9Ux/xwC6mumgw/Q8n+1tgudeQW05RUimh
wkvzOCc509I7ZIti8z6941HUEXCqf3udVbCF6ZHjt5n5h6D8FCucwJsEkWiz
EKRZ+rRH8pgCGzcs+H+K0Dn1BBNe2CkAMZ1oDyzDHfEGsI1UG5TBx4+9RiFh
lm+r45bC5EK765s89OuSSE96HpFwu6FO8YU5Md+2629HTOrDyi05DMYap7q8
E5dqBraJ7JLcVJ4pya7Q9ZJiD7VXfpFMUNzjzcllfUCNiz/UQRPwzZtruOp0
pBNu7nnidCuaORX1lxUQcUsqoUCjGB4/o5SBnWWFHneKrMruQ9AUK1nADsXW
bPyPOf9hpeKRtjSP9FwlExzi8p5e9beLvrj0sk0ZJ8ZUmUG5KNC916LlxtZo
5j34cqwIR5hVGZXQ5SEHzCZVHe8VghWu6JEddiS4q25g1EiuB4q+oTtlnT+s
/q13ORvb0UyJkZaEeylqOEmiQ1rVDrT46tK/1rTcXdMmis9P609tz3lrJg3B
5+BOiowAHpu5KPWU4McdHAlC14IezS5/1jxtWoM7mq/GAcU8tdfTMwMa3zJf
9pIstjom6hihqL6E25Z8u2A1HEcQ7GeQYmpN2ZE8gjnQtvwRB1flQjeGdtMW
6ZVN6VrszFZXduSNBJZb2aBGR4AoeepOl2UV/uiMdPgu5B31hcu8qWbgumH/
C7CkWFFLTyGodzw4IGRaxaV3ptOlpUhRecvw9z4aFEsxmKrU51mtkcA71lbi
owDqBLLn+sFGQU/DytNUUW/SInkhPAjpHHAhFZ+b6w2viuMy0JjPvqTkYuDB
wo/aj04JFa3n7KUqd+932lPRZ0OBw6KmvOe3bmGqMzLX3OPjlgAYFj+gXN+G
4YwSCgIiI3uyEUXZvwRbY+hfkl3HtSEYZhCiDcCBEwr6D+wdtjR2NJBVZ+2f
WtUlSjfbh2Qch16m/ZPT1/V5WA/YCmejXli8FvcSbwbKmuwH+eZdnfLUiYIX
95pUdfbF/0rBIkdkX3dztXVljYggVUzzgdQVhZSuEr6fTwmjZ4zLJCqI0tZJ
TrNRQAmuKR8XI1aThKnIBCv7chgbqSvaKwqV18CcfTa4nf7oOJ8KaPSGmIZF
LlVexk6fSe+h7EXS8xsUuzzCjtlw2ifNpGD6LDxxoznSgUAgAjiA0koTEjbb
wEJ7LESMDsl2DSf3HFDhc6fGJIUv46gwUzyQjpoVYdddkRla1IG49kww1Z8f
g8BRL5USstYRZv1P5mjQJwuvnCg5o/HEL5eK7t2S+nq78QMtOvTg2bAtdZgR
qgpRvGzF1OrVLiBJBavttjduNfapo11NtFgdx7qv8hUG57yFpeCPc3jKQuPR
WTOzzWkEZj2oPFBwejXNvT2wJbaWiW+F43tKnVVmcwtTBded6USJRBmHhhx3
JSMCCzPese9EG1Q5BkI5NTSZE4xVByNUmWwAYKsikSfXSKaxGL84DxYmDh/f
kp7rAXZrKgM4Wr8VxLdM7+QnB3Y00toUQYqI0QIbYHnOEbgeNtA5GOe9oBiH
iE9ELk4nOzIR2UFs18Af8ZqnSITEaUbC6kNAT0HxXjiu1maPXSCeh0BPjoSt
GddVngyXA2n0MPnHY3h6v92sIHnbaP7olN0tJ0lRMKa9ifBxyGSM5oiI9QvZ
u7cpeR09mNVwXFzZJx94ZXq5ryicQGO+ucnoGk51f+pTppvHG93hgYXnfQ1A
XHk2ZiHYXIozakcSHvOVD/T0tTW0dH0rGIC/Q8GtHpkLNKqnuulb0QAVF3c7
rykCsagj62ZcQDsQ4obUqnS9dBQCiW9gywyL+mw4zSLcusvcKDTPjdxtHaMy
GBypbCQRTsqaDGMluIdbY+37x1hY/L43nXE4kUmGSKj3ATynIAIVAawveZX+
wKpbyb1DPh27s/qzwrGfxydCtlX/eRHgFOEI1p0+PG967s01D8+3pxJxnrsi
H8arfc0CdbXIc+kr3E73AgwdMljW2EN1HK4VLHMbSzBgmlxSzhUCzkqKbfCT
u4HJVD3wjzifVClhKd/kjr3V5TvXMldbmr3kS/fSdw/zMEKGGcMwn9Ubz10s
KyKMgFyjifzebXQ9/jL1YssBBAXzyP+ZpQZtFI/ddquOyVxFrisWoUfa2aIe
Tc8x2wUR1dPcspgkDbNyPhnUyVamgnYhe8WSXYzBKzPrkP2VXeZoEsw0PYG5
ytCpNJEN0D8OLZgH/VHibf+i2XpgUd2NoWkBY0shw+5VaYoWNetE7p9TkAqs
qP9USzw2WIdznqRYOFcPXAoY4ItMXiVyE6cd92fJZIaGokagmBy5PetPO2Ge
ukOSpRHC/TztXpMplW0Mx843hT8n/1Kaa2V3Gu6bZhWun8IiVX1qy9lAWGuT
o8OT+8ve3k4RumTX9u7g58ktVv7m+BQAFxxLoAWLoVQL2Yur/oACBguBBWHx
NX1glSMDN8I3kbKqQiXPJmcHbpp7mFmZbXriNPoEBuGUOuLyyCoTWacKPWSq
PuO8l/r5Hltll+rgT+0Le2RxzwbXRU3UaDrZRTVF8en2y25YYr7AmNODyj4m
Eh/eOk+nscM1XVDGw78K/fO9LA6nMRb5eWwLVRR4rQBYrttSKeK2kduRlU0+
0wisTaD478DnOMJzKjTJoE+CkG9XgO6fv7DO+IU5zWHq3gp8Wul3Pjs1epQh
s0hw8jEzikmToJMfEilWzCCbp5J8QqlrP4pY1+jcUhvyVAfzwLyFImbHpl6e
SCexg918JSmwwTNuEnke4au5dZrBLIT9SM1EXMYki6LZxZggnnK2eCqMt/lT
Mf3NV7jIlS2NSdrGBgPewYOvkxG/8RiDq3m/lfpoVl/FNO+vmRsqlsgMThn7
yLGodm/Nt9W4vCmw9g5WfNQaV1Kala1FJF8agAqht2HOwPzi1KTfLUETS7bX
O1NNRKqnUZq17JoenMXamoB2Xv6gQ+nqLhnCTcUX3Ilb2pSIa0bda8eB0GoP
QWy7Sn6RSwb7AhP7pS1EYhQQ+u9aCqE2rZ9zVvis6BOzzIPbAzkCUtF8pC+r
Iu5cTUYSoYFMuE7DhDAPOSudk6UL5YP/hViUewUoqC2+EFMjZMQqjbPMfwn4
54/tWoppTM7h+KaUYUhmj6fv+rmt7DSAsNivotaTGYnmJVSCMDntw0BRIj+r
8nl1xdzax1CRJCRtsYdTECeTK75KF7Y7TYCQMbhRJ44oI5B+uEj+Wenl7xWD
fJ+N+HmGgifpXxWOqqb6HWBASXy2pQEBGl9I4YbsxP/ozSy5J4CK5a/RDNSG
I1/ha5NXVlA6CuRo3sMxGF+R90mB52UnaIA1XRcqV3KyXS/ymhJo4/IYSHes
L3CqF0MoDTL1T0eIWIIfLEYnE06uUTkXqXhitsdZQy0SaoRTImsrHogKyJTY
Imm75N9FKiUQp/kYgqLuMBKuHVQcjW7XTYsNhg/wQZPP8yONj0GfrYuSpN3j
LvzLh83nUtW7V2/jy02myNAhR2g1qQGHzHiAezrMRvGcsyOxoygQ18YsVXYM
jJcGJXKn5/sC5njvvStYuTeLFtm+j0SbEXgXohGb1l8TOvhpMVRjHm+vAADs
yQGWTTHAGN/063M6TmVWeseUzkDWcAQ8Qz7nujUEwdmP42p11gRIDBooxxC6
DsfxEeclRjSTaCJnFYKoRXlVJ0c7kAbyw+biEXNJGPmlm+upzb3P80X4lKla
gF/tO6zFCRqteLbc9nNJ/rFdgvpFVCR8fZFgQv7QP/qpneuScpq81lptjUzz
t0XI12NiSDSLtHgill8PL+IRmISSnQzcLND3JZFu9clk9p/5cycCTg+Wjx/d
wjyJGugyQEhS43mxIjP+tRoS1exWooew6Oa8jhMXXuTaV4t+sOvK2BxYxr8H
KIhXOl9Deky1HO2TEvGuPg6zFUHzdk5FVGDbIHkGvo7QvpB9LFWvXR/9LQQ6
emEHonG774G/ryPcd40odHHC5IKwjVcDsh00zYx28syS+KQLoB4PP7iI87/i
FWOlc6aw9EcqkChVWcpaxMripXYcKDSQ5JMYhJjipb4V5/3S0sjYuRI53AfV
2mzD6GMc8feHBhBZNkZlljVFY5pGSgrqpwYtDR5FvhVC5gMmav9zo1+n+ZJ4
Uhh48d7OsVgjj5xZe/YBVc1o9qmONTP1847JzbwTFZCLHqmEI3npeKvfFxyj
ewm+EZ5QdMHr7Ym23Mi7VxH/5tH95yoyd6GxD1rlV5vfA+r2zbCIdSEeSiqB
8jEAeJuxdRdW1FLSd2ClDMeSZRBlNJUc/IR5tj7l7TVuNeEhGP03fzzapP7g
al14trkrryqlD5AfnBZzktaw9y8pM9P2xzjDGnyCMF7W8lwgFBREtldNYbe9
V4sOdT5/PiGvfS8bVquXt/NYwo7I8ojB3xP+vKl46TnbD4X+GXnamPwHbuv4
1L5lfSWwUa9FAW0lqMONrhV8HOhcgj0vuPb6rCPXDQ3BOuLzM27slwcat/fc
gdKauM3whSQPZuno9j7YZrr0epdKwk+9nWZ3kZfuXF+MByz7nGWtD8w5sbnx
vNcBoQ3wl9SUd3LqZGJ5Czt5w10LRvqxicIhnpnJQi1X9kkq+p6rXLZYoDah
N0A2ZZYa9S9bROr+ORAClqN3dP7uvInfSmtlnPARciKKM8R5bIXYc8QTP5l3
LArehgfB9JL5Rl2yDLowOrPiAwjA5VZu4y9pQy1ipDbLitg0Xi6esih2zus4
1jxNqFzIE460lD55/uGFI6HqFTBOqOlf2U3xUNJqowmlQfnPmnvs/kuaT5ti
lqxhvVtob4RtW8H0VlEpaehcjMTX1NyShH3mo7DnEx/zDhR7k1pjM+mpLz4d
HJSrHHNJi2MtSkoyLk+LI6psCMMw7IQIGhwl091Axi1xXFgJMYbzFmkCBfjq
vN5ah5J1K1Em5kypJf8FNMIbSVEDOFOLnvxRHGOxGjOlWKtHSgB05nqC644H
3xObmwm9EJn2G/g8HZy5Z/J46VfkqkoQdOmWe+XDidkdPQCy6xhxzUEW4pju
8607vlihVem8S2wp3HwR+kceAwWcCtw4M51B6HOjnbyx8MTq0QLkV5ixyWqD
qqx2/5cgfOuUzYKQpKMgmJxXu3JKeiMdJXDtOFEBkUgnEjkLLx4bQLM8tU3H
MikjOjKG0Hvp8KHTTN90Ef3HDiTeEOFru0j1J1dv0vDXS2C0WeXlf5C079Qu
VA6YBTJzU4GnwOhK2is6AMdTeHpO6WQod8zUuSz7LpNEubjs2LF/lpheEYH/
ijrcgLL+i3u0FrUWjSU2O24QmEJjSHCeJ3pOgIjNnBOaH9P54n6pTU9T2T8N
A41zYcZN977NRAiiC9KMNvYCO4Y1NROi4pscUwoCG1sB0uAdmomCe0BqLaww
oo35VqJIT5ORGmkFEbajYHT+saITFM04bjuQjabt3uPlcAPp7NMNiaN6/wxa
h7o2/GwOtk+p08hMJeZboRDlSVDWoVUPO29YAUKC8RRgCGtrDMtbUhUd7Hhu
wQMiG8pemjmbJE3aRWj48GpS0BfWkMQVjq+cKXyb8ULS4T/utCVGJXRFrRsp
KUOKyv1hTReYKAMa/x/UB36sVkr3rffbHkrUmjf5vDEw6a8Wh1A3aXjpU6Yk
9eLfPcrGju1Ai3Jkrl6r6B5Tpco4UU8gFY9W/t1WmJ1yJ+tzHlUlDBZXmygw
FLJxfEQNe5r0bec6noaD0jGYf6DuRl4nVscQEpu1vdpM1ivpipG1dLFdRoSE
78PYuEfg+EWYQb7DujaaNA5LFveLuomGNlg2W/VZgjaDn1Djpp5GWET68J44
KMJSXP/4UoxY0MrizB7smno8dCQjLTnJWocwb1CJFzF8hNVaCBna744vY4Bb
xwFgowGL6EqfUNqFeXH0ufcZu3z3vjqLPXpAgGxEdtyPqtRXJVI/RqA+M8Op
IEvfuM01Xbpj/6FTDqQvTNbpWCOWntge4Z/Z5LE5XNlAB3Nn9j1H0XrdMmfc
+ea1gvZUVk7j1+wjqn+y9R/3tve0jvIpgIL1Mx5aeuNkiB48LmVIbTSFjCFc
zkrFzjRHLGi9yBcVBrsK9DJGxy6Y6OB2SYPUAhX1yYALWbwEKy5m//Jd69hZ
BdQ32ndecca6LKwFqFRiHchl9o8e3RiPNlizxSujcli5TXFw4p/exax/D4yS
hYWCT5V5zE1290bNLXViQh+sa8BH/ikdzw+EXY/OIhNQ61m0DLrYjmP0gnIk
DtGdW0YT4qkKWatdIu8OPqMLW66eHSpoxZGIZF+wBwqH1v2ViOmJQ4CDS6s2
SSGGqUUywabMBNg1ZWbVSibirxCKowxcocJodh4gwp/H138YkkMrmCFS+RAU
cjXHPeDax6f8/0pDku9KN8FxzBpH41T0IT0ZhUCvIsGWB9qCsf2/salU8LSk
h5JcjO1UVlof/xaUX7i4kiX4eaDsedcU4vSn6t3i3rH6jWK6Y3vBjzeqo61i
6MIY8IsO94e/HFK3KFtRa8lhXF62ahoCVNz2KPFXZBqtGCfAJ3VQeZSekF2e
pNxDb9f99lEHrIbkU8ha0IZHpOSYHPr1vvNyi86CQ0IdxV+08jPaOyTTiBIe
A3ZD0tL09M9q4agX3YBuXflc+oKj5mhQNa+Cp253PkEGnGxD2YMGbitivG8D
8bGHj43RrrzjHCHRC/mS2VV2ARxEbu7/CpzqKBvqFo1UrhmQzYswKB+watVw
f3YybAyjgnnPG4hpKoJeuj5F7e5IJpZsTl1vk/mv61QQ8Z5lckbCqYjh1Taf
Ir9coaRt8p/cYHAt83++63ZbaqwMtHxLDPAfnIbcS/Qtzv6VGJ2O1jzPZkQP
Gtrav8A3xqLADsp9F38Z3kZxouv4lElACA3CHIUNnHPo9znLOwsCyYyU1f82
GR+xEEj3DWkqfxJEJ4eCfy+lrdt+X7KwOE3VLB70gLu4+wwK+/j+FH51ktsv
AwKvTnhrPbGmd2UTI6wXvQsua2Pq4T1L+JtLd53oEgNdey2+1Y6UlWOx8dAO
vgv0iOjERsgDLXadSElL+0NJniMq9ecSSEbXdgQPjZRiBRCjfaVsIoLN9XDW
F00jTSsJqGjpUzBTnD9Hys76GEIwT5jfYCW1kV6NQ11mLTvqSKx3soVxkxsc
hsrvpJkYUcWi0hYecVd0BkTont+89ov3ab2H0YwSAuPnrAYKaKFe51gTSVgS
rZ+fWyOVwGn1e7VtgqNWEU75ioS/SFXBo/WLL/xMfvwmKFUeotaDpIB17J9r
Qsi5NSA7g97+vgO5RfrXTnSpgLDbQr3mcGJHqHtXmx/qnYYrcJwPk4QSu4iG
7Ck++YqIQH7l+fqu3d3VSu9gmhoM6uJYnn1PmgHHaxyxmMBHp/UaElwdVB2P
bGl1hEGHwEmucsU0ju+Ct0N3o76Ht9dlXSSNVJCY8EShkmi5KijlYlz5yYIr
cdhKs9dqpG6J6zctj5T74qREwHDBfisemWOLADXFWmYDQ5vYQxmpVJ6/RYeu
XVr8nXhk8KH5XO7Syud0uHgLPDIDTNAvHCb1aieboGCaWbv/SgMl+alYmcs9
y8aM7YFdcxI3EE1FnPSWS2bEQkd4qskEyEVfyX9sSDkYxc2KO6Vv3xDD84Mo
mVgzH5m3SQViN3ioG8uuXDQX8Zv82a6Ny+nLGwnrdHRFiq/fl4VYMEVeBQPP
nplcBWfskWf2N/g7Uds+3MiE5hZPqhmYnGElUkXKJ7c/U3VPa7ljM3H5KJXK
vMzhexGQLjfo7xDOjKqVQajpyyrSmzU+oX5X69Q6n0XI5EfwW+vRyCIWNgBn
t7WlCf4h0zNedFbcRyjval+Pr7AM7Wt2tJ0xr/28YjqnKS+L5VSmy4CfBEFi
yvhry4IAv5avk/IpKwKCQrYqUHDCwdZqsEWf8XzHr8xNH0eF7VjHpyNnfPRI
k+/AlLIS92C+lkUDBrDvUiS0O9aWUBgzSVda3DBZWQkZGAs0hRaXcAkLe8T8
lXuFsRA+M25fC9fI/qEzxX712HzQa98jBS+SY1WyYck4vvzlOgDbAj7ZOP78
qoSxaUv94DAAq5OqwcxSPJAMLWQ0VAotUs2mnKX3MD+ALtkL20OYua1aKlVQ
Oj2+/T+etUBYI8UldGod457H5oHoWwS+j6CrPa/RGWYYR6G+PWjIm0sUP0QI
aKdmejSt4NNl1sugDUzDbIr8g27DpX/6qYYNNMaeATT1LFi/dlLsTEtb/udv
i5Efu5rQvrARU+FlFPz7OOTUIslGorYrI2JSAQSrJJehYcmig94vllc021wZ
NbLWsdRPZp0jCdOXuBMcz1Zcsxf5Z0wWfLa7Za0ZFWTBZImeB3HzvhqZUJ42
tYlAICvz3YbCawVU5Tc7xpNEGW9tEhcSDA162kL0jLRzBUb31vd512SIQHyr
J99cvtyiGXp1dVujGHvIKPJTgLDUvVPbKA7SDVgddK4bppa/hkLYl5X6a20q
YCIFanfDbdyGuqjrcuVBu/80Jzeh88FMFy6iXw/iuRYli65yVvN62saff8Fa
XS8os4xisiH31Rybjg9pWuviIayV/rSja+akpFQE/FxRv9x10M70DUKy1sdg
LPVzw2onAkb3Q5oR7hI78bG37PJISybOFkPpVFL5+I65+i/ylptGRjgSC3p5
U1wtuapL+tusxUwXBNNVVnDtA4zezzris7PoqytSGymkx7uhUX/An780ZI70
xskjU5z07VeUvnJX+FDUVqBe7NoPSFMJdSdFHxMCY4ZVJXqNsRzWE3SwvFYR
qFlVKud4HRgUu+hiRROpxkac35y9o6mwYzAa9OgOWQ6Bud2cn2ceNJ8bXOYm
FJ5kHFWDmdJJLM9MlFFzw4fjRMk0kt6GDx5S2TI4L01Xgu4OfyaMlrk8WD2X
pLSpziJMi1HBe0mvfoWnU0xZHyfapgWeB1OXGv3OIIgVUiU1qBAypf3wbZEE
at1c6y5pkbON5DFsGbhepaF5hOQxwnt+zu/9V0IhtG8+eKKOqVWifwpqt3sm
mLR7tp8/IPnBe8rILTFfPTsbbIK/zMEQuh3J3rATxd9ykLmNgvfezJZYS0oU
ASEg4ZmrePCqS3pohl4XbtlAZSLH0LdBotTTKFozOi5qp9s7Vs7TnhOEYPNF
54zNOzAEJGEFD8gRFFkM7H2BJMp3Qc35ipdq5UUtArQJzweUTYTM1Ftns7zz
n82BSzH0TdGwE1GG0NrQKmBptxvrZTB7DWcEdFXcWeNuRnimDePJwaDnOiHO
cO0om0bVA4Mh4BTapf5e/rO5J0dwi5/xMjjvNThEewfTMKLLGAJ82HTG5mk5
TgxBpPB1Ycqzv4R4G+s9RwpgExtw5fEIcLknzKcHokRh1VlxRMAgzQm0bySX
lIGNaKI/BhRRnTUfsvb9n9jWpvamHKdsQNv/fEePd3ArQE8AhvLvA42X9ycg
0csi+W0L7GuvblrjhW+j39WMymAY6KgKOKFcLI++X6+inCmKLU4pJKFpvFHc
1s5o10Z1H/WtuBLCKjlqFCMdYZKf00zfhuyZwTF9+d9Gl5pwVnsDWXeYMn2r
ClvOHmEhSzCBWu2fnUkZGfI8gI2JlkwyGGLGb1U9mqzd/atHMTqnel6vm5I2
GbuJZOIxmFrpK+oWI7e4DgQcjpPkPrQguyQuOiDxdvsb228nlIy8MKrrTexP
SjRYDnRh1viXs4xPN/PNVypF2EsMwnQmoxddvHW6HpyNHMJgy6BvUdQzHOcz
hHUb1aQzmfNtgoAjK6ZYeTiBuOpV55JEdB9rLA+h7uBQtLNQfIn3/o7ZQ73p
hxsSUmC2l4WqmnQD8n4Pw3D/nO6gn0zIFHFoL9mlM+8T909TL2aJWBJwjGGq
kBlTNJNUyI63bztMUr8qvLlFePwC1FCPc/vSlrvlQaMKkf3Rd8WWCev65OLO
VxPdcInT3f0Q4JchSxhG/GUEnfCkw7qgpkPVzZDDVy46gHJRnks47JtW/O3w
o1NrRkfUjrPKO5H5u53/nCb3tgio1Zn0ufPV+Wi+Ej4oQdP4xqkywUwjUfT5
mq9RL9O0Nz6EVpSyFL6Tqx7BhNTXC3Vhkr1S44J1JZKP0AeEZ/p7RmtNVgk0
ymAyb8nBR/2HQgyPRGUhAl0rvoSar0A4vfTLmaw7SFwnCisL6+yJn04pD6PE
1RvhnvvcbLfSsHC7FpgzIs1x4f62ybagBWYqma6RwOKnIYKFal8NaFrv5q/b
8FY6oT/14xoHb1dPFwBkSH+uIoqjy8dPIDj4PrsE74h5p16DNx9rZmIkeocR
WV9PzJslFOb1ZDLuQc3DOPGvxRaH5FIvPQgTpo7NwTOCueJh9m/yFJgo3U8h
Y+/3imJceezNwVgGrf05OTCXcRfnMD5lrkCOz8YRQA+SClxH69XUcFHhvJbD
Gz+u2ojAy5TSfw4LWPOtNXXGFWAnrTkynkyT/X+5c28T6DgBxzMZW0ulzahZ
zj0F5Ql1era6f6j2Tfv321yhd98mx0rQ439vcBDZgwOI0H4CwpU3N6HIz2ja
uWWX+/Ls9RDRZFn9L+DTyxbYxr3bH6LZf/a4Faf4jkK5yCNB4BnExNShwyVQ
+6AVxo9QascvTalqU/gUwlXFnf3Zfs/gIC9IcBqmz87MMcUHI19YXt2jVzvu
7IUEZ8Cb+YNtqm98rld+izb4x5ODlo7uMxk4HAv1nV4MMK+k/6XChs964fL+
rcaHhp6LCwTdbLdfg750AfgZihE6XNUqwOjnwHSG61um/A7wL5Qpf5VqUff5
w0y0zsR6yNXVoaRTLQPceskndunNm4NgWlLLNqlemKtZiSJ+5nhoNLuHDs4P
y2QBAUPKyj+UgR6rHnasPyBqaji/AWgSWUouyVUvLAyrJ0Iqh/tZxfv5P/mY
9FBtcKsYZfZG+J4IwK9SfEmORM0ASeX7Nzqskimx5YWwWJZ3cfy4ohVwLg4P
n24I/CEVwfrcd5jK1Gnvc1U5zynZTe+6ErhC+diJYW98kNNOhAT9ox6Yx7j6
rZs08QgcJazNwlpWxVDiYgdxL6YaLEP7qJo6dteSc2dh54KH4BWUuyWjJVam
oQzQZ+JN240T76HPGj1eNHL6n1UzJXPQ+VJ6LWHnCG2A15EmQwm0266pDfY6
b5QdYJnr3tehGbSHj6I49iBzylwXzT08MUBhkP1gwa76bqy29fAOFwZBDcpf
XdulOyHt17/DCe+Qh1t1SlGsAxn+Bs+vZ//1pqsHm42jjUkXl9w5hmupOCe7
oebFduitZBFLqeXSFla4ZtmdX1oG8t0DJXGBTz3jmkQDs/DHXeFpAWmJZgI9
SJqkhl1wUPmhsp3UYe9L6ArQ2iG1Be/2ab5n0hasCsvN466fJmMdsAOku1Zm
B/dRmTY8w63a50QjtjS0JpfA1TvCvLq7ZS2qp2GYTU4qL0sUCwuHB4Dy/qH8
+kig5OWrIzOGWLDxo4utiOz3fhdRlgLJmQWaDQka8NJLIE/1ue5qvKrBl4DU
/S/PRGnMskVtlgvA/Xn9IMQXDubp9LSXtk1AZoi8DG5TU8S8/zU2DDL3vnLX
2CDTZ0ou1Au1rgsXVKvnX7P8mn8u8i9MgPlSdzZFja/ve70zlu9KW21+J5MF
feEtXLFGC+NkLlRSORn3B9SNHCUpUgWWMlmJUWeDrXifRST8MO/WqrXzpwcY
kyz4fzFw0gBnzwPbEJ6t1mUEH2sjsl83/wYyN56N/b2Jh5/Qv7ncsX3RKNEA
YS5pdc/+5g3BIGP4nLRogEXHz8gjJyqzH+ljcOK+LCMcNNtT1yHOdqGIytPA
FXFNoPwGeowN7ZFuXmADrdjMSuNEZ+prLA/eWEWcHth9xBj7A4um1YQqZiW6
6RFOvpxUdQjJnB+GNibnldp2KBQTMwbnSyK5u/oLY1yApQi6szWSg35xOioI
LkXgVjgTl+yxswtxjeUaURmEqvu8kfpZzbHZ27pu9+U2QEYHpdRwR/gRjEf0
svEfewkbmfRedaFOiQnAUSNyelmtwFpkIfykP6WC0pPdYTnptUdQGN5SOSrT
GA2NevO6/uq7aahwNNy/OKlgdV0n/Im7BLpezlmHOnh7+iakr07BjT7WyCtG
p9TUgDZIuZPyP6/Zp+nLtOl0Yo8XQB+tePTPCqy7CMImdlUXJvUmxLeovcWr
Elg73tdV2KHyJHWZqtqb5pGlfQC+yOIsKrUlXapduumvMCIto6z8WU2G7x9j
4c48TO3x1cIbXVTq99iiF1OBnkPRC8wiaZg/nACBxhZqZMFizetI2vNIUIEL
Ad2rsOnwugFHAnkk4LDtSm0ar4I9/4c+GacnISh+XMv/zyVu8NWiR9b0MX0x
MyjNom6JUUkTuOvtZOWuohU2WnsEJEgUl6frUcGufUWbQZi9OJUajrxyqL6B
2+cfVjByuW8ZYEgHpQ7F1FFnlsRmSWewVFgYHUxCk6Dk4d/5YV5+p6TmuqpY
n1wHxNwFS7be+vZz1DZOSP+t1vrAs8H9g+4NIEbHf8eFzOjeOidgltWpQkDR
5BqKOqV7j0tkXqo/KZCDTqSsq0Ipw4Via+5menx7X15O1S1/rfYJVK86XQY1
eARFtnBnzPQ7tq4aOMgHOcItN/t7ilifnpkXl+yhQA7Lp/v8LhdTd6T5DjuP
Bq7O/A9tF9TUvlMJv6J4S4KxRVW5Q3gsx3/nH9uBkiLhlqM3aSgB52FhAjPy
Oev6+sueJhsKXeY6ri3jXzFrHj+sQVZkSZ76HjN4WlFUo7D+uJ9Pb/+VzwSW
qVWpXEpMbWMjbCPGcrBXnTH3ewY/0sQNEb4Rukm6GgB0EyfXn4AEjtngUizf
09nWLJY1iPSPH+MQD4FyonT3qG82frWXNzBp2c3AMsWYKtykGN3YtpCKdM5y
TD2TxrgvQWsq+NKb8t7YxUL2QDE4jpeBLMoaiINQMWgTt2DFe7lqjDzeb+kS
BFZRDpFjgMERmi/V48r9dvrkq8ZozYTdzSR7LVZUoM55/2w2wCSMGqKvouiU
ciiBvvizj2mqgsaQUcvD7aWHSbIgwuDsbyEcUk2jqddGu0ee1ky7tPVlLD1K
3Uqk/AvsnJ9PCV5ollH+pWXQSTOjXQn2X1lpW8NP02UyTUn/jcHMCW/CAX0y
Xvr3bjZMQxbNxSLU7lxWAsfHRipmlrffe3sdK7tVpjz0rWVb27Mc0mNMMMss
dM8dBtEfsjGUl5Z6um6A1ELTA7hAZRSFxaT81KnhgE96JWgMOR8zVMmeBpU4
jia/BCLX9eyJWvCrFsCfSUn8y4bQaYvvtQaosJCa+YTLNPIvTyFkdKjpj9yX
4ztXO7E+e7qeVduuXnRZk3mdjDx5dOCdcohjciJJN9NHZlyZkZJjnL++G9de
AQv7Iz3xln4PdZgmsIt1B04UOwtNoC93oZLN1NXlIvopE5idgSJWAA7ezsVX
mHVRC5ONLX8AU/ePu2A8luT/C0a2qtof2+S1cMIP0Ui0Ey7ykZwxeF5SuxEy
weC0KkZ6TLlsGtZBY/9XgzEzZW2i350Ob11r0cxtVVdrv21qugOOpzaEI5n3
spglJDxR8EnjWC8NST4+VbU8ktxzVa5kh8g3124vkukyR/FUFK3t84+W16Q5
/UmoSoT+i6Cc+zXAF31yYs+DzuHmXDxZ328LcfoXTFFVLOi+sdtKtCeeckGR
Cn3PqXXkZrfZj9/I6RUEU/nnh4AQL4FsFEIGH2UKrBOJeGq28X4KtzMPiAbM
P7Myc2RuqWEUD/eTRhLhAeO/YXUNzkVEx/5gPxbRtdAXdEaO1cLYlzytI+/T
8MqkwYti7d6BLgJaMA07U2ZA0D/2OVfj6rF/rBGkXEBDfiHZoa1BUEHKRPuY
o4QHDAPGKvGDr9OmricQyJxVUegplSvIPvWMazWbUgQLgh0/Q5gqBj+f5p91
98Dzpwt8L0JsFm92I1Y3w6Sh1bsMb2f0nRK4bdJja45fyxXdipbJMwYMJ/s/
L7DCFp9bOkAvwUJNG7wZkxcwL3GSFqdlmT2HLaRIrqyNp/1TBfTYHfa1kfE6
zIWZ8EqrdMLukuntQnRqtealVHr8Oh/OdgAh6uCfKj6mbvnp6cc2AUFuRXo6
ER+d/SIWTrErCUwI6P1LPeMkE2oouEXpIPZfmqg/Ax1q+QmTHTQfQQ/X6Nri
x56WELxk1YeJrCOucxqGH4nH0gOr2VD1WgzidF3nF9GWxTGMR+Iun8mf2Neb
8u3dKco8uqvJ19Hb+LMJ2aplCeXHfK3F8zNuCuMCcBhIeKssth5CsXSs9z2L
UY8ui3l8pI9kW6SSE9DO9T10dAYQUucBWX+7w4SHI0HD0K7weNrAbahfQsx5
zq3JI9oMs+fPVuB3TdjdlZvSW+CRdgVWZEnmTLNcOND9iDAhTXowDaVXhKzr
5RZHbmRWOFg9VJcAi2xrnasFppIICXSsSZvdP0VSUFOxT9L2y21HqikMffpG
wgzgKG3Rn5hVrbdK9tHK8D8C1XpLlyDoIKeLKQ4KseyWQ3N7P5ZaOFq7rG50
51ZF1vESgIrwxQUD/HUgK5QAzzseLOvSUa+yh7PUqyNx1RJrIDijwrI5MToz
vErRYcgG8JbrfQd91v14p2P+2X/tkYv9Sk+Ae611EjL5JDkqVpG93DRBAONo
y8c9fMjyy/by+J1MAg5u3JtrV/mRPEnyqs40w2gGo0qd7hGpPrRThuOM+Uzj
XRt+bHBiPtlQdzQ4msobpgCvWYSm8pjM39Vq35w4uQT444vyHX8ddjcax9zg
cKZ474gKQNXwRkWAldX2a3PF3hSoVjsVCag4k0/O1LEXeeMBarw66cOguNYp
kWoOQ00wEFZc7Eogy8tu9w3yNbTpakkUctCbueguC8igzmTY4GJvYfxzmEoA
lgEXX8MsZqYM1QPsiF09PnjqlooIxbJDB01GLU3Ff1LRHI3IKrV7eqeYqlHh
BMwwLFzp/sgGoaliQ0wNWc5/6fsHOyBSh1Og3UGpnvsATb3GJ431p3eVD+PQ
cIizpeV42Q7xxi1dwe/9X6I5q4nc6cjskR2pLPht+/UMcO/3muUHO5H4o1YL
bSNAmbQmg4pFPvsfRRx4gt9STg2Z+7cHcbP3Pgs21lVjsPpNVCZyfxZTFg8e
vaRKw1gEgGmvaRLB/Pf88vrNEjMcjT/3ORtmRsz7BxsHIysTQ0smYDgFfqY0
8iLTs7M6q6QPGIA8C4+18exd3bJmE8b6B4lI0ifG1CPx6NjaQRC2TvVePzeS
jveZRrSPchmhVjWBOk/X26ghKYU0W1SvIOS3cXv6f6xBaczWG/zUKZ20Uoxk
sRM4MPrMPNk5VuhL6rzt4ZGiTSD7h0AQlRKFOGLY4JudqeYCneGKksefVIN3
h9lm0tn3/QkwX7Wyk/nO4wTRlS9CH6jTRiBb92eAgbQeBnu9GEECSpzT/0Qc
MuCb6MY30rdMSOwWJhYrxjtMx33ceLkXWV73FBxRzvmeFvbTzedvcK76b65s
EHHvCc+0oUcfjJwXJ+Fe+lcLtxod71L5XjjaePLhr8wx8NOw96/5XIrlZyM/
kIunbwOdnz8zRHTzBBjCJIMB4ifWuJJQ2PqUNfvxrxf02fiqyX8Cfc8Iejie
Weo5OXqRJltm1gWD+wmdiRhBwmeiPlihIrmU4VgtFUFmfiktAMi9zhwg/l6B
f0qKIBy9uyDTJZfR2iUMq+HTTm+i7VHaSwVeMIfQ0Pr4K5j4B6yukh29UYpU
0pSuP5LjRWJ95xeC2+A/ykyLrKlCCcwCCn8d9+b14U55zLIVpdGBcR4XpCwq
dyRofWpW5//U/gj5I14noMxu3oWhHD3wQE4z63ri/TtyLzWNiW42omWFA73G
1aIQ4zkpywya+LsFnOSDzmYrMH+hLnltnKrKSPXMr6yvB8yQpeA3xLcEe+iS
hbx71VAx9wJcTQ5YvmLwuw8YQyPYAW9B4d3gmT1f0Lu2s02ex1K8Yb2/7M3Q
2zvJ4NsBcxkfWPtp55jOK5rvOAA399LKHWirRnB8/K5DyVrfMv7c/2BR/dIA
Dzi5DduVtQloivPgRCNyrd0mvaAShXCSKB8OnyHVNSo9j/TQwOoC/Nw07Lw8
zge/RMa00vPRDNXButvBRQ8JY3QdzdID7+lZ/7l+2vjbhaT0FlRps+geS+hh
4nz9BR9qQ/oCtozhzvWel9pwBwqZmkpqdWyEeMZcZleAzfAS1pcbayOq5hgT
sKRMet3WzEPyeOpHL2VwF+s/58XPYVzbW2RZiRfFS4iZn6vUP8+FSzv3p4Ac
hAAUow6hZ1895gjcqslhjecgLWySRQPQGTLbaVJVI7GdLoS3/oVSBE3ACnZF
l4TJNVekh6U/0+AtBcOTyBYYD4Amt8LzcRHaM0jF0he5XIGun1A4i9Gvs97x
QD6ptqzJuVCGcSwf0tYGXrpUVTh9e49OK74dRiQOe9iMm+Ne3o+dOjQ5C/LD
SQcY7Los0JjuUxLZDp1A/z7bQN6aa3nbmmw70EpfUzuD6QQz7uM0nmijisgZ
SP9c9tCvK6e7dxYS5tbzIphLNe5qUy1aYvUYEJAt2ngfHKJsGeZypmSp5PJT
Iy5DCP5VXc9HaUJzPytVZDkcm9RpFDMyglzqHOrLsrkTCPgOgWhP+g62iaaj
dEO/SFGSYrwHXLp145U4V5kzIfEmSFRtD/HnRUGSmvxF0U095SiQABZP/5U9
+zX4u3yDEvAzyy4nIF48S0ImnXiFgfjELNvGvmwtz/ToPzsiV+vPO4DWUHz/
w5BOA3h5RtJnZGSx7ISoLfjbXT9vf/pxQ4zBaJWRwijhzv1Ykuo+VOr4/80W
dafi5YfL/cfdZUuSGRgicEJobLLvGq0kDU1Lj6kiPfl4WnHUXCSxTHIX7zlb
E+nfUy2xxx1Zd2aUvPbXxZgbAmLSHrOjyws90glM51GGA//p8vMF4thdqDxI
UYYbJ+e8SjzE4x93FuoRmZl6LQO8f3qOirRowFM1/DAw16eRFWl5q+YXHZ2p
yrJ6f7ydfvKRyJwN2pL4iAU05x4e4UrHn94DmVkmDzz4dAk8nXt5Mrlx7ehS
IxxfpgcvhXaPldtMKECX3kw6pfFR5aNmf82RfCt3v1VPHLsZPQBzoG3tp59B
pM2ctEn+PklpjF97Tq7iv04wmWVszGLLn1yxgyMnVWk1PDyUEG/aoTmY4+RS
EPXqdbiCEZsKioK/fazWFwtrvcWavdU1KgVlNGYCB2lK+f0kX84ifNczF42n
gjuCORM/OhiZmSDmDqgUoJvMEVt0eIDnHrZrDNkqcomC6sQ1hvDIFPflIS6t
lNe1wiW0ce2HHlCITLOYp8DA/TL7QGNO33MJ1uWu2mV3LpSnFxLUrYfkd0Zi
jQuoJc2eqbkFCl5KPgXEKOayy3TRmMJtPgr6oi3a/y7kQCkOSsywskc+RdXQ
bMev7DzAdpJ7dqNZ0/3+nJbRadTQEjcbXsYwW1ALc+328Ujjfy28ouJ2YbcT
crlu47wkb8sOvdvU53WYtqxLrIrsL7mt4FYfV0cgw21hTc49DA+05JQQxsd9
3oqquesTyNvWKNZMvmAP3sV5CbicoGcZRIeQWPzk6J8bsi9mW81/Y9G0dn2U
5cAgjMlM9PqP+0IzcVlXKalWWzmHBQdAaJVIheQeoymoKdsl7V71aGxCqH7w
E9FAt+tCT3nqCZXbtGVE08fkxzVJpAht371ZXJseCVqTEqLjhykCAK0Yr0Xx
A4rqDIqGe1BDtCG53bWyJIsv7nVEje7HDlnq/BREWt8UtwjchEzfa2IaUpeg
oN9DMoU2SRsg83MBir6z9LxfyJQw8aH8SHlXMHIGvzeTTBZY3V7IvYJ6PmoZ
ZpsV4hzpFT3KS3NlCk0533e16tvSwREkTQ0DpS8DTuipo9U+ztl4lrGEahIH
t/dNePM7ZQ3fK7JxyYehDDEOswE+f6JOaXszR+vuA7nK2vLdP6ERkJoCEdYL
2P4mbR+Je1ZQRHoJOHyJP+aC8Vv1M7jEBoT5Wt8El33qb0wMC3vWup6tEqTw
pg3ZhRG6a3sy6AkXaBTYEKJqH3l/tB7Uqp1ZnAqBeIxGubLl4HZ+lWTGrDIR
V5Wj8O0G0r4E0E4tT2x+G9pN2Qrgkum4v5lufUApBLdh58EY8DcjE2g5KE2E
H1tkhQbMVJDEyuSkU/xjeoC4ImjRumGg0TpmySkDGgIYyPmTgOCpxxaqpSp4
ySeXBy8dGCgQvH2oBsvJNPLXCvxPiMXcSvUnbZf8WzDoyalup5ReC5Obl7zK
kHmm3AHg3X4Nr6YZIL3W14IPRzDE0mmsnyJpFagg0LKu8k1JDWZT7n+lhSdr
YvPKs52jORzu1DZ29iZmwuOv30T40aXMfA40X+Tv2f1jkJU+H8hO9pHj8aDS
0I6KWmglFb6iabSYNhHqRJhEFWQ3tQSfcTlgvTOFXul63+MSSWCzfpOSRahl
LbYFaCaEqbIFCRRhPNpHNpV7t3gI0S+y0G5OkRYiVy5IiSYfe7WFJTEaGday
dTm7rWF7tJPk3BI+kDaQ5qsXAXvuC3k2z1t5u8rIM4NCHfP9RCXMmZ6jcJ+Y
01iLm3ygO99eDCWkdBM5ifpF1eno7ggF7CrkA27XUR97NL79ZQ7mTUddZKh/
fFEvnVG9zGWV36/raOX6n4oj0W/5X9LPifmZ2EEMCAS3bS42NgkkUKMu+l/A
iVcZsaHZ0sI0ZPBXj1GBCm33nsEwwWiiXmpMs1QVv6NfjaULthaxC5A33YdY
JOvjd4V8ZNO7dkeeM0YJnCUFm6OrISiU+Nk2fZ84ujh0ZYRW1ibEX+6XtjYX
7aO3TFYIYzgXoQfPp/PfkJdBr2Rzg3FC84Pgqj+8OLEcmo2wIvuW0yKEQVC3
bbtOrqymXKNd/X2bCZq2Zfv+wzK+RlB1QfyyvvEvfAOTUKSVdHklrk+JBQlp
oXeyNAlTeg3zjUfORVGCLXSWpmdJ2BEoW+fxBb5zTcuJl+C8nOKYEJ08X213
RdsR4SnGSrJF4ZbYy+8O4Muv9lpk9Ltw621hhCfZqqPs8dVMOirmbUqDdyrJ
2ErI3p+hqFy0wMi3rKzDUri7GQofYTQ1b2rSGaoA6MYCDPZh10+3/xo3V1sQ
0nTeI+pYMZ3BZvtOEiwIdsPN9UcA5t/Sl57ofWe94eGwsjNzykFD4Dnntesg
o7bCCxc2jl0eERWmvZyDAg+teIDdu9aSfYvBRN94OQcVWtrSmq458fW1Bcxb
OhYSE6qBGTG4XomcE4RVccJOyjHBm/+zCDj9Fb2NU333+aBu/qVWK+PG88CD
7GmUaR4qr+reizcOa/efyB8fWm/po6Lzxxa76IRZSQ66ceByVB/fT3ov1vSv
+l/ZkTuNflHJ9ov2/Ulo/729XYRQbCzqR/+1wH9bMEyizC0AO97bKQ824oGH
l2E8lwn4wS4HURyiwlEY1/hTke6fCr/gXfMjHxKQ0CHtOXIpgzHlzU10e0+T
eb45VcoQe9/L0upjOkud8sNytxVk4YeN3o+fRaED0M2ERKaZFCiMMlKjVbZM
a9Qa6fT9Ei3ts/MCecij4s11voCV8pbdbeXJaVEMUz/b6dfHdms6PM8Um1EX
F+c77jD+XHoFh9aFUKxNAudAWqrFW6bx/N9VCYCeBDRb/RgE5e9ASQkQ76mz
erTMBjtjPalFs0DFtLhwrOhEYEyzPT+18S4q/pHBory2A6v2MARwX9PmThO3
2/53wAJPs4knM8UUhQ3JfVfCeMMshfGd+ivmRqIanLwfVp7fIzOhbnFlSFGX
cwN/ZY9Gtm+e8ATtoPmJYRv38v/vvztKFCV2X6Fn+LI9j5iV1CqeAyasyv6Q
KlHQF1w7jzyrbRcvwGW11FxzvOuQ9AiA2JvDAw7W4VgGXj97v1dRYWhlGVer
lL+0zvt9s4ySh0i6HkUeBHHmsODlBnhrP6rHX0OMDipVXhDyTcBnhpmgjMwf
EBFSWjW016e7USYGqNcMRA5B0xa+iUZzyrmf8+joJBkMMQJXGDoQywtB3GWy
r/pxKyBFg4YbC1yD20HPpLksbJfvh/31pSTqnUnWtVFI6U5HWl0B01NqdoQb
6ESvQypOFLSlpMBLkuSeUdbIDGk3xXRrw/Kj4YtgKpa6V4epiunEOgiIguJy
WFwvxjz9yAGgh4OmzVtPvacTqpCog9kD7EMF5gOxakF4DKv6tSO/HLmksTOe
vJWQCirRLRlk03dI+oA1xtVvWTRIFGfHfm3jAP1AvWm4RRbI/ufUfb5HX57a
JtV8SDV4ktVh2YdzCThpzxMdyN/HM97X2flUxEFIjucV4c3UIebTaw9kvhku
kGbjTAD7NNTtGWgtOPcHjZWtAqn+Af5rtVG8u8zjBmy+g1ThrjPybRZXOF0r
pLquO9/uCSuFBtz660z5ZnnBlEFaHImijjCwQ/1PcXy6de3o+nBDYsWEwfFj
CFia/jierCV8DrqPWS97p7lqCt7DtodJmEvgi3vPgaewr29KxwccaDFLYXIU
9XOIQKGn0pYl3yBlHFeIgm50ML8/Pf+pgVj9u75/OUk/PuLZ34IhO5eoEEqG
qKvTV9bnamOZR9FHVE80FD3cQcDXdeOHQJyS750rwK7kpRpbb/M1NmD++VRU
zmF4eMKJMgUiE57iwbU/vet7QvqHveX0T/Y64gbp1r3KnORAwe9Nbf23VvFZ
vsR8jbalX3lhqTAwghbLrBh0korJu/NgYQolkbdM6HuzFXgDWmeI69vD5bBi
/fTi5Z6sRtaazTa7S95wpl9svPZ1I9RDJLoSu1HhurbXnQU9Ol38ACdqfZlJ
Z3su4I/1y53/8ZLK3/O2QPz7iB4iPvwEo9/fi6CxwShmoX7xxGNgO42NvrgZ
QP6o27bPN5vEAHDyN2xCWYujUKRxe/7i0KBp4B2JjMWfvFKwxjLbmOdYlmcf
khz3TQNkK4bVG5wZlu/rheGykOIYHXP1lPZl3VpFiXMhnd7nugwepqMC3OHp
zw4hSD7En4iTc+2l/TlayVVZurGFoq4bIMzg3a8yKe44s2wsTejVsx/i/laY
Z01hpTsN7DmEnjYrJPII+Tw18z9Wl4s/8HQvMUBNczU+BTbcKjhVk4bosjod
A6CQ1gIYS+w5Hg2UxV6a7TqU4tTwOegIeWX9LPm+5msUlExYb5Zh4u988BFm
QCogfANnAoxp+jrlNA2cnUzCBvJ1KI9jG3vj1xHkL2HC5I/3keGqJgQt8Hku
7RY8jx6hYxQL6FgoTJZHuo7JwF3VuUfQ/lAmwqBGv+lB3glT0WEdBu2q0iP7
RHObmQ4NPI4bgOYQOSLHzg9qSjk7vxn+9IM7hxoK1XbS9YtISXmyywZRX/Xu
QQ95tYKJe944XluqU72fAqcd8Ei4IEZnzPcn3RorD6I4dKPMoMZB0B20RLko
h2DTtDqjfi0poNQfv9RPEckuECipp/UktTd2gq9uIyK6byIV3+1pakHzXyk1
19VigYL8ON+EAw82JbrlhYfsLRraHLfWVM85RLvEop9P9CVS1Qms9+ekgWZE
qZVf6OKPpkFrWwhYftJIsiJsYyay0D/D8L/yn0jhFdZudjS0649vDnQfRicE
uoWg7/fiuQyXhc00+l5xzd9iDzBSNjl8rBBuIum4ibL6CWERL/qHfL6CX3Oj
Clk5CxY+T++t2f9HMhWDjbwJKFuga0/nBv0QkyOGXTh9FHc29rkNK8pGNWv+
ezrsQYAVPGlaPwFW2FrikebIEZaLWR6Yu1ax4P03HtTreZb7eANAH18bWnE0
5io7ivJHjrdr2WwNu04R4QggZZL8D+zI8kLk7j8mMkjFVqZwrrg1OIoPTvwf
sskfKpoZV8iWpY/1xv8Xc//qjwGJYRklR5bAVP4e0B5lavhDFGkiUv4OsMDj
/wtfmSZoG/IQGWPgNLzbjgR3ts/0+Qah6ywJRO2yZB2zNQiKxbi8fF91Qf9T
gF569L5YvXg4gqarz62anGLbB74DR23Cpa9jO7AiQktIzTkum6AiZwPqB5iM
tC4n2PVYntEenxVwE+ha+EQoJ05K9VdocE7bbE6iC2TlSH+s1Y91hObHdOj9
Aq1jJVrXq4IfN1YQI8xro71bK12/VfN8WZ1STiy1FWunl6VjLeKuQ0CcrNQt
cQ9vrQ4yeslS/+TpAJs6eMyHpVE6WEJkxd5JoPMxCsikTJhDsmph3cR2out5
den6pNJtnQfEcqpo6hMPsAQ4piw4dlMaZbHGkJzQNrlLPhQXSqk99hNwdnPj
zpjJScxQzqZQZgFu2fKHqNVOT7ZvENFjIBoJkXKim6wXxBvDfwrVbpLEMPLU
e1AEy8NTSnOJ9+/5TQ5qDXU2IZoQzXktdiGx/wIUiiTdFH/O6v1osqaQG/JR
oaZ+MeLFjhXXuwhYxyNu6z/+QPnSHJNWq8p0Js9g3e8pC4RfkGvBlc65ExMQ
RRCV1tI+sKJuV9c7KsgZKYFH7dmlj3kyG3kmzkUwds/7WSMhTZNxbbUjgOS6
CzZ+YgPfy9lEKyWM7ov8isru0680RRi6Y9B1mL9bxfw87lrU8A+Bi0KovNiV
cVgJ7R61ZMitad1OXxyYgg5oEof12vg5XQZsbcCmA2+tgWnC/3OidY9lpAAr
YY0HRbNYWXcnMN+z9spiDUrQwMqH1f7VJQ9Bxj6tK/pw9VeREq4VktYa9WGN
pmGoNS+p10zMlRzzoc23JCwRnnodDL2rRnjB8PkIu189HIZA1o556WLu3Ga0
yU0VH8ObuQ0a8Ms4yCRe9X6I5Vwo4NF+2KjGr2eYmM1oX765kaCjGyIP0Nlt
2i822L+iVOiocxqZEeHgQDaZx3P6RC3DJzc4oafkcH1ozlx/EBobdaqd37rm
2nKxUlp7ywNsEbHQ0TIa9WV0O7SjvCS7udsXYQeCjhbPsDu14c3QzyAOYwLC
GyaRzcDpEGVra/k5yPoXzf0VpmlvyNw0zyE7cnY/5oAvIjsnJYCmTfY+cWbH
FqqlBWNOiIooIjwSTUBl5UtfbVOsx2qhXuHexB/o0eyIHOFldSAUKNq+Vm9R
dZj7bzWNH/KNtrWtNDEfn7E0FDe8DduzB5BI0O5da9tgYZJCKGcsnZxpx2L2
9nGESsVPKzYYehNmK8t3Mc+rLqykpdg7PnuYq0dROnV1RAFjSpG4W5rs/8Bw
3DZ2+5+vOTgrNJrMwpgtGPWGygaIT6nU3v8Fvyj/nk572UBCPA+ELZR4DLcG
Vq1XPTj5tQWLwe5+jJEHmGtyUVZbQEabWJzoo1EHH2sM76MmeNYAdZb/CDX6
R1EpSzy+lE3sHuO+CvMZr1yME1WrerDMEkxgA2gc2122gfIG5+7OjUoyKV/D
oYj9KNupRemmVrS89Ect6T8c8UwQ9Z2mD9QZmRnkAE+xjPn5mhnY9x/NZ+vx
zTaOa/qNFeTn+xRSIbY4yvEDvKP8tx0saJWLmI07SRhfmvVYtCkjXBdltbAm
Q50Bf2NPyo+GmLYyWx4ZtQsytlFKEAY4V0waWNqnYIbSPi07Io9lIwQMbj59
fIycm8oHhxdGgumaiMc4lQjKsVPn0fiO5yiPtSYNnUjqMccNSRRkoL1zcACo
YvN6LYHzDL/n+4B4PeF5sjm/GvZVNlq7nOu4W4bXhlG5aoE1JJesvDdF4Mzv
q2poeZZ89qFIV/lxPOt5hVGP1nRFiTfWC5qacw1+5hppdZH5wSRmaox47H1M
LQeoadbdBMz1eBSzzNDc4kRK7WSgRmMXw50Om/qKTnRCcvrmKDUF5gmucc7z
SEBjwiSYRw4pS/JYjKIX6A1XgYlcBc61A8RLGMpdLxtfmbxLwqwH8RYbAgwl
VCjsJPXX+1sef+UdW1Ko1PSn80FOlUTklIdzuYZur0MXDJTzL62EQu8D/3kt
GGDf6rgKAdGpeOZfWEw6yu8/buVsM9KYUQsAJADXjA74oOJ/6p6OsKGt1/Em
69sfW+Eso7QxGYQYue1lTzVP5FKIZ7fxLcfwbdoYIhefMm3FN5w2pe/Y6DDC
O/1Amw4u6+dOg+tihniTvcuniicS4O5PbM7fHA5PlU/9sJbble0jXsdcPZ1h
ipmRyDUqs+9rIBkVG/T1LjZW7kfugZWEFPeWFx2Q2W8v0uzFP1SrPaVA3N7k
WQagmsYL52HWtTvQUXs0iQggmYQGAGTrLpqmmWfYZPX+88BlVWEnA3otfDs8
g/cXBcMaXvljRSkUkvxMbOnzEusI1X8OP17O+cSUwNeCm1T2EZnrvzSQDCds
a5lYzYFSHcKqR3n1kSxZHK6DaJZm4TBWr7bJAThs6OSa+gCE3kxTIxn0fI5Y
q2iU1QKEGXss9Il4LcBxOcYHFCrpWdJdVe1hp01DL6iJ8CIK7Bvobv8WvHKo
yJfgoD0Fybgh+g++qEZkf92OtrMJDRHa6LpYouxx3E0tazEQGDeqelLI7j4p
c+dyKzBIpPpyLfbIQFZ7GsT0YvInvy49SsUYLg2G8go7al8fEAqF1p1RNhi5
Z0HRONWGwH+rvRM3O8x1+IeYjuUXiWWLd+LFHYuHZwZQXU2u0i3FK9DqgvkC
1yvfdI5nPh0mUR/mNVYP3vWtVy3rEYwsYxJiPgP+A1ccaEeiLaxqKijC5cza
od4fhzasYL/Cj/6CgzOrC22rqoQyWcLsg6AoFXKb+Jwf35deDLR/2pZ0+/vK
4/lHoR2jiRFI0o5i4qcjhVB9Qgvnn30bhNbWVZ13amad+HoCNAOBPuvumpcW
UaSxJCAymTxnwX6zd/GBLaEKgGjejLJk3pIC6prsXCM3G0hDx2CcE1S7i/3y
gyJ3UV1R68dWQ6Hea/M8jaonb0s1oy6K89t/ntkSwGFDoZkj5PiK8zFRcVvo
CiOvWgG7kaYLCnDF7PPRvYBm305boj82ps3fLaeGn0mIB5dcdd3JYG5NwREb
d8npon+bOtJrB17jYKag0FMjzeXUavN/EMn+jvY/7BEoFEPsWO6yefyHleko
qX9JmDKL+5GwRbhV76+FcsJOqb6zCzaW1EzVoVLUDQinkvnhn8FJf57rU7CE
py0bwmP+KFTm0RpH5cOOpb7Zp5lF8ks8/WiXbBiy1TQgCdkTErb7sLw1DuPV
A1N08pa4dsMXSU4F33AGL0tRxICVTTz3j2fiQp7HwGF8k5l1PJNNcVl3kna1
y2rKnGdZ6CsawXc+6E/H2cHnYQ3gNVdd3SF5WHCiT3HKlPzaNdWZ+iA8oEAy
R1tKPC2Wl5anCJ7sfvwUvZK4+1QCoGaTgNPl3oYrl6T0XRw0zCzFVFm2ogjQ
zcyzTurKyawUusq0i5EYpm7XavD+5F1IZF8AHvnJQUHGSfZ1zSTNUToSOEcz
eygXTh/XS4CrYjoU82k/PTXJxo22hTLypbDtrnYAq6XDMPRB0XkFHlMDII6S
4BfVPCnmz6X9oMb+Q8jBKFJjmhGbiAgfgbJ2IFRQYdcE4uAd7gC8rtiP65yl
djv9qyEYdCMQAYrMwqzGPn/Ox/w5woHO4neAWZJP2eTy5BTGtj43HsNU+A2K
TJMIl7YRMGIiybbMcLZFCJJevjTnmQ0gjlA2/cFkzdger/g5sgy4cFzq1Sum
1Tedu5gl8MOuY5hkajQKa1K9SOllkhTv+WtVEO6TbVSIxWI7a5jNN1v4ERWF
nFhK8nKrF1tWtf+HCMap5NkGfD6xU3bATonk78VzeYYaHh2T6paWFrRjUQIU
mMUdCI3HiiQYlgefRvprUi0/VtuGwVLMWkLGGpSOnd9vcOgbIyo9Nbgl8wtK
sa9/cyzH/XeLoNIB9gtLDjaAdwxHbm/6pk6vRgQOQN1pwtM5I811mjqwH84o
ZzXQIz9s/MMGd12XfuaPhFbsk+P2nt3WxrAtQjjymuk0wXoBA7tdoqnMyBSz
sZIzHE76uFVzMRiQcAw7N39zujR6m1e11ZLHbZN/jTPGhi00MAqcHEJaymfQ
lVHkjXM/49h5xhoHDD6NswQ52gmSdfgZcRv5E98nKz0xdPEEvjW96cpXkNt0
2RSMDCuJpZWU8jNmp9oekSLV5r58tuin3cdwnwB5kJjSsNJhQEu2S2l+Hf82
KCWSMvwiWIQGgvAnBtRNjX8Eu9LlMKlWtaE7L2R81KVR9vBqCkypnaz2njY8
A23yqOOswhlPrtp2voOToPaf67fhngB6K5+3QTsjBKlp20EQQG5vzQlvOcJg
r2Ss+IJBTMa5J4KZ4EW42e7zL7yv5JzUYwPkdNaTrOqItVdL6POsoocsrjKV
Y8w/cbhktkzOeZsIN3Nr+306Rm/jYwkP3KG05b+ALjcC9gd1kGcMmVn8OvNI
wA3M64dznCECR4mAJd/aHmREi1P3/yc/1RdN45q3pIb8D1oZ4+705igjQ0XZ
Vn9tn6q33McizErRtFaNubiUD/FVOHdtz79JkM4eRT9abZRO2bjtLh3zi6yT
gSWgMkfnkRm1qbTPuJXBO3Tob7WMr9KdpF79h1K/FIYPT6gj9JZs3H2eJaqe
IGJ+dMp0nXtp9sW/+TSigYsnwmt+2tdzjzVtMR/B2ZhTa1NHML554ZRzKU4o
pJwXQvsFFso6EJkIgWi8A44fI4SECERftr6uWtCP4tqv/3y466LDyAcz4PHe
tw67n5iTeD8HYCFmdMsH1StwrLuc395bswVKhBNlA6Bn+ukIPRITZGWEB2lz
RjIBsaCO6g4/NRd5IAN39CmcR+79pMWofc57OhLEnoEG9ezsJ0vclLmk2Pnv
QsiZ6ygh1EyHASuPw6w0nI16QM0hsY8dVqPd2HRUXSMm9fMgNJYh6YZHI+IQ
FxCLorGeYSsxvpoaI9K0SGN12lMCx5aMRcpp58Bu730EGvcV8LA3VwEkX1gy
41kTMYfGA8DB76C6YVkKsDCOGLxdceV7aHF/7RY+2mcm9PGh81i4XutFiL4a
0JzIZfBAdyXS+AESerqMrZbteZiqxgNgU9Wl6xOeEDqfhdhIYcBnf6hbfEPF
pERVLKLFggIklFQoJzoniyRu5aWvqzN+pJNbL67doVDNeDjjb2dcXQtFOqgK
yLriU8RBZ0UA75ajlxeze1K6oxULV+HcXRxl95wcDz391CniO1VqD1l+V1Pn
tVxCt662wVlVEzwMzUzlgJw0DBHUR5jNWvJVSGaLfi4zwLy2BQs6XiVJ4b1J
MX6F77vc+B9qC1PAPv2/OYkWw54nCGeyZtuGdV+HLh6zvmiEiA4m5tfSm4lM
NR/kHGium1cVEc+7gVtywaon8j74gmGXX+qGOLqrgJPz6henT7wNPUPD9EXY
JuRq7Fw7eFP2jTEh9M2A93uzDGrbWhOcloQRSWCHDy/3JogjUb4oSFe1GOGx
pC5/BJh9AZWMIA0s5q2j0fX5rUTZ5UglllDpgIq4G4fyKqRW1mbsJZ3s4PDy
D2oTi7U5EpD5mODkeXHLV+GyjjXQGgd15bFJ1LOeoxXDE3TH5Z2FCcgfcdpH
XXcydIeKlEm/7TZp/crLoVHfU5W8BWfReTmuCv3APz+cUFwNqRlqMdBndbNx
dKIdP6TSLislkzEWxZaEyVfKUqNh2WAp58dMxjm0Jg6qJNQrwGQjaWaIrWzE
hnNLZpG4XOzYfOsaUjFSU/TQC6Cse3AzAnPOgLTY5PqKpvY01iG+fJ2rOfNn
J+oW9S/KU/B4syJlUrMT42YqHq2DO3E2KI7D6RALv6ixdgH/cwNxMxvRj1dP
z39Ikx80Cdb7+s/O1/2V4NyiROOnzY4XV65XmNnh35MXJoQvTTYXaE6ujYQQ
q5T9F8BF0MgsjGKwVJpBA798Mw/qZw+MvRJ8iyBomZd44fQq8Wdqv1ywZjDu
7TzKIyQJOekqdBgvbm0xtK6Uok/m7cLVXDZOo+jvLGh8Rqn7lnlTxAD2z1E5
HVHtEZfZm9ivhwNY6JFiiK8LC8/QY3tx3/bj+VzdBcTPxXFK+8umaSFze8Hb
7QI16y1bts7/vcQ8xcFEHksQuQgkeP5qOrfA4x37k1d5pdgSs4nGU67XweHX
sUGmRs+661UGe18+OhGeucFhFwONYZyHYRHWAiF7IHBimraEjyY7PEaLu7sw
ArG54cg4WG6DxUYXThPOj+lNruKXWnCEiSvOcERN695ffzSjpm7b/t/RW++X
8f4VDTWHLtOXjwzBVUzj2YVnrcFrxQBRFgwEYAjYwTaJ6BGLC54kzgT9Bym+
zIoBGMdi9xFkJoTB5pg57wiJx/cnM0uMi9M5itta18p4KXgkaj+bcaaT8Doe
48dEXsEc8SxwnEz63DmuPy+h1CZtY+e+WB1qJOwhFCLIe0V3Ga0CWAAroIA0
vYfe3niaSom7Tu3H6O+V7Pl1UCNWAuEeIwyXrKoPiXZC8kWfpO193edA3EEQ
9kT/sPYg8KyFfZz6pwKBvJejlla2vWlTyyzNJqgd8XPSmV4idvc28QY/ZYZf
rxB350oiu3v5T8z2GhpWAuEKkkAtjaJ80rV4qR5MokdhataBhsMGu8uOm80y
zgzqPJhAkQ7F0iYI6g4HEa6qBYlkCiHvXQ4Ls87GYnChVf5UrcBHylftdcTr
gIDchH0aZxW67zbWgcGhg8BAyTWRkjt4l5zzN9j0jMc/kd9c7PnpbgXuN8Vk
g26sYbXlRh/qM1PnHd+sN6173sX+s/pAzaLREuNIGFxWZszg2vXsO3po5XfI
Sx1vvmFZvWmBARZAwzqazQiM91rcf1LoeQf/xAnlQTnHyDbbBgmUcHxIp3sa
8jzyReco5xdvkRkcBUcD9wjnuJctpvYQc6py/O2ZgCR8xjYVPyCf5DMWDKJZ
lT7nVRvYUrYZPYMsH7karGTUqKJ2V7Su/oEayI7JWAPnuLAagsqPdiDiJsvb
U/7/6WK+wHpES2VNUUS+lUVv6ieCG6lvBB2kdno9A3TBQpNUcoUHbPc3Dedl
ltHeyeGqGoAP++MT3sqzmfg05EISLDi2sTW9ugJEV4XD7YV3y3+/K+tlAE4S
q2sdr1eoOeW3wnF6iNDq4qMjkjLuIIIvmiATvRCBZrsOxrwad6njbJODtkkh
LR4pQB9gFdsgIsbI+yeThIV+NtNR1LZkUoV/p47BnnGygjaaaopixFFer6uR
8EQLDCIlXfj2slYQwqRVaZugBbraODj/xQy7g2iEJ+crv16+SGXLdPLlYtZQ
558i5t4kyBCvZnP7WVUf93R8AwMKFrOMd6dU9exdBzHah+iFqYhXhlLlXZYA
//ssEk7331TqYY+WMzntdxoiDArcHG75FgOl6MjItH5vEzRh+k7DD+hVQ9Mr
uGamHPr3srIjqlF9kOXd8N6tXYbmmLdCNHZ4jg02NryCLRuoNItrWu+Nq951
JByhegee3BvPVY78Tx+phwi3O83yFWFAT/eSfrvY2sXX64hom0pSqcumb0d8
kMzxsb53tvkxmxDK1wMCcclxxZLWZ6ia8z7L31zmHbOAyRCBiG1vNzLm2yrY
Qj5TiM2baimFh/MMUipLsQqxttVCSVxt4A+6MZybBm/YNmkui/+KUX50CZsh
zsX7Yh8DOAyDmL4VaTnDzMQC0ynFWeWlOzbaeQbedmS687Dw8A5NyT54ANgZ
exfp5jtMGz1b9pyjJi+5hiHpeYEa5comorH2NbtUZb6jJttEbgnPo34t7n0D
6nc4OYT1OVJgCLc32lfH1Xeom/3x7fBfD8gcD7tSvZundG4mzG38Jz+CxzaS
dNeRxzIxe9RuFoCeLs4qHEgNd7rNvG5XHbaGcqJ33TsIbI+JpapQ/5oSm2Il
KIgdzeO8LR02DAmPisX+luOgS+h8DQxC6imvUixIrUzwQxPbGwzhx31RhIuY
0b8KrNtPTrQZFtbrJWaXij112Be/s014hvxVNa0p25Mi2G9c9Ij8o/jeVQvF
j8Yedgp2izwhLCzv+AFyZd/u1J/XyGvLMSKm+OsftrUapiRG2HHE+OmvH89q
Wv1RmmavxRyhhZH/H0Gy5sfY9kt6qFsxLWYqq4Cz0AAB/h9/kCXtM3kpThC4
V1LLkYQgY1Lfyg4FZzAzF40Pr47a9yeX40Z4RqBWBoEZNoPG3z1Yp4kDZazo
dWiq+KzCUgGHKxb8Xicg+PF7zfSYvGO/eZSHEhDUBEAi1161aj+crE8NgbcU
0ZVNG5428Hajv+abR9uMTBcmLWED8N0BXQqtnqmSSAGvmXUNRy2VIiqf+4Nr
wD2N323Xo0lENPJzTKKJhsKPHUZOnlPp+KSq0a6cAcRSueUAkbGqZu8XT7YS
/1owxsli84bHY/44VVnDfpIVN7dEqRqsIS+1rVxABuGr+gN2Q+M0WCIUtr2M
ezZwO24a6dEW2gWKwSEnLopZmUQufXXRN/+3jUrS+cZYVNHhs37U+QUkY3uD
ZxHNgJWDOCtExS53pEgzwH4rPe1hhmykoaoLMoEelZaZHmAZ4WukVNQdStQs
N/CFqi4HRCG+Gm7+OnnsZLQAbXulEiYPYigsdzdCRAVsGj7omyReok1HeQHC
kMgLdAfQiG5a0E3yILbD1kx1DD36dUK8VCc5pOdu6kudIi6vZcajwV+tanDP
2xxBxzFCcRrDuLbDfeXFL2jFlhII1JpEPUkqGIH7u/jReMFtHhavPszgATpK
On3QM1GLPv0xCnzJav+ZtatxTePbvO03nKm8/TwO1KqPxJhGXyi21bNah85B
iIdBHMWdMGBbuq4jisuXRJ50w+zBbVVgaBL4Mgtz0y4shiCZp4aGiYNeGty2
iVGQCHGjSIpIPIAJR/GlO76VRbCOxypsHnpQKUYZlNtOaCvk5WtRqDnzG+Rd
AMlBW2WWREI8UZl+t+veRUD+gm7BxVa80cn06g9bgj3CX7QwJprdbOyiA78b
vm6XsL7w5uPmDucuu3XHzIWPhIcGK6zI5QHecFgfyUzQDqc6pWgHvWrzEY/z
UUK86oiC3nbzlt/34SM+qafr6LYw4eekSyEdwGgRClI2g3hunophuXMuy1ks
4c4KfAW/AAgzdUAHRlJMAdlkOldaKUBHXf7K6zPuH1c2SZNOOPeR2DUuXITs
R5l/2kziD2KBTNJwEYpCLPJ7UD0cMz/DDW2CXXi6qI398eQfbmEJvSEkUxiX
QxwA8YonlhzXuNQzFAJGnWPMS8/uV2W5Uo7R8gxNvDsT2xVQdgqLfFIlB6VT
pkk4il4V5QWwaCG0UxRKtPubhwuRvvpGiASDbSdp4G2XsFpXMjYtDTCz9FFE
JwNqvQOhIH/Xh1wNRR63ma8lJA0sfCNe/ZgGmkI9fI771ysorldFVcM0+0sM
1Sz4PrEe7OwVJx663++9aj5VJE1KtlsDXlRsIv63O1WKBz6Nam3hOBDd6ySD
DFZwzx0tmO49BAn/LUknVB3BRbWZ9Ase1NKUWiaAcF7AIigUIK30D7mGrm83
CB+EoBQT4OKIhqrKqcxvwpoJ0n0sbzrY7W1kZ7YDF208rxEGo2aiz3vtHZqq
stuYp61M8dYzYPQApY6B/5xJAG5yWC4v73VzaWgN+rvc5rt/oNlNzsqh9wqU
SPGC65DiwFGRisWrqMzeHq9mXCtIxc8N9GdN9T28EFxr+QV8hCRhocpUTdHA
myuvP819CZYevCaiCy2wiZUyxaF5O4CAkcfDLV9KPGM0oLyTdGIeo1BiJpL+
pZWlk420zJfYbCeU3VXyjI9dDXLoCLpq2zo25ix8DOed8LccWbD7hg02opc1
C7vYMTVKwRwvlaNkuWdz6rWypZAEs7JHX9S30n/KHTYdSrIbvEvQZqX2Wion
slwC+j97DLj7AMX/iOc96K5Pr52a+jB2UGjIN+4FiIByUeOdmtrMK/N1iOOC
/E9rBAIaYj7nvnpvL0R6HR/Fou5nbx9w4dk1gFkODorVnE0/4gugrNzvkHAE
dIDBU/Ahh/pMrH+1F4q00vseR3GaD6Rk4yMSjqK7050H0Q0jGX6XszvCacLO
24wg22nn5juHwUtRqpVxfeixssBPaH1aF9UirIG0dQyxJGuqgxuoZA1jXG5A
C6RdYjhIcwPUdFwsWZRJTFlZYIxHs/Q99q7opYGfVqq+8+3PtRc89x8PP0if
pbzy0Fiauzlu8dzlHfJOsKJVwUJAkuLO2x5aIlu8bbBesO03T3laro9KovKZ
qbZo+Ne9EXmpwoERuNqxQVvwSB5TYjy4chN1S81Dmv6g3qHB5Ldzs/EZ6P1s
WkMjlEJvhIQhs5YcKjDMa+AjfllCA03HbWtNsqJ9YUIkLUeYP0Uiy4Rn6BDn
7uRTbQdYRglvqUbx3ohaoRcooRkC7278M6pNPvH5nrFQnatTaGjDRCbg9R6Y
IB5uXF4xWCSoXC6Rlmh6De/BCqn8utWLpR5dgWz1IkOjZR+bx5J6gWpIMbj4
uAjkWd2BKkgvTgncfXNsIpYuT5lHp/tKXAZrGqXuFYk4ZUJNDvbAOj6eZ2De
siLlXmFkCrvra+VfmvmF4Sk++kGdQEr8L/BOb8U17h9zsv+xUi4L9cD+Lxbg
a7WPKCql8VLoukWsjnrWp9+OtzfoxdV4bJ0JbJXGxZZ2jtWjPnun3ma1Onc7
+ZsRHNyzeGH4sJYYVB9sinTyUWSbXsUDlUNgG6WhEXZ5MU62f8e4v44yo2BD
eFk8LWKvDT/0j8Bg67+rNPO7s0F2jLV0MJg7gOG4Cq/S11wEbE3cBN1F+vTa
cFUSPElHmB6IiOoDu3k7XDIEtVPukFa8AoqCIc0IpAQeXgQDuI6SFxrCJzzG
/Ej2wWuuNnvy9GzOLqt3tV/TP2Xml/zx5vPayq0ZFkXNqwktxhWyXIGEhATd
YGd4Dptm8ouPWRX5DHzsVX+ScXsPBi+CMSjreqtUXr3lyOYFoNInJp9Htfk1
VWIO/y/zeNO9JRm06sZbCckdAggsPrGZ+CseDwAOub+eFJiVHDwpUFqhz7Hb
Nd07wd6FFNXaA9D82mVgG1FOb0sEdr7ZMOZr8Uy684JjOuNUg8ak1DJMp+l7
V+Ci2x9snreeDA/m+Bs4dpLeBFi0R77qrdc6C/N7C8FMvz++DYVuGHxN+CjX
0P0kPBhxFhCtovIDQBlGcsRsWYxDYH2EyMT9h/DzY5gOfI4Qga9AC7a45xNs
NbU/1HAj8XQtoMdN8aL9c/oLrnt/1onEom/xW3d3K3oaeon4CoRQ1ljUW47R
J82Z9mauhUHMJblSQYyCUsbrVt1p+AysM12QRHJrvBjfLHBCa+IsHkKfQ6FX
81vGT58V+VimnXLDDTtzGJ46FsSTUeDyfwV99USNekpC07cJrQG+U4CWrLde
ZNgREc0a5yGHHuJ70HQmro5gSeT/w2HTEKAK86K+/ivlx4qPLja/pV1i1k+x
2ndB3Td1I4CdWHN2wDPfUsPHvzS3bFGLGq0W/v8EOFrIK/so65hk6pNobY3G
eSYaBKYpojUSBy973h8pv1KmsrR+JLTWrx5Kw3H69i45g6cgs13G7MPPznIK
UY5YuvKl+wwCX8vtqm2RxOujw2ue6TJjG8u/A5veL/LSbTUZ8SnMtpjzhmXx
0S4pZN2pCoawmdk2U72mKk9iLKA+m9Klc2BJ8QWexalGQwaaCe8Pu6hMUu35
byGOZrYd3I2C+c2BZOoi7q56T1Muvi5mhkNGgjfzTZtZWilXw+Sm00+HSb+S
QqIAFqPxlzzIll9jyTLEIe9WqC1mCs5yyFmeE/tex8mzvECuZHas9cTlqb2R
0vP2DT3j4ATrc6OQNRNlYbjJR1bm6CqD8dzWusvbWXKdjp7mh0m//6bgr78B
Fs1yedF+pe09CCE49C0C3x7iIAjW3AHNzum4ivWkAe4Q8l6qNTE7ERk/Pm2l
nKt2JpboLsnGciCAruuc3K3B5L/viYY5IY3FZDqtfQ3WL4Ks84lOY96bCTfo
Z+Z7T9sNFX0DIHnvDUqNBn5firwQENW/HQx1tbhe6EYCAHqfUAxG14NgpjbU
OcajulieoUm3U95/OYVJ6W8HGBEDtoFj8hjPYCEsVgL6xOyM+3OL2UgzwZXC
z4IIJobuIdoFLdkkxJ3PqOAPR9ZJNZbV+xpenouq2co0PEfYMg+Wawm1ss2p
4cIwiGH347ATAAaOfPFyzqKgdde1A2MpXQTDaYWTpWljIykZiVV2B+VmjIjO
Oy3TxRc9zmc1yLyRtg9hpabZK1F1zytX9SAp8SEo/dtbLk2jKyIJyxMLgQUB
TpVJ46yCxtUy54QK3cc8p75Fim8hvTLGZi3TU2bs8s0UndOJZaCja755XGSd
wfv6qQf8uHmGZs8GHDuWDGlv/XHOX1L968isZh38wL8Mc4xAI0xA6cxqydN8
Modj18pSCb7WLV4NO7RW5O3vmlg79DFWbMzUhONYR3wIlETRv787RJmYh7ss
E9qlqjfgKB+4XCQT1fB+BiEngqYUu/+GSweBqd4obNoasPEsaJgTTAdNwzGr
s1XEdpZD7FAv5+4eJ6NwattTo1rhO4bznDkmq7YUjDP9GyNEH+lzUuy07IzZ
e0bVP1XGpN00qimaJAwTIiiYNSG9HyxiEH1GjmabD9YL3ZQUmtW674d47nNp
quJAUgu+4IsMbN4UK+bvUcv5FSfC6W47Jh2janOtZDNcbQpi103qXRKTI7HS
r6aqvbg4NInH7JRGHeVdM+r7MO2Ej7isij6j66P0IXLcii5+q+Sk8EOizGNH
hVPwMjRQ1qFn3gcuzSu4PTV7tXpgqvJsdK9P3vCd5/koOVoq+g/fKxZS7XOT
GfChWrKgpdpaGA/5oxi3mZS8O0BLuTYmBGzRTZg24dCZARcEsaTU7AzyJQl+
eX9s1rF5KoMS7k0yCMyVk/7LSECSynzrcRciBTVzKWLFZkXWnaWRWajoWh7g
I+xNhg+KLg79oqKPXO9StkfDtUaxuW94n9WHGv5CLH0ISKYOthArIYAZtPqL
1p9NTPBqlYa4iBkenptJqy/UPa0lU3EjrsomeBRhQWoFahY6kLaHaFyMQ1CA
r927HiE1uzVt1RxAfQ+qul+Qvi8TVCf6B90JahdD0IgrT5QPGtVkEtD1i+yL
KiwuL/7sdyceDtMPuwrSmKZxR3BAeeIKQ5YiCYbCJWM74NpNn/xN9AHHyPGA
7UtZm3C3RBXLxnkpqcwfnw2QkFZVusi5fDSTVUZonjpJ3boBGJTTKqSxEapd
xTIVKJzGx3Zi0PIpqUVTNOdAnhjZhdKwIV8g856vJjMRDLQ1+bsjnRC7cvSe
AOTzPMN1bMDPxT4UJuDnsRggoRckccI6LIrMK/cAMiohvnuGT/259mXK2L0H
0/8HqNc4HE0qeig5hwJuHfrJUxFaT2jEtyhvuijnPqvbN+bY56vPiyGCNjja
xaE7/uBnLDUCnwFZYG5THfScXu7GfluWC89fDXigSwULwRzI1ViPr1IEYDXb
DUxEm41tviP56drNvBoFdzcyYNa4fTNw6Ld0NcHtWSlygPQS+0RNcym7eDbB
hYexYXfaB5LmKmQGJTlE0sM1mHgm8UEj0sD8mHmf6m8mqBRCZd4fMRFKkNNb
Gy6QHaKWcyhK0jt6YYBUs+XocEkhq1te+ahe7jn2ccOf+aJpHmtVEoaTVWqn
cUDNIQmmvYXgJViM0nvxFb9e9VvyX1v/iyBnxKd/7ZmFnieZJwYN+QPq5gkU
RT1K1e/ACK1KEy5DROpWdCoMLxDflsMVs/PGsQJ3IfdGZjfMKSVOZ1Ju5fF/
NDD/QdvZHejmfjQbR59qqiPR84TNjDoUjxSEGL6Y1XMYOjlrZUyufkx8HCQh
xdtW2ZE4MFRsQLudoPPfa04lqMf6dg+2sGePWN6eZJSf4eMyDrJLOpHNxD0U
7WiLUSe1FHxMHnvuWXK+krAUqy1ZjlAwdhwGeL8pE8huRExPeV/DPROGIF9A
ZGxxXr11ksw4N8Kzw89FWvR3AeNdIJgmuzKewFQGcJNwEg0caTdsE2FCEUW4
AnkIm1WEFObm6puZdZyP1jCWnr/ZhGKK69szflBw1kYLtXp5f6wi4uOEoOFD
eWER1MssidgzfUp/SFuveUy9KPIuUP/duw2SA6VMrZ83qYQh7r58KJA+wabt
XynYNKvVAvV/nqUu1nZMMNGgm1MsjRDEReN3fUa434LJsqFwc6iFhFAmBb/K
YAmmfCOP3fmKDJ1K5ks0659iNkyhvldy3JsbDnkkfq9QxJSAgTJPicPqDC/F
bp5ew/eZSsT8l88gY4j4oNqPgir5Gl7LRWPYwr3mYOcpG9Ri5feFlmjYsYSO
lCiyvGWCNnsIEzRXzC1CFxknkTRLOK1bLDiA9NDiu4Q42c6N70buLSQ9kB94
OlhcW3wR74H8nGFvnP43XmbMWl2GgHXgJGmJtOm1rAGAqCsYlLieallOGrBY
DpIp9ffkmwmJVVPiLZaHLgwssSCUvn1ve/1hl6ovyE8+AtEETlPxfkVtMIHf
mbt9A2r5JSnMM/+XapF9GFrj9lvSK+nkGXBY3IIvhw28K3SAZ2/pf1YDLGZT
xIBnkpqLFoZetel1ZRAjvqYPfyZ2lHvl9K6afWXUr12y+Vw9Bd0MPR/ejHq5
2o0Y7cJnofwnFim5s7KAmneMOEl2iUW60jY2HnRoiEV/JRP2iCsweIlrfa6R
qLnWQhHO1eKZd+hDyhzQvMSl+5hy/NVyQ4Q/IbwCqoEUdFTnnizfUQjXCmH/
GRBaCI0ybDDaFFtcLD6RK3gxFRg/FbJxx7e53jOMIt6ew3TkxDeL9ZMlT4YQ
wJLE4P2E2nhJ/t7rc2tXid/woF0jaYT4+skDtFh0R1lYuxuIyh/SILfTh/qL
oD4ZHsXP93XRiMwWlvNDC4fcj9sP4eGhbolj1jhPlGkbauc3AB3TnzYyNBN/
qOdKb7Jboms6TzSTYm6svzU97b74pHEo9Ws517k+QfC6SYk+9uuMaFtfK/di
wREaz9aYgN0hdBPo4+cBk3/IqYwDs1qMqn9mn6LZBKuSAuUIZcoL/AeKt0ar
Eta5Hfu/djF43L/6K0TE3AlLm2RqCwTlAEHCKDcHoMg/+StLQReyihv4+6h1
GGMn/iaINlrMB1iz3Z2Pg5/hB7kiZus3ZJMNEkrD7DJeoVHBxyNF3vjdABcK
2SlBC3CCrOmXGiEorohXx8lNkrBfvwRfgDFS6a8xtNdm6/gZhnxbW6MWqj08
hgBxbb718LhSDnaICZUsYLytlPUpbF50IauM/mlDA/WnNSBm7TmqCJZSycvl
tGoiW8ceHJlE7DtwfAe4CKe2D4xWucoj9fE3Me9O8XK+fqqPbZe37Y7Z6h2P
ltdboXsBituaWJ4npJn+vwzwvyN18Q3YkR9Oh21pNia8VN1U8fJsRFnBN+HY
5XhZqn8RTqPShfopLQlgcI7NYDYjYJmt/W0xTWwGzteufndHqfIPNNyfgkK6
IKpEOhHy4QhYONVy9euxo+D7zCezOAkIQLrQvglC1rmbPj9IYU3kCwZqP3Ka
8/qXEHfuzpJji8E5iKjOIGiGpXhMYPVACZ9z18+vtMPEpzKu5Ut7IjYxGp6p
4kzOQ/lHK5ocNLmSU0nYUbHfcyibH9YsaD+iSpf5MhSS5Ihuj+PY//N9Zqae
1/pANuNPJdyZzknbG2fIn5r+Q7VHp7oOCeIQVQxF6Or5VojZOv6qgjorAj8f
dBWAdVqTFuP3HbNxOw+cFYTPrFxqwWtOoFZ0z64lZ4HVQUXVp8A+h6ziHy8W
yKRq8zfjgQ/E3nasfINVeFbdIikBVGAuAYAint9dBqBVvjx8Zmf6vj0kQLJL
tgXkQQQxtjno88INYafF/BkK3eyiAfL3K4w0g0VD2jts8APj8e0k2uueOvFl
7I2S49Fbn5ByeV50k+yxZ15t5vpgPxQydbLXSZQbKfLeQSKy6C2mhyqBNcMK
q7xWm/AksqdynLATi1EVUCzk8e8h0GRRC1x3Sj9ZSe2qnH/31/BbGpO9KyfJ
kGeWtaMCbMwZOdOP0hSxXE+RS/PzpNx0ednNHsNe6uct2ScDivsMFODCkOJ+
IMpxoM2wdhsyNHdU1FcJv2aMIm0O5hlXrfdNz4foqB+bOsK58ckBsqmVPjAz
fWVutgozzO53wxSdhwZdsPFCXm1HG1Eq5zmXxgLOwSzYawjY4S1W5YP0Hci/
QWqH/LDxWzCZXzpsGkdOyD9u6DKBgZxHGlPTun26z963hpQ0cixDJ7l9ziBB
BYjZNVg+Rppqqg+b6U3EfI5CWAID5Va9BDxj5tknwHpo7xWV5/mhuZes+djR
wkJ4aD5LlCfEl1NJiOniJVTJH0JwLwiemH8oZP31IoWCEmNP0BPXmflGWxdb
F1oLsboDDMwRnZwFDtW+B1drN21klW6+oJ8fak3K9Ijsj1lMErtxiKmnLBX1
3tDrkPx9fJuUH6nPIew3trrywK9cc7cl+bGO9stHMsUigf5vhvG5gTwWmAPu
O2ZRe6erZ1Rk7QV+3v+ncc73zxdqy1LTVuo3f3uDdZP8eURJU/JL+FOOj3da
qHHKU7b/rShYYYYEcm0/6wn639zUIrvM+7fDnFAFhcX7SETqaJU5+TIZDRnv
oZdoHA7VFapft7S2rYtuzJ4Ust3AWbpc0KInOxRkA7FiRWgMf7Cl/7iU+b+a
VhDW6YsE5cXoUZ5Gy1naqvS+iBeGZGAs91I5rinJ5g7ZbesoUaqMA59/v/IS
Cw4Fzo7pYRO0o3XCVqOPHfM1BlFE5KO4HX2/K/tJhP0tHN1l9QOWagDt7Ipa
nyLwBbR8YzUmJT0QYcLlNhbgazApiD3lJrzTUzYOODHc39FwG6zp5busMWd5
Kb+28Tc08973Zfoc7rAaPcE7ffeFmMke6ncOPGnk0JIDkBw1pqBWgqD3JER6
WlkDpLQhvosW41bV8UDo8+FDGt3np/G4gu+N8UH81iEyfWkj7wTEhYF+oCXI
m+eLKE4Q9xCKAkEr7XiOeXIUvqiA60W+5ldqFVj7dnDodZny62RiH94Gnziw
3aJZV+IDf/MrOjHJ4uLc8bG7iWXrXiwxAKstvnVoi9Gv8YnmONuk2EhHz2Qu
l0AxsOOdwLZVqUBls5wF9+tmouO3fVX4reQYX1jGLXeHMOH3D3PceF5blbD1
7sXQcoWHMxR3jg/LOFLwUWfISOwZKzIXHGtb0OCacumNTBCxXQ1CfjHDj8g+
q8W6tsowQsFL4BS6QbU7VqEipcFFh0iYpELza+L8cGqRgykXrXVMPC4HFCjo
YZyRFTZqK2qFHdFpmVyH++E1+e5fy0eIqV5fVhDUBtwY7ZewdW3l6Jf3dE7N
l/NvXMtlkfPsjIqX8f/wAM/pKIQ+lIi7pexEFbCMkGeCSvhSRpnQWKXvQVkq
B/j4l2db3xMelxnucNGh9n2Xp4I3Gcbi7IYgL8QDIbQoNMGbEUC7QeTO/wwU
TOx5ycR7RRw0k0B8lntibO77bLo4WTB4yLW8AC73Hv73K8UX+6CdQvV2NCz7
069D6yJPdZpQrusJDZYv2LWjZK+Ai/n4EizWQRfAgCBlxY8jVjrntrJmTm+7
whjmoUvyOAnAg6PkKWdDNorgpsXUV+OKZAN/734iPKP/2wjS+VJ2gYg2uc4o
JQHpbwRN7ugkI2WkddeDuhHxClnL/k12l10iELoJYZbyl+Y7Z/UHPS8McX0d
xgAKbwNHp78peme4avDt1TkeOl4kNu3uN1UIiSXdbtmk9L5b5JLVqk+Vsbgd
z2GPfuJCxt4sN/kJSi+Lgdp48CyFVlugBYAWDLy5hxFAoBRDnA1LcoabumBe
gDvOKD0Ik/FjNDcGxKX483wYD8Xm4ehLRP8hYRoloFRCg9VwlXnEKGdbeaiG
V6Unc4tP8OJnLigBhOf+ENp1vgkim+RHl9wy32PueuwbN4kh40WFXxBw5SpO
OfhOewiX4tt7RebDgPNMbQx2Czy8yDiwrSTkp+ob2aMBd2PtT30URNGSllPO
vcQCml0pyzyVtI5fVi1C0qlM0e3KtSGxL2ujIASY8uE6dG3HmtheNFB5jTy0
W8y/SACzaKHZaRbmsozZn2lScNMSHBy4sDKkTryJJYgi2zKQcfGJ3h+ZaWjY
IeEfKWmZs/2ffnSdIpA524Fv7Tzil35woZCO/wilVismbCsR3WE0r0R8MFAq
ej+UjNG23WVw1wSrNBEu0i+DrSvKfp46+a//dOP6pvgA2gk31g23nZVSVU16
kqKIpFhv2o3Xat3GjdtXHvZbPoCozgt4bz0Vh29fEx4QAeljq62bNTmGKvh8
c3cIV0EB6Rj/M4HOW8bmVsRODLMkautDbqedTmPOODV+UErehcJMzZrqVERt
eVHeIK1h+870kp4u3oYnfPa1x9YKn8TYksfx/DluX9SBWiDgElqMR7euQ67E
QLo1nUDjoqhN5AJIvdHoYk8iIxLoZZ7ZsafE8ruTntq/dOZyhZHHU1DpHdA2
/g2eX7OGJLuDdCDiQiRwFgNRcpRKRvXFisUl/9j6z1zS1+8TSkC2GbUQMdmK
BXcJ3sY1bt4D8sofKT4RKs2nzxkxqhL5y+gVP5im6/5VpMGV4rqV53MHym12
DBrVD2r6YWux5qGPSa6bHOgM2M0rIySJwd9Kj/6oX9RRIz4elgA/5Iho+Dw1
kkEPiVOuUoEe/VpX0KgUqSJW0gWAGhE8e3lQ6ED6NzXjgNMgCA1HMVAeWN6M
rwqsAoVMUMBeTI0CZM8rWwlGXGH78u6dZ8uGkChMJCkobYDjZIxPcqHGa4Rl
9m28kUnkFOrumQbBW5Egi7L6Pm/Ys7goYA80IO9aAWkZMAtG5wxSCfrhHgPL
xDMaWCObg4rfcZJ80SzcXHMNfrwORf5W3oa3eWCHN3g/rXvhO3ve5s7Z/QnP
4hIZaVAKnkhmI8m0PDPZdBIdS8IOvEvdKacO+i7uZppKYozl5TCkhqG/9VAT
DyvWbWwZLKEZpNm/UlpnvnvNT26mMmat9CqtOKNMDKQMy7RX9CpOQDn/iykb
pDeWia4kTObB8/ga9fAx+/jkLb+tTVsnxTmxqe7HbwXTlvr0YX7h/AmcwdAD
PeQS3ntJIUFNsDHR0SBMp48pwilWWKVtVVWa+7M25Ib4cWtgLIhV8z7jQTgy
zrrwVX/ixx83Thj30A36vJy0CktiIOGJqn4jv94Mqj7Rk4rBWGXKaHQkHba0
JRu79ysHI9AaP/N+YYwI/bHKCOGdbhUzsqpuIAcI9gAmQSmd18fO+N+J80s7
9Gs41IdUk3xPhWZS72eDtU1ZUSIr2oEzi5lH/6NoYAUC2NN+1nypgGwgIyV4
blXnu/EdaFbDKbJvYKpT/djt4gxcj60sp0zrbp1YK3dpMWr1Em0i4GshIG97
SSBPL9e9j22lP3uzlHEZtH+koKqzkV/6AvewbGxxSOtKzHcv5sihmO/lEWNg
Jltz1738TgnGBgUyvUOGml/dZtP04d2O0M6ZbrUGO2I6C+JLOkT6QBI9ZQSZ
OUgup8z35WPQAu6wT1MP6IyyHQHcMO12WoKs+siwIeRaheNgE6uJmKsq3+jO
v1sllrlFzG+uMfCTkdwciSRskGYRoazb+XHH2nXjNrz8biR2TbB6fE0R0Eby
KqayEj6cCzoRFboGrVzxkQRrI4wdf5GkmW33MN8guU+y5+rsPcL5hx4zM0/w
tN1XIGTCzR70m5ubFCpCcuxs1wNSy8G3+4kK2EYqTGLVGou+rWFm9eEvYGP/
xRsnHwKf9I73dA55oCL8hxDReVRI2LU4JWUgpJTmKpBqCbouQg1ujsmSBIEZ
iEBiE7iD288gg6k/UW0LlLjv96ONJfJBuYWJdJdfxhoJOF3c0VR2IS/G8DXX
G8SvNf1+qCMlQ2K38INDzE7DwuOy68PpH8OKXdO7z9BJ+sbW7nTMz+xCQSjv
ueIDqjVR504jBCkg1mSi2w2Htcr6+FC5D80eRQmCbL2jIFpBuVNevUMddj8w
DmhKXAf4lW+Fd2pqJXz6gxD7CLtQfLn8jKbMmEkmXzBLDxxiEwvN7ms1VWsX
krrhjnW8nNFdkg40RLh31VmgmYP2HMKdVqEqaduyEMnPGR7+1DnpPnmz28ha
lLiWlAE1Rvb3isWCfWPxqQS7ox4H/Wk0auoppOtcX2LkwroqOcgT/6AmRFG3
+fxrdLw+BLQb5sLiOmTZiCLVxZJ1azS5XVwul2v/SKkeH9J3GhLAojj1bL7u
mbZEYncyQKN9SHvY5r3+ZXe5XWyo3tAr58GbbUEodaQkd6ZClnt0jznMcexK
MBEfkwJS67v8QHMxUiEvP4O0Jimsm9Z8rTCN+yOprhVwa94rUCNlZY0nllj9
bRMZDjMYdajrQcaAxk/sp+E7femrAwY04CX0SLungjTYMljUQZausiL3IuY9
jRoTck8Su1zzClGxzLF7psXDbyPdNvEC1VfReu6BmgbS01nGq/2MH9fvE9iD
7RVZ6S+bN2Gjf8roYuhvoU42/uenqaScPXQRkQdn62MaY/0jCDW1zyDG5axD
ZLIQfEUXSGvKDfG5kRaTSOYUgmnVU12TQAYC37vXcQZvhHQnHMYMX64fjkNc
ao9A7C92xcUZa9PmLhqVXaCcdw5rEcriCtaR3g+XYNGTL2JLksc/jigVz//X
NGsDBMcg0V1n5mWQYE8JkQAX6vcVZ5RvYO2knR+iQvU3UZF2OmFepHuuco1M
n8AZv9vrrrwmdqS7Xg1nt/fD3cbHBA9WBKBhGK5pn+OXZOgULZNJgnhAY6Zh
ECsHcR3r/rrCMAZ5AI5hdaxK1K/Cmtr6h6YfXjNFDL7iPwHRzH7Wk71Cvdss
ipAZYEUbe7EYpLqia45MUTrs27WStKR2/XmcFoIJkYsLibYFG9kNIeqk1Gv1
4n56xaS/03f9amD91UH+kOI6fL6faP503scWPMnNTpkIYUxwOC5D8T9lJ/ig
/qjrFbIBEWFa/TonRJhqDvh53ECG2lN+CzNng1SLm0Px5PGpZLJQH9BaPGjb
YQtIUP95AhCInzooOL+XJWnZuOfdt3ZaG7IQvCl0SztJNfdLOgxjlDMyOuQB
MCOj7AOg/mlm2aFkdT0pxmaz9DkxbYn4svs1O4xtUx+FtyY7rf2NOw8ly9Qu
4nO/qaaOR6uLFHp8XQV/l/3LStBGBQrF60OM8BrQqJp4qw5FKtzNX+JSKkhv
xc3bsndt/fiJsZFxyKgd70A/Gmq6ngz33+bezrrAo+8UAM1EDAapU72KaROc
YtDgk+eOLrWGeWAw8/MMtFhoFfbV4j2+lQpmsUj1b1eYleYUxWV5gEEJDLM2
RJGDbDT1QYMr8b3cVGWWEqkgZXqTNG3rkS+6R9FWbTADjvo5+9j38sG7w32q
dzxev3qQ41geuFwVanRSZLlXZnUY2TKjJF6R1SyfPZIHUuMe+rZkLMV74Wkl
67g2/tm+xUSAgzJr6tyqoe3TS5SeCfhGaqPTXrJgUMV9wsb5yHxgUmdxNjBu
xYYoGCg7Uj8cc0rNCYIdaTjbPHLOCSM2P6HcJc7Mn3yj69/S91nopXRsf08x
lr3FUw+EJlp6sl5t1/HqqH0G5XUJTa1tMNMrS5wNvCEiDsVYgMmSrg3aTZ3j
osXkKeGE46S8+eV0GtOTGgxeOF9BLRLb/TcWhm9EMjaPPqDTjbPQSiMhyG/n
aJbfqu0hpHhxZr/yjISGZlq+yIFMFcx+9LgC/f0qq8X+4AJT4FHAIMMVx22Q
79DrRo9CmCzkyYu0PwYHca982mCCPhhnwlpe6rYKcftdQH+C+DT8j93DJy7j
XT0sR0AcSz/EenXDZ5eMWbEJNKSwPY4/GUl2LXiHCwLAHGDawYi8FgA98ZnG
34cMyW8AEsgk3rsCY4RRR2uoeRaMDp/GcI0dv9LkKJIT6Kx+KJ81ezO8dUOn
0eWt0CUDDjw20+ZwI0KnmgR+gI+0X3NdJ7uZWUk228BOW1d0ltb3FkSwnR2A
PZd5mQRf2xDPjGeX3Skm2AaAGRTR31dg2jai5e6l9WgPnQUA5ZLMLGpai5PE
loYlQZkt+4DhbYQ6xc8Ii/Bq2vWiSfmX5kIr9FF6DCnhP6Vqz1Mu75KVsG+b
OF/HIlypFT1Zek0vnbXF+0vlY4aizhORZjtMa/rt1pLRwFsxotIV16Gcu04F
rhsnC4Mr/YWuuebc5SC6Rmb9A0Nvc+3Vq/dXzycyPsthSK81aaEYfRfrQhTJ
Kq/XAhU9FC7lcfP85JMhJamkF0IZ0z7HvUJPIUIfC5jvJZoP8YpfFtVQ2xlx
U90jEp6n0nIt0CdG3Stfg5gnuMBdYz6SXgcX9BGDc0DSawQZjCl/xnD/w7Dm
iYbiZpfy6W6pM/At6VZ1cSI+ZdOBppnroApGa/CIb+0hC6RE+StSXE35MeHu
M6gmktsKBp7PLKXDEWztcD+b4mFCHt0BHjqJQ9N7M1wilY2hEAxy1vUy8Ssh
oQAxJDvMFIz4F1TNF9TkLRwvzyN0Q+lZEPPNykFGKeZZGFwp/2JBguwROI17
V5/1T2kzkwikTiTGRA4wHAtlLr6nkB4excoWqjcgA6WKJGVQ6FsczmwCUofk
cscLbV2rfB8Rf5jBPOOgRv4/UqHA4tpWCDKKD9aW5FTULa2rAFK2fyR+u4EW
m3i1aXRR2Ff01X2Wff/34zOPVziU9fUYFXt3RqxYV30VtYGYVUvaEdceFL+D
iYsi7DwnTAefkF385sAkxkf4TzRftBvSXCgs/2KuFXtLe/HW53QFo+NJLK+L
lLz3FBk4VNxMofx4Jh+c9r3uADe8hZpSGYmISJh9TqgpbMZJP8JreArrv14u
LDozjOmX/ThYoT7r86IGOreE9bHrg9SInFGyOG/zPTuSDA8KPIRomZKsMAgn
lGECrhcxr1AYGUXFv5eoUtaUM876wEurBqcyxzlZOeNS30xypkgjC2o9E2Gk
qvszIs1cSYKHTr0HyS7AmDA2Psb5qzjb849CpaRyIhBnslxd7RqDQnRBo35H
kTvZ9kHB5yvIlMxZDwPz/Lrhwp8RPoPoil6D9NfEF61k46iMYsk7z4JS6dC4
d/ptGO6eg3pm8pdVWhe+tc0DWVICf4dggx2RY9hYHtI05j4TSxH1hp+If77k
EuS0RQ8r5vmdzfnjruNziv4WLBB/OryoxeIJ2hwfHTxyMhsBHH8kyg4gLPuq
SgojBaqmlXiHOhq5mFAWEpUa7mnTtO0J25BoyBezyGqTvyGyDLFAjipIv6hW
Yp1GkaioGvZEKr7vZMFld5Ukg3i3DrGyCcmYUA50JmDh5Of3TVytNCq8rnQ9
souEK1g1T28fPYQXgiiXQCHaDj3B5nKdtFLmJhqT/kR3rP95Cq0vZrLJ4iYl
lb+1fGKcw2HBq/+Erl2B6jv7nTy/2ncFt58RsZNTL4/u38XfWPPww9957o2g
1Nn6oeiEFxbJ2yPuViqd3G5ys9TbDKFshPSEzvtvAMivgvpe/nnU/sfsfFCy
fbsg6Hts0AEvjlfo9vFkh9XIEBHndmWXw99q/qPWz1vGPXQX8t/d7Nq3dbYC
9FN8K7ZD2Le7fZybPNZMomDUJ8iJPPIgDzWUEktIvPi4okY8e/lB5nTjzK26
Ps9RFsmZqXlPNxGVQphNXS/5XsgJoZFcU93g7gXXrLvyhCVtSxd2kqt33VDV
AXHl8FBUTSKiidz8NT6qVPsNAHp0PU7hIVRKb2bQorPH1tCpnNPjWlwwRjAL
HqQQ+P9XFqaMO9WvLxefXPL324/I+yxUUmQLU/Vsb6i9GN+pdBcJW3/QrkPR
+j3yuLq9FOHroUT4xrCyAXJJFZPXc3sKSdksg8r9hqJi8eY31okGl617j3Fj
l/Xx99fJ1fZU/brmtYgQjmnVHin7wyNa6dGpwAJ3Tdg44chkpZETPMLAFt+2
ypj+7aIKORPMHb55R1iDrv/R8q1xIiPxos0bE9CdEPRA42DxrQEY3lBJvd31
T0keuIsWq3q787pfCuKYJjLbOA+U8io2GAlfSFtT7LaQ1rRaA7q6okG3V8aW
en/LhTma5imhntkVW1D0o65/dzwM5KO71YiM4DW3ztbxKIKcRcFpQ2qLjLGj
v0ibojBLEeAzTy1neMwZosCzbIupBMKR7ey/WFEH3vdqdV4fHlyZ/qWqrbKl
yn3NPg2zGRyJKOw7fl0DNa0tH+ek45tRCxgU+kB5Vr86gToM8+R5SNtxh07Q
2I3t1lKj0EXUXbV5UxVLhRTc7SD3zbHJs3SfnG1NV7bPQ743J8KdzdwQVN+z
5n/4JkzVwy3QWOTcagHTnPJ0XkOu+M1F1Y9TCzOzhjPM9jfY69sAAnkqM6eQ
nX/tGA/81h2Bur4D4xTuSofrcpuZyY2xdwEM5FwcczwAKvoXn91izu+5fyEv
bP849GO9uaI6GEK1YDw1rM+586/tJ092KxVJcHxjkkmARRkgMCQBpCpLOgxU
4MMjWVOiIEcoGzMt2djqdNSTexrEjHg93r5oadTi+wIKxyvVy/42dvOOinZU
mfOmVSKt9m0NsN9E64N1NTNMgnZLEMmNMkCANbMYX1dKNinleEwN8u5xq2iB
rQg3Q4B+qJe9jXqCeEvbuxNTilQzrOqpUqp8Q1nBS8m83O/BtKd5ulgSdyJ8
i+02lwgkxIa+nXfoUjNsvmRGx39XHfUqb1+HlMV15ZbsqiMPlezpGEPFKali
EesLx2PQDMQ4XuX0EHCtDEnt9OsyDThR/xt8+dvcK+M3B6qSux/y6ti8zS8P
8twBZsnL9GQY0SWrinPSoF2p/36TCzHniv8NwaPFPvHGkOgpR0HVV+TupuhR
UBBwailFjEky+2kfFJlgyi5bkSubVPv40A7lwlzj+DFkxrf7qaCBeOW92O0d
jM1Pk3m7Ninvxq3z84U3r/S7OF84XCO+Rg5jiZE7i+KLx8B1eJ6c9urgq6+X
CFvw4GO8jtemXufgxT0E/N7uc1LbnMVqAQGaNar2BYfaM1tCYzR4EGNCfmTW
NfXh+pJfu45CXZpJ34KxhPhBy2/V21Mw9ca2tleR4HUYPph2Yrrg4G+0T8q6
ljJAJNPBzFgPu79hEAeAYGnl4n+6cZalFRo1fFBzX9O0fH/uM5HwrAsrHqBJ
UqLYAJrIFVAk0G7pX+egZRgB60iyltnzPYwGVkNSCHWYhyOHNpp/2chvKFRZ
g8D43cqRnnD3Mh6HSHTXrHlZZkbyZvJ9o+6FYUd/E5QuQEpH7kAD8c5qSXlp
wwohwNsk9W2aOwE3OoqHiiOz6tN4kZEF96PHIL4SGlxAhjjDELriEwt1oNMh
bve50vDKZS0k+SgHciUovYj3MLZcy0Zc/kYbTG5FB+3SL6qbcFAsFhABCLH9
V2Fx73GsQ1jLJzkD8Z3KcMoMxpuPS+F2M3/1gGPULvJqa8JDAaVTyEBLW1bn
vwsQ+DlL9Iun6ECY27xO3+DxNwLkgb4EWcd7WcQk8ipdDbF3LmgO9PeAJSci
hbZ4zwYFEgasCHM+gVOE2MARd5IQQO2zqA05Xe786qxA09GDy9bZ649hEYGX
gLn1/qJYGxqzfAsAVNOdpnzBHOeaBIwIUO1/BQEPgOL0eNkAUx16TsULAiMy
yl9z5KTc1eUfkF+ykru1Yb+KPmkXnRoReTmsCgVxIK0nngW/Cjp/W+oju8A4
sPLmWTVH1MRkNa7R/k1NTItLxQ7Gm8x/MPEOEvmlqJed+zyIXkvLrqejMw2Y
UuzfY1iYSZeMovk1Kz/fAu5oFo7ICuAVuJtJwllO5IJ5Ip8z6gDTz00LO8IQ
9zFayL9mtN/YLltLm575/Egk0sGeu4a+L9ESNkN525YlPv0WzUW/JawEgilZ
hVmeNk/FRNmz7d15WYnIufUPHF7jn2XvfWZALDR6OHjIgLV5WFlOrX+NLIMl
3Cbetr5cn4Ym96mZtKk5wChfL6dJK1twxa11KeVRDKpejVBm7Yrait3ZOW1K
jpYVTfi6uFY0pUmcctRKUjyhNWEdTKhpHR/+c6DJj0//QF0WXtqvYRJYfAw6
0lnQi65XCIH60W3ZNj+djYIyR8CkhKPG47e5tZxtZs9Txwgn70UA409i7DC1
5bYKAT5vOz0QQiDsSdHGaVbHCsUV+KF2yK8oqFKBAURUaysO985spuc/W9AN
LdlDIfneIDj6zMCYe85jP/VoSHFwYQ5h40aGDJOt7nxF2ER9yhu84H9xrxN8
Q+Me+7vrA5p4Wngzul6Pwb01zDuZFaTa2WzPrl1DNnwO6zkP5oKmjbAyfjeR
FYXU6ijntH1sDpYpA16peVv36pt/p13yUt8oyUiiHqOzmikba0mXXRSvuacs
fJ8dZIM0zAPV2TBZiQor9RBbGkGhhdxULUbt7Ohggc7JlAxpURfpUhJnmx2I
92gwY+h4bWZRAFnY8yKKp0jTcHgg4/YKQkh611jT9Jvm0zLW0cacDpYh4Yb3
Zy/FFl2h9FSC/XFpTVAg9p9I5eCucfGpjxthWxLmqIKhSpR4aU00so5XuhFr
yxDhPh6c1aW2pocCmyNHkIH6nc5eqE/0qWfACb4vbIymX0f1sPv1q/Otk6b5
6CbTHCe+PIkLSJqS7soDB8BmRThF1NvriZVrTjQqQAp9PsvIJDVDAgFJVJ9Q
aRcljGtq1uuqzdoJj1tkUTiR1H8HsNIEWpRhjn6Fik+pNxl1auMXEFn8QCTr
M1vwZAtsdTnQrN24QYsdL1LfTjzFXu/RPK0plcSr8E0jj3Uouhmbp0bCTO6m
X3MnY1NRQsEtTwFaxwOBmgBblQUssNPGa30aWngOP8T3TU0gIbzfB/6up1YY
ROGTPlV0EgvXdBpyQycN/aVlA2YSY/e41mgJGvHU8YjmqNA4ekOAmGpDuBTx
nSr0dx8+hsZQ2PTLJQfoNyTVJ2YJ76n+xl+b5oDoP6P0R4Dy7WJ5NCurZ7TO
GToaG+icZ5Jwlseoo6LJO3/V6OTcUI+NBExRhwo+jITKJwVD0dAA8D7Vh6Kr
bPvVFUkWm3IbHg4Y6F3ksjRefFPC/mG7jHlFouqUN+VyzQrdZum1ohnkbZBA
HlASWe5RmqhFoa6jdIX5Az5AjeBNLLSriY+cjB8Fpnrl5aBa0BPFmM3FhTr4
Rtr9HV8O547Pv8MWcrlIe086yIFPT8pVhZgedEqUr4NLrYaYSSgT/n5hb//P
WMkd95t+rv5A0DsiYSNteb0abVMvzLzxUiNtspXN2WXx9Zwn4WC0fPsPITK9
/yM0KtCioDiA2NgQVzuc2UcJGIHyFFCbccJZ8b9zRjI6noCiqfjJca9GcwoF
5Ey+kEav9ZsxmMcg+bIGkrqOB1RAkVE+gVtZ5ZWNTya8f0+eBke2W8Wc507z
hT19GV22h3TnHHx7fjzM7sJMP42E19lZ34FGCl0LHNtaZfLtSPyAIfckwmB5
/i19mdN1Y8C0YSNCcojUbP1zi8ZD6nGW1JO3cthU1f/+/MnpkPh3pyja0SQH
woGQYuQ7H4ZumDLI0qEofB4XAC2Jy5C4qKOQ5ZMRElO3oe+WBCC+MWfW9AGC
fMjcrNaWBPgrQkRuo+YeNCNzFVtEt9OW0CA20FXLVYuFYGO8s4+/H54l0xT7
2Oon1QG38L+RTNuDa8Z9K/D5kkDhB9s90UJXP+Oa2ZwPAc94BuxycxHDUQmT
0uOOKJGMmDp7pYp+8TZqByJEANvwaDG/UtgA8dxECQQP9RhSnaEjAj+/tlVN
BpPrWaCCVWIzVouM0LKhO78U6cE+R+R/rTy4xQeYeegLG9narrgrU40VJifC
VPb86B5Z6CjZYA5sYPecc2PG67ObWwW1dt4AjVNE3UREvfqfL/M0iTnzz+Aa
FQXU+KN2e/I3NE87/e1UVgN4exy2uViXLTfzGNJkU8D9NGnH4zoPZdADutQ3
MG/9XfU05dXHNi/VNa24vz4jnToCFlOkubI28xlLzRXwa2kgSNZm3B69/UCw
6c74aCDrvre2enTvfcw+T2n+zlel6wtUAKV/X7KRjGm3S908xbJVa1L0E0LK
SEtuMh2fE101TYw1zuinf4tZULWKwiaeEqxFqUmxU2ASYPArlaisctO20Ms8
K2nVw8AiwQGFT2n/ovHxTExJCNJpimIcip83oNTVjZ6OkQan5FgD9H1ZFNUS
2B1RYA5oRkpBeppuG2omNoptx7cJ7IjZoYZ6zEXt5snvRWcvRYx571k9b0eO
nLPdu+UOGVYFPchi6xLBvt3xA1wkHENaeeptd25te4hXOpji3TEvNDe8hU4J
s1xFBJw/0RScbBUakMGYxWATDMeNBDwITqftgGecPgMvoRoB6OgShbQYsifB
XAEdvhc9c3xNQCfvM8jYpySu3n2zeGS+Rtbcv/KCDWcrR2MjLF6zS0qlpI++
aK0Qlmpft8voZfBBRHa9U588W+Up5MO3mPsfFkukpyZbqFDG47Je5grRXGeW
XLah3ictL1vQ7ZYanvHTkhZ9gWrOm4+vV5TwRiPrPjE6jUVhzUFOvZM+cSax
QaIxdOjAPkDZ5pBYiA1gnta0js4NcjGU5LtRL9SEisnxlbS4ul9eccdLj6eS
IUKeg65DXIdBN9vqGLPzpFkVvc3xGtN3CzUuOYjo1r4mHqT4hqm+JN/Pzy0w
UdH1h2cqaxCMDYSmesaDS29UjAQbBI5TWFQEcIdTD1MW8D/cR5fsAlnm1jKq
yxnBEW//U3OLVdQEYoumoH3BOXoBaf9H7Lrkcf4P+hqqSXoCyLu+yJLrS4WF
3aoQwEMca3IZnOdN5MO71KncdH22UbYXCdLsVYmOJ5XWTvGiSJj+PH24fAy+
k3zL7ynxFDnbkD74c8yDDaUiaa+gN7VIBqVR4WKZ3Juf3yUMaG5oLN0NPH7Y
/PFfcUTpRIwG/aPcJPQiQKZjsoKUhjZ3snJatQzTmG9QbJYE7oVTwbIpyeQt
hckGmHF603VHXP0dRG0sb3vIIXAG1r5+7q0JOhb8jqCRmz0Km5NW19Ru2p1A
ndGU1hdOomg36DeDV3h880Tf52UFTnNbgsA38kGODJFIJEXhQ6nHLWRv+yNA
+5XPd19vw9859xZz/vCha7jJaVj1Dmpw6q8FGAMld+b2dfGMs3NDvooaBiXM
OWRFaKmZ0/DfnCY3glNAAThRODgMcgWQYBSmjKMwP/h7clv7MjzPjbV7/v3I
N/N6REJfaw7xYlSwWayZuF2SFsvUlCxBxmF4zlCPfKQgjPAsauovq8/p9Fl7
943knVRNV5p5vP5rApP21diBUgZWNZjHa4QLVJdfjhnB8OVNtuzNBuRFma+m
AZk5deD8DnaRMCoZz4ATMg0eXY+sduQtSsJ4uKvEmNuCe7lunTZO3SH/7zxr
YBfVlP/stziHLUTshZvkVSbyV/cL6tqT91zVnTfvx86duSwwzwDdjbrnoQ3Q
RxvZOL+jGgdAZZvJkjHYLmxZPBEfD+xkR31pT89jvGJv6hFvkKpcsImocSnX
8UIHYJyZhNsxqRDJeWx+S9Lz4QI/oSF0l5VXEc/w2GdcqGqYLbR/tAKSkg9g
N6ghUkG8jTXUhOO8qPFBQ6cYm9y2H2rQXGS+NW3/lAhZQ461n1AkcfOviOLl
iA3j1EI43ScnB14IDCUG5u+Z9L1HC5d16iNQGmZIx22G2K70/3nh6PF2JpfX
uZCwJ19NZP6UjT5UvWAG+93j16CJWpEeZA6QSYH5aWr6aiB6ZkMefmYMvrrD
ANSlZIAIoMQTrN0We0eMFjcKn8pqqOUadsy1/VZdmlvkqeDGuPe86idyEnbI
PouMB+LdE25DF+09Q1YWBGfu4/qKHuiYPskIh05WcfMP1uup0sM0ZodzPA93
TmKmevzj6hO2U+OAi3yUuLzBAOG+WIEhaZywxGehSycsSDRjQzHcfNKC5+6p
ZON2hooJil4/mn6Qh7FD65mI/M93Z88me7hhVsZP/HC90b+xcKv9NPdRBAlf
ALaB4rCs9ekhjxmIzZl5pAJjON2z4nJqNG0yfOLRLsaOMGawTTRomLWzm5Mr
AgoUFdjDLGQ5Hh3i+ok8o/zd/qptPo+sltkSnMIpbKA4ZfllGeNEttonaEIt
FBKqzqv02JIGiCROG1fVKfc9JPpIQl+RJfYqz3MFkLmrvdWhpVX3BLsYnWPs
JsTXrCaKhVcrbmU6mmktQjFz8MT6IogVFAFH5D4nOy2CkfhLb5ROn2nTW0UX
3iPJxoy0Xwde3kNNa8EGVLMNz/N995WNyPeGWdEeFnKh+dmUgXgs7EZ9CxFU
TSoXCJVKd+3QCe0HZvkL7/iMhyEqUu/Zk9P7A8CbunyNOVkO4Dpz/Qd0l9xQ
ymTWrZr4sgmRsECN4G/f5PMCchyOjdMtEc0PQKpmqNnFvirU/jDq88k79ljp
gkX7HerapXsUufoJaPqUH4VkNUiF/ZI/TO30GRnwJ0rnzyVi8SrXoISOZdjC
p+ElDNn8JLJkCVSGUjG9ID2WB1Cg/v56DsMSV1a/S3dxb49nkw9LBStJ2ocr
3RefAxZLq95K25GKgL7Ue+WG+GHR4JQcBkxImtpEg3q9O70AeaGozzd0c4yI
SqZDRSgewGJhhME/hEr+mZe1NsAx6xn7A/E6gpDJ65HS9EI1RqZnnacEMeXT
MVJJg4qyYD+VGUllyJtycTpps7T0S/mzvOdQ36HfJClx8VIZUL/Mk7E3Hrb+
97GfoHwcYnc5dsRElD7jMOXkkhz9WjASq28qVBDGoTvlI2H2qzui1qQFJX68
q/1SsaOQ2fLckcA0UhClWbHEQERBtTSik/2dhdypjhAWvpLXa3tSX7Tyh5QP
WqEDdqa55aivfxKFSj1McE68vbblb15eMNIjd+2OWkWzE6Atg27Rtug3uN6G
WeEarR4G0HGt3U2c10GiVZrin6pk6RPzk8RXUz6poHA7pnCRniLDbYUyA39/
kwxPEWM4CGJyO/TXTnzyYA2/Z8WMB69DZCs54JXzVfjYKndtU0lnKlOEW6Qz
k8OGn8qiCbox2NDCsQ3i8MNhURAwcVRxj1UqI2GHmmspCWhpOjbnHHET7+bl
N8kxRU+jdynas984gVNM+fhuSnBaKpOxZv1ye6duXuEr9ogcfN5Pxgt77Tqs
OicVvpiLNVn2PpxyPZ8UrKRXPiJE9bLwmEquzzkDhnoql2K7EWwaKmZg4w2i
YOY2AKyjMcxf6faqiN80ojeArU4Zu+ia3Dg2YXv2sXRspqf1ClVaHuOzkSD1
iKKFTuNsrLe+9VHlRtE3pprrytzTqjkh/OrmHxt9Tki/qDfM4o+rh1ujOdAb
rSi6gpSc9dPSkdwQCn1lmqRF99+j3siW/XMtPxjJVE5r7zpk1UNb6arJnye8
dd5xcl+IPAFPgvEnKgHe6QLed9L2zYDAi726dILG4jfRp49geJBPZQ7QTNW4
F0Xrj8VexbFwSIrth6TqfGw7kKtVbYZ/Rrywwql4ZEsKxqeou8JO6CWNDQhm
P7wCxcJqb/vbUjU+k8T2QeDgtutJg1sE9HQOajYF/gFN5+MJoNrZKUuQ+4LZ
hDWpDPavwX0vABBNmnFGimn8bA9aPOmdkjN+xG9r64QaakTrGhJCAA7sQ1an
gBASKzEKc7lK+o9GtYltzMfk8WonnBiQu9Hbef0vWLHgJ2VVHmdZWD6NkW7d
agr7ea6VqzYNZ9jvN063A/Mfq95uESoL8xpokq9WIGlvEutUpD2xx2SYxmBn
diSQLXG0neqW8E5PZW6wsoemXFOq+WzkSK5/aSn4/ey8thB+gSqYglY6p93v
F+PtpKO+0lYtif1TdYlnguAtykjbGHz1xq4lJvUZS6b3ilO5fNsbyuYZPdtL
RxsSs6bmqnXV+LvKX/aUQDhKUgK65/o97dbBmlQyZqyZaPU00umSIw5BXN5H
mhrPUjmZFpJSWXn9pHhwZvEd6t0LOwyxpo4EH7BcNTsd6LGbxgGnfF+qsvJq
O4+jzDQtDA4bPMIJcCZG7zfWXXkTj3zZj4UtBclh4Fyb1VTqZM+jouRGwaCE
/mwm5TX1Q59OFm1BC75IOz6ubfhmzMIv5YHtrgHgJTADfukmhL+rvt9j40KY
AtGxcyoqNZ1MFWDETlglIRIZ21Zw7Ih7ynYFu7SLtj6tHJreNyIr/EWvdWU3
Umwxj6UMvhYCswpLKdvZuzzfMWesk6u0DMOb6zdjJFpJGrz3qvmWUcgb+Pa/
0OWovI1RIch6zF0MTTnwksNWS/5hLUEYmWiJsU9IPoMogACKgwSCLWCxOGLN
ahUpRVIHOaHTIpmsUxGgsu1mSeKb4knYc9grwKz6OFjtmRFqHUvIbj9sWT5R
sj9jGi13DiuQ4s67N7AMwV/wsQ9B3SNZnbLPdC4IqE4/eHaoUonMsFmuHRaQ
HF+hKZ66zOoL+oztuCopkXybsWNm5CZd0eP3viZqJwLfew/dYeRJ4Vb0/cC5
auE0ZVdbzlJNVPdsZImayTAqHaYTOPRmCReX3bdOJTdtisW7CbPeUG2kalPN
USZJ1+3rHGMfXSawwNLXojyylyBIzQnu5XEsJ6MUwMVn2ChKWMpGtcfyVpRe
BHtbUQC1R5+qrsI382l56/pGUO3pYzsVRAT3H0F2PxzPureJy8UNMWC5LW6F
/MC1YgvThu6ukx+m01z1v5nPxJJpIAp4vu+0/dlX9M1sb8dE4SPSlP0NLaPU
uz/zWhtdfwAXyT2XjEel7CDwXitrYjoZn83Q8nYesgAzMcgCQUJK/NU6RNcO
fQf8YnMhnpB91gA2E/5sOqfGybMMoEfLC0MB87i3qxHE/Wgclefgrgwv3+2T
nMdh9I3EKIRSOrHsIe8ISEYZj2dHhY/Twtrt2W+1HrjusJDhEDoxu9D1gbje
jtWdxEBL0Aq1/UkKoNcDDKDXBgAzqW4E2ZyYPh7J2kbqF8wVbOEQPp4z114K
JBbxT+HAoxtXCO2G26zgKURvI+p0VgRAFoLK1voEyfdbHHBUHgcwXw88TRUg
icaxEVYs7AkGqMYvMYK80ny5/1wuO+L7cLbCxLCCTnSjTtGTBMLPNyilOMT/
ZDIyUIXwIsmDcrzUzST/nzaHONmGSmObaO4KzqtDifVL43sYUUTKpREQ4Okn
DXKlRG3a8cRpiBUouLHBuiaoeydvCg6s1EwgDwy3xPEmAyxToKhJI7XG/msU
knhn4YPzNi34vk5uO4Wr0o7ikRQe5XT1R2DZEJvCCqiGZxv2ASE/R2oin95W
ARK29ve2JYJvougKzhOKfQR9OeLmgUDAhwvzTwI6Z8X9wXv0DjbIiwSKcw9U
hHnGuW6i0DeGjx1nMPVb6unIl+WgVCI8PNMU2ngZV6q0Uj+qnoiwTPoW26s1
/0Yf78WHLyVRsgedypcC67hBr8+pPmQRrj0qBHVQeJCSzEYOcZ6T7SiuOkJX
xjtj4lUmfTcWiuMUIKGD3K3ISU5cMbvOiChRqUetxJcvhPFiClAZibnCsMdJ
y7VBU/ftlNb3pJhJ0JsumuDuHSNQ2RYlAzmnjyqpg8x0Ik50u/eK6oJaJcw8
CnfQWz8Gow6fl4WWveW1PQ2fu2dnMpaGae07jP/FDEbhHI5fw2qH18V+tpW6
OhHR9TCjVi+bUfTj8bnB3OnrfGeaU3FNrTXGv1xS4Gwkp80yPgwOVFXnd2VF
VP5lXaUj19p6dYgaoqO7wXqGrRZhvCR81XrfgtsB/6KslF6BoJaDx5fU1X3/
R9gWgnHa3V+414gxxzG4e8O9wSLd1LI1cJ8l49QPPBtvZkNV3GIGK5UW0dzW
3Q4JvnjXEYIz+82a1cnMdU/HLOAOkLllR7PrMZhqmbVbW0fVjVx3km2T+/mq
qne6JwSx4t69sfiQXMahkwFjKxvjgvVUG8aa0RZpoj1DGWnHqFGNrYB7PubV
OXAR9FgF1qSuB6s0jpjAU1WN7hMDTaTloKlVLfJao0njAYgc+/ectYGqDi4T
r573BpE3qDXzaeeDMK1ps4dNIdQehW64OQGsPRpOLOIKcxjB4Lr9XfEEhfRd
Hf38d/Sw3EvvlB7D/t+zfkdmS/3lxWAj7vI3n3u9FlEQSagQa1yd/YCzq3cK
SAozfeGmtXPtGC4WQyY6Bews+3bi9AA77byGPDx4RBeNkqwwfpCaQd7TODrZ
FY9WOgTPvAetwWhocRw87AEMJEGMnJisqSzF/3Hjkh1Xn+W53y2rWwhQ2vb4
f+rjbrk7BduzyZZr49Cnrabwcui8jzGsC7qZRYXyYWv6GeITMTol+iEa3dJX
Z7Qfwp0cOtyvOQsk5ttKbtstVdC/sjWMK/oTzDw1eFZSf0tizX8Pyireb4+0
/7WR/UDs2xHWvGBsp2oFNXI1FjwZWTVh5pOZ80YGeeRXdO/duojGwAq9Wyw0
0KFvkRao35HBVAzqUOMqOjxvfsrua5gbxbwcf7ADTeiZ1iv+mjcCfqy4bkCE
SVwBwUIUqpt08lA3Ire6XPAauxOzecccWF/Agirg7ewZc+UqKJj7Stne7zLZ
2ZUzzMZD4s+U+AhMXCxzcTroJze3ivKbWH6pnxLZdtjw5Aap7wYZ6SJePPRD
qH+9pvUAOiEye2JmwlwsPTHaEWDwo7NOrEpmDz1v+VUrifvsS4JFJxLWZQM5
mhQYrtcdwCiWr9TyoK3ETAigx/UBtZ/mREyVYWOQVFTZeqAHG/XRw/uVlmBt
U7J5RgN7GzMIvO7MPyGlvKUMEHS6oDQZYQLfOpkOOUl79eYmUZ9wVfHR9Ktk
x0coFjSiIwX8vel1gHq7DbspuUwSwg0jyplvQIit0OeXvHWMlpJ4O4zrw1sO
HPr/g6SjdzmHpYSe9xz19uHVYCU7WsT5FCIPQ+YdOISPo3/nAR7S4IEz+hRp
pjo7RbC4SDwWeqkD5LwXdfVQzAi9htaqBqXdmhCax/1JnScaSjyI8XN/k4oU
vyzOgcj0mY+s46/NUep/YPbGjuQR2n3tUhJWWVIKNePMwX1Vj71l++Wx3Z9h
XtWRsZJ0z3CdY9ps9k1tWCMc5mM/7FYWDYGixt5P0HrP+LjnEAv/Z9l6jFZy
Wd9fcd+bKVt51vU5VeGHdvUhhGenHsiiA9knTEZPDDwV8QDlSmgG4RUAocOB
SwxP1rojXs6khrpfulu0q9VyAzFo+pBFYYLJdVz9mrH/1PoIaixKZF5PBGc1
M38bDotZB5T3oXlOkrCSzhjdzNEVKRFGhPc2TxPhzcBe9M1ZB8q/E/br8dlc
IyToB/OwQ4UMCAfsIfdDNzE06SgJfF+HqPCT5J+GW9ULkbbnFmeiF9lL6Wve
2HpV5ETaOpxxEozvxGQcrbfDAaQp5JEwREEooftBytGpwx3FRznmGC1FMUC0
6rxvufjyt9e/L8ut/bsub7uaT5ddkjedDC0NKg03oODFM0/rdmsBV8+2Zts0
DdSus+TF7feI7fLprRVpCYa9QSi2Umdl2dJeckcje/7e3c+buF220Bfiz8zX
rq1eP6CEFkEJO9hoBFjY0FkPTNm/w4TeLQ5UbSfoRte12XSzgGfevwTRO8Q0
e9B9gu8IZjNatFENsEwlOWhalgVfMrEmIURsz4W8s2aK4thcAiUbbl8TNkxO
VHbfDS2Xm9IAwJ/Sxij+EksaL6SC4H6Jk4SxR/20g2cwIowsStdHrboA181b
11YRDjJAWT5b1PmeKxhALsl8Ky0EYzJzSIl1zw40Mj52q9GRgrmMUWAUNfY9
hi46DABq5lIUiFsPbjsgq4XocdZgT3Q7xQgG9zAdIx6Q83erjcGb0g9Th+Vh
M8RLZ7qpvcAy7Xh6dGL1E+99QjlW6vlXZaYMlXTIYLWQwcqWfvvUjRuF3Qc/
pt01vsR+NOJlU9qEbDy2btm36+eEtTRpWBbEWzNZqT1S5cRr2gKbehDX0HzW
7sKnx/u2jpWI+EJQB9MtA5ZfWDZOOWziivmkqAwGBumq10H12vc0ZFuSZz/7
l/XoXS+aEK+9R9Gw3B3PTtKQJtIpZryRiyPWl3FS0/nISLD2tjZoQ/dprSV9
VKumZIiyK73oicVjyfYZTmbVxZTyu1Ue7Oc0Y1PbRx9gfYlJ8eEHjkypqlEY
qjtJRVZP1VVfnvKgO6ozRmbwcZW99P+JL2fl6W7ZQCW6Gp1LD13UnCXXMJvE
RH6jj8xUHxgFF5b/EWMNRPXmwq8GR1MOfYWMdbEfk0wucVARyG/qJM+gTMWz
u2U+KKmNzeaQCj9yTJ0bh7H7Iw7Oxil8BeBlqWcNnNeTBM8mVTEAG6t7ytnq
ZBDeg/49oXH4OFaPfvY+h1Sf0p37x2P4YJpo1ifLug+VGvfjEm3+PlRe8QcH
J5VFrU6whYf0N1fQZ+iChk3gBN5+/VBuNbaAGTcwHY318h4EAwP6x8hfBCGl
ip+SPxnFvH+lBRmtXOf9ISdGbVOvV6ciSUasyV2Eal3x1MhpiWgBqwLLtRAb
FJTGVx/Urrr1jzIR6a/yEDEFwfXpTS+6CaSe3rJAvTj18RRwxN/ypj7hUoL3
wrFIGXkxmpAwZwiZxmDszeYZjFqq3XbU4CABSip9/5vnbk+E+U0KJprPE0Zc
wbUaIkY5JNOCZ3iH/QVEctlbOiypq1j6099RDoW5xSfyVVXQCzN8bygqNKrB
/2Db6PiEtjsbjNbbX4ntTqmY64NwmW7wp+ByQMeyVbmCW2K1bUZxt3VHUc1q
shBoL4RQ8xWt/U9hzgAnlG28VcC9PY/kYKfq+j6QP4R14SIYbISDE8jXOHmB
SPR3t0dd+NwalOm4blkA4kqJmGY6chyEb5oxKWe1hCc5IICw2Ug84h7iYEbh
KXaW+nhoTDU3zSgf6kP6BPB8ckeUx5N1rYwHcx3pPgJmhDlc0dIiuWjB1H8l
AJb43o/dHIpSUO2QCvkSkeI1AwS9tyQgu3rFSi/aS2B4w/Eqfk5Ryd3O1HId
s1AUwZWxDAyUoEwQybCrhDpeQTaGrWcWfa0zbicjF/2gAMKZpQPKS2QpmqYX
o6tF869sCmm5cnpAGlhwZXDCKblsGERRDsdx6rmtGedqeXw6Az68Ik4AoS92
B+UQxp2m/cqixgohXpsewq/JD12G+oNMELiZx8Ykn4idLKe7IqEnFyyTTdH3
cPZcW+OBj94OrgbH/bKDuNMS84CauyMD1jlKUGUxubEaTDE2rggcG6h15F50
piU85La/CuqJ3sfyNKwAyK2gH2HfNji5ckEL1kl3DIy93VOP39IQQPYJ8MAM
7M0UIxu0FMtXeIzGMDCb0kqRQzQyYvld9WvqHF5yV6X4/n9z3ZkTa8KCdOGo
cmD7s7WG9/3XPnVMRi0pn8dsUR3hL4jrMkPPQD21NNr0FuNj16MvAvDKR3ti
YvMu+cLJqBrAPHcjjb3wiy6w9b8fW4G2xDnD9UAA2FAJYpVhxjOru6qZMxEx
OCnjg36TBcJ3SyQiI8fkZTxr+zZJ72uQg5s1R246oWlCMxbiuS3qc9zdyFXD
UDKWJ37bbsEfknpU7daNTZLiSp0JICWzy+BgF53/j+Vb8p4Y9HvNH2GTeKAQ
3an27nGcLIbrM81i11kf8qcXBR9Zar3pCwg4ZgPltaAn1eWX1KtY11UG7Qcy
q508jNGmQCaPK1zZZxEBDP1LC/jY0stwm47bynrRzXyt57dFv3CfvN8zJvD1
vgq2kZZe0FEe0NJsil0Ox3bIlAHPoNws4AaN6Y9nTaICzQVH26iPBkfgjIl9
kWCk7k9n1VIoXrvbGa1etPgWm3PPjoQ6DUbu0xodo4ZnDBJroUJ7lRJhuIhG
Z68FpiyQZ2w621ng1Wfqs6wJb+xrlRLMD4+nB/xoaxuVTmqZWeCLmGhJehNH
xGGkMfJKQZ52NkFozwmiVAfyTsAAZjhpEERCP4m7qHWvh7Z2LRFmBMySvNJ6
s4W45x9s9cxANjn6UUB5QI+SQpkqj4hTLpaXGaM8YpP7K/0zIQOtEzIfGUSI
deatUGzSgrLSLPDutJr4sCLP9GeugFZtZR0Y91UEEFxsolJdmQ9miJBiLFs6
zSrGv7CtPrYp1XkHHoHpRUW+apmCzFeWeHU4eZcee1xZDpGEMGWMgrH5bOYP
yJpp5OeqifwDzfB+DHA+JmdSNDEJ4rZhXuPGsHwbwGApVQ0jYt7laVg2TgJb
9cCH0sc736wQXq6Qdcp56pxjNLpaYaJXU+ed5SR3fScYamCrwqHAoPXwoNnB
YrB+0WsO+0JC1uQFlNoHubsv1uQLWe/u7OKdh7VEeawOm/Re9Aso3COIoCC3
yAQPrp3JpIIrWOAqrYv2aE00Q2A6He1tW43nv8ZnxZ/pB+hSjL/yDtIXuhje
2gamL0x166ICbnYLFY9xpdr8A1j8y6IWBXYdWVAXrscX+smr7jXGWYS4JDGb
sS1sHrQeJqGx12LI689eR0rJaFnyGaSoKHVBcGDsx5IaKVXWu20hYOrpp5vi
lQdhJdnJ8z71V97U21/+RewGuT+Ut41BiX9Orq2g02AUd/IoZOSv9UMYFAiR
6+C0ALMmCBwSm/+VidNWYZ6eUEpaEtP+3yl7Hp+n0Z/+OdXPknInZ97skUCY
11ntges0GxTRHsnguoZpseRCYCGTMd9JFqW/4pQIT9D4jAPoAYLX09kK1Nqn
FYzqI00r0XI3r8UtJY5OOBc5YSn1N24CNJw11oqPg0FdeEqVJqmUmO281bf7
bs8Gx182Mh4Envs1K7onHaGkuAGwE7RpRI7xbD3mbsBj0tEIAOX+D3Kpzffd
46fhpj/g0OmjtyPF1nU2Os2HDf0SQj+gxFc3C1Lmj1c8RWS/vglBsqQaFrf6
DA4FTkUN+50/jPyfOKpgjEjmaQOMUyV1Bv5zfdraw5gg8zHc+rdj6/pG+K/g
6yltB3JxqIuJBTCqyVT6tcBrKluBprPeCalBicubpIkllufngzZ9cfwsYLBP
yOcZlCvSyK3b/0P7D7e75ADs7xrpkuT1D7U7ptCT0KCidergD26fNbML3UgX
lECyIVj6iUBn06Y13bSrlaOCBz+Ru/UUNDUOynbTR3P30UJPAsWlzijV6C9l
J6phmWTZYjR65WSWv9bwcDIPk9BPecuM6bPqtljXQTebH4/gyCpx/2y6PEPp
IgJWzNTZk0N1/QZAXN7u9ZEl5LODNss2V2xOTW/Ldq1wj96o7XvABs680OgO
UPaQU6b+EEA2OQJm3PYJmFLdJZMIm2NSKtP7XK9yOphT66c6aih6am8s8PXf
lZKRNpYullBjyWGhNtH3n0r8i6IACVkqJxbxEkewR+LJ3TjwO/6cpQWJGm9G
+1Oo4wb/nRBFmhoZbPEgaE/ZBlSJYuSWBgUuiPjZ4LQhtzKm/VYYNa08F5RW
oAQeZaEL/C/ErDGW/1XbjUeL0Rx5mntzQip+9XFEyMwiLUZPuURrQf5VWAtd
ssl1MsgnDpjVQmbhYRySp6AZvSt9UKVl7rnfkj3MmrXEt0uPOEMeytCU5Rg6
AwiVOKgFQvdYhuW+3uR5tsvTdYPgQ2OuQxf9GXQ9A06/e/062zEKlCHS4Xc2
cS9/vJ3i+E2GJibJ7E+hTeNeexJSZ2BBqwag4/dViBWY0p34x/x3gIZr5Dg9
hsTjxc9t01Kj4qFZh9/xyBgHbEUYLLhkVUt6/E90meSouUQoOQ/qGdo2DMmR
dCs9Nx/yfw7hD4OrBd+QjLGsC+XNJYPuZtcIc1k27gWc94S0O1bgOCWeJmaX
eOjStlEuqC4aqWJRc1deGRy2Nj/36ujMATBQQixHQW1R/j3Kezr4kl0Yu14V
8awZAKsvfpNAUAztpJVbm/FhpdzeXIw9eMJRl3531uu5KM3Qj4JbBV8ycqY5
fAimJ8RE82QfSmDJ90cUJjtCoEbK2zJoylqgYgPr5RzZHSgipMt6qqb3kSjl
OqcwtSjrp3qVX0GepMFDd8BEIADgRBHjx4hcGuDAOgem/o9wzEhxwUjFedHx
h5U1BF2ix/sz9tWkMrkz+q2cB+joigOd3evWfwtUMo/x+5RURkp3jOftAj4n
fVbxSu5KeEVO8LO0FjTqA2FWx7EN1VYBaII9Ns98lcDTDGVOwQGDXxMftmwq
n+7aUfkhdrQJzV8/3orSd0mH8SyYSPuL+B5Htz2jIUYRdLy/ah69919I+nHf
Y6T+7u6cCef4djfWaRdHE4TCUtgGgHLbfURw14K1ivLE81EKFIyf5qjEcTAr
AJGCH9HrCDRUi8gaTWpaWy6XAA7ML3TJCGF6MCdPRzEWxrMxalwY70upDgcj
cILfAIRj7pTQOpUH6Bqy68k1SDk62kT2nAvsKr7/c/wwkBE4dpfTmhqwXjll
dP3Ey32vje01itUU8JPXidW3HfdbvVdBwAZbZKE6v0T1yMsMRUqsokRGEMNR
Dq+YOw3MXdJlmiCOLfnQcnvcIjBDgK7UgmJO/ZX/rLQHehpuZooVpFzo4D3p
DQu5bUZFQbCiX6q2D+4fZMUvVkZdKeVC1hosdLItP+XM4eExXeZQac/f9s57
ZYXN2aY69fIX3c7LDu7P5etilXdEAhP9fXZwuydK8SXEyYSUwYroqbD5nBot
dAAz08sq8+nr5AdVyyI0133GbTUgOrbPqFlOoC8YkX1xqir/uG4vqI3tHCSY
b0AJZb8C1EK5wIdRRguPxuUglVvagJE7bUsHykL2lyYe5t1sSYZ+IpOZEG0z
ql+YTLckGF9aJf2H1y2TW/hpUp96hfY0zAfWLimhGlvaiWfScUrf72Eo25f5
viaa/9yW5Yt+pSPOl5SoR3DfvfXD4YM8UJ+bKot9CX04puWsNDwgye9KYvSi
a6dLIO+hFS6kIVoxcnVB7bCcfhRllQ6rZmN7sMwgAbYPmNsPhMgwqxjKTFnx
aP7i4/5cQhV+Ary6r3kY+DiSHJ9ehmQTdibtT3d+uOd70NF9kTj9jIJIQF23
3dIv7IaUkZ+Ov6ELakCBXDievL/gB8yXVNxBu3YU/h33uXawUifSQ3bA+14x
P4jJArFRZduhTXCu1rjPpPyLUWIchyeC3Ka+Qa6cNMGCzB0VcV9VZL0OG7zV
ClXM2kfEFCjkOvd8x56HbXwrns2VQFl7SWjA5PHrCzB25MnAMn5kWzFknpLQ
xg/SLoKUcMMOUUc2+eYVVeE1A2TGkvV8Bo220ZDE5oNX2/ez5CQFEu1Pg08x
ga/nAls48jgNjPwtP/jNOqwbaYI5X41T/S1m5WFD3zdJYDl1PTjNvRF8AY9D
sIVidnFKNg/LHsw+hJzwl5l0z6S3UJLbBngJI6uzHiaIQDCJRD7A/7jNoUPR
hDXmZWq499xp1k4LcgRPbM4IxzcLICrPJHpp8j6sZdiGORBWpB0jPkWbFLZi
j7eUSvxlWtKjLhKSl8lVK7JlGn0apf7v75Y7THlXRGWBfbph/QL2WJaLUDOn
4IWAMa4YKOMVq/RA+yg5CC4lqquM5RgIRRqnr+O+p5SZHtoD9/YAB1oWulNh
BdtXIzyYpvuzF4gK+sSoxSOevuQCmXGjisfxC/+r3VuDrDoc9gzY5mx4G5tE
66vKlWcv9R7HwaSGgyCGdGLReuV+h6t16ud5u7o9Ykyyyyxcb4IhU3yWuSly
maFu/oOIS8M8zQ+vE7AAaASIoOoLmyFTIfhkKohitzPNr/woGI3/CGmBdnio
V5a+kfLuKkkET4YvQJjGbe3jmrSvdkhrSXGHV4W4fYaxtVv/AT3H/onRtuhA
ydLAEee/4Sf1zexvj6c5geGgtTKuiCraEstlobehsZ5Nc4R+1K53Zm03w9RG
Mtf7uGZEiAY82bHTEaiRLgqUkxLdojiHtRS0DDKkTkQism0fBySLxCuZdmjn
3vGgfj865EiJTrr6S/Z0bz8oFNi5Ib1ewxc7EEyk635FLzY9l1Bz+Zt3LWHt
J4eM/WJIDkgEVudD93PhvLq8Z0ShfbesKFfEElmM4ycwQg5SFnwq1EkPZxDe
CftW4yrcCttKRWlC8RD6MfibxWGeC9O9dlaotdT0uOLUPs9So7uo/BdyYARM
UIqUxnpusTySmK1GVQ5cw4YrjDP1Wiv1LC5HSzn/t1vWoxGGoXGpit8mfQ1Q
P4LzKdhlooeH8dD6G5gQAhBZeQoZn3wn7ujAo8dCJWXt5z1OR4l2cfnPXEl5
D1Tfkjn7ecrPLiy8BaQR58LQpgWwOtBIllxz2LUQf1jaWzUDtXCC9qLlbYEJ
Jv8YmCGm0n9PqS1AWFH6QLVuQjnrIkaEpq8/sIrQiWS25Ggz1SjeuRiy3ZIb
zQMxZK9UDA0PmIPrs92E/g/HpUrbuBWy0dth8QlqZKTSTFWCfD7PiaoVZmAS
fSYaXw22ZM2MyYT2EHcidEwk+X9PGSX1Q6UdFuPQqOqp2SUHRUvI/P4SoDOC
o/Brj6k5uHxkN+QFxtA1na2mRtaJdTWqqJW8wbj2rv3V6eRLbA6UtyxwVKxS
SzqRuAXHWRqeIRlaZCulWRp5W/LdTgY1WmxyrVmX2k892/hNNPjYNVtCz/KK
5qRfTMilC6whUYKTsYgO5kripPM9ksAdk1ORgNVn3VA2Ly3rdy/hn/vwv+j2
8lAshFT7x/ufhzXujJMvB7T+hviR2Fbnrm5yth3SE1vlDm8lPRp+k3dS9SQr
x9ODHU99zQFb0naHY3ZqEcojxtoeE8FA+o62f1t0HXNxSVeQnqwQMLF7dFeA
n8QYhWArSV/s2qsW/W3/uN7BskEmWJ4FANvj8P7c6bJskN8kMk+DG1sxsQQ5
1R4Q2lmbZHZQTPW9T/qUePejRBua+0JUjKIzIgrhLI63itdD1mCZZRCSoEoi
u5Gu+AIcoxfkL4yTV9HQwvuPvLzUbrRXomXWzuoolvbnQcyyPY7VyhoQPn1e
+1E8upX6yDE4IcUpRUV5K8v21apYwtbwbktLLF8ZDOc2Win0ZYKu1x7urUyn
oMg2aXU81W7LBA/93myEiY7sNUcRX+lFTTr4LxW05NL5xblvNpFQLKSMrrKM
nXIlGj7UQmJ7qWtxPMxJMpo9IFq+KpuGfhC4XnF8OIPXh5d8vb+J0CHQ1Nax
z+m79F/QmC3djAZTMzldoZWEexiN1pRgRRsb7uRZlXe1++CLj2QaOlSf2lkU
AhRKz/9skRrMDkvoreASB2JzCn1YHXnVGFfYeTf+AykOVf45A5u20KT9+fj6
14us82vIWPGlkUV5mKhLg2VxX806T67uSxXgJPUqpMrRAvt0Sb53CHd7a6or
ySCFsMknEyXyNxSeXoH/aFc0mMrHyCawCLXC61x738U68O6W6egzwDCEFX/L
iIHPlblGku1PeEWwlBH3736fP4YKI/oj7No++Vs9/xLOUCIhW4boDh+TzbaA
/JAa7lFnJqAxOIinS9QX8AmSYVX03s6KjAREy3GyKeYms2Z3oDoyyGI6L68O
TSXdW6ALw7Io/wXwuWW38j9r8kRRib7NsTwYlvgUmPO285H6XGlifk9LPaBs
e/9iAW3HZgzWdS+FCWSmwGsR6Q/MLsG0gBf4GGfRuCyci/6Zmp0duSoALscD
08849d2PHFEZ53hndSwYBOJqsobKcef37Wsb1r+TB5CjR/iv1vIepAdR9Xgw
iNTHGNi0gypO3IQys/rTXD3ADgsmB4wRqXNMyqDWlrY2W/Gy+duutfVFlpXM
a8ZIllFQ+wXdpn+lDXI4rqc3GWWSUaIXi4Fr3Gp9F0uOwTnEh9APmKvqVz2Z
GCahsSXSORmH/VwB2FKynlaNVjut7OOhyeXFWwuZleUkuJbdhdKEYUQg+CCu
EdWIG3SSf86WVlcZR5DmzxEcLvp3VN/Wlye1B5z5ZTANf4qlarpxxmCNLGst
fieQPGMM3q3iIYbGYXL7CXu8AVPqIgTNGO9v6yzoVNpvADt7c9ZVZ/ShwpJ3
KkCgbQmEQ+/dM64zE7ulH0eHsSVbE3WqciuoQ/tXucEpVN+Gh2bsiBKEUXIO
yh/m2IkZiTteAr1d32xNVctPPVdCNqtid9ikkpCEfSvWgVvP2zeSXoFKREGX
u6XMFisFuo0OZP2yNfyoNODCyouvR+ZFlL0287u/aECgmvk3QsaL4vHlFC16
UiDdpMa5ShoZkjpRvqOeMldlbkJiKb1dvOZQWOwcT4IqPoYoYxCs9icI7hI6
iRilI2sKZU3P5Zz+QggytNkJBdSwYYxKuxUu6R12waByLYoThVzDjD7MPW/L
aYmhRBP2vxwkdILNeSmuq8KSXwjuZUMvSTADsIkzHW2FsLrO7o5HsJm4ZJ8I
YZ0zcONQwat6ONzS8R6weyJ1QSrE/BiNn0CJFjAp495+OEgP6fUrcEV+muCU
K0Kt3lLgKr1YVxTeALFuVi7DHYcrzPkIEutljwXreqAwRN7VIRiYwmaOC2P3
HvbX0wSx6ELlW1DOUDlS9dy1RHwYDl6sJjm/8n8BNVNvKd/tn38pZyY6Pn1/
4JBRF3CFUNztnt7E9T48v/2TucvNuemz66euLDYxFWJXUeK4vmok8OWQAiek
qRGyje+TRgpYtg3FshMq7Xq0WCOcCCU2eq+ib2wJs1S0RdodDEci/rXmjM5j
OSHJ2NbnTLCP2zODLwKK2FIM6mvIJfRjpZ0MfX9AwCEz55b+ljmuVBZDKedJ
xFmu3V3Ym44+9bDkayejhqggVPmUXBFxLfgydJx80Yj3k0L9upaqpQz7PrSQ
1KdcrcmePAOymhNCEyGuWxD+Z4R83LWTqG7QR83Xq7UZrTAD4uRRjcsFKquq
QtGRcpuQmwd6cVTDH8i03y3EU8KygtMdW+0ImRztbI3dAWm7R/b4FKyLObpn
X1qC6a+LAmJ2fGNi6ZpBYeNxya7PE4bdbU9Tx9k16uxc7Ah4AIDtnX0vMxhV
ihmjwhwidObKMCFkmUBagLvjm+17Zg4jzQScjXksR+0AqrXfcdZ/OmZWLpn8
Wc+kKS3borbiuejOnVLK3LoOCWuXEEMZ+78dMRLt52afjbCOXhpO3MPOlDZ2
0DH/GHtgvezL3R4EFpDlFW709z6fWrZ9RHYygPjjYr6ZAWlXhLVRbsj08evk
7WOMKh+TDMyCk1y4C/+U4/TCPe2KriqD7EYI4Em0cPs5O5sWVnA577lMd2hu
NK3RBMYmcihGAG3BKn9l3dbgegxvwSpyPgwRIg0+qy86nBzmUOBTs5SU2lxN
F/aK6y3rxdOgLsNuVX9mWVKjgySo49QjDQt/nC1bT5AgF7XtWqemDJ6GuH0L
zR5le/k/laq3OiJaKQh17s8lOV2rp8K6l1VIBetyFAwj8Zk1Kiba9+cHxipn
mOodqpUahFW5dvIjLOrrDtWznsqf8QF+18j73MqxRpvEV6ndpyXYwB3KNRGU
u3s3udwqR3IekUvPIFsSIDxLTzbWpIJBObER5uobBMrrT2aqGYlcbCsKugfZ
dIBAGtm0LjRm2oy+mcm3uwywhMzwCrU/F+4Z+tLCjJn5IwpmLiruMEy6VEkq
YmEtrOseosCupWH016b+KRE5cg1B9Qx9+2sbaBCdpGgt1J4//JB5hC4VaSR8
trdON309qraHMyUgHLNdzR6DfcqqGgGkYgLVZqGYf9eBefj8VfAPfEvAFTXn
GAmhsu4G0vgrhnj53ZTlfyQ3VHsLlJxEdYvOGuzEgAM5g6lwCIBiRjmGHKtj
peVny6tSTX9JzZTxaE8BqLf/+fq1fX2I63/iOkRRoss2byn9BSb5vOCYVIjG
frfb+8GPk0zrTXP0f3xnPJJmmUyRd1s8iZq+MLU/AcRfJ10lBqCcJKQMYWkX
bRsm3+3yxPNR57rEtF/bq+C4XrNFvImp8ljJpmPq85D20Is61kviC/wx2FVF
4nigv+MEK0PHU4BQHJyoskdbS7M2E2oNnp3/+6ORCXejKbhPswae7A4oyDs8
P1Q1NbNB/uZBHhvX/ERKPRXbC2poF89IsjpxxZd2eTHjxRAHC7yK3yja8DE7
lZpAVnCgM+5vLf/EyVRMKbx5unfa3swY9vv7g1F7JWejer6nDGa+ml9vnEkY
soNfLtby+DYniP/0S4lwT8n/XYOqiz1TcYBsfABKfjRs27gq4XWedzgukS3y
+BhYCPl4ZqoPpQyw61vRaO7hXxkOH1iIUBex/OWNZkepwo8bOSJHSjjmjTf8
z1UFpk3mZXCR/h15PgpzDarUgLeHrCkQPLQjMQwXnOggLKPN6XeKFbdpR4Mo
WTH0iK2nlkQVjlhziX8N2HqTU6fHRsNM24xFfLyE+fXEbUMOJvI2/dTi+aiR
AnyHgVZsxAfB9Yg5fSdBdwhr75YIKE5yX84UfK7pPgDIinMb0s1zdE9c0xfy
x6Ls7WZ5gmAZMylGvg2lWGOKTqsj30QYtr3AF2J0TBOZ53AeKTgHBYV+vzt9
Z9tF4sw5SMcp/zAxEAlW/sHJ0+hHSkxXx7/i6EHpaig2bxq8HKYI0A/3ZU/w
BVD0nZH4IqsaOdYJD/0ioIEu87KaNJ6H6f96mAIuR/La1smPXi3cyGNBB0p7
oB8/5QTGcRJ/FTum8nVBvy+jqjRw+3KJaLM+zEyoU9lgwPhnjybX5ImQHyyJ
cVJm5t0uBgXMuXarz1C6C5A8rBEFaHaZrx7wDMMlnybeq1ov6iNjw6Tu4PQ6
bMgzrYqi11uQ94R096u75WwM2+WIim7YNa8NRDZkaTkI76nmukKJheSHW47V
rbLbddXiBznR1lWG0ib04dhOXxSDz+DA24PNNJZbGwZs4wfr/RtIKIRgG5kD
tS7bi3XFN+nI/HJ4ie3UanTltENfyrVhQ3dXssWMXIraQN5Zrtq2Jfv3QB9e
Cu+IheWnKx/4ey0TC6hSIA+AT+mhl9PZCNYFDd8Vsv7TUFSdlAvKHllMIO6O
MlMNhyieIMqH3j99EsWgrYcUXgFFFnhTRb0bckzUFaD7gdzWEZbpBEzy61mU
MZcJs3ccdaf3oHQz7eyBFRVw9aKEyV2EX/AcX86qb2QeUPN+lLnbEV+6SLmH
zRDeseS57lunh/yBGraDQN1bJISOadgIcJkR44bS85Kqvzaymy1c3ut5ls/V
VWRsoZI8CodXwHMTUSMHPwt2ZSK9tKDJbDoPmHKHEkeOkwYY0FOdA2prKdyj
MqUOB6sKTgKDzM0VJmMVF2e6dVNKa68fiLw1SIMyI0sd6XGkfGhLcTrSJ4ZR
5JkpZZoe3c7MgsaRuTXqHSmCVLCy/Uk6G7jF1cbElY5GsfgGWSC83WAyugvx
2YrwvQ3zlM5FnE/TQf32QFcamtP5pEG7fuQ/W2+rmcxQsrNSV+dt+XV34mAk
H4+z+Lzs6gpFbH4SD13CsbvcfTpXS21MsBL4cLdQZ8wrFFCLx1oCuAmY0/+j
00XvELP+MwfukDTTR5J5+POeqwDz+ma74uemRGXlHDSsWsu7hiv0bYtPUeBd
tzyANKAOEB8aUUxBmR+eH1JE775pHsAv/vwVY9LO23C8g7zBHeOP3/mvuZPx
bO+jKX1TFwKPFkW7KqY+Ed6BREzGqoONckZRFpjm1zPpanNuuYFx4tJH1PoT
EdKZB4KdZ8BPUsF1R7sNCsiAO+6WWaBAtay0KGRJ9SXT2bZgrvpWiP03JcC5
VLzMaKVFrIuqvoIdC12mNnXNJlZgJlHOgc50pJcQHIXRHL1TDri84m+W3CiK
EQA7fbFKV7CYUGOgdKf25CR3mxBdGpdUzqMUppt3XB8507FPMMJY/R3uJKtc
NIYx+W7Nos++PeTbWfZhjgSIEFJFb0IZF2BNLcecQoWvm5Yx0/yRtehf/6N+
r6S3wbhWZ+buQaP3IG5BVPWLhAJyVTo6PdPfySfZ6Mgbj1zjqshChUMIlCIl
uyJ87wHtcs9x00KDgQEqVtlzfEbHaagt4Yl848GVIKlJ+rjVJGQbiOV8nQ5n
rJuuZc9VmgzpNqAZ6vBgqX6kvXohPn/AggI5n5lq4ouoUgMu9q5+cX/W1rD8
CNJm5MGxoEi5Htk/8w71B3BNqAUTAzZokIVDlbzJJiNYMphBmuDqZ8CpOP7G
tVtyXiV7n5AqPRMNtl/iNGhk912KeISZ2RDtoTCE9JLRhbI8pI9aNzK/cBNv
0lxYCaW91ihGC9tG1LpMcsydKB53C4SuZoQBn/+AbpQ5kQj1tF6TC+n6clhl
RB7cYpBq7a4rfH3t4FbIXi2bHR8two5hTg/e0DJovqY6fUsW5I8UV60yhYcF
UygXdj90dtCn3PMmrvLZzU2+1PF69x4lVkJ1gq1Ajh+xjAYlorFWfEo7gWow
WbfJcQ4tdY7yZZpiLauTn+HPZU3IjWtFc2UBs5ebXEElpcKL7b5yl4XzNyWe
ZkUfKYUgKqsvkYlVibXaxHPA4aw/fMl5mpc9XZftIZ6zD0vCPZGsuMhetcTy
X2XY5dN6ghP3ZznRRZHGe/WCkjX3zLv3C9pQBfYVqXA7bfluhGWsNisABW0O
w7xfz10OYz1FspHyInKVuyUjZo+SlHg2MOVSPAckZnFyHTq2Y2uNunx1TwQ6
N+zxN4z7iFHpKR6kBo0ilJxryLj8GscIaWNzkhIZ6XkRKWUAs/4f1FL17mHb
Ul+3NFUSa/j3y2a+unezI8WcExNtidLCcwEnlRQC21zU8fjuf8guC93CYs/r
iWdRaSeIyjKfdsIASR32Yo/ikJ/Oj5aIYvwiP26TNHx87oU3YcPyVbCXAGti
UTQUWk+/jbh6USOf32dTGap3rRlG0Ge/VEepGmN+V2CXwzrkZcLulC8O8vDZ
HcEoo7HK7lNZHBf1L5zdS/KhIcyAvBYOqPfgD3x9bq8izb3AwWhV6qpuCEDc
ilztQe5uE8Du0H7pMrt/ty9gMMLUH9851OrVmP9uUtJAP/tIJoA+AygE1X+F
THR8a8bpxKsuq+JeT6JK+alnXEboNabvw08F1V8ZiL6yGch37X0Uba/EYurB
SH37TB79HN7rim47yX9Xydb4eUmqEgSBY1vT4tIb2jmwnnF0gvh5ZBj69t28
jQKXrvSURADx6VlDSjhzNbQeFml+KoDNbevbdhX0NI0UuMKTKtWiUoihlWMu
nCHwYwQk4pXMDQd3jjEWejajHS8C54n75sjKSRpvcn9McySY/6BejeRUcukN
CkqntGlXhZugdroMGvVsfTYX79rcOwgYUjBEPd00aXrVDJd5YzMyIlpcexxL
1ka1dgCI7+vVtqH8r/K/zZHgakZdOS+ahzphXPUevb94cp0GolNGrsCrOm58
cKyLKHMZ6XVbUKbmHDw80h4qEiuHiP3+TNpis43OxQ4PMLqeBp43jR0AJxJF
Ip5ljONM9MYbInVxkJXI+ZqhLxSe9iyt/iAEPihy6tS71MUUauLBliHdPXOb
9769m5hDetn/hxuZ8n7ftxwDrrnDj+zInUkJjoyuOq6P/AM1R+v67AeDnIPM
xRoV0dyRSg2acDK7Zc+CZC/h+/Qu+vXKfoGhPJDxa/sKrJLc266GWQbXmtrA
2zpxKmi9TG3fHFFEvBF0kI3coch0lgNUs/Szy08dx/gUES4ahralW4SoVRze
+IelCogio86DO44vXpBwE74S5NnxhFx/Rm5md8mHvutHSpfQrxCH7NJjLypk
xMpYYS1XfbuSa5gYBuA/lxvtYl5EhMnLfXUFUGhh19B4BXoCRjtyBGUxvYXP
7JyNQdIAIN44BuNcSJwV0dBzuSSwPiki4YhW0CUhOMpbT978P1NFMUtuvp++
ThKoyZJI0sgqCTEjfYN5tU3UPaJbDntZUv1zMsnEWBnsbxNPxm0VIv2fESeU
NzIYnU7iRUbSxxQDXRisF6TbVkCBBftRbWtVa4xzlNDNJZRBmiiUWy19yxvo
y8Y0tfEgOmagzLC7FcMdHH/8z7t5jP8alZaHyzve/tWiHp+c4CEUCyVIbcBb
2AlYW9RyMNWCOSqoWTPZdnpP58mmsRkMnA2CFmW2bSQQyZ8lpxZKnSqwlig1
rx4EJithoZxCcCA5cH0jRPWwEcFC7mF+cMTlAsGAsjfWMiARt9TKv0oA8UE9
VNBRSnGge8qBoML92nltrGzlWhLPdgGUlDOnsYhuscezxg89O4rIFpeXMVFC
Xni7iraPeBpEFYw6iqu+4x/v2h+O9iU8iaERkktdqYtpHK/Q16nDRUTrt32Z
K5f2oW+EAQ/M50ZYruxw5oPvTzDAPHf5BFWv5T9y0oMJqjcEy/Qrl/cHQS1R
Vvbbp4ktXL5IxTTU2xcJF8Ce0LCEvmzE2pOoVGzysHlv1KE9XRTuYmLfurgk
cr/48ATHCA/r8wfs8pZGMxvgudzcUxomc05LRg1qGcf/4vZIbeh44nXjW6Tm
1y/7JziMfQJRwk8dsSVmkQwu7LCVWjmIBEi3Dpu61964LXpCWkHLKDNfqo2u
K/p7Bgxqf8p5KxMMFf1HiWyF+ktkAaJu6CQ2+AkeMf5WYGpDGgCTEGcCr5k3
nX1UchdQQOc+AOpVS9xReYDcFpv94AfDlAKWXJmj19qtnyjWchg42KhArayj
U9blDSbvsO2hgER26jhNbdiki0KnFUpntoh2TlP5Fua1x3mittP9SHa1L5Ff
3eZsRc+/fUDS9I785EzokT/Bg5whfr+awXJ+NgsaRECxtEKnx85fovXfifwb
IZ9qOZkRcvmgj9fQABKHysMhhAoPEogVVnynJDBiEEIJ2NHTsUexAwLVparX
KGzm2JUEEavjsmK7+ootSmlqb3E5JgiQs6J281cfV2fjlkb/YnXQYwR2jV8+
vqxcjxGnPr8W8xRUjXsyMxAjB22ekmG25mP/4RkwZZ3pO736LZz5mxM0wWTc
9Ig1Qh+NraAVSRp9/6yRbFgezOS6qESX3PB8Phfzxxpw217u6aWTd9THyrjc
LBDuj5vnNSaU9UMqM55C4KNGGw44b2/cXrGmr63JawZDvgNxw9lxyNcexWxH
CObHaSfyxCipe+yzHevhfAi6ch56ZIPJ7qt//w5Kv1a/k8dHgiRnGrQ0Ziwy
oNkaawrSqn/56rIOq1e6zXyC0g7NSIDdCSdr0ZCJ+RNc9gwRP9wQda9zszoj
zM0iZ+F/tYATkqRcEG3HoxMm0GTQ2g/MOmWolZf7v3mre9leSlG3KIqstIdw
RMZeUSNGD7sHhkaAj425Tj/zw2B7WS6sSh/hdUPieUvC2kKZQXtww+07cixv
7B2gucqsGDVoqNlyu/ZysxYV9EWPJeee1tLFhZMVUWSD9/K5GXsfWWbh7v7m
VEQzK8vIHC9O8OZKKYQPENSawSS/i3XtYrqEfUmDHsRcLbQ/jzdzobcdzGIC
gs+ufxhz+cr208SAWXYH1eFeM77or7vYO9FMPAQZ6bvY9P1jl9rCuRdFZH7E
Oz+ZcmCdgGrpvtBt1inClEgz2Ir3L5JGgTYu9XPovkMqwoQuE+qsvt7gw49/
FHXtt1lnGzjZ6PqTagk8sUPHweh4/2R5Kwr+BySoiVS6R9EuvrWq+PnNZLbt
hfmjo02cjvb/8xmDv8SJIkO/qsq7MVnLPQ8egJQyre4iomvAB6NrnS8Pk0zP
Lx117osopTUh7PuU/ieItnLrGvFG798J3zvpgXt+HAv2zdBsQCfUqavWO805
DAB505fH3+DcDTkH/gRJrjJdsRIb1B3uFY44uAyYhhj7D2X6sj6KB+qhvxxv
hp4iOQLFZ2D8ULMzQtvYwdUtZbcGwyQFOSpt3S2YYPLV4rUb1fdwh6ILbuh3
1UODfF2RWfXP53P4ZVSIzqGjb5PRlcIsUbn/mgvSEuSdB645Aytmz7KDh0Bl
jsNFbuFNPX9e+ED5miaWTY8HxAcuNkm08t9ZUgvfw+yRmoFNGgqAJ30Dj360
gh1+hZoniWnLQBTOkG2RkntK63QLn1RIfTO2NeRY+dj5I0C02Og4Z8+/W6E3
62EvxazMNHoiWUoVAcvCb+3wHeszP1OsMAPGlpfPNtI9JOxgZ1wiA12W3eLu
sOtel8kWc0EeA+f6s0Fnz6zt6xOj++BqiOcsq5YpDPLlRdOOZJGgyKmBbS2o
xZSOKt2+jeSxNogp/jaCyd4EpGz17EtZooB9TcvJJe9F+KwwmgXhzc8Wjt7D
0dAh4mLC3/7Thz5Moq+ernLqu/1ogdbZREDvQNSzabZb6hK763FH1CnosAdP
cjZkzk3ZrsN6+Dvar/uVmNMEVTqQ1EXXc1jBFL2NhcM5rqWxFaU3cNYa8G9+
+CXrnFwsfVC+gVuSJIsZGeUv2KbdHaPKOZKNbLgRzYDni/jvc4M+ZXbf47R9
tewHcDuQp07qN+vk3CS1FqpaTIMbTS9NyDdaJ7qicPDhfdOjDnB0Q6pAt0/3
dGs72+ClfBFt2pnBcL2M1Nstc0JFcF/DlW93B22+dboCQ9AX/zYEcT5lG+Nh
N4IT/0biB2wR/Q9zSo4Zq1gGrPUKJnCHpnlppAHiuZbBt9Oj9jT7PQWjllPk
Hm1XhJ6+1j9/LA2JLsCcXxCkcyfBzJmLotcPOpTDkvrk8rzzqPc30X0FXM9p
FIozqASkXiLttDTHHLjzqlZZ+F5xiZAXIp0Z9LTcd1l04pyyFzNN1+yKVq2g
hC1SK1AJBEO28WDtSBKsEcZ8s4AQQJ9y9O+7lfj/G6Iupp2l9ODqX7MAIIvT
BAgN+EljlN5ga85r50OXy24SfEhcHPE0kpWzqpfEQyVNvOu1NfSp+Q/CF+Zu
KVcyk0AhgsjgNXvMp4Ol4JcUobPDpcd2dPk+DQdH3FPBySUdIOX2BGfreGdU
mExJQxsQpPSMLtOS/phf0DVG56Vyigex1G9uEriRi/ORxeoHPHin3YJXlKZB
L5VtU/qexEJxmxlmH263FcHfxq4+x9Z544k1CGda+juO9O/ztv5s4uiOpK4d
knJk/tqfo4gF4pneIEWvuvDo70wXBRqWBejAm9qPNOhPDJyzJ8ikQf27Hnf9
jBTzwBM3LkvbyfKahY/ylo6H6Glu7Uj5Msln9NI4qFti4PDgGPSYyex6H273
XvCtie1caFCQg1BhPdJsISFo8BHNsUXDzNlHSmuKAaMwCUr63TiXT9FvdSpL
W7F1u7jA1/E20ya7GnhXgSItxEksfnTK04u5cc2PtWr6OqCK7YTlJ/pT32xh
8XZ2qbc4WwaIYZsi1EEf7KrA7ICpSSPagXX0ItqJgQBsmwhb9PJi5MDyXEK6
/vqyNEIpD1AXmAu/4mxerYYtH4hFk8xbU2NpxTSpEGXu3IR0CD+wavGtKa6a
V2kxLev+E9RVv1cT3LBrOfeBRm1FBJxQvbAlT1ElMld3fYilSsgb+sEgCEcg
wbrvA729gq8Af0w6uGUVkpf/0QfONj9OgNicJGOv3TQxilWKyPx8FbgP09hP
yaqiGCAiig29fb6c24JSUT5TSxvZFClaHivUKvRhi6IIL/DbcL7gjhmOYZm+
1khnKi546gzjfVDp1h8uS8rSRnMWgbxRTkIhN4yzmuNcuzs+fsBiqNsz+gLA
RGgYbKLOPWrZKyb1eObQwZLX+wbQiFKdNMlH27K+B13StAbveb0NPV26/RL3
GpU2Ei9b/PDj+LuujDSaD4+41MIxZ9bdH153voOd5m4mIp0p7ykW9o1IgG4W
nwNcZElKa7OQOQJdM2od+v8MvBGZf0c2nZX57EEnDPWPh7i40lj5BoEqWtbY
ISBlNmh5R/n+fS1YjqN/s6l6+axUiEE+c5G33kz4IXW4bb3Nnsrw/N599lkc
W4dzstKSTk3NfCYfijp2OqU3Jdbii1wRlMoA5o5/vU/IHRGCFYyiEGroQZB/
QBmAyWLJz7c9+Qxbm841Tf6HuHUts2AEJFabhCpaPYcyOmubKE0Khv2V67at
M+h0ljLMMeZi4vAZeUmwLhz3E54to4K0jjFyMlIsps4ItBl9WzaEEhHWD63q
ENJCh0biSGoq1IkHS7igPeK2tYAZnPCKFfk6R+Ptx0pnkru/86f1RAwo//in
b+LuunStrNDj7pn6ShDaBUrYWnUclW0kwJB0tjvAGqMabBW9CrtHs3+b2fSg
hj1EIN3o8kBEpfFpterOTGMwF7mffakh/AAf7RUAguzTT/ZGmfug7dGl/XxN
0gv7JRh/6dq/74meF/pVJfYjNm1L7mrkl05oGCUhhS+/gcUU7ctTgwFB109T
Tfy0X77su8Jo4OliZwuy5Dvh26ox4QZAqgGTwvcU+pYiWYFBlzkylNB8qYbF
6bioqxQ/rElCQlb5rLq/O+6pMKvpsWjHGYFUisKMmQyabOWhnlfwvHw5K1GG
YdIScSkF53SkxyGZ8Aqc43TNDlMcZYBe1D/9jOAUh1mIghyk/BqS9g84DiAl
W0u26vuFjt4GDNhg0X2zEeM7afZkNfvI46XUdTIA4lggwsO4yfJwwJS0VGsG
EEmHkK90MRfugaz7SiGxtzdTJT4aL6uDHALMb/8bcll/Koyzx0gHeKF2zejn
/OpF1LlSJBczRyLUbyFKoafvUDISasAXj4YrbY+ha3Q3A5zDKaA6p3zdgwQA
B8tiAZ0itUn2oeu6u4I1ZdFEJBV8nqx2WqZvsHEQ6TZDzKuG9FEknlCnauFq
TSzmfUNXareoFwrgReQVTtjoa1k9pxg7mNnlnryOmOnyPIyEZ1vIGv5B1sjr
9UCoKHxgyAm0Zg+Wq60vLM1iHh84lOyVrBlynQL16J7RxOY3pCkUBxZwbHNr
mA1nImQJxxBvarbW8wuL94GAAd7ytHudnZ/qdaX+SmSGZ21T/Mj8k56y6fjz
aVn3LvhacHXBSAeQuJGU7MYGuSbVrvb/lLpxVybR/LgcWI6mAYiSxDUe+PaV
CtTJ3LNUqQjvnGH9/n9AlcFuWpPtcvvZPyCPq94JUXAEOoirtSB31Rh0KBgd
2xJmGW9ialw7SIyea0oSBDVNZnta4VqGEXhZf5+xDPZTpL3mm0ZpvI7bc91w
kpnQFFmiBlaFcaijHq5BKDwyJ/rbqYar8RzcDke1yBA/y6KuYKbmbf1bKAGk
3FHHoYzusUDeJofs8gT/+OB8yvahDYrjjR07M7PREQu4qTdSPBjxP2gSzlcC
S7N0cGbGRf4bKQUAezxZLzWjsoEK8VUWC3j16P8hPpAWvVKIKuof2RxLp4HL
B5rR/20qgr01farTQdouZEOjtTzT90gDIXpfFWgMr5HTR6H/P8DAoFA1xdH+
0jqchJ307DxQbRf53Bm4aWat+a3w0+76MNlq6N9hspuHukdrGq/Pai7tEeZx
Mvmbbm3HHI7yIx/xhrSY96mEb2F1tXA39JP195Ls2jJt8avuV8Mb12AOI3M9
ilVJ0ELfoFZ/C/9+LZYVLKUxCx1xXdCLE88gWK9BQbM0B4d3HWaX3OHa0KKA
9GzoyW1i7xHVtbP81Rkd9l//u2sEzjL4tjayOkYpZsn2ZBx3mlLnahBPLfva
+JJ5NQ5Mlxsye6glTGIOwze2q51qO3yY19lL5GVRAx+onMTf5pkGwBfruFak
JKT+3sJ1UDNzmUHmaxt6dyZl/3x89vIbvDivkJ26bhVzq4ya9K0CwfFlTXTg
Hxe3NgvMzwigBj1VE+nX/nSi2gSjBb4P86jav0c01fiX+Tr2fWNCyPLJpBU4
fQLycrX80pZnRQX5RyjLjWZnK5id8650EVdGXq7fzBePf4v82ShwfvOz1FEK
Lz/fIg6+UGUsZh+Wr++Cqhj6x0rzQBxTwLF/uILu1Sn/F4l0IDzljTv8pVoM
kFGcrPPapSIM2l2Ruri8NTzOd1QN4bctfmslPafvymzP9CQAywI2/yNP1C/b
wRKGmATW1CK0+g3cp/fElfDQEa6LTklz4BwmDgtlsuVlmNAq/v8jiuMX+sDE
bf93rKW91Mhiq5nIkhn2/43r0JjuvIhpSn3jRAiyq1fAElgIWe1PhEkm3xVa
3+Nd5w0STqdOWaiygdzsgmA/Y2ZTQkBuimg6P+Fe3RmRm52d+3syPq7I1TvF
/ITZQ6IXCtFbl7/DVWAHslpZPc4ALrlf62JTu6WluymSLRN9zi5T0FfqnzC6
dl2y/O7vj7xrYeBUjC1mhzysgXl7gi1tDZxadh546m2eGaZNlSVZHNx2YYNl
JGJ7zI0M6MOqnntwf0NSmL84O79f4UzIKFRiZx4YbYa3qZmdLZC95dbHkKT7
YHuK1sy8jtslUWKH6GAc27JEpLupReBBSkGBc0kro8JysjiIM/TpgrRA+agK
xhwQg18yd0updqoq0IGEw51vJr1z9LKMbzULDwj4Rq4yTWA3u5tAqjQt8HxA
/F4pDfkrcIpS4Jt3BxFe2mzCPwAbrvJpQ8s3Hx9/yP/xO1CtOKmT2uKTaGOI
KOKdhd4rQ+V4pW35LmKwR9Xt0ch8iAlaq/WWF5yxZX1RGpzpF9yDTV1Kv9nP
pKZu6Ypgf9SET5CLuOAp4EngfFhun3DJfGtKj2UVgaGymvySPGLbFrRJR3SA
DBlPzCidtPc3JujFfUvONv5GWFv31ThreG1QQ7zWnSiPeYo4Bqz5C2l4LDXy
CGe1e1Gxz9fFZMoeVVwXdo/05vnDhdW3uelRc6ZpBW6s9S2KxHQDprE2aeLO
HyGk6lA8rmT9Zfe8CWDdyHQ7BTR/WOpd98HxKrsqUr2JFpZvJJIbmPcgrMH8
k//gPATZTpd/Js3CsOyg8zqWJXYPiOKvy053QiiCQ0Cl4UEN/BVOStOHJf+D
t+q4sWb0C6WnsxiToFnT0wFkzXSBluAuZVL0SmS4+g0MCiYkL4p0uN9gjBb/
Gr8LTpiWft2iYyEj6O0Ltd14L2Or/IWmdvbCaSgLaft2HLvRH1aMppMaRhlH
6NgFBUqV/Pbasiwb2468GZmLFfKyZuSqwUwotqim/BhYTC9rvsdp4bIrnn4g
AQb9O9hRFpqWcfFlJrKgIVa/KyxJXGlYANMzcvbF8j1/z3zRAwlphS7/Rh7W
8aoYhDc1e7gtpla8SzKuw1B5D1+qVlCKm1mflIJdbSM8dSgTXL8H2b0iIDsM
35akvHyp/hmJD40/ZDdDyZ3Qd5f0jie9D5i5OeRfWeWRB+OzzHUUgQDaxv9b
QbsReTKwpm4VB/Ph3RS8mbGlfMKG4++8LDfjdh7M/mvMMK8oI3ahnJrPt2TB
SxSrhiEck6JGyv1DPX9fUFdGRw6nDipvrs6KbUPd9Cjs+GZhp4kzaOZbbc9Y
MP9skQP06ivbYy4hQUr/BsBYjf4WriesSgAlza72pJGhxMsOhRf0ds8YGMWL
mszf2jMQDGqxffwhlEi8w+MS2Y+RxSvhMWKtXNn81keM5tg0SQaE/PIze89m
C7TKywuRS4z/er3GMFnb1QL3yh26QQNmxgda4FlUx9tCzO7qCBNRPl7nqGcL
v2LmJJqg3XykOhbEBnYPdakKNNLw5OqDA0mEgKPDWiXe/tc9zsLY+uKgrwIk
jE6EE+lDP2dKfx4SSAEkC4EXJE4Hole41MLQF2MJ1T+zthQQ2NPPjn6Fsz/D
x2sEnGT7iMZJebuPE9xpGRwxMrKgIxc7LiokybtjP/16wnPgcWLgnbQXIAEQ
69jDmAv6n0j4Lber0iVuyjeHiaqFRVXEqZFyYwJcMq0aJNh11cwIwUBHtbr5
qQMw9ijYR8GKlcZCP2qvv+I+cvB/lMiGI8GrOheQMjPha46HGXPsKTBZb8eG
lDbwGcPyDKlVA6tsE6PiZ6QrzaNzb4ukQekHJCOxSIPydNBmq+N5n9+YvujR
akAFMGbsksACUKJx3VgiMCy/NKY4ACkWlZG6RatLgGbtNDFtyLTu5qFHeeK/
K3yTaT5JuAQUR5qPJa3I/2xKtCQQUcyTRmln3BK75IBm/zegjHayNPnEjQu1
4f9oCgdYi7iI6ZUQQ59wcnPI0eSvUxmi/72xrLI0qqRt3KlDcZn/6vy4tlgC
IKD7LA6d59L7aFgOnD0QFNgDrQSEHjpo75vZEedBH3vMkD8IAT0SD/BidjrJ
aFHrCF8jAUW9M/cj5THgRDFN7WV8qCnIj/VX8fMFPaOF1gD4K8Pero/nFtJl
osxKPBD10dydxyZqDwtDARw/m5ClOPV7sZCIVgpOjMH+hsEgW5S+eFQOsTHz
EtyOBmrAGL8MAas63YaYtWk4W+d7s+CE4YEB7zvdoBUwynFze3yMzNUsOiza
Eka9wbWlAAr15xk4zoPT3IyVwZ3shDOXFQHH9H58zeFDcNAsHbD9s7IRyByd
UpXSpTjCvOknN6MCviW4OjiRVh0DtZKLIAZEqGIHfmZR7+usI5kQ7YJ0cl4W
R8SD3qCXH7o1BDdi99Z1XlUiwk1NhV53+ORQOZH6j7JLb4bWLosCNZvw0DsE
SXQ2E4gZUxBx77JJQLJm/j20QfLbUbiwwkYiBiNY0avizytR0fbkmR8A3IxY
Lx0cqNTTLXtcHtTzve2JzuX/bCQ+6ym5iL1KyTfQytIec924XFIkW3CRqC4u
W+DVvffvdw7zyG9Wo5td2ZJLIkimaEgPTeHKbtsFA0orgxs/U3H9KLzwUqTs
1uzD/66Fn0A56d1YnUAzyMVy9J9syh5DggdttKFyTwJ3EVs4yz63ZwSojxxi
I9ubbzeyk+d2iTi5+laiFIVRY9QwRtNsudTDsU9fvqos+JRBUpYzQc/ipcMd
KSBh9TZVS1Bgoh+AZACBRmJpSgD8FrUzAiwCt8/Ti39H3swZgF4PoZdsFoPE
Hp/aY2yScvD2wbWAEjXtBiHkuOBlSFwmz+DM7i39cEJiO65misT8JESGJTgv
A+nPkm8WGSkv2zt/ZLlJMXgL4qEScALXPC4f7SY40lUDiCWJ0hTz85nfDKg8
R429hdOHmhsGrYDHU21ztyuGkCoPYVnoEYnYB0zxmLMinLYv6fZhfTixM7I2
yMIyvoL54+cALoRB1FFc3JOsAma8SO6plS0cdt06sQPgJszoiXUfzAS6rky1
KXACEVLkHia10pAeLUXKEMIbx7VwLEzxIn7FsNSR6FoMQizRVH7BJ9/6NM9J
fqJt46pq2wOsEWhIzkXGb/ETqipZxRE/Ur7PI08I71RWhgSjs9/rJQkRfjj+
58V2vyYaLk1b2ZPC12UxgmY0K2w5UyLoGLhwAoFDlfB22OXdn+Z0WU9gTN16
lVby+YJI+PxDEhj2gfbTZTO9ygmX30d55S6D+w0I3oQcem0rvIVXTM5JCPbu
GexnQwB5h0m0xkGC1IGdH4KXINLgE0OULVj8uh4M/FzFys3VMKmn5VEsU8jP
5U1wtQhnhCQJWnxtWrmzcF6RRE0zNDg91DcRZCir9f6ZZgLMGojiEBENxCPa
14LoZhqkKWIcFjCJTjJLUSihuI1VKd8KfwXYBhElZ6e18NGOUhcP8aNSRVaG
OOex89oXSQZ2YlKrE5cJu5Q6SQpHc4q5hszohQEyh9tQP8sPVGXcPT63Ykfl
4xqHJXXKSBkplTTvNBHlJ0wh/9aixvBVwiQbPFMcb2W84Mj4nFjUzmW8MYhW
6bASQ1PVa60DMnIB1jhMq0XFjdVmKTLysWX6oKXxCeuuHnFqQfQkqPKfkF38
SbBj9zXRvTzfskvI3PoV+xgOdoQJSoIZeC7lJJwFfbWAuQGNAlL4ie5S/4cY
iKNXhGTJz1yDLkrIUwBFh+IqyCkv4ypa5mUDyaIyVP25DZt5sPEVSuvHqEUS
vSnrVZpzxasqA+uXUih/edKQ17s6fdBEYpuaS5dnEjY2m2lIfpyX/qvrIkuN
2KkyD6Xce1dniTeNps0+LVTbySrGdjoyJmmKOyisXJi+ZuGQsnHRWBFkcsS7
PeFUuwDQmdkmHz7pCUzrbSqf9XPBofqFNZzkryOFMyQNTXQ/V8IdbpRqLKVC
l/Ic1mxS2fUgqPECArVOs3jkWZSPg2dPQPos57GiZahzxPoc5Hzp6Q2bf+qu
Rgj8V8McW/tVkswsuJgPBvaQz+8/+PUQT3ACD+DWTdlL6kKacgW5FixGJG0E
m5FjcqjMPyqxDkMxHE4iMzpF91unsAgkmaiAiCTwNJn5sUXmhK/7Vspq3Enj
fKy1B7lwf4uIfWNQzO7Gqv40cYGZTtrifzEFog1/3ButIQIAhHfixQ5tJ1Ne
Co+LKzXjY3Sw6KZITsiAEBywvuEKSsvNMOfHF6dDv2P6PZNaw78UklUxFm/8
pbKfYSvIMUIWciirW8WnS8It2GUPGmJD19kvIyU4qz8ssLYqIixGBzNOYsM/
/DgGnq6mff/4q/PWSBK9RqUZIw4lwGxVf5UYIUzkIwuC6SNFcZfzYUZL44a9
+3NrVMhEG+pGYUAXL5aPvFQUjFVa1JuQPghxcEaQdMpboEVDZUxnwmoQIHKd
VjJyWrbIQdHDPGM4/69DyYt4DWtDdmvsN9KRAdNX9Elcb9V/I64NfvkCztKQ
bPJUvVLrmTElasAReE64EGUGsl31KEDItFqdsJ0+97XBgQwV7zA1kUlMRl98
rDROej7VbBbRfYOqSupr5semFPEaBI9ANYK3dSl8DsrEanup8XUrug+ksLxl
bF4jdRI8jEvg16B0QyPs62ukRSRFabPZxnx3HkCf3KgPRuje8lUBv6jz/1dh
pj9sMWyhFWu8TCg0xB0nQgfJablocyO7wq8AHB5etYX5UV7WwbnqybhNSpc5
waJJuDVXPz5T1CU+7aoXC3Mzdh5QC/AGN2hYp2dCy578Qs5e/5iK9jdhRqZ8
o0Ix0y9JzZVin8ItTiS+MNRxBLFkD4OxB41rjfoYhb6594kbBAoJX3922Og6
g3a1bA8B9H3G+E1llsfJTQCelC/+qD2MNg27k36HK+YHxvb0Alx1dOnQMALo
b1l8BvCSVU/LnUhaBAyQgwr6COMk7z5ULq6KIK8vjVPAMFm/JCk0UfHaKO/4
x+oxmU/mfDuADUw40H7zq0J3oiXbQytb3daESxLAadDN5sPjEkMutNnVc6H/
xAk0rSSCn+D8JM2XICx95AAVQ6W9jSZ4uUcenHzmHu7OpPj/WrVd5GWoT7z9
jE6L9OdCo1Pi5v7Y6hpDH+GT5HIwrlhnNyAKZJdZOaUGdw1aNFtAicfdYRxV
e8Gs6dqZaXY+Gsk3SNWe9IjRO8uxibGHlcgnBqEGdubStSputaCcNoME4D0+
7Wt5K8uG5aEO2kBxPBBe3K17+2086Fye8fPucty0mLW8vKRFugHOng66HYGG
8BwGMfSK4efkhSvsKzlPjITjAY4ecxBo8fBWmDCPULwbcglUCvcc9/8VGNsS
t3IHtHHciB+WFNNufC/nxx2vDFpIMAR4rBHgM5AZYM0CRlV43sYEC0a2lljc
mMp5VcRlAEvDg+FoyIkRlfUfg0TckcqI1uyBZBxRSImB7vEkyAQ91VkUeRgS
0xBBGGlI0vY/cNj/4dHmQjGVuuTNSUtlAeDHt7byxLUzUnEzp1zHedEcTxA+
MOZUr2KIfKHFKvny/WpqR5BMNb1WU2Ig1c2CyLyA2CpTowxdY78DVXYSU+ux
6vOCdrrB2zS9QuEtNmaIzQ2RqwsnAzGpKHQO9b+03bCBuDDgjnJNPq9IGH8n
qILX+pNMt17MFbb1spLslYNZl1NKEQIlsUx5Ec6enAZo6P04aGe8zfyndv14
FgyrJAOHYq/yvhi2ftHdp6Fx9JqBPHOpzKtHRiVXTBzi4kXCP1uteLs1ISU8
PJYriBcZzMP4urSX3d4xbcYhW2mN9rwNW074Kt58QOWFgSwxHJ3ydvuzBjxj
Bq9TnyFCy9hi5liNTlgaWvZuLZ1EQRdwdtfVyUPOzVebKksoxOQRxpdCOfey
fKsxFQIkFItp/Q47vG7BloYXcaK+B6AYc2/yAKU91rniNRRF9864LIuVMHn6
Wz6FRNNK4JWee9sA/u3fySsmsNu7ONoZEc2kcj2UQUyoSoe5e1iNaGY+1Cxk
nAHaf93ppAjPgtUN8SXvnLca3pkPoVD6VDen2dwC5yvuxzIae+BC0o6Dehui
sgRP76MgwI/OI0gtLsWPB4twDkPtGjtuLeH3of1P/L6Gq4C3OPrCuqnUI666
wcGHMy/zs63EcJvLsJzy50EEEDV0TYTU4WGG03nTQYm8qJSxkFxqVQv3l69z
MUuAoek2lowthNTMYetuoaVNczgmTdeVz3hJNrADX0P5tv8Dnr+wCAgZwZXI
G7SsuVqcrYkR1hdX3AOuN3VBG1y0Oso8lRtxeaJMIQGjtMT2JPz6HjBv+or5
eag6jAHcCX0vZH10Ueyj+fSkTJGz9kXaSbf0VL/GAU0NuCt8DeNILzc9x0an
Dh/poL92Hw6s6bdF1AbMcGPf7n2PyxO3YQsZSWU+oXxyjlX5UG0hYORKXiYU
ROn4TJi8fCwhmVktsiesmyfeFxuo71+NLu+ZQtN1s2EUUhvMgyNhchxSf/OG
iZINaJxbMmvlU/BVZVdRxzTWIUSQtXpKq/c8ubGARvnP+4osqLnl8b37hgvp
p/9Jdx8SwiWjxqpGeAgqoK5GMB/ovzQIpx1YQDlRez+aqcdBtHcLLREMJ7/b
4eyxhg218XzGXfmWCaRo8bfMN69dz79+Em2BkEeanLOHOAPdKToo43hhkcug
py/502K4CuvTNiPvbn5dZlhdysO3UpVIFuSNpGrn/WepI8A8gpcwJWlmYvAL
q9x2KZenE3LtbU1JDgrSeTzaiU0b+eA+hppgmf3LC2CnesgoSy98Ekuz4sIT
j5LjJ6ckCNpkdP2V5PM4+6AO0jAJOVVjvIIRUgm1HAzC3TgO7AJfrNS8/phi
QYJyVW0eUTf3BghK89q7IfKJ0PlUWuZr+1fuiz2bupVM7kSIZAIn9Z0esWGj
IPzUDwQXAW/6m7o60+MLNjedjAoeHVo+dOpy+Pyl8aXKEeFsQPKA91s8RIcJ
6QIfS3NS/N6FAs2WhE4p46n8SKPsdBgDgffONnCnsAw+r4NhertwS3E7lyi6
O2BpsT4rhpIvXQ94aC3GjNgwl2hSHAaMJVER5eF4BNQD3J04WahQ0sHk2vO0
c7k4Udh1Rx7KE6xZpEu6FrEzYb0PeKY0jSKJ+LkX73cKyyIN4XZ8TNGVF82F
ANftSLusRJs0f3nem2T9/M0rHF8ptX6jqxf7Uib16lul4k4Wmq5tKq6CF/9D
AUK/rZpAyABDUVjmvV8uzqLfutmAZobRxykoha0zaKs3UZR3Gi3RFqHVZE0E
g4DXdQv/s9Jg1r/2jijGsBgyGlIs58gltej6EkM7DBlHgjq6jDZP0YZmCw2n
RO1tPDZPH9YI1Z1ARhUQGwqKlT3elqMBgVJeINwC5FTVhpvk2IMlrXjGzixG
QFLbsp7Y3riGVPWc7MCUHV+EvOtosodpkwfr1mA5pVPw8VqdvN4DduU6rfDB
urm5KHIrq9pAbtnvQPYJNqJw3HPDsUrOZ/VEwx+gVXK0TEbK78TMLv2W2EOn
ofsnqnSFVy9k0OqE9s0J3qQplk2QTcteC8zic8LtcrBMT3NuVVpPzS5L4UJ7
KDTDr7z8N09TCMbMW1cHv15ir4zT7d/6qh2M6DjakFXhta+IfC902f23CEmj
svBLNy/NjxD27vJoHutej2aEnWeyhULRfJe2AZMX6+4XwArPmuo5PDKbzusG
Cfc0CwA3f7UmSiDzQl31l+OmM/dcPgK7KFl8/dUWScUivdztCB+GL9dhmO7g
lUgzB9iVMO7HernyyL+cTf9p5XZcsZSQ5rwT195XRzEy9Rc8+MhGcoKMEXom
HwQbSJb1Lgcy8wrb33XdwhgwUqpR8yxIrKg9uMhY8PwZyuch+SelKK4LtmHm
Bk1RqQmmfS0zeWFvqZqjMMnvcWyGcJXDx4+r53cGcpFFEjgVeu1qOfT9DC6C
pwZ06LG/ThCNaWTGc1Qc5AsqzDdmdP7hckxqyEmpodJW5U7riYrBb4tuPf+G
IZwYWqqu5Pn6tzKLG9R+etDwbKN7rW560w8Xv4hN/H/tktNxy72iRHiS3lRk
UOis405JL52Va2iGtvRW6rALfN2L/VKfwtjdo4mzQqav8aUAOsBeYSmjVwwO
IrRv37jzbtEzvHpKI2Yphb1ak3cvk8cqeSOmTWH4hW3S4pLFtegA+mHufeLA
njpT/IvfRR7TYIgCAZ8GZ+O8zOcwwEaXbglZodU7BCqWPhO3W2dijxhIICpX
74oh8stmYnpXAu4aolals+EhDtQ3ablq+f+jhekuYEsIoyz4wFoO/49YpXwl
KI4HmMVj/vAOBS5sRrOt7cHCGIsb/adyGjJyBx4q3iDgX2jlFI6yWAQo9D+F
3VcGCtEJk19FmsDD7m3oCT03NzmjIeXjQxBq5xc5iaEaVPfMBgW+Sb2VN2jU
jvuXFgV8/VujGj9AGHDrKhHzknI6D37Z8VCoydMU5dKuwUwi/U1u3kE4daZp
3sY0NpZ404ZnnqndBa30jBwFHJJb5DsQEZhEzpe+Xsxl5Ejb+SYoLvoK8XwY
05b/ylaeub6YMReufek6smgX8Qjusx1rZ+jeT0WX7Ut7FO3hKhGgcZcsIYhP
3dKfri7CXkMii0T9N35+FRdzhpXdeRHonC7K+c/zi1tDt/qWV5J5Mro7LYXp
7iotnlhma/v5GM+stLAVOUGLHFqaCMEIynlSax3ffZ0glBXjD/sh3XY9Uavs
1RK0Umchbyzz/YXwph7dRevy4GZvGOSq/ypTI2T/ibhIx1TpRiCddxQQ4TZi
TU9LpT4K2GIqQR8QDHhKM0Sgh9G0fkUBNqHGIs4PEYZtYkBPlby/lYIkNvlK
FKA2CN/k6pOGScBIaDnwdGdfceFjDdQ5+f1bXePbUteANDn6BMaHvLwD0DFl
YnAYGTZcSX2+o7v/ehcW1alBID8HDgCCuPD7/otQHt3Li139/Q9dcND+ArRZ
o7y1RMbbRu2jnOEc/kFEkXgGW2vc9cuOYzKrbBJ/wQ2Xlo6ALX0aBoNmtIVv
51lQswY04BeISsk0NEe+8/Z6bTkq05dYGGLBLL8dVq1m7J7gO37U8hOTgyjP
DaWpC8gKM42fv8KAhe0JRPjnTbkhIorRwazKKM1MD71+C3FciM3LD25So+2w
QG0QJBOOjHuSRIETzJWExV1bziilI4Acxp9iUDnOXirS+eARUh2KAqx+MqFE
wtiPdD7eSeE3YlwMjJdAbDI99RAtoyVqrQHhF/Qf44OR7FkVdXD6a+IrEx9u
WJHcd3jWbUEbAK4brw89nUZJrW+jovpYSrSs7juXjU5FOn6LIEVtOUSkzPn3
rUgo0vu+qt8kPOSamUOwKW7DbC4297B5acAIq2sQ697tjz1za4i/foHz4FnZ
UyZROksJ4cOwizAdL6GdmWJTK2EsVGou9+dijcXE34jZdPY9gv+7YGTGhxfb
bWnlOU7aXrAYHFGvN1g4BAPQqPXQguFI0YyHas9AdJAv7GsKlgfrvDur3i+K
MLkLFEvfKkkxovEItd0m5vAemENyQxhr8bvOWOKilAfPYkH5r+8dTbehO9OT
bO3mZYnlLRnojcLgOxtKjDIg7GsACozQh+5jxY8nF3zLnu6XftSkwBp+rarx
39im6Yj0y/jWZU69O2YwE5mWkgRhJ45MYzIIQIg0y9Cd/C10iSx2dE4Ttoqf
UuAjtTlwBM4PLtDo/WDG5jzEY6vHcq4KWBvy38f+ehpsTf6Pl5xoniWxSZsU
IojroYwFZmp4qotNUoB2MObdrH2ucuRu/X0vdvzrLWNrFhvUcut33Yr1GjKj
qgoo+D6Y5slAkCwU4lVCrwDpn+CzGuurM2JH3h4Ycn6iuv3mEetokjzXaP5P
YtNEOF0F8VOxhRwcEXiRSzFGQK4dQuGRpvps64nBc8eY4tKiGtIdWMBOhGRG
nQYXLpxfHKoobQoznt2bZMMZ5H4FOdel4RBlA4kuL/kXlV1wS5Z1sgHDpLz8
dcrCTucBoZwbtsTNFmHy5CcTh08HK/F9/230PD9snn8dY/UhjacA7ktoy6aw
gHJsKFOGqs7OGSE2XxrNBZ2PnnpVcJTypWMOyouZFczpwkZMU9uRa5kV82fX
KjBbXjTk+lis2DeWnx8NP2/fjjDTTdo8ff8zkxoNqWk4RSAkhLoyVRTM+VHO
yOtXLLZwT7RWRiBpqEQ4jzS2qHRucwcL5ZTXZFJLdkI/EeYyN9zlhtConpbf
IIY7Q0UNxqBbSQXZe9MhdZRnrQZnCN4m7vOS7LGKYXvSJi1Zv96RDOhh9kjf
+zu3clE13v/vpyX/Gr9U9Rq6Tb0sgfcqj7ebTV3/WujHHFU2IbdnylcSGRjE
sRWTcxgbY8A3YEe3XJZQanoH5ZIS9EGNvW5m/yl+pOn/ats08zudqcY04grX
bHlZtdw6u4mAVMehz+eq6iC1IRju6b8IDpEO5sPfCL1SLKQ8t0MSY13yx4KA
Ijfw17N29WqGSFyiF2x9gzgjsvyY2o972hoIQN0b5CdZFhVdRWg2TwDuiZgW
zQhJij77E/gZJIhlkCRQECR/X7sYaxFHM2cBq3dtpdqhqNcRdH3xyb3CN6Pb
hKfxN4FvPRC19jKHysTm3dPZn1loHE30rxWEdjiRSlbOlNz9CJYhZRtyDgCf
l978zkEaAVQpy4QTvuw6BswwkoXiT757VvCGI0nqHOiO5KQmIqzHP9EH4q76
XVsA2P1FccU+13ep0pQH6qCMj5vIceUQNlBl4ZhWmGw80Fr5JuH1U0hy+vum
5VTg6gPowwZNY5ewi4Tni4KY5OAa9dR+ZpKg28zTI9/k59QJ4qj2KRe+XYqq
h2o7eeDOecMUFRx8ivvqv0QrjrmcXh3D0W7AOVt2Wm+3EX9Sr/P9I6ekujTc
ptg0umq6cfGf9dtZK8IaNQZfyb/Hii83ZtSfuifR1+qegiEOPMLg+kfA1SA/
VwgrbuO4GCJmwrYzITWiPm0C2YCyhW8g1+zXDwaFD5i9S34B/onMgWcf0RXc
sfyY2nsKACxRf/82zgoZxqbQWvXfk/G/Uw3VsOh8xZTihnDYDNvkQpXF6p7c
xQVlxqicnkqlT2Sh+iBwije8OrrGb7ictP3sIxH53n8FWeBywVWtFObZ/Y7C
5jpinmotBL69iKCTHtA0m8/fKnR3pRMQodlLQof+UT3TuF45EiJ/UuwINc5D
1jYKjqqe7tiClVtY7CsVWajnnwyKbOcMkOrn7fpzguU1oqb53ym/jAVimNWX
19PFSl0JgDJqZAr8YVll6/1X0WbsA/YcfP/x9h+L8lrpljw2vyeult9EPOCH
arkYDqSsdZd0dXjNxJAXa55sib2gNpAloSNsqIwtFhiek7XKDcHcMrBt4cAC
srlIT/dFiLRaq5adRR/qGfpYYtr3d1Dz29kNIxuSVjJ9WIyD+JdsgEhhI883
+TcNzfSTK1mMhRxcXCEixW//nH69NBartdBk7cWvDzj/+d+qJASNBr7ISTM7
5TIqUR9FNvu0bhNLKAbmvG73WUFJYnFr7DNAyLQoPYvdSqgxD3hyB5iCB2Xj
oKNKUa/EiXdd2vc02iW1jQsfXa4MPyvIxnjgY+cAuNcxo5V5cvrbr+OkXJeK
ICsLPwVCvclOrEQE+ib+Uk+JXwtmi7WTD26b/jXXuEX1eW/48g+A0KXdBnCO
oBmsU0kvA80eTGQsqT6X1oiXObl0mMEw0QU5ZWqcKgGCL2mxRpUGrx6qGJNe
I9XRy4q3xy2c0keFhw+ofMXi0V6Bg66JwCNG6DN9fb+m6cSOdIghRGHX4Uuu
FlaO48C2oV/R2A7QtBCfb1UNeetW1EM+Vz4fBFBe1IATstb0DZqkuBkHhOkD
hh+xWg/z8bBfeP3pg5It8Red0EEkTCtWiaycCsWSvua1yt7QSbwjcy6dfbEL
GtI8l/KsbCn8hqx72t0ABUbsLbVg6xv3/C12PUhZmEKTfOZCa50KMICMtjyQ
Ln01eLWzWLHhB+OP47i8r1MbstcR+rFZNj1XKT9aqkYmekAyUlwGoiZTWO/Q
ZVDxtttLqm7rnoY50dutVxNRFMM5M4+lv1PsOscOOqF7m3btE9MngIbnThPs
qbEVHMfkgh4KrNuzqx2mp0v10zhJdaWs7S/b8AS2Jkr5yQ+qiq/N3O9okn7g
PkrGjlx/udr5NDCudhC+8+96IbQrDXotmMfYv3d3ozEZAoWPaAYqmSjvbbVA
gpFuxEdMZzgQFw6h6WU0XLNc11sK6QP4wOIbHqf8cvP5IuGVg+mMkQ7O8YcO
sLUmzLvjw5+h1txP91H1k1i7hxV9kTxvhFw2z5m0Tj0oe/MM4Lq3ZrojnUhP
kUCaK7Q6h8X/PH7OmBn9Bg5FxW7HUiT99tKReG0MGQcplFOqAHGCCiLQSWrW
F+/WfT3CjNAYZTjlMcmWwO7ORmSKv/eFB6fR3AM+00oolmZQr0s1pUePBd6C
hHLe+uauistQ/+p1nOsagB2t8mYHVkH3gZHzvL52hXgHab0bex2VKuvrH53c
bfYS654sfeCE2IaXKMmv8Cn+RKkyXsGRU+0AGy28l2o8AK8mdjKBBt74qj4i
0LF32Gl14d2Vb82CMP20nVAQ5YADjOa50HM94h2c5orqGooNC6pQoH1ReBgO
Bgp+wewrWksO0nxBLn80q7QTZnpF4/K7CCBxbAgCn4MZ3Wtb0VgCv6XCaBYS
7v/Si9916VPOhaQIToe3pof9xsS4f8t12K7KpOIin5uYqXWVX0/YIs4CSmuj
yePy+bsb006HGrqg2uQl2WpdpXwke+/yzu14ZwJPNaXvVlPs9Y49zDu05/2J
gdH/iLzV1SICSR/fad0DvEkUOKfb5DhJKs07RAoejdiLsJG+Q/L0al16XtSC
Jp7MYBq7jePsjaXXFkSs4dbZoBiosnkUB8ldhkMNZjCf7mVCyxGwDsoskENW
FCTXtub4JWyVeYCzdqmW0twAu+/uuAiqOtR0ohRjLr4Egr0XU4krjc7mcT6Y
yO/VdplTzAMXjCJ2hbkh/Sw0AUBKVSp/9DHnpaqO1TSBT8T8O6jpg07uh7yo
zRhoyVsTd+RRMu2TOvbu7IrKDZPq+qBNdBmLtUBLNtQJ9nVoZoTt66s9AUnC
kUxhUykPKpQhMdPRW+FJp07RFHGj+46txq4ThnvneB5pPEjj28S/CmZ0RzNe
WwUSJtbd5AGH6v/KPlaW/leBurQ/TeOgJs6Hn4bNaenBK0qIJ4X3qpRHBPK2
AVy6TxVlI8VbUBkjLN6aiEk3AXB7JYCRtqtgdD2SX5tS6K/kyFx8JBBFa6YT
xnfZEcLxPoxVokcCfYrjn/pQrmweyw2JmSd43sipNtaGEEiwjVtQiq6yRIOt
8Trrf8BpX4VFRyYIs31QSiyhOO1cuYMKJIcj4Ey/rAbZe1Vj6ANJeqX0b9Ub
GWmAcraDoKKzUNwSQ1MauTUrRiTCfrSxzmo/3FTNyL6wklKJIcNjYJIILL0Z
r4D8qeuwraVIac9Geb4VJPEI42MJM7pvwdOpGoVKYsHs29cuiD5zhM8TRKuu
8rW03Q/BM0CS2UY40JEFmdXMi5jw9TWrBVTZiU5+J+7dt3WpMrEZ3H60oxmk
sErZkWW5q5TWKm6baU5nuybVWO4zHNcvLQczvj3ZKZuLzIluQ2k7Xetm1Gzn
4etlsSz5Dgryy/fN16QJzFwJL7mcg7HLRjjSocO3TUxcij9kWWNp+6sYAvSt
a7qEI0+2a0H4BQca+xA8lri7K5Z3qqdgzUhEM3EuO7g9UjwKyLjwnEa7TeAU
4nCrzQj9PdDF24sMoYGca5XLemrg0pbFpRuOeIKbJ0rDA3ceL31Hp8uGLyTf
P/tu78cDg+0snSAXtFdbrPrxafNv60sa6ZN99mBH/Wp68sPnki3t3e5/3V6h
GGvZAFWJAXcpRKbPQJfYm5xS7ND4onqFrhy4AOVWojCM01FYWqkcDL6CV1K5
qpVr+RXb9+xEXUYfaOebFPFcsNhVsSYkxkkT+T43855hwxptnfl9CnV41fWE
hV1oAS9DGQ2rbYm86m6za4LOLA4jYMmNdzVSIdJRoMcdZD5V0CGaRejxC3eq
/MTEoyu0oh7083QJXCZTcZmZnq8aqX6SFuV2eAyBt0cQmkEwhQoVGJYgBCrj
m1y5xsGWUTnn6+wL0RPdnDRJN6I9x+fWi4Ca24C7R+QVl+Q/L8G9E28wkcRD
PZ1JfZRyTTGNy9NEsUue71M79+hU61aPv8C33bisMDZSYGrUHH+4FHuvPGzS
PNuOTvagV0CkgtcuovwH3KqMCMXQKYIfdeKIY3K1gAixZUujl/KL4nRgqy2Q
OH1Eq89nWfEDwtZlDoaYyh8YBsEHw6CuWBP0ZqPzjfL3NMJgAS8OYB0XSYeJ
5xfaJ8e0dL0BOy1X8KRgv1gP/N/mb2jKQm+7i/doh5/M9+cjRjh464R/+DnH
NiTmcIwbtqpifO+wiDwuLelOEzZfwWWj1W7D+9yDDjjDetYWHXSkfv6THJnd
W+iRf3lo3/0qbxjgPayxVDtY5y2AdG3ERJnrutmFTIGYO24B8e9fE6cXzaZ8
+ahmqsmTw02VGRQ29UhkxBkGe1dqnJd24G2DHPj7Hv2dV/f7V6UE51CkQ2KV
7Baj6BVdM6bJIC5jBIe6gbmSL7Zxk1K8aJE9aXFyjWbxt7YPNP2qRu1es0dv
LyNglrcRg5HhVXuzpIIy/mTBF03gZC/XqesojfjwrqPjtNUGV1XkppWn6/lP
kfnuoGK+o+ECUJxQilBoU/GgOlAktweoM/tPSKZ8Jsng14E+P5arLUVi9ZNK
F5E5ad3iCA5M90AG7ZhbIFDSAJtx/cDzFNgqeoBYtxEtsPATP7w1OPK8tGB2
JjHDQAcIQAjekKk++ve7WKe4nf77jWBg4pH5Ry5sn6ZOCh3AsZwmDhK2X8ly
/totVziboEQcW1/vmuuNm/Bfgbd0Ocz6Mjk3BsdNGqHb2G0/sUhD2b6zazHi
GZ3iWV92oGPd6jsDg/OspNmvKTqcN+J+k0cAVHo3TU7/BM+ZFgi4biVVdvwz
tVv8vAkFr5P1SINxUeUPZ7RAVFPP1vN1BEES8FFbLwIXtbf6junXelOJmwsf
fkJzHLgqA1s6tPUFAIQm2FgkLh3fULuTIWoL9mHsgOK+xrb95elR+xjX7G85
oNA+zSfucT6zlZqAmn9bNp9EO06FcEoejvNYuu44Fit9bPPSNskzQkUv9YLq
sKvdOkXM44BstZZsLLP20dUzUwt9f5bWFFnlO7qq9T/l10icBNu9g+Bi3MKv
lIPy3aFtWY4+s3IHviVCknwsnZOpyrHdJkYzaaSZc3tDSBbQ5v0b2lcQNnXs
0uw6WGkAnrdq0vNo1bjo3LM8qMiYoczVgcVelwrIGQjqYsyl/eP0aqKe3TiX
lSNAmOVAVzDtXJdAhWMwkxUuYKlVpYkEllGRJSMMLuSEdBWB6At3zutqF2aR
ks3/lPwgLID+yY9IB0W8zmxEoq1zc8Vy5OAm817IJAAhA60UugdP8MNfLyT/
Kv2cXo7wm9+rKqag9weThLS5WudlScqo7qkTYw97xIlIj3hslR+sucq/bxVe
oJO7b/zDURnTp9PjkIbkuwCsQ2u2nBS6Z/DpbJ9CnkrKW+juNrXANjLmHiML
LsxrouSsiAAVrGxSf7BdEPnwdZ35hYaVU9dYEDgDlQxsbs6hubKIqWxlnyPC
eEBvp67wd/TD1OENQOfR4q4CNFQuicbD/EFe03guZSrOlngjlFb9+Bt2Js7i
veEb/Eh7yW8hlV1gC5slYnO/bTvbV/lAAcGz8Ta6thlblRy0lRoRPzdziqdj
vCao9CCmyyv5YBmzZcn7BAnksAgmSVXdNXeLzVq1Vv5NDjCKlrs38nEBrrsv
FlGZevEewo2BmAHsCNLgCdZXeuXu0u45FIIKuNBs7aWJuYTYXZROD+uQiiMT
yVVzeqwe5min9WwP5zrP/BDyDPDb9VuDIwbJhEwxE3VnTnW35YGIFDnPf9YN
UmYLwiqur/RRU295TV377Vt31Xnxs/jQhMm/orMV7OmPE/cJ2dULECIOklkK
L4mdBtIx6Va6YkM0Q9a17SE0oN/2F3vwUQZC8uDwkVYc3ZlxWo8Vbziv2eg5
SL8jY7kRrur+pDtNrYBFoOE1m1ScjkZlRnumyV0stod8Ej3BfaaLnwCuLl8q
gqD88O19+HhgtOPjKfohyHypv4MQOhspKzEdnL/7atL2z4CAQ5GfutpHwxPy
BkRyb4tJunTY82W+du24j805yhVW8xNgfCHmbk4raSrFXcfb40SGIRg95LRL
dQRehxpLp0q9trxgPSnD/eXL+7qk1kWu+PSyReXrO0G4tfv46l1ys8LJ4oSE
YM9NS39fzg7vNG+9S3rzhFow38qtPViCfBf6s3Rnil4UgHI0ozp0nzTl2TZX
3VEL0s+bGs450jX5YeMBsR6Fmmpl4OBJLuaynma6Fs0gdKuOSf99+F4hs5w2
3bsBpLkl92iZEotOcqXvW0sVhsrxEfiHwZGRGNp5FVxAsBGg6GGRp/Qna8uE
zGf4J+PPRInaf3zZK3PTkHzwade+ZRIToX3Ur0ZfP0jSb/0pMa8+8lJhC0fV
F2hZzHAzVbyiIm4ev7VuutSh1U26Qg3tP4UgKPcBv0stndyzP3rW108VAWJ1
9e8ayfBoXfz1T56hwiSVMd7OmScFuR70mlCHXC0uRlBm1mdGBbZit2FisPsR
81Wv6ue+QBKbfa/sglvaNX6ohrvR7NlUlCkvqHSXFpZngob49KwqTeIeuggD
5WeHNkwDcj1JO33vbs1s2F4N4pI1J2KR29fLEGsDjhekSnPWjrgW+SboYkRB
32WihG1xbszmU3vStH8/StadPTKah6XpJzQj3auIC6qFZHt3do0OjkVTYVFS
u1q2U3ShMfRJyt7J9LbXbBF0IUuowZxA9C0FBO1magFU9ICwZH0qAPENoAS1
oUowCctAglBSaxrNZYyr5eziklxwboFO6d0Aep8/aoow+hhkDbCWjZujiDDt
AuvFMnfdPepHSOef+fgE590X+gvfhXTeRts/rGhn3oN61xlZKBsVYJSTuWnf
zwox/OHYn8xMPv38rZTNzvx3cN1iio8IzZMeNH9muL22gW9a6T1/TaSZGmBM
XZmWvsg8yZgbSG7HNA2PAKlQBNCFgeSRA4mvdgA5oI5dBz8dEhl2Q2/EoMhQ
HvnGLA++MOOWvZ2sN74DVSGu8Bpn2o2PF2rxPLNNrhrDTluGAVEgDqjyrnzo
TbYHFHKAfWAF8ZOAs7yKnNl3I1xrZCkyNaeM8uN4ZpIlMscA8tfNRuYgCwQ9
Y0X7A8/ZbsFaJTITF8+oqRIuvOLNYya3D/c40HHjYLiarszEU16SBUJAOD6E
AjX2GzAvgz1gcevYeuQjk5j7T8dH/qBIU9PXnr3b4f4/9WvJwamv4TkM3d7L
pcjNWC90tNVN5UUjd7bTTjY81YN7R8M2lc+Ypp/WOe9d1Hv7QNDopGXTFGRN
wl648HoySWhrA0tApsR5yZStQau3blcF2Y/x3KWOGAdNevFBwpfTfeiohjz2
Q8G4IKNS7vkcIysUykjPQ+6kE88mXQrP3JKYA21uCgbnLCquWfltEop2mdHm
pRRRgqdpbiKqKjHMbgzFz+G32lOeLfi7KjRSNKnsKM5/uZoMDd7L0cVRvQr5
FsHYCp8aOBbJJjdosnRsULVAM8Gi2yKI5l/T6RnGBYomdLrOygeswMuy7+tg
FIR6qBLmd37YJj+hjhQ4z48taE/uNuy05vtGB08SHi3+ZVRrzxfAYJNzGnAb
U1h0gBEKwO8ybUKMMiHiVKh5V7BDYMxPndf4dFieG24tuUFOslzkMfeiwrqU
ma+s3Y1MhfnkzelMdSIivhfJ/U9rHWSEy/w6HOwY3xbw48CnRzO8Xlo77fzW
mE3iYjhjOrmrjKmrofcuk55r8NJMTEzSqu5Mi5np9vrDhqrsEhQIhoPhBn9e
waaQpSRVkAT4g4MP67I/JwHwM0PUZoCVtmuzhq34+CHHJ9KC3WubKjy091W3
S5ZzqH2GGktTHYFfcgDylmhyMhFzGeTulofVw1QkJ9VOCmqQnc8qv7Tnv6ZW
gHzs0buhWPiDdrBkRVo74I3Q6P7whnY14VlYTqoniUdPUDQhtr+XomgPbyQi
mEOQyx/UwSOOTjlkZYI83BVUvyG6dc48LvHgVDsISbjLgeEPASVr+i3ZLyf9
1losNRtJNCzbWqpX/wPcC+C2s+MqnoZKeXoNVk23BY/DVv/+LR93E1tmvkPY
BPx+6c86Pki0JwX5ems7j8lHjv79/ixAdlIgQxDCcLMlKxPwYYVdeFmtt/wB
L3IV6RjgiZXaZOeKzbNEEB+tFOjj8zZUUTsAiFCy09BJFjYUY2bpLSzM74C9
84DoCJaHmBL5GWxWFQhaeA7iL+GcGh0rVJpN4VgD99rzfHD2iPyl0BtTypDy
6ZZ5tKMdEsFSjFA4d5iucQPzEPlfUx5C2KStxbjOvNhYIDE+ouuDcAJFFvdM
yveiOm6Pe6WnS76BpjYppEnO+uOuGYnBTCTcKxhkk6f8uBJW1Ua3Zxx/+ffL
CnmF30Vv+mvjrKxo/MLy6z516H5OYCAm+F2xpJWeLrYJnwFdVstJDkhVfdCp
+G1pTDuPad3D0wubEGSXneaF/BqzNcT6slwjzYI6yGIz5VpGT8hUZJnBAMay
Iv7qNVDiXlJoFhg4HAhJ5LPjyQzA4BWSVCuOPsippKKQcntU2cKfFehbP7z9
R/Y1+fb4Vc4fGaemNbVuTOQjtm2r3shPZ26CQAySgAHZ5Oik4aiHnV29QeBg
UiwY/IMyPqFZzCe6assYfid/7V0Ga4alWw7Od2kSp9d+BOVACe0yqMGLl2nj
d3AkhYzR5K0SRze59qc9/HHFOpjfsXWbKDgwceJukh5p4bLaaPqVTimHt/Y2
3bdrmaQcupKi1QD7a+zCyDT7o2k2078fryLcolccMs1pBEpH1Sy502nBD03O
w2PxnJkwFAqp5gVSF+EkbZIhrurc0eHnRgLAsMgeBFaKbI40orAscM/fdKYG
lm5O9A1n47ovww8Dv6/SMOTREm9iu5aQgVlkz/NMscVNjgMMFJfvu/OVxtI/
TMnuMiqm4xKAC8wBW9Ut0OG3raEEuealYbhPywaFEcHLIXqde+xBAkJr0YBn
wCVPh7KpNpYa2KpjJAC4dfdxl6fdNbuSL2a2xwMf55QjqaF4kcRnkPczVPwN
Wjqou5SnkwaYOXQZBsGEXkzEH3sUdPo0LZPaJBUXvYfZYV24xosTgVmzTwJa
oe3nK7q8u4u3vC/2E304zQdr3T7DDHmxYlBveK2spMOfmcpskLLoB+L8JEo6
DvId1TEbaqbp6FmOtS8TY9y0WvCQT0P/UsV6u9APzhtx4MSOIzaXiLUxUK/Z
mvisD4TKh4HmesuHxCHlagFn8ihjmZqstR2kGvCtYwR9OHPCLUYAe6JJADH0
spT0kuaOeOCOsRAq8xn1nsNaZsdFQsWwXqECyJhmc5PlEXp2SVqPp2ZkAJd+
eNDDdUfFidx86lwp8VhpwB/uxlOtW5cP/YI+g6kk6lUcJz6wN7ZF7qS7dmuM
ksW0xbhJwRtIJ6d9fOWq6qO7KxcmjL3lExhk7ivX4scnTqmkSYbygDObRNvN
9ltaUx1V+yNNpBvcjtvnaFwjDi+thTvEewUCJzPqKXECUtb/fia99/YPh+hK
++NP/eXcCREMKVEsD+U5fwo7TPPKPyJc/KuS3LveUSl+gQJ88kNU7MTScXtv
nprTwFoD8iT07cy8sZ05PEVSZWFMkQDEwPC5A9PHsjt8owauI5Cgx9Hme/bE
+5qd/AOCODLe+OwnUO3Vqw8wQG3cd0A49Dt8JKLLaujKOx9RhWhpI1J8KXgD
fzOTGq5nCLhNH9cEUgAcZy7DCFy64hqsndwtbjI3xCAN3RwiH/Rh93SLypLf
6dYEPnECkOxsyiY9UfjfkwB32YqP6PJg23TB6lDeC3wK0fToIhS94GAZQNmD
TkGWOM7tPhBqQB76jeYC8sC6XwWVcVrf4C/y6lTNvEB5KlFuNiUy3I4er2GY
uUwgJBeVuTjTEId6wUf6pAZdwsFtbN+/bfX+spLz58hi0R7m/HVTzAtRo03r
5Ag5G3HlCDMB+MeQLeijRIk3pCrKYaL90nXWfnnu5U3Z7dgLVuGSxyXR36uE
wrApB5YzgmF+7yuAh/S9T+SSUEsVsEK2cDeZ5HcuI1n2oe43+z3iPcI3tEi+
n/3B5Xo3AutWZv20xoLYVZ3gnqAZuPijdmutVrOH2/xVm1m/asLEe6sd6NOw
kogkpzL0WdSL4+MHWXuQxicuJzSnpjCXruhj8QnwP1VXlsN0DdYFreXE0+zp
MC2F8MBXeiR7exxvCl+bzAy1l1cAcmKvfARmT6ScuDZ0Tjw8RL3koN7ABPG8
fBT/OWstnjsB2SDMmpYy64qRkA3j7ube2ea3GKqZLOur5FFP5LZG+Gtq7FIw
/M7xxQqn4Y7gKNPskqQTdhStrjNIZIcucVbjKxLEX4ZAOFKqubf9Ef/WWGSZ
jalAELpGOJ461bNzE8soQQDUgCbPI8aP6aNzt+miKKURkAcEirVoXxOXxsQJ
fMmHYIsL/SCn9A3rCFudTYBpsUWt+BhJHSkAmDaFZTDebxceJT8Lsh2XQ8kq
7BRXEiqjuA+bhsHKXgwE+YUSRWC7ur40zMo0t9Lis3Z8AkpMvymc170rcWTK
xay5G+SWSt4VkpjETpbtqdWYTc9p8Urs62tl9/fDOI8PLmSS2OiNGVDZx5Nm
Oi91Jumh6Gc2EhmbrcBwRnPoe4TBL8SODJtJ1JGNGPImcdOeYvNYVKU7AqYg
Nph4gVcXYWYD+vUSWBMbwVtAiXVIaUGZvEek9jXTJk6IfDuki3H0Y8hSadNH
wvs1ByziySCuPd9CjUlbLKBuR/xC1d4PQcst/82HOQaQUzukyZt5jK0xRUot
eDB2Kjk1ffCIDQnJMg2QDUm9yWkVXAQaWW/6L8pQkBU1uHjlZ00KFrjDH1q5
TivdCxCWv+e44QYtOVsJzS7cbOIOi2WMtpGmQtX4abjqp5+xJOPr9geadcK5
w17jwi1Pcw9TIL5pU3soYbB7fKddNM+5G6ZjD8amaRj/6QmxOcNEnZNl15Fs
qSs491Pt9HXgue4ja7oO8GpaH0JCUGjcFkgJSxbA9v90Q8e6kNrTMtn6i5Md
ieZGZF5jEDoCXqBq4+P7MSM/PuRXvO5j4AjlL+UG15BRLTlW9eQPgFpv8ta+
2yhECXl9n2MKSSBPoaE1xjBbq5QN81UFUoLVLEq8ADtODM3shxnmQdbe/ZbE
idkwol1JW5QVro9UqQ/32gDTc/Z/q+8QHnjYrZPK5wGK+KpejT4fUzyMOFFI
yAm0ne3l6NCWNemapcEgkZqQQzN1upv1iufMsbTOxuj06PDXJxnCK+xT54iO
c9+UemG3LriTAFo+tRWAMoaiH4Z5ReaxNQb6Nf7zKJINxV6jPBgbmQBnbiRE
wqMA3jiebGMPwlt4dmd1PTzqGO9L2oci/7prEOreg56HQHLurhIq5Rd7wA67
Cw1KWoVaKLgUB/xEJwNPls1L6muixuTMiBEmAB1MbZBoLVpMiOXigliQVaTo
ZZcxfoNS90kfo0c9Jw/Kc0fSt0cvchIg+yfs0/O/YVAHcaHFe9kYTR1BoK3R
hB9zwheuPrrZSExfZHbWQFBhswWPm2ikrRMrWl+I/AMc/ZbSCwySSPsqaUd6
0XdD3AV5skDNtLHExsg5BFiTV44/g005WGuvZcakCg30GoqnevljemtdZSIL
onSE1JT2otq/X59zVyyDwDHKhOgvkjzfzNjd2PR047/olFeeFwN3llUZGLbp
KPBg4pLkqRXi6B8epzdaj8Od+ejsAYxwle6WOuwAP3E63FzMs3cQNR+MZb7N
aW6IaR7CTEDt8BJKsURPNAq6tsGBJxByQjearEQP1Nlp23EdOysCLbmhAoLe
u54iN0hj/GKBgCiOXXtrtUjSNpAbb+kAsrTag0cdP176KDSBj3ZuVtssPvc+
VAAkgG7Yj182vdqqHK84rM4y6B0K9+EABOcYKoepUPxL0wmksG91a+UUjGzm
JvEGe5u3N3TIE90YGmbw5fhbEswhTWacYNPDC7l7A6+TD170QXH7CTGqNpKb
tiihRlq4qNMYRAvpYkeJXF+8OJFtpXxLeDjxxXR+hG4dgihfPc3q132IfBvW
DUWboPScG05wakDBI27lqkXvAzGgJPYWoYAn1oyaMv8COvkmeUv1ShjfbKap
n6BGFCTL4qfcK1fHuqCo6sS4TBmVXwGLAGdxVUbSMlPYm/FCdPTNwfbjnxhM
yziXU1H2UN/t0ZjS/u7NOJLvGfTf//OJqMQJcyDxAfGrNXO//onOxPgRQKJi
b3lULZY7NF5V3ZFkVx1TJlnxIJ0qGi+UiIC8s4f7oG+lm4BZfFz2HcG2zjQS
ZrA+Mu7mcDJnuC756mKJhguGYq3U5ojAztqo3w6vlLTZZE0gyv8wEl+Oq09m
XukU4erIZcUKkPrDBBI9KwMdQDrC7bBPloZI2PQro2NXWKwFjcgmY66G9xUl
zjFMbK7DmA6s9U4h2wJymwtjhmDcOqC9J2VwpTKz6YAesSrXbcfz5V1iBRoj
rK2EWvRHphgPP/GXOED3QbToJ8rc1ShLwqHt0CnY9dKO72mzX4kgyL+Ef3FQ
NrzhLAZE4HwrRHfH9+F63uph7VoNxCLYzZULhc0wJXjvjgp5kVE4P8Zrqk7X
Nve1mVpaSuVry0LR99ovkmIsDY7sWMrHr7WpNQlJCEGJBU/j2SwDwqqHjxsK
BE7dec6q6ahUtUhx7YMTrYRFGuwSHulqx2PxU0PK1873FxOrA2/fBpdfKQyA
tjI+OFaB1mQqKkUp4CIc1LwORYC1/sELUvI+ykQUvBJRAtpMa/2dwCmBVWg/
Emg/5kBsuTG5AgwN5aDdf8IFtCjuutnzVeTtKUorPHtFQEhOANvLt46sBkCh
AflViY47Gun+/69Avb3jQRUki0U6J7yDukX2qirCIhe4XiMgw7jdyLWQIupS
xBr2A61HujSb5AcqcDmUsygUgQqvk7Xl3CHUfZBkm4SJbs2hpGnlgPhOWea7
08xgHJtlZ9KuCTFgJpUTStvyCekbEYXsiK1rbgrAuXV5CKG/5WY9B5rP9iGE
PWL2YpCVXMyb6XBbI0943JrQKKJ+RK+wj7wZ5977lkER7Y/MD/zzqBSJZI2k
vBgqnVjuBu1gqmFGfdQ7JFlu2s9spoX7d3tkUiGOtRNa4GVyDNVgzR02PhdG
ZpLN5GAKksIxRBmVoJ2qqWfZH8S8e3PR2cszgFWS9H79dQGBA2+OcZqSbHED
0tsLOOEBRp+eKZ6OcWkHG+mOUx6M8lpuXLTUNMje7bU7ZMpcEhzSU3RGKNeK
e95xzdcPP1wZIZTM/znY1OTHwDonrtedfqKw+jcgJtHewqLTDMbdEYkkhf+9
MHV3oVPz8+TV7iQK82bVmX6fAwgDvgk+VoSdT4iRUC6YSoHXVWITK6JtVfiJ
nkhPB8vmu+cdFR3oepKKigQfqQl0qClY+dKboXIXsMkNUkMAxH/yS6gKDVrx
312TKF72v5epTq+d8NAmhB+BGkRQI22dyyHqg9jC+Qg5/0Lo9dfnRoIxUBQ1
2NscvtCtuEu2lRCzB3NZdVenXgXVZKpR9aAH74QCZfxnMXYJjf6ZNJFFtvBV
bBWfMoDpBcyNiht0wbCICrbauP8Hvwm/Gswpuzz5rq73ZLQ+Yvz+a7Ivy5d1
BUkRrCFl7rMonC4xQIaex3ktiMnHlK78ljqLYkEOcAHEWNKbSN+0uM0pgVsv
KhjehV7i4t9FHrEfzu+NFkR7FGUCNjWkvwKd3YD/tSnP4YJkxIl5Y7p7kcrs
//pGaWUL9La9OB66d3MQ5HfG0Pa09/LI6twiBIqLruW9+tZSSTKtFdipIFRA
6ifqH2fwlJVmXOlZmHcbJHh9DOq6ONjWCH1jWhjhR2tHnpD7izEd4VaXuxEn
qMFCr+hPKbZ/SgZEXO6Xi26Tk7Tcs4TBIPTY/H3FcjU3XWLo1GbwdrNslhCm
Y6pA33/xMq3H32SFFG4xhXP40c8yICRaDuntKWURNrXdm4Popn4obfhh7xsF
L1noQABEh+FX7JSyTtaFmsBdZzEWj00aqjXbLVlOSwslw+Ve+MBQ5mAExd6A
BAudLjlmF4mt+M497iPrLXV2yYouMHnviIyIZuuYTfPNMnYbXJ0J5I6JBqD4
10TLvk9SOLRjwIrdt/4d+WiD4+CqoCZNzSGlvO919bd3Z/4T0sbh3SpS/7io
8Yz2d5xG2aVp6yCX0ei0LTv06flmhEsg1pIIYyLTZzoC/qqTiYVpMDhVpsLq
5pgJcBfNt2SJDXrM7+1d88+H6MfgRjYeoiJIueFZ0zBrJMPvrO2SO0x7ux5H
UHT9ViKlBF60bs5jcC0+euBfFuxCLOyPo9n6t6v8Fdlg3LNg6drxREykj6uP
V6n80lUpbcXvbJHlicBm9ZZaLOR2dbwcRr1li4sCimUi4dBhB+LrRFXAiOE2
3JX5gCsWkWmtWlMS1f+gCnZqhkhIX7p+AYGpIDnWUTkWoaswvupHBlbeasL3
2qbVUgKkFwMQBmXOfeG8Ai/AzyZzJ7CAVa08kJjuQcbmuDWzEFLyeSZhXuAd
kYaaRHpJxMoqi2ZLn+aG3OXyBfakz4qQG/yj2HoSxmCTKnAo/xh3zvADtOA7
t1C62F8TKzX/0/+OGQz8bo/7MiNNgEmenUEF5CU9mHgwg13mFBRzeZ2G3o07
GYwoc1VUuGOlEzgN+YcaS4/FwtF7jZQHhgjtp4S33hymIKyrsrlpkWJ2U/c+
EwXJ3pgj/eRoZxGn1kRGd6EOHk0289jGUbnCDWqwmSP+JR2to7AyVhyxY57K
gvOnSmhqGvYIB3al/lUCeA0IDljY+jZ4L5vVMh/9OPGE4Kv7o0kR+oleQ79t
H5LbKPeOFn9HGwSqxHfVnWvJ7ztLBde/uepzEXAM1sRGKPXG2N820LJRV+B8
cukuZC5sevAqpGArJF1h2sypXdlB+NDJc/5FzxIKkNGHtGoI3x+/U9OVodWq
xAG5/H9/gTGfdYBqdYMuLkqIgbtvlfGv918aswowa8HBqDG3ng740ZyETClb
rmRni48HlCmsMeJeX8iomFhHejq3scdG+ZC0Eiw/Tw3Z39q0ZwIhQ/BkdrSh
jwSMI/amP20oY9OCTydEDbnISwwch+KA5jGgjqDZDCpPdbOdLvkZpqnzEwCc
+kOYfK/ur630i/KeCz4pVd7RiZ5kkSLvFH3d/Y+L7zd6T9Cbvp88sIM3srnr
lnhFS2oWoZytJmGpOMP7K5MBm1z0ept99Hh9qOMfquXb/gDi/uxOSqtlCBBr
5kER5hz2F6YXTmfnb0OwUOo8rAyj9T7sogGAW/fUqan11vz/u8r2h42CfFyG
6uI/RO8aq00OJz2n/k8ECmyMguO+dHoErlGC9Y28r5OMWZyyJp3chPJ0KMIk
U/YXjkyR+DvEwiEng4uPgCbnL7ZCjaN1PDrGLh0Da4QsJgAolwRRmwOXiLkb
G0bcjQL4sqYHuKXPHIsvsiv/NOjfRYZrFvSsyKud1Y2ZTPkmP3L2bKjrLASi
mral8pmXiPMawTLKdHRc2xZRnEVjWb+gYXZpzBfiiwsmTL8J0429qLD1LP6F
SAbaUMILTo/IZywDM+2y9rPiYDZNjAzZQ8TNKEicg9Z/ryN+8bu47TxJ9rJt
GJ5fe/pDq8M1XBOFqPDMYpY92mRKbs8hBt/t7bEkgZ6oxDIMpP/Pd+WysKPz
7I9Z7XdArr7BHurdC+fKxJVjNk99nETP4NupnTEhuAh7TtSGDpvYkXeGEU1X
jpGaSXKcErx+hCttK+C3J8ov5kYX0I5339VXPGEM1r9hLhmmik9qamIWNSww
AHfRKo7SL1e1Z7ZAhb6TGlebozFAA4CFGEoMzzExMhz5vAamqrUXyxyjZshm
Ng3gnIK242jiKhQYCel73wl53+zY2hxMupxhWT1hfa73bnO9HQWHpZyWekmq
nqp+GcqR0AvA4MuQ7OcGBiJqWF4Dm0AsiA9DrovGNrgz37zujtbLlUUV/q3O
/OO8Ff3PttG28lvsAjo+zyYLFei2kiv6mMiwfKf7PWkuvuFDDYCkACYoDDWW
i1uQRqJ8SC9EVKZf4fX9fTcXjtJsBPJWSfRhM7WZ6U2cuEKawuY5O036Hkjr
U9IiCgjtHDFAdeBI+GkfnYbY89KOQ5fXQT3goYiV2BdCwKGIDxzMUUzjqPlw
iO/+wL2dBlfMgl9T8bm2HNr6QNBT1fZSOrLieOnQEG0OWDJRlf4Annyr6cdQ
ga1YL9kD3RNlNL1bkj9JoXTDmD9Df9r3RF9tJQkionwTtlkxEy93QU2NOBK1
6Ixt6mhZ1N3+a9oD5PxfAm06qGV2TURZG6Prjc1AuD3GYvQqhpSmRcrt1Tk4
t1gMFediCdr/bUl5KWwWthc488MM5+i2B0wIoggpLCCLdd3QkoqPuOLaQYTw
X/Otetg6cIlu2+brY1x+Z1MgbZSNwWTPFVmRnpIbz7cEJgtCTplJmQxCHNuy
B09cmJ5SxIGme+B9fQ1fWlA0DNx9UxLex6KBOT83pME5qkfryauSIg9zxPDm
ty7PP5KllyI9QJDdsRW8RSWEh5lX/Z/98s1jo2yu924N2aIWeiAE6nrAo2/e
r0J4BvZ0nnuwlhF6TjYZA1474uwrE2Rd02aI68Ukf8jItUw2lrF4ZtIa1Rbm
3YKvtBJpRmEagVVNj3xjEgXKhDrtUFEjqlPwALexrzBJxxzZRSQuRmAsofNy
UwixXyNOmjhJnxvVhj5w2YpmMg87qjavHq/e6cTN6HoYSTemfgtu8MA0xgIm
RMrwH2gej2plTkk/eTOckFW8GkRkmF/dUpTqeSLCeINSqhgcd0SVlvUpOVFp
Fp+zbt1cjEG0TjPoExvr7JV3LrIljGHX6IA9RWYcEkF0qL9gd2jQdRZQ6NQm
PH5mNhblWkRqQDGwLIm19VBVCAOnGjaVGFDD4f/8j335aoRx4uGyZCYJvXV+
FOe4kSsqCM76+pNzv405tK5VWOYcygOia2lndycIBYfjEmQBdA9tCM6ZiYeT
XtTQDIRiCvJds8QgKx/cokgtJw0kB53C5rblJJFeLqJQHWq+6pCpisbEDoNo
V0qPJkpWaqrp0p7+Tr/NCr+4i8hHa1Eu+pl47K1uZnT4tAR5DkJgaK74aged
xy+e8ThkP9cHb0ZtKiWQ6cG1oT55oeivawvTsS8qgxoiatT4kzPu0euhdkha
KixwHArSHmEShYOPY5tStB/lr2ClLt0rat+K3Y2rMwW4zdtA5nqMUt3mYAet
Wjrf7EXh5S9VS5XGB+q+gmeYzu/1j8rI1t3NIwK3DMbgNgQFcMh/xyRgUl1I
q6ZS6N8H7UWgnyKeOiV74H6LIYHr4sPPgpGncd9eg7IdBDMfaCCZVwOMVzqd
pYawP8OVIVv3JfdryC2T8RCXeiHb/7AUZT8+cbTr4bZeyWVZp2/mv2Bz6Djo
o0BoXuxx5E8NNhzia5fIlzj+oW0xR53VgdWburaaaSOnhd/zwfFifcCrTnPV
dpM+uw9kKJ6nM2qUDzUYKxcvEFQ1ASoI2UYdTr5zsD8mTWqUlwezCUxCZJ9S
OLiylhgi7lGd96bIjormLuagJhdPKejdGbQJQH6LNlkJDtbeVLqxR+cIrZ5t
hkF1adJzgMXFgI9jmBl/QuRXxcBc8P+jcaK1z0pQu9yzftIuyLk5yNQ/iVVx
1C4uAzpc1pdtsIB9Q2MsPw0QrwGmX55ItTmXVj52tlCnwaQCqT4GFa1c3NcG
nhJH4tq94PI5x916JsBZKs8TRI76tfMOknf7xsRiQROtAj3/AX8X3NWp6aQ8
d7gTpd/ItsViQ9kXm2fchBSgFdrx5a15b4/r4/XkG7BNYQyhnvKE8UFpoKrh
E03zlUwY2fpkDfMXSYUdJCYHcwrF61PlOHa5CQGHDBYKaH0xcxdwIzhdeL9x
zw8WarMkaQ8RzeMgWJ1o1ToI2GenzsJVepdjAhN+h4duZavmcjjZI4AI+CZZ
B/aT+BZM+K3ET6/gLCH+qvozmd/Vy8TEPOaGnLOWd+shvMqMZUb2yqNPI7rB
UVBIXxc4iXhe23H/FoO1uhGVyszFuVdVp36OLR/ho1weJEdOyY1Oa70lxeFg
Uy+TlicELkaJWC2UUyZh2Tj9zGVjHDJBkmskKY0rlf4NlERCteALWTCLIejt
kRiUClx4gd7iW8xG/SPVxnjT1snTzJdgiRBSWA8K32o7qQi/MRKbAHYFgbYT
V6fWyqc7wWfbENAi2cIy4GPh858l/XKtAqTi/SmCjmjKELtop7X+DX7A+piS
ogssu3pnxO/H002Eu64wE4b1Q40Rtb0U7G+TylZvZwCcCITJcYSplTEokvsl
VgrnX6+MXdzOFdRnKjEcn212DNe422lzAbtNSNGrKbitvyudtoijCeASkWR8
3Qx5sY1H9+3qK5rG4/aNH7oC4mTJoBQG/hLUxGppUHujegHG05t9feHROdtJ
0Icm+mVOKkozy9zelmwCN1/af8x7kljTiH9ZCHoDLvYYIpswnWhpgHq57wOG
UQLDve2TxaDAoASG77pwIx9HEyzSuTOyvNuPfLZtrKdLuCkXnk4NPHkN2n3Z
babjs/lCUPSPNV5caKIkB79ncT41jOjc+W2hqNyCl83fI9rOxaPW6nS76h1O
RP8Cqp20IBVnyM/xB6VMWzFFeIYDEur3n/gVuuVuY5U8IMMReNBFWXj7eBlK
fZ+BSryHGKNQ5N9IdbWfWx0/T/wvBBHzhgC9poolRYF9wqT8BbCvkM4Vp1Gn
3dOUSYDjim2H+flx8TD/CJo6Jx3vcXHppDmP0DjcxzY0Tx9T3gE3g5febZdl
m9zlwsFUQDg+wFXl4nsWb1QupoTQryS4T6hY4md1i1KsImx/mTY05u0alAAu
5PTioJj3wvm37+ThdlVTlDHWYYCqaM5z3uo0d9ZzjXN8bii0Kr+9J1alBFhl
kAnzVX5tdRdymriK9Kp/Hq6T7FPfvdgJucTEcpr6WTa0CZ5EngEq9ld1mLoi
rQBchHYMITbbIoF+FswzIJIoybOeOgGmOOVg5MJck/fHK/r1L7oHZ5zvhgTJ
lYKVoyFfG6b5uSBcrAOSV5br84CYGjBsM2iP3+G1bNQCC0AW+ozqOEdByMHs
xDhaAoeawOfNjWsuGfOA8uD37pJPpYLsqzMi3k5kRlKuVKu9Pu4oZXOBEjRU
gYhnkl/RUxETJsrpJJ7CjZhfKyCUClowJAYq2lv4PoJsV21emTZyRsctTZJZ
E9lKeNL07uIkDQN7vhA+hTcaKVFEYcBk4PCogeMWNV6csfzJTuIsBrrquH1P
pZ6EwVxJncYPmn06Gw6A7s9Cp1gyDlGMMIkGgzG5iBwvLhKUCvDfukR9e9Xv
svhdjjBbC34iQH8nA6P2ISbxTuoxiLpFXOC2ny0suI3p5v6BTZHOsvVudSgc
Up78r5kbm/zqBcIXpSbepilZXcB5Gf4pcq8BStP7/eICxIqduSx4WeYDXDLv
Gd0Xoou7AkPKymhgIxm1uq6xQRiL5qHKaf+nnTzXNMX3hz3qehpUfpt/RTtu
zWJ/ZViKnybY8xGOsjIUZCqYO0aE71ZgUF0XXvRMsQ7xaJXKrPaBGlp24Udz
bq/+YHQZjq3zrXp5iqTn+ok60K6XdGTVm+pv8WmI4gCXFX1A2g23OBEZsTe2
KlQ4ZDSXELXfFgGuNyaCnvgKvbnY6Fcu7o3G+ed8wle+YadMopc1wVZJKGGw
NtNiMQJ9c8vWqoNpiX7gUrs3X/eLO38a66CPcmSXldbWHNravn3axiuDmcZQ
OLEjdR3ZEgo+fF3JqiKkvAQ6yck+IEI4bzclHqT82vb9U0Nh9P9lk2HTPacT
a/60tvVti2AJEygpHX3qHMPlCTkA42d+oNVYpeKVQQ95rZqX8RKjy1+jtfTF
zXW6QGGazw/0U/KffpTJT8lu9NaQCYKAx5NMvQaR+lY9aWoK2UayW8YoU+cw
1cqLHaM5NzDgkWCt7/s/LEGEh5xFJx5swGi4jDIcIjWE9eMm3/U+G+yuE4yA
ssL7h99q646yXk62G7GaGeu8sGwdRRxX7DQFHodIYhOhyXNIQRPv9SB8dttj
g6CZRW0wIRh4TLk48i3HRpE/KMk2Oym8d8LQ87du7jChXNcfEiiShufJvWCz
yzsXDRn8UUM/bPsZ9Q6QLkgT4/r3BX3LKWnxwz17zj1dcL8td3gMbICnfno6
AEjMxtbwShZOIRidGOuO7eBjf1lgOviAk+8xokGUoeWkzUMdOx+7oUoEFRvw
hWlTHH1CEvKpy4mG8YKk8wnABiIEMQ+2h07bJKlqRXvXV5bB6cmP3i//GlGn
VREE/DvccnUWLodpvon6FrtrQ6RzkAk+HrUCU5BY7VAQ1xK7WigZGg2dFZm9
SHYtyIey2vypMV0EGDCg2NjedhFro4tHkaKWtBMhYLBQYunPHUc0kLSnt45P
aBF01sXmv6mVT49q2o3v3PySKo37SlXhj8TVvEEgemDfuA/GScSEedr6HXv8
QHENW+MyaxRjQkf7WdZB50772WqOhmvEAHjEhQElSX8U5g8EryHnyMLBvpv7
YiBhUjDeeXWc253bi1nIVs8hEkUdOCJ1tTHWwNZt73uOMUjzpmFa2LShcDjG
2ylbBnF5vA5z2kdUGBEvxVC8muc1dC3JEMLaczIRstgxoRlXJLNLfvUmHLt1
D3AqwBh/Fs3nRvOJuPfKMQdgGlwpbTFt20/UROKlhLVfAExm5GxRskAXx2Mx
9g+H6+PpGpdBDlm80ctW36aqWlhRTPx15Bwg0wRRi3SK684HQK0+g8+kd/aQ
8mVHEErYUjmXMjFswex+CmBI9REKBxUzcVPdpv03cdqUXjZ4+fj7afpdbIzN
cDVBTOfGh5HpERoc93OLKxqEConZNrSZe7+5DQQE7QB0BD1EQ8nbQDfyK6AW
4Ii2+w4x4CLrNuQvHAwMgBlBecnWXB+XVmpk73Fa0OA4JlPvr5wWtJV84ZSI
8FiJYsJX5HRkVQgHlQVRMcPYTuN64oRNHt1Vsi+MzJYCRlGVUWnOI/HbWLV0
gkbDOoX2XrEh7keE81XIyN5rdMWJbO4XSVwWsg3bztaxEzgWNgJEjyb9N8/u
MX+p5ThvRFcpSFt6iN5iCQ0JyFK7JN/cppekGat7c2K3O0edVxIEUKE+BCcM
X8vo0QOdySf6I9BQ5SFcTPumNQ4RKbGPtwWeQZOXikDKjcwpmfxb57rOCM88
P4anW8UdSh90bba53mtOoLA4VJD5FejKk8yTJoPnYeIfFQgMxHFW95QzsYuR
2eMVnyYNqo/chJnQGovCqepXCOaDUg59kAn7Kf9888R8TGZU2dDjmiw90x0A
YUGV0fj6bPkXGCnENT1Pog1tY1Zvd+0Me4/TeVeS4SXrSoBTcZXAhDR9gT9x
DQyYiMzEaD/PIkrTso+Xkg9bmL//r2WrtxlyrLPkhhEAlwrhFwkwWa83ZcGq
rigabB4BMWJZFQtVeqjB/ewNCsQygHJKp1FPQMS9r+wX1JVsdIZHaBG5fWrq
pXicztbTqnOTls+Ksyof8v7OdpBuz1qze7Pwd2JvR1h8MHUghSy1duV+8bhF
KIOUi3SB0m2fa7jemBYyza5a99dGYgrGxe1ijImwuoFwY4pxlDeC1g9dyE6Z
pRJyyrkXR4cDM8JwkVFXsbEI+AzZYKE7BWtxDpqu+j05JGgXxVmBBl1sIrGV
fH1sDhQDFdsNJgD+OZ+61MmUFm1nBIJkF3bST4m7wtCY/BDVlCbFIKWdz9fN
Mc21gqgmkEc9W7xipcgeGZtcsVfWFZ0X659VNsHyKwJySik1iV76YFxQXOK6
L9aTXhQLUG4qMvm/7iPec/CG8Rzu8FmP26ZsShvgutWsaKvMJxvznkt255by
WFw7puV2A8LlHEYlpTtkV/e8G+5WqXCHgJ7i385Ft6oYrp4xtumzrF5cx70L
UxrnVBj2sAiC5m9rXjzinwdiAFCXJvM6Rj8Kcv3emaUCV+vQYyHZHsd974S2
1Y2tAY4FoEuAw3CJAzPCnBNaOYc5NNx+JFt17jAs2PBjzR7b2zbSDwvZOtbe
BtBKysTX+de2XxbU5A9jQ0ffYmCDKoPEb/2PG3VRKqnMIJzRuOd/XREJoJgb
QAsEGarxHHvl+aWBkY3pr7tVuHvR4wpTWePmOSepS1zCjwdBX9xBF9ahdV0C
s6atAN9RxYC4ky8i09yuWO7XpjP7Lxe6EU9GKssZ7eYx7/GJU7Y8YJsKDklO
QuG6Ng64VBH02pzBHl4gWInH2lvvehQZVb+Ql255fjS2s4JIhwDaAUJ5eDie
cZ1zTwydXZNaWlKy/Q92HAfSw6PXFEdSlgHbhBqIcPHI5KbgqkC/45v//WTf
+ah1uQ/Jd+A0nhVDG2RjVWh2XWeG1gUEbiIB85eRmig1/D0QC48jyDVGzldB
XY0X/+VV8HBE/RnE9o3/3k31g8aWbLqwCJm/tFXz96LFx64wSkbaex1tCqZT
Y9mQJkYEhxL9z18mIS0F8UuZ0gRaKZypD9k+Eb49XWmI0ZGMw1STZxyy3YU7
cRYcYvRKMC3vjVGO7vguIPaqnI1KTwLrOfxCM3e+MpSU9Kbj4bhNVfeE8ywS
lHZwGgl7QxIOS3v6+kqpXLu3vloo8EkSGpRl267UDJLMpemajx6ozFBcDxUt
KWECJqIw/nmjlFruv2LblMHQzUJS9sh8joyyyTH7AcuGrtDN1G6J4AWBK3ND
NGj0H7zRaqtob/p/cav0PVz27o4UHkrwP3289U21eFrIPvkF1CIxggqCT9wp
vbbHFGryKKJKqk9YgrYT8cRcq16i/8WGgJrIQFCCDVfeIoPJ1S58pLY5lSuY
ELoFh1M8N5jWK6Q85Q5sZ67DrUzD4Wh+VNuzzlON4WzIn8mEWy4F65FGzLxa
9g+d2j586ANG2uGATGF4ECZF305QpsSbpZTu7Zu8/Mr97zKS+P343xBP+VDI
Eb/7OrGyWD+uKHnIxGI8vPnnOJ68GbnNK7N3Wk5CxotEZ22KpYvhPHvh1Y/b
hd8J7n7iEqzZmXGcnRu7Q0U5DXv51/3mYvJM0SBRA8zRa590YxUVv9LO3tSr
+7lhdrfvJWiEwla3Lcz20b+Aw7Tkwbs/QIwQ+x0mOLUZQDnonzV42vDe1Kyz
k1swULebhsqQviFrZ8EZYC6WooBGVQvGTC9ax/hf6rC4I7vrbTgMxwt9yWIf
X0Av9PvbrBaw10jRikOYqRoWBnnJlZmIiuQuhtiba8TOZN5s5SkfBvLaKXTr
Hqn9wGDrTHT6LpX2CJZFmaCHIYixua5OOeSMHuQ4RQX/qyTPjr8enCIrGD83
hhJrpc8wL+rXmCuAzUgHot1i0HRhgtRQTeU9cXQQXp/PxdgbLSAahjWxaOqD
Pii99JB5AGx6fHOMg8FwHoVzjqrVsjXlJMCuMbISLYSeZeN2w/5Wc9DtTVSf
KLsk6BNpjiYC1ixJcuN90PTKnJLKQthRTGMQPifbKKf/QMQpxkYLezmNXu7d
9i1TMyB3PVLb5LYjnHYeYzm5hIuHGqv7/Lgo3h+IP8BovzowCzlg5fEmJ2I2
zORvaw2HTOjTfUDL9P58/IEz8x/8JLVhbXFexK9Xy8uHXs2w/NBm1TPV9BoH
wEz0t7GZb4hOdcMwPpITmdWFB4x5vf3Y6gOc3zQn1U9Nnu7KUjIA72rRFTw1
uVuH5inaDnA9RnUL31XtakF2pWSKm9AIvPs8AaURZ3D9eGa7KZOYZ7+7yBKg
yD4G/8bR2dM8i2YdU9Gx863xDeslQC2MYtiM2ZjxT1ELKvtcE4KfClcHlbCN
is3CUDY9mxP9MFa3hCNIUHfgJ2zezaKZZjBEvs4K7Yveqkz4JrXExMSjza/n
SWlTv7Wox2DWYK15D/cJxu8AnJujln2XMdlg0JzUNSLMr/9PahmmkCyrfDcs
i2fVpAlN2pIlR/CazRGEpddJQ0vuo5d78Aa6pYraKhDJLC0mE0Bd3ri2MFIS
SxZMQWTQYNa9CzMS1wlPJDoKkGrhSupkQ2fps4DuFTBkBAigmOqumKbNbC++
y3qepesXz+wVDcihTVEAt8YScdYc5UMYXc6Qm4ipIfeWc6dJ0q3N1bwjgX8J
P+8TMNnVl9YlMxd8qjSt6onSV36fkgWa13piSZBxUnpyBpqd6R2sZeZIQMgv
nY5B+6DI4c9J4xXD5mpmO87Ks+M7+wVGWOmUbXXW3Q6PGkGkCzT1rTKKEGJE
pccZ5cAU57aR1inp1C4MOvYCg/hE34nWOICri2C0F6IltM5vIGb1SjnFTEr4
9mGXGsLYA8kT3f+OLkwNeLeyi1XNUfctVCgbs8LA2eAxSGqbOwflWyzck0xg
x7WAcnAxTcCGcuCMnZDaYEd+iRqHsC4b2KzTKRtS6FuPYiswqjsv4kiCc+qZ
3l3h1dc3UP/FnghMljUP5GjeqtujT1w/JF77VP058CX2pvK/pHNiDXCabBOV
SFzPMGN9yAs2SD+UT/Z+TBB5vbObxhZT8VYYcjJ3PyBaIf9x3a2awirBkj4J
Ymg2JQEVTuS2/n2hsbcH/pfy3q76UcQrjqpr4SX77cnPX8q+8+hykxwCeiKv
/+rhsfKctVshcv1SxDWnzfV3KSCQuwgRUGg4KsaKvcZYIEqIz50rFmbtxC6O
rjPomoVia5Amjl2lUmuzHHXCRaiironF8fth5mteyJiPM7bFT79Pf8ZRiqyp
hFsf0/5SWL5Dn+9EA3JTzJOtT6+grWqEe1HGSE62V4bDirrQHSg/8/vHTUd5
stMqW95uA2j7fNoc11SgHrrs27BNXyYMhZeqxpPivf1xVz3nkki6tLfPWNj5
5f5OdBr+cXsAeuzjSDZ+nGIo0XerhXskOD+0fdBEERRMO+rhcm4k1ql5Vx5+
UZyLnIwcKYSzcxXXjFJLjBqlZc5aKp58tqj3QtuGiMAa+EALwPN5/gjz97PI
FNXf9gpjnIQOQ9ASFOxYWMIyaYcIzAH+gcwVhmBhmfHpvjNr7NtjMkNv9puM
+RHNGY8CPkMPPEotYxhQ6id+8IUHzTL9SbLfzFNxlAJ3mGCESEiIJoa9A7AS
BNtc9i8iNo/L+h0Bg5Nyj6mG+QKAJduaQXbOwddHj6goWEj7/lL8uE752njC
byotOhfcz1o3qfWqvnqgkkc3xc0UrvJdcCcRmLpMLpuqIyo4JwbCGnoZR1f0
ojaFiKZ4Nbqh9/XKeD2MeBhHlJUI+53uho7v62iU/UtUK0kzpqRr6eXdCfzf
AbzQtPt6bo2aSNQt+lNMwApQD1ROHZ6DrSUj6dOGlEo3jC6rY+r9nU45mjNj
obpVYMCVEmGj5+wG7u5zMNSb2kedeakxafzx9m1tZ6uzkE2duEIEJRD+a8aS
w1RUZfiYZr28AzGRM7MAqaUYO/8ugSU+JemS0pZQ3Q3CuZ2iqd1IW2Y/18fb
R5op5986WBGxKcV77Mk3hCUB9u69rTVqtYnG+UHj55nh75o1oW3qtWbkpMYS
gdHAgdCH0fj/jzNNbeIcNox8Wt7xyXBj5j1x/Jc61bNUG/oIhiAk+w8W7Ch2
496SxPjyWaPW+VqGgZGBsnpkCdERZd8UeusrD9m+LPr28I54z+olbnA9xYch
W1Udtf5k5+joz2HK5mskVdKvuitWEbbsRuFF4+JdmIVxE32/1C6O7P0etJNb
iBu2wQuWg7YG05LjPZEZqOpm9t/VUgY/jRwBv0OnPny7mzMkh4YN6wGkhjnz
xVEp2jBr8iHkgvHT0WbwNyBUqJOGdhGXdFpNVOnNxqZPlGzFmcr/e71Cjwb/
Azi9P4+0e77JX8yOqGFnsmqkMaAX+HaISwARzJSbMWdizVxmAIbGR5fuKzQl
ijmP+4Y/b1GwBWNJqIbqHeq2yxL4s85he8qy/QHWHzeB6K2DLafT0bZvDCNe
8tm3mdmh1/i7fLktMYYInxBKPUg6Z44DPXoNqig4c6a/VTh+SOVB7UUrVW67
7jcF32VYx9ZnYQvdqiYyapzJs+Lx4iBdIiYiHWj4EynvrPk9cJKgod5kpB34
O3NwGTniH1AHCogKqDi2xdsIcSzqu4qjjUIbKlRu4HUuVlRh2uux22trg+PF
dPKksX1iJZ2EXYZ+/8CWQO/RDVGd5d7bf/ZOkqmmCJ9LPhI00lpPJOwnqiV+
lffWodeVvSO6jHeV13tLf5rTAlOqIkXkQjNqmzQjY9p+aw5PNq586NolukAS
Kv10EVDm9SWAzFGPIkikTKE0VQQ9lBGfJR9FmAzsPWjlLxR8x+pTMFeNqLWe
5XJ5BIDn66X79TSWt9Udb7SXZwMMozhwA0Iroo2qd6vj4+iDsICILqoJ2ARm
Q95BBTLwmKdELPPcueUH7wH28IyI/8agiAFeGoTNsZtzRfAPCnar+hfgJE1Y
51QgJDpdj0SwhiOA6hJ6JLBTNphNooTjoPKXmXwzCX0AAm9CTxDprwTUrra3
OhgzI2MbETzcXxoo/ly/a/CJeRYNMAXHhNzShUxdA6yU2azkYHAOR8pf5zQm
AndKx+ROgIV4sNOEnN0qhHnXaYezcW+oH2Uke9ziWZCSHLsXHTwvKJozOzlK
3CsDxelfrmZLz0jgowhjJ6todM2rixat8K5nM7fqPWrGCz5fzToDQv1BzJSy
FhXpFqbdDUukvJcMSpmvhUIj8ie3pvaDkZhXPkvq7m86rbpG2CwCc1jhGZ6Z
BjC4UIsrV/4BZXYjiBs2dqXqSzrZ/Obdls4yJ7dyc5iW/GsNpJhwedfchRS/
R6nWudXe1gEHgPNAHWMPSciw/bHavlRKsLngb6kSY0X7kYI2B1aSGNJ1e/jw
OUSPbbhIUiriuCI/EQsd80kofghRKVJU9bCRPc61/mNknDeKt68pV8QzNKzG
sDj1CQDkIyNguIyQsKSBPjBS6fxbC8cgafGDGRBBPArluIdCJ2V0Bj163W1R
r5AnJHTjN7/MDiWA/LaUZLpgw+GqVLFRqLSAvmIler2wlC9pv90vCZ0T93gO
MS93XaAtXZViaUqpIVzvry1XPO/LDf/LrudI0MzX2utMJcG8Whq5bLG12Z6R
2Zo00KTLQR8pvj2g+ZUZaseqF3R87PhGIARwCL9zy2RbTqgPA4ayxAxhr+G8
95+MWB1Q/OawcW/KVEKHSOmn87p6L7BL1gas56MMlRA6cHcUfNZ0u8klJluR
+H53a+lzhrzzRLUaK2+Q8hLnepg2hiHvmDZYWpgnhYjJ+3sRlX2RYRE4P9V1
bxjhiM8CETbchdzvg4W4vr1FY4oP6IfTrUspRlJyW3B+0QUvagOqZKgtM/l1
00kp1D38xJGUxea8XxkD0B5G9Vb6iiodI/ARaJfdg6Ngs/In3+wxt2jEdL33
OUREFpxijNwxRrka0FMTqiLltf0LYk1wC2nVrJiy3NfH00xS47dYsifc5xga
AxlzC70rFMsY5epJMBl3/sPUZuiUufbSh7/Sdh9kMD12aeWhT+xYNUqBUipt
vd5BGdWcoilyk4GhQCx/UjMMqEva5EDNn4LL0xKVx2jDvMxubtJuBrMVYVUr
g1XACkGXZtw9lnHD92sV7s9CrpApwENoiTrgFZLDd7kowLEvA9xPpWLtYI2N
hnz/zoMAo7S1/d9XgWBzc295cVXPlBmON/gu3liLbpWDZuKUwSqb7rg3yNZB
z9Z+W7xwS5DEhYDEkic8kapNEWV37Xw6O8Eb/ySvz3OLKHP9D2FfiEEu+VGs
8Q8pEsUhderyn9bVmI8BQ9iE5DrXjI2IqhZr7+CeCCDbuNSaNBA2ac5FpZbV
nJxWobo0UV/gBN3JfxynbfeJQ6wde7KN4P1DK1v5Txv9JtTX26cIrhcw6on1
rvtZ6j7xvKlfzrQWNHHPSVrJH/MpduNMshg/LFnRfMkPgcEWSWhN7Oct6YeC
OXa2HvrusUs+fyVkdbLuIfHkbnq1C9tFZaW8WYzw5B3K7Smj9+oFEdxNairu
d6VDEa2uEt3nt1+P4ppVO7/PPo00eIW9WO0kkTf7mZZBoD6p+oDhVfDPwUBh
1vBB33efWe9nPoe73NsWqKligtutwIXJUPbPSgUMueekG0A2cjs1XWQew5Vg
ABSXlNNqeLL/U4gjnnMewuhOoclzAtQ/BYsXOq/uAYapngMYyqRtt0s17i0g
6rX0iod6xN4Y3yPMx2itFttw5zy68HBaBZJ74dErZtX86gKlJvoTDM2Xx/Re
AtRaBB465UeSbrIFtsYRZYXI0ai8AXpDpFSIpzLqeC54+9leFZx5MEoAL/Qn
g5VVgt/Ah+vx9IBnR9E6Ea3NyCZJbA7WaGZB3nfBUc4F53ZuoS/8mE8RriIt
bHU7ThQvhJ1RKWtTQ3UR40o1OFTQSxfPG+MR8sOqZ5NB2iIsSMOIdqtlikuo
iYoTmxnn6At91c9QuX382bd0KiSmccF689TY2YCykhjiF5qNEDmuEaFHbfaj
XxbNPUEHgSRI+Vr7+00A95kPKb3Lay6EvUp9UfS+lJNQUdFw8lRbj+iqxm4K
u3U0VyKDteDEL2k2EvS5pdGty5umkfU1nShwRTeuC6p+wDZGP05SlYCXUlFo
1cVBe1bmxaUm7hOxTOfP1EYId+clahD+myNLJ1P90iGosJJTRW9Ntjgj7xQK
r7HSMgxbrP2uGNVXBixYAyO3SukPA+o6RAyvmCNrvBjpzxeZjVFI8ZrWcrg4
nmZVvhVB1bx5YvULInMcUSqLxoCAkpXC8mLFRV9uK+t75RReU0Uhkoq2NOTB
al5BQOyk86IiBwqt+9zp4dTqv2XeUqPPPSVVOL/2iX1I22I391t3dtO8Obw7
CXW5xJFcD2bIf0LWj4Sm9uHHnr8GGFUeTqXOCRYyHHRTXL1EN+ajDdC0j4y+
OWJxfbeBewgBV53GbZXFKHVrbcYqZPBXY5ITpj3PYVJD0+qjBfzuocrX9P8g
4ZzA310/mBJx5F1mOWy+TFYHk5Wz/i/DxtrJFWE+V44/fpjTVKG8wfNqj/aM
MOYOGk0yJX49mjG+86hmwKSFYrv+uz54pA6cv9aY2mZLUD5LwRmavOImB+sJ
BdrdMMRtEc6NrCFE9j3C8VPBRFl2fccKltapj2bij4vXSzKNV/TJd8tEzzHN
cLX3SAdg/NNeu6Ur2MIOMJYA5erhPJ7zbL7nbZsAQwcxcwUEFsxOJH3isby/
T42r7jtCg9PvxRTdAUt3aVk5CbPrJzrX0+NKdxEw8xUkQOnh8P0nw5BdGYfp
uSjJg52H4vgI5hP/dKSTyMpCeK6LeJO3i0XH3l3X9AfWUvjoawit8eemk8sg
Unam6/JCcn3MHeV99KFllm8GSAr9oUzB5Lq9TuqXXghSVa9kLDkcZbVPys+C
37DRVg2E6RvIu452pQn78Efyga950LvohDDPuCiMsT2eH1qHM4T3Eld/g5zX
amNTublglXbO+l7ixLmtDAUuH0sIvdby2KnjZ798ErcfEl49NZPVMu/45BWG
G2PBFd/vOAhmXPJI6lzKD1dN8ii0vb042NPalWq21GATEnUXGEbYSwW/oko/
PKVP+luse7cr8NmBWLO6ecNQkFN5grbay5e7VNjRaYT/YFSShK1ytznAX3/e
/hJzExPEcrbYhYKAUmKocSjRgGaeCw6THw2z+pkYc1XT0Hlgd4BidA58hQmT
l1HyUaIZ/Wyb20sdxim7HYuo+s+AdTRc8JGR9vcYdClrTtmHwt3/4uqSX/aR
YXbJEsR1mfPcZwXo9YP8sjJd4FSKeqmzt0n5b2U4nbNEQCyAn8L12Tc1UmsR
ouoAfW+/ZEkjm9HTqZ/w9EEUHxWr/r64JcbDq5znqK1czrPTpJJD+pG0RguP
kQeJbi7Uw7wtaEh7azwSDqqOEtomA0KuL6Si6kMS/lQxgqR1LAoqxk7K48iD
JDMBRJd1WYKL07dtagmR8Pf669pSvQAx4h5XROEpwI7xfZIX4pV1E6q79bj2
BH5vXyHWkzQQYNUJ5Vwn/po5LE/FdNBLyBKGirRZhxAoMi4e95RcOKm2smhH
WKqlfEEy+MeoYc4Ahzb05st9ueL1izzOtoAzy2g2TlWWzSuicFRiJtRK+QHU
c0L08vyuvzpD/xitcUKAvES0AnLgDKet3nKPc0g+AQQzNPx9PSRGRTFdb7vS
/iedgpzUcDC3qo7Y3AQBnxiDhZ6VQMVt+Hy8LixEZPIO3niM2XEB7lQ/I9Qr
xl4cEiYRFwMsp4goMqGBLAc/RV1nJjXnSt6iw6OxwRVoZ9Wh01r90YeU7G3J
AYbuoWFMdqWftWG8X0k6yCNgmV2vcmpc/vhxTmIu0cMVVPf8yoODt24L5/BT
a1/GD5gWeFEU6eAbc8GyPL+4XnkwbAoLVKpaiG6+PpLpkRkKegexQ1jb8oH5
/AntZ82eK6Gmx5VL1OAqTVSc4NxjZBqhM6prGIx5gseH4IJQzEDSx4gWax6b
Bq74/nX24fM0yV+gyUxvaGE+HLPVPcq0FcmsBbPQnzaoRoTT095M5xN4jQQy
BK4WNrETibHPQV8H6mmYQJwtXxgG+m3mUNy8xWwAoWe310bbczCMBzmmnHn/
wGvhRSVonScx6ZJhA97K4aRQAfESIMCUbKkJM/RUWTbb0o725hq23EAt5BSg
reA3igzFdKO5DxHylwRC+jbpDWtc9TuQM2UktNc/7BuQYKeHokvjgHNAzXMa
vVCNhudyQ/X+P/bQdHt39a+5UbwjUPuuznAsMpamohWziqrsfsXGiVfzFVXL
lS1ute3gBr6KfaR55QU2TzObMSkmlLQ+A3czDs2GhNvRnHGMIVhFIvV1o+Fb
Yon6mLeaEWpwZbI/PakSBzyIebrjiJAzoJxpsFVwdWiII2t7XBnikQ+sD9zP
ZcJ8obKSKT2WS/hf88fYktB3lTJFNgOUBkkT/Rfk7+BLvEd7KRo5Wq3QjSwA
G+V+PFnFbnSV0dv5Pw+O3v4DZEwTh9dEjyFLZ8UjPf5byQE4KTFcZFfT2MCi
GfIuutA53u7yntCQd5HlSr4MvqoIno0j3aonxY6dcgF8i1cdP95mWJuJA+Kr
KmnB8URaUaTT5+y+kx6ulvRA9qorsrWaCnL9XdG/APWG8rAOU56bxp9+rOPr
rAc735SDnpf+7CDR7z0ctsfQT54lIR0q3yVqKGDRFO4P4z+CainvJv6AT1FM
5R0lX3WdhI1hSJ6PHDEevcAcpUid3SEWsqaxsh5e55RkuHyLrrR/6zSpa9Bn
FM+GuDIMqwV6xV0ot4ZgXubT4VNGkXIrdwCt435QFaG7Woa8QY8mXkE8lm3o
CFs3ujQYt4+XxmSzefF4tLeRICBWORd0e0rUyRLxpRp6R16lbxHoGacZTZxz
Sbp48kdAoNhoG1/sjZ/BUa09GJpMrAjfa8aTZz/PzW7k1yEKhUnusJH/Gehv
glQYAtCPqR+0qLtXV2hawG6jrvom8enAu99cSatXbkuLfEoe0T5N2djC8M6o
s2nmz05RZsNb93ddzpIR9hRgZijkA5e8WsQRmoqtWzWBAGQJ7IkkEafobH+l
MGobSfkyeKMO+/J0XFNFq3VqYltT+UILzWU4PevrbvE0LhXr6uCwAcJUQF8q
g9L7wDD9UItJuOHUFkOaPNdsY221fEcXLzhyraLtLfVi2NA/M1/wZVYOfxM2
PM9Y5CsDMlddpPvnPRaDK6vaHdShwKJAlUwCFUa/wQDT/rvq0y2hz781v4iu
DpfAZEuPag1nxM3bjpJIZZQ03g9Ug1nMXmtclYhoxYNMwGCH5Vai8K2wH+Ua
qE3tckgTf5jI5IXr7G4SG8JsAl1Bqc32kW5GDJZsSbyRn4zvBJRd+LhP00HQ
XIyL68hfMyaPO29dguZ3yEiJyUP2gKHbd+s/SAwHwdCN+ks4ZufFi0J+yE9K
1DqC4GN84ee0BpF2N+GzFSn7zC065gdyqF/Ea2ZmDybIw0PdWzS+muWu2wn2
27WV/rxXelVq7XaDsQXYsVSkIJBXUxTrSzLS5zw82Q1OxAgBj7RqHoa7PQ4j
JhUWHvsXW+DJLXX8BpJCzUav8YpmillIif5mcJVLK7uPg9iL47szq+h7zH3p
oLq7/PsdEF5LbGiqFzBT+5wmuq9DGHWk0m+oQirVHniQXC8QHeN72yOh6acE
BqzbnLMmdjxNTsBG3VLS058NU2Dnk7tu6oM7+MrIzAIBjv2Hs94D0Zmwjv2z
MlPluIPgpzOpR3VAX5k9V1PgGWj5zsctybzk5qvq0tASNtB4ySbS968wN6jP
c3MI3WUhR7gY28j3LpD41Twa91xajWVDkAr/xP9nmylnyJGvL0j+i7qVZeJi
3h8ihy1raKgf10f0WbL8h+qDkgxYznxyzf+nwYrAjmWkwrPq09oRTZkl1O5J
6PhfqybvKogrK3c1zNlj3SOjRz6T/gnHo77qHJ+0Q9lzQq/1tn6zvV+pHeB9
KUBwW0fjvqmL9GdIXOq+8ZdJCcG6zFjNIQAx3/7Eq49lLOTe8E3nCSaJA7so
dkBvYiCdZQKfmaRE0SLgzBYWXrKX0HjMmIoA8+lHN43uMWHxBrpJJbhrSxfQ
T1ejrnQbrl5VF1DTItV/HGmLSSxlwE14YdZiIxHnJOlwhf6zDwCjbCL26U+m
iDK9RFWvJfvA3aWbS2TevJ2ya3HBgvN3pc/qUCeyx+6J3VUrStq0FLi/jPo0
DSOT1zwc5KFjDJO8C6ALcxT+TfuI7mFWzmJEiGJ+LMl9oBeYJrOSAeNB797u
mrvt6wOKZndCJKPlKjnFEmJT0GM8vSGP873pSZ2zNHSoM/300IElgeLMIBd7
T1F57fNEci6IehVI42anpnY5MxDS9DxDtJUjpx/yLUG0VrfoBECtvp5qJuA2
fFTybjd0L0RhW2JCn/2Ny7mD4sr9GM29KSuXxsxXnQbbMB4EeDloy1e/HdoO
R565TtqDd/qvKC9lNXYhalKCi+rAiARFp3+MxhPkGlfxpyeZqnwI2Qp/To97
K3GH0ZjNqD/goiStSZU3ZYXIiGmGym4RssvxKvuh7y9u9EHuEUv/xRNfyvoP
Hp1sbRlhp8KL08oCTRSPhMOWhrsolf0LUbss/RTVmvunM4bcGTGKLQHvK+9L
wYl+wBo86i1xJVdUb4BKTDcipEdbp4Q3fpJLzp5jJwWN/OtXQwaUBxrjWbvD
LLqaoueK1dxk3SQAtWPG5R/GKf/pUeHsQ85Zr0re4ybV+3hMKAuF5cu7POym
u9lJ9frwe3uZkteIFs2qBYYr2Vds7hrttabqE8+V1svMnmsc5Mc//mgItKOR
YUHHnxh8+Ia82HQGIOHSrV6/eSKuWZRU5MQrFm8ZWXW/uiQ8dz1kSn4RW0Fa
Kv4EHfYKxeM4q+rFD+4A5kNK6j12L5XpNG7xJgZxZDRzroGzebAcC+RN833r
dH9B7JwpE5C4rnsXw63kEmyFOJ+59ci9IxdVCYXWy17DPRc5X3dIU6Vp5UEH
dgw5gCuSXEfjeF5E+vW9ikCE+p9kKtikRLA4U465sXtxHwhsHYqIpRGW5HyZ
rguRWAFtjsI7y4dXfP0hT4zaCsXvECk5Wy4/NdQO7KqM7R0a1kU3Cz+4Klaa
d57lYbmxvz93bsa09/iJ/LlaPYbHOg8dub7tVdau/p0uWkLGUEvhkNBvd2VX
2NXMQvdU0z1Lcc5ckFgf6VK91pon6w2Z4+JiO+Tg09BRmhx//MxKCLVbIFO4
TlnWY5LWKOE65DaPJfhxa3pnbMRhZ+MlYyjooyxsJT8Z4xWyj9Kvz0zI2TSW
SDHFEHIzuq38D4BtFz7GW7Zr1UOGt54IBJM6UvSbQFksL1dI9rNKTnKB1Ig7
KZhI0ubLQCUSOA9TQje/S3JQN3f9FvtVtWv/taMaKbp0X/Q/rsPn4055Z9dl
KGmY/rWCzZe9/nDPN+X9d/qO++3frfFskxB+y0jVEnD6TTnFbRWGs2jTJJ4h
YeyKtKwD+7wW93DsazKjy8vzlZebEfJQvv6y7wwsMe+G+KII6ERa7y5V7OiR
aJ+1xWJO/kqIi/2/VOAWi2dvJa91Dacffb4jmMIjgpidrW4dkEuSh22+5ZHs
ksH7AL3N77cgybQ+n7S2vbYsjzeeOpOsFNes2B4zEI3wONhGzKQsDWnxwTNl
/Xz4mlrKv46Mc8YYmt7q+YBddyC1bjsFLRaq4zIKT11nDni0uTl+6SiXyenZ
qSnlCvLloPnGqCrLWxrgN+N611uCdoH6ndwXFz0gMCj5p7/zkJTBewtU8lTM
pvROcx9rNLSVai0nbN4O8UtcwCcL49TM+H+o+0Jsi1d9qkUNNvj+8OyfG2D5
iisKx5XFbISNfCzdQYGWuUKfuOnk3KHmB+XcSamMPypnqAD4aMKFI+I6zmIk
LVy4h6TY/xxtkgmKtPZfDHSNn8hxYNp7Vrj832YLMAa/lpRzLGBrX+T1Mpp8
2eSpdMrlCOaw/zQUI4IKahk7lARLDhfrJ2agg/rQE2nAy5hbK/ZOCstaUL0d
LaraLb5qkF7nP1XGlwYWN70TjAV7KFRtjtpgIE4lJMBrrQC07MmPv3qghRV0
tPvnZBcbXX67DWu3ub7aeUq/hCWlcXom/03ogA8a/fpQYGc5fl50x5RNzGlI
qojRYSmwHigqTzQTTiVibiJcLkNV1gP1FUHaX1queIwKb17KyN8IotyfOKDW
N9x2o/YYmLT2TMdTzK4U71yZ/kEOjmYOGuRFonRIkApQmuqI7lc/LBbF9vvN
UaR/YMUpHXo+RMl7IFJRrgveFXetkju6VtcH58NbbXFsVqEeYDDHtFFHl2Qy
5AszdozLG0sZ840vgjpy8yKabvc9MiuXIFEIxyzbC7H6WMLDeCTWPAAfKiXG
bQkxCrw796vmacPXhEzpLhvVbaB/GFOHcsHYN8G4FK2QPuNebb9S9ki2iDv3
ozpbOY9idcR4s6XBQpkXaVS6EuzXKFVZDSgchvfgro81SJCNegzpoiQKv0an
CwdcemJ55MQVFhwRd7gDKrMTHv9dNbg1sOaWmA+P89dVMN4s9fERKFR0MjZd
DV4c5woH91y7+FBQ+7EaZ0LbHzHZPOruzkzYyNrakFvY95hT4Tk+7nbq8xRA
ahHnKPqDi8twdAvyfVYy7xs4Y2ZAsRHLy2rswk6Da/Q119CoNW7mZiC9cKRN
cePiG+D4civJ7U2CEVwQZFnJ+mO5I7Tojv5rercIH3v8F9Hz+f7Il1aFM/rF
ag8q/dQR2uvY4hMqzBPFp4HdU5rpMay17aFngCFhsCXRV/hc78G8Q3v33ihA
XpUJlhf7cZav0IXXgKuoAiXFGyubo+KI2c+HK5OSWMy8nB9S21V+8frZwz9o
UIYiaCGmUV8ofMVUw5tm9tFzGcWsy1LZL1MErlDtonU12fyFkezMTR1Xcb41
Ssfk1TwtM7X+9ESCxzul3RQa/GtAjiAi+UJgoHt8u/kr4Q2rcbAR9Bz5bXS6
s7JOLQcgXyi0UV52SodUBtfP3Me9Zeb+x7cr9L135BmjnoP9ACMgya94UoKs
DSGAWMY7eF/myws/HzFrY31QR3y5od0FC1D9GsjJM5VpkhoFYyVVfnotSVGl
FsbFXb7ixvOP++F1BAlZqnAfxOtp7lZ/9JurmjN0P/3izunm44r/YfvRSoQY
BeiOyNFFthkbRjk5wbQyQ1xhWpuEdTqlf2/+r9cN1iLXpSUJqTJP9ZThYs7S
eCm4DgE0R/QGKoAlcW2NbNBTqKj8oc6v9quRrFHsyXxhpy43uXY7Y9zhmyfS
mETfjK/00qLF7+XTdTspmPjUklbqRkz7406uMHv2qHopX2x6L6fVVt2jfhQN
oGKRdmIAWrr0NsUYhUI4mNUQ4vRnqeReltXhOXBhD8es4/ndFehl5QstKIPj
bdBe8Xy52jwtQ2EmupRlWt/DzzQlZAdMmbX9qpJLfOfXiZ5Y8IatPGOrTUxQ
ZNsZdyRwfBnlIBjJH7Kd6QUFlNFfVGP4a9LP6BxTzAx2QK2bDbCKFnJsphPJ
kqPHstMXvltEhcKwdoADEIlRFdhVbCP0MZHwOCu28Takr1eACO8TeKP8nmbW
L1/7j8lm/aUqicQSTefItEzjqg9nZssBMkDMGKk3Jfw/ERRccmr8pP5v9Mgg
j+wGEohz628za4P0skHUod8CXUnNCillFZ3zfT9kojFuatIniHETJ85AZPqo
UCy5gM0doR6+ggjmD1FIEIECkrLkEiolYXPOBCOelp38RRrqAAWcsCoRLYVM
K8Y4gqIc/k06nk9pBP6MTMthSPWiZ3t2pDkoM0fkfNU8NlIkJseRAO5hvjMR
BG/vJ9TtGbgIQeN4Yv/5H1aSP10CXTHXI+BeeOpaL1yp93CusaRCsTkNWES+
WaTBiVVTUR8veQFJy0HPn1wWb9v1O9bBQHOLMA7X6wZ0OP4izWZ+JKU50d+k
N7B5+O3yODR+ThK0g2GkuQliPchL/oYJJIW+AKrFz1On5QjFkm4vECNIIl2S
+1xVyfkOOCq47SRVblqyOLS0BsTAbikgMcCvrqATuCHSWyZy+jnE01+NNfds
3E5PMQcb2nmFOIkl1Pt/iGxq3VQNKBdU6WsufvGzXcVfUuui9fdDOG9vIMZR
iz0aozrEyCT3XrVsoi2kVkfruaJqiEczrHg5m6uI0mmmnLgmFUDIxJs3zK4o
ZBcFYNQlNYM4Wh69kXnDGC9YluITVjGata8CF8V6At3kJRSmTpGGaMKEJN8T
QKIS/EXETmygykLPIa0GUvEckrj/Q8RWOsT/ZwFhEMUKSt8+RKHEHofwx3vx
vHBH0daAlDOTJjdOZ7bZ+q4DeGfjCCzuO22LpBZa1QGMZIP4Ifag4wwaPSff
itWp/rro1NMy1QehDee5XDAH4kf7b4kyhmq6OLIOG+bkPHwbMgfFdSTMrKBm
2khAqOrJNbnzPK9Gkk+ZDeNX5RXHLetqiQUixPJY5fuk0KOhlhnLC+NVVIdw
hMtTt4JmxqHPT8dNdXgQmM29mysMeJMb/oCOMCMgNMm5YtJtvUNHQmTsj/Bq
QeveyMn5k/hwxMooS2BpNrMy6w2RJPkZaML+WovCJG7fSrpv+f2z7/z43u/T
CpC4KVLQmDOiyk7xSon2w4ezAod02zg/G3RpIoxDgHCc6ijT81DkgHZYsF/0
o21A663DHZQ+taz8FKflSwH4FWc9WkvkRP8Z3GVmj9jjjevNHhmFCPrKPNb9
mdZWk+3Is8hwcFiIqTlQmLgLdqGZ7Fm2b0qdZ6jOkVjPj3o0ZrXUt0Uof3w1
3Zvewyr8FY/GKiRrZdzViUqYv/TYGJrZMavKadv7tXHKu88xx7vy4WRgOt1m
20aFwMoijl8ixdyyF1VXXcNL4qfR35aRysdEm4+esUUx77EnyfY0FURLpxkJ
s2GIbDlfv83C+hgnrBuGVG7IeeKk+svkS7l/kAp//r96X39sFzL1qEoA6s9c
cAwD2dPlK1nb7r7Lp+kPLRfTNx4002B46dPEEWIOjh5Su7CzBdNZUbbyrDrZ
HaHaa+wNbdhoNQmmwA8IAVUVfg2U3R6fBRAoi6txgAHfUBOF+ZZbjwr3Zyru
qhsa7oOAVTAiZCDXe6sYWDckMbpueV12m6rS/1y1S8SH5DK9RF085sdB+ik+
/YoSLPl+yVfThcmRHEwM0MoY6+BIyoy4xEMckFQmZTG4CDSCtuWJduVDo/C8
8wtpnXBZpPtzrlLiEGT2AiDTKxI23pkrSrWoZ5oklqBBApdHGInbkIVx0byn
IQlGTDEpDt4PYc6xx1nbOYeIBDesoF5g27cdEN3Zjqy1r0JCgOcZHZaeTMtw
EEQBm1tTqMBudcQn4XSKQCbkpqkoYUZaEHUkJjgePAuGTDZLA3AqJlw3vjam
f1OKcllCXN8yXPcAcneFjk/t28otmBlOdchFgUZqJSWOELY0WOc98ZXyIWaA
GGy8riq19VanBJZjBOMHrnKNJp/589FVchqPY2MsZr+Bi5i/pE+21wqa9nFL
b0wFMRRK/vkDt0Qn+eN8RLp2lTNwv73Jzd0oerGGHdnzqFC0N9BceypRlOUK
qY7qq/sqGTyNCaoFzsUHluP+RdbBDNTxDwmUk2wLZqU5Pqm22zuptcxaHMBn
FcGwqTVzWMS4xjq0tLUnhNwelgR9hyXNtge1qIHwBSAdm1X1fOgPYuJYsYjW
bTP02e4qBRy1tVL7eDi7tEEBHFZcwmKQn71VP7AVoya22B1+SCX/NzKhbzOB
lqmMizLLOTyHG6QOLHDXAOchGQRAzhU6dZQxQedxwpKvDqr3MQuyIuUSp7yJ
6sHLVI0//QJKlzKs/AikiQ04UC3l1TVrxykavQLyglz+yAufcjmyZq0cpHh7
ZBf1YFRZs3Xj5yEJt3C5j1XVotWoPJW+C8hQVO3aF5YWNkQaFoRvPnUfO8XA
chVCZgLEyy1Xsqn0/qwwkOIif/GwVSNBsbgXd45PPmgdZSe61/n4sGPRre0R
j5cqs87Qlkch17CkSnlFcyNcirUgjemhN+Ud53CY9ufj+jVX3odfwq7du+db
KuVsqo72LrjCA25GW2wSDAaRrOPCBg0YgJm7/R5kX7vRysqQ5liCvify3Gaw
jFu52xMiGZbDR/5t0P0ER8hyB9YBiSyc610QyheyqqKUzMFcRAbKNiBqOG7a
Z1KfgGOGRd3+8VOZYwpYiJqFEmGobbRDKj2vEoO4dgS24NJkwjG/m8FDKif1
h+0Kr+euQgfbsxrP363hZfk+GDnfPrAi3As7K0Y62BtdAnH/y1mjiS81onzy
+PFcIpbYKysktfW50A9Bes88OlYSS6+3ZYd8d8ZodcNEq/4MyFi7kOaQtQLl
ois5d31WNHJi+NwkGEYzt0mQ2h6QMoGd4AcikN5+6sL6H5ijsOzi1dYUgqXm
9eCUrtGYKlxelGm8zpSRP/8Z8cFEv19CdRsCZBsQZKZqALgtlJdSXWF8FqhU
7b4v6Mp0dFIQ3cNSv5R36eaDxfQAiAxIMo6YPA4K5bPsapdS4usJ+se5mrnc
pm6esKFrpa8+RR/UoErZMWZvhyNwlzC0j5QbOw8bNyM1IxyB/KIJzCxg+Q2S
kYRZj9NSaxjuVFtV6FHGcwVedlWYA9ff4GhXn03UnsEGFQ34mI4Cfre43hoJ
nddGEbgrlnuQo5OPdqI1nCkDTMn0UPn3Qfc+0NcRh+HUe5oMneeFT8IBlfjU
ReBu3nTqakAsHFVET8NQ+TD4HZ+KU3ARKDDWqVWAW6NGj8M8I04AKslxrQlb
R+4Fj80NV2lxKwwzHsDAVi/aVMJnwV0bLgZZocNfL97fDrWS+GgLkvjPVNTL
T5r1Ws5ghB/kQSCF6Won/RaTvBfQjMudo0axjxYWEpKRnLFhdKhm/4Vi3Zt+
0DsvyuMJCX4fns3PBuoTOzyR66R0ogdgI2oHaQ3MgRAQ+FXHAnAZcWw6k2BX
aZ9OEqxwDZn5/61+5nhuxlvZWARk+m3p/ZKrO73Aqn6wsqhLUb6CIcLpCFV0
ADdr5UoUbNbfIhQCgJnAPnt6oZAG8wEg1MXOlbvtfyVE6Cs0hb+1/w3N4Bok
h1d43bD9QJTxe7fwbqQkvKSWD9tIkgql5Foaa65U01biRpkI58YZlPiX20bX
eDSGX6FHJtoIiRozauSLT58/UEKgc+iORCJudtQ+PpK2P7y3Qv9MZWVlYiZc
rdHfSBylyYWcK7H27q5FnHYsrBr2Ma4WF0T5g7HC5ea/wgzwM2AQG88eErm1
HQNs8m2vYeTwSV5AHArm80jZ4cJbSV9oCCK8piaB74/ymj6iAJSu1CnyCDfE
K2EYT3C9VmZAEMaOIFYxTfBHxsWNndiBRRl2fhogS7TpyfebHWOAQeEtdMjF
mRnNhGaMqf4dwQBLVNXEBKtAvoqlNX4aPfANsZA+YRtbrf7WGX0O5ACXdWky
9LNvReY4ayGSCUuGXBk69jPoSe4E0s9eVJbFa8uT56nD/j0vwSsgeDhkEBeR
3sp44av81ZT0SZ2qGHfpE4s3ME6S4OLGnF7TnN2wRsSk3hPC1MzzohgCAEGz
9hxaMsjsE5FhrKp44aRgNE/T+eY05oTUrVZgOxyS8WMvsqoqQUqaXI/QoUmJ
Y6+Zitk3cnf+TVKwfva/AwuKIac1Kr4zswVpwx/Ua8oKNYgI2OU2xRjBvW56
BWE9NDa9ZIUqYeJl/W5OVMtgH421K/79tOyXWJJpJ1ULZYqRUM61H5mqairz
YqRDBTiQkjJv0qlqExAuFkrbGK6oZkQN97RikV++V0FZCmLO+F/D9TL/Bjhy
kRson66AUtUb8JmbsoTIUuQZZrIQMQEyUgvu8MuBpOG3gJFKmL2cyHyju6af
sbmEeHVD+YiIgYvv9y2eIdGtpae3hLKM02isMafs5BxWsVdbNCofL6oNH6iZ
5VhvHQHtFTqINkAnOiVUC67wjz7gI6ORuLaR8YdNgWOTY3hxp5q2Wgaecjqo
v0ihhhwSv8dQo6sMFi8oWZyd/0cMPbPg7wag5116DLQ5dDOkd9uy84f4Oqbs
WlUScwQr6tJaiTbI569uzSXiS0z2pUskShrEMVCklUr3yrmUdWW+1znSvUpp
PD8iSNbc6BJS0g+DZs5f+wWEB2GSNUeexBxrarpDCVRrG4fCo/We+1x/TZbd
LkznGc7uWHkzR5O1B2nB9N1p5m9LjMx9z1iOvGhS1khWCoqGhAM4ky2nrXdj
ljT/tjNvgkJikJwaDMuqgx3ke41+wLthVZNeJho6vp1HUn4U2CzplhREqRp0
XVE4K4OZXKkeknHojH7cvGvrfaPjGeWaYkidgKcTaH+0xGRnjuN8pWRh2777
BeaMnA5OcbTL6yAGyj8oi12bvyRYazp5p5/H2oUBsCjuVeiLYrp7vm8qVISj
xpkKQ7Vk4TVCuizFjWsPC44kIiKiI7bqKIi3zfMd1xp7xlOxbaWcXzTK2I1d
PVlcep2QMk34plOEeP9d0RmUHdUsgmRST9osSdXIEzWbQiJkPLmLNeqDO4rA
OUTUG+zNn0Ck87aDUgjwmCjIJXEhYvOeRPLVytr6A4Vrt8mmy2cnXNwHtmL4
FkrUwyuzyoPO1nWxP60MW+6upkKMrYUimnWoJ2MdyRNSybefF7MPjwbOpw82
imUKHKtrmCcI4fB18VGZKJV0ALGrFMuu9AU+9euOptQKj5SIoSIhEDXRjhPL
1asrhbLSLu055ONGhTQ0qSwGUbrYbwwbvU0gipW56WQbkqLpjPWejj6AnrX3
THIzJQncP14LPvTKQvPXszfQEGnEBEjyd6jwP+IqOaliNmFKJf4mpWctzVT4
nAfBLvWF3LOZIHFzC335NjUrLB7kaJabMeDEOV1VQROurdhjdTj13qH8oq87
Ku7vtd02D5eQ5n6uVREiUwjPex2y5qqMxxSQymkYcgqP2yn2pEGR+lKztaAF
isadUMphGIygxsh3UnU3HjI2cscxMgMDfmrhMZfldwMgT3Tg8ySMpyE7jA+X
UW8WqIvSanzd9mf/q7LWaZc/lUGGtVjpHL4XzbvfplMSv09BAfgsrpEeKKb8
vlLJl+OSa4w6PYItzmsMWc7Bo+Qgy3wHlJTgUQKhDaWBxgZ0e/QXpqIZsLko
nLZesS84Jxx4dMsDp0iSSWYDx1zivTa7ItFLY/UE6yYRkLYnrtT/NGo+Qt9j
vFXR1rmjsnBph/7UqiAHdOCWqFBCV9KE86bUrslN6AUnuOuFK/3QZYlQPi24
UGbIy8Vvcuo7n40DDHm2KhFbWcu4YL+4YveVXdfqyDJ7UDderI4yFNP1cJts
T/lkwAme2FwIZcZD2/8UefyhVITmmQipfiUGrWyiGLypes2A395f/nZswGMf
ghiA9NsRpr8QMbJqDA0ySINPSH8XIYHcpnL+fJqMxjLlastA3J9L32FxSTuE
EJoWyaHArImfNk5P+8aDU8RRNLAkpdEvc54uk5btMopwQykobjeMjGtJx12a
pfmXJYec1O2WOZoELncvSA2OcG5IysT2V6rncs7ank+7SkseyldsP+OAcj8C
VqXxkrCQWxtnqtdoLR05HPnFeGmSEHeaESaaZBD7pwf6l0p0x+iy3TZZR791
MzIamq/UPOncG/G0ubgxkHfSOChQ1YPBN4/Fj+vc9S5EalFIl7CgzNouuu4h
lxhhpiwVvxpNNTLePpNUZBig6IxQ2Gy5wJ7h854oJY9dGPu8MtcqFi9y94ip
l80OQtqwLDyGgFRe76P4LRopYZF/sxPJ/Y5NFAfRtnkMUrYrSDtO9OavH0ZL
yWe126kTi3MwJ8E/ojZhtifE0OjO1TVq+6XL371VR+9EqRZePDcaLj2otTYv
7YNwuR4EjHRCBqFtLUs0UoT+Hhfa3T+8p9gEQPx1Px0jUU68UUZTCD+UeCq6
CwxyEmbQ8yv2pWHitbeSvseX59L/N4pv4ABxovGSb+j5TEF+kxHnamCK6CBx
UCdFtApA3bYZPYggmokvjyWYvGAXHIelnOGUxM2A0KFNjkH0uKMV6Vnzc+iv
M+pjUA2LNvUNCWQSXwcgc4/c2APF0chYwCXp2s4GlC6YiDVgLCCEs0A9KyE8
m9j32oZICVKO/ooX6ncELC8uKNBW3JBttNU/0YbVYqQZVcwdNCwMB1L2wixS
Ce0+P3og8rt+nzFDFGI3YOents82ynaVitggCbh/pZ8mmf5qB2WsHVr1xwbF
0sgLAwQRDjwFfM40qt49zf40JGzdgqfhDhddbEe4XtflM6oifdtARcI+H98H
bNtjbt8phdLi8NhTRDeHf9LEYhKinrchoY43z6VzDDzkx7SV8TQxse9LNTnX
1SieF7XWOKDDITxyK08kIuOQlvpi4pAfZJ17/ucN3g+wkk2C6M8dS5nFuO94
Ns8hTjioilwR9EiH/TufsiTaRPf0y2zFh+418hZ6HH0u4tRCw99ifKiTtucE
euFIkbIHPTA28QJGn6/t53JzfOOaf6xYNqVor0fh9z5HqSuzzp4oSoI/LGn6
wB6R8gsfVVDVW5LlbEBuNb37tz1d60qG4LbY9fgWCHPhkMRKF9a/wimwYsky
STvrR6Z0RVuaKqvnC/kcUhUvpkXqY/KLeRyTM9UvGK1HE+BsgvuxDIsKJEfF
hO7hLXzN69mMmOjASFsZct75siVqqY4sBiKS1d6AIK0NEevV3o6d+0PfuQUv
PrNrRyNlASRrHCeYiy8RU9ttGY/8NPJ0PCyQJlJRJCipo4ArWE+2MrJA11hH
3QwKqiHXDDxvUEKZW7g4voINmhT9iCaAfrQtzARRFJwOe9qF42Of7Ud66kL4
cxduZVT7WjZR2MGTvzVGm9H638ZnO4h/WsWZUjtuiIh23kNpJALQybR3TcaR
ApGB3EzSKkcGOlDqRtjaM831JUeyACKdxANTs9gOyYRPPwDd9EZBWIjYvHO4
g6dAB+GePZ98LdmFVXETyHhDxHFmKkb5EpN54Cu2YyOomCarMTg/bvu4D6dn
mnxjvRYbWkUNCM5+RkBp6sEkD8XHQ/fv4lAYqShfEfNFEHVGJ96tOkETUzUO
aEL4vwgcyILBQFKYD5Ih9sTfEcVCGvZZrFZYBjD+cfn4GPlbvR1cgFHPT3hU
l0a9EEAny2vF4+jR/ocNA9XkbTc0baF0Fkkwqi41uSxy/sI7a8eb6e5UmbFh
b6BjJb/NZh6ysVi1049+QZgcAhX4BxW1w0tO1O9EL7zAa1B//SB46V0jakrX
Q0VtbBbDw9ZM5naeBwtdf8nslef81jkWxoYeXu2ZqWbL2+utWPfMnQCs0TbD
j+1yLoXhl/1tZ3DpPl9jxIfLYr7hgliN1yWlfjnhLTnLCtBOtCyNspaAVS4R
h893F/6VHux9VkGbLWrR5NVl7zsX5IXfiISUCoS3FpjisvYlsOy2tu16+3iB
giwbv+KktbNoqubl6yEcW+qLcOpxnEy1WjnmKAimCEl2bbm4PhIwK3htbAXA
A44LiWr35JMp9zvjEkxUDT1J2BTCZwWaVoajXBDHWdGnpbN6+boZo2p5HTnA
HXmMPpe2m8F0G3umClkLoYIh82FZAbtcL/ALYBUuWjl2QHwsDRcHzbrHkNyH
qeXyJkjzPtNG1sLFo2FuOV34wpTNZHWORbt8slZNVq5LGtdOaCSHp7Yan8Sj
gI130XLiBEFYi5HLWYeK2IjZtL0U00GAy0FxHYCxMHPkNsheArfhsDOxi/vp
P9JeyIQvBa8cLfVofDbLnDtIgbu8/iGITxSwlvxx3ZZVrtaa5Cb0AClj3UpE
S6ePg7us+v+gG/Zf9hrnXHmPK7EMN3D9J4GM+qYczcjYLR54RD2O9K6HJRuo
RAi4BwEgh4tA9si52oV+ZnmsnjfIABdYLhOQKDkzRihkncyE7xZ/im6oBw6/
6yW9lwYJCUzeWozzG5xlNjwcfC+3V5WpzewGXfxd6aPulUCKUSVHOFxL/BVt
sFJ5wW4CN553GTSsQrhh7e7gZRy+uFVOHSA6b6M/6SwmO1fIFq6zbOo9HJN9
TxodoE/KKtPwyLMWtRbEbkr/BNfsc08MwiaH9ZqOH7Fz0G3dWsXOzkFUd8fq
Ur23TxvHjJI9KT8GPmS+pHEnGrgjLWt3fcMVeG8e2pWNMfI+K2uB7KxbRRJg
K1t6y7evXJvfBpOKSzmz73TTujGnu9KfTWUicHh9NDgbSRRxDyveCnakfeGG
DKEa0F6sYTLxIa0jKC/9raW/70Yp1LdDRoEuphF/i9PbAqaWXNeguuyrlLlO
+C8x6pKrqERG7R52ibUBRDqw6P+nVvoG19Ggkuehuq+LcZjyQ1ojtaLJeAho
s4Z+9menct6ToItf1pA60D96NnVYp4i7WNEm3EOm0ql+/G5W8ddxTXTC6Yir
FJOzHRykUe+ypiYhmRCIbb7Vc08borUtYFE5TR4JN+TXMqfFSu9M27BlhTKG
pr2Q1qcj9oDCrTfhLhTP7/4Qhf184oUx63d733DXg0mWTyRFsOyIWZFAzSJ1
P6SG4h66gfLuXKsrrV5mgwbJJlVUYGeOrEw/ScGY7z0RFzq05m/uOvKuCnyE
JfToTdI1nlaiJPf7Nodov0Ph58/oh2AmkABbEshLuNae6g692CKcbazqXk76
HIhvZqlGVhV8erpEHpMOw1kW7DP3A/tkNPfVBOJVjaLshAbC3NsvEbM74SbI
wE/C2bW2jWxfkkY7MI3wO+otCmobPBXzCPM6EScpsELbKxSFoPXu5t8T871S
QoPInaG/1LYv6r8nTTDnuNk4M7OCeRDW7squ4a+rwzivf/EjHScgmK22wRbN
goPBqMGwIZwFu/b4cj7OkI6g/Mr6t/H+qlVly5GOHdP4ROSvGnNE3PPzCUKl
f0DyzoWVcJMSL0vtSMY2/JHhsxh/ryhd4xAGDQsss771nIGDzHhCog7LwVLB
VLeGYdks2OJEwIfqhIyDWHw5BV55VEU9LPr9cbT323ks6qh+rBz/FQWAyBP3
gjAUX9RMHYSOO0ZXyfUoA3pGZT7nkskVI+3DPmC2O756vMfP2V1yyjsFJyze
k4a3gT9rQysW7dRyNQSNYwfj/shZVV4YyhO/upwqwX8BO5o5DgCbiUBFHVKH
0Wpodk3uzcAhUg0+/Q0ViSGJRB5TNL9Hx0lOFd+ma93ed0pr8NvBlPYPStXS
IwAa08vB37NFdVEOiInMYJ8b+a4FtCmzFhCyXElveWqykjv6djlqjE7rO9J5
O0Nka3UgkGhouWAOOd58MevgBMuizs0VTd9zaWithTtGh/Wojc0gVIdbxW6P
qXVmMclidVcl2jMR34Jqc4Xx6HyBTiXyjBd8cLFCjdFBD1YNJF8iTFboXNZV
ctN7SpkJPku83hoBaJvGwqV0ddAhuU2XmdeiEw6eIB4iu6nPIMUVRWAiYL/L
xep0YjnpBnY64y2Kefi32rAh8s413TrcmhnFnIZwz5e9xGMY5M+nST62FRQG
xUsBiaWUztPxToFSfkmuSgonpZV15oqAlVPPyTN5LQsP0MDdLcOm4ci+8XOp
vZPjb7LVz8K9Opxs/SKcTVLkYnAamcnuSa/XB3lILe/gUPxPzn5FfiVl8UFp
bwQdHBK+JpBStFTrH6bfw3RqVNM2OuXT11FFnBPd1rLGuyfqWhMq+AMW4ASx
U1OA9cvVJXprPo1qp/uXKqVB94UiI6aYBnHsfxcvFOs051xmlfY6tgcFIQla
ELfm6Fn22MTvWxPr8dt9nQF9kB7VEwOZqeS+BaLiIYtWqiqgAD3VTKW2pPAQ
EcOU/hPz20Fjz3IDMhRT0rAlRfMzRTZtZ7ZU6C30vtd0cP2So1SsNKyrQKmY
ZPDmRGMrvehN/70LUblqAh7RPBdFtC7cTiN09fzlUcfYSSGN6NxMlu+5/z08
oFB3UGeWZ7FhCTJuYDQrl8RN672Uj7vHBC3MN5pym+2GgYbBguc8K5VfFbnm
xPmxAryBoEBqQvQfQ7OLUaKm7pZzHFYF1/O3zXrVy5JPeCYvJf9o0OJYhQrS
B1HzHGf1uPJOCJoXN2bUCm8oAZnMhQhurOsNNnUPbS4nr7nONPRZlYiazVVC
YpfBlNIyYxdVt7MrVkt6pBmH6PX+un4irCZ8idOF/ovFD5rOXPOr9vuu9GLt
zjfMH89i53rPwakDZMQRJNEDQEe27DrYQLpb3kqylI5KPXEFM/T/yLMLz3i1
nyHpvMnZ9JPcX0epgNuGg8fkB7YAwxn48x/FNw+E/eYiHc4baoOZ686HBg9c
J+FHsOYb+DtZnASz0MMF/U0dA28IUu8jhPUvjofu5ADTiKzu++zOBsblQVHz
af5L4UirdL+d1NJVeIOViYaJqC6Je65mc4OHEQ3HMzszu8Nrbkg8NLoSaSol
+1VCL+N8IFp4INt3ODCWunjoptcMRL8h6d4A798dXWLDurguXp6B5QHOfQZy
b0cQsbg4lYJ5cJxHZqzdzmzsKzwN8dftwgTejLTzTtgECllspD22DbJuLymu
RIbo1TMhEgiP1LBQkzmEOif1VSnezkeW0RTnbY9KTwhtAYNGrK64tG6AFtyD
MKOyXxKDp6B1paoD0wtlZfWJpZxZZ7wrikhMcSMN93ewie5CHgIk7gv/9nwh
5Rzskfza4yMuvj1hf7CGjBLBtK961fc5Iw1rOQp0A0zSq8ZJmiucSmF/Ng4K
+SHJL5xU8qGCgUCVQEJVEBBf01amctziOC+tgaAP7bIC/++K59L7vhwdzV1f
bU2gcIow8Rdit3AHzfUT4+xCi+KX8BNe0bLAMAiTKfZhkgYBprr8nhEaZ1j6
JOsv9opMImdBT6jbY/sjLARF9NGadaayNY6zO2abHzp4KqYhSwM9P21dLbrw
qbgnowstRBBKHjhU71WIuOQwt4yjQZKxclUO+xylKE+7it9Mq0frkJanmy8H
i7IQajgAJqy5V8zSPKUL5Tjzdy690y87b1AGCjrDOIPfRIalKXlFmfmy289w
PWFelCCjtz9RS4li86ShjTSMZlXJiWRcaYEdPv4Sj5Ifc9k1ZIJM+yUOJDSo
kM5FQQl9iIWnxgSlWbzeOY50cwj4K0s0AuK4H2g9TKDN7LFOfwlmv4UKn94b
s5SIAEg2m2AA4Mp2e0O3nkd0WO3++0L3l65B5y6/AQrIAVh+UEwRLzomI2lJ
6r9wh0uZug/0DjV6I0kadcyAdxFmwDVGTijATsKgyrR8zwzb8KD0ePFo4bkH
a8via9lxynUtzU5PhUIj5X7S0XVfptuIHJk7JlfgBmkermwxaDQn9xwQRLRG
8b4GP55Zh4VvI8yAeXcDcZSsxZ4z2xqIsAhGDedLkPvqzgLKf6EyJdaNDzSm
K6hFijYd/xp4mb8igidyVenYuwrBMmxWY2saSMCeOHrq/wGgbgKSSrcTEKxp
4HrzTRSTBnDg5gPOjevWbcSt3hVA/P2NGYeirSZdeq8eo5O4ec0/6haib5Uk
ok1xVrLz8g+McIEBYXxZECD8kWFK0qM8hhaI+OQfJAuRpvobq21jyun6XAUT
dq6X3pmn4KcZgAFpyTzMEOpaIe+I1MIAX/Tut3kpWtjVjZRDAof3BE9SEIbb
5lAoPf9p/kMz3fUF1EK9l4BfDJUlP/ziMm9uwjApJO9QG1800+uVXO6TzrGP
zKEfK2zDJjnBE08hMP1GGWHeiAt0KGsuGaIMUJ2s9AiPMMcYUFxVCfWMDWU1
dpK45MKfg/8Qgn7yIR+yh3W2X0WOlgqjn/XF/vzB6Ro2P/HimTm9wZ+UyKk0
mkAAQnpG184nkvqrgcu90u4CKJI+kjaOzQnhOwFM2hnTMAYzR1RKzCLurybe
8C722M6yOYk41MDZwTzBBSO0M9C8l7yVxZXmUfH2uH3ZNqqDMCiIOpgRPDwh
014TMVj6AwNQKcvx1vKeMfR2o72ku3EopewEWol1IENSmGTJ7WVv9uyNXsQJ
9sm7ngMBbdqEck7t8JOfv/rbNC6fgwHlSQLTzE6qdKhn3yAb8zadmXB7gLDW
WD/52XVWWXeulZgDdf80no3sqhGC5DNWL03R1EvChYBO1GvDfoezRqZraRoL
VdoCRX+wh5fOd/jDOVJA7lC69dwRmLxuUy+9tBCRJiweI+eO9K8hIqLeZUhc
PUzmR+uOfldXSkf4U5+yxnhuyY+x1t74HphiO8L/djz8mTTLEt8KwEpZM+vo
P72E+EmqhbLL3553aJ+mmMJa4dh0LMjNsR7Du/p4sS6HWkNlZqK4yDLT2jeb
21PftdLKz2cfr4XkLt3yreRtvZmVfDzoaFQO87CNu+HqRg49axb8fn7lVIzk
mO4NvE72Cziom9xULAFZ1jA2hAu2qAoJao7uShbpN7jb8B2XBIvhbR3pq/Lu
YXCjfSkle2rn1NGPPRVxB7+v6KuD/ooYQ4DCVJPxBb+rE/zz0L1q40DMnGpA
n5v4J6WuKP+qIu+KUkNTplVs/eS37BMYQ639+OPUzgB+u5RtFILtHFlthUEn
IlKHtWQwZThjDqQ4SyLUnWlOq/OEGeuWTs9YAP/43IWDiDaf9WHC/Q68/b5G
yekouOxooquKsiuS7uMcwbhxHILyOl/G6Iygr18b0DfGTQOxIjjAKI50PJBQ
dmwMmrSmkva6hk/eftLnLQwta/GjeZlqLlMYf4dWiznfpnRbJSjiWOx6S2Pi
tkx8LuLEqN7e/XzrCaCpkrI94+2NY2wGw/1WfwlAnhtBSYqkLB/XxrFSRjei
oBd9HXD40dYV4BNh73Ag3VSyD0ufky9g5+Ovd7b/6KgY6BKMaTEg1z6SyzZJ
rb3yMtJVsmywONV1DnT7LHDb+Aoqr0gQ35WQSzuvTMsHWkeRTg42sCejGIDB
sBJYn8U4EE8S64VBgwFGP3rGsXTztzuMWrS1qLpwQhsV9IWB4xJflSQWBqZd
6CYXk9Xfsjlql5HrzGXzwQslVX5ja3RCa3eL+Qt6nX5v2Bwc71GVRNztM8ts
Bjy7ypJnAzm4D6A2qavRNS/11RHXu2372HhathdLLvff/fIS7gbI8oEh2aXl
eb1HHuj+Piv+SbkXhQktaiJIQ+TIfnWsmbW89nJKgDHMw7NljfqGsMEjlqu/
FzYXuvZ66aUgi2eQZWAs5x5yZ9UQ2lD509QIT7wV6N9fSOrqtr7enJI4NhXr
pldr3T/0+R84/NsbtX559jy57Eonyduzs01lOZvtRf2njhFRuHXP1lFQ8W/Y
Mm0JVF7yGpWUPdNQL23ZNTXdivyoBC0S0bTxnYHmpqhGhFks3n6ybRkqb9zs
TzgbnnIxPjc9gY3TS+Io2ny/DFssiM110PMVVYsH9E+JK7mL330vtE12pAUb
fAUJTKOo+DTak3ilMeXOj3qemRpz60UNUMpGiUCVfGeWF44u2ziTEk8pJqfA
/ujtwYYcSPW6ZGgnOSUf1mZHYntBaGfca9M1o0hNdoUyIc9zjiPV5p3Cz4ZF
1eZhFf4k3ZpuUFBsHCR5cj3g5jUzpiEnNdMrGLk3FUf6aWqZ1y+jE2oEhR50
AfYOv8+Pj9chMWeavfXbIX8qbbT+EyhgRvW2swdXf7jbgLWirPLon+DqSLDv
OrePIWTI7upSyToclaQye6A59Fy/vNu2LG4pq6ngMkeqMZEqHRfvGuTiVeVK
cUmZa4UK0WY/feUIgwr6kgnMdW8DMpZD/8CKggy/O0odfCeyxgDOsqyh87Cf
rTHKcaOekZTiHWjKZvkYTMhvNAd0FuvzKUIhAqnz7FiLRCMpFd65mz3YI2vk
uFRsfO4X83L2Zpvlg9FcRa8425WTjTnLquyLiakHMG533c3LFISm+HCRHfQs
b7hRFNNXobQXIrmG/HaL6NtWmffcVOXXij6UL83ZznAuf9cVzx5K8ZfNJnK1
z8NzgfXAmq6xXOxeXHUluhxj77y2dVYW6uzvB4rmiY0TENYMkcNM7hw/tiM5
TO5C3Ylt68cHg8bwyMK9rTILI/F+lALPnHeEz5dMDpgZJ8b3jz5/pypxV9gM
6P+ly8YTHacukwYcejQ3xh3LD78C4wVQ7BmNbs2RAbFc6A/3vh7rsQwECQG2
cXX9xW9+dP2bu9VVATjA8zknzJwqflP0fXgJ0dBG+uyWtepFC8GnIaX10aRL
mgcyQ93hGOddtCl9jC0cMj73o++OG/k9rUk/z1WhoHpEVczDKSf8EF9JWHTN
xgmSQ78KCJflMwIzib9s3ALRBysHLdZni6Bd9jXqeAC+08pGbdO1Q21nUTtH
PemRP9/0BOn/m96PygS8Du2KDs/Cj0QMIMviP5OaaqvhFa6Q7HzSeYfofl+w
NLABfa9Q5J4BVeWlC892cqiH4l90UhzBLAcPEAVE1xP2GbXeTKUwbnFWJOtX
i09IQpfxLvc1JrcF/+n4jJB8wPy5xs1GdWwlJtg5SpMPhSnk9LVhFTwRdjfY
UbH/q4ZFLdLj6b9YQJIbagF5ms3KRZMquMLZZVkmY0vgo9D2nc1CZY2ctGRK
QQI2AKCWe1cVNhWWGhIDE15nep9qXFl5X7/G5GHtUA9u5kx+SLMyJnbyybhR
+xJ6e7ANixZCb4CJrfM/SlT6h9bVkSNq/AaWwIzBf6PrsZPFcFXq/qghFvZ9
o/gcViQrdsvB9tk/wBPmzd2zf4HXOIpNL5qbukfrylNZwVXejizVfYAqng0U
z4STWccIq80hmPUVTptFssFhGRDMJ564ivqhTrViD1Q1OVg4zfynjnaT3v3m
WecH50Avy/V/0ph86nv07B7i1riGLEUwLqOPSJIxaFCGcPZOX7fqdfF+gPGS
u2RoOPdaaqHZEG6WqoRuarsqT3qxofUST+eYRwqjH5EfJMmTLnmmL9W3oC3J
ELG2bp0lxFXSDwShhJBJYMjjC7YVNLkypaQVdHx/oj0IvFaMhYZbAWJVI1q3
OOuGR24etnjx7HmVWi1Zq/MOJUYBhjc4r+xux12160q9/riAwIhCBNXVK2ca
ZjjK3wjZGAXqcu16bUXaX9LI3d23PDnGqydNcLWoHqLOz+g8vZ5QCa7mxrkL
SbMNHgQ7ih6PrzBHFSCyUr92RK4Px2g861Kff62pqDxwS3pkic1REEKRd0C7
VPajDJH28YRWwkMplJCgae5vXRAEW17JjWiH3z0yrQZhLkWWSfEx/bMMMJ3v
Y1T+rawIRa+cpRTKSakeHOA2TzsoLOGsqZngRJy86o+BZYhT3HbswGPwmvtQ
KtaMz14nfmPyUOpvGmn5mLe0gh/qgUM7pJByCiZkkE1gfP2mK2k/BzgMnxgR
vaTLk/D2T9IUtGi0X2x+harFS83I1m/J5agBb1EWEAtIa4hcgAR5DsP9eO+p
nAg4KEkOgXj2uQJTfwIng87eJGTsDpGSGnbXx+cgpeVoGM6XFeiuP4dEfTTx
T8IhdcnJ3bvW0+7G/0b1tHkJNufcY3aGhjV81ozrenXmKoqHRdFbWx0M4+5O
5X3g1pnivtFsVQWZY4Np24H1RVpHuCEeMytgGRgjQ07APqLxCw/N8xir8gHo
katj7So6UdZJJmRIPoj3eD7eoxuuooM8rfy8Pu6Ht7bn1Eh28tklECCF6zWR
KeBm6zPjVoiBWA7rrQR0+CZ4qWj+wgpNZ/B6WfqKRr65JjcSkWUrVF1hOe0H
+zjaMQ6sm+UKAINyRX/6aTWea1rXRuC3r6+GuqnKzVZBOCOWY+WPj+dWvoe8
PPOug2xBVDVD8WkdVvhT09Gwb3Pv3d7u365HHH+lrjh31GpzjZgPKmR1KSfp
NsgeAkisn5UFfrIz9fL9wDjnSL3dxqKVczRSZNBwNPKpwK+fvTUu0Q22WnDd
wb0XAjiRlXF9J7qZ5305h6+zrWMuy6r2QAV7D0qxb74YkB3K86pC9lAMf7rx
z6zFXHBAbHauu7oaZvXsToQTsshhzbcLGhQkxJTk8ii42Q6HCp0N8Lo4MfYO
eoRfw57KXq3HbCwejRZO4Yv6N9K/iUjH5QYo+yOHJgj/CHOnpRL6FMwcVNNp
IcahDOfzn2yf+Gr/I5DvDV4Tl3LmVxpjduYDarurLmuuX5Iv/+XsK7WUNTHM
cvI7aXB05mvVmRphjEIA9MgUic+QxmGrhRwrP952aD2Mdyx3gr4Y9aDqmqKE
k7TpYAeK3m5RQeBpqq0pCzXIffzfZ6L8hykFzrkxiicZeE2TPKqIZqWhedJm
W7Y7vt21ElZ0RH/9oek85SLjy6YaXApg4WT/bTRFDI3xQEqx9PKS5t+DCGvJ
/DoCvf24XKCUY3djIx+XA+2EnVtV1faKpYZrY6BbrbD3pBfunZlWOz8DaJkD
RYvSBRgXYHk6wgBhz/UJ/OVumdRFgAG+0Gt3lpVv9OZFwXorYbG0i3GY9AJv
WBbuxyloVMfJn+vv/qFRLhuNG6hMgo1KIxFRNqOxBu2bN4UJDG0T3MrGp1ZR
XuN39kWAKSBLFLlOTu5yEFVU29SshTEUw9YlvbDXw9Q6t2Kmm9UJtFymP72I
TBVKHxdkvHpAjOceJ2Cf0BNjEBF0YCbdE/vVzXGvNuilt/yA9J4+V3SIlOC9
wezwcVTbQz7vYkQ+UvDLVDkV99OoAPtBt/aS8pzscBjD8X0AbZPohc1L5B/b
QXIB/VQ3tK2l4XRF68jJRLy1NyhZK4GrRrTOyPxFSHzjDx3VjpXmjCzLpYW3
pFX6Xz/Ii2Ci0RCL9XukL5c+U9VUfS4/KS+3sZ/iyjjgcaz0L0pRNJPH6LHX
hAli7/3oT9ceks+z7eGwYMjXTHQO24Bw4X+enYC9iNDdhKkYX5NRFelCNkEc
CMAwa5IlRf3Pt/epynRAWKxsPK6tfHvxDVtOh4uO0L9oBxLbBYH8qm5BZ5qX
Rgk+cxlbZW1+Un/EIRRwoRsOTyu9sN71WzRan/JVh3jGjY42SA2zWa4hADpe
gf0guzD7Az5Awb5SgRZfMPvEfoFGtXUWJHGkldqXA9vJ+bnt0F7T7rZY5qVH
pqQAXMsYFqxKeavf8kjfvbtUs8LERWMv402GLHP09ztpvMbJJf7L3nPVV2cS
UN0l/lf/J/hZ7Aig3eYWBhsmVcgSooRXeNjUOrINPaA6/9SxPUXnyEK3K0SY
kCEyEobLN8V8hwe1pi2y8cJe/ZTTNPwPouKUGdebIFuUVvlYYQCKP93x+Q5H
3ElCoeKD67RX3SuVLek7ZM+Z7VWIzEkH8fEYpml7ZWd2IoiibI8DUdf6rmpb
TqhXIYBYht/OtAqK4KYfmtvF2Gi9/s6V7WmrG5Z/Y5p6gw/PJobel/7A2eez
v/ZPAVItr8LbzYkBJ3s/I/6hdocRDaMpHozAZDFBMP+kHmwAbo/qfRxPUxXO
g2svbUK6+NjLt/9NqpkIUPFpejl2nAYhFGaOep3BfhXZyJRX7b+zgQnEVyPj
rMXfBmDbSH1CnY83b58bGm+NCRYZ+c+aVeed0oyDZUpvwCK2ibzwH7uMlPnl
vH0EGh5kYs4zUS7Eb1AbukuNtyFevc2KWRPwgNjuTrmeH+NOfGLsOLCs3Xxw
03yjyKMLhMsBTnNNPyfxLIdvd6b8P/BN7rP2baPSbGKldW0LwI7cq0oCAMhX
xcua94l6F96iOO5esHFCsyyTF2qFb8Ay/QFejZGjdQ3VfYMWWEnJbWnog1EG
RlcnedhW6K8tmkuDN5SwL6692uPtCLPLT0B5SuDQXlgKjCenWGFLMYwQ5ubj
hdtNdxD4tHY7WxzO/XahcIeANSPad+gDO2Yd0Gn0/hwGJ9v17i3DrJDjviGF
jrlVp++62zD9pNqfrIkZu5P8j38bfg0n7aDSqI+9jb9NU08SsnW87ePKZKy3
dLcdfCh2MuFB1am3zlSmDQwEBRrTSyCLW/vBddkUHQu7yX1ytH8imRwNj1Wl
ZFqf58KJrwvkQ9h+UOhd03OlruL59tpB5Cfb49yygDZowTzmWcSaXYkWrK9W
zgwmiKi+ARgQiSVcXhuzSANrhJZ0tfSS6d2NBtRPhYdDIgrikrNMB67g2fat
23GjSlc26PFiFjjoxV7QR456GtVR7J4FQhVTH8BYSjckAB1laA204qtyOklv
P3i5rKss9PwkzFQZo9Wdt8XIgde64S4KFScr/6OGO24425DvAGqz0jJbhC0i
/t5+Py8cmmakWAshPfgTAg6gk08kz79gVuyXtOrR04H5eUvfQDHSb8oXZIXO
PfehyDsM+tiZkTPOb5xi31ML50zhUzQXAJws9BpHC0IIu97SX0LnDhMo8K7F
v5bqS0uf6fmwa0tI5Kmr7OvTpzW6XBIIM/pQXv6njUAL895cq6BWDPPWRb9i
W5Lqg9vfk6RFi/Wx8PWZ3I8iL1IhZLUBz3Y3Jt4bnlcnvX9X1RGiiOJKfT43
qS/wpRxnPsnqb3/L8lwQz0b5AknIpcqxCJ0Lko9+l/6X7K0trSeaWkPbZZCS
7B3d8QiIB8iwzL3IRPAeqePpHWsDwZslMDTPdh2jshOpRyI3W6kXewXmUGrc
+TRTU96PRXcv0jFs5J5igxVOg0kAZRNnxt6yCbMjcsbQjvAYd7f+Z5wFz0Ux
YCG7mf2D/I4+d9sEy5MCBNsdqYTK23od57FGh3i6wOKfcS+i4yoOFBlowQmb
zW9KpqOeNlBwZuJ6gWFtpdRsyaw8bVhfx7nzQWFFc6hjFiBj+2NAY2ZXceaF
7eS+shE3S3tP+8ax25bvOhpphTo3WqLaG/0gHgMGrOPEQeOd7xjAvmJw3TvA
BxwEocIM97RtL6cVFChiVqkHp4HG+XwjR6MhB9EAOaEEhFhQ+Al+NLS4d7HW
6BgCCoBDOMCk2m/wz6kL2q4EKY6pr4/ZboipTrT8oWBjwEUmRCTlSLbD+KjN
It7R1a5rCMCeuhz1ZwewvZpsPuJZay2U31t5cvlFt+Sq4TM6mYlBk879LVis
a21qIQ5GXW788usRLCSZueuqsIm/4ndZyB2GTvlJNqIwhUM450/TDKasAD6I
+Pg7+gagQev33CTKmoW6/rCO2QYgTvJsuYcgzMVdRbXVWKfID0cd0HdqYwPN
SFEcAoOayKk2jkm76yJZ6OD+KAiXcqTuLC8Nyrem8HNCIq3Xud75GLgfXNbA
pDDbvJA29IcTT9XTlgtkJ+wdfJ8KNOOxLQY0jN7BVK/7IkzlHsz00Pe5n+zk
MgZ9ciVDey9wMielt/IKl0bonSV1zm8+DDJE935YSynrckWEqPZam4nmsXFf
npp7NgurPpyzbeK4oK1o/BVqlUVhkff1bhQRvgi6nzkpOhzBKlgSXvMoil2k
wgTxgQkystT9g3B1lyClqPa2KPOluncK/0pZJLBrnGaaq9ZkW+Cj1IqfIx35
yxzp+Kx1kQi60CPwm+9hDtB6vBoVab62uLMvO79HA1QSf8Fg6BbNEarCqxU4
SjgPZ1Y534ZFDUhLCIbZ2XIMcUglhvcEgwyknkAVeiE3s2rY7lVo4LLRAKFK
ktdKcwriB13+fmr0WaSwEW89khRDmYnPLBDQBw0cLLE3a8WJO+u+Mk9we78t
IQkggAWLQZQrFr1zUTrBF9FhfqESY+5pPjvsy/IBpBe6CIIkLOrJkqKaqAOS
jr1P3InLPiJDkpO2shG/lCqGAy677wv3FWm7l0qjHqV0IfxlLZYvOMJdcig/
ZyY+Gpc6lMpcWQqA+uGfSs9CTVR+fr/tf9HjEo14bxdl6BUoNGM9FnnTsMm2
y8WRn/r1fNTLXFcKS7d6R2ltleYjBMMiTF9XtkegojtF4EU3/BeHydoPtx8o
LkScCUREVKa7HnDaqazUDla8UkNadCcVy6tM0ch3/T4i/FIHMPCabJjhYWe8
IpxQ07c/LTW8inYGC/NfDLr/xoZu9DkwoCEyhPTQrsj4cmk1clXRew7X6YQz
5qED86/d71FSmxBYoXHrGomUA4/p6ryo3VedL7PkgAHgiya4azP4Ifio9Qxn
5EftUhI88tVoYZuQEuvtBVstEPYR34MLtXuuu3q/6vHcVqOnc9RYyvwEolIy
nAiEO4aSzyzu7ANLVQrDd6aBwVQkune7VXu39UhS6R3xqx5+ceIfMoRWhI8N
U09xl4GywF5RHx5hSzYrvjpaVRVbpi3VWSrQIzM3isHjwXQFn+eN0IsKrBik
30BDCY9ButTOrvBh/hd+jEBpnA/l5w1mh21sEismYFMT0X4Y91uyPF+r8FpL
QNApvyQy27wAKrQlHMswrW3psn1r0QYpiycWOhoWgM4YxLasoMfza/tLFX38
Y8gCJa6cVRwywLTuOx6bP+Kmw4nNp1RWMQmRXJV4CaLlRq5iyDNizYxQnw4b
ZztHAhKv3MBZW1ZajMfLQ9sobIqJI5vgV1PUJBbldapGi/RZhdeN7nqFhe4D
46k7mjXW3kM6JcfyBcTEe8iT1FOitM6+YfznHPh3FdoSiPKM6oUJMYBGI9I0
QvMqMP2NDyRoTSJEiUUTph+pFBj2+lRdkTszyR/dLOsy5Nflh3GfKFHXCtcS
rTgmUPcir7kp0BumOukb+bui5X/LkB4fkn2xhZuwKB51cMKgjb2mnknWRhZQ
rIJPfasg22OMeO/bHfzTjiru6NHXaL2n8v0d8uR3jdMuUvm3VBMMjOflsdvY
d8mPNn4drcJOyQZtFi7HZjsQ2qjc+pwD5TsK1P6umzEfJlwoZe1LCmnJNu3C
/p8nYkOz5kw5RnhsIougFUw6v5vfcQgihMTzdvrhRVP0zVAFjojeOGEhXXdJ
P/tRKStHDI/R29uL33S5sgJtp2BCZ8OUffsZTaCyPNIoh/SHcKQylBWsZllZ
lKCRT7XwtcGHEAdZC7xXW+fRqGIPnOfottr9M9tay4YXOE97KX0HfkK81C6G
cKKx//JgoRh7vNaRPD6bjYxnrKX9zH3pWXLwzmSukWr9+zZeZv+XRr1AgYI2
oX5B2SMUI3Ywd2WwBb2ZC25lB5ErTHI95dTbtCnHa/Jz8cGYpXshN5GxOZfO
INoGbc7SpgHDEoOCcff/I9lZYyEkAD36teA58SPXWrMbJFN6LY+kGdr8tMPO
yf52Kk2UrPnROrPGaOjZa64uzp9ew5orI6RPGCaTDxO14Og7NZOhV7nQY0T/
MxqEEOzlovW+xl7us2pokrHQy3cAXgjq+6ojT5Da2Lrjmq180330jAiuLUR2
Dby4osjcKjVoVb8IN2ApCWEem3VxB8yAcA0o6++paxXNC2MOsJqI03+qla0v
Yn+WAIyxFly6stRKdx0hB/EZZOnzlhSkk6zhDdbyhvTTxm/w1iFNatqrllSI
I7T3h3YX/90A5CU50xbg/+t3q0BWdAErQurFtrN+JnnQM/CspzTYbx0aBZwq
bPSSiTEdq/0/KychHmhP4fyFmiLeUHS5O/YFES1X55sFNxY4hm1aa7XaIpYo
2LaFK5K821sSUxxLqJB12svV4TPy0Y9AVYHYLYSDy06QoxQQj9QYQsrZABBd
Q4PMnRoHOEZ3snya3vcdAh83Ah58fi2nmd8Y4xpq3F3TynYOJRuB8enb1gTX
zDoBOVGYj5KBx7KF8k8iPsR/jnKMMWPBBBykZ/3bB+d4ba94HYvRcwogyxwi
xQFlIz/c1+phySlf59XnHtDLfVH7LtbYfR0TFJzGv6kOdeDYcZTzPg1XRpRD
Wo3Eh+U3kJcztjQqI5xlYgR1UnrYpS7NXF0ubNNw9IH4/cneWpHdE87iKWU+
CZJj2dxJsmgfhl15d0FcWILUSx2XcNLuXXanrAw4TuIMjNmIBd/u7oKfTgO6
TdODLBwpqlavdvnUoVxSZHOCazBNlU7c8XbV+coE7+70FLTsPnSR0yP+FbbU
OeQ1Ps8Lg+/VAn2THhKobmMjfUxuw5V5l5+cfXD/GhE6nV2PpF3MgUWCoHUR
KTF99VnbBT3L5WFFoIZHQSq1tZt+jbYuMMPB4gR5l1Z9HjHfaHUwOYPUEF1h
mZn1zp9HlUAAaus0IlgNOMsis0cClfo/l1AG89BkxtU8Ouzq0HN+I/5MGSwh
cXqAVrBHv4dIM7LL5aPIu8/xfu5adnSiT/t2CnUpBvisNvGYh4CXfyF5wRlM
IybOhRh+jszQdA1FIyT6xMSFZETDOR+ifVgcboAgzyIBaQzjkPIKj4igCgHf
hDrr+vzV03k1H4BmsnPTd8mmDJYzWG3bDbb600O+eSJuf7nI/IvwtVgN2rZ8
k3A0Q5V4o2wIlkaNsLJWGz4z50VhlRk8qOTj4EvUeurJbTK53yXneTABPVHT
R7SiiRTCzjaIDLl7+147DCNK5eTGCzxlMVUHJITrD7ANEtX73Fh2rgBQhcSs
OdR5EhbU/e2LiLoeF4AUAFUr71pxomN1XOFA0GQZws7kjdqOJwLEjN7GE1E6
dOl7tskc5b5fTBCIikhxc6ijHaRbkRTWGdWelVAOZL9yFycZ/rJDcYSjrGvm
KTeafN1ai5D1Y0hKKIpIZRFYPl9t7C9J4vlgHux9WMFny33U/1N0bzoww3MI
C2OO2aJBeY3vqY3g5ALfCSghBh6f3a4FOIxIqh5EkOwJL0re4/ec7+/ftfPd
1QTe3KLpKgvvRjRTmUpcSXXEJ2uUSOjhP5riUGJerJHnTOhNnXvmS/eFyUxV
zw3lfsSAKCbsXA+PiLF0cb3o59RjDz+Am+CiYnYULIav3Y7OWvTGLD7PmGms
3AD3s1lgweCLHNkot9TpS2hT7/o8EfpfpRRGXTsV1prkBoWTdy3EOUxnBUwh
yWblluBbPyjbvAqfph9DbLKWn73QmGyDI/ZoT27ZV02hdEBTmFl8WQzxCfD/
lj/iuE5SNsTfYLkGiRjB9o0iuqvUvais/a8dWesa/tAW/qlUPkYzfBj2COst
yGld4V3VPZj9nxtye8SENR3sFOR0YwFGfIX9P1kfI64UsvtczApiX+RoGDD1
OZC8AF1sI7w35OzXVTRPD8aw1OK2UdvQg43vPS1SVy36MRrV6Idghu6w6GcY
0a5Vn52nM+r42GSQ6LhXLZBNolXygTbdpm4bV3EWqA+cW05t9IURtkExGWAw
xZPS9uOU7R3HWrmjiF6xBskuHyHtsPCVlUeO67TRIZyoe1/UEJ28GdLosmzk
TNWnJRp7DtbEzGyo76CUDWjGKssW6846ugVETQVK2rClx59eb/eTNLKP5Jzs
HpTJNQheg4pvGNhNQ29sMQS+BouId+D2G+vZjEyAJLk6XoZC1lut7Uqs1U0u
QYRMVDqfsfDDsuDjnfzq+JCwHQPIHh/hbaEvtxB2Qsqyc/P2Mh8/TlUCXgtt
SXHBSk+kgFx76hSR9wWYVLUfjtGrBtklQUMlOK8W8julm0mePqRcImH/xicH
0DbpKY5xMFBaj3Gu/+tGWU0hREZvgxjA0BmCYK73RQ1cihiR2G8eod+p3hZq
k+o1vnF/ST1onCIx9CFMelNEZoHS839uGcrr4uLrPjmV9jx4AQtqPpdkqif1
kTmh9ftJygHxa9pV9vFRZKFkOjZkG+siGx2B7acopzb8HW3gweQQjAkHccXK
4Z3VnTKpu+v7CDkpojNr78MDiYJSlZwVyjXl6x2l4PYW6VAjvI4O8nAPf69A
gjw48uxcXgqgOILssjxQyXgpXtcxK1hD3JXcmjZ8iRncI7OIdPyQO9wHhTjl
tmz4BP9LEHNPwrxN2rxLGSrHsz7LF8wnLvZVW2EdD2mTZsno/vHl77nffGP7
gBG/EoAh0sTt7KW7AZppUiNHzBjUkDoDs+Q4EZbmb7psYbGLkaaL+IYUbAgf
ZTcHJE9ddJOWgYOXKGtcblm+y6TDAFKOGO53JtPzX+zUlezwacfJGhz5x4/4
yvpuMnoD22Om39dgC7IAbATLl7LB0vOQgKtbbaAm5S9A/W09CW/jB4eeroli
KSdTdamFvlb1ZKmxH2i1Y98qec/XzpvzskGRWH4I6q35Uz+yflVNuubBU4ho
l5Pu//cIS7KMfa9bhkUVS6cO5xAzulR0Dj0luzd7yXEz3tYLcVfPKj4kXbJK
w1Cz7yre0BPRFnTkrwKIAUHPharHBUutoS8dlwTzqfweDRSRkVq1DmXxB6Jn
gVVJIN/JKvRtq/B7UxaiG4kWZmOzkksctn1JBprZXuOuh+hHp6rw/+41ZQEN
rl+rHciKu91qmVnY+tP2/d+ur8qoPy7xX/zA9uy5SEiHU8vYZlWXm4k3xvCX
ny6so8L22q5s/2BMUukLWuuuzbbIQXTeQksVAEQMkv6xyXACyoajGVT+P6eS
QqEcGwZEPGLsw9wxRAnYSz4XpgZvoaoG9gJfzsImpJ0Qj9cWxDGaCV8Keego
NHJpA3BUp9fUhqYuaZVd1A3Uy03vS2uQoy+u8xPZbPO8CZQogBFxDQuADNe5
PzZpEnhvAtnpMrxWm8zZVGQMucSK3fuVFMlV9rW1eZW6fAv+d4ANWofFCcpJ
jSoCx3YhJ70vhhVmrJMjLgqyNeMagwEBX/Q2XsmbAWnsdbwaXCGpjRNwdzfr
pe3rOOUviv4lwoEGcpz9lDYCdvWcg1UBHnysb9F0JC1oXQa9SNZqlbo1v68t
yV48hpmv68Gq+C1ZpBiMeMt7KZLg7HkjJxut7PUmvobsuynTj0gXQf8AnM5E
vMv64Hm2btQB/us17hsqJOQXVx/5QENP2gztLiuI+mCb3Yn5Ro4zia6nzpTI
jkCSPB6EuIqWoFDV4ttU/y9yX8M05bONs67ZorAT0EGPay9uqszpx562fxZl
GyWH4R98R58OasbYHwJ7FYhbzdNG9GH7Gin1iQ1I/dezyXLZBqML6GjIqqyi
QRPHmHhNjS7TZ0EkhOmEjbSBGV/eMsaibR6KPJkSMyk/m0+iQrQ3ibdZS0rt
TqlSbpz9FLpwiX1sV/G/kr/SrooREo2YIPXPh38OA2z/oVu3QCl9nSM2hm+F
YUd5+AgBJw9O095MNHYa2fr2D32tVgXujaEHDbBG+CiYQOox/631y6VCr9xH
C/E4ghxuvyX0fz/IWEmyvr7ltS8w4Bm+1N0HCVGmGYePuxUVGYg0xh7Hysvt
BDQN9HxRS09CB0NH1Dk2749uNIyjpWAO0vNI6cjvUHlLRXlKJF8v6XI/TbIL
U7X80ZUEZVN7yxMy3051C65ao0AiZlu86A5/vYJzd0SPLnu5Leus2pF4Lpsi
OCDlxkbvevn7IFirDpS4CZj6Wh7tCN0iNrBH4R5gFnNdcTy+PvGXl8h3uXxk
v8nkrGizFJ+3pBe8a/QVEwRCVD9t7ivzK2Y36TUjaZsInM79QuejLVKiX631
12xyJRSYAVTJZbYnHgbi59nWF9C66XYcxxVrSweWUzzzabugsWjQhVIvsdzt
kX+cN9ke3KvQMur49+z7SpoNxAGXJJ/rd9Qjt663SWaOo95tr5//m/Gj7mkp
D+MN0X9ENaxTnLKhNi42v87JdfA/FRLvs/ovNcKF/cDwmvuBkPlRQ57bS2ul
KnhoDYPCKzZI1RaNpI767zJi/PWvxGgVhRL19MeD/QeJCs35loCrCQyJk6ds
6yDGXqdq0nsdZbCfCa++kpPMiFAtGIyDaHJn5E8vPqwa2k/dLHaXOy70Lovd
PDvFXgEQeDVMckkbBTwCCcVcLsNcX+6gqu55/ZaLs96PH+keCm2eOoT/6Xek
Ux2y9z1kQbsU5yczbp9ZdDivHSCckG5bvU2GiQNM2KXt4ybcmUIrkEJyny/y
KD22t1IzCnvQW7utAhL0Z6UOd22rWOuyolCdd6G4rPOeux9lJ6+qbFrYqpZU
776SEj6wVPOSOz+gnjxDB9VQ0GwN/UKNSrKBD17DkX8oWVWA7aKvsJKBSFZK
B0o2kpIwe7n1xevtY53W9t6SQ/vzoOxOTSxZRuJRVewOFhJH+ma/dUiY5y4F
2R6IN8Z0hKcNmaO+vIKzEeyFe9cvd8Ub8sE/XauI+oFaik/rJozP2WxjHq3+
1jNYYCOztGPrU3K/281uEXyt5uEfTgt3FyqW/vqGYRLVCC03yTzRuZCgbBN3
tsSC/n+BmLcIjhMNiPLaYaAXUJucDw8WH37zs8uB0DvtWoz+hqswvblMe3n+
Fw3Ro7oUf2GPteEQX2TfNNBpuQzBqSbHbUiXFFdqeaX7XklbUp4PAbaE41/x
0aUuzniNCgNOjjWt+UhJeD6E0hmlrtWFlvbFxsVvnetCU2q5zhxc6K7r9UBi
XoqFRygq/clOye0CcFQLG+h+xg/KoEFaWhSprJknA9a1ze0EUvQ9EYc822hn
sczw1Iwtp6aef85FEgq84IwIA7ux4RVw9B+qnY9FFNO3LchMOgR2Np11FV4G
gtMIp4d/1MFvGr2kCPFjawpgbzDzD2PyybUIaOxWmDoev0Mcsa1s3OoUoh4j
gYj2eMeVJ1WVVxPOATA5HA/qFkEzpDwi8D5otYQOafCVvrNDihGOPjzcVdnS
gQurLd3qgGa1GeUBleC89j7N3b3ACUjqh6AYkRWVzDBSMv/qcPSCNkUbM6yS
yQZpEg78x6QppoGdcKZERmeusnHrK7wdMZIxQAV8ik/YM+VkB234HnTx/au6
aeA3CfmmfN1KeIIIoJhTma3D6u5qCaBNZs98sKk8MNNIw4iaWvwPCepTBWs6
Qi2Q38JNAugTL11qWqYn70U4QOnZCu76SB7Juj2OzoqG0F06u+JXI4z7a0GN
X8aq8wX92aAqGuyD7lKa4XLrb96to888ppHeAest2RcvXz+BcOsvlCPKFLJU
mlPqe0SbDLGZuDnRPDGzuT9L38Bwhnt8/YMhJzlpP6FiC5SES82tSnYYesNe
vDf3iYIwOZjdDYx+npDMGsw9GUxsmOMY9WIPJIOP6rYqK0YcZ6X0g6Ow/V8x
FASOri+ltAh/mrqscUs02wxMLcV89GfnQ1zMu3GcKqj8Shg/T64/0zl3Upjk
9d5NyDWfW7JS2hV/s7Wl5GBoSPI7tXZEG6eofQA4wQL4CbGq/41wX1c3IOnU
a4Gm9/Qm5/whcM2IhqBpfbMYJd3fwpzhoSY4uq8stXS7PaGWa0haXb1tyd3u
6cP9t8o0pM3LWv7yAQv156nekw+duzz901qDd7noxK9wtLyGbrMZJ062UYir
+7c9Mnp3Ea1qYw08joow5o11FX1JnxKfzJIDhFnjVhtLXN0PkYBmEGxCe4Hz
2MSZWh3lvmcZeOCz/BoPIEs1Dc8ydkf1xHAWTtRY/nR09tZk9z5G3uOeYaxS
W7B7KjSQ8F6zMe9JbcylY+838SbqH6CDNkYZqnxjtjsT3EDtOYdyThYJhZUz
CBmbjuMEx5ixAd53JkAyHrEST+k7azWbNzeKxmkiGY+haIJh1Z+a7px3IobA
0z2Icybt0B7eXNT+s9DtZjkZJD8WcGzpfGijiceRbTsLi9sQOTbKT6iIpE/K
LxiQGyTMPlQXRiZIcBvZ2Nfgyg+LkU3F+3AHexQITQlVgTJzuvecNhAaXklX
9c3iprkc9YjeXbSLiC64Wb1efyisJJDBVz/73vSdAS31t7nJpGBX8s3GnMq/
Z5aZRRIzl9QBWyX6BhFF1bpazXAom3bXhVyGRXGUFjz+Uyh51POaczmGpYiR
lyX88k/I6G8hrrlfGW/fT5hyxxz/OKb54VptBOSgHQG3INcluyytJW2/lZwA
99dut0ohwSNkEG0KMXpdS5I3NUxJuO2LPNydzb8hXfLnyIxDcs5ePUicjaoT
CP6IISR2GexTPgJKfoC2WJieep+nt0wY++XC+1otDC3FOEwkc3xnHhfbBrHu
a6f8P7KzmOaSGn5GAHBFygGhbbBVgQm54tcD2U60yFf3dFsu1PGuH/b4Twok
2ABq57ryAAkabaTo3gMYP95cXEDmo0jmtX4wCgqDkNJ6H8VE5WZbw0evFxGL
kqvYr0R5guEoKmBLKVf2zUHDOHNMRosUj26Ki0vH/ka7tZdVQcXS2QhEEhuo
Iw/8C1sogshOMIyG/x0bRMjSqnaf+OAyB6Zj9zK/Pu5IERsXMvCWzIren2ja
XBtmMUybWLl2x8iawHMQy2fVbT/HsFOd9cR8XHvl/rtv5Dr1O83HzX1OpJHu
geo40S95fOS3VRC8erTQtLWdqsDFrmUk83avDB1jX6x3ACfSZHDspASciKQp
PVQgpvv3u48eI18HpdCVULUm3o1zKynI98J/i5LB80OWlNjcYNWZoWkZmxeG
0MlQ95o/tAXyEFNgyVRd9fsL+2D8vDgRs3Y7tHilLLP3JT0jBIcNw+Fa5e9t
1iQi7+Id7HlDgJRU0hHLIskXisrxx8qyUHOVFm3Ro/KaVzhiTE6hQR5JcgGs
oxtxDYlbds8CXkpPIlW47kYCoPuqNFekro78XAe/vOA0c8SqdKr0VYO8G1NK
nn0acbXxByLG1A9s5UI8RFaHKF4xH2r07myyyBFDgCYfiL+HVVfAsgChs1oC
K4FYpag43c4WoAdlQ/zmFVhTUTAvv7o9qeUB8vVjDg1q77y6JxuelJzOAOlN
+W5IkAJjDlYK+c/II+rrs9+4Nf1Fj/5Lj3/rcwDXbyOvNjzoi47I7N4gjJJ2
0tc02UowuO8asMvLWh0tTH2qlKTVIwKHM6HoQG21DOuqHcxWa9ckUZNTsGnp
C0+pUJWuirKWXPx1bGNEn+m8Td2XXBWKLLUxuy3Nb2W9jTEAFw5aagsVU9Ck
ICXyTIXbh6pTSjNWEDh5BWIxbuMCHPJ2IiG3fe0RVz7H4ZBvxTGdbTsB+Uyn
wL3B3Xfd2GXAvBPIaCgnIxDPdmf1e1EqfCCa5hxtWzTdMivG7flEmnSj+o6+
OFKKFJL76crbiD0HNZPoqJZ5j9dR0WXGZK/3h8tCFatlTtzqBSQvAfq+YT19
IvEajkGWAJjegnqfm4LnwPORWzA22ASb25nCF2LnjGLpd2NMgx/sduKeM5+L
GumgIK00enoV1IP1wyG84npfRT8KJbU2pMwQrfrWmdRExbnBPIMoS6LqwNJS
ugXR/RzQF+brouGv847v7POicnT2B7cwIGXPzyF61rMcvWnV+BvLQGmll4I/
c0Q3T7u1HCGXrBCCBLM6oidZQyXnoo+AIFhwgYjMc7yxXTQI1YTwFaqSFBmE
5XFlPLZPHVdpQ6G9rIA1TPQzBYPMpzRylpq73gQOTXRCZVwCUNImnUCAHG/V
Vp4oxZDe0aUM2/nEF4ZwLKDlHESWgWD9PnJINWA7ZW7uJHyxiQWwe5V9qITr
FLBleN+q14tAuys4T7MU7pjt9lrQQ8/io6nznbtKhLxsvOaLCTxr6hA6rGGt
oIu8p/C1KCafz5lKlswP4bBY0BGw3VwTkasbYy9zBrnM4C0OzAT6D1nG8i1n
2WvQiWSBBupST4MUr+2hRNLaMnD65+eOARUCT9OCGVOBHVFOQLcyA6lAxGD7
wFO2GxDg251tEdHKrZ7ZfS5dBXmlKU4tab1+PGtCL/VvqGaYkbax7NOFBb/z
CKn3gUdcvZLsVpalOc5ni7/7OtmLpoarX80uLaBVwUyNpgheY/QBRpfpRJXP
EJ0R3E+i7VvoVRtQ5bveAUjT6p4QocsljM73HWIJaBcnYELYiOKKFnkiYv8n
lulUNCUGdLjnYWdJiWJ6a4KZukC6bKnW3GehIO+9f6fMDPzpyMvuTm2ajoG/
dDDLpm3a5Wg1yxP/wX7tcgXnmqZHu/jysV6zMG7OGTyMulIGyA+23T02Mm0h
1dJ5sWTGO3PXIal3VoOeTUEOYIQoZmlHtMDT1f7Ob+ZHV9WHoo3hGSNzj1PB
m6/6QIM0eMbDS2lJxyFcqpV3YVq4MsYTKHWnSierCnEBq7uwdqNp0Rg7cOtj
6AY3jBV6SmWmY9jX6tmHR8irQN24OqHSeLMaIqMhx2AXHuWy5Qfy1lv+tYpt
E6J4obYEXArP73/8k6LsGCc9WUDHoeABeVvyngVS+opka13EOCc9VLiHZx4Y
DJwVCzd93ajEHVTgPwCCNqwYLR0n95NpbI71/WL/e6MLhflTuSKGZnDnLLXR
e7RqbEotjHnD4E3aEh6c1NFY+Rz67payXy3KyIMq+0GZ5xjMMj06F5b4GpYv
RQ1FssNw+zWsvz8Q8GmI+NwGEbCZNQ+Z6otDthbpUuBGN9pXnj6ApbTpJNeP
rvFpSVpD27ZqZgReFhms6HrTaON+34RCjLQLb6qyAPlTt1HI4w9wC0S2dMsl
GH6Al+NXMJpHsq9k8VCTjD/CkU6MhVSQoa7AELCY3D7gXohCe05BB+QTbU/C
l3ybkJLzfWgQ9+ez8PQ/GhagGuyQOWaH69lk+FT6WcIqRNQpp45bPB2FZW2C
+sY8IElEXUC6R69Ofdugz408KPI74uhGdDFPKgvqetxmgo72jwwzeOeyLclz
SkBNfhmCcQxpcOWtLjamtyhB7Jh1VepyhMkTCHwBslDCO+23rGnUgNdhhz2b
2QaMm8bKzVzXyqFYr14Zk8bwmLZuCP+lRU1RkPydzHnu6rKu8a2dJAabaup7
ZmBfbfi/doe30PiMq7LyfbAxQ6rQ/YwbmgivPHLru3mjZXpqylsL2QBVt3Es
54S0qg/ccTntJLqoPDqU9PT5/X27zRjJ1fe3QFQZvCDQ7JgSWx/x3oBHeWlS
i0MS0Ano5E5hRHecELQDRGSDj2QTiGNAvCqQ30/pdeGDCg2dMbOLK7VHKdjj
qUimQCtuwYC1aDxRE1tnuN+e/WsD5HJEvUwX3t70TIM25Kzsb51A0WQK6roa
ZSqjIJfC+5zeip6BNX8udiwC5HT2kGG/x4ebKZ/qG6iIHjypaMfEVp+3JYh6
V1TqLTy583r2972JbVX6Cbf/EAx3Boyj7myk2MzP3mOs0JTdtEwt07wZF8ld
fF1zVYiYWqAPdqPwO50+DExcFV5kenZlIFDlHYwNEdl1FW8PC8vHcxS/CZ/S
s0lBSY8GdUUFAWqtZQOVrxaxKZK5AVnbFxJ0T4IJ37McQUI2lNH8N9GqUON5
U1EY0eRkE7IQMOUhKloCwFk+gDNo5XLRUNdJn7k6n8FJ5MF4atuaPfHZMGO8
nKBNI0h+Q9sa/CexprPDdoQek/CTxROWEXsWq/1laQvmVSWR8ewNUZdaM1lf
4rOiO5NakNIJsQGnlr7OJnriCpxekdPBTZBHLXTQygQlHWyTeuIN5xsXwNlQ
S/HzfLguwXipVedo5Fawa++eFIWPf78Bg4mUEERWv7uoRz9Rh24yaC10PGHf
N3OXsr7DctVWri+AnRkWxR/Cn9zRnLJRKW7BgMYu0K+lGcRqAHQY0W9STm8v
zcE2oC5Wct0iKX/CHsczRycVWddSAM9YKQz7fkioNwRJJKw9Ad/eHXWDn7iu
G5kIZ+Fg1D9CYNZDbzFsI8uZwRCV7SUqRNPMhTwp1WGpJH/zPvjYL5Swi3WD
Wifm8SNV2NWvCSX7M27fg+vc5zVM/M2W1m/8ld+vcuu/unBjxdOiUX9j41/v
YxDIdpeTE0qw9Q/1ySN7S4gZ6XI3BJtYmOLLbHJiM87BPsGMircC5XnVXBS4
afBkz2inPB7Ovqz01kZvYuIbxRcNx1OhjFGmh3pZ7R04MVm52Zws+nT4imrC
UToPvWMWuS0pwU7457LgO4BtuJeo6veaQm8RhaqglHOf2ErYl1zy3UsAf9wP
uTblucxy6UbMPWotTbw+QCskj0+tvgym0BQXvgWPyxcp0yf72BAYbWL3pjEO
4Co2dRPgQo5CMB0uBXp9EGoheCD31aKD5JFGSKCxCOLggajeAYPof6POAVOc
4hJqgMAQNbFqrGQBNi4SSChP4RGxKJ40yv4Zc9PirrRTKdqxZFLywwAFyMtD
rBeFA+ujN+xVAbv6CLqFQsP+Q4sh32cRYOcfC5L31o9gSnodW1ibMuM8SskK
jk6FgXf3PTWCcKyVhI2KyMcB+MkOhD27E5zd5iAlJ6LlhLj1QQ0e8I9gIE9A
5z2Jrvrk6piI5rSPgyI1wpid+2Fx3Lj3jqjq+y7G4QZgmptMaiZLfWQJ1h34
p/JHWXuJfuVcClcpGyZtsRl3Y+5154YadDkkYpAUPd+Ga9ikxgq/yR2I2fUN
JOEYHy9xkH1jMuzGjCF5SdmGgnEaHZb7OIqGkZz494GycVamAimI0SZTO+n+
wCm9RPUZniQII3if2H0wkgXRvycLqTDsl9sy8gyRAz2A9OAg1rAmbPh7hT2j
VMEPTWbaUEmSQyI6SIaMen++oC8RFXn0jAszodMWIbDRjTWQlOOnvQ4a2PUD
tCuuilOBiZTZ2zhTbSZQU10XA6KCfTRUN6rSzArdlzlwHCaOHLQHR03qz4KR
d9u4jsxn5rDZ+PNiH6AwBBxpnuUgG7lwNcdN0AtD66Y9mgVOWNYVSAjr7adT
Nmx9c7URlY3OHr0XvUpHN9pVJralmb9nZykA7rDlU2LPVhXI2s0whUK5FIHB
lJ4FkTPdmlO5zSQMN41ioXb/xAlzb3714OpLOJe9ltPft8TMOaPmtFzwEN9b
h45fEQH7g9G+bPse3YisQIq+xcwAtOr4P3TBU5cFs4FXUSBYnwdiiTpDE4f0
Z5cJlZvWh7wMw0+dQ/yqssYAjrnhyOUHsZPnKwBRMGXdDBBNNkzB09N5yf6C
ctW4aNCWK6a1y+ZXviBp8y2ms17SR8gUTga6C0sxkT/6ceSFkhfn/cKT3ctN
ONMCAaH9ezMQJKx/0AHYhzIVKW2U02BVIB0eIfkQUEC4e/IwqcUyILQUn1ok
YyowRkzvD0BHhf9eAqCqkWNGe0YbA0FHN0ct6m9Tl373Yd7nxzm271jStOFG
7VgnKs2lCb2/W/DbseqCjAveD/j3zfA0MmQA/xq8uG/Tf5uMqDGOADC5I1MW
eiM0/rHz8aOgH75RKy/n2p+xmsl/ZdM4lLxOLHlj+fdU6eljZXaEP0fow7Zr
rqCSPBPmeQkDdqRF2Z75Luzb/3D5yJAQNgoZCSCxucpebziE0EV77XXNjieZ
4YPhpk0cgVJPYJuVKUUIR8XJ8n+uC0ZfjX/sqmopjebCMosIEMkJdeiIuTUG
3/vOqo6pJz1w6SPzwea1STqz8jtzm83TNT/V0wckQP/Olf5lDK18m7tY+4CL
4oia/C3Ttui6Zk3sn5oMoYew9pxj1d9VNuuNAfDwoExnmGrSK3H07I1N6bnk
8+hMVuuO/CZ3XCNs55srFUHiZS+k1na1bTndKUSy8MYupz7nzuKy1Vy76HPj
Mdbo5t8OOlxSjR44b163qkdoqVmC3mFNnKFtA0Lgra6vnfvZvAbgOPajT3m+
McJ9s7Ua9Uyfbq+INpvyshQDS7hq+ysOY4unLk7ry/OLVBllzQHOgpFP5bj8
BuM1K5cMJ4abP1f0nmBSoTlTRujgT1VgrgQx84Tu2OjyUNkoPbTon0r3Ee71
fm4SMRuqxBJWJdDAaAvlDKLdy6quMBUB0gnLmwzrOg4TGqnZhIbrHnxTH40V
cjOGJgDBqYhCLdqdFiEKVcxCxrNEAZgzPP2GrfRIRTtuTOLVnPxCQBsWvb0S
MF/pqXEnwPDe96pIMNrfRnB6GTRkGUxlWrfRhSINcxGRBew3mJj1yhnQaBgR
yaab9INI3irQO6uQzItnGn3xDljId7v+/QdaSuyFiH5QRtdUy1lSymltiHxj
Pky5qbfOED0quh6edlnhrN3aaWEWsRKHjj/nDh/cZ8T+c/CIatVCY3F7NVjC
bDsX4i/m6k0HkhvIkO49D5E0jBIJVQ20PAUvJ1COplQRFysRe2+jPtS14odR
9Dj2hRLttL8lw6LfkYgL4BJd796OYk/By/9h8D8VXLPsF9h+KnfBeV6Z+PKN
P1cja65fBxxc+2TsttqSlMvvNojKE8pCLYuJFQQVS7tvdUcSwUEkScuCVsF3
IDI4YjWeZMfQpOPQ9FXvXnEQz1HxzGtXbhn80+SHf3AjA0ECQDNb/F6TQ/0N
nAb5/xDflJ6OQD3O5qO3vzHU+oxGv+zUdbNywH0WYA7BHTK8UxW7TnStoBvi
+AakRGW3DoV8XyOW/rPR1Q/WY8cKom5oUxSj8vbcA2S2mX+jd3Ov+DWdt8Kf
1fx+oHTbjBrWY6/18GypbBl7TCYLnGDltqP3BxqjfcKE5uAavTWP3j0Yi3ff
E2wvUMwj+f4U1X5GDVrTZK2kFbic9kisHJGtafSRcwQnI7dJrjey8Yrt3bov
yceNlwy4SpPLKqNR3BHCv6Y6nQirSM6nOonP/XqkDInjw46qpBKWrOB3tQmq
BrxPYh+hY5/NUQeaYaGOuusDDR3ZZRo7AEryUL2G5PhBhW1jhONf4tERxzme
FUT2gznPVNN4F3sGFenfqn/gdLX3yROoF6NLsQyOw/AaXODaV3CW1b9TQ232
OmMVLoIwDyQEvwkF/WbznfgkyQjq/MIVb6kakLYzaqtbM11YfW79Vi0e9xrG
njIEehK8NQd3nPOQuUrbsijcGzPWphB2mq5DnI3PaEadwk0eyFaVNo/Hghzd
U88v5YgbPmUK5UxVwP09NnuZOQwJWO8RoUqCQhzOjYxklgF1LW3n7zlWOCEE
8MTuTIQ1NoCM9RrT7+0OnltF0Ar3V5rNyeODKdHxE0meSL/zp9vERxrSwAJG
kvA5or7S6ADE+RxjFCfNg58CEHI5Nv6r5bd3RypvgnvHZF4saWAS/bbrMktQ
zJFke/uChko6jyLaAfqAlVF2o/OkoTAd2GQwsI/EjXHbMP1giNIceSSTs/JD
7G1LYgDskEnSZavefLAuvW+OCqujMbS9F9p8WhcAMLxNowKQSIVPwFGBroBi
r2SDU8dcZFkuA35mE80fw9TV65nDUz/BLR+pgNniXJd0AHv+KAtZ2ZmGbd4c
G40QatCEpcC0N44TVX1HSba9m3ZVMiuGngKsgmIicXK8PkC9tMwD/xSO9Vec
RgVTd3zAr2Gju0Mtlo5C3EcoNMZ0FWnsgG2yYlxwB2wyyfgJOi/mncu0esiD
a32W7evy19fnbK4bDEogey7ivyy7n5XA4qH1dBIp4g0J/2Ujk5xTi/iEsuJO
d3Wkhx7Oq7e7po78T8ndGn31fknFc+xz0xm2Oq8KuTE1EW/mOWv28QnH9Ip1
YhkCeDgsErseKcAufga9/DGKVqrZyRdnaz5ybcfDxmPfrmRUh7taTRtnsxxG
ZeVwI6Q4TUX8QQUSN8pwx6+kHz8KJ8nmrRfe91Ccv0qNpiuAcUb5Luk+Dfyi
N4et7WwWN5bcXZibnSGxCy+gaNCtGDtfSUYX5DrKKpYRwU0XFCE1LOwtISRz
ZM8QbFWzLfB2AFlYzzi/fmC3pX2qbYHrCcA9fFSiVBu4T7OELxnTA/GuVHQE
S9wzEctDXTdWkYpZxR7astIrE7RvHVHFYTWxarHfDpIfCefcB5+/D5Vulnzr
eK8CClM/B1ajM5e7SteVqQj5pC3AEGDfmXI7Hh4CCT9wH/hW617/nVD9Tl4+
XNoTT00sfDmbgHhdxRy7ovXzwZBwsSHWZsJumEdEiVE43vqnYFppZY4RFe9l
3d+SJTMz37J491ms8yn/edd961nsqymjAFomQHiSYuZUUNH+aZuuJWDtpXbH
EBMVO9qOARYHoWtGFCY1PP/PwUuFYneFwWXtChCqKEqJB+NUXCK/otkm84xB
3rUHC0ckHqaDKwz7sFW4qcnzVuMxc0snT+2fGE6qk4rSPNUlzroC/d7Wbaey
oez4kAJmCpSU8i4A7xpiVqRXR0kxAbolS4JH0NN9ym/MTp+O+HCcd9FXCmV8
EGt168yiO4YeKH7XdxMof5JGd/1GS70/GGMZsGRFR4Dso7rHUtFbmd2XehH6
m8+kKXQ36QqlKVcxwpLHtR8oJLYOLgVqkitCwIQnX77Itxj9Nlb0GO/jqu4d
ux7HpOwZUqs+mco93VE/hnErYb3x7afl8WFgXrNg9XfMV0nTtkbimdPzTe6V
E2jLkGSMCVLUxN3E/vbZzDk4MBh3uoaIpoz0pfQ7huk+ffJSA99IoeK48npY
7OQ6Xm0f5Waw0KMQbnlLwNXJIP3XkVEySiuFCqt2gULQwKtMtXEmAC1lsbyx
Igar8MXhcjSKlIwg37F1lqqgomXhWpK+MejUIXqQ6E0wSuJWN93txAR0Xg1A
0fuP0+wEkA/UjUjXAqUBIJWsSTrn2/4RL7N1X+3KiIeKne+tg/y8R0jMUygg
rzEmFtcEjpKgM7UYqOpIaK5m/Yrli36ujDXMmGQOZpBMSS5Bt/BERz74FFQ1
quimxmVKlDyzaAn1cEq8LVuvC37l3p+lJRRNIWErAigBHywi3XUVrsi6u7E8
6MrGvEvmcNOZdNW6P8OPE6cAIRtTXzPM7I89FpzKktTC/fWrKMhSRZLokDQt
DEA8QEe/zQZmP2PXKF+rpQHqHwnQCjhVWGJMdeVKkqmA0bmO6WuqSme8qGGU
f1ybd7L5SfGrnYsISVSx32wcLs8ASVG00PUhlN2qnD6H7P2cE/urXKR3zXUb
kxq7fYL5Zw9pL30vEME1H4h3rlQCpUC4KmFqvmPTjP3xxAQDx5eSYWdYjyrk
CA3ccMyMD1hEo4d3yepodsWihlhhdC3JPxlPhalP4n4Vl1WLxOZC9tBCiH4R
gqwl5Zzp+r8bRGNqfF6KDrTy+gEz7VhzDY1w1ZaNh0hAbawAG7e3dbgXjVP8
8aDoXh3Yk9xrZwc8Tqoif2VqQXNtcc3FY3sc1UolQROIY1YGc8XhtdZSxp+8
IZ4oex3m3UnQ5/kxbyL1QjBAByhEeXT6OnW2uOPcFVWQj4L7CDRJSdN/eTMC
M9uANg+tUvZXdZuRqxJNNvycD3IyyTbnFYoKCAHagCtWGZyYyf5EzNm2Efkv
PxZkDmX9pYVx14fx2ugFmqUjngmg3CqIeleb5cv8mrZJ7J6PVE2FRygCq2vN
UFxGsc+BFXGFMRG6UYWG7qOzu28brFhK8SjbZDmYQJJshkFs8pz2zzpgpMlk
Ycvod8MoJJo4ylrRWa56L/F+PEj6UJAItXTuQxG+HTEuDny8nrmeoxJT+5W+
5bcxZM1fOLvjx+movkaLSsfao+bRUDyWP3wYXbhYkZLPHGceln635THJ0PlJ
sNTGg8W4FDmvpP7Fe2w3t5o825RXfojopi5jImkN6wvaWNhxmIN5njZcjnA+
tZ4vQJc0JvZ95POEVPFRu3Z+rbw8hhc324bA72e91gtyXgIxHL8s1jickA+f
eCeybgMO8FjweOs8FGo3cT863Q4Ha4crl+OF3sGiN+dOll4zXuVIw8z7Jm+M
CEf6eoUFfy6vcyVz0kjxLvYiAyvTf7VGN+V3coDjh0iBWYXJy8jPfa6Ap7tY
bZAqWEakrhDD6F2nMbcNdGQpyQAefO84BrSEIcohiD8wHIx8U4mc6H1HWw03
m7iiyahUtu0EfUTQBi/Tt5SfeaX7eU+TUDzuzSYsN4SNRVid9XmFovu/4/fi
t6O0R6H+mMxzH/WZuBSWhfv2hUAJvUGV0n7h+NSNvG3hCA5qR0H8oVbmR2+X
rILt6Qhi75EZjl9XQwRl1QQzRk/6kNzfTbhrQ6QU72Jhbyh4zEDOaeEx6Sfj
C7MS1/FZgsrOPLV1LLXAVgLEB5iXTBv3yfV1GcBDfJYqlmTbFnueREusfD1z
vBvJ7Bsr6hDJqXPtakuabJO5zGCsKWqQ8LTpAjs9E5RL4H6dkxBOVv3j0wKJ
tEp63Etg7+FKhNpaOQkJlyurpigQYc7zQRtlpsfN3uuEm19Pc1HZ/JKOvl7w
NMBBwsHaVlpPKYZG4K+G+STxyNaj1FKgZrQ8OZAmLqYONcjp/JlKje1b/gU8
TbxyEs1d++Yk2wdkKitbwyJhku6MpzXvLqaIZ4EYM/Xh8rUodm4AR/aB9peA
ICEwCaEHqagBBWW9V2N3mQdjQ9ii1ItS64lpOviFQSJJLZaNxfw3RtVeWA7z
FlMHlp6K9gE9IMjRCXs66KAYAlmHNgvOThB2okQGVUBIVw1mqyF9KkJQhO9E
F2GXOGlNZXpxk2KIjv7loXAxtN8TjJq62nZCna2AutK47p7wMBBIsAX0rPTE
wPkvEocbo/yWD/xNgzRHVbFkK8W7gzY5SAEcGPqMJ8LEpo4pudX1tmh5N0rE
iARIG7ADpnPvMYx1P6pQSqifPhw6+XdkqVagTfxIqYI3wv6PKWxnaL0VE9gc
002z2otH8zyXWRt6SBDDTp8JDw+VD1Vao01DPvwlB3tfowyMdp1KmDFt+eOX
Y2ifLSZIKcAoFCKBgSAK51b4p/h+NpLgCZ1TkcDevYD4jGIY+bs0FplZi2Jp
9COPbE+mDWofaCLBv9gn9Im91j3u1Ivxme+9qkviFOkuEM6TPK/6+bGrgf/l
YzoiU9xQhMEYf6yicj4SoSS56sA4OjhYOa2yswOwGnC8Wm+d5J0E4zJ0CyYB
2Zrg02avDKAbZTUMAwTAkRHyujhqVjKuoFGWRA9UtBOFAaopUF/x0i40ZHT2
7Wel1gRQJlCV/Q2YPfMZiLpLtLMdBFyebUNFdshpzqaFMhZpY3Md5jI7XdLm
1dWVSE1LwXYCwU6Hz8hzbSVcBuvg92X6Ek6iLobLp4pWy/dzFqBoCLE6Mioz
xCFnGx2RDKOjaXG7wM3zj9t4ZU1S8uOxHYsPfV/4g+7S6Xg2kwJeRD4/uzbK
QGLEbDJxouehfBphYUiLxPJOB9Ck5CLNurOLOZgfoLPfNuyPU1GB//Su8wIN
NOX8f5PwmW7W2k84aK5vmFoeNycE3ZA+Wp5fjpY64vCQQj3G47KMNqpvszNH
aiBhOgjUnoqFGunIQy9WrfXLO1pHZYxuhlmH/SBiARXrm9I8E3lGVJuBEvTZ
Y49liR+JvNwWXEwWQIj6WdQu3QdxUZ9CBQL8/0KiEJp43+nQwfXomoHKys++
++mZCnWatOBSy9iRASyJEpfpQMy9U6kLQtBPIwHoUPdost4gC+vxES6WbGms
uCt+SA3xrGwSozjRhVbpObz6RLhl68nbxR8APY65mzJ7y232iFzddCuuU3ld
75qEUSitrJL4BCNoT6aXsHtCf3PCeLl3wk8N3VooUhcrKICX+yXgDMFZslho
tdT0a8BnPfxjuYvnttUylPTdgLW+4zUnT2AwIG1oJHrj14ys9zIIXmNUkwwh
VEafoz92la4yXvc1WmBRY/aT/k7KNMZLfed/JjxHr1tc79oKNAmM8dsoYMkX
lu1LM9me5zQ0yOSPbGtDk1iyg1dxk0jlJPoAxmMKzxK3/bfkeXly5tIXcsYe
9qOUcFt6HM9Y6ugvG0tvAZFs26HBXRXuytHXlFFrcHWY2MuZrvyBrEK5kmbh
wTyxntPmPe/E5ma2OtR6xZPBAr62fT+vU8hYcIUIBzik1fPsumJzU7S0pyhx
JQ0QUzTpFxYedlm/8j9s1MQ6rCZnfxV1fxLcxZFsW9cfCkL/fvmKwE98vfaM
xiSl6o7kvzzNezrw/dO2P8lRIj9EAc6bwSp2QoQ05eml2afpOvAti7ry1I3r
av1vs12J6PKCytptegkJN1jEPbYzzPLUePVDP2+59Ps5lae5MKrA09m7EMVg
d4y6DWyeN3TvnGjiU9jA/5YvAQmIl+aaNSaZP6qpcqcJCrEVqDnigA4QIL5C
PDA8rWUeE1nX7TMgUMZ8aD9m5PPmpUf42xkmjZan7cY1CnKq47zBk5MmfgK2
449pEeYPoacftXH1+HGVHSSo2bQ+8w1/dN7byERaigjCmicrFFNkE9WBgW1m
Ws1wv+ORaO0ky7evP9cNHhVu36FHBPhpnScKRuRRK91Qh8f+wn/TYUEoloRd
0w3OfTxbpqSd2oxA4QasR1fF4KzWm15aB6YqUKzoZxRvPoBBCSyoF2MDTwZQ
LjsSUgOZhihsbkYGMlh4eCyKRXz6JsCJ/Yab+zjOlO4av+kPhb/+k3+wHprL
vMGvkshW28VJ3amGXJ4GPNZpMf2tMmKZghyalIkbgY4+waGM0TD9wpQzrPv+
mJEe6uGPkzVdgcxRzFmwxV+McwGVXgZpVIbwur9xxEQ1H1l2wJnVaqROTcoh
FZlNckCMXqFmX2bwmx+tYVXRFIca51GFKgzC0fNr3H6Skc3NpReTPA7EaAtc
gCOU5YmFejHgmAgH26+xcDgBboNwoTgGmaOQ/PG99bu/PqOJyIuvFTrHuYvy
3+XFU+r8leVopCLxWK3ucCeK/EIkyGDshgQAr4uxsiiLu4Uz+CGm/T9SD8WL
mPlTQzhA9VFBx18ZkRykxP1pA4thm4w8ZeCJ5fKrYqHtKjPmgplf6VOVvnV2
R/evBD2anLiQuRuQcfAjU+/VjtYHuUsxaUrBKrpZNFIkkuZSoQ9tQGZl94IU
qNT4BlO/+hZYSCmK/fRiRNIemjwsmTluIRIyFtPtnOIXmbGM2HhsgLjaXSTb
GkMzqzPPVoDSx5BpTxkZRGCT6k2p/AxJJrM3fgL0k60qV3TTjfwFkrlTAI62
yJeid2W65iSXD6p3K0M749jIbLRd6R2yTb0eGNRwqZ1gAFrDKvAUF1GGPy/P
++PssFZ+Rrtw4DVSe3l91M6vhpoYUeAWw5V8RZIuO8bROdZoPfjiOHOo7tC2
NTM6mmO7PdoLaap3pVv6GBf6BE4L5DzauNmdXK0Yc5LLIRfVvEx4d5AHz/wX
Wvo77MR64YpQnajtNmZId2bWojtCbZeCPQsztcNkrrqJ5721A0ZYBOYPxMcc
Uzs5pf4LQWW4tun0KArOdpdCgyc0midZCpbuwEYN2kbjynK3zYBgE9HQLzOT
P6NhUeslM26g28lj7998aJ3IfMZFwmkVLUdboI49MdFRVs7XnTcYFpp6UgaS
bAZhLTSGG88hSty/Qjp3u1/LW79XbEpmaVzyl19GeTlyUr5/1I0Es0InP4WB
UqsEcIKyGip+UikCzJmvTi2JbSrmC1XRkKEHwdm/wQHfNNvblUXAXRJ/yWew
4zoH44srI2c4jBIf6lBuV0VprhcvdDgeWVkFPCBxIg2j1Xuu4y9AR/S3EZRY
aHNN8E3AM+xkwTruJPDKZ6Uj9QDoM25OctriYc/SnMlnGReYYaaVWlKRJI1I
N4nMZfLkPiNrBJfNAlfCqhwZwkUMJ4bT6T6ZZSV/hLIIRzrFn/61uoCKiew3
BZYsybhsLi39jiHO7lR4WhUppXndLnUjApnXJl2QEUQedKCtd1HjexylAx54
5+dqOoilEgIcBoy7wRxBUBCb++EcUhhBEtagGdUFTrN0jZ69xiP4spcJzEqw
B93rWpWGhSZfsG7/5j2Xcb7PO39YWJLEnBgi4ZnWna/bpK4Dq+eTuBGxJjZ3
OWanDd+Vx7Vw/IPXmc0J902g90UPCqekaHgTZJhmbgiFZv0gp3ntR36Y0rTF
MRMWGNUQBPPadHyhwQazAe4VfaOA8rvT6YaWog35omrjb81hCAhZcDhX1tO7
cfldLd+6YvF1/qrbsV9Hbqlggjjs4iPJyUoF6twrug1fr1SbR8abmvSRknrC
JEdHI2eeMDPWYBULxVMQnyL2D74gx1KioW9FPaXEtZ1HUHh8Gf6l6lpdRfDa
IUOb2TzYtaCgo7uMevcqGR1/KmpJXw4WLmiM6lRLu9K3ZuBcyetUV3CQ1v+O
CzePGZjIdLjPxbuRPb4RpyQ3o1ucrQFDKX45QxNrPxrp2TrdhaYcsX4jvRse
+owFaCw2eSr6b4XscP14qJ1w5br21XBxUnMb7MEgJGdzksAdQ/pmmdbokFpE
sytFS2hk0MAUtq00tmedddEadE+G5lY5WpJ0rpzcBWHHiOU8qAIU1k6RXxqU
joZyVVxv5ZmUHFgfTG4pZIoX7v/5qiiOM8M67Ie/bcaVjA7I1XXjWzyPNlMB
vKGjuyrv63ApwrvbbYxCMCJn1hF5bSj+ySXYNy9G4m8ibQLHKbGuKDJWeFBK
gNKgY3+EMvlfB7lHlp4YYS++hNdUVUKYcj7vYs7PpJ/Dz1svaJmzd/ZD88Fq
VelvDcIg/0ANoYsC4WGGb4PW16nkqRWoRCcpqN+QcAdOzUe+CjKIalGI/1yQ
3/rNdbSXxDfBtsgzoETzIkuaFMSivqlwuzs+HnvngwKmEmgU5gpzZc0nYlSF
eAWJDhEM+AQDxZRUOhgEPZIBWb+U/vlNiPYftSWfXhpByC2d77IgbqrU7AXs
JseH8TuO2QCJNQk0zqeRNQhgYL6lR2Nq9gyEAchFANoQDPqA7WbVH+46JHhB
2Pxatujz5nQvUZRplYjiwPskuuQhV3t0HAYt5k9FYxLGRaEKYTWhcYP7aj+w
vsFgfXe4poo7B740sDpcEn/EhkPLUSf1iFBxPmDOIIoStA1bALhWg665yFVE
hmYdZ9TKPAatXyT1BeEMpaC4vNKi8VGgcuSJpy8jL1Owwikqjp3GJJXdaQKd
QATe9eZOUnDsWSJpo8RRHxhFFw5sHEMQUmTGrPkiBBB15lQeiZI1bDjSjEin
5VtQCEOKb+WDvmGHmJSA6EpKc3Kf8eaY2/eTn7jJTF1Oo8LhG4noRMabHTNh
nuAcjoYp5ZvZipI5QVjnH5Y9Mh5bJGJi7l1MAnZA1DXAdVgSv4m7pUZJ0Btn
ZhLGub5Acm2hdRcGy+rpQzqxxtc4uNvo2yGGucHTEKtwI+/EOlDXDvRzpQnC
d+F6+q3gKWswZVrJHhnkLtdsZ8Dz2UTqPUKWuFYoEHpdveGtTs8Ap0pVcz2d
r/WPRzr1zzTb3HHcrzV+N2/bLm5NbkiLlDs0A59iiclnftOsFWvIxA/dE0tv
SUdtg8mPmvoolzsUykqBffG1GHPd1DTtg7zKiEQM0ACdKfyryEUNrRTrfdod
EwHBLqWYSHWMsiZdgSdYeHSQC/4De/wUtJRJfvuNbsywW1xNcY2YhNzA1gcw
GwB17whLPgwmTayIsMCXnmpKi9+U6qIO7ipysAm2GuHv1tE5fqjVOJPe0Xpk
Y/Apoh5xlU8Du13s582obC0sgh0knz3mDomzKNw7lr2oeGOeP2A3jLrvQJj4
FKLupN2mWgJnpIe4IlLhsK2KqsBwn7f5nDwB0SGRA2R9Z20T/I6rOdXWUN/H
kSFNXKm39Wsc2KctAtddgxLwFD42Q4jusCYe9/EKML7JWwG4E3g1YOWa1t3j
SDrwHdDi0dhtSynyNafMa20yH22ppRQk9H3C6z7W9I1Tmggp5qH/vgOKuM1S
gzbzsoqA+HTFel2rGlNniDbtnbL0A4Ut4A+ZBxUTlJGUHgO43Zn0FMkgDJ7s
6epzYArFUI2595znKgV9BApkZthdG7rvxIIHGj6QnZaievr1uX6HIxPk8ouL
k9wWvWY8FmWi73PmnkXUUsvf0HLstxTXWwQXlkZq8B0zBntCy6prvkHjVPsi
7gv5Y2u159UeQOo/Snfyclmt7cKV8uwmJ+CopB1BNDKS6CQs7KN7hWDnUE5h
KUnOCOci1BNXF2+4u4w3pQfTYf4axkcTBWsrTHz3mje4ZpkiHMriZPWvZff9
zD0I3AlY1zQZblmG8Sb0IpWlNQVwQI+aGm6Zyy/uCcA1H1d8yvX+ruukk9HU
VJ16wOJTla/di9MCYqp7CkwFK7pCNzcQBeubQbAV+lbIESbraetvWZ7FlMzM
zAGN4RwK5HrWlgbWDfHuXm1XCP/zyRIfSTeAT1bhIoq99CfMHK93x/5C+JHR
IP81k5Df2/VFN59+GIREr160asbTCpIwrKyzdQCDiKJtruKMTdJdFhV3fnBi
1CX4xfDPzyP3erHYtNAyLoEjXsVk6ZvAREF33Q3Rzj5VJgoWeRcyw3PKlpjL
WopM1+spb/9qpb8OesIwYWKHrQhUp1VY7SfvZq5X2WnicwunJrhxUQTQ4Sof
NakyN59f9kXq690HCG0oZ9wAKbiyz+u0tF5ckYIlKzkJ2ikcEBWiQyDoolu5
Z/zVNg7x+p3B0DifxHplth1w0caKbxoG2ixCyka0QLN2aOAZHiho5YQqv+ty
BpL+wsCwQKtzHeuMTw5+IW4IsjpmkyJK5eBlWD0qo9Fh6iDN9VpDIPy+Mg0+
w+ijJA2UhX8uFJFsbaPNfyz/rRIFnHWk8x+4WcCOP9p2PlyMcEPxw0wWjgf8
CJp+r859MYaECmnMqHnqopopl5+5pWLn/xEWQt4VF8WGw0HD9nJPIyDDNYX+
DBVsNPVPE4Bz/93fBhq3+FX+hQqHL+8gg+24Q/Pu3zRBI2enWPOXy00LXxt4
CcGLZAq1cIFcG3z6rddUgc501lhuVoUTJ8x2uBdcTt28V6zuYRuHXPFGD8hV
mo0GMYnj1rEN4wGQqE52xt5ts4uPFuYvvCM+1LdGGyIbh1L75r1lbfVy7+BJ
dK80n2a6+chIov5zhNGgeJ9sUfSnaQ2clqTnZh4s3PU/Poh8acCbVg7eay4C
Z5QOzoqiChlGYuVzYjNuvp+F+8VBbVAwMBhY6b7bws9WQwB2H/cvIjN5oE23
YpeQyAOBQ1nNLH3gOl+GqtivwD51UDZPLxxpsMQprWUXDt0hsZw8TdV0I1Oe
t48IAFgg4GGmeTEZo0fDiFENkD/AhEtE7m+y5MntZoRwyMrIBPn6Hi1hkPf4
7scyCAVAsTsf6kj++7J05gWeSFaZcAoXIYN9l1pETcRtCOMbbUIQNq2Z5VXW
Y/8Xybf+Pj7FS1KcRvEEj8Gi1JjBkwbEP/jXIQP2yF4QN5RAlfJR9jDrvU5K
lTM1SMGHZhYG1Sm3N6PxXWfqTYnkyJooZeRR4dgM11pDXG/nXkhzrKk5+ono
3xMrwjEghsf50+pALaUd6IoCTXRv7bUFOVi/oD06WnMU8SVSFxtmdrFk10vm
o2a9kFSHyOm6GG+MDl7pdNnF2c+PuWjlJ1CGZyJUdBPAMfvs7nDVwqAQNx1C
2Ziao7xssTpuCDMcRn2wy5yc38rxMOf2GaMTocgBMLfQwqU+xGk2FyoW30/M
KQpoi1F7NkhS54suseUbloFtOD9Km28e8mpCR2sl6V2OH9QQJGOYjsa2p4qX
QxcKgmlwN7e9rwXlSpu0bUSuJIRvMOHa9lsgETKnFzV5sCoWSnz8ZQyAHp5d
x0gERFis9gjH9PAUxf7koFFBaCtIF9+Ufy9IiEQ62IjNErSWjsrBOXJ4Ktjx
uNHezYrdqRTWWAwUd4SR+p/fsqbcX7PLxc9Qc03Yc1xx6rPnd6IMJbT31Nwn
1flZYOy4HQAGtdNwuOZmszFEYXR3x+L2EvhasjkPqyOtBnmqiZcQMjeaShLY
39XRIOnNxHrsSzskGQei73jdq7F9QSfkFYpk64HSUCjBb3DPruD4UTDWu+cq
wc6LopP5o6JAkkutFYFZjSprS6416CFUUbWU7gO5iOcswvsO3tqsjq2abpW2
3uTYg9taRCtfKQSNpGrcW2AHp8kfGs6CpyZ7Yqw71+memUZ0nE/ceV/biVYr
RiayIv+5wHjB++eaIZp7ftJOkDzz5wbz0uOQ/J7/5dFhQa97pimR75zy5sFR
I73CXldFIwuJX7cKeGlLZJUJcNXDfNFB7kS+mM6ewe6v+MX5N3ONPLfwtGFu
kCJzFmgtLdRPZe4ua+Ay2HJO9zw3QosQpBkDG5+9kfX3HdoZtNc1Y9BEczW0
7RSBGZVPXFkcKYnZk3Qy6K0ojiCR3Jee+xh1fvqqkkCCprCHIIpDQvvtkIZK
YyLF2B7ckEqy8D/prkRg1SDxXVu2caN+JixB9BaJsX4NoSBmUj1ikrJJraW9
MIJ6/KY8oVMu0z/xTsPsIsxoteFc/TjcjzjxPmGu8DvyjITmOdY8PiFrK8TJ
Xz/B4B/fY3JAzYo66b100OBv+j8UqWhClbcvepETo/G5/sq4JF/CoLaod7Iw
aYQjQM3zKAmTF6Z6Uvwqi13U06g+q3ftnXCM8h+LpjLgMg33026jfQzK1YCp
AMx2pUNNXupw4BVWF40zbbh8lg8Majli0wUZGq2Ab0qC2ezEK9TlC08s7Hmi
K9zyWQ2eHfYk3tlICiAV48U4YODvrcw3x4uNfQFRCbQJYTEtC20JZm5fj/FZ
Siw8Omr3CpE370H/JZwOnk63Xui+QEe7mawcWhWmVW3skpJzL6HgaIrO3qcF
GUKK66+/p7UV0WTrXLo72gd1Hs5LwguFR/wyU6DqKWKBauS6SwkHx39SPRgs
z2g1A7vDZhuSaSk8+Qqw5Koqdmd+C+0bOwseMmGiMb4KQtGghirrJ9QjGytd
v6qi4ZJnlXLXaxjdQ+WBFoEgPjZo/F2iqW4zzRR7MhWHCpzX0X6bcc18MyP+
uskSErWN+dGVW9uwqt7u5QxNIzo6HIeTvKL8Gfa18gxMbFaBaiUTl8cQotF4
RALyXupkX9NOKDokXeq8VZu75QqrCpcUlQQrOTCxfG6nu850pTycaxxUd/s+
K5Rb5wO4CNgKW0IPZMGRF/dO3FRtVJMS/975J+cU5xB3QwNlNPP0FYFxgDYe
fLc6f8jWrAH5luTVtiB3SH5mzKUbuXJeXCDD5MDg9oIfMA0jorM9GNnI2QkR
xLQi+yFItviS3MfZNjcdmffOlElm+3BqkpnzQM6QEx2H8JH/DKlxDoEibEDm
bum3Pqn2eRiy6aOodW30DVEhvApJ4tyw8pvVblS/18VMi8BGR7aVAfweiHva
8pSOg6fyJpoHVZNuXnJ00JQk1vv00M8vNLfe3ZmY/O0AVCmsCa93ZuYPZHts
5geBLjwGcp5VwFqdBrG3oIT9ILDXtnq3HxbEBtLe5gtr3aFyKqNouahozg5F
62xApUYdJROgtbX3xf1aIU+JscavOd/l+mJpMXst7BSH4WrV/nVmwxrtFIAL
u2GgLrdDMIxYsYoE7s7HKX8GenVIo4mRe+DUreoWqw790meAeW3UFA10DVo6
eXDI4AG1tccd91zy2pZh4aj6LBx7MZ/R9rUBQKUBVawESa5Ko6DJURqISHvd
z1le6dUs71wRaCBh7mLHeFZfDM5mrKEirHB/uo/sblHl8JLFhl2mCdpxbcye
Hk5b+5tAn9riZCZ39Kl4QBfYv7pAibn9aFTJNtL7ZzljicpLg86H8jK6iH14
LIaKUtE8Q7DtYUKgbYeyK9d51T4RRq1dYeYtkVZjzp7cX5NgJJnwnZLCLNz7
Q1YiMFxMp9e3KLIiEAbWHqxR/S0RShUqSKPpmqknnOwZKvu5HMEgqh3QvJYe
Dy4wyuxh0nK5f2aspoSCeQtdPPvXSm2JL1c8Da5eNhqvvvK0WclZsPaMTy5E
I1p8kMdZoYeqHJ7rtE4OYs8FV1stztBxblQ+bUKKa7qCz0OImB65f+sh/wpa
D9VOp3h6++c9Olol1rhi97hZBL4r9Pt82STpRX4j9nACSQKkOYQaHvmOCaxH
zaE7MtzEv+uH3NVQUX7wGSr7sD58TMy+oAxlQDi07S6OPbdvPyXXby3bySfB
Z7qNUNLY0UaW2m2+dCkTBDUokitAzPWu+YC5hFYvaBUCv98GcBBnqIqGXW4w
0ZmQWMngECCiQ3G7KefhH7tYLpXDa653R7SX2P4IFxBOxml2Y03vJE68oJTj
l92o42vZnScDOR2otm3kQEyy7vvEyJb42CGpLurYp07a15F/4/sj2HteHnMf
0e7c73nT6atD+RObjn35l6q/Sz2xfNofA+bYwvQ51/P5pqZFT76FxKyDj7XJ
DdMVCTEabJ+VL6S2stpS7+zZ7txUa2PSnhlXsjwGxaqaO+SYTxBkrY2L9Dlx
QjMYYvPfV/2m8tJJuLDzQWkIOARS95cbTAGK0llPdO7R5McRrxnDf5avVb99
afh+aAbEJk9JjsI2yiHagiV+mm7WQWL0fMSzv6CWCxpLbDn0Y7yV048EXXAd
TKU3IShhhgCEg0/M05br1U0Eo6HMd++UYTLuDWl5FmjetSaBk15PsjFIZsl5
aCPThkEhziZwLy+mc1kf68cYygF76TFx7AnInhqUdCemWgekr1tMZXsIMiID
z+hef5dfuBedNPksX0vklKu60fc5/jY/jIkl8nUVF6Z/b3C0ZWyqD5o9mUmT
NlLh+MhLwCu/Um77HDFiPcD/mEI1JnHueE9oYgJevpnT/FdYlAMBdRRRblYx
3qlpKkfuCaBjRA006yiejUQJCQOgDEqY3pZU0lRj7zn+3k4sb1J0QWREV452
SGYdMNrqLo0zTv2dLl9Ca0jgWLT7fj7mepFNPMw91GRe6zAlG0mGTAWflH5o
TNtjDKzRtzwR8NqX8VPd++uudY0AwYiYzKyBaJgYGOXL/ka8KXpAk8yB0evx
+pxox/BvcEukr00jjKuknmeOqCUAqK33O2sX9xwsJRzy1zTMAv3TZ6E20MEQ
0kpQr4+l+fkeIJ7/KxZkVzkxMntVsepl6q+41J42QiTEsoz6DZ0vdJtje69E
zGTYY1qluHq/GBueXhfsNa+U9MFCO9KBrQAix+CJ+z/LYfr1ptwQmsnWUFC7
kS2MS/cLkD/1lcTJ2AtOClv/WIKC2Tu0RQJSzHQX450Xsxp2KXq9sSTclFML
VnvmaLN2vItLtXcmg11MMCufKnbBsaS7hjINnsCqyllINir9vQffzz1O+aRK
9C98fyxRBdUOpZPnbdu3loS8edsG0zyN8FjDHdWAKHHTplBNYob0FF5dS0kH
fSEu1fpQ/hBLWgAbdiaQ1Ds1F0hu8dor9Jz1zPrNxbPoYlJfdVAW6vtevZOL
Fnup18vCxbzQgRKsLMGm18UMhfJZYOpnZlN+nDY1ABOt839cYvaA/3INAh1N
oGoUQtEQ9JyLbGrg6YwoqluDaQ/XhF5Q4+J5k+W049p2ucqPvXEeFMVdaGUg
vEogrxz25LNm1S6X7+YAzdUGOYo1mDiv8EE8DuWlQD+1SRc8bvk1AQb9nBVc
aDat5hk6EICeXYpZSMzbcbA6aVeWdakCngfkk5WoxWWaMKUm0bdIYg5RgoHo
0J/q+Jrv2e/SP+e0aqKj2Y6PFxSxstlElGItrUpVl/c7VkAp4KgEUQORGA0X
jbiRhAxPyIxEpWaB0miy/LEEQmklRJWbs8he1wEjQlk6wmTa8fuT0m2G3cjb
GQ2YCUWPIzRNmehpEqnUqYF3appin1/a0KZ5UIzatZJfzYWho60HT1WXj+lo
Z/Dhxvu5wK+IQPc02bsxkYuQ/7VBSiPphv3C47oSt1UCx2K2LY9wOLLKQJOW
nDFEUnPBcjgcjKvffY7zAu8rgDvRM3q+yky/i/b5b1WSoideivK2VPAypOY8
pisaXXGsKru7fymQeiTI2aDOzNXIwYfbsAbBKis9P0GFHBGn1CQUdjA847tn
Ik6tlEpuG/Qn+q2dPc869i8PE99myv1Yukx0At8PVloi1/SHWb9yZ8b2eCau
DRNhVIGsrx9hAtE9jBP/Tvb/2MaHgy4CuGx3Q5B4PmP285L4e9vQCbUErote
Cbn5oHYNxMS0aiSg4KAVvzQeDF5S38TzHv0OJwDGP0otYerITxG/p+RoAxxy
wKxRLTP3ZESCDjhT3UV/Cqs9quv0v3U88XD3uhjXN181J71ilR8pcXtYU+TZ
FBf6mYWe7SwaPWxbTvxRFGJRXB9FUol7O9R2n243EGsEhfqk1wMs6liM1KiL
ylqqejFzLB2IT5aOaI0Q66U85HU14IY0XC4s76g1PN58xOM5oIb38Trv/HLM
rDdb08f94Hj1ot7RD0ZyM1brOi16I0sjOa8i3ws3r2mgS/LW0eRxi9Zt4tkk
365VOhO/O+It7yatXatdK+wWee5Jwp0e3MV0D2BtDwyjHeUwrDt5TmcrMri8
0AxBSMqftSYWi4WMxdf+kY0TOjtvS4NpHSb4Z0vuB1lySRPHEQhaUjvaOYCy
XaFa+K3qvGv9s31vB0nZJO2UyO4x+T+QHuMfaG2fzJ6S+igpLTSaWinxn0eu
XqqpgnLGJoHXqPivCBNE25vh8FKm4MoYfVQ1WFkXL4x0Kj7A10c+NJJODqB8
T8ZR21IBt4Zd6BOeLfqJweIqM59UVWnLsWPiOCm1NoOqczVz2QZsCwSft3bh
muGRzzNmLu+Nv79ScfDsKFR7vYIjASzXwfYTKdLrKPi8y9eNm3Mx+mkG29d1
NEbcrj3PY/uNSVgxXFrQazSwr/aPFZtQT53/PjBG46RpGsmT+k5/hvRXVR7g
QS2P+bLxscj69jESUFizcGSr9CoQpcGUdQbfZ8OPhV/0KiPY7ppMrRGLyjqi
g9m4Ch/S1GxSFrz3PBr1F2XjG94MmmidWe0n8RAt5WPIVw1zfRXX9ev+2UqN
mbzxWaXJJ0AA8Ucf+h5Y5OjA2/tESt+6IxRSI/614sCnxYURqapQPpJ/aZCX
8be/S0zKVjv556cU4c9LQlvJtzTuewXFWv+S1XnddfkCeOTPDZom8jplTyt0
CsUJSdqYz5cFs1rrSUQh3WiLpN3Fsq8Zd+aWYVsxQ7k7HJs5OmCqOg4bTW/0
0bm+yAeYifXYZ6VtG51rjVb0JgAjVrlti0wf03gIXS9HUh2gJL93Xh7xBYZU
l+bMnIzXXY2GvBooSEaMRK7HMAP1Rf1kS0BoVEa6b/j2HeOsyGr1P6+QsqET
PmrOrhoF5KpzcE0Id/VgwSHERbDcX7u+crel2+gDFGpbn7xzYu4G4LIaUcxX
s5DCaOAQcLAEsFfwToGqjTwBDe+xjiWr+qVqqkI6nz6oF1j4gOQewVrTX9Eg
wBUn4FcoePL5qUcJ14E7VmhsCjXssVw3b1b6e7/XTdX1rlwbLBEh3ohb3y0a
YO3sRGnWB8zxjTd0LyWIlZAIftWZpRLerMXWWjJjGOtqwu12ikUVzmBk27sZ
erNvkKTF5Qq8UllUk6OqlpHQb89UYJKeuXeSGnzxCQmjc1bNehRQmXkI9aZw
0VT56N3gA9lAEQrd1wip3tU7h62La4uKdz9fgkzGN4rRG/uSUxQL91kd2cLK
KBcdOrZBSK2hX7FwofkDWltcF3NiYaKkIonMkyGOI8qTD4W7SkZWIoSqIfyl
F52mn73QZGZ3fMvIktqULMcHYaeK6MYNaMV+md7o8ZxQEUAFosmPtiHN6t8f
yvMtg6nnjpW7mhLrMTTmp8NRujjk7jhVr9MjYNrcLqVIck2Zii6RheSOEDy9
jzMyHUMo+MTSXue1ez75yuPF4zYSaWbRBx2oTJLkjK8L+GvqzSD4CIN+q47P
AF70/ZmtDSWnyRrOVGYvZAs/cVHvNXYOOqtvJRBbrQFrg+5SOClfx9/hLI6z
1lUgRqLAHXEoBPxOVVHEPXsu/do0ZtpDnj8CEHoflE5hta7jAiY8gMLmFI1t
xeEL21nUUW5RXVuDg4y3wWzEhTbkam20rzT50dOm5ediZIEUNLa4oM+q3CsI
TFRCA/9M86V5HkF9/XJXpcMtFfTJ2nbfe1pXh4iQgbAabHp5IDR7+l9QjYur
NwW1U7KeDIlwSRiw217lSdVMLoyFi+3kNFnrEZxeuYjmWCycffqC4euLamsA
H22vXZeyUX8oRwb2Knos1nkP8fL3G+peXWlgVbj1/oA4L9w0cGqKnhYgzEbI
IzZv+q8VDNx7e0DMlkvb/uJZVMWoftLvH95SqG4Mjtnr2g5FcNMYQSB7oPBl
zdPdwI5INEvGzuPirZLy8rHrsb73DlEYxoaw7oNOvr5njhd6mwfO5r0ix6cw
V70dBZi5NGsabdOSrjJKomDJJQNCnS3zxfdWXfZYZvqsykcbiOVZGe6CZWqH
88bnd4abDqEZV/fDnK3Iek7kjF5Wli0KUaZJN4qE7jVY3BLtgK/H6vGRndPd
V1N0DosraEpVV4uYSwFlPIzQs9VErmAcSZBgO4ElOTXvnduCbeGHZjVJNYPA
SzuoXifJUUhXHtKqbGJNzw77fOh11oWF4LrLef3t2rp0K7hSSxbJwoB2dPMb
HvuInFkX9rMDa9XwVGhRkd4Tf55CuHS8ojUeEtLaE3qhsAmnK8rH3itdnz3Q
E2/GtJiKdNoKvUtJ36NSTI1cHtHlUiQmCmLWch0FM9OcTOlcaJqVMxuB4tx3
4jOT16zawlQWEfpyU+d50s0F+IwAjBtcB/qfzr2mg87aFXA3XM/MwsrTcOgI
o1mzeVhU3fvSm+84A7WReARtiXciFnwuPm0PbFZn5SP3/PRm3TEvCtdFNIig
v1PKO2PmPKHk5AkLsZhkpFiAKGXHpdfahnd+/VqiaJyM1EiyAlavpzJxswcb
KRt9iUwL5hGP+3LJt1bq+z874Io7HBgHNDSvOzSj9uuJnaU1GUiufvi+DpJ4
pRh/d0uUzM2j9scIQnQsmh1DQHzyD9r6p11vd+I5PMC3mUYIT1CwsXV42N5t
uJ/FfmAtOLJzEa+vVMXzu3durc3AzpvezEo4WWmfXprpQDDoQzXbWks/ZZuY
6q7qcHKnn+zDzrsg7OK7FtPb6UzYC3TwI21ReA7s2wr0/5KrNzq8DL2MooL5
/gcCb07A9AMSXtbZKyfEkqXkZ4PxNTleg3ZS0gxiCqvynDwRqCV+FbHTawm2
7S1x/vxgTKPQTdaQ0EInkqKb0Ud2YXFR0GsvjvbtAlgMtYXBqoosblMpl6ai
ro3qhd/i2HO/xGigfK9MH8QEd+FxQ6lD5iiKdUji4ow8xhDTs5weq87FIBU4
iC117uONQlZEnJGzMZRmnhEm+M4BsfeUAtUVkfQi/BsV3H55Y/p4L4JQfRtK
/f8KZZjNCkjeRmBWL+V8nkfdhVE/t3Z3KnvpCZF6Mp1CJI0tQZrndTilWsIX
efiiKEPGA99cmVTa+e0WqW4nI/obZO234DvOxhe0umsGebq4MKVRqXjF2Lio
f6tjJxYjLcYOOyM+uiV8Fxu/fBdBa219pQZFY5/lyYuYB7ZYxyqCb7f1r0vU
iPhNUm8v4Jh+5gl7/1yavC21ZVG5dOLAW4TOQSo6eC0K9T9tm8hygkV1gH8q
0yODe8cTBNUbRnXhwGhoFj59AL8iQHIFOAlOAbdm2SqhLD1tn37HJg7m2XOw
aEOrhp5fSOtwTZ0cy0K+/QiF6d5SmwRcx1LrWNBAOr1uhY6vTHVhIvSBWKrc
1lA6NyDkeI+X+Y8OSbPBCdTa++K3/7NdlDSX95rhkZlYAenrghgFBVm3VTaS
EP0fRpwWkMcZXHrjZG6XbRlbZEPuT/lOJ4uYo6R0oAPmZ0e41U8kRIksbCcn
gF3pYEBKbmkEjG19KeNCe+CrSj06Zd0FpFHjFPXrz2UTwk5eheueKcwf+U5Q
tKhut2UTJQK0yLYwjGvRKckEPvivPjMktHTQXdImAIORxpqmWEuUeB4ggmYQ
8MMgVU5wPN2f9U7sCqDpHiGkxKYqwM+IjQY18hCTOZ6ddNDs2rSnKUAzNr79
q5PH5xiJ2CDH2guEj6y1Qk+TgIxNeoN6ZfG7eC1+jBElY2tQ/S5jC2SJ9K32
wIiIxjNPqrt8577iQ2Je7ot6xQhCMfUmAwqik3IXvR6ZmRyGaP4ZMyiwPRJ5
GxzkxjNOyWU9Z6EeBo1QcJVk7637biGZBE+R/DHAGrRbbpGBzlnI7hoy0shl
CHl+gMyvGylfY7PsiZzjC5y48TUOMvMTXtAwUfxNUd9QH27aCLZ/lbP7eofC
jRSvOJ9bghFpvOnaRelJMf7mRnWwzeG3RGSBe5F5yXNW6+tyBwLWMtJVcT7S
nRbk3UWvHSIYC7UqaZXHQVrjQKidasZAyY3OFXkXf07TInWHOEpI2joz9GH4
ccrxj1lwJkb1U8DhsMX4zHgwk5vB8ZGxAXOOnB7KD9nTqtHkUjbvHjQ1boE8
Rjc7yof0+FRLPXADiEIoYUccvU99Ru8kymaTQYriY/pn/fX8z4dz8wkfE1dt
C3g/eTiVLdBGnA/cJ1RPwlbTzsztXRFi/tJlE+ogohkMX+gvW67n8y5vHeM5
5+5uQTspBhb/b9kIAhkWdvMlWt4+c1YA7xyHsMiV/B/hVBkn77Pl9b27FTbc
Y9cU/lZIGMSYhEEYV+nyvqKibxZzSlUsnoTTDjmX9fyUBAwlWhibvIrmlAPY
HZdjasRSU4fvSrHaPFdZXeu9BgoURhHU0alIRt4VS13m6uMAa3g2J8rqvW9D
yeDfct0OXsN6zfyRsjSQRj5XhA1qMyx24k0Eu8UZPaGcvfdD7mx2gAYlfmzl
9HQJ9M7KuEEMqR6CDdVCuPxY4TmFYEK7Wc7kyByvxNKPAqFks4U+paMUoKxV
I5O939NwAGIjyrmXh6XRyxrMwG1PaX42XgKUJaa4mQv1nIdyVT7hNNNBMXh0
edMHauA55b3WIVfLLwXv9kuPonSXoEKfQNCvrDOtbE8jAvEv69EB6hyEyXqd
osyk31/M0HoxY3Nxa8LCBUWoBI1gxu6KJ0FNcnBKP88ASEYZDqy02wQxyWzP
LjSODCsYJAYL5BT869It2h61zDx4G10IqhGDZAKCXMStwsrSt1e70GxJj06w
3vmaEMKCUm3AmHMtbYdkgg1fql1Lh9nMzKPugLDzjda5yn1JpXmvk5/YI+C7
RVRieDvXGS81/qYYoZaD3PpHCcA6nPR3xrsjqtEQwLQrf44qxABOb960ppOE
XznVulAMcXZOpkqDuPvp5CFYAJF2EPYKOPL8p40YIWyD/+MoLVNuHg6pWkjp
ULRTLk+r9wq9x12iN13zCCfGLwqN0jQIAYUxJOWae21TLOCW8uWaSS+u+uTu
lixlf0burUEJ45pcret88qnhsuNslas0S8POnTyXUzB/Ioe81RNM9l5Mlewp
DK6XKP8nyEIWiUjK7ARjpHATgWvGcJNluf7TcBfgFP7kn3o6PyN4Uy3C8o68
Ft0um3Xv132jUSJbj8uzZg9nSIgfYMjqGSVoKcaZL5EJScrox+IvYULHIP40
WMGjOBYOinwbaJoGRtH2au56EB3WcR9GVTg9Gzr6iMQbVBjei0Js30w2icfs
rOsWrqQjTMVqwj7ovLtb2l3vdZhfhwDsIUnHvF3eAGuv7DEb6DQ9YGPEaoHm
kRbzXuz9X1CDt9pxhhXVBm2xCUpZdY9cHObs/PpPd/sd2zQCEjz6NXZsuO5r
LCsCXfQp7c7eI5AJq00kR8UMzKITEwXNYSSlQYNTD4+NeFzr1WQebqjgpBMv
zrlSoUbbd4wzgaRcyZxsilwGWvA9uXCuKwNuRKY1i/Opsh6jzMv7iPXL34ds
w5O2a+yI7FHLzzGV7BFfX613kmuZCxJLrxEakojUDad0PvPmr8pVdn1MAW8m
R3VJ7eM/QiZmCVAUay8UM+Wps93vYWz0FFanx/Zd7vi8BWYQhcLysPGuKh/h
FhXvXfu/v2EMXYruWlPNQ6Qr9e2edIRLGhsHIxI/s7GDcopEQzIoPnHBZq8A
Pl0q0mFshVfgHtzEpBrfAe2UENWaV1ETd2CJAHoObpbTBqIhywAVsD/TZCCm
jE//4I41fEKCmbvyn2kccPqTS/7Qs2n1+lU7/+cA7S0c1mxQW6IUn3JsYfqA
ylYovBcf//zCc/TWSiALEYayXyl5tg2b5ICjGCfkcGkUD5kXIDyzr37fTJ5N
ncOXf6T9EDkFSW3s7g64FWL+bU3FwZqjcJkiVY9wz8PVf+WcILbisOr8f5lp
OPSOn+ugfRjv394hi3axqI0tc6ogHPBN8PwQh/xzGzsEcf3lLbIfnvcCyoBk
TFpbQ8de+hx5yx5J6RogzJjzL+f8OOXF2CDEuwXiy9gZebYWERqipEdKiCwU
iWJs+MBFSHX9Zy3fTqNXAnjzeYWScZ1wILSvPnyDOkoTJGFiwXtN+slcUwgf
6EYnai40CXeI1W+5bVXPmG6AbfRHqplVK/UvrNUDmNnteWBSXFt6eVFjJO7d
1121KU6uquoGSzJv1xQEe+pnZmM1dgNadiFMFvqX6TfJvryzUSme6dsG0I5I
cUvmoImf2CxcY34Q5G/PGCqdz2eFsqPHRmjh20VjC6N+qB5GTDYFNciAZFrO
IzZ/Nno5kfgFEzgvfR3NfK+ess24Xo03sHXt7emONijrle4EkFPbdU4QNsoj
Xn8bbFjwD3QnrrPJQX6HEzeStcA+2pKSTxdXYG/c2IJFexXCbDx8/WLEW0zA
NBb56ips82JChCH4B8a9U9p+V5qQ3DOLgDHCLTOlji3TaeNnmpphvHJ8yLD/
d1QYb2RdLJ9AayPENbSoXZztYG0mIHIYUFOpf6lVTisJF+YO/AbRJ2nJK56j
0SknL0MErMiS0680T0eJTa8UjeOIpUHGjjn/dwiVAt+Kum/g+7YyXfrF4pt8
J1uGBSPAoe/AOfi4Msans/nJ+ja2O22xt5MjH2vFy7YxrnKZefQy1wm4Hbnw
7PomzhaSwy1SpXD1FsKZB7nSvUAfdmxTQ+50FyBHsW+nY1XU27S7H4jqJBhI
Hgcm3rE212B7hopGjCFNTXjm3cZn8wnx8WlRd0GfhqW3wLYv0p9tTLnX4R1c
UsfEP3lq6RUIA8IQiYAHnBn2xsf7z8m9mYQfsrAZ3jIRNbuDYJImVAapeQht
KUQvLm/Q+b/56cbu9sjCndynUtMzqq/4BShF3OR1sdnhYgBQPOdnowdQaix9
KoTQHFsTcaIJuI5perK3J4wERvuNO6RCH+kK7ko/jKDGZmxXrXPdCq/raI1+
kZsRGR3QEf7VBRjAFscyGTad63DYljO4/eaqHodMV38mS2e6BN1dGtXV78j/
JxN9dsUxEJgdDUEv/XMA47sGC+QzpeWVybHFaqSAX9OWM9gTt1aAAD0Ousl4
lLTbCgXztY1t7erXOblTFy2i6T7R0H7gNF5IUl3BBt1/RH5IXV6pnWmyFMi8
tF8pJ0894k1a8jR5twtmyTn1/MCItX4fG48Sxski3fyfVzUndF4ZP4p7DhHo
uflGDXq/PTYbqEqgDBOqKEpShb8eZm7guXUo7FkBMYAbwruW0v9mD/699fy3
hZJNobziQnoBL8VInyskK4Xt3P0cIn8Y1zGuMKA9JyLusEdDS2+6EvjWHxPN
+yFgGVncPoafZhDajr/KVgmxPy8eigGG2TD8s2xZskQpMuapL31Tkp1THk7L
cZZ8MPRCmmSKcI4LkVfuQtQl9Vmd2vQab9KWPdnBNUY+DmLbpvJ8SXs33t29
Vcqz2+04A31YFqo8dao0vSITuZDyhA5v8oOARKtml+M8tbqWdkF/DJSq5cBH
ks0sKO70tpiHO/fhTT2LPNMOkNGZ2QgC5c4W5PvUeFDyAb/QmIil4KH4b/+c
ZCiscysoXCtP5yLRr+izOuIuJ2rr1T9XPTfTJp6SOfMTNCxhzWBPWHIVVECz
OJIyP/+InK+0LtRz/fsMhclDLOuAXSaoL78+RKI4BESZkI+ZkVAky9GzEGNC
cIRFPZOF1LWfRVRybVZmTkbof+tWRshopOXuxAfdwteaflAEEQiGVBTDVzvu
QGsL2kz8inaMIJNAPz6NK998cKrt+v9CVre1ilkjQ3kdANfIwk6dijfQdQZx
yYdnSvo7BA9+/ydGFklasvvnWz4RhX5NUzIuLUMZZqdA1y5I3nA6hQHDDkqN
pgXk9W760Hkqw4B0MfIfzfVyL2W4rO0/q0alFIXuTMMtCcBXUkgYl/+SKLTC
JtGvIctKBI3U6hbTnVC/aRor0vz1iITvNqxLmpjSXKD2RJH+RkOO7B3jx7fc
KqWVPE6sH3H0OI+XwC04cpoX1EalKkw8tdF9lU+HWDyM2MGJ3l/jkKde7yzb
De2jMZgtA5X9fMnXE5IF0nGCKN2RdEWdcjzU8jwYPPi9PRAbrpEKzm987auD
J05hDjnwLzbH1CYbLadzN4ITD017wkkvF5yPHS7pm2/KfYe2cBtzCyIrObML
Z0f5ygHsTIJ4FBM6uUYtbJtKvs7T2RuCwdoZzbOBFCpwDe5pRmsdhczK+gLu
Vf+HBr8ymrHJCrfYB/NBrqNJatiJSudS7XOflUe/JBbL/X07EozPjq6hs/Lw
A/n9S43BY9CkLAZEErNbm2G3Xu+fQtsznGEF8BjnXTbFthi+GA2Y8etF2evU
OPbrL9JIAijyX94xV9if2Qa35/z/ywkBAhzl33J2fKL07PhgKo6hbAkDrvND
1VNcYx9YrZkbQFN4G4YLVDMwHlgsZKiqqfDBGv5qFdZH8RgWFc50+wbUiOeH
6D9oHeDlc0z307iAi25vG0ZyumyFASNMFvaftRvM8Hc4ReSQyaL3Z0O4gPct
Pap6SzJuoTgvfKjBWsqfTSKASPIUDLMUTfmm/Svtd9RgbeZyNdS/meE8IBsR
QA+Q5suRaBfGesUbPtOzgF5tboOi3RQ+cZOp1Qsv1fIf0k7KvfGDIUITDwfr
plsj62x3vNwdVUp4sQbCTuWu1idyPNF2jcsymJ7WXj4CThlC/UoOPhUf8G++
soXzQO706pztnAqhYxnirWvr90TBLfjZY0NF1swBPs12ZDC24VRxRxwsowTI
QNeD1xOM1J1KIZp2cZF1STbxUkP5jA+egCFpVg0GriSijUEZmxSD12Hkdw9C
8VkwXbuH6/sGBiALK38o7ZJ1srr2src7HKJfPpJr5qyPL1roDUiMK5WfD+Ek
MgLEsVmmqOEgQqHUwMACPji6b+yExO16n85Qu1pjmkxvNspnQKdBcEYNQ6Zb
2GYrX6qtGi3MHDMqzS3XQ8Y446+wSIcwAivJHVkSKWNLcXEyWUyi3/hvnM/J
vLJlQ0E/OCP5vovVYnU3xK/D/8qq+pjf8QRy4GWBhNenux2WDaXIZcCtRVOr
yj42Vt41mnuSufJ0maDXOtRTM2cTLgxkejHleEMra+ASUk2NCRcSYlu9MYa3
Zi6AxG3bgV0Y3i7qgMWbFshkfHeG/eXLG+xGQ8TDKdlhidir56Y70Hz+aR3y
dyUqTStOdAgvpRG3HdmlSXMZzVdI+pAFzNtrYzkLfPc7r7CQROmy+cth5Wjd
gZXOEOsjRlNfiEtPBnjMKBN7i79uLGZm0T7nDRb4RSaL+OgGG2LbbP+ySsob
YggBP/x9vYXDiVRoVxJZ5X5k4FVUu9fw5mbmbhKB2wwlsRN1CK3eKQfjvDNv
z5RhGtPqgfPvX1RuE70okB0mtSoZh7LES6rOTwp7EPa6jMhLwpH5SGme5zLQ
LRrhihr7cOU9Wh+xBKHVot4Sg0fUD2eOBerknMLX0j9efXSFr9vVDvmoJk2g
hmxATTJ4jPIk2z0CNdbZp4GT/l3pamzRHGBW5FMwBpSUiAk3gk5B1YfqJIdo
Dm8jFUfvLsFyFvy+1nE7zd2RWNgL+QYnatF07EC6XTLqoM9mwyXlsI0avc+b
K7P5zSK9Ewp3a00hNVyIMPKEuZHdpYnmz8zlqk4bq82fPTNoSlVS7oJNekjX
eeIWRCCNtrtileHloVhHtgmpopzPc+Qm1DsbDfShg8Mcy9l1NCr2Wl20D0Y+
2vwF5Q1i1reNVYdD3en4/s3k6K0E4gUCyvw5SVgjQPuJvOWhKv6xHAYvVGRs
A6rUff+XZYy0w6RX8l9z/Lda1oI5wxDVb+sHwO+PmW8JNqbA4CuSgADcWoin
mQowbEIi2tqsqhn7dATa6vhRf7kxBTp3KYfn7vVYkIkRkVJ/SPwjhKSRdS6c
TwqXTx9p9PN9TugC/UzG9LnKrlPs7oJ3nykzLtsq+GYE0/+N9hFvZDmEyoed
7sDy9Rg3SPVIbjIq8xRbuY/b7/E29jNLzlaJ6TLuc+gZWSiE+l0JFlPeAkxO
J5g9G81lzB7Ll9RTQmvcDvfi2BA1G/QxY7OZAULAx5otsmMdd3zkTNqVb4o5
3Ic4tHq3PgXhwp/8Ti9B1yWHCoe9hZkl9uoLHzfaoX3Ubn2d5g2mstRcFwnf
cHy7qKhUUf7CWY/3nlDHKRj5rRAuY2bHihDsxO0qu4My2l9/FxMGVsiK82hY
RGh8EuSP3OTlPnKjg8C7f1S4vqon+esRLxGXkv2iKHSp+HPnILUV99YtZ5lA
G4rIrIYKa7P7fjZbuaGGgqgEU5EsfGjrbiPpfcX8DcCMTfDTLBglhSMeNyRJ
Aee10XxVFe9O/ZTCv5pDeHvA44RZKyFaonW73RPt8tbg7ROSUgjLQnq7RieC
yOBc4WjpHPhMOB7JMjYl7hI1ZhbPHGGdVjcZK9o++zNm53C7tDDgE9McpGFa
R0lmUawk/wkmY/V6rPsoStBctmqeXbjbtqNn2bQy8nlqKjraSIEt+YGLoVa+
EpbXK5Huj5HI9zFenvz8ot48qg8kKYq314nvLRBcNWrQCW6o/uwoR8waFZhF
J+ACplfxuKrg8wEJwWbKK5nYPgFr8r5+82GykLhpRdsTpxpAtfEbltRKung9
/NlfCV4Qsul1WHZ4mqlYpcjBjGFHvMiye3f5xGibaU3wkVgpKoGo2ys37aLn
XVPi46gsOKVfaBtmJTdAcZaUC9BroWx2hvkyKI/sFa53LcJzrMSrmNHWztdX
7NNRjIeVOUMZjKir95CzTji/ykkJKZozZQCaZpQVhol8bWrSIBZEc7OJq4vS
IJcy+uVSccLPlpcU0QxRtKjsx6tKK6IhgignN+Ai8yKIdEsk3DLMkaxCEHel
6Reu1mMyzBXqXPMkWycUsLxsSr+hqZ80Cj98XtU+LuoZZ1SIrCsKacVKkCAr
yG3r97VqTv+bzc0HibJyJlfkFTVd98KUDyta8T6u5yZX9dxcDS7zPilgb5yR
/bruGspZMb/RJkyOrBa1q9ukIkwZtMAgwdT8hmtDC/KZpJBZ2fRelcToyk5S
zeY4ZWu8u3xEB/Z1HlvV5rUiDDy+8cJK5B9pLDtgep8Fze+x7ZuTHjjjphcT
o5YtZtB55jm/Q8aoJ9+Bz0zbRGrN+TgOK9ctanQlc3FindpyTQUKUKE/fQic
ULVARga1gxTklS/paGyO64y1a/g5R3khmYU/ba1KXnB7UC7Kr3ingMMshdUU
m0tKA5W0+5eIoeeqxM1x5h+abxbuzwgrNEF71JCeKGIIboZbznZ3brKu/0us
HpCkbS0qMVba8hxi2fhD3sXzNo5ILxCS/+iBebiUMUmZ6nILv33r8CvSEXnK
q6HUxXUrBqyyhGrnISu2eVpNQg8oXXFYfLnNTYQKg0MK/yVeIDe8eemIeqUJ
b9zxSj3EstgqgZS7Zl5nvriQjC4TUhGrfbT6hdUv0OBXI9ueFJZjCT///ID3
MOFp2xtUvltYCWiHh6xcdGawbb8+p04D/fL/9tv9u3s149m6s2XsaKvAeJCM
vZDFYQGSEW+dJScsde8BinO6NSzNRVl4I68Cs8oCV76xUrS4WKd9/8TcVFFZ
0nbWFSkZI/TR6FIz8mJurITwI/boKxu7FOq7vN+E+CofCIKxgoK+GRkfNBEj
0bHo9Ef5mDcMlhZIb+HL04JJIT7cdzQYI2gt6ANnL2lXmwjrOSgF8rzYOw04
KPYZK0h04uFwU1F2fBKoZi1n+I/O4aGhR2QX4W7lfuUhiZ90md9T2OorIute
h1RmhbaBzK8VexS3qhvFPnTUJH7VlJ3wpTvfkT3Iz3SjBw6Stpbq46T3bPXT
8mlYQzNZ0RO6uIFPEoqmZojyFz8AJEbYHsgt2HCw5wOqxXmiz9pffwrhlP9f
PJ+3cHqfrKn6obxbwv+SNbtXqcPTLgR6UKVeRdXnjDiiR+WDFrOams68JuYC
Ree/PCKAZ/Nif6skc5H0tQV2dsaNtEYDDI50vnv+dJSwfxMI5TjCdfgOD2Dw
Ba68WerT9vdlf/Ohlz2UqV+9lVPICcRseS7oj2tnQDCBcEgs7f8Gtl8gvWM0
E0xjR+mQiQnphpH8O1iF4jxKCDYivk+BMywfc0dg+3YJZBPZiFQ3+Q5JdLET
NRNhttehi5Zy5fP6blaHpNyzkfr3MfsIcS18KewsLgaiIA34MNvbZz0Hf+X4
K7tAc2jSlSBdpUFO0KYy+0Lzlz9MUcXzz0YgBCugBHtTeMb7VNVMfLO8kTQi
g3aSvM6f+OpPdIPhwYUNndqJ+gkcZdSNI65VkY7bdckQtjTcXMlOXRID6UYg
IkhJXjal3iuqj4FnoD+6uFHwP/8ek0aFEkA5+otviIQzxDDk/hf5I/FVo7Ph
2CIKv4rCBlzH1xwqWLwxmo0tvx9I1mtyRBf5XIDhRsD4M9tkZQNiONLRDg3G
HoKlw9/St901ImdKm7R7WHsd9D6/F9GL6NpXTwXSsD7pEuWRl42aFVHrDt4s
Stye2YByfW693QBywbCSxWjU9jcHyK39JItDcyBqtivBGI6yGKPDAPSM1x12
VKjyGzXhnIxuLJvRImBsQ2M4dodduVInZcMSJYwl3txDXDh7ZK5Cq+lhvOCJ
jgStAy2Ec2VdF3JoUyimvaACB1tioBAvbwEBathCZJSX9UKfxVtwrgRj/tlO
xsOHfuCZQceZ//oVLgMfqVhRkqZolph2uCCT6exXpWCtuBcN9qK5Re9W5wc0
IMEEZ4QIJBm96n7ku+MGEPZ5wzhD+tXfIwDiRDLre2njUQUUf/BXm6VKBjYg
QD83ThyX53ZqivbCpS32CGVzdKnKJWuLqgGhGT5iidxrvwrSbZs/cEHitdsp
7pG6aOnEeVt6rIPTB0hJ0gmdgrKeGUieFwdgCxvXUqeq8DlmAHcmTnCrWkkr
u9BW3RForhzCHA2Dkr1h+btdrn6jfinVV5keduncxg86tBylB6fEasUDcIXN
Bphx4aePOhlsedvyaA72rP2CaxGFTXKJUtM6HH4+bvV692MyKJk6fQQgnWSS
m8gQKllOaimq4WVu2iWmUFzbbWYTSUQS9R7y9/q6FmLa7lJQ9LoBFQPzBU93
H5Ww/Oa1HOp5d/CXl9qxSMHnLrzsFsJ9EnRy4ZuDcM/LAZv1Ov7J6wBgI8q6
M+PKHyQ8sdF6Y9X+YTDXuuQZv2wAeS3zBFm05Y25Xn5LvpYi/O68HPizVbdH
TAvkLhlPXdgEYk6MS8I+fdxE4Mv6cKRc8LWXjkK3BaPqs7rUVoPmvBWFR/zs
dZ3LIjKMSyZSV7GrRf/INCG53HAaIRTgYPo4T3Johx3zSVVVD923+FDiqn1t
O15HrWZYvP57eWm5iwsH6+bCXUXbP2gfSUa0c9CYlUOIM2u7O37kCRtca9jp
0Hgo+QiS/I3X+2N0TAYiK0xepQNlTo3nnCKHoHsRzRMxHWH6WQ3EBN6EJ2vD
9qJAc5Nz3IaJTkOUw7f1f8YIbXPhynqPiH1Z1O62sVWs9fUwaMRoezMoYARi
Y7o6W5ina0JS+EL9/RIGvrhL/XXnse0GzcXQVtb86iwFvxQc8MwDcldn1yx+
yeVS83acJ1tS8fkLJQI5AVkFd/IPIYc3YPXqMf4pe6A+weua9OzGE2kz40uS
CCI+1nhRT6s8PJ+W6Lf/MtQoEQKQcSr5pHcum89mibEXdo4EOLr3tGjtvvlg
qVcMYciyKoS9zerdD612slRtYRbNLIojAAKMWndIjjkBct/8salwILfY+BrM
IsEO1vdwaCgjjrfRFKSqEO8zhwfHi71Oke4G/YJrFz/qIuwi1t7E7hrtsER2
O5bHUxaPeLd62k4hkODF77rvSfyx1pmHv+dA4gq37nGT96RoAiuKAb3UDcQJ
fiSme2O8XQveMrXqPayxEUHw9bGjVS1tzmF+CdXuSlU6Qv+KK2M85S2Pv4vB
3r3WEe117qNoWybVi2LmNPLnXXYwkYEsM9OVwsMl/lOqLNGaxxHNqlBIiFUT
BkhKwuJvSIgQqrOWnneWMRT2MmxnCMOy+9Y9WVFUIUj4eqRNpON5Sr4G9EJ4
qH2wFLILZ3HxOfsHJV6EUw7HL7m/vv8pADPbVgx1QX+VpN4MlUYuLmaZrm0A
+CA6ooshyqZfF3lPlmH1nFhBJfJ+O7Lc2Bg8v4A09wGCsU1qgUgQ1NFQHCz+
/YahIKS4rqy6ac/EwnGB4VnzeBNB07mpaYsigTAPPIE3Ytxf6ZqAFaywcg60
MVnX7Pxple7r0KCUAm+oIH045n0KL+Lv6xp5XZ703HrG0eW+16PxpgH3bXDn
m9NhOQP8+slM5WTzXaDbG6x/jOEUP5xBuRJ2muYuMo7HJd8S1mwhMfaPFAmR
ycIlji9Q493FRnWaPoAAlEFKlmkYo9uEOz1pIluUPBmauz0DJgYUzosHzLHP
dQV3wNA2cwaUAU7CJPIgVA6aTbCFUg3fT3OaofPSpDQk1ATyNRccXFKzGMwU
8lH+7CCJ4vBTAN8WU+tvZHHM5dn/n540f3+IlGI824xw1elRkJP0auWd206b
divOsu3eKjeJldicxFfkgDISJCOoLh13Q8TZ6tgsJyvNKqOghvjBohHCmS/T
4IfHt4o8AibpBTK1hQ0uU3qV9LfSbokwr4vu3JVuWBMfQ9LDuXe5RhRWIfpz
J9RMXoc7cpzDhj9OCD//AGN/sAJEEfF/KRz301B+OEgT8rXrfLe2y3pmqUvo
pTIzL/78bZ1vMAriqFxROfbbeTrd4RD3lSwDbbLKiJs3gpSl5LmiLent4JEW
WIJ1kHlSRnWi8QpCqRCUap71RAv40hvhYkQfl393aRfYOEnxo8mmSLUfyVYx
mLJwtMkK1NLdJM5Ot2l9WL6MlIIErh9t91aLpRv0tcWqDG2WKZHK+U25TfPO
kW+erInCZ0r7oBEY2bOy1NJ7kFqUYugcZEd9w5CFuY1jwdR8KDtto0Sm6geW
2/DreL07e1ts48bu2xnQ6eT0FPdLXGKwXaY05C7x/6FZWCYbF8rIKFWPBfb0
SKtxTuEyR+rUx4eRYv6+qYdvI98tVgpbkdENTPtPw8FsPjnea1PL34VHXEKN
mCNZrlzdgp6JGvojRKdliRNS4lM7tENfjv9AjmQICMKouCWw6v5q5fef8KyX
nelJ8OIC4NykFrqI6PZFbucdxgtpP31czFzBXkVtCfMTM2/283vqksul01wu
XZcELUBvzP2qwYWuK047yDItID4MpuysqED4L9dPIG4HrE0hp2svAojCQihM
cGYnp2990UP66ecjk2f6zLom1XNFk/btwOfsxqmgN5uS5KpB7FeJ4PFg7DSn
5/dhhbdJd/jnsxRSZwiIc/mW3DWodEc5/IoSQwagNTBzdRlnq+Yt4vuS8WbH
ySuKm5HPOk43c0Ge8r7T0abk1vK9U6NkPwlxFAcOAl4Me072u8vt8GtTM6fz
E2RjcqW4W1+/NZZM55BfAx1Kgm7f8nfvHMl91HeEA4tw9bMlwfbDCm3Rw/rk
990wW9sywxPosBEuIzalj3Q8jGMkg3JiA3ZjEE5YrsSfkjzIFJ916JuD49xY
DwtLVJylPaMQTIgFHvOij3DolwaJX4SBw/eCk6XNK6QtuC13oXcWP0T1dAXR
jSbtXeG3nxcNZjFfE1KODZGZZMvd6x6scEEyZfzj6yPmZ/LfABTweCaGqFWm
8jfx1kQgFMGmKbajqJgbzRNGZiN+e2ngIq3ay8VzXYyG5az9OH2RV5nixE+O
FzYU7NesUPao/fwCKHBQ9NPuZDEm/qKhFDGpOxEejGIDomGe1BXk867S2ZYm
063K3OS3F1UA7PVZeU5SrvWYmWCV/mL9YHZr2sPaoX+/17U47I4l/Yr9aK4/
nm00zQv9KoAVf1+BUGROf0J13V0yAM/iuC2jzEG3pjtLWqL3x1mjsk57nd+t
cm4zPKXwli9PS2R+iEQp9D+sBL6e2SI2DoU1Y7KCkKUpikjEQOCfk1UkV6lU
uN249hgeS5RTgvhdi4jGrRzHBf7PElzjuc94kVGkbVpB0qyp+NSqyhdcxjYN
+aZr3Wq8SPpswhpfjRKSiUH36VgE7YpO8v0TVOobDimMYZkEEaPc5K/IXTcr
S5UNnOAqUlHlAziqhySq8tHXF0EQY+LJrnIruwT0jGb2AwkklKim5BjUWKlo
5g3ICz6ElRDfYLbU0ajSIuZah1WSarD1qP1HcbFakYe/8zmzyMDNNhY3Jm2s
PVRyjX4FeisgBxW+m658noh+6rlcbUVpqDqUIXTRnEngtRf4Jzc4M306Prex
FqL5gVZj8rVYi22Hr2AqIk7JiBL5jnbZKNxa5W2dKYi2/cBOXJveiOLG/ePh
W8BcDL/Yp/27RXSgz1XCDK6asWHyTa+yymz48FPWXH/UgFBTPcDAbtsF4zRO
XtYtSqWuTYUB3r8a+u/XuIyO+35ZyOkiOci72J7Zz4hBOeLTRVyhX7bDrMxG
nUAlM1gZQCkuMGZCYEzsFNMziGhEVs7HJl9aKdkCzhJYP2BOHDrncIl9foqO
fyMlnWa8nnYZEsanmBIdd2C6X0zXUC9uZMkI0Tzl3jQSEex+yrSTg2fYEwqH
pqDpajKw6AcXHigwcwylWR6Xn0l4FVCo/D7whwP5BZ8Hn1O4elBfv+0dROfJ
8YJPETgZ6Twm6JaTFoTpRvQmZWafotZENVBii5ToVHxBS9C7rSu5zjcL7vJE
J6Me+pCJAyp3rnu71J2edd+EIKdkm/APNbu7f1e5cx/eWn/b0EGzlzjFYNiy
Wtjv7SAL2cmtrN0fmAzPxb972jVHqcMrveRUs94ig846yRKzI5EM0EtvAjeg
TOQAWsr/OBI0luP8ZsE/v1AZq7zGATOVCx1so+++4IRDtx1zN9R4Pq55kjx0
Xo6k+FUfrO9ew/9uzpv3Leif0j0khy1LFsBWTDVFCW+aIsQLcoMlT3XQCywe
UWQB6qIFh+XLVnEVnb7C3DnbU1N8dprbIZm9PrcTO/5ilEhuodaumaf6aO57
ePrFUnNJxLjuz4o54PTb+pOhqWez0iBpAkyDpk1VYJib/fb1prMqaLXw3XPW
CLKz+Kcu08ZM+yrhwFN2PKTXIrBk26+WlnjyTpmlaln0RDKfrJKXBsu6qPPC
nWo3FmssNvku67FfJb0K9EJtA48kpzju+iXHM3FB5a6qTpBqgPM145ZM3EzE
4FM0TiEDecSuOV17SHVlykdhYC8D+KzdfYmveDzaDJB4lkYXtwD9lZbk5qoL
CLvVEvWBvRbqBZbRmjoIIag3mnkomLfe1LNaafqwVJpeulM9QCeZljYHletk
GSk1Lq8CIelp7qJn59BocPF9tRdFjtKCJCg3YNvmHu+lm//emgwN5wKpjjqw
CFRIe8pVt6GsP+JoQ8BH88Y0wvRIDTS98UHgdYq59GAEtFkoJ7zo/tth4et4
0tMYmggZ4M99VuJmDZhrCxFONhXkjvG1ZCm7xBXWefTwSy76+fQLzgIq6ZYH
EVJ2J7CroPb6Su5wn4/5yAwVUEgjtMB6fsOtrz3cAcBlriT954PtZ0YmGByR
4jfIHSTh/iCB9Y+HaDVw3xU4KcjIoeirDF7HbjWnFN0rTo2rfUDaUQXc5/Jo
d7hJs33lbLuWJU+o8LnEMcGEAhkbWiEla1A2iF0m+blxTl81qsTWqdP+LDnI
rDcfg4mK65NmFchPhkiC7IL0LBis9IDWt0gfK8XMGzfHtxo8F8e8qHoJzlKr
lPNV21YK4zTYK4n9f7xG4/7Ph4eNBm303QoTA5r5SLovlwnApLVo2Vrdlj1R
0mbm8VGGYtPfj+fO+IjeCbSwedYnNK78D7GcrUPcluThpSPnrqNVMVnY/YAl
L3wk12NeY5wqVuRyV1Kp349iFdapLayHDBw+7WxmhBZij/VcDq2XzlCpn5XF
Lbi/quLtosMWvnZFQyWwfprQ05uxT2lpQOWU2z6N+Lmr10ng9VtpvN6uwxtQ
CQlhI4SIg9TPsZpfmBLm70GUp/e8cvivmnpFlGBMbNf47zENXUiNiSUq5U27
Q23ty1a+TQcaSBOynvxHlkdIHfiwelprsbSuUOpdtyb4Bn+N8IKgfrG6c8fM
P1/QP6mBOW4P0z/b2yjWodzQNpmA660itAUFJsh7Qin8Qze3reVacgGaecAH
oyDBJHyX6y6LWauk4tbC97ZNbr8vV4RJbNL1IPzU5HCgo6814fCJhPlqPNiX
IFU/4N+bL6NygVxLU46f8u/CSJmP9th2qQ77O4MONJVWPkeqoojZnvdz2igU
hDr4xpxYh6Zp2HuBdbgNX0yz/MFvIG/kO0nSt2S4OsbczuG63AiAFGDHok8y
zJq0yoCkD+Hhg7TNj9LWIcKQdvH37goOeNzlIyBsUi6OJdXNXNx0Kqz9xYV2
U+sDA3J66HKNVXrkXU8PUlC5zbPRKE3vsHD0cc31Rr9OohOeqcOx8CN3/E3h
wJol+dueHvWhHsDolsWyi/0fJPL9JpS03da6wpM9vgyH1rYWIDp3Z0jguqmE
HecPlR1h3EH2mxP2CfUryirKabpzsyT4XdjDOscS8owMcNMGhoW1qR6qQmkr
cCfZtRAGKtcx/pEzF3D6Ukfx+7HSfZAJwvDrbZkINfsFwtnl1lZNwy0zCOQg
rypu4vUCTOXn453aDP8zkd5zzsvzubqLRz1P5Lvv8f+cci9cJcrTnmi89TjO
6oAbXa3ZL4oNXyY8XVLm/OaRfnFXw6siSz9XhrEv/FOF/7bSVMwUZbZPqQ3t
U83g6JfjGFa813o1Q3QxYcepNN7dAvNEGrF75lRygpjhhFHR8HCveGJnz+/6
Yu55OsM2CXCAQZZEr0tGIS8kPR6cHtPPQITGLE6W5ScPZ5umK0TBuvNvV/uh
V97UDbnHar7qvPD90tP+dSqLpGS7U156OF+etf7j1cARCODdxxbZ5bAmHxyI
STwUgsXYJGDS6KD846rh9vf8hXWG3yXAlQ7oen4B6nu73FiRccvgjPc80jiH
qemdEDKivB+rfa794cKPGU/ffJ/t5xj2qsaeVQp+GeE9l/QMy8WbIqf1BXQ9
OhdXlIPhjzbLukkkXAMotl2GBIITMnmIlfX5V8fbsnBAQeeRaUe248ct3ieW
/iv9e7C0jjkwzPOqgWzUDAz0gk/Eq1sr6orOGAdgw2HdzRTPAC1gvTo0Qt+U
1KbXuQxQwF6Ug61zYd/PvTp62QNIAlL7fTi56fHTkTbhvRrFE/WdsPHXDQk3
zVqQ38jE6/Bc50XeUNorDD3PKuKR227s5E4UY2Z5kWowKaKwJjHvTsDdi+sw
h7gvYPWaCsYLWvDT3UH24Y2e/xcA9RZ8detFz+3955ValtUFapFRxHuJ1Sgo
ySVPEGxW5bnEn9rRpsQWUkcUdoj4Ds8Ezl5lc5h/H+c6QuTe3JPF/BhFV3h4
wKLqCj+sqCXFBOn76ib2rDMOlsbXcvywxe4EYJupIRAGdzjLshFGxYNp0pWx
WsrqVJIuksKtLibTv762isQCSGIT73OuPYQ7IEFMjUJdcqy2jbgXoUEAlCOt
DmmuVqm9bitquvwF4exAI9MUNM2A9LwQ2zF7p8T1/Vijj4t+rRKCTT32Xxbf
zZ9UKzGa6ZyEb8baarkrW10y1ctGyrdZ4U6ZGN4xSke1tJlj23zG2TiBAL/I
GYETeN2H56QJKnGZ3fY7auw0BAbhUeSb6jU5ysOkEewYUZTZ0W74VMhHwH0B
8Sh2UyUeY9dxF4aBmFw0L4uLtwYiA2FQCJaOKAH7f46Ed4OD+G6yDndvtEb5
83oolhgfSaTWJPKBPl16Et7e8sxm4oUs5X7uaRJZHGX9oguY++H5N//9hnkZ
epx8xv8rOUb5XSgCt7T2GdvXjNTJ9qAN5uapGXcyLmMfhbs0t09Y4ax+Ng2B
QYuw0jEb9fKtGkuyil54D4S55XVx8p3IKp461wMTpKxdxRe0VO7TaH/bG3Aj
K8aCLMdGwJeq8Desg3wTkLTkp8H5+6/m5HCQ2VLegW5QpUVDght65dVqmkmD
F7kEifPtjXDFESKS9INz7qjUPQQqDXBLVpZluttwFiQsRb2a9o0PoS7FLZ1d
eqRHgNiTBdlNezxCOf9bf+d8XR1KieeEhS/nTwgMLFKq6jo8xNhmDkO2lCKX
Yl+TvkQ5KonlnyOiJco02O9GJNBEiBUoshEXxMhN3XaNw4eiLwyL8zZjP9DC
/eEBg+Ov8a5LXwv44hdWAV228ZUPEowaxGLxJ54fU2VYX4vS0s2PJts1CeGN
N+/5MCS819+rHIQXNCGvBsP1Th+VUYlTnYU0zHccyZfJwrO/c5kgGVuJbykT
1+qaglVWXkSZz9TdS/pLiTv+8UhxlggpPdrhQQtEsR/SzxxXk7skNY+yBMgM
qmiCKTy0vXANXqFJGcdlCnDWT9gwvZYswqTMO/RamgPCaA8AdoOhcMfKigzz
Zqk0lfSb8HFkKiWKVUvbnRKKDzyhKf3iThUstAzlkuhD8ADL6/RA5xrqxBYd
ett4PetoQ/l6OjZf97DMn/l2liu7kjP6ON1a/Vqq4DdXrKwVx85S+mOASe3T
HxCRU1t/18a/TwFfCPn6zQZh5kX0wMspAe69A6kIh4sn9AOcq30YvxjDwMrm
Vd//QBXJvXwfhnY1/QTgcvk+vq4XxfUe9VLze5RDa6e08TeDll5dxLwt37zv
G59gq1eypP3+j4yav4xex1P9p0XNdh21VYAGEpYHmgBTC32WXUEjBGfHjESd
ImjlXpImMm5BvoiJ7Pb/z/lIgHWQAqjUs10AIgOPV3ijTwARBSbfg/GYhTwE
yUDe12hSGrNiggp5GU9lD3TaL15dgVQuTAsWM6lAbw4JZ5U1sunLKcBli1eV
lkB3FKUzZJL7h6ROQ6Td7lCzOkTTe6zGKbhsCBc5CGa6XM//mHjVlfQqQbT+
xOgWIPuFptLR9PTGU/iD/uase1RueQPq3VwPaUR9idWwFC2ftfFw6V0HUkPo
fE6LK8HhnmV0X1aFSJBnxssEC5zUPxWQcgoPX9NVcdW6qANJoc+sN4B+81bx
lCb0ZoFfNImxXl7tsXO6AnyYLqOo2cXk5bKJj90nKofmRK7r4pjnqSr3An+/
qIKRzEWhvXMb3F5mJqFWhC4nDMQ0L1fS30g4KjEmCP38LdTMHBwmjemFxQDi
HasBr8Rle5NKlQ9KJtM8PLHU/4yh+5gAkQNIbCDr1quztaxzjfzv+y/1oE6x
GkmJGIGWpnd6PmShejAr6iIH+tkOPoWCak3QqY/ZyHTfXzHOD32wHxfZMWxD
vTkOwCPNhNq8su7+YLRCLZx4NJ2XSdwA0116tktMbqZqJvNzm7ETmbh/x53p
RTRi2D88zcLHoMZDQtyrMoelCg//O+LmKAnnTVOEIu9xjTgeQHdfu/qhfiit
zuyK08uthYbKrRWXv3MdeZfzHH3BrzwI5ojfyh1gI0rN2fNWOb9e1EzpmzS5
ZP3fPtncCf2LM5/tERbpU4R1vFc/Oe0cvhEM7j1HMJaL/NberlzGZ/qtrkNc
PmSXgKmldUucm0gD7aAJeVEF3hiOlvWEbMnOlg14w0rFnMWwNBGhetUPhR7Z
B7TPs5Alf0YCzaCh+I8YYQIwgm3LfeGeeWgxYwDiX/Y7M08XNslG6z3OR6qt
2N1uSs6guUk5/Qz3MhC6GPCcpYedHpA5dIYLtCXYNjITRi4Iu9WPV/+K3DfI
cfTyC8bcdvvqYH0ekW+o3Whuh+MlA6aiX+ZK8V5Q2rWwVEn648fr54bkoPzx
pT2B9GiqxVWlXeLMrmwz6bWnZiJj4U5BY4H9bRQynwbiB5peQSCpk+6IG0um
aFYgZNCr9AV1cckFPTHKp1aOjh+xPYYamzT4Qmkl/t7PNgDdpzIDlAw2rOpN
CnNaoczr7f2YpXKJgW+LYMkjBFI6exHpVFOX9cyuT5GRyEFwICt3ZveI9wSx
Z6GxhRUamY8o0DUm6Hv6wr0QQrquwLZsax98t5MQOb8W2WUWFmp7wZ58hJ/l
dEu3af3XecEGSJKAoWaW+Vdpv7U2YUz9b0HpNUIyCLQSeBn0AM9ktGgvxTQ+
o+kWyZqpcXwvn2BjA8Lhc73nodRpTgJkG+KohJr+GeXcas1BAz03Jldx/FRk
b6YqYuvg9cEkT/1f9DCIQ751z1h6rn4bP46gkUfPQPvwqItiY2BxO43yyCCR
Y1HA99kABGOqY8MPji4fSaXZOPnDmPkwFvqs5J7LJVXvTIFURPaK44pSbyr9
vigRrL1GaVp/fd1a0BykrNAoaMxsJ5DjU5zl35C2wkwDPPY7abmhFHydmSln
s6aOaNDGBkevKzs/6/WF1t/umZgvE+6pu7il9WeQ9aPkLW33tpLhMNV6UUfC
9RT6m7v/z4gUDycYUp6zvqpwtmO9gqBIjGbCd2S/Dnf+6vFs9X9vsAtz3VVT
9eN60luJwEQ6kDigTpNeYNeLYAqEyo11s0u1y7MFzN0HRQKLseMqfIswcADr
k3tqqbnslhSY9MjPSM7dx1kktv5hSC2xtKXiwYMr8656lpjfKetO6AdY3++y
8sP9ZufGkHqBr8WfAbFE8/5O6RJVSbxp1qlWK1uZnbyVIA2pjfKdeGGCWU5y
vQfkjtEfKOVbw3W9DyQzmD8iy/HeeeEJ5XvzxTjrgZQBkSeqndZmw78vjsya
/W7G2CxMIf9f+X8IpoWGh5M67Rf3AAPe2B1fFFtOG0rMgbAOE+Idf0qYuSuH
32ioNVoDAVNOq4wHoXt+LJUmpyCAmYYZCDQ6bI6xJgvZwDAoiVUw4HuFKh13
RvYGSXeYzyYaKAS+lVg51xX+yHKUmrk/JQe22vhcIvqZJGznE8j8m/evrzWx
GvfAHqWhkuvexz8px6ojUpPWN/ylCEIsDEHRs9+nYdwWbkCt1rMp0DK5sQxb
QZNS9ZTtBkYjteKbSYsM0jWNVOSViL9aOoctC7Yc8tZ9OHgJLXawlExfJBB4
2bqrwLrD5+nibIXParuQ97GLpRzkdFHeBlPvZ+kKTrvsCxmVMTDMduXVs0bK
bifM33PXz7IOuQpKs29hDDMfKoUUEK7Bifl9L4KUBKVQZRapg3qb5NSidVSk
vTJBBqv68zlfeobGwqEDpjuXmJdZZEOCP7ijrfdujDaKy9ZKNf/FLSlzWIlm
uONQHK8sKCo/Nz5kHKrL4gsJKWqAt6BuLwH+cR7tkj+PqFxwR/2Tfm6zUwPa
1ri5PxY/2p5ErjxtbNHjiJrrLNJBJd68WDHUsYVjRTvKqQs9rHtgcUbYjbZC
gAcdswc51LGW62c+fPyoxQcNaLAZoMAA+eKbwJEMsRN69TSA4A5MQPtvoI/9
f/i7znWa0BdMScOWOlckixbDtVTh2M4ZQyk+0IQ16FVUwJ7z0xGWtiXaz2AH
wMA1p+Dez8qFMVasXh7YwF8FwquAQe88Ulh46FGc0Ri/Rwl5yk5cSJkAqbE2
zkuRX3zSqalDZJ/QRZM9yhrjm6ojoK0dZnN1KLQWQ8MmUio5mffyLLEl0dLW
KBr1MqQvpcH8ENzFpDrHYmrNwwZT3sLWR4XsYoING2JFwM1tWEPO038xxx6O
lhd4Io8HBMPaSsMCmixqqYNx/Xo3fpLllPSj2z3zixGVC3qvvOnL6PE25P8r
YFdbY/yaqmrpREh0mquerzLmar+ip9kuks4hZZVrIep5DcsDPc5Y9nG2wfJk
7LLytpqKhCnHYPQF2zgWK+WCeJjAhJTkpZ+bc6J2pM2S7PiYbWSWCMF5dr4B
CXcYK5yFq84Qfy8FxphjBsvOG2T5XZcHTEnVYJWLX2AIz6cN8WYd8H+hA95L
jiSCg6o6g1QYgC6b1OUIhOu3dgFFRVaas+6ZClt9LR4YgBPphNzsCSQeT3qA
RcgwdOVCKmUnvH60Pm0mEzyaxq+zmXW+yhFrUqHgHUGck5rCMBsWLG8iAILo
5aTmifZgVIdbFfsW5+FHnnhlkgrmjOlNBAH2n56oWnh6OncY4ofemHfzmwdp
pGSy/7VDKGgjyLVRl9QjQ/pI2xZgLpsrD3ymGka8c02k18u8r2eIrYJx520D
7tBETVvcoe4quuHXmy8f+b6Eg9ubQQLdLgE6SIqWKaD8OLdmk8z4W2Isqv3y
pcNh99aQKaYR0bsPUquPllkdOFtiPIN76eRAr+W8MdKuVMhNXjtMKzRZ773d
xuBqaJ3YBL2Okugk+iBGZ52YuDRQRPdMMeJ6wObZO1N9CFQmZt57CDsJwKPm
2xBAsQvr76PT4iUhufNCKOzmQSabkM4g/Ol2oKFJwqhBa6XO0zuhFN+mWpnl
akybCZdk+GzG/SNU15I8Lvr7uhOv9WmfMQtKFZ2jKnd3qdYpzAizRMPLvlvL
Boq8UlV0F97n+aDX21kkQMGl96VJl+J+erWQb4DrM9drCevyrQQTGSVc2Etn
D7zUaP3dIIuCJOXavR1LcVxG+ysCqRsnrStneEKYuWXQ/s6NHUzR7WuXUCAI
1k3q9QpETEbgzHvqmK5JEoqyyRO3//3gDmy6AVjYHoMWdGnjwyUu6wZph8In
gwBPJvfhpOQGd2oNafLrWcb6gy8C/Akp5N+8HUNytrLNJJ78+ja+nuRUCISV
88qtiiNFJ8ofLFGUgmN2Lwi0iRfj66CZDh0GT9DVm67wexl70ooXLnHSpUvw
oukapKFBQsQ9RAQQOGAyFCAwBdnOKaxJBHaDn9cotlpWM6Xe+9S4FpratTYw
xxru3NpzIREiSKdIQFPzjCG4EzNDcFGhhjnvXxkoWuyEiZ2R8D/mO40pIfaj
2YzOnm+m+XK74rBBUJV3xRv2DkAJD4mPhG0W6dQhxiKkGFp5dOLRWBD0OZ6v
uU3l8n13VdyU9qgyVQF5+vq6PUlKMCkFYkCNAGxGNFiWGMCDkc3pANiigTIv
AHRSd5h7Zl9VDUQdpANjm9ts+r7kJttG5D0RXDHcqrXKeiZEfOGfEVdcqBVL
4+NOF01mLBSwRwu2KxWVXtwZKl4K7hR8QZtBIdQijyGVVrrzUgW3Qa98m/RK
JYaLtw7eRJULREoJBp1XLgGbFrnw7lNlMLjp15D6E46Tdz925UOteFJ2/ItS
cSklVQK7+SYZJBG2A8O7KO4t4fRK4LdJqexqjq/jvfBMFHFemMGsvyJ+bAPp
pKmH0cKmx26Lp3MVGcE7VdknWaPf+pH/su8VDk7Dgc0Dg+KEaTeu3dNmCaQZ
FY4U/GFyM8qSjMMPE2DVw/twCvSPK/HWCIqhPMJl248kyY35B/Omkit6YBZF
LB48suZzU1kY8NdAI8Wma4Y1Antumm+onvUsXVZ08FHpF7dhh7I4WJvtDmJU
XO03S/z6TskhBu1c/3Us96/m9gw4I0dlfaTZxC/HrCSE52iHMlzjhm9qcw9Q
h25Al5a0CxfF6lIaahP2supzP2EFGoLdbFJcNF9EGpHW0WDjmZhLQ9lM5aGx
UZ3DEluIAOUXCA/w/aQ6pI/dLG7u1HcVTYGzaGBARjF1gO+23lgLjUDXrG3M
QYOiRnHNoldYWUmhroZCXnmWu9NRH/DRiUctDDSHzLA/gb22hYtlHi3cSa3+
nOOlxXm0+tpcYGAxdaV3t89OCP7DNIGN6WM18tsKGdcBZ4xLFIdHJU9WM+6B
3DO0KPW1/Ll7hgXul2oohAprF22/SonR5L5tebPH91kG0NTdmRd+j4QfM+pn
ms5sJt52T8CS6iQsJOplBUQqsD+CNT3IKX6N7oW4SaWYVG9lnSFHQ3M4NUYe
0+7EWA2vokkms3oUEZQMIa+WIhbRYuzjVJTW4Hpul7z1PYCjUEcpDwlIIZ4v
PIzI5/FyCz9eCezHgaYwEiAcpT0S6fjWMeZWFHg9qRiVbuu0GQc/LhcoS5vQ
51qg037ATisRL5dDoKE1A6oHiO9tR/UBz2cVofNC9hdBLhwOKNLA/Z52X6k9
Yn4Ed8EdJnIlHA4JsIiH86OvPfVL9ygDz/zJAT4QhBiHQyuBKUCdx+QK3Lom
siEUk37DkY8DaveBs/v9dM0B0j4V1ceNTIajCTIdfaaYCQW9dOqwu73jIMMK
8TlFjC1bvOs9Q+NbcNH2RDwtUWbPHt3YAzHGsehDbwT3ZsBa3cUsMe9022yC
8l88AKOxk4y7HGpwRWbraobEurEo0yN72JFjhNHJ5Cvu3S2ZIn2i6bhlufYj
XPWZ0sMNY/5smFX+FEdGVsiQXZnS75ejesLoXP0OwLMI7WgqUpMRI0USjU9C
wDhHSxnM6OywG9QikCw1lb3UBRjRvIIYESukxmIx7DsUHjYKQLKkQ+b923z2
0PPHvGD8d4hkbgi8rBsIVTF6dxdrAi2iqSUCV/m6btLulI+pUjS805bOn7mY
SxxZa/bm/4xsynvT3+F1ElmrLYeWyoOilpoEKr8ettePU5bpd18kRWsnOznA
UZXn4Wu98md0/Hnn8OxMU5AGydj83pO9MiHzMT7rMqCod7LslVdNiHMLo4uh
PdKiPSaaP7fjPCElopDlsNvY7yJ0pU8Gx/An7f6y/Gwp9bDwR2pc0O3yjer7
GKvWTA3yI/PeiT8WSHVPUxygDISpqwJ1vHqyI5ysBmzj53+EQFcasIkmpZLE
dVUAOdP/Kch5KLFiKRUHzDB6UvoCFYd0lz7N8dzwwsOOdZAJGe12qjkVY+18
KgsIMVICk1T8Y+r7uAgZBlRqpLUf5dE9QjdR9UWtUMgXRLy0K8FrcQRkVdaW
cTuOvkcXGXCAzvkIkEDdEm8zZstxEyyA0Xsoe3hIykI+3amg2w6RKQorXXvT
ub5IKN3iWx0B1CRa2rnIZFWK1rhI9m0YeZUTD1GBE4n1fvza+jUr5VR1XrZ0
Mf06WTM+uBT2Rsgx1u8UPnQubnQuqlKNnx7tyos1OHB4uHwqnajz7CxBU1mV
AtRbi4JAgKWgKYcvqWzrCzDuI1C9h9OUlrpouEoBSjNMjIKo3PWRYYCmh/2x
Ir2QyjgUz4p5ytYL1jOCgt/mHJN1lQwica6N5LTgV+8JzxdPzzHrcIdmhprf
Yb0QA5hJeLfWTjaaZAl2/4IKbE6ol+ka+1U5IOmMu48kfm/MEyhrYxtnP0Nx
muIQrcICokk/E6a9zOjSXHFiDwEUM2e6J7Tm2BProirk2hXHfK8SFR6gsdFd
r2FLRoGYcpka8WXG8rL2AhtHwHO4/0BiC2J4LEoeTaFzmTBB8w8Nu+FuieRw
KpNdyN3EuEhxCmzTDl12LtJ60B8AHqAA4bqaAUcR0OILjU4t8RFxg92Ha5EM
3XVJ/HKPTZlGaJJY4lZZVF30lEsqfGs9JV0nrJtgii1vClp16S5yKjOZA9AG
zBo9wwsuN6KdCLi/Pfchhj7lcSlGd9+eSNe1fwCYswRB5EzTzYpVCp+cZtIn
dmX9PvXIFTvLLAwVq9IlkumvQI94DfVqfVYz5tdi+V9Lkf2ed5iA8v6obFzV
TuVEmTMF9fVRkvOBanr8IZkF4qeM95nKc6mBadaU+8pM+KlRBMwDUrIpyOt3
mq+doawo7u15IsQ1Un8RSJ3UZxsr0DtcmU/ECFaFe1QNFEL23D8j7fLv3hL+
NONTWmPsOzff1uENVP2iM2tkKy5LNuw5ABja21Hy8GU9Ir8O46/tMiX+dkz/
7+Lw6EqFyH4y6Guv4UOECuUk3uCu8Vy32aLd3aGZHQa70y2z4UU8vuLSWTJQ
uUY/z7GJsS1N1YX0BdVNGKjn9WRim4M9elPVKIsfuA33PAMUvBXoo3k9t7bS
HDbrIFYtIUZzlp2Wtv/6LSWASiDi4PannjvpYL9PGQkh8ZT7XRUOMjB50rQ9
m92Xy7A2XxbLwb49Q0hZ3krphAV+H1sKjYEQ0qMVJ+oQDxNySgDkXwdaK6+T
WUXvZz9y12jHi/3Z9wwc/rY38ppeXhUKQF224OB5AooesCMkFZlTOj3/UlK2
muUmGdWlta6967s9U80t0z4YD+BmGmGKKGF6hxa2gBmv1wVvl52mD9NbuYbp
Kd1yJdkSGBDfPCgqFt/xWE6n4PZmYopIki5B0C68CnSpXYS/H8rTcBXZo49U
j5yfznxmRKMImnOHe+2liKk38K5BIXqQoYeG0o3vmTldHOUOHy15QNiuXReu
AJeZa+nUECHRC4dM6R8ucCa3jEqXeaQLLZZ8RedWjtsX1BiDrRjbLHt8UHgY
b5mkVSjWV4qmelZkEeOmPap+Q+831HyzUr4wcT9FliTltXqv6PusodGcbZ0J
/nPmEsRQhfOpo9kz6ITE9Noz9KNf/daiqxLVEGagoZnpv2w/1CjyERGDl5em
FhlpUF0YPCXO6+YE1/VCg8uRAZ/Ea5G+PYgmM7cJYrjH/XcvJaM1ZWOMQ7QT
8EFwsDqZUQvXK8zYuQhDkW7Kmx2jooZNpqbhT7zAuZv1SsA0fp3uLRd0dMda
8Skcf28yo53+Ms0pwGKPxaHhSxMllGsUQzUFwAz1Jk4g4coQqyVMZd2PusBW
a+uSr9pstfdhkTMOMTDcyzfEobRb/GA+IIRWnJsuYHqecsRJ1oZYQ+XiAfJt
juZb36DUICcKsG+6hlnfPIF34bwct0WggmlVDjkVHE0RbYsxmcDTbZAWxmn0
En2pIaGYPM0CkBF6rBAv7rxeLZiNJyMSRlet0VM2UZyiPkpCYO8QNi/hZ3Ij
hkCXbdpkS7pQidxjUxdH+L79lB53Y+u8a/Gnue4dO5pFbR/NMPronvCtPQgB
uldrYbDWZ+DhZcf2cjpSYm6JewJInooS0W1FhXBJDACKpU6P/WGKg+YD/V3h
WlRhCzLZBEjrlodRUoNubc4IzTwuWQxD20fRv+sjueTds3mgYe8OS2N9nPeO
qUxmhs6BK7ckQdH5VF1fwedSsbRqp4hNaFP1bXsWVDFyaeLzxAyoe157O9k+
Qpp/sInti+7DXO+JCQJyu8J8rTZUdMOyowfbl4RKEsluh/luJBcXKQRGg1ZE
zIQDul5CaRN/5uSt9YS0yotdrYzO5Irwxd74o3EBVPCept/cvRA5rZBXjfWB
oL6+jV+/5C8TWR5jFWOAgQAjmAMqgt8e7DUrEJ7TFyrwQ9kwbYux1L//LfYV
qI5LNkOxDbLor7P5dIiVLHE9j3kmIp4CydeR6utPnHskJcBlYBxNFeSdtuDw
EBe+hwgoSl1Uz3QiPkeuTI7DnqhrxG8SzgfTiWgYvqJVYG07diTBrjMAM6zt
4lwyM5f4grBlwk2EKqzxcGgHFqETTBpsaQ8Lau9nHklv/2dflsu8Nua5keN7
kUWGtSJw3/yk4crt2YMRUIP/eUDTnr18pK3MvHNtV9rSi7HYJHYQixiJWZVa
z5ed7plQ6Er4EyKbfzEj6fX1eq18VatvPsbOAaVvnB1pilUbpkzS1WBiO58b
kemJpPcRIE2GtfURUba+x5GvZmWgz11Fv69lREhKl8FpDTosMn+hkA7DO0ff
cfjY807HHeVnF9fG2FhQry2+a1h4mgXM3kggSBtYvaQkQXZp5v2tY1wTFwge
d2eNOyTEnASyIMRB4kXUEBPFK9XomIE4Xu1LHLLM+G2DG+oYsgqCLruCwlmK
3AnUBUcFs8gLQ6Gwjdjij5+WGnsOTSV8OoYXvbPTi/vYLsWxE5uHCKeM8pSY
7nMkJ4Uv8jzV4LinoCrPR9Ztvx4hQOBsL+v5dJACIeATQFSdPr+ACCF2Tu4A
cLa7jr7dfSP/F50g4eukyb5/+ciaH5yR0UUEhZkYEtmumSkASDl5mX4h8wqx
N7ftwmnhW+SI5P/bqY5jkALM3fOAvTPT1AXweb8rdIzD5kmSFgvhWrdDNCTg
hYGLB1sJOuGbiEKcl4bXZa0sbsssg6ydzOI1yhjEyjx1Vf3k4F1hH6Ka5Adj
o6F23UyJThXcVpw93q03NdoTJ+9dMUrBk5V6fkjSSASxOpl+iL1aoAlqcCOx
vXrUxsBM8+UkeDv8IEEDGsdlnKzqr0awNZBS9/Soqxi/qg8UlBCen4LT+A47
GQZLIvgnEYs61COeoW9lKyPieOyc/lELqTZ4E2da6s5sFbWPb3APGk+JifAB
a6i793hwKPvZILjEBtlisVgH0L2F2bybo/83mRaY64pKn9Zvy8JSYlfNn/Qg
EGdmG+REFDbrkKBvFnOzBixECbGAs1Z/YPt6Y0B3UybJI6w9dkvl1D5iQiRi
bE6Nad14bvVb8BTN8ferS7p0wI43qylHv14d9U6GmGC0VonxLLRbaXVembDq
VKn4ANfa8+90WzjGBF0PLeuleaqxNWR9TJVRs9tr8WcfE6Is5dlwFxA5YG/v
CFbpHcMlZH/C1rleMHQR9tbxm5uzCBDVeRhcskwopEjjFSXZ0kw9TVf/3/Rk
wCZRA30TYTWTX2WFoTRJtfCc3DV63mBsShjNisCuhM9gW0SOhP5JKHOzOPFo
9a7TH12NLW8mKd82O0Sc/w715DuHuF+vsZTFVMO9ol7tOS8bZs6kCXqiQEAO
wZ/JUbOfw3ROWo/RqhqnYTCuSQT0W4MaBD4vQYLjYPlITP4UKn7VKwdlLRmP
0UO8RXIQUxltiSELpKLSMCUA/xLFvBAOAmdSBLrq0E46DmQqVlTgrJ4Wj3QC
v0UcVkInKComZnIA/a2Z171Zo0iuMSjBk6xdIIR872wtGwoK0ongchMiCAAF
mKyRtkNArKjDZEkZYyDOVwpU3NNJPsN90O2mGGeUaa8vriGCn6wLQYGBmmOE
xjh8VSoVQypH0YHz9yz5Nee6DyJj2z8a+LmWTIljbSBX1RTz+gNJUD3brM28
9AEctp6533MvyHCsI9HsU7jPjDxketMF5gBsIpCliDtOq4OtptUEpHYjFoMQ
xwV+9+YQqw7eBzMlnzxrmR1E8tt4lNSrUFnczE8Jed+encKobAm5yAyOYzqk
DRCEVD9iHnhAYj/HP0hXAOWbS8DzEhk09lCc77lHt31+kL9MyeimsfodXmW4
866BDAUguWqt+0PHnsNzPvHnsEwFQEj0eMRHyAsvdEspLBLJx0rTO1rxAFcK
o52wE4gAMEhEV/DS+LyagAH55tuWewpDT2ArUoMBRo58YfqVZL0ALzmri1bv
Sw1VE8Nv10q58rzkrxO+ww2Ps/tuBWkUZebH43C506f/30WykfkZxbMaWTrm
XiE/uvdPLEULEcu3xWzHQEmqe7XppJe0HBdMuw4TRcnpOYO6wxUaHfUR7Tm7
V1wECg9fPS22dE3u81cmSsHS5Mq7fqPT+bQLu6orolPw83xfX54B7rj6sPeZ
rUipLE2nANw0Tjkm1EXu+kRjmRjMzlSBwqCD8RflWQJkMe3mef+keHbXpkwq
ZLTFGarRep1FdRubXC55cLfp3IDM3P18Ws2Kr6HE6VNd2AcNTaJ5F0i6GPeg
xTNQqTdRGIrHZDGF/8l+/Kc8NVdlsneIdEmhvvl5Blub1Z/jbQM7Ykyl3Yvi
FFSYlS9JOYCspKqgc0xeBQN8DpT9Zp3xcFfkeC/3KssWUV6TIJ46/+OHrCKr
rKtCp9DVbRKcQTWhWth04JKAEnMVYV7xS5idwssP+N5fvH2wZreuFak0nxkg
VoqiJBe0pX9bFdJyx2PUhTgryDCDxhMI9v/opvPpb1YTVbEziWXhiYI/9QHD
awkq3E6/fi/78Q2zWSsImgCA602GUhIGmUy5iThdJDXZiCgBxKKsY9R1UKPi
lDe0PeWjo+clo2Fja+ZtkVl+Bi3gwaHothmjY0hwkFDL4dtvm6lwnnisL8Ym
RlQ2HDawcxGBT8WpMI7bOORy8Kw23t4LZ7V1bdG+wzPmUdXDQDwM9jlaTLU1
G5gl3Gdm0lbk6HC0Wq94pr0QEkvDKfIXJOWLfMd+wOOccitZP8br84bmdJrI
yV7L86kmp5CYSAd/e8jeebPlrsXWSqGpOVE8ehe51KDTzyCa93/+ktnWARl3
XEjgkeDD7c7Qsv4mDEe1zLm7wM+xh/6zof/f8Yeubj9RW5NVd7EJwGvoVccB
6YkIQzCiqs54zy7UUG+UhA00iZZALfwXQGUUjn41yXLgbIWB9vqSMXL0AsK+
Bmxs4DgzScVlSWLl6DTqU5gzxcdLDftl7glBXE8lFkhfJGNPfqQMaIqU4uiF
FEMzTm/6K6n+IDFj5qP8Ym6U64BXml7Fs6GN7zsa+sQqJHRir7/wp3wFYNhX
meW+c0hh4KV781MCXodvEGHhmB/HWOwImSXqiYP/z6O+5v1580pw9lkrSEz8
iWXuuAkU1bRxZKu/58h1wX1YbWP/sHa4gYnB2/un5bfOBfUNxrurqMsMub3g
Du1GqwrQlb6xMRwbnZE7lPUifOG3YzosZ8YKBPTRsouRHMAB99PUrplrAjCB
1MNXsq/SBaPPtnG1PJZBGRIfYm0IRAHEz2RB1ylyRle5/8cdrGgQaUqRKisC
jEXXyR/DCwZA7uhpY2CO33KqxacQ9CmgZ5pnBuA5fjWWDHufQiCJj44u95yy
cW4Ne5LmtC6AIY7xfhKeNSvShAY41TuHZ6Z3GGuWQVeZ52vRgxed37ZuW7f0
MvWSTepWH0cF4tYQV6gJSQVgT8R3uOsazkAQa/7HecyL6LpA5GuWA3udWcQ8
h8SWA0OFA6Nf7r5tlXma/xhUQ7MDtUuiXtvucsG7FrP2GWphrd5vaTFerCr3
JEWd5SQvQuOAoffWflcdmN4ecoN2EutCaFH5iImbWbwxISJz8fjKl5YY2glk
uCDbQlbG6NZ10pS4CnpYtCGMBoddoUNTiDqyO7edBYOamYbpzWgRCzFj2cAc
Coy92CyI3FGrI6QMLj/Ly7FXVwRrf2yymwbKxHLH+eoWPYSBx3Nc92NwaWiN
3N0P6WaXAxBpPLZkybKU9Fk9bKblcWft/7PkrlUXzKx8RDaM0YTCAaC2GDRm
mjPSO09BiArxURDa9+Vy4UPr/tYnwOi+wnFiNg7GoUsVFQlVvj+su5cc47XX
eLvMjRZQE3smmu637ImBEBBra88mDO5XeyAPfqMQpblyWm34BkA3uciopLTc
cnnWKgKMisDOwRqOMoT+uKO1YlM4xnpPCejEQNWMmUecqOW69RLypkRo8aNB
wTKgckVvKSLhouY+FvBd0xgSbsJYLauKDS3Z4R9QLoCHIS76OdAh4rEppSOv
Dd3gti5tCZiYvMu4pSS6bxBQEDoFhUOC9b04Lpkr4oak2TO3l1cPUtG0NfqE
BeCwsd5Z/56SaWozmJo2Aq2Y+5/qqpUt6pmL9zZoeVXBriW9sJhZIVFDGEGy
TWmy7+xIyC3cy0PZeokQNB5Rv8NVtF+ZZCTFem1y75T2ZWoBxS1EGPi1w5e9
Qkn34z6pRLInhyuElggtYAjKobSax9KUSI/XKSr0EhgfW51nVx55M83nshp6
6Zw6UsMAqMLtJA+gM5Ix7Nwjmd9Z+I3gAoUg6atwb/Y+RE2eMvtN3T1feOJc
MglkFgZvMTPZPcK3HSNFlrPB2r9emEk2uqgLXgOjTDOupHjYOd4nWYDsRS5Q
K8lbju4KLswW1a3L6TWOjQWHCkYhF4aTTTn+ovw5Yldf0nJtt8PhsRnt3Uv5
XTRNfqcrdQw25Abc2zJAC3pMN48UETOWY7NHNp915388NuDHatrWGit+2Wb+
wFNY2fBvFnRqoSYfrf2LTJDaDsB9diZ4gs7T1nl2JxFvdxF1+kLv59KWDRvs
vbWsbMQ6emevJwa124OlWkQMKiiaKZBli5ll5RMR/x8hFFDvhXMdycH4J9ev
NAdERyqf4fUhk/wQZjs3LwVxzzv6+E4OxbVNq25PUOSBe+z6c4AjqYSVee8Y
xqWe7w56dmCu9Wxkj6HxJHmTjidl/Rff+e8W0Ottahx/abc7QAQaHOkEkwhO
+Djw2XrT3ZglJcImCJcrFyyuoUDK75YlWpdNYloYfQTc4zjz8/mpe0XLcGEm
aYf3sarfnDTVH6iZUKgjVJcbp1aXHF9linmY4avLKzVG2ao684Ahcxf14rQx
F9b+dXQ4Oi+D5/JnpBWrBXXkVBM6sGzgxzflRASwya6aSk0YGVovBOmkgmAC
+eZYc5P57tFnvBPgQbUDvhKO+TaIktVP+j/ZH2raUMM43w68/2krPIdDTNIp
rGKIAzU02B+yyyxj3RquqoPXfuunSklRLhPoAi09aN7/gxEBzmf3JPdH0YqP
w915Ir20G3/wJU5pskDVXV/mQ2PA9MHZfftDLL23vJt3RixzKAdIDGl22YRl
OdcwhhGLbSDWp4f3zmCBOj9lxFJoq4pdZbJwtrOc3nmTNyIVfVqxQucqqBp8
SOnkAlaqo47p2Ai6KVF5LuSQn2K7FZ/Y5paAE9DtOQcnqa28oLE3f8tQhArx
sg5IXmPU+FlnZVTcem3te0S2E67XCN/+0gtaLb64K2JAdMD8DJ3Ck7TquyVr
02WsZIL9DJklG7a6VDltGqW9zHkC6G9yBxlu2k4J5OpRf+Xgr12pCc0veCQa
+UGCXGuX8xvzh0yM6iwqRBU8AZaUDgoVlJ9YCZG+GUKeF9zVnKzwpGDl5/TN
EdGFIOvxbg2pBMYxU/uh60ei17SYs1lb/MSULVRLDdFBulT8acHct+QZ7eKx
tVo/doYTbife52EgNFQabw6fQIB4jI6xZB8Z9WFPRZoRpxTtbQx4CyBZJAT7
MdXNod+rej9nORoBR/puxYIayZn9arcAFDNIGhJQ5YAcz9ZJt2kY+kwwbSwY
Pu44QLymZ++Ve0HyrEiA+VWeclxItRlGouXDnsTIY6PCU2kQVPq7to8zqxf4
Ysl0tGlhqOuI+T8UBQSzxpBMPCRCH2COfwjnDeKaPZNcMOX9KnkOITF6WwU3
gWpQAcULpsBIeK00t2GZCYNJvoG2ohpruWoGCXrZ1lkv96lStQUdd02b/+lL
Qvdq2yOLmqF+u2SAGcsoW9QlVwX8G6F38Je5cm51AJjqVniZ8Y/50LQvo09v
uLYPFpNlrhrbF2JKpK+fTEX8EX71JGq5JP6diMsxV/BkBSldPII6IrLPjPf4
2RScQ6dd1oeeDrR1tPWaKGITKUECd+zbk0KqrmCTlL33oE2SI/R/nFUaWG3j
/mNLldr8K/tNro9fcXk9H8ZsYnxEQ7YVXNEEYbaOFcdf24EawhsgZxhofHxl
vWxvmgmobMVUMxmsKpJsupRxhj+K1zyGIj8HBmFkUxYSq40witWhfGfENr1S
lSYzoIWSCv0e0g+Yq8diTsoUbrhxLQVwnzxKPfKb/e7I9LxAVcpLKFn4YP/0
FK80BPdYpa9PnHYO9s+RSB0n8wnzGQRE8/MAtyOXT/msDQJQWhhyc5dRMDQu
BrbzJ/tCuQTvQ8GfcXJcWSr+bAXxQMqMi8jFSHyJeNcM3XlP7M1zduyEonns
9gFYu3d04j5LiLgWl6TGIcr9mqqXEuJe7v9qk1BnkU1sI5EePzl0ASmlgSkL
alnyK6+rNwdUb4AwFtUcjIU3lNRFiSobT6hiO5iLCUYH7r8Nzvp6rNkAfoqX
Gda3NUUTm9duWmbe8QmTAsbrOzKmYGpjE6wrteDDfmWtgeKGyYWNqV8Npw2k
Wo2YFJGfXSfXoKBInpuGba3X54rNx65eZhBJiNwhUCz50cDjLmdZDdaNmrDF
PsKO9G+HQH/fY9FrsZXaJ1SFC+gmmal9edAxUsnP9LxE2WLiJ9ejgXCfIEwr
lrdm6l+XHjDss8oPzKeWrQAiqAA6rQWb6YkOb7cARMPnXmPRqe61uQKYyP0h
ucn5iSt5zoQVX35ifPJnMeXYLWmIAy93me/lstJbDOcaDSj5mXzOVQteDtcu
3G5Cr7QPTi6ycUk6+J/M61PSu/HseGHM8/9iCTJj/9jqj5ARc3tr/uzQ4blb
KH9cdWBSy/gBmXq1J0SvjpOpuYGE+kfutSbrDQ61k3oNTcOb86c4TBC2TZN4
HSXdvadcV91pTk1roKSx66TSFr5uqrnitArfnCsb/RGAbp6qMvD9vKa1XSXF
3TYYnP7yT0iRaxy99CL4ZHqf8hvVYBwyj9/3shfDbWpnvRGdRXx0Z+6/m4cP
WhkqY3yBdJK43iSEwd6pyUleXgAGmAhA2Er/HbSN1pm39asyVjJ4O9MkIj8f
xkgDz31YbZtF8tUXa29HNHR+Kwa+LhyC1+sH6vwi+ME14KKT5hMi2cNj8zHN
4andOjEIMlGZQoZfVv9vPCti82x55D9mazudw4nfwWtgbsGzlQa6uMkkBMh5
nAYanMxlqqtTC0c4Jjg1gWMIJOkjhIX/dqB8OZOph4RWEx0NAYRGU8LkWWLO
NXlcSNDRQqDykDzuPDVfIVEigZkMHOL+6TUkj2+0ao3IaW/iJlgAsCKHyjFK
GrbeGikQUWvvy3W7YDxibJwRrRxRsHHM5MHTEcBmynEETzsiJIcJKYUu9r2V
f8vevkDE0vX9MzqthKDgpwSmVl5WgBpN5HcMhB0vzn5a1cJodLnuV+kUC2cl
dGSvB3EyAsb0B6cEiGLp/z9C5Hsjn+xj8rieqnmNtPS5Oa/T+n8XjpetOZnC
/4ryrVpAh1gMmdgLAOKyRuRF7iutdQD5/wMlf7OwJrEyHOQBhx7KkB9J8wTf
sHZ6RdXIsR6AjdzhnURS5sP1lSDmzeTeYZ/Xkdqb82xvySXf0ZWuq/wiShTs
ne0yXcioUkzDCgp/sCPGDy/6b4g9+W4KSXQoI2MRIkc24aZJWpPcor7A5ZB0
dljU8+o73prPLlmfskmFxWsB12hM6vdU/FrXJ88jGqGCdeQOBlCxvadib6wb
1J6F3Hhst19PB4RIWP++huTRUk4czBhsofCO/nj/u08Y1Lqh/wV1Nurx/+ig
wWdRxWlVhlkD76c7gF1awLhlI7dZzSDlOryXiA6nvFSlQwQtKTeCT9OD1j27
+K263v83sxkiRx3c+BhI223GIW5rbHIm20ioOQMDtHR2vBT/m5COlERnz1NK
yLO4d1INul6U4okVus3SGfI/t0eoSar9M8yOlkjHXIWpifrB9fdiHde5TZUJ
lFVwoSKhnu1izhU9fa//YdpyREFaP31ghnySVrxgV3dqumD7Nt2SrU38W3Bx
+h0UpAytTwOf0GzrIrFi85V39DPmOJY/ueNiOdchKDA6PRyQMezo3GhvpTYc
ohgMrQlZZdJPkBH3IUAbz+g9ibXPlQRNWLUJaNxJf4Qyu7Jay1BnxgMFKnyT
zEuPCGIWy0pnnpjvpg46At9/+kYQIkwY/G256BRiiQ1kH36trOYOqvTuanpx
jQTjM+ypPZCpnZecPh60gzwWH9HpLjG7dP+mSWUv9WMaZUWhgSOKZnGwjUKr
eBGoCKC1p76s5lnLQFk1NFqfgLLfYEopIBxA6J9GU1hJax3m7zCMuFnUMJEp
kpUyOBnghkZkURE1nD3Ap0WKU+y4IoAWzNsxkN7FYWsMVMf5P2ZBI73l7wEU
RPAzjMIzquy7LDas2ySGxpdsdpSleJfD8BbP7OjE9LIdZ7aHhiu4/+3FmZ3G
eBcIp442U3DVoXWHm7x485YQFqTppnOCULbMTsGI+3U22XeJJDuifbU+w4WA
mq88wGxZ1GXPcr1OIjMn0RYYspLuUXt92+njoJh7ysT4YcO0tAjfrchla0Z2
upPXWVZfZG/ycPPClPbCX3c/OwdgqK9bCJ5EBOUytjz9KTyaGCS90mZf8bKP
7NpnO0mYfjJcI3u4vJw1DOAef6fFlUuDN3efQiQ0i8XGWjqwXYYUasqpU4gL
aliMyNOQuOOvcJQMRQYGOqBo9q/jHzGgOw7mLqpRU1w76czBiobQIXPGjxoG
1GD7Q8cbV5MZpXt05WYut74xK6QQXJwk49q+N7xVfBhIcRazWS8v1HCG37Y+
b6lqhfqv/9KX/nu+p5hpf5iV3/8gcsA+6gatNQ8P1i/Iufrclizn4Ny/5mx+
EO9jGBxk79OGq23tAkzEDDaSmO/fXq1avaDOsnMLqD2AkkYGUzrwpt/SstSf
CTmhVDfIDIyg3zmUojSa5SJT/CSwkQg9KMF9t8HoM/mXMhQNVdQHntYxA32r
UihQ1hjW+SJ/em5FuP4f425B3dK7huv0c/IeYxhjj+0GiQg3vUZw03nSolqD
Jb4grBuFCojOqfwNrgbVGSpHAhlF1cyQAVdnSkeJ5k5UAkc+4Ji/gfSu2gjZ
ACVoYc4cslC3GbChJYsQ69xUwNgHa37K69Q+/onrqQse5a9OVi1UTVWIoxUI
Pf11bimuqEpPYC3bIvaQ9uwXr7eaGgpgVgqMp72bz5jfzMVgyIfcARVxAm0a
5xZb5ATbT36GvyimSQR1F00cbkkz21mCu3CPOk/Tx+4+EPudhE1HcRP85Jlm
hFoxFTXeyfltRASadf/kQ0ii6+nDHWk0tPglaps7JBxiOg3CUUC9kEYCBBZ6
HBR/ao0ddCG7HhXB3Iqq6AnbYO5sY5EQkYdhtTH2eGQOy6pqO0iDwhyLBvUO
BEcaSa6A8rhyJgz1B9PQc87jMvu8OxhvUrD9ZiDRKIx9oIdS83UVaBQL0F1l
+Oiy2uZ0C4HrI5/qrcdt9PwNY/d83POfveaX+A9RWDzdGcqzhmcekqJYfEd9
UtHXYfzqZxEUPtNJDiErtKJpAKXE/2tW2sXrmogrxRXisxSVuFRDLdOMQT88
hVHOPzvPbrfIsJzgOvraT6TcDrPyIk1N2FRzR8l8wl5G4n69HsJOWaLqWf06
qcD7A/e80ZrKvEo4NOYRIFqRqbm895OFU+zrbsGR3yHmOoLRO5hFn0zRBLuQ
OgQf43sjAmTau1+Rsk2hgbYeCSLnn/sjYhR00tsC1ijvESZZ4MWcCcEoYKll
yULk3Kh+s8V+O8uZjzicAYJajA32KPp8LlOXojwt5g+3fhcG/e1J7K9n0jSz
Qdvw9dC4D/uMRKX6jSLiXk6oo7wNqFTArLVVVJqe0+cd8pimRsS0jdSwnOQk
LpSD0Zqm7J0/5Y4+7U5W83GWJWStnMR+mc/5e83CHPgyAZcEUH7b50iMeE9B
TiY5I+03xU+Ak1DsCIrvOSyo168y+9WjmkcAl4U7JIBl2WKq+vO8on4naL0N
9NX5Jd1EbQLqbLysC83s6zSZmZyBcN9UtEby3GzKYAcP+rC30eQVkK3Nz9Ed
Y7v9kiBM9GRZoxcDZB29lqapFnVOVxresrMVXbQapChbPnYhGyqE2zdZJ33n
JkTZ29p8NR7PMdIbkicwRHjTlFkk0t6Hf678CyYQTgCPQyfJYniEOKRfqr0f
8dIf2E6FuFsYO2m1dF96dQA3LTlBzxN0fvd8G6PeD+dq8sas5Goms2pGQaLQ
Mnssj3u/ZCQ+svjWE/03wG5i7Lj+PW57J/BSyZ/1Q+YPHwlPm22bHSGYXULK
R6d1tFZaqmqCsJZSQoZk/8K9TavykXxKJJjKXcdAeBirxahY+JNEcHcLI4da
lJOJsYNlUqiREU3KPrSoGbjNLQp4RZuA7jm6MX2DIvL9CyhKnnn3B3dx8HA2
8FlNjYlrqHAT+GizHHbvr0VPzExyg7j2EMdsyzoiA0BTT8W8+h4vEKZv3XsB
kRpJrmEOhbm1lVePgmjN+c/8nSEK+iSkk/AtPbla0mc2H2gqqfBkzAPuORsD
y0IUEUhb1jB1PUBVF//qDye4nj3h3DCB5rswshcOzqT3q5yzw80LH/aBuLBP
tpGCkyJAN6SEu+jYy6pIN9XnsTaB9vQU8UGTZdnPnA7qGrj/OLGK0cxAdiAQ
m5XFt1uuwM4jUNSaA15LNffhgApOEr+q3bMX9VJ0fGhzvimvUcVsvox59ypn
9gKwl8XnsI7+50Wxls++R/DnRJe8J4UErhu0XcCTNmKyhgXlQJcJwAmhAGBf
WU1gedoQ3F6u0L0G7R68eZVuO6EzFlVnfwtHX9ZDkgf9kvJqfx/Gb1rqZJ3H
ie0vUIKWZKVu3Vcy6RWe9Pc3cJ/p161bBuNz2/3QVCFcVWR/suF0bF2RN2DA
0hCnLaiimvi16Xu/B9WiX7VlobqHKNP/FGiAKPSdAgQ/c3n4+BUzQIFuTbRj
7knPTeG9SYPYYKP6aTAO0OvXrLARoK8aaYnr7dRnlSUkTWpBmF82YUejYNbf
QkxJVEvJs4gLXyfJ6I3c7qM/dpVr8hoGkgSmiygAi3ReRmXFgADbBwRe5w5Y
F4RbVW/s603bYN1/qJCi+YWr3XlQqZkG/n6E4z29x68u2IauRJdoB8PKjxyD
ItiRmHASYoU2Lo1gSX54Adsj9j93fjypqWH79yzgvGNOWi7dg1moakvfpHfv
2fcO6HcU0wL+fM8o4bKJhGoG5IfSYoJZ14qA9p/wgfEkgmsr6THJWhoPA0ZW
3EOXMgZyIYJzx8zct/YMu8F+IiYiy3fkKLnsSpjtP3KeQWwoK8usGnBcy+ca
O/B2bA1cnJaCh0igwkonnRXSUOYAMhKrfHdxwSjcEmyKJ0oXvZbVftzjHt0O
LJvAZ02WS1BhH2P2NunExySwors/4xfnDi5Jwsz9NaOIYNKcm0td52NePO9U
vWNoFm810NwpNnEEL8EgHbyfrgeceRjuL6jqjKIIR1IJxQGnt0oDtUdgTWu9
hGJGj7xpef4CGWdDtXs+iMEYqCDNoF9ywm9jT0Rl4W5TNLpf1g/8tbGLV2mC
0+xbYLUnfXfCClTuQUU+C0syg92AVVxIPUgCNzlL+wy9B3QZM55IdYgpjG2X
H0NnzG2DJJKCzaJQMzpqMuTjUnilP25q4FzQ5KVo4A6rqsNwFdW9zK9sr/gp
8YubVFT8DELvmMdhIAd6MgwquNtT8M6SmKuI/QYzrgmsMqsZluFLE/R57fah
fa0AuFGc3HSprNoxgWi+W9M84NkU7LGAJ90QJRIZ7lLEYxzPGOaOVh1ZfeKg
nSlHSA9YTzVPAtE+i2FnCar+6fjz2NwOs082OUCXH1fDtbpjUIKhVtZIZd2V
Kggu4jCp4Ygssgzi8Mu3eKj32rEQRB32ANQA4++Px6kUcDDL1XZs2B638G9i
IPE55K9mU8FzQkSuWTw7dtGqcp91IAT6ivWfI/j75Qy4ZnZirkrMcZAl20Pn
e47jFmHtNDM9klsWRaLJrDc4O6SK0LATc7/DXTaOd6tdlwox+x9HmrUw+x1y
cR/WX0w/CvoVdt4utoNHdIp2bleH0RBMtFPC/GPwTx5gBlpE+Q2ZElasoq6n
T3uoiDa/JnDBm7zeLHSN0t6EsZPOUjlLQD9tyg87t0fzbSu+5B8m/omYIe1k
lGrsC+1U8a2gP06+2W65U8jDeozDNkpzKPSv8O/7Sj9TAkxl0XsjpZxLT55O
NIEkktCAtWvWLFmDRNcMGT8j6GvjcE3B2UfzCHKflio2zjDsAXf5/KCewvAX
ihl64Iqu7ARed/3jAK9nMkbYO1u5GbteGj5xe2e/LPWR4dT2+sNPxZ3T+PtN
cAdCZHKZzbYVRlMX9+IDjRJfgChJ0Zt9SS6ddBv1IEyZ63QAqV7RoCICLfs+
AX6t9HyKGuOOLR4+agXU0ANeOiVvuJ+anvr9pQjZ9Dj/Hr6d2kL1ZwqO9edO
QzYa0yE3ipcdYi9T6ijvj/SJcpy0/Oy5spERxvuA0bxzC/wuEE2sRFe1lQ/m
ZiikTmYfMmYNNaYO3sRfYZeU1aqGKHLqECre7qNd9vj8bM2K123B7WJ39DD0
voVfiVgJxDcxd55jfPoOzYhlgmg6UXNDPX8UGeAuE2EEMeouVxC4HbP56w/z
mnObZMq6E5g+6gW7VEPGKHnWg36DWyPFaVxMsF6so5CjlsotbyD0YrMzy3Xc
QnoUknKT2c/RejR+7814cT0OK1yyhiEom9D2Idj9qQ4B887sYWx9aAJjZjbi
yy9mVFUdtleTVYoh0E7nIh5QsvljK2YqrSFN1cid8Gv3GJSwtpeclntU1mm5
hr2G5uSYK4sPodKil2QKNq1b1GVx7jwRikMIRe7Xu5kpWEm2t7gFJ4aDe8PL
EQtXB4FaMPHPgnGySu/P7zAslu1vwBUkm/mfCElKZEM2daTWumHrBBxqb3uv
bwrE+P9BXcIAMxQcWFuNiZqqGcupKOvpyrjg+f9rK0XDJmM53eQh0AQ+rrN2
aoEY699CuaRHRmWIphgH2q7h4e0H9A1uE7+ozx5MYFovWhM8ZbZvIbApK2Kj
nYmW8/xcbYVh2ho/YaANylFqdYKC37VedZ1U3ZVuorchMUC3M1lLolPcAF1L
3ytePINxQPaTh49OYtyseNtKAufdGSNVaKkkeI5EQOF2IFk+rxGZDcA97ilV
io98oK3BXSJezq8BpV5Dd8gx2askJkFwj+D67VNdi/umPhL/JUW2IYC11XAC
Y1L31OfE/llt3d/fTd+fhgxznR+XjrJxW7YgNuc2IbwRhfhsyaudGIsAQ6rM
OjS5l6dfaYElaSBSgB9hk+0fqJ6OEoFH53cZ7oT8FpektW7me75AC2gklmRu
8tDMWnwt7/PCq589OTQ38jq/39fuSrqheGuDPdamfCCj2jJy6Wbe+xb8n1AR
lMLlX6zg49FS/9HJB24SuWFChUxG+zDXlZYc1YwDAKGE+wajMmmZawN1fwVI
pOkpqDukhdm11ZBPi71+UTYuznOjvasKfzEGHR7RwrMspgKE5MtFjmg30Fng
ZKiZs485nmnycoIAn61buoIqZCmSOtj+n93z/bUj6Iy26pZrTsyoqopx0N6W
CVEj2qJOf90IJPAIQf62lokhHzS8edpkQjNPBZdKtsJz9SRTEMIo8G/W1dkI
W1TlgDzP3Oaw2v6MPHXux9+UHCJVACe9GiDgqHTXKd+g9xsxjpUN0icn9ecH
0FLcULosBwfGgAdU4h1YSLgQHTZg/PeF8bYLr2q1NWmxqCgRH5xKBG3vAirV
btHD6aKciBqpzcqRqYRmCB2bNyQMYBzkdEze2QT88EEDawNZxctwmm9/FGiX
zbtuxsTrSlPqMyXPr04vZlxSufEhg5Pq59dP3tm2EQ3qxPB+chhNlIPbhW6H
aO2FqrnJu1a9BNsZ5NK4gXCVkvqaCPBLF0avqXu6kumE+aTlXT+KudBCH4oH
ODUv/XIgkl9vycMcvg3sZ0GuYE+NFHn8g2I8hqc+hfDrVj5Ed5+QQFu2XpTN
2D+y5Ou7q3qXZdMoZS3EM1bD2HjH8la140jvXZuBaV1rx9pCvdAYCCI9wxxh
4yIshec8p3/A3cEP6HP7kY/l60amL12tjmTS/QJKQb3yMAZ2VaepaqPUEgO2
XhQRgWAcdEK5VeBKX33heAdS8PhaPWaiQe/1aOqsD+Ua8pviEAZldt52K4i4
YKNkEikGTXGJgEoqYu5fwe/CTLBLvxBv5vMRY9Zr/utwX/p7Z0k3GtUfDTtY
t7GYalhcMYexyIkCHuI5j4pD06gDDeWybImyZxfcmjp/LYbQlCd9/v6pviO/
ibMHw0MpmSvTvjR/wnxQqVf4+MIOvG9IywpxbbYeewQhX8CORUoYfr8wZ8BF
upbSvK9Cj6MN7SVt8b6eWkAsIlnEkDAM+zRvMzaHrfgM79GxCX6An1HMP1Kb
9LhayyS14yBey136sxwiFQ3hH8cncEy8VmkNT50EB340dYSqnrpOFDgR1iiN
GruE1+wTto7Ij3gIAKaYeu9d3CrhoKRzzXKGqAAZFdbwuUjIh18Fp2HzyzM+
iEl1ZUgInmSiDGAUfdwdR9FBhVEyE5UXxKoc3LXwrwp9skAhvyGQS/38rwqB
A3GWOtN7tQXscSTigPGr4ETspuB84xwxJIi6g5LTFp+Aps4PtyPq9dbnlBbR
L11iakXNIeEciY5x1QaRlFgDjzD/WvwHidR4DTu/gEeibfqy/OtTuSdVeE5/
EMq/v3wy80iYTg8KwDJ2O9i8MHyqpAL+jc79JGe2J5ymdf4hi+QNyXfIlso6
m/JbcqHF1FIY6H7Rofyul3sEq+OGk0G9dKGCobJHkBcl7T32KNHlyh0uerAv
Ey04GNyJ++qU+31JrdZal7LDGjBI+0cGvZ/w7f5diFlh6B7fwTdg1qkTQTkJ
5GLLseBdE3ahd4qkBujtMKvYQPKWVMNhSyL8zbExZ1aVJ29K4lBQXljZtsE0
yXuyPvG3OVTk2s49WDXG976mc5ZS8U5sDyff6gUnXxVIiYWN+IHer07GipAB
5UmIIPIt00/uLx/81fmgrwmIkbTKXFJq8VM+sArCLXUgbOL74ZonumirlkzU
AWpK/xNydSqIklJQpboGHd2BTPCxPERY58rY190oLb4jE+lm1+Ogmh3M+xuC
dVonV/z0KDchnDTTqQOZY0jCDRsfnXundoEbPOxyzBO1+3ggaTsMFW+EA1va
nyC8C1M/EwwsJ+l5xQ4f54aWw/y7LQ1tfyXFnWOSu5UTwUpN199HdnojJpXJ
cbTL0WcDYSjmMgNLbiC9E0vQq7D4dfqBYxRC2kaZxSipZav3s0ZgyDFoQPoN
lUNUEno0TP0wtBwOZP1tSt6aB0JkxYK5ewK54e67QJaZcbZH7BZffW6YT8By
q/wdWU8TkCUtInmIjMFtAA8nKluoQF/Fm/3dg3MReOGgG4VaiUSdJgi1yuTx
v7iEp4w9m3gzrLVk6nmN/HejDuyctHaCc5JiOvQJ5RwPj+XpsLEYGTp0foFA
mieoGHFf8EF7MitjaRxY5zpdEa3x4/3w4TyNQmy+z3zaEwTa3+14vUbeQvWM
yUDBCdmwjQbX9ClZhiOppYzf+tM9CQQ6+n7n99dkGO0jsMgWLu3JRx/EU9RC
oYUKt1+kY7wqGjNYXgqIujThOsmTdMVvSrg8aFbYgq4lZmmRxALNmbr/CntD
V4N3q64Yye9akpY7kfkE2X5OHneJWnv4+V5LV6UjDbJxRVhiBZZFJknnFmOj
B1jELFm1gjr52ZM/49Q9Ko5AawKi4vY2KNrGt9rTAb2naf1GVrUgsoILm51v
Yl2/N7CtbTHH+Wcjd1etBlIOSFG4YqBUMCal2/9+5oKPJp6oFyJVwBLqG3Tq
y+p48x0AmMRQmbhg3S1wzJyF+QeJnKTerwxFZBoKhRQzjZF32TUdVv6xuPdc
gs9mqchavYfBo7HpL1ru0xJ3gjH7ltSisW/SM2T5tp0vC3IxH0rAOBeKyqA3
Z+aOX/MnxkKDh5fnmptZOQ0Tv33lXxzXo+S1mt/Chk4f48sP1JRuANg5qWcf
99EAZ7n5mWhWhgwGwnElAI8OsUx/fLifOCWD3Hp8GeqFjBXBqkbcbdiJZELU
7BPmi7veLihs686CAWKB7HCghhTMibCB3UIqdF7L5iKLnFvnAlXeE/pE9aTk
RmfhQcuKhBKRFr6nd/Wa60VWDeTd0pqb2fwiyMpLRzGmLp/kBo6ZE3AJiK/Z
5NN4A7n1lV7C/8FjsMyc6rraZ6oRy7pR/vtkplWqKbBvZeojlfGLCqCu8Jae
aOjlerrIMYuSilanywHNb+Nit5IPfumUZzL51K6gfL+AQBMMwRORkdhCj+oY
zrBn+7mPXjCLFUfk25Y/BBAfcR5Tgztd6d6OHDP8OyTZGyvt3B8MbsmxKW1G
pWlB3TcoAWGP9hmme/k8HKbGC9LzMTUiudv3lyWb8PK3JP8WouEgzfJU7mjq
kGamxBD3jYZF6+ZQRyhmM2/5+zYHN9+U5PMS1d44AZmC5KMJVpzDCpih/ysK
s8f44WrK42cuS7jg5lb2g7mRkJsTxlyv+FWT5zHgMpQCRE44WMNVwUj8vw/p
TFgitSZdybHjcK2Gz4VNgQDc2izpnHUmYCUR5o86JfArIAjloxW0VlerzMWY
vAxyoaMSkhng18md7NT5TQzKU80mnClJNxsCHnkcwhQ9GCPhf7lrChUdQUTy
pRFvYH+Iv7nSi2jXWWBPh9z0fB3OVkGxLEcgCI5XtePGvna4giRRRxKNkuSW
jJMpgLUsOb3FkWsCM3E9PtpiTXeDftB5MJpPRxJyCkN69mxN9tAL+Tb42910
6q2CJB89UaMgiPepf7qHHCDQOyuBAwNdMepXM3OKp+cSm3G6qFy8gkhmADXa
MwIKe4YZZfEtN2YlOmDml7tYU0v0t7uXbKhJZlhxlBSlqeGvCQi65HnfHwgP
B1upieuKkcv4cvVfa9laKTp6X+4JfCzN7D1j/Myo9K/kjwv+Vhxrbf3XKYtj
XBKFpwnh/HoRROF5isEDCtw+N8dJf5nE1QKRdYF+AI5EbTKFhXsluV20z0VW
Ed4Z5o+v9mhjM0LUT3dMBe87HadzECUGBuryLGWFyhJ5s89q+becGypei0Xd
j1yw0g07JjZl/hJnXovAZfXz/SPo2FQrjITu3HaC1a6lWS+ehxDMHaSOheOM
p02Jv8Idod9IrzRKJpieKyp4KcDDDwSkndubvtuzw9VEZpfEa5mZRqCs14Vk
26NY7G5kuckRuhPL3Y8A0M9mlUWRGuzVJOgBsGJ5J7R6NpBkez9vcx/yBZpt
nlzxDwejc1EzYpc4DIS3LqiAbCSlaBMpu655FNtwe6/OKfdx1dfEmlbs7UbG
8L+ekqZlq9/rU3qRK1sEjQbf4uQ2UISINAtFT/i9CBPAo3zUPZubLYFARtCU
ewOEyIjVsQp09AEcSr2d3hjwDq2RfogscyByfuza4DQuGmTFSO6iCBJA4LcR
NaUHVTSCPdCaQC/KPph14Y2GRu6ght9PkxluruVBvMHhp3IZ5IREGUXkS8bY
g0pnf/aAioysWu1moExTxIltCuhDlExvlVSY4Po3s9s/82soYJ2cxemoCfFO
KRDO2wLJhXUQUIN6SSfy5AndKaGSQwfqLT2+2EfP3GBDB619j1AjY8876eE5
3qqXLuHeLRjkfIlwT6GxgNfkzxcFmhb4VZZv5JAKZMj2LHTdRIYNEwCsC8qk
/iicNnThhOlokBR8cc7xU+l/x7cndsdbyMr/DjPUkmWJf+Dk004uy2CmxjmS
CxeGDV2q3bzzzmGmKfddbZ8+ymQFCoAVsYGE10TueLYtDKpIDcu2vrbMvE2i
3Y/76UTkFoy2QGHVobvj/6y/ODAN1msNK4yvLgBoKaEaA5x/PbGopnQ5eUW7
aEu54qHgkkdGJK5p8iJ+lKXxY9Ma7SEafn4bnGsbbrUpEeDsjh/2vSNNNlmm
tbL8BIq+k3RHSKSt+IsqxJ8d+rbvCdW4t7vxHJQ0mHRX8owO9QJnjyaMpHbD
nWcfnZ5Pkn9wqOHFlH3Ut9qi7q9cd7pz9auEI/xGluQtTg+ZyAi5Vo1fsar7
xZcroOCnMr0sdbq1hoYgu26jAaJnWAMRhSuk414q0nBf9lLEO2jHAETZgs6f
QlfYFXCFBr1svZvSmmYBWUxzo+onnUW4daENIJrDkOY8u8PtXE69ZcehAxh4
5qW4xE/ABsWBqb698fe5DtKuIh8gOR39O3oJtMfxI/MLVMPabkZRQ70SPm+a
SejUGrr5H3QZaQpd9YGQ0QNQ0YTF9ksmvxHBjQRsBeLA2D9eMqUE6z33huXp
S5yQ0XbsQ2w0tOINGd9EFgfYbB+GR4YZC0OTUfbWRJIBBb7YanLCpiscBEKV
HhAzOJxzSHh9/jc5Bnbg4jbF12Ub47Dkm41jPTCr60ns3RTm20inG6/0OtIp
vVPt3SlUatHzA+lTr9eb5ZPP760FsG/4aqtpRTr3+irBlRRqlf5Yhur2Zyuv
xjIHpkQzter7oVyKxSEUghvNqwVr/DoCoEJDnVsauAuv0H0VlOEPfkLAvx/9
ES7PiL8n6wHzgPYey0eJhIMeKz53EPe1ZYC2Ddl9+oVTHPg36hwf34nI4rRY
MukXl/VIgHAqzyILiTPJDRxqNKjWFYxBXtQ+BUDiFFw/nSbvBZMWz45SA7/t
DU1AWu7PT2qrnEUSjBhAG2tu9o4kEJN3/hSqL5u15Cdr7oxR872Gwtu8iRyV
/oBV3kNxDG+OmKXRBGr4RPWAX54ogL1LLAjGqCJ6PshaR+WCJI0U/AJI9LNh
UhId7QqnZGwYJ4KF3gmJ9vVj3nTWQsRV+bf9Af+NKCgydmX2cwzUXMYJCb4D
mS9z9XMm+9u1aTYKprr6U3cZBUOPDcOwnX7EtchMl0+hXsbgDGoycga9osPy
4gJFhq6FgdnXYYJ3n2qQXjQvFJHjavRscWLcvdHTkiH7JzTSZXfJAH44//nJ
4+O3ViVwnu5KHXGCoVgHKOdRBWK8uLwVNzeog7eJGM9nxlUT4dRvGTFge6rc
wRibIR8twPXq1u6TuQWVEVtutM4ODpx4+fCm+HvEtWrfZA3K58KjL6O1lwNZ
kP3sF6eODbhOqCLXryYo7ac+87GllPlGkZHYigvMcveyRGJ1np+K/YF6mpsa
CrHuR9RRxssCkZWk2A/G5PWI8UT8AdopIKgi8quPURyawlDvN69hsj3vRYcb
PL+gatLdOKCTXwy/sZkVXVTpdoW4qjGclXNsFFso68Fs6FJ2huBmbeEFldwY
MydKX7wjOI7lsyJEuQ9gVfqjni/5hQkS3JihvPv/vpf8DB2peovGcDgMTRIu
MuLgiXBBsf1ocJnh15CCS6LQWgDKw8yQ6PcRWwWHe4DNrtga3cV+JM6SZ4Rc
7C657Az/+kvCEY1seiBb6x6bi8gehJY37cUscOx4LNzM0xoGmamStNWq7mzF
M6F/Fo5oOly8UFaZyag6nxxrRsUZGHAZEnekkj7UyAmzze/O77LEFR/uQWQ8
RKtIFcO7Tac7FEAZkbjLZLqoqNVCzVLWBCS3l65ylXVN/xt3yz0bfsERABY0
c57Gq2OSOlqzCl4361oEOB8pkdneMREDgU8l+QCVFSgqvrkzNA7rIg1OtZWy
0DzdpLLksl7gf+NnJ+ntIkGkNoTd5huy8ZZsONGeooAD6xb3KXDXhXfyUj4S
DpnW80fo/j6b7Epoqdrihr8WAHS3Ylw6QfK78ZA7OrbOx3DeHJnDH9vwpbpc
wIURHHUtCqz3mVO9c9AeBy4QWXsh7rTgNGPor+7rAOsFR9D8FqYu1ACLwJ13
TIgdzI4SYEb4jVxQIgO8WXOqf6Oa0OxaddnLIdrEDGw9sdW1Xq3lr7Blw3km
ENEw6iBbYZ4JeUTqAPu5ykjH8/iL2YdZPzogY0RCXOUPKpT5GLasuiAxziLT
y6giINt2KIEKTBa4b9g5TncGVRgM7m0OD7be86+PeYd+TsZ25CXsyTQsrr0A
YziED2EtHtuZ6o3RxnEZxHPJRqR8seuhLBZtJTN7dPCP1ztv5qsn7xCz/sTQ
K/AzMG0ghgZP03fkmS81dg4eAUoGHfH2n8QJtzsheu/4pwxakEp0UFJ2BtXq
Vtttmr97y5uCZXIgo0oBfOeGIBRRpMpEd5ZcxoINVRCiCnrHMVqJrlRNz9As
TZOmpznVVPyVXESVEM6U19RJwxqMfFS2fHmIE4UhfPzwaCUXEeQxxzcjhRrd
hbPTWs2VSZ3/s4dqlW9nDQ+5l09G9b3Dw7uvt6x4NZ9456c3hpPUYyWN6N/E
tZL9R2NDXHlgHe/rcOMVASS3cNNyh37IGc3dKykCsubHRVtTxxoP3GwwKsg2
wxYSeLDD2nuksylgCny5E8zVTRv2BGn0XP1TS3sTfNHezZi1F2HmaDwhJPLc
txSx7dHJvQQ5yMtKrp9yNPHBq0IyfJqcFlSfvYdEwdhFDXP0h5DOUNMVjDKD
f6gJkXpfbYwiqWWeuF2Z8aGQj+LzzxuOXlh6Vjuc8tWFgktdx+SSIg6iGGMR
Za8yjhWjQURYJmAL9d8kLrRsRYSAcv0NG880f5Di1cvfd2kCOpEKnyyCF3q8
xnTyKpS+pAy7hLvVrcPsJPmOc2C8/yI/g5smohn4wOBBi2fbWavzXaCfQtry
j79n5cVoaQVQ1zT3X3GFPNhdQCt42dEqb+1dcFAZIw6lv2PPIc3/2xBLVqhc
irF1wUlQWiHnzVNj2H+phrwK57j0xLMymu+WS5TPNzNDSbjyw634Tut/FAE5
sWa7k/GaF2VxyzCUmcDKQCUQ2VJKqD+93RhPaI+JpdcHNIYBy8S3yxfXNRD4
xtW6ZmHaeOl1MTrzl3n3zl9zNEkZ7IXqDQVM0VCh2ZayTh6u25Dd9TEs9+FJ
S1YsUAtmbRVavPFQtdeOC+2iu3+zOemHviiTpLxfTz9u22vRknlcV9JZnsvg
nbn0uVr7m3TdxI6vZOpe+b2ufb28xm8WukOkayG3ez4O+4WVUChhb0MJXhJK
1icSGwwMpK+jv4d6ahvEXFC4Ul1KUaFILJhlVJC5Wr3j5IEcPaBF1K7rvI0R
mf66tnWR3+lkzf/GyfM5Rk2S+tNro6LqfIrv7sVZKfnerxirwU+Dn5Bk85in
3NLmJOl63GTHB91893YC0IBSnzkTFX51huDAXnNPPfnK7YkwB1dlbh5oxtEC
K78MoTvEaYLjPBRF0SH8HcxBQnJ9SMGKokZXGcgamuTEYIApLCbNqIstGQZV
xmlP2Aw8A1UuIIsIYhn7FHHp3V2GUYGaEsdMqUK+xoTLmgnc3Irc2WAnMkKk
aiHL/UkU9AcnRoYXa1nQfFs6zcUavs3n7dqACvjFJsgFw4vLt2r0pJ4FaFaa
Npaag2TTckBOZUUSgW7An/4HlNp4Kxx6bhdZR7nVgTqiQLsxrF7X2wZTe5fv
W3sYnkweM91r/iftxTZdtwLgCRFUuTVy45YCr5E8+l/Q5bPKt08gl+PVX8la
REqQlEs01tD7MbloYc99VR1D06+DeYtJxYfa/aGPvVQpYIU4Fcb+bfhmAODO
p5euxKlA3Uw8bMTeE0VpjwmrTZk5YcZO4hyumhWgTl7PXdA0UTXVVnnFeU59
dUcsa1ZdXxYFQpDVMnh2jNENGTgDuqw5Xhu8qL7OejY6JAAgUcRwTA9pGDXD
vFqf1Uy6m6fAGuVFRpzXol9PT9wMnOHhXbgaGgC1qLBHhkPBY1MMwNE5Me4U
2xOr37ZD7hFw8Y1UV52AjZbR6GA7jYz7WMXGVWKze3fJESzylQXx3n/ZE8Ap
cf/sriBqBiSG5lgldEbz2eNEYdxIsYbm8k6+66BVzPnc2+85aoBFdgCnZSSh
rmasiORix8FQFEKgxgNBXTExiXRnWRbTMV69/rke9GLY7bNm+I1R6gB46Vqy
jVQ4zQ42JZHsPzSbYBdPYlT/YTjbvzCVOy1VwJuP+U8MBRyu7bVQ8pHKrLCE
h1hvBXya0arNTx2kahtJVi0uQmhJ4bTw28pcd+yMOR8EHGIHrKKWgHXm0ba6
GTG7rlPeJMmwktK33LOvpwDsPS7/X9eCiK8WIgCnOQ6Ei3Q4kzYIEna/fuQ8
0Zhd3EF5n6eIBXjShzquaWkTGAl78tqGR2pmFtpWGXAiHHczrbaDSKTlofEe
twtl/oLjIgx0uzmdfZY9Pq9R4rbcGxcsEvgcF/kc4sPz1b+ypXMktZS0+Maz
Z7rbLdi2qgQN+vmEt2aL23tdFfICVCA+hNmnUbh2pP3BkR3s9g8UayHR3m2d
vNPbKhb7nsacaDwPxIZRiQYaU6l8MkuzccC9LdWNs2OUrJLVeFcFbfr9bAf7
z4xojOq+DZ1qOhYnrRzsjKdyoQ4LNjDMoJ2TYZxffz71Lksl3d21qokzcCl2
BEMGporXefd+16NgrvZLEA8OU7rRLd/glUM5ysbh5tJoBvrywPJNOqoUtG6Y
6tNvXM2rRCNZl7HgsY7VuNXg2IkUnSrOSBUd8ZeREuYlojpCVQ+Oe7XOjUoJ
HziCpuSLX0o9B1LcksK+jYdHMSsRkY0lEHBDrlsCbYDpQc+g2DYkNPYbqUgB
MjUCHNpST4UgoMs7WMr30NCZE1JRIAPCg1Kdwz5knq/Snv+Gfe03P1pqyqaU
XOqS4w2O6F1hthEHW4bb9dPR2sHLzniHmDFde4Pwwb37bYMvKxilwTtBRVAS
WP7Sy9tLq5KuAygQt0OaiTWsz22abWsOYzuRhLwfBJsurEqsXuKgE1nFHuUY
G9/CKda1/xB0OGI0gUDMpoQ/FQXoDrihL+pgIrxJN1VZYtACD4OY30bSQ2oH
QAyYYMM7lSQtGigLzi+Fo/n4lR6zW0hr5YQ+qbIy2xwopd8CZIN/lqDHm+WW
JpnlcJ8bZQa666QGpYuP2uQkwPjwa/MVsDGiAzXnx96j/W9VzIpvnz2ezqTF
j2VE4pQGhXGC143ZFBnMcEwkGO3x/xU8aN8Ex0o1bzbczCa+CD6fvlsog0NL
w5g2zjuBmHFLx51AvOxzNsvj/4TFSSpyhKufij24LgBxUoyjHugLsr7I7Zgl
tOJNz6qz22xj6fdCsdVzkmf/uJU3HjBhzOfktiHA8Z+XLemuQx4T+76LMsEH
O12CrTpQnfaJZB7t2c8UBLrDpZ0v1V8w5gT5+kj8aaXzBnjgm/P7CvoxXCP4
L1zj9ynjuwYSIIeNxb/7/xS1nxSG22FobRSowVD3YqjgwphItG8nw5hTRoD6
doLwjFx41NNzk6puyGuUXrFW5YtumzjgRu42xryS39tI8qDWxxNrtP1v47CM
38KumlkELMhjqpMrtdNDhUtp/OtYLgoVb8f5FKsxPSLoHQcvfoR9EBcDGkkL
8AnZbY34FBqSiDc4ifxsjwepGXZE6ueSOrvSXWetZaFdfQfQH9uUgOqv0SLl
/er8GXvQcHU72rIgNORkMAToWiFr4GgMOKiu5BE3MUcqdYOC8VrcDziNC4Fk
OqJ7ZfP8SmsOuqQOlviKst1vRX4jwjy+/yzZIw9F2ZcIctB11vvBA6G3F/xU
z/C8KCqZQd+74Z4nujvsHO0zB8TILdNG/oVvd0Ders8vmPBuC8/ADOkMFpTH
AkcO2+hScM9nmp0A/V2c2NEFvf7m/0rb0xOH0B/qNVt8Z9S3zSEV6zNm/4d8
sARvvtbTMTNB65Ek8c6egfu7QnF+ZSyUBJ1Ws0DNZH6QnE6H+YFOhCng1Z17
Heye7I2IwtUf8GOHpLFuaAoobWXM1n9DwbIbE+LPNKnUwlkhh/LwtemeDoPn
O9B/HhWyzBe+9dN8j1VyWmCTFKDjigd4GyEvs09i9TrwAg9gin2v/kIKrWKn
VU/U67O44ZofxBUvEMA23GgYUwBzGzd6nIhHOCWd1ee9SCuafdV/dDiNYGkR
+DbtL8Ac2HJp18emdZyAYae+LnA+cs/5rd63mOKhpSnlToJ4y2UB0hNr4GAZ
wdmunkN62JQqAZZBtHmUN0gZHF22pyqA0ENfO2q/5FLBbDUOFjoWqn/GRtvL
rKJdjJkN6eHpkFtB4SlsPiI1vuRXLC7rMOXowUWf/30Oxn78B/HqVvRmFxwA
yX3NvKiM9Pk4E4zzet/OLDlXeFmsobCNVgeJ2fPWRD3E6etiOupyPg5ZoYKw
uljdY4FxwtAm7/wB2ohCjkq4ohEVUKRQVmne/M/aDOv3CyDmSTr/yJDecEVb
WyYKNa01cSMtRrcBPG0qsjPqcBrHrHKcM1aneFm7Sy1p2E4fO5AaY50BAMbM
RJsMbzORWo88tkLR0DqBz9QbkOU2XAJELubVR9wChfFs/2I4h9xFEFyT+NKK
96zHeyOXHObTrqLiIK3FZXkC2GC0pHQQjqUcTk2/rBhN5Aa8JHr3RDhiKMkS
EjvyLak8/tUvz6clO3XLi4fd8v0ALC6Sy7rw2Iq5v/32t5B5v3P+MaH41fXZ
I4ydBVYh5o8/XAbNjRKk+hMI10yAZz8l5kGeo2MdVFdGb8KpT8fvczVLbeJe
xdZ8JFMGryPTVbSE5YMFpxy5f2gKDZXUac/T0TGtYzDylSPiChVFtITulb1J
rjbvqNsrfNrVaXV5eh4cNPHzHDhw8gwp8MDDii9Ov7WTXDNhUqaqahvQzmXF
rdZslYXdInQaIkDd2KAqEmKKBFQb55LbqZPDAgts+qkmKKi5xQQP/3dF6JFg
+H98nko1EosYYQIFEu3n8jZFHOR8PeBkwSv/3pGFWqmfNWSj8nBdh2KSqSfQ
xa7qeJPAXZ2hcS3SuhcN/+Q4DrkW+knL6AXTbb3HiFsp6AfNXNN1P/uyjY0F
LQ/hCrmNeScv1APC6FmU8cRs6MY5qaybdZkjpgiT/RB6c15zmROsZwJYMGZy
4klA4xHxffNZeJf1m+UDXIeww4J2YQ5JM6iLw31CuKJyIrhIvV4I5pXylh4Z
jZRePAUMARHjuBXznIMMhNGNUVaw8fQ/jucfDG1N7uajajnUA0Z467ZMv4OK
Obhob8hmAJl8JK0CnDvRcFi9XXGxydedD5BTe3kVb0iidN/ZvNfTJhu4seSI
MkViqrvuWJdM40weaBi97o3nvSWL6B7BYTHoKaWtJsvT5cSe+x8yfJIWbXWI
DgbyQDdI3Rwj/32fRYKpbTflg0JLQ3DrRMJ6IiTpiTvrULH32XKUtSkRoJRa
8sAYtsmxPmMSyFUHpHXw5HecTNLeIfCln4trWP4HnchnaWcsbViyoev112ja
lKLiodqJXoMev8Zy3AZz5eh/Gd68HxQu0F51Qv82cLW/2LiTmcixxhQuKaQ4
qF+OqZ8FMay1ZSxRKWYlE7/PGAaO/sY8awcXJwtWoK29utHrFThMqnkRwvsN
Gy1pCC+jMD7fAR3VMODK0bFMHeT95Z2LotBxLvt1PLCFQspl5iuQmB065Xd5
5mZmfxc5SnkPf2HyRwjkFpVGq5oHgfU32SFFjItTA3ctM57GJqivBNxkAhsv
kUua3KOFz6WauYy9zKCcrmIxHjAxw9VkICU7pUTgzOHsOef5vQm2yHI3ixTl
OOtqwOIk1sEjc7VKoK0Gi/diK21u1jfvyzKbOaXrRgRMr6D71VEMr0o2fYXJ
8AvI9+44dvXAaZKbCpP7AXk1K4+G/ksGb9pGxqFxrloFQaGWjlRFxRJ6zED8
zBLLdZ4ElUdiDl6blUHIjYqUUU9MDHbPZzC9xEo1irLleziRraSspI14qWoI
BGjcFsIxJEQL8i2/Ljt7sV05LdcHKuazvZ1dWqD/+bILXY5njVV+woyLxTIX
6QpkwDX139dQj0lq8X0Q4dankFhBYApcbdTZ5EdX9bBTmKi0y9or+Cp3x8bL
i5m8VwtWVSzRzFBAbg9U70jv3D9plbLkT9dnP3rYXzKjgiUy8chfb0XLgCrU
G1Anzg7f4DSWhP5t2kpxLpnEeabtdk9SmgUtBUW4e7Colc6iJbppxplc3Tj6
P4Qn/xEA8ZLGgamL6QezOFfa6GjeLW4PsY5fMGBL0pNsdFRauxkTBhQgSsXw
D5QBpuJjEtj+CU6KwHMKdoFHYv59JVpOeNNuLnFambHtyG/1H/IDK3TZLM7r
T8Fi3zh2uzXXluCGPVqpdJjBOgDOyng28ySX4qGOX9O7QZBfpr/KOU/ys7yy
vYkJQt6KRutz5Z7PuY7y3NwUDTuB20MHRf2NpPaQ62nCryLSVVQhWIKdunMJ
rgb5aPAYomCgb/DK8Ja1OhXWDq6uLs3hTE3Bf3J5TAJnobY8ViltQWyF3n3d
wXPczXwUfeS+q6lK5uky5lYJcmsYqT1rjPnxtdSqEbzQfo8xGVGy6fAvnCRm
iMXZKMl7K02teU/jvC0HDEvZIJSUD7j4kZ7btJlQAOgHwdyLR4c7wvHXnS4e
5CP0qmm6VooAGGOChN9E8JnhKrNG+BL080hyhsP1JANyGaeAt3fobQeWlmzr
huj0n9ucOZXDVuaVZVTmgHZOUWMRTW2GyZj3/qyfRZLjCGWuIx5r6ElonBEz
+iQVyo6IM2r3UhGTcsWWRlcbWW28tOCXW0+8KInbA8I30rJpLFpCQ9TOo42O
mK9bAkB90HGjsfFhbR76TaGDQs126FnILThKN5qT+LHIb1e9r/a6BaUIpmaj
tIQRN26Fj6IR7hstSlY0vCQswK/O+7irSuxe6O58EK/mUUYmXLJgVKz2jaR6
xRqC2BbptZ90R7d1pRZ2BZ9UsGQUTz3DDZ1gydWSNc4qpOZ1PFHpkje1Q/BW
Mk25hzd9WJyRUWlrMtHKvJlez7c6MULAeMJm4PNter93QSgOfqKXvsGeafY9
1bM74SSkhxFNSmhawqneaP32SXKilrYRK5QNO8Ds2R0Cp3051DFOskM4SL/v
UmJVT6Yn/FjbKTKGg/Yv8sQCf/kTWeV8olVuf3uEMKne0+v8819zmY806P/N
Ro4yx8TwC0irXOXuQqnDDBHhM8AJ2WZkqYkkdlRqV70yRpAC3DPF2u4wABVJ
pdhF3JDCKeYZnH6idLIVvvDozHW6KiHPNHQnyngAnBKRalULec2+afy0KQei
wuNeN4HqJGzz0Egm2HA8NCDfOJjAjw73+1cKmX+rw8NazrtGzHeTxdWWAMWx
lLCjVT6sht1T3tQMzUM160oApVHMf0fydwpwYII4QfEnjgNsrefD+OWxYJk0
G/yp5hQRQm+Pq+mkJRJThzFSu9Jca30DkY5OjW4yooa49iR+TSU3wNeRkwlt
ORVpOb89XsIBhLa2siThSj8JVB5PAgs7ezt8bxwP9q3jPel+25wk/tAag+nv
/fxAVSzf7cRI3zdKLOYplr9YJN/ZD+1jsFWDHgropjNxGx82HxuO94dBIVkF
asD5WEtMsii9yK2nvs5x4qwMKvzivz0pRyonLKknXXX+ct1bNVp4RFyRmS9x
RwIsdNnYPk9VxOKrp6S1ayOQMXZ4V6MiiqnM9KNzsJ19E1W641OsZxhr9CbO
epYKeBUVQ8rdB+selsk6obMhl87sf114FF6cggW4yLRKGyd60XyIlBjby6fg
gzU2WtNE0b1UpoIWXVScCXzIO9NvFs6CWC8ZHyq62L9DuLJrCV7dffkEpyh5
NIMgbOfjTKphO7x32V2goYmZP54ShrsyDxoVjn+74oHqWmgCHfEVELWZ+skP
1qxR4NkNaaPAvPwPn79x7PBK6Sgxlo6QvJ1OmKW4jUT6c4ChLGmO/hCoP4Zx
KWf9miqId3XvJjclUG7Jiwtfvbpe7GpzZPgnQsFljLXBP2WxYq5jQkA68IzP
usYJCRJhWsTBEnYI3WSkxbCXcJIzf97Zu/Q4RehNEyrsPmXllu/8XmiQmuDb
GhpU7/Tzn9Safvn7H7bS7pW5N+BBRWgTtrIjVooHvKG2YjfdPp1zsE32B0QE
6vFVH1W1WE3+GMmRYjmglaDucXVV57OgGfqqu3dWcHpoOPR/r4P5SS7aQzPw
DDPoRZGxo57eg6tjatAREVHSnyO7ufTKRzY1dmUIVTxVhfOOTDOmcwiefpud
UKA9AJo4ui0LkgSc5ZV3pYNUIHYZbHl+/i07B0gsJA9PHxaUk8GRMi/GAjyd
+Wb+vPKmbedb0izcT6z0d3j65fr2xdKnJ6g8hhNudCIFDlAMuUIwXCOzvIB7
N7tuWJ1zzHxxTW+mC/ioJaxn3c1UBHlQ6F8I+QP/tP06jRmHNB24T6Hgl7ZS
OqOpjHWE7KHyd9hH0k1laq2axTxAIPJrQMFIQGJfe6vFAMI/7FUyDeMge09D
lnkuerisGaYxXQW28S5NNWAoVnrwqsAei/OWDkxeIA13fFu5m/9Gu+fFYZJp
3Ej4E0EFXgbwJdvTgiL9reHgdmiZKJjIcdBOUZOANdR3wvR3xqqTi9zVul6j
y9fZyK6BbygPs9pnvAXSb/Cua9LQ3R3cTwzPDLLsm3o1B9gHBftwZINNPqCD
HDM0JL+G+Q1YZ7ADWkviw0j67RdPgyvXhq/3GNHZ2WIU6rryjKsl7tpxODy6
e/QHkkMaSDGjT2pl6AKimKO1DdYjMbQcvylCWnQBHQAzKjl6qJ66eImji9Kw
EegkRcnmtSZUd/QCJkPkzXeJM5k1RttnovAwi7D5WPWv2kSSOiHnEdtR26Ex
7lBhYXW316FDxuGMyRGB8CLxVx1tMVCqeJ8GWwRi7Wte1zNLD84ubl5wunB/
uK8cwP3EuSsnD8cikwf1Z8YLNRJc9/GTnrkoxD/0rSmzQH1fZux0EqoaBgg+
Z6vvoeX6Yd3wtRHSLv59fwh72nKUhGVvCpzrIBMfCjzjK39FtuUNiXZPTU6O
qtoJkW6da1vGtcIgkmlPWW9/nTWvGnjWSfLyvX2PZY1bzvrzibwHopcg73C8
Q0jR/ktakYfLDV5tiRt4NRzZDdTCMcMNGlIkXpdH38CsSz3tc7js0sL5U90u
SsHZwOxDBe+4hI1nQG0CBt1AHv8Zt/ELGijZ5sL3MbvQeKO/E6NYNEPHAS6/
3BSTCDjk1nY2JBDCQhEIKtbTTIndyHoxnnLfyqCmWloL9KfEvhVvAfkeYFaa
0TIMyRDUP3cXWxYHOlMRxbmwgF8S5bbEjHIaxFwXtitgEFvTT7g0qeq8ZLIO
5d/J7Nowirp+kzD9d7plMZ4Xda0Rw2F4rM3c+dxK4Xbj5vhJjxZtpQ7PKuJQ
PulIN3gmtxUHK5i5iq2uaS4oQw8QkiuhdMatfImKQCXNQQV670tnkEbXsEj5
nvF7z5fsaGx5Js9lc7K2bqRzbtYxDNXpgrq0ZtAjoRQ1ABIBVZ4v8OtYQYqm
CfEjeGDRC+DdtQ2q2ApNOyrLm47f70JuT/ITqqpuEBzkrP2DqyF4jd+i4WnB
7Ynjx93Iv6pknFtWiTiLLBBqSX2JmJcIcESndjpw/wvFSo9DEXWMiTcJXUis
DxEVpEYPDIwOKVdOM2gB0eb9oNGK1dbSjRgtEHTYVzmi34huqOnrliYbeiDJ
fZ+OFJil6McJ0TkN8WG5kikEoApmTg+uxgyan2FW8U1XSHVP1HDcFfiV33OP
lyN7zvUzlrklQvmoSsRjZ2QWqMhqaWKK2Sef54INFFZdrDl/zZo0tjCbh2ZW
TAAo8vNJ/vRwgx3HgsXwB/UTnNLD7QE0bhA/8GLDUXfEnqYXnuGSQt5CWRYh
rSWmzqf2TVk2dy2LvKN3MXxNQXuUbxAfyfQ36tV0oJ83K0QeXFDSNEGYmI7Y
q7QV+pug7iiJhz/qQzZWwSGoLdjhXnOJoZHNEu0EP07L2UAYsumsUsxLCcBt
LI+Jy3Ug4lph7jThqTG0AMyNDp76DLTy26Z8dYMoHF8PciaUOCh1k7LSbb97
x5SMP/mfmcM5qrKVVcYy0GXDiQ6NuQ6WxJwgEwLKAp/4VBwmLF6epvvCtgSh
l+PPW3CZ/FgutACdJl5TNBEtDnAR/2dI7IBq9rORmWx22kdFPXbFfec0M3Aa
IrUyIF/VZeGNZbmk0MxQeykY7hZ1ecEH7n4GnIz86CPtj6zQPnGYiuk9Gxnk
ezlciv2o3trensx2piQGRNDiQFncfJdMbCoqsMAsAme9KVykgd5gzuQ8bjtC
mz9n+uYAAtqweSGvB1sMgSqiNVmw64PFiR00kRZxpDgNEj+Qi3drCCKRwS/1
zg85Epczd2ayBN3bI7b+KXCXNu1I/vRbZ/RkwCueEPbOyAmOzj81lmW5DHnP
0LnAM/RG2ZiB/6+yVtQjbtmWK7eMovvme3/BP5UV9sVCh/OyNwbCOY0AttuW
GVbIqEWBCc2FQrFjZDOuHf6BEwDTRRP38MBIGQCESwCCweDzkWsScsl1eqnM
Bbj4DsNouLLHJrvOfD1Ah6Df7H5AVIT+Czj5SVh+LwL4FsAoSlh0Crmn9Du7
THhmGTYGc6h7fNqKf+oCulkK/FNbFQYyxSV6d9MenRisNEjWz+mdOX0Cxx41
UM5jjHltBzWEbRSE9j55TFrDUBg26RuH9D0Ho5w1/neKwfUtfsVIRespDHnm
qNGqzf7eJ7JYCF8We1RuOnggmK39Zm9mPt9DjGGy+duCo0UhggzAKTLKlVBB
7owSkMMnGiK900Vh5avu1G6onUtkT3XEI4GHAXE8KozaKQNZoRUEz1t3A3dZ
DppcjItE8W6WOz7AU3ekC6fyoiSES7Hzsf7FxZZLef85CdWyCBhjg0EGxF6W
PdFH5Xd8srcodoaV4l6xR2a4SrYSAGE9sSERjMkb98nIwOf46OI1sASpowvD
kxlB+NcL4DJiusqSs+Qz2JYdt2boPv9CwmQbtKYynjXCRt+5UkaCuA/K9vzh
rGdNJBHseHUv+gzfhhSpV6frk4yeSGMbRV9H04Oz41HMg7MbCRsAP0dEpwBG
YXjkltxmnZUPxm/uY9xpUf2FXC3OKSJme51WrXNsIHE+vW3I0liTLxWT4o3/
hKO+esPbTzxyu7mlYEGnPACKahC9XMNWJzsgWtLPMe/J4GENS4Ic7eZ+Aw+k
UifPrWg2S7PuackKgQXZsIebWtNbw6p7Re5K8FhjLKu0EbzdV42hRBHiWtOu
eiFGrjuH7nTlbkSlylIUz9ChTi/OBkVB1BZbnsoMbBCnUSfPIvw3T/sKnnBX
aFYF3m/GclQaoVDXdl/cd+j90DBB3ecunRGZvhLAy8iSUHNqVl8h8agjGwAa
CJXmXbgRZejxQOSr+YEM29XXlSFRRm9l8GIhmF18kw+FUsQvmHbs3JwiDeUV
enRvm4EJUusiaVYQ9J9uUKBU6ahWOHRYUFG0DLG5X15S7msG6XjY2ue35faS
iDjOiIEb5tWa2DMe4ELZU7vw9QJzt8EAqKNpoXPNVM5jOHQyT+P+dgtgQM0U
mhGnZc+tSa7iKjk1MMPKNJNRANT0sfFV/mV59HfslFqqSL8QLWtypV2zz7De
bFCY1Oh7r8GtfwAqE+MdezO3kuv94g9Hd/Lo9JmoTXo+jaoQrDDh/RazI6Gg
sd50QW/ipEUD42OUdb82JnVKCARoxSZjKbaSR2bC2UeWy1ZRLs87IrKopxCt
35vs4X+X35vUueaac5BcMkR21+XmPjmdFW0An1NFtyyk9ADov7z3n29pELpW
uIcIaf1TmydOHTydoaJxTcC9c/OTETrUG2+vIfQ/VP1v3AKI5nFihJ5lYw9P
ixOvrtYIdmOsplRGQhx1+a++WZi4Z0/ovdkhqRFs+77fbS2GQMlHeaSV+Ygx
rWdPaUPaPZXAWLFjCCtjD5/5X5BS7Kj789uOhJdxIRw1lYFy+1kQfzfdX6Dp
ymQD5BEdMeUXTImT7ODmstf7PIxO9pRUybfEAlizQbMojniu438fEJHJPuMO
8xeQcJwcZRVKKsu3sHxTESJEacNlRlZZr5soKl7cxcDvYTgBmqeFz10QMfXm
8Uv3DWr2WNt99N1KOBt9X4XsAGL1feWfTXndgbqJ0AqutMSvlg/z0apYEKkn
3R8uGxqMwivBXQEZzloRNczfEEaJuvTqkOxolpekI+uW+RAqy3qxDYt2JP0S
3BWyI2ehBwBMqUaewMIn41Xt+AT8dCcGuBQvosvHK1qGCzZ7edz6gZcZ7bpi
ZLKRrX8rfRvLCMsfLxJdfsxAwPAKEpf4X7YOnfkCaJ813STkPNkPCfdDMFhd
quazN6cbRp48vKCbnbxJGYsui/hSFSEYxIUGbybtr69mfsuc9SEwW+uLtAVK
0CBRwWkZ3D59FWGYOdkLs49KGNdP+O9t/0fp4PnauDigtex9durSWdkcXm7H
hSN1SwmEnpA3nuGxchQXNdWwTWWolKjKkpPeHd03wmg7cq/u4wrjy/wg2CEe
6bBrw64zrTLth+o5yV1TkUavic9aj+kJnTMiJYTBwee2uo1bzvjy8oCzU62N
CeAv/Sg7BPBIk3/ZTQgV2g5epVjnh5GDr1wB44uVtxiPzmZbNa0Uwv+JmM0F
pA73H6GwZbNkhjZ3IjXYSzNJ42EIWmp/NrJPJW8LV64hckAfabHFA1t+Y7VY
cfV8vvOTfPM6+aKij3F+KB62MN1pqfGl+8dRKmIgX6xW6QSUSHT2x+GlcAXc
T73JrOI2BO95TrO8Qzqu3UAZH2YuLv68+QSHI0Pmph7Lb/15fBWqi5FRvz5m
kvGOORH3I7mfz0D+yVby9GO2o6su0VYqhJs50+sdK63QjWBdoTrsr6hBq1b5
dM1JNFWHhEu6NnytQ7QliqpHP3H+xDqbZ/+6ANr/GereIEj1276zIl9IWh+D
UsKa0deiv1WfmoAIiu6gemH5m69/6VOSLLSTzjlv/nPkM5byrGtzPMZahr+k
I+lrfYoW8uj1+tN76RBjQD+4mNkZqZvHWUcyyXPX5FsdaYjaTiDC4a3uH0TX
P+6psddoD0RVH9nFOJC0ZVMb+qB/5ajGMnR0ECmnwP9ic8kV2bNi7eaj+g1A
0wXIzKfGcrT39gANUFhn2wKq/v6ORG22XfxZnHNZvNbHbN4Bws3R64q9SfPD
54sQ7l2qle6oJJj2cPPJwyb0YIlbscBjdONcjogn/gvsUBFwqX1QEvFW/GBg
Q2zC9tzdDfHf5GsHbrGCeVZzg2Dhe4PxbB0ashxSyE9iURJfSFyu9L3CA7c8
axil+ZyeAo/xukGkNBBJbnGNrW8aMK6Wj/5y79dHLK3TlDCnkfnmVblYbl+z
Zeu0tShJ4xhS3bcfYl95ixNozANANiXh/J6gIDwX5Zw04C6kVQOU1gIiK2WK
r0fd3lz64nwhieU3SlpwSUh2/apEvEMIpbh6+ERLSgAgfl9+djRQQpd4LZ/o
jbLPa+xAyuIsxPnK7dQSKjALIWnPLEYqpC8ZWfjK2OoBad4Zs/KM7/Mx3SYh
ZiFs8EXCN1HJ53DsihD7qMHbMHUiGf4Xd9zqjqC4DL5QedXSOxdF4HJUVEDV
buIoMnpk03eQmJL46rVTChwMEJNjo+gi35JQCEguH3fNZVJVuLS9fEW3siwJ
Rxoc6jXmQcPo5lg9nf6WQzHcglYiOvhtymYgZdlgpuMvLnfVW3jUncokR/ir
QcUEQNvn1MTbgEafLORDOqEzCGiHS6QhlVRb1hxGcx6kecoQmvvV8ppeTaby
zf6UlRf4rsp8Aqm7mGV3ML3zjvs0Y5GKwyCMWItnLmi70iMbW6i7Yhe6Q4Pg
dY6wwb65+lCMEXgT9piC4KUZDSxdUDO7kaNdabMXH7lBl7OTY0RpwNtBvAVL
2BbG4nHRh7/NZ/ba1tEGJhfVdBYKZ8S8G2Fp5EvaDRNRhY0YBRQ/e6nNUu7j
zCgQsEQ9jNEthrry4mQNeET4t6AJ1dz7x4H4KDrmc7KcDV8zMhFqnP7hEzBX
9ICKV/GdcYjmu1gIaGuVgL4+woAWkk8XChhDkXBEjEbQmkENSPNX/0kCtw5a
Xau2tEW5e7uXTTs5YDMMsh5/IQmYLai5Zbu0Kv2FJy5g2yGYm6m+QB5eRZlT
cNAthFcbDqsY6J5nU2JC4gxDPWuOk387r6wLMH9zdMO7CBkxrV22/vBO+Eiw
cli157sGvVEDFAG4mMSVx0tN0JP1cVAjtoA8mOD+Jk1qcIve0W3lqBo0Ru3K
8YAElCqHWhHBw8dJzJIfewhwaqlTXAp59csvI4QG4vF1p0aFI/cJuJbIogDJ
GUg4e+3Tp/SqYMqEQP3C/FyMXaQZEwxYAF9X7yBt4ktLoz0GfAbIkRghTdKW
Jz6HRdofVG12JL0aFuxTQbvbTSPCTiS4QQGZlMGuYPhHzi+7umH/XqwBwnVC
Io8Dgn5rZlG2Nc5f7/PXsXg1aOrIfv2iFnlpURzA1XwVR/KH8SFdzttuykED
5G6jvXa1PtDwaGJcrW4mcNFGkM4R27xI2j40XBbnzwa89C5NzvVpFcERgsRJ
krdQIBgBKOEGGG1ZQYX+Ic9W7dVyuSuCWLLz/JrDtE+7XvRqAFNc4LmFcBMe
QBeZxSM1RLZ/ogpHZSc0FB/CpTe829O1GwW8tuOFFKqUoNeLQWrJrK6bVR1A
IfdN9UTiP8iPSv9lPslyuYUMSvP8O1BAVojHC04TmTj4JPMlStLvxKd7O6JM
r+C7l+QpURXDL4WS8h8ne7pNfHWo0EjJalZlGQ2nb5PSTpkR5Rp3l0nIrIpa
jqApLQpOkCBxFsMQmXjBegmbtM4qvI46fZnyK99LRQo6fS/6xVKlP29fJgLi
hv4V2EDnbNUQRLTbQ6EgB1xtc0rb205FwrmdFACf33YKX+Q+flpGND5ibhs+
ylEXmeION+avVo1Wv99Ur2Y1DRclEkAD+ACSXbfSvveMLJDNF0nXX45lhhMt
MeTWQDILU1F1/LWHZmy2zjRBLmw1K1p1PSrKW2TSjJeCazukvXTEdRa31CHW
t4DGlCMscNx6P1+Mvugss08Z8MmZYYoFn3Kf7AudQ22YkyiSrZtqaaRaDU/y
2LTRILTJKEF5et9UFYXB9+zmheo/Hr22aXytF2xPiwpqj868L6vH83etrYgG
1qrTEpA7ePuqa6Uj69H7pjMjEH+MTkQ/gZJ8jOsSeoU5ev22j6ISkXV4vT85
Bo0plOVW+6WlWlwvat0QWgIzNgP82l02IezsJAX0frmniEWZfrYsn133eRZ0
XNhwS6Hka7c3f3XmXWdppbkHWiO2aYNGQcS2ezyn1f5MYcA4Yr9fCUioeGbI
Rs98d49CWoCp0q3YOxpFngGDsD+9nkYk9arF0TsG1afzuFXwjuEZnotAsijw
PEIBpz+JM2ytFOilSKfc8fl7V8Tt4WSNoJ2pMd7fT4mzhprnewG1jnjUGlns
2PKPtRlDC8NME0WVYXa+ElhDfAVOrKxxyCjNawHhNgBQy1Dqhah+LAsYhhs9
HhK98346mHPQGW2FHEKyGqcetLCXiE6Q2Y14ku2uE++rnQo8JFUcC4wPibFG
GxqM43aoDxPp4XIVZ4UJa7iWbzypzTexWdZwoMU2RBeYuF6yqdMe8rT9q7PJ
uOE5QkRPycGztTrGpdCQauYFUet4wm/RCwQuCzGQtHYtUqmoktqnyiV216Vo
ErMci+0ovEdFyxDso2jZHiMLEO7nytAaSdRiivtLoJaYc8WpJ2Cy+CRFxEWu
mIWKBingc0ymcrcymA++9We8VVh8DQqQTh51NF8Uz1ArxbA9S9WR1Y+eBxUO
th1B2cfeVjjU4jRVj7JpycuPBqXFXyaxV/0zVY/88+8yw/hur86YyZ6XI+YQ
XvUEgd3Qar7DDpGD3M4iyKbXFY8TseZzlCvBF3KwSJXDgS5IIajrcSq1jdvu
kvXiqNWNHevnNFJdE5c6/97/w/aFMTl9w3QVW92J4sSLD7A59yw64DuoocqN
d6uKK9A8RuaqqmD5DRyGibKCYXESpSE85+XlTYk7kaj6+viZl5RKMROMZj7T
5JLG/v4Fnv/YvaI+DtLheZcls24y+mZzHFIztIqAQGzuK9Y1gBCQ0sFeJxmH
MgtVlcKdlt0SBdGhyx/YdHh8y0+C9Sx8e9m3IF9JnnKBabNJRXpOUwR366Vy
17Z9o4+4ZgPQRlWgwxuULITkboYUzeM4/ycSx/iSPbMcjOsbBbmt0XNWXtMu
02l0OlfqhoGoYx4gEGSWZ3VfnZtPwWSR9xhNPWgGx3gajTjaEt5ffuV3RtDI
6jkIb29qKZVJH1zvgGfOwZl+XbtGIWwRVq/Gt+nspFmltGBkCG75MJZyKJmV
QO2FotJowOhrEOKHlgjE9BNMkhnt/UeiWhifcPzDrN3/PvjLdWzwKlEWdawE
UYFaeyWVEFMQJqdddcUfA+uzvJkYpz4iQQaPO/QzkxLEEkzR5PzQ6GH+KToj
FHAW1dN+LIeV2c7iGGgHgpWjYL8kXCY5YTjUeDtUeob6HPDMwVhAqYZWp0H/
rn/+A2rsPmpgsU5WFh2bVl5U87KBIToAEZ+DJy8nz70mylVgDN8FqsvbA6IO
CvGHX047EmK2jGGBEHzDnUCcJO6mv98a/Ff0HSiBae2QRXBldc/qIpgt/bMB
CLQoDfCYtP71PROWZTSC7n5pMBsKW67XJB5zru7l92h3a/vG0xua6Yh+RcO4
7k9eHLDlsHfSkyu+tumamU9umzshRln6LVIty3BzL6ysxbJZN+ZIudoH8110
/UZgAWIN1i6awj/n2wCrodVEq27C5QRtvE5pJsga/vzPhIVVrFda/xCplqRh
LX/4srTZpHs53XOanMANzNz7QLT6brZ/DSZEnSSs8Gs3V2B4tEADticaUPUG
8UYuR8ZaFuJOZN5DYheZcfHQ8xI9x6DNsu6HPVOG6Dxe6vP4IaooLFoq7rPx
zzhraLwa6CeMEXpVIryqpqZLeoBUOcRaHsEFZQpJqqEnnn4mUgejGrEixayJ
LMnB6Z8gh0sdKhiLU+RkmVgsDDoqWhdRmjJR/yXSFqFetrNZVrtSPolf6zz2
rao+elavcSZWDm1rLoqkd7A4Re7p11ThZmaRFGVR5zjFwQuE9MCe0HMEZ86b
FGRESOBMq/x3Ih4rB5jlN4HxrfyR4V343Q5l3Qp+kAz/XnX3yFAe9HPlfC5J
dQs3ZS5hJrAfWbuVPYG2PyWCpuhJTy40MMBnL4R6vhqoaUUPnRg7j/X/c1be
5NVycDOXktytyJWvF9IijZaHQGN6l0OMtiQIT8UyT7LmelPhePhI5W1S5uNe
Is19SRFY9ySPBWMMiEES3XuqU4SbYYDqgt7tGP0Q8PfpayYHmGcPKnRP+wHt
yrVnAUVUNWB7CWpYf0IOS6GGU9OLATCxY//FFhHOA6VTWYNgmgbtbvw250A3
Y4L0ke6sgtoF7TKwtNm6Wllm0hqQJ8Wj8WmOFAG/M3oZfS5wuZv3m+I7CFpP
fCkBXLvPkJK44hzmjpirztjCAlrLzsbkp5eZAgCMcQbYUDFPcMzXUz8zbWZZ
zcGhhkEDc2mtaUfNr3Khhgq/CwHAlV26Ze3+8uOEFOE272lUanKpkIo5UOkb
895bxFL0e1EJ1rsPNTWDnUt07D4nh+rxjRFROBmei+Zn/Jyyo5zEan2w9YUH
Ha16Ssy5HKLLtkGuo98KqagIcB4ynHq5aW8vRNIXr2Ugs7Lp+agEk8o+pFGR
Q/IJ0F2UqEkDS5Xo7XaruxzKB4MqpXtC2qCh0NQBwPS8xcewSFsdvIlLFUps
prGaV503dsh1vvtKargW887hLLmUtPgNJTPReo0IQhJo8c0tkE2nmQKtYr1D
/MmB8n7rYVP6u/M1vnztROnMs9VoDJy/A8Xytrwco+2rtA7PcRbIbU7m9qbr
l8/FH0J2QMEqCtpwA/crQYX1sCQhpzZGvaUa/n/HsJGUJOCSNyNq3QclC6NX
qKQgvGrUWREnpkd7YOPS3eOe6dKqVWTTyg/9Cve/diLiXgf6097UPV3xcC1G
3HiWInhL4Iwm+LDMRPRsowJG91wybLPMs5/Dl4Hj7cyFcdF+0coePB+L+SH1
DGU7N/+yd6omthTmIVNU2PcsQcNq1E/R+VCAVzIUonDX9zhwVHaLiKen8m+T
MguaxjrrF2WOL1w9Nha5v21faBWCX6wm4eLCeUI7SDNkFH4UDN46MeKGXvew
9Du9HsUqLbpPASwP4ba+1q05EPXgFOoyWRTMn4k1uaR5WIXT/VZ8en8CsLH8
fqzyVz1RLt9uCGcVIqapjMc5+SQLANJHg4FMAoJMHo5GkyMjbJqbQTXHzOuK
8a+iEzGvWcSSbzbLs0fYjDsVZTRiL9avdP4BKSt2IE4dyqpABWzU8mzXQowy
R8KJ3/ODL0XSqNgANBNfr2UvoRTeAQppY8/fNxaehj/RMDR77ug4Mf7H7hPu
bMUmcGxdplXEsQeaaRCRADxthxu+R7n7khj07Ll4pLbfqKepfObMZNO4JCal
KsIIyFNEC8q1Gj13JAEhD6mqtazP8dCrZBiR8uxQVxjtTmDbakQ8XO2rb6Al
q1ctdwpVRuPKE3IaG93vhUetfufv7RElaZIh2eObJX4ZCSLz92ceNB0hR+5b
e+qwGlVbw1njm9BWnMHoGCw9/6OUYNU/mCGYjNNydklhI+DLRpjaIcSPnL67
h7C59Ea0KyyUID+z31UtLtZAqOWiWrvHkLgwbzrXrBeiYYL96sKCQnKa/S8m
i7iDvw1qE2DgIpQ5lGm/eeT1F6SpxSTuXT1wkhIhdj4KetoZ4giB35s2F7Wf
S0RkCzdpMbHQupNKvMMNIPpX7VcpYW+nMTy22UVNGzArlOXaulICsfEsDrbb
Uixldemk0/mzmXmqElkyYm1D6jJBG13H9Z7ZSApmEBh6FFeCrOBIujJNETPU
vNSQNyDlcSXvSnpACP3s1ddbk1fMRTHIzqAVMbpKWnKfw/oYOrtbljxjeODx
aAzq0b3Loy7Tfyn9TE5jfOfV6kIVxlx8TXJP29OKVS2MOs8cXCtlKpBQXHP0
iBXJPygGFiOG8L67n2sUOb32YLXwzKGSElvWjOdSN28yc52rUOPITWjaU25z
KLRpc/TJDhTb9FInqjNbdF6oI7NhssiOQgh9Ff8LyrxkfA9aQAaKESKyA6HM
DZHpd5OJFHs0YZK2sxgUAuIXIi8DKp0QamAQh1RjEVYO8haoHjBSDfXdZZWY
KLgmctCdEhqTXuSEw+fJY/2SlWb4ApphwTNB0ibc3WqwmSmfP/F4ny1ZnH17
mlATuI0/ARJnADOqEgVYAD8QGUGYcZLit3bY9BPTVH6tzFA6bXuFVBuB3Edf
j9lNTLMKKJkgfbinRi4rqec2mbST1Fi700lcKUBUSmn97KAY3GokCTEoi5qs
47DKoDOtkjfCySuz3ZavXFbXk4jHg/4NiBeUgfuq3IPFR2y9q1PO7UlMFXk7
hHUbVT7A3chFx5CRRuImTgaE6JwXhqO1g/VdAeXzeNaWnZGzPsnwJbObQ4oh
G4KOjDpHqnMHtPmfn7mv/O0R+RsKAeFjb8UzHpUxoysKfugfxcpFTOxWKN++
HYMuzCER0nYOK0TUKmcEi8qLLi+nIcnouP8BDUAjr6sxk/OEadcQm6YtEi85
UI0vLIrKqWlbMf2diS/WEe6gsc5Qzxli7Rp6W3LX+6HFIMpijRi39Z569VMu
kRhR9NwWgAzSEjh9i2Fe9lavYfnYd5aoONHBdgJzp6NVRXNbfqdA7WPkd3SK
NvlB4cP+P1ei3u+Ht0+qv7BX8h3IISoNQlB2y7g348qyIroe4/6Mc3/tICEi
hCQV8fBTY5NdJXQXlsXkPeacrcZYAJkMgHK5USA2wde4nxNgpFdS7HvRTMIZ
hwd12efCeEe0oG7Rf6gpcQs9t2n4TM3zPtUdZeYLLnSKB4U/4NoeIG7+4o/y
6F4EJcCgnMvZ/rcyoVbjWQl6nqpR+jsHe+4GZLK6VQzWimXuC83dqblh0doh
DQwtZBjNl4kH1nUhGbZ+sjWt1Dt52VU9n8SqQLw63/IpvoIDHyupll9tqe00
mGCyQWgPIUdyBaSfaV34D2pmWcr9j06ZJLE56dUxeXsAK3xmMjG/ZtYHH779
xKG9DxoN9P29nck78l2HTquET0V95dg0tl4A2Kli6VkgBj4cJDtiX/UEpImf
EKoM+YtEq4uS+S4zXDEDmV39//H9zw5vd4cilLEH4AbaRVcd6xh6VsPHJtk8
JqhpD5ld7+XvX9cKM39Aq61RH8ymCBBV7eVDCIpwzJq+vZz+Nsvjqy+P1YRw
QrrvZoI3BM12eTz4+pk39spmQ7PfWQl4TgToJ64j4AkKbvqXGIL4iFWcg/q3
6DHDYnnUFC3eE+wYuim0VgEXXz8dwM+Y2JpbbVniH8nM3KHRpD6gwFxszEQP
BXZQeOZuz9SoY6cQ0P6FxZoNQTeXb7ifqhAzDJ7fTScijloWAoo51u0j/MBj
W2lGNlpOwIm8HHmKhFCFSp5U902Jm9uFnvjQiP7UKH7UsYl6hyOoT7FVK1fp
xTf7a5hp0YO7mclldUtsi+1xRIfvlNiPWXjcMvyYiT+/WeeDNhJ6mYa/rxhI
YkdL6VqRT+pp3mXytkbki3Z+8t98B2AHp/Kq5FNtgUNJF2yVNOrG8n0mPf2y
FhYLbXq3lpH181+avDLITLu/afgGY4xZN3YTuDXEBpSTxZrHMHFN+AZuMHmy
yN43ENIrZ+rSHId6i87WnMaJ44CQwV0QdKIa/1Bnc37afwoigyWBWIWOpY2r
n9LkTTAi0R9e/65CyEqqo2fsqfkE1EYVAnXnJwaayJE34H/BpBQenr4mssrE
72EcOq5k2F671G8UTYpye/L4lCdy/09TqvXZCbhzuVeNWhkXFQ3z0p+HFRJg
j0W3savBOL9q4u8+PctftT5Nms9djNw6qC9rth1YA5zxHX/o2ii5rZMt/Yl+
dHXTkYts6lC3QW4TJXNlPTu8tayH0QRhoWABctynMrQ9TbImu4PM6NXZWb6y
uWayVj5+N1X6HpVQtBjDQ3UcGDuwVemU0ZLoBnBEJX9JQWqH4Hip1MEdo7ki
aK3cTDp3sguWZqErPNI/nK7HahLArQDkbjF5nDVPv2m8I3RxIntaAFxUSd0b
Ve3qbbUhhK+B7VHsyzUmDoKHKJEjISjDd5P5LkSzl0atqECzDkzyWD5p+2iJ
4dWCVqLsh8hAyPlQNK0So+6GawIbTzEpEV2xNllR8fg5OynJJ9r5bVAdarfl
950gsaKNKjyE9RIxaDOOCxOKDLO939pJu05MWx27z26IDXOv9HikckdVNYZD
DQaR8CALV9xIEcncTKIhgQ9Lj94XUGgX3Ca6uO8f6CkuzfrMDO5o451MYrcY
xheV9BYceJEsybQ+dVQLoFeDoRWrWl0wyy+fBmKEiWEWZycN/sIZQBs3OaD2
5cvXR+DmfXv8IwK0IBgA4QGNnjFERbWD58dINnHqIqMpFcicccP8NhnbD8aI
xa+fRX/HE2r63I1YfStcw94LWwgep/E0TYwjn2r1UgTYleP3wef1j+P45KbG
gQg8fjSMBYn8a4UFnYwtDXWzvX6CLR2nguAaiK/eA5wF4fhUtyPubO8vGZQT
giP5dWHeW9bHzYfUqaqm+zclS/QJBMMxgIUi3KXrZe/a5sIlPM74wwlm+wy7
zadOfEHzC/aBIlWE19cvhRvwlPnaSa/yizfUNESJkWGrc1S92RRzzZa/MA93
MoarMUN+/q09yStg4zc44B65PZ169vervXwww8HCkLrm288kgDka2bTOGbeI
g0vcYwfA/cyzbZG5d1F1lvg9zB0MZBV8tjYUCpPyAdeVCICFQITbpGkZklxo
PnY8IRhdrr0MoVEvFSeyM6RH0ZoH16XMbNQ3hjdah3QM+VD5zGnQ80LAMa8N
y1kdkLc5fngoO8btPC7ZTLPysaik9AQOXWq08tQ613OPZm3PH9yFTbkj/SnD
yeKOCrDJ1lWmkV0nKFiEbAZ+IJg55ueS9jK/nKkwT0VSUVdv0n3mkQ/xpPlS
0314xIT/6PpbmbB+qZmmpoWhbsEU/KN+uyk/Yg30akL+luQ16+xoRLf8rQtw
M7ChrCtVy1nJEsh0FSQp2fkh0mzKcvfxRrbxOwmnirFZcVo2yW5RqeckCDMN
W0IbVOFSw4DOScRkuNmWFk+0LeQYsTFp9lNsFKnPp5FZu7iuFmAGE9SZdrWT
59LyB0bdBIbpEmC33jkU6nX4iQLxkPjsz9ge6w2HPey4I/Ipj8r87z6VD+0r
iyXdqHbSZE4tms0kkBjjp0hjuIPYR7eNw3631S/GWndSO/LzpnzI9xw6woS3
aTtUqNE0pP7s4s1mnh+2dTTiis4TwzBZ/S41rKpEJKRSnZmhkIESg5C5UBlc
xza2yWPGy4YbcSpu/RBkRae6YOaf3bOfqCVJp3QgjByOr58QJXvS7zQCzKAz
KO0d0Z78OrSYF0hOcdguKjte1QMLSOnB3MRlOnKBr3nIS/Hh4DGDlMlvfxYL
NQfAItdnO+HQxnTeJ+9idjirOuTrDFWIhbUrpspaRsTKhh9nh4RldR2wGnYF
rprmI1L5jAPXMdaQ2rpug1ZqZqN1q97oS6Kvi/5Y5TEsqh0Z+VOKvwWHD0g4
53czrJDQ17Td0g82VVdLth2LD3Sglbvm4tziWwdo4fy8hOCgCwNTt+MEWA4r
AzRREoeUYjSuD+IOLpSrxxkf/C7zdjFqmZbi1p5DMrr1lL/p01rujsvrBr/1
485KgW4zwNgaPFT8lc/jT+Y2NlkP/wE3YQYl2QoHukhfVRL/P10yTAZAQ/gq
SQH4zKR+/NEmTN4RPROwXrdmMhpEnA0lp5tixB2HNavGbqdHVYvECizTI+lX
cyGTc/xlnH6i0N+CovI/RXErC6E4yntGACKAIhokCuX8EPweeZUE5/GPx0Dw
WtijILxPtlwl59yVXji/vxQAAB+PPMgW9TcaC7RUrxOHSTaWKPRZkq8g67mF
Qvk5q5IHkaA0y5H0FU1TWmX6/avEWtQqHvHh6HMH78kBL2osQCrl3KAMpt9f
Wnxxw9A+h+m4Nmim/guuu5PytpO4+3+ebUafJ5PZVpp/3NeiQtrEusAAFt+3
NgBzzGOcyMCsd7f9mthcUL4213qtCoV8yNNpXBH5f+AzuePMXFX4fDEvcYl5
uYuRtEn9fmnxP/uZtB9hhPfs40J7aZhjJ+v8KqJ7LCtXfEQYRn5qk7o/X354
mFH7btJ9nFeb0Ac90569vQ9KOwtc7x6UyrdhTrkWp5G/jLds7DQOnh24rLgr
qm1Qje3WglbMQA4o+6FgSA+JUKeHImU6yHrqXZHSe7tVBU+91gwFUB283rMo
RldUGEXlTzmavAt9bLxGf0+vELWbsPsavt9Fo9/Dh1KozLtG4rKu29hV6Cdo
Dl9U+EEOCAGTNQJw47Zgx6wXsEo0aa8Xceq9ysPWeih2q+2VmEqLHXEKSZmD
Yhz1yf4yqUhMPIBc4B1tBYO+co/RBdNWZVkZqGvwJ0kmPqN928sqbDWaeSk7
/+gOU1DMOnTxH7DHr2WG4hcC8fXz7GW29NLddX/4KUqoiPV7T8CWfbbcMaJh
W1yfJWxsI8pGjUTsupcDAgAb1K5wOXCoHy5zHtWutsYgrHdSwTSDVOfLSG7T
WA6yNYAE33oKcKCvQ1UXqijNEBHRJgrfI8T0wiWD1wJHvs8htYRUhSRPlZoh
TRxFgCOBBXyGpyTBs/dZqlcveKNKX+z2LTN6gWdvRzI9hXKul6p5njc/ACV0
6o43BbL+7Cl63E6B/z3h5fIluTRNmPmwyj+mYpDM4WlrbedqvZbQdrbEBOgD
0YYwqEEEVgK7PljONf748wur0sepoRYNgDgO0UrCJgoV6npAvbirwT7xIp3x
GKuv4Pil9RMOoP2bJcL5AByXea4xMw/kz+jInv6nFyvqnezcj/6Lg+Ds7dGt
JQPwltfCsge3QM8p03WZ2O5c0lpww7HgrzuONQicxVEye3Mbvj7Bndd7LCGz
l7LlUoJ4LAmv0/3rjsVTbGeoV8WIj4bR9MO8RLC2OzJUkr0O4FEcEotyTIKL
7PWKpgzV86FOecBVCaUjyj2O+F2MQQlz6pFxdbM17NR57Z3VCCY+GhGxuA9P
FJyGC/IUwfmxvO3irLDLThMF+7fr9GPj7/I8zwOwJ1Rthuzp9cELbso/BENE
RK8ZDRjcWMtEANVcPLNWsCAEfPPpIRxh7AdKvsymzsQfG3cZHFqHVRdiJOEJ
cAxFIR04eagNbEgXv2fYKKGXo0auVw/283Ed2wcDJETV0HMQ84nr8i88i+K9
d/kWSjKg7YvSHBlXULK7GC9e94orB9sJUMzhelnTiDCexvk5pw7inzTnNxjM
FJ53Q5kFuSkCWpPUb5YTxYapflm+WwGDCLqWnDE1XvJfhVofv1gyQAkiQj/q
QL1d+NACh3TP2CTS2OnoiWwSDwUsyZhX98VCnb8tePM1hzK19MNvwOQCJuHs
eZZtepXap6NGYESk2woarRX1Rl3fxtWfXGa/HojCcp3fQEF38FBOBSiCLt/P
FIEQmSlWtB32BmIKTRXmOjfOT6CWxXUyhjXi8NMHb7E2uKewNUbhRefQWVyX
RY2Tzqmc2Cs8hwEe1OBx5qzyYWtfbUe5A6gOSSUXCd0BNGih8m49sr2P3M0x
i11mglZ6UkFYGiCYEAe284rE8eMSPPpuyEA2xguURU1Ig40wP/TTTExgSv7f
BFKkNqH6XZGXqtO7RjxvwQEifO9svaeF43Fjtu0lEATheU/V4OgpFdc3gGsi
kdS6gmOtdykzG34y6JHQUseYRSO7dzEw35MzcTYpeKo9veNsHspb+Q82f2m6
7GUCa+PedUhH5/0vGFYqvK5qwOEZgNx4TJywEblSBP/T/s7nVq8VhzhlHXsW
HIjI+sHnr6cq1NV6v2r33UJhjm5JqdWKNKNUh2gBFiZe7VrrD3dmTYy0CAul
pKygyjf+Ov3u+Lu4zzWwXTMsVLK0dsQb+vc6xWpmPUqxZx9CuPuW1eXTB6XU
XXOM1AzPg2uGXd7UXuAXvSVyQDqEhDR1Sxk7P5B9KEDJb+V1K83Vst+1ME2l
fGa4aRKLiKRRTRN7f3866qna12MsaV2skoftz9LfuJJ2sQFMJWsa4ZvOtcLa
BRVyD4jCcwi9M2e7OtYbyHmsIGwxSuvTgkMOMtW4aUoTCgKaRRCjHT0zYQ1V
SgPmEpqyP+idnE9qDaBFDu0URxT8g7OIbdUM94BOADO/i8/feNV8hd+LdkAQ
M+oD6KDvVYPqxWwuLTilKSeryNJKOcPbCpy/FXGiWK2RSMl1iLLbwY80hXaP
tAR62tQKLMwcndBmHRkVXOv/yDCzQEsxoI8DeviV3aVQrYJjUXGhhrGo5AfH
EWOy/JPCtqhzn1GrUrAlXevYf8Iua1AJgpW+o7aFkE5HyZbVICncVeOhwjGR
2XgeAb68C/WQDlTH0wFs/cU+8fLpcFJis1Wq+JaNDg1gZON/fE4U5sb7bQvj
1ZT4yDWkj3xq+OsvMDRUdywcEnwsHPp6iV3Px6GRj/dIAiuZyTqOwuvubrCC
cVzVxbL8ehVr86WVh2nGjZ1+K/3fMEyTaAk4EJTo2wKWHF25ALPEaYhSLQV3
AYHGSS16lX0+350myQwClWYjc8uWc3ljiCpEqJaxCIs2+19AZFCuLwztzOzX
B1YCe4tlCt4U21LqDVPAx47BzCWAtuso4xlXk+gdarLzRdFn8BuCEC/OYWv7
Ck6dB9FckxECJx8x8xhUuO2ZezkQWRsJOysVQbccxMglL6TnRR8rJocDjqRR
apvHMbuc+ezW0MXf1NL/MAAmdy4JrFjqVk8miBUsgb15wsakCdzAkmnXR60m
RHjQCB0tnH2y5OG6J6Fa5s6ZBbIIdjyPjw0pUfC+EqCa9rvFdnjAOc4Dmbfr
Gz6vEjzPt52ThGuc2mTDRnHsjLT+oAAS1TjPeXSrXAdhucbjRuBGPNy6fZTf
ByO6ia9eZGlxe6Dbq/pGkZ1R2PoY+p1lkkcy4epMYYaQ8+0rB4ZlzfCVQ9V8
0XMVFYG0XokLOIqSBx23munCwsUtY/qEVKihVx/5p3mOnG/DO0lAHI/wnbHN
HmGfzV9zCjwHob1gfxiUneQKLZVK+dEjW+gn5JfnRFMObUthcx7GD7T+hpPY
GKOtHVh57y4CJMuiuz5L70Jr128Ut7gvqyKugu+LRDg2Wd4sPdWjG3mGBqSt
oi7bInpvDyBM/ojS00NwhNG5wArog9I7Lyrzb7dHOydakM1LnbKDERnEa6Ga
+b/3D43BekLN6hgRzoZwklEZ/rKOMPgOXz9uFFHZwLboyj4RBc1dzBP//K96
QVczZrIchU+zcSgqnck8SJu6wVA5JX9yw+4ZwundyZ68mjNnN97FhHLyDtQe
Z+cNu1Y1En//JgLaPVJI/p7sYJ80PNpyJexLvvUOFrXVLXs1MdWnpg0tLsjr
spYJTylK8ukh1a70A341tYIy5p7Rn5zpzfFxw7n5AgVCPUzfNjPKaTbAuFX5
vRID8YJ+GquXj5PyTp78+TaxQjAjDyl6pwPpP45gyc9icQw3T8J8T0wpV7T8
EC0inpiTTbXpJoL01PP92Ix6SO2PU19dcHb34cOl07HnKH2T0ifwXrW1++br
uGyGc58bwPp3x0Ux/tbXJSzInwIK0aGhjWzs8/GkopfB3CNp4oc2X2MmjRxj
P5j2mB0O80tHWOd0c3lhkyErsBU0wIBetNNs65zm9VOGbLSBCbPTpVtrtxE3
UOVK3b2UtBn1nRF383sw3TP21cRfBgYFTdAu+ikijpBPa0w9mlWR3zz01pK0
8JSPUvxiYyUNPSI2wdJCKJsILP9qiSV/0d7XPsLNneQrf3alcsFtc9qQx3v4
oaLtV8VehgdP4QqCGGktipJE9JInCI22hw92mL1r+GkZCW4+io2zmx8uyyVt
YmxJaYNSO3Re2qfG/0kfoZiM4J9VrgcZqEXINWQlXJGx+rYAuGWDPf3XV4gS
qmUE4e/Q4y52DSC30vAVj6orVEt1BgOSzl8uFDi1cU1BEZ3y/buqmHMAbr2P
TWfj+nf0uQPg9PE/QRVymmJEbzlVbeJ4+07Itz80jids0AKD5whOFbDGf21E
v6lTqOG/0oiMpvNDt7KCtQ3GwrPOKdXqvP1H6nLim0bngluRLx3wc+9ZHikb
7f8OpPFkp2a9wkeZdtShxRj8BAyUTRTsfiozbzvXq5Utof4WvkpMUpHcbWb7
ah/1GIp7I/1jCBli9uFzk4YBkvrH6TYxfvKvoDmdggiqmmMBbXTKQQrKzTs/
m4r2YQLvTioghaIhcVCm0FCPi0C5nkGSP0No295SGdheETzcsl5ynruv3o28
DCGmPQVthZDlp9evmWpZrXBKxDiXwyDlL4Dccxz9mu2cIq6qlieYlqU08+xw
NXHmDL0AAQzV57sMRVFwXMKO4FNOv3sonJBiEgpQFJvkPR9kTN3/HpkZTJIH
lNMLJipnEll9Ru6VAO8BEfZwK420Q3RPBKogMXDbWp/vV1a2WFqnyw7mAwV9
IVN6tlJvzQMsH6ydATxn1wCdiw8aCwDoINb1+DuxyaKbEbtvxKnjpo3x3ErG
qEjjozeB4FSIZ3+hMhj0A2U7uMtaiKFxzmeCujbE6XSZKF+1oA27S3OTEDjJ
mBK5uZCcbGk+AdRKHNAz5UFLL3CAI+lq1Z73E8YfCJJKr8eOUgWVN8rrmt/I
SLb0OpwA5ZatVoJ1rJFlfQ20RBsqF6ekQBywIj3+ZvL6tUHIwozMDAmRDaOr
p1X1LLody7EenG/kHaXqxqr/wc2oHieUpoB68NPzhPEjZ6CyByh17ZWq/YgX
DhsXj+njz8wqK5mo//l1Wl3jHPW+XXtdJ6RDjCkuZvPrcje2jMiktikZlq+q
9b4LZWmikeLkk+lZbO0uLnnuUb/Ml60pFb7bPKPDCh9Y3i6vYwi8AJQjLFim
vgYFIXzrvfJ3Ay4t6pcIpRMbl08YH3/tCTvYIOk0Gtf8eXE6mbIkBdMJm7fv
XNukPEoD6UbpKZ850teOfTT5pw4lUv7Z0r8EgVTqoplPHmTLCtd4eBt8x8GS
noMfbQOgEYlyK977cDVIw/gnKVa0YrqRlFQRTia6oHy4QFgOd2Eo1gwKYvtu
9JtHcaO4juv0GcGvuDfTwcQ6T5Fe7h4FomQ5IWiKikPCK8uYuHJPUo5t6i9N
66s+gjQ1c8TV568nvGBFWHq74g3oJmy9qcIBIBFRsUTtDX29Wzl93bCFUNUy
h+6hkyDnTpWM8vzLU+yRiawOqT4wrasowHGILId/K3UMqwl9RIVIpuwr2Vgo
39iWZ5SpJX8LjWQ6sTQOhHT6xAE05zjilu2Uo/3GlhdXd7S5oxrgluUpWCnO
9cROgtBwK1KcMYbiZLnPLgSknaHmT3JPBUjk6gme8EqMoLGefkZXPkH/C4Bn
h4rR2m6U8C6A3Kz4sSToAdfzt1o9SZv8m5JJxTvjUwsqZn6eDW+iQZz2fSGp
TjIgJcV6tfDSi4pLBGXVsFIcSNvBSbQgiLiFQ1kvGBzO/NoV6Hs1IAOdigrg
EWan7JPikGfTZVKoqCrLdyHKD6VgsQq8ZEPWn6OCfvJ4boKOAkoDVOXZnaCq
NzPXMLComUWlDOZ7hPcbtkwR81qI/77lTEH50lRg2+lHUmpd26nHu0xg/PwA
PQb2rD7Qn7He7a+SlQb/m/VdT8qFMb2M3kUUE4tVYyRX+PQiJKcKmdMNG3Jj
MLjJ7HM7bsV4CBJfBhBuMUgS4ozwDdwkRBpIKdPaJwt0Hc1aWJ4pWUh7/1fH
MmtU+teuLt94GPZ36xnH6SQyXaTeC9jU4Q9OYFzfmxcWc96TAEp/jjWOQdeD
wRY6QDF5t48HPPbDl9nn0/pJvxb4U/PST6mlSPfoOihxGugNCJ8RFY5SJDc/
ru7Mw8DfJemJwb3FnccDMZDENkYCmH7gk3tnPEoI0PnbGAb4s7n0AsB/4sm1
AfaPeZk7wfX54Zh1/P81i6xNIvG0w09rX6NtpxgBEZ5hiCXwD4lW9dtX0p3b
cJhDd6kkcYewVenYzedx2ElABnJ38Wzc00dtbWRzznnBtOX0x8gEZilQy92J
hiI8FfCsuezPy9WURQry0oh2KJTRCTViOgQIB2bjDSVvOqi+f2g6W6SFhHAN
IoPFRyf1YHwfHCoXH0mP5l+iftxm1ubrKMcWnUY8XW+L8l7ZPS7QpPl6J7lz
hmSwiNwzRnXW1FhRve+8YtGqBe5mUv6gbixzDWoBCyBtMr3WAROp5UEz9i+P
b6jYVUCX22jW4kF4wElkyKSzzluI96uZnP5AlqvLMw/uOfscWIT0wvzolGxu
xtswT4bHVmE1ao3nPyEMluOicDCdpbV0FbUoc/JCUJn0vTr7BhY6t+FCo6cD
aXmQq0x0f8Dg5L0dQO7ocsSS9h+zUF+xiA2hyJdRHnGW59IAi6olDf2YxL0X
EAqGHY3l19RaHj5PUAp7uDbk0YK5MwEyiOkJ30osXjAJa5G1DvkNCZtuH7KM
Q+Ld99nQZtc5Qi2vFVMlCYnbU09rEUFQTde+VLaq85Vg3l/WUpqYv/JyUSNF
mL2HVxtD5XaHcUtPSkYWGdDY4SVf3IqhjPnMwVdRFiaHbF/OfBCxJ+qO7HDa
K/K/E+tlh0qMaBpSq9ZzGSQbefVlRbaMUC0I1vwbW849Ioi0AHb3eh1CGKI0
b+oBnhzFc1dkspGNjouXO938fm6tKsJMVoShlEKS13Csav17FL8Rw/MJVr7X
dzKlhtyTzA/YYGiIcOpaJLIo8I6r3C/R3BEkPYz/UysHeQuQMFdy3BKzqMGI
tVKazdUC+JVrr8eDqXF4WWXFoAgi3LY8sYXTY9kLf1IeoWhOfDC25yMWeVLZ
u1UYvk4wsedz+ueIEX2MlEYOY5TaNr33/kawRCIftvlMsF57H2w/X4ysEccb
C7/1kP9Zv0CxTrczKK9LwOu9w1Jso3D1t3ouoE4j1EvdiehiwF5K0rpJHSuL
M/X0AzkEILWbeEFV0vjVqOP8SrXueo+J/mrX8C5S9jLBMzBA557cbNIE5p3I
Y9zaMMWg3KQCDl/J81rHcOufrWybxDwTCyzg4HsfOOz5WT6cAmt4MYqinb4f
QNUpJ17nQoVyuym6S3EVs4nexqNZIFwKqZ7gjUc/zhsvjmp+TfdEmrvi2X7d
9hGxWIRnbedmtM9MAIXYakAC9dyEyCy/OqRzHqCHoECOqUNmM9yt+sr5oLXN
nOCXOPlb/e/mElPGtSk4cEE1srpNg9zlzOdOkIauMtHv609ty8jZwo4pdI+E
tn6JtG/2IY/3yF6rMDo3rT8+qsN1/lw82jrtevk3iYiDklqRok4FiSZa8nfV
9BvDIX/HkS+dt0aa8dXoIKwrNwG/Xhq2N0PB0LlSx/719NBjg0xaBCMJjyF0
AItqV2oBfroJ3gR5ZphMf3KZpHObkGH1MNsVNaggIPiv8acJZV9SWBvjfbT4
M8MzqGk3zVvtGmvvUON5jmVkwmSBABmkDlBovnoatoZ+oB0/Rk1tHCaosGBh
dPNTw6mroAtyNw8lKk+mKTuiO3/Y+1pqdW8O/UcInbJ8376bi9YrAwpDaRrj
MS5h0BxZ28+cDKIDDm917cL6iJ+qt8S/uaoM9qputjw1u6OLDcbRY6bQFiGx
U/OkLgSh/8QIH7HJeGWYdnG2/qcbn7V3sUjUNvRaWjRhiHMPCSPhAvh7srwc
hgBDkgmBgedO2eMnc2wY9BkYmJxS1ttpuhuoP4p728IftKM9x+56DFedQzUe
5lWlHnQ4glz4y6riURGdYRwcr29gQJ/bV5kWAozv5iFC4dWsDsoc1dqDq49m
3XXlV7H/dNZQkIHJ5xMTtUctEoGXDqx/NaFqPxSgKfl6+pN807jtVK2U3byE
tT1DJ5tmZf9Vt/ZNPi+3NqRzqX08HBQ6pBsyfdN/5d5BFpjfT/IlS3v1RaBG
RDDN8+lo99alu9k5/BR7XHBFRbgGVmhMxWBuuJxOtoKAEK+UiybD0OEcE7iE
AnnVjTKgmjGaVclCgFBvxDeD8EI72RuhcnfLNt8oAzSyQ9igjKPpTClgrFJG
05HKD4rpOOjyXkuO0S29epNTrQ/9N14k3au2gg3DlQIqoalwabK12ShJW1V3
3STFCB+X/mf2xS1muA7qZYpTd6tt9kwXMfNNRWLZ2EOTZSIzXyO9SVcAdFs7
IgsMciDj/dzzvStSaefPdnskysVI2w8ov6QWgU2npN7uUlvOpkAJVFYhqlLu
mBiuQAL5TXEjrSbC8cgSFF/3S6RSH55EoYsZTMmTgjvqUaYzQWJcXq/DINcp
RQeqlJUQhpvHg/3hVOg4DsKBJG4545lLs1aqcZRYxqs1A0g3Ztfwg4Eijw8c
R+C4NLdspaamBle9jjU/4n4P4CF9mT/gbFjZCT3TVlRm/15xTY57ehRXRGv5
ogie7B3lgE1KS9JBRqJARlnX6l44QDMr1aI2g+JXoY4N9O2Z+8PJ9RcWh3cs
gDD/qtOfQaw4dWIeDyYuzncaK8JXqrA7wqnxV08K+LFlInb1OmmSRcW2OZFi
pZj4AtUq3Tkv2GK1VoS1CbaXI9e8TPYkir+rnI3seQ0i+vIFOfEaS13W59VC
MLEAMUsf+qqTe1CsooQj9FPkisR5J3rbFd2p8LEJaXDY9kgATm+hHVifXBtR
lMLwTIpKuHAd/LGEvFunvE7u7v8AJGzdEXHc0W/3aZKIPTfo1ggRhuHAGkzj
qOzzEQYYOrUhTrUNijRHyZ0Keboptg3C+lRm3rHeRqImp6zNmQCDHALY+6XE
Hxx35xU6uAbIlzg1SKxI2FbOFEWa2q4DCcJaid6uC2Fq2H3kPAxfyL3Pzes2
0qm8vlG/Ff7Qx1IAaxW+j9baIszIRw/mE9Ai+HYWsyXqmlQiGAgI6ZySlFoV
K11q/EqYEQX3YCFXjkENNtFT3U48N+2r5+YTM7yiYtp+kgtAr351Jh5IO9eu
xCyQWBQAYKHvvDg09WF8RYQWL88hk0h+X6j4p7P/4c+5SyfgaoxR3rKWveUw
BZn/G3cIOGmwZyig1z7EPQ2lZ0YuoGfMtNsdHm0l71fIvSD8txzfUQIgxQ4F
8CBI8ApAdCrBENZtFE/O43dX8MST9sFXzHPbNHGbaDbFVyAt1CmN7Zo2friw
zAA6vO5hGo3GXDEkIBwuNRetP3jr5WM17OQzzqeEj1XAEEO8BiNJMVgN/IMx
pDMTmcQzfhUT2BjKR2GmZsZM65qSIUiUfnl6iEXoFfXbTYRfRF7G6DUhxS07
sANs0ohVHA2/lwjJe637P9BD/e1qeEbr+PzXyU4n9tNtUlb23q2MG0gRFYsn
b1UsN6U1weIga4GGs8l5Z2tDXqDFDr7h1t+J+enS91d5oQ6tDKZL2Lb6HThf
nwoM3SeQOktfD1pTtq4ZxNLPEF8M63I1+BdD00ni5PKx1BdMcM9wOSxcp1CD
x1BwQOX7KtXNWXDATpf1glgt8gbViKHCgB6KZ2Dk3YYNR5ZxcbnIuTD0dPKF
G6Mj1EsfrG/dmxbo4hvk3U2bjg0PXh0RimuXuoMe/wEEWwuorwUcss+50E7c
rrjkSSzwO9BDHUomA7Ka5cI5Q+psv0r7KKs58ZaWmiraTXgGHlL5XLJYsrrp
2GfuoVLt5xiAReQSHUAeICoXeaPz03panbSGvrh40VwjzIbtKNE15vRfmQ8O
NpzGDvuSy9Xdu9iVrKDYxjnd5BNgXk5lL8OOTe7/wW1RlLIwtJztouOM6Wgd
GDbOIVtSts2cY7Dr9F01JHbTZDe99KzkiarDdevh6tMRlhrVD/ndsGwbgFen
FJY1ntv3iGxwgxhPxhh9zW8Xv3uvM09DyUED1GTqKJkaSWmQPHaJHddDrgaV
CgvMYraEEA/fS2KM6T91rBF5u6eWeDQx0QMycf0JdZceq0TjoM7+KHwU5CAg
QCGOPQ5mKQinyldYXpsXnk8AXhUimqikx5Lth2LVzcetMYWz3F8Y7RTQP0Kb
3CVO9hnGNZphlKFt5JzG1h4kNPLOJFr/OR7jP66GaoygZVVOfmRRJeJ0ukY2
dwbpw0u5QnNXVn6FZtNYoT+RE1Y7ZjFeaV3atQw36ffh/WDDLr0Qk2vTqthk
zpMzqp/jUU8ZUZzjXCJR+oyuYaT+aq4um2HbVzs2j5eAlrDWwmnsFgyKt1vl
B1jwN5VLjgnQZOeF0TVP+vE0VLM6rhAKV+5oVdb9urrGchEjCD34kXQ0rS0p
3tmr7y/TTcFHlYd/nxx6m+QpK94bPIPm4ZGzd9TlEjLzBB9CuAvcVWRG7HM6
R5QUoq2Mp6OMtBMUVJcJAEx+SDjWmRwi6+u9qbKBiqw9hzsN3VTj6qPTKIlF
feouwRtjWHX9TjHsUOX6jqX/LTs+SlBe+kHLfZkRwN2uY+o9nIoglAhMTMS1
qaqo0hsmid6BdhACsuqhlWnimdLo5fZ5z8fn/8AXiSN4n7WIwmwWgxDC6BKh
yPGV418sUU9hxSKyRCd0f3ahI0n2cQeDvpphDk51lr574gGswCOGjGiUHmlK
iuTue1TYCtwLDT0jkrZiJOEM70JB+SV++BZPzWc4FTuovKfyFuRMi9VOSV0n
XDqGAGAuLSTNZXXGCcCOJ/Ur98oTHZyU+i1CkzbKW4xhck/KUCT1GY+jcEaN
c+vrrUKHg9aqreAEm4uJh+O5TxdsR5/IPojzkpca+qi4c9XBT1CepcAd94bX
/o/FN8++BMZVxaOxKY/YQzIEs4fCyoddCbXQxdoh9oRaUhLwdFwx5z1l63pD
QtQd8nxmSKExpqZT1102wTYM47rge9a+aL8ODFDAeQh89v7WLH3J9v90D+PR
l689u/j07TU9U8zUDpKWB+SCZlA1OnQYfHQmnP5kiXmyskiHwNwVvWnljKBH
I96nC6mO1GyPYyKx6fOia+MFhFJtxTk1RkZU9CwfIOAuAQ//XIBbYN+UmRJa
4H4Rl0ssPoelrAW+UOp4B8yCtn559b+L3gEUabTIK+H60hix2K97xWm0nP68
eyJE4ys7OzgvRksDuqKxDNrFRfMRvcs/10miLlHM1f0aUdBP+EihPCvhlhNP
rdvoXubst4AtJZSCv9GfNfaTOOAQxhK+4vsF6UN9TAkMMOEN1PvSUsUUPa1Y
+jmX42jd7FR9dRwsxhg6Ljej1Ytbl2iP8ssBX0goVg/nJ/vg/aUlBvnsmnrl
zh8Li8j3/eftzNmvZONZWL1HSSEM3nWH+EOqD4RBnLq/XnCs1c42GYzsCBno
b948JBu8Lh/zuTpJbYz+n2B6T3/aFPgfP8T0nESOGKUXRQpbefNUHjg67LP8
F62iNh928YXPLBOzcHp4evbefA0YULGVXWVm/zDSBg/8fTSrKoQ1k6XRC45b
OuUygI6AdLUTP4zAbYldxAFlklIsj+ErSR14bZoczsIRwuhdK8BomE/XqDJ5
SmEipAsBgU3LYExRbBZ2OXum8YNjSwoIVsLnf/4Ehv/wuoOlxNH4ONInUiTa
oLVYN/ZuJk1YHKbeMqzWjQTIJ1rrrI0+Zm+ZOogmcI/B7VISmuRbOa9heU0r
UZoAuwII5RjQyNvis+R3nG96XegxmR8mo07Q68tr6H9+GbBDaBBcDwQvUjR4
ODJZGVvyu0ILzCT0CkjgJQdQ1lhc1ozqMqQlIgw5KWWcptdzDxRreXqZbpZf
GKMmLS8+E0PR5ISxwwET28tR6/MDRRWwQIZmg1FG1GdGomH3gMBxrSTpbCPH
L6PXRInqyPOMazi9OaxLus4lnHmb/OKKSEKiFCOEcA2wpk5j0PnAZM8t9bMR
APd0VVhSecmARlRl+PKmfxwiX2VFyHb4FXQJnQRqX/s4l7xKdO0+/MuNjUWm
0QsTDdRVjiJxoz/JNrf6n5wEKkclPmkXCj6cOJ9b8wf/nsIp7ifgGBcQFFQb
SvEVTm3Dvto1QRI9PaIx46Gy4RRUCEOqK4QRzTDuMdP3FU3faPPL/W1Bfc4T
iQoVKzbV5g7D+Vxwki6y/dR+6fj6uOe8ueA4PnOlHtM7NI5fyxFTjM/LuECu
zaLPFSjkXnh5JoBMoOc9SHUlFKza0TqJgvF0kYc4MI0Zk9Jp9txKOyujUcBL
p1hUk2Pz43cilQ/kJI1pQ/dkiDgFilRYZdUR0xSzaquHuBLTnto1Jik0f304
E7UpV4FjxzwFVruz7d2VcgsIag2/yktZ/B5UiAm6fvxXsZghFBdZl6u/Mss6
WUbfRBCqb3NK4ec7AJcVvBa2DqpgVpBKW8TBvjz7F5IuXFitWo1OHn9PrFuB
LtX1tKF3LODSsP+E/wY9KGuK1yoKaYMnJV+N212pBUfq9b+76HZ0e/c16oeV
NwfboQsp60k0LFxswBshBxVJw7My83fyURBXCxuXiOLxN7wiCBuEvRaZ0hfU
UHydsHqX7FICIwn4hop5GUHB8uv/7wGP5c17qRF0nHrVGjOCKQbNdn5KGeVN
9ry0h9MoPNf7Zg4T0MQuMD6YFzqsysbNYelcD/gJzdIs22kAhafarCYEbKZ9
woYOWGhuEzysQDgLefWFEipkMlSGc0z2LsKbMyBEc/3EVGBwygcvmQg6MG8P
2XPVRLOLoMlYfMYDe2veaJV0hb46/n0wFaakVSMmw90gNlV4B17df0KvQeDo
WoJEtDOorseEbe7O/8iC3Drmps6ky+prAkNOEiQ9FOu6TLYBSHfJ3XpHgUTc
H/zyuyR6AkghC9B9SzZFvStU0MetYYCdDEBB8J2Xamlgs4Qb5QxF3pcKsJLf
lGqGyXgBYfF7rdj8H4SIvLS57X6KU7TFA0lgS4lM99n68Icn7RZtqNBbLjg/
9C5ODc+uXIE3+wyDNAY5FFpqAkUPZ1aJm41oep1sUq0F2GGmm2iNlCKzV3tk
IJJoPmhWGve32KjLwweVXy1Cl1VXsDXgVZD8DKdXVTNiiZ+LJIfm5UdFQmJU
I1dFfcT3G8pSnLxQRtlcPy1nXw6P5/sKbKUij6hCqcqjdOmnMMnzB7XLk/5K
2Ph1xHLXftrjbBBzXP43bPSbPCyscWysoKrEPw8ThY1ULfDMxbbO1Rkec89S
rRraPVVK6EuadO1fUTrHP9vqqPBzd4dNyc9bj+oBG+VERO4OxxUow4pEnVi+
2bPVJX36S5VSQ52Jv7ZOoeQVY7PkAZ0TFsXUxllBQcQ2uI/7LWMBmM6r5UWM
yI5Yb3ljCvdLovO/aruknoqGKsMjl+kjfWoxlvu04u3jsx6JVLQ56ti0mqGl
PdcUebAMO/Hqgsl9uyMfjYtTPsgfEDho4D0TT62Yy0cxjkiQHs+KTyuvzd1E
g05zMTmsmIDp0/WB1J+9bLS95OzCza3KZ7x1/dwZ+DqUvmD/8GADI4u7uK/K
CENQV5d/PC6PiXt2iffu40UCBZ+7cHiQJUiUHYJ8yaSeEuXVmShvcvTpkUXY
j29/JbyO42848U1B8jmQX3BPPlo0xKkeVmj0ET59bU/fInx30NscxZuJgX0x
APnrl9d/9IA4WoPDMnqOTh9XhtZyHVCrKJmDYolhRHGLSodXvOSQzru0wHZy
qpJ700woJiqfQ0fz99ypZcWyXl1A4OrfUd/i7lg7NJIOoQN2XmwzrSEAatAb
RN9ofG0slluvMK+H2tlla9P2WjDVO8diaWBCgMJQE0CpDNNUDypz6tDgSwRi
enPzSvfDXSynqh5U3VS8TzpbQV1S1IIne4h+GrlNEkR1IJyhwlHzsUMAGt7S
FCH0/4GMyEQz5wRIIYFYNfjunS376czNS2M/h6jduDreuyk3nfQ0PY6soVOJ
gIGt50o8X1fZHRoxft2xVzxGrz2n2oxcVthjz5ybUnznKJRpJqPvbTWxe7hA
OSNbU480ar29xu/jZa7fgGdzFcWyqZwWPivsCguOoCsAdJXxOEcamcULvEhC
bJVIOJ4apcwHL6uFcyJDCos2krj+Ob53babH6oFRarqwc+DgIJW1PFCAQ4sm
k4PKww44nD5JCcBJfgAHIIF47L0sigL9lsmDNXfgj+EEyvXLy6/sfR/hOEuL
kSxlNUggbFljscwGRZ9DqjqNOsZ6mIQUdsHk0tmHlWUrgRreZ2Ec1fQQUuKI
lOMxTVL4zkBtcxrlRaalZBlHTiCi34vA3AN2IGrEhXWPxL+1z63KPJZgBGW2
58ZA6gOkW9OM0PBHxR8qYvKH990tswWCYTHJJVPRU8EK5PEM4MTdCnRBCpM4
uMlUVWWYQ2ZEHwMb/by8u2k9sE2+q2I7wSKnQA+m2RCJTSo+PNW0ek+STKP2
uWYlRaZgQNNHPUswD4PXoTz1lXIxGUoAU4AKfnVyVp7WgteKTVX0uqn5TETl
Y7/DotmN0UO7RVAvVVKoq86EnuyMDcl5zkeNazQEWaTCEMrZPDZx7dMsCIge
+pOmgAUj2kY+aDxTZdmUYv1hJq0O5zhm8x5oTUv+S69Tn2bJGCxLv929rh6G
6N08sky5W5Nf+XhaTBb+8OpZfrjSrnmbMM+mWWbLFdvgHGIZjM2YbmozrlEK
wp7fOGSbbBkxN4htL8K3hKhzGMzYndMi8Kj20Ig9boQQHdspM5oDG3D52X9Z
+zSOjUWevTBYQ87Mx9iurl028fR8PF+KXyzUZyU/y2brhv0e74qdTT/uyPV9
UKsYYA4C/W2vUEpRpF8wA33nBjNKdmIAMvnNVuHGZUm+tm2wQGejGJ7lfYCV
sjtjSjBajtqb7jrs7n/qVPYo2Ero5eNb8ldd2BzWsDdPM/9wWfjpG+YfxVLk
PTF8Q3QGIGDIqDOrtSkFO0FUfPXwJLgiuaxgMKKxpCRBhHiN/+FgCLtCt/Og
ADF3hqSGhyzus0rOTgyyQknjLdh9KB+urzXLa1wPQRddNhyeymerFsZfzmi+
aMz7VfhI5ssASb/idIWYRyLGkdiv1VOCAY0q98TWjReFzmj9/laX6+na4FW3
avLtZA7XKW6hNnPbrG2DqBlsNTbapWSXMqqxToiuTZNaULj3hA+XsoZ2w7Cw
faEwhBb4Exj2rzpOrzaUa2pn8ccb/oCYXqaII3N/dWOQ3DeGUTB+fAOS7Q3F
+H4MzNsPQE1JbOxhSZQkH+VHZL+GebKNXr9wNjcRYhpvRp+hmAENr4LMkvDK
ByJwtaAMcdn5OGqaaIb+Uat+Zco9ndNgx8Kbfafw3QCfCH2RBZL85r55guG+
LsXxwCeOJqNVr61PuyGgIiK1kn6Nmk5zTJJY5T5NfN8cw+VfCSFUDbJg1mY6
Bsjb901CIA2SPpSE63DNyJoHnMNFBInXYfkuHONd4dSfed5e7waCFM7lIefG
QLlVgvMZmY7aXcChiM164LOv7dUT/h18sQZfZ4ZDmAE5x2D5YcOO83TGPVsd
OghYYGpA0wdjQu/HSiwrNwlj3JH3rowvWRRQhq6dX5HVJ0lbSJLqlJWVaji2
oSVDh7VVNaBoYl0SySlQTnhl8KQxEZ5qtlmqC2Fbdpuk5Ry0rN7UuRz/adkT
FeE9tqmg93aj9u9jUj4nYMmYy3HTHUKX+s/ypoAtaA5Fuv/hA56nWqQxqAtg
SPxk/8Y8YceM6cL6W478KXfntnzo8cddVkIqo9/oZZtKIqPwjTfRQ+vRF18X
psxpvVqPm/PrJHK+V34OMZzmNPRfObvd5sBbG02SHcqb9+hkHjKFitmv0pCB
5r5J5Z2z+VsqHtrah7nS9GRrEzM0TVL9Jf3QhkvCevdDWYdFnRQo2v+liO6d
aWJY/lywAaWc7UQCEet9hoGNSAE3bz8jTcuueb3KoT2QgpNpzeUzSQMCUWV0
/h62hBwtGqTOr5yD6QlJwOdmlSX+XUWfyrFovXJpCHKUGc4pf2qzb9ydJuSo
NvRMDbmyws6h/xxBq6vXC8RuP6DiYNZ+ZvZqLXpOtkcl4Yt+OSMF00jBnEXl
TF0XvULiAWD/Xf+uNg97RsbFAzAPJG7mtnt3ztiSOpqejf317eoy/l2KaG+9
4UOvJhABHMc56HYEZNfJkl8oTvvSQ4TPxNP1C9pLuJh1AE0N4GxgnfCj8/bE
DLXb+mzRwKq8I3A5CZEADm693qvy38u1JrZpBXV8F+LXwATgYRZBCPP2o0dH
cipR46V6x7YKjDSI2fKeCV6OIFnVBV0Zk/O2AZdr9NEOwyjqk0GoqgzxTxc7
4qVJgmULMSg58gva/euXFMdj1pPUiwORXKIxdkKv3DitK8Nqv1Gvpdn5HAi/
ETw1a8X8BoYglqumPz2pR321Z7KbSqMBQnXC2VtVEpB2wyJm9j3XAxnT+6Kx
s4X6XieJJTNQkSl1nCbfGpBQST0eXv9D3nZB5PPm4Vr7tO88uAo5Rk08q+tF
AJAO4Z1YKqrgUns6BXdsoh6943MJB1uPymyt4cAcc2+EB6UgWAwWAqimbPeM
KSYuE0p0OkL6d/xleybqJJ6/tNHQnv1lPwjsxWmKv3/x9F+ZfiZV1q++nIQ6
+vRXXKyUXMHs1+ajRYwZBpp00CXvSwVTWWlAd1Of2FpsBID/53SIIEHrhCVg
wECsyroxr2ztRLajvK2DwbXOEYKMmUhIGDSwtLzDCd5YwuLYnEu0ieIx/BuZ
ks7kczGJLbTCddKhTSYQleZS5XdAu9lgCUMRtOQ1P+3lw6AZJu9Xn4W1XmwQ
gSY+BxdzNSfPDGB+cx3vJwq3MCpYigzoIzpSWuPZ0VD5fvJ9DMNjyuKMwCeI
7R9fFbItaWtaQjSs72fCy960ujIY/0ntqMg4th1LRR/B0SsG5kAOggUgAAnn
4WEeInqezYBGOOnA18fBAmbV9UlwEJ3ae8EXYdGMMyzkv8x8nOzIZ+vrR29a
oE5wEUR6WpgWqM47nsygSwVZLUd1yTt69nzLRu5H7jym7Bcv2ui3NDnIEDr4
lvgZ5ybyqMBk6qi6POLacuEN41EqkeiQX3hA0GGmTeKI7PWkBbQahOHCiplT
MtiuxYDCtHjYzMf+gbzCFjmtdC+A5HBzf6NSMBTM5NzEFj4FEBN29VFVHY1z
NhE08zXz15EuHsCe/f5L+XHeAbMMeKP96Mz5Q0KfUjID+dEn6ERxy8o8m4jd
rtNDIdGJ2rRz+XnhsJUapTCd09h9zGoMDG0cWBMNMtYbf3KABmk2Qwgsj6F+
NTgV3apEAYK5btCsmatlvrRxvCTe5az6WlQROvWwqcu/lOb75i6lFoDYGNy5
/MqPOTooqo31EbCwsQveLzZjtGqhg1unWdsUa8MFtRznPaDLWbng/0sJI/zR
mmdajdn/wgkFVJW7V63nqFdPJ5jUxqDHzxQI/EI5d9E6QwbeQ5QO6na1xPZm
g/DJqxbWdpuK+vJDxZTBaERQj42w783NYjAJId0CbG+jLWEO/5QbxizI1qnu
1IQc/An7qVR60PoX6F8gh/JS2lDUmuERXzIA60cMX3D73Kb+XkcnMMEaWJCu
FPTkr7iJWT9Gv1KQ1hrZ+8chhdJGlOLWv27WZoKCQC6yDN4BEHWeGQd9AbHc
mXZXSBapMYN6PrLDW9/PVQEttMuu2SAYnno9EkNNrvkATh0lrxwK3xXC1wkJ
YiezzwJ3q/5BKGDiFWTTCZfTjzIavBTn7lDOv+U4hGigNYInUTS1Yp9EGtUm
h92CtGa8CdZ2OKJ08qQVOk901m+c3J6uARt0OpBw2WhWb1YThElGJNIV7EsS
NpBcReCRpe0hEsW/5/qfCxSoInfp25WmGvjTbqq71nyeOzUbmt37mTe5Nua2
C1WcsRb9A+MD3DFQOqjA6xP9x+SSNYjk9ir6RyFdvgD9KTrije1ocel3Eowp
dFslNv3KdkT1P9PZSebVW/tMIK+pY/vkkfdhnJ42N8kcf+UVcrH0hHW4Pp4q
yLUy6cvdFIqPaVaM7yGcD+CY+QMbmNyEYqtKkPxkdoINgaZYhGpcbdA1jy9l
3zcyUVbDQl6gITygWtFe1VCDMbxGCPknd6hzl3CW2rZMHmtPuGH64SovnjSK
alRarY++SFlwPsR64JXXu0uGjGky7xWn4nIrlK19UdAsyNQMeRPBTO0f6AZM
NCh0bW4vzhX4VbR8rZMBIR0JvSRDXELeI4yZXbKRfyeCZzxqdSe2RYCs3xy2
kz40mc0+1jXhGgE8GV5hhGBT63wewSMRJkVjuJhtZMtEi9PklhfBHvDSsv/J
w95LO9EQF3zAXJuLqhGXmlOk1mVf8T31tD6gwxogq9cA6jn4QfIJW5ee62mF
OLCs+FdQyeHwsQQXHQqLTJuAJPqWMa1u0z783kF4y5qp4kJiSE65m1NLAXDs
ko28sJnE0bly+5ZT5P4W2pRW8bjuCsaAISCgLnOvxSAaLw56fQWPOI41IHdD
2QrxAqXjnZWYg8F9WswKhqS5W3iUYbPm6mCiJXdMrVGcspMVZ/I4oBq5jyus
xQcLaJZlxwnVu0TEtsH2yt0AEYnbiobqIC3fGHp1UT7T1lsHsaCOKbPo5ooU
oVS2tydtZarEupOJQq7J3NXFFoshrIPewgfC5yxLTlnjIMSpSTRc4F6+afTm
zG7s3d+ml7QTdxDVoZI7KqgXV6Dbsn0X1DtMNdO9bf/O6u8WgQiwwrxJ2hzW
rZLvgarBLV4vtWOg83bDguCs/FP68d6CvS/2hgxSHh8CC41IOVuchOND8o6y
763gCcufTGk8e3Hj5Wvwo9SPwVSQ5OTHh83UyHkv1QzLKhT4gA0t4PwHsspU
rRiOmuAzrfwjU3Ebp4bxzJrMzFlT0eTEYvdvMzki0haon+FsFzshBOG2zSyt
WnxvzfQOnC1Ugj7bUjYW3LyjeLIzuXz+MiLjdYaWaWGp/EaWMg0VSib9gwa4
dqSU+bTYJID7GLxnvCO29FiRyhCEtzYPnGtZzKrYWFKPAaWhdwkruQ/Ofh8O
in8Od61liL2Vmu7dfp2ftwOHTQIkc29oEuzILLIfdpL+jZlQQ5qp9MyPkrv0
PvNWUEsmetdJiEx677f04G4iRTDOWeZvX498OzwCXo450ftb6z6sNeKP1/tU
Z2rfEYluee4sxQiSZRgNurUKrCrUno5sFMnYx/PFhkyalzjrOKKQWD9UGTj3
YazFFH0k7S6MAbiHWAn4rOqrz9mOQwDUgB7J4hXNC7grk5k+yFfjKaJjpVMo
9mZJnV1v/HNHdqXQwpuKGcu09W9ZvREmYORVS1DqWgPXH4zLKM4lrbTl+GeW
uqtlxI/MWB1fhKjMt4qWRc99GLso2yWVhiYCFj+FEb49gQsYQsGQ9mI+DmwJ
9bWPB6qFPtB4NQ/aZGkRwIjRaKNKvS+zObSxZsciUhKoGmzPRn1S/s1EDaAb
TeCSb0JxxlVTfcABK4pIVwYvLsbMiOf+igtglMTdY5Mf+OBzdZ3g8DEde+2f
89eI/SwyB0k9DRrN30R0wp9HZzdsh4nfU7RY4dYAUJey5HdAFgI5FSb9hFeA
eF4Axzmk8VBHeprRFNdGwCEw+OOMD80iI0FYKO2ogL5chxRYYS7glA+Ofxdr
Q8TQYF+voQ6nkIy2iJZqsVyuZWl1g9OQ3q3+1Nroia7007p1IqH3RIunG5HV
06EZ/eKEI4gcxBcEhcdNq9zZtScisR7G6ATOeEQ/qEwBzQ+8ZzjMj36ct0Pv
EisvYnNLqXd4Meqb64QpWpRXL3ZDTezknNM7aTpG0DX4dzZa11o8m/fBAxyS
LJ6+E5MugIvb8zL/3qqIgDHifUE1qktSB6is2gmw9ULqw2+tPd39XRW1eIIZ
4n3BwKGJPuLrlz/OHDDCkBKOT3qaFRp7NZs8TTlVqTYkKYyXr0porDMtcsSD
De0p1oy8YwBv5mFraJeSznB2NS7J4kkA6kl+UfxXRDfnC+z6ek1XULd8EL5Z
8H/YnQ650hCe5SyUAvQxt9IlubolxoviYbOCMrOzvVPdwigknBSSVbV/7r6z
O+6DPV+JudmUO/lM44O4PNqu9JHKiAJd0lbjnFjEyzBceTjJ0eLtCSUghdJi
3r80/h5sgEnS5ldvQ+Y6pOcfPKksTtCqCE4RM/nQipEPqOkoKDPq74vwxD8k
MQrM0jcWdc1hwaJnLeUhpQxKpsw+vcGNZfcTk85wRRUCDzUcwyh4T/elwWSL
4BFmxOcNTmo0OJ3ViezrGd6WI/OhWWhCcakiphgayDNQSf9IlDANvwxEeFld
CJp7QicruK+OrzScyv9WScaO/4qIsMxYkv/bPm8SFcD4VrXDwLv/ivznEV+l
Ed2F08nj4MGnVd25XUYVwVpyiFXP5UQQ4Vew2+nqJ+JsCvEZULVOYgYtLzbz
BXP0htiWZXJKRuvKHUcpmj4GCPdyUhe2i8yYxdOrXJRsrG1GAmqTIdvQmmV6
T2CI+bh/rV+yTgJ4/ZjNbH3TAv5vca+wU8c+AA6bJjiAp6SGp+UNRnwDfxR/
GlQQ7o0+RvxgBZuTPt35meoT8uKixF1cx+FpfaY6wUIm6DNsnvC0UIg8skMq
/0oijDmSoUcOiwOOEArEYFYdvbhHe50+p0Q0psjGANE3qVKq8XH2KeBb7u0R
2f5ssV0zNo4CFkr+aqonQZpp1YGIEQtVnNMz7Bv7a/wukF0fFC/eH16LtN1x
GJVqhJUXii6fr2+WwAhGsHDMJISkEuaxKfxGz83zYYHM4XMuGjZ+UbOFtbAE
eJqgY6xPurfEUbWoZJBtNbuOAXps+emlh5vBwcZ8hWjGrviaML/dqm+Z/E2B
tejLJLHTrg4SBATKWqpnLEy4r/Uvei+hs25/aSN89qG5TCuM1f+e8lzGfS1L
JisGvSchMyGwo/6EOgyCILcfK4lmdqPZrtzrTXhpR8ok+3yFDV3j5yegTuLj
3XxTejlYNptQpXp4JK/eTlmI7ECYonORan14rf/qABks2TCftcedL9bBoDgR
3VxoFA11USruc21TZCPqhSfMK1YEb/1cDZ2R3yVxEYY6UYoM/TIKuISAzce+
MJReo6ACTug7GgVx7Y1FjxLkGyd9y3tHw7Sf6d9Tn0lC9RwWP4MawcGPRg4V
bv6+f12Nto+pf1zeIRb8yvBIUWgBZcAXIBBehcv93PSalvmP7xfH5IF682XF
waW+6UoAjLcw0lzSoNdQIh7V3hgcMFzi29BHW86L7QuOsr9r+16yXKSHteIG
1KKqt4u0Kho1FN7oRluYYq8jvaNny102+M30V6Ye2ERxk40D+FWkp/IAYmhE
PAfCz2md1XObtiDMxdBYbCNO1QjSVSXXLPBcDw3FmtRRKOF5Z8MY5ITwFo21
SpBOoQMDYgm9cLdH724GBtBXlsLM5ZcXtaaRNcUMBNfONi8dGNFXlrhltxBV
jjQp9ArESz1pjJJQrCq/981oGPX+Lvp1cbcuGM4UNvJUPRb5+ky3+yQ5o8/u
d6PlgjmulYPJN6jMNR1G00T88yAg6e8yTH3aLwUkVm0Htrw/8L2YCGd1/ukr
KW2quBnz07j0ZvJk3yzoHr1JN8xzVs62DHm2Vk+bVpKV+412BZpM2alneizX
55UeqpSNKRmObZpFhiL3omdnbfKaAWNYVJsy0Ob9AFu9Gk5DKA1MrjVnwDS8
PpvPQutuKfTtP54x315S2w4+Jyx1RExa0ctxEilySNySfpqSeZrCmDJ5YdLo
5AKaqlvqaXt4jHC8pE9WZ8+Bq7X6a+azRdpvRclM5f6Qi/c2zNv1bOUyY24J
abuZvQ0Put43BuM11OVNRAV3yFDbf2AmlrZVU8ZWeLz3/fcMJKPIduhCW9Z/
ncqfUTPOR1Ywq0MUex53/VGRY6u5ZixLwzgAajc9ycDkOE91sAmjt4z0b02k
Av++LyjK+l6AYbXDzWmbk77h5DUEtiJ6noxlDNxx1hidY4PPrHKPWN9uXtew
bsYprHWOAykk5VjSSZe/0l8CVhokYn9LOebJpJwYnePKyr5DbsHtVHQJIFN0
Gplhwh+aQSo19ABgtZPmpA1wSW0lxyvSIjEUTZ6AE4PMaX4Kao0Xg+v1H/n+
yGQ8pBStMMZ9w8Wompb3hqB2uprixDC7gribSE+5e4sYxF9L1u/Vuok5aEmf
OeOXTtf3Qbs8ei6xI5dTHEZRoD5iHAM6EJVtB+nwCL6Zo7mnrejgzftQyk8S
6zzP0oQsLTO849F93GUttrhvAZTE7yRrOOB1tfMpRtGGrci72HVwu9XXFkl5
UOLY88zj+D0ICi73CePALPyAT3hm4Y+VTkjWK19zSOXqmv2xdwykbuMJZNg8
eqOlUuJCnYS9GKRuVgC27uz4CYSVzjaw67ZAt/Q9LisxePIviWiqTVrNH9+E
QFir4uYLUYitsUR6gbGRHhMniy/A/0S45kaXizLEiRTHiB/DHP1S3bJSd5rP
3XSnMWoSxAkG9I0rm1JeECC3iW7wCVCpAI55YnKCApTIgzGf+Z1a/CZ6yT7D
5xmmdmGWIurUjTxxYXU5xozqhp8xEFu87ULEBya0KgQE3avc0r4WXDrJZwHk
Nu21FlAkbYB9rhQdT07NpnBXXBM5ZU5sQaidNfw5fAUPOhtBitCtV2BHuhNr
0sCrC4QHEU7rscG6x6lxqnzrxqr/0U4PmSwte4RzO6/aF+LN2uopEVIXk9gZ
Dso8Y0wajbBxo+qrnzDXjaTXdEC8PP6/Ad1Dxw2eB18gASeMYm9Us3GbVWhu
4pqR5ejbZvs6X8nNz/gCvZNs8EUDS89i71M14vz/aWABH0St+8xkgFs1hHf9
bKeMWi7/nWIWHUqXBw+s+8/G9nnrRT1+kb2/qwGnxFWAowF0YDFBHLObjG6Q
JgOuToZwg6yIJ+6KN9SOEGM3VMejORd470PpLGYEMZ3q+p8VuQWmQMjHMB4d
/VCX5juLszaMXyeJ5rDQmZogMHR1X3VIMx3/muJrXDjK4riXBFOMkGBqtzP3
jVtT1CExysjQt7SrDSB9q/CrV6Lcynva34djx6B3ayqKz14zD3fu6bAwzm1E
9B3NnS7Pg2wEXfg3YWIfjlp5+K1Ayo5AiCFvT9ptODz2Ye/8+gJCac1eyVLc
4viTtZF6SOkXZE/5uPzGrotZoF0ZNyaEbR6JV1EVpORKo00ZkiwIUMlbQkhL
c2KpFTgxDwrA3j99Z8Wd9oyiXKTv/4zduQ1ZQwFH+MkD7HiSFS+rVpLvLJb1
f2BNrfZE0HC7mj7OiKanpLDtNC2hTI+DWUjg3l7A9ERLZeiyTCUGryISqIhw
cfhiVpvo4LtUP6igNn4ceNvjfhisJQvYJ3VN1O/Z4S6u6gTk9SMqWmhSC3VC
M1QNksVBlkxFIYBYboRb2/t0Ev2OyjRlPGbfKeQP2TYqNo89gMyYqXm4UG7s
Zhl5ksEP/pY7uoJ8Boy4AG8dDW/kRnNknqsBBu25TK+rJe3rT6/RAQwxwrFX
r9IfSyN98KceJIwnVMu/OmEWr8CgTt0mLofQRqkgEQmRME8d4TqarP7hD4uq
XQaZodQGSZ4kg7aR+uUphZAIaYkezTnI2h/NAvzuK3yavHA8NlFEQRPcVlBi
kFA2Q6ZUwrhsHJrDQmM9+2iNL38M10WX+7RtHgSJX1WqKNYWHJkF7iysWn9g
gbI0n/YkEDKKxj48L7992ADzbtUspBWrdOZ0PKKaw0MourIUhlvaYdUHTCwi
KLMBjfoQAY6MNQjKYx8sAwHVS8kDFJUN8M/W02QLmqKcSYoTZZN3alJ9UMu8
DmYTkUhPlQcY59MsxnNSCgKBkzgkWcb7ArnT0dQtQU3a9MFkH2bWX2mmazaV
CuqMEIaDIsSdLacMxv9k7X2RLPiTQFIj/NbDwXnnElEjaWVL1/mVbjyGiSxV
AM+IjseF9McuHrHF2NHK5iGOEpnT9amVzIy00p/e84Ts0lxRl7gHjyW2Wqen
ohP2HIKnnTPjRFWAc56sHpNx0bk952cUtoVRlDRMCFUAc3vE9J2eJMUikP0K
AkHrQai2zkYJUWBlaxtlOhN0ewTneyNJh6MBpVqGbteQSK9OvjREGkAhHD/I
u11TRXUhf62f3OhTQqU3UIF1Y+2OstVmuZPoi59qT3WWsP4lvClH9F2b/Prx
LATW07Ob0U2Q+QGBYAYTyiq59CN+PvDnJJhwlKBOlaki6uGWhH+Kwzj5n0FB
TTyiO5H9SW9E+5ArW6gfv7CkX2yKWDz0Z/5Tf6p7L9/HJs4uUz0nkW+ANlZm
nSAdblSembdougRidTAw7vr2uGOy/89EALBy9Od3W4tJTyps6jAVrOk0JPLF
0FfZPg4MWLhdjbBzs4PgDbiH1ZaN0tziUAqYmhBVFCR7jhMPYOKGs29+931O
d4VyRTeUFxgV6CZys7sl5nvqDp9k13qBg4PqVU+WQodVuIAXwZrCkocY8sKH
pprgE73xckfCzHAzvhrkwT9bkQcUzOgmbLJEAUPKnVyYO/0c46tIO5wxoFUK
Mqp+J9ssfhvxb9Ufr845P5HbcO/vjOlJct3cCv+SWH2fGW5xcaOZ7ji0K5di
2by10EU0zgV2z7REM7jnkADQwU/ZuFhDmTaNlZWmYfMQbxzpvLi0S8nOi72K
lKwxbMpoh3IYYoqt/8ZmCo7gsODcGzVJLZ5nto4qeRn01jQCq0NPg0tI2Fgx
aN5mFc5KNhQ6iYjWG66w5KT6X4CSwVLEsmayCS6TcjZFzCyDwyttBDwsbiBa
xPHPkLjONMiWzP2UI4iyE46SqfAuKhpGIsoAlVCbtuc/N5ERWoaM6XJAJSTZ
r6NN7gDgKIhriZLvXpJUm91iT5eL52Qo+KP9rS8Ri6eiB46WU4WvIpO9RCYZ
wqDaigj+iC4mOrkOfxtBCsY/C02O3zlMxqUjlbvRvrMEOkfNpVO8d4gQAdaa
WKmM85PBDJBMzt3wAqAJetIfhxeiE3FCNv2pddX6UBPhtdrADSMkxQokInXR
LprPBM9eZHyYG1SQ000iEwjgqfZ/hVgr+862AbM+nb5b2Xzt57GiJcrvLCVP
1j1kduAB/KX+2speqeqtfHeKtsfVG1mYuCHjjKq0N25bDLaqVumyF+1UxcwU
DbK3HrXhKvS5sLEq3auKbo/fP2xDJepHIe6eWvJUD8u0FTeS9u5xa6MODuci
24YsOjzZt4YCybzUkrLPAsi92z9xcom4YjHv3GDUiA9dlV1a9yl+csmZzbRe
vtL/vwWNwlnJ4ktCESESXN598MzkApmAZQ9HvLoyQi7Z5aDJMqHBpMiuqEt+
huBBeENgG5MuoEftc1pat7qY1hTJZAfa0PasRlWO4IMIJ2cesP9gxOkjS67H
PCGKuWKY5eMfsn0fflmgtPgLXmZCtSOYCcvb7Hm4b4WYz/TVCqnEdI3g6Ykj
N6/ersY+udCIML0Jm+8xQYB2dzhC/cK81Ggi9fg8HR6SLERRNzxRx80W5A72
CcOQvyo8yCyobgVJ+15dxszp8xnpbC6q6v8+zBwo7GjyEuqxxrMWSUKiBGfv
Uf2n+cIRu2KyN3cakQWUG8M+qOSAqyyRkDDv86aM4eYYWHuE+L8omqGqWRRL
c77Tyo87UbqGTOvpETRyQX/fQUNGCCvpTq54ZU4tnj6MDk9R5iJSY0FaGhFI
eN7zsuhJvLVcwTqQdzAEDSf9giDls6fItbEMMUEZHmf3dBP7I9cZJ7vGmtJF
9YHLMxUXZpHiDmjj3xKmrXgyH0mNfyXLMZ7vMoV6YSRzhC++FWAI9aKt1dnO
JwM2bzWfmW4qHBcRFuTGjv+ThVrEk31Z5SJpJXPR4IhP7jsWUcCi1pNtnlyZ
4GsfQ9ZXGrq62rqYN0JsuTQuXKCEyV8nna0B9I9sETYszlXuDamDezXDzFM/
9uNX1AfpFoesAGe8OdAbO8DyzD7lglY0rSStmqXd2yqSpMQPeob3XIYVRJwA
dVc4nBsZ8+N11j4atTc1VEINLO/uZ4DUA8FXg5xSMhh7fIeijFVG/G4HqBU0
4yDGIfYxH5VBSnx6vx1GWdDT+gzjBqiDbOci/gnLBn5FiD3nC5Eqs32FWRq2
rO1+du6QZxcyx8qZyiY2lHvCEU5sjLX39TsWt2ixPwTM3OhHof/a75MCIKAX
YO5P6QWNck8A/wCbE0TWu1JTgA8KIZhRFvmCeI5sA9rroUDYpblSXvor+wSJ
YwoTvH3O4DLgPR7LXtB6zpqZm/fCkSQFrY3ZzfY+sHur9tdt7SPshxrMwVC4
K3b1QnmJGAJf6idv5HTartG7Jx1zORussNkgS41sRHkXwNFNShc5M6xHCqm8
YcsBBpO0eNCsr1tADxAZpHitrC28WphQkULu8b2RC5cW9w3LRAJxTypHD9mT
jN2LbkLr/rEzBnzgnxzFIUpg9WOIsDsEZlMfuShX/zUN9zJazzOmKoLKANjM
xhd0aSDygUpwOVZSmy4QrNgT9+y6Yry6sK/sMKxsmiSBtwa/c41VTUzD7xqj
LVg8e7i63GTXxsj2rqXLUANLhUs1DOIA8frSYrMnNinS3w/9pZzt/ni5cUBh
H3C/rWKh6GQxlbtUUeoeQu8P6ScGV8EXPIb3XDWQv5+/GtkcPlbDJr4rrQRb
dCWXuQRP0URsPCvlWX30Nw1w+R40pUPhOInxbud5jYTidnUWu2Aq5A7p82Iq
8Gt1WrSfwuXR5QOkFdBkdMWPMeDvhIzVAX3Fxqj/pKysfj1jIkg/SHzbGrJj
PVz9Bkd8H8aDevDia0o5NRy5h7l2wg6PGkcQvJhSXCPQXGyUOb9RjzC7g8Z6
qgIXYSieOrarnN8DGYoMCEd09HjORcd54+9a3o96tkTCFSvSGn+1a6G4wV5h
pdmV3OLWdi9i9R1FwLkJXVRJOuQBSFX4LQBaLKRt6Iqti3XvI5VkVGSz6NET
fLrgdbRElbuKyUVC9tvGyr65rgqgI4AmqklCtQ7UhTc/lfjt0nt4AKGixLrP
9BnAcDj1TEYjjdeFIQ6B/YlQ/CzlMoJAy6E2s2C+niTKm+hKa85aqS0uTpHD
Vl2QPG0o0KHvYbnq5MeZ6KKGolTr2PjcX1REWkYuVO5GlowYVlUTHkmtZAIL
2X/4Mv1Zm9i3IcQ+bNrabYP8T2ZoTQYLWtYN7fMdQnWVHwGgiND4s96fAKtD
atxifCDsHiPf3vFNWFbtk2pG1tgumVTiSOfabDCOfKjywZTb8nPA5uJZoUPN
z40tQmObLr8/TMuITsDGEJbZ+bsZaqgZhoHrLQ2nMsxmqvTAv5TpwwwB0sH7
ProRvYWR6L/yYfE2s7YUi67efIJ4jQppUVo0wk/6EIlfzd4TQFLVmHC7p/Ab
JXiGI1Pz/xGbHKDm7gty2YitzxyySBqZ1D/x3G1xc6tBZg1noOrk4k4G5X7f
dVP3EFqGqRAoV3Q9qYHzd4+9Mkny34CKT/fYiw7DuDXmBgx+UaDAKrVNWItc
quCqKhoA9mTJAuetmxU0GltbvbcNTrIRN1FzNteiJYGt8l81g6i3JmSWumzW
P2q1i8RQshlbUtdi6LpizcFSPatWAhymNoHa1LghiuQkXJM9lM8G1aNu+5/e
MQbaHGQV6dokaW99DMOFlBeF8rPcgDs3LSg29yKF8E+hFZkxMeK2r7540HhD
f2SUtc/Ted37dR7ekSMEpo8NakxruoKWaQsvyEHFzty0LOWFzi7/7vtV9P0/
4X4OidnFPLyA4c71bb3KLdaNEj729qTIGQsLR96tKJPnsE+e6QTU3OyPnkyn
pBmh6bixz3A3wP8/35gzqBDynfDO/AVBdj1o9wRvzw6gCB/+cxcn5BsT6oU6
qgOrhy693KucgRtWFFEYfokf2ES551oVlfj7v9MeUp0J6sO2hXcoRc+my9uf
ugJ8EGxuvZDi0fKkYSQ0zeo1Jgv4C0CTrRUZ+mRzX7pmbhcX63PLWIgVsqaa
nXA1nmI4EEwR9T/jk6QZcumVWpryw1+gleNv6BCdFeSboQiOr16rDObdGg8Y
J//iAoVAunFTPwXlsYTV1ETQ/+eU1RI1brGAxPprCFOA2LS2O5fbRQuS2ozp
2Lc60fxTNL2AI/+Vqtt1eDweTNG9r68eUkdx1otBb7T74t3KB4O6BevQWR3B
FmiCRsn6DB38SGAv+pjJVWOjfsWQ+3L4kPccDD/0FAIdCtpo64As/ectMnG/
Woyrw8V2TRJVWh5e/Kr3tU0QBMLTnXKoS3VTRiK7YdhLXpYDFbGIj7+eEOno
X7idV86wqaTT9uIho3mNETS3/6564M+tOdlGOSoksM/9aq9DVRntkBHNqzax
ZAKYGjJSPXkhY6+ocukmuLFVQeSnxUgCODsFNhJ6zK2sdIq+Jh8j3QZOeaGZ
boFdXiIfJeB5Pixo5wWnEzZ6I49+eYtKuLBinkotnBCbi+M/WPoRNhnsqt59
amVazJrq9RVRSZji8B5SzkuDxchVVEBJkzP2OXGPiGI3ala/7ktTM5feIWN8
Pk3LKIK3O4HuvgKaxZPIjqqL5qUlrdNNTzrrng6LXRAvUB1of3eAG4+ct29l
/TK2o5cUeEIPwArkRVL33n/WXUtKzgdUx5PxQcclAADL2tnRrLCwe6AA65gK
ugYjUqgsF5WLtuCOcYnlrspOJtxoQVPNuH8Gc1p1wlY5P6tNUJOMBbVgUy73
58ww6e2yJuHJu1GNACozHZXkELkovjt1Uy4tqYpoui+ZtP2cUlQUJIgvD8hY
zN1DKoNbcotiNj4r88vCOwpRVlBI3CqVc+kRbDLTcAF1MmDmDeFuOvQ0r0w6
iBTbf3SoFeIWruhPPIQxj+OIOdtCPnKvIlJnepNuChHJNkz3muVPll6zK91S
NgMDbWpdn1jiAxrtORrUSmSyZJozhAkyN1VwPUqI7+LZoiWmCdw8r3Gtp+Yv
e0IM05P4FgERqKbUCyipxise/0k7mzYuWbBQWCvfEy0rOajUItmGKhcBXA7u
pkJnSNeuNLBEi5ouThbgMiznjL5x79zyUlqP4gi2pXrDKV0jXEs1raBTjC1+
6zYvl+bkjmHpT8QPwJQTs3avjxUjMsyjCVv1ve1aD0IfvAXVuCie3t+G2CmV
7eF+R8DhfATELGy1YBKrH7sVIZ7boLURmhMBNnoH9gdHwqiFCDTgq8oBt6w6
mF6GfiXqUCMhgq6L+ZN+L2CglFuQg/ptd8qv8J92Iugi46Ro4LX4r1CB6sav
u5YYmhHbFYrCyj7a/lALF6n0yKz0CgjBokSxIh0IXa399b15lnwa2qWaixpp
dc+1PGgACMFSqTdIdGKvi9WsQQa4nMddOLdshxUNJ+lzqD/LjiFLktbxIM1O
XQWxZMnJIU5DirLs/RTA6EgKRfTmHazfrSvKJSKk4j5nD9YGWUDTH9AY0p1o
yMM8zBrqyP+dpdkY6pLMEz0mOIxRdZ+8CvGKbGY/Yt8Q6qv5nCObHkH8RZWh
UmtSk8IOWn4FWbYWDa8Xnqf62U6FvYb8BhR8MUzV0WWiKCTT8m0sbm/EVRLR
51eheTIJ9f+0fa0j7wt+fKn1FjvsGlL0RnvFGAbc9PQTZTAi7wTMOb+vN9sG
MMD+ItaQeiBrVIlLVrkmAlil06xQefo2lWvH5qXQF3JKLPZJ69fORKBLpWOy
JWDLo2mhpesi1J3d11S4LPom84kjNuRWHE+rFrf3rYuoS3YDM5Lz2pBijBX+
0e8bRrZFSdbTaFZYioAfkKR2tcWyK0INn+DPHxLV5+GkYGmH+01l7OJgl2VM
DB3IEfgLG06+9Bhqxxt9sFdxNFU8gGLX2JEMmRqOnriK/Ug0vv2zcF/Z11FF
UONozV1vwZWDDRW1FnsCiCDw9lQbqoZifzCwf+by2i57sqS6amlS51c5RWuj
B3vg6GUahnErsx5KL/RXxC9Z+CG5fky8KJCNDlR2zG2tsb8Rljtbr1isqUai
H2kE6K2BShuv5WqZEUZIe/QEnT9A9YHKiR0gRpdrKEs0cudSl7/+vs94cWC2
pTkn4BTpOJsXJ0Nqq0wZ1ROTCAe4QgL+ucC4CR64oofSPfueJUIGLoFTXSpI
frlJmil3c71AXS7u6AexJYTII3vV9YLAY8+kFYmm3FQS2EwPDlFLj2DSTk8J
7xsrixmoDTiPkR2g2TgpZWaUO4VVhsj9jZndzLyWVO/Lug7VMfv8YNfNpNjw
enAdE/oCuew7QRn0S2Xdy9opgA5iAoSxDVb5uvUP3zGhyWi0ilbJ70J+EAIM
KHDlft0WN4DfFs43vSKHCNN2FhKBLuXLdtl/0MM+IevyvqPy+AhtM1zrsM7S
xyiZLpkBF+FWDfC0evPtY9RMa83041n9ZB6SRwJSHz1Mqq/ikMew0GWJEaI/
h4M8nGjI9dOTXIz/SXKbpw6L6vhtkT+Xx2Jk0VXBZARAc4B3l8tF9FrKXSLF
3fYgFBk4SxRqnNajLychkhB/b07hKJvFMu+FkAGzX9B3m90F3yb49HPaUN2E
1hkJ4xUVErQ+WauJiwTajrZwEjGdRkDI/VirNJiY8w6TVRIbsfeRVvogBsYW
gBiEo0QiTL8Nczrlg6fHGsFd8ld8Dva22UaYHvn9pgHbbbGDzr41HauStBSn
WKW7HG+NN9ZGRsqNejwdYCyXpvjWAvlEiDYg5yrIPx4mm//NjmiCtlH8I+CO
OQoobpTb3hx0b/TrGU6h5kodQXfmQE+nZFSvFclQalSlZpOh+hHWpEDA+O+O
fNg7tRANTghH38694enibLrrO6B7IpIPnPDp/DDNSm/4PTFTAeFHaD7w4kAa
gL+1Kxc40Rj22eHwV0gJT9wQFQL8dv9PIaCgROVkoB3SCZM2z+nn1kmtnWVY
FFmUmRG3R5Mj1OXwUfh3NYHyE8ZrTU3Ag/45CiFhUMxtRzCtsoV7dTI60JrH
cQhm432ed8aGjFH17/uwDNogEp0z9IhP4SjkEASpuWUDxSkt5Lfg8SENWIGq
bgjgz8Sb57FlOI3u2eXK2ToAR35V1uZb8xMgQeMZRTOBZf2SkWOmKcWJS+Cw
F05+FW/b56j3SjO6sJ2xSg2SSndTfMgaoFehEYvemsPvcpemBCEm55Swv9Dn
hFElPQ3+2wZ2/2eHzt8dfB8UI57XmOCWqWYKSE1ioyrd2tkbbSFad2uSd+4c
w2BYVNHHTv0X5/jZqVtoFbX2LrUeyj5kDXCLCACncd4C8Gij5BgEHiBKZcQZ
RW62NWdcgH9aqs4IQgp6ZlVWkh+lRhCvDT0sIPnH4DKrITjSBcOlj+szs3f3
R2Qv/iB9SG+JFA5dRpy25qPeNRtURJ7ypd2AqKha7b6Jd1PBvoYH9ZXw1bi7
B2F24SGvdexNd3gKPwOvxd3r+JNyf2Wmwz5iTI1ccmWN+Vf0UmU8l9rLlqRe
x05F2GJQrXe/TDnzMtlwBHZFU1GatcSw5bbeFbXSgb20dnOGyVS1NHJucatL
rlSAJnopZSBj/zNH6jvG1V+tnZr+hbM9rtyVdQAWldsnKog07x7XkErcyy+T
1WdtnRx5YS2tJ0X+PrD/otjCJthFrmzcNZDgR/K5D6ssewczFwuHpcUDMGPV
WtRYi7nenFQkpc6Pao65GY9lAusLRIhEE4agh5cJ2QFWTW8PbxgU4bRsdY78
8Xpa728PdO8A7hjYXvze94o++JnS/H5hyeyCTiuWoj6gB5IRjYsZWRrlT0Fr
sVQTpbuaWhg4es7SEsJO95Ye6YUBVo3UfHSObtgrbgxdJNKMaCpscEEFNJ4T
KOEhwSIM2lxmJATlG6F6o+iTcoZSjGhqmlWw77zEoIIH6q5eWuCXaLE912xA
T90FuMkG5L0b7jhh3JPleHm2wi72wr8IrKeA6ZIxGleEEtQg9FqUbOWi0OS9
nibJxbxUhDGcjhAYNwS8PdjYfY5TaoWEowylhInbryHIJaNkA+ji6rl7zdU5
7S05qyfNwxGIjYObwvP0NE7fWNUAeiiM/ZKXvb7AbO+0MN5z0N7//wGQA6HQ
zlgQhnQsTeP38N+W/nuLXB8YlYJtkVJPX+aZsEFWvbK7EfcgkMT8AB1vb9MS
niPHehvRHxlLzIzqbw+gZAc6xvvBVHlcY1NA+BtKUWFy6Z18D02ZptTm5P/1
rAEZgmxe7CejRmzkRLLz32Irx3abwkR7GgY5dn9P1c8AF25z6f6+YVRlRLod
DzUoam7R67wPBHtJ/HRlV0kkqsIKNc8X1WkssXZH8SELl2rNXMAiwEZBEw5x
yV1EFg+fq3gtPEXJxCTd5LeAaNlYQp5yCR2F+33GzeledwI0AgP5WhhtGg/Q
netE0MzDNGqpMa6foV8ueRChgaY20eWHtzSpFDf73/4vU5ayX33gtaZnGvjH
A8/Ee0XG3mKYSTUeRQCEBJUhXfyAROm0ta21OfyroK7xfiWpsoCgl0kuTSEu
9DW77xFqG+XmjYzUei82/QDRr5GxESpxXTfZRPrbA+rPuQdN8u/RvBEfWY7D
hpAvShfwnCdgv6BqyC2ronlAX98R45wVLq9i6csEOsa3zIzWN1TSsyYEDrau
6dzQOnoLzcT4btWUZQDSfP0XgyVH27xO+s1uLbHa6eXKC/JfdXI4ZhF0lUf/
2Ox8PvFXNIeDWBhuMU38iKcWtf4+eZi2rYeCkNwsYWwRKYZnIgnSRDCvk28n
xaUTJaOUs9uN5FiSE+oRKDO1p/mHXv7XL57tEqSshGlNI9Uo/qlhIJhPPiEz
F/zOBjVdsL7iMpmuBhHkKvNHTAywUyoYxKnwZHtqPjsTXmM9JTBUCn3Ef8J5
8qszDyjqyZ5HJmjGlEQCeUAXNaKlnzvg91r7NW4tSB6ZxEeRXD0jOWQ4NuIm
jktvHcI47bkOI+N9fINJ7uzpUPert17a8GcPQWhvBJcWtyaAU5pailCZvC2o
2uifZNC83vQOUK5yABs7LKljQ7k1lwJfzdv3cxPWhqsop3Jul2K0f5ZqTV5U
uAx7iKJxh6PTRR0jSGFBu0w8kczS4Hmf8p7JKw1d3X4y8WleH3M/IU0JsxoO
Wz2pP4HTCqOhLXz1kDMeBhR3Bx9MMWQhCHJCoC+4Zf26EPSKmCvzSnYv1Ztv
tRDhao25F8BzBKMCvsc/MKOlFrwkpOkqKIKcMRKe10ktBguSWIbyy8raEuvq
xqgD8SXB29XoQjIipmDD+MPxvuwKwLXg2KJkJeM3K9tSuWy666giLynJzZaC
WTngWH0plPSqjmAc/4c5D+Yu5pSIz4OQ8hCe+BzW4rJ45yiJ5yopUL9Y+qtF
SpHujE6TgSbCetj6//MshRE2HwBnKglpnJzf8ZvnQaeNqg93V53FdyJwN7Qs
JCuLfDepSNmYAMKMCjw7M7o96kcpVUDrT+cVlNLhcbrl7K2U5lZ4N1d6Aytu
5DOtr5D806DnM98b5iAziDIHT9JU/VuziLvuA443mOIRWUtOaOcXWq/ytPQ8
UOV6vCJO+SAIZq/Qf7PpEd4etjwuK6eq0ibjZojHn227Ecy4lqu3RNOTstfT
CvTgHuBQ3wt1r6Bh+Fje8BgqaJKXasfVN+ufT0ORxkX4y2zwBE/ycJsH+BVH
XxFOXiCHiIqrOh+gj3VtzCvRSlZKH2cCgdFts24ZLdr+l6IkiGlBEN8fLxxV
Y+0Z29cYBMN+gcnaB34Set4eLcy6inWJ4O1ohkSVj4hV2lJWBYcV414X/j8V
sezbQFeBEnIDYrnIcmU+TIYwKslA0YxzcD8b8T3KrA8bHS0BJfyd2UuBrjvb
5AF7yWvCmdnMsqeYXhou42k9M13cgDt7DCYvdwmasBjQHp4MK+T3MbfeJm6i
VhP1KCugsxoXgYQHn1M+/LZHIs44c+79lflwsCn6aJ3rJ29gDIfKlFdZwVxV
9uNeVMHIZKK3dLwFZg+7Mu/wXnRYyRq+MgPiWxG0HLM8o1/Owmuh8Vkrra6m
4UgBCbYHGgliIKvuT54Zc4rRdRvt0l5cT0g6qLo277fEtpj3SCwaMLqIK3iC
gIeM6edlaSUBG2XXYv+1NBabAKHOLdA99INIIFz0yehf4sAw+DuEMhETSQCG
tUQHJjZQrNMueuRBjJPsBN9UygY6xUhmOzMdKZYGcCRmRDjQAIe/U+A5MbzN
4T5IaShTVAqsV4Ai46wKWcONWeLKGq2tOcTYLYpIcRv9d4KbHTEY+Mbr20WR
H9pYQJqM4R6McgCEznr1eUUUg5VS0sdSojXVG4WxEfEq1zIe3AHZurUTxKRO
ooGyaAQLeex/I5RItu8eYd+GRz2WvpbO3j1P8DD54EkoAP7iWaKnacs08Ncp
3QxO7P/EQvvnUif6/PhQ1CQs9Hjw36yWBCk8Wfn/EXwJxxbsiMo8TssWTUgt
g8PxiwVHG9nHHyUwBUHn3j2yPtLPBA4B3wRCWJ5YfcNlPDgaD0+s1c0qJM7J
P5u7KMlJYgy7r2RFns2+dLa9N2IimYLqCFrLGTnMdOk1F/s7T0RKHbNcUz8W
gK5VdsY/2UDXS2WmElA9ojewC08qasQ2aWs3MyiVHtkJnZqiieWOPXDY1pLj
1raQIw+r+tcKqBhrIvY5YiT8gz/aL5aqf6qEBR6msUnhVEv5gk7cxUDf7S8/
ecTtB4o6eKJ3+ZOGUJpDB+dSu0yBEw937RQrikJay3fzX9Xh45ZlYBfSWy8F
0Sk0/mk0PRYOJXFCuno6XVWfHiVlk7GjSsbh1z/f3gfjPRNqRhvXFzyrBT/Z
hrkcxhyaWyUrN94t9pqB7WSt0u+AStBwo7nFnPB/Y2wgnDSYTbkfZlplES1D
grP6GnjSWalFwyVnVbbWksZKSy5+XCR38b+hZNASCuNf9D+58NIRIQMj2Y6n
QGhqSgT5F7Z755NhWaHGydqidBMkfeVhibWOpNsGfshxGkTxCPvSc7Btt5Q/
vnNdd9gY/NYCPNyhS/Em4qV0M68UOwuu0VTjjHzNcHCPivZDQCLcMjTJMxKZ
4hgCwNsx5/N5Hg+T2z2Hq+JgE+CvisU+zxZ0Q+cXopsv4BXwr7gDjr8a27fj
xJsjRagG2CKTT4FWN9N85RVbvhcCWO6FCeXC5BkDNBTwcLt5Nd2wwKi0wc/U
JMnjp9soq9TOSHHNJT+DRJ0Ub7bZbJkRXoqQsKTBuF4NCfZK6AQ5M8hB7leZ
y1yrQq4L4pTWk1S10JFwW/lQ2CmA5OZ8WLMvTVnpzvEqKoiEJzoRYeUHbu06
L6AYBEycHVVvkm3p9aab9bsFsxxCMnXFO2fP0cDwyt+hmTh1bAbx0g5tGwnt
xZKkFZoJLKS9srISdlk1erQEvRZTXzWYl7Fsbhcb9LFD3otPwUKFos1GIqn/
+TaYWz82NSowrJKX8Jb7BaL67/byQw5ULwDb3ACn3bDFIE06ry+Ic2oLNVPk
uu7nkq/x5b4rQuqoN66psLTDSWJJ1oA8BjR9EgdKbRWEvPquz+6CYmJoLaV5
QET8Gct/WLMoKiLPfafnUNVKTraJo3xxCKYjXqGuFUv4PP5Xk9BQYWEUYP9X
YvB8seA82PLxsvxu8WnifU0kuui9o581/gdfx2jwHD8zO+E0FZ72iTybm5ux
SzNuZ6eMzVWVx6x1zd1bn7EG4Wlwew6T83p2TnutDc/kzXm+reWZmwbhgKxt
Lnn6aj1nUT/BRtpTdY2RHDvMKC9P6OjOkOvifVMHJy8P4vyEQjI3RZDn9XQN
BXg3LvXww99yPcWLnHgBGf0ckFn+mXKpGtggWZkxcZuVBappc3sU9dtZfgnz
g0Iue5jZ5wJ+r1DLux3c0aWTwor8WHkTOBiGXLQ+7aKQ1IajuXfvdl0SZmQA
+YSElDYI3AvA7gC/9WA+SVEZfdZvFo2PChbHvDkieXF/RPgZeOlNFJSSIO/4
/srgTQCV1huGK7U46EAEy1P4Oalo508VDjWKC3lC3qYQRe4sxzgOnwbFiVW2
nDndgDd6hE9+/l/XX1bmjf0Wa7jZnEd0AT+rDO89qWumGYCKkqg6gKLO7WSe
AG/mWX0A8gLbXIN6zIMVED76vS5SKOGs7KNpCRrGUYxZVppql05+6xrLG3/D
wO2bBBK/xtSJAbxCfqVYUJ4RDq0XT/+likZdL4/n0JaND9ehWYW8AZOXzCf5
W5WlXxCZe8WSkMn8PC69Tn9N6tnWHe9wvqaorJiYaJ+VbS4UtH3RIUumI0S7
cFtBK1a94A691R95Y0eDQ51jgXEDvbAvxJ674NEQLODTEts99hdkexomAfMI
XnSoMeFTdn13b+WXENnDd9upLIrRn0BF8n/AWtP8FHAB9Ohl9AAK68XTB0y0
uz+IhQtQ6Ot2hpeBsEezebDzcgiH0jLyCqrSg4cR+u17QA/S+oDNSediR1TL
Zy4fjFLklY6lC1TySX/CH1XCo87r6OpoJ6SrbArfAtOqA+QqKQgUveSO1JeS
T3WJNC7calBqnmQhKRGytggX+CJySob8j+SHtuC2zaU5HZ7RdcpFBt9CSc7u
MNXKhlkTJnOrwSN2huiGYrOTUH0LL4pc9wix4KTk0JWwYov7XyXsvBG/h8iQ
P6inpDmYh557dUjJtzl+9lPP0ID6BONw8pDGykf5IJrIIjjs+TuoSFQrqRWv
MoP76FkuX42HTBSHn+wdB1Y/wb3iEUmiE9lhXCB2WdZg2bY+quXGUceSbjxe
fPp650u7dTn6noqSXj5S3L0RWGxlo0RV+y8WS60o80UPsA7C9FI9yr0R42SN
Xq12iBZna13ukYWp46YCBv+WDR97RBvrhT+r8zsyfLXgPQavgcXeS5eFaRIV
tRqzoglcCZ2vKLwnp6rHmsE7d5cfZdIu2CayKf0iN13q9qnzBvHSkGeSsE7j
1neAO3DDexpiigqJLhe3Bi9td9iT15LDQgb8r898Pmlalt/qELm54UYdKHUw
f2TE/gHyphDYBP3z2wM6vj9gM0J9A9kXHwbAZbGfeeTqtWv1uSD/4D+6unsY
jy9YK6DBbYLYCrORLQvaqqR+fqeefuf0EhBn/TgS2Q5zzFJ+ScmjxRtKT0kE
qAwyj/ZHR5euCMCtYkWVourezZrolLDxnOmDk2OFJt3TPZze28Qh0w7lXsLg
+PRwnYzGYlwV2A6qGjZipKWvoufAvpWNvsoQZpuXcvEGJYwOvIIG92IdTe61
dsMbaInwUK1GOjEp7nFDTIRP0Pgw1f32/oOwV4f/hH1wZ1/a6GjirFk7J46o
hET0UEtt0wsnthTl6UMs2pBouPQKYmPtg9TJ+AqRv9nsmr31tOZtHaYkXb59
YgaRtKRGDo0ldizJnOgocbswwW2m3fKxV2FbfJ6VkYnbFJXDmVwXVNT//s3u
7988ueuSH0q8a2oSHYHpFiPyrgqgnw8rdyhv8XTtdmqaP40p6nq8RLyigYap
GnyGb88HxRTQc47pHbcQruEu6SiDv8E7EYoWTOhILoOCb3iqB84YAPH+TNpd
yTWFEiHxTkxuJs/WLChQ+DXcdHUrOJbKz/cXVeX6Vt6iOZMO4JFZoA66kLOQ
zl3puVe2OFYoG/0kxZ+owG9IvuFjHiY7qja3yiWrT9U6OFI/RPk1uZ0g1XOR
Hx9BkHSCB+QZNQQaWSi36iMw/LjkVR7LEH071iPNwZ2P/pB6vaiNgmahHhh1
ULiHGkg7lvwxmGzscr/fWWZlnZi1EsRHWGIOAmhlAlfa5IxU1Be0IAbUZLwu
ISytp+rNqx5/hHcdUj5onChmx5Z4LxxMVdPYsMmvEk8WW6se2ThnQiovelsw
MjgYMGi6qmldKHSUtuqNMjfj5aBZWqKzSfalysS2jY8FK/RHF8hN/WdyKwlD
Mk/jPPhGxHlmZqk4NWshLYb8vI3++eZL9Bg0jYboGOSELIwpdJbfaGtDaQI/
8UjyDFSTs8e2FY/ALqqgVP0Uw907ZklqgmhQKLb17M1ddhkty3F6kfJzKEXt
jfIqG+KILH/Tu5B7sedtv50L5l5+LvEwE8vpE/+GswLXLxQ5qNPUQqWRsXng
gVXmUorj3DPLKnMg/PHjIB6nlOCIDBjC/TrW/Q184yb2Lnf3mCEHdkQ0tRCQ
O5ouL3XmSWkN4de6kDug9qi/J3btW3uei/uDU8HNHTlbGftckx4obDiaYTEU
ize4XoAeOEb0XEx7L4WIwVxx+TmWOBA83a8vsIubUWUDx3uB4p6kp228z+ij
escFv5RkdumpFx+jsQEtardBxM9F7/Em42JVZ+ziAO0x/rLGEuErnHFV2f2x
CFKsYISFR2P0bmGuQVT7QYhUPlgVLOLcHLZ1sl+tdnhuGzoO4VbQgdTOp1aK
p4H8/KhgQ9kLE137LKlC7ckLvYsFVEm6aoVOMD0JggpSljKC9vwCKy/ujS/l
55z+H2GIpI0A2XyRU2wZdKG/BUyksLgzd+CsJD4Kc8ZltKGXp7SE36FvYmrJ
v5suVskW0YeJ2viCgVv3C1BVjzJJGj6LdFxgzOVyR/ZbyyBuBDNcXrSkirDd
aZVCueykct/dEF0RDzsNoOGzZdR4baBJRqOPE7TWAx9vwEQHQUph9FbLD4lm
8cEXT7GJgfzlo068/k7psqQTRaPG4RX65ZPpqj2AadLDCqu9QSOl2k/1gGL7
xpvqESbnd7YAhf2gEo56DJ1z6OgZa3uR9eJwQlIFNcmH1JdP9BIPUnOLd9uE
3ZHIN+RJh3NrjSBbkbybFatJ2C+XyKSRnf90lvtohix7PIV8f9EvyugCk9pZ
0op/rwyFETJ/H27nohKuK1AdhhKPp8He+EUZDt5D/bLPCxfyGAR24fPSnCur
tZXKP2pDXaggO6Qp4plSYK1RPNpdZxEa+ttoSPZVxga5pw6keok+geT1zuU1
KP/ddHroSdI4Zn+QbRNHAtqp+RFJ9KsUc0FIbkd3uL4oemdIBJBXAWamllXe
FyHRCdO7s/3K7dpPNfyBqo8oK6SPqzydOUD5l0GP6cpS2XYSKgKfpfZzbH7A
Ni+xzjenD6W4dJr1cqUMCKoowv4dppatyBXCke02vSEr+3XPriLIEjCAVzMv
CWgJCp9P7pi7/OAFAqdP2Oz7ZsxUEJAblhcWoSlhu7D9m5jZj/Vi5jY9d0o2
v16o68a3q4cqNIC5wiyfejGq2cuj4BSb4ts/t9zM1qlAnnnVgjPlTYFF+c4r
mRq1Oen/93gQO2XiEf8v9PiZoO/RyL6RCi3s1gQcijNMacZnIL2mI65ojnzE
GUiIPHulTc4IocD5FyPhCHogPr4PAGx985PkgzY4sf2KXgI2WVhVOoJ118dZ
LZtTEAlndF1p3WexAwKoHVYu2aYp0nHjIan5KRvmTNGGbY8Kc+eZ4+4Sbe+V
vb60dPq0hMV4A0MYrUFtFeHnYH4xuqoALmiwZHIRbEfSTtDLH53kcYb/qxDf
ktF6mABIktmyl4E88/JvK61bcXn3/0Y2IlDd+ReMSUI0h1mdN9ig3CYErMt+
+sAjkv+OTy5ZR7coIeZN1fq/FECZx99OGDKI8sRzKykaCI14vmTFljlJWTLB
ChGCWyKtSM0lqrYXoy103pS7v/xaNEkM9ZbqmRYFJdOJwhHPT/34bZdxay9q
zUrwh+AqMZW+5JukUKk77FZu+dk7fNygLLIaNZSlUOEc2v8vxpc1forO2wIc
ivvuvegbMxKunXW3UuUYVwWwCaN0ynfpBnPko7YVt3B105Cy5rxGYsL4XDQ6
+HMsZ9xDIe4sT+48/2rTqURD3hUMVxDvG/QRY3HFJzRBTDc5bcvqqeT2u9L/
TkVvyLIILFQ3MqMupkwqjRTfEeuKxkwA7e7CS4YAdo0oxUonEjhwk5tYCP5i
Oyk7Cl+RzYTiNdyyk5fB9ojaHjIH7CA+rxaEz0xg7CCZNYzY+Ac+B6DaADlg
R/haXddrP9OzdjpCjuFSVKDBHFw8jx66cSc+0kVZ82eoU0Y+9slwoW0pcKgu
3t3h8j3F3IRXaxwej34UJEhTUYiUIMow2qVQTM+XscdCw3FFjLYyWg65wxlF
FYs3i4ueBpyYio14T2xlp45eSt1Sy9t18itb/kW+/a92JKk83+Gy/F2qahV/
FkZV5vUj1X8rj8VpTxOdO/egVp2oeqcwgVziB4XBarkTxa7hNBRoLp1KsM/Z
6yulNC06pPZhI7JFfnoJXsiYHe8z+AVo08Jhn13EpusZaRbe9BBdcJdSrXN+
gPukJ1OYWgBNMAFwYvzlM5oU6NCvolwgwFbSp/J6mNkMfXbMyCoEXj3TBLjy
vMwJbHcWPTFGeI+7etqPJMCd6QTPLqYDeQciyGI4uVJjib1YNmF6r9BC2PAz
wJNx3g9zt1eXASRkVPL/jvEKwg0VJ2HWg3nsD7uAaT0l9T+LJnz2+2RE5ITz
Ilq1k4V76KOoYfcJkJRFK8HHPfHnU3LZHq5kEan6yPahkssGX7sSeJTadLit
ofsARFV9ZZY9Q3hXnykEVPIbxZ8aDKv2CD/cfoII5o2V5NWwQhdMENRrccnt
byQM3asy/0tmV20+QWx2/Pr23sXY1qKkq3RSwefhNICcG4iGZPYGV29QD1PI
TCtw1YJPjze4nu/2XAqdm5tlP6xHNS6j62yxJwbWQXkNBu9plmpzKeva0q9x
3AWDrW5ZVJdaKIoQAne+oi7kyryaVpaGqCFfR18wpplYBswEx7Jt/hd8f9gV
q/XdLqw/svjJESfb2xyRcVWikz7q0qPh4UWRq2GF+5T6zze8dPnVP/Q4JR/S
JYIsWm9+qnUDbv7iO3y+khNFj9aGbZrgCCG2749Aq+DGJXrg1EeS/lIC8ExU
hu2WIkA74VpXxBMkPEOg0+zqVUe3E8naYmn8MI1minZ75lx48H4m6Nusal9H
o9hzqLAZS1cQ2n51lPmLP9aYm8a2IV9FKf6HPbnNswrABicLbrZxA24ShLim
km+0yySdpTnhP+6FVbAoXVaBeyOdQomRHpnz150fOx1V4nbPBXQr8ZMPOMsG
ValU5DRHhM1S+d0T6It+N+f3DHjieey+96EeaCEillDEpCSFqsdnvEfCo/RH
oaPLAXvoW00+rds1buFmit2F2R3+WP685OSgYK8dlov9w+bdcx9eaWkKU76Q
a+fk4XLLpWgwXPHYdWbC8oXQxmnKJSyYgdhxdL7f+gn9IJuwEmSML08nSxG5
V1OaOpMNxW6FYOFXwMWxm2MJHlQ2EdkI+qjk1Oe9fSlpwXYEzj1MWTr4wmh3
/C6R3cShVKcLQMq7QOtsi4575t9mGCuSWbt4x3Qnt3ImjJ7bp9FMfGLmpxFj
DOpzxxxNnsU8OjSjrgLrLda3ZACEnU/F2ggZIqAmBNATMFfmvHWm1Apwxurj
luq0sJ3h2zAS7NzR3c08A2lk3IagAYKqy74sQHcwNL9nhRdp+TfHQf30a+/4
uSIIdkCfiHaMYe1p99g6+fuomqo7m3Z1x2tUdgMHHmJOWSkk4bsSq5oVtSYc
EmKw0dxpINnL8I9JjJbQihX+0WUFWVFDTJYLY3p3iwmn1d3JDVUH01GoFgy4
Vnu9rv6X4A64zwYKqpYFooDFD6ylXnY2yx7PXvcUKAQeXDWlVRhENKbBSNqa
X+3mJ3UKvtG/vwCy/ggDHoVwnWTvxBWNGVE5tQYxb1C4dd94/MXUdQKQSGQ3
1Y5SWRyJ3U+lYmdnVdhjPfFYtuI7A9MXptsvjuhnbwk7MTp0+dUK7ERfgrVY
wEuqtp8XnkvdPQF17F2opt4bBIWAhInguajE6JyizufIzuR0RunlO4lc4zfY
XY/s/6iNj0HduIh78i5uH8nw3CjyaEQwB4ZjQwU+HbzC8tQqywhj7FMrly67
0DZKc9zpJGP2iAHsZ8p5fN060WkBw+7/dobJDNYwYygTyI98N+rtW66Pouhc
4MXtReKM12RWhWIodSxqmjqgZDJ08m6aI0JfkHmdIKqmaRolLAgNlNvK5p0e
yhCJbCStjwWYGvSFzwBCTRdl/kQUac6NiOntDjL/z8QJsgLbPdaItpn7oNLU
a9Jvxx8Ociq60WiKtDrpVGDyuMPDjMRvr6HkiuoTXvFhs//OSPo8yTp7p9nQ
Zbp5TxbhDAvI5gOIXjLbaMKnSZvaPlKH/6+R6TDhkTN1s28rsCqZnla/ka7m
BeZzzpjjhTxTUNRn9CP2c/NX6iVnP5nMRFdi7BbsCwlmpfpxeU+C/0gBQtHn
QOWvhHRYE0k53hb+44e3y0r+Uj5YqAWOOUkd5y81byTaTSV5QNs0ufmUNAJG
U07D7ZBkii4JIkpE6PGLdoZ7YIysTHHB8uFSazHUqs92maD7VNA25Sq9XtCC
lmjDsyAAdjy2WxDwNsZ+totrcPW3PBy69AtjDMLjtPhJ48+50jT5Hg+ai479
T5dO1QyywFjy2U2bW5jhKU/O4/HRIGno42eIrK6mG3EyEL4aWDpAEVKifSKk
FdpZgdUdh7/9X2nr3KgfR1Cz2f9gcFL4tohNeNdYrE4lFAVCSsVfY5zKJowE
ocfB+f8HnTdbFFGJvYtjykAQdHhVb7FY6oaEu22SebkTcff3Yx7eKYReyhlN
TeYmxrXnBwSTxSfQldAA0MtLutkkAdZLURwulpMT9/spn52YO2B/7JJ++ATA
4xdJO2F2lzULzl4xlrYlxzJpOzSogzup6oHGEvrlbjcVA5lxNdlQwUS29ieP
8lybTbtonNKc0vNkDLpglWCjulyHIJePk/xV43iR5ZLAT1kehahzoO2XOLHC
WRSdpoIJv8jre0zBx3HhxJyo2deG8QseWQPoGG6ffANLqQtMw5J+mso2ro9C
BTVU0D7YGlAYwVkDkNPjIbO8enRPNoCngIbpMUfmE8cC1YmWucx9wt3nfPC8
szyZ/rFSUio3pa7BfHTKtchddmcO4P8T15pMm77lhbmRcbhjv9G8f3VyYiYn
hC+/0AOP4bY8UXX+KCCWxnXlZH+4GPGFBvji+U5DN2w2aZPFMQw7QmfGMDwF
XnV4hj9fiW3Q5jSMsobBWnmW6k6B7U1//HteF4obaXGdh9bdYCWBcy/3jotS
JZGx97SGHB3ZDfePqTqvTOiq+nntuIFiIwCtg/LyVjvsUXfvf2KQPNC3EwQ9
Y/qE7jim9ftNC1863DH9RBAUeDI8B77qwBUHW7FhYywAEcYtMNPBuwuEiHP0
kYOtyA/12jWEqyiEFFT54bI7z11ApMRVuc9FSr4QI6Nf8ZXnZad21aBcLKwV
QKefytRCLWX+d8M3mkVzcEK6pjFSbzYWc4HHYWC/ppYv5DxYmfm7BYiKjmgt
6BA5FgH0oOJWenuQZpB/tPy5VWgl9BsIMLCVhWMnMWFWjzUNEFe78CNSY0fV
8fr2P+Mo3tjXC0x/5aOJgoVy2xQYKjpfgFf2aLNjoIfUFRYs1cF0oPG5c9Lk
84BtvxJjqiC7udxijOdFIm/nDVKfLcevOwYPbS9aOAsvCFuF/sR4Sws11uoP
s8V71xwn+r/4avMBTuN7rgdHvEd3Jj1njdQcBCbeJfWt2xOgVySpO0FwTTPx
8YEPaRKsPGhfCcMzPiBENGC0ja4wkEifyPCD5ejJKF6JQG4aQNA5P55XZ1Q9
5JL71NmEs0JEVCa68bVj48MiyDakheVVJFgm1dviQGxQEOMZ8Tbz+Lmuomq7
bVk9/klFrzuBh1uiqCFn5xE55aHLOxj6mFLw63pb1fWnaswMKhjH+/CJn7cd
iii+TmI3Ff20TKypCRotO7wT99PcE+CP4QcAEpJzGJ4u/6CXMu90HB+AUdph
2SEACa04L2OIQqhjqt5gm2Y2qKA3sy8FaRTf+oF118XgU8425C49+t11Pwjh
e2e6C5GKc1YUoAPaY9gg89/AshNvDpjro6DkwIQAcgBlCSKSUXDJhEkh64On
TjQbki/AhKJcsRzmpe9Xi6U9pt/X5w/m/6WT05k+8HTy/JcmJVHQVWLv1OnC
i10Og/DWQIV6dt63rdDGIw8zydSc7D0PATA6oN19Pw2aemXkESAzQSuEA9iC
qdz3c7mMsLZR3YdTtysp+sKbTdd7ucZS68eZek8aJ70DjvKfvLMuhgCfAi2X
WQKfLnPmqLENCFBj0D1r4yEJ9LcYMZ/0lKzpGYkYf2Dwwib2dYSBfNrHNOIi
akGvyuarHoW4v9LFGg1LFE0B/GvbyWHzwpue6grgIWw3VERTfmgGs8T+eN3q
+VG6F49iP075TMvBUELrOhtTOxM32mn5NZX+5MXXprd1/ID54OPLy0UdXnz5
M1X7syk+1IlciJxjDLPHQYf/FG7PGnYeP1LAbcj+c7go5V4OalZEh9heBFXd
lNJlQ8yha80hxB2MecCha13UWhCp1Ef+B5OvgTHC2h0ljcG08AVyrQoIyc/k
NL721CpKGaXYumbXw2A7F7qGpOtfVsw2asDMUHKTMLSxcSzB9WIkLTz8MRpj
zf5SK8ejW71Z027d/ZAvHv3w4mHjF0bGBRMG2DzkHmvWu68Pg3p0v06ryptT
sDbYdgSVUG552HpEgd7e56ftR5ZjdNCQDiuZY+9o7j3MEL3f2RL9z+yjLP8o
4BWvD9DtnmpvEvxAwYNr/0ZVOd0sO5KJvrxRg2MfvKmGYRVa2uzRnlAI1Pbw
EClsnRxndzUlWeO5SQ31xzJ3/kW7YD6iu1/kW4CS2PNU4dfE2x38G+xhBEQF
DsBTB5D2pOY1L4zNMWnoqj75KYOtmLiSCjaGNveXPgmrURbtC4tooQss90oB
VR04tj4ley30BhaHHmxmKiVP+Obt0HTkjYndnR0/21RYJNqqDh42eZ59WxMD
cC/vJh5pKH4ueE4aHj2qG4J++G2or1xz5aFigE80veGvlHogwU8qdxYvc7aN
sT92ECQTM6Ws4VdVE2tl77qhwkENFdTc/aTr51FvnUjpCP3X5YDHkBRHkRGn
wyGR+eTOs1E8R4kyC4oxDCabp4+hEwbJqn9S23uMeRLR5Gzdmc6Ah11j4pNC
LEL8Ut0d4Ph/E6KLkuXGB0zxvFkrLIU2DXKH3nNHeka1s5NKhF77XnSYZnY5
fgUtKsyzJVgO6WUpNUo+MUSYJUZ8iN10cg0J1lQLd+M1LafrWt1zPnaWUCij
EPMYhMekpmJR/WomXXT91evunxhDVtalvTaGOWWzKRaJ/v1JQeh5pPdaWcxX
YgsLeoWxeTVW1XYnwaVzMMFnK2+yp3Uhk4jbroqUgt4GFR1Zs90PkEzwpneH
hgPQ56dqj3YOay/jmjOOST6fyTxwVaCKe5G4+wr2lwjtJBZ4k0Dp9tsw6wmI
BuKDB5tCPOpwGCLdEEUgo2iC/2zVtRX8uQ/5DH2Dzb9eukUAk6QyoFk4CcGV
RuwPBxOWs4PKbyYAPn17nd1bts52o4r5bM6gR6JhGaSgT483DvLyq4Q3pkCe
vTl46DQfcQDacvdOdFNSkqLbr1dNoCBbbkZyQTk0+PB+Wvog75oJX1FPaXuO
1Hcm+Xh9K7yGSGnQlNz+ybuHT9BAsjlz7f2SQgO21rtQwHq+isDK4s5wvI2k
5hjcFhJZLCaegGzppjEAQVDXIOtWGC2u1MpfmAuW6vvIBYWQVUKnMdGTROla
vWMt5jyjUWDWsdDPVZnGqjlsYuYeZbAZyghjVrMPfFUYDXS9DXuTjGcrCCkj
hGU4T1G0HNtrZUBNEGEla9I8fVpBmup6FiZPKeYolPf49YHu5x71JJsYubfW
xJDnVh4iYaU59/HNpO48Eb1pNZbzRv2opRN8WxhA31kiEFzk81p3MLfiFAP3
qmuv1WNnu1va4Vdk62+o7QOuC6H6vndTSY8nqoHjnHAof0oHzIxyElPEL4HP
fguqs0REO6sDmEdjdEUW60+mShOskUrOGORN0HwJjRY4ExO/cbZXpWZKeA1W
8agX+ohC/rIfsy9DRnElSSzAWtwrVAf9mG0CmUMJodahPy9vuNq8Pj7rWEG5
aPsULrfe6KmDMh/m48PgmlIBONHJDJobX7D8axFnuC2prEB3+jmevPYs7wVO
cT7fKnijfMXrv1o0MfL8QA5I560Du3aw1L+qO16VeGLqhOQeDMK6Pbt8kooi
8UsF/aav9iAOFsfNUVaJG9RRc71DSeWEF5M7pJIjQc0pvoJoMfwLXTgRo8hf
zaJ/GelsFiOps6HeXgRRGnpAKlKEAcFbHXicSEZo1XJUc/2Nn/f9fndXY6B8
4pPQRny+QSvBVD6uJXQukA1wkw8KOx7yJFLRZk5w40gy7Ew9kVRAwyZ3tz4h
6Uin4ZnORQ6fpn3b1R2j/bHcuzuPwZUUtdQxOEfBhl5sDt7mlD2hcSCe4H5l
gfTCQXi8OuhZhAFshg5JVBON45BTxJv5lwJqChddqIntNC6bmHgQzla6XiBS
U6vmB07ktyCqV/fsdDDxNhM3wdrk/xrbDfdUeFprRYEIk4x+5uRxWkNcAE9Q
YDsgcU3sUAYU/mdXnguHHADbRc/uM1j7447Ip4blofGc7QSuc7MU/6kI52lg
vQiSfapiRxA621f728LTpk1g2bjaQTcVj7lKwOc4mOkYqo3bgaOlDvah8yg3
D7zyLX+FytC28f+ES9VbigWznkw5p24qnxMz7R7mr+TsX1cBwgEeZQBA0beX
TbkeEq/6GNLQupIX6EyQhPtbUGQjavY8CckejxSt7ejQCFEYQ6MmAxB7VoRK
/9+7LdyScEHgpejZ3caEZaQ4BD4Td2QvsCEOkl1vtFl15eHMN8+iUFMz2XSI
DfjmiXQ3OrhaIBOV37A2dB9QJEWrAyGSL/rW4ly6Qzl0tqpQaaVnViqF5qJW
9Afj5pQDAuWekzqAwDv8zTsqvpg7WHy6jH4KjcG3MPIGXk7Ah9VFVFyBmVdx
uUmEs8syZtaH8PARHDHt6ka4sbBI6U9vEdqfOgGed64y18X+RqUjNgjhJMSl
boDiRfOhee22S3Us6rZAcl2ldYHSVwfcMzt2s2xmZMqIBGOMJYSDKFc5HAQA
wMuAW49IT3TUAT6zgkqHiDN+NuNvMYluSXpqHvi6960y96aC7rLzDmDeocXl
54ItUOHee1Y0dKg/sD5A2doZ/7wduNpsJNSiL8pDm800LiVWrUZccGxBkGV+
r8tTxflnGaRQlGJkfPpq/hW8ZuO/o+GrdaOKeo9m237E/jYh0qGi2jfkQx/Y
cBdM4D9YjwZ2dAEOxtHs3+VwQk4kaBdr/Axeo29TzExC7omY8melZlBf4u/t
d0KBmNkvwOKtGfxWe4HEcZuimlIsPn12ccbLtsUsxyHUE1qrwW+r+giEgTLl
ZWkcLdJA/V6wXVMCzEylaFw+IU2tm7H8xQe5NJ0EgJ7wrW/qi67WRhiKqLln
aR23g7WB3ISIlp9qwuYzkq/xW5smVxZT5Lk0KFhAOWlmK53/XP4m2D+MoejM
eV3q6yqhWZbdRstH4DrXfyya8EabitCgP7aEcUWc/5eIXGv1WSQmUAnZB/t4
TDc5GBajGNUPKfW0yllNNwCHNGVivcqFWiwaydtKUmUfri8dujRo3qI/fowc
L7C8lPrauVpeVUhAXAiqGu9gAynw4ULiIlvbFTBLQfCCeDCjH/o84MRNtIoN
UQiuSBBYnr71mGAkOuV1/t0P6sv6YkMtGvBdaZ+cLpwhO56IJs3Shvs/kf/P
A+87IgDpD8PI+Y7ZVvoWbjPVlrbUoT1YAidw7Vo/OnevKnct+4o9R+gpbgsc
fog/Hxk3aNKcX7urkoAg/cdnpNAIV4+Vqt8sLopI4mqiZiaiSV77i7D4QRMg
V16NT6dbFh3UKCIEMx2K0reuCyQuqMQyfPBQ98TXqCm80R6rXi8HLkqj1dko
N6KhyRvbQmnNqQKh9EtuMX9d/D8HDaUSrUXOC4G+G/rAjkPxh1e4F2kX/uin
ifPSz6bIoEVDDc7HjucW0emTnEJ4vob6LwLFyWg2i7yxYgItxdF1WWUDQFIP
9cjnF5q+CD6965n3/9vATCgRkTPoBR239dLOuLlnn2TIQYoqbZrBsgsvtlVQ
msYJdxTJfvKAD3zEkdZ/X8h5keD9wfoJiHJG5xHejpdnLtEqYhPPVIwL46ds
yMefrOMzBVcREl2IWdbhBGv0WinUZ6WP2jpTiOsumT/jrKfF8SOiqlDQm7tU
ZjaeCjFtp3W3JNnv5/v+c3UCrdLko1b/OItpYu524vj7Wh7KlziM8sKF2qJK
G0vTRIOhLb0lh0WE35UAra+CeMxzGcFrJesMTZfpHDybS9ircm+j5Ew5FrLQ
o+dcuyPIeCFr5VosgNJ7AVfyljYCKFfXVIurGrxc6NABURxPdn+quoFopxOQ
j+g3bsHuS6mZQlBNHYw6vXS6R1jtO4Pcqsds60LynEcip6l6w5+fxWWs+HE8
7sSdEartT5YMdO9Wbjx2ePA1j2Sb49tELSgEqap4HmXfn3eGUoy4leuPgcV+
66nunyzKzF7sIZAKOdbrfEpTyWnJvxYb3GLMvMHKIhU1nKefVRE983wD5KWv
C+uh3l4NGpOCNdWB6tyR7w8JOpWnACumBMNqjZ5OJY+2uKAq5MrtDdljsMKM
rbYwDmwlyN0Rt8hVz7r2L180vCeKGRcrP7xT1ALhi6LpsUG7++NfHqDyZAsT
HUuDn8xUkuAIVjm+vb5HdBPtpkqpgCF+4Ho/FOiuNLqdUpNOadS/iZ89LS2Q
VgxbjX54pH80z/LU4mAmH2wzfGW+tJ1JHgIgBmxcfV+RFo/IJI201SLvCJoS
MU+EWTn6Sptc5JHIdxF1kJAO5n3djfWYeVb8+ZKxx5zueBFwE7c+TAcZzkIB
nufMnYPQpo8ufNMu9KGrUty8EqArCP19I/IM5qpfhUYw8Zo0WHgvy+J3cV4F
t28CcIlwN/2eKJuaX8LS7ZCdq5V92wdNQ1h6uMUJtkT8bB8CIrAGVDwTIl9P
eXGSojnl0+ar0iuNqrLwfrW7N+Vl9qa4MQbJ9PRyz/vla4oeYF3KmLdYQEIg
D/6SCDXnPiWZTSdRnAXlOwVZ9RPrPWzvou/XUMHdLcoHqZVEW4zLtk8aejC8
bvcdsztgll4xn/G4bO9yBtBSQZnvpbU6wOn7ESX2d8MAGMFQqjDIGPB6rF8Y
pLmivuapxlF/24JOslRqW07ucG6sd/swdKWEkX4RwH53hcwU+3kGdocMUBdW
iRY/cxyfox7jCTfa9Ks5Tw9yCBPJu+5tbxiSWaBMsAyGSrwg3ko0mwXcAWnA
DKXDKuuid2BLutufAR9YMEoy5tvVS1jSJ7vrbn0eMHJXj1hhquVNfgKecIyh
mkAp1MGld1kYRnIDtFdiPgQQ7CMlK79sFIK5O0CRiAJzlGv7RoGdi9+ckIeR
4D0SGEdtrIdtNf7DHECsJQO0JtB/WovXJdnyAdy1gphNsNd8OKCHQguVzTMO
oX285soZs8IRznKehPeOTc8CMM4CtvNWgro+ZN9X4LBYdgEdNsnLon6xtnlz
8ssDtDb0aESsRlxDNBGXOCw1tNX8HYkAoshq+tU5uSDxJiunD60cZNkZTIn0
qsup2FK7Lc9XadkKOUX1e0J+9T/bp0+7Ijbjugsg1lrQs4d3Spd6/hEYKF0P
CaQutiQPQTcyntwUuxsfiOxyU6/y6q3zAZQtKfSNgFHWUXKTWcCxQZWJCPhI
twNCWf+4Tl20fpJ7b0LkvueeUJPBlI6tNQbxk0ws+K9++/zIO2tBf93gwXVc
iMlQI9GCiWnu28x0EWyrFV3GDpR3joFK5UIZNOKAssQxa1OXPgkZLemu8/2Z
vREhQ3v9e6gwc/NFYtcWw1o2hOYK+xVdGketicGlmcOi3lZAa1Qg3uw/vcsS
y5cFGFGAYLMZlh9+mv4oJrwYEJ+qRY7/UQRw1QZwGr6lr7vJKXyMqhi5U3Ur
otHxe2DD1o+UeMhr+FemY/bi7wjx9dlvP6N7JJ4gJysZzFkRCIxhyniY9kqb
hBX7/RqvBaucOQj+X2hCj4mzOoFiLNmBhRJ37cfzxAy5EEarvGeE8PJmtXBy
AgzYLhVbv9UvYq/1PUfJUtBSWLHbF1VUNbBzkQvnNjnYpzp2Qq0o6R1UIgCb
lxqXTkaSRjEXiufDNHmFarEogKzhqwxklUpWKedjzYlRtmzMJ7jZaI7Yaosa
3seXmIzOsoYZ1SXIeuMFrWG1l6amJEZXCoC2aH0y/FnmdZZQrSjXOBbVaX5l
8jdKQfbTp9/kKM88L0ht7GBOQVCtgEbtGZlnaxziG5wOmxpmqwa2wVR7c+v7
0Fjn36xP+k4UmODY3EKLAKFI3bnk6cgVtmDp+MfDMvLuscl8ZfhIsXt02Smz
/oqH61ZzdtJNST6lQCrsG85gZ56wDHItDdgUVUVtqZBTb2YPT5xj7ibiI3+v
QK7mkddGb6rLYSrZiP2rCLEmWr9apM+eNg0h6M57lAxlOF3y/owejubX0QDa
mj4UQilp3xH5qiV8w36hNYQExiT0FS1dVk2SMlZePT/uw0Wi/2NFFAPsp+l0
xoZB5h1mtvZ0mrw78OuzcnusbzEcuZ1zeUKTsnoupVZ85yVXYYmKYrqeSAF0
OxYQ/SfOg2eJXscVKEXm87N8+KObvhRnvh+0Cy6+UuOV0PQZAxddg5zCmIjz
KR8C7aN1AkrxACV/K1C5ZRRrjNGjE/N9t3Bily+dwZO5skFZsrDS1YM1ZgGI
9jTmFfdGKfv9hppPGmMlcU2Zo/E/e9wYXk5F5J7MW1vquppkOYmJf5Is7fLj
EeHaAdO2+iQSGQPXsnScdjKWFNuTJq4+CYToBVqpmjgl5v5kUu23ZQGUvBJY
VZtpgMED3clIj58FuKXW7RjvVjkoWvFVVD1STdqRTplPvIs1OYQm34BdN1FY
QO/b3M+uPitRzvJgfTmCWZh+epaHQARFWHDlijNAxFf6OjIQ7qHajYPknqUt
GzECRckJ2BYf+YXSc3zzITwIRDFMPydcLVCWQZ0e1eea2urOwWM9vFj6XQiH
/dCz9Quw5dljZV4ldhTk7dmwsd50AkbzPM0RZTscNkw4Z+VFWyfQHQeHj+2Z
GukpKS7oOOijl8zVt8U2Tkh0tP5dmAcKk2c7ha/rmKLMBXV0mXJqwbhaj9m0
S3GF6immA7kMEiTUEZwdMiGXGy0QKKnB6dlzrFLz5NFjuJ2FPABJPr8NksLQ
vTwlqoiAiS/H+X205CrJm7f5trBm/9CRgsE6HmiVF9JRGekaSD/kyxKrpHoO
LTRpDH+8Q6DeDmLvLK3M3vAVjco2i5RCclI3qinPJgHkBc/2R2KYGM6CtfIA
2LrxyZFlHJWMgQOE6w2M5PEwsB3bOCVAN+gRMKDZVr7ISLwZqS7uf5+gH1h+
UQSXnFSLY62vLLC8HgqIjlNoVu8WdWwMGNmVhGjTEsiMHJ5PHE3EuxEY7gsZ
ae6FdvXxsOTSxCpofjcjWCuK1q7O+v98QNrkyEov+M/4pJcQD5ighxgE2F83
l4zwdG0dWff8n16l0BfZuOuwO9I0yLLaiuxpZV4GVLnZnXfSBao8w1Sy4alp
p8C37T8Bx57DjJqhVA8nbDNAiqxsIVUji+Ap4CDTBXdiXLnz803ug2Eqp390
YyXOYqJH/3ZfhJmg9Yt2BVvqK1jjwRWEUHGj2aazL5tqLS3mRLTtJAk9BavP
qiNAkqEA6l/DFHjbAqzWBp2heIOmAgR2Mkble3dj50Zfzt1rEAJFYOzO4nLk
8CmCFGZ76PYpZ1AsonPc821G3Nw683YQPUY5cQIAyYPSu62WcpOUCuKzvVcr
/D5iTNQUOaZe9O4FjtzHrYhiTRXiddRvdJ+cRX+ZJr3H5tBJDu8t1KA6Nrln
o6pUDC2KCsmjjl88s+9qERyq7Gj6spdWY2OGrvHDnM4MWxtYqkeFaOa/2kJV
v0d2bYLTWVwwncihZlmLnED/+491IARHZJlEnRSFs9eKVKGESg5zCghwxilv
yS+en5D2wP/V2QE4nNorZ7aXy8DmXxsXWcCSRbRPQ949t+abm9jLfOE3cteO
/N0U2mrCLZWZ+UoISyhLIgH7D7/mJYe48PnKI4/l8kzZFRt+5mg+iXJUO/t4
0chUlSL9gPqQpB9hOnEq0+FHbajb8FNqwSErn4Gc3sPhKXkg4wT/xhky3CdJ
lYrUl7MI1s4r755xfiOfAgQMKqhI13CCzQUASw+UFSIjsQlRjcHL3lY0hinO
2O0mxhEX/Zden7NVcfNQtvrltpzku0BXCWK9fHhRTtmH1RPrkPGVuqXjjI0u
J3ycEzaZ3eWqjB614NJrm/BMWlCQ3Cr0opiCzGoH++BVbU5cWiu9gnCrn39R
HyZ+sWMzxGVYjRCLFN31mP+Fx6DLt+H3hPkmeebsgDSrgbTd2RtZu9kUnkme
wODEb5S15KHYh6AHHIMSTkTJ3xHQJBc7Jxc00N4VLWkJLlHe/4E0n7z8V8ko
UBCRK/baRBCBN6vFQ/zRvsSDRf8CkMTIoERxOPTwFsdbCBXDnaBn7VfhbM3f
0aSy48dsSGpGH2lVqugS+EUnrSxjjNnppp+34lNzJPRCsqykFmTSo2f2eSk8
Lv1STtGlMZEa16fWBtV8mKZI7BL/hTH1/KXyjUtWuYNtQ3W5YcvtOyU8AXwH
SrOtuDt0d1mE0rBMdVwixGZlud+Us1vHO9E5o7X6nJclOckA2r5vjePZqnz8
XWnSQMJynECZ3HkFuTyd3ghQQfMVskNTxDyHWdd42DgLOgJjvCZjXyo7hKm+
N1ySU+sd5SowdcCN9xlvdTmTdIq95pbet03ggFhz5ElsCZbX2lT8mHhLzJWp
szC4Pd7lvVzWY2MIzNJv4GwX3G3sZrFTu0RABg0Vvg52dwd3vwikxaU9RXJt
ANVY77SmXL5tbm565J/M9MLkLqzIaJbk/JWywRrD5sGbmX/4vrwlAvMEC1MH
2oc1ZddsG3fCgLhxx0rMiHdCTWBlO7m/E5eE2WU/C8Ngr0ToDJd08cKE6lq4
2p16U3Z4SJazBHbNWbDqNqiukEZvi9KJixyWgaPGpnJRjWqu8ypPGs4FhqIl
0gFcdxk69mGE2fSi0cyFS6fPGjLkV33LU7RPlc8ufWHdeLTNJor1K2BuE7+g
R9tttP+m5BOSxpTWwrdq6ofkAuvi7QEKG6TEXTD5htDl0Iwq6pG8GfpUbxoK
DyiuqvtjKGo29xpkInD49d4SQr6ay1isM2nl1wZ1dfqV27E9ArJHzBNV1YKK
ZPGYItgjkC0nIUaPqLvW9kb5Ydlrm4X+7b3Z03qSnDVH5AbdOzj6sq/bNja6
P+7NpDyJogdshFAi5XAPuhpqSG+okwh3fWhP6owe24q1Tf7syLXqHIWkDRlS
PfA1t8e1tkr7u0XwC/FNnN/Zt5BaNERuqapEz2HWCWe3brlokge/WzYk0dMb
e6XGI2GS96l9NEOqhEDyOXrWTotFKvHK+5IgiBET/jcpm1mLgX6G/yyLKlPY
v/BNf1Wr81rzC/E+Kq2WA/70xl/bS6WFuYZPdWJWWGSF7nU/QG0q+S0KQZYa
noZMY1C+dmxvnzfPne90grYMyRkZXqBR1m4VHTvyWfIGkw6H6GKRBqRvZmfv
wMuDsS3+smolfChXSG9M0zDkWAw5qyyR8rY9hmJxAREvjlIo3z0M6imuuC73
LBPZaIsIZ4+DdbWeK5bFg2Mh2Xe+24DiLsGkYbcIJpwTEOwrpnilmXBI4EUp
Xl7hqUe+72xQwqJz7ODUz8Ml/8+sDtm7HhtEL6b2EpwiCEQLQUU4PFTPTkwb
N11zpPyws+LjhgjSsEHiYwc/0EdmwfdGCG5jXjIzZ630XrowwdNVQn7ksqB2
SLuC9Nh60tQIvVP5fEg7yirq8fP1kWjJ50SGoLuvvMucWm7F66KtxRQQJjTG
drV9U+d9I5Iu09rbDV6a7rpwl0m9DLGU5UepNKglQltNrQQswSI/aJcWBvsG
koL7zcPcFuspZ4Hn5xiwkhcf/ogHyarGa/M2XE/MddOzASSngLQEBVjiDhSt
6NEBeEL1Bb/eRLHTDf9NcNtgCB0dR5M1k3Lz1dkBjvAeq+RhNz6cj4R8aSNB
R6aGTNrWi+K3l1scdBIhLL4qj63FIeJee3W9YKl6B8mQttHVGTIqR2pUhH77
znxbJKwvES9uc2mRA+JW1UkU4cxfkM7q1Y3QZ/hqmAVCCGbEtxA/K4EfJG9u
42WJqXckONmNA9fvChip3wRn/2Q+jAQeMXJKCzsa+sYbGx21MysnU+E0guYq
a1tUsrZ3qR05X45yAuCrkVNDtKR6oQ7IuD6OcL0cDbgl+oeDSZPBZ8GbIcWR
Xo0UIcpgMMUfEdux4YsLzGxh84totN+EJwZHOo9z4dYxvDdNVPZHdlhM5Qtc
975eDJv0ryaWDm5cpfGLBUFjW2upfA6lfKNckwWBeDei6yWvGSVznMTvubxb
z8DkykIz2aPZrBYAVbJa/KXSY36Q2pmdOyOXk4yDLysd/Uozc0P0CoMqFCaZ
KY24Ocaf7qnBGakmyJxiT20DvMnoxFneBSKwo/P4WsL/Xt7Okuhnq0V3PkbT
5p3ROsHiKiL0t6gbxpeJVcYGL6AkcUJdQGYKm5NpYE59wHcj4RFkYxDz7hcb
i8yjZCupVaxrFOucaBqJ+ygnkvXE9zPQG4hXFH/YaJYbe+RnP4Y3x8sTH/Rl
798Uxrd+gRf6oY8vFNEaQ54bT2fXIUsFznNRtPih9cqnlbB+ItUnP4OtJklL
yXtlwjWqNufygMfdemb1A9joAI6/kKKU+lTNBmZd/qrUsh/ZUmpVlT6lNK9C
eUYcv1pclkK5Xz2GguDgEaCGcgOhfR98zlAGyORAIDVYCrfXBIg9k/U765Nb
cSO5OrzDWmEVCsRxNzqoxLs2ypn1qIJR7WzfC91h5PeWfSiFoaGwWsKFnYWc
NGPHv9nOYcXvS8GLEpr7KEAmZjpoeSehL/pzWHLmYtc9BtawqDifJ0KMp06W
RVxZVgeylQ5iEHAim0NVcWtjiG/tmChWG0til1D10UrVaIiHRJB3tpaJ2Xsr
V5noH3+yfh+YzMmfjifxvIqt7Lq9svoUIunu/KGNmn9beu5dWW3z0/4/VL7a
CHSj3395nJTNpxQ/2esMgUUVmuwzYbrKsEpL/TiHUtdbePajM85CD5k0KOVp
KGx4F7bF/m0QNaF4Tme2aZMNRpihOM2hhRFfq+5gOWrq0ZdFhZRe0LEonDfc
fMv8a0uVGEp9T1waJK5uYB/3IiVcST+wuE5sF9d6BWYIxDQLZ6GRER71lmap
KCKF4MxKxJ+KJSIXdQp6x66cjaAtNZGgaCTZxAXvykEu2yV0xpk629rcKynM
e4TyNCAn4HM9Essvd50y3oHVwX35rn65XrVUFnu+8mOdzCUNN8FI8/u8rbnl
6Tr145Ld6DkgplIUnNMZROxn+/LEVnq9OsYMKMfI+Gsby1xgVW+bOMXsDhP4
lPnUgnbu5WAto+8fBKkXi9ZD7X6PtUBIKUQUDJGGilzrnoGGfREMXwSW6ci9
WhJGCtAmRQmU9k1z/uVmm3kEQTpLSg9Q0swznBRWGBJemLUf02S2FeD7hk6s
9wiGaKiqEXnZTZ1HBL3JxQGt1nNDocqQB7Bs2i9imFNbSl1pALJqbemCC7Ld
A9gJM34bgqBaIOPepdZrcINmrnFJLS0NJha94lBsuRfn7qOURMJmYXkE1Bfn
wi0CdVx/O+W5Fp5aWLD/ynsoWCTgb2Ujz9NPcftyfqEHKOH/4SlqTO197hkw
h3HmG/kPSb+bnW4+8URn8jKpe1JPX6UPxGSFchUD1oPVtEPTIqTOJuw+39lY
sc1A2y1NR1m14lYLQzvVe9S28OgBtoSKv3z7ZgOyBGib3IV5eqirw1r2QK9h
xrstfOTFM6DWlyIqtaL7QCTUWcScMv/PqLQ3EsrvAHuqm0NYsNE3MB7C2+VX
cEk5GAHlK4UnlhqTo9Ug1AvcUG7or0iLZaWG9zWZ2EKMiMTwKNmp64vRl6NU
bPvUQDodg2pCV7LZWVO2csid+5UGVOCzVlFWI3TLVjNRzj01Hnx7qqa/ujnr
ka1N+BjUq1+B3u4DDAAxFlVrFf8GeVIOl1ac0gc+DjdyMoy6WYuAN3z1DfQP
5nUMoiuQvDKo1pOZSANlNf/CEKnIMNG8f6KLo+Kj2RFEdNKpDxOYnzPd8gDl
1n9Epk/cD+owgRnY63lKDqKu1a+CdvpucRx2J6T6pHPDKLf91iCl3npYrp2p
v0X2jH3BeJdny7OPWNompFs8Vrw3Z12G1D2uPHsbAlAfe26awCq1HbsviMDL
d2vo5ICRAJSUQ/r2LNRE4SuJLQ2Xg+vScD6Aby4pTUlDZLqfUtOzuYiv3xvs
/zUcTWzj1q8VdjgTZzmgEnNt7AWZQFrlZx1ZaO7tPYu0yN2GDd6EUkj4SY/c
oqH2ieQ46lyiur8HjVjxpX1InuwINYDUr5QTa+Q/wIycRoj8cDPQQyLKuQVv
twH9glZPyhkdFtCrwBgauE+KfO/cxhsxVffnwXZHtab52iDyuWYPnUMlo0JG
Wy6AqkqKZWO7+CMV4hinPHfFpMn8CeJbUWnmUE0dhTGCzzuhcw440pxHYj1o
/ayiMMrs4Yr3Nj/EnZEkigL0R3Dz5cXnpRC6kmnZuviCoTns/aCk0iaSnt29
68XlWHCZ41lj0ZGhVHtDHMDGaAW6aw1IQXUyyVKKT81Qr3ak2XZ/LoQSnU2/
naIHWcodUJKekyVOJSG4MVxAQboc+9JlRkEPboBOpHtTNYnM9J0W66llgIMJ
kXA9PnLrvLv8pVxon/m4tX6h/9mTWvE3WGUqTbvQqRBy36uGjXm4D2EvQcH6
GD0ApSNYxgyyaL2XIGeKrtRLggJ6aVMZdg5H2EEfKcNNX0HoZN7lJxDt51gz
hDQS6binJ+riGfs9ajPD8PSTXN+eO8/hR4m6euxdhsoezsX8n7C2PJWX67Fp
6k+QXc6wxUFdggALuj2SIixvy9mz4Qd1K5rC2847QOc8bxF1SSmYYNIMHKY0
MV+k22Q0PmeA0ZzXZHcfXvULoMIjNtD0+Mwx8rxImFqo342zLpUJqSYcOxCA
ke2tfRycF7/7yykpZ/dJEG+h0q8CsEnu8Ucbt8asXRYQ/5FyNLQeWicTya9A
Y/FFuZrK8O2RMqI2weG58XXSThf6KIWI3nYz2PkjlWqyX4RX5nQb2hslIwUE
+wK5W0wesAlLGWmQH8n3brA275mSfWaAIoUEcXav7yZejvu9LD+UilzFGwac
2rieTqUajnFUh/ZJ5MnddlOpUccKvX7kU4/LX3I21VZFdQIn6ivAAipRMVwD
eLZ8HV3qdvyYx/UL+9UAUM2LFNNXc1y8KwJQtq740jDDgl50yjgiLsjuc2Dp
Cv/ejXdJ+wYaTV6Jn1foxJPC0FNSCY6XqnQuOr458uzBU8teo3qs1uG8m3cL
cqUC4pqyederOnMibkT/flsHi+zNbC09jkRVchsILX9ODm9Cj8mlCl8NqU00
WueDhgx/9VybKUHz5GzDCu/tUD8pbQ9pIVVdMsCa9sYynynY+EJOYHleluSf
g9Vdt9vK56jozLX63lox+ubzqX5VLKtr5WIPEjbMQxcMU1XBf2LgaDNk70UH
qyz52jrxZEzYH5u5wbVYG79CIsQLY3gjucgpiVre8vdjqVFQJR414L8Hht3S
auORqaayZIUyJh2SqthCvCWGs1CZZ9n3P+9gYNh66dHQHpoi4cTmzBkqhofF
ZgQvt6dX53twZ2qQuXKDCWgMZXI9W3K5T1XVVeAWlVojDLTwdbyY6x3mlpfh
ZTqlGSbue8qyOT1NobzXuGDgOq7f/k0V87CgQUmjlgHrrLkJtSxcPgAZLfm/
O3ozaqXZ8MWu+MPiLaGQe1XC5+foLml8O/g80SaVS5jnfJCSi7FFM4Z6MReX
xubYhFr6+H7vVTWp14WTjnUOZgf1Pd/4xnjiw2gdswBp5gV//KcBt1zOvOWQ
pv9zeXsdqG9rVN9SfSsYtzGy8PYTj3oqOj9seipmzwiYUtKVVxzNUos4n8Ir
9Z6UpQF+JDMxidi2meSVtb5cKxppvuWZPIUS2tktnnQVKnK3i4HV8sT4wU4i
wHb943JDzucdssO7s0F5MhP4djsgSsSVUMDyWuqxqUyVHKTdYbNgSqDrmseX
DnqcCdFaEPgLs6w3XtvSHL8V3d5XHWGvwsRPxDPPX61uo4VVs7/1wngEcjv6
vBGbmgwIGxE3duFk4ePVKLtCEvpWZiT5IyXd9iwbvsUQvTm7rF/8Bty+tzfa
SsIKx+oMqV2/Q+uuZUg2lEnROxqX3DfqFI7bjWD3OkDPmo81FvmvpkcqBpr5
cEVnfpaDwqwjT3FZ5Xz73DMnhDO/hqy8mjw8sr0aC94UVht4NUFpURRmqcsk
Yz2E5a6pL4DHm47f+hRC3VVHOj+k+vBaFIx8M3QFnj0UtgQqxd5bisC2bXKw
GnTjMZH63EeRc4CHR//c6SPb3N9MyJrf4XGSjhzEyO0OFnXKrpP2psW79aZZ
td/STo6C096OOaOF6OLm18BGTLwpNON5pgFOdTYHsi1RCsDxU6IoNkhV+hmR
J0/ZwGpv7YxGjEU/UC9421+vhYBJBJdhQ9YMHaGh3FkbemE0YNT42q2iaxf+
Ze2w25gFW884jjmgdj72XN/nVzsVGcxqLYuL97vKmIcxgCtv7ucA/DMfnHid
FctAoX3ZbgJCDxqtutAPFH/UO3WrYf3NBeBZ36bE6ZLYBdO0ctpOzluvR6oM
W/Z/83OjUvI5mqS+jyFKpBLYQp9lCD8E5A/kHcwJ6kdqXO3VfMuGXM123YVm
o4C9RiTstW5aoDhgJmqFpcU7QJswMswWy+YUwCPCpe/PEokMAc380rKdKt2N
rOmsuEKmtm6MvBcDCoeu0XrcaZ1CSQFv43zjdKCozCwGKG6DN6r/3Br5NMI4
GWEkc5WQmM80t2fsS6biu5dQ2gqsR5JazD72QYpFkuj37jC0APFV5IhqEy2i
RG2wDSFYwTxMg7ObutxESjK01i1/2gcotzrePhICC9KdRFCrjiIhtDjkQi3r
+UsGMaBZbTJ3pWOGmwqQUolRd/9zrRatB1U5R0UwVZJnthErpY0bDY5AWFLy
QoD9LXkptOz/P0Rru1jrw9q4ym0uN3vnEoSFwK4WVLb38YbJAc/m+KG6ZBYS
we9SXzuXcnv9zuAn/KAqqemtN0xS7bnGJ6KLU+qtyhkhM2AmlDid9Rbja0ZO
NJGOUlj1wNK9NYjpMC0cOAeJ/PWiX8LgZ7SA5wBD/ScPwybc2QJiomwZ304r
uQIo5f+tgdYYcOeXAfWGoeklMCdyw7eRo0Bovg1ly090VC/6inQG+fSdOnZc
fHSODH8KQbeBkjtfEAZutYuvSQ9btlDkUyVS3mCkBmJEOf2XuHcuiqSsKnch
vTMGg6kY5ea4BdU34BnrIevOW5OzVk9Ki2/xEJtohZSnNDGvDEzXJqEwzUyi
Xnb3gY9RbBp7jiz4hK5JvmLvF2XL98d7luNM/OVTSZXeMjpudPF+Sdy8KOYc
7cjD9blo86A3BOvLP5Fc+xQHNYe588wkEegLOg2n+q1Yq4vPRtU+9gtbppHn
xRLzr2zMVJ6yjgHom5KptgxoMlC8UWwVSmVD8BPn+DfMOl1PQppzGJja3ux5
GOYeeApJJD6MZLps1gbofD6/tVt2lrWoB2/9osMWQy2vsJrBe1qmMlJ4CGau
WFOHwULLtGgFGW7UJ6P38PRP7RhvEkqOOPCb1z1YjpeB4gMmkMWIpZ/JWsSa
UaJNliFYMY6WHoKgIcW2W3wOEGwruzuGAYznwEZGpTZb+5qhDdypmSzAmfdo
0xHfqdMNswvzWl0T3P3IlmbmXQo71HTbhE37iivSLCehmD/A1+TGmQecCDX7
zu+TmKv0SVqVbRsW0pa3aG0ioj9bF+Dcs/ZjHaTsN7UBrgoV9vg2z+kw5BBZ
xmg8jhPU1I1DAMVszWHLAAwvXq/EKRc6VM7b655rS2Vf1KRwst/sUU5800ij
Cb+TZszJAHHCFaYDHQM1pLtxvCi4wG8AkflqSzCfL7jsQ/VxOi+sN8jCoKSA
iv70HAWV8vFn6Cs/FzPVDwXiYAkcB54yNDPfXcTGL0+hgWEO8VWLGykkqk05
8NWoFBpSqW/zKNzgKEg+rwnv/59u6mBGK2dHdgk2mnwDJQxS/l5sa6AFebTO
vJNb0mh2MYtgVIL0qrNWPCidqZRIxVq6YxqhQZljOHIoW29zJ/VTEhucNOt9
ssRv0Uz6Rt/IlFDhgSbzrfpI9D2IqgZy0burO2jqkmDsFavjPoWUCPxGwWRQ
H09O15Q9x5cw8Q6FSwvFiJ7d+PL3Ido+DZkxbn4GXPzI0oM/5yQL4tSH4aqf
kf6itvidxY0b/IbL0mogoaBzxiS2DCfHKPKucUG24Y3t+W3dHkHYVcXrH3yC
ht0QTJckINGpn7rOgwp5qeCuX2zCxWug+NPQEslPeEZ7yWTPKrJu+X/kyN8h
2J3PCgTgARMX9KE0ldzgcvrzIHTYW0pfXVOz4Bouzzndqeyla5pg8dYSdFvG
yc04klA0hbzT7drJlYwOaZnjJi347/7MSeVdb/kJUoDlTElknmHJWVuerQZG
AgiOBw+JS+rrJXGjxxlbwb4FJcGITUcLSDp9CEfFlMZc6hDwfIbl1K1ngbqR
yl3gkfnbwFe40GlHijpSTzQS7S1tQnl7l9e5GIr67pncz7GAgFPeEyOn46rU
w8P0m+QLy3xMlsiXzcMF1UBaPHcF/6YOiaXc9zxqUYJoedT0Nf6M/kNw6DN+
fNupKzUVmAtozcQc6MR6FifdaV96Mcmzn9mtMHSLVFY00kODUu24cLMcLAIz
Ccpa2J695TUwTxYI/CP208GeHD1ds8KjxtmC/4iwgH7Ta6woojMgBsOZOUcr
W3zX9zueKV1JlahjMM8EUWv9gSa3z117TMIlEhbgq3G59f5dvXGr4qtP0lxO
GC3CTQEWAHws0N7oIp/YTzpc0ddA/1xYSapIUHnh2VMf1EhlveHSJzGfk3hD
opwlkzPCqJ5mUL5LFgj+ZkZfV9d4EwVqoRquqEbNXzikTlTAOiNNssJYNc0b
DfH0Y7tKNAGjr/dFs2MzxgvYHmBcaqnnojOt4FzjSvfacAYJ7/WTPpLy+uom
fHOZnfuS6RdkCSwauoob/3snbFaK4VjG34FJKUIA/GbUz9Tzy4WHMoYhfUU0
pmpODk1Pt+Z4kKl5I4Y8f+9e/2GP//i9Irf44fypKiwtH6Jfiko4qrePINEO
PSAhVHAt6BMORkX2UFJ6zuPqrp9LP8mB+FcUIOHkGHVK6H/9yzPHJmaj0sd8
U6xYClntA2eMK4fCHQtO48KkXoHp5KMtprcCTPRxuipzLWiJVibv4p46yIEO
EpLiGgOMyZ2Qm2emf/l9Zt2jp3qsw4X5HZYnUi+m7OV90e6UW+GBlD+sZcRC
YlbPCHeeoHddNfmfMpOaDF9KH0L+7tPXvO5W0TYcaicV/0BHeTekVTFgEcmm
iq4FKOqXmRNuqJNj8YfQnh0fAxGZs6C0g5QZ4fprsFPI0fz1/14/hCz3C6p0
kenxDYG+X4T7tNwbwLFJt3Hs51+3PwM5ivpNCbc5TfcKBfo/cSX8SLllIqgY
t48y1ZEabbB2Nt4VXp63qy5OqpUG4a5TmSLpWQCLO6tp9qRt+CnFKTYXyf8B
LXrbFSmNi3aVIwqrnV1CybVP+hBkrkXfJFjZlFnaOs8MuLd4EaFr8r8VhWOq
246luzmqOIhwkP1nMWbB91N++iq4MK9UJIhKRv5nM3hstrVzxC8E4T3rKsVQ
raax4aGiBQ1uWnNuZm3DPDDeZV84FOlDoHwqmFd5IWXYWiXYrxzo/TlUSNGl
+EghIdhi8kZLIDyns81i9Ik2TQBaRteu6NDwOvnMv8uXQhrSoRrSCD2WZKrN
f493CNvi6wjKE7PoE3Cl0GMCmK5F6w5dIPH9piOKglLMqu6V1TckR1YsSkOg
65VgfWyrRwjn1HxoMTRQtQyoYytIFDuZT6VSHG96JAMrmwM66yZ04oeZNvKs
qIBOYHYOM11NupBf9HPSJo5qfeHzTzHBrhIgGFZhl8SsEpnZW5bUxTLWno/t
uqOXan95gpLJRmo6PzB3h2zRXcHbAVIRo4U5fkwebDxUjSB/fo5hBM7oq5xD
yuM0Rw/hBn8rveWt/X97FTCqIfr5IiR/mIMMwPcZtDNjrDWJSfyB391IJ28I
f5OJRoUltiR8EWxvcafzDOQi1/U7zi3zza8tPTKCKh3yIngTa0s85ODmPfmb
IBibuaNKT+iZB4P2mcWmPpa9q2w4uZ+fD3Qf+wAvz7Yu13O4IK8QXK30canL
L9OVAqnThe9x+NIezSxnuZP7Ac0cD70VljJtX+cfItWxKZE1hjbpzFtF5a+v
ftiJosW+yYJ26gx80vB37kXSjTSbnRrvIyTGDHHQz3/NCaMjaCl1ti5ujeT0
Qk2Nbmhv59h7Bto0S2ssafaYUbze0bzZOsLJnnoSUMkfXBMzCaiWij5Xt5Cx
FhZ3o58z9ZaE30nv3gBx8auG/vXXNjdGV0O5JRffK7YEh5TmeSvByiWyRO2+
yRj0aU2jOKrnxgInrTYNYSyxDLhTC+ByYyXPkwif3lzcO8faDc7xUnZF5adg
iLfOd/7npBXgLQEkHcHT3myGHJ/N+VPn4+QoerItwcy3b4oiAjPEfRh/mz/9
ZEZHCMSrFLcXj201zCsXnTppwgEILD5BODasnm4SogWgLgDAvOejUYBdXHQf
agWhh6bxxtgu+P9kD8DRtN/nFsgwiHCD0vWbTUod2TEYBXAQGJfbqLWasnMf
/oNKnFSTwzlRCkspbV1rQAYwCxJE+JGLvoyLUb4ayOZ3bjhbcXlTOqTS8UsX
MEuz4hmAFIfOiqQOVW4WGI07zDvtp70X36RQkiLrG1lgtOb/e/S3cO/VZAC4
dT2C/LldngWw/uQO+O1e6H7ZR7PFzSkZU1JYXI4rxOFaTIpXHpYyqeDaih+4
h1+SxUlQ6n8W4lgMlBFCCGemSK9Roc9/Ier1Z7KNDepgv1YinI5DWXHowFe4
JGlZbwEjkFDdfl4g5RgzaxmYlELxr9CBp292j1TvrAFcckUI3dEwOFIxm6q8
4U27gE7jErZvcAZp+TILpnaOQ9o+GkHlVXFZiA0EwXykr6SL+S2+/3Ut1nhb
To2VN8OEDtNr5wwL8B99RrCMqrJoyc0PywGxhNRPUyDky5tGry3AL2qhCDqS
Jngu2+ow6eYRVPxvBImliSOEQHpUIkUEzywj55j9b6j1NBHCXg49sjb1SSPT
O5L3ZFySFdQkKkDNh+jLfmOaxzscE4tHpcE/woTwMOFE6Me7cPuiHulT3T36
XdS6vi8fxPNHqCfHAw19VIcL1RzVezuSSe7xutlDrZHuSQpPBTnq4otEhdHZ
5wPp/YvkQmW82oyHuVlRfOIPoPm2nRvxLlzAoWyrDDHa33jphS6J5czjoH6S
O3GQSEinJavd6jg58pxGxDZufTYXsVzq4zj8v4vGVl11o+FWNJcll5aQYoIw
grQzFehopx3FDwJjekkAF4njSzK4Ya4BvH+WkQBL8jc92L5r7Isd9xanVFlo
BFtVAlJmU5SmYQbqhIpj7+TFKoo6BUn+J0iQ8KtBcbg63V4VLpx5IlHLuZYI
b7eE38dHj/vBMnhivinmLja4K4KeE3xof/TX2XDuFI4a/JfxP0/FcnYN0t9F
bQ7Q/JdUGNuV8Z363f5BsdlOuSzpxWGnm4i5xX/dMgck7oLaWokU2UW5KAAg
j2MBgqi7Zr/VnHONVEA/HILyE4TcR4EEzZPcLuFDkbt6Xz3nWxV0sE9f/nLf
BFPCG/svCtm+7yQl1wimmnQSNxAwp41WXmNm7pwEi4Sgs52shMej/k9d3rcd
N14HQ4o+QGmVKgi3I+duX8P8eq93CQLO1Y4jF9TK+Z9YwHlQw9luzKlnInDA
T8btO1jGltCxcT9gHMQPHyqbNG/KSpNVAbERo0jcw4LfjrlceoPt6n1GknXw
S776jtZsFO+1wSaMtciKMvTqON7H/FgLiGHxHHewaj4a8mFyl8fsr0aItnOD
oBg3Ncs/JHFmUd3kzz8LGn6NrEski97RFff7ZZq8aBUaGIoKw72sPErtjLHM
3ad+3mWGkuMkFy3Uv23XaFf5OTBWeN5H7AdyglRmmdhOpfT1BAtJa5Z38fng
Y2ZyZU7hDHthJ/bByfKjWkK8+xC4s3ti4zpfKBXQdo/q5vWxIsX44FZUK8hN
5675IgJmelLLoK+oEd4lD9RXhmkL2H/grI9NuQJRdvlNzmklzlCGnIWl3kPU
lBCTMPU2KAB7B+YInDsc6z/I4x+PyndwR4DT18r4jAvPbQ8RubvpgBis4JKx
1OySQPr/LWU6AneXPzvINQXB8aAdP8X2dXlEKpeY9f+EIk6NQynbbGcpXDux
Ke2wbYgdXB2+TtPi89bspHE3LmSwYM1n+uD99+X0mG9yncJ8YAsZS56Or/C+
Kxh7DBtNmMt8gOIBMJLQ2ErkEDj1z6eZ1uj9+0ISbZkTdTDv11rKJuX9JCAb
SH+uQKf3jNGJp+5GRrvcP2ZsVj7x0EE1FyTVKSmDyF7pLrmNZSadWjKITDxg
i/K5wBTaqvIhj60fvZ2hhpq1KWkpR5iPZCPZ+9ZL1sV6w+XTTlThIRYbBue/
me+VF0rBnrjwcmURIG6slbBYtoUiCZOj54TZRiACoMToJSkdkwD7cjkla0vt
7euR9+4NtyYdTatSOHaywkQR/j+a9ydlb0zZ7ocA9lEtxCy4yIwkDQIVn8+Q
1oLBUMBW/Q7Tnn81ooGHJ2Gnft2sqt8LZfX9YMW99EbNdPK2Un+TlgP3x37Q
e3Z7qvK6vpnAh/40yPMKMhD/U7SBsKPv/8cAZME66JY+JbiiSnx9pKjePf4l
vx4ZhB3NQ2hXrzRmPudMH1/PAAoPryLglq7seTpRxwUXSFWprI+6ZbxvWubK
02HPSkP55BokMnbF0o4048Dw7uS8IfE3MPxLFdvd6EIhBnWPCxD3j+DDHwRw
ohSa/c4rxpRfknyQCNiZTyvtjO16q4trdqQB1XzC/DiwXF4ZHX+ktp7sZvg6
+/NlnqfBGh9d5NlcBhXM+JOjZKOaobkvH3EV8G3AkSz9SWWzmQuRu/aY7Ekl
iVWo9hb9E5HUrdjIKW7ptx0C2cSaMB5fTwWJ9bjLpFFG2NaeunNynLmDOihJ
EySKkGFg8m9QlzhvRxU/xuPMrjWAMQKaDlS4TM1OP+u4AztEWVMv+2LWdWZG
hKfRHQfnvXeQIOdQuPajDzdtWNLF0pHgtN3/4OyV6dP5Fhbo+V1TkC2fRvhD
4MH51HfuSM9ChTq9NZDDOX6RBpfebzpTfsEJCJ4OzUPdqXvfwR0gpMVrIuR2
gxTsS4knxNw5Vlh9q1rKkx4GSAb02wwglRRf0HFMG5uzUx7tl4D6RUYXL1wM
c/N9AmUtL2qttIrZ1hj+sHQXhh76Ibo7m7oBIIkRudLSkzUAlQxADzsY1jlC
xgnONfCyuJN0OiHvdEi14h2HpHY2WhtJLZKh+xhJlFZiUj8BfDC/tb0mBgQG
HmHKECzDapCwfEU/TMT6v3zUvouHKtgJ6f+MeA2F9NxTEk1hf/kUkTVdcS2w
XSj6kxww1XG4Q+hJoEVWilaBvc9sgcvzsZu+wuFw7jL2azKuhDNrW9KoI4Jl
Z/Ss4unXO9BooNA1+JLe/ry6tLKwV8/Kp9MUT0jhOixMNp/Dt95oOdbL4PQO
rkbBKdLzSiGgz6HKVnwfriEFiP+63tOBdVy7+kPtIVqylgusWcXYnsRfDTC8
qvh5Um0uzXIBwaucqmtaN/ZHjW1QlF+UYuwG4IM+LORQX87KR1WOfEdAfV71
C+7Xe17E3YBbsDZMpMJhrOAeDQcplolFv2cXhfzi4PH+feEtMD4fzlieo8jv
RMV5lFirC2EnIqjCfnM+KAq4qShgI1wwuokc6DYHIIfLguuJZo3mVKVBLVIs
LAVEGcHPg9m2mxLuMbA/Bt4Nxt4us7/dw9428uRSuPWBJJ/qLVaUoHhjsBrM
MTdhK9hf9f0ebzEJ8NuhrM0u/2V+s76jr4sOk8NoSMJqhd5Fa9T6Fb5UEaRM
wIRq1IKK3IE/yowbEfQnuZFN4mBtSbtmMA3acWAsJyffrne8y8MuUcbX96SR
rQQH6K4IH9la2f+1k5G4TrvKWHQNDfRrQn5xy3EH0RiZ9qVtZ+KMBHR74PWo
qHH1QEuHx/zKcAdMVkkURYNQ3kKL7K6Hv2RQbcB7vX9m/sF5oEYtP+Ase/ey
H058b6z3dhHZ5BAvVP+uubMhZBQHK4illNrIZJuYx5nGcTvJ/IodQb4tdBGM
dzaX4MWQBEcwQYsp5r58Jfqhuwe3hLzBKTz/AcMCXUCu2BkMvw+jP4IKMqKr
OfxI+S6H8XpkBzR4iJt0raGJBMXD1JcH8S5WYSpfC1GU0/QkkFsh1g9uwuur
DW7cN0FffaOfxmbgJ8j9VLcy8oHpllMcgI9xMUfbIZ2U7zHvoyvfpzhm29lp
uwlOx1DBVNRH0MOuvtb/Dd0MLunATSFIR1jmPVybATP+fA4lIe+IZZOV1BJJ
JhPgheyfV8F+8Jta1ObgIGbF9W7kyctS6NL52AFmo5rq4vpkb7NUbixHU8u4
94FOlsT2TPv9Pg5GP8Hu0s3OATtFRK/XbxRgm+/73rpzrKrP7FrnoT5tmKbx
H/sLf9axMLZpIw+nCtIPsOmqQae+JIKTsfR0VfOuWCpSuGyjATGVUdABIuAZ
Cs9wdLsJ3jqkFFASVlWvxTYsUVB4pMqiYeXmV0DFcQ3K/2Ei9fUOGDj63NtU
ruUC5BmP+NBecq/qUJoJAilb5kozKmy+5bZpMxC6RoslUG8pFFa/41SQFloD
7Grh++BSM/hCeIiv6/waGpjeM9HxPVowYuV3S0/HIUs2+29mEAgata0c9C4d
7vvz42WFIFyKtBkgpzHjavM5IkCpJEtM7qfUSx3nLknlbVwaUctGn1vBlpQB
/YuTVs1XhG2TT7/cFwjzghqBut8PrkZWWuqiKPZkOsWpTuzcFyO7xYDZhVxK
dUmOSBzFq/dB/62D5F+CAOf8HCUlJxtBSqRAKYYnX6ZbRMZTj1hfafyNOg8Z
duuq6TwqpqelHijHJi00nR93fNeiKub9ltO0r8SubYfvteqjpuDcxKc8LpSG
8eNggoFD2K6whgw+14IUi+22WEsx8mOYaJpVaiLskS9YM9CVdIHdAETy6DRR
4d9tuB9WExycLZj+IqzGi7mywfZ4aezNjODHQft1A6SoZenZtwgOjvvAsVEZ
okStIzoiotLTiQ3b1DFHpzsZ/wCExxFcGaB5NouYnh95BDfrUT2CDDEjr5du
Td05JnWChv0aDHNmKC5zRFqGjcACS+gUoJyeH9g0Yi6CEZuGidTvqw4mpfss
/04Z7gSPGfOtiUJf6jDLm2sPJE2mc3DDQEtyHf9a9c8Gbhfdg+IiR8xb/Jsx
F0yKno5GzQKQlujxXkQeoXL72Wbq448EeRXRjVLIdYGJzFhcCd1U8/J05Qlx
B+YDsmXPyuyMfG/83J706nh1D7QMo+xiXt8n9L3jcL7XpBdOWa9R5FGPXZgS
9y00ZvNZ2J0aa2cXj+sEe78ZyaqXWyOyKicJygew3iKteVUasbRMxFF+HA7J
iMcjX8FowOK5hczD0wZza7RbnQS1iEc5w8zWSNKdUsmhAQYqaz42AP8Pzvn4
D8yD3C+QaN2EjLByrmsPy/vKuHIq0SaRbQkdnJmQWw//wKxRqiATY+STEeGs
YvijiYAjIh4KLmcGyfKhivrwYtA4cSNH9tv9a4TFjN4CAH1ufsGhM0gu62Ux
a2XqqfgAmfkJtxTIJw7nMJtMKXLb3TJOmh9Hf32Iz3k52+SgZb+fsVa4oYIX
Z31IB5qF7HortOosFp/gm7hJ/RkBeD33D55L5g3hR6LInF+s/riS8Owt5h5B
2404qOoi8Pf0hKU3skSBY7GS3cPbEMH4Q9bZT1OGLJCXVdM+oh3N/J89Teul
XibG1ngZAl96ekGaddx8xk/Mp+txXVCNQEoR1yxITCIXhr06I7n+iiq7hnfp
AhjqNRfmERKpL6RxxEe/kfSgCIdkTjSpOpVs+3qNRLv14/BD8PvXf1aR0ByW
r4Jydp5+1Z5+ryFxCA+wrLfhfvlG3NBJqoRyCtvGV/x6EoWzS6eVMSphIZ1N
8YQXEPQaiF+BOt4/p0+hoYJ99UEW4Q2ZGs4vc//nSn7kyYltRtn/iI4Onrap
Xv7YDLGIdRPuY/1M40OEWVDlyGpRRIt/Oqykr0No+SQOfpzW914D1TZH5Y+P
3Kl/uUMd+tSmqTr0CZT64vxwlTsXJs+mZZGGYVwzo3ZRD1A3R/AwU7ojETqP
wbrQZCAUGvQg3JfyM5mXiJbRIz/OiDlW3UD0ARyGCxLYZpWkmcrt1+PLfUtU
/pAoMb4EJeZdan1nkRbBXQEHN3HgMRRHYCyhinBcEZYIrSdSxxqqtBz953Hu
kLS7JMCU8bM41v/EFWi1fFKc0L4qyFLyYEo0MlPFZX9QSyErP0pPTtsrD+Ik
1qPm+m/14Ebf3wzOXetptaE4w+uUI4+430ErcwhpV27yJLj4ORMIkXiWKTX5
Th9dmPia1RiuKRYVrHXwHkPupMKa4ts/Vwyw3NzzvUzD1QrrOkzQi/OfucEc
JBO62WlnhDePam2s912R6zzhqUuBjdPa3ydJIP1fa+JSZhyPlyek5uB6XZhx
iOxjPpUqu+uX7no9PMHURz7ce2HJdx9dv3ZKojVrDgnOAT+ClYrmnI3tvIb+
Gc5ylFLYrcikEUaxyOnHSubFGcYY9FrO7vhg0XeI95S/g1j8PxrUTgVuFTd7
UHvVtfS3i+CThCf/4hAYZ+qqLqW9yvfIwEMw9uvsSfRDvmqQk1NodkgVOVcO
QAioPg0d5XIpldFxlZpgwbhUz/j8+SMvgfiftqaKpgMg9A9qGnskGxOl4BRy
5pmsFy+2fIlSRAs9DuUgRzHb6dQ6Vwo1Jwk+HBkUmQ+Z0M3ag03ZjIWtZsrT
FJdI40zBu4H38OUVUN/ukB9EphO9KrxgAfUYaPCa2SFBWJHtuhHlwnwzzkjH
ij48ICnFQLGnv/c2P1snMV155Df5SCD7KTJfDVRZn14+xq8UT91yKbTwvGPW
lFvZH7auVBDdHzqma8+p0kpUtS5n5kIJ3oMh4oTWLysLmYi6mrUD1FYnLUIa
IiStkiwqKi/A8c4nD4n0Ye7pRGeChAAEz/OXnzQ6VZKEf7ma5c26zW812lHS
sTJd5VUv5YZ6LgzMFeQN4dJDE5Zk3gp1FBmKFzsHLxl3+yAP/wtTUcN2sAKv
XDmFdK3QDONfBpe84xCt7uHF2Vf5YOKMGia+JLrwstuSZpuiWyB0Q/ZHwTRv
0jvevYuZDYmtvIu4uDbovsePHqDurf4Ch1b/bupJxEmUTG/7TWPZr2VHNTgs
EkOmvoj88oDF/e8ilwvW7O1h7UtP1+eSjVH7wCA4sDW0kkMzg88GD2L9+ReE
4EsWkGGkUJgWAfkj08m1VyCT/6par4LYqwYf9O2QAGUPY0W1H3aJhj/2cX1B
BlEthAOjBZFT6L5yVtk4X4yO8R+ovkXkRZ//laNTbFLlNuGj7TAugBY6GMzj
lR8xerlQayTbeNqRr8DDsRC6kNEIggzyYkBBDbwiRcwUJNNP6Zu8JhnMy/sQ
9UVIqGHm0DyYE96FjR0hEQjWjEDQ++JGPK00QMWlZnR9PoDB8QjvxSOu55tX
sc/uifrCHt5j/NPB0LEhyGTellDK6H+zgb+kPA1jKl4Wq74CqPXC8k4eyWBy
rC1DHL/A8jG2mbGj7ePYv0yXZmnjGUFS9jky8a8315hl04aPDy95+zqNdBcJ
f1zjIHCMdRY/hYZ3hQ7ATpE6d46kZaL5oU0J0Jsp+Qif3LUN3rsGWKyWAYT8
BcdKPKmuk3EgTD1rxDdEgzM0smBmaio3TTRdfZVI0qlNgE7/ubUGpIBpO9Ja
pJO5unsRCnfUdbBv6KB3yzr2a5OGzX21snmtmJ+3vLViadL2ApPnXjtn2OAv
Ba+nV8x8cxIAkcxSxmKT45GgJZYtiPDwQbwf9lPZFzlj2T8MWKTTGyLIWXjY
jV4ut2PJBepABW6EGvLVq55HXdX1P2eHur81ufMR31/aQu117JlUkMsc0KTW
eCX5gCwAQ2EoRdnoPuXxT9Si1jS4Lo0R7l6XO3k6NNqD7gPmToOFhU+2Ckts
4aOBB9sj0dii5IBF8nmFy3ul7a0lxfV1/N4Zbsx4XdpZ0APY3DgoiE+mdQRz
rgzS5ZFBWgqD58v+FrMuAZkUtd0/3mVma/nNi9eNeF2QXIQhVwSpox7Xyfjz
9GqXGDZFECzeIZ8NEP4nmBGgAobBNPQM1dwGwmUbdEQ4Z+u2DjJfvo9MPpvr
g0RoFrtGfJ4YN7V1JUtZi4G5hWhlUx/tB+sT2TkDP0QV5Q4ElOZcnHugv49h
S+NR1twVLLGpJmPi8S1L1w6nf02jascXh0BA7XSx+jSz7OP0qt3Xol43ZX4d
qPox8+ZLvrVajDSHv+XLBhwEeCsh/SLB3kaw/8MoLfEqItAKzVVRRNiS+Cua
f5LjnRwkJQYOOU70D7DU2o+4XlyL7mkVP6cVFSmvIhRJMFpB8jryEhr5GMjq
pgN0aOT9P6JpuU7Mg8lmfQKpkzhnqUX6RjU2liHgC3YwxHfhOQr11sOxLvRn
CoRZO29+iwNXfekrDET0kYW/OJzfxWaz3XgTfYqbr1/5nYa8Y97R2x/oI8yH
REx1jPEZQE4azjT7JwWpYhjcut2KCBls8D5BVM/g/Es4zjFVKS/UBniPpehk
QEv3xOqVECgZxx0iqFjMaDUEL9nM5VI9gSDbRWmPlkG1YqiJQS3iYQrRzgWp
2Zb9DHawIhn1KhDDKb/A/WYNGmUk/WQGgva8bA7HBgt4HS6oiy06V/Xn08y9
TiJ8EUpgQKbeoFSfWoODKUM6UxY9B/n0FRtT+xs5uHJ0vv1RCpaQ5QXUgnXT
5FWU1jSfmPM6x5y0/iUErMfZhAlzfjoQDq0YAuxavAONnBt8stHgOSV3hplV
DUmSuNYjP3MJmr6pOGc7onzUxYTrFdGl8obeQbuMkL4io+rdxFcc/D2jGnzs
plK49npnK2+41UFcE43hHpyxPfdyhRM8dJsdFeYw/9ZvmMcuj6taJ26eVIX6
NtQNTD2E2IDnnL8BEsjSyQ6JMqgvLWU9NFf4ZpbuuznrvqFFHcH5+Vx4Pu9B
uUZWGZQ+KO/Ku+WuQ8aHphjKpHnrgbZLsGkXScYA6hF8pYMTaLacvAcWdItG
smVgdTsntDz5HhxJA/OPQ3kLtSyoaLHDPP4WmEUYu2VHqMHxRMnvuJ9rX4Bj
bub7N0zBrqt9X3FVLwDQF4VKmWDUZFXdD7ER+MHvR4XoTciC4Wnirgyy/wMs
tPpnAiJvFlapF5Z8CxKQBg+Ylpjvo7zWl3PkMrADqvWqPG1uQHwocn00evd+
6PtLRCaBVBEOpniwrQZMkOEs2p1+D07Omo5dSbYDnUMIju9kP4A+e/jPX41E
CO9pNP4haem8CNmiPHN2Yvg+BzdFLcNRbmvJ2wrq52l3AMMkROIVjJLSsxuX
U5RVYdYhKiBI1+MgqNzZlKK6gFPS9iIyiIx30GcDZT4Vw4SXtEv/fwhKC8Ez
aNzvJozY5mH7FmZEqSlHO2K1UIqi/+NyyULaT4uVauXidhyFWcG3zYJ+68JE
qznP/kHBGTYUQR2FChG8txq471D8UsVhzdx5HcurW6EQ11FznZqcMBckWibt
/559zO9z8WH1JO7VdqDSpvTwEpvWsHh6AWjEFVCns+SEb6B5niLcW+SpUuCO
ywaFsGbEquRQBEX6ZsSsnwpQZkRcuje3ENQC98/w4O5JgWZl6z/UzIdJ5IaC
gW6JtgHblYK522fzEk4XFEYQLzHIfEXEUtsb665t58IjxxRklAF7sC9NDe7E
EWVQGgpB/pYLFQe3fL74nFLIinxyaiZW8KYEQhzv4roBCjbANuFmowTJFn0q
MLBafHIesu/bDPZPuNMra+pMhaKeZxaWiPg7N4ShxSSX76ulO4VZTsa+86D+
G7Du6OkjcpiY3Z+XN4XEKRApLlHGCNIZmsfOOJCa1o1vOSotV2MBEA3xlLod
P1V1gOrXOJgPHiErGpXR7ypj2ThzXJGRiYzg/w1OlbQ+ldP0VZQTiqPhOd6E
/gHWg4DektKenRtvKToG/yr+KVCQG7XcfffraBE/4JCmNqmGhI83URE5ke2D
Kj5aEnuINHZSj8A+IcbSznpLhY2Yzqq+CYSqNr7wQOHx2PyRmCD68YcVLeH0
2uVRg/arW7LcHw+qqVTQP4qaEgADV2CA2cWgwt7R9hDqkyhav0QudlsSNaHT
MjK9jax89Xcx3qx8Xd1MHo0QMNm4xp+ODDOyA4CY9LcsqHIYNopgbNEo+I6T
l/8GtsMBQpYG8cuTvVwvlQap2c9QdiILMSE75E4zp8G5/JaYgI7Hsdq4YDoU
ifJWkYmje8VpjJlkrzEWP9c2RClZ4eVh/s4U5/ZPEpk1sWzF001CPSv5Y6i4
bigIkW+FKz8M4hAeZanTbeQeBtZkL5TvIpbQNQ4vpkYzcDywxMSDpvnIAygr
4n0MjaVe9kSbAf7taKQu213ktOHxBZgaiwilRe2mNbU3P0NrtQobtxw9Oly5
09MD9XXXcYAx/506JgT8zjfvDlvN5YCJUKBlocSbL7jQ7dJsotYwbBTuLzrq
/OB9QAt4ms4quNgFKt7ExpkDToz35/hlR8iAYbqUO2/j9tEoB6e7qVgVUWI8
NLJS6lIGCSTcnxJQHp+thzYKQnVC6mMgzyf3QURdFPZqhXXRexxCPiq6pJg2
o581Wnxuy0MmkiHZTdrNUwy9oKMfAsINA+eTFw0aK9D+PA9sQZ39VtSy5DvT
MOCO3ekuPdO0L88kG8HnJtMAqffkmDgo9h5hzyWyDF6MQRO36pD+A6wdb0hl
VOZTLC1+0A+DeTnjEMJkTEKZmNwX18032zzCUj3izgHqeb31RKcN3ekZiQR0
E3mxT98KEwY+VedxLDtjXv5YUJj6jpGi9py1lcTqe6z47xS1lPUQaHyya5ty
uPTs2cnbUeCkHjoQkN7wL8GBEveMxIQN+7++/OH+Z1D99YcUjma5wdnyNwgo
rmpQbIvVQkE9TcAHyf/x1mqYgSUjIEy+O6U0JUTfv2Z6cwDLvj4RldAfVVMX
DAvP6qb2cRa00OY19gVzw0SdInU51abMgNsToVWX8tJrjTQLE8eRsSOpp8ID
+Ycs8K3qjQ2MvYqEZ85Ofx+No5ZWRcxyrxTFiKl0jFQoBZ9wDFiWz6naqpYo
Wtz35ZPmCNndQKVHjzOM81MH79qmJTooM9jYhgPKR0E0+TphYt5xTmnkz2Sm
ZV8UN/Izj0oNKMFPazWkwJ9Qtzmo465VVknXj/tTuKxpTzLC6/zgccHay1ah
a/oIc5taUFN/pznpbFJg2ZJb4PyNW2X40H5WROdJEcLzFpQGfSUXlWi1Xe3f
hcYtKY7M/cgaH/8wgzdWXzGG0v8UOHQklaoHUp5qVEZ18H119M2Z2oVHdL+g
rrZhEeqxXZr2UYhbRQ7a3QXiS6JGU21AnTS1gVBVB0LYM70EyGY9suxL3KYe
CLP/1WCOEbYMYLGJMrT3kl1Dn1on5RKVim80f+HHS7XyHr/ASN4udXCpU5zB
a6o1/vYi3F3+muX20uVJdcCS9HGCuQn1RlCzhLwpVwa3nvaWF4djPuATXVnV
noisIiFI7k8AvthiJbYpC4F+QRc0G9dhnPKolus7mkU+OdUhWFY71P9Yt2sh
Uj7a2iws17cVR8mVD8L+0vtfvV67qQhOa+j40vODuDRq+qso5QyXy5GzmWdG
4vr8qkkSLa1EWd9oexsCSqS5/yuSt6C8QpLLh1RMA2ix04juvffkDDz98DlH
gyCTpnW1TC5iKR9fsYR31EcVumGHYhsiR1tHWaxRoF+3clUaE1NZLbefGitX
GzDPyYCVRlYE/JgBUG4Fc2cl5ecnNrjCzvq8LRnCd5vM2chjjAOnHrNgyZvJ
OvPb8qDJ7xe/jc34kLjMl46G6I7lB9nR/dzM2XbEVT8+eqjmu/cQ8dEc0eUd
MmLDyKCym6fE7Cz3/Y28PTKEQkv2Bzikdn+qdXnkSgCwGb0XNFP4lCBV3K+W
SkF8tG+aOJAz2RdHWTLJALDijKHrKUx2QzlF+NPcAEGX2E/ZEsuRShYkLu8Y
T5n10hJFvcmKW3wlaH64p3zkIjy+43aEs+bCJVShvElu0Rs43sCsPSN3QAJs
bcvC0k7dzyXnPf4O9fiY9twdXj3dxJu5EkUbtjHEJJwqNxHzcS6ujYsjDScP
En/hKEXnjjB/9j5rrtnmM9ay2O6CDrNQzQojqyWzyBoMVxMU0uU2/1avDGag
mu8F3w07JO16KH3fuZzZGYiKO+GZphNvXhcna7eDXJkdLHfz3dTyBdwWf36s
w7DuAhblE39F1PmZETaeafFqUei34VfrRMYfQDpH1MW2VEF6Yub4J8fXA7b+
K5PCwsVIvqq3KzlM99EBohUjl0O/BGYmkaWxu+5baK0Pdvp/9IYBK70R8Qsc
pfF/z8KuNccCxOoHAt8FBoZ9GJeotpxswdCZE66Fscv5DohbO4gwEX1Gb8AV
nleAN0ZmI7Vx4dVQWDNlSJPJG1+DBGMS0ieaMmEv4ZtT0zvGK8+5sRS7IYSk
3xr7bIjjDPi6O3cexcmZGz7t0MvzQcU37AWr984F0MKN4/tFHQzUk7gDqQ8x
DNSGnTwQ/sSsPFYLdprxp7mDhOo1i4qwSeSejf/XsBqkSmSZVcmSJHXv0Ygq
8S6SWz8hN//VrA7Zl4VFajo1QTjUyt6vbtD9RfvfjYdcfGDDw6tQoAcMBEVc
1YXemOW9Kaho7bpRBMjTzPQDt3K+89SrgLvOY3RxGJyScMkjNQIkBiDxuqkk
/ZaFzQjqcxnFgLahHJSwu8LL5YH88a/nppszemUkAy6SS+x5fGJQRttjGvnq
U3j2qfREVjBmKva6Hvrzva3tLVggo1LEj+W03lfMtHY6AHv5HlObCKjHZxgL
91lwuHMMXXn3YIh8a1eYxRSMlzIGWXuLXHuCZTwS8w9J90ixoYJHEV5iK8DL
dsNk1iRpIkPPmPy/Dx+e4QaZui7Cmqz7x4j92KbR5BJimevEvnRCnEeYzIXh
c/C4lxLwP9EPuC/8I3BkC3Skpv8x/sVX1FEvEKQDwl56JP3zBTkGFk7BL7xe
x2V0CuJLc9ebh0enwTQhUhUtcJaTXdC/j20EBqUM86vs0DOl6GR40raaHb/D
/fXGIr1VAoBGHM6COIMptuPBmwcZPjcJ41kJqtFXyaDhjUHWpl08mbNEXOpE
nFjvA2YCOS4+pkTTCIukY9ifSZ1F/5IHjQB9ByViaeAknliikA/Hl96ooy6B
ehBOpZVXBRHJNxmajdfW/Czc6CvkHoFi2iPXvSqq40QarYYoUUjVMKafYo6F
jkJiPIYV3gp8bV2w59NEGa+PnbltxVO4gy1X0kzw3GwJYwspQH0BoRGyeceE
viwXoeq8Xz+8rUkcRj1KDSZR875dAOrmKpZbxJL5joOS8fDjSwkBt3FFFK5I
0IDLsfoPuzCU1V8lMTn1Q8CV+nZl/SvuauIuKhe4IjIZGOn2fdnNjqhtdpzj
45ZcGOdvC7U02r6QvDJ1rTu1b6iHyPMWpH2U3pBBX/+zrt8dyOZUn4tcK/t+
i9ijOPksSPuH1xeKZc4TouE5erCc5HN4Rkf1WGX/wkaoA2hWPK/pb9v7sQq2
hQ0sVCK1lIZoENasNqlhpSlH6qAV7pg7Q7MMH9ckb/oP/RYFj0jjYSjSdkL+
tfAgHQVv8zXI85pZG5ttfzsO9dLX7FIPNiuOh0AoOphLWbK2vEc01GWueyhJ
XCMuTCj9IGM7TPvBqCLPyAVaBBgxM9zmwFiJovNXE7IL513wNTRL9fa5bmv2
7HDAuGQsnEm+wtuUP63qLBhRsTQnL/wJyJb45EQr2Jw7W5q8wp9y1QVya3XS
OV/dfuc5w8UcbGYQksbqpEjliS27FTsyB8nzMB43lULX4kl0Nb7mMP9366Tr
nUvwus17aCs0W0xOG8AURRLzo5tqiETWMC7luYpH/oXGmLSyvTK2m+zt85pw
A06RJAL6+uu2PspkMsa8lpMg9bWqEpQyjw1DPFijYkTwYuzy0Y/DnHM+rYzH
zItpAQaXWA8QqVBhZcRyN6u/TOmlYtg1QJGFbbSBSLSEqw+FlD6qjV5LHkMD
/J17QOdQ86VfqmL9vCvYuUN70F0dwm2ub0cyTedKcGefKlj3MAZVJfGYPb+M
BpFB3ElH8RrQlSvbMxFwsrRdcLbepFYwZ78hsecITdnB2ZytFC4RxZy2E0FW
8H98uYrGgNETpftAS76Yoc8s64gmEoqsJ9CF0VTpLTvQXZjYS7a9IAbMXGHW
3aLtVTdCuBJzHsgRdDL6xD4aVRCB/8iHlpnlx6XSmbEsxYDvG8R29gEjeIik
2nZYfkmrojObWwNAZE+Nu7ct08eRR1Pl9WrMdOIbShWkqdcZouEBmQtBwClr
CsovV3v9up9zcZqCNyqguHAW/R3lNx3AbxEa4JIpzG4iUPeLfK6oBPTx6LtI
ru2iKDGFPSAvrLqJEgND5KkSfawre/DdKCeCido820VBf1FarJNgcRoEundC
scehxSqMwfYQ0H4br2myg8IkMJ5bpLUBk0x7f7Tw0hCrLp5Nk6PB1QEhdyuh
CPY1yi4tMQ9cznOYMpMK5UyXl62jWOXUguarE4bwyH97Kx+aYQnqxJYcbzio
6NsuFfHYUKocqqHx80sGWCbZ3KR9GkyYTX9xBNcdmCX+6mJrA359ygdQmxAf
Kl82jz1K/UgmqBVdcP/D3T7r6UJhxtP7+YqkFQAfUN8r5z1t30YUJ7l5vC11
2dGLqQi+N66yVmo2myvL/96o0D55oEv1OikIVVgia5CxwmTi8FuESPF7Dn67
fFuh8PF1nFm6SaqbidrsXh4hWasOIXKGEBpJe5SD9JZRffrvrdndLfH+wdxt
fNDykvP9+SUqVqAWWO3i56SrGjfxrFNlAViHbG2QNYg26ku3tYrE8es+S5V8
DuVp+4ID3UT9LUsUiitDIjpmy5MIAsiMGCQj1NosxXwroVetdbj/ci0at/nX
2hErqviAabzge2V/HFUCgxBCw9PmPJ65BYJAOeKUbTgLD2H2ph9Vnf32Ycwl
oDViWTRFfuvGTcO9EN3qdIDciEePRS+aF/2BZdmc96+OheCUHbAOxmLlGV0d
ejFAFG0/8mZIVD59OOoWhI2JPdQRqZhpfJ5TmD7KhPWzcPucTQhxd2ytUoLq
gyQ8vVHozA4O017ruiD2d5YAWbtDx0YNHFp/afFUPGYGnCI8UaHBJST3mm88
Y3VT+AxtaC6Z6jRTZah9+J1kk5rUhFHeQ8f1tyWJlb8uRm1JFC8cKBQxDlUo
aKmx0kGDhEwnpXfuGztGIbKYiSvFh3dNDraiRkTTvfKdOw9+0wbVkhaI9REs
uY3Xxmg9h5sprrC0yhszISti8iiciEER3iA7ODa6JvAPH06+sd+HrA1CRjMS
l0Bh7CI64UN/kJ0KprO57OfMRdX0qpsyQpHklLF5PXVtRWgLHI1ckVbNlqxx
WXKuPmLwkXJPvp3amIx6z+RuvX5dlRf8h2bp5IAuZqc2ykkHmtDV2wZ6Cs/X
cpBFg7zp2dr2DUAD0FeL/cy9kKlij1M6WMkDAj1nrfyVirxkUzBgEg4P/FR0
ebEQ4R+OlVFDMG7Ym7I0SB6Yfow9X5KLrTA4OIozV7EJ6O2MEbYJkNUn+0nC
FWRn7VGQlL2ih9ThSgp9sR+NhAyI4sS8mrIJYILiiK+BK1QhMCu8lijouEtk
rd74IC8dGndVhN4D5ZHY7Dwfgqx1Vj8TE3NG4EC0JaUNKpdktgNKiOCQT0pY
l9gubBfN7OBJe4kKbSWOFfWl1qvGGifm5V+FiUE4a7GoOuKd2fLCnqY7LWvy
Ri/LmL5oOGQ2ylebfUnNB7hSY3XnbCnYb87Dtlvd5Xl8gnY/GlOX51ChrW1Z
ncIGSWl9Ce0pPO3XZHbsBmDhomxZO24BnSY3DFAV9oFsUXdhgyczVNhTf/Oa
jvg9F1FyqSO0gJU0TwLPiCVNjbKS0BE0qn+A2TTFVkMewEaGHPCtJTNTj5z9
elHQSFh2SIzN7RcURhuJUF6EtjYV3XxEpHX4gu8xyBaabOA2hRdYluBtqdFF
Yct8kjhQpSWhqsZ5BiTUetKsfokPOtP1ZOoXZKIHlExaL9kqGTXm/YEdWMAB
YD1my8Ew9ztD6QqSYn3LkAlvz4gnmisTfdNKOB9h9U88DrfT6ZeoLpyKGWqF
qJhtOstge39WOUY1j3u98lwXwY1f/DnuV+v3zZsNe3ZYmCoTMkaiR29HY38v
xGWbsh4yAU/TbMKwJHEYeEGhF1yBhTJbH+vbsAiveW5J9K+gbqrytYSLF4Kd
HFicQoYcLuGBpbva/qzuNlaQwOmuV7ifbDkLYmglWpUy1ImM8PUojsHRIBP5
mwDHMpieI1R7tWTZ2UpdvAO4KGNmfiuo1NoJ2h77s9MVBt1YxnczLcW9NqHq
30MIN/2Y46rqTg6oiriYuIGUZgTewsq7qSX25yC8ifLZzDkLM/JNbhxraIKY
qN7p8myjMg1wxMK0v99oFWSc9xozOqqMB4YV0elL4FnIn41KgI5NkXgvgkwU
gm4J33dEFHR92iNxK7MQNBC9Dgr22zCjJzhjJmLlnqsE6HGDmHkxdfhQLS5Y
ujaiuoyBQ8sgvKDMX3bcLipObeK63fsbpjZH6OTpHDIvJn66Kmm9eSvZbTwJ
btfiR5sH5c9AP5P/8clzDPIUdH3vLsqt6Vyvw576H30/7UtMIePF7baByqe2
Ot4AdxqTIzq1JIR1kaEG+Dxlm2mgjiDmwjPC+Vn0Z0mjKguON+30tnQ/pVdv
aotSRxT0x8HZkhYxpiRI8N1IZrAL4RclRXIak36NPSI5kbWh5GH6znEWN0A0
4Dl8sWHINyWsh7TXoI9dwjsZ1itoXysVFOEyhT4KOXB44jS35UOVJsiLTe57
EEx0QriBsxydyzxcbHY60PToTI/2+mtZWe4BRuqPK6XSjA/rLeyWBNkqsH0Z
/1oaSaMhoRIoWztH0hT1bsQBjI5AprC9isroNu6X/SKvTV6DljMEJGtVTMh6
uTyiJQCGqY6EZRJANCxn7VtO8Ab+znr5swYHzXwPZMO9K/JnIdia9HnctohF
xSv8pPgByfIhHm2AptOSruXX/NCtdGD1ynO9eUzU46WQQsbzRePDnnc+Pknt
C4ta7j62FngWxIoon5R4B5EsKkEDRy+r8tmjuiZzcVsHJykI6Mt6r3kJbAKC
P52An/zZi/r0/7L3WN9JubT+DfY4KO68waBwUEcdZUKcF+i7xApWpX90QKvG
PjFdJMs4IVDfC3quFgpAJyV637R1n9uo9Okl72qdT3Ae6C+LgvsGM+PqLQBy
lby0GAXPdnNqx3PTQ+0uV38n32ZhdEEmTTY8peCQztwARVkpgrDe4SZljTbC
K0A+TuX+6vxuiXsHxT7mf6h0j1ZgGF+vizYV0/quSJAEttlDI/LyiSm/vSAB
H45qrkZMoie9YY4SKEpAjL+E2qhl2Is0bk0Uk0xAGwREhKiPFUQaUSUu1ZZs
3p5Y2CrKpPM1E4dUUnTDC1eZLU5LMaVDfzD9GIf56/bn/Tbhyhq2+UZwY2aI
0iz0TsnELGd305Ki4S16+XCAOe04LTBwQrw22B/pfx16JvXFlDUokp8rxuJl
MZLU0NiJ2xSgycrDuvU5GuSKhvAW8v/rMXxWS+NI79JZx3UqQxva9FTXwedA
atn7NbYN0qdtxkuZp0EEaJ3HpxXHRT/ubMliYQwydBSFLgfSeANjO1zKK41P
86a1ak3VG/ejB/hrJRgwwDW3STckpCT2JlN2Uc5lN44GuZOpe88wSkKvnPi2
XDPViT6ACZTdrYh5D3HEup1+sDUsNZuOZP5PS0wt7kmoHzVlT+malXF7kfSS
J1xvrRbNmWDMCZlVwfDOH4FZMhT6JKqDH+IE6/aqcGeqbgF5R6GY1DGCOoWc
05Oh2Qu7p6r6EbCqw4aXRyCOQCwfFOHZZ0W/Z2QtavscjqZDjAKBWd3cWKsp
SepjuJc/IDTojgSTVDH5s6Az6hmdakYgnjtppP1o7XM1fgXk1udDm6F0esFS
+IvWA1Jxb2W8Gpm7TV2WiJN1BsaR3XK+LaZekiWonX6JIjNcChen1SYiFTwe
lQODzWtED6DetjKulOll97DdxIn/pe4D63utXWL7P6n5YiGioQuGae89/TJY
Frt6E3Stn/FJsfumkjh4EdJvDBMTI+eLjKTYfhh37wxYi2MYywgSXLDfQJCJ
xHc3CZGvkbql+LHepjcNwWlCZk3RF6aRAWsYip5Jm0ZoTbrC27ko52icbhIS
Jo20LKcuOHFs8TE6GmakwOb1rX0Mrh36Epbceu1J+1cMPA7GipeAGhgfH+Qr
vtRBE4b8Qrl2pkFL5AaqeP4D/k1CVBAW46se+bDpCDw6AqVJpoZsbb/7McNz
+GlKPh1uFN9yJBCkv+f1Orxg8IFktMRudXof7fFZNNNOBTBwOCoQSOXg61VB
XcBlY08kENpyMT6bO2SsCXSBTFQvYxwb25qzl3YLL5KkvFjX51AJQyWMbso9
Du6lKjBLMc+ewJErymIJBxoQKZgTHiwf5BRWUzE1DKuWQMQ/EdY1EoJihVyS
BJM3sBaq+1BgDN5qO4dZd9n81sddwqYTaYctODdVqlvEg+nz023RN861OM/w
MvdTUh29C6vztrtBN6q5QPUDhrmQ2NyuM1G++SbWzv/0osDOIutbvwvByNlL
ibv4EP5XgT56Dc9T7U5KqIMhTceMtp7/zK5B+prQQGYeZsQ3w2GIrexBi8+m
O0xLXt3pnVheFiOadZqI+NcJDtiV3PlTXFeWJcHEcHiDmgEUqqt51PFdVdZx
7UiHceOZ05bEWxBkWLZRVwLpYcRZumzYO6JWw6abDiqjirW2/9liHf2Dx7ZX
meUyRX9R4sjLhnQwhXZtsCSsScw7hyak3S0FAZu7RSY6aW6deOFqLAz2hecn
sV6WIQGNvfDbrMht5dkbrl4kDE1rcFyyQNIE03Rvq9N04MBDow0SOY4nOWX7
0iJo9pgiXLzOFrvDOrTTKZ6ShNXUhQDJnJXOFue9+WUvqQSUGpwIJtHvO++X
EIeoLwPvsDHU5vMe6AmD2b/6UU9H2dfweKvPklzE0/BQtFkQZzOZeuiaR0dZ
/BbCGNiR6lE6yu4uin1J/W/TFalAaO4W0+x7JmsZE0RoBplndYXlFKCQbjLq
NOVtW00PHxu64WHqkn7mqZgQJtqXIftyJ/FgKWItfaSntRuFYe7Tl6d80Tld
ivFfE28SLuM7SiLnnZ/mZAlrU2a8qe9OBBDeCF3T8W6tWV6nqNjeR6wQA7iF
VBMKxVTBMxR5w5zVP/8D0ifGWVMKLB17qp0OkzvLBQTyw6XfmpxFc0T9GVdo
xXp9G2rd/XFfD332/rr6p6t05S1YIY/wuI9cTRZkVjg803Q4KzT5dCWpLMTF
VFwSBGSxO9/8sPKOPvgFqab0vTDx3AaMw0Tx67z1k/wvw5u8K29dHOetSSCu
Sk2I8+sDuimnZwd6MVo4eHr0O54Qi013Aa1+ae4+eIlkRZoW0IQcqrq/VryF
aoEWcGrvBbAobeweIxryzqHSD1TiY2yBTWW+aX6qwb/pa/LgosjAtT7VyBQf
GIo0dReEIzNOWu45dPkdl8fm9eggR9khVPrqQO5JBtqkyt5a4Ql97ZMmjw3b
3WdIXKIIzdqKU9fA1r+u0eND4lcGEXdolnnIWRdiCFiGivaGJnok2uAHlPmt
FhxSxnOqaSarFxzdO77BWR2irLuZLOo6HnqJI6d+fYcDp0eb8kEu2vXuJlYD
7qK80DohJ7B3GZC9RUJjyubprTuWqpDmltR1OuKk/rqZlPCWc9kW1CZgGKif
b5bhPsieUlWnqVCy+CqxzkpBUNCABF7cZUuBPXlYyxwY9FQNPXH+GrR2ikpc
uhKS17RrzCbrKGk9OQdvNRlPZocd2WiUVN0rMSNvuakScgvbVhi37nyuCf1b
zh40kU/rjc4SbDEdL8xETDXP2ZfO+CCPC6dz7Sb8TTd2AIaPTbx96o/tk21H
QfhcH7DIxVFhX0ZV87z8REk3S8EjU8iYqYrDKObt/5z/SlYaL/ChOG6xhVND
JIdbkwWh+DqXPdvKMd/HemCH7I21zXY5J930M4rg79PwAaLhHeKcsUAqa808
QtZDwPt+oSstYO4oFsuYPOVUKURjzKtmUTA/0BURvNH14X7UkrHzmvp/2Mvn
uSx/35yg8Kq2fATdWAHx+KQS+WcA9lonGxqvCoIASRFBbTj//tgwcQSm9oUv
cKd6oBnYAb1qt1L6psFKuPMuoF34HV5c9k/QABydvf1LKwsDCkNOQm9yZHQ1
XPmmc6zyw1YLuDOAbqIvogT3ooct0kLGbJM4oxVSdSKRMyz6rJuMo9AfF5i0
PccRb8czHc9paHwCp34pZy1bpGHIkKbnX9YXUhUD2Yl1ZzcHMWuUs2qPEbKe
9pX3MQqF6+knyExfmzzZXgD9p3dcB01z7u9DS1TtjDI+EMRYLUkPYAkaoxY5
gK/hjv9VtQGlel3+yGLR6GgMGCnU1/OsTDmkpFPkvmdji4rBAmEFzcTT4PHr
xN3VYSpq2gzs3Y/7F1Ohda/BCO0cfeZBe+GYQqkdG555MUIyZCtsR0kWhBgy
zgNZd6w+6RtXqw5OuJir89SUy0aP7VlLvDe38EfnVweaO/nPPTV1gH6XbKyv
yIBps/pVr2yPYcA/Au5wzyLMlnQA5Ruuc0x4Y1up3zyCbCDbRUHPX/fLE6nf
6lWVLKa39dwJmNAZjU37yT1CzNjwNyZ+VhsnmPwTaoAnTsosNRNdzWEUzsTd
knhUhOEq7aqudgIqQ0Q1OFoDzR2vjuN92e0IyhJ3vE/fLiNHiDth0i+8rHav
W69hqK05VJKIQSEDAUnxfaSRIYLSuZ/Q/H4ZKoTQnwcQ53qTFfqyZEFEqIhK
kZ9JYg0ljh1SOZ3WdPBeqo0FzCAm+uRanNSJER0M/1djGmldM7mMJXMTLqqh
4HbAdK6Njc2C5rXmwC9+yNjgo6LZl62rOvRWSBNv1CEJ51r2+fT3NUhv8/ta
p0bjdeHsmzUh0Vad9qNGa+Fu35Cp6TK/Oqv8JP6LT8hTHJlkqddRKDi+EHEc
FReyMP8w2VKxmXNt+w8TJ4O9EHphm1Xnp7fk5eouLtdO8aNjo0sOanNY2eXF
tXjO3gq+z4rvZ1BIjhzCy5cM3XZUx85MjwYCWI2hnAFeVKR7Aawq+uRKyHps
PqoblN8nRd8hjOfC0t424vc6azPiVSPcBLSBK8M112qypvhZzXTYI+EO8IXA
/gx7wNpC7OU4fys17oEeds+IPjMxmH6SMBgqtcAAmK3JJmkYPW8Vfl4EzLw7
d0djSm89fkIzgOgS4I8r3tyKxCih6Ie4LgV1aAQm8wosDbduYqYP/U06G/z6
yGWdPVzc9fhQqIXdXyOrVNiXA7924v4jigzHH0f0fDL2m/aj1USzPNDCpnWC
O99UBpyS0ATbE8h42CRadF8lPZrku9aT/L859dU385mErMlBQTbg3LDy4rZm
aITUsHWQzqZo5SlPVCn0i13s6D2IsaWwIQztsvw2tnZ3BN3QIgAx8fEt6LcK
6TAZwzMjaRsuH6ADKQjJtQTzbVsmc+04Ti8Xg0g1Y2PD1H4xeU5PvAUSFWp8
3a5QjMuaHhFBlwXxAtfWQK00Yxz75WOkBrq7fq3qzt3ThUgwaVQyg4niyVKs
1OdobpdjOSfzMdjVVKLGao2yarm9/vXvzdD/SVQ3PahRu5EYebnidFDiuHkg
MGe8SWxLOy+P0s23iQDZUxIS/o+EjhfxDAHCGH1OHe8ub8Q08Tjm1wzg2K2o
PgRVVoEhgQ/Y51l6C5bjVYXhyvLrZVsAa1yFpzfqnTNDJ1Qq+qopddqdu5jW
X5YlexGD1xQwSvozJu0/+SJWFXv5sqj/eohk5sgmG7vRglyPIbX1k+Xdc2si
JuS44Jvxg/ykHUnKRatog0WfhkRKR61xWtDR6h7hSMMDWl73gSdycaivziTP
UKMDqmL+eVd22MuStHtqRQMOmjmSHi14+smQ3Ae3C2ikk/LIfu32rJg7huu2
HG46E4kmYvZGJxiXo5kHsfqqpzVwgX8WT19jbTEwDkdhfmivl+T3WGf2+vSB
4zv3E7QGM1CaMoqkJLA2fLlrp2ZQTPLYoeFDGngGKGP93hNyIeu3iY7bqHcT
CS5LkQ40EJnGd9v5yT9E0dZyDjth2WrEIvGZEfmMGcYAHEF410NNzuwOPAHC
yGGWYOZbIgnxfydWpsSUG0ewhNGBpXUZZr+VsbZVCIyE9tdnZ218CyUL9U+Y
x9RtAva7PHzlGxfFMeR19Ktm20BTD/q+q1jpk+Av5ksjNp5VdSo6dBLgofna
Fg2+LB7Wgzs4GyK44Cph5tF0EJCgM6Ex30GwDeR7VaDmOcNmn0AA+c7W4A03
7uJbYeNw9ew6t3RjjZ4SknfxGzkk8+TjE3zXaZlzUrpFj8+xHrFLv794iUwv
cqXKNnyX5jGXir4Lx91oMiIFaFgPNvqnaCxslDfAUpqoEaTVp8BuCXV4zx2s
K+TGjM8fz/40Cce3yA6NiVu77R3CIIQl9G5oMrm+e8Xqk4Lw6/RDwdCISKwQ
QVea2IuTtEb8LKTiStDMqyk0w32f9EHaDN7W2KaV1tJec6+g8sOmmujE/GPq
RpvgWQUivYa5AIbSHksJ0SGrfgctb9kPH3kJ913WPLE3QbDqNGk9E6k3xW+a
spXR7+Pvj2++/zCyokBwjJyvRpro7H1C4u48eD54aoSBme4SfkWPHkIa87Wq
cyspEKWqkPecTf9MpsIcGR7CrSgAbmIbbyLwC99gAw/ARFOwA/JUsk1LsBiI
YTGODFJB3et7dpkwWvwvdmxVNapFWdBTb6MyeXFzOZd4RC394QsnsFiVXEq+
q2fdvJq21tMyq1hG8kJTnCvXPa1qijQhhLfBTWzDQ03YtupCVaUdsAsVyCFg
Wu0MtEnMbvUSouxSbDWSzH7zDDFQm8oO/opn0nvvtDs7lvu8ILTxAoxjxGcf
+C12CFsZPW1Xd2t4ikln/AExnq9zK1l36VuaZHoCJVnYnEAgwF/DVywfsXUo
WoEE/DlGBW+vQvCOqqPkcR5uNUpnVygu8P7qKbWE5W3fQn1ud4uiY2W1GFZ9
OQEU3s4c7DoGjOCoDc1wii9ObyYwWxvnU1yc144YGjXzERAXvCUcYrNmnJrt
52KnLiLwNgaROauhhn1E32jqAZUL4TEtmV/OCNIkJ2+PnUnaMdUetI2uxXu6
X7R5XIFYAXX8+hT67a6F0+4ywk2VnS2wgduB9hYmA1fahpnscTYqvQJhsxc5
TgoUpolao3eIm9DteNY12QcoLQoFx8WrrpTBQN+O3XbbJd/FSU/p2d/5Aofg
shmn3XG2yx6y8DSv5OEtDnJGZQnWdSBef9mA7lObO+TzHvG8wOe5H3WYDIdY
XxBYxgtES7X4IVhHM0dAaSExh7Z2S6VqJrsuJbA++L66HTiZWNxzFN1GeORr
5lWpneKKgppASu1Pfv6F9+D4SzXYVbEhzKDoN4JCNLESTrj+4EJgJ4BqFvMc
LqsRZ+3MeX9kkzwnLoJ84hqGAcLmwFi/XvxW1B2995alUAWGTWTEG0UB7nNZ
Z909/wkd+/Fmj7P9tLcZJHM9MMBwGtAd/fy8225Nx33d6QjkStDmJ6hwBtHF
wnZfDIfjq3DXlYF4zFZXJEF8WXmym5fkyPWsjeFDg1O3HJcCNgCW/IxVHv7i
3Q7W3vMcicMoXiN6TNwGTKsFyaR3BPOB9D1F6W+w3tYxAXDQv0F4SF+bKJy/
W0ybIxLkp26jn54/RTD3pNDlXpZW0FdUW9o6mD7LIN3jdHssRrPSWQUIUWvO
PY6ggnQjPGf5pkFLGJmoeghb5hC2dBpIM+M6hC7uYGC/LrhZJZtDdIcK11x0
SRhavgjFAYb1tKBEw5cOy4a8pM+BNCkQB1KIK2n8203Sff/49w9xpeYGy5WI
s2m1RtoSD5ieZ63UT0xFVbE4sIMOsMsHa7048XdUjodSIqt/LPUjLzhvYSVP
3VOIukVSj44BGz1/d2GqRbdMnFNb+beUfl14zc43s3S/uQTELoj3WFONK/TV
9P8DPyHhq6Q1IEt2VB9yOrFE6zExPjrI52GQluhlNrB8hX2Qx641BSP4XiU+
nQyibCPJ23lQY6pAIijLBjTOQ9Ppd6NbV3ZCX22JE+ZC9ynH+Fs/8CXdGGed
FSgxREBB0JRXiBcxRYKRVhdKJwVLUpmMlU/puL2d5xzmJ/JA8m6VWMzEp+ou
MNK8K8f4+I/mknPi2swt+K5+WzBiblTSGK1fC2E6CuICGvthnfRsIM/n2i7Y
saFpPcCjQm8uAEvyzR8VzRymST95BNDPHrxkbd+3Nue0j/BAWMUjngNz+ZXJ
jNErPoaEk7f1aJ2ssN+4phOnoNaba1S/iisS38L8mmHQ9iAmCbmmu7kt+bMF
E4Un7eAYPOmItOjW0ubnGylYqr8vf3SwStCRMJ7gdSTIiqIunzGTNb7XbSsu
SoSAA4+Lii0eaM8i+sHng+wUyvEbOPpSXnIqUPATfPgP3xVlasqlPrVKrfa/
AhoTVjkHrCSUDaOVHHBJIXpZfccbRfg3l1x3XCBmTB9nMrZUE8+JQtoR5DPM
kO66EVQ6q9Yplflzk/wGOCKjgEGBTbNOZq3A5gPpf9kGRXrIwYglhEoYXzvk
PpHXdzRz45gQAOGFcRd1UXzeNSdkVZKsmzeVisB2yJSdg8Qmxgo+5yUqjs7X
AWRctMKf5Q9iH9Bf46IrGUwLoQ49k1F6W5OoZRavqTiOFOyLa51TXQLIMIM6
wuUgpsiCCtK4A8EgnP1n8mNFy9SgogGXkc2hAMyZIrJdm2uCv6OKiembWUmC
yw/zbxXQ/s7IJqTWFwnvnOzKGjV5ilN0FjNybEcoBtDGhfyRlmUUSG62aMzB
7xLO9KZ1gIIedfvJQzLCbnPnUK+5BS5e/+a6sM8lyjFAlz/MJqXdhjHPQb1j
rXL0b6LlpPkkNbPvt5oeGE78KJghAIv+PTf7DW2oDXglZPEOPIpx9ylkdJcg
Wu9UCP16ID5L5kIu7NEF9X1XPaQEamCn8V/z+EYTlpS2IyVcZM3xu5D/KgIp
Nyhzjd1uqdRdGe5Mn/dbOP+bPOy/bMVgRc+QHjkbyt8q82D9oIIYfUcpFSNV
NzGDLlS/AMB3M/CKwboSXttgyvkTo740uaOK0lwZynnHN5sW6mMeAycAiQpn
Zizp7b3G6R7N9Snu+5EQnMmj6hJX/voaHJEcnh76rvYVhSSKJt0EM+5n1tI/
whkwoY3vHK87miA+yzI7lgCxs/1QrSarUzvRISxxGOUDA29kt1rq4WZpet36
ObfBA3kJ3YJnLRg6cjqQI4Tq9PDT1ND0M+vDjEcd7z9Sr51Aoc7+vh8X28Ie
gD6P3nGiie6Urm43bw2Rm8KsUtW7sV5gCkZI/X8d7m1qqapIviE83tkUQI2L
nNbrzVwT3n6JFgo/LFL1VJR0+xlV5Q8oFxZ0QE8e1ZZYv5xheFs8quRvQp6B
TqgrIElfP3FeNteiub1lL5um+SC0pBWOKxKNuUXOjyFyuj/iL4iZmdMrNv3o
futiHh6GIbQYLlo6sPllLozCgb4G6jfd1CAnSBI5iFMLpZjE8X6lHRQ8+Gm0
qgKBSyZADHkwAEXsYcRj3b4pW4TwFmYYBPq1V1jG9gnno7yyYF3PH137xPSN
qmdKJ8t3qfqTtH7NqcBJA93J74/LUwgNmF8OMgu0C+zNQKrRHPf5ZbEfVVDE
vA+UMb5zhsvazsp3FgtOqze6JKdFwuk/DJzvQYpOAJ0BiaNIo12NNYWW2RMC
Ybh9PRmqFoGCt2BVjBqZ0GRfBkzI6twqKiQI8FrXEnwnjumxnBMHu0viJj1U
1rbWD2JZu36Lw6PD5HL7efqBGLb+SF/NdQg1Ik/GrbzxzstiRT/83rtPqV1L
uPp0JcU6wlStnO6HQ1V5iIhCs1/KChxeB+6L08uoxvx+jNRO+CPmlFqtqVrp
FXj8rCYa3PZmtc+XAwHT9artNd2+qb7TRn7uMx2lRWFH3iJEPgPa3g8Xbp9C
pMI6R1wE3WHk+pajiqaZt/wKuN8pUvGwTg1rnERojj93bODpMhg4XovYD05y
EBrhOYnqWqPLCypWqioKuz33wYvXIXOx86be0HBhoxmlZpxdUCK3KKtWxlQo
d8Hult1ouDbwOQf2buhvbw9CeuyAOnSlgkyWB92ZCA6W1repG5ttxeWN9d2G
UKgPifmRd2HOa0XMR/YNmci+a9Nvh4/BhAQ/Z5S06txqQ1XWX+e/znOqm3ih
fxxbe38Ups+hj/LnHIiJE0XiyTBsC2R+Xf7SVMeM0HzQDLYld/b1+XtbJNju
uoi+1YQwAvT3+Hr09fbFTYWmcmdpKN2NzebxIeWqULCKmRGfT/KsWKlf+owp
H/QJJjp/th5arwrIzZKgNUK5Hz+6ukw7L4egNZ2CvYXw/pC8eTC1E5yF9XiR
odvXdcXn9ewDBpBpTWV7PtxOXotS0iUVzl5P3Ate6mx0bd14NIMNo4ggCpfU
HxxGbz8qlZ6r+Ck14CIK2Xyh/ZooimI63CGmJEi6H8l2Y4PGi44/dQ3CVUNT
gaPRJuJgDX33Nnukq7XDzsKFYFP1fcNB31Bix/bhtvgtSrIpcorZMOnCYyHt
MhXhOoeMItQ3/zYYAhXODcHBPS+RK5dPVVv/DiOYDrWHmu3pW90wslJWZVwa
WZ9K4qDNcpZlYGxIofaUPyy+FUhC6tsF8qfEpG+L2awIMLzCLdx6BvjbsQ3g
PBsgZP7rBbg6Qp8kE38Oenreh+vSmIRb8JSCVi6ohNFRX/eXDTFWB29xzT4T
7u/WVxPqEcMLEJr02C9zKCxP2S/LPuqoE48oDUZHBYj6OBT+SHX85a1YiyIn
POKURh2c14IF/gVou2Go+x4XFxbNISa9Cmv9x4UxXw7bEyClEw3e7DENds2j
E36Zb4+0hpTZnI4aGauA/XkfX9eI0uDQaopnTTuAycPeNz5iVQWN9Kvqj0J0
agYjcz4tUwxzVmhIDVnqW/IePuef03HbHRfWTKT3oW9i4l5dY5RHUN4F3zMH
vuAFbJpJN+UJodgzZ8rGvQmyXwqMiL3rLsWuwY3hyw80V1TX+5gCnLrwicli
uUfB0yA4+B0e+RDlUrgNe3ILHsI8yrZnjVCSmHnB2gBDVf4Zp7MJ0vkxKil/
CWFpDN1DmEbiU9uGQP/OYWVrPvTnnByl2EKzHRqeGXp7K1Iim6VnGgzL8Byt
+i3Wz+I/P1n9Hvq5qpxHYk/atCkQDmksJm/CfNHoHpeVsNvLWN8pIQ9G69Al
32ip8KAKg7ohe3A2TeTVGvMDAtsNP697TqSK4mP9a10XN5JQ3+u1tz5jQp2L
u4zo82Wo+UkCJMs9Gbc8jHuFjUuLrj9hxGCdmQWuXbBptbaSga8RZ8iH35Q1
MJNJ8BFi65R48lktAFCtYmF2s6ZCO4OJ8/7E1kluxWDUJe+hZQcg1jZeWtm3
cSdZzFacmT7h31j6QWyVEBdMYBzVF4gPYKLIt/N4btCbUB/CjjpOdpcU9/YN
ewmj3N2wadvp/NCluwcyQxRfwiVRMqYz9Jtp3t0jOhmoC2Gyp/dzIvALGo/U
dcdqxmHtyI56Mmw9a5BL2LAF9LJqqbWmKxgMHrWFa9lIojhf7n0PztdoOf6N
fHYRlHnfDUOrhuOE6SNSdSi+Tg/tncu0AAjTDZaO/HmaEKvZ3jRH7iFNuLWS
Vh5WFczb3RYieLtz8tv3MLT6qauEso7jMZirC1VaP65ZcQGdq/+aBB8LohnO
1Rnpm2UttgbBPigu5atvVA4jcsHiOzCfMd8VxK4bOJjHEBrF9GK8DaC5NRFe
hEfjdUCBZLCXTXqKzlQP6qiSKUOijw8eVuWjsOlW0yGyFjt16/5pEFOxAgd/
bIVea9/bBvV5cM+v2tGynd9dS9jln8eCLzjfQLfL7dJyWWlFPcJwRHwyR+xx
+AC0dOGAiKgNmVEB9T3ATtRkMGhnTjitod+JrtFNqf+4JS0yzGtZhEabVp2j
5+YD3p9rPugivRpXeBSI1e6YU7iJXBujxIETyTIM6E7VzF8Zt7YiLrd4oLXq
e8pAMPE8trOFNb9cASZNBBDS9PnH7hSdo1Jn8bcomfmhz+ctBGZorrOoA6LJ
rLdHgadVn32ytO20EUrgiQY8+Wr3DsnM/TA4pHieO1l9NO3uj0VBXasDYp4U
fYX6QYUvwXW75b4upxUTVILr4p/ttjeUJl9eNTeqE1XaUZSNrsE2Y46TjDBX
Br0iSeykVLizo1Cxbz8F8V4YIiJDXmOFN8EK2KMF+LSIQK+hmV7n3KTPD/VI
zq5D/XbxgNH/tyW2r5Fbbaxp2Hh9nJG4oNsM56tPnb1T6nrs7aYwogQ4n3oP
BNnwixLiqTHnuG82Qu24ENolgTvLymIBfVieTlHBSmxVzhb3PJNalDSnqTpB
OH8bbOZn5Vn2WhIVaJsNx2/mNjZGgUrhivAnkOJ5Q9ox8bYTvzmWr+jtVOLO
RhUoxSYBk/4zVlsKMJyd9YY/2mBLXKCOzGxobuV59T+kz6iLxY0DQfI10iBq
AiB9TYtE2B1waeaQqV6WntSPZq+jectnrAC0+xI2Bpp9VlIU+dAGt8MqOA98
b0oe9Y4ivS0X0ZIXC8HU2rB3fF6fTDrYPwklTrWVMDCz2PWwp7QYZucbmSZp
Nde15f19RrMSefwyF08hm2p8o3R58gxCNmxbEyHhbqFp1pKIWlllSYqSbcgZ
lFicUwktDmEw58LLTaxiYTw/8MCV3wS/jBCyhz5bTkUn81N9wE40ShybTcRw
aijXHIX6Hjs5JWxxm9SlFEiU8vKH4hTFshKSeEPC1s2aXlKkkjQpLZvnEdLf
8HqvZOy5OTa4iqNTfGJJaW6jHe858QQgWRBKxlGHwGQojbFVJoYzKXF8BRt8
RHJR7F9fbCD1uB+VCPcqY19h4Dz9mFMgz5ECjWui9ajTZ6MdfE6GhigXa7Id
UZUN2W1EykTJS16m4ix6lgHHnC10BCpsuKPDK+hqopVe7uUEWwYpJjm8C3Yq
yjCU5eF87HUz8lJupD5EFtU3+D5zFCL4ONM53936KQhLB4rMPX4QIP+E9mgW
09L2U+6XoPzCn25TuYeEt691v4+T6CqKcQcoTMYI0MsDHvs/A6/7O67y6gig
zurxQD6ksRvt1BZ4LPy4C+NcXk8YJdKltS/J4eqd9gU0+CMRcRtmrg6eBymU
0FYfuExaLi8xQQNi15WnF1Y+2dJ9/8Gg9ZjwPf+Y5lqmJ3+0NMFpeneDaTfd
1hqAFatt+HvBPxM5QyaQSL1Mau/4c2q+8MMzVXjaMT8uliudgpkV4O1b5tFv
rLLRVPzkazWYfIHvKF2K4bEMvv4/RWsEEA8iZOcG0H/ZzGB6tE6ZLW8p+fkY
SGMH2A1wSxyrjuNWwZOFyCx3N3f5xbhhNOfqKsvhK/OIguWfmitz3Z3em0in
dsKj8XGhA2ikmROooBt/T8Qtm/A3mS8RdBPySy56cLrLFKMaksa/3e0Yd+fY
0UgoOqLqA3whojyxl+x90r6BdWgZdAL1+de2Lld4jK0q1/uL9qqId2Em4vrk
XTe/XT9Wc3pdN6eNnezQK5J0tUhDwSzRbaPdE5lNhVFbQ75/WWQdNW9650O9
O4b0zv8OqoBrEQmwoZXb5SgocfOlRAFxgATuwHJ2r6E3gKsZiFNC5aaYBB6D
qELEdweBe56dof3UgODbkKDXSxZZYm3mlwYU54K3QxH/sQN9bcmS4UHYOyLZ
3EMXlfvU9H/swqg5ONhMszsKSVnydd9EjLgrJkjtjMW6cFgYPNrtApTH+mpd
2mLM0D4Xt6HbjgSAYOO75ui+dBvVjiCG/XDktZ0lZz6xXICgssoBq7WFNCK0
1xjTZFA3PKNkoCeJ/qmubjF/cCp7dif1dGKi8krLuccee97FMEcr3PR6PBkt
CU81iwTN2QnC+2CWwjB8OxwDfnTg+jpNOTnSJSlslpEYOTzaJnw/xLLGpv2+
dk+ZNlM0HZIIksi1kzyRx8ix/VDMt4y7XXdeIs07dFtGZ6zYDNHXcFbczL1I
KIqqji/QW6vRwqeOjO8jpE/tHRHSs2mv0Z6MbJSyWTD8RlipZbrh6ETGrNUp
30Bw/mGY5G844i+RpkfWiAqt/l14reFmkawn4IVGr5n9vhG6Z5jxki+hKDuZ
uWVdPoa+oyP0+W36CCV1a6mV0AWooYN2C+wysD4PLNEg6F0FdbjSep74sJvw
CV9Z7etF6yIXwZvm9GI2W0YupAWv2ihRWgV6xWokV0ERzO/JZFurtkc3wcM6
VPkMpeie+vATByf7pzt6qn/11RNOUSnp9ejSP8/uyp83lvwzBMVaezF1Uflr
tQpqlPt9zaSdCHuZ9URMQIFBPtSjxsUi4dmCwYrDZ9MSerjo4YyXD8BOb93S
1ytJyuBK0iMhTS8TrQqzt89E8GZcTVBRAGPvMrCSw/5L2FFMV8AFFeNIVlmF
r5EX9oJgDRLadXo9VqfkXv5yR0lUdUnv0T+hlWU8pcRhbx9wZIpk0vUj4zZL
iYohCsp+EaWq67YRW3NTg/u5ZpXZUvhaymNv8z21Q/ncXWaVl6+1+MV81ehQ
Wi/agPwhGQrgyvoAoAECZ0z7GWlscR6bFCsuf3ZVnhp9a28K9R7JNl6oJb2U
9NtZPpzsS3PPRA+7fkGGOr310zO7RApSC75RT3kcuZOn0zzJ9dxT07PhyFxd
0xoaI1x07mf3WCzUT5Y5pFBL7JPTmv9s+xsoEV6S7sbyUE8YtH2zsnTycCqj
/qiLMNF34HH0P1us4IhnrQfr7yxlxV5GQTSuKsLwO8pEsSQZg5U8rLMaRe6K
3hfefhOqvcPRHgFGMhZEhECxthdeQOO5XQ5OYbaX6FISztafXg9Fd0riJeuZ
Fb6JASbtujYYFB5zKemYBvmrNo5PXZU2OMkA3yz4/se5LwZBJUjIpr4k/HXr
XT74LNBBMR7lpZF/QJmft0B2B4/sB7UklzH32n4ktCBt0JW6HET0kcebhiW2
w5cdE4vKxkW7wbhSnXIdfiveg4BIyKJH9dYZXf8qlfXw1t9nxztVVE2Uzpcu
ckj1ow3foWTLddhrD4JZdwwQEM/YHUVffyeXHXGxz36pOIggMdasnyxajbIO
1IKD+Vnc7R0gZAjChZp4xZ3bGPv+ZTvbVH7iJSRxDnhcqaghtezyPr7XJU9j
IeUDfKF4bGTz1pNwkjUfV4BY0CIEIYsi5EKI6ylZq5Df8bt2pUZWPXdRdM0j
EymMbSHA7AZhf6Y7VwGrPs/jmbpO1x99fQ7MRBkfr5ON7CG3sSBXGXi4+80O
NniCYLt8WjejighRGL7LiKr0yhFL+H0nTZodUfx3KSYUjrsdCKKQJCv4mDA4
scE2+133te2t4OVJvtitJ2l/qrN1iDBW0zsNp9oQsmfj6kAqEvgbMaenTTcz
CVEVjMtTHaKyAgBHFpoMKukbzWKLiBAbQKYiZeNGaOHReZ2Qg8Amu6BF6JzM
ENZi+TCQeKZpXxEdBFdu0Y4kqcLHb6EFpGQzXB5m4pxp7DsM2q7iujlzBwRe
CZPwYIonSJONJkhC/X+CdXNpw4fylfVFpjzWAn64IG06hli6qseMKRAqB/jJ
laGKJahKy07ZCP0sLxC4OkccJL9d7udevn+HAbkIgYwu/VGaFj3AnLnjF4Te
ZH0BE0mrq+nYwEHGKqVf1wU74H1KFDv54qzQkPwPz4OU4XCLGQGHdkm2PKl4
ZtwDXWxXZLYhdJLUv+DR0V1cVOaapTS6AzTcol70QOt0zPammNcajX5eepdO
9JZLbwCax5X/VOx0qmg7nwLUOWd6AFlwwoy3Q+Y/FAy7wf0OOFLrc60MPvAe
bYQkDU4GijeVnwaC2iMN7jLPC7dXDWGu7r1rB0vtld9q+cSEqRGo/c9VMGRn
9FvJqKWEcJZNM9aUcHxystnnBbdW1HWedkGa15risE/lgPE9rAFmiNmlUVUv
dIuQN7b7Dly7L+h6fX+F1QQhnpJwC/ZgpEgr9S4b4Si7zffhpMkEIYLFdSLk
Pv2ojomNLrb1PEfN2kODpv/a5ZOo9NL90e0p2tdCmMU+Ji/GfYnMgpB/Z4pb
DIe9P8FVfOZ/NqfDGMvrWuT4BN1byPqkfPqaXBVOkWmpGR8KGHyfqUYrXwgH
zfJRHpK5IdBnT4juUFVjedEuYkjMxvyUFCC/Lzq+jCYZ33r6VJy6d0EBFy1G
ADGNCus4feBXG81bWfwMr3NK4v2efMWjLE427WQc2zxTQy/QzKI6qLVZgOXm
znfoV8qiP8M+D4L2Z7F9n/hXjsY+UiE/f9696g03lfcL4LVvpIp1AR2VMI/b
QQNR1J+e+BL9gZQCWEIQLFCv8Ogx+ajnn2Ypbq4RlNDFJzl5xypAmWpJnlwN
FXPhV3BB2GV5VAUuz1JdZMFzsx0FaWT6nLBH7PGGSzhTVpUoN1XV3sa2XuSy
smz/05ER6zknDjDcsNvEaEVAe05XNwARqMd732MUk06J1oiytRTtWYdKKMKU
m6nq5B7EC2AF8W3h7Nme4ajutEC/jX+JL9+7XmHcXdIUxhVDS31fENQd5JHO
JdoUxmv4S77zhVFfpy29uLAFm9pLyelmymEV2D5523Wxvd88yBtQmWqfRo+g
UGcslAy05mlGRi3ixVnq7zPNzlxtiIZ5i3+8mYs5CsvvEPGtCM35a8IrIrg7
Uj6Z7m3g8xf6vV98HA6c8gHXQ15XF0ALKE5WAuuKoQw5dBSOL2yZjyW47thX
DEfe6roBdIqcx7IYb6N9qkmSrNRGWQ29XhKDMO2XfwuiT1GL0PBVkGn1sgK0
qSGDulKsrbO4eiBEDdeX1LNMoOMPzAG3/0UsQBXQvkIMBaNpldVfqaWq1piy
+i2IW/M+WtIrsarFNvHfYpI+APfXzCkGYaXjZPQ/75RmUwGZRxX9lvxE740b
X3lQYPBjUM/UrIvfz/e6+Cga8qXaSGvJbc1hSbfiSkAk2VAPb+0WE+d0LtXP
hfJDn0OimqUTDqVJsQRkroUn1uzSJl7YZm0rkVZp6HWdtL88DIICDIBb4Dy6
XquKYNtR58bzYDYBp7bHeIIagWa/Pe5R2f0i7Rwvqm34kIceiDA5yczp2fOl
i+ZHe0UE1Qm2i3+nGjlXeaZDQVGM1yfFSgcmJKv76YJjsTHGAfUa82uNt1vc
2Bf29TFdSvcricWhsLR59kSI9E95MQ7P2z/k/H2iFw9qwp+X3fqcxgrt2hAv
DUYUm+vD+t6b/D2Db+CFzBZtwgtMiQqOZTTVgVA6NVIuzo/8Mg5KLbYZRCPS
TeMWQufUoWzx4PGYndJ/nBQhTIRM1YQPFeEoS0jJA9AHb9+SJt5rUyLAtG4W
dTv+R61C+pASnB1Yn0H8FiRVgb171N+PV+AJudZr+OzqBH8tjCw1e6YhIgli
kIRe6fobg13sGz9Y/2Fa3VCbybzkub4GoJNwdBZBiP6HaP0TnH//k8Rt8uLt
d4m5H37gOa4aYu6YOPqT0EXL9ApXhEeLVjfeQHiDtQ9as7TISrNrR69jHF+D
ysTVkrf46X3KwCQMU0YCrQvlkn8SPlSOPcHSrET+lDEAxHmC2Yi7FwWEtwZL
brwLB53+o020fp04VFjGT6nrjwikmWG7O7+E9ZN8IyOnLa3YxKo2A/iWe/rZ
cuZKjPCYuj1/gLmAXFZDXk6k2AF3OWbjfAgdvnBj/jeXcbYqx84Xs7pJZYAQ
ndJnZ8Ch8RGQZ/9U/15I7sdDH5wE95VPBbxdj3X/mbv313dGpDQrCntONe1h
nfFGHK0TEaCf0ERFcOuLefblP73J7tdHWNs4iJds2uHo1jLzwytdm8UfWWf5
ebkSWnHj4HNToQJ56qnFd3SNNM1rO4v7vxbGstKUrZsW7CcAWB9jFjUMJfcD
Ogg7JJsSLb7BDOOsY4V+lshQHpLNIl7NF3JyqCdP3HDm8lA4rFZZm/ZXcQBN
ehzpwd8COJHrkgbY0O9GDLAqtmcPRLPOlN1E/oapunwzbu4yExJLKd8/mHfr
YxVMcqnIBmbGa0cqxAe1JcmmggWnfBUpGiuApO9Nda8vSSAwrND9a3jZvlih
vDARBaRj4bUUKc9pu44vaPJVMVVR3xHJbZeYjJwdRyUJiGuv4AZiR7T0JsBM
hxjzXw8v2dzRe/AAMsqMEdFu5NnyvxY9PVJ0CnYFmyolu9hR7SUnSVZsnoFk
+slpc4x9KLVC/YuBeKEtKR7qWr6eAg6kwXpKZBul3A4DOwRhfHG8o09sPdo7
LOaoE59n6uvSTMc9oe76wyw6pia25zH/VX3EtWC/VUvGZs8SKi0+ymBED0g6
k7tfyriqtS3/AiDbTHqDRcitBS4m9TBLFZpsvl76SLXT6CLUMPXz5MVgiWge
aVwYhQbj2okam8+SvbugL/3zvRsCk3/YXZ08EtKg7qOKsj24jI1LicTgHlfx
DNHnATbpMUgzcpNc69v48UYxMNPWYQp1KAwRn2fpEsWuoWOKnyMn//GtUZ8g
oXwJqMoy2Pjj2b+7y5L1JO6Z38lZ7+s6b3/eJi9AyR+tw4hb3hKXOOozjNPl
Zu1k/Zf7j/ap+bC84aXcmZgi+oCHZ9TfE8q5j55OeHNJjt5XRfJaSQAi6vRz
GmLLyUtUgpqFmCH1fLu7U+/ybikiNRkTm+jPigS9cDcwIFXMnGucBmYpck1Z
ng9n1xaDkNrR0Q1h47tDBDDsinzNhK08rJSZ05WUYkPWpNtQjj/oBKBcSFy+
BNjrSOZj0UFfjUfKXxv1u5wf24802zW5WM6JwJFzv8g3uFl7yfqNFU6IKTRb
/sdriSSq24D9lCRIOGY511xb4GDh3nb3RsWQmae3tlfviTk2cXoGglHvnoiL
ljEgGOWfiE/7/SrPzgNsB6i+bIBiqrfb24IuKLnCCNr5aWveac5jClbi1HAL
Lga+NCCPiANCzIkC3vui/U3wMn4FaSMQ8aJpz5rherG4TtROddWk9Z3TIy1X
rwEjYUhMNIrKHZ0QXm/10QSbuiiGBXkvCRVeDq6XOPKWbweTSAgoPTf86EO8
Y9M/d7LmkFsM9MwycCwtX9iNBgOa5JAJaPY73XvxQ41SxU81MXieRxC3wQM9
IaaZt35nFlck8HgaXkb5SNIvuKR78QMkZuZnv+QUCImJyywavZOey1XGvwyq
cpa+rlasMvdII8YzNRU/TTh6zdIkYE8ElYMgcRZYIC8c0gUn0wb0kI2WAeeL
9prersjztLteNjHIP8kXdZ8ZSOkIqbFW7t+VZnGzqwtZgUW46NXh8qwdFrB3
M6/lIOvErIbvWfR1JxvCDPu6BcjpE1PNFS+Rbyy+qtb8gScqU5RfrS8vvrms
Ru1aUqkgAqQN6kn7MehLbLquFbw8EkZ3+Uz6Gx3838LdiGYnSVj5d8Xx6773
Nhm2XNWLLVvei1Lxs/2kr6RPQrEZFX7fbFqzASoOv911zZ5ZZS0G0q8Gaoc/
CkwbCIO6XvmtdPyjmgRF5yVJTCbZLT2NA7fn8yIyhk6dsbt7vGN2SENYeMN1
wbbddkW/qnv1MZ1zZLk9Dv4uj7xgIkBraoKPqZtrnZY+/k+sfEXWIJnjyea1
LetIg9DM2FhASa1Uk6Ljq2Op/8zz+Ggbl9OQimntqTM1GYS2coI4DAu7tJIJ
lSs4ylx/yVXrHflNOUMYU5i8cITu8EsDfGKuMGKcVcgE8sC5Jheh7e/+sv7X
B/Fb/4+j/QpEzB4o/nP/xS4YjLTnGLQ5PrIG6plwU8Dwdf6z8ScdfBhfYCoI
4q2kVIzn2zPLb02T0M30O+7TPPmbMlyJMreNfBkLqL9fTQwhZWkDVE221/mC
MBEzFlecoJ2Q0wG67n0ig8THXs+niq/CzPS2DQC3chA8qA3+IByA1lBJcSEi
d1nhlqmXklK2JBQiYSY+ozVIQ+pRDv5rKdPtLtccFP+c0QvYamnqMM7M9zWd
RNv+wlWurmABCxLWY/xJ4yqTyTV2DR71e38JUILsS+aHkIBI9czhdhjfUTPC
cjEEWohiejRP4VPo10UItLlCJ+vZXX00JfhmfHJ0bmwtODhnzfP27lmb+qxv
sOqQYcAvpAUfod/TxZgAjUVA/u5Ke5cqYM36FBZbIi3Fg1OSqlrf1QzD4OYV
mLMXF8+VRm2abHXU8u4ROGQSnJ+EYBjRvSTQmfW/4uD5aVmnZHcrll3gRpuO
19FcnLqcP35NuiyAWfmmS61o4PoG5hk3+lvy4Zwk2IeR942+BA+1uX7ycI0e
i4WIint0bRGX7pu91z+tdKNMAIV8wP19waAgS517ZWOq6BXtv7x/fK+Z2zd+
Au64n3TgnbYekDYo8OiwEXYEiE7D7h6CD9am3UxdJ8QEhtQ55NRFVMOwlGAQ
5jU+wbgO1YUnAGjauOAVKzBON/VJNUcT9ptg1WXWppdMsO3mtT5Viko+UE0o
nntkoSy2QvdujLMzeWL8zNzHYP093imSrZC3c4nAGQLUhRJeYwjIiSLCnXty
bL1DO+4vUZ1xps2lA2Eb3JgaClDnLWOk/75leBGkxcKi/Oll0gwL1VTvBaVe
Fgc4l7ifY9XyTrPGBtrVYlGBFrWHbZSnAhESdvvQqOWTi0PlvksmVHwoaBDU
wExjqyuLP/jayh3/wmLO9OgCOeZa/sJ0GeDlf5yv09jel66UOlUu0/BjakxZ
h/opnvGWxNk/3aZsID/chS52yjlAGzNVRmuN1C5KROZt2hAX/6ZWAwTKFpHh
wS4b8sl3/048zmGn7aH/+bOHlVGmgAXVpPlDgurb1NPYtGoMJNwgzITR4cN6
O/8LXxYhx8lLfjXenX/gPlyjTZAW3U+/Bjb4KHINJorSzilYMRRa6TYH/BvS
9CDp5XVBGm09g4/bK3ksf7/cianwPHoBS0aJG8x4X6yNXE9aEgZQQX+ez3xy
GOqXBlCRQZp4I93vB6CPBw6UVXPIx10S6j5/PoPk1Rh9bdMeKKDJ2qX5QJLf
ZmVW1gQB03PhV0YuTe5xIY9wvFo9Z5H1OHnEYHROrjMof0Tab3FJMsSIm9Nw
o3dF9KWfet7vpcgscdTQNeDEtc8yfzU0UkCLzIGGDrqb6ZpzOJxL9DWtf4Ji
dtbh1iaKQdlSFgZnDxTKL/3fXaTv3xYWB6K/0hTcGG9OPK7+okXqbGLR7gF6
xcKisLajl/nnJCVnakynfJC/2YUQ3e6gdD6tIfXm3M9e1DEkoZnPzTYr5xK2
0Qmt4eNi4+ij3LlfvUgmxR1aRyGlxlPeXCSo4Lgw/oh4ov7/7dRiWvJW9LTa
rmghIASnfEghVqUliu9gzp6KmJp1sSqKr4EEyzJLfIYOgIgmHJoFGeqQaiWg
HZfPJw7AGePNpPmOX41YgcV7FkD9kuHxQFY5E12ZILf3UpT/iD3/ZuDSmzxQ
kPbfN0avAilEmPR55gP/lAMHsR6VtAuO33L3XSY1p5q20dRPnz4eioWuS0QR
JnISrLyrn4ibErWMILtjiiG7vcyN/ZDY61K/cCjs7Pou9sA2HgabSPk8p5PH
CgBAL7LiqBWLdhmz5ce5oVE0KIEiMJdsJ/74ZpA9K2XjeH+rYwsxuucIsobj
aJh62hamNTVMh2OqaO+iQw9yAdnrCfS53LqvqUr2/WObJYUWJAIbqSba1Z4l
W4DgAnyCSBb5duI11R9qia+W2kLSk4l6/R0Q9D723WcZ/UL+tp//FvMsyZts
tpeS1yOJyUtaMPzB3iA1a6DCzCf2mi/wsOtk0Ohk6Wx3PIVi3h7nNiegiN59
6PKeW51VfnFaU24Yx67pMIuOmHJxqxBkdnTGb98h7LSPeJUaBDJi1JF51rDz
j0DmOH09/1pFoNYt9KGU8r8nQv4OYv8p/WcyRhefevHKxpXCqSDS8hDIPZPT
2MAwKTNnY84iZreHB52u6eOqRsqZcdhlNjOj/gk7GF3AJ7VD4cn8yCmviSqe
gK/WEJQHIAFupkh3342GAjZ0wVRZBdFDW/TybS88cWOUJT3BSk+4q3JEh4Rj
tysErWytvWAfxS30NkwGaIe9wtXo4tnXxMW0LQOD+OUaFoxJfth5kgScx8NU
K9/nhLzQDhaMhbvdcMCHC+iBJNF1xLoB19yTmGXmanbOScX0K5sQHeidfqUf
WLa8JnP7M0ZvaYwEWzEJM0ntPC0Hd3vc7sffinNou0aLgCp4dnqMYH6C8jQI
REbVtkbl3VgaYUvZDpIWBXuDRzkiAtArP4x0Nt8tfOWZ30UYPXQQ41LDFhpE
xgWctKD435JsThxsxfkIZFXchwfoZ5c7P1jOYz2tLfgvUK10vyaIaW1E2dwG
Ju02/0F+2njA4Nz/PAVj+rIcADwPI3CWEeusp7sb3fWJ9M3qMiVHAJuWbh71
2eUJD8sf/vztQmM2q2uNMdZ76dj5pI3lwD4pFI3+7ckqt32b31750i0eqkIo
RVNi2MCTQM/C8ircdUb8tjzk6+sdvJOsHlJbIl7WLjPgcnjGEwrbHaHW5k6A
nS0N9b7HPILbxQUYY6e6lVHmS+vTg1cNJ5OP4fq3jplAwi9yof/VDT6q48MC
wIpAU5eCPvmiR7ox+jqpzQT+kr0tYoAiCu/dalb3alPIOCFCkIZyeuJ4iG89
eUKZOftBPL6+ZntWxYcqktY0id9070CVeGlYFyhZCUqVrg9ZAE91uYSszucL
RHr/qbLOqK5dwyz0qpv4IxlaZegnBMpvDLQwgFFshOgSNp8GxEZ+pSczpmun
jfq+mZaqKfuqPX+sLd/D4+HSxA2ua485ux5ZH6B392vB4RNo6II5itRf2hPC
75IoWcN4EOL2QggeLCMv4Pc4G1s4XDehqO49S7h6BgDCEb8sPdT6E2NlxppX
PXnODkGM2ddxqWGT+yG15iJS1/jwVtcgqjtVi7ifaoQJEdTk7bwL9CB5Odsk
z5Urlm4Wqb4wMU9c2M3gwgD6z9SH+TLyRigQsCZ24eQD9skwRRgSo92QwhtT
k43IwDk1lLUG2B81JCa2MCdDtewapm+vIfCsgw8rMIv4oVpKV3nS1N5olzyW
jP7+2EjLPl+TpqAkMn3WY8nBXyVZqkzYrKOSO2uerSRMkY9M/2kf0OpqFPyd
pVDgXEkD9pxPYnE7DmEGfKN1jRE7udMmrh+A2z9CgQ1PVwXr6YILGV6vDTdF
PqyGjxRYkP4jcCFz1/0t44FT6I3Hu/wa13oxUoCeBJdxxDnEv2gbnNR+REz3
NQ4Upo2T9h4Bm/A8tioQuJfxp7D0MvVNixlE2G/P0o1JWPSnO3/MGw2Px3Hu
4TamqIC4wF+bOZUfPcsgaOxpzG3wcn9/Pg57H7eEwN5feyE68rYObcATztMq
2fNKN5LaPMXVJKg5FXbMRyUsbn5+puohdakZkxOnBOq2rv7gnEnIBZYVKRSS
VHIR9M8X3Gju21glwRTgH4kX9IiAj1iXh8K0V+POUjFgfFb+iYqCLVVN0yeP
g36T/yjF6fBzNSIsEn4BHp/bR34UYhTN+OXN0FJOxcfEInKWfgH0v6DYCKoy
KGBPWXmpMxRlGwq/jpJr4WusZK+DLjGxrLJCVDHvJVMkhsOE5fORUt+bTLkb
rfHejJE/PkE41zMqeJf37BMnBEmmWmp5PYZ+ltLwKO1PIon4pxZVtEVoMSPv
xJEbQXrgFs2Qj0cHRGeNG0+FdUma1EbFsTqrp0aXr9FYXWFocwDcvYfbnLZn
4JUac/VbBR3HYF9MUfI/eAQx79czc36KCKEWJ2k9d16R3sGjAPnq4/rQTOLg
aefnCzXSv+cQ7C/RsqMUF5WCz8o9NPDgLMJDADkO1lWJk4aO5iuzZ0n7aVdo
XcNIoEluwQKuIU6+dUNe6SU5LYI3ntYmzV10cUpY2398opHYrLCh8RmGQED2
wgT9NBM6lPR16q9fWP0eIf4yWwNRE7uJ36iEpsWfeUVWvm2Ouirho6zrAPIF
tYJtJIPXJPeZkeaBZ+stpjnL6w7tWV15B9f8VxCx6FaDJ8NiEpAhKAdIq0n3
giOLj361/LuNkgADiUiksRokrbSiwlc7C1o56XdafKBOvE0kWhaI4PPhisWm
1Yk/m/QNScitLAwTJEOqmQMa88sPDDzVscI1B6EXwqbyzM4kWobD2OOpokZZ
ty5aT0SLPo1tj8kvo67Z9C22NRxQ2p7fjnXfrWzn3HuNuedLtZH5rqzLUPtp
3dPrPg1OIsZ5S319jG7vyDREruq5r+zexK5GJhE+V0G9tGFkaslSg2pTfyf5
ajjG/XgkDoiv0vbxbaazmbipNEY4UO03lqV97IoYevfE5IP9w4s2ZCQOuRWm
RRM7HZWHbRBmybCGANYd2CNYZEYrfpTgDw90TQtFE/4X1ahJUVvVOeqXjPut
6+VGPJ90E4eQhJ3aD4EOE4EGA8c0RqEow2fD0Ko8UbrozPeBMYLSecr6a8z1
A+Afw/8zvPc4TKLmSAKnZ8yvWpkzWCTOyg0moeDnUNvPm6fwbP2QgkYXJktf
5T051uR5iXkJQIXRn8zYdyAw0o5H0fqa2Wn8TJPuNP9OGF3yJghDF1B5NVr4
+FHNxwSOZaIeozhOc8S3CoskXlKbonZ/eeTccGMr/2+1qVz0HP3PaLQDBdh3
p37ZbXn1MxPw/eg0iTdwlW519fPEj9XPAnpvplsQw1uT/S8khQaLaObXoN9Q
f6q7l1zmhPBVrhsiHO/R/v4A1H57ehhPYMfxN2NOvVuzo52hQnSNwKm7OEI1
l+zyyNiTAsUNZPTyGWONedMnK2sg1f5kQjH8yKFf4MOG+nibHtpVv36zRQlN
yrzcUBeyNZeYmZZOjGvec7c7NH6chG5Iw4LCvCUEEtxDk9sCNo//moB60o/e
9jSYopcqkQqD1SDc/vQOshiYbU3+nlAOqG+9MmP1jzDa1KmjB9irW4KHdgBK
s7l/wqEq6A6Oah8hH+tWdrn5/czb1w8OL+Etg7tzyGL81HpyYjuMy1XbVI+/
JwM5TKyPowtKy9HgYlsQjOdVN8vw8pIwWcPYY9uvHFfPclYDIY7GUaT2NfZf
uqxZ7QpHzApiVEeU51zbVG3/OZUh4uDBF5vFf/XNi6lSTyqzck7VFLyK7rek
OUWgBwx/pr0DW+SQbaAXiffaQ4UBhz4/Xq8DYAQWHDPqt6icqfY4aV/SALVe
6MPNpUVYWz7C6gxqOIdhZHUcHxhnO+ourQbGiSvtQmgiJeKGqQBr/EcM66z+
sCfxt9nLkR8v5SEkvnTJGSQTpuy/Fa+UfXvzwONBEA3UTn32I/Fwmc1k+ES6
YaHPu7+uz4+QLqb/MfZ6PEFAKos4HnbuV6WqslWH2hnWhL+5Pg38neGJKtyZ
npyozVu7hR0Jl0RxNdbR9aPux17D5UDnWXxXTAyGhLg+pHjQ8cWonqFcBUTc
6uEIj+1l9XpyO8IwTDRJ+D4lqC8bfcvQHKJnCANqdZA5gJgxNzBOHBIokttG
5FSvmu0PAgR9SnZ714RdiP+l8yZRirwiV7upUAxRejiDUKO2dgVT7ttUSANm
AIXApVzt/tavnYBbiBCqMP5jBRI6SS82/NEfYVH/GnuZkUlMJ8PeTmjOnR12
z2eW67YkxxkvWFybeVU7JXyMefU4QYWeS7JiGJ4DOobWKsdS6rsYWHaqW6TZ
m1qoq3BtJ7ur6fWvKW9K1MltmCvchx5op6p6jCy9r6AYW6wbeisvvi9A7a2y
L/1BGW4tCUM2K/S3FyJjupMi9z86lvRU1QRBffl1GyQZdtZnpQabiUooslmt
oZBqcEcTngmoysV/kPNwFvOFudbwGN5mGCD0WKj8a43ET1WNURf5wwH5Kwog
GenIeAGQ+Aji0e07bykPbe79aTsHXcRE31habwucFkE2yURb+e2fQ1syPmPC
Zb+w7OD3wuBSH9MyJfX2luQsXwTIcd51QVejJt4lfdtEXfuTtFo8kyZJmqPu
3CnDq/im7qVrMes1qc8YNTOmbyJEIdSkRq+17Adw4s1wNYnML/JwYMiZzUD+
vTDsQ/i09WkpA+mCvLyAswgc1TSYuerEYvuRuWuiG0uP81ExZzsJc11HnXPh
H440F3K1/IHrF1/ZI+2jUyyxQiw02bZna3ATIwGSJzqSybpu9SmYaEl3mUwI
hg4Hz3iSrKNICYG6zM71/+oj6j5jSEDOVJifxxiu4C7LPy58TF4HYFzJqQRD
zKICDWJordjT7azFDmypnUNpeG2AJdQV5tbBNeu6/MRRHXyGQy/J0siUUK3x
OssxoJIrOqprgxpsHKEcHSnslotmbffRPLoRgoxFNoGMrrTb0qWZS4xx3GmK
anRdGt2PMC5ZlhaDPqzvkRTqa76wb0cZHfDJRuAfHMm4x6/vd4VsP+BlpILU
oBwgKaWCEbdMcnwKfAlCClnUt6B9VKgwPnZ4ODzxloESMIFDAKKnBpFSnHPf
P7IIm3VOGVeI+MCFqIc8n3cMUpSHWT1H4EA/3j9Cb8d7S4IkR1EjZLafOGS4
hOq8Tp4O/D0dIFa2MSWBM+cK2NyVgmlu18EOHRNVdz9BH7N/Y2f+NTrXlfzL
mc6bGBEQOzTFVv1qgs10kVYiIbbIFkr+xPDcHKJ/On+W6j1anJzJ2gODlzd5
A1DJSZGYoSuIPusG1WlR52H0gnDvDZ8cj8IUOpmjK8AO4IpIhOfcX8nYivXI
5/9xa8Hs5fIf6VGJh8yIkmT+KkDV3sBy0PNHV8gcCny5ROAZ/o8/ttDK+Wbi
GQld4DUWGLKbZkchhx4tQJE1fMotBy4Og8jqBxs77HOUw4KcDO/9i1v3a7SL
JWMv286iMRRj7QZP5EIbGn4fxTPXURkjgOPO+orirlI/Kqt4HW+wArW34T+Z
M9K5jx4jTOBt2gz4+PudjH7h5m+nM7DG8moJm6myMrAkK+njwfpmifmbLhs0
b42GJGIIDXCbBVLiPnMOi099DD/jUnNcGubL42Hlvv+8vT4msrnFxVO38fqY
r1o02IpCpNuOBnGn0yOSS1B4YFXGIh8XHPYzSdPdSuzh+EAx0CIGK9CHsM+N
aEeH1WMM2azfhqCk/QmkuO/Z3peDZ+S+aAoUqvYyBKR4aRFU3QZJa2YiPDO5
pB1yQOT9adqqvX6GNCE+7THTAu7CMULjaVDC/LnjrEwYZk15OmXPL/bk+rfl
iqX93d9wda3jEGcxJldE4BR/GNC3fhiyH6AYqA8B2EGBfIbAEvahf1Tj8IAY
fPzJHGnsyx9Ng7IkaHWLSP09rgsK/6qmEEg/GM9a5jlxHObmK9mcpZ8NEUEL
m2dd27xbgOAryJsK5xjdKb3tsmSIAqSqoEDQEp/gG7SRCQCJHaMcaCoT09VE
1gh4ieeRdoSyIQeKk/g6TLhl6+pyvWy1BNe9plsZz52oq1Ad32G9onk0L3nD
cvHUkV+1wcuqIZc9AgKhMk271phEkuaAQb+2TkX5Tq+fMPDObbSKpfAB32O5
3MzVaIBIqXmMEfYO+8Wnr8+efjGtSpqvFJHlGWcG9M0qAtvgnm+Pb4hpnUt+
x31SZ96ookRebBosPQUaotj+FIBacwZv6j/i+QbufDxntmd4nJTG4GezVYs1
NV19fgWpjpAeCOdRhYVLkqAOCIQrq4/PmpQZFBkLy7TzL8RKzaT9Md3dq5Ki
rL+P+bDQVpZQeXr7BWSDlcvmjvjL+yo20u66OZnxlmpnt9OnwXaSsO3hEbX5
+kFb4jbLKLtAZgN51zN8E3HnacKb5x2jbcYVQIrpIgNWXoj3OKqNf5UGHaK8
n1CMOCuLbRTnviaY0QdNfrtOVZpvi0LTa8YkrHqznEDZjVubDCYTIkT9h9D3
KsMBiukZTbyRt+HmJam2xX5lJJKxJ48miAywk1tPdaMhZHMPj+kTaDIFajxU
AM8UWp7fT/GpWA5SaKGqsxNT7OvAztZ4kWqL9LwCA+7RRXgApggGK81nVQAG
E7bZkdTgWS7pHE0BZRfqDRTHzfzzTml8osZMnEN51YGsbE3YLsFOyDELSv60
OACOqs1Ct7qSctG6z5IApLhON8wtKfcvmpfYD82K/nlAO7Xt07kkK51fTVQY
2FV6ELgFDZyxk9ZK6sksQc/78Yj/pPwuDydj6Wr4pwynL0bhn5rbKeUw0kld
np+6ZTPFUe/hecNI/iKtIZNyDkatMg42m5B7E+8R2Pwa4m4R1zf8J3M7O2XK
pX9wLAw0kzjAfTuZhb1uBPSzrX0Ihfi7L1C85jzoycDtfFYhmsRwEhWERmfV
+Y7lSHqP9G5s1kuWRcsIG6VqDZBNI5FZ1E33EDrC2pumN/CwpVFzGxBj9lLv
tcvqksbm24Els1GQfzbJL3KCr+NsL9wrI7tPe66aoj+iovmaVce7t7hNx72w
wueLr/qAhKx9xrtpi1Y1UGuvujQIPVIflq1FbmDT792e4ma4SOAzp37zOLQj
qX57K9sAHA+7a+CwZa1EjmXl0oKuDoXCtry7sQwLJ7vBJWhhNKIjHLz2n6to
qeKNgMnAsTd3zM4AIR1pbnAfrE5QReL9jX63fE1XZZQr4IINquBu1eUp3GGA
pGPX2NjkHYiB3ewL3alt9p4uqJ7qsJfOMnC5y0xsMZ689eGbK4IN2izeLQNM
0JCvWI7w+KuvPXj3DwhUAPMy/cvLlsQ/w3Juzfzune4OQDCMdraoxjsP5aJG
ITSMyfy7m5eR4Vt+bIeuE5+sNvkpA5OzyR+t6yohv9lQG4i5JlMK3JP/WwWq
L6la/T2qiTyadpKSSlLOZRI7dqo2EVIVn89QyoI6tjRHCK3rXEoXEZZbaygN
gc3H88LBEScACs4QpT3LRA7agP+Blqz5iyQSpeoYiZ7VvJSI77f59Ero9dtv
sW1JAgw54sSSEj/3Wjybqufm2cuBjPjVhOrZgSAQKolqwJlV4BMl+PNNLTLs
NVtpFXZXkj1Xx+vqasOHeLMiItrt3NTwTunJ85yS929dyrvX9EA3eqi8GxxZ
DYw57RMpuR6ZUmn2x+b6kUAUWmEIR+kEYSjomzt2e2d8myb9s6MwLbgYkr62
zwdJJ40rAVurozBdd1FvbvnlfRd/ksjO1xhyRwisVvi5I/A8MLVC4DUnUHKa
MY81IdWIhKIY8CIuoW8YgfbJcOg/lDRY2WayJvKCBXDXbygy3s6iTb0BGJx6
VactsA8xA4EO8ZDAVaJGcxcD6XUYuWr8nVvyVxk0ttymHerfjuysSf5RaVm9
bS5ROtR30LkwBETOkL6JTn0YJ36wlFqLpsL/KAuVABC+jadZx+ugvwaD6oYc
+JCW7HLYiTqIjUCbvlIWmfFjmgBzQulWHQSE+0tQSolFwnpLXAz+TPrMvpaA
UXTqQGlDOUOldFL8b9pwoTQHDqN4GaoCrQ0COWgeE7Vgyf/Lnwtvk2agnCKi
2kgDtQ6lNjGQ8ge2VybveoyD7F4et4HnsBn764Z8ERIfQhcaD1A/aaGLDeDK
KD/l7UAO7GhFhxlJG/eP9tQ0/7fia2Xj77dVGGsZxXvD/eE8YrQ5P+iD8NdF
2yqAuB/iBYW/lbF3BfkigyAsec4j/f/EiO462EqRLUCQwIZgd0sZE3td991u
3ui1951QfnclkF772B+GvUx6iuH+GqKwSVfzR+oFM1G0cNpbo0c8VvhklT7F
T9B6DX0G4MLHJET0aptKtB+hblvwKtrIXetp8J78berfA5T+05ZrOC2IVROD
97qAKe57fPflEcsD1GA6ICjE9/+nl5gsf/bDr8Rp1M7sQWf84V5DpCTruiTH
fxl5/DMUTlJtFMQk+ARUK394UyNQtObYjmCz8yxiZcQix9eSyTtjaGEi1PDX
TKA7ApFVGqSoNDWlz+RcPc+igUiBM0g8X8sAq+Stkm79sOdz+UAzCBpzTOnC
A/tOfTshlmY6K4rDJ3mSFTH27bIryEanT0XrWDIWTo2nvFKuCF3RVleW9ElB
aHvB1ImnvgSvDTcH9ZVisxHpr7tVJfbwUKfaHLmRPu/dFlu5BxcPEXM3GeN3
bEomCZCS7079etDIB+HlQ06MROMRrMLgYtzvR7Ir2sJ3R7K9ZXc5DWsxBajW
zhG6gQSkleu9k6uR79D+4z+d1jC2UblqGrgb7X1xWXUFt/XvpjqkFVi+4LSp
k07npDrjr0NSOEAi8tdozHkomqGJISze3Gk+UnD/2trKe8f9hOhWI4P0krGJ
IZ2zkuKCCW4u4FLqp96Qh8vNDbhiw43MnCMNcWKMd5bn+qgsDc3VjZtwSUj1
18kg4RJ3lxYn2/s2dU/JnhFB0P+87aPPRnvJfJXtlbotk4cb/0A6Ke3yVMZ3
gIE48/sj5FvkWptslc1Bg5fCEhYir4n47XDk0Fpc9DPK4wksjmkYBlCXRf49
0t/5rIyO1Owv0pvwJxNCnhHYQetQx+RBEx05Tbp7BpYzsrgqTh0700vWOfdW
YT+1wq/CYy2PEPC2vuU9FvTFONj476olPINvUSKQ1+fEZkCKmAvrZYSifrYr
Tk+3ORwZrp5muCR8UlweCZV/R2CGuCq3vrjGdHpoagOiSBnv4B9piRJLOElQ
IYBgsA04FPSJb9xa4rdywAmtXX2Q8pxoOPmSpg5I7khY6nRloeX6yfgk+3Kg
CXA3t0Qt/bJ4PgqpMxCf1scdz++cHaodIifaoKFre6CyGOkH7gppShzj3sbP
AMvbxC7ypxA59em1zqYtFZssIV9JAevluMKr7mWzOnw+OWqG4U70kqCXAZz5
5ULC+2dsZAFKIujnGGPYpQpItOIyfT5W9tRk3SLswFFwnGNMez63JAoXLBFf
rfYNPLfcCFixLYNcdpKMZro0BdtZQ4A5RoMPhVxSWSfLEQlTsTn94t5KTG+9
V3aUdlvbRB/gLWSErvKIukXlWMuGDpHYGp0oYoxKlzMEo2NVhjiiopAO8U+8
nH/A1AzdvTQe8mShgxKWdv8+YdAylg6Rws3hRNnXv54tL0QJPbk1eiIPMjMk
NJjIlXUeFfmCLATV4SyMPvacQm0JexyURVZTZJU4Oc/94IqAK5ak3Rr1ofCh
heNNM+94Jg+vjWx3jxC91eRjZwJuBnKbZR1/Daydnwq0MM2QVTSqrlP12LCF
cKMasMLQn86EyBzkYiBy5XvJR3R7VKw/PPU59Yvw95M8tn2g9CIyZmDmqwna
9cLLzdaxwrWuODT4IqMR3raJ+mSmCrOR+G8H0i9VualAa3nChufPhcLdQIiH
tU/WA4uprn4z1mDMAJabQ0iJBNKqu/gvTeshGqC4/Q/VbFZ1zPw5QZ9QLQK/
zHoTGKMUF+6SzrKOeS6qlq+Ao4XWwGFTsK4Oruw9CXIcsr5/hxzVl5r3Ta3V
h6pZvrtdWG6tvWfKmXiE8ZVhXVNY7wfB2G6FI+P1FdmNNl6Ydf6DUu618YhD
b6/jwDbTaetk+ILmrb9+X1nTI4MowXFmY6BZNRRoyysq1X1ixLTqMCkDbyhZ
lIEp3bp/EsFekQNTc/lxg+LKzRt2UwesCXCixyLw31k5sOGsfLsk7iE0oosW
wpA1cqIJ1VLullB5jRWwdMOnIe4LoYsbIm281aeO08lEX1jPPJdD5TYYDYkW
k4Sd3ryJYdb83gOtwsA3AnKFS2yY/VMIptcKIaSqIgXA0jt40dPxrZ/BZVeJ
+4fs1k5eCoaYWO4eS1VAwwvMlqRzjqFmX0rrknlOA5GnEnclmDdYQNCeAd1x
1/VfNfWFu5Ap7VjwfFG2lZ4KZvlOD6s2bkYIevsg/+a+WMGcvZNAy9DLdH0m
I5aQwFRWVbaZZARlnFQ3pMuRrtm8sNCkwIH39ndAtUlKznWDYrrVOv6/wz8H
coiKCKwuCamTDfhQHB+TLaXaVcGoVgYw30s8zpVEnG9lPCShALTUoPNPdZPd
uYz9yHrXDN1R4MojltUsWcFXqYnE+ViTqzrmoUjwGNMH2P/jqlBLOM+Y0qHO
fUOJ+N1KYA8/upQywk4r/HWRDp3IiveV1ilFxCSLOgW979DdnTobCBYf6OgC
UDyn/DPNa53sMIvJOgARM7FewaD+k8n6Kb4v39P9lh/sROwQ/29UV19yQGWJ
c+YF9p3AzALYODlwp5c9qXx1CXxfhWeoNOvHY6Lpu2O3fyh3nIoUNKp67UrL
WTSnIUg+eKJ7sGSJsX7bdR0ITaS52FYp0MlDVtRUNv5lzep9UtDK4f+rylMt
ZxZR1ozI3Gd2pI1tXIQ6KaxaHxs9BLS7DJjKx71VEkM0lFSxP9VUEgWiyFrZ
MtfxXtSf0w/5h+2K5HLzFDEgPUO8K3aSwuNZ8nX0MPw7sKWmbNii1N44gd6T
74SMNILuBLe4Mfr3ZAxxE+EpJNtBSQQiRrMCiM0EEe87S7H7pOX0zRHftdsb
YMDWDpAt9s2qtp29UeMUcg+CR3rsmF0PN5u5lITJp1rWybMGHFW808pJKOKJ
K+IFMyw4hcYR5DBVyusSyo/4OUETt22B3dTQ93M7ZAe9w8hv70bgAblU2wMS
z/HVp/roIAP/mndTKIP3riCsKBnomnsnbnf+dEo4FdY67Z5R2DpZLO6DEIP1
WVNGgRqo1pdifTDUsXdjjOwX8MC0wx0qeOqCCeral3mHKrRCOYBRb5kgiE5o
bpyiMDolMqwT8+fDiUOKIzmO2hfv12DbOMMNIXJQTRhtLbExjLDjW7pP4jDG
uCU8uFl1xMI6G2XZJ3QkomcGR/YrMBUNTvK/B6PF1WUDF9Eo++Eb6+xRpQC1
zi7+LE2tdAUK8KsBWGz8LlyI7ionvMTs3M/dIh+rIFryfSiSLRDUIFL6CxGU
9tXb4MnkViaOZJpC/4Ug2sqTWSZX+XSYSwe1txCEcIrB8oTRJ1RK0u3W0GNT
aruFIxkXkooGJwHa1MG+ZkSwrZZSWAezUfHmnzzuVaTe0OsUG87DsIXeRMLB
iVvqW2o02TlTljMIFJHZp8Bge5tvIgW0aKdZ0iQij90kO1yP5SiNEbxxHklL
zH+7gAKQ3tNJyZhwZFuIeBgAD0reGb0zlA1zdgMGiC7A7yC3KLPN9qMOtAh0
ZaVNTk/9A871BWwDQ7P9RSBdfKMWPnZiAC91H0KaINn9j1k9fBQ5jE2ZY0Pw
qfT2Wm+NFYz1LwC9DqygugpzyJ2/XrJByPy10nGe2uHev6zXwCcqsw5mNRyh
HyiqEaWTiNm7nun6yyxXRv0cmdcibRAdVOKiGZzbscVOHN70sfr2eYnA2ofl
myKQ2bHa4b8RQsFHVvhY7m9ur/jZyikzLouGH9gqnikGucWBRSUBWp5F+wzT
rkRpKFFMa6f4eCYleGaDsKf/0yp8GghpfKmOaWfXd3CTv0whtGhHoDHV/ht8
WTvL+fhkoYzFyVMriEuTtTkK7/iQpb74VkAF4nPWpfggxYknlYMbpC3KC9tq
PTXqDIJ2URuy1r+5VMDa6+LNTDFcfWKOowg8k2wCG/P35k3X5XZegqIvmdma
3K1oNhxDn3qRqNqWVOBsm3WARaPONhrSKtT+Ugm13EIOx5BqQ3Uaaa7XUwwn
VDi8/MXKSSrpCTUIFVR6VUjfRmV/PrbXPAp18B70vQgyFGkC0l0kRE6JMRBS
966emHkyPq7RTQuIZ++MAQzAk3hSFNMw1LsezxGdxv+DfZ5oYYSEZC1vKuO2
g34+KcYnE4/gxO6ZN54zZGfAeX7dsfxvk5B36GBi8LQz5Snxwl50rA0u8Ag7
w+mTJANo+QF2MD+O0EtSB8W/Y09tEZGloH520gtbAef4G81mzgDxzyrU5zjI
ItCAcSFk/pB3Cm69XeRMCo8Htlt0GI//GGYVrOkRha1lMW39zvWuPSQ0CBop
AtZvrB3HdgXprJ1d214QePPpfZXrn8jReYBNbuXQjGTWMlKqr/cdt2y5SVWk
/2wXpsJ/e8BZ/k3kqqRm0cqhgrHbHrZ/g8fdqCM1cdHeTqDnMzCHnY8BpVTe
sRaEfcMDy3RgD/VOuLQ7xcyB0Zxd8JsJbz8Bxd3+qBKACy5w8E5UTiFqYlC+
Z4BjyRYX7y2boWI1ZfNk2NW8eaNfvKzSWgKiZ5I5X45f8YS5n34Niq5ka74y
F9bZaZFK7Z+0UMuO4nPAfDiRMUYT5HaKX12Zh86xmGZPGh9BscrURZi/BBnN
UpLV26aIGpU4qr8fC5yOhO0aNAQ2w8hTKXnOhbcmRgiksv/GV6lR3P2R2IRI
IVWtN+51qvVNP4jArJAqlrSyqccVm3hnBe55w1O4uCT6FyXCwaa//loqIQOL
jdl7AWXAdo70VqWnXPhxqqMCSgpfdqLKZbx1ivp9TJLQFEKYrITFMwyvjc8U
goz8qDXbQxNReKve/RqbSuuaUAETb+1K5VKeBXBXklytLiIb73Icq9VOPxFd
DghVHBQK/Z+X+zGpjgwcbgvCepFpvFjULcYcWCCFKoNvpamIBVQsU3DW4GFT
wBfZh2SOM9J9furEDaB5zwjgUOvYTuTJT4OXcVYHswdE3x5Gwfp/Y2zszbXM
LJE96d8B2h6V4WjakrrnCZQCM50m+9t588vNrCDHMgcJfuLObOwppLCpUwJ4
yTDyt73XxF+viaWJoZQrDEontvSfXIDQ6AvXJP6hFdLJj9jAzNoeLgEf9+qF
/3MhrSJs0ShHKutmudj8YA1lVnHKTIcvVEAcWE6RVNMlVNXUnX18UrpkJMdc
peBFU5EQvbrIXIx7SgojoxzjEsW6JB7LFNe04X12uxmRwdtnoYhIxqT4/hmI
vAkJvpibzjQcTrOmVBkvCIHp3tDzlCkum9Pr1eqQrLX/RW67PQDPMsu8lree
uCE7t57dO0NCNlyP2CWxx9LKfcTjQpT8Zx827ACgSMbHCCzia/N65K2M3bZE
CHzgJGk3/hWSoo18uY6nHJ3ao4mGXEfK2LOG8M7KUKsji8H+Jffb5qmkfVXi
E+MNKNLtztJZeIf+pf5GolQs/hzLqes94y1oFYWh2T/oq8McTaZ0oZKN2idT
3grcTM9hdhaJ4pEMFIeXhM/8KFxLLjq1lP1u7XYP8x84+wCwQjEWcKlMyvBu
31QYUQh1RzD3oEe0BBnXKuxeY3OSaEtRdZOWh2U8PB7T7PxP+/pUV7e7rXoJ
p1HMgyNVEBdKYPJzE5Acus6WcPA460CJomP39J9tlRNTp5l4Ml5gvO680AyL
VUEX2j5I3jtjRT8wmCA/hheWxPej//UaHs8jObRmzQpB9g1uYkuPkiAPFvqQ
TdijXNmy+nRsN4EAbTTmBs/+bQylQrrvn6ocwnbd6ymlHwf0587H7bvbP7+D
DYZgPL14F/r1as0+U0BzdvSEv2q9JQOCVdLgrGevFVakocgqqhGM2mTCoWkA
etFN30x/tJ9vtj5lH/IEbQ6YCZlEs6zOAj2CFYPrO+NGAf/nlng4HKiQUAOm
rpiJrocePZLpoPw7Fm/Kd9kMYsTvn25UYmsfj/177dl0iEe4Z7Si28tI86pc
8vNqx+7/8ouOpbZoIZSYSi6LvU0skKxoMsVY//tZO4uiA44MCuCsbnm6Y363
2wza8oAnbDZPBDtM/8pw/3Titg7CykeTYyMfbmp7SOEtCBav4V/2U+jwPm1z
9HqSx8ncN3gxW+Yy9jqxN5/6Q4MI8EdKl5BkprdKl8V4qcU2v2MylWUHel5O
f26galymlUmQRN1SGp8EySd7epiJlnMrDeXz3VzDC8vspqneEp2NcZ+mv2ho
sAzsQM1NGIT5wMMkkEdY+lRBg09BPyP59ZHqiLgFQ5NuFi1cMHZwCO6i+R5j
U+Z0kxu7OFkcWasyHsDffJfsS3Ac2QU7oci9+z73UV5T3SlIV/t7wrCY8RXy
tZJqYayNd0Yjtk4t78gg415zKpsKLHavfIDMWoYS5O3ZPKT3uwvI9pSLb1J2
0zI38lAIhIiEIe74h57rUthxLqz3iGy8zwRCWNqpWv1dgdQCMUdYwJ03uhKx
v/yh9agnDZlyzgaj9uQLgpConS8TPbOFfXcFad/+545XeML9tzAykTxFmOn7
h6YKzorduNtdsCCOUS9bVL670RVmyCGjna2/9TloRasIAEnvTmrBxtApJahR
w0E6q+DHgiH9VJah2gcF4NRSbCbBvXEe1agRUe9jDgj2cw04yZV5cjDrB0k+
IfiARL9xI2L2N983Y+b03yYINk+yTuDTJlcK9cAPFIYb/0N4k7QxVw4HA22C
rrkMe4qq4o2TjO9Whx6n+55ddRR6zExoWVVGpfDYfEgGkVjjEn6Q2XVmXAqp
1Onx0eRVlQj4SPeOnAcesXmnqYLOMN6YlOia3qzyYDfzjSJSZO3DI01gE3Rk
9VggVCDerHz25OOQvdfLUTqZWxUw5MqI+IgMFGfJlTRwN6NdmFrx7KAZCOIy
Hd2OCGu9OkI3qICCMmlT3u4sy11xKwpccK8FnFjB4vC2NMxwR1+vo5tA1hNR
UDA8LqKgfjy7lOBKCNArxOzwcgao9aTi/rjyFKmY+ShsnWHBqivPLFWe/5ti
ZZJzGmA13NOqM+6XivTNo+8TOMzIaWoIJupTyrnR1n0+1fcN6DNQMnzzusyP
Z29sKWfrvqhJerxDOsohNRrSyJ7gDQ7/wkLr2pAg/ufxwFTxqHQr10o/Jh9n
5ldoYQlPu6CGy4sITzKxsJPrDeNGPMtY0QKKec7I3nvwfPhrMdLWbqjcvcLv
8E02Q/f48afe4l1pR8titLYE+fZ1qEt6dGB1qrlRuMUUyhteMFPivkXbLtyX
hGFx1t+Z4o32r3K6XwhyCc/1TD9UcDgBgEm3kNJYo9UPi2yJaSkOKggRCGPq
qTfOz5Z7jxYHDJufaulWJFoiYXEAyWpiRNR8Qv83j5WCj+kiz/kQpQl/Qcb4
9F2XZxEAU1O5Zct4S6H5/QxwcQrnUQMh9uYlpF3m26FUY/12QFq2MFUqQs+g
I1d6UKHcYhiBUx/9r1QFL1TqvSoXiOyd63wZagjyxeXjqyq0NffZh3avXhIR
lKgGleftayNzDkppIC4yiJ8w7V/yXMa9mFl3gEJk8KrjvGzWRLtU9VskDtrM
y/Sr//4aU+bbJm1i0HUMTmbPSofoioM6hsL1uGVBMpVOqcjRBYTcZ8f1gi07
k5NRGmz4B8p7vDPw8JgnmqQF+dsgAakhJKAwggruCmuHndcV0XE0Bxpt8zQA
MoY9MKLTTa8npHeu7zoi+xZ4doQtre4raKs18REtqwDg7biFSKCJuRJsbBr1
NPcIlFQ5eOJpNoX/6cL+34wkoPBVmonvI7x5WAE2P0D0bkgye5SYsW5vzU+h
vkHHnQlF54aqGzsL/BMDMmcD4pylUWHSRV4fZXOUZJK+7esDwrSnvClcOAw2
abT88vKQCaFn5COCjiJHlL/tUAJw8M7hs3XK3Bqpa7YGMkX2L9zmxtPGxSiM
d+LpX9LjHmsW91scVMCbRK8SrJjo2ctyk4GizFnBiWMEQV3eYTYXGNOUTLXv
KFYAvJKerS9yXbV2cD4w5phPH93p0Je0UiqOc/ZmGukGxNCKOXaN0tCKdTCu
53/5I+6FuiuqrO7PZx4KISjtyrAq6/PIpCoToGSpDWHSiuzHCaJu9WdFuSnL
YUeDpnp/rxBCvkOno39bA0dgv+4YWzHpx4iKc/GH+Em84ZMUNzUrCBYVhxRw
MQEe093GsxtP2R6JcvsboYU8u7IEJS/6nPpRKOf+kF02xdpMhtBtXL1P46Ex
5JBihl9faf4ZsGN+rs0EBYosjJeFwc1L/0GzC6tAhfgVZLWDqd6ixdhSb7MI
u0pK9t3YeatVBwmEKVwc7xxdRqH/zRBW8ZwpZW9TORLrN1xva7Qm5tLJbAi/
34gusGwJnkKSlvLx4Kf9RGFBtYE0+UESYO5hT7rrgNtMI1g9MQ156jJxGy4M
gaBU6jUxLHDIYyjmEVVXqNaBiTMnw9z9fvdTgKAc/nSjb5oL9hBngAhWq6Vs
g0cgmMj3tn7EB6GX0WvZjnXBMYO/3cOiSWptOcCorjMXMzICNjKSd404jF4j
T+wI/2TNgu9em8iTYuRQ6IAPzh0iWnfLAlxLqp83g1iWc77Z7p6i12Flm6Wb
mtfQRuuT03apNdtWtTuu9dx4Ay/gAJvOrEC4Gtatt9UDjgrAM1oEqltk6oge
3D49Vfx41+BHT9kjXzo99cH9a1kTS8ox1Ipvk5hF53mTWlaZqmEvS63RI3/E
T1w9w97eToHTc9YmUxNzCTY5dC0/fR6WRAxUomKbcLEfYQP/WBXueH6YWUR1
gaPvC7u5bT93NzzNZWjbIeKOXzy/Xzy5wghEXPlmVArKbth8AkHB44nD9q/b
+VfpFsJQMGItQpKqmwNh5GQxDhDinmJepqEv18FPJX34IZFWSwUjWVuCFRZV
aDAe+dLeLseP6C2aHIAIpZgRY3Ab2/4M4Wn2YD6PN/REJO5p789dZf1ZG6OA
cIOHggSwfnLCD3nLz7Zo8/LBvs4gOfqFRJvrQgavHoiilI6k1z2L4U9WwKm6
Gx6kwYsNa0rWoJGx2RCyGyop1p4LYf/tNTrx26O2eWeDDiihtL5oO6b/OfPh
o0Yj/tfmW6AJrc+dwrP6VKLMEhfYSJPcL9O/uuQHK5vgDKGJolAwN4Ke2G+a
2E9ALWT4x2fdQHoiNtgMswny6AuW6VHk3QQALkTgEaVBNBlrnIUOxPV+gbbr
NY7FnaD3gtpBCBbhRB8hIsCUon2zPpHPmoXc9ka44tIhcPAjx/EKjfSkvG0u
P0fFM9WFRkftlFHYkOzsOsVVzyD8hoGq44m0O40KfUw1HRA5uba9q186iFI3
AjtrU6uBtZ6AobiYTm6oc6LrJ1IHGvWdfKM+kmo2XgnMVCPNsOx1XlmRBVIo
3Sh4JYBUq9JskNSZ0EWrzXkOP5JRNBzYAL9S7Bs1DsHeKYgz9knd/mrQo045
YMP1oPka5GFufFZJuHgyxEJEkViXhIEPxlasrrQpeulpZuDH79Heh0ZmvDsp
7XC0C+D9XlRStvjdgkee5mQ3d94yLQGVFFY2fah3LCOl67ZT8ckIrlC9CgxA
6WUwbKj9tzquKj1Lw880fxel80UqHNKX52UM11AKRW/nXWtsM5+O9p9XQ9dZ
gq97WbePlV67HTmJbCUCdcaohIDpN4ihQJEi3qSRBvzotHXsG5cZaZT87lGl
1hkvb3gmG68ZSXo/ChmFPk8OoBALNI9/Wl2bk/doWHQE/L/Cvmuzvhj3Sl46
gx2E7/WiYSiQJAbK1hugG5pomP/Ah/4HAhtXwdZlDMNMfV6HLYUSVidMrmje
ZfPX0rbwSucyat0onetleGZMFWYQ9bNRUPsJZz0iCYH5qsPe65ClTuxBwW0V
acNtDSMHTf2C4Gx6AjUl8jj7/2fZQj/YbGxHbWoz0zYbZvaoDgQ2q8AmwIfJ
auS7C/zB2RwwAZlkJw8ajoNtzMoGNvleqxZJm7ZFZjBx4AO6YMV2hpWCxfNu
DqHn4n5XcnEwF08ZfXd/mbMGklibalyjB9gtXkeSJw1mUMLd+ge0LUcdBqlZ
zvr7nS5Xf01Qa59ZpUdG1kFeBykSjUDz5+i6l38LhTPoAl7t873Tmv0ageOg
7hR2qIoQHr81axC18bCJsCWsRmTvB9bBcC4VQLYqbGJ/FJrKDD/5BqQ2XRxf
abIQ2UujhnuK/zD69WjYNOffj9heCjHr9tgA2yh50A3WFzsSEjfSxrzJQBZy
vS01+E1Ob2j99hSQbcwRe2T5dhc6GK/Cxz+4OyEZI+CnQV+Qc7AsQscziQVr
qLBFyc33Uf0kpv0FRlrZ/7lJJZsJ6rQ+YDs7sO6JA92eeApzI6uYhTDrokVz
JIFgVmMzG6xNkPWjaLLEjFB8oF8QXsEZ80v9EoiIbfczXLdiK1oYHh1HgfhX
Gq+dXWE2jbWrLREidhDvD64qqnfPseOUwmXu+3iCioU3Q4j+5e3Ahz8LSIzs
IYN74FAoQWHIGzLXb5xGYqvc41LQWJ6apVjpX8Nok+Prg04RuPyGlf8AhElW
rIWx2+Vpn2i4ecWjamhYvVVmiQTrzggYsoZNnkvtrTu8bYDzFQSjV83v1ol7
Z+02TWfX9jXrY3/KkH1wkhb0M9BKDU6CHNOGDx0lktqxhEPJBzs/RPOHyqSk
H3KElV8mSseRY8pXepWbVNKWbTgPUephUPVIUVIyGvJsvAGN/Kg2nnUYkiLZ
SMn7A4epIW/XZsDIZrd7acwFw6VmIVyiCicqRkIfg42nAwELp3PohCrEBQHR
/iGeKHtl2LwE11gOVmqJ1x/QAKO/QzyXjtQSbAxCYjY6cQ3sB0yuHKWuGhcO
NAdma23g7QJ1WyeAwPIvwblc/6/NcW4i/u6CjHhWk1CJlmcK+IrsHT1iVXGJ
RKrCszvghAK3ki0PBS+efLslBPT+ffdJFlx90+pAEFERucVsxWhmRZt+PuaT
S6hb1XDvpdZ3pFlfDWSwy7TEHk3pWTHU7oaHHLiowXClnMWM0Dwk2O4YMleu
iZ4RLsnFOQ2ykMeHVn3ac36rWEIgUrDqRXJ7EVj+YCaL2qhhLKzYh12MES1K
9oDeFAZqMdNklZ1ckyWuPuXVTmiWOgtTzzqFusspLmPnHESkN23QCiivhi6u
hC+3rdMTrScuBB09gapD8NfqO+14CpNPRbw1XjjEh/vqepVhRCbqIsJw6EpF
rR6Z1pN9ok9HjysxYYCxj9ITdarWL4JonhzY8jMnMimEbD8ChlQa2VOQwNS4
7su9V/AYwUSpJDq+pQCO10c0gLSxDDh8kuZmyXf0yOPDSPnH+52OR0IcI0HS
qQ5HcL/ByJX0vBOZAPmrBnpHeh+PpJXIHy+wJZNTXsh45nprIVBsJkp1XYEV
Ol5TIT5Hm6klr29MB/NrRjm8T99Es8aYNSk7YtLlo2gIz8nO678M9H+MIc68
IQebTIUIW63lRCPqiPn80kXkI46FeSlU+PcTkjHYqQ7ffp6AB7Kh+AfnkvGN
7UvPbiRmfLzq/TeRNpxMx2vpcO8QtwsnawLj3aAg7FcWFOz4UnUI/PwrrNIt
T93do0AqHPQAAbUP4egrYVw2G9t8vZQ4lURikqnPzX4waoZ+CBQAdk7Ckkr5
pJFzF1kB5RYCKUNIXBM0uSMM2ZviDfHG0nU0cTGJchfUGyjcp+VUv+hXRpQt
Mgyo2vBjkGC08cLcHjJMxZlNAnd1vIXC7QoYpXk9EuG2NAR1iQXjzEDt1dWp
XsgjFra36nglqoezHQNS1cNY0D63uhK3Q9XgJ+8sLbOBCaCtU8d7J2R/8sCV
5xme/8awh05juoyQsvxgy4uIPcu9PiIHiCuhVW3/mmjwo1jbmv+JfDtZe2U0
XjqpOPO1STbjcLSkCFwZ6USj+LRUWUHt++i5/2fd4dvczCAl9tBbP3LBUQ2N
QWcQEdCa6rXsx5fxkujGmcU1JsJu+xnH8GEObVPw6ZbA+P8yc6Ds/8iqidHB
dtwA4STQVfFFJ+VZ/BnuDgE22ZXX0msYBN6nrY93xZE8Ha+08C5LUZzoVhmr
CBKwa6onmPekX+19ue8pCTIDTOY0JeHlA42/tZYVvBYVGqM89GeJhW+y9YHx
xhYj/EFEFRXBs+w9RcciUiGudXqplPO7xYXUj+OKpFxkdhPRK9QTG6pkd2NE
ctfkHpa/vGjzmT1y7cOS7jD8cUaDCbnXUn7o3RXsH1ShnBShqYXA1yMLRGku
5f4K4VfN1bH14GmxqLD7a9tedDmg6nD1Iao11lB8jjO9QoL8FjoWVA7X0mIp
fnXcawFz6UrGI1nfW7H3y9z9Tg7LE1LeiXM3hNunGSGwOiP+AHKzZdz5Y2ME
aTP5EqF9UgRte68H/Rsacp2puj9L3Jo2JHFtD9C4O1GSEamNVaA+NuNvE9SF
PvdlTcXQi3bVBLetNK7b+hKdgHQfbZAGPZTJjVyepBgy9fF8PeV438bUuGeR
wtZ20SffdwSKLNEGKLn+//RZbKfqhiNwYurAVumc//1aOvucAVgUtTcrvxK5
rrTVQbH8SolkA7nuFZc66hgisY9ClPcQzEQAJJ4yWC+1616QL8+MefRqE5z3
Z9vuco2j53upC9uPZ641CRbiKh1BJ10RxyeOffcAjqydcsf2iQbKjxkiQsCy
+2ZDsPW7ESbQFtnnPs5IEKm0BeQB2QxD0N7lcVW6rvbRiRUz8L+n3YiS+6/c
79xnghgfTrtMjNXk/UIVYq6LwfawYALIQHQHRus/W5+YHKXEF9NBLCO/1Jf2
M67nAqg0fjGe4RIi9hMmlO6+9tNn42lrhGdlcS4TEYTsEeTJzwRgmoHOO5jg
2fY4TbD7gMrj9rVtP9Dz9cbJAk6xqqJMkgpqelCvCCx/c2ao9Qxr78TLLAvU
pFP2t5B4NcHEo4jI08prGxB+bFKF5yGcIyjfLtTVTBUjrdUAxZzwhK8EA9oA
qxB8jT5xuJ0CSkxeEtmNhDEuubV8o7XKFdYOiAaG9S+HZwNNCyiLxmsbM1z/
NMqBL1uqbvUiDKDtz+UHKHgS3OsMvOI8vX8ef/Gpbll1b0xAjfHwEEnHMW9k
oC7DTfRZFwoZ6HxZeyxTrCX9qhZLxtKcIaCzCMQXL2lgedCwoc4Xc2xsLzko
YrvN5pILThM1DPV7j2oCE3cGDXmbmNVHaLB1TIA/ysVZhMc61HCkFxMNv6Ov
p6Qeyoq8dpDSMQzBzGAGWL8eURc9QCOb9I0c2vcHqSsnjmfGUh3QUJGwwsIk
VMsJM+CVbicZjOlDurCJnthjelsjPELnJ05I31f7nLW7pxe5VFLWLonW4Y0t
/JoFYE60TfplsN6X2Tha3qmVeg3ur+oRLsM/eE0+QgkLx8ijyNC48Ow30uYC
2DfTgWOhLMXdLW22nfowBKNBcSFifXHD1ja6L2TNBxtquWu3ROCj2Hr9oPU4
zr4oOYpmKupUwVs+As4taaUSRdCjgFm3KKrPoBOle/3P4InFvJNXUg6uRrT1
0IHsJ3HHGQDdi44Wm60tgIDcXMV5yXsS4y4hWBVNzrnBrhvlv2Bx4NC+IHLL
IHc7CSWjySCW6ZXSYvwnK/Q5b1bm4RVhEvR8+CG++sPO7n50tECZyaN5ccnF
79pHUFMr+z8kp+4y3fDyJJ/45EzGtNYgD5Z5fKYyOr2FGykHmmy0/tWCRI1+
K6jH/Q54gitQMwXqgWvRD0MCJkN/pxO2EYxGU0hAr/WtOC8AXfWGOi5nL5VZ
sIvgV5h8erDy6aTdlMgvmspak/9+xcT5jXAkvL/s8d+iih+dw3YwQkxIF5+A
cDEaPIFU39/KXePKSgSasj9aHSQDPG9TyrQQB+aqGDRSXHoR1B3LzI/l7XqI
bcwX5wrfY4mC1em7IVa001+Nri7cXASW4AH5mLc68N5XyFd9Z04QY3w/VYzB
GALozu7hK+HwC8Z5eBvW39Hu502j3eViOc6pXVl1Di0rNAZIcNCBZWxUtr6L
uwABJm0yz9y8JURHX3E3yuCM/v+Uo9zpWP+Hn0I5GIl0nzWo8b9qQRK4wT43
kJFlvHccuSgrIb5QcdFKwTGAQXU7nCJf/ElHwR0ci/PotTvsN13jO01R61wn
lPE4/8qrITZaSzC4lO2mbe8w/1etTZNADuhAxpAEtx9FJL0+4OkVAxAenAWm
EScvLNR/aY+x9b54Bgyrt+VBC2grlQTZkdEXrd/r/z/cZvErEjT0Hoz4Zf1/
+gh15wVZpWYrZbHc9a2zjWb8OoNq3yyr59bBAoU/1cIttyn7S4sqEZg3x7bE
oq6BUT41Ac6k6Wrs4+oed2P/iCaV6N731e9rTWjpBibYWA99/14cDTKdzOh6
ELSaHE9yql9HPRmlxIfkI4AkD+CQe+oqRYWrQ1ERLsKgVTbcq20yc/Z7VSRz
ZObEPVGyNFhXeSfCxOl2hnsyyJhcBqycTmVvAuIx6leouq5vsCxKvsuKyu++
+sWF535noe8CUVNo3ZJjTEWWWrkL4WDs+3Nu7V0hWS1D3YifnRv7qX191go5
jwzRrCyKVM6nIpcmDFDOfktJUWtvEzYgBRWJxtGx0xSW8xZU7vyCmCaoC7Qq
+30s3Mz6yCueobmDlwYQU9kr2ErPYV5Bhe0PhN5f43eP5bhFNosPOWxayhSh
dY5datECjRHC1coIKTi/lrhucBp+e/o/urFqkKQwNHR+9UQ9a0GVoXpL5VS6
U9hia4kVcRaUl6uj0WmkboeDkDJ6/7VOD7ZeI3J9E03/n3Ewl6gMPSz1Qqz1
cCiGM3E9a0PQ91+dE/U1QNZxXF6Zu3+X4z8yb8GsEQ42EV2HhyonozwzEm1P
vmuQWbrxSn/MN/MSExoroPf60yEow9NtcPNdMjl2lnQoCtd7Y54CIiJS3tmH
xUe1SHfNK9g20PJo8nSZDdRcoJZkOz01MYv5GV2NPjyEzO499Vwa8FyfPeE9
3KZCX+eTSapr58kZN+KInj4Z9HF2txBGjsAeLihYrO3Qg0FRoU9/8+cPuwtF
1JCumjMDWvBbwoCerSk4DesBsd7STsoUHyd0Hfd0zGV+jdKoNLQDi73UsFxC
E8qaF7SbSYvUVnfytomevzQJhWemq8K0/JNSvR03GG2lZiDL8UwRRE77w3Gp
RCiOfcVqFZyqWmGYy0PLQXjYmDWg5KfZE+A1loB1KSFWkP/eLRIw0+hpfkES
mM+XSNZhZcyvFv9jHdzBm8IsA8piGmU8pWl7w6C6texpPQaYz3msXJkutYlC
xuoTw93gnyNGU7M4vVy/8fvzw1YnU2xO8fcgAk5pBCfTpMtSS77IReQz6Ae3
+HNz9MTtCfDivsgshQZATetDAxqF6LnvPXzn6N6GbvqIamh3WJnytWDPawKE
3MiMC/+PV6DVESbGl9AuO/iuKcyBF49HZqW3MLUMTxzSvx08zcdI5Q9CevhB
ldymeP549Hj8Up4oXcMS0PR7hu1LV7ZkW9nmgdbXgCGRyJUE9t8xOLMHtbqP
Nqv9N83kAyEKm4ryoHPw8riGECXuaaw7gVcXNBAKb59mNwLuktISNxSnsNXs
pBzRcQMWkoS+wtBP9sPtKEcDOyk9ax/3tasmQM35f2bXHbj2UJv5cXBgVdRO
3WA95aioUjFJAU9DNBcVNkyYpUNP/xb0DKcP9rkd3cTZ/gS0axSQ3/006lw9
D3z1lkYG1TdW297V7OPHwCmGoxVspD2eZ1gL5WdtTdU+s6v8JnR7esN7lJ49
S4pdi2Agg6poHKLFpMg1wefuuogQxop19x8iiMdWnLEKpacsvrBygAGi69Bi
s82dkCRw484lMwGBpOTcBl5W1i35PaVmrRzAmyZlKydUvMGZ/ane1i3HufJJ
QMv0rkOC6MT+vEPlFXTaWqOlnAXTAZMkAxMz+RePHfd+TBAkWmIO+bx1hYxg
2tHhpnVu8gWMIzgpDTCaJjS+VSda1SofT98y9uz9mtBVrhRu1OYjPuP8/Fza
GHN1YfILt640xv1bnNPtmskEU0ht4lAT7u2btonVrAIb0XU91XVWBsBRDzx9
XxwmA9XGy0GS2Cgj/XWIvE79RLrrUO7kem4MyU6OywYznir8yAWk3aaYrHe4
TOlnc0SlxQc4LCA2J2sDdV6pG53hgKQXqdGeJnnF5KSacLmY67F3rv24uDPa
EprIdpjNExKNuGyf46k7RbCbNfTg4SwGAV7Nt8GeThsV9EUbyIBc/lILQn24
CqJ+CO38c7DnNya+SzHVMTsGU6xVvaM6io5SQ+G1WDaSu6qA9b/xEciaJ8N7
iOHGMtT0s7DNiml9KJsdO1onGkxUsyje05CFaOQ4JTD24AUhmKWIFoD3dSf0
T5Ba/l2BBKqccrIzFdeny5TPat/z8DNqU7U2HvKotn3NXi4XWU9rd0SO/akn
Tjf5DEkakPqtkR9cm3IMm/U/qLvf1K2u4R0Kz+vIZdY6WjBUlV8uGnX/2CLS
h+dmSOegKWvzLiA/HIHBvjWBzC+YnG/6wFVaIiTzvkSkxV7i+m0GFjMmQMtN
8reEuTZ7YYGC9W41MCg8swU7lEx5lUzm0D1MJ07N7iU8PQ4B+dU+lv4e569l
cShu2YyyGohh5YpF+f+Mhhwnx3gCLAc7FTTs6Nrw/mRF3IVEZiOTQ2phqV3X
UKy51izDAftTn8YgqXiAn29d/BwPxRE5B7rdZCh+5kNnJIq1IYwaly0eWcms
j+v4NzrRtCO/ELG1kUzq85sJAQ6ZeSGV4kmmX6qhMN9Q5ep/eyp1SEZ7ls2L
yjx8wSgeRxNSkYQanIGkvU8f2MMZJ/aJgLBUTF5UKMsptpZKyIFpaRoRYDyI
KymdALQoS3lrSRA3Umh42kle2mj10VOEQCDC67oxCzVVdNOO4ioVcWiTv/vF
bMzAy+1dFOuBulQeKOC3RDmbNecxsIiqLlNE+zzS9fLeoDNRXSbxJoBTCXvl
951oHDTt2j0uW2+WabAhX9Fn5rpRkjP2INab/qGqjZ1pZu9v6ChMv0BPKeU7
695w3Qckc+EJGXgiUsClZsAJW4RtncbT89tFenffzm9yIqLJHGb/A6q/puYc
4vtAFeh4erYwQ3v6uBi4v7Ve+Ug0oLBZFhotYvYKKqSSGTmn4TuxCmBUEpBg
FB12QB5+dHFvsUELSg9fm0VV/m3fp50qrnWFi69emzmWnLeedFwLmpDdQ3K4
NwM9ub4oE6HzsN5HJXXrfHYIR107uKZMxKgKGb7wBREKkApA8LF0Az+dNaaW
ODmTdd4OzXzMJDIcq59d286UaRqS3d+ZqPwX1eAh9JWDBMfxbA2i03TtkK70
8HXdSzEhuGr1sYZPy6MDQBoMRuLja+ENgPP+8J6fkb3RGr5vUc8GHAq8nUT/
tqmSXhcUlRIKcLHWZrx6z0RLaKtHZreS6g2sodpzCu2tmG3FKCB0raFkjWBq
MZAadicxmkWX4ydEqAClt7DNNihxjU6p3shsKw/ok1LgPUxurFItynoLuh/u
VCQJA9HyYbaH7aHTCULHZjbnu/8vhHnchXjuOed4Y+ph7mLAj8S28tfgmIwT
j/HVIYiFhixrhL6boJ832+NWLmj6dWyq5wdiuMjyMw7geoisB4lKagUNPoZT
Jnxae33Lu1gltDwbr9xaa9OJgygo9rkTU85YpOZBihMoTvO/MgaltnR/TgAn
Uny/Qnhc3h9BwM8HvQGhDe3sQgachuygseInPJU7aVPP26uSqGuJ6gxp7C2T
LGSTOHFHsb9KdpCXg/4hsOlDAjkZbTwmhVZ9OT6USnQ43EQcZe5MuO7cDTzy
XJi7JtXuSfY8LNZ3FW5QbVin4iCUvbI+VnKguR/lXM//Wdq6ftnX/hQld7Fd
ssHsSffwxgoqDOuRNUkV6qLYifO00DDYm7hcJLUlS8VHZ4PF/1kr0s6lXK9R
iDvLF4RuKiZNEgKDv3ppwDnecQkjkscSbi6+VvI2nw+00cxtYNs9tVP5jUG0
JIMnRfsy/DRkJLHyA6I/VSULR4lZi6blk+dzCiF6YiF4VShVAha1seYZscG8
5wBygXJnKKGCJYoAjdJdb72ySYVL2uxvvPbMdi1HLJg8coUxBw9tU40jfOE+
XSdiG2WqF+tpsUv79oqIF5q8horIu6W3+FCuOPj24ShPebeJGJG+S7aF/0rr
jflz/gIIZV9HTKTl7uR8MKqQPwcfz4ooYfqFh5cQh/RMPZMxDKa21M7RQnND
zkdeYTIhh9f/tGlK1fl/XscPRmDQRPF88S2cmEO5JJZ61jisgghWXRnT+TXS
j6tuHp6AZDqSIfs0Q0o54Yd4gdFehSvjwIiwikPhVw7BK8m2y3sUxNradSef
WYSrz0Pseql+z+StIn0R19QwP++uojkPB05YO30tJqhtDVPZqqtq1XxmNf27
giuR9PU5gUErQ5QhgZkAUIyg73r/BfR50N9BLkbCoM5aFTKc0cKewES+Txse
V+ixYQqVUp0rNiwtyu1ZoTJ7MKDaozlhEp8E7zAdOkDRyA70jyQPqqCEHPdk
BFP+217t/8+5yZwdPPRbCiVJYemtSdwQEdT1lcs3zL4qdDvk1dZPAE26HwnI
Ps7pdwogpB1LZfsKMDIJCOH1a2voYe4mlgnNhfBhLcVoTF81vIyjN35oi+BA
Sz+6j5ECItof+qFNefgSonsEdnSDFTn/QYzB761HAaUgwp5tExdctRY3TWc1
TyuxXjJg1Cb1Xe1hU/7jp+OCdflf1NqqhppPH66/2nSdXFdOqrjbDMZ8m1S0
Rt09eHSlEF5g44IAdgF60vWRTvTamkRXwxBXPUm+igIUaRRcIXVDGR3dYc2X
2gOLHLIdCkOIR37+rf6xydlo2VoJLVtPE2wXM/74Md0TLaHe81TCoKT2gnZO
NHXQ+BHinZIps2NosCUsJli+pn9T95xKUk19PPWN95h9COnrIvQ9r4+V2yRQ
g1O2tj90eKK+2Uz5Wn0x00G6GJ/gWovH54a2tQ3lSKusfhDr8vnJqDCh703Q
147uzT658c2/f0TAoAm+HhNUe+zMxBbHMb26/dEIUdD80NLOQDhpRRnCPvCo
FIThspU0EVQ57Zd2meoBcvuTqr3vHwcABBbxEPSgfWkLHsCb4pkr9mZYhKHd
da1FoQmLMWo6ieY0ALHQC+WsGcDz5J6JNELFDNCbDY+82V5Jdh3q1nO6Zad9
gg2ndTeu+IT4g8L5bSrwZtbnuUxCZyicyWOd23KDG4LSiLYO2HaP5nu+JXXj
u1plBcTK1MuYoLUsqzSuSZx/rZJxsm49LMhTSxgEyJsaooc2/TymuW4OoJbY
x3nmUOqhMWZnZUK77WgIVm1fZ+sBfaQlOiupJQ1Qw8+4q45XU3zoXycSzKIV
JA/fUqI2alAnmWGzlQ0ZKiNM8HxD2zhT6hkIZd+WHninUHx8ftkbsZx6ybbI
Iz3FvUoI6tGWrpbexjrn7wO/9AOhukSbwFE+Lyfr49ZbKIN61p8l0XYbm78p
b94OB840yd1xjJOnvPRIxWl8UWVnS3BT1deR5R95YKjhq6gGpGEZWvPSyo7X
o8T2iCzN4Ip3VlBaV4Zhd+N4d+3A8Pt5eORzJTbGV4nf5mFiC+Prl+9U3Bm6
UgsHOidTrc8SePnDci56KnKdSoaHqt4bYe2ifP6+ApY9NrCZmWf7nwuBQj6N
FU3WyOdvLLC9vrtXqyY08HHEhVKdiGV8/PP2PS4L+isDB8fkSJnRydqA8YfE
mWIkC3i6cBaIX8iburdOABmuTzz7Qmup0Yc+CT4B7FYXyIC8h+/IuaHunDtZ
stf5icybZiM4s2pog6QJs1oZH847qPI+Ji6vd6BQPqqRUcwxy/NwbjY4Vy0M
TQf/ZdA1T2Kb99Q8YIO5d4LbFN7j98UBu+djk7jViq/HIstRTizYR0ALEwgF
ZI8OLEEHqTR8Ttc+6YPMr0SpWOVt/2nGEb3MYOTjGqFb1jqvKP+opOQa2cv+
HW8qyULHqVPDobxw3dwiJEmVwK0dmv0ZvBjwpLbIRx7Xg3y21t4gS8Rd6NDH
QIfu2CnacF+1BApAfmNxLOD9sXbEnHrMWTLLLGe7rQ2tGawEbho0wYFcrRLw
m79fclfs+49APpfJmZxGQlYvhp3PGPu2M0US7ho7bCf3JTXng9GwtoRbAhhC
YMm3tPi/JXBDyP1YB7K7wN0N4bbG3D+Xl2Wus9u6iN54JEvifzhy+jFAc4xw
xBTnfcGfGthwG9OU1FJxYqtBVLgK4QOn5Qlpu3uSGSvT3+MqB6JycDAUItls
Mzm8kRI7mYqwpchYC31HxIYyR5ySjTubhbnbZjNjr+wn5iTwF+hRcG/oVlxL
xz4Sni2m5T1vAFhniHdrQwjSNKJJFjie8/vwNrkq2o7OG+mN3z7BLzHG8jj/
/M8xnpSX00ZR/3rv/XGuKDc+cv+3yC135AJV3SC07jrdAM/8x0X2s0UvxDN2
Fj0j/nN/6chz62N8bq7qTXJRMang6ONXZA2evZFZpzo0jHLo8ZrR6KpeD6QK
N72xq4QajVaq6/L5aqF4JjMc/BjYGoUwWn2MSTlKyebi/T+gGrHd4rbTo5c4
v+zJoIbF0gvIEynKPmkTcdQLCl62weyH41o8T8CYAtkLtKiPSxTI3p8ShHgO
ft0akqPmC4XBGY9+5Pt54hfZHEeUOj9CIyiwkgKFw6SxvL0Vb2Ni0RMQkUAH
Dfw70jk/V++FezwYCZtd2yNzX56sQmCsdZC8MK08CTdEvVowoAOxJn7J7hn0
PDeYzOZWMc98ySVm5BzGNis4V1iQfN7yGTspv8UEQ2AwxzwYdXGBGN4p/2Ow
VcqIIemoVKSg3Riq5w86mnn/LTQMy9DN1jBxEe67yTsnDrJh7jFs4qR1rNDy
8VtHV3GtW4YoAwchMLEJRSrwL2ICySyfCasnxUOfs69HEhs8/dS5gh56skUg
6u2xo2z27LMMwbVYkrRXgXobj8SxGqcewbstZTZuR10vQG9qfc8EPdydwVUd
Jd0VNVuEH+z1zOzFtyUiUbQBV7+uWB0paLmpWUiYVz9g+Z1WkIVpwhR0cLnf
r8NOUTP+cano9SoRgLnfUfMcI978sUnRB0FJRhSETLfwFtHlUAZrhBO+Sfrw
twy9etg3VPQEQ2OvCh91pzwTCrbD594Qq/+XV+wECzaCXryu5oJwS3SW19Lf
JKzIqTt71EggNHWuPz/hU9758cjp+tHiFtDTNRb1pwPKJQGe0v+hIgbrFQyP
i+pIo7S7sLFw6Kg27FNYb2Hw2fWD7r8AjfMYzeOmIqH2QDkQtS5AyzfZisG5
Z0nLNWqqVAJG+8B1UQ4sF4wNAVtHv5vbYnJjjqXTbNFvVNMJ53r5lErg1/VZ
8rNSS2NzhiUk+eV9pkhsrJCNwtAscPcHiXRrEUpmvWtxB+vckqZD2rREwR7O
9vLQprKe3oTccQHL4ZY7RBJWILw0BIQKTpheBMsrmLjfij6Tu5EwRERCRNoG
rxIz2o44aUbgkGOsBDCrNYWllDG3ykCVzhdovRUj2LoUCW4KSNPx5HhFsmiE
1Zg/oXEC0tLPfeQG6F3JKUD4RbyBOKZdSBSD9NWp+cPkpgrMe0FLQ4YU6tqq
Blizr9gTQEIM13WpebBzTZnMMmQTFZ5hudm6l8lv99njSJ8182lLYAf79n9J
WsGheQapYfbakqdAzn6kSkyPrJ+2n2PchI5qe2IXHbnVw5mhdUa2LPfyUya2
cVYdmkLJ1F04MpoiMhJ+bFlikWaCDjUndGvgx8fJ1dNQuv7ieadnLOYDMn1H
jtdkRCEl+PAK/W2ORT4BFoTClhDE0ZxkwyxjlQabTQ87staq3EE/Z/Wk84NK
LF1nbYgs6W0/rnpkpZ4MYQQ/9S+nb5u6CM5j4UNHcHx+Sx8i8vPkjNNq3RNE
cZ+fw4703T1+LJAzNvQgADFqbFrU2jqaE65BymcYZvs+Y0l6PUifVArA0PvY
xFmTMF3/n2AezyBAzw22lzw0hgivys2MHU0Zzl3cVDsBjZYM8hEQwalnv4m+
3p3BBm9cQ/tPrq3vh/PR4o05ToujgpYhPu3wYzxQamcllAVWNFXEJ9Zm9lmt
coDkA/vtzIH1VHzHRDIBntVYRkpZp7Xe9rK/nVMoj/BOQtatLe/oWEhN1Tjp
qaP2M66QVMeOF+BzLEUfSJOrdNaD9B8AphrFy1T5fDbgpfqN5DDu/1fxD1wZ
K7jTl7Uy+h7q/cKwNUcBKD+LJk94kBIHNetekrG6lekAw4ZTdddZYv/Er3WG
0DYpKfLfyadRBs9E1dhpoImBnp0V4tX0T4Le3Y0qylnaQwolx2xqeqqK33OB
IkYeESHRcuVzwbRB44gAwOTFOgDWtpf0oTC9SyTu9oaRDw9L0N5csxBJQKXD
qEiHxWkUMtGEuhCWOAkcyNSi+JSR1e02hhnAWw2fatW/bDyXH61XE+XpFO0p
SVtBa54fY9fbnHl/0wWFnvX5ymDbRsB16oBDA7gRi2TUVIhPIwwEDosn0m7u
HesPcPHb5UEwF3oCnjGK3hz/pUyfIwWPUrKYbZcwIeG0R/csx8cppF6He4Bw
fVrQA2dC4vGgViQL0Dq1jwV0oYQf8eFBDcb5dZ58HPd8Kjmftkf+q/ZG5C9n
zD2LrNcQ4fR/7EqBsWAv8nHpP0XHill0fjXJ454NPO+Cp6CuLT4/PtdsCDrU
+buu37eIsIGFz6NjroGy6EEBJF5/sA7QL23HdThjrs5ADvYladrAeCPTT+s5
S0O007f8j4s9DTm2f4PgdG40DM3vElBywNuRzmoTIpKxCt+Zf74ZAhFMM+tF
2hUzhXR6OGSxlBdOsuKEi8A7s4LXg2o3XfyC2z2KBIVYU30jHeXbdEPgwXME
YWc+9au85eUcvQxwo/mvc98CQZWS+AwllRP2EdzU8zVkpVXXeNt4NRwUEmZX
r9vDDh4VwleTzG/wgfYLiwUsHMRjAlU0XUZdCKFS/3Xdv+o0A5lHL4aakrR1
BGWEOv70MK9tjLbSU8f96DCl8n78KfaexU3wO0IdrB1SvWYA9eofT+O1jU7A
b3jJ8M7M//QEFahoK9kfyXe/Ml9uLouHer5LqX+1KXM9n1pdOF+gn1FDOQE7
VLo8aI0KBIjRDuZa5MR3zD5UOB36DCzc8yZGCOsaVukk768BnZb+nvrgkfPO
/YLAisX2d/hMG9KWDj3jdRqyskWYDI1WugP1hw0GytDdR1GVtiX/Bl3aPDtK
hhMBv+vg17scRxrm9RAuvL8IPJaRR/OHZzwfQulWrszBiVnY1VeBvUZuIX09
TMxQppJPDqEdH5zF600kir/Oxags2pFu80522fCwDkrcKBex/uk8NfcwGnX+
nthqVHh5Y0fOkFOhTy5awfXVeOZv0jP7St/Zuj7PpJidoKIv/kRdxg5Qo1hX
97p4tASEo+HhC4SC1xTPw5PFgv13zVOXztDgH0u1WJJtRXO1ZAZgpVFwXskq
/B7Dwg/N1hIxbaiyhXfb6kZ0Csp8OGTfQYQQnFobN8p+aPodpZAClRemCndQ
qW6Zp4fzWxEYNYJRiDO6tJGnjEsAWEZTV3ioVzrjArlA02yLtZupmvUPFnKl
fHDukG1f2kWPvNeuLIiuR80hP3umNzxbu9Lh0/4utYP47B/Piww79BPXJU2Z
BCY9xKBjW+W9qBy0ujRlo4b9NeavgQoslyFvHuyIIA2OXRN3nev/YfzaTkXg
dUyD9t4XYYezA24pGfn1ZeNMrpOfkwutrvqmNaBjec//rGUiYTgYNgaQ8ayO
CXfZupf/CyNhGqsxe6JfgG7NqkIJfL0hQApwsboXfKXMGZLfSR2TMODpvHpU
ayU87DqV1jBwBVzyW/ZFoSUCmkLSAcxb4QPHXV4V/DCqREBoXIyq7/E3BlTq
bmeoo62Oi4bZ40TAR9c4hPjWuO+6gnkzTtPh904+YLN8PTIGN6L5hvOqNG7u
2RQztvRGsMnufsXSQIAWWJMtl0I1Kj6PXK6oMa9b17xxFhI/o0GMAQu7qkI7
0zkGqfjb+r4/6KIx8XWPW7dvtEIApWamOwqSMNS3Lwkj1IFUs57gkFVBBj6/
uGgtyZMlcugAZpEy+dCb9BeWRt0joiUadfVEg6zpcyF0qhYNTuVDwFJwOjfV
32+fCJbFtfOnB/syiNHQDfqZaIc2PV+Nh6jxrmlBLAR2OT12hxH/X5QmiSre
1gy8WSne1vmzCE74A/3q3O8YfuHfpCMnjWwOqy5Qu2v/DUouryZ05lKv/cd7
0UGOzfvAWrUoui+6jQqZijmnzXK3l1eZK7Xhsm577dpq06NiNb+KicESU3Vw
s+gclZjmJfKfjrswqKhngxv3u202kz7iW0ztv6wBlbEmJiUA5BWlBTTgLUCj
FnDZ2um0gXWsX4t9l3e5x90jfXZ8p8pwIFC11Ow+8PqFnTdkL4XPvCTnAC/g
FvNxb7oYb94vB/BXex331mIyzNe1QWmTr1d7ETYLnuyLC3Q6qB2jDcfrbB99
tv/XErdmpwOBa27V+KAQ3EYBEPDXa4OmyAqylICaTtfEdE4YnL8tyzfcUr2J
NGK4UAQonePmGr0zSBb93a4+l9qLTGZ/BLMGE13s9LwTFyhA8IaXknYsCe0a
Azxqb2umTdQC0pCaj9k3kK4tICm0gwYeSQ5B+3EqSxYggDhmk74H4l5FDkRm
mGrPf7qJpvdv8ZVC925S1LyAUbYisjtJz62KUEzBCgie2oA+5pS0wAWlhpjW
2DFf1rDYWWtPG6WQnpoOoddmJs6ubAOG4f4fvIAAAysnAJXoeujr52eJ9g4l
Py9I7XRFPOCfjSd0st+tYwnNmppkpvT7Ob0pq2gNixZVeXBVuKWez93qE02M
CVMT5sbmygBG3/eJevESvKbNJp0XBuuufdeRRxu6xesErmnJOouX5j/njM41
WBJQlsvvfIeIpoaqeKm6WlEjfxuPaBQt6koelHG8r9J7pvJR8quFNdgWVIuK
SWOvrE0ZgNyY6jLB7JyoNSbnKYRUmuQ8iEg5VKxrKWCMP7smhndMm/J4kUGt
X/OjpKs1vc5OwW+5JENKNy1hdX1BRuGWkxMFYBFtSewg9++VB8vk+ZNaK3Vx
BsobC+5k+cfmIJg9pbrmjqikHpZNIBOFisLszAaOhooqJtopOpEg0FjMOOSK
RAvIDtSqnEIaXwgstVlsEoAngQqCjzDKViodR1phccaShCxVvR92pCPBFkzs
jibXy1pmJAkp9xcLYBPF5eA5dJPx9CUr3DJaQyGpOpx6KmUdd2gKqbeXMqIE
r6xpxfMxTt1eTuggdHz5zWYnHLKODCHrxaJRxdXLT6wPg9ayubh8Qb1N6U2e
HbnbaSNXqbqyycXfUKk6+GPBWsz+heCziiJG6q/Ozr6zPA7sKUDxVn1JbZSQ
EEmDdDtuDH89r/cgrwygtg9D1k7fqJqHetBDMwzu4MImVEoT0xWUtYZHEGK6
BZ/5QGjCJyk135fnnAwY9DTrsaT80jbc28rXGfunm+6RcGWxdDzJVQL3ucVF
a3j2tIkHlT9Yj1S/vhmVaeY60oDUhbu/U7Zr+TVIi+yimcMP8ZoQTeiwjj2c
/jzqNx/B1XrJhOe/pwzsZuvi+yTS8/HDtWRf8VycIRPOy8OHRNjqeHCWC+iq
RErVfs/VIWCvARWd5M1SIx9BiQ2/0CSDjCDRlNeH97WTm5XpLfZlZVDVwowP
7MzGIdGAimRTylmBY2gG9RyBcVwJan09nLoFOJbyxkHALlWCKkzljzl2kw24
QspwOD2zQpR5S4VJ+uKWave6MagEerQZiNwU3RYY1Qu57aefFGQ2a4Bd2NAT
GS5FzdlCVXn31ygyfil9uNYqKjrAItg9EuPJofpLRRjDO7h5mLqfZjKQW+ZT
nLmM3VmsE3pDve/JwlhPOBJvmZJ2YKL/gjMYsAo0Bjaz1RpgS0T81j8tdQp+
ghKhNiBVAfEEv9ZsJ6Q/4R7EV82zlwcNfghDm6Dcb7tmRr+5yuotUqq/mXv6
2IJMe59TAX9z0EWJl4vqkRJbQzDMAo71cCB31dfMYs835ZLarrbUELDmVltJ
Ywhq3d5eSbaNnR1C6c3Dqr5EsOrhPc/4w6NpCTt5yCFlZJA72cpvrJ1clmUX
SGpQYPNbhTF3Xlpt5344iCbzbtBcgTqYhhNBCDSsA6vFZDCWfXxuRLIrrB+w
aATVYRkarpOe4QN16ZeOd/Y3/hY5+wkcbjges8Heerw3UmEZjE31Flj2Zwlo
CEkzSurkVzjLWBm4/mmO6T3ZnX1Wkn8yZpr7czGPd2rLQIR0G9bENYJp2lS8
IE3DgiHKOuE8jfHpctbPohSNldFZmy+rLlNmfy8e+3hkLQ+LfsX3p8khrjcs
kuITGToq72VhpiByTIsalSgyZCOi3xY41Gh2y7S5irUu0gFM0J0CAdR+AIQz
PCsi+ARvkpYlfa1Ftg5AK80B9mZehZAgCGGqygHhP+7R1nHI+irRVLc2kUV3
igJnX24SxFzpi02kT/1UWu6LExLY3JCIVQTaWz65ET2o24d2AL1NtJnjN3i3
yglJcwUUBffS/yg383whSMP6m3PYiXWMkB4DMWAgsY9JG8DZBEn5O2tdtiC5
ljqNffOBqGYz/npD6e3+dtNwOpBnFZY0emP+nMv0mxOpjxCY4go5yImg/Cos
L87HteLEPC7pmvn6wzQC5mCBPTCbt+QGkxIVpby3nqx6C8yb0IZkEANQOyzA
rvHDTBc5BF3+UPOb7De7GSbXbXt6mJyiilHDy6IyFR7vORz4+RZjobTktKwU
BNKkFxZrrs05KvYNVXqmuB79ZVbdbLdqnc7U9m5Abmi4HRVP98smDubqJaV9
0TXze3Rh1sLhFea67n4AyWlfCpj5v2uumDSrMEDKjq5OccUDTZXSSM5e9TOu
SVVfATNhaCf5+26NyQq/JQfAiCcKibPXK+nm4Uj10oQSaQvIWdl9CYaCAYrt
oFw34eufEMPP3AISownjb8kW/McbVTzsXEvuuknr1ms0qn1XB9VU91FhKUTS
3Rk5AWzuRrdJ7I0YY5NmPRBPnU2tTRs0ggpmgbUh+hCSwWy73V/pAW8YnkSV
1tVFWNBhjIQMmknoj/iIFBUHksO1qVtK4kxduoEysYz1lZ4as7+t+YbbzXBG
l/90ArJrmqgQGHtNs9gGCTuEyjQHIEM2T0h4hbCMOfxG2efhX4zcoR0GdQbQ
Ao2Y0N6Qi95bG1KaRyNEislUF6bWBWpLFkYXZeiHCeA1+KHaXJi69NXYF4xn
7XGn41WYnhBgi04odsF86hRqs5eIKdiS4gxVmhEIjDSUzd5dufj3comPe3YP
iaayuEdVN8eCc9Nay0cXlzl9qU47GZVtcX2d6vQqnYpZ0o7KboBAjhJVaAOy
k4lg/MDKkxtkdYOuQ9mJALixkokzMfsX47e+13kNqDT+QyX1JjdZCludgbeq
ZAUd0OOnjbnKcWMsuptD5qIRqW30EV96/fuvfeYO3SZUq7ClpUrOwhw1dX09
mFpNj4aNMIk7gN+3sheGWBjtCsUwUptOuZmBysAK2sV1r18Rdl90Mn8WxPE9
T+/77jd13kj/ZA6N8BHcRTgOBLaDuWn8OKvy+GsnKvlD0JDmdBv2/FvEeYw/
Qt/wR62qdn7XhP/d58XBAVWhYS/V0Pe7gqIuKmrewf7tB3Hy3iWtHNNVQ7bO
eBG8h6hiZ1eiWBy5hrOYgISC2kd030YhN9gJHG3UOagFtFhmYmjYe8tXUyB9
cLhVBFcD1sGDXtYQ4OGC03R5hTZuxAWeNY3Qhft0CIhDaCcb/HLXqtZYoduV
e3C4xDJWVycb08j0hfW4CbTMpIyGHpQRhd7kka5nhmhsAoZdbZPiyl2BWAHV
tJnmR1RZsLCUC0hCo8ms4ysLbA+nzeoV6yaUclZxflYndQVRWED6wtt3JaAf
oet4jJaFcVQRqto1hpKHH1+SRgcTHaQ7RW5nQMa2srV8a8LVd42kF6QfJrK5
Zs2YR54c0OIhXgxU17KOOswraYe77REPm7DsxRXcFUR1yLwAgr6fVkSCrwzT
No2biykIpYpGO+y1crJU+7RehZE+VWzOeurtmlphtA83iiRI7Q60lj/0uvKE
q/kVXrqe/ZIAj56DcCZ6YQIBOreLlv9Z4UN+k555Wcg8ml6XeVrL0D3cTc5s
hEnklxhK6I4tvmO+/eR7UXyz0+5oWyBGcAztaOK3rrzglQS4uk0qz2B8PaRO
0Ul0Xm0XNuspWBdbhfYM5clXGiZT+r9umWeZHwumbWvNwV5rMYpWcDU0K/8s
JqFdok2OTFSDjw7nlyVCOklQ/8I9h17wuSA6W7OVQf0ZUz4MAkySAvXm2SdT
yy1uxfS0Vf/zWy7b7/kFH4W5vFN8aaBYoU0TeRVCy3tEDVMP+PwLaGI1r5za
xXydhLIauz7O6/D0XpCx7d+US9KwJXVOWfWn+8Z19JEBPwJP3IpZ+BW8rCot
Jh8ktst296JoqLFyP5/FQRXkxHP4lq+D+9XhOLvDDtp/2bBN8xVRT56TYUtZ
ladWCr6J0bqNETuidtfBv6cwP33IlzzI0MLYopT6hc3nmbbI71sN/W1cPmYR
jQ/vk5KAoGKAkpx9/1O3GTL8RGFOfHhOsmWW/6MrB63ewOgVmzr9blB4BJny
CxCs7WRIVTfLVwi+fXvHu9wUh2k9kFls5ke0FXfb0mpgdh5XXPKNI6Ol/lSG
wlMAsjEVoxyojlgm4TxkuqjblPUtG689klujZEFCgeel2Erajqzm4/p1hCkG
puJuQCW7bBOQZwTzKdvbelPrXTHPQi2JccZIkwt39EbqhJjgBOc9LfQlQRgZ
GNtsiW0Z4JF2olaSZvOgXKtu33usCZktYF23NH8hoJZ8aJVk4MiAKN3dG+It
2WmcGf4pRiNCAzUlBIYELgQuEV7gt9HfwJqlP49+5TW6uUrum5DjjoGR/90z
DMAuyyQZUPSI6mtsmam101MRvzCL16LMPl5NPTf13f/C3GDeM13hpofp0itD
WBWpu2aCYKQ+B9mbJwVVB7tN4b4tcpB4u5DXMgTMUpVRTfGUSVxeRN73phrj
iRDiqGfJDpiD2YUkrcWPvEw/QXsUrzyo/DaIUxW8k/dPbtAQoxoqcES8pZRA
z9thBahXfyXMKgaKwJ3sQQkQUcXpUkglKZw18P8SoAiNDemxlHpz3kPbrmmA
Z7YHGXbgbok5Z0XQyy3aeNj4qifC9AAO6CvJOPaoigKDt2y0DkRZl+Kw+eYm
01WzW55vKtQIuN0GtV2F+xx874qYBF1OJAMet2xgTMJBOJ2Lkx2GubyRktiq
aZdEbiNssThiYsSfyW9uMm08Ju79yqMca8CFdx5wi9pJt2pV/QSGYmNOCqJk
hXnwh5sNQkueBo7mm28jlQWaSfVeKOwBAu8bPLFFg1HzXAnOBF00T5IzJmbD
33Zn5+Ulwrmw7p/tZxWA17/r6ad1CTcGQEQphHKWfa8TOsx7Q8O9aLq66L01
k3kGMEUzV4+kL3C20wgkFQfBr6pTYKQSvp5JkDXEz0VMt7PodOkYcQmbakYl
maJY+EBEYxMzK+uOV9P5hddLS7eN2tg/NY7nQI5ESZgDiUZZz2XPra4bUk40
Mr4l6KXXTWqkL8fMyQGsTt+lHm4eV1to2qh/lXse+jOo+FngA6e8YkiFDZy2
UB5we7OrgHRb4el7jEQZvguRPSDVwW+rwOf5yWB7zs4csEgknHAznrXGM6t7
6S/ucuwQymgiYRwm+THCgfSRlcrK0rB2KJ0So7Lf7E93sdL8KZAfv3d2UXFr
hRZ0tUnDKJe7j7UNt4CB+HhaED/GIfJyar1c/u+2zN20864iuzcMXHeGP3NX
pwo+YxQaALBQ+HEpUX9MpZnyxpY/OmEQUUU9H+xbBGdICPMOJE3E7lQ4JWhm
cGT93cP6MIM5ekLqML8jaYckS7t/MWBClfwx/UHon8w77V7yrPTduMje9it0
LAfN+cdqU3aCbvcztRf3ZOGfD2N+TPrhnaBJxOjknhHBvUccTW8l4OYccFBE
LQEEac/hwAXK+iu6XmDDsSq68lVOzpWZy5m+qLKlLYEfR+x2/K00T2s//I4m
knCUul70SjVqZcBsanceBsfrzU6YM8E3v60aiC3cgSGStFSNQaujlurwY+iB
HQkV5xlITwdbESO6zre3S10DzBJGOJ/0LFSPK186X9kyV2ye2ZeIEuSDYxKN
jlgiTWSogpXmyLsvj3GJIvDawQB1zoecOkfsaYyIaw7H98TKKekda9CsXbdN
ed7uEA0Va7j2NnSy3+rOSpKKQvqeiT93zUNFJ67b0qWmdslEmRPmoVB9ScKk
lWKu0eqrKOaRqyB+bNK5itypKkESLa8jUB+caGuyFeLzUl7SRffXQx2T7jY+
RuDF/wrnNR+599c54ZkieIHkz7vWNP2tE5NDHEb67Yca1QeWQ2OFHbjU+uhI
xkUjXjS1oVEF4pyD947kTbXuyCUgQYFyUsorJAX4qvOIoRvgMU6JApRbb03t
KSSVhqUlao3/0zpkZzO4LuklODV8SUQgDGOaNASSLsw+MIN5ylsUiBiPcVK1
xqBRmoV8VTiclQHmrfduWE4B/wLOpZufOb07Z0h1cwD7tkeDJ4DHkq5yMbU+
AwTMFwVQ3v9IvRAjRr6NSgxmEhulCFwPebBrMW6HI4lbfLZJvK9GSGvUFQ1R
/hQqdW4XNXVIT+W/Py3a5LAcDTIWWDvUFicWZs6cKTsUPoGawzjMf9eauHHU
vPpFXudOR3MSJk3hScfBMlpqzFBpu+I+R/kspBJhE+RY+FigZp9slhiPMxNi
Hf68Tdk7bh065ZyyMaHMMEmaWKuK6A3v4vvnWn/jEq2oJXcy6+yIX4IwdBJJ
z00nAIQFUEYu6PGYrKnorZhPGLDtth5gdNFa3zd88adJGg30zO4Mt2UZ01qQ
TufF7NtgAkppL5VIhovdrDtBebLJ3EP+MzKj8+Hqy9klwcPXJpvTYatqlf1Z
U2GDvDkU4wn9kHH9LW+zQ1hInC5jcO8aGarD0Iz/gDwVSbyRuDjYH1YUDB5M
dUU+z+k+X+ZsEB1qNgyx1XZQAn2LNIlhCHeAcuVv/x6pxiN/7FLt7Ipt6kRp
X3w/2+dOtL0xttEuwEISueffOxauFgX3cwbcS94YJLIaHvAwSzdYTYC0I+Z+
4lZ8sm97lfRByV52cKch5IDeEJWhX/SWozXeg2zCGtTJFpY/fW7TD3/sa2hp
bUj9Z3iGB7iGsMR1VTeIcS8Qjw1YnwjS5f8/fi4K/UHAStdmsm66QhNRdzeH
naHcKW5qxO0DZLA5Mt29BrJnpJLBTAJpjLmky5PsiNQWPE89jgiizIokWDJs
e0ZKYFEg3MdW1K+0CxG+Ctb5h0hfkUFCEVniJLh5wDyGYVQ6LXJjvV4Oz/EP
KpycKRAuMJXZHhN7xw6jVpFxz/HN21JSBS07P4K2tXwHDMhK9DYVOJc5tdfN
yT7CAYw0GRA5ZLWFr5qDprarwBvCftzvGnUfxn5HkpAF0bJN/eAng+VxmEdf
PTqM4FwvvZvFOXTTzzv8zZUfKJ7rSHyC2bMiOFPsxypBiEDsl9qcVjYTurJO
8iZQirLURwTIKjQdb08lrA8vGM6SXOxFWuNXJS+rnSdeIkMiIyGCOtuHOVdV
6i8WwwddLde9RDYIxDIjFXlzXko0BtmwczyjF4rF9MOGrasLsbyrE+PhfCYd
VtR35YMWERHYeDnNbqqELXf2OKOfScq1VnCx/L0HtPwq/OMTLfe+dd78kGoU
RjjrSTzw8Uh8d1xBgGrFN6ncYlF6nlJBpbvREP2cKZbfTDqgnStc25GcdPcl
UfKAtVi2n28LIYW+RxYp4wJ6gxg07a6ViJTCQnltvjQ9luIBYvER+8HLTE1C
8vDQZU3dcNugLdF1wVe8d0AlqUTju1iv/vAv4qMDelV3lHlk7LvDm4vb4eW5
YCou+jRCshfe8uVf8r6rxECSlh6IzQyUnh+oU/JzCF3jESe1FMsqFetT6Qqz
2+8uG/AazSDLnPuiC2cHXbkvKZbY3aKmtwnzNpM/RWg6fnDKO6r7wZpZShoL
D5/K75PHX3QBKaH+vAsOYlJyb7MCBM0ET0Hc1Q3yfQ5LSV5PTRm+pPdGufrb
xnrAUs8tslSHsxoFrI6SkA2PfZ1xqOuriYIS4WLN0l7TgwAB0pmrxk8qxpOR
xfpAlthMq9uy9lCjJxAAGJ28xbIITLAEWgWeNuknp+HBDlouca2q1CRYqJ7a
Ln+Kpk8LVriHEV3hlblKWKCfwShij04V3W6Ne1xY/C6IWP2T18pE0ckG7S2u
Jy/Hc60CK31m3yBiua3fP7F1Fw0eTmU7YIBA4A6vBacwJgTQbS9aGovOSJ8x
dPcP3vceq/BeavJNLFvD0ukWDVKzfgayk3CYvoDNJvnx5zfg/2qVEYQ6n5hP
JL/oIpNw6z5wDB6Go8OYXhpqxWkG7k/k3gd4ZdYof5hWB2R4dgRJh2iiGio3
iJtO85d3f578C+NUTTfY5XCzX0aZ7kKH8AemI2iBh4wXPIoBUgEWZBXPKbtF
TiB0kj0AsTTRsjx0qR/cq8zFKWg16teKdsYhiSA2SAY6k93bCM9Bfzx/eg2V
5eYHxkc+Jiuwfj0IyTeKWtd22pE9XLRHvVB6753H2NWx0xusRH5lMtIk9YIk
fpv8j2scQVEi0SkHI1N28UQ+P51UMPP5XghBCLqU70py4s4nNCtdVVYNA5V8
KI2q+AdvCbI+flc0YVEMHRAplhsVipVzGZJywPmUuMcKBAiCkhBFClBPDFCv
heHBlu8DiELk1aBtgQUb/FcdLBEP0bX6sHymC/wBgelXGzi/xsDUBmuKgq03
vMlNZhLJb9v+ltFe+mfWC4kMEbVW/6r2U6RuiMCMnBMDm+/DvScFt94w5Ypk
nF/EkI4WTZOJ38zEl4hMDizBuzq5DGNLAHn/u3S/Yo9/A6c6I4WuMDIpHkez
x2ARgU/BIj7ItPKZeVx0z+iGzVoLiyrUbNLMyZTzDTqJ8ip6paQ72jwUo/QR
QmllVIQHyBW8NGWk6Z8zP6fyidFrIHnrPJZkUCLbMfa2FfYkU8Hfoi+qY+Lt
LRE6YdqI2PHzKZRY7mjl7WZvVkCwveow/X7aEQnV4NIYcsHLj63Np2CqWKAM
3jv2XHz9jaXl8lPISriH5Uy/krzGkdLrfiUmfOHioOjzqADHGPQza0W+aGUt
qIYZ9XgDZM1OBFDMunL6ZlmCCTYjnIqU2WXnYvj8/4Qy2gJBsuBAKTV4vXcT
VNdQWHDwpJywuXhylyHod0qf+pRJ+5eCmfTq/2lQguOtVpYXdHnJzpNT70oN
ay+txzVMPtAMkZBJLjTBTukZRxcPLtkRgWMNTl/mKa2XuFSvO7HZ1V0QDg7s
lHh3nUL9ndkV/Gi2PdqzcecBGOdqGVxxDB7VncgH1+ROBs4DGw3dutjVjQf9
l95aZ8xMrBJjgtMJdBNfSSNlNuWhRYC7fu2Ad2zNSK0SXkUKpvEtJaSFbhAt
kVr99kc8jtYbxFh3jJ5LZRSqGjsFFSzdvWqSxqx8vjMcu4Y95ukYET72m1bF
uEcB6yV8BPaLh7zbzkA4zPFAFMYxahY1GntGc9ifl8+y4rjnO4prVdv047ZG
iK2CH7mLa0artV/mtQ0CPEggxKMg3AvGafwwW9tOYwLEA6OOU7dBJhZAWKiv
lU1ur4oFMi3d6+KiNyV0hUCBw/b9n7mizTf/6j7vtKzLnsNhY16DaIQf/SZq
TIrwd3FUet9BtewtqS+QIiC9mmjJM5ivsBMiCrdegtXRd/Lq6wE2maBuTSqV
0I68MwfGzr6L4j2T29k4fyzZZhVGx3+7KrixYH1Q3TwqnvE1cQsmS7J/lvEY
xl119dRUKlAtHTSGpgr1ZV7Qef3AiUmckRbqLMFV4S2WkKLDkm5lVPwPsp5d
thZR+ej7Ld7jkWeLktEJPehUX0+w+pMzCNJubyR6L7jq7mHhQsnzxTD6Lck3
Uem9UjsHTuru+ewyBRgULawWQrJcH7WYACrg4aBmpQoqtCpBSrOZ3dT1kyEq
cOULuy1nsznYgPZyM/PdO9DTTlXF6eogyIz9b93VPASPVcaj6paqyF5oo3mm
Y04Zw2KEolXJ8wMr+BDPDWsgwNcveUJ9ue2j0kbPx1Nri32fOfedIEh3BNRF
7hOAfwya8qodhNYGtlwc5vl6sl8P6zNRmBCCeb5WGwX4SGnUaFnJuRnJEPc/
C4PiuD94O3qQlZ3a1FaY4emWQqYeiP2ybx52Z8DKubBgRMa3sEa3u+WnFytV
JK5dvQ4sv1JIUmwW6y/XP6fODToSvDGf0uNcAFWsy39wpzJGo9Q1BnG9aHYu
hxdCTs3GfNqvvWDpF+Qxtlk7Qa+FVKIqKY2GV4HnOroMZBAe5VN/Hh2GX8lB
wTrsCHPTZWKRtARz8TWiJZApXFFKw0/CN/pYKGIrb+KvvawrMCH+XQhHAxjb
VcrTrGJkb6/lp763L0Dh+kl/qsVb5jNZycO/AkBkh08p5QdYJHjwhm2R5wMc
IAg3qo6X8sUPoVM/h4fK7t5rRhgPVJzZPMhEggtd0qWeSG4cMfUf0WNKtZWv
eYr2cv4WqkXkP6D1KuZ5J5wDvPlf0mE0wF5K94WeX6r+CmS7Gb7L4lGCYLqw
mOI/PDUYaestrrEX115SjokNdS9Ao6vWuwTYIlSY7HsPcFdgnu9FpLES1e7O
dDQCkRNefaQAxDxhuikR0PdkKQCHk+FDFEgdUDYtM6SN0p9UbdvZePri9tij
2b1CbWWtTZDLhgdmZNXzusVLBFaBjmPYup+FSu7ic9gGJxsCZOo87MIM1JLj
8NueBGJHmu1RDreLDjVBo7IBOY5oYHGQfjeHvIfG5JQmeRtCMgQr4DtALOjV
S7rF0JvjMl5/BLemsojgat1o4vLjgzj1UnO1HlA2DDOhiRhi32Ml3LDz7ua4
LsWtWNH0tUQUDH8KmxahM5rQ6cmQKSq5hEhCVyyBNrkzeNaD2lnVivAXUK61
X00RT/5d8RXwa76PcStNkXDxu2GRQABAkteng0FmvcediS891kxzQUNo486S
kvtRNKOequ/OwjP1RNA9ae0mpOZbShbwfwawvodR28X6+G0zBdLYuu8Qw2zD
/1iRhbJIMQQ4k05GW682gFVQLRijlADI5ur7lwNpVwWjcOs0lH0y990OiqnD
RyqTxcqXe/70i8Jy2a+ETBahYv7NcEHKuZoK2JSB+GXadQaPzfIzkAMe9FNP
QaTPYBVV9J+Izkbzsw/dcW1Cyp5UOdhjJWg7fxzykrGFHwQ6z0414yTVLDGk
rsSnsILDniOU/e5tHbxPHsAQPJ3pgqLNe1+Zm9rcbH+7qEW83hSKOaVrbfUI
8+W+ox6xZt2SA0IqY32Q6DViHGQbAIqqsd6RahMor1WF3b2FNB/WSQT0mANe
nGZf0pzlcra5559+jkRkr4/18H0S6LdeCnKKUfOfze/TJs/HTMAEjTEOLEHu
R6mh3uzdRjYddBKxb+spJ1187gXnKxkwOtmIreONrtoNopNRadW6PxVEfqGp
OevxI6b/H8YZTH8x8xT5UFbZqNKcjN0oAo9VrBnRp6PquD6PZaT1tvY+FxhM
P0m/KlYgIskgrNcqxI5Qlo5c9yAa9byewtZhD6d6aPoccNbjjFs0HjiTyHzP
G7YLLlC2H0M0riEO65HDbQSR0RLzfsqH5jXWJb3AhYwxbcM0DFUJXMPXm9UI
OC9vutU1RqRZzINuItRnWE89PZn0V371LKEsSAMQlz7fVAvWUEKXPmfoBDNA
seRIGS9CaFssA+jaBL8P3ytPZtFgneyj92DwtVotLYbkCN+BXWOtzxbEJ/NT
m6yG5VmCbEu1w0KeIinuoI2oRRwXReEq00cX8vGOWKqvoG7FSLZkjc9qRtXi
sa1PZ92JQ+km4vKq9/dgQ2eWfmMudDJh1B7czb/96XEfveszuJ/+gJf6Cgp0
zcEOvm44IDlTg21PL72/dohHa5t006Dj0tNJSfXRnh1Fqrat3+F+LYKmnLza
fP8FeCNhffruPFctcRNh6o46io7jVgI3yremtPmUK3aKfNZb5maW6SMOqzBq
DsJHedTTPNtUFtWWxyadfUrksS3Nae1Pa9Y4qAoXv+0OIkpnP2YfGGlbrsEj
yfMB/v+WgnVu6kbjIKX+1Bz6J2q2I/GXWbKpjNPezqrq5Obcx9t7SdwYU11A
q5t8b8dBU3sNrYsiLzeGJjnF9vDSy0sG2LjOR3LyEE2A5mOLbNgoL9Vubyf1
9rXoE2labezBdJJjktaWgphdecZmvfaUng5FDI2FUcnXHyuYQFy0jCduUd15
y2Jjb5XGNRE0RHPQLzvGgzheQ/LM6nHvPWWprQ4aMeAAB48VzSDrTMhzhTqw
nTIkD/QZOm7Ccwp6ORVr4Amo2RO11qJ9NI+K+k3LgvJDSn44r151hRMblB9c
Rdv4BxHs+egiloYBmf2jT7OGkeKOLLu299zr4KaPWEZQEHP8TzyFhlzUqCzA
u/yeEdzBkO0cU6vOKJ6nW49qf84whAn3eyHONVQFJcTD+vQwqKP2t+zWRYPf
7QhovilmxDMlKSzkQW+yc++7DCarYfsctkTbsAqMZ6nToSSU+mq7mrYVizKQ
esNx8IGjQtQ04N28ewpC6AlGh2KVBpHqQM8b6wnMFcI+V5yEeEk9qtMxLzpM
+vIdU8tUjM4JhPd3abSpUqPE8OfKSzwn/3vBYMEdDqzvT3podBVmklGZUwFs
J7KsDQ1id5QtFpG20e4MDrc2UjTtd2UZUHcs7iQ7PjRzebdh+LckrJ1B0039
fvlHG8HGMKA2jdLgrrHaG4v9VuQUZHm5wAJcbuHI+HmX+/2n2dLuDXWCwcF4
sQ3b0hupGJqZurKEcYq3J9/2McOEzroJPNTV8T9EZjnE7K06ghVRLXnxE41x
NPjI6mUMoNJxtjmgBMv8b+vc72KMTKyKn4VV/jFFo2ANqI3k58N1JnpP/YKf
Nx9RLCzk79WXu/jf4euXTtuDRTdpLgeEVLOFPiEY0Nvp4boaKv06WmqL0nB+
j2VbBU1l9L9C72Lwm+vjCfA5U4voUO4b+u+4mr5ovmhgeLHV2IztTrTieq8v
JwkbKjOdZejNXCzMAeeqca38rdG2HE3VHx13wmybHq1VHhi+ViE3yTdMVReI
8MYYJblQmnZWi00AQ3wr3BHUhHHqQmty0GP8GN8w6lCBTJnTQ/XG5xDqhxUy
xMXkD51BtYKUF/dUx9eAFuR1rkEAzQKfVcOei1yAkY15Lu/U/NLJ2bxCtB1O
/4cjWOHl4B0utH3Qayw67pTQ5Fprrq1r2GNaXCQKjRTIcuYGXsqZZJuwZSvE
8FeK/mpvqhcOMDXrPjARHO77+GrliZXT9Rtmh1puQmxQuWwUhowXb0ZU2+F9
fYSEZGKrp0tsmWTs/J6fTuYx2fkmWeFYM8xlY1EjiSgPGdiYx60wynGqwjhg
ZJnuI5RrhX1U8cWEJIGDO/MF2ZBtQhUw2+v/fGr+hjMiuTjwZFyve3JO5316
3hcY3zjdI4p9jrzazLgzIN/HbJqB5cPDkdIw2tPryGCmNA5V9DekoM7/KMkD
usQDv+SCGc94Ppe0IIRwbBnv462fXophRjBASv8EI3lEYGfy6IJw7gnMkbdZ
dGmgIbuXujeq+U5dp2n27hTV7BRib4BeGRqdQMe329Z/X2MBixLKakxyBPSK
VHgKz7wEo1sn0IGVCZNgX7TlXpmVhKteHJWtL2I2yxj0ltevuQACm2fAXvyT
hOiOSVPlZzn9mJ9Suy+fJiE8/hPi1YsNC/wmg9BHKSkXGz84hAZqDxLGMSBK
CzkD8fLjxeONYDMgabK2teNZhNVuTo7xoSeJQKF32Je6fmbAFhXs5GrNdDmO
/3886voKDLnkTJUbb0oZWAqz6YA3s5BM6N1oBsxkP73tgx9Ry5fewdJyxRT6
xduFwO3eR9VeRHeorkXNea9Q57UumEXxnjeCe51rqZPn2ewXACaQTxMXGMIN
l7PMHeafOHflRY0ZBG22tKyg4ytxYcpbD8hwlJNnw5dCjGFEYMzlByQC+UFw
MjZbiFghZJU9l3RRxFz8TVQcSqD+mve7RIRMYC4zfkOaBXTIfelU2IOaqjaM
KBFCg1ba0XHvUqtHPJnJvQXrmo8ie1Xh0DSamPkoG+Qi0QnbtzgehdWcgJon
Io4kCfOxKXZ30wdnru+VedOueXMIWPtJgsNP08a7pOgk9+oIxmMMiYNe3QmM
KTxCIekQnZAGywgsMx23d8igCuaNH987CGZ4BjmK/av0Y1e9TPIEzhQBBpWr
Q8Aep68doWw/QBLSRbdPYtHAKbc3OhDrQS5y1HDkrGwnhDd2u/8cjmF/CMks
II2ptuUFjJ8A45H3coVa7vdefXyk7loEBVDrXgRhXBffnJlzMC9EM7DBBZN9
ciLBuoJQIF97lRWUFN0CvVBHBuFcQlR1ctuRrp1rv+nfiQzkWLe8f2Ts2cD7
UmAQib5uJj7lSn+p0emWgsJF6hjOhZxvdiKH/d4hJfoyrAiQndljmN3tmuOZ
uKgaLnWAhMc1IZWhDZW1VsFQM4emmT4Xa3iX3iJx82CjYDNyjLq4f7eiim2V
vsBqR8xTXugt3zcaeaVtRus9Jio+jz43qtHvmSS2fWZYHKb9W8GGO4X9WBC+
2QU7kaR3fZ29vdhHe0e+mPxvozYzjmWYBc5/XZBNpfTSIXCoIhrISQEIkLyO
n9zTGlqKhMP0aPOr1X7c6r09puFtOfayoRJtpzn44VJjc3zs13hwG4k1i5w7
jSYsAn6Ip1YHI66Jovbeg+5C5l4KKyVQ3G12JXw9au1U9uHwH5OIAoMV8qaw
JLqAkxtSA0ZC8EWABKocDRKbTAR80t4RUfzPPek1LSyARVbw/5IQo4VmcJpb
XCRIljjph7XEkNFjaS90fywmcXEttJ4B7/oZ1AeKdfKyiNx9Mum6I6Vngo0l
tXylwiUH0uXGyo019nknroA56xRYyLQJW5p6rY6Q2YBYKBi9HS7xbFsAJ6Ge
Opky/OiPWCkx8DGXa67h9EqUu0p8JoYlN3s1l5If9YXpoPdjMyI2LyJFWmjZ
7ItLnTrMAwvz1GXK3mSdLWWr4qdpAzLxZQj9DG43DgjtME/iCoN7JlBbcLNa
tsGngaAlIr1lzjbHsGXl4lqUJemm4fsWQQ78LvhLXf6LDdb2/ufDw6Spx/T5
/g+dnFe4wY0Qa8DStxSM9jIacLZR4DqRZGr7ErhAIdNO92LERBEzwX0Q20xk
fQyy4IdSaZKLH/bLeRBug4B68wWfTZQ+a3a2ubfWiQKa+4/lec6jtwoe5rX2
ejtorcx+PL580iWIFJVIYCHU++SZGJLcuDZc8e9cncenp/w7AaV8udeVs8GK
XaE0VC9u9uQ/vOJuU1sTNXyAmgWlSxsY57xkrJMlcgL4MJSks8sCguBP+giI
cCbCjwMwQ94i0KSCW8mVb804Vh7A0d8BA8uN9ZB/wVZChFTa/dSQFPw5GtNa
lQzr19MIqgWVwYdBy2kEECthFM2Ozmbj2KG0X0LWSaub/+2vbNWesAv1DEos
FUim/TaH5UzqYykfRuA9QAkNR7PZix+LMRIMo3WrWoDacikLaNbdzD8XEmXX
QfuB4Gx0Y3zh1vcvNX/oRvPRL3rR1aDpaHT/5CJFSnYZymSdyF4P3NwMFSNk
uP4KjzsAHcAK73bBQtnXvukVXDDYVd3xuBf5AZJgWyEthoOeeSpCxSKuv6eP
5dcYttADgfp5O6BXvj12Eifise9+fUVjaOh9sVyyBxktnJ4c3lc9Gi5/+wSo
B76rEj6SKJiG4Zmq/pZbwlVYtSMZNxKCNJTzglBIPaGxFf6QR2sp3r/SiitX
JDdS7fwpMqtutrLKOLyfPglm9PG16Wdr7gjd3mvVG13ZhRW6qpsYnxK4Ohgj
LW5sU87MaZiHtIG10kwAml8NbZ3oCs3UFAtthsNTcNOzMTZ922lVC36xYFDZ
n5Eqv7KibGpFDQ1nosc3DtvY6XZk9iuJ6Aj5RxEKSo/blZsDkGJXR96sqmss
WGxhTOdT8S5QD2vsODTB4WxK7bbBu4jTl1kKw47acQfZCdzQlqfTNcNlkK/i
oOQY6/6vhzC7jWZtDkP4w57VNdHmgVJqr515JKTGqRZrFBUPFyJHlcydWYEm
aq3PlR0KS/uEmhQSXjJ4YIQjXfTQoh14O6V3IwuyeskQDsxsll+PChdg4SrQ
oFgkAtikwSs1zBjXMMgpkXVQhL3GXNdo1mn/Hy0y+7z/CzacCQWKiIOPj/ky
TCk60F1gnLp4uBaYTPE+rLPtNhFnkK6RFOdOMxsAlJnNl1FCt55eCAP8+PWK
W5xtgyKhQVXqKma687cTWZrs0aS0Dy+4FCP0nByRq4oSjoD82V8TCvpRjTrA
2iPRLCyqxL5nZIPI7QF9jMFrM4x9JDKmq1XdIZh2X3Y2lkRKPkLyRbtFqU+n
iYCD9YU5GVRfbkEPGJfU2eL26D3Wu67dJebNXJsMv+d3eKHISz5XeaTVRLvg
I273ywqgZ9huVdnclKKgqQXhfTKQpcYfGk9z/UwPosaHppsxt+VS9kOTsIsY
vPEZdRgdcXvtkmnaJQSdWygBwUzat1W8gavuIIPEptIHXggbVoDAzaoEiNCV
8ibrLTy5ljzf+6XL7VFImVoFOWw17MWz/88nhfoJoodU2Zi2ItjCyBrErysV
M2lJ7MZolH0gFJ6G1zE5ciL422Gi4tLW7tlXmO3VgAtLS47vErGrtfKBXVHB
mv1Shihk5I/1El0rsl6VBPFCDoA9MkkjHhw0Ycr9XYGg1apXZypYSXVySg5b
SI2RoTga3DbbLPJjslr4LbboPSqOdfv8x8QTVtxVZMklrF8Mm291U2H2czGl
+6kpmIfPpQTHX5wXA40E0pFtRCDNJD7MQVqd3n/MzxRaySTLUHorNFapJGOU
1Pq9QkFJD0uCPSRmMuf3up/+8rIUtnTZTPFJ7EYBgl5Xw8MFzPkOgVn1oXi0
lHXQLWS5rj1uyO+TNVcubiTLjf/6nBecWE5R7ZZCTIhuR3WBSIyFUOg9bdKB
M8Pp31nGgpFRA+6YrIKYt2kTGY3OxSXXAYpLH/vHIGaPZcribYMDqBuorcNM
nz9xqmgPxIYz0hjhrFwTjE7cmSrV6I6pmQU6dOxK0PI3X9jgDWYSVKUJOfsS
QKbDrj/KMqMMEI0B64s6G5unKwFNeBTkawdgtbi7nht6AC/jmcexYgjyzUe4
HV9Zap6xVAGBEYrtdvDEGvKMjxneuwDPwkMIwU4MuBQxKs3y81TIbwbLqLjd
h6K4O2VUUOyw8VQvv2fY3eZ0Fx/eGy7bCnfRVdo2DBssNpbQpbbZo+o5QaZl
8+aoNQv9xbzdScTB4OVECbkiqB2mLN0lXGRnrjukuGYCgrPwbhSzOG6XlqsA
NqFZtW5I+ZvUy1/0+OZRfqp2zHeovHA9G13IchJqPjwhyoHLDwSwbeWTc8k/
i0VBy8gVKCchl7QaBkZPovJws293+Mit4TdCh0RNOBKQmb76Du6l+s/HihQf
zCKxalHZxVwlJtwZOwQNu1S9Bt23Fmx4+jRZ4eD7YrSTCrIDzN9y720p0vbE
4MdybnP6bD9IrnNyJ0MoCDNITn8nlXOIBLclMY90dqunLibbOfTap3skbuF3
wjph42qx4z8oFbNFAyONyn3MZfSqE1YzDKnIbdULkEU0UUztEtr62JfupSdG
D097/PWhm/m1W42BmLLjxj1N9ECNtA51NKUHIt9EDdiI5YyntSm9tl1ZSAuq
36EyaQXwLGQplVn2+uYnFQT76Qg8gnCnRqnTdW8buYJcM/i/kqtBELoFf0s+
f0QaR7ZBVXhltyx2IApfYZ11kgw7ewWUe5TkUp3BdDkOAaSDROGJH1PPB2eB
9GC3f2qSdSv+vvd444yS8fjly/gTbMVNjB67ZpDV48wyMHCcXDLWVFfB2uJj
sXr7UjlV0B/6Oh2KATythjU335m30qG3JbFN1jWLeg+lObVahoUi1RhRl1Am
sdP7yanCYTXbDdXnurmT4g6kANPMQtU/0RqaZ5tKvdvJWan0CjvvbuQJrKCC
JgScf8mvX5mynZ44us0mZSyD9T7lLG4zyV/k0pqg8BLbZrZH3hvsGIud4BDx
OdQhPlMaMAc4qRuQBTiNA2dLmQWbht5PvineRNVtv36hBZRJ8tZ9uoUL/c23
UHD5m76qQS5P1cXfJ2NP9OBJcTn+lr8f+kDcm9Z3B91ma5NMky76ZmLy9pCj
o1wBfq8lcfSY6ZcgsGz3mtPrADHyL24lJitSw6idNlRPw0z9V+jZr94e8wDl
GN9GLbEA6Lk2g2q1P91OFotmZ/E0Jb8JzPz2s3mFdgXeiNdFTx2hpTXjxkhI
4Wygxxz0i8gvboLKeRkihOPfLviAlgm3q1K0EOZnjGON03x0YaPCKYtyFHgy
wmFy48fOaauN0waRUqX2DTFnCq3TzhqkFHIXKpI1JdzxVcLDh1OJ+/tQ5Lvi
MTprZAOPM07Vf/+1LCXD8/LCUSiFGoy54jzsp/at4rvIpIwpm7D13o1Dkn6Q
MxfoSb3w9JJe2zmSl0GtXLKYxvvc1gLk/FEMHlgPN7OYRjoISAX+DX7AMvAJ
Y8bdc1o358lECHEYnyxKJH7Pel+apEsKKOKx4D5TPsLzqJfIALnR3D7c5dn/
1hqHUf/RdNAbStN6F8ULGnpTHmMEAN2WCXo6HB1owsYdCv0jQsu9AJpFRGI4
QW4CyL6Lq1mAmpoqfcVl7GUmxTGTLTouhCtjkume0A2CberzkYw1WMyVnraP
R06CftaUq+vTQwkQWWvfTYKK0qokYAhvQKJYuMOfi/orH0UT5y0NXGXUmGlo
suvs34wyGYw+S6hhVtDLqFMFezcQVBqcHums4CfpKwNE8M2OHylLG5sa8L3+
QIBV7WlcrsfCAio9GZKLowptG3EOUSSlCqErhBIIKVw0DvEk+b8t5vrtyEyh
3nRWHa6r2Xpv0tXiIlT7ZsXYdE4g8gjxdlUorbCS/+X0weo9aFlWyGjhmTA2
pn4JJgGzPt2vJ59Nxwz799VzM4ckF0qqdYIbUkP4SfYMKSeH22HeNrtz9BGb
2jESBSx34El1H/V1aAkgc9D00k9m796vURboyrzz8lzbKCHTJy3sxzd7ao9W
RClXXId2xXf6N3tR1ZYcGx1fP3YaL4IMv5P/hOb8xOUfuLlUGN04Y9PAIyuv
/lduWaqBH7qe0I9C9k0i0dcULkktg8UQoI8BYsjij2AklbrA8U45VGZDkgAV
dlzOR2GVk5l5E6o50+GJ6aUBuz9v89NIWGXKHhHX1k9I6mv/D7dyZK3Nr1P0
5PkaqzR30RoF8lTKU6gDcWfLH0HT2dUmCUPPCLZZ8SdlG64fqokvildhOBXw
q/mKe1FGKBoXzmbgWrr0jTU2xWz7cHHfJLMg9hwN2251BFTP1O3yPNLdSwyx
G1wfVVp/SVq1kzv9TBqPmj+FdqqMP0Z7zKQHNAvxg4VFCLNBK3i2UJ3zcQ8m
BwOego0acuyMgbeStQ/uR0t9bnrSEuict4Gv3rRjrTKddPwB1bvIpBsQ7fFM
XOWT0mAeGB3oQICQRv4ZBj48PI2mxwi+tkaa9cho22xGdwiRyTzi64XzJVh1
ZMWG0kTAp1q6l4+XOHMaBPnCVAyzAI6fVv1/Ok4xil8yWGoOsNYx09Yh5wmW
tiZbzYnK6WOctPqKmcuuVsUZ+HIxERbaU7u1SXacg80O5dGp30+SresPJvJQ
EUm0RNkX3dpuwcSzf9KlLvK/xBurrSFTuY4SPMiERJWoM7kJoDfBL4fR6i3w
aJg7R/B7CSW1L7tCUuf4vhEtDpy2mzA4AHJOxIXRqhqPRWaS1YGlqfvhaaDE
jCeU2ONp7m1UZuHxRlCTwtKkREgjSaxDlOc3RN/6+26KsXgAWa7W0rtec9oF
JO0uVX7LAFWhUVjrMw5ZweeI3EM1jp4hpwPfbVW4dfNF74T1bXSfB1Z3MJh8
j0uNKu9cxuSXh9BYfrRlHv66r/xyXsi8CQk3URix3RWIDsY+ou2xfedn7eP3
VLbxbt9CF3q9QbtgR+kLD4xuFdMkEEVSmAxI6/JegaInb6/8Qzu/p+d20jgN
E2OxQ3qtDAGsgxyGhrXQrgTE3r5Wh+LHUqkcvdusTqJT67Wl9JNIKD7IEvPw
6RXN1NNrN6gvS2fYtRK8C6tFPC4kgsjwmNV6d2If4zbWkWZWXkrcKgUE1nlH
CWU/h+X24GYiSijWaTOit0p2RLnEIdnGpzp/17Cys+WFkY4TkHr/z2Y71wGv
HHWHazjsTkLRtlmljB9OxTen5ds9mr3xxOMtNBSh6JAIkxxlKUMol2P4WLDI
7vTbUak1ic1P4ZPjkS8XewWiEmmfDAIGy/bX1J7T7hh6r0CgKLLZq/644apF
syv7cnMuQ1i4wGlyQTEOGkC2u2RyjNQPRp1cT+HFjHtDPpkJFkrVpBjZOYks
dAayVgPW0Q7Gn40eADrZEDgHyrRv5aQ6OHyPDZ+IETMeDvXQ4cvpDLxcS+Tt
Vt55LiA8gfuYrM3aV0zkwaanhYk//rawG7RJcwXWAVV4aWCAP6/6jMDbtel+
p3AbqwV+pFKg8VPIFMk9hRGNlPP8VPn9HmuVXZLQn553wc5m1GZ15E0OFvTh
s6a5DAtBGrwtwEX0Xv0EkfWS2GyGruwU5t/L88WwDH4oKOKbDAuiDhzlFDdB
GsuL6ZWLpoPvyoHgGInMj9RWjhnPkW9KwfDCDzvQlieYPFz2Nekh9XpR78vU
Rkk7aC+l6Czyyv1vk2IX/euOwjGsT7qMwkW1lHNwcVb9GVaRSFPlXbFi0OA2
ySG31bSU58gJq3JeQn7k5Nl2YSLs/WeSOb3C0EA444gmMx44oTV0xsRXSwiB
r/XWzfgYoHWlfM7FklqDXrusm0gVflXNQgmycXAw9zJ0o1YLBDNoh85qKdWV
tXAOo37Y1j6lc/tRQf1FLfVKDNXfd4JXKYoFjDTb6aCd0DcQp1Xvrp0RhcGF
g3Pudz2ksqwvxcUJev6EmMOgd5sSYM5JvtF9RBGYZPhhKg8rMIsIqXtyAADg
4Sh5E2Lo6W9lmsRKTYac1B04iH1x8zopNmANr87Gjl1EJEnKOhC5j/rZIWv0
dxv8OBz/MScAVBs1Zg4sRDefGulCu5RRi/rTUn/7kuOWJdA+9BDrJw9oql1S
I6juL9OmwcIhV9suCOrQiWwhaGSM5H0i8vP40tnlAcyMy9inDmz63DRdiYIV
paSYyW3AGNwvIfDpTEKRUCFUKYTE9oSKCPa3zIMRooNdDRuySlz/GQ7VBdkX
r8RavRcYsQ1w6Ob+0bdgf1MkbJB6FSxb3zZTTxQW9IBZ92UrL7T6Y8nUYDFW
trq7B1J0foTc3lkYbpU1JpJP09N1WSFP5g+QIm7Zp7E60pj5DlvEp6K1nKcX
ycqEAPseRAtu/7lz12ClvgiLgnQzmtIG1WQUWg34mw+e3Ktdv9yCI3gsoun/
/rgWHLsZnzbs+AQ2KLSe5sb96ST5u0gTWz3gocW4UcyG3qqEpPFBCPsLykBT
JCCyY1jyAMH5FGgjU90zbFQT+Zz7w2t2t1GlIAVv1HfJ44Cti0SS44+axtkc
0wg0Svrupfe9ZJdwx/+nVyD0U3HA9onT9QHifvzhcB6/Etk/MEJkWFBA8994
BBhFzx65gyaMYgaTa7ME/Pu56oiHPfULj9oMO51u7Smpz6jsX+EtSujtzIOH
eTbZ02SzAg30TUAbFZ54oMbEtMqz7WBPI6ZdON8xP+j018wPOXx0KbUCqsT+
md3aKkc4DpRL51mWX1D0l2euFD0fPO2eU+Cum8uFBMa5xaOlcqK5IU1AKLxG
29pibtEMy2eaLDu/oNgifuWcOIKcr7wnilmcsfa8k6PB9g0nN0kGVtSfj/Lt
OLFNBvGy1JF+ZJl/CMyUILe8je3N8hWU618wyEyNux3biYkpWgWr9u4KsBmf
hxgv9JtAb7zOmUR2KdbZFdk8PkxWVz28VVTfOgDIPT0d11a4Yqj9+WxjrteV
7R/0yUyN16wsPb2BYnxqAP2U+MYaX0lwlJEg2LphxhADEBiH3BgMhj1bwbCo
dGPqVZ4rCRLPheAJ0Xf+4poSvgndiJCX8y08NUPjmqnu7eTjPokZxFzMOQFp
jSwb32q5q1WvnqBcbMc/rVFAijnqyAYfTK7mM3s+l/8CiKKh9RdQw9MBHQJ/
ySboebMsgjEfmjwOq/oGgSeKr1TXqOdRoIOUlBs6DxA4puQdnpe+DdXqAT8d
3Qyyc+2oEZsdiubShPXstZMdUvVEdjQtPHbC8DkEZFKQoWhU5lQa/y+K/Lrs
ezcHfdT33T5qZpUow4seADsjuorkUC7eaaNPz5M5da0dEekELllw6ZPsobnn
xrUzjKEqmGXTfel8HAl5BzAOnjtnOGhnc/xVkMKJYsPFc/M/JsPdfJ66WYF5
yIVXB4IVT9NCfU+yzkTPR/Pv8avrM+NtIz2deyXb5MiMc+OClxencC0ff8S3
zCR4RC0ylHNAdpLK4qX4LV5Z3k9oHRNM9s281+hgObz25e4o9MDoTQ9XjHzi
YwiMMkESWxIM90DUjrrFesKpzp7b8oYW+/vRBmBw67AnB/d9snqo41mkfF0S
Xutdo0bY57r3rn45+DM92MnKjEiT4HiHGv6H+pZnCifF/zjqEwOUJlnXXQRJ
+0dj85m+uxgqx/zw+HZV/3cnUttfW13u+TTXME2P8O2mzpX/WPlfC4etpP0q
3K+8SMKsE6TnBwDs7/FfyijD/OhhHkci+squngCvJvrQMY2+bdtmfPaX1XjX
2K+n0niZqMGxyeDWylaROCBBsfgyLPCkABgVFzGOo7HCCgPJ5/2OPQbndbVK
xc9g+zIm9TKTmnhXKQ3BmBvPvX2yobU1bTUr6/wjWqAlkokBA6VHNRdz/I1o
jBhevStB/QYr5mgRWACg+MA9C8TqkGuzgzC1hJYY8skmZLGgKVRe4E687TxT
NhKGA69/EcSP6Fb3Nn9WW9tlwE/QB0rW4WhIUKh3/iI/vldv5AXHxrhy1fw2
waRowjMHoTEYWlsKJV3WYiG197aVxYxov1q9NhfMM2KiDwppjFJvQY/GX0NJ
ZGI7mv/godwgXpOUWkU4jD+Pc5I5AuRwpKkMkW0VpkeEJNhGPkzkJEUD+2sq
1qbGc4ihAWa8KNS8rjx4lKKpf741OleyX1JceifJRqeEQBtmtfpJZsvWE+Hs
E5qCP2U7dw+3asQ5yVOzZeyr0Zar9eGgKHpwN2geWjOQ16Yl/wrKvmgjrCIU
nLL2dce/o31pqAOp9ibve6FCmvQEClbIv9cHqxF54oHI9FkRujzfLD/dJcDZ
99ifoMhEK5feorHU/ZcKjUpwmNy8iHW/W4MWCilApNSOyMZSr4IFw/j2WoCQ
BDWrAK9SQzes4Lz7T9Bn1vOs4vDzkEQRl1ed8btFeyKzlCdNeORE8EWtrrKL
Vu4tjkze+PVZjSET1N4uaivoeHZl5eDqiNtqxJcm7AzgidWCIFdy6XnAIGCj
v4WKxDIKNafJHwPJJhTNf7hD5wbZUZfEn9kLbI1rWLDFZT6aORLPKgqNIwtI
TXhrkXcbvvQwbKrYIE+P2W7LbyUMdYBhFYF0eAwmEUPHIf7eOElBpmEQlu++
c0wLdOibDUWWWVHxStnQvQ19b5MmF/UgDNcuPn/T0mw0qIxz9Tcq1N8y+sJW
2Yu0b1YlU4cvQ7rHzzyMzftIYcT9Ciw+ZCN+KyPxMdhbUjGJn0Zn+0NPS7vl
SPq2uACaTXg9+ORFmvCiHF2W7CnrLHMvM5j4ai9wC+CwluW1jNWiZQoOeXqN
Fmzvs9jd7ozyW0muRQmWBdZzKsIsAP9RtbfyzP1NfIcvsCNwQtwWwgClf0As
ZgflOA+M+QOs6eFvdl18DevAeI2EQZmpZk8RUIWNGGxZIY7h4Erd4Tw75S8f
adnKWZ/dEb7jy4YiFOD2JIa4WFbl9c+ui0X5tIZnRC9zpQL2mgJ6o/wmWPWK
iZXA+slnFZ38WjjwpYgQIILlhBimlZ2T8noIUc/Kg7Rk4D6G7mClVKUCE0Vd
ydDsrv+APr87NMCQCtGHsPK8zlhTRdAnmX5n9fVs9p6GFEdd01iP9UQJHhEK
At3dHG2cHLz6jvD8wGI2raunf0UkZXu4FAffncRYXSAQqwjuFWXI42sVPcKU
liqdaKzYISdOQLJkeBdJX/0k2+nFI4Ha+DjbhGpoDeDvqc5D4oyWuO3r/QQq
k+mqw0ooqvnaCHQUl/6N60Cd6p5VA8auVFbJs1WE9JEkwoTE/+SKMtBA6+4p
E38hUKL3lLYTVixvonfpSwxDL0aLw1Rr6EmC584vnjSsztyMcO4x5VXc4Qm2
WhP7hawQQutzm2dKPuigOjQ/0cl+0vqjj9f4bmM+qn6CGbzXwL6HRIK1tZZW
OsxjVhGv9LpHDUybwdFAn3EgNj5koJcXI/3C+W/NJMe0aPg50mq99VXl71Cv
A3qw0tG8uW7jIUpYLc2ZraKB2ePM1Pi1FKDgIOxu24sfyChtQ3+UyNsWh9dK
bW6yaezmGax+/tYCBbSYDioSSBcb2KvQqAjJF49rLTjWixiLiGr28yhk094t
5NOWONnJJpqQUX/gT3YS/yxjcYfVHWf8VTRSrN5XKrnn2KZ+7D1px9Qopc8t
sM51bQIVvN3snCfO5PaWiL5RuEXKpHPyHJeUX97XC4Le58YEu924iR+NtPuK
nIRC+ClG9K23CnKJy7ASbwcUyYXBY/KobroeEG1UeQGDztrWGaoK2IlqSpJ8
shKK+uKOWhO6m1BIlsKoQl/qGeFtK/GQJCcobEgGTwHF1HLhSk2FpRGIiIsu
TqWZEtn7S3xXUxtKXKAaLHzggOCmXFa46kzsorxFHEgBjIRhYc2b97EbAlKl
vDvzxS2NSBCY4UvSX7HxYpFqKM/7o4WBYGYY4uxhFdwhcoDneghvJEl3ZFkm
OZBwCtFVRPNdtMvi/uO9Ft4Dz5uOLnbJ36VBtpA7Z1X/Ms24W+LS2wWdeCoQ
m+RbBGgfyxa9IG0J6uujKrqJX7dGMmQXgQArCR65xZyqAKtK4Sbzei/AMMtD
mf4aHXw93dJPOgF10kzx8yI9yQWkPDP2xFhROHIJGIxEQ3N+7LXBIfRHOJgY
SCo2xCkEdakcVraEQmphO43msM2q2VT8dSWzlwuO+cOAMNTyYcmZasNELJ3k
Q0x7XwxE034cBI0tNOzQKhGAYlbzfjEN3uIHAmgRjwG51e2XsVgD1Px5JAG5
1jvfI8uh4piTaB63umqRuwopeHU8JET5RWajOd+0QEMa1dbW2OAGRL9is5ms
WKy9tS9Y5B2xEtyH6+LqCstHYQUrH3s4rW1DNwMEXTSGlnQCSCp48KHQ1DNs
fxcGFdE5rFap1SMHnZG4FzsAcosC7uXdQjka/hmthfyOFc3t4VZedTgnyig0
kciLOYfhkttvTmh+WnK7CQUKXlCGGI5gJQN1ytzRBBGnmnA0RCL3kRogC4zB
Da9rospEfeYvmopqSN2eAQByX9JUVBqkzVd/+dt3NZU0AhqsBA+l52UzOnFO
rbmmgG3RZLzXdRRrIltXOs+exo2ME+Amya6re5QDzXnryAynAbwt56+rFDyu
rc8rA7j6Iw40V47EEsKde5S4lRu1+du6o7A5Cnt2ka0DrBWb/6UyUecuhUko
qW/Voh0l4mvxh1F5px2FanDVGHR3KZMYC6rcVDIrCI+SQrlTJxHhWBirCSus
yFpCGnpfbNaK89uo4LOj4l2rgKp+PhTHk+JtkdnR8R1TwGxE5m0rKT3zoxcF
C3Z0MJwO7OkyJdi221fPpQGxxaTJEFZaa/21ZM6BGutybbQchjVPFN8qGiW8
1rW4V68woL86K+aYGvjobBE6AzFzmIRQYPtDCjZACSfSXjsWyuFcEXeS9+Vb
1f5csyFGbYkEpzW7HywNsQLWMz7KCVAiEzDkmKO1FtxK0g7RJFQFeUk7uzQE
prC3Em1JT1NIFBlf87XK5xmo6BK1qOU0Gkj05JKS/ZXvQ/ePxkQ2N48J0JjY
CDnhwnFDzQCCqqWJocHB5NlRhTzz7UrSU+uawM7pEqce7s9aSXHbkdNfgQ7l
gvml9ofQdHeDSXOTqqf6KX61oKOnL23hLZ6xL801sqCcZp8Ed0bWwLC/w4Vk
KcIGQ8e/KyS/BIdxs26rTqDsk8QhQUNargWyA0+EjoXbW2SigepIuQFvgafc
udAHdPr073tV+LYpAahAobSHVs7gpWUHG2Xh5/sW80wJVxrLbsiQ9EhUiglM
y7MrOFxLJSmPc06FsWB92Q3p42mPF0u/VMZYB1gT4GfvmtHFXmcupv/jtMGO
S6o+FMpb+6HCbOFQojYenRGLOL7xEWnHGZEFA7zwGK6BzzpGLbRWHtxB8Jcj
/YTSBzK8atcaTKDqoBQ6T3Ii0Ouh1X39ZZQRE4RHQYq/d1rPdNbRL3g69IeY
6xh1BoaYrd72qWX38LzEXfV5X0HzaC6SBs9t11ACDEZi0Hb8SqMbHR79ASCl
24SJ9vj5bqAwXYZD+BU8aEIwE33hdIYJZgPF5h3SAbSimrTh8PHw8UpyJOsx
as329M2/rGpVlgZ5sv0Rt1XaN4teAdBFmKph9lD1ULmtc8NsDmZBXIutC8Bc
wfIDU6LMco4Sk9UJgPnAAIZuqNwCT4j5I7SC/jD/d6BofXRU5q0+QnNfNb8h
eRC1aF2IompVY5bTuAvrSr/XjMtBHEI9TqeRKm7G8xYF9/S6soJUs2wJfdBE
PFmBetpPSYU2rC2xhK2aZ6GHnoWiW3KTmXi1R2E8C/964ynrU61q+myxweXB
bKv9Q2ZdC0Zn3tdAF/wm9zkK0GEyvEF8tc+8ww9DnkykbM+gFtLLxLvQluuk
lcMXNgqQ8c2R1GhGGR/sT00Ey0D5PgU4R03yVJhx30XK4cUNiKRxkdyG7PtR
xjhOSUvqjEM5loq5k4V+95VVKA0m1gz66oChN4q0on2ppQ2HW6eG0jpyUPvO
wo2BO8JUThcUb2EE6LMlzUC0mR/potiYzx/bUsxrb95fsWbUbXiw+9SwyIzE
QbSasBmV1Y6obXKWRG3P9HJSKsFHwB6yjt2UUPBc6faekxCBH8jR0jNCFxfB
jzyc4jUBM47vKhBKKgy1p4HLus6V/GIThKM67NkIV+rfTvI0188/RoTAI7L0
bLQPd8kT9Pvkj7K3/VuxVCC9rPguOhEvdpdwkN5snA7QPawhn4fATwY47bno
urKQzi1kFPQOBEEHXcO9nhryw7bZ22k/guJ7N71D00qYlxirPRiMHEXWuWr4
PMiOba2x/eW3dauhUq7uBrH1yTTuac8MCYTEHyyEL+yXVHWLrb4gvuxQN2Gx
ripRHflzyKVtgyFx7UCBCbz1Br5JkA/ruTPWlhTH0BN+PNezv8CQPoVxkeaY
ZzG6XdYXzZTHW0ITKxJ9afXVUo0tEFRdwras3NyEB1L0FVpCVtjWp75/kccf
amJ46/LT27OQT3k6huFw/o9AcFEZHL8YNai8iK9oH9UkCxZMjYJX27QUX7Mx
fuQHPYfTGu7v1dkxbiccYbp6XHxUNWzEPNoKyx4YIT2MIiQgRxBE3bTlWPO2
2XTrwIRddtfpgMLAFzn3073aJecrr7Ve6H11Q+T6plHpKsspelBsiwpfPWnY
YF54rO2zPZcpzvCrd2EaIBmUzOhZFwus1iPNdCfr9IgOwFRml3Gy0rwb6mLF
byFPBAkjjRf3tVfT4ulfi81op9El0DU5cX5lHLbrwhjUkG/joImw4zgLvKDV
a4P2qQwbBoa4eWKrwNYv9PuAlpZzNHUzwEGLECp2SU/v/0Cv/BRwCiahJJ6z
MzRCqD+DsdxSb+YE7uUy1AFle2WKZAdnx16GGCk3gEd3ZuhATX3l7Cw6tnfq
yIlKUJFpa1v/KRFe71GbOVVdDMW/GTju1VVtShvHxBcREpr1IP7q5UMDLA+f
BF4MeK6PW9V7f44ht0e6rB6T0cDRsJGtmHqWB/jiLfPOsHghn8lYAaCZEugC
9aEF2vVjGdIQH0wU09TaTWZt1O8hB+JCtY1EqkB3khvX8/gQGXlqD0uRhRU6
OSrcRRYG1hcRpcTvgZvP8mrKO4oddqvRoC2U73I4OJSitlRCh1fD0ZXVDysD
2K1302byqOzFbaA+EO+ZbbiV5SmqrRoI2KhE8MswW9N5DW+urCMTD6UEONit
X+kZ6JcILF4MJMamVH87ISXTu8/acjyrC0Mg6rcm7V3OkDACAb8Z4BLrAJzW
lORjS+EV3LyilyimtG2IvYVSAkhc/PRn+60VUCQMdNaPGjCGMUMk62KgqfZL
1Atspn7mXfbeztBWEVHAFxw5SJh6J81nXptJxsQSGzuPx4Z1+u2kGf2weYt7
U2wjER1zDj/tNIneGLgcywQ1dQwf1MmkaCsNGuv4wf+s5kfXEP65CMzrcles
xmlrzlk/mAFkcwy+BXaw7TStsYB1TClVqfqEzU9x2kEcMq9qGexRrmwzZSZJ
lPizm24aXVehNhcGx/t4KcO4PdQr01W/YQz0Gw47nDYIri45yubGxj7etPqD
KUK1//YQUz9mU4rk2FY0fwGPmfOqvmknhN1jTq3OT+1zrTEIXPZHixQYKSmd
nnS5WJzySWSMED0We1HrIEI3iJDiXPFkXsSkT//y8gChjoXt2IqjaKEEAlv2
OBpDAagjXrIr+kAWwv3tUAtze3/UsIK+nim47kGLP07UVBrci0/80G3v+1xR
Wt9ptREq+HewWbVLLHtsNytOsEbE4lQVAlv23zZ+o++NisLw4EN4XlT/MTFK
CyM1INXr5xRMLWR1jE9ly6C7Dg+Ybwsw9ZbnSvOzU3e1ofnkQrIfapr/4tid
WKROq8NDi4TQXmdTjhhQZQhjlFFw5nIw4LaejEb+FxJmMprxP5/gZWsAj6X6
LXYPjSkaQO4ZSgdzH+V7TTlHiekjIhoeoN8x+df4MYKuu0tCMfSJFY2D8+Yi
evi4nsFlAw9GKhs4CZk0Od+qU7b4Fr+kUJA5f6ZL/k52fgXFqKJvQeUAVNNS
8Y2hAd+HkVIMfWrN8c3Bj+aUPoWWMP1JZElFiEObbdWVrZYGv8LIj3Uz3M1T
OUvMQFpCmOB9+Tv7v5oYiOIAa3WKuLk1gLV7zL9fAUOJfyUTtot7+OAKA3zV
5zbq4nOWTSNJmOJTKDYL3sSwFyaaPM0PWHPp9eNmW03GmTYQNDe9SWkhog3C
OsT+CI32ASPmfk46r4HHPO9n84Mq2L12VH173Hg2X75pZ6hAoh4X8qWtRPlj
7i7xQh78OIhoeJIJSS0MLUoVKOgKIOpbRLd3XyAOgpY9H2ebdnmXCsmcA16l
Tz3MFy/HnPKAibVlyLruz4+Rg5mrUZEdGlM4Vo6AWZ3/W8V+BVWDTVIwtkRS
6jm0aj7QD+6jB0KM5tKeLoXoWcA4IrIkQ+Flysj5O6KxFXQRAWmdYuTiE22/
rbjeKyI8ogWMsPTqWbylagSxRU4JQ2fH61gO6G5IqZFx9PPqq18lyYKCO2U8
ud/scMqlutp7tjHjQeyr/wR8Ev/sNmiPzfNNyCg500roxAxEbBmc6Bud3JTu
JDH8LSCr6J//ingndgN5QrhQsOoWkhwANXNRB3PvYqwBPzPqr2e16CEq2EG6
MwVIdVDMMDbCQkm29porxFukU/RcDJLcEOZBOlXPPpGwtUm3+0rkHAnt+zwE
iVH0gkK1ir9gNJ56sn4+nLDP4rX2kiag5hkP7hfd2HpwVNsyOg+7RH5AxvX0
p5h1fMYMbLS6m2jNxEYyTtQ0uxsE47a0RUNbsdh8I6k6WfxpJ/ir4FbFq9Hn
bEAGlhzZX3oS/ghUFc9H72JkSGKIVIUflQPSXeVjAEyX7UnXffrT0Iyz0RrV
LJLY7hFdf3Vu1te90aF/45XCQmPu/0vWm6I3MiSWUtcySqMKMsdR/VD2X4pt
iARJ52r6jxGEbyUyBW3+B4aHon1Wlirnf3hrVipH5SXBhKp5GEdhqLSlOsF2
8oeostpLxTXsEW5oDkwFg6PkIjf9OZyjUoFnnWx21Iqodhas8ymNAABEUxGo
otTKX2bnuS4dSQBm08IAx6/pLGsRN3/LVYPio+DRRQbJKWJGiioo8G2NkrUj
lqYbgc6wIzmjIRRIoAHyBJoVATUGN98TIm1FtlghVSoaa5HFsVQt6zr4j2Yg
ez2ITUTO62sOEIXXdZ381G63hyY4XgQcpyKoRJhJEh/U7zPLTU+H/pZ8tMbv
2SBRjQhdY51wQAfcl+DG31zVWM4/GoDjbIuWW4vafmzhsCOIc00JnIPc2j54
GTKNQ83JgVx/4LryB1Q+z/gvjQKVEPZGMlICAgDNFbqPmWaAen8t67ph3XAO
wIslAFBPu9vowbfmMGdFbGLk3SupJtiU5rCn0XMFQosUfoW96WHRvcqbmF08
7odrCNwKEIcrww52amsogMJcmWFfFJD3n3emXjvRBw3ziwvu5vgLd6w4OnQn
aRSqOo+zhNm1yriuYp/wYTdeevjCznOS2j2UE1XNre3+PNq/VXuRni9vWGDI
/eV+WlqH4PugwrWLzA4mRVRdOUEE5dUjKF8kbKAPB6CsgPqSWk1H09R7hevS
GqbORunPszIMyaUMI1mU7yxobJt79jzslA1okEipBiX8541MSTC3KBXdhrGe
NbD3W/Q5QFkyU4/O9W/4cSseON/ZK9uFQ0gm+yPG10XHRrh83e6K+W4b/Llk
XbleYcsqGA5pKfBQE64LuHgnbyUJnk/8gkn9nA/DOmT9KvCn2AGndsANyU5C
O6MzSR9mzjKnfCEeF4FzTeVJ3FsZXbB7dXTrjzFdqraTairwLgT2xYfUuUEk
9g0NppigvbvNDJ/L6+uWgUQLyxnTNnG0OhcjEFVMludxcuQnLxWGUw6Cgccm
UTzfF5Cu59eGgmemVzeVqXb/Q/G11onlCiAI5z2dUXIA0y0d2Ndg8VGH06bZ
A324El+XP0EGmOYjH7CQ8BTyuj5poVTE1opmWVC7UvpQbx0qwCrOvaWr00iP
xD4X7+LVb/++rAZNYg3xM7lPHaqYEq4fZe8d+FYFxVCyy61v352M2uEJf+Tr
6hjmDiN/mEzIhQWXxGu0nxtlFc2HGF1Tm0cmZLVPlmbyGkgZa/CH2tjwGL4Q
hliyf/c4GiiEQOo1ZvSbCpBME3T9xQt+UztswqLyOfbUrU39SJQiKSfvs1Gb
eaYfZhCrNX2xIkZVtl5XQiRkNSvq6878lJeUmZUGFzl9GFL7cRy1nAShvbY1
CZ1rClSFm2uAdtaMpp0u1m7qGR7K26ImpY9JDUdyGrHUEwzt0kd7pSDSl/2L
IAUhfjxoH9ji/qhvITElApc2Y7MeLFaGscV/aGSpVLfb5yabmaB24A9m0R92
IjNJm53uvCDBGX4eCQTAwgc8w/DqHP2A8jxRjeBR2UxBJEIRvhVUhsOIJfO9
+p6E2TZ0ZDMt9UzJ0QvPBJlA/lza9YHaEk/Bg0A8dWrSv7gHathnnSvTvrPK
O+SI86h+Tn9d1xPyWAIsyBnuQbQ8dhw2dvmMOOGK3ve9XUwiPZ0B2E64ukBo
V7CyKshg30ArAnrWpFJnnlI+ngbcet7cmrNfMwMYcCWLQFAig0E0xiftfABQ
ZRvTYeDoUda5UGqeUqtUm6yBhHhukob8FZhO1cwYhEFCDq7GaTIJt6iMiysq
vRwqXVYpTG1RhM+k9aVQXgTHCz6LVfqPF4qb4FuJa6Hz+1FQ68PN48Gps1FF
oSU2Hemg+1qyKRAkjHYPWQjdNuFcaYPY8Vc23lDzwwtkBqys04tGzgWlripN
N/4jDuCVJp6A5QXba9t9VDo2eNmrdGDXqntO3Rcly8/kCr+2PtRxJ5i+pOcP
HJit2KUY21OVWOR6V5CRQAUOD4JzCphEQHzRRkmXLMKnVuoZHn4rHfdKTCK7
KSn1Mh57jfx+w9FFR1su9yBVXROocupI9rJ9IswbI7DXcj/av2ZU01KkLX9a
hEn1Nuqszas+Izl8AozNZdR5N2/CJrjM0u71jqB/rLVf/xCPw51UjJ7Bh/Mj
xXrRa0/ssgST7fEAjEiyDD88xQGIhu5TOpIRBW9smzFll83b5OaP1hveftKr
ESyKe7lQmf8x25n+XhZqGjIL1GeatWqlasdYA11/KUqd786CjbFM26oCfy3u
oLmJlETJTk4EsKLa7o5K4mtFHwXdt97yAGIdCqYf1/e9xEGvi5XrO0u5RuAJ
wpMC7z4mULdauaY98R657qN859bY3FDaZH3u8p7xAsVv4HOIJf8P17ijrzau
DfXr8vmktIGtr/x/PzbkBgATN6TaQ3M8jDKoSteEF8HZQe3HPpcdeyWGLlvA
sOPPq9nEul1IB+IFL+5tuira7FinkbGo4pC0sBa60Waxd7YsYmcclwUgCLgu
WImXffp1zEKd1aumgPkZtFSFXETB628qP10dbmX1gO2s2ug+L9zExr4KLMIX
e7oh8SkqoT1MjKvIWi+ql0SMfqBw1rgPxgCOz2NV2ogIY2F6j7PXpM0MRLIe
Pr2jKz7GyPkwqUFTd+pCpH2PANjnxOvkOdVwzT2d0zYf5An1pKMbLAjtW/kF
Af94shm+uR7uIRfak3QvOpSZ53m3OOYsqpkwr5dJQQ0ZRXnm1fB9if6QSkrc
5PFRiFJOlp0HmRJekj6V9MEXmktDYgPaatwJD00/Z8VuLirlcUoZ0x73vE5a
3VFVDgnoOXmn7hmvGC/+n8zLZG5aS4aU9BEqhHFnXyDDVqvvMYitGe/3Rb9o
oCWH+ZpUH9aVpGvjzsPpw5liMBWF1PMrZfj2JxOU1ImSZwTJFF52TGMZWv8S
j/qxEjW5w0KRuX1BkyLZZ5UggGxlvYmLpFifRDvogKBOykNCsiq5vGAuu1/T
67DqZuBV8jdfy4HKMdDHY7noRvoyPxfWlbeDmYvTe9IPIlBPxvKaaN/puS/Z
Mk2DTSrTo4QD1AoVW+bYuFGTLwx4QWTpnTuyoAOKJISiCv26Vmxd+CK8FIxS
OAY2rZL8wDgQHUMUeQxa3zY7MDfjE3omuonHNiPj1+BoYhJ+LIh7lDniDFb8
PQ+rOxXsBkWGQXLQVA7Eh+s/2LqxXehHVpTpLpPnzGoYIUvMQKOuBUAOveNv
D0QqpV09Rj4jeot3W5PuX37gnzaGBFt+PTGci4Z3pYlVIdsaQQMQUcwRtAQR
BFsHkJreEtD7bL6wHHSnpjWTuVJLx05kwsGEfNoa8YRXroEpcll1Wtt6nRjP
L42Ft1Fy99CjMSY8AVMpFFY2eFcck2/4ZDGOOyZmhI1Eu9IlO9XM2+l4JvcZ
Ww1UAURg/ZCoYGnz+D1G/F9JikUZUqyib4djGIbonrnV7fO5CTEGTukCMpMi
CMNTLbzgAFkaV3le5yL+UNHJ7bAoAVTVOKboKyH6j94woSIlesivNrQQ9Pie
unMNqOQMyv0KCjmLZsNlmHl6ykDXcwC5W4lkJTxulVJKxkqnRjm6d+DNg5mr
G8lIkuW9iUHyihyG8v9y9aJkN2ntZcNLjg0a3QewLXsBcNq5v5h71gFTmU/r
lYBKfdE7GumCAXV4oDh9BCefBYMrRExSwNzcefPRqb+j15WG/xCVgghGphw4
La2H/k7HCtMKQVkyBie5zzc2DjabBVYSMmlPt658Kvp02fmv5LvB0C0xJ9q1
ItlGlLxBPBBYEAgQ3HRoN9JO7yi3ir0D9sGJmPNwA28dzCcaN9wli3UwiE2w
aB8bHxuCGkhlUllzFUJvZB+lynfd8kYDbSMWxEvRSS54lYiAuYQKWLaBcPYp
fz5v/eIHMnpunm2BZTzf5cipi3zF8HeEExOYN/1Z7o5SHC6GOKBsmV/pZ2Nr
YLLkAzJxT+M6IW5Tg0HnLEfBKIGRxGh2oVwAAktaEar6YGgc1E0S4vufoPJF
MjipnwxBr9CcDWLIiKlGEoKhWf/ggKmLfIXlqMaEaSMC4ZetBRdapkRIdBF7
ZcxKsqskVC8c5nXRQHqEzmrSy5CpqW74OCbGnbVzqfyQXzXDUe/5C34KhNi6
R4luO6/DC0xaol2uMAWxQaUE2MoNKFSlg82zdNGiEwd25uUN+z+vaYsQocPk
obmXi1pe4tX4xvfpyxoOnRNRGPHOwiOHKui5ux7PSaG+330mgSpL03ISznpH
40Bw04+au99eh2DKhFrlwn049KDxm1StSSU7FsKaa42vz/euAwWIigDEhT8U
qbVj885sfqZomeVpflJyrjBKkUVyuNCDzqrB7/M1LGVHnaciDMA5sgoMRw0v
8AcUcazSotZZyJpzwQcrgvysrc5nbS4FSVqrvUrTFY6Lt/hoKE4CflXMOT4x
ON8r4nUbmTJktBeo5Z+iojDfXwwRG8nA+xlmd0A9F8Dg3VGbDbA0wu1t8Ov2
JiHlCGGD0euKw/kZTsDXPtPoQfXBt7H/APze+qCD2In67QIxk1H1YpKVIVro
fDtwCwLV/vy/q8fqTOWwzUjAX0S5mosH3DJXlCkMmSEGrSB2ElvXIJk5lZt9
G8zmdOL6UR4VZG2sszYQOReEgNC9RaYwYSU//q5jvJ4kUNF4Q49Y6JDIqyFl
9QnViRdsDTJXVsXDPgHaRU5TSIyfS3pa2Jm1EjXnUP+N9kWW14X3sDPPJ30b
35BUK2MSkFqb3Pdm9H10lsu/nb3nuYftKpzd8K+KwmANe9rYNVcN7/GikhgT
2w93PFPotPPURnKmzhnqAADj5fcEit9GKJXCYg7GwsNPwQiekZgg1qHARYuz
yeVHq8tN2Wm83cS/E4bXEFSTabFj9ZuMSGISTkNuZuDHLuc7AOosB26Qv1cS
6c/0ClpIKxq3UFpRNb6YAZQ05q50KV9O0+6TLKny84IRLMtqf8okwzkzzef0
0hN7yKjP/7pvgXCT3I9h6mGGCXbyHLFvLvTMf7kmsv/EftEdVNNGSP8CoGnx
D/3kDiyFM7aaZN0GcVBjgcc78+vQsVT9FBaESuNwpbKrqPPZCYjqn6ucoYSf
NjNgjRZLKKxRMHmxtWdH9X4MpODQ0Cym2OANHCNu+ypbXc2rLpLXoLUgv2h6
2GxP2Hq7Q2DDZJWS/p7dDnO87fJ9yR0hL0/uHQdiz4kCSlb9rsOC9IjOZaoM
fl+Lm/lMJbrfOisBGerLtLyPRT1LU/KwzGZjzVzfPKkNQBgx8O7bZRrmxAGO
6sSKqf3FpSv56BW/GIyX9HudERSLKBY7dLKhhGSVuRdOMd8quspuufGn1kpW
BGG0wfhyR1YpyU3JO9JjrSCdW3/PbMebg0Y97doGsyJ8K6wgRub8bzhpRUv2
X4vtYLYZV3l/GUGBt0huLqZcAiyDyuYghIFwRkafbMLx7zUS5Cw5oFJSwVop
GuWU6JoAl4VZDMZgUGNhd+Jgyynj3JMRk5ErBf22FgxfxXcSzTGb0msnn8z+
PdLmrN4+ipTzpknNGTelwA7jwZPKUUceAvmxD7HDfbqR/xAXJPJ/61MwTuTj
vRG5VgRJ0yvW2eT0Jn9gHD739BB2vY4r9E8W/NHBpFjS1cNmZOEtJyadz4DJ
SN710Kf3Vw4lhrP6u3l/ap29ghIF0+ua0qUQDKBHGoQKVAsz5qRvcGDqOom6
0jVsSjMIUZtlwK5nQYqFtuUkxB1CENldsi08dPYMRjzyjvw1DcC4VVp6niB7
6IT43a+m7f6uRGU32Ke/MKgbmWBSFDeQVHuNZFbo9fqoN4Bw1sIY0l+zkAU/
wtk1trUiMOLP+KwJewyAVZYqOiBRUVrdnZcCwyAcIoca2buJY7hxPnIyu9Qi
SOnNAjRvB7SooYWCJlIb01a1BbDdRR6sAn4oDVfpQ8dU8QNwy3AMLLW2XNp5
G6PxUMBRGMDlGdnPYILCremtG+luowpfVRyQGTmg93bfeY7ZLa7PMLVA3vgM
AWst8RZ5p5T4dGKpMWPjt9mt459bPFBPPw4A0Z17AsjvquLh59As8u75O7/w
Msa9seLVgwIxQj9r5ux81mWoXdAWNnImhBHDxXge2Cmj7+FOG7r3NUJdPlNS
ZPFm5wFmgTZOvH5ffjkXKMuKBIncGgkiDwp3Tp92vKd9yZ4uSnXwC09M3oRX
3KsG2Zaaxoumm19j9cP4XVVfXsrg0q6TVZyuzsTBgpJ8Zv46f7feZQ84Oql1
GU69i7/ElH2qK/KnalOTvSEnoboHZ5glDAjR9wmdMqjDDSEFUD4rCsn0z60R
285JGF4VoomkvsfPzuWg6WirDgBxJzBniKpMwL1+vW7YjYXXmzV4COmSkVn6
SkPu5vb/1wvILPify77yS7s1mxnmdPc3iosiPLrSJwtLBFIa1/T/KiKuCXDK
Q1Yqg4+RsokCaiCGTKFXB5RF7QUCODbSM24L17E2lfu7+bLKH+3WX0MghlFJ
nsn9oF9RNkv6oYPfZfj99d8O5wNztdJMM34kMZ5u8YvUD55d5VWWg87P5Cyc
gF8+P7dZ1F4T58SLkmimBZYYVJ8OUW6iKJ7BC4QdasztbfJMpBQt/crHbWhK
4NQZmIf0YtfRkaVM92U8KYiN6wQ6xkPBrnH/2nH56OskCy3oWv4JjFoJPzoJ
gYvFPZxDd+EmEhGvqlyQmYjyjYdxyckXmyZipTrl441K/TSWXRMEj+DdNxl7
/lzOvtHw/+I1ckBEfDX8sY0fEStCYAIamuIlJygGgxUC8BosB9VmYiGxFIsA
sC/RKBTv7N2Vc6T36Xp0F8Zw4R2Lfnh01nKXlPaLgpxbPEpUgb8PWpckv3v/
WgehnXbNbdDJA8QekTtgqeJCInQlCuBlNlqmmCmWCD4etyhgI+AP/uN/tIAm
LeOg3lmYvsNDZKIO4yGi7DgVFbImTLG8S52dSBP5LYZhO/VghEBaG2f8whIB
NM+hvW67qxIX9ERvzlS6g6ULD2JmaEL/SG58JDtxC7zUY3Zbw3fXLLZEyrjN
UqX8Z202e8xVbAQztUanU3Tv+kKdvycWEfcq0/QbEdXKtRGf1dKAZaUUq+PB
rOYZJYq9dwJse/WXHxGwKM1YJcHYXQGqkyR0A3M7UN0NfNyC11SyEJ3SAQZF
4kxRi6pZvriGaNvDzzN7RzB5JNbl5bw2EMudJuC5V9WKDDo0CxDYX+byBv+E
OmYym5VDRzaXZmpEcysnPidh2j/BziyiWwA0Hn4BtGRmDRM4bGX8ToW1lz9N
S2EVToQU+iqD2b2prB3B+084uQAzYVwRW6z95FRzFxsq27HI0kw4zwwdBS8+
mhdOA2lvOu4Jdpjc96O+NN7c//Kuc+Hxi6skuxymgA55wIiMC+9wA67JqtxN
UhWYfg7qsDpkJ/ZsOnjH0/iNHcvxNvuzy9RiYIAdXnmDIXDzgjMAmQicoDO1
j7xxg0FGfHxJ1scGOqVCQ0rfWs9S2fzPEgmBe9ugEgepQVByQCytGZ5H7zDi
YR2iNhiTE+6/AxuYsfmUtbsWo2mUU6dyWkeOvubzbsq72Xyj0SaB2fmgYur6
XCnQnowavLu28Yvm7gVsFz1U63KBO9JEv+evAUo9BxtZn2NfqUy8XEIGIVhj
NncpVncO8pe7DOTV3W9/HrJh9GuRcKzlcsYrB1v4mdIK7vg85b1gswKhV3rA
BKZWku9eoKsdW4tPTGQxE5JWldTwHzCBEbWLgu6cSbMpibjmFPhbiGC2HOB7
rlwiIaQ6gZImZK2dspbmn4dTP+nReZViscfC09XfCGZGM+MtNQFzpjV18pGm
uD3AWUn+VuogrqCjPczACak4/B15UHw2DCieODLVsDoTKPlDYgPFCTFmIUu6
GntJJPhkEwDi6vC104ocOfXnALVdNP7liTiPxDhIH2Ijv+XD7IwOewU9Nw/K
J5/SQdIs6MW5NN/P7nTpqOSSeRf0dOaV28Acc0Nm0Cy6MuB6xCOrEh4H6Mb4
S5pqrq3Wl5RzSY+C6Xi4pWF8aXJDyfAep1z/EWgAH2HXF1Zggoc4SuLGnWFF
voQELoepVJ4+Oye07lmieF6qozZ6UqFTUtFciZpGzybgsXDHMhgPldm8Ahd4
j2yrlFCsVfGep4ImaWK+N5nleb06GAdEDfcUZflMJ0TYdSAQHuDnjAPi75jr
CK3h5PwLhbX4w+/pVyNRhnPNViCOXtFXUAz2N0eDLbE40ZLKRUznwu8YtnZ5
cSQvqqNhcmd7Upse4sS1HbeRwQeTDeUaBzLTyOl3aXjuBK1nGYQlTTIuWzHi
pG/DcrSeu5AtH3peu20vTiAynQL8dKyNoDxlbl5gEdYNEhY/Gt+fhkg952bw
dClSWrlm9lcRSOY0hB1B8rfnjENFs3qBBlfoqufzcG3zjs5NdFIW9s6C5HXO
CPueZjjMN3epkJrdUFvld4Jvo6fdq0OsSEBQpCVhN8MNnp7P7LKKq8qjVmzi
2xSrbuAAbTO7mgFHAOUaWuaHjb9Z89SiWvNN0BYcB8PuWeUe2snUHKxjlWzf
Mw3o4vXzURnYtlcgMv5Kmf2ch8SNQm3gqhF7lTZFpPNjTX8hQeb3c0UVTDsS
JcnAgYJ+sG0gd8wa7f/NwTIGUGYZLVCGsJl4/ewUW7oReRT2phktlbvTIw9g
PyYQTrbAjCjbvtk1HI7lLzvtRUVkEqK+0q7Cu9CyUWoIuviTXUot80gx2Xo9
KYCz9qNJVXUi6u176njcxUj8t2fSiqmoMnGx2lR5lEdGa0sPmt07nvJo/7Kj
D7qXSd6/bbFTuNDYP13ff03n5qMB/eqaQpBlLfETvJOwNYFSa+s8jEiXmTKX
oJWwRg1rqSoHKLa+mFbfX8KhT0Ga7sJUdNjXfu5AwFP7ymlGopC3t7BPcf3w
Tf58/UW/g5TdRe09KPgzbtJY5CCe+rDMkH+uYnTRMNEGl0/SdZc97kMGller
GTT10l5gimHj5RV4wMRvj883ZS04j15VWr/bFhQXtoPatypYIlXj9QN/F7/W
jN6YPJ+Fmvh86vq+L+O+3LJREUrOaElaCDBsQ8xmo5wwHu/Rb3z+7dHzNj9y
tErSA6CmIszOzh60mmSiLg6TVEGFBOWCU/iSMqzvmzQRZM8y2bFgGX3M73Ml
LX292hBCWhkl3P69Q7KC0mFBDazyk/GbEF9JENFT9HwOJmv/Wy2qpHutBi1h
+OnI9DdGU5sRx8CvJPVQCvxB74e0+8+dMufCSWGACe7lWwyhTF1m1jD+hB6i
odhxm2eisjObu011ylFYpKeuNjkWBHJk1OeXpMaCxNkQQ4nXhx8NrSHDd5yc
lJkN53XcLjurIGstGNAJJAN2k0EKhGLOpWE4VRtW282Uf2yAK5C0mkRuvuW9
ofneTDXbNiW2y7RKCYRPbPNX/AbwdWGiNkvnNiz/e0PlYse3FGVuTgSKJdg6
cLVrW6ZtHC+GbCf0cmHN1GZoQQ5xB/gY9Nvrtm+vdXxWbXYRujcYlZn5Wm6Y
yMvwn1SILO7irSzPGvf7GLbhBuW1VS6cgZpLPjOcT+qdnEVS6F0vq3iZZBe1
EKZK8fGEqmjRozRB06j8utUWnFxEHVFuiyy0GYbUWwkz4mb2UiKmHBNjlv0/
mBYYGBUtdzQxN8HyyrPnFf4Nxacfx+U0SrwjLnf0mH/BhyuxKtTytT+ItEr8
7CrxEbIuy+jNclultUPvOEoUKiKQOnFDa64+E6NAZw3BiQvv84WZDOmgsAAQ
D2Ic1o5sK3CPqRDHvbZKsXnL+pNfeVL8GLnWGeAvlH02VsKBsPSf4ksLRaoI
AIoOu2LbAnlpSTaEWooC3BdndhunHeXsreWYoEVgzzgyn1qGcFNoswHcf3th
xpP0vt6Z/8IvomtFZ+rx+epkHgyZAtPWyUDLLjmO7Vf6uP64bXNxUfCtTuUk
l2Z01k9zGFHBcN72WW9/U/VRkv4eDltQ0s8TPw/64wrLuAAe3XA3cWTKDjaD
B5NaJs1y8mqI5myjhSX4XiUIP6LTY9d5skrlvKaPnY8ayLdcCas9hSEYHJz4
amuMh6V9k6ZEWVMlIefe2gSiSytivrl0N0y0Y+jrZtEkIkt0VPFBJpA56mxT
3PqhmM9K5YBaCrgHfz58MqF+HB6DfElknxdDe2ksV1LgItfBOmL2bNG40547
54rc97bAP1S4t11ZaqxrfgbMq4gTS4CJpN+vS4oXl6jTSp/O5xMw3Gn7TzD9
2sRygeh8NClZ/mAwMehjmUmcbd44QMUIRq+arii4hy9gLo+LeiZGThLu5tgP
OuzqKLf87hTH12M9FRHL4HhdTcCeGKbTgfpNUM1jTcGp+JiUnsHW6UBsHU/Z
6IBGG3jMOJ5ylgNBXT9lt6HvwJlkEfH9rvOt0qkc3G67V0dqjw8/bPKJ2LVG
iSGfcgMRmNiOHQIBqTL27xVquJWUwbbREIllfV6/wYtcAHPPfEOWJTPO/9u0
VWqwo012Npq2JnGuSUtDDECHSrpMu0PtnR+qkx2h/NTcFTqHXeZCs/H55p4J
RgXi7fYuHkK7i4EBJ5xUn2zDmTR0VY8PYatx097wZlB3W2+sedSAaNwu/NTM
Kc4/nBexdLdAzplWaAaIQfYl4z+T3033eq1r1wW6+F+N1QDSrVvq5V0ZqvN4
7xauqN/AoB6hsoJ1v9YXeo5UvVowCMuJabr9zoMKvE1767NDrhjmH5AmyQuJ
f7iiLyLya0tuA9gdXac2QbArxcxZR5uH1aUBC45Nk1GfEpzRqzRVNGNv4dUo
SxCJUwnaC089cv2ZZL2U8vUaES2HiDBMTH0CaBckfNRF8vxJfiK1jhffBwTN
gRGRTfDV/74JFWbOeAuJO2b7C3vdZYzDkVvg3Hahu3azCo23FWmT2TTlvGCE
yQCuFHKgKjIp+ummiD/iIPZBB0Q06WFaQqUSq+KR1bczDbKxTFSqlx8HLbO4
9WCYSjD/3YvoxmAZXp+wfsAhaRJsxjs6L2CR4XMtzyWOGZPrHqkO+iJVxfEF
jyHA7kjfT24mp7klTcKJP8uinpQqLX/MxxPNIiNLGU46K+IEu5KwZ3bGxEMN
ffUxolfHivoWVAaM43KDuef2UPrexGdmYy3wyoc6YUiDUBfsFxsxtycXryPd
5zdA2zRB/IKkhYqpEHkiPSjeKG/3DcrtpTh2ojX+jeuWzhUcHqFTSCyYfKpd
s1IIP1Xf0FNIBGPT6yhB/tYVuVadPAbYN30NJBHAB6YXXVtyLwUokyXkXaWW
fXPxG2G3HNSv8wIH//lIpfNVMT+SFVBKVDWITlgvwSqkpX7+1yPJxVvWkE/k
cA4Vks5p+xp5PywfLHxfoqiM1WSlYZkyrRNBhjZGysDnU8VJu7Q8UPruuktm
LHH/e5o1Ba7CJ/OHzxynA8FGL69HEs7DZTwUX6AxONKWnKZBFYu+Ls2pCJzF
fT5pfJk9hqOavKhbm8BYZUvlpsdNbRF5oEt+sGcEdk0hVLrTf3XhDHHBvOvk
VIW9oxnIY6E1wp9ehm92/uYgefWpGtXeTTCfx/oXF+x1KBzw01Km5Tefe3C0
6lUTyr5swJlbqL27h6KGF1hSxR01NhLcAE359y9MukqlOkegOgbj7+Mzy7CE
paX/QLIUE1rVyb7NUAYImFwF+BitUrsd1hAzaJW5zjJhzBRZ0dvXbcziHvBr
9co0NbeLEeFKJnK0WiiDHxprwaLqN4yLnQXFS4DXyNmGVKcVWqALXBmKzTeK
9p+/atNt9yA6WYLpuo7zRfLh/qD4vim0Yc0kCJz+J18/psNObqca8LCFp7cA
tI+ZxyO9hnKU8JEIDMyxmxXP8LpKF7fzujNDVx89DqIeJF7cvFhp8XatlKqZ
AGFfvmSMf/6V5vT9aTVflkCEe2j6eJ/pdFqlwzCiWq+LvKi5ibzwUi06JA+p
qQ54FFCPGlr8kz6pTpeTsCw4ohEu98YdG+V1Wc8LIq9puvtsSzenyC9LUJIT
OtopcMTCoRZjt8Xej5tZtcaS7cnN6kXs+rtbEFNcphAX6yPjVJn5QVCqkdUU
gNVjjqmdfzQdgdlMiGCawK2EOQTy8XQzB/GT6OYd8l13aiP+HfIykf37Y3Jq
Dc857Tp5TPVdirdeA9nZ4X1LaoR2AupydMLQUwQT1e280yGYsQTni1mHDziw
BH5fSiZMc+VTqWAolduVw+X9U3AQRDBK3KfEOTLXNsaJQ1e9NZe9fFXIWjO0
qaZnvbqMagrdy5+PVtiQnDQagyp/lNkn1teXVuCEtxDqF3URSJO5IcwBVjg/
8cLwDn3MQcmow2p7aENWZ6UzpUlZJNMd0dxaKR/x1LGmCyovWu9VBnPRVm72
IEPcpl5ntn938VFMCj8yaYuc6V/GxmwIZivX/xaC8W09D/G6bsouTkKITmaO
NmekOV5C4E+SY11ZWIlKEE9RvGEUONzhDcyL7S6kZ3fxQF3OW/Hjuj05caHX
Dn7vanM+gomZx95ivzBrsjC1nfs34E/H6qSDTByJVxWqGuEm9ESwjjCcypJW
tVvNrAtaSVBnYKW7+P+cGM5O6IB7Cl1+fKfinpBqdOTrx2he5r0Ov+yMy0k1
WXN/hZIVIca5LOGuJSxIhv2UYNtxU0gsstSUgWNLU5qEYyXmqEVxFUMxCBYg
r42CD//t8tVnHuabejTBjFWawtzzHCjevchE0XHtf/P0zZAbsRFFBJUD4GrB
6Ip9BUeM6Ib2giuDiLcIrtlYCYPFScZG0LqmZnwX34mq4xgG6r+u13UQzyXy
wTlJa21Zy2zrlsP0xFQi/bF2X3eryqrmvx5WnbtTKdR2ZaYVTxiMUzHgDB8c
5VBTuk6WnWmlUUETNHd6XqOQGC/d0vns+vKlZU8GWd7xfRMTw1yJU+fg2yof
6WD4fGPZeWS3IMRk1jC9L4yUv1/8S0znhS9DZKHS7gQTq8ug5C171HH5xuL2
uMKbRt5JOZknMpeuXGorFpVHyWbhbOZUNIPgo0dhLnt6C+y2tEsxjVUo17hG
3zUJtpuYBa4m6zTT48HdgbOFS+vzsRpPemZvN9u4K0BsDzWG7VYpDulf2LfH
u7Q+0Ds2p09H5THVCzNM1SGm1hgAo0INkye7wEvHpD5Egd8LFpR8w1OUchw5
crZtr5NX6tON8qvImGQu278QgeYvIPPMYTgy9cQrtT2aGAFBwbSeetesOupn
B73gCWywd+ez2z6AX6tGHl6A8bMI5c+P2P8EtIeJG9PJYVNprPKLTK7mo/s5
gZNVAozccPI3yoSX/UCkxoT1l6tBjOnOzcnJbjLm878xcy9ZcfjQ7nyMp2aw
EhflrwC1ZVKUkyaQyUFcpYrIh1mbyPpsit8VYESt4CtGy0Ce+hgEGRlCkr89
KYaswa2sktgOVU8HdJkEPR2MnA5b+ECt/p/MmJDW99l8X0englIfPTb2vvfO
j7HvCaHR6XGHJAzendC8c//J75wy+NRFfLjEj1vjPmeQD1E73bpmHKjZWcBP
j/7mjBM2NK7zGvgsBtkRBcF2iXzAEZRpie6XTgtVPez2wZKIud2yVyv/ZiAw
+ZeQiNQFJDW5LGN8nnOwARgAXKNznsL0WpXOm/TkjuioditwoRDyLW2Ga2u7
isEMJgg4G2n4TQ8CTiSgzdYPvJGDvYvKbpIgqPaTSOjpohXtp4KQQ+gsOD1l
ORHR+HydxrqhUJNVKLIa/LKbdMdAoYh8Dol4e7dcyv2RNPjw9QblmnDF3vQT
2lXnOJVKNJDELoNDlBSVgZn87toVMrQA5yM6EDlM8JffnldHw1ly3xitk/FK
ytdGL749gP1LZmHDOX+htZ/BUfASVnaPG3BhCagbXzXN2kPJmvk0XjG2nEMs
/0nT9Baw1jGqJGkpAo3khfZCL1jwvTo6ud6tH2xSJCgfcdpUkuYnxS7V/mv4
+NSyh92525khRS9/pF8IlJsHT5d4/2wXrWoAdXRromNaV26VCGZpX30ZtMSK
bg0CT0IiWWYO6aXfsg6Y39gLCwqmzVHVrUrb7uxFVkXNO8CvDNEvzvS7LoXY
wzA1IpK8HIEPX81Kb1osuqZBFZZE90nCsB6Jnc3q2eAo05sYW3WFvh+3DKnv
JyECHGbwRsjehiA1YSai5bx/T+vzsM9t4b18JC9hUmVfpZdCwv62AZVM5ahl
BKsv4HFfDaZAuJxVwx083aRoXBOv3GxzZ652rkRYLm7y0cLKeyJ5p08ZkOxm
yx30u5RyEhki3qUWuEzAxhai8JaP7oWmM/jspeQU5N/v1o6YT+OE9+VqeMfx
Mh66P7gV1IePWYun+P1vBcO+lFBmnwp5T1+BvFl/VBzv8evyPDW6UPGuZVaU
61gTrvQF16CQgO52fQb6qxHeslWJPKfnBGw8LRHI+3pH5o7N+n15BkPVfdYF
uAjwoF1XUS6VIB3L9+0i+n1o9iPMMlmoBPsP/JDGJWaYOTzbDvt7zvmwZIb3
QaM3HDUe7wmZxMqfEu0Z42UDfE9oHyuBWe8xhn7Ehj1rU0ZgvnWPp5FLmls/
T8trimNhcoAuqHlUBkgnqmGsGdIYjb/PwD5u3abKNWxbPaWAQgtU0/0zsFRx
eli7+hgZMEe1SCBWZEhPjy0w+iRTFssmN/pO0R84bX5vyft74Nf6gWBnAyGV
PfJioxpF9zCnWdRIHxi5RqVmbbt1/2Oy+4O2SnYbk4aPiayvDktiIXOkGj6l
Qt0PZIUndzMnTGArx6vl3I/ER9f3iEPaXuSkvEvUFuRyJHex+VUI5+tCcux6
cTXf7BHRZRhE2CMgwJIh3p6CNNbTpZURM69yymLkR0FMTh9mniW1OCvcayhr
qm4Ofb9P563R/d4xohpV9/gjRMtqZxFYmzVjmq1Fd7a+1FhyUdgAknjj1xcr
/ejnfSRKeKx49zsXMJYnSFGifdM1AArIGfkm0hN1ceBgxXgFvCbS6vkfMKqY
grfmOJTa0uImC4fBikXQfu5jL8TvBVGQCw7fVPTtSrfr+QeofhaVEK2tDGRD
5FmsLHgMSCOthIhBb66fZIKtHVk7whYQf5GKERr5yPg27e3JuroY6d03Iup9
5avsfZ9dL5IXj6Ei4drGEUCRxUZSSshRvFCPNu6T9kCbeomCTNjbo/qXM0Hp
UVGBgLD+38l96jHTqBlBHOvl9/xvMfzTQkfBjEGBsQabMS6Dfl1svD+y3fkO
/ztkaQQWVs1EKBWr98FoKdHFDHaZWLMjdXQSWKIS7gGSQFqA5UHbRYBRAax7
X1Mdd169FmzfrKwaZjrOh2Tz0oU1U8Asb/T8oxn67twOYsuIjFBrqhBqRwTM
r8BPWwA8a0CA9r7hciNMMTYrOC1OfLQr5YN5BRniAHpJJJNjCNc4iXeuItfJ
anlzDL6stA/iAzYQ3fso3v+9kxMXhXiyga8q1V4EnnyByinEBgpCYweB7nIR
CWNQkvS+VOn9C5bOpa1X099F6+zXagZiAEGl9NbsAeIm2vi8bikGJeF0AMeQ
GGGzivJPd6o8g4caQajP1cNoiLiI9SonoZTOo28zY/0/AXK7IhD//gWX+4dz
BP4Yx96d3qtlXNjSWDKgIkcZEL0pXq+E3/Jx2t+UvUASPjFxrldo0KzcaZN4
UBtGMbGvf3mVcIkFjqN2y3mBzAVyftQUK0ZWKGn4b1BWhGXVSclgUteMgxku
6QZrjB/lULdp/PLQ4p7QDmdqbB7FJYsigahnjmj8XS8/gEqQ50JCn4V/O21s
GoofG1JDARpSfK46GmtVVKuFDUsHHG0Q73Ll4QqhtSwGo3Q+v9OtptNeTNZo
uPNMVqixXRpxJXKyBV7khPoA9b6bwmZF+sRWQKsla2xaWGRoq1Ejm5cC6v/T
HBIreKQNRn/0Hnqn36oZJGKU2k8yL/AZ3NwLX4u7klqfAApSYVBxnArN+8Gw
ckEUmFd9iNsgaJ148hCFASOJD6SUvn8I4c9BhafUBEr9N4pQJJUqwtUsRCYC
IkedA3umRDDq0xIMY8XxkXnmrxS8X5mifjP3gZSjmQrCUqHzNcS6wkyD1s3/
EWKfzFj0X6kpf3LykEPiDVNz8/KhuKJkVFr9946M6TTlfS8G8OxSRF6Qd87y
fbXRTx8WK4R49J4FwE1flIcOb9MerlfDjj3RNxQLOagufVbOpwPbpV/3aFgG
+yVUnY9uPHcHmOxB2/QJgJ7aPuv+I9J0egrnRS8mR90r1cspoZzJJ6EicoYC
CTspWM1uK4gisPSAgibHeP54nLSeje5H76JJicPVHx+oKwqlET2Pyc7AujHj
L5luI1nzmB0H1VdKEoMUaUsDCm1MAJXYiAXTIyMfKVZ4kTAoD4ymvXw0ds8n
vOonQdKo9QdxaZUN4AZnj+M7fjVUjPOiNNwQ4ixcoQg6bjNARU0ByWZAg1rP
E0rOiXaAbNO269zl8tedgXjN58TqQEagRHgdvTJQQyqweSHD8hD0//keC5VB
Tdcy4dL/qcS34+2JdMLgSnBFiQUP0mUaJAEOjqTj1pjOfnKKaeKbEFk5o3Cq
I6iij35KisYp67qTYzhvTpjKSQgEAskf9GqZrzs0fxdtf4HChmE3tJIdu3d2
rCupdrcyOtSlDwkRh4kzH7sBPkMbXLllfpjLQBSQUbacrTN+2vGpvyzwQVNg
PinQ4r8P71Bug+stokqiDbyMiKT/iPHi9Pebff18B5XjjcrjcpYhyeek45kJ
c+YRjZdfv0fl8WO0I5q5llJkqKFTiXECkVIUqZzuVAlj8X+BGZKnC0g6ri0y
E60UqUi+oUzrZOuwr2gYuIWJcsEPpfqqu1M54AHh2KrKkvltqCPpEOqu0Ay/
7VAhGEBihNyIgM3oaH7hb8rT42PBf3Wp2fxFHnaQOeQleJTglG5hU9/BQihf
V2u+5pVH4hNW6+w5I/dFGvQL/jBuCdT/Ih+k/iXdAfY6faV5/K4UPaCToVam
se3mp47Fv9VYecJEJEbdvHaTIPFTIJiar7C+aQI5+kvRlhIX6BxzLoqKsZ98
oBmwwgb47I2RMneUkLFMRlELUdr3KpfXLmZdwJRBsN4n0lR8ykB4/Q+V/cDq
wTQXe/8fDEX0IkQ2WmhUtxwrb40TL/DBpueAL4SYONL6d6FK/Y1ebRKJfjvn
W3jge6PF9GKfoY7bFmXtBAyR+ZHjK2ThsJM4yXs1OLrQF08fUDvQtGipQaCw
Er51UhQ9aW/iHeV8LfA/QxAsLp+UFC97V/AFJeGGiF0vAHevRVBn7Ru4PbOG
Q7DYPK8gQmxDnazGUVKcrGMlFVPS7SzqmPahSQhpW8lfwxPY6Q2uC6bOZOri
YqsLZg1QQ483/Q2Ho7PVZ6cWerKSwBZlrAfIWOiXna9zSZOUj/WNsPHrjd/y
gIiIt0lFTVZkpDxodaAk3bodBYwHCVtzxifRgZ9i+p7yQ83khdz8y4oXP9P1
9CswPk8eDi34qFkEhVtT7eXLkwxGvkmsdm3v2HQsicIDubPTXLK7npm8T8eX
qs9qM+Cr4wAZmAsA24TsleAzMoZnjmNziT2JlRPdop18lwpqJN12il4Ds3gw
RIyUGG7DFLzJwmdqcjl94m0nzMYKLKT1AXyrLDLRPL/TTPIGtVACjGPEmpEs
RYLHB3ZzK4iLLhNmjBCBIUyKH+AblH8SELZ2mWUq2LALuizVTg1a7e1mULjM
Z1mM/z3NnDK6sNzTiNoQBXOjFlCj0/g+YJL82lpg8fXz38HxkVYLuJ3/oF7g
jr5lKB/9PVD4sNx0zVAN1xJflr8o2S1ZQvx5YwW/behuIQjs4bWP0b55U2FY
Z8jCDGjMsheLfCVYT4+Kb+f1X9URl9T5FizGDSUjahuK2CF+zlkgI1Hzlhfa
htOy9iLU8ISj/triyP3iWiTSXUZxy+rQB2eXOxok+t+tZbzYx+TP2TB8lJM0
rptutEbjRmmMCfkbF/lsWMFDc48LuPLRekWHnUUD3I0p3K/slN6X0a9R4mOv
Daz1HNNSk9p8FRDx5DCOtUOeR7+I62B28W5GeTY8WYtSkUgRkDVjFWypHzkv
QoEksGqoGAj0DP7/BfmreTZUTx80JrIhV/UHsycSB6VLUv8Z6TXErDv+sbTk
K7RFUmyJZxkQuGLb1l4Q6FgK/l+gqaNMT5Rx0xZQUJvxyK7DQMqz12gefN/B
J63iBTX13Ck46CyEe5kLJ6ArXsmp7lCxviHqQpPymIe59bPN8oVQornyQ4Sz
36UxTweeXC6uhCNFbs4JlQv+TkMpA1hFv2c6q+Mfbz+3zLLnzy/FDNlpa7xb
k0l7gPVt3tls2u48KnsPKgnfTfFtiqgylSbGQ8Ohp94K9tEQmaQODWgBCcJp
Ak/GGdxNtAVYO1x2QApJhB+LoNH07y8cTgO6wVVIowF4bNtpRTBvCr64daKG
usmEVwrFzl9A3d+kmqW0F15KmC8M0gML807u6mwXMI/meL3ivntyrAHheIkv
WhG7iEAHaMCpPDy9pvKoJh4/BEnZoGg2ryN70ijD8gQjcwA7PpY7DCAz8657
wWg7dpNgmQul4h3oV0R4agRTdBTgI/ALDt35URMSF3LdsZRmLCh2HKIoSv/1
Q+Fl1EYrgMvLtNMDOW3JuFNviWHmkphUnsNQ83mzmTMQRdHT+4quRh/msql1
voG1B9FHTAmbf9bJC8+DT1G1W8duAydYm8wiHxV3/vrHwVw9OD2ezmQ6FUI1
BVs0bBm5nJXGI8e0kO4X/m4RdCeODjOquedDOfQUiNE+4FKxRB6yffaSER4B
Kbys3A7KBES5yjaP1wfGPKyiMUuCVGgsNr1O+YjtyPxWKokDq0nifjzb30Ix
ixx/nn043g900MxZMGoiEH2I5ZQTKC4YJHUuLChYXJlCin2iFhU+eAFBsbxF
hmMcfOawCegFVm18Dm2/ctGO1PWgBSVJvnUSO94hxDX2PaQZFBZT7XzCNZTQ
OtnHBq9l56o9VRbtDTM/NvOHPccxfFGEQPU40QPbWQDRytxZncxMUWt9F7OF
u/GQysOww/u8JtrM78HlZd+3NjzK/0wP2NL2rTZvlf6BdNlnvVUuDbpKXMv2
5eLBGTJPApxPmo0dLcxz8AFVi1cXUaUkkzCdNojk+nKHwCOhffJjeHUtN/uZ
a1qebjZseLxKfXEon8yBvRUyPQFDtolFgUOVNlgByUCSsp4VaRHbx3qcTMY2
/Q27duzYrP/swBy+U6a06L9Ca/DmiCBFl3veK2+kX7sx3LiN2o2Ush5rOrIi
WK1fNyO+5voBB7WIRikUNqdLU1L9cfu0if6n8/uTZl1nmKLKdcV22f7lhxBu
+goe1cQ4UV1+L0D7SVLKOT0dFcaSsCR86KfYMn+692Ecu3AEvq0rFR16uB/A
IMRlyDn6UNXxSFFkuCIW3fSD/h8L19ifwQ1sKEOAkDLDldZIR+7Cw4W1TRdp
1r+5DeqYbxhmRiNbG+FXk+rwajaEru+fpdEOXugV1qHRc3WkDCoSjsa82VP3
yMC5sYCvPOMAQdXgx0T33xuqMP7Qiigefm9Ww5hqAz54Yh0oG/Lqra2BP0fV
rKQTcq2kSpmDE5eM687dDtXFplmP3Su5fB01VVseeTZWu0lTeWqHDdcnEfVx
LZaRfHI+ZCwymQdHargd5s7lYc6pkQc6IKETfKcBVET3dwvVfFZ969mVJGHq
uFLD3dygDy3hr1eb3Q+aC1wSgIrlkp0zIrOBIIFFzbE2BMvcgQ0r7H/jcFWH
zGhth3S4b16T4/zsvjEix6N6PZqcOBVeihBUY2ZK/7jllbuAC89J63yIWcoI
cMw+lhJRzkaCWv4gcuYrijuVfR24KgFDNfs8NXDcRY6PhmUdu/VYjNs5fMjY
iVLJa8v9A6mLjbV2P8uUN0AGLgg1DhkfCiwp58HbrrcKNoXQrbp5WUr3BtT2
PO8grSizlLSuM9DlsgjSkDzReDawA3oOkpD38aiaEVSalLa92G/Yuj91dPUr
6hhzx2OtaEvsuLTQQLeAdJJJjMhx7ttYaUSiraO+rVZCFv4aI2xYAyGtVkQ+
jIJnA8xUGw8zcfsPUyzJP4hf/SOZJqSQvIkKVH/C1RwbsId72Ii55diSIyMd
4W+UAxtSuP/xV9ErOZlHVT1if0x/j56r1ZIxn6mEZntaNhbYNYeVUMnTfqaD
7kFwhOjiZzo6pmqdfAGGoeT0TeT5S2gF5/A0HmrXti5+mRdj8X8JhyRijcr2
/xVbjUkpQzNVMZN7Q+CGAL1ot7Ev2A7yx+ZWpiRIZdEWq0VcT8B7VBijxdm8
277Y9yrsP/f/EMoTEFLP3my39QA0I8yePDAKzseOukcm1/8hJRiNAnakgRt/
3oH5VqIbA0ClKmzzK14Coy7ivn47GftPgrFXFxi4aJZV7m3aDmawnxlfDmpm
wfcLVW9zq27cpWxUrw3hPct1gJLkXiGIdnPScBKpZ+TwgHIg1JbfoNRxv6e0
rryvoQSFnQmYO4pir3ZqkVo3MKU5GwvMjYkrafmfLCmgs9B+ioAjO3vwgdLK
nityZqp4eHpEriiTNea/dqo3QXQnmhk6mW6dPtKe1sroLiEiyoKKQ7OWIyyR
g1jLuf+qY5cC5WUlB8HqVxx8ovnLsc4az7rbaFl1kqsBk+rNOMLvM+oZteXn
hzfVxcgqovrSrm4KKRAPIV9cULhyKe/NPtmPIMn1MskSo89Cy3jvDuGp8rg3
dlPwi989hnNzqHS9m2zL/eyG0zaKzTfETBlG5kcw8JNlmM6s2SRoz1sXruat
Ju1XkJ0YvGN34Kdgqjj3mVm/1WOPOgGOj0lHhAaKTCRLipRHwrraEkshAEuJ
8pgr/RcVGn4SypFzL/GkVR3v0nPbsJDsgZ7HRGHFQhqYknaNVoRidG8Lxl6i
Opd+wWmU8A7ExASRrbGpyBQESm1QXsDMoMdgdJWRpTvc0wjKHq+V4Q6vr9Lp
p43hYOhk3OIcwV7BvuXYj7JeD08cR8kukGvRFnm5j1o30xypDze8M7kNl8jo
P8vqsNOQaZkpWKG1a/ijVdQ73vsb/n+BD7+JCI9hSws61rUAviExqX3nbf9D
0MBWQp5aPfcLhPRENscFYnldzzJz9xTkAtlsb2vVLUUilRe39/x9eeNr05YK
2+OBTCUEo4D61xUNi9yxp/grc8mwhFmXkkN7bLEr/OdrXkd7KMJCNietma1S
jPH+R0GHnihDpiTjoPnIyllGY5V5x+So8OmFrdaJWFVxxf88eiRybwsEbkH7
u1IIlUt3JIFsjkcyKTz4E/c2hUuXZFnb8MgZFlFvj6EO/tALRuJfi6/4aB41
JLfC6xyqcHZ71ip4aLwCWUAKaZoVUkwyv0U2FaUnhbzW3MWBZLvQlEOBNlIZ
HDwpcIe2Op9VbpZQioMvT46uPQTwQiUpZYfGtuAis2AWbA/uGpwzcUl2ueLF
41efYJWB3uTv9C5CN8wCiGPKh6GAizojTPWoYqanqOQxf2EJbKLaY0sEj2wB
aA73z2SeqXxFGjEB2ZcQED3DMO7t+c+cKfGIcMtB/2Rjz0LGuXtaSqzUMQ09
E14Zqh98XuAlckB8Uc3K8RFk1s/+mTSulI/+0aUP26KCaguH9lInEs+2CtBc
6gQ/BfefnI/o9zwvBu1l43bn2/LJeiGYan91f+gR3GkqDeGRIiihrRXgV9V5
6x38F8EGN0n5izvRuAvfYrF/rpi6HEoOPHIr28XiAwYON68P9XxqvraBfj7B
tzWRq+Sq7PtaImawtURO8HnWxBG7bIHdmcQLK5xSMb0/psLqxlTvyUdV5TxU
e4KZ+GlnWlsoGpNFdmhFVRhnD8XL5H1SWim0VdIXRVK6vuuw+N1DZm6DUuTb
Ed8wxEG6ACb+lbfdbL6VKcLoqbfsTEl0JqlTitxE0p2Vv6fHjFYmhzuTiZKb
6EQjtv/62h/EhN1AnTPExaXByrPb7PEcx2DAWgUy8T2SSmNlb79HXtHo0KKO
dkemHpckF5QUmllUwn6r10a2zMSjo2nXppmC4yJsmexKEvIXHVMmGeXZ86a4
osJCGtFk2Ow7JI9jg1V3xqFoLd1qzPq3Da5/vSKe6amoKLQ3bzoceomkxOYW
65JlxG4s/KdIBPl3Q+kaGYQQD0HdF93yYPi6UnhzAxuhWBySdpZD3qQ6Tx72
cTg09UBX0+/Sq54u+N0kXW91albVQuaRs8bM1zekNHpiJkcin+IffUYIPdNt
0cx/BvHh+bg7dDBwCbeIpM6R76t4GPYHK3rXTaAi84+cbrOxwN+WgnWwNRBv
WGsXOMNTQZoMRqWqU/DbHJZU7ZSsGzGdroNBiCCpIHD1U1zeDvt3Sv1qCd/v
H9PsXeqKNqhIS8SL6kgGqZKX08lQHYaNiGkWVXS6Ht2RbdRlwO+4gNkqT1S7
OZoyR99tTyPUVOi96M2sSFMaEP+6+vjp59czedm6eidck+vmhPn9+oNl8m6O
PJeBb5A4flxE4CW1NJSdMY7EBydsEawanuV01rGgkL/vkw32YUPX8I78DPag
RxMRyhHW83k/Kd1622tLFYk7ZEoeKFptJMK5a+c91v6EY0aLfqwPLxjEzsrw
sgIwFRygnLV8YRlL3aLZ/tgYgwluj8WFPPMVm6FPEv7hZVfAXlikuaG1OJYU
N0b8yOi5n2CZ671G64yzaYsMTwXlNPiqMkaJmk6B/BSGIrKJDjMBjSt/pp4x
NKvF2svrEs/U66z2OulzxoJnro75eCCWlLqCPOg2hkouvMuoBGzMN4cb7Is1
EikYVG2X0d0QZgg++2OaRVRfOb9bNMI03dpLZixcfNT8QQCoMzKPd/lPsbqT
7wMCVmulUeiSTHAr/MI+IjuNUpre4Npgsi+PHClAkeK7DSsuEMQrkDbBWjyO
uLiaGf+b2riUuGpTLTWwSx71pd7IsmaLx3V9rTZEbUhFWGu8WD/m4WKMK6wV
vJWPPL2dMd+LzY40osOdI/CuQPMbj8s+QYq8LeKoRQXpC2fuMlALxKAucE7G
oK/DnZ2LJ2u4fsKh5DNODfzDXmixOpYSWrqBCocIMnfdEwT1bI1JPmpYFq+p
TpYpXXKEsiKuGIvSAtsrZAY6vW578zEi0V4syQe0Zlus10e/psXzE/YVPLxv
7hhNEoD4cuEg+AGh2hqF+aG+5GX5hTdy7E4PUbRNwBOOlAJe4NJ3p/nuZsMC
SFvWhxux6NGZTvjDZtxVrtdCDPYtvmkCyiOGlgPju8kGoOHmz60QfN/hUY+T
5ii6Ku4tJ52PrQjjykTb/bodMqLsUyNha7w/dV9i6+EMOzn1FNjZL+oipfzb
MtP24jjiIfRa4okkvKGd3LvWKr+npBCdi0oN+7XWfdzdNj5V1AJnpEBQRrMl
pY9yCcFm+lbrOQrXlXFc7BnNH3dlJQAmzlmFMGMuVjIyKGQxwLK/0k2V5ri6
3IhQONvH9eIzdXb+1tSVIMLe8tirHgq8OBfU3gsv9ldhhni8+F2smxgLz2ma
2s7RxkSO3AKEdBmcXaNdq9TiHCID5plq3zSOJO1A5nprlhVYvhIjIL9kaXqG
t4aaTrlf3nrMYgUqWxvGvc+/fEFH4AlzLshIjs5qm7ohzMiAL2APHHD7D3ri
2FzNol9+N29ZVzIcB2Az4o1EKVBlvLallpKm5iF3XVai6tliW5iaisiWfVAH
n/Rfef68R9GrWBam7iCbW4HUahysAEq0bQ1jRj2moRbgdd9P/jMJYrQ6kRu9
Y01KvuowU7iFn83KWYX5QkoSSDHgR0e/RKMYn/JshcQLDVMRcDPnnapW/cD1
Cp2p6rejUms440jeFErJsfkOD0bYkKJZJdNeKZzKGwZkmbXVMTWdWRU5t93n
rrw5jPNVsDhA8aZKEjUFoUlGVdoEiUyMjaQeF8UC5msIGSb2D+ioL4dK38gf
QsfYwXTFgXBdZHrmt4fEk2ZIc/pG/qXy5cG5xfv5dLl6u55Q6aVKeCKvZVzz
yveZi1dzz6Zz6sBOXT9v4WFoJBPXGqqboaON3WHxY3wIBcGCEM8S8RHnNzN4
RwuRHoi+FHOppUjQV1l20RlX9v7/ElcXSicZMiYEfxlbH+oZ8WlSozfi+E7e
hPboJqJDSnGWLrsoGlU1EKU222Owu5j2XUW3czpuebY47iIW/B+k4owUApOj
qVr1mokzCl+AQvk+1Cvw7P3XG6zAlXL6YfAaFpFS+dNUH/wlVuSze6kTkcBz
/vgsXfSLFx0m3WFKRZKO+K6+D+5UNpmp3xx5P7Asli7xcbijlV0TAoeDiYWz
Dpwg9QLEzncZNxT9qZdRFZBwawF5SOzZuJO3DVds1nSXMpUgQfeO+ieEixxf
3xr1jd7TqDpt+RuPLlKJJ3OZkYoV38XUX/EHeqjKlbDe6NR18yMHEpegaKTn
I6hvKol9LK/ie+BRQYi6unaVZ+3b8ScaL4JN9e6VI9cmCM09UUYwIMCoy9J1
VcfjXn06HOWme+39MtBdeiWA9HFOqokAKmPW1yoAwlnbeOZeNqzhafYLIS+l
m+Y9804pxF/1/HUOAqmjaMV95K9Zez+oN0WeOYc05BLEKJjhz1wAbye+nuQ9
PBymk3dt+g6CIaH0SQhFO3VWljqRzOIZSuHmIpSWOOwPw0VHxxD2BfSZEgWt
YiDweoDhbTxKbMxa7C45v6tZeVzDeJgEdCoxPt7avfJyyQqRZMlNdKSPe5Ko
LaSMGF6mMFgUwotIykdlrZyMFxzVPsAbLQ4+X11IsZFy6flDQg39cJwSYLgp
hez+cN7ndgwpA3ySWOJmdX4m7YO4TE2QY4Lr180EB3O4aWqkgq1XF9A6QaoC
FLUIr32KoJVDsWUxqiGWgl66XZpeQm1+ygNhIx6x2k5KxuRJF/bnjRREIBgM
rpXzBxgEHiDy7D0YiqD9S/mdgthrOSEVI2ejB/cZDOptV/hK3NWG9PuZKAmW
ZzCLg4JrvFcu7kvbMYm++xkrJEveGKXbORfF2aDW/CWO/ot0DVz6yc5KOfBN
NIbMmqCzoEqUr9tutppP//sMWhzDg8KxQtzuMKDG0wzzuNqSWXRw9AgIlEYU
U9logD8WemUvMVqpbVg8CZg1PcvS/YyDJmwcB5SE9LTKpffygvMTeUjxX3Zh
wu3qcpNxoayQffBQ55C4pd/MXz+YOGGB1A0Buiwz5NHYK1LuR+2YHxyhODDf
ufl0g7c8r2QVCqYSo6AxcukUi67Ik/Ld3isEMLBk3SIWuMeo/DibC5BO12eA
zVDJUoGCgdYzyU6ojdKUGov25uRkDjGUY+4E35e49cIB2F0SFlNZUB283tkd
eI/yKvo00zBwuBVYdt0/UFvEecbeIWQI2ouWrHtsLABiPxF5WStqthQQUSEj
2n1rM/kf968nmOQT0Tj5q5zGD194TChOQsnQgGh7faj/mN89a0mGtLlp03Gw
aU0+MVhiWWcekDszgp3aUM8vSPVx7Og8nH+dEPIs3PgwUdgAT8gTEitJzPaK
I4xstmza6jbbpzCM7xAWzCmCcAG6yZIr3gDGajKJIbxyQsF50Pt1dM7sEsK9
bf/ZpRydfluY5k3exN6A3xbBRQsp2+Um9E1xqiy4tG/+BxKG1wYNp9di2rnL
y9NbNixV9JJnhhOL6gWAndqqSyvbeKmi6e7Xha8dlZTT3+3YBs+215omCX7R
eCJ3tDQqlxYkzfks/n2pnU0I73SvSAL9NEkCl9oH3ISdQ/moAByfdcxTNE3Q
YH+f7MhpPuuuVZD67RY0M8RJwW6rlkH5aXDRBaXbQ2sJb8KmwjIrJjAIMvk6
96+70lWgVUSLvGh6Sbsrc6cANKz4qhvuLqqpda3mTIA5MfwvvQZETibjo345
DrSjusC2rcsDCktGfGzhA3MqypPvjGJnTdDQie3howSexr07AEIlJsE9g5hH
ebwe6vWfhKHBcotSsPgudEp/w/AvM2jdx3dJFSRe4gzz7SyTMCOxTvANjBgO
PMVQD/I2qtBsViv+YCmQs0/tIi38uTAOiYobMobvh20+J/aqUY7l2PbjA/mA
1NkFlnwtzYAMMeqaIGlEiH8Ebd/warvBWaE+hMRl7KmjzQG73M0mKf1gSmTv
wLxZlnm23gGbNpEgCa43FTSxllBxrAETFaZwQfRJEA+jyksDoDcybEUmrQNw
mErCz5Ohg9O4h1E7jEQlvqHfGanG7ofNqIBo/7dbNxXgRElXe4S+5fJm8USW
kPCylHQDxfDX6Br1f4Iy6yvAM2sKOO/GsqdHJXTW2WujecD/Tfrahx2jpYCa
MUxZS7X7MHMKwwpgaM6eEAuqgaRfbXlO3nLVeHrKh4AAH831KIvQa40ny4bW
GIlQWWDpkofZoxIHxU+iV7qrwcJB1Xp1Zj3ZWr0zY3G3dfPQlZAmS+isTLCQ
k2wqqCzSIde3fI8+GiNfeTt4wfm3I3RPHVwK2kR1//aLql5Ss6c8AeChE43o
cAi4gzk4BE7EX3iTGQ+Y5HVe5VMX+ie0MZQThhqchF8DhWqPwXWq46Y3e8ft
q1ssAKVyZ2wb3B/SmXJ8yxDLTAmW3PDWUV2N0C4eyMYtX8ZRQ8f4o6nJtTzQ
NQ5WynWf+ljGQdfgpxwXC5dXGFQ0GgP4V1/B7H7TmM05MwG+2NWkAUhnqXcP
5bAmd5Hfb7/UMT6kwbYo+wpQfZx27PMovYQvEiG2BUmzrHoSIKGkd4wluiGz
Fp/JRa1GcZb0pVDHuKml2JrXyYDMo57Yph3g4XBCmVgZODMU6TNTkfVfOQLd
hmOJIeiljMKkRYKML/0K6+FAID7huTy3kJi7L5NB8ufHYdmCWwOrM1fOqVIk
VtMQ9GhYcCowLOvzG7KmM6b23gVOrCvkK4jF5f3rlwP8s2EmlwbDzOmhZLEx
vbffvyKsGrMAnmZS09qx50bwM0K46uQLI4gJvqKTRQqMqYL/dmuDwrwOKBNC
kAIIDZXhmMkGK5hEO8MDyijK8IAVvCj/i+FxEvmAzHPROyjsYin3V3hKQRie
njGSJ3k7axVP6D3KEMNLFmWKHgjvA5qAvtd564DbAZP9BhjQNlJPq47CTKNd
y78V1Oz/7uTxT7Di9xOfcI0ss/XPm4dyICvVeX5oW2M+/wwoZti1GlS2YTyE
kuCHLxsiGcMC9KHCi31wX+6wIrXMYDf/A6ATbjRUUW8OkIZye0H7Cymwp/Ds
nOtyrI7mJ3iITfAAWCuJKdE9sq6eHG35HM7L0IPm6fw18ugYoGOaFPf9spwN
RakkdULV7vxTgMr80PROKoYB3o1s7B/bEQJitxYDtlOvSMti4PIXHqVzocMd
Qv54TUBk9LX730lQ4GXQgO3AKI/FAHJkG1myOBqqAsbje30b+P/RCdqRc25c
hBiyt4zq+Xqd6EPDV9AM1gpMKqO3Zp2YPmbMMjFX0LKjGJbKabH/xTaRw0mq
UKVxVLaPe+uL0INKT6GlcABoUdqAr+UI2ciMuinbyCyuaYn8BrwGOGHPAtW6
jMst2vKBIXbeF/oHhS/h6SOfT94uxOeaJzGE/XC3UIanM+kIIYohHDV79ufO
yLgqrrz83mBo9Q38Fu5ajigQIlqmx3g9EYlFbxrgRflEjX8JfMlZzK2nfG+/
11cd5dngBtnxmJ8M8AoqJhHUSDdM75GWYeWZZFrN9Kr9b1Yn7Hrnxy/xe1sc
YXQa/zJ+5SrYFkINX/0j3R//0GQ+U9Uhg2a1GsGHGeC0BrntFqapFf6uckFk
XPgRTWfw8wZkj5WANpOJSC14iGYeDb8sBWX7KZsF6yrkp/qsQItskrnlv3ZL
Lj6ZtPLj1jHVtiA4NVINkUjE8zSSDfz6T+BmRjsuubLoUHQyxTG6WBbsgmMH
80AuOmN8nB+y9xBDnt767rEwiRKUd1nG4lfIyCEP62MRSGHDtUZSNrEJdVHK
9Y9F0U02FFPWG2bb01wnc/LOkQCMcUoWALEcMPvDWDZ6WS/J8Z7+S59vFcjl
aBgzIpG3TcQmHISJK5zpAebiVfsD0z0GI1zOqPBY7M2Ak7gJNnELutAo5Wlu
fOuqzPqsKSWKnthu1KXWwY7JsdQrStoDEykSUp8amWxkdbLQTbOughyna3Am
T0eBr1OpQyePmv1lyfmqtP/kYoGHnbjE5FGPViop76I1N2Fvpz7IcRtC+jr2
i9B6cFJZVXYTVVVtMm67ZZLSyzyIytKKOKlKX9klfKpMGCiyCBbuxaG3EdV9
r4jaICdaiE5rICxcaBUk7NSsnyPBZQJNZ5W/Eq8ZNmwv4x50zrM+J763UmGa
XBdKnthq0cYFPypQi/TuSaI+s0uhaajh6r8tFOB1CPzpY5OBdn0bLzsNXLDo
mh8fw0earcbD0z1Akaif/OQez77hQLp/U1FWkkGjYQg0aPMYSHklszAEmHKM
ervHFvb0C6vIVMMG8G5woKNJ+N5qXUqGi5yVygc5yVI/xsVsYuDjKbcZFecW
lNtU4WYiA8bskO6iuw2EIT2W9Lv4/1aRjhGquF1O9xpdWi9/JVdxqEvgb0mP
cea7n6gdFMIBlAEB4pyY5AqF30tzflYUADng+kPLiM/u6daTveYGWgDFBaT2
rtZHo/nprC70ujMuYt7KEZt/3n07gub3jtyOQ/GeQ9SVzMSRb5z8BNhluFwX
Z74yqAch9vXfAgSp8faETDz4dtBXvOPkR+NIwRAmI5KLJgtmsq7Rl6LurayH
pOOAINTn8FaZNjEANj5zP6snuwNN6mEadTxFG+eZzgvPPluLnOyCAjKEFHsy
yaSRm3KQOjJiWhCTPgZ34dJ3wQrn653v6DPlT0IQZJOarxetbHHgIzlRJJya
r1W7LGeFh8E8Zx3egNlFB5ZYD5Oz4IG1h0h00YC1Y5BR7OWMSgadwvXxmQFz
PvhsM/NuY/oB5H9hcI+chlOAEgOe1mvpD5Rhzi8AnfJmJxQYearUkSTXOdXY
RTUOUsHCi1EVGI6a0EnoFAJWatWs+AnmYkBbrrjSJPP9Lk7f/s+VR01CVXS/
hDl5V0A1qGsknY5vlwHd7roIdlOLfKf2AiYc902CTHaRdFLTdAtkEQSvAwhw
oMmFkZ3MeBWhZsl7ZehGyUybRs3YqERg8K3MJq7Ynqq8F5WrdoAyIXT2AxYV
qz1nA3C5sq26Y8lZ8HKVh4pIm6r8+Z4W2S6+qpuo238mOPossF2Avcp4Gn9A
uORJLEO3VkvnVEHWkd3gnf6Mp5gELwhU/Y/KqiTr5m3+1+JEsaQ9VU5vKHND
UvFBGc2FSjt/ahSbI6YWVJQg7NPamFGJ/MFNwiR0ce7YlxJGhZkZM5VSVINv
Fw4b31c1lQ2DwbFPhJepz4x4ZC1hUH6NzX1Yyu8P4sGoTNBNFeJ8kSJfn8A1
knbVtvliUQm6cfWYTodUgYrEB3x8oI9rDLsqSeXXnuwZpnC5b00qddK+M+ZC
K0XMvOP6R7qEbqaKbPlY38j6JVBSFNk0S7JJDtjTshwP91ENGlgqif5VBXmK
6tbdsZexg5l1CfvO8yv5vqQE7RFNIxAeGeyD9wH2QMceLRBhz8iMfURZV9XI
ie37X1+7RzRx4J+ww2Bnjf2YX1+eZuJ9KM3UWdhKuUJOA37pNrlpXf9y2gp1
L+2YVZ2ShVlWIr8sRgkIpRqqHKxxkbsnW7Rvx/S00iXUhHGBdrYLc/CY/XQh
Dr4sCJaGy1j2Ac87LXg6uPBgRty8hozsJEkgv7J89TbzTSmj0OoDNIfFANyW
vbOt2yqNYVy5WpN7VwnN0Jjz96RKveBb134d8kpEBkDBJvZ2UEPIjCqR4GOF
BkZn1SnhaJ/olCxGEzwFOobStkuH2oIOLzm1HzF8UAXtb+0Z634VOP8YnRRh
t56NCZAKDQMBwb6LLakiV3i5zq0QBlUF/lOX0ivl64aEoIUfK5lcl0CeA87f
yxIBD4tIRO02lw9MyMCtxhBwUhNXktzGOmVBfQ8HaTWqU/OGWaV1VpAFroyz
4quYOzLzDY0mB6w03ebxzr1Cu/WOMvQm9eCMOFHYgqfNQb/eyXS2+yu5rFrx
TjjNDy0ztHSHBQUMEMU6cS0nCVukPHchk4ixfq83+5W5wXZ47XW/BlSmrCxM
H0AMDnH7R4Bik2+h017VfOeS6SOWGq8+a0xL+zFsrVSpov0JFxg62BB3vvBx
fcfSd6I2lU2A6cr+XyAEmzZXZkTaFh7uFuG9OsUKSy+7nKhACWTj4gzp7EAB
53ANzHG9NaOIoZHdxzPD351/3fS0Y284Y7ggYhqY6Uf/INOicpT4QdvZ/9ae
AndRHQcLyqMu/bxkuN1ZWXngvy3+VieUJxfMVpYUcdh0Q6a/ixaIC1iPZz9Y
XA7L46dPVAiLTU7T33hKpVjV0D59Ch5S60MfWY6DVQOF/ZFtccpm2w1xluwm
TkOff8NC2IkQmWcsx+F1MoA1gpDvPG9Q6zBPT/oaOdzHEyyg6FDcEt3MuigK
N5rPLqpkRyKSSAv35b72GSTr2UFRdmitAJISXbfsNUUnhgQrmzjIA2gm2OW7
Hh391hVDRO4cJX9ydWRyWdVwVC7BqgZ/s+BhycHTa3IsI1l+jiQEABrQ6KfB
Ums02Zb/21zL0zSzmVEO1a5cVm2ZBgF1BAYokK0uaMRprfUPJj6Z4vaEx63V
5uQMddzzbsEynYDRdsTnpn/y4s9Pfy8lXMpMtDY/KhBLKWuglrN3SkW2qRUG
9Jzt8NbDC/dZEJNW+xIYt1pc6bf/1kagRrhBQFg0olLuzfZC4aP9QWza6za8
o8gY7zapccH8E+vR3A5+G0eBYCQ6DuIFeMTrkzLqzM7+PbRW4eny9x1gu7NX
3c7wSCQ7wgnHVJjNX7/xDbH0OzHb3kPvvBlPqGuJ6AEYZMAgvFKwRCED7OGH
9HI0fAgw8tz6Dxi4Ro9jpa5fLt3hdRWUmgrFlDpKWSw640svyAnJQ2liqNpa
NLAnUbiRZQFESt8Z0Ox4WUyKes8wK3JUVV12ElEqwvduSdQMyFAj805N2ZRX
b2KQOVCXfDhpV1cJx/WoRvxXPKDZa7/gLdD/jtYWHettdibYpgvNO4mpwzpj
NTIOBivsG5WUmVG/RrNDPwhmGyW9hFI7hOPC4m6aSbK9XRt1Ri2AsadcClFS
XbzDgD7z2Lbf+3qUp6dGWu1BSfrddz3Vpp00e0gjkaff/X2iOxeKtM5UxJWX
S/015w2BxwtOKSZSY53cVbga5G8GmiL9vQj6J5+OQHmXgG4KghvfoJTiluJ8
T3V7cqtOj8rVoY3eoZ6/WBB9kNgBDz0qggK4SyjRk8RQJGKU7uR1Ds5a6JbX
BMhyabuCpc71yOcQvaslyPfi8Ev8Od7eX5H/S2TXQDEF59A5CNm88h57ZtYc
wRU2GfkauLK4FfvCwjyCY43Bbmx0WnuyDGk+NcTbZ4eTbEsoJGvZ7867w+eE
Go58iKaVDFYlSau73VAtgsrYGoQP4JTDqUe8dc792o7b0zcyLQVkXLY477bT
+9+gr5FLB14ozfMDGZKv/Ik50C464VHt9hA5+/K8wFF64xTkNtqVHWgzUL67
l0ZrlV+1rpDuqPH7jPTaqP7wM1T/9o4vacw8Vapn6ZfxDZTgkX2d3n4Q53hi
uudFDWItuF6yf1WytESpo2J3VYsa+dN8BMEDoGHUvscwmcrhRuti+lRhH9/u
cs/Zt3fkP4cBpqQEsBFhMC47x2uzsPgUv5Qvl3sOXYkKK3bNQFDOn2/qVqTO
0x98DstB2GDb/TSXHbyq997zS1EWMkBAdWj3LRFcyj56/wCVnVSwzXgTGTlW
cUwBHf6c5b86YfbxuSeJQzWR5NHbWAQVqgRIvhEcPxaU9VCnVpOlDcVFU70q
PkBkKXX1vNaretzJOfPvsG9ILiKoEH0XxkCauz9IFpFVxdDDn5W7tpbl5xey
DKW5x51G7aactM9yhGy6nCQ3jIxtjQcz8QzWJ1vgWnFvV+WEB9ZYuf//pjuN
kLe665mNMHwxEKW3IcaoQnvtkeb+uqTMRGEqYuyNYF73w8mXuZO/cUtcw6nR
KqmUSytOWOYiuR3yOlSbVWKf4vTbdE8J+4ab8O8ZssWCQ5mD+w4NvFrVDivW
ddF31qGk8hXor5cUXqQCUv3ChQ3glhI9EkulSmoaTjsda9RxmzIv3mf2LE/6
DNWH5U8VlvsJXVt/N2tVtsMxrjFidpEfvo7Te6v+m/E1yf7RFfUgCC9uovfU
gpLzEHeofGFObtyeTSmzRyAgs7PE0sn7YMcaaPC1n1bM9KQLU2jmMdlgIsgx
I5wU1ksZaIaGpPwH6rWSFramU7Q9HPXoE8xXsU7JTpkTj3jw4U1Huxu6pen/
PF51U7WQzzas379y/g2/thJENUnh+kQUiyyBYWEld20uG9nK32XrRO9ru3Ti
tvIsnpOHgss9Kx/kisf7Ad8p7aTwWHCozB33deP1XTu4mm8Vp6datlA5cWIV
Hw2XOhioZY6WljFo69Lxx1HKi22InlimhLSoZqtbpI3NDClfWQXecN41DwjU
Dk6tXm4ZSfA3Jpit+CAs2WHfwKBylvDlz/H3lb+WrchAVThwCMiOklTKdrD/
VJiPuLf+gabVQqW9vs2tMJ5Tz3bvaUhdnYfEiqoUTtgqPiT7EJM36mDrDfLO
QFOQ6xRkz/73Bexlay3Uj9isYgNyytF4M0mQrBExVIv5E57gBOdJoslj+3P9
WfqIvumjG//1yoCRG07xmgGyBcUSc1e4epqAWgZz41khaqdxpIqRE4cneyAr
ixc7c///ZrUKm9PDw+NP4Q3L/3LCAT3F7WffwU32Etz0CxPSpTFnNPgVkBCO
GTdraz0D0lbd/J+x2FM0fOSbYA9WtPQCP2BkFR6iFYqjlDbrrRymza6BeQuN
r7lYaG3Uy1Ve5/tkotCMjXPzoBWdtiGLMkZs3WbgHLhGhg9tJx7pc7b/leDZ
zH4FYMPhhbppvQqHAaPTppKDg24E6uuanTyWkOoyeefMBrOA0uU3M0xSDABM
NJgg3DHE6jxGvsJZn1vr6WsZmePthzKEMhFplX46ntqNe6f03tNgqDY3tuo/
MVvYorSlCcZ7ZcXcwQaIem5MEeoZJfnncYbvkFzvR478nRauXz4KxQjPv78a
A9gxNhNiatIyKYb8AAsCf78c6UG6LhN88A9NK3H33+CXyyHwVrU3IR28zd3N
8GoUwCRzTrwQg+ZyalxxxgjyadNgEEfTDw7TRxMLbVLCPG0EHDeQz8Jqbrci
oYHLO6JQnBeCxQyo/flLrQPlB2Yn59pWxcYdmnN60ybh0sc2T58DTSZtBhgj
PvUrHB1IN7NIR5D1k7LU1eAP+QgLs3IS0CEv6GgVTOqC/DksvM7lSHhAQuA/
SJXKd5rOpXkBJq1URIpDo7MlcYuMl+Fi2CRJ25GuF7xZHXSrD2c5hIP3UBFN
fyJYlaS/cclSuesoxffME1tKtxNUO3k/D5EqAgRA1gpJhYVdeONec2sF/6pj
laSMpQIkERj/9uaLo1ZahbE2IfuiHVXmrqwcFEZBRev4bc5TDOjU4XD0/vmT
yVc4gWsHQ0tDyvW0OfUUPFnlyrUQmAlGFyN2yC07mT1Q4BiNwxnQ+iH5M7aG
pfWzGkvxfCj1FVdzIIZ0LJSnLsIiJBdmw9rkmJr0fqoMOJ17HDw+0QSlt7ro
mdH6okPZOCxynKxIYKA4Wndx5Gzgi81ElT+cRBoccPtmX+pqdpZZTAoiZI61
2p4T57e96xZJ1lnTAebrTaJ3y2nFk0xvIUwELyGDaci/2jqNkHqixCe2FgGK
lNGYrL225nIzMjpWgd+KDRF3MNah3XfGtekjVoVR28Sa/OU33fTPfH0+uj24
pLkzEvyLRayY8DjnaE6gtJsi0UcV81e6ZRUfNiT24En2roQf1RsAYCALxcLy
R5SC0tMyo9xCvSWki8Y5msm/UsBPb1+/5+zT6TbMp27hhhsVT7++O/7q8jM8
ewcHOzklchBbWJjfE7IwXOEjwpVKXy6QXSpcDiRFP7RHZP/iuojYqWnUe/LI
jIf7r0xLhyxlzHamuilsbsxzIO5AG0R0n0XYNSqDnEKsb/WWGyiaGj5FFRxP
U1RESHuXEhjWo3STo6pYtl6jQgGFdyPppZsgnTQves8OBcLzskVYe6VwwDIc
WkAGGWZulyMa8E4/gqEIm+gTOyiVPQufQH5iT5yj8Hp1l9bC1o7oGywnCh4A
M/Wr2WdlYkSMts9AK3ujxyFKhgXUxHL/xsEHEGXGmvWspr0/DtHJymhvyBFP
3pektqJlYU4B1eKODImZDizDRWKIHFgBUzZQfa7uJdMUcSdZEu9nDn5POMIv
tBNZVOkaCQ6FYQlFEwhHsnuow6E6H02/cYIR/Dv0eqW7Ku6DFIpWTpaneCMa
jsTOrt4JMrzLEHr3QjrnhrZd+77NwK1ZC0f5R0DrR+elvlEb288wWdPZFtxK
W3Ap7IB/TTjhdwqXV4Q/nPjVOc/+Mmky1IXbH0eJS86uY1hJNcJMrl/zMisW
WmWHZy8qk7QxhY06O0j243/05cwRN+5gm6WHDrThFcXxMQQisnkaCyTynlZm
15m8HZwFWV3oWyDnKOKbWhWARdR1bI4Du0Wwk1UbFN4/jUhXfXPGsGwmB0TG
525t3rNN2OumPC3SrVWywoJ71nnBAlV6MRkAZ5+QmUzRRS9zMrpu3sJYihTL
6R5ZdXkLRfkUmS9xWVyFuf0X9V2HnSXH/ENeSgfQtwZPgbRs1y3oH3vZffDP
PySb2p2nkclK2Phv4Gpx3yfaT8dBhU9YC0Obq0GYofFPnD4zZi49/sD/y/eG
0/jOACauSsmfkBgdPwGFfulWAd0fiNvKvQd7+RNzs4DYNGcma26ODVm6AamB
AlKTAVfPO0FdnSlJXPyrOnOr/TvoTt9tXBzHEcURGUc7b5ovmVYhrXGHhVpl
sbBtLPe+7H6ELHvha0VXV8IVIzE6XXyyMWGJOvwQgM9dGfGMPka0oV5c+sp8
fIjaiFKT+uh6m0xIf9yLD/WBHp+rglv12TR+XDGNGk0yCchvwVmwsHOZGwKb
AtIyUjXh5ypfgvCMYf6QnddDTMH7yDTJQ5DbYRtXsWhOSgW1TMSh/tAVyrLR
ujNz1DRT4yJXQFQkmj8MVFjyjK7oJG+1c65T6sIQHWGD3fcsxC5MoE727thk
oeXvjDyrNuUxCberEsyMC9p/CbZ+Ac6RJrkjHunx2hSKCY7FWTjgrbuX3DKx
iYTIs0eP8beWC6cYn8SB/mbdwwS2oXs4fltlA0QfZWLkrAtTFt2PNnYEVoFY
bXY3aljONinvj+8bvBzz0snFuiklntGVgYrX+jFx7M94aA926vU1+1OLYwvZ
xt2zrxJM5pEivkKaZQ/HQyB+R+CtsZfYHIREKi0AWWTKgq44nTRwNqvu/tW0
WJ5vWHULR/sIR5wBescYB/p8fy5W7jyS67o5+vbrhyu4XJiOoH6XJFRPYDm+
FfivUZUpEmwoyrcNd9udXuQpRUdPCuuE/jCcvNbHaz1vtj62e8KWOSIbfU9E
G8F6sbAssoCtT29QJpw/zBgzC3ZTB4dyr62Hecb6QQi/36ZmEvyk0LkmoJFB
lmdnsIMQNS6T+/qhQNdR9g+X1j3W7a7mGJupJM96SS4f58L5I42xTKfXtZ0A
nyJ4Ao2ZlbW2qx+YWEgvM472PuvahuMBYVA4CO9LEjwzYHhULc2P/R/uupci
enctFzHsxprmWcTFdoeEuR+BhYSaxDHpF/k3ZB3x5tDVDtuppryPONnUjwSJ
PfqpGNysvXkwZrHJLUYzBYGuNbPVTsmFAd6x83B+A4Sgrb8PcgGbjAYc8Pec
0rRaVb5KdnEv/VSFKkebDmnAynICcVvmQxeb5SdjJ1oqr6WPRfkTr/stIdcL
BSugyo82POjFaFHcf8Uy6c1lsPrc8ieN3MCL7jJF91Lyfvoy5UFmfYM5CLOi
nM1b0Mi+Lk8bOm+ZPes4JKT2lblc/LTfSVHggBXIi96qWmJ4rbU71opLVENb
9eOVkiMhqaZwPFn1iz0gNI1JWFfbWvC0b2ajodtDiwG9IzRd54GuCaCytdeD
BWmiHhoDEH5nFQzSneD1N7oV5FSKZ9EXo3tFYZi/kjklbFZS5mNJcOhGLXCR
xNgmu//IJNt3HyMIyTey7PZOeQ/hX+IhLWH2jb/PWF3TcZqPsKZnTTXRh10p
PKZXktaZp+z85aaY1wP8qt6hdG8q3Max9t4OdrcYvhgoPKA8DxKEa6P2BBih
WNcV2xNNfA6XmcquZJZg73UsD8scBFpPAfMPLrcHEDwemwTazBp9tkYe1eTz
W2fnOqLIhyjP9aZ2eyEPwWrcAjpS2NPcW92fczXi8X7i2yO5AuMn7gB1gEsh
71CzcHhr/sL+u/4miTgjQm9KKlNNgsFAADlNz0SnAXAyBTAJgLbvrCeeCLDL
hec7xcrxUiLdDXOCBXZH2AFEJalEL0mXZOLqTtGpjOTY11wfqF5q4YmcT8Xa
76M/Ab/ogIuQ9SHPSeVe0ynoXGX0bginQDBEOV6PK1ImqMefKipXFgawI9Ds
j8kqFdpL5C6Q+W8CEX6MCjCXKAAPv5P+ebRif+w0hqE7uMM0mkXESDxlEJVI
XKwxGoAB4VvlofvAYTaXdQXd8Pj9s5dQLM+aWmzAiOtlskTpzLEwQ1MiFYxI
da9Pb0ViOKKcJ5FyN4utyG0Xn+jkE9PJoSWKbmQKm0WnjoQX89yofJ2e3elc
SI2LEzbju4k/cro/X32dmJ5OAFJXGd4bq/n3pmeji+HW3KafVrbYo20sJIb7
TiyeT8rWJ7g0KkPWdCqbe1DzXaDx7lT4LF+JCD4Ax9FwQi0CAxyg06Wyfpsp
rp9UTmYMTw9oo5+KmUeZD/4DCBqY85hvYKEjBkJG4IVoVm7NZQGYdiuG4KkG
uzD/10kjjkFrJ19m9ftsMAexqkvEzg1BIT5xTPXjs6ZJ5d3qTj9TRSmJsnSl
6zUJeVJhm4wsSC7ArfEU89GYhVXVHHa20zVHUgPLdflRtXXBPandp1NhthO+
Mm3tt6P4hCmRhONDaZAHGSoyUARcvHB4s7UGyEDoQH290aMdhb0aeoI7xBlW
+zbh2LrafkkeunRcWuU1LuMEJL+f+TvkOE1FgETLQrpSHupWMt2i+dxv+yve
fHLqAIs/8mInnFOw2QTy2hiGHF6yxG60TtOgcosQhcQ5iOOCXtLkRJNlE+Sc
zqXMuJg4cGjptIpFp2erA1Yzi3/lkZAVBq1Ab04qbTDt6mEQFFCG2drEDcgH
f6Ji/5jKtUQihkZLevvUxUuQENB8PEIbFZOvJhZcVk64piJLF3EUCAQmmrQn
BbeDMXRiT9cik7pvLpUOgnkYGaP0JZyDTzSj/RZvDeKmGR+n2y8gOtzeUY+9
c76rO1l9wUZKdekF2LT3A2ESox8MwBK9dqqzhh++BvtVUiMQNwapht9p66K/
us6UYR5azNpcu0PVmFf7TfjpmLbq6encnmK5q2C6KPtytVZHJWYGMb49pzpU
Tswa9RR9FQvHaI5EZvMgS+TZmvHN/b/gRlAbess944wy2TAwYgxU9sEr5ofA
yK7qI5rpZRhJ4A6Ufy0HVfMYBHdas3XWDfQChVHqkpNq2YBe5ke8Lu65rOIb
sGG888X5BCyOIGSV5A75Qlbs27/SW6mCwKYWrYCiJCkGHe1d/VVsSEGMB5Oq
/ptf/o0sNSxuD6y1lJ54K0oMIy1iq3XyBJkpiIZ7Sd9ZgZw8+KFSxxqg+oSU
nKNKtEVMwEIU6HkStDeUGO+3dCZtwDPq1mWcKbREqMb5QT8uwNO9dYZ+cIoQ
bk4VdvvK7+Pg3jnFN3Bdk1dOC880tfmprbGd0AXYKzeqd7zBaD3AfdPQp61Z
hrddpiir7NcMWhNHUHSz0ptryibyAAWsPRZQpHbGcIhKddkOWPQi95P8rAKc
OhBWkJZX2SHgJJAd+kQ+yY3gOpuZ0ulCSnrsJZW0JuHAWQUtJ6zF8GNJH8V1
Awb5s6qnutdM5vFGUtSyEcreylu+K32Ay3kGTJEg9c5CjRcYoCSwH1104jmN
fOtgUGFyPMbESDZo0gcLEb5eaOXS0F+u+a6Gra5IuKgez8yzl7ULtJVAWqI8
Wh8OubtFxefsbnvWrsiHzgJEqIchYITOwgCBXjJ9Lbu/w2RIuZ5qAvmY+3wK
fqLEr4JhtvtmGOTHLax8L6mkZmezYjWj0vkH6Nrg3NddiUC71MjjLS4eH/B/
Bc1gsDFQAFzzspHdz65fETp87ONN1PygyHopI0zWaqDbrY+6uELK8oDekGCF
zJlgwosHKJJds5CjEf6pkNAqrKfvGHpaG716uuPQUEr6gneOHgasZgsvg8mS
f805/yPPXWfgwNa6qXYEilW9NFeNJ5VEibp7Oo0uHa2tqI6o7s20/eCpWDkN
x5a1V1sOt77I6SCDqvccvKShx6LLpbTzgstcjOwdaZZV0ts172Du+nzoM2Fm
k1cRUualyp2kAERccMdwe8YdGpZwvPPZhhrRwioa/rf17T0bt7gmnMvJRSg5
zeKrKEvXfvn0/XCFGXKG30pTTP3otHsUe8+UISz5dz0i4ckRnMOAVsCkEQJK
hn/9Locj7gNKPnCur2c1kpk0+asePZF6Lctw6JBfI3pFWP6vnQ+Hd7AGhTKn
Zb17Pdu9/Q0IsbrOuPoeKqfuaU9aCQZwWMFc6igsJTtx8Hu/bqiHKglUwt6G
QW8XZW3quIBnGZ7esGFUoTB50W7UQ2nhCaAdRJTVwXLb5/4hbJwC0sWRpQjh
qqBEujkunGgeEckxLYLUAq7s2VEf+K1FVhN2FU76LKBeyMiu3WEY7qQf4XXE
CIBhIme1toXDae7tLQUUqvYo/HiQVWHRfGzXgGpbFzvYsvTLWrCpzeRH+xbH
PWGkLWtDssurEgtBqv1HaiTr7CAeQKkdcGBRAwu0fygx9Q/zYqpommV+oo3A
0x9P/DlGrdbX2Dq+XIVlShRT4gFw8L2jqQ2EjlbzL2hBIoEEq6dyBSGbxy+B
r/o8UeEmzHDD/OWDQqOhih0O2nnhEbMg/N6ycGyXabHKibe24176zToj6TMB
/Fn3Njq4r5+oQulLOsdzbXyuf3BndV8pnU4xiAAS+CT6qzCEbOWx7VH3tH/j
q2ICcocjI6VBV8LOYjN/pzYpyZiOjQQaZ6pFNTTCTSU2NGQ7bTqou9/7tmXl
nIkSp0bGHc6rqKXPtCsTe2fjpJ1rkxNnV3wENFIg5qJbEB61LmXeFWc0HsUG
+E5oM184UH0JypwCunnlb1JIjiy6roL0Wg8nwJvVltCHtGOcH+nLUcnoZMs1
g4Ui52bn7a3F10qSas7wT9WIPRRnBnQY6hx+R6GWDO0WGipXgo+C8K9ki4hr
XhSo6cM2HZD8gTj1KPb9PHfGcFktMtakkBW7qZOMIOFEBHxyQNZJT+syDH0F
1AiJK+jJAo5c6Pi4GzIKPDd2lpIDZ7QFjQDYkRjKie+snaYhCvaHSgrfIdwT
Ln6+xX/AEmkB90z8jSxSApPmPCduHvYmI4vKrdcN2YtnW9XnARZv7crMOThr
Py1LUSyG0fzDKcBJdTMvpr3xZ+82t7pE3AOEY9ORdaOUIJFFeyYARR0XwioU
uzSsqJO4xmBul1eQkd7mHi7CBn8SyrItM4sjCk9coKKC1y4y+ocWO5+Qotuc
RoTHTE3kIfOsQKsCBcoahvI/NdPNotzhkJjZvx1WYCmJZruY2UfGR3ThS06z
VHxc2eh2yxx3gTeyjUpv3ClgR9y117GgiPPSLPAXg5Y8IZBuNW8RRZSDPqoR
yuY67BWU3bVITo1lJmeY3P1Kv1+UC2QGUaVi8LEKawp0OwxrFpKvpkoMCqsg
iVu6y7kQnyjv+c2sMhVBx3rxv7PeXO2hdbmTfwyVnmzlnXWET859u7ZCL20K
YDTG7XR8u97aMMG6InNS3U8kmEBHu4uP12lTl0BuCgnwWJNnZZ458Y+/NibR
uHqSafMzQuNk5LI4wj9dwLfjVMUXmVTceX8CHxSu2B6BbKYOB6wXvl33VSxW
YNYDgtlSTElqz+2WcLOw8UDOXwTmnBaceigjlr+FnIKZXGLVZ8bihW9EEcuG
TCk85CjDFwXdUGfZiT/0fB3fCvyZEfSYy6CVmxcVanPZ7VFzzB60M5hqCtrb
B8faZKlzWkqDpcBo+5LUo87RyZk74/nTN+MXs2PdOC3NXrUINMLFtQE42wt9
zeBFqIt20OdEaAwiyTbWeftTYytLwDkvYNMil3pQ1CN6Aoj2aIP5SClt9lI1
TAijvoJiXNxXQn+ht4fDgUZjdabpiog+Cexv+j7oO3RNj1jfLoWUMSecNoer
jE4eGZ3MUQCQpJYhO+Hsj+wadJvTMyhf8MKs5F7MH9aHZwPRU6xJq0GxyeHo
L5U+UYrkO5VC7HcazHFEJ7sSANll3Ors0bXRH6WPfxcTgtIhsIBw3NYPHa/T
XA7FH3Qu4eoK7FentSAUdqLM5dzyDNRIkWMuTMA6oUQd/QxX0kiG0P/lBLCd
EQSBO0EwAnxYjXFmDQ3wSxJsY4fCv9sQmqo+X7aMFL16Z5Yr2z+0wWeQlQey
y9CEx6gnsWo39sgYOqfpGHvV9sLjydfq+mgDoYYEDL8YJ3bJA4py4Ae8U9Es
mAUhb5eQCnvXx1xgE4titRRrW04UTvqgd//oojmI4S/KSK/uboxkTRCaU/Jt
5b+VtVxgBlBjAkMssdCs4isv+SAX+WIbV91Mss422lW/Oeb4lmgeXGvX5zVa
XJSh8MixSVR1aYeFOiREQi4p9+V9Ue2dAsuz5GGnMFvybMRCpFocNay3FKAd
Mun0oCBY/14qoU9OO84Ank5bkjQ9kCNRm23HyVh3ju8qxeGuYbL1SgSED4ed
w7gsug0TRJY8FiJpu2JnrofdntN4HhRVlI3iDxz3BmJoSa4CYtGEsdc7lbeM
VTbh+s2CCaAQOPFozKl2PgOHtvdPQv1v9wP93Y5oitKM+dmvy+4juKYCrk5k
5D4uhIMz0WkAEE2Wd8oCkX9BfzKgtRi0sJB1VgvCZbSPb/ZEkQD0LBS/rWnc
ZIPWHgkSZ2PPIJH6/XhdGRycNN5rVMHbKrFKNWhyw+fGNTZrGiZYuiQdt+Hx
GeJSM0rlkVVs+ug41r4zhFLAjkkQypcY+WyPafHtqunboljhheEbx0Nlz/5q
/M7ToQ3dFfgat+PMI/qjAQBQS7B2CMG9oHRAtMiTbVcwv3tu+iGraPxzuSdY
+lsxcQqURjOf8TPKDJqoGpS+N0Xg5gDR/+T1BfrAuiDEZ2Etwr+Z98mOE9BT
cPRqACqE8+l9OxSpTXwxkJ7ShlWEgau7/jhlM8Pf0HnrYCsRcEG9o3eYygqu
0EmhFVYoIxEuUekVx+hkqRLS56EdWvRnuR14DPJggF1vADOw4pMpDNDYQcDV
MV0TU/3wuAnqmcgcu82D5McbtOlMymGm9Jn/K5VtpZqzV1f4mZlS+JT03uaA
Z6T7eDx5dHZHueMh4Qco6lR25Xfh4XbO9uTDuIoeg7GYsVZwIVG6dMFTWnu0
HbMSKGeQcNR1a0H4duerRadMsizw+Zrv8E8q6ZTplkE0uMvjXDJIEKTH8HoW
J95WoE+gU92KDE6vEOAw8AyqH6g4BIA8RdB0IDjCh3TDsX0IIchD+y+2gLfg
ngswuSvVfKBHx8H6aSxk6NSckUaCct05PsJYIPakuoVkHTWxnpP8FDzRk/jy
RR7IarO1NHNjQ+eO4Zi2Ew4HhHA44x+xWqaN6yRa88ZQlCbXolhLbKVfVEM6
PleUyZ7Njkk8ryE4TMeeqwvQMJuSNbqOlKkCmUMPs5tyIgDDT6U7ED0FdD61
+58TU10vKLq7klPNs2QXfgyT7QGEUn6ELgVWM05fRRbtwjfCoJYKi8ijRheK
zabF2QVLPbwcA7GzbZ8NcYxLxyX52AyOllUf4veQuE3AOW6d6WWi0BRqbz5N
u9RKuZNxR5PQtHCbvPkHqFAAlM8+VnK5ONHHINM+D8lyYyDwcJ/GxYMsXO7G
JDh1nC/S8WC4rg69wmfeUcCVBixJgpA4FidTYyC4A5d2Evu8Ygj49yN00RGC
jBdNzf2SkhjA11QhZP58CR1f9dmQbz+WfN8ogQ4cxvMULihYd2JAUKmsrNPk
/WjE9hqQoCSiV41LVgNH7JME5gj1TEzGYNGVgORDANQQPheUNj/+/+07U0+p
g9m8JshUp8kBlI6m8cb/wxlGvSBrIvD8vTApQxtu/IRsmRD+K7WxEBjD+2cP
palRvzZelre/GlI/M2Z/gQH6DxyuLuUkIncl5hQGXxN37K01yRi1++nKntx4
1OPmbmZ9g5roTq378hQg5VK70ZzupxiJE02gk4D9txtviyrmL/Nz28ZZPfXC
4BMrLY+CXrRmVcoueTJ8gjRl5zh3HRuctCkRreUfQhaJcSKti5otpHYuKKAj
hdOuMAllS9VAcaVvMMgX9+PBlrw8K5V7DpDo4T4nIQT+ztZYRSJLxC1FICZ7
kfIO1xF8ou7arFoDBZrulha/iPq05LH5e9e5a/9AYBYDEjW3TsIFXuitb8xE
TWPWI84oqapbxFD3WYkaUo6knuhPzMspqEH0mDNaG/FMZ7oHFRSCseKsto3f
XWN+dUtOuc/urhhESpNhSWwJRQvVvqePC0S+y+Lh53+ETnx95ufTe8u+MCxN
bvpy3JY5rkEsYOSDLjni494ufXh2oqg10aFOVt1umE7YHtWA9LV0uaNOmWnu
1nPjFj6NLa4Fc5DTso7lxRziYg1YxlePeT9NQKFYUzroQSin8jFItiFBeXl+
2LgZsiUs2ypQgIOxDfxmBBuNHIO1HG4rdkmg6akHPOFTMmREeL9rf2x1ih/p
pXOknwrL3AInLvYf21WA5xg1P4RegXtp0D2sSfPZLb48LWaCuwBdNtYTltut
JFnbLtw7dDDBRdU55HyW7gO/UNwDsQCWX711NR0bX8zN02zOaIXpcHnnzqPm
1qls+U5XKnC8khJibHfI3VJZsiOSuo5Q30cIwQ3Kgk9T2f/hA5lRqLEf6566
1xyQkt4dHSzv+U7Rms+DqAgYwcvdzeAL2K6ueBCfLm73QZCN8hXl26F3AtA/
4HvZfaPtZyVF/kWraZrQZRMnRrsN6JZT0JO/9ZV8Xasc+30Nifr6TxbJcYp7
VUU2o3CCEuCvAjFuAZOoYB5PBNpu3kWzoHdeLQHoAReIFQQhHiIP5BEXa7ef
lLEi2E8E71yFw4mt4424QMsKjVLiiaOHWB44wkY0ZAFiknX4d9Q/XLNldido
picwIAf+jA7whDaOqZ+CZiBmkOdt9cBfwkt+ZyQ6PAQgSfMsexacE45A5K9+
VQUQXsp5JECTZiuvMkQlBi2/Wd7lRAsA0opuw+PEcLjlxquF01owJF1DeMPu
L49vJ6ikMOpdqibhrfXIJ1GjDmip5iR4QFcWJRQq7nCbcS3YkLvGFAYwbqNJ
7+wipog+sKhWUiF0wNP+P45a9GFWevtwf4DtECCB8IVfY6BofroKc4ef2Lmk
2AwvxHujXZsVpsyawtQFT7j21lbmPJYYHDNLCQsZ6dEjqJFTakKS1z+SM1ER
DACAmczIelhLfDoqzRcnoQh7zcFGbic6OnAG3KtCQIjWYxagHOiOidcIcYuh
+GsZTSlHPNs+8bZtc6l+9OCJS3vCHqHFQKzvLP3IIFCTAQylOCZjSV5JcLud
8T+T/raZmWKEihSJjFz8/UwqBFR+4+a1j6b1wm6RBToqLQB7phn+Jmin+eXL
GM0hdDOWXA/uCpOeFjBZ5lrPnUVCBrJrTP/eNdiNzhxI2i5SECHBcLG6XkJw
axW6yZUlpamErR06tX1iCB5KSM/7PtUWxs5jCaurFAQNu02Pzc48nyxLIBso
P7i7S/LsEfwBDMfk0IM0XSYeMxqw1LK8yy3Ay9NLL5aDfqu/SPl347MMoH9R
a8KbQySJzNYOUvnrcHGcNjbyug/QqVlAp69ghGJhinGbXirewmI9q1mIMHEx
nvo0IcGdFuvW2c2gqGjZH1S/vrZ2o5taRenl0NSWa6UeTKNq8H8q1txD5qTn
sF1kngty33RoMOodDccl2PbOL7ud90jnv73PK8nevaJ0yo0O5W9qpAf4vS13
BBmWSBCwnx4ZLNVLG9+W9oBB+FQlNkughX9Xf/lFVHDK7ZgDDeDtpTSwKmzi
sEXSqyAj8GjBYQNNLt7VBr5v9TRiW5SdcbCRr26fLmKwIX8/o9Myin5Lik3m
mxZjkirrdeUQfwb13vwPS8mG2pK9pd/EF9T9CgGSsLQZIY3AX39ftQD/dmN/
YhHkkGsTdkJGqsYCpPPMKeUq1/6DcFnhGHWOV0JHtiLQk4PoOmXzNHd5+Rul
OIAe3pH1zWIXYEyOpotUwCvgyb/fDF4ynUMDr6fyZAwauyFv66RDjpBBpblH
XBa/XSxddTCknxiSbIkbaeQpaq5kdFOw7qw14wEIzighgVYqd7qdB+raR1x9
G/darpMpIJuwV7tYwW+4hoY1WEm7cUI89FWgPI0jkEQqYATftKzx7yZZTK4T
sQPGkwn1wkyYNWcMHh/jUHpPH3w5MAhtBJSF8MQQmMScxuJuaeALj54+R+H4
BjGqZkXaoV7hm+fseuvTSJsoBENEZpRxF2Q3JQr83FXlKFF1dgh4TguT6Ylt
jL5YlBYW1LrJtNEMk1sbDYaL2IVgPzdILZV61AyWkBBenyeg3no3jbgZ52Qi
WzcSpOOCplr6ROZSrC3RUYvm4is3kpwFuOa6cES9N/p9QbEGqYM67mq46tjv
O+lRqB00iJXhxNb5xHGzufIyQS01kSwMYbg2ARj++bBo1jdh/M1ja8VkbS1M
eq8jDNBO2zioPN4orVueCSy2yQwVcr7VQI1kjcKaA1lqtue7HJtEK9ZQT0G0
r8Ypx4/I7Vi5UvrKzrb6HPzxfPf6Wu0Nfl6FyibkL9LW8jC7e8PKYU0zWdlU
BnG2AemjZCM3PvsoYOiRm/37+OAUCmsoIcSSn6QoIGW6DmIR/IE/JiL9LBGO
i5Fv3BlncKkrs0SoJjp1SWsWNYGQS1v/0J5blJiMPm94bzRUtH+wjESY1JwY
vIyFU59XiisFoOjnH6+g1Fb8ntg3hC01wdoxCYThPZmtxi45cZV6XaiEKhan
DA1z9PZc8qVyzVjT2WMIhA5Lse16QdylOI23WYtIbDh39vGa6GldclvNQDqu
y3wRMOhYSe6uBB5iV4V8GJVNznbONDnueLiwB5KvArsKx8a6JGmEipDSLYWz
x2u0MVrYleX8YhCBEFSFVKAnS9uHpboOdw+5U3zcM/MvQhgvK+8pRYtkhaIU
Txvx9xWKtp2EJKxrclKyOlf8Eab68zAksD2vEPKqO9EmNano5KJiMgkZ/Hfp
fPc4uSDFKPVMrrb6IJ+SqJIZReMBi5NMH2DAbbRTI24uU37xJwZxxNDcSAYv
eEVn4SPGUpNU402CwTDDAnTwixPxM57pMTlyHKy/q65smmb57KJBs+83tiYx
FN6ouAJc2DKRKt1lU2Aw7ClwIfjdRfvjXy9P3dRytvroNG+6ReyMa20fGHGU
GbI05TdjTk9kzDW8AeTOJTmk5agqBRDjPkQ4OT35V3423vlLl9S00WHQN1Tk
BYVsWP6RSRxAxtzvuGboTLV4hSuXcpWb7iJX6FG7+bQr1ISwt/DDZsL1ZuGJ
veckY21vEMx5WjAkACDRqsdV/yY0SnLYoCJoze1W19JbhFDXgg6TGJJXjZ1x
x8SDy9IkvX7nSIWkQxb8iKcfcxCs/P193rfGF6QzQJpycL6AHJltcQu4fNE2
aW0tYTRvUoG816mHZZ+LIGcmtRFT2LAQU8xWkiUBtZr6Je00K/dzq6ob9PJC
5O2fVyf3xeGB/75GMJ6o9UXZFfeK38Edxi8STrM9yK550K+0Ae+YSzHqHVs8
rz88bWlmzDPoEqVppLdDIAC+mUkrxnA++mr/KiqyA/8FO5Yu82HjtojHXX9R
HAEmf/MDka4OuuvjJDwJF9xBjjeGm/5i5J9tcoMLJIP8An7XN/kA2Z0+EeDK
iSWucVIo287xpzTHaWGhIIBPJzh9lBlIJotqX+XyalwOw5ecldS7HLjtAuZm
NfJ2hRi4kyExX/JOQRHTH9+uDMid9px3fik27xJpYYKs6aPZTcIwZn2kZK76
JTJsVIqmG7lOulvJXoHefBOblXT6nIWKZqRIsfcsBl20dg9hv4/aU99oqWgt
NKk008n4rHiQz+4zUDdy1nL2zMjdpwnJg7cnhEowKfCiT9v9q9lnX/QeeyL5
vEvMiO7/kn4lhS8plyH9cpnEtHZvbiegvGs+cU6jx7hpERfXVJM/UVqTYpBP
sJIEq3ysZd+wJ/ej0qliJt7lz1JgJt2c1ZorhYTB0JBlF9mwUMFjYOzH11WD
/DICoOF1iJMFRpEOZ82s5XJlBNkMIIN5XHSHfXM1Hum2ssOazl77mdMq4xaj
HLNp8XGmSgHPbGgmqtjXmOnDb1cPhMGGqEj7HGyLJvdNPd33Dypvcge2Udnw
A52tcuvPZ6W6UxpTqnlCW4dppD4swLnKdaQ0bIwVJtO+7fZz9Gkb+MLsa9X8
u3RoALmr+XUXnKQxQXttd9PLmUVC/t8JMJUSEau2EtGftL5yjHrqYBq7/Zrr
f/mhbpLkyqL5/PIOqXEp8Jr8IMx2jCwnzF1aULtmwKkHjJwYpjip61kAV2Fv
00DTkYL2mshh026O+zHRCoNHqfE2RGH9e8SEGmvY+tt+q/VrDfoPmiDr2Yn8
Zk5U9jTIxncXBy3Bta2rz+UxwUS4xEpRXZ6SzMOXfTtLmAPCIUunE2oEW5kJ
RFrL8pFWEJfYOw3TZP1m0zqKsfiduFwdAqjSsDS7WggDXul5wyiciZyLVCSM
fHxvn2g0sLA9eYH1l1kEO1TpwOTCVitVu3q61VMXM/d7Jsy7P2+OB4L1YS+S
DPYjOps6kt3eiEKUbkliXBGy0BW5caXnwNLUruT2tq3KfmD3XnjJbWuCjB8e
e6g4sgXCCmpWJqESnhN+bMr3gAYIdOCdGaLLls1PpVcJJ/WvzPs+Scza2A02
4TDeH9c2BqzxGN6UGZ+q3Q9ZhApXo0Y4ekX4pMTiLXiOrtPVO089CEsB1vmf
/5FNfVgf/KH1iNsPVo36aHOj7Kuk5UeQ54mp0/ouLDI9qLBJeT7vZ8nY3w5k
R2xFhNT83ctfR+42u3kavdYjHC7Vm1HlxCm2XEyWFq4dlehQlcq8cw52YOJS
Lu9hyoDqWOXdJqdZPsDDsYlLNFb8JAu4XmfTnn12UfH3er6n1vsQHX75y18d
vGpI+K79sIteeVU/1DEdJj+u883a8sNoUH2CotR438jMMttuj/hcJqnMVah/
eHMr+wVei6G025aaq9Idhe2eXelxzDUs7pQSnuIujJpvuIU5FIEoWGFt37zO
s6DmKy+sShGfeACnv/pS9Z8z/iqIXSEayDK4n8mgTmCDiHsQB2y8PO1aMvLW
WH9CHhn0C/MqUBqM3GZ5pn977IrTFXm1XlDmogEdwO0P2Jp52laEWYnYXFbn
3Mydcjv4SL9i8HDow3Sl82DslbSIO8Ej7PNLyF2kWcppPjQ3dMja/a51IWH8
9YIrj+Xa0g29JnF/pUorRAb6F/Xjpghubgp/at3HKKaz+AKprTbi3y8vcFNT
XkVkVkop10KZcU1bYCf4ELaR6kFyUfN0e8yO5TvYT01PpMoYUbR2AXt0WMm0
YY3/cNh/pL5Ltsfc+3h5yOJa2x8PrtaNvWR9Uj4d4ok+WfTq/4jSfuRx9XDl
WKGqKx8n2Ur9biQvOM1vZnvuAAfoxlet/t9fXrqiiSSuPBcoV1uAxn74bTom
0RX+uRisSYgLoijE/x4k5niosOSr9JZZs0ysD4lSuBskOlZ2qCqpSQz+xJvg
Ca0E/rAPZ/HPWCXo5YyUeDYGjMCbt6kaJrbVU0w3tfa7GcEbQ33X+HC1ry5+
6FpSXCSTqkIw4fpcQ1obTbYPggl9vRr+mPEcz2/qoJ2Nu7GUEPs1UexzvSm0
o1MAlUsRnqoY33kmn/wyW1IhN83chxPUopoVYtaqovdCKlkhXOTvnJaL4hq3
lG8RhY6oDfLUrBn9R0S1wAKY1DfKzed3v03FH4dd034wMQ6DZcx23rZJZYEo
1MuKbLegdFz90p/W9HchEXfHW2b0dsbC3rIVeKldvuXikQMDBUJ2OZ9sGbdt
kzgxqicn82hw+vX/TqKwCQ2zhMMvqtqUX1YyGydo6wyNhNMg4EbKTvOVCkZB
DK++dR2NQe8XP1JbemQ5CwnRNdPyRlSu23XjrYrtyVg5/PyM7phh+J9atdRu
+evT8RlNczgANbIcCSI8l0Ygul1+uxYyvGkQEbFtTrIDdC6BeD3lO6Je0CjV
LiqY/C4pLo8mux6187Jou6shPnTENsYQVpHwk5vRuohS2LhaxtlBbK7yOzLY
QSl9cMun93NMgrJRj7IXFPZWJzEXZYfra7nXRUwp0mJts+NryyMcK122AT6w
6L6YjI4bLUPr5EBl9e8L0svi2CVxdwlYm71zPEcba+A4FkNp1F7KfP+jP6rY
G8yRLeNsvuw0u6SrI1xAPxZ3vpPmaVEFysGg18UqPDm5GK+wLbeaDgTcnzI4
vKuc4ijwyhgpTFZpt1AwCtdKXa36kUjPt+LFIQ1VTIJQgZRuz02O8c+bNODt
PuxxHdKGpKNk9KC2yp+zgjYvGq45D6pKRxevI/AB6CazTjETBYPL4MAvYy+U
dagFrle790BF3nnuIImz8H19uZZ1OZcp6tXbktDynzGBTg6ykDbT48QsJn0Q
27KGjorMB6+5R9SCOnov9aJUjTXs99kyxRpv9o6ZuXOFKq2Pvor3uZI1+iYv
TlRxZV/I5BdL8h46t2omLZooqC9SJeV++PRYrJt2UQUMRfPP8yd1spXVSOBv
t9RpuzOEdFWcLpRdomZ2WoSDufkeGRtt1g9Kw7hjW3cK8A3sOOxcUf3n1cbf
GFIzXfIcpOm53aU9SNNnO13A/p5KWoyQg0LX97zBlb+7qqdt2zLcGeVFLbLL
7y0llT7MFgHoOZAWpXCqtYIcgx66qxgHIcH3GFnV1STgYYx7Q0Mh4zoHdmdD
BMGwkArhrlwbn8NZ6h7/pSywKb+QN+ec+/YCm/1UWUeRlt5OHh/DlIGvU9Hf
rq97aeFZNWzi9JFqWIR/Hb7jq24hvo4BPPFgDhDGcphR5EI6znEz6lXIRSLr
BWg+/1xqsgmtWBDSihsdiMxyuBEr+b+PLoX59+4uE10d3DHIcvlrNwkTrtfs
0N6TrY4qxx2wvQlmBiFP+/xTv0P4oxI6CMGJwzu9W8qn2tAcyX5kiQuShD9P
ctikfmDl8xkdkYWePk3Ol9LEluNv93cuvzV6LFXH4O3Ju8LacJIXR5GWxnaG
R5WvVVYSXmS+DnR8sEmK+5j2UVsR/ZkFY/kiW1+zfiVxlkDvV2TYNPriXbr+
e4ZSiYriZ28HZBvGdmIZ/MrNgcdVE0bRXfZfBNtMu7nEZJuRVptlQDqncCBt
9hQviU9MrrnqpJiGRuNUAgPIYtg2k3RNA9K2JXpGgu7yDmwHjWpT+86+6gZS
f/1/hhFEhzv473X/6eM9GjsNinF4Mc8aXHXjNg4VNMsUQjzdRFYwURY/bRN3
Em/+wGyzcDot0y7GmGiJEa5t+UvWLchowlag5mGC90rp/CleAV8gLGLXm0IT
GHpVwvfS6OLuq96gLOP/O0G1BiGZVTJ7lgXmLPvDNGdwGAjNMam726NNYv2C
ZoGzJswaluLReFoFQ99N1UrpWIiF4gKBSVvWvaIFGhmYvn4VzoSaQgJkK7b9
bUaPyBFfMN3JjeVYxiAiLQVcfxrGMwIPwNYvP2YM7b7G35nDfdgdvVCAHfxG
WeOpg2veVVLiiu9lRQtWfRwv/tp93hLFCE2Cb3ZpznbQhNTMC366SZ843hrY
fb7IYB9psupYHoR5iU79RGcTVlIS4DK/mfmrseAGX4h4cN+wivqsyjjSyiw7
H3LOiGY6dPlu1RhWtJ3oOPdFZyLlPdTnfipypOhLcZqLDro5erGad0ovx0EP
laks1svVZvJSDiSmQQqWrmuFcMFx8G4ONvZXhnPektoON+rFyX8w4dl/IGEW
zVoqqKNW77/7UrvyIQZhPUnFXCykVbumFhEfBF+N2YMnAVwgWrd1ToLRq6vW
OAUcTuLHhwyO81CydNYhk8OpoOJT1MvK+Dly2Bwb++gEM/g019T+dY/Heo84
pssC1JY4nu5ECojgssJDA/eO2CrpQLSNX0IYd825aGDo/QgdpvujAk2XJJs5
SyEAhinq8OGIxggs5I3Rh8Ow2YAxct44NkHMSlwR49NH4dyrWV3XLjZ1gn1K
ADR8aejaP+iSsq7arh0OnSJRGLF5JVB9RQjAK6I0GN8eUY2DhL4lhh3fQrQB
62jkNy92RivyTpJeSR0tLMjz6XHnEC2628D8/aJ5JW6iIhBIPb3I7Mn75SCR
4u5brR1XTJiUV8hUR9ihcGUpbdcewfCh3cwCV8SuhQkAZ6JDXYBizYHArirC
j0q66cZGErF7zLHjFSSZEJcT7AWeT+Rp3C3odYi/h0J7JrglYBnehEF0LmB/
Hg53KxL5sFNoJ8+PO8BO/XdOm98LeTyvXpFdSNRQts73o5/NoufUUtZmhmuJ
M0F7U8iWiAcDTDh3zJuNsLeQY/FOWpJ7vxVztCT7sBPRDWgrGoXe0MyCeB5L
YTE51FHdClPXwd+jA/eTp9BY4weoeXa4TRbEbmVcHs1ro+5r9kj1sqYhQyBn
ey6S1LxidURw2Sb3MC19A0kWBiCAV1AoPPVzfc+PWRpUVLX5anIfGBDmPf9+
Pkh5WG9SowugMGf49eUspkdrXDmCbM8XZNuMVH0+6jglxAjdVofc6Xuz/xTr
nXvQ2uIEm5fxQ19k28kfwpEViAhnxAK1PIhimrJ93CscPYa3wzyty0jLcZ1L
h5UAcZClzSW3Aqyr96tBnKxk7Vtya9aOcFlbk2hBxRyoiuxtS46sqd3QK+m3
KF359Vqzee91voh19PcBy6MPX0M5EKfkYnaizBzXCsQHHT6YfpDRvxJSy9EP
YW5euui4ZNiN4bQwQ8CI7RdIVQ+iiiXT6seu2EDKksoFTcmSEKUBhJbWb7Rb
HyoHZy3bcXUMrlzdhtzq03RXjPasg4S8WIXb6LaQMn0pzrEigsPtU+gGswC5
tfsjc9S2yGCEZPhaYnJAV5PhGq26PyC/6odnKMVT1gnsQa0FxeyaqrTo/2Se
pNwTV4SomuE3xPYVMG+E5fsHd1n9OUNjQ0P8mniM7cKthxHtlByX9u/d9TeZ
33TgsVk6EXbjw9ZgJcOXMRGKSCs5PPSByNwi3B4neKOSGWsuCuQLx8cBgTJi
fyCZUNqPnTJ9QLjC7wSTAXkvmaKiLRbnnIvOnNvqJn/43SdTwyKD9jUOuF5k
r5nwmcG86CdwG2rcI+/M04+xJpiE9CE3y+u0RiFB2ATsEF81gyhEhTJiSRLm
mt4rGbawlIrLnRpT4kwg71Ag7x7dCa95frTYcs5GSrvKZRHaT0/LhrmQYFmF
TWwriyVaAuclvbhYVrmGqND1bwci/WeTu0El/qhggY8hGf8YXdVz3gheNDhh
P9Kbm/uSJPth4ms527uweoDbXX+TWvs1aaXJbRoQjMd1fBryYT+eeL/SzmA+
cPZ3X+DT2y2H06sL6v9pm/dMHNPRJ6g8bAfiOyerkK1qXCzAEVnVrTUBT0bR
m3074a18JpwVwwoPhRBgRkC7sD7W4k1bLAwRJa0DcmWtsc/raWDFaHnRt0kU
Kpq2i+RlhUKQriRy9hKMTrMf1bqfCejdRExpOTb2xOHPRebOQUCouXwh2Dvt
Dcf9BS3LRP5KD/7bg69OVwTWz4a4MrjlFMCNHiC5bIdEJtepSx6RTf99+MFf
3PSC9iF/h6kdO+8Jf8n7KQPrGYZL3d+PFjpkmmLh08DLI3dOQ/rCkDVPg7MB
+7qXKB1iji3a0rGiZMTPRnfSwJX+RjeQsFPn9T3Z927ayQ2DxAy/NICB3VK+
ZgMPXKpwRTq6oOpleuD/ehzSyxONVK0NbM3mqBmFrcXKWxyR/m2RQZf5Hk4K
CJIvJRqTwsNMAr5djI9o7EuPCGq4mfAjrkLrwwLlB19qr99AZdSOMiaPK3QC
tQtQ02wsJZXRPRl6S7g0StMFp51gsTil0ZBt22UD+6dxN20DjFVhawzpEGWx
IZG/G6rBpzO1fxBjpqDoRKZY9SGq+Q9hRp4CrNe7qFZi+CZiBszSdc9KoQhR
DjSaf/OAq5jCtwsjh4nuARbIoGY/8pYFnmUPNJWGahVu2vEmm3R35IYURBun
xP01iX4ER1OVZrj1er835w1ppw55dCHSk8ABIlVGUpnkfmMZFGq9p0pUCEMl
dCXScvkpoMhdY1W7NJ8jrizJ/qnIhlpwM1KDXIiJd+c2PouGO654n94mBd7Z
J+E+OYImLmwY8aVkKPfCXvftO2JgwQJFZZv25QKvy+UMPEZWv1AW0avrEhjS
FI62CtfFdnII6r6MQ+4VSwhj/jPShTjTXbylOUeHkTdXU82eDEAgpc3E5N+s
WVoIdhbKFD31mnUxVVXA2M1cEIzm9iSSzw89hnK1Ps9huNeWBxmra1kbiy66
jkHg4gWIU4SYMbk5jaNLFkhPDJKljCpyLumY6x66jM5mlz/cgDVkovYgecmx
5nzOrxWXxBoF+i4sapZsTQMG++TG2O8H7wplzq4uIevjnf/chZhyk5rP1qBH
4WEnwRRtfHI6htGiCnYzskDAlnoqx8/Q3/5xWQ+tvdmM3iyzZQPvICJCh11F
HWGlOBKWC5vLX4KM/oUjl5cgEU3nYDP9GqUqnKDimTzWwREbvpv3tbl53Ebk
DtzvNSQfECk1kSxTe449rqGp8SNmo7MuQWdH2kd9hpspG2O01JbuYPYpbYyl
ZSBeEfJyjhOiLVJE/uAj6/js1RF81DM8FOxIV7yFBI2M6bbOEgJ/dMKwpA5a
Tt0WTpSRQGe8TQY3eekOofWsMoD7bhRmnkIH/KGp7na8mTOHg9/FmNU+Ns5S
rq457JHINJ3bTmtrRiP2zdAB/9SDDY0zc47XgV7EZTpctwg+360w/6Vnu80y
k9XjKx/+WcbtL845mpQ75EoLpQFXWE/RayMk7AL+jSGLmiFnXJHLT+bWvKv9
nFz9fwAwb6sOZ9Bmp/ssfC/2eIOsQx+j7rx+tUkTnjiGniyWTFIAGQ6t43R1
oXJeQ96fG44HvoZkhgwIH7m+iFXg7nuhUPuL1cUYTY9Prp5ko8bMqY8dQ30X
zz/W6P9rENt1NTXLSKAsKBKLznykOks9/YoDryZ7dJbyCSlk+Eyxt29hCzXy
ZmQNrP5fb92LZxqLgeHdkQIoRtBbn4I6O4dkPLnzF02pryz+B9/kc4Q8ZDYT
3zgNbrmBuOsL+9B1xS2eQN7ENjsfTpP5gCfS8iAtMyO2md2EYY1bbhF4Y5St
/1uiJXZHAT48KbPkvGmHoFycTsggFt6m429w4dSebhAa0uxqAZy6EP/z2XsK
/pNB3aQO2EmzbtWv/AeGv2/E5i4uY9mMkrxDYnffOt4JdcAoxV2/FBxUv1JT
N2/Ak18ltXbd7szuufC0OXuBTdueOfSCOoSXWkQPI1lQmiggCKN+OIgNNmeZ
SxFvNNLXyDh/2KC/Yu58cS5WDaVh4+s4fEztQp7PWJp63vy3EvAZv6kgg7fX
JXiEvU7QwonBw3e6ABkZdh4kHkOf8RRWNHlHrlbRsVSaDXbM9BtrQJRGc4jl
/gV95mPa1XfW3hQi+e3hCYU0a8PpJBDMMSEHdPzHq2VJAOZzK2aFG2AbguRr
k0i2hbA2nyPt5UDmhUZNhfgLATdleItqws+kNJW9A40DdaGKJEf+fhtChERy
wGm8AXtTEPoFS3X8gvwcAMWoLtkjKfvPUdqT09C+BDob/Z3UY5rdmdwKhGr1
RzNlMrXqEi77e1n+8Nr97R9e/5pcWY+yoX3cBzrhx9FDrbiAJpGLnGhb3KO4
AZ6AXWfCacABtV6QqMiNq4I6aFTA94u6ISFNtU296RiWQ4i9ywQVlXGMdSkh
yMdyAYFlZTso1FkRa5FE9qmt29ycNVzv5ZHRN1haMmVlA7iIsAoKxr1sHSnr
Bmd7CsmH5bsDx1ajpOtDJUUnbQUh5Qk+M8MaPNIT5sptOsSxURuHB4KTDuvx
XoplD6W/9UE3ZkVKUVuQHd9aosUy1f+wLH1OgVa7+dSbZawO3ixBxU/z9dmk
9BXslziMe/xK7BO/I3C3H5wQtu7gGP14xDtSDlsqY+KayKoJOZzXJysLbOZI
tUxf/Gu+38RqyXoqTAEdvE7w9fCH5Y87tvX0WocJ0jLvMha+w0ePrmgyW2/i
FC2M0YMoXbEW2f+oPMc0ciC//neFo3WuiqCcTsAb/G1lGE3SAJe+Xr9ogawq
RJxyAxSNhbqEH3Eba3HbNPL4Qw4LiZe3v+tAlZVEeRlkOEH8gJO156g8O24F
F6TpFmtkAAmVlSpmyjs0RFCZf2L2RDyRfnXHwsYZ5y+tegSybq1+V9HmYYO8
pee63IHYdVNAaPy1zb7/7ave66StWyjuMjeaxDpFKS7/u78YF5H3r81d1BEV
s+kirtNKIxjMBurpH2PMQBmvuEu5XGss6s9shWXtXIqUJl+s9fHv0n3gfh8R
KZ4sWg66eZpKI6+RYrRh7U9zW2hWyPLx69iahiR8NiCYgO8OyUoUhANi9fyV
OyB6nKarH+kpvuXl8P8+i2NGOryWkYcE+Vma4gWMhvA0AzbKQM8aSHv35hIz
mf6GHZPY/4NdlW0ftyge56kCexMknp4M93VTcJX3ojVinVsLW464O3DTY7Wf
4YtB4f4sj0gA669R3Ej8EDpJylDVil4D45j5wolP1U+Ssj388n7j+wYdIWmN
wfRZovfYJu+YuBB4Gug0Wtc4lCGz6L3RLuQKZ32fKfOqvq45EFF7860vMsdt
28SXh1NHBb36N2zLBqKoKyt77+wCJG9/k/aEjOylz/K2Hzvo9XkQ+HWE08Nm
gWOuqLvBWD0sRjt48tMJ3YH2ADRaTJeBB5QC8dhvztOI+NNz/rWcg3UyRt8r
9qfyTmTca2jvWt91MKbDPctrxd87eCqCq9WOUPY7we4bHb612K0vRblDaQY4
EsmXWhWB5GDafdLJrbNGOQ5GFOpHSe8q0Ba/4hoSF3c0Nh4ex90ZHZTonxUi
cwgF42entv+Mx45byrl0n0Zo2WiwbkLr4Wen9VQ1h1wdY256caOplZELbOKL
Ephm7DkwM35RrdS3+NN3NiQdhn9bNRQbi8VTqpiXc9vfeHfNpxdrAJKRoS5U
nRB4owHu+cyJxMc3NnbVNbdB4uq2Me4ScfOqFMjrmRon+kLaXXz8sdiovduO
w756hjpoDQqjbRa+1MY1vXsYbfOEsm1WPhfF6roP+jQv2UEEasB8rLGC4xZr
YxIQ6ph1XkDjR2qzr82E9e6VinVuKXMUskC6NTdX2rfxkFaA9mD195bIlXGK
L+taPX36OOgjhjBI2MZUXJyVVeZkK3zMQYIF/ty3+Npb+qyngudVsOBaIuIV
7LnXpDuTskuijW3CLpaX7MlUafUzC4xgEO99u45JTOAfA83wrihllUwdDSuB
mePQqX/ZonmXCX4oGR0lKGzo8SQm5QQ+N5B1ogtX+zSUJDQn7kHn67kZo4Ke
0OWoZHMjbMrgPOcKbgEYOBfeHevjEqvXrEmBsWGXf0hqSpSOdwe9HdxqU4Yj
fBFl+HBPN9jCVVQVWOs93Hcqh2Tj6uBGMnyp1zgtUjF0UKVWlD8yvzSBqI82
PyH5bWBMT/5lMaZNo0pH1FI/ySAUAMkjgarmVX5caNxEYvxTqR6hvT33cBrQ
QeqhYODHpYqKZq3ejIHL4YoN1jFNPRodIY27cB0Sefw74/lbtYupON00HxKf
GK+ot77W1Z7kJwR3kudmT8mfu2rugQHTPMffRxhJQ0Bdazlnews+U92aQv68
m0tvChz2WWJmyZV/ev1p02hlZogpcOpqmQWZ8Yw+Et3KheP5iC5qGQperohC
7a5ma3PA+eqWziGYeUAHH3I067+YhxE/6UMzJMiYGI8uXR8ulYB5WbXZUmnH
rrwz1NS+TRu7m0fvrFmlauhJvdWN/bf98G7j7q6zAjbtjLMkU2Nn+0KIb6yp
C1wcd858VbGq/weOT4zXrWhJKNq2085GUWNREHhcfBz5DHjxrMNnnrcHt5FN
ESXEFOGr+xvUGIEujI77Z9Tjqo8jYYOtJVVHuEClpMUl+POXaWgQl9CY2Iwk
8ZcBD6Pk2nMR8uC0NPWUqOdbvZeAOKHKrsx0XjZFTxKeykOQV8o2JWYkQeHo
9p9q/HdzUHscIwhKUrYR0qQgS1WsgtdDXFdTtoHODwTgFT4qx/CKZpHluq7f
7tfrWBW15YxE5IszLyKorHCbWdYrDpm80o4pgMiKw7OLjb2aHupWBB/oj5ZX
empiLsFcMHUjm0ROvdUkNIykxDFne3izcjSi5sQZkO3jLRr5UgaDFd8vQGLd
bblJnbeEvcHcx06paX6pqOIQzr4pbj1zncK/FK55xrYP4Gv99Y1eIvi5nj/p
8OP4kcY0c7hxioQF/JMBfnbdTctnzWTRIzkiY+jIGD+svhon/HInDZZTYLa7
QsN+xnZASAwFLbBNN0CK1vz6rZMHXjM7rbeKIVHWfgv8r31kdmWQdhllmqlf
AnY6O5m2Q1YejGgKhvAgWgvh/i8igJjE23tym6qr8pyaZs9Og13KGRwmDqvV
0f77pf1OlDrKo0kJWjH8WHwnMu7VGibCLgwnDFi156LlMkDPu0/XSqgyiZYr
BQhNStMJzts8kppwD/n4yWLzTLqVu5/Wxf/XKpr5RitvGLdcQiNVGNy/27sX
dpelnD7cwycYSgX2g9l6QFMoq4fN9678KvL+ngyjWwAO1ZmZF5Lz714mSNlY
cCLYAN6k04gSa0Q7LtDI3vk9NBV8210OeH6WGBZpBcgcxuV5BmkSAINxtOPd
GtzVAeHgwf520TLUuy2oFfbcYRvyP04VOoaLVLsdvOqileBJnK6/Rurm0/YO
A02dnOml45UJ8PQ9XNQT9GPLVo5gr0JTh8seduWIiAlQMA2SHfQbUp5cjaPG
HaEo+mOpA//4P+YjJFU6wUpLcDkfvjHKIUq+covCT0edIfOGVSMNpx5AKYC9
BmUxwvVOCTBuzP4/lLsoB4YUvGbWUS8ohaCFtMeRsZyIK6vS0dOlVr25SL93
+vk8CPRyz79dJTepV5K6Ie02pQMEvwHe/hwMM59qYOOHb9vxQdG1k6mZ2RPM
VH6kF27hrnOPTcJCH2cLVRbad090M9j8i576XBFCCgTNpPCm7U6i6kA6UaHr
pxoQ/22OFpH7dPr88ElF5XrRP7psQhsvnYZCpAOpUARUcS4V+10XDlZli4jB
ld6sbcAg5My+hIedD5cV/CW79clEVYr7nK1u2fvwZgewbBZbufQ6sylByybe
KcWhla3pWpLJzWZoL/jx2HY7N/+kuES8nbDJcCOM1v1ikqEvkFDgBNZ0QqNS
3XnSU82wm74zN3hew1k4S0hsunkNJw6/NXCKAhEVXCvtyqKIc16rvLV7GM3E
iCs1j60MqDCnlJveAuo288LQfNqO7rt/XchjeJh73MU6DiyotJXPmElLD9K3
65N5i87HkTbdZKCS/QCeadfAHJZcsRaYmOdqY3N/FS4xoA4MVSEkDmANHDTG
GGb7/COpjWxgYiyAjTZp0vHBfRdCh0RGK3Ma8lnLyjvEKPQT6UfX3ryiU4V2
4g7UnaLCocSUYzkI5Cm8FXqPjMGpBtzWZJ+MyBilPGYplqraQxgVZ/PXIrn3
I3t9s4nZWj9/RNRsLVZpvezYpqsky1fhm0LJI+2AO2F2VJrKeZUAhC59gyXJ
dTPWqaAi9PBFLseUXtPUr+Vm/jOXXoDEgd+O5cu+iRrANy1pKgsCUekxV7/1
KHccWyi0ymrXiye7HMrEGcr6GkzzjHq85qIH/nbkL7OUVwPzI2IFEtye4EDJ
TYXl9cc5eC3lS/dnnU0j/7mUwj8jZJHiGxb/INDw4dKYFc75q6rkMihRtAQj
IvjiR1G9rwbRHnfVWknq1p6hMI5JACNkqoSGNtq5Bi7za56PY4W6rezgOz8O
anjibtIooZ3K0l/cJ8ncM1Eddd3P46KTn2yJccaNIBBQqeyt4QP0ZMgDkl4T
Gf+OiwPle/9ynsMN4a+37kwtzsa7xKljj/PtJKMOg4oHCA7GNJ7MoeZsRqQ5
xYSaKlrESQd9+CoxrK/p7rC3G79VP1btEddy1BM9uB7yuyIdfGCv6hvoCeXH
YZRnLpnooCcDNW6bjW+s65b4XD+s0p1nFs7BcaDZBzNry1Q88PPM5nqEjb0K
N6d6+s35pb+A44/F25MSpaCtMuUqXbM/mlEcqjEst12G4CaKnerQTWQNbNbQ
PiiV7jn3murbpp1Mv4GvQxVJGRxS/sQobc2UAtMySttG6UUx50BoL3RGBwXh
Ed0Y6q1GM1/isx/IJ57l312iE5gAi+tHAReFWCy4OoiKpZUFbkCL+ykoU/VE
lzCx86kgSFH1bjX6LvZgiCgekZj3ZyGuFxRO8HeskDZoEQSY+wM8Bgz2aS9V
We/M2PFIcCSjOxOYgfQPhlanQQLxtVSlq5P8T66Nnmwztp3QXMjaojwBJT8Y
nfX5VEJo4fMPe3hkFuz7DLeqYZBvaNbCg5f622RNS9o3BBUlrlLLFA0TaBxx
eljvOb/j27HGq7KU3zjcIzOcRmuEXoL8rGpGtKHH+kwAjxdB7O0IGNPIUgqh
PZcQSg6kMQTl9UnJ9LF5YsBQjbmnGN4INZI5cXNSQ9IQJJ+VtB7xg6lB/ShP
sPam3LswowuO51fwUjrMqcKdsxSdMXqDQfHlugV8eBAycDN8/XnjUSUFTzGU
gic3A2JIMP5LkgRe+NVf274TzXhlrqqbz5SdWHRWIte5IQqtB6FP3P7B0Nv3
AYW7UlilTSF1i7NMwlChCaO4CfVgZPjhncQxIxRg29OkmGxV9nHdK1jn2f6t
b3LJIpiG9mYLMOwRd3IiYMGawsBa9mZMUldiuPzZZp1UbWkzRTDBkYfHJdNg
idKeukYR9oySDYJq1raWGpM8257DplbNdB4NB9nj1/H4STgKGC4eiR+oZL20
8pZgjy9Y3rJq6bFLGA5K0ZJDQ3ReZe7Sy1omBP3Bmns0re3l65NgYa2ZSyYr
KB4btWulWlq6kZzYR5wesFvij1gVhaGBFDFgjDbW0eZhmRBoYN/NXr30gsWi
1BmDeFx/naW4EQowQeY4RhTwEqV6S0ishXH4Jdz3L8FKNfkm75+GjJMI8OCk
DEPtepWfaGPhVeSDSEz3WR4eF7SMfCNtz74R0P5smsi9Ewa1gtosV+VJCtCn
Lguui6ABorW6To5lj4loEEyAB85j8w2879L9khJITkaQ+F8wNy/V9wpeLB4O
05dAzbFDaH2e4BXv1NgA0a4IZdMwMpvWc19QA1vZKrgxKV3S+n4qb/oEYvkK
ALcAKJBRamDV2UXX9qTBjanChiEgc1rt2+J7CC6dqjg9boRmZrFZ4MJNjviI
sdhB7OSM08y7JlmpY/Iuv27p2yppgeQFsZgfaJws1GEsJZaReea2p64QBce/
bEo7RXlD/joZRFS4u+vBPVWim0FRD9n4hB49m2D+dP6oDJppIPK+mNPVXOx6
hhz6qMmOgTCjQSU/QqWodsWBhMNXdFQ6KfVOsHt7uy3loaASOfJVqqiccQDB
AqHpg5rIBbVgDX+qjsX7teJdSp5miQceoLNTGMx+pgj/FB99Zx8VOn8auhp6
nd5mF1n9aIFr9Co0c7PQgNt37/koZ08u7ABf+do2R6VFgqx2jYgIV4jblqr3
kewdAC0syKToVHJExnkSsGbpvrR5sZzBLfKooOLuby16hjSmGfBtMRZiq6Gi
YSZuOfTtmHtWWpFh45hzaiEqfrrKiIbfEtCUwEbuWcZo4zXwhE7FKeWhXqFq
EimxoiYtLZ84LREmIUgakqulC//YKtsOrWMg9q7IxuxHSump2gTbPxUp2vie
/BGtap1WjFnUgvolJj4IRglnfvvOjkSyE4tJ1zrCPw2w+bUr4AyYmTKCkyJU
rquiuptYCFbZtgmXdA16JTLL3a+/Kp+ZMaow35hPI/SsDOYdlXPh2fzLJn18
LhN4h1CKYKMBSeuUtSeUlsmfnFdDZAwlW5z2MWG8XqnCHxST5l6s2bR3mM/J
Vz1ISOR/j6TZsQ64HC4pLJFuKTAjLH/vK1g0xXWhujeQmwUrRCIRkGLPPWEY
djo01+pRKI1a1aiGw85bDYeO2ZfzacMMBSNLAe+dRNZ9lsxJ01C1zy0K/gFq
5c4CcKObY/RN6eCYdSSA4Xh/6Kkn6i/uyjaTxA+SYLA9yNVljUkQ2t+WyyW2
qFOl1tf5FLmyCjRWauWueDd0Kwu3twTUMAwruNmCiZ5m/b6yqNTY6Kx0y+JB
QqEpqwwvZJn6o8R0vq10D/rCTsUd50Gqy0ke9gnpzwg0tf1qxtDwybttmNh4
spazb7AOv1HXNZg7wbRFIxWSRE/v33ujsyKHPd6lmGhAzsrNere8G+gJkHQU
A+rTNd2Djms1Ix2HSNVTZZ9hQYBLofF6hl0XTFFMboldJYuWL7pEOXh07k5z
Qi6vU4AIwRPU4AA/nlPakRCnu5waRZipHTLLxUvLKzrsLRFpe/FZj37JegSS
yPcWRIW1g2cei9XP8pVtPKca52c3pxjV6xaCmN+ToYqsK6OkdGdi4d0MEc8/
XTjHT2TtPYeSOLLRNPzuYmklfguduJ8dtKRm5LjgjZY1kb4omQILkcL3mbFo
P/Z5+EPQGEf9X92Eaqnl+nuTtGdEGV31V2NIYP87G+HMXwwpahYq/nNP6tJ0
gyoJmaklyy62GySDq09+5SMQO6r5wzB+KWLBl95Pb1lBjzcSodCkRBNEIP0C
lzQ/iNHS9EXoGIoGN2lO74edj94h/6lSyIxmsuBJbPfj3Jg9u2pJSH50V5N2
IRv6KWqOAn5pNmdxveOV/fZzh+SzVmpUkcJ31dBN7vVZgOQX95nmpkEOcIP0
9eyAGB6w0F1iztqecfmufZWhBC6TLqjb4dqRX1Je3R+Ls2SEmk6LKqRRXqXF
7GL1Un5kvD9RdePqzB29Jts77e0sjJtvB8vVn7e8Z+DKjGx1AGxrX2xBBPel
8bSeHu+MszlUor67dNUVAePDrlvYECKtHdNRJT9oeq3pepjd5zsiwJDy06ns
0eNcP45tWwpYAK/sYq/1o8PoPBtRTLLGcHaYHmDZ16c0H6qu90SPkCtHNBUZ
PW0qMUOWqMzY0gUTla3105W2Vz4G7zYLum4KMO6ufDWs1Bia5MEfsT+PS5bM
ApZxxzaGovA6ZYqgIgQ6CYX5SeJhFe/AgdYGKm4GYsvG1VdTmExLKvmAeXSk
FAz0oSlC0nzZtS5Q9aK11L642TfWjmBFtAQh7HXqaVHSu7Fxvw6KRX5/fgfY
HP/Y/A56Mgich03T+O/OOua1Iso6Zf7s/z0iK46JybfnQ7QfIGEEJ65hvOwt
bTuFe5kNDs9Ejh6Gjka9ksczfcvKLqAh3sYyMkBQAVF5Rq8mAXw3VT94MZhd
myFU/T5x91CEa56qV6eATZOyyOl7yZKvQt2Ddi8Vq1Uz9pRIp7ajPOVl+695
nOqnKBvGM1aWKGXWYH0jFh3PNNLNzk6G2IbQ+YNKNDJ+/vxgHBYT3fHRoDWz
r29ogWRiEg5O95wTOcB36lXYCklUUTgVX184Z/uF5PxzMBJCV6bOFPUCygzm
t2Eu6iJBvXuaG+D+A94Cdr5B6wmCy8J3EYxrbBQ7mYXFPgLMp8kbWLpw0eyD
W0v+TGTGIrhIdL6oS2RtcV5rDMs/dDu8vJjyyG4RCdPmDTCGFHvPSHZWGxSq
YIHMkBnPfTnNWtJQ5t070DN4Q49cx8LKOMtApEBfsXLHAHQmUCMJFyJscXV0
WancIwk3bYH6Eyq7O8e9UOttqxnixN0tBX6Xkb9z6UucRyWHcVoQDP71FroI
JMBYo7M+2pObgGtJRthyVGZWaymEQJ6B8w6XOY1NCAVLmjs+3eOBPEUY6gf2
roFmxIY8GCuEEQ/6UTXoTDAHhE5YyqhlbJPEen0Tyo6Y+Y4T5iilwwT3jKAu
ZRmxGyBViTsZBYvzOA+9590YjMVXltjJfRbHupL+NRF6Alf3neJXmGx4WRJY
uGGALxfbiDkRpePPIJ3lx3IKMaQgvOzMg2Ce2sZuLTise1JKGixWT7aS3GTz
wDL8ZL/hI8QSgBiTraiJ9MArMZ1fxsGNzG7D0Dhqo9ZI/JSMdDtbdeK+RAbD
bKDhJxfp+44gaLZP1Z97Q4SUmy1DBBQ3yKen17yWowO6VtNSE3k37qkaS/mQ
d7xz4DXUwUVwliTMLRzzAUj9JH6iuEYY6FJZpptHkFWDH/8+nCge70ohMrPu
3zRI9S8UW71WTYdjK9ajfqTAzcT4uemX/r9DNs6JXiQ4r+jKMF/52Ds130dx
LyptPBx7OrttMKTuJ2yAef5C22dLZnt5bELuaUyetuoS7w0CvFqHJgOSzobq
Xm9FnuSPsO3LWKgKMZWR7rnzfqoN59hHFQnv7JCTfgUsTAgxJE36XNAkz0iq
zcG1jPYwI5uHPNOHLeVr4bHJ5gjs6veAsIkFYfXWfGDI/ZeMnB/F7e42udMg
iNv1kqE94bjwdHLU4DFuuaYttR/km+46BvtDsxy/AqT8Te7y0UnHCBYQpjCQ
S/X+GZ45u1BoUvutPAKZIhsG46fodAS/qJKYOfbmPeUozyBDVYtWq0KEDGOO
HFM6NQH+pOuyZnfR2jO1xZ6mkXzveVA+/OlzLD1+QXba1VdnA4SIQRmQrTA/
oSfzfXL8gigU+0PS4XMKIiRg50Su5yI9EEbimdMght7f7jknQg0Rh2q1PX4Z
MIm8Y+5zTf/S5mJLkpMoZ7/cjeWeFraXSu3ejU6efBhuupgvGotK9EZ6VnrM
pSrBlyKkzlFVBvTWZ5bHmUP4UtJtKtNUqJZGwbF/8b7cIW8L6Vwftlv6jUgg
Ll9a6yvJe1ajxBS+gdcXjK1z0A6M+bkfw3wnFbEsbNrYdl/VONziJLRHuq4G
mod/WSYzUyPlN6+nmbiyTzCiIJwjtD93AYdKaz4GrWDfjXH4cf7mwkeWwilp
fSO1dPP99tSm1QUzK99pkYlFecgY8qnD0ybyMIQg7/k6/xpJakpKJt/+8Lt/
maqZEJJNR6y0XkJPUtrAI1HraiKLErl+P9z7RpV1yjk8uEUbWEwNyToEGoff
GgF0ryaKQAxbMZUrlNq3LECbxSPBwYTHvwbPwmRtMqHFbHk+n3rwxcwDVhm4
KaujYRNhEY5v4KXmCoH62hhhR3SoS2jQFPb9kByW/fq4rpvLV7dNxyr1a0SD
jXcln9DLWvKJAgVlU8KAZs3SOs2jBA8bNMxif64ckR45jBwuyFSM4TOhknOr
xbBcGxIo1lPe9m1Hwrt4cE7CaHmC9oVzBa77IipblC0vztvbP8yLaX3uxl+O
x8ZzcXQXIapQeGXl3SfsPX9QnxiZ9mMtZMxBGGEuCR1Chvz6Jh9e9axHZrby
/E3CRd4azskknLCF+Kps6FLf1bLl9YVSe0Fc1uAZz4uQomcJwyP+8Bmnmn7k
/j7SKA2VbS3VkeueGAO2M7oNOmr0R+Lp+HsRRSH2W/VQwWFepvHtgEp1OXy7
dwof3YAl524/NK7wintFYKg9UEhQB/cMBo1IqxHWBAb+5RgVxxZF3YcdUvut
HSbrMV4QPxkLxW9tpS5/AyQg1SGZ+W2eX7/riQT18c7Yxyo2gA789bW6J6cR
SMKZ+wubzeJ6TI3tbUn8GlmZbcTVvuIOHFqtmpY8KnKVNBEB3jurE8LT2ks0
HRtB+OYsEkeIoHhzM4HTHo6G1vsPsdvppLrQ4N7yo2AkMTlqKx39pJ2HjFUW
lVn5QG9fkkN+uyV2hscBnu71E+1vEwQi6WG4dCaNlnjFnpVib+3L5B+NixO4
7MPgeCNcdNddwIOBEUi5ixQaME8MwIf3ja9UNhqdp+1Gj4UdY3uWF4nED+QB
qbrpUCYZrfNpvsXLKNm0xqBOW+OsSdH/Y1BmrqQmdRhWfpi+jqAj0vDOo4mO
lPdvgesNrZ+sdnbGNAaz6Pl2WPNo4tVeXwHyXgtCwCVmEu+fhrn61ga0XiWz
Cqod8x8hQ6VPsGLER21fxyy/+An6Zn0a+8LuVOqKu7yd9I5eBC20eNcqv0Gl
qef6fQxw1IWDN8suXr+SMlEGazrefnp8zvFTPnt+FQ7jkgkNcBHdAEF4GTfL
3/j112L21fKMT2zwIBrxrsgM3qpcrr+XvkTi+NiJYEVi0Ay+Qleq2VCuzvE2
kooBM19FbzbZhSZIbAV3fSOBq9BWScnX2TekGd2PLOXUovR2nkyGE3gfmw6F
4pLjWTNJ3ZVjEawKmIj2dWnC4kc2R7D4CSyiAbKBhIhinGZybIf45I7SbbV1
rfI8DAT6q6Bg+SCOCqCmjDJsMVwx4Oo32vAXBOeKlzNLat/23MxlN0bSncrn
EVXkYOJgWHCz3dM9pWRoBjU2c7WGjeIs6E0XDrhmtaB0cP8Q+xffZn9cqhfl
IzcW0osAYF7jowmT0Tty/y1BiGVqt7WMpM+baoSMUcS3va34/cWO//EDLy4j
059INvhTeGduo38kJh5WMsZuqI8UmUScDymahJC3co3zsar0ahxEfGonlhDj
WaZE2eFY4OYzAzc/CYTKq/unofpL+AmTQRSvpVcalt9/OWMA8QJgRahYAxu5
iGCp46stfouk/+wB0YpX1iYcmqsbi+Hf8Eyago8cCHU4mWktAMXhdZDBtesf
KhyYDbh3hhzRVTgXqqPM6YRmQAIpKtOdU1tFUt0s9UXiTtXNc8pqVrvKTcb5
B47a3osSnEkIY9rw+ebvwMiAl/ycp8AZIALmY7E3H7FEb1VTEDF1tkzn8lj4
tpMdv3UNTds4ONp5GlFOq0sO6SBZPCnUSMDfKDJWAOnxObBAFwFj6RaB9GB7
qEkSYxK8UUNz5YjB+pUgon+deGRlyp/Zzp4Tz7QgobBhhpK5z/ve6lkh3p8j
AdxneWxwfKhDoiCITBzay6745LM56Ks6SQ2UkJR0/pQw2p3twR+noOtHtVCA
I+r8iO07F96VYwv0FDjWxCkf2jhXFUXKIgtK80ZGOiiIJIe/yCHJW2L7MyUj
B4DZ3q6WCTu9BnTLJ7HpUvn/noOEj5giCk6awnbxebJRfYUNYUbV9jMHgiDn
ONQmqQ05IPUcdXKxvWVSb3Mb4KbKIIksvwVye/o98PwfM4D+QmydL+co+1dY
F6wFN3zduCnlStPglUiXGErue51s1wVOamHSPriaJsYyoWBba5tid6866fcw
3R/qOUlcO7k3L7//hIKiwJnQLmxZDYxyxZBFaumjtipx5saIPvRJ34Ieh6P6
d41d0KMTUPLdBUgCoAXcvyeyAuLfnk3UtzbnOaFqygTlXEtfMyyLBe8xlvXM
ooHUm2N0d4eZ8QQaaLzkQx4+YxLl59TjCeMH97iAj78CoIU7urHBafaYWFiT
Fs+ssXKfETpWJupys8hwFEZUfYRxFX8NfWELvtsfC9vXHh7zgNNtSGPHsxnX
JwDpceSWQP6YqFAYc8KEXzV1C+4JSkCT9yZt2GUM1HeesYcUaaandOtK+RnL
OtLfGG3piiw+/AlcmuWsR2yjk6HD3VARxdZIFBWiY3BgJYfKKzKrZwwmQjg4
Wk0VIsynAcO/jtwz2pIZjnPRCG4o/QJfp3qKKaBE6GnwvwnvaHyaz28W7ggs
PaUn9ACmPyQEoHxPWrGkOvNolkD1e82C/CjaFXPDHpr4vpeDtuABltvb4/nI
5tIYBRhVEj2p3VF6mR3AVXYeS4fK+SrnuMuPDwk3FXvWs3oWiexsmo5deDeu
ucQQGeI5h5YH0yKobcvXjORaGow5T4w7/na2QXRpFlc+DiJEKYWaMBJnojcA
vfO5yK4qK9tzjU0xXA6X4mY8ZFeofksutvBX6nGqgmJHFhmpZebtvAUKzM3A
oDBmkME+FbP27LMUcAVdxANamcWzvRcdY+Xncu4QuNvhbB7WOH969xsJ0/uZ
Jy7CGNJDMMb7A5OSqwhhqHfT3eauhMLVpkrNvIM9r/O6Hxwe1eg+tn1NQKio
2Fh2KRveyA3V0uhnJExjrgQGtZ0C3Rz35ySIjuCe/PbFdYpC09H5ZHw1j/H0
Yp+bZncPxw2yokagvFcGIHEd8RgeWoVk5CU3a5fvS/DgWxPuOgKHoBj7KYJZ
TdgqlE3wY6wxbCbsuHCo7nr6dpEPO6SL6YXoLkhliGKpc+vCxM5tqEDWT5j1
NcRWOO/2u54+YsND7p2w6ZsbCFTIPCOE8rzGqgGpxmnzJnoLkWT9C6ueW/N0
r01yCtQb3ACCZPLedhezPBrV3EyqGsrA9EV3Qes4FzzPEUs8BLBw0WnlaLBz
l7mKOWv4y4HeY/DbEnFvF+S6pIA047VPyA38VxQua4eWpVGk06RWNk172oHP
tslIVMhztBBR57p/jSoQ8PgGI/OdZTT0IwadA1mu5UcOd31x1g3jj3+rbgSz
y4S7G6+I+FvJM4ILRjuEa2WZDbCojaa3k/B5p4e1mgRoPJ7p32YKOfGhjvIF
VOZ3IWu8ip4wsXvcADQ8TT6jOSKPy8Yylwn7gh9OC6gn5MApvJ7/dqcjxTQf
R5PQ+yglvvXiJdqJyBUoLk7Qqmp0PqkYI1qzrTK09Sjw95pPYMI9WtVj5pVD
UpwuKntUqg/UbVgTSUkZFMNXxzOGGnTbEGbXNItDqiZqXHxc2KLiFlugvSPa
0Xeer6i5QPROgzEwdujcGlcTWs2BfeiaX5Ggbz3St0JT2VcNTN66FEwYHT2M
i+5WZuCrF+2o455tmkqYmDkUtut0pQPmffgQmMyq+R1acK9mY+kshfuHYRb5
AtVSPHF4+xsAQa39j0givQ6StTTS1saXqFgJlAam0N1TvNX7q5ubTa/YtfRD
yZgQuW/4H+1VGlaKOeYbBsM86xpYMBroa+O7skYomRZbUTn01QV/zz4H+i1m
NZXjemFYNxCZ6GP/GdPY9bJcWxH3lW5jpsTrGMOOrowSsRSqsPrZRulVJJgx
/s1LVdSKbFU3FZxRPfmqpHzcp+eNDjOjl1d+Vo2TWVAUKxIL0XxBE+wvUPhs
AnUqhtPz+f48qtVD+CdCSMuRwlRu5+iknu/+ZAAE4iKPtiGI+LgnX86IsuSP
uHS2OoFZuEJM0cZHkFCQ6r3kauma620nQxeV34+V8SlcB81ypKDm07x4av2r
G3mbLMDhyVecAVkj1crIGv2a2C5YihhAmminDsUkGkPCqW+E8CuOD5fk5GTu
iXwtep6UnY0A7Lkj0+wlP5Y5GioCOBWY/VY/Ek1s3Cn1puFDwBOMnNFPtSdw
/zgyVFfOYB+PKVaFlY7/XA3Bs2ijRdkNTP3yPthSfSEn+WyBDWqtKQZ+nyr9
Lnkmjc3xC7mtLR5ms1+jJuR2GR3mVCKQVPXSAYc+qvlIqNOaD2qG4LQZ+iSU
SrfBNAqfOldyepzsAMEHypd0ljsAIe4i+C7PDB0b5d1MtSzw5ZcN/1qZtFK/
VDU2hTG4QjH0Ymo4j1PhdyLvnVqbsHx5t7ruWjB1S67LSz5um+qEyGxtztcE
iXlt1RDgwxmoJ7Z2jUwVS4+HXY25cVJMKWSqDf6lrPA0vbuBmk7/T1BHjxDQ
cO30fNv4TvT2mxzvWGQj2SNCuqAZP7fhQ/6I7QQ9/tQibiaBTZ2TXgH+KQUZ
Ew1OcIzhaSm+honYOFdeGUnx1+S12bLiL1DHp8zi1ZwwhmQac86Fgvc2T0Ao
IfrispRd7c9VIav5uPGWNdPEpkbRDQMk81bIKtdiid2I37r4dpylpk+57iI0
+ntTH7XEGriz0u4VBHe4og5SgCXF8MoTw9FhnI4MkxJdKe0QmKiqqZBkvG2j
y+L1Nd92NNw8234zE0vgRxnFQHSEZ3cA3ld5YZtyn+qNuBVmcfVCQtYyPRb0
D85ZKBnHfFJ0ZStQBzRUVwXMWBFteIg9DRxtkyhMep20yLFSuW2ZP2OEqj9S
ZfXRIO/LgIoc9GhMdDsBfYeKujwxNfst8BKlCeUooRCKnqr8U00x9Lj21aPu
vSulmgR0OpCsZaVv/VXK6eM1H+wEMCZeXSqsHQO79Pn67xV57bDgtBqZHQ3G
smYcZrHGtQa2osZxqGHixy29AGb65RYmDkEyDKbX37be1vIil8prTaJvOByc
RcIR+ruqvCmFhXL0Rf3nJ8NuK5XWsXSV1bYlBs2Mhh8RSKYN6agJwdyAqn78
fzEQk9LPrRAVPY2qBuxSVJrLTBpfHli8sRbI5IotMUPCTHz1GvKPN61dS85r
Z0Ns7Jt1Y16Ws0U9EdwDpLWQP7L2WJpnt6C1lNubh6sWD9DHsw5N7uhLDMAY
en/qqllyCOvgnF61iJu0oosikE6HaCINS1BV8q9ibGGakBCqUnu5yszGUubP
CV5WjLYsBqmzhFPEeJ2EleBNjVDtBTH8uuVodgFL3MKp1SE4nDe0BU88RjUn
tluLn8RDQUxGraL88XeivC5XqFhssSi5eTTwuJTYbP62kV4aeMd+Cczsra5w
+Eh9d12sivOiZ9uDipthtyuozo1+dUSBf0LbY0C4yJWJNVKpgPiwERPenPG8
8fjXj2jCnmJ6bpygm85oDDDJZL/xgREMQruDq/6nxQ2JNZMve6hw7zoeLA0m
C7KvZgGu1jFyW3f1NUg8t8fs39aQz3c6KT8I6QIAvzD2N8ySZMUVN+F6VnA2
lP6q6cfTUeMJBcKRv3TamCywi4Ms/NK9/dWK34IwPug7kSWDQ9qyoojavlNj
zZtbTDAO5RD8UKJg69ks5VrL00F/imJtLqW1Obd+WrcWop6WMdUTsKGj2ny7
kctKnFIBauRjM8OpNIgqB/SF56Iiq/UemO4y17z7Rv3ujKEl8bQIcEJMFtGD
YS91RZzWAweDSTh1pUHQakOgZLJEj1FJmtduzOtZbcc8bKxByljjSaWPFOQo
sk+S3HaCK/AHWbKlQW+xpSsaT8VZSr3uv9CCDpdSpMNyNXeoxwGahGyvSYs6
7nJrkEVvX3jcb/vJDUoSDjTrE3kVQxaP6ftWkDq8znsB3qyPzQrScxYRl95q
2KsMHkH4H9DxCj6tdKk3T28Q3rsIthF95ZtJjAaAVOyiZ8Bm+bg8hvcQcaXu
H5bPH0PPK8FAkxXmx1+m2U+H4jZFkN4TIk9jLIEW7slDzzI1HPKtLRjYgR3+
/2AlPXHMeVNc2ZF/DXZlMWh189k8+Q3BMp67pSUxQHTnko+HpU1UKbZMafyn
w+c+GvzrruLiEZf56LLb0UTvn1AM1ULL5byfGrT0lBAwOR7ll92uAnc9gsX+
ISG1QpRO4k11G9NIh45J6JVyv7wk2BPKNKs7rdmamL/ym0yq9Ofm80rpm5eq
Y3yQRVDxOSAbWJP9wxv6aEthOBUrvtD4DW+huXBbciWk5S+ZUNUvtFSLEiLZ
dXZdfR6eNBO3oo2CwfPFGBWjLG2lq2QIA7dxIzRYp9Jsz/I81zVJ2h3bMtT3
IJd4Iy9AHZQbQoMNJ1nG1e/asPqMjumHJPmnflL2qHhIuaPqWSeznrxikT0U
0aRzDBlgj5cPBx0iash6A+j2RmZwXJsqmuiy8gnvslU7LOu4bOVE5a7Aus3d
ROBe2Oq77P+JNwnBepHNTOiyDaCOxL1aPN9Y2qfiR7nZ6BIYVQqQIfhefLS4
0mSVP+CWoOiolFpylUKcyMkinWHvtRyfTCvRompi8yRpFvWmGU0+H0yq23Jl
RqpbK1R87kdQFVp4jWI0mKuv8FmYP44SaZ3BCy93R6zxxLdnQd8Y2zYM9S5H
7CL7Q5+Wa4x/u67ZAT6sFtGmj8Fw9k5tPrNeXqc+Lq7wrMnVK3acDcPQ1wff
OfH6xv61ccfJdIvPb/83f2JvP2b81pwcnmq/xAIG3yEuJ90sLmxneiEHUmF0
ys10eWggmhfTF1Om5ZurhXqh5sE/ZHKNHZ4iy+N8k0HeBJbApS9dnfFj5dil
J5gS8g+N6W2U0VcjkgvX+IkYzLsqX2XrtqMycgUFq2ZhtQsbblxC7LHuy3yR
BXCPXNBBYa27C4gwTNP/sl6xo01E1XzoGYvay1ZqZbDs9TRnyGcHAkZ6v24q
BTtpNQ6aO8utU8Gj8XOGPdTCTg15RCuTmxi6n8hVsH2ruTibH5+sRlMJ7qD6
tllxeS4GiOaj39AFcSit6hwgXt4UPY2sL2o6bNL2wfvx+jnWq1JdnALfxTGA
7KuwFHE++KuOyGY99u7MXuEHbC1LJRpVKOOFoMCRohWZsSbl54zbtkV7qyq+
2BVUA//l/QK04eSt/ZvTKvLzAtPfp1up6cgsY/xva8N+z/5r7WBnXQyTbVCs
e37kGhc196Q9YfpGSR09GiF8C1m0aPooBBNkANwGtaDQ4dh2cwXL+4fJKYPy
xmA17UlUqK3bMLDRCaWieBgZUyqp4pXoMIp8iiYn/NE2fhzgZh1ziEDnglB8
wdDXpLK5S8Y7hc2sF4Y3FQnePVt1TKiz4vcdEXCHUzvbKK72QBSoQRc+nZyn
Z4+AO7bORGIHfJOET3ugmhoDApK277IPeAuXG6h2N4t9BWtRYMssJafcZDZC
yUgjTTZZFFitdwdWTzz8SRdvi1L1cQL0cU6xYn57K90rKy07fNjacOTSwFY3
eTLRiyi+sOtr9h3EjH46y/Z4dIEUx4mCq/YTPcFiGjvh/X+4liUXKsjJMHGW
K45GWiZRqaaD0KXLSlhZXJuWVGyKunAY8hjxbSIy49dtqibm6KVOqYEtdUzX
0b8afYCz+FOm9cWYRr92vrOAel3hqFHAWJJ5P4J6ia6MW2rXLmYeb/K1v7Nk
MgBa2iXSlYNJYi+Ua0yni9sDQwP0Dmc9mUlYgO5cgODdUBYxOaq3kC+LgT3D
NyRXq2WkTZw7jPuYczshPb1XlQoQWg862SOIJ52xMoNr7/S0IqoPT8lthOU8
Wd9oONC5u1YlTBVUFuuc4IuMQ51rFPXc6JfcBp8HhBzR2fkZpY0Ppp7vciUg
PnFLBj79I0mEtPUf5N+ArQV3u3IGgUdd76vHUIHWWF5zoSc1M988HbMvl/3Z
gTfjum0J0lZZl3rBQyoPw8XwWg0L87w2EkcCn0KyblNnZdPD7OY4/TpAkmwV
OAwse8lGernrlaAE+d16NmdWPG0niV1BX0YFnK8Abb1U1xKMzRRZ6DZg93+D
XeLqC0BsJcoN6mnBUWt9+3s7adZMebPUBWq/uMwOx9ds+7NlVOktlXG9ABX2
OQY2rmaWTqbaMD3WAbJfswneShOFWNU3x5hXAdMtGwfuxkT5eqdfcOKQmy77
0PVkq+czpBjvXu/h2O8yD9aojKmo+lO8NvP8yh6gg5wne6N1ur0O/4Duvg/W
sGswqMhCGDo5GjIp1FOzhSvEwsG+csHwzTdVMFD1dBk2Z2GejbUdJqMmMmk7
Etxh+3ZNdnL4oBzUjq1q2zN7JCVKXnX74eRYq5U2+5z98G1TCWuObvqMabBd
3pyGuuzREB2Wgak7o0wVDJoCUKDIj17/PSptLNN/Y4wGE97gtSpvbKyA6TVH
NX60pQNP9wpRMMt8dKdx1L5gb8Thjtb9jg8k/EBXq5iLgbVM8g/7EPceNkUG
8mbM2Af7RtHmeat9c+NqoYAPnohJP1jScJp0FB5FsJOCaHROG5W9T+hqAZxA
lsq5G4TmbR5ML3uJzNasZKJeCZfb3U7ikJNL1TDis/LEuGqzQ8nwxBe8+tTP
icwEJtvSTWF+YnA27D9lMiQ8vUW+iuZrQ08/6g65dvNvRO0nPCUP65ev58Q5
fp+Rr3fdw1NK1V3ruk0IdQ3vsBX/+YwhAfOMnkmshoDHQZWPu4YXGBxS7QzU
+xSjpzdXYVRNG0YNUIURQ1CEQ3e3ttf6SmXiXoOCj7TuDX/1xDiAT0kD6WLD
U9pEFHrAY5G1p1Xu63d5oHwsIX1Z019V9pYEJItrmN8SV90la4yNL1av26VR
z/mO6N00CP45x0X8Twwenq2PZYdYEMdkf4FR/Syblu5s9Vnc3tedWTXHq4ta
81RBcarjlJ6n7S3Z85f2jT0w+5Lr83/K1uzWK9pVMlZy394ebUWwwHPT6ltd
vE32rCXdlpmKciGp/ODqUCwrwGEwOccTV5A8mmEX44l7NgK8OM5L1Mzp81vm
cDlaFLCy95iTmZOIhAGAydCb5suPefq5+x4bTfQ3tzLY0sv/vC8Riu9Qxlbu
EkKl/Ew3XshKMRpxczfVL7mmSS7XrK+i1EM2sH0dz0Z97EYTKWViPwkZkwCU
O8BNvHQMjG7iVIjAEm7XqgKLvKJkvN5ddL2KyQQAd2AgsOruon2VuYEv/gBN
gvFrzg6+y2FCTagEyM7dEpPk0hiq/XHJ7G5m49GypWj0YjztuhBxtb0C+9Nx
N8/LTx/y6u0bg/8Q+tCyoWIItaOScBulxU0oh3vcSVmQlHgTXf46/5e1ukS9
7HC/bJJsYtf5jDQv3i7VmQs26eoqzGU1AEnJuFVaHFw26LGf0xTAD3LVuoq6
c88kCTrwi+a1ltGvxiCEtkQWZhb3cV7/yLF6Mwzol2gyrQQw0J+f3BtEiOWU
mIcLMJnMmlIK4zUmW6guOeLaSlncKElDCmhEOh6w2sBR5lbHR/uMZh1yxtJG
fYok7LYHWRMX7I6MamHbCJecUsXrgQe/UZO4nvVgi61L4yAJNcDI5POpLcxD
GF4Hr4TDRyolOYXBEXIDq920D7fZRuUXs2YsSXNMCxcll+QqPdIWK+9HxH2h
SBvR02fzIoqbFGIpqtqoZtgbdiRzvaOjCdePZz34OENMOz/rarVAcR66WciC
9aJbUgBUDMH7GJGaWwTgjPFpu/mSVt+M6MPjzI5mb2G7jAmwB0em2I+f9G9b
MS2BkWrIaFucJVhw2s6YFzOzaiELEris5+lAIvJatmBc6kAnTNWp/Nlbt7PI
FsY2ZFwn7uvrpiBYVmCCH4kF/ByLUk+lmUHTEKOnq/G5wcSg3VO78wQSDyGj
urBfc6aFQSYq1EdJfNfOsxOZST9x4O6kjl/kpsnAtnmL9uZP8T4UIBPA0RNh
2rR/AYht04msKKbDYHzsIMTVLw7ye3AyhncKp0rSgM+teJuRA9qEVkuAh2+N
pf0kYlBgZaA+X+uKrzJ6uIZNSNbryHOtl0lK88GhEE+nX6pYdb5KRpvJdKxb
LuGb2t/OoI56bqScP+nEFqO9cllr3GwUN/09Sz0vg5LZ+JUFTyKVfVRm+/TF
wZLeO71MdsQTJz5MxOk5c/F/BeRbW6EJoiVQZx7lENUSu3OMeIRLS5bjJbcj
CTxD/CyRQS4P1G42RJsiwC9SdGIZIrmIMJtcNljVFcbTwg4Fjf6mm05nFbXq
5zP3gkpkiGSk2gBKOJeFn/rQHpsw1xe2H+5SRNRsQCs6Aeaw12GB5wnF1dM7
nAnhmgFyl6YIXZcPHeCRqf5scG1X3dLn2g9ygyS40jlkg0rZqqUtmEMk6qVA
RvCXVl0vaysTIsby9zFcSg06lStHvY3ZOKRcGAm+wyKbIvKyEs4RFhDi33jS
mpU8roe+NkpYX4LixLmABFkLD+DPxTgQj9MoX79MCLxz9QafIdVdFYR+97JK
/i1z5tALVZ3+1Cn2Ram7wG5uWlnHbzE47m/JVnJ2957tyKgpGiGcNTv9loJK
LkbIcu2MA2gvujZkoH5aigEIosqgOe1oUX9ck07de46BUjgvDFRkwMgcMhou
M6k3YAWMRuHQ/Jc/ZAFE9d4SGkPocsprI8OwXyr7CidxJt80ydRjfkXgd2V3
nrkAlcvjA5XZ5EVGAhSGXROpQZZKHINmBdCGlUfyZ8VmdKqgNLLtAY57wGB8
0oQl0ggmrtOjPs8wrO4KTW9OeMZhSYbVKuys0OX5vT8tKV1RCSDw7rXtEI72
VJfIwdeXdRkvWKnavxEhdhnEgeVMvGf45twIjI01PuDw1ruhaJ/lldWPhmJh
V4CoBxNpUeohQaigw2cFO+6LU6pX69hJkvuA0tEkQf86Fpt0lU2Z2oLUTJT1
xyRNvsRxMrwpiQIEJ45Z07eoWF8uoEMZ8iEnve3O0ANc8vbnDivsH4WaOvp4
qx4yNfIZeARpAI0uTunFE2EkOWITWgYLZtTQqY5z7Xdep3qQiJ9/GS9hmLs+
ZlIY1ZMkuFc6v3/SWmb5/ZNNu4xFRn2T2PgXPnzauLyGswYOykfULaY2VQep
AZTGcfAIEHtEb144IdX3Cb9jTsfG+eyllxeP1IqJIERl2I9GIeux6OoSqkU6
EoNg0WGDpaHVm0A+eKefsCJ04TEssQNVR9dnLYFBjB84YJs7JV6R3ao9zLw5
Kn7uukMbsaR6MyLQiuv46XAC7TufujKWEv7/37UcunLOJgLZ8U7S+J5wKurk
9/VWXyzipH3oAjwHc6eHovmtfRdYsVXdGVnXO3S5bVEF4CW2JEcEo5qiMjP1
Qps8OeGWrV9ysuMtLuOVqA5vGfbRWI+cxoUV0GnSr0xD7b/g/2HdTSHkgHyB
/YchJ1irfiWgrF9S3aMMCaCmb7xQZyiLNuusT1RsNtX5AM6jIe598AFGsmmC
j1GrswFBlBNPYMdu+Dmy/zGagGn53DF+a9ipdGmOI8IyXxYEpdIXB1Is5uzl
xZoGntDTYxl9YRr+NGjelS8r0SRm3Oeyz7Mqcj+cU4+JmlOmH/5IpsbK9dfk
q4A+ecjBp0HPi5WMtGSC8/zVHn0DpCI0uNAyg/Z8s5nRxoYDQH1MMSs/niWn
cQbg6EV4UnXdrhluYhZfTXpmqpni90EbV/LyqxvREbFI2uJ1H2HZL7tNvxyL
1yVMNEAmZmFrzQ9IuU8QLE99NfZKnZPHGysfc5z9Sm8APxYvmb+q28EiI7zT
e6U/GglOcB8eJTgo17uEcuIML0T8317sErqldflUd3j3YZfZQ8tRh8Q64EFB
1yNxFMRumkOJYV1AjZyH7Que8w6dhVT+W0i92uwsOG36KMPa4ZS3/7dmtv+i
klmuqyhPszcMtSlGjZ/qx1GFLTB55Dz0BMw3OEnynohC/1OJBCPusGNqejC/
9yzSa23GtIRUu/egD44Dq7eAOTk0BQBSvo0AmlV5cMPaPvMJk7HVymTUpnv+
yefWd1Gxt6fBevnXcKL1Od+J513d9ltjy53xf+bEkEajdcJOsaxtFbytciIE
MKWySIG5XZdQyAXjgUSDbXpQXj3FiMEgZVXnrPdprINAlQbCZTU8ZxEEzPKo
uoxer97/CXR42BjBGDPJjF+qPx/mT5b52HresHLlj1MMFLqIqWsV++xGJEou
KzMylhFIOk+mby9apZ6kuWqL+3f7iTL4gmTCZInlfElVUSekKaJEA3ICE8aK
NLeMRVDQhU1Awb75x3gvQcGg3oBMhZCqzx7paI2KdYX8i6kqyc1TV0VbeXFd
AfMKgko0Db5rd2GlV/sdM+fTlAN9+h9N0NQCc9oT4xrLcq82E6VhLEDty89L
eklTeNFXjdr3Tkrzv471dMIuje3pc7Ri8G7GvPjUH0gcKWVgrUmpgmhc1OQi
/Ptq1btupj3Gpj6DHCU/A0YP3dJ2YMh+zZENZzpvl4JvwwLQAYGMSIusReAb
sbDCH5cvVCSVsjrDGHMkmI/f4bxyPkmL/r1VJX1PPvgS9erclAoBz8lJshQ8
yHNy4ny15d/B/Rvb7CcAOWbdGJ1ej6mkBx7n7EcOUc60sVw4wDRQrMc0CdsG
9hwojolZtGSprXJUiCsgPxuoNh+yOc+pWCNs66uR42sgru3nwtdC3KYGR2Gh
2EdRFnkVEUFjNaVjp1JfXVj511+TuJIsK/NF6bPqacNdTOOlc/GJs8K3Q++U
/mGdrVGrws17NFAka+BB3sNfRLIZ1ZxoRJk6wt751UdGMPZekAmqT7rEJejT
qifNfngzYBhZp/AQ589/iYDU8l8hj1X9hydfZm+HW2wNVwtw5kcL/zANgtfZ
1Vw0+ivNozFfLkAr/23FA1KhIgkRhu2OxQ60uYQOp/xS0CTSpl7kQJdsINst
dLsYoFyzPotMVTN0IdyFtw9VhcLvLAHqJX+hRQCSbQHVnTrF1dbNdrik2NQX
lbCedwpvSQy8el8H1q6oAZXtqRRQN4M0zse5xL2K6ZlSCzlnfkdA9iAN9LrQ
WNMd6NiTqstW5VwFo7apvH0Z2skDLPTFUnqJA8vXCwnE1i0Bys6CCy/2AkDt
jlt8+KU3BbqKTVHWofZqiajt/OomoaQ60x/5H7PIZRxqsPTkb6k5/vhE8kEs
ILDK14L1VGPPDd4C910kBhVusp28YOP+odNZlIYZYEUhwUQp5wzL9ASzYPYq
qbt8BZyjozB6I/oQvoN9+YOp7uNVeoOH8snr56uHmI85jSdv48InTWShpflg
YnegdkLmlRro9WSW9dbux8QEumGWA5WuKONRuwH258emwc2lz5pBwFBA9bog
zz0sdX14FS82BY4yC7F6FtUX99I7Pi2YFG/a5/LMehENXrExSwP79Lwcm31P
Dtl3wOTY+aZ50R/ldqmF5fpNYI0GXWF/sddQqdB9fsIKep61jqPdbvoJvcHA
i7mQNS8+Qd62FsBTAgtwvX5yQ0WBp2VA4QAQ2dMtKyyp3DHZjPD5hsSxrtd4
xA2PF7twgwvUc7YDlVt2RIhSPbB7cw1OgzKK8+LhQKD6EKhDnIrhOZq0w84g
516J+GwhoSoS0v4QP2ZNg3BM+Ae18Czw5mwYl61kZU4JGV2WuqcDNSmLu3DN
zUKWGTFLQ444f1Qw9dSUu+Ve/kZihusXTWnPPIo6WCRUNV9Xdi98Pba1KeA2
xLgNtHUI7LW7b7hBQSjJc2Y0rCwxDleudkcWGQfw2ABAMRcsyk0XEqKiyUwJ
F+ov5pN7jppbYYMz+otSOCVq8T8LS1SQw9aOcIH4hTsCXD7OfwLy/Akp35OL
+/1DB9FIgNReIpy0eVPsAMd00gQ1vPkDJK4V94qw6v2BUuux53WhirSVtXOs
8bcQpnv3kduh96z5BJ/1GReWLJavdeAAlcGZsVkpV3kTDArgZDgJig+XQBoy
PGOJUh9JFbD+6EEE0nm5foRctAI1F/UjiSlTAnvolETTNOiWv7pdKcqDKF73
Dpc0SOLPz4xUyLYwrhONfzfQTWQcM41oTPENqnCli5R6TyhTv2PSTyBplNjI
7btLji2emfHHF3qQcO1+psm2ppa3OVSJtyVg1p2/k5SwYoA1sdffDPWyY8Zw
FEoTX4rDKT99uyNe0y/S+n46c1afXWaGeQCdfrl+5U3SIEnuNfrFflzDJISW
sbJiRLnI8JcIFS5pcju/EWXeNnCmePV8JGGgeCJgZxBzyICHJHo/ATsBJhBf
/JTv2IZe9uzaYQEpKFMlaYZe/Ibj3F5fDLzXH9hzsZdifevsJ9ExlfWfQwb2
EiCDy2noujZtLTZ9kiUW7bPgie9tU8xmjE1GL4Cx1ZLJVzhczs0tulfAkbM5
fB/1MUrQcA92Ucdy8UbLlH2IfMdUmLwtn52Qy1xRdPVfpoY7hjlqgQiyp2+j
zN/NTq/ANGOoTkM9VHsFuxe5FS4IbmmengeVvszoQHhGAmHEUfdX28Qo0c0L
wteupWWex7VsKU/zsvmLkSfYk8gg0A244+ifYN2ZTUjIs+/DCbSmIhwLajgJ
8xG9UHanpCzlAuKYDbHYS4brf/kgls1juWaz+bOK3tPBIlovl0SZvLbITfr5
RQJ0JBIZxC84W/RNGoXUB/Z7IMDF6bc4aQ+oJqLjvy8POEQfq+g5xx1pfGqe
rd3Ndb57FIfRhCuCmF19TK99z28Q4kmvjWdBmVoNQ75Vhvrxc4J7ks45vXcS
7rVyg2l8Rsc/VHQwdOs3whMJSZEWDV1vQZGKYtHUT/2DumdykH+x58s9ZlgF
oyK3zK4x4g1R5VRwpvpxWu8bQbmKUOlKc4cLrKwHoEr+lJP2W5jrUvArzfPf
EWy1b/GMXwDkyfuR1f/krCz/Br9YJZdvoBtIMF0BezgxGSLgMCJpI/z0bjs3
0KFjaNXRn8xm335wzc2jtrCd0aaA28+v90Lp0hs6SncifdiZQCyTwm49qNFC
2HEMWR2Rd9CqrIZcWW3sjVf0+quERIQcC+FZjQCRkUUkj+07EFWPc30arvdW
yQGj3JBsptCGFz5fMr6Sz+PWA1s97XpQtbzjgsEW3cPLwZpEZA5a3Eml2Lk3
0CzmjU0zlGgeHj4brua9wUJO20RImuZbCOtVp1DoHCs57E+R8jfo9Ey5gjyp
wxUQFuA6BgN36pFNdWtFDstD31/vblPSdFO9J9aqbW2J78eiDmFElQnQi7J+
rS8O9XxFJUxBzizJdt/6RRDeOVkUMol9HkYbiyTT30xxsS390mRdZL1NHYvJ
uISyIVRdktGsJ9cSJRd2P8e13sB7E1O5+xidG0ICe78JxKGp0Gjnx3cJ9zBm
JAHa1yMsrCjgmfbNmy8Zv7KhYow8UHfprAYzku0QOm/bpr7mRy+379Fl4eOI
9OiDbRXQSIMOWcJtmZnrrtipNMQoovjXP3/HnLWJWiJ6AswoXqAG3ByBAPHK
s5s2UYomFDqNx8CaYivaszb0YVzPfOFT8vKFlmqua2LXfFlM7E17Ge+uSOVo
CoAxvsIoDJtkKOTZ10wL57Pk4c31tCVEe5+JjVYXUt7tuN7VgA4UlFnz+zfr
I6qEF0EhM4TeDd6jBzn+yVnV5SW8yubFrLH3tr39NXAaz/CtH96lIaYWR/WS
CqB2o31sbw3a9wdNNzU8pboUNISGiziTsTPnN4L9Bsd3fK5s7ZmNFEqh/ZKT
tAIUhdbEBiISyv/H0QinQTTgMCQum8f/cFYtCl8iRblpz79oLBWp27VEaYl1
dLHojXEsE8ilItVCOx9IuFdKniSHIV5DFSzYK2SnLfljUlOXCxK0fD6L34ET
PeAGTrbuuqss0o6VtxB961RbNc5P89oaEr1pklwoAV9oOGuIsRxsUdP4+omi
C9s5qqHEJ/3wnxGW0F+mRZc55gvrXF7AUHpEzsWeKMMMZI6gpJ32EHjKyBVw
C+Qa/oK6fO/Lj1mErJUwBAccZMfEkuXmci3wTgIpty6XFKG2cyfEkm3ZR/Pv
o/IHvoVBYmMol6jjh37AoSW7QF+dqIRWUjGzOszPfEKYnDF/xfTFkC/MAyFA
H3I5JZVpImlhteMVTsKkyL8AWNnn3RJk3q9UI58/gs8U9ZH0Z0u+w81QDqto
Ah/l0Eot0SBPaGiBiGOeMQCcKKvGQyQyL4kaOq4I1f2xY9g0khBOl+l/KhQs
e0bdR1rELNM6BymRVol9Qtkt4/XK7doo6AnCFpZ/b41HPZyGr4SxmtYQ7a/b
IVJmoj/0qzll/GfDeT1usesXXHRS63UvJVbatfr1VLfl1Qvyj8AfuOgNq57Z
NGLgmVJEkhr1TEHHdw8OTuwwA2wGpUPP9fVQsk4WDZrGhUT3MzpBN/hG+UBf
GTa+W+pKDAK0JnFQysYT3yEARP5jzviWAcfs65N10SsfjnZ9X1sQ/rPOPMp9
FFWe9Pf42r96IBkWerxtCdop1LH+CH9YPQQg+IByTyed8L46rmzhDKEvRpmO
N2JowyTDcpiBubp6876p+yI2SYju4LWhfJKzX46TY2LaICHab7iC1EA4Hn/b
NzKro6R05i3+/Ms4DopIaMSCzj3hkQTU8V3LKsLsNcs/VbeJJitkrXloJKtM
J5YQlkPvGSWDkOEoIUx0BgUr1gJHQCpVEuNqAmggCU4yNw9OOKN9ng+jQDMk
uKtsUIRIPVC30a1urOnGvf253LqUG8z5Po8wHBTAIQbz1uymlUXjMSiN9QuF
YdiN0RuHuTRebLqy4IUdrgEnStn8BjiERgv/xOxo/NeJcdjdWW59iIm4qffX
E0GuKPlDpClVn1bfLKI9Pv47og7L2ccSdOS5u9iRG0Fc7CD/kuKaMBl668Vk
7cm9C/bAUWQt1bPC8T5xlQ3L5MmLmkoWGCGY4u8vFSKlTB2oHZmKv1ody9jj
F7KrQTLS2bXUAJkfQehV3dsu1fHFbLSaAygf/aa0UYZUoyVSAUAfRogs/vL+
KYVSCQFhaX0sdCLqfdP+mft+jCAx1JHXb85DSNlTn9WIAZUcyBipur9ACyZR
dzejzPsVv/x61wGchLf37aXUpodBYHLCyI8yOsd9eIU8QmC4rP8nDoKUTuVk
+ZDwZ13DeqIZueEvaFGMeCumHemzaShQv1jATvIXAU8Hu4Ed8vUl7UYl8scm
b0cpNBd7Vq3pxYJu6yYNpSc52RTSARKkXq245HyGECty66q5uzMTdUmPzHcp
M7rnDVMmP0GOvDJ1g/JgO8H39s9XSmPxpMswbCJApBsU2Bj1jwQRGDp7USj7
3XGiHo8BTrpgAxBy+Feqjy+qsE+4gGoqhdLgzIT4iNrjTQRQUEOCvKUBRN+L
4crEbcy7rJwz0IVDK/62hMuew9EaTDKBnDaRbQerWkrveVTvzuo8sYpXcNzC
yVD8Q+rxEQCH1k0N+NhKRcUq/z6oHJlKGfCfgkzoZELmg4a/WR/7zlGVNmhC
FGMrX+93haUwV1DhJEQwmSMeYsg9NR/YhGtCVOttWXODrCWMukLRitJrLPhQ
2scABEEM7kqnlXRcC19MqOhtWmVVp4YZRb1DGlJqoC7FEi/JmXWOHnwezcVn
lvWY5IqL1JD6oWvROjx31E+/awwFcCysf2DJKhU3NuRtLemjMY7qPMQxVPS7
QxI6JYKbfhtcobriA7J8t6oZAJUb/Pz89xc9GHEM+66GeW8ldbfSKG1w8+2K
yrg4VlJOOwRdRCZx4H93WW2MQNLu1kaSSoCNpzS12cKtMXEMOZLjivFKui6W
RB2HfAYNAM7rJWPTUoPQOXCl3fQN0AH6IMDz0B1uxMVZVvl+/md7/d5gcoDy
8ol/0QECZuq3nl8QjsQ0I6MfSp78pFTOAGBVRzWctu7bhTu1DwPjzZkRwvYa
8JM8tylx1GZ+Tq9vrXWkmxnmyLHd7Nro84aRtXRIMG64Sn+vBXPFIzo+uM+Q
sYQx/6koxhyqUll8TODZPb6bguY4J0ZYs0/ajWbEKcTGj0qm14WiMDBFexEt
cqH+r2xoXQhz9nj5iDIO2Dp6VPNeUF9Ku84lHpKljWbVO0FbpNIUf0ZyP0n3
2to8RKuOejCRMXq3Ql30SmKoHEAF1rDDFPSoG0mQcZXG/uvA8+uV+i8qaVgs
n8R7mbQ5eM6KQjcMHokLzlubLoxChRTvRPTwpp5bosXkvwbLtxS0G8RVdYbc
O7mOomiDBIyBLbtPnJ0j6HoplKVocRMXXoc82QyiXUoBOudzWsf5YVxaa9BK
g9eKtEfhHGJTvwHorgm7PEnR6mNw2veuKF5afwxPBr/gdivlln6CfKtJs+kQ
OfPD8mfSCMYi04HwrT42QbZQEDbp4tC/MbEmJbMJ+h8OEHX+PuWMR4XE4nrx
1MclRgov6SgA+NSPY/oF/EH6ii//wfXpAzeNrQxWOXtg6McqiPylvvELrBa1
KTpGpH8lIu0cGdDNx+qWrMkG1/7UZAdDZj20Hx3tGDuCRsyzvrI1f2x5FijQ
hx4Hk8vSX7GE4F0sDWWQ3Lf/l5CtH3wOAq3bhxs4Vtx+KzjAQxUVc0HJQld0
itrKUQ56mK4+H4Gp9V+/i24gEpDMwfeklBtMIfKuXKZUoyiar06BRPqHT5RO
9CUXr6V5H8TTacbMWbwHafqcNhVT719dwqsJM4ri1gw392uKX+fBtBQw6B1e
KXNOCJbQKIWdstbppZbJhd5BCbFOKXbt9xMGMxOVizwF/s9fznmHT+CgqBtx
WSXaTNZuEBnxFliQjdAVatsFyiAJUhqST6TbbL5fG/lG7xd2jj99Q+L0yEKI
0n31zRi/3KsULJ7ELdzPYksy3XEIVsCQ6P008MhsCCiLIRonROJGqtURZMDd
P2ZT04AjefSd1U+KdQQWsR/aj/pbZHPzCfQSywKa48pnJURty8REZZBigcOY
/Oo6g84UVqP+18MntgYrzn4vI8SvulVD85EhHK2lTQ8QmGgG0a8cFzNEUepd
gGdy14G5yE19MIfkcLjbolZ6Pn4K29NXlAsVLm4U2u2Qkq6NMJd74yF4hcqH
zsMj3eV/2GZ0p1IUnnGzAjgCroWxTigBK4u0XPySd0UlvO/P5wsCvagYD7oN
bpfpjPcLOaTbIt1BheopWOmLXFIlLBd4096Nr50uHN5yqHguUcSIZmCptrTC
DYE31AlCX69DmdBBlxnCHTXfmJ86BmqyIUlJtrEPoTaQSYD0VeXnjbWE6Gvr
8bsj+nQb9iO+TF2WPk18aCsT7ngb8jRe+V6z1EipmcwtfU4MayMvxeU/y7fs
pN+hbOyctTTSO+DZINQLf8Hv+YYWYwGP5+Fd77n2bM818uWuFQEZv2XksYoc
GKv3JVTdwMoH/CKsnoLX62dFis1cl4YdjyXOS0R8PT5uuqyXsji+cw5CXAAj
Awz/ivYo8tI5cmqAn+rCDz1ANqbGG/WnpGiZ3bOCo1iHKo63ezMBaFLXXz95
L1QITq1gQGWEGev3bfb2t00ZSeCO2lB4t5qd7+/JtJooC8BcXjZrfcdrS11+
CqpF0q9EqnosExTqhCF2+ObBc6pfqci9xCTe/RHhtj4teeoslN1mQ6/xdrd0
zc3i2vc1g0gQQkzBLus/iKaGvmsyrJ/id22mDqXT7JxGoF52X35QT0af56Gi
oAZqPXCm+ddMjOi4n5XxFHGyTad5Wh2SN54tz8CjLw1qkRVqzwOztMKwbP8S
lH1jWphPH8N8Rqo+GVE+hg+zUhTR/GOTNwkBYorVZPxDVzEdnLyKdvCcI/Se
1saq0IjnRmaZ+FoNtm4ORA2f1mzcoDddEQueQXDSU//X5tdHTA7DffwBpt/R
il5uvObGnCzCeNu1ONBpPbrIGWik6fBDjQZGp5rDm7nGPqEzuT+gXSPUdcVl
ylD88QhGADaA7gQDK5AydNOWKMe5gLTnqJcylUc3Iy3Aeh2akkL/mjOV4CEO
RLiWWq/FahFrfi/QwJcP3NNPuxoOTtN48SE0HjBU3ceEP+ONOsB31FdqlQja
7c02vFa7xUBiyx4wCtzLfKNgDjxCwbFG4uNGJW34w+s/sIGOli6X8ks02IuR
UCZ4OmNMfjeHsdXBlMa8DqETmXG+2JdyMndk9Vk52J8+LIelGAIeoKDiE1Gz
b+JLnqapAvWzpe8Cv/PLzon16DL+IAtH+T1CCD8ZiOQZAXSdRDaVljiDAVEw
ww7HoQVpyTtS3rYSUAt3hWgWO1Woq1cgDgqUAUUTLD/Ued2+jADxhaRgkrAa
EM+Th1OoFvSdhMlN26ukkDgbHiqsHu3PB8SkQwOmciHTYCGZRHEWIXHAE+s/
KQ9VKlCL6L9eKR/TCkZ2aHaC2T8hy9kFNjopqictgt7X/P/XXONnUSTjpJ12
73rgzBi9K4ipKJfDgDHNQLR3Y8RosAMDNqqdK94iK2pelONXm0TXxeaKlxtS
2PojNSnVlX0osij6joGd39EdPUqGSNEBzCBaECaQ8j4j6RgBvoDY+A0kFC5h
iETfRq+IPXOqQPewua8Z+KLx6ZJ2DePKcjLwL/0pRouhFsgVFKEfFJZBbF4J
SZnlCTztE49QtgIG0ELmZ1JG7hj7osGc8bqmSp/ojg/lUnvNegeuANtJIxBb
RmrP+YtzoCzjM2IXr1mn0jNYWjasnoi0ljH4c+RNCQr41TPBCEWUGMy9aYOn
ZFjVXB6UavpLTJDHYgLZUOYW5twAoCptjN2Rlyteh1DK2HtVqXIE0C3VcKQd
vRdpb6xAHzCQfKvHq2lNwbkyS58k4PZrLrOsY+7UCNMG5AYoRpA/3MPaj+AA
GqIVVyqbZQIBArL0uvbFyqbHpgylBwO6KpfdctDRPFjOCbe4wy1kHE2PuxY7
+/Vq2r0Q33eWQLpDfGdbl7dLHMml9/uxMxDDbfVQyfQsEshlcdX0/Frr21oj
PINAdItcNkYY7RX+lTnwHNW8ej/KjyThbcqaNDii3G9gNC0IYjWIBPikzlI+
/R9pCsvKcBKshuHrfh/vTFfYN3vpmDkZXfri/w78EpT7r3H5jlkV/ajgQ2ao
j+SqDANsJWB15zt2ODN/XjT0PlzHgBRj24rwyAdSHnjA9Fwgr7gi4D6z1BDS
0I5vJV1O3ZLuL7N/UdKJT/22WSNNkbv0UroASX52IqS2sFO1oL8tg28GqUGC
RNUYJ1cakl4ePm/kKQDrGNgyzdCVMZJNQJev8/U9Edd7HnMvlKZ7A1vv3s+Z
xGp60X3WC5bBCguz0c2QUzfdFESA+VY11usQsFfw4UnAOXBjGc83BnJ6MwLc
qCWo/ZJysbxlZDinYFah4S97TgMezBD3Co8+lAjsQQG6cghiq4E8HejShn6D
r8Uy8r1V/8XtB1aTQBW0xBD5+TnTHRl/TOifTFvZTHfe/7P/DVET5n5KDCgJ
sFR73tWtVs4jxDQS4fOxfesVMrI5RT+PPILrK8pTPo2s8mJPZ7pHXVjAR6AG
7vbVJVS6FO8pmQp1R/JNY8Cc8Qzagjmu6s6WRgpe9ADuNUs5xfDXp/ixpCsS
vDjW/9nPp3J8If+o9D4jAuyft0jXC6/Gk0fMSgyAZpFkYgpGv7twh/rPcqks
sc8v/1kOpOQwXe+C83GovDj7LDwK0bEbX75G19IjjdJJomifBmwjyW/pJOyQ
2bcH+LxTLxcweCwNJ/2adkP0K0jJJWdhYnZwipHAqrBX643rXaNumaCmdfvM
7dmkqyjBQ8slJsujOJ0KFyHYEWWxPJx+p4spKRCpZIiui4pb+EZU0Fz4mLtj
+LiAd/hU/GaR/I42tiH7u4fZ1E2ZCN5NG+uFYZCEZUEcZftX1XiguyGLutD0
bnWfyNYYbRRj4aM1rtLKNqRh/NG0DHWEHN/lbeRbzI4mJOGv3xY3YTskew+u
U7oDFggQBAAqfdhgDmVPVErCWOEY/qhSnRP2G+LoGs8qj/GQP3baTQpBhCgk
4uOfa/gSn3hLtPbldII1iCwKqQV1qbwUeqm1DRuGK38UP7v7yIOIk/06xXCg
mKF/UBhae7RLRc0fR3JOEvSsFzYlrHfptfI2U0pOWJkpzELqb+RVeqQjB+Ts
6ogfWu3pCHvm/10lUg5Bv2rTRea3mhP9s4u9mGn7opmlF27HKo50kzrfO4uE
iyxiMN3lScl0GNeCJRUimLinyN/WnfXulhh2z00BXxwy6QqP2/qZltXcyacH
VZc9SoyJ5q8wIeUMi1tnZbvT/WmcxNkHwVluIWpvhPsGn2fKPl9GSNHkQoC0
237Dj4ldK3qLze9lLOkGZh52brc79I0MDNeuwPcyatvjzXOlhzgDJNCLfnNB
8iONGrEuCcyWpDBKUUVwoRGl5C8sVHuvfHHUF3gwNBGocmoY2uSfSGQld5Sg
KmDnx5dXWNA32s4gFVZ3kA/TyLJ0947jyW+UnTOob4RHD6k4mR/uDCTo64Rt
gVhoXEGQ/wqHzVYZlQcNVAzIqEEqjHLbJN1KPn/sS3xZsZoeQePGSoiyIgDo
US2E21cE6BMFmk4xNZ3y+28XhimvT9cXfh5zPBGMan96GRIbCIgkqHRgXoJw
0Pkcis0G+idDftQpExfiPzGD0g2TJ/wfkbLth04ODcmG6J2Y2caKI6n2o2Ly
WYCiMNsuwm1ZcKnnAWohSs0qlFaiwF8D9H57BNa3Oev10zAzlff5HGknhpSG
5pHHMChqqWSBikj8Z3LXjNnQF7RXGxo522vpNKXTqUESBfeR9ijh0vHfAJsa
R5EAtTZWcsrPSeyw9krvanpF1ft4y2xNf3MpZdRVIXQEadC6Lzmv5n7lJH5+
dekLdE99r8vkSkbYLtWGD4iK5adM5eqsex0CMNVrRfOFEPJeYpApfGdOmS5Y
QjD8DT+s5YL6tAfw+7W1tigqSoZJClzvrVhFAzt/zZ38RhWC98JnpE6aSMP3
AYywYQHCSlcTwPnC+TdUe/wkREnfBaMt8ifTpp6UwQUjKJBGNtviiA1oV9HZ
ZOeQKGctmuD7/MNeZxWoZbUROkIg+k/5w81RzUCbggl0PPDdWX+WMlvGeAiw
Z8O9vtg9UqvwbEt7gJpsPWTiciFbB6PVVH33cINxlxNwBIr445nN2DUvhoyw
ITVVFGjF3e7acVWgqAm6UabdYrHHoqplraocGXn5LV8q9iSv1X9TpArulvBP
laROsr0MRFxbW+f2PAcSauAtVFVJ5aOsFShVdMPMF7M/0T3aJ7Gmigwuvrq0
8dgJmhGq3x6KNd3R8q63xsTfJqdeYPU65+MdO/+IgfXLXHyGvM+mYdU/qWSI
JELxuEsLtCZ/q8ixakM29GnzwHNEHrgk5vjmNQXX3+NjCTlOVX/LtDPMWszA
hmQH6p+8je8WDd1kfA5KkOBojFsuAyrMgpE0wUi+kMn8rQ+9HoYd60UpqOuD
NHUAguUdXLbBsvJU17QbD2OzVn4zTxY1/Tz3UWvqPaAYe4NWCtz4y3wAT0MI
+ul/ooGeoZ0t7KBYS7Jwb4lVmcIf8KbtzWMypZ6k+uJfq/kmrNeCYdB50F0i
0Wq1gSfG631CnAHA/RXwWctbjSfpcEhUgK3eXmVDsmBEOMLxGWG3qxbvm/3x
j+KQBIWixAbKmKQEwNhwJBS8slQ9v8+Sxu3NT1lWQU+H+Q3d3Z1rMAvWgyR8
q6KdwDjs2p68Yfy9jLmncKRB125t4jDloKgTL89VEAZl3aeuLndGE1vj4SZf
dlTC+wMc9lp5nnzofqf4HLWzk6z1tPta4Z6+bjoxxS28Qh7ndjloYs9+7MGt
nFzLFkqXj5mxxQ5s5WXBEO8s46Q749QOPCXGPWovcxpnQpYCVzthAx2v7p5M
DVryV4nkK91qQRgrT1wX9gozZHyTgeoHsXjOXvUNuk7vgCExXN6EzsZewoBW
CfR6XWHIn0O5o47BN184lePa4DEpGmYyQyHqZAzhpQwu4CvXbBsUgi4xCY9C
bnm1bQYVaNjk2P/vcKwAA4V8AXav9Ji/GgI4BZ6bdIhH/FsH4AOY3OSWOhYe
GJLv9jvkFbxggn1azxNFd2J6mfwp4QwgSh15XYoZ626561ZwiOYafvnlfpwr
taf37H524LJ+SBs3HMVN8DN8KY7Q0Gojg1zvbPJpj15xpcvhw2xvkGJEa9s/
B4qiCrlYp9mlv/Wo7GDL1quaqPQ+4vVvgWrz7tmEcrdJS/3v2/8yX3NfG5nG
ZrrgD82q4gPTzPYWcciAaO64kjniIliOLVz71BATaKmPKkpeqdqSLIyqegT4
QeTCAquT7wgZUDTJcg53LE2Cag9Vkxgana3x1xMHnKSLcfyxcOXTGEGMnmbv
h4odHYWPbTXpGuCIb/WbyGJ3cGYpMyjxNh0Mj210UX5wTLIw8mchh2uctDCE
iYMCCnp0PL3mULNgTZ97C+8eHEWpr4X/N22wlA5Dfi6g0KWlT6ZF4dfFfMoc
IfO4viEwa4HcAFU1pTLFEQtVeCLGXtf8qpK3Ocf6+6Lcn0Y8y45PrSnoM2cQ
59khNHmQn25IFXbmuWyKg26tkFmmaZWWNdyg6GqZxcrqSnJF4KqlI9v3QfeC
pR2H5R5QGCAwMBk2de5vtO+vHxzkJlWzWVpoXK/T3VYC40YTkKCd+FeWdvjw
x10ueas2wRn0YQmwsXdTWrCiJ7AG+a0YCVV13WZLwPf15kw9Qh9fgYf1wz9J
afNOPnyHFJP+/g9Dpcm+eXowB7s9YVNLxvAh7mn97pnV8NTqX+3pEnR2Sk1H
mId6SEr87riaQKPxLxBukgv2VZcEqSQm3wEyts2hqirhS2a8+hrPTlQNH5Vb
65jSYx+XmafcSWk53Tavqt7jjHqntEuOpKNqycnvY18OrGOsHsDr6fhbuc/p
UQRQ5O0Jru39mcTgjQwIq7XEDgQQj0SMnbxPaqnkPXg1kpxkavYfU72JaSgJ
ktTRG1nrei9bl6/2gsbpQj5h2nDHhrU7HdPv2ftw5Y7p5n5twcjUs4swJSZj
EG6vWxnjAZ14u4vcm/UYL8U0PM/Hz2NhFO81Bun7z2CHy+cRki+T8ir2/gtw
eEo6MJAmBRddpic8qchP7MgeVByQV/QvHflF+cPwGLhZTlC7LBKNvFoaLrKr
rHMTC506TNR9e9eZUy7UjZFdjP9LDk8l3Pn90cHnb6h+YJmTnHbzd73RFk/I
74Be49UcoJ554vPCc4FQFS6jSIWCnVyqcXIyZ24bgLrETwWyVjX3PMrWcTvv
aPS5bI0in7TxYJgsHPQxdMmztrbBHK/SVRrJw85G1uxz0ewtYTEWqqacLAkQ
eRqI219ctNhLrpy9CMPlEAmJxxTWgbBXvqgiyQuu/VqYvKHqAJ9qCSbA0ZOo
GuH1YYLdayq2H09NTtzvpgOtJ9fHIUsuVnhBZYh1z9JzOZ/Dh1PDuKpaiYXy
vQuGHZ2zY/b3cDf8povXEdk2iLBeDbnffTE81FZbZxk0P4C1m6nd3UJev1Au
k+baxHqJrylpKOyvY4jZ4M3DGEA1ZBt887V4zyaQAmQhBrrFkwKmozJxOUmG
bg8E6D3NppnrfjAUITgX2NbtPIL7TZ+l1j0n890OaWkRRZGGvBvG6HzsUFwk
2nxVR+uFxNBmo6LV1qyA8Lpc0dq+v32J4mgM27dZJiWZTDeArrkQ9vRTsvWA
0vZm7B2324WenDl4AXKcMROnBfMQprNND7+m0iELehL3mRin6n8pO9A1+xt5
BcPjUtM9CgFIsDQZ+GdrWawsdhsx9HM9gmTHdCntgsu80J2CbZTArM/VQQNz
rWOhQ2Q7w8WBZJxqDfvP9UN852FcQV5ICT0q7COQm0xGzroMR3hbmqZuJ4E7
w/o1+aUtIeOgEbRmkC+U3V2i7z4HbdFeUdCP10uw9Uu4AIi8QoPSMGJB/kml
288JMUZe/NSl99mHK6ygSVjiSpASG0Ytb+kvECleuVHWlZR88vFg3jrglNZ8
/S4jcgj5FgcbubGSzo3e5CE+YLvd/X3l76i8whfwhqE14+zKDTNuoMdh1F6m
Gde4ExGmxczzsSsrsPq38tf7fp+LuGwZUVVT0KStP1hM8gGIjPwE49KtoeHb
npPOxI6r5MyfY0EEfDcW812SFgETQM43Mg2oTJNvpANmdR+FSJgrArsQ8kod
FJN8PUZ/w4nOWUJvhx5sleka5p+AY+nrBcOPsceDZmBoHWPoCG381qldKhBG
LBaDA0Qw+PDCRdK2q5ulUnHTXsVU4NBI2LoSPWaU0045DzmkCjlr8w+FdXrb
nxqKqKGpj1fmGOGqtId359K+0MRnU69hAqV3XflWEf5KmRtrwAaKpaEeOz2x
SzEQkcSzutgxZNRQ6sJVcznYmhCfrtl0SS6RxY9rMGZ5/hMwmnoYi4WJ7QCo
oh+i90YAAdZRQNF8Pxfz/nSVr0/7ZMDQOr3qoC98yeCJx9CqB/NuzoKDpPes
hebPUUHco3+RHGnknixMhQNdhzAEGt1Va6mUeRBS7W6si+8lC8F0MBJiwCpk
F6CBAEJnYitpPg5eNsXnM+oWidCjAomQ3xLfzybkCza1MeOKwt70fQ4TPnQm
a1sVJB8fkfdcSPeiiGAao9cbHTg362WksIAMdEQYbyyN2uSLYwF4qpZmlGaR
zawFOQKC8AtzbUI+LnhkG4mkT6TfgDoajiK67EauY7hCmMZjxEJbIvFcz8ta
4xxDIsyOAZc/RYt30Y7NZtMDZ38Q+1tw5LyvF5ICZ/tx8Dm8N3i8E/h/xq2r
5jUqCYrCpb+TQPGgmKX+uFEmbUgSfJEQpUgNiOp487IAVS7m3Gq8R8vNG9pT
9cWvn5bD0lJXwpKEC+h70s/5OvA26wuL7fbMNbygj8yhNmbtf5z8AIDY18TO
Dc0xhb3ypGzmkI1JDEoEYveBpcdHrUQuxFl/fSRmZ4H3r9yLmcxZoYXBYe1y
5R03oXRHIJg9nM35nh2TftHXlcF3DHODoayJC7QaWGGM2fm+eT4dRwUX1ksz
m2h/kbIOzzD2IuF/JepY51DZMtEJLbdi5DHLu1Wf/NnHUFNiHyYxAIfTf9vn
inH3xx71y1gCqHGpyZ0lswgZVx163i95gc34TwEJfTFm/Tk5LOEKaja8B5E6
g14hcIS0VMG5sFDRmsiP49ope2Mg/9eS1JRUoBJVVvZXqVLWHkALNJaAfQqR
ClIFZtymtj4IQkRxUadpC8ej4nbF4LquVdTwmQGmF1Bzxtvfn/U225gjF1jD
EWLHbJJtfj19kDUrO6XYtZMHLjpaVDfRUvwT74xGKUH2+M1OZH38KZBPfoR2
sIoqokmhY1qPJTB8+HOLqk9Z0NJS76fRJEbV3cmMGFaD773ttJBb8NCM7wuZ
EQt9zCMme+TIJ/vBM+KaTrrez+g7JkrLN+BB/1bveDgVIRqtFSwVqmHOkDxA
7f4UUZBo419pPwwwi7m1bb4Oskj9RONEhdsXHmEzf+r3qjB0ZpQdLtuj5eIT
l3HNbRnrUACfD9JIJh7et2vf+7sIlE92ZGaFWFstYj2wrY+eG3A/fsPo4iMK
2Q4DOOJm4vMV6El0CyImRkImXgxqYlew8gnXvLsutKk17rbW/5t6INgGkHis
8UThbzKKk5wWDmp/YbcZnd+3j4JvG2EH6BU9z02NofuudIGDw7MMVmkFeS5x
+PsFYjKvTqpL3vUPYuXxxyOL9I23I4iA9UUoWalztWQ3drzAQMJn/Ei8ntrs
ysp7bvN3EmpxFwcKaC17ppZfdkg6CB0LopA/DIEUKpr1EW6xZaNUl28O1ieh
qyJG9SlEx2zfmzF1vfOH5Fwif0jXZTTWFFUAOohy/zpH6+9R+nTfbltY2chb
uWI52rEqAGao3f7VzYt8bRDE4/lZ+na16jyU/mrMuXA9yPkhKy/RPEZVREjN
lAAk69DyRzQJ14iakcBTL6zQrJEd1/oFfSFu/Ic8nkL1dIGQ+joXVVjDv64c
XhJwKgJuhBoHaYAStuFKI5QSd1Lpj1FgggenDXZcBagpRPsrxq61B5boYMK1
+Ks5YxOVkbviEaVXV1r/YKBb0Lz9umTQZv9aobQPYHfH1oFrU1OAoB1FvOnw
9U1k5Tx7hNFzQ9PMcGSAtyyfTvnD8YMlvoFzebJXTcCb/B4AK3zqOhoF1+9z
aulo8YJNjS29FKdWa/PNDiG4V9WjXSNudczJgo0Q7njONZQBRmmI8uQfpxL/
3yDaMJLtiET0FUgzF1cejLZnSiSJqKIIfHhaho/K3I9efUR3Fo2NA8v/pvIq
7uZgSLG7Z+/tlHeFdlF+Yi8UPG4G1Ndb5K0tUlDdA1MW4jkD6J1Gx5cmrPIj
MvDutvzNyMd7XJEnakUCLq7v5zUCg19OlM0B6PcwUxVTIDJ3WmC3wKSUG5xP
28OY5h+dqlaGtU2ADBFZMKLab7mCGtvE1MlkGvU39mmVHxI940cN3+mUvvp9
BJif+K8d1hr2OAJ+IMzZDfLZPp2OLLjxL3UTQc5RA/YBHe887GYp504WJOw5
EwpSG6yyQQCE4XjwbiywqMesyZyuds8Yb23rq0fUs76t8MG3y5QXP9Vz04/Y
yEwsHfmV6RMBt989zpx5u9BwKTNyrIY7kj5qhGFjCZFodx0JtVE9oa/xPdD3
Ghdkq919cbFNieQGlMUjRFoGekoP8A+8KSo66gLLDpcJIYoJeDGSNvjrsAFY
jS1Rj+2l6nwhpM2muHGxeBhua93ZYGgViPifiDdiOXUJuh0C8k0QL5ijiy10
vSan+D6klr3pGWDNblhsb/vijc6BylUnSEcHrzaEjamNy4rn88i8ClpPGtSr
6+KM+H8/c2Ky48Fo9tbVXy8LeRqPBkPl6QzlngJPIqzdCFMA94H9ppQNlj03
hPWt2jbxCCSUNUF40JredgpERA4jPFnVwHG7l04Jpa7WSYafqSgIbwYW0/Yz
J//bgNT+fcRE++69vGMphNqFDQNGH+yPuDVGeTqbfZl+uyH+kiFsjDVuURKY
Vkw5KaUP6TqYID/00yeJa9Y+MlHuvq/0+TWf98dYEYCK64jeygZzjkSzyqLM
rcx0CU7jiBfibvculzE+9Pa2mOIjWy38fHSWSXf95t5u737CbBxLfXAamLtU
3Ple3mHbAkMgu8vR6tfLREbPB3Ri26GQbWlo18r0k7gYBRF/SxXI/XJ9yxKf
fxrn2YKTkQHNPXpsHFWpFnFYZN0remdUYOhyCs12Mh5sAZSt96dakSQLkKUq
1Ps1ALWupXg95HlyDB8bOSzhrDemTonZWEccyx9I0HEyeHiwq6e9iwrBxASL
pv0SYZ26fjHrAa7a+Mf8idx37psgKi3PRkBLm4bU4gqA0OpYuHWwvpQQEIiY
ewfjsqQjEJ4R7BmZ91JUnLqCwqaM2xe/zgubZFB24u7fVUbExk7G7uAOA21C
kFJ+nHwjWNb23+T8hIPmhb3m1PTO7a+hQ/KBzR55aMc1t5JKjvkbfdCLZKuz
s/if36rkhnxLFl31drcpaLJjS5XtUap3BMGeDkmCGE65qT0DOPBSMt+6d+hC
jJ6g3pcAFGnqbu7mJG3C2/+o3D1wxws5qcKh4UwA4Y9uauPTMl/RDmnZpoRB
vrDpxTp/p1w17xoC/eHAGumCFXIatVdOxlKC/ZfpLhyKbI8UgpEhVeeUr4lb
GwRqBpcvF2PSd79XpAdg3F3EOY09pZqSolWqXNSXCEEaMNqIgRgsgjFYzMX4
NisfgamLFrkl1XKFi8tZVnTFlAGyYUzCs/wHZQWKR4rBpUOdMUlVuBJLa8ge
dplWPD0Vsr+wnaxuYCXp1cb7q9BzZIOWfM3/RyHiwpPnGXi4P7Wd7bFz3ZNf
mE+s1syfjc4XRW+gBjk/uqs90SEg4A3Bi8Zi/j6+aYeZe5ozscr7stFwzEA0
J2zGCCMJMe3NX1r424lG3UYpCaYE1jHJCS9sUWKNmM6kIqweIvYqHOmySGU1
C7KdXabznKefnG4sdMaQZGgvoFx2XmcON3XF+5sJpXuMIJKvjLayCqnw3oqf
HqXHGsWcXD8srWm5m0BxM+1oz0s0iGSwxJztOhCd3DvhJrEWySzz1e7BP4M0
uo28xw4C8LvTlkrOUCUZPEjv52QVla5U9KpCN6OrdwAuYUYC7ebBwNZJhsib
m3IgPiMXpHjfdcbISgXPc8yBXY2ySSNHGRxWjJnuochXqiFQx5+z2SHaCxE8
W7GIM/iqI5JBka0b2OmYt8aoHddxlnfEbgML0F+4xuD70cWRApkqgU2MmPB1
u3ToliEuUOvOET/N11V3pBNGR8PWEyWDD2D2ozlqNT/CLSzSHiaNXMnAUKvK
TPS53p6NJLTjk8MG1Lv3HwGUdxPQKH50g56xJAaAMgMzpLwLtaEHZeDzN5L8
OBferrOQjzAXiyHPLt9k3ssx2ZWjcwhM9ur1cqOt3w4X/lnQ9CVlFGF6YUOg
elkxP1TVWMoShbmIoFGC8/jOOTJvCqu5A4B9VgNrQtO8Mx5k2nHK2DUqblUS
20QLmgm/wW5Ww7xBA2QPQPSa41ToQK1KXLSl3nnnn8fJ1aUJ50dXjclsh8mC
yuEMrOTqfBY+5/ta64H9PHE8o51cVLYqia+BiiEJisuqxY8wRjWtK3I31Wff
m8im3mia+5sE8ZKP/TU5Qwxz8J+isX9MIHNoQlMVQ1+hw2Ezx5fe5qLvG2Fa
IvqQ3yXd4rUuBaFXF41WbDaNaXSPFAgXwrRmCRJpYNw8PaaoxlPxV0W4kTq/
W6Y0vcO+IXcNax/gwUKcCf3W3fJzuYIYaCzzK5HXA23pk8vsKcZwcJbShetO
2ayQkjqoV1XRpu97ozOCRojQ+i261GXVl8EnDtJOYtdJMasS2A1hmdP2n0Wb
UferE75M/Aip08rLlyfHrNSgO/ZSgNb0wL6IEKQ4O/6EK8yfBTtmvAveRbtJ
HsL760unOAGuCq7tGgkKbkw/Xfb4byKYzjjagIqoJEdE3UeEWnAtOSn97jRT
cFF5QLku6dckBloeizDxQo0XiJmcQ1wgAhXFPb9hDWvo+5Qe5ZQnjFX8/dSG
BktVZWUh5BNqMdrCux06m3VwVUDluwH+Sjhs4DDIEihWc16VOMCD5L51k2Id
E58KvQRBy+MsAn5dbzNsf9ivUDiWXkiMsxL3Wkjhgu8hVuqB1R5rpQjk9n09
hmKIrF6zUWejfdE/fhzGnu7I0vJriPl3zJnhrwFXoRNzQ3kWdJeuhE5QsHt+
8EKu4d0tioMjkEwd/K9JQqXZj/Cf9UAu1cLe5bRYSLgB1+2A1XPo015YeY8J
LNq5ChgKbii73ToKm422a8FYq0WrQ1fGVusO+fSd9lr5HVqlOUs+gx1zWbuo
WtKGjRLVQe5SlOsvO2js1Rns7mfV446iAcFL7NfAtUedIi72cebj9Wam/jCJ
UIgdd59yd8ckwQjOb7FhvAWtBa7MUyb4BC23Ep3alHRg9pI80pUqyIPMCVje
Q0RNfbOMH4rmDKLrb96HWh+TNfBiIQ6bYMdHn1bok8YhijRnh0oFZGTaE0Qp
xgUMB083t/tVSMh+poqCZT+3tJlsgCDhmoB0yJCqr4RmqZeYHsJgqedK3fft
QnvqgH1fw8gTxVfyRy/WgZUrfiFRCuKJCgL8vo9VHMKGtj+x6g/d6UiSMfG7
LUeJfpE2TndMdWfEEbY4rD4+S/6l65AZfI+YYPGqCtwPeXmEEaumN3DecgCX
8rf03G2HN7Pz+y4QQXJzuAYQScS/ERvXFYV7iRQ8EGBwMOoP5gdj1WaZKBj/
Xr6QmXCc9DYz01U93Pj/vRSvJp3FySF6WPsm8P7Ir+GqKpEL2JwLcyBAibuI
rC3ESQ6lXYc2goo0bZnB46Q7i7aMTF44Y792+uRNg42KvcBWiIpxauxmfvKX
vRpEbnK+7YC5QB1PPJSQVbnQgfwWzxvfdjjt3h3QtYU9s7cfM/oRf2Y0VvmP
2NPMRUZlS8Nm7+m3I7f8Wr9vxxPCMaw4YMPLo1VUtGoaFNypgWphsnwKiu1k
qbwr1Hf2Jsash/jAi/sE86kRe97KvwHYajWJQl+Jnh0nleQBEc5mU6glXMdL
xlIPVX86dtqmDPemO0ltii8pvC0yreYjQ7c29XIIgG/tNPZhdTPHc3Bl9uWe
HTScGGQz8fbS8hz4dQVuGd+5Z2sQ5JxRJnhQcwver+Wyxubp1Ra/dIMGLAul
zexYmw88uXiUCb9pCBl6uo4s7Q8dh1nI/bBsLi9aQICE00+eWtghwpwk8q35
1cS/1Z0xFMAY1ipp2TEV9ChszR0K+1zI1/tWQP40mTXCBYmxVulqaQanMDrw
Sq0Zq9BkwIC9RWTC1VggTGygdhp+TlexIDU1Rf+R6qWsj+mm9HM+qtWl3+cH
roE9dhMSDUPCyN1q6UF6yYXAS30tBR2D8Tqu4n3koLzvhdm2TboU8+cX2TUE
9M0/erYqETELMDWN1QWTHGCXUom/8o0CVsreKkOOAvnvQzp1FTYgzSWv67qv
rPtg9QQGrxZmMHJzqZ827UukTtWOGc3RFWJPq71UqDKWwu/J+MiKvugnnu40
6qzcPKezyJ8M2mksWsY6TTbuTLun+Wu3ZCHvlnuOSJ+eSDU5oqlLqFya20mJ
SSlft/pUjb5Y3OngH54uXlkGtBIG3lOyFVrKi3keuPIErZxivtT/x8Te7LOy
xeu2uIKENX/Z3feQxPW2Jh1h4goE8Ae64xWsegvESFMvATzHNsktEmw1134R
V/8rV1TtbBd22+CgrfKr+iTY4rliZRWyuSLnRgcwXB6YpHoCAylDS0aJjd7S
2hwh0q6hvNWP9Hgf+OR2Alz/rtmpphEabG8glhJyFe0lJi2lq8MqVWiEreKr
gVvTeVuhOVbC4teKlhpNWG88oS9LchbhL0asvI8XF+uT7l6shpELCkbAK/tL
f1nLI+Cy1m99e4sWWcpFfMTc+KVTG/LdqwHtZo8vf16AvYrg9ydVh7K3K60f
NepRADTdUamTp4KrgKbI75I8k+K9aMKUYh9HmwewQ/KDxkucHORP7qQmHJKc
Qsw0JUWjMsUlqU2j/pV5uTecuePQUfPuUU0j0DF8xkHPobzm7A2BqRcx8gtG
2dRf5SCmDbugv1TqGy+M/7qYxjtQOaRM3MWA9QqNec9gww1MwkBhGepsfz6+
VRjlNm7vY36U6eb4Ikyb8VkZuuaaoCB6X4W4k1EgxDKs0zw92CB+AsxotLIR
UvGb83t3TNBUBJLbUzjdyRduaSroe04w+DRbwG93Z9EZbcN6uUfmlp8Kblxm
Ec0wzsJuoIXEPq8YoJIzMzwLpjp2JsA+4e/dXf7W1f22JaU/hVarDn+rLfpx
XolkR0AcAAn4l2aSm0YkLV0HaSQ7rjb96lSnspAWLObBO4GYJ1jCfg9Qw/QI
/I3feh52NEJwP3cP0eex6tSK0blEKB8HgkxlRHFr3UsRHnk8hs0tKUwUoX5y
3qKe6N29O2XNuX0k8YG0UhXF5CBKZqp5SMiT9WUXpQGqkhoA839fj4gk8Tj6
x42dYpfliv8Njnebffeo40+Ey4C84InsVcqPzW4mSaDZ0hV3XIk+EJQSGh0k
AjfNGuagEDgz5BECNvxQnqZImxH/c0YwOW6uLnrAvoP52QjYJwv0xM7XC+Sm
eA7MYmSpt7EwXJnezLq7ZAF39CFYAmlC9ygmgbi2+JH4GRIC0Bmr6Q7cvI5V
wzi3RFpCCE0Q3RW4ltl0tJ1Y+JF/nNrwZzfjMP4ZrLLvC2HEIGQj8c/76IsE
Qy0BLtPIFZK0N2aGML5wxPMog4VD1iXedweDTTEW/nPdQPFL2AXc1MIhKLlJ
14idyNebtJIRD/e6LbE4YUHdV1TQKeyVYIo7+lLjTVxiI2D+LXnyKKZqLPUm
PH0kkbrGg4xWxxB9NXYPM6hvF3VDKloaaREny3cycTCcnn47lyWPNqG0/AKm
USssVndEEzr0WA3V5bOjK5IuBfkMxrnswpftRwSpwNf/Gd7LLbCaf/8WVb9Y
Gl1p/XGt9kady9iyD961RajzHRCyoiCfs5PjRsIhGk5GimNamQL04tNIN8gB
thu/ZzVFvobwgOutx2ZtWsDuz4nc6E3aFrLh+WxVbtotBVnMPyAexhmk1yaH
bavnzyNEI3BuYNamQJmU8Zpoif0eYfW9DP+SvzPRiGQKkEZRfOpLBK5tGck0
w/jA2wGVll/jykWDuxfG3LZOTL0Ze6lmtiAkU/iy/5pm3S6LiBk186CbSBGc
c4Wg3PqwCz18zMrVt0ym/R3fawGu+/YhKSbsoKaow5sqCL+2Y6bdGEJRZ7Lh
fy3j4G1xfriYePPi7l4Pq0MAikbJ41AlEO4ZspgarNh+Y5ucWGxcmCdLxrVI
FoU3vSOeFxoNzppDS1VwO34A6HXlttWqojv/sMS5hEv0y36vLyXmaxCnYyc1
JlXrO8zkKqSTz7nUMXaubTX+xA0dMaAvZYeFIOeHJs4eGH/BcrmxPPrtwIVS
53wpX2fxh6O4IK7Lfkp41VtLCmU4ehHxZOpEN5m8KCjFsYPBM33xweA4xylL
E1XBAMcdNlo/Ngv/vA+rwZV1N5q79ctcgRexg1aw7Dg0MyjZiDk+VfZvGaUD
161+sCsnKkiKzxjMVFo+bgUQafVD7X9YGe0NDwhlgPc8ELqVqX6nBQ4A83oS
mpJ2TcEuXVUdXF1qzLMAkutYs1GpI5QBehkld4atMFmeEU1zxbqSuZChsHbf
UG+A79K1/uL3f63mE4u/seSIDzfxtp1EE8b/wTXudXLRHSx43TIWwBHbMiJN
Raln/pTTpDDiZPivxFj/rAUof+XHCKvkndl5UgEl4bRQVRx9EefFQojWvRxG
5Hp/+KGLeEvNdSGqeRDGSXNFVnOb+qNAVEsbWmCdjHPaYX59cIAS6x+F5CHw
3ph7mgLcreDf1G339dYeI6nEd4MAxntJ7VnAA4aaTrpen6AcUfKZ+MCkw3q6
MC+gJ7UjALCQjdpelV2ZYWAHkvikJfgM6jQ+F3LCKWmEZdYp29QhQQ536eQf
wDYjyyhMWliBrtsCk85BnaaCA6pipNRNdvmTexhlM6DTUBHjdHbOOGbJdm3b
IHvtiWrsc4W6KbwKIW01KuHjhWiAlodPrwTwcjzcgTmjxANhZnd9BSS27/Ci
Zrbt9DrBKa9Qk5j5XU9GFxS01PvFIyDX14hO4n0P3tznYkmLlxklid1iJstC
kx+v16MOITAF9wvcarasPiC8guorv1NptN45swUaFEJxuQl5/C+3nT5rFXH1
XIF20n3/SOniADujd7PSUb1w4E7wkGbbvdAitOpCeDnKOoIFEbVZJD+GUSlU
S4dsuUBLzhxdz6Bc+fKxt2yfAqDDcMPbkIUlYu5NoqubkP3awoEQ256mZ/jl
lL5OQsKymHuq7sGoNRBbehmcvulvmzVl5erbrFbVBSCevc9SsLK4RweoAojA
M9lrrX8RwhRD3rH7YvSdTr/hwGnwINyANEDsjZJKUp4CS7YdWFUOXqLkop1z
GO0/0JZMBxmKoxkEs15Us17VQ1j7Li7go1JNNL3/x+pW7EJOZRyY2ijzRV6c
etCI34oRMkzu5LG+Q8Zm1qyPSF6VfnDa2fab8/aLUMQs9CxsjhtmFlQuA6lu
XuwcIAYo4a02qRlS7fbqZI9KEqFXbpU5PhlDFIip5aH2ieomiNEFbucOGz4p
T0h1lY+oB8Nhgiv51dIh61GW45vlVnT93osrwsj9GcPap9hJXl+PkC11R7F8
WwinJkurwGPbHWvYjMdO1DHz56mt8Qrz69a+y6ChHNQMEKOCUgH5PcEXJKGq
EnmTgeIptWYqGGcn9vq3pNPJFIcHL9SpC1vKiwpuSwlup7E+G02ZokF+CH7t
oClch+zy0J78UP8KFJY+2/IvVUdF/oRFchiijVWWLIyE37ofSj5j2dSQx22P
NpaoVbYhdMK1x1QDtC3F8CaZfrs/kMV475ifawnvM2RtxXd06NqIRyphvr10
2Czmw6ML1NlTcy3Vv/f8HfJx0XMObNT7NlXh/o6WI7rI0vwSI2LcW1WBep4T
G0nuZ9YhFcJD2zJ/VnUqy76IBovY/kdZTE51qpeX2VEciSRGIydoJ/YDG3Qm
QUAGRBXqV+5/vJrY9raKE+rgnZdOXvW1g0+OjvEEgAH7J/TRNY1gM2TkdUiB
5NvfQY/+lZJLLCyEBe7GYqIYUqmF/Jmx+J3WMH18mebbYDudRwii+UmebEES
eKPYfrrFrizJddBWqEwArJyeH8MzrjxxJkRe0iX+yzyt9TfS74Fmcu28FP2+
mHGLxkLCDq42WBmExf79M0AUlniv6/H0aX0+guBO0q4TI4cVhEMHLeMgJmmT
anhyPNr4skHlM0UqmfZMJ/iuvsHpXbcPlJcm50/0e0RfS/WKrOFcHWMMMjWi
IOo8eCx+7tg/9uU83G1RPJBxTwXlpvF/G82OpbobngkNOWoMYm6TJhVTdkXB
ugRZN+SW2aU0oTaTU1hiCadNmYKjPKgVNh5YLV+T5hlAasKteIQ8N3E8t5QE
FBs7l6XhjBLcA7FQ6aaaeHoGywmRCCTybPq55o3A7j5VHafMfSu4enVXz82R
FR278XLtkSGCv8pUSVtckPr7AqXvP1BP70IOys8vvr+y0etNjlTQJ2z2ktLM
ADejNhnNqouI3+x8UOUkhs5WwMjI11UKgFuhCX0iIOwD/d5ygsHIKguvJjwU
FCKbv1xr8d2vEovbl7znspyC1v17k3BaZKs54mmiQetWD4cq/W0leLWGb26C
wYpPIwFArUsnnrLgjMPZ+ovujgZ25i+TPwq0DUGXPhwm70oax9IdZVvJLmzU
20/xOrvrwKVC2w6kk0K56naUZm8kqIGXb16mUhtV3vJMBQ4J7IbTi2GmsOr3
J4ckLKFFofOnJXBC7rVNgw1rdQq79OwPddUuvvWONN1AgHjiXpt7Lbjatanr
GitUQlVpV/Q5+J6zAgDr8sMiO8NVxtdZbFbu/iCQiKAkXiuCBrY8Jw8J2VPv
JTKwfJ8ZRFSqsWSthKqvGmxpWkKFl8gk4gm5obxDAOUMErlC4AuzYwIuQBz7
92u1eyPUM6Bl3dhczl5jAi+PE0Kkr0rbSOxzklcVLiQXG5ugC19t6g8PXviH
9PWLEqXXqn2aqJIO2XEyupr8uIjHJDrjGZHZfQv5TTWCVQd+ydI9jazGPiAM
KpsAPpinYo3GQuiihR1PFuthbqnxMUeAEVAGI8ml5Fq8c/I279advyxO2h52
LIcE1z7w+OktBYzklIS/0IyNBu4qH1hq2yG9nagdlvApEjA5s0LkV/wfdEle
wKTiQtrA0Slo2KLKvI8Iqph1hdSaIVFOGkGKHnjMCIS4Q+auHi9kFCkv+/sB
9lp2p3uzZVKuFP/LJX/6In3bEJpVrsHvdIsqoqJO8GbOngIwVt7wcFITCbnA
10L1AafKN93LQ5UbrjJeXwV40CH3ajJW0qy5BLS8WtrrZMfZ57y4/+dqOa8k
EiofN+dGELeij3rjb6p2N9DioUTrI5dqTw4pVCMl+KTBA0/zJQhykCgpxCso
SAevOHN+029YtsZRp7go/vQwumFaDAEuc0MatVjGsE1ByYziQ1iK0uOwdohX
eCauXA3dYrPnqD1hmVqzrthz3i1ZFR1Kibh5ZqowZCu+/B34HKd2lsxGZfRV
0HtqDjk3GYmXH0/7ZzgE6KxAZPF6i6UWDkAk/6YGjTFMAGNOIyPMlJe/dWxw
/jmUEKocruAY2H2u5cl4DT6bj035gpwjbfa25WXqnLxxZ8pHJcvoBAo/8COk
A7R5Wiw7uWBaNFXi7Bv/e+qRw3fCO4qWZHolaL3sDxct5idjZ+hSQWZ0Ih+e
0Zit0854Z7P9t4dNjgPT8HzrdKHXub7o0gC3F84ygqteRap6kgIrGvoewcma
eyZqcA+AZuptBGjHTnAV6bLiCnvYl67jJrHZSLP5LcV/5CvV67MWjQmLhGUq
Z9FHWTXOUbUuqeb7wR+iszfmLJ+eY1VlWA7nEE4rmgKdwwensVS9St9+C9CX
rZYIcoXVeQO1yNC4UB0qxGtOeoSO7dyrbyJBHwhpHmjzOmkG1R2UXFG9P6hk
4ojLWlRGag+iSR4onwK9llg/smjijax7by5iCOBujK71JtwrJBpH9r3JZUYT
/bW9e85muFKipJuhk03ej/CWih3xViGWUi9w12IXYxHRuTBpkpEUcMhm6VKY
9SRfGH2whyTnrh2bz48Et6u6fE792JdsFiNmaDPV3w/apD/mtJ1njmLK9SPb
dFE4KgKjGpRqaPIaCG5JXfOUprMmT9kDDmEnx1gayfpsiZGni+NykxHhBcQF
aVjAUJ+FVk/32FULa4Yr3KSHCZzoab0zBVsWfLvJ8+3ARdAWe4nhKmzP0YkX
E7IL/yxQAumoL92VhlG1Tq1NwQwd7Y3YcvgtEzvbdP8jlVZ8GuIp7ytMVL8b
IxTdBiDpQCwyaiYDd9NfT7lMSsC04KPONe42pqImCf7EYkYpPSQriiqatzGA
f/rRrXRd902AMNMxYl4aopaDQb3J+peWdCV9qQ4bMB5705/tpj6Tna8/gjWZ
am3cdC0YTOxCSzkHP8fkohCs7v5GLw54M4L1RZV0YA9O39QHZy9LkGeI71vl
05oPzJPufdIKpZE2eZxHMgp5Y8Q0cEQq2GltHSoP23LMR7xfqntQMeTxI77Y
699XJdIF2EuyD9ilSW1m8bMuFx7w1VY6LjAC3vP9UOrfK7T5A6ndY5wuga+W
fX1MyFr7mkOnYcyFS1LFaJfi0hpEaaGcHUgP8lWWeAIu91OSpl54xUFWItxS
3Z3RIf5TEL70E5mExJB6UIDYeQ/HwbqL4RR+gO7WeQ8yGQudmb+xgdr7SBdN
fQtIaZawOm+/YDP8TpaNhu73l3veDWIniHhRp4FQHpbreo/k5IJiQtGHEjNp
F5mmgJEX85cWNzwraP/9olw70z/0WOlbXBbIcNGuYlf1FM6UdCsnhVhZt/kJ
ADfEJDkxNzw2RQqIJZ4gCrgH6EKUz7h7v7BdCQ/cPpuPgTtIDdKl8PGzQ79U
Jqkeep6UMJDoW1CzkaXlaAtotrU2SNTDtDYQuPI6GT4+cJ8Epe2hDWhT8D3+
QWNK7VKWZuw3ulL2yn6plD+iaXi7rGWso1dbLVVMDyNmb9VDa+88de/Oe12o
YF5bcnp2EKjdtXFX9F/8CckUBx3vzuWr6Unfd6uMUpuruFk01opxaqFkYzJi
4ABFp0L3Y5Zim/0wvixbAGrMR59koDX+FCXAq6wAhupi8AJV8as92ANxbKyB
fjLOcah6Y+STgejJv6vbBdFtARVdE2iGvFxG7vDG5xuyZX6UxtkHxmIsS5n2
eI0aqyHSiEjFlGRCgfZ0VNFkg8vZu7mnTJbE7CCoxskGWAfHz69Rd1shBvKC
v6kur4UL5eD7YUiTmqKgCJN+eS9ABYmUwhCXir5qpC7FBUORelgrJajSp4B5
v3skCyq+lBcrEqWoS/x2VXBGF+z0ARaP6r8CZJuA8Ce21DL/bXxgaFbTQkkw
nDGGCQ4290skh6NdZKozxtjEz7A/iAaVHgs9qtP2neFtlMePzmr4Ap+FKPuh
OlbdcBSxLTQwPyKfVqs1gntmJtZEoZwv+WImVCBPnh/qclInpX0zV0tU4gkP
mtp7/RD5Yg6sakcUuLZXP5CWNj9zUphZJpziDpAUtAC+i9UnrIbDUg9uS4Ti
D0VqaSgvVWLV/HVKs2PZkQNuirMaxiWW137UlboJtV8sCZ7GMGST+KhZ7tif
Q3EMv2MMerFBlR/6p+yTTIFe2JxLN8Eu+VxDgucvM4gw0YcvC0gM2WEyU43T
c4iDj/El3K4FjboAU/Te6eZLKVkyh9j4SAhmnaLLfkwtQsvNfQcHkm/Eks0k
gSlMAvlp9leRFiLPIFdepLQ9jYAPJMmRNpY1pTrXEkSiCedG4boS1EUjy5Lt
7h7QKKam82tuoRXsFKYTTSvDLBSkQffMhvr+cmLApJB8Y83ckXlg8CWmBZoL
yAhG2kNhrckL/UwS17KiYzBsIE+wHBVQvzkkxg8AF9DcKK9l6U/L9Kc2+HRN
qiAUpXBT5YXBepROozx3bkemY6dGQjQ6xo4S13GQVW36g7dcN48bfDTAm3JK
es+RHP9mefJpcsMeoVRWGF9KRH+tSufcUBieA82pFv4xuJ6FTLNbUgNO6nih
WZx7fuINSz1h6r4bjqXMzHQDs2O7pc3PKWfkANCLXAW8xvLN30n6aOgpQgUR
pMWjIZF9ERKeWlqWQ/VsvDYFxk2diaErBPYlkXqT4L3FIPLkXQmlxaOY8OAh
rEn0jx/E0Jbgy2X9JEXcn4XwzJAtoGASYPoY99LIR1RWbCEt/9xSAfdK0/Kd
NDtw/CbdV5/0bB4VSzCFADltvDuDKqusVfMxMfB9wDIf2FN9AmS5OXmuFy7U
a+lPxBAgZ2AO8xRvCVuW6cwvV6QiyJPErNBKv45Xz5SsXkhqGlRVY7XuZNuc
TzatG1b+6Kk+SwUuYblW7lGuWC9VA5e2M5z5mb0wHy6LH8pme2c5HOAau1sa
LTFWQdeg0W9YvNWxrX5x3BQ0wFpgV4a2hIVpKQ74n3DIsx8PjoBJW2MUGhC6
8Q6LuEAlQdf96nLVQKhr62zrl3JVJTh6jD63n/sL+JrLr8iN9d0VP7h9orBw
qcoWRviXoCLVqGd5NOy+hISz2U+JVZijk5Sz4Kr9AlYwulMr6z2f0By8Rs1a
e3Uc/OnJEAFzQOA5vvUZ2Wrejp5o1+jrBfKMTleraL/vIEp3nt+KB9TkUaCz
/XycY3TkgxKnZ6HAb8IIgllfNJT/phuGAc2deb/OQLYo2+KrdssHD4EZbe+a
n8KeG4ulT+snME2u3oLKABl0Hu8DWkL32cORK5t3FivwxL4P+eJkEo87rUfU
JLVEi2S6lQpxtwYgEVRQrdyzPfVN1n/9TSX8cuuLPO6hbtX/8ifTmgiMEZTq
pUAq3j6sbwTDYmDvLCaRqza7xqBRgfwZfEB5Ejy4U223/FSZG7dLFrHSYrFB
NNyJBFCK6cCM+6ymJeBJpbyr05KFRfsStJS/ig5v6KFNTlg8prpAR1XUkQgv
l5VFT8n0mv3p+5jJGPpjmdv/U4DzURBDtlDZ+7Abyy6zyhztjHGDnXGnpu17
7ngIa9cB/wQ299TDa9FUhYnjeI342YoIgjdWa27Exlnsmmqd9bPbmEcW5OFu
SZ7f57eAn/dESFSp5hIayInhPGSDh6r3VewwPl2XjB780pc2Wt6mmNZJC6Gn
iNe0LKhYoov6PohFtvnI9Sl888jguSO1KTydx3ssBIwNkTXmnialp/JoQty4
Yo55szv2at7J1B7ZPCPFf5T9nVK8dPuTGTI+GlzAA99/TRGcF1xuKOZ9Gz9c
3zIM9gVTXfVAWgKE6j5Gwd7f6CK6HBGI5CxNEC7x92s+hYJvxPoAjY6gwKKJ
OBCyML++ItmArKJgylkzXYexxVRVr/ey0u1MiG+Lua4srx8tlrsQ1j8lrNF0
LCoc4tW/2B0WLgGwDg3fK3N3AFhzL9h7Y62ycwuHfqnpKMit2SZNo5DBhUs5
5RH1Y1BuWEZolcRCUY7LKq/ux9DVfPice0tDJJ2KKzPNkfiOEJuqaoq6zU7z
UIiyjoMVP5rfyBYw/H+k28YSqe8c6Dsm366wwaEpuGr8PeaCa9cycCgKnhh3
6Rn19rLOdcRAXsqNspMm6oQXPmRCo4si3uaVFaM4/ikiIqBaFoncz0P2JXwj
DR1uUxErxN6sx4smeL+i/I5mIn9XGOqzbXxTILwGBTLtS8pmToI+8Yw3orF7
3LdUbGjKxznpnu+MUGIRlilzs2bqZrKyjll/J9tet5ZbiuCGpukCvX7foJL0
2HpiG/yyZJfk6xmK+wtNwQqLngIW2fky78WTIYxb/3TZkqDdBlDXj8afK80u
ZkP68wUfWIEJ7j0McIRA9T7rACGwxX1ENgFkDveL93A4TtmNt4VlxpvWYDUx
3qKM06prtx9FIzuiNnhai4E/aU605Mn7YIKiKjGMPxRtI0UjB7ukwHJew8a/
YYDkScj6GDHwapIA/pfKhAKdQ9u2HxWMxUZe/Opu7y2wppxK59g5mAA3ELRS
2bIWGKidpmRRtljk9U9eA9rUNzcLjMi0MvoS6+kP89RkyiEpX4duy5Sq6EoK
uxcDcL5g7jsZ5zOdFsdErxD62QO6vpkGyms/Z7/BwS/ANDHac6322WSq+bnE
1KDs/Vf3ltJWpgPiTmRTLQd3IXIEw2qmuclQMz2KdSb+/hPkFXH9wcpgX4LW
ZvwaucQZ7ziwIx/BdbYKbBBUHpnvuGLcjee3iqjjQwE/S4EIX+F+K8Zb/ytO
Pmo/vjhVKwD+aVs6H1jnFzuztKeROJwgkFvzzDsd0C3xN+v/6tsXTuIYW80i
RpCJw9kSFWe1T8kpzd0wwJ3z/d4FdhvAsoSAbA2gTGbmPwN/2na9jB7xzidw
pNnJs4fylxVFAmV4AROLMV+ZZddBzj6H5TWvERczdALoS5hEtok00JwYuhwh
lT2mLz6PYIAKctc/OphVQzh34XgeT+QQ/ahjiD2Bm6J5jcavsDlIuumtxr7s
pgQjIrM0LTmTqdHiy2B547bd3Yn2yPjbrFrBKQh2LNYLQXBTfW22bsJH16MN
aLxAb+VzhcCZvJ2ns6pzBWV2QhhgvZhxBYRSZGnm4QXR4kyD9y4RoDbOLl+7
Co4WLSR3Lzi4zl1g70whM/KD4BSFmblQGXtxYpzouWSAZiIeQqC92yZoOhdP
iMqHa5PgH/iD+QgKx5pM5Pma1kXQQF1BJR7RALk5QBR21Htcbru5MZCdgQZm
J2/BpBW5TIlVepYdEMRLLgpT+w+IiYMeU6bymdh73Iv7ZUhzKKf8bftJ3Qmu
nTQ63XR3gH62HVpAwX08rVTLI7jd1PXyKE/MrZrOLzXuhIUJsom20ocKzNV8
m4K9FmKRr1rB4tkMTwxDD4wP5fFY5HhjNdugum3jfXAIqUtQ6MXxjSi3A2vU
q4oY8Ad32DBaUNv/ihHHxOi04EV3BMXmiMyBy8/Ww4zhG3BzpzYENmvl+4Ys
FE7cnBFVkhvrUUfo/EHzhLP0VjnkK5vkuPcmWknKDDDv45t3p92suf1z+HUd
d4gwC6pJYvSdAWCPmMByxJTfNk5VcJsvh5NazBdIToy5Q2zWz4dgm/tadufx
BJhFOPeZgf+KyKFFQjqO+QGm0wiJgyVNBBOiHzSrzdAIuBdXI/37CRTr29eA
nBYuxIdZ11j7tiTLzyJpKUGSsyU/ocL80XkOY7hWHwQhAWyarrMO587jRSel
1DlMCTFg7nHcJcrCRn5v1e3Z/z2/42RSZtdsVwbD+PEqzX58aC0cjsOzOSPP
MduMHpwHWrRRktAmB7WHAbe1ytOIex+f2+GiowL5XJ3+al2Z1qwP4Y9ao5WU
T/KZaEdhimrHNWeShQ7o/Keiqn3ULm88BX7AFS5H1AA/bM+sKlfy+egXhrk5
9+6kOCebLIP9IfrgCCyePDtYMyMsA30UcGK6iQcudEvBecxaekQ1fb+fciVD
+PuBWfBJO3PbCWFBPoDe6JuAIM5srBr0se66sfqkH8nOxjbNvGsm1h1g0Luy
9yZZs5usbbpc2RbCiT5DM+KEJUxSu40xNUV1CzhcANUEYzWDqJqP0RCZZ6Xo
X8OH4wketnqi6YBUDXWTfoSH7sKYsxAS/FruoAebC0zzTsI5/NCRE+Wcc0Vo
XICqmyDhs0N8Bg6Q6sSu80b78lFgTMTbuZmjzSkkAkcO/oxN8OGSzo73n+KR
3FLvRQP8dxzqDEaPmZVWSwp2RovQbcSFUFAv1ZwG6v2TTSI84OF+/JCCSC5t
wif9mjh9n8SKA6kf7b6yg/lb62ga7woI1wE2kBr78O9jUm6CKceiwe07amDY
8nMY1IlzsRnltzMhjPKOEsCdFMZuS3fJ8y1uQhH35NP3aPRFi8C0ozmq2r0T
s8gpp8SyXrOMaUzMZuvr/6Nj1HdvAjo5C8lQsZg3xteWVQwe7o8uOsxm0x+Q
y02txb36rcVX0kLJoFs4802nktZGUpfttuWa8pl7MjdxocELNz2oEPz71B5r
jcPenRl0QJV/GzobXsf7tk0uDgMDzhXdhw+omJGFrjMWXs3DkIV6jOV8fzGc
/9OlcTuJvUC2yS6L5s12peMKNbdtpQUZ1+OtGMabE43MkgiJwqA/HQzeAwmi
L0VZSqnxslxA0na+QdWoqAvoiMtyd7yG3oluCeGDGdTNeWjZFkNuhHXbRSWH
yxBRHNmyF8Mgeu1fXMoHpbyXFLFeLsc3DOx15AfUaNtR90cak9aGC8dxWtEf
w662V38tpYYd0A2k58HsIt1Y8smk4qroZfiiChoAHPeLtskf1ZOkkZQWkNtj
J9zYHDrAng7Sk5mZbyCoZuXDsVAHP+gx6yrYRqMtzy/AWc0KE4heDEFj/oR2
yovCtll1c5vV2IFWlrMOmgu6P0YE8GCxFIJU7XRNttcgnvvo7IeCJuajqNnI
P1MqjqmXFceUav5sHNf24siqYuuwfdpIStSO2UVO6+C74krydal42iZK7iHP
xIRyu8h9hhzI7w8zDDAM67GPgxe1wF0PE/mMdYepSg7UnOckaoz3We3fjg8K
Z6wgNsIqj8+D9o6/13cPTHgfz2ZRQrxR4QUEtTHTl/B/WKQQjFcpmwfpbIe7
kfSu4TyJnwuEPiIO8m6HU1Jgwwn8sEQlOHQUiJuUUa9LikULcWKSRkiVJgjn
igp1qhDSwp1Et6WsnoRFrPpQon3yIfHLBZ1aFlTlzUCPlt99tCsIg9otKOXY
/MNtmAGsvYBdSZ5JQovvcwueOWxdn/RQaGOrB6qOnAaGnIR3uPGHWlJ3fe1F
0V8TXnxomzQKSVTAvmttkF/x1hUEtUrosV3bFWobEA9aJPwWQ1pbfzs8R9rl
gEDGfyJlqOvslsY+gXPwkHm3eTXxjAMopf067E8As8WcG/GSXEkrABr7jqg1
InpPBCrlj7SDA0DQb7RGKWVqbcqGWwE3j9TF+kKpCDIMyFQsDTnT+JgKwNhc
HyAgrxXQlw0lMtktdHqfGWfoEfuzPAglgp3KSZZVj+QsHcSgG8btVrmwJtnW
NsRLK4Q/+dD3mmsK6VPKlZ3stbLNQECshIKxDxc2MpF8yuotjHBVfs0IzyFv
DfwkbWlHAiRkNlgPoubZedjCWzE+UWNKLr4cey/r7cOOi5yUByxybllpzn4e
uKSJquL1sXRYMQWSMucqCmf2/ueemwDjnrh9fob7ELJ5tky6KvuAJy2yuhNV
E28p8ijVn3ltdY5G3eSjaMaH8VmSAmAhRXOTPfWns4EX8auLp4leA43H2UG8
Z2+ovh0BJxUlskwkb4tUi6OENU2jGGHMHjMnjExyfIFOlOMv6UmAFMhp3qks
Dcv/tHHlgwnwqt2w67Q01bIahmKBTu3yuJiulTGCzMm+C02BWkH5AjeANt2d
O8b8eeVcD0vTgqMwY8Mjnh1YhVM5zWogpHcCX3+Bg0QMjjCO+9TQE3wNuM+U
RaWG5zqjPRL+LvDOYvzW/YqO8iHYSosAitwI/L6FbHLayD6ODmqNEK96P9nk
xn7ZFMvSBIns5/QoAAqW9mT5+edyBAL+uzMn1Hhirf9uWV7TX4DGIZlVsTj3
aBVqTcSk+U611KSyggx7Y5VmZ8VxmQmpOHkP+F+Y3uAT6QZdU5GOp9DqS67R
uDfWoVJToTGNatnDzd24AIhyG0l1pNbfHYeW6X3tBaEd4UPFeaIpCmxDkn57
UBGSv7+oUX04LHs43b0eaLqmBiimDHPOX69J6XKdZ+COtBde48L53m+ps4Cy
//7DKkdgUsr58F3V1CI3SIIj4UKa+Tl4dkQ73JF9tYG+fVhfd+iT+tTLa9vA
mrk50oOmYQ2Dn5sLyvoeFHW495hz6NWnxMttjUq/rPaafG8gjnf4EqEHfTnU
mjCho8l08t7oO+WhgcgUsmQ4g1pNX6FDA0N4TLHpAkDAuuyllONbKuQt7Qf/
LmmDskrQ0OyHjDoPybWPybs3uNSPU2cG6eosPNntLMsyjiKXIRA7Mi+Bv9h6
EchJHBSIWNKlxjB2ZrO+Vu08pSbe8oeGrPO7UXuzTMKAjpKcX5+xzhaJm3xv
I52bw2oZu+oXOwOcLEbqfhpb1Z2egdcRh8ZLnyohAk0r/3iNkMWzMO31scru
bOSWus9b5igFgsAyL8JD2HysFy96J/OYjB6CpPGCNfh30ByvIP4+b91N/D4Z
ZyLe1otkENiE1WZyaoaoD6DJmMcXs1Ii7Vd2zHcFAbQh2hLIZFSBQ106N3xw
GozOyn6hUsh6c0ChK9t6a5ER+KxmW51xkU+UE0BK54RjY1LLAVWaUqJN7ncD
PGTLQVmqFRX3rBYpoLMC0MXpvdv0sDASJRp8FdtTLrc9H8nF0ciBr3bPvjrN
pFTH2K8hlIC5AYiDfIirMkBQ1hAu4KIYJmSsKJcg0XtJ9KY4kz7vEkkh1+4s
GUn2M93L5bYLdIc2u8aynOxhJZQYAOm6biL/L9U2d290cmU0UL04aJ1uBs9M
b0Su7jk5WLmCC3VZe4mX5bK4Ka2xX3YqwxZyxZ3ct4xjfmUV33LCP3F/BKY7
Kij+NW+hejXyE5EXiHTNGwtjYNegY+JPRC9O5p1YXpT20ABNI59qp23g4wnc
D14tyaZPpYzBBywRX6XvZVLpKswAoiBw8HC3yiWdDSlZH5qdLakI9Bw+p9qX
3fMgeOx2sVb2/MbQHItT0fzJYeSKjvcaOoUdZhVx9RXJYIxnrMAdZiooSYez
NhRYxoik06UN0DXVxhKsEai0A60+iLiFDvEW6VZtHgm0pCFytiuWNdHFrtwP
cjV/q/c+eiZB28krm35noIUKo9/q3ODMJ5gx0TjrN/U4yGTZ3BgtQRJaPjKY
xo2pN6FIWLicDghQ7if0F0mBO+ViMo44E/gfERzI6V6uap8UPe5KNusMA4nn
7KJMfLyZ9euSIuNCGEF3hYdF0bEio0jXO4tGpXn5QemhtPHC13z0ExjCG69W
78d2tBMPp7zJRTgLkW1UVeBdlRhVXk35Nw8M2VE7XYOo/apfbR+NBwEjemzU
HzCuXyQ+FX8NXn8SZTpzOxQGoYzeL2cPeFgJwxqeUwhkfjYICnOOkp3t1B9m
33m9DKOtLOIsRraKbMAr1VlwWeK6LqwXqrnZoX9CGhbLIJ+Et5raOcBjnebA
KjVB37X9D68axu7Nt0YmJu053gIYXuGOiOv/5z+63MmJG9ZwkjqZHaLRVMz+
TX1sO+T7WItIhfeF/gjFu2wkHQkAkcqQII90WBtAEADZMD2iqUa7ojkBubFF
jEggS+AzKYN0b99+4+Lk8NhdZ3f1m3oGqQJze2SwQqgDYFCHdeodRMctYR/T
ezKHelGBfGSQ0Irh1apb2qrHu+S5xLigwIOPj1SZnU0sYiYqjFWnOR2PwPV2
OO6eSGzUHRkU7II3LO5XPBwHbuM0KCrGekHoPwTqDAAckutt+Jg9j0nT2A3x
/sb+vy837x8+ZofNyB/q1Aslj8Nbuw2YKeHvQTUl/FfpNs7rL6Q4iUOXP9FW
R8InYS/O2ngkRenfXyqTpfd7CplR8gesDC/dD1gYHq1PXXgYAgY+eDHSlLew
YMocsxcR3X/ayg2O4n4qt78T50PUQsTvFvICGvv7zC+5FeK1GLGNbbLuQmIP
roA7p9xUKFbfWYDajJ8UZG2N1SwZOxg0MwwkzCjGVrCp2CjmJvZ2RjiZvrwf
5rdA3m7TMWKcpUd8CuyDfd1WbWQl1WKslY6tKZExumdqWpWHWH4GG9PFEK/v
TzHDRbggmbdJbxHw3B8Vvlvh0qqI8gdYgdF1q6eQnL7yoFe3hTerkcB8iJnC
Etb37BbGMhuRAZfEcoSqDr5ZkvNkO+RDGQ4tjbMz0ZKdpSFT8MSESEYABi1k
of5t+LAWtAKUZr45f3EQyiHmnPcp6WK6FFsWnW97ru8luMt0fIoI0Mo/W2DF
xNigGRoBVhy62StoCGctugpAfdkxDeCQgm4dDfboiKb3qEuuGPdNaSOxxr+h
1u7cJXFoyEprT5Obn6iZYWsCjkzlyQbhHFzDc2DqH9ssmbo3U0UlFCv65EG2
x4TLi0LpF7EEdcJlPXS9IMvMCbjpf9c4CobT+nVpgERj6YXfpsUi2wmHPGVo
8eMhz/6co/20lE9rLoXlGakgqIuZYw/w6a2E4qvc/zbpTOwfe/u+yEsKpgbd
wbF8eHNZOtX6xq2lgn8U+Qep4SgLnD6hBJSFk4SYnCS8lHfk5Ru4uSmy59OQ
PouaiCvWt54Z+hB4JavTWLnb7S+jCTmiCuB9Fy8Zfxvz+0JWAQpSUbjTuVyg
y9KMAimhoYObMg4meD/HJO9MaokPPVqy5YNuxcmYJZRFqFlHtquS55dAOOjT
3nWVJEMYfvt+qHMeLtKNqXsroVOwbXqu/R5BGCLwoJ5FD2IwxfaGxPSlzwfK
dp/oscBklCadvugLCY7rmsMtoR92RF+jLuULvl6wr0TY+ktUznjEDAbD+PtB
5rUgavBQuezwyQOTT8ZKTCrA/hWieZH+SrkKBsUKMxh/LHRC7/6QK7csD/mQ
YibrPa0zNFaNLHF7rjsbegxQdhKt5Y6u/ol6Mtwqbn3y41RvH0XN4HQ4ZuC3
TmTunJXMS13Kutjug6XcrJK4XS20zreexfp7wn2wmbf96pCVUrzvdGC87g6+
3H2D/5oM/fnSFMHZ+Oz5+cZ+jG3iEafk3q4/IZC3HOwKpL+mYuhmS9+q+FkF
86gWMOJMKh4YdlXcADK87gv8t/Z2hu8UcdQOZB8bq/aZbKmB/AaNQVKVEdoo
IfC60tGA0eZn6bHWjV86uRoAyweyiWvNE1qiIOpHn2rQjX5/fC6jGQ0arJuE
V32GZYMuBeLJDezL2ipvLSR9SedMx8ptv6WHLscSGL8p2eW66binKxkRSgOj
3ev7uBoLc5A6Q6QvPqKKA9KNbvEUQIu5FOIhoTPoh/7SwoLES0WoFKcbsdID
FWNhQWUP/eHKfY01zf0kt6JH2JfyJonB7ATgPrGEtBiowYiluqhteNdcJm2v
acveAlYLHJ24G6OHJCzQVKIIF7FYK6fdx6hr7Jxi0OjjmJOh4lqE6dvLgQoP
EvzPdCkrcFzzp7Oq+UO43XRSbc/i24tjSl0I8QFSeDJ0p9lefIwf3k4zW46k
hzl09r2UoYNffTXOIiBY0GBBB16VJqDJyvPOOqA1eFy1P9N+qR7wymQ2Vadf
aSgNrpmBylWrQzH+zYV5tCSAQN+GEiXJDlFoyxp7jUmc8AfW6URwtYpfVnRQ
Y/N94ETSXJhHD62qEq2pJh+M6BApY8pXjKDogx1E/I3I102fLBmb1hRV9qtG
9wYT5vkA7mE4Cm9eoCLkt4qU0ESFhtmlKzSbE101Pmiw/UP4z2gZCTKVKaby
OC0H/WbShaPcbADbI9CjzNiVJIWLmsiQgI1DCc0WT2Q/jmeBuj1OYXWLRLef
K+8hRBdd0IWZYxTrQAVHes9eGL1n0zw6RokHlpwaeBz8tnYAL1iX1SEgGUec
ZUsYes5VULWEm50ifVH8fi+jjTm7walMwcMdEHGBpeD775d6kvpoJgK4zjve
jGkui5LoxkX+wXdniCOvaAUFW8NMeYnxHpckwWhISaU/atCrVk7cYPqvx1LP
5s/Wc/w0BbjxTmSIBR9aQ6NNbmIcfTuSy2dzCM6HwnW0wMerLP37Pc9D8wsW
T4KjfmaMdiS9JSgX8X70Es9yU1ACo3D9Ie6q/dlvT9Zn/Yna2qUgIVX06ZO0
syWRfNCwJjwTlzqK1EmFFTyj9T8uiw29z06wFogT1260NB4PEieAe9C9dufR
lQBpoQ6KhjBF4RD2c5tjJjgSTdfo/NNz5GO2h6fi96Y9O5CxHQ5LbFLWvm7m
9mYFHVyVHeUJQDB6gxAtlYFybPqOZamA5v4A/mtHXnoO8TVdtWbdJLNnJnw+
9cvof/sSILz6z9vlshj4NsKAMgMhysev4F/kpZ/sWLubpqn4CangWvZKQ9GY
DPxuFiX3/WYL/NXgoHJ8UUxQOHbxqRVlDs9Ty6xWd+GpgOxK4gY+t4yYbRjL
FOuF9dkmmD7kzN0zXl0R2aaSaObw/uG0I9p/9PLvS/szsgRAutilWENj0bXW
TcwKa5HlsaIYz3yPiAXfE4TeeSz9q4596/7Uy5a2wIzztZjIIu6IUBV4zSJo
qfIKUWtXGkEds+K8zfZLwQ5CDAxh8ac74FGPSVdMDzC2ZG88pP0QIUmdStuZ
u6+jftmDdOf8GQxIV8wtecyAqwSNdiyzjd3gFa3ADlpVJsLUbqRILV4Or9t6
A3AFM5vxDTdExCiJkAdiQf6x1H+mFCwczjJZAjHVODdiUsohVZ2HBWCGO3Fg
6cnsiIdlMEIaSOXQM8aQK6igDTfLdAA0yv0FYM1ujHNEWq15On7qkpoFguAP
tAVjDJEeU6xhd4fRxM2FsOnPo2nYmUyyLneDM0eaQk2Ct+ERtPjYPm8dwL4K
YWq4O28bkx364mh3xphGBtZieFOEHDZ3bKZMZSR9LS7aqMBJaci4rARTMgnB
5f0WgOMREMFJPxJMCLFecpteyiTw4l/fO8KjAsRyfTbmVvD3rNY3Czxr/AGB
CEt7WEiLKccjPEc+fDQni6ui28t2oAJ14WF6z3JdecKgQxOSY7v+j9ra723I
1qsHmED93DJ4pga0cD8kxv2slVxVOcd+M9XqEGLcdiPqzbiygp1txJGuhpqc
o3aNeGvgTqUPxeGZ3Xm/uVZ1cFOJsxbm507rAGQNAf24n0nTNr0nmUbChwdQ
+zIJwhhRqUvwsbx9wMwT6/NlXzXIOf77FN07TplGa82LIz5rrqTvnAJUBbrj
gY5J2InFU/XmvceIOIx2yJN8wngVAVY9PihCPVSikLU4huTOlWGa9UGAVmEB
RdTT22usK54ECwTsDCBtBtQXqRbdNtnumt6+h6PLCVZ2P0aoYnozfd4e36mo
1XQeqqG7c5D/gbMg1nMfVQx3VDzUdJZIfYLeRgWEYz0pygBTothxynHC2aJa
WTcBabZnqrHDue3+Sa4/UmE14WaOT+3zTnttZWPSu03IsVBn0Ub3sgo9hCdZ
q9i2vbee58PCsTHebOwogJuXUfXt/p97k8wQcg6bI3mFpwPKR2Sk7vZ2ZFyX
Rj9WtLT7YO7jgPu+FdZDrn3yIm8KdLPBpaNYXQLuhNo/Zjcw7Zl4xtyyIXTr
GbuF+Ke2efDV1kFw9VjUIHHJqn0vS8WsK5Cfz2+2W9KOC+MPV92Wu5eb/3iU
UU8Svmr5m5b6uWxwwgNC+qVE+anW3zmDUHqtAPQ5b8gbjMQn8N7SFpItgiXc
os4M9z6sUBPggzTBmcwg4X3piI4F3GK4QlhwRR3a5TVX++1K8JZ8FsK4JU4r
XRdPGU1uef6lYmeh+kefhdZtem9CXN3dqQy2Wn7jyQm1/BgWa1chEx7ue00C
MdFKFxVz6ugvWQfdP5CX4POZ9ZgFQ3RAp/wpuVdZtUAYij7MHtHl0N9+7zTB
OWqp4Fs8RaQ/0hYcV98Whp8vdtAxtHQ8bdlTjQppF9+ZMDJuiI0iZJ4T10sK
8/Z1duOJPVydHhOsMvm1oEbp9+/m8wJnorLN06hGjQxP0xwYz0FLtHaw9/nJ
vv8JMo80u1qSFMsO4ce7T1DCHUekT/EpvY9uThcQesdtYWRY7ELrKdFgpG4/
r7P+yS7cYDaKCgnuZhp3LfAp8yg8QQ0zmWufIT81e/tzgzHfZLIJ/rk9sOl/
NtpuPwkK/gzceI+QIhuw33AWwrwra7LtNGfYck0lvkCllc1oruJujbNfmefh
GfNH/QV95iOiaJ8sStyrRZ4avMGIIs240l2c/ndVsf0HdiHf+WILSAAfpckz
to0QnWiHfn/iGjENdPb6GqSVfrLu1t/HvWEQoCBGVS/mdDf/JT7xAhIlYYwJ
J4D6xh3cADskLdV6ktxxsCWAQtZamznJ/yED1Y826qJQcxKjgfxHlrurgh9o
BjZnmLKwrYE615BC0IgbxdF0mpNpSXy0uP1cWs4bS/tzKZDZ0fyK+b4RvfFX
yMISJwDYIs5osRs6kOFGpeEbrRyX361HLAX3xM17SaeOFVB+V9CYZ1uAkIOA
EWEnxqAZyCMwPVnAgaxvwBKQfXgsD9rSpSkYv7cwjnt5pMJYCM0J9k+hWUTC
FCaS9R988rvURpcTshxfDxTXS4MRm+N3TYqf62diOlPEq1eic9xmjzfsOKyf
Q43+khMXtW6cOmf9V2pFhROhxWX+pY4My0mh9nuuTup3EuoDoQO8K1wRJ14m
raVz2W5cbHPhxG6QY1cKkgo29hYbmrqIZAlkmVE76+b0PMLFPhx5mbr8omRx
UU7FJccAR0gO2j1ExqcfJFpLfdgy9r8oKby5SUxekySDn1cM8GBGWsqtulJV
RVZ5vJpUU1swPd67LsDEUMiomxwRBrjK7Ec6VCHPEJEIrzMtdtgDaSWu/5C/
39MaAIaH9dVOK30qGpujVCtgN3Rwh3HjbnqMuGnIZgU0P6SdGtjiXJhNrzWv
M8BfzF9zav6hmH4U1f52o3Hgro9Qw/v4FbUUtqpgwFKj5QPb13+jp/n34YYm
w706x3fNJO6tXFE2XdJ22r2zMAbSALzrzF0gtXH+lMKmVGntLoTII0WtcKsO
w0kqkM/sBzzowrGtkrInv1uSVqBvN9BTWxEFM3UJ7tHQJbueHBce7aXmIepu
D/uL0DsJij494FG5DuPH4Q7ZwBI2Ha8OUHtkU/e2lXN2Xx6s0zZQOOscw6Ri
MFsyPIzTK6m+i9LL38LrQbB+8jCCJHmU3HPgAS5Khm0G1DsZlGYZs9Oqw8bq
MMzx3V39efKyp11UUpDnR8O7C29fVldStjRseJsKcWWLXFrRJuSWlYUFTUGe
xHSAZcuHuF4ou2tYe01Eb9SEZ5feuFIUtrhQ5spAQQjcBLSV+2bCQjsqH8f0
8d60ENjsu6qWnhojZxf9KGxQ61gCsyzUJeLKstV+jxlQc/EqCpNbyQf9AJXm
e7kqOcJGaHrqPy2u5kfE/KwOYG0WYuyqqb6h6PoU0DaDYx5fbAU1vUhGSG35
7sRmnVm4K9NZmEvydqvr3xPPwzXRqv5rbuAcFU+8OjRZkN4TQz1cyxPL7LsM
o/rJxF/nCoCs/FbrljHtbWeVu6fPEi7AxVuyAS1q5te4HrGfICaDS2mdPmR4
JNO0k6a9DkV9/5OF48Oku4wnmdGNo8ZPAay4lzjKEii371zLJZ2fKziYXPo7
DDxEhDIYGmoihvxiqyQ2L5WxZKTlRzRDyPhFFRxyVTRrG3eeMKGE/vCZoOoY
VEftlN3KC384g1uFJp3+LJdg84FXb6nLLvVkDwM3D5QLcdI/Zeq0uouERRhK
WZBele4eKqCXX5PADKUWdTdVeUOxbQhdI8OQFCQlhxBsHLLG78KF1ts4N9nH
OPkHwvq80m6eGNGZ3WgrM3fL/aG9umJr2mXY9ljfEzJhKCvMQhL1UkhRTqMs
a0VoUmKNSdyFDVuuhfy6FcSBxAzOyQ3MRW9xeIWZhLhaye/mAjDV97MXZS/X
KGQ6TO6crrF1bperOe1c1a92243iLz6106IGgjhivwI2LETOfPbicszfGOMM
eP6X7dKEyihhrqPaD4e+SbWd79BzVuZUDLf6unSnlsjCL+VDK2A3BZcS0H+1
uFsfpIRA/2Cq8NvXds4jo7Tp2c7X+A2zoq0wmQ8VCsj+ocCF+Pr/wOO1tYwW
h1r4dwI/NAmJdohwmwv17IegV2okjG4WckkricskGfeoUGbHbr7l1D6N4PkI
NuGaXQkr26+BT1iBRfglmlcwshRO6H1C4XmqGMAGC2i9R4X6HmEaApXGbijJ
DsVhvlMFdtrym+4Vzn1vzfH/BUwul9taAutfvtL9HrHF6r7gFqGDkL+4ohYB
6EGz9DuB5ViYmpdMXCB1Hz0ZlSQTlRnrF1j55h5QatJ4qL+anPkC5tMmf9d9
uGrq3WDo9+PLNbW7IJvE46s1JrQzT58IgmzTPFbLzn5h6TBmDnhpTQn1B37Y
M/7Igcvq4ZKeCgdPS/O/purGpAdNaVDd9arrz0KkRMg5aqeERR9rdSj97IwT
wiFFU2HvFTyOo5OHjSRI7tA1tYVCuarLlZmv+UnbpV2h6dzcWzUILYG3GUxD
CKHTGtpaQynGmvCm38VtgQFHBqcE0MEqvisl8/XwnI2Ev0YEG/32HLx0hPNJ
Q3iIirsOtKQXMZveQwExdJl/MI3hSaViug/jCDrbC4FeEHrDhG39CfAp1PBN
CxvLGhRrv6fIJizoZhes5Ir9uYAJqtT3JbxK4P95EhIFjbgX5wZt+Xzs8/k0
dzibPmR/THPHtow6Kie3rxLLYVKldzV+11n2gohZ4dueZfWaZW9/fESbGVID
5eAtTog00Z56VDFiRXnDo4HV2c5JuT4nLaaoe39lFS6DPbvs1PcPksfL40zj
sZuLVTv5sbXeczwA4C2z7h0/ZtW0Rov7KSyXKgwC9wt95nWoO6hczVH3CFbP
7PSSGFcUNW8ttLe1EGKulqj58WNY/bveaM39uawTotmzmxEknK3KsCXdxKoX
3IDnq+k9QW/BHKYBpH7KwuK8D45HRv2gopxazkk3sbEYu1Q3VrBYapi7zUZn
jxaHeol8sgAu0I9pswe8FDWaKhW5JPNwM9vHO8Aj0ZDeAWAjeqAoRhEhQBc7
ADf9BBduiNKZTqeZ3TGD0njkOjgFsXIhyJJhX+uezoqw8xymApkugX+WkwCv
6+3C5NidQQSyw/YuOBKoGSz3j2HjXBLXoGINCcOz1qiCLe96oPyg2nv7gI4e
ooQy08Q5grdub7gezhctAlOFtpcWUA5QWNcYaJAEyZdrUFVWFW5MEFZOwq7i
1ri95aTsl0Te0ylyVOhuZWeSZdkayce3e6UVvGSljADSYa19SoFWVi8xIk2Q
snZy4xEIZSJKwdUfzlHy0IHj0JetEeY2RZQs/0zS3c7cmfYkgP/IHOxn6szf
z0PnsIbGcZu/xgGZ02qvWpGvm/TxW8yGjCRAC1dULAt9eEGRKtS9gypPbOiy
+EfdBGB4Y8XIMT/i7kBijtuCa1gKfzQsS8yaOX5RL5/60A6SM2hBhrOWNkPX
TDJrRWVWtuf+qHMLMaEDdn+TC1jOwLTOLjud5PUdmKnSEHop8g/dQeOWAw+f
k+zrAMsnHsCGJhuM6/5CUmXXJHHEoex/PU/usgM36WPkHZL/9wd3eaFZNrU3
fDUK13fKasqzTtgevNTdqSJEqiKH8cvFSZgcoi3Rslz8rmsRC5eiyTLoZssU
6gUCOM3eeAkTrWkqJcLQaMcyop7az36a7ieovu20XqKm1kOG6ymSbmuF5kdH
/n+JI2pgmGueJGRl9R3ajtku6sc0NB0NQDHweEC6cTXwrM5Dq+1CWC/SFE7K
joherxGqq3Vie0q/UZCjZ0bxfBMmOUvOI6s2yPBWxlPxnZQHD5ETul6FfANq
KtmzeEMenQY/sMk0/Z0wlKZRUvEa1T+HbImW7D8owmTHinwzm3k8b26C4MUf
8Xj2KSJXwsNf3Tuoj5Ri5zet7D3CS73ylVQAcz+jl3LBaD6lnscHlCxT0JYx
Yu2jZWQxkzL44D/sy32KJMJHxlXuLOR6cxzVZxygO96E6M4zKemAXA8cWJbu
JVwjFvutkMQxKiPTmMp5h36hao/VHp6Jser3mlKdyUGXcq/JCIRuWyCC8B5J
5DE7m1dLfCEXqVL55LPJapN+3sXUCJ8Dhl1D/QI98LH7nZ1753o98B0woZBC
WePjLiIsUKo9J+ww3UbVTFVd1Jrq8hmb2NffhGkm6N1a92PhPgrAazEXvEaV
w5RoWKLoP97TCoFmonH1cVdcoaUjh04edkczVbpobGixl/1XFaClWOrXBhDo
otnPphV3OzB+utEN8OVRNILEAOK12yrqTCVId/jQolf3ONQC7J5PWJFncQII
EpaI+EKOwnlzkVPR7Zk7mW4RSl+vd3Xxk/ToCXX0WcD2Ddi/VF9Y5GRrp1Kg
e+qG/+9Z5CwHcDgkyVhI3Ve5p4Gk5+ezplFfXZIttgjJP86VzpL8L8Lwcdl7
h5PtylJtXdfm+BgmM7/eF6WiWE7tBClmwMyv2jQc0zYPrr7J31x3GDTMw23d
HNCmjpQtR8luvVtHEJuXwVz5vDHvg50aB4IHMTY4Vu73Z8CUeTiQScQ+M8k+
3+5qD1wkclvwDTxyR4NCi7EjHcTbwOC1D7OxbzLKdsV6nYsBEJnOskAthz7L
s1/77ZfuNz2mNPV7kwjX9sICNrlrh+C29COGzl2n5jUwsfOOKmhGo+yzG5pQ
Ef6lwAV4zJZ1uTMX0GTjNygZd9j6vc5dVmKx0eSkSHeL63L1kuKtCOe8ivMn
AtRmUlYGjPB1gepETza83vHPsJOxt4Z/am2UM9LT8A3Li9IBGcfK/qIAYXVd
eLL9HWtHkGb9kudqG6LN+1IFkoODEeEoSiQc+Dy48psuSGeoIHZhfQMnsS1F
v6NVwy9E7uHYup57+iNDCvKpi6OQjiHPlW9OLEFIWOQvjcL+H27hRhRGVzZD
kX9xhzhtf6xEDzagkzgCn/F7ov1WeTwUEg31r+bcUtHNh0LN7xqEpw/+jz5l
Rm/E5zs8bi8tPzEhaQyGJsJFHh5s6WpNMdZ9kL1Ghee3mxbBtOkx4ExK4j6W
z6gtBmVnaVwxXNCNk8dCNLASASq5+x4kVE8cpkzoEupYKrD4zz8z5gU9RJns
+Lpf20tK2+mhO8OYXsGjn12GbPHRmqbC3Bgx9jajGKC7vaM8vyMam0qFMFqg
GJOwFawEHsXKx/KapitrhluY9SpP9VbTY3NP5jVhXA0w5MnyFxfWL2d/e5Lv
ePVj4fdlJX+QZJm8takrJriIgiQvM365y+qxpmrVNmMypdwl91iBVgpfOYRS
xV+x1sflKLE86GuuqZeI+kFpKbdV8MaG7Yv/Zy8OVjvGH87tDuRMmFh+DdTy
Tm78Mx1lLcU0jh2y3GGsE35mIliktQ4D1rlEolO5qibwsAifvoTWS7rhigyT
MFJIldYOk166hJuSsLzM6tzBKOpW8f9XwBJskd3mH5/imERj6c2HkImUCC8E
dE6/Gy8wJN+g8YBP8pavfFSJl0WJgxHMMtT99Hvur1Vw7HInfQola2vBE906
LflhnmZmkbHbFtNy0kNGK24MMWHJrbxL/pUwMULT4WzQq0NCHaiENNeLGeug
NJsjSbQlqm0oobUWq4zT6h+U00UTh5sYGO8prrxoxfpNFkQEIdo+tklgSaHQ
PnvxtqdC2nBwF2u559U4hFn24Qn4gWvS128itPNJMrnaRtKwJMz31pIYRBe5
RfRrBpLrHssXlb1debCnhNuGeJgh+H18iDoaIbfHer/nPgcz/IGsXnZ5JcRS
Ez9f8PRfG4wchX2JTou+AXQuDdYih1+mDeczYic5lkMuIZxAsDjS7TdPaO0F
a5OIX5tDw438vyxPxbW3X9B4HD+n52DRzZfYkS5mQZrJdY9Z06Q4zL78nnv5
mU4GIZwNid3kPEASXdRkDvM9rBpL/jigIm5sU16ACoEn91DMphJQwureaWcR
XiuvE+JTDJRHgysHJ6dD/27JzNEEPqZG5NbGvyPXrs1rV00y4BWcGI4g9AUS
AX6VkFjgMZGnCrk7rfTlWGHNRmdE8SnGFEifhGlIJZv72pweyNNtsQFi98gc
iumv00vk1VfXbrCrmbPOaZeX9cTGA7UvDI1r1lECMUNuzXfzSmBNS5KfzK3e
T6LbEmxN3VTGO3NWtMXkixhfDwtjy6r+EMOydH+182lOPjinkDLFmT9yjQkt
dZTjS0Dsujaz2FPLanXLQmwEK+apMqEynCy5zNbFxyxzl0h908wjheQpFg+z
76rgjDTl2V5LIUtEyrmK5hXAhmguzNMDK8QGhzy1C8/5pyQQ+SuZ/8PViZeb
7IMgX84TSrsEDRDaBTgbHCcb9O0KqwR4UA32y9M+W3GL3Q1WhwgMUesdlF3p
85E3fdRmzaHvWIsAUXGDsqsZUbODe7CQl6nljMdjMttBTArEUealwwAN3icu
YVa/BsL2SdFsP/5+RQ4M6kfqkQujHHFIFo6A+aBnGjhtFFrxz0invxy7jBNn
0sQiHreEW09jecFbhD+15oatcm9g0qEZ51AhqCJ+oOBHY8aWSGYHCpT/geaP
Cr28uI4948PCvuumc5BumPvEWMuacgSDX/rkJDX7VyJuleWceizGCshhsmkL
55OKAbCh9WAPNGQ0V3vEPdCDXISsIICKW1QUhlPSr6dOVbz/GFx2Fk4ofWk5
SdkYHM8tP8HS4A1qhOViBj2XTVObwEe1Xn4aUf8ah2GsHfoM5SyhbYs5ynQ1
mwNt2Sd8aPA2Vcj87JDDlQTdJYCOYV0gAXq5Q/sI6d310j3KHxonTF21eL2M
s7R6LwcieD6UL/Aa0ZxvU8wCAZGINwVDVbDTal1zKCtEICv0ueGMaB2ip/D2
BoXDWAPPtU3hiCmxow0vcFFQf8NGzs0nmLc6jqMdPqfq8vZnKKSQROAIfFP7
cmzpx0ZkXQP7Kgs2bz4WI6U8yC7F+sL3Mxi7DN26ISdegCn8PkffY/44ND1D
WIuA7jYw4Qgn/ZnQlbC3uymyVytmqjRSS9wyHf4iLKtY4K1xQv1VvvrDD3I+
v0msiP+Tvo9VI3PAD7iPVOgdMkE/tSUKZ9YjomjnDhmkClnOMhlL8ZactDuW
H0oAmNgOdEFB/f3opO4I9MjaF0eaW2X7sCTtsvaJfhpMKn0w3J9wZzqkyJ/M
vA/kXM6PfUbDdiwyfXvEnhc2YjtwL6WjOFaWtFV3PI5WyIZCHcQG7Lguzd0I
kB2MXR7doEDLGV9KcdjjqbVY1fXI8YkNfv2yFJlVjfCPH9XAKK42zqPV1PBO
kFc2kqq7iOuxcCfkThA9IFEerReAJQLWI8R848pjzsirG4UbdMc2ZV23hnbE
x12a2g7l0MOWtZbLzzyNrHdkyxRyQq7iu+X77myeNwwEAMWwl+75KOdsblzO
8dro0tJSZHq/T4dbe6Td/r0Qohm11kvWHy7TmDjxGqgozkKQuvernAnJjj7z
rK2G2RWQxghcRNTWcSiUSm9+szbH0S+pDvhcp15BfEctvlUsCYFajryVSoNY
Ex67U6wlfJbm7uyaTkBJ56hpFujgG9zuFUl6KSK5lBb6yCM5adawTqAQ3FZg
JGlj9zyYrZT7hRntY2QF8YUQq+IeQDzMvVFMfn8i7J9ly8syZNxqwkuozLi+
XfppO09wOvIfijMGuMQNb2m3vO2Tx4utMAHldiHkMgh3zJZ47lL3pzx+H1ix
z1fDB/HY9YfvLYOwyuNQOQGjdZtFniEklCcy7mQ82pRgwNAViK50Wg6PRUnN
pXAafNSHuCHU0DPu28xLSDHna3W5zvDkeNrgyvFIWdRdmbNkGJ2KCjaWu0HJ
3dFqR7m5dQzhw3nEMSZoDBBdH9XQOreCldv8Q39Ct9Ji3qgm2wRolQOWbdxJ
2Xv1ppTAWwbKYghTDlNSxNYBVdRI6MWgaGDPb7M3tB5WOzyFwn+1iPWsP6Iz
d6GvDO39tLxsxrJRPsiOknq5kWQ6GYLuriVi/YYY/+Qe2MeLyJ5Abv7MOkiL
t/x5bQhsEvPDSk8RZZJ4ZAR+J2mfT9YWMJcJOU829No3XU1U68UAaexat6xn
hD03fQODx9pSgZkAJTq/DXmnu+8xzj/4fpVGSK+/pz+Q8DH9KDpV5id6H8Oy
XKXFQM0yY6CkZHF42s+kVmRqAVlEbM6mwxsCS1JH1NPPgfm5oxl9KTqLLvrq
oONHh5Pxsnk5diPLo31djhhwK4IOWboKFLmQLFAwVBf1LYZfukCGZAoYTyJG
+kMGzYyL/ziw549a1+dz3K5gpNqSh2EI+RB2DGLfeP2hM60p+HNMqvu6FiPl
Pvuo3IYYcfznkCVnJ6LW7AzjTSjpzgTALpbUyVg5uQOVrV7hv7+PM6W9/CIh
S5DKQqQUlpDzL5WYJvpX3i4ibkpYmya4cuIY0/LLkB6mzXY1D5lgkBMDYCvH
1LJCJIkOo/znfKYG23U9kuPc4wYzjZD7Ma9L1Dn2MVfvT982NvQ51PLrpYT/
2jIqZMd/Dsaz4JbLOhLAj+zZ6PNVFqbx+aPKVFqphJx1vyv3bsrXVBVKJ0Bt
YjPJ8RzkxrbdsD+3znmU6/sLnBphHRb/A+0xlqPd6VXbh9C3nX9nHy62AKks
r0W93w1CqrIi+3cCShjjlxP+JaWdKqBJU7fV6oAlZHivMBtBtt7V9KLviHYx
JiQsNlf6UxMqZ1jytn0gYwPFDyhgIrlYD0CqUrtcj4SI1Uxh/uqS7chtHgb9
5KN3MGqN5zs/EvqfLe0BA9yCg+dk5A/gfHnBkczskN7s3B5o2HrEmtnOkdnx
b88GId1ORJRbwn0kJZCa8noSzz7FxWqTj/9b7T+gCwd6w8/hcDWvcyv71Dzk
P3JeFb5P8aeDdOu8Hs0yS5V4HFK0f2RRYjVz12XTKCI3pV9m7jQQ+OCzeyob
B0XhV5RcIqtVtK+uXMrqZLv6IP10B+oXJvoTPHV68XiNYpyI1wxkrTzsH+Af
R1UwjtyOyLVcX+pgJuSlXt+qOHy0AyRKtmZcT/uP4bKJm9Cii9AhnmxJ2Dwr
rbqREmD2y6i2Yuk+SKtDk1IAcXivK8XlPGO9b5X9jpiVgUr4WqbCTNJD9XM9
P1oRwyIEcsEYSnfGt3H8Pkig+BQbl/5pp/5C2YzF0OxcETLlEGdSMMPOu4DJ
mNltVj3en1HjF1xtUXX9AmaiYYpvYQ1YaXjXM1V6cd4dV94yLY5Bik4XLJOY
jdJc1z/JI5IJy3HuOKA7987m40gH4ZJ96CzzbWbvwRdh/wxuShDTeZxNE8bq
7SsSILmcMN0xI2FM3heQdSqkI8CQ55VhnQxJiTbmP3aiWKqiL+PDjHwFW8lD
CEG9WypPtSJiqXXpHwhgFw8DWUFchEMND9+Q/5XvB59+9GXKaQwDe4WgynDj
3N6a4gbwQcBMxScx779hemKZOYp9uqRJiYJrJ46puiVasFAUnsEgp0rZ2e5E
rGAP4aS7EKt8glCcFhB1SOm3uVix4HzCVD3b7PZGI6ThsL8pEgfm2UMB3DyN
l2R4Wxlea2PgENF4bt1euaCGRSVG2YV4tWnGmgx8OcvBFe5vV0IWLv9Vtgwz
ufgN6SFDFEmr5SJfDhfR3y/XTID/u3iVBYGZZKzOtZFZGTTIGzI2/CSIzBhq
ePgYb0ha+Fk6DE9IHUS3UeFyQI4IKigcKrJX/kpyK1V+zkx0bAroVgHFm0mx
6xeBQc+1jL2dVNk1R6SXQA+ydFsuVGEyEk+CoMRvLmzwiVdPcGopoKxDQ1V7
0SicETkfWDuT4Eq2E8JGVhzUNjAmSPMEW9ucHgcAxYgNy6mpZUIN71/WiEYE
1/x2wy7vKBq4asBfhDphZQ2W/zBiWRxrY600xLRzdHcskJdQBClOfkIsSBc4
yA1hwgwnyCIdOVarb1eOfazkr/QDiAdd3kj+kBRooCJbDKiAqeNfeI7tz4VF
Ip0Z1HsuMp5ppodPLk2KZB+9aIP2nc9nLlGgc1SqUljwwTm4X8OzA+6I2220
oZMnDT9yli4LUtY9SKTJQHax8wTzB8UahHNrwID0+VFy7/AdCO43QvF5y+Mn
kHpjlvwvUJnoH12rbbg9bfZoMBXhb4sLdUuW1+7usjVsJGfsN50CNlew9LOi
0ofs5n8LtoufKF7QXfIgxKauXJcPZ0PmO2iwzuhzq9CU1JucuJmN3qZIe2mQ
L9k288y+/60FIspeX/DUO0CxNATX+E6iXB9MvOo6qhtPQpu831XYotx/xltR
IK7K2+MvFHxifQUf3vpRNC8EDd9hrDsze0Wvy+iLKtmmrSimcjhOhWOAWkxZ
Qk10v4TgOUpUVde7srXIWVPe4Exif8FvDf7+M66o9RCC98I4l3rYwGRj1b9+
RaooGfd51RNtADPPgcD2Ua6S6IdxFx6bsb81+va0NW5+O9RdKhSBanJ+8yTT
2TEknSZ0dSWQProB/dAsIc4aUIVnDd4/ZyrnPHxcA+4ZS2un8x01DEm2+OUu
iGJOYJzc2StucYqcLCmf4pDk2XVsQwoXqaXlPmdDXtaMwmJf7LWl7rsrb2vA
DvpoPVY9nyC2Ve8IqflYLkfKTqEI91PaU6pCRhQ5zB4AiGC7cyRG3ryJ8rtk
RxlZtdgE3pk3jEoTIMdKAfs5SBWW/anqe0/6KPmr6srkwxhX/vgCrUG4Csa9
mBZPDJPhgu1TD/G2fe05qi9AvF8SMiQv5MskWkFnk8U8BnusfAGn2REb8weF
1oK09WKMBN0l+dXSKzCvnB2Jxc647odR/HPHR7/UPhdmMRPuSG9jLs1bfmFJ
6yBdcVSLDCnHw1dLAPmuKWxaTh4Kg8onKBIEikKRgGYN+IaDaaD7ZHj2Wjpf
ZyK6zU5j7CAp1cmLZfHzzVgyhJLmU+VSWdCWfxOO+NXQQfBBsVAfylzztZ35
XWIOubHNbydaYCVuEazfbFvxjyf76c9vD2HogAlSe1froAR0m2X7FVpoZBQS
JtvxMQTLKUaQyPgD2tncf2vb/dH3wZ8gqs5dTygtLx1Mrv51JKwTQJCKV11p
oZpDBNISQc/tIKOM4ep7l+EJFXHNcrIs2q4vmIhlSjJTR1peB3ViWa6GvNwn
CYM1Le/JBTOofx+8ws5CQye6X6UuT0QgA0WK+kY9W701CUgVfA2hTqDxcAw4
/irmf0nzAxU3IwB5czTiWj4FdCueFv+5iFso0cGNTKbdd8GUm/5q8nv8OBAw
JxSQsaVh4VwNogIxDZIrqgyIjN/x/HyEfD3LleXlnZ3JBvu581brOD7eDp61
h6AWbh/5H7qrZ2cI7WOBPf8fZfgU3QRB+p3mIco6UVBZYAyVUFlgTqwJAXZM
8CBX4oyYd5Q97uOIBnAaGS7pVk7hUh/9VtY564v0xjKkGqX4BzbIOyZfEmXS
FHKZTiTzYXu8xlmecizx3azoVDu8UlAUa7zFRyoTZF9ZIoE0YN1hvdz4/iCT
IoGBp29nJGTwfD2mB8cIOgtK6sn3cVT3RYYUcEJK7jL71MhEiHN99bBNq4kD
pJ52fyWXwbsbr3jCGBLGwbB6dFcBN1ucmhnX8S49MValnUSVl7xUAvN6TbGT
X3taBRnoSzh6/k9vPuBpx5aTt5p15fENMVaV9LYwpiqUlQApSBCjFUK7cERZ
z2vcLFbi6MosgCe4/JtZqwGHDn6wTby7x8J+TX7u5CM9tzrhvay5pottKUqk
jfSkrILipTwOjpVH73Aw+6OEPGis6uXRvZoHV/WstIr7Y/nBK/StLBQGnoxh
fkIb0xtWSvtDSrpT0aIMUFxjwTpP8ahN/TQ2xj91MEki3GIoq3MSufLlf6J8
rx75gaMw4YJtaMoIO/aa4GspvajG0itcO/3I8jiHYCqRKwt2vykBDoHsQani
46UkfR9L1v+OBCwZz2sN6H+aXCMUzGiOB7Mdf3R8R1BQRm/nwQ9TYr99ePnK
yeVP/roryYhPkbV6xKM3JwykOIc9JyYmtDzmjRaJuw2j/HGe1s18WMvYM7nb
cmC+Pj6EnrNDaSwwGn1hJLSNGWAxCIxrQOZAzcvjfWs8+ok2utNywCqD/Nt1
dmzelt6psrkjA8WD7SwfBZMBDJIEWcMHnUzjYpD1o7D6pql0zPvidq1g7euX
mw1BNaaM6ZyovJ71pXw1VN4oAwV+hfEqKP8n4LTa0xEDoOlw/XZRlCY7xv/I
x8PkF+r/vydrg1hzz1NV7GyAaKxJTvGKlePcwzqbigS2bL+MnsdC3lobUcEv
R6g1REma3F/b5NjhKtbaweeSoIiSEIj/31y25ziTlMGe8bCzBocpQTbDExGj
EWaOvzEHKyL+x9YB3zHU1+o/VG8V4lqi+ZrxnJoBYTqPpyFNO4JaNry2Hx9O
jhV7Cm64ra/MazeaD5fW5oriMurusybpEMzno+fCCfaCblw27IY/zyW6U4uu
PWQcMqJ+4LFliUuKpvdY8CKyRJecNJ+BlXGezVDDVCIf+SgZTGrtOKZ9RWJv
AxcPxw/Yoxi+I5DvOSknhTBAjaPHlZkfsCX7yRUoT3WvMltOF13dmK3bHDY4
yoBfpwkf32nKT48sqoCfAGKFkSf/IfUiksI80d2RZ4Kk8vcTrySFUZy2HI9p
gvChD2yPyw7G2/ilLJXp5rawH7nGX4YL7DCpFVRW3604N40qfShXDjBbE3Id
jCtO/a9x+ODJiUZ+WZow+OVCuvF/ySIHk/rTbhBFxxeNNn+PMK9ZltoetQ5R
0prKjmttNT2zlsiNGGOpevEbNCYOe9+frRIOerkEwFXPeCfW/CbD8x6dDKtx
B/0HMRFcAUkBGwr9A5wYZDn5hOi3QyDO0BXsmbRbEh0GbuWxxH1wqJNOnTZs
Ag5ln31G6qxWeWttmvGP9dQvVhs4c4kex3mI69qeh3nXvBjFhrNglAEEdZKt
ShyNONihMi7vy1h46bnqnc4ztTJRVJjCsur7Zyp4JnnUhYZEj0zTdf/8qiz/
mmD5/UwsvRm4G50OhYzW4/KS+odf4nHK9OMdr3EOhKdEj/8D1iYvzb7K9IRJ
4UKpo3C2xfJWxyLPP2vHoyv0axlboVK/rH2VuGhwVP89TrCThdWTZ9Yf01DO
goUQqT8OpYuG8gc0VvkoXt79rsERH79/kvi7mUWq1KXNwTPC7jrR4HR2e0Rl
y/5vNdGrVEWG76s4kp1uLJJ8H9MBYKZBwiOQ0+b4Qm1RyuZSSU3K5In30b7X
91rjGTCzBlubf6KAbu+pUhBLIbARK7z+mZ3f/zlnutuxxPKfDRAjgGfyX66Y
ecmLHN2VZtW3tY1BWAqchqPuzbGqEbKd9EWshLAhsH+tPLSTVXVstHyJJiGy
O5aKw+14cfKtCi9lhPx/F0fUws7zyAoJPnH6+q9TwoobJsC5WF65aeqKgIQW
N93iyO56+r7QOTI3wKWSdU/0JkvmmhFU3HJX4ZoDeZ4TkfDfhCKQxgYp4499
SimANTcQ6HLYFN+i8CYoLeYOKME2G0Qd9X91M8kV4GGnq+T4PS8VoVmsnClg
x108cOg5iP+bNJ7hYLSSPQKBD1hI1UFSJW9/4PHCwR8v+FnFO7QMwD1Z6XkK
lv8YYDETjqcmqX3tLLg+mQBpLW/0tAK8J8ms+FqqA6csQRSbpLqN4jk5z7sA
ZeFn6vgPd0eTNcz4Z+DNuXIL0N7hu2fntp+/TWUpYFMEWmv8JyB9BTEJpsUH
Yp13OP7YYPyGu4VxlB8Ez3DbtVE7sZrJQshcziK6AegpSB2QvZL4SFY/IYN5
KpV0EM02x8zZEbt8OsTns2cVMtKOuWiFeOJHU7X4YHM9tFOQjRlfG17oxGGl
Ya/wdQh/+A8cscR/1tVCXoBJcgbp0mx7+XsXrX4Ad5E3IrliV5mj7RYPjaYI
YlLdD+giWBJqYX5SZ0M3cRaStlBeNchDmZj3hE9GMVsap9d34KBmUZF3G24F
G1BcYUfaH7YRvqIAXNVYRq/F5r1qUJNcfgcXRSQz//+sElJY6Y3M6b/amxD3
mxg7ibHs6TyBRCwIMqdfh10pa8pPivJTnrkNKclg8oLlb+r7mzAe0vlzXf6f
F0Bt+fNzhiCeImriiX33ckmRUvwEuu07dwwUbpLoxDiXrItmgGVRRGjh6e/t
fIktRzJWohwrLFa7axoh56ki/LLpOuEztoIG1PidNA073LJRa1NR9ShN6n8g
JEwpfzSgBY967VIOiA4iQRB6+Wj0ELKATsayFW5FJ2nBZGQeOOa6AP3PKzqZ
XcjDcmPhCjq6FiXMedN/54y29mi6470//1L8HyvnOk7GO7Szkom59zWM2Eyx
ZmfUPO4xyfMKKYwS0A82qDc9/9pg97UNl/gkqI3uXIX7+mqO9o1EK6LF46Wj
aLiNLNB2aYk/hJl6urul5+CnN1lGM/ZbysjHfJgVRj57XgERTIIGH8fUjCkq
/eNnWvBPOxEj7Kxc+oBtxz3vbzqTohXQuFIwuQuqVBwmjD9/czC6C2EzSkxZ
/qftYv7hr5AMzAFRxpGJbK6TrMc5Z62BzOMeQZXHmQObS1iVlEGOZK6aG73A
p0nbocCpG0c+4q51oQO0S1k5JcTsQYDm4F3rIKq4+SSMfk5gldleXB/Dc66q
8myI9TjxJ+3+ajg61NSQx8UdYLfoeFJuitTH9N1X2y8BgIk/VIifJD1A7L0c
082no1oCMaqRBmhc7bj77Qh6tUL8aFcXPT9qcy3F4tLAijD1UnAnKkD5bolV
AFQ5d0ptO2h6gsYAh0DCRCvSdgh+Q8cvgMG6v1bb9WS//AmPCJpqEq+W9UEl
B6XTzFOVON4m8rAWBJPLLk4sNigVmhV5gILYf+StnYQ2oJfabpJqzpoQIfrA
xhLqCkwU18putk6XOTpzbwKz6BbZOjzvKGzoEpUU38qeD0znLjdzN8UnBqjf
VBpNobWWHoTU6tgje0d+dZHXIw0j/BAEaNN76eRylIolFh0kUHhPtjc0qnGS
XOpY0m+pilHNQwPZoefTZQqZoM2WVb51OEbQ59YBc90ySvLhmwED9jgKgurX
FxQIqNGk7x07hJNlON6OIym+kXv29hfzLoc+W5S4aZiOVgki4xVF5/A8hbc9
J59uDsEGrMOGrd80Hg12Xcb6FMI8j5T8FH3qMD0VKBL50DdhIuEK/006OCXI
cV+uSucEIfO5IZfw6429qV0X0PvJMDx78y0DTYGcWKl3bh1XwgL1PXeop9Fz
4O87rJhl8cPAFA7yqbfKzcmiQna2ChclrOdOfDS/+XExWKW33W6kjy4sVqKn
XA50osEYRmaIGplWtO+HKQCzhEzaPljGgKXJFAhYobZNFoztEQHr44RoDHpG
Cv0+xm4HSEYluUdW5May1Km0BHhhCdVaulXMA+d3f1kDqKAkDDkBEWb39/MO
rjUG/gxl7ASeyd6KyihnS9l8OAdENKnhKgmImqaUleHBP+FQ/jPze3ydWpdW
5GMgi+3WjBbJcWUP51ViQzvFbDs+4aC+W2/I2JoLqbsdLtOUKIOezrfkWeOE
eU5KE3p9fT9f9pZSDC7LhyfEEMmP6LLCj7ZSe9P67/33hO7iNWHbpq5i3s8X
pyxY9brj1l+fNlXTdubBMN2aIpR9uy9d2+3qnucvwmgncRHU8FV0piL5riyN
hOp4ndHGwe6E6BQuAKigsqrtQnXTyH2X6ns2PQtgPelPQYuMvuaYrciL+m8c
aNSiCuGro6TN7Ize96MMyatF25uoZ3aHtCypldcLE85EiEigwV21/QEU/woW
l76KP8bLdS+nrzL7W3t0RBF4kjtT1McKOMLNdVI7iHcDSL/kKRrfcQWwCJ4K
A097upoC/VsX/XfB2XCycZGr2FAVeUcNbwV09ulg/eE4zt6xxqAqNbC9+e4a
QnWzZCQH03bUouNwBwdi04vkAXVS4LAO19TCCoTGtsGpNrzcMN2jGqIyG2OX
SC2dKt+JAIAta320DM34DpmjT1DRiKzV/0lFW0gCFDp8LbAGvlRG3w4DGGbl
hqlnYqvAWVeiF4/fRIdz0PzMxm6IhnODA1jSYQA9fev2Oa91EAvLRjCBwU4H
0cf6oQ4GBZ2y6WwFIHD2MA6OsnZilr4t/7Jhsptu11xniZXsqnr78fGYcCuM
WaVY7Fr4DvXAm35VSrvtwsSpAgmJ49WvISx7Re+TwSh2K6f4xnUEDDcXu4LT
xw8oxrUu5Kf+ZVYN+4/bnIKkVBh+2CPLpgB5hjaRts4k+n+vaYN6nqsVe3Rz
3VSG0gn73CntsOMisnAE/GB7a0nZr+EVOQ3OIG9R0uSU8iPURPp+MVTbFfIP
GW81mMvuyshne1kjpmd8/x76O4R30uKyrZsVyOqtspUz+FYZwbowYapL3n5L
g8Trs3MbEaZcWIGVXZW7Q1+dLzMahYd/QKsRKr1t5Lr5T5NbT1t4o0/sRRzp
plIcF4RL5l7qRimnj7l5WiPazFhs+nNbXwh0JkkF1cv9KEJzo/YTx5PZdJBv
9rrkOSnyFZdMrFmX1lizeaAWlf690O0JKsWwjcg3domPGjoL9qzKPeEGPUG6
F6q3N3L1DWP2BwutrbfjBCoOVAN4zdxoRXE6Fr5d43KrLRlxs4v96wX7Z/qG
f/M62uYUBsJJptphug6R/0dU7BT/TnNCxXthR+et4rKv+zNE+TmP39IGeKCv
9lekjmxvcJNEDr5Eob8F749AANjyrpjYcTUJXWyyeV3YrRNpn0KLEvuTfK1I
Vu3skq2RSPoNI81jEhtYO1CsOz5hYTfItnH9Yb5mtAZp8vrCKqcP0g+bz1en
N1CmUC/TEskwwTiFCBeNGoxTc6fy1UyyVXeu90o0oMxghYCIHV9SXA7CcF9a
KyHyythe8pYrHbe8/5L5vvGRbiP+/5OiRNlzh4mPp+FCugme5sbWGCOHuDeR
ur7ILha/OmaGEQqmXZhM0NbtEyiBQeLRewRM5QXnZxj+jdak4Bz6KBAhzRMS
Cfoy3JbYPtVzwv9gJB/6e5qvz2xd7ylHcD/SCNPz1wnRnMpFfE42xiyl+q4k
Vno9OvL8SSLXPPGLYR1sULbWcw9u+4xxL97XPzDb+9shp18axhJo7c0aq81J
HggnDEVFYm5pqxaBL2+JBiNUdn8qma1t4Py8roh34ilMF5ptRFq7gjmp5Vh1
MZKN19ICYJFoD8f9GLqZocVUJRA3UAd4cmkczOHr5BGbASoXTeAYxilqQikR
LQobkX0LDbPvAvDA1IrRcC3+ysplhS+SpKF0s95eQc6amJAUUpag8VMXqNN3
gaOx8G98vzl+Guts7893kKg24Oy+QbRRh+URegcwOC89ie1tfXhO5cGArtDZ
r9G5qnvNBO7HXiBg/JOV3cpuvtjxmJ5fKkku5imLfNzaQ1r9XE4YfSAbmd5o
b97BhHYy+o1Ay8J++0fTpg9mZIbD8O8GP5GvwY/GRMRYllZx2g7cb4/JnwPc
UMNgzHMl8TINc4ixp622TcUvzFIF0CpWEW2rZ7SS6Syr34oebJ7q4tiXJqKW
klrxL1fNcE7GGLOE7vMSUzB2ojR7g35pQu10GFQoQ+dv1+IGFbdN7iddQzTN
sLmi1pKgFRvUa2i2HZpS7jUBUldDo7C+uaBcd/qlb5Z8oO4KcWMa1t9uMqo4
6+Yqi5CK7GtFPuhEJX0m1qZFr0Z/Inf8CUKV8HmYSgBT+utYK7dTma2GJH77
69L+Tm3/tOE6uSKVyHmxF2r7vaIgbqBBHfrKzkPCKddOI8iI3GTA6HOlFgc2
k8AZjH0EyE4y6rj8el1h8VnYuq1889wxH5cLaIsoQE3EmCtpHW42VIoWkaFg
ZKeszvmQOFwLDVpPuulXM51knns0moe5SVakdtTSTC2STinNK4fmIU/d+ZKu
j9CyX5b4ZtE7txKokMCOwtuZkHsxfjI/B518A3upRzX0ctQUuQdPsMB+W+NT
Q8f3k08YKslG8As7sGmySBA9OU9bM7kx+Q1fuFvfP3HU6f3KB6R+ZwrMmZLL
PqZaVoOoKJyVyTLLFf862gK7DUAMpNPIgeP/6C/eaRBftle16aRP1+EEcTES
b+jyF3Iif+zLXkul/oHhicrXTCtmPb0Dvcvg9lRgilsi4M7bCyFj0IphavlP
JmZ8fS9HGVDwLnebPlMijHeB6QQ6gGTyqgpSt6klCkmsf3Ktb3d8O6WsT94o
lLMYQE1yDavY6ToVPy+OaDP4Wa4s3JYDsT6VDZJhfPgxE/qFA+fsLZgzz4/6
DIS7h/JEEQhg7xzpk67AyDg5yJJXTAgmmyEmoCwZcuRppS8FbhhGxXyTcHiL
9lioi1n069+J3BWfWrYNF2dDZEsHoJL4hd2bAouXkB9VF3abLG9zaGbbqULx
9+2z9xHeWzzW0HsCVvWWi+rcB7w3iXH7dE/ezwWDExyX5hJhLXquGBKt6+Bn
93ka1E/ekNGprVIHGmC9rxR7QkSUYDEg82tybrSsBFzBmI01ejrycBddELnS
J1crrLrcDHv1fvBlQxW6VDXMKQOgIwvket4b0LLUXEOOlAogoIiSct5ZYdpc
vHz0dOLZB01hCX4hNy2lovVszVyTVA3uNPRwta0iLa+02mboucNuiXbh/Tv8
3G0Z+mYosOWz/60tUVq5axu2P8FLl7z3br/C8/T1zP4tCt/rJzHAbPCt/kMQ
lmHdv6SMk+IUid8ltn97Mt1JaGbST0QlsgXpTSQmJ2jJ18OMUlW74qsU2mgJ
gu4bXbJ2eL8s1n8btpLi0wSkv9nzV9H5xoHuw8XySMsq1iI3x6twzqSKbav1
wqnAze1q7+5HJVIFKq0EUAB8Af5VqTVyvj8arVRgdsm71KjyoZ+fcsroKV8M
BCiJhRP2wuIkEDfKHAX7Ba9JjSPoP0SgxHBuItDPvSEYhe1U3W6eg8ayof1j
hW58GP61f58VzKX1rLSqF+vDdc8WnjhbTN6VCHNOCruuCdDOZo3ix8Z/qzy3
xMPDwlM/YTQQuG1SKe1d+sQmKntmF5bLyA/ILcnvoW94Rc0YvdzyH7843k1p
mrUaJbCqq8in4fY64CCwq2xjYuIJDiuzVdgWyP+BJUEESjNpf0Uboj1mgqgw
Sm4DPQI7oXEzDEocSxFz0lMa0V4zHwiI2cFt2SaWn0U+5C3Oe0ZvfUMjJwvx
wp28pUNcbgnlublLz+ebNlt+jXPK7rrBPAkSmI5C+Dk/cl6dStLyWPrOd+p4
yUE1NTGDY/lwBjrj2M8tDu9+WFRRWVUEdu+KpPTkr7IXAwV1jKDjJ2eaxpLk
9gGJswb2/ry3+Wt4bGu8fpzXULo+kBFkks/uAdle8RpGdm9dCpMAaK4gPxF+
ETesmtqhz8WGJJbBsLsVEaLH80wzlPgB8I2izD7WovRKJUVC9PYo2n1UgUE8
H97DwwV1XlDsw4BqETXEqn5tWchw1x1G0/m1st1e7G6hrMYwq5E9FgIOpEbf
E29CQD7N+8jfBwguzUbNGeulG/NaJ+0xL75GMhUwTALmdLplqPFPj90hMZX1
o+nr252VxRKUQ4ylmFX3K3+kgBO+0my9uXWZm/uJ2xRxzqAslIUTtJttah1T
PY0yeytHtPBbkGuo5tUV7R9E2bMZUUwzCIGov6L2tdYEFm3Z+k2hrSlhpqJh
Nu3MaaZR5BVhr5GVn4qM91MfOk5ELTJvZGu5XYGUJUjbqpCKTE2O+nZ8Ty2l
9j0CySdvb+to8iKIaNjJIsjS7FNgPopkZx+riLSJfW0s8ZYWgr7jc/JuLwe9
W4/iTG5KexsYZ7OpoPZGXfSBmvbOPJ5KUDnysAkPPGB/sc4+V3PhRA32Q+Nv
wTwi29uTd02jb0nkaPREQbzKfOdNYY5dlCIMBe0hflOwZgJKz9yK3bmSajwg
2MFsVVJUboYsMYEp2cA4jcjIxWN1ogCWTbgo+gXYBwTG7lv44mEV/XukQ4SM
VPTdrAvFfPgk2V+9bW95yMvfZ4Hcub19tPPJtggIsfBxpdm7G54eWgIi+Uat
c9AdQEBSfPJ26cq5quotUUtNS9dfZWGw6yIHzCR5hAZLXaKn14AHarndOKuL
ElR7wQMIaPfNI0KU5xN/UT+ZYLoCeTCVpaPMGJzaFdBezkm1UxnmJjYYeduO
ZwxAnfzrzCEsQX06hoZkH46KG47cuilpo5vFjxpyekmIYWPsMdE72/FBN5mN
mDnPsQpvOtWV1gT/IhJLHvng9k+sbyekWnkRZ+dTXF7iMiw9+r4bSnubxjbW
0qSJhO1UdIzpsLPqCx/1slnHNaEt3GvCBkFpOKqsdTWHaLcfr1rhXwmz29JV
8A7otPFl8k6YfT9u2kbUztkWl6LuNgbU8qkJn8LlJeeFmJGrRyqTmbC2Jy0H
D3HvdrV3BMLPZRIKmOvkhAFifPO8UPyBbc9ykBs4fjJdHftR+hYGOJmqtMOw
Lz86PK6/I8rgnlQIMWGLwRSk9Iv0ipAVqqCum36S3lxzgXs0rUNtzDUGL072
ubK75eW8xT0gKhRxpKjI0CA8+KAiWnTGVsfFg09t+68RKvyIWFdk+IHgEFgO
4/lEZBI3TJva2YUtb0V6ztQSVifwIOgk1j/RCdBBVlyIgGtCWLh7LjMVbb8e
eRLPTboPuSKOrNK8PoLsQ39GpnRZQ9m6OrZcdXH8yN88SfXWLafnl5Ci3gTM
RZT285X+TiIWYipvjjR8UMYOqTtrndkN36p+wRSUCIZuspPsMB64bO0YJ7R5
M0qrQ4E3lrlvS/o60MJCmpxlUQ0/0X45pAgEOolM1uxgC0YeaidT/lQ8kMHx
GTpE02YWIv9f8wmj0mJMg2J9skV5h/yB1RviYbufsDbjeSKYHYPOaZB09eQs
PkYJdBDTf84qzpBHuWxLRitPGFWrLT8HMmsWp4hfRxVQLPyV0cKzABhyZyOb
KDVphWygpeT9upgh/sf3Z3mHKftLZdeqsGorOydRIDeJ8297s43wJm6d/aRw
cG8Ry8IThKbnWasZ7LqLu5eUW0XW47+QUgA5pFbRwtCSZHbT7gCFXzFnhfug
ep1t3sssQ8FehfieQRianyAmk8wGHVE3YS2eby4ymn3/lpk/QSwlw7JDrE3k
fthQUzBwkln8D7YOKwocftYlN22e6ennxxJ/Nc6ZhwIUYVzFft76dqpHjdBL
UIarYSvGqZOhzp+9INXKXwcm0DApnl0SKYMBCttVg8+ENWwRrI9Y2WJYcfdT
xyFWeoXd30HSIInome2pRAA2Nzqv7XjUNVkjkJ7Qy2wYGQyvdc5ZPvNvwQEs
dSzE5QRMgVBPPSiOPgEYWCQnKDIgBysc6ogvGKIB55wdGR9nHcEDNod8z/Pw
5t6fLuTeY6AYUh3P6gSKrviMgw3q75q2BYvGjNjncH+JZsfiKf2BgAEHofgM
NufSi2T64esSzL3B4UgEAR7AsAVCurXbKf36vmJ5gP3QLbEAl+Nq1k/Mkqj2
oGxBUSya60cuU+zMz2htoKauOxLwTt8Mdas8GQpuNfw4VsiTrSVjE6Jrq+NV
fJlTT55svbe1ER3jRwj7iotpz+pkWI7sjaChSekDBMIUqrcCurQwsb/thPRl
fnsFb8jTJZb69ITvVLzf1IgxmjAfn9T/rEDCgdWMEs9nfpWm+bWdT+sY/u9S
VXbYzHR43c6iI5iG1qyyomPpQ2JPjFcRSxYm+LkUnz7vV/VW+6aOY/nltiCk
Nkv7WNcVpeKghHY6TY4Z4ffldbZkzPokEWQdHf5PrbMbVW7hOmBFWA93cFHN
kLer2GBCKc6KmOAgrDwHLapMFcHbIMJibwpW6sJ473w+saHZnlJ1omPGvZsZ
c/yklzAIqQPRawFA5GfnpExf6daJB5Qq4N+Nk7ZwSwxIOpYLWNa0xQdeyG0E
uzZIqkyQ61JmVnhV7u67rp6mqvdJmCrRKYAFWgDGGabowCUPpOiHsndkiAmS
4ermy518oUcNB79B9DQ5W4bH/TZEW3Y3zcAZjPwCQhh9759JBN911lVPrtKb
6IdIMq5RFntVarUJYcGdCTMoiZ+q9JUIaFyRopgUf4le+CEW2AOSgeCG+RUX
R1Lfn+3RnS1MkkCv2CttHJvDwp1vk6fgPyq2HZoXrP8Xa7lKyeMJQ9wBvIaj
OpY1tORbxn3l4bK5iKv8qxTS4gbA7YHoaMC1paoWvpP5xhTwocGIAYXVreNG
Q77RgcTElinFjYIoyq/n7ZWWCMzzxIOWqQraXRzUyOEGguoLr9ynaaGvOIbR
QFF3vg7+IFazZshBqUjXfNafynR5F7rNY1cTUlj2wjXMrtnc5gwOsXvBIZ22
LTNW8tSuSHNzJMKn9aJDdZc7NeSvL7RlBD3QJN1/upgn+6i5g1NrUp7lq+LN
cz5SYMGbg+vQc5NErMGpR0uZqVmsTrHXt40To/xYG67NB9lNm5m1mg8eL7g2
BLlTqkw5Pd8fcLenv33OZ5EDhMZmyg+ThAOvtDllhaR9hNk2yHJMtUSGYE55
dmB6Se7MZyI2fQw5ddZuqFrP3yJuCjwPoaLBPTzKBuzvWs37qoS1wpyXfXb9
9tO0TS7rwUZ+2Cn8zkzxg2KQNdH1cT4zdwadhvZ8nQImGlC3NFmRwbzYR6kl
431YDnzVRaZqMYTX5ILgdx19ivB98w8qYiQSkqxWshFe2DuG0fnbgSFZZyS7
s6XHRAA3v+dYLSPjzsCBffq+bCpoKTLalnNvphr4hIsYhmdl/2fGDrE28Gnx
VwNzwl2DuWo9adF2jSTnoQONEca2JnuzcmyEhv6rUfoMaLWEA9dhl/QZZkrK
Jn4+yDz/FwzA38NMyIv9KO5dLIfdX6ngk703thUBsJoFDabWWrAgPVZzZ3sP
RGc95RA/o4lTXM5WQSP5F/BBKi7FDM1KmjRfMOwtpd5WFRmGSDOsX7EZdop8
FGabDKuLe1/rSU4bX5m9gkDSCCNzIQWuEvl+nGkSPtle5ayi040JNoXoIeeN
nUMoMrunUb6q7qsgHJEaWkepcyW6HDqfHBH9rI1/RN35qSmXxek044auv+nZ
0KWE5ltD2hUicwQFWNQ2R6jXYX4BkbQ2Pn6P1MSjzTNFXgHckFwF6/F/JRmQ
IqesrWKAS68SpYz3Jt0DOxpEOIj67BRnHXoiRLHUQSykIfM53FyMoQ5NccF4
C6YHQxQDjrb8ewTKNNYbY2ex6eOUhv0zwqyzCxOl0/aoTF1e9C8ibJ7CJYjG
wv6HUEjtPfyvYV8i/jDXPD6HY/+MtDb3Me6eKB9XkIil3h5dQeOnNc1U6xqC
NcwviLeFYN6vh4ihFwF16TupeN5CKxBWqluMHgj2qUZ1cHCzdBfpNghZdBdL
lzTZGU63YSDwwha/XFfeVgdsasHnBjBh2qo/wjlTJCJiLc4JJplfklqdRPce
5W6to/qEOBarDw0LaElX01dNjqB/Yj96OPWIip28mpFiAMj2MecVidwsFxrO
4Jehsflf1GkjwtYu3azMpCdURVkszbILOqD1I8rS8fWncBO9opNDNMbA6Psq
U2VNwgo9GuXmyDFiLRsctnjVWg4aNo4WamSd0dnHLJa1q3xi3NDus7/m58La
tRJOG8nOFI5+LXwzmmfF78CJoSx6IznaKul1hhYtRDa5TbsYVvknamxvtUcE
Mhju+9unWZoTSKI4ivTLIp8++8WUefkxeYmbrk5OI1vO3kw1+qw5lImmrTZ6
aDKPDkliz8NzrEsss0rpxQB7hJ6MBm+b34PNuLwxh8oadmzz6TLW+khupob+
4Cps0uSKfz+Xc8fp23keFt/1WN3k5XfXtvJY/ThyRX9zkhNtJmE8VpfEQsxk
gyADTUKOOPCXqiigT9XVh2QPPqFJWRE4Kp4eCqM0DaIidUH/W8wQ6YAHjZXm
aP2Dv55Mneu/C2RMOT/QG7sKH3Nmbhs2A4Jm4d2+JpRykOnPtt9MEQS5RIDE
A9eazvbd7PWIzz/fMGdQ3eKUzLwTpov7UYueAClDIpZTirTzqoSW0g9zqcaO
qmmg4bdO26YPvAazdSuKUokCYnXKspJipPo7mO0ibwUUIA/rptqNwHYxFK5E
xsnE/MHGQf7JIAjZ3DONHe7eW2hIgPNNCglSdA/Nv8TIqS0u+3ihQEC4/wOY
aEJUVjbawrD/LbT2pZMtkTpJ5VXjW714uv3dp7ak6M/Y1ZWaQZ7s7GoougVO
4b0wPkmUFwEfWPzWY0TlDGeVaQYoOJjqMM4SMd0dWbqKQmbwaNRzdeQ5UTTH
t5ktrhhLSBZ6C+U+Xrs1Ig6mZEOJTrkzWsKhNO7aK922XT+plPi9js5KrpL4
fSwRlURaIO2OcZXMSPXYacX6wkPfw2dSAj76IWpddeGTVttAaK92V7OTOS8C
BkLqpSdh1X7cHEvZXBERZNjlkw4ogiLsjJohUIGRXAgVALS9zRt9v/yFZmQn
meAYC70AFadCP6KXQKXqOFgjLDLGkh9OutRl/hQQQ9JRAhalv8ygXqvS9Wj5
Oxq2Q3WmPkmK2SGPYxdgDwqoxrgxGEGZ1C4GaUjl4ruUJVEG0ZprWmk1C/ZA
Kzz78dn342+ChpZD+6nGb2D0PqXAfocmaf/SNIbvP/7PlcPvdwmnUOKToEAj
E+/X4oWpV0n6ERfWqaEdAtZORsJJwVUQoPeYLFx09SlqOGN6t0mYqi9a6Ilx
/59KUysYyutOnBNqOX4Q+0hgD28z1JY6nIbYY7Ou7UY84dthWhm6odRQte4Z
LJMm0s+Ju9qKPWmm1SkQwNvSINUotRucWvKWoZtE13qYSkLsk0p/mZ2SYrj2
AwYr5JQ0vpPmA6kZdiaatixgjPgqCA0o8D07OsctbBz7smO8ICDebopSZO+9
mOXCch9jvrfJ3WtGruqnoXEEHJlmYgMbtYUoQMZkgogHU1Gh7oYmj2sT9Xvb
f70qtidH0e2jlTf6Aatx8E5s1fR/yUar075Z7u6+MuxrMVVMusJTFzHsgadK
Repwj+lKSL+pJ121+Mgll49KUhMmTxe5KBJAfRsViOpL+PJ+fgl2sZwF7jk/
PdfXcEArdZfzLSNtN+YeJo5OFsqpaxEXnH3weP+nLDtBRGYflsPkMz5CE0Og
pLRxwEPYe56E/ZV3n72LkhPiCWKN/7vRkGv415oJMFn7OqXsXAeEuBdg+Tgc
o/fy80HyUI8RrMlyVvUI3iztK3qFtJbOKcNfRkdOaxVzjWqWjCjAgiZIdQQC
BX6r0dET/uY489bzpkacJMWsWvJF1ajmdYgNJsS85rcLgHOs2zqvpGKPSV7B
AZihNsdIqFCgp+45IPnrNTYBQZDVx0qSPMePDS294J6yi0mRlEvzzc9sYagk
r2TSyAE2B8KT9aQ/Vzt+lOJtcNnJrZ1jd00z29SFtqctmKLchxUvOJ/F95bM
GW6cpZSEaG9ZkGsug2YTQxzrFLinVOqREjUtT7/tBlUlisHr11ntj5ECqLnT
Q6gIkDgt0RHWMBtzpgprpfyIRIkxQETO3WmJrjtzNAS8wX14NfpEvwgBPHXY
vGs4OLuY2hjBDhmQ3/Abb0W79OxnMSp1WAWY114d3vx7ZoSzJ4MY5Gk76vNU
snZHmXaKtjFa491mK4OYttoHk4cFW5uQ4pTMMcw/tJeprnHMZxPOQN+uQdMo
2WFWt0cLLUsfTybOZ5aKWTj2ks97O4hBsJ1wKlmKK1HuoG1b69lGb7l/dFXk
YLPDGEpqjMqAkIsJaalO4zVrPL9Dc87tGmwh+DU1vhbo2oNKGGjY4avJ8XrI
e++fNcdqhDbgmU9nvPu+WbXTfcWfpE4je2mPRBE2Vi8tRrGpJrWX7TsV7gmK
Ta0f6F4jY4/16lo2ADwjdP+NUUmrKMwh5dsomS8tBLxAY5/nB8skhltW5QkI
gzDBDSjHI/LoA97xH2O8x2WqQ2ye1SpC5cZMrY42vx0yVdubsMvOFnYe+OaL
uHg558Yt1ZPFr+yThM7oN6n8eL0MXOQ/jmRvMDfVCMSqtV3DwYBc7rQaMdJQ
9wPGyMHLUOMDpl9tJOy5GHoKIp5qRWjggWpmB/MLQscm2YXKoLHrwGokM3Vm
J89kHb5Bjhfm/6qBmlAd7dyMEZENGWywomiw8AktSCk2ohQ9nyX6iInMqNBA
XIagMQl3PG+gSsONdQUBNMVCpVlbY9K+mlaI2m+RjxfgOSuKGQQgq+sZWJ4+
wXq4Z7SZl8gK/L1cS1niKf5JiWv9IJf1JTxG1w0b1DVDzEKEuuxQsmHnQ1Se
Aqmj29d6uwpPdkbwk+yLkjZOf2h62plSn7jOLYuIej5RG5B7Gtw+QRWIUJye
4OSwAvzTlRCMmTnNLQvbws7EMcehnTJbz7jkGV3wSMPUdGS07L4jpgXCB0kz
ucRnPQ+dnDgGKC86qjgqddWYpec0/QE5uZiNEBddnQFVjjkElNuDg4Qs+HK/
rc5XomPGcKTeNvekq86U8cykTmqgQhfNjltz/+qFSfhVHCU5Iz/uRy1Ua6Ji
gEKUgc1tcb+yNz3Nya1FiupmlLaVy2RQlBEgOdTE6itzCa2cw4Z4qYzUwjx0
AS+H1R9fE+tfED+92sk4bYAX1OrSUH22AYxaEvBd93jEMgyPGPPMMZgOVbLq
nbxUhGUWFc5Ztfz/BGLcu5mm69p2gQnIVFFB47UkOYZjIkGBA2NK+kGf8wjT
o29E8+zr6ViSLS8KwqYvMctTDIdVPwfYTNZBkSMOqw72AzUIZ+1oS4GH5Uyk
7ISnj8QH3AxkuumQGlHrZd/b5lWfP8JfJDCJLThZn/Wn9/YyQethtyQu1HNg
jfo6AlB12eUQyym8tsmgWgMdb57lPzHn2RKCAyspbe8mIen3/lWdVSqNGGHa
ocKwnt6e2OFQc9m/Dz7VhAg+7EgLD+iqRFc7a/FYS/ID7RgZQ66o5pXMziUv
9UUWR+UifWSG89IIJ0K/ZopCgY7XnUg3aODgV8ooQY1Au6S9pJD0EX/xAhY1
uCyZN0MH7fpBkc2/AzT80pAgwMQxjcZGESJYeRE5Q6LmVq+i6AYo1IypIfr2
3v8/F6/XubkC0L1ATiIG07yiu4OlMtLSjYuYIc8cwvJgTek91ImeKvd3uWmX
hEi4brm1fiMqxSq1JMRO4oW8qg6iZdCUaXQCv7Ilzbappgf4Enp92fTQHfNS
H1oU8Gma9R9o+kUurTnzqOHZ6U/RZE+cYUqMbkc6+eJzhh2/8Wzq6fJNvSRe
M3uVpbQAMdG6m9d5v3W5eKqwHRsxCtNbVn22u+d/hmoA/BFZtjbkdazWGV+d
oUWg2gmGfCMk03I+ILTp4Kdy70bXbwWJUJUy1sZIGEGVVWkOs+hovsAcnTa5
QrUGphYEYqfmnXRXzhtV4JzBcfs/IyPvFTu+V7sS++G9KCLwbv1rDnkYBSig
CLzwJCJCD0cz9GlJT5by9sJNH4EqejCaFSdLi91Pr6sTCaBESCRHIBLcoJlT
Wtqvr/ZoHiKpxEbtIwftULuIvoTTX8KbfPYvcHYe3HUzspSXhbSFELgZi8O9
Xf9UGahTncQ0Ss+0Ibld0DgVUyU4mO7mMC9wP4Mj6tqmO3QFMfPyWBEirAcd
0y7mjEBh2YcKZa3uoezpLOtTaU0C2QqZrEP+QXdueonYfY9gSyswdQm5o5YV
XMYxVaiKtqKs/IRkqaJu4uq+HcfFwBWkJrf+7m9GndXBb9YACltawYqgAUp1
ncgVU0o3yvDkUx7vrlau/YsfOPn89gJy9wYMGTusiBlSBKr6oxPBTAqELeuK
apoAcDj54jPFPWGJ+plFm1BfaEHSjKZzHlF5GhIvbuEVcenKWoJZTOW7x6Ad
AGfMFQPJ0z/bpcS3rhBj3FDMl0wPK5A+ZsKGPsTvre3+bBHWRoQu79WZMqA/
Y0h2XypRF67R5dhSZc6/gOZSomyCffCGuBrghMspW9TSzOI7e0D5ikfW0lgo
iXMh5NePVee3lXhq+X3TA6WZgGQYWmyIAMu2QunJMLQYqphqN/WFpTeTju7r
40wqFz89dczlN1kVYRMRfF79nrDlEE1OuGHDRlAwl7fZ2tkQc0+jP3RraWVg
TZ127pUE2zlY/iWe3p65Hx1hOnKTzWVHj8obDRNOE4quaT5EVGQ8RFo7C4O/
+DSjRDBp5QJHulYxtZT9murNzL8uzW2vh40Ks2Ha/KBcWFhdVlALbuVtXThj
Xg6qNRAooDcEaKoV3ewNIRBwHE2LPA/wn44D/F96xsIlhi5o1Zz+twn7MmSs
5SCEXFUjauphG4zvwCUoR49GszZONiwBt5fQJU2Chno2sMshb9qyI4LSPIoM
j1f7sW1tSXFi7OjeiSi+beElzvmY2OBRLKkFTNQ83wh4WDKPee/vZklrc2q3
GRTtrTzWauqCj8Va5KAtmZAMUTbYxmbTTC5XinX/W8EVblDHTPZtVElVA7WI
BcypfsDlCBSBK2RctoNIfTDKkYhzZVUV4we829qrGERNGa6edKKkXQN7dHUN
6YPZ8Q66qwSgT7aRD/r/3gR1GKwCdEru3MI2nxrmo5bezyT6pOmyrurTUg3l
8KimBHnVbg9xnG0cuE/BEsVVmyvIE7QtaOsqx/+XMeolUy5+HDkDvpqkqkdA
LwawmylPbuJATacwfJZxujTmoI2CKmpX8piCediVzTsyjmLpIfYL/hbvhcMu
F/djYdZx10h/lB7A8k3nSZE/KqNZubB9I8Jm3Tiird35fSlt4OEpWggzhPFC
/gHZZF65ErwgvXMOwNn0OddMLPEivdxGilJoDKf4uuJOQrzsT4r8F+dQpPCD
/edO4kETZpjxL9TmsFDWSXoOjSnrh3gZpA75pDcFKC5TRMLVyimulecAs5uV
2BbSbfrC/GlnpXXB42WU5mk4Kkp08lwBOx3qNV++5EnFkAZ7k1b/btLwJjD6
WvjWHZoDqWTx0rejzl28fqU3Nlrd5QYzBCPjsQB8T7yEnaRZDx8JDPERrsQS
rlgUv9XvizFDGW1020jaxG9IddukyX1kKusq0+ELVuTK6aRmWj+sc3gD/m3y
9PSG1J56DWA1+Z1WgY3NfBUSUPISzX++txpTU3WCBDClDWDdwwajFEJRD2Q3
0z2moV6hnIZR8euCE9nVSBWPK+NHrPbruTp4CFt6L8hWD+VCA57G4Jbr27Xv
T0+ryNNHVhqqtAiJIpnFaVm+L5+d29wkFJUy9Z8ZFC8W4O8ipkVxrWcTrRNd
vjBwkVHL58HAuVqj/OTDf+k7I/dNGfsMMVGjdBnKUZ9VEWnfye+KJcQ8BLez
oibviqZbJwOtylk8HhboZr46dREEjHpIc30MOnYt0jYxmYDmnFZokGRVjXYr
2NL4z/Lrrchnp1JXBuEfnbEwWms7iQbW5M7Pa6Fz3NwqGOxKCCHIj50eN9bR
lLHQqwGYu6jKF62sALWmYsZ5Ruz3+y9cLgU5zejMeUaPxVLeorNvKGRiH9du
Xl0i+8iaNy7JuGj0wsy81CM81Wy3c1XAtRN2GhFsIZo5KNlwwIYRvQWdMPhP
K4tl4dCyenUHtS4cuOkIUKPBrNmO8N14WKXrJMbIy4b3QwjP+eQsDYDUnS5P
i9lBcm/R5jzVH54wUmnmTK5D1Ce4j8XQJKSPvpBcgRM4CRN5W4VfTc4lV/1k
b+RyFKhi+Gozfe4/ArZ95ruPpXCJrwDip//c5M2ZjUON22S3qHpd4DUh9nnh
g+zBlwGw8RpZmzOnsoamp8mGQtG5sgYGeBzwdeqqZWber7cD+lplVYecGwHf
iDaE61kQiBTVpLBwRIzXwui5WZIPqpl6jP6QC1tGafy0QPjKs0YRL6IjUHed
yORJ+n7Wj3s6Pmi/Il0KaSgpIXeyX8dBV11I5NxO0V7HX1ai3D47ypUDzXuU
3ZyQLkGnclwgvr2hJRKry2E636kXj4GuCy65zS9OBXpRJStE9o8Kjtw7+3FW
6py2eDZicfZGzvTHlm0aFJRQ0TS+Dm/niwQlK1DvUFCxdtpzfvpdbaaca4C/
AZN9ZL0Nrg1eL6PI/jmqLrvMaY8IhWrBKDQaf8doF4cMzeCgoEENG/zRtdHc
aQAu/Sq8up7s1zAVu+QSF0Ay6+f95EZRg11UtuSJSuUm4V5VVKpWEJ8c3yLn
pu/eYHff42120x/fr7S7ar0G+23i1eCFcO7a9R51D06xWzHebAUKUG/Xm6B4
BJl91eHqY+gcTbEj1ChhAIL0pnFbkp4HewnvulAMHIqV/3DsnV7E0DCWJivk
V1Panp/+s31nh0aQT7MUNh03aiDxVdzgJIES+WO+xzeZozLYM5B69AemMwiR
0VBmmQUyGWmhj6KpGSMx75dJzaZaK4Zs0zptWIExUy6CuzEpBSrUNoL6AU5D
itKRSAoU3UuxYAxf1mr7eWh+PBeqereP03hNvSFt/fNmeyetTFWwODN7PBVr
5tpbCYw/WZ2TGojPiCmLxu21iewLGaky/ZVoV3WI2iRTts3F0q9hbcx9XGH+
pL5FFxwX91oc9kpmv82FZ54N9FBsVl3M+Pdl54muV7Ckfvpiqqal6psu304G
Zc2kl2f0ZSelTpWL3Xx4qUutWtdphwdFtM3V0CU62lvQ2DoNhDiFgVktkXQF
mnTnVDbabyBrLhxK9Wu3ibI4hvYVpy0hOHdziuJR4eCfyCHZtxMlNjnzq9J7
ROHtotyB3nL0bniEdGoDQwhIE2m29V24C5i0NPLAzuy5cw5qgeGSn6ltNaZw
EMd84fPo6FBokjPd1H47l3zCsRtJWc8lAjY0RmgNfyzTKKN24YNwnBqQqOHQ
QftDhV/3Abc7VqDAez8yOoJ1Wih04n2x5o33zOOx+RwamZZ4df+zIs6JYHvo
3+iN439O3RHNilFP5HnkoUPp6VPiNkpnzC9LpJopAX0AnlCtrX2SnF8OLuOn
b3hVwxk/rgPylVio1edOaJgFlwyUBA/ejWQOktUo2gejtagTlifvaQyO6XQR
ug59npop5QMOmf0c/CmdWTSHjEQov3g3y2rGuNuxGpAfdjPNVYMVyTi4AV2U
JtEDkxtE8zDEWFwDEAmhnMT7g8pnVA8a8xKq9VUlXPl3vJa1REhK78mz5mew
sQpMcrxPuUlhxrbTvgnkL4J7O2LSJxPaC+TWje4MXq/T9csqHLD3BM8IbBRN
qGo7Vx2maxNHyvCls30cY3cISHh3ToLBip0laT18Qr6wGgJoe7W5kof/9IKq
61A4e2LSbM4WF1aRFZut1OOLqETx0ERiZVtrbHvVtKZ8VnEk7j7IXfi9zfY/
Qa0gWP24EBXiXhNwB92Ezu9SKTwwXIm8qIPGB66kLqKgtJ2akhOrcq2EG9zi
/K0jT+9MSEikE4rY737WGLLz+M20JZrLQWFGcfxPIUYdPNj/pb4o8UPNLlQd
gOhMKOWwmYR0b/LVkZri7mDzukuN7ENedGz3BUIgzc0XfgT81wQXRnSzhc72
9AbTa5NGCQSXu9qQMt4gABqLMIWnGE+r9pYCd0i5UNF2WKGRdQvtwVLUL6Ue
oF5DMBY9Qq8xFDsy+iac297bdG/8Q3DBL+BW1iSPnM39oybUZtsZJqWUT6nv
AbQ3okX9Paz25m17EN9J3Xd8SYKcBLiJDIquZkn5PE7mUhj/w70gyrf/5XtO
zcLCNsy1HivjfmJC8o0taE4uyeM78YXad0AL+oJ+oZEp6mlIYd0RiroQqgOD
PWYyObGmK0W0wPAA50dJ2NxEwc87Z+vDB/MlghLrxmJVhesOm3MVdGfOYUEE
UNka9tCofwJEQD7BDhhjXrUjMj2QDeQX9N+x8CFo2qfIKv+ue1KTG1rFw9zv
aF+OeBbFB0mrefJ81Qink7izF+ZJ4cUzoQv19o8AvB0KK7idR+DfqsAbSp5S
fFosGiSeJZdyxGBgN8q4t7CwgEWK8Eua18z/P6L8Lu1rsPSDLmfqUlDU5HoN
UpWq5YXWWVu2HWv6Q2S3w6ZXuClCSDtmfbmyOiZBgzr07OdpcO25vsLb9ZXJ
S/1Qj284Df0dTXtlte5sKsYI2rmb0QiRU8RKwJVubZU/qK60chIeu/VCNBW2
8bvfshaVSvAQB2itFs7Y+wg95PTrKb+e8/G4cNOp3OuFuUqzxdfbwCuZVscf
6BYV5vsdzcKIpyIUN5+6VgbPrW+KRws62DPHTEA1PDRrx85yaJS261vv2DZl
X/4DrxQ4pETf3xyM8/LkRmeJUq0GFKSzuFg/mhvLEhAQDTJd7QSiF9c85ZXJ
nHP635iy2F62p0pcIuNI8m/SKyRCoLwty5C4waua6BPp5sRjjXJ6ZhGcxhEk
PAK0UWWheSTuNlWqfLZ1GCxVly2z35OHD6A/+LNhoqq7UDZfZx6kZvVqbbTL
mRr6iBFGwf1l4gV8K6xcWhZfOZ7m27A7UNL5NJjm3GS/yChJyjavkuRDy+cE
U6y0ZQPWvh58jbPYVhhuvYDfXSPGiNa55Gf2cgckvCpZYxpr1Hsaqxjpq7Lc
32+QCWswTAIWTGLYm+ZGrYEqpk5tvKvLZ+++BPtOQUplj6/u6PmlIonrACXr
I0T6sBmvUrX1dqTngaL2h+lsB2cciG55/kZloHcSjHOjDToWoArzP5JGIEq9
PCXs7nGKtk9HM7IJWYuGNByDtBxYihdefECilcjLRiTzn/HqquC9jv3Tn3ck
WFGEGUHznGIuV4+qjNOWipflqEZ4dUx2mEuomDFK8BObslllf/Zv1VQK6uCC
b9MJQvC6EtQ0NQm4WIJhd9od7op80R+hu2Ir5Eq9OT4Hsbny5hXBA4ZccHw2
TRqjz1G7KqCqt0LUKR73dH+2TuhVENGLfGNSEgmgT6pB7TUx/mrVRd2oqGVQ
q/xh0WnRoZtr4niiQLQf6cfU7SfhKelZv0YAuTzwUJzsE6ZjrnDeHRARvAC5
vbVvzYq4AoFKlXFVlz/c1+7IIjpEBZqG/bPYhaCD0J92aD5Gz2Z+3fdltZNK
KQ1DSadn/LW7GmSdx8evUhcwUudawMr/Ky4VDXwsCu5YmRZHo/7WGSlSEX59
9WktDIFB0X8wbQkq0rc5JIo+au6cYyJiznd2nXdahAUCrMsDqIz6CwnXZaM3
K1hOSi9zGUxpZdwvYcndVCsa3gQN1aTcB/x9BkD2UtFE2NTT1JGtFXhYc8R6
vx5r1yH0n/fqYAsh3CZha6rYMDKdlTP7kkXxeMOFkcI6N8vpKxlafxcBTW5P
l2gwWGRuWtflRx4dvho869aaYNt1SN+s0nHqaSw9W41mtUfWjffG01JAABTl
MNNIKTQeT8vjEke/xaNtU+sXeTQ67TgKtChcV4yr0xtJb6ZrkOzbtX9Ke7nN
kOyimJQiOuScjH9lI0PWJk+zW+ntKYSbQplVBBKoV4UHh+R6akbm0cxi9rFo
wfPWV999sjXmONUf5Vc/6Ioq2IjmPvcjqNZ19VO25IoSKXawFqn10eQABQ/6
n1wt3+PePWxzi5QGIBdi21HTvORQ/hMBXgk5zS3tXW2Hz26YDQiJ6GCWMacj
EuyVk6KxzR2hTo2UBgCLRzCxJWIi6uPfoDrRJx2eWEFF/B2peMom5dkmx1is
UWYPOU/zy41j2JdUHGAoEIhrYX0jFLB3Z0yiptdE0im+MzpRTAsWTWlxB5ZC
L0YGo0rYALzzpjjwZKehRUFOSE5dgnehWBwOPOC2M3SlZJMJhDoM6sXwY1Pa
S0WXRuqPX9eL4x9N1gHOuK7KVnWog4qhYJESYqx3vkQh31gvfkkLx7bLjhXE
iwjc9lofJXEsa/Ep0CORZ8KR4zuogie0eZghsMB/AuDigq4l0TndjScKZp6A
lTRO20pMf+vd7NmIUSFohd5FaSBLJiWs2X6VbbsuNxxmsSQwTuG1j0ota/T1
6tGKnIOQhd29lbkZ6Id3lFifewJLizmEMDoB3PLRCeQz8hRKRsznbzA3PRK1
Ra1VNA52PKZsfK7GAkeTMOLwtg6KCw1oLiBuUXXi8TVyggH0GiC/bnmkIIXC
mbNxgpClJrPXERI7gB/QaUh3/J0kcE+L/2sa47Q0RH0WGUeRUkYPrmu86qwh
Dz/pTRBScY0CRfTMKT5hkBShg2Dmb7iqrwKg9xavEH4qox6yGyM+C1ze/H7e
VHMpy7iX53FYtl5gve3kTFfYNhkanW9GrffJVu7eUt6tO28vvRqWdFTOnqEB
n8bg/HhaQuyDiADAxdyL3Ust5VnIt89tED5bimYyT8qCt3SxOuUJWFpKEZFw
3irEkBdDZ+35ODdU8WRXwUtBN+8TSPy0i8ip9OfwN22nwQQIWah2/JlFd4GM
PP9wssQEayaf7T9r1+gCbxNb+ucJHKW44ubk52QtoLRRyyk1pRA2IgXnJljP
rzpzZQhoqOv+41dQZx76MqcF04fz4A4+nbvzvDC8dAYToEcjAOZlkvIQWya9
tdcTi561Rm3tp/0/sUIf/zFBP1a6cGPNTNwTFwBQ5+QQ+mib+AlK8hJukV8G
U+Cnm+wuckqpEu/zaw3MPWAAvfz7R44aBvU5CWos4pvN6Y0+MeQfFiMELgmx
8h0xPzSD7JxJ7Q7ozH+rclaGFAvD6lgKM31Ml2jgqVcir1CtJ2I19lwfxHYr
mEdUWiLb7D8jCQ7YDsV4IsAcVkxC4DhdLOU/TvaCCtgXH3ywwptTueXXklGh
SXbrra7H1+XWr75Q2uOWwCaWYC8RZF4gjxwmgxAE7GxgnedNjGiRfy6A+e9J
dNA+3UtUIaPFlY+/pI0cP4OZCoeg+fSTbcE/wFhZsgYHVP0vTm+ffxKsm0yH
TJENm44lk4qOPpdoMfKFlhft0rRK9DzimH9NnPFawx3fbhJ0ihQ3hShizmgv
gbwUBoOAdIjCbDrbRi4a90U+ZB1EhcEDx09jx/yhCJtfqgRgmVw1aCEj7iTQ
dOZlCoA6dBZf5jXechB0o22Pvdh1ktkNGcugG8DN7htxKsoI80jnmgq/pti3
smuJ6wKKxyfCPOgOEQCyXSObMyH8YDBUjlxM/8rQHYStpTU3p0X7YKxLx4Ve
yt9C6csyd4POYXm6YJeV1nL7UbVistzvT7Y9/Pb+zzK0HvcMOaVr7PnMmx47
GtyoFD01+anw/T9dMyfFBLzANRd8vpXO41BSD80BkQr5EuAZbKxeOPx9jAkO
/MKe8dQ/5Hm6XjEMWnvMs0vfzBt5ksTlBXulR0X2E0xsm8Qt04lRCYB3JCCP
Kv5mpqbeFm97cXWsKCfXkIgXIafLMcf6y8tuqJc3q7DdnsmNFha2NTDQ4UAV
SZUZOjqKXBuC1/cBb/vvIpcVolVOe8aj+QE0988ZEyCNdHO3ra1EY+61hUMc
+p4Fa4X3UJqjyrvt6TDoq+L4XTKO8HWjDewfA/yu6f+0Jpbdjponk2qumutu
FcxblB+R1RWbsD/F3Ty8l6wDRHEAIOvxfT5/cawVkqM3ukCZJOZf8fpIvIWt
q+jpkqXCGY6Iyg6DmNMIMpXJSRv8Vu3CzG5la+6EUX8rqZgUNYdc7Wk4FTPi
pvjpyDNJwcypiyXKmzQw6y+RWXGicrm40yvI64aAa3jHSw+2+9fKyZj7GiuY
MNEpG9075pCiFYLu0Cz+l6IKsiDQtF2F38sdlvvENZjl3nbTB5KvdYWPj3Hc
5HqzLD68TfCma3PpZE4KHrlmt69U8YNhZoetz6/RfD/Fq0MKmgZLpKRsj8Tr
AceKGsbRPJbfA43GNeMiaXEYO2kBWkJXT6UezpTrCMeKQVOPecdxgIHc6ra+
0KLmdJhJOKEI1u78+z+GWnaEoqgIVnFoVt+CX7equVX6tO1kleB5GhDqw52f
se9tPQO3bXQldD95Zp8sPDouO2cAsEcnHxpuqG8qGU/6gJuCmz2xchLKA4iy
eICvcpZbKvcOa9ripmy4/nKnQOMeuZQjQDGB84EebQ/PAH44QLuoRKEeLezv
IXhx5v4GKdRTDqRqpeV7jFShyS8qbToHYaCBpLB5zgdjcJBWQz+YwNNQZujW
b+RwxIXuU5UJFHcQyiAT/QXSQseElnAVBlFrwLjssKLSRP9U+JoE+InVdCkM
XN46b5eOoP/U+0qZPveI1NV4e4WBlLhQTDCjeGAbeKTkD/WNsRycaKcuCgHn
r63jfb0PDUA2WzhOYM2h9tLISPc2NoY+R3YXKPhcK7CVi41sZga1pROxAset
T7axW7z35mvToza56Z/4wkUXAlaMjT3kks9ycPtN3wDo3xr04g38lJPwULpr
v5/eLjmAMDJbeYbStbpnPOMaUOv6IgCTMqVP3AIooEaIcCdUjPfft/tc/0tv
3Er0vRDQOKPMKO4Df91w8QgRIiGn7+/uK+DLbtnEvq1fdsAvxAcTgtutmFhe
JCR5F8KwAt2eamLv6k5bzuAt9cBbngEU8SzoDHqU4Z36WEm5U72HlcQBWBId
7WA7gvL7OF282B/PpVuKPsv2Uw+S+MEWpXPKaSmVxU5R0BF1eqHV0T1IjjC4
vu9xAAqRyao1Rt351Ozy9pSt1lFb9QuN5riJ4TErrr+tO9h6WFj5bTLvhZfk
Og/Gzki/Eh0KlGxeQTiBgb4C7hVqnQR5NfyIkphYZlaOVOLlaPFnzNE9iUmH
JcBcsuJfBRPWEB1sbEHYCZAiYm/k7uRYquv/YQwJL4dcN5KwfYERto2zGXhU
PksemH95UJhDgwgd96kyJhPuhLYGuZPX9JcpDOJVn5x2HTU8OQuR4SSeMcia
crvO3ph0vUQ0P1QaKoV4DclLAWzu4N7lFpvc5xxyo7ODp4V21jUx9BJXz/Ck
eIwEg5sx55uPXbEYK6BG43fgvvj8S8hgVdSQRue33MvGpYj1d//zY3ZWL0/m
3b86qzUsu7JVnGvd5lekGv/anOgW1srjegVGGAUAQDK2PvxylghhlOPCcU9L
tjBMwA+6JeF1xzgQhkGk8cCgkqBnhGqtS4kgpMEB0E1hGvBV2Z+vYXGYXPfo
HrG5kF8CUADb6H3++BXVb1jlGU8nUi0xoP4HK20gYrhZMz2Fn9xBz8ftfcl/
5AMmNbRYj5yQM3hLPOY4hFyEoFh111D62GAB9jNyIlZUk4sGPRqA/4JcHvMO
BoZlGD6MaDs6ZDmUlYDZrEZtqGBGI8Q6C6rJajkja+tq8W1fdoabVzyfLN6x
cZ88FuejkBGH5b3yxadQGlPRuoysvHAW06Xx4XGEYC/OvjBfQhHUBbymNhnl
jtphw7RPXi62QayR7klVGVogNBQgzLIa/W+vsUabD5Hngyg0itcCmgsX9j8/
1FLOuA3Yeoib8QEkyQCfFpdF2LQh8q/HaI3hdjZzYAiSnSbDu71YYMo51Jdf
li/ZyIiBkiz8aSANkN0hyDyFdHDOBfasmXSPlnX1yZ56tIDDt1MHZLYj+oa5
aXaUXpbGogiXRFMsab4hf89yA4ods9C6IvpLm2mFcaWyl1vmpZXmfRyznIch
eMJ2XAQmouULMWkDpYxVCERUkWRM09hToqdtEYF+0AcKyF+KQ9sSpNe3svAp
q8ENB5uo7DMbzYM6u17z+mNEaEfMtT5OeU+1m6o2fDj/j2gUzcP5AeY+LXcW
O5Nwz3eDEZo7fBaXHhG/IPdRqyMNtdHkYtgZKaT1fqThTyMymTZ3Z6ykT5oP
fa0S+xuCsOvxKsjrzPKa9BpZqRiWHmROQftRKglWmSMNsvibGfsev32Ih1sJ
h87YRD7hL2FAWFj501em6vkxERe+WWGDmTqbWklxYgnpxnkewhfUlk2lvTy/
qxkH2QjOvUQx5TI4bzwsS3E2BTBS8r/PwTEj+jOU6pP9ewt/wmLYmlnJ3rVh
gyPVVPC1yNhF48SXb2WHoYb32bynSc6mwJ5ymuLdpbITRZDzDk/s0ALSmzLC
LescOV3PhPfdkR/VVFQj43j1HiBp6LZmbyXdejp8elTDkbMfbbd6ZB2LXCVQ
5/ABVeYv1YUMYTj9X7wi36uo17hyfwytm2fzRE7A5JAIRkArNrvTuCMLrmrN
POW1hPyqyj/90vteI3+cUTymLhqCzQsS3S88AYHIiK1lrXzEy1K3wSroTkVV
GfivFio+Ouu9fI28ifr1xjShaTN/rwlSL0SvIN5p64qWv5kvLAUj6DhqumYJ
M0JvaNaZK9HZ+xOeM9mmQdFBKloEIBydJ5cu1sHbX9ZHNbxiQ5tPOn/p3sx8
tvN4AO4fj7G2TeYIjCk3w+dd3oR2kTMjwdHSgbyRpHPBPJ8UyFyQiecN1vbO
e7e0Crn+J3TGm1oaLg9l+A13/ty+Dm7/tHg3bZS+Jha23oy7r4k/CxU3RNH6
2sK0sIQAWy3tSo1cWSpObqHF5xwyi9FBI3ncnA4X+RqaR2N6lh27vs1ar90K
zpBFYLfpymPIbrQMCK66xzX6rCSvoH2twPSSZFPqDdrJ9FHsUOHovi1kXZEo
wFiCrrm+hodIMpNBKs+8/9r/aEw1OfgK1H31cHskV5whOtGXqkSPSAs4+M0W
JpZg02XPR6Sgafu1hk/M5SRyivLtYGRbWAvv9cpgTVHhiHNlm1QMMA8KCwJg
xO/Z/SlxophrheKqC8tYkImOauF3XThEfPPmAYF5voyCofiHLGEETdA7HIQG
pNgpodxcD4yFV5lP0tiKdPfGa7VsGzlTPGaLVzL2cFKUK0DWgprby7jHzMc+
WYJg6O1aV16wepwPvhXmrATGyLIH2S5KZEhY1+nUUqI/ILeEygn+hnxr1G6b
Sm+mLFjZtkuF7/cddDSbzNe/7mZAM87qqSGxrRRCTdskW6iCOLX5jDJzuH4s
LRCAG95Vz1POqDiwxRXh8SrtpTiPN+Jf64/wTgiT5nxBSv1rhopQrr0JJ3hf
sNa1lOdAKI/aJQhLfdeUy7riATQDYIdnxC0iQcPpZq0IkQXvMqOAO1/18mQj
ZqOdnMEiB8lTycqdgIuiq4HSOidwNMdn39JvShQJUe3PiQCLyThvHxfhmQvt
IuM2O2OygKA+aeQJjI8O24gCfBPtDzHv97l+X6p72Rc/CwPLpWiM5WbXQE8t
sMDeNG8XSPt1K9fASu+nSp1kV1Q+kycS0vHoT6yQlO2kjCi3WvQHKzpr8svN
38GZyJ5OYhGvuKzL8kG5UiAT0RP6lWB9Ydx3Vfy0e0eMY0KTKnOZgAZfA02M
haGAyN1uRd+dhObaqeOKlL4KX0TWizTt/Tvbp+hSusp5/SZZCphITfKiKOD+
AvRTjYdBaLbgv+fVGtVS9TeM3MmZTDQ/1wqCJYb7xnaGpNmkczljZ8oe2/wE
kmA7Wm/WzGJk6+gKa8lCN+NRcWobgC5oM/LpQih1Lh0FFfCVbbgugJ5gtstr
hICdZ70Y9jStSNuOsM/mh1G580pG3ztmIQ3K7VccE8d+3nyynygQyNooafiG
PQSImrLX+uB8tduMPnQ+7Soj8NBmTZYM2QDRz0WHJ4BPHDYV1NFYQLzkoO3I
cOXKbFKa79ykRRITJRp0pX3H1zTLyFFoHzzVH0aBXDfMuVnCc91OwdpShFl3
lDEgnx7wCWhQpEhHFs4duG+mm1AJ7jQ4DLgRRmn9RPIhwMR7eoTECm7oN1lY
3ecL88LkB+zr7Kht9pzwFG+lgg1b1tuW+6iqxjDIqtqF8ZAYfBL8KHtX89PP
UL2UdFBjcGwePa3NEB02wSgsG0MClCqJNkS9Vm0/cyuYEMwEr4BbURAbZtLV
y+0ppKZgmW0Ql+CttCwyrGuej8Q3gNDbTGV8BYBNhknQzok16eySUfcismHR
dUNnQbe52/QXMAezbpgtFeBrjGibQbAcsEwRan8m1Z7WPYKpwcydYMRKb2G4
t89PcVEP6MALgZ/D7tfBm16On5lA6gXAHI6LOszP3+hUoooBk5JyaAVhtNSU
lhXIZuoS03GdNXxyNAfOE2YPni6/ahgsBOBBJz3r+fZJqq+yrhpQlF16tFwC
rflzGWv0pw7aJ4wFBt77QvDtdParLI4ezKe1Gs2qINvziQJNCozwmotIQLJv
MkoVo38P6VTJ4QostiDnMXmbJ0dbztbEIq7anL58BplyIxRUr3CQCmRisW61
5ZMe5GokTir1qzIZ+VhCiy6jU9Jhu5YDs+5BmEUzK8+95rVoDydp8XNhFizp
9GcRSP3NnwrN3ZtJun1qQ+UTqjJiRAeQh0I25fVOS6UdteUno83WVLwW+d9F
XXQ262K+MsMDgOhqGSXACoDTbeSCCfmEUYvH6vlshVio07YaT4jxvJeNYf2k
oItrlh9NZLQIa3zcMVEF9k6RMri9W6rCexDzMbf5LbtZY/KUYUuYAfrVJVTX
vjSNN1vtYHsY02wxnngVUdSla4rUSyFYN5W+F0Y2vUyXiPcpMpvti69dGHLL
6qb5oaaR3kchbuSBOj8TjVcZ0KWH7jzvr+Yw6WerRqI+lN+Mnv62XJuPOh1m
VnCrx2blDau5LD9vG6BD1zS67vVID0qeeLAjsd6FaIRFCIlMPTfVImp1bOok
J68FrHdygACHMo+toXuMwElepoNzpCeykl+NDRhhQv/ZI6NpZLwFULnlmOsE
jU6jCJ5Z/rr3uWWbhcFd8k9ghIpsGgPlOfiMwSeGgoauGKvDAEIKnEwAbbwb
ov+ff5advfz0huVFURIWkkRB2tfW/x0zyByLJXDePu2/fkf4PA6byiVpQ02w
uOvS7gIXZ14T3tZwCO1PciLV3yz0Ljd0TutB8BSb+2dmKuTtjdO3NxLEL6pK
zdvsgdlmnVMKK2K9g0Sh36MDeKAtDXKcNiwqG4N05vPMzOvBYOaKJ3mAS21/
h+8HzwiRj8T8gUbtfhljgzqZSIwOpU2CIfuzxYHW3YmTKxobQ28wR2O9FZQL
BwBj11g/o+eKzOckQftMovaf+zkTOpUC/2xG2t1IeuWJv1EfdCt4jABeDudq
RfuvpGeEwOwMLFtWtAWagTbHUxsfXgH/sNMZIxoupyZU4aAg5kNvDZ4vR3ZU
HuoIEyIV4RhMSx8awCWHtvRpRkLJKVBJxiO3SDXFke+UmrDPMJc7smvbAOi7
VrELs7ZMwYM6VLdWnMwjzwuB4fzLNBbc1Tr2c/J6IwGWdCCmoHWCx+ad86pO
wJWX+9QMFG/5kAmEcM+Ph+BRTcjWVfgJOYZJ4T3imeCPr/lbZH7UOlDD0HMp
cbZHCg0u/U6FWu9Xh/1Phe6N9BapYiCG+XQeuEc90h2WsOWnxkg1599IDGkM
9mobPuiBT7YYXPSNqKU3lbmQr39J4x4UWB2PCZHLCtoKt/rvtM9xttMW3dDm
lE7WKJ5jWNwx0SzOS8XfqF/Wi6jhNrrVsKRZY8RLEtOo91xVL9cgu/79faTY
nqGQwsLxyVlLKcum+i7+whVotrhKEHaO/egFi9NQT/QFdtdzFVXOL13XRcfZ
Yvl60lfWa5hOqR6kQR4343dcCx7g8w0X4KGSVEsY2yajUK1VxCvFwYLT+2q9
m57gvFnA3iXGdz/RGwevirVn3xdHFmMxergy6tN+zpDBqUmalhqMrp7B3B4c
zsTVOmw2n/uomwEcc39qm3x1mqqm4rrCf0OMunKnVt47tt/haSm88n7bfVhY
HYh+PSe7dwSy3XRJHf9Ye8B5c8iPHeRpr5XbkMartJHOS+CbSvD//fTIGV6c
dE+4/KkTQ3kstOTXZXllzSKthglUhgCgaVK7sAJyewzv3cKNoDqbyem/d6Z6
XxZNJpT01BrlYAf3CXcCNv367jWlJwITmv+njvhIs8NH9eCGQPy4LMNRZ1V5
4K4GF1rFTk0M/m4/7DL2VA/gvnAfYght4POLcqmJwDQQKeTiauHIgZeHkQcD
eZumnI52GcMFklAwcgMFbH/o9sF4VINqX/3H0t2HHZZr0C8QILNfevqMtBAG
yBBZEv8ikkMR6Ck7Qxni0/nRq/oddEN4ymZyh7f8lxIexCsIMzRzAiRtLyz5
7KUcm871ZOyp6Rdp1UBL3wBfegSpSxJPw9/WeBOWUOtNjcKLddFaQqVTogNp
u4eqrvuCW/vv9Wh/7A4mjEarI36K1a9WkKRUnhXGq6RhRJAPefuoClfTydFZ
j8UAPZn2e7QT3gSel/Bx9K0NQbK1V0J7lYx58pqxrfMxlUoBJHivxjQP7oVb
WemHJmD0QusnSTWsJFIilaAuef/Bm+yjFARrMvJGMaEwqlGh5y3kghyD4ikB
OVsIOfBiTkOAegS0ZYmY/wXlSyZS91SPSGq2M2e3iO+dZwtHrd0gAAJalrJP
nRFCnJ0eQW68NtZzCDuQm+Dxlm+gJzgcl3xTJgP7GIaPl/3iuNyoTU5Wa/MA
6iO5EBCas52QMdBp4RFK6zDwaS9c48CVP/Tj4rS1Q2f/C1W075Os4lPfvlx6
BdP8Pvj4s/Bv7g6804p6aAZ3q0e/azGXMUr3keoKy/+GZ3HgZycda3wXM5hk
1Un2P/8MjdbUCL6v47ROw2j/95vNn2N4f7RtEpbjdPQLV0LwSL2Oo50mIhbj
hgeKut3+N2P6x0a4+R95eB3Jz7GfrNTIajG3RRT/nEB5Xudyxmq7rUjoG6dP
sCCIMujBKzUqeTAxgsqjWA7dZPXweVmrEHMEk365i5EbnzrbQNhCaEsTfSna
0PwGXubSSNhDjSKGxhpilrv6kOotL/FZ6Ns6HXWyrUm25Q7FPniu+3AWIdGa
bLIjnBdVL4EJqwRae1km06nk768O82vtHIFGHTCKecxfw6Pzayl0w5axj5Cq
efizeGkVDRBbKIJEtDdMI2AgQMfE11TFODMa0W1Ue/lG6lcXpv7hP9rOWzo3
LNkJTeNbzXbZcN7qjcKENM1FKb9uRJoM1DIY6ZdwvQ5l9UMdoUMeOxDDPUPM
UgHrMb0HaXUzYx1cpUiAzCRfNloYUOJQxbmXS14BAOON0XBNz4L/xQcWSGBJ
9kV+vOB0mb3hJSK9dMEoSLEFrj3oIjWEukE1056RfCCpnvrWbbOg7zB9lyH2
x1n8Scb5ZO3h4azIW2Zvvbz/Xighm649Reo+gpQEbyFiBG3PdqZSWzCVcZIA
bXEtmUfYawYGtWPj5rwLT3ZsmuJ6pg4+lVcln9Kkn0dmqV+gBbQraP4f+ach
US1EBJUIgnrxLYPILtMqjjL851lEUv+hayB2J8a/zwldS7EDFKZTtRntCtE3
A8M/mZs0iT5i1FcIHV1m/fROscLaw4YuG7xRMJ0yNkmdUyvpUVw27pYAplvQ
SrjdDuWtReyr1pUYvZAT0U1u4ur3QwHbJdrL3Y2muAIkrjqUGFpb1ckM1te5
6d/iYipmRL6rQsdwF3ZaOJn4Em/w8a4ZazJe7emsu4/7HUsksy/aNhbRRQO/
ucMwv7Q1W2EOTqU+Yosj0c4qgXKUvbWsVi4qDX4PCUF1GFS7r6ox1vqHXSjs
r8YJduxswaR2TsOQ2ppg6c66413HjPUX9/eMzrl2bOtDSnftT3L7n8zapvQb
MQKiCPbL/OktyGxl0qV2Q08xo8/bxUBD2WubUlhniX7tZupsJGe8db2YYiAu
gnI6VWlYk3npxsoXGAehE7fWeKkIWBOUZFSMaznlR9EOOM6psFkYevNUwyEY
tHZ+gx5a1iCU8CVuvnhdLY7aH7YW3/rIquRYfdk1twZQ/2qCI8pd5DEjXzhP
bYZX7fWdHVU0gyanQ/pcpJObGUapXTCpqksMTXv9biwV7yUtR13T/4KyPjTS
SAsIMs+RXd7bA3WmNztyl+FyYoxkFXAfOuTi7FJaW9hdsS2QctLnH/wUNDQI
rEgHm1Sd/xN068t7bwMG9y3tAe9/LbriufJmrQQ87jX832gjPohLmyrv9zQU
langom0ZYQWBeulvK1gVipef59j2ZOXq+urTpzCZ39sannHJIPUkdl35UYKT
S8dGV94//7tQHMPave4utKW55LJQU1NXuSXS64u+lEIY7sEGuQD6Oe5/27ll
Ez2TVcbs2eRFPpWxnyB4TRn0hdKUQHiYb8gDv6FX9ae0qNRNlUVhNuq9hnf2
t02VFbKmUSitCUcD+3jK2EjsL1QNZ0QdVg223Q0ysKnhaHT+ZxBj1NKK10u6
nA4FCC1YX6LUGH/UswSkV1Vp/pwEDbP4oGEpRW8DlO5ye8LTxpT3XSCTN2yK
mFilUkMYO29PB4PXyUQ2hnxJNT3ZFskxSsMx5clZ/XcO5gu09M00Gg9iB0aS
31IdDyzdcCVzcDEom4Oz/uG18YA2qZplBrgp1ZUfM8jdo9/K00dg3WqVd9kO
gagCP4TUv7kfwlxAa9Yk4jXL6vXVy4ao41HDqsLfCHUJGVCHuGqWH0Hsb0U4
7bkR84Qprb75QijfE+8h7G37SK9LjpXUONfB2WTsqEr4LaPb07g5Y6glwJwd
Fki/9ZfkX+nrCdVAHs0RoWiNejitiw/7E7aeYBYf0dNRz5MN4d32k5RSbkAw
PFxj11HNCngU2/9yc7W0eVfxKk3YM10vvAkpvX8uZRn0rV1LbgyDv9RIed4u
1IqxdZSOkdgA2EU2mxhBPGIN0uPy59NJUH4drWveht/nD51SrAauQXmvTwc3
gFhi5UpYJtEOaGCU420jQPfkHtw0BObfNvvJwyc5hQOee3t5jaCfwIvY+Sz/
IC8d+m93LxUqf/dnsz20GeX8KM/RMhTj66rdwjz4yAgvkDnZuFWlcTRZw5IQ
RJqhBVAVi5MqC2F5guAp/EzaNu8AH1buD9g+QK6WX7IzrdA7eCZ5vGhcQb82
cjoGVGtB8H6x5l02wGWZPZiLby9FYZm1q+Y4L3VztJKPYHuUCB+UKx0xNAlg
Wz20KfhC4tSbI5H6aR6UppJTahC88ih1fR+cxD1nTfhV+/TNrkvJNLr6bjTi
McwlUKIvv2ACxVvnkLwPO/MhShFNTkVl6lBvONVL0wbfr12+6UbZViNCN2dL
WS8seWMI/+2DRREZGOO51t1ueu4YEFcwIOrZC/F9LlLF9HRvYjc8BHAMr7EP
R6LDW/ljprzafe2M7stmwt0Jm6/2T6Cy4N/T6EpTL9D/D84d6P8VI7SbJDCc
8uyAlH+Ufr+mBO0n2C6zyi3Cjj8D9vva5p+Prosh0qv7en8/B6N0uNB8C7JR
Z1zJ7dQKE41f8rJnNUyfOlrLAc0fG/yZZyiB9ufvfeIPsU6egLhmu5bK/3WI
lew8w1e/rzXnBkbjTdJhmNRsKfQFoLhbtToVUiJrb3daBtxUUSz8iSAzvWuK
3npBKKYCciUmyfQtqZ7LaJWPJYnpoSSIClVkXyTKtF/6mwkaMenWqyrlfwZg
Ei6HjQkyoCbS/pzZPwNlnUWYjv5K04iGp7kR3kp2yhVTGFZoH4ZwZgQq1Bbn
869a0okEeOZ/22cyvjeoZeox0OXeMp3pcwuNdnLIuDG2fiIA2CRwfam4ZpZF
4ZFKPxj2M7GehhFE4TT2kB2FzcQ/6FKKdrgmSBcgMISuYPvv8zzXTDeB+36+
QDX+XFQu3ZHGGm5w03JEbSls2bMqmN+tmlXEwwxoS+eVTCX3mlA5pd9Gan8W
KKgljr8S47U4F6wLTYyvPbUFj8xG6a4lX9n2NjaGfODxsQLyXk4jK5pPceXw
9gLa/zrq2Q8a7cJ4sEhB9QxG2PWQZ+9laSVIuAok4iGfyYnDFgn8+gIARmb+
zrhrzbFKcUvDc17Cs9Mqo3OAkHhYc3Oy3yuKJAc9sWc0RvixQP+3JZ28ARqV
IXdV2qiVJEe2mietkHKgw7nNCdYwhd2RV97QcwqaeIWMwJJDh3xCJfpHaDCQ
BjQopiSh3vvZD+7dxBDsl7NRk9kHzJ2crQohXAi6C3hiLfCeGSO8MUAVYwO6
/FJA8zYE2/obE60DdjFjVgWOUN3biwhLbnypLf5HZIX/QthNnUWFWoAKnbAG
VpMNI1Es7rf2B3CjR8rZpM6cogFZA4e8XQ13M3GS3VXRQ/xnRMuSLQf6Ncnw
Soflj/vXd37wxPVB+bk8AYQpuZJbSykLFGNzuQGnraRUb1mz/CxhWG741Uqv
jfHzKgBqNieOzHMiJK4pw5sX6GiW9GWZO2yjcVRlPRHCA039MHbSUoi6lI2e
DfBLUu0J6CkdM964SvD0rOj8EWvs9hQrx52NGZXwBMdJR/m08Cpc37VteGzg
SlfcRXQgcPtM2Cb5ryYzyAtDlB7NwrYiEisipwqzFTXfOCNRsUEqf8jjHJWK
SRyWnTmXadZpBciifHSgjB6J5fJOWoe2Ug0KH1i/f+3YNK5c3SHhWB5eeidI
uRXRv20c9/wGU/iMPwhSkzfoukgcDcdsyfrc5lZqfinVYq9a4nlp4rUdB18V
Goel2Gi8NmhoY7+IY2vJ4Qfj/SOQaaX13eyOk9EmbN/cANpC7bGAj1J38wlS
YCNFLRrimI+ylclobws0aIbotCobsYTZvMCuDCygfRshhuiEw0xruEGfWbMK
qEJqgrVng+6wQCmHHUffQa6vxcBwlSWWuxDOa5N0wdYzS1Y05o6ElgSB82rC
Yer7BSiD1H4sEqPhQjc74jT+PNTmZMXxbEvBkyVLc/N2zy2FvLT4Yl2Y5C6D
x9fsDeiaUlNuwj9QzetdaS7y36XcqE3sIOnOcZhHAguXk6ql6SVDvKd/s16Y
2NYR3l7wDRzYU1bwv+ndqtDN/aDJkHGng5ur7VIJbdbt5qRM1H1KCHWHVOIa
DsoPxl6rLZWDk1ITp7kQ72DlP+zGCR32uWrjSwS9G04ME26NwLzPTAOJ7dgN
AzjlMJ3pnve3tlx7U0G3sJiLg0TnzbUbJ2W383UaJ5osd+Uc+1DzXGZNCMoT
BA49pZUTzETW8W/HQhNoQf2ybkFxBSu1tEh+56eam6v8zo5zDDrM3FMzFZAT
cmG0xPpDUgXoSK8E8esdHgYv6rW0OsjaIoz5eqmwadL8d1TF3JnGVqbma5oR
+6jbGRZt/b6rNATmGqgfgjXHST1iyG0lEa4kkaE/lkHC3FaVTuQVpokMfB3p
irbp/1e1mC8zx5t2QsZilAHYIX72QryUFyK1bVuZdpfLLP3+yWsAozSJ3P0v
p9c5HzhwtF0/jv6rafli7W2toSnZ1GVmnCLKduLa9i6/qj3sX6vWj0uZ8bVh
btTgmOr9HVxHBlEN+Yv7Djps33k2tUVcjMjmByOmDAVCl5DYLJ87vqFFhojN
GGbuk21+eCz1AamXQdqPgjhJgZCK3b8ZpWx+ydKTTgn3Yt3yTCXvMhUI2hTB
P2W4waryjzV+mJ9f8nDshXZ0RmC8k6viwT38NGmlPwmnCv2CcPDRvzHusEXQ
YSOzGOKzoecHbNJVf+O08qyvT55vlZQTp9bnt44OqC2juYzdYrxtN8LQ44HB
8PnbZNsffiObuEqQlpNKeTUiWvyNMjfLdQRaPU3z7GdmHWfyrGfnwvDV6P4F
2s4aImPc5+8qwDnfjWePlTvEH+nNL2CDRGAIKJRB4enH1kueePUqPR03PfLA
3+fxExp/iCTXCFq+TQ/GrdOBhXwgWicHnrSf7XYSnl0NaVhZqa3PGt+VaT/0
+VIYejBfeS8BCLrOv6XLwRPCgrpGVCC7If5k73HhKTt91xX9wrRmtKXUF3pR
uwWfPJJ8aJq+QZ/TpEbq0U4rG7/ppvDX+9lto3GuwoDDdS+73Gg99ywpQRH4
nQcK7xQTBW8x0j8qa8b2UHj3l4KxZqBJhLougfNq1+g5cIyVANxPjTLXLfte
JsiTKzIj7oYwS0i3x1D0muXUO3Pex4q0hoiPn3Pi71rDJ6BcLi9y2h2huO3F
5dZZ7dzXpxCb7/xiVs0lYy3gmsXdtTM+CTg7DFUq23hi6MJa8EMPp+0WiUT+
6N9SWK4LUUFFcmCFZUkS0G9pSoEK9CEc09A+YLATW5m6wbtfrALKShb1B8jZ
ot+qPRYNc4uyWHuUlyL3oeJw/MgVnDTZqxZZHmihAIBziB/4TVGhtZIbNYL3
lgvMTlVQCBggZJvbelyl4XnmSQLZ45b3BExuXgd/dAautt3DC/LxPzclsk3q
0k+S1pYgS/7BKmoUJAp9J9iDEY3/BtHe2N6YPxXgc2upARjKz4m18BERCDau
sBAYk6a6qTKTXVoWu7xjUFg9HcU4cCG5sr9MIDtjtm+LT08VvHrvL0E5B4Bg
4FyFBaCGUUShKBqN/HVaC5SD3xC8CC5NLZTbhbrm5KfnYzWG1/hGAmK7lqkJ
hK3YlFkA7G1oBuTITz34hy93GyF+tpUWXCz7JF+KFtnuV2EQ9Unhaa327WV9
ln9mPo6LG08aV60Qx1u5iP0T5P27nPFq+vUWOBoUkgGssZL+V+wBjU7yYZgT
9fVRgfxe+lKfMkT06CJwgOqSjnkh94vOkb+9hic++wGjjQDNWhaPnyzio1BH
yDJV14GGDi8quEnfYAyNoxZ3d8RshbmiggJEyxgwf/PcRkd0iaJVNpJNKu05
oiRh13mNr7NLF6px82lHatsOW+5gqGE0Qp7NCC5/2E+mOWJoQHv+wC4Rgn4Y
GkVS9GayjHKKdD3jUfr7qPJgZGZiMFfu4p5OJ/3AjBjLL+LEuQ7JTYk3WdaB
F3MWUmtymIssRtexpuM8tmkaredFwcO/gYXdiTeQ3ptJHbRIDGzyc7r8yUKR
u3TTjdy26Cgb7kTln53izUD/SMiP3mCWFa/oC4bYkgjlCkbYsfMDDLf6Lm4d
YzEf4QAxhC5Fg54+V42/ks/5Dpw3GKBgFxEoB6L0JfmL739//lDdqk/hjybh
cAKiAwlodhtZO+a2S1Rea1DuxVezwVfTwATy+zYsqu41PBNLhWIuP0ajv+k5
nFT6ydv6E94p7HR5FEvOhmO5nQ4JgDV8pPS7BbfG7reYcjVHDMwKmKLtHJ2/
vucyQbhK88yHPVvuiXgdTp3BNIKmoLqQ6GulpRHtPhs2QIf/n1fPh1hJ6SDL
aRZEXWrl9eZZ/TyeVqvg9b4WQazcT6P+LFmNiwAagdgW70Dn4nvfsrO2IFmr
akiC6ls5Bm9cJGAbMhuytoxSliHQAA88ETwr1Rs10o+RNrH9G5g6am4BsvyG
5WwbuUIxTQcvrzi0MnHGkseZu3L2Wilt2LDBGOIBN8FLLZOvBVVBNKw39UEb
xApNv/zbd3R8wGIM12a1uLd62h4NZFuLkE3C1kkBi7rv5Yd6b8armjOYgMRm
F4c2xMT8GIzugYv8gpfB2qMT/rhFnysiOdft6ESNpuZ9MAjg2aZs6qxq7aZ+
ZR5I9TCtmrEtiYjJ4fm0zoOsS9CwoQ3xQiBBRo2l9Mau2hHqH54AoOZowEkI
F6K+PrGamvU9SLBRoN4Iwizxxgu+vE//yoVI57E6L6qGXdtJuFh3VTcLZtf5
3pnViJZl6LknsiovA3twXtFtId4Xomsf4d1odkbeosc3ZR1DjVEH2U7gaC/w
p1UL+uhjYdpSFoyUY64Lzz7RAP7T+M1sA0F3n4eaZRgOnzDLUfOPkfnC7KAo
vo2ym+I897/i48pIDCYdHw/WaBijEARlvhSVuuvLWDtzvFiboBPoDQMRttHl
fYat67Cu5CDdhotssGFuHqsem1N81MPEQ2Y3HCANBoffNaksGbmiMZwpTVv/
29FTBmZ+ilWxcggpvxEX/CpoySqTVHl5ufJzfvRQjFAB+sF3ZAvGMSYaq0hf
bwKpvdniJaDoafmD4QylSUyBWf++YS+euedpqfs6Mibtq0wUkMSL4T4dM8fC
HOhz7bHFCob3ywQ8eMNesIoXOKq8pEUaqFV8DVkwA+kC82TqhVlBKZrMKHk8
nyuYOu5Uc8D6zv5bINAt6ZHspF0Ts2ibifxr/n4azk/jfj+VTmYwhkxj9tzI
h2QR8uFXUk7q99EJv51xBtW3N6t4NV48bWq6wGZAAycYay0SsJKz12e0ElFV
7ujoJ9qEQNqtxuowzn36QsR7xa8ccxC7QhpVth7tJhBjmkdN+sGL0j4b8eZW
KauLGurHQL594e+QfZ3mzxMPJGa+irtGCJgNhvXUu7xijIA08xDOdhNF9V+i
eiEBo4qZCUffh7oV+vY/z9+IJQGSDGoT/1wv/onsWtDhLndMEEra5V5Ns8Kz
4gkcittWRWnNxOSmEDGma0aaS16UbQNSZIot1zsLS//Z03YnnqJ2xhhCsYIS
URbQnoU0HHqlu+lI75wZM7+zoZzJADSQIrf2lW+AqRKFeNo5xpQP40S2RGne
hqFgQyS5oxdMXh5R761cshFEyUlmxmrjzebZpaFz2p+IpFT+vKDCuGOthewj
auvmRL90NWokfYqa+0y6pJfzdf292SJHlPzOoUIxt2LEKCuSG8dXomycxKzq
mr1CgN2MbxYAV6ZDiPy7oyFMaRXmjo7AyDWdxsWlhCtHgf749GLO4W8x66yr
0ZncnTjyZtVwUUE/siN33n2zbsMYDdQhV0+s8zgKOWo4MVPw/Vl7jgKDQAfE
Tg8wTsTVcX3q/RB1conEbhEIJ7ew/haNMlx30LsPhi0hicIW5SAo78E0E62D
7DFh5kXBi2Mx5dDu2+kYNRZSyh4iAt6THSB2TSWP2n2YqDnBq6eXj/Jlyatz
fjmi0uulePwxKfzZ629N3cycjOk4VGa13s0XnugpMyUiLpJ1yj9X+rZoqmgT
GGmo6bRz282PgiC2LCQGvqF0wgZQcNZ80waHcFq22RaMLSbPUSQuTHMiuSwW
1t8KXLknX35rWyRscmgNTM25N7Ul+fDBdwNxnj+Q+66oOhY8GAClkXSchnpa
qolVXImUruB7bc5RRUUbXNTRN8CfGCmCL5ghZNlxWX9cmS8O0psxBNFaGav2
wJdlobvVkO4vjYamxP+GNXEuTL61UF5v7RAKG7vKz4a76DVIMxLijtDMLgJk
uS9Re4QOG+pmSu+MN0rIbN9zWthBgD+JKZn6ExZ9P2l4AmtQ7WevMBLh6m+8
js5l2PDcZ2q6xtYfiWQV32zk6N+o+R5lt/CooeY6OZhB5ZmrbomSyCnXR7qp
2RQO+qiQETRl+V/bgL2YTBfGlH8o7XoQ4Jt70lgI2FeKtoFOinUwMvBG83DL
M/mbuYOVMIh6LQ82ZG0V4MUFNbg5uONn7kiTol+danx/MLzkV8Q4mAskNZDm
gFkmFAK0dbscav9vcSMXB/Rr6rtj52z81ApHwx/0TJmghnsvpqJvjKPdyun3
agOaAudHuuZ5fwWBtNNS2/aiV4C2JRkdErSIiIbe/5coxpP6T3qzC/mY1XHN
6USZsvLcQwCESQdEp7x0hI6X2mvyEZo1qnvsXHAiSmjTT863D03Z+WYnZF1U
TDUfagZiOrhCdX+MD2isrJFD3axXF49fm5LwtufXQYAI762/KxCn1PDSFu3x
FgueMu7RZLrOE7mjDYf0KhSNtqOT9h877TA7kpINwocW63gTknhsvR7VOjsN
pZ9YNAQ8dZby19tJgxxEvD4D10nVj3IcWE+M6CCfQhDcNjAexSE551rr8Orp
beZzsoqs4oGNP2aUpFf6+YWuReC5BzR184AFF8GZU5TT33gPGFSlnRl5Sxcz
iOWXVCBc3rBB/QUMgGbGYui1bttrOIH8r7Gg11Ztf3+7QpUSfUNam/YGjDfd
iDKxE339Kl916riSX4yMU07j9v9fkHOffM6yO7pDgRpJdZfAgj6TVJ0LvhJJ
MTPywl/9DulZ+PDEwvxAoBlNp5ZeO6VC2OCLQ+DPDd7MBwoFov1Y7dY1ghx4
dbnMW0/NFxNQiwobh+DNM6Mm/LdWaBhk7InLXLnOkHFHErqvhEgk8LVmAeIv
PQ9BQUcZjjt5ZnnfW2l1ibgQIcjyCAMi0Xqt2pX/1DWA1DysoqozhMRtjzJ3
2K9nVh5vnMaY6Wm0AE86i4KY3H1XtWvduWNePYSgh8ZmAKc61ym+t4Evqlti
f/PDaNezkxEKTUVwPtxkQRgVvryqwkEjy0/2QbEpVtQeULEsuefpOqzzhzKf
8JeCfH3kyoQDqOmMK/9HqPPeP5VdScfAeawDTfc5uL8R8dH7Og2m0/6fIp/2
BN2xCv1KINcuVx5Ht3avKRTKiEkro7VL62vpVjyo3+6XZl6d0xKo75ZXDjub
KD/HGCL5R27XL42J32b94hi25F+g23O/YfDODWcle66yhjoH0m7HU1xROyS7
DBcl1sEJEHN2YRStN5SzmtaaYATIpkiK0As1i7WirtMzY7OzmMlWLocrib4a
i13wrSBaWZQGBzzxMdkUNFm6QSUnTgj2oju7RSfe/0lORNqoRiPCOKG+hczh
9aHDekkEjcWhcAVfV/yYBAAYIZqgrLTdpbw00cr7visT7moR3j3KC0AzkIyH
X+dOVJftmrfBWMdP9ZQfPVhThAfrQ6lXMglP14Hdm26zuDr4D7npQOYj8Ykr
1fnmAGTt/LcSvG0BleZxpn1mVUG8htsk+QZ+/xdUSmbp2qSyEFP3OqKOmD7g
5LDrYka0dq1jF34zIn9gEnn+o3M7sb4V67sRi0drbIfyEKlUlj7DAmRW39mI
UixWho9MfavplXm53eac8IW3Np6mZlko+tJar8WFwn+AnGeWShrgLGrxeQu4
oYbp3nshSDzE3DpdGa19Bew9MpiMnhAqJrhPasEbGLaB4hR70kzzqaFfR4yZ
hFxeWB6AY8yDeVS8s5cM8e/Pc84AA6F79anvx9b+N+eLcE/yVi/K9e+sDveF
5Ku/L4b2NUONq5jMz3P5AklZfNsnzSQoRfs9j+Po96SjIsfYORP4fQZsHxsD
XpbUE1OXcfp8Tw6kJJV1Pafpap+bPY1gNZp6fZ5st/MCalA/TMpg0sjL3TFx
OCy2lQEqGeatYtQp3ipupXYKQrvA5XN6YZuLQ/pgRFOnwiplsudtro8hhFBS
Xv4RjK2zMgxY/n9xUe90vZ6RL8vwuEgFre2QuywqY6FxpNTmK/2kFjBXWzHB
epy0asWR3sqKs2Y6PVtJFw6H1IbM0MVXwdy90qfXI7f6x92cAnvd6twi4Nd8
YXY6rSHMH8AU1yNOayUONt3y8bZD3JEPgFLUcemoP7x9o6UpBOpWnoijX6Mw
DjXfNyUqE/d00E+3HxxPAJh/Ft18LYk5m4BN1ceck1dnkjZ9c8dRB25WTBF7
AXgkTQ99/BoGvP37xdZgj6PVXt9oLnv5tV7XGCampImSmolYQOpf5qxzRqjt
HfMsCvoMI/Uv0pwiRD6CZuV+ojfNh+NfMU9BasdySlmgeFna4OswjOeMXS/F
cfyzZhnaMglgeyewstPcH18g6cX0U+BS6GMm/A+Kez1eNzY2YkvSevfZkDmZ
HCPRA4QmGF8hdgvLRbe+IeTU06Qgmxv2hIMbnpFPoQBUZgz/SZlOfL70S5bQ
BXCcHKSC3Gz7DPsYq3fgl7lEHwpBy/5F5nsuP/SS0m+OCHLU/2A2eT7OsHBD
JUedkSFM9qyvRt+UTb5SJbTd77+VcSDgiXBrjGku6/yx8M6CMiwYxZI0IRhr
I1/AU0s0gzNNOZco3+ic6AtyxGN7oit+KZXU08+6kkUwahVx97mwWgZr8fUV
0pldPquRywJc89VkamNXVz6kPcc91blILW2VE1Z82hnXONBxQ4FvAolsbDNj
wlCWVuNPnrDkSjv+CDXE+D2/aQwdZtSws+Bg7XnbL+7s3wrY7AJklQrtAfW5
hOPG8iNgMUvqVR+I6hhC/IarenZrT7ZIOK2WVEq814ATlnCE46eHOdvzczc9
xbA5B0s+LXCl60fNWjwe0SX+V+jZjRuR8W+8VVhIkj2KmRHcxqiguf8HDeNS
BXA4aIYaLubdZiNHLhTpKcCWWViNMmFRuhxn/VNGGLYvsBLBCANFgBOjy+l1
g38gG1H88UbPcPIctrQ/CD8/TrVVt/QCxOuAMhnG6NM07yxD2c8QwlzIOT7a
p9XWD14ct4yY5K2BIH9qq0p6SE6YJC4R+YNl9rNnrLdE2u454wHH5zrnl2bS
KJvveGAkdncv0gLbKI8T5eL8rxT40OOi7xFxrWUNLztYzcq8MXK3WYLkb0rP
wF9+HOTfPiGdc+occJ1yFPqC5QpEqfQYSiSjHy5hJeKI60/lwrpF1/q4vpCG
DpQJ4Rsa1tJolje3cWdDJ6Xw0Adna7/cUI9E9wb3YxTgzSpRuzlzGLGRciGt
mDZW+pit99r2+sRwSy4juk8hFXxZPSshsvrQ1T8R0ljVtKf7RYh26UeaoI+8
66yWEsLe3HqNvZV4qS67BahHCfSLTIFf6Yxf3OhIMqxo3QlVCjBATcknkzQ4
GMfzCgFSU73brqRqxyDp3fjVN5SQJvausrr7k3awCq4jn31ZQlGOb/5AM7Yo
1qfhz/HjpQswjCMIgRxcsfW6UhXLrD0mSrRFgdV0HraThOU2bsB/+v0Kep/2
6npAmZWThug2m7087Ryw+5ZyPiJBoCiNqPZK60rbZHT6DZ3LMvN+kyAxuTD8
PwDUAguzvREb5WjUHFNIwCn6WvKcO6DZ699s11NIBLYRL7FK+G8ygF2SNRjP
AmDb+GXr0rmkEnNNye467UVKr4TfrOajoJjEPL73OiRQGdIzUxKN6OfQDzvA
jqvzC1i+uKEBKYGS5sM9EPABcZCvs6H5DRrRjiZGiq1hIgwSUyWngnQPp0KU
5QdfrLcawsNSsOEoh8rSY4gq64XGw3cdw5oTMVgGJjVnmJhPOxQDPK3drTxR
0J/ldAGDRPqI3rUkqG+DebNHLEn3x0tcfAqJ82w+NThonGcxr6h7QT432At2
xRedGgtHoQ96xTa4MfhZr3Syww1QIJYDBUiAB/ZquTFW6p1c2ouPIjQEXfUh
1+xdbM4teDHf6g0QktmjkUWvgYGjRKOnYj9Ctpk0U/21rYzcHc1OyxU5/4Ti
yM0XScwm1hQXJt2W3BsYGJ4HxlIz91PQ5ZsJbSk1kRJ8cjoKzqm6ZI7BmJ81
dEIZBbmJD81XqttA1XmElkSm0fuPypctSwZglEjXffTf7Gj2rn2iKqY6cHZQ
U1escxYCaIbetWLk//2XGalEufXhGN25lSSA+wnDgBFkx60Z36d050v+yGex
LpovILFwuf3mIjJJEFbVRVKkp0TS4/d0t7RJWIRFSTPSSfO8QJ6KpIFQvoHh
HG/aPJTUHZhzWg+I33qVJIPC6Vu66L2T1F1oeovq05DFP+zywd4tVLWJ7M8N
U73dFFYdArNn3xBmNKtgZMb7tDdB2eCXrmq+BTVpO91KWfWZaOtK7ZTa1jsM
HNwvbqtzcAx3uw0jM5ow0ndmzovX6kYt81ATW2P3vweK1kjxWbYt88W0BenS
uvbohkTrgMa9RV+pJ5sgPmdFKkylubD12cn2fUGyPJkImXH7zwe35+1ZdIB8
l4cn7ofPEa7HkUQJpsMsQQvrrhkAKKAe3z3r//ayEJdEkvtQOy+scfpVFDes
1cVYS2qg3R0JyAZFcM4Ygiwk+VCuPxRmqGNGWQuxliu2kDiJuN+StOvoMEtd
aq3/dca/iMJDpQFqnkNujQPblurtXdABvtOs8C/sRN39BjIPVgL2UPO8a9Gm
2gdjDVa/4TlEFwBIZiboM2oZku7xMlHxlpM1WRH+8LKh5z1At2P72TXTppk9
ZIyBKGF557FKIUTXrRyWbn2XZZ/keBLrGY2StNuiXRnJ95cfDe2AsL0gHUOH
BNf2xpnalXTxZdf+esZDx5MNtmMwJUIRN0ghqc7LVsHZNG+hP0pPdZjOC0kw
rjh+GmuYrYNVfOab9XPObKv66RRmcvkmIYQlr9YSbYu1IFpfyH8eEi6R0fx5
4akZFnCpdPZuHE5f5CucIrBZ3sNCWbJA/jrxeeQv7tClnAh8e/dSATwqu7Ut
5Dm2wi4vRNaiRQX7Qpc/hbyRGKpPQ+Cs5Tb7qC3ZCOoBLFlY8sWSHw9z6wiY
ZRFYir0OSe6+O+d9fMXzEdlv77zM/KiWXf1uy2qsRR+plC8cGW+Qcc3/coS3
AiSfCvN6AjUbK0t05nLKs0frV5W2rVi7aSU+r33rJljbLm5DDxxczNJ4PPzP
cbd8KqzXgispzF5fQ3zXMDoqFzxS2kb4f37FqoZDsRMEc2sH2Q+smPsqv5o+
NxPUZleuFlnwpjzvhXXqbUnbQDHh6H0ECfm/2b6fOS6TLuXDB0hZbxVtE3o/
tLDGIYlbMQTgBfP0iZ2xTloZtwRCrnXw07TV+1QzEJQ2U0GnGtOq1EJ0a9Aj
gt0rjjyiuhctZbJcJQVnrS8ezYJY5K20Z6qa+aZxg7lD29dkcXHCxF+0H4ew
R8YuCOS9F/YiMsdi6Yx7Ol4OCw0wCl+gQ4pr/i05wNviUz9aKEKC/lQL/mi/
wuwcjAlFr2YskPbXRLmHQgTsUzSU0LBDUxhSps26WESa/jb4oHOFOsllJM0h
PB/Nm5lj88DqR/9070xDLxO8W44DyYLgIBV7ZVrJ7lbrDkcnvnGwGLA4xueM
nkv7kfGoXx3Q966FmOh67iUno02s1LjKimCk98InhTDtoBX73wOhLcm2Ii5Y
buUjKyJXK1MVJrFxAAT3/HcWMxbPRswYnemhtZ/Oae+oGLRdFsC/FecCYCBx
are2F6TP/W6H6ZWt0goE8qdjQTqcNz/IXmfnkJrXwsorrSuBxOrb2jqYIkY6
eESkPw44rqxKFrlgOrlbBPwN73tLLBMSp2j2l1Pn0v42sH/yf4jI2FIYa0+i
QydxHa0p9a5ZvQQMe8nu9HzdkhlxDg69VDi90sdPs5ta8fMCF/kFT0qYfJOa
W+NmJaMbG3FJbCAheyZEKZdskVfvis8/gcAhVjqAwWdeXm735NsjSsaqwV2l
Q3PhdEc8po9fXMos/1F55L8a88BLdjOaHqzGSIfyhi6/2PEhdG99KHsuYJ7C
CXh049QJR10PRNdx4joPlXbpTdzoMPHCbHQ3DuxPc9OuzjluIcfnLiDfK5aj
tYHGel39F74zYYKVcCFLplCMwITUdXgYcxXrM6iq5GcL+HiwR0vRcsLb3RI9
txvtvauMeNTrAdZIx7UyoMyW+F+qeCnR4BXXf8T6vsRevv0GvqqIIE0ZW2eK
4+CFGpANvERHtfrOxS2PEU2o1WvXKOtmknVJDZSHWFNlgF56aB7Ai4NsfRJd
Ku6QFHtCYGDvL2+Y8+Y9kqZG/pMml2HIV8c7vLbY1Ctrco8DVNTWZo5p3PoR
1GqasM5xwSeOMsJ9xYw+1umVAr/lub32mOQJLKWFSZYrY3Z+dP9e1Xopnpd7
B29UHTOHlIaHNL/A2QkQcNK+XT/WDYa5HGY8/uK7pp/SEZON1PsoNt+WepkJ
v5BzOyLCEVFI+89UBZ1h7E/7JaLtVTyX+GfpYrSVLtiTGw+eCcpZj1sbTUzi
MNZZz3+uxfPaU6GO8IZTDDRolL2ucvI9yEivgvGQP/3J/iGlecBd2c/F8r+B
KA7ISrBcOOHiNoPYaejBRAFoWvoSdBW8GrurJyKk2SmgZB9zIxiE0mNmp+IM
LlI+QlxnNRLpvCUYZIodfXsJPOVfwIYmAeFNZ4wsyVowbtSgPNxVeYLaFBv7
aw/4sdcjuQDQ8Xq6LwG/QsRY1S2FuodDfV6Bh5xWpwriIthpqXVW4JYjd4Qu
MWW8DnFgUJ1R8KOFSvXurrQsssnPybg+TA9L44TJGC1BNhfo90JNo9oQ7ZQG
uCCllU0+BV6iHY7+yLva9oNNz17iei8dGdyCcooH9iPPt02+3nik2+9zkIhX
LGX6Ao+wBojjfRW8a51pa4O06WI8dCbAx+9pWiuivqEJRpqjP+1/kh4RcP2j
JhloxIf1VdY5QZJSy4ZRoZYwOGGKVIVKGGsEupBgf35YEjzZecjBwE0p2GWp
mDZp3jqA2olXIjlVQsnIdRd1KtdORjdOkEhYyXrEW3HQjSX968GiahBIoY5+
BJ72C4D+sVfRxojCNwZVMKgnHiUAtHrDlI6ZO7ffQtSIF0sAoClq9baMqGaa
EmbfMW3Njze637bOcAfcZm9iFlLWPYZEN5sk2nvSa3MtmTi9Kv4nyNWQbBEG
JijAKn/FvBUCOwFKJc9b8h8jQNhS575BOAl5IG6I2A55ZjAxYs6AOruXVgLR
6JoC/339bPSYZbs1yCHaJ8EB2j4WNwSr+ixoLZMZcdy5NTLyTNEXk1DaxYAx
RF2P6nUM4DoEsHrFOu/2rh4cbmFkWOpuELRlL4qh7VFt+f8Ux3+Y5d7DgkW8
s6ldysqIfoM6VWa4cbtiJNdOr3bOCxFUkUGw58HfiJGSuX6GXrFjNtZhNJn9
7A9d3S1lhBGViv8iHs5834j+c6IX3zy/o14jGIi7xDZqanI+62UmUNe+KNY4
JEV05qoQtIfislUSsr/JgLvXFFYtTiNOcMzlSR3zt6fgYpcW05Tok0vYgAVc
fdoy5mmkYfR1TOQTQiArWrqPr6EGOeV18jT18QL0kfnbgnDP+P1QZsjgEOkp
wxzj9BrtrdI1D1m7RzQFcGqw/8pmaPIjoaeZ6bjQZ5Y1oTQ7Jl33lT0jOYNC
+O6Gr7pGq4HndZNi8kO8v0z/vJOmEGhMCzCmZRV/oAiIgQIf36XZjITlg74r
tS/4hEzZjh2NcluX6SbQ7csSR06nYu+LN3zyWGPPNGPtLjBp3rn6nNySd8Ha
ai2Onogl8wbRU08CrBVEjgqyPysGlNp6NWjhSzCH/Jx9Gg9oOxuyyD4r1Obk
MOYLQ4GzbteUz3trjeDLPzuSV/bjSXdbE9D+wv9W27yB0FqjdVxst3ZjImoM
fPy5X3Lz2aqNrIKaz/ssWYgqZ4lCoGMcpgDGqHRQWDzOFJDVYgHlJFXfK9Of
6W0QZffHxdMQj8TRoc3Azzf9/6bW7eElGnkdhNLD5l8Xh244mIgOPCSgUrX2
pxUecXYgtNJjUG9mFvnDoBa+vrorEWo07QbCXMfkdKDzLx6mBV2DqfPIfuDQ
0v3Q4G/vQ6zBAFqYZo37zLzuQMzN3HsJutUQvTCBRraR1+/hlFPy98X9D2zu
QZCJwz83t61auq0XeL88qyRx8zudE2fslSitD9kPtBS3TDLbjb32YcU9ddxx
+cAzmWMqpsgFgKa7/V8Mta/d1P/GTSYbp74sw5fYHu8u9m7FBgz34jkteT0m
gYDsmKRkBkPWYFux9J2x6ALi/pKWqdVRVdwqiuYEymi7CbA3lvoU+drNzmPF
LCLBoP4U5bRECqEgKsjOwKOKTjExUaRHaRyp75idCugM1JRQgV+GDiMRknkV
/3n28NmeKuIfjItxPdUhjQTIOLecKDSHP3DHvBcXO++SYvVCEP0iAL4tUn5f
2Hr9771fvIMf2CbLL7rz8ICeOFqipSupZ7m6+vhNQYSiKq/9I43BgexpMYu9
AkzUmosu2v3sHA0KMw1fQLtOn1al9ml2ycstqgki7wmj3IiNWpbNu6aawMaG
FXhLAd4bovy1kFz2iZEpXatpSsARftszCuWeJ7jzeRAQjzzUT5MKY3TU0gpb
dpZrTphvR9FN/C3441xHypOhFEtkK9TmXY0V9l4VvyLDzjmsI1T2OzOlzIcE
7yhFxMrDbBc7K7kn4f8swDRmsoqQgTt07yOOycZR7yfF7WvCn+xL3zR88EDa
EBYHsPy7AtzDZWwnshnRBj+1cjkbQe0kU3M69j+meEdzJ8gqjWGZL/uxJp4Y
nQbufcS/7uCm0wMM4BS9DsaHXClDGwbtyWpfH/0W+cRx+ReWSJg3lVkPKj2P
F4ZgarBfJnYHkol1VGaFnEr8Qsr4ffx8gErTf17rrz48zSy+DZuW0GXyLeSq
OfflylzBXucPn9O5mw4x3lozzH9sraD0/dAPHab6+UztOC2Z/lrbCyoXe2VB
Cq73IMepA/eJo2inlk1Vn0Y401ObJaM7PMET0duQ8BAIwiz/lmwua6mUeVy6
H3nYdG+CwPHaDGHx+iOpboKlA7KbEysWu3cnm3NQXuw/p2DSxiCtSMF7bh30
nfdpmYuVAwnG5lqUqlOWXMjnrITje7qcU4MLvOSO4fDkwoDXejpPhwl79yKz
V6h9f+XZPb2kQj10e3yF0CqoURsMq7Ck/IBPlvP9aoaoVtSvoBi5BsxkVWps
v5Hv0+ow1yPZp7/r0x6X7hHfPXx7GyXbbwvjkzPC469+1IjpRAEQbApK/man
bH6vQqkoVVLvNzoofVnUcB/ihJ0EujHhDhIjMY5sU1B9BbJWGAiaXAfX+1Rr
w7/tLfMSVUArBOjZFQXgEoAOQwfgVF4CX6yioaZJibu42p8XuvUv3ctn0tqc
RoJDwCggbU5i4xKVW/FCM2l91jzFmPA+DxlmFCSsyunytuQrRygSOileczqU
AkJdKU2AR7syl6dMv46evTLrAmpo5WzokbdhvWnIJcI30qVojkWyTXmyR5DO
YxAj8k44TU+3QbuYFOYKiLN6QncgFSFMTORgP+tDOkU/yhm4R6tKu6FNqeFY
CGYGumseQlVxHlj6kb63G9L6OMrAI55yg6Rm9nUQ2V/ltRhdkA1IGkMdYIm3
AuP476N1aF4gdSHLRVRIZRt/MVddiU0eTCWwvZzckSiLjzNkChyfUXd+13NC
Z+4dkHDp9Ql5hvgGwGWZUrMXc2jwymS2YcihVLmGDTSiHruwJMA0hdgabZox
l3tjlErE5lu/prHYJrdJH9i3mpe5vc/ZqB2OWEWpuQNr5iikt//PwyUb5nt2
iupRnPtpX/EGOTVjwOnsz36JVs39x4Ve+YyU83DGo5/FJwU11JX8nrQxmPTi
sYO55vuAPjLLSA6h3OBcuyfMND8sKYr84DGwghX2fSYEpE0Z+8K0//4oJrxY
O+z60uwzq0R3p094MueVJFM70n5dAgaojAn9iJX9RXPbTl+AEXb/QIAI/ePI
d1itNvNQ568Un2ru8X6tabXfmDSCy63E97wrW/3fPMLculKGQHe3qjh8X/Hc
uk3H+4gEX9Z31fd0SLqpe263j6gkFQTYKmA/GJX2D9VtPKjoBc+6Wo7MPDsj
UKSN17nGZY6xAwBnKEGueSQQWOYKE8r9DKZq6AXDkm9Muj1nvFAyar6MlqLr
g8dGGLfRtfIKK4HZzXdn+EUOu4idAicxUbxRS2iXun66XlGFKUWnGlZI2NL7
iNNS6LO0KYctHbKAO64Pm8lcpGxxjB72e8uHRmQOqgyZb/rcAQ91iqm+PxHm
q63L5uzBbynlh3+9PoEX2AxRyFef4fRpjVHWEsJRbph+0oBXcNiz2IHcE+Ob
/tF2B9K/WcAIX+cA+XOhkf+BukND+aDpJOJWxvcHLNUJOG4rhQBobO9hvxaV
sdYGJZOyyHonhfp9EHSlxfVj92u3VktCwSOSJV+imbTX25PdFuqLOb94HLeu
SEOmBc4aE14xAaxTaXWU+Yj8GI0BfYnGhJAyNvGD86I36WAoAdWh9xWjgFlo
7tSc0tH9+CiyVFUJI3KvHsvU4ZybnLKD59sj7eO9WF2dOAy5w2L5LIS7+850
k0r7UD/jQW+lw0dI6mcWCzy2EYsCDjeKUnGgcxPRMJHLEr0g2nCxDxR8+9hi
GGKZ2X2jvNXq1DuMKsEaUQ7R8RotBKoS+g3j2k9nvxUfryiS8J9b4icxdHSY
DS0EIQtqX0rtlCzMX2NOexHlg3kEPih+r5plGdol3cmK2kw4A/OLEtUlQcB+
u2K7ghsTKlZxD3ZQ00r5HULACMZ0pyK0/9MRHhSh7xBoroztVcZHbwz58rrO
x5JbBi6SipC9gvcwoPRwqKgSyjsyr002zR6eI58k397B/qBcJAmn7HyOA/gi
n0mMMPlcRyQYfQMWAz7WKwdkPkPOh8JiA29GV4qauADYy73KJZSqSKYLdr3B
rt/eW0KDBzB4pbkGmvxLqmdE9sA/EmyI1DXykpAYriXbFeuJPYN/OEvx/zba
BkkdlJW+OQir8t1TfVDncADlfZBLdS8Wry+4NRJnULXCFmKXWuWVfra4wleP
zLVYNcHri2GBbKRHcpY5xuIWoHE4amlw80uhAtLojnZ34CcPuiXb8E5V/UIv
d/UkcKAedUsp1icjuFt6mG9cSadBFD/dF2AWsqYaGJZt41qN9uN9VdEOpCAN
yLHDZFx61UCS6EyN1uLuV0QZlykVovei2LXQypKwquBCf1/f7kb73h4Cio74
NxS17hJxe/gBUT2pabyWgqYKtCBDYpjiIPxzow/QyepsPIcWaZmdstTnRXi0
24iRGHSpwrXLQZ6C9VyT1i1YMyJ3bjKOlaZAKhuPnl7UUUqUK9Y5OMfnclG1
385xyar4bHLoIqVHByx9U6hj0FnPgYbY7D1z2fioFg55iERdN0sQs0pPACvA
kHtQEqqJ/NDJRZz0YZsG2fyYOdSUARRYTr6uVtDhJTvaomD1hDbsf+Cv9tDK
FAoW63Tppd20P/fKXIgG1492Y2F13Bu/CCXJhmyjJKtC7qsNSiomsUtDFKTX
iKL5cZPnYqdyHVrWQhyLCcdjNn4M04hTGm3qM/OqWCOrE0BB4CysJCX18xA1
Z175+ZsP04Jfl25GUMsN429Qu6YEnUtZ4Ykurxpr22gSkUqXkMij3SrY0m3k
3sYoo+Mi8wd7iLQvdXOnZYFEmKv4EPuGwX0dVTh+O1ZD35/EMo9JqaE0JY9j
DCE0DrYbVSFjbaTpbLyOofUZAakl5FFTLqJODM/4va5QtmLrBBsueIxf7ilq
hDF0LXi0bHAZ11XzGl4e23IS+BeGQ5DuF20gPyWC23/KrKLnhHUKlJYkmca3
U1k6fiV8MCABV2xmPQ+5zxzmr9XWxAYu3XdXzPDNi2U1fpkxsER5hfdgcP2F
0BQOhARBgbntMOgNVQvRwexJ04DZxhxOCJZtxVsOfUuN1zxPerjSAkARJ4FH
gwy+cT9MxaAIN8rALTRZeFr4gqDTYv0NnRm4RfAdK2JItOH2J1qVXh6ujosq
TZMgurgHJe1nda7NoHby6iT2wivrpuXwu1BbXFZRhj27fJz3PhcU52xwx/7v
brrEu9La1onvYvP0ro+kPNTitFBlcJ5aUL+rpMZ2gpGUwRkxLfSQ1Yjt+OhX
thWM3DDHK+4yRCcKut83SzSbcna0qPMSUqZ/ntkmf/bFn0Z4iY70GObmqCYd
V2PJfk9M6H1jrEyjHRaX0oMJIFAEg74QvGf7rcQ5xN/UJKwOctTcCCPN+KBJ
tAWdyJeCI3GfdFqwor3ALQ1GGxcitG/U/pm8JfwksYNiGeyZ6hRAKsbM4IGC
22gzWXkOZHscKpbUd19kshmfmNRqFo1G6biKSjy0vk+1LvAmCbQjskqdeoHn
aeYLxmIZFDDQUjfJYG9DQzeKW7+gKyF12r6qkN8PVfI5gbbdD/pK9Esq6S5v
nRQZd9oVk2JHuLnXvAiAQ+s4H/DdoJgeFS4L131d8vcbCujYzrLCoIv2eZ84
icSQe24xs55fuPHljDUvP++aFPVH9oIJhz4eN6OE0jQpaomUv6oZugTxbLqM
9rIvZ+GqINL/gxUec0kPIuhTLpK+KLn4lUfiQIVHC0dd/ZcLTn79Z0w49NX6
6UxM+Jq/Wsl/L46w/dLPvSOBjIMqCg6mOFmXB8qXE1OxIvOkoLBWUuokRDCU
mlvLhZPcfBv4QFqP9NePJcemuK3yjsQeoELu/4kIak/RSvgwyMQ3WsSdsyd5
bDefAYqXuZPYYgLIDL6ZDkpJYyazNSLAAxUPRJO45FsnOdQbECLlDW0jrMvO
vNk1tJngtdrfm5a8b6PHHiaW7FqIhALUKqZzMoCUeHKt8nSOl95dNdNzzi7I
HQTZ1LpwcCPsqJwdV+OwiyRAT36FWHm6I7Ee006NOq/J/djm9WNZv5+kskfo
CSlg54B88ce1bPR6b2EfvL4tkfNBf/IIahf9g6yngpfNRHbTkHPI3SRlKrVc
aq8CSbU1PAe5O3/2oiXvc0Ns2+DvVm/9nx/ow/uxnl7CzWjwg8kc9Heofkrx
8uQUq6MHkeD8J1/vY0XFZtO9NBY+6tsKeSXgr6TFdxL45WR+Z3DmlTIcNnHq
BDR+GWtDHeBE2b+nBFu5iyQ98aclQz5mcaOew8TiuIDK2Rp6uLhgusa1YZG+
0KCcQvs9n4IGusYZ/8ViT/Gi8xDRj3Zx9mLQeyzZF7FMJcry7oufk4oUv3iN
KXGGPf4P+EhmGt5w1aCKE6Cv809/KJzOSHw6LBAsrKp0JjCuJlHbSZnB6U7/
O+nKodpOj2xhS9HVKnOfEWmvT9D1jSDuGOw53ko4ndDmYnmw1LjWhnqxH5PZ
A4RfceWzKLrDrLHYfB37pIMBoqaeCpdi+0WmKrDeELiM6xIE8rQpry8Nb00m
VqD9Ms8HRgalQANLchHI0ZbJBfA5eq44DVpzZ/Li5OgvIjtGja14QYxCUhOR
INWGo86F+NOAGz5lB6Bm1Vq2/wF4hAT04U6yuh040Quegou+oI/GAMhnO5g4
lD+UaEjKUNX84jMKCihU93ZR775dYukiOjzCwP/M27ER/EazpeVG1Pdw2MrL
LBFN63wL+q3pOvvA4KkCZ1WRW3ifL5lGQUfqpHRMaYObOj7K20SnR6Gobvhr
VtfoJ3r17UOuSWTE+ZUe13fFcOc3M0VqHBB+5Op8tSfnB/jverTJfcFvkNxt
l/8ks9RHztppkr9/xw5+jGQPrdVLBcpXTZTLGMX2J1guqS1HtljxEG+rkzfA
0DlDyZDo4ZrMgV/S6sT0xNFWFTpVIusPFu/39bwxlZSq78uHbUfwAaSIqUVH
qYAIMeTKYGXb4nqSZVI5xPfN6Uy+xag6ZsBVhC/JDfBZOpp305tF+RsJxjhY
zmZOK/kM995euP1SPpi7mtaiOhDi3DrgEzqOuJ1Xu86F6PoTIIXYMs9peqU4
rplEH8H2jfj5aiR3E/q99zotM7TBsaFXpUm7DB2CVIRbzP6l8rqeqlXv33VI
n4wHHwt0zNgqbSSq7HopqAg5I0ryuPjFJDL71xBMyHJ8929QJkgJBQU3p+e2
b8aCWvPrJsuLZD54gVGViI2n/YHj/DBC9swMQeuJ3bSwpNPmip+HH//pRcfO
dFpm/9VrDaZqgXyB+7T1wO0zqvoFF5lKzjhEvgXCghgIGFw9/w6u2RwezAmh
v4b4pqf7Y1njq78Fgn16u9FBPkabLjoYOyeRjW6Yg/IBtrr8PQJz6HOWyIhi
SdAcQnHMrL/b/VuBwg8foYTae9YhdBdvhiVQm078+9Od1uOdpdAICUIxZrvK
0tHBuC+7MdVRiR1Dw1O8MpYLc1sNmIN0E3cgHS3BJbcIwL+2nVv9EOCY6MpF
6QpP5nmNLjvo1lo0B54PS98h6LblEwOlDesr9/hDNfFRSW3mxCyxJmemUwKN
i/30oBgFya1/Uh5HkkFR4YcDZL13AfhDTqaEMf5IiDzY2Y/DxNS1bVn4ZM7T
k+CeGSMautlkJZTheUQxrZZD+CJ1P+8IzLl8HChREZvf0hv030RuwRydY7mo
uPGz1p9VFAHlLgXAn6xi0wcVLcZbcU2AKqkLoUlIp0J/Fq0IsTbROHnsQ+AI
dYYcPtztcc346PSpsMV5WLt8CNJ+Rk4ZFNO4KAUpjZY5yLMMTD/aj32MAsfs
S1xY5lArmS4HsASg59HhHQg3qAHsd4SIJqSKo4RIIAxKAGzJRWlL/U82xdvw
Rzp2x9gBoyLQhUoR5NbUu8151iwkuE3T1eyZipO6bPQnlHDv5hOtv3m5HcpD
7oiNb+HpeSX2gSKb0gNvRjSwKi+m8ow2Mdk7yw4zOZ5xcBDcLXNIIwRkaUXi
RYbzkU1D7sXrz5xUHEcZ5mZbrGisoXvJ+hqjmJmfJu/N0dkj4m958ovjry4O
6klJ1GEbixFqNtzTPqwnGPex33KvbNXJoDqIsf6Zw8E3PGpy13736gQVDxkH
E0ioP1ipIUQCXOEIhlgOLDMKk+RMYe/OXyO7nj0FizQiHXqYVDpHPggJlajc
NXolag5429WuECMttp1IJxSzw1pJycGtajG9xPxkkTYe2hQmSmTKVfbQ06Yu
9f7rcdgGOfVj5qDdycUfITNBGNOUTkTgz3AReLHsNllFPCK1sJErQAinIlxh
MSAlKhsIuRn2x4DqjtfqB0gtK1c9UMLy2dI6tESTaWc5SClPka0se95MSafY
70z88JkPQSQsreCCaAlpu5lPLxWe+F0jzuUciee2WTmwbqs35E7GHBle9dMO
4nIpE1peey5wFvgNyqUAauWi1dxS80U703wuQ6rW5cPKI6IX0/ORhi1Po5QZ
+VV9DliyswMwLuR0t9y7INJavQ785Htf0DFFl/uCOCyHY8y/SAQx6pUpo+IC
1NqyfVcAff9YsK1wr6wc0jdnInZ4HoyHW4VcZMdh20xXQ/+q2fzVX4P96tcs
qGiZaLVXBAE4RDJYb317Ukp0VfEOP7jcOPsLFU4LRUS3RZL6tqB8IeJ4Y8IB
nc+GmlIgLftSiR9Pj3GL2tUBX0GoaeJacWHMZ358L7pOs34knAYSxZdql5iu
JFrjzrKyGtwhWunAkDTVZIiisf3j2IVrj+JkH1lK5sO2XraADvmwvFxp9gnP
fKwdJ6A1/jmq8AjF0F6YsTwF8H/N1Kukx3343LhLAUnsfHZABwA1TOiUPA+b
WLN5mcy96DN0DZLDSlgRbLZvSJAE/xyf2MTm3FvqVj0sBaLiQTr/g6VK7gb1
Ok/WdhjnSFKMzkPX56YnKK5h05YDCGuZAqPYkyo4Oz55Bwo3Upfe2bLffr/s
M8tivBwxgpiiDodUHotTbnM10gaKNT7a+syZXpUCJTtWYnWfy8UwDSylfubZ
QID5+w3RetSl2tA6rrTBh9kRaBj/7nKqVTf3DEHqbQMFcdi15ghDOqJp5qD8
xNbDo30mfGSKXrF4c94faxvZWa5Fd0ruQFBqwK7uvYhp+rVhQ1ae/KTO3o+g
m3WGoZURaktPMYWsaEGZKNW/9p/DX6toWsO5Fzo8vCah7HnEysFZfxldIj6P
1IgqwT84Kh3d8+0e987G8DIOVZk2I7Utf/E7ZJ7/Yiwfp8A4ohW1z9Umq8uj
zXqvT56+pmODq/1dM6m9XTfZKteUWEJJpHHAvxd7I/uK6R6TKa+QnryynP0D
eJful3EZrph7lWUmsuo//w14PQRhEX4grF77WYBeV+cXK5BhvuQtFDiQZTTh
YjJ5BZhCW5m/Aqz22xd5MVR4pNhBadaqLZwIJsCIrHL4570J9X6aaL0DdtxV
ytM8n0z91u+NL2/ZpiUKXNVlh2qrsMtJfrSZoIZGq5QTCGHwoLSy3qGZE9n9
qDq6UJdTC33YNXxMr2gz6RDRkhgHTIpnQ3iqyDsG8SHukLOzuDlgTECqMJvV
fW9hkub1dsugrLGtBWuLAZUcaoAHOFv0L5ornmOuwTfkbqGiH2vrRTZwGaEG
+zjw6KMqAuWQt9cH2wOGBe+73d4SKXGdLmBekdIei7kIBSZLJO3/fer3MTWj
A6sfI/rJFEOP0HLLk5y+8TqPjzwh2ykPSz2wAN09jj9T4Qz3/kpBsVKhT5bZ
unR8D7tEHo4WY4OUpTXKQ+pELn+wZCfdW0Ump+CFPRwGZtY9ccKyGbxEltOT
xvDR/WhQDd3An5nC/6Hcuj8hjWnvgETJL9wuAZoYPrQpA0gBjrtCJ0HFZgwO
skE6gEPhQ9ebuDZhg4+mC9XYoXMrUTG8eFVSl+kEmjfMHh4fmxuz4C7hTUBU
qsaQKk6OgJlrwHqYvrJkCu1uP3YcBzkPyhDzN3UEC3hl70ceowQKTvEWyOQZ
9eQxZY7yt4ij726WZYiQilYWMGimAgBg6mZsO2s+QqIJpW/qnShRZTm4nlXx
GrYUVZ7hC8RjZQGY6ah7citoCB66Itslcin4SmPguX371Fb+xzyIQLYZmJye
ktcpTr8z070M1hSdfWdIO+RQ0lEkEMzJtBDlRj2l/u6VhfgSQAzTNQenIldg
44xq123lzCDvSDVPI14HKhUMYWwWwS2o7m41cN0DMmGQ+JFU2rISTe4jOb7W
JKMJaWCCxumK+K8z7U5cPIgJuJWQqsX6b3Yr3Eoxx7ESWnRz1KxRmbKewEbZ
XPU/F6HNCE7hSH3iwxu6mRNYO02p2yLPOFn/i5ePjEuYGcRMibWU+awBJ7Du
RY6TV9fFvZ95IYkc/gKv1LHxDKhi+BAtC3B+lyZZP5btsdR8yjCD8Tm0BqzY
10r7d16JkHJhgdgPvTOO9KKFGGl4pK+l2/fGgrtyrcMOEtlnKQSpWYpVHw9k
JwfQ2A7Wp0fhFXp9NFAmvo2TSD526im0mMvemkS7jc5Gfc+Q4//lqWlds3/B
gsMqI1DpHQXME1C6POkd8rkiXN953rQe5P8EGBKOO0/5PzQIECd3Z5Ggssim
SFLsk3Jt4SDVCxjzJJh1W85nKQ/KRZc/ccui+0c1tm8Oakg8UbMMMYhikKEb
AwELk8q+EGbHK8lwwULHOKrZChLUGLSiS55sgcmEjizwOLQW0vNZ8kZT1NSC
jqHEDszrWAnLvlWcciUU9rMcl1lbRVZ81jL60dunNcqu/776O2Wwh78Yv7lu
8HJaLOdeOXc7NJx+QOibPTW+MQc7aXKQVvdjuwxEvbbYfqrJpVNTaYRdueTO
iuQPtGSh1KQKsV7k5nIu/MVnHKGHt2vQ+xARbDl42nMqsS3IpzKo8S2oVjOp
qsdyM6DPpeKQJGLjxagUzYol1jNQb44R7PRkFvU9u7+Xd3D+rjgN7pkAuCZL
hQoW7B8V5bkGXAUWOltVLZM6kN+QUbyheLQ+9qtxCjPPKlXltMeJ/Ln6EstW
20HOKMQtA49yV9dUg4t/MiyC+2pnfflFGfSPgkaQyArm1c3NSo50KssUCHBo
NRuedHtJLcovrotPXPFSNqe5R8ZzfgFwuEGx1U46EcsxI2afcpvHeBkbhQMn
bQjYV5Qi2EWHpHeSPgBYsX7n9n5L7xdKkhsMG8Z5qmLKVAYQLAvGB2vfau/V
7RH3+W4xnwSOt9dnlYlD8abKijru0x2arOKFblo0uP8GqBl88PrRj6gy3Gbi
33/qjQy+uAvAjl55R8Krn7Q5S8+GGcRd/9P8QfSTIHdThyWLYandOnlNs5PO
tzqaHVvPrjQ/77QmNyI8+ZLF4dp4hU/7JkCHZX560sJ1JlD3bdm6Odxmji2i
XW7h1i01GhUigCzsFuNJTM6CwRELLlTWZGS1lIlKgafhMHafV187vdTOWGqa
d2zjj1SrConDTLdUnD90nLLXwC9JKJ6+8D8ITP+2X+VIFMhKpSb3EcYFNtWN
UtNbqggOsHOjpqK+OQ/S6axTxbpRt6icDU7v1A51758IRK2c7HANfqPJfLN1
HepUduUCoPqbNBg54YmgMYg7d5OlDaRoM19n7NzPrxnWA8c0mn4DFCM6Pf7K
9EN1lS0cJ6GqMCUYf866nEJxOVaDi1DQFJ0T0LBkltvgMStrqiOrSAEQ6KWn
FPocTFoJkw4zuao3nwC1ay8cO4ia5KGxaMfGE5f01ttQamitZSHQTSV7DO5D
yZn4TY7B3e8OeKsUQZie6brc5hqNfqM4qV/idOJXLBxzpJl7MOrAbcm2077i
VvvldBYGjA89CjlD7/BuJDgHpuD48Pd1EQbpMMAIUYl53xPn1rJUcuUxu5oo
2I0KrM44z9nhApJ/jLsgpv722YT/nRUj/TWdq/MVQiyEep1z9+DLrPBAYSXz
PAMy8La8XUVejxOVRN2cnMGItVDBBmoKUl7FVDBO11eBZBWlK8DGgXBZSFj0
uy9bMe/THN8CK+zlHbTv8a+j5yyQsNMpmuujcPj6+ZM1axXsVCJy0SqtGqzk
CfbDYXnXafE8E/ycuJI44/iex5oLBfUluvGc/+X6w8IjB/ZBc5Zs94MqY1od
KJ+HFcvV2r87mxzeQmcuops1YYZ1Ke2TeF0eadThl2GRy5vEfrJlbGeUbW1x
XsefAG/FtQl1gBeyHPkGJ44Z/Jd7O3pscnny/dFVPW+p5ldx4Y8eWE9MkWwO
8MET//Kd22AhUKQymZsSm5vS2qVvTY0unxGD2C/2ZOgiKfy75h1yYPKtWblE
E6SMDqtIn+JEzd8FJr0VXlfd04bNiswTmCqFzGNi06C4HbQLwHmtQqAMsLwS
ZM/TFC5rHHUX6EhIUvaoWsMz4J/7hmYAJ+W0jB98K/zMBYMMrfrLJs7/nO7K
PWkfKM60NqzepEbZSgstMKO+u+/HhHADXInnOHjekN7ZuiMgSW4fKxCM3Q58
wTdAkZ9pQbqEWT5pPRHlW6nTPNN8siRRI6v2gisOAyfgQUFqAAiwOAqNwXD1
8UTmRF67IlT/Rd0AfmBZjEndxtR4KqcptRu181F7x1Qw5vc/7rohzAsB/Ytc
ZzYkeKfLl4ZOqHYSTenE1LPNy/YPKhcB01t1dUaXzr6ZY5gpRXqjclF6kfvx
HSW3BcfhmB0k11LzZSExA56pTMutKHlO0OyxRVB84BgXxSzVl5KRfDKt15T5
KeKDg8LfqLcr1DPOk+T3rcn4sN/Bhy4knoYRz5jKZolJJoNHkK/4ZPboJq/0
LdkWHDgoVTjkzvCxD6bDFnUHBkNE/CMqecYPao9YIipGXDsX6NVyn14+v9hc
BcQqRW8ueqCjgfiapbEmoUE3caNkqGIg0jo6yHF72P1Y+IjMyndW2m31xPJi
dUh8u6//joudsMooyu4Std0h8XDyJCIODDnKgjJ4mBV1PcpthoU5tca72QDF
rzO7cEBRp6R815Z1FNmsIyl1iXVY2iI7jjsjwnEOqEzEEDdcKhfv9AHaCWka
0BtYtujb6ZTwgloQcEj2IOd1x5rAIIC8vDIfggegUNFWcOlZ/j5lyqYCJP4M
UXhVanZdZfoUdgo/NVaWon05RIiUUv16MrhQ2RBhCqb6nImFNZ7GEBa9XB+p
We9uf+kuKMQu9wkk8I5/ZxBmS/TEL9DbIoI0qkwVYkPk9Nb7aIP0GwArSWlE
c/2Bm3w0t/DkA5g8jxXvUtjQQlgwuHiB/ajbr7Grd1QDZFcDX6sfK05SkTEf
hKEanVAOlhazxik7kUauQRjB/eDu8QIO00L8r1VE6QwlTYin+566Lsv9A57v
q5GcTv1+eax1ZF7FvVfJm1WnQSKp/8ZwMNrl03103/Zf5NsBg/DjKAm/YnOV
7+zY9HBz8IxKkJpDroCYEcdP0H0Q/FgcP1g2vfcdQGTRysHA7nYhtHqe4o9w
fuML8HFzrq4ou2u8RMLtFwJ8MV03ro9Rf8hpr6UnTVNr1GYBnOMk6AsmGjLW
pOS6KnoClQA6qb2veqvVDIXxNlmP/rrHEvfBNDPl1dWEkdfjPGFHDp28F4Nn
WW3Ha3HbymrOyHlFDdJil0maDI8/s7HrTo9JGDDbAmKcw7KqnTxM6yOpWBfj
yAfe1CSiTmAwWT8V684+0cqsULkJzPMVNHetQO/+QXnZqZMrcXJk4NqpY/LN
4luKvMKXQLZL/lIe10/x0nmkk+FjfStiO8SaLr/YhyTAPCEsf1/uGv18ACGJ
qr11V8JY9TZHiePpGTNPSNAuM97BRxcyj4SQ0cRahpj1dq2BmcbTuQZVcuNW
71aghQjQ/g/aRJyRoGXQ127RP5m8d2PncezNIooUksvaz8z3hSaYKh1uyPCX
hUEDsow8K3flyKHyJsp+WIeXcm6XWIArFoKqrgjTO0wRvjvWpcG7KIOcyxZi
SmGSaxf/mQCmWd3tzuUzPFfbzT7ltHTY7EONL9ymSR5XB5xy91D4YYiaZ8D9
lqv9KWQPE0mCqKU1vZvi5Cv14fkt7pETGDxhiEbU2YHu1Xg4GFNOY2Q6i3Hv
ubodqHbWGOhumDM8+RlkWPcU71Co7qoD/fBSpXwUQeUyY3pEFwtzGmSXRHpP
/4U9NO0DU1pZ95EoqaalnCnCBt02m36qenW45D+9/79Wl5x3FwcnC9wCy9oY
sNJB8ZpKLEvpnXA8d3DoMMpwADNdpnZq0j+YE7lEuiSismVOyhdYjK9o1nGd
zMHEeODF0fdWr7wAm3Pn+E+1a2K8kSeUdd2ZlgYAHWwpXUEtZV2hN1/2BksJ
/ftdKQR8dLQzvS+YPXKIa9R5UO2Hnx3hNLvU4ZsomeiYv2OT12M8I7S82v0j
oEgbojOjJTVg1hI9cN36felgquZWCntctWFQgyGSiA/0mtTu4Jsns1qFBXFd
7ErxNRe0ND/1x6PAX5jYk5n8f+FoFTFkCqXzDAtbUbp8C6FEGgOSeg2BTR56
aMrlQqhPgbGzjR9DvjX9kzbr1eYDDUMoxmTvrZd8DktxcE5RJuR83pq0Fzhk
BLunzuf6RHIw+aYMo1c7v+tneVoU151STXk5EP2U70NWZqDcwnoow/dlLOAj
h/eII34cndKpLl62AePSow3id6jR28ZYzA8tAXly+hnccP4MtZeQ+gq5VM3M
1zXy/2GFASY74F2hpPCHc6lWj3t89WGJzwT9MJ0GOE81CCqmkhq9+65i5uZL
MT/0Kd1I0SetdTdbPSkrd4m3Pd+VHFLvaeucqhkyyrHkmdkLQdTvQXWVIsML
gES/+eArOl2ZaxTUS/S0FI1E8g1pWwl2+hh4VJcQOMHL/RKKQURmZmTaZ6Gs
UcEi1abqkudIhfAyY8TUK9thgQDpEJSDgQXDjfgTCUpi1ZYCmYEtUfqrIJEC
Hflv0Ysl4IF09V+5AlBQ2vRwEfEBmgDIMW3jYIjz/h9OEIuZ/VBfzt97Q3PX
H0cnR2ym31KedWe4jMvJ4R8PtDsKxuaguNxPimiBL2Mot49dnfIruAcWIVLd
QXepLFKbVVON/gRA/6InonewoCzuLLj2zDt+HtpYcXi77Pfn1xHAltDYewam
/INdrKGwuygF+OUxg1FuaD66K5EPEEUEA1/H8uQqTMEMotk+hIslD1QLzKty
kOfzt+E6oXrUAoCdFC2s93vjDJZzLWZjOmzg6/JfzCLMB50Ien4cDZEqVdlz
+Hmu1/hKGMcaoYkrwJKClFYkFVOrqoN0aHPSaDUiSU3+8jSRjbx+1Msm4M9r
ua1iJVzXJ4+cskg0I+xRD0T6PETDpj0Y7i7oHNlIZzTn9A+1SV5DizZtp7qG
uhsuCvo0+kqNz0S4OejjVHtRCwTQwVTZuV3hQRpGX9RRu2eAR4OWXE+5BnH4
l5qgyTHec5futiyAWoWadtrri8TLD3HBEaLarXB5LJnAf9FVTW2m/1P72mKh
hWH3Bws92svmHNHU8gi07x81oVsH+lb+akERTipVw2ZcwDhNxrLbdRAZ7Dp8
TR4xJjttE+/GjpVp/Luu3A6ZW335eaDDguXy3PQycSqpMIJqgrwVNxo30K2z
ADcvfFgsIFoaFODsZebekEUTKi1mndKVx+O44oHxco+L0If/wWJsVztS26z+
x57g0umjnvMwMSpYHN2BxgLvEz4CEI0+V10VxkGlRTLqR7FgmvXpQfev+peT
tc2Qc1s3XqzzM0dWSvd99cdb9J0kxvkdGAuXBJ33BhuKcHvbNO1wMdCYUcsW
SGwqPvKvdyJerF1CuUS1maSBeMmOPDXITgsA0CoXXPmtSUwE9ZSn3RqsN/NM
H/vXoEFJ2XFzovNFDQ5qYpABe4fqaksqU6kv8VP0oqFPR6HIuWVwV2Baci5Q
i4njsBliSN2sjnJtAUsKxQwCFvuZfpDYhF+HsEWbllGAXdq46ZKOnKPJabdQ
Pmf8fDWKPDKa3cJ2fVVwhzyVhqMk0LjJh66MC0SkKxYo6pjpbylTRETfy/ho
kva2N5eENjM6jYpy4ebsq3JXy4XSOvv+eAxguY1kD1JJYSSiG/gSq3DKIkvo
SyI6vYxLlzcIYGZWD1TrmV62e99LV+EW1kw9AJFgizrSKkyESM08oFlA80kZ
TflEP4FflIksIVwWkEgjIRbDlqv2FhOBEJu/Ktxeix28lAah1+ybCK7rifp5
YrjqdzXECnMeKGgpr4lIc5EHdAaP4cstVWnzKFFBro1hMvzgEQYda0eOB8DB
IMaI9fiGRFC4TlJ76P3oSEcR+rwgASAS/VVw+o4OcVOUa3T8xKz8kQ7Ln8H5
Ol7WXPZBUYAYw8bNxV2VUTGY/EjUPywMzTAZ6q93bRJ3lg4BSGBz5ubsYA+F
0h1+2ihJcMSwWkSeQ/CTFXIlYY/moglcDDfI71Bka9pN4OPgI6h31O3tQ/fa
nB+9ENK/hqAsNKBER50o7KcM06fEzjDx+t5BcDXybiNYRIpvN7ztcezoEKmA
XHlc8nXzGqcneXGAiydMLu4+w827fzGl6gboxNV12ICNiGpMwwpiA+nz24Yj
5kG/CHWA7DpVCHXm7F115FH6eN3UYApD0Lhoq9CVuttnJbpKHqHxjB9eQGzm
38rwzi62myaOJww2p2UQ6Vx6C6pRrx2Iv/WrHbgHUD4aZT9QmuER2wBDvgI/
eNhZ2fAClJ44kllV7envx0FV5AmF3pCqUfBEvJSlQFPmLS09e3UOczooynTa
YAkvW9GZKEdJFLojr4wKMvjaFuKU75IVAU+TgYqlq/GfT5WojTqdfPKlvvV4
0WsKkCTqLULv/smzsj30eqXZ01umdTXVpRQP/4ExJJhQ+CI3LRPN286PqY1r
PCBetNUiHacvcLvbR+Qbxd07Sh0dCtpst4ZgaWjkcgEPuIf59SVJW0SVHXJE
WvPDa7VuP//4aHvUb7NTAtON19mgan4zyafmZSeJJEBWpBxT5BEJ0LpblYo8
pJbUX5KsJGyIej8W57er2xuXw5ptnvXz5EIgtKfSCIxLnWHuHRhP0CQ9QwUq
MrsVkA2Qco2APAPUClTolzWPLs0biy+qEbEp1296yzpM1B5vKFdbqWG4vE1K
f9h2MutYBB6tn9xsklLgdeNbcXCZ4ItdNybcgoZ8HS2flj9OpfdxcWh/Ztw6
QeLWiLY6NTiZw8fxxk3wXmH6R1uglpzIsELr3xmDYxumujMlAhc4CYX2Ojw7
xdAVcMbEiVXRJT/6qVZGQvmALRkp701hKQM+3plCf0AbZCVb9rYIQHz4lkqJ
dmBlefJWi5gJGBgQMl/w7XxkwzR1KLINTKv1Q00PtSY9luKlbYjbAvFJs1rI
Wo64etQZoERdb+Xyr1fn7maozG8vWpoOk7rpvtqrMhwEPQkteFpRIvL3anvl
p8CXYZbYaMfmDGzzUugo/SpBKcRqh3qGJ7CK7HJIAyspu892c6d73CcgpaSo
kljBX5tX7jXDhJyrNF7UFl2ANO0WthhyRorlJmN0lNsmRSy7D7MVp/OSFjcR
ZIMRHIB4NJVl9jsrlOlc9NazH7iXWKiwanR6sZ5v18qpkMwgwu02ehU5aVNd
Bq8/pLduBf8b/p2vC+GurBynvkpzkmGN0WMNeaOg1jfUWuC4Cmfswj56PVr9
3FDxMicDzUV1DX1AzHXc6LgcafDW7+OtiSj0m4oR3eeBSS41zBG894Y2oQpF
suA+7vMJlBit/XxIRfpK5YfWDNqCG/fFLu5a3fItKisvNfReujSgNbOhJ1+S
qrG1zYhyNzvDGvmBr0V2BV9T5af2oUWMZzjGkM2tKUoAJqowZwVNFG+Dyqzy
jDftSOkvkp1qEAPpj/mtK/JpQYncfIGSrGUS9sf2/FBrJsO7/tYRPRQ/2V0T
t9aU7k/MJE5oLW84Hp0mYyDdRHq3LrzNaCw5zb4pxaR7SGNbPsVpcm/tqNSA
8+DCCwlUTwl/6iZ1KNeongFGw4+we0G6adJP6hCDCngRUmd4sgQ5WE8TPh0a
9HykI/zthg8Zq6PaY9HQZhRVgP+uYviVThT86GXiYBsOmKV5KFctvSbYvbQr
J1C40bsPaGV3niQfe7Xp+1fkRNQAuoDZ3hU1Gg/hBIn9W0S9gqfjuzfQBJUY
r7AzVN1fpYo/yjnqAQNGQUOcVJfBw2yL6qo9WyY2VXu0b1AloCSaxWY96Psg
N63DnwlBf9UND8kUOLpqUKTLtqRKeVkve60H4Xsx9PC24WU2nbDn6KhTnCkc
HYvisuJiwDoSDamSl1ImBW9Avk8xNbpnPN64N6IbC/EdaI/ErKvI4e6ieKfu
Fa6MNTy0cU52vTHBHuSDZ75eNfe7W2T/S++QTkfEothAkJSuMMIyTr2ZcAFl
NpZc2oefKJ58lRN6tM+DA/WkHcHLxSD8UrMwg6g/fPuLRU9A4IMMNMnHwYF7
6iH8O/AvUFhZd7Y4eGyxLUq3pDoJGO8YgjMqqvt0YZ4jVVXXdHY2E0rN0Bn8
CmgGrLi/GzFCduwie2vczROyiuDcOPdbNsCvT8XKW5hZiwsavoXQS0K8C9TC
ASL0u4mAA/31tqQXRsxJcov/bOmIS4XjEz8FSHaS/9jTxxkgO9aBJWIc2TQf
HPI3UtFUj0/mQcDf3hQfSaTxIsrwRvRGsdlo/DTrfNk3p32Eab6htKEF+lrC
tZHUI5MxKUnx7+UIwlJyFDBBY7CeEKCW8ygAc16J2RKv3Cpa8dzUq1scneFJ
ZqURdQgNCU/uj/M9TwR2tFkN0YH6KgYE92v+PCSpwFl/+K/UjAqLADeYvXSy
FAmGJQJvzOWx/HClVAGo5becJNoUhGXhFF+zt3S646+HfZLV5Oc7EeiSbjJu
21F9GhClw32plEfSAzhk2iCZ6FCPkGJygWm4InjZGsW5HpjOV6lddjJSYUMP
ZQoFm2WmvcuDuiVa4Fpb9Dzy3D2pnArLrsF17X5RCvu7//unHK/GRmTdPZEM
Il23UE4WwIIEyLd9hlMwahg1QsAhzs2B7YkqeFaIW1pjLN608Xw5qwdSGPZw
TKO2tgTPjwFBIxJ6BpeQ4dvSNrmRNPptffeGn5KH3aCXlLEUopegGfkn3k5i
59pd4tTKPn7/nKT8pOjuVE76WPzCYNK1l3ysGoFlvRa3nZ8aVVDng23d9xcx
+M8rq+hm3emlgybaU6Vzn+06XHfqpn+42Nu/XXGa5ji9uuyDXFkha+RJBKJU
WWWx1UA49Q2rCBOlc5PD8zxIPN2CFLkSpX8Bqtg9LXpokEr1LYf9w0/V8Puy
r1dOMlpHGRKWL+zBgB/vZdzKEcFtWXPcC7twjghzAeCvPWHt3k9N3itbGtvT
ePur8QFcY4rY67easfcovUaLYJIhd28kFNXY5osd37pSIprFJGv0HJSB/2jr
ziDuy4yjfRRZXcttjBbFitLJjPQ3OSJyeSkAIHImrUFasdb57ENTBbgY0RDw
derKlQ64iPUF2o3LCCBboZnoUBk6iE0T+7F74lKgZ4XwJwJFQxVx1YmsjOHT
Gsb62Ydw+oEopCUFKkGcewlJeRqzN2xfzOwOXQx7eJSCpvK2iWDGwDxeNcVt
ai4g2XAkGJtY1kC2m8WzNRGw6ae0rb/2TG3SfNacgrcW5aGDtPYCNFIveHRB
1k4yqM10T0BheIYJ+d1672NoVpEJg5cBV6y6uZiwpjtI0GXtiyAEjWvEBKQH
IaLQ8PNemVF4T3+v82r3O3k43eCHNk4WvjnwBW+bZ7durxukNwd5dJD4FgNK
prdQ1Uh6Jh/a9y2jcrcm6o4FR8OBlqBe0qMWOOmabVhn8c6zWqpTQxccMCNh
HLpaDht42thsgZdSEDIItYO2a2+/FYYjkRXs2e7Yw8sqfxKVDncR8LBYWEZ8
1955Qxb4GcatofVgGe6kHkqe2REE9YqsnXz35Vv+6M9Dxd5AUOPZJstNRB9/
BxxOSX7qeHpSf/y3FSv092upm7e3sI3ieQuEIaGykoT+euN8ZquJ6VcqFfng
YuYVFE9baAzTis4G/isbJjWBo215Y/Iu+MIi5brMOWCUP36Z/tAX1vZhYAqz
GD2UZPVANPqWxHBC2ZkofAq3H4sDu8ar5ZMLAreuq/vOs+vk5yp37r6d2D6l
J8WW6sl20dvk6g6QNRwNZGkakXfT+mdniwfnbYtOm9Ypp9lFFZH6Q7zxXXLM
7zZIJZMoH2wcuPYnfMXbksZMwmtfuRVOmwENhskvpik1/obp4TtgIQqn/o2d
dSrE8D3b29yWirmRbIoPBz8bg+Ne2eBCrgz/D5PbcIpNebfsi0yUIs/7b/ok
orNDUmfkWNjpqR8asFhcM3Lv+Hbfelz4EeJxUk4atHu+AcRmnT4pqri4MUMn
Cvgor9NXkZradBYfa5EcnDp1ljI9txHnKYPeuKVV9W2i0MEZuZdi8MaNOMdq
WGHb0zEHpj+5fBvXe9xG7ZxSuC2TK+j4ElyDGwQuFGfff1nlFOM1hMI8m442
LTeBSqW4dX11Sa8hTlS0iG5gicpVJHWmXdlKZCS1Th+b3badjTYj3yGL4K28
NUUj4xcLrSEuxUxQ63OwmkkR1t8L6Y2VxDjcMFwmGV6mTBB0eThlrvyAEVO2
roj8aMv5fFXDsh1RxENHRo9ToYl/ESgUB4rxyjGOUGkNEXlPODe3fvqn2Jcu
Gtezqp7naX74cPTEmHuPmTN27nPgZPdnE737mn1fkM7woVteP53EYeu8e6Yi
ZDfvpE8bl9CHbNQEK8srENwUzk87MWU0ypjoG/NxSCXq/tXjbMZgxzCapP6u
T+crui8S0XOGDMZ8lw+emx0JpW8TQA/XG5UxT+WopozANV/CkP12W/gltBsL
EfQvBLwWnWDHcD+Dw4/U9vvH97bTXGPBV6vlW8MOthNyqzvJiCLekYhOf6RY
NzzCg5KAJcnMQNphM1PzRNjZm+cv7tItEq6l+xvJmqCVALbDQ8oeNJVTRq77
1Ht0KOkToDKdi1elEvM2v0ei4Z+DRJHtmJDTjxe2X5tMrVNGWK5vJnG1jrUL
DsKrLK3tok+/dhYOsmFDugZlCFT3BvEwuCuoyE1NFgqwQzHl816UPyEkMc3Z
2+scVQSpegm/OMlf0vrFIDOMT2pF5H2potLjTgvvqCO5LA0CcqpTTke9mMGm
LWJU7zQ0ddHM+p5YBOLGh461IdgMERu0xK07XeQgHza4GRiuTUyvjmziC9Ch
+D23irh4M6xj6YUVGzlaAhtCRkCyx+rht4RjluLMys/CbVc4htP7Y+NPMsb2
L4Uy+euMeSf64iXtHlIw5ulwrvKcSwENGbuboNWSU3w5VaqN31XaAUq2aezT
aPp7EXSPNv04mTTSaUhtzdEc0ozlRM1zHL1ve6ceuxtuurWkS/BwR8/TlCzu
PXzjVPJL0GpljkXs6TUAoZcweddrZ/fKQWa00uXdPIS6I4rofXy3mYUAMko/
jWhehklin1XnucTD9kkHx7AufINqesoG4YCrdKz7eGHNwfhFYwmTDvPGe8ww
0o2oRWjRAdetJ6oVosIMJFhMnbg+PkHxKo/oTPnodUV/NycpLQoV51A2RiJz
ItEwRb+kEW0A0vs4RZOAK7ur6h+enj11rXt0UMKq/iw8gIHhejGN5qzWcsPr
zjCYA5qtBPBLRQNDsjzwvitfxQT+X5kQ2zw7ePlCBrpOyvghNg1COFE58chv
Fg+MxKsJyNtpGMElkWeeQnNV/+yIvgJDfhd2ujywfaZS5Dff8k1mERc4u3Br
1oyJdjXhl2i3D+oAgdiaBH74jPQECEyuYyACWS1D5pTL/xUau7RDq903VTIU
HGoXE/yv2z3UBHr+FmL/BoqDIDfapqEFw6uGpVnwifduY9pHwdMA1fc1OJFD
L+1s3J7oP4va+ix4r3T31CrMKcE+gLkPPMZFXym1ktDc90o0+BmmM2bykypS
azjMwuHczLqwG1zvahOKQzSFhozGGJU6L//ntipL7xs8RVHWxK3D6FFFZDNV
yUcLawL9b6Madq6yBvYKkP+BZBVh74FyziAnxM2PlPpmGItv43Hyi8L041u2
H+LzfBKgrZ8IIxHa4HuWa8md0FTCWzjRFHR8Er/o19yfuEQMX0MfQiV5q901
yKBob5/MalAi1d/eJfwRdfBCI8JGYV4qVC7GhkQ892LE3XodANNLll0n+fN/
BtHJSF9kwhWQWW4JvYdJTYNftHMAreTt5ZOO67LfJVaZ8q4I0B8FhE/N7ioB
sOR06qSs7lEyHPtnM8Voi+obluRTiEaCa7GUo1FUJ4t6hwle9ht7f7CjcBL1
ShomRGHEQqcXZSW/oHT/wzXSRBOUY1pu7rsYQosyWrhL0ypL/BKZh/M+akhf
EQg2/pmph/PQcNwoX/yHxJKyFuJSFjYxfDKHiKmuacokO6vFnug7tdNTLQRO
DTvZ3nKFTW01BI2GOOvbt9HqgmRx1hRENvV9QAoMXgUueC6dKwu2XnFVOjif
/1WEi5ZpYSb2pm9ChU2or8k/1PzDpIXN/LpVfqbbLAlGOcOa0rJXR7ObE2ZP
KizwuVEsWE0jCq1NybR9H4YSkZDhLGXjHzfdEo49KClTC1F8PGfWSzUV0rta
/w1j4rsdsnUu2TVTMv31OJFjSUFw4/vSL4JjAvcEaW/rnDWuXvAtMhZ+Ie1m
M/9ZC4f+JUvBSVehxGPcEXcZIFy4qSJ8sZb0xeWx5kn+nitqoldk+L92Xse3
QHgWP5GRy3wTkd+YofiiJ1gObBEvNqykGHomselPrbcNWYfVWQHNX6l0twKA
mMJPzir9kPoDHK0Rf6S+IR+aDZRKcTaNGagi363fpiC6O6x0a5xLAOUgd3WA
CoFWJGQ8s32qhcylt2SffpjODQ5Rg2yEE8GP4lQlLCgvqTFs7IHnfhKCQqbt
bdgJ4XShRns/qe/bpQJty9hJDIS3E9SWUxkLFlYc6vpMfDuqJmfxCqjrZ1UA
JszP5dA6qzFbB4HgxbOvqv5u+Kw7MZAnGKUZZEjLwdG6RMuA9GDmxVQyHunp
8HZq3wBTL9yVcpGMWW4pXrtgtmFT4OqzYYx5FqkWtKmQugN7qGvbPLpxtqlF
oJWBc4jwPJVI/kXxQGy8rn8qRr59cIUIRZhk5pe9wXKTVMqAkLvnPtr54NaI
MvQnpVt8/hhbHgn8mgLX+83RsYP40EaVs0TGxZt4DAB/4JFdZHpb65slFCGT
7O/FuNoiyeySnK3u7J0gR5qgTJOMsHRhgTd0rsp+S65dPq9E0RPXKOGMhiVk
3taCJZ9/yu6Y64fLyPKUEKJG+eFLjRVNYwbxhS+oe6yG0vhUa3rdrOmgJMsL
FXDw1XId5Z10i+mSQMxZ4krXNS145leEtFtJjsqy7rBezYSUd7o43GK+ot+r
n6JtdUXfwBPHBLUqgBBxnog4wma+ThH73Y0+GFFXv7sw6qMGpRxr25vIe1sv
Hm/Ml9l7C/hg4AjYTw3cdKnRXnxQ/7k21/uU8VYDU8sKOOOSQcd7kT7b0dwV
tLoSBpNUirsICsz99hUZqrbgmux2SPwGiANyqq2CjPupNkRwET1nVdBvL84/
zH89gR8zbLwX/9Us0h8Nf4zOJxsZhSzx2NFYHx2znu2fCPdfW5Hs3//OkGnH
PPGrEEt25drKlvGZ53Jpkfyw36wXGOP2ibKqC0A2l3aoGQ/Z+Lbp4AHgLpJb
N3s3F9nuSim6hpSeBAQyIq3kJtFWAGwQiMe+H4s62LRLtQ+ViCwgFPG7LCYr
Tt1IyUIRuF0xA1O4LrWxn3mTs/nfr3vxJ/PdOg8Ej373cMo4vvQGcL0+/LOk
9FPgOENMyL1dDsODycOqosJ0WovNUa1mfyEDEg9XXRwKmzwlGjs/U7AY0ip6
MziscwpyFJeKJcYvfbOg4H1IbKFdBaKs6h4cs1iqMaDplt3e/8Xcu7WBK4zU
lPyezxjBgNnlTT8XydIB3aVJyaJH9LCKmBgNTkcCs7g99GOGy7Ls4bZUVv98
otmgVJ33eet4kB9BSytdnvJUzJifRtk607qpPP0AEAVsyd+F2BHdRtFQwJkN
91Rr8FpNZsDIdyQ1we1prTOGDyY/WKmZhENfQVVCNoD/ZpUdRjbq7joqKnSy
/sxZtE38LY/K0h3oMp1Z8xnJ3RpaLB5XWSmso99O1n6Stqyry2W2G06slfFX
2hi0RiP8acuBE9Z/wa7C8S7qKmZeeBPlYCvslssKgXlljCXcupQW+XYpxcBv
X0f6xgUZuHdT4ylUL0FzX4qOnlHK2b+RF7SgGpXUPDck+smSQw99RAG4I94k
Tb2WK4qYlutjPOmmVqw8XWYX2xwtfTYmvt5Wwb2qqKzyCTBZJ3sPJEB4g6f7
ajB634ciH59rBn77/rKfc6VnN8ClhNWTOvT/lnxfIoAXh5Ecu19LBqV7Esjs
lITtBOXiUqTleVukiuUWioTPmfeNJx0IIXzvGIU/gJYTAl+rbYCW+51F0YZ0
n9NYyCNubLKCc0AhqxMBkzHCkvRzi913f7BRc7+G72n6s6JjHu3CvO5h2SH0
Sr+vBXRcXUFJO52LH0bjJS5E0jAeFCrJCnJd3m21gWgSpvVfD5mVECY/RZnE
u1ScBAT+zfuLGdxs8+srKVUcefrY6BVMblNF4guKTNVy4VckASYsRaIRiyao
yz3xLP7iXPj4CMG/ujObjSIjA/q5x6/aV4eWRH/j9eZIyZuDUDAbbHbcSE1d
gL9TsfiIj61pf8o5hzSKS457iXJG2piOYAXW1+2k+2SmUFubSBvryc4i63WM
lifmk6zHl+1LJZKGguofInoMRM5CWPKS6jZXCro4MZPc/bgXDRDXH4+IIQ6q
VsCaZqQnCmiM5CRqxuLiVuluMDqAHKCQ8GXo42V8CQbzvBJI+v22+zUBFyF1
q+uHXEMNm5zeFal/F+ULwA4XBrJqjbw71j791W0/BAkFBr0WYfVjtiqqxsDa
Vw0dgFwrlyLSS9ghJJQ6laOQLjG9u8OlFNkLkD4XmS+IL4IX/ehV65RITgnE
T9iEOv17V2JHSotoivWwMBdlORvR74wvVp5pHWWnkcPMZVG9kjXQeMxnXSEL
imn84c7jqj9TxAu94gVlRP9oFm2pA7tTZImyBI52vBEyrken6Y+IbHaO2q0W
PtrjjcJl6NGo+3H3L9qCX86qsc+ydD5Ts2Fz0Juae9wd3FutzxldGTnOFGJ7
wDSk+RtTYby8+TpFY5Sr5XZCcCC5RSbYFsfRniBi+xRgQc3aFeZ4+8uYIdYB
7SvRhx/tc+xbBoFkn0GI8iBRuewgAc4k2q9ic06+/ExR0QUn89dSigKNOqcI
vwy88lXk9HhZfR/HHVi55V7MLSYyw4Hx+HjQcjUayWL1jCE2XWuzvewSffE8
ctPioIQuiMMXj/j+lvki5/WOUwceWvSYvHI1CJtAes8VhdRr1Z9e6S7idB7m
fVRnX7GXuzlbeGT9p0N86AlNgj9EXJXXGgkA9kweCk9ArZRWoAmE6FW5s57n
ddzSJnlfGYnyGNPNA9Mk43s4TZZuhP5agz4AzNiIi9Sw7UFZfYBY7JmmErt9
1wkhAoPC8Ks9pWNc2E+N08IqFSorzZ4q/t7PbO1JOi2aCi80oJ0aF6SuJlex
SjE+PR7ccXznnaFaVB97P7luejsAOCDpvmPskxm1l1/w6lupFyYm+GNFPByl
MI8fr3Jn05NdCWIcDdwgOgCf72INFfZY8M/DGjcgzFnvYLpgMCiAMB5ogK2c
f35XpUl+fpl3nIkxztkKl3kgCBtm7sr7s85Qpiz3qCBaYLIsqJwwIuTY8Y1W
lM0JuFI/TciFZ7UBsPzqvgmGh13WBahX33cgwIRN0VJwqiQJYoFD6W6uhmOk
wpiWm8IGx9Ru77FlG2MsT07BwVOvobIuKWPRcYUM1RX+8IE7JEWUbrRajdQB
6iDCNVduFs9adx5MldXazw0imyMayOt88thinWA3ccfLPMNhMPqUMcObAMEo
9YpC21IcvbsQa6WTbHe+dT62QTU4S2jpujzacfjtP4epHnqYLQe87h+vWzvB
4LcpT9oDGEQioBRg6ZToGxu3LYAnPlFRxz/P+0ce2vijt18PwtT7pX9sCs4H
SyV4e3y1+gvr0yugaLUqB0pui0bxZrasLynRDvbV6fAb2ZTc+L6+lYLPqeaA
nw3LNvPptcIQ6DONjF8wRu6WQMaqDziCC1JkMDodYjf5qi11u6Ymu4X+2LmR
FXcfEjcq2gsF4nPksQJQ9HS78W9WHlle1xfHvLhxsU/fCAhJezpMKMdMjDJg
zC96MNwir326oV8SReIJEvc9uy0o9ihFB1Zao503Qt9TgHoISTa9yrlJ8KhN
3gQSVnzWMfU4zSs9CHJ0wOwmLnZiqyBp2atjpYxNL4EOJksakwuPCs+/bJsi
e8S+vHsnbbTgm1IFMo34onCYHoc2+50K94mMbewgAto5xE2kHYwUf+kDYqrO
herzv1ZaYg74pn5v5EhWh5xBym7/8RqMAPZot6akP7VbAfXdt/ocD/AKp2J2
zlsTZUFH4g69hHexMjusExHNENqCWP5THp9zwxl8TjePJJR4MWx+nWY8W/K9
0+WPudSGruCwuJMOdZadEr8f6bLAH428uw0LlRMFsIY/j+xrTi0L/EErbr1h
pT/ghd7zvh08SSe7c0ciMYyjpeTklJZK6iHiMcSJbNDzJPsseyojG1LZth7J
YMXM2i+7jJlGo9m+/etY0d9UJOMeH4Z3Xxw35t5wqTMwSTET7r5CEzNu2QMe
AbanUtWXRfJFZj2xK0oVMCkEZqtW0egWdsVkUP6mY3Oe27M92+/AazSG1mmF
zIwSzUK6D4/zsVkIYY5B90YQ3dlfveIa5LktMafpNEPWC+zI4GGAojsu69An
6m/a5VBLkHGGD/jrtuK/nNkdA1zJLDN320BhzjctoBOCuyk87pncU2/k1B6U
sMvqL/WqF3BqyeR0NdaF5GKTahcG0zkk7PsZGo5uxjUspiyZwfg2gZi2Gweo
n+0TfBEJaJ5AHDUoWN9AQkj7SedETEyst1Vz+ly1SgBiPA7Yu+b/fWVes33e
jLIHsgNVqBumLfO6p7Wh6fhLQPpHb4NRxJPSVhTPgYkKIksL1BS/NOGvvpyj
SXAZ2FiCQWqUhbjJ/0KJWD6u00IBWyr5pGg0x8zLWGl7JQ8cSAo4Ra4Oo63b
yWKr/txUi/yqMLWPzuW1aqm7iDNxlp6Lppupj4RISa3pYQ1RglFgrrgcygEM
zSIWm7ppI894+iZw4MJbuUeL3s2TWRZf/8jmyJcZlUS5MGhNxPEZLyH6qC9d
uEx3REspR6xTye1zrK0cM9KcA0TIO57KDP3AwVzivNtNSqPqz4XkGohEppVP
cWciQg5HKaLvEbr5pEIZE9u7I/YrzPHHXRosp2LM3ZXPm8+iYV0zfnKAPIoZ
Zcib5/BbXVkMn95I8Lq9k4oUDE7oQ8c6hQnyeVu93l2SRdjr4S00y4JCyS2Q
mzEN2SRr/ptfsbrqDixcC4cUlsvDlwURUoGYhSBd7wKInVuYVIqrQko5fnA/
YzlU9wmRqY6vrl5e7nl9Hidk1snCGPWUbJ6aOt6oWtBENSYUXF0m5czAtLvi
sXFIctj6QAvvJ72RnkdKPQCZQPpAmfIwbUw/dDJzxymuFECuo6WNo9LqiYSO
+OMoue6PEeBoctSzsb1ldX/QEbzrR5ipQac2G9pHxPudO0dOVBDNxwIqTau1
7gyDxpU8xxgdqB9yQV95fQVUjM9Pm4ILNjoAx8YC0dBD7Qb8N0y0ikicmD/B
vD/9/jPAe7vEPqUAwtKSH5PldIFuZRNmZGTcYMgBi3tbWdv6EoxFNRyaj/7x
b0RUx6ryAvVuR13TpjstISDcbWh5C43kcNILLiUxP6xk2vAF+8ApuRBda+Sb
CC/eT5dLgatMD8x/4SPEeKEWhUfpcDRDjiByFliwgL+kpS55B5hOyoArms5T
AGq33ZIRdsBWXiok77dOwASaEQu+JmjbxRh9B2j8C+GEGQWnXcnZC22BZFGP
2qgazLnk+pZ1bFWqq9xErE/YUkkI+MMt6K3vUY1byCNINxaY2SrvNhhC58vl
0dz2nd2m3YLULBTQL7LczSZ50NPQ/Z+Qx2KQl2mStcpfwJ1JxUTBwlo7DClZ
qjaUxwh5JMcr56hEQ9RphEUBD7NVLYY0JsSkLOlYRIWSuQFOeuxU2f6FZtR8
BVH8xvGvJFY5WJsv0HLwFSprKIpEVakrS320+9zqd3gQ316qlJgVvjYikzpe
gHcNL9y7/esLmIxijBV0vGS+JkQadYW/7W5Vso+tW66V/7397YDhldjWRsgT
u5oUflZQ27TP2BQru9PQDae4Lca8exm9WC2Qu57tOvYMLlzYzE1AoAv8uPEt
hG/S5V33oznngIakGNNrSjxTU3p+729gUgnlokpKSNIkbGFFCoFsSixiri/u
yfFd/VPUTz13lz4eJOuGBB2qW+znizXUN5p00PDaX64cq47VFA/PLchi09RT
nlT7TEBW841w5EJp/zJkQ0SziyeGfl0g+U5wjhoI3X26CooZHUvc49X8xfqO
BMFjXc3uTgxvJoqzZs9KxR6/Tpn2oYEKOsCHM5f7Y4YdvpxNgETtIIyA8+VM
f2EfIKzs0HlY7+k4XBXjpz7x/LIkBHkO13ZCtA5GUgL/ZOqVOyhCTtNmTmQ/
cdStEribJPl9J3zm1NSMcnFdRcso7fQppvkzSUfen8mxz7oshRsPdlwzojor
i3Pp6PoamRAOl0EVX1H+4TVnobd2Ci6hE3KbdA6kE0aZuoce0nULUAg/ewm5
uuVVQD+x5ZItGnpLyIwDi84Sz9GgbnE2V1+/wfieqIim2B+3CaBdkwCqtPi2
lHdiqNEP97HvA5su8TKcxAcPSlweOqEUEGRSLh9Pt2T8TgpLv7S9bQ6fHb9f
oamV/DB8Ayepsz3E6cAPouc+ESo5eJ+5VnXGITRJLZfS3+0rMRV+wIyYVpMp
JyIPUYrecO/l+7V4iG3VXj9r1iclXlu8Z4HKvaoGV+wGMIb9vJYpwoYN6VYT
sBIHllpZnx54T/oiXyfhQ8870SjiPhO/s07QI84dCx9pGU8/18DPPhpmHXEH
HQwv+7F7FHGb/Yo9bKOfbKQbgK3ZyoYyJJ0vGNGKgcIs0IzdDQVQj/5MtcaW
p5N4uIe6o9YRCTMXntRmpXsF9YZ0PG84S+LNLs0M6kujhtyFmDHs9zESA9sK
8NXPAL8Pl0S3OdOldPZ3dyBtyuiosQqdZhM11CwZ9TTWuTSxjuPXXoFZWpAh
+ERNdJtz9n5TOIf9ornGGz1XS8tBKRK5cx+nMRtrACEAnYQ7GUajXQehE+YL
TnUGYwFFyxkEGcYj9T0qpJJd5RkMcTIvtXk0ccypI5CMmGSan4Y5nvV6SCN3
m/8bQcdhUxKC49LB8sWRw+Yk/8DzCHQhUo+zNbkBCe3S2jT+U6RGOO7d9rrH
Y00Hn0vhIlV7Oa5s5kcmAR2GzwDZOuGAPl7yntBpuDq0GNdpYtVsxWsHlG8C
M/U0gFNdcIUg58sKBWAJ8A9tbtBQC3quo1pZuSEAuqj1FiFMFDkOcQVVTXiX
RKIZKa4yOCYdZP4xlTIT590j8F/gicsZrWH5WEH1O1VJmz17cvuZh3Yp7eAD
H5s3+N3RgtwOsFX2C/jDFtLk/+z20keH69h35PKgCr4b14PKSisv+gc8KsMr
oU/i8DSVPq0ncUPBDmRwqZQiui6K+j6hU5fRnGzmD47owmv8p+kY+3IK3ob4
5KFVwDbHY3M1RRKOtuo0p6bI0cuxJ0eJTV5r1VLRf50K8eCTbnH8OmvHO3Uy
RuoHruYjZqTDjP1WGIoAdTREsd8d+MXWUzURDF0gLEGF0jkVADUIN2LPtZkM
CueaTEu8LVoy2G45d+cLuj3HmSiOffl7YL12m0oiuHhFudOzMBNGLVrhfKIs
pG1sd0pReEbcQhIr1d5TrRmQFxNpT9hCtJWJL5o05o3rQHxpzg/VvtY29fMt
a7knzt9euKHp6eMufb4p3imcVbQdOxE1Gg+2Fytfl/sTj/E2++VTRJJrv8/X
D3qdwHz6teKlhY5q4aWaGgAv6CrlUEZhXH6fyRTmUxWuEMPBt/KtdjdV+z9o
QOJ2dEJYm1gp68GXzIt9td6gAV2zF660XKUV6+4wDklMt/q2FNykRh6mVLBe
TGR2lK83nTP/w7fSO0S9IydwBi2QypC5tJPt5v9jyRQPKS2rGK+EYzFe/7xo
Iswpodz9sO6AdN50N4k1cfj45UhPAl+peDQGljIXj6zv6y2WsJQGCPAsl+Fn
mD21kg/rps98eJyqoq/F6KT5CCumRNPqViBLIxwGIPlpGjOps4kWFnw+S6ZN
VwRLWTQYMMCHeAIARXHR2aCdv/4pFnRj6N+XBXK4l1ApRfK80DUn68Mvj0+Q
z/khO/fvQK45QLi0wDSQgvTscgqqlJlle14rfMCXK4ynmi5X0N0E/71j7OIp
cqdwzk6QatGxFJryr+fi5az+hMvM6wW3VIWgUUL0q0xcNy1hhR5V8D1iVIfM
16ZBbUW1CHD1OtoFzfEp557U6oWRcfUtRDZuZiTzvqOxFFFbdKan2zqvBA8c
rlo5HTQVZWzW0Mx3gTrou7C7GTarLHHNyhCeVIVxU1aEXXuy0yxHX/lFMong
mjxkMT12x28DqOrVtkzVz+ppVxbuyKnjfSyB5KX9ixmo+CJiDwQjuLXsER58
d7QKHlVskrViEzf5lK0mrYuCRFO8e5geJRWvpz47O9P9eIoBVz9ubaJcvQC4
g1bvYln8Cl7Ycefi2ObSVxpkSuKyX77vRpq+O1BPfRU5fYKq6XHv5BXLjX3P
whNgV3Z/9vPeSYr5TiKPyYIYQFW+faDh+JToWFqRBsMWkmF7ZqU47naQmnQo
RdIJ4lplHn5B+omyehu9B37LKhqRd7GEsPEmDQOYH97d4ByzZS+PByqJ5E0E
g9yTRp2M4+xRjIo9vbCiymYA8i5EfyoYkGIe9ONEZs4xwdyrjU6i0y4bUast
FyydB0E5JG2l6VGkBcusQ6GuLZwvWqv6p5s4weKWls1M5fy9jl9zjhvxTGi0
3raaHLpYrZS+BYw/dfHKU9BxwT5JkHSl7VvhRvMrfv2GqjqtGnXFtidc+r33
xUQUa11qahiXC97YvYJmNxtpIxJf2Nrzwe3pxunJGOVBwlf8kdOw5dUO+PmK
4kXK1z2kvG0GA6hW7u97YtBmoxrY+A+WMQ55Z5g9GLPnlZn9w8CjYKbAhYez
ykgP8Olcjd9x792rk4wP6+Yd0KfodA/QfEMJqcgDbfKPu7NqjJqRyzp1fdtR
ubZ488EtNaN+KknGLM9/bLM024nrvOwWGpvxctakGy7YlxMTJ3NdbwCYGmhH
QC0yYMqZ9wTRNlvjPfq+xsGf9O+iLRKRzhBCbzbnAlVvc7yG8LmDSfozJ/BP
24qBFc6KpH6PRCa6R3eGnsK80SzRRH9AxU82AqGx1KMBGJ5P5nIk7QUSQ4tZ
yz0AID+mt3sykeyWnsOY76eyw0x5/hMKMeJCpiaWr8X3jfs3U5/PFeKpxz91
rN5fJKKk/EKUDq+ljOyBL25a4XemxhTV2LqI1v27+AqZHIUoAAGKWLmU7kCo
bNRB+7VnTKcPMaUFf4V3JJuIQKe2simf5cvJyJCUzHSbcqIBFFbTUsXt3DhN
5eszNL2IOYrZo4IeEbOzkNdZvqE9vJgxqC8+cf70vk/pKCntlLdv8JmPytPM
gi90jQkyu686QLwSVshDrf8fhpb8RuH6Tnnb8XpVWvmbw/j8yRCWXfYx/xJc
u8fQ/bLOnWUaigWTp1gOfF8zPLJoTlqQn18NSOw3wL5hFjTbai1eytjdvfUp
SYOM56Hn+EwK380PUafBBoJdh/iI9sIEu/VZVXPFugEQ7Ty6pSgwGQy/kUUy
gD6MR9ZTRFdNDL0ADGwAGTqvV8NI3JgiMlt02gpjuHBYmTSSZJbbZk29HIxA
f1pF2Tv29nyMzD0W1YoQQXhfe2qV7qoXAG5vT9mkFSKcjyEeLWY7ush1GV6d
ig1RbrR4OCpX3buH3DwOWBTOa9oJOmGYtG+dGdc47t0OlOeos4JNf8VWUOUt
nEEFFARvUMxSau/JqYv7n1t/UQv3Cekuf1ZysTravjQ382l/VtC+J87gXlcX
GzTjm76HKAuHicuYel2Cg8HB7fw8SwYsmdhDyS5ZUIABppMgZzxsRI3Z5ZUM
l+zvQJEmptEXrVIFUz38oAOOt+NZ9VxZyhVL6gNevm9iIV3arSTjEJ8orKtf
7CMXsFO9WT65vLkvwDU6De5hBGoscytjo2VqewXzuwLpVsRkrnhwA0ILF9EJ
0R3YZs14SVleZm69J1j+XfGTs8GMkHYmLxB3CV2iYEJsq5JW3A6RzcJJeR7P
EwV2Q0/i9mvNCFvOG/rUZ7p60blQVaW1zlpzSW+xHmFtWQ1Yy0TGFEPiDgcy
+AsdcbEr3vZJPJK2et0qFcYvD/no96Xfiw6goQ/678bFzphHtn4wQ1dE8OvR
NM7Sj7oNQtKgjCQBmHL4g8D+7EWRJqz2aoildN0yrZWz62fp1MIbt42dxcvc
gJVaQYEZ9U9pfJy6D9ChSyvtBA6w9Z3u8oTOlBxLP+HTxTIDBBYkOijBU+41
WyXct+7gWbU4tQYHBeDX422weTzAgCLLtK3ChYxhogsDVWCcCkxKpgjmFDrC
wQJWtzQ7kDOK3pCPu+mG+Zxl33oYwPWn0Pir8GDK+N0d4LY8NsY73VHwo4Sh
NMfDeb3r/DP6eS3Mmv6lwXG1Jy55hRR1qhn2buT+zeD++yJQRm38Al8+Y+Sx
4khYe4O7EI/HLkBrnoedsN2Zmed3OG7PdBStQzoHVG1hKWacvf/7O+RBoQ6c
qeBa+g1kyEmvSOowwe/JxbcDw9RPttilEzxagISQ7ttguYo6Ri9PzOgex1IJ
Au45Oeb6BZ/eMTfD8P+gzjStLFiYJPpZNTttMQ0GFupLw5vsTQLpZbqRIv7F
ruJIEbazz++K+087XQb0pfceO6Sjun/08RegFNvD4CI2Sgo6wtW6z3LjPvE/
r6YUDgiwlgdfiu/La97cC0vwiQ0Rz3pgjHNgSPvNvwlPYyx4ZOmk5KeSFQGe
vovsEg63juuN4gwNje2hxU+tAd1ETTTPowQQbRwoZj6uCq2yBgdNtgkPsHJM
oMsa78qD9d5e+mTOI1LaqsPfrxiOFLU6qa6B0iAiIlPMlZsjLkzAvXod3UMA
9UiwtRnIsXGTWFgeBhbfAvw/uMfHjyN27zMsGgg+MFo5dvJH4QTQqE02BSW6
xV08gZlbSHFd2VjnYbJ1eEGNH07mzWmiVYN4deusexxQ7ABCzLx7P5jV5+mq
02fYMSYj6yaA5b/svl50RYtg4tSJyDa+hkKssZFnzRg1RJWhtmYAHxYcgbvu
nfO5Vz+zH8OCgFZka29hgV5BShdVG/kL+uNUFPtp/5gKsXHb8ZcygK1dJRZy
plE9hbal7keTu0mhclvfFpPBFw91JZNCnKMlVyaCOnoDNs7H/HllSPisdj+M
PJKVyzcFoUNmx5VCILPpfSqmtVJgIM0SjrxU+R5hg7mTlherqJVaC7ZMO2QV
2gngkoCAEzXLYVGJSLDIsRiSW3FSfHy6FeKpkbR7GJPYZeLoaSwz3MMf6Bpk
eSYYWMFbPdKCymaQBUWWZ9c3FCexfz2LpVKl0SeFRELHLz065B5Tnuj1uvRa
CeVBYgPYi/du1qwxE1ET0My6sV2WQ3Qat6HbVrubV58rJQxDUaC1Iw6Z5ADD
PtbI78wPE8O0lb/6A7skpdeAVay3boPiEXuuGkooAe5TWmbnOmWSdi9Eo+qx
XKmp7RuehIrUwgCTuImh/dHKfkhx71mhzclifsIWOw1TaJXiZ9bp8Iw6qvix
yCcO73iUhE4pYpYHv76QE/rQHPSwIFxZ7W6sNUycHNw1G6wQDB188//ugppJ
RxBlRh7+ZocwkEpGHiIQad+F+ujtdGKDg+inOF2bxCbn3DHhd/EjuLc3ts0m
YxMoY3/W4Bl+1rPXdWKpE0bkPAiRyNkv6eMvTnGWaM4XmwyClUprWQdMlfJu
sQjZWXkEYPJ8VXHCm34By05rFoyPBp8eS/TIV65Ox2dQT9f+yPC/p5+k/Y17
nRtbzblxFx/QFGNazRznQScE2Y+24hu3jTsmDQUJNvwrv0Iax1a//04xCSVc
yaGIZuBuEfYEP4kH1HM7hrBFzitbXYo51ToqB7Bcix2C28KawzNf+zNE7pfn
ra86Rk+MxrANm1KMTECLIGNscVDF4SMn0STZjgoKEtkLB+568iae3H7cC+pn
QaJ7ydTMFanVQVH7Gi3KkF3aP4oAMuwzUwiwoTtu+3IpHux9EuDrbde0MCJa
lxs10GQjcw08jyeDtbGiO9P2cWQjxNb+4LAJUqjThvJGAIJYlHk1d4misoOy
wlWTKJmeJua+B1Bvqv4XIiBxehLTZ2drqB+Xras+g4C4H/HdcZJzveqQYVUe
0ipHiQs6jUvCJaFmhyxoX+7w0Mpja07flwYacJVBQYe7AebIVXnbPjO5Z+Qe
kBaDczTHE/Sv5bwZYI2mihYC0pgj+U7bq9o48cE9S0/l/N+o3vZm71ghTHiE
J6KlfppjG94cQejN7u2FPY7y3sI04+edXvQf+J/kty93kqEXy960wOnpulb2
lQekXMt/5ax68Df1BF4RnN7CW7ql2/AxKS+7DpbuXSotUDI9p/yjMP1PXpI9
InwLHng5IJ22Kom9A2FmCUfskFOAKN31YmEEq+l/XWrj+Big6qwhEe+OCG+N
QQzIoZO8YNVZFUsHuXn0Kl4NEzU5LAstN3Jbqz6CYihPkPcjo4utTFmX7kiz
KeSgFfSTJlqpI0A9HDso3MHSvs7K6Yfx/oaIMA+WyhpiZv36LAgNnej2JOiV
IbUkL8EA3GJZWRNy0hI7JIthZvJIgEVQK8kbiFn35esFL1jLzhlC6zD6vmWp
+oE41Jl+8i03d/QG69CKIeUn9OTe5hUKApAEzJUBAFLCISEDrGEZwxCtkG/c
OnR7ucoQRabEpa1SBWhMBgzAPQNIxGSFKkkLxP+NEKxLGx2vK7F2icr2jqgp
osOEOPgTlxSOlqJ4OUYnH0StPqmsTEaqEvy9NsHFbS84uWPEyyIdH4sWrOT/
emU6+MiXTxRL/v+UMzDFt9n9NETnXlxdzR4N3+76gt/R8u2hjc9XWiLdFlQN
2Ja7BHZbFLwRjln+zWHTNb60WhuJ7U6D+E9RmFaqgxLpXT5f3FrYI3J61fWB
bWFZU4Q46HvLdF6aPDtmO1TOw6zRKgayFv5BjdF8Vrg9M0/542MHD+O3i3x3
zRIfVYFTAnk6tA+ZatYM9ET6O35DURiSIoM4vwPMh+R77MC4BLZ7WJlwC1LE
YFLgjQACzThQK3xJV1wnqUbB1u3tmgoFvITXSWUwiv7FWMUFaZ/K9Rt6/pZu
mSX6pJsbV9mZUyjtl3ejXVTFV5DDZ52d1l06SuRcwxnGkDwLCXIWa6IxQ/31
Jt3BXzG0Mk2fhxA1Xwuzee6iDgJq5WpvSH8BSwCTsyxruLAfdwubwljF4q3c
Xj3kn/JgyIndxyRwxh53MR2RShkgGHmCXY9wScezGgL74gxkQjThTVuHx75Q
nIeDXQnRlFInyKyUNf6+1uv2BmVHjz79cwYsEgqnnvHSGw66rQrJ/6AS3f9m
YpAz8hwJb1Mt0+m9cfzlhdS8TJEYMmXgFCBWGA2MJ5bNnjNbBEdYvQ01Mqv5
0cskAIQNAH6OPW4+71XC1Lfbnas6ixrVTRrqENhX1jCLaA3C1iKpj8bGhPTg
AYvZa7ik4HYgDBfayZ7T5MCJ5Msic3tUjdio0GyrmgXVxEkiDjVMNjDiQs/6
xsCG9LQMWpzih7iahMxHKAJHN1gCYWRwmNS7aP5QVY8J/C1UhOnfjeoBXxDE
Ookrwi5gtMnI5ihBmFvdAO2PWYmaEbNwWP9XS/arMz9XAirEQR4iLz6/mKrs
1uEBuKqiNnQcN1EcH4iRWqmDjn2ika/1C8yuvTJSqKF5dvNpmuSGs9fFLZUd
zJVUMx1e4wOMaQoFAyMW2s6905oePjztQoqjjnnHJlblDaph4oVAi53FounW
c3NR1Miw8H/s5xSZhX7jsB47NyuIOzwEfhGEgu50u4OsEyIDispIi7gcXxhN
q4q1Qu5eHD5XCR5oakbXqhvrem/sZp+qyZxN7N2TRi1d8HfuDFPgwvC24+Ip
UT5vBWSlv9GEvm8N9IAtJwnNFxuseFU0FAcKLJ+1id4wW6f1ZTn+tfwYdl7G
LB1CyAKKgBdy+m10/eJi+BhJVjLKObpR1AOGzpPzSOKescB/ertwuzeV+Bo+
SHcKDVqFS11dQYmxqFIp+s9E8s34g+zDP8bReQUc/ulasAjvdo0M7xbBSW17
cJNcEY6MgX9fRinZIG1OXFU0EcJRTs5OW+nwvGsHOR7K83CFW8ho1/PVkzhw
lslH/Z+cbk1w4ykAG6SCTm5ZqlYFudlJ7IEfX1EVlz/5q32agpcXbXCcICIF
IjcGxsrQc73wQIeKXfvfnejC2Qfjg9DJnyZr9fWqO+f3ApH5CuDCcfthuxfd
g6MACkB80GmYIcxNb8bPSlAxdZWfSZBEOOEZ+PLJwIdWtym6hWQHdmJ6uOWP
TBUczjTaQ60eoE6k1/CRAKmbwEoWzW6NT5rJp6/Gc1bB71+nHWl7irrBWtS0
Huax+63+fSM7FGsndjMNqOG0FyvR/wrtOAvG4F+TgitlQa8hDsBpQ7oBz0W6
zoSoGBgSXvBuFuNaC4wATG+kfGvLeF5FQ2vq8L29OvupX2RPpraWu+Jh2gVy
bqfVg98+T7zIAxbmpJCA3tX3TpwhXqyHEFTmq3kqT9X45BRpsVQxAWzFFpVi
kDnTLNDfOxXccysRjib9cxGsm72w3Qxf7bHsyoJ0u3vH/O9YCiA2dhGdi8GJ
lXemrl9Qe2uGK5gtl8d1pvB85NiYX3qAAanYu9VmfoN2yEF6lv4LoNIWHyWi
H4MbdTYzqXSYpVZcgq0NuBIT1iWHygpBQmjHHZxx3i4T8hMD7doUKCRQfZrp
8MWMFZngLekfJa+0F3WU3SLN5ZUOxmb1WOfXnwezWneqfmZpzIMdfvU9JD+m
yr19MrLNcxnhGAej2ovfIUIQgUQ5YnsB9GLviZF8FAM8LwAI9x6R1dbfpi8F
J9lbn1xc9brwsVprB+HGSyw7fnDwgvJWTIk01F9mAgn/nSDPblwPuH5LYOLz
gdzBUfbZeodzuHzfgAYYOHlYTL4Mx1HG1ZsI11Cb81wt27eXyw55zIzY/3d9
H+uFhTOK27Js+dtDyTzjkuE8BLz5GjxZ/XaytA8ba4ksR/RH28aP+T4QSnxR
pNofbtptcMZ6gAB6K2zuCOvvb0+p2ytkWzGuIG5lntQ6pPe8zQpxu0sZIUwY
Q5l5qVwb/t/U6Wqc3tZpKgrj/TSmDWwX7vaLYgBLNPAwyaV7xwd2As/v2Y0t
EnCBAjXBHlA+bF28+FejqGKfIgCA3DQbBRoYIq0PNeRiWtmWQXKwODX6jLqA
d8PugYeyOZoKvKDFFNSl9iDp+fY3vPFwK8xaP6PIYKn2ANxRB+8h3IOmomnZ
vK84zrk6rpvt/x7UWzZGKgkt1OZUPhJan/hq4mvbwW3LuMjxKayyV3ymzxsL
VAwnpezrVfmM+f+sYSdqhCNRaqMxlZO0iqxm+my0O7h7BxjGT4iznQGI5Hj1
pfEk7bNbV+wuaD8vupuZr797A5NwyaMG/XVphV6uS+LnQ5n+QY8hJHdEI51i
UUCuvtDEPD1FN685jANN9lm6Eq7R9kkZCLwtbjyVFKZqpw+ySWHdlTsY9lvL
QvMrcTDlGffe4a4jFnAA9ESNypkVu+rKUetFiPmC+rLGPgTPDOKVtnl/IN+k
Qie6hkxMpvX/SkreSL6NXg0rfzdaRCTSe6d7yBFdZs0cQ5QK6V+M06tGA06i
A28xMq8dkWdNl/LdGVS37BByOflil1XClWHRs0pDA+0PSY3wz+BaG2ZXSlMT
qJoWdcHc5Kwb14XW9tAUDyx0Nwg/KsLu3vqaQzlx3IRH2PlRq3FWcGOEyuXN
FWqOaxNPqGoL1/eXfq5orBO9IIRaUer6oKUO2HSEyxOmDzP94LQqjHoVVyGa
7dcakH0fih87pfhEYSMWi7xDA9BcSelICcBKNc0IJfKM5Evk0GNcOsYi+f7G
t62QCKeqibXVq133IVrNKCm3EbjmRME+7+dd88LLcNRpAt/3/CZSoYMcAKhV
1K/wRxINNZa+RDitBIs9kosf1T9ZOZxMFozyc7vpukatAmiPZfhF/jGM/UKt
xU+XBI03vKBThEd5rqK4xO9g3QmLACh8zLh5aa3tKXEMhZPWQlz6Uik42imW
gO6S4mhzzolS0Oxh8oud1SK6K5rS9SLCUgs2pfJC+an7DppMwRMhImiFmxxe
IyT7q3twTWATBs+e37iUmIukXOkJM8JhnzWLkP+2Avb69CEdH1ZUqYbAA/E/
+9Ic+g20vViKaj/KB4Zcu8yL2GKh/DBYtZyHmgzdg2fBR6ylJ5XxlAvd9lH5
O+0FQ5Lgp+JjIDsXqnDRBm9hr4aeG0UZFqpVOMpjIk5kRZT5y1kO36zejpfa
Qwv9XnWrtZ4t5SQDb0pgRSWq/B20AR96E+ZJIg7b1w8pGPOs2L69mNzLvqOM
khzrc+oVepFhnnc9x62BqJN2E4IsJgDh5AMZqOgDEsyzFtepU0WpF//RtuSV
rux7cI0uK3l1addmeq6/MOFBNFj1Y/fin8z1HpUr3mZvtfmmWaYPZj3ShE7C
2u5qtIDfWgdDsvD6qwImB6laJWMK0XQ7XSjCCmqLDSOnjsh0M8RYjMSm7mdV
KkSbjx3uTQuALo6Lvp/H2rSOgPfG/2/dpSYGximX+tra63o914wR9AmvhXgG
uPhyV80ku1EJPQpxUfJK64mQElcNiW7js9mMFQg+LHCpCImI7exWC8a5DtuU
m1aFZeJWZXy7A9hPL+VvgQzeESK3xJkac+BiQxfDGs8hY+nmCzZAFsAo7Jty
85Cj7jPL7C2s8ZVWE/mQtBYyNogMetBZGnNELIkRymZ/byw317ClxfLTXMPO
kHPjIcH6gW25UPV+w196wpj3tjvt5EEFBQIi2cNyUQwyM9gyROmNDSIyEGJA
UVbamoQm+IDN8spbVU5QnXV55lFGQFfJB2YnMm/6VXJtDaxUWRAm52mmDs0m
CgrD8VlaPryxkC3vN90zPVkBSRwVqO7ms3OPBi+AGiN1hDUswOsAgV1N969Z
tMQCThOybzxml2m/VbRavrfoVEqtEytUv4z5zS7+idudhVjnUVM8W5qOgjrw
I1EdleIpnwsd09OLLqE4s/32eglFts7Pn8ueW1avgv3HTJpy9a3+zQL9fkM6
g7AAKq2WhGytYeBCOZyuPw21sOPMU661o0iQ4nWlwe+n4PVn8+YbWYV2qRCP
joYUA9CJgIB6z6S4xrpYGkxaJsFHnETsg7E5g5dZprut8nPelW9CTm511Mph
OVa40gmCe+xA6cG41phxY8YonFs7Pit+61TxSagmGmMjBsXeV1xLNBgAWYkb
YGQcUIy9rnIeb0cxNJnCgdGynWl1XWbU6ngAblZNRJYfP9DX9/gq9iVzTPXD
vudcStd3QcTGA5hpgbF2HxhXDalA3dMvqnQLshM4OkwvNGTCmko1xO7kPAaS
1TemyZloCy93YzvPl434PsV5yRe8LFI/e+Ju32oPqUAuFJDqbSjiR8CPmlPp
qiX8zheeTpTWhrWcUpkCZyzgJFn2qQ/WMj1Tn2/OK6cJxHeI5c1bGGZKab03
FEGU2+7wyRji1CGeWg685pduj3BR2rbrZcLDaxnDtGaFzQlfH2mN5gJDUiVd
0ZeXIWSMTAD8VC0WvT6MXm9t4fr6F1VV11mMw34yh5/LcMoQGXvttmagN/8u
S8us4RgWHI0V/0Aqi9tYBxFmTZaKjLukFoGyldwoediIMRjmfPzjcI+h3HRF
z8VL1jgCP1zDE8ZAPMf5soRpAMNn1NWaLe4QfZx+OXdbFs0fide0X4iCl/gh
RO+CuDkjJy5X36cJ9YF7WJtE+N0MDgLUapy/Qcs+yLP21/WobCOmL1ogWGXq
QyX/RKHaJF/n0yZvLpx2M0+W1FlRBwd+yt8K14UBYtppLhLZIlFvGuXdEKQU
T5wlY2EKarmoD+EFokJNqYtvT6sw9wVOX5QZA2YKK/e4PQBCCfqvkUgJmsm/
uLfgghlq2y1qiKuWSVkgOzc6ileSF6PFNY9oc8pdpZM0pYTJb1Ta45pK+77d
JRJP3O9TzRDzq/gdx/NodhZmO7mf6b2okffFUS0KTrPxMx7RfOBFWUiu3Tu1
dmyQzv+1DVaPHX14bRhDMJSidriiz8rsI/etO1h3LgNxe0IA6i5XnMoAlfkx
pU/+7r2c+7wOUNFKhjGyJ3urM+6YIi96AkZd0kYaRhEoAP5JJNp1jERWXBQX
5zZFoR0kU9FD9EPwEsqgIpE+9zUsf6CirXRQ+FOZp3ie02yH1OAy1euSzZCe
TgLBcg6rq/bqEQdKOGmPvfkDdpsiMR94y79Gy4ArFFrsH90BxWcEuk9gJyp3
iqvZxaERu/+I9aLklHBeqZTRvZ7yFKhry2UJWcYjFpk4LV4TnYYyMs3LOePp
zwx4nEfQHlKzuokktVso+u3Or/k1fjeeaMI3plyo6HUADWbi72kDiCQyMfO/
3ZRqQRlfyyTjRCVO4Gx/ZDv3IMUaT6SxdRPDMObnzPx+6Fvc/FjGGTEn1xlM
wKZ1X62KheUryuu0YCVDkqTpFHdJg0vS9jp6suR4ZWRCjYVeYTq/BANXqIK4
+zpVuPEHn8Ia7UHYrsv/D6wXW4cysnoJN51u44wuocfdo8PmW7LTaXtSMeYK
XTQ3ln7t77mT5c0VMlAL3QCLsl8rp73Ig8zF0uFWzYhGEQtTn//Ri/5Sasen
8oPlxroFvaIGdIfbnFgVNeeG1vZqmAcJ63228Kmr7XYJKLfDvOzojZAvIX+E
r6o1fG8YUsBxkauCyTK9venYLUbH6LewFQI36EthOTHnGztaacmpHEM2cRmn
kCOHDSCE8awR8oLt89f1XePk8oG/esfOwz3cOyQPu6loUCSRSqaRW3h5UG5o
yDfrMDf2zeNPlmEdhJC22oPCXXRmBZCf8UkqzCT04Pii+QscgFKLI7KrdE3R
jAnn9/d07Ws01dt9aQ4x03uYcqmaBVIsEEFn9QeUU693pl4pfAi4rkAIiH0e
/yrEwzw8eLbgZhxz2QXuq77YEXUS1/cpTESNScZ4FkVkiUa5eV/cPQhQ6Cxu
FDojXZb1JdLUMO/TlIA6MstIcJasatSg7lrhtf1JSgnnl7ZQfvw2dqccOoyt
Q1X0LKIB50chOGQwZga1PV4KI7Ftj/qLgjNw8arXwlPSrM6xC0b3M7ElSTRw
zBJerBXGPJZHMPStHHFMX/OlMPvUF2xI7g6N5Z/gK8qWPdGLbqlBHhiL+J3q
tSdTz5glMf5LSXUUkzqVbdpdOVG8dYEQLQQKs1KF+OELzlxrzuawfbzHggQ1
zyRTlDIkWxMwXrq4bfcx1i0qeqVyuWgK7PQOaV07ZIRkdxfmPGybvylluGTG
q5HGblSbjjs5lV77KbaNgYWog7M2jlzWF20D/tdVpcivkKlMdWocl4zLn1Hl
NNiviHI+UyADhmurhgYC671mpgBESgmOmNx7+2iRL0UPA+VH6R3sWt3reqQX
wd09Q7SKAU9Yp+8uuXEwGu9PGIuL2m5QKYFbH52sKbIN23SUzprPNYq66yez
Ov/HpkBBgybnKioictLgY88/bcGNQ25Hfl/aZvGrAuZmN46DNJV2oWylr3BP
AX8vekqACiiAWW8jPdFjnpOd4TF8udnIZ7C/j7VfRF/aa9c+XWZ8nmEG7alZ
tOLprg8ebeePn7OMugSvZP21Bj8HC6HMSreXyZOHdVZsmeqokjybTw1PYDcy
NYqRqcqFCVbWz/fijOMU5y8HChQCai6rAfbFpWiCGMFXJfOyLuPrK+G9x9uA
FJJmiwlBpIP5laIGb7MdkrqEqwt/ibIntm3t36zOryvcQi0oYPd1nyGp7qNn
L6SYkP5FpLLR2B+AJOTQcoabbsAtCS+0cHj1kZFefoTkS2iZmTHVK8jqqQDs
1pyXYIRKvb+dHaBoSDWeyrl/7VmYfkOMzqurOvHkejXndrrKrFIxFimHmZHq
BShlT9AqTTZXR5ap+uNGQM5jdxFYJRydKicwX8BGjpYd3w/KK3+dG2IBwvmD
Wy3WH6Dl/AYpr378s5xYNJUubWSTldbV2CfB3ykxPJfXOsy1D6o7zhBmIyC+
uCIH140rD81d+t/v8FHqeoHRcf+Vhl0d4bn5qs6SwJMY9pshYDmTP/o1A1Ny
Hhnul1dTK+7+q9nMSCZaKbTROpkHvmy+aTDZmbGX2AJ30X6lRR2rop9VGpOp
90qDMPtNTuGjPRmyUxng7EIE3mKeGnOTrPB6pMfs95roViSXZJ/xSqR/29RM
qhITOPetedrvazR+hnCS7ApPvbYLXlftjeY4Ck4B2xZXS/lB+x+ebVydpkB+
nTbYlLSoJp8x4lN9wpZJ88TnZcuOkLTRHVAj4a+0xU00DGHIHE3c7T5CMBQG
Bte79NC/R3gvTLDB4V+utnqHTJTTXC9tugNm1FhBEEjWM8D1TQ+dZXYd55oa
eML2JIoshNmgql/W5CUakEIuxMb0quZRG7s2yy/P7OnIfCpkIk/v77c0DmR7
3q9HMaFwjDR6PyQU9GXhFvDYd/Bef+nTBJYInYSxKTp9Vmfk6Q8lO/1tdxXu
ToWJ71EfTTNT36JuuUl/ZQ7OFIthWtkDJaXeGEbvIh89Anzij1WYezhK8RtU
R1T01oyj26c26MdzcSz0z1rfUcVTIQPMgrf/iQPWMl5qgm+IEHAdfx1LJ8G6
uEflIWUH821Ha7CW4jUXgp7nHOcMyfnbCPXuXlmTtHpGV5iWyxwZRl7u9EFy
t2zeQ41ArZ2ys1mv9bf6ZRROrSsXuf9OGNqeX+irG71lUvazxFKP3vf4SLCU
kH2kNgXC8OO/OG4KxkYs0mKtQVbOhNP+/xE1yv5+JE7wHx4bocrsXG1+RAIJ
ZnbxpCJFNrcABL1ja91lXHSc5u/nGipHe57PvDF+5tlbOufgP3+7BUpeelxu
+q40ix0RN3gRZtXLZbopzebnGDng9fsmJOO8QgfxW6g1Z/4l+Y2GfpQjMO3A
+rPDWcRmZH2IZlkD2+yPkwdRtS8fMTFDUE2X/6z2ie3e6DubpwLRKzv/uqc+
21hOTr8i34EvBcdIuuxLHqisDVOpfFPEQX05ty57ZKYjP6Xvd8tpzvvvBLIv
Dvz/xYsHPVa/AQOUFIbXKKKL+cJ4cSysDLXnwwPxDmP0wHb+K8g3OLpYuRhg
thl6U3Fc5lfHpIplSGdrekOXoPTXqEar61YuIw5ZjLd+Qr9hXGBSEJmwVUt0
o11Lt1VsSaOIg597bG0smmYF+Y5EzFSAvjcESGCPYvhP61r4ddywT4tY4Gpu
l0Pf6n7XFhIr26NILsa9NZRMJwCve96VlU16z+Zqfq5BEN3dwAk9lt0gfWm2
XJ8TBFvyL6xJoXDj/YlrAu/KppwzSDRjP4/ESEQCoTxjX6sovg2jhI6tMNpF
55cvGw3INroAHH5WxYayWLnx7zJxOUlXePS6O13arciB9Nz4q38h3OEyjjw8
IWpE9COkkBceIWcf+ch31lSWN2xuVsCbOdCZhIV9Pa+7GrfphlFTUcaCgpI0
ypTAIcKeftc1T3aybb7sf0BXRlpihyvAd1PFPaj4mG4ye0tPl504Bhz1Q2qy
CLWINZXk1MVwyMWi2zbs4kdL/wwIzkjZr2hTnlD50Z/limiEKifXP0uNq1aG
vekrtguqupO//NhSMRQNvOM+Fxna8Ruu9WNFCJ0JALbcRGS0ZKDkcELy+yOO
0Pj1A9IbkdHjlSouAPMS1XC6dFV4n9n/AIZsbxHMCE7ZFQ6zA1W3+8C+txg3
yFg4Bb3EloiI1Tt7m5xXIuJ8Daex4ctOgh5S8zwe4YqZDb5j5uiZX0IBMODq
4suPOETHK+bwIhlkYW22zSwzhd4iMMZPihF/sg30y8gdDJSlrd4QiTAmg0C5
FLUIo6oH+9LlNeuQegoI3R/+o4S5R7UciocmVHxHo218RTua3ybd++N5jBuZ
SmU0JeMAVkFu/jglU//cO4owmGdF7+9kwdPhg9uW2fLGgSPzTfBK7bA9vW1R
gjQX8K8v4Lwy8d2/X0gXH4Q/GjtZohndTdEpyTSrk9kDLVTaVntx1Fj0mTCU
+PBRi87n5Mrgc3JjhnMF9fW2dnVjPRs1fjc3pG3dxLS8Ex/6yCvJMR6U2bix
Tx8GrZZ7Ww2WLihYk/MxjVu2zBs70tZ6jtTWKTYS8Gf76i5bF4cnAxQWa51F
/Jsudw4iGESyIIIsiEPPn/pgQTW30pC8YLAgDKV4z1vtomIu1x3ik3NbZSXz
LrsTRWe93gL5GVAPdbvcPG1eGB6OlZ+Fky2brmCQ/AVO1UiI0IuloUxdBzbl
fKDjgaOpVYsc/MhBfCcKyQ+5l8Wrce/CNKL6xldCqVbt3ucFbXi7wSQJNRpj
YzBNOF7lBwvnlJos3Y0KSSPomuB5e1fyBiV9vlc+vyHkeou1R1H7vFc4NPgm
t09j+4OEGRqFoldyZlHpXauKmRj1OOnVmJAbcR2QSJ+rM0Qknacfu+sybhqD
sea9D4yFCT/zqVWGg2nrBJjfGKrMSn73ARCpZm/yxfNBzjjD7zObpx02cFDO
i9n1Dkv9ic/+x6Qm0bva7FslRqVrwZ5JpieeMxEBgUYkipEZ5HX2neI5iCgc
xTj+e1aX8OiUcuN2Cw4+ZsE7ofmdgmj7l29bl8crEZ5pD+PnN/CdcWQ0c+Lx
VsGwvbYBOElbPM3bqsMDqtSVe6p9HtvbXRaNcoMmzYI0bJ4RWzUZbazpOzkn
lhPZvoLBhi90HhS06sfEeGJcoggGUfJneja7cOJfrjf7YmLeeOpcSL9SOfDz
s6WLIcBurvrXHeie+G0lM9ZQr/uFKE+dR+Ru9HtHxygHMrSrQ8Lb6lMy5Ojy
fNey5qFzs8/kQLF93ex6eW2hnVtoU6mJHa+J6cohb827WCgs29htCGITi+WG
z0SQFtIXLfN2wdzepeR2dzmfvZ1A+yWYxEQhzo6FfSOYlX8hGNcKgBHMPUk4
n4Baf2W0K4qdEkU/aI473Z1TsCfW+n4jBCVsjwhjpCWeFYkVTEzaS4BOGLCq
gTzHV7dEXALexQo2Ses5ce+dIMjjPjTO39gGnW/TDP5yPmQeHInDZ445EsB9
Md96uHmNfQfd19+pTN0HccWXdvZ+5BuhEMkya/j84oFMurYuL1BEykGvCBGq
buTW+XvtqFvghTN0ENSsqxVcv54RuVk4zfZk87Ju0aGSbxGWORbcvMEWlNsL
iU0vd67S94gpoUB9bQ/+Pw82N1kb/4dn68ftfOdA9YN9dDRix0cG2V1fqKtZ
u4ht6bxNwGA9mDgOYHSB286hWrX/IluBLiOGIZZpuZbn9gtoIaOVCYk2oFJt
cxNyiTtBMjJrgrnEyTdj4t6jgzOeVjzeC7KSShPiP2N1McZYcz5JgDICIokS
W8YZMwAQlDTX3/36vCA2SZAsNmLN0Cs2Z0OjgTDUh0uQRO30Bw6W8oHA00MW
My3P1hrWHhhkYRugZkH2yd0IOtPH4r6UUpVBYjhI7AGZ0kJPHmNB5nExdza5
oM9bmo5LzssNX+FumvZnJWiu4cbMEu/MPzsZ2nxdGDVPfUs+J2iGC08gd30t
K/PvbZgAn04Nygj5AuyRRstVHkWWIeZb/M8wtVM9slaZRmNbxxbjOlhzo5WH
gh0m0jKEx4L2oCq0i7W7tmUvwQokIKPJSHCuKp2uNe/4lDsdC7k6qt0cW8yB
uLogQ4j4jhvFSDEU10aKLNUJiKrLi3KkoiVJb0dlHKFpcqYGbJUYiueasui0
awZf88r+VKvR4/jBR72vxCHtM5vb6H6daQehASKdJfv03aXbMRsywdVOx8pZ
+7wgRKoOzuY2MErswm977J5I9qqtLDHNc21grEURt7YWGl7eqkQEvRpX+Y6e
HrB9waAyE3AyhLBAFi+k2afVU7JGQ7kPA+RTCJzcL1tbKMQehXq/d0tDbt8I
8KE158tGJIYfSARi4bQ22WZem2csUqQca0J4Aj6BN6AGkJyX64ryH6VVl75f
+ZN3bOJbxTUCEr0BojlWTtSL4HqYXR187syHMLYIapi9wgo3w7HM76zwqXR8
7E+8xke3in6opGUpsJMSQg9ZMjobOfcbjzxZZcwgPy/S0Ro0fbf1Jt7bvyVd
zUE7J1sXZEuV1UxaYtPw6DajkFGYU045fmudvcET2Hag18Zak9zgKsuLmpRm
wQImHNs8hOL9x36Chqn9I0yQSX4Svg/BNrVFnoTvJfmiL14H8b2FemGRipye
bzZJL2Z7+3v4HXx1dYTVIAkBLEGd6XsoS4Oi4PVivITHCFvFxsEiYgDFpHAP
L+4CqQ9X31JnnreJyMx/mcpWCpjF6uSLlHrH1pwbSrCO+S8fbSqmqIDvWKFi
Ow8HQEXJ4LzpNrXM3ktsE7yzZ2afgzEOyw15ggEGq7VxojWtnW2Xamhjz53h
313lrgMDMugX7+1lIZMx/pc/WzihTODGyKs/DHtqr1jwlzsOSX16GjKkrluF
Jo1J0SaH52WhtjTznh4pepNtTFfHftZx3WCwVG6gUy3lgEPF7uaSWiZjtNeh
YOrEKL/kZHloCjo9P8EwgWWET7QXklcDn2rmALmD7hZTQLVbEAh5WbUye3Jc
kOzw6vakCjz3ihpcPbgQJRWzB9MdtQqKMcryLbSh0b+lpbybOIZ/yzqW2nPy
+vGxEJahqqcVxSABO/zUU7NnqrDa0HL7nr1n6DHI1OXsO/m7AaMdpHnkHSAy
N8tKCC3Gf1fa7dDpVcmh6mpJqyV2+APWN1nUeusHVm35xbiXrMd7QD40GtW2
b3YACFjovrBmK4ITk194JHIbp0FRwfl0xQ2B0qlsrswL81Ixw85GlenksUbV
cs6zeQPa3MJT7O3nJG1SlhbA8smNFUvUMVcX0kHfcvw9TsrQF4fHpTrdebVt
cnRF6h6FPc7yt+8gh2ICcgAhglKqbl8PkzeDuGmMRBe7913A5eRYpphrjaoe
Dpe/WNzpu8PHIw9tvUCNeuLayJ9Du/12ktj6XA0Lhk3cgvhnDL+i1h0RBk7O
EGqbXZ5fIHq0df9SpXNrXo/Cb2VFGlDuAoxNWtr46zu50Q6Zhe9i2OhBy0T8
GVpuWAlQK7WrNE6cE03kH7jU4hf49dxF0rYNrW3pffjhCpqWr9QioMbaLHQN
6otsVpjY587kXRXnDA0CcbW3C0D6TvBcyZEDK2nZoXMY8tZbV3rKEWLlH1C6
yNrTyaIYDDP0zk5LD7GSjfnPROOqje30tRs6bzUBTaOFmGWuTM4w8Gw3r/w7
pLYgSgmFKWZMVMmFp8UUctELvk9vIF8GAn1xhWMke7N55/0BQ57p3ycrL8vR
NxMepVsK0D9SjBLJys4yvvq0cSTBW6ezHwKwXgxHSK7pCaSjrpvY7pw3hMrj
c/6MAQyGbRuSNV1rI1bDdpFpqqSmIK4EPLQpeN/d6j/djqI4JjVdyRGKTwcl
nTk2prKczO4yPRjRJ1rrR/DzUDBMpQzwMd39Brl1n2HuihYbvWm2yRo/8850
+pklTh9GX+CQPbnqPvfIF3q7QoOKhn6hlDcDmPAHOW0Jcq1CsS0VM4jb5gnJ
R4XFdJnur2wR+IEhYmx8HrL1mCjodZ3LGFgaQxrdPQ3IAJ76vKK0h7NaYqi8
eZREhNYEWti6V6nsCk+bfijL4XerV3oicEpZOrotwv5+z8BnZmbJs9vmOEaQ
iEViLAnClpsIHBLeqT6VhT61/lU4fipvDsECmOdRCExLOGQxhdVXLuzhoPtI
y8p+rG+V8cLS9jmL9C2OJgXRgtXuitGZf7ILRk3X8lm9VJ3eUaoaxuxYQc6K
1P0t3PVvIRy020HfBklKCW6bl3l4g8r7F4L+DhypnzIAs1SrSW8uAwgJyr/2
Kx8b2OL2IXmLB1To6GjFHv8TJC2u4+DLk9FKY5ReXdBPeME/zcbz3zlBf01r
B4Lu9zDQ9gqhyJFUbh3b4ZHdT+Ratt1BIcacGP4Fn6IQM+XN5AB7beLvbIdz
ID+aTPBWC5XA3o3vWTzwwLoWzlERUDv/QO4QV1vKHP0uDUwrXclW9ZaJJVLT
RUQWrgt68GfouyQAXWFK7WobrhbNls3vqy1Cd5tSLZaEzYAcpIZg097BDQpE
YX/8X+5V2zxxPKwBFlnptgvyYZynVRDoT7hrQoElnwp2YFy3PFl5WU7Vkl0K
h7QsOI5ZL/caOHUxJ768T+ygtfK3N+vkUZ27WknxOCDorLOmCyXyEShrv+jr
9AzT/lMJqiPPSxOPdPiM0A217n4xwzl1KT53QHv7AJKauforrEXqGOtMFAbn
tnYEwtj17gFEykjjNBw4Wxk2j0GalPwvCj5Nu2vbn/jmEi9r1idB/fUU2QsX
wT3sIgV5dVknBMi+kxvJxZF369G3ETY74u47FQJu/zjnTUn+ZhCp+wqS9c4n
gcXCIdQHA02Mal8AI5aoaBaT2QCM+HlQ6V61hsJlZB2SC7q1CZzMUn4XKfbC
OK1d3rYRfDPqrfnSFHeiOATHJewRZnr9ETxKtSgYPX3IKxC4wcP3ksU8mI9+
xc2dViPNvdiLD3zODGk5zltIdpILtilv7WlRS0LXvePNGiBtldAQ/ClPLiG7
ctIxmwNX4HskG8sf7B5+o/xWkAVkEWM566fI13C2NLDAIfgCtTwr8YWy312J
V0265uiajVTQ/IOR3/HMCpovYvLnHQ7s014cxss791Bp8FJeCG6n/qVjFAeg
l0ZtmLFEp/RoHtP8nC6CB0Fmf/Ks76lV/QvpRx0FQdPoWHKV0ywutbdb2m7E
30ifSqeOuJwIT58c7GlJVimm7rTyv33NNGzPugDlSH3yyprwbjCjn+RoWyiF
V78g03S5q7o2fl99U/82EJvOv3FKd+AQSAh2+zYJVxhhleIaHo4pJuPl/6uA
e1/6Pu3Os31xvTfR2VQqkDIkDIHGNILIMuCZFkCqrqssOUEQqVXzUF6maBeQ
l4eUaQcudW3X8f+JmwEyJmhwxmw4CHw0cdSPtcBPwxrLawLiMAXabzxIztp/
engON9G2wHA+Ejivu0xDMRLRcCX5sDuPReVluTNYwZlZbMF2s0WZWAmI/ilR
jvTV+EzIXPLInHkk5w8aXqeyvJYf+rE5A3+V41MYK3+tWLJkmg0M+qGXPKL1
fQx+PHSgNrZPttsxBBI990u4lhl/p6AUeK37fkDZ6f+6RfGllFNI3KcXXD9R
RlLpvZk0xUwdVe7gs5qgbpH+fmqMovZd3O4cbyxsbXD6F8gpeYEF7MZDGXSC
09qSgg6UFORtdUHfeCWNHvze7+PKYkTTsfc+RjqaKSDIGGTRu6M2XjkZRjIi
ULLeg3B6ddWJLTid2YJNDttNatujigUr3Y+S/eSzSdGk2G8nG/AilbT19xNV
yNRda/mD2oc7EycQ8Gh4s49yb7m+J7XlEysE1Q12/N76NYY87jo5eLFW1qFV
df/+2y6rGO3JxkQxnXMs6emE3yxguoVHylAb1gtIS0L8LXl9U3LamQm5pNNa
kvcdZ1PniwdEAfXLDRHmr/2oMySNlE5pdVCGFVrhEZAzVZxB960iGkpnlWba
XDjL5l+IvbLYDQkV2Ya6GAxOFQaGXrgKJOm6eCrOVPTTWMUrCqJjh+fjCPlH
IKa7tkLGD3/SLm7n3iuH/u1SJ3tnuskclPVnB9oo8ZOX2qT6/jpZJMesLRSh
ckKPJvnzO05RvEGs0tWoEYQM51cfdkGv2LqrbRtdk+dd+qWLeIuJmln2ZfL5
VqiUimNua2Ci5NC9Rg1ISrUiXnAVYToyl2iG65W3umh6KpM0NyW1XvPkNwiB
wSkCUEDGDf8VIq3Xi8FU8+jG5KgfPcaxHCEfOnQrWVMonS/VN8ayHWK47IDF
/YsHk5by2DBWgL4RbiMzdUyMMk6TWJibTjMu4S9vG2TbGKIUFcw2785qmfwg
Hyw8J3qZWS+1kEVeBn9Mh/Z9IyKEjtWWHA+h/qRPbfLcBzrTLDG53noBxYZ3
TmpwREjxxSMHPri6116ikXykNuzX5TwSI6V9q/xcM7HcF43kYg1t0Enoq4ii
X0ZVT0A/fCsbV7GjYsX+Td7Oq7rFIRVSrHEyowQB1nX0x/ohROtCwBiFLyt7
9Mfqt1Daq0twM3nwih9gMN9rrlmY+GYKRXppcLurX2TubRllC9/xozBn7hFr
YRzXw+dBKh0eK7CzNV7PjuZ0ngYKpo4WZT61lMPKsEPXYOYfzGxMWaYgcBm2
BQeLEXsX8Z3QxKRmIF4E6kdVV9piv8nSi51FExdm2N+kmynhlpgEoQ7BClzc
lg4l5igI1GwD4fXYOcxzjXBqGua+pE/CmqE4Ceomb6oD/WzChjztkuWFBZ68
GivF0ce4ARWDb1hk+T/+fhl6zL08v9EaL/wjv3I7RPJTRwOLgWh8CnyYWj8n
daLHScU9LVtqOznXMinuZJBGXbFEgFnSkC/OSWdJW8PDnN03zkrEs/gFNd03
ZpRKoY9m9DgrpoPFSYdQHaNWj2v2dEdDjJHa7w46hxtR6U0sbT6AsIRTcs3T
uROBBb39fqU/bnN5fFBoR6MtLMmEJ5+8pEvPJcQ0SEIgI200GHonpjt3oEQF
LJSZZgDQe3o/YchFonIn2UGLYOU8PY7ComIhR6QyynTibszkD37nuQ/8aCog
8kMK147x+TuCkn8wpc0CibVKdTUdB0K3JCusmeFPP0HNo8G82Hg055dYM63w
ffvK5SUiQTaQU1kaO7gHoOOZQnCeAfrSeRWl/gybfH/uo+JnxkMAR0aYyd/8
DQkzEd1yDxejsO3cKC9E2aqldpvVGrugr32lEgQ0MaGGivJ1NaFDRSEEIoUQ
RXv8lPMU4G3xErSpknH1nx5sqrrOZe5r7+OR8FqeThXel2CF8jWfm33GpIcz
eEKYxT9ARN1oUJJfNhCEOiPuW29ZuPpxbGOEqkzetfg9dIb3Oih3tbqTjldL
Hn3rs53rDsTlwOmmXgivwjAWfF1kKYSpcyLAcZRGAd/D8srWytLzuyCJPVHO
AOJDAClptHxMYnyyfrtE7yHu+5MhMFgxebwXfq04n0EEoTZCBtDncHqhPYap
gQVbzgb3df6ZrtB/fAJSjp2wbHI5SWAHUeR7DY9aJv+iHufUQQbd17B11rlC
oeUeglXXhCFbWhPWOzFFQ6bmPQjYQO1RW95Y/vTQgjg3Q4P1lfxUoVNIL7cD
QI4nAkoZGytWttELuaXH9rMgDXrFv0lsjxisy07FQaeNSKLqY0Yav2YWFJA0
MLZ/ZFxkiOuyLcMm2yHSm/hsZ62cuqeFdAPJDPzxDIVg3MT343OvbH8TCgR4
hzimJxYYG7Rf/iAtiYRf5o5SVOeVaJQC1OBIsZ8k18ZPXsW0My7UjFrC0TWy
cvtwzzOTWw8fomij4geUev24zEVeIG23/AquXIdaQX7+hfl/ngMXw1Sv1Twf
dsudhzt912NDXb0I9S+miWGmiuiCB3yYhUWyFLp9c3NYKa8PpW5v1vsQndK/
V+8gsTUfGQhreXYuARlWATpD3jX9ZBnkL0hTFQB8hRLCHfphtv3CdPfchbRj
7W4dfbZMZKh9cAFyAFj1RU0bLAt6MV/AkT/ERbiVP/Gi78E3grZWi7OcbgTE
0cZDrx6Xi0/RbB0Fa071mTt3dnpIsOiPkJIQ4OdSF3pdDz2zTzG30KEhY5b9
N6s8TZXjTkxXutGeBlbnNOp//45HQN2vihqnVZ4oZHWflTZW9KC90ryalrcv
dyj4Blx+jqYEoQSjijn1nZJizc98vkqSzFeSeQsmD9jW2poxVCBOz746B0Vw
EgGWOJKE/GMfXeX7iaOBbTFmNE49u23rJ86RyyqkYlpPRWxQyxSuyG7Nl+az
2P2GOBoVOlLEP5uMIb/gVuoNUf3bmqi10Mt+CTsMj55pSZtCKTKJX3PPXQhj
kYdc/mYO9bSOlycHhKT8JsCib/WYmbwAyYufmGW+mvUdEM00cQ6JPzhFtiFH
scQEvVxERNdAOPPlvrXsCJPkDvTHn5297b3rvXACEqJ6AoRLBJLeVSvw16oQ
jQH7btO0Fn0sYIb4D44HwcfsFO6PMDaiSBc9OXIozi8fRqppikZE4NrorQMq
Rp7RX29mybz17gXIk7z6qXHkXM3nWPoTg5+FWR9viEaSBeIb7ShPe/BrN3LM
9T8ZYV4isz3LM/KC0OsAlm5bPgeMqD11NhsNzjqD0tug/Jb5teXYfwGHRDOe
17MI1y/1niQmAVC0c3U0Mc9mZHXYkjJewZ5a69jYWBssrGLPzx6RHRVxsJIZ
dhVZcwrKlZYpbBB1yZBKdBSjGEWY/D871Ug+A//L+nK6VuJvYX8wp6UPSaZ/
buycm3YcY44G652PWjUpkkyE+/yQSYxo9qq40t3DmMRvtsS6C8W7yp/1Wb5S
VouQMonEiNOSMNRzsVPdQZyLFXJ7Mp4Hf/QUejQ1NUJCxW6GsBsLGkU6+bXZ
KZWoyrHpDDFQByPZNWIbRXqDGShN/N16vCZx6cLM/kiHqJcaC2NzQG1z+9Y0
Uf7iRberl+SeMEUnuzazy/60vjbFk0rA20u/y7p+Pd5E1xWTXn/U6Q2XhTxN
PktLCuBmYdVvRteR9wnQxcEBghm94qGEL+VYhRukr8uqXjJQ3U2+5Vspmtmw
e1VFoUMVWnmc0W8u1pFvNz10xSy5I7YgbxblVv85mbud40SFaXMXNwN+WO/1
w5gHMN2h/0im/tG4ZA9GlW6443MaSQ/L4+ZIDSfwgdcsF1lJhm8yVd04dcb7
xHknjll8YmpMXbMUXgcVGxnq7cHV+F9wfC0nh3Uh2/02tmjLa7/Tta8f0g1f
JPdXEqMH50IawCAUc+1gMyEhV/5+Of8bFCCEUapQUIjw4hxQ3D+LsFM88OJd
YBLRjwlju99Yzw002z8uniyxFsrzGT3xn8SFY2zH7DC0J0leaXy2YiORgYv1
/NU6iDGLF+Oq1iilkk5p2J+XLFlE71tudAoeZWbDHQKrwEhxymNjOlWa9xSr
HyooLebFVkU76LAraprUz9b8Vf1D8tSZk0chpni5DMYfuT5Eju8QFpf5v5wj
/6OWxONt5lxTpbhLhhfRrMhSK1Z5AawiDOyvqBRoBzLyGz66V462xneDY4of
q0gqyBhPn6q4F+AmRv/NLjSXdSfGz2vg7AQLF66+jAFF3fIuKhr5jt6Rb+FC
eC6t1DtRwy2pfVkQ+F3vTC092G35/4PIX3mq6emYcfFDJsMhr17G4/hbjI2T
sORuk3o2j9ShHYvZeBEzWJyW6WtbyMt7G+rL+547tfrM8entl5imrQP1hqXm
1By8cmnkSHU01sOXMH4anmfgQCoPvE77H65qIJO/1vtrAgWfLA3puu8XFu0O
beQ5repC2uDy22z+LQguCVuu8/NKlNncBxidJ6f4LSAy8/8MkPmTfO0QKTX0
YOgNy72M9Ws5Z0diqgp9G9WtS1Z8VwMJMoDBdhJZkv2R0s4Omabvc5FdYRFL
QwnlCf1FP24XMzrTa3m61Wav1pCBgePS2AN8r9ZqdwbS41FDVxi0F/HINZiI
ppRnn1M/sX/WETBdXgH8rAqEWRfoIQRMLyFPFiSXW25xBjKtS9VGsIwS+rjw
XMp4Z7eQXBGO46PzwSFDvOIrbYUA+89lLkvVsRcdCBA81T6JDa65z0386I7B
gr9iVyZsSklABprzTlesQ8fRz8sBrvFs15JQu4Tsttl04TB+c3qdzlaPr5gl
owjPzGRWQtRfMyhUINiJjSM8vs5VDqzW6cccJB9YajcfxqhZHXIrIln7RBXK
QESlZAyFFBhV5EGKSCx5Q+KKhWlLAV1mxwuProCsWFYtxrzvKmyMw9iyMjzC
+eYifZNxQE20DwfvBdMWfm3W3u8gE2DUeAoovILa5/YAG50mBI3uOlYrp27W
cVR6hSFBQD6o5KnW7jKmOvDrWgGWwf1vEGQfiE1VdaHurVRyKNPNLQXfNxCn
Dehexik3yZi6/B8fBkGPSi2Z5Cyp0dOqaiW61HdLpTzcEtmUJRy5J7e4aC9S
nh8/Zf6x+Nw6HSLC2cNQ/4uCJIkmocXJGdMcsDmo9gxleOqp++Py/Y1T9ro/
Lv/le7S258F+EE+SopNlpTt9DhdIFtgJhxa4o6UGVRQB4S999ES1gaJPyBjb
su40otKYEUuGIQxRY8dhli/ksCTFcgNmVI7m2Gz5d7RqWYqS1jD+M6ypK238
9Qtx0LMGOGlfhlOGeWzPdCqZytMyu5VQMgfghZgrLmmO57RcevoCHlFkyZkK
cYxwj3afx8H3lcSq1+kRn3u4ohSLcH2Oy2Qg3ytlF2EsvoPFluk1bCX3InRK
M7AbIjM4vHA/mjATSTTMCzS/iz78DgJMTg+i7LoJpjBJ6dkKENH037aKfV8l
CogKGt4kxh4KuzAxuPJUy6xtp/rjoNzbm0fRutEHhlwYsHG5QzlPfS+zCv3Y
Tg+gOY4mXYxwXG0DlyPuTf+zqfT7RuluuHb5y0xFQpJwyJmBPSGvqiEN5j+E
jW3VZmpEe39L4Ki9+Fq2MMHpotIHiIjfwXAhNOy7cOgAP+zNXboc8RNEN5lD
XuFEjmyk7/ZgLadx355L1OFFOKtSO0IORhDVBrI9Mfvs4nSbclDjprUIfdfY
l2cXyvODr7To1bHAsY1KP3j92K6Q+jWmN3hwJiZ+bAyw9eH7MqAlMj9cHPly
OPSE9mW9SyGvm9e774Z59SoNGPp9ESXoTfz30TG4oc3AhQumqK/XJrRHRn97
2BgSzlZBx0aD951F7IP/cfF8hap3K5DRw3kMu/p6J/jAArtgv5D4h/gW/4/f
7HVPww2nl9qsArwx+QrmvIs8JfURKtl7ePm5J4bcAHd0TJn1BfvtOs0gINf+
LecaLaNEZMZ0L7LbC+1sS72WJpYGGcyGmZZ+LHU93YHqNvx34XmFm7tu3PA+
62liJRDFtDU/g+APw/3R0le9/7SNDw/w0+1+zA03HLsK6SjOFsu1x66q/rAe
zv56Mksgccv9UVJ6BackPwwhkffCB9jNCNaPsiRbVQk+exWZ8ghKgq3kMmFS
/4jiHmt1SS+eQOTt/vyUqdswHN52wd8Q+D8jeZfoSAqylhgGOOiPcHYHjlZv
ksr7wcWrQHQhMTYStt9lDZKbc7Ecgdb/Pfx2L7VU5gJmhPai83ydzu133WyZ
qV++6YjPOCpDw9J8NoFD23Q1rvniIPb9tFZEOPA8mgQCuBMDLvNgZYiF5fSk
QZN5aIo9tlO/B3eUqwV7fRWNejyNX0/ZX40Nlzd1O7E/OYGexzyhhvMSe1id
AgLPm5Xat/msBj7mqDzlCSiwpBEloASW5HLzbabMuI1VzC4HqgB1NWzD1Fkj
HcIx653zf11FgrruCWcDLTSvU5ST9w3P3WZ9K3g3BjDGEmJQrxmwjWaSkYGp
pfag2MGIylfVVcjuoawo8umOy1WrG2FicqyB38FPaIXBGYBqTFQQStgaj4Ta
yq280j/JXRJWKmvG9GRrur/cyRvIZd7XblkFu38ItGQNhC15zDcqav90WGj4
haaYAK2LQK3uNGpxUvSqyEfGbftg/0SUc4zXBqy29eQhBJ+vAE7jjY+EsSy2
UrqUtICTOkOAEfdABQHba3sYimKk9RB4OFalMk0FuvvZqEkrGq74XbLFuR2d
7k28zlXMDjzVX98c4PC5bMikpybff7OLwbxDaXDWogfF58y/ecmL1qBhusc9
xCsMdt8VO99x7RbfZnIY0LaqPrvLBeBETqlzb0+iCDJQ3+Qq/KPNEnaSctm7
A2rHO9WYcGDhkRXqZ7YOgwvMUFkJiH3Ig8PZilj7xD99Qe+dJheARxkIs/Gv
Vf263JNT7FVXAG+reI1oVid75H+BkiJvEls/tVv422Q0c9ihRfhMQvTYOKJt
sPAE1VYX5RynfAifHxtTyhcFES+lUeL3xdVL9zCOwaN4gS9H4Yhsy0PfbXUt
fQviMUIvnNHYmxrvhuNPrpC5bYXWm6zeDNaYWpISOQzc7BrH7T3clLJjzZbB
zWtjGZHPKo4VgevubklOIdG2sTjsUhFMXJnB8+xU7jyhpQQilxudbBCiJZYy
wPy6UI7JvOfF9fBYqswLzI5NtyTXudVV5Xq5aXh+l46Tfi8WwKyDcY0nDnCj
1AA8U6WZiDvp4+P5Y91dEtq2NZCMT8MWnnSkTKTmIlY/hLpdw+OgeKIBWLMn
miVtfB6Yr1FgiIlGVUGRh0wJYUMQPhEMF5eTD9NJoTKC1Y1p+yo+McT3Ba8+
kEAwPdQTSPZN4jdHDxuLTBAzKmBmMko4Rfqx2+gNRzOmti+ZiCW6kbL20wyo
EXNpXggYrbifmclAfADTWXRpDTJPykP+XP3uIX1jrAd4PsdxS+JRSAvQiWB5
+tvyL5oBpDYzY1CQEemzdQlglME8wpmkP18qMT0GuOfn2EbKnB/CMScK1FvF
yIpslvn0kmgsMRpnkVVsfAtc/9jnKFJrBmHt1LYhhdOzfaXlqd9XZLw+gNrx
koMjtQfUl45iQ+vohU62QcznWn+kOeqZd9RdCrImUohJkDIl7I/2JzvmteC1
SPVQ4m3/LKcUsTVtlwGjaLElGVFVVpGF5CXyyr38h7eePyXrgnPjWXyMmpMF
1jEJCqJTy0ZMzRYMi19LR422mfmfKmvVIJH2je8mrxc8L38S4jLyypAz9xkR
Dl7KDVHvbHtOiKChHCm4zpbemu1DJKaIKZHqGFX4lp3pils8Al6UVHJkKeG2
rdrmLvAniGwEi1quTabgGyhA0ecJLmaj9r5t+OjqQiygoUqWbMp3qC5ek3Vk
fGI60P+1ytdplfnQ+aco7DFv8ZQXJLh+v9/cYUSnhl+rDemgCI6eoSkE2pOf
g6Rv1jCQFzR/Ds15a7AZPafm7P31tvrRgR7FbWs1ZNoel9lBmLM7c/ovI5Zh
QyhcSOiQdr+v9GubgjC/rMWqYkHRGJ/I+n+83b1YLtViLNWK6xN9HgchNhKF
Wa/MAW8IuwI0liZzbegJTm5D+T7eyf2WBtfj+BnVocl4rFn6OT1JHR2iMNFS
MwneRP4M0iTqW80G+yVb2OFsTiuhK6IM4jDshaMY7QUJ+etQqId6lHc2Oxny
Yj/VQl5M6U6q/3Kag4aqjlSXJ2utElVDK9Ob3AsHHfBld9S/JqraKStkzLKt
85TfOCJ0aYZ35vAU8DqVlEJrG1ClRxAy18HaQbIpRmgX1ent0q3iBryaygGg
xiKWxpiSsnfc9c3ndHNuIOco4f3/e9pGsUIoo9K00ygs3LAarPovdDdeBnFz
+IP/RQaFDSGxhbPyILl7ElCdOLq6wW0hz/gCFdypft6iYdc/XxUDWeIdNu3M
3tF2HP228w2YeppN+jqTNUWhKIWLQk3OnOX75IQjo2PGYvg+8XJ03Nwiho6I
T8RVIR741Ie7hT1azSRbxbdu05OP16m7C3VzAIydhZof08IT5C2J5nodVNDl
7qTREaN2np2jgVSzvOBuS+8uLTtcjGH2NchXzqGrHngbMguXRTSemMZs2afa
Dm+DXlPi427zPaq/CW7PPN/ZGGrkYhYGEbadRwd+sO12PXIo/hsiigL+WObJ
/nAm4OltotCZyH5JMSMB/NT2rD6Lup4ojFagibo0nOKHg00cfcFIr1Fz0SVi
i0HQjjZVn9dBdNCGmd7Azur3gCZNH3JqbVGZOV54wgEaprVNqandshQQN5qe
ugd0io1XbqVOSsSfyNTodrVY5CWrcG0E8221CN7Vdg9X8JWRI7IdnbeFH4X1
u5c/ZW+XAYxtKwoYDrfaxzBBtq0IDjjtCIpoiCRIvtexz+553Ye/l7+UzhdY
1xOedxYZJvJWPC1tKLinePfoT64uZm8CzHqdluCV2op8PdnRGEjmVv192U17
SHf5vZqGlFahYxrxmsbDJuLMnZWML9KpMNjoaHNC5B8NoWB1D/FwkRV7qaZ9
ccHlnaCxMut8rJtQ6gLUOv+01VnuWe/YXJNatx3t3W2rdffHAkQIdwgONOTg
x3KkxZZabcwUZIMkzbE/dMjA1kUTD46ZdvE7cbuwzj+/ebPK/96RAey2A3kf
cWaR5VVR9BybrxgkAKg8rXSa20vnFsdCojqmO+iFmV9tnmMu70KQ6/dDMGpX
ojyfSNvObTv9uFeqR4ER/r+iqYeQIpPUzpz/kKalnhb0e/ZHryUtWmtLYoYF
T6R0DR3oD1MilzooBqdUif/P1pWQHoYORRsb8RNK77lDhk7y4KHWF0fdkv01
XNd23qG9BcAv8iqReNyXcpRer5pZ7x9535jlSK6X9gm4KxA8Rdk9njLaJa4I
5Qlryq2pEBKczcCAGLFNQyoIvYzqYQKaNhr1CyzQw9BTVzWTDeSOVJoGKJgf
ao5oEcKlNMUBvZ6z6Q+zM/g288405gO0lJLgz6cgWfvBLtzm/ZmPFAh7S5bI
IxXTuUsXMNM0olccwOortrZ6xRCjjkRH6UT0yigTdx6yRqEbsr0slS8GfFYX
MO3nPLPEYGoUZxo2/43FBjZW7uWU3RrUGduiVkaKKrRuRC6MrnkZ6zgx5G6P
m8z9vpSsZOukO17DZRI2vw8HIHYqhtr1l8dvzaPJeBxuc+GFVSO5gGMrjpuF
1r/wH3PhVXpcI+V2hD3vdVmjiQEd7mBl59+fEQbEUdB0ofn2H8Y2dMz9Y04v
e6mD7U+fRWKQ5AJkD/DVas/Z9kpFNqoeUkwPjPYOFeecqk6hTnP6PeM5dg3K
osnEIRupJGM/rkdT63wCuOULwV845PxQtbooEr6dOkgHh3UvE/cGR/h1ceLN
OIq4CkqQK4dggs8SmWL9Oc5zEaf3PzsE8aVSJtBDSeHHmNTWeC1fZBMeU1DJ
Gw3swGlClzRDvk2I39AnjmoKeZaGUgL8ATkXV57La30DBINKlISk0ZYct7PU
FUMsViCFbgr0kQJMaxmfQVSBdIKrRonHhA8NDV8COQcMO0keo6kvK0ML1CyW
QX9KsMimQ6/uXX2gwQIrid4T8kqPD53FAb/uzB7IpL2yu3L/ONS8w/32dUbb
HLKUE+BbFH7XI9xyc6OMoav7aSXGi998yMsY4csb+vETOWxdPzzpujVPnChV
0hAP4HZP6c3iVd0L5rV8tpQZ9vm42+4FH9NZIR9ZYifhnJO2Ig/3bgQjRDfn
wOugJAIz9E8qMFJYhRc6vtT+Xx40jVOctdReAM8EIZ8eAidB3+CInZa8KZHm
1LQk4OEEQFAM4gE2Moyvjjm21q9eVnTx/zeNzW6loXXzADZEdmfwMhqo2AGz
bqByKax6ppkozV9ys1JimXUKqr6YDGZu1G7p+faUBjSvyoh8urobK4KwRqaa
yHxnBE2AKjVCj+lRxWKMzoqJtPRUvSwdTz3YDLQsoqGQ4HOxbOrVs4aivMcv
/dhJazJaBVPRyJxwtz9hzWD3SqHPQWH96MV34QjTZnOxdougQgPKPjs1TeQx
L1N+CrGMLAGw3MdMXfS9zJdwHUNoy5Nqc1kApMLP6TiFdfGGIPA/tDlSNvLA
zkgjFoEa5f9zedHgGU840ojae1jtJMkwQ+G6vMzPLDsDLy4ZhAOG/mbKqhmT
drDiq2j6G5oor/yRE/oNyxzPRc7HbZFj9I1TYoCccF+72sIa7aQLLhIqdXee
ds/YKZxezIrHEpGCmZMxRO7nC/UwbrqsblpBvMqesZFAjCudu2xR+l9tW3J4
i8sBk6HiXsmASimM6Wiv781hB+figCpdXuVr6MiIwLw0V9xHOhS2/y/MDtGt
N/fMop7FE8uL9FDFqNiNhrelfwW22sdRBk6M6bQrH/k+Oh30vhAlYlR/VAoK
e1pooJzxIaM0FtsrP1uW27TVDQJByNTDqTmlBFHuI1Vdvj+Xw5B3mEp65CuR
iinfbGPkep81Ta0pAXJEm7k7Myhmhr9roEaVxh4Op8030DOLz18k7q/h5uqH
RcEzGl/Et76w5ngjNV495ReFqQ9MkGt1NGaTHvrBT7XT8EdrCPsTP7QjxncP
snPJtITHZH34/GY5kjlGf7yoLhxGQSrx6UqvasKQj24a9eb9eDtTQHODlubO
52h9maBriGWniN7waWRI5amo/HmrdbWRRp0Bmg+QlH0NCS/zPwsHxPCMTwJv
U9BvmsPclaXIcDFtdS85QDw5Bs4u8qEFRLTu6GwOkFW/JyW8ivRnGN6dQs2F
HMZBF6eScfLOtg9jtmaZy5W1omhGTMbPjV+Jowwv+EQQIJgi8gSgZfFYM4Z5
WVUB27Heio3GzO8x5lOu3jflaxDdDh7xzxofr1ixv/h5/dgH4ihdBroE39dw
+FFXRg/PXROEBqxMHyBOhmc3bPFw6+uiSZoSBfZsOtmW0TlfWulQuCy8K0Ji
ZLx8qQqPnW/p1LEND8u90M6/DfdVmzFXWqbP931wLsbESaq59/R6t1tqDC1V
bwMBeoet6DIIzQl94yXtdFHEk7KGgXffDRwdtRpT1+IlByOjxkREOk6O/aCW
YQ+XckF2lgnS9fClgo9bGx44nHw9iaIMDp3rB+6iNinerfFxRnSqk31wqc36
1CxNCx2ct4RI5xWaR64d2ktRfXyCcCZ0hcx4Otc6KZRjqk6RMOBaUgtJsF3u
EnhGkXXdH9pt4x2Pqr07OmzlE3AELpNtmee+I0bmIBs2mb5Tn4B/LMq2ICON
gSwcimF4D5SN9CAJJDncSFpucRku/WkW5CnNNW8UPJ8bswyfiEy7oCE68gD2
DoKkGHxTpaBgLaZESGwaXSc3UYeapLOe+YHU459ezuTBvpGm7hLDjihKs418
xjcq1z9bvRPOE/evvpls930qn4zeyj1N7ORc856J/geL6onnBBj1S4TLZUsT
6DlcqtlnV9ajnfZkgAqw5/nt0IiSTHsF4MSNo2VTc0e7JdwqJEW0chg34/ki
ilzEI7gACGewjwXYaUwaSMmEFcewnUfHpzQIY43TRoVasra7jul+hO/wFH1i
xYZDSuohetfnROdyDm9K/Zvdk01zfcot2J/E6dgXiTh7LWaOjP1vzyuB6vCd
AzVDNwQqnhtraxef2jiUhmA0Souan4bhJQAzqSASAvlKKW83Y9Ac9gLyLF7m
a2undAm8mmpPNuEeSNRx82uRfFANlcdBy3fUtfbEkRm6D6sdRJaG9/cmA//S
BcKmxjwS/kMy0yclyCpy/95A6AGBeduFuJndRUacrWCvCwYpa2G0qmSx3Kjs
esddZnkc35AbGTQRv/DpPumc//CoxWJkma3u/K0T0SCNffBY7/QcxhC+wNqu
ivQi4+SNyzWgMS2o6QlF4oLlhRm8nGhuQVKqr4JpN2tobNznmRwcOUZjxrO/
k0kby7qhpHpfcrjl4jBJvD9UfFnFIArFpwFf2vwYJHif97BxONMF/JpJQcRu
/UhNS6w7b80bk7jiuO1i4v/afswPIYcq8j60gRi70lv8p0SWZRcphMMlby37
Aji5vvCapGhb59yEcmpJxc8522uP2obtNzW+5BJV5mPEjVGUfBbDcXTdtwSP
Dv15RuSFP8RXZKUxdraguDG3ka9QHWMjBdwHHwTLqaqZYmLrWosWzkNzPmbE
DUN7KcMNJNjZWBfWNf3cJUFa3e9EZVjjZF5P7sr0HwHijgO0p1Ydo41eGEGO
NT1ffHVE4szTSl7n8M/lrQeILgdyYDsYcJvJ+KZbnTba0a287Ema9IxW8uiF
tY63eA8vt4kV/namGxyDFYzpcV77TceSermk+143i58e8lpMzUjG4NKKLCYq
C75R4yNxBSYb3f/onBAxXDH/k6IDQH2CO5EeNOKLz8QtspCMqzP+4t0kYJoN
eDPT46owKJxTAdczGlpAE3GlofxyCL09FgzypYhUDV5p0rinEu0gyIXzlY+J
uvZFn98PwcnOhTvHo+Vd5INBpapNhiyEdFS2ayLhEDYwqUVecqo5gjFSzrVX
ETSw6kJJvF2cDKBUv4yLwm5AMHcWhesKX1L4YrApW0jnQzSjfxf7np5JJJfL
Vvbs5k4lu3Ox3YdcbkPBZh9s4bd/eGGHElD7m7QfJjZ17C6CNUuaRp94ewyw
GRQfFmyHRww3UgAIi7bEb16/C+PK7lCm9jk3ilDdQ02dyml2EZfiJPhD9Yx5
EPZCtv/HfNG6l/x6Ogm/FWtfXb47GzKJqjyZeacxeTkZhK5Dm1PRVsBDtMEK
roTAVcV/wsgLSyck7GiqKn5bX6SyPMySVrLo/nND5uAK8GUwRe3v1KbuSBlL
MbxuD8wEz/L7mc+zYcybRk6W8m/KxiTXwMyLY8dMexmXUJG17TOrbMBHnCjK
6XLQyFeWInEQ/PVQHwiO/Apq+IulYajdLyVuPU+Ed0kic1gW/5VUxh5+Od4q
vN9zzD3TNWsJIlh9kxQaN3M70OLRsxW1+0oC4uu2N7oXmU0ct0JOHOYgxzIX
87gEo4qzL0sWA9MbX6wVCG1dPEZL/0w5W5pabmmtV5mWo7Y8D2NlSMgEJpSD
/ogbq3lrbBj0s45BihJsC2QrQdX6MYGu3OUzQXeYgekz2mLe0ybOIAEvZzkr
WQTQbbfXQHRky1vzXPfXa5YhOB5cKPMzU/oUpPeCi6XP2xe3Wrc3RHm341nj
7/SaUMhwjlczg1UDwAGrVdCqaRx1pcxuANw/vA6mXXQrJOWVvlvkoa6nyAAG
Is0yPaZcPvPDdaCFuaowRKguS3gOJdiB6DE2449ZfSP52RGPAGZLOHB2rxv+
zWeCY9FKqT84Kb+nCQio91Y+Fn3R7OJk2P0Q1U35g08gClqDyTXFJqmiHSKh
McusmtcUoxYmQBm6mFCSMSAiy2robbBjMJZpuB5X49cLcrNXIjwHRuaoPIqC
mS8Vi829DtLzdjaeZuA8RTb33JcJXI64vz1d8jEB7h+BEe8fMyLSEkfFoLMN
jGWZu2+QUzgXkv08Jo4OsQ3g70gVoNQmByb642CjbdR+P8fUnOe151o2eopJ
lmCFsdT2Gl7MT+K+39YWe1tuH+UCWA0YeaJMAfr7nqqRWePK79ZgJN38U2mi
14SzE8GTz+mGNM/gTGHoQcg//wuQ2lYXGq6z8uNK06GkryzRxMm/mQScWIuH
7bycuU5spuK74A9SKkqn+s9h5VrCQ3cL6jb39KsraJ9WEJZS8O9D2h9InYkp
RnjKZo0BpXzU4V+bF8s0gjXVjJOw69YMFpXCiit1tN83jYN+sQVfm93Spl0C
RZxxiMPaNCAhtvNI8SqsPUb7qNC3ZRyYNckfW9tScdYF2eHoK56byRkze+4E
1olcJFc4FStQGKlmdZWi6OnhdTH/8MbyB/X/lJ/qnERBHXCSkI8oHVDT7BSB
F20BAIEhaN4bTY1HADo0s9OqIdYJEnMCZdCHCb1L3AmEWCDtzwk7dDQn2V1H
TBLiB83IS8uNQaVfuULG4Wvki8W85HxrTbbrW7LyTU3KDtVkBllzMk/gYWg5
BlcqmGmKtv8CM84BJQJcmzYMBVzv80d0Xmvt8xsuGrjh222mexjMYSToB5/B
5VLEIfv5QUWA0fFO0Di1TATLAi2P2ZJOCwbJn46MdNp6/sRAquwc1MFTSKx8
5n5yO6sBaETmDPbhGLKZOhzUN/dZCw0UfPpB3Qgr9t7GHNIpid/aOvZUH0rd
8iGSrGwVRTChPXYSfxsGvYadKz8taEPgqJWPk8QCEA4EupmJhzS3x6EpVT3q
NVVguM6r+oht1qHdoSqk4KYlUYoJnOlZ5lBRzrbosQ0wKn1diQwy3QN/J5bp
BqQnItfjvH29vfbZKeyEYq3v75Q7mRSd+zeDWthJridPGQHBpvrlhv0JjKqY
w1cujqn32c09gSFXTzVADOHMvvkm1itbqjOpiIld7/kzaBH1te3KWwfxBXcf
uDt5z5+v/oI8yVpbF4zPcBe/wUkOezOiy1UOg1FsMI7cTpRjcgRFUZscTWYt
jV9yG0MyOsZsP696dK3j8nxrEPa9NHPhZBKEpG6sYhycOvmmh1pJlS7PViEs
slDaW5vz6Lw+o/ARdunoknZKwuF4U2YG5R4HZi77ToK7ZnkzrFefc+QSWYw9
QzVK7CLUxJBLpGq9SWkq5uAwSkyc+joANZCNq46Svd51gjMWZi4HoQnYhWpB
XWFsYhin9it4jEzdIuiSOMFpAdeXbtch2So52DJA8cwdByEvHOckHrisCh6O
F/fdv3cbB+BUkuZaBmggrjry4hE9IrpAHCNwWIR7Tzlz1dlQVXudR+C6GWRh
7ulLR83/I0XHwHSlxalb8He68DjtbdqIBiEbbmAhJdrW7FUfv6hd6YNtHtUO
K+N41cXhYL7O71/qvrcd0GCHJ3Y1y1hd1yWrJ58nrEmewDDFa5X4shjUu0t0
RvVQT6KybUbrlmkjff6YIEE604AyidYiszRTuIn6knoe3LKANY7V0YLHs39y
Xx6FuO8g2ACMjtACOEtraIyh9NQbVizswW8mSwSjJnKwMmtWN/m+gy3dxVVj
UGrg15sHFR7trYmQ0VVv9fLJc45ft5/wLh00ImQ5l+B9v00wz794/6yof/Oc
wwVKBAx2nddKowFBmCMhdu8ZGmpfQgzRbmj4uLw8nyVo6C5b1YfLLUaEbzRt
n9U2r8lQ6RSy++yBgATzh2AgZVGIvVNGNGbSKcQHT3HCVd/lrU26GNo/ZB3+
vrhWMf3+1YDiZPbdMkBV/gnlp8o4nUv4RAoTxVuXwVlWB4LNK69JY2PvFe8Q
eYYTxZEDynIDSt74RfP4jER/L90dHb5d7L4ZHHNwKgINYmczkUMENY4lKwXm
goUV9RMM8Z4Hx1XZ/OrTXDPcyTatt+q3eEhQZ/0aajm9sM6P07WPojDduK2+
onNNWfMaqILKoPsAyGH/18+vrDjFp4Ukkoz2KZc5c6iicuG0CvyQBAIqZQBw
6toRZvYKqSe2S0P+BVAIjHBz96UkaQkRQUbfJ96+E56NelV1rJ7xJuQQLvrH
bkKleV86oVRWxmC4PULn5FxZEwGXURYo+ZBsu/Jf+FJHnxWXDlUDzvJEppTw
Fna0L3DS98YCaBNnIzYZeNcZF1+6jDVgyAaOV6UwxIoOGg5vDTxzafsLqtut
cMtmd1F+woCBxczVhdkkJwp/Pxq3FPQqyVag75kwJDXKIwP8QumYqWRZSA1g
CzsG5WpB2n8GALeIVPDHjlzkiPH+UY9NuwqEmc+VyqFFz0E+eBU5uHq84U27
VRZbOZXbruYywLAiVUEztAcVMkJwSiWbtBDA27bIW3yunsWX9OJomrSFvkNj
wFJhzR527ZkcQBrtKIq1+tsiH0U3SClxKfA2jDjkssBYZuBOdqzY8DUMiVT0
uX/874qkzVIRrx4ht8lwbEi7PWcAEmUUIRYnkkMg2zA/KVwoVIITUntGw8zu
GuXHyl7WRggM1etDJFbCtQuKRX45xzSt2/n/4WQrI9XblFXD7OxWJHvP/Rs1
GSCcEjn4/d0eXvkTKuVrVoO0ta0XUTTzT0s0eXQICdD6ucx6tE/3R2iZGzBX
UPL1AtdZHUE5fEMg/RZ7ciDkHNP6d36GPsx/635X9ulHQvLOC8Z4RZm1cN0k
wbyM0rs02CGaIYq0No+zI/JNaiZawZoqgt51VGXWovj/ZRVLy7e4b/u3/e9m
R5AO1PAtSgSzKqrlZfQkzw/vXeqUEJAxHhk2fNzThWs/V14phnGscewVeDt0
WLYUse7I0Zaand3XDODJ54N3qxv5Y2kQp+2AV+xVfve0Wevi8lPXRDiL4UdY
1p6E0SWXAuWyM0i6Fkj0VqqHDp5F6ukzp/ArvIlgSTqj8LOoOoMrlaJIPtWb
n/p5+jfFhYF+0yEPT5PfrbyHNwvu+lG8+6tVnVQ4ggF3MaomC14WA7UeaycK
KNbxHBv/AMNfQGqcPlL+VGuuVazVDYUG6ZvsnfLuTX/BXBRCYus0edZCeatp
Zsk1fFNdWAGz+PPCsTjsH8I8l9ZSOc7iUBXhEjqrarDl+THc0LWCJ9VhJ/BI
zuZPhIXCDO1Sanhx9QZnELwXQ5+68yN3agSd57nWSkeiAKwW6vLDvjQIrk2U
6V8rHC8ME1cOQZ3+SiGBvqlYoVNleaKND59rMuWmSRfhJ5E9IvJPI2NmmZy0
cT5LmEL8RzG7HnwAHGqhnYmQt6aHr+ACll3W/tyB2Sci5DozpwiBtdlmVqiR
+qMIuc4Pml/cxgO3zY9Y9FhnU6l/bVgDa7I7oc99K4Pk7dr9xt4YoJi6SiTX
PJ26Q8y3E/q3wchecVAVpqolQIoNBchshooF8w8UOKh9PxxMiMPBi1bpkZ98
o+VRDj4E8ABg0WwnHbo7tHEWNSwL4AgvnS4BPDVWZjLOqSkl5jZPwpZ9xdmQ
V/nw6M+sW7r0lUMqzCWRWcu1YSuLquXkXv7ZRbF9KrdXNOLske2RBLs53ugB
airvAo43yDuAXHxKhEiJPXfe4k9x3r7K4B2mo4ZXFhS1HQLX2jkhj4EdR/Ii
V/cvHlzxbwrW5Bdm0czKKENm5sy/hMMdW725nN+2FIedAVp2qkFzZ4maHtJB
dM4oTWVeU5SMSdWMJ3YhRN+hDhgFU8JDYfnOCzbWIL+gwGmkxbQTevXHIraN
E5nliqzCbct9BbAu03c/3CNvGTh12o7h5Xc7IgZ7WYNLtEnyxPPtyge6m6kg
3xPE18d6EOk+nR0R/7Ba5FwyIACBX9BAyt0O377hrCfmG2JDBSqKL5u3xdLE
t6uBZwtggvfhNlaVgUW7QAxgnnw7gqtMd9x2lONZfBmFLAtO8KUTzh0pEw+s
Y1RMikoXqzn6W8u8G0GiyrKdB35UUvEauDh3tW7wBthwLjPln/6XCjwfWv93
5qTuuPcktKQeCmvHAJ8kTlQTwI4GanUXZ5dfi3kSsCLzwaJEceI9pjSMKXlU
ggzEY9fWgbDIe+6odLMSPd1UJxWmhiITWktf4sGVt3iFXfv1EDPZ7v+9CqFH
MmArm/3EwbhCr0z+HMUHeU+T0+1TMQf9xSrzifjCHrrxP4E8nqZAlAouBNUo
it2fxe/un/8kWXhB49wyw/nZjqizWwgGIzQa+/eLBdeffnobFjOwglLV/v9g
K6GpIZkojCua1TT5pUkarTuHqSIOvwTI3uYLzwAkpL5tr2IdM/sJDPYoajJZ
IxROsr8nJ+FNu1qIsk5/vBlWiWQ+IkOrawnDPJfXaitTywK6vp8ojBcxbEKd
h1KWZMeIiJKZL/u0RsBsDtL8R3PAWh/hw8/6xYP8opLiiawtaaJRND259RXv
1NWLoZ4NneFenRcDaXLNd/8B7i0ZhAxO99yYyLW0acX7xQaCto/mSzvO4AM7
J5jQ/w/ddcozjCWuxLtnaC2eQ5qSv7h1SRoeD5fTe2CXAj4r/vSa/8MWqjMe
xqIBefxJqouUXxpBzv8lAVu6ugzU7UnOOeqSyaZ5zEhcCQXXupGCV7goFqBy
NipDsArtC+OqvZk6XvQwGhjBrOLtKIpvwgznjHgBTND/kUhP/iVLE367NVJY
AEGSZjrrshGJXJHXuXrkC4O8iJ7i5vndDHnpslwCMuyD6qTeZ3+hmerp9GmF
3yGub5tUJABWgII5vciIHEOI88lDsDBu+GqB+NmuSCtv+YmOd386GxLqrfBM
s6NEAbaUtdUtuj2h/33daXqIeGplcrQ3aCiQDZq3P/1HBWi1wW/kbk+Y6oz5
jgDcY3JhEP4oEs1XZL0jYGKEhXfF7qjb+qvzV/v93kxrU+Amvjk/bq4twXAA
8G9cWaSpl88RS6GM0K+jsm0XzXT/ZzQbNCh1MLCAygvErU+uwJ/yDwTOw4bq
O9e+AWTNy3XsVtI4tek03onJekwrjAsm4Ns6XlinN+0WgiD28QhLoNPcAi6t
eiRhA6xsONZkH8jEx8Ww2YmboO0IRWMA/jylZDS9LqnyVgtFc3jp1CgKoMyR
4ICtfv+1cPJ3qdPbr50gTeTPoi31BrevbVNM6cSYMh/MvbWZ8s08VDpTIjam
XyqhLCMXYQNuOQ8RRVB8XBHr+2Zo+hl/RzHXwRZvgPcTzGVzSVUm/qOTkDYA
FrvxsMaWMAlcLakAIE1Ozw43xdRey2+udE6SC0NyuA3fDGqTMNrOQolkvxbH
P3gXgl7wgM6SPj3ONVT3SpjxTuRCqf1QfA1oXhbtxbR+rPhKOjfS9PXFI5C2
U3h01G8vmVtL/3HG/ozf9jst4ydYkWLWfuMrLEbAGbLB2SzsdYStiyY6Cgmu
ZvgDXPA3/iiUBydgvQhGwuttvpxFg5XDocnkyuZRIMy2WyXkAMfDLRFHU6JP
nD5VkuKy9sHN0koLgyAeeMFVgiS9pHPczQcK5VtBR46fDJFxk8xb2/cqHUtV
LSo339CYqBohxo7f2tJWbTODsL3NZ7dWRt1ZTQPi4a2IvYuSBh8jAEzCUNa5
/XfEvlRjk1ptZy49WD9n5Jvqg74rNaUcvdcd2OdcuhrcuQh21uK9F0wxAkU4
DTcvra0JTZAqbJKj+zBEDuOzScFchcrYy6HY09RESMd5S3BNyWTzMg0KPYGa
JExOpEbEkEwc0qlkiRMKbAGSNmH9jBR6BZRpw8LHor1zmLctjYhLgLC5qzhB
qsZ5GZGCgVLc7to14TNPfhWSAg0n4UZ8s8LYbWaK06hpU+6sdRS5EEO49Ntd
tgOmCB4A4DV5p9FUL5uV0MIcU2OfyutTb04HfNn80HpX9VwULTYAybPA3CxM
iPbTHchyhsIcYgD+Ib8Iih4REJSJoWhj1vpbfOq+Q2PaPvxxCRx21IW0j0ik
ZPi7+9qQ2CCLEuCvPZm90Bqi0lOPHisIt2dYEPonslXADwxT4PkopAEQNPXL
entMbG2wwrz6FrIXSfZvBbSG7sn1njkKL9CV/JlpX3XQbaCNFVyq1+ZMthfq
JaG67qilcW6P1XVdCa1HdpDkLoE8kPwSwCsXxPkKN/mqasM/ONidWwNHawxE
h3rbEsDi3GmN/kJskgG9cn8VOboa+7OxihphzJXwmOKdewfxdpu6kPDB6xtT
2GzdtXCO1um5tw5Ib+WPXBIJZ27sm15PHVIlsGvr+vCtq4PMqk1FyGVK+d/C
DUFzUpeMwpZmtxjKka7u+10MyX4wqIAI5JCs9s1S8J0Uh0ZdHIrQasanBrp8
k8AB9UK+owZcvELjGdlR+4sS/6w4HGJxT9dvHJ92QqSfuKhAwDshKf4UgWXU
5BNdRsB5Bl8VQRxrvpFfDxW3vSTHietH3Ye/I/9Ii0ZtEIQNfq1lj1tqvzvP
V9ymzplOtptrhV4ZcGMhCmdpUqGXpEQpLVzmblhM/2z1xcYO8JdRI6FTCPJo
BAYqFPKxeajHoqxLtP+m+HPwjDut9tsaovAHwl+RCqxvf+4znVkej2Wlz/TN
Ok+zIuSdnNA5gwfGxcmCWZ6rdtUhUHzItvZtXjmj4KHwcBrpI8g2LUxvWFzH
jUrffMsTOFk70lEFWKg5bHO1VRo3csw84izx28IMLYl5cEnvgfRGUS14TYj0
bpPCpnh60Nl8AQqCQAKNt2zkdg1OXKOqLIDgIdzEcg8LN7xWPk8H9AONFONa
/V4hO5Shaamz0jKOfNe6rmdXPzxvXWeFDKiSdqIvMGqagbkeKufZFCbMNSF7
kiTRd+9il7CfBoxjCS0JoYc5v5AmaRTHSnIBBE/CpM0Zn2XrcOjUacJcVr5y
/ei6GuCinNHk7peVexpZX7Ww948TdVkrea3Pmcf6mQ8bfjopdxDV5CXR16aN
6nnUaKBGxh2YnlnXXIBw+46Gky7hZOZHUdWkPv0+4d5grEGqEXcB3hP9fmH1
w7bMENV1KhcSsF9bQer+KwOYIzhKwVIIn4EI+eNZqY1st13zm9BaawHU+7ru
Y1SxmrUFIjWQnV0ssJ6CmtDmTqrYMxUIepqcnbhmvaMDNmEdcyUP/gopWDlg
BhSlf6zWSBrIujmz2MHsG+3k9y+qw17CA2QbY1ZF4TR8d/ZRDwysBha/GZsm
lboHehrpzWn73kPrMOsjVc76sRiSkUmxHiU5B979R1b4Eg8+b/yqbHP4QpeA
NyKiMfUm1hdE8CJuCmzMC82X9KGDbGbpij8dv3AcWejphsKlgAZwydjeo+PE
iHEL9e5EIMQ46nmwB1uAbzbAcczll5TotjUeu0Ok0sAeXTOoAk06Dux8oZE8
HeqPB62qFNpGEWkqvoJ8jbv4fnK+lByjgVzt/b/+kEUZZesUeyoi2ZFAtzIN
rh22bSl0ePXuZAXrL86W9agzHpItwx6X4LK59+qVO0HHWglOVpZb8KeLn1Kw
p9rZt1Oxqzgjf/AbhXJg5WUCPrOE8hpB6FOUExf8nuRCIxj9mpbR1yq7MbCm
HAnOFrNTh+YL0SxOwADStS5n884T3o/Ty78FTUjh+TSZgF3FBvUsSu47pSrB
lr5OvzQGwOXl00wl+EYOuwLMmMIvGkeTm0ULyFF28eGrofOPASwfc7ZxU8Rx
jLlH0gbYfAC6si+/EPka4hxSdws1FX68JAJLzoltTIUpYM92ZM4c8WvOYBeT
2XsZ8W0fdiIrLImItUpSw2iMNd8Dce0xj7JY7hs1VEO/H4Cyzm/bJJX1cuIa
Ae6efznxrIs5KGBEVogdXmuJOe6iGQBPICUrP6vwhyKbgN06JxevOhRsFC8N
hKcZO+Uviro8tbmpI+iZyry1kxCHL/k32ZN+InQnYacFUyrdLfWcCfJmwRp3
OWZPzkULwva+C1fw/6xtcz350+Xs/fyBvaK9Qjg7yeiHPfN+mUtA6Tkr8d3Y
hAc182m3HCD0YqRE0V26Ns91XDEeP5FXwtkZXPDMi/6T1APsVDW7osv7dMRu
7P+SnT0LdQLhmDohjRySqkdLrulS4sWt3YbwRfdqjYX1j3pZNM/IkGDovH32
jzXJ/NfmYK4ERNePbc9WPJEsP9n6cpvoSHj5X6I+La/hHLmbLJ2TnolLSLEi
74D2qWvDxsgQcpE0V8WHRJg5+MYd1XpF7ovqNAOCvNKiblmTveKizE7eKZw8
08PlJ5YI6Qs7bgORFgOaZEdbVw4OzZ2NftBXMd02OEMEwC4CN7nM+nRUm7Aw
Uiw9a8FpgZGyN+vVcvmIJb6JZe5UEkR5ei2WzVqRtSXL1UfIpGGCEYXF7+g4
k1hZmWVRSRC0cLGrjWHgwh5vl1atJI+5V2/O+tkNaqut2iHNhR3QFuUXzHss
ljcU+DhbslZ6LfzcQUn9+4OHPcEzS+hAvw2MpJr7kksE84eAt1vGnS2TuOhg
3bjbolM2aysbWphKpAuGKozTguLmXpD6FaVFwaTR644AhFFpMlvfEsCj3acr
ztWjA7QEeA3Yp3Ukg23Vj4Lxuqyb5Vnyz7Mv/V2t0mBBRBZwqvETCXBWgSli
O8NaRfFnwVEtEu467NvbnNGK/Bo1oziA87un/KbnpVLaj589q5KAgbRP6EYR
QD7uTsY9kj+ZwaKgudX8vDIQXhIeeU9II5fRi3ptfu5BPdWhu2vpdRLsAvoq
b72X+nt2lB7ZL7tutJSYUtyMwMn2lsEqQjpbCMFCNeqYAl3d97wm5JN4riVp
2PkaGwEibrCJvH3H/ijlVHMIIkRCHkCNJYnA4mXDCVD3ZRmK2m8R3WUfOyLt
2xDrv6qA1Id9dY/BIPXqdBNLkHeFojrMXA7y0Y5NpZIhoFUOVum0Hfi5B5wn
1+Hk/kOiljM0jTCA4uSH70BSJVYcq42etpW8mxlVhFVwqjGCRFniONuIV/d8
WyOB/kHB8TCipS63rhnrA87oQoAzMgTKqAJnJNRT/bQh5kKFjhDN8lmNY4zT
amzyZfFok/X0/nsqmtDcHIGE28+tBFgeAdO0oxKSvW1iInbHvRkKIjG+pNb3
OG2tExj0mD1qc4jUq1nhpsqCkpIKocHS38X6EuC261MnLuyoJ7er3Y1KU4aj
ArxqCDdJk9J0swjFUjlfKciHuTjv2SPpuEw7E0hQP4DahxwCUdLaGh1tp66s
qUNprO6REfBkgLDnIYj2h9uhnK9Wbp6MIBt2ONrvp1lGacb0AWZkyO8E9opq
mQJ7hSZKTnVDZLRGZse4+y1y0jnE5y0NfMhxhWF+2thI4FSISNR8AKvbzA3O
VknxLOJol6uPMSiNgTymwixHB6c8rFUEf07Bi4SCjY52vsCv+dIRBYVrYakf
UPqlUFU0Zr1I4c6spWCMZ6RPXSDJaAUvkUQMZpWXd9lldZSGszsT1YqoWY0O
RyJE/+Lq/VCNYrA31KJKB08GB+XD8k7TIUJ0ox/AnsSz0GWtbil9JfukPIky
osQHtW4jCsGj7tOo5wBm+nhVh4oSdMaKSoqTn8IolmsVV80fQ/Xctt4m3QM1
YrXzyxldrhT9rdb19YiJzjditWCzVYHPCYkCPMmmx5Kv+lcpXqVcWyRIqFIM
avV8chwNO6l91KxdtqIYptQxTvtoZ1bOkJ07cyEJiFjw+HMSlsQU+JMuD/mF
lQbT/SyChLvDRZEeF2ZE74IvnLWMDNuflO83w1LmjD68WBsyGjWD9wFWjHQi
Wk6FMbjslVTQHH1v84EQKKxSv+E/8VMvxkACdWvOdFPGywxqlJ39yPbKDQf6
rPpZsaR9rwoyt56CXeQ36ca0E6Y+F88CV+kt0lb03J8tyh3LOsfs1y3mCBXa
1DO8rVBjlTVm9bSK1FmFnb0M7BoNVXqjoWyycj9PiwDbA1xJ2RGqEB9LdQ98
053qULh5v9vKYSM8dA3pu7mfOX50E4ayf9OPuU149uxKG+Zw8uIj1jw3y1Rg
9c/U08pc5at9urgTL8ij1viE4fFSO2vC4YaMvBiqsU+g0+j/c8kLW/TXI4R9
HdAZ/XVXdQXZ9WpIstNkj48Q5O3OYSQX0eyb990uDmbM8zZ48V9G5ezUu5zx
PbXi/cMOK/DFFZ4tV+bkLmiDDTCq/cl/EuDLoeEDg0P/B8cPL4XMfegGW3MX
RCFiOcnAsDmwtUce53Gj1Z8Jec5V/97u+97cLMlo2ypJ/k+3oTWXoPwf5+P9
xMs4im2BDOCh3TvLFTo1AwH3YSEV3zK/7JmN4Zr8K617RnFPEY+NLRZz7GFR
D0J6m56+W+DBcq5g6ThmOHuaEMB5LMdoMHPtU36GXFaQQcyrmEI+jRYURren
skrFqC4gt3Ch5QVBlQJou3VKEtzfNzKNTYhDYg1mzHZP6RZVF0b2i0396Srv
a70jVVZG6bAmTWXI+uZKw9oNGmAVsYF/kw0mppj7EbLCpPtE12FY81pHCD0A
357Zrgz9VPg4Kft2JKAgvxLyPQtnivtrLnfRqHSj/1eal+HuiMsMW5DoBy4a
AWskRh2ub+oH4Z5ORGv+yUC59Of86TfJTvpqq5T6Vqxr9MH0K/jgQhZEgep/
hmc49as++DkJLgL6qeFwOQeHUrJJJxr5xB3Lc/sEFKr1YqeL2y0Bs3rZW3oU
0DnJVNbE4xDvhrTn7ESg+Pu53NdWJ+pOnG6K2/hQ3KYKPYEYDjhwP5SinDm/
HkY2uVlz/q4ZkrvbJeCp7jigUEszh3goJhX2BtqJGFtUMPjuhPePZcv619Zn
ibS26rdz42rhdV37iTzk4tHZXiTjNh5c4PsfGcnMkcqdcxnErR3MymoquXUW
S1R5cJi9ehDZwCrpqaGMhsLcS5KIXKvSu4Bs3z0zA+wevlgfsJKV0V4aSOmt
oeX7W0CXwWQyN4cWWSSeilVF3uvZtJpCyIw3F6K1BAlwhH0eIYs1Z4W9PeYC
HgE87ggrOd+B7zhMw5I51SjL2WH4LEK6yI88ANEc1EhfLOvLPHuFGh1wbIqd
NEvN43r4LtMLrmrPIdDnOCymExcIE6CqIMnEIyF7yJDyc35xBp88JlNJbA7C
WOOJk4EN82Qk7XFio+pGcvvplOUDomwqZMQJknK6JhYpkrSshpf+Fj3geERA
rsRdc0u5SpVXnyN2f3dDulvxRJm7J+AeeYM4817yRS7iYUW84reN0hlUfSYy
GneGmo62CfQmUB9Nb5ooae/W2OCWa978e+Uyeo2YMZn0b3azUoZyOg2gQTck
QFnZwEppKe1u39NHJozecLY1KeQI12P6c7TzHBh4i0M2TQZGlVa5j//uZ2zu
nVVi7ksyNP8id25BGnkDzlp/Aa30oDnsI81TqD8PrRhOtRSOv/zGTAWM5XFn
sunYruYHRlSUZ8tQymqrD7GEx4lkwWSEe9ehCBRN8tRYZfjsDObLvdVSbyxA
yholVeD+JBs+EexzJ6fb/Ej2BgjinwD8vVZr+sr++eOdHHGSOuDd12O5WaAg
g8/G//wJEa8uLNDVM8YF9I95oeMR+siXAVl5IUWjPIDBGKvuDjGRZe7FzJP/
4ijvfgyUxspsqOpVmM0aSt4DRhmaH1s3pUkY+wBz+qsf7nlQ7qB1bO/DLg+I
PT1ovr2D4q3C6zHrGeQwWcg6jisTWLtcpI6T2tMHoiHsMxsvBdvzab/m8rSL
6Q5sqoLYj7Z3ycjpFpz/WzQRpcPfCnP7jq5gwEJbFj0XSFxQ+E8vK/bXtAjf
mm1E33vLOmTrKLJhZZ0ntDzLDKU1ZVuM+qcQslmZs28+CiwZ4+owU3m7Uv3u
Uc5D7Hp52QQVWlsV/ETT13trriAVGDEiNK2p2aapwLT0hJICv41/GiwT4Bz8
EEMScv/xieSDqAPyEJStKm1JGCHxMbPNTErSrN0WPcXh9vz5kU9r8NjcWHDk
rlPakW0uTySD2ZoKggpAJ0gSkLNZqApoHjehSrpoQJLMjglq30vob0oG3TtW
1ct5KknYncs9m0y/gS0xa+yEdp2mybUMFvKcqAL9nFoRxcioQyIvNpvnfyjV
QtBJB/lpP0SjASECvL68JWHLOrrwX843scN5990gwPHSkkbkEfeqhuM0Uzu0
xSrvbYTZ4AHIV6cJlqnQWMXHmVK/P2eVUU7ycqdH+eOzMeGlDWMbZLwjFl8Z
CnOJj0WJeEaXZWmIxu5JvROqYPyRi53cGvmELY6CtGAg5gRRT0Ex7q1lKDZD
O4bfnpHgL6s52WVnBNUfJBU0pEZFDEDTZ9oJeTtjOrRX+ShVMP28NG30B9Hv
RfSE1lmd/sw+jfF2Xv5CJfilSXnuUyRFHCcT3fkQBRPngpL1a635Ad/a7CRb
C1crjMYqK5RtFLs70GNxONg6a/j0qiCLlPK1pMx1jHF6iTqxEM307yA5DiR7
EF9H0QCBPRN2TdE9eelbavPbjep8Xnll2Vq6AOH2XfRajXuuwG6i/ZGARmXj
Q4B2bxQTP+cjP81rwg4t70gPeg48G7nfasNVXKflBJx6eqsIA2nY/Ew2Iwyl
Cj4spkWgJo65/DA6WNPqUa45JnPmceOiPODjXpANhGTniwcpfbloY4Qkd9v0
wFWVvaJziH2eIhJZisSJDOpY47vqV6lHqWibOW/049XBjtyz9Ekq4vC24cIX
kOfTv4PCBqihYZFIm2635MGVPuukne/m7SJudp/V4wp3IAlLi8GFzduIIVsN
yNA01vWGSt7pIQtp2JkZxO3Qpt9bxFoDx7T2mHnW6dO2CQcoiuD80DzsfoSY
rs7oSDJP5OOpEKCVLyxwNV0mVt0W+Ffpwa/d99TzwmC0oajs2ak+1XtpfHPf
iAJQQNO5qa33+j2yUEvb6kZkbtkQ4OJFLQCZjRjXAjBimEqRVZzFhGl5F4hT
NAP6LMbHiS0HSz01q6OKdzjjjWeEZqlJXpUe2qBpveWraYOHC9Mr5UPTaF+a
w68u988rtipEryxqie+92NDh4o0WqxltTFZcmmqOGvTMICePtGDd5TH4OzDY
ZYpU5KYUP+4SRyQ4fmTeZZKYMglWG9qjVgtKiLridWsIEeZKPFG83iYTQl03
Id0gVEvIU6Z+Cr6V2vmGad1JMF92dw3Gedm9ZTLr7ikpEVDsF8tlN6Xo2O87
2o73c21cYwGY+sfV0XRnsf6RpKZB4mj9Ch2C4hbyIyhhBMon7oe+Ve7qhGqh
6QveybX7bpAXWUpZd3poxqkckvCqonCrTXAxvb3WFfr3cBTIBveq9E9e3/8B
W9QtXIyCivTY2JOSxRr4HDrwVEWOFtJBNsXiYpDgANTa8C181jPxQNAe/mAa
IHeMLE7/my8P31o3CbBEqfeK71aY4l1wnG/voqf2hQVvEk81uyfcUGCBfzEa
OYLIhJNV0VdWN+jWWvcnVuSXR3QAOGit5JMR95/erEAsLsqTDRNMgKbdAg1u
Wyk4phLLh57sO5RN2Vrj6vO/vwodUoC87Yp/0GY9P0u2Pmo/HNOGD+0yQIlb
VKvLqN7rYSXXS28sp3rX4Oy3MSEY5j2MZNRfOEoSjEW1onZ4cxtDo70A89gb
hxKZnVSv0bv26uF5zi3f9PRX3o8Sq49YrHNaoiulhTyjh7DJF9M3Lyf7Ii/F
QiP9A7UPjaFqHfkwgoyB1xfEj0s1v2UC2FrIpABYCQL00PX7Y5wcrqyX08XZ
80Abglqo8Hg4LOg0ixUvwqHF+9cA6wzGXjABcQkG0HGeNNLwIOy0SK4vvb0M
ekp8hiWJxn+JGpm74W4Z5A45f7rssDHkBLphB9AzzYiP8gnegH4LR0VQD/jS
tqQ3xaxQExsH4XtydDyvvOcHr76ACCXpJrEDClhVVxySBVl8Hhc3cEwoyf5I
XaC28lU+cbP1F3llJIrz8bvfnESgz/PExM9bfqrfv2HxAnHPn9r77nCs71x7
ZOo4iOLGuI+GM2XNWEGMWlDdb+4bNoz481x+luqfhpXnQBvE7xXmoYzaoslj
fH0Jb0GOSDo91tAP0PABxN/9xXC8Z4IKeaHxiILkmClSYvYDLLghDkJkJdTk
XQ3z4tbY1PoVxUWt5h1173IdfEh8PKNHKVHgVj00dodX8iCwoqZ5KZs/UIHx
urKz3Vp2AQbmrJFWsiq8olvjfpQQrV7F2XErQlMUbIqFOUn8kxh2EfiQIwbi
kZoxgn1mdU+6gUj7LmiRwuDq1Rp9oE76UjsbtaGH36ltMOU3+LSppkRYUGGa
cQY+K4gkfuWjs+Ty1+ZM1dv/0RwM90E9a4k3y1KBBHHYRU85rk2ro4X+Loec
AAKqY8lstBJQQ1wZge2dzhuf3EuC1BAwVA6X8TEXW+RBpQtFmYmdZoQYFYW2
jtResdwkjCqJI0tZeG6sPLbTvmA8vWtFkSU/NBtaBeGWlNXle28tjBPJIt9+
EfQjkq7kUKPyvGue6Y9nUvHYLSnPLXRBLz6/GubR9k4GjpRIfgcCsTFwXOt4
jF4FRBA2AyZQ16XYGKH6/ThQ9t18MXon2sj1MwAiDqmxrFFNG/ljU09JwcLe
YCA0Xz+HqtFeegDZ1AEZQBrZ77fp/y08r9GODX8HfoMWBWJZ1DssUtm4XVuR
B3d2fVdG6XEbT/dcPi4BeQ87eJn0oxbhLPJgJ7+BURq8ToO8LOylJPAffPUY
eu9PuxAJx1LeX3xKrTdHgXmOGQDYILsa84YWIEKMK0wpbOqHt+DkBBgFh2+H
+fYkXoj8k+b19IMGmi13aiKG2mp7NoSQOTyc+6s2Fuwtyej8Hki7eSlCl5ih
obF5gFvx6uLwlD1RMcjJFuYo/2OB/nAmUNHDtWAcfCfgMYBzilpgDs8BFPsY
mZp0nNIgEecst/FIJ+tl0QM26ioeUQYiNEIFOC0sj2fLC/5ERBykbca0f/8d
PwgW9LahvElc/6KAzWa+6qLK7aL9vfEurrjWjyZ2o68VR20r/d5JlNBRGdv4
I+6Uy7HWHCZrW2R6dDC7wrxaiWn2yk/tY6hjY9NfKe5WB03ZEPYk/BF+EFva
c3UvxdtZtJ0DYVCBOlSwHFqApHyXkZ9mx51SLbdBRd/Vm808w9X2fsYEC+Iy
Aw9TMQ4FXpxXoZzB3foUT3w7jTi970KwAFPRYEaLLsWTeMZz+Ed/g9Mws9Yq
JrcwELHf3FRet816XUskgn6yeqTzi0NX/n/xEpCm9nK18BJMiT/AM47c6ygw
14dMz5R/GA6xe7RcR3+lzyqK3YlxlshsF79D8aDiR9ftwtgERcJEeilhlNhv
pbeCXO0ANBvlm2JRPMMYVgtpT3ep263r0AzZBURVk0ZIB85G7846z22vQ+cg
zUZjgcuqBG9HizrxJqZdGJlQGk3WWXOEcVE+6HtDf9/o+v3odaugsu7XQ221
t0Dfb5gUJ7azE3sZ4xkG8hMWwrmRjHWwYdJ072vMBfICF2LfA0u3qSsAazIt
kWUP3ssqUfHRHVocOKPV3HfIV4xhal6EJ3WsJz4hdhznq1KcFillMSBjD+u5
NfayuxTheEGWXSkioPQKMdR2csWmWJUV9b3J6jaL30aBdzIXBSP8Nt3F+O2r
SH5jeg4Vvicdh43BQVpREwrE2zdc9YkbAG2QZglHrADZENYFUfRgDCRI7Zb5
GcAuIaxbjsIjsT021VZM4cviCa2C3MiidRysWOSqdvqveu1nVngNbMem0T/r
79PzgvRscq5zmXP8uR0XcxW0A5lorfV4Re77oYULCd7WAJwVQE9q7Ci7k445
/spoDMKXcs7zF6JC346BWGkLfRgBPueljWGUVnxLViHOfSfsvYWA52G/Mzf3
4S0PlPjISg7zBIGmLMu7V1YBbQxae7U0uPPrCYjeiQ9hrRIoFvbhuBWRnOTz
MGJG8+kNJ60lSpxwBL3Wwt0sCxhPChN3yeYellnpa+n9QGxedIPXdE5wuziJ
Xk0dFPqcT3eP5JNyNrn6KR5/obKAt+iEnxbVIt+0gCoQgmVkkFg4lN0TPw34
FNtrgd1FU8lKZbDAT4HZHXJgfM19qPY39Ye3Xwe73TOSXjGlQXKZrqAeRm31
n/dLzaNdB9vi4KDV0USsZHvdF/tX2CfjB9YmHTo56EstonBtaASyD5gEt4J8
iVCdcK6SlS7ixS229JN92ehQeMxf3UlfXTVuVtyH7UrGTOryR9vYU8X9xdwB
kUACWM4OAh4OsLFIikFVOl9Peruk5XKnGObS6/3jjRkRTMHsfyy6s6Hd8kEu
HqnU8yAX9n07VE2L4w5uZhWDV60WwZ8Gm23bTj84Od2+AAcWhQOPit1mNtdY
gnymonxzbRru8EetHx5sCk26RiB2nG3hdvsAsXOcc8mDD+fPG747VOg50bQS
cueNsPajkSptdvNgMWJPt29ILqLMwYCVb5zLVJKPYrioLMT04M4JSCk268ZV
iilFGBOWdgwMogHOO7yWIqkpUl4U4DnLS8rzXywlfdd5EyqHFsE3cYTEtE1A
J9UiC/o4yfvhLOuGNuF+fZ4srwNQe6UJGSh3jXJlh9CBzbr3GCIrRTHmP3z6
cLAZrvaXfcfMQM4wuPXy5Ek93S6oUGzgwgkrSTifVJrC5N/PFvsg4uIAHOzf
asVN7zBfs0IeOmasE5FXsgJdaIqHqxkEA2qu8N05yOoUdgwykzTHqbuDhRWG
BlB4ugYRXBqahEl7NfcrAzodfaFAAcHpLqnN+FLQqPpe/76b2rISH036lac8
BT/BypKa6cF8oOP1u/jaAlh2JuZyi/x2W8qfOgziCnluA76EvSN2efWhswb1
4SM8pYeIqYwNXID0aKReguePDkXbR5OkihDXGicI/zLPYo9IXGrqHmgef17I
Rgg//AfQEMsHa3oBCWMxHngjLWeqo5qXNFoB70S5YcjDo33G18d+CHS2uJUV
kEKK4iCHmzn6HhyD7n8s510NcuxnjthDrrN8chprlAYjasSb3vIvP3xz43SQ
a5Eqk4P29zDPmZa/DLJIfC1wWi+IfXv/6gveEQUQw4mAcI108JMpNcSF6WwZ
Hcjpcs4STIgw7oJOo7Ki++C1QwcVL6txr9Gch5ciz9d0GlXRpRmd2TgRWnLj
ZhJfHTgH/JmHHwstIQKzIdJp8/l1W0n8h4bTasrTF+jACWrWO2a6S+ZZJvs0
HJuO0B+RdDRMVdwrHs4RN9LiSKj7Yfmc2TkNPsiZKeZ7841qwTQY8KW7vaUo
cErTDiTENRyghKyzjkDeBSIAPOnka6K2C88VKFMzC3H7wZh/J4PvOkQQRX90
Ata2LKzgHq83IrkC2x1mFPyvgd004uR3xRJ8CaPHSa6L1+Hd7INVnSuOTKNl
o0r4hgQGwkcbgBsWnGnYhRphTwSQLbngLSDFzQ4Vrc2pVnM0/+Hw38uUNFjX
j+U1Pwp0zYbPl5VrT5wQee803YmknUpfa5WQVyCvNlbh2ItMNg++3BwQ3eZH
z0jDE65IECv7qYfNBMdO69XQi74jtwjU6u0HvCMUmcmLutLThLmTG+R45mSI
Kb1B8qot0sFyjE0UI3reoK0kvB4d3ScTTFaLzgCtAAY12ATDufUccwVXLZNe
+e74zFW8GpN7CAYDKqHCZee0Ibz7/P6sZcnJmYwJ+7J4s7zHk6pyML1aQsy2
OG2nfbrzt8kUfzc2Fn3vSd0sLu7AXxf0ehzSjjmug+kMzGQif5a89IoJxgiW
ugcQ85DsX5zH75Cr+BhPMFDzr6bj6d4a1I+z0oXmDbxCJjVgSbfdvU2uOBBU
ixPhe9RfVR4aIH99hA5xWy29DqtFzvcT53/arUVhZWiVhvW09dN72WGOPHzc
BWmOVMuRIPWpU9YebJ5sURsuGKhcrT1aMtnr9MJTr+2UcKhLlStr/+CMRVjJ
cx8WWawRtJZZDl9wnTIRcnZxW6t0t3OgxpSdR4EJBRknCY5eW5k0NpTHqYmJ
WSjVobLEhhjIxtFH5AhxTf/kB/TvmA4jp6svuc4bcqRBZbj8JuvRbYsprX0k
TeLaxxt+CI3Qv3hphOjGWFLMwZ8VkL61lGVPttfADTKKTZnWaUUSYo9RENhy
islHKi++v8nOde5qbXKq+My/dbUq8968TRUennpyFIJFpgnx7mv3ksKeqV4V
jeLHceNNxPHhUqOpDM2AT/HSqjBkf9nPCZSEYcPaE2SiwySSjuJ1hGx0LkZy
bDV4zkXhCaPHwDEnYbXD/l4qQwVgwnQvxJnV7OoN8WJU2l2bQGH3844c0ZRE
sUHxhD3LjOBlsp7vJcAPxdjSrz3MD/T3W07wRP3+c5JHsiSv84mxPWEJycVE
DtUyLDkvU/GaiuRXC7Rb4SBnjLLzRh+hydWJDAojww4vDpIqBWF8Q9tUWEs6
J5f2LpgSIUQf3bePH+Z8pbeywhayLPq+n9SMMfOuyodhFcLYZR932yJ62EGv
MSJnnpZHG404K+per9PrVAJ8zNu0sc1zs3bm7H5IpA7nndJEWAEkCweZuQR/
P1rLu2LNERt4+DHTUtFEqTDnB9aOBqdrNMY9C+6DQY14DjhkYAbQHeWwO6TG
5jes4b1IiFxYJOuq9jpaY/E+y8ZwYXN8W1F6lMF77CoviozWTZ/lPSOlauDe
u0hIJRbWD96ZjtJ92ivsXNpqc3R4DCDm4kuSkVtz+5y5sXM9QlQ4O+TUrFky
plBuV4LM9+IsazqqSVptobMP8/qJaGlbjIYd+xQnCKurDGrV8/0Ze/aCUYIz
O6SF7ZTLG5fiS3CoLP3DLX0ms64/S+k0xSa6KiD/Udc6sZZathgEsOX8jrDn
tXdx94SyMnuJAeFXH8JmVk5pvCROXCf2SGqKB2BS0G/gH546tEnAWl/zz9De
HdJqpZgAAEDyPZATuYOvRAUm0uMGK1Uhh575VRf6xzkFcsvTKVmSVESJVet3
nNlqLsGo/O0qXlRqHvVLaY7l1QOSLD4T+NWDJmVOkIR9TMtyp9cwEowbnh1c
MstV0xTWZD4nVvWAZJNFqbDry6ZKD9mVtsurvIyHINx3EIegLtDfmj5OHN/w
3rHLVwbXvv0ml8/zYwgfX6NBbVWpoNN1Di722ar9R++UPDBI7E8+Amv2z+OO
5lRK3u2TDiB4JC741S84oeOWUUCPfZSjoawUaQ7EUs4O0QJRnFwxvVcXjD7e
dls6SPId/lTu3xnpJRsKESVMRIk8DLa2Rf5zHAP2fp8OlSiGK8Bz6hfMPF3Y
Wc9BEVWy/SSZhSaR60AVziB9y7k5KcIFYpjokMcMBQHWZrRTIepPjvjIOUwE
ZCy9NU9ZRn7vd4K8iriLIkqWzSU6/w49V8uy4b1al+BMX2h6c0kCvBEUtM0F
MimPmHDEIQG/40FV8GWg2Vji/Dxz9g70tbFxrWupUZVpZFXYPcwlrPKMhYw7
5nerAZtXsir2UO5TIc8mexySLtsiNIX4q/aeOTZ0EwBiuzQ/1uJyVWmv3CeB
hk+fi69iyNnndI4Ppga+xBQMwFZlkrXyDue1a+F1v2f6ctWVeMgxX/WQl/Cj
78gwFLXxQ7rHQk1+s8RN20s3x0C2abRE0F9f3v0faqsVDZTeOtqlfMlapDOt
00nHD4wdVb6z0SaaqZ9kXGWq6ZxiDaRsLch1hp5zN3u9DV1AwhQVJS65kiF9
5LLT0htNjNRlLs80LlTLYy0Jp+BwnqT5g/O9qVL8CoE5DVJY4vGs/Y+mwy8b
1bFthUGlGy/RQ7knrZUmwsKGjGgNMGWW/5j48zb9ojSJ8r7uO2/YnxARRLOS
x3onT6kDAOnrmMHLEARzQ1eGc0ICo7CGOTzC5UAkV9sNf18FGOeDZQrhxGcd
j0pj6gV/mfE/QtcAbOkIN9ocI3phZxN2QUUrAGPL3eNzgMKg4F0f2BWvCBs5
raK9CLP7MFwhWv0x9Ty9kSJ1HMPwAZaEYslycpsTHtBxL/tzJFpZ5KvUc51R
XX9vtnfrQssPkl+WXi9UxkBeJ5bLEU4IFRo8gO9KjfbGPsdRfMZXxwVW8gnI
Bjt/n8Isf1jY0mfWVNm74IaD7ke8cioDts7frCrVcnBMUeH4ZyVuaeMWM4zX
KQDrtuHejMQ1oBj0UiYSiIIGf3Xah7k3RgqntHrhw4vOSW36v+ipICV7OUYE
n7D67d7susMiEp4z2iuHrGmZcWtRp+jUjk/UtSvopEIOMG54vhHzUwQxMnp3
xQgJi7pbmjyWtWLk7CrgimYcU8fzKy8RjqKI3Bkw+M9G85e1RK64jqmQ/hVZ
+L6QBkh8FBbvhb3iVUMVmVIhtS0edECXAp7OlrW9om3V7/i7PMan/71uJSxi
4GDJ9AiuhfiPNYWzRSG1HvMsxgao0G0TAL0bYu3xzl+l29yOnD4X08PIiDIQ
jmLexM/rwYciv+wSFmoJqhfecgMzKcnCuyNDgE45y36HPObeFW4TU73Q6tdj
GJ/PhFlRJlr9K4ebPv4jRbTNkXV60Nbick20bTxMCefEeobN/lWBVwKpQOa3
67/VB1c2kjXaMVemRYaeXjdEQigCEeBBuL2wpNidDvC12dZA3vo2c5WYz8jm
46HhEhLHpjB06oXwh+euAtogKo63pozpPdIy0GFVHWAm6QWEK5pcjGq7u2PB
1puAN5qhdGY6GFaNBgvtQtDdeD1WWp4j1MIYEL+6ChUeKne+nk3y/TY42W1j
+fEKZOOpBtHJ2y3dv8UXU73XTCqfAq92RJYt6HTHIBKBtIAfrngL5h5APpcj
oQWQhV9SCvDnQVgTpjkt8mDqzuT8cHD7Fw3EFBZ7GSjdbHMTlgBCb0tZ0IdC
ce2tSmpCLFUlwFLokSM+C1yApZm5ppMxSgPoTv4QgvEL1hyXlRArMVerClq4
cxhjGOKq7ldVMUJSEPdHUNUsSQ4NQMOLdBCuelmfVNajomOQTXyi10tMPF8V
l6a6KX/8HnOUN/6L8p51qpk6Hj5x8igaEYV7eiNo+edOu//p7ITTvK1DwMCm
qs57dnbAf9pFQ1UdyMLAdvDA/Bp6wjPXHWpSMw5BuqEmTXpDaCWR0CJrN5C2
oOmYnhqjWDDiBjRKo0+f8Rnga9vLhheVBx7/9Hj7aPZObpgQcmJ4Rl1E0+lD
7DHWEghGcporkyK8b6dqFEUjFJYrYDxVZbroYLVRliSvdnM9Rl6oQcpE/R/N
Lwn8zdCvKe4nnfx7hhEP/K9RPQrMFLJF8BQs/PQSkkpG+s5gWMnMTZ1ZhEWg
yf7NYx1dQSZ6w/4Qy8kBlYkEW3CZGocpt4YI29D8PLiZjHlNECVpDVrxqASF
o9kgzNncy/YPLhCvjwp2rBpP2th8tmwNX/1d0npj1YSc7vLeVEEPqNKZCei0
atXlopwH9PQNG/UamcQIIKtpCmG+xVtcyf7D1IWI8GB7jwFt4crvKgf/qoa2
1O7kC3aMyJ6/jLw7tQPRy5URuZ9lJ7i2I+7xOTCtOHm8jXV7X4P1sR56HrIN
/GdYAD2B0Txbc2nN/qmYmrRv7UBJNQOoeuTF2sMEbj+p2uGd3ei3hpQMscWx
NWSzShQ5SamAl5bj/NmHVmeDqni/BqkeL72mf+LEuaAPjOooaJFYGgCaA9Cr
hfXpXapU/ByAnr+3q6jg+7PsdouJ2VNyQXDRBjdiJ1FQIm3aqzqROmiv+V3d
J2Ujl5MewZmvsxAaDM8cU1iQCOHyCfn2/iUhHXsChhBuzajJt6FdYN/vxa1W
sGZMYlD624mMacZ9yH5LpzkenSpUlLIGJBXigInEGvk+puUsSWUhugM4NA1c
1gV4l4+kFbsxMVFzBsoAVEVtiouG51TudAmmo/c/lAfvTyw5vahAEkUV+WtP
vTT3SYvyPTIDY9XR0hR2/JfchPaWMg3RBzPRy+BlZfbxprYDKRpPR4ewTZbG
QPjntW0APTiwe2z5tEzZBZJXZ/q6dITsFvFHXv6sXlsfa9tgixgjCIrvJ30I
bHxefdpT+Z7NTacPYGLGGFEFUV2aUJ/+m2PVrEhDzNVVz0h+xTCsPgybHfGX
GFZvMei4r2N5aZlKVoxCT91SIfPn+F4jLXIjdA834LwtZOzYCXZHIm31/5ed
WSkKFBKLOZ7D0fgSPd7FQ9FpuKVGPRXvXzBrnoTsNLM6/yNIgOyYdx8irQJn
Xo8v+l6mi6Ewyw2RLE9VBqW4tARxIwE+dF+g9TSfjjoUItnnER37v2Uhn2kJ
5Nt55ou7qPCY9XypQRajqBtW/JaPR9R5H7PNRNO7mU6CjmwopjUpK/7VrKIP
NAuY2+oOXfYwBNnTqUra24zlDcFIOGi6iNYras97nXkQfRwJgI6HxMyXp72N
8L5uLstCJbtCqiDkI2k+JNLYe93be2n/rirmFAT1JcT8CH8IkWD5gjGtU1Iq
DHyJbeHSpm7Nw2Q62eBUy7hH7q09DQk3sUd6tCB8cAb1bktcbaYlYDN3sWx3
3oJMjXz1vrmGivf48c/GQJ9tNuLYM2jszXXxaTrp5r+nv4a//9mRZJwfIei5
+q0y+J1P0FHdLx6ayo2THD9xurXp9DToO8aPllbSIYfsQVZcUG8tH8IliuXA
6pAAE49fNW2TjoygPB8EABWA/knA7Rulh+8ke8e0wRt7QWpSJvKRGcN0rbNu
zEbySA2YrShj61fCkWXgmkCp31pm9dyXyXcjmE2FwKqexaiMAXHxkmjaesJT
t8DXybdQ7TiiAGBM3UVILffum8V3Bf7mZGc7+m5y0IwktByPMqllsLXNxF7j
OwPggvZLGZmXUmYmroZdtgJe/Zdu1biSajKOl6fWENgH9zoma/nElElgPTka
tQAWhz0N3d8egc264UM9caNUXSjP1QfdQzj9CXQpmJL+7vANbD539qNbKeBC
AFL0z/rwKD6mUod7BIzQCJZJVGaqS0aiHiC8tdLmw5t0l19mF8qYjNFaQvVz
vIZoopMZsWG1Z4BbqsJSBAlPv8o4E0kQrkZNWbQF8z0PuqiwsdGzWXzbNHUL
9GjP39niDQ1OcQGsBw5+yY/OonT2PydpQ6yiYjmB4/ORTDwwcwqQewIcByRM
v9RRFKLzLSkKwuZRuDuE2E0N5JoPjwQtHJsWp40PfFDxCd5NdqTZwG8tEpHt
vuN6I6mhucrJDuJP2Yr8Fhbf9dMbLwT7mCvC+rwNN1tl+klPe8irhn987O3x
aGyemg+bhEL7yOikmGcR4utrEa6QKTfnEA4FSjEGA6VSlfqWJuP5rM1DViP7
sEpZcPLCYBeJABCTUgwB03/wQhH6vpTPGfUvC8KGznY4V5ZHsmZWJDyZZ1LS
rS679+6RWJPyEkh2SJ6F6Qe8RMgCrX9k7gAVk90VGbueEEQObCd1J7vU4pXm
lk8YZRjs5HCQF2hv3CoaoNzdqPNcZjso79yqlklUr0BtLck3AFZCGHMkQ0vW
4L8AxmfHXjnpNJw6DHs4Bo6Oz+dyULkzVzX0fVM3ak5qHAKgOdWfB0FfiltM
mQKnTo6PdLUF2j+/Rmxs9bEGrjMPqxgNPAm9x5MhT7DaUaxVjPmLpE3/g1d8
ZAdXxBXCoyuj03UIvpQYdtg741N0SRw8unEW1PzPaPD9uiz578oDyB3qvQ7z
xrhHyHcZJ0VgSCR/kczT6V/JA2j73HKfEoeRtiqUbAC0fSsoaDhvLyT9I8/8
uFNV6T72VuzXX86h7TzpGwZraZ2Bzdczo3UEBzQBDCjm+tT0hhLKCy5SPYIs
ym7df39RlJg+3YrfIvTeHcJZTtahwehfGTjNmzeozZ+M0fJ7Zm/80GxjXkVd
w/WMx2/Y/vJcyPfzS3X8mRU2LX0ZIhTlU8ha7My6MRY1iBwGb1SqLnsFwfSY
s+Py4DHHO7tWmWJRY90Q2P16nRPc6AHHtne0nDe+Fsr4EZz1f85MkxzfPOOq
nk3xvpppzr+P5W1VghnEQP2+qvFkR62UMp7U1zArEhfQ2zDQR7AW8oGkRAcA
hcaWJ33j3iFpQiMMnYAQ6E0yoykCcYnv2q4T7DvESwTOtpgrDA1dZ0VqvdAS
qzRUDJf1LmwTUWvGY8+a65ZTOQsFkQlB2k3nR9ZeuqiP/wIuJRBDNim0siIJ
siFSkhLPnZYxwTHLa6tnne4wuaPHUsLL8RQ5IFcR3xLZ14wsYsEeuE+5EtUW
e/J4zdTQ2o0Fn2cPZBFxnr5XxFsDsBL0aZvTmyOQYEuI1d98ReFbXmzwQ346
z41C+TtuF7qX9qxeZD2etw2ktNSRCjgT1xK3Zv00y6Ystc1r2Q1qfdZwL6r4
aLAUnFFhLgNGvS6vzNx58P3AUecI0DfLDa8NfqDhepj5lYseqf6RVKnFUzsF
8bL/n172C3jVe8RZ+e20NPBEQ7dN+5jbgYOAkQLa665DwP3nY6VZpozyGuOR
i/t9aZRSm5KmNtXpSTCIRhMUkDRyn33EaGLpoxZAgYmB5YoydcD/VB6NIi5O
C92xsq3L6V4eazcc0En+bUHkiqqNAAoruP7slKRMYrz1qYP8Lo0cJ/6U0g7o
KXB761DYo313ixiqat+yfvbISkV9RAtFvaQ85CQoHTez6H0EPu+uTvUENxLw
7ZETrI0nY9yWkBs3IW9S8Q6AVuVspcssHFMC12XDcArMlcuraeNi+k9gWcQY
RkOxkLifnw86FnzRrNGFURCeKmkB50sCcPVXm9jrsSdA8CtYtOdVHNOzk5Gq
lNHtB9wz+8Wr182ZIi30PhF3PHCHp/mv6BUQKWW0Jzw0XbwCZQN1MJ+YCPvg
cIUnmf5qp7tM5VUQfjcCLPekgqJEG8ZHyW5TFxfMbKcJIUsF89jb+UO7lRwR
RCqgx+1+JDoyViz4sDCPhZeaZobc2yZZueI+BFde3v0MNvu1AeQpwrrZfUUy
KpWD6V8wKGqcmQQaIAdbjtcCssXVhofhFi0sksCApksud5lSJWVGjGgfVjkm
X5ab8f4ez3o8nDazdG+YDPE1y4BhnnX7tS6UoVBc/wMBmdoLgr9RTuKHIZiO
44FrDVnvOGPtEjQXJsMgXv4BMCHfpSSsrG0DxRi6KIz1p62IX759SDTcVyut
6jdGn+f8nC3+CdlpB9trrcxdODdxvtK/0C80BJWBJLCQeoJnJqxin5+equbt
onN5uKNRirfMLqNtNgoU8x/oY2xEjz6fx0JmoyXWqbsIbBbW3tmLeVs2xkU8
k6zsRaew2tuV2V0Sn8BQVxaCAbPPjtkBtoQfAN9D0/2/t8bxY/gQjs4A7rBQ
hiNznC+EEGCd+CvTWVxrTq8MHPIr14PwIkLxBv7/OxNU3gGz3CaKKBZN0h/k
nnMKNSFIKR1KkKbuWxi9lgxPsab7simbSKXbrvRH/OqL2vHFgEwGvG4ikKHB
73ECKS64ehXqcOU2x7klqpGlMeqp8AsC8X0zcHhUIuEfbCOaHPG+LmRB8lcr
Y1oqm1jPKFb/5qX9vwNZ2x9FCY9l1kcxHDBc340LF2aLz3m/9eBatGiVD6Tf
epf7RaDdB43qGiI92WvH0XEVUW65BFN/SZY9vYzmfZbmBfcgGAVTXXUzjfSE
GIsOLvfMFGlOJ4IQHX1IHYBwnQRp13qfa5RfznEQn3rVue4xU2/EWDbMg0bj
gO8q9+Xt/3ypvOz5fveyVNdHmFmcUR5ox6WuA6gCn1GhcjV6jCXA/d2gFb0W
Y6qjPxka35234BhHEtSZzsorFgwX/eafaWiZ4yJh7h/9bz0se1Yn4pdaA5ie
55lbHD2/2WJpuYaZlCAoEMGs+LI8ll21zeWz6cxrKNiBCmMLSDZA6Xiq6wWM
e4nXNGhUUZd9UgjpWHgZ4Hdek+jACmbLKrvY+2YtA1KXX0ClehxVF6cqm8yn
YDUER4f6IwZFe1fz7eDyyvVLCbNE35hZa5olBbtgCqAatkdITYVgjBhM/7As
OpfZirRDQAQTvb0mYvqDUT0nk73BZVIh45DSisJZhcKHVFPtFjdgQjtOc1dn
wpxzIFVOGF1b862Ync4HslQwM0JmftlAw5WFj6NyzgNJySZoeiELphQv78ua
CSFo7C49GAGFrKsorbh4hEROXdZyipff1SH99+b+fgLALpJi4kTHhSo4QwKo
b+StH7VptwY/IiAKTD7uFc5aDXeaAjQ/I6mHx044XL7sXXOfNUeYt+eH33z7
AogR0GT8F6iJhOa4RPxA3KD0Cgx5xUefGDqnKjUTnih+N8jvpCMcuBD6slld
2X78G3FZxvgFjfNRNm2aiIypfBGkpJ1Tfuzv0xrLfINsaLkFYELO7gqW14pc
5fR/gaFY9tG3Ckt4VN63lxMpOpfOHLhUNTkcr2yNqEOVI3iuePO/StdU6esJ
cbLmXjWEzKOa48eBRygBs1CmEpxqvB58upchRxzDdHCTu6UNWGm0uMXQU+Oq
z/QOkqrx+214dhm7PIU9HoyjVt4l/iR1BsAMVvBT9Rn18ebh8KvEG2fO1fRy
04MprR489/oOJPH/slRGrQ4xK9A0mv4oP4tsSG5adPmsnlr6Kbv7msU59BT7
Z1hJanTthFT237BWU8p43qTE2CMSSqVGJ5JKgaesNbwD2WU3hD3qihZBzT00
thONaeRdIgOM6sv1SzTv0KzdmqSLxjwqdoJqa7N7+hG+7BtkXuvkadyIBpAz
kOGu0iFOxFG3GPHJuXjkPMi0a0W9FDMOTX0KOGbUzLxAfGlrZhSIInRiP/ar
T80hpDIX8jSQna3KidtmHU+Bpui34CAaYei4bOrBRnziLKHeqpZvZDJRXxwx
O/63hqODRUZckH6OrRcON9T0JGm2WuSZ2L97pqUZTS7viXAy1z1m2I9ayVZj
3HKhY/+vJxygMkdniXwV8y8DUm+gD7/rybT9ifo4DxSiAL2xQPeum82j5ajX
H4j+m64aykl1iAMKcWexYo6i45dM75dV/hOd7CwqwayfK0HA3wyBw7GVt6Sr
Z9abRyESlpk4QZLo4ycWqeF9hze1A3LDlx+o8JOpWHlXrD9Yx/XUNmIWQeYx
iroZepHktKnmffyPGFB/xpsDFUq2skof//EEETWXE5L8HbuPchNnr+CWmD9F
cV/2z/An7nyT+zuEQJ0/hyQyHZUTPYlyjw2sZIg9f/ivWXXB4nm9W+xTLdpd
KcWJ8S8Oqd80GQYUUxDNJBqW6hSW0jrVGC6SAxZsblTv07EXWh1ZaHrzKu/n
Rcm39GDHsPQ4lyl2KMRQSD0VX+h6q4pnECi/8jR3khztHl6m0fqKtdV6JVjF
rYeenfYQF3lGl431Kg/w62keju+9rqz9/27o4y0BV3dEPiBo1hdeDtAAi4gn
8jcB3GX/WRRxz6cz17+08NXxbyK/6muXu+vwfBh4cLPUNScpal4bg4sFgUyO
LFA6d9NqEBmFAqy+vVbKzl8hEeT8RCX2/cCLbn8M3fznfK7BMVTwqbkU0BZC
5hqbj6sYu/UvIpT/57/jWuNFn0G7SnhFs1VEqFHjmLz4q5pA+A0z/gtnL+ZX
QT8+AqK0uKSKni2IvqZgfySuYJpfkHjQY4DrkwRULsQ5A+tpR7sjENUrtkeP
O5UeArR8jvTunkSiQQe2st6pG8fZlL+JZOZCFUK3KdDfcPTTRKBeac3FrVRI
AWsOSMcHLUDreT9F+VHKbBDXrmLVq1SwuInd9tpgDxlrZ0nlEu2xUtha/eEU
8xmxScI7NkVG1IUyJAopNr2uIST9/oLIACLxowuftFEj+JVQIMtOCWj4+VuA
RHs3c0G/KV5TyHxb1g+3LtPtoKn3b+H/wST5gr5f2gklpzLa1d11N4KU7APY
xXgR0nMIVzvTFR87Pnx8tt2q/fKHGCcDcwr+IhNz9AACMo5Y9Qlgx9nePFqw
5zII57lMMWrmzTqen9fifqs9+ZTzyXpSGkmaL0MNuYMtWZgIL8rf3dy4PAj5
ojzbETKgCsptUaat+xddE9BjcZ/jyygZ4zcoCjeV5b/A5qGUmvC1o3Qk0qi4
QA7vX5bsuizWyFOFWkTnYkm2l+vc6C00VY4KzyMupMB5hvUnL6eJmMo8DxWJ
tas5GLTbUOYkXmk5TNo0tqJaKcERh95VlojLnkb3Meb2/HMiG531eDkMuyxF
VBi8bt/0lVjAa5hmM3TGrHyruzygSCReNxPQLQAraZY6rLkfdrBpnDdn9Kp4
CdTjdwEBT2YPP+DGSo8U5It5QSBsh7k4Jyfy9bOElfpu1ScZnH3iZZU311pb
3Y7tdc4XdmhGQueqpiDwXfks+3wGSzI/Wp4m4TXtinjXlTKc6WE/fsb9j4tP
dC1dDfou5fOpPLuOJr95z8O99g14/li9jG98pT7a3MXJj9IvYDaxhUHY9IZh
NkPYD3bPZ4GuM9/K0ehWnejfl4Bgck3YxUiyBg7JtQwxjNK92EvFzpcFy7pz
Wg2V4N1fBInE3kpIpZnWueBFzhuSr238s3oI0zt5+KCTFt06YVDbXVDquDgA
or1evwLmXkULwUd1i+DQk0ftz665sANPHaHU6QaCw4QkhqrihvUNjapXX7TY
MVITxfASKAXsDqGa9rABtCnwiLAkMTW18YzB1IigOJvlVgjiyBqzaMnZn2TV
zngV2BRuzv6ruBcKhxGr2je2QFsVv3FlCCKADH3ECOsaq6Ptr8cb3ckCNoIi
by/Sz6P/mE1kR5P8L9wEfUuzngh43J/4PzXlh49c6SbqaKsDZ5MHVBv8ovbL
0rD5R1lLJpQkAaI8ExFf3eUy7LogEh6i426TgWsuFDkj6w1jBaBGiBYfsVRo
lIc4VozbMyp8K0Nq435Xymx4aWyC1qEusbBKmJi+g1+pKW/lH5vm3+RQR8xw
S+10YTH0arpMK2R6lhGxcpEELI9j6LcWoetRsLd+lj3gvBBCDR6Pljm0h59E
covcDWKfvOnhkHPaVhcu1ZF0RbazbKW6PvxonVb0OnJlnEqnEH5iHr4CLtig
52n1vJQbYYe8YizJoA6DkBy+oK58GsIsgwVZKnru8HPdU3BF2gxxtHQsPpT9
dSphlJf8umHkKZEOUu3SxSsGwpSvNi18dyYCyic8D2b2YnNOCPk06uGJniIK
V3qcO98CO8+i2/4ScPdsgMy7hey6mAdZEOz1tBb5L6F6k77jjWSwvoe/ci3q
Qez0IJkGfkvQSUIt8+7o+C29Kam8bZVJE/qVKtPiKOidPQlgK7rBrBziSrCS
aJkhrCL1s8QD+oQs4UDgBA391+HSUJbb8daGl+v4D1wV5DAFq5gwFMeGOweu
FpXRxlI23lJcnSFb1o2YRhH/uoGI/eZlrI1Qm5N43jzn0Y63YXgYVZqzpmKe
a0XadKQ/vammOSzrmU5UZ5lr9IrbzWagXgM8gi/mywrBb149vB9kT9IdItDO
O5F7NWaSeqUlMqVz+GPzbnJ2b0OmQMzBDXusM+h5PCwA9esk8H9MjCKTsM+7
IQ0LsiH0LYOA5NRKSbf/HgF/bp9R2dcUZcGKsZ+9wg8sqgBYLpn0tlqhaPcf
qupG0dLXybO4NL9ge67WIjMSCbFkxerbAUK3VbFVkL5pU+uj2ZHaHToiyIy4
coQj4G1BRAQ7AGa3x2c7UzIhjtdbNdr2xxEm6j3AG/sGodIgWtus9v+A8bhO
zR4hEL661yPjwcBOeQikLotMTkCz9seutwP4wiMv97MIskFZT9My8HwmUbLJ
loxg20HVAE0ZsblarNsbv6qwfZ767qI/NOe9fA0dDcQ2Gdq6sS7zO6NAlbqd
+qhJTmOYQuSKvybcktbpCO5Ms4/Xj5xrgEMgbY7kZETUppSxpoMA7ayqAqhB
Al05ElZyDzRm0VoFHdLHycpooibenkcx4aDCoSYD1rQptHwYNRtDnEPqBZgz
YToYfuiwqRTgyOfekGVmAfwJwJ2epDQvgrV3h2qQ0fjQtGxisy1gfVd0kmEp
t3qmLftwZ9M+SfZ0go+03G/RScX9diCy1TlgOzI5VGj+ZX3u6aHbRwwsSKLs
vrZl6++st+7owDW2EQp0ULG866lxlglMTaaccK3eUgG7wIg3fTtnyodZ7sCd
BqpI/Pvqgc784TedaHSKXYSuniTtktkBNsQZCAT94CiBS/2KyFjnRmorToBm
fpRoHe0YW6qio1MiLdFdF7w9sCLScbU6wOKcTrTRChPv7aQfQyZ4Bsb7Dk0p
tD6Y8WcDKug2dPkX5aQmCvlDA/Nr09bE3q31IY5CgmxyZkr8ASUnZzV+QYkH
mczhyj+fvTrKMkyqF2cAfjzzWheMy5ovtHk9j9zufC3ARgShzdrhN2+K+/hl
mVHAuh8EYaYwlxpm+hXueRI81DWtEx2X1D/Q5hCKpAN2e4IC6hy467ybJpKs
jjlOWupRVHxDbMH69UYTc2HQUnTNIN5hR+i+ABg+BK7ei4gdLB5XBsGUWvT1
xbvzswJhvuffGhK+dXCmgbHyZG+504aBtk3PCzKg8ku5IOQf4OsT2E1Smb79
UQ3csvf4+AKI518haK1a8WC11miSOWEGXfqQhn0FTCn1XMtxSUxKQLomxuv5
vkruT1MVDACBuCoi1StkyI2kP1hfcNVmBS1WA/0/kffNpPZpeWL4g9ssW2ZQ
4klfAyaYdpnWReTWl3xxo5tw/dvHpSeGAZlhQ77sH9vgsLUC4/I7f+0A/c5X
FBqLsvJTflaF+YNen+ymKXhVhNmuH1EdBDRodMV3EuYfMXoUjFKx/1AtPg9H
3FaFV50dfCeuk+cF7ZNBncC9ytBa2nO1mn3LsL5Vi0ZnjLSb+A7TJxarGurk
3Wx6SZwn2Qtzd2inXTCdhA9LYf462KivUpRHNPUqG90dP5DsOqMyaQ613I3r
U2AODq7H6q9isotHPnXK76/AmcU11mXdFzi/g7W67cMLaLNEZJYKvLAlafPX
ZucKecv06B7Q2mx0q4LgZ1O6lndV9wP25HXYoGU8sPfgyMG2B28oEVJoDf30
XCPOMRmVyEu8SMVtMD1qbTCxXk9TWNnRw5XogYmqZLqnKFrhZfZQhEZHL+eL
NZ4DDeIzvJsBoZLPrZkVPo+yJxMxQjOlgFRHWvMhH6n0LVfpYskkM4NdDt/o
uy9i/2ArPmquMefFP2hoauJGfFmwYDrbDvCt0BEYmUsB9IQbJE9pOQjL/SbL
lHxnPGdh7jOWwWAsu4t3Pq+ZytjZXVKMpSbONk6abVU2GCNRaMNxoh4e6D5O
IVbXucT4uBK7rkoRBWJislHWV8zhDyatdgRiMYvbw++7dHJvqlu5X7SbLbsB
COoppYkyPVH1MaQjP5/p2yJA6MqnPS6subyB5UWz2Y8dzKJg6kO+InQvobTw
byaTLpaH5P6GwTFlPt69biJpKtgiRXjEY38VR8g+KtLnt3sDKV0nztVYW0nn
WkHkq6xq6HzNBwvbZ9+vN0xoAShRXiXyLZiwVdep3ep+n0vTyq/pu+63vK6S
FuM5zz+vZ7OrLwytfuqEJqgAEW+dd1LaFDSZF+SQR8E/JYDZ/j534l7GMuDh
Cg1W4hHxeI8ZxvUQ9lquFUZDMfmTZfN6AMNR9YhdP+/CCuOnXoTHDS1AG0jN
WuTGpSHXhMPfLIsGu5tP2ayJ+1uFE0zELe8pBM+ZyWE2N78GuaQH4kDONRu8
7T/YnkQ4kOlIVlJH8ivjN7OfFCIXAA0iFZvMqZwI7F/BpbJD3qvMynSEum1i
oqYsy3TupktX+Gcp2Xy0exaku0qRZ6lVEh8XUwjeok6HPlPsnEez9W+AU9nz
RtLzlU9a19r00mIAPmZKXayXaiXvXvm82Trf7DOeOUK8Q+3kvLAel2nB6B4v
Ok98UA83XDZlHN+JY6uh62Nmag5b/YuOR83kSU+sfqaKwIYUbIDfVc6hjaIB
sRV+vBP5I7WDyvx+D/Kyi4rG0SLG0pG3QX7ZM+a9k8jNEMBG4r4UeDNVwO/k
girwFmGds9wS03o/T4bUSCdcsHCUPKktsN9Dwk7kNdEzgqs9Soisrwxmtyut
xUOeGzW5w1LCa1MV8oPdDys2jpHxaRCiB1xi7bakhN36U685LQd1Pai03SvW
BQxhsyoXHMRIg8JWOnekmy6ln7A975XApKCzMRGD6fDis6D1OUabtnaAQWOj
A7CFH1hp3AFZu/LtBl+y1t/EFb0KkvJ1kgAuxp4KzQlxS2lzaDRB8aLTPYxE
rUundDtyc563cGtq61pe/7ip0Rbii+ReBLTMaTzAaa1zRYFPAgfs2wPcXFHI
qZiaoQ7aXIauzb+k+4c/po0vlQqBr8CO69o8jVWw6E8Zgbsr3TzC2Fu+KWCt
kkRLW1VqMGUNcXo+8Q8E61zDxLrU2mr0DrwehQ+tDUbktyq8Jp1+6Sn/12/T
qIhXBYIXbzgJUM9zA9wpgSuJIZIcLqJcewGQUCETIzW8WrZOvF26HLmR9OJe
TKLtU5NCTVcEZUpmReAd29dZyux8YwrVC93Z/btQQXcVVC/XmO2UyeCyMDIo
woLhkeMdXxIMQn2uCI3MjA4pZqAgs9WxOj8Ux/07dfrxVuQipAAW/3KKC7B/
/6tjfrbnUa9HWGJG6O6A+6xSbNCOSfBCEYMc/+Ub3W8L+cIbd979hRCNNrjz
J9ZeKZgmDmv6hfAOuro9ALYt2Kf83FtgnnlrZ5Wfa8tUvwMWCGMMwjG0McS6
JFNidQNnAcpHNwi0nKrT6yccC73/A2ZCkU+srwkFIyJ30hVsdotdhwA7Ld/9
fPGcpa4/JnlEMfjmKIL5KUHMcqWkxTStMlgrHuLNsJNjxeWNzooX0hRWfOm8
0jet6OY8lb4nz+5UZCzbW+rrmmDMSykOP3MXOHvoEyZ3wiO5AtMOxkSzCRYv
wZUlktNjl7daDqSh6hXAkUUgFgOeH+f6Y76FzokQH/+0Qsh3Qto1sHBeIC4g
xZZUnP2DG+CSwwD3ffi3dTGouJ7SZqNKjn1HA9P009Zr8K+AQRN7H3/UmmmJ
l0vBm8fBt0jADRkST9iB+clU/mYIXmdCfU52vnN01yX547eSVElpZtQID3gQ
u7xFnUQqcV/i32/JTw77Q+dygEIrmUrnPGTe+tYbEJ77jMf63IdDsbsmJKM2
cf4cVRn+BDqtNBC7F60FzMPOn7Q3v96U1QM8BW/7s8gX5iFEpBXpb/M+1sfK
5phMRVS6jvjiDHN4bQcEz8EkcfX6iKno0nbnrIJrnWJfJFSDcmAXcdxd+zAA
bs5MOG8DdR29ZuPc/YdvZ+nMz3C5+ZdrBehbrNSlrhqISgd+4KlR4kvPmpAd
l1qmbOlfPYpgwJYiIrlxC5atT4Jaq5MlqGsYKfDfB8fars7QVZjk70E7K2Xr
FyvdLR+TDEV9QbA8yr+Zy3Pd9k+NcZzWzoXJ3GLDIcui1APdih1wbw0+dvlW
BhMr90YghlS0j0m9LDDS3FvYDo5zjFLTk0cgfaZDTJnIcFa/OsnV9KRZ33Mr
mFJZbnG/YboAQ01eCmf/iyP7cSMSPkN3bA0jcoKIAJ/GiWyCi6MbNRUm4hGr
c0koYp616e9Mt9nkGNE861fX35QkTiPBfqUW3rJZeBLxrAmRyiI9sLboUMbV
QAWkQrbPQ/3eCS8ZBiKh8E+BmuMKgK71ILrwC/lpv3uiu250B0moZIoMy5OY
cWx2I9pCHLDaOlrSGJAxCOX+bn1YW/pEi4ZRmPaAAfCAdjZtK928EyZ1caY/
hG4OfR4feMY/pp2e2UTu5bzWydPpA2skceqNvqHiuXOuoCiH5Bo8R/LHpxZX
eql5TRnwPbigP0WnjVC6+/AQi9a+swNvMTDGdqxjlfn7yVI9xeIGu4FOtBWH
xMY8se8umoI/oO085Rt6G+kA9k1Hk+t0yziAiOgFzFsY7RD/sQ88+Q/Ac4tR
Yc+KLDCWMMbhpzBc6OgNQMVvTU0v1MwgWSn9O4vcX2DNqtheFZ0qY5iCbWtS
gMRPtDS0fe3EgEIYRsLd+bqacEOkhLEM2p+Na7TaCh+j3i1fd6x/Ps2vDeHE
ZxOYSwq9IbjNJZ5D48kIv6GQWTzjT4G1sHDEAfXhy2DPCgDCu6mz6Z4L91QJ
mj3x+WdkJsn4XU9rNxLHnypLDZXeYan3bpbYbCpev/mdllBitE2OSY5kyfAw
hQngjBwfb0TnSOQozlNmGOtG2BfEhgFD4KL3Tw1T9+JksNHh3Q7QbbiFWsO6
GwA0P9ihTMeirbrhFqK29TbTV21MtWmSsN8WQMeNTZvFqR905c3NciWo/Ujf
t6ETREnjbeCGsni/NNXCk//UBhm3Vi3qrdYwBj49RRlgXTqEQhy4rJ3XcYzl
qn/bxT+8LOW6Nij7Q1KWAlVgUcgly5GZlrkJdrJ27VYD5zojZMyLdvODPJdC
MldpXnlyV74Lm9O5J3vEZ1ZhTXhNlANm1069S6kKo6hoUzcNR9hKfpIHZLA5
ZJiF00OKbAGpe8XE91qBi7TQ1/Sjw195EW7AqPC71p73Vp56cNgIIPF9pEGJ
HJr2y8lIWxIqPI2nJWwalF3oP0kzU5PGtACZ0Qtcmwn70NH6FKL2yMbLO8Zj
29Khn+MxKlCIm2zUawKpDe/ru+VsH67hxg5jXbXMM9S9N01Mp8h+PCtCm8ya
J+Ppq061a7ItKTidj6mI3MjykZ22U6f6BIWva3QacKH+qgs1hZMfhWGq+yAh
4m7Bg6eFGGji53lA/QMJSXseIIQUBHwPuiOfp/rS6FMs9/DoRT1rdqQloNHG
vZzTu/6kCNrL1UnwWR2g2SBnyIXhg4NqKyob3mKzFhhVs7Tjm/iqiVFOjJPe
JqrnFIqE+Ceh4bNCOqPaO2k/zZ9vQwjv40RalUqEtIlv4CzIBYuVooj6tfMp
5FkWWxSTw66W4bYl4xEF8AQh1vJL3L+rAbzlqN32Wg7DBDp61xjxhFK+OJYI
Xx8Wc9SMcdRcjIQq5ZC8UbYDhOKH4lntXzV225DTqZWF4pbzbtlQ/QR++4Wz
LZdEsd2VOsar42d5zCFuaWUvnP5ojR1tYIJTLdkBcfXuPyDyg2iljPrSb8gr
YoKKYFtNcCvyT0p5P3huZY3n3Eo9+23VmLjL7x0L/YZTLehrt/ELVYM1bTz/
5+SdofLRX1OIUExr8iF0IWM+Io/F4uPrQwSn63RnHQn/xGF+bQfR2Rz7Deig
OlmsmgHf5zJmBOlvA377jJezt3Q/bd7vv9fJaZadzhRpqYE9NpYH4YYW1NbJ
plA9726xPHSGAHKZ1bxj3P7bdi6gROCJ53MHzhy/2+ZfztAxfgPNGRtdQ68v
ZURo6PfJRnIG7Z5s+mM3c6RhxZshTqF80V/1r0u1mhAlH92lyeLc7UXcgpRJ
IsLFObMX5ZUAf4ILoLmRGqUSeZLxgnlKcMExqUEFs0uyKo1xn3JrogdSR0IN
2Djj65n1oieyK/Q2kSUEevKlDpWoy1bbIh+87uT0B6FqPfMz48T/OJzPgDGy
ubjHgW6ax7rWFyqpLmBFNruhF/m4GDFxBkRCXgWc51232MFJ0uhGQ0OB3z0w
8QqdIXoATtyogjjALvKPST8W3fwCJtdLTmiCoURdL/5pQptNII2cVIjbrAPV
d91oLA3S1hwByMvfqhzTAEMll+ZwBbUzHywFdWXBUzj+FwWQenoVIC9xB5ar
M4TrRjFUhI82OuQaB+OyrweUkU0gOqNrdXCA/GSinlA6Yc8VYnDpvnS13JN8
ltCeAGnvslNM05BMVGDRxz4A9iqAuyUJCbJqDE/qitxRgid3sZGNrWBnIXJ4
XZ9qYEpjaGpoOZRU3nzi7YHtWKxT9A46nmxdhVlwkAvozLLfciBSFqiyy3rE
nfg8xDR/aWIsW3t/G+DTOzXxG9hnwOLRKiTOGWb8RNX6p6X/sa/0qkIe3+nv
6E4lxXglCSfbgpkFRvACVNAVWtl3fBNnkuAIEOwWvH+ic3A/i5zxLpWFHGBr
H4iLMwApIL/k7SW9PF2Vn7OcJasIyUZf9r2UIet1pA6CB7UFPvkpV+SJG5om
gTuDue40Q4rnUFk4LpCWKHvrLeCpypjLeB/pulNQyV4ALrxAG5w1kDakcKWT
YLkUm5oRUkhQbE8BWngm2Ob5HERfqti34cyVg1dGNphLivA0g0ZEkBwFTMpu
0SCxDwiBovUsxy5wKTVuupwv3YKKHpMysJARKAYZ5M6YMRp5m9Fy5UwhhP/S
caaak9EhFWwdeltIavaLA16O2U+k06n1yvwhJsSfq27GcpdIDxjZHVD/qNcI
/rv49n81odBn/vru+m9O3DM/950GRVn6LFKfIdOeubwj7skZGkGXa/c+ettb
cO6R76vOk+YyMKzWUG/TKHU7EZZAUKT1hgiTvtde3tc+zUnGPRJ0ftSgXZAU
RF9imKwL82/FrF7+syQlrYvSFfvHqYNhy1Ro4smsAkuSw5FIu15PNDH2mpBZ
DpVRJ0nEJJq2/3kMgJT291/mPvsSRzfMzKmJlrCzqLzaqqN/+XvNkQdGhCeF
SFdvFUARX/4nrgkVqXxG4XxouX8n9DXpeoHTmfpSA82j5u/wYKkykJCnHosE
JO0TzQQa1Osoqv1cOFa1fdNqYmqdPOtDTVnS0R8b0PS37vOPh9qTmAFoiwo/
BYP2Nvpyqb3iTmFLMd6gxYwJg1buRL7O8lilgbPmANrIsyCMFPFlFNXSG1mg
kg1uDa60N1lVX+HR6N1cvOqaQeAjFI7D/RmZj0/e1SUoLcIA49l+6PdGx0q3
ESpOP58pugT59TXU+q/TtrRd+qmAwPwZ1C7m0C7RuyED+U3fs1FysbJEu7nR
6r1HpyXuCC2M3PJ0JPt5UDrfQQvR51uyzmIWVYV58GnLkMbqrv6QHhTQ3gkv
7vRjJzYJfy67lgyxHLYxun8ANBBdvHBXhN+Wd0QqdRrLih5Iy1K7FAyN8f/B
gvxC+x2/vqaPtRhqbonHhPJTfjVEqSfqpWUcZ7E9omPlWkbmyG2p6jyPhTmL
5nmjKxHhokKbOTZaLyujtA6nymofdImPpDkYnS/APQvFBA54a8GeA2BOzPIR
4F8wfqyj0xvq51IpV2Kq28frbeMwAOE8nS/1xkHFNr1WW3paQl0mrthzJeWM
NXCzoOjlC6AL+EjYKpl3PcfcsRpgwFWLFHKHhkClfpqUXEaBZd6vMCHJj6uE
1Vy2KwMcZF1s9BrBfw9VWHspmqe5Bd9yiYA+uF0aww6VyiKzpBOCKkuKtvhu
i139n0Kb/aoYrsSOmwl+FVEnSJc3RdrGKtjfaCKs7M4LjkDZWfuLTuysxuWz
AZ8g5XNw2hv0NeIYmeEKNiK+2T+b7jg9NUBI1pkHglCRgO1pH/S7/+zLdPvK
ZdQ+vVIPaHdqKWpePwrS7zh4uYEhx7ouITx2DSi7nUnp658Mgr+PiSD5aopt
FhrW5GKAH/d22FYtjzc1HLw8KDTmH8hIC09NdT8a3sT1NjPp0QFQATLAdWzL
TG7SDVWyqe1TVtQKEPsBNodhPfHrHfEFpKg62/wDY78K2SvuK0P+3fhIYGdI
vE6X8pTUI+OzRbz0m4gCTCsHIr1RsETZZHzloAzRfFQmz48Bqviix7H/6nIB
tF4HYDVNyyGNz/3iq2TdRqTNL+EsBeTsPWoLX0ap/LHITbuzkqKefx6PpX6f
W5qX6j1JYiW57x9OKkRML1sVA8GT8zf/O5cV3VxaEwN+hvdjuOaHFjiz9mZn
RX018Dgw+DCUqe4de3TI61X3P49/hB3ZnasI2bti67JerKZWLKw9FqqVnT8D
OOwGCY98F722GYtECLEpkiaPUu9udcQzkNoL/K9orbX+hKFo7l8/U73krxRy
pSGvqVJn3vq72j5m30mVtecg/Lq6inR3uw2C7L5qOoANlOFcM1UxK+r83VOd
txouiAYyxIbP0Br9TQFPF/iAiGSYNdeZ/jwxItCyb0MknqChKmqeBJKz6xMD
H8PgFqBNHFXetdM/3XrikowO3dCaWWY3VujLJPQJrfARuGZpOZ326wkGMmnX
8uz1fyZnYeRWkO7ky4Zo/6qUxh8JUb6efx9H7Q0ls9IP3EzRJbvLFzs3ZQuf
PdNH9O6wMOJAqWVmzBxJ/vFcR0hx/pDCjcBzcQ6WvjArNpKkLosANrBAlx/8
jAI+NQtqWSNB2i1Qj5cevUJ4LgEhXn4oPDMWvD8nfNyfsXAagGGOgtpcsWGA
dsD5UPGeEpkQyMn36Nc7B6D/RApxk8/M2qNp5IDQ/mIgQOhX0Y/MQBnVYvJA
FzPhcq8DNOYfOwjj4a4ZAujjugSPMdGZxNQXC8TYDiGmVe8DtgoSifxLsoO7
S3/RrOCUR9dGhnpnGiy812QmOMjACYlTSnjeZZCbiWa5Mi6O2TrFiP+IN2g2
50DZXOHFLnKhezN5ieN8bHLed/oeqXzu0ddOBhecnGJf4k7WJXxUTXRJR/O6
tZb/eph+OhIzWA/G5rjb0MPn9cxJjaT7blk+7DUYiX2nI+tSEjQe37s297zS
RXuOOhJQaoF+332GaM6DRfOyB0CDWaRUyZpXSnMUL+cuZSeqXhr23oulYtD5
WE9pZNmOlckqx7Wb9IF9mkD2vrJBZ/pcuZ4b0SNgR3zoZ1s2iI98C1m+dtEx
gZ3el0ScaUSjDfi9PSc+gV8yjdIfHArOTmuAgwGu+KKGNqBMeN+CcKp5Y3uf
3W+vEuj8BZPUDg6TpOzYcxCiFEJAVLR7dzliA3CfmEKcsBPWvdWClFOCThFG
5VPpLSmx81YZmbpv1zCvVK2Kf/BzmFHz2D3savX+SpJAGhfbDPmp6y5TwfFg
PJcanJ0p/PRTnEBBVEUeZeXWTZ8mif41qiviSAcHImURvS1m+PLd6Mii1Zcv
wVSQpb1W/MPNtyHZ5U3PgZ4/5iyp87oCBuqyRQGQvE2yAF7FK3kyF5i3S6Dx
bjngMZpNH2pmIRkLnp+rBcflI6UoqW3SAuupuB31UZ6CGgrL6UwsJ8XHo3Ry
Ortw8CJD8GPzLk1Oi9cesHqZT8wNqguwO8LkfCFGAJpZdi4FbD6PrkWpf9iV
24iYzGzBMlNaEJTDEZV0CGbwldGUH1Ok98rvGkOOQYy9CiIL+x3ZR8mkawmV
i+uaDiZ0l0slRulVsbU84P5NdtU1xnxITrHRMRgmk0LBPXRLqa50OaocuUG7
mRU/OItHSti6WTms5gkG2+js4jKyIrKgbLy9ScTO1D2VYqeCsJqUkyLAVUxc
vWf9Uch+u2Va9uS7oaf49P+p5StPCSeAPR2khSfh+w4T+wROL7VjzJ+kLNXA
OxsndtQ1clcJqqv1K5SJtpGyMI/S/P+7yjEnmkc8tecpxZ9Y3Y0ve5PXY9Fj
7NuuU6m0DYEMXIlbNqUuerZKsvbIdevJr9bYSswM0KH0nehwA/S/Vs5vm/t8
mmN42KBp6LiTL1hHNvzd8nHVCzlJPW4DPGaNwO28k7oqmknygUnhO7sN/wh2
kw+u/pdYtJ9fYBUplF9Bo6l3C26vOKZdXfIzSgoFLEG6CMHumftj9m2JvbHJ
1ymwoHL2+4yx3skCO6VVNecmP539vSfKW52hB+LXGXY0AFrLAiGMbj7p7o83
e1eMuFqaaZD185BWAsg0/5xXpYwQlj8ylbtj4wy8nLOVtL4RbcMBpxKaUlzr
3XgPcQ/t2qW7xupkv63LEAqChUPV+w/AagJe8BiQNYqmT/KdvK82C375t9TD
Y8fb8g5+aWWllXbv5YaxfO+V5cmNCoGnwWMPdqfvncZgkD0AazmvVw0pfxzG
WMFy3yKbZLx8YtR82c/hmfMZ1PKfrl77+zB5SzpC/FwatpVWUVu+iZvnmmXS
oHng60Yi22jiVeGfapUHr5OS92snQ2xHO8DwYyHTx22CczocXBSCvNxjHJ/C
43G/ZkTQPpSoA7DQyFRIuMNdvttuPX9DvLAEcN/Fsz7xN6Xw1giP+hgYg1HR
ErY+zXEDQLPc8BV8Kc16Xx3S0KV5jnnhhzpyaQeE4L8PzwxYQKhY+4OOBGYg
4aXd4SqzWpieZV73bbMMTd8tNRGtqpxKAF51s6aZ3tNMqkvWnGn+mOJAo2IC
JW28y2pE6Wkuw3pcCIrtJDF88ticixqAq97vh3S0hynvwdUJPkb0H/dKgGXw
BZyRqSMPgGyLacyNFDw00sPvWcBJvv6c/DC+GKRSMnPQfXzSXPf146DVRU0l
4W1Om32MymhaCZdgToyJ4/T+n7FJlZbZdRPj1pIPBhKty5nzVPIbOqbM7VHU
RMMPnT5euiuPbYk0Nzs0MaFIJzD3P+AsQjysWrCB5u1LEd8Lz9D/CyX+q2Ts
HBrltaJ90eizp21mUxPjq6sDnvEi2XmJpHX70ocYDXfV/Hw0z5bXHOgLmzUF
PDdPHdthXOqa3nbQPsm1FUw0lPj2DU/BymM6iq9xu70IRq7CsD+zCIoV4BDB
f6uur3Gh4BLCiClg23hWCjgMpjZP7HjoLnuMEpmI9AY9uZH0i14Td7mHRnQR
FTpaWNjVxfqg7YEKJz93m6Q1guAeyQFly6u4QwsOqDyNIe+QU9yK5nwDN/a7
Oihgee6x3hlFZ3pjxTCI/alFmySvK8Q5yBjbTW30l8SjwjE5Do5p1YJEwdBC
vsTmOOdhAa5lD1RjorEzAmjJtQwnrTMZTSFtYBlHVOXfnPCnHuBnwDsGwqFn
kxBw1ihJVpoxe7z/5EPbePbhIpWEtnV9TfBkiMVejXCpaHRBhSGDsjnM8WM4
CGn49EF4ODPWK+jf/R0ss5ODQdt4VpUjSmmHhzrCKppody4m3tHKMutear1E
M2Uc+j/QRe0V8PBUGxT4NE6de+lvXs9tbLCQkLXZIv6kxYAhOACAjHrjrGLt
bZZ9RVo0JEVO1lF2Pvj6c+hSPtRnqHjXRAXIpo1JOLEvdye1XmEfgBu/TrQM
+UGlMFeAYebZM0tic0nYmw/yM34UqndHNr0p9oJw6Bgn10a2bEVHbN8Sj/Ik
uoS1xXOKJtsdVtUNjbhykto20KX/FmxLrQdECIjcqbCDcXzvvreQ32e249F9
RtYjFNwaNnsxmAtoCiWfhtsfeMnoJPCZIbL7jZe7CJ7zoxE5NEjbAeeIV8qw
a3nb7Ia49iPUDijvZk/QE2mUPfFjSD3S6se0ViJ0GTyWQ/qSNh/GWymAfznC
d/CgtJoQUoxalAFav8a0g90q3YHMSxIQRDpqezyh95jGSfcBQoOHGirc57qZ
U9O7MHKoTkDkFDxIxnXKJO3iGmtNqJ4SQO4B8DT+GcyVnz/iHrwdz183mVqv
/FB5CmQEzqs73DL5RFEMmpAfQo7sCcUWHE51d9Wnl+YAxbNG1NdWeLbHHT+3
eYnn9WpH5Oak4jiPENaiL0tGJefFg4t4aeHqPJnlqcmQIq+0/d2hrEkklA9i
PyA2XHafBc2jTf6YecAZK3Dd4tpBCiZ6Gq6VoIZ5pS8XnVUCczb/UhNQ5eWf
ydQVJWRSnk5hjKeQkMxxaKX5nzo3OcRggtZDa566Kl4gXDiHkfKqglLrBHYy
KOMsg4v6mTaOsJRN4HiARsd8J51HuuZ69KcL5BEW90OssQvB6tfa48IHeEzW
Jx2HbGmPcTZUvCHJf5qPJdxbb0qbfYGxTzhwCcwtYsuQTzMHi5HddrQqVSeT
t6lYES0LEYAacF+rAb0uzsJepNr0aNFhe3lvMItLO89T7bh/6MZPIbZfbScV
VYGYbFWQYEB44PdXM/Mtu0l3PD91KKSJLPAzbmwrD0riIWaUB6RedR/Ha97d
ZmanUOg11+nGEvP5Qs42nar7svhNRrqBRoc4A6f9X7jLzOR0PHw4sID8tMta
3TqkHbtsZsMB49I75MQfK7QLZYFxsCcWa4aECZLfQmsFvf/PBHQS1m90PWfQ
drheG49oV3MajIgb6kQnnTxlJZHf7rza9yuCkdvDiMdT6CjXw4zHk77KD7Is
NDoEweNaTmGaS8N6kF2L+sp8/pR+Xf9tJGAAihcGxqKMRhELf7pBqv6WAMpn
gaw9U38IZW+7zV8tCo/KKSm1nVh8mdCL/Xd04tQl7+KaRfEzh7NAGMJL0DxC
CKjiLgzBco0vbXFa9OrjKVFgvELKKCRv3eQov8vRESWFHXtgu2/ipQ/F+ljX
Pw9FtoLff0B6mlxQGLD71954XYn2WNvvDt4E/6D3SgrLkayElcqHvHQV0j5x
SjbtUo8KL1kkQIbC/mP3sN5c25/7yZdZ09R4aXE34xIm/Prle+F22Jd4a0GX
2xNrPUXol2IMS5hMa8NTvL+53PrQdXd6D3awQsOqLByy4yxmTIG721CW7xEf
/SeJ0dsC1Q/b6W84pu298iF01eldq1Rv4IVPn5yIOvVrkB4qqSjljeFMAOVl
9N+W10ZHkoREhbZmN0TqD2VGHAYHjBEYeFeshyQxsxlWSATb9bx18Pl34DNT
S5HucA0w6LzrGhIVtp7N6xOKL5zDAjkpOORsgeBt0xC5pVfzUY7fbfLI12yI
786Km9ZB0eu5oYMAysg6rb69V0ZIC+6pczV8S1712re/pxfreKMXA8AK+dPz
EIN7BzwYHq1On+R9KHXBpM/LC607X1OdinD7bHRAzW+AtRDPIQErDn4F8pEB
nJFJSeCWZiY5w2VmnBqlKldFt8lag1IC1lMpGTTJn5xp1dg7IxoPegOfxNi/
5L0rgnvxpu8zuKhMxLqit/490QJVBq+NMvBmMi4Qiv4K2aJfd4fQt8wSFypZ
Teo36yWy4BpQqkgihk9TmqDKuXoGvU28Twe41YaM04Ze/eM8BYdZYhzWh6Fi
RFaFwpLyuwoxIkaVDEejAIYuW0XaMZeqph/8XRNCE5meTyaVNo46lob59lqb
RxEnicjHK86CxlfSZ33rzPyE4DfhYqsADmhGPmlNuJiwe5U2SRPtiMtkwgW3
EcwbyJDgLQFUE2fek5T101JXJSVVZh80GkBvpk3STmJiaslaetSESD5XjOxf
wCgeCW64DKhbX6qp2kcR7iYyaEA32AfN1mJsz0sRFKnM+ftQATbYBkJo9Tdl
P1boRxdAXeUlUjjZTOeIKSdVTrYzW1XQqLKu0qwHF6u75lJO1uHXF+v7Zg8Q
pcY1kO/LVHgsiMMlVjLcA/cQfabbIovTwYq2f5krbZw0TaOy3Hayj8vjFdiL
+SQrHwznaUWcO+TRvIDhrajozecJwCumgZAekkyaYvx/ZyVoYx06IvNHxyoo
bNfSXLHk2uZkIRXvJMLz5yg5UWhvw85Pd2Ohup425O/k2FZ2R4vY4kDQTjF0
af5bGldhEjZgNNYp8KWObrcYcVAnPvOvlYqiS+LWBmw8Lv0+8GqaEhoZKa4P
6oqnnDBam5DG3meMbABDyLuieWe6WhU4P5lmRKesedKY1DYuxEH55e9CbtDr
tamxaoNvTICn0SShcYfK4xMF7FG2zQpT0ux3CL7qDarN7nLpcuTwlKk95fg2
WqfgSwZ2yPK4QQz4MbfwVSIuPntRqGZixzzZtm5KdP10chKv3vUfOSBsHxAe
AMyLJ6I32V+P+q6X4zw6nLRrx6D17xlJAPpe7Is7F06kS5ThKsAsOMrDtTFW
8o7nK1hsnkXDi1EUVMdyzHEzHYGyTQgzgZn5FgNHheYYRbbG3G1f0mlvWt2u
iwhe/lWs0o0AxWpyXa/XHnQXRezL1uSYG1C2WkBTuPBr1+dX1ldUns1/L6oZ
9pnKutFQK2rvGyloYwpG1wSnCpJHRsqJm1eGsv5Qq/kbnKSxNsAP4/QL0V3t
hGBxBQBJh+rIwfJX2GbKrtXPkbAia948QWhOl74DRncFq2PAkJ1JmTv8Dwt7
hh5lLgG/tSqiBjlLODAQImouhApcHihZqH0I9u7g7ixpaL808Puw4jQ0EYhK
hTtnGG9dGUGUqlYhyy8Ii2YW3UpKtDMLYkdyIjwNyQlHj7GK5po4HVqZoy5a
Ot8nAvIgF/1oa8Phef98+B0v3vkTAyEWTFRQoInZg2klqV51BWSErhzGtVOr
/Kct4iefMGQOPC2L9rKv3FXtr+8HMhOkM4dmwZ0TN3G4k15SsAJHDreLDQRy
S6+2dOS8vkTk/hz4LucDygS3FHdzSL/kqpxux0C7fJ/EAcBGE5qSa08cvtkQ
G/voAIf6+GaTwNisS3/oS6PU1RZVHulW8nhMn7g3+2/sAWf47xXYYrrybwID
GghmvRysLLnwb3GNGgoKNqr8oxtuOneW9CFpkx7IbpzyOkL5+WyWsrRfKenS
obADkx0dduKSxlkOZKFsLh1CWS4XtBHS1iCj+DJnsvZz/cLXxfU8zmZf9nen
pPzUVaj/v7+TT5OWELA9XCsv/dfr0xdPJc9LmOWfsBIsahPXvxGDhJ+oxeSU
qxXEVphZ0mCvviHcccaAYLsWxqaa4/xTEFFrBd2S5tGmZkeF/OsTAL/v+EgO
xvCpOdoTwdq+0jS/ktiLXTCueK7Iv1kDIyxpjiBBr99TYDRNOeN8dVY7E+E5
R8awFPS17G2A18Dz1TUAUDDJ8Bmz4bdhMFnwwpZAo8gt0KMHSmMnetvQIXQD
h9MYGBwX0sSrSKNntF4VQGlmi/prCVRq2dgdrDDwA1QWdu39/4d+U3B7CUUP
1cTuOHTrVKS6Kz74x0mcQ4cjq+StGgpblfSCaoGYq3x+CyyDBlgplCNScMIL
3n0Xj2BKE0U0o3JpNMvSb6vzco43yxtH/OAMilJhdHyHek0CTFUhk3/vX1QO
cWQlp0LlVDEnxqYfeX6BUqqPPaV222f0dHE/ugYSi10QKUIt9fq1g7/USXYo
mBKAC1m7//nxpa2HFxEKuGffu+56CgTu4d41SR4cgvVRE4T/odWWK3SIy7qq
jDTzLjvlLek0NUGy0vSnFRIatf2RBbBxONtjQQ5BiqQuD6/XzVYakP5H468Z
p7h0MbWoXA6mj1xXl/N18ZuSOP4pJ12uOvuGyrRdEgIEZGk1OF9qOZ7x8vZ7
7Gx7gQ7U08tHPO69lgrN2T7vfyUioEiGFdyAQhP1ZQ9kKxGlepujBNKSOEC9
017wV/dLXYQa/01COrmdSB2etNnh8zXG1aud/Nlyd0s3mQ665EmQ19JWuvI2
tBszq9oiuHgOIgefQb1nq7elB/ZjxynTMyVZDJJqNaLDCYkq80+uQGMgx8ua
lzfuahRTEbG/60Fn28nRXROLzKlT+k0tM1cDXDAFhYg6bp+5tSeAOYOhcJkG
R9e6IuyoWGbmCsg0YYxneN8S4eRBmEep6gN0Q56xIEdEE0Jd2E2+F7g04bp6
2CDO46evJPY2RwJ1pw8/C5Ok8Le2VeF/a9i3L2ggPShoQ/v6t3Yuc1E2LCQZ
dyvDc9P1NmS9+OwWTNP3FtGAGOfWgbwTSTC84WE0fX1Qm6a3d+vdaWFVtIDC
N7qZryPswXWR8MEDwlB1LyM7AfmmHDOwDx8100kjclXET8kemyZSG1TousHX
DcULx23dzQGhrlvLWBXw4X/ZkpaSaxhL3Kr//5KnHn2zochmDlzxeZRZZHyH
TjpOH7tamMzb6gwowCg652iPAsAv1nx1xzRINF4Qk5c3oq0agLBPqbg/K37h
ba98Hey/hKcLa7SXrZySecy68IfaH0p3grcPtIn/UMiN8ds3GDkg8EqxmQd+
RfE+/gEUP5W4eSY8KPbRb0AlWMQtn5pGG13YhWhBB5WXt1NfYmTjOpTCbmEl
N/fbExO9ewTGytXmsU/shuSozW60VhYqiXupwqWb+kZSjw/L0N4O3BDK+f+H
LZGhypB7/Baae72RYQ/2Nq/7Q/+7SfsM3/y8W59BnrIKJFyKJ+9qv0lfRwc4
iGhvv3Yx3MeM8M29vP3Rs85KBv8BbZaJCkTODu0oLA4Go3j9iLSrkQDsZfPy
9Y//kndGFakA+A7fZVt4cPgQ9UcDSpMt+4MvrNFUwiL1ByPHv5RRG9BFrPtx
Skp9Wxk7jPZwXYf2OoS/qbqvAzNte8I1HoQ13ZeS77jRTp+/w/4/29gSMHmx
XM2BUE0xQkhhteyI/YE/DObeTUDYZlkJUwRLyQsc2q/xdHbgJRN351AY3kiT
u+pOKciybQzKqxikYxyEbkxIDXPRJpyWhiffyFjdRMYhgAGGqngvcY83Gx5f
m+B/AujuGciQJhJSa5zD7SgG3Vo2qYRm0whhFcH7o2eOF2hxD9o7V3vTK4l7
77CtXjneCjpK8xqGC8CjKCpOt6KDPVDWN037aULSt74PDaOVd+5RtjgHA+T9
6jjYS8oE4sfw16fhCBHzIdNBQCIKYKW7HeWfmWHAh/Dl+dsKSlZFVc/4auiN
84PYrfdslmVGGgWqg/uk7xbNC/64Vn4C+LYg/fS8tu3m8gox7ujnPX6DQDqM
g0UGqEyq03OE/ZHllEbnl1RqgryyTLBGIVYCXR7CS6jfouNvzwjXyAT6pq+l
LlWVfKLcwVgbN04fg/I3R4w+gcDu8PSVvt3hCLgAoQELO7SJjRNjKJSKmEw3
a9zn01Ezh+1gCcMnWvRVq4anr56dfC28Wzfjs+BoOdAjyTeZQxW2AQyxlP9s
660HgVvlHxnJqS893ykVmMSHGs6gTeurmY1YQvpRdck1YO41advYeugbQOU7
MZODtSNcaRlYg1KUg735YsHsRVoOVgtuKLdKr5wPOIAopnVn2dRpgl/F+ywO
j0ECF8zO6hcfCn2AJFh0dOLvUOBMi3W94zuAtt8YhEBJjwxFkzxD3WeYvxAy
5cQTv+TXmSjNbR+2Ds9aDvQRd+gyJbLpfEZriVGbUh+mDyeIJA6GDDAOakEJ
KCMU+/PziDDWABox7ga7WzcgeOj92cGu8Rh8A18l7Kk9bSYBO2x9rcJpTrVz
oxfu7+pL4emvDRIV/7rhMdSNZ7qY+C2ZawdSTN97fLyThe1wzc7i5lcSMr6Q
DYqh2QKgoZVASQ9wjroqPi3qIEz2k6SClXA4yCScsjdTpJSAEGWSAZW395ax
4Y5xDdeOPytiEmrTjhovGu2mq0OFHmsOIcnvm0X1XFtCJHZwgmwnmZxwG6jE
3VkTFcCymXGwlExNmFEBeM2Z7hHlQALnXO1UXwwA2D3zuUbwF6glki4nQD/y
2YpaWag7ARZbMp6dhZjBh/TSCpMqAs0gqEsxRHzPORWckJt+eX8S4IqlLSkx
r3oo0IC6GHwhIG0XfU+SjpcrfdicSpl/VVZj6SzfwIL75wo9XlyG3CfchaF2
YecbuSiWdIJ4WLU8YtLLulXAomCK8ZBFdL/4OCz4nmg+xmkQE/RgCw3l8jaG
OhsGUGPr55DcbE2rp9Y3ZBGxSfVRnAF/iamTLyuU2JpDfp9PolzKPyLm7iwx
2H6NkQWThSfR7+49sq/cv3bVzbomdA6o6qxbU/M8E+EG3ur0xB4ENpomhUy5
07wuzcmio0Onh7nA54LFBNXIVuofWGf0KXMmshDGPMD4TqfqIxCCtH4et3I4
t6NbM2sjqykA7gkt5pRKtR/YrxclyWM9PO0ZQZRepTsiQevP5Es9IFXkxRHo
1m7FejVeMktEgFePd60Ya8+YGJ48kEKBVRwE9TVDlAHed2JN5lxkAiho9fBT
J34IrvxtTYrzKEdugXj4l773LjtA4RPvpEe/WW00voUlY1VAy8u3C1Fsc8kk
Q1Y5N3drWL185w7I9iknnCT3m+Q3YkfLvWmgZp35z8ECrlPRo7HMKz9q2DDg
YCV6z+hxNgjmHK7eOgFQM1NHdzXtcLBBuM6cU+4RhDCrSa0RSKGm1KsOukDV
S5CDxeW9MhHDnXzJUCuiLBcg9XJWfsXhXnypLacnmfs22Z+SPrEATrBXbabX
B0/TnnsZ8QRBVt/n9gdDXJKnbJ+DRwkVa/MHCdiAZAP5Wc5pZFlOSDQ7NdFO
oS9TjW0Bg8FkMXQOJ9vQEAQTJWAgGCeydUsiImEni7Py8Vyxd6q7byFpWN6j
zQ2IPVyvQA9Wp31i3vPdBShsGwfwm8uXYt3t8rXCJPYiHtD8unuIvgyKg+Ca
+XltSeJyrkFAbM+lVpw5W8V/9HQkqd7N8z6joeo7UQNNPpKYadTTZtAws4V3
5ltGYaLW4T9R/RDIbtfcOumYo2a1YZihPC9tv8VAmu56N7l/uvc+zQOXzNVG
RazYsF8572k3rO+cWlBqjNQI5vg1O1dE7yUJM4QfkJvbSlMoN+Gs/IQcZ4FD
xh5ziYiJ2sbVmheyBRUiQd0zBwfLyyuNsFozRBMSnFNBkGmgTcVg6fLQcT8B
ELdnMIyWb2Rhpvt9UJYd0XfNqEvlrRSmik+wuCRPUp3x0di2wbgfOwlR1/NV
7CAzT0Pmc2StNKwwoXMzN9jKjJPYeOiZymSVg1vxrt02tZwDVB7effaJ9emQ
jLuUWtW3MBAP50IH91+mBdeULlacBk1AQTJ5F/iZyC+HaEK5NsHTvKFLjppf
9fsYpNmkLnYn0biAseKvmuvNujkAzmsedbXHUfIMxeexv0aufGHJ0RJeYDMg
ZkDjP5nwm+fektngm3Mbm31wWKI43I5AEyQb/Lq/lZjFD10gORTM+jPKzjcf
HJerv5zkHXS6VBhmLLtSnmz4CIevKlcElDPvsfSERyWctILJfga+1aZXXUKG
qtl3GinfrL6VVkblas/AqL0yl8wgj6KKi408iEM9XMR88lbZuTZUKEJ1RwVx
PTVChZNU8ohWQ5kbg/YwXzCX+pYMlnqNDGiZJ9usQ+t4gW8kq1l43lGqLjkZ
H0lwLWrJQI/CLZKGX19646SBchgw9ZEuYfxjPQUM+x8X0QjvauE+QM+s+uwY
xOsGvzMqMW1ClDF3cqrKVoKobqWhftOxF1Wfoh2h687cyP+rSqIbe+lYAzNH
aosIsvmaNV5ViuIZn1Sx4CAfVpWPDs/wcogf10FkNIn5a+2ECOY6gF0EVa5Q
N3eQwnN8UxjUbshKg9Ig+NIt9DRVabkMhByeYIl1vOssPJxnKkPBnaBFD6PD
E192QHnNzu/cNSyvK7Q8fodKZyEheHRQ7g+N8PxpwU666GrykbMheefGzCuA
tMYf5rXBx0jiVA6jtr8j/9+xdYw9DoXyWHP8FKubUSKSizyiwm+/LtpQVx0T
HjeEBvop8XWhlphpqPxhtRU+o5mwJ/wWByLnh2uVWXQlgPRqufopTfwD5MDJ
EzF4dlID9g3+5ev1BQPZ+y4chFx67aV5aL96Qhy7Bldciol4DQF+YokrMdML
nJxPbLjcA/QimptoVND7MeA5H32xfPYzLgFVRbcD8ohZtF2jp26sO0Mym4My
EGAWecovw/8GOQQxdXD80npaHTC4LToh4CBpYdeOm49OEPMBDKxIwDow1cuL
YoOjJvwZx0jy4hmJNicB6H81voDNJo8WIrFK73Xo32x2jpB0OVEmxBshPRof
Gyck5NxUDFiMzHz7+iF9qh7Edx1to2t3V3ocS9BoqVK78qjhLrr8uD1VpBUW
R7IiDxgglZDWoguYNlY1KheZIRpYAWWg2gJ25EK3JcHEvo15hHo9Ru9VQAve
2WZg1jKmmObS0hFKeLCv680Ax7XNz5CdvdOfVwXsAayJSW2WTmw+Lny7+oo0
x/DaXlEiVpfdFHc+DO4LaI4P7npc5MPXkZAzU1LVoOzRYpKeJdTp79Rh55Mb
hADzTFqOEsgeru8UVfmZGIHuELcIokQ8a3TJ6jB4APdkwUe3sggpPbc8DEdr
CzcXCbBFprkIooPwDSnLSo95VKNjkJzNlQwhvyRbydjg25GzCAAJVl9GnUXk
7B1lAJ7dkbW6wPXRobWSPUQtFFcQ02fo7hCGyxtYbmuZjfwDCg6Wdju2flmJ
QkiYMlqwROe1srus/cGwTYASOISPZh+WtKJj9VnQ460Hajqi34qLWdZFwXvb
ZVY7K6Ww0MkEMpoZ+UG0wg6V3j5GfZh5J6GFIsLAzL990T8Bxr+A+CcExiQk
83Ss52Tp/3e6kPd0C5kVdAGwNWm/FN9adyaGAsGcLNp4adkExyeXxUggHW2t
+EInGsjqEC5pqZKzU3G5r/xy3wNCYDsB/x4/fArtBLUgoaWzIkxfANL028dp
yYJrqloh2yH5+EZrA8umhE3NQAabuVD8KM2sB4LZtuUfNyKlToA3AB/NQ3RN
pHLkHz7WMjoZnR7+3YmprPCnrBmtLlcX2ZxWgmlY7pxbmMM3AnBfZSml3NsF
PvkUnlRKxZQp2MkwyDRURnALKmgZsLgvo7ZHlwCJinn4wnnUeW7Zpyf3qrKZ
ZyAH9z2380KRFLBr1iy58y7PtmYEcMfhF0BZCUcE0wHrvEkrfkXACWAVh8JE
/uasFjUAf23W+aAMdebfruzh3XhLKMQ9InrJU1ep02T0ghAwCZNmxC0zxMGs
dENoQKu0XwOYF3HPGXvpyw3zla+yE1kb5/KrX78aKmB0FcCtmRWBWE4Qh1Z6
hd1ld1cdWsg+n4mdfEs/Rz8MXRFq5Xv57W2IgdSwrCVxQzMkVvv3dB6wob+d
TuU0FcE78oUQjFW5idXl0plrTGSMX5g6b1hyFEy7yxFHEWX03Aa48eh0u35X
5uHbTf3z0b7M6xodORtAghTkanqxmjsPa2ym6NkjjEpi+us8Ui3aAYhzL4jK
CD2PWkcFLPMEstgFftg52wnAg7uT8q3Ymlu0h1m1Ly+MzTa/iIqhFOg2oT/J
H8SL2wa5eEm9FNDgkZp4ibTQaySDtxtOXryzweRuW6r+7mX1mhuf5Pu+7d6i
3KgUc5xNSurWzVxHDK6GTOIVD3au2nKOw8TnaQtvimdoa2k4rBLm3hNewVqw
TqIPp4xLr7s3L1dByrbyP5iyThcEYJAgGy+xOyxad0O26U/+aVZdv+/cVxkB
ZjXIXzh/oElXYKujOI9V2ram829HCtqNtDs4C/HYhmIcqTUyOe7uy8v4te7y
YaQAicmBfBNIDZAwpQBNH90Y2Gu4IR5n6CBo+ce/gCmuBR9scJd/3eJgDL/9
H1C70qeKGwNmviNBdTp91oZ5XKbqVMpgUNKvxToGJMPNwrEnQdOpvsdu6CNi
aUP7mpM7R3GWdN1oNTI2yBWA9uABtsQ/SA/LZgm2qRVVA37+ptGHDHc92uoI
rH3pUtr5n5Qd4AOhou2UYOJiuAe2d3N0fZj6TrNccpEjb8mtyrFPnjkMizln
rwYuowfrsJH7GQQiOrbdzeB2ajBOVTpAwcVhi6D3PaDu0nx/jSio0zbd7ZB/
8ZbAp8O86Aqt4TpE8BpdZul5ERE8+QlPDGiliYjA7yz+lzw7remz1RHd5TLl
FxB3Bey/k9qXEM/ALpuq/WtagnEvCDDazlbL3uN1RJsI2heG7K6v9Op0HYxO
N1Ok+mjd7ha9CYHx7dsnbbJ1spCgaLl5QVWHwDvcSdvrq2MyAwrq/qb+iqyG
cBEqrrGEQfEo60U/ES/AdNSgkNZnTCYtkDMnjZe2WeHDjbIAzsq+w4DAsmh9
ncBwKS6G3xJaaWxQtgYBNuicVcBtI+DdXoL4eBGet8sM+GdxghpkzufbgID7
A/PO412IC2lCYG5uxXlnLmi2OZ6gUZOuPg9IVDE4vLlPwydphBlkrP7UnGu2
Qzg5cDgCUGXyNr1+flLp3lm3GdOV+jP2S4Sp+3tMvizW/t5dVt+Y7nomcWp3
7dVKIxxLgFrJxOjoRwFbVudwZfpCc0mI37xAMoP8LlhFCHzw3ISaDo9XPepd
UtjO69cIZDB19eR6ILDFeFIEEC6ujHAvvPH0hNZ07S5H1jw2BCENQ7do0SBV
MX3nAsS2K5Od+CPZ2HEcENTSVgaAhrnJyjS3EC+K/ndP2aCpLts5FFKvVk+S
/KyneSklycPxZulLtm7qBtpWjfeks8OMWocygNYfqc7fteq/ox7d6cvMpgZ+
RY2KJDGNsoenQL3siLyQQjbbxuOLowee8i+LQFM9Feq/R1CkzI63tOM6hbE8
aD7P+3zFPdLD++BMlAg9O/8fx637emjTbNUI8b9Ac2jfBFrOnbM81QyPmUAK
gyAXrdJ8LbsrH86Ijr0/Zy3dVFnEB8i3DIDVnSft+pALCeIdRfoJiwJrM29d
OFHLecWQfqYWdZr012466AeVsBqGY6gsWLS49Vxo+yWCBaZLDmW+U6zYaLlN
GlAS8TRrvATev0q3//LivZx4Y3Au1NHkUraWWLYi4MZyWczrqCjMaNVBnc4u
cOzvW4IRuC7E8ZyKFCPfmizaUj533S0L8HbOsdIHZ0RfZOZzwxQrubnLZ8XP
TgHXXd3U6EKO9SXfVB0GtH3fMaSD40r9WRRg+gyObjk7fdngEGIIVwmETwAd
GVfOWoxLu1pfloxPZsx+mICu5byrzbhVzskTDZf/BuGk9cEoWaCtfl6+kt4E
dMD4mljD0VDLUI2dUdqcsI2M43PaMJ3oqYSGkVWsGwb/p5gKBexVRqMI2+oU
7rDbFo1krHgbCn07mVzqSw4kSZhdyWk/MelKVv8rvnhXU+wbFFrBdsI9ciH7
YKxDDbyBlNaCSznLpQh8lq4/wD0BE2oxN/wLLpVz18ONreUfXYdz270yaKX6
20E+DjR/qRpC3No3D6ng5P5UDb5t28xn9nZTCCwkqrLJt4rgPWq09dXMqUaJ
aa5U12Aybwky2tRmTQy3irgycYhiRTTkAab3ITwMSyhDeDWposaGAkhX7qGe
hPf2lHbWnu0Q5FZZmvY5sA/KMpiy2jx9gzdREcdT7EYbvZfFqA+oXfYACTaa
VdnQ1X45Xy5C7Mrbv2Ab1Ssf4kDKSLZClHrHspiR16L6buhA6SX40rjoNywG
GwwvvO6+6ijRVKd9MrTT5d2LY6LChHNLabpDiAuvzUHQjPs2TaUJ5/yc7EUf
vQtOZxeM0jaNYiFOfV31f+xw99KSLXAa9s4999lDZUOOdUmDewM3IJDwEwKR
4kkOu0hBDevsA9ufgv3+R/IMH7Ao2ZDiZJBo7f2D261CBVbZsYIdnd/xIkSO
YboftkpAoUDAfKevah3Gtc/FmCTWU7ul/aBsTiI6KOtjCOs2zcukdNpzW324
uKmFpdF0lCDh6zLy5xMEwaKHQlX7LipiJw3kxb7MdHeKA7iZAbF9vC3CP2pu
08+ZNIY5hKuc57rV6OH5aiClEMCimD1FtL1JXW8pOt1fUtNY7UvY/cnqOoad
hKDrIqyrWrVxHlq2cskGEJFLTYmRgb5DVpjhgq3zxYim66a08jOq8vuxFT/H
hS55WzBHKKk2e0yFJkhuuQIXqYBxQPjccz3MpEkadQSxfFRECg2YRLSdTw1v
VMKR56DLC+7Z9sxlbV2vnFnfJKn4Zi0GkTnBnzm1JF43MYFPI5ldaRznt2dz
eJ+dD1f6pUgVYxPvf05GzHpxnQADU41bPugZXHBcpjDjCyhTw49XR/e/MlZE
//fuWePDg1chQq19KPLsd2kGl4unSZ9l14c896YZR99qaB7QJpBrqDQIYZ5t
2PJNdV2d5SxQc/Fu6Ze7xFxUzIbGMb2uLwyV/MAmP9RNmHvnuVAWoatKS+jt
CWps4wjqSP2PUSU3LV26k4TLAhqt0J24iVzaf6yArLcrZvAdX8EpWHgzjY3E
+ACAOBzbDWQdIxR6gIpH5/cFg9Kojl4MdZp3hWiSch80+/Bi4u/hj06nzzmh
5l5OfgPTW0oCsRFBhjTfY/yIO+psMIIF2TdVyudDO7o6x85W2MZYZ9f1WMeL
5YC+LwHX3ipPsaEHhELX7HUPUzYAAsoXZkboKyB7y+eVP97Xnj239J9hSjrR
cIbuGyvgRMxT+lk+c8lkky3hDxppW95pbg3Hib+gj8aNi1f+2RlUqqlopII4
i7BJdL5th5uKFeOW19it8XPiYzLKUw+pJ3MwLCeqjZ7ThiXTud5VECHrAknQ
cdVVYL0zUKfQd6JLydxpUMciSQw57hy3MeiG6JOqfajRzgDr884NPG1vKcUf
WWoF1s3eGHrBrBugslgtAq0gBRwfOFAXRJQUmpL4zz9QGC1QJtqR9EXehoIo
yq0SNTyrYdbiMbBD3iXtceyS3DjqackZTT27QKsCODEXfW9f83LZ22B14Avg
uVq9H/mSLQXdWH7/RtIYPGMwY3LKg4znfXMYMvmSma1SCFtwAWqQAKBbihRJ
BQLos2P6MliiicoyObfNklb/0TH2+ihRO0zUvd3T5uxdfzrKq3h50DCNseet
55WGC+jxj9BrmyvOsP4k6be8RS+g4MKuWbuNOlKy2THIPUi/tHgMtlaOBUXD
f71eO0N+EvjYxyGfabZRKn+gOLW4LQGzUibW3OApfCSs1K/FMvkhgMBjA3Ov
CJM8t0897VRvfvZsm+2r9C/m3YAMLJWb4Lp7qWILKYGzNs6BXYxq6Tnjywfy
bhLUFJFHsfueAf5UDpN/BOmGMxxdlbgzRYv8whC+7EGJn3EftVnahlsM2AEx
lZXM/RrnsjBN97bGaClSPhEwIvKmybH0fGrHslM1b45FDT61Xe+mocK9VYhC
1dcx1GoqTL93kwRrhXl03jKzSRrzcwNqlIQmOLHtwuMlZGjsMVf5bpjZJqE5
JHf02dRtKcegveFmHFnaTZyWug8CaeoEh/qXdua3q9nTw/jozL7zCKGOye/U
mFidi16XJ6cuFxT3MvNyXt/4WdTQ+EEaNimYDGSeVEkbRvz8jIRH5BLC3/0h
iJEfQYLnVmE4Rf+s/3rCM75UZuhGkPmxbX8gy/AC64KDeAylN1tKt+ApDh59
CJkcuyK0rxNwTfByLpZsXIrX8UNx7Qvi7zXzhGsLeyuHq1neG8ehfUJDcWDW
x9K3LEQL1sanzeqUnkLMabY790XX0UbwpXCHr7FWUZCMrR0chjv0gQzhNGUP
U2iF6u2LDCgiINs4tFM0BFYv3462idLDeqAnZrIenJE8X+G+MTnnJlc2qK1z
sArlzuEZFg4GJLhtzO26twnuVHt123PQkHvw83xF9LuXcy7peNl0A6jimAMd
ZD0WRu2BMDftA4EpfeB/8PH/z8FQc+Bls8z2t7iJAMio+Z4CxxzG1zBpaN7Y
KhRMAGWg9z3OnR5r777E0sK16WxL+W2jdESaN2wxQu2o4C8EoKSkweEy+/zS
h+cqKrnEBARgsKXz9/IMjyppY9S4rNIRB8X7sNJuGFBzkd9TXDOkPqf0+zH8
L2QXzgMjhpvH/s1BoCk38AzpnPh+ZZ8ybKCm1WgGnpM28iE+m8azC4fFfbf8
okS3LAY0OcP14LUWDK1qvy+R95WaYV/OzrLdU+c+DTz+bxR5RkAnnwWwmtRn
e+F5qerQSS9Vjt42WmuBfSyJZbdxlpYOEdQISJMA5zPsw439IMLtdZI8KO2t
CeWnMQ+WIKmhwRzW2JmlTzOaviEex7phxwsK0ERpVdve3QnatIRJR9sDPG0d
0e/qbbK4+LmurgcwxPxNmlpjOnNyiwxD/FSvqD2tbZF33pc+kIDboXHG99Xq
Azx57ww5RArPyMdz5DKmDshV6RGptKvsQGJK40LvTt4n9JdUtqZWc+WPFeyk
zcvVuDdbsBvTL37UycbUzit8SZb6hqBk/MUd5J0EW9LAqdKmYB2iy3rNB2Mi
gM22o/+DVkdC0FUEaIAJ6M5GsUHIw2rPMGgc6pog0TeeHW7oXK0UrlIWWYJp
rkmLGziTYeyfPXVOJKoPZLvD6u7Tn6apeWaVLLWfMAG9n3evaLaZR+WgqGlt
jdK7qPozZwJvkDaIUffObYFDj4cJjktp8NmfjKBV7zB0TLc/HZ01GgpR/0ce
r+KNY8Uyz6QHlJK7dGmgctsGaUSG8q4UScdVKic6359Aqwuk1qzbf77a/hk3
M+KcbOW2XXuftA6y+DFLB1WWilnms+zli1NyV63gssH2ArmRvr29r3VmSLWB
WmMfw9h0jMSFWjOU63okNPYPQ0dbGrJBgr+P5LOxvm6f3EW9bakpRSEOwEBM
xzDWs83z5Fw4ulEFgj1VaYmwCe96LFUnqb5dWLmje3aCrgviSlbM5gnFxFwN
5c5hMw4FkPvLKPNh08qejFM3pxhNSciUS50FTBdo8/gl7SiVEtRRErosiX/M
uBETQC5YqDQRS1M2CmthIcgFf3dp3mgs8iIgjaGP+W0NriAwQZ6q/WXVZlIe
YIxdc/jHbHRMxsb2BZbShl/tsePUD3Xr8NyUQYzzkjXu+A4Gg0VcqcEDt1a7
N+tUfROc5qCcH9w24w2egWYFo+uuhtC9QcbdxkKN+8gIOnguPs86j3Rl89s3
CfZuV1bkz2lSi/HepQP3CllemkGJ6B8HSXRFJPqKMbLaKWNOn7diiU43gUJr
4C1odUXOMzHHPG6wONkJUTrIJiT71QUnJFQHaAerBwRq57uyt/fPvtb/uSXu
Uc9G/x5Wc0wh2SD1SBVXePQqJGovXPdEG1cHNzbT3cmoYHieAjvFQoNk3AJB
klfIqnzT3C5Yd9G3raMWoBLAOnqnmyLljfkiy/NZeWvUtXvnIlgPQSeoWNJ4
x4N2IaADArEHZv6Bmxa1cw6pte9g20K5gMZVPNBNfw/HLgjllMyNYXF1DbtL
1yx3NewiDPXLkfRP3Jev7iRU6gWRP2EAxrdo9+MlD5TZ4w/a28u1BZnBAszF
EyXcm6XGGzJpiVoJL3RQLB8aZOdG8wxZ81Oc98rLjvamGAcvq4wokczyybcb
z6GcJrpH/STiyW4EYVoMhhu62lokNE0IXgEtXMVXFyQszB3X3TEsnGMAzAIK
9aRSiD6ExLSh5Z8u9PYzVFYJOKzadoFoq9naefpmp1aT9cprAZV/Lca6J4Am
jCu1zbg8Stv2D38iOh4Y44d45RCdCLJzXe22vzwj7ZVzPDBw/Npqs3v7i6/f
2UHzLl9dJ1HiNBOz8z0bO6JZQVD0EUt+73tsXQZpiOnDCfc4Oxkh/zDiQA6D
B3+O99nGvz+a7XcIm7x+DxVV3vGY5OogTIIb4iFbRt66PZlUu4SESqE4LOr9
53AHSyAaUCvLSdGnJB3vIoISu6/Cn9X+jQHnWegn/8KUV8wCTLOB8sw0AGfr
9nhtf1AkBkR3ak1E1EZuzxyBpAkBhWfJjKdyfLgUZ4ZrUbqN6HNojAbbM6y8
rbJB1MskA4413MZJphHZDYk22f02lacZwVXx4QYToFPJuqdJfnLyrP+IhTmq
BgH7Wd34jccHRLwDN/8db0vohXnDfW/naVSXpQY2FZ6CAydVzx2B8/eoRBA5
qrIi07spLy8wQ8VTu5TPHnuHFggOv06WhhYskJ+vOsfDlETRVhvi+FkP1hyH
u4G+9AA9dEKEjUT4+05069N3/rVXcMvTsrpW7aV6QhNgUhWcgZ4uA8Ikcyly
zJdJLL3eLX/sqmM8omLFfsPkPkJnePjeVy3ffdJdwsSWOULc+E9NCxkhfAXl
segWMzX52mvRKaK4XoUiF9L5/ZtMpDcGrMXmsoVJgaAQBHlwLCOrn6S76tgI
EmAaFVRLAlC9z3X8yYBQFCrE17v+qpYvEKqGYUH7kgB/SONqWO1Lwtu3U7+Y
S6Jg8dDwWF03oWPMdYoRdxGqAchkfH5z0S7zaLmPGLo7NAsStPMHgrDQ98LS
6dK57HdcPKqe44WuSZaFnre02qhXPInGAdvAI6rZdQ3IB9pEuDboDuD8Vy2D
5oDyLzYrCUdxYat5LQDTLOHtn8Vt8ww7OjZrcoHpffT/FhnYspCFB/IBoyzB
8wJO9FlIaoxlwwYMqMDoWnO2fLpOYV8LJEuyzRRSgIKDGaVzGzYawqI/3wIG
pSsIUmvxUGvYxaSm+jT/7VT0YQKpsF+79ZTXojx7667bXL4HCQLIvyhgGXCO
CcRhNp2l0b3tnpA5OUkvRoeWUY0AtcZO+zTGS+bVSqa48M42HdgS5zAKNrbx
2yl2Z4RjzaXFKRegHpBEhZdDyDq8eDa5uCrp5oGvhyosd7cpsAY1kOxuSMdO
m9j8zAEXQ3ThpSrtEaxwnPIEu+MluSErnbG94gduUx5tABUJidlXTbONTNUg
Ar4x4DcA+bGWhdmyoQotrQrFHqTzU8W96xBd3Tr7Jm8noQ0WYFXcn++fxlsY
0b0Ufft0WV59u719urtYeAQSpDBo3RezCPVYfnKjFv3jZpodPAxFYdV4rrof
GdbEcxUp/Pzvfiz1RfeAgdUTxxY/h/MjvX73aI1yhuYcUM3HIbcz1ZA8Y0E/
tM7NQHwpsRyqstPFX++uHALpeP61g0JaQKU+BM2ICmXTezowxOdwzPg9xSSV
y+DZuJhWoClaTWKNcCJOinLZ3sZNiOgR1WH5L5PAKsAvQggJt7dZB65oxw4l
f3FhS6F4Sq6sEnP5XRv8z+XoT+kkSoi6tNWc98qlWu6CvhLF1teEWphcafFg
71wp5vip8a+KY1gWAy5FZ01tFFkjJXhw5Kjrbjrs7JH3hURa0BXhDNYCmY1b
+8NglXJFHigKI6XBmVpli0Kp4k1BCgA91UkwuizoM8dChJhtgkqgTYtaaPCU
Qg+MBEEsOX4xmwUHDjSndNFjiyclE65H9guUwFqL/Jkc1B9Z7biSHPHTyLgj
//qCSf9J0HF9AKiY1wQxDOhUE+c14cGK8+r+aHLbheNk6UQAu0FhrYMui7iH
AlvIohUYuH4e87xBuigPwzYGNgAIYvsuD5iWV5uBgMmW9atlf2XTIs+nYtg2
nyER+5bjdXaoG+t9deWCxq+DqD7lK0scNvD1ZSov/rp2VjADD6zWRiSLGIIi
6RtvMrzq2GAosYb1ZC9m2tkMEwTiJvT/3WTOy6t06KOSiq1oqnBiWQa/kWxV
8ZjhNe/L354Ax8H2uuzZB8p+AxpWXRX90XU3whmYo3DzrrlJUdJew04E4AwC
hxgFt7E7tNDAZTKWuXoZRgo9UUIl4XGUP5FSnOO9nV54wVP+LcsmaGgw7tKK
ulZjP1jUlPzTcSJK8Cvs6uhlY6Q64HFp+8RfHeK2tn1TLUpj9q85YeN9/mvL
f3e77SL0um3v9XY8UA/LQMaR3iZGm8wehBSM+T3iL9aEFecbGdD3+7+6tH1m
StyGSYIYWdwlNTarUr/x7yxMeN+H6kQLRXvvD1WFwcgxKhBntXOQvnzg/ZdE
yJWe7+isPk8ignDO1oYI5xCNDVZvwJVsdx8BukCVC6bRHySSkaqpngt3xqPV
rN2M0D2SJp3B+UMfUUJmd7ygQhOnPGS3g5BqvyelSNbDyM5Jj3I08kZXPqM9
CnxHdjHPBAjDdUj7MgWd1P9hb+psst8Jt+q5NlQ3hila82a3TiFkqae8pgLx
N/4lfJ5SLWJn/Lf6pHQ6MguJFwclkXgmdtB30QPoSO0PXAvwi4rUEt/euAy9
oBceyTpdJBGgMIcK+3neSiDbUQW/ekdOe/mTgJhU0GWhupXsv4gRsX2tWgCA
zIR71CpC0YQwdyqp+dzOZuPKWMtVkKdLMWeNlmgx9JXpePBIV6jDTIIpJJOz
RXLAXzt0mK+cw7S9i4bBM/RhmN3+ORk6wpmD6rE6VFTweo+QvhXIhNw4HSCc
ShhjlUVerBJonthk3e5j10hDQ8+NiVTF1PAZqGzgpEIVLKuj+499QbpVOYsg
8K6kyNoQh2xH6WcbQaHaSDaxRXCk2YusovnLc/fPp6bxMzlf5HjJK1AJUKel
wCTPjiCSK5LRA+N5itBzvNrFbLqQ+X4aLo8GzDlBVS+Msm8k7IxFPE5sH5fF
JaL7/bfL3CyagkoZ2703ZJJKTbC9LQk+Xs9ckmf6lqlseJq3lUGbuLTVozIY
4C5pLr+ct9W2+WFs9kY+oHh+HWGUnSKUpmkBDVwWUiPhSNAIjqujDOSPUomS
7imDj+lqS2LazWAc1W/9DrC88HBIY89jePT7o+ZZjQ03qJkb2aCsjbRvcZq7
aqRR90IEAkqNUnnorAEv/S3TeQGVmdPoTQBHu//uMWzZdtEWhvfSHXA5hEv8
IW4oUDeZKf5IZb6b/EevLqL+YORCpS253srEjdKmBi+hML2EQMfS/jcN+1XS
AZ1WUAbVSgQpK6rnXSCcejjaSSCDntL641ipZFTKgo5/ym/kkTBeVGevtDh+
c/OXfQdZlTqUn+MKn3NkVKMw5BcfPFy3qMvc+LWgUlTLMeXasSz9D8EsF+m7
3oXmRygUnq2C4XszP2ff3frFCCbdSCoJeyk063LBQ+K60CXu+7OuLO7mK6lI
U8Av7WjKhIEAacmyV4Qjn5vxEEkIwqQ69zChYkq/cFAWz5fZDUa0+Q+CvODk
rYSFfZc18prbhKsz5enPmMf+b3tTw5M0SbVAK9if90hWimUH6RSwcQu2yQs+
kgxjpW3O8ntkM0snX6Cl/Thwj1p0RU1Xth8nmz3XsSvirWVEmJ/+RUyfNRLr
igmdZzLQ6C7IWYuiRYCYPrLrrL/XXltsyxuBrA8BlqNsHiQkbG5nDsq54qqn
/47xLvdSWXZkgQoEr0Yl7b1oBnPCK4uosf2e2bg5jIS0urqHNfzlgQU57my1
pgEOBwMA29TwEk00obeaGc0dkMj6Pdqn/LJdqjBxJzC6jljCQN/dW2P40ABn
6sSivM5TKEs3NoByp2R5uECZq3/JN6ot1YhRNRnO7yNQ3yZps7WaEp+5AwXp
Clm+ugQVGSv4S+P/imAMScpGH6rUMTlHDgKl6JhBAQMD8yvrE57rsqfwiZ6x
WqR28tw+JIjIxrdz6nQDSqMNcaEfj0BRBITb/757bJJZPHZuMgmdFaAryVZ+
RiyQ+7t85TWwDoDCj7BLS8aCJLBP0WzopbAvjx0YHbw1WCj1ZS5SuUqWVdpn
sQ2GfX+98hv7ytjd0TAotPG8xsp74gaKYNDQJexH6Nc/iXMPpSasc7gCGul7
JnTE2bHzvEswA8pqFiXKrK/I8emLxeo9erTFjomxfwoz3BE7OItMvwcwSThe
K61Njs6GSyiJmjc7xpzFJexQw79fnanD9wgN4V++C76y4FZkH+cXub8mkq/N
/dk3G6x0bjosJNVFiQguYwiPW5STyp7pck9NRUKMlYCNLVuJCFpnQ+ew3YF9
jF4P/5UDllSc5PoBBxmwRHh6U1cdExnEOqP9KlAuu1ph0EmbYMjTd27RCqAe
tuFTOAvd5mrBm4Q7MJEzkBQoexsOZyJ2gztQOT9XXvS4o0ZFFAeWbBJQbmgg
PuumHji3Cam6rNfvGDSa7E8Vsk0lvxDajw1UD/iFeD2DwMaCmJYBrwUKrJ9+
0SHT/nedmoVq9JRnPafAScVRrQ8RTr4KLcMoJMnqwc0tuFZg3toNoqjmkkZq
UMx52sKir/jMT9G4MyNrpxZqRRGm0tBzdp8qTZIcYAGluazifKr4N8b1Y0GN
GLKqVgK9NLayku5oVg7NgiyhjhUfLlCT20GbO90x86BJjOBIMMWq1a8hGiD7
mfmkKIkM5slKCTjLnaneiyc/IGR+sd8hQVDtLXMYmakFvADuWAadQqO/Vvbx
9vDhxvXeSO/rY265X4aUGTgiYzFJYVcShAX2fhKaqtxRhXOWDyzX6ikfjnRn
E+Nniwq6GvPmiVPrL9XrB8ZgdUnxjd0x+LRmEl95mjz0dHDm9mq08Em1NtgU
hXFSV0cKsdy8rscem6hXsSazeKRzYAGCmcwuKvohbbH9m9kE0/8m9hLgL5D8
lOC6QH2jSsO9bqroYT4hAtkioHfIkQybmTXJQVwop7emad8v78jgFT8DCIgY
TgYnmtO8ilndL/3B8ApPu79b0be1cTcVjAR5tVA6d2P24kf3FBC42qPE6Iov
vJDSkKzVYH6b1cghR1ZKNDqeA4nohPGHJn5nY3LWzxNvHS0zBkBXSt402R7C
deibVfQvGFJOB6iugmByeJv9TDC9aiM8z7NaZaJUdsnuVpx2a7ACEhnvAVv3
0BtOoZQ/RJucwlXtaIOA86EZjhCfbf0cNRbFYNyGX3gfTfHvbW0NQxhBBQD4
jrS5ke9O9gfR98UTGBH+SF+DTVuz/g2bITs2ZFuPexgp+YmIZQzAcsDJdfBL
GG5N69gbMUCxnv/Y2T/jur4crlTCIR8rr+dp73jXPNepWpXxytLhfi+dGLpj
7RulCfFK0BjyZvEikW1aSOkI8giZosgZdDrahvjHeG6q/QLVsB1V1IbqlKyW
TrqZAIHiMzdXirB141n2cJYc0f01ZLCCgpgHnAu5uVn2+WNYyQxFho7FPSvz
EzPKu0uHPCioL/OAOmZPvrHanm3JWcsYt1J6sCaU1THI3JWD9MFqd9UQpPQF
485PilVV5/7azPgaYrdko+e+YaoEI1SYzmkD+yRI76dDya+rOo+LxjjdtyID
F9MfW7Ziyu/gsmFrXc4F+iKepRlYvfhaJr7q1nfW8lJSfFZG/Aj4qVHpswJj
2LYR2aujzbw4EQOg1NUjAfcZ0ZmePZxzJDQ8DQpXJC7yI7qjmgOIt5J9atLL
KSBS6c7vOnHaQvpLmg5e8SGV+WKTR32TZUU0wDk25+EtSMQxuymPqcGlmgEm
DSXn1T0Gm+miVyF5/QYKE1koFFD2T1jtiNvzrC4fpgnkiJCV8jz3mppxrmUM
gXKm79IRU3yvW2kohA4leKCVe93XJaeeUGtmG3u3CUEdMkOVhH3z+j6FSlvj
XWD/F9EL5sr8FvCx0yUQpX0X4tycaEu23DvWjuaPSL11VLVKuT3VbwdIdS5r
3Y/9bXi85wZvH56yNbTHvuOrahcmGkg2XekLRxET/c7pf5ta5ZEW1A4s3uBE
nbltXRZcN+CNSQohCD0RNhLbCQ0t6DpNrG1NxZ6eMebJL+5FhTbtZDfHfFUN
ROYql8dLIbfUXTK2powM3EN375Geq7ZK+hqV0lVfmtP0R6qx2Bkluqgslvxq
+EA5dkGF96pLzEV/makqgFFD/1iOt4E7Z0Deh24JxuKYXGHYpk3V/a0O3vXT
UP6e7cArKZKqqMOs95L2v6whAkr9ZIeR3w0RXv8nnvNI6T5yRp7gJt821BHM
UFObSIx4J0A2QoyQNDJZPG4W4fJCSLiwrV/2USzO8hKNHjUcdWpzReSNtJQW
RNaFQ2xNZsRQe8fK/R3p/nn+fD/t1D0Yy/nTPmE4+8nshWNrHjcJpwzJzs0y
7+Ga5c1pgDsIXui05q7HUcRrUawvixXYdx6xu2kVLEL/Y4XWEmI0V3UKAb02
6jfXPTBE9L9tJCrfamJBzwbLoT9iZO2Cy40aljcjqydtuhI288vfUMbSjOtG
kezXv+Mrg7LZIfKRGVTJFTH/V2JNu/BTN7H1Hc/8+MItNSZG30FKz8Bn2B1/
It7jRPqkFZ9sQ4CmBOvWC65u1HmhEPuXWWLXDqfUbMf4WBBLvkhHcHubiVl5
yIhjQlxTIJaT+usZns9G4mPqgAqc4nwypyR1Lg1vpD2AADPpokjrSt69a4T3
YSs1RvcRbcmo0cqIBGkHVIib5o+brQdiKtURj2PVcamcCHaboevHO3NTSshB
POCqNY+l5xURgEKmOGD370ArcyCXSqae2d5O26W/yxHgjeZsU394GO1/j0fn
ec50gQupxU3cr3Am5f20BeZszyN+4aDDwGvpJKfkE+dAzO6uO4ynQG5DWHcQ
Oom/zV7OeB524G0xjoS+dnpRF6eBVrl9wHl+DH16/n3JiFc0OUxaqtiaLA51
ck2JlAGP9QS6UJDYnVyBde/nqvlJo6Z3e3viTPXXZODYaXUega95zFRCX2+3
aFQT3oNFvQJm9V33YYezhZsFe1C/PKHpBcqeSfWbisn8fcmq1n16wsdkvhnw
qzYFfW1p8TR7GT9E3iEVShuIkfwt0CKKKnjhl6NDja1i2qvFlmNaMGVLzAx3
qAiZ+/k6jvYGz+VJS2NEqNs72yGnBO3RPm33TyvICLEAWcD8nwqNwdFC8hV5
MbV0evSDjjP3+Xdu7tpvmdybF6rcWSX+ttz4OrDFJWN/ergrsyjNL2NL9LE+
7wya38hTLOxuGGbIPN+kzVlhHJ+1+yA4AhaWSNw1+unVfHr8nXTJD3JFqBUh
bcQwXsnfFf1UwU6G8XTdmlYDVxRVMS80yCnJY5/Hss2dgDUVXcuJ7T9fCbL5
P/yhS4AeTKIM77I9Kfn7t1hLyaPQke1+ZkZc6nOaanNM5cmE3M4+Nh/KzR7l
qlKVgjifERkrn3ndRvVCPTiVqGaOHnBk72B3m8WVI/J+kLUUfnGEMmLxsCuo
nLJEmaG2QpgRJdtlnQo3bfN3OOsQW70f0rYXBcHyjcaDoEP2KilclVR/zJSp
9nKvufqJiC70cjmRget/Nb5t7bXKne/OBRDgSK1btLdmeFuqp+PydLBcqFXH
ZrYykNmipAle2hncQ7y0UYAl9GoSE2/CfIN47HQEcBsQovN2JmugvsXFZATK
/wT3guUSEv/QbL45Vms+p/pthUXGjnXyVcRqjBEwqswHTT4q8k5bDi3IRw0v
CA6MlbJLZGJ+oEKbVERJxOnpJ0clRxUckpRGajpvdniGKvAFW2cUUtlMP+ig
D5GpcYLtR7/daMEISDmChsgc2qMBxdr3OP0Cz7tHfgtRiosCPqhtOqgiqOeX
K5zDo/kVFxPnTtNeA+SiOF/2qLJj2bGbeLvQ2RueA6jf0PXdU+T7WCKwWueQ
UeXWd9BulIuSUzpf/BtezkL91IuZz7RLL5eoTztl8JjBDTHij0lgnowQwr+E
RlU97xhLhgdv7x/mI76C1cwfwZc8hcQsSVQjZ8L9Mb+1A1s5Oo5l79PIfZLU
fNlx/M2wvMRGBXtB2j3wmXj55xe8UpysvUO9/FamFfRgFtP/Wv1LxzZIBt5c
7q2eYvfoP5UUoSnYEipLGOtC2s8Ml/k9Bw7FNv94x6PMPxSEtKigPvMyok+v
a7ywYx7ateBZC+ycmOXR/kQx6gUk7BWefYBgXvbKHpTvLPBxhN9JH/zVC0wo
ZjpJFYy4W8F/geD9rHCiwbROxGuxMWJx3d8q0E6m0lTd/Ex+1r6xF8ILdcc7
d6N8dDrT6FpJ5N/W5vR4orxGygfTSy9xZUF8kTaewi/uJYxh/U/b42uynzBB
itcqi1XerYnWD/4kJ0jsBMsyUu3gyaHG1eVANtDGGBOoeHJK5vy7ydTCBd9E
W1HU74PeDqnZDsy/QS3z+/EtkK4y+4WxYv6WK+2fxUWdSrW5aTGg+xRXNHTR
ehjXwtNRgFCu5mKdzZeybbF0u25sW5xNDsEH//Xr7QFVwnxgYnXJ8mH3oaNM
sfaS0MnNrGjlCVEom5E72UWnwj4P9FKPjW4OFK7u8pGREKfIJHdQgDBNmn9r
5jdbxztSZv/c+vW2+Q+7SE5xPTp9VD+1g6xeCiZGwRd95nxk83fDR9KrxnHE
nsuWkFwESzpdMsPva90lZm6PS7y3vYETWcAFlk6BeOkx5SuWLDBDdkVxp9nZ
jIkzZ9Uu5TXC6G1EPzb2OEuBZ8Lw3U79njjOGtPMQuo+Jm1q/M0vFtEcCbDr
XLvgcgGhDQS6pIotwzKFS56poZI8RwT+QtGZdTr+/t0eGQnBYa9hyX3hXr5V
CQeuYr6PyHF+KuxHQo3nWLGBXLFTolggx3Q6Yfp3Bs6KkhaAgB/Pp/OOExQg
K5iJe3dYuiYmEAVYzDX4wN4Xw64fAKr7YItqkYC8a9EeUVeOu+2aKUqa2zrT
emhgV390HMq8rJMvS+7C9Swedm/vUwML5Ir4pOvHlbLngAoMp+TWx2SMMZu+
I9i+64NlL0E7cI24nzXTJp6MDsMJ2fyLJH2wK5rP0K/dHDTbMIlttL+tlrqc
eviw79ilTXGQtnlee8TkDTN5+DFm0E9iRmx25DE6gHpyePNkWyehiwtb8vOD
gKdJ474Sd7OLxxBLs6IkEu2X2qpSsfOZPRbb+bffcanyZB3DZyKmfJqNk+C8
k770ZDEmSP4Gww+kKb6CXX3R6oeRQNiZd0J4MrALpN1kjnkFsnRth4+stzUd
MgqoytVUAmfeifizOVf+VV/OmE5dDegzcE0BFqqxAxk4QvsLqi2i1+yDBhnC
ncFRha5AguXOW7/EvoKeenjz4ttI95gXF+UTwK8s22vJ52gAXTlbls/1ye1n
da9IDcbShSgdH504S/fU2gj0+rxinVR2h0dnWV/ieEscbhpI3OCFgH9e42Y3
P0LIgsK0wyklbrWaX0pFd/Q8Y6VYjRrDlOdPOwth8nGGPImEqVIcPfdFlesw
I5CcA5zrBn59D7C4FVdW+0FFky3NfS8glTx6zS9xj2Bm1go/wW2dNZgPuxWJ
6FgHA3rmxo4/g4zuAF1faa9h/b2ZoPoE+5SxKT8oY7PQhw+ZBkhd3lJqo98k
zhhurTfyPqXNsPTL9S6e7yslYyAhPtqdrqli9aV//9ZsG7vSsIS1TN6ymOVr
l5x7JaYXa1mlbb+Z4V61rx8yz2uGbd8KNgVT39wik/T5m6nheiaQvE4RCNZl
TZLh+sok2uifzPkSaWYli6A9FL8i8oQUkY9X/yArZGM8owTGl+tK7b1OlEJ7
O5HERS0chSl4/kBIiNQpqLefqvnbttdMslpPYKrhniBlldnKC9nUVGof4jQK
qywfHsibCyYGp17cSWtc73P9ZpNzyE0DNldc9jFB5gWcwjmxk1CiWhjCI40W
LOxGAul3OO+a21EeEtgtyGYT7vHHKVGxyN2bJELkfYc5aAQ7WeP9xl7jqOXd
wyUTqZniuBXv93qX6vkutONm9peGkjd5ZjMLUl7bqXi8n8K/T02QjLlanWb5
fk3Q+UgIYJMYNlCu2X/TATn5gQ4PjcHPn+b3kuzvaHTohtA2rIKFLBIS2Ftj
SaVZetWYQiLDs1iD9o8di/sz6cP5WUVsiArLJkA5HdSOwRdDKEryuKr5LLiR
jGTOrJ68Mcp2t+dbcg643YoN8GaHhAL9fOB+m/69bmkNDRe9LqkeRlqJz9KN
2+lvXIAe22yGyiO8mC+hs2dC+TrP1aFBAltPCip9uwa57IFVvs33XH6lZjCQ
s9kPFLOESCYeejNATT0j1t3QaAwlJhQewXaF702U7s4yOEfVf4kQmXrXfeG6
Ja5EI46TxeJNq0VY55u7+deIP5F0fQjF6RoTtEb4kCZ+DqW1n/0A+nDRAEXc
kF1GrbGI6xZekntNPsLBMMdIebYGeplKbb6y+puD6pE9MXEcPzmi4Giku5VA
NQN8gwj8MB86IBNVEGGTfRUqhX+RjYlgILaP0hGaAAKjIXVTofny1rGyFWj3
+BO769wB7LInGbG9mJsR1isEoRFehcXj1OXPIBhwBr9mXL68n/ycNzdp2K1k
thPyxKNFIQM1ZHZsFKTLnmOR0OAhzcQC06orj3axi+uZL8Fu3C5CX22abX4y
bleLBvdr7l7rz+0CWXIXH6PGUAy5+ZXkGwDNXgThJ3xZ9SOKTwd6MPCqf3Ep
PUzmDkyVskeV/pM4HjeeFGd7bkqkmH+zjDg7YAM6opbnXqq9dzKsW3hqFNPB
XhrmWeybRu5stN1PtpkmlAgCzrGXzg3ll75CLWns1zVsnnI7mgXAHeFWutR4
9Hg8mZtR1gFap/XNguuTWzD8cqhptnJUIymEqzy0NgpFCkD52KxZOA88AdM7
U664k9WktAloBNwQb6KEfbrCRffU7+xpIB9ncwa4o6NABHCf8ALDFalkHITA
f8O/kUItFsKdtqIHu2vANki33u2xtzDrjMVRg5i1NGooPlNWlN6aPCOaUCYU
WcBtm6OyKfq6F4KDvcvAwV3WBgd208uHwWnKY0kAOTG9kl3tl1pRqF4wnMN/
1/FGPD24G+j/CDdCE2PKqn9xWcjSo50VVrObjT2VaZnnCfA90gof7M6Eit67
FWvCDL0SmyROwLNT3Kp4REXceJVxa8wyScDYIWFU7j92epNQjyxbPx1gSOvp
NUzOMMByOgkPDBHYznxG+wFAH5YxfG0imJnSJphs/mZeHdfNtGNsSPGAoRIA
CX9Txi6eYTom6RfKmk/fWj64Bxo/NwqLW3sFNYMl5ZrYivDuEpON2FRoRv+Z
W19xPcvqvDyL8CEdvp3fTaTk6urvkw6uHmfFulANKVdGV5Vna1EV32gT+N4l
jHa6w2qKs0+Ap44ra3KuPfcufubtwLMjaZavEGeNA4Y1CNIXNfTJdk2CFtZz
yTeeqjYCOs7w9vRZmzXM+nAvDgKqBanvsgvTZSpFIi2TQYxOamTLpxQLcvDC
u0e5biBor1fQILRz/HkXEcQahNmJqnU2Fxe8W6kz1PdlJJnp9lqSe4oIssnR
XoJlQMxg5FsoWZJGiVD7qoyGGvoxPaRmYGoexQuc8skHWTErE0bOnlPA0T3j
bF/bxB55ggChkyonXuQOTGHt3nzD12w9Y6ORCEWoL/L0mJpMvqzjQux0RUwr
9l3BvpCLA3rch/ZX5bgjjsMUVUCHGl8PLGhidHYXvvedHeNNHY3p9qMo/BsW
hUEoSfvDZpAn4f6r7Z3bfyNwNpbNBMoxJWDnqkwnCp7N6nBqP5criNNs9hAb
gubskeATfUZPmOUxENxa/V8gZ6y+29PAHDvH8/ewEuIY5vnb06LDfB1124IC
AomxYpMFWLh1CUauISfZGK++MghpLnJnnC5wLJWS2e36iRrx0MpIJwC92cpA
qzt4Tp/UHtml+hxEFFfGtUIVYM3xj6Qw2BOSUPl3W0hc2TgqT6Lw3IZ26kYp
GD8YpiACb1ubtT3bAQjdxVXfL8GKgVf7jX6SPqPMehd29wK5Bn3mQigP7x/N
vMRvU/l58MGMhQyXXLoOV7dL0ZiStodEpcx7+Fk8h1u2iLqfQWPs82aASzz0
nvj0v2vkdsGEiXlxkgqaa7CU4TUqDMsKpMKTbfBI/GvyANS7GOhq7EWIAsUV
C4P2ugwXyDqtIvbxmLWAdgrbW6EURDuMpuSXWLMKBGoBHfz5MtE25Tl+u68M
htVlyFNPTrsBjut0adKFIBow03jRKnCUwI3713Pm3NBkc/OOL60ugOBui0pP
c1c3sZFMQiY/dO+IrFtIQZKxnrFVUbf1tkyQ0bmM79zw/AZfJeNmufxDWnZq
fJ9b9NZFyGLAnAWjn2WErCrmqhww0mkhH6aH+qerFb1Teosefzg5gpfobMJD
00VWIcQFspbk1Mh8K5ws+KaYhKg0VhqwOcmhj1VE5GBb0yfnHAWpHvmy5rHe
+15ayfyUaDKCA+xDlqJfm2ZORhfdyz86HToZuYOKwlUXUM92WUybS4KlCSC1
kU1zQR8HB7MR6cLJtBtinAC692jzUWrB2svfPrWlbeytyRTXVrMmDplPK0Oa
WBMEKZq9T/3kJf3mKrFunkjpw80dxhPSdv6DCnQWPQX6BJ1cNCL6XieXvW5e
vv/oS5/txYlpXTUkpYK/UT+LO3KtVXPdE18oF0KQSgkvSSmBoUro2p+uf0m/
3IPvE0wta8+f2xITei3E89jKmFTxIbPYbs6XEWI+DmHErkMzLbj38cmaHb1r
ER1utKc4mIhOlsNjhP6GtqXqoA8LqHn99PKcaMNh0rhPdxGoSGaypasQIKt9
1AWKuN/Lxocm/FPp6JJegs3P4RrMio4G2mpdqnCz/J0pBl1+KKtXUpItWYSc
Zmiu6Cc5Rq4H2AUTPFCloiwaTUIZNuJMhQdoAStKBRPMwFcvfVnIWbMk/9zw
dP8dvjFb1dRWDuRSZNVOnRKJoKcalDKjcA/SmjTMRvFwgSEPcE+KrYnYhM28
mqbA4dIcYPscOepSAAvzH3VawEMlGGQXRrfN94g4MPbL/QV+XfyU4g1HjwTn
XH7G1kq9q/RL+d6M6286OecuZvuCfBVDjm/N+xccnV8rCfccSWWTjuWd+rpB
c6iCzASjQ9cknPCSjG16SfcqPlxbMFkNSLt/taXZYWp3UyewPwf3uzbTb1Jq
ypAlD/KMnP8z9Rl+r9sh7QoOKqMDEtCcLiDCq586EpKGt7FocoNpaWSqRvlR
CiQOnHxrGzD2uUCpxPKC3GxiTglxLmjkunspv6EHXvbW2wfEFfVNSHQYA61E
zC2bKYVpinhakICi5Kpvf0gJJY57G+hyy7ZNzlwtvZ4pxO9wrl1B6p46K+NA
Wsj7j7ZUg5ziGgZZHBUPKkt8rCrRQCGrXdue/PgT/Bxl3WlVEPRLFF1OGjAm
ctizsa2wHUtcqVFrSfVlY/EHDq6CfGjsk0UfVVi7DOYwAKH5ZRughBbddqDc
ta47s06Lhh+vhMcw9RnNhfHqsBCGXf6iD9tIMSZb/yCle4z3NAnO4QYsuJgN
koeI7Lsroa4kaJvd0QzrJzZ0ABW9xXs1YE8DmWGolA9dGnnIvWsz1SmQnLR7
XLAQAQbOCIoWcW2s5gr3LohPVeQ/V/T2vMMpB2FE8ez6i/J/bOdE5e3uqB7+
z9WLbXjX3D2ISVTYtvAPSmkRaWl+WX1m76bagZuKsLxgrkWTlLQMuHyul94I
Jqo76yZY7I52wA/aSfGl3P7mAngU15iWCEiQPa+ADnl5SyXoLzhGK3DFUxTu
XmNeOllxGKyet1FgR+QF7pbwzpGBch5BY65WOwuODJI7+DDh7Jvy+Pr/S2qf
1qmrtb42DMTR5unXttM4H73s4WGxLy29lSQiJdsrlT86QQf8SdL8nxK53SAJ
1pKAh0wbQbG0maqHtjx77irer/exADXqEMn/bfvSncm4Gp3PmGZ1IvA+++yL
JVDiPr0GDPcjLPqZRV41dgDhbu2lLTzCF+Bx7LPzcfo6XLIXsUb19QElf34S
70dwOdb/QA84LpUGE+WMGsVldMSa5jWo1E1Fqlx1JE8ujL1ciScDTnHZ6MG8
DPGaZT4We38wQyiKraHL0tKb4UiAou3+XeWD4Ry0o37MPJfBd/ZaJEgECAVS
P5kijXoVVZhhSqANpgT5gKrDFud6at5q5wAUpeoS5KDRXw7sLGJadjoIpN8f
+jUHGAZFXTIwa3Fg8YoV7Q2UUVpz0n1x/yLiIueQ8Vh4QhZBaveMMZliPQKh
2Zz6HRZJ0cGfOVHlMAN1Dot5SwHs5LJl8tebfexxHkPFbjmGQYdDYXNZwZkf
KP8gm8Vv8/b/+N2YveNdPefNsfnGkU7SQn3mMLHtaFcwnz9YX4f8afUMzUBL
o0L1cIWXHDBIkbz2pJ6KXdg9DqsZL9mwVtDXyjOCKqKe4jZ0bgjUnBVA3nBv
omjD5EZJOVHpB0EZ5KYyANI9dr6pML0R7aVghuccBHf/JPaSTgbPDQTeL+Dk
YfoqMHlK3fP6Gxh+OKAD3HewN2WUkp9rhgTkzkyILW0KoNnmSGviIZT9QJXN
WyCMTmFywy0j6W0ZWWH8GruiYdkQXF0YcW7wVM9/PcsfTvRder1/t63K3bU4
kKT7H7e4fnbMMK2ZRlAU3wXFASueCbzxoN6sGoU2vDsq3lJCzjCWM/9CuXLZ
zGzUieRQc/7dkblQ1+DBmEgI9MEWoKUYFNqU+/pFaCQAGFqfu0vLw78Q+uN9
wg4wEjwkYUu37wXELVHIUbLHqjZkHxAB2YrthllECAcDvSQSXiVLffZOQ9LK
AGqg5ATPPS/OXxomEDcoDk38tbC3OeSvCK8Henm/0nGPp5a3xVQIVGTa/rtf
B2xt+qH2co8JjQGQf7X0KUw+MpjyG2pj3dkhX0ld0wxOrom6l+GrP7T2RZCH
CqkNnSM4qYJgINMSOJRu3C23kihQSR+YFivWMIHh81rKN0AVrwnwG64uJbp2
mRpFZt12AYGOQhLEKHs4eSNo3t77UfnMq7tnFM12VBc7UQ7q3uYHJbWTR/iQ
1grgZIW6c49KdN01V3YPt5jyE+Pt5Xzvd3+5kjpIU2Rr8zQcA0fWxEOYO3cX
bvy4P2AwF8FLxN/BEKnuXCbZN1T6DCZ8dUD79KETJl42X9b4CI/O1xcklX/4
Ps1TdYNVA54jp+26rk7uinB2IoJHYjXVMqTr+d5k/2TrUGf9+soz5IiXqeVE
xIzFL342n7GMy96/U9TMy+q46KQPXCmfVsGNexRkvpSRl5S0gdVPScC0l6jA
+YtFsMVPg2JPk0ZScI/yF/NoaTqfQ73l04euCireDC3p67ft4rfQSj5gU0BX
oVmmxEb4TUnfKpBj9DfXldLkEibKm3VEvHnpkNSHGj0PP/yNVlU/wVS+WF40
ZqxwL7hvR+WeZ62sxjYFelVDz1mGQodAU7wrkDXzrJUUmdFaRojjDPDUCWxT
ws+D1ZGgMbT2EYXGhpSzJzP4zkcZ+KjCa67KCwJ1ccHR4gERQwwOoERR+Mpi
IfvUEPt6ibtHtHW2og2vfEQxOhPiJ0uk/Gn0xy/eTng6UJJEm4b4BHcW8mh3
JFLBhSXABKRuq2JRKghQHoyH0VHMX3GBMM18vXfGWLv5SwzQAYTKox/nT1wN
WbHXsG+9ObkaexaQODNmJd7FMUzc2LGAnRDxr0tMv2L2yOcyZpUXGBGhqs6d
U2YvOzwF7fs9FNcUJD5A/XVXB7bzjAqSeN6nkdgIzPhDL0NJll/3GuEhW8bC
+BxWUABXlXeltZGU/cbfTFCxtkKaoDSeoUwH9SbxxjiJxbXqhF/3ehGV6RHz
yVeHgQK1YOtjqJa1Ea0FdQkcmbNqy9U7ntgZ8PUuqXXnkoSGYjco6sb6FtYs
KC33pJeT+DM0mtDVRFKM0eTxXOx08CDCD8bHHPgo4QlJMJ+0lWmwapnFgFM/
1nibEs1YxvsycGQ/cJm7I8R7GDnDLOzMnV1trDTXwxv6DiAHbcviH8G+Gxd4
GksuuOqPnmFn9o7niwT7DOqXBmI6x9xraGDKA6ge7hF1NgqlCWg28oLfZV3m
j3Crzc4z9oYQnbMf3oR2Y+JCpxKt8xaj8jE29zbLhnEqMs1VvHr/5pJlc1QQ
enAU6Rr9JO1L3ZmeUmj099ofPmGf5gyF/CQmHtt/Ld2X3Mq6eK/271D+etNg
N/KmVcx7pLB2Aox8EwDWeXJCSfXist6spLuJtDBi7nsKAGNZ4XBKnDYpuxeS
ByXUGCRVmN6JLNWt5O8KosPXUh0maapQOyffanPlMmR2RTYOCPVp6FwGW23Z
M/4cpZ9zsFS5sB2FazSFyt0+mecbm9Z+o42PmQQ5tGnHpdmbDVzx9ykzM9WE
fDpqov8bYMrSI5CcRXDrunpQIxeiYACmX1IGNAkRvockSGrxxQ7yZrmw94aI
Hya3A2VHcWnfmxmwvNNJSJ4Kxr/rOMRYw/6pK31Yw/HKqORkFINPr3ak/D/4
6obUAZJy5gkCbs85nTNuJr5XetvRAHVU/6hCyCjO7mkOhQQyQC5AzH29bG2q
BA9XqpA5gv6yG1i/hUALefrQquh02jovM467tvHbT/gkVKEjXVWy2JEShpb6
xwwLA8plEoMlrgQkZpDeaoxWqgyXH6sUZ+bPlUQI8k7iEcWaKgFZV6eK1w/m
f2JbXye+nN53nwF6XkDa1VxpG2tOoECiULhWIX9EA+3bBh/0owgmGTjJRwmc
P98ab24ixdh3RTMSTm3c2sXQaD5QQmkmVOIsIbIB7ojkzLhhnEav86hJk7l6
MY0AlCJ33ONtsLWGSd4r9iYvjU0tn+eEQzofUvWCGH+ltuT3ExzXTFpIB4Yy
EKrhRXDTk6o3USK+7SYD2/8mdw93cXsTVmcoGQVSDWhoOjjHrtKCr+X2Y9nP
eXCe0cgNiAd1BEEO/63GoMJbu9Rk7Ofup/4ugJXRmwxHChlfTs1aTR//PiAh
+/HGumu0ntYdI8hl/VU9gLxum1fRl2jw99VCoD0CmbnB/ob17wId3fl0tc9E
Zz15NURu1eGt9H4q69usK3nfi+zvm8fQ0UY949iyngEECvWMYjVL+kynD1E0
D3aw1jgI8xIRQUq0wyEH22VGYPdle8GnDnlOMeuG2BkUnXVsCbP8XmKJz7Ez
gGTlXNzzGiRjQR05KmX9r4OZ0yOhdlAH1sYsmdA/0EyDkwk+n3OQnhe4Jajq
eUD3+PvVKBv1Db2VUAKs9YfcHPVPs2nFUm1c6DpsekzZHAQhtrggtMsEtQom
VEafoNv45qGST96ADMKvdQu28MaAqUiQbC2X/qqubidmGkJZY8puO8+iWko/
dhwHRQYzwrmgh3AOYC6mB3xLsDHW9gJCuqJz4EuzYSTrm4g77IQn+BVMUbB9
3vD+UDIkXf3FmG5L0NT5UfUQqPCassTIrzjip68CHwVmrAqXHs7pZ4sKMdnX
xGOe3sOHo87FZtuILyxXzHdNAFN/NRm38nD3gIuYnJBulll4/V3UpnIUOh3Y
ApyATA2cLTQesKxgI4XgKMcUdwlqRyg9175r4WEsLCb/uQFxzZOzLnZGfaBn
yiPyamqzd6MeUiisllj4WaiPkfdGQwvDVnXPWQf+rRGcPnwehlTjpDKr3ICs
MgB3iWd2w9d2f8xOgySEmFWAheyHl3YeY+E4m/j7FYj16D6dyjQQZYSi29Ij
GvXIXqBF1Fe7Q7a1lXE9fBKWWBk7RkFdPX/RZXSAvvbTiAdN0qVuf2yCA1vG
U2ydBz4Cv5tMN10lNdolDc13TxONJq30JgR/cO7An0/ba5RKM7hNonn1mkMQ
wuWs7//r3arTMsebmv63lWQx1PC5vUQ3akqST7xFWsB1hheo/ur+LNlR7Hhd
hc23u5Sd2kWBGuv1DvHCsdkdImmDcV50/m9rqsez/kKkBo2wTsTFevzAOpFX
+n2Q+5ip2FZH3uEgRxCUFm6+/fwzGjryhvSl+D7ZUe+Cwtj3wO2vOZ699RdR
/WhHtHC3UFBk7xJ1bSY5ueCCeEsvmBgsv6rQ9u3GIv0UUdoT4RFtl69TZrfI
aBcHSqs9er0nF9luu8azhW1OVDKBNKMHDfJcSpXHLCVhewUUv0rrY6Dfxv75
O2fVzMn1UWX7vzGKU0bB2yrXvEqD2jdZEqk3dCJpScwsJWRIRUD/N7xPjnFM
SCKLSJkNSB0Yhu2mjZsk60Nef5SIJRXSYzlnbUswpgr9P53WNEMdVXFdfQ/9
ia/0a6I8smL4D0nfYNCHMsRQvP/+k9EWfVJ8jJRcYjqtcFmTT9dkgXF1LTWe
Z7KXhYMhVHUo1TFZxxV/ogNUfWTWImWZZM5/7JUfF3I0cr2w3C4JganLkTAm
2I/F7BdziLpudrLMFERg+cLCo4ITNZFpv/PxhDsgfcrQTaowX34iO6sUamB7
JbyvmuDXXRuDoFRI5mLCvoEovep7q+Rx42kC7Jc9gQ1DDuv89Q2Wl5nB+jhF
sbbeerjpn7FXE/5I0BhWMl1pf4nEI7XwKFMaklHPUNCDhdlVn+Mp9pzvaZkH
pchNE/Slw6lyZ3NhnSlvxLvxr24+Yi/wV0bZQT1gvS9Xur/Hp1byNAUjbMMz
q7un+g8cg0BOxF4pxPtTDPU4+fhljXkFYOeYnoBzrHBCKfVJO0APcP77oUqu
XrNYDx22I8hYQQuxZkcWGOzGgicdEFDDU/UyO3Vak300h90AIH/C3dyrieO8
kmkTvOBxJwNTlruJdJ70zKvRXi6MuPLeHmn4a800AYfrnOuECkkq8iJJM66V
OZRfTFCCxWJ5hzGY8k6A9ernEw2CJTjJhYeSLrfTOlRzy7aciIFDW0+wbBKR
zAWGaKsQqjDnRghnoZGKbvQs+SkzI8q0cDNV48Mpo+mVphQZ+KhyUlprjPF1
zcXwyXR40v7CS1Q1e3Yu1aKSXmBu64X2Q63jNxSu5JHchq9Js3k+TG8LME+S
+e5BBvP79V3Y1sCyVUAIqcBokXJTHdODuan4vL0vn7rRHxZPOS4ATJMmlwHb
sCFFMPGvrL1YXoWs4MI5VXr6uYVqLZCJjKE8ygr/HSixIAdOnVrk2E4f2qPO
mH25mcoW0rE9rkS+CvEznBtlRfyNhuJp7XjiBa7rwkOtO5/X9V9Pe52D6Vtc
oDD8RzoMhTvFV21whqJ/rgGsC8zCRNwNa6dcTIyf0WT4Oh1HsrRjJVCSk72O
MoOjm/SqYTbUAdjVxsmG1BcutrXJYaULCWqgZs5aRH//r3J2EmvcN//jP1YY
eUZFTVW3qN6l15Y1pHH75knq0DkFxi+6ng/QXgI/XcLWk8qHfvHQbCwJWkmC
Bzx/Gzvqi0ioa9TbQeesQ7rGQurY5FnyaPRMcYTJNP17Kivt0bLwveodtlFY
R1aVdZXvnuUVxYvPlC5uplLaZ8NQZO9gDA3sxpFS7OipJL2qtn90c8fBQtGt
T5aWcC0UW1N7zR9ROGDXy2cklGnteCpHzM6gUhSfjv2V3ULd5dYJDq0GTWxK
SZJwo4taZ2YY+/SlScjX+PkBi1hT00tB/ow31nMtoMySoqf4DH9ypL7BrSrz
1YAA+q7GvbqYl9ObszKHUocEQvs02opqeO/lfa8SHvyFtMWrxgq7jt8cRWpp
mfBd2StGhPGE8oNRTJpdj4jTDlpSX1nLWzAti9dBWQ08vTb1S+HL2pa0ldOg
itP++om2J1A4MEeDoxld4R7V3B/uQnu1SXBDSnek+27jn6Xxl45PUkt+yV3x
KxxfbpgmtGs6A97y4OH3Bjpp+tUHte60wKk5GS60z3XQzNb6jBkGQ2fYKGL7
FwrxXzar0FOMghCgVbg/UEGaWiSDOhg6n6iGd88E1c8Q1zIW7QDEozndqDVS
92yELKJUZWuebsYF6KCE+8dhNAlJ2ezIsiq1Vnb4MScsY3jWPES/gnuWrwOy
A9Q1+yc37kODGDpIJkM9N3MUabySnlfuDBrgKICLGmlgJcd1kbeDVEkXUJMO
soicH2Ma6C2HRRCuKqfyCvkixSWqsMoJRIGLeHqWr6+/qax2SObaD8JWJmu1
bzYrB0rmdi10nqXJpsxuAifrU0MI6vNO4+X6+hIugXlSJBOQVfoiUp4kO+UF
gUvYe6rzIDLLWSeeYwblz+KZvcRo+viD6BjXJkDGjKADlGRupR4Kdfl0Br1h
uCfW0YsoOnVNq4qznJoVM+LC/4lGm7hxfEH7Lx8uab6hCN1Y5YpwuI+kRJdG
r79YGADnUDO3d03xXgwXPeEz8sprOFtVLmTiDTuYySykiXppZEuYfZqyZAiy
NFv3QUTk3f/Ojce3IzkMDTDMoT12df5a8qUMdkx47WHe9rclDWR0JBZm1En6
mdKNElvIcWZsxSqhBpAx8DQZn5wc8QpfzxDIZWXWflhluLPjH8t2vcFPJcSz
ZH64qeR71Qo5/St4kwd047mT58WBrRi8iZzKQyxT9TQLij09Tj/exk060FNj
HxHUO2QdiLcjEbd0kbzAm8948wv84rUKPOCjOP/EqrnLtyCIQSdiveacxY8v
s+VDw9CjhYVdQCFAAU8a/18+rPUPv8KAW9In48E4ggcxPdkRhDXO5dKl+89j
77NR+pNkLOZ2X5ucqCkWsvLEkl+v/16Yaw+tkniyVFtTRpvJND01BwSUif9D
HP7WrsrnH08Oo4KIHneOpRrTEHOh5gHa3gzoAQuQPX9R4QS6uRfkYTjboSxf
JphG2HSzRYsYu/bwqESmHAXFMQ8CHQjnm5shpsmpDwLW7DMaEt9PPCqpQ3IV
+J1JoiHN6h87kvOjwdbIVtJT1KvTAQbf9V3O/6ZFqmSkypyot1o++Dc7/e36
L2MIBqUBDMyc+iC4AWZiqHb+9/Da/QRnOAyKJvBc9KwUL4la9cvD2P9wBjwW
wmcKQkxEI+hT0ZFShW0C9SDAx4ZIuJsRpdZdTIS7nufatlLAJQx0kI/E1wQO
M1uiDiccc51fFew9alaN2Qse7v6j+Tys/3lY6Vm5tTQlTaiNdo6xvjNw8ZCF
EGgajme7OxM8dKs9i2k/yYI3hrHU/Fd8u/HBcSfZljjhS+NJi+QEJwVbGoXG
GuSZ0DTddqXbch36GBzqkqXCRE2Nl+epTxlaLqy3n6zCWBtxIwcRaZAyBSfN
Za1apNKMfMp6lrTjW9XiC50WhrbyB4vpxFdYRR01IjGpNPKAr4jkQ2Wx6Bp1
LBk6gsWzOlBtmOKfGv3QpKNUabhAMLBQFMu4mVtvPWSq5mEWpYObAJItawBO
2XkgeFkYvGkQbWbi1gPNg5kuyoxL44YFjppzjSj+9sZnUEyLq5e6Gyd9+i7s
/xDVlfm3dxhPxkFNTZdyfRJSU+j1S/QrC85Ko33VL54PsoM4fniAM8orxshn
US4FzVjFdhgJ+8p+uTEwn/tibX1MwKQCB9G/q4N3GdBfleFC0HUZlaxoy97x
nFFxTVMjlI3wrRlqpa/FBflX2jq55WQviqZniAZyRvqbmyNVzc8h+EZV5CYB
eHhTOlkz/233NqeyzU2/PBbono98k4WqZKYDBkr/QrJbl7IV78NXZ4vZunIg
RzEm4s1/LeAIfkYVPDOR1UmIIKSmzYmgOBiKqLmXA4XVpSXvCsJ37hq5T6Lw
Fdy7byHgrpoG8nEK3ge+ihBVlb5viRXgZB277STm0Z2Igro1yK2GPzI3VTc3
MB/L3Vf1yD1FMSLzx0sSrTAiJjUFO4R2iBu4Uoe9aM8X+OAwghYEty5GUgvu
6fm/a92s7/OWeg0SJuIoNv264Pp4p+OJxR1vivmvOvl9KoWQUSTY/JhwNamH
Qe75fn/V7/0kBHGEwboKcvJeC35TuoT5Dqp+QsaY7vu/YnFB206+QhSH06IF
NvzkvMaH+OBMlI5BSyHEeQQY1JmpJcWGLsqpnSLhQLTOjExPf2iW1+OhlVe5
s9XePe3RqBaYxw3k0Z1ilW+f0EVtDk3qb3dX58kOyCWFLiF2kxkF/R3vv89b
4YdItqCmYfZGozugUm3vuzaDu4YRo81yNckLPpbgmihhtIsR8bcpSo9q+31W
8B4O253N/cPx3A6cATFHcWMjVvLraFNdWSG6s8KoClndGqi+64XoKi/5E2vF
Qvk5ggFKpTzUNSHUyUVo9mbMp83s4kUbf5EGdc0i6FSGJsT05K4Sff45pnD4
mWM1E0PFUP2dXB65ae3SJBHWegj+qMZeGlyvJRb8uxiKcO13xPp4oEmtC5Mc
br5E/uMEE3JX0TlzgdTTjIwOBLLUEQmReMVlOze/z8+oShXnCDQMjrTy2bob
OxJ6+4H9A5LKgpK9GiYHPtLyTqcaNRcJet45tMc8rHnca3UlpGCaNheitdM6
zPyVdMewI0SgBr+fzOg4hlPkYBQKdcZYe6A32zGTv1U0ZdA4aiZC/GJH27gm
Gl1zxkV8Nzmz3TpAhwLRC+LviPAIw1qAcSGtUwPnTTwQkdeTMNFAgbP7Fi4j
HUTfHCnSk2FQspQeILuphl60tRvN4bIBA1e7ofCrxG9doRRpxgvjUrvyb8/Z
wM5U349I/NlzRkkzrpF/IsAhdDHtKfYXhc2N1UliSDhVm50prXd3xGo+rGSE
KzZ5EdQYKk40dkSRtDUL9fH7B3xGmeBRF2uSb7YAUxqkTRUMbrvIhXIVA6Bm
OW02DXtJaQTnoM/LHlntVmv8rZ03cpzy+ZR/vwalQ7U3gc1hFOW/lLRt14zh
bWU9RDhqM5oXuyYCTUlVn1a0DeZsQAeuN93v6Z3xqi0bU3ZMOsQ2HY8ASd+j
v7OlyOe5z4RwbuSnjG4Qvx4qNdm1fmA7pxGj6yzKQcaApfNoV00LAfmTdCNe
w3I9jUVLHxhq0PEMVPbHTSrGiYkNtVyiCX3cJj3sd8uIdPXozzLIHuqgKrxg
vUvmg367fSIczAzHOjg7C2Bcr1EdtoUwfzZj57oCFQotOJECaMz/ne5TcBeT
e8qnwJgkjVjdUfM0s/MuEtL1pCYKWlhu+E3atEO0JfnPz4IKG1mhKJnhIqAR
Qq3v/37zfGKM+FNo0aUObBMR2llztVuXoXoWX8S3u5aI7p4GYpaBR/E9R35b
jl8DcSRA03luZEelzKQhK3SxWp2SzmKAxoiN4CE8P5hKq3ZRmrrko1PHiutv
46adTWnBhCj3SgmYTXRWksAYqdYk+2B99MDli/ITROKTWzMYfXmCYt3MKTDV
qpxNj64feEYCNt7KVbKvSO+EaXvqRRLU5/j8wrNUWKFEDiwPcqwEkOgNk7mO
0XdhB0iL0OvM/RcJXxANScqk7I5yJthZ6JHB3rk3Vm8zj7iSe6H7blrDwl1s
Qr6AomcSleEiCbnnu8+3PvB/xI53FBGheDNDPId+CZlOEBfWzLI36LamyhLV
AwV0jjT+71VNNmVAzEXJpf8L9YyUzJCeNKsZL0wwqsJk23atKME6gN/03iOs
B3nA0fyjx38C2+rweVmMWQzKPgBmQZIbEq6RnFzM4IRpsvShukCrBpPajSvd
hjuqj7Dm++6/2cOcanVttEb0zp80d2NPZ0D7I/jfTIHaaFBRY0kpV03wiN8Q
883TMphXJ4p5568jGF7K013taml0x/ZiTZWFd10fMOvrsOJnLgJyO/N22d8z
gMvXOwo3sKS+tg20NXp8gcfZodEvzB29cGIycbTmYfRo6qAAYn9rMfPJ7AMR
7R+SgmjaNK2I4ShoriLd+ErkMHy4vSlvz5aKG4Jgya6CXCWgn7CdlPGqWc1x
iL/hpNs0kaXwNJYBAAzA5wOSnqkOXOAJpLJXqk5/vUD0/bnUjiqko2duI/vx
EGGwhYG4UmORyXGKVSmQNuBUWF34s6Bz55xM07+SD2RYRabH00F0HksP1q3t
6tD6r2IEe7DnBDPccPWXIlgMrPOd8KwLRFP0UeY4WS2r7X2n0jD7auHaTZj9
QTqcTavOTu7r5NrTa/uo+rYvQwgdJjKK9iHB4XmkWxFmB80s066Dlt2SND6V
NCmMVjdSZRtZJuqbWLu+Lkukn/k0DpOaNnr9gF/1jyAP6RVEJbm2R/LKl7gD
PW56BK+YpZhr7AN21Up8T+chBhZvQ5lHItCdHorz6O+JYm2xVtplk0aI4tLi
GiypbLZG2WD3bK7xrCLWdRdht8L5V0T+7YIJmpSmhXZb4gn2G7+1dnJSjI9P
ON7x5Oozl3IT5pqXOQ9HVxKa3fBLl7PFPdqDuHAcNPIed9aJoOylutBtGyoZ
6oLUJSHk2hfKc8QfnO4UoP5+D8w7tBmUXsufV/GZKOmhbSKmKOa0dhT/l4sp
g4/nhPXMhE5+E1H7v7rFwYzXiO16xu8yXgxi6FfBhWy87yNZXd66FI0mHAu1
3jXkDuq+V33iLFxlpo6R+IEfo1mA22CtVe1MbWqCzc8aoPie6XxduyJtUA6j
VmuvbQg184fkBlIbIGUCH+Gy68k7gtyctDw3fgR79fqIcJBoBjCSwgsFkz2O
6MMGUlardcpoms/LGM4oeIH/yEeSji4aL4D6iCgm63KXIQHUSoA/tNLdRZuG
BQOBXYQ9KFMgD3gH/b1kysPtMAsb+wMiyNs7hf4eKP1PRXneD9Bo2BOqM7t9
pImtDx9zV0hjGAUQeTISuFtqCV8+E5SqiMeVqFX2bC1fIql/5K06si/KSKfT
v00GfoPFZ0pHlWqBHv+uPsQnXMwGskw0hU7V2K3t6v4Yu4c35/RuqdXQc6mw
J59uMgjFGt/j7V0g9cqTXswIMwVKJv49y1TIi14V+fgYiCWiPfbWYARgJlbY
EioMHAjQB5TSF/IqHpC8etmAOUKmKp0zYths8DDbjL0HzAQkxytoZv3j2Ia0
Y2jRPDwe0ozmxu59sbM29aBSzOHdidt1BLMkdKC/LdlQLwHNLqpz0d60/qEQ
m2YlqHXwlHSrDmCKzLCS4mEgnUeKPpDsNAssUKcFLcjUsdMwqJHiSx2lZ8Ne
bVRorzqkjER0etdjEFireFXrtBlSpKa3FWeKstU/CORBM85VfVSyu+QD/xjt
elMYd3NkmJoMOl9XO4WmqXTQ27SGV3t8K/IN7vaz3s6Dqf/oqnQ3eXTv/wB9
xmUFQ1f2VG95ww7bxXh2qHVwlqOjVxw7cVX/ACq/lzPc0QFvqXbiwPpZO/w4
gsgbotjBXYD5KSvTuGEhHFWXNHuks0SB4sNd3Ndf9dnlakNIapFvvOeTwJX0
aLKZbugSJpQ+pytObZqTefFejDxwaoJ+apVxB3gnKtF1tvf1WTLGlkM831sa
3nlJtirFkcJ1V40hD7I8XTFfyBmUXGQ7EXrgmI0rBxme8UbMRxVXnutIP0Wo
ptBq/k2/QEBY5hb2xdEogiNn9KJgaIvy2TSejCN01CqGbBnDoMuvSMlOqHFy
MSfZ7SOFipsR7D1FEfTR41eXusHuS9fQpJS4Doc6V4YCasJTytg7FIHKI27p
97vMxI17WyW85xxbur/NDkEyM6pXdgUO/1j6B00E/EtLfDNOP93MeG/tLa7W
xqiLf3QP9Hms7XmN0hBcCJ0Nu1iu/W9gzFxq+3R7kRdLnwqiEeKhJWXN76kL
KeHZzPWpK4mbNQVh9ULHXEqkCMo3fCOnoVHxzQgbMJuqHk3MyFEV6CawK/Rw
nZtvR27QrHqWdMB8yN/6R4csHKVpEqP69i6+QAZLgM3kXKLqWg9b/FjmELE+
45G5VzgPExHE1VXuqXfrlLDgBuigk37M4NySMlZ0BEH6+pTvn9Mgg02I9wob
OzFRN1UY4L2C6vUvpb9+xa1HD6ygscYwA4X2fvdPhn3B3SrtQAP3TxJK1eYt
6WHnrf/KkJoevAt+zJr4lu2fDT1BfEmNiXr+li/3MZmYiZIueC0ICpsPMLVu
dtD4fQvguaEoHEpyesdBKFXH6AMvyrct3WQdaQI+fRazvDO3ofpZlhGaJg0g
SxdytEFiDRrT6SUZLtpN9J7dtp0EePdyRbC2gpDq/u0iCohRGI+Jt0ZfD6fr
Mfch1HDhOC6L0cQvySaIyjiZY6EFQHgcxIWYPlsxY9isNM9Bc2lhT7Jn6QzF
5l6pZ57D6t7R87zOYhAblo2B6yGSoy0jMBcbPA96hdXE3wrNysEL/LXZ/mDK
/C6tNhG8+8Yux1zgYnXASy4hh++LrcLpsgUUmwfoGZnYwgz5BdPcD70KiysM
IWyaLhqeEwAg/UhFwyuCor+qnkrhXvJYASC39FiF2QJBLMzFuyX8bL1w/a33
jXLVewnJLz51bdbEjBBLavAFJNGMluv/o/oQI69iOhq0l4WMt9UZyYewnvBE
ySqIXYrEGWW2YfgNy+cY+EQhjb1zHHiB6QjXBDuu3yeo2jId7d6BCrhA8n+W
A46v4WCB0BuudzsnptgvE5g5IBTnNFay0iHvKXXlC2NvcDIGOjLVUu1v94vN
ExeuOzfNokzSK5U+ZPAnzTdcw+N92keKMIIoHF5g9JnGX9HatMwwajThmuL1
aA5S+fKv6iR8wMOsXpvqb/jBKQV3/V9dChEUogYgHnt8r4O7gCxDPAVX1OXT
ZFuRfKKD5r95Ob7KEkA4OJxfgZ8Y0BflP/72QX3p3I++oz3e6cheVJ+u6lw8
aZEcSIcaMPS/nShxbLdcQIG6FMMZoVG7ZBgaGoBFt0yfAw5pqsCKkQVHwU59
QI3ZkLMM1HxPfUUKEpN0Txe8uFd7/TTx1dJO9iAgFco1moz4xoVzRPz2wpWS
32t2dwW4sAAcjRZVdaxnSSDdG23IpY6gGp3cU1Ir0uQJUaogy3LZlxdVCjZK
iumLWXBZG5C/XKfi3gbvJ/4eKpF8oSG+/bLK6xaH0QaGy1Is2M/4BEuTikF0
o1DmAJcwFUtSA5B95N8afuPPga8oQCC/Ub+j8mFUKEqZY7Zc1xXAoi9aviqG
X/wjWXZbskekYB5tmZcHG/a3hyyBjariMsC/iCHQXvyP5t6773cwyN+eT41H
9BZtMvLYyoXCHf+uhHAVfqF+fEp/Ww8SNGSqAq4bwBTZlCWmefZWTfaNAutx
eVqcbmOwtxRZycNU2Wi4VKbwtKPUuwuM2hFM4fQehbt4Eu4F40wXDclLU0UD
rJBgV2vqTY8CMBdr94aCDwVU5ti/ya2RuprowYRALL9TO7fs5lrlIjNP2LEC
jOKjcIzSl0EHZX/VNfCARhQ0XcnLqsQuTaRnU0DIBLddnOZ/wqnRQjKi7TSe
/u2fP9BU987kqRfHdgPgzdxNWsoChjHAVdqBrEpYm2Tsr1P+kM7F3OlYfJKJ
yhcH+4/+tRF5VFRaJDxg+yANA6nxDx9UvCNrbVF619XkXYSnGAJQCaGtZdMR
iA3SQU1pdti/vQcHVM1jJGeNJoQUUKQ59dWUelR0amG2MuoQWalQr+PmF7RW
Dalwd2OFVGBxKjT6pD3VEctYdrRsLqinsHOscc2EcmXb5OuOfAW4TkIw6bau
KAIte3x4MQoSR4U9uLwFTUHME7y9tyXVIIk2ANamR4uGGjocKGWHLlXb5u3W
02ivPooNydgqyv7AhRUI3C4LhAUHLoxPboetb4/TnVdGIo21y5xh+95CfLcQ
KpcczEUF8n0bcuxsz9Q5mYoLflbFol2bbHYLL26SYnX3WRpZWzGDXGIqAtFn
yFpHdWB8QewM0TZqsgLBfq+v1nt+6scj+YFCoW5QoASMwLxKXVRJGfBu5n0O
yU3l44rjoppUYMgDbDKyLWoctCK08d8EoS7uKJumiL2Oxuo81FFo9Ekpf4/C
dSgfZlMaTT7OwoDpfge1mDsP2UQ9HwmUBL1bIM2mVZgbZymT/MB13IOU4KXh
5OMqBOqoZr/qJIibk90IUzYhZ55uBKQ8MHuJ3Jg8W7+ESsv0LnODWaPhEHd9
f3u4RQ5sNvSsUdq/vSdBeHQ8gUuQq598pDxOQD2mf1DnnHi6iyXnBkwW/bVO
yEsZkCX3oJnhyk0LGGCxvcpFqhTsmRC4joXsQgKLJzN/cEK3Al5lhMZvCfKy
gdhXUSzOotEU1ksYOvAmMG7SW1vneV0Bp5Iw+NE52lJ/P7n3vnshLcojGHAX
wtJwjPoXUQsLN251y3vvYI/A8PspzC31xEpp2BoYNpyd4Urt+GyPjp6xqfW4
zx3JpyDGRl0u3yoGmSkKmaWPYtX0T1GR6toyIKKzQ8ADozMf+N7O98nFncLU
jM1Mhub6DMYWnEGJ9sS9bg18lM31JP/faU7l0vXD6a+bUA7Q/S99Kni9Kqi9
jejhFt1qSGXALQ9ME3IHAoyIdHvDUgvNy2sBCY1d1tqmM6/+Uk2JsrxIwq/G
h+DmGLitFRl6Xdsy7Iog7a1hG5dQ1FSiyy7yLyOv/7JbmfbodF0sHHIgH5Yi
0tPozzOvBVsGOtt/0yGTZ5iwdeAltYQ0BkjXwKBtaFWXaoCxldd78aY1feH7
RvKk3ttxRg3UHwUoVr+jRZXaYhH5sH9x99m+pmJo8eCebVJ8bK7ED4ngcyDj
nQ0WrHJfMJ1lZgQBXM/hmWtjaBvsiW41FFpXs3mheKhkeKd9O/syFKqI3dnw
txK9XHiC2E8JqUJdx1fALnTRlG1khqlkOkP1hzgDnR01HmsBBXm8FyIXVpy6
vX99+/DnV9ollqBO4tjToih/9vOojTTD8elrUC40j9Y+VhRVqHyLvY7kknX/
kbmW0CvfvACbCPjRfbhujac1EmNLf9i+oZ4IVw4mktWsPPnRBTEsg9DSK9Ha
NdfhZqMha3BDN8GwcusHo7+9vWEQDI6aT0Y3hj5Pk6fuolTXlcbU+6k585ro
w5xDa+yIVw6P/VXDzguG1CB1RV3xo08cR0hwcEAft5jmJ8VZqQg0m/sicTqT
rkhfWrs7RCfDuE1s1/WdbSYGqlg1ZZGBy49TtExwTgXGLl0Z8cP8i7xX/soA
3t1UBzBAN58bAKr0Jzjvyefzsm0SEhV4MjxtvadBrGIeSu9Wy1sukGDYvv2n
9TM4aAvwuqFwfduKPZqqfUMt9wgDL1qavjObNByLXggKRW3FdqgLh75CH1l6
UXJ8iEWZVe0DF3WHLagSwaS9KvZHkzWBCwqOa7Hz5JlTmYmHwTt7nB46fcxq
CJmSeBi1V09p4k5R4L3mHQK1gRlRYq2m5GqSKCsyyPvpNcqusPpQV6fra9h8
lIp0374h/GN8d4mNHnAVhmTKNA5uFwDU91SJM7z74pa1Vh0OT0wyPge4kRpW
UaEXgFt9LXIlmCzYjYOItQ6JYefnRX/Umg6pnvoK2vcASG6d3Y67MeteH93t
QON7Dm863Yj/CMIurd/+77xiyRsuVTsWG1Ydjwa7DZr0Ec9sCB9taj3Ql6j8
jmt3qhbpVitrJDLZpE8JG17psBZpGSmAECP8KRVd3YL2sr25blNHC/6sH63U
wVL9UlMbvkUjp9KehfiehhWH6SKWOKUlurfwsmdtUbydWgLkWfkblnibEYlL
hAHIZ7KmLZKRjdOTNXY8F3cejzjtvurzpT03TNaU3JmJdazqkORCHU4a77gQ
1TothXE4ZZ+I0MOXJhlNxm06f2n82Ez0I9AECdOd2RF+H3A/KNp8c+5r8zTN
gXwQuCY/nmQKDFg8SYpsT3DQoWT8gIlKwLhPt3w6cRG/Wlf2iALZgyQF8cIC
6lRrR8JwGhO15kOA6/Dq7Oho8PvhotjOq7FI/NE3fkp7MoiYuuoMta63BZ9a
gI94sMWfZZ6RpBOJXeOgaBqsWlz+ehCn+llBCQTswA7g+Kxw85+2vLcxwJeT
M+3IP/HJJn5CVr3c8/P56FZw1CnUGGk6BCk+7Ad0gUQkJiyKQN9263DeDDEZ
4Xee4qTpFuKLkSA+OGTsgMrcEK/cxqlbY5zfp8RlkzSJkQW3z91rL8Sdqry5
QxrqxfdR9Qq/dtYpXf4OpF0Oxohl0jAgkC0gzqhkzfQZrdH8vewQyaWGdbVf
q/kdQ0LMLbC+4B8Jv1Im+eIiTiQZ6rBXo/vLV43j5Bk+kfsOToW0Rdt82j5k
9BPAZXDgDELAlDl5hAB1z+JpY75bYuqjWelcOwRpeVAZ+DjetynATZkqPyJg
78iT64PLAAcAxULb6uXYublJy0pHuXD9IIbFPteexdS8tzKlLrDRywQ7YWng
/EtC0dskqidkIoe+DrXupVMYMyLaklWAlnFjMAL4MKHSEaoMGnBHU6VaI5YF
0FVi2xVU5La6xEWd7Hzh7TGORT4f3udOBxD0HCAg9w0l5WXEJZi3jVJXWFQ9
T0AIg3ejgHQXznZ4d/9Ao+zLW+51Psl0VkDm7BtuDxDxwDKTavXIDLziJ14y
RuxQ1E7JixC3voTyvVbpuW59yz58OTSdtw5qXib0KR6st6bYqs+wmsQZt6U6
Ozdp3AL8yZRFgB6xfyy9VMzjYn39avvEfrzr5GGe6X+SzQH8pMPekQF98M/W
18gQMisCEiO0Rv7YMRVasbQeFP6WfxPEzjqU8kJDJYRiBpTAH6DnV+M91rP7
gqKIAoEkClcoVHgTMkVqH0v/Eeu6+/JeRZYrau+13lqEsijy/TQDldVlu9ht
tpGr9BO2AY+Ak/uv55LHbIWB/yJaUtP/SiWLND48iEns6JUdE2O1QHJ30f7P
XKebWUvwP8CMVTKp1jvZ9YTTByhKtzWJxk+tzjpy7icJrejlyw53aTKXXvXS
VILx1H0aJ4rXIhd9C6j4YIuxqh78sOgJ2Qh0qUdlpzh83bQNY1+1+aChATR0
lWwe5WsCPBzf6B0Zjd6cC3hm3N1uJmslF3Ht58I7Fj6KVT3zVFBM/zxDhkZM
45y3ynbejcIbvqnHN73XbdJtjhy224cYRchFk0U1w2Gv9VYHv9qpRyfvjlbZ
KvCgU8U39Q+O6DDZkxmgooLk1Ki2vMr9KKntSC39onmdpIVYQIEzmYOmuGmA
NVJ9fi22JzrpDZSc4kr6YvwwQdgbKTijeidl0mzkMEmCh/D3UpvnG/Cz/uDN
VgfzOIRSS7mcObQ8F7blfcktAQ/BRlEC97IjpPdhXVSQIjFIq/GmAISi+lSu
S+IOQ3wa7Yaw3GblZ6kVcPRaDst9cg0tBoTQ1B4aoxkv1gn1D/tS9G62ezD2
+A1wJudOWoprFIROUJ5I9g3hW679OtLbtE28zoxOrwCG7v7xU7fB1WlghMe0
8blrqVlxoI73B05Ax8/Kez63+K6e9C/2flbCPLhWfFOCVpOqPofs9pj7PDJx
NkElBhUct9B2qQbUoh2vBduaXKmKoPd1hLmYn6A/RRMch7YWpDV2FIl2SafC
xxsIPJWdBUDFORM8LRkxISnDn78dqfST59Tsb9TtUEU6fymWYzf9Y8cwmVn/
jVCcOAyIjz9/uMLC527vV2ipr5jU59ssenj9rIBJu8CKEV3vKkB4v9/odZGh
fMq3+3uRf8AgLh/qy7xxXGDtZhXoJf6TODRtacCM2RFgDuekrBI/i2liiLU8
NVK/NSTgSZ2PxAQPupKC5qY9JZQFqQO0p/7i8hH3Ex1saixzKWlwFdei+mvI
ZwFiFQUNyuLywfiolHabSwZptyVDKoTHGGAOvnZFkCWfypid7Rda0q2Vfxsi
sqVPnWwmYpxL85+H4seARvtGav6AXYZbEU4AkWcMZQa5OJZbZnCFDeLwU580
k8hvSc7rTtsDIBFMsSHwmaBOi6ACRa6h/rMF0CjagnLUOtdmmS5MJ4Q/M8hr
2CAlev2QPbD/2wQHzJhPvO6+8f93NePKIKHV6AnCOnOhsC1mN2MexLJXkhaM
vmLGGm6Ixqpu7LPEmhtj+If7bKjJHl+0jmYsXWU5T6ortw46QhATlJ6yWvPz
so52XKJ5kGSeOVfBjDhC8+vFAXPpOgmoI5UWDvLHkpO5/eeuX5Ctik9ttq0C
jqp+CbnOzjVBe3ECPIemR8fqS7//2WgSddJl8U58G19ozg71jRwshWxYqV7w
KnOCVsMOwvHBveFb9h5b6nX0V/M0upMRyCEhp0c+B4C73Ue9OFrDRjcoS/oY
SFoAY8YuMe6sfgI1+o8jHcbwPhkoX29qvBnrrpncrYHu9YPO3/JiuQCqy6Vh
4vVKt7ZyoyI1JcJdD/DNFaicUsZk8/6hpxVoomwBvInT9dWw/KWN8Rz5L/Qu
EzQo/anx/9JDR8sR9b7DWf5GXwB5BHK9TIeU220GcEElgTULORT+AmfnHxlh
HTYfck94301EgSAjKMFgyYQEF2pYP+Vka1yRmA1qPyz+WoMrIXH/71au8ScD
i/G8yLnkVEJRJRwXTeGEycm56P6Zq4RloM7xU9IdYnUiGeaZybn0kD2ZiO73
GzA2Psy8F8DcYvAwoSAOHoXKQ+H3biiSUrRg/Bm6neE0c8HCA+K9v0/LoT6Q
HZTPp3DjsEi9HpFKB25VWhSWUGNSnBRVhK0YnZyzvBa/wk9PBnJ5Z5iGZ55C
wqibIYLRjwkGL9NRGDPSdcUolkWf1g040G69Lwb6hWD+g1yQJ8r4E0S0AqSK
hPcUcRl1kW80JXZIAraHj0+Kp7erTK8DGPVsDf/HfTdgnVysIQbQOrQdfZsU
ye2yAxgO/zi76mXJM1RzUPjhv5rvCXrHo5WW3mx8t5eVCCGWslD0SRj33ylL
xC2gQwbkGPqrnScmKxciZUyixGmEhZU6i/gFz6bi8FiiIyaQt1g9V4Xlh1rU
MZpAfIkC7xEgvwwJbsoAU7QrCNgU4vmoqKQfO1iosvZdirYdJwQCxs96a55d
Krg1mQAHfjncnfegBoEmH9xOztQ4NhCizMd0oRlSYU2L40Ccxz9TtdZGYxJP
qqOptzfZ6umhOh59Q5bk1mfzogqazQGnU68GSVBzXXp+4fnVSleOiAqBO4gF
D4Oy+Czi9KIvOvobqsifp/fEteTbee8Rmxy0Bbw6SBO1u8LcUIS59HCcJZde
1Ss59UTDrHzeynOJ3Jti0gSB7pZeD/gWiOlUsMCrAuG1xQd7dOBU45K6JPJX
RmBLUunwiiW9X2c6q3P+0p8+2pFgv4yCaDQFf7SJ6GJs3scaJvK8G966peLC
oBIi7Y5L8h79mWnPgw52qxHN/hn7Bz7epCL85R86J0C/NWavDD9ISLohizmn
EKthQDDOtzRNOKMPaSL/JIJ5y+Hzol4UElX68oCnXRUxhHbQHBZuGYL/3nSQ
LnB4UMkzsxXGcc6IfOGF5k/N1fWCDDp1liRrdIe7LrWPUfOZf3M7js0WGcVr
xIQZ94th1+75qPMIt+x+zNsjG1ANfsjueNcF53bQSd0BhQ9GlIcCVEZ9WuRw
egVe6eEXkPsEM4ZgjhP2LgorfiQf1T8T1GCuIENGUvoOBhDD2H+8yIIkD0sH
mti6fD4sZisC4LhhZUa/ynClpQkRZdAeg8LWQTmcrJsXCXZquTiBJjP6wwFJ
q3Hs0zIRpQQtFjQfExApA8icX1wIkK3YUAZgMd0mAg2n27WkG8pyi1p9EprH
sH9z/zyrCnEvFPvsAnnO97N7nmMXyNeSaINV6h8QqPl4xr2wwMc5hEhONw45
f30xxBpYJVs09gq/GDa6c2yq/Ipcg8i5fySZct2c7QGhu2zxbOU9Qy1SCFxf
j+HssCaeEMx1ABhiOXuXdciruVZSOs96eCeHr5K415Qo35S+XRHeAHY9DMQW
Bb9/iiSfUkb78xfy4duQ1AJ5YK2kEaQjGBdUw8XzZGvigGiiLPRuOxFDkzeK
4BcSsA0GCW8vXxgwBBWCc1JL5xn3WyERe1w4XogVf2Nha0bKypsnhi+evPMh
Sc8gPMBzJf17O5+yOnDx12/K4w/WB1DOTALBW2MHyY2Gp3Tx/f38QHz1uf+X
Kvp3G5ZQOTeMVSEtHFqh1s4nmnC9lXQ0e7TX2EyxFrhRygDj0Qzs1ruBSd1v
7cvk/IG7cuXtfjPfkf3ErDcsuM3rLVwwMw7wDyWgdAc0YOPMtzJnsF4FU1h0
pd5CtiUWRQkffPJLfP22dSJGGguxasnVwDVntH5TDb8cJtTv7rNXi+bgL4L5
uzBPXnPcOU2mjDQvtmq/hu4t9YGpaG4B81QYhLdvfC0eOrXqmX5Jjr34J0un
hgF1ldxpbGWzTHVKD/M/PYWAcEqb2VNkfY0K8XjkilhtHt63sDHldKFzK8kv
hJYxm8vEzX1PtA7BYejKeFbqOSw4fyklK+5vkpnwam5s8pmrvV4HKOeqgYTS
ZgUJgMK6o+FeKvG7f1PxIeabWeNEOfaqHnBBWqDiVqN80zVijovJgog6PCj0
ygr39ApPlbu4cRoFbAz2ndlZozakuPefMX3hjkgRRIsjxrxbkXuvhUTR8gMn
Yhzdb74zxvTbF4iQuPK8K6uRrUaeA6vTMbhpK2krRQVPCWXJ74bWWpHl7WyG
cYFGLAcXIHe7EZxX7AeJpvjt1YmHWvJnw7ZVS+z2DkJZkJ/9IECpQVmWg+eN
ck/I7LA09rDhNEcr0ZbN+2EE9fnjpHDbynin1dyP6q+Sa8mmo1HReoppKFr5
q1ALJ1uBhhyt9usRBse8lyjmJzD32lAIzzz4Fdx278h01F+6X9ODkhWDQZWg
7jvJyDppS8NZ0/1qEz0BNkErX34tbxQwxQvH45G4h0sOOZmBBsAx/kjZGZBf
gt/gq4/FUeos+7oAfp0hVQk5MWBrxlw8/p9wCmL4qt5LkO022RxpM2V5ELiU
K0RTXc841s9/Rmqj0GMXVpBJspTaza8Pc2DBTCvSZm32Na2HWxYh80C/ANpG
8rtMojzzlQmA/06D0Gbh5IRsoARF7tA8HwUFLbJWrZV2H7gS/Xe6VOAKx8mq
tTxdf57XI0lchJ1s39xOdoM3VEc5Lm8E9q8QJftJUFiZPLci7yGJj4IiOq2b
F4HBZdKw6oB8iBROMqAkL+PfTwzpt9RItRLcmXFF0j53rzBHlK+DHwQpnQQ9
T4mVF7E14XctxbngDV8oeP94j+XyShyVZ7UkPfoPv90SGpyw+sLUgj+Nfm5C
8V6iM2tM2e+pZmu8HsXpb3gCBAGBI+EXtiIV8eL4pGndDU8RA5fwzmkuCYPT
mLAGO2G6NdNqV0HLyNC1klq3w0eAtBYRJW7y2oEccyGfEnTA/UZgAa586waO
GFG9nIisJwRoOm50iFMzrScbcoUyDpGKL3YZAV6DQl53VxGBbA+4IpcdFqCz
cZrG4RM/kIvcDMvhPqQc0WtMopf2dIasvySAOn8x51QN/a/N8CeLWwepS/eu
45NJDZzoLwGu0Z2YW10gAs3O5VraZhEHRfuuxL+mNo1+tGmQH7PtE/BvN8jR
5FMx1b/Dl+ITIt+pJO4Nu7RIsjErqDyzac6W2f+eENK7AARB4jpDet0TTpoQ
sz01CW5uRS4GhkWUMHlkNPaiPNAsAah6IRfsDcmmNCr9/k9X1Q7nkOtkI6ks
f+QuNf9fcjXNeUU6UU19sPkkymVun2yS4zpvGklrxMiA+SJCk4LrpMn5yudr
hBS2ZVqyl/fdILj3gyykm+ktT6LFc5KI3TlfDF3UszhtrusDEZKeGZu5ylWb
nM5sG16D4TXeH2e3CV6Qip4WZYktp3jKt90bX1LuOXZORqWYmcw1Pxl1sHwZ
0nIF57/480eawhRbQwGj0d17nrqnyNoRw9O8scPQwQvMvJDDutBejlVMr5Pn
AVXrNyC5KXinE4DjkDxtWY+S7zjdDsRiHAQDwagQtQAQYvXWz/ygCeirXgpr
ffWOAqkzsPfWeFlJqukN64jH48aP/8wJv8wgBtBn12Y8WFhJSbn8EruSbQUg
qp4Il5Npa6uHcw3zViEnjgOUCAUZQxpa0jFsMhyTXdg9VPxbuuH8hu9rdbhZ
nNou2ev34KHuEScG0aPLdvUp1QAduAnZ/Bg7UEX7zSP/XiY4Mc5gR+fqvjlr
F9KXkmvogFZd97WfWwcoEoNC7U8vnky7s+smn/su2OA9rOpwxT1Css8vYf9T
+HaaIDAsCJDiOANmdGcEF+cv9t3tsgIA4OF4kiJlc3WBFAE9dwA8KFKOVTf9
UfIKmsPxf1iBOTlXQUqSoisaf1DzCraEIdPvWCtavBcCMFlbR+e+eK2KEgqE
hwfNpnNnb4svD+a7SC1tk9xPXRM2wp+GWtt7YIw0MpltfPXZSERZHcqP0yTR
mxjLoO8lGsu0MityFvQcoa2Y74YCO4Ej5ZrA4eAyFi4pfngP67Vpxqs25nD9
/2nH1T+OZnqmqowaruchbuwqUXY5dxrnY92oWJaMyTDyifK6i8APtXW+ItGl
8tbthbDLMfJ2We5N1cG6prsZTHfnFseJVcAlLMk2PcedM7nrboMIYgWp2/pP
Qi+k/yctTRf/Nt9W09lLHXo6eQs/x8HGFaAqxe9RsFtH/sU8k9n0SMR8HAk/
L4XXxyxIIAE8boup45/kt4l7m7Pw9JE71t7lDRDzuUUKxSn38mjV6giyy9UM
MlOACCQqi5ipTFaBh91apzs2Lr8/lf+MBJbT+1eGASdm2XCep3FU30DeLi4f
r6ib+RYdIXYCvIN9+Iiz/u3kS4271US7WmjW6SAyjXhYrlMT4uEwkvLHlikM
dEY8PzpKgbdbzTGXvLli3wxJAKEc2vVlftYm3Z5ztbrEQqTNkc46dChoaobs
+GasoMh+KfejkVU1ADN6pI0OpABvDWCx9Yew78uFUsLqLOiTQ8hh2VxaQit4
1FYZN/5zv/c2fo9M5cr4kNApJMHGa8KqQQWxIH9T5zUio0BL/0i5Otmme6QI
Y5wo2vmv5Xjctut6vZ8yFMaLmEfl8NdrYBcRxKd2ZzegcG9JiYdn6nrDCNuO
4A7R5yIjw0vRRctjBJcoz+E64CzVRVLENPJZP8gnDp8100hZ/7IKMmQnWqyZ
1zL10bWRE3FN9VMcIARFOCm2ITqwlDBuRWfqfG5RfdZXxiDnYzDFwNQWjzqb
5J+EUJQa+LbE1P807SewVOZWcLF2hcMxcAOaSLGnNwL6T/FZKmJCiIXHic9s
PahWG333qKqlRglx4+lvTAqk9wrGNnTHx65S8SlQwC3KRHK1o5YRAhRjzans
D3vWYtfwbxmFCKfpMnS9XnzUA6TxHX93h6sNzGw77ZX4VRbxty74WAj8wjcf
tR7x4CvxAXM9srp7g8xRU9QOhO7peoWDu1aXHPRUvYQt6ENVde0G2zivxUI/
Vq/ZsVVhbYY8uWSsUjJheuw1eksAqPYlN4TLerl66b/tN0RFY2bDwFLIrkw4
kAjIht63t0X/7wWM3+LOx8Qy8zyWJxi+8hXSzGhNjgXFnyTa6Qg/xJqvFFNW
1GfOlihESdRHJTPyZ602RJVsz6PibRu8Mj3I6KspTKYR/W9pz4infX3SyFi5
L1XMqhbgO3/UHrcS/BoqXdeha2ifhZroDgL6keKpJokRqy5+cbfST9YeoH8s
sQNYwD5JNQP6hXQQTyfNjzBN8n1q+30IMIPcbvJuQyaH0PZIf+AZL9BS67UH
mzRGo5/XeywTZ55E1bTX3DrRgAwQ9aXoUmnFmc1+uaRfGC44rUW/BZQrdgN8
Pd3xMbA12Xd98JLlJRVKkewN3Yle2BlKaPiIsUs4HYTxB/OaKwRQUtt3PJkv
Xyrip32+FqxTDyzIRvLi4WiytXsoBfRNU2WHAaF/Gl5fRQ0FXXHX6o6W5Fva
ZVMqm6idwRL0vpb8dBd/5g6Gu/iWJO1lLdGvaCZ0wpNIiAnx51vwd4XviZN/
GcUeos8UV1TwM8IBFW15LFf6F9sfJnYyIWgcv37/mTZKF6ayIijhuNgzgl0V
paUiAlA1TUszSpoj2DtNSk5Gg7pVn/+VIvdaF2WLqPOjthho/73ByaReIt+A
j1YIXjaYG9rD90moMZXgeLJBQqtVEHgKKqPTWNW7cpupSZUh1+l6ou0ahA3V
WSsU0qWERTUJ9T9dRwMYy9gfLIIg9LuAm10WGBdNzXl5+QXLJa8kyxF6Is3r
TD9WrE+76bXuMFsz8yaSmgKtb4uxfV+fCfMonmXgIoKVMgK5zjVzYUNtFRKW
YCv/WtqMblCUCKTOpnF+R1oxAPKUUaBwKpdc8wjJppP2m+8QVWCSzFuAo+Kd
OkkdTEUw867ItNlx0WGj3TSVBjFiFLytiF+5e6o9DVCgSoJAAGfp4Tpw81DS
m136RLPrloFDDZvjskNpk2z26ENPkqCX4aWIeSMMAM2M3OZNq9AvOc9JjbEt
fu3ojAPN0O7QoZTkq4KfRVvPa339wDDsRM4OvWRX4hEYovciSM7tkGQhYn5p
DnyhAKyshajN9FUwgsJeKef/p//rWg3+7gtiqmWsZMkAtUvxEuSS6a/zJI/d
OWpGAd46ThvBxv7v50yrMwwWKD4ijL3uQeTTrQZd1rAZiZFUk6IMRNk+Job2
uqxDPVsYoVdwMZstVgFN9TGroRg5DBnFFQKIE56aXi+ZqjwHvHOgPXpM68I0
UIeoPtO0AsMNpB+//V/zVaBBH1Su/xORG5zDajNLYDHh85xRs19hf1+VsqRs
g5L5UnKXwX4JYDWG05x3Zfn0JmOUoR8wWKsGr/XcMNkDeOezqv8TDix3iqVe
9uBX3QmeB/UHXXbCQNVpx9CZ7BktJlwbIdIyceOIIXEq2JbGHP7rN040fp1Y
xQZvknQxVopH9CKsEnOc+3RH1BY1E69cQoRvNR17JZMakNsUOLt2OMZpWXt7
7eOepokvjbRiXII4i0wQ5+2sCN85CDHrNsUYytK2mY/D5nLUZIxNBq9vWD/f
WS3QIZG+/Mcb8XSnrqiTK0IvJMb7hicshNPMEcqbN/T5hYkWRNp9ZnrrSgXv
w98q621tpUrtIVqczHc57IB2lahflkg+DrmbjYU1HzDDnAAT+hU8/+exS6Ja
vW8Rdl0o3LlQsO6pTQRGEoS2woDvaNj1K4ML+epfGxij9UN2IcFRcVvy4ONs
mf7wWHCirCLSOscD7pDEun3iXfpTK6OKIXT6bJ9bs7DV5Wu4mZkNJRBgV2ns
y+AbkUtT8nEAeubyBxnveNUCIttTWMfyHAwbG6OTogAD/J5ToDmQsmpUsUry
AhVyTwT6G2de0XSuV5045LL1YYl1zwycHAIQhdh61Ra5rKa/2CdiikdpXhXd
CngPuh02qruhwrVrjwno/JL88zAVO4Ou1gqPvt0Wrl1M6s3tJSrkqvgtTBAo
/YqicaogeYH1r8wvUFW0u4/Sm5zNJoXtF6PiJVGj/lO+VYyJGaqiWfuMsxFq
qf88tbSVXEPGTMidByDSn0/c97ixpaPm7j96oSGbM8uWEFbaub0E9fExEjhP
VqrMCFunvitYddsdcexArikwzKFSKZDUb+lX1QCPWgg6CnHqRbpcdxbdqhW1
x7bSVKKomwk+cYp9fgsfyWETP6+4hb94GQTyt966tIjBK3zZNqrJxQufAPD5
60O4s7DZMTgRHREUZXs0bjsD6K6swmXsqt2P4lLUMXINxbPNtR5BVYdeb2Om
/cLfZoZKDdvsb+xDYazw5CIxMj6vrPBrB7NKau7ekwFEl3yHhFR7DqsIlG6/
Cnjuasr7lAEgdzqnXPcUtEF9vFG4rKopQWVuKFiLNORf2zjYdd14Y7g2T8LN
pREsrvvMnI7/AZaJw2Ac0C/rJVHgSYDGk1ZVV8ZngfjGmF5kak49vmRPbElg
j55X2QmC+poSV0wssbvCWPbp7XfkuBmch6gHbaU+w1IsZ/fpv/bEQtIWYQe2
l5ocHVThafvOjO+0sVCQ4ttTIvHFnZraLblVzFOi+35AHy2AkEEeZJJMMV3j
fYGJYJLDJfJA+u1QMKY/8z8zpcnMTatWtl2wBAV+8A0Xih00ERqqrCkzp/19
2H6o7uwgwmm9Evy7Se3O+CfK20iZ1YrKeSMYWf8Q+LRg1WtKFLdaPKpCb9p8
6A4rPapyigv8xD/3vZ3GXxL28gaM0QAFyQV+Zz2mB2Ty8LiZqd/2EavmJxLf
HZerBSivNvXZ8aLyTooxk1SgayZjmvG1wL0VHzZNZDB9ijrn5KYETh7s7E4O
wSRFIW4ZtBgNvikbgROYRxSJlEfC1nWX0xFTZiKw4uLYHI0SlNFgPh2lUVVi
B0GH1WOpWZyGM+FADEt5e6yE+x61lJcYTa+lo2uJvOGIANG/mYeJ1gP+22GE
jPp4bUTjK7GDHTjXUoN/hGAi9avdpZpBFydoMY4JAdQH5PfMxIthVvVk5Puh
1lpizYDBnkdR6bEq43/kQxjHF+E46a/+RM4Rd68/P5KXpeUkGXhOOi7hjRBu
ULkrht9fxDDtZ/m70F+gJFn/t+9g+yHS6qYhNwPxbU0waJRpHlwo+pMtA30P
i6zg4LRFLs8c97SZGv+QDOmNCCGqvl/3hAYIS46QO3RsHUj12IiX/s3Kt6g6
ohTPk84JQLa7ohhydgnavzpwGum/uscLfHC5oARBt/UmlD9NfBQe1Qa6l+4+
2y//1TmWV7Ni1OCWvrhWUPIhAPgyLq329GoJUpnMmuqEmeTuMK8Yb4R/5vGt
MXPtLkvx8DOaQ680yXoyOyy2k8/i8PSBrZvyhJgoWdQznX/eG7f8S+AAiMi5
oDyRzzYL/KCdxSnU6g5FYoHSj8vRTHRRTka7cue38SDW5Fk6Imzdo0Bov3gu
zODT4w60ZGcJoma+Ninlhc6Rwc7vLTZqZyH8Qna5qTYZ868OWQkDmzUKJJiy
/Kj6WR0Xc0Uv20IF6ugF+1yr5aJjdhL0E0VFSrcKir1mm/2zRXUl1cvDRWqn
9/ukRaJ4vBXnxkgIzLR7vJtB2h1m5xVMcmFo+tpxcDhSdG/LNYBQq/4xqc/G
4+g7Cf0KFGixeKTnT8VdLtV986K5cI984Xe4MduzLZVVcQ+HyvuUykx6Mkqg
8ivZXlH/kWkx2glB1Glut4YGu4sj5hVVS1/tdVo/IV1JZkeae582uB9bd2Qr
Bb0/r7acdHGWGypKem+SR/urwA9aRYlDAcCyMT1sd8zL93FOcVLw/VseQ0QS
fCG6I0Swy1gZ5c22W0RGfEg09QO3wtgQjStqcbOmyCCQeomC+cQggOsmwOJE
BB66peN+vUStTCJsbCMiE4/YYlCV1xnahfSyvPMDWf61ZQ8Y4Zuq/y5jupFc
tNfMZT4QJ5ZHFrBVA1XyrnKgiwCCZx4o0G/RwCFRsuGk17kpyrHJ8DJg2NuS
Vy9sjvtOGCjVvd3fStXSLcX7ow4lzAbEBoeI3j4xTvUqD5wlvO8Jk53oT+kj
IKBMTpVBHCYwdC0xc4/VKZFJm41SV/id//rJftaYI7UBHN0ejBAauLv76lhH
jyGaZnrIbe9qoCBRwEyn0smQeydUZ+q2DH7cnL3OVMbhLIucVM6qYrL5O6Cc
X8jjb0qVFJbCidL4ClSDQv7z+4tRjF6xGYqaJlYJR2AFyqohU043fB/kCXzO
iSne3SL4nb+lez9OV/sGxWUup5FCQZeE8e1OFa6OIwGt7zjo48yAMIT1lCZp
GLZeyaE7FS3N4cJ5nLEmhXSF2itbAhrhxOmvO6q2mwDthDkMIe90TkY3huvT
dgk694lq0xJZuPg4GP0jWCjLGexbvt1tUNAYs/jMutexirkBJU9B2twZe2BB
H87R8b8VA7EfpL4cW3H+Z6jnaOBwAeyJ8DRVK+JzDtfXJDP/vzgKoc07ZwpC
zkCXk5LmJxFTq3s+EiRgcST+9S5tgIfS++sLaD7neVi/7BuZIggHU/rXF/sY
tmeVtJsGnEL9t9zVj5NAPmL+QClU3aQv0AtIAP+Kh3YTTMutd4qsmPoPpb9g
jhSXqYsssbI0Rlzv2+uWzxhThVp2OlBIgC18LvRLUQfdOg72CJHvkQlbjllE
embK4P1d2/QTIJV2WAFTgqulEGdMPkFpnYealn950O89mQfo2mlKI6Rm54Zu
03muQwHadt4hMa33yzbpMNc8O9iCRVcpHoKuJ3J2LuKeAlHjbap+cwlgoKCo
eZbZHNSwgnKOmEu3MufbBfTwOHXnh40F67MA7bM0WzDIe4NQH6VBvqNu3fGx
8DLt35LcYTy9Ww8fOh9hxxUe+U0FuzsEVzmF5oGOTGfh4SZBAZwEbYcpC64x
1qmuaTznQJv3x07vTDL22nhbknGrtnsBjPSzB4QgL68HfjJa/ZmN3XvPVD1B
pUwVIP8tF4pacWjs/+FDYqKnUQW0apH5NL8jGBt9dUwHbvECCGOZjIRbnd0c
W5JGMxE9x8ZAF0tUMz4PSpEjW4ueVrG+i9zwZ81GEOBXvjsR6BBA3/kLnpw+
XYaPjb2T1vr0JSoHbWt6FrRNpPLCCVqtKwdiaXdNnWf9sBWZvWlFU4HR0K8x
Gy/XEGtoJ8p9GifvlUynvsovWsnkrAMr5CyUrwLM25iQqwJQ9neNtAmE30Oo
qJtHO+1jIT4GLD9B2JLpxM9DXVBwcZjNn/au8ypkbBJLIGOqkBPqghbRYl8E
yul2I6ugtCxbIgXsAK5oJ+iLXn5m65yqLpPpVpiC26nBgGNN8MIPE+IZF5ZO
bqlCcrvBPw701/asYn73x6UARz49ScfcrXAsjvdMpt9Ix8Q101m76m/KuXk1
kqauRNlHFwYzhYY/N1PTgcffBychMSEwnPLfdjzDkUO1neoQ0+4zoia33cKd
iL7YwRjYL8NFrU0FFyxIcpac8eqFCZcQ2ZvejBgvU8AeIkWkJmYd9LT74ETS
4jaXgorQxKGm7VBqTkZdYoa8fUbWGyhOe7c1XkOJOMWKYPk5XCzoUPoa39+c
4sZ1qa85GBc7ZQooUnZGRNJjXIoXo5UAPd+ZCNt65syMZy7JRrAUqXa45NB5
bgFr6jyifxCBNc++wsiVWY0o4ktIP3aFMK3xhgcRD9bjp2Tv47suzMvgNIv8
+cTNPPj/ZmbLEn9cjZ6fQhzzo6lyeyDfHj4voV9d2AvTtI0NlsaDXsi3u+bC
1LxM3L9taUUafIhA7G/kZjSpQziLrPgDqEHM8rC31PuAzkCWH+VBZBbC02mG
a0yfF4hoZJRvRSEs26SAEzZyPHxerIjRPSbSAhKIQW7lhml1y4gOxDL3Km6P
yGJNcYDBIsEId3HDzKSUUmCfe7nbt6RESPOgPxSK+msPyfusw+pAEqFvgz8O
mGSF4Aq46aI+kMP+/VHM9qKaRQg79TFXdppJqJi4o9cg/wHm2e6xOfBNt8aE
2WD4/12RhO1g2kSnhOjDL6m5MHBDqnJqys84Hdec+lNnIbjNyS41rI8KQi40
ts1J66YoGrz3TWXdldSM9FZpwZT4R/lh0bxp2cHpf7ROI94UQLNPZTIHQq/A
Zn8+fdea8B1THzcF4MqSY1d6+HY6V9HvY1oiZPXaPiYihiUZ+yOT9N8Q/EoL
Y506dYCImAuq+oq2rKHztaUuB3cGrJsp5l2rrMIuds7RDZY8LLkOHeqyD0+u
xK5fRHdRNERB8sRnR5/uWUGfl31m4bUUZ97EUOVVhqd63CoTACK+4QJCNpZa
KoYGsm2n7s/EIMZNdGU6+1+C7trOsc0VII0hVsdiBsrQfj1/TxYxlDIr/S1C
XmmdABJ7XkXOez6PNEIfagn1fV9XQMSruolq1vCvIsPw3bS5F68/AwB3+I1G
j6ptS5vkUkWV5SA9r0Lgj07fg5A15cosTaQFCqcxGh2Nd0AfCy9KTfCFRrRu
2qcREfABvsCwKwSQxgU9ZFv3kz6vz6mLVhfvEoEc3LPL3S6s4Q69AEW6yWsW
GzNx+Z1qt0KgVbHb7V+ufxW83I+Zzy4NxSFryYNIunUYmACxxLIIuthCf5Bz
jkk2vGCnFlsFTq4k02B7PGhGVIcYrguZPyzLZkpXSVulGOFylIWVAHx7h/++
4FY3BkQi0js30Nog2dMmBSFh5ck/M/MSxxhxvu/4OO+9f1mrgkT7eMpB8cdG
P10O1DVe9lu6n98QSFZBg76CmxlJWlAu98JeAHOPNuMTaheME8dqpFo54JXE
wBDGY4+rvRxNogrDSpSyghK25qNp9KPxwa7LThIwTdG/h5BCYxJIh7Byl49e
Wv6jK7XIo4xtxFFDb/X6xwcPt9DeEJZbISz7wde816C4NdwCrRAL78MHJvgO
LxgyLYFs2M3UewwGImxHk3twQRuWaf5eoNHbQbvIVLMd0pRod+Mt6nsTEqJS
7X3uQ34X+3amTynJrgUYnD2gOfH5AQNRmBB9/rtSKMJHtI66sHODfKpOhqCw
Q+f1Pi56qD5ZJRoe4AQIk9VBhx43K/etHD85siQGM43i2h8UN8sYaWZZHvhU
nBRijITyGRGQ/3IMrohNpdom2ylLeb8kn5uJKvL2PvHFRm1UwB9pt7KCvB5g
tf/mIs3xVCvH0WAVv7jXr3tosmhngGRjY3+wNBrgEKhajEZOildWyNc37uxf
iCov56hfleonlkGEycO3SfaBPP6SGLV46PSw8+WzQj4waVGrMHAOFaUQY3J6
5PZG97bw1uM0ewGAZbXlSW1uLrjq6f7XFnZUN4PXo/sZ1weqODYv2ytDGwjc
2NMuu0q6P8m7bIq9KVTTaRuUrfoGl9GZcPYT2Tjy/1HeVMkEsZM7LgUKp5Ig
VeI3AO8H+hoKYw96kt4bFQIV1Di3IqrvZZrnyVH7x27m/42XTOdrD9WBDDk7
FIZwv7Z7pXisRSXBQex/NMNLcs73SUbIbcQBH0tVdRNmlBXzmoba/mxu96Wh
okFJzV5KCKHH7uu+oBVg7y3C1xqxBIIDXx9fMBUMxVYnN7lhL8G9tqe0aKMx
fuRH6Q50jAc2Q/jDgzU+nxrUeBsSge3P2C3pooIeeHt6ufTDf7BEXh6QWV7d
D+LEjpZEGImr++Db75lMqNFLl0NKIYqWNYsmfFABFPJMs/sxJSD/CnXsQcTg
o6XRN3w6JDYhRs2HgF378IMnurQxQ/zQaL3yTOlcpv6I9B+WdZfwMjsk729U
WU7lQSxDaCTGgI410BCtyTjQxXvu/Dsep/hYfyp6vY576g3R3dcQGnWlXKSv
FawzCoGqqgbH2Qrw4EJwAum0Xg2h5FFihG9FTOB2f9h9OaTc7hyBMm0PbLJp
gp+LlkFprEKPkE6slbRqp6wrvolQvSIB7Whgo6rQwefJeiiWSjACNB8F4eFi
RfiM04Z5BCnkpCuof21L0WfrQsAeD3jc7hDhVNnU9tnydIvvIbYsapHH38Nn
9Z9e/UQGmfxCHoXuQVoI4n9c7qpWrWLEHyLu4zL1NkJ1+MQPVoQYJt0M1n3P
N0ljxEGaMZiV4BSJ2119ejkDqy5ktlcwTRcujlT6GDBbOfS8lbP2QkEAinyM
o1tD9bRp/NWTi061yQx9JI/FdlG1Zd0LYq6qL9YMmzw7te/KEISY+cc2ESoL
eNJ5XO7nUvyKzzz82V9u6RxOt3flKuqaCcqIFTq7QIBREFlRrJWXxUcU8beX
BLK1/FYpmpBRsm+kxwozimp9V2KMgJKZ/skJjKMA8zQmJRxqfID5o85NLXti
/gFyaBihB6yyuCn0/w8LWQ6PBs+HfBnr0pX+eU2x1xSbW7Z0fjdttYg5uScg
zkK2CX93IFO2D/H6a5MX6ULUTjk+J7AAeW0ScoOWXVuvlU0YdA6ao6M7X/5T
hFoOslOcnw2y+HDIvYpo4ZOrOS0+lKbx163E9kSM8g6JMqi8gicaYRvAJGBI
9aWzBdwTMtNAxIG4mZuFqPGBgiyFY6dr2rJDwe5Qfs7v7nF3MFl+UkfrLLq2
EqH/LQBRJ4FH0obYa/XzhRA3ZOwOiyZFRVmj51cbS67aclxjQVvfHI5THQ0V
aFcnCoaPDckOjaMvpVhtbMdCR4b8uIZeJaP5CYJhileBGkD4ublJyK8BMvSq
CVRItF9M8QTWkvcCy3T2V5tpD73M6aZgJdQ6vk1qzeqlXMYLq5itsAnqDpgT
t9ZSnP3gLnQSUO1+TPTKEC/lixRssiO9uihwFo6zSV5tbcpFY6yD0D47rhWz
4JmwYa6Y+9Ol6aPfda6E0N9xa8BwWKImhY9crev5g4m2xCFujcZwLQKTnUgQ
Io91A0NLRGmV2vvwQ0ZAaPqLsMdBaPK+7BBMyoTvLyjJcox+8lxqbDtecxFy
w2QXiI9MF17Ts1GRukVRWqiiQTSRik4VbxBz9ZLNPVa0TPrDP1yo2FcUYeKl
WwML1AovwQfypMwrGztjEALoleyPILhYahGEi1gPkY9V5AKoR4+PL5grznr5
rxdrIhWoWZW6+XQecNE4hlHvLV/cI5946/6q+b6FszG+y/CQ4pC06/qZzC7C
J0zTDh4ZgNhDw5sTOQ9snKXSsIbERyYihBhiRM8HZcEpbuXVdaNKUDPM4yl1
ApfzSCM+EsAQ9P838xIYnboecC9NFM7wEyu4GEKTj9DheFU2kVeT7nJaqFeA
ufEUTMQVfO8ansGmPn3k6B2WjrVeigO/+aKllPw3XjHqoTvV7NV6O//0x6JW
1qF8oFxn3KEkGpqpbUhFf4Qdq4XIk7Dxq27mQ1pX3oa7KcDRMCdMVIy/CnMq
S76VOM40TEs2A1/3xIHkLCqTDEClInGrfjXvlG2aW4UuWKaoD3SYzudkjxik
hu9yWBwt03LXFEY/y24Q+MLK9emNYNteotrh8kv/EGd3PzDCkkwbm1J3MsYI
OB/sqlqC4HjEX1m/E5HovtWG3cjY18LNdTpANdY5ph58cbQl04jR6FSBJTq0
Iizq2klphhsz8T06c7Xzr7HggaQqpBO5IJuVNHnnzQM5EeyrhMeQtK6uGOSs
hANoUYzYy/Y2oRhmk5wX+ZWnY2LkE3o5dTttOz2ud1X/+kl9hkzvftGjm4yQ
YFQKuAYmqzrolvIVdqS0RUyMihJENePhtJUYsv0maucy7hfgt5OND8X2219l
TxV3QdIk7odJq6Fg59nwNkm8slC4NTXoHTWyUNkawhGgT6BweObn+jtEGh4D
fQujwSbJtPmm4805D5IkR8qQH3MAyocC+iFrhN2b6luoK9HAIw6KqDXJGlLu
xYpYALbDZlwSOXVHzlzqG7LXXurbC9EfUxO2Xqdzec64XrYYbEaerulg6fIo
eUN9GeLhobudg5a7N3d6Ilqg075/FH2Gzx5OAacG+liLWfVtd7oDxfMyl7R0
wfy+yGf18k89M6+hrM2Hc464Djo1h0oNjlEatL8czIcd1HheTqdtqBvOzFIW
t7Zcs6YQwjt5xJoT/3llV2teQuxu3yO3agc/ODcOQSChyxTc9uD5mUkJqmBq
7kkdkmWhbQHzFkFv96Mip1DXUVoR6xwxkUciJULm0cqBJZOsajxBsAJjCXf7
9ykwrSryEgcnkQvUvpABJl7LfYaN6byoOEHh5Y3Rt9ANQaP0ZObBF4fhE8uM
wjjcw+EBpV/PKy4DZD1wZ6B1Qh9tDENKyza3aGO6It8zM4B/ZK19d6wM1eei
9k0/5Nr2gBqPSa0q6+tKtTqsFm142e862WBewjdPZH+XZO7c6SKsdrsz8OCj
zhvjhRhdzF1cqgIJ4xdbB9lAOa87JgFiX+wZXAuCP3uTrkK1Ke8m+4zUrVHt
/BrbNNlHLl8etY2nftCUg+hIzyXW29oY219OJad+fTDq0t68FZRz7sc2gXaG
jpdTrphFy+zCO3pnVyIwKVr8JxUTUhaMba0p1LbWnYzmzjDKCz+dkA1Vuqj5
qryLojD+acS7kK8xEkFt8b+zW5e6W7fhQh8jfzAgyrrwNJGUWBzA3REmt3i1
pKmLSKi70qFKiHRm28JtMGqDW5wyXY1KWZLEGt+2NswpcLIqwPdwkBaGkGtE
nFe2ZLXgkdfSwpN/FXTexR2SRD0mbSTQU0ICVApRRPkAf86hhgrotjLgqxdx
mVp+gyOLjDUQiIhsbYzXPOkW0yVeYMnene9kt9+v3eUqpF6lqPcqFCIo6TLE
tJxvM8YaibA71D8Uu8ofUqTKBNDwDHHfnEUAn4AWirxWnqAhVQUJUtKKlk5c
R2+hntGYUUuTlKSDCZP93WUpY48VaiU9AabHd/yT26Z3/erkKJSpK1KtneXv
R81jm2lX0mWiXW0iiWIDL5w9eN6HTUnG6qM6OCkZLf9e8A1bKKYYZrN1u5FR
4WuoWJUtvVEtqseKC0PSREx10h3C0zLatiVmgSrGLnUDZ+tmrg7wKmxNsqVJ
PgShraB5UNHzahf6n07ZtfnGyzMd7h9H7wdzVODJSkdbIn5dhV6JUc1RZg9d
ECqxbSH1Vxe4CqZ5CIB3XmwoNGgPdvedPRpOTkXWd1lDojbYLZeJYcuNW+UW
nefupJ3XwuDKQhf7CqMT2TXSvvBHBZVuEMoa3tXySO8YQr/PQ4uvG07GkncA
tn3bKxiKhzfacPrsAdwK5USK/cRH/SEgAIYW7n27eFraK1I+B9RlAS4nPfSM
B2Rj4uiQEeC1QB2AcPm+ovOc7hobY6QQ0nrtspxt9L3uYiLjiLkOIh4JTLTM
7tKKRJxagK+FszYXAWuyQQj//GsbKcPJTislsdXYyRvEdYq8701O//KC3DtB
+aU5WRmQFUBIc5SzyE+/KdmKguFaDTmUUqPnPtzBxhK7AH5KXNCg1C7K21YI
n9LPbJ8h1pt4FyCdNJlEzcPy9zskrnbSxUAsVGH3dF7pLkl80a/Be2TzGIt4
YKsrLpM2cG9amYcvW83uj7PG+M4kzrexE++77S77ELJxOGH28TBKx0piUzfA
rk0hALvSuPMzcJlJ7Vl72TqEbhUlgvVLjszPAMSndH6Q+uJ0rwt3skCMlyED
0Cot6ii84+7TY3Kkzb+QtB6Ra2CqPkVlJK7N6klYQt7GHdkgdfv3vkoSfEQM
XZBoPqwLrxvArbxeuf8cTh/xuNtAkcO7QZS+926QCYwP04BDynCkSaapS1q+
g8nG826RVn6+4D7rva1ychTjy6ikW/E+9WO/wNzr+w9N8qjlVjx/K4uyjBfV
FU2fobGSkcSuCfvZabGN2NhpS4xrbuT+XGPsVNaRpghKfQiaBBKZGnS4NXzm
Vcil+QU1xpd3OlY3wH0Uwn3ToxpGRW9Q7UKfBO1vuLkukQBvl9K9RZo0g3ib
iJDUgMt5io1hPg26i8z/Hu8ukH61N8MDbf2GBmcy3m9IfNHoxag66yMjWq+S
oCUl3ZHJZ0ybEK6Y5uhZvGcRYyvFwFH/hKvRoe6A4Qiio2woLallaQ5/CFuV
Z2WueZ9CJDf3jeDQszOeQv54q9+FDaPLRQm3+VbR3DW6TDNxR4rxAkeoUuN1
rEGGwExBZ2zjhPpvRza//uafApKgjqTnS9Ky71OwVZYcqn+9JlXjaNzLXIjx
pY0tu1vL0w5wZE73DCnpz5VPemRh108EMR0gvMBty/ZO8mXXfs+EssvvVh7k
k/sjl5/pFZY1MohkpvdgkaQ42KfSi5ukEPA+NEz3Nc7F2z0M99hRBfur/tez
CJU+QTtdku0Yoj25k88xA7nnAWoSbWsVj1XAAcXWh4YRkuw3WmRps+dzz6hG
CWfyGyCsHQnrVsohfH6B8ml5iYa46gMZmmJxCgRZw0gAGOEwzlQfq5uIQu5U
+u3qjgmKbIrpVnakGtJZZl8GSZHYsW7MytLtuksFWY/jg7UB+coZBHIeFQU2
a/vES2gsmrUf2cF1/cqJT5l2iA9koKWc2thQIIKWHhiR5bsPDmn4VebkFTbr
vOGLHE1xsAnt86QDCUQXuRk+U028F2svmRbXvyWpxNaoP9fL24vmW5fkPsL+
5KFRzb8OqywiK+rimNIbYt6uH+WP5LlP+bFiQcSk//wImfmN6tMB7K4diHGp
5PzWeaubqSeog3DtXE21mqYmY3sLPPJhsIhtaAmhjzTG1OWGFVkZFtwZpyQ9
k4bZumBuF5xxkslMdO9veVElBGvn/cOcx7ESKKD4ETeko5yDC1CexsxOxDaW
KwHpD54PS0DYCBhZdFtFORuykIEqbIhx7i858sYpgpuY4ge7MUe9Q2i08Fdh
xzywBz6+r1VbFI+wBsvVUY0eGmop85Zn5gW8ltL+uqfn4MIfC5Vmnop8DlvR
fQVa4mpMXBGO8Ovr0ZrxSwB+LRLTeUwxBb5a3ce+ku6cHZQTfFIkIb+Y4vwM
yY3FxJAjaDXGqh3mmHK9rc1Hh6CmfmEaNcZ9nq2efqn/fHg7yqk/+V1E+Kys
3q4+Aip6VkrTvRZaoLto/INJvvBRlha0XszuB6N7MHP2Wa+tlSQLK28tiVE+
zkRTwp87IjvUE61PCXiA81oVlDpw1JYhRAu1Vl0eVqXhY75cmj8RHURBminV
SAa99bbKnRpnog+wgojMBb8Buhk0GS2Wk/qwYXPAdQgrkQa9ToPOGBMxiMZj
516EJwREqNxVZU9H4M57MBq7TjGViI8g/Hw1J6mRPVmlGrMMLDMeV3QdE0tZ
fyyKHMG48ZgYoOAIP7ALWvXPBXWqMbmDqRz4X8imiPRQQBrICuuwmpQOizEK
8LaoglQ8RESingZJzMO6f96CQMjRU+QCF0gAwOOfL31pHb/9cJMs52d/hJrE
kTUJfPK5TlZd6AMPGzF6QkiHFtdX7nqHmFxX2Xj36n9aAW95q7eMUvktXPkJ
RWXxeB7ZNIPPgTwA+Wud1RDt0GBKsxq4Rj1RanobMFYdWr7FKwvMqZskwweI
lqn8ET3dih3hROjGJzznbm6sPdWjSLib03RupH3dwbSHh2QAttlrrn7Ri0za
fbuvimO+KYeTZ+Nf5CX2zyzvXFjo8pv2OE0l1GUTx4qg4Y5RLePRPDbEbMoS
ufOmsCRixd+9u8iiTGbyvnZcmurabWSVOX4zNLgvNzx93nL1seXEHIIpd7IR
QsZDqGbmkMQldwszhHfnrCL+Q3gwUSEu74jYTd868isfsYRa9FtgPo7DZdJM
EzdUPsMj+MZ/79EhJxq9TlQeiB0HukrzB6e1uZK3wD6MFoWsrL2M5YkL3+/P
V/UN9JxbGP4ynd/qLFIoIK40Qo3s3iz+5/4BiEahLQSeBVeIdqGZI5+TwRby
zO+tqRGgmbF3Yjr094IjrAuG/R08AGqE8lnvFwsSHfmaXaUpnzdujagKPHFK
GplAQ1dW+YGZfpbRRnTQVHFqVkO2ZuDh+m19hCIdokbQ9ZJc3H51yv0NYPav
0589P7cBrdKjD8COiKQF0OWal+m9KwFR+6GO1SKYIa3JUyiS+Xj59qDPh31g
vwQ4FXWuJ0T+vn4wJHViHbEBa21r29HkSdJ12Oy3xiMi1pi9xSWEHuxvd7sD
NsGFRHVwi44yvZBOmjxhtNK6/RxZrd2UOSggu/dn9+rR1L8NgZVZWkaRqTkf
pL/O5PHTxm6xlwf4C44dWoBaJ+aigafc4uxJmhpGPY/tHn8Zns5IS43W0ss1
rleMFuXxqwRj+tTw0rlyTN8VrCSymMCd99YKf3lSlvgax465JPiNgruQeLsM
tghQsWYx4IPwa4ykYGcoAZxGAG7eMtn7BxTWtW8i0OU6Z9NDP9a101UVUr0Y
PX7oDdkcNVAkyum3XkDeTDE76rZoPnJ99bMESMVsAquhfMduE0hQVANJu4yS
+OjdegwbwQNFlURY1KXtCQSfJB5zd09jgbl+dacnDkoTg1QiQ1Inu8/E5P0Q
GCH/MayYsbA09cD6Hfr/HTVUU8I4mXxO8U9AmK0DqPU1bEEqVKAEoI+u9mgW
bc/9C29CfMRIG+lbp/d62Se9zevPkQLvvyYZjKqII2jZeXyCJpm8HoY/Ezuq
UtbZauJlV/X4W8yVjSig/gxxRFz2g6O0vVhtQObgkwd5+QMvFhpkEPKm1QCt
IJOV3pao4539Rglh2P96CloRIconiBbqw/mnqmQE3nEK/SPoyea08ufM8gXd
eTsKoOHECg6cw3M/KSnbwij+TYtJb5xNh0K6anY4k2NlJTz40Qo7HhaWPvb2
Wyyk/Y8MLEO5NlejGfirQ6xGJO2JlhD7Dke4ZuNBbEXzrWNz73Uz4OyHnzG6
7QtAr/fdyl3/pxTTGpOet6dyjOGv5HwWAsK8m1AoOUJ0q3Ud898m1Wll5Qz3
/td9xN7BQHDVt5YVRjRyma+DYJ+a06JUwR3gwFdNiIq8PdxKhN70LPwhd3Dy
GIqphScFT/fJI+lSVKwI+GrDvM5aEEF72ycerTdLEnkK7HazJIf/FqX5jqCa
ZbqmgmSwh8qpb4xxR6BzY3I42LHK4XedEKOfTqihKYaeaYMlKRdva1zHpMXA
bOBWWVUiqkSTKyi8wdHE50W2T2hkVCzqDC0w6rO3wIQb9LeftKsDUYPVjeor
3+c8y29X82NdMs0ZvE0NptIQ84+48IcEY6JW3KvtyQw9ol7l6jMmmeJDzA6r
LHyn+UfcBPtrsSdLsWPIBvC9hvXtCzbdFEPjwiDEOGp+/UPg/PZMMnn4uBiL
B9ceHn5xIhgbdsiHNK53tA8wkFncEe3Ms94yhPqkIPoCPUHTSCfmsZsLim8n
GQ8SBYtMPileaF/stSgcHYCxSedTsgARaUUzRw5j5WKcKQObByw1q4VdnjwO
9j/AD689OlG3UZXHFhO1NmyFKxTQgjlvS0rmCFNBHptJ3k3tr1E5rv9agIL3
PfHGqYeEdbnyiobYvEbRk60KDgtqKjNMVoPLJvDixgkIprZls1TDhruNRjL7
S4h+T9qoP6ghMkGyealQ3qWHSUWMd8PLtguSzYqaUm4aUvWJF4OFvU/PwPbY
Dn8iYTgdvCwE4NVOhXLyyseWSzTORBOaJrYiRs0N4HzjSXfHb6x9wo8uJMXy
597mV+pdIEuifJ33xavpfIoF8WgXNgIHlBeUuiLuU1y595RoylxCklIChsPa
IHc8EcL8M+S4wZtdQdOZxumY7OjE0r6OKjYbtlGrtxbCNG6qQPrbnYsR4RvI
h1H6/o7jlPTFp0gMuXTGeXPfNi8gMQihqXJjXf4V/nfU7WuX9PuB9ds0tftw
Fx7v8dL91sf7KfTxlNmqruuQKrR5SkcHldGAiMRKhrUUmSo1ayaBcfniol9Q
i2k1Tro82f11S63/1cddcyyXP65NMF16F0qUPbaTy5z8CmuunuD0GYEFzjHJ
2n8uxUB+mYs1daszenzHkYiiNpWZ2Lwzc5bfQxwzTvrFHtTX4LaKqzcnLyId
BzuDwLFlpVPd907rE1V2a6dpLDN944FOgv0wv6uEppp/U33Z66IoORRdscbI
AcgABFcH+lSnWKkWlG5KSX7lzpj90gt1vDkInXyd4Xm6pBaZ2o0te/AQyzUs
CSkZClxxFIrKo8h7cLcgTrtq5rUkNx5pha6qIaVxB/HaWJsZrM7Owvxv/ekl
75SlTOIGsmyXIU3zBPMfaY3zPkSVsRSsqHmhPpDWAcL2LFL4A3ZOrVlY8GLg
fBttywHnsubNSv9tl9Zqe77dKEZo4YLUEYEA4xE5ZESbWxju+94EtWnmc+Uk
drfbuGLhI8zk6XvcfZ2KsYYAgNH761IYamii/gkSEB4ywZbxDZdfmwYowcoY
0EzISmgBcMRFms/cCxitEg+AwnY/aP7hXcpWJJUOLVLD28Dks1X9V5POWZuV
xFMXucVILMjDt65qSHKsVkUtPczczB2B++VGHQdPPtgW9EpYBiEHT+8R7KLM
3tWsc9AUkbGeEmX9Hlznzi+lgWnl3HG1IcKNNA453bILAvn8M4UEgBbXT7FL
+CRfM9F1Wn3Getfp709hV5qbuODXoJPTdtAyzvA4x0V+m4rzfhsk00q9SB72
mSP0V/ERjtaqQG0T+EAl4vuC6MDx7zY8LXlE8+3hJ8oU1jgVGqxm380z39im
NSoOVTNnQw3p0GPtbZZz9sPfzz1QtooeYn78+PvYj7+30RuMEyqTHJbLJdhs
NLJtF949aIRySC0qGecyfM/vN8y/MgyZ6fhqnhkLC8TA1eNTw3xRoLm4ooa1
kJYkMEh+SrhBFWiLwesMtq5JHOK2CDLbPfr4nkRpDuuhOVXhbyrUnDmL4W89
AjacDgmsyS+srG0XbAOGn5oum1oKzPfwGa4xLIzduMDLRs+axt2o6cWu2DiQ
HOwx6HMlQfIQi9oKobF5jNQA6nXIcX1WXwnpETaeNV+hv1gun25XxKt23JqF
FG7cMpCKq+nqHcfA2FkGaxm5C9MMFhIzheMmu5JPVikLUvMphzR8UphWe3Gn
/KVWHlfTCRhIfj1I8T+ig4Rp6+1NlVC9kJzsJRVCNkq+/Aj0sEvMSDlgSRCH
wE4NuKBU4lbTjQMLP3xgIviv4AfwHosbrHIKjHcpAdZKx7KTo0cJPFRRy1kT
XOqrY7JJhsH76THhaLMPdljrFgV1t0OQkddyVuZQ2BWfPCuuB66shdQdlqOd
GYzbhLrE4nmKlSdgWXTlrulfwWi7ZudNVeyieZCP5GLEl+irjGPcEXCnZd0M
bvE0Bf+uhnXf4xAfR1Z9pPQtC5ARGjtSl0uxvLqUWf+LoStTTOu+JmMpph3J
B/sJA+Gy3tj3rMsv8SDEyE/GasRM9Oe8MAv+HdfijCYr6DUwXAyAjRNyqUN0
e4H/ElEJBUX4OLWFj2Fx3VoWa6OYWN8id06ZQc+/Jp8X4+ChjS3PN6PB5vAT
7905FpolKUCAQDkDdzJXhs7My98aYq3Ab82ttkEN9gnYFU18yzaDI5BlCEgP
gAvzh4UYDPTVSnLrtm2cO9rU50FmNWVub1SgGmF8j1K6fgruCnmIs7TWbjJv
YoY7UlvmlCPgiG7DVb+ZNbC9QG71umZug01bAbPpfgX3eGdK70WKdNM3YkZe
y650/vf56lZInUQBZHgzZ+dmfU9XWU1MNlba8Dvy/uegKrEzNJtCX0ib408H
XzaiOX5uXxSXRps7cQQwBQaub+2wJ21JIg5GdmtsGxp/M8nRn/SJvz3bGHfg
NyNZWoZ5j3n1B4BS9yTPeTSesTtQeLLHzpP1EecjfkrhiIsV2/d7dwMDN1OX
ykn7IOIKJoW79C6x0bohIdskHuK4ZeVNVBH6CuyXzKN+n34CTuciReXSB3aG
SdY4xvj4QH9VqXFYvfh1fNU9CrPFboUvRuWc9bnUqvS1KKeRIXlATgYWNWGa
k8kJP9cpWTSgeHsDEA3ShHUfhvZGNtOqG0jZp/NpGCjppkHRYJtyJyR/W+/o
2mr9VxBX/DYIlQI9Zc77BLSbZhkfAuPjqkDKTDjQ9lXfcYvMjpmAgdMjeS1A
HFma+7sfMIXeM+XRwpsn1pkWA/CxU2TUGqyjmlhm94AOUHDYxfMHp0xCK1qk
fJ02ESPxKK2dxJCt8q6uPHHzt/KH6TBnOO762sZfUE+5jZNK9G0lcTl6qHrM
iCgdIGUQ79Hz3q16Njveh+ExpxYV+rlWAaaA1h/q23cVSNLYIDAe2ihAWaMd
5lfjWp7+zQd7n3IBhk5W/pxRanBMIiURZz3038m+IuAJO/qDPBltE0q1BzlC
hTyNlejfTX9o0rDFMn0XCbWJN6Ld2lupQcH7hM9pZDHaEQBALAS/8uDfqiPR
y2W8YYC4ai9RSWCRs9P5S+WXbGDCknQyxmCqIgKfYBhlvTg6rdlKIhC+2ZNZ
Lv4j6Mi+DrByND1iLkAxp92agEyAdr/FvhNGbRWfLfsBdecYNdr4bisDcvqc
lwvGQQedBdlSeCjkt9rkOBzXHSN0zErBNDjRkzEO3QYdRzJtXqiOB7fRhBsz
954j5vB9wDwf52519hjzE5NuBZ5KXvnmrx/mqx/gbrjw3GcKARI3RrM7I1JN
MQYcDXSIfVDXRxZWLG4FU0p2NrK+rQY5NgWcEqh372yY8Z0kNuuGLQd63vwf
1jiIQ8XB0EbrvUoY74We1I3t9U37xZNnKVdkJWsCV/vMAp+USSqzpFcklBcG
STePNE13f3vMFHY3s44w1pcEKPtmPMzKSrkqYUUnFPWDFOH7r82QJkbfR5a+
gWIl7kj3QMIVaoDGOcEexX/JbbqCmcvBj5+gjVkFBZzLOW6meE+F8RVFYxvT
ogT6WMPDD+2AqPEf3SArBTSDYukyoLHspFz+AR96OVlOX4EjZu/uHqwctkT/
PNKZxeahyy99mXxUPSho3UoRXmS69CWyt2Ld857VzkXpN46mRGRO9W3Xu/pV
2R7Nr3GPM4AwCaumXNUo7+ZeMM3Qk7ou0O37F2wROqGGX2UKsxavVXu6dS5n
GvFScYUJJusNk/d7ldemnGffRRRiGBzVfm+fslji/HEj4zpjRR0CNsPKhFtU
NEhoWwHJ0EwbjDVqXOGx3ZdwAoEaAb7jjihO73cleh8p7ZsanIZrthjfXOYm
ZIfZlHGK0O3krbnnahpzDI0OZ9Xjrvt4N1+bG/skmzgDxXKMAYJdxmc1oio0
7czK5pnnXAO52Gdu+ZGY9p8b/3kHVN/8beqIsIxuVDL/jfaJRiTLfYjhEm+A
Y+80TUKlAD8H5df1vZ2ujxguLl7VTMWhXtzoFzkS2i/ohVDWR2F+p5NfnU8Z
ciyGsUQwDWJ3XeyNgUHtSoL+9vOzTnycKntj6RWX8HtyCtGm4ed03g53hKpf
g4qCjD+SN8XpdgFSM8DGmZ7RGLHB3R3K5agPu4WQfeU0a7+PuicyjLFpKW4N
vfNnf8mES5iQMrRPqy+2+ne7nq0kjByEkatJCdrJnVgs5soKChASzVYYHNbR
/Hj8lZ7nB1dEZDX1uWuOyG6dti8/ymfH15Wv6mz6UUzWH0bLZl4ZFKJbp0S3
sdHc+RJtNvTjoTvW/Q9GEs+CKawRiAigC0SJMrQcl2mswgPioaUr+lnSxNjC
9WSyHkbGNqQ59f6WSil43wCcaBBJcKn38GrwPFFC+i3R3Mkn22jyv/2w9YjP
ySG/xFDkdalPJv3/wglX64auKTTF6InTD0TZhJxCGGmUW3jV0PSF3C6jhSS2
1MJ8RAMpTm7X8reuzPFecV+Jc3oh57vfPcSfw8QWo/XruQSQ2DmSRIoU+LIK
1Ix3jsRkhMT3gWCpONuzXIshKgKqXmXYPYB8xzG0Rs1lrR0A/hyJKYiu5hJw
hVzfYsZWQ7AqTAeFjKcZWU7l3DYEEJbaFLs8iMK4MgBB4sX2guUleOOERjjJ
RSUlEadN5JvSLyRrUF0q2spOyFTqOk786yYuVvhPGryMwwF4HNGhozEkQxup
gRBQjjmDgGlWwoq/Vb7ZjmbNsfKRfHwivfbhuiYaawbZ+hj5brlBpaGax4YQ
S79G0lWB0JXjOKrfKvicZIshszyEPTG0TLe+oS3iKda42INBXDdGf51XSgfi
A07BwCaY1iXH0wF7Sbj3Vw06nGNIsT9lSzpjNKIK4UY7bqCSCz2oDx+bi1Vl
MobahxU0w6hPV3ao2xj/Wnpi+K+7R1/EE+ELBG/D7pS3hGYtmU8jWFaFp907
muE7mJ63lTLvl99PCp6PTj6NbiFyajwwQGuB33kkmQGDSk1q4UI5DaBu2GdV
d5QlJzCTMUvL+vlZ7MTRyCjhZ/ZirJWZFo3Ifl8yAnBZeQKRu0frplONcvra
F+lvDxCzWP23VTIPg6dke4k2t5uzf/SxyCkCmvusJiOeZZ2UA0w4eUREP9n5
rHxySU2QgmGFwqCI2DxIPWU/Eq4egukMh50Qq2egYeCo35ByYX/TU0HxihYe
s/4ksJcYKX5m2oQY4ca7B4WNqNLh9uT/LDqyBYicBKutQ+XeWiBPST3IOkqK
fLwzzWu/IKmNuxPidQyZliic9hm4whFoAgHq/92iefCWVApmz0y3JS0UO8x1
1xsc6u5s1XvxpoprMLZTaaraaJPkHXEQxVEG6fQrvNGXSNwLN9JV/FGm/RET
jRtMCbGbkSIRbSKOoDuPnECelIOoXhWkCYgQFw48Nj6n54VF4VweCJrBYx3G
+R1+jKfqCHGkiMsRX0Lnwc5GofSybRgmGhOwOJPhB/O4GVmUvF+l8ZhkkBLX
LZcUVgx2qObv14IuAD9N1zrDrXMUljLJNGDOcHe4PVh9H/phKgcwOc0NbRf7
9IRfg7eqK4+FIf9X3/hrZ8IjkG4Hej0uwmTYTdiDP7dttxDPmpJzx4HEB3nl
z8ISeVd6H++89cCd3PN3FSNv0vTR6YCFxsLN2yBb2vo3zGblmt6jgdSF3jN8
r+/IztqkJ8qIuHJRXoQJTpofIayKu1XGBYrU8Sh8ny3VyAmga2M8wtSV8EwC
xRHrD2+pMjjNbmwTYSyVSLlQVI6XQQmNKyjnVJJ/h89kjW/7q8pQW/ijzBu1
W61aLjN4GF4RjgBVlIsMwjMYsVOOMyBbPAR+gWz9mYBoXFGK70pD5HktTF7G
T7ooFely0FGCk7zfYBDV0bSPNDSH6MVQACdN54WpEDc68uelx+2nysEJQxrm
/QI9BeuJX+7P3RhlxQYZybknXQhbroDcZXYVOzRioV94Bhb6veYwLMWCef9/
YZvJJeezjVJIqiWkHhI9a/MZSxqAxKX4Saa4HxJbVj7nNYVxhWy14d+q1oJ1
bBqjrSg/VXMoN9BckTW4tqx6a/7F1sH/nIT6mi2nAHfc0gTh9Hgd6agm1H8w
OUnV/DeSDXL20RQtXS3x3X3mW4UvAEQODGU5NTntzOW70dCZ12pT1+PHEVia
ftPO/upSZ0RCwYUs/fYt2k7oYo6ceDBFWFyIBmLku30H96yHJMO7ck9Qfqja
D9XvnJ6LlvInoq/7SQRgAt/DxEYpIQznsN52AWy4xAN/Ep/SnpT2CEPaevLU
ZwuCSo1EnJ2Y1Mc5FVvd2KBUcLDu4ChgRgd9Qs0TFgIrtBuxfTnZTzPDP1su
Fzf3a0ILx6s0xG4skNLrvLbjV/hF2XypfKyCY5zORZbTftNFEOhgzYj0Zeg1
xYw12MYsqYWhCpM1E8XBnx/t7FN+pRaej0HrAc4/eGXzlG9/mSTksYj8lS3o
uW0KHal/yUU/nkj/OBH2i85Qd4tPVYEe6YsmfDSZ/rwOul2HWBDAcVKutSlK
LIVUkWNSRHbGpHfUgFOHBxmLRbyOAEiP77Oa5M0yhuce6ixRGSkaHiQnB9MI
fLxPTUS/UEcIg+FzJL+DItuwC3OxbJFriFgYZJgAfZo9r8xuYHwYaVfPEjuM
K2AvKLqImcQWRNL2P41N0K1gJanDwqYveEhu+EswmFLP4S8KRDhRnbm7aDMS
ZJyDYoxB2gVpEGyvyZIUTnKWyLWBI8k6f7bfu7shO8NcpFJhqcsvUu14EeQZ
/Zmchl/Ie54iy4an5MOWOqBSPnz3S8owaX4AAZ5PuW+WEihYHeDNRsVVqW8J
ohioC+cdnS2oLrOq6DFRC/F0aO1eiUSQgSz9bl1SqNIlXeK9JeEjaww8DPxJ
MfKBV1a3W315wh0DOnPNpC5cBNXVTda4JTvEU89ZgIdsqVXTmmvuXKyDjTx5
JFCIt8LISkjMb71cVCvTB0VMhHKaoJ1dW4kVMhJSsD6x2XxT5+8NNMiSmPcd
vMAqo62knleBRhtyFPXS4iZ3AmBEfGcML8IkIyihMnYgKUl3wUvRZpgb30uA
3Iam1YhLXzoR3o1RVA4GSsuv/4nk0uWUsMMG7TvHae3oF8qpDxrkgxqvvetW
bMp9n+05eALOMCF+kTHKq7T583DCsaus7X70XegdL5/I6Zacknm/amcsERFJ
kZgWZJSAUGHK2unJeJ7tESd+fBBewg7nESRp8LYWJWEeVlyb8HqAN7XToN/f
KTbVsj1FSQA2tgYpwXdtDhghMH6KP1rukL0qNxL82RE3dN1o4lCnuido2/5C
XMo8zw0YcVTdImUFrCiHVcOe79MgN7i8CGBbpjjQE38+dYBrcIFeR3Y9xbR8
X8Dx3MYgOyVAz8z0Mw1F8g31HEqkZahm88TuwRP6nyeFkVyUtp1Xrfm0Mbcy
H5hQ79BO45BEt4k9l+14uXIcbrYNeNwBhdGJVAyl89o+VWh22YLHArWd7vl1
OiOy+PZTxgzfiAt8tagEdWPaSOYTO7GP9YlkW/12uAZRGWyBCeWWH4HLwBJV
K1a89RcRNHM6Cp2KBwm5lXQl4KoyEbOjqAIIN5xPP0i7fHRsVYx+p/lj6NGE
zQ4natEWxl4u59ISEmBL1ebIEGzEeR5bkigZ+lYPqZVo8Az7Fr+jpaGfNkTZ
ElAlQtc5Sot0skq9Y/9LdQ7Dv4TmTquPdjT8nguZ/+kq+WHJGK1ppxNKfFe+
Czse2IkFBuadHtcbbh4KlYYj01IS/xt8B/bywNlMO3zxmLfI/e2ixuZUGT9M
PgCy/dyjR+jE6yboApVIMiYYI5uqQHz73eqqWvCNnAmhJuPH1gmfhBIcUgPI
vZSHkkrFcEKYBFCXGeRX/7fIQ9MrORg4WOPtdsPB+KoP+lArxwfK13F3uIZZ
mEXymtiplYel0ckS3Qq0Ir6al73+F2gDTEd1xiBms6G56L/VBz+5ena9cNQo
9zpkkmycIHep2AAqwxK/HnRd5FYtMTlA87Adbz10BP/nWcGlgw7Z3nzEyd8Z
ta0r/MqUOC0Iv7KVrlQ5c3I2PFW/OSNaVNLoW7wpvTTn/oTH8BUbC2vB3Qip
sVWeQ83XJPNh84CBV98J4V20wC1Wq6CI08R1uWuaGolMlxP3PP12kdqmNaa+
p1K3MaFPxiWOGXg8s8MyCY7d517CIn7fbdI+43qohz+sTbSoOnAdSwNR7a7f
SjafVnY6J1xK2cJ1+cvXTUJiz7762eBn4Narq/qZLBSG0VYQxd96KjA3DYRA
IrbNNfaxivZw9iwvF65CIZVJfzSOTCzrUYeRcwjibfmoOhHcM+3bKPaYoKgt
2UueDQvZkr+ATUYwXUkHjY18Kl1oMZecV0C22+CIFFBll9QcK1OTyAB/ESC+
qAPnK9xyMgIKIQoh69ZYox2z0cCELQEynUU8DJfNNnhpzHhqWRnmgaS8kYNg
UBljmjj2VSH/jHuGhoKpGRByYjqWQV9Q4bVHUnyFDn+2pW+5BVfwIRW03nS7
9O9u1QYOy/AiXiCzM8civ6vg4/hd5yKY7vLTdSOF55pvD2x9wyAP4mnQ6fWw
DAwd+9hq9Qkk4lqmUmu8wOND3Ode3WWDw666F4LlJKPij6wIYbRXDjbUNv83
EEYW/DPqcXl5ZcNVqKQpdzC3MIsI6RpxfZ4Yj6L4F1+xW69149w5e13P+7n5
SrTunHcyyB6cMIYHElP5yZkZbiGDVtSD8ZBU5e/uAJzX1vIjFv2s6DBpQfDK
K6xrwY8WVZYyjRjPboAOSTSCWGqR0a2+9n8BiCYAmnDUJ/IeYNgr7w/MWSPK
98D7Fmn7r9WNK5UqfP1vbpkvGqczbBHXZODijYMs3EJsb8DlaQklj1L+nFz3
xzuR7qOzRB01uF8CLyMj3vBxz2qadreqTSWTajVwXX3pvxXWkpPdFpjpnrmB
pKTWLjrfidp9TNLMGRuS5YcCEO3xrQYfMUxFxKtC4FQclyH+cHIZO/9wKvgX
6uZUu5UARuIbc9MaeF6kLw47zpss36JNF2tW20TYahjEda289ZjpOo7hO3Cb
1NTbVl2nKwRcTxEauZ6r1O79VORJE3XYUwptZk2QB3NHliungfoEGpq/uvGG
5uACeMl5ggtR1SfJhDDvvwmXkK5jsFGwTRqVNS1gWl+grlqgtMK7CgctM3ov
zYNVpiA867BUKMAY59h1E4kLfrfE/sQV9qWGSEYwGeW5VTrtjeefQ547m7i5
I/jvDbruUqdQtsHzyGf0xpRfZZubuuWsuVf8/JyIfgv40I4rx+vaWUfIUz6I
co/d4cJHBP1qqiV3+soZGrpPTGc3PxCIhv/FlUffK4cjIGv3PwThgbninM3/
R+lmEfRr2zaRU/iTZALiQAuu9Qk2xM98v9CljxgITG2GftktWPebmsUBzlD0
ViQScTEqf5/0XziCYuyVUw2HGTrQnh+e7wN2Do5JbIQZJd2xzgHSlXCAH/2+
3snvv9ctOt7vGO/FvCYoSP5OurxgITC4OaVUWRk3K4K4n1MGUvbfqxPNsdfE
NClSstqf2OTAx9cGCsRvRyLC0Os3kwQp1UqH4JO9KuiOGEFfWVARoHs79yIS
jhc/zr/M9fBYAbW/jTMyz6aG9bWO5XFTXLnY6tZ6m4AlU10ZqX/fNAuZIcNI
hmhmdbuDtfB9dU2ApyBNHG4Jcs6IcwvjYMW60LHHh5D0kukr6NTOO6kCGgZc
lBOT0TJ5Rxuf0uToTuGSeIKIs8Ro7LyCTXFhDjLoTn1WbWmvZPp8c2xbCPj8
DCow3OOpbwiqRfPtDGejVfEVum9YJB9JHqHlhEsDvaSZ8tDVtmOtbjBiKLA+
i441+BKwP77vNd9wFOYNUCfGgm7f4U/KoxYt+hd2n1COA+k63N2/dbhl3KcJ
PlP5p/266od4WxVvkCWY3Bo4ehwXWCO1rwgCWMwj3wwtwwq85Eb+eCQFWlZh
RMobtUykcQAjEyd2V2g2jjPUaccAxtS38Cl+J3RdhF4bIkQXsnan5vjcaq+t
1j5PFmGKN1hQ7HwZL4TB8IAVoH8L0pu3r5u3XKnCF0RFTraAWWDKRQArF2lO
oKExUWm0vGJTF74seGiOZURNbo4UD2qcaperjXlEQkWbXEt4JyxusmfEDMTJ
EnkufdxQetDyuxGyENIZ19YYH/tgqqBUc/G7/46ZkYfF9ZPasM+Qi0DszREs
07hDEAyZXoHk+i+AwTVVrs1AOWKFUxDFZ0b7Qo+aj+/NQ8aNyxzz5gJHzEoG
5idrmgiXDjw4dhxvWQ7AKIo4nyer9Pz7r905MoFxZ2AgP8KnBqADkE5bmr2O
j71u+RvLcNKabNTFWq+Xi/Vkj068Z9DSqCYBEN4Yo/pBnUc8m3nIYZd3KthD
7QMz0KeOkdA0KtV5H+K5e9WcH1DhKJYJmc21/VrdqTm4d7CyiBIWNvOCfNLP
nr1uKlc2ViXfeppgE/9xybFRDo2EvFuSrqEBhI2KIFRpyDvSpB8rA84w2pj8
kiaF5FYVaXzj5lXEewzpN0zI6LFjTBqoQbOhabxUSF70LabAbYDaMDCuCePw
cT9aTGtrGS7KhVv+U3POM7jwzCXGz8GdBIhc5lObywzpExitb8fN2u8/WE/Y
W77sS8xEUjWMj25zBrozXQHQbQH7EQWuZ3TQ/myC83CWcCI/UPu1CVOyRewa
qpdLOguVzY7skQRi5zFYOQFg277OS1RzBocNOfoxlYKYypum7hgQ/40ygXP3
0s31c2FTdz+G9VpU2d1Q7FipUHm9bGhtvogoftMd4ugSOe7opjo0hGsgTgrV
8nu4XqQrITKzA1XcLkkdmOW67f4uussgX9Jlaxh2zXvR+OKyyaEAeTSxly7f
2ga8nauktlAh6q3x9aU0jbB2H8+1ZFLZFSqMr+/lzC297eFj87U2/YKVu1+2
gnJkcikL3KFjvkRghNtFkwsLaP5ZSkv82HSHeNhvkYvM5ZibdoPBUSPn5lYn
atys4IHnkizruOCPJz5Q62r/iviK6DZmyzYMfBlI12tKkBXnku9apdkKApFr
ZjjdKHbG+VogZZ3pYYMoJOt6FtQwB2pv/UeC/ckTDv2ZFuOQyC7LaAGuUNks
QlVC5M0V6FgdOIa6fwurx3g3msfrIxqL+4zlxVe0xtvUt0J2NFBezlgp0AZK
KqL5s8zjacM2afm5CGwJCM4r3Lo3Av1xcfIYBr+/bHq4dJEcifi3i+mdcstk
keEd9WjsMZy+UzvPrI5ldDuRRSGHitKizwgeBsX5WWaAmkfWlgKWP9LmPD5w
VmsCRmGc3ApxdkLbE1KTq/Rmj5EycPmnjkc0OMp2Tbe8k3iErKU2GdfwYEWI
NCB63VqHACQpuPmpTWSns2JQZ1egCifBsGbKkA36ZI2VPqSB+ANoYO2AQStJ
HVp9IEorybE+Ow+HxhyoZfdatSS9k0j7+L7oGqbG0Tk1oJLruORfXH6+JnU6
YGZJ7qSqmAi4dWRxvreOSMp096//Np1GctIaJhM/5m/kQ6fJtk4zKId4AACf
9/PKV+VrzzG1MZULwDSyQLZALZyZPAJjoYDxAfuAPqZqwYX8051+CjIM29x+
I8FsGHWPG9ReC/qyTg3cyj81AWKNLJ/L0jUrjhbbEoSJuGtue62e9Llny/zd
LqXQdlChKZuaB7WvbTQREWu69FuRzzGBcOkF/5wPgKhVoAUzi/iDtIS4FRHF
OK33U1XM2L7ujP39EEHRfhq9q1gd3iOgy1C4+onnmoQzhgbv5Lxy0E/3knEl
P9/7GQGoBiEqv5hDc5sJnT+7To+3A4LuLy7ixqh0fJSbiKhmq6sIp/BngW0g
n1eWEYLSslGv2z/arzkVuNnXuR8DjBltjCiF7sAjntrPIDVbJ8FkiydkdpAw
IUBIdt+0/LnXU30W04zLbtnTShFwqzHI4OH0X/I3C/U2MAUC3F9og20eVM31
cd6m+RH9TAre65bSBx5eZFRS/hqjpbds8sVX79U9ZhVFI8VVnyhytVLBGdAV
9YIMzBLQsEQ9uC7fnqbeUafmvEdvEMTs6m8n0trK2s+WRWG5XQ5CINgREXfj
lqcKXLSdBEYXXIngv7RLdf6ngiKHEUZZES6b+6pMS3Vhvg3KQprqdU+4hZdx
+VrW6WvMs9fejR/WNzeud8oAJTohsGV+wgzXGZhunbQFJQt04yKt2aJF/tfO
q90IcDnNzunLjhMMcuBsZrY2DZxvVM56r/8dxAP3v21rIRgEEyg/rSpDkmr0
TSD7E5W10jh5QzG3tbYYxmE1mqXGnkq3xOdTc/uG+8/AlzF5bdp0s3KdA4zO
QSJIXZ7Xw3JDlVzebTSAjiRXWckosHrX1ulDVQClAoTp4/gwn2uQpFzI8Gzh
VMfJTVTlF2Kz4VW6huV4dPm/XUG1YV19t7f5FNruofI/tsfG6FDxUxxkij8Q
Qn/ba67fUp9G085MtCBGzMgO/E1yM0ZfKxmUVbPzqZtzuHh0IPfSaxGaPFnh
7Llip7j88l54EGWeAdh4y5KInx++uRfz1bXauEXsi6HkSlSXbwg0TBBtGjnh
sTTD3nsSqShr2ZUWAw509KAKQuldLrblpNdV7dtvjADKh+HXkDgN0g6Kwweb
XbFX9PV5NGSyI7M0XcyJzAJ1Kx+CWnCFWVS3O1C6Hgmra7m6OXx0IMdZ5KK5
A3M/dzw6Psw1NbRCNnyRaAmeP6cTaQjPehy2DU/3MNk12H73Esjzcmjwa9DK
GmEtnw1PUJq4RNFxoTKtsjwFDYfHAgHyEVkyjAz+IgdZIIxO6kSXVa6m9wo0
MGmPwofyU1tw3qqstquAqZMHWZKsJcZW3Ofa1RYC7sEnBXBK2+0J7ImujNYh
ob/IGoYB8o4DuZMm04PtjX2mePDYeo+1bFwOBbmGaLL9QTqgyEEeCr/eFJan
nHV0HC7AsNg0/VpG7KtlvDFUBugvHMMZNL+Cd4UCyUEbf6h8DaSxliuUiYap
VEqb/6sZ+z9N66frMbk7/fxZNgN/M8/8pRF4txdb9OYm+JWm2y1qgK7uHzL9
flRx8OtyItEWYkI+8FvIg2aVzHwYFBozJVan0UdcYuHfNWJWVMcMwHphsdxE
0fxmfJrKlWp6XGQKpVO1UPIi87EvoqUDsep+1bw06OMrdBlLuKAPTN//0TGF
fvCPNQRpR9sP/SYjwmiVBgxtyxM8fJ5l3WoY8MPOD8NJhgXyk3yr0MMzCNsy
IHR+nHmtdvt1EvdTbY3c54okbIxcKh5nku/agyg3yFAcfEJ7iAF+XnYEPdH9
/+pmfXjD7MnMhctpWzZfXa1OyR9cgfWjCc1+IirgrfZpj7BrQGUwk6LEQlvH
FpgI+v8AsLwun/Uu+/IXknK1TnY68uxNeArbdFsuXOfQjXyjtN8yTUFDw09E
PpWJoQqR93av73GoPaImstJ6C441qM1sjfLdk9iHTycT9ljLh3lltEs0n3Zb
DhZvpooRjrw6p3Y86DVGKN9RZzkPZsVFg8iSfezjB4iihXF747UThQiOiZYd
9BUqmPxw6Vy5roBBzpNI1pHxPMHvpmNB50P+y18JnOVf2M/3v5IJkZ7OXLNw
hKA9R7N4UhziGwKKsh1wB9GTt5CrBl5/ZvoxsavSsOqE9XziQTTR4lYKWiHk
h6TFCGPtNSUEGfZlwrF5NFATGKY5Vlt0yaL8tYLHYGkYH5PsDYAXS2Ahbkkq
VGrFnKqF+F2lqCMU/vumjhWIrs6rsClNFXtsQ6RUVnawoFcZZAliGPNQvlt2
PeyZJ0YtLYOpaGKxAllAe95fm4AcCdIZ9t09CxyDzfVBM7LadSNL7+8nhQf7
vNyQH7Yarl8Mb1OSrZ4+v067LxRgdy7PEqXFgcdu0Uo+qw63o234RQ8vVuXb
0V2RBHe1nneqXvW1w4KCprVgr4mrQXpAKNSY3WanTkBIAOxJ8mkIC/iKU7hs
4qHFQzzgS2ZlDXGqVeXBKJJda3xZbSsWARNxDzTsHQkrEyHdNqLKTsFtHAD0
6PutQtdV7hyGtUvGZ0N9BhenLpymOX/ZsuflLuC0kxqfuX76vU9qR6xSiOf4
lBVUxQI3lBqyVl61NDAI8Nj6d7RbHPVCjl+SRI6XZwl2cUDKPDotOt+OhWlo
cfWfzxCmBIcZM4EP7Oc3bgQEPl38AQwO194MUk/4HxSgULObd3uUZOtM3pC2
3LPeprtXuBAjilXQm/wKe5QdmhkRAE07QsXOmgPZapQ78ioGf/0q9wFcd4j1
nEJZCpZAE/dvg2XnTYZ3n9QUeFkOO64IKRqFxKJDZEm1aN+xXHkhC00cLUKV
eltJwLdyQFbV/g+Rq8PBSw0LWssEZeT6D0DjE63N1SWFmxr37enNDLO5PX1c
ZBRP3ahyUoWc6PTAafy+NTBS8Z+BLK9s2xY8uh4ev5HzU+Ek8VxE+vRtkZst
sI7mdrI7BPjzUE1cusnNVpKjRvjjlKH3vH2c5TdOc6SbYilCax2Ih5Jmi4GV
+hsJF8Fr0r+nQkBd9AIOLAeLbVxY+bz22vYfJ1bIYu/BC1yxocdy2rj4tBNk
IBOuuS2QVM+ItIG7FhE8ydAn8fvtbJ9Z75+ltKIzt5yLFtPZ4vfqujWcAmDL
+P+hzNG0XkIySLYl3lXE6vopQW0ntMMP3QWyudAVY3ZMr+KhiHcuV0Go9cx2
TEjxz4nsDBl9YcWmtNmpTzd3XbIcJ9hELoYRQLX8IKVOelWPixHsSi4QoF5w
U1SCdLoVKKniDuGVei89qPSnaw68q09JgMbbyFnDewPy0zoMTxcOglA/fDRK
Rzq5A8wgG1++JqN4Pi+PpYRvdnHEdcPZK/L+ZgnCQnKPNkbwDxAWPLl+wvOy
h1tNlV2pExmz+8JSdxxb+D3Qu7nevx6XLg5jMuFnnt3Gnh4Wrd6n824xpUXy
xrNmKDhMl286/mODvQukLKlH4M/ahrAeXN/jbDYMptCXXtP/RgMaVCHisl/e
x2jmKSZWFIVJfgi6ltKP/Xj2RomqtLG3txUmWxy8Slxl5T/8LNHV/7X7Mpjh
21p4V7G8bTTnXvQYPJSUqfh72fIhGhrJjy9zyohPfiqDTbvH/ysy/5NdC6Kf
cvraNt4ZZrKOwievR3Ng8cXc9yRgn/ShiCZIGSP31h2/bvLKzSRtHkT1aLrI
7Io0eDZ4TPGbru5emeL6b3xIXcScCjCPlhWBOVK4Yi8CKGVPvUFudPtoILPH
BEgUF9QepMb53q8O9/SXAaBriGwiVqXG+UY3m2JEHRlTgXV6phAEZaNZg1xv
WLmBanI1SGX4vglYnA52YY7/D2vWHU2hBdvcU3i/ACer5rTp5v+DDk13zrmT
BDW2npsAcnWaS8H5LLUvnE3bTB4wSrtZrVo+W1AhokFAyG4xqE4aCt/VwWw8
LKmE4xBIo350vMP3km/UnBVV9qb+6c+beby1AjhARRZCqEhhtkQHAl6lPsfp
52cK9g6mcS/5a1FpmqMiKMBnkV/AUo9Y/7J1k6TgN90B4THMi+RRzXKVQuhm
1vUU6azGkcYteqRGXu3MHMclk5bO85rAPQ4TnpODlF6UmFK0M9zg4MKme+6A
buhblLO7lJ4dOUrhIFn2zQ4w/gmwyXrOqD2nIw1RA2L1I9AdyHzblLKjEHnv
Fbm3Q5nlLBzTY9xruC1BxZDwNx0CBv1Xq8VsoWHnrvg0vPAvgcGk879Srmpm
nD/LBuzYEcZCymMNeKAODdUQTLMrnVXsWieRIvu4Jw/5lunae9QaNLkO6dRL
vDj5DYb/HNfUU88ZYwgLWaTpiyo9oOi1zcDwutEp7zcg7g9pVftodm/y6wo2
LVQtzH7x54uQn6SkmkIatiw9Y9Ua6e32mCAADdh85GU8PzPwjTmd3IgwqvR4
Agy4rSpDTnMaE7MJNH8AnKJGMdE/BmZXXUIqKK6miIuhyXeefg31Kzr7+I63
ZlZpK0D717Z/Vo065PycCQPRYtTR/u7js7lA/RKm+sOY1FyHtwabRE7WALKM
J80GVfrQT2qyG9/Jbfs0RbcAE+fNbl1h1q5sQLTBsr0yp5hBv8Re8t9RpeOk
OuTOwQR6CluAmDzmt9jnX3uaFkavveTm99Hqjm2sAGd+KXvqIJJT49FExg1a
NZAdshg4LcVUfG96UpeAIpQX3WOvT49r9uOr/10KuC0VZnUDPOJTwZAXDPCD
C2E7VRAACmbPXokOXNYRNZCRiU0ax1CcFxbsVxpam5g330R3tgQeRPbVCXWC
ZqKYpglou8pNiPbS1Jy5hU8QIDJFhwDJR68xy+itsa+B5vscl9xleG39QlcH
m7u3kSyFCO6k5/qwfLoNm2ZJOIO0XZ1i2L8eerg9YxEsBYUiDrxndDbKIcOF
Aujm5cDZ0IgcWH3EMXrH5MpAxDYuVdls8XML/I8qLGj9hV3zXru4//c3+yDc
FfMIZOsfMUpQtLxb60Anr+ecnTbdh9EqIpGcQostIdj/HtChbQ3O9ZJKz76l
xins5RxLycmBE5YVF5YoH3hq65mssgzUg6vrVSx4PEX2grbSIJB1xf81RdOY
FV5csd/+ZWRbdV3wzesdPSW4G9d4QlTPogFxY8677vh9icKtFRZp06jFAvf6
YooWbup6EVFi/I/9s0Ko4ZQz/LkVym83+MWVVQD49bLnPf4SH9sqDqFmT7Pm
Qm6zLCJ8WhqC5E6lxYRWg34uTGSboDUcxH2R/mWW4JSKpYkcwYGgIm/ZeFhh
AsrBgAzeQP1MM9d0poVMwogDXeFr/iPdeXn4wWqjZBGR8xkVogQuQ3kXSLef
1BIWSno2FV6VQaCFy+cRO5B0ktD1faZp1W+GCmOYQ2StgIZortG8NfIE7pDd
rEjmaqDLjlXy6LxXCaLKRC+WCCR5vVMjDKeSYaPAUpmV47/STCBDToIrdm0T
kSiwX25V4NpH5iaaMMnVdc+nEyNQ2syRWpNdC6xDqq5Om6SwCM9Jqoulmt5M
oyQBCCOg9vZtXLKn7pOPMvE4D84peCHtE8nRodoe+ikU/ITM1ewcD2TnkSgx
deGIXKpZBYiDH8dRu3tjEuQ/nrTDqhwyOsn7zjM77u4EJiCjR0kHqWWe18mz
nTP47TJ0Lr2TqSkjw+vBwJVX+anLw939kYVVVMDGYqHf8UKBMxQrSPiuW9ZL
2Kr9a4Na2PUvWevSo5yajPqO0HeFtUilOxCKXdeGMIkwmYOLQRxQ0Msu0ajT
ml3oXn5zgtponORxVo7rVJ4t/dlC9cCH4z35eZrIDRjp1JZZjhKXrIEoyYd3
GgIk6YuY8T9MrusQUL5ilR2v9UKrXun3cCrsFig7A4yIoJDTlBoNUYtm8ziG
KKACz8gv1Q0WRwOhTpW6c1O7U/oYALNj836KK0omfGA6XeqqrMgXOSGdbEcF
Gvw9QtIp4wEOxIQvIMODakIXbc7c3sUAXVKcSCTyNxYdH3Rofs+pMiwC5jMn
KUX+mnrX9d6zB5dMfZeL7D3/XNlCcLHQkTFOra1lOToDJ7pcZbx3Ibe1f+FH
SqXfJ2AWf7ad4GY8BxLXWaG/Lw7jzdx5Tzv+hvGxZ2ZjI0GUni/iPe/l2+cW
mBXII/FgdcWwL4D4QuWBaPEwLYPi+r4svPcuecQX4mH7r4a8+u6XMrEJIM0c
iEYlvqWxb9s0CqTQw45s5UziYdRxF9FXyDfer/H6BqKWEtynG+6p2hKqlrGw
UI44iu1Ukf5qOyPcdHFg00lmAy9Axi8BaM7CTMJDlIotKoQNgZBb/e3kpLiL
d6EQXUvDOnOWMafEDRR36fq0nXDVWcz65Vf8m6QGUfzijmlYIUAIIxMl+zw9
YFeta495Z7Z8f5dSw4Kcj3IrIezTvtVbhLnG30Lu+VgcOHUWE2c9CKcOpSq1
D5qzf8RXao37hIDmuTUFOvVRdQq+2WlD3/VfaQtAkQjFZg8hhB6pTN3EOqic
DStqxEqv731/MiotcNJPLbMgUcLp9GQTeF9TIAmgoznoeVfSuMYchSuxt1cN
XJDTlLpRh2lHijUUhlBIy/omSbSwi66QhlrMcTrzx9A/TQE+3vAL8jxp9SA9
1a1B+xE9igRr1DOv8JNtqEL4+kvFsrms8Kg0KQ4CPmfvTWBnFEVyf9VDdtIm
1RhuqB91orVVCSQrDozQlIenVPnoiiNICCvV9zuaJVOW6UNLJzigDhAgwPmx
NjIFL8n5LXXhaz1OR/qf7czkpDy6YWGGwOdINUYXUfWDriyPgxGoaFyORl2N
37XQjmKwCRioiA6Lz1/l7rXGqXN3FOKf/nXuY//DBEMwA/qZUMjAp5QnpgrQ
/XeIuyqECH7ahVXMiBgwieKPSm0Kwo0Tcnl9q8lKWqq5U78bWl4USD5wktnz
LSXI8q8Um89gPAZ8Eh7U+Pt3zeqil9Qa9a3mTs9bma10KfRfM+Bfh7u8Oh0V
202cEBGiIOEMhzYabsZJjVBdQrs2n5Mm3yyuNvuyLhD6LXdp/Do7R1/1S3Va
Jg0J4aZKdEl0fXE5tTIwV/Zoy3KxbxCqNGsy2VofOQlJgrruhtNXvb6citGD
CT+QakfpKAPbrkcihEDR6XLaPVAgJNGRJgxAJR8YGYhh4U2Hfj63RtghTsfZ
ayletQ8i0GQHLfTAuOIGgSPwgYDH1EZ+fMSD6YXFv7Icau8ZAdCdbhcp+UcN
4z8zWZW8o8cLNvNaJSlQ3C+FO7zLQA9NTB8aDFS7D0nDK4m6rGu3PeSnD/wq
ZDmsnw/z56xFpQ9ndztNFSBAWwKaEH6XoHf+nVwvyBRXT/jW3Cd5Bcio4NxZ
cHtfW2ndPfBoubHSfx+xcW0cwQXa74R7RL+woMveSMycGcU0mCpp7uaVg9NO
CheDuYPsHgzNGth0tSBajESXBU7NtDC2qNGVbu2qciI8sW6MfP+yepqkeqMl
QTmdc3t+uFUlO2RTkgM7MWcamrwXSrbGySO1pqL5ipZwWOPiqGTHBW+0dd1w
q7SIbNi0Y3qoZqCCNo9nO/2bwmAzkusCUHxcRFzipX21aFkPEhJq5u3PiEBy
bXpFVOPmMB6u8/tKqY3tV7sC3HF2XxwDEajA0Jp9hv6KHivISq3Njwmo2QUu
O9aGYmwe8uXuYOzeB1tkD+M+lvBZ52+EbhQCpcu3PgTET7m4ehMQJ1u4ugGb
NreUqCgXepr93cI2o83F1weqB8706jAmP/A4P/P/6wiZdzCDNCqX6WUKaXNA
ZwRIXIFNYk3KNwBiCh2VaWdLTwiTCFXL+q7fxMNigxvnPaLLDM79KANV87Au
Qm9krSG23RjUw/TJr2tf08D0jekrlDNu1sqegdwypG2qHpmyeXdDjsvd17Ft
98R4/rVNTaGlB8NXlmTq8XrWB/wGt9ig0pgjRbCdIyYwWFPEuhCKH6bLjfh/
WaFxbqUQU5MTEU6h9Lk7Zmu0owahlsMzai+dlTNpueIyuFbEoDALmm+Ae8XO
VSLXK3fFptfuO/FU1tECgOjgv9EAnZuEvVuZwGzWEyqQ5kKC/gc3sjsN/skr
MuTcq3y0eUogybq0Y6HmwbvCsnpWfwS2rtdqtoJS7E/h1CyohMq+QLfoyd3g
zbMgHHpBCWkvzEKaE52UdzXIio9mI27rlzoaxXTCjdcAw8UK1IrrSvjLetqe
SwZGhk7zxzCDxPCImX6jKPm0tgBC9nKS3Dy+pyuydxwjf0gxSeBnJHKW5Ef4
KWs0CrFqHLKhHmoauOIfFb4uNGjxldxjoXoJh6zOVtjgAlwQ8VI2ZSGwYGpG
8lNo0yZBj+iAnYzwj3WFw2S/7Y7VOpN6qe9W0F02MsLqngMi8QMkAXuH2b5/
xF6ODr3mJ4Yu0GR7Z+aiahUVwVN1FAEw8sqCVUao7ZoaAUk8a3QbA6RJaTJ6
FHMNz1D8D6JwO68NeIubycMlPUfr+o8T1yr+RP0vTU3Qzl2J1AzfHX7OGpOq
H2NAXpwjMaHrUKjJ2diiJHhcCOZ+n2LikPNzz7/J3B1lA/UprM/B9tAPUv7x
1XIHJ9MrJpMVDwf0GJog+Sjjm0GbcB4N0OcAeAOx83412GqZnyLnbz6qlXTm
dcD/Wtj0ar8WeMOhIBeO2SvleFAdO6wak6ht9P4BNuqTdsD8wh35vXrEHQGg
qoVruF4PXlPDbcUc/63HEV2Phg3l+IwkBZ6+1DhYXOOdQ+d7fTa73iysm/OQ
vQMFQYAlayXX3MPjhBZ47OOUb9aui/wOOlA3InVNbkvuBE9dotS3IBK7PvUj
cYHGOv0oXVxhRXeKkNhGJqlelW6LrP7TYgevBLgFKt07DKPwSNjJjDICU42L
i/Ocis0SIb66ZGC8h2ZL+ofiPqvfvGgB9id7n9ZChtS2NF3lhl9TOSnAjPc/
tAy5/qurSVB2dkDKQm6N3nC/hVd+ywIYNwYC788JL33yRjqNjOSTEY6gwHAP
iQa0UUfQ0A2TtSQHB0Fw5LRKgrSXai8ix6XulneEz6K6vGdI8Lm3WbC8ED9M
xkNeAqZT73OWvWBNXl9amINmFaz1vDxVwGEv94laUUNh2uULX6uc1KELEQJo
vJXBJUDAy6yRnINToZgg1AKXf1bLvCUGpyzTy2CgTyYFgGo5ba2xGDM5kaGr
z3njC33Hm2r+fLr/mhEb+wK1sXE2cFIbhsN45hFFOyL0pNDpAW5Ke5c+tJcI
rcz7GDIVYmCx+3juPdQwRPipiBsW5Pm34gjPxliXZxsThWlJtS7CQW4blIdG
F5ECqW68vPcPtqGNbG9k74Pw6EGhlOHrPMgkPUYCTYw6HP33tLbMtk1COM8P
s2DT/UkRYbvmhQRE/69TN9JGuGbvnjAoGQTi+jrrwgFp3yFwHD2MX6b67Pju
9Pe8adb58ZEHC0P6KV4DArPty7bsxvOSsNszK9ab9B0o5dxTxVByPajIVW1p
hLoXTlJ/5M25FD4Kun+Zb0GlY8apv1wgQ0TJVaT33BCtmH85kjp/7w3ObHFi
tHkIRWSOdEt5EVBqUaQa/f9pHvKBoEYx449XIVKh4JWy0IcKCaXAri+pdDZq
u/KO1qt2okp8HJSJzhdgCdKvox2EqeRgKO1RreQmMYtx+KJtLMxapDGe3VgT
vaBoLmQsGf2HqHAaZJEHLg1lhtsn/OBKTF2l3It0qkTnPEDJGpAs4TsFno3p
5/ZdRodtV7FLiORc/ykHPbjKA2ay57HaF+rJ2oO7CmITdRn7trULxDCUYdWp
MxylbQscFTZcm/wRVq5JChWOHc8FLq1vOw8qCVcniOqtQw8PVm7ZOEP9XGaa
RZ8QGmNvfeCPyE1ESDz9w3NV8ikX9c52Bbjt5+2jTY69MEE9wiVjM3ZM9di3
XR/IpvhIeI04TClhM1CjpLL9N3J36y1hFBOOoJx/DJF8Fq/B213UzKbZNPiE
6edNNvqvOX7c64r/acqVPr9SZ6BN6rx+Z/jUyTqAbn+QLIp1YpJ8GZYwS2jM
IS06Zb8fH2b6YyFx4+f5lcvJTB00fbBWTcVKCRr8C9F7Bvlxl+eQeNN1zQOr
f18sG7uMSZ28FZU5wh4LutPY1E/g2biHBBCurdPze5faOOlpQG0n5HJlWho+
AvdKmRMf1og0uGYW+FPI8vPfion0sSzVDIhFkkubhgniLPq/LdXh9dXHbHJR
3TjE5OcB7L0cniHX0qz+tcDsUpckI5UFOYKBX6aVDxHVQPGkwCXFnGQdFoR+
W/nDM45mS7iJguJEohku/vvgZXWHlKlkAf+b24wU7/OQkzCYvBAthbCwNmo8
daMYYBiRm87PVSwy3pbwTH58kM8kL4ODHSCcAwRYYHD7B9D6eqGatHxRI/xC
s623Gna/c254+woTNUDWoRBcPJDthviTPoNg4RROItsM9J7qH+bDABP2dwCh
F6PYIZsJVurWq8xFGDu1Oj7IX63bE8pO9MCTYKTA8MWI2N6zjUSe8eNAGX78
PXAJmt4HCUrbEQh5cswFjm76txocWEdOak6IRWwtFhMVXLH0YTiNbtREBhUd
eL5YAhSIIbYoRBuOgAN9KlKUqNcUuGx3ycLvpQ+3jMR+g0wpVSIlyx28lew6
tONAfouf9gMxP2XW+qlS5FNiWCUJ/xAtUsW2o1uKlZBmPIjMvqZ28wdJoscS
RJVJ4xChIY2Pzp3je7j36lGbLrSYP6gTCYWLBDfLeGc6ThsxcwPLnVt3IUrS
fdUOyW09mCFSBKNbgXC6BtDfUNhYfZQZlzcEW+j5LVYnfISHCNcH54gmCXUg
RvJ99yyE7wJPuQgbVQuKAWaUNnauBTaOA6oy89q5YEnpsnNW7sOtO0FjJc2j
wgmkkzS5EDlRtgb3onkiq2li0V31/CCOYxYIgJvsr+DdVY/jztqILLsiwNTy
lKNtFwMnHm1Y8M5P31UVuHUweORTgHPr3o3pya9E5NfVvpnZtZ8CI8AKZ+Db
eiZLN5zkhZUjYR8YH3JbrMcWpe+0YcHuy27DbvvmpvZ1BxPYOYFAxhaIxAsO
pbVdaOOVAOIN51hQsLRlfiTmMly5ncsD2+PyOP94VujDXY6ExxEAMbMZVs2N
7HmrUjaAqwMfG3uNbg/rugEFf/JT/CAMpg59HtxJrl0nUdKm/m7SFJG2RKak
MIzDCpGM8kd/Nge4Ld9T/P+beI+SkVHy5lQjf25LFvaDd2GMpqJW5tOVtCvo
VWtJXNP1nJ4cTFUkcgwSR63ut6GLu5c0V07p/poSDsTVeOvaUFtIFtBcxAR3
3p5bTHDPBFymp4P6QrHEs4beU8WRi8733ksDvGyNt2bpKNbUneJQjUPeqBQR
Jk3txpdCrXXGQnLdgI/F7WDNQhwWOu8jbSRVwKOO628g51hep2mOkoc2DRRW
KFDKIaWQZ38Fe7aEaR1k9RMQ1Y9EoAcVJ1VnD9dcm7S649GBy2YmsZ3na4hk
eOlZYb0GTbp0zDT0D+OnIIU8zo6RfGLcGfBFpUlKVBR0tRcGS7tn3Od73vuD
i5sXe2p/mZtp5hpaj7r+bF1HIP8hSjssibbAk9afOh7F4auikUXJUStTWLzj
MrvnCj8YZAfdWk8Y7eGAne64rSvRsqKtEgrbvkMDmUHDD1Ho9RDaWKIj+YPO
80qSFRtFGndFBYHWn3qw+Oc968VBXJuGXALsrvqj9sIssnCtvqWt3Oi+3HN5
7QHIr7eNbkMgzVW9MM9pYAkzWbSEbOWJp3ClxeRE5SZoszHUyrO7cDCcDYTe
OrKhhL4wmTBAFdm88NKBFX4L0pqKjthaEnfb2ynPhnGYHBg2eeJoarV/r+8L
E0cpVcNiIvqX2CjS4vFwa59e3ve7Up9SMOMsIj41m0TrW7PCfbXhNH+ErGts
ijMBHFujv1296UTz+BVNnTGquYs4/k7bYb7ILnUI5IYxfOh43ES+qbCvwvAZ
YjqQ5DVw9yVgTU9LDN/AwoVGEVESgBwhmyEEPmJHBRWKQdiD+sfPiVAfu+Da
zl6L3qngjVyIdjrXXQrDyFlPTaHdum7sTyB4c6YWgZM6oszIgkJHL1Qh6XQ7
7Xn6AX5fLeJBimbeRqUzp+lisJKJBTiFoizroXpKvnkLah7KNpqw2WC3GU25
C08cUxqf2vGrREqvSLMF4K2K0dDyxxC+apqYhaTM6hJJFs87iTKDzMb0OF5T
K4GoLRmT1PztrB1Zhh9XHn/YhlA78mnUWcRF8e6V5yziIeB9/6sXgeb/YZON
lyTKfXQ5LVmvikIrP2o6etXB3Xxv0xfotGll3aGmoOoxk0IH3/8YWO37wtME
AbcTNjvozK6KjGuwPUdSVp7foOXoMvxIkPLG1ltKHMb3gakXdob3Op5r/Lt7
c5UaZ+ixKNftV79WWap45Jxg8SPis7zwd2yXsjj43ioNQ/qRnYcpzPhMKJU1
oh9ToHPWFcrMDkhF8iqd7z3c/qtod9Fw3FQ2tNh6tzucb7TIc4PgQBU7l6R0
ANAOdRpMurVBdDQ/XLSCvTp1wGGpO4HHXzUXheTcBxFuSFtKSBf5WoP/yWG9
wLEA79FqDuolwGMqYenambe8fglYFoT238czs6z+3hDqErI159dez26LQBNd
/5JsFTvA42xyaxiXao4rwqAtjYL/RJePMV5qS2EgyPv5isSLLcL06qy7nb2Z
sQHnBIkjnixWcor/GFv9m+vBSzbCPRMaA/eRIjZluZoWLB5sStxkArTu3h/c
LDefimRVSsOfrbDgsGy+OOq0INMBK+k4836R5zSIrqL0eKa7Q0o/ASQ1gcYg
rxZzIE8InvVmGFnm+WNngb8yzOcoO91ocoo8426lG8LFSoG4Rf0tf3NYfBTG
pEzs+zv/QO+JIGmRHE1eaC64Jiu7Atm52cx3WuG/4bREysx7nqVESeRkUvpj
iJPeCGImfKrU/3zDUq/1hiJjxehE6EZLgTZcEWXjZxGy3w0F2UdKZ93ST+xz
sDSadD1xFKvypiIwyIFg/2CIDlCC3yCrolIMBWB2e/kxbZbeWiqqGl0WQnaU
wMCJyUFdG3CCWcCU77AgsNsRBQVQRzFr1YymNQOqQk8UMLHybFmdGIHGtLlU
T48P1XTKQOqIlJq64lqY6clJS3QZ7EtqoWXinlV7SA1gGU+XgAwnkBSlCc+f
7yfiaZEfne0LNY/V1CDGrO+p1R/x7ILTeL8K/Fa+5+FXOjAL+50HXXeCKP68
Tt1kiGofVHdu94rmD2X2dkV9hQCPJR44+a63CyBOuG7QxiUTIurjWQXnF+M0
eEWk6wLJ2V9VJTdk+4IYHNNXjf3UEKxZ9253uaswCz+8l6PaROmB1jxKpGKu
T1PvE3L8xtfCGjBMCipUSNvHOET/4GjGO9K0e5QUwIeP2anUpzd4lzLM3CQo
LJ5aubQpRjIf7+IJzIUftUqE7O+IGV7y2h91fYyIEAvlcE0hv9gAHEW3OKXt
vrp0bzKBvdyYrCls9Mh2XBfYhUSCVphhF2waXN4cBnnOG0iIlb3DySH2TDDM
+vzBMwIBFKcWMjSVpl0eW+r/4BKfQXGokzkO3VxhFzJ9CcQBZTS3z+7NjP1o
JKTdaC4lFY4tyyjg87DeRQjTiuGvFGXLUW8L9++pPyd14Wnm0fUh7rjTMsd7
Kbh7hgCxybDbsWisAxZB+L6n5HWzP5+Zuj4EbgwrCFe8Nz3B1BecP7ssEpJG
bdvpaSuzvPZkeOO8nlGKTlfcqiPoXwl/euPSTVBxmTZcZ9fs6Ejh1foPLS7i
feB+r34H9UScWUWpqyfGObdweekbgjMXt4lMLtkCwu9e38N0yVspYCaP0S31
V3d32u724ZHDSYpL9VN4NH1LNKzAjJA2LHrzkTPzK3Vgvexkr/Y8YAptXCPE
hgOpQfsf6f2X7OKzabhEDzh7VauWz6NgHWiDr6r8VnvF/s6aB2BmSBTCPHJO
2+gWpZcKG+3IOMExLL7nTZCpGT65QEHjr9axBn2xk9yAn9fFCuxv1I3Qn8Io
xzA7qKqlZ0pOKXtnEdhVLGgjLWnj+Jp2gbqVK00rZIrRNd5Fv5JiaNM/OuFk
k61nE3QysrGuGcgrKAf36v/92YQRgX1NPLs8SnbOb0NRIdupRrnezb9yZs4P
kBfUfzT2pPefAaTINnyZHUGJDvZh1OOwiwc45ZwJKInSwOfFBy0Iz5oLtEWm
1jNDpld6Hn6p92QUk+PufFhVStTQrtMYuigaH6CbGhSivkh8KkNt3m80GQCJ
OJS3Aj4gfGq8+MQPLI59AMmSfu0dDR4mFwbpiB0jjJYXAWbDcOjSmIP0G6Xq
Nzg/9Yl9ACTfu7XusyFAjmmlksnf4mnUJtN7/KwMoChiVapaVXNBHmxBeYGM
yqJxaX7s/nYDsQAzn0fU6Uk+k2HiWf4bUI4Iz1CR+CbkxJq6oiWpl0TH36VT
zYkvy4ju5fu1iufa05ePFXiGcS3EQPovFPPHEiMyAak2/0Mq1NmTz1ZsuhCI
GwJ16rrPgOLbOtp9WRfu3cz5g4zIpFmXEz36ukKONyusaqWS4BpTQkcPBTjL
+CdmJ4HbYxEr9dKm5kiECNE/uB9EeSmWN6J5ltB5SJmB0U/voBUA+Sikzky/
LuMh2xPXnEKTxrh1YcEVJLkEVGcNX7Kbsz9cZ8iAd5YnrZ/S26BUOSaEj/kB
X9yBaJIqDPCzonFqKMEOW/8XvoKuMl4/vV2+J3y+jF4+0Jo9eBXNeaKhBQIW
e6f3JnKMGpUGQLHOpkCU2F6Rc4gdmzM43nF0ndfgqudRe6Rnqf2cHkQQoY8w
qaG4yRzc3XmI+77EUBKmlkwbbB1m+JIptxmze7msd5flce4lpxvmvFRPZSyt
QZ9ECPAEFffrDEiiP+m3FKYBhohsIJX5V1QjWYuYp3XsN3S+PVsve4AQZKvK
Z0lWrvnfBjfHRsDs6v9GbwRScnS8dONnhjBQEdf+kF4n/kKkfLLWB1TYuRBv
65Vdhdyjup2IumCOk4cDSDl4ZkYU+svvN2M5V+NPaVRgeWmU3mNAlOhSMcRS
batgL2PHxkhpJOyuLRLW4m6f/PjmZejkUtjtPp5Yyq3Dgsj5wagHJEi4LBnw
Ii1GUxNTlrO/KcFaiolZtzE6U2S7bVT5v7UOgR02VjO+QAp06FiwayCRSwfI
2SVvWqiJVsYntcmwbct3LEnlfTM6M4ZXlskR4OGD8XZ/fSVLzQgUQSSgTg3j
FxnJu17bu2GNGhhbEyYxrlqn1ZjhcMZ1erbcd93nZzQPRizzoMZz6scU8dWG
MSijoqsQ0ASlOGLBFEof7Na3jVATNbbesWb0W7F/zm7Rgac5eFDJMY/ntpcl
hS7bgd6+vg1lXr3BuGAdQ8RKek/0W2/4vOZRYHFzMHOiRyetzKfhI6baFBqQ
htZythaduRCGAXlCV6EeMMVaGj9GyU3xLt7fzZHv9WrhUYtWKtDIjtePI2YT
xafmAuXpKhushN/ywWRKN3ShA9dqBvPscJHlkHR7qIqI/Ff7Im0NbYFI/6Wu
WgWsWhypOr6qot9UPw6c2VdcTTwTOa7XZMKtAmG/f0fHpRVVuK7KsbHiDmvz
5bX7qdAYwc2b/MU/d+bR/KndMyeoEmbv52mP+PbU4Ur2FhmVTZTfxbeSYErw
46pl0gkiv/bsaM7dPcPTqefs6x9NQGu+i5tBlQE1Df0VKeMijNPnB/wWnVL+
Wi6zEx6/dUO8HSOdz1P6o1XHcM6i5hTScn6iQj/BezL/+7bJofW44irumSAW
URMr/dZTlM58e1ksdxzygALA5M2yhv4j0GxvZAi1C/PPVdutT8jX7MdfL/vK
S2GICcgNuEHSNk3QsPp+Pt73oZfnaw3Pksh3bUAj9Xlf6ruue6s3J+lrxUMR
I8cqtoUSBgs1JI1OcxVdyFxVfic7TomZUWVVjO/N9GXz2DwsZpJytQtxGq/O
toBLielAGKW98vJ4ie7lNdpdIRlXBkrAir0S+yPNNZY+sS+6YuYUXHqG8IoL
gI5JeUmMgyjjyreUV2K6fx6xazftcWPBein4v6kNwsUn8zZhSm3yZgmJHWI3
IDK8/2RSHJeeEHi2Cu7i0lSRgKQRY+ft83rBC4KQOap6pU/WpErnoanRmuy4
szllKPd4pPFBanOqiC6pzL7bk0D0OUT8ez+3aTtoWUKKBisV+y+2lVw6DZt0
Zf634gchAaRqMkZEg9GQN1f4fczxIZinPC1Lc/swHmUCaOI058UhyFffGgLg
JDujAM9AKAsaRQN1HRaFrDeq4HlKgtkbIAel8gv+FsK4I9C9Mpi1GA/GRRgI
nHvUT+6KijJVl/2Y7FYwdXSJU6WooYMovS28zOxBIR84m6ZQxpKCAwTjcEi+
VWjtq4Jf8gtwMiJDzSwXIY0G+9uR2S9+VpWuksM6mJVQkHlp2LHfhYq5tg7Z
WEvGDnrtn0UlV2HYEhv5DlJxOv6G569rwcUVnxAFW5MtT2REKk0P3cNVdW8D
IrLq3pLiXqnneqG2crqkO+ZDmdLDAgNAbEmtZhKa+/YadLhAmNW7p1dmBjpO
rlk7gGNIvCcs8dkX7t2k5GOOkiOzC0BkTdvPozWoXbtB8/uUjDJEeTV6sC6r
x+/dvAKieJMG3l3OzgdA/S82+pWBPgBmjgsM4mXT0/aADzY/jUU/Xc1z1dsA
pcUIdmlmhhLAKr097C79pCiMzAbZEbFi8lNMhgzIrAPlhVzbdKWCo0Rcwntg
yU0LCmW76UeGICkHStMSv6hVmKat44fT9oV2dA1Wd4kLgFHyXtsXDNJDgCfa
Iv2ODhxC5++P8k7z99CsvyHnaSu00SwTanCQfAj8hu2Jm1N5P/5niXpJtHR4
3kUHrkZFQejtu2vnMxvn6Rep47ttd3ssN6C9Ztj/q+8CRsexghB1sRRBjDuL
1AxdhJh9TlEZCkaymEPYynug6pdHDHhqj3FAVOS2Qbdw0fO4HhxulVS2y1MB
I3LxT+xl3K0YfVtFEo52TfRdoKfqf731Lm9xmwCmbWkmGtgwYrvnK6wG+9yT
B97jBORGDPCj+Ibf2FSLTudO0SvJ4Qep9KLtD05oXewqcQvM6lLe8LHoI9vI
u8SYOX1Zj54HYp0cAs2myRI/TecoT/KwcMEgdYNUtxwbz4jPVw/pK/tYqkN4
FKk4EL6mzk4/AKsbjYTkSvd1m1dbXJGoz60/XcLQPa7VTB0FfMXQZuwUH4cc
p7O9Q+KkxeYG0vZ9b/sG3az2dAlYIcn/gPUnnF0Ko/Izp/pPcxAuDLdMbuw6
Be5Oupa9cwRE0LHZrxZXqI8t57TjnOsyiDkoF2SMAmxIxGlVA4pNV2df7PCR
iGU4lkaFt2uPL1P1+ayPwJR+6yfhQ9HzAusAHGm29A10iDGi6wpPtfsEaUIr
cQyEDcPuLEh1zOma7WNLCFqhz7hpeTr21sInYOxLjpATR2gCeWkvgp24VQpc
QfUWATCIY4WR8rGeioU+R3zPd+gVk9WNqDeI7PP89yvoQgBdnJMHG2mmSAg/
TVtbVFXwEhVULhY71c5k5ArZPyx1hT2pCzxB353R4KWk16Ee6Y0bPglhHgtz
gYCb2wmFcVcOlgKuM0Lox5c7uxFQcZ7wX8QlgpP0Bxxn8MjIks3brP5oUVf2
V7ibXRJdabQuXAazYf7RHSd/2/KUB+qEJq2/Jfh86d5v+RzpV3IkResHuRdP
D/Ze2iBmiqsuQPMsey76uP2FKyKf3GfocA/9e1nmNnxMn7RLuXX9LCE+HqxF
TJnFxXxjLEHRw3C3t5JrQM67xue7WwDi20pL8IB78ddHyw627ka4BoUxBCjj
gbd0DSnm0ROo0nicwJ4c7UFxyLP6BbKvUuMzXSO/U78V33UusifnCr38qGl6
PBQ+nhQAoQAom29lYclmAYuj8HgINfWKG5kKppP9E+oEu9mgP1u1RFsZrwnI
Sho40yeFR6wgewRdg2DP9MxVJPnhiE4+xFeKa+Tn2B3PPmNU5FqzBlM9KHYs
flJJ6ZjC6kOSu83KYSihihA4Xk6gGOtALsKfyC2UJJDS6zqA97lcu8K8tfFA
BHkJBkLMIQa7GkkhrBvUuZI5MER5qrlLcTyPJA/vuRPXOpknDYiOjIb4rirK
fLPcML02mBzF7+dHXVe19yn3+XArwpmH09neZvtuBeeEnBnJu6KOpV5JdFEv
CeX6gF8kFbEay/uN3zaAhZvLGCXNvXvYUTgj81uw38VqtnZ8jhdvdU0aIyZR
4IaRIg3urKIiD1jQX5lw5PvmhdBHEWv9TSqGQBlcJzBZh2qO0gGGV4cuT6p5
3CNZbas0HerX9rgzGi5RqbREL5JTPEFNFhSXlyEJwNQRIQ/Nn3YpsUhAWqk8
00cCwrfVy3/SgXwqcKnbhgT1cowvdLf0kZP8+Kftu2PVHMJg4lSF9AT/TUZS
LSCg4Pc6Ecvlqpl+ODwgvkxI2NF293t9YRLQwxjpXtjCN6Oqy9cs+73Pl+r9
+pFTYF9+zGL4ACgqKuye3i24bj4s/zITvnlvBv6A9/gkTkAAZPEGb7JB/hHg
yxXbzxy0uQDIR5eb60jY3DJFSZqGVkIyE2J1tz8CIFzaFUO3V93kzHzxrNhW
cSwrxQfcLdhCjw0nU/XzrC8EpAyS9nChwAXvF1IdioAHfwdvJKYi+jnlWYHc
WIL2o71PVk4B0tCzl/7T3Hse83a0K4Gsehn4xtAsXv1Hv/0ucn9mUWhnlFmd
1liiPBSQPt9Gc/DrD+IWovn4mcRczf+P4Zga4B8UiYJ4vOn3xJQgDwyVrHD9
P/fyU91Pzd2Za0WGJ5Sm43yeNAehZtXzAn8/j7hn5c5doGwEUayq83RrDM/p
d0Y91bgjP1dsJMWAXGM83Zn45XG4bchJmuiwErgYcSUjKGCQDkIpQxYmZLC/
aXdmRdR5CtDw2N88y9G29g6HtupZDaynj/BzcLTkka3i+S0MgbvElwaMIkIX
Aw8ycGgk63U2Xlk6X+uiTKN+5IBhls20bn0+2LPcoViP9cp3Psl8hfz1qxda
cHqwxjGELrBQ9J0LQpsaH+q+FWr7IwCRM1t9ePu4cJ4pz0+E3hztCfm5d7jp
JMlLE3oQ5FJlMtkc64p27MTnC1EyAt0cGnWRJg7YrXrItZatpXLR0zl5DFSm
dIgk0Z2+KgnbNv9IGM32Gg1SEIC8LoY6NtUsp6oGuEaLBCR44qkgmzGHW8y3
tN2/+JcU57LLKaPtITXff6e2i7WVQb92eZ6PjXDkYgZPWMBgNl6sMwccgaOJ
n25OPa7WF+zEgR50ynI4Z61fMAuiwOD9vwS42UN/aJsO5UnqVCdF0h7bQQa/
7Bv0vZpSScg2z0gNkrM9baeDxf72QfaCuYz1M4c/yqaiwg5/RUcMxWD9HDuj
dWE9UrfdEtS3n38MLb5man4LtiCzLHz77zKkBNzmbuer1X81GT5S519TRzld
+lzjOUoKZkZ2vUeoOdlHPpJdfH1OnL/ugtk10uX2qBVHfnaOq2yyefTInp3V
T4cDav//7y2Pc723KkoZDuYo30to9uBu81tmSyxnvW3IhLv1IHloqDYKhyfC
MLA5ejFPPPXH9qA3SDMprmiDSaI3D7zyhZyb43e/vA86TJjDT39HYvETmDIp
iOy6Lkx/D3LUAq7ipHrpHpSmrgmm3MdXAKpTcEYGkKjMMUEyS6vxWPKpDKOR
XuwdyukFeTHK2LbvlnjwTOVrhdBltcmIphxgTxIUc4BD6hUf5iciB0XeJnHw
nOLC0PRTB0MQiqOPX8mxH5CjJexKuXQDf51fY1hOlWOhowVvIPrH+vSj2T0R
0hWZI9FNOaln7snTv1QKArSAY2e+FkfGS10/W8KoKgZzyDo2nLQqyxMMFr8Y
QT4GrPIXfcAHM0kB8+eswGLt53x3ia2bxyDc96qJA7gkMSkwx1CRT9MNmBAo
Pg96e+pTePnb3+HVnAmx1Pdg1UZprkRAX7bL97jKd+mKMQkvT1RDdVewuxOA
6QzM8iKc51x/dBTL/VXPOtzsM46PkA1YLOTRcMEPQonTwSmB3zFkQVMnkTaN
WNkHtoshxR6sDIufCr1di8BVFUJoijdAtvow5SX0+WhqLrPhOkMkQQ8LC1Fq
f1kVD6zzDPOHXnf3zy4jHZb54zVWsK256DfrTmFpCF1ivIzoq4q21LzKMKHg
gQcb4Td2d4Eth0r0yZUnw4B0q+x/4M9WF97GYoPLaoGLzpMcUAXXbf1ljxxw
cQ7lJFoT/NWJZIFOhV7j6madf7S5Y/sgkIDQXpCuGAwgr7tLUhHcZKw768Z6
O1Vk5x78uGTJObWzgh+nj4m9hpYQaqHdubcs2KQutFG2YosPd27cHR2CrJVM
7orKJG1C3QJJM9rN9Lm2snK8fW0drDilXHrrLnJppUvos3H7I/5TahDH3Lra
nJKXrzSezckUfXReh+JiH5/WLTecXPmu0X7FZV+QGrSsZXtk05W3YomN6Fq1
x49mOhAb++/rBq/sTjlHImx7vTKDiks6vntxMER3mSco11qLFNZeYt86F84O
q+RRd9lJjNzvZc/23HROBxlABKDCxtLrUZhIA8yk+bF4KKlsg16+uRai/vj1
fK1kY8Ic1VSrsFqLTtjCgcTcjvRQk/dtj6aW/GQpbJbXVVEoef1w6cAzjZl7
JzwNCfxFvI348Ufljtq6DjiYjRlE/lNHbOLj1I+OFE9cCRMAYKjjRTjbWrvg
MG+DftedZpK5oGEihNvAk0eLKbwc72GvFnapFnhVd/z/QaP42TxWDoSRvqPQ
kZKFS04payh4ucKyP2M7San/T6r+W2qvwRhoFNNiGCNC9KLG5Vlwb6iGMN5Z
lCMk1VotvliUqa4OBBqg83r0NLFaO/ZFC7NsrlDkOI2bf3bkgbOl0XGEU0x1
PzYcSdXod+oO2MfHE9/n4UGuxAHbUK1aKIOksgvmpavRBBUkL+Phcrd5RDY/
Jd2+1lHXXpssZmEsU8r/mz7r2p3MY1khg2BeCgL25WCHABb69ONf9reSsuIf
z/V+QvVkWpPBuQh9FhQj2nxKfkuhjljmlqXNFyg4dOp8WjWkzecAQjPn7iIa
JWixmJfm5tkln4v3ThnktI1DD4xiSTK+l3uVNo+rqAJygQRZEloBuiD3LQJB
DkPCb6SwHX5d/MupifHMCRtgKFsENQNGIRpXc8OAft0jfl8Ds1TTSyHMu4Kg
e3OSKuQxLPQFPtux0D+eEOqwkLxqMNT7xGqfBkNSntgCJqdufbajx/vYu98b
vZUxVKluM5WgIRtcg5iwbuGTXYLVpyNW8QnK+8qIQe5w85KMbIDBUCQ2k6/A
I73KFCiSPkOnx8h8PRRD0Wydtnm/1J92AigAH6xzuO8VqXZLdrEEzokwrGmg
MtFKBDMWJfJ5I2sJP4MCLPCC0wUmCfwtEDsPPK9zE+kvzgbtyIy4fxorX91b
B/LNQLOLk1mveMXvNjo3rD0HRDJbyer//lpaAkegxGx5J6IlYiCT1z6rlhb9
SZ+2pQBZetkw7eOA2UnOjEwaFjgj+/QY1G5x3rkbZIR0ChRhf1GyTwO/5Fxg
x+JZqvFbEVDqIQqsU+leFnV1XEjzziKWfA0DipTnSKA/edFlr65S1zOUCMAl
XY6XtOInV2D39IVjqfrGhtfqawHLNB/3C2dq/X5F2G+zzuniMLrFp93Oy8kW
mFzH8YlrFTUGuqz7QYZdK4Wo9vBGa0B2F16IHAbjl6gWbIoWu7FW0BgCEpwM
W5yA44FgjGGQuLKeAeX4aLXtRJR71lNE6AZBp8AW2zrPld97gOHEfKxxurcP
4NI3eMqvlNISQE4L0JFi8efytUuYKxQIBMwT5pYJGdw9oqVra1jz0D0ZAtLJ
JLjBZpdAkPQUU2gdkCDnD7yKHkOL3uK7rHHPL04wyaA0nc/w+QCOaEnF38Tr
AZFspNwIFAuUs/9jgjUyEWxsYyZqzjH1ZvN5bi4Pl8OPFw6NFuGgCJhMKtYp
Fop4yMQu4opCZmvthj+Iv5ZhQbmtfgRldZs9oCydOrvm0INlmZtvXwRbWHzO
GKnLpThleOKHprx3xR8sGDqAdMtzYvWVE93p0F/w7nN6dXXAVktafbLtColI
RKPDImlJl0ToGOa8rzmR4EF3AXYGrBoZEp1Lbn3a0I5E2ZXnQgabJ4zbyP58
gxVeulvUtEWSdVWey1yom427REv0xN0Q8QHpTD2ElfeU8mBXxtk8gBVqe6jG
Iu5uS5+1VacimLvvXg7cH0ZmOocuxPmHHjn07bJkT59m6jbFBEI1bb+U96CA
nyDZsCEo589bQ74oWHbugMiYlz5HXU3tManEuqylfbSITOTaf+kw1QD8hh5g
kJnX3Zsh8n+E1mm/jbFQP8xohf3PYYK8lzNzOQCghacPBTR++T66QzWrZhLw
HK/xLdeujO+Nf1zQ8jmRiciDCxUH3paPSSwcPFhJwg0zXaEkyf5EKdJ9P7Py
j9cdQCIXJETRPNMhlFTvqqcYBdUgPS6Rx8uDHiX/6sVDns8MVYk1kd6qokSu
zx61HIPWXoKa+1xI5n3uROlSWqj8GnRa6vUgoHZ97u39YiyPf6lhEwdcHdyp
SbOk2poaoCDCT7OLGr2L2VZchuozlNPFA9lexJBL1aCeQl0gNhtKsgH1wlXz
dPnZ+lekZw7w6HIrPTUYP7GTGB+PPyG9hYu1aYOJIKF/PJwA4NJ1yfTsJc9X
/cJZStF5T6DiDz5BLYboUnwN1tjJCurKhtiME3qGgQLnfVFkDkIE5fh/YEjX
V0zNICFXOqsKcQt3HIj9Kp5oqs6qE3wDgqWllMpLCTS62Np7MjsMJiouLfQf
zAN0sObCvvZp3QjRBYD+m8pfZvTs3cH9ZNTQ5zVNkaIEFGJ9fW3YIqeuhvst
sllN9EO6hYEDstqdIYwpEhLpy9+lC7UnwzOIj1Tz+ZhLWuHrUitAocNNDQmy
Ae3KkvRVtwHQVNBqQaUvyXXZL7IvzDwgqKGVr1pN0rygO0TogUHb6+BPL9rQ
vFLKPdeABTlvvROF1irf9EhXTbXBl2aatnoxDu8PRYgZfK8HfG8x1nlE/DnW
kFGkDngzizJk6s1asBxvfZqKf+ASOu5wHfXAJLBvQyXRwmaFSvnzJjtIis5w
Aw+KihP8Haoa1xnF6ypb/VpCVv5BdJ3VI3hvJYM8FiGtCH3WxE2kZRjoWkgV
JO2zF3CHHmkldbEhP6ky40jbLTe1T9LsUFjy/LniiqHJOGJHUQ9HNnzXa5bM
HitVZv65MXmLEH5Y9zojIXp1/s8iQ0iuEjMV2GMGovR3zv/GBOFse8/COpop
2X3RlAk29GNDbFQ3OFL42TK2p79l1bb3aLKMbGe5bM/j9fy3vmhiiZyHksjz
Icp1928CObthEM1lXcMGcl2sMY4vs9ZmEhQhlW1Petbc6JJWpDRqzI5k3vNL
jX6ylh8gX1VdJPQThOWIr0cLeoTzRe+Fuv7i66piBI79/s6/W+VQgssuTTQc
WxNszxgLXNbUxradmVPmtEgVE3qbfCWizcEiEWX4whixXwgw2sZlantws/Mq
mOzC2SU/CcUkNMwuQOerj2w8GHJXa/q0TDr2iX/b/6x9A4XOjtrBAbpioCzx
j3Tt5RoLHyaES78Fuymp/JuVuWJuYbyukgWccTi61TXalQQf4hJ37aREcUYB
kU2O5MMV9zB5Oa9eNPxCxkBvKl4JJCWZkDpVmHZ6yP2WaYrtjiMDWKseC/5i
tU8WH/Bu6k+psiQv7UvAUecCz8+nJ2Xy9q95tEQ4ZHBnGINJu73xtkd0aBz1
j3ueHOQ6eiOzhorAG8KZUMOe9A9rvAT0SL7Tcdbrrwqw58PVn6bnYat7UC/h
q6ZkzomZvHC2QTMHBjEv25mrzCgKfyoiypobQLpjJOeqkq96KTvHISu8ZJYD
dR1KfJUmajU3nbsz9pu8kbJQawxMk6htQ5yAO/6p5ZtYejJNKcpYtTYMeo5u
+Es2GgmdnsyAYwP5IEH8QD1Y/2/M1QUe6416AkrsZlcBGzVAsYhW0XjDZSDj
vwUhkBQ5qSwrNx4wG3/ID45ss0aMwWpbRwPJMlmXQVcz2WPNTdaWtfJlSr+/
lsn/WoIBNRhy77xuj9llf78eE8205LwvdoPiPpMIcBtU7iRYXjkiocCJkVNr
oWTCG/Jg6vaBBjS32mFvwEOE9g1ogxURja1r3ql21iCzEL8XTEL8gM24GkYE
HIslewtcVNNPkKuwJlN1RIgihsmbthgt1od1qvk/DlAHI6xU2zB7dzTl+bm4
fL0nWc+R8N1OSbM6f2WhP2OUMatWSfYZUgzCOcrF932VkctgfK4V0pCw0KVw
PrHfCuAT1b4252MAr5hZmHWp0OPIDlB+zGs4P3Z7A90CXPa9rIHecz80mnlp
9wxJsw/zmiEhmicz4lRpCEKXWrisFKidLreI1owZBfSriJvZ/Flug5o5Ivwl
rSb1LTqJUDyT5TxfCUH5b15Dmq0EDLgV1jZW+LozuvpsjKBBQMMOsdO3H5N+
5JK1RQa7jQtJT8acZoqL1BcsmdWFmU0EZVG6noBJjUi/c1iviAYoR/I9GsBs
GoCt9OquGDFCWlyLKi/BDPUloRs1bbeNKdhLXj723VnZBxPNMnHq2+5UnKdP
nBZJiOn2vXdGa5nDKKL1jwrkxqNW4bRbMZTwa7gBvPxaYhSokz3xH29gooXL
YiuVimaY5LjpnMWw0SHaVIeid2+xNJNuPeEMHKVwmNolDKAQzvcMX0ihqxxd
pBBrKFSYwdT/lX/cboTo29cm/njpkig8GY2LPqjOgW/FK+xt/rTOIhOQAndL
1B+BEOqOHdonQo68sCH66VkWD5mqgq3evWsDdd1fgSpp7azgfgA3FP+h5iyS
XF9jfEQV32AKsrMQcZU6U1nde+mJm+PBb/dmUCbOqH/KJVRasY4Qc8WrXzZR
sWcwKu4WECHbpucDg2eADMXvy+C5jt7DZ6eK/5P/Q/y8wmZ4ivm1QdoxXspY
HqVDB3Q/fsPRtHTtqXIJAwd+W5h3FZ2zuphQ8W2rd3orOWCezJWNlc/QjDQw
XA07FIe7+FHNoRMUEMry7B2XTrZYXsZqEuASOOvdb9KEJuMq4PkXteuZFSEk
3xmFcUdW2O5gQ612jKwotoDAgAgdPRPi42ffP/i+Fm4e3KwIhqKQ59a85zer
HB6MucV1MtNUbiPk6cErmI4WQ8sXoBQNhjSf6JR7/5UXz1ISmbUCAgzX4BHF
ce6DCwYSugHoKqd15DrLtFyrKwzL7/Lj/zMNLzsrkymnBmiPpXbXsq01HNX3
O2//+8cqOumiHgyNIoRoMuE2HSPel9PwSXAlnORWZpJyU0ZBlYW5YKl9JayT
JTHsXH6gYA8JXP2CNZCOFuQo/j2v+rGWbOFeys92V7zfgUI6hPB965dsxE75
84EgkWbLhlw0C6No0FB1eIqK9VOT6U1iDcG0UqvDH4kFbHYZRQJYHtfoMTdU
Tpp2ActVxiNtB5HbsEqTYY+/wELlqcqWHaAgSj4IiRJjEOKCRbiMnZQ9NQjh
FC8xTc7g154tHPeuLrYsMD8ZRZsS6ysMPsYIqSHIdkX5oLDCvw4FuLtSE+fE
EsX+24jfl9C3mpE5AYNxPc/l2Jr4LHcPR+3TZFUZv0jT0mOjpese6qbztmoo
9BJhKkJX24LgzcU3dQPznCpMJKuV64VPDgE0FLk1sYPNu/LZ32bdWGhUYNTw
2Z230rdlcEebpfa0lZSB2YUqitH61TA2WDXjo0OQVpZc5zYvCDgaH0qQRZ1N
j61Hypbrp4iT/1cJTh+86LUbsdgZ7GnrRBpAv6iMUV1xhnTWQFIiHFc5KnUw
EtLXUNu70dy4nKngfA8BBHqDvb7CgrOcYYCdcbMP6ny67YKPwjk3H48jsj5t
fBZWj6l425euOfGBV0LcZOMyCmU+hmQqfZS8pfGIEqiGBgvpbd6BXSuLiD6l
jhDJBSOrTmIml1GL+J4pH1+GfBdT9MFUBB5u3z/S1nXPg9CPVtdZj9imFTee
l7QchLXR7tTCDHtkHfEaMWnZQy5ld2qP4sebYBUpLx99TZHkG8kwRj8tAjK2
oJQUW1gHRs62spq3phbqR4iMcYUGwrjRm1nwD7Tw0dA3kxkEpt8oDqIV7C69
IuVYcOER8zDPcInk7qijsVbaA7ZnJf1hPB6qfKMVazedtUAVzwvencPY1lkT
cODVNZf58byibaUC9mJpe9ditx/SlLIUZKTgat72yBi0RQZG2XALBuAGfUrZ
W1GNQOd5uiwOQqBnhDQL79ZIJD4d7FRLvCW9qODfqBkbcA67MCB6p0c6mbZa
omgRH5Y+4GfRVXkzANiZ+Kmz55XrI1uXLOVbm/Lr9zXR17T8RfW33J3Shfu9
J0LZiLiCLHdfZgxYizPwZviO+VvmCK+DUQSltA9NsZ1avPmTxey7q9KxInlI
2vbNyXlaSmxwZ5I37KatvAlYQMpMS1adhWtBziXAopo4sEfdlOVpiosngf8N
Mu+CDii0Ma2y/2jH4QGmzHl+LsbnexXd4IFlPmNu9BToHNh5ucooPHQfWpbx
8kNLTMw7A4StFoPzT/L5ocoMa1oDDNNf3cXOLlrrhpYIaDofqeWx+vvygx9n
+c/DFb3Lwq2EVutQ4BBr9xFbOpeUmiQBwEPgsoESinsMbbn48LHRBNLGVhfv
DDGcAZmvFrbyNk1PR+k2eu+0Ff7NMYytRCS/ooTgb5v7MFyNj9a0TIFmF8JB
vXt1rRBw5hUvpGYBYVxJTTK3TjL8rdddWQakQkJqXlEXulkUCJZMDaBt55Gg
R24Dm8G37SYkqU3wzS6zEs9D3hu0Y42JipRHFrRpHa4RQ9a1iqBkChkHHVWW
empUMt/8fX40Be+4XX2Il8o1KtcAWNOKOKEIMHd4oCim8ZKdEvFBiKwATbqM
zkV9PXMJs0+ZIe0qE6dsRFR4uVY9JeJzGyUXDrWRQScP9piQ6sHVBhsZUTiF
qJ4w4eqX0WnOWAYKmFtlSJSd6FUezGepHNw198CBI9+kaaVIL1ayDlQtfxAI
5gU9D2VA2BEZJL3YZ/w8Nfa276bhNZpc0bgbXwFX3jciCkchAuxazdATASXY
jDk8syU0pjRwD7brR1LYwwx/LJNz6AiwWlpk/Pelc0KdWtN/RhNoLu+UwI9V
74RvpF0nwYomWMxPMhHvoOeTWn8D33nlyidy6oAEtqezzNDYKE8V/b6QqHCo
TNHWmfM4YhmEjnygF7frMQlb61OLTIWca/zZhlp43is3TyAVdfTvgzI92k9f
h866WG4FveYp5OFtw0Lxzoyj8naFeMPRWh++payv8I1sz9zmVIKTGYNEnYwM
Djkpg1r50Xvm7SkOHB+3SUmBRv1NI2q/qfZVB+LCUqnMR0C+zWK7NBiRXc3i
6Aii5Ewk+VMfttTRiGcDTSmadxLrfRD7+z3vGlQTot0krD7w6yRJN5556SWO
0nGoZZn73U1lxdsw6nDUpAsPj/sBuaPMucL8Fl6ptBlu5jGvXu133a/XeVXu
MI+EyGCNuy4GcVPe0HlG8YRYEo3HYithafoyOUukG/+ytfPphMe6nZC9LbeB
/ymXqjwf4yr4pShDqnBD3sAJhPrUks+4MNPLN2FApZJRfzCUJCsgCObtXmue
lmAKc1WICSzrRH2kNCkxk85wuUqFlnLb30ZCv0lBooH6eS9s8lbnZyaL12YG
6VA8oIjvNUO+l3tPDqouzj6MYcqZSGf7HaDZNmULD8ndIHmqtrqNDE1si6u5
5GscfMaIGPwjpAXtJcbyWViD3T8ZmyADzmOZY7VRLkTHdkLu4MR0IJZBikp4
FTyjuQomEQ7H99O1osaXg4CqB7E69k/84MUanh8L11NRSXIKxm+RSqWuTL27
xLmGqVdtnnfvF1E5DSGrrUXp3AAeJ/q3FwGpqWyugSeNTzsrrzLadshL3ox8
M4TRF0NnDXo6Vp5l6CSrE1qGShmZouj7wowRiVImN4d4673m8rWhFlLFiEDw
kkXeWBo6iRDqN1HTY3op9uWzz0HSWX8FuyWYTUwYVY4OcjqKLsjxWmFlhnJC
umDQcOfQi+thPrnqwH46RytvIkGWJiis0NqS37+rt6oGeanblgwMsPqO9mD/
NcWeEnTMFW5H7aHcrcyCb5CV3VCoh0GoQrYl4OIXil3XODU7d3J9F2NHZcF+
68EcxORRnt14QI71rQ8Wwsz/rPIz+XKsf/KWT5NMnzVXNOnEBW7EVpqYOYC2
FEzM3XenyamgYr/WOdRpdoQ9xRMA9Fd9F59WBNUQnbWRn2kYNGDEfR6/aSTE
ILJzormWjDtU3rZ2Bve/jwBSy38mwhbtSTXKcFNP8hUjUbhKK8JycTXculQu
PP0Sabik6ypdSX07hSwPQT0daUqaudBc3bdF+VEFpi33RzhRIaMrSPJwvVNp
oMuMIBmv/vsYPxkgRM1IozJumI0nShvuxCsrl4dSmG2uE9gz43YFQIM+1oAD
hWiar+P3OWKS1SqIHH7yTqIpDk2E3aOl8oEn8XEc5SJzzM/nVmWs3MpHDVYp
tGKKPWCw64NcqqIt/TRpO2G21ItcWTYLcB9CsKzzFPeYAx8QAF7N8wDoVD/p
tSLKbPcpQn1/kTxyzv6kkDPWubIHTFwwyBV6sIyD+ukb5B9403BAjuRvyuXH
47t+P5cuUIl/tLPJXhsKF9n00QCHj5Uu+u2VXm5krFmyuSLUZyW+aJ8sup6l
lpM0IQIMZrIZkhhCo3RWRhRyOcgdKiZ8ZgjMV1+Z18A6Tf2boSorZ3q7Lg17
UwWR6M28eUHEwMocs0HrYPdgy/++MRx0NEV6+yXTvZ5JfnRl1mDgZEomEMCR
qwAcZxIjCdvu0F6Ih/Pp/FV1TXrwb/inWdyz7e3CO9d2P1sdwI9l+z0k3lWJ
EvKfs0PgYh36gQhNmJ0WIa7ftup6j39+WZCjmSfpf0fvF6GFUS/3Hwi6QSO0
hNNufirHD+MyW/1R9xhTJazJkM3CrEyYJzl7/Sj0uKM06IwUWIT2qjvrPilf
xswgb2gsAa8DL4ZObiszJOaFCHxrQtiTga0HSF+t+na/Gv7YT9pdL16wLTDc
HG8GWgWWmnwh0TzMI5IqvVjvxDzfECAJYlokY/+CPhl/QdAR1IiRHY09VAT6
LlXFeqSHIFJsUOcM6eZVV/oS3sLZzZHuKO0Dhe8/hgK4JvlqWEGjDYuNm12v
sjzuhTNHKzdPK+URjYmcei0Z7ucdpUFuGXIjdZh2t2MxldGGPXBVHgABxZq0
5Zi3I+DJsXYn4RAM8TJLKe1DvoglpG9yLB0DTDWBPwbsV52R3sLsRnH2pcPS
OCGqfJhDSENnQZFKDENkwW7rMiF98oMd9rG5EGuaCFsc2Np/aqKFIMZvNxU0
SdebBPHSwo37sFDFdpogX8eA+FatXq4aJ3VvT7BwFvaGEXZ7NhCLisqKVJty
Bq4rvre4Ts/4lI+VsQ5Hwg61wHrQ51zBM5/qvy6tXXR+teVMU259+6pN4I1P
TFs5HB+N9x9dbF0v2tmsCD6OrUAPQNX6uAWK66BPWagrsdwNy9J63WcOUEwa
QOE3c+x7G0ZHVes2TyAI7wI2/Oyb4OmuI+t5s9ABkx70Xb8ZjR7M0PLu7BZi
8tzTYUSbcJovHMjU5xdF423HqlHkLxvRTbijhIidQ2khze+MHLE8/cHnmwr7
iG+epv/2/3dQ4OeqHRVs9Cogdhstg7JVdf4qypHVqenZIgOC9MS1QZTu5hxV
cc5j6Jxfzfzs9P827OJoCWAiHzCzAZbQPDoSO8bSf0ePJnCZJmyYrW6DRBdk
2oYWA7VoG2GJ4drCxy8bdYXn2zDypIAQZgGXWv+EbvArwvVl9mKVQHr3+LAl
Moq8UKCXaGylG0RsmR6bU2/Kav29lNwkD4HbINVkFwz0ZVNgL1+WMuQueb/j
Yg3EwpWMmuddjsQE8Q281eeNaKnV1pNhhnmhAIXBbiUs5+mD16uq6RrXo85y
PUhlTQLi8GXbsYhHO3bC8vdHN3JEdzyZTacGLTEFro0J/EtnHF69uvjKDSgL
4B8szv5Ie7w9KakDUubiipvUxeQtUlEDOCzI1Ap9arPyupZuirftJY3E90nC
BvjPBudd+d10XNcaYPeuz9ztWLCLzcuSxAuLNQgteqHHD17NcEIYPTNN3wJ8
1pzZZR9eMZ0zC0g5DL72+gSKOOsWLq8b3AIDjOK+xOTntsePm3CrD3yEby+C
BO3qJNvlEXWy/G23uQLMF09/WVi33y3eFJMIcOt/SRASp2eKtnys8ngzg35k
CgFpfCt/Pdn7C6T8fOZtnEgkiP6xC3mJ3FHjgVFpORGEQlj8NEVgAqrBM6mN
WEfXdoDTOd/WQg+62Y4Jw1mXhuJnxKUOhxmE1sBoLD9qS7PaypPzJhlPJXZl
14sp6R9uKLWs8g73ucbIeFkxNWUuNeph/XVbNP2w7vN+VJ1VDzWoaTVYh78a
u9W9J9Lxm44BqV/hVCHcyc9KoTph+ZRx49IZ/j2HJG314SmoXtN4LQ2uTJ9D
zQzpYhJ+MxG5R/rQxcdn0Rf38AXJlULQwyoAXmSAXZICL3JlkNURZSVLTTzV
Xc4035SXUD3zPCBYRMN3ueAmdEof0xmsLqNMhX/7yxjRzuHPDNBOzxvNVVZd
AS5RANN16+AeQ3r2YWmG7dcAr/F/+2RHh9BoLjR8M/D575nW6t2Xe4qMpyPG
ryZEMjuzSoF4ZUW3PDL5FHuLKIhvp5f1J/ZmD0uuB1+2P71WGeQtZgwLVqw5
iuGAFeeXqf2qbVjtBM/ny+VjHOPfAKS/c/ME45fvHhcWLmYxTuaSctomSezy
6hfwT04J/Qjp6Iu3K/mhUXI+cgXk6EWOaZOlO1WL5H8zec2XB6oJ+k13IQDd
AOoZjhGEiFTJIEfMGXCys3VwebqKJPpCYMT7Erq/3n5tR7xLoUiY0adDCtJ6
ugliBREgvx4anaRFNz4pSMf9xekw7j4rFBc6Fht5D/Y7CqkzgUmoekx8WkMW
BzLuywnAzA9WxVu682eRO+IsN3mOibSeHgpvtNmVRe+z/4zPduGOuqToYLdp
3zHW7W9hsssZkpnm13qeyz2BmkUoMw9V15O+HvLUn3729wyYA2+UeKxcdIIB
XNu/sqNj//RhCTeavp/Ef2kAxhTX9W4hXWXVpNTOm8GMwgDF+EPgsBt8k+L+
Tj1zi+bos6f3ortqFMIczCe+NFFVvw4ekBYeE6OsIXg3tj/3uFCZyakkL77V
KbuZEY0hg4lRrc6GeeFOrCyfqZge9vCADWpmjGKYtdUOMNwVu+ripixTbmtI
O5k2nrmCIkUo3a7yWbRPTMTHhcMK2C5J8h3znAm+3ggiocvjLFDREYgsk4nB
wKXv+EjTKEjSKfQI+xA97htddBGhj8mRaGEGahB9egZJ5bqsLsq+kBIuRQ0p
7Z8XKTmvY4jMXZWt68Oa3Y1QEoy3Cl7vGLT752UQZecbfVgUebOjRhUIlMWa
NdzKRCcq5u4nZ+zv/cF7PEsEBNWGMltTDYr2PWnIEl1HvIFQxLHUXAannqty
xahzyRmPwfG0WZR3fP4QeT/WuPtnkVfA/Mfr53nW/ylVeewG6QNJCuX6NXtn
meIhRRyyMbPKB7YHrCyZKyREyQ+9rLYVrSVgE98tvNYfQNt8gMSCahlnkOPV
OD09UH6mi3TWE48N0zQc/WcUTJcIxYsZlo9eF1zUsUWCHwmalnlKtAhxap7H
cOJoXBS1ZhfefZpwuUtPbWCaUqvy16GI3uy4v2oo1gRO8CJat/5CfT0sH5eB
MjlXSdIn1Ttu9+Mn39N7b7dopbSHGHepUq1eo/vUHOafvcOnJKy9eqzfglva
ptLM5y69xuV77T+Zg/NTxm4K45E0zJ06aMwppNaIx1AZrUMg1b0v2hrDR4P3
8ntIwIIh3yyNmAMREGXsfrv6+xWIZc9fuiredNC6ZxR/VfQJfvJvuDGueTLL
hOND+tO/He6+ObHpzPP1XUcSwLZq2OXG69zo87+has7dwYQccdY5jgvb/eDn
F20bFKNZHetj4UeCrOAPZeiX7AogE4wduC6NR8cc4hRylVsiAKHGbcZ9LZOj
HEDm86vtXEbc0O2rwuN95acnsOgobDnDYfrTwR8twPaHlw+EcpxpkGH+vAKB
huU+YbreVKbcLZFO5lzgfvjWNIRBCumhNlubIZ03PNHYz9Q+2dfl/+Y3lq+C
jirC1oFZsSFk3Z4CQXcljSuz1hhxb0u3Srt4kGU/58MEj060Qn9IDR79UPQb
SJJAmFf0eG468SNoXKJwIb6Qh2apFdDbXhPZeiH9Yj7Vb5+8hKm2RSxVwTT+
hQOSw7EOTvbVNmp03ZQ7veXhBy1O5iPph1ispksaCMrUNFFuNUL6Wmc9gEr5
VYEuFsY9NYvcw4/9p4QgsUfrIIpM8MfuinG9bL0mnvOHG/CA+gq8NMaRkXql
h821wU3Qgy0jhVew5PvdOw5RTQAZ6OzpINwVcfgQkDAjYKqFwx5LSlM8+txv
G5WcGi4trBk+ga9jGR6vlwMozgaPOPTRs9pbofLxUp7U8ZosaScrDVQGscB7
Wb1+qvHkZRISVUlMmstOdsObGltPZByaiYGoj7JQ2rydHoPIYC+fDQB071Ap
rTyJ7i6WD5J6ksk4wul1RWQyxEKaswBMoCvVpmpFnEl83ZQqCihuj7+GZkSp
s1ZztNcLP52Kq6Lbd4G1nzz7uS2SsS7ofLU8g8z1alprA4XjHhexlM6BoNWV
q3IR8XxYUjum/nplbkv04wPjddOqnD9XZUlzPU1yIMHes001JlZqf0zqBj5l
PDiStU57QRT+t2IV5U+QiSOEklYFbYryOhbsZVzmS3qXcN8A0CfpcDzov1J7
+lGpe+c3LTKF88hJusmDL3m/5/dwMRh1zg+kdNbHk0tBUaWF6ZxTCB/fz8sV
vlni2G2mxI0XBwR7S2QIS0sYhMSoKhxdZnf0mfJtTLUz6nXt52Fdaw/nZTUY
As2NAYo7tmWMZpsjq/AJwQA6MyesxbSWwK/HKEz1AcgTe7rHhf8CDLQQHHHu
lNDZydmlgAuTLk1jXSRAK+ulRynzaAy9vRT+aQy89qnOLKslR6XslTcxyK3P
RvhZXE1jozCiQ4ctrlgwpWWAUSAD0kiw0AHfd7SrhgWkwp0xmkKn7ZSyIpEc
aP+GDjrpEWYKpoplpeemDSNW7eS14KduIp7tgKZ5k374rchGjDPzunXFEnnw
9rOa9laQlbAsIp6INLNq7RZq76iN39eMO3NySvYpKCdqMBesA5HZ+5evegV1
seO2t7ZzkRcdRP0Q6EdIKnj6q9tk1rg6C89ldg8jEaU0uAdg1H3XnDld7xnh
/USIYjY/AeoRIUpqoioQCJtKdWRxyBMFKxX2aJImrNkaKaMk6igcVtbshHlp
wSE/h65gUTBpHVqR3hjwljvDMhmnyOZ6+woyTPrzghSJZNKSsx9584eOz+ef
KIMPaEpzY4Sgudco4N0HCcZTdLulwb/7dF37+VxcskF7tKCYwUlt2tH2TW7H
+QdiRuJfIukwXozUgMk2J0y31Ax2shaM2bqlTS+qg9GPfpSwevMFwIPpNFbi
zZZukHF3zyRjBcU6W/HKpbbEEbkz+NWBmSR1BqTc/2zL17L0L+nuctLDfX6r
N389alIU6Vw8/1n56wMXX+y3QWkr/JkXJsTsgCd8a+OAnNG7KKc+hAF5nqic
hOA6lAQ6JdQFhltoLdDlZcsQXdE6fAZUrnUcJLifC3AT0UlkGQHbOmf8q5cp
JcbJW4p7qMbeXAUOCNhiwJUh6Depx2/fzEq6cyATMWBn4q67kJc2DYBSYm/A
4zPuNAh33jnXbMNf1TxN4M8oMo0O/xH+IKQOPtV9y6IZh7CC8/TtCCnP2ytM
5GmSw5eF9iWfozPrrx+fWzpwVheK8sAcvUNZydPBXGVJqGspsNm9ydxn8FOn
VdBPuWbv9ol9vlgQabmArdSfIG+gj5tkO3CMbze4X7FCURo4aO5cDPb34K/W
WqDM2d29ZrCoA7gq83efs1gQrtHKLgQaKxbv072EJEmdDUvLYVcZR0AmRvr0
nmmOsg6DImiZzn8gB5tN5wV83YkJECNqc1A3dd0M+KG01cd2rnQmWkETWE8b
D8Zrx1SFE8LGmRQO8z0MJe7+yttkZvWTVOVhu9pAKZkHr8iWNps2qpXfg+Qs
3EOV7ikT81Z4jMfA+9SgmS3M4pt32S6GkjYjjaRRllr48xLcymssuEzAv7Dq
IPNQ49SXu+yXfuRU7K2bgMkZVUtTH7eznRUVUzHxmpOqpbRzuC8zMi6cOY9E
sfBlb/XgBxfPPIQybLbiB034X8k571jgAbrFpmfFyftKHSClHoDrS6X34VuA
hA8xhNYoOMre0kjV92JTI3EWT7/TzwQ71PjdoF/S5eOdTGq1nTzhXYxDdlYs
W9FiagW4Sq3ttaGOX4eKw+1Zxy3VCnUJ4xbwZ1A+ySQ/U8/NPhskxoO/sWcE
CgfcTSbuNvxlZhFqj56/7YvXxY3EiT+SDdD4GRgDOf2aYLUkyZthhbX8v/jB
BrnYmPdGyxgTyhMnlRQFqbxcmEwWAP8UjBO9Mu/Fy9PCz+pQoGIfnzD7yRPY
zhzW9Ql589GF+kC+VAWlRU1ca2J9izv3GJ0aMdbWH4+iDAu3Bi1qGzS6PbMv
qBVkOnL65eNgHbYjFZ1o4encTP5q9Gcn1e0WVlgouFxk1TAGS+kNuDFSDeAN
zlTLIxu09iNq1LvDSARsPgX0FrnRHLiawp0F/155sQiXUPvUl0T4MiJ37bBC
If+VI9MMlhe4phn8BWr+Oc8addUY4nemOoS3L3d35GYUSwofJFRuMpASBYNV
9jfoba/3/TSUWb3Ue2QDqEwTlPctFHRr9KnE5igiU0gFtCqpIvncBK5RDSLI
orrokGg8zVuYvSUTWXwuBp1Vbv7MhgyCDxc800T8Mvx+eXXUOK3x4ofrQLNQ
TsAKuhH0aCoHikWkzLltWn3HPbRLlfDQIIbLJNYYa+0tDc/R5iCmy/6ZWL6f
5ih4+NM9kkWPlzUBJtRAEkCEhAA3t8cbJus6MdHPuRn6ifoxlytG3uo4E0Jr
DRbpnKo2xlTHkY7JkPCDgtyfx8VjeVdkSNZRJvRIPrTjj52HVwUZFfTk1SJw
1CoKKT+FEnkeuhe7TNbeL4mNxjNJTz6vUuz2UxbgUg+d+8pEpRvhrfoxGjld
2Jq7p3V6SiQe8SBbbd+RMB0bGI8wPvZN2mgdJmorN5XPPdKKGPuBTz5bMhw/
TlUHyYxB54uBBNr1z4iz7py1Ke7OI8f554MvAWp9u8ElNpX6389CsRnyI5xI
Lf84WpZE1qm62a8vn/jxOV1nxNuI0CYsQtcNK/RzISPD7vrX4DSI/nQBsQbg
bJDeZt91N+V+jJXtgaBPumexGG/ldAkOrpq2HeUB34vaehuptgjWzV/6798I
FDClbj6BhLdkhY+H+fN13FxsY4xDqJ8VmZeqx/O9H9FP0TJk+iaDfFV9tX/c
V4JyRZn1CC3dZJ5+Xc5VQNZ2BW9RfGgImA3vFV/B4MFVo4BEFBavQhncXxo+
quzjAoUlYtFmQSSxbzjqhbVNzHkNZSiEzl/gFAAIs4hr7WX+6T9CeQWABlG+
a//8ak2PTJE/AeyjWdOsabQVWMmI5UY9+FcvX4m8V5Lmv3owlBd/GLtWB+zy
1paQtdYXmXJMzlfEj3ncgIYHtGT656BnFJClJnU1RSfPPVMn6DsE79ZgasdZ
gp8YYFaQDBh2C2QBYevZyCp/nfCnRjT9aH+q6GWq5RuR/hNs9OmmkvxBO6aj
E4921LSsNkw2tIDzD+kTvLV89eepcAsOXoIp2TN7Y2lnm5xOQZvZBA1W5Mx7
T87ZDxU1SfmfH11QWzUITeERa2CLQDA1D/cT0YhSTyKZixrRcG4sZ+SrCeLb
z7R4UrCRNv2+T0ysntHdcssxNiqT0YVbO+9YFp41ZpRrWKLrKJaAOp0PwKNt
/B9kjJq3nDBci2vnSAHZLCgF+cELozXP5L3NZjvOIevXhfImhkJzQjJmgHSb
3PycyzzbDbtq9i5LGaL9DGi9NqF5hsrgvhz6M9LmGZUjrDa5EFJaIssouQbl
SVRhaqLna5KgM5a5Rx8zla+qJsNoHBuuBPtXBSKFMHfZYxtgHdB8fGQBCcq7
OayzLZ+R6vieyMrY84cRA1x9oi3Q7xMLQfSjwfrd2tGB8AEIKf6k8wFSYNlA
uIvlDWMrg+DYhug/eOBYKKjd43FU72vqs0Mu/vTumnlI+iuGUMW1tblS0LNb
V87q8BqB1K+uUCc1e7izbQZ1fYJQVunVhuK7utJEpS00m0N477HP0lHTenPH
lukk4fyFaVzAV2OAurtaCmqL/1GuE1N7M8KeD6q+ydc/ZklLG1MIMSF28TAs
8EFED4bb3FREnza761p2DXya7xsoNxcoxf0qd/13+L/E1FaEhdszaToYBkVS
GKjDI50wJsdq5x2xXIZsexpqD8rbBJlFkRli589uX1b45MRRNBsZKdTQFEGL
tMFf6xynFEyPrwO5jRmwmfljfHd0qdVTVdw+uITdPYZH7CVp4j/OgHjAXkVy
a40UAMp71m59x/krnw+KVjMUhkUQoe5OAC5Q50Aw0tzF9nAFlOfQww9LbQBE
gPAAXnF/C4GAD90vu02u51km38M0TmDGLIXcrOC3744YFxQNmdFWXX16U/K8
WQRQtF4fNmUhMJt/Uh6VIeNe/8tFioP8crB/5Fz02orF+WCDGWJw/zL/Tf6A
bT1cu0scqGGadI0YC9gtTaBWVHhogytgArvsgQcAxV+j0Fdw1/SndtX0Rnqj
a1EirRTi6l4xrvPyyIWjoldqyrgs1oQlPSuIfT2Xl4GmvtdYL/WKZF98Ebss
xqFSiE2b2KBy2m70h/qoi6RKmKuqPITprisW3xF9nF10IuObfQ3yWwfheeNW
BEUukIbp292cHFiMp+aTZsl7SjoM5xUqAWFXZkucN2Q1gcFmCNXc5U4CV4mQ
nZTUPQ062XZDdm89Mp9eg0hwF7uVb8ytOkjdPQt2EmyZzpySIWzYjV8+ujGS
L0Ys6kXrxFqUm1GE0yM9YlfToBiD2+EZvIs283/ID/cPwldbJ5Bl8Obbhx2J
wN/xEXrqtNteHHa+tvQO8R7/Kd6QNIHNrkOqKbicVuAKHuqNVHnJiYD7BE9S
7Ts0Id6ly49YQ7s9Ry+GguoFUHHshhV3GyUyofcHkdPIC1tfKCrZZSFbMcf/
tSEIGakcyWWrp6ZrkyW1y6xwH1b/G9S29+3kZ1hPfxFHPJtNXhdbwuXBe92k
N9nWdvPi5gKxRQXDaW5FTqMpmn7Sk5vAWBdiD67oHVnXZwFmvyxrOQ7kQScu
1+qCo4AB2SWUL0o8gv8Vy8ELfCFHZHY8bysR1RkP1raBPa9+UsH6GUCMqujB
vUG1mr16MIo8NCYALvvpFw0w0sYzgHiHLipaoMRKfaQSp/7eazg9T3Ym8LWO
F4YcMjA1S701cGin2d5sz9Dk2/OT2LYIiCapgZ49YQKwtSiqh2RhfWX351mJ
IJ6wtzsCsS1fOyUIr2n4c9hpkNFROtUIKld8R8NuvwrJG8H/dfIy7pVPAC63
qnMnEQJV6n5JXkK/hONH5HdcjINYv4xR85CkvPVvM600Y1gFpyY66db8fjJr
JgGo4vkFVus5uiUOY2rfscsD4ByBL/wyFkFoNQucXXJSjhkuop/YaUJFI7jF
r2RqQ6X3cXhy38s3+lnsY4jSQtGYEoAGJKVdflKmu9QoyOpks2U5v8icHqmZ
1Dv5dFc+Q0U02sA1SCpCiw5JUfU2IkHtoRv7N9jsuxBgR/cBQq/g0zUUt5UG
p8ZAgMvMXq3nIzot8fITsipOhmQ7Shi9f93H++yLesU9sgTnqtSNJp6LpSCi
x4M7mp8LEmNTTuaOS1kGiavwpClwwUi4LiZe25HmLFy9hY/sHF6cCtV6ohey
JFK0dPecYEUp3LtTwCt4HjK5UGaX3+bMyR8Y0kC0YOZuk6SxwY9OCnmJ2Q9O
N/L7abgtMTAfiSQiP1yp73aCQ1E7iOmebJ2Iad/rpdBIOoumOwtjGqc/1InY
uBNZY7eO1CLuR0mJisPRSuzJeojsliS17A/RDeFd+LiT2DGEqh6DH1dTVa9y
pW1R/9C6c9qeHHnSk3oiq4iyCvT3pSBeyqJvJd6/TZv5rd+dt61B50aoxsRg
dMunltzmLgf7UQz/NRrxS1uqJLfr8jEwawQgnjB8Z7s2vkZYMO90XugFP6vR
75TV/br2hSVSbqhQ8b4B6ygMFzdPN67z+ONfqa/HHdqsv8KA7bl5nJp6MiyP
3p9x1IVfSy6iV9zD4iAvrz39HtYO6q+gdzf+OZ4LPsZHIIJTahJhU0QXCkIQ
hBa3mWl7HftHxlTlqWGaiHpSBZySs7SPj7fYj9qe+kVu0tn+9uQbIldVebKV
ruzsPhmp0JFbe4hPcKX5uccKhi1E43C3/H/QR2lQvy75rtSP2q1h3jPKezMF
omIFCjQQ7WLjcyxVhd8X7tmr7+zLPSqTimS6bMG0GROtiMvTBwThqzEdzm63
fbrwUfOO3bPsmhe4sJWtb5A3XNLBbGQHxV3Bf/3VJTwnGWwht223ffxHfJi4
3o51BIt6oY6jE21V6cAiiM7v/VMlxrz5ZGr1RBuV9vOW/H0ib5lFo0tNVf+p
qnbc7/5XxtDTm6xuDctF109RkLVoji8i5xPXVOqoI6pNqD0b8MvrnltGFPlM
5Fd6l3/4zvTSiQ9Cu2BCvya18h8viI4aTjVhtewWjekg7ZOs5JZ3uymf4Vl2
ZG4ISA6CKVhudc8EXr2a7SziQXlt0v7Ajh1OezmXQG3vasEMYB6szpdhtQSN
vnjhfkKn3YAf093AVSU8WbL/TnqjHk9gt5XpoyPodzwBHm26u/t8ILxEqvIZ
MoWWQXyjBQR7jTSUIXS4md61uGMVS+1dtPvZowczJF9NFTryeT7syTQ+gQZG
YI8k49ZCap6A5CIykwawyE87RcjIwEaF8FIW1BV41Co2QZX1sNFgG9D6T+DO
EB8y0XIV+Sxm2KzYhE0vpvalwrn6w5GRT231Nqn6wCGsYHpzEbxXBdelm5eT
TfkHW0DWqNbixWmxlstiCfTvItl6KUQA6sPdN9lXKnu7J3Tf8fXG5zxTxJ7t
e0c4XmVEUlcRrghrREAe2TvBMUregZma3rc255YHNmhVypdElkF7rXOdiOGK
DPfysO/VTmx9YTQibxrRbWJMX51st16aBu+cc0CtoJOxci4AqMXs4fwtzaUy
AIz7toITCgGNHCiI9apEbKfYeO6QYNKc/i3unABdK3x6jzLkGLVog5FvOicN
W8fMD8jWgHoCqj9TyMd8evAzs5eLLpCMmhe2O4TCuQ+7lLZrTHfzByEuWTW4
E6JNYwhn/xTGXdltCbZ4v47D9RtJjOxP58zfaTzdRr1bfIuj8ISDl4HAGE/e
6dcDiVOgleCZs2o/q2r64S1MrKDRf+s45QvcQG1pZ0XDZ5D7t1YtXT4nWEhw
kHwA4f6NFviMQBuqb9npeN/xkUWuwaATVS06O2yeOvEXLfHKFc1nia7YxA4b
BUKeoi7YxG3DdlbhR2SDo2R0gowk2JZf0ZcSYzUyAn7MDG08FI0I7WnF/Nte
c74aRHer1ja+pnoCT+yW20Qh2Y2AP3VSU+3BmD6Y0P+Gh4wECe7TN+U60Fi4
2zv3Hggs+7pze3VwoEF8z920duKWOh5rzjFiPVmJYwtutl0w0vR940hVETwd
HkMzonQiUwemRfrfddGlWAdWAsoA9N+vyUUCniN5/RGH4GgQvIMyn5sw8edl
V5yiml8IDDvtai4UEq8oBZLffJIS5JaLFWoGgvv9pWUHrdqde42Uv7V8iw3U
aYEpFEIz+/3o+Q22Xnk6G3T24Exwec/7p+4D1e45A9Zyv/IeWlrHI83BoKXI
4UNfl2SlbEOpHP9eJr++7Tlbpj6TMehrT8ZhCj24ExkkHbHyouYdfy7Gii0b
6tZK5O2wo6L8+QEV0nsxJq1bb0G41Ij+ZqTofdmY0oqJJCK5/AzJGSA14lIa
fswj/2z/xNBQE9m/MMiPRKSfYOH1Y8118LonZXoVUKLiy8sG6OdoXmxTtGEk
siOIE5oAz+UBr4xM02QwGm03lLpf1UreFJeetV9fF+hqjOutFsiJyBdksR7M
bfif4sSGrMnAJXhduQdDeKCz0mBbmNX5KdtiFLDvOBgcOCEq5HTfiBjJUwLr
Om2Zqi2PdF1L3mkuYEd2zB6FQa++UnVniXTbD308Fx0l+NqQiS/SFYRXnGw8
4l8+cb+IlO/Zm3e5YV7dvtQ8ksGUQPfFvtMRgqC4imbDYcBlT4W8ddaMmmHH
2Q2enjlUp37WtXaFmf/SKHHcx3sTQa/BQuZ2D3xHYVyJOtheC2e+clSEr9Mc
1P1ev1/Z8TC/apLIuc7MCXFGq2MT5lcKbXRdsGZwoEO5Oc/RrZ50rv01PXAj
34Z8oBiu/Oppk4J80QCY2OM+qQnLTiWCwo0euD81R5jBVvYuoiCgUC5HJARn
bs5Xj84IHkjakTqZ5vRLt/uWTrzXAAQ0TW1xauW7x157RdTZxvS9eCvpONZG
9xlV6Zj8jTJxGldCVE0pb7Z2ZltY/yjeX1yCOGK3y2HDcXN2i0gWDWcSfG5x
TO5DA4EioIcngIsrTHkx0Q3xL+aPIuGT+bEMrBBc3mM6EVi8jhrsH7LEnRvf
RLRj6bgyjecBmHy7y6l3M3FeCyAoxbLncQ9RZi6PBFKPkVWkxxOeEw0axBgT
i83of1ZxNifszdpSfEVI3PbhLFe0Hv0LvVHGmLzpqdkj9TYfsoqMPs2hJHla
U2sbt1oSiPPHa271GExrLj79KBBs8pQjjNGqAxgzP26/XTeEUeJCvfiUjkm1
6BebsCW5JSAOdmnalgYT+Oyl1HKhXnTDGyVEN086zyuM6Pvv/evXpURNoRqb
IIj6XHaL8O8UaHxy7NihtoiCk2THbgEJJdGGZXaPi0e3f//bo23Bg1FaIm3/
wdPIsqfbt9Aj+ACrfyZ8AnibN0rBLy21R4zTcCjrlcbk64lqRMyQo9LnipTl
7ZmwziOOJjn/XxpJn7uJUR4mjMeoIF/Mi8lIZqE6L3+TD1mahYKNzIkOBSOm
X0wfxNUxU67sYCHHadkSGFJpYiwXdo6TdPiQ9hPK8zsaMUBOt1qiZFZP/0hK
/dYp/9W+Q1+xDNqg8sGFOP5zl1vyElmy3oPEbrfU3APErM405YxkHQwrHVpE
ly94TJWClgT61kf5l8yMBTAWF2mLXIIV7zq2akQXVSQ6vITZWoeZ/gYNsgtj
Awf4NkEtOW+PepXLKG4YbKXkY4U7Zj2Pjin55rPud7io91dl1lP70oaXNWlj
vt+mmjdFFYP8AXB9Gjyq+E+082M2ErlduZA6X1vGFkbWm8EnPpSpWuCiDw2h
FK7yJFPUH0+OPaLc2lrFOXCfUm9Rwa/40jAjY6jeCLB/5j+CW4a+8ndjQDf2
Bu4woxDdaTJvF0Y9Yio1fnXHDVuP4Xv6ffj9BQiX1uy14zqcP9CTiK7RDt4v
1h3aWyAZjTPD0mcVR4VsVt9ORu8w/thQb/LlBMs2ygXC4tN37CRJRKhS97+B
9VDTV7cJcNyBusW4WogqlUXXZsppqHQkmYyqtfQ5+ESPbFKbJHnEwXB9K0A3
MuBTr02QuT6gLwu6rTPenUSP7psUh7XZp8IiM3GfkZA0MdweMjU3mnVjHTAG
/Tas2Gn1GDWbAavh4UN3QMXKiawL/H3Pn5zRBjPZHxh7DO3oNYER6cMbHrZa
Iwg62kMNyiZLPvCfhgP5rm/EaNQCKpgT0cmVWnMLkKyLE0Cl1gRBkcfzyXA3
YXQ6+iEDM/zrCliTOAJCS6EVZvtJZN+T7vlHg/LZtaqmOyIg+p0HodAqHEJq
J299gHh0psinReAJAFUbDNqpBVZwmo8tKHYf9wvsfpZ0SqEh47NiVOPNPZdW
rKK5gyY8W5s4GQYAoJprYN7/rFImlcjw/Clj0Leqj/+OFGgATjbOvIyEb8Ap
AtH+AgnNIM9LhzKWQ9w8COZQtbPIJ3p4CUjjl1EMFGZsZgIf0PH7OylTH/T5
yg7IhCVo0jb5dPFpbk2MzI4U0QkW74dLNSeAmNwUH0OdRmOoIO7BMreKv7lU
21RW6Lls09egl6ij1u7Iz1iW384QxV5J+111OR8rBNGUocibkhacd6AfZEEz
jZiWhDSOaOAN802Kbj3LlyHHf7P5wNbmqGVfAebjbcNACpmtZfYkwesPuLYx
q0CBNII4evEVcffpAUYOMmdmHC5krY3tVLtr+SFDgRgjKvKRuEtL6XUIcJKP
FNZ3C9zjaWGXtw9PajTFrUitluTKmLxZufQrtMYcebZTLmBf4+sPKsrxo1Qs
+NVoFiyQ3dYd3EgeyvfDd3V8fMK8KAtJZbUA3m77HpPFHRG22JMuL4ZOM/VH
0CMmC2Jyvmt0DGmUc8lhOgx382IbxUM+D4PzkvgmKNXHaCk0ZnnfS9KiIoKv
dY7TXFiamKhimdkcH8f+rA8zBXnGX5jHd6/G3JYZtGWG4J6BuYRGVINWSmhj
ca0wF7noaq5ofw2Qk7aWYcUj5ev5k70imowNwXP+L+P24ckeBaJs70tcDdCW
59jOdHvoB0gJVAi38cV/dI2ehutfYNSaJVqpOU7nU3KL+9+m7+aZNi4v6vu4
CWuVEcHOedDhqBGwLvbybQoQYVDhC2ep4J1zsLRIQlE5eHb6Tg9S6O7ItaWx
p+VgJM7+OoCt7ACb+YLSzwlYVHIpuxkWEFdApZ6lcWPYOoWX0mXnyFsPElrl
TIoJqX5JZcD3+lXF6mlAHvmaXDXKtaehLAQGGhwIPipsKoCHf2hoOgsi05Rp
54E8QifeRpc9OyFmSBTVJWoDF2vuKxaO3mlabW66FBnDLtVhXnluAt5tbz/i
9GD3yb+MfdwGIKjPyrQ+1559dkgbtpIvKzZk5zCY2lQsN4veHRRQcUe2qjNP
+jBSc9/gaKiCfY2znctBr5gly+YPoMn1hBxB1b/h8dPq3Z4/G2tbTnHobafU
zAZ53URK71iKwnoYqKlLzuVOaDOZdyVl0YfIzlUoa/RBrYiSHvJIrLeWeNWa
mOUfxFnCv7Z2M4eZ/ZAenhJnaEbT7AGKzFtLbB1CFi4p3vzrp8hdzAViebqb
3TwFgqsXZZZ8TfVIlxFZrNEUNv3h4LfNvVw+VdXxIfbM9h4cQqBoTVR8yqkj
wPjxVkS2GaLONd5pzFHRpyiOA5/7ElMyCZ0HHgAvWWv28pMlwaw/OSOzf/he
rrCsw6WuhhWmeOr1uErki7KwlhPQctFmynUmzi4kcUmfNF6kyTDZAqFKK9MT
3ATrlRx8Uf+NmlxMxEL+AEEXgHkQNVToLNTFsuQ79Y3T4KJvtLd4dqsNXj7L
ga4Hw8AwrMtoDUJXaiyv9VonaSXqj3aiFCAg9b3XsfJRFMPRvW//9FKcpKwP
VRoVHjjEZFVPZcKC9Mhxk4lFmjI5UIDqXiYIYLDhnpz4EK1lq1ebeip2xRz2
xuaJEcV2FvN3ael4EhiGB+5QwGgpaxpjewxonxnqa5Z84EKLlNfvJmvDpZLE
S8WyZUspbZKekIXO5X5q6xBxWPSJ54AwSQWrlI5hhSy4VLBlfD55TGPW9Zep
nKydG7lmGvofJfeJ4IL1VoXK106f9ZlR48TNb0anksTQyYRlWlEnAZh/mQpL
wpjo32RvdOaV+8utw/KP+/0lLVrHzAF1xiycKNhfzyhazUn7od210m12xw/o
aXAHef7U80CzjfIdtPr7qGy+wPNIKVOl0pns/ol8J2Ce1pCzsiOjpo3OmBNj
ArEgIwl9BytlIvUP2szb9g1lEh3LDhuucK2kx5IQKWr/CeHGytuYThqEOVkw
C0vez2dMzVgGhNdEgjYCwjP81NUFKDFSCtLT9q2San15b6VrNw5KZUkNdr96
0FItJjPLqd3wfnbqU/3QjH38vh4za2ADNxUN1Khz1KdsNcJ298dEo52LiJNy
OktJeyv+sRwldf2hlSNT6OcP8q9Tx1wYb670/Ai16HjV6tGevX9hjUMLj6Cd
KxnkhdmG9Tg/fxSRV1ZXckOy9vEd9zikzORI8IMlI2pazb5cA2mXeh7K7bQg
BliqyJllUavICJ7G/zdZ1D4718O0WvoPLel3acy3p43sBXyB/r4e2jZZYD9C
TaoyN8QTA61PbzSOitI0byeaHnvMlfptpSYKI8udJ8ZExUg5vy6flmZTk3V/
wP9JLQrNDr8Iw435faf2GqE2DG/ehBOMpL5bhni/noeZuAtbIE2a1DbO/oiC
QwovnfjBLXqmq92QFRpnEyD24BUm8hA1Cf0RDfHZwWBflzQaVvZ5wTZox5Ik
H1n41/DcT9sAUZF0VTHdRv+K46sZeoi94Zm7RTkd8mVbbavTbmbupGojVfMo
dWoZzsYo75HKdfNOPADpx1ox2agyxsQs2Fx6PSkFPHEWEYEFlBpUc2Wdr+yq
rG7SLQlgLY+iG34YDSP1wga7k0gevpUO5HrzmarneN90FKoog4Izk5t/IXdm
chZE8IqLZXiMiM+AQN5sPaOz0P6Uboj8/Wb4BUBK3m1cofZDnHaPtxqZCCEV
ffgcOKwJl/0nR8f95LYbL8fiMbZMGKD4CcENqXkZkAzVbAzQPcVX9cRtCj+p
xvtNKN0jqg6WjmEz63OLk2Kp6gGiSHqhwQ9akg+lU0sTiOY8KxcU1ZgIjK+6
nRZZfINjgzGHdkap34FnKRkX/ple2GFJy3ozT5i2bHgPCjq7eFU1D3n+K1Cd
JN6D38ojR1GL2qL0uBYfOJnadpQGVqWkWUZrxa0VZJb6gBOQKTtR6lDa3Lxb
7roDJ8Pm05lDI8JirQBobCdIfLTaUevqJxxRcLzIZISw1s1q6oP9qwj7BSBE
hr+6A7sXYBbTsGN6X4mBGsCarv45g0QRoqb98kY8XjMhwXtjTcEj036u2gZ4
LS//bdxyLN0eTdaVDd/BVxrRTWoQ/exjUQp5EwRDphTAnFAmeEq0ZLDz8Xou
A3LQw3/IgmStwj/GHv5t4cYXZ4ThKkD2MZ6H6oh5c/sZbjNVLGZ+LI4wFpaJ
ob41WWecCJVv/JAKU/wXI43+AhPeU9BUcCKfhnOaIZtNFpKo5R4yvaoFZ3V9
tEDo117B5sWBB3Tp1M17k7HfqFqPlebA4IOGZau1DpEGB2SXa1ZxdFVXJgbm
v3hAAqkeqMCpN0oKKjyIaJvFFSOvuM6mkS5zpN1jSrWVYp0W9wqEXFLPC4/g
ozm3FCjKssx4MBDvjjidYNYL1zjbeoVZ0hhT9eZbvnoCd1Uj+PUOE7FVeJX2
ixImzcVcKZxz4alpybcYpXlB7yfxO1V8v3IyL3QwXAM2TOVwAy4ZzylclF1b
1DzlQHlnEKqkV0K2ZSLhRg55B9ccC9U8Wmej5kd4kjKrJjtgNGbOCy90+jko
zqLXwo/55FzNyNo7xd0V/x0bbWVSd0DakGMk0bKHLti8+om2BgtL0dUOWD+Y
qSgUe5e3ttsOEnf66y+YNcJ63risCXaMmxNh/Eos6BHgUmtAp9Sy1qG6ag0F
a+n8XjnVauNsUn46nveEUT5kQPQ/XyELlG1fN9BgTfNlFTuTWCg/GkvLCiLv
cB0h/wlKit+a4KfFiKbJQHRY+kX/uKa0AGpvD+2V86O+qomBwFs81qmsetjN
bU+imlLfMg4NDqoRP7rXXyTGAFYzEnbS5jYW0HSejj37uhk0dO0QoFkIwvYc
RR8IRaKMEK460JqDZrn8GcZAGr4mq0Z7ft6SnJtSfq8WlDFoLNDjReg5jYFt
euQhDWoQy5596s8FsrWlf3k2ZePTu/xN89oa1YXl6OOZY1wSH35CijX/+4mW
0Ow1mOzKEAk7Qhfh89+JsE+0mGahrJxVbi4ZnWTbkaLtxkUjMxURbwu/TcF5
uiN9HFkVqDTBj2e64WQwSQ7vWipHCVG9j+J3f4QyfK5OCY5ZNdLyLhkWjoxf
T0CqCZauo3v+J1Vh1S1RjOtH80NQg6bngxjlp6xhGNo4nilDuRXJAjvXkcgC
22EiYvuRfTCh/j2Z1DO5WUwbGWnLshTfnFKAsV9ph7Pga4AplgMt00YYUe7Y
yUIxyKJkzIitTnxnHe/hVubDmDSwTSoZ3Mzg9klMXdlMhIdALvq2ccYWyJp1
FOqQipdw/Q7fsAaGU58TTD/Ebr4/t7KIKdIztgGA12wnpRqiW3DBN8h0u66V
9wFyTj4cYHCSf07vzOk+s2U7+MY+9JRdS49fPlvABYo5FCPMWsO7N6r9LT8f
Lt/5jCOK0L07qHewjWC1gN21qgs+YaTAOp3B0RYEj5Tw/XS1Hxu2ylHGEp6v
z3oC6iKGoY0BjY+IXlya/wysirDFELxK6rD0jAKMq9uLUFd6fSZgBf0rU9W7
0ZxfuRTKome1BANNdZI25k0/+/79x5BgdNIcdpdTMjfSuDQjXYWq9l3UI/9h
xqgp7H4d4FwNxn+LlAIS8jV+v9yP3rLC9ftlDDSAcaem8yFJglNRi6deczqE
mPdaZiX+TKwC6Nzl8kpcOmlG6bphP9tClnTK7IKa8eOpu1x8ov8d2IHC7wOa
B2GGjz46QjTnhz7z/xNtmsvt/p5X2dY0dJzTYMhf8DVSYmt+LRD5OzsQDzxU
CZr/0qEDeD+X7iTOjMXKPcX8tONTpsCAwAKhZBTOGFJIpsOpp090okNbfUxl
hnfC+34smfix5+hkHVTJ0hJXs/fgGS+SKyk/M6OPKSdQAaU+Az9UDri3jG5a
0fNcOsROPshvFd+qG2IBExZymrRxe0+WXHawYARSac3gvHhLdjnZSw+5KFEH
0YQbjvJ6TC4mUpmfhQKqNAcg0ehQSVpF1tSv4sWRf2YwdVyPniofkns6nGCu
BZNgB6o2Y4G/TnwXqNG3by6UFIW1rm1JckFT6pJGoYJEx5Auti83+jNMg4/r
dnnXxS5pWD0ulZbsVMs/SPQwcSJJ1AR8RDMk981sk2tHsq9Z0TrHzeqk1ble
gZ0Ii7WJ/bbQvj/mQ4alChago6Px8RbRN7qzNkv6G9Wh0HRCzWb6MzzC9p0h
Kt/PJm09gEGzkUAVjGyrmblJwUUViGl6jql1XVzkKK9YSwNRcSW+kx54uyfx
NcAT/mJJNuEJGs8V41JE7EP2K69wza3ZNkxTMjqxs0IHW6Tf6QwmvLMeqsW+
tgdSRo6W5K09RQmo0dDWZWrCT21P45g8Ugmrg/QFEDW8lIvT49cDJ0DstOBt
b5Ej5eY0TdL/awtR6TN/uzd4wnuMkMDB08dFbDojkZpdTPzm9yRw/cnBaGMR
mEFbxqp8b7lBUyVjvZk7nVN6A8JNf2851ne1WadlZEJ72I0Edy0OAwkRhC6p
IHOI8eW3T4rl78UIPXmqFH9gOUTyQNdQp4QUl3gQutgbasoiyGLDz6gLYWqM
Hug6jyemNgZ85Ae19SRZXR7VHKqhA4+UkBQOSuCdnHp9liQ85MFn7Ue2hMYL
FcFrzUhgT/9i5CbQpNjWF8wxVHI82njECfuUElw3giJ1KbtXDUdUeK8u4PRm
d87emcfAbagI0fLnfA1dcbVp8EAK0fLDpPvIzp+p/yF+F+YxhPqzikoS2tbK
TQBzPXMQxK6lx4lfEmM6tSDIxCH6Bo7omUDqXZkybh2rANAxh3cLX/hxqExw
zJJO+w+H/0ob1+3EuAHLK2kcEEiYQhkuGZTvyIQKbCQ2hfhUQ4Al9n7sDsgi
qDjms/UJOja8aNUhuqqABZ03VPqyX3KdUGPFzyhIRqWtnqE+eq1iF0rHhddF
VlHOmY0qh+5pk1P+N9GstzYEdCEcwsG3uI+trhJHMv+M1Ct51+4nstCtBJE1
pulRv8HJ5p+Q38iviUw4zaf9vUJ/cMGyML/uJ54rxLVuS6enIOBs9n6Ds+CP
fBPQSy8JhQfds1AmLuZM95oRg2w8yEcjuc+UX4fcluOiWmG78MtdYY0/vFvV
V73ncdxI4QEAYVYt3qZBnwceSLGYnF+XUO88kc7Dg8i5gVOLm7CNzuIKgdmX
rYNIhNhG0EVL7Woau0+tcoVtjkXPKV2xy3uNYiPvJnCKZprzz6uHaIMfFOzh
nSPesyfrcXyO4lKqE3fFXxutb4hE35SaEwuui33XT6Oh2euUeBYC8y0QtAqb
JgQdTk+lBvRrn7H1RjLIfp3KXkSTeCzYyo3TtqE8IRgLMnXHmJ7hwQZ+Hyfn
tsgE/60KDcYbgXii82XkK2HaflRtzDIA6avAbMGs0CrSUQZcomlLC6QwSAKx
AqvWG6F8Uf5HF4zVCiiX5MJZ64Upjc/zwa+BJ0vvCULLzcodxdsWgSTWcP67
IJxVyQRSBPcB+MaXVbfbgYekJGbXGXoh1yosnJSOmvrEF+OzxUc7pciSYSOc
OUDkbpRnFTsoQWCxcrq6TS8RJ1c3J/hNAe3INMZAG+I+DEMiHoG8lvC1yThC
HPrhEBrxvj86wcP79MXC7Ln13VzONlMfBQxaCtGq4w+koOL462zSR4DmWiux
0+qbaTumnTQML1u7yv6OravLdFh7b13qOPgkl1LVsn+SyqbFlyTIL1OTgX1J
xXkIoQArkA3WRl/fX9pAL3BxFmFcw1cHItRSDGUrI/7WoN03Wq35SERT58DV
UE6SxNzRrCuZT+Rhq6RBDaD5rHs3suzQ/QWDeXI06PJhpoWMkYkEdNx1K4b9
1MhOW33fBWxJ1JJkCFdkmY9kVdZTcaBjFAZu/e6wLXr8stsc9PMpOC9upnCh
5Z8eRp08Bc7gPE59CJgTkKaTsyCpihconej5N1VPeHRKgtLR3dGCNyw8pMwd
mhSO/DfZXiBkYZtFJ9SE14Tf7w/7AKK0AuJmBxPzLXitCogMgF3edwz83Goe
usjknJjzr17gYo3Ha32saMn6/e0CtEpc28cKr9KWEHmkv34q31qre7sMP7Zi
jLO/1MnJyAW1LNFSHb4o1jjRMhdoJ1PxKp5YEuSnCjZkgQgYM1G9tcvNyI59
1g5kgj8nbUh+zITUvfK256MgXI2aUnXbzsrMKPL8ZOhWI3hVwMTjhzVel1Ro
6qFZ1BMCXiI080xa525o6u4Rxiur2wg/ACpemRbNupJil5F5NALL/cgocl8b
+ycxhmpPUBGo1/6XuQWVs1bvak7mxmACKj/WaZrygWLd66OLyTzdZGGjRryO
JfyC+1PcR7eFe0GNGDzezL1pF0+41m48LF2/+FFhDZnm6gE8X3w0JpVqXJBt
lz6GTbQwaL7oSCono4Ucwd1anyd/EeQb7kCXVhm+RLYGktxsOd1HXM+l3Y56
lKktBUWyXAmbQMjVG0DUDJtOPF79MU3/Tgpc+v4Ebm/jdm0HpjPty/lG2f0t
9GV0Yo+L53rS8wl2F5mXqHCDspEgQeNiptTnvm8prpnXKiBlWhBijn5gQ7ux
i09eYCfVJo96yyy6UC31CBLTUZsCiNp2cN5O4l8Cjcy27dqYCQkylr0DLdaL
r6j2jASk4OTEoRbzeU1j4rd/N1mg3EMZQQmSZl8LkTc8qNf8DP9TXZo8EOGZ
AJ0fk/94DnkJY5a6NKOSKQJ/Xo+z7LvGmvsf+fm9iRG9oa5WPW2R1Be0Aito
tDWmaqDGYo06sB8OEj8gUU8jbJ3/TC8V61CXzg79gxHzrYdiLH0XxGGv9zY2
EcGi/AdsOVCGbsi55tLwWRNKc2NDaERV9HK+CP14Pw/Js7xz0EsToyTca+YM
OAs3mrE1NrhOhQyRzOE2YOjJAGtBSMVD0syUlTKy6sYHyIYyf2SKTYoNiljA
lwuiGMl7LVmc6kPAcUa1pMfw96NeclNQZ5Cp2ZyNO6DtQRx8o5kIham0kYKi
Ah2JC6Ydt+pq9e96DlALZbzU5iKcUW4o1A1LJ6bB4efAku6N1eX2/0CvocUP
mWTpZbFb9fTS+8h8sgruUcRVa5BB3mC6figVnlXdt93jFNhOB/fCqlrW3tQN
10oQBLMZNDcDufMx+txr7gprrxQUB04fHspnqtbjGnC/ouuKLdE3EVxCg1hn
3Q3xFspTPeu26oBh4epOcl0YOj1qmL2Ks2w13QohJAz9f8cOyAzFQT5q3UC5
9rn2yjyULnhiaT8c/yWjZkPT+gqydxrnPVO7zi9yKaiEW82J6n0GXdMvTFKc
GJPDyz9bZmUioY6xBHNgE6B8dXdwqqCIvuY1se/FLk1vG2rTX5cx8ThdDF1Q
1O0iG3eebiB/r38e97ADGZwoV5tIe85Ip2INoaOGUkeco/KV60yfV+MecGEN
VxN01fRxiGEHwCJPvMYQMd5iLjhOYVwUlmq3koUEbsRLx3eEIv0l8fYdb12l
vAnLpOGye8H35gpH4BeOyUqA2i7or5fUevmHDyEjnwQxAX44yea2KY5NTlWJ
nhyDCESNmO3bSigs9XGqB90hFy+qOXQelIBUN5QdqBS7easxuhhPqr2CM/Sl
CMM64J41EEsFiwAP5CzNdePp9OtrOLGg+VLK8uXgQgvc5V3pBN/1DwDVpCUQ
le9+EEtxSMlI1SdDkJNOujsVi4sFMwoS4zHd1dB0OCS9I+sq2jjbPWhCF8Gv
oYXiu7Q3KjWe6SczxqMdWEwLbiBUEE8sLu2x9tUrXpxPR+ziMNV0lQAR0L7m
9OM8VLEH9z7uacbq55bpLMkeLt29JiyX5AfQeY9uBCjffLQ23M+8a4E8DWiZ
4AtttZOG118/wtVlwLUS+wYz2FWbxJ09n4t985Tah7/2HF/JjaXW3TIVvrqU
E0eDwx3DxO0/H9un1wmoNw9l1t11TbxmtwCIJiXEAYtCMG5I6vJT2hsetL17
zjVyc8CKg0fZw5seZ6v7Ww8Psh/G3YLFVixyiVCFnHYNFs2ioekMjHiAPstF
8vGQtpjiWvl0nGFVwbN4PdJu58w3PECJGShzQqM5UEugKSTtQwn8lXiARkP1
bmFxh65vKw3fk0Z1AP4Yh2N8o3s+zQPra3giXrNCeb9IQGSFxf0HzwosoJyz
j2LJuULhifdhioc8C+G0qnuibdGqKUTjdl55yGLsO4JOTGSqpIOCsPg3hgiK
oGZ4mToGtGGo4mZ+yhXaKDgKOfEypYvjGUNAxxX2X1bMz0zEFxaDeG22EyOy
/+EQWuaoemYdbfPjsQhWXqGRwZEXAwQ+ogQ5el3+rijdmK3h9lTO9W178OXs
lib7uJQiiktJvyx6DouTSmymPfTwjPavVw4CSC4hLubDBySUGP6rVburl63u
fgENDV5czzsYs554qJ6MFR5QAZgQ1UpjrfZSk3aS/tLWw31i+ZuGigluzkHA
YjivYu+GRpJZORISN+vnT83pMJdiorU27sjhpZlqgQAvty3D92HBtjIfC2lB
LcGyWJY5+RppdlI6nbI4OM7tozjipSGHB33wfqadnDH4aaA81FuOmGQNsPdc
7FjeNWl8kR5XYiZdY5ijzzLUYdVT8uotawhn0jqtbu9dNVwaTlLzG7n4/ajB
DOsTSzt7JPR0pQhhhg63cd8urPGCrcgvs1FZAfHtUhER6sfwi0iNHTzlaHnJ
/jsyWvP43YIhJSIYpE8BwovaEhsYk7xyyb6puyxBqe7x8MdufPNpArDem5G0
LC8p5ZAM/FxuK0wvP8JH74uv3PhAAIRtcHyLbF+skl1XvZwo6Zg6x4ELs7+P
t3qJCkbT4zjtUo/2v91uj4/hjhR8qu0W0JIALo6ll9ABZindII1AnOiw+c00
J+QkOMWTmuJlKKovXCDqLgIijSk4fydpbB3a28IjplADEKBw/9Egn9B2baGP
m5o/1pz9zhzphuCblKexcRmie75U+UOAW55Q3KnGPy9/QWdPKJK31d4VbR7p
84A26GYxtdzULrvwlwQCrMvpRU0Kjq2PnIMEhYL4JBqvxlLpzlw+VmKirKcn
PmgdRuqwnt/gfqUfEstF6v1RfYszLrQC2yjY+h9LShmYNyuEVKDGWoKCfdXh
Io379NDjzCNBzD1AEYWQq1sDXz9uc7wLfG8d3dqwsbq3FYT5Tw07O/RbSLWq
/5xtuv5ZFB+JtlGOJ/+dhVNc7G/8Xlhdk5jm7MQuWB3WKC0LMxWbcF6KAKiC
r9Fn5KzncCtHrou0JuW6yRPUmLNxHYCwr6YAFEpPiqhu3+bumYiWIqtmyUdG
bK7xTOi6RXxTgvKPr9JiZR1AqxPVjg/+V6/TLd6zBBI9Cj6Z7xRWr/+r4//e
hTwvgNiYY+ZGUY21rdtA1TGXG8iqYFScNYbSQuJG+CHi+TFyZe33qO1tSQsz
0WvHqpFCEK0YNfv6OQr7AXHem5KO2RGzKseDtArXjfrRXLovMOa2/54i+5i4
JUw01WXAqtj/pZXg8/7dlj5QmJLXsKWSJsQf/SU0nuV+sN5fl+D8esZg3eID
/wkBHOHDWa/0Ybt1OCdumSZWNWDB8ZFnrih3VMH8iNbGlMhosXjxc0WSr+Qk
x4RJkSrp7svaqpahfyMfaL2es7GpO9ksn2SYAgdYetSqGIfXOMVdjrwrFya0
cjclTi8DRoEyMtcy0ke2qb+KFa9Qg1tJ0AztjkBrChJpgfn5sbkZ52CgVLSu
UHo0C+7H+MHf87GPURrhphbIATAXkT1LhlxWbR+kr9UDgV2bQK5qG2rXAkIo
3BcodrBtU6uEshrmU6yZEZBAlgYeviCC22aZzOO7YwNtAaUnEkli/ElJVXqx
vFgu5DvoBUK+wWR+rcgEHXDdiS0I4FQSSnxWy3VKVoogrka+r56h5KZsSyAC
4i08ObwDF+QliweyTUdhBE4I5kKN7sX1IpajCvZkkSLVuoHg2npdzEZHy+dD
UAaART2njC26mec6X7u9RUpS27wec5VQBq73DPr+rMahvPQT6vgEjqoyQjAc
yw3thNwvqm89tbefjir9Wgf78zppPaGG2OJI8Q6A4/zVsyjuM836NxPrzKcC
rMvV+y0MLB/BXkE7wFeUVo+g3LP8tGoJL19BCErjrdbAXH2CVESbF0yTDjxr
DBKIWG4pmzz5ruBTcFemGj8ztl97EORuj3++LX8HInTFpHnijs62gFcvGoyb
Fu+A0yMC+SiuiSLUWh4oNOx9MAsqjYhI48ts3NQt+s9hRInh4jS6Xdr9M6eu
IDKAEBE+EhWRYQqh3ebmaKvUsw9dLw7I146DOwJwiz+G6YuZxhit++JzTXXF
MVvkXnXcH/d8a7VG2roG0k3K6dKTKBx/FKSm0/3ErzTcSJGDc2LABNP1Vn4l
ecFG9PxFTwOPNuNusTiH2X2EiqjYOqY1lW8BoT4RiA649ho+jbjew6+5n+Oa
dDqBmRWDHX4Ro6djjPGetcJC/02TLJmxP0d7lm664dKwZV8U2Br/2hpIeHXW
7CKnPaWtUPmsBUBl7BJVeVZgDAjir8bdFznz1YNEypSthsW3kCdeo9vHR9o7
tLKDoiCBRgECB1IOIMIPLQNUuKPQBM3Vk4nJ7LoXvhaxrw5kzVeqjqw+fTcR
zeEkGi4uqub3aSoAg9rQdjWCc1xA/vqV3aCePUdIpchEu6Tp1Gp7E10utzRi
eTO3/6sdHTNZA8uMCD+F97qyLlazhjFF/bi3Av8l3c9VH25qPbr8yp4K1/Jl
j40CcWizb5MbWqSKDTcZVQ7SvRc4cgQ2e5YnKEez2JI9rGQqinfUVduGgGjJ
mj4u0SNTGr9NH1rEgA6mr8xx0fGWeQaoYUOhI3X6eqRSj9yDLYo+7wGvT/Hm
Y55iALEVdv6ajW9AFMafpeVxJgcFmV9egBj1LHSoZ/cfybBJOJxmuGDS+YLD
em0vWQy9gGsi8lXXGcTj4BsAWOc++W+E2JQXIdJRg/pXAHCJWMn/vzd03mYT
XmbimSedGJ2xnsOxUKal/4oiQSbWbEH70cum6wKJIjGIF37u5H0Cb5dDuIr6
mI5+8xK/SnCMXp3MlS/sv63Q/vOpG5qhVDqBlv8nrjBZIz32eCaDQ8xFs0T8
QmDVfKFla1AP5+KqQL3NCGjPSv/9UeRj73+HG7IcJ23euaDhWHr9xvYlNNoX
mYzkl1QtLrvU1U9I1NRQKrYZUA/AJtHy0686T0Z4nJ3p9IIOoabPPU27HNA2
gXlfVWI80jBgNs8rVYs70mKvIKoMUQh64wYCN6gto5f9hCn409NmpiM1rh2g
k++hc7+MneoPQ7QMZB68hqUAcK3d28ut3E1P6EpUnMIPx9S93MUCAnB+rA7L
3sGgsJQvl04UPN8XUPuA6rRvFY9Ob79QnkEGkuMoEzLjOmx7s3+3JLbt4oCZ
W5OKWRUJWttlz854slu3MPmgXHmgbkPrCrUcaiQWzgUE9phgzCV1sSEm9jTp
HxLCheHBjtxhQ9lhfWyMBmvzYwQII0mCtEZufk9rOMAn94pfS+KPuihygnTe
1YhbbJAJmgDa2qbGTj9I+ZTS9FssjOHPy/t5ARIjWaAfg6HqPz+gZEUUTaTL
znqHrBcxDyfAhJmH78nQtA2o+j2GN3vVCXfUr3X9xcGXtQvQM9c1fCGm0C/J
WnqLVAUs+/Htr0SH9yRCqXgh8tDzI0gcMmyGvJ6mZ9cVl9i9En+mliWX2XP9
V0kR+r+VCTYsw9OR7DIHN36xKZdfW1vZpeoIvxpDXRVVmProLozlWxu0L2mA
30fUZ1ujuZEQFRIEOYWJxSzh7/1PZB/4N440zAQt7w51jieismk+RiJEAUiO
wPSDMDvnmHxpfHPW+dbUhd2JIRDVll/wToPxeXxU8FGML9EhWUNY3JbwOedO
lT1rMPb9x84dYKxOMlkx/rIGcyyfbDTG+TXL9CEyF2iEZjj5itX3wedHZhjH
eXUgFSxYty5A1/Gq5ipKG7YOMkraJGr8MQjRtZ4SBSWDI1pe7E8Z7LBglO2I
s/33RZ8hXQA1F1fD/t6Qo8iOPtKIQbL8vAqKUktu2fhSEgUfXNwxy0JEjzpu
E5FaMaEUitdmmumJaLN8+DNnjD5EANTnKEH8DhoWQi1SBcZPtXkxe1hdJllV
KOYqO2tR58YfmfRHa662eoN3ujCnFFsaH7/KORHyUvp+v4W5gaWflePztqpK
vZXtZCm5O/YbVDIP/tOBi/1jlu2ekWY6J/YS9NsGELra3Tw57l20FO6L9ckY
xoJVR5MDu5V4TsheifJV2MHBWT933NGdL2jC1EyEIBPeF6XtsDJvmGtwlKvU
0w04lEcYAhaIj/7G6/kgG+jcOB/Ab9K/ezlyA02nXgXM09B6BWMOfCn4PmSK
OMcC9ha0f7yYf8i196ocjlgWu+dMnXoCNlStHWivhqEwntdH2vrs6nI+ieB5
ZXG1fL7rGrIBJwg56YC4MWwfYBIDDZvkxywi+W/ULMLUDjFtBhAS07Gy1b7V
6+gt83pDxk56uNk3j0h0tF2D7HSep44b/ZqNpwv8nD4FaPL2cls/MHqI1PGy
sHNux/N3E+UAb9ZUdtQw40xCu61VGURJBzJS0eRg0KVYmOG1cUR5vVCS6NDj
4srdtSL9lYqYT+ZmVgbYCs8RizWqeYEZT2QFWdsTn2j14vwNdIOETOzFxzSV
xZdYrLFNi2PsCfxJFtTWV98tuEsZmmVf8JMTQdxEJvh/ICtWe/TBtQsuy81p
+tGtjQN7Grvuw8+zyfUuYzqz/HUmbrcMQC6LsIEMZVwBrFu0i803z87OF6Y1
Tohf/JZJa5XzlHLgTIGZTcZ5vU4VZR/XHdHorqVDWZZjcBAAGd74l7xSg5Iv
jS8kT2C+9m6d59MdFlTQMrxldsjPpz+a0OOkzTWuPIEk2UKDOWKbN1mK7a0U
wuGlvzBFYWafsqSzfjpIGT1QQkjhS2ElR9VY2EUvy6V5h5eaxqet5IvTSiqM
0UiMkMHilHgS3LFGeVl2uwudJVYB/z05ReYjn4VXAKmEpjgW3n3Nah3mXAGm
fllC7oB5uNrK15JU8vD7LaxiBTjAeofizZUVG1dF//dkqwYp8xNznW+hpyfo
sPyL6GVMJ0t0m246oSSMfDssxZm7XMPcHNTyljIhyFu9MFgskuU4t5gYD2be
PLkYptfp9HtzayQ6Z4SLYzeT6rsyePaELKZVCfjoQy46t9cOSstBXzkH3RyP
yqDI2+VmY2EchPhggaxU8CSc3R6sbSn7SrXbpNPxkha5EaDOm9cjU2MxtQf2
NGyQF7LAqdLmaUU6xYqTFJlL6Zomp2RPnM8V5zxlvkqRAzM4BwYPFMORTRv6
vx0pjBF+a4heZtR1/KLbTc/evwN4TFBOhMOzMBGjc4g1D5/G3/IVgSXrfLmj
kwEJ49O/3QvpPSyfbVwObD9orzgOoIGsg+lhck/YxA/XDMY2rPhOhHL0QgcC
/MQlWY7uM+ldsWFhBa0gdBVNtbueWd+3eo22U23VjA21gwjZiVpMMi9HpHhG
FZhl4Uv1+/ShrZ3Mm5CPYbAfQHWTaKyAJIgkAYW6D9Pcwj7QAh/3JKqcqb2t
xy27vdYF+h6JguvZ2grV0a9p/J+IIRwL4ogMSkwqzinx06Wb+ciKA+Luqybx
vrnt1VTU1q7JkqC1DX+x3FXyNEp4TWwmDHrFeRPldv4/SBQkaKDis6cqFRKd
M+uGphShLfmwDRcEBQE8zsOeFGyygu7Afy6Ha3BItKo7gl5wFbYUOBN/n6sR
HMGHC7+d6qkszvHv0+kv2eVhgM6iiJi3qClJynVaIht3bMj9LzBvlDlIUe7v
5lK4/jWbH4b3y46WaM2SyAA3X8NhgI85aAT+bl4d69cjpPKmx5vzMGJ1Cvyo
h/AHrmqkJmNKARRSejlFNNbPV9zzb92zn+cJEw42f0r9mHq2OQnDaF8sP2Z5
y624rvCBeKO94WJsyrlBLSBeP+PleobkCi6GME/l/X/sp8tiQurATRqA+CWK
7ouGNgdiazeZirbS/sGk92H64/h5ZB1LdJY4WeQEY9FuY8ruH7DtaYKLvKEI
EtZIHybOYKnjDcQRx8KnrYcsrG1RoVT4meTjeHgVB/ciOfenkfYKpLQysrzg
jvagbLKCw+mm7reiu9ZK1yBpuBtuaRTmxvj+X+KrvFtv44IYepcWxslSHdG+
uY6h79DKqNHRXBL7XG3J2GNZQGW8InzsCqfW3NNQkYARtJnHaxacEuxcg3mc
B4dr7Sen6KjqGNbB2OT8wWPcyhSftAxkvGDhPuixWQ3wUkUt3qiFLJjg8dJ2
W1LUVc1KIbO/EVhhH9Sk0fTOkkXhAhwULbaEjj05yvd3VxdfHfcSQczl+r/E
doauWmKXwZBUUDCLzW4VBAvGL+yERLRaMR0RredtW6xwrYDk4wruJyBBlwZL
vvK4AGSc/OlZyqguIcqemFabDina2nsvkoyCcYQK7VNhmqD1hdTvVvYNtn0w
xBCaQuqL5GzWqvuUz4m9wuVqdBVxfpKO23ECJqCYeS0sBgzrH3H1kbcCV1gj
8JX0kIRznrrX7N1ggzp6xo09MLUpMQsOmwhezc0qICwQ7ghYVr/BPSU9tkvM
nDYtJ1Wm3+qsA6ZevswwRIuUU4Om2F/+AQ4nfAcfDSCSZyaxBLkM3NWcK125
oyXJXAEwK3Wxpl0S39MFTRjzuIKPAn9yXN1APhsvC1ptRN8j657oi00dDDYF
Hro8J2CnOPbJSkKp0eGqY7aKczSPB0NM/1gYqdCtInA6NHrHSOmvMTsVFtPJ
yBqVT3ZV9+/DfAtCIC1NcnCcCZ/cocT7EjpoydXVPffNELb4xbtwHBgQNSKi
mEMvuYbVvNgHczRiYr2pjSw+ei6ipv2OB19dgz2LOjJORN5FhL3vC3SixBfw
mtOJ4oDLvZWWxvtuDxs0tKJEsUElDadwAPbEgBh2odnYP1k6lTosEpWICrjV
hGq4IrvWrIaZSh9a222jO0YWrErgXNAOQeeG+OGpeZ7p0uTr3jrTh01n972r
ffX2vTVyelH9pNxHRdU2xZVgDJz9MTMSruQi+O8LeX+x12pZ0pUQmltxAwP3
qcgmlHqipPgx+ZtVmeMxR1szSTZab7rUsUvzBF271lNkvYaUqfHp8d2hpUtZ
8sAOAD9+wT3+d2N1LsuoL5RQwZ/hqU0H2GQIWU32+unSEQcyxIUxVJnuejei
3cxhvSDCzv8usWF4cM2pOSpPnrR2Wxqgc+AjyWazqd6Jn5XjhjL33n7k3Rwb
uZR3HqPRLTwg4KVWl6IlzmIeIqhJsi6HQ/EayqCYEW0SRz7xvEArmbXLgPg9
lPSP2nE3WTwKwIBtiO3VHX0WFUpr46/UYSSsLmA5uoLNxQSwGtu51aB1ulq6
3Casw4sjdKnYYM/2bKhOBHCLrnBS9Q1Lfx7HHI8WL8dbw2FOuhzdwy7ZlgzN
ab9ehzh4vi99XejaX41hxy/EDWfqmlJgMWU07hl256sIP+A8jPb+/70+7wE0
ovV7IZ8p5nrdX5+r2r0+4uLsL5UqsZM0U2jueDaAbmJmvSPejrDHjIx0MN4x
VbOptzhy9XJx0Rn1oHxVjdmCv7gf59HY5sZpa9u9w2QMeX4Fe0nrQF6fm2MN
sya+kLSb7tqgCdyUtkB4lEFkfo/mOSsifSFzvDxJMGH67jRi9z5XUCoIefco
zbx+jIIRI40oug4vs1Xy9fmsMfT3Yu/EAExIyIUuT8rzoDKskF4gd2/bjpvR
pn+9Hy+t7hd7IYXS52gL4dpmxeGQoRBrj1PSn1vSP07aqbH+PIC3VVw4nkJG
tdeV1/dudWh03Q0H5kwDgDXPvc8RDXQhRisA/WNgkhlEwmgG1YBN7HO8R+nL
iukSqe+hMBnQnD1ikykShAFXLINmf1gu6eWk6H1JmEIVYETzF1KvdENoGwCC
7qqHbgMY9pAZGSjRwslG9YMpzPUF1Ti9YbEsgoi68eUiSlNQ9jDHKJantZT3
n3o13icZWT1DZ96wMz5Lo2gMJ/4SoonXHubViBF/vFx6cc5+kBUpMCtwpdjY
Z87UD8GPd0Di7Rgi8GBXApi4/hiPq7YntlhAJGpYECeqpU9FfsudLgYR7NEp
hG4sTxcoamwrotIKm3Do3vZxotrW2ig9NIOkV3IqsmbnLeVHUzm7i2Pn2AwD
31yniE9JQifhl2b9V/UDZlYeShQY9MCcpehtOpAjvLz9ctVN4BFYoasqvyjS
0GvrGyQEjIMFV/yYDva/t7MP/Da7GLr9Mdg49/i4O76Rp2OGUl8Nsb0b8ijY
WR5RGtW/HZQTD5GLS0/vnGytoBv4pmkEhsljzPq2zUfF38DRybGne0IbrMa8
jx62bN3b2hzjCr0tJNxmIAOhfnVLvCUbPRuUGyLun20t/lY9AH5sq9lJFALY
Su2dt2/5Hj/PQWJbpHnKL5diFxHQSVpPdwudEwlzmsz6QZUIozoKcBiQj7Cv
0bfoswYunf5xl8JGtT4oTeyw2dkw2U7C1mQ0W48s7Z6qu/5ivwKowW7VKCO2
coOLTenxsAGvTqdSpjOJN8wJoZAVnFhO5Xr4URymOUPe9FB+pEJ2K82I+fjh
Meo2N6Tmjpgar6nUR5jB9/15D0MiITGuWj+JQ9pv/hbNE9X5y3ev2KIaXfHv
7T4i/WxGawDhqCK/ohr9AtaduSgTTzQHj99zfYBWDecwEjx9O1b6p6qE1KXW
46zPn89jA4lKEPwmTHQxmugAOnQsAC7OY5LnJWrA35GTiPk0j2g1x/z6DTxo
JCChyEUy7+eBfi+bLQUyeqf1RsN2u0QDO5NtMPbRTW3ylUVGkIIzoda/bSTk
J/rk2WroRsP3pPz3ds1kPRtU1osFYB/yQyd0yGyTZ/qf2SBiJwp9uawaRX8S
Iv1bPXZ2dhnxwgAq1GMv2j6cmymAEyU1+OcbnkYUVBXuLRjYHp458ILdUsrw
gtcSTORnBsnmv3K3NV0RtAhFbQsUKGhlt9uYY2EjnXrypJHpftuzxFiomDr3
miVzPpc2eE1/lhkN8L5bewLS58fHSUelf28AwftxVXVehvoW1eurjr/DKAkf
S5BegH6ClhrMu7Elt8wo9T70MMM9gf6jo3K3BOqZrAuRv88CPshR9NMBy10K
pDOeWrX5iPcpoF9dPvGdWxysJJ0292+E+DUVTGhRw9SSJlvQNwZtYh95uV9V
IUw41wNVAldZHWdMjNeRXMV8Ojz9nEhcrDbk2va3I0Hktzhh8okREvwXta2q
ohrJ0I3UpiVK8O8aG/Q+I9kGqsU1+EfF33qyNMZ9CS+GcPmIj7YPqkhb5hcG
EEGBaMnpcPEDcvFPRqwrsYjB/pGpNo5rkxtHFqIM4bqdgupQjh/erTcVRQYF
8z07Rk4hkRvPNh7XglMFBcBEzK9vyI1Q0VrN1XTjTrJFqiSwneoMUymX6/t7
j0NyztLGCsE43pjOd5dsMWWmXid57kralVNoy4jh1SMfgh2EI1chgFTi9WnR
ptVR0KmDDN4znhW3c16WJ1kjyA4zJsh8/ynDJs/4zraop5K6pzz/F3gJoYFv
LMZrIPckKYksod5OwCLQvKkxZYBN5QtPXi6rS20Dj/Emh+yx2gfKei2FDLLZ
IcbD8MWAd/+h64Yw70DaG41y1VuZizner5JzMpVjOYxOTUXcHORULtwaWsjr
mTsB8JcGN5dpf/YuUwasGh178H0qmkRRGFR0hU2G7l9X8YjXXoaONoJG9pvu
OgA5eqBA4Vad2YQhqjvqweK+IOMZVRpWBbehB1ecWWzgcOtlp+U5B9fRG8G+
mZA0FKNKBq6cet1NenBv4/OcHq3NTAn7TDYkYvXhKI60s5jeEmmyIscMpKus
4+JaHvRxC59u/YJD+lJMx92oLO12N8vrEvAZ9RzWt0m1uZwEjh7AEbCqdGG/
h5AjczNT98qetrISchys/FF9tjhdLm8R+rs5+EMF7EJDKGXKzmOjMNsFbHB0
wt2h2X0znLjBZItpw/S1c6MyCwFv/3EJr0bdA5fI6F2s+HuruX4zy2tNObyf
5pi2Iljt9bBgq5kdz+BH0WC7rimD+1qJtOn69X4eLooFTH2Y2APFIsjMJLQy
AAnKI/FN9d65nTqvsXbRcPKSUGNEw7syHKMu3Wq+kOHae/WVxAvjYd50m5GW
3cSIv/d/UyLvwHgmeEJgrTa24FkuD3T88LE73el6l/zcy/hVr08EcBWyeMi5
ZF6zNzvl0J6BfEwrM876zGYUiT3OzKr0CT2j6RG3MHc5Iacjb3Bl+4HDcN34
K3H/WpH51r+O3O+jkd4vAPDr+WC9b0T3+I7llIrpoKXF8gPX24UNmci3P1rN
DriZ53t0TFqQ2o2GuMzUPv6sNryKyfZro8ZERDGO1R6xx6p3bmvqklLiAwCT
Jxi64yOklh/Ic/085e1/9ZV3yO1YL1PnByLbsK5y4cAiHqgV1Z5UZDGA1k4c
jc775f5wjCytNNopArNG3v24+TKkzFUvJVft83Ny+bNCTGewCmnVhpxkfj2V
13kXS59Nxr3yD79DDs7M/cykd0WcdSpVIdQP1P3KbN7wNOZpM4W0xKDL4Awj
zhWFcbARrP4h8r2J590XKtfsYGW55IXXfiCTkasT9QerMl80PEH2yCy5fr5a
eN16k+dOdm1hPAGsIUc8gLg62/trzK0DuFq2YfHZ+DWJAARRzO684APZN5MQ
qsRNEmGSZPg0rk/0VLIohPTTzBUaM5HHeP/YD3L7pB2528VQAKekl7LWqJmb
GPHIumVYL4Kx2J1necst/jkAfcl9xKW0a/a1g6nvA8+bZRvz9O9rz/AT9x8s
U/Q9sTgTOHuNEh9qiSOf/p1xc++bW/RMlfTAPvKhoh25Cisx1TZNNhjtbY2x
nN8UMHKCAeZlYJ2WeVaWbFx6xnpQZ9XbbhaBim6VY0V3oePlYqec8QLIFMMC
gBjDLevdAkCgD9nSst6IwWoEpdfjeF4Eo5msJAv1SJaoYpmadm5ZBNM0GNGB
cHFgQva4f7foxl7tiQCNNwlL1bQ80YJsn87PZ2QHjGGPZ8bTiKW/BZZtP9p7
aUhl6h6CX7z5MiKae10ZjSVz3hwnKH4e3DDJ+5I7/VvJqD5ZtJczqSqnWRSo
jZDAZWDPRScQzkG0217mgFMPun9bF/xfwlyZZnjBZP6+jRybEAV91xDe1P4B
Rktd0tROwpGUTpfb0l6917mdeu7z8ruT4/za7PpQr0c3DTnf+qaCq7dsalq3
00FVMLsq+sAjBDOCd+9vG/dqAwCo26+Ldd1bis+Ej2OHPihrmj6JZmHuj3ks
/zzHLzBw1BBu16c3IBBN6NXgvt9EhFQ9bOGnDnnuFqPRjeyGZcHNd+1TaCje
SVceoFFkXcJFJ6kXgCcj76+ZPBuJhGbusQVlWsKEkYSSy+tpHgdujXBe3IgX
76H2cHK46NWN6J9T+QPkNSMW/HyD0HJcuTkW2tX310iK/ZAfdhWYQhzEBwYS
lRFW9B/FOvGDyvWNImj5qWyNk23yQr8Co5e25xafrcOCyNc6oOrDJc30coah
EwEuD9KKvjRqSNqW6zocEOmw8Y1YPwVIVJxruya9wK6U+9lxQ05xxw/Ak6g7
2yz4UYDhOCtzJnuDw4jX1CYDGIaK2quQHLI+erCkgKKknAbWt8fRaVZbdK+x
yl7V9mzEc+/fhqLx0n/YstoZr1Sb6b+r9r87o1MH9aqGo5bLSTWoIBLiOzkz
x/ZgeHkHarUe/dNf0Vi0pBraS+BWObAwha/bxH3V+yJ8rDHgw5LM7eceEM+g
SXQblg02/W9aP/LeronxO9h2H6tdLUqydT+yq/jtghYKx+Y7K6YWLP3vsZqw
CsUZ9qCqFDYS8fhyJDrWl8Vaadni3gE6kUoIDaokYD8LGwAp9gjI//dLvHXQ
LEiloDPtlOkQCznMf83VmQAPkClGyTzQWrOAHyYU6E1MVUv/TrhauS4TGwJ1
Zm5Ld0olgFRmYEk3Wa11ydgnKW1MwM3oazHNzIA0FqSU14ke/bhdHAA1lN0x
jzPSYBr/mkC83Ev2Svuhgjuzze7w71sZiBozN+JFz0DwF/dkJP/BXiocAA0B
/syBQeSVRvMRfObaFxKjPwUXysf2EzGxDxAyu/AvB0WwDACYmmoA4dW5X7K8
609QH+4mjJvVm6zPYUBLIek8Enxo73foLyE5QzxTHmZUL1U1QoavC4uj7Kcy
esDvVnI0TsEUw5gnxFDPMv0aLBLwIjp0tuC+J9XBd0pyC5zZfViTUUG/3J65
Bsk9wTqxf6pR0Kbgp1BvVa3fmaBTNsYKMyWNjWGwp1aT952arXUB1ThHyAfR
Benb09vc5RIL5CYuGbwWcIFU3lOJWgU/Zyr7ttjDmInRvvtt3YqnH4Z2lrw6
CiYbZJ3DkYKppUdywTiayWINIvXy9SyIdlsQwBkmwtFa7veyYawgqTTXIcVB
aUaXQdnYl+ZtKlG3yrAOmfw86er4ebOURP9gJkL7rELKNWwwRoymCeXjirDd
lnelJ5aeCC+vs063AO2/Vda9y8pJZRoVJ+bhsofxSO0BPL1eYC8MbqO1I0UO
OWaRZ982sEWuBrDjtmtGMsmZ1ZlpTIYpMJmhvdXyIz3YxFZiXBLi51YcFRk9
EvXel1Bph48qsr5kKtdTy7bn+DoFGKYmext0lqh8oOXtNH80R1kPvyeQ59+A
QkKegy0KtzvuDtPjkX+Y+pVDQaN5vj5lE1ogFvu/q6QMeM4Vj3qz7maQVnta
fDKuSrNHxgZBef11MaI9g0Q8lnjTWTZ0TkUxgSsY6IumVK1ls19j11Nk4liu
/PBwQjLflxG2Dfjj5VMegusRfof7msJ3SLySbhlsEMJ1uOLWRInbBWULbA/x
SGAOp/SNkWfoLIIZCffCcXojw2CFkvPNyAs0d7L50pdzWI2x/j2X17TWgYwN
XPJSivztRPqkuzIy1bAvYWqAL9zJ+572LmvcqTXkvmaKroMu8ICS3UpbtBN7
doj4+RQTQjvk8Alj0Wf9edoNSL1AMuwqkGQidPJfpRJoZjtCKK045NhfMOCE
6g85ABMknC8dAKmWZuY896GdSBKB2IG76mZmEZVW+adYW5jIIlVIdaNwrY0m
CZQCFaF6Wr3YPOhS02m2Qh0Q0e+I9i7HPAZQeu06LUTjpCBB0rJnT0hZ2vFN
3C+xynoTemXkY4jBUmhDxJhRtwNQzH5IL/3BZ8wvMvuoCzh5h590L5eKUX1Q
4/p3m7p/oGwIuaXMntBEJnaL331k9s+Uq8UpW7a5FArUSidMybZt3xMhCx0T
liAH0B2k8uWdeuh2dOavYTvqNHzPOC+MtG3mC3en5TGi9+2/skwYhpM2NPwg
rQ/B7L3RjCBBTFbpnjGdPqvj0mDPPOHIMgSu8mb5jYD+yzPsUwoh7Ll4llVo
JzBTfY8BRHI+FKeRaJ5rP/zx3dznZYJ29jzw4eR1O7ffhNl5EmhLRvIET+rs
B/zBAStkVZXySjzO4vrj1X8lI3NLfr40XxosVqEFXen98pKxG5fwF+ewJF2k
1OcEQL22TSObcsF7dglEs//M6wNYRjXkDmKSulcvcSDbq6QB0mguF9RQgqWo
3dQq0S5XTj+1hD6fQRfRz+gWqR2VLEovnPq4EOSmf1gblS7VRZ/vT5G71mhi
hpDlmZpnwTVSkZ08Y1Xcsb1rewWDy83oCRuoqzDx4lHFvTFeoy4Fu0kmkWqx
qJ3rVbgXPLqn5Bsj7oiRUVLRIuPoE4F4faYwKvxojFlo63/GRNZ1cYuAHuT2
4lFB7weCZ1Wdxl+3HRA0hNohOJMJaroPWJGSY5ZER+sGAiBJhJ3ygFcjYSVg
L3FdCuy1TsZM4wlqkS+5FrVhyOB+LVMwSX+ZvLuJmERUIwLHteaV498DvXnx
k4ygFTUNPdis4mJx7f6nmZbAvl1yBf9+Aa9LIjzTDO76yRPi3+CsMaHlALtH
naxxRQEkGkHdczh7FJsMOAA6ba3X1A1M8jQdUm3V4BVKIVZcV35FJ4eFS0Fu
thzkdcDp9zQl+ZdNXACWaYidCoaW5x3cTAW1TRpx7h4/qKmVsEu4+4KA2Ivc
ZhqttipFiBOtDMd3+9jmFIelkAFI2B8liQkUQzZmxz55q9Z2UFg86BCMgqbO
poPWuIfcLaBL1lCE4eE1c/n76AZSKyy3YZ+kIA+H/uut4QkO06XNDfVgsApR
xLwwsexiKHCAnIS4woIS8GjG5soGGMVMALs5+XdLpban9nFAvB3ys/Jvoncv
/X1ua+Hn5TOpYt3gUsTwSeBOByt6EbFa/q/gpcmNnYVJu/E915FBT9qCnrrG
VtHXi32NuQHuKJwfkXNsNUqVVKdi9vrRn7B5+DFXoJfXfr8mJwu/a3tAyK/P
8HYJTgP7mgCebPDE8a7lMv2hver3eAYLatp7OYYeZsWWw62qIB42dQca14s9
26pN2ClW0XuefjYV0s6KeujUg7MZIdL0GOLHXkSZ2cs9faXil0Fp+EmCArl+
h5CT9zMBcRzrD+FDqtTnhkBbKiaozksDT0XHsV/0rQm2n+5ROToRTuDVPZv3
PJNQD3lOP57ojAklXRQWlv7uvOoWn3tqEmDuLWE1bQhfmi7Ap15bArFMsRu6
SQjJ7Ms1eusEv0GtE0Vf/TEz4bADmrLeFI2t8aOvhg5yQl1G9ygw019OKz4a
dEdnE7XX5ddcl+ybnHgci6CkyXKwGCKtON51GGLKISFww3lsNdd+oLA3Nq0f
aY8l3CS09bj36J2HOUu9yLx/w+WEgxUj23M2LyK8omlWgB0OdcdphhkL+Vgc
P0IKqUUnqhLoZyq24uZwi/Yy23sxyjwOMlEwXLEWSLLIlhmsMtTKwIJVLggx
+9sxmwbQnmYbD6OrhysX+AvbT4wG9BvJayD7c8h+9W6DtJJRvHoM5fjCRcjd
ULGS6YN6JtJhRoOIW81SE+A3W/zgs3ImfzZtTu8V7STheGARjfEfWmY/MUeM
2l7LddpWfQXsJUMcysmIjA8IQz4owTpcdRuWsyELfJOfc9V3mlbYc3ppsC1F
8v9jBb/Uoa7+jvB/L46bcuX0CzxKdWYsXz85OsqORBy72DU3djUXz9ge8yQX
fwR+lgQK36LY5/6ruB/olx8f5K1NFmniTcH41wQP6uFrYiqH5OgfH8XBS7DC
oOYuY44i7zcJ7hRauO6PWRgRIan+5JcS9wg7ifo4GOlirMihMyW8MBi95Q/f
Q03+gpcX1NufZRQ7H68XUzvavLdjupahJ7/QK6AB5CkmOuoTlbcBrsDaEZCL
gRF1/kAeHAF9ULg/aZsy97rdPWa9XaZKB1HJpJp7//CoQ3b+Ry3xeLSAkhLX
sD+3OeK34AAFj46nFp3Eq265n4xWj7MzZ3VhtDJ0GTiPg6/tDbMqHWUsQaxE
MaF5cFQXGS7j6lbmru8vw/VXMeoOtsB0NE+z7eQBIKHWASrErAN2664Q8+n4
SzV7QOYf3PI4fmEtq7A1HxfgVh7Rnf4aScBSY8AEYbQdDHuUWg4Lnko55Ntc
wj42aOvaijB8nOQoK/fi+Uzkxqq76h2C0zf7XDRu5ZlwbkkirVmRO87aQfSa
Ydp1F7Fzdla+jVvjHit25lKTKFohevzmdpw4Ggn0Y/ikJPLxNAS+czKjR50d
AVwBDgKvgtndHThlZ2smpIn7q/9T3M5wFsVtynt3+7lanfHlKHspyvhCbnZ/
07F45VGCiWTUB9SqZ0Y7NGFXPKspPaUV7cHGBRysmrOgy7tR+9FFG9792zDS
gTNiwHKX3rWPgeAy74u9Z+sNuOEV3DyzGY0B0cEONUoJHOzGuQeXcNnlDt0y
iYZG8Fkad9zTlEJN4nRIC5VgQiZcE3Hoe8Ie2W7ZbJ4+Me3HhVckSd7OxQuI
ftfiCKjYoD6Y7/InEtGweGV5GGU9sk0x+DXf0k0aPabmvAsLcv1gmEed8mzM
Ff2oSFaSLJ/0B09NYhGJSkPPM+MuvMghkfHSJcCA9mFHJvIJNU/XGXf5hwXT
pLi9yCn7AoxUAuZgb74Lc90gHgcQhgVHS8ph5A4whbLgmTu54meirt7IgF2/
kc7u+aXuIccJ7OSm9KKeVN+8PwEEGoXY9Q/PvcMjmuQGOQCCkYc4aeUemnch
fMcOF1Q3QAWXAUX9ZwmgbWguzDB3xyXlBg0rWvmp447iGAVxqyhtRmfmmHD7
MQiJ7WNu58fPRLoa5rhhNywlfZ9pD9dayu8HTfHEFO4aX5jNqdToNLFX+14Y
0y1F5u83Dpllyvoc/ili1Dhv2ESUXCohD0rsA+VHdcQqv2PcUvUvKxSMCF3s
9Xixtrc1cJcmY7IDDhHu3zF7qrW1ACm4HFYxzGOqhiXExwh39Mu4V9c3jKZ5
Iae0IFMaVa6Tsx0M2ACCiu6yWlAg6gECmXsxdgDZJ9i6ds3YCXlf9bL3q49p
Xl1aaP2RhEISvLfdl41TE41bvdS8/xwVVzCZ7SxITTBn2xPgfidW3WKvJ0po
WP7RelIzA62cu6Lwk0AwUO0xNaca5g494gIEbkC7cA5lc6KCeu5DLdClTSTD
nPq0INLdMChgvCwDUN6AekmbS9ALpngWR/PCRc+FP5jbzCL/FV+GF7sQX3eA
Jae/bqImCqtfR2Z/sdPwHYa7p9Y0kQfWqkzPDxLxLcOY9qqmAeko5A7LPGcV
7MoNERd0gJtB2KQM0FRR12bMz8w+RAquCnw0aka89E6YFRcObPhgx7XYEDwa
kCdEzQvDP8uWgRSNNUzT+zUgOwFmXyI3T1NLqIs7Er6GZivuqTWebB40CxH6
XgS8E/Q1KByEv8rv11hDN5ff8cDcCCPWJBoEio93nitJ61jCGhTPuQcS60lh
RHxFzTp609/5cQVuSSazSI5/2M/3sxlYmyw7vJhwX3aIz3SJOAftme3xwTFj
fn2A3Iz67b9sIC2enTeo6j/VMTvTU7Vynhgc8ZCS2K61u5YxU6Xr63Pp4s9u
0v0PHq8bLTAyOwr0RFDQbskNJpKD8uoxVBNogq5C2CpU5eK9DECKNAbHX7J1
wxW2wltvEN6pWjptPEkNInQmgTDDamHzJhcgSEjiaNqM/67dag0FAowu4jTd
zDE9Z68jW0wE2hE4wYKuru+oYqYvAJ1dUlRssJ6pzYp9tfqvjgU9gZVIJ7Nq
w5qYY96zZgqLpgPQpN3o+rhZtHch53+QJh/77tU9/ki9zPkt0oq+wmFCIwC7
VEE5uoTyjuTIQz3fIZNZk8SuP3cqEdN/ifl4p+GNTuAUWwW7rOG2Bea2h2T/
HCFqkXOnIrffst7DkqsP5iEcUmOiHPpESF30RcozF9fIuHYBWSUqj03s0NgV
dU9HlJaxFJyxkEtj9rrd9AxgD/IZD0Y9LlFicQVcy80SH4GNpG5TOqyN9WUi
IQf7Yn88l0bLH9cW+H5h3GjivOnVVUu8r+tT0ZTycisWdUKt56BifDMK54RU
s0HHgOjXO+vcTirYnbhdtasUuDqGcwTFRMhXAQ2AvmmyloB7zdrhw41H/cdm
JpCq6Mhg//1VXYhh1i5nKLAsvMVaEGVK6gFZzTQV0RfqZpzfFWtTe4xXcXo1
gX8zejK2bE3F4Px3xef34QE8Td/j69mEELfrhPDMMCwkomKAEj5gLbvR2vZP
giAh2497xiXvoWc9QZkRyjj4WGnnsA/SHCzNscg/dv+vmFGlWJp+dQ+fwyaj
6AiRsqCv6vPtrIOBe+smX2G+FrEFBS6AzL5XeW6ggXO/ELz8QNTPNotmK6O1
C4rAM7qOea/JVOsA1rg1xeMAzUQpSorA0NXAU0jBy0MNeke/yvIVO7BhnkyQ
siktH35ZwmUoT3QFKK5GnMwGy8p1YWiCE3bKWbIptvrrHM2Njq2j+l4ROZVn
eO1ySJw8eJTHoYCtBPHfOgQaMq6i6tLOP2owLNQExwJQMTOWcI0NOrg5xTYD
7fCePC78Y50EXbNDDAXDOTXRPiqLikAB7KQgCx0kRe8fXD3e+0b+y9Jh9Fd2
5n1Cuh18dxsObthMTjHd50MPVcDTNV8WUHtY4NHTLnUKQZ1fKkMrsKaUrlrt
eacwXLAH9zPz1qKyXmz0mKIGoIj2XdZ7xegFYD+WwXjdtr8d+3E4ljMeW6wd
+iPJOhw5f4sNqX/g5AvKmuj+Jti10dfiBGokyQIV6t74I5d16d0DQrCSmD7F
WrT3MT8ikX7z4uUkmo4+Ycqs4gDW+Fhf326ftZqwyY9QEBxi1QcGz2Ym4GlG
LwoS2WikA4b4La8SB1wGhviWOhpqYbtklgfluNLqmlN4GxrPfE8hxc2NssDK
7zfQKWxB8ya14SIXlSf4M/mOneBb0soLDgekSrYmAK6JviY45/lpZ9qWBC3p
NHSyJKjAQ6eXrnTnXnIEnaRxSwb10jC3JYn6umh6k8BiJ8WnUyLsZctPMHTz
6os05VTkxL1yhZrWDON1isSQtBF2tZw6pFzHr5ZQDxi5TFU1oNGVdFLh7u+q
nyZ8B07BhxI6+59B0m1sFH54mBWDUo/r3bUT7aOFMZKa3GP+pTM6v81n2hK3
pRcItbTRxLDi/sFIWJ+E+BaiALS/VjxoCSBiZeQjYB4AiSEyH1tbNTC8gHTA
Gta+XuXKeS1i9D313Z7EdMYT6UVh6rg1MhmNlj4D/PL+GjskkAoafT5k0vEn
D99PWhOKC271y+Vw9L35M9/kGh2uhPIcr2dU2AAwpOLuXCzebkwE0u/z9SYb
W4H+jyoiIjFwqnxpZtL19OFdXHJJNFoyHy7hLtGAIbnrx3GIOLH83UV+pmiF
GWKPkYCehHJ35QIBBSqv0KmZ57fIYt/yAtfv5eyrDK5xFY4OI1gEMwgpbuO7
3Gkphx9PLwIE63gRIKB1igr+WyyyOn0D9LUmuYoYwKQBOgnAmUiCTcrlirib
DYkcFiTUhnmVswN0Wfrq+MlkfU8q6O52iB8d3xRxaah8bmKpddmCv9uhGRBW
9AMYHSXUN+CYlYrOVZu9zUT4JdtAM59bc/FOspTQVU/lYtuw6WSeL73UpI7c
9c8gGPsyL8PsZKeGg4bU3aqZegazlixqRHpqrpT+ChUlJ5cjh27Mj3gAtAM6
VMwXprv7EYHpLoPXKH1bcDVwYWrjsnq7PTl/AGmxp8AJkq5X3pDQCBCqv1wu
Fqxy/2iGCPBeMza/BLbcWk+YBlv+0sgJFVy2ZeWkV9GM1+2eVDG1AmbYtiyO
dws4iEKHfN138c5UxRx3H31x3Pvp5LByQD29GI9Y8GdmUoRLJsDJDD74o2+w
8XdriZDrT3Gwm6GOnRhERsSVMFImQ/cv8z4z1ZF7vqDcEy2ovxmYweyUz2lL
pVjmaORX2S2IRVosC2m7jYdVv5le3p/VtsPkUv5Afgv2Z3q7UFIHMnbmyGZH
uR9zYGM+Hau/xj/TED6QLAOeXkNqtAyAQQ7ljW3RhXg3TVVOJSvBYB+ZI7t0
qlNXB63g80GkobVPVdFun4QLUoaFPugS9+7vR2+el2z3GQkOSSEYK8vVaYog
SvVDSqHKEPkqnl++YoX1GjZzp9yWmap0i5HI4FgAP5lrWhx7k+CoUiQ0fVs3
hmbT6QpficeSashDPYj5wJr5cUdK2GlHFrLUvPCbPtPjAC9sqvEOPB8/0kCt
/wqVcpfOc28lHkJ67YF/sJNuTkon81J4v3aUQ+92tv9cnwEA1QLthZcNJJla
yprf6V/Sy42JQRiFi2M1W4i6wayizz+bt6m7XDpsaDq2ZD0fdhe6t+bqv5Yl
R5UnF7y+GOAfYPuLbTgm/QolmYIJ2NBEDnxB6pyogYHdfjbSsiNce6dl/vR8
TnY6nOK28jOfwyUs9RAeSRe9LEeqI2qGHtFtTVDv4CXZRbwOB7y2BoRQ8wcx
3mEA5jAbsBKoMWc0cf5+ru9jGYdyOnFzqHU3qNqEqG8C967yn+es3raBvY0Q
LkAGXVPtNcYFCQaZVg+QfTg8FBIOlZ4wnrUbbox7gOrH6pXt6vwIJu0B6BtX
sEFn20kzRims/3wa4JhWesG/Tp4RWE2opv77wYvHVFmfwnAjFR64+cpdLutY
wrbDdRTZAQPJg5eq0mAj7V1YXKiDisWGd+kMYXNzw0563JbWFio+T/ZzCG0O
Vu4u50MNSshOThk8mW6OWi/mdtJjVpv59oHijHjVTBqPaa344fb8DR//adS8
ZqS6BpS6vlNpU6t/+GwyUe6HsidLIkccnHFZMOyiMI/EYsx8GewS7qxZNhTu
oYLYOo83wsrII07rdXBfa0fujRUmWYpiOFq+lPQQKoeXho2ccaDV1luTDy5e
9mhDip7d7Oe/RlPfYndzEQVmoBuFkvgqzdi2jVaSD+HD44NQqwPhIC22QRv2
LU03rJw57aRvmlpw/2uKvXkyb8GSLWCmvCbwzVM6NHzaqCXDJwnwgUhfGevT
FPFAhIPzzD1e92OJ0BY8njwJ2Jt8A4vXDxnzpNJErzFQXGhNaZhq6XXYpFma
mK5rkbqzTLaRHW/ZOCOpQUBnkOlTOmElAQndrhDaBe+ZM4E7rrWlNugLy9um
Aw35Iebz7+CMBHwzs18PD8EwqetwJOS2UPlY2c7QumiYH0RFXsP/Bgh4ele9
mOSI6prlSvkCoJmXiBM9ZCsgyt41ovESMnmWBW2uyJ/NXZUXY2GGcHOvXAiC
MImUjFn76vBjqLXhY+6dV+XchNN6kxclsJVJLoFzqzOHfMhF5bBEoUE97GDO
Z8phep9EtFWa7iRVf8lAp60Rjt64cO6JA8Q1/ZjfmrwGFqC5dyk+PFgXQKtF
knf6FEVD4cKWY9V7lh5OXaCY1CoBje1MtrYBY1SOBNoc3wnC3N5n4RwUdNvW
1bbDfZ7+x7MwvdTWh1I/6OvCErCCKPgXpN0805QHWhT/B1vNRrK16hy9ykst
NcDqMB2Y3kdwgDV83d7t3VqpUCX8KAZvvgfEx8oOafUooV5n2N3uW4canSNa
KYHHV3Z0QAJCRHqwtJHaSg3Pc0+lpNnPOC4b6M38D/oGdnfZE8uvB1lVGP+I
Js83Z8RIKLPhQHFzdXIUXtq0Go6VsqBradsjtJDYG7bGZ1+kDjHlDLLLEUUD
KZYQxb4hm3kz3ojCyPzZWScgJnPoT/MEFQXsPdFWiMYux6v6NQ/cBIis9krO
5UmWl18XBlVynTtYVCe3auR5KJo9Se8dq0eXEJ92OR+zaifXttqxxLbNc8lq
icWaQP932Wybjfb6X4O6cPdWlT9v1U8mU8QKA1QvGUchneqXe9tEaIOKF8vD
g47oKduO1VRfMJdLghXb1oYtTgUTRQCVMp5+KqCtcNRaZ8Bw7GVYHt4hyWcQ
miiERKFyHPReUPumIkGFoGqKma3CPPIWOKFlF1HUK/z+5utzI7qV/oVN3T1c
FVb/H+69zlHfFWbxWnrZMh4g5DH4RMODnB4p/wTDMMJ0w8xCTYYjHbVjWjio
GEQVRu2DOb3y0zdW8Wi1kF8EdMfQOCICHZ3ypdyW/q0i4Rznv0wRlCYmCFjW
cH5KUzT/Y7uNfne5z9heDyVVhhXe9QZ87R02qbL3E46YXUOCrCuT6L8oOL99
FA2CIXCBOZ8X1x5Q55bhGa5U0yrVKk7x4Pd3ba8VDiU5KdgETUgwlAzkQBQt
11h7eW8ddySds1V/oeWghE5+MCvUvao01xNYoCl52TxmChpTda0Pkpp+bVJh
DWhxEaBvS4ngeOYVybzvaUNygZQ2KhjTiw8/fhd7TDi8RedlAa8Oys5E+kLJ
qLtCH8CLnuOlV8TjXimtrznxEXLE50d5M6bXEE2WSRTaOln39B0W//5YfK3w
rX2jcFou65TX5CF1Hbgn68qkfaLf8L+4/DemAZagDQndRWcB37+D1u4ZdnJY
8y2XJc1pxIyuKSWdrBMZAm/fL3Rtp7ydA0e1QRFIfHKobkTm7v2h4rkvi3EJ
5+Uni4FaR+o2COuBS8Wa3LFsZZvvx7OxnJm26Pi3YzSuoQVv+6g9wQ+NAgl4
vU1JUN9PO2N3wzhveYBrtOAMVBGCU6WoSrkJoO50syKu1TxL5czODgf1P0y/
U3467vlk9r+tlDvVThBRSPGwERndoTKs6dcJoek1tY68s7PTEeIXBmWYoKTu
VUw+DsDaAMJzLEdoNkIv3Sx0zS9JznOdXzxHsurCaBkKS6NPHfjfh3W0Vtix
hXMX0Y0bnsUoIhmQHFAA0c5BbxMq1X4QqmyBOcoAl347jH8BvQb2G+0Q26m9
96Zc7wAusJnQ8JRwLNyM3TzTWjGEWV33MuFi9eO5bB7WbLmnRxSoupiWES8f
oqGO4dMsTFCLP2SDXDi4fx5qG60KCQYSI3V2NhYD8WpJvmJigNjy+1y/3LCy
brhc+ZxKk7vbQAYwmBVRJW81GTNMD0X5/54Qilz4nKfxVv3gp+vCcGCAf9EO
Dn7RzUy8OgqJuR5Ya3Ewm8oLAOO+D0rBuyu4TSH5mgd2vBXgPt/WxTJhdcn6
YJyz3ETOtEAKHUTYUG938ZdXunyYCoHg6gEMBbuioRPRtmY5HZaA6l3G3911
NnsYhrcqTz+q8zdbHaE+6Yg8Rm4ermRCs/RglLRPhbSdRJgpQlnZvEBmty05
cjPlTnS+Dx/Ivu1HtC2zGeBngTNWSkff+0GgM7DqB+BNXUvY6I09IFGYtAj8
BF0SlJG90zR8HU+wEfgteLFSWdRNwQyip3LIzbq99eW3ol+DHKe9jjfUOh6A
1qhs5WuDH6qJxe2xFkhDfReoQkhqTq92jyJp58hMq9PzyE8Z8gOwWl0PrpA8
CcJNGQ3J4XrCJJGxWIFdHWP29N42ZqKrrHwFRvhjaqEoCKIkSzka4NJRHifs
1q0EtKzSkpA6OyUntpNvRspxJ8iogf+SfTSM59cViIVJNPKaGeYeKHWTtfeq
iS2M0wwcLUx2vYM4l380P7BRA8j9RrqtZJ30Qrvjytx258Q52Y2CV5sHmGHB
F0A69YgWB3P3Lsz7mWJ0gFHTLEz18X5HgujOQVl8uAvF/T4GyDVa3dkZw0pA
3/3RLmR0bb2Y6CABX3TIjWYDPNK2BX/tsN6hJ+ghUyxZgZfevoLM+bpQEJmI
iEZfu/SsIxobDEK4hlMPDZbLHBzOXW1ff+kO4f6yNACdL0igvfJxCDJTirmS
1hzX1qZd1s6fLC5qZZCvKbzL05vgbKpTwuskT6XpKlcEOtP5B0MPsvew4tmc
TWn3vOB0fe0930GenmRb3xlDb9w8t3fnpmd+jPgPUOqCOmvhHtFsQrZnDBvY
RLYhNqg6k8JF9b5kv86yNcaK0V1goXUUC+GvrEwkwlvSxkc5+OjoMejEMjC8
cdPKlpYhJ8Ggol5d1bEnD6aRFFdvai/ogPQ1aeRwwYvNe02LlsnrWSky2Lfv
27AV1Vt9/b2MuoCYSFa13QKPcFzvW//WRJ9eJSDpljAf9Ip0S7PoZDrXl28D
iC4HZ58Zxea4ZlwcDBujB8rP9Wvoo6CTZ82lnjF9C3ZwgdO9Addjg0dL+m2f
q6JxGMLjp+9XOaDEB2YNHLjHYdqbigrir+0YbXL1TT8/zHOWlWKf1AYz2uL1
9ydu1hDkorS3AxkACzASjwNzM7yXNEUoK61qtzh16qB0FhNF5ogyOlv5jFgw
BVzRueilrvjXZiv/bZMGj+6glqpyeqaedksZuMY1VNb23mXVaA7sXNfPJ9py
W3+c891o8yPuvUnslaeot0XsQwxeVxUmtKkFaY9mnEghwryvyaGXyNyRJQUl
C4pyQV7/VN6zel61XWSqlUrF1cFOmatyOeAid2DwuRRgQ7VQMevl1VPXjKjg
OUDNznrHDIFFMKQc3c9Bm6sMGvh5f7tksyie/cFCShPSHdT9dnuhtE3WCGuo
i5Wos2Xzmu3e3mxxzbrh1gVK4R32d9+gRryYMsrhNEaw2MugDOeHtN774nqD
5V+jsG8PmXAZ6cVkfd4oVkHweiWn0yoNYSC/GbJEp3PQY93Vf5k6U+wSe9XP
O6cqllJokRx0K8X/GwL+MIiZLrkC+QixCxq3VDzWqutY77WXscMNIqUZFdKk
d3nvWi8gBK1qxtPZLS582AbMfKU1BJRQ0vn2TI0ssYfiTDEducK3yzvKHfNS
mVDi1IzQdbaaBgTOVVWRG5rLBF8/NaSq7PkdPBKkKTsS862qDh918a6FO0kk
9D/cK9uKgZ5qMQLcAtKYpECBiuilN7TRBpX9bKLG3YRwNZD+zmMFFQARlEha
4jf319+H3OHoF6jGhrOw7W+IcBz3xHmnVa6T5C6hjdyFTx2gpeEgHh0IKwnL
1HWrvjhmHeKi0l4rQDe6PuNId3xQ+iGXcTosNaGDhjWgnw7/l/hozjQz7Kmi
m6PptMBqZE143HCvNRfBqBgmtdPZhblDU4s0e4G/7JnANyRhnSZJ/9WcbbEy
qIJpKRzqlJUoY3GuuvUOhRi1g5z7f57+A31cN/0pnbKWnwpvnKJzLkmNBOa/
oqtrGH058KQ8wVfpNRNa/CEtgeyuzWiAR4eH80Cn+JXerAqHtgAvov/OTbCp
3ZYpmBs/N3hR+RzbvQZXo6KkcktlC0nX2bel2q89yEal34A5qiZzeMAo4yO6
0Z2/mo4HpTc2qseW3hQOX+C0Jp7R+MYuwL7rGuyUy8Ism7Mp5BHVRzxvy6jB
DaEnoE2V86oi8kc/1xGJijCi3zqg5TgCNg6xuVBDLfIBUwi/MmnkOeISmMSt
9IRzZD1PyxTjizeqLDO3DvXgYdoSDf1ID+okdv7X64S0MKli1/zBS1Ehq7F2
EbxIR8b5JpxzEO9orJuJL43ZgpGNTo3Ecww97kLe/lRO2LvWRmXtAlcYoB59
QjI/ydOmRNySKEdfl4hhyv3yQhX9xUZPz4S8YVttSJyXmp0cZUadIoq1GR86
Lr+3wTg5pCgYKptiXRo1T+FHR3HlClKnPc6IMiGG3tgWVlh8/LlvBKcULS+r
M3qkqGjsndU3p9iY9pxILa5gMldrOhN/m+ZX6KKgdzzftmPEspPVWXn7YBSj
LVst0rHpl0CEkvhXpvwKVuXu8lji7WJwxFujstJcdOaii7ZV+vKj8u8GwUVF
U29J0xuCNwIG2ATynXD9Y/yjWyWqNT0OYem4soYF5VIXSBbwCkyDE13nKz7F
do2HoNREFE5HrQA9VE/X96eYBBaXhzsY+mweFrzbwdJC9028snIbcxTvT9Lf
oNc3GyCCxo1jBRpvJvU1X1gg2LKmUVu5WjV6RXaK1aA1ZJ/7h+V9FvVXFlks
3VNdb7YLA+5uSJRq5mQp13Xg1meWZv2W83J5+A9/4jatthuyNxpPsAIHi2B3
w6wwYqdPb2QLOTRldzgdr99wApKBomrBLKHq+cLB6KJPe+aLrfNwGB9jk+fN
bEA99CknRuZmQTHqfPbY6D0r3KvSo6Ckbkz/zVAaT1o/JhVZQQAzxAsxCx++
Qe2FYhen3RcT3qHoTl8XzhvfbHIR7N7YUfGDptQl038G5U+Y8NOMl7LPWzXg
FZ4IiDnAysx+kAl8JSo+uJ/zn/MRdE5iXy+Ga3lK+1qb0tsziqYjmaHSQWxQ
pTrCZvO8QhUJi8PYHaWoZthK3oRkWYWoq7ZTL1x4Zqz1dnZCnOYjrAdWDq+1
cKwEF3C2P+URu2fAZ8cK3qpjTBI8DV1hqJCQayUMm3TDmIkTzeFX++4nmp2H
vpVWDgJKB2AZYH3uXQFJiC3JDCWnj3tXTz3Q9MGQ298BTpUO9NXtTBoK7PT2
mEW0u+zMteSwnlY8nQcU74rpD80ExLBxKa2in8D1vVIPREumzGAY/95c6wzH
IhUUb5uSDuLzmVkyPo8E2gsiF+/WIskxX93F90MrGrtchqnf//BaqAoRjNKm
FhCRNu3QZTWFHawpvLjZA2ta0j8Q4+U4QFND7vneehpD51x9sxgYa+uw3FgY
k6Hs4VDQ8YExeXKgV0MuVq9Nl2vHjlyqdn97QEKc0seFQBQgE4sxwhOwdXmg
T6JmwHt2j962Qxneq3zra3W3Hz/BfcL63hXyJQKyG7qu/IPWTD2SGzrgw4sg
nLcwxDI/z/cw1n3sGJJb3ILP2kJTQJH9REiXqPSF2QkVHHAeiuDl8JWWNxQp
3XxK365rBnwjuAYO2UMV2kIeJ8iz1Dp2Ddgqexnoz+YDkOCNx9CpBDja9xOc
iPj9u39EK9iVYrfQpWL9ihWy2Gn162qSdIIM8Joy3lI2NQ3XPoDC6Fu0QDlE
0eWl2F8qZGcatOVPq17wSdpTySfVz4aFb9tj9ohe8gDgkvoNNEuPA7tSoNrb
BxJydlMlaMs/gNmPLdpJVVTpWngl+4hAu2Yl5SuifR0SKrB1dlBh3+xVuOgJ
PHUYtlHcaH8oCPzfHkOFjy5i9MdXoU84tIJUu+wEeOgeSGuptSRs1FInaQa7
uMhzNgnKtUnvWWtVlf6ja1EllVmPMBBI0eVYQjecTxyQMtB4nozAsrwd2B6Q
FRG9yt2jpYPOm2WsBBXsDBoPPfDup73ftJIjUhRkW/Nit9diE78WY20UDKlQ
RPPiil5pW6SFT/6hCHfZcwG7yJjWFGvsyZ0W68NxET7JBsUUQkIZU7TNNhwh
B5b5DcHohW2k0XggVkqWNaYdoysA3RJjWyntTNQ50LfmEKkk4RF7/lw7dq5B
5jJn4j10g7OZEjBYLYfghOLsg1gd84L3j3I7vWmUQI5vHXT9mAaq8hPSiu1Y
doV1RqCaJuJz2zq6UlDcywdlNSFtMeI+Ux+SBXzkKEQSJD+O2qsO57MrK24n
4F6xurtEdXPE5os6jtW3Y+akkaCNhKNs433YB48AmTbUKzLBULaCGvr56E7O
43pSDm38pjGwbuJ+XjjGaU+Nrt6mzbW9FSbc/8i3V1I7vr/a8QMcrz85TPpx
nTjmFTjOWMYDYfjhJJ8xZ7DZ/sCTY38NMOv2ep9KdthejubgppFPOCk0OJk8
wqpdkej5RhWolV3BtZsKMwML3FH7k7WotaJNnZBx4EAcjsSg3Fk3qeE3IAMB
2duvhor37y40h6nOUlEM9m8qdsDXzMXD4iA9bXAGutYQXA52D/64Wwnvtn4c
i/KLSQrVrYezpDUNUGHjDkhKXmDkhotg/qbRTrXvJp2/kQm9eiVy4dUpOlDw
iEyXtfXIUngZsAXnrVLzi1tliBy72AtdlYpIDAWEp10Xe362Y35pzwyPiSUb
WsIVg6DY1pnJjt7LNrSFcbYoVxDG3nSNoqev8oUFBPEM8J10i+Zm4b0Cz2Gu
jpVqqxYpX6w876En3n+0Q67lEBth0vZoo6vZ3h+uOr3XYuEgjbQbZ6y7sV8t
RrwksJninjLvq27Ch28eYFJtSrB+VGrvuNbl8pr/AfYfIAnL7oFNOCXSvZmR
4qyHceYcY7VlPyshs2ZVwhhbXi+AqTNzcj4GdSwG8ELfABURbAl5HeGPPqT/
whcwYfOel0lODAQvhOEfA2rAV0akRqQvhIGCdRpTajtDhw0St4YRJX4jQelT
3QvLVVfQMnUpQsyS/VtkYYBA+ofAu53pDZBkWNzssODRF91zToEhnXLq8Exj
wKSK65DawIua+uGoqLThlL7qMwv10LHWLVKHbF5tTeTp7dltXKxJ3zAppFrg
3t7SHRhIozLippzheI90tMfWrT5ZsA9HfvVgW2MpZ6/0bVOvDiw3kc0+8KMm
oejDZ0RZ1utaksmBT6p6i3jYKEx5mjdMmuxMq4iZsmNuXfrvSwW9b2Y6gIx3
brYCilSaV7w65we5Qp5SjnohsjyEMT7812GViYhWgHuw55hFdRtrv8Bq/Xkq
CfhvbqcyENtHtKhPoSn3ltsr2P8nQ9HAXRDJ6eeWGD5KHiFZvnBf2iQn3dlM
k1zkiJPBDuf7Cptw8MLOoSzHskCo07r/f4affQ2jj4sTpjpDYIIB5Wo2ZU2O
vg6yCcLE5sXNhhGgpjPedemfThRdVB362WPct2ZEDcZ4AaneQPnlZERZHoJx
VzdyeO7gNrPFNThEkWDpQqya1PiFdKNb3dT0A2Zs1inwZkRzOAm/WSvPgGYg
LJutCiTrPrXRjKXIS6Bel0/Cuctt7a4W7rSZZRm1DkUgXhJ/vFegInvu5qaB
7oBr3ohxznwdR1waP8rozPGVU8mKi2brgefZcsF1bWgmnIoiPdpb+n89ET67
LV0kzqxbYnbNM6Z3XmkE5KJs15GVWysEaBYqZSDW2gedEBumS0F9BmzS5h+F
D3SZsclz3+FJFrCchx6XeSqr+Z/94W+4AOuqK71lmo8L7y1gxkJplHKSYNY/
uGiA3SDl+s4IMSC1341JAMz/qObWMpjkbnAssYauNqSlwKsyCzixRd7QDTNZ
5xMh2+LZVHIQyhYCiPEs104p5lIqS073JGXtmMvvZZwA2BEGufjxj17pvmg6
Tthy1o0o3sJhj9D1/uzBSXi5YniFKjYYnr6l32CzA3itoqlaj4+BuQRyyPEy
VdSwXu8WLfu7wwa+RSKCvYPnkVGts6WnJM6TwIBfwVPuT3q98ZFGgLPOMjk7
eGvOoiunosWYw5B6OSSXWrdkCqxjwDidBvXXd/Y3FheXZewExbBHoLcN01KJ
j2IctVbHHIWj59ZSGOwps4zRKph/9+9EjDaIAtms/ywAy5y7hMZqd2jvWKFx
0Gsu3VIS+l0y6hpWqrpSuKlot5OmwJI6DLFWiua1b6YJtdNEFuOg9MXMin+v
My8aUCB3hhOqyf9gyVWqxTe14EAKnhjKWpEUc1PPs+MF4lbgGNywcNq6f+CB
59L3up6XKQOeDIMWPQGuQmZR+5kpPtD8EVkWgKWR0gIjcaVe2rHK+atHe51Z
eflsF2+yd1nrBakFAHvXQnLJSK+F3dMWrOsgdz3kDThWMjEJ6Bp7/oxCw0XM
z4O10VQjb4sZb3uAW926INg1F4JAk6sGTWf12207Uc/oqDLHwhurmCzKNKrL
Q1CUYysCSkp4BF/14VO3MVBydXA1ffdCymUafghx28qDHe81/0+WHrM05k2g
9YXzZlkhkMYrLca8e6rnweAPK/P/3dOu6fuLEKyovUWe0lNbyofBkgpJduRd
yU6p5sBFPXfBjKylzbRXXgRnlPRtukMYbkB0nJ73+6khav6E/+SlUGfTB+Oa
keE0LqMx5G/A5Foq+SVE/0YMSpNt8wrKFsetBTbS/TyswcT5V7uCYTG5gUWP
NItv/E7FXkwlQLi2zN8jyEfCvNP0VEQtJt9Frle4IQuJKdktn/QzZoY1WkJ1
R1wX+vkDX9i5J1n3/XJ10xSXFPMu/7tak+Qr1SBzCPb4QGiFLRDqgwQpZ1FX
ATb+2eu35qnbTlkhSQUJfHPt3/NuQ0wL/f6cnc+VxVTVSqHXwVJV+Mpf+2hU
tMIjhpUCv+TyjjJIJqqGnaDNw0BSD42ikkPvM1NCE8S/TUaAjhMQwKxXVp8n
LNeCzUQzpCxOStXb2LeWE2fhm1m5BxnJBaqnFV/BiBTMc5XK5dTedWdL2Y7y
DRVrijpiMJx1RTrSCMiqWib6PCMuM8+iVUs5rCtWarznwPJsNpOB4D4JVkAr
HJP1lno2mUFfSz2HhYQld8W9iH6wrbS0xSTMA4XUr0wRGxezFHxqR7NdOQ6l
FPzp058huTQeQJMOLzH3IWypm31U8HwcKBRMnMt1Yi6dd3e1Cv7g/zKzyaEC
+AwmOcrqXPX7KqMsn0gFB9ao6po+J1J2+o322R/hn9Qf08t0i2hNo6+lZ9Pb
J0Wl1rp/1h/3i8l0bEf8b74BzbJhcx2xGbPcDEUrHysWiDvTztfRX/09/EOO
e3bTYHicxUnM9oMrdB1Ad2Zgw7mXVE9aGirJtl343qWTYh7Zif9m2o37VRa5
AyXEUPM/okAS4sWNRyWAqsLZpyd8HXLA1ujsV/9+6SgEkieZ5xsY4HXDN88a
5VT255jaqNDmq6EIpaLL1GoRKCIaqmNl6UpcqC05cY48qbLzxv1TUgluMG2x
PU8P9REb5A5QOseBE3FNDDBRXUyKan4KzMAPCWz311IzhjA12zmRoI/OD1H9
TviD9XVHtuLWHC7MfgL2AvVEF8xEOJR/U3jIKYN0HHe7OuqoaMsCR5VP33x0
HQBHJOOLSpafR+it+M2smaBweyQVkgEwp8bH4cyq2LpTDxg1BmumxAcoAYm1
chpWpbXYW5uRo1E5lX1hAfeNILt+HfLkwGjueNYx9uWHvKmJQuxJmmcB6d/3
oLk5t2dZ/f/vZUDyMABHh33fJqI7A0VHHDSVH8f8X+dJdaXiXc7AHYI0RJlG
CnMgnJsFgodmRkDHw8tAe8H1AyKJbuLoPUnrIhrnEZkdKuMVGUZXT4YXZr2U
MxXN2C6SBtzTamnBR/w+Q/VRLI7OaxPFdFt1axnCKX38PVulZj/CjKfb65kw
s4SMjPzk3QpzbZjHA3O4hRe+OL6J9tGj1c+H5INb+C99x/35NTO28+l0b2YN
Cz04HykWBAYiR69T3+uiZ4qBvASjgvI7heqauPeqZPGZ1oxKDepBul19FtrG
4mLsutWAPt44pZG7ft8kg+R8X3pSm0mDZTpNZZpr2f0fb3R9S7Mp60UBTlqE
Ml0cGv6EVolK+YE3jm+sba2tviEiFj/wAjiWDyVLmRygD1loSBClAyAoK+89
jZ2YSPFla92SOvTGXea3KX9Qeyn2XzJGty9w35dAxNw71kg4GKVVe8r3v8+b
j87xvq1AqII5CbN/W2VBSSxyeyBF/n8L5SLocxsGRTPekkAzvJv6mowu0+aL
GvlpldCOZr4kvsulyFh96nWm20XI+wkfrnfQdchfbb7vP4D5JkMmIczbOrYy
dPq4GKTi2xNByoOTB5vP2qtdyvXVwANIx0n7XFa7HLe/ODLt10UEYKcWySuK
KfNy2WiiAdoEpqtvNjGl/AhaiNHal4x946ujYZju+m0lQr4+J3qtYmCB1Vqk
beHep/nLxUBffUDTiWhqCQ0NWMzhBbxnkgHSxH+fNJdYdGCpsYV9I7kY52bC
uzUTKu6EpxBAWGMQ+YbrYRCa1Hh6yoGtrLB2UEYM9yIKnsYUV7XQqrIgmBET
cGHICOjLWtoWR8l2TOpsA06oTxKphH1mungKWiLHVd3OvVM4k1hDnELeH95N
gF34MLXmexm0WdlJJtd4Yry8+Uuq5ZarJak0I+fZFtbulMUy5MVZqVU2zKIz
S6Hbwu+MmPd9JqEEfxdI0Ld1WEHZeiNPtU9uFKJF/o1a8556SY54RGOwYzg4
yWzdaaOm5n5IsUxyPIZ/moTNBlPeaakkSfiawR/r2241eI227ZpopA/eJcYE
f7s/NRib7EVq9tnNga9fJNg4ayrvqjR3XyYmX7cAtonq5fgRUi3eRZQoIhXh
TMSZQb92/0sebTQTWFgogpaABaMzaaj6tkmfNCiRKpAberNQNJqzISY1xA+c
pPnPjjqFpy0qazFawrv8CaZgBs1M0pUNZK4qFYzVDgAIoHbSiF1q44OnzZRe
auwV00Nhb0L2i3oTOQg4YQ68nuBt7d2Wvvm57/Z+QTjO+/vguYLFlDO3ATbT
mORU6cKdA7vRb8cHnZJdIgoTQtiAYHvAyNwvsZ1xUVX5TEt0gZVANbouIhxn
jpJq8t/TF2WA2yS+hwIN1LbD9gm826WGH94HKJf/cV3rcIyRmnhFTudQTHim
iTWdHJ03tU/WZnNU/RYjhuGJq3g0hNDg0hyb+2H5AR+6mBS8RLAz8XbvtVSF
8p3WjaiWwo2jKCm+x5pYLfsqt5LETojGRq0csYH3Q8cXesBZiJBqIlnKmuWR
NJxsa+3E+cg0STTr78BvUfTp9xKnFWyMS8NmyeYPfrWzYt9uHhozWpG9n7JE
RQrqU+yifhHWL3k8N9OVUhGrDS4VcI+wAvsVQluBi5cZlHRup7O5Am60uve5
kXhXF6pc0ljUa9bT/RAN7P+z1qLqeIzBLXny3KtbyCYNVExcTTO9Ys6v94nx
KzWGLb45B184on+3+n5YuZZf5xeoOe94DJ+6eNVCsbgDKgbAVgfYJpsi/7/z
5lmJkqZA34sQfM8VP+AIkePfiXWvFViDpcgNT3vTkmwexjzzczxsYYCzf6fH
Ku9cz8K7HN8rplgstpAOAIEvq+jG2bpnqWxD9sUugfYBgehE2Vb/h0BJclkB
QcIicmy38j5u75TpF33cgQHcOII0nxVipxbkOaySoHSUNazuBtlNtcXup6IY
3PCvmOCCHKk+ooUUyOfaC7/FJHkcS1ZBFO+rNKTJ+GtqqUNasHwS9l/GySAe
InBZzME1E+FYj8XJpb9HD7zWZ4f8E7tRkXUeHUKe1j+g/KeYHMhvwSBt6QzB
hSzwRbfRO2nG2/huGigd4N9Gu2z43kccXwbswxM5VbKVPufZDKSEvvCMsvzz
ABHNfJBIo/e5xIj4Rke+D/XiyhPB1nRElnj9GGAhavui9TP/OodpJ/PEFAxQ
XVMDxTY+wv060fP0wYZwZFw1S36t0V6vOFuLPS6WGAkZwxGt9zdfbznijxAG
BkPZRgL10Iw6ALWsdQhvrMqZs+b8wIzBEeS8ZP35P/KRmTof8ZW0Sfkbu/4y
KWK6RLl/QnYeSGLidT0cbII3Jb1ftrkCV0Eo3rbJSMZW0pIzB6hlRd+68LlU
H27vYz9j6QNy7jekWt0ILyZ5Xrs0cwJtkoxv5HUr9cQ/A6WF5FtXNlhcybG6
cpFeqYvFe4BZE6WJM69N1Sjt1pI0OI1+NCl9vyhNmGGnnD2p9aqnMM+xRocT
jH2cBdTTU/hgJPc2EZumia4mz/tK5Y30QykzBnYwH+0bZvRxmpu6Hr9Ua65O
ML0iaIfEOfzlafAQXUbKGYsQWmpoEN8IP1reI01LTDEs8oEoytzYr1C7Xf58
d/xm4JgA+V8ixZgHJ+xQ24D3YD98OqSyazjNd+6mjve88Qv9BohUIdAq0Mvw
zWeYZV8LMmnVXTcou9hcMPGfO8hbO2sl4Xm/T6zO/0+FB4o0L/7YEvcBC9Xh
BZ3bRFLQ0Qx2vrOamEyZaWvPZw/sJPrKOWCGU5J7qJM+evuTB4W+O11BCNZd
l7EnZnQEmH0N11YLGF4wGccUbeLC57WAGAL8Q91qGhm58Z0TEp4wR5uB8AQ5
gcoGcZ2eRTW/sq7Mpot0SEyoXDpdHiaQYaLPPV2ZuRt9R+/7ztHd/1PyQDjz
Q7kO4lw9gVKUrJfykwNvsciyOqmoRbSSz0ZlZQxcnQxO6jQtRkwhoPlWUPR/
xNFe0Wp7+lf0RC2QweA+4yKbzb6Em9MGpufT58FGTZM4WI0olu7tMC6Qv8YX
YgoO4mqkhC15kHBlfGZdfMMZFCausVJPnvcwrI+YHLIfM28LNXWJhbytcl6f
bA1n9PoMCiVzpdPoVxv2WNuSQW/4PPLiTdMn/BxvGwf52o97MmBsgfPXRu/4
QzlTqglB2HIayoZGyoraettVsyn5xBwwaFEwB1CXQixeGJzpMr5CST85xb9m
49vS+2Q9g12CJMf/H+OGBYO1icq13zZqpSpBVZ7O8+Jl76ElsIH6kVnEfBU/
qzlBBm2oP7sWMGXUDs+FCR8xh8clFLmNLJ/InkR6CAFW3AALzqqOVJ+XnD3t
Cfk7rhXLaifmtvAE0ez4n8NpJ1K1bSR90dsCdORJ5gdHMJZHck1hEbOlhL3B
LU631RJwmJe1/VuI5AhjZjHDkXGFFcJvW4Go6lj4ts3X7rPVAx1UkkDIoV58
HD0Yu8yGiApkreFfY1/4vuho2B7zDR80Mbyv/NVYeEZcQNnLl4ZhNmwAmEDr
Hylvy6YkuDp6AlaqSlAnr+okOnS5fcH+T7p9Blec5qv+95agYsZkviGEA5AB
vh1tm7fjupiqcSouT2QiMN6Bj62nBRAKTnPpz6dXpFQh/Jtt3l9lA8UtJsOV
zDoRkdge2UYhlulQHV7xI7ChCnwF/weVC5G10nC8R8XdTT0fXO0+DHCM6lIV
Ye6T/an8nB52JkwYV22iA/QX4q73TXDnKJk8uS8hmWw/pMw/4rLBerOr03dX
40HtuE/eQagiuYw9ADqI8Io2TGHBDXCjJHSVICCHd8UswQInz7OvgroiWrF+
qqg6DBVpq61h7br4eI32gU/SNdSN/emHa9mTWuywj3vv6gjR+EZhTda8jG+k
XO0DIq8iheqX/gmngfxKXhOoclGfKu15eO6IBDs6reOHnBl58xxc45iXhEOx
pdpGSG54anFiEOPc/tF4GvSBt2XjcMXN1zXvUh3OA11INme2BeKxEKEOZ68j
llH6Rg+lQmuqYf1BSQNMDh7JCNs3Sp0sWCKWsGch05J0zFT4stt94SlUdmE9
5gFpG8TaCyL99Bd2c9+NrV3Y8Q5oIPU2T4fg/D6Q9DNmuCTO+o86kwmOgE7H
ipRhixiWQtZx/WdlLn1eDVEsc9b2c5oiXlx9fLZ73pxKNSC9/RLAeF3OnfoJ
zZCf5UOFTuN7lZprd0Gr42Po2hLBFz+z8sd5idR9rKo1qgpndULJG3PlZ0Jh
s8W1v7x9a7QbQoFW8E41Z7HjlIurzZzQCGCCYbqEMvS/DXj68igctn6vRs/a
wLaX4jVDpSpuuua6ALuvaefVR9M+tq3tpWGTmf/q2Gx/1Pte/jpfdeQXu7/P
6NWN632gJ/j4gJv6VTW4qDiblDR4xwQj/IxODxgZjdlTNyr7DiYaJWRfcrNY
oKpoC4rackho2wrzOGvwsS9excf4NNnmhrxuThBUDr7EWW3X9ASKV+MWOyGM
5DG9iApYatEAHwawTP5M4bX9KFXxbh2vjACl2cfF39jxbClNRepJv6c/R8h8
SIEiSNlmlwfxpQw0rzFxH/HDo4KGSQ/rczkAjDto8moAEGRIV6O73BMOWXqO
Wju2xBSpPTgXM5d299Qy2PgTCbn6J2E7t9McunmNyQ4/d15oKM5n+fYiQKTm
semVUgPvTfSi6p1+l36sK0mVS3E/XvNgKdvY7k4aYvxUjd/6hCYNiC6KC1Wk
PaqPvIaqHDu6D7aPTfyqqnpnw8GzFTxtiDj3mpglAOow2imO/Dz3C+7mmcNI
GyUeJfYRCdK2IvEMHGAdOT/O4EKX3yYSbM+FJbqAqw2Xc19GfJdfyBq7EZyR
wh8Sce1VFmSzJASVJ4Tnssb0TK6/gps42XWcUoMn1MWbO8+XLVj9McLN5ahj
myaaTUaQNsldusbJYNXmrR0EaTvw5KP1YL2PAV3SiaDJeM2YG4/VGx5EDWan
3yHjRgR9KNwR/JoxuUsInizczsznj3uAdTZ8Of5Ps4jbOVYz0Yt+v4aiMTYH
/vVf7NzOqzIFKDblgZnPWQRD90XfP6b1zwwWxr9/SG0pAUaTcNf8KZo/K5j2
sCyoWoQV2WYGLOPExxGXW+144VMUUMVkKTAVDlPirMeL2RqF394hByYhSxwn
EIKxU2JlBbaWtXV19kXo4Xb8Vzg34rGu9wqx8I3+MStOX2vbK+nYGG5guPw3
bRVn/rg/y3g/o/p63hgIh+Ooe/39/HqcWXW9df7xtgX1/BzWaJ0gcfS2Kwfh
gL073xvnpjzjMpo3I2uY0AuX+AR7KEfA0fHaPo6DR9dTmjVapW7xdcy3LC57
19Cx3tR/vbiDrOVuonLEJ3zN7XgJl5nldtiLheALmlyiXhiyDP5sk+YodqII
f6DPhnR8GfukopHsNa+n/5IrwdjD22Sn39eP1uaaLq64I8CB1Kw8uexkq1Hf
RH+bn4w3nGyLfQveQknYBkH4nAcg49j8xs3ZH7ltaQZghA+Ih/L3EpaEvp/m
0f1cLiayo3RlGi2Xmrsv/Z7Tu6zXqS0OCzWaPFThRo8QHghWSSdBt1FBZnCn
KMLtdvn7o1pVfWxXgOkhGrBXIK7q3M1Rcy20OeyQkADaNZsc9nX9SlqdZgzp
hLaJv5OxFPFMuecenzxaC0d5BP8SXDBVDaGChHm7pyrhYjqbMFV52v4ZdlgJ
E5cAkhYhlGEcKq+lJ0abnEPbBOakePVgWxoOER4/nJ9y2HIW0ELrcoaMZxjO
rH4NOd4djrsz8+wBNhX5WZxU4S6tE7c5F7XearYdH9OfOTjoBXk5vGfMO32H
s4hwYM3Tb8umol1JuIpCKLNP1s+THkcbMPpsctMuZnEmmgBieEd9EWo3csWP
hb+KaWA85WUU2TV0fZWR2stHeYhLcuKOQJHZTQSG35zxNSnDywesRZVK4mJ4
C2ClHE7UhKIl3xjRTS/G3lVOsT6OXzvFvRy/Gh+CtZG2eK5znCbGxxpIuUBf
Gr9ca1ZneG4tYNiCMaupb1QuOoMw06ZrKJN95L2M6dkG6z3KF+UeWEWngJm9
JFwt0SPoOzGMxBiQJa8aq419gzwU2p5G4EHvGUseuCdL7ghO3pZmmD/ciz0Z
7YRwdouQz8hP1QaM44cGDloVP7KS95woF/jLnt7lfziwSzqWkOZzimi20K6z
qxJMG3RlS4QFWQxja1tCJn6835+rPaT9F3bYZfbhLRJDy3j7DFnVziQCqLUo
pqTOm3LY2VMDm9Kn33QNE6s2A9FYTQ1DVrXtwvtuoUsSMCUrXo9WUIwCKUwB
+fH9EdpYDt3ec6muc5pEbpJApNYpFFK/JY2H1ae7oTOdPH39hJBayzlbaRS1
+zuoqVXeiLEse06SFxMWsaOuCnv+TZY1H2yfMO2kb96vfeKQ3G+gqG5wVzBh
iigGUDObGbzNahrn0IDOLx54cdxSBxp343duOspvVEz/Kak2KI9EI+EuqXnr
2SkIWaZRyuJAzruQQ6uGIa5+OJ7ncjW/kE2QY6lh04M/pjWsm9m85mU/AOWI
iLARVtTiokXZlVBXTrPS+4I9qqPa/q2Efd0aQewD9yElDDZ4fyvXyWLoQicD
dfYly6y7VR2rPbCYwaWkmXI2ghcZ97yau5VNgE+Mwhx5hYxjLmHlb5HoCsHs
k0kciZ4M130tnCW72L9yT9hVOJIFs6chRuWUAgeZ0WnqAkSXYpj0nOIOolwj
QwVyAQqw989wIS04E54zjbXkQYiGKFkjUblozTccEZFej+o3qymIETwLtwyr
z0DqsVg0xMmacuBvrNKu17DB/YYiIwtno02jQ0yQp1GgmBk5lGjPpP3Hjgy7
OuErhwaU0eXrvEUuf2sFQ+KTSZ78IQidsUMtFjfh5qb680kTdDADisfEoJWk
fFWc9KxmVkgXOFgrU7ynx4yFJUqatzkkDpiTrv/nN804cxOU6/vNaGxu4QZ+
b8JQAt+6sYetkN2YP5Pu+m0iempYiJ45Dsl8q1gG1il/jrYpyr1/pBNLz61q
A/KJiRPEPQlCKeyBzQXUJSECUz0ymRIO7tf5hO0utWe+rs4+i4TgAd6i9Scl
v4xMyhCwQSCFuCG8DD/stLVQpZPys4XQFWtHSBOsNqMuB0jbRBpmoOub4fB5
YIiPO2DcLVoQMq5i/iHj+U4X3Bi4FYqKy64Z1KjZWN9R3F2Igi38lGxwoEWZ
7PxKJ/xoDWhxkhHjUfexQ/hpFfEys8qP54UPC7QlxnxPAcen4iNMhG+mcsyY
e/rrQJPM/71Z8/ndurc7Qu5G1J8O9yhCgho7usmptgrW4dBYKcG5DxAXtm5+
GAgx0SD/E8SjP5uLLqVNaR9gIVzcdTpugudS4OiDmKpbDEbKw/58bHsxr4Bt
sQYTSRNFv4f8pkR5MQ9/miIrMJRo6A5kERDisSHmk78vWwW0ZOO7BanqcGHn
ZgthydGn5zPf6KV96oadHDo43AP64aLVUFpmVaNN59wKnElwwD2x5BlcOXXP
au9VL61XwzBU+SPT3gcXkuD7oVOi/XwhNw+MWnNPm99FWCZzb089zriVB45S
rjQj4N/qZ6ST1A1VYbpO4+0kcRuhu+k/4VFhy+mzrePHmfTsdu/XoOYtlPTo
i3Dr2vn83Q5uOYgPaZyTt+Efq+vb/ZjKLZeOrGDvhBV/qIQJlVj2RAz1vec3
W9wpera5dw/gE/NuwrOeGhofTS92WvkKyJ1VrIZwwG41WHLUEw2gFhFJiP/r
Zz6L+hblaHDtMQFHaFyeCZ/1cfXg3nTRChhjFunPdelBMQrP8S60+EXzunyB
h865EY/6noqgDtgoVzR2L8IZhrfWHr7P/9ozZ+KcaOSsmnUBei+9ofqWaI5O
/4jp+MlvdT0ArflmF6me8Kbc1P23PQ2lzLyVj+2AT45p6ru87FN5lOiFPKWE
0//ocTzyK1qUa2YIwjtMbQUg5/Fc3N9KosdMVNZeY4DNDAPbmAPk7nI6rhAE
pX59oYo0Kx6/tD+7jZgYgFoLFHQZJ10tJu5jrVJ2/y//8r3Ny9lD5Ptz7zW+
BIIU7VlxjgKG7cMDDlNsZy280UxbXlirN/ghc29TwG71Y6rke48KduqXaZRj
h4LdsiaD5TsgbEfEf+uDmTki05NvmO0NamAUypMX4KWCkAf9/4UKTGRHXM3w
QdW0huMlkhW3HkFv7g9dKYMx7Rg/YzBY/n64kMxewNli1+1nkJqzImJee+lB
STWoPImvCd3VQ6m3rlI+Ru7x6lN84Kxum8esgBf+L/FIUnVs0qJ/yBe5vT8q
TLnvCwLmS63Q8aavt/kWmKgPzjsDQweoGsPb9Oaq8GN8GcQOHMTbQTvL3+CH
wqr0AMlWG7W87omHxE1xxbYfS7k4tCLeqXsVrsT3UIxSpxNa5kNM4saIxVq/
TufUw7QIj1/mge27q+BctPlXLzNsTj9gqVAHa8NRZN/Ly4zzFRQwyqZw3Moe
l6wDf4qGVT7r0vh14aXpOPZ8EDK+CoykjuECrt0y2nGn1F+zc2zP/cpABUTr
aaxU5VQ7ernlRn2OB7mOxTtgmqOS2XH5L/N4/FOCkUP3+/jLVVTtmXW2PkO0
Gub/LoI3D6G3HgExfyJOYP9Uh+z44WOGyGfdpUdhbrIQzohgGum/YGUynSOh
1EOKkxJUnidrajOzdOc2AEChfeyKAiBZy2OL7k2nN8zH4smUiSTRFxC5MFM0
37j7ue+gFHLH2Qgdw/DzTveKwc6FG4klr070vuX2lkD2/khReWUM06tes17E
Rt2rT/J3/ToTq0ggwfBfYzovx0ph47fjeWB+/U0OHyUNTfwkhk/2JBtn5IMZ
j66TLHghGfUv/Fb6MEaDttVWmb55XYRXhcbjOqRkSs7gUDX+OcsTNJBji/7v
bBQwD9J8kGVM94/LEkmITjv19aAKD2dzYSrAeA4byyFLm/zG47jbWyqc/NtY
8ZgQHM9sVeCrI2s+vR78HNBZDzTfqLviBkZso8MKaB17j/CzZOmQzR5yy6//
2RvcmaCBJ3t+UWDwdKPiToyeYM00VJiYLvnxDA4G2AEEfXyOGDrf51/Ph907
eLBzWBFkg0jxuds6Ck7YikH44CL4LkTLtFz/nHnK51Fszbm7quRUEeuJQZYJ
pi4uBHLtQ6aiASdRKHNo5HQXfdy4znGgpKUQNXQBegCaFEQyICVeqaXzbzNL
jr12Zu+lNIgRIR4jtSDCvqxWHhOZZiw10FmiOOq1ExqCWduCbjm3vTarrc58
jEgNwUO97QoNeuFJSacuCNXI/znL2CPvs7eXWE+8OMXYSjreaC8SkLxtscG/
VDkTGz3d3+ZyXqyFRX0weGhWuswKgee+p4EyYRLkl4es2yZc9wOiX5Y5Krye
RBvcO753NtdNaZCNi6OpoeuvSUZwr/h4ffkqrNWRzYq/O2WZ4fiebUT6qeN7
FywaMvuNAoWDabmFr3fI5kpYN+BLQzbJBgUJhyoQ30PoIBoir41hyaj8ZnlU
T8HWBeNLVeAQ6CPB1/bTAca41CpRxMWwBk6IsLuR6uIY/cTVcttdbg1Y8cdW
6UFfCB4cusyP9tVSibrGP8oi0XkXszkRtnmeA5zxApiyuBFKXt07ZO0FnSxI
h70ZdPvtkgi2isNu8SRjCQ/CnHvyFzTso3Ph9m5+DXx9g5AmtDzPS51T1NeK
GawpfD8ivBpbslp+L/uLqwM35OGh8E+rHivQZZQERVOLzKkezWURwYEMPG06
h5TyhIGDdV91CWXAg2bKZRpduyN5S2XRGmQPiMZGQzJM+5rJcns1ZympeBsa
s5J81c8UlEG5UXUiT0kA2wE5vGKWnAkYAwLdR4l18X0zBQjskj7TSsOZNEyC
cfOnXble0a1n8VxgWxFCo7kklGE7ArV/DqIBeuDjzOcXvpG/cU9vXHWZ1RVl
5zY3G7mkEM+raEBniCC6H/CPZLx/nGDYyoIYXSblv70aqCfZbroFc6xy5HG7
I0Rh6EMmmNjb48Axj63B8CgKHWfFhy9lopyapxxpYz3+xvSC2HBBAHz3EhQS
KiLQsepvFzPmSaUH6kseBhnUme+px89ahoDfO//Ftu6ggvdT9OrAQyyOlfSc
HVk4HNRtse9nzThhgdvBDZhcNdyjv+Fdn9k7LubBsp+jDBjLMIHWairDcUTr
9X4eANZNrCJ9gyuQjrJPtQ/AgxPdxgMdkg/nBkDYtPYp+jeaNa43ItQMNhMR
xA1vJAVRkgEzhcQARjOW1JmwxCvroUePxKOq5V8TDblQTo1fsyWFdFu+PFR1
uhh20clsz5rQ847Lfeflz7lP6w6hvvwWEnh048XCIvHz6Cr5aR+ra5YX+9Ll
eB9JxFirLqIlBJkvJAmRXP9yIFQsKxKnIs8R3YqC6KApTFylHFpVEMGivAoP
Pl26EHhiimFxa1Fz6tQKdKPz2fRoHRFp07G1vj78P2eMG8Cic1QWLN2QmTW2
bBkSQUR5JW6Jy7NfloBI2UBbwjxx2UFAoTO5fvXG5M3JAEN92kbO/6kjS8yn
yFDjQFn43PBvEf4VK9+S6VaAYYovuEaWrCTZjq11QfrFySccdsja/X8XMPJu
hqXZ6a5sg6zRm9EyiwEw0om/CdOLYtwfibRAPcBbb/Q2H30PLecrSHGoz3CK
w/k7llnqo7IxUTKNE6k7a+tueXr41C7OELWRAha/Fi9XqE/InRo4lEByouwn
aSzR/QQ61AWxQr1YPMOh2GaxACj/coOHSLLlswjKJwhi1Ak26QQux/9GJJhb
7lLeDPkCJZYZKMZKq9bB08almwqREme5iUn6kkRYzfcV+Wq0eTx6SsosUMuo
y3m5ENPfwlpZ+jKJEKj6eMou1MCZx9V1YKFvXM9mzKlRIXf9R4g316TGgctm
kxtnPg8gynJWcqUJDUNNTnFwnKy8hKcahzNlsqvFF6F+hbwd72WeHuwHjCdC
lsv3P502H4+eQ3eTuTA85na9bnFb68spN4PVJzUcNJJWx8bS1y+yQXRlrvAs
dHjdNErxfnMaB0xu68zVqyiBaSVDhLIFyxia2XNEii/VDic6WRmBWz6Qbyq+
Z35B4Pkh78fD798Y1RGjjWrMHd3UduOmRkKx+mQ+bVwvhqOovebfOcWnmd6c
xUnHntDpgFo80D1V3Ysatp75AIW8Q9710bYNlyvIpaz/CE4TTb4mgI23MxDP
idgJzAzezyt/p6JfmOHP0e7e9uaUPmBqBQE8pDDQwiN1TfElp3WEixoah3zv
U/YBlu/hRLDNJmMKWWGaHTZlFYyuHQDYRR6dbE0IvQxvIYwi1wRcZZXl1WO9
qI640MqcSIyUgbsIBCX7TDc4guJ6wxXlvz8S5DR4KtO5Jxzi9is97IfMp3m/
mgrhgvs9qlhNhTQQR8InCQZjK2FvTF/lan/blclg2YjaAzw2nKFekwl21VJH
s8jr0IiXImFzMg2CWDgks6kwbccy7mgVfxXTfDMqxF2yq+3Vx7WLBXxvHEBh
9uVDoaY7ps1/kLeiYBa5YgyNOGz17k0gOGANGHFLXcBfsotcvCVR7MA+3M9A
FNCTvy8VFJFrwje+5d9XjVVDvq7G/sbfMO/0H5NacpYv+nkdA8CuESK4QAPM
A25DoAI2houbsoM1UNJgRutNSWCsaPCqua2py6n2EUmPo1OWDnu6Rlg65oMk
LdxJU9dOlg4Jkoe5S8+j8QJqHSedRZYdp2B5f2HL7yVYOA/g5i5HaqRBXB8S
OtKl7GdR/ZpvXoB85WX2ELDK72nIUFz/AhrWNr6kVAoMZF56W4RChQ84gFJ9
opSqfZ0O9bkIWD8/OYEtsnRBmkbftqRgaFUEzNVsVlWI0/Pmqxrdf6IGM/LZ
ZRyynUViYkVemXy98utXYIvAUrQMDHSI4LJiRA9YZ5HySr6wPAaB1jMZF06j
+j4g8u/zd2/S5HsdBdsmIZNbn+tnQaV6D2myAbF0NUR2JzPevIwOwOHdhvrw
HnZLn34TR6Tz6y/WaTVVQRTkQSrwL0Gq0Jq7vLh8n27cWlZhh3Ic+NSwtGa9
pLDCsbY/jBecU0Vt3BfkgMJP/GBWm7XgMkjXSzlIfbsQa87rL57HenBcg7eA
jHlGxKE7BXCWGvMujYu5GVnasoZPatvNH9cjqm1VKinLCTXS4Vvg61S/7Nlc
/Py22aRM0K7UPGAQEKnmO1s81hdB9EYGmykYuTD/llH9RZXWgLfFXcJgrasC
2IRrl7ZuwLAKI2ZnQlg8vOArkdG/skspkxny79rUY0sCPaA9cxId4FS5D83e
xgYtNcRVIPNam3GCwbczElT0i5nEZOu1IZXUYkXtfgE1PhAJJ9tslXxpr9BU
RfK/g6IsPyj7wDrryfJM1su2RJurbl1cr3gCmWD5lprN/Q8tz+doKtsBFkW4
pHU68c0DFsw2uTq2ti3qLRqsXL6Z4bW+IBa4qI0EUQ+TsmUEnHb2iqEj3i1r
G3iD/3JFY4VOnettArep23FbDM0eqmbD75ETWabUf/ol764kwQmOsYhc/3oN
c33RLSOFc+w+J+l/f1eKyxlE+NVFsWoMg+WdtM/FKBXoGCJAM642AtJH1/aw
U7r3tvmHWCGYAPSJoGdpKeg7RwvkkJhOh08eHGdoempZMPP+Vsb6K6gICDUJ
PkR/NfCprx00eH/kJfS/AcejngFrgG271xeH5omoyug46OG1u7gUYsYs4yza
2WLkfszoO/1uAZbkuhBUOKaJGRKcQx1dNmxop9w79O/LHHYu4F6/4e3L9juy
HNAgEWUpC9fPX8CcVrQ2bwXWzMw1vsidPMtAaV4dyg5k7yYOwEru/+s9ishU
dR97P8aZrxkMl/dzOoPI9iomjmMrVsnAY3K3dk+WbYNQYm+U9bfJzshpdWYR
MKnShs8MpCqvV9mzxBcJLNu0bHmKkHc5AS3nErhox8D93YfNKq3HploVg8wL
h9AKmPFuWMVE1+ENxW43IOWZgRiCyJPWjRqYW8Kx3atwe/l4ae0eN6s3IVkK
7ZL70B8uon5m+31hj83v+KOOmu/RT5sN7fUk4GPOcVVAktu8EBk3VjD7LjiG
zpheUBe9wgx9fV5vFsqjH9PDDkq0pDHqQ91aEOuR26wMQWBvE5gcijOg9gU8
Fnhyk5qfPOwEkNeoJ3LAAYgLejjuFpt1vr0c3d+2+RF2TXtF4wKW03RiF+a7
5INo2Q+Fk4bdczRZ9f6N4PE9aGEQn81/edOM0xBMET6n2Zz36xlQKtsTgLg/
YxGT3eBnhNGEhP0kC2IHqjfTV1mWykT9IhxISoN6A5bkalka7Kq3hESOpcpF
EllAB1D44eQuJD/fg0tNAhEF64qfoHvSHyOTZ7xrxWhkzQomEMNfveeOYcSw
18tMfUd1g/bdXK0q3vki8GNTClmwrs1zl1zHKl/6v95ED/b21kuf4a2QaLJS
DO5paW+nwXJBWZQFMEGKDh0scaVWkBy5X6qO0CtHgFEwoxP0guN9cGUXPUlK
mG6544t4d8VGTG+sWCkoRD1EoSP3VYnpN74KLTmJAQ4gbrnlUgFiEEn09SM6
2frPLLccYRm77gA8yBHhkkEkGBw4Qjtil0YgqYI+mAuKqLIz9h4/dQ6D4WlT
7SdMdAwXgDV5iz/SqtwXqcir+s+mLYxnY7H3JwItznq32FOLLmGd7RWeIUWt
/u96Y8uQQqdtLUz9FcShbAnvKsmAnOp2a/PmCkBWWyE+rNBNYJr95ONoLlZ0
e2ZR0uNx3XJmJOhOhojCCVOLbp5HWpHPTW/mhA+EjA2ZbMV5nhLlYPvJIxuc
fmEcqebsRgLTsAwTYbub+JZJxPlIqg8w1ksefsjryQBIUcemX2ybI0Z53Ten
LBvr3/XeWbshi0xRTM3dywhcDP/unNgFSrK3HCcQguXD4kNZz3i6b96mLQ0C
LI5GiFD2gjbQbmN7P5x2dHfxJ15uNzBNBRhS6IR2kUJsE72ooWQNNDhoVoUF
t0e3uYK0AEcMJntAJoNtDO51oh9BmjAMZ9n7a1GtuKLYIn+NubGGQRwdayv5
H7UlYvPCQw1tzrb7DZxLoPFqHinopL113MEw+5RXL3w6ctYvGQqL5ZXxnHnw
uEizeC01ejcf+4miiF5GOvWOYxfVyiqwCwPD32fyMSdwK1kN4dcOyzVlc9TX
D4CEt4avTIYRFsHuj8y80ePKjd1Z4sn9DvmR2Jn1EvXzs5cJC5Lk5PhMUeFN
DOD5ViuVBs9B2H2JVT+7ke/LPuit/Lb08SoBhUYMuAK0cErrcEJtjMjZJxgK
+vnG1paAM95RIuAHBxRz0WaKvcZwMXqq2BLhvfi8iA2MK5fOM7sL0Bs45d8L
BMTEaDO8cX+3y3fiLnrgYy2F4tK7uO1j1ABtRRZvk4C59UFV2BODMMU+FDQ2
OTKOz9yjLCRXvGHYEPmugQoZELotI7mfDwc7PLmxmzPLIVIvyyHptjhcjjbh
eIWX6/gvdRUHDJLlGe/Pha1frmzZaXBzWr1B/CfGayxrZvq71K1f93sWvoRF
goJc0BWzzc+ma8juvwqVLp65B9+1SBPjxTZ3GA9TcPzNDfhpjrmMQEbTOs8y
JN1futHKbWD2fVkUr+RDK/INJ2l6QHvB27+Z8CBnGAHh/QV9t0v0QmrlW8CW
OKaTP0dsXBbt+v/p+KLS/UzllgAKgqVnqLKkRA7Vn+VaLtUpSo7wiwSQtHAI
W1bh7p1MIHsW4edJkZOi2SNGzZXOMrPMFEpvytocbn//dXaE4M07yQbOYyet
EWc0gyfBhdAb9YEp70ufW9QqLmQ4PA1hYb/PRysT00z8fAzdxCxuTm0KjoMP
b9x+BvZuq25NZ86PTyO2TDNGtSa1k1Bi5wavP30Z8Z22T6weKTGRNpuoFyWe
24vD8hPi+HRvcqISmgidv0ntYOF140J8ZToOb5cO6Z8hqeamHbR2oU6onJy/
Qk8cmS2yvZD5t1ch/Jx0VMk4latBea1p2ELlT9aYev2R+GVbhYoyMmr3HcN9
O6JxXhdwJ5YnL0IivtECmQmAGSR8A9oIxZra0r1IB0yIW4IDobRUi/d4V95Z
dTc6kF27lzn8o1F8HYM16vJHc8CCuMGOKkvvWPfdBiB9PptQWLqe26Ynvu0O
tHVA/Jq6GJ5feBInNCU59yy/8cpTXiNmrfh4BE7blGFt6+Y7G2lE4TaMGXEW
F99dgF2+/uNvNdOYHCBE7M1xOB7q+H5nTR8ZISBY4uobt4BJtu80O3Uu0LbS
v9EWdBtS99AdBtGflSJs8WcfLv0WxIaGYgoVdlnxbp1NQQVGQrCwr/BygvoD
BOZ5e+mfiGdgim3vRT1v2QkJF48DWtLTDRfP9KRz8yNLQYbZEJaB9NaMGhRZ
v7TeEuOv4AuC9dukyhp5oIZUku9yaf+lom3G0UpmDz55Rwq/60Vak+aNnD3q
3m6a98RzxXOy692wz3bP6dx/0myl/u1gauFjFOU8HS639tNo6JH9pYf6ndXm
i2bkyZ0Dwax4brSLe8hAO4pb6FtN0emyBGDkl6DGNLtiRLQgz81jO3MnV7oW
ixTHEx2nFrGYMxxWXmM9Jgp+OJwWxvG/ufuQCrU/AWXR889E/vrFFFZBtZwR
GRdXGsSbbLLNV7OOi8VOleyTT/UEp2YQpseoEboiiBLndL3RIkRmhe+4EJXV
LvF1hlwrN0nFodAFrlDi91PfgQbYVkvtHyvyIqVYZhRMtGC9wkHa1na0jGfM
pHOYnbjbbods2ZAJ979+7wCuk8VCUFCwrZv27djGuOYQanj4n95iXsJZgGFF
xSzm2iuYkf7s+FLGxZBkvIK2otaVvdU/CSJpIvpl81y2qDgyAERcSBDP8gai
p514MwOrITCHJBCWREWvoxg36hP5W4ImCTaYK+wGacy1XoAQ6Ta2uajTLa3f
9av6xGNeZCqdde5eYPYXNbLBlZ4CosxNvclKPMOXpT8/oY9YIH6QFqGrg+ug
e/5BYu0N7LiSIyV+tMME34jNqXi5HlFm+CTS+EijmTXu5A8vPUHQlNRunyTW
LSBZmNhBJjwLpc/G7uiE6DvUvyZ2LxyMyzcFcOvfhbub3zRMYRQ7r90g/naa
YTbAwITnAGli8haAqGEbMxPbdKaneHMpAstL0anIxJD0b1vFYJH1N+TrpRPa
Kb9zcCp0TQsZFJFlNew36K+TDjlAao5zp5BalTM+uqKy6gZ74EBFKvkfmh4j
lkGk6G0nBUefM7mGCoxZZia38rCGtBWoMCnD/T8HK8Y0S5WcAt78ZbNBA0UG
eUzcwR8sHTOUfoWiONnk8B+C2awOcYvC4KI1uP//3O/07ajVXy94Rrzsw+WH
0eal8jfAfP3jXmDuNtJscMD91Dij7Zf/6L8ObIs3xidjvSlufjladzY4cKZc
CM6MAJWOWKEEVLnOa6pNXOjkfgXJgJh+ZvNC9eoiKKQDml+Mgd+9PaaUo3uV
1zV22Lp28eYzi5vYReiCrl3+MNigI7GtiL3XdpPnPUPq4C8I5p3HnyGG/jI2
3RIRSamfa87u2cfW69RWivL1v5Zme6ujcjORtyzqJxYWmPNjQTmYx+shvmCG
CsDzLF7WnNRbg3ZNnaXntGpRxbJTvrO/1g1mxv8uJeYIQ2RAm2cv3S6MrV+0
QkvwuuXZVWvMOIdA4OEPSwH9xeNkCIjdWvhmXyyhU8uuPZAAOuahOxWnfLcB
XKbygWu+3zsuyWcrztV5SxT8jojN+cylh2U85djZSYcEgk1OXmr7E2Dx1psL
qUI+8d0t45k/LXhiSEbHO1907ubAQ9hK8TrIrGDbnFZeVjyh1LwEu/J8C1aO
zYdRK3RqqmJAOU/Fzb2jqC+p9IXm9Ku9+OOZljwG4ByaTriA19U3Vp01WeQg
QJ9RvNCqv1IPpvFSKnFIjvym5ud4D46BVup5miJPA7d3QHIZAHsOC7M+qLNA
JnZESh3FiTZfA+se9J0PAF971YM25M3QcyHAwrVFaoKA1Jy76LspV1ARNpy7
ZP9iRJSno4Co6YQzSqA8chfo4Ss0j8TritSxCpZthcm2zkwDsynNESfinxyq
B0f5lp42SEez/F3WzpRpIye1kYCEsPAFRwGlMZlcybc27HsglKpEh/M73smi
qseHGbI+8p5XUfgd8fbNaV3/uVPgrjQwGxddHUm51mNImW7tw0Esp6amQ6Qd
3N+dczp1NLGekxjOupBG9Gk8BEe+LnWzfymnjEv6Xks6k+BSbkA2b4RBreq2
Q4hKn/x85JQ77Yp+xuQ1Zi1JnYZgmoce/nYiePAuspprP1VEZtB2gt58BEIH
zbABLjenjLuahl5iDPcbddQdBQ3NEf1laUhFu2JyJvItGVE4fca2Efo4bcpN
9CgbCj2TOoe7vyItzW5OhrtqEZpYywJtN0nE5z84s5ryNROvxkjaV9NzLZHT
wIQZ9Stw9y8H4AhzX3qobA6ZKNTt1d7HIdb4nWlRUJ07+85aClK5tAe2dqWU
6QwJBOeTiskeX+Q0AnOD40r47SKeLMOKags4hO3jogiuHpOvBNO/67ElvPxB
nUPNz1B7M+PutDnfQtI3+LXY4hSBaExZzNTmAMOyN+1GWCnXfhd9r9IoR4ph
8ShTO4uVRt1u9yQlqATVPEgk14Q0Uf4Fugj+6DZpInY6pKiSaXVYyzci6p/u
QOidKsaVW0mO3OV39ODoZ6GzqV8EJRVBCx6cd+D+fDSxwc2Q7V5N/PKg78bl
ywRDj6hn3az2vWbdArFnTvyc+/SeHf+a0TwjLdmusVAIM/FuFZtdDUkuqT1U
5LvUmg6E35U678hnpo8ZXF8Z0yzsqygHk+1rDG8CgDhjN1qANIcTrEa9wLea
+BtI+/Uq3u2dOwPUyZJmhCGCK9HMsJ8aKmreQr3mStW6GJuDenMOuHSFD8HI
FO7htLHOe0yPM9gdxeeRfU3wgKVBUH5d7Do0SWO+7onkHh4l3Bd2jwBlIxWv
MmAhZwYVsopbjMsg+zQqbGFOX6EVc+jPa06O35vnEP4xmMxpBtUhld3YvZAm
HQb8JaMGJa3fLyPoGbCq/ars+7UrH2H8mIjOot+TkWp6h2o82T8ADZ8ttI3o
q8OoqNiZIdtD4XFjL4cV/UHV6MXXUhQt/lbZs8YByq9tOpAKUogLO2Fv/WGI
5aZ6I9fOFTsx3j3oejGEpxVjrGytQwuL/pXRW4YDi1TWVZ289Zb9Cuygp+vb
kgVHKuhEfyy/ldFQ6e9bO3+NvukzjVQw6KKSqEi808AiAvqDASIpJy27UORf
5gWUYf8jTI0HOzZ0sGgZkORlJuNSkeHIpA3hmVNJr1anq/5xLSos15cNFBJ0
X+S7xllpGphOXVv1z4gX6ZNhPY5T2/oWYICtThpX+XgVUWDbGDRP3FwnQXjD
9dHTFoVHRU9vgOYtbiibfRWpyIWUBgojhDlFCnKtqEPIm5nCrAcaMkOSr5Fi
xAX9uj8hav0BJmZ3gzFxNLEoOmZxVCEI4DEf93SGNlXbEj4r/7p8DCahprAd
3l+qqQ8DhvM7d5XAiFPyqCJmLSum9e1oQHGn0CzoOPIfzlJe8Eo7zfOTgB0O
bHeYy4gc886CCVIdEFlJhSTwU49iGxtKwcMgHqXJV7NxMH914PQBxC2DjkM9
J5C7TPuXvs27GRVK4hP2E0rDcgI8ZMETbcknWCPIxEcmKTxxuuAoPLTAKHzg
a0d0CetRZxTjaFWNpu/uZwL8ncCbqCx0OFnZe6p2ikOHps3Jz73WTq9moyvq
kcV9svc+WhOL+dieOA/3cK+tMB5FHB+S1mEFrJ5bTu1oxFgOYzQKb/UZ4N01
dC0Qk57I83axkpvboQM+9wH0a6ZLS0NozzQMfUNTKXyDcu5kV8pkqCIKUPG2
5NBfAE1fDIujurAgo/IHEyrye5b9i6Abj93ermkE15CRCoiYN0GBhi2kJj0P
UsQeWC+pEOTcX+FpG62L0HfpGc+C1dH2vyefAXMRS09zwnhlT708cOoOp5f7
+kc0WS08HLb8mM0gXyifCCv6ESqwoGio6t2A5RJSWRu3fOD5pa+29XVTqS2U
fvbXepozjDOdQR6norI4LMLrahExIt5+3YqW9U9gHH9DGe5I5/8zFPFwJHee
oKgUy3VPRYSRweo9N44kaBT43N0KJA8jAz1sOOppc/ldw30JvzRiQQwFWb0N
sKXQfPQ842tpzOgzjB2Jo4UQjAj39mdrv9WjAbFs/BkJySByRX+hcdeWfytE
/uebsCGkdYFPDv6yBAfYdycIAsiNatC+TqGgwGDte0ldzZQGh+8x3CxGRIej
OhfWM1rpoC3Hx0ky7B9vQzKJI8E0IiGkrErzWGZdVAyfoutPfSDOXHCt/Woj
Jmj6A0+9wYowzdTkHaMXe341gWdBgu777gusDsogVu+IMp/Enz7t7OsoHa82
NMFphUUz/vTWaqLRqzdoKIJBjYLz3sPJdcKk3PXc6/UHX2UNkz9C3LhUTcSQ
KpYCDknHjkrXyiW41GJ9Ltd5VFpYgpFvLo/LKurQypAnOwcSAS0aYPqbPxbK
kqbgE8vNuge1Y0ntRexg792bC3EMf5EMrpEs0yvk5bf99ABbPl7AkWN3/9tu
LS6hP7RajI1Rp+lUH7lGZgzJm0dUwLAGeaa9dLfNh2RMYTVVpLkKWKNnjNvn
AlGMQmHT8SYQchBPB6d4smnj6lRo5NxS004/s3MOHY95mUrgz6pNa1kR391n
6xsX/lVWQo0AJEm6s5IWXqdTSaGqCcjnlhO60fWcpq/BPmSYjplPG6fihF6I
mDg9/0cL2NtxvGGtLXoZ78+Ih/oRak77FpVNbkwB0DymNKBGR1fPDXSQlCA1
zoHR17c4lEz4H6so9ZzWkALTMYI5SGbixdE8W895qgaQdTsT56qN7drF6Amu
II+HjeSeo5452eRcbVtNga1TKDrVTw0tC/urV+KD9nGvIksPC/qffAqnVVnV
97KAjx6hL1pKjmSG/6v85m+Jy3rYDNl1fLR5nIwQ4XZhqoiGB+ZTEVPHu/cp
sFkpz3zvYe9O+yVnK0HrASisGV6th7vb2buF8GyNXG3K6EkIErkjOa+++igY
mSDqfaW2y5BL7Jjbw8XWhhjVCKu7WucGGMmO21i3po13hoe1Rv62tjFUfK7s
jUF8l6eXl/tkjrMBK4X+FqlmFQGCq8B3+eY7xo3/GZdM6ZGhRNcg1hxvH2J3
ILYt/ycGTlx1CCdatxnwKVMzdAolk6gJ3QJdir9np0bBspHFiV2KkwMLkax5
ugWAFx5Ep2lmAmAxIAEOmz1ObHhuo0fe38vR59hU2dX2h5M5+0APnUHhHFG+
0RgNohuVJBH8pRXTLn975HeY6Wa5AmpkaELFNVkMcTuBrbkNPmBc8n+I7P9T
hT98MPhJQRpRGf8s5DzFGZVOCswPuxCS2NWLKiQh1HERfcoxM/zz9I0j8ZkC
NU00APgAko+hFs2de6AECcM1OUTLrV7K9+fp2GSfu2ZK9rOQ5nYxsuZxtIzT
eWjFJyHer+xkWsSvPhA++dazJkpI4wdUQVurAom8pw+UonQrMRLpb1cE7XeO
26vsiffLL+zTGAaXYuZLHAE+oSjpNC4GnhSYn2mKEiH6pTquWNy7aF94lB1D
fJ1u605ArBvmCbNl911JHYQD2+Citnds3mCHTdmRqRrZ0NbeWTlhi58QU0Ey
jIjzs/eszhivnyBjrN8rcajmb0RLraJ4btPq26u5wUyYL+fShPZTCCPd0SuG
9J+8qjzKPzK28TTVAdiEViT7wWCMVTGejzP8eGoqNCWIDE5SlydsuKAUlP8j
WR0SEB1fo+v9ZyYo6PTyd6NBTWZNPDAoHP0Z+uU5588leqjqOnnB8zhMcFTk
SPY1dqKVkYx2rraoeWaBi5vIcPVKmxNvcj4mf+GC7zPcQrlYMuX0DFCT7VnZ
H5Z5so+9Zsu0MSHUxuw9oRkRv3t2Vr5Ps6o4s9jFp02CDmZXKogPt38Cm1s8
fT/Yp7OviLDcwstCa38y8obQgAkVydJyUQA+6dfgUHDxg+r9F2aEH5dktMHl
XnEsK/tPSpl63O7FVmS0yYmb1dosNyxIQkPYrQTPWJ4dLqUHO7PPXrIE/pz1
0WP6xa7zAqum/KVjJsx2X0AD31c/LDYWHhf8To8qek8CDiiMWDUyInI0k+fJ
l+jVowvEvVhjC1bZm/XJj+dKtrNvEiZuor9p1Egwx0553n+GFsHVaMfjZtwu
ryUSjZrj/YS7KYyxiXOXXd7KJpFDxNsHfVb7tWAygGJlAQ/KwysTrUpFHFxT
tCf+YI7b3ais3fAC1ZlWk7vPHEvDSQZvwHxzbvxv6crtwq/g0cSxMbzxGu08
JHz7cj3lZfNwLV2R6UPd/BMpwMYV+OUEMQGLA/F1aDG84FVM1nmbBC71YJdk
3srY4cxb1cMwGsiMdgpxAZMqpPTbgjSqo97JfL/VWse0b5o+lAz19vlqW7kj
QYFR9NqhHOFdn7+rWkYVkipljK+iPYVXYTVtCHl/B5Jp4PaQRw1+BtaZ/d27
WIBT3qVwVviu/W+76dfRus8y3jpwH128QNGM+uH+HjlX5io+Mqt5ALEasi74
Tssdp3urRgFcWrled/+wa6+MTHNEHsAMAcvYscKmAF9qQiJeanwxU7WqBaWp
OQRgMxDcCrvv8TGDq8Hv+7/Ai+jK96drfkKDIHwvrhmOxbkxCdOp0MRakqNq
kKIZj9IQ6OoEEcFfTjlHBQShSYjsXUzC+QfSoc+23jSoXQgHVjPCLwYx9kYP
2ioPRUP2HTVLbwiwyP7JL7Foew7PiTfGFHUV/C6GqRAo9CoR/4nGFlfHhgvV
fhTBP39rJV3m2hS7jj85YjQDinKbKzOXnvPoPz1EEFxAhgEJTb+KMhhIgcUi
8v7/oawzj/bnNy78T7H2FVNhC0QH+xWgF0CqqjUWbofJ/bJPTXflFL7msHG8
prtcyVstMosOYTEhSfOMnDB7YhNZlx30Agl+makDsFIPnBESde3Z19jBlK0U
yJdhKnWbO+9Hkvj9kRE2Zj1S820X7Bvy67qEagXTg8JBuW2hffe3WFitf19L
x1kHResLb60Z5We3hvHwCSmcRq1j0Dnsu8UOloWd+q2RSI53AkyZqeUur3Cu
gWC54YSoqdnGdROKUgVOZaKHELJ5MxYiSWBzjhW37jSNljMNmi8ApBStvnhy
FEmImVfSgO1i7SThdaQ41F4RcWYSahyBrdkY1g4VpVZl6C/9NSuqDYuGU25o
MWEj3CGcKoZpxevMtM4ceY2GyPvORiZOLgd/a1OZwIm1h8o1IlXEsPW4sDNL
cGyeFW+MSUE9HdShNhL+1gCSCCgf38nebgXncvuSM2Qv5+tZ7Zmdwa7hvlnJ
Ik/uEEx+y+Cyt7j0R9+ZnYXGB5NJMnPFtOef4alcatbByv6Cg6b4XaUO7HXx
sQ+rVAv2uRPKRmPf5d8w1xpiwTCw9FrygDbHw+qc7BALw3SajDZAsGp5l6ae
//h8Tn3COp4ogSI3rYvlqLB+VSbtYl6geKZ/r9aE8KKeuDJHB0OUyEAj7w2d
Bs+N/hisCAtOMxIuzojHL9Pi0uizEvjiVACXJqOc10lBabTBGuns9pVoLJRE
dODnNHAS5z26hw5XmBah08HkE/o4QhJD8kJOkEgQZvrI+ZdUoqykU/g24hd2
hzCAb9eyT7BNxaVL37Ao20NZjFL19718XiAiVROkS8IRq7ZPYUC/DcvYVymL
U+mGqSLWYKYR25AQGhit2wMbEpWOcVtrSIQlS3YuREcBmA8utLHpleMciYDW
VSh2PFjT9EVJErFSHAh13LUL5ldHmRVF24hfD6Y4NATxuJLN/6nnqXl++R/5
JlezEI02DqmAqbYhS8eRpFZh4qERINKbrx1Q9XODs00OPVg+HgS2sSUXOejF
p4+Fq5rKl16WQzL8Ydysy01+W0lmaHTC/IXe1xacXy2G3d4SLgv7sCIWGEP1
1Yiio4xghasaglgiqRRGYtOoe7QR7gieT4GkX2ouHBDZoqm+Gy5/+gysknCm
DO0U1WeQvEhuP24FOCJGeUInBqYqR3WJNktUqVGMwgfQ+hvqu8AoG63xXK0c
WVNlrLDv1x6ITrbFEW3l5tZx7oATCySraT3noLY5jxRBrlQ3vo+e7ieQcoQy
LV4vSiitncXA3HHTVGHk0wgpJ2M67OIYvvo+4J1uPN1X7ugLB9B0IvxMuCMb
Lhbm0floP3+NGWoyW3dsFjnVlTJAWydqTRsJM3u938MPOPJV4rccDMMtNwlv
LQ3Jwkk9y/4HFvqxTRDT0sh7vkBcsFHJM2GZDRWLspmpH4nw05TK5mqwUalX
Akr6gEgvXs5XJEdLJmYB0m69aBt2zI6fUOIp7iE9xpgZ8MZzBPA24JOfZxER
Y1YK1sn9ZTDXi91HcNhPoZgdR1OprSywFsM02gAzWWrtoXWzsu9Gn4z8mNW/
2uw366ZHX7rRjQ9dFddqLxhItUVZWdxMCFE2ZASLHvMFD/WrA3FPTBJdQ9o9
VV10LNwqVRJxCuSShgmezACIzBeSEbF2igtslTsqHK6v0HVlYRakTfpymCNu
uVz4nph70MEj/Hdl9ajw2Ja7zn2J0avbsvEStWLlkdVV5b0ol5uAlf6gs6P2
X9zQVe9msiVfbM6jowJHs5FQl4s/H0Hj8VpkEToBDh+K6njFVrc9zNrrly0r
xssu2AHkAFj2FywaTJSzWE+epwktcQmMcQdxK/b+xG1iYB06r8MhoTYpHVZq
UKZmWz4/X4UcKCJsir+03hgJd6JBFYLPBceK26KCLGeIkf9Wlzc8uqH2wnyV
y19yQpnOGXHm/FhQBNTr629d81x8z6oLcv8HZzOSi5SdKkh0WkID+YkVUyX0
QwbOAyD38FXBhMf3d6jQT9SQ3nS2/8ZYAxwBw4rDxwe1k7YqAMvG1Rf1j4GK
Gfvo8/9XhkMIBK67d5PhjbP0d1N4l/p0hC2QD6jbTKTD/EmaBohcXAe8Epn0
PgPRfHIBH6TQ3ifBWgfdgK3gwgXCAxWjJn7MGrk/fq9bc84cBBISZipMQdQw
LLXjSleh7+IX2xrcgIcl9Z4joVG5EYJf3tXG5wXMtWFt7H4UwG8CHWykNTyv
0WhVqKB8jZeWUpO2xwxFR+eYSFPx8Y20GPzY+EZ0wp45WvMeaXx5QoMdY0KZ
NMBZl+MZWwIt5HcBJBxHFvqHw6tR3kM3Ml411FbJkEaD5iN8+5S+jXuDu4wD
hMv7kWQACgBG9D9XRFPwhwn4H0mzfO01bgI6LBJYi+AzCG59/3BwBPptP1ti
Y8G8bDzEiiCEe3rPNfiOjCG38AVY51WZIMkx95Y1lCB05AblRHVzq5sZIp0c
7MYCio0VVOYCmsxUsfvRg7RAE9cIhvfy2iSYNN5sHvwNOlBxW0LNBZdJcE0+
njFtSrGPR/hv8xBpqLh6rFv6FK2MOHaLoyOw4MbmHSrZLeYJViy43+Ixw6Ih
6RvX/KM592JrTxq3nHAK1gjqRpSUdgNIRIbWB6fTg4l7bdenu6n/x1kP0A33
oh3BWz3d60DqurnKBssIUnDol9f8T47WsvxZYp4rNmVUCvsMu6lOTZqkcDss
HAaWhXQaAnFtkeBIshiG62Ae0/pfdQEqMgkWqmZntyBGr+P4TFUDRBz3MuXy
/U278w1k9AdiUHzBKt0K9OKWJWY/rnS8IA7jS076/1+2rm3sWBE3iFPnbaXZ
0spBOf3OC2BaHTwL3ywa2NjDXYe6mPHVmaeffX5DlPqDOK1SddQepFwA9Wi+
M2c8wb+ZnDSUkIrU6L8K1FGbsD/1VFtuENbtpjhQzcQvgMmFVaizXGEv2wN6
M69NhDrAKb4gLrD4/1ft9mnuVGojmMKDEbs5WxyRi0oT6O7VyOQ5pqU2gPgg
nKNmX/7MNm3vs2xKoULC9hc3SiivPCK2xwV9XLxrz3EY/M9VY+UMoUc43yNL
KaLHr+g5VGPb3JYQdgoNkeNaU2zva9fSAqHMn9M8Zi6egIvlZKSoC6OQHfzG
MXjfbcz4WPwzZwOm7B/ZecQ2Qm8zUUga4KRNHXWCGpnSIc/Jn8g+QHP3KTmr
ZTBlZHZDBRtdPfAEx2lO11n/GGw84GBb1H3FsgTrQ9BsHZbSIiVq39yVLFBV
27vQEjP/60UjEL4J9/10q6va4I0ISd2qfyF3EeVrXs7/KiWSMe4UFBL4OwiY
+4AlUX3RN4tZhAh6xo7c18M5H/uWRLyXFyj0XPKSiLoiwo8/DASpOTpl2K2b
SYXKrCOJyWe1KHUOqWbPv/xlrJ1i/9/8X+B7vHCcr4YYqjFamfVggGKIqAX5
ICr2yi7wXlVli0j+ZuvzSdJnQyhPwMqVepGdmmT1/buqUeGSqPp0QIXHoZ2F
C0a2vTNs4pQREZcqEggMzQypxHSuguv+KgvsNI7qmvzi7hFj+x99QpNumeRq
vz0LYCtwAtYkN/TB9eiyFBz0gcSQaNZn+NREL7ifcbuoRP620g2A3gZ9qLbZ
ax5NtxuyEFdNEH28y+An/ldUcV4YM1T0omqEyJTibgnnpdTNO2DVXj+oIyze
88gkE/3OhRvdDOYLGEQGElDfFg0CvfHhauawidty78PB0/b883t4C8gU5lU8
euM1D89dMoZbU99FfnxvscOIXoxcNE56hxpDNLRGprefEo/NPrZjDM0//f+1
pOEPHmiNn463riGOiJubTAWW1YtgtbYVrpPG1dmAsaNEMWbBR0ImxVeENImw
X/WOulvJY8X4q6LwunatPOomfQqY6mS5QPPWqbOu+sVm9ueE3NLvewVxz7x5
TFp1Z9q+gj41bhLiNJB/lN5ft4sKhTRCBCNcwYpZM7FYbKbo5AalTtF3LeSH
utj5WW6dZjo70SgV+xZAbJ2QpmHwT0YHmprNCTz1yHO/rxuBtn234Z9c7ZUm
bKTYxcgWnELhy0MK4Vimw38lRg1aOPmzXk+MKG+Hh2hYsOsUzcwq60O+qyrw
u+P9nRH8HoDTfcUjL4euJmPCsPF8gidrQspDrkEuiMDIKZH2I2LAyxXORASw
PvKIeGvXG92389o+S7YviZm7Rr6nKSG3gKcFNi7Xp1axz5idQ+/c8l2IbYV1
uxUY+YdoZOmfaCO28omr7Wd5N7DTEJI1ghI2GqpUvc7k6it/lq7AMDmCnctp
XAyZIVa3YevBV5Txic6n+ftvHOOYQaOwIvJX8FgcorMAjA0QVO5PWVPUULAf
XkifTkD3s3dltazVlL8KNdEzFqltZvN/VxqLVTOrKeessGgAlojBjjffHI7S
L2u98SNUSXl2kL8/Y9JVvTM/IxKA+x8F3fYJohoulI2GRXRGR5Hn/H8xnfOg
PZeY/iKgsZED7FSxKrYpoY74h9sMOdTEHJRaHefEqW5U5h04lxO7KipGdSrL
sVnX6fBHn20OZfdY3Hgb9xo2LPy/KVY/P1yG+NwFhbI6VmfvGJzr1Q1cjzGk
xwVchknGwLT3I65p5n4RfcSPrdbzSYcjIY/CoxQCKGMOgzBPn5TyvhgSgmF1
VXiS6kPnBJ6lp1Jjy9V5Eqz34L8kFaJ5LeoInby4swnC78K27EMwipA9dYm5
O4T6HoUg8ea8u8QlpZlS9kmif0IbmYq028L/uTI/2lYmgTRC6yFY1wqIMs21
r1es/LiXVmELHfZEkJA6pE49m3hUIAQng8G2XaJ7NNB/4aum34KA+goV8Pk7
cvRARpcuKRegxfBK/5t37TqRsX9aj5mAhutnhS0KUiQ2pHMACkS6UVlca7sm
9SCRxiX+plv1uHPNvY7WTBu52L8rwb5SsWILuiANroxUnb/ttxWz6A1JEoJ2
WuPr1naS84noeF+JvVec9SrQUiovM3227Vw1RWhE7JizA7je1x7pFKo6fwwd
/u7pQKtueaKwyr/I5I5FjxI9adeEp8HbgR/6ii4tQeLyYFutWfxck113hRQ8
TSzaBqk+iq15gr/2pvjJOGebrAO7o9am29L275dTartgPqxBbw80lRhc91yU
L5+9fMrP+wB9kuWB8Of3h/utGZ0voejFh3evg9LBI+IgrIUsIM8wZSet1gEr
BgiwapmFbBX3JTS+aG/XkLGrb1RvTjeO8ccyZbHKzeI0CGC3gWzaF8oapwJy
CxuFiS5tv+pqmxj6By/nGvaJ+4Mp4XOgP4CRQqguww1rxqWDn1058Jrzcs3s
3PNhP68ER/kRftXf6CMKv0OQ44YAs4WikUUy9sFsTOwF6J4n0yXIcYbxN4bh
gEATwUJPZUdJ0aSPSXUL92IYY12hmhjbaF4/Aq6WSWeF/wEO34gYJmgwXXAu
2CSGuUtl4HS/JJ3JOzzyNNF+qwCnf0aIf4wZTxE1VuBw+ZZy1jUA1s1wzQbl
7IPFg0Gr+ruibWT32AV9WmpOLVJ4pJdbrZUReq3+BTj4V4flURncLeHtJILb
sPqzAAd4YdjJkQ+q7HZtd6EwuechIvTunhPVGpvo7vycJ2sreiJ3/ihmJ7OJ
EPz9rceMZSmyOouJnN5lcw6pbRIrl88XnB+LquZEB3cgVPvXdzsMp/8KhyBX
ZLWg6/FsJVplxsrkcbZ92Ec+iRM6zN2rsaoet7mPDmebYr28RI/6e+Fn+X6H
N0QS+CMF70WB0OdxCUDNsoOR7C+l8tdu4qxGR7jLlh6BvJQA3useY9mELVra
9z6cO7NlMCZNdhBXNuBGpKrh1BRrlPzWzEMaqlS67Hv3P2tz7RhqlKqqEgkp
oUJNAjBd5fuEktLiFhx41Dl4C360wQmsRlHThqrsijZWEsQV4/kMGmTKP/Uy
KmnKKFbcB2OsmSTIbcdh2afXl+ed0DntVDhag40dGStzgV7d9AAkVV+LW3+s
zH37g5Dq18B1OO9CU3rAqHxuDTX6p+QeTgAfTRxfRq5hMMIaOkUA9R/ETNY/
aiMWWLUX3ZCDJtaT3yVvj1GSQew5SqlJeGaRuosrPJFfrzb494IgkeKtjq11
igWN4UJgghYKPU+cN+MNMY+i0oVpSJ5b/WuNxfEE+e0zc5nS1mWDRZHhTJ8X
KiPnbTLN5Fsk0D0nudJbu38b4GbLD0ZGezwmKZ7/rtbSlWHfU0Ko4RC/Ek6s
xPvoxk6vbnkz5R2i8lCG98s/etABLAr2V5iQeC9GuwmuvVUOYPBN0hoRnqd+
5PMo2y4Yr/18MOKtzLjbOLngthAWrvhtwWmXs5YG4XHvlao2WbkAlpZrtRH+
E7dOiAFIM7Y4FckUoT8b0isIJKTKwvjSUHgueBwHz/m/z+2N184SterFLSib
Z6vZFzfCYScKfXeblXZFgZgvVF8ohSGrh8spgrJrZYGw6YERo+yZA3+4alge
AMz6h62CZJvwIYbGWwHU57bD6biWRiCUd5moFf7XYKWOVrGm8WNoM5P1XoU5
8kXKVXspWwUoLB8pD0evKViovWdpL+umt7pvOkMcILia73GQlbpKM+CEz+n+
ScBxwGUp3Zyprxfwk7yA6tKQak048pfJfAV8kMuNhlyleyJWHTBGW8VU5Nhw
bGZK66wTKguGWDV8ng9FIVPbu3XB2TPoUX8+cMsMd6XonpZZQj7NJrH43jcT
vQ7TM1nOD/sYhODjMJcNIgWhDsp/pnpUjhipWZETxiyK3qOtBeFBZ3Vno3La
yqLBP6KEifzn8cWgUWSvFHGiNCYMp+0HTC4qUXBtkmG9fifCbGXaFhzbQJ7B
uVO2Tgxt1S78ymPVgzvdftZTMBZrOl+C+FH/mGlHEQaTFUtfNmdu/G+lXkd+
jeQ5CUWED4ttpQ1vcWb79ztkYba+CXP5IP/Fp+ZeDdCUuzGjILd7yHwN3ed3
5DyIDGyL01dpY1FXSdIBN2HBGPzUDGKDtKUVkb7lvFMJCb1JyIRIncr2tjMn
OLXl8Dr29NLFYQYeJMtbY2UDZ+ygcy0T/nlGFGdqEbuOScWumUR4KXjahU5A
dqqIy5+B1naEmAAD8Cg143xDBCKWM8SS35FrelJVwk4bxvGWAkm/2kTclY59
Su5p43qnltBJm0I3SHgQiKeL7bOq4qd5pds+2qBnZYTyZNecCh1/fuqSsksq
Q8N7bjr61jowSk1WR+43rQ8u08qPMsGPHZ6gbhGKSHIev1PZeZq2eOU5lbVb
VBBlA9uSyyUE464MihOj6hXqoS1S3PFPgzDTIzZo0U0YC6OczwxyHyGlxcnF
7sj6krNVoLFNCH0M+MW7zplNejg+e6Fs4pXriTUh8uux8l8pSWh6g5ahhO0x
Jybcf86kDrfVDyK3W2ksCy1X3MC00gJtqv+OwSMIS6ywBftkrAxTwVgxRCDk
E+vCo76+Y65SNRHcuPFTfA0jnNYC6mdrdu6q8UhT2BrK5b7u87FiEsbxS+YC
E6dMwtdQkQGD4yaomoOLn9thE7idKJRXwqhHS2UYsQbpvB8UlJe8HESbYTcS
0WIcHCkQUd0/0qxpS+uBIkz5RfJStmipbtXNLX0FTMcoFQzvVICVrSCmTUTs
mRdQoRA9K/WnQmO/Iaph3e6VCBKDRqeG8SbtarBNZG1jLEeQwtLt9niZroJc
H8XO1TSb+31qZqBMwdIbvu1q6nEjg4o4DGFlE5YpTVy+4sQG9MNPzY4B9knk
JmAAJFW18XgjzZK5i+EyAFoFBVyth4Q9SatsdN9iMGK8GvRnyXiuDinqvh3w
SRm3Rz0RQZt9tuSdlelkPUpBBouCAYssm7B5eGIcLr//obhnE1eC3k7Bcg9s
a3hwqHBKUcaRuTFNEb0UD4jPmymECKWRSvnOMiXM7URtx2YxFh1HZBXtrkQr
MFp/M3lUlA3qTQYV83X8xKlAJwR2yQ10X7IQoj33krXliEQki3vcWmsAMt4F
1UVvfbwRAohZIFRLs1uyVEF2GTEa1BHKU2Ucva07IIyHW/QoicUQxY9CFyiE
m1CW2c6HFr2BSB8OHJFVtH5X6Pf4PaSisLU0+KDaO769Rkgq0K7Q2OpHmSyy
/bIHicCSbhprG641uo7r9OuLydm1VWrR9C/PDum31Tf2zwu5I3FpjHAap1VK
6+cFDircxuroIDPXMj25zEVAJ6pCkbfF2rjMxG8RhsaZKpLMwv+fl30kO0D/
i4cSlANVpt6RrMqEtHD7EAEBtRpgI2jVXmCWioI5sBe6vodjspx5J3Kh7ZRT
xOvb/3oJizipMlM0wskNZn4J8K8sayiEYBx+O01yY8mCMZQalafbP6+eCuBn
aczsMoAsHya+JiiAlE6PgvN90UL8Gh5ExqEqqGT1gTq/l1qwOVd9i/Ugao58
4B0sr1BJGQYDubVz4D2jv0AivY6qiNGYumtH+Eezxr+PLJHTUoVCveq5Ql41
SBRgYPqnmWWRWyTFBeq26uT5e8E3VsUNtk0zIJuChqCbkH8txI0Wg9rumLqZ
rSJBj+a4x3DjiUKZyJHgSelh5Br9Tg6hLeSBDI8eWYAHok8wcC2MHwrJhV7V
84nBwkiMvAj4AUOh/MXj5fVr7rO1WkaVsGbRMi3JQp3Ybv3VmH56t3Y3dLtQ
JfIuKLqm8INOCSSNmq920MX1caY0SWF/DzlOBTk8OVw9MQCk4JFVfyHrVFOt
0Z05/iyAs2yxA1UPXxv3bve/LskxeV6pp7sLiE0cNCiffwF40IxdIdqlgQ53
A4MMCdg8VEFPTXtSuTv1YvassD6GqfpHL8WmuXR5NGQ5chFoU0QtcqMMPlnx
oU0GrHbH+dHd3I36CcZH86L5YBJJ7Hzwufa3oReytUZpiIRbJl7mfbDZ9YKO
klVVmPwXs4/gs0skB1cLiWAzjarn/VOHXf1mB1pLbpU51FEdFWExvi281kcD
nLzRbASbFdqDX/gXNEhxrgLvUqLt00XWJ9aJs1C3FG1HRTv36+SssJSpV37t
xBHRwbmd9/TgXXoREHdPFmKeHkkB8+GswGpOk1RctBV0bcerkYjN6eyPt8dd
81Eb0U/SxJVcD1xgSsaJP5VHBwW5C2Y5q7/6i3zG/WtGEIe+k+5ANEm6Aiwo
WvOITWw1G28vlT5K8qxZ6kUipMovPssQanXU/Tb4d4GRkuGCZiTU3q7MJo07
t0yr1bDZIyToa0qOT3E5BLqos65zXCo8YYmiQvaUJR1u5dtmsCrf4kuugZbE
pbVOcsdmS8lzG/waAFskxb13J9vgWZZ34vYtNKWrsVa3pyGops/R6pRmBvqj
rnQuqMwoaIlLyJG7h8FdoJGww7/M1+gIVkVjtUfX3fKKq5GPZjK+x2HQ60/a
wNC10ahjk5fwmkdxKzDqO5MWaKPHZeW22s2LMLbLSuclzSwxNjBpq+Y4zG0+
zdopr+XE0WTfMtO9Nc7TkNEXCAMb2bUJMf/RWoyq0jNCeACtck72Rme3Wc8R
BZpFe5Uidx4z71bTO/iVwMReDmWJPWAKoSp8mLBNu69Rumw60W/xB669FTOp
FK31oHU3khF4sDb2fa/CYgVxzMQ8qNRbbzkS1WqNLzvXeDenvKD64jCB7NZD
1H5tZAX0KEUFKZEu3jYzBJEyNn8vK6aJ9+vLjwFc82q6l63jaRmEuJVa2fla
0InwG/Y4ALyk4BdpwJX0J9HIkXa4od8e5l1kWsFXgOw7eU3DQKTEXntNTh1K
N/FrKrWRU5fmRXmjLrPqS843N0lbcUi9cRUHApb3FBwEAoxRXERUUcYmCEhp
6+AulmV9+ZeC7+m8+egXCaHiXJwLY7O/5N1oDzpZTauvhEo26do2p4MBsaJQ
Qoy05GhxwuaRZulx6NBcolTAJPMcSqJOLF+j7csi+BD6Uio2hP4vOjtVn7nQ
XD5mgIFuaBMSm06erbEXnd99qFxr1cmmSQyz8emmqKNR4bmFsM+zdqc943ss
rawNgaXSbV49IGn+pxMdhXovA8+txT1Fda0gnQCQVhPfF3NT/l6ljPdbvpbx
6AIi+8EipJZ8jt1PFfQ42iFjWydQIJalA7bOsxo1Q68MNgrA3KhYW5nXS4Z5
ellwoU6cQVDbTL8IQFlfDZJ6lZIkH9L5Oo6MkgKH5JVdXNejSFunUJuaOOJ1
SUTTST2h0PKQwg10Ch9aQnAdAZ/8QA6aG/7IJIMpItyzP3QDLg4NDkUSDrx+
rcfOLOPl/afstX5OFkpzMsYcu0OCC5Eu+zvoKZiWBxCHP2Gh9+QfIG/pnsZQ
qru9ZMBy4rAgNPwSvb88msO9qPAIolat+wvOgZ0/i0TPyQycyHMJ1n3vbkdQ
gEFKUSgE44kuMHOlUdyOoh87A3/PWDDYQhwvpwKQGzynSWM9R2giZbeTgNmv
IhIj7iN2ABkke2K7dLv8DUAn9Vvg0ILxGAjLQDtzxyGvg8tZdcxzOZgicY4d
24IH/JQkX1dffGPGw5gE7vlLevpf0ClHjypeFV1ZMDX+cvve+ZgqcSkKL3uG
Fu4Lt4rS7m5n/1LBOF6r+7Kw9zYlNG6sO72XxM+OWOKbEs3EeAiQtbEtJ9wU
hLVWgqpWLLxAJxVDeu3y65BDAzw8jJUwxdMLlG/zDr4YchiY0FLB/xgitPp4
NDl/FLt8cS9o4gUtcOokBp+7BuSvlqgqiYf0qT71apo/Y+KyEkZmLtbTb+0j
wC/tOtSC4diMRZ+EOwafmf5tE/s6H426lT4cjNixWJlcxBROqzM7PVcjxMGi
YyEK6W5NPTIf0xtafd7OSLgwMpts2g/BHx+qKHvSYXHoC8Fs4OJXttFX/O+l
DKaKEluaNpdupc8QfwPwbMEPlnclMavMpUQpE6DdHAvHVB8z2Yv0NxolcIbQ
gW04fByt4ecZo3RN0TrYFHrtjxoI22aSk33z2oNqo8C72wdHhoh0ZbtdBJnV
XK7yYhTHzND3yanh3ubvtpeevJh66AQZOxFiHxnmG3ZbeuvnknOjo/X7LdKF
wgfFdiLgALIWyt6cDIu/FnSHLpC+utzZsyxrOr8Z3w12b2Rn7q1MN+1Y5Bdv
HEsFNZkHQluINJ2QFE8dTLeWmcjG589ZVyP8t3dIpYH1n/7WI/PZEMDlRR1/
1RiDUkr0jj2jThurnJ1xiK8fp6KG6qgcW/jZdauwUhIB7wubf6nXR6ffPlnE
sYen4Qt8dZZJiXKaJt/c19D6b/Xuw7YE8UkJrfiQ5N4D+5OPwqdQ1EiyQpQL
KLNEiUVvhPRHllD5f/M5l1pSBido+JW2vWqQR7ZKpYpgiS8LeLnoxTas4+bk
LbkiE+H1NfDtm82+4JdebEFVtsRX7GTbHwFfQ//Vw45itJWiGnQYqgv7FJJh
0oCN3Bfl0c7WLqfN0oYPnQM4bh4Dyhrb0LZjlCuvunvBB8Tz5nOC1/xKgzig
CYdjLF9m0c4PrtoU+izKSeME5g0c95wKQp+oDd33sJa0sXCLJWcOK+8BRVIE
T3C4Stwj6DMh+Hznd1JQbPS8pZx9OqbMOBS+d+mB3grJSJZbYCFsNfPK7jlv
X3dIRIKe8U0Fz/TqErjsANZ7MJQY91vw8DbaksXqUsD4pF2LaHATsq2w2DWP
e+1kzpRBkhkB7ejj6n8bx7k/CD7Lmgvj9vXuv6BX6mnOTUbs+BvF3e/fIE8K
WXjxJ4LYy6bjS7XaW5/lWA2r7GMZkMYRYEx7wPjekmdIMS/gAugQ8Zd77xa1
az7lReycEQYWi40X6/GbKZDHAjIzwJ5V4CiFHnhckBksKMyMPUNMjP7Gujnl
WuNPb7oQQykRVK6ohbooja2TK65o9wx924SpEJLb1I1JWKazbKdOO9SOBYNZ
V87vwLsSfxhXAlc/3ob5iy4iveKIsDuMUAwaiOM8/w+WdWAluulTYX7kzbNh
R3uqKQ9ddZeiJupm+wRl5awe8puAQNkXqKImtxcFGl1CoWJgIIlZVULi4U82
xudC6gYCBn9LHEL7txQlOAZhkJ7PZgt8ZP84UlP+LtdmkZEqiC66VpTRVjhr
9yD96sMJNXsfB/5ElHbjRHz4vJ+KQIWisZwTKQW7Q7SusG7Hgszz0SnJlJBG
DsbBAQrwNKnaH6slola3Tp09VenBevJGZR1wzga84+okqvzTTKhgDa2jPyw9
QEUeno9laoD6Ts9qcOKcOyWwYNHv+6kVfM2uHtLd+26O0uQeA+XG0EjmjZ8b
w4NouVovZbf2wRPKcR1tAmSObAZKWpWzB5FJ9ZsJ+OWzLalheXATb94erN/h
7vyk51VfhN/902x/avSXq492CB2omx85wVf8eIcdglcxQOivtD0FAJbR/sm4
augiGbfZb07JxXsg3XmE6TejLsHzqp58tIM7r9JpWZbrdYfAojddHLjbKSUq
U3ToUfSklhSlfBCt+FxGsWrSrZJYpWHiEAAVGAjvdzSL0T0Fy1DHO8H9+GO3
rbshCWcdZ5enkK+GkfzuT+LX7UOBNsxFKIDu1ucC5e+6mUX8BUg2au4e1Nuv
97urTJo8MlK+ruiNIqmyE3nQ3D5bYwgoTpGnCqST8bYGHv/LUCJ64qMD5yfY
Af7QtUUHhxpO0goi7xZ7BrD7Fe9VC+V143Au0B8Uy1UPfnnX6L7hJ2XiRWhJ
zaA2gQsmxDlHkMl0QxKva1H5te7d6H/tJS835GEl23ojtWHEffuxyM2Q1pXY
0pboqcCX6pafeiIED+AaOpM8g6asKbF5nKTYU+Fndv8an4RmO+PIsNozOCOF
ZPd/tdbnyYux+Syw8odpPBaU7MKzSpwiEvfHmAdg/NTgn5wlqB39HF6DFVbs
zGVoK6vCfj9NJWyxytJVbgrRkeUsctp0DmVZ+NjCUmr92dSBs6xFFCTsmbcH
f8DQ2d0LvNxDHhMuXaHKNUANvEEcFTMXmyX+ejdx8GJC9mYGHv3AIzvBOvBr
S1y8s7wQd3LOBrHk1jzdQaOuhFIUsYooY/a3ejfaxoJoOjw1Mlv79lEbKXhN
3gOQZYZk46uKWPk/rX/U4ustolz5wf762/O+a93GflSXZDjW0yJRJq/r9JPr
sR/AexSPWoDjJg1uUaUJB79/Wy4TxvVRSVsmR5Fy/R72pUbHWexG/E1BfOvX
VhoDFokOMKMOwzpBYdrIzlDtVtMzmji6YJx82Oe2huYXWajGGDX6B9t/1K5t
AneBzPMyVNB0QQXqoflD9gGFDEGpeJa7qQcROVTQtLDcAhXygyzSh8GeP+SW
UKCzeMoLFpLSS+i7tyFImt9IZkOLgZ0wi+RVV3+0zfcolctHYgpFDcPUoZkm
3svBIc7P9REFGrkPaSqryx9RFzV40DeQY+AbB6DICF1om7bPoa0HgxV/+IFQ
xK7V703wG6K9JJiBxl7aghvZMJtpzavNWsrZTzV5nnVta0+ADGAFTXVumcWU
8u2dVzbspm9qKwPmbSIVzESfTXnuubRZ+VQB18E8fWlSRNw0W0udR6n934Vn
idZwsCq7u5yggLPmEx/AUofxH5TMo2uxphZgEokNA2y01y+dURPHgWXUfb42
MR2X4lB/NUTPIo/p6Rabq1ZEhoHrwvbe5NYbSD3PCm4VcfqJ0Poo3gigDf8L
mkoMfZezuT0pe1sOMh7F7ko/67iqFVC6oLEw8TtUvlySVzU+0PXGjuaSFIya
xQPKu/DfSen20RMFmG590c6q38KpwoECzhJGbd4jGy2dzi91PyHV7eGhUy9F
Y+ERlqvkQ0qBvq4i9UMDhc2WbLiCjyddo0VY14icGrYJhvxxbUwzDnVEv5cX
0Ga5zJ9HYDFCwn7gCkerZwYuc28BAqo0X/OGjflblQ1xb9q6j4vEyMyy5PML
isKvAIUzBdXvMUFn0EsHvtcgEULr8OM+IrGMg8zMvKfTewqX5WnSWq7gqlDi
CA6yKXOSx47rnuQEBICAht0tc3UahApIxuNuVDIDWq2kRXW+CDOsG4A5e5gX
xCVJ7Vhe+QEMgWCIo8VLX2ik/kndJ/ZQG5rLO1rUlAwlhQq6CeWlcg6nXo3H
zyzFkIJx5LUoK9E26X/pI726h4a2B6Wu+//3iH9igE0dVrfOeZbVMudUOwhN
H5gmR79ZnAgEecnfBHD6m58jQtJ9SgQkpQH/owIHEsAdYMOmexPwnhqOHHFV
uj3TzaKmWU/q96Z7sDQoCe8/7oyj96UmqCveapDe5Xs0ExpGEJSgSHXqNHs3
I5Oep849pxM+RcpNSsoUTdQhSTGdXBJ8iO+NbQjbVZ2dQ6QSZJtf6D6d900O
cTwPfRLirmAZOylNtYTibcl4/7n7psWerSRD8cEFd4m/FYArJcFt0upwdfR9
dpKHLPvWP70/gqqELEdOZfKEVOFO5kI09H3dMwM7xFFL/8V9F4yO/FvnFeDe
PS0wN0TQ0SUAg6xmNiAZiY9WI2Wtp1Fh0W5JjM4mSIfIapPkE39Sqy4V1D0U
bQer/LeEPyAym8I/wsopWOUy/K6ug9nFyKs1QubWTg2H65FcomO3gNKaVtsR
evUIhAxGh4IglkF3m+Ra0Ik3mnqGUvjSL7qls3QdqYzSHHz63kly8HO9RqL2
Hb/ze3wcfs0QWO/UGgwWPRA4T1q2vH3bMh5NXIc/B/YuC085WxkFngsVgXmS
lFVumGg+g60+L3rM3mfbVAXhdnLlLNNSq0ehjBTiWxxAfUBCCbp3AALr+6UF
KFKon3T32kKbegfn92WjfTM+szwxqIrH9/QkndYaNkfAH7m1ClR7A4gts7up
elBkeIZV90a1akWsG43q/k4l1QHUW2oJpT7z1DKbJYmzw2mhtcnqejuAw3ZP
QaLM2Ep9h2zrHJJxe31WGiFMxJKoW92yhteGMm+IA42KYB2BwVVTGeZvQlS/
scyRUTHycZoCPxZymAW3/emodrzkTpa8BuWkszgZHWSoqMSJVluVQi/lVkyQ
ZBL2ahxBp2tRS9QijIdFUa/q6Psv+5HnBex45Gx+p8jZhiiOgfcrEx64EUV5
IbMwXA5vfjTZGb3i3ay2ezsrWjBVcqk1wIUF7/32nYYVjMMqJcpX3h4Ax+lw
5Opcx0Ya/r1JCafdKOlyB3suRm3EBYBruj8qa5bL6RwMjxPYpGLjc0qL/oto
zZ4gzYHS5M7BxsUfrlsjyQ4BmFAeuXHJ9frXM0BDzeIfDYKoT1TfvOclzKdZ
scaIDGSZsAeh7TRU1RnvJyEqO2iiYuhHAtnd0L3PwuG1QEZyuubSOQs37iLn
TeoSKHCdmwE7MTpLTqNvycloGyyXnRHNYucz5FNCneoM4WTAvh2pM1Vhlzr1
I20oABqDNA3auRtdwtfwGUgMMvbOyRqM+KjxdrlRrJM43pgWvp4y76G2OAlk
j5UOAIRh0XcMF4PgqxWQ5XuG4s3aZgSFPky2VVUSPVbzJxMoicsBu1mbm/I6
4UiPE9aK9xv3uKC4PBCXQ5hy8q0hkC1/zK9xTi36IDm/xMYddrDeSrdmNUsb
KsxTPGEjMbmJnRNruqu42h+08HWYbYYt715mxg+vlQEvIoCUd0tGn/dq3kjM
20qWtn5ihPqCFeKnAVT5wLx5dk/IsGgAUkCCxIIvY/07zv4R9eIY0rdywqBU
GcZzVyH0zUaEvLHX6Whf/R323W/BO1agUcpL3gQ90OTnT28wmN/3GoILl+hn
SRui8KnUxqIk57UYnilKA2Z41HKX+GBHyFY4YIZE1a584rLj4IZdaICjJb5O
16o1ODi5rRJhQYo8GNxwGg9+fyLHQ6LLRNcU3oGNC0v9I08L+sSTK8i1Ux3G
ti4Wjw1JL6hBEPhSrMCofL2SsLhke9NCT8mp21ZrBSTk7u83hwcN5sjfnuSA
k6qPNjCXEAYkjZMAcBQSH58Te2sN4be1e3+UczRvZFAraX3T5QQrcsPW10FP
w3/oqiZpcgDFApNHf/iiqjBWip300HJC/b7RXra0CtZhKmoDc7EAg4nDqrJH
PHvWoqXeDTxpqz7m5b2QbmBi/CLH7DQq9v6Vm5OkX9VfJC9u4vE/S1VmD81s
m3TmLdolRZGF8lmUwoEO4RcgDT5RA8WP0G39q8VnPjAfLWFVi4rqjJAW4jxC
7R5jpHEkG7YfdXcQfcUVuq3dng/6yYdDllaJa181zPyRe+GQL4z0Q13Dc69H
hxk+3y4+VMm0kR3OAnueLhkwOpR8WWNmr3wo20rVzKCgqNKygpn6aWIpyn+h
ATnOYJJSvZAdGwGwdyY0IeWHzXFcQqF84G8Ua64XBs6lwcunEfrn/Z8HPHak
NbYzCdZrXTP+n1jJPB6shltNMv9Jc2jAE5tIU3tp6xbFl7UzpjUSV+82QPYp
ycsptViBmx7L1ALSCUG0lEJO79BLJEsQJu/qC6ljo4oR5uxLrYX0dr278w1K
4OQ553pLbX6gdHwWF3DHrFswtI6kQpMO3Bt4V3UIvnH65glcqyd4oYo+E+pb
ODQ5of0GsLDF1vZNTo2Yh+y5bnEU+aQ367Cru6t9+SpRiro2r68Y8ivhxxx/
1iY2qvpL52a6TS5EKHLWOuYX9ZNbq/krlmWS9God2RxDJMjHt3Kak1zvYfNw
lM15LBGAPuJQhbCyMbaSwrnMxoP1fQFzlCQ2GdE2mNVKv7ue8dlG/yvopShV
e+hPKGgmER4hSRztaHn0D0vy12E603X60KMwJBPH4HWPUOHOL1KK+J4KvmqP
Duif7mtmiWMK20M+FFH8pmSycf9JOEFSLBDAkFAW3esU4d/cyBkfb8qrVDYi
YtbBChsQi5ZW96VHQHSSasw2WU5EXg/FgkNeqy1SR0ASQvjjJbDUCZ8UXyjp
d4RtlYwq1P3YKpCmJpR+JwnPEZz7lIjAqZ+TwgYOFkKOH3IH9xtILbybWy2U
TLS9KEZV0vFpHKIPp1VZcz4dQWmZWVBoTJIMp2GdbnstwMpgFPtyTopokZum
3xDmh9Vpwimr+UOt2X34+UNnnvVQ2F1+2xfXyFi4ekL3V0VSXJJW8EyM+nYa
qmEMbWVnF0wHF2Dc6dZnHAFqcvZlFoho9D4BPQaaL8qskLWgCBm0cY2IQYv6
RSYSfKalJS0qMc9dnUPE/7tbKEv1t9+x7JbSZ8hHt8k07dlKy+woFWqWAZzD
9XL88iG+HiwiG5m39AK1r82PNCIBqqw0SyNuLudHcxwCG6fmEyDyNNO33cd3
ZtPZHPoWhheGI9hdoB1nzu6cVFW36ETuYyUGd1v3GiLdHvBIN/y0TNKmilxM
YThUu/RkPKGT8TvUFsTcEap2aM7ulprIPkl1ujiHtH9GXx+9I8SaL8jtfsFR
pXIGV30Mbjt3p4Vjyje2aswQllFId5bss6BJSrtZmItPQ8GSSMY101YIg5L6
qXyw1bOZVwb4CgQoBrL4AxtVKEje9xoBuTNICibt8mtK8air7V9QTicyRH3N
1AATwrkxLhm/qNcCsCQzcKQTwhurL3y4eSOA4XNOUDhsBr39O4Lb+LrM49di
NxyiXU0bzLVe6nQImfKZEmFn0ikRJI5LEqEVbccpzzRN2d788uuG8w+mtZbI
lBaKNlD8RhFYrSUW/YTLEl7FRL75hvHGviGQWVMJgE0G914x9ssdfqJt6PcR
F0X66QoxCOIve9p7g9F4qQT4WWTw2TtHaiLBTVjVqyKh4o7L7BV9tjoZnRXR
aHcGrBToNhBmbbPaiMmynIuGdt5Ud0BMlbJyxaufQr7c93CclnfeArlwglrz
Z6K1iI2sLkkDh+HWYEQTxJjSPSq6GIKZaJqgPhItkdt1GgI2qV1sjydkHXSG
+FBgVVWcmlRJL6ioWXSRBdN6oQKjTxT6kpN3YCgdMfVSNquDZxzb03bP3yfk
ItP/BsoSdUUWj7kQQeaTrTi8JGNEh7ImGSQMxD3cD/SGvJWZsOz7upET7Eba
+fZdsL0OXniJLLIjw9oRzMpvYzCuL7hnL78z5OpLCOeGjw2QZStlKauuy711
1eQ3gPyfRvLd8qPis88X0ZkmfhmF1gTjQWXZ0lfuGNAtTmIl2yTPPzKAK8hR
0sNFgdfZBdLWbasKY05QFAz2y/llSxxETi3N3KDsiQ5KgvN+Axsor6XgLbqf
F9jMM9g0hIFhLwut1PSGbXyatRv5c5L/elT7+hfnXdZQy6lHkvwqi8N+vOKE
6/clwtEaOVhMncrdO+rA7G820YE0aAmo7quzfcQg8YUS9Ef8Mr8XrFE1soHx
fksq/5Nohs9cdvDvy1Xxc8KrDAj4oBYZi+HB2dyf1/kO7WodlpuMueqeaTtM
UX6dsTN/Ph6OcLJ7nwn2q1RmQV2GZ1aoth2xWLGsSAoUo64mEAGgDr9mvvRn
EXlDs15BrmM7xTQvOhq3GgrTPvGOxMj1BlqhQk+ImcNYVA7LGuZnmkoG9me9
C9udx+q3GUZAbSxyyn082bhfOiFN/xzx47STsprczjeP/cFIMfB8+T8Gxczs
sIb4fuiRnyIzibefenaop1nWGN13npPQMPshdKc++8JlWgZUAO2P531Ye/jQ
zZu/oLq5kqloP2i7hjL4ErN0fgX1KI08y5CdJT3AwWLRd3gN6gyu9cELbfMC
JQhMcUoxSG7Y58Lj0BWp83IMEFGS6pr0DOXWHPPeP84jIQRpzxXcnRKLv1hq
mSTTmix+sdPUKyaCaepc9eoNLsm/GYF3BdToV5d8oqpXvBHMFVGpdpO3md/i
B55wA92apCzAfKpZ9sm2KZkExwhNFtXJ16qGR4V7/rNcGN/Wymh/x7tFTD7g
R70sGaxL+2s9ICRrU/d0j1fElCpCLW4y0fGT4zMo74H7zowABTOekHhZKeIh
WOBaJHdwP1BLj4nWdGW0EIv81nuCLtVdAryrZTypJX1X09qWvWX0blF8Gg0Z
+XQQOJxE5D6v6cw2Th6ZXufugLRVxMwQvj9oJnfw+6zY+xKK+7Qb1shVboQR
rZPVLNpfga0QwfjwjW5Wd3+Rb3ZJrTMo7YRBrzEIUiyNpakWYFEkVkUvHInq
v9HdypXPxdpNlHz4cDgAaBZTbnVDe+hbotWTu1De7zTJoh3Gd/Q+obXh5d1+
d+9CLjQ99QvZS6VPT/rRkONr+OC2tO5+TuChau8olHwWnAI/IVB5xn3vLMxm
mXpcTRfDwYhET+nt5oncrIOJ8vwKWGKkt0+YwusszPD9lrsdQlOsQVSN+i9s
U30oA2H+M8+G8fuVE/w7bG31FfUyut7FBxr8OaC+29NZpRuZOBxCknX9aSGp
sRDR2r2mG+4v5U0FH3N7E7Nh5aBt7ghSuLDArO57n6yMynwvpQYV68fsSYZJ
ZTSByu5ppi+BJzQxBi8vKNYwMJ8CROKdxybZhxeddsrVL+MBjMBoTXAq3WLK
1uiQzAAJy1pRwMUmCfnsPBdOG/V+IRYzqN8rlqMSFsmhZHSvKErZQC58bILV
fKd1AqZKNvBs8LqgYstO/27AOuDiGnfU0tu0nNII/t7sPgCtKZRUPlH0/4kL
cBnthdQ5FosaTpkd94k6nVTjQYdtecnQkXepqCBNBQbX8+gmBWOUGANvwJ9w
tUwzQrlTf577cXNxRp5Hx1LExRAqwoA6AmAMN6ZcnM+vjwTKO1FWdj36tG0G
y46S4V+9LaIUcFSuGFaiBKrvxhMT3LP9iXQPu/sKXUq1E2DCknAY1rJDSjYa
i6NgmfUEmLPZu8+YLxIWKZ4nx/u+x207uGZJSZJFwJtrDe02Fqi77ekM0abh
q+hOmyoHH3lsC7XmEjwCdlge6IM0K/MKfjJLUGeIHKzD/xti1UngsMx1xKNR
rZcAYa+1vYRj3X9Zmfu/8nMYnE47z6GiV5DjmETjuCpbZ/laqS8qwoxh2ZFm
Myxi1ZzLwJTsjtnwuIzu9buJxjrtQeXgPQPmcufFCHyiYj/ByJj85k5D7D/1
zyOjesyQT0onM0f1s84cMNIuI0PEFE4zNKdg6aBC1mmVgvz6/0M3fbz5oiJF
FOykz+kuABc7dgMwIKMmW5pmE2GgzWrqFBPtcDwna/iLql2WUjmC1u1hd33r
447AKwR03vfvUua/jPK9Zj2c26meg/osQAHEexKz27a6Wo4psgTqltOBsLhc
7ZPwJMZ+XiBmkO3aYWqi0JA4512lHzytMYyRDPwICAFB2iBM4SqySFvcSaVf
1Cm841kyD5AfzxmAfo+gTN8GX2ZsgWl6e/sFzhpCElVbfMWrrzt69KypNxTs
KXwHwseg9ivjQuEbErRnZah6qOV8HJyNjwTSU+223zHjltJ+8AvvwLR5lanX
otvHqGCE8FSd8t6uxOCPI+Ck/wJtAhuIRyzzmXBWCBt3yrOfJT3KgDLgVl9Z
cxTOg/ORv67K93icedcHdxABtHM9TgwZaFlHEw+jc+cVtj+8kxZttz+aAFqG
Tp50KHq0+HBCZfRGJje9Fqs88wVXFFerJuxLNO2bwlciDA18tD/NRILFpX6w
Fbj4o9b/1xNwqO67yTzCv4ko7HKoDs1xRkxShS4558KRPg7HK0EiXkr3TylL
6s9WGUCpGPAwXajjvH3Y44tk/e95aq+CUgx8622tJRx6UzQ5wTKowMc2TZEW
bGloFUKeegydcuTNPpL5cOMmanIiKpd6uTgPdYga9iY5B47A68uX+3sDvThK
CLfldEx5/kCALngXYy55PwuVM/DoJX6xUsZm/U+R7ZZpu2l1qarc67q4XKuL
nJUTKTPYRNavctA7ub8eB+UNtN0dWcmCg17jW2LDUzIqVeNYXDPNE4xco01N
1cLF3XXTHWD9BnYKS3JDq46m5d/ToQgGZSwtFCqxMPX3EPJT4iB+WVKk9FsX
dwY2TxxZoEoZHUKKfzF3MPsKM36fBsm4Z5oICY00Dq0CRm6KvJlMgwUCugks
vRdIzoggyc59qisyujqQCVhRWYUoaPp4GCVK+YWBFzJPBSyv9JNxlBbSbgyY
mc+z9jTC347BADDMS75QNOtDiB1zgDmyP2iJoWQFlPusI9Y/GCa/n9LpY2yt
oY5D9KI3lIWpmdo7B/buXgbtEf1obvogeJC5MEUdCKEvRmkfYr4TQOU3FgIR
buPKhzw1P9U0Fcev7V0YXs5cMKE9dRg6t7Ai47XP/gfBSZ9isIn+ICAQZjbs
2pGHVB9lTi/f7Dhqtzdl0f8qCxbWhOgrwWSQaQKQnFVmoK5ZJqJ5zSuzALtV
LDueRwoysIYAvISA1v91hjYNqkQbTgdRrKayHN4nyv2xlXrK9kDdHkhDutez
bxtg/MxRwBw53HNZYs2uOAL5OkxmoaSjMX2m1jh8Yh8pFzsX4Bu60TBWAkke
foLvxD/37dzptWHWehOT0yzvYLGjrH1dKcXPQE1xPA8bFKTJLadC6aUrB5Ul
INXHguzdUYwEPvSnU+R3J4pZiiEQV11E1yN+qsQy2c42GSMRrmmA9vn6Lhoq
1cbFPUd8Kjclu6pzqkmNgHAQRXwzzqvERsnyVmklNYSFHC6H9heDSNGU1PSw
sYQk69z5isDTMUb2KpDsDLsfoV1Uh5OAEMC2LmPt3jaIEKWO99xJ2jt+MUJ8
7IP8YV4CCbohmkcXJrwei0Gr8MyoAKKhyhcvS9njWd7bgq+OpMXmZEW7PrTh
nRaO9N0bdSSmy+Qft52cXIIXLeIkaOs0QXuCsbu25w1vsjjy2s5fxqi4cQ2E
+oDuTAcNiUoZUrLW5XqoxEgOOPztzj17l4cGPhrcTUnlHh/9B42VYltWkR57
0lJB6kpF0/XUsB3/+dwKvh+r2KQkebe0g9jsOMtwqXTxwTv5cn5P9oZTfNVS
zAYhPmJpYYRWv+/Ahk2U9GProFzYTijVPktrGw3fY/UTf9xmUKbgXTnofrF4
zKXC50r+891cE2DrGmVTrdWx6S9Dh0Xe6wlezFfqKKVORMmxrLRTV+bJxzkg
NGYPe6z5b3EHd6MU7QhAM0Mpvxl370RZXk5fR4DRJBeUbViNDkT+vrhwkiu1
A4EE/v+iPL48qaoXkAxTGwkPUruFUdpSq+Wwd9hKMRMm7z1y93GotsIgogIo
Av26UDg70GGoC/QsU4gX6L0j5NtGeT8Z2ozq5N4XW1xQUVe0GhaqeNKQJrwD
rL88s9vMD/SqwjiQ15foGC+il8RgsLULKisdlrk3FOAWJKwZR5mpdUy0wWRX
zmh0Rylkr6US5o1nXfAZK1mbND52dsXEOowabab7gPBtTA9TncBTy2QgMQbz
dycn7jMdMljyR0KYqTMZiGcSjZUeixkECjysl3pPH4H4U2qpKhCwO6WW1BIK
OvD9+1T7jlz9hXH03Hkdqrq4qF7C0XxiLR3vlS323YQV9vP4lIMWV3LORtM6
33ApgaVugvqnZQL7rsXDFnxy9irfb1Isa3hv2UogXN7lHpEvsIKgnskV3vNx
UllYo2sSSC9OHL+GWFsemZSPJ5LUFXHaU66eNDAr02AwhyGMpb8GGqdFoy4n
e4qMREtF7yc2/4rrwO7TfmRSaO5gLmhRoCIgfpZ+m/vnb9Oa74xIO7q3MheY
5YAhsozv3ouy0wCS0nGuWgjNaFDa6DM2p0RjLF5XkHfwvqkTbANR4iMY/rOq
9+GCjyv55YUa10IP+yO9gR8hbjpY9UgIlWxYqC3e3t8hDy8BlGjTmm+mkJ/y
FufjfEOK1abSWefaUj4gYclh/tgjt7sUDsz6xHPtA9k55Bq9QphSCGTFdJr9
ooPFlc5KWCQGVyB6jo/NJ0A5Q9RZK3lnKdeB8wp+hEGjc/nrwO2OGwThVFJf
Sy2OwbUfjTvFAXeLTu8T2+/1/7vWcZHqEWKFOwLhrNXW/pJajbrZMsoiuk7m
ibmg9coBHAkZmIEH88QyZGsrUYUeXOJPruswf+/VH2I6nv3+8ajdeeO6YuBW
HoJFtSiVRfF47LnbLkSXDtp5Lrk3sjPOneoL6QVZRMShUdsP79N0/asxGdya
Ze/pm8S7N2HAsOcNFiZvHhu/beq6JBC1GZ+F6v1F5LTN3M70KAtLU7LRrb8T
vd7Ss2u6BqUi4SZ0kHe/uLoJ8e5hjqnJ63jQH+HDurklt7RvSuQl5tD+l/Vm
VGPwyHIhgPBC0vIkkkmKbaM60FLG4v7LalCQQwzkfitQVbhondrg9g4yga/1
n4u9kgOKpzkPeCUJ5Kfnw6di0TTIOynxoWs6qvdParriLDDxadbGu9L6LGMI
rqP2i35VqspuN67SWWJbnwST5dmSBo6mSOojcjMNdDeVL6ax15fmnM6ZpwWe
izQHb+pPpxEf/OF3xyiSldRFe84agMS7EmtnK6XmZHuy+7d0orVfhNnBnOmw
SjoxMh16EllG9YcaA1l+uP/0OYgeygB+cqM/2MEpwStFQuzgC15msSSp1Md1
kdGOogBqHNeDQuaxdWW45G4ZRrwIADlT1RD3R6IJgVs+nB20i4FePs6QwQe+
wFX75/omtx4eaAqmcSkOAQSNJW3ol/eNWRF8s4z4HRyYkSZJVtjqT3f0h0Eg
wYIz9qqoCC0hc/oY5M87AJRzW81WmQl7VJyTElrno3y67E91TAVUYKlglvHz
Q9cNi2RGUkwHk6+k9KrP9yCRw0Uzgzfmz2A7yvrHIl4x1LrzLYCq98xWt1Ej
c/D/OKiAVu/tCe9rXKdngOYyaEuj0/5sbjGlIKCtQy04wGqHWq+TwuDWXZlf
m7PL9myGFFmUQ44KLrar5Q9l1DOONBlTboYRCcFJWpsyVg92jH2iXVzhbxhF
lkc4WwGM/xxnltovZF8ujUxzaIxQNzntOqhLSpiSysndj/dFJTSVFaL+/CcV
1bxwrZEuZHsiOh+MODSD5WlMq2zefqo1dxd0dkeV/8I8jZLAEAmcdfmJQ74a
b6vXqN3aXCWEx9Xkk8i+XTy81Lmbe3+j8fHgCiL4oJ9hglgfewqpXTV4zWZi
dqZLyHRIh83Of1n8LNjjBFX/3yf7SWXs4b6gduIr+EfTTiTRvRpwGFW3rEn6
yz7XUPLr/6kSmPa5W0fZ4IYeN3oVim9JJiUvxL1w5xbFE3dC86mP3+fetjVO
L9HH+iKcle9aCaTbVdF0htRqljxp3gZmjATDfL4tWCz8vV3qE6wIGqDPfOhv
HRSjhbMHlmEEB/mnsCu2Uq0mNkyPqzwdkDk6PyZfWfuKEJf1K/CqaLTAQ09m
nk3tMMa8Ls3a2QOTqdswmodFPwGPGlK064C4T3IxZ97zAd3TS+vSiJYwNf+B
uxxhfqbvpXQerNm7yx3gIALfXjBo3NXdjfbMpx031/K8w2PxjGcJnuWXhth5
q6bvx6fcB/zTZdeveSMJCKas569GEWYu03/jTbfn7A/K043z09LRmHOw6xiE
irOaJ+UXHKTD12f+DqvSJ68hWWQqGkpQc7aiFdUISab/JH4SMQDTlZc33rOg
vQbS/+iBSl27tJMSQbTVcKbs1T4T9hpSY+7TWo6Hb2BHzEu5os6WZhMFat7Z
1c/HvBMyvfZodtKu/rrJw6GNMgAD0KSERl3XQMcSFfw7uzEm82KSEp69cqz1
qrN2wZ49zU4cHwvudcV71KxydQjQigutMbu3pQgE97fTw/ffxTiBFCTA2rOg
3aJTiCQnsSVFBIiPFAPUZPRbX6DA4sQiF765jazzwg6EUjcogKQrm6/ybysx
bDrR4omnzNWivTvclOMs/Mgk9xkkgv9BLV4FuOY6m8+WRRBrrhFxDEXP39NZ
fhIiN98qX+X9i/3IxYGt2yR+RLsjTljdIId3KaphyLHWuW4LXjZuj6kaSYsM
NEzmNKPm01U/75VhA3zQ7TjXY+7GxpabS/E10dsMQ6fPOmF7FNshaPkBAWE/
UaVy0Gfxr1eVHvoa/zSwxCj8+id5W5W9Ejai5ElhLAEFHsggLSbZ4+z5kHU2
NSest3HDWaeVA7ZF9dydmkzqlmIFOMEMCMHtG5LIYNJ5L3vx47as1LAjaONS
lK0Ughca6bdgvXQ4VnzZS+VHN8bFAOnYyR00oGOTjs6Mp6LNiZcoDrTqns71
bsPaYta2k2S8vZrVZ10Q+g5ha7anZXReFze0jTAzk50ctNGiXwyk2GLCbLNg
0dhXmPWzcNvzWQNWEOBc0fpr+JPAlW1zp6fTh4WnWVyq7vpsfowZzaYehh1i
yXC/iaQT0RfBvlSwml+Y03Cjx3dGwG7ulxHysgZjngtiqz7KD3DtPl2tVtDG
bTuI2IqarQmsr/JLIyOX5mjyVdvXv2beW/OmgODGSKQaX/suj5LCUIIF/3LQ
gphhAeOlj2+xfQcZtF8r9GuQT7XqD/kjPuTQ3nuiPDA56QYNruVirkSHdcG7
LukeNsUcHgfyJOVC1TK5v5YT07Qohu5gdyMnNeaUDX4KPxqKJrwVJmnTwj5z
bznCqa/Zc9uP//1fl9xTpQk8BFUEa/mRNQ9Zic+bz65zphgv/0d5jDSZQ5K7
kDeXdVzGCnNdz+h958SIolaKPzLlk1+yGEbbZ2RCVGKosSkG/3xpqanSQmka
oIk9/gbi5R85KayM1u4I2NU2RgtapE93sRlTcT9JCnCPWIjXIXhHhu0bPiNs
mWXqWKWoPxwd17PXBOg4yqTgvkGnXZHWcXUoV+DoNgXc4wqmRNvKcouErnnF
bnluHFe9OiGxCIsHSrGa4r46apNmbUMXnnXEdBmm5gDKQp5ax/ZmX8PWfb8f
ugQTig8VRVT/VsOB7xiwUWtHzg0GvWVA1XgcCoR7K5fohGcjGOdXWGEccOF7
+E8My1E5/g+DmUU5Wu9mJQm1xL0BdzEZelX7yntIjIHOcGJoM2pXYOTHa3Nh
+3kHBux4Pg2UiM6/CyAg6WNN0k3ATaDRZDK620GrwC8YNDrXbDGWkxQWENG0
K1Yu3uWmXwFNL0NZG4uY3ciRubIGyx6HhFtrI1FeLqni3+vDuetaSLJtcewf
huzKGoQd2Kn+6Z10e/6v0Y23Je1A/QFWpP3X+2dC8l3UybII0S87rC6A5gcg
ZVTXZ/ghxHit3seWs39scs8vwhnh++JmnuTMsQQqzyWVlyM+ZXUtn9fjpkEs
WFb7K+a6+v14jY7Zdacv4HUsw8VAyKtrGcvE8J5T2gCoWjfxe9ew0wEHp8VK
F0JhDwzqW24WWplFCrxbgzx9kBU2ViteJmN3QJhLteptUO/W8VGJj9f3a+DP
zkKtxhEMyoUVo8XE5SayZ2yPXi3IpE4c9tSyNbhkoNb8UUA+YAOdVilVFLL/
QR0J9oCXoc0wTjBzdlXNHleOCngX5KbSvoLlwuGTDUViMt24ibo0DAGtqqCh
u/vOgNXFtPvulMxTKFwufizl8qft7a/6RlXTfnikS8CZuGrp4jaFeiyicdO+
h/lEBffy0et7+pTjY0HosgzwX7ucSwfO44L8G1EHpBjuFJOjqdT+oe53UOcg
yt2fEwwHS2krO+sqaHv6W5LvK2dOeOI/uE5nxlpvyYWBpgVnjfIkuWNDA9zk
joakcbzlkiK0RFK6TC3pTdsCHQiZQcLJxhavEFJJxfmRFoMKbzYGgulOanXF
b9NZ9Ug5I2JlA8va+IRKva/+7oW8h4WNYG62UFLvjkphxtqg3h2+9+khf8JQ
nys1XLvfagAZwaLXaYoHYxyQ1o+T2BJWQrnwclByroQJAz4o+TiJ+fbuJwtd
bIIHJ8Ze/Lht9QHK+WAns3rr29lAcwwvwvmjSPoxIAlOL0myKAcRA0AmxjgZ
zlaNv5JpOLO0e6SEEnM4y6KBtFxLlpuT7WqJdqBypaaWwnuNaSDAlsIzoLaG
iGObu8qEwRiu91akYegO7kbwwgquDkPv57wt5LXfvDmFqwxbKvJexQVB3+Ox
EPBNXm8BaJTfttQV5h/cEZ1jrlE1aWvlxzapt2mXjkJBc5JSzJMyKFOBT5VO
4chJL7xu9slXhMYQLWF2Iy+OPo1IOv5VLGlI4DMYkTke9B6r38DHZ2m6lia1
FnhiJGhiOzWs67KREERN007nqRa8d3WohypHawcRBw2MaxtrXV+eHDIDld0c
OJ9YuqvtTxQbkX88QTHipgHmaQRHLjB0WpGmLP9Rco85YTLHgl1U/vh0F9Yk
BjxNcVJjqNNJqCw+RoG1qGLSxh/neykiwclwQnRUKMDISUh333139mEv+/as
xaKTtlwmPh/H/S6lUZa0t4OzZvxAi9i9pX6EyTjPeZJoO2PQ4oDl0wl6PN/F
56ucP5suX3lR6U0hWESipDSdG91h045XXXoMjGrZRezkLKmuMVpSkgS1YC1K
o7foeg/IDpWPxlEI2UGflJtBHZnEXWNNt3PUuNlc+f3N0tEtO9I8ho172HHU
SknprtIn73r0YQA+rYOc3f/NVA/VOKEu+oM03UlclcWQAo5BP885gjO56KJB
NVAQcpLlgaQt3svlmj2LdhDcwCMVaWZ2JleJrr7PAbPPZNyZmHzXzsSAscIa
taqgMaDZ00Gg5oj18EvMvPnR0+UXjNWR0Nzfj33fRB5zPZy/nXNPPg4eENAz
4823Zoq+5abOgfFWN7PulZrXOFSxYcS+PQhDS2yzfM2DTitEJrM2NrA2cL3V
En8icnUMljv4y0yWQ2Q7Om/c8clOzxNZVUthKvlmDV9HJmLPAUmcgXVgTOmL
bS75u0pAvsItMPgHOao9rWjPSHUvar+A1LH9iUMCd/WeCd/BhqpvSrtjMBYD
ZQ27ZlQZqcgTie2b6NSugHuBUxUslpFVtHS8El08m8hmfOqcmqtcGr4zB0JG
kRx03U4pPRMbpby9UEIyVfBYlb9RGpuQUbW5ycvp/u8J1s2qpDsXlKKuhsKd
B0sqZIVwmuDiTNmV8A28v4g9ssfPjK+Bz4N+4aAgXABCAOCIpgarBPxhNwrW
mVSiF614qygifl7jYd+BDJmiZOua+X/ArvhSpi/L5DVQgayCtKoq+adt1IVQ
m0vtUzQFNL/GFbVxAI2eSOvcEpmxUWZZZ2F8Pedlr2GuHDrwBGzFIo8HLYhv
W8dERkqIwBEugHDCDFjIrBexCJDrhmrDQbYHoMvmnLeCfmFIladInEEJFFhy
FTneQ457IZkdhbLpvEwvAvV5GzupI9EYwL2VXI5LZq6+M/eQeX1kI4HigVyM
rp7ZD+GZat4H7RwsXEWPqK/BittpmPWah3clWGZtjFkp+zm4bz9FKuLr2XKE
0gfm6RxLvX+4bfYCwZsfjCB1Cq11OCQNzyY3/RSwyRL2FzkSuCGApa8xPvqc
gQi8nBNf8UOOcPqJffF7T7ggfriuOkCzN5UzbJPoYISCiEcV698Q88is8ycd
afBZgc1NSfdBskLec41g/6E7n3zDQFAw5CjbIXFsF33/4UQFKpYHsCOICW5E
Jpla9j0fMgvVvdpih1NqdY15JBtb7luMlWVODUhbiuQ2knWhxGK69T/G8CdN
YH7/eCYAZnX84V7zt/4tzRVvmkiiGC2LwmgtNr8RX6RsnxxASruIw3rGMnE6
mUG6PqNVi9ULwmcwOHOl169evMVKE+yyOqb1xj7nCUV/6/WBOcqqs45MjmRo
TqQOGqlZMAdUtYRh91wLESjf5yUFHjDE/SorJgEo5WP1Yn/qxbeRjJz6gx1Y
woHj9RIrtym6uvbU63D0ZiyrNSF7wDepeTiyc2lKaS7/hJ4h+2GwodcLyiLp
nXSfMZJUktdfk02uv+60g7uwSYejkUz7aM5+U/QZeXY1Nuqs1wppPOBsIzEz
hj+c0f6JUqud2q9ti9j0tWKZMATuIDe7lt8ITVKMWGpqWVTriqkvtJ/AXISx
m1CuI/seTKaW9+zWSn2Va01BUDVxpRSjUn6zCfR3uf5MW0fVACLSs88vXxf3
7FRk5jC+3q3ADNA6hnfNHZy9HaNDsw3Nj9AVnG/xTgF03tfrIqa/zy8ceWfv
01n9UUzwZndBfoT9M+3bfKjQcKMT0T+1BWd3Kj2i+1NbpWxoeq9ch9ryh+Ni
6Yh13NZAiz11Jewa6/JCQb3d4E8NFrD4npWWVDoFU6h0GJYIgrc98syb9zGc
cUFTSfnIUsy+Mv7ZR81F1cmjgdrp+Acw5pH7EEms/n0CvqE2bC2dvhffYwlv
o21r2EkWsLmgYDLzBZMrpGG1Nmw961vaOIgb8EOdSXyS3qS9q3r1UiY822+O
EtojjcNEpzBh/kiNTwbAXbJkInjMVjVClYDEdBSz8duBARhw+VKuq6KNEprO
FfsIQ3dipi1Pd7A6sSUzRrk8IFopH9ikiT+fOqQWlZITku6TpT2Ou/ijGt9E
+NUMgpuZft97NtTg1W44RkqTin/IihbeV5Bv6hSBJLyGTg/aPgnouUhTeXJZ
dwxBY1hxPrUQORARRa7VkNVN0u2Y9ufSrqXChujurHQPgtQzC0F0lQlOi83V
BaQYmPWsIgEAr2CHoN3ws2BDTrw59RRDBpOwLNfzlFrAK1ZSczoCpYYte44Q
2XLEj6oeAl86r1JDurZ3Dqfx4ZNsSnolf5khUveplvxOj0hHB5V/+SwABLZw
9HH6Lsqnq1FFeeUgE4nC4OGS+IcTwCzLP7+HEmy3KSuS514VQECKZicVEOph
PjFH9lgRsaEVs+71xH4RpEOvz199suTOS12REHQaZxZtFSbpur5OSY8TJ98p
DN3JsI/ZIvrCZUT5lE2Pn6RxkId24keUmcQr2N8rFZ59EzQjsXlDz/+qNFaL
wZW5xAml7LwSlPCa2ciaJ7J+4mheKSD03scwrl/ITrKAKVB8UBi9ZeXslURR
Ji7kvoyNn0hWcOoSATpj5jHVHCKwUuDy5cYUORazx9UX9Bz5MPwpc4aRggmZ
0uGXZ2Dy/5fnYIQ1yufBNf5KxQ15ZcO9hGGHK7O6cg9P9z6WSbB7SMPH7nQO
XBzceJf30yC5r9Lj+r/juI8QClZq7/tKe6aAIVkRckQXOVUbRzs84W8eK2uW
mECEX/Et9epqvNUSon1ajrOnRjB7gW0zmFpFglEPbx1XBAeyd6Qo51MJ1U0c
USye6srWmbYYhwVKRSE9j0KMJ9RkuVvW3/iJ9ROtLvBssm/ZwiqdIhHZfQ3G
vftcZ54OtPD+GpCh3OJSQaxoz3m4NGVtGCBkaxLo7APY7PNjLaH3unJQcV5p
1om9pMJz9vbBjPzVQfLqu5vGGx4FCXwxXdoed34pKdnDDaAOcIj/pmymD4Dy
idscgMBddxU35H3WYIb8O1OlCKRl3UUh/7H0+1pKFyvDJksaN8JajX0RQvtw
9diqQfBc19c/q/rkErJX0LNxUuY2ILcB58AxfqYWyLpL+Lr+jqii63eyf7JZ
I7/LEVdHzcu1m2eKuZn9jAJJnJhfJ7cCx1lEzWidkIMUyMTnNhEwiq1Z24ej
rfwmUMQD2w2puFWxHs4nOjoltBmY1yEdoeJocEGz8brLg0gZDOW7/uzjVdXi
cFNq5sxh8dqBybWraTTJ8w726iiJenlVzj/ukf4SVTvtk0L7EFdBDF11m2oi
OdUUG6N5LKr/FJqWqx7UJCzUhO1F38+abUQR8/lpA/HBEF69dc9OTG+Y0Gmn
+BJ1YWbBJqqr87iBhk+e0XbDJsmBhAH9Vc6v3jC9QbG7qaSNrgHoDWydjdEW
xxcZVof1hd2DzlAKWrvB1LMW4E/AJ7pvGcRH+FRHIycxA7ujPuB0gnaaw8op
hAXIMEqyZpN+bLTNc3ZDc27Mn36iSmCmHmshNBbgrdEeOT9FG3EybELs4XAP
cR+Nf8Fwp9MA6gda4kKL+bFy8s1c6D40ZAPBRntGw/KJhXwSkshuIhBw3gvC
tGW3IywN6oYjCI4I++Vjl8SBc82kjXNvYJe4siZRYSd4Jgi59pnI0T9mR+Cb
gK8MoTejqZOoD2VvgoRKhVriBnz7yzwqGy4EY6GiT57NvbHIBXO5HIhaSfSx
ZEIh5WmVmULrBOdCZy9t4AflAxpdXgAUrgmG/QnbJKwlDkFEQtjgp28UNN97
iyKbncnRqGn8lOnnlGwJG561qJeVG28jKLokWvG8x5AyNKLYWG2X+BVNyoLL
zwPSlnVabbFQ5SexQugIYnVTQPAzkkQ2teC7KyBRezRimuVvJ23VP6IZG/cY
1zVz3bTv575eoJI1G0rYB5ciE1Z5TzHkmY0T1bOo+G0J1yssYp1wAen2LM+U
9hNNVVAekcOnunbsfdRrfyFUCFPLaXIxeL1wBZQLFKiqLqJ4fgisRtCcl8Gk
lBe72gpP6A/TmBQzUtT0I7jiHJgN4fFqc8BNxYwJJ6xCcwcndJ+fDcz4FhMs
EDa01quho58gTxZhOSNxKgrBTJZCoIzRlmRr5wdFlai1nzdW+qndK+FzSGLi
LDMRS0vuUOIq/xkovB5eNYS5s030aCs6kuM8Al18H0GjvEU/ckHMnG0O194M
iwbzn4s0/K2v3ibF67LZW0ncuwgZVIQGeCQUZ1gwPBbL2Zjv8k0xOdW5QOBp
MSlSwgk+e0C//2M1cUucKFIAxSj/yNKcpzmWukDCgJQJIJTT8OcM+CrMNOyv
Fcq+pNEvaTP6kLvB0NeaK2C73DKypid9HY9U0oF67pGzsX+wGA1WC0uWlwVw
d1ucchKJ2GD23uWjQ611PMPPxRwu1s14jAK3VdYwPPrP9YGPgi6nxldvFMcs
MS1AT1GbU0hEQ0xgSGkGFfHC6+qq1CnWkbr08lGLVT0SbQIuXJRgwJ0i52uy
FyuBQ9rmxqeWJZbZaD1bcqgy3rOwyWu9yLRYWiVEOc7q+7fInMKsVQY5tPT/
bau/hn32VE7QGEGb5r2tpmBYxju+jDG07OwLTOxkf3a5+OfbmYWAcFWb/2BX
0jMMlz73Q2MIWd66I+ncOCE773OKyXh1h2AP7ixMVWdaxrfiSEGp05Ywu49s
zh4h/wurcKq+YKQq3sAT6HDYAl69MU7ajuQB6a7Ox7fpCua1E8u45fCrHdVd
36Ek40sqUAcbQdZVcAihH67H1x7xjcQxopvnEp3bNw9jSiYy0ybG6NdFQQA+
IfxAjZY+HYs1kqlJXEMrZNXLy+QJedrZ2906KgndS7rcwAVNk2Ch+sIf0SEn
BHsgJsezzkzsOyL8NuXKgs7tOH1K0+eTaH8n/wDcBNmHCE3UIFf35dTdSt/t
yDIRVJVM8LfNEr7l0xgMxB2Ddszcxn6OCvHUM453al0jyWkyoZvpikOc2Rli
/O5kxW8XtqHjhttuX6RKWvN0Z3+ojHFqlWO39/A/VapCacGu9PQrzzr4Tg+8
jJJ8loyBzfAekj9Yfja1KkILnATFOMDg0rNSsdgaswk16/+E4fQ4ouKV/Wsx
Xii8AOZlVHjNkHlk+E9m/VbYWJBGdd0PVilelD6kGKdI7Sx0yfpz3EYST6Km
icuVlKn4ZufCGHsk9Jlt+eArXId8wamB9aUv7RfIRBebhZslWjM7PfOjBZaD
qZm9GXK0ahf85ISv8osaCYan1sMKth76L8PwCHg9SpyCnDGJp5h7mBmIo4Gx
4PpWYYMacaYn+DY2jdTKw00TyIFJJZ4YmPYGC5F/0HhykqhGRSB7D9MDs9Bn
A1bCNIva7rx0UD/LAu3iPN3Vhec+JAQ8OS2vWVPA6iui5vHIkPZDfUEbaYN7
14QTh4pQmq62qx91tV3KiPDQqVyodpDRJu2LFFERTMmhzQguoRzVJUPRY3c/
QYkQ+YOdjjbGvwYJ44rt6Vj90X8i4U76F0GNNGjtBzSfOaKDGKe4+F+vB1VK
bdUfZfug4ACqqS84m1NXK31+XaEOaQcevEoXr+pkFe9POffgBesldKJUSg02
nXctECVJ6JRvESZvwBGHkAqeJ0RZuMLNYJvBncPN3dmCFvaTvVb7unFb6aZX
yX+ICqwiwDP9u4MuOKJcSSfQ8/w3zXWNicYqdAuzPyVcaUvlQ6x9MXXvzhBo
/HlnkWhYAjamimO3Tfvwkrr09gmujVBsxo2/9SYMVVDARaENOly5enxzI3K1
uVQtxsybP0R1r9xKdxyvl5wzPD7y0YUiGqCX6WE5fdik8rQVu29GE6j3F6Dv
Gqz1G4LWCqWU1pkiPxI980JCqBVS60SA0tqoqHadbep+bvP63NwHEIw3X9P/
MjRuPQbwFdsTRatLTdXOJh6H24AXKYnklhgIKQJPhKbFhu1v6zlX/qigEhvt
lB+l7+yi+rAivsK9+CSVTXi8CinqBrned3N0g4m1du/pHIzD7vQYWhrxUH4w
u1PfAeL5Rf/ppoljzj6bRGpJCMFNOfOdnX8GQQMGQ8BWeV20LThLY6m/rh4y
MTynxXmw6A4whhrM7PkRkxcjpPrGZvPgsej2EbdXsipRwqc0sB5W/BZt5Xsv
tLPwULxgK/BPLzaiYw37Vzj3Eh30MaXJbiRFpcsdU4y6Oc8yeN2a0x2ao6vl
kh5qXlhqgDiHbb/h0Ucf6KlRk79HQOBWGwRa7rJJPP7aKRYFCHhWey3vD9rI
GvIu03ZL6Kv/SKy8BLWIVZr0rm2gG+W8r2x4i+sEiT8fw2mJSNgGPdTj3PyQ
W83sT7UX7Mln3bq+jQGKb+ogFky66kKESPhdSBM74Sv6zLdU5hYZU4OxDLpu
FObRfw8dTmEt9pDsEkzUhAO65rgU9TPappSI4q40MmxhZVor4d4vEMCrUcsk
9TouXc1/hfNZlOt2YYMjmbA5rKYSLRYztdLk/Mahbb+UavWIB/+Sw5J9iLmj
SJOU44waz/egNpiqEhStGPV9s/T1qsEI9u8MgvcOO6rXfoEFdHK0qHsBjplh
zCTpotBNiH1PbHZA7ZLNoCT4R+ZfyFYyY34Dz31+T6+Dc2X0KLiamBSFtJox
P3kHx77IUMdfDAV3q7LWt4dfbT9IVLHbtYGvyBqAHDpH+QRixvvwWd5i8HFe
YwhuV1Q/8gAGSxFjRRprTT2ZAI26knRnGIHtqaxiqjtNoXyeEXt/iIvQjv+j
igtUxWDiRdSrB2dbI5H4PK0MR0cXnN0Ml2KuvS9PPFgBOxMWitGraeL9P0kW
mtck3DXJFQ7HSPQURc+meYeVkQqvrwJjpQZYVfzfdDq2LMQEg3fTDJ6YuwO/
0DqfMiIXr29W0qVNRmG962m85E/y8adLHuiLIRNRItedRG35BKN6KDRmORI3
jNDrowpuZIFangdKAz0q4Zn5//AZfzUY896od5052vpgzfn4/X0+HaSm5hnJ
FTX6B8zHht+jjNneugPv3mcJA/oLHycCBpUtds406lpdCCs2sdwLYCz5U4be
v9Lmh1B2H/0X+EfZuT9B+BAkwl8G7eOj8TwrwlD4w3GSLGPJ9kan6kzcaIdN
ihc2SZuBCnQxEfPrMGE16C9MP32XblB9LyMDJWbybGaSLeqwtN+y25Y3n87W
muPSIekppFLaaWKfNHn66bFdk4sF/UvcmzoesK2LtTT69+sk4PsStj7as1v6
c0kAhSDMerdbVy9WEbeWOqouM5v29V0cji7+L36QhjaYLmujKPhjYOWe35dv
GP/FcGCrNmG9I2T9W1TOixQYuTsOO2rKBwfZybpfZPVJTFAkxz7OkclT296w
yUQ4ZEtgnYMO+InEqIk0ViR/E2bc1SUqYISZ3aMU5VZlpohGF7nKZ3O21M8H
j2gQ9sft21Uo3Mw7TsVbCdq3Y43/5w/bdSrgSUb/jlQ3gBCjUH0GsR5wlxfC
jRr+XWnZzi2zGEenxQngMqlEvwREAjCJ5zbSuEu/DGHOncUthXeSsvd3sLj8
t8VzmLgTY+EmaOpf//4lhVkb6U7Eqh93Elf2MxnzxfG+Lpg/ahALCpFJ2wVY
e3CP/mmtxoxilSMB/I9WBntQxTMZ6D8ZqozdjLdtIcKi+9rwMNCEA9rExdjU
jd6lErPDzjEj3udDeumrfTx+zjHgFg4/Eg2sW7Y280vB6H/wtNTJB2l1z22J
1YtYGOpxSC5NA9cNBV7Q22/lz2NzFK0kf93VsDqASOBK3aMmlDsUa6E3QzWH
rniSNhQoRQkzWbCDzIvLkFBGHDOdvK+SUStHsPfp98i6t/yipiJ42WtBiWbJ
1XXiBN+gLxrLBFJSrxmSrziw599Nw3nS2om7fR8R3Y85WdpbNb+bBcGjKQls
3mTiZf1H1rh3OfeV/in1GQqFJ4BURbMAr2aE9L8L846Z8Ndi3MBPvZus/AGh
R/VMPd78r80lo7UVhiu0D3BJQXy7FrdWB7Txa2utqpaYmREna0BjfAuJ0GwX
gZrl+gY1OdpyFfv16kltO1dilaNc+Zi7+2P8lLuYutUZr0Nmzc3zt4m+zMlB
+74xJIA2WMbEy1dY3ioHfQQcazvttryYdwSqOWfPZLmgy4+ReK5w0HvOtfj3
QVzTElOwPF/Ws1/6XCBHZrcVCE0X8s3wTwhaE5WcVapvQcFu115SO3Txt65c
r3LDzZEpfioQ44O4Hcegd/M6bQd0tePKJtHyfIPOVAAB8X8yRy9aQ9nVgEZW
6KQJ4AljPu9knT/3fPhdwp7Sm4FcD9YQz8uMaIcdsfkOYwvIhxWb6Jmn+hPV
LzoIBJqRe4VCzKsyaFhUD1dPmMjCI7YqIVUq18vjDCifQJxACiZyPargV8EE
xOBfQazr6XozQRoghsQhGV0PaqZ1tZHr5sWX9gE1grpldeDuzNAoSJV5dJ6O
HfKA3SYBS4HJCvjE0JpbLx9Tf+Pdjx9EZCRy3qtKwK1xG47S7srKWEl8DOqn
gjW3Jux3BH61kwI/cBXJJKg59MKIdB1phWbhBrV3f85PpVk9kcn8P1laxh82
0tk80qFSKc7SGP0VWmn2sj7eufRIkJP4ndX5LNDuXtsHLS9k/hSZ1fM+j3yn
8/FiybEQZWm3BtlpKWdHojxCivTG6tHApGrZRR9ZudF0HMVfkDiY8y4nCytg
OQhFIErbap1lWUNwCLOKfEItDHcnUBfA2Dh6JBZCb1g1zs3U7B9eDV9AOi+v
RbNxQr6NzjYoFe6ZKH12BWXITRcKsX5gj440YjYAY1V8UsSlxV0Ix9ohPfr3
TjMWL0LX/iLBCmUzKAUvRNqxsAMqRbPhliaFYVuhZzMbombNX9U9ECio81WG
fmf317BqAjWyVGRTgIaN9bIazxXLjD8H6FNTjemPSK0WftrTggF3JIjZjnik
5n9dBGdfXYkHBWMbXD2Qr2cd7dUPiJF5zrz0GB90Dg6Xqj10KN8VZTpOzEho
bTDT1k3ffQ6uiIGSKgSBK6DEtRo9zrs6eAQ5CqnLBZ6teJSY952qCNzzn+B/
UAz6Vukdvt8+vy5I2VlctjIJPBD0Fcuq49b2nj/Dn2GG/2gPuLd9jvinMxLu
LhPkIv2/arKNVmW5QcxQ5W8+wOizvns+hp9yEg7x9zr6a5s08Qbzx2kd/eTh
K5Hu4v0W67s5YieZsmYaJ1jyWmrvLTLgcWhWRalmN2IdI7jY5Tj445wQ+Lf5
DdrwN3bFvylJTlm5TljqDkYQeVwANJyvJg9BPpfDo21ES8b3Dhu6WmvEerop
MUf25Okmt0IO2vfE+jXhNtNEtodcTwiKczKSgMXdxrp6BxGpTHvS1ZVVcEXx
HcqiArpNou4ykYhRZtk2GSknvN9vbXLPMpebRXJ92mUx4QY0srIiHQ5EtJdx
Y1VKs7uQClEfhMCVNqbn3EpkiCOLD4GioRV8E2e28aXaj4ndxc3/ym4oQr5n
yi55ffQNWFGNQD77ah9F1LEHzoraTNxYiZ1DcScxZJzJlVwdOV9YZOWj97cK
4uACI1HO5+Dn7WdcH8TecE1S9gh1h6U2htlL9UrJmymy0p6rQhv/Hwthu1yp
Dsw4MKHU1/qrw5wnP8dmCkRSaWJdGOINafER2tckXBLcvmibYj6jdpcfzo+R
RFgHBCuyhdKE6ic/GGaal40nSnnANmqL6DlXYwerlYjFrhlf/9RdkBYdBxlX
eUK1Xs8MbsjcLfaDiFQuunkDMYZENM4LWnAdofBCiF1WpPm/Hl6S+dTkKQ6b
HxKthiZBVRXfAhNles8MF/tQfqMTlGn93KwZoz/b9KLxYvXTUOVgH8kunTrS
C2GKomHKuZQ5jTaNX6z8vnRoe5YtKLrU6NKGX0jrq6vAt1jnHNXllAwYgzX3
zuijJyxAka3PIAu8eJac55OwcvRk4q5d6rdpHKGj/lrUv5cn1dyANhomUoAw
Al28QEzTcgZ6IJV4GV0L+zEHuyyLTj+oaUSefpYM77yBoGUdkvhaOAptOnwe
peZgTz51K3ctfpv3D0wXt+X+tiJphKl0QqZU/AnZ+1a8EXtX2xU/56T1Om6g
nUMK/1xc4RDfPvvPC0BbqMXeEBulyXWbvpVE9zfqb3HKAAMx5KLQYa4KLFRe
LP0HLWKVYYntx0j4V2IRisHN+sXn+0JybgVfIiLh8Y6qEJBhZJA0tRLKWBkG
ecMUPWe6XqGwlwfriCLZxI1qYK2WuPeZzeFq3GNLUQRXP3RxES373K1Tz3zw
o2w3P23D6NwFmx934+u6PyZA99weecCzmXbbgVnHStWX/3qgl/o9i0gjIgfe
bpN6uFnjyMElD0N4wGf2M+kn5bbcbMZb09T1fVzWl6un3lf2cyzjVmxGRQ0w
NhVOK/4JRPiZ6JsxeiXN81LZmKGA736Kvhehwu7YLFSy9ww8NGsfXCQVcaPq
fH4TiSEypdI2eAMZ5hNW2bAypoIVkLl7lWVJ+p6hmMXWGtUc0RD83is3gCw3
tERACkCsqypV7V2R9UJBywmUPg9aKjMZjo7WYZ4ut7hi8r7pXTUz7m5Q1+ta
wm9Uyzrv9YVM2CJRHmDL9r4Nj1Ts/tdPwS7FXCvk53ZIOoC1WZJjAdVCYf25
/U0B+AilO9y4yQBIGDaZW+bbtwaowFT/zYnVlK+bz5MAjU9eyZz6WIH2I0Rk
/Jw5xB6GiwvvD3VL0VRtK5KZCjd6CK/bxGB9DyZQGPeIQir9xpNk5vNetIKA
jMUfaAS/oFixzQAcvQSTyGgeG01iEPTIoBBNwybjpiAP8dE5yj0rf6foY/LQ
WCRWC9KMgQEkLS3BEtmCJjxp/zbxNN7VCYDy7nkxgJY/epp5zq2xQZ06/oxR
/dEB+Qg8BIeupKS+X0944IcACTzgvPS4ZXhDyBzOdho6V30FS6Ngnt3ZutyI
PujHDEhiUbfuY8vXeC8TRCUCbjbSJvCsM62v68VLlecjY0QhGHQIR4s7xHKo
ol7y+x5kPR49u9HdAb+XZCWwwFow151/THWdsVYqQYxBjFKNgBI6HL8cgqra
KpqL0ZlyvFxW1N8fPEi025SjLUvs0P0+Bw/HGa3BSOaWse2DgVai+tTWAj6Z
K/ylThNzb7EK+ZLgjDJhySmnXJ1I53TPMKj5eM47am14nz9PFwmEzxKd1kDe
fKo+Bevc+ThnDHJBeOi8pMe4di9/v/iGkcC95iLorVk6cUVNQ8V8uKvkbgDc
gmnARqpFOtX67E9dSLl/y+8se3PUpZs/WjQaQHgzH5cRYB1E0OU5tI6DrGJB
rt8RU7A1tgf3SgfWelweu6IOjWMvn/RI3yyNcYLQRGVG54fT0XcNF0u988KB
t+WnCEpuTNQcPrnnu6mx90cNXie0Sbz3v6sWE9wHp9YWtzh300KinPIR729h
fLRFdA5WE7i7AyHNy6xHKif6CdyFcmY0uOoW4frvYy3KxeiaSEfp81hbDFkR
nVKX1nEVXyT/ObeJ3mBCE4CKpVmHSxskzjaLz9ZWDvMVbO9CLHvKb5RcLi9C
ffdTQlUBu9jbOm1VbU7IVyk16RjsMIK8uYvnVi/6Sy/5DbqQ6NZNvtKRifQK
ILTUYxU7CK7mZpge5ZoiVgRp69pL8wmFuGQjoSHq1pJaWWDPsTuHEn6sOWWb
UoZ3oj2R/QbXMrIJWrgUgE5UIyvCZg/mtpMabEikBYnHFa7muT+YBz/eVbJW
G9o3qe052tFQcOEvqKRMF42/3Hxfo3n8U0gdDT1XpXdcg+BGcIp8jqge20MD
KfKkO6/rldUnaLxI7iDfjj4o8qOF9zMBkBzF1PFzzlN/TPDs0pWIfaDGFiyH
SFXpFpBsaQ7OYGrs78ekcdbnBdgg9A84KE5eqJTx8yMH40dwYUTdeZmN+t1Y
avBtCEijifZSteETUEs3pWvkZN5i1F1IgijkQr2PmmpHylT8Re0QPgUMEtT+
yE19V8Kga9Stk3xDhJwCLoWjJU8crDQDu6pZekhLd4ajb5/ZxkA9K8FZ2yhI
OxCLXCyb8p6smnwLnr3hhY8A2kOx8UBWAfKiTv58meNh0btbJlFFtCms79LI
e8hkC2DwQdt2KUwURcKDO+Khn6tf/BkgIAsJZraDJbU/wh8n96YAZIXID1nk
bbb8RvAEPNg0KJ6sqtHfivtAPU1IeScnolgRx8eWXMpLMhOKvCpJ6JqXTvJk
GIJDPvxEKj6fOzKBejStk5FisktErj1iHfyGZVTv+cgQ4ly80gAj4cimoDYY
ZBpB3qhFetySBryrJPIq8XnfFWcFl6KB5t1Qx0uPGSsOmfjClxM7ttuTaNTZ
uJmNDhf0x3rL4ql3Y0Tmj2FJalGou0ORWc6HtQE35R4XqfyQJMDVdXeXgEA8
BDYw7Hcy6guOmPgCrOVqMVh1vx+onHuhcDgCVO68kuf7MbHser+xSmSp72Oi
JZM8ZQ62WYv8a5OEEaoqEBOrTI0+Xa5hN5+gS4n+Dl4kfwMKNWkbrbBXs6U9
sxzYKXmyp4MvN+xbefqfRk4Evh1IQEkvgPoERv1j8JQzoXDGeoyPOX9st1GH
/Iicx8V2xKKCzosS0RYhdVNwedoLWLDgWMXEEjD4SqHt91VrwEdLw2iF79Rz
JEQuP5E5wRrbkT8Hf6FRWnRm2H3RolggxoMqYqFqjOmmWAjVTPxcR4qzI4ZZ
lhDM+cw/mkUqralUmQtbCijRMUYSdh/L0Qf8HsEq+pmbJ+e0WfE4VaD74Dru
6kKwBY+WrmR6Pdr/3/UQae1rSa4STxkm7Dvrvt3jk4r315ezsZrjMtWrigbY
R7qau8cjwrds8CauX0GLDpeNI6IwsG+DureMBkFTos9ZFDrg7LC5N3LDO1QB
vW5zjyZZinfLExNp6T2IOn/bNc1loHMfmaaVNynAROFyEFwyV9pQ2bObBQjI
fBOFaXDZodj0M787aBWB6SC/tk9DfqnvQv+tSM/fIYMgEsurJ27YCIspdsVl
1je+uc/8DiB68+iYYwRZQ+TaLA3mxsHYdgwfGB9cgmGB8Xcs9EcluPOkH70H
C2tDAJe1ct7tGAQ5GrwBPTs+AvbjYC0W9XT+BO9OlyNfkDLQXPr+O7L40OYe
Y+md+dWpLIzMYoh6Cah91GGbTsdDybeOt5XVlE1VCY2lP3qdF3Ljzio2VKGT
/xuKEGW0chtzxoC0AAezYWxRU7cADHBK4JqHifgga3NUK5amHB0fd92C13Uq
4VVJnYxIVF5kjJnYVrHffaiMdsqPSzU4oI6zj4RGoCnoapQBQl2Ep0+8yPn0
DVUD9imA6+3MdN/634fqntEhj6paQWK/z6TNOIbzPVYIXXOmDhgLY7TxOdGG
A7JnUPy3JLDwctxQZXKwu19z4thwytM2sgSWYiCeZkLG8pD10CvuqxnerIL4
AMKM+TvvBApS0CInkkvsmfbZBxPeYBtBluheLQwyopj7R1WD+A0GKuEjrC5T
4+wtfKA/A3uxVd27QCjONkAcSIC+rGT9cosEADoo3f7D8yH885y86yG4LEMs
YA8x23l11vrMvhVO1oGdNjfv3MAGqtQMLb0Is8ZL0aLRNrobfb7ot/5SCkHt
pdBay/9cGLelRI/n7Nj4C3b6fbi5B5VwbaJIxqRx1k3HqqSexb/hSVrH8R6V
blB4LBjY8d2Ll0DuUVLorYOSN7R6kJFb4U3O4J6zJlzQCcnNV9Az7nTOSmv7
k789k1lUymzWHVeXQiH14h42LexDjuWI7IUpaxt+9bAiKCbcSsadDVR33qJ2
IQtIddVIxkhJj8abR/DJNzEXUKf8cspslDd6xpL2jmNrOdwSEBOpdScN6WoP
2CrkzVz7RDEeoIq6S+WG9eYSqH/yXa4Aaai8zcMHtR3wqnV1t6oQ2z74CUKG
tiYQLJRYUSYHSMi2Mt7Bkg5EDLiMbXfIf+Fel6dLUS1TcIKV7r16uoyxR7H5
h/nB5jiPQcAK13aOEV+oraInuMg4HG34IIT+2ZHUkEYB+LQ7aGvtdZHaUROO
PATu0p26BZx5zLM6dZfS3LdPoqB+d4+W34oX8QiFffTsYfiOL2IwTRZCkhTU
TKvTL/LYreylqfmXcpOqWLPW9B83dBZ8w7IuojMwxYaZyg/T7B/DHjCEkWYH
0kNB0dJYoZs8A+kXuvMAK9roaZUiM89+i09RE9FqpQeD0roSBKRrQMTFEv+f
N5qL7qkAoFt6+F1Sq0UsS5q0h8uWgU5SfUlDw4tMo0JB8mCVbNeNz6kwcWuk
x+BrLKRMqAhQj26EnpuYn3bqjNlv9+2MJTXJ6cu2sabmZ2leLUP3VTttze6B
8qi0VXHv37fbFYfGBXspsD+LcvW2knHQnz/FEX4T7RIHZuLnTW1Ju6aLq1FP
1MJi79aXecLrzyYT9K96dLsNwvwODfjq1rq5pLp8gdaOWfPE5MS+o/aDVDsk
IjfH8GUTIOTs7gq2cOF2h6AJHHO382bos+9p19UAAMMon10U88wrRzEi124W
4Cu0sMkP4eRIJBuazQC/I24kvHbepV9y8X4/gcd0c0tX/DWoRukbbuB1m1gK
Zpm1id/+vauHptyRimIrsbHU6O8cncuALU4csOzaLMFBMsFSVe/Lmy4EFlin
iA/aYumedvk81GGr7To066IrsJj3W2E3N2z9ZN527BQNbhn0L4XnEctDm4OZ
ZzDcObp0nQB+VhCjGVNaNFxtEBof++5+SAWReWFMl1I76+TDVod3P6GmPeQN
g9sRQGtzknY5ojnoxy+BaHNOO4SNdzI4kfwROZ/bsUwNG5srQ+cOlthWlmg1
liGH4LUkl/0Gyxlo3DOq4LynI5gVYwYZ2kSDd3dQ8OHLbfFgYubiwP1KslzC
63XZZp3wIF+rSEg22IhDJNU0atZvfMvhAZ+J1Nq1tpIpvVj0hBsYF4rmcWdG
FxGUgT/ivxp3CvoANWHvM4RvsEHPqeHTTNqWPSfBFUBUrxt0DSo+WF/13ByM
WxQ3v0ogpjqM4E7pmKwAS7e886EYEPIyJxIcahCCjnuSaT2zQnVdZjjJJHCP
y6C+xU+F+AnoH3arEidClbFR+8reKajWoM3g1QRURLMSmwgs6asN6hRpszhg
Mr/gFx9jQJ3YP2LNHX2mWYRfCV1aJ5Qh9OYk9LU2pod/hFSAA6TLvBRCZeTN
Uw4hVBn17BQZYE5Y5rxqz8nuCsU07YoMxiOeONuG3REuuKlwb/8m0GyExm/M
qQRDQcpbtrRBQTdSTEMVN7anEPvcadjB4unmAS9lzo4CdDsz2q/cl+fr5n3A
ANZ/fpsda6vPgd+s6t1X4M9o+Z5japEEI8DnlU4Cj5Dmua5JnOz+Kbk4uc4/
aLSXxvd01gq/S/oqe88RV1OXPcE0Dp4MX0pIjpSOwty2myy0YINOfMQVha85
uEnvlsq5Wob8NDM4fh4ZltuyNXiH+YVMhBiEIgg+msgNcrGt9wyXvCelBzte
l5HGUI2etk4H4P3ZVDuFIARUS4pmhGcEH6NN2BNutOVx7Thvsia5iFptDdsT
MbGjKtilv60XbXsUDCgSP8l66FSj06p3Chzyo+uIc7UTbb8MY2nosGxCsezI
dSgRlBmYQ6vqNUfPDReuPRC77QSKG42l/20mArkpdvwyBP1xQeiB5OTdkhLl
RX10YO4dYWN3iGDE9mYAxQ5rouoD1XM+Bt6aO+4Ewn6N+DyArO7qwXJCqQNY
jsCZaNzzh+OvAt2L/VfdFa7DkmouX86bXDj9q8M47gAS9utWTC2LWchdr4WF
frXf9WtOYbj4ZVdcCVSXmZvDGVAFqbrjTF3ZdGvKpEJ3xWK/MGlx65OKFWaD
N9+xkII+5U68sfqDJ+tD//9gxnzgB/NcCJBlgOmNmU+mDXpd/8idCCHoht9h
/FujWVvyPDGH/w7Nei3at6CGVikZlpGfXDDiEHm8OwE34s+UrPmtWDct4iIM
XfDuGnd3Q8h8uxiGCK/y8W3QivSw2H8S0yy7aJOHjwneaB3PehWZ00+Q1aOW
0RzJpsE7TPpo4+xgXAtAWAn0DjbrRLUZGJl923qjGX412vrNoXH5wXc1pglw
W3caCVsNlLKx1bfIrV4lw3iPDwd6EqFNVi660g+mJyCjn7MeSJdjKAVTlT02
1rX2Tj0ko7QUoNwxQd2JpocrfEhbxrCK2jz72jji0AslY2GNGzXUyE3VQULh
whA+2xJcznMQQun6qQGvppEslRSS1he7WB0gqscXxFWV6D+lcSsekyhvHBeC
PECuXWGcHjk6EAsJdQlQzhJQOcbieM92uuZurEp81JWMxBjfCcGyLktIBgFG
uA7Dj5ev95+k79Ms7NSA8ypsFqmwCv2G0H6iH3cbHDyK0+lNRmz03T6RtWCX
tCzEWLR32n4sUc8jH8IZwrPgwO4axgUFnFzddwTBRagnp6HJoJRsOERj7iLk
sN4ZLq+E+5az7pjdTR/GSMpVJjh5Fof9eQ1JkbX++OQGLZYdTEJXFz/K0cOq
aNmSyAYiKmsDc+jssw9GzBOlDnQcehbl7ERZbdKMjkJG6uOcvROv0TwKC19L
YJb0c4eHw+RbX32Tp22zUfXpg4pw65Urjp2zt6XibyRgCj34wFsHuBpNUnkw
YuFPWoZSBUIKQ5ymN3NsYgbFo310G4S2bHML+/pKti85avms7oAvlDDYMPyU
cVUbSngU8vfhQ2Yo8tZTPypHp+yHFRMMSYnbPm905h3MH+AL/W2EbFmKnkXg
GJfuG47lexwMckv4yc2m4CmTRP0C29a+V/g2E2sq1I9Jd/U0CkpSHbxv39aH
D3nJzGaljzATi9CHbu3Z5WIFE8+a/NvDuOeCyCMp96VkRPm+/wDv2KQN51GE
HkVu+rNE+y7zjXUl6yN2CxbcpCCBVWwM55dRN/c6ISnu81c0FGzosEk6PC0u
ei0BS53AIV1UKumYdswbpQahLJd01U3T3ejnzm+6rQnWGmt/EL5IlU3Nx/wF
BKXSFIXxu6leco5qCJ9nYhcJyqUZWekfti16ryUNqIiaxxKSaC8SvDS37NEQ
xjwQKzlkXTuud/yXQXpxiVPcd0pI9etg4wbqAnBdN1q4tBMw+CoMtfWcZ1r7
BFm59pLyDY3HGvnWcGzM+S5P49Q2Tal9XXRUDq5uK8n7PRaVLKa09v3/1T8n
9o9lBo6CKzDgN9/zZP8YFlH89XoXLcj3X0mJHrUBHioFkyKQ4F0hrN3tF+TH
FHPqu4Pj8/BAJYZWu4PTfSB0/wh+JxC6s6SJd/xcTG932FZAwDNoXhVy0r79
pSOo9d6FDSVrhpK0GZsZkr3LMmJH+zRIgzLUtoizKsrKaDRyte0S01miEq5e
4iT7H5TgUnRkoeYa9GGAQ1S/aTUUS4oeOPqiX4bRvJ+U1KUoPlcSC+GfGr7w
zUyXaKj7MWF4bKEHJwoKa2bJkk54WLwqKgtmBLsS+5J37hJ0PQAFhouw5/a1
ffZCYDAHg65xwc3uKfaiKYOWOs6Ma4d1GpZ07sSZOPscCFKPEfIqcmJ0zQ09
xqYFTZRj115bbIq60huMNUI+qFEommum66PRxmzitjoSsz6gaH0l0W2VMf0m
lHTvnl9AoHEBnd49nC9GGUG//IiXNU98CQBCTOX3MdEPv1ErPu0wN2kqHW8J
2RMc1SZllMRG6zYPFhgGtulxizztk1YXH5yJwc8QA2dZokciUOrvLelskhOP
c11Ug++9O3jT+zuK5as5EBJFYWob2EXLtd8f3G3mwOR2SGCM7doN08E7ABrn
h+vrTk8eiRAfJWkjYSja7JqYxm7KeEZbQKdW98VUSTC0eDQBH5nWRhZXo6nf
Z0NBSGrJZ0neGQncjmg/pkZriKAXDPftjVw1QD8u8NyQb0YXRNpeRQ0kruMH
GCBeQ0Z+cj47j6ug2UYoWEaEPCsXM4T4z49lyYuRu0/6lVhhCgCoDVDIKN2b
dkiZAF/UF2qEE74vwbaulvGjILX022QkOlh+1b8Q+9rqJj3FiUH6ihnd5yCk
TIEUxmLvqF6Pz+5t5xXknwx8Di8kZXss+UeHl4twPqGMOgBmEtrXqGm0IdVg
bWa2OaKasG1+fUpHBaZNi1sM3saeLYKO2WkUyNR4IQTRjx3IaSrysnF+bE2G
hmk/5DLIGQ6Q7ZCMndeaqs0BADVbj5Dyyn4uKheLwJTKmAAvG5CowJ+TkDYS
QO0OoCT9+fKy1yJ5wF1fepsP07LsnvhVWMYKkbyfOI2uv3asDPjaHahgMeDt
OfEYixtUzhYpTepar7unzXcIXZG+DjZSJp7icAl4KPqV9hgM8pKpyetlOpy4
gyiFX83YaW9KfEq8/4aIcHR9iQYhn4iDYtsUZmVKxwk6XrZlhx1QXuvF2c02
4j6ca8bRoQGgHdIyfVgsmuGm0wo9qRMpmI064m8tvg7yAF2wiGy4vVjeE5+g
mRJeOTDhTBbmsi97xVxOrUqLuXDRI2ZURRGkj5HDnOMa+P3MR3Z/e845zq8A
+xXRc2KB40KEB9EckUvHW9JykUxzZXCK5M3To8G0HVvPTiQawk9OGxL1Tgqc
9BIfEREa7+7rbdIrVPgs6RdZEIW+zcNqfLy+Zare6wa3TXFSBTCYSl/w1ONB
9dRycYMsWrPbTED3kqDmwlSFa6f4K8wEsCVPDqFDUW5p5HLexcCOqUinN2e/
CUq2KWyAcBaLuI6jJEx1+A5YoYB3lCB1k/1JootqDzWDXTmXFRmNAB594neR
H4WJ+/8NorGMyyzbpP7P7tMiKx1AzgYQVfJVsmJFo6r8F4NrsEKATlwdPTTt
gPJ1UQPyetfaidbfSNwmjFb4PzNrHCe/gXHORxyKFIvss+D+jmUWebn9xwER
uaVvaZXwHWVtHUaBlhX9ZbV8CyPuYSkcKvcitZ3tovi6JXjI77Ncib9/rP0W
jd+XEBpboH+xTodNS4ybYMMgJpdFPWZXUq5Cw2Ok2CD29So57rALY0ycGXA7
jTObYtDeNeAQltnyz7qcVM7YPbRKkcqsjhqDpYpRq3n6df2hB5E/Vvxo41lI
eyI7/tZpugq68qUR72NKsXsGXNsxMrzG5qrHreACPbsty32SxlVFUf3q6sG2
HcNCGAyxyT1h1W1f80F0D6FftCIcg3bSRiOqrtyx+eVnCf5Yu4tPec+wSWlV
Oo07Nlo7cMWXZtPhN0L7M8HL4kb1ClPcQnNkIQP8MlsSfJd1PJyhVA8rvBAA
F+ITwFc2pJfEd7IBDIImz+VHY8xFM/TKX6jbDvq451meZ/WZfO7/REsIKIKx
1hBdGiSTmz3A9xpK6mG6zyDU0FWTid4ZojOnuQBSY34DV80ohYG2ASZMyRr9
gMUwD6Ivqoxjm/E7uV4hOnRKiuH+F5F4gePxWPLECUVmQjQtUST49JqxBhxQ
giUNxvtbASN9x8/Ji6Ahx1+4YqpAl3Xdvv3Mo2yBmYtcsF/2/B1tBOv8sOLl
UnnDCv03RwlBqTJ3R3zO76/cz2t1xJgw2hR5iMlP/eCPZ0af4xMz8qpPogcx
L2j0Qt1UCPIDSKSLG6V8Vt0d55I7EvTbjy8s+41euvtjsoQ/z82+qBO9FcOq
Fx8572crJ6XQheJCOcM6Jrhvh8NF+a2Knrbb/5b537LHKS2nTklE6koLLxDJ
Btc2wWlaGmGs46PmL5L0rddt8+8d19RqKiap9bfjhQ+GZreDl4wWrtzOSR5O
FabCdSMUbZMwslt3+YTQ2uKz1ARgGKZ6jekUZsRUQzbAJ7uQ1drNPluzdGn6
3BC/Der8AVlKKNzL5TxDvVaV0W5GT/UuZf8nbYABwiRv8GqyDovIbNCGOiJ3
rrWhSwR15Pk3RHaUSxCuvGu5L1CZqtIRRMC9DZRLP96XjFsQaAowr1lmQq1F
GmL5G6TwnZHRqjpPUUqZGaw8qwPzuGrVRU31o726pJxug5yv3BM3d/4gTZpA
ygGvygbEXRtx74Fhj1R8STzpkZLQRFX58q38vAcGkRjMKctx9UvRC1bdXu1B
X7CMV7ZItd/vFLFLqgrcUVp1v5VVP7InifBojFH2WFwZGJNSFpxUSWRtC+0o
ofnT7RroOZr9aTZmHJ35D/4ysixDdZtGs19TJlsKUsiz0+Rlxq+Qr9QkjTtM
FAoCdZFbj9hMdCdxwXgFUEP0+CvCoTANotX5R1C7h27sA5BdLMdi6dp2/6sG
cB8JzESAa5hmy7QaJ1qFtrBL7NVq6chtjhFCJaAsKL6k8HXux11xW80e30TM
yD0hU7JJr3ughmBUamH0FDDQHumZEuuj5e225rM4Cmb+/quvqvDlLzu4qjhN
rQe3+wLr9j05D8ZgG+WIWS8Y2adCiZqQB9NAHDsz1R2Af0rZmzhEO1i6gZju
G8nahzFT8HIH316aZLWW5DZ0Hy5M+6tXUGtx+5nmYLhqZL+V6Lv06P5QJ5F2
C6trTN1mTXysykgWODLBDQealnnd4FoLaneaqUHPaCeW9WYXl7M34gLEmLuh
kKSTN9CztRJkcz4dSVGZN2Acdn3uwqY4MIWubeKpGIxHO95fMgVW8+vcWBRU
qoZMqwmPowPnJw98fBnSmkUpQ4mw5kII9FJieMF7mDbUKCblvtr7NRTqGxP9
6OggNu/VHm+ZsDw2uQoL/bMqXN2/ugtigRJfBCdKCDYSDPasjy/eFdvuOI0W
2i8U3G3dHegP3AUeDnrAPtpLfVXltsBTvSPUi2lsDserPZMs371K724/5d7P
k2qF0o59d1YQj05KAm1SCarmAcuB6dcLIpXP9Vw2gl4TDGtzzYB3Dx4NayTF
SisK7o2y5Y/DNDEU/0gZq0clbp2Ta0M8lo6hjKX4AL26mb8cmXldjX+D6E6m
/B8yC/UK9kb4PzTDpG1U0Ewq/0WW6pSHAnpioUJRhcin5TdQ0OglCYL5LQVN
Kx5xH9Lvfng5KKja2KGosBoterae/PkRIrV1ZTZ6d6izfXdFc2ovyG5M8egr
7WNqkeBXWkN32SWMevW9GKUFr7KeAaYChS1k38NUzVsfFVPuof5AfpcArHyI
5P92ggPuLbdi5BJ22AJohQKZpuhKwGKMkplTORKoT5U1L9JFRf/f+8fb/kw4
95VIK0bVPv3jMvqy4KKEBWoUGXXb+1zDkBxyJwS7X70cQfbwCpAGsUn515L+
BwEQ2H2BY2tZvUUmmGEQVGRcp1wbiNsLTm3SCgfaum/oH4Jp5SvXGaW7m7St
JbwsbtdluTvSAmC6Ib5BK1Jp5Fi7AGthqEjKCZ1Imj8CaZLs1t2xL2HW8wLD
BixiJWJEmB7M7llCngBmWDtdYA2iWIAJyY8CD0QKuRLhxeXWSgNV4i8aEOLF
Bwb/hDhlrUov3hKLlSw/MkQlOhiBb8XD+o6Gota4/V92dl9FxFVBCw7rdd9h
bUzPNEo6ravGh88xABTKOL47Jfm5TmEBCtoiiDlHJwCsH/aNC5OlQ++o6NGJ
fIVJS4Gr2oyqhHIMuQM59yag/v4PziiYyz3gPNuCYlpuYs0K8Dq+K9LEM6Om
iJwQr+R3BQbScAN20RpAQ8I/j7XRCh7LdekRmoQ3uqGROfcISQ5HA6IqtkHA
1vCw1mASBvlpO1n3nWs36CpHI7/fbmkIj0qP6E0flCHElNwojhxYATME7fxO
OrhvemDcGChKY6JNInEvt7gc24MZuSX4vhjeI1j2JB4p3+SSwFYrAhabu5la
AHmY/hd53pi/qldtoZsB3ND2AiVrj3oHMo59bLXR1go7m3KuuDaQGV6w1pQw
Zcsr6J6TQbykYNgpZ/dl97gV8XN4PqPh8c08X1Ac4eKjJmoYiIEVEYXRcj5a
KoScoRRikL7Mvib6WFTloPAzrE1K2OPmbDjaVjIW11yoxug8h5KvLqIfezpe
yBKkCUvmaagZSGTUCCyTfix1p2WrWyq6yJF1Om8LCVmaSKdtkGtVOxds1qZF
uhRlIpckgwjlwKjYefqcjgoNJuJPDO4JkV0VSgN0j1rIOEH++MIm5Lv1x26w
vl/vKkOxuHaeAzJ8o3NQfYrBWWDHGGjbUf3XkwBW/kT2//gIhcS4AxIsYOxv
xOO3IGsrAsGb1cmyeoT6YGEgW85ctJgTu59xiIf0jMHc96UHE+l4TfKnB8FS
WWo63Kt3fSEsBNFx8l6sLaCHQ/9U9E1jE0tPcQxrzuqXR7leYD9Znvgs62WR
a62kXtv76lOHKnInCGWgX8QPSOEjrsbYo6MrfRvv59jpQdfitzDWkv8tPsxE
wvZ4CSQD4YU2tbfs0C6pHZ8HHJkEduWC6bEa6UOURdFiXGwRDYZAlBC0030U
zarWqrrA9nFy8k/zSI2msXI4p7Ms8GBu5MJEhf51isSgE/p2hZjPryIyzYSm
OvLgrtHpeaDl9W5WCm4R/nWHY4Rzr9uviV6yyVMMxKrZP1JnELcUjwjubQn4
45+Gm4GL9ZYWdQqkHSf0Tfq2Lx6f1M+Eo+Q3iuVIG0TSUGx4EvfgU3noKD//
aEOlfLlo8PzjUiNbmR8oXpPa6c9+/R5BTy/e2eEbJaOpxe4MONfHFnJgOngd
Sfn27WCdAZ/ckJl7ADDAOy1TKnXLKgKyNUjYl9M5/oz2KHi+38W9f+v6OnYl
S/i2b3vdLEzhlfOjySUszXevSNIWY/aR70mkBizDPayH9JUshmAdYCJmNul9
70rErhszGge+nzwncguSW0qCL//XWrsDebsI4mASTaQTiExMaf0IDHLqzpvl
XPcURUPjt05SZM3o9wOuKqLIcl6Uur6Jo07PFRcR09JqJzVzTSEpYAp1Ok8D
e4nC7RHpeT/SUt326OO0iFT4NXagrxNDpyLQykr5yqN6L2vPU60IX+F5MafG
wsGh/b6jlfrTdT8xJ2QkizHaWSaaCyAUKXAYSbi7ux7btErr1imQtY6ggvXp
668IUdvIskMvxSNf4jBPN9vjIGz/tMpWGz7jfwt1BFaANYs3Tk10WpI0xnfC
7HfNx9+3a5dYgeFxo56FiziayJv+ILps5iBbs3Hx/OlTkkBcOOzbvlbooKma
UOSOnMdpQv/bJhorXqjDNHVE4BgHyAJv0mtCvyeNPX9DID+mXT2q3ejHELrC
ZIQw2z/LFszFsdCVAqrxTIS3OLamrJcomEeRv0Vm4pRqwLcaGnbn5rGX0PkO
pzzHatxl6RVnW3Pmy250zA7CkvRyDE0TT7HymTdl7beTH7z009NSJLFXvXmA
cOp+9VoqgJkhmwkuac552F4hyU0bFSM00Pn9SR+xBx82PnybZAEd5soTyU4V
/BHjIl1kt+x4RY8SMLUeh3TR1bE9Tm4DUe/ggccJBSiMHXchOw14D6V/9HV5
Axf1tezjXbP5ax3GfNSXI6yGEm3qpxvrWYT8YuG6SiR+el3/SVCo6oX9SFF3
DKiSjjeAqjBq8xvBkao4gJoK+f2y2brMzQBbNTJ7fjJq4Z7Ar5SfVue1iEoF
6/8LDyi+LhtJQeIwRxzyU485aec+4HZ3ZnreTPrB4jLnNwThpcEIS5oWvR7K
2pmzdFFZ5kJW6LPoYL44K27fXf89/Spe30FRafbHQz4rvD6FMYjznumt1hgH
cFZGiylRpbm1jeqBbou4j1P4d6u+C8i5UoNLRPe12VaPOGvR+l2qQBuk03XH
3NrfoOckUQRJ9mJq3BTa+drb9IGQ1YhqzZkdyz1x5kinr7japHF0M0kkb1ZU
OIqpFmV7N5yRjWbnS4Udst0URW1IbQ4oMzKYQvkKkvidGUbU5Ne8eX2VcqFp
cDFRHSHAnyYOc5XPWTBRcUpOJy1iwF2UENAiwVD5gLAmrZeZC6UXlusDklX1
DlzI7bmiVjAikQW4BYN6yNRVP/r5nsg2NQJjhD+qlGtSIKuhHmn4YuFOGr1A
mxVNsugk6Gb8IrCJWRTjjaDzNVoxqzovrPxylKPf17486rMQ5cRnB87ZNZ27
DliCrsTyQEBQxrwDbKCJkeKQd6ZZIkwQJez4Slo+8ffIkC/NyHWyXs9mMu0c
IPPj1j6XD0gwuozTI7r+VcqgPbQJGdzlBDtUdcgdqTipsCm+bBDv+BQ+KFT4
MjmWXwOFUQb8+DN73eY86Y3gc1OLLxNaVl54dhdQA4lhpy3xcdLCeJtbTtdL
bvl4WuZ0hlOooMZhNrkwJ5kCv+0A7rJ0fIpE+vRIlsgtL9guhXonenfQLtGw
WLvG12W/QRwhzdZChpZClsgkUlyntN21XSh0XvRB4GFMTMAp5atb8Xv3h5c0
gOgfSx4k9PbJ+warikvnCTotziTcR15PQ7yyYgwjrtDgD0ANP1O8637+rTyz
5JNXE5AK0gBLciAmtMWAr+Hr1vaXSnqMrFBU7gvuvE/xyK/Hvpm8M1aKo1Oo
y4p8v+7rtbbvx+PBYlqTh6Rwu3TRsiLrIGWD+py2rZlcqR2y6Z0GpC7yiVB5
gWIbfaZUt6xKgPHOO1IDoDY+0iSfVksqoChVmCe7Lf6fmpG2WLVDSF0uuBs1
HA17W8rXUwIhr8a75K43I9fkXCIkuGxKaHyN8vtPqvpmMbhLxHuBAxeu2P34
Dw+TQOvRLqVyoLG2nHmsCCflYXrQUMIs+QgzHw3nxr9hdc6GYPDaosNhB3Se
290fzbp40CLj6Xt1MIN7NgNsnX/4wdJ6sYt/D2fPwtWJIOi9UcvhwBQLrHP+
i97eEKrWGIyeUHhtKqsXsWtYHG3XKRdJU2hWqqd/RzcYB3oKWoGOOBqZpQ4k
IqIg7a/SussQSGlWhDAhbKxJ7t7fxo1Pz+SYHrLTqIpWcWRt/xRMWgK/qPJt
hePTyb6Ijjquhalij1KyDpo3qHSoAF3V55LR9pADbrY8Au9JumiCiW1KoK4B
iV/EOwsKbcHbZI3rSHpbF7Pyyw0wNtKyv6eogWfb1xfh2oBW+SMqd47DjwqD
Q+JBP9qNvOrHUZ7gQb9EGb9i+WeCX5aPDDCSypCJyojyWE5Uf9Sga+KrTVxf
+FRTjOy4MQh1RZO1Be2jJVAoUBVAe09Pgb2nGIdUSIOK8h3YajPiCz92X+Qb
gZhEb/2FpkIOgrdM3HlE/qiScETemynAGwAmUXeHlnVlvNXtNKACjf7goCNG
CQs0Iy8IcNwmAEuvwyq3nYY8ohdxemGPRrG/LNOnjH0VXERIjMSq2BxPUxhX
S5a91jWONfE7tRUPEAYkocuv56W7Q6RdZUf1PAIzPmkkD5oy5Ax+4XzT34mO
bK7S4ga4Fieip/ousa1xjVHT0StpXrMOrIvAn37i0p4D73K1X6NwlYCypJDx
8u2DbCvfV61HeISa2zuWruiXSzCjBAuN+10JtPue47YW5YYKfQiStcRy8xrZ
CpCgDI+UKfZsr3iit6ejkX6Wa+IB9kwO1dXOqDo4/YWoJ+054oeB+L7zEOkY
ksWDA03Equ0ho4BYHzifEjYxE7YcpWnqo02Sxlx+Sm+yAifsnjiHWYNk15Q6
5GS82SnVpp0Gp6qFQaqJa81sDJvRRZLOm7pVYaONz2MM1F+yzkNIM70n51qs
SHXPPVEtvG8iDfafyn+wh8Gf/B5a0uJ/O8ggiHdlSocsBNWV4tGisS2Sv895
1gJO4aYa/D2Ug8qqkHBhWeOP5N9pOVahu2Bk1f1nzD+oBTVrErUiF1njI7pa
+TcPXiDqE2+lgZM+9pq2LlSJ8f9hK5oZh8kx93TLczq6nGzy24XoEfOACsZW
Ej/rcfle0mF/zhTrIGv1rINpXPpNM6NE/zEcCGu9VjWcobxH66H6Z00d8Vln
Sdll5x5iFYLyNOmWutgK1FaAOtU8ZC+IBf1aYOlSZNF8BJsETBYA5lF9puWn
vOjEDUe/TfmC8MdR9P7qtSdjmrxFE3hlJeLnk6nKp3FCcQh4UJcVyD7B2s4c
/jceeaLOyDfSonn9AtiM8qAG0rUymtF7kaIjIR1EHtvfGmzEDBzD8rcRHLB2
/IaIUwiITo4xG/23+6cr+4numizxDNrLuuZz6nch7Kvd+Y1Us1OzMkx+kxox
Hzt5GR9gh3OxWFaqXBfzj5IjatBB/q5VkNIdBpqIqba3wJQoJqq6Ssm/5kil
EN8jw1nF4UO5W2I/YwxDukHE3OwcwFiryrXglyT1IucN9cqtkJ1Z43Du22+C
eL5w+UbVRvsafnLQTfgE9GMGF0ND1SxO1flbBowmShkjWyu8a/V9tLdeG/AW
Wqs2Kwt7/q5IefA4JICiIF+Cnrdtxrttk0dojm7WHOllRxnFfUEVqfmDpu/1
IIxVAaxp6uJN5OejFU6PMabRTdI9+SOsDR9aOczOIedGSx3KgEBH7WS6Ny5f
+o+7Y2JckDbXeRGgnlu03ZvMimGxehPjGNr0od3GcZ24nspyeDoY3ov6+O4o
6297F75t1NiJfVV4bBVlbGSCDU2SmtnlXek5pWmauGw+k0qb10wbtlwCi+6A
8r7uDKGDxiww6M/XlNMtmXOQhd2kui/aO28nZWaAV0a4PKoQN10solPSTsbm
k40kjJfSZ5jKbwAT8EsQWLXVVEN04uxFZF7TkEyFJuuE60JVuhVeVl6fo1lb
8bxoWUVc1xQGHII7Zqad8uWb3UQRGR5FpqZJF5ygXqqqKxjDeUcUrpi+IVx9
q0xTdxjyqAXMGxiwN2XzilDfp+U7RLCjxNSjxoMZz1LKaBr85ZStamNAfKYN
FZ++siQVrIpf8l8VfN6h3P6rVlEhqIjipFHcoMJSn7z5gsbS9wlD8VQzTMEN
fcZMieLdDyA6Tk2BFeiELJe4nTPC76L83iiroE0NLAZQOGzW4N2lyqUbPWAI
lm4IanKQ4T+LHNTe07LLDPSxlo0kA31t/fVoGfwDTIDKXh8AHlY/IU+9tcBm
vdR7MW/P32SVwHBqvv7vk0SxJRbBe+vSFLAGkmX7OLmNoWbGx2TuDMG1kh0M
QLvdBaj2SYTHzH6r9wX+Sai8Wx1/rJ0tHd2kuojktXGEtvTVLvdgL4RqLbS2
ZQ6WabNAR5VlzEG3l3gioZ2L3i00IsFnlagWuOlMUF3uWMUKuj9cETTWilO3
CyXonb89ppSbCko88HOKW/GZ1QsvDbIq1aMasoxFinMQ/9Q1UxaahuGItcr0
U9CJuwBpoa6C25DhafyhKinXefXndqji83fSVGAs0R7UGrfwMLNNhA8KT1uT
uQghFCT6AQGCpWNsD5BtWdLokQdVZ8mah5Xd4CcgZdWXgVoEJJb/kt1HfR95
CdoR6NNJufxuHqhFLgWYU71RIDkfUWzw3sonicsehLrdQPoz7TYMLwLxgSAQ
+ksZpNj9bU3Lx2s7NLh3R2qydAPqV4WlpZvA826aPohepn4ODnYafXZM53oX
oAJFY+VN7SGUxCEugF54edvlbly8ZsIxHqtZciPmpI+gAkNprRMOJGYM2AYU
OTQUx1b6U7ZiThgGoADTn6HtMwlpiEb+WrdmKDbKHwtXHdgMVP03M33LmqvH
8NBdUzzq0YypfzGITdch7oLCJzj+lGn34nV4vU7taRJ1SGoQPCDFWjGX4faV
05cyPPKEL6vvLxDtwLjV+KpJ3Yq+CRSM6FHJ3ZqiMNWJKgcAzu3FIfN2kNl/
hy8XsIGhQ4CCTkPw+dAzrcddfKgbM6NSYwpo7oOOe36ZobEcFvG1dMuNgw70
hC7JeL+pWG59UME3g9nyflaJvIqFMFEjmK4cCDlps2pxykMzxnbg7WyEl3oq
22JiFzcs+RIN2+WU6aK6tiI6F1iBOqRpyZT4+pDpHPGu9syefarbLX8/k/MH
pgfwuJaJuQU0bxVAXyhWooj55Mtdh5OysCqMg+K6YM2ou/ZiCGClR9+dgI2R
/xVXSycOXpGdTAH2POWHpTr0TUvdLIcaGOan1kvy680wgE/2GzQsZ3a8WHsU
ftzu927Q6FooSNlEQ7x5rEOG1C67MJ7IJtuEmlL7Rg2MB2tuKJhy1QabCT66
oypdoVA7M1UhDlL/5NBTP0oWYmKvqIlDKmTziphqssKDCjipsv+DSJwn246t
v9ywMACt5Vi4jkQ/dLGYyDL5pLeXLGxOMaOhFIxx8no5au4AvqXgCojJ0OQT
cj0019Nv40toRygL+IV58UAMPmGFX3rWYPkfivkGEjSmGPLl0YSQW2DbuK1U
dl+nj2LBg5NLfMOF8EWQn1xHzQnOD3WAnVLEKWBHIpqOFKEiAqB5c8JYuBs7
B+GNzE/54IS1fQRkEdc5pDJJz6qDoCnzlAhRDrQucQMTv6TDIa8GP3E6VLmh
IZqCjD6mfKM/HGgM5jB321V0MjFZ8C9mY+QPa+4ZgZHwOIriOve4BmvzmGly
bUK6I0PAzkiF5yOxJhwP3I7VXQ7VY13RZdG/HDruoPLxkV8pvMZH6pL+wYLT
IuIhI54cDb833TD7jrPwW7qMbrm1Y++1gilrsyYECxU9cPgLCbOs6qMwMwa9
dV/njQYpc2c3OEDuJGBadCY1n/eAVL+P18DOfo1ioMmgH8YKnyRC/EzPwNOx
En5dr7eGv6hzGLChcgYIdJedZw3PVo0dQIk04F7I5K0E5u3oOE0Ai41go/h/
7KLRwC78wh6L8R26Rljg2fkpl+NDEhKRz/E08tlfO3Zz+t1SDoA3YfXqZ+GX
OruunTJ4rwPQmiSAin28C6U9whW4P5kVf26g/EzmG6kgSSnG1CTkIW2LZxfb
rW5rkNMrh6yi2+1J1HlEBe33JJm2fRd4xQProuZBfei9ybd5wSyxoATQOhK1
pzDdJqptyHd1Lf9k8YxuzEM2vMNBgetZLh5tbAlfBaB5jvjdm66KZWZtqQBk
Ok5JMhOPFqxzSfBUyj12tdypb5UIMLHaXVAFjFA3aQHu41c0i7BMuqhu0Pxh
S886A8MI18AucYGFGrklZLqzlQpGuu2MFTWTflKKALDwpP5/WH543Dk09eg2
lJIl9awHieMaqo4VCCvFI7uGveGXtTGDJsddqAEH8wPJL3Q1msPrrnIHpg7y
aBDtqfKrEg9kTUsA7s09yLBD99BLGKBeTTpNMFw8QyBLt4tAngz8dNItAjyH
lalXfdZYUgM73JVTijd0kh9poA6E/In0RjWV44mYlkyE9tbUFe72rGEPmpjp
K01OCqb0mw5P+X68qsv8QwJSkcSDG0QIMOaV15oVjB2iDPUwc+5c9sNi8LXz
wLqMpSbruez3rQ9mXt4vD6bIIvM43703DAupunukdxqJ3sUBp+S5Y05RwfAb
bldpJxolu5zka0imhKqLCFFlWuFCcsd9WsY+uP+wpViBrr032XmxVYcarvvP
RQ5anyl3ZX6MllSb2XAoAi3ib7SbAhviFSIMAI5nGqNFWLRImOieaT9bwXz+
RwkjFgZ+u1XpCDSToycVf+FI7FbHzSfkGUIWzuIrKDtU6EDzcDSDAS3DY7Av
AJ2WDMURYQG23nOj3BM92e1Z91w2fKstSrzP2wFTcHkb3aPNFCIZIAF0gMnZ
iJAm2Lco6OgAbMPgLEk8b4913+fqb9JUzct8l/GxuFG8OjcabD0WSssp6RKo
IHsfTChJn/LsC29iPHGQEA/PjAPZUAQ1VhM+EM8YF3V8BShqX27NhW8nFF/H
lIcADLtiAmkSubih83yIz71RtNWYL8gWPD4fGx+dUS9RFG2KHB27W3jITH6+
p5wlL7EVtUN6TLMvDIFWTIR4bzRH3gPdok/ILvCJofs9fk7s3J35PF5Qpgvn
2XuzIiEyYepGunxuhyLYIN77mnmAH26rxn8aTlD+QMwrx30a87hdci72YkKS
C5ncj0kwXOxNX3LfCl4VcTI2Cfvp1oVhlgF6BqLnXPtBhK7cFeJMquTnAj5M
zdzzFoBHmHqdaMLMNhfeNvKOYJcY6TftPqTXtZFa3NZ8qXUxs4RzHY/NrGAr
qqCiN+EJDlX6ejGj8/Fb+/v5UEa6DxAI6W05FyNxdnJ/rzCFSOPzcb/li/w6
l230u/aF8ueUZynLo2B+IUGUTEZHJBFCDbIrFFFp4DewtzI5n2nCF/lFcdyX
NuNCfQEh7GmBJwUOftk0T7dZnCXI2X8QdfDhV2Re/4i9S8xyl42MUzsDJY57
QHb5Qsoh9VznTgOhU/hYIDdc4prhWxD/xPJGcEUpfXz05P4cDZaLCmjSkvjP
9bXxsctA+u0S0qnubsYv92ZT428P61AkvFGVkvuz9w4Opb/BygPBjSnLLC/Q
9ocdAMiqoqk+qpXX5k4zt5MNlEpLObgW2ueAkPWDi0VUTCuRFnICsWoUnGnN
rGRtHrkkJTa90Nr5GYeQRiLZMabmXDQh018827DtCQu/m/6W7jk2/pWoI68h
8JTH3RsHNHcEVMXlv78ulGy0wL3B6A3ooazS4GWPc/0i1NSZf0CCyiXPfkjT
xbaONnwnrJxawOIKTRn1xiRLdfEbHKHwwilllMhR3xOXk7FFGO6VsL2uIiuH
pdTtCngpgLf/RsYFIoVcRSxaOS4+98ReWFJnx8LgLKsdYkBfMqzUjBd4SsV6
zAM0l07rAMSbv7XU32BGKa8xgKNsLug7OpRLJ+sIlEQtTXn/WA//EJrc6b3W
/Ze5J+7nK8uVOfj/dCrTwQFDAH76YIqOxW8WWqjXy6Af+DuWfTuEqyhPLI+l
Fk/jZC/gct5H2wOhIyAQDILFgtKenH+tGUH9UCuR3cefSaOb5vQqjtUXQa7x
NWyRd8LRYZIEFsFmQjO89vXX62seqhRl/rxc1eNWlpBnghn8WTOYJ1q19Edl
oxUgqy1xX1xkVFeLY5wBhz4TvbuV5Q89mI7PbInVyLETurmdf0roA6aITUO0
+7vyncb9zTsE0t5P280dRw7x+gB3gsQJfugYtw2KKToDSA4ny+beeykb1bvs
izm+Q56RMhe9Pha4FYR50/VJNaOA8C0WyMdQTAFd9G17rxkWT+IGjKx64Krf
IcQDvc4SWzg44h2hj3unSFumyHZ8st1uZO/l2MxcrtvCJ3gpgWdqvjra1vcu
eH5OUkq5+efAIz4FviGbiUnhI3YK0t7lI+Qq/BIr8rI/Xd+Es6/J2uWOO3Do
kOtLuFytFP0Kn5YlCMMNzOL3e+W3NVcKC7HD0hLPINYmrjONEYiiOE8e9IZ1
KafE9KiMz/MjRQqGBSUHNKw2afjECkE05IWnIFh/C1OlFWL9tfVOZQMl9RkN
syjmY5DoZKsmk+KFXlLeoh/qVxUZOrOLxfa8e1kP1EcDCYymCeJIRvJulUzJ
dZtTH1m7WG9ej8ZP2RYji5H64h5F32Tbfl0qwFjR4fCIqKpcn8I5ufS8RXzl
d9kZgBr4PWuK5KuFDoPesG9CW1r8V2KObxX1DatFBCpk7OKF/atH6myvMXvf
EEkPmnuFPfFAiJ6zI7LGAEYlMjwk1Rm13VC5V7Vv54tbQ3tAjuV/+1E+FWga
bAE6/qT5UAacp2rg4aRI2h0uLTsjpdvRdxk623BKIXQtqvmFPMJgvHp2NDZW
cQh+V+dU1tcV1Xf1eOoE9x6CadeuFYZkiq/puAI5BlpYblVrM5b+bzf09ZhY
7lPDV+6zVJfAaFGXmfMUSYPt6+lW/LjZFWsRHUd7zZbckzl7its0dxPAWP38
lHoLg3iZ9r+7f8oSUmh0cDMfi2mHa+nS6vZZWraHxkwu/hIRU/N/IO/M1QyH
1ivK8OBeAZxQcRVgHLKNDPOUZadEbEeiywJhwcX9RZaeph9SAFPL/TfT2VgX
aV9v+53tF8TXMtIJL/+ljiMXU4b3iWrBypxyCkzYLK57hExvc4kwO2pk0INf
vbI4Q6lZLpkVJXZXw0+kme3VuSZn6OqffUe6ZOy2M63Vo2UOZvl2ofoR0wtR
RALzxJIiKiuFlo4U0gugx9dqGNf5QPsuqXCX0xuVVOVhj04gjY6yfjy0+4xP
DprHL0OWFBUij6qzxaaMHuEPU5sOcprBsWgI+pYblocv5YX4BlYCoyJ50w8H
9ImNvuZhztPWYbXkBYL/kVd8BkihWG8BpfyJ4NY4pD4sMxy/mmFp+jV6OjBQ
UT8a/ZbEim3YINp8EawAVgGfSh1Bn2D3LYuXu9p64z0NBOkKZJlh94cu0gN0
LPfOqZ6WIVrCW7wOK0kFQwHiGvRNNlHv4+dghDqLJFq7dBrE64HYXrjmcU+Q
Ukuh0bY9eKjulZYVimopcOQDHPu0rAvhdFOd41DD53U8rwZwc2OcEdL07XRy
2JPollBqE4gm4SQBI5ylxQGfHyiyfOEWRvRKIWzJ0iSZE5dHUvzTBhTN/GYB
TOxuEGyS0hjyLYVRWUpzp5hXB53JgWhJP6qz1hAR0CefUKOK8kTTS24ALWIw
NUwOibtmxJ1aBP9YqQfvxXd950q6OUE9liAhIDzjoc0DGtzI6nVmjhI5uEC8
EETqSytkX7RRfCmOThrwCRVZa1htGMtwhrSQJmCzjOUp0mxTZJYDJpdiaPbZ
lESyetXK6xUjp/MK77/AjXyHvtH0G+qnVNRdVqAOzWjY19FTvBqQDvXcjDjq
oglpRRWA8UJ4KCGAA6LEy8t8TFUR9iHPHoBGO6IrLIPdfPz+z8IVozG7/6G0
ZGQ4kV0CdABRCRocPyJ5PYvPVUhplqOISVn1S47CFMre7/90n8fCZ8BFt0xI
9OYAxQZ2GhOKyuN1gpSq+XK2IzwIlHoorPWYI5djpbOd274yBhQJclE+3BF/
PulX1o7zj84fwn06UknmuFIB1W055ZvywlJ7kEIq7QAu/4u/yiuH110+ppQZ
tUG62bqK+l17sgB2VkdpNojipzvOappLUe0mxntiNZIXtXapEpPINNjpIIGI
9Rp2HdfHAVta/Upp5Yn2tppHnpaBOwQ8Mu2gQ6COFf+qqlMQkh5faIS2qgsv
ztBYgtzmyhelsQKcLVAOEUQPamiM1SH0tblq6MoCnsJWjOcKtBrCW0e5M5Xs
isTfzNtHeoFzh0YTjpaaVAG30CWjN8Az1r8dxMzM7bEFU88kbT/zt42uRt0f
7MMb1osf9GBBgnuc0+nLZ7Bdw4q3PuFxT5vbDKd1zpZu8zWR8++kN7cNCtM1
E8GQzF1D9B2ugMfQ5fMqdbSGsRPRERDOgm9hJwJP7EcoBjjtlrD9vRhkCFSb
OnDO2iT5c/MBPx/CUmT7TGBilk8BPkf5q4JYzAdcu62IOzpdzD8Rde5q6xIj
VKSdOXmuQvFjkxv/p6VMVaeZrwD6A4lCEKH4A3we5WCbs7+41GPSNsVrPHII
iqGFp3G8efFGElSRzsKpj3NY6bBDTBTPO2gZ5lxuZnRGzNhETp5fKsaaaiHV
pmSqYFv4+RB4deebCA0Xw/tp9myfOkPZ37n+ZIg8/nesA4nT+hq6ya3mHesB
OWT47auO9RLEnGKJz8K3XPOO7urCUhgsOjjwFb+Qb6WIRa+KxVgDiofug1a6
1KZl3QgDG9cdfNlRZGb632xaVIytj0vy0e2FXQw1XotwJIx5ozkHwdZA2lyT
PFzAaUco2C/ABuHP73x8oiwp6YitEl0BuILWM6D5PQ5uXlgQQrU2rQ48hu16
LbzYwV0p/jCWTbV2etkD/FLPEWUiOTVPszHg+iL8TzQuDVgtYyjZrOwH19ay
dlOA+F9V0hjNzzv3W8QzXcwLeiOQ5MusDXhfGTyehrSi5aJDdAuZX6mT5gsm
SbaMc94gtfgwl5c6x7mVu5XulLeLFtumKd7kDXx8THE44Gmvm2VezH1hgo5y
/GW/oy3B56gScSsEj51VAH2hV8svqPyRMR9h3eS9CtseyRE4toZm+lKDgi1D
Za5OAkWtTrJoUi/UGql8LY8SmW7ZWwUbpHqcNccmJlBwOrP6mdierMeL10Rc
LvS4kJhIQKrDRyYf7Sc571ZqtWft35O76Yw1f64iy9s4Cp3MVeZMumLNTK7w
IU87Rl3FWJb9FHG/Bna4gesNy18P51nJRSx+5Nm2QmeL8MGPsP9D0pDcmNQn
mEEYeEcLHfwJpsd7Z6k2xaboZ5sJF9JvyT5A0Y5jphQAUatEt4Dvf7u0uEcB
dsGyShd1JHpW9p/G/IR1J714O8IMzKxgQ87vZJmHB1XINwa4JOz8MtSGxDn7
nIWKKwEOUEjYj5RzVm4G7RN28BOfWeqM46K5GOvZLnsrLDxD0OjcSHNi82mX
cpM6MfVmHAvJQMJrb7Dh52VSmqIlQmjIaY9faks4vTP5BW7QrNnVqeD+MoG2
v6VqRmB9W/y7kiVm7m77oHK1JXxAcq/MM+oISVA2I6ebc09RgJIsowjNoup0
teq1fC9o8NLEHxA2usygGndBMe8rKAhlmsv8fT2u1MxxrdVjm1QxNurcQrH4
+vnlINS/1R91mtIT93XAbwmA4GjNHLzVyAQid6vNQyQ/dBp1ELsBvbycWqnU
nQK8UkmlGKYl7e0u76LIZD7dmR4z9ssPLdrhLtYlb1/13x2qKKGUW7Lcaa2/
WmWQNxjEmyI9xp7Gmd4euzKzv8qziyPZYZiAW9ZpKPw4SGsd8Kn4lMqexmkY
pondZ+mCHPrZ4vaiqqafi9O9e3dscX+UFSXJ2GEFykxZS4ULwdJclNgnP3IV
lMcKEHGrxo76kEWx0uifFTuUc+O5XR4SvWhCbQ+A0Wgn2ITYwS5kb5vspm/h
b6RpadAldbB2f1YfD6wYdUS8Dw0Fg41nzCHkXQCSFpzbbh+ihCyPGomb3oUQ
iDOJOVNuNMJgCh/A6fHGmqkwO3peK65kdmAELpSP/BUSgHO1HiPioFdupBur
KZnn4wJX8ulP6zut0Axbm8mONIrTt45vZF+i5eHyScxrUaqnVirhU+LliQsT
csMfSYE/8OR6nHJWg/i3P945HlRroWybkAZ+Ha6VGJPE73LNBu+9nZ7IViI4
muDshUUMYaJZqVE18qG8JZu5O60jdOaAl54DmMa4onFmxoH78O0J4qvtsxjr
aocnsPS8013iVl6x7bUXt9ctzX8ri+TGdk8tywysX1yRo4xnf098PtHCxJBC
3dY79blaMC7hHeDb7rlgwXVHhuJNB5l7SJT5BZBUumypu7JKBCHkInzoZ6Re
oFxSpyXtkqr/Gi9/B334QdSJBcJn4ucTPOHoVuEMOqn98FPIt7INUtnEhzxN
GMc2ThXu7oTrnv9xMzhD3/fT7cXVkWma3S5um1bH0pHfhrk0ieBjF35QbOCc
2A6SXk+bGGXZzwwuFU5pLptiUNJYfGPEO3nt5UVX67p+O9R7ALasJdEMgWrJ
UM0bH9ZXIiu/K5peTwkjFULFVwLLKs2EbjFaG0HNi6fo1hDWF8ytcecf5oL1
PzDlpGCFl8mRDm3V5eegOLMbdmvfBJv5521Fsabkjv82k2+Bu8SC1cjCIvgC
8o9+SzgZxyvC2jAGUgTSASPPjFSX3kj4+n5AKUlkgc7ApNOA2+uICPCjAazQ
u8x6fN1tE3bNUskGuDIcRp168SpjUmTxkVzDJ8Krw8AoId5IryKPBos8Tqk4
MYWpEFJ6glaunfW0X49CobR/BCrvu9IVRSBXuy8egj5PMvVy35B/3wL9pLt1
AIWIXPf7ClEW3nzITNnGfcoo5778ZUMrThXucH45jnA9szcLD9V7Tp5TpL8H
ZrvNJa6gZ4xyiQXMb9SVydazrlNmlr3WXHJ21LcDx+L4zcs+cKkLKnbvLGXa
16rxVJU8uIzw3UUbn+JOL6oaylX1MWZUwt7qNtsHYd88mIiRsKg+ndGOUplg
cUNCOLXjA+hfictoqYauaFoYFS8YC2RyMYNszEPYTVm8kJraP3cgMsvIShO7
6/Z0oewPvG3zA79KqCb1P/NMpc8XZh4LctJA0GaxHiiXoK73XpRZlu8jAVlr
oxBQUAE7XLTxFkXXmHpCInHens9N1WLR7+J22+63f4+crrmQKOjmJGg8KI+3
41Ze8pHnYOYMgaaqwpFIxfrNMcWpccUthIt9FQmMx67C3UZ32t7/qcqMS97B
/s/i3AsPPfhLHq2qgT9SCKT+6Roh8OcXb1Q1n6Ra8xMNmwVziCFiZD3sGP49
E8oC3Aaj3yHHQXZRTipahuxXvKFB7fO8KnMOxiu9SOrc1OwMqTZngz2Ecacw
xf37cfXM+oxqbJ8nO7NYIGPzIUwW8KYtOVjfgTvW+PXWgS8kXksS8Qh74KN6
QRZh1DG6MJhN86z38UVWRo8xNzkf91LNDtZH3tro2Gcaze2C2mhGDH4/ralA
c51RV9vm9pjgPeCxNJHT7cCnK66h9JzXkAupiaDyQK6fYBuCdcuOJWC0fuwp
LiERmvA9hjc4S13FqynggSHtotq0C7yXgGoeNGJRzSZqj+b/5YUeyK9IQGVf
ZMSB/7+AM2W1SU+T16NbWZClzMH8NYzEiBZB/8ad4I/6ojEgtkWR4qPvg9CK
7GsoYc5N8UnLIzzsi8DCr3NlRQug+7XdazewBqdpTQrJHaP/L45hkl4qWjBR
Qiv/UsPT527COQ+Qux6G2lTizxzi4dJC4nevW9tfXVxfqAi//JBnHkmlub7s
O0Y3DHpn5jl245HaEYt0UgArdtC2kl9rAlC+brKnf1QxSDqtvGY9hkknkuct
FpXu5FXxu7rJpc/Eg39J/fNBan3xSWRSwmAvB8xZK96UX5F2kfcAwjh5GpdQ
kKpKHaZ9/39fl81zpM7Fv1nWZZ2x08o0pOr+QRaLYSfBr6b510AlH0hdHww+
XztK2aYFYPf7tY8AX3LpdaxeppIgrByLCWYbzMJH4DouhViMPvdZ/Zfoc7/U
Qj0hXk2FM+7c1Od3sgdzjRAtPPuNr5131ieQYRL42uYqK0PjuETX20m7oR5B
OWJT/YQI2RokY0lIWprEr0jDDnHKPG86jacUZdmB2HMps2NpdacXMrmZhzgz
cmGhsx9L16tm9jnNG60v5PCTrJ0bhuuYI0a9qX0KbfiH13VQkKl5Ays1zZbm
XEdfhXRigCuq6Ya7AqjqouF6ow/ot4pp+I/RFSZE/WEfzOHkcjgUaDbRBHsD
I/twnLHwndrz2dvnfWDPhrvsmPLxgNz6xwkkuK6sYs97TFcrnUjxVqDwWi/e
O1KAP7KAZbN6H5oYCm949phgoFmNSu8uCPHCj/tvAuYW57lSZhhmp3O6N9NM
frvYhz5MiZ7EggRwmEpM9/XLx3LfJG0BlPdyFBRIux4hC3TSMLhPbypDCJhl
T392U0pz1qoLiCjqhMV+NAB93kBFLkyaQBwnnTG2B5CvscRZSPE1wAA+yngn
Yk/W84XQwpQNqvKJJAmwtkpBl64yvaikRqoVnUJWldyrS4HH6h0o2Z63fgyk
KT69bs741xAzl8Ip9sEV2qqgOBtfORhucV8rAtberZs2DJnGapvivk7ecQLj
MzzKkEDQVUO8l/IJq83rZXjMjLXOm7bVCt3WKFQDCa7+uq82+gcKmQpU/eIT
2shYv7vwzB3j46xlG/uRGTNCLAXBXkmD0mqnTNNlUWCxEbWwL2o9x1j2BBFQ
a5v0c1iLK+GxeyJrBeWCiDyKUcKPusJcQtaenMPm5AAafQFa9x7uKtz1nQBN
udTKY0wh4wkd84x3jeQI5RSXLtiKfjnTOm0frANzdB/nBxLuTACoUwQILpo6
iFcZCpv0hLjmhWcjX81+Hw76KvwKxivvKLKVKwxt6LAfkunkP47FkKpP8gPx
UYSwrIGJ3kEvX5IUooawtvmMUflI8CL/4V2hQHXc1hi06gpdqz9nk/GmB5ph
k7E+hotxSnaUuz6X50wbl6XesnqKOmX6lZUbP6g0b4bhCjmHA6yDUOxfOg+R
XMzdQCDyw2UJDRSKiFIu+quqqeNsd6xpLzFQMvh812moLpw83sICIOBHytno
I64G1hhjOMamchELHdUb9Woq4AAPGZFCqvpUKaMJN+lxiYRMTLr8g74V2Aa/
m8TcQUQSQVd/CNzMWrO0LDgB/9to4I7w2L+qNYX67F3K/mmwZg+v2GTv4HGQ
v6HhQ/9WeHMwFKq7G4A7r//kKmn2VBAPfITSpK9bipQFL/ldVBuGgtlTVFks
gsavRIhQX65JRoD3d5nf25gKoryY0zlr2rBY6MYC9a99u5T1JPXqicxrRQI4
uufQdFFiZaNb/H4Xu9/RAmsS38kCxOZfdIwXZ2DcnF4gBJ5luaEhBE8NBCDJ
jrnEZMuXMqyenEvzQW7kwQHyXBAX9dELC0WS1TgjP/maMJCLqenBl8olwnlF
rB0U426WxM7bq/sBp8yCRGcGaGlod+GmHfA1J9MCu+XKqLuJnl8tCdNtzbW1
Ga4IOGOQ6ua09AxDNPyMPZJ8Ztjb19mXV9J/twwHpctcnprd72S0q5FytVsY
vXTx9eEcbaSI+z0CAgwE2TkzRvQaqXP6ilNH5yFDfqOsGipLSW+hF74L0JtV
/oHYqlSTpUkF3l3OmiINQ6Uhqq5vrrMVFQ2fdNbQZnwHU/R4Pqrq15tM/Gwf
S3jcEa0uFP/fyxcRi8ejvo1TQ+9kKowYW3ERIQGG8++4as8tbD7cdojJ5Z+0
e0zPXpTLTVCC71ak7RpdKx2UA3jtv1TMdOPU7qbyXsjusfwvKCeDW67T2nHK
LgKbtDMmVk4QkRrrPSNeUyuef1+NcBuTVh/Wa5QAx61WjjRYJzWbNDU/fZJh
ULaPOwTK8ziJIjSm7p4eubF6U0ljDKUQ6MumpK9HfixF52isOeDfTQf0HXu3
P+Yob33S45f6qv1RnfCjcCHMuo7BrmVkmibSzuaZsG68I1luRBUwqUs9sFJj
eQE9rufnNMt/dRrzjkylPFDfIRer4iiMV0baG932MWyQcQuogDpUKlPBGr9a
eI3+jtXr7+tO33tM8tFd9L9m82ReyGDkRSAzBA+ZsTb90GCYHC7LyUMp5LUj
Uj4b3o6Htpy9H2N2uj31JmCJ5qomsVDvn/0Ur5NCHmTh+V7fkhasVwm9ecRo
0DAsPpn/V6l/0HLPav/TME+9v9akW7GkUd8fv31Cl0KHNedTbQeYF7KxgubQ
ONvUh863MsyIOcj6lg9yTUZ0KTHa3awZPvdzHXqXTqQ2exjoSVpYyefy1YrP
s7D/z+k/lD5vCjGtKJRMevmnLpWTDkvhQkcdg17XdjhqXtXO911DpxWLW1lC
+QxUbJTtdZOLHPRyXSqkI0i3k7t4QSxH7DuLUrNOuFaRBXYcZ3Y/zuigRKS3
Va7gvVK4E8XZDBC0Awk+tzUFUJ4TLFxReOKvQJ11gW7BLC+FGGPneSnsuUZZ
KTOQjhO7v7inshnbDQkIyMy4sEt8dLGSvWvxqXPirv9eCHLHWO3Wyr6fWuse
f2f/WF5QbVb+63z5+hX9EfboYR9C8vSR3dzmZ4L8hm4rTwDzWHKtuPPAwVT2
cTwRGQX9ocNFnOH25cNK2FpbB52+uNCZH0XaXTVkBn97U8qmAgbhl2ML0m7r
XX5YeoYXIILHtPmcPgRAXWOYohNdlCWDqxGe+eckSlEnZlarVh1GLPLH4MqN
INNjrhgM7WtgCwTKpxJeuH5+V4Mt038JOJu/2UW8OSwsvheksJpogrV9ilqI
HGzHJmAvuYVrFVRsduE06ZwG+edx74ScztLQ/lZbmxM2Wn/YpUYh0xqrVv0X
YjCTQkwAnruQazKh4HLQock7iBLmYpMjitPzzx2ul4Xejbrvp/StICNTg+Ij
oO45NBUuxDkuxPxIovDz7TbS4ZFtQZbHIzU7enpAuE7ueWAYhMB4E6RdrWgw
YZQymB4Afyf9KibHDtA+7ATXb1XlrWsJtaxV+ioHOIFI1xDmX+cCPsfQpBoU
ZuUX/NEktwTFndIKimpyLTHYid457VQUWZgSI7sWDy+bzIADnFeIDdkLOMqe
mEku6Rsgztvl9+0CWWdnAd2CK517lCF1OhNuitHMdkkNFQmgNEZpYRjUCOpt
PnyXanDXmcRE+MOcCN8V7f+FAhGSPhqGEQ7BxnrWqg2bqOF+j+u/6kbyKq4A
AA7h4FgZorZZt4H+ku1kZL+oXwOIBPMUC8gxwoHMJnUK54DH2Z0RdD1NbPXs
LoQOP9/usp0QcZT8Fp2IuOzN0AeWOin0L4Q4zp1cUVPcVVvr2KsJbPWYArdb
B4o8A2fUx31uqMmd2S1ZhXz+FtV51FRZ12p7BWg8/W/kqkoMUQvhSUk+YNeT
M5ahExHGpSdcG60bnOV5clmhf3+oQ4O3dZCeEdIcpird4idi6z4ZnAGzqUFk
560P7gNzJ44EYP8cAwpOzsGKismw/PDErnsSP34Epdset5aFV4BlDZWoUzZe
tJ8rBK6IHDXoYj39P3nrInsqWcbu7YE5AknHf7nfd2rkj1Lw/599nXasT3qJ
li1wmGGfX3Z1as0Wxj09KLyyS9SBjdx7c/HHWw1s9llA2EZ/gQ8kClaKtV8y
YhLO704sWnyU0T3XUGj/jt9rFKiSPgMzT0T7jqhUUdzGhEiqYu2N5TsRFv3m
TFN1SNVnIkhgEe8Md66XPppAEo5bJ8zb3TuCKzaSgCjIjNTmbvSaJiq6aSbc
j9A3KL3dPZPGSyW4SBj2XosQRUBWU3nyJgie++71UsgTpN/CFljYyk/E39RP
AxmnpPHDNIWnZr4dEOQbH3RaIx12E1LNBe9Qc6DYEEw9h6SuhfhAFH9rfuuK
ANf6V7WqWZHWXMsaTUhdYkEXfrzm6ocWUe7CVtX78NCfOlZTfP4uJsqzBLy6
bjsk8l85DgxW1/4Hfbu0fbv/Aw3mtLQwVC90rGepSHJV08ITnu8BX8nzV+kF
9SKgYFlJ//xVWBT9bPl4aX9YAzFXGt95ek6WLz9/4s4BbwqbE1OVd0rmL+RY
aDgNaeNc12ZuRERqiIDR0dpQcWNl+8syYZ8f5EeWMaqylRiZnI2I6Ffjr6Ah
1AesGkfA4y1AbyQmhW8xZhqxLy+Is1YcBO0X6v7k6l0bzyc5LMvIoXCO8MfX
pofWvVQ1To+G2iQXBAIeQSDLPM76DysLKAsFg3Au1fgcFz4X2+fTHBXd4ljb
wHl6aPHhAozaG8zFDPJNoLJlS5LwWY5Bvv2U2Vho0szZQ7ZE0hc9fkmaGmQ6
7AzqtobeMN+AE66b+/VZ3XregmPklDdBQMMUJe5ECwDZCW3B1L6iOSl7kZTb
7Me5UiFARGkZEnBUkFfSJ6fKFWeWI+prD91+g3vnruBRr6HqJjez0Wtc31hO
EqkULo8VJ2ZJRBdtBFFPlpOOQvLltg4XHp1cUsMmo+4nsiOpv0bT+HVfNTwe
DMmns109FOhJUyNV5QNCLq5+CpupZDoVO17/dP7pJ+4MAMqmRHJu3NDC5KJP
YQH7hbVbwg5akEsaKNhptEpjP6Ws0Ckr4sA29bTx11XmXWiatRJ99lHlrW7u
msmaSfx0IcR8nypZAajR1BXYnJhdrCQuX7F6UGo2if9X+PeAirOK98e1p4Io
PicaXZ+JN7EmqeOIaW6RxWXjZscA/mw6MW/6GBmsLvri3SQvg3N2F/CSyj2H
HI0IMmkJIeXPMFouvSQ2KlR+bMmDX9TjgeVGfKW5TYjDephxCZZK8EVnqZGM
yt4jxayT5KN8y/wX/kZbJ3vPdjkFCPkbUULzT+w1vw6GivTcKVSr8GjFoREp
nU6DtuZc4IrovsyEAEjT8/op+OGc9tHGitfJh3bzSQaJEm/vD3h0VvvM2m9q
rueAW27WlHOf/Ecm2MnSnvTAvPWeAG/jVVI158pndvcHhRPFeZRCIpMAvPnE
WiQse441a0P8ngLAYb5eFp6/gdvcnqXA9OWwNTuEJMUSmRglTkpgmM/oliE/
EhlKqXQerV4m96yH1dzI1NgLOXPwf8s9M67jABa2BrYYXq81/e4nODJjfaVI
C4zDYVBWdSWZF1YDQL7sNNwrZ32m15dusKRZsDJnhe8tM9X/g0PwpDrQW5O1
cBaPI9kTjgUDgbFxHN5xju/Bmyx0hxjIQwJ9o+ZQFmEuYD6WeM98OEevvf7y
d8P+y2LHz4KBZaaqpr2O+y3MeYFGQoK8VlTmEUNzaH6G4MEJEgrv0vc4H68O
z2GWXl9nYXq+CP1/gL+pQZpHbmU6WnWQLag1bzYG4d01qXlCKJh/TeNlEfT0
LiIRsuk4K5FNSs5w2aFKLzbUkHMy1e0SuNMR0ZODiGkqYqg1ICKdMpPBo40l
zbE7bLNFaYbuoQaChziVUv+452hbc1xx148OFh8vwORisjARgm05eUS2zksK
Gv9y0VBmjcXm3izSNZ9Kqb6U3m12ugQE2+z0wb5PlpWBS4pdtzTOrMCfwKk5
Uf6IT5uEDsRpKTJUYGGGMwFoU6hNECGoQJzM183qdpm6zck1Fm8o0UJGunEl
DrCfkFMB+2Rlko0tHuoOGcqPu0F2hks2Dew54oLtUCWZN9j5ieDXFGZ+fY07
olJ5ps+/DsgCB+Vejd/BXF7ds3I5GvwtmhivY0X/uWita7cTVlusV90Fmf2x
fur+GHTkzuiI124RZFCgUlJk9MHI5zMOhFSSKARyHKXSmdr81jtq7LfzkdEQ
udGYIP5/Pe9CURD8PoP3lv1Nm0Yl2fmV6djuN8n2mYFzUhZFuv0BHMRJCPMS
JqKRzY1zMbyjQArD6UakrdTJxrCLpH3QC3VkBZj1lhZk+W9Dm0mzWiMTAzEs
jPeltwxyOjP5rSw5Wp+yTYgNpoXOSjQoHHxGb3xjVea2BLZ+mTMvUy1TWL03
nTr/CCaOMgnqqn1qldgqCfdKSbpN646b+BUHiqWOhndfwztvqvsm63k/kx1S
Gw3ta3/nH4xywJyNk74SiOguQRPxgavhi1XmLEMHuBDRaD5CToI2USKIK3Q8
xGiTImArQc8zdVnfHeey2qbWJnzqa0BdP8GKHKbi0SiF53PWZwoenOB1vVAv
eeHTmFyff5LAYr/UEgzu2TzJvv5OCi38CeOUBvkLMnJEaQffuoLkjA8GY+Sw
6ywGpifg44Qz8M/sCNYSeLJHxHz+sGg61QOGwueTBO8cQbfYTRMTDslu9rGA
SihvDqlTA75sNqaeaiofq1WblQJ9J6hrNhIk5/3sEI3dwxc0/MquRSqW9mmO
67v5KDNmqBjnIMlH+BCcmMUa8fBK8gOkaPN/GOfylL7g70c+xkQGdvRj6Vk/
uK5s7hhuB/1mlAFk+ZNQYatJsSpSfQUjOh+yUKu9ZTh8a6U0hts6iFcJZNzZ
XlMGUlfva61bsxAl0InCtGHqHI01A2Kia1GIwnZwvkOJRD0dgIeEOersedTD
S4LZQ5EZt/AIrUK1ctTQUx5FYgIRGyXDit5PY7dlbjcrgoYDThDBQkKe5xdY
cXMAJFxsU62/T1UnFhZW8IgcAmx2l8Y6cA2QwfjZ5lA2U8lIiEJ1XLrMd9O0
dBLv/eGGboMuFEPcPEeSd2vjLb8Wf1kTN0bDzZ0YQ/q7Yba8v4N5Gl7Rfz17
s1JVm9qvjqp2Q/kpW7MRadLRQngG86Lr/Qs0qZkNOjQcZmcrZdRGkwXzym8E
7/mY2M5seR46qS0XEEDqz6RMWQgkArZq9jryG/KZ2CYqe+kiSPrBabTQyxC9
oGOQ54I8m9L1FebGCvn6dQfXfzBrFsd8iMjwru5sfkSbJ+ZTOb6qhK5COO4u
Gae+MCV/6baPuYBnPOiQrv0dw3a5BLxI2m0jzcZJrBgFEDZBbMpHFzh0IzUQ
YakG1Nt80ELbWFl/0bPmwjGdMA6wr6ik7wUm2ilyJKczxZaeqYqjf22svfN0
CYOFABMnR59PXvdn9RCKm9zoyDAwjriMxWO8I+wcpSXBfEnysn0IvoOMqQFa
gU2QhV96/SnGBPNrcezMtMPiJc3B01elsBJrpLj+osnNbCMncf4kIq3Hgq8R
tEyIzwGKZwnQsHuunhHU7WTeVHvVgq6HhzIBnF5gfLdRVMaK7hGd+r78RRYX
GqZ3Yj+WmUY7su2BwaCFkmXCXfCVXwv0vOCHy04b+Tbj6WDx9K0cp2wOnFuc
mVpk8KtuDCx//Z5rEaqkZvAXN7W4rwxVdxEYvLpo1qMAuY4je42EnqCnqXOv
YD5VtFFLrIoT+3d3sXWlf0Y0iac3zIBvpErysM6ByfKvbHXPbCAIgtXkm0Xu
isBmIt3ibQHAgyUm1Wsuu8TncwsnLNz7vQWtR+6v+eOyYrstEwqXMGWAdj9s
Pxos/X2OkiYSsDRk0DVbJhWUbbUKlyqo/XnRsmylzmzfz2gYjca5JV0fqtMa
/826foMoadakAxqZE9w1KtytDLD2qXq6/wE+myVEXvTCcxQTm1qKI/ca/p0J
IakMqUt8XK/mnyfIpH967DWjquqxVU/dAAzsLqD7iQHJEsS+CIrhBUcjDQR1
8SjlpMn8jyaKYyhYjMn087DIgC0XXH98Lu5JDjiqT/S4r5FnIrNypMHTmeQz
JHLaSzeNkAv2xpsYGPMg0+FSYwSGDv7Wj2ZqtmXOXiQezI6x9FF0Q7hA6q3/
9xsVlZR4Xylg3UAZR1w9qaNtf5x8vkEEpNMLyafOgYwmSnId58YR2UN866FT
9ZP5+973laoJKsiuMIYDNkrUffquDs4UwwVQQctMo1rIXKYGluPCzlyHTEh6
ttiB7fUHszLNJvUThyCoXZXSbAg255OkxDvNzhr7Zzpn+VcDGJVFLMzULaiu
UVKVXwoWJx1veR2b3IFRyzCpoFUONsGifAxLIm+Apc22xWkOlNGEQuk+BRMe
Yg6yv7SLj6EIOOq5fQDKCcc2RXuwmRyEPGvp4AZVtjl97fGs3iNdc1TsKEZT
e/YcVF+nu+YZM6/thzF8NbjpZgznh7oi0Sj2EfsyFQnJw4JQ4IwEfvTY72nw
CwtaBo+BYLUSDzG/OJ9dYI2ctZ1stmkF3fqjl5WeL4z1Lt6887mnkty5rjMk
J9wkWSpgu/mzC/Bs1Tpr/Ej2Qp+tZiWZ51RR403RzpdYEO7N4uAn9hSHp5AF
B1++HPcBXc92IKsPzchZhUjxkvWP9ROrib2f6/lPYnn+lrGi7Ef9N5UohjvJ
/n03Tek3gLG1KOHqrvdJV7zqllabU+cE1dvHUuVy35rod+xq6FrRnS3QMVEq
OYzWcPg+molN61S1d/eEzSZo2QpV4OOB1jPDKf5CGPMf4FEPeua8R/8JMZuy
ABbTnj0/vNBzBHQ9watrwqekuIGF03LUw96lM2LCBjmnZxiSDcwD0wBsug2S
xWTCx146lSWgJFAWw9iRUW0m7OYd8+yOaDqSxPiFa4BaL+z8t+AUpVCcxLEH
hOcrA1mHldoVYr8v3aBAVPlb4sT+Y1qn2/ZdfzSyNLORSFJRE/Am5me4R0+4
XSja4AGDWFypv0T/VVQUmioWmU9x5tpPk66bfHtxMRYUhzJLgeeO6gvsaAWU
h5YpQnVHAD4k9CF7yLuL3kr6jcYzWYRwbs4rD5HgKUxv7YWq3KsRX747rsqm
Yi0EJrhPhOruGogMb1LhpdexzBz5E/Y6NW7iTIh5/PTm/9eSqLCWvvFguc0z
7p/xek6NgtHQTHOiLl1lmtgkC7KeWQnSYvjsGqECwe0GvYy02vQ8IkGJGTAf
V37BnmEGYTOeuBHul4cFxnRDUUY0AcxRARSxMiSxF3qb0nBxa2oHNFB4Qkg5
MWPEOucAiM9vFLAGOJdkQJcVjoMgZj8mN5ZM3i5YTCmR+J0cV/WLlRlj3n26
foLazpS6Vhv90gT1t9qZL2+2reizdRMqJX96AjfAmJqU2oqiUmjD1TTle2q2
4RT4nXg+A7w0NK3WKP7aA6+QHeWrDm8spnsHeWB8AlpkSeeNLYNbOqemu5uX
U16YuSBNi5E7f6mqHkucgxcYYdl4IXUGVyuLqXOJIC30GtQ7bDVN2Bk1xxNI
zUcEsHkYBdcNzVyQfJQ3MQo+9kEE2vCFH8ONKD42nCiBNHyUo23nyf7W14yZ
+rF1bGT2p9gKrB0naTwp42NtrZemEMHqcKHqM0/muCDmo2Aa8cZv2p0Tr9B5
v7N9VDszO8VPobAFH1nprufMl35qgJipfrjjaZUp1m8ZE4bxr/WrElQDS12H
eUjKzi5eM6XEU5jRkQzzmROfGISdPXoGbjf5x12JKX4frDevcBjgiLEjqKeX
B9cpFbs4KLC3qM8XUvS2M6auWytIbJKCUY4j9Tv/U9WhlRDPMzeqrlLVXRKo
6dhGXnoNYZ/KH7SIsyIxuByQTQ9RyulogkT9ghh7vQinlawjhGM1q7A1bWX3
CkjGS49aWt6EKOLC7k8sHEaEu/v6AfV6c3MyQIOkt6r2o1Tq8OjkQH6ju/Pg
tjTx3oUDEVlCRfpivj7aKDfBDF5fWunadwVJTO3YEYNpbOku64cR4l6q/4qS
22WLU+7VbVqdalFBeXvNi+Emtkp/X/JsqV/tWOC7yZIfwJbZjbpcBVvb12pc
jT16WA9iCNkaXgKEGz++2hT744lpQqjKs84/QxvA2HTiIRJ6UNQYOo+6vjJZ
KX/bDjEhuxCDfSAKTWJ5JXdoDaYJQIbwci0zIKJC+sW21lDNqwJxWuoQn0Xd
BFUaqfV3VxbSLepvdsi1EcEltLqyr5/fzM47iGTSCbzEm+O0AOftWnLXl2Cj
zB9zpmkLxV6wuAcwE5DtIsT1wv8NhVc7jxKENyOihrCmq2ykLySSrTIse5o+
HVbYxiXryg1wipo5kovd2FWnQAo5y8Zj7FH9MgVHLx9y8N6v1IChSB/TY5nQ
frjFwmpsP1ok/WOAKZqoLtqz1RRv0WQdtP1Rr8AFw/3XGrTf/jfufOWhWrzl
3vS3tW31SmpwL7UEImfvXf7HRUoGoUF793IcfbxVZrEUzEb2BVsdCuCqym45
Tk1Azo+zxElMvFOL+l5hgKOJRyuEDJK+BBOwHaY+PVMtY5DjNuUSEzY3T/bt
Krbj1quf6BRL1bQVQhcz5HLQfGeKHW5Yj8qT2kVPJ+s7uU0ZGRntUDMJtoDO
eEuZqakxBQxKQRol8okc+UhjIEEiMovEqQooa/ynFQQfbFkEkI0TfdNh1xm0
1v6t2B8+VlzJzhPQbxo8G/xqA5xCTg33r5uGSMn+ngSaqlxc5oddZ1lz97EX
cpIvE6fNCeNkg6E6yxXPMJ2ryXbqPfa9XBpTQRaLEA7TOB8vRWK6MN26pGw3
OlC4Bn5octQsR+Gz6R8/EDA3GGLfs3wVRXCxqOg67X4fDkAleMftKnxu1+EK
8ZG2lodCiO4pSi/XlccNgk9yDoHlYCcOmq42LAPKEgOgiRJI3x1YFY45l5Zk
1Hj+crwVuMsJq4SVxaTKRryFJW8yx9H54yvr2PqrfS5oqi9Xt54R6VgVu5AQ
PGG6J8VtuTThDzKRkRtv8b5q5Ow3OImmFizyHU2JtAnQgd1JzUES9fN4F7n6
Er2tOOFTnR2CglRUW9ArKZCVXTl6qSFb2X5egVN9VUVSIF1NMDfafwkGbwSs
6sujuYLJDdSW1sbCubBhtMWdlcKeY+Bg7LAtUT0H5zkHNfsuVTT1rwpNc9OU
3Nykyy67GV0iQAME8Z4iIIvWNwNnXMcjVoXvHKhYsAIKZKiJaE8/l+/Fvqwf
4RKpwvroAtlWjDIcdhvihgzXhAId/3cWYq77W3iWTZeSqTID0Z15gGcJk1T2
0AV0BJNS/gDjO6syDD0HRw6IYAHaebufVH2YqqUoPNQn975LcGGHJziAUCqJ
Z4YMcFgDy91xFPLgaX3bTJekqGOS8KLdNT6ivrG+DIsg0CgVYmolov6EJnjf
CzPo1UBOsLa15XrASlmMPKRUD7HdKpoxKuUcHAzOI5xCBykgcMWqjoSOViW5
7Y0aEhDWEf1vy7ZFfIVw9ZGlQY5YK1FJ6ESF8pQFdVYufyZ2fhuHImbbQa4O
uaIXiTxbKRESlZo6HwB8U97mlPrVPKktGyjLeiDRt2iucY5cQW+6MkJk+oCM
H8acdu7/hKs/wYI+MRU/UpLy71n751aNIVLDujMjtx0hAqqq3KD31USqLoji
X99CSHPg9mgBx3+ew0+Xg8hOPpAKGKn4QuzlNYXd91P338UqUZ1pvOrLVriy
ab49rKPIktY9SXDRWjuZgLDyvy1L4gPiqr3mPC4q7JOCAbgTjzzW1AyDKXvw
zaXVGd3OuWMIG+bJWxO0cWMuDaZl8mlhNnavslaL/rhWGWvxuwiLNUMtvQ30
gzjJyGhRc0H56nDLXWCS/A85X0dCo1AirBRygH2mEw+57TRLbSS4hV7PuzlL
luC413I0bF0EzJx0AkSHioW8bs4hrw+q01jJ2YyX1xVj4LsaWnV5Chc7nroc
kTBVTJcfj53pLzxw9VOiNP/PpeJeLeTZljizW+NNBWzKC7ddXFX78zNGq1r9
+IT7lZBndOJTNVz7OFJ/Onkh+LW8vJxUO0r68Lq8SPqA42Hj+cuN0JCiHHmw
rJ566ZTf1eV/wQKIr8yIgeUjLNLeKLI7ECMrs3Om4QBWBG8HRJFYkRagSEp1
ThvxpITAt7k7Wj6Dkvh1Kt/5Ca4KnJWab9HH7cLVHTjUbsCIm+9G2LKVJEow
ZabI+6ni+mFV2z4jT/EFx11bFimow2vOhiNgvPwAwRN2nK4EJvoa51M9BAjB
MyjtOZ2egt7dRUPYoFxy53+rjRB7UB1dsakxq05YhgmOeNHPfmcapvYDV+OV
cr4NIAAE2cffMfaESGFvGE2mjmcyEvOtS0QJK0feO+uTVjhL8x32suYpO7rw
IuRXrgvSwd+kHvT4DWFjRaMqZY69zo6L+LTLcQnfquTE4uKFLljC1MQ+tqIf
5RIKBncsuPK7WAL6SHZB1e5krODFD2AaFxgg2dK2pzpiB0uYXVhNJ9YLT3J9
0NqJplQ0f6qo2kzy1Z1z3DAP76Tt8QNYGGKXfes52piPgp+qyW/Hu2kskW+6
OsO56qg0L2UtqOhfgwpOCrxDdxaCZQmBk/TAyG+18p228Te9NNqCCBMhwc6z
eUlM6C9NSFeSPCBw+QMLVsdmUGD1yJi5ybpJ5cS483vP2VbDohZim/9y2STq
t8Vl4fBpQlyYO3mGIZ54747uycIuWWR4hlXmdsdHzPy04+Ry9CvoRq2SJN78
ghKNMq9ukD/m5lZf+4OnalNWG5HX075WfGPc5f5RD6fCT5Kz6D0FvjDnTg0U
WIIs0T/Obux5/svuZi+3nSIvj5RbKy3i+rQSTHhr5/enxSEZLys7k39vWRBW
qmGoYE8keSr93JyP5fbr4oy0a2SLLjuBVG7FP1GZoIJjGIeQu14NnK3MGRVL
wdDIYVxTCYjAnTkq+OFyOVXUVawLCi/fMf/zTEaUT3qnyEFhZ+HOy66BOwJw
CnLJbrrK4iHXJjZiBJ+aRhAAMJ7iJ06PTDX5Ys3e3b1timZTDY2G53CE/ZJ0
0Uoarsi8gUejRd3CmpU/OgU/Xij+sYwxHzCEk7tk4MDXPbgtC9C2R2DyxSGU
eoEuzCeO3VWq+9qkI73EeWTdIfrstW2jxQcgWvDO1H9GiN5aePRci22pKfA0
0J6qxmv0vC5ZjABoWt7R2hJT7JzraKC5V+pnIrsn10uJGMKp54avjyO8Q5Jh
wWnD57p9dREMwQULhgVUB9fbhyDJ6go4g1nzjEQvXnDUoDenQhDdHV65ho56
NdYdqBPpQbpABCzbXElflXMS+Ep7apjHFmWgF1PLPR12LNDFOCl5FjZnQGyi
P76Tj3fKQ86dUMNVe0J7r6QE7MZ/Y6bqxJ9Somf+bNprtfW5vVDp+URe1cl5
PZ4MV/B2lGE+tLnhfEA/4nzR4zfpQWwZ5cWZug0UjyaZuF7qkY6YKrubcu0s
6CW2Wljlc08HywuF4t5s+V5ytW31e8WAop0AVgACGChGFg+cYGprlax0dT6s
2vaiajBiSFcMSpsg/egGltus7Q5c+glkhabx89wNBScsa7V6qp3lR3Ky0dLV
rZ4FUWZpWhOnCqGU2w6g3uOwlA3uCM/aG+2MKpxJC6Zh8xV1So2X7567BV0L
F7hN5v9RtNIdQ1WXC8JweI2jGTTha2+jB2GEvIIc28jebWTc4X/0rOPQ2K2I
woEPWcLpRNWx079ati3cUyVKMsFRLUZ5RlBT8dnSQrG0qJN/y+WQLFEJ3ZBg
gRDgYn4wh5ngl+lj5QbjrLLu6nKyiugnIh5Mpcoxfui7ZdO+yIl+Yj5AEIYC
AsTmrnTHZvl4fZYQI4ULcmdVpETUI+c4+qRSU9vNb6dYwifEnf//cgSRvzci
ABraY70i8VJyhiTy4oIw1MyFuthJVXrjONkcRrasx5PVp+rBctQNswSad7lv
M+iJMlwEXYHWCsuwzILWkpeA3O4QXKrX1O6wETOIK9bFfK5YEk6rhXIilV04
Fj8O2/DIy77UiHCyTuJOWSYMBC429EPasFOCJhmvBdQC+gPPeKctS9EXo8eg
5p1dPWWei/R2QIVPy8SVKvAC9oYr430q0CTh5ZXZzmpY1e/EZGHHyBeolbB4
rx+w6JDK2dlFmOxmDSS6326WdhxR0gkX/okURLclwteHvN0iw/Ea+e3hCEDI
kGkYER3zDtfozxHnoUJQ8G1o9yCO9xUZqXw4+xX2ES6Yd3emVz6vbOG+5IFA
YoSVOl2n1hd8LHXpZJBOFpuKOsNGtLCY2fFkw8hpPbie0m76ww1iNkicUf2x
SFzA4TeeryGmhomVYTqsZVTb/jOq1ITZF0/wsvbfTe0YdwzUUy0WRD6Te2kL
Qs5LnZpXr48gzWrY3ELUNXbEb5u8r4jd1bFJcvrV815/D91ghkQrFe/+8Mb1
zlyxiuhK4kWPrIas+7AOhyy9WQCovwr1cfm8d31rCn/tuDy8Wrek0Uqg4HUs
Jxih1E1uWoD6qQI4h6w18nOS2YXX99LY1pvZgB7vpKkc6twUw+E6RU+XSKcD
B7j+eemnBkaUoxJXE+fNmB0fWoDokt4KJJkP/xy8/V0H96Qd/PTrnTfaM/E5
oYW+cMtGOcwEzh/7aBLf8duJLtQNgZRy4XfdsZA3T8/ka9WKyIoW5vSQyHPL
XuwIDYsY5n9JLh2CkRpwlpw+Y17iKwLwKDku/RAECHD0rPsPv1GXUvyIJnqD
UMSRhPUiCpKAttTJwZtyRjTxxWjOnedjq+KHFPqWv/k3hAK02BCjHRN9A4Zg
k6uihpvEgTRxAdMV6rE/jXR/6G2krp6bgC0PtuXsQFgXJqJmcsmTMswuEkW1
khLgHO14xbcwbBvt7xDBOD8kMgcTHhTN6qRfKcjysL2dS8UQ7m9c7frFXMR1
Vb9To2uZjxlpRdQX5QnnToiM/QgTOoJdf/aG8M2nhOgozF2oEcR3wFwqlnhv
H3InphWoW1631haN1YOIM3L2M3u0PMk6u4mPjgz9EJqp+gCYbUC77nfosUTB
D8ZcLTJLnHln33Xs7mYCThPrdM+9dLtWb82m8RQeRMhHk25yx46w+fpmVd9j
+IXW4OPLsWvTlQmd+nH2000CYT0eFgk2Y3JSa69m6ctoEq3H9bQFhcd/2ahF
D6rU03eZgH4JKi59oHhrbj193mvHh9yR+uUSuwk1b4W52xtsDS3u0uC9H8J4
lRy16prkFpFWRrvyoWU2am2eVcldXJjPzwYczfdkZANL2QEcpJjiSeRKs8w4
Oo10sBJS805f4x7HJb9WKKBoyBiuUGZRLpCuvcMPaAHnEvowMeZt/eOAt/a3
sTqcGuqT5DKQavS8TchtSLGmVjSDgOjBLMimJvTG5k8G/taEapn3dtYuRGtK
OlOSO24RqGKS9zUx3z8g3trhcyFiZbPgILEHt5qkAZ78tp9AzHvG0BV3iBto
u+puFtH+pOMGsix41f7jpxrS7/ejndv/WhYANZtP24aOvicmGN+4oHsw/pUu
RG/yj65sixd3PXFjdIsXDhc83w0TpOZOUH4JQC4GDppUQIO8hZuoCMBnhLjL
8yv4EvapoRrofrvQvdJF3pX+YsCvMj46uINurBoaU6BPlG3PocmvxiIVt0qP
gak/d9BvBar88oi/2y3uQLKFuzTuK/wsOPW2CfHQYaNvaHWbWGc52pAAM551
4TTJgXiAauOdRiNF5RQcZYzbBB2DhIk1iHNLpvgyPBCsCujQJJDMhOU/JLxR
y4skMsijrUio9AOPe28emMNs7s4LwSO6hWsW5IrPCMqfZIuJsl51bH0bzlkA
LVkqun7oN8a8LFcgNJWbPVKrDvWxugQQgobgKK5efztlKDSfsoW2zK6earCw
/RFyPTeKhjgEwSfS6p3+PbeqKNRfhVXLm0mF7kWRzt3iqeoz08YU1xWyZ228
2RF2U/sWQk9rzcEA5PScaRB1B1kqAvj4j4o6L9rx6/Wq84gCUn4KAtq3dRZM
r0Z5XXG/vtvrzSwRgtV8xl581WMZKglFshFnPG1d1eCGZIe+Hp32gYaHyjbs
rfISppgqgdYe87c638lAsFUTPk6a8n/gZ0bViGSmsqPyjqNUyAGgv5dO2uoy
saOASKg3PFw9HczV3SBR00E5ETO/EwUMjI2NrkY8MWRc9Eei3sytc23NNZwD
/+/sUMbo+D0qc9vxgOZR1eBzybRY4KqqRDKvct22D/AKfl0eSu4VYFMkbENP
GJzQm1KOK7hQ2zG/hXVhm7afFp2SCy8l547FL5//FqWR4EEmbiB0Y/r7mbr4
zvIv9gw7RTizpHVoDLiADxVBYU/nx7Yrq2valb1l5v5+SU0+joH6TInHd7zp
lR37JATvO9vJ6PUjXtlXaJCH7/kcdzBa4dKPaUGgVBCsgEEfdyQYaKnfvUfj
cPzd01m/LNVC60E4J/g6/tUDTyOFLADtTArIEDpOm4q5AgAuWyOQLJM0AjZU
DZIcC7/5MLXDcOk+zmq7+1184yRkOdhpAVSuUEYqx7CPZC7DKGIh1wqY89V0
N7h8Og+eW3y3Fi8FUcIfBX+5tugRNDpL5sfUXYxvFaFY2FYqf69uYycolZb+
3913HHAzZUGWt1iPom0C953hy+z5ckgY3ysggUdabP34+aFH0DdgSr0nL9NE
1j5W0xEhEAiPomTSW/n8HNh7Mkh84Xn4Yl6VO6okNTeQNGzY43QnUcrB0bog
3MpMdlID2k3m4hpUFJrpwSA4uF/TlI3nbBHPzFO9jCWzwnG2v3MX/3cVWmVa
xWCAGX1Cqpgob9mtUYgvW6qvihyDPp7hmunpW5wmemtIWJo/t9sI5ESH9ATU
S8j7nbgvUdiIy1SL2qgXFsPMDotKRSGAniketmeiHs7YJBWf+rjjoXXs5lGl
QCIEWKtDtfHL1wjq7cmCd76p4VGDgojaHTlR6lCwD9/cQLsPzblyVpW+0Hc6
z0t8PufVGHrgfX9B9AbBnqzQ3K1/JufvivUPsSt4FwLIJa9GWomO8o44LJTM
XnOB+H6kuzQjXnUDBgWDLQ1M1PVWoK/W+znZdlKZ2ryCQwuVl3cKNwCJMx5a
zFDNfYg0ueSv+XqUIwOQPodsVdbwOIBNea6nyb8jD1TD2DeMzZnV4ES/6xiG
NQI4mQIYLYuk11gH8X3u0IunfqXhGQcrRkBV4mNMzpTPomm3rAwN6QkfCZxn
0XhmdAN3eqzw79ePikJKMgD2stjOA7s4UXr7p6/hJ9C7u2lAVVk5F6GB+KIk
5RevCZ+j6S2p0VGwztstJhjhHL7UhM8AXdyJccwCb2/xFqjxpzjMgVpNxNJn
dujpQXhqyy/XvS7atAFr1TcRopk/iCgtBo4vO9mgRgSg8xaDi8cjqmr86h+D
xVsd3zANtjPHC44/9y5s1tFwiaameLSAtdgy2bZX1oL9tbBEa6XG5tiYovGw
ffNz76/QYlcJYM6sP7dha5ZE97C7C+4AmFgnEnKtgkAy7a5Y6qsb6XKhbjdQ
V3u6f5MMb4FseeR4+stHAl1CdiWHpqcg9sAJdneeOXsDSvtl0HIcc4wcXgar
lIMTkzuTvvJ87ZIurWCvt5lHhHX71l5wv+pNsYtvYjluY2F/eTn091VleXiH
04aPjHuuEvpMz56H5hZNycbYZXkG7B5J9PH6Mf8dqBGhsdW5WsiRgDmKWUGq
xxx56mx8s6WuHPGPfJM8MgEdpST2ti64GRE30G74ttcECqRlMeE//spgEnhm
IU3BbsfSgQJddESTuUEVvypfrEYH+MuHLj4f4wueKEmYrHXsm6QCX+KD/r+O
DrwarnU/qDVvIFROFG0WBc5LW00giLBWX7Lw6oDJA1QVY5/8lGnEFwgqhq4w
ScoFuyVX6bjKC5G1SwasYPxE+AjhepOzLIiJx7hFWDwEjBWVqxA2arZeTmB8
OLf8spagGkXPOYxob+/W5FuNG2gPoO/z2gSdMHhAxyqn+kNQl+vWqvLq19+M
wWBZFP7s52esvbpGjtEc4sxX1FGiYgIvqC7hQrf+DdTl4ST8jHvDoD8hyyHl
fGm4sio+Wlwp+piAbMIj8lZvU8pFTA5hCWPqwVm6i7QcZgz8AmpmLBGIj8WE
h2/ZcXjv0q2hhfxSKPda5l78rf3E35NmDYdRsQjUQLQL8FrRQvTBYKYdSwVW
/mw6nN7Fdkc0wZleka8/ivoWnmWdUR7PIcG9RcXLj4EVlYyPfWeHgif4X02G
43WSayOIMYcp5Rr0c3WYPBF2m3oCHkcn8NXCGHbBykdRvQZAbite9c9gxVfH
T4tsnlZOsgaTdsSfhDuuT7gUhm0M5603F5PC1dw9HRT0EKbxY/0EwNMgngvq
rq87chmcHJTlo7TLATm4FiYnPcXPvLWpuLo/t2Cr573+kTkF7dMYXzq+gV8K
7t8wbSMUo+HLPobBwptW792klb22aaIM+vrRjPCdruI6p4GJne1mt3JGuBes
xzcWCLqXM7gbuTE2r42hfOsSewR00X9JvMCMetVXrkfqrjvX8hgSi9uY6yqy
U4NvLEcAWMCSZunvjMxBFWacT+4EG3PPS6FVNYiD1yxzW4RtpqBpCK6EcpDo
T3oC6u/QV5BSLuHtwY8cCSKjXBKUmWzUicpoNvfLNgA0/i1ItWDgxXHNR4dv
oTC+GtKJnTFieClGOQdZJ95+M6jh6qKa+TidjjgQUHv+Gb6swsz5f38k2PU/
sAu+KZiGmnXNdDhUS9OuTxy4WM4xU5/qR2uZfC1resHGm2xN+3qPLgrKqxxt
g6ThfBAKrC4zVZEPTMqeDsgYquiahCQvqdicMBIFFka0zD4F4LcHF64NcLss
o786fLAt+ByCr007lv8o3nG0RsFwxJ/SIQiX/+YnCzyOoquh7QY28UUMGLw+
LV3yFyUVU1iR1ifb+LUiHQfi7BN2xL0pb32cLU50e1jcMtBikYth4Cj/YCwD
FbIzLFye/hloHNUNZfJFvMuiO26pQ9dMZpE6JuSnCDAM8AteDWmkvskeCq7s
kNSnumgMmXUm+WXIZfKnI2BkAiXB6zjq5ZwwEymUZHhF6dSvl9S6jJ7lSaP8
OSCpSWIrhvjiMZuZh6I50Y5C7XRMvNqfLYlRmfFNiJzjpN+ltNW2X4xOjZBx
CoWxHIfwz4SopVDNdIWOjDZZYKp7vcd8oQ5aoiRXIubOMLMX4s5xZ3Q6k7Kz
rc9+fQkkXt+2QdCmOKusiDTws1XgAqAmWvPeIH4nbxhwinKvJ/O3OtvSRZ9/
aXwpM7wnXFNNVAmgq6IYA5CfjsQQLfChUCOg/MyGyg86W++tJE1G8kdSmngY
6cWIv5d0iHBdm2aKPLI5wsYrW3dyzqfvxJ7/gJ71esPnX6Uqyg5kLytoXUoO
DucJjxQfwx9g8POa/2aNmvl+C19A0rgRIwmjOAjlyY45tJ3lCMPsRR/84fRD
QjYERBsHAUI5iIdGkkuCyax0M89Hl7PuDUXRqnlCHzbjAcmmz8Q9BdsGnvB6
YDSOu3w5LBKI/AAhR90VHPvHZdQa35SgJQDKFH0vzoDUKKsYJGLgq9qupa+p
FSI+PYgaG3aWw3mVkhTyrb6xSx/5ruSGHAWXX4QrdKJ1GSNs1EwwTTmim+vT
WShiTwyJZbHyc2wqRRlYLFqQUtE3bq6GarNf/3cqQpvaOJhdCdtTIe1Vqbu4
2gv9O1Ff0FtJMXSEh77HjHvDCqI8CPPXY1R1xGDIKM+QXYvGsfHIk2Om+lE2
7bsVnPM2JSM7LjDog/Rfh06oGCMd3ewZWBj8Z9OHAYEZqTtTNH4LCNeo3bLj
WAooBgRyQ7gupDzu4IPAAy58gwyI0f/ZmNV4/Og6RJ/cu3677vvAc8UzmhG6
jOL9T+1RvOfBjBGJ13ODCBwnssNEEd1x4ma8kQiABewegEMeODnj0SPcWV6Q
DkFFw64xmtZlQR06M3UQzrcZO02jQywhAIwWV0OZv7cC78hV2eJQyJ2JRU8O
FCOd4WYFBlBdvprxb51ntxgdNMdGwpObIKcO13eBkm08a/2raSrb0wUNDzDb
G/1SPa7Wt3YQjUq2gOmpEQWPjmz5qieB6Jqwl7TYyIs0LQmPvHeXOyCte7Ei
51FMuA8N/76OE+2zikSTAD/C+/iMSBByB3/C+CUcy9cZzaGR606uMRJJI2V6
BvduK4J1LSQUXFyME5gZMdvh9d3wOIcjpsNsH8zCK27a13WO851RuXGKx+Ia
hX9E7UFhLAM9dRYAyuTzvClq4VVmf6HxVKmpnKjJaw+bOa8Hrk9GqWTQa+22
tB1T3jSZPmAHx53LC5nSUFKI4/cf5ZN5v/EnZlsbiqLhUqio6iNefLAaVlju
hPDe3nDFPZ8eu1lE7MOMfyZPMF4JL7Ur9a0S4LFNLrDafoKgaGHL1NGjcEgB
BC2KGMKhtYl6hhOS/wIICTSX3rIYIcVCnxN/E5UbFzVFRxfwh7Dt6LKtCqpf
TFRR+HpDL31WKWRYV/iySZXs/bVfg9m6cfKKZxNTVrzzvFXdqdctBVbG3NvV
iTOCYCYaJtUPIjVD5NbMbrH6zVtkWdDnjnWGMunuvnuluD+x4r/7mTkK1tQR
Qo72gt5M1LRk2twQ/mbf1qfR8ue4DydtUIp5zkS8e1owOaQu4ITT4WYgYdOX
wCHa6/sp55B5aYhxN7zrvKwE9kfPPnNwVlPzLEJQdBDU56BCV2xZdNwsJvCw
kBx4Ku9FmNabGeel/UO8/9ss7RfHaEOdYdgw1d3mfOUYO2yKp++uPlKO+icm
s0sJ2CW1fAw3rGWPWlr2zSBNgY0Ide+OPK5Y6Mn/bpzaZCB5qhb3xBGbryq3
mFWgkUrf9EuXfcIz1raafxueRmLL9VQH0ICL4zz2qkDilNhpt3DpnS8uFdPF
z9laPC6pSnIemts7DV+UOgigcl33/99C+TnkYEixPE2ijfFJdPsnyKLNWg43
nBYtGhmI79tSPLCBm4pHCnCPhFfvyQ0rLsKZzMf25PRTGwySSIIPwr1SuZOj
TOFRnNPKnANvBgQrQX8qXhZkzWj0MlVJ9lcg8zTM5fSNZWbJQfNwPIHrn77r
wMrKbf6mz2BGI1eoCZ27LyB0FbpNs9v8blVgED5YgePrBZ4A6cwPQTcX4QfL
0ccAgatbVlttyBRUJilx57+2ESOfL9V2nmRGp/6q7s8wHtBe0J75r0LpDMVb
OtZRkZXCP9wLIpmP0s46fWDEm0RmuiPDE62s+05sPbcln7hjlAlXHq+X0kcU
IVhdbBKfxO7+vpItNMPzSo730XlvmSImj3jReGIdZmTIFvktmKsQN7FojJsZ
cC8N7jBWbQPROR57RpWuGCtfDFEANv+/mm+QnkxLrycb/Ir+NHZVY5TrpN+Y
vDNRzS0CZZ2U5GuAp9AZ4mzwkt1yxdrUCP0NAoaO1mi6sNlbKVfmZy9TuzOX
GQ6cFOOCDqz4rYmr8pyRyl4wI/VVxDXdpv5pX1bP/DY5b33U/sIQvfGDhwKz
vnVVt9QDRWK0nNwSplC4u2SAh5uXWOUH7lKsE9q226pleDOw/oOdbpj99zlH
m2X+zMdOkxFZOobHBx4vnnIntme0h5n+3O6u8rzx1+ezeOjGdmvqAF0R3jeD
tpgLU0p0SH2paRUTIUU6NBcJ66mWVbaftVJE3H5b6xHVFlNJUzzzZzmuKmK2
2jl7nb2UDMvfmAIM5jiLhXv/ARaOm/PDYbx/gg3HHo/Wm6QcNWWVzSMUSybk
esKVOSlIh5FGnyOjK1P5SdVwGKBc64fNi5sMEluRYlhhRPl6V09jZoNxeDaL
WWfEAJdl7Vbmfzn3ZsmB1MgKndS2kITlzWTc2siVR4nrC+qCaHrSDtHMnsQW
oNOOmWjOs4l8uyR0HB8KoD1F7mGM4NKZMHoKj9oebZvyezv8tG0iLyHZJ9Dp
cV5hLOzqEIST6z6bCCStU/lcrC4UrIwZfIgfCqBEXgUdi/rNCulxItwTHQir
53CRmVeuIt1Vi0+9LgnmUaCTNGRHmM5+N9V2vSopADTLcfqMdVqCiOVZZVeZ
m6gDJg9nayfBCIy0vgW2vTKVGBGuxFRJtSeP2cT/knVEfoHvk+mG4TevQNVx
QBrIUL3bvwTm0xZbLnSDlX94iQTCgz0V3Du6EQvcCMjvYohdIWSnbCMDKOKs
3G+o1JE5/TtGGR42o4ktpzhcNEttqKlIFvGHGrKRClKB2AGQtLPXrbRvBG13
SWG1HvooyJq9TDCSViGPDgz98mMVOqU6FJB2Kyiz52JOEB8v4FxFzrZYMjfG
FpsG02AYra/JPn+sGbycfSd0y+viGrV4T0GRcjSFtK3V3g2TXeB4yUFiK+eo
OH0NU2s+3a91SsNoiLaL0O7ypU2keUvq7iFFgNd1kag5d6MK7A/WDKmILD+3
ODXn7+hUiaoMnqdHqGNYGLr7OofOE58cAbI6DMUW+tv68GwmsYDj7hVDGjW1
ev5lnm5nPfYcqHvn6jfafQZO6iJcmKDZAru9aD1aJwUBz+YGoy0Pm7WUOjCN
HKsmUr59recs4otcoqYc3Xx3Gw46l9nYjeP6+seu23MMNstm+spO22xYxJQn
oc9YX/wzkiPJyfYYr08b3AJcspI8gDUJNAR0xBj3Xl5nIdB/L8ER0tKnrHSq
2GioC1sOvV0RExUq2YIOQ2CFlV49V1dFiUqcVpi/B2L/aQ9UJl4jjSHxI359
6y0BNU0mb3QvCUrCkL+bQG9vzcOUnm2azySj1X7531L3IWseuYZXFycMoxTu
1DtKoKGlc/YtB0LN5qv7Lr00qkY/CYJ1gZc4Yxf5cVqWP6Xh5Ur2HkUH8u90
hOypBLDpqA0ZwGzL3qynKwFKs4sQUltN3bmhdQmecewyb6fSKdeGi23L3ctl
pHtsfoe4jfe3mLVW/MPPr4gr+TBZLzTH0azbvQiMxY3oD5xFTDWiHiJq4ddP
FeBYMRDudZzWKwjYHXMrD7uIk09GDl2UyMAaSAdHQ1Ncr13O6uLb9QvhbJEx
wexHyzxess6NmzAZWBnPpg3IH3XzcdURb33eLdLgjajMNz9ZdbZMiKjW9Shj
UL0zBKrheWJvWC28BPCD2G7SXmI6E31qyTwlM3axURcWTOaqjMUwBZvqCZDh
ilFxVZE28um3km+KPZwZJQGyZalAYZ7P/3TqIswpwRkRqUlJ2Kz5/qPkrWIz
AKj2zkY6g+2XXw+OstLULLZIeqT1MUYPccJwggHlH8V4WrCrJSfKaenhTryu
DtSdWjk5w65q7gauJALARIK3cJIRQgg5EdydnhbjnHaJWWXVZ39pF/5vMTcv
jRntbxAV5wGp5qY7EtLoncRZyTU5szqykaWWNgJ3HQIkt5GrO4mBju2tAPHB
EQ/dyWaGUC2ZylgSMNmwNPPFsy0GhqPmOONlLpi29yYC0gUISU4rlWz9AYkB
XlNrNwBXjyrratc9TFQN1MpznAp+hvve7tudgFEtuP2TWY6NCs9sC629D32Z
HC+WdsxclUdbYTYGY6mAlkKJ3cCrN+7IdBR5UBTtdpK+cFW6ctCBJCngQXQY
iHkuNzScSmRCKC0MgikavRNECwls/BPhDkKxzzC2Di5rtEjXRTPatlMzaqOd
MFUPdtvUgh++Q8kUIU3NjcyG2X1evJaMWoQ2mUoIbSoIvTCCxAlJOu4E6eKE
6kq1NGh1OEaOb6MQ+PRomjbGhZKUevWauWmWASfyxKdPpZd46CRt1p9dstuX
W+UlGhGXgOsZ9QP4BJ1vYma0p/KUwldiqqYv06F6GkB2f8LvtWcb9aEUw46G
wbBbwLhhlLBmVA1PfuQvPElZN9ZL9x80bhUPZKHU1SjndbYmzvRc1YLKM6pG
oITFE0Q3H2FL4Dvd9oFomY3U10N8oZJPypebKeAvMzGizoiFu6kAmtBDHCI3
u7NhxirNa9d6ijTwv5JQ/ZSBKvQ2bfeOUW7AQMPo4rNfZa8IlJc/Rs2Jk/y0
6Rbu1/csf+lMd89YRO/SrlF2WmYj/qMYPcMXX+5pBpAEVskj2mLX7FrUa/rp
QqC+CwzzrMW/Wh+JCOjvGOJVpjSb/1GbKuhkl3cWVZc7Qyh3eEOWduUCHL5k
KKlFlLeJEE7PZAH2nT57D6keQQ5AhFS316YtEsntrS/BFrTum95L5tXgSn3d
K32D1F/ZUpY1OvrdXrDwKTlkjCstt+zAv3LjMoOQ0InEIzEqCHtmGW2K10Kl
vO9rC3f43GVmfbsjj1Uk2tYxvauc5n0FhY9IfDF9SSn+0Wudpkf2CJqZaPN/
rbd2T/8T31TVzVvI6VkcpvBx86rrZsdRioBXnvrGU9QWWoJJc4HPUyMpcyxI
gqtZPypOVoPmAskU+eJ3Cthr7vLVcSchoRXw7sbo3STT72MpGHeGdh1IJbpD
ynVcEz48jD9D99hEeK8PTz9sxQijw/oEOXzPpD90VCY3ZZKSJmOe/2GOnpEt
e+EVV8kxsZir8pYkSnsiivAv3y7vJX48+9OY5BQH6qOkXM5VPlrkIiVAbBv+
a8ixcfataA08UFjzYJiIaOLyRxuszU1BoW1Y58aJT61SXbSfxZH/1SYyrqK/
hHzHJMndIGz+gBES4dGGYYO/Q0f7wTBAeHLwITRHmCJj87q9YoNzA/XvNf7g
afhhVLiDHjXn6+F8AEBBMjHntG/OpGwYxP3h8w+cGt7uj9WGk9SNbIyeYfdB
4V8Ub9Dnxk3GNMgzJuzE+rUBHrharsnwlJNsvNEUlxOlaWtnqsDyyNIll2KA
tZqbA7FmfJfoXQMGGO+wotab/CQBNH6ZFn7zzHRcAvF0ZtqnH7Ll0+QP9Jyz
ttWZagpQH3BFUOfUgeG7PGgOGTW+cLKhbv0F1ZeKXi3mtN5DryRnpbqAbeGT
2HpxL/A7CNO8ioT0h+GDivEe4EJwrew0jFx+6RozTn18Wu50EhvQezVcyAwx
nOGzI3qs7an1vPvpiEKGCk+uAhjAcj/bYvZvQm3PukyEESw5j/JfhJ/g0sy7
D7ES3DyfRpH0w1q8127mWrdvv09v/CGrGx8IhCUoFCx2LedOM9rE/5T/c8rL
q4z3WSKIZZtV1ai1EuiPFirwt6gQHuTyW6SWOz32MaNVo47Ifm4X1z2MY3Ra
OKGuVl2Fi6CHZEoDhU6UVuwuHFnohJqltzgPmre7WhZ+vwSkQDz8y/qdNSeF
1EbOpyIYSz06zdBbWLUyONydD2gXkunJtZwRNHeGZKnd/ZL2eUc16Uuvq/g3
dp0Q5nCC5D8xXe7eI3KCVHii+pQWbrX5Yu4Rvio/o76KSfQxGXtS6Fu5BD4l
KBGrHtrVIltVktuO/XUs80VU4qC0KPqYIikQooR2/O6XBwbYWKXa8MGAG1Lc
SJfCdsxc3poZSjO5tbT9jqF3hYuD+kR9z6dh3z83CcaxWrsZsCr9aalf12h4
K5qx/XZaW+WKQDflTuaCszEX3+7y0aC1uLG4Mzzrg0yBQ8rQzhCXIpZFG/1S
V8a8enERPXBlAcsiX1n2VxhoSFkPRcTc0YMp9BPAYoC+zNwKXfOH61OMly1m
T5faNfGdb8HAORm9sltLMwBV3ICEcHwakF/xV+NPUrP7qPBUOhwTChDEsEwb
GM5nnpnS+bZsf7/SgeRXYqJ/wLqFE/sRCvQgbo1obroOw/n31t5rGZruB7tN
kD4iZMAwkKxLw0Dl10swWEgBPCqdU9QBkDYrRccqakOX3DUHIrqArMhRIr5H
B4cUKm6A1TSOLSuzvP6RDvlCns8snizHgL1MwaECKLtR2zI7eohC62ap0UeD
X+UeIOy5R7xPJgyN+N0TwhlxPbH9GtdLgJVCQWwCUdIRgE0fPRWmND1Zs+9U
eKfOGTNArWVhwOxtHvVk+ou7OIFUeOlZ9htNX9Uznn2j//L8Xswxdmrx0mr5
xxearmQ0iZl+nU9eobPay/3K9iYQwUSsiDR/upXpSMySB1fc7suFSGhpw1O5
0jyc38JoFRflNzfL1uqZSiFpwawdcs2gcnPEv6jnD4KuLyaqv3yb1FcpMXKl
mCTd1P077Oj4XIiDRCUOpLs6iRsd8ngEWALIuYG/8vzFqptwSFb/mqWqfjAC
k3BJY4qaZ631RDa8f5UrlIoTVUlgDOkpgpS7MOKnJOLicqp+MxGCovHE19JE
xHogAZGhddwnMPg5+2exb5wDe6Io8HjS4cAPhAGphxWRNVjoDk6ImJixhWub
CE+aRaxAJ9AKEBS6jGrST0U7DXOnaoDmKxHBDN8IfJwfWwKIPdE/iNoRS0Hi
LGY3J7M3VXPFKqHqHUKg1GzZ+z9E4FO7ugNadx0HVuzPbPLrcmbzeyyCBaCD
ZysaljLC4d8NvRcJoI+StAT4XsckAQEiIBorgMYoUdZGf3Kz+PaN8IPtcnVk
OjKKCyfEqn1GjsrO2gwM0LmNj/iCJOiaTZnVbNW2Z7lz/DZPZCChOUmtwlA6
LIL3v+UOEXjTfBaUEflmuCGJRnBsW//w/91yNe6MZO6utauzvzD/8eQJS8rv
AFAhtoHpn379VZ6ZVdDH84CAk5RLtGr1UHlEtVmHKIbBwqnMV2sOhpe2xCtm
Iy6CcpudMk0jtPlMsdxJgPcNlAinvW3CW/KeOqTdPrKeAOuDyxtI5KSR76Kq
5kQY/+U/3ewsjrRWEMgPVTVt0x93ozo+jHrtg0Y2PxqOAYFxwYEjKLKwaK+L
959Zqr/5VrAzxUaVulqLaCm0keHw9sBoll46dwZD0XCpSnktQ4fOo7yJJmRb
xBnLjxJN2BH5jIoaeNtzS3WlgiKZNA5RXxcN5oteZknDNI9ajg9ZO1QEqvbQ
jEuD5i1vP4KcPpuqg4ybbMdzppk0hckS1r4NNsGWyxU8qRWA9lubprBXX+t+
CQMP91kJ4W2gEE1NRHQRDcAzkefMfkmug8EBqovzDuzIJ+tH2xrYDiHv45w9
ri7oGR/tx1tZV5G5C4h8lFsjgxZwwRpEAGWas0G9CTIsxpUkCDh6Yi9kO6Fc
NKL8zLFdZvjNMRPb4qgDc2kRck6TDk7zJsrma9v2WuPkqnD20tZ+xJRHg02+
IhcIyameYAAWooo2zJnHBno7aZGciSFY+Pv5ns6X6o4p5Fbtt7FFWeWQocdE
DvqpiOu+9GNkmHsI6a5v85S8dmpUZRSr/N2rLRsfRGFHZUGVPQuBU/kywnfb
IbVpuuLmQeU6SeQZindndvWMG3K+uy74UzN6Z1TxELBIVLh9mqfVJUrYbKou
Y9PN0f8OyCGGCCYfSh6bkZaLALxvNX/tajaUQ4RzyrnOMa3B3W5bDWuJ1vbg
ybzSEwKVaw+p8wnCRlxUt6fKsmEGFv1C9Q0uHGB6GzgDpg1OtAeqAzsv+d80
BhaOkPxtGxxhjqAsrE9EIHn5DLo/Mx/XefWy6Dypwd81Tevqkh5S712fDCc0
C2iKFKT4dv0i0GnO+QMxL9GfD+PgcgJmYkZDXOn7gWJdGZtv2a5SfX1lcwTx
dnghraid9wuV3rfK3UYayVBUVHOebSaToowtcmMSOgTmAGQbPMTL5EdAS+8+
JryzJK8LcAaQ/1hIRbiH27TaDvR7rQHe5qnKXiztGIOhN2mPzGmCW9n77aDk
/FV8TZLUde+2daM4rr1SqJcVomMG2zZ21oAtYx54os/jG71RzuDN1a6nPBUj
xlCzmuzqEmAQC4MRZxiUwIQ02rE7j3kp43k4w+tLu+t/M45yi9Un0V1e9TWT
BeonsyF78uOenDQVpz3uPaeDqSQZ7dAyLuindFqjcJ0VwruA/ci1ZcYkuh+J
uxpGYvE7NJFXkHoHz6iZNXpOsjV4DDyD0SGnqORJ20w/iIx8qAtXLP3cs/E3
I6WzZKGPCadc5RzikzPJBb2DTuECRqlBP4sFWDdsg+JQAFeFpB6EhKEOnJXj
A052lDfUK7l/ppW97PyTDfcuwRZOf59jXdv7MaY0J8eY/CZtJyK8ZqigTMFh
Q1EZZV91pmeUBDotQd3KzAmGzVVX4OFHMtqMsv3u5XN5t9Mg4CE8UHLJ6X4O
Z+ZFFrOgNI/ykXHjq3o3PBQYhEUfQALnlCw/X48iNs5wwIIQY6T0Hvo/raGy
ycieu3uQqGH3mUOf7Kqyg4rhp+nBU1g9xWrA5ohs7+X+xjzHVb0BWg6w8CiU
SKW8XZzUFkfDuJU7oVKk2IBQc1w6DgeAHY785yGGCHXBnM1d3MvCcLwiZsV3
HKvRSGCtG2Vn28jJwCrHtU70HZpZOg4Imb0a7ESjEatVT96YgUgUEpv9QejT
dXLk5ggpkBvWITrXx3X2lroQUuULZfdEjH5mKpE5+UGVAHK3ZBRkXF33nEKO
UAMsLpn7s/XMR22sD7QdJHwKbbzsEypUbV0wtc9rHcwe7DSBCh8tfjUdH8p5
diIt4iwQ4+2Krs40HzdMZtekmF3/oEmwYqd9v/BtwqvNQoZFbsrs2/kITEKc
Ml1EJ/jBTJEBRsSWF0D5T80EbLDb/AgBHkwXb0qJOn4tYr2YsmpzTgP/QxhX
2gZIsHXQ/RoiCpAwDR1JRhfvHvqnSz6Bgo/2XQxQerkHOx3yF68BM77AX56S
Z5sTeoZK3keFtMDYKmEVJJIX7vqz1dkTMiuqxkKJqAwFuR3ZWEfsbxljeYS0
uFJQ87DEXzqKBuYcg8wpnZy4dJcfZ3E5VKymW19EFzSPsGlGIGdXL4Ms75rs
QgOWpcL7evB9ZMPrXudcpLK8FBbwxyt+AOGPKRG/DcTTD7C44jKEpO1RvFfO
wls8ji6uRdVo+n6OeQYCl38VFvyk25cj13Iy2VcwVhowyhpti1oI6GEtUeFL
ODZNQx0j6I3BYWMz6TwrmKW31JX6aG2AxAoJh45oOgHwUmvgzpcztCifwNJk
jjXnBOrRX+E1x+Fjr9NMx3EH97m1O457HseYDChGbW1egDvx47XdavraWlft
/mkW1thfPpq5qnHSUOar9vKyenUC1x31ENBJbpoYBLgTaKl7l8m5vJl9vNll
detHL1bpnjtmzybCk6BTQJz5brwrP8UwIWDtefGFvh4Ce6Dq2xaKLNUV96e1
98UHaG3rXfSMe+UCbAWTQ7uY/DUZQ9SiX4760ITHEMLEVUB9u12StOCbpD8m
aRHyA7OKfeDuc/goPY2uwurzasym7aVX074cEbfLDG6S2OMQuNPzHGs6ZOKn
owM9nBqDxTEnTu71XPKswWVIxTqWZD+dgeGviYudsJUTUkVeEilDOHKGTCST
AXctuKt7to2KDJs8/qOuEzjFUf3+gouIXet6aC+bj7oIhzL5u01zM2nEvvRY
NQ76izBIim4b3M/YR8p2Vj7heOFH3c6qV/BTlYePTRhORwMEn1ubBH46mbQY
d8o9IrFvtkF3MFSGIhA5SbIwvFPdYP1H6wXUU1tnbZRJbdIOD8/WQFgNKH7C
k4XKVKRR0eQZdRzsupHljSpVYFkPgQBWYarxbqz/VNCBbRreipb0SUSC3oKe
ZyAWBsZg1T+pX4uQHp5lGHq94kxL5lKuvZRMltS2UEIPn3f6IrYSkvFm4LGq
K/HPgdH5CM/ZZs/i1+H9xTNrqowGzwToSJB/kZu9m2QC6iot1ZrZIMhlEOr6
2tlK+R2b3nV6BHWfFhzQOEg6krWpdIu83IpsL53038LhVOQ5WonE+Xf8z+ts
95JrnE4I4Vz7iYRoQGxwQ5na2CsUMUGppkCDccU44351SCT7OIoFi73A/QIj
MEUPN3S3ot1B9JVPZQF5OwSGmxascx70a+Ivw9hCdPwg623cH/QvabFYLdeO
hgHcBYGLiedWAtvZ7yN8lgvBYugTQ69YIzW4b6Pj6w1zmWYv4t5weaClpsWT
gN2sWXfTEz794W/jGrseWCGrR8MG6NnaLVbpThj8PJNW7KxLnrbq0WpQLSkl
QZFt8acIg6hYq6Q4cOXx8gQEJ17fO/HO4OPFZA1jC9fjEx8jqb+6y1nINHOx
GMTQzzyytm75Wv2mnerokhHe14GAZ/FmPwQt9AhfEySrM7dnMVsl5tAgSemD
czHCQW6NBWMhU5Sth4ThoVQUWtQ+iOF9Wc22bjrqzNM2A0adnvAR+sCvQuZc
86TGPLwGUOdS82HDgHpWqUZGfU8BbxlvPZv6DmHnMbHNGa/jM44XwTsczey4
6yr3OcACZ/eyR/dvFY6CYCA4NIU4dBsS2MZt7/CpTFB4oM2WpATfbJTVVg3E
0SryVjuwzfT1fGI4ta7Fig02UboTFRGf6jlX/MZL+bTIYw1EAnxeVVZ3Ol9n
LSx6/MHwxUaX70ITB5UUT0JpAnzlYgJG4eJ0qytXxdM+oMWrEbqmTeNEXTkO
BVB9ryHKxun4gNMYQSUCTe8pKAKvN2SapnNYgrO9t936Ah1bpICvHaEdLB5d
KUgwNW55uOallZUlbDrlk9IFFQ1A+9Hcy8VbJNL+StyEUiq/PzOAb/f3bg1k
5QPXGAL+7ifFS4RwEX2sErUdwzH5XUbKkIFcLLLSx3SYKyqnyqua+JPuV4r3
tKtuTjIl2hwoDYbKCI4SmarxdAKlFS5jUNoTllQ6O5c51igrd7ZlSKxYLKP9
pl9Y9MXH3ssz7Dl54wEgoPSOrMgcC9Hx21OVIJUcytsXEEapf1pZNiv3LVMl
X1My5vwBCfmToE0zJ6btLrFu6Bz+ZHTyijhnqYitCyvDfWPy4fT+bF29WfST
TW3wzaI5W2ALTfTU9kZO291T1TLWijsSEY6CjrEq/+mIce6wspbruWauTg0q
oAudYkN0Emf7KL4mZJuVoT8bY4XQ+TSXWOe+dFKbK+KTy2HFuILepT7fUPzo
FCManBLINu2+qhFtqNN1njnFF3N2BLRyKIhBgzcVptArreSIANiHxChXh3b1
oUu6TenfqPDsK7LurygIKpwwdJrVioDJYUTiZwstHa4MH3aSu78kJWS1g2JQ
GoOBlvfkqF9c2NKpqc2m5mcbv4gmDCQXwVkEbRfSISrRUHAp/1KsAw3Xpuu0
/ynXwyPle+GZ4vlc8i8ynQ7SSfypLwfFvvuYDMeg6qLq9wc5eeQYqqFHLIXV
ybjNkjAoAyHOMY++IVd+vMg9z7g1BZoicq2gCU58ekwaiQVN4F2k3P/wy6+9
XgnUWkTXnHFLtCQh6H+h/rflBmRA4mwJt3HxyyrMcK1a3192244cMLtevP/N
LiQrDNge4Vf9K6rleuOk+5uagtm5xT58dOcsnFbz6bOah8tCO8VDR5AZsmQY
OLSh8vJskZM2dvpA1GY2TUSQ/3c6Jb04v7xA0zh3hTs7F0EP1t5DYhOnjWRN
QMQzf6f1rC6PeieYEqSVju7Btl3nBwk637HsCmjk8Dc1+0ZoZWLCAeiKXra1
W+9kD67yGda1d+5aSmGLY6pX/sRkTbiCv0TE5vuta8xasgm18S3sTnXXhKab
SsFHXkODPgwbIJymteiTYfR8uEDL6QapTElc3d/+ciPW2n9N7cSSj7qlKCw4
MqQHMLOnVEL0rPyt7mMvXmYgyrYYG7EM8LTidb743LZztuVKWCTf3dWYOD01
s7dVIIzuLliK+UgeQQ9VeH6g/czQV8EhENUMdODFxJAkwCpaLLpQuv+2i9m0
MqflC84OFrslTyb4DsGzVCk39PSzBP/pe7coDQnvh97p/K+NV73aiuJmqNj3
FEVZ5OglIABF/jL90JBwxXyqsl6OVKaHmpjiAkvPcv2zLOArXRGtVUoGwKV0
a+Mui4Vv6676BFM+l7A7Rp5BlJyzBXHuMWaIJJFqz/CiRWQtDFmaOqz/QLpn
TJbfQ81jnHpeJD3tFPSunZuOdXTJhI4TwOwEzoLywkS6ZJlp8jBRwNEGkP0V
Yw9MWylEw/1YXXlOjTeFNkiDRzWA4ZSBbBnMn31QfCCI/0V1M9uDxQdLpojV
rj6wINd25D6zlEi9lOSv5YekpSXlRY9qeWrx/MfT5q6rvz3e+5XLKNn0Tm8b
T+pT63S1DB91zHMo35bZD9o/DqjuKwqBSuFNJrNF44xIJ/3ZrV+D1aCrNppd
6jtsWOwizqzJh83D18kZzsNN/u2iqueqnpjBNLVdvmf79s5sS2Ykk1U6fDAF
fh52NA88y5PYqLkIDQon95QJTrpAdweLSZFQIaVMxjv2soMs8CWdSt9Meo6n
SQ+/7rY/An4GN4FrGlhpWnFMBEHuPdOhZ9K86FY2SmSRXE1kurk47cmj+HDQ
3MjxuEQqnB8SY1WFUBPRZFzZi0A+KNuYH2ZSXLXtX7MXugM1pw1ceWFM4kv8
LLGDHTKgXriMEVIjmxC5V5vRUas3g9UFOl1NL0bA9722F1G4IW+ubsej4hx1
kTdb5kYQxixWBgZzQL0yUtpvlE6l3l7vNk9Pc+F/ZYP4ugr1pCcyrJIkeuO5
rnWghZEZGr83dNqdcCCqFsUEmzPcSQVX9GH+wH4FkiZA9z8O5bgMxhHYgH9g
Sbwp55j3IlJs005yAiU3VJlfdylO1EGcwy3pD4mbSsM80rXC+2BeKg0AkuU4
TGTFYaAUnDRiXQKAaE391M8cfa2D+w3ARYJn/u7F6nj7YvFWTqHd0wpi4WYz
qo+Oy5dlATe8aabip3GvjbAEx6UPlNDn9dweD5abdjhlmwQJ0JdGkAgX2U2R
8Dq5WlxuaFgnkH1XGr0+h+9AxYZtBqisJhfia5HVdKhtTZVuijG1qa7gk9fe
bxdhIfAmfJQI3VI1q0wwxY/lEIgfn/cNH7Ky/k5aqEVVIv7UkUG9nX5BnGpT
aipjLae7iZg5WckwG//DpqvCZpONaws8yVGkjPC3aHCIeZVYtFUCK1yhDTyW
64wCWC1POEEYzxUChDYPrEVJJt2IgC+bEXZXz/Y+U1U8+cZdOZpfsC80Tzo3
LEFA8AepSOYdgssOQnpssOgMRXjocr+drbvuQjJPlRax13T01VJ5RUmV78/A
KzgBEVRkIS9btKpT+UXxy3HB2OkErnzQ+/1qUo4768fVzpVuI7V2KMFvQf/g
vzpSLOZBEySFO69zsO+oFX3P4UmrqWPWOJ1WzyDgtsZhTxzaNvbpeHPFn81w
gFjf3peyAdNdjFCpILu01J52wN+0yb2w3WOR03rRi6J1q/tIB95QXAKgu942
ksBz0yYNGpyiZr+08mG1SIAG3x097kSXClx4vxgD8Ey/y0Cwz3au3RfniYZc
mQVxR2P3Y8gfhlKS/NYwQ7HSaqzUZTWl3IIbMAfIcc04H6UwUGrH9wB930yN
niCrsWQK2CBsC74wfTgbrntCPw3uQ5qqJ6spSbFiZ1FuQKKQGZHDeUU6/NVz
qrNYM9Sj2ACsaG/YSDuCwcOYtuTZU3Tjx+YeZx2gH1QQs4fpWvqgfjactWef
qma6sp61r4IVevLlEqztuTEmPrKrMD/nqRZRdORZGnrEHs6M7XwiPnf9x88f
z4jlnIiQyJSYaEf1Qw8BowilvjbL5TZGvKVi+34TENLiJvcZ0+QdpUcZDh8E
rzCgGNTuV9/JUCBDxu/d/319WifdVgicGbemI1b+W/uZHKINPN2RwBZeaWYI
SxRYlPaQBKxJmbcRn0zV3xJtLK6YvgVnnXeH22Rh8Y0qHpLObXZNGwX6Yfoa
cUQxqN80AwpKiIksJWeKg6869yESIMwdX/DIquIppBRAc+dUFzgAmpHo2NWK
WUA7Z3mqLVYINeXBu6OEODzVct84yQXg8KXy41iD1q2pHdyMH5zQvMiVKOjs
NghPjdOHjkidTjsklQBybI1g/SzXSK7+PWdbA93YS/06Y2ZznR3jnsfRIeR5
uAX+RF+/NaTFeZV7tSduVkXlUVmsEcLolMD2rQFw4OD6Fdrr/iN/RguTCoZ/
2j94Anqth1ju1r0zNFTXhuz3NbG6dCXI7FokMQFlHAok00e5RfhuyHWu68ko
CZWxPzROj8xnurJJlfzJLE26KoS8D7LSx7cn8JTlmLNdyJ0W7laWd953UCTa
5Gh1LiN3dPuE0WMjAA9gjGObnq43NjH6SOOVizmS7i+uosJZjDiw8J4sniQ1
rRutPDDDIwziqnjUrzbiPe8Smt8Fi7xqfmUqGFZypKS9dTB2omjporg1U5r6
w23uxRkl2TrRTPx6mme3vhq5Qx31CBjvg89OF/X4pHYjqavP8WHGOcJ1PFWD
Q2RF2N9rTH2411DAA/IFrs3AMQl2+HLeSQ8jxIpAGcwMrtnxvJRKDXP5IA9L
WgG94aVwb/ZJ/VFNfZ4trvZN4AZ/IvcNBFmnEamiXUyON/6Ag7yfGOu7RwiP
+r7LoiDSKQe3eZZwLSa0gdcMSyGD+oCPoeTlKjmbTT2kt8Kaj9zcXfqPM4sl
d5BSXb3rvlaSKK4aW1/+9XPhhDUDx/cJ+rG45h6MKxVp5aiLMYg5cr+n62RE
uAFgS+SCtVkhKL8g/akjP2wjL4NA7IAII/W0vOrLoCcdpUnAvqnKrICzLegw
VxcUB4/x2Tw8ZaJCGVKjXUHZ8Qxi5dhoNR84macYBhAmdUjJmKIkx/zv9vou
aPteHkMfmF3l9Pi9kPh/w0mTTb3uQq2BSmWGaFaMoFdsfIi1GHLqG/1sh2iE
bbPEAJ51FnxRLPffJjBjXr/Dx2GMigoqphmZD9PdFbolHJAAr1IiyIY96uJC
FLZyZo/0yA9cJ0GyGk93atlyK+JPiJTdxmdcC1QIyjpSDI+1ZmHMdn2dybfY
t+QVq8ACH0qDx4cqsA68ZS+UtJBFKF82cD82SOZuNleohgBMZi97uABcmfo1
CJAKVWN8Jj18m2u5h7fqRgeoqwtCqXpxmakNMyBaEOjjaUVDvRtwa4ksFjXa
js/mk//lEBo2dUu5dC95uRiZgSL+RRPX/f+vkXS2evL90Y05Rw9kg3dguMi2
jvb8eBCuORLs2GxIo99yAF++Hjb1hWYE8x83oTU5m6KEDk8tSOU2RCtU68oI
ZiKYMP2XbBNDs1f9yHsoxi3nQFblYJulGC9S2XteF3Gtqeue4Ta2dBVZWz0Z
0W6l9YniyFULiFYuly/D265Q2BkrgHD8A1TipiYtBPyCSYT2TsU6v4N2QLrp
0S7eiAz+Ob6FMGXYrpqy032tHH4BUwzMtNksjIe0xP8uZbufLqJCzrmTRL1H
vR/CmIPM5wEqnEBaIp6JUxVxSu0rEPq9fs9Zuk6nOjTv9+utzdBnW1jBFVJH
UHToLwKw+Q7WcqJrWpd70H1t8/+TVHCSX8KvdhOPPgMHoSzBQeZQIo+UQDAa
jah9XorEW2EQnQUSOJIZz3sU1uVxQ3WcyxPZs8j4PVpwqTdwbDwSIS7vHvd4
JU3ut+3mkSnlGE1tZSf37B/pyj7Hs+fvd1I7pZXvLi3vdAYuMOdQfUe8SGkv
2uBwngDJEcKOESwYvNsGIzvp+Ovi4ABED4Df3rdmwtKxVxtPklUcMsz6ms5c
QVrbyaerpQK1et1vjtRyl+rdg0LwCM2D9qh/n+sbiv2QEeOULSr9ZCxnXh2s
uhYWoPiiitRNE3D6Bv4rfR4bX2j8tOnPqrET6O3KPfOlAmW+mpQ2Wz3DxOpZ
q4Ug9o0YvgJsCMF2WvT9zoSXoLma5YWhDrWXKk1C4gEnyfjv9Evqk0UaoGfn
8zSntJnVXY2PD+iku9WZGUQ1ExCorsUc3SBFBuu6UFtGk5cJgX6iO71sjHNS
Te+3+t0rPRlZYcNSu1YCW58kMmwdpVQ/+PqJaspfWr/8tod+1A+GdIOZvHVk
8Mzb0kFappvo0cv7YfwYQZfVEjJFynrVZjfTzvic0/D4ULgQN6E3e8ppgWQ5
Baq+DYM7DhY0FVwlxW5C8H8nlM44c699G5PheTYOoZd6WFyqHMo+M67W4oqS
uUC6ckKBygXPURvpgm+NpGberac1zSs5PGgMsxczAWgHYCcS2kLeynIux/yN
5FX2UvSEr1LyI062eUnJVtRoaoHyAoAA+di7afFHQSXUadxvDu4m3lKB9DG0
+M4kEW6bKLSrkPS4dNgyxQ6xu3f/CzTWsb9hj6gyB9TGxC2FWx3iaNNMdGWu
05DvJW9YZM/0pUKgzccw83WxuJMKjvTeDSTuUB4c9k1003kwGzh31ODad0dp
hVsspkLeApPGRS5WG/8YASp1wth2g7K9NvxI1ebgYsdT5mj13pYL5EVA6jvA
Jc7XP4AX+HHFWSmG4Z9RssiovSK+ALts9lIec6vxNH20a5N/LbLEZNXNqeg/
yqHJlM86mg3RQZfYi94tRrPFspcSmx5CIxqogsSfbS/ujQzhjrZ3mcNZYdVl
wQ6skJ9rTouTKeaGPRouZqOXLYk71j9Zi0pA6qhd5u26OQLuI/Z+BV+iO8tD
bI0dvNGwwVMme6/TLZk4H0pjJ39RJCtdo6Ab/TqJVG/KlSvLlOdMFsFIO9bP
BzcJMiT0WR9OKRYPl72f1xbZaZDo2qtERZpBCPauWmfhl7RI/A4F3oyDWHS0
Qc+HjlE8V+BJq36vftkkg9cxex6uNGHRxfcBWruOK4If+MLSwa/WnpUp+PNj
JZjyL0V6fzmo8xIvAg9WiziXi5gw9vEIQw/EnFhaPzoH8q3UpbEWcAhQCMDZ
4K3IL9AuVWSFYDeJfNuDQ/I68o6s2bm3asJY3dWG4hAFDpDSDTUHXPuKbYXh
tjj2/NzkIqSM+ydaR2odxk+5cgaqRw/PEphATM7B4qclzSc0Ih40ZD6pLPye
vic91L9jT6F/KOKcaxVZISIsv+LtUmtTHpZmAqMBOZpSAEi8V1vgElk+UTLo
+fjwyEuhkDXzG1cR2bFuPnddJgkXYOkJU/7574tQRWs5zrgkRFPMuM03pxxU
fyaHHIFzpy2ZrRDyr+29vadXudgXRgYrEUbivfLA7XWn9gA+3dIdppcYsCQI
6pdt5DDUZLXh7rd2u8HWzWv1Xgd72qxrHZWY5d+Lhf7ZyAcIOkpqcc4v8KqH
JoGIr525yKrdKVq0MWgBJyxByk5PCwEZ92cO+wAtXgKAiewdvEuoxfUj3WYC
kSCmXV2+yQzxFa0Ps0F0aS8zf0+sEaOYErFZhbUO6ZCvNIDhXF70z/qwNb1I
WuqdQBF9mWVyWKXHg+FLCcs3m+yO/i1gqNZgX0IReGuD3ckqLy8OwM2kVtbA
6GChAwo63j6ewurmwyY5Y8zb1yCdZXqSBvJ0DLzBvDuaMb8mUBhRpDZZ2nqn
7JrqapO0WE++IwufCnk0oABPCqkkKVq2Zko31dZ1Mm9mW1BiBMJvYWkSa8yi
C6t/OGcn5Ka2A8S+ARlSMMyT+gNMvsrcc7mUMMw/pgOk2giz2ojp6Q66v0sg
XBbmcKV8GCgnEOnBV0VLRyB4iGfOJIxKpX3sBPBkI6eBZeN4LTWHCesR4wrz
I7ufhgBq8iH4IxOQCtSTv8yzPQbNBz6jrdDpIkvsLn6sOBIL3wfKw+RKeIiu
A2/pCM4Jx+CfcOlq+2wmiy/xTEkXYz4e4v3E45XmXJnTiH6I1cB43uReeSK0
TcU+sJe3inO6nDRSctJQeTeC/lwZkLZRQLajxcg84ueFi1Tuz4Hkc+GPPD5t
wbbIVLlljwlNVp21UnrD5WesI5NTb5Zf/FCPJmC26WZ52y2NeSo+vrhsfEzb
ntKLnfHVZhvTY+Swl7rEEw4A2zEd9PBmHIS76T7alEdInQTQPBnptEe0cid9
ss6/c/jK14NN/KiLUuhXlRrqxOqBpX2zn8DgUDHRtT9VgjDO9hMkWzUi9Qnn
hcR9xHoIvi3mC2I45DZi3NTzbOJbuEIunN48UNhO2EgjjLbsZqTZVRReqT02
1MZUzukkSv4s1aDc0a2zkQ0Js/VW28d0BushVqpl2NkXXbs9ubp+eHWEV01Y
9YB2TGvyf3xK2TtlOQJvx9Ft2YvqBKU0yC5bSXk6v9c8GhPa17zevVbfGUea
foveuey0Qb7B7tR29qADocAa4TG5cMuC2d8BM0PqgofmG7cWrZjFPyKioJBY
7n33caJ7EMghP2aPhtPckql2uJf+aFTD/HyU1d8OuLa4hA9atxjl63t9AJSg
G0M3zTxBG9FDrF5rE50V/so64eq+btRgHhlmGhHLU5hLxRPeFr3mLpItj2Mg
hNd4iM4+Dziur5PALKwdOXYzOtte9RXcvHx8RRuk1a7eI2YrItZOCUzowjMA
kTbfHcy+AHpTZCwMssmM9Gf1Y2gNlKe433iPUSlm5PF/GUNY7bLWKnOQQ4MX
Z8u+No7pIayqvSLDDnrK2xQoddgYJfsaAmhAioXoCLiidAw5vvb2lzi+JMZD
epCwHAeP0JEXPn+7OpyXEoFbpNv5cI8g71lLIK+cvpz6VsoA6GRJchNxqRPa
JnFWqwi24Q6YBQ6C2lYfQhBAZ5hnogJzVN16m7YQ4dQpxx4t0hV1nEFpmUk0
SjBpDT99Uc0NY//FCHUrFIFDNmpMFbJNY6naUGTFsakI8ouqFKZc6MHDZONB
DkdPHQG1IHH4qnhUyPyruDS6iAyoTzNCGdS9+fhH4BYZzEhcN8LKU087sCbP
t/1bvrcqpEmNbAyqF7qB84QPoeaRcCmY1oVVqRiobR8lxmtD5Id+8ahbGl6B
K2dl8HMqBPmDSfDWRW/tJiCAHUsuDykHZa3/sle0NeQJrgS77enykk7MIYJr
4OPaDAuPgQ9FGciC7McLl2+EOOZGtmll3rCaMjef2rOlxsrVIYpWVCCCGnug
V6BgVWRQJzULG6Kdk4k4/fUDmacOl47APTJtM3cff66O7ekbepgsUemFMksf
EnIlB7oGzTJnBn5w/CU6BVt3EsTf4AOTduC5ELI8PVjj7ZEXf+Jkij+e/CsO
uXywwB23F2P7Xg2NTH+iaT411LRLQq4Wkw4IuiSCQrL3FV446weKg+isChr2
Sn3onA7sgFZBDl7k71c9lfs0HccH0E6e5DhyWWckfPL6r9It8BKQoj3KeX+t
5sYydEPVd53vRFPru5TbcpvAj7K8xl2hnfOo1ar1xK/3VraV0W91Gx7g7bqw
4YDeKue6mPgsYaEAe1ZE++vvTd5WNv/p6y+5yomYgpRw2g7vYZHmkWhZvdOQ
FCD6lnGL33wtt21Da0L+OMmWUvHprMfZOGAk8GX97fkiZtUeES/vYQZRiwoo
X8Wkv22PK4wuCC9j/ATB7TQYqHTasDMUMuEvLiSxClDZXuylnhU9taSa7bVu
LSgh6/8ZbcNVWRqC5AQZ86noNULhGAXh+3Wpo839smJ7q/suQqidrmUAfhBV
z1j0udEQkfuVpV5L69/DX/ZjsXmp5uTGTrz0OIrZf6HDS4QOih1PXps3fmX8
9DgZG7m3xGvsHFZhJSxLhGr94r037vKAWVhKG+0FWFB5iyYqNCPcfCdL1C5u
oqeWWz+agNqbUavfD1IRLd1t24DJwI5anEfsgrn9J+U4dN+ELhDXKoNHq+m2
5lWXO2qHpGW5pnQVZbZzlnDmg3+3qvQJwS3Nt4T2XjOOvccB13hCK38lSiKN
tKUWEjjchQzQ3wnVkLvjeSx663W9s5bj3MROpCZCOJsut0Kw6JjworXNnQZq
4qwGqdyRfQbMGY7HfrEAo1VEpc5Ik6hzAurPiraNMY/sw8AfCOyWS/6Pk1MO
9r1s56igrXo0cfR9XHQD9Lko7F5kBAwyHllCdFDebl6k+kGnDx3TUdCe7njE
dX4DdW35NokjobLm7gual/UePAaF/0nogViC3m02j0kOCXQAIUUj8og4AEY/
BMaSqjgcnIINCwu6efSMWH6bMH87ruJ2KZq5UK8kIHw1E7TGUlmqSx31RFc/
UY/OSGldfusvyLsPRi1Q8nm6C6DOi5On/hb21gpbmPEXqaoBhX2VKFMLOdgZ
p3MXzcKzVizfd0OKW2/zWSx/1kn0G/q2+cwQjA2RmhHCUZRGWkcRFjY6Pv5I
OH3gQI+N4V2Khv7RUTFKEbefdtd4UwiqyFMEs7X+2/KHhYdDtfMZuLOCXbS7
FUdgsAY559I3Qn1sdJgtaxrHqYDbo8mqutpouIYmB1cjiMxPbq3/er5yPpBP
ld/IENFRXZhKu39btGRjsnEAO5p/GqZ68BqVFucrXRpISyyhWLDlvF6nKekH
NmnWC0DqEv+BfhdrAko5+Bu4L8AsZUmr5fnT7vppt5qV8ga1gRhi1Z0MuWyO
P5qFhgb8SLJ2XzPoZtRd5fB5U6YrhVuSxHxhTQBsCN6y/Zgg3jhfF71/R8Nu
IDBfxC2gyiSyumlrSX2DXDJ7FPuisBw/Geku0M/j5ZmDJW3ZqYTYE6u79IOO
ksOtGaAI/b4UmCWo+63Yewm7jBN27WF2G87nHPVh4uv61IJ7SKszDq2lqIg8
6sS5/tMYUi6fK7a006Her2SQEEm5odnxUsLBwecQagB8vxi1j7i1WfnpBeTp
LLdaKNAeppAgP3KMwy9iI5GM81X9CtmARObGCyENclBlvmVTgoeoUEMDCDwr
u4Dd9zH4WE/VcxRvVSJxMcs4HMqP84JYh8zxnt86EmH3BMycP5awS+E2bYpG
984tzyTTWBdZEkfdH/Z5TN3M6Y/PbgDTtoo0q94x7j16JvFwOQkhvACdf3Ra
fp9/99lr/4nVPjt7Didzc88abxcJwXlC+l8WWBHWnVA8f4ZmSYnZupbw34Bb
Si3g7HPN+fn/4qh7W/hxq90Bs+hHbd/+RCpAq7vLiBlbJUm6ktVWCCh7c/ZR
XkPZ+5+/iQEfdz1o+YSs3VMSnsij4ue9oy//iXxuVUPUIOa421wXJlJ5bXHL
qxEiAb5Cw5rG9U2nOA9aKGY5nYy/0RTXNAK2StUfKg+7Bb9MsckAhr+b7mG4
Y3MCnA5t9wHtFJvi8lOrgG4P7PODy0JJVhh77LjQQvk9lwD/3czkIhwrSYIp
TxUUUrC+259rtJoKGG24fLOrAgyw8NkvkpmwVEsj7+Vg6Ia8wjm+bl1CA06m
cwbdMnZ4M6dTE4rCKDXcrEqCSE2/DK91fPfB00j2TBiarrcf2V6eQZNqXMQn
iVIh2H3DWsLAfusqPxH0a5A0iGhZHpycYyHfJl/iSxDoo4capYDMCvOdULnJ
RYf1GDkKv7hCkz+fV41Bxeyipre2hwo/L8QEQnDgPyCRBtZb1JcN5j5ww3VL
BY6Ri21x1TxT3wjzmXlmsq9FKFK8wHkj5a8uor0K7YQuXkn1PfvgYt3LDd5P
TVbccEGyo8joDuan8J6dbGJFPstG3uTVvYtcze6JMEaarouKbRUnRRCm/tn3
BkeT83LEsxdIUx8qALkmcBIc1Jw+GhKfFsXk582CjdO0OfwGIvPxIOQVVTPR
MKX/HYrfQhclCTnuejLCYQ2SabrUGieKyRLAY8sSzVbuU8/946aj4roQceER
z2YI2CYcED/0hwwyYRCO1y7LZLDNmacza1cTTR+d4yIpO/0uO0MDD7ThJBfp
K+5jEkiUaTiKWFSdi9Bgk/rdxBUWCVwVoU3Le6MRguRjDWUdbJfGkNu4bfXF
CYIi4RFaC+xv5jrRZ5RdrZECNSoAQiXEXDjC6cfitwAFNvFm7IC16vykhFg/
RLCYDpHj2aegceom9FMWDoo+YNrIIVOsNOzwH2KxNmDY4kQlfb7LCa0mvFAZ
KsId259kshZLEh+mz4P+RdoLmXYx/49gJ4TsHTPE5eZQwnigWU6QfuwpqUKi
h5+hH5CABS6MacpMh+Oj0JcjFjONJODZU3Rx2YRPdBj386umVP91PjlgoTBT
jKA1Gypy1WtcmTMa4wQSEDW8BNDlBsHsSzlcsCuSAtA51RHz7DiM0sPA1ELi
gIqVHScDlbIcaVQ6KWeothrUqpYLBJHSgfvGyl1IsmxObQogOgg3la78+Ks4
uKFWQxQBj1Q4QshlrU/WAwEMzDJS/oroYvTaUlhU47yPAkIi2ablAIoDQ6UJ
yrTQVu8MKvhryhxr1D2rQCdE5qQ7nBtymaRVTl6hU4ePYsiwiOItjh/nnlRO
5/eUwGuu3kcpzBQVzxFbqAd8bA3cSgS53Z0WKdV63iRNH9PInPkg52idIYRT
O8tmLSVuwjwlBpywr2SMG/r/JePSxaO+fcKB01VpqRJhHq7NkZDYSFOHwqX1
BJ7Bm6kQ9FdWdQej4EPKdtQRJtznOmpmBu1MDJEtG4jwxJNAvsgP1tVjR5Uh
LZ5xdfBSRCH7o77X7ecbrcLfLCP3EAZiwfwdC/KGkJVQqquYRiAnpFsi/AUH
5afLTiHGmnRf7r7KYEK4W3wcgixPOMN25HPj/xnDMrDGHytup3tOGKmkEbdw
a6cKXXQQM6n1uSKCaEJ+xAZQXRo2hPAu1EqaK2YRgrJlmFnw0dZ2OY9G8FyC
IkNl4gon9xfCKiNIvqX/2PZOKIkx7nqIkkBMN24KVU5biHoXhQ9YV0VQMrH6
ptLw4cMh2lXLwUpXWj4Ws7ta0B75datLR2EysYIsOVoVcqQhmek2gMPrgIrr
SjRbdebtB4+p7aAMpHXJrecBMSEN1dipHboaVlIZ+1iq7iOozfVfXWBpYm0R
S34az88jUxeskhjXVxIF/+A3dTC7eev8PW2saj6xTRjJViQz61lyap6hw/9H
ZEVwrOAz2Z3DoP47U62x5V6wd1ZCnLHMEOw00rL/mRuOADfIP/6+Nzrpl4Tp
p9KniI6idsF1CpGxo52iKuVkSMcCAPqx8K9zzn0v6VbJrwLcWPhsJgGPU10f
eBfK/KwDNtODo70Y+LwAv5M/gSUg6xQmZAjXLTqMj2e8XNDQJXXbXJq5DXaK
WOS3GVYwUKRtLR34RPoOn5Or32+MCtxE+OS2i/Yb+HEjIfV7qO08n73rtwjg
Rvm0n2I0IAU5OlS+9xiHi7sFEQXIGt0TPphELZDw/qWSgECXUtj84BCY4XHe
KTkE082wLwXKUzNGbkNmCuYUMPLu42pK5Z+PqQa+ipAxdEJ8KG+1gfcKwsJA
RD5THWhTHVeKgHI7HwZGJiWfRhPkDGHqf7xUYa53d8dFKuMaXO2L5qC3MdVH
sY7FMXbWT+T9PUduEh0qEWVpM1X/FyyMdJtr8tYWP75LdhjWG4A6dfyJ4e6j
ifhL+t8GWzWVxCFMaaaH4I4UYcxxodvk6QIISDCwXzCIlVUU5lrm6A4RMD8n
Vus/KxKZNhgRdaf8kPsaFxsUec30wkoteCVPYBgV/samHNxoB8FJORuWmpZK
pQ13M/eHxnvBzAh5RGBtVirGGSImWlw/4oZuqkH8Q8p9fc5bGfay5t1d/lBX
ySU5NxI8IvFhcxv0Vu7mSK4dyEiv8+kiz6M8zCiRtSv4JV1J2VuTiGh5ZV+H
7lJlqSdkx75IEK7aYr0sU1OORyVeN/AkQCwgk2utmZZjNMf30cdu+SqPBq+i
DEkmz90NSLdEUMn+ZtA+NLRgWShhUN+y351uIl+aawUm/qGwjbXYoWBSpTVQ
qUc7Ob5SrxoR24A/45yfb5n2fBGrgNwJjdZsw4G/gho2l/79QtpsnCbaLzh3
GN+gjGjQJTXDBzvpPZWrzVcYbZchtE8FLI5WYNqocYYYkRmLr/eAdNkKKsDz
DMf/gRkUvFKke1kUiSlFlqJiHAomcAQYc0W4R7r7H4lCKPhFOIdLlLFBPgUK
x0UeRkMoP5vTu4Z9xcGP5XwClhgheRKitSSl8mwk7AQDWNdAQ75N0gzjopeP
6zajTOeYETf+D2oPQV9vHGaQbf1MM4oEMtgA9VzCo0S+V6EXE+YE+zVOYfgN
/aOouiEdxTOT4TIqD1vjhxSa7Jxd/50ZkwAlmmUgndRz21FT+QnLR0SKyIDZ
ZzoOfNwYh7FnEiyH8yVMCcIvgwHvE4InysuM3Ba8V/Af/fBdaOt0lyuamcac
5eERFMLUolWv1nNTGMKebT8LXfi4S0eCpSkztMgXyJNu0dCG5cBA0Olf06ws
SUQ2imD5Reez27YH6nKxPDnzoAGo/s6Eh7gpntbGT0eHlfN8iJiE9O2Yz3cW
w/X6ci6V/xKhwCzuJ4Bc+oRBkVAUl5GAk0yOx9KEPJX7C/LJ23F4Asr1Fdsz
L0lu3+pDEB5QwZ1rb2Uyv6XcXT11c7eF46zO4/xYf48Z+umk5iXn+KXTiTDT
6JSV6iyA61WD/PrKtsEfhn2cHbkEA8gqypDS+AcRDPmDHz25aY6dXFVnTk+5
8E0zUp7+dE9qF41/p7ayy/SFrl/D/K+TEu8GRhCHPyWhkj5vniwNZOXkKnPS
+NX7TBpCHTKWVSb9Rly0vdWHaU6b4hM2KklwAfgsygijDDOess/ZJGJOOWgQ
aoOoVztBpy1nk9JYHpqczlRBaJlRJCX4rmRT4A8S92g1Tt9dz5T5/m5GfrdH
MlZH2D5xyksKGIVdWpAZyWjAHvTXJBQTnw6WAihQuAPEHW012dyAxBHP6h32
/Kti1+HlX4Q7pib/99nu8gA/LLu7wvLFez5KWiNXvQMa9DotgAr19bpdN/kZ
X0VXKYcWSWAduZLpDFdOS2+kjyEk85Oljp3mYnbGkL7bWL/hv6fv9fRxVvD8
cO9EEUCXgziXfRaAEIDYw4BeN+/2WM6qIDWBbu2J7stxCfINImnz+gf3Ykif
KzOHevWHhy7QLrOd7lAVD+RnH7oW3LsmnJPd9PTxB9xvpT7E0s5470GriKEk
t5fvrDO1UQkL0IJ4CEWKtCzOs3lscbyIUWCZSC1cmHnssu/E+20LaxPYLeqH
Wpn0Nmr/GOKNvZCWWMJo6hJg2gES+hkyMkABU/OJq67qUruEJo0IMBRXrQhZ
TlmMYEjuoWGQunLgP1bhd5Hxmcp1fpYaKVyHmtSlSZr9SVCrFBZzWOmLMuBr
9QcAobyTF2PpTh7VtmqzIZEaYquB/zAWsSvoH3z0WBPeUBMlPGqti45Z94wZ
Ip1eKnJYrG9AlHE+C+TX4o7gq6rc/nHCQX4/V4++cNJh58czqK2rps9LH6wB
ZSHuUkb72vz5LQCm2/kbS/oy27MIMySmVHIRTLsyK9LniOjEwEMbQ3qNflqT
gWwc0VKC9MikNJEegtFkOG1Mv/Gy2RX5nA0duS6/fVfnTFZ3IAOoLwvh2GLS
TSRcj2ckOeF6Hz+EzYoazpokKZWDiuuF780Yu9y/4ncCBaSWPHKjky/6Sw3v
R6KFBawLmctZa0Nl7JyNTR5iIQdb/OSGV1sIFf30IQCgH3LsibHVRp63CSJg
aVonMVi93hfSY4G4dl8bHaIFaobwoYkN1/AoMXvqckrMw8ijUJYzfufthVnN
S2DlnGscTmjYAZ2ruzrahpzfV7RDqD9NCciqN+EoRtIW5xoveXzjXSTxEezK
5yqQsvTMliGBXuL2pYEGhslwNqGz4xFSkLVof3PKHU3ZTC56EaWk0wmt8xsf
/hd13jP1XEDw7IL8nI1/BTP2Y3tddp5gZrhjFCDfDOGXT/qGQGVWeqQfV8zv
XcyU3mjNFMZpvrPCb5u0ieJEnGunITSN3i1alvgWefsF2w8R4VUVyQhDs0Em
AWbeAZTlwjPy+5uUIHVOVzA6F1ZuFyfSiWGbs3z9kV73KxKm5WbiM+l/ozO2
uQh8iwtvNGCy1B8vAKD4Hj7/7KWi/3nCsGUdD24e7ORCqZtjM6GNG2DHZDfA
QEzJbZcZmLdCqfYqs2W5mqYMzvaMFWcOx4J6RCQ8y+Rfc+PVdLF+Fj97oE0Q
4eKsTxLNEO2hyzJGypeFxH0y4TPniug2fYbT7rjN5J75a/mZuRZlJY13HVWq
c6qS5aYARme5Q3X2fEoM+d7bSkAdAcniMSL+3TJvl/OXtNqU2YiR9/eJYqCR
WlRkSNMypoW7y8MbR916142L6TIwtsXV/EU/VxVsFLbjZPR0NK1+L1/pKwMC
BE+vRf7hDYBdOg0AlTqrlp0bsShXttKeeYMF1ovtaOFZAqMb9UvLXHOaPNL5
8HXB7D/hIwPyHPOo6BK2WK+kPq86cqyX7FTiwIp/neIu2UwJ+TuwQD3+Oj+b
H5Lm3nbixowoZ+Bdj6HCPNoizBBkq8a5P/vTgfvYBSYlT4TBy1YowXR/7m7d
76Q6flSQ9MP7ZonNS5i3EFQcnOGktWJT0JVmI01B7Z5LNbUHo3r+Cj1vywPS
qlAS4eG0fGslMUhNyndlh5bWr0XObApow1NHsRx0KFH1BeXaGUyH4Cdx5uzs
6eKn5QpaWtx2Gh1wiQvggrcxnqL93W//Gzh2ODCHl7MIIGEfAREjfhbsXBET
xxh9s8fuU+plJ57Zxhc2UhY6XJyJaDkKnkh050OizHEoXtDk4WII14SIzJ7s
aEuQDbdd3/BnKNZ5fsbCLMvHMV4+q6egmJBsrdyO++qfhF9qmXa+NNsTH5Ff
D9fLT/0l2ku/vnnz4Hd3LST3WM8Vn5Sz9sXPYy2+iJiP0+QYENyXZmBeBjiR
0bzits24i85qfh9zm6L7doH5tugz+p7j3nq8pndS0Zk/ovwaQRRkI98TiydB
cqDQDRUrpF3pHFzkoaiLhdD4LGOlSYQZxBnkExjfoFme28Latvx81pXvfq2I
Sfta9u7xa/nnTq3+OMKsXM3aDYTpaDErKXKoSPwtTnPNA5jbR+rmxtk36FhZ
RSSREjJiLdmLQ+V4qjNgrGdaMjtBDXxUoyv18l9W0EjyKlT7IjU+YrJQhII9
50/vA2TRrEfR+5n9mDnTIXCkw1jyOCCL7k+BNq+ed3W0QMKHMu/3G0QW1HRR
Nuy4tcF8Jmiyd375Icd9YPHS7RPeTkyXTIPetjsLwObCZHwSTVjlSrNIv/n3
4nP9ja/fY7OsESH77dOv4/OX+VLs83qZlJrgLGlIpXHElToEoa/GUd6+axqA
cG8A6XSSKXGo+GrdUfLdC3fuA8ZgCdFQfcXmTHD93od//2DNsmZdoaHwCbzz
FataDxD9p7og0cT8wxmMseUE8wlgixmDbj9DyLXrcyaRLKOm1b5Zj3EqSN+Q
lxAQYOcbXIlFJQmKtfr/Ih0sy4Gc8AY2jlT6o8G09SKp+Uq+9U+z2SnwjcaG
NJN2NVhAhVux2AyfwMBH+SWcpRa/rQQlWeuwFWLB/T7Necvy18fjFpyxZrkg
ytxLiZ4bKCvggRO1tLOXW1irk1vq8PdMdE7oXXK5GHhlzJKyz2RXgse3G2hs
o8b3F+8lF0RQPDyBh9+UpCESGOEPDfi/D/m1gr2S6rovhwF+Wqv/JAHzxWOa
HXP2du51+wHTTjuoa1c+1orb+4BNc/rj4ArE0LmFRbLC63bgb3hO9osJc5gz
Mrq2zBpTJUhugsE8zDTfVWleaWnSyCOG5D6S6UZ6tmP6RFius3rfzLzq9Bxv
KkKg/MMY004B8njNXvpGvS6kI2gcXspqMisWXFDkCJoAArIi7/TLSfffzSQ8
4SQNJruec2aqhnoj5aomBtwb3NHxlX1W6J6PumkIkRS5YIoKYkaxgyTbFZl4
YWUO9E2sbpIiPxIE8Y1JQXp+Gaibz8TOTV5yoyBPjXrj4+cij4UQFS7IvSOr
2BQR8sd4x8t5Wqtk9ykPlRPiOWa00AZ4DIXAzW4ac+OSezrwjkhtxZm0rZQt
sGZdEk61EKnmVUQO6K76XxulIXG/2s095nF/1HrctOYZ3ynKVgzSP3DNe2QI
Wg7UHZj2qNtZBQu77DV8WPphHPccH2wGyRRRgjifsRxW6uKGts8M1FED00Nx
akFZsLtD4TQq3FmGoRdnIaYiKcEu8p12NB1K+XaapjLw4LkGc/DSkWYrQ91s
YC7BdvyMe1TTCL0F8ZiYi73YpBzEFryC8GtxnRNA/GXloPplQFgqfnr6pYxN
QvRW0MeAtgnBRExQrQYO4OEY7XBrsQeDWgVVbmg0R2okMkbh61pWp4hWSYCZ
LWjVF0Y/ZRStTa42av3LeHgqQdhEOUXkwW7uBNvI0vwhz2IhJjhOa7S2IqYC
QjPnNH+XUQ4JW8dy/VPqY0BJfcVnCf7Cmg5mtZxNlWKgyqlSsPLuQmqkorBN
gNmmwzk0qKqmrhfKSUPH3iDwH2RV+86kuL3GrtYsb/BgETRiGNqauqHYW/ky
TLtr78hWJVtRPWwz32Z9NVipYxmDDZtYLe6aM2P53MCmt9xnRQ51woHVf9TQ
/bC0rK97znMqMSuMSuX6SanK5/R6n8b7iodYDRpKhktIPTtpkTyRThuYEogB
SMdeSMS6xGhB0zFPO9/qvONY5xIVJelXgaNlbDIfyxlljxPu9NclvlRHNuyI
6JQUbkFtl8oHTTmeI1mLWDCWmEcsUxHyOpAb9qmrDSodXFzfzAMvNnvifoUA
5pC97iXCFi0UaDee3POEPOz2LIbmzQAnGJ4Z2v0q5rCFOhVf496vC2Ea5zli
6Im7k1NAyu06VU9El4pcCDmbsbNGgjvXj3DhJIx8EUQZ1+tYXUhxOFYH1Z57
ktJLOVeou2WkF8NPyevZzJ+ilpheeOrvsDE7KsWr/f0JV/JTD1Ss6MdpK+2Y
B4EDfUxF1bCyhvZ1dZyQJC0191htbwKARse72qik4cBW+Nn8O2N9wWqK5EEa
pBRnQT5JuHsvJXxl+aITY+0zWzhDo9BVvWW0XCMsoCQMyZXyAc/JMpA3rWuO
PfKly50YSP2QaTMxfpxu+07jKQSSe0oIJ3h7pK96rCtW18SdzZ0a7J7lJm42
25fsqXGCTRtyNXcu6l3cq4XIDiVJ9Nft7PCJmVin/MxksnOZKxsV1T10Qfs3
E3RpV4boNdv1Fcjj0JvrUXYAtepP63T3kF++IGvQ6+mUSfNV2+pZurTPEkvX
pCU3b6WXISnaP0KN3zGVjVJjXYIxL3psaBWIxGKjr6s/V54BElyXiw0uOa7j
lQ4r4fZMXHKMXjdU3Y2ao5I6lkl1Mh8g81c1VLqUf3hGfUYpb2js88QOp5AK
lEK9VAqQ4miiL9yfsjCg+XXCD+AcWlJD4zBpUTIPvMAfPns20pYaF0nGN/9i
KQ6dQo+wgpDswswig3vzbhv8993VkQAJ4d9jeio2J1IReWQF0Xz9cPd9Op3n
1Tsc8D79ZEHXe9uspQV6MQD/PwItvNzP8kvtx8IKdfHze5b/nLLcVX2GOShq
F+R5BkHLhvUErBwer07/VfqRJ3lVfCn/c5nO3S6bN+IkuxjHAiutqTBm8Eas
ek5tBD2+31ISXCOw5iFxf6MHgPOto2v3h/8TvnduY0TL7OZ45OJpRmpUsv0b
4NJZGcZkw847YfNZt/2SkHrd5ukmYIj0qoPfP+AQVlKISSNhNPw4oswVo5uS
MVzDVqOrD+KnL+vMS2wp1n40/HpO5EQXvAHOAjby+zcFkKR9T6zYohO9oblh
1ukuV2c4or8aFSzqBZOf42sJazLdTaajUXw5wQlAjkAgjIx0jdQ0/UGrEHAO
kaxueCl+xlDqHKNw4PmTlqTS3rrg+UGA1bcfTVOVmwgcK+UT/4OJDy6e/GzZ
gNf9NhFu99Wvg02YidABuqC5z18DNr/5Sx1dk3l51QaPtISOjYcQncOt8SMN
XnaHFMgqyVmFF7avZjW6+AM/GduTXM44qdp7vZeDMUcfcvE4RofOP0XF3CQa
vRptX+y6VmvSRDjpb90kI4y4OLR8T9kBydelOLjXJtVBlNCd36vI4JzcpfdX
bvLDU2fkDw1K3aQGXhMIv8Bb1jwVp/xN2HcVnvwGaJs5HXleQ4KMxcCF4eMz
Xv0VWAWqZ7Eh2yMImQ6aBmoW7rA0zfpizXT85T1v974o27Ecl56m52RZZrR7
ImWErY9ZjGAusWk7yo6W2DIPxm1eKlHagqynlgISjZAV9E1g4S5lP0v0Bjt+
lV9GJY3bwBjPBhoXDSE0uFVz/765McCnzffmiWJaoVnHRNdOga+PJ+rEQnJk
WQzEsaaGb0jnFzpYkvOZe//OAjLNg19crBWBsF9LKs2FxR5ODHK92jHaw/ka
3tI6Xm7b9mS/yVaxXgkow0to8h0me9qtRkVCJP4l5la7H/1KrNr9cC2KM8iZ
2E+CCnL6hsVfFv3DxRfaAsK9AWBctOwSi8+sdo8hhFAfqd5f2yvI4y/W1d30
cSEFOyf+WfwzU4nnzWRHY7yFhGGVKo+xnmTqe527H4LlxrNwgZRS+gjgETaW
0QNHHJrNL6BHBuAuCc56o7yjywqrA+yuLVxcO04E2Zax2673AVdARvJfwegz
q7bZCgeWr7V61nqPdN+h5gl9Ar3A+to61OC+EJwnbn929soSNYXZ9jbKEOYe
+3Pv4gWIBNNUDoor0sdn2P5efsmOIbR2s7L32hfTpnt90FeqECE/yZz0oWzH
WcOxHDkjnd9UKLwbRaq0x8S8DtFYM2p+bhyHboYBR2eiHP3+m2sIekonAqoO
GLN08kDTVkqK1EyQM8Antc9f7rskcalOi6wGStrZWWgidsN/iNGGHF6DYHAi
Lj/rz0u1b0a9nUSJLLeq2vPgbZNl1veNZv75W96nJnUhPJd6VppFdBDmtfG3
q/0zdDoYjrbUiN5kHsvRAq02ciyZUSJEvzRRyf0MWmw/UYvFaNl+zYWx2Ato
Dtyy5N9Q+fg6C76Pkn3pWr9Q+hwwpQklnPSZHSUelSKuPWAWytssmnEOUCgl
lkzHki9yeI/Wl1QS8juuh6kPtuz4RVzl823qzH0MxRcjeMGmNtnsBIVmEqPj
MrcY9ivc3sd5+rNy/C3qJIMT9HP60TfWM8h28DzASNFzVSx1nEh3TOlmC7RJ
QSDYBC6Mm3RxaagVCKM31Wonm7oI9aRpLTQTZLgKqzWx6XgyRoz/XIynoA3y
7/yTaJyaXrT8wcsZ9Zy9za6ED/yMoDRk2R4cSPthpkOwdI/vkRALFZHSqMpX
LO/arV/IFj4NsIApk+Wx5gUtTEYDjWAMt8fbAF7LNZ+wNHmiP/awUiTJ4ZId
gmn0PB9nliQdNY2IwYgLXo23/k8rn/amtmYmmj1IAs+e2IWyd7RjHL1fLrQx
iNf8EgFzGerK4kWd/ifrzZCSHi9AepzjFJC0MJZEtqgKqS6MRMnBBByI8zNZ
8giI/9uFZFNhIvLtMoINyw7/tQTtXLF1xxSyI+EssTeb8jQx78C1uGBr7Qui
344Lla9YpjVyoYwLrKS+FxE2uAvewO8GVm7c/kfCaEN0JwhNVwYlxgS4oTUE
YcO03IUoQa2jhqBDctIlEjODCqbXaoRcIG51eqGkYQMiZnJ1DFW6jDWWc587
6QTj7XtHlWOA8H8WLtRtUlMxzWnJLJmUMccytTh8zAtxaaBj8Er0Y6q7vvjL
UwU5W50AgovhJl6OcZmiFEJdwKFVRWEPfMqMOjxHrooMIBRWJwCIHYPdzKAD
UqmPiWEd8oRVjt6jTX5Wu9EAbN670p7sDjLKAvAk3GmpB4lOIz0aVMGlMU1g
yJprZVBCMMHDrLWrcHFCn2cwS9RiWwBlDPtcgtWyyctuK8qy2aGO5QYNQ7mq
PyGZd9yEVdkXDQLlttNCfqX1aMoqC2rmJOhugKw41ZvucWFriKZBjcqjKyK8
CyzF2wEPRqgBekbYjZ70XghvVZZCa6efH7denEzw6FkCADgF8caSUji9oZlY
XI3zunF7SBdx1AZnbTuZ4QrZvHlFGX8n042zPjvS6TruGXbJFrSkpxLM+4xX
GJKro/U49n+RM3ztBa98zidMcoTno668ax+dtQDcQ6hcf6Nv8MO1BU3Ml1i5
4PedSAo96hNbSxrUVDpqNj4Fr3fC25O7N/pZfHBB4XCT6cBwuMDq3Wv6oBL9
ntFPGxYgFVbYxDsq+GaA1f/irZHFYYxJI+qxMKn3Ei7HtdodynpogCNs+fT9
Lvf1cylHhM4zA6qdwxKq+jXVVbX/R3MWeA60+D2ZNUOdUQ2Gy4yvSKZTaiZw
3d+R4vYvoOLx3vyWRWpJBo3qt/PMFi5gjODUxGuUNJTuNDGI9m1pvjJxJzA9
X+JKclc+N4awE+m22jcKVWBlqyAGrHnuoJRFCxjUo/lJIDHtROR92O9IbsOB
kFewJrdaxKLcs84ISbKTjUUtAg4nJ+enywMKSESTA3/Bc8DpyyYlfSqhKu7h
lVZfotET3KwR9bPEWsmqiLcuZ15unEz8tYAACRz91x5fvoNvKYoWJyls7bNR
MafTgIV+CGTEwAx8ThROB4b29ke1+6cObO1cdIruAtwSVKFvftzWHN/Uz92A
cTJrJDMXgjr3BBB6Lpg0OjwQEG8p1JznfW+7EwvuaQtp9yDnu9Tkf49GxHQn
buro9Dl/hQ69XdhTYXiP7HvAiIhfxX+qFFkcmx0+QZGXW3w0HifbVKTknZzR
29MQFPW1/Nyb81F2A0nBJSzD3xHcKWdkLlGtOn1h5Ig2QwqIM6a6r8N6pmLX
r9DY4YG6Sv4oHGs8j2a5+CILbkHsvoFbD6hy6Q01Jtjv83usIu25TY4mK5Mq
O/EJXYwU72LdWuSw4a/jm0fV2zVX4lhEYrmPxcM3yRc8y5UENn9exDoBjmn/
Y2A1iLatw2UrEBkZE+eryzN03CL8JkvYW6DU8wRHrJq29ZO1ybAXm13SwUfQ
lZOaqTxR3HmNt99foaimBC8F8c1v9zDFN7p+04FzpuoW6gWwJb41Sm8sf4V/
As4x4k5rYlpCrDZVXF2S7O9Y2JvMyf7XTLnavXMMVpcSQlPJA++lT7HwvHXw
F6TR6gt7g2jy9uAQokhjWaNKTmzD4WQQ0oT04URTGEPp3Cx86EGrdqo/73Q1
G7L17Ms0K0bNi/fO8ZDZKRnKudoIJY+6GDQzoQBpQu/k8rMyGcMYmeso3+bh
j4rLKtvptX/fLZCGb5LRHxj91S6bO2TB3up9ltiJHWNf8uo1HKvp7WhgNLGd
+w7YphsXXKeyEoXkckkZ+hBBEwj71HWNRlQGOrm7xG5wlapAO9ZXDvElTWdz
4oiP24Ac1PBRm9UCzkPZb0LupHoz7QyF2nFzX2tdIXRzhOJ2t2n7C+84t8VO
cskM0elfD6k3tqe4I9QecrdIe9WB6/BMcbmvwcvQkzIV+ePOyNf0MH39QWnJ
iz63mvEd1Xjs6UM0SLCgaLVYjtvBf67cFZ4kvwDbN0qkbAFISYubQszdp99T
SJQjjCkhyT6s1rl+mmbb6VshYAmaWiz0ZU85M5C5ZXfe+Gs6XiloK0lMgbbH
jKXpuYjjXn6f2gbkLt6Tv/rGWipE+d+SQ2apdVz2pa2TL7+EFlDPNTYkG2pJ
d+X1NujGTW2auYHnTNGB8HbOu/Ig+A8PfkzPHCtVGnRy2Nxl+jx8V7H/87LK
QqvHLh3i9pSyoRZYy6zPtJG/cSg564JbY1rmBY5hP7/5LUARD/lLc6RO+JDo
7TZZiv32RKey5BoghhKAwlQNlrNssnKhTrkrm80Gco2zO3UX/12M23atkM74
ySj1BAvuSwMM+pTL6RTcYFNw8h6Y54i5S9sQNkyRP6Gpk7JkjzUPmoYzDEBf
gcQx58CZXI7yuDflDEQe5Yg3ewrOduHzMGghhFsjcX5FFC6z7mrGrbF4hKu1
CG0D2kmezmVHnWlC4bDgHAxTsvBC3IJbYQuGvMfLBYkgdcZ1UKVkrLxUz43l
XXfBFI6VRJtLC8bAH0OyXl3NXBpRuwwwn2SUjuovlYZYlD2kLcf6uSLlsSvw
ZZzH+jqE7Co+FUWU/ku3K8yTvb5aijjkxTdgQ1vG5dhi9/Vls1LttYfcyXuU
fpFYBGTERfFQck+n5yQY0lML5d4nimIx/dPRfru8okNQTTjSgm71xcs4+/eF
HtUFqB1wetCnoIuszGw0dLzHz84F48SYnC+BiLj81VVOiVo9XHPPBvpqcLMM
N5A5eeSYJUijJh955k4B6gx2+vgc044VlzgS71QUOeuTvURzp1A2eN4uywNG
7vUpn7EUYERAQfNEoOVMHxpaGwaBd21KowLRZOG0fj/S0ZJkTTV0lBbZwVg9
9wYNr4CGiMJivNRKC/X9itM4KH5TcV5Wq+0RfXvmqQuiZXSQEtfq7lyZ399p
SbzzIGHmGEHjABp8O5i7ir/bElH4jSL5I39sVQVRgI/H6oNyDynyiggATol4
/K37f8Ug/zxKw7VYilj9kI8WcGVEgo0PwG8Ha9NNEipbtraTMi7dn1GU49jO
W/yP9eERZBFYAnP2HFyYHs7J6GXG96t/Rz5ESotWBYAqF2+TsALzYCRf8YGE
V/X7Ark/TJHQGYV11jaqgg9/7ML1bFeAQv8hyhZV5w2mCkbmuN0v6YcM/tLv
MFJVz02PLT79kqFRveHahVBVFjLsQCEvoKI3kP+O0AGqiwxNP4s6GyvELlT8
oHMG/+uuO4Dk6Zp9IHj9xiJCznH75KgecWml+TnJO+exhbMRyUo+fTxnJXOL
2lK0H630x8NOD7aT4U/E5LpVBwxLLCMeA+ofR0R2nLHBZrNVXgwsLFuA9jp5
RIncmmU3X4dwRGB1diwjKlonAh0xGRK90AK936yEyn4oMzdKw7421fof22AV
WK1imcBFatHP//2xegnrA+1xbMyFwDoFYmfRwOsaVxNCN2x5BrSJ12SzmznP
BIQXuAlZfOkl72kDSIV4EbOyjGqecNWQt3R5jBSQrQ1nK/wiYqdHNPSxFl1f
AWeHXW1vMoXkx8qYZtBcg3kZs2f8gAsdOMw48+jHxk6dlkY1XTC4OF+mpnfU
oVwBzP0deRBgbuQiFML0RS3jvD4PGPgSAbcS/zT2RaCiRXGSoURImwHeRfnn
ExpP5SniKZoPELXXOml3Bahqa7hDhGjE85V1e4hDXED/4CDQV5JBc24rLMT8
xdvzQ/tln66JPlbEIusuEiRZL2gFJbSjXrHmWDd07t2W27tM+unuj9/a0Kzb
TNYyMKJjvC3fYn0MEYeGWsts/e6SGrnA6wavd85Q1ZDVua/M7RuwTZte5Dsc
WuKxStw0v1OgD8RppD/oMiRVpBq20CJnH3kDHsyv8c1iHTNS5QHDL37+QlaU
vHJapeiVEJ4ZY6O0N1h3rpZdjjIUTDSRgwoRrF1pRafEcNZy5ZQd4oSvDfjE
1DymprHxeifPgURp+5QDsGv41KY9PubLmOMdhJIdeKL1wBemm8t4XquWxORY
LOne+0xOfH5k3idPafMhY1JtLeCuZY8Us/QPfvAFMzQn4zwEIwHvk9iDMoIm
vGQJ/gD/2Xhw1nAmDTCXTxxL8fveVtTQjKk3Tj4Pk19n/phkB2Lb0q5Lqjbh
cyeb+Mw/5Rv1p4CcDvF0eUs4CPfcRErdL28xpIJy++kHQK5KEdYBHs1y8M7G
MgvT1fJyI2gVaTGbEtVmb0HLoD4OfiwZUX5SSruI5SaC8uVbilyIJieFc4Ep
sRXwTdEc6AlUfKQ/HrLjHBfZIxH6AALOucxmhDDq6wvTfDP+kW5hJX4vIecK
vD2w8pWLGoWXMkEAvrfn2heo2vV5SuY1rID1Wru8hsb+gpyMGo0xOPZietSa
YLUDaaaXPPmmuuVQ4KW52xj6DXm5g2xRwzpT0hHflalnelfyh40ulRcIPKiU
stkcTM2p7JrG3yWyi3TvP4Lh4qo9KFe6SPNK5mLvqb6Y04qZ61llRwJCNW4o
CSjq8mDorDFmWAKe98hzDPD3prGtJ1+2kFUQUpbPeutbPB+ifNYWppXGiMWb
WTxyFlA2nhVZvryuaTbRASv1sMu9+z7x+shtgsCl27rJu2qtgaUS0iMJaI78
jnxk9gCiiC3oCG15+qRcNvupdFNZPsd69ripewnHsdAkIrwZgh9VQLkRz7mp
6qEASXWf2PGa+bXd4F3/3j15fJl3gOax40To8z56v6f0+RdSFfjTyunNdJph
8CfTiA9JWQo0Fjmr2n4MAPMS/2N5gUgs0udiL31SO+PIhcYfdtcgNXGcQnjR
lKpw6glnFXe6jh82LSQ36iqTl3ELdreNI+kV3r582H+djztmPa21yYENvaVW
LtDNmSvBgfY1b+yrJrfjjw6knoNMGZa9AHY0YSCWIbXN+CrTnvrf4A0O4LHv
ElU3gpAhv/kMWSbeyhWztdDUnJWQTlH4M7zvzDyudno3N+fIxcADMsphAxoi
sxQ6Jy69Xt2toZCvmIrvoKEaoKr24mjk8//JABwvaDTs6Jo/3eN4epdLHWWd
FhgvS2cmhnD+VtaGm+3XwD+IseGzvQaYpzwDSJ3BEfLM6xnBt146ofOnnTmw
2byT+J/yZlDY1NVmDWRfO0gUqOux04BRPo00FJn021NvXba4+WCBwSmCb/VN
OWxPPs8OvSiqWe3XZ4JwHICDnz2r1FsSa9xA3Pu3gU+tBx/UZXBgxNFS8jeY
klqAAVdlG9kGA8gzHCnW/sW/BGn/AxOBf49RmRkYoins015Fizo46tcmQre4
6kALc4jBK+8V8LuQQcceYW8Pq/nQr2JlIi7yEHh05wg/Y+6YYzPTO36YB8Yt
DyjmmQsTKLgjqy7hndLYW+uBFx7sZqizj4mcInD8ig40nPKdEs6W/XvCQNSn
RWuR8cNcwo+vZJc00hFXoEx/b2VXqf336hB4P1U0K7lQCqWwyNdl11GiJJ+e
CWEGu6ROW03Fa0k2Zdhr/4hJn7jvL7ojCknDjmkqXW9qYSGKNwbA+vBQxvTY
ZgqOlrITB5Vcxe1UAj7wZJppaGoJogCNR80ThBJaV8uHiIarK50OXrCd8H6z
yEsYylbI30zSeiINMTrOG1+shXI3ZAweWQu3bfkCksW3dGnPsSlo+4a60wAa
+i8SEyhnLAmknTi//W41vVyyAZXMlesf5roLi07rWQqu66aoYqb4/QHXeoOA
qdlQQvcvDDZOLIJ5VGi8oKwodhfCjdNm3fBExqpz1GiXOfqpKtxiWAbJtFC3
XB+FQDjHTviTHIptzTADmpLIJ1CQS0G0sWZaCkS2EnmX7c/O3YzbUjqj2B0K
soADBi+QhdOw1ohJAY1/6Z5jAuNAsFwjvnyKFBsNOcjqQXgNfqJmU/P9+faW
O0Y8v0Ywgb8rifDRfcBOYIyxda4igF0crK2zQwUSmj90+NQgGmtJbKo3uN99
3Z/jG3gXCYqkeUddlumoxxCM3vTNmQENMvslU8hVg8w6135/pG31BV71hoGh
xggxX0Yh2k4vp1ta3hZzpHmJ3ZJ/c+xQaEtUtsiW2Ji1OXdGK1B3dZXNf7/K
AanmXLQcjD+uwp7vJL8rqLP/vBPVTLInFrj+OKYPLrC+uqOzlTLNUPmp/TGn
Dxni/PUE08l6rVn4veZvBj5Q0lhsaq+IBNv0js2E9uf94GmbbH+awG6VI8M9
IwQOnf8cJUAgUr1CfVktmcpX/8dreKyB40wuYtIYsAo9/o8QPMyYdcgHyIFj
RLr359M98C3X4b9G6ZpilCzgTKlbWkMQrDuEDJkBOTeaeD6qsJwdOzayk5f9
FgPFzgj09+XIxphoqsJyP6LVCy6NmDzuufchgGii9JBxjCGfYtaxoVuymj73
w2mVfdAKxV3ByEUC7RhNIZvGlwOC9U1R3QB+daVT8UN6oq0K7ZP9qq4hBNoi
DNrF+tPC4WV5tbD0P8o0I0i9R01mO0CwWtkDiW7jhRPXsQWwpK48+WHSP1hc
en8VN4qiSkotvn3951rKMV6gYgUJQm5UMlFrpXVkRi7HcXpFo9e3HXtgX6vY
0UV87wH9ZCrA/4jk98ttXeC/sl8lbnBneDFL28cGZ/fk65ETxyasAor+GkC8
YzgvBjPV1qRLmXcEk87ry3cVWBQNJbh8+7HGizsAFHjLhNYkwD6TrtvUHnEn
XMTUlRizneVJh+Eg60Y2K+2CJg31PYTvLN6HLQukD8NOH1aR8MXkXaHr7YDW
Wy8gow2Xy6HWTmZWr2lNzVn+Q0QKqGgVAIRpJpeMNw11Yof6tojuSX60q1uf
UVvu7gezE2lMNSnsWpIcCGbxAOWwdhRwWRm6EgC8T2EME2ouEoKI2BvScjqV
KzywG+T6vfwxkwsxD2MjaVjhhxnYG3DJfo6LDu8M03hf9HkOsp154ppPCVgg
LOAarp9hmtBAEgEXcR/MPAplLf1eftbjHAAQiePbvpkDX1ElrY71Hg3onDUo
0QEYmIPjuKIWFxlW3NNJuvbUalYxyyf+Mm2ERdq+WG0JDu1nbcy7ip6lXzQb
v4UWQutpJYgizojIBCFomt6yCfVBE8+MJFKnuzGY7IrozySPqdHd0M62IQw6
NNRw7rQmQXYrVJeBi+MskbpmJJjICPoMXUB/4NLz4gVaUyyJcA4MF3rLjB05
OUgPsFRUK6nWwCmi+m/QNweFdZ221mBqnvihhloXUtSbGq21GNJwc2Dl36KS
fUiaKOQyg3NmVW5NbrH4KcVEEx2tDjviPOv8K4uoyM3agGMMO77RQh9caUBu
MEQOzR1FYdKzKAvXOMhTMyHcQSEfAa6WY4PtuxVhJtng/KQZa1lletI7s600
m882QM7nqZHkgMqWTIvA+B0UFpVHcTYv/uzLVaqZeOxgIHYaoSW0Y+SbXFAe
Ci2dy3bw2tbPT/73+e/mvJLwFKhMYELXis+ioyHiA27maZHOq4v0Y7t5sHzf
pC3CB/HBIY5yDhJARnr6hCsVtmZQQFWxdBkkIdGUHUtRHucomnZ0oENNkQYE
H0q2C9st2/9ZOUHRCXDI8BpkGDgLODHHAIPt4t7C6Z1vGBwK2aLxu6XSJ36+
8qoVM6f0BsjGwpuuzRZomg+pSn921ndhmqKZOptUmfvT2k2L/k7JtqyU3QvZ
WED0eoNsaxuO0c1yaFvfjR6/A3OhYplKHwEQRAcg1Ke8w6w6orkntW/goi1E
b4BS0p2lK0VZEW+pzk9MW9HsSWRsZBwnZZxvhR1B4AGGQUA4dprbCZ+6DsNf
nWRL5b1aOoreaW2W9lHOslRMylg5jGHW+jRZi5td8ICUqbKt20f9JL/fdWAp
5rdbj46blwEwXOa102EFVqqujHSUcT/KAu5Kclsq7h3VkUlUvSyDVn/5dGkS
vl+J+Ps9H6o3bU7EW4xuE36V6ret9q2uw5NDY+91YCJ84lz6brk8ShdyGb0o
bRo0DJVsBtmLsfrfjfNamamk+21JoxaSC2GfrhZKARl24rcmCSZSnmSl6uYD
qNRl7br+3BYj+1XBHeDXQYkQ8ew5+g02M2Y5Y36S/A8WIIrkMIolo67zSjKm
4gTmzS6NRKXaJyoP1xdF6Z2NgHjjODCoX1fMVJdfhWoNvId7Qae6+YRie/jT
3R4MQLdWoQbCJdKPqhY0gkbdkuJJMGzDjCGUmGYg/InIaMjblytLHnUakEem
r8VwQPy3EKZk0FBE36xbsKYOWSYc/MymX1Subk6LdEusrsnbgU7WIK0A2JiF
ZcEDfQc582RXX2mhH9AHASC7OEW6DKC3X6RdZmJEFYI3pGDcNnnF3IA2vBE5
9VaJKOLQLqn2zcY8vqg1GxWaNonARNF1gbmJJK9askYe9osc/+LcKB9avfGw
UjGx8VO3Ur2DEx1MwWBq/XcFC5CZfhODbKMmEO4cCGBZZgWi63pNt8omEjYn
hID+/dCKZ1kYUEFfgrLeOOIcfEmsocV30ZQysgiXiTRVDblXDjqsvZR9gbVd
RXbCn9MYjzCRXuUejSuu8fn9H9ar1GODgfPS5AvK4dvdVT47updlhFIF0Z/5
hCSicmpvm03KmyTylVqgXj1GuCEJGyTqrqnJJCUbMjzNxj8PymAxkW0f/+V8
ZwaARbYUqCOYygMyPldRuDoSYTGumQ1/9QHFClASj9QAT54JLYoBt1Rg4nV0
kPkjwTh1HCzbq1/xiJX9zfsjKkr9GjJV02jvf4xtl2kQ7Lp9XWtV3C7ie2/d
iKMCBs9ZSg5KggWSEqe2bjSktM9lo/wzpPoy/phv87rGVRMfEhmY3RaKafr6
sYlcMA+zUpAfdOuLxIoUSxxIJ1tZp99o0ncTCBnQQbXOusSeOb0b+dwpDxao
tGiDhnTF8gVxjeGAtUcT10u1onrRSJZbzHHVu4I9YJtrHPoQS3IMpNZnmW4d
pdeGrbJXgg6zbGAZuTob1+GYsYT5f3pXivbvYKTAEXJdKPGL8u2EN2+VEppG
htKTB3sP09O/AxfKui35Px5H4t5UKN921KAMc6X/MYkU/DXK0crhdfKDYqqq
UuHsh4N6JJ47J8PABbs0mSkjO2wigckmr+32RoAp0X2Weg7k89zOhZwrqvHD
S1tlxMeLAQoJOAoufajHENLtJ03P81DoeE7Wk4l9iI5wFTkzzRgVfFXE/tKj
Y8HfvMxSU31mcjwzpSzGg/+KrfKpAKZzcCRhq2we/xtDZOdQFMAxGIfzV5lj
VRUBVAg9Xlldj5aNijtZobkPUbcZ8z7Lcrffmh24vV6CoMpeeu6SF/FVuFTU
zmP2CJ5mHWhJPUukHB6aR04dyZSsXHcj/y9iO3u8eljR83u8mtJl/pw9Ww2U
vo6cNpFWjZ5zHj4omaQsvwO6jzMD3H4bW0rGrCDHP81ufMLmQ35ecO7N3I+A
iI2aa4POj+LAaiDh6fvc3G3PwUX0BOjDo4DmOnW21+3FWvxagubMIyNdmhXt
1wcjDxD7NCLapQMTt7VvkV+GQjEm57fQ0YEWBnwO1AEBLS90QDecLIGMlbep
3845Z+RQLtK4IJfCYz4QdjHcbDdKWuHN+KUuQKDF85gkeENUQEjDJqdHoPgt
e81ZEEFh8/zzxHAuGIjIpud8wQoUxZfzTV7a86DOCIXqeRXgfVdcXSu2Geqe
tOwxi4ESgabifZBhJ3gUoygRttjiyXPIWvQ27N8qKv3a+USmL11JexrCoTS/
GUatysqPc6BWuZqMkaFaCUtStODP2+y+CvVO9IrqdEoVVoTxUHuHjrmH0Oh6
1yoG9Udzatb3rICr9jM75vlEf3/fAYLn6xxZVefk+FchU6bDDRtykkhidbJi
sHLuvL/zosUN/8BbX0g26GgQQbmeVqITy/YZ6fbYXO8S7HyDE2TGPvxWOSF6
fiTkpCvgWkhIDzJ65GSt84U91mEvWot7CBn5DAwtT9Ja//d4rgNndu47Zs8m
EFEZaEMfZcZJRGNWDbP+0jnKDvBmvF6baGYgJyQIaxEJGpoJMzULnVW6tauO
mGdSmSL/z4+K9OIFWFisAVuhyhrVcGXZRKMyXgJO3vamt5lwVrU0IwsQwLN2
CdlWhrhkIR1bUGmLzvMTSjm6BFet64MQZLBmgb/piroYJ1DCtSb5wub0bzVp
0amzHANWTUd6WdmE/ENaoFcTUc3IcorVf5rWB018YfMpbMyxAKmEKEqGiBUJ
Xw0AcUJ0pnYOABqTq6XvocAa33t9QppXDf6i4RHrIjyDuaIv8wowvMTwUnRj
U3kHcR3Sa8kmqB9kbgC4kN0/lmCY4ORFnM5Lk0Qiz6lSlSrQn9HEP+6b1ZNk
VzsL+IHLtTafQCUuUrUUVoMi4rx3UgHyTiWEXd2l0BbQ9lt39S/GDVk/XpJ0
vxIfi2ms/TIC+oJ/o8kCU53F57X73ypw7Nc3SSR1A6TPZE13yBqR1jhQRBmZ
bQSp08MS5iM0VkQ+sf7WevyiFHS2k8F7RXNLOBPaS5s+yOuQlB3vp7r1lK62
cH5fMzYC6fj7uruGZWe29Vpo0ejivu1zuFPa81SfJDs/txYEzhfcJBV1ZfxK
XTDYXEqkuX/qEb1qNeWwD38nUfd98Pk4ry+sYUt3+s1ihjUSL3HYhpic7v3x
lkBtyU/FWf95TlTm3jihOPbQ/AGTZPLaWStYaJNc4Tx7GhDG2V+Qhq5s5jaX
bRxbksRkqK9XU6DNWzC0Bc6ktUOvxJzx0lmyzIRQ4Fxy5u/50uYRQa7FvVo0
BldX89hioOV4l5+foxJv0dQOGyoufFOY3WZiNL18QdaxkWSg/YbBeiJNxkup
0SSIYOM2aJ7UrgHgTRjtcrbWVXZjgCePRuGDm4ffv1vw6pEBW6gEfCM19fue
2FKivp0/U/NULqbPsPtjdZrIJbo+PJP+7BWSZ4ADaRSPjvtcKZ7gLA9iHH5R
catKELLxWirHLs3Iv5UnuLq6D7gXcyUTk5TgGNpQjxVGa0L5IqPwkaPdY4d4
k3oPfrSDuedK4Z+SnbGoebRyVLqdduF1c3PjgkYtMdBwVKoZqUAVROpSbYAx
qsBsKAOhbOlZmtUineaiagCMrTyKN2/ag2S6O7zhOw0gLW0yFhTbYF4a1scZ
3eWfkgVfEzr0/ZudO1SWQPmS2JeUG0qQ+56v0MC6ZE1QArju3WJ0POU1aaS3
pFeqVMrA66JbapJO0M5S633QT+UuApN+AbOB6bQg5HL6zJBasKvQDv+uayl2
P2VOpPWxMAN+BjBl4Nwxk1Obwy7m5OuqX157hOIVJ6hBCabL9gvNU2hI3Qji
dn9F3+6GL6G+bVPIxye0H+QHlJ4iqc+KlBEbgvLk8HGjIlE9WMaLeTjl5Svq
XWPwtLHDX1KQ4NHnuYHKUY5MqYI3LrpVDyFRShSX9mGu9mip7/QnB986E8DD
1e1vW4TNFhZKRwm+PMt70SFcLWVu7Z11BOyesIe7VQ/dy7MO5uolgH9riarS
U0Us8xJ+0vJMXNKolMjTsz23iTmCLe8UO58eSiJOnhNBD8BOeM0yVvt6To5/
GN0YYx4OZ8H3/7Gv9LHVjE5dVg10WuqvYAhoH8GF4KlzCL0ZPdaI9xUBW80K
/0YkrDeIAP+bJwZWShVu/ETtJd7trA7eaO0SbO3S6Bsojl96wsIlMwXNHPBZ
7PHsFYsi3s+CQrFO5dI9iRjTIgBDy0ORXTeLcU4LgUcNZR9FY7hzhlTzja7g
eTKiX7EiHdhYJSXSgxA/2BMsPAeuy9/OJ7z2NpbsmXxH9N8Lc3+PBnMRnhZi
Moh34vzTp8EHsvb4WNjGmSmfcSfS8RTZr1wEQQjtlsTSB21VRLD9D4F72TSG
0m4eMKeUsl69MNMWirHkZksgXhqo2WcNcb4NmnL1zNSV/qzcCvineN23Tiwz
5kmJJbvpmz0q5DjuIQ1yvEc6mxmYRytR9YVhT2Iphvvs9KV3L73Z+cY/JxOo
DNsaOAd/Gu4iHhCwhtvk5aP2m8p0l4c9DEXNyAt5BHnre/uTjN8WBA5Cpg+q
SoBa6ZlXfko5yMuT7i3Pqp8fs2MJ2F8n8cyD7Sgw64PHaQVhLZnWyc4vTEHf
UNCk/03M4uJ0+Og3J8vR+hV0FKHHSaEsC3GlxE7KhbJ+PUqJMlwaujk80taC
UjqullgOLzdSqPxVGM1DzHbOBLMHSt1UR+zPMiP1vVjzBPzob/xtbr8iRE4r
qm1ew1RgQVmg0/HKt8Q1jNw9URXXa+KW09wG0I5Cvd90a16ZATy/yJSW528k
nvR0CNHIpzadLcCpMCaXpMPJdbqzEb+1Vp7KtgsdVszWuQM+mSFW8M7hwTm3
58Ckv+JuNqWO5cfDn1Nj1aFDaFM6JFFu4Q06W87ugslKJSO1ylGKB2PEKER6
JXe/iWQb9Rmnm7XzM+Qlbz6U+Nf9f0rVDpMjj6niVtUzfwwZWFuMPPXVvIEj
BdV/EtXOVw2lcMFG3nNDPEITdQn/pq8TM0/5DMlr/nv28u/2SWevdGmMnCLw
/n4zzIU705aEIkGJfLcKvaZTcBiqF3DsZY1Nl/99WXJuWtkfH2DnxkK8CMCv
0MDGZq8/tQNZXSLWBWAywTUNGjMLV1qRV5H5ACQgKgeM8vImXxXCBKxBLjKX
f929K8cdvKGYGWoHTrjcTjYFihUH2AtbPR6H0XFFQFp349pGi1dDAtviBg5p
q2gByOqpAQCX2GYUGUh1vIgj0LVW3Wujj0KWW98OG/Le8GES6e+grHk45100
1dxfJHkfG3l32ZRqHirwYLXWr8WjPg5K4AnhZcgYWvcFdzlALSA4/A5XgbSj
h5hsaGtG88ecuzXDA0DrS1AFlCeP84jpIySSsfeWnUUlRPfMAgCO/WNNaCZd
2vmYvRCX1iB1zeJ0g98uL7jZi6zyjJcgZlE23b4Xd7Xuc2AnGNmuBwWOkoWk
cXUoWRMZqXKMIvlj1dQw2v4b3CDSHhlotTDyJQysk5cxyBtq9JuZyKNTUk7A
4Dmsh/IcpYaCFavZM8PmnpD/udHjuJHA63T/AWTeTIdQE402w498XHfynJ56
+Mut3DtSg0LhpQm5yxbeWD9xDpfVusPirEC8X1PvgQ0Sr1cLE+qu+RxbuY3M
Y1ne4Z61r+IyzHyPAIyE85BZm8zJXs8B+rPRQIWLq2Jsw1LhGJmnNS5W3Ra8
dOqMoLsaF+Hgny3rXOiPXMUOfVNm6VsCdUP1QRxautjdgapmDmRkdndl7nwd
pCsIXZxOcMImO3yIGtfopi+RfacJKzejHKcfVPEaoYy+HPR//utisPX18102
V+w8L4y5a9hjhYKodb/QIV8LsYxAZJ748HhTJaKcBQT6fyNJ4Ypadvm9r34p
x0j3X+soVA62QtRtqUwVDb7v7e15RWaClI0nCem+DCmRFOgeImY1cCeWqB3h
/V1xWh2ihr6n1xrZBtm9zBWHWdcAfT/6cb7ibSi4hC2IbHwsKOEJu9WS44Eh
eVWUW1p5DM1Tt5K3PxAs/8pm9Fw0IoP3+mPdjqGk5MEvigLBqTq0v5S0dfpP
H3Hg/48rAlWAmp13B4FUSNBHLp3or40YVf0lNyZol4pA4eH82CBK3hYBLCRc
YrRObetisWLzGmhEj5FKRtTw2eX9A/juocVnmhRXjYP2PJcvO96K21Zim8ai
bGWzeROGxa9bXiC3cLwfGAlWrC6hoevFvbOj9WbTm6ZBUTkQZT36QbtTtc0p
fF0vtOF2daFdYwPQd9iuW0gL+N41syvPvn/XADfOVWOj2ipftO9ilpRO+lSM
cMucuXf4RVDxcqMWkaa7dBfOuQLrsALg5Hq2aLJDmpVxMW0oSeCvLtZvq2/y
wvitrCRrVvTa5vhx/JQV3FT2sri/Mdg6WfJAUs117+jL91AT+qAtcu+2ZsBa
MBQpumjakj9G+imjy0ntj4XHYUcDzs4AoQrtT2dpYscUO1vQbzVnWdZtOuEG
igP2+Lbr/T64aJXD5R8VKBzRVIM4YjyGHuQWNeOBdtLgnpX9qYT/WUrc4D0V
xG/r7N0GHkUn93VBfUxefcg8/tHR3jzeOP2ShtK6CvtjubVE1xbtWECqa+XG
em854ydaVi7Ow3RgLbjJV/tA3FXpSvklEBcPxkMzp2dV7D6KkmNxrlriihiW
ygFPFTcNjwD/YpcW6sjMdxGHZ1VOfxR3zliyknkZKICmu/xamfBa5Ph+7vkl
Howke50Rl3arP15M48ty7WNKvCLd08SmJmG9BIOZnjh3C+nrsK/pFy51+eIL
w0bpsP1dMzQaqaBexWkZFspc0t7RYTeTGFUv4RGF1KS1zQgXpPK8wY13RY/4
i7fvzZXeehky36wd/o3fkaX1OY52JlHwTFki2s0IOHLsJBSh6VdfQwNh8og8
invYY9LKjCItR7k8C+sSd5I7q5LPknVFGMyrhMtxyJVU51DthXkwfkMk/Gcb
68ABRzCHJZ57ekA/R0/AAJRBQjtc1E70I9z6CnXBVlhZFYx0yNxHZIukEQU9
R0aYF2CFhyxMrhanY2nyYnQBim5dFXWl7IdVCKL0SGNshgtqv27oLXYuBoXK
4ZMHnlUx7G8a3KIANebAEwLeB9aFiAXOCS8QTD1C+92i8JGUdaIl/NyfGanF
RVxHNEMcEpT6hwW9UcK+HQS/+dmPlfCSdQA+TsSRw3N82R9SwYOpIB89QPBa
ZK6ka3N1QpjHNVNg2knb5NA8Hta6OL4JLIYQg8rEWRAxYNXpwYJc0O4RLszu
0v+74UzInyJjzila7d6yXK0X8zDQCYF+owDe4hyNaZRFsCCQSkZ7nmVxbthU
upJOdpDcZhy1kR4D9DAeNBwLqU+gak/MDCrcLh1RJB3tmZaFxYe+21a9IFXC
yFSAsYXBh2OKDHNF+9YU0BdORn2cn5jR8aLbeHfQg8m3MHk+adtEb2pZAYhi
JbI1YtBquqfebpYI8/gnvJcxdQI+IFLYL4U/hGjesT3KuMGe9fZmAqAYblob
n5mu6mYYnmcXer2UQy2TIGVv+qEjQLhDM+L9FnngWY2ZosDigZCOvXS6hikg
q9K+8wNV5owwfDBqMW1F8q9xHTa9o9VKJHDRn1n4TmIPwS/fapetLl+8nKcT
CytQw0QB5WX1f/yWv+3L+zSU3/DHGAEY5LaU80vpC8PVNzWeqRf1EvngMtFl
Qm9W89vUwXU1iuVtSJxfSjsD/hBNt1Z45dVEWn92f39TTnOR1pCqHpyTvJMz
tLd9qaADfF8AUPjebnVVlzbjTw7UqCENWyKi+HINOYmlJ6mi4O9SsLdoGGID
7IMPwby8VzeX7LDhOGc2nCQELhhnuXiafG+kCVpKP+CwjPZmelzmCALu4zhF
sSasjFz3OI0jNsG1ncpaB2PUA7ugARMOCCVjmIbQC6olLl9WLKjug1sTle4Y
ybL1fC8YdSjKZoIelNxFkNhSZHkGLqK2WFQ2tQjRuxebae2M6CmcJBR7QLED
LP7owTKAQR4rIYI1HhVRWlmpXopE3/6IFs2fqYItwmfv3dgs4eK2SmKBtYrB
jVxUp1m/RAAFPfF+ynqq9BwOKY9De0gYoB5NYE7Jl7yVm37HzPIXZJuSMJ3O
gp5ZnfWPkK0ZicuvO6wbpEYHpSPHu8J6pn3UIm7NgwftYebbrWj3BbwAijBe
sUtUVfwPpp0xMngHWvP86xOq4bBnuIvnOiIigHankd+LOMQGM3QTwcfNkeGq
nN1zosrHRJs/5GE3bWaqND32s6PP0hAR2O9WQ5nB7o4YjoAeRf630vSSXAtR
19Qbyw5DfiBtDXtNqkkxjHK+Tib3D+SfqK1uQLuXpfSLm84sALi/IKyqMoGI
k1INQ6j0a4Oc9wF+R/mLtesN/YjNed+EGnHwc5++HcO78owjyVlt7a5l/64z
RVlTIcLZc1poBN99jGvs25E5vkKwG1sT+CMol+1VQXY/NNw01RMl/HlsfrDR
sKZiNFj0+QYgIwuS+yEUeAcZRMB4xGolW0KdJX+maaP2ODzksvgp6L8CXv7y
z6teJwLrqbEccGhH9fasOuPfgyBWfPRpBdp2iXqB1WDC42/oaCNnoQcfd+9b
Z2hLl38aZUR1RIHGBsgLTE2p9BpQXhWAyyq/BSnPVtM0i982Tj8VEM0gztGC
E7dHJyZvAAdryM1Md+w41G8EYo7BrcEzXb3n787u/SSEhMibmP2+BG5bpo6r
y/9CVh+rDiyiijKKKu9DRvg07wYe8kXFn1U+cifFoAdHWhwSIaLGM1H1hV0z
QCdtfsUMSfIo/128/x0WDRbXAnKIdnFWX5G6OqCpfknplkGUYzpEyctmg1HQ
clrKIkRfLzE+f2zf7uR/VD2M0rPKj1txotdvI0Vn74Gd3/x/lZ2Fso6NpY0N
q+/WvUFsrHUSCA3AeRE7j1mW0UfIJ0NwsO1+5M9B35k5JG4faTNUcyV45yys
KDaOOOb4Yey02EgiuRG4nmcyn3jv+oxvZ9rQz3i737eneKV0i15lk/WI04qb
EjmZM6+xvcgYKVIGkK5emjdbdctY7sv0ldj/aQd7SQg8XN2eIm8aTGaBeRtR
MhkDELdQPu6JiFTnuqVX7smtjn0e2qCQqlOghW203jzDUjJxLJWj2DNTLu7L
zyOI973UJQy/IItBh1f4EOH2tgYabi9i2Yej+pa3jgiWF5uZnotfyMxGWSoV
Nh5VirHJg+w7SxELJVJVPekQppChuxmzDjjCS2p3WL2n82OwIJznaannBKhA
qI7s+ltqRwvkNLBvE/QsUjcQbrOv++jJdTxamftWQhHLg7zq9+HB2rp6i3Aj
+gwnGot8HIPXMHFQp7U7KvzcFD4AHljI0339rj42lUofOz0Z871HmKAVYyNs
KLuvZNNdkPNZJuw2UAQ3eiKJazLY5NaO4e9Lm0/PT8Uwi2NTrwtKzWBGxKQF
Ti9OgTKo7bgXmhOA1w3D2Jrzf0TUSY5I36EX/gjIpoYvy9F4gSi8eLAe+0Cm
z1YdJWyl06vddizyHJlAsXP5GvTHnOtudgT4MQ74dOY8Ob2BMO3jtbzL4ZaS
tuJ36Gq2BXP/97T0laI3h5wTB31n5xeM3Lo5bRM4B60IzV7chzX7t3il5nii
42jm/COqHmtC3mFVPp57jNJ2dhNctGGkiFqw22hObHh3Am5moh43W+nAxSiz
heV8pQEmxH7RFQ6cM3cmLYAS9qtlZeVfl1Y3B5OFYpWzC6HDVBoD6JwoQCVc
kJ4cnJsbGV6eoWZojisY4Ig03B4joixcKxfGN+FtAaGYELcL70t/z+gO9qcB
iHpdGpt/AR0Cla5ixDPzhzr0rxqLa4/5cq9qzSnUw5s7WB/tYJ5l9aiItDq1
kTaz3S+JUhNfpW6Bs433sfTjjJBegBvQwEKK5KZmg8bgVvBqDM11vwV/Shyg
BGWFttuoNZd7ywFx9LZvaarKXgI2OhPfiaDjh/thYQsm0v5J/+ct+xBQ4DmX
Ns+RLrTX0LIx5mb8yW+lYkbqfw4tg4tPJM8ar3pmu2nA6X1EDO7ylNWmcper
gusY0LsEFJR0ZQPNkCFRprMYXYMNdLZe3uTabIJaPn30zSM+0Hl5Fxvpluk+
qwJNEQ6hgfU6cqClKmfNZ4K2qKpwqea7kPoCwGD0aVWAgn1WeKnoBOzWK8hJ
6ExThBrqmI3wRveG+zlFo9aB1652mWE0zGHT6XTA3UgY1J9PEGed/ZfVURkd
S89UUHzM1kT0plvb1JK3VHtY/id97ateAWe2jS2nWlSWAiVJNu5UA4drsiYi
VjTel6pPycNd/SxqZ784B1d6Dogx0SBCVpE5Kzg6M2v/jgSnVNPWvgMG7Jcg
Oy58X9IiRo3+ID9dUc7CvwRNYQ4ZkVPe2bx/+8qC27lpPDDVnSdFyRGVxI9T
Apj2okWtc31y0A87ZhLdtm9UGD0IUmBYY4reV1cnmDnoWAvpm3l2+aEzhsAw
8ODaTBWvXvtHAstEvuZcSAEMwfamTpJ6NZClW4zOXwLcxa9lfRLFLvFujqON
15JJDpiQnIi+M6ZBBJVs41ocor3RkxcxLiz7krp+6ibK4qsMclT5tvwTQ4Eb
ydowXei/P7r6bLN74PXD0mQ38IV0mwN7iqmSSx/BZnt/NRfEjZpv9JDx3mNZ
ky6xJEYIklLItKh27fVYW4OdcH2Qvwe1UWN5h2NiVJRmsrFvaGApjQOxRxMb
u4nF8o6+OlNqn8XyMHxmvd+BaQm2pZhhlWawuoD8xsfAvYGX2vyLgwIL8meS
2VcP/mcPXipR0e3GGzPmRj3ausi1N1g6vXhoCZe+HFOpxUJ4OONl6/+hHKf3
cgusNFxSNO4NUr3IIA+RrsfTnSvlxjDpJtIXu9LNPyrNWR5+B5dSRI7Q++vE
iGxtnXZHAWZHgayB9rZYxzu/d/4BKiTxt1vPn8BPKdvKwfFs4A0ElH0j+wfb
H7VVFq9uS00Fk4Bw5Ekupz+P0zO/lkxrRk8wzJmYknH+VTPyhsAeiwtnI3hw
W9ccwWtiuRcxvy17qACKFIvxweuYDA/RoyrajorkBKm4vjjwjoJd3GE5mMdQ
u4y6NEZfwT1QrfImltT/1K2xQuW1CWnNAdzeNElgfNdHcE34LrGQHDVUH3Uc
vGh26Ws+TWyG9KO89xKJ1QwzKwyrrSZp7pWYIohZqArcIqrTIK/OnBhdyacG
el4UEhRvhRb15T8+5Tp/eDc3utEC7ZlhW4rBYHzJJGB3uooyrTFaNsBhd82a
Q8WTD/MV8R0WsWzlyAL0tOP0sOtC44K/TNpNKocfczezNKKm3ACCiqbHTsTJ
AfQxzQ0Pw6p1MavLHddcH7j9IjtetCFvOOlExRrFf3wGE2uTDwFy2NT1ncho
mvd9mZMbUpbAqLNBAKyisep1nTtAFrDkPkKdGCjSRaLzu15yXUYOuAoxF/P1
tk6ZCE7hp0gijHsC+DQiEUXkOhMKdfob05IPNYfeM3/1tGONasULgNSfAOpW
5vznLwvvv2eAEjts/KHZ7/Dk0BJ5DwYdDv1mfFKZUwHptWfnykOcNFIWoypP
l1ZSGwiJv9WpmVmpIfAzQrynUVM4pixgZC/e/018MEck+o9ZJ14YHKz1EWns
o1UceG/eD4KMKAAIQQkL86S2Y36+ltV1uMOSfVqU4VE+GD5Uc19qXNOROQo3
RVaiTTJuCR8OcbuBv1MlD+x/M9E2q80HIhtH51GFtfU8XrQ7Je5eIb20UtCR
zdZhgb3iox911d9CtYLzQvcHuGs5QZarreZ+7+1eONfhUnY5WT6bpM4PBdRK
Dd/oHmKCRQVU4E1tpJ4e8JUANSRetOuINKl9AAWaDhtCQfnRKixDNhCIwABI
qgR+dGJzn7/c0MLrcAdhO0YwBVUJTx9fmKPLWbQQL5FvHmTlJBNCha9k1KZs
iuqAEY+FA00nQAGXgWVDln/iUAMuvsZBdMjdmLfrAS0vYxarark5s6tGzZ41
E5tq+50MyxW/RlemkJR+o77QfE+AE28lTVGatJ9ws4RlAgvWXzIanIP051Qt
+ZyWh45T168kJY3nwPGg9XNLHESM+X9iVeahGq82STarrxjyIanKPaDDZaD3
geQ72cYxhiYglVC4wb06MRqb66GTlKeG06bC+5Ii+RHxcOqatNZbFvh9pr+U
OhG6ES2EXDv/wJFq8I6OtNuhzzO368+324X9SJwHFt3ul3kDhZjP/oH7zC+c
xl0S7ZKQI9NcmqDOxD1drNGF1PHmnIIjExnEz7x+v0HETd/D25649LWFLPDD
vMKpNK4PSmPsASe6IoV2nBUqFer60kfVk7jaubyy9e0mVPHIn7ZVD4h++7P9
oZVfATCQ6zA0QK30Ev2V57m37auy26ZiF81CvAmuBtIALxma/0osw0YRGiHG
JfrDQc5wqYC61RU/UF7DL3D9DxpnPAxJFJLHcyoC/Gwxkn8ce4vvpkWP+CDI
Lxm5S1GsO3hkNE7pdCCU9gdgkyX2Ulv7+yeI9CVa+7sSTh+F01BKgIWtBfOP
GF3wYuCzOOMdRHCkj7ehVjNQVaICjq6+zN5MccxUQ/GvYS/nClRUTzsK9+sn
gHre+mk8nnc4V3XIbCbsWKQVPWndo6H51ysM68exkMP+LMPBHUzflJoS4ozB
zWiV8zsgjYEmTiK18x25WszlS9ZOGhLEm4ogxydFlap4VZ9Fct4rh1b2/eO+
AZwZLbrtpH37Vrmo1urkMG5oWEjwYkoVDyg4MnwA1FMOiLrqL3DU57CEid8Q
nmidYIby0HFYhBEC9Ic4+TmkWvVKqn6Pm4zzpkK3rtH6sJMh+usAkHrwXyks
9y+le+DD/iCO+xN/Wvxgc+prePmWJrp3k1hAPqxz6kkEN0ke2Xen/WdLtQhW
nALrsP5fSmCnCcuk2X6qAPxTDMZXnMdUlmk5ZBhiKwnee6EpNNXZlH8MoopP
rghJoEA/VH/wt1EZUx+0WyR6wqalRTu+4Cds2GtU7EKDLkIW5uIJC+iSFzxV
mqPbjWgD/ePi8NrkboTpLSbXuEiZ/zo1aHahnouyK5OlxXb9CaGYLLnTKlCV
3tZ9RMbaMwdsNgHHPcdKksZ9/DxpjIY7SRFLUDj8y7Bh8/PsU+/AChcyDZI4
hWXGjy/97DinQnnVwthKZN40rYDnY+bPueBGYe+MgMY6ToIhJSfMmRyrBg4K
ibST5m9xZ3R2BDm8rUvGvPxyVbX0wTEzhARAxwkgDlwy7rmssWWS4LS2dlIB
GQXHb663UnDbOKmB7e7weqxjNi+ZYLfm8gjhJPcDjZ5JjOKJ8bMdlBvhCWVL
gd/YeXMCd8yMNNdL+XHAfcydlBIEILQAg4WPZOthYb5Rr2bxLzh4/z8gQ4xA
v5h7GWoME6jH73cR7jK9osCvKbWeKBJcZd2TeAyYzIYz068QAfMfb+Wiur69
nLHdrQASO50cr+Gz/xINE7lVFdeNs4FpQEiGJUWC7SkUmrqx12Hmn9VbCCB6
D5gizpmNUnNccAOLVuVjoTJnGHq4yNsmGABQStrbfapnJlepJCQBtHio9x3k
3LcFZySYHCDGDcLu6GTERtq6Cs0R/VtuPxVUxNsM6Gjv3HD23nCtkl+Rr/Jk
/JV8q/g5CLmE/jQC+v8lypMyN96X038TkdXWmA5IPqCrpLsUckMG6CgqQiUf
kk8IciaqeCvB4xJLa34tdSrmmf6Q1/ZqqGae8JEKlkS5NDvZBpnglR08d/1h
BJqcmejel0SUOEHx8cCCRgRR8vKk5HreZJh9I2Yv9CqJZTFhFUnYokl+SbfM
tw1mQ0wp2mjcpSG0BBWS0CPm7qDAlI1vsVIex3lvESHhQM05zh2aH2+Gc8zV
g89ImbbhapFMUHoyZq6KUBTzAvvzs43pt7So7zDzt5b7dLeRP0v5OpyaUZ57
TmftH0c+GAQPohAdTGMm0ydbM9JYcZ8gHTX3Zc/YsohQA2Ob/9jCA+Dj2206
IMWqbj1iNzTCZgm4VatVL9fFSLp3DNLZfzNzlixQAhaBe2Oj9n6v8Qj23A3C
YBqAstYfgkTeukdBG+w64ILwzuQ74Q4qmSLLt5aLNYV8q3lSb80VINo4k5Be
QzZGoVZsbvopADTgjPszirk3Q+3PkAKDwR9xv2xVy3tNonrtstIIdm9fWvEX
yfrGpkpzbjw+eJUB1wiVARfVoM0Unv00cvJaafR9h+tOElk/Wysmdf2VUei9
fb/yiRo8nh6UUjbPa3zJjxYDsA8+ZscP3kKhtNPp6oH09LRW7HIjmwKL6IoT
k+BQ4lQRM46+tv9aPdkgfupOB6XZbNdys2jf4eTi1JtNjpatilECgvt4c9aQ
aZlz2NIVZD86tmpI7n4polnMheVnx83Xg4+GB3h/ty8OV7Z+a0r9ILF2kyHz
UGLsOnhoggxpHy4vBU8+hSyXI58LodmT99EtqgZkMEsMXPLqi3ZuxEoT27CN
jENHGSthRNzNVN+j+PjbpYEtJ3bZudh4ZuIUeoZg42BgrdECVh2ud2BFpRZp
jqsVG1DOZEnVrpPFj/CFfHsIsvKkUnsexerYIMWwm0uf97Jy5gpE+mo66BRm
XlsLTiFawUpvdv4jrdUGmuNk11Nv9s/wcQTelG02cD1si8mGrO/bPIK3f766
VkLHQ8ntFmAZJ5KaEkWQDyQ97/WD1iSgtuytcT9ZXCzwRQXFSSnOMmFg7GM3
IuzDarVhR9rUjQw57kUIolZp9D+1ejMPvAMm1FKBV9CwFiuBsEI65xnZrqpc
h3sxMpMv6PoBBMMOFn/syN9qLNYr2tGDeOrn4RBRYB8BCNGDgyhxVs7i3oQY
AVg2i+1+DI8sALKBpwAW7LNM8u+0MimJrTovaBUTTJvG/A1cvItEgxZ2QtVY
5fgzU5bbc6vCDi8TifY5QGsKpblhQvTZv9Eax2MYgF3hR/M3xZwvPrGGrONG
/5UlnavJ+9yIcuTfriYcYOFresdJTxWS/+Tz+dGWeMyY/vmuadPr76vxrCEc
8c4Xtsd0WcOeh1nYTTuunzxilvZhuXI7BfbKtB+z5Zdyt7dMuo1lVl0HsLlq
oxpKNjbJnPnlbWftDAdYuQmF7MzQzBNEYkZ+8SYjSUz7egUv43rxUtSsZHbF
aObA3FTdaKdfOsNtw9R3k964Q6w2IWwnwL3BDWq9AKDEgZ8187XHhgiJd017
WyZHQ65q0r/iLHRT3LoWpnZ/+7uhNoeqTVrYPO+uEHX4TCGYg/7wP99fZoey
l+hmfJuK3P0KYuyHPKCd87wKTD+CveidQn4L+0ABrSVbZyDXaNUvwXDVR5/D
E1rZ8UPep+rHWLqSm4aLhfWOJCeyuOmRYBjYFwXUyX5v9ZTgmuXfwKCBEGdq
2N2q9IkOIghqEhd08QAI03OWExD/huhZLDhcPEhwnTqLwiEPFyWSqS6YAvVJ
Fjjkno9xh//edA5O0pFe6Os4aNTFxHjE2buqav8eeY3l3MZkYzPwtowqoXqO
h5HD5/Pua+ZAYFp74b7Mv7VJvjVL1O3KtGsT3gqDvVR/8LbMAdOZNyewzXDO
go2+oW8dA5xSyl/9/9ecjOvk+eM1xora6y/kL0T/cFsb2eQNa5KEFZpj3vMk
OJHlX3tpHPyuvohO+N+zMq2FdiH0yjD3vERMuFp4r+ETMUSfMKUEum1kFjBU
1q3tGCPEMDRKfshRkv8N6d/uP4ELduArbAH+hSr8D8wIVvFSZQvtp9gVzVcO
VhI5x6taa+QGcQfrnxyhXTRe2vp77rEB5J2ibe1F1l+xWoRqfW5g4cvnq2tv
7WUMUfN9R5vkCo4GF4g0tmMGYRNnOR1uQ63Z2Bl63qsVftg/V5MPkrvjbsNb
uMRoQlZ4rRk0Q6bQtUPa2aQuFPrXug8Ia3nPym7Qu+U4xo+taDvvznlsL0Ww
BaDj9lZhrmnaPxP+6FIg4XFboD9PYW0hxoYJpk5bUnxGTxPjpHTHE7riTT5Y
4piN+tmhJ09rmbDFk3S9MTLljqB3YX3QX4Mtj7lqUFP1FL1hFp2pYPPitGZG
WZnHZZdvdYRECwP3w3KaRdZdt4j1W0euoDp87U2GOC2BXoqLUW9nW/oGBABR
45IdxycZOJBsUdfAl8XUN5MwOezCQ6MJJVK+3B0sWxbRwwtQJypnYIR2UMzP
aZrbW7ck2QeU7Ee9U9xaGvCWI5yEOS0tKZG4ByUII+szmSFIcIWv2EcVaVog
UYAWKM4jC3ttmNrELzkaZ5okXRviiHa62grccAu6up/uLXP9mzQmSQqGU0gx
MBzgV2jLncMb8E3jLnziyOKsExdUAmnsyBCEv8Taa/V7NJkPiBsLYYlhFTwV
i4Hpt+uSvV3YF0nrBdVdF1nKzopzIJeJV2wB7FIUGjSGL649XF6GfIQ9kHrJ
npoNj+vIQeaqsGR0KfFY65wVZrnEVVLSLeBokC7l/yNfI+NCjq3n9Uz6gzh5
e1u/dcypwCyS7xFNe9+O5WSNnsR/zOWwXo4DiaLBCjexBL1WECGH4Fl/vr/N
ELcbp3yQOOdF1gyAsTO50Z1VUzY7Sh43vO8T8yzYr29t5Z6ot5IPuAxD3F54
ixse9Fa+gKjvdVcxs3v6COOHNP8H04OB0nFtJjxQjmW+jSzrTvl4qINAYI/9
JIR3QN3wJzLPD9JECYW1fxVA81DN1dSTvZY2C4Anig9WrtSo5bQQMJd7KMIH
TTudVMk9mCevjmHRun5WyGXNbW1V4W/vlqnlUB5xr370nhh2tgQppami4kVF
50DwV5bA9z+FoXT4mLSCIMHvStSb0PjEBxGVZrriBCdyS/KlThbrfpADMw/f
qQNHMnlKvChWN2wyF0rqCUAbjiFuRIDUAb/aRrydzn42+wVLje4M8dJOpUX2
PiW0RR1o41rieJBN11FEoMIhLkwRrmlyS8+qhhJ9ZzqUAQGj2oH2BIr0JUVr
9YX1po51mA1TYYcWCKSovJ8BFDEgenPm1LdcsVgFUIJCrr+bYaGRmmWHICPd
D+WE2K6csFhXL+nN/RsMl6BJnr7S4nvmTTjFcoomZu9J0UAfPxkvB4Cn9AsL
FOuhugjjmwfrCqimF7dNhwUUeoCzycb8yU2EcdIVBCM4uUO1p0IOb9iw9Jhg
lfPm6K07t1lbVMVQK+LIXg+MzWSZ/IYWJQvoNLKOAh2pHEX2+D8J3D3VE2fJ
jRROxqR70E6brfhIMT0+IkcDFJUeBl5ssGuXHrFkh65htHZak7lxOEFpYggM
roifvAAQ2q2zd+stbJZUYnWM47yQrvi0xR1orn4t+6gcVcxLkfVRev3j4kEL
/mOyN9fp6rDb9ps3Suiz8VjKbvD7ocr7SVcWim02Zb724TGmWHjePtJKlZAz
cjeO4sKVEZIBkeXYLDH9qk+lwCKJQ4XChCXHlJ/ebh39zMGIpfovDztYC3Ce
Em+F9v0Gs3fNWA2R3ink5qEtJ58ABQqIhyQff7YCIhc2t6hr4r8HPj6XYPu8
jdmYSAV3Q0rvBjvOOt8uy4OlXeKPfSuzxTBGrK8gPbBmiv8Tmrpzc8d+nqm5
NFzBh3xQvPGcNfg1OAyl29YSzLmqDlw40yVmXv3/3l7cHHQnQO1sWCQTC6w+
TDqXHOthje+WvoeHatB0PIsVQKto0ViuXzaTevnfkpFGg3gaR3ZgT7K1h/Lx
y+jx/ywUGmbYW4ZxgUhChayS8VSuzBu/ME7xCGi8nj6HF+fSGnXNhNcl600P
8XMpH7q98UDMcf9P8PDg7kxjV/1TkXTVOTCno49ogpTJYfM6ffejjMfT9dwg
GAnv00vuf+W4tuOCe46ilp0KPqjR0nQJ4HbpJqbjQv537IY/bpkDDLFCrUet
rvdi4w7v01axVWyeFwQbX/n8Cjoz8vN2714mnSFE0h0pcUtAQVFOfJBC80ql
0aGZUkpvEXmmgnTINEmFfRqCb8zgbQOf0HWqeb15QtAXxTd99eUp+N1ZnJFR
iVtOJXRrjuSrrljXJy/EoH/BoO9CjxzmbTHOn3JIkajgQUVD2/Kuf7tRXghR
EwNywELb/+s3vIKbrX8NDdbPJ+XCwOOnbmFimBe94B0/fMss+jvAkKsGpM36
z+L6wUcZ4szTSbqMWGcddJVf+bF/gkraAb2zQDNUoRiKncBq7S9bkG4XsE74
vaAz9FyVC3GLm8e73MIL3Bz+/8JfKoy41T6ho0ZmsOJJh4XCooykgm0B6ta5
Rtn2p7fZfsPi1s1NraQSgVSzIhLGfecARgzmP/k2BrkTEkp6mVkMqqxphrtv
JKQmbfr4ioNlzm9FfbSgR0nRqfNbJhxAfaukGgYbSOWeX15DcG88w1zikxrc
cRAi3IVZ1ez0ksmtjBHg/TlCF8Gogjw6tlL5bPe3emV9vpHlqRAwepk1BLpW
NALWM1nmLX+77IvRNEgvR2Evb2tlNJaDOBT4K3snCMcF7vyryC6Qbge+mmeO
n3hotipfPQfst62XXLYxnpy9bQqfDqaC8vvL8c/fmVX8e7V5wTt6kqXI4EU5
if2F1C6NqFtw1nlo/2zdkz4N7EI1jR5vnQgS1/jL6Ud2Ic2mBDNOAi1FpF4F
p6klbJONAbTsEtIRHqkXRTlLGF1sWFLdCSMSu8pqZaHf1bTMFkDZ/eFYrArB
xfJtH3EfP5cxHLgHASC9calgVci32LryRVsm4h3t8ubaXhKbQOvNLluGOnBS
eUOuyQd6cDlSvrBvY5ugjCIIZOIiOPebPEfEnhtWxZBTxAu5SFO84VLQxIHx
Dq22TN0sm9vbzLQWoFXr1G5aOu91NkB1KXaX5NRUN2sbRXw0Gk1splXYtj+1
RKnNNeJPM2vB5XfOMdW2FxBXCryl19xpXmvz+xgu1pSqeeDCzB+H5zjROpoq
UE8tYpgNGMlzuxnA02DGdxlhC5TMdYXG01xrUD4stcjO7LteA9f59Yo9eKVT
EY4tFZ+ciz8lFPEhwIUV+FHiCHNPmQ2qH/D2SjSXs/MIF/N2/9uwa7hTM9Wf
HtFoSGNA0fFIy7Q9uV1sDi6P/CW/uLu7OPTyk0wDLc78WOwM4ToobX7cj7fd
4jXhwjzL/upcqtzy9DQdZKuX8U+AUAyuGvRxBkwttS4iaRBWC/ZoIUkCyT0Q
XY5uY3zVbg0x84FmiPBlq17mL1zpaXE3rl7OKCCgifK78y132yFNNYie8m2Q
NCv68LeWanBqInruiOtAVdC2hTcyhcr8C1tb9QsUt25UzFqvuiXXgafHYcRv
NcfzfQIGDCZtBtOcRNEOJMlUhkGXwbWolkvzD3xxyjYqBSoJuuKD0ZAS0C2O
C9URs6BReflpTpRePYb96VpishukUd5Xt3kO8LKz4bV5c0afZE1ItNyimvgF
LO2Ryz8lMGS3pLtugkHlUd3yYGc7ErwDH47nTZUojftEvylic1CwOGu4P/Ra
cLSKBbl2AO+cv7yucng9npxakOxsNlEdSb6BW7p4ysiBrX4b5ZLzZUAVVjld
k10aDeY7NPJsLxG7q57pU+BHVbwNIUwpGP4qikPn6UKtu/U5aKylj2W9X/lw
qVoWu/tCab3ZrdSIAdaKdBqjSDLOFb0c8f3g6OkPovYjfyLqNncZV22zs7pM
ExowA387bmUJZcmWDZK/spPFOPpcEpt1Hkd/fqAlKhEiNKYB7/8TNEA4KsOj
QctWg38agCDqZz3c3ruZCUqfgC+wgXa9BjzD+5jkjy3/Er5NAJa8motsLFVK
pjyAzDd3nvn+colDgw67TCHQSmNxpA36M1OIWOYdjwSpQHwkoLQ8CJhMAEYr
wFybaJYewvfMHg6n2fvnHptbFQT8g462vxd/ZrkUweG0/N5vD4wyzA02omHp
DGk7zqyH3llVVCtovyb9t0v0EgWe6SfBHGtE8N1hG8UciUfIdKl3vGjfBbe9
ZR/NVwzySmAMx788PYydSOrIwDf0txGxGYeuMg4lsdz8FJ/vkBBGs82KiShX
Xqy781ohaPGcNnr96O2cCbZ6xzv3KnXiZ9ELrk5ehtrkbzcjsDyegGJPS2I5
XsaYdRlVYgXA5iUWJu63jW45KwCWx0K+zyJIT0l/jh6+GxkQrNAY4B/tHR5A
0zTO+iET8lbvtotUBWMQxQkScNCiZPBLeV3lXCFwEsynevXdR/22KjssUy5Z
ECdqHDkQptvuv40tSLqCMPfSjYBOkFCilDVt/WjI2d1+O5sdkt6/caohWi0y
Jj584mq84krWdqqi8b/zxK0c7+WbqpylDWWSb0AlfWPMdhprTnWHq7pfHqCI
9FXegNXG2hZubM0W4WSMppnQteorZAIC/6TzP8mCT74JkpnTC9iejgXbl4wa
ZhsKDve99DSWVVwTF30WtjBcNjw5GYSKLGmuHgYoknWe5GH02kWZOLz3tQ+B
d+/ZS4+k1E1iJ/Tn6kiylknAr1xZrsPd8dKf/yGUEkJQjioxTc3dX2AYZaq9
9qFotipDSeFFUcosr7aSJJT15u5vIk1xhrYnzxmNqMRrcxk5upMbfnsbOqNk
n0wA4nDrSDD2eKA7aI2GLIkDPkxPr2glbyf70AiTbhR/IVuMf3Cev1JzTj8M
OMjBS7HdQD4+wMNaKbibCPzEhQ6aOhSWKb1pMkHGl7jXSF5n0s3D0unqfTy1
oE+ISyOtn390OYHoPL+IEWwiybBkZUk4CoLF00td7N4ZraHuG9XlrIkKocMB
Kv+v0nIXEmdDUUPNG84aBs0Zt0HQVWqS4lKjFSNrZkbgTaH9OXxTRYzZdhM0
yR5v3iw5kit89r2rm6gqdUBAFmK6yy+UT4xvBCSif8OkHEOQEJRG9WjzrpfR
cd3CgQxvVk6KzW/643B6d7SKhQIwIDQ54Y/GE8nAwwlNtFNOu7bC2JmEXSgK
E26EivkJFnSiNOzcXHlDws1dFFh0h3o6+yADP6zs4TDfyaCRaW2A9Sx6DgVr
VxRj8NIKoDSslsrGOc7rxsoMDzV/AQD1u1XqB2ulRx7M8lDI0lvGMgG+Hr+n
ETDsGfRJx8IEMuzKCGptq/NrVzffQXVGFSf+iTpkCjUEjAnlK6eMXmPg0x18
9RZYV9qEHEGh0itmW/MS0wcPGxb3f+McOAlZHiffWjQgGsNus+UjkcrqI7hb
SdAX8VLLup9SG5mF5o730whDTx1N77RnUkoyLlqwqmkOgyVxP5CJocEVYHp1
dJngstv43im+MRRQ6iA5mZrOBzCpUwQIB2Kb3faeRN146YIO9XcKTmvZ5V1K
CUOOW9jHVNx7on0MNpvGyqx7AsQFl3sWL7PjLlIT06IEHQe3zBzUvbrthrlI
RswD307TlJo6ZFlTzess5UsPWGWvl57xoSgG3IOL06Lg6EDMSRpsvJY+/Jt/
VsPa0r7RJxFMlqjDTjeTHiuyU9Lv8e8ZFEY7vRctIGup/T/VtANbvTO6xLAO
dIj7MMuhjKmNIMJbkyBNat8Rnse2M+trNpUntl/XdSPKhtc2kArRFl7xP9aB
+EIHixBRctMm+xX6H7wUYUQgsjljOuyXdKCWnAVOvmfrrFTZY6Wvc076h0Ad
88MNTeDnhmywEY1PiVp7J16LSGFVdFkWZh6fnzxNwKH6xVwch4uBy/NcUe3A
nw9adOJvMSzlxvfVzGJ4oCg/PeyWILLuucdlGkpWVcMNCVtINmB7Ub7AO8Za
GQuriSOm93zGxlV0uhrvu3zFPCqxQoMdsdBLUFoRgccX7tj67bEdpJEwZe+8
tpA/nTTX08k4nsu5EYlN93FjpSeCjjknXlO33eN533h7CIrxGXImzNkh+bIt
iVcLBS1fKdL1phk8ItdvNlzqAn1qUcR24zeo1RsCt1NSQr/avlCtnaqHKslm
X6XftHuvsyeuhHhGksHlSxy7vPl2yeABBdSVONdcRrVbkThJzNCVD67Uj0sK
gH3XHKDf6CduqJeJRUYX2JtuBLhOehNhvhLFyJqBzQGagqH90YGPZynsJ2XY
y/Tw6XmsAuteVKXVwd3xFhXFhejI2p56BQpEI//jdykd0tt8TnYbJK69a9Go
+qMP1MfvnM+xDERSdQF31usxDY/F6Fy1KeOnWqibPaCEN0h63jgUh2VQFmX/
9MZfwYZJsEEu1XY3aLZXD6LR7rGnJtO95UCbuM2EGiuzX7bLuqc02i6SOfe/
kxoa3YP1Nld2QqOWGoKj43gK0tDREkXRihlb33KfHOFINPpTdjPKUKMc/nH9
fCTxF62TIXGeY7KaG4CiYb0kcBztxEVeDUMc7nSupxa0uQnVUGTk7Q9k7pt6
6U7cCcA0fsykmzP3er1zgvuPf8yUY0ANH3/c1tRd/3WzOzKEM7iwL3ec4nYH
xhZi/ZN+KZ9M7rPwlAl+W9jC7CEzMKZzKJzWLAFh442HFAGW89jEic3JyCar
m0XQ2wT4x0Xp6y0/lqMtiloM/tz32/FweZDSWu8wWDzfgepwIi02guMpGg0Q
7jfoqkI+CSpuBrW+vPPYQI/B0QrOQscc07cTO0tHcppY+eRYDs2/LsESHm3J
LSJs7WDXT5XWoxe5KzsfCORISzv0oqZbyvguqchGcyTtKiDVsIyUN+rxho0X
XIaowyiju75mBd0deh/VJkeyVSWxyAunvXLb8ExBQ3zmbGk2ElnG/b865J+f
q+Kc+C6qr2B/sDpP75PlNMZMAClcR0bdJRm0VgFHcumYhNMgYeq1ixSi4w+n
7UMKIM6XNf9ofcJ/8dTWUa5vX4TqFrCQyMLrRKYgKn9dC3OJxCElCnLr5JAs
4gAWlVxsowbvwAljRvWrConPdvk3EnKHEMNev0w2D4pvy41XAqT8JEXe6KvW
fk4S6kcXXx6meH11aDMWhP1Vg/gpyW+7uyRkH5qRrw46Dy2TOzAF77/8JZxr
5Pa+Fv2psHxYrjkO4Q8rnjLnLRvKOXZZ267uvBDVnz1K/TmwGc0AVdcvobM4
rWkzG7PsjzCrh2fCUT7KQKCIE8pcgowOSn0FTwSR0romTbRFbL1o02CyUHgg
bSsA1d6K4WtKiGmbiIple2xc3YaalEzy+65ULTS0UAssF1dPcJ/6qvDHELUR
MYWKFOnnygOmFjvFh+S3Qde+WrYlSKgN4xMo3gjKZ0KmdZBx3MfhAWp4fEB1
EBlaACxWTR6L51WaNidcYlTwBeuMNcCr62//s3O0ntTXMrD5Mb+qkxq1t2rd
rkaPxPTaBWoNiDWTpyj2UdnpnAZXypnd76RmIdPshzXcJ7Qw6yfy7xcwcEus
ozdk0TnmC0Lvqt2mskOu5lTimlMpiqDG+d2/NWLExTzCqQ3ljPd6Vm4CO8pY
UkvUM3/T6PgQaXYhQnprFcQJKswSa5p8rxmUTcc+Ea33a0rHRwJ+2zFWjdh1
ShH2faFfUmB0c6M0IRy2ViVa+N3VONX3E8+hhl2CIzjE/GJw9LFtgju5JJCv
JKwZBH2lfAarVEn30fjZ2JTGn9kziTLi9nPFMmaRQk4n7Hh2h16idBXwlgnK
IystGBXqvl9S5rxBJX4tvheD2G3GRF72qhUlROgkhNiCsY9AIP4RkrQlnuaG
Lz/A97zCyqzYR8x6VjzVMDHMrzEDmYXj8Pe7LPNDFwHDSMuGhVE9g22e8+7c
DO9Ot0C/kmd6XUyvDNi9bfB1A2I8Ah0cvnV2ElSK32xDW8hVHheOkeloQSaN
Dn/CmhhtwvNltkN2qhEWNDdtB8jYt7pEJoG/k5Pk76dRlP8A2AJG0sHFOEin
0AJSZR7f41tRyjFQ+2NlwzQSxrJeIRWBD2fpiCObv/J/ofDikQ+O4W2sVArO
UQwwyXxvMM+qiKTVcCd/qRP7SMIwR7ljDu90YTRzzhsaoLWXqNEcZtDG9xYz
BWjv/BJLo/sa4tAcCui6xo7qnBv8Ef81FtrAiz6QE/wcBTp1YGbaZN/nMEqx
7L+bySJ+lnvWjwku64yCL196RruG4uytnqCOZubiJQhhwUCJ7YtCAJsU28YB
Y+rXQKhDT6ksyvm77d7yMebAQQbpFCPyCbZMfG7W9SqEbjgTW1O9P+Mt5Mvx
GWETSv9q+86y/3I3odYMzgMC5kFM7ndPP+H+uzlfARGkgl7QGK0GezrgEbvr
7EoUklprfDE81sEHf0GINl/nm0/JTnDtrjWYNoMWhrjJK1dBa2+seMfeNpbG
SaNamcp+F7fTxM1I0xdkLsZK9KaOQDf1A+/ppTBFk7D44W49A8ikiSfQa8he
NFgRiC3WnIdiuwUIqwGDBCNJZRphgfX7r8thUEVKF0z6g6yY7BP002Qt3qFt
0VQ/q0BYK1UxaP5ZDdsEOaHFi9G0vkYmITFA9UStIJrke+3K0DvYCE9mTmY8
rafc0johT40wzix2F/MF1g/33b/3jEv3u+lKdozgKKXzwnxy/drc87eRxsM6
iaGeZrd41JOYEpKikQT1+WXXNhJExN/xsyv/IGojRxfIE3ZVXZKIXKvXMK8Z
H9pxJEOa+XcAJeeP1rYgcxBXTcDiQSHAzK5hKG9OBlukBOcRlOZ9+TzQiJAQ
zTtM7nG0tCBhTx0Nx+auszPuS2jSjSGxdcq1l/eoDRfoePS+R9FhtN++RgT+
TQso+sZgi45OUw3W7xQkzc/Kn6Ues6vW/1aRX53xh3eAqpdM6L0oNWazXiao
K3cS5WvIewYCDn9aUADi09sneNHwDx+9FEcaZBNQeymcZtRPZyioYd4BrbbJ
S41qM/fXnpG46MRPAkIHjIGer+OYP7kWD8ldYou4iLdGYNIFZOjYiZCdl34x
1iwvNWsnkym5kJEtoupPZJl0dr47LNY2s2BSj68eAsuIJ/mWKfANt+7MXlbY
8rROiQ8ysq9ho5iCHBMJdNpdZImucLNNZVR8vGDrUAdNGs5UBeWuMKMaqXtP
4cdVzxNt/h6EiHBzjEL1ZdsqLIT+kvUlKfDlih2/rge/O5CulD1WVxxRNcS7
VViiezbWLyaZk743wEl2pP5dQpN/8stvQ6o+s0EbbKgd2VUY8EbhwsIvOMQF
F6Hw+UpTtekjNSx8YAWcvbz80TjFYITQAhffJ3HkhBUIaHqV/Cz4a2uGl+v3
JBU0qVCi6dWTlLsIxvcPkzT9ZBMTYouRKDvlej8UW+sarQlwWoJmSFwW8/0o
tvYrtCwHbDZOiGTWxer4b/6/TrdD47CmaB7+699Uh0PFFl7ZBeeAdeRGLDQw
53FAiJpuJYtqtUQU4z1HwCGJKprETq1va8Q+Sluwh4e6smwl+htrsIlqbSRy
4YyKei1VMzpjb9K72noYapIY+r0ypS919Uf9+fHyct9Cb1Q1e72IBoACbdHu
ZBliftz18xJay+gNhvcyqbz5u3UVrM3wk3JdWgbehRSPZnbPrmfmNOu+v18w
3PCA5OsvfERAi5+aNnHtAVGOHuVmK0ZNM8t6xW9iWgsKB2sFSPD1hlFrsPcs
wZSrCl1BcXfsfwfs3L82KYGHtYgz+pZJglApYFcUYxqywdSCjYPk3YLJQRkl
Bw8M+yFLSwOOem5n39Pk6xhKCqrneb5nYsVE3q/vjRJ4duyj1YiL5vrdHboA
bK2eO4On6dkloHfp1G2RG4UWo1fbhAeVYyX4iG/JRRB7rtTZwSpCfCqSJlYK
usnPaGHPIGbfNa+qK9MfvT5HOEcdqdVK6yqHFU96d1sFVxsK9j6l4uqE71Ba
t4EeIRLUm62k2OnpMSYQSDOTYE8vOtTLALhl6l2LeBX+JqWvCrzUHxTZQeyB
+D1GllCNksKqMLigZM3T4Eyp1xa7ooiSIgybVLDxXlFNYhYuC0QcR+b+6hQX
3geGg6E+Kyi4L6+c7rLGmHTnPTu4QDtDLyjgq+Kp7ogjhXXCerIPSfUkbsN3
f3x6scp9rt3lYhwmkFPDGUjVlJuBHXUIYR2rlJglaq6eeRyLyqVxSclNweR7
Eqxf894BwQkWd8PE70wGwLrEcle+NSFnYemAO1hi964NkGZugC7OeqxdEfDc
QJ6khCKQihdL3T0XeD8rRDj0CNeDRNvU1ulgYY/B1hRJSQTvx0HcvUFhLKUC
LcJnEDKJAI+ms4ppOn8LryKe8Rc3dK9XLsLEwW/2H5Z+hXGv1gQa49mPkwVJ
MfYxI3HgEtCkTJqTDI5XyrIrAS8Cag9hFe4zQJXW6+xW3BObMFEZT1qaUUQe
WQ9jKk3B/GcEQ7r5PH4uBOrQyUz6C+FS23WjD5ChRlOOtp6udtdPPqzfhlOD
V9sBJryR/3KlNr5nOdi+X9AWoQU8DIR1E2bQLlXpplFyrGgKoABpLsFOykmb
Q61576N8p3HFGga0JC6y42Dggd+p5uppzN1ppYxKTad4Hz46N5/edWnJX2Q0
schzvKw8M4ajrph5MhUfbDxF/O/tnGaqQh4OpYkZYDSbW/jOP4ZAPAx4SciN
ROCLym4GAKOsA/WVKe2PEVrODbFyZm1pffDacHOiQQ8Z2vaxewqDhv9IPAVb
8r1x5aR0sUG5y14jFYQzMjscpRhyhnCjAT7lMT7tEOUDxoEZ63nhZv8uwYmy
1j0Ji8rJOqRadT3KJtSPgkfrzfn0UuWfjqEJpwLJfr7jbsqEZs5SNDNvNnaj
MkzvE+QZz+T17CZI2olo9o1eiD/SoIYKOrh/ratF8vzN6PHfpmrtxqNc61rD
Tk/zMvOB2J5CiiNSr/VktbD5BOGm6/QE2cUqS6RgAzb7YFks8TL85K+q3UBq
tl4XWXSG3rdmedML60PvzEbjMwZZfs9zqqexX8ICv+upXJwNXCL+5RW7W2kP
g0kvOratGPI2sm0/ozlhmNb/PPKPdhIqjE7GkQ+amVCYi6DuzzgF5vOBrUbk
2a/BlN5tpMHSMnwmpQsT00Q18chnMaXGdxvN5XEBVg0hTr6ZJdJA4fVJfVbV
95E8ZYpXLMtpMSw1LUnpx765Vvyo+D07lGOaPKh/yhH7JuNQ4n6WPkxbrKne
xj2DcSHTMD73nISiqcj7sUg8Ekq7ctOXlQu0Xsah549QPf7pyx37Qub2QgEQ
7KCEbdHTUzKFLQjXMp51f3vavQpWv6oSyyXQIL4qetVxxyiG742cwZbaD0Jh
5b2OCzcym/MY0L5qNt7EW0PO8+Syvai49DO8lN46wJJ9H23rmHCUND9Ju+Pw
tp74J1QmFzVAgeNMVmxpkgz8wmqgh/VHoVqTcjuro7CCWgucnoU9sAOx9LG3
ohOHWbBKe2WWHfBk3+tP34mj93stPN6XbxeYt/G/u4zBuz69VU84mw+A23c7
k5wx6TjKckBFe0y0R1GypP+9Ql1mLco/yHWMm/U+oNRIL0HERh0hmfeV2xCv
ebiDr+BVqFVC4V93+4a8n2das0VBTQEkpNgX3Uv596tvygCdE6n8q3LdT5ru
0pUYGjKYMnGLDolVBNIqaxI87iNopvLqrWyazkCGaVJ0X76XBMVqnlHIo7Ni
iJaZgfIM+hZ6mKLhiFJ/4XORV8lNH2YEwyAvCCCd1GBJvV1N94C4V6uLfq11
+32kpZqJnSaOop1IoKphhcYKJVtntoNNYf49D/dNfG7Dbu8fVdxeR9aq3mTU
Qywni49FRIB5ou8XnHu4iEnQfUTikyXQA0POov7bQ1PBmv+PqQWeNWuwxg+q
5wfx4XdwZwFO9rGQeeIhnu0WnmcZcWdScgJn+FleF7pLWAmvLv11YuRpJ1zM
wxGy9TQ/0YbOsHiVj42D/W2diBFcjNQTo/TMWiqYiFkzTdU3yQcGxC55FyH2
0spKMmr7JslvTCF27e74bAVKQj91kCNxq9XF3T+af5yS//Oe1kmd5siFuyvE
BO7gx8gam1FUj7Og2iP1zQnSbwldgIKbXuoERLP2tIwsB4FMnQSW8lse3TqS
nYd7BBonaK1UYHtgtQOoY3gZX93glB26pzlZPf3mVuFP/spFJKmALbPo34u7
bFoPglCzQJNONSYSL3q3wS2Qnx6hICndp3PG4oUs5Xm7VY6Xl76gMPV421SN
DavvHBCBkkDNGQlw1avfaHGrlwkbQSAOehQgd8GXe3+M3nmmv/99m2/p864a
lxU9GXouFdmHV3eO/FpS/NE2ogMe6NQAAZro4WRNoxuHOSO9stpAH+Ekm9sJ
rCXDpVkcRXK2tpZC29VyzRbBRErsMPrr0F8wWYV6qg/OYUMjli48jpQVpMaP
JMHYRyjuLOTlr4ZgLcRDQgwGlIzikEiO334yvZw/iQLr9MVQo0osVKOA+f6N
aRKTOnIGEoQ39KWwTSmTVMfUlGjAArHI1y5/0nOO3UHvKncKFE1PtwtED3cV
gnXeJwev6rQ+vGu3nyPfM/PekilBa6TtIdGUk08FZvHYGUf+zETDKUnfqVF9
INRTfnIluv9mBCObBVCjL0rE7X1ZnmIQgF9iV5clwjAxjLgkQwKjMWBWFxJ0
vXmtnmoRjbA5lMpn4ita1ZQuGZrg9IcVW+Wf0tTKH69q5B1QTUqL6Ohf6KW5
5EN5mol308vu7UHiNX6TsarPdNfJ0BDlCsEhj7Abnvqgd5bKI29LNM8RIUpN
WiSS9zgtxFkLOjCoMq87bNSOWn2oiUjywCZm9HbZph+kJlmxmcWbMRj3pP6w
pUopOVSLRy7QLxFBkf4wmmJt++rIR3bIOCh4/7pY3tqneGHo9sdi66EHbmBX
axsOwQOb0buYskAGWt9utO7FAcgOI8n/kVOhzH7gEzjh0k+dZaxknF4h1C3Y
AEkKrSlQa+xdP/iMosEEAKQDtLtVIq4Axu9oLkANm/gfrAe3X/8MazIu2+xW
NCwi342yLaYl0fbj5txqpZP+CRum1DKrBp/rmYVALEaLdY9m0FuMxm89Ic+Y
JuH11E/rT88cSq/vJCfO+t+k4ffV97cBrjE9cG4GjxOtJVhnBqbiwqWWQzWS
r+3I/wwSvdTW4+gqcX/9vbdGrkvii1F1+1jI4TrLmjZ/PwicO4jEGY35FkB/
u0DCv054DEsN0l9fo0S/FwapTac1U8XbBc5EBpsu0nAv9fh6DSTtbOQ4JcEp
oE+ppPwg32JDanP4xZUXWfLlIRmBqPbCigXmJSi5yjElDNfvO24V/RGlVHVO
yYLa8TlrRpSyXmAM/9LC1bYfgDRUS8Vkb/GxUA2Hby3JMzuIsNhZXwK77/QV
lH+3PLq/OxwGalnw2VupYpA2LoRZ6XooMqpKoLJt6PTEi5KYzIs8pa2HIIHI
76gGE4M7kf22axWwqV7tvG9lemyo3wR4XF+24aTA3ozahAWDNDaieZUJ5T7F
2f1cnjx5843b0TIxnoer7n8/ND6QlJ+icFWDzfOTr+v1UNb8eQoUB0YUmEJk
YgMq2W61KIgEe9950YVIXtGcpdr+OIBwOrDzeTJVEmBz4tI/SRad1ukzFCq+
bTAZgeUS67ubZVy657BJ7VK5EchIrfyH+trsX3hDo/FFCMsMHyRE1RMAfuzE
+RLiP1xQ7bNuoCCMOnJtyJ0gGl7gqjM8y00vrCFGDWRlq2Q7w213wb8vPZC+
byxSyp/0o0madkH1pTW7ZJeeOTdFlsjWhPRDajK9C5W1U31Lg+HmGLyAtrV1
8S66e/WBueU4EZ8YYLaLJyIqNNGsRCLT10FMHq7Dm9WWTDC5DqI834KuANel
ZEQuaeiPSigf2YuksthtZF8v/3C6Q9fYr9XtaI4zP8ymdh2ak9e3bjCJDlRU
oB9bhhK1dHlq8BjRCB/7HrZIft+c2YKHX9MNBoOk7ZyDgLbBiDNYV+WX76j3
8bRGhtnfgzIJ6jUJOkU1FS38a+hQwUAQFm1funXQQkqQpO9jCD22bXkFo9gg
DT+m2oJseTwD3JCI4Ys2NuMqGMAw/3WeKsRJrD7P5hfdQRcWGkkpFnFx0EOM
haol80sia83aTovVh78jPk3oc6I1DRm3quKRHjDoZicNL2rjuUDXawdg0AW9
iZmRujPnHfGC2LxnGH0hWVHSr5cGCjvTrRRNxHAL3VN0r5hQfVsTrS27LJmt
cINN0b4ABiRqIwwaBBOOyKPM9L9wvdaINq1xbmgZ4E++1z3i5/hzF7P86FPo
5bk2U5P2QkKzRJlU5oSBXUHzDtUDgv/J/TRkYch0onzoSvUDOxsomVP6cnrB
4RBwogohVMqNEHXXSRrEc5q3hrP5ZbUvy42arKPjyBpiSu9e+N+9aBEpVJON
jYLj8QJE4fiI6VxyJPzv1lmZNyF2MWJuLNuE2xCnN4087C7AJeS5jIygKOqU
zHJNR4VH7ohdjZQ8hHgmdgV1QqGuAyh9Sxmn8EB9Y7aZwR7hcixJ4ovdo/ak
K3a8Qp/5zn5uUjDwQDrdAzcj8k+2i6sSrmVy3hpqKpZJoo1F38oZ8Jw7OJ56
PibA7az/vBvjxBJj8G0QBms6QCAT2uJ1wTPPeMaSCDk9bay9sLGP9FiOQuvH
Hl0vyAGSDbhthGqb8BA4wPR5S2xyCeWLNfTnhWzy1f1xefAUnjk3KT+jqpCJ
0Jfl1r7hwFaBHpLYntDzWSffpkA4ZFWEAQZJhQT0rQBBG3vAQN2hw7pKLx+X
68CDhypiAQnV6CceviCeyfj0Xx2qq5rfGdVb/5IE/CZ8dPAFy399hG98Z2+U
zIdD53kUdiwZU5QK83PnPOunWVR9epzLaxxVs/78j4oxhNpxpaaVSgXqBdO2
FpLnv0oYEhA7NjpYvPzJ9ekFBE2PX/sOlmLVIoJJy/+826XBPFVtOR3ObfhF
LUq1LRhQavfXVX/znlGpb8on3VvwGHkc6OXIWquFgjNontGZB6+gM9PVpIXv
txok2OeftQX6M4vIo3T0U/bg4eh7VlRbs2i012kb3Irgl7+/wcUtaC3gd1wo
RX6aPmBp9+eN8MWOvRBOgvJeLqVYRdv3juX7dKZ+yO7lLGZpInoO9lk3usNr
3QEaf96xET0F21PngMr7CZZrDQ9TcNJqdX3xdG8yU65rW/Wnx4gdzGZs8vQH
La48yG9JrnXHJ3TwjvR7ioH+Q9YJG8a+3iZwY8CoBrMHZg1QIy887jieQHOO
1qp/ReFs74m3c3CF5vsD56voM8kvbCndHmRn6j5YmSzHu9MTVkvCHBlGPrmn
0Zzq8U71VKLsnrMNcBQBy7knJQ9ygzTXijJOiKZcbQEF9Hc/FmtHF/G7W1jb
0rtQ5L1vigM6nBTAVaTMdMxJjiHhGOB5KM2nfEXhdqEaPCaQKTLCAWTJ+o7R
Tk6czeyd1IOM0VEnY/kmxFS/NQm162BkhxAyxv9LbNN6tT/bsv6UPwYmosFG
W26vwGlr5ORtAaeX2WWGa85anXYfgjnZT57dwW9G64BneTXq0h7f4KFPcdH9
XkqNiwYjW9gI8Zqg7ydl3X/DDbiKOtb9tmuBKsB5JdF2EFIqzVJUplUZslF8
Ic1sF6KZpzlnNYVjflIxlimECe+GCMDhBek7aMSx8fepsgVBk/HUuu296nJt
24WJdDPcPTU04zvca7Zb3s3U/e95B3xeHmpKcck7XCBpOxul7JITzDN2oX/O
UoLu8cAigC/Kp0R3XMN8t+Z+Y++Eazd2qmUsipsuRRexfAe4T3NlUhCr5feo
xUBknFMQwzT/VCkmMP8dj5CYMcqvK3twomC8MezArqtuTzSEqL4CeAjLNhJX
3QyTC4Kwh37kkfdzOrISeS8b/CehZbeKx6T4bzzQhuAkNLdZWmyr23Gta6g1
Dl+Xn5cGoAJGk+sdo5GIuboLbSleA3dihNfpcWhDVnEcBvikYo3U5ZJWnWYH
YdFv2nSnuDEMlMmLX8gbF0AXhzEGureALHtdohTX+oKhqkYyDqWez1ykf/Vv
c6q38UHIVkpn1KHaTlK+xyAeJkmHB8RiGM55sz2GZXJ7Rnyby0TCVpQiXggc
WhqbyeDarArglfdPn0U9LxRHqTt97C+UAGFy0YJZxgerP6eU6Hh8nv9v+Ph3
gwHC9UGlNzJAtnopYHiQeQ9fyf2cFwT9RfmHjs6SBSDekTo/reJNC6/eRCdK
EWXFHtbxBWHnhQ2fz88KI8ULgmkiPFRkgyGwoa8ybVc61CI8H5F/lke3Axgr
2noJL0GQ3AKF9zZhXDhlY5XSXT8uxiRIumjZGn7skmHWlcWnndeDzhwn1slH
5e8+lfVPYqNRCNTmHg0qB6wH+EpjHFqVzzSaqxfuuuYff9V+wxNutaiQFI8O
5+UyUN/zOQ5CqKui/2KbV2OwFSNRFfVs2qSCl8BPzEtiuR9A/1xpUX79QiVw
kcFCWXbQvew0Q98TYmfBz1QCGkVIib7xUNJpR6e0cItnPDjAr7l3JZ9BWFA4
jIZ8tO9zKJj+Ol4V3A0LZ60mGEN1hzfpb07vh1fpQmA7wYkbm+M3yaWJ1dDw
ecEch8XjqsEUjmlhZurHPmoOjP9dhgoLPNK96I517k+2kgXoum+MUESmaEqm
klb1tSix8sZ9YwF5piQNLIrsHePtxzebPrtZD+MtT7GKzKt1uP8Odg5kAyX7
VMEh8d5kDVThG731iaEFNL1Dd0ecwuf0SXhxPmFH86m24MyJVnGTWVwHC+3o
ZS31vA2+rBSz7XGUXkLcs9rGG2esrQb+V78RykoFM97b0hEgbkORh+Fnh05G
s5oh0xjSNuJ9yf6wpTSQMSLkVxnvU+2GWHTa8YaVo4/dpNyxuWGM7mGXMCrz
WJ70KhaanPUW5oEo4wkr+XUtlWnDg9q09WHsq4ipfl9YBu3CZ0tcFAH6dYHt
O6TLI5Pk8nZRuF9LIkLocEWPZKqhjPMy2hITVV02HaHSUyLoz6lDb80B8dHN
71j1AXeXm179IcKTPk50FuTuEPyxDhaB5JG7uuaYd2mXhKcTOAAYDEoxI/yR
BLOqof99YPNDN+4hoWfobnAm7O9DtvhaX4qqRNQBF4EKv22ZBDeLDQIgydlR
cZhwS+wE4AA5fqQ+/LYj8IlJBcJvWIO1MrmIbWulB9LBOwz4D8DCQQCdZ/MG
9yPzm3RdELfZX6FcZ9Hp/IsAXzXkZET9ZaxvFSTxNKW3POaRkawA7hQsHgJ6
Mvkf2EzdAKna6T7m4ZyN7scw1E8IQOegJyWzF+B06fqyEWfJHcNsZ73N7zj8
ziO13lrl92nWxRX6yieWiVyJlAyV2dDrasMa49jx/Wife4jr3vhSC67Hnb/f
aSCCBx21XDI5GDlw1BfBATGH/t1hKh+ZVYfT/2/suRQMKQJgEKx9gnYQtGsY
ri0eM8GnORpaaT9mbsRRkUL3jmji4cHXt0sSx5iVpUO3pEm8Fq6mWhik0/eR
OIJvQ/ygaYOqnJHOibHRBS9LpA3TDsUjEp2jlcTwLZL/W/Qy+WWulTq01etE
kzssTTf59L8pa4SO0TdTVsLQ+kLY9CaBThuKLTsYj4sKlvpcEswaF67bddNv
cMhfFTHfd+ceNb8+F39Naet5UhPA/Wc09u2LZIviMBoBKs3wW1O6qO7j4U1l
tAllj+7iioaMFd8H4uHeLtePS4xuk7JnzGvJkCLaaAUJQXATdwK0ZboWuZlq
kXYFw4XKhB+ufUzuEHDdE1PqzoUs/2MTk63QQ8goAZ2gyZCJeUx09CZHjG48
/3QZWUFvlzmaNqK7/cOkcVGTu3A9yLDVcW26cshZtyMETMpjdEt23iLsibLR
/U/75Op577Z1gj/TPFmokuvbWXCDiVoO0G36fQK9b/tea3VnkIQpq3h15Lt5
ssOtU6LXg/9yuZ3W7t1aeNm7V+DEFVeupgZZYH3SLFJQDS/lTLRizyobgGOs
151Yzlxkq4qeQDB1VAUr0K6VPS8YC2vmOasRTWsDoDFkZ7Sh0BCLe8iixi88
J4zvtQBHfPrxQa0rvOYIl/uyUt6oNB2woLrkWnwUm5JPireXlNBwvPHiB2hB
mTRNhqwZPeO3mSeASqnmXk/N8WjY5HQYt9j+8IiDa2a00y0YI0U+teK1l6Mf
9uC6H74IPi/0gvrjRIfW4EY+nEhaLTK7hyRFKbzCzmlSEMGvXYGrNasT8UK7
T3WbXFeLLVuqBDqzMR6y4Rl33wEhx4vzkmhLku6YdP/irBOSOWDFodNXKYn+
ehrss+yygeaRYCAv4aLCUondVVpL4UbdfcmsfTCSAoAdAoAuX496X2HvN65g
4pbDpL1ARP/DHxyLhE8L+qgC1PI3ID3LaleuV+jvo9VnKXjTHEW2jFb1huUG
A8nWpwjZ9b0/VrCHhJH0zGGXea42ajYAQpy4gNV7Rhum6bdf2hkpNi9QUSBT
RygO4zS6/PX2lXQbupeq+yQYDbg7EdEtd+JT0SVP7BxLyMstUYpRcG1ME2IG
PHOv5AtmsD6JhMpg0YY2Y2ycp7ZhYWTzFH0O5IUzTjUKO1eR8+C/FdW5fIRo
U7937nXCOTvkds5oRY5BcNDCO5Gj6zDdGRSyeVMxzFu2vBSZvjQmCUEFvdZE
DkiEOAvTb7bLPWNC7R9B1fYmnZvpAUikuFdfGhoahuq0M/JoQa9HTl0ttaCd
m77tzcoANNc4YdRkCi1mA/YgvDmha8pngKabSb/IghRS6LXLrSQso9/E732+
dm9RjNKk7u2G5vKQaYWcw+chvoJChr2G/uSEBWd0RVdTe2bq+ODwWFMo3hSc
KMN93pHRpdSK5aebKAchnhjIPgKedTcOLgYjk2+n+kmAyiMc2SMGnSMsMgSS
zj35cPaKIJPzuqOMwcY1ledfWzX03BSrDQH5iSdauqDEPz5qE91eNeUGpR8U
e8wYsOX+9+5GStY49MDO//MtqKnNINqh5JT7AdarwhKaaydPkRF1puVowooZ
4wT2+lDfMAm6C+pM0wnQJnNAv0PGomZhYgzvP+ERw4nztj/OtT68+iUjdj+h
uc1kRNqAsW3VmRU5Ohbjg4ZpLI5VJox0iPrj7f3h9U8sh2UC+Yhw+yqJBFVU
DlaXw5O7weItuzzxTmur7kTZmu/WqK1ggBAK7IztNyzQFahrxBh9hxZGdmQ8
pHWCI0UDt1AKVDkjkXuwq9MuxDCUAISt8CZ3wPtWW/MbHqWuWkfN5dmPNQP8
Ymi163Q/bio9sV03iTyJ7OycJiASqMOqEO2Yha0+ZAk0iqJSl4irxuljj/k0
pN3DKkcPnlgbfH/n3jgwCu7BzNIipoZZQ+vz2Bs8vdpGSHTpcyw7oM/ONB6p
PX3xANd8/v0hOn2J343Zk8VFOkJ6Yh2KCErpUgkX3fYhbLCOyB6mxuegB1Kk
P8g+fZ2D/YO3v3SmW+W4bV694l40MBkNM4mF/asY3L2OcrW8U7Y7zZwAWDe5
5aEQxcecSqV/O1+O0g71NO4IjFgNJceiBvUZcGHrBKSioeXRg820Kq/RLVJ4
d8nUh+XHA5NnXVco3DvCv8EFAVhav1auyphXY6ocFWaceFLLNgha9VQ2NHbY
yYvfMuOyVX3J0MsJzT6/H07X/KiCvNHZhEmE5OAhSjsDHYKTH77kuhILH/3N
xM60GuHZr1HEthb90VqrR8Rj4Zb/ExQYeHUMcOf9nZVYJpofjOThgosbL9tD
A12ruI/vSqFFNnUzTouNFxasKIAloyPdg5YLu9Y7dPFW+Ijokxj5RcF+IMh4
pIIZouLu0sccwCTqzhqZx+pBYP1zDX4dg0eP/Em5/wVyFCYyQL3JWVBhtL5c
QGfN/6Zh4H+gzmOx00NnYKNguNYGSYIWqeMp6Qfy4/0My4Oxe2H5d1CzVXyF
GgSOvs6L7pm8XjJdu59kJzUcjVzPya06wlURaWJnYgRgrnt7jrDUzDz4lJHc
sSzP3ESfk4zVMfJP54ydTWQ18YrGnjZtXVdG9UlAyztXRoPorBbNEXZZehqY
rXWirC7o3//1ezXY4TrL+ypwEw1THBjQl9D5UPgG+D7h/WwNs/K1BpxOHlxe
2/cUfTBP2ALbKgRi2GXQmmpRYqBJJGKRXgXgqPlr9LibM6Gc02bktqreEJMK
7o6eq0Q9oLxwZ0OG7Z/Gs+KysWpBAg65MTya6FYt6mxOh3+wMG2Jp0bYLR3X
aTQNH/PaTxyB+SVr0Jf7CgNC5saI1/YVuwZ+PgSKdw+n49ja7PccucN5t2dT
XK6qoyuAFQWGiiRd8c5XspXAkKNaZUiZ913YjWndapQrsva+cm5fuezLG3iI
e7DGrVPbYevbm7YUG4WDjlnXDhj8yur4UjQsLymKa12CigvqzncHxdKSHjko
a1EUUhTkWaPkH/aoDV5EAeTzZEJ17SG5buT0V4lUUMLUEweaFRv4BMRqyhes
ZFbUxaBhIhlrI1VdEY905hVzj6UYQGl9rJS5CMaEp9XS/1B7p4qAMajBpEOI
qtpWtDijC1m8k8UU+fjW8kCnnRwZulSkMOBt9xc49LrRmvQxSoY7ksuDN5Vg
muGk78HL2h5FL7nywQxC/WnBweV2uIpEhr4hZqItVwSTxuqhxpJk92Xiv6MD
hATo5Pirllq3NSlQAmkWhsMBYpLnmzzY86kUVIhZV8EMwFu/wPvXCpES2m4Z
WSRDYJlu/4B/ex5KXf0wNqf4v/wM3KU6FzfyFnO3+boyJoIiqw1mY/Jmgvfq
0xgPGRNWvwZBcdinKeQd7lyCaEJRrL+cVlLiNEVF48y4VjWlxo0dO46Zqj8u
xpyG879wDavSLMAqzR6M86dEzVD8TYi5IXOV5x+hoIuyziTeqkyBkDfq37uW
lnOQBCtsGfTVuZyhmlzKaOMv1VwgdZqGfk284cfrl1lK+GAOVb0F/obfkJAd
pnT5ujGglWCcjdLegAPfuUzU5fjERsntcXuWFrBxH/yTNC4L0GG+PYQhT5P6
Y0duAwTWhnK3/WcYeRxgREe1aOw6FAHIW09d99N+VVg61tCjdTpf9mcI8iyr
DtS9PaMFixPJAxXBQWhbDaNm3TNCbX7dYs4OZBgCBe/ak2nrJ0WrtI6a7N8V
AhPfSQ5vUyh7MLWMfEjslYCRr6dK/NBdvPdYqEY8RhP3AwuDvjMiwb8n6SKF
EtI2fG/QMQY2WNSgfuLrHbxjHGpW1j9DEf5emNqY2OmEdiGhEN51otCP3SlT
fQLBC8dmxlDYgFxBe9/TeoIJ2qHX0XneHRfUKo3L+Ybgzt9Rn7SFq9c4TEgR
2B8n+PbBsJTEhDmhsQmFN+YO23qJvNf2wYDcXhhzzCJ7FjPLissiwsSRZ0U4
vV3UjQwmkwEGCGfF3IZeRrK1vTmQvCkhXumA9Qk/8pE+LB7xrSxjw1IiL800
80XYZmc/rWrXB2GQTkjiQ20W4msxExOgvqojaH6/P3Rk5mNzKew84vwTO6yU
hdWGXUVjpGY1MU9fyQIfQbwFmPHRfCpHOkWZ4LkvFzHNpzk7tFd+gJ8K8Yp2
EZtnj919JIVeEs5JUglns54xTrSAQqIEqD+psDMlSO0FQVd0A0B9fQd2W67V
kKX8J/CQuEHX555Y64uHqaiwZPOXJQaE2C/39++dk1MANGEKtRUaq7F5sKO6
Dg1fJpiIiktoGup2FG9KqmCbNrnz0o+gdsvfl3bge3KEQXTLZFIxtD3OrHu3
hX5y4+Hn8kqHOlKftVWBTQECpSQWt0Lto+kQrOEhlCUicJxfICQOPoyhgJqX
VkJIYwc3Rep4pHRsTxVdnAiFTPE4XAe5pmyLafm44r1w1upInjTlCYTF0lHQ
QCBrf95lDIhRUtzi8SRqUV2wWB7r+EZZ1Ay1JnfiOsWMYTOGaUiIjlQr5Whd
ziK+DDAbqZm0da3tgvzrMBOtpYCj1clBvyx4lQLoCw/+PmkJVMwrUH1Hi0zj
tyYqOhyINeuu7BBu6sOiXycbIG/VrnD12+0X8poY9KQ76gWAyO24THAEFznY
qNWTlNpwpWTmm5cm9ZIyTeS+RTtOLpwRpsaQkOw1yOwoCjcgLdOaIvAUTMfG
U+pbHQcwwkUJ7p//FsQwDVtPRFEOMFpomKir1ASvd5MMkdlg6pMfXdo1Xmh2
ITf1iVSSUCJBmFyd2Xch4ZxMqynd2X5f9xwOj0PiD9xOsZOaCwRKGouT9/pd
j6gdvyX0cbwm8uEftwXqHypjYXdQ5HLWV0qEBHWEu95WVu5qEaAZTenMSSBM
GsTgRsoA2jrxVaDx4FJ+UoF2ObywusNPIjw4/2dHFu3raWR9Xnr+2pRN3Dct
xBdsE709rW3oUT6RhKj0AfaDPy8FEqHLObDzUPE+uLHosAxlawYUBOdUtBr/
DL9b0WJD65hxMVqo2s0fbziuvK42mkI1kGSdUpoMYOkgAzPIla/dCAXOUvDx
bskI07BXCjYMuDUUsb5P2KLA1dSqsHDJqa2yORg21RID1ctm2GtzCk8YTeuO
O3x2TBbBMxAYpd3F1rVHrQS7AdmIOwh2/WLKhK/h1lMkMKMHiHUDMVKwdT6y
Cs9be6tm5yTyuCr/RaHJ0kEeTB9+UTqgZOQr5WFbBAFO/Xt0CSurUod/ksNy
inq4H8OZUVEd/aQBjbwm/VmVnMzT0oSRJGN11C/vmh/krT/rQpW+WPRMsbuX
S/VHLHBn//L+dp/b0TnWoaUCg1dAFSM5eYMu+SUZty6cUe3eKMnihQmXBG3t
3wRwG7DTtmQHpqpVDxImriLXlqR6lo1Fgdz3m41S/d33Fcg4//WiGYZruSdJ
R5o+2szLU0GWBEFveAWyY9KCor3Z0Xb7fHtR1e4Wy10/qZwtXWxGmSVbS0jW
+sxfQXm7QXuDT0qZP6Ldl/sn5NSHxzDq1Q94+FFi+nqSezA+A+VHtOz95wlV
7qUE/kFs6IwZAEOBZBTyRWRcgWkDh9OZQ66a3yrSHyeCaKQ8rjz16an246nB
6pQl0894Oanctj+ezWLhb4DcVjSyBOoDzHRL9QvhYetKBmHHmNOsnL3DbHdQ
0BMZoDQUIk/orAt47GgjlOROJgIY5Bmgedcj/zxj3DHPExAi/8iU+/dGqzSG
NkfULBNLVp+odm+gL054yar6dmK4G1av76tbo/AMzIjFESdI3DWSv6WXhV3C
7qsTvetlasvlmGvbRkCx5unOuYvl5wnsJO/KRnPKj0+3HYmvcjpAouoLQ/xB
P/ydPO9rzKqDw1XMedU3lWU9xgxVs6DXa67aHV1TDhk1pNRrq5RaBQht6qcl
W9Y62Eg0iBDicJSRY+pSgpdvhcYb2h6E2GKQgH3l1x1pIuXavSCUTGLS/zea
y5c6sTGdk/3A0GRz9Ewu2oO0U5UNbKGYdipb5aqKO//RDT4Htst4kUcLC0eK
gkGHALwScvnU1/lvdr3MDNcovFPrdnmvJew8Fut86OpyJoCsOrgcDiMd/v3M
1TCOhOOH4UYo4H5PfXf9fYahcpa9GFd44BwGlKKtwjZSDXxXAYpkB/PuvfV2
zbQVI6hSazYjgZHinMwKVROyQGxlgOzO97KGol09VjNKp17gpLIqgRPP6+b4
z+dBPxTwDb2leYmkWIHzF0PAex2OOCjQd9vcznX+hpOZb4swNEWPCefZnm5s
CZCfEtgH6RRUxRXrxiRhnU7N0VEPF9trH+O/KHcY+ipUn/EKjMg7dMjsx2Kz
wtKYM7KY4xBK1WDzBrvqrDGVuWLJZAQYEQbO7clRbfMr562EPW2rh8RVLJ/R
zpyCDSdqkgJiri6wgGDqY5+5ZWEEnNdGPcfjqPcPTWy3WR/opC4RjGxLyk5I
lFOng+n3tIEjd4/WpnCn75dzVsxnG0FCcNIXnqrtaxmuXQG387HYHOxOdIVN
+k2hy6wLwc+Rl10nh3czDKZlu+kzpE0koYghHr+iy5YHm5q7BOWpNAkkdEHU
AJYCArCNLAdZvaaUWgT/ArCF6yQRGSa2+OVbLV1HMaOQyDobYkfiVu/2OrrD
eQ+YGAyAyeZc+SVpqOOFLESht3o+PvF0S9Jo0WKahqET6JPNPnl/AVUVWduI
CWcC8Z+JDKTJvyXpdcU58iAjqxUDWeqNZGJg9H1RndvWKlCsWzr2yHL0pRPu
3JuDvPsjGvBE/4/5FEm9FVwvNu9PnVcl393dfj/wu+nYKtwZmlxLQkFNu91i
rwjosPPVD4QpOd58+0tSUC/2nZE7XypjPxPaCFUErbhmq5TMUiBHVyGkg1NA
+Ta2MTSpLiTGkk0h7FmXVZ2MhvKzjNBzXHJSR23MO7OhK67KIsJypAWpQj29
kIcHe+Zp5y5L933uxaloZzLsV2OzZmDM3bCKhFfucwaF1UAdHRnOnK8WVB6J
L3D4ZEd7nNSORIQ2lvjrImvJBRsa7EWt434LtfhbQCzMW8Z1jCHX4BqJEFRb
YOONCx0lSbr86n2ctApX+jX/r/yJN5IiRd6Nc2Y31manpqq52INlcbjg09GT
vKsrPaqZmSaxPBmt5qyPjQUeYbt/UeXXgRpchsDGl9YFHMwgGMCK34rVnM73
Cpt+VOWcyN47pr6mO9+L/ekyrXRs65BGSROrymNBNQAvpQYuG1ljcTixBaEJ
9uRoy0ZpVhnOfss1PeYDISoWfW/Vi+lKEDl7oO7rbCQMBge/k90rNiz69F1K
wjAjT9q5X9tzr3QhkQi9yXgIi4n8Qno6zhWMyN3+1kYdMho54HPQEGqMoMw6
/zC8FKmlWGa4xdLVX/FTrhO6+0efQpyT85IDhasVxh3XO/B9CdbsxOC/xsi2
a92p2DL/sxMjCPV8IfG8G9kEg63MBWO0cBb6m3oYc3LQYgab1dACD0SVX4pW
pwQjlyflPDXAT+BaATlLZXhq1ZUDXDu3OqVLPU0XKxfWPurfupd2RGxG3Nut
+xOIDKTH+RfTzAvdPyolZ9Lgft7onHOySt92s63XwbXGqS9MCARh+9PlCTLd
5xaiztaJZeE8HILD1ZT2uIeh62l1CmBM3R5ZQMlEYI+eCBiy9DfKw9S1bpG2
XHc8yHmQDcm0zu94w0iPcf6GE8nSMmvajWTCZdP0xZ08byyIn5OldHmzciNC
CBSxnMJ/Td2TY7cOmSnZ/VrakeBLHIk+q67890GyPvIyhVjHbZH9Qlpn3i1J
2TW/7/KHWIYfJ+bKdkndXs5/CiT0ThEUR2izAn5LIEBwix3wkXm2YIzRh58a
8UGPtVt4CqZdS5Fn22S60StyhrNx3vJe+nOEXefEW2QAFZrcJYTUJ+8nD22i
00IcAScObXFjIo8t8rDUbtOlfXkgZh/8vV8PcYUk/qXuiWj0Iw6zkd9Gplkd
GT9hE0TPOFUe/QhLV/zVS2hJ1xoTEhn5yk+ktYngT3A8oAClVQuqVkCBV4A8
TK0HFcsur0/EjzKWhAJHaPs54d0ghe82cCbk8fUeUykokJ8e5ZDkBlRH5xuJ
DRXCay7B8sclOKlxe2ac5fVkj7qecwCfaUoWo9uHe2mE4YIPm4dHamGK8MJv
mu8FKkFqEIBhNfBqXw70DXPVVAh/x7NE/AVCJAK8liVwlsd1bAdJqyqNiIvw
BrckMUdmlYCvjk+4T3K17aNdVlWfvYse6v1ONLM84sgZonBtyTNNd6YS/Abv
+XDwJRgGkz6uFCmUNhyK8cst24Emmr5wcazm3k5WgM/GW7evXB/n8E0W5nDa
QMmgdsrxOypPLfrFZzgVfx0TTRWF2c4qfZeFu5yPvgvwUOq76SNGmF3xsRd4
gvYh/yDNQYeiJUrApatAZ/z+7ZE+SmTFlliuSrDIW6sUh16ZxLfaIDETg030
6YMRWCs6+uO1ODEpC+mxcB4WpTLYyEQyNLn7qlzhzS5RbqwvZSlO+P0Z9aNC
nU6LXq3JhdGP3VEtYwSuwlpZLAigyV5j41JGTSBbyMDKsYrcxnZdSGZMO+HQ
lyQOSWnqh1N5hEzHjlfGvNMJ7TNS15a2snEtHPsLkWSnfp6IGBjDrKCYVhoC
DlzJ0xQ2EKE6hqivJxdSIK5qa/kiLAaAS3p/AdrPHzdoq8qs+fmd6vw3MMQp
9GDvV7WXwNNcTAo59bQbyJOR0xGNHmcJ+7FX0CnYktF8WBVmzqhgGrky3GvM
/pgkOa4qqbN80ZXq/pJQq1vsZganVN9qKoE/KQ0bO6s0ZaR2mncnj994Em+8
nolzFuCZ5pd1Ujvqu9IcOrYG7/t+7b+tHfIOBauHvCrJ90P7WCCSqJ2j85Bg
MLMbcWrc6DVYI/LtgRqqLNN4Rarf73p71rw0ZBzVImkCM45lmL344REGTS1F
ogRnhtAh5m8hj61W9Gk3j0UBQlLV0b7zuVuJpqs2/6KaMN79YRf9vW29tbD9
Ki8hCXqsNnR/7HHgP+OIepTgmaDk7Uc+neim2b4vdcBMfGowMZ8uRld49wJZ
Zyn0dW/oBjaocoJHwHwk7gq64e1GMtHZJS1l8N6pplE/QiW8abQPjP9eDRSY
bJ8agYjf/+aaEXLoCNDwCGh3+mrBDwsPgmnnRSZRTLJaj5/pwma0TjFn6C+N
xDsO5uUWV1WTY5o1mFrui6Vpcq9sbF7x0riZhJK1wWhq3DEA5Yejly8WdDCq
KOtCD2AGfAO7IsdCquAYG8ndptRxJeUas0dBFhmsAha0gteIf8wr/NNZRxcG
KlrsgWHp7yb2d+ZdwUMBywD7u9cNfVLMpxEvtjEjidwnKwgHzmxFp3O39lon
Lgk8VRMor1qLnmsT3JYFe+HQpLBD71HRzM37Umb1GhWSxvJqBp/qZ3ddfpke
Wle3jisEhvu8ygNyXIp+HmFuyfoafk1mrwg/J4bWgH3LKgBGNK1CsrI9junW
fZdmnEOeeWq4zhx76o7VO7akJyC1rFkS+BUrM6DlTNWVhZp5IVka7CvGrQ27
RQNn5shQ2JNZUH6tL9V8PLY1OaHn0iDRLaitFQMya6qeyHYudv2uOojsbj5E
4GCH4u/f4AMlzu51uSs1Qipv46o1Op1u8+vh+3iwymvZSfuIiqwySxdvtoTk
OZNunITv0jT7tLw4/QAtY9Qttlawl6JCkBfqrIl3bG5IUVG4elHbwYZv/Zji
4wQJUAEl7HchFCB16x4g5H+8cR8Asb7uasb7CUzZGPMwlhnFmsSuyfTXuiBi
7Eax23zQblORbyQgckkXJe5twLFFB/+GKC6uYWBgJdsjjBPGtFfsRZL+BFjo
WQhzN+qKFhMCZ75ogaJgNZ45j38GCA5L7RWx/DVkQvGyWbPPFZFYr8GMLvRN
xOBhFstSh+p2C0FF9YBRHfZMBkfMk5LPFQzUukG/blVyfaTuhwxMYnVshgss
HqSMHYlXMgkv83mP9ufhv5/jxRXWjyFvuCVpTiPmXexbqyCKSPmT53G9y8H6
3lk57Mbgijq9HEpFXyk+PlX1ydulMo2qq74JFHK+zou5p0U37nLsGGSZ2Pmu
StVWj5vN2QBqrn5PBvyu86PPp09SMn1D4PeBhy2Mip1FasqLlUoZnEwhN69l
u1S7hUtJ7hL/+5ZN0hdJeu8v22oH2ERnDoQAbvB7fu+t+xeM3H/sEIbIGKLU
u4jPaVl+lWa+C+v3FEEky3BABmzQlBkb62xzKj3tYaUqLqu1tIbs6v0agaHt
mMZskzYSTb/QVELdAXcx/gDrvx/FOm8N2Eo9928J/DDrYB8dj6ikhEyOKEXJ
roucxEsuM9Lfwk1SCqpMA60Rxi9gtAPYXDLWiMLjA0cDyFleiwUakYZ5KPJr
+GxPKXCOw27PquxnondNYfHqr7XeVS0FGvgJyoqIOvWAAHDLXUuT+csqSTN2
+AyXoLb914KjQhlBrVgE48nMp6Un29g5ifvHyD8L5X7UdQvFU6MCiA5/QdKK
VOifjVl4PH4h9cLmmNYNbpc4EgFz9DRbgaA+MD+9PRAvCk6Jq6dS89oDoP5h
D4W86L0PaBBE2dqSG3n/dFcSmhoWcVCtz3+1EkGey+WV6rvRgNM27joaAbVv
DNL40slPgFQNYRypRz8HDjp0AKui6Gd0L2Esze8INOtQ4/uqaSKHQrxEgWeE
fiyArNHWvHWbWPSKE4K9JycxbiPXh2w27gOVb2sxz4BewQVqw0KJCg6668FO
JCu4omDzh0fT7HSx00noQ78+Ma9P6iXUKI1gC7+/hnaYalgSizkHOwE4418G
sx5TvxpuyqmTvYh5BDgrcJNsJ0iFuvbUW+GzGlQp52hLNIIdQ/WHBj6pT2x7
iQcPALPdlmJQHufPk5jA6Tr4s7ObCkFZowsnu5Qqls5r4E6+3mZ3gvjTUw4q
1gM6rIqdXpCnS9KntDNXO8PqgirXBBVHIHd773h17mGiaLSiO03ZlFTvn3LM
B2jT9oo8qNUCnxy9Vh8lJtmBo6yIzDT9Tx73T2ErGpzRhSXtSVM1pJo0jIam
8dkJsphiFA0FFhZF2DCGpn0vXJpFdkIjm477uhIlE/pcoJ0k/dwIA6lsgY7y
UAQT9THYNA/Lua1rKmZPCAmDdajj0Gm18lMjJDlJlTVop/EDuTDqRdIBlkXM
bUDbzFQUoYS7j6cPw3r/ZDd7Brcr4I4NEWBFUbw9SXIfKUqs0gS1OyS5vpQX
PlyMS+xVUaGV7lVZVZT77T/whC6NwsGJotHzMbbaPxg+7zBLvI8LLX5YAwAi
3b+PiKMCBMgbrVFyX2OpKmEfYln8bTkjQcRJu/31rpzNYr1AkWuDUnDOUV3u
xs7jVWFxldafjAg4YTe46xljHqH++b/M77gsYahR4QVjMayFLbcjG7oYdXcF
cabo2JHs2UdQFhmrMXgDOKLI0BTgugenGdz0ln7e5WCTzZWRG4CcXc9tzYUT
D3k+36d9O6Md7TxYtwZriFJcg8Nbc89x+8pJLurzMtQMgzRQfZwqyOVSaWzW
n2eh9hY9tp3HhF9GJvzdm+A8vcK4L+1I9R1ons20lLDHwFy53NWjdPHWUcdB
BGoZ2wkS5uKCI5unMCHOGbK8yQh93aUNaIZ6o3LYR2V/vnD8Rbh1Sjv1DK35
xptUB5Sf1Vv6DYG77yDCTrbr9XeZrz5KeDKxTWxzEfzWBWebkwpemjmyexBv
bmHVXTMzCzd23M6MaclVUjtQNii5p9cT8PRV01X4PNWsdhJl4EjXY5yZOtzs
8BA/8lwqTkUK/2fhu5PiPNT4fhlc55aMWCoJfhU2IS1VohoNX6KF5dyRq4kM
r5HhADgjuqclNI6OBnPCrTQCpG/jzc6VkXCruxshSkjFvfYIo+8PscDQs8EP
BNiBWzfVkzF/8IVRGLHdn7W4StXpYW7J2NZrfUge4Zw9/dhcOiY/IJ49l5Wb
dA1+/vhjCQnrJvQMHwx6q0NV9JmkJ1Cul0HRCHmWwznBwcDoTWM/FKrXsRvs
tgKwGpRqUo4//fbbiLBXzXWzxF3RFoWM6ETiqjmDANWtOgG3JZoDFcnpG95x
VX+egSzjhOMKXHRKbbY742uCBBtPgdwUckuMrIl3CRTuPZF7nX91mLvqyt8d
N5B3YtclQxu7l5HplIhfupPp2Zflp1wCR0PGa3dn6Co4vdBPNNWfPqCvpABQ
glU1goQ7SzZn/iAS1+xeCOluGNnQEm2hs5Yk0B9RaxRITbNeEy6Jngfqg8WF
pq/vV0DZX2Fq1fmniDeT4hYd5lwYgx6Ctlf9XT2hmRVMqIoYRTAhKsR5aQF9
UxwG2SlTdwQ/OmB77cgNOrg7ukdfE3+r1jxVkYLybuMZFZidV43oYob1QvPG
MtBjS8vOIAq9mG5S6wNAth++kEhmmuR03qH96hp0PHRddG/Ao3+7GBBbtQdC
C5CrXl+FyB7/6uRzUwiRYvU4AoQy+WXIy6GOJFfwKd8AKeTWUPZgDiYjMo3/
ss1xF7+gTfz5aQ48XQRRdYRIqX2T8IHabQ5pofjMNjHClyctt8M2M+8NZyYa
Y6LiXLDEnIFe6b+NfJXYxE+aHe6l3fedbSAsO1igGsQhwlchNlDJYlUitL2J
dgEzgNBEk5w5LPMEY2qGIDx9ZfnTuNfcke40pEmXOzf0cplFBzPMxQqLSYZ8
BB8kfAIT+i0yP2m9hItxsGEGGMusvBHoogWzZDgrXNF3GG5Cijv2anLv1MEs
2MI0HINPBSP6z5HfDLCg4WVrhCYM9RpjpEbE0M0OxSxrbIyNmiBPdEjRy/HK
CSz0AQ1M6mLd57VF4R67VVLhrpB+VlguO/l4V45POl6y+ShsvrW888TPiGi9
r+ctSFavI03fkjjLQTy/fySeEb7/ct5PgRzx3sVQgc3tLHrWs5i1BeKQ4F4v
yF7f+vZBRO9991ZnKdOrM6YPNEXqmmFtT66xi23MHbGjTqOc2h0PjwVShLlJ
bUbpT7PWKFG36SUibPLKLCyp+bs1cAMGW/lTM8P3T92q/7hJCyUw4pHu5sYU
FhptqhLHyEmp6hF3oWjiiaVVGjTR9O1nXPmf6RXm0d/lKMxd+aRbO7iKlv8o
uWdDuZne+JcqvGEUb2EhCHMydXNhWIx8ToWh40WhopfllvgEKwUjbgWjNmEP
OCoDHPPhntlwXEh7fyX9EACRe4q6K+ov9PFZdJTZYVzvhGksKX2yXHBo6DWO
gvJPz/KCbHvjOjMRFl6e9ZWfJdMiuCG51hmO765aO3nZdcGwpULAv5JqcyVV
4T49TRASR5m5cXCs4g2SsTl1ZUbeGr0wErYI0j5SXrWwiGcJCr+69A6pSEkE
P0RJNF4L8OT/LuBm/WxqIR9JEC4duJLTAkEni9QfIIQA03dsvaZf5n347+44
o9U24ijrBEgv5/xRI9OsEbxWUGmuYc0q2576s+sgylwpwToWx4ea2DhKNqhD
7A2/AYAttRxGvXXj6+3hq45+Lpk97U+SLQvmZfZr0xlX1TlEsVRCLSxCxnKM
i2HdLfCo3LAFMh4K1JWExCKYV8PqXyRlLJ8cb7q3ZOAHP4uzm8Zpi62lrOAU
3ITllAVuJ/DyOkhQlrErj/yvOXiPTPNWKXiVZh71C70k4a/YAPYsTURtPfu3
LhJ/qHrj1cIP9PLi+Tky4DjwkUZx2b2yiaWTMCyZ0ulv9GDUGapl4lcfBAwG
6k6obAxfQysepUqa1dJMTGDU7N4iYBFxInXr6Kvg+pAnFYjlRucivXBXVUT5
4VrcuXWC2kOnevi7qpqABJc5aljSbkPpBnZ2Utp2fO1zZbrFXI9QLkVmU9fR
UJNkQ3e1bCQmNzGVoaHDT+0I7Atgix8Qq524Ff/v8CQDQYr4DHRf8BTJM0LO
c9qpbEmYVzVNfCbgNxqRYn8mB980QAW9xFz1E4rWWoqwnYd56qPrhP0gRFct
azX32ju/LxgTa9IP1ajuPlvPt8emj6y4/LYCtG6W5jcIdy//9jMy/uzFz4mY
Oy+XjmJZMogZOdTdSHKsNy2CajQq1Iy+WN1quJRTK4ensIJQ3BIB0vS5A7Z0
XmWduhfN2d/dtwVC20t09K/fes2Wzm5Pq39jHyL9+2dUae7debO4b9HdlhGi
XWPzvKY8c5kZsCCOaPg2tICcGMH3dBD4xx9lCF8aO+BMo9Hg6Q1LSykIDnpH
ckZjXzHijAVg3DUg+gIGUZUG9qL6HQERWSJg66+1SNcLIlkuNKJ9zd/H5vlC
RCgbZxpABw/t998JfgAunT/wwY4a6zEWLfIx5V/RQu0R2Y2sku3cSVH9EdMG
mPkGE6E0kvbZwL8WLNNo27RDrOHpaPBVD/CSMnIz0TvuL+rN9vDbAVnqrSDI
2mPvl4DDG+1NZn3jMPDOdL+kwruYoNkTAFYMHFTcvIJ04Dnad84NAmBeADLM
Xrl+K5BHr26huQ2heH5DCFpDL0o4tJb3A7sCitJtBVdW/Evhtr4i4cj1b41V
r+b26r+HJBVHkVAW2n5jjXZexepTaLA/YwzPVM/Obnt9x3IlJzSHOeZNPK7w
iD44aG3Q/hE6HpEtXlO1Lp/VzJQDmt82J/2ySXgd0C6EeUBd1E2hGpK3Ql1W
SgOAFSgs8049bd/7dp/dda6yRVDFlUmrrctvKmWKL2cCF3/HdyE7jhQv4pKt
GO9SBKHRglyWciQRUxCAYOgPlgT3/KcKe3puuevudkoXscFt/h8q00YDOfeH
mm7eFbiA8UxC/Ne5yNSv3xPzACxZ+BQsklGS8lP8rveHWKJAp1kmrbcDcuwm
bfGnKme/tociwEl/65hrUsw4o2vI+2phcriAIxfOLESqzsS0dtp/cbTnTRdv
sIrEfG5diVGJ5j8fM6hLDBu9K2HQBom/7d/bLtAFXB3I0PecBU5n/nKkU/uY
DMdx8e8GTq4s5HiNJbv7TcZ72lij8RJo+iOQIbtxmPhYpB2Ww0k9Oy/L+LBR
HOg0WqJNy51MsyA7palVAaPWu9g1wqhH9Hfs/Qi8reVHi3qMlaksiBQZxPcJ
UQYm7OzfAgRMEUsUFsVuExtNEQoaaWsQwZ7EGoLNUEO/akCBSsaFb+JMZZ0f
GmP4VL/M5EO7+y6KriVT1rVYrCt0j21VHCj+XxoJz2jNU78di7f89gFeDmZX
SJyxgXfklt+ALqMA1iTbNdnrUPS+50VAvgFiAUlFWIgoUibaXOomYDjQ0tBR
r77vy40dzNDIUmT79QZulxw8JTPKvoNZ0ZfDlrPhZIHsYEouNvlaxZbiCyKR
crO0g9709pJyD/kDNCCCE1tMM1BsHnSG3DiW6NkTGsoFpIVxV3EqOJS62MJX
H736DX/fKYLOweyMgfjO0Q8WBiPBPBwrGE31/V7IE4URoN2gjeOA5BuHRdAV
jQhcpETM9RFu0LLsb3KlEuU5fEbgW9qAqhbeMlbbb+/SOAKmLeeuBNh/r7Ly
VycqJcrsYc34EfGq59twlEDiQtMZXZB9rNUUCMtNaE7FDrkNzu3kDwkqyyTl
5iDaiWAgtag2aG5Pu6NHPqaeiCwXHjWBv5eU0+wbTdKsrQr6E8d+zOi151dm
obx1n3uSXGsHml+c/Fju/iBiosVefgFU31ogDLN5BqblKKQUK7LdY/oCs68T
vkUsDdbpd2XBN8S6oL245lmX4ziWywOIC/1LUCgWS6sibCZtba8N/QST4aCA
w4QimlEBCfgaOzb3L/vHEUUeONbXlm4Yo04jyMMlWZix+wqM2Clp5cOxe5x7
dmsoLV253En/46/7ywYWARrR5poxh+W40R6gLoPN49lziAjO/vGpxH7RXV0I
WhYOswVWS3v8pEQmugokWm99ID3+UlhX8gQ89wpP+tC16kl4KjNwL/onGxVC
G6CZxQqAEyFNnfp2lTnopwAGySB0LLgeNTNw5+n5DvrKMtz8n0kK4riw13bI
gB7pk02BF4yL3wjOWhimrYTilnk+QAstdosUa5sdgtTqGjzcDcEGdSUR8T2E
HG51oH3g+dlqLkhAKndHh3n0vQJOZmbYBmnJPH+8xYNEIuNOzpIpTXHLLuQ8
3KjHHw8N8V0w6d+YwNNIbigBDHT4T5AdKHYyWv2QtYYr6pDvHH/9DDHw+vWb
PplzGlMjcljRhQ1SL6C4AibZzAwYUXbM7YSbB5pO3UpydTW8MM/yMTsL4NYy
ZBUpBDFiV6KLImkwZKJ6Sb6VH1du3iSoSzhAlC9yP8nuuFFe1NTeiq0vwCzV
13clInQbPZpMoArmLfRMMBpWSHl5P52uzmD5618OCkRmrnis+B3iRBTOBgyr
z2Tuvaoxdgev4uw+9cBlo2dI6d2I2OTtha4GYmCuZwAOk0ruHB8wkoRLMCyN
PJVX3LzQVZgexeItdudqiTE7pvbslqlcIkEzesQ1oQClN719GFsLGVi47ciM
AAof0I6YyQlWAEJOV0VTWgt5MT2e/KmH/J5qWuxMeA2ZQnZn3zICNsMYNcMb
Bdl5lFCSNrEmqVIrxUQBljGaYVkxa2N5jmDbnnOfL8Y26XbX9HJOc1R5ftvF
00DphP46LWu3pJVG9zjKadOt7eMi64L7GcKSnkaKVr4Fn+/9q3q9X/CRwMMU
hX1tdqVeXrx9JUcx+MvrM7CMpXo/eOluKvQ6v30Yf+Uij7L2t7RuPnxsZMm/
8spjaGNo+5isjcptX541C4KNAuONM61jCoMpQhBkd0D6rFYtPDXXtkRlHBve
aMirPnBu91Vx5LM7FyQTEpMReIYmM+HQ9r/jS4q8gqZufsM65eUfuz/OucNo
Bou3APjeLOgn+OkzrZLWPVsOfPhRp5fx2WThcdM5o+xxnmHi350tmlpnDFg+
C1b8mfym0yGT7Vyot8lIZsEBJm6LCPJX48F6+gSxjSbiGLYebzk4k3duNj2W
YzRZ4GL3Lu4K3/R+1wwdz12IRmVsnaQn9mk/sXnq7j/EhsCAY176c0kGlZKM
mWvZecg/vDGSdmE/yns/ijGboUeO2p6qUXdiveLtcafWzZLw8Ut8KjOU0fx5
09e7AY0rBB1Oeg+oqWB21uV9aKM5ieWUnsuSyxm1hpLVuOEdfU8jV1COBrIj
gVQdds070XBM4S5/Qv8mBoYn7uqjI3c8aabNHmnGTgU0s3sI5jv5u0qVAx8T
gIVnyFjfKL/En8ZVfwW8TbQk/gNN18CBmNLefFj0dfPNg6yeMHyJvcuP5JMO
xDBUbg+QnzqTI252i8hBR5MR/1xZ45gA3WVsPFFMpp3YUhobNvoEj03RkVrd
1EdWs/ZJ+7hoDJkb+QdAYA91eFG31bFSgDkYSCQP4npRZPBoYHUSZZ+pw0Vb
LQZFvp6byOSqajUqu6c81Zt/I/1VMpZeDG2iX8PF5oGhJt35STI/VJ2N9nCz
hSy2LkkgBJV2yrvpa22K0LH/VRYg7WRgq5TVkA6ptnhtmUZi0UpKUuKooP0S
pPIv+uGFv61U5SZOjZLHQUtMhBAs9PNH35V42qScFri5xXMdiFYFlJMOLDHk
RtG7x1A31tldFF0/iQNwTyl/nl1VYrGK4PErqGx4WpgCa0sYQiHJOvC954dl
n2wpN/YOiMkQ8NqFx0G1NHlGOeVjs0LJPWASRqqykrsGhSoRUuzOM2mhyyFA
o+SmEpUuBL6FCq/Oq9KbXRsr6Pr1Lw7pTXlDDGTG7Pn7+R65xOASyV7mYe1R
O9KaaIqfvq+X94cWKBR2M3aG05Pgso59yOkIIrZ7R+u6vzdCRT7I7buxYBmY
KEMaQYAV1ShYesMQ3y1qq3TUkjpCPKwtKoTXm1zPJyswga8aQVaG1nLsmOAr
tBTvYMReE30dU6ElphHXycXL21Kp3RGVwfCgP7L6uX1L3mZpohsRVGVvXs6P
jeVlVIunfcMMOLKQFmiwFi8cqYlpyVgvlDLvifg2ZQ4Gg52ojjvmJKeNv7hm
fvuR2NCyK9f1w49zrEy9qRbLUKpGPs9vLd0oclnr8J70kVtHvIrebLvJ/uTG
6SJ1GT14zxl0WaEqeIR455dqLKHjzIHIp9vyMS5Z6eSdBZIwpyQinkoi/Iu3
u0PDqlOSU/2dnwyfUq/VrUJ9xkS/AzTn5zMJklP5ClKyCXQd5qVM2tyEYReA
hx1l3X+sVhg2K4uB1MimK38ynbQf5VgOLLmoN3xu7So+1JYWGHpcxQq8qxZi
9WYDBDxxQO0HrLeRcqPzkeBif74AVtHEVujaBOuPCmx7MqZJsfbSl8APvqEY
Kb9y+0Mf/BhCOwsnKZWhauYdpDNEudXz8qt6mOpIrzPQKivZc2+j7tzqmevI
XdNRFehGYC0a2Riqx6gsLnTwUydvKrzpVTMDOssYcr9EdlcmERBasYUvL7rf
4AIpTOgRnIUWNUqLKqh3djCPsSEGdVg4wFl4U0A7kHC+eBjGDSWEWMsffRwQ
qq6b2kstJatHrFjOj2agi+QnHyw/bh+xQ1m8d6bYjACtw6OdEOAVJAhNV9U2
pTHcLqqQmhTCfHBc3C6qTaAtIjniJGOA1UDmscAwll19xR5zyZ4kkxGRNkz1
S6/JpEXlNOj+gGu7+MZ1G5PROILnV99Ego9i9OUP+LvG0RocNp9qX4WVSS/Y
U2hFEKZ1cXbZvpmlDpIaP9kdehIfPZQVuo/kwJBESPVr8nism1k8a41lamF2
8thFnokg4iRht/rc0rzGR869U3u2yIdjv8v268kAbWqv/eo1qjSUrkmIlM8W
ecZ2R5uQ0JzizgvW8zx3DLE1O+at04pf5wQE45jZldm1ZuZvM0TguiRH+gUF
Mj4uh6eAca7fYB+Bcmc26/4ohaACczNcAid1NquvZNZktcMS/mApkZcDpOSi
1mNkDumFiuaaO6XQ4rW1VGsYgqNw6KP/7edOf89NFflZa8DwfKXzGuxMs24F
4KQoiso3D0uHRgC17RWrRONIjpHXhsSS7n0WGv2wETbcf68YK4d4w5s2PMgt
Zzz1tkVoxzUapjzyB02AweCop1NcYJ5LAA2dYv5ct/HDg0PMdyLRhYb26Gj7
hmU/hR5S0U3a3eSQ7tE/SMcy2xay7xJlQKYl7frPPybqSn6IMSBkAiwE2nfl
soadDJld2hEVKA/1+JacjCLT6Pq62a4vcahNaMk2aLisiDyXCvYLY0dsbcLL
OkSB+JHJ/jZk0d/FwZn1PHNWDGCr5/d/Ar4oq3NOH/SmALQN5Ln6sDLdTf7i
FiuH/hkHo0Asr77yClH8yZA06cU1fIEdz3Gl1lOhz0XxeQUrJwdMwfbHB50A
sZwCha1go5XbhQgH9SnD5uF4NeoZb3C7LXgsul38+1pXV/+42LcUuGtOzy0Q
kOC35DPwocVOqrmf93DeGzX3dAr56Ta8cZi5jeZkSMjpq1YLOI1pcMI8xZCd
N49kFrgctaH2IK/rgHQsqwiFSjkR8wsc1xi20UpN4wmKeXhGDdJl+TGK1DSD
a9JFhU3NFRhujecSiWYuzckj75017SA4ug5+v7EoxsnlOVOnS+2EBdTCAthl
h4W5/UNegNwQvtbADKfouidlwHodPUnu2BDo2NUAmQQJ5uaY9pQzXUb1+nqb
Qez49JLzxbDWNF56WMUFVj37+cMPRCtSPdgBRvONWy5aNbW5KQvFb1dqs/VT
SLNby9rgyFjCSvauJleaqbk3rvaiVrYuCu9TjMJEvK49iI4DIPljqC9v1tjt
L8PAZKMRDAQ4CfOqBzjJ5ScDExcO9Vc8AqIv2/3M+fKeubH2BAq0QvunYHOx
JCXjaaS54hE5Tll/+taZIiGKpUxjLKEZmGEQO5gzmSL+omOmMOt5mu7Nt/+j
RjHLosfR32Nf/lHRtapecJ5scIF6dyivQn3KhGMMfOG2qh8qyoWXLFmkIy4p
PIX8BEOkVRQnQBUQv92nGlXEhZf7hVS+DNhTR2MjNikLDJWypudke9TOcol9
sPNJecx/F5649fU4XcF+EyKMkZ5uqHVoP+ohCI3oIrvWGJPjjVE6AEE5wY13
2crTF6vUncEnrlFxGyk4ElpeQ24S4bXGjjsoo3fDoKfK6F9r0WHsZ/HMKYdD
FBJ7RuNFzPt0vwWLrTScdzNNYV9vQv5OdMH2m+ATo1k6ypBaaP5Q5+CSjTxv
x3VbVt3nGlpkUfg/AS+V6duVSMOO6pKGBRdNl+FvSqEga9D036naToaacXu5
cv7LYIGG4E6hxuEGjnR1VhO558SM8ZuY+h7zQfdQJzOIWlnEVdRM+wwpZSDB
Ljb2q9jjkw8uxHEbxtrBMSEx3jyvjsiPBtQ/LFOjNCfDFjhyIrPp4tRSWudc
ttKKHbJAkol3Vi9/KeDaYu7oF2uKV6IxXHWJ6s0PmcfGOoJT2nXU2WvLS/Im
qjXQ918Sl4IK+BiQ+jsAjkFAyXjRmDcybgEUc5IrveYeY6MHWEkfHE+6QEnQ
V0hB58JNt+PGggeBHVF30p2PNWc0TjnEOgantzYK6lrerAgRdKRY28FKgn8x
nod5KxnKFPuyalA5aITIkijUQBPURywcvjiqT9fJ7SRct0zOKRedy1ejTMwU
vtoJztzvAH9pH4s73eGmXbeV17P4waliqoZ8q/lh8u4fGXR11WUAOaomjG4a
8XofzsiXH1dSeJSULDi/X5EDBHax04o0KH53LRqOewoZi97neB4qq1LZdw0i
xErYloucNaaEqECnBVNO5oLjxUC7uJspElLg3AliBK/YNXqJVF1oSF9PSocz
O2wG6tGHHKK9NXgqPm3bH9C7iF9q+IHHC+siQdjKY9sRSGW+VmkBuXtuh7rb
Gr1nL4y+ufrKcdHVK869Yv4kHwrEwuoF0ueYosI2Ahe/XoZiax30VlCK+tk3
2kxAnBZHxrT5g/Yy/VN43Ix8IAtnA69fl2i8v9Q7wbGeFyKcNM1Bj4LFk2Yi
C7ZHKCbeJO/FfGJhLe7dtlydispSgfStr7S7/bS89QqoBGUH+2qThk6K+mdP
bhhz0dYnmjd1IniM4P1P5rD46zvarwT5G8D5T2G4X5UqSezJwIlUoZOpuLTr
QPDziDm/aqbq3AfTalCNuJUJvTmjcZWdCKUB2jx/6kzZufySyw+joYVPqTPD
0I9xdXtNo0czYlELwDfScyUAFu40KmAAvkhBJWK4Uf+GBvBLJGd3XblbB4aZ
dT7njFw8QOytLXLiwzymQfW4hIGJGklp0/iGF4rix5fWMJiDh88LqJUds/cX
tx1PRMcO5CI+a4vjS7qyElHSHEVBWLHysoZOwRw+VDIJRY7V5abe2h/ge07f
HSD2ASGVZeewEFynm7H5VUiR1Iyv7K069eqG0Q8J8eivzXp/tE0V7KY69mkz
O///QzO94NYlpIj5ZwApMiXRLJdKymVl3stwy2azYa7kIgajVA5QiRQHQCL+
NPujif1HhTcHPjI0RJCpGdUyhec49uH8ZBjCJfqitC2fw6Dr8wm4XV1+H5K+
sG+FW1zwQm8Sirj5B7hmD79eobB6IGrdPkqRwORiXI00RWxZpgZLH9rjWzuq
CVfLgFk7rvnQFYmZTXprSCN98MXAPY3wmE/AWsYcrzg/AO9y43rVYa/CnmWZ
WfZdwZnN0/+7WArnmwNbu6+hNESEdApTpGHXmF05sC7mxV/x8a3qE0veHduq
IFUQNUNDsQ9JptuzyvRCeifXkB3fLn0tHfq9TKKynIJ4UV6+VyOi330zcMHp
FM1iuRPaUsM0JQ99GgGJ/MikdfsQp9JvwCaTZC1jHljGCUW9hI271T1D55iU
ePxIHmLrNRrBvgkdbLJ14bi/P75mZlQVfzP5uPsq+xneClayzVfbQ4z7qloM
KpUCE4v6o6gPNcEgYO/x/d64wIqeV2NXcJefwkfkIm5BWNkgOq6WQf82gfQw
aFRd5w8CRvytriE4riJB5rfLN1lADePcEe9zbDFIx4joINfsIfasxFNY0veW
6ZskMbFlrW79L9OF9YiBYQoghXAPriUWWZwC6P0lkkQVftrcuwnayJGo9fJv
WKg0gfCXLwGRT6cwqgYwSOkGdU0LbM8PlZdS1yR6+qULYYfLsJfAO09xoH8/
7qX9X3t6i7LlvXIlkqhrfM2cG6u7Dw0ftQJLbJn714jkSMipLFNitMmGaBLN
h+fElZERCstWfZQKVFsPtL9JjQcOFi627tAqP+miDCUId8GQ6oYM9YBp47Iq
R7T4B5gY2jMT1JMHUWU0lBvVTQH+qjszGUAuuSyJY/G1UVba1BbjDOLcJDgH
dR1yDqq30rEHPWAL2yCAxaq/im6LQImrbb6tllXI3E4gACO6pGPIIQV+EGcU
EHEY1FZzjNvIxFALHCX+7NkAGvcYR0eSwjBSbH2F9cbv9tGmeA5O795xKRES
vqvu5g5o+U36zc07xq6HFu85IOCghPvujvtLwspJEGd5b/uaNZkjDUe3pt9U
MOh2+EAbwqCcvtX3bjbFtGwIYvYNoDFG1/ym10/ZhHNrYen9fGs4DT7Dsf4J
849d461Irl8/JFFEWbF4V+JXUazHUnbQoI0kZpH8mIWGIJxrh+CF60pzh7aE
WJz+tzZLyle4jNKX/3Ws+tdUgSw2vb7vuwozRx5g6uK4PKeGowS+rBx2ebD/
uHVEtK+AZC+flWS5UsD2SwoEyMrqmQO/NJ+jwtj1rqBMEXZxhNdeEvFIP6H9
JggCYtXQ4pbCldht0q2qX9oGk/7MbPKJ/+sOTfA8li3JN0u+86DjoWodMeqN
sxx/oj8gupEpnsS+YWDJLyZuii1Vlb50udORdqdVVMLr64Vy6r61QYsedMR1
8Pr+LkjLDlLynGiLRji0Q755RauvTbuZ3ZTUF8uuOGEosjnrCmPNjNa2Hod/
TipugKwZN4funi4aQtQMxJDeQuquU5euGQ+Js/R+GOJhqbeL0kKydR7yW/Yc
2w7Y4aSZWd5acuVNq6wKWZim1DWOrwGApSgAzky914aH/fHOZVBJHU4BcnAV
pFbespCS2tbOVU2fUrkzxtsCOUEc65skPMu5yoy5zc6LtJlVVBjVtir9I+WU
OjWXYUulBbGry5+inqVde/gHVn8sq1Ss40lr5forPkdfqkBDIn8J7Wh/dSZG
eCk2rrtsVXVXhfinSt03zCO9wS1IDudqPX8lnbW6tUl3bLurjTIHxRXQR2LT
CaMxbLLPcYauKdXC+La7sM7wlOXtR0sALqqbZy5LdMAfavgwmBcC5QcIvZbw
D2RDZ2msDSB10QLsrTULLYhKf1rcYDJslGGhRemqJwXqlQFxKXB3lB6gdGjr
rXKlQiBxsXAkltfP+xZ1frAgPuSPBuww/0d8RFouZWsIlW3c2ny2RPI/Lhq+
k4/WzlWKFuNiX1nzkWrqApO5OuHbMlWsrqNNMjQNK70xPrQYtFe8BH2v3rZQ
tcxy33XSjf9QKhEahoTd8EWom/GOJZI2edxIDaIL3XKQoL0mowKyDBwqpOdU
Cqb0a1VF8M3reIbVzq5pa351QiyRGcvHO49AxHCWN5LMAVbS7r5ojRsXsHG4
fjMhfswjahn65Ns4OllejuLtDW/VIk4GSmQIrcDs+iUWXC1mJJhgskDV+r3T
B1nADYuMLIf3VZkzYK4a30jpd+xKfCI2dSJnF5nA+KjT8qkedR2yfck5XZeb
rGtW6jml6azDdKVvXoxEyF6DASQUZ4f1sb+dscLb0u3rxvxn8Dd9vIISBUHD
cNXYFEtaeYr5HZbPlu+Lfks6z7sK/LXusq3FdzwpoQromNZRJ/UIP4kSmwrR
ij9cqOVVhBlLWG6cteUE4IvHPZZ7JIvvRDMY9J3Iw2ZzeKuQLKPWo6jJcqYD
L/BOA7Nj/3Eq7m4zgA6t8kttTyDFuZ4BOD5v68cwOUkioRhuVlTaP13ZToG9
GmcYfpTAUCoJLjdQOO+t0LZ8gf89c87j/geLDWJA7VQH9NOKN1pGZqjTi8K/
VnXKLY53c9BDQ8+Ob/nNCUuEyLs6Fzvufu7Q1qW7odDwpDn7/mhIevsYXK+l
nrsJ2caAQr6auRbfJrsljE9AQTXGBnjtGRVs3lynyVRQX1TPgbvvvV8Y5yGp
ZFVS8qGGZNoegn0b0lvI8+HUoC62c5MG28JSdqwllG//+6Ol1CDhHjytj3Ru
lEy100c0wURCqb8eJOu1iQcJYmqDDA9uUURR+BKyVAN4UMjSruiaTXJaf355
aY+hbnv12eQ/gBT0/HWYqPauvkbGfB6MCmgL7RtX1hIFtJ9CX3pVp77W8jlR
uowOAQVVhhkHv3PSAiJ2qbg0kO7tas3MtkTW0Upb3ID9X8PZNjrhU+LOVQQF
N8+Wqgv5IrtOYLyNDkgtbiISdkdLTKesl6QtGFaYycc6K0deUSpWs7BPhxFA
7ieB+h3xi97YiVslnANjHo7jMbyw9DQtGdRWaVPUDkWnmKsKPe96W9iS6+dy
skkBnSnPYnJdbxbpnxO2OkU/yhCYHDcbINuQU6VTX8NO6Qe5HIrSYGf0PEa3
ANc40mNHAW15eOK/N1qE3GVEeq4KE8RmDKWrIeG2p8pt65tSNBNdR9j/GADE
IQxhwY+e5Wy8IZEW+wuZLA3uQQMO+rqcD3viswg58NxhHL5ke2RVxS7BVHxr
RIo98ULQqwyXgn6xV4fRoCeeS15gCyfv6mOc3fuTnfVeIEXlHcgEhRh1NdBs
zwZLRitOBABSRop+xIxWVw5Da/XBB8+tgegtQiHtrLGVkYdxTn76vDsWxVs0
J03hbcV2MSHBMa3lRrbj3JNttqI299u3/N4oTW51a99Jty+FbSrkaRw2aPEY
lLR3zhNkZ2CUWY7st/WSyWqbm2bcZUwouOw/ip+YALz6pB0bxqzJJ7hmer+v
UOWskvwWkkC6TKkhLqo7vvGzV64dg21Ud9Cd0ikWNTRi+B3IZ9v9X8fu9oz6
DT6j2T4Rs44stFZSNET8C0He2GbPxaF8VmRC+iOjQh2Aot9p+/JBlfDfut8y
K1XQB5bAyRhqojs86eowas7SPnujo8Wk7MaZPdsPTMKDmPtH5E4pYdrlnGcG
DdLa0KWXhm1rHlhF0cHm52M2PNX8DlU1VMHLv1kc9dZPHqeuEEH0lE4hA1FQ
UY+WMMbztJw7UmRFiYWxrwMfr5dbfSapPE76LruFXddATy5fBhMCWlpUWCeW
vHtH60FU0itB1flDXBRXNQe7OenIHMKkNWXzv1FYtXP4gjDN11JWq28uZBEc
9B6k4SsDaG9g7V5kouLZEW2kPilhUCEJAQ/YnbKNb43WRXFGxruZUgon//4K
7A1cfEdxk+clx4CN/YG60Q58DHKCOakQUYOFyk+u1uqBAjZtLYy15wDMvmdW
NW0+gx0kY9uD6rmbp8ieyS7Bk/AHMpLlQBuUSLcfgztzyO0M0GQk0aVlV/F5
BHPrchGyioZpBZCG7pB1OJstuBSbT4uGyR6UPfnvV6FrcQMcxPPEXx0lWWrP
3ayDB67CQ3mreAYDnT6aAtwou9HMNiTq1doNIq/0A88xUZQoEwSs6meWHN9g
gWS0LhkWgsYTsO6Mo+L1PCPr5tVE60hwyO2vZPQcLcjtPfWgiCJDfQabtL7O
If9dJfTFU6aMFmclh8OEkCo4t4EbzOvm/dCPBxJqeEpyYoKCju05lr45Oeow
z+pEUcJVUe/8N6CtBqGg+35avTq+OZ/846drOISAbi/54/BkquJEEZOA/7tZ
KEQ5Ymwj9++imRqwscfKJQkQTDWRSgyDapWtIhP8PPsA2aL6O+ux9Pg3l2Il
itowXI34OJFoMme0Zl5u0ZfWaP0T9ymlU4E41FiuYZNMr6gDZa9DDIGla8X7
YCcU4FDd5W44SQMRQVYocZZTB/gnmAeFFOMozGLu5q+1IcQNKmeh2dyf2B7a
5BFi2V0xZyS3ZvKgY5CBHQ5x9Vd8/ZNJPC3g4LvM9aUqUbv9qLZ9PQH65tT3
3lQQHpfQE/lhfzGLNBrFwyfqj6gvgGFAcuHzBScSywaJMc0ete5wQ1rz/cJg
pfzQhnotYNXDtNUrcGKJ90lIrU4ySyEcdB3y4J6o9FnEVTbffs6EP2CvVQBV
MbRTQ/itdWgOxb7AoKQr2n0MhVESLToHZafGcq6xCkxVgbiAv1u9bXp3g9hH
qPeeN2oQq7hR+LkgYs76dd5LCOmSLFYp/67YzR9XNIajgMJwxtN9Qx3VMMIZ
/HDqCtZzQZuXC7p5p8TCB4FO7xDVdhTgqHbqMJSAzBzL1Zyuadm0K667MgUj
zL0pD7G6Tsc56qIWkefGs1MIOuSEU4GqTHSJXOnQIOdg3rsqq4qhFce6Jdtt
eDGhoSX6f8Qf3jQ6GykDsMcYIj9HzpwYm2nYs3hU/Ts/3+U8X+BNA0ntM7AO
802yvFlrD8kS7fbzqKBjamOyYi5YB/2/d6ozm3izlbYXJzzrLWgGKMISlOFq
oQbPJmZJBZXRUS3LoKq+5UhvwQefg4hbBB/4Xrz89aemIbAvd2sGsyLr0Q9/
lzsKTbWZIkfvtOubAS3PMIoCn2p3n7jphKh+1Vqof+014DyK/aOe/MAWmg1b
Axj4eYrqzGU/+/sP0bFHSd3YiOIPPBOn+WFredMo0Hzcv/z+WekrZGmYqJv+
oZMvBKaAXx+bcGhlW35y1IFKtjkWv9YlHbCnaEcQamZxdRtKYSdm3ftG7ge9
2SBBKKdYpW+8KPmwmoWAA33yflP2zZSvvOFGzMh4iygTish6KmazlaZsl7k3
R4j3qp0tJU7iHjUImbOcIwKrYGfwJVjL1FRN8krohItpiIzKsvIDk84V4O/P
5Y+4HsApUcPRPmQp6rTbWyHkFy0tg8SMOmbFPeo3IpsHrZe6dA+PsHEVjKSI
2RTgim5gkAiJF97PXCSqpUkgf9saE2K2hZ27dHaPVQ9PiVyoX6SobHf0ERJb
6rj7Xnjd2awm088QnCvjMQES8/BT1HNbAUQaKgofxMWye2BAi7kziQGeqBar
1k0C/YuaN/VZhaCHqrFKKwGPvu0asDHI1JGJmLesb5AZ897HbjBnm/Qvh+YJ
ZhgpjIyrz1VEDFZPD/9RfE4GjT2bkrKp0iMGaj3CyWPIMBbhLSrIUUCuDJ2n
rlLcZ06+PbAZql/qVG4lRm7uHnWpXu0bbzIRZ+xfeMycHStAOts99SuYuoGb
LG1sRSRmm14OoU4xTrzsp9dtBbkuMoXIlKEBOcCKeFZTaHJezEedJuvt1aOC
QHseIwwxXq0IfvUVVek3GAKXoZi2JgOaJPfi3vW34IER2PI9MrAV/yG0RyNo
p3HwVDvJco7u7xY2MDWP82LZ6R1bho7GZ5EfvDyRScV0HijNDGhMVvXGc/09
+WeSggzVihbWEzBeCCiNP88k1gCoRQ2j5hrG3L4RPWabZJeN9qYhhJwZh6QE
+DeEyDVkMU/woPNPq+0nrwpbvaHogrAXfOe6rVGgoraiut4cxw1xis8uDSuk
JmBza04eGF5/wUADvKfgqqz5mTb6THZuM/zCkLqtWpN04DdL9mOohPkdk42s
vNr4C57Bp+7R6xiRMUs2dJgK89eeiPU7L3PTXmNpzqLxISwX0d980ta+Sqxg
LkoJVW1CQV7Kz6rRPHjolSqqJm+NfVg3KxfFHQo2uSJHYkK70VqzC6As9w65
A5w/0Ae6jzIRkIuf4zdDz1bQ/L+nRhBfo4CU3p0rVtVBH++d5hzx8LKUvIZk
i0M7YrunS3D0ygAWrgvttF/NukWj36CK1fqmsNjkytY/ixhpkVPpuyk7o0Ld
yyWBMPaVNSkzYXJeFRTrfa8AiksE/HN1rFFXKuBfVSqeeDZG/lBH+icM27pS
+GbW/e0VnUCA1jxczn/6j09LRLAeMuEWWC7pCeqwDyS3bgsyRwjGiFZJ1ck5
u3xhuR2moQNfyOyvycZzxBxIhbTHP7WRF2hijldGOo2SgDkubBlC7t7BLOq0
g54ycb7YZHFND9E0TfFNgYn0sTby8Agyi0uyPGHmugBN3aERJqt+Dly/X0D0
9c335Jq/aLrE7wEU3v00IrmuJsQJQCs3ZsLs9zknBKdNGh9Ata+oZypggTe6
fFCDVfyPyiovDjFgLOUm4iS5RJKYWArAc6t0a8iTp5Kc6RzCQW/884tN4Q0E
kAfkoZW0rvkuzk9/Cbh3SkZPX6x8+8SFlpvo9C+eRUV7l5hvF4vrxAMpUmn8
gSx74PRImYk0XjCOFjlUsxkSp4AkL8REOvvQOUwNzqbCqlphPeqwfHDMzDQ4
YszOjDzCALSJClTGcs3vl8AI9r02LOco/0i6S/5GkevrQJ87QBhI/kLobHTa
a6PZnE8qwvi+c8N2gpIUioNSp9w9bPabu46992/TXAHPN6yLeoKq+sOo96yl
1k4crQzCkcXxhuH9Gd5usIZLO/yaV7WOCBBk9ztc72Z9Ie4S3argUAU7eFix
SWse/CVn9QXbw/C7p4Lw0vVkN+rVnJZssXwtHBrdU2fPnk5vWQX/Xc0wM4Ah
WyxkT4LmgACTxDdOHGFMtup+nEZGddnmxzTwaqwq5DKFtebaPRN3uUbL4y4g
Yp8pky4sKXZhMg03qhC1wVBDDcAXts1DHbYG2ptKcmedDNA5SMqHBtBPSHuZ
EFgqzQOP9o1ESIwB3LP0BNzyV4OeaGEQ5gwGdqppCiTCkmJJmHnpjol1FFUx
7VNsTqherPYSj2v2gWiPPeUuKPdGgK0kE+PkUsNF2jhLQ4uidHdX1SQDir6b
EEMAiik/45JtoKJqUErDXKNdhOm3iS5MLZhHLsf4Arktksk0kfEM2FTw3Gel
hlOgYeuMX1MAxiQb5lup5VEgr8YnC5fnLpKhJIGJzCQ/2q37ctf3Lfiliiqw
uBHWCi+817dcgPPgDPR8LG22b0UFTsppUqwrJu0ksjV5uo3+oskpOJu00JAh
iCX8yT40F9CL9SPkyJm+3qvr4SjQvdpgmjCTl447+fnLoCZIc7t6mIcZLqQn
S1SFRWW84azd4bYDWkQwOAi/cIT/+aJACfxcNY0gGnkOQMK827eq72jqR9mT
JwXhApfXxB2EsjkXhdpxaNoCuD+WZKiSTFVPcm+YAekr+2W8AwTt903ZkND+
Qrlb69vb5GJefrdBbOjunsBpEFT3NVN5EQleG/MsK3JNDOQ8bHbaNqLjBur6
4KXdpEpCE+vAkOEWjEB5vAETW1mo77YE30hfKCCcsmUR5/nZ2vbOCkHO/VrZ
+/KOFdOcdgxLwgxX9oHEXWtwUWpGA3/PQkugqmQChHSzOFGaS+hQVgdq2rr6
9o0DlpqN99YYo2H+qhzYwV6Upz7hnsVjYJALk5mZEQRjxn9wyEEiReVW1VH5
iKVnJln03Dd9aStw8xBYSkDVnRnge9qq+WnNQnW6XBdFYu/K13gH1QDT/ynT
0qE8b2vYKTn2pNiQUHf82e84HzRnlVcnjNMcutOMNm9z4IapvoeCu862naLO
8sIWPq89uzTEkZBZMCXQVqOvqNXPW3rTdsGSizBQCsQQ82wKCGx0Bkc4B3J+
hhfIdnbe2TQQUqIZYVR4OAQH5YKOkBptj0g1pGDvXIRGs1Jk2bTi8+qcSOuU
ggAm1+SbGDbgA2fjEFgeTNAtZHTRYYAQur5Rrpnxtbj4/h7SVtjmfuSr2sTu
8rPdtrzhcLeaPenxp057gQi3pVhLdsBQbHNI1Bfc6WnCndgGSkOmiwbJHW9m
taGVGJHQcnPGOHmCK3hov2Rbyz8ptcKSXlx+hey0Wr9b/98Wpo11tE3Dg2Xq
yR0TjjPDzfVLb3onz3CmXJpoKQ4/Gr5+jI/nPIA76RHuj4skcRI/PAFVGcnn
BgKxkYGbswXloa/pN9XXlrAN4RzAVC0l/dbpeUBZG3jOXTion6M57T9oHmkg
TtHu++5iGBZDMlNt7OF5vq1gOXnBBkwfnKTFVgS8kIzUz821Qu7fNM19udGm
ADFYMkybLR8Yzyn6EeoC+JADeo0RrkW5fJvl/egJ+lBxnVn5Os6N4MhqbcLc
K/lZm0zPPhi0ybsJLnKhVL8HooW05/ynFxfjCiA+Or71kF2sVfFRrumbGLAj
qf4LakxkceltE9EnrU/YzWhqMfboeJDC0sb//Xp099/mWVG0z5IGPbLDxu87
pSXf7kxYcNMlFvC910GpUqYdmHaqYtWOeFJDHB+haItyYTv/CFGOUehfa0uN
gtK6imT3RYOafmLikRc1WAsTkTgKIQu6OsN5OwPek1sN6sgPuh4PlfKGg/eD
qpeJ8UcYEOF+R99H7eQ+uK8wuXjpQHX91t9gpvq/NVZvkZ9dy6KeRt/oMNtU
zhwTvhRYCieVnwX7IUr2T+hTR1r9o1ubMN4lB/wJw61/ZT8eg3N9YAOhQQQQ
gWrMOPRcgcwx2d715l0dnUxpOvfzLG+4gGql8jjHvH5Pjz37SRGoVJ7TGyFB
/YEHQ+GIjQtKW6k7CPrKwHl0ZV85K4UX5VYOqvatnihDFtsxxg5CUa9e4tCx
WY+pp3r76Lk+AVPY1Vb4h95M6bmlNqaMHwQ96WP65IgCNl/sJky0bXXZR/hM
AlFiS4Arwrf4jyis/oA8uM7Yn/7g96TVVVmZpSeilMkT4QWfND+/YufdbXZk
1B7sPs7zSdTpUvQFF/JlMd34+cH4sc/UDJWioE0aR+PLHyAaV6B9TQLpdCHM
Ctb4I3rU7WgVxUsB+QnouSZTo0vEYhxajzLo+Ber2gYwcGLWfxYXHGmmNH4H
DsCmX9thMleQP5Ft//ew03vijL8K1WCtJn7oFj4wgXo4uO/wyQ/4pGtGoiJp
XRnZLQg7WfTpI0kKDDXcHxyOpe3z78PbIDWSpgGV7ciHu4cfCy6/HRFEQkw8
dMxzAimJ1KEeVWDbT70qrsIgBMU22IHf2nfXDGK2f2aLyA3MAmHNRJ8d+F7+
9DxQP+6O/QjlXuNITYHJZVFBnvaJXKM7U/VyXrY5SPFQwXwWyCfU4fA0D7eB
hzC2Ml6PsP4VVH5NNkhOAjZV93dxXLXl2GEEvch8hLN6qkHPOnZbRtVChu/l
hlum6owFYxuuZeE2iKTIK33IT+JwqZWjKQPQwRu9D5YH+5igrLujyAzm2rEI
kdq6E6qEw9/Xq26sYOFcqSWTLAyDVgZPvLGd8G+1emWaWKMxLhKmHE3Mo9TI
UO2BVoxhiKXqcXQhX6VhKGQ5wVxepiepjkK0xWiVW3nfF8R/7mkIulHoBUD8
DOlLOqKyX9cochiUHdz/eZqPwCyBmMxDmHlQrUJ122QAsmgilvEb6o0DXc0K
frKGlKDhkIlQIvYbu2H01UVSYGN2f7JiyWYnG7gaN6tG3bnUAwRQA0s3/3Ax
kHHd4Wmix0JvBHpCfEpTGUlc7vTx5NMimjZrv5qP/S32+mieRqcA/2Bkr6PZ
BSKUQNpIm8HgkdSVbkojMvPko2q+yu6MrYAh9U/qjtrNYaehGXJ0c7xkCMl3
EA/vM3S4KcpntsdKgyejff4Wg2zDSv0vjOzFbEPqanhvoGCajUEudqOM3hNR
m6oINBsgmCB6FHyTZzb9TSokUNVtwONt8TTy5QwkqiPKnIhkkeSFBrZ5ZkpR
bTfyLee0T6DsOljT30SINO65Qy+r53U2dSvT93C0hWNQBU9wlrxhixv0dayH
IXa4cXyENaI+WuWi3ZrYE+EhmEB5gEW41ssm6GNUkKFJ7xKfLMnzJUPVgjtR
7PamV4pgJyeOMqJaSxb61NdgqWMj6aq4AfievZbLcZtTIlZhMIjSw1/JpkK3
PbH4J6pg2aeRjv0NsO7nWQV9W+Jj09cwyYeO3+aOyQZm6rffwLiSEgg1GqxW
56MzCRG9JcZTUHJVKUmyPVc99gHTCHWUGr3Y/QvXqAv0RmoF2GC1GwyTg5aO
ULK4c3NShImsiwg1cUl1j/8AflK+l3ME83PTewJisRuOhQSqYczWmuiywKOI
KBCfIO0zVO5IA5YyMm69ApZ53br+YrlOAqxLxdmupPzx/o9syyyAd3EhlGZ9
eHXCOuxLE7f9335RhyfdXFNBvnYNgWJB4ExQ9+S1Vk67qF6NIT18ZEuILMcx
/e/2Jr73jJe2lzPNE5v4rNClWS2CqnXbJ9OJH7MCvMEj35mqpzuTEXVzvgJc
/7Xzid/ZyX18EkbJtwl13Qc1n4UJwlOQVrmM3lp+NYzJB4VlRbqRFMk+uPO/
EaFuAO5n73mf4uE0XJLqg4Gc2/TlCVJYkrhI/fVpoKisoq8ZKBiXGSGGW2yI
fpygKzb1GIo7Bz8am/rAy0jNzc/oBXdc/ChVBlnysFCU1UeX49kOytaDgx6+
5UyfBsBfRhP1Y0e59y5HfRizU9fNJn2L4FMhCpUO7IwQ5Ld/Pe/RB/yQoCWZ
gRxWdefx5wPn2MN6lDZ7+5nHsL/laEJhbJXydDb91LlrtefNpu5qCdfSYF9f
tTpsyifLyobXqPdCNp5ERatxD5+rdoAGdNpqTzlgtPtbr4zGABI8qaxyQARE
JVOBZ5NZ8EJcUVF0tXAD8S9u7jALnSKspD9D3fLIy6hp/A3nbbngZ9yR6Owe
/59Xq/pVAA/mzOh9bfzjj4IyoTwCXCnf60H4tQZ4/ZMaqudG+jKgBKkOJemF
pu+W8yY1XyDllX/V4uv55CXCcbWtGvXFvBZbETqM7h65EjKwklTZjOgW0DRZ
xV58DHqkkdiBGQ8/TULzlNCMq2bFRZQj3EuWtyx3g5iLzCbm3QrDoBCbvmWs
R0S3ICS1YXvRxk5h7SrBsIkIzRvqQnhFhjgJ2Kch4Q8mscSyND1ugnVEX8uK
+mBsJxDirUrnS4GpwYSElfgeiGIXUgvXhJyvcnniDmEHtZawUFJQ/0zOYPzQ
yGV87TG5mK9swCC+EYKPL0JZfAumwouUE2Mu56faVO5WS3NcQYADGujiP7xY
ftaZ+s7vwzVWOIKc2pN7xrYBTEW0oXqf55QD6S9cqbcYI0ueLtQvkhwcTZaO
v4AXX6erhxi9Ne2KgiV0EVAm9xQvhvYrTFB4H8uARrTF/QMf5Ol0S+CvGvA2
55bsXaUkNCAIHfrT9sIhI9lLcTFLWJjud/TLeG/0WoplYGuIOhxBm0VHT13I
/J9jVfl4AHUAWHdMmJTtqt0IPnlKGl27yuC/jofpnJrT7bP3+36Y0+0WlFn8
Q0C6ygtRlcTH9ICZDSdwcoxkeQM8JEoX+tsle8IkB4scekhc/90JCHzkFMEv
w7i9TybRuRqeGsZozQUlBKipupwPmWmy5g59CJxr/sZSOJ9ePo3l/ea1UqUB
zriJT1ecfiqqYkMx9Qr+D6Mx3ZVXalfwoxuHet+6zc63pz5DA4ve6jm6UJ5r
LIjYB5rbw+9IDPN2CWhP5ve7et7yFbN5ERGdEg57L+SBZBSP/H7QibFD8kNt
D+XDw6z1rltYbD/SAFkSA560GyEM4LJTp8og1cgmEkkvEiM5/6FoB5Eb0hyi
9zcqESZp737DvE7pkH2VRZjk3I/ysAOsTN5UlkeOIcXfUq29EsKbqDadG3mG
njiiHJtD2dU1ym9Pbk/9OJ1lDqgBBRtOw91Zfl5b4kNQWCKiIlUSuelykwy+
22F0iA482c8398SmNg/fAukurFKPnQam8m0ZIlS1g0sbuYUFhxVEWsah06Cu
ktD+vUI/4s8XcK6LJ3ZCjslGdNanpqHzebKAKaLsSZI6+knxHypDTDicJBDp
8iDOIZHAM81K8inbLJ+xavD61rSLlrYotc3+XNjcwKtH5TKNdOtbSTLqFXr4
0D0icO0UMb/oejW7ifdIFMZVudyLCOKzkjw0o1mda+IAxZNjhHKWsL8wRK5L
y4IcRm/LtQ06FxsjHSmjTuaa6ZgRAEcAD6orhDSqvl50fTQm0l5Hri1xKv7y
ElRdg8Utf6SBetaUd+G2NYKgk8Fzb7zoPKM5P03gCQQk/VYThPG7o9uy6tG9
c/LTDobaL69W3zi1m+gNmpZZNSi42YqtBJNsb65Z/riTzyo8VVCh+cOWEEo3
pZnVk1VS4Tneo5dpranahTUSzmMEQtfwxOpVAamFzBjngJIhASurBBrh4dHe
/iGY6qANqKtjnzamPjd16R5mvyWjBvlqcIVTSv8zhvR+iGziqBpox9GJOtqF
46XtQI6aENOfvFfv0LV04T51SmYNyCh5KblWwQKGUIemQZjA9k1OSpb2CpVs
E5Dccw+/Wc6Qred+mz3H/iS50exjICAaXbE1N186UjzoqTUP8/0PpszJLHOr
bx1HhsjhXlRd2Pml/aGc/ZfoSs13ISSWERM3k3ouPxTBPOVmRArGPtYJUghw
ZoThidvrJ0yXFUCb+eYuAgq+C3zPqCfxuRkaz5w5aYQCT/X/91UNgElCl0Qy
seEFu7I9aVestgf5Vjt5tRn5N3k1nOEmQs2cJHnGWJCDg502tqE+ZmVH1/Wb
FrZ+8ZUoNK0m0G7ZfSk4a7pPaPv191KCgkL5p3x28/cv0kouT7yCsnSSDOVo
ddlQTEViySKi38UMk1k2v28abO6zTQk0cdMepqyyoiBA0nYnLSKiZ/j31eBm
R7PjS1dfcLJTekZY0zz//hkucSh3KASkJBGu2i297ARGcw2PeEMACFMiyPN8
2M09P164vQ3CKkuWcje2qH74BLC8jBoIod7CQ1JnU1XFQRwWZK65daurZVjv
rvQIi9ZI6gpJLq6tkc6cu2zdy56gEMbtIvn9P7BIKWKTZgNKu5OsIgjJhE+/
+4jyZ6I+1W9jlRHWsvzHrX93e0vCEB3IN82u29bHJKy8ctE7PshBLqL76IgL
6lkksNtkpgiH2zeOcltOAclkQw4UlTQl5sys5G8RB3cFwYu7e3akbVyeuz18
gncWa4iTzslmvv8MbvU396DUj6Hwtjjwp/czp8xQ9DFPVCGX9OBOf9/YXSDf
dKW510uhwKBQV64nxIvFbFArfLt8pBC0RbiDnk1hTvObSXFmEJSO7hmwuvbM
C3AaAVGgDq0aRV/jUbPtiGAlFbQhrwdPnplr4ETGsESIuRTf0ZsLfJ1Jx66N
aQQHlVYC2jv3Wjejlzl/3x6TtA5kQt5KMrO5ZBaCI+nFqv/8437dHqNdG0/R
lCLgtxWa5u9bMT8ZSsX6aLAzdSjFWBP25qMf0EGKmFlZDtkKFPG1aYU1uRTC
obGnizEHGSEjt4PsCZOgjZfy6qTWo5AuT1NPy+Lz266WDORlp92ZQqxzjKnB
AOlLwGHV2C4sEGc9m0apFIYhx70ELGFLPvSzFwS3R4vBcVgQUpwM+kIU89aP
SBDtxPjTM5J/AFsMHCLFD0TXX/pfgk7/LRv5XN1743ghL4+P48ySf2cyn3xw
YzuwgzCpLxB3geJ9yCfn4zVL1ho8N8knKT3IoN527TcAfYO2TevGMLp5mDBE
8qKQRIfL9BrjQuagZOOyGGksaDefzEat8TxYFSrAvaVRtdjeRy871npxplLL
sAQSIsZSw2kpDgKMznmVr6DoU0ASxUn4hUIyP+OK4+t/d50zCnwyWW3DAhgW
hVsn7bK+r/s4vzEZyWtRXc2tWbvHYs0SZPh4M10CKtuNIqHivGHlOerAjeHp
XlISNQAL7NYov+W0gda7rxbdOpzmT2V039qv/nxbDTCp8Q67CULVsejgIViZ
JpatJoQ9Mj5d5bulAn8NM8W4viaXuKWwHY752VvPcekOiPDQDvI+Up8qNLFY
CB9vNvwJVcNzEdpnk50z8R/2YhKoHKrYAxxmBlzopd4eZDjmluHe5fGQ3k1r
LWkSQoVFnC0bidxUlwVGg3saCCvVKxqs9W0HQCF01CdO/L2rIACJPO182ZkP
7bNGtcFKMMuh97JK9jWi9/JJOz/wktJTwU9Cb+Fkne5S31WyTCDP8MmRDb75
iBC5ZqlohSGnXVD4r+/s8n2kc9iBANLTD4TtBTfSp5RVkggO9WE7sHr4fRLt
CHE9JpGJpDQsjInn0Wz/5MvxfHGcrPRRpqpg8SUwqZKPcBGg2eu/FNEibKR4
ueAMTCxQreAIKNWz0ffUdCqZNPuqklFsAlaJ5Je+gjJuc/OAEprUIPZj5VPi
dxg06OOfbf9QjLy1XKAz4jEngvIwnBXjv0HoqAWW2t7VZg0+XofrE2eZK9FW
Mun+9FFmT7qf9Gf8FJL9d/ygAToCTWB8Agx4ge368XX8cxSzyQoetB3MZKWv
F2T/HUf04vscLC12PDZiFGx4xDp3uosdemtvqVzVaF2ID4etz1kgGVVgSU82
27K4mQTgMLg3MbqwMu6jsobq33zB61IVy66G2RfjKQK2JbTuSKLjYs6O7C/t
cFR3bVG2Max3dgHrhjc14fZZiFBHvmpOqIDHa4+QFqLlzQ6k+mT3STX2vY9R
g1NH+LtZ/OuM6iFkibFk7tyKTXX5NDBF/ViXAs44KKuwuiQXYxetXOYUsOHT
xu83r6uZE9/hAesrA839n1FHAHE5GD90BEBYKGP6kr59/JJ5iubsW2D3zPot
/j3SkBZpZ0FOT22xsouKrMiienNrznLcT9XTfFpTuygtZCLEZ9p7A2oxkAPj
i1vcVOxVXHRHuQpiNi0KuyYCySLPFQeFeRWlz5lUaXJ2GkzZpAam+VTrOe0H
8QzwjdcBSfbu55IATNhvizFxEOr+hMNRNf6CwveWTVarOb1MsCKXf/rjJihS
4hoCFdk6hVqtmoSyDzoyk+J7lNRqyruwDF1fBBVLU61JMsN+P+ogbuIK9gNk
1QDjGM7yxa6+i8reY6rhaJ5zLPY4omEIEUfH+ve4NjqHFpZTh7is0Lnqlqdm
8k6D514RVndHsVnPsb0/8p0B8cCUhQwQ380fYkefKa7DRuDdQRJqp6A1Hku+
83PNiHZF7BCBhgZ9dDdzbdEt+SSdAMADoGOfIUj4TVqlWdeq0cqIcUAgiKya
wzcFPBZ6OoEaSxpit3J5W3kB+iVi5jzeoPueriiRGz7h7GDhFdF7AK2+R002
yw2uUStWfeSYVbvoAKoetyNa9BoZDExi/CDOlHOj9zTTsUKU8vwxfbZIUXAt
7g1QOa8KGd8VzpVt1xSmxpqHKTzbsocjhjrHqFoBBHkGOXavf5WF7QYAo0Wf
hfTIElwnCRkmh08RHymFyiGgZPmN5FZ3VuRV7D/prQyJQIGaVBu6XaJvmpMk
enYp4CiHUFrM7gL50IjYPGxBnu17KD1Hfh04i3vGIXeTpZUbsVYrDpP/XhLX
0jv0gx40fJF/iX3+o5jjnmUBC79EV99IhgWdJpX60/JvoOx/uKzzu/YCzf6G
PHZfyalOsheyUwPLxp/BiTreHl/KR2Oz5L/b7xCEyvdyATJELJZvu8gSyswV
R8a9olWkZAIl+9aZ0uR+3mZxpIixuZg/BDhzFmKEEa8O0JnvZF+cqV69HZHn
alFJ3EqBI0OHOzLMX7v9bsgb/Hrn4x6bC9b4hdTci3DIB2e+FS15/70smSTA
vvsWu4Pdxo0D9TaSZNBu9caJqichlUaT0YuKnFyV+0fa/wcYYslKSa/SphP4
Gfm9KB+5mFbN4jc//BoYD3QIeaZEKf65O9QjLlG8yLkl+CA2sTViAgGOSVtH
axuHo4Cy+k9KSJh48HzgPncV60Ow7ZUAGqKEjqucCnP4Kz9/PI9pnlsysbd1
bjAnHtQ3FVAM2LSRW2RvO6I/ohsZs4INkbYJZAZTc+1CasD1MRWeu9ZgcZsB
wHeMcLM8NccyiSuhWU43Sl7y3o+PTkMgUlCtytoWgjkHcQkbONXWYiaLREXa
OA9gsI2Vjr78RsYrFUI+PJefPLXTA3mPTal7QzbfNo9hx28CmyvXMKRh4vzT
7SmW0e2OKwQ/x65Bmf/j23UTVD8TAbf0UEYFnyHYHfTDYc6RLsoFOoNv/wVp
A1ix8SdEKbG3tJwZyc2g8hQ9NiLQKeO/OsfYDtIS2RYc5JwfzZDHR6X98B8g
2ZJ1NXkCPGxCoM077r7B4S4pK3RSnf/zdHEiYix4Xg0aMwQ4lKx5fJklDch9
NJgA8qN+dF/fFJRS5c+WKWeqvrisnspwpRLkBXyv4ccPi+kxmyz7uwl3TPXv
ATPTGNnbHV7//jpWFd/HrKEFmQAKdGOMAkquak1xEGX/ryS5KGn7EntbEsvO
q5pKNKmUYVeJuoTlRIJAjdgcsY9CGLpoS+eAZ8RrzY7JALjE1f8+G9Iz1OIN
IayFoeSdYjFXYFD20DDGZltyoeSp2Lf104liDsAHnn66qz9hc//316D4QlA3
hfJ5q360BVzJaR7tx8gYVXT/OooWS1jvxjavOCV6DORqnFTum1zYA0yLQIqt
T/stPaRZNXJTxBTDsjrokTUfUrIm0TdBGXRoR9xxxFppfaHBLy+Vbdaqexg0
g674GdtfohDqtlXJykq4488Gk7vZLtdKAh5r9H2+FL3jRAvPKgGRX2nK4IHs
Rlmi4LsSvNuXKnJrLKM9rMMVrOnxowJBuSZCOTpK1dp1NnfoUuEV3NYYNIBq
Xus13wdzg9QQ9qv8JMXxfur2byil0Dy8V3ojiI8XifvUKdzIDtA4tyucVomF
7hSSJzvSbhwUP4Q/UhWDhwCmMuWMvQJ7W0b0XZxNq8hfV6oMr7zJh+FKyRq6
kP6l177ZVnFVgLFMfsfEoAUJDPsnnuajb0AaaRp9VBTbl16/eJOVBxsP/sZx
LvfpEY4JVulGMLh9AgeDFTp/bZSl0fxbk1LV3ddeN432sdxFlQPx1sCAes6F
d2Y/EjCh+j3pSgqR0N2JEdsKKntJnD6sqPX+2Ra/WmlW0VVb8nREM/+qxIxx
Jw2DyD7Hxri+iAwIoNDlOQYie9rZhxiL6QbqrldxuGQGlyukkvpwFoK2H3rH
F6XVi68j5JmnD0XFF0hMlRPvycWaDs4Yh7ij0jRjg6BFHY2je8V1qn7Ej9pf
lfbODPfYlt991UT2jrtjdtkbGj6ZUSI3MAVNIF0D9u2+7A4nBU9X0N9al1/v
bAORF0TYdOeoygOciBKMABog0JuRx8y6yia9pQ/M+Y/omTp5vSZLmLmP2U5i
O5BVydiuoUhbZ1kd0lpYy3p2AJIDbA//pPQ5Cw8U9n4gCs3Ls24eoKeUXJ5w
23mA2Qq8vnwnDCTx9tYNb2gF58VAAOVVvEE05IVEMNRri9V7EavBFb+1LnTJ
HKImq2Dyn+cehD4GQGDenXfaV7uOoCDLa/ztIdp87fr9mXoIwhIkOaTKClIl
1OTu+R/d+Q5jlMjscYVqQt12TaHLHW1kdY2TxWDeWnQFyBYLwDWBco64fHkK
N7LVNA+pT4MArtPee9zmEZrFgZPACAgW8p/U8GetMMFifFNpvIHX90YgRHTc
ebBC/AD5I8rarRvwEyGhfHVsYPoXvlSTVA59RLgC8umORcOXCbua+2qO8KrZ
pJA3dZ/UkOt03Esy1TQqAD1eglmyOI2kOHBSuF7Foxc5o6U6tvJPSiD56a6j
89NTtxBzDy9FuPX59TOp3rUOdRfhogUkSR1nk9EBPMxMTQiAIPpq3YRWlQ0X
A8b3YWRSlPYAHmxVICDlR0PjLHZOVJwvP/H0LJTTZpY5shlQmZb7Hhup8L8j
1uJ+hO24ZoP2q+tG9WRQ83lNwA0lWWXdQB53VUj8qvOSQvgIVfeIGSXjO8Py
kJat/I5f9WjN08dADVvwPHnLBfsKj6TpXyMm2q5eTdBC3sWtPYo4YnRWQY7X
f1w1v6RMPsokSLCpjnTUkv8xWq/+sicpkLGAOuauJAag1tx29Q3oJUDuCpxb
VGwm4xZLyOngZPnez4XLUbNL4IYR1V9gT/72PExqr/fZIdgX7S4t8H3MJCCK
XuSHtYkdbKff3nAAQY/MmZea4+jiqFjhHuRMRAauKDNsSvZ1Sd6sTZv2+4QX
OQuZoQwZNGdNrzB+5P9SZptB+rB+EBH8YnLKz08+Y/biThiR2XeYOT9FAhqB
+eBIQWmfrN5VqoNE3g7RPkSfQ21RF2CT9NkBcXCMbq98qtJVFAEdQT+pNdu6
gyPKxCq3s9RYefYtj/TAM8fyscwm66MKUdSUsLnwHusf8Gpvryf8jeDS1E7D
3ZnvcstYZNeI0V3zRGvZJYrPdvZhzI2hEo+1s8DFvWY6aZRLSBqrhIEUGD4V
Wdgh7odP5rj0iyti3yR/us2krUpeLIOh4XhfSpvSuc6q8MHgooJIEHFjcRdF
oE2MdQOXUoB8cjYVDlK8Jf8RcbRvuI6+djGcRcXUC8DhhJzOF9cDZHKLs6mD
wP3YzcX1lGI2HcIwGDyrFvEqJ2Pf8YY1wile5rVR1Em88TyqCpn7s9+u295c
AXJyvutk/z7vMxtaV4GRZkq7w0sMIIwpXbe5ROrqppPhFtVqzKZqKuL8SZKr
sHZ0LwNYSjdPXXhv2Bug4c/7TBDyMGmpgvT9b1+4tSj1T8FXrJe4VxoJsfVe
Cyka+GUTyLCvEJzqr3e77onv+RCW8woO/ZFc72rfT1zs/izrkbXFon9XfHnW
HeCFXv6RqwBFPkCEQbpKMHSvugFFCJ1ugeNJkRbGMQioD2VovFoDvGwjsvgi
PNzNdhrV6gR1KHxnzqwgueEuOU2OnPN8M8BiXYDl7VEPClAzTxi3j2QKQLMt
wOe1pAxj2X4dtbe+SZN/CmAJ1j4ioOXxoOWrP0TCUyw9xLJrH12L42dVrr3Z
fGRW8GTqT47lqszNh0gp0k26Ss9UEN4hmirlQpsnYg7h3T0T5gWYFAQkRalW
cVR0muVU1vqiGpm3dKAAUu9ZKycTqMUXnNZ+8Oc4rAzSQi+QEKniiwTz2lnA
KONo4i6doTO+qRBCTX12wzsWZkR/GHRTqXIbZE0CCLL18CKJ73pYXajzY+0i
zoWF5xf8oLwgiqTBIhclqItuE8wmINIRUIulYVqUqdMV89ShDre9tGcuBgdB
117YWaILLqnCkeV+RptthNKcjfSceMrmRjX9Zsh3zmxqDNSDMKqKdoWTHIbX
cnHGisy89/HLHDAdr0v31oqh1AQmYQqoQd/RURvt3mxcSN7TTH2MgC/QrqGH
6RwVilEqUcfhnfpVLdBS3y3zrnHhYk/dxwdRBtR+xQSP9eW/WKePl4mJ30MW
lXUxv5Gu9WtevYvRvade8y1vj30K1YbLZiuoUNF9PiQxr6jwPo5o6hVVlTdc
UQ0LOcKs/qWCyz3N/z8R7PgX4Ry4BHTv7k0DbZiYI3VPTGHNwvgITUU2A/Tm
+8mPV8xyWNSlZekOKoq+07BCnGlBuGEYmQmiRUTKObRJ2l+bty3R7ccYAame
ZfjJhkq4TvzY8bJ0ufqYufj6WG0q/eXUwwYZNBzq+vUmDMBLUdScAu54RAh1
Q4oSnpoQFi0eE2LgcQR98gVwvHn6vCFQfOc1Zg3ayVl2CxyWWj/KuWTcttEm
R0qpS6Dr6eX8azpSb7/cz7rn5u9xnqOQ1Wr8AKqeYCyj47GvbnlHYik74pAs
PU4IwIaY4oR1KbG4ClyWToCFSOqMv5+VeFtW+4nqJLc+SO1tYRvDkvyb5bc0
Qb+oYeeQjMrZanKByb8wWy0at6Q+zpjqwe+wQvUEaiqpdXl0F1m2DxVzzx/V
AP7smTK6dhnkH8pryLlhEjlUVdEwP9YEttZ9Kcea5JJCCohCpUHgOruaTZV4
IVnMp1YplEOmT/+fuXZaD5yqs0XWEE2qraRLIAr7g9lGsNFSWFfl5aJzdYAv
oBtr/vF7p2GLvd2JROVKPeJZZIh/fFS2IHJn+XeuMJXPnzFopUJruogjZT4O
ndnVbmZaF9jRS3toeM2MqYcNPO7GbeHqq2ImAqGS8Y/kx8iOcrAgwlXt/BHu
2zflQ6hYMg3onkTJGigYlWFQHi/Z1Iu2+bEsyV3qrRWdqLGdVUqKouNntGVD
hL03ThwzmMPSdGtbIQgE2K4h2WIUtBs8IUle3l17qm12V/VxWXkd23/xT8fZ
62Y1+tKMU4yTexy/jjFoH3BFd4jFLl7q0aDAssGe7iMGFCy+j8ll4StO1jXS
swSYfTQkEtGT05k/uraeCn9We9zsWwCgnp6OfI7liFxdENZ6zoKKAWw1qBKd
08opsF0OMCC/z/GGuFe8D5VmwBPGk4OhAc+upAu62pvQo+IoNs1+Jdv5Fw/C
m4ZdSdxv4KJsQHTz4KAE92LNFja8OdSkRjoSIxzHEFcZidzLBhxOIG3Vwa5y
y0OwJUlcnrFuCeIuKhLvWfsXwSQSBWW37UcIXLt2smnTR6dzfkdCZSTWzNPQ
q/f6Pf9Fzf0LrDIaDBzp1LnVQdfWc3fEwSP4j1DO008xwR8kB3PPVD7xlVuz
G0Y17CFBqXbi7SdkhtamMHcv5zLnh5DTp+pBK2+pIZzCOtLh7ZqRxfKizwGl
C/nEvtBMqjcNXIjT7tvTrneDNXz6yqXc1WhBLIqXfflnEDHqQ4bOIMIFoaCv
gDAlUhtTqI0uPhmKobxho7ViYGcih0qazaWEbVtYo3JRU4Tutqk3iZCNKCog
iLiKG5zVHV6gUlTyPRq6BlGVHcYCAaVvQujsgkYCq+iMQKsUFKRZ4Cwyslf0
LwG5sA9rtPFCQFkxo9uE8Y8KGibuY+lzLB1sVyle47YZXw/Ge9vNSi1ysV1m
wxc3ix2BK0TaK39KByQf7NY7WS/CjNcaNytiSBNJwIbdRsuNWVyM9F3v1f0G
mvYO69kxDJlmbyt++Nw1OSynuQw+1zQtyrv8JndmHf/h4eHIVd5WutL53Axk
Kau1rTH2nxEHDtnU4N40h7Q9bOL+8lJxWn39nsPetVd9uJKcJTtlwppJ3JyB
u/21arkbc7YA1bJ9MeABgi6L7ipmnUdghtT/cq7OmXLfYSkq0Vaejq7SwBnR
nxXw73XP6SbaRQOBdCFetCh79ReePX937EEq+l2XLlxgl9j8py1pdmvACFlb
AJgScmqR+QFG6GTwYGIv34FLzYdQV8zOkwAN+jANoFCL6vD4ArnA0zOjwFcW
8RcJNZgGIowOWMWeLG9j4M1plFrs3HJm/wp/oKB8ah//X+oiIKZ7rl6zBSaI
0klzR58jF/aGzlbnb8wNmRF7Ou4HbBHgazQqnloE9CegZSdn555YxnO3M5oO
ZH7K1wNimS3Mv63GxY209pg9ITGkzYi9h1Gaz37imNLLz+cCcc37Rc1saFHy
OX8zhPA4OmYnLceDVsfbWL7u40J8TbhQwCSjA59ttyTWXzwFVf/A2VfWrElI
HcVp8w9kBTbdVUfHqA71VW9qmxekOE9TAJz4o4nbUKr0KmrBDgVFhKnxyn3n
AjMkcYIwEZBwbm7pY3+g6q+zlMplkpHgCdxx1+XmCLKu6d7YhfmpgkYQ/56u
kRxuW4ggS0fgu3Qd4v7nngTCYpboS0V2ULMo52btWsUBtvy0gSr4r8DshJz2
U1wuSLJ78P2SBYwsZRwGxllis4s67E+LNaUJz7LLzVMdgMU1+kn+HGOBZoqd
XFs9xqejXfKSPY4EoW35MIVNhsKDzbwGtjVRb6h9R2NO1x+tfQxVT5PkNBw8
JX5SUWDsl2LkV85HBpRzENa8CK5B37+Dje3NB7qosh8HegjCUBgRKeuGA3N9
19fyKSTatk5YdxdpFhHkENBuHCtsmMObitfbiQiWPgbWp8wzKaQDM1z6lr3L
l7xJ5Cp7jUlNYsgTU5c1NOreV13ES3iOvVx+MoqhOPMmIH3EX2niHHg/uPlI
kA2ODQyv9TtY7m4TP1+UuJTLY3iQfr9nSIJSCQq/4rhg6Bs4anJmpxG1fwpB
MVNuG+DaYjiagfKIjV0FoYIvsZlM+pyN6YYHgMLzyVPG8+AT/wvsjrSo5Hbv
JjytgTog9ZUrEd0UCLHMeGfMU17lbVCewjB3ofIxAkiv67W6bR8hV0otvMID
PUec3ea79mbHvxTKEzIKQcUg0x1ebPDC/fj6b+fOSJC/FxFyJtTaJ6DXtYQx
RIK5ktEKKNK1OV9wz5dtbJ7jXJCGzmkrkmrAgZr2k2y/Nuz26uziiAOIsiqI
mg7R+/iN4aRy/NdTrUt/G+corOqnUptkF70ZhF6qDq62/piNXoqmrP++xDt4
FZIe9+cOXBHN4xj9cfUn2q+M4YwRpOLl9uVDvsBEJM9JgUupr9lbzt0wpRmz
vc6iRI36fgtu0xmj9YyYlkZFZuCcn/BPS0Vuep5+pXq1TABsTq+hzLnybwgo
YQvKjyQ8tvNTZ3XE9TXQ4F4ke5l6efzw1Sgni9yf4eQLg+fbuDuz9d8gUDto
Lloc57ABgP5rBx85db6q+PZIY1/9p09JK4mAhn2wqnS5Pm718KBHsG12MoAj
nb/3QF4Ayn2V5rQlr/YISMVmY1W26RpVOsDN/kIXhqujAKhBrTTrzlA5ovQE
AgID7sZNphtCLwDn1kjVG/H/7cS6fPc7hu3jjYsBMJKo9xGAfxPLJcuMLKbh
+Z5QXs5YxGH60BKQUbb0gLubZMo0qLLILGvdZRrZiCeyM4P3hjkiz4CaJfHY
i05fOTmMfuODQ39UC0/HX29G6Lrn8YoOBpGpqzVLT4CuG3R+HhxnKPg+SIFU
qDV2HKbr4qgdgCD4aLcsJ/m1xvfiGQhxr0JmtFgWN0RuHL9jUw9hkoIgsBAn
GyCEEytgC3HplMBuyeoJ5CbL/fvq466e1oLgcxOFcUpru/lSVM8lJuHZhG0b
9i0oQt9Y1HiYE1v+bkHCVf/B9YJNjoX2tfqCoRMT1BX3byX7YYqclKQn37J3
B2vzrBzv7ryBaPiqZFXP9MY808pDNyjW6lBjesv2rvCY2wXWxARTqtlhzHAh
6LAKT5O70/XNd5BCwAzEH5Z822rSj6KnP7akt/T+dh7Ubg2i3hFyavlcXEZp
TC2gXChSUjZnHyAFNBMtjz6LZQF5dVmv8+8prTS+MKEygkI6AtpAeoZGCFR1
06F538z6AhPAkjce4LiVgRC8khHg49KDs16u9/cCwc7cPPmqtTSiATz6ivJw
9XzpibmtacmiopWa6LcC1fziwXYkheA0UXlGDDMOutxopIcsHkakQ2N/NnPD
6LqbRFTpYEN/l3v8Vbdz6kODwUALWTe9seVG8JjX/fhiF8FEZ3JD3XWh1VWJ
2LnJCT9BwZBXFyrRiy5qnZlhPWLENEOG72bQ4eeI5nA1d/nBij7ZjJxg55m8
GVwI4thWDpinHJ20q9Y7jjSvFC7zj6OASknGfyxqHl+OLuNOHJ8HljOiu66z
Qa4KseMLDcvq6p34Bo+ZYNbXZBUqnRsbnrdrjdC2Jj11RwWjxUsxbPoBpwJs
u1zJ/YmR2geiaqHy15bu8ndJ+ePWBWpD5YVtUVo8zjHBog+BgKbpN0efa2zW
9s3yEuaBUlB6WonJvhw9hVj2dXAALPIqapwCMVSpm/rOFPlSmZFFqmGYMoxl
tzJWcD7vz06Fi1zsQPIMa1T0AbfEGABDdRACAhtfw3bFDsT7Vata31AJnx0f
tiNA3J1Z0X9hmwxr8yZegIJUsGGICUZwdDZ0Vdm2aNP2c1t+JuIkRDqkFQwH
v49AXC2zdOR5QbCrggofeZ19I9mfpersYi1Z8juNp3Bz3jJUIFRPbyI1vDD/
t3Ao4r8PrTWCHgmGvkLILBl0yCVyegQlSIaDUWTx5Ti2+18RUFaVhoxXGk6X
aA5zG0MCsjCzmjHRpBBkkBp+nNhLfNBq+LBER3fh0WDBzgGIPlU3CPGdZFBG
vLaQuRN3XTRNAQTE9WXcoxNUlcVLHMkqlakIn5kOv30+fDhxRAnwnMFPRmJT
kRn2Q0DangFfCEtmu4fHXyPiDfrUnUYJd+zQBfoX+eWADMxUYyYfMeivZ1Gw
WIzBpImdNTD65tycD17rGPEWGLBispQC32fQAOHAlffi5T+L0vUlFR0Ne1Oe
K8IzddFKrpqHe9srz6wWIaBC0ZS3V8t1IhpDZHqQXBbDXU2kAhkmKG1xsXfo
w5nxruB4N3uE0G2HqUk+IyAs8fhOy9wWLZ68ZEmEbF/noDVn/B43yu2SqtgF
HR8yhO4cTQsKL4oLS9pyCsC37ppirBctz0K8oozfPoFFNV8wQ7r77S91nSSU
qyQr+gNjyDm6fVMfqKfgjU6YxDHXwcybEo/JPfqueueuK04wwiFLuBgz1ZBL
ZvVFZWIeYyVJWF2U51EEBlnR9ivsEAgY62OXTP166j0R7vvSapyKrkhS9O8P
/nWxi+ehmHQ2HqygcXH2Fo6E4fqM5HRkXXV5FENBAEhVisKR5xRjXKXWQYWn
BeX8oi59quz3qW+PczSP4nZqcRlsV3P7YSPjlXwCRGwWAv7yL9ATQ21/Z3lL
snJcSnQDpVUfWemPRtjkDCwh95TZ6X0L4qGUChBb7cGdPh5cGrKXdTXYCbwt
8fWcPXbK0fZpRdtnvn22CKZpLB8lBY/ogCn/xQdPq7O+hTAVcyZR0IRc9LBu
QZqZgqkuUOg5Cq6+VF+EprpuC2+3myTBijGjUteqEMccZX8zP0LSGegaO0Oh
9jX01xNMLx/EIth1BdK7UaSw9ySx/epOj2mX7pisI2QI1wJyAZoDSrBLLQm6
Fk60xO7J/bK9AvxiocgJ3Ua9549I1e/r1SiMRdm5CfkTAJE9dsvlf6n8LHrG
D9klPDNqDcT08zlEq6mn7Jb7aCFbeiOrJ1KqeGmJEjms5NF/Z9dk5gyiI0Pq
o9p90sk25m+A0V42C8mzyX2HDeIRyva+rj4+7DuRmsRoxl5CsxdyEAXIy6Dl
NzeQXRzoi0lzYnUqZwb4eB0Hyt/TC7RxMDClFpkmILbIutd67mJ7Q9KKxNWh
2X7WQ3qthZnqjT07czrN3LJR7tnRddm2mFkweyVy9N4+/a6Z9AfDpqHbyfIm
3V2vxOOict75cEo47nG7nF748kW7pvHlvO7NDw+N+9ay1O8gPWyd10WDnLrl
HcqqI8X/OR1Q95IkZhu9aj8xCl64CdA3byEtGUHd0N5LWwvB+KAi/o4ZcxyN
wPzJpGzgoxOTsArlVN1rAWisHaHnPKpROUAR6UN1HCtUXuNNcy8Kym3zkaUk
zos+R8dFmeUNoLj7esWts2ApWVy9PxnlmEYmY3y+wue3MO31d31LV3cucl1k
6eDok86zvh/arWdfr75+aQ0R3vQxZS0kJdVEcR9pHZABsCjHgw/prpyPlv8z
KkJXbFTiYFAuR9rlSi2pW0Phy5T4SluV8s0c4Va4nWExrIm0OEq6dImKwFPB
nJmIfmiwQetgZFYGYxkPtY07P1AsXLnpQah6533kNUnqsp4S5G+QqMnhyVlG
X+wlU/i8S13UdofJM23TDNVgG7WIduR6cLpsyV1TECcq4CfZfWYizfqkBVzH
KOLHqXBNJZpswXPV2qcgldL7W3CwLamtos/cLwS1R1AwRUONwOjhDqaCzT97
jXZ4+TsPQASgX30T6UYOYlS8JxOu0vj2w7g8WUHNHBUpCRmDdUMZ4N76ew06
I0Sjg5h2bvIQCWW3hXSFRE0D/WULplb3+SZGfLMsiBePPEnGpl8RPHHk8V3a
P1PzCugPut39AXVe9Z2uvVgQzQBrHCURaOdLE7eD0xG4z/X/zVgQdhSbrR1Q
3ZogY6I9fpQQptpIBV2EWpiP3+/h7PcMNc3Z2JG3WrQzEN8OGHxTRzRcHAxw
WRKny1DEk99Jj+sFwNVbN2m9R7Q0aIOAvebiSLj9Pg+jxjUXEgVR2P72yJTj
UA+iQP3LQA5PTiFBXNjHXQJZmC3uJ9ktW+FCOOlFC4Vqlxsbxnyexl1I/+sY
TorY106u9Dl4Ca5DG5/bf87F9ap81A/sORbw2QestgWfQIxHltcVkN1+uDDM
kDN70dBBzEy11a25q6g/Ztnmwv/QYhXtJeUOq2UkFjNVwdKFffrFTqvdg8Ao
tVOltKoJe6FachMW7RNMqIgc7E48+QFp6NIQ6sb7rXtcBDhhejlwL7zXiiDh
X8UjwQS4+QD2aizW53/UDikXgxOwMq3CwpAr8jeWS/rPzIJdW55you2ZAvFk
Vw4wNdM1mYZL/eANV9XQ6I4uKQGheGq+Fwbkv5ryzvYs4LsYYg3lTDD1Hzx5
2DrHkRjFrqpFOSn8EWwY3g8IJQDAdKt82MkygisRZgQwAi2JzXf7NCfg/X/L
ZFcIgyJ59kNNGev6cG6dSjTE0N1DC00yBTNpSH8cd6wM0AQo3kW6gO/qJm5v
BdQeXqxY1XeIS0x0d+XcLjA3gsa3cMcX3NioLmj262rKj+QwGQFLbkYs4Vqq
CC3ycGtQmo4y+/rCLNlkoto8UVBDgB4mKDeu6GWvLitsiGPIQ6WE1mB6TqGA
pZuKvfEFeKV5PJ0Z1G9ptF30TgUHU/sNmUURdLcnYg5EO9t/WkOvRLK5nwTk
1hoU7FoMuBbTQvKp0q+jICapHF/Vtdu0ALAisOlA4/mZsmuOUT95DeaGIapD
iMr0QUWO5khv6d2V0nb2AyeRxIiDRkRPSDTFVNvtGYU8rLOGGwiTlEakuPrk
5hDz6ZT1YtrmO4FApmDMBS3+M3UAK1BnO1XlW9BWCg++oeEaStcSUeV2KMtz
+Kv1kCe8jJWbSYLdhk/mm2d216qLX+sYmV7WuMx/nabq6ENuYHGwnKanFrup
n+9Fm9obn6/gBZ6KTogGbnud7RqI7OIpuZAY++mB6o8PNuLdY345dVGbD6NY
bekYAZMnp15kpAT21E9UUNK9rDnKLza9Gr4105t+dYeBodal47xp1siiPe6M
kNlJqQSa7Z2vZXyWRqSC7yuxp25iY9IqdNkYJhGg80wcs7SwefPM4qO9NL5P
UO2JPNQA8pKPiXT6HULdR8PFiDlXF9G2kQ3bfoE00ytnmr8S0PDXo88bPvjU
zzO6WFQaCvJ4qOTlsSxYzgr19fpr8IeChjJRh77CrKJFBvjikulfIkcHCSOn
+085N8nUc9tQMHPrEHxhxrsXoTav6ahuNrkGWdh2+eKUjYkm8raCDo//kVJx
o4zE/ChnTYIhU/hRsPGVCcRt0ScidNwG8X7Bp8A6GtieumOlre9EqiFcWnLn
Pi7lh3LwYFqY52UOAVotvgfMrCEHM8eeLeM0Qv2Rkzlb/itk4JMGnXyFkc9F
stWr1fQYejYlIT4IsNOQxNlRPk2XKDrAjd/nlX16BuitUennDiZxAv1xSn4J
jnrWcmTOQkqwEWBriX/Vq/UeiPBKeKLv/75MWfDi5jxN1+Uo8hauPYgeNvuI
c4fl/NctsBndBFSTUILJvfRVkpRiYhLuIBui3gh6Gsadp2E2wh0gOIBHX+Nq
B2Rp/XpJFRRfFaOQ3wCRzH2by5C37RM4lq2ABJyX1kbD+ENcVzGn/wOPsUZO
Nv4ssxVMHVBk0UXiGKEhg41KfaMAQ63EbpQ0ZHc1DtzvQkDAuIryW8zxNWnF
urMFrTpEo8aSyeV9HFKKfz1BwwoNdq7IeLjtZH37nPuOVVozIRM1N/XMKqfc
RyZHtv3yk4KZWKUXQco8M7DupPt+HyGOnVtzYDZ25Wgq0YXTxT99bctvPDcF
w3wLFzXc9uy5fjawuOWUl+LYWqlc9ABIPvTMElDOhdHQBN07sQEU9HF5Apm5
rwUVpyQqftad2zvNvD+He1NN6R6eGAhKWlHV5cHnHKLGNxB4bTaEgGGPwsQA
RNkpP3y1PqSr/JM0bpzvGLWzX2vpG8BTD2HfYxtZ9LLZdPyc3bBxhSesQl2T
bj4xprJWcqsrtqtYy8ZrNfh09SExfAi958bwj8NqUW+d5Ta/LS+rLplRXBs8
r9Yd+2Gbtv0DZCn+Jsq/SFQ5KDSOz6fr8hlBPLQEARA4eNjiDI5PPGGUQmyA
yojsx9PTnbl2I8GlhFg1Xp4u6I51wEIA7Ic82yPhdHZ0KfjPjF0GbXZu8MaV
I5KWX6aw8+p0SckSq3Ds3+d+IzOPwFiVlPrk/kU9MzHeu1ExMVDtlKUUROOI
oG+PW/TdB7Itvhv7IE2unaB1g0SaT4pcI6gXZqoH1I56T+tCSxxR0SDE5EjS
FkWKPZxH7hKcuDGDg/q4TZlPKRMJ7SJh4yY9e0KrSz4C1KQmVnl2+GP2rRmC
zUaXcgpECAZ3nJ2S4f3D9Lzhuc2WCCLL2H39zdxQ8MdrhTyG9wA2PNh1Hnff
Czm4Q/HLGHFhjrvSh7lvLhgKXjA6T08oQkUW2+ZGtokZoaA/bpm8YHmT4GQL
OTDL0jKdGUkvpZDjnTp4F5UjaiLXOGw5C3YKDRA9xTqR6WmdX0PBCFvJC5x0
j2TLu7AUV5AYk/BloXv49JQoOUWNMppWJR4s0y/iEroVy8OE+5Z1LYmiGtRi
OfwuXoT0xw7rVLOaqVK3L9bnVghcj68YCKTwRlgrG3tLIF2SooTI6a0h6x/V
fM8XKGfqnnhTaouQwF7+nExRH9IuPVPZdoNWwfAWEPuNV3PdKM6czsgYYYJ1
pCt6kGX++kzrQHET6zDTwpvREGTWa3zlwiPyhndTetW2W6gvjXiPwIAL2cI9
TJaU1P1Eg5AhFxGoak5GV3Xir22exGgTPt0njToCIb8OXg1Uc0reJ958dapl
RRPQr5B2bzLfhmUbJwGG4i0gJnAjigp5eYtfcpCX0/+pNVRILdxmPsnz9KaX
Fhj18Gv2h1prnufCRM0erw+SI/0036GTsRVqIqMt720dNtt/ZVdIEyJe6PWU
ir47mIcnYMLVCdNO4xiu8v9QJsDPlaKpMb7ZS7xvIbFXL21lhOC9Mzn/Un/1
Z6L3k2pRSK1Fyp2g3VUJr3pqIAMZgCuuPhWU7VCHEBVvpGY2Cvb1m7fhN+XN
KpADDHXQAxYeWqfju0I7v4DSqU5+LnVm65NTdxD+Whi4W8A3tT/01a4klqm/
pvAFQ4TWZPlbe1OoTRmickMmA0d1kbUKRsfX5hpCdy+iQ6gG/e+YA+dkli9H
Jtz22yzU0POp3vDFC0YOuap1sqyprHV9reWdvOlDLDXt1bazHzVvGbGfm3jH
D+Zaa2EqU438brl39rbyHghmmNHVMbASM/LdI4XqEkTXkd+ZSStj+jzXd5P0
oGRdcBY/w9Mcy5Hpgbu4TihwpaSTrr/Eh4AkXWNIX0thdJ+zevX3onetGzfy
mZAzfNorE59cx/LO9Dl+iOPNlpe9ti0m5sR/r60g+JA7hdvwSROD9VMFV0lP
A3n5Aoi761OjI+YCR2MVc7bYiECb6DuGmqwUw/WXGDpcK7QkicllxDhZu8kr
MejPpBd07MuBEwTcUQ/sYFVNcWFcnaPu3kV4Q+bDE+iP9eHFVbtZ0s8FNn2H
YJS5GctgEbqZZddQhlron6nrHjUwFwOEciD6N0TbY3pejPj7E8bkkSTXQyGJ
uPAieP+/1nQqNwtsD1D6PLBIYmc1s2ekQocFCDjX7NKbcAaOo0BYnYFBh299
/uXsjx1zxZaEZrLTT7Kpwbdhn+ws9kK1043PNQNzO5HtZsVS9fjSsu7FTr3e
y49Z7TVWMaVwipRMGuTSwXu3wAn1xDHWDFRPle0IGP3+SYksnkWlS446vDnF
umnEIcIbmXMI0O0fOrBMTroZq9gGZ8I/n2RfZipULHMN/sV32KLOk3j6oaJK
0bHuV2wvwhHDHCoQgbGyYXuxKNmI0cWGgprxUZ+SBqO7t0duZQEyaFX5qSpT
lKW1ggZL3AHe3Zf+UFDj2C57H9NoPabk0pW/mHAyjy1ny8y5G1474rW4rhbY
e3GVeixrnh+Ozr+mIPb5BW9SS2didcAvhJdESKwmX3FMMpzX68fjOqSK6RfI
3Q/mIRBKIBLormUTbPpExPjkH/SaQWwgnPTW2lQUPivMXksB5sHHTyzgdz09
1EXRrTbM1UhCbnXxKjm/7Nw/DB9yFKH2jNXYTunbtxiju5fTtrDqWPzd9KKo
O+zHHkJVbzKRlb3r8x2DOsrhp2DHVz3NQopi4kmUEnPMIpJlhwMS2TciXEzb
YGAuaUY672917CbyeIu1vPDoF6+Cw6yn7CEUPVc/xO45bwU5isfW+mJFpR1u
6IUvnGHA8NL4Ylsa4YEmM4QkT2ceMoPra7UMvc5i+wJTNydKQs6UwgVajLbn
mhiUad8ydchvBm6cRyHdeeUUMxDMytehur5/KyNB53TEH0Kk4QJt72sUYVZp
hKEvF+cUB4e1f8S1hI21ULokdo4hprwyPhnDYG7BQxpfN7MlqQdkjgm+MEwi
5pfkVyGFzBkkSnXTnkB8f2d0uuA9yNPKMpq0WcDpU8ZdZPP49k0YZ0Tyl4tN
/qnYBV2QDGTq/p16Qa22bvQqgrE+d+rL4WtPIs3VbeZAyhBjesbEsPlH8/N0
Nxp7qQh2bBLwYIiQTFg1gcO9vftSuKipjEfj7BrFBQqeWu6d7IjVtDV8sp+6
cHhrq885CnJwOtawjH7TawqXdKWhxKRdIIuxbebmD0YigSyzabBlCjzWs+Xe
XwpXmLv0X2UZrMlHmVWcxmA55vJoaq34tD+4hPuBIHAqbPvh1XRj6wDSjVdN
T78m8YGaejbFSQI1Ctv/TY6pbuIFfYKoWglCDfZgdeBz1iTWx4YS0ZFepIv5
7RqHM3L35JyYpUpxwEsAjvaUrsJnZK8x4SBBQh9W7mkXwQTMoWNdjGZMEdUZ
f0buFAnYnNZUKvbW3IDCFfOWHXa6W+ICBgdCMWWLexO7Exnq31WGlVc7ktOz
GPWoI+CTY8GonXM0Ch57XldtE5oOrIRdTBb14BzK3Kl7uoqvr1GNG69tNX2e
LWZr1LoWFG+8CTXwPwdkcDVmJzEteZvTLkKUHZ/gOIvlyUTfNbuv+GoAzoJ8
v69smI/kK7MzdFGcjV51Hfh/OLMGgJE8tdRXjeO9GMycKIYvVLHP20pctj4+
Qi33rsYCa7/SxWKuSZAjqjGGS9rvK7Kju5gZ2SvHSOVBEGl692kLR2mt1PID
Z60IkeEaBK9Bj0uIOeTyaAj9aXnK46/qLCexrs12dC5yX/BGdOiFAkZzi0QC
+mWA9cxpGoAHMhSD1RJyeeuErDA37rZxhzxmi+O2GHWSWe/k8vO9ZlLxwgxl
EfTvPhsksXw+Ygw+ZIJItrjjL5ZsCbD21N0+8UD2nlfnmt/Xyh3EaVKI/9du
qbpE+qBrY0U7qtTjxnNlH3TcjpHVy1G4R+r0KDk/TKDRXsLJIpxhVhXUPPlj
Pbgs2W+2Hf/ikjthLKccSIo3l4KvOyfn3/i08VAUIGZ2ndfr5KWnaEICy9ky
52ii9VSVd6gumJwRPwwcsuIS6ePW0tOEq3S0PQ0rVF3DX1lzBgKwNTTL2b6l
nkQu6UsOq4N9NZFEQ+Oh+rcaUY1cu48xZ17OIXZLv2PIMgtoO2JysOL9oB9B
EFGaJs/SUSMXbopqCe7oK/ZB+59JzH1SJuYMrtsYfxs82BccIgh/q9B3FUx8
jQRvaTiTwcLQgWa98wBavi4ZEy2TB3jECA0DAN3Kc6MPcjyqzSZczfA6DQbH
f5bCTI1eM0kla1kWx47IINb+O0SDLduHDiRu+HYK0TDLofnHpPaz+ABTyR1R
k9mNS2AZqVoFVkhZH6hNpYAGactefCUhRrmmluRyge0XAzwDwMS6a9IT9YRy
i21N7ZVXAqCfnagrP1o0LNsrVT9HmelbNgEgOmeLDZQ6pIBzHqR/66L2sL1G
9qA2QyX/I78nthr13jcnghZkAqk76Ez6dazG1V2/UJgLqcyt/hSUj9s0+/Bw
X0a+O5MKwFHHEKpvLux1iyoVzqwPHJF4jqFUKGuCl3chXMfLKzrGbugiEXni
iO22397vpViTwOM/8fBBdC9KFT6b9yJ40Cs7oksc1ieTYCcB04k+khiWN5rJ
KLZ+4en+UH0zTFrkD4rWrjZE056LyQWXh0gadNAAkMRdeaMAnbUidcmMp3y3
wAHUmkPLGGcQIhYLiFyqCirr8Tw/h71tfRCKdS9YN+y9uvy20srPrQOzVvYI
TKd+fw6DAvnMnHg1xHBLAsSxw754lgk7WumOIgYdsFpq00uxgtYq9Be3LRQ1
lAHZg8MyZd7NwZ4TrJqNzXEg1DmJFvWABWcQQT66re+J/zVxBM2C6Y6xaMeh
fRbTfyFyUPAcPdZvFjbzIKePhKkYTD0qHzACjN+NwvPxvayYD5Kw8Am1U1YQ
s6PscO17IWUMEL6AndjUw36hKAUYowCwhgwrCHMkr9pHCrYFGi3A1tJsc78q
+/1c8mFvTmp6m06eGCAEBQWBBHIL8RxFOyCjWNGFA4UZg0PUnJSs31J5LXxE
FNiq+P1Zf7NijRlDAKlAsvGYi+hTIlUCI4RGkNJy2yp5uHTS2HwLFaZpPxzY
4gQSilJRhQBAfeHyQgULpruBjPJTZNKtOwt8UEYs9/m+QBcFm9i+QCJh+qjA
yXFfNQzBnFstGl4I3cQj274H2/cs93fkA8AIYh9bolclLkdN0k7h5Tu9uGDV
MspSXsNx3ZAu6inGvwEM/0uHRLJkiWny+5LLugc5+c76dYsHmXB+VkgtZzDt
DSoiEWT3o/yZULY8XVqlOMv4v38iMONi70JeRrmjcCh1e7Z/7HrVk43bJvlF
RQfPJYIASKaRYQbw6QgU/xycE0AjyNBTac6uhV1ba25IZ9/uw6CjOyUra0zQ
MW5edearX+GAbcesydNWTGroV0ErSBH5wtH9UAEb6HRJ6oy4DeLsEt6emkUT
7uXyR6HV/o3yAg4m0g0T2IN38a0KK61nxTGShwAVKrre0fStP0NzrWujmlbj
ElCEhrAQoxmKJlBUcdzS4cG6/HOe7KuIz9xxjP+Jc8Vl3l3OLbXlpenCe5u+
Bap5ic2pF9Qj6r0HwMKKttdTK1S+mDDNQZ6x55HFu4zhpIQ83yxKTash8N0L
csW8SR0WtXEORqXfINAhLmJUFO0ZxzFYcQaDVPG+IXRj/WFXJZ/gpDQocNBG
wO4QbM3jCgYAZKUPaqOWl4h1KiMqeE35Y9usbs64eQbSRXo0yOTZpLktyu8O
oYSvpaiQfDnKe5lrYJ64Z5uitciXl9qNS1yPsT8+1YJK4+zNFIXGkaVaAzdK
+axvgN0DnWDQqNiShak1Is10pNRVPqMXq4Ap/atTBtGLxGcaA/KnwZx6M78D
mgWwgfio7YSTvx3lQHcz6dMyePUYCDtdpuZq95O9YsiAk+WUZbgv0Xy7Rgnx
e2kIuCD62q4vBu5YELwiTtMiN2tQ3dSVHNjKFPDzYzTBdp3FresSpoImAtgQ
hG1jmVOfRrBPwX3wUoO+XrzmBEkj54mIa24x71iJrtwlQVry0pjNrqP0T9Ld
ZTDfRkbWQ2gecZATuGylQDB+KhIoJCFXUe9flBMXEC8zVHsw2lH/FBGEPzfb
s5GS7bdhzGr46QDdCnB/ce1bQs3MOJqeP9UPMZQjdVxMtuPIPtBUgEX+OLCs
KD3+BXYYTgqM+6d/QUSzIHkpnMcMLhAzt/1oh18FLqM56khTtdIp+4aZdbAC
Jc/yrzPZDLM7NYnyQBOirXoUItfjTX4/1Xm0txTvzHyodRSh12O4E90cr2Nc
zM9CqAYt8bcPI+9KQpTH4i+KnfpQ8uLzB0dZ4iwxJuaQuMX9y+XhTuuuIBgt
GaC+QXzwEIq8DHcUoxfN/l1JN8C5S5ZJl7M61XChpL9a+5kANrNh5rBawRii
nnDjxdvboib60zZqHFaz+kpLz4tBaUHkroU/V38licJ5H6a8nauuKTKtO8Js
5GZse37EPGWGL1cPuHiwzDTrYqnT5gjAjuujmTaw/91W7YnkmPd9L5frGVgs
O6pYapTV6l4nbSkbqvq9jq7i4Wx6fZn3QG+zPb32BdKL2MSREvnBuyGwtxsu
MGNR4b6NE9WqOan5luLxhnzHlJyMbnKRpG4fVk4Tm3M7arfZa7w++N4qm/So
1cDMeD0qkxADD4DV/y05CxqDYmulRQAiU064DJ9Dzkdrri/uCz+WS0Bm9B0c
KHscGrLmS/iSbhDOJ8IyQxj5aMR4WCb1JqtqfLa9+jA9CLbQa0/SMLm9EjHN
jsvKpisGd1FHNHjYao+bEOFBp+hyVfvVvN28af0izan6Z171bvMx5eWyiUSe
THFYpDap/J9E2VYGU0jdd5Gs81qqJfXD+j2GpsRpdH2WWeKXjGDsKkJM0yq7
/7G6AEK73n3yqhmuB0tAVhIKlCCDrWEfQQcpFnqKaD296cODIYN8W6PaiGGU
St56czZAFIArWuRH7VRAlRH/2YTOtJBvcd2dpGUymToV6yo3MIX2erzbbOqP
NJTX7KenGQRJPVTF4xupcNC6DpZApIfoJtdZbAC86gVk+AY4qBgwcbPNzhpr
El50PEk+ZJlhvjhwn/4MEoj3M9uSGs371cAhajzM9TgT2SM20K3x9OIWvFqd
QFLKMJmqlDnAr2BGE21XCwcT1ZypAHdof3aRT3skkdKyW+fLkHfOopVuAynx
52LtAL9Kb+W/b0H5osYAuKNRxeYPJ84vmvCu1KUuiFXoDQJ0PFW3jDazdSxV
Kum9lhBwLhOJbJCMCvdrj1CivWEBVqcUlNI1+8xNaELrNc69QD38EgmG8cLx
NXm3WI1YCBkq2rMwjE9CB56wks2+niQlSqcvBNQHDCKLTeJcGixQW0bnSVqO
00RcNMZ4epMWhw/zEMrzKI7BHUNMFadMCLT3zcgfLVV94pGtekhwnYhsbNh4
9jBmYPlHd0hvt/ELz91KELBANBxQvPaC+8hRPxvqMJluxqoNeVpEENRLA/mi
T4umlMK/rmkpwgy7N7ithN0plcoBA61ZZAQo8+9ZuUtEWMJNDE35u0uV3TsL
xczlZ1Rd6Tiin5WXAw2il2OAqZ7CBr4Ie++5cMouVXqq2kR+EYameGmRraBq
/azANDpqpPNqLM2cB0G99TIrnVNEcyYJ+mDTM3IOHIsAlN4kPi2NkKjcyegf
FvCsad+5uTubbuc0b4MzSsGvfhr4r2hX1y1XBol44VkJL8G2/7lz7/Y1xNT0
cBDzULIm5vQ+anH4D72tYvLSLA69ZBEZU36iYmmch62AN51Hdl9rHzuT5gzG
gaEw3I5XxZFegheI091hNkKcjLn4yM1v9l8sOHlggDWs+j1e3oOVnE6ZGULh
iP6FrpvMpEKLcgpQap1Q3SRNkEYe+YAPzeNQ4Y3uVgprv9nzkOMRa8a5Fj8y
FvYL4DuMH+XEGnZWuSIqZJNFlQ6EY+F/WQY9JmDlNMMcXnQS8OORws4f4HTj
h2OQhAsOkolqP58hsIimaWU/diHyz9QDj7yYgWTuj0wKu3+Dh39x/ZtYT50O
wu/7rxHgx7bzU8JAz9mj0+9ZuZA5RVd1vPsAYFYBQ/WSH3Rhzn9YlZbdudyN
jkev11FD4iZ3p5AcW+5VVNuFBaHJmHofvV0ATl7pGJcVkuTKhjmKnkVtmtKo
LxhtjZN0mwq05h12eKEWAmChGh03LS6OrwZHG2m3Gtbeit1ZujCg5xs+4YwK
br4io9VQ0RIIepCIKmQkfGYcBl4nAaLl30+Ly8fF36qQqQMUPKSRjks2WFRC
aMwVer1ZbtSJKX8jsTcgKmlbiNeSBQVHxZGpi1qs8zvDV1KfxSJyUtoABS0j
sBjqMKTUq2tuRVy0rrw6k4qpyKvBcYuWbJqwQxuCs861Yyk+oH2eKikmTlAx
l8DB2vxgB7keIZ279+ksAlwC+Y34hKkI/mqk8N+YjHgvLPxERW5WA1GOxDdZ
mQV7TQGSB02vqlPQRzBc3dWUl2EGFbudeb0peiquKpyQB6fSyoRDekmKKkLT
aBpFAxxbNLnaHoNlZdjvrxoxf1Fz0JcSIDQpTtN+o1oFCepT8Rtgbq5tSOlv
YSDtn9j+gaMpXgsDsxMdVKORut86gWL3QRddeHmM8WGYKmF8j6GZ2Z5dXRR9
AQSwmGABKJoih+7gVDJMPZrgr9SLdEM8a2U+uwjhjdsK/hWsyau7q1IKjt06
451qBWH93D/iLwUBSrKKXMdfdk1TrU8DBvuMxrGucWt/6a0HUToektbM26nC
dODj2CIbQoYLMbr2/qhMnhk9yIuSrmFPEfo074IKHyxwfuHS8WC0hHrqjr/h
qw31Uq78NQapCwIq9jOalQTlGqB34dSggQ4ax6W/WwUf2M9LXB6rHxIoAMYR
aFjwwov7Xh1RvgwduthbOJB209QKwOP/PyutHy45FfCP2CMOtDxepZNDAR7E
Udq3ssGXVNOqKu0ur8kclNMdVk+BHh8gG2aazpa09bOlePBDArfxCcfnaf5r
vnCg5fdDZcN0Lp+ox0XmowylKMQjyoz9st/a+ZOu14yxs8Oel+Gpg4Np1Mh5
lwxhbEjIEQ6CCdeQlwjItf7BO9eXIzDAAOSpRnYuHFYC+kGlRO/vvQEpwP0f
DXGqa6DftGo8ay0h6Izp8iSmY4u4i5GKqzd0/cbeHZi9MRTqwlcyjWxLj3Im
aI333WMcuhP8whjOe1NZwJDYV7V6IL3W3kMGAxBYjV8spXLW9vPtAZ8WRhm+
0yfs7i7wsE3dVlUw1hMmYbUCVI8XxVnQo4f+YqoX/r7HYP1K3PJKv+D+olFa
EtY4uzCRrt+qivGe2qfzghqSpl/byi6FizDn8n+vwz/TmXwmwRUEd7OSwLW5
btU53jp1R2rtpu3r1NAtuD34Kkm1hMoJ1QssgnILalMDU5FH0plx1gzp2XE2
wtTdEW40qb0WI/VsrYX+Eh/wd9umlNL/TfvGAmQ47qEyMnYjfRbeW6WBG3Kh
7xaAZP6nVU5fVWRCcgikLesy/3XZgnBbHDNbxlJQw4aZPecUC5DOm/ZOEPYN
Ph8K6OR+OO+8cWPqJsfl8fXDJI14Njd6Xx7Z15bKPplGFMEzvrbKTylp1oA4
meHkGEW7yG75c0eZlHCsOyuaQhE39JqNr7zbmGAGjWM8JAFui+JonI+FuJ/n
3Ch6qokh0zivdNmEftuQbkOrWKf68dndPs5LH8j8dvIRHZHcVWy5usgmAh7a
V1M8ZmNztmzvb1iWUAbEpVgSiSHR3u++/ku9MVp5QysXYExAMRWWYp5BEU64
ZN0sEOE+ggR0JrwcI6AdaramqzVEk/zFMzFKRCYoi19IGUv91OvslfNpYtVE
fn0/bVc32ZX29r87r/TvTvFdYJJfix8TDrdWbCRjn1I6Zc6o9ycyVnOzC3qU
sxgUa+BcOUnvShwItCwQ/oRU/z9ms/MbsIO1rnjXr0IDgcra2ZgIiXpmPPDC
i66UwnIYJV5eGxT+dDoDqBZK49tT2hgR+LV0QN7wm4AAICaaBNvFbolNE1PO
OUb+hrD9TkfzDDlN2DJlgpsoT2EKMIOiRhQkQ6YTB2iTzfbhJje38jXi4gIm
UbIXx2gghtc2GoGOkjAx5O3Rya1+jb492fbVzWgOBGqQBhbMEoJ3HZiFGK6t
1e6wjx2VEuMqzd8t4wMYvC3RQDaq3AkVQruB7R6Q3XXYr7DzdghgvSLJE5Tg
XLlh8ER6089iGKaWXYqASqCC7PMCY68WiVTNV9qOSix7osOdQvRGSP+F5urY
Dzr/2RQ5C/qCUHJZm4Hu7l6IFuYEWG+WXL0bAgAh/1cfwJcgHGZu/oP/R8sR
MObJhpd87Y8tJ3LHeqHU37BYB/XiXS0xlLmqXKnruflNT0kahR/iYvbOObfD
LAOMfNPqI+YzBcUBtuXFbY2Zxs/pZhRtsxaxO3jVL9s9MZMpYPvIIlyBaNi7
J2af1LDBf2+Gi47qpaiUXnOGrVZgsLW7FE1J6q5N5yXrIqaSQP/ip8xnBChK
jz8tamLhY0SVG6mUZ8HNEapIHB8r8J47FO5QJXcVTpMq+6CUv1jRXZdDa9VQ
2GZNenYsr0oL/Fa5u4K6hqUAyKt3EZRf6mRYGn4NtWn+pm0Gin2TeAFD9EwL
lHdVlO6Lh5NU1an0Qa+IomOnA2Wmmac2DIfa0PGMjElWugsMZNAWZgP0QXeI
eZJ/H0j+knoHNAnbKe18tIxfpBkPnanvnQMGuktAtBiZNrIjDyUuYejYGPzD
MhlqA3+tRXBYi0RYewYE1MnH5bOul7Y49fxhOE17pTAbKsXaAu9MeRugOd9/
NIrCIAAMrHwK/jzNQjGNJtGD98/lQywMfHv05YiWIwWFlNKvW4cFNZjiPlXF
AchHv96BeoHnpjRKKNpokEvH5MUVVTWE+FCdoUBAnAGvi1SLnufqR8twQzLZ
Lxu+jnmYaKIUN6pnfU11lQmG9juvfUHBlDy9gOkYvYtUsdl9+6RCXfZN0q1E
hV8AQxay/TCd4iBmtM1ZtY9IUuhtYdNIbG8xcxkxY+kIqZBdjIMmxHrUiz6l
UOb3uQg+TLaIdmTeM6Jmu2WWa/2Ek102pdZC2rSzLxn/Sc0HDuz4UVWtD+UO
uQ9Ai80nQGJr9ou4b0i4j8Lk6jlUtySgN6NdY0tRRZYiw9YtWMjrU7mVE0IF
n9Qw/4wKGnx8fUCJSIfRQRr6fiTSG0UU1e3QOQNPjM9ohPLPTYA+Z+tZFydT
c0mwvGw6sCYaBVPVsloYxwwbkcWlmGtOhNafEw/v2XFja5gj8KFZOHmktZcF
TwCunuriPUJfi/EE135iaqggvUu2iHuxbTKuPtf6NrDh1Mpd2y7/l0AR6lcu
CoCQzgyCZfuwz0DybywSW0NPXDhMpkg5q4j6l+FTiEfga0jQBL3+JfrOppzM
vRZdKKlZDLkgPtyMVKhWEGXlMDSWaarxYbzB5PWJNhj7IquerZfrVsN3uWfx
YcrDl2stLsxnr7aApaDP4MVkUENjQwXo6hHjQk84rh2H0Np5kh0ASARh7tAE
nDLh7+zg0AWDOcVTC6ThaPH0rjLWnT3GsizOUItulPukLSX8l2nep2/38Awp
x31yQaBmDZBX5Qb47hX++t/RYDr3S/+tBSIciRPTbC42duHFEAFKByyj3tEH
b2J2jgVFA64tpkdVRmVgbWDd2+9AXq54ArnCndaIXnBE8u7fZqh32rff2zWB
YlqqcxIBCe0bGdrJjp4+foDRSHvGeOaaFqmXd19Yf6/6OiiFWKz5I6xUwSHF
QdLe4JYS3mzDwbDe/37W4GD64xJpjRN9WXfNvehQpgVzpYod30WhQHc9rNF/
hm+JYSKV7DwvEyfaBLfpUJ3c7BtXHB5ktr6WaDiBrgnbxrTDXZDPpiP532lb
mVxdBIeosKmGWPuJSxx5pj/Jv+UbzMiN/hjy+xFNuLS0rvqiNRK2Po8e4apr
+uPTcj1EIw61fIsT2EQVJH3U3he4UyZLFoZMtQcItOoxyQ8MXRLQPCeYLb/q
0TJWbwkwpTyO1KTjd5DxT/hkkYYd41U+tMHFeesQhGMvPgChKmYszxoxya20
RoRYTChkRPAoYgoqjmA0KwbUdrweXxE8at7NIZJ8mDfUZSxIrSeF/WBgR7c+
bveYsweNXFV/FZpy+uQ42viQRIhKkenexQrgZGGOdnGwd/+ZA93PxgumAAQ+
lLpFE9UGod3Vj3DU8Ufv2iTcEhP34vq0FPeVu0v+pYm6hL68Ogs2bN9RxRpN
hBpLM4fWB9Figwas+VTgPvmysIacYgSc+1YudT7E1jvidvc+zMjNQOVd6us1
7SrU5H8vdJsLpb0qSMJi1zgnsZhdWEhYEIuWuqS3QRokmWgfm1woylg/KoLD
Zy+ZZ2xDWXQ9R7cwI7hKi3mxkW8puol4ZwPtQ0hMDRDTfHgIebS6ydLUNvF1
sD4j2qtAMB2OFDl6hBU/tMkmT72MFoEz/LE00amGoVLbly2mbWSIis+192Kk
jlt6LmR3JyFi52COo9HOB183OTvGUG1TaIApwy3ysTqSpHtRZjbK47qCxDpC
Ow6wGqGzKl/pDkU8poTliHrtMPDMKDVQn0cuK7xzAOsrZAVM4dB2WSS8DWzk
jqECYgvvgT3gCxus7XYEYKzT5WBfksOR8uHUEzYtYnZSAFVa6ruvUioJ2466
NaNZzTJM54RcTkMiNoWDD1KcDV5Uyf4tXuruJj52XMZibeULE4DxinzPG07l
2PU17FtwfuE8dSELpO8/GNXY4dUrFdxehVLjYu1uxocS5fM9gjZJc6OcmTga
dzH7GpPL08aZmBcvLjEL03VQ5FsLwdXmB9xnzfn1vWGqlBHkgNd+NRGHNoU7
4Gpr46Ssax7v+3DZoANaITx2VtPvB06CnczGVJPxVvsho1hNdyJxzd0xTqVC
p6LX0bPx1u1Db2VSlts8MQ6R9Rdgo5YDxUi1YrMlg/mPVDFYEXnU9FHcGChd
uPayxyGsKSJ0/m2BXrSuVv//Wv+HCflCdy7OZmdUHYWTYOmFblZZzLT99eSM
il7loyAFR7DW8/5/avJgtCCQOVtKBXJV/eD7qGXOwZsZMxyuEzbuAJRwW9u8
O9M7XsC8VJJojXUwnkofloRijc1Gz9NuKQtsZAMzMPp4JWrzIrdSqAraUYCF
zgLX1aUPQP7tdlCQIaIc1OaabMjU7bVx7Brnbxq4rn4NAr7PoO5BwVwHLRuR
82mmRbp/0BAaEAi2+t78f3yIvNOkUZTET/Uhlhi4fsmD0oZEzvBrDBVl42ix
2Gjw9Y9gf1huvCwr2hWr4iFM9rTVACMXd4//XYh8VbvHP+Sfpm7nX7haal2l
t5+c6Zr7/+aftSQnntnHMIojz5W6u1/r6C4/b4EfPL4wdmYa+Uczc0GYmzBD
eYmkcIQDOgIRxJwGy/lBMr4foWkJTLw7OoWiH+qthrPLVhGKsNO+N+SsMhE5
l2nFJH/HLtGrtTUCneWHXJ1BGyeVe2ebToKay+VUSa3qgbWX4huy4SkD9LMU
tW3KdFYT0i/WDoE122vhprZLnrK+SN4q+Ug1Kfo+e6gJeUkE1oRNobzicTlD
/2QKvKihoSzP+swdSPIlOX/iuq/yyOPo2Xtxe/TCemKrvNfEFi56emyS/HSF
eAWm+P1pJOGQH9PZhtlEEQ63UW2paDlZgKRcmBk5OTplLuzYS0Np6J/Cn0O0
+Oe/nmRm4WAoyqMxDJy7I0dm5UCPxZMmL/0X9ZNwJPN25NWbzzWS7zQmtEqf
NCvRLl6L1O7oc09WeiW7Juv3sqrqLzCsmFvuixWBf0OTqoERq5rM6PT3mnix
+mGdeFWJgEoM6tREgxZBs19iIsTErFAveSPX2mM9xIwxLymXuvGj6UASkF6n
rWXbqcnRBQjzymNZl+PW0EE4rpnGO/U33+e/gfIYL7WFoW/b75ICumNU3ory
d7FUhSeeujWsI9iEikxDQVVmbm6g+qmO6v/H5u5N2OsGTpX9zCrW5sM7Uo/6
jheieatJtVy24CLuK2c2eXRHFpBzxLbXcwEzynzivwdTbFrm6302rPpnkGIU
dzbQ4t7if/B8KYKH98uCIRnVcrzpqy1ntW0OgzFz0EIDA4Qo4SkT+OXgrFNV
+yVHX7/4cVHS5xKCzZC5qNe57VYYhzk3k3ohxNA+D4slwNCndN0erOeq3/wA
c1kxwzu5lpSqxvwCx3R5uhQFz/IKgDIrpI0jkRdrkA9PIAclQI+JaMsKjH0W
rln9z/CePUTjawWW1NTGYeDBpj8rmJOBXih1JYXp9SGtggmIGcHI9SiusLK/
W4OWsY6Chuq8J5FL1C1yvpvEp5wuYf5Rlz4tOyqGin9ZzAdquA+GLk5PXJwY
zJiiue7VyI7/YjXfWg2mUbKyhub0JUgfBb+Cj5Sdy8ud0P9E5QZNcaB+yZp+
bDkIZzW/MY1jlOeBO2RX8/1sqz+WRCtSBgFb8+uLFLqKmgZ9hi8TLmYa/Ewe
wKQp0uoSZm6F3H65lo7k6XI82vNg1IRXdZXF7R3KMHL1wBpIKWrPNHpqj6Zt
WkTzBeQcUscZC3zNfBSRYK1q1SiDyXg4dGICPlAxplW+XpIfTX8tqdARd2Zt
a4Eoj2FFakykZsnufswLytO8pNr9mDoRJy8Z5nyGJN38xbphZhc8t3srIHiS
5YLZtOf4Lzjg7yN9WEJaoJ364nc7BHhpfpAoxcMnNluMhCAPzJVBxMn4NGBd
IEda0B4DZYCnLrwoK8CayPk//b/Nx6rfw47jd5iCVqT7xSSmZqyNhSmh1MiK
bW3FCDbi98holUPTYBISlrVFKkDkJxPTmUAliBuWXW4z04BQNVClSsyobhtY
S7GOwc2wbpnhSIEGQh8EbX44gZBJTpPNiZGHkcZUviukTlDmKi6cp4CnaYpG
mOM5wZdoogKmas9hl65OFuB1jaKQOk0e6+pt1uEynhvpXYdo7JekLagMZ0wN
NiertsAXKF9MNDI83nl4VHTUBMZZrV/cAwR8SVv2NB9EK4aHgEC16LOzBmri
wsvJ9nK1NyfqyKGEAfBxAxWzP2P6I9gxOYhnoQOvdGuJCaAK9Yc2ZOVprFeQ
ODz0ro6xRmARMuUjVtnsHOziTgk4+IrykhLUpx7BJ66EKUPi/I9ZVI+JIGEG
svV++flYvkGuE/Ca2A92DiwZ7fFKqc6HDz+HqxOtCz05xCp3uBUMSwbZHwNV
ZBnUnVtmHd7UUMcdm3deZgD/MbYMJV0Os3iF/q/kTWvqc35uzjeF3smJTS38
2kC02a2+oTa85SshSFMPzoaXsfrYAyOleWoyPAo+vAhcFEipYb8S3FrR9xQd
pHCCSAMFuDmKCS734mWKbjKgizftcqj6G+vWqvXnXH8Azf2WbzmKsEiP8OK6
W069KLwMoK9IBDFDSMm1JbgHjrBuB2hYcFay0DEygHylSgvEDgCG0U9mb67G
bL+KRVN2w9P+hUOJiQ3dzhOZP2lWThXmGMSW7ODwcNl1qSnUU4xFmuCHaM0w
jcLLGEeqX8/cp6oYIfNKS8nHTgK0luMUCNbX8y1Ue9SuZBsZODOZuGh6ovR1
jv64FLs9K5wj5NXCgiUWRLFPfyJ+TLEfzlk+gJaPN3V2wP8Esk1ZCXWUccVP
sI5cxs6a4RD0vEisQOE5xobj/eSeMbP/+vyvBXhYvvIM23pr2vRKLstCwb3+
erRL6RNm5SRACQ/vB+BgftnhjgJZlPcJlmTrsMEtKsUtMFAZHKGo57ce0wwq
0VI8jYh7Oc5xmQrVBsChBpmdQqY+9jbRDIeBraOArWDjzQOEoRV4iAa6v8/u
whvGcnpcYH8kH1OiqeDV8g1WBBvFdEpOCRLpfhEwc4I3qiNb7m+B8JUFtPUJ
YmNVH3wr7iHqoPEuGCsKeHQSIhiZmIf64JfdhfVSLQ5HoDBsky4xj12jmp1h
S1noGu0yKDfQkLZLy7bKJTYCdrZMbsSH/nRtGPTdNDcv2HCtJXyTXnzy/RvL
bC3XKRGNowSLsaOB9G53jE2VltQnkisESHIQ6ibio0lLrHqfcNOtoLEXwzpE
TFrloZ545I5b/onosaO6HrtKVdvSjuF5zNQos57RfXwp00M7Oay5xpt7l3Od
loFEu1yaRWYk1EEj7GhTxMtNhIi1O+ZOIz3fyJAn+3yBQr9+mCXT+nC4j09q
SdQzURLvA3niE+cvV0YCt2VOY+grkaWsxEsPdGm3SmnePrb4WpxczfxSVGAh
qjoTzCxsXg48e1fo3p0nKscM5bmRdC+qvYmlM7SeeQHU+2qARjQVyMEeVLtK
kmm3yS6pYGMkBX6WH5sBLj37vXDV2uhVr8Z0aJx3Wv368rA4Q92qnUu9UeX9
QJLAizDio/iFFWeCJPCHqN6LBfqqeP4Qx3lUQszUnF7CU7V/SsIJ1446lwbR
Qo8vWUFp8PP/Mgceid7w0Bl6blHhWmRIY8TI1fy5IkQ0W0iqRgc64vxMAIQD
kX9XVlqXvCh0o/kIVklXbCcegcjPY2vJRFAVN8f2Xw68T/p8vDwUGBrL6Sra
taVsijd98EP5E8RfDFTW9J/qkLWMQfZeqF+4wLcJJVLno6gT5t2rIH5xsDH4
bawOS12+TLjijekoyYxddASzj8NMTYXG4Dp7fQgAl+2P2+xSSFfqKjCxbcfg
ceDZpxVPhxvx7P4HGXmTMSBwFFyeSkoit2/LhfGYFzYcDuRQ79dK+M7CGMdC
04mAT1E3wm/QCN7Szjll5zcCwMafhHMddBcsOU+Q4lcKALlEb3M6g4cVMGuX
X/Lok8yVfPTRMXoHXJQwS/lxgJl3nPz/eRFpax0Ala/3V4E14W9ZHhtEyrFa
yEeJruUgIex05X6Eofk6yXBw28vp/tRnpNabv4JX7sbhfr2DUJVpqFlHN9Po
6Bfl7Zn4FfYinEIcbcJL6nKcsdygWCta3AvbAco0UECGhXBBdnEkA97S2e1+
ZHETEtqRC2dDE+TjpxE4SSsfeEEicSMpNmbwCNTI3RPnNgd1H0y266/c72iA
VRq1EcvHVu2SQVlgFAkttq2oZlSW4MTSEBUFhuMMCppWWNmwlGwicUplv36I
as8fJ7FWXPrSUOyd50pUlX+ppGHfnRId6EZWnaYQwz8XE02W4OHesYlb9oaL
evHPpmYd13kFPnEOW9XjowytEvkCeo5W0xEM8mSexJM397zFSK5xAyqFUh7S
EG7wUrFBHjyam/65tgMmHWRXlVKi23BXN3br5/lx7thJsjcP1TwNX2sTXFxn
FwIKahj+XQR+hBH+UexG9VyS5gEQ+yScl/N22mh4+34SUylFRf2xl9xRk7j+
28742eA4uf76Q6ZRDltcF+dMholha5ou9V16JXfClZ3f/8R+7PabA6H+9ya0
+8VncFVF9pFsuD8YirC+oV5zjiojrJA4JDo/T/kXVXX9ogPg/txaueCVbfYT
O9NTbvJfucK7GnnzBNvjgZY7W3LLtMkQ4DaUdQyb/3HAFPWHtwdGVg9USHzG
1rkkEQ2NNCt1N8OM7vMDZa8grbSJzrSPZu3eh9SIciuzVLhW32P7GotobHT4
bNVhjyp9Mx7/91HlRl+Qk0LqtBBHaNMR1jvKCDffVK4q/eQK0gm21/afhbcB
3MxmZRmqGtOhhK6uJTtGJZ7zsL5X8P2KZ4eR3hc/foxEjrNCpUfsByRIzc2r
zNYXudVRT9YH1JjUc8ccm47I5kF/x5rJYI/nm++BrKXZ4iGIJPVKr3Dh4wkN
TkbG1kS+1tHW3bpWnT3dG4Acqut776sz5fDMZ3Cg6yROTnVatwObAeH4niXe
jtHyh9590fA+2KTOcaxg8msxqjPciJK2FquFFB1dwOAZAD7KEs+keN+5TUIj
EeQbu4VE3LHzWdZ5t8IeoDs9HdXn1jd9edl/pshNURiKgfIBGCByOxIOe8db
PXHhyQh3yBGela8qRk5it42XDQH30y4Mfg+FzDXHorC36QkAxA8SgoLocokv
C/dVHlHi7pooZc6+UrzmOdTfkOYUd7bY1In9E0zGqUuGoV+LufdJhFmtYDOC
UDgYgPHlkoIDgbZxEGfogTeP52fV2SvfpkDnLPORkgs6kygMaGSl2vZsgvwf
m+YkBpFpklEPCJgseSGtRXYpCurZICdHaescQrwy8wlZ1TL+X4bQdKSDQ9p/
yR3VHAVXgmJmt02aIIYpDn3+o27cUg191RT+xnRqTuWeRxLOY1tLuBN0R9iq
tW2hbZtvYjew9AKFZPT1LDkjKXCFqW4XlDRNCbAC7XvBo5RCiyjtEi7Dhw3U
xRDlfRJMBwEcuBjtHdgzzx4cHaKdsWbHHxEFrfP9YOHQ/Ts1KU1WcjMGQLLg
HFdmhxWsu06ZHvCv78U2R4dJMTLCWMWxvXs9tAgMbUha67pqjsUNRdSsfiJc
jdX1AkHLYf0V5CMDKkk8E7JcLlFS8XNIlGd/8PXfU54SWWZX7dErGH4GjO5d
tp9m+JJpWxmNDe9adyK4VoTbvK58tsqTLT6lOQ4xp1Ve8hnaYZ+fyHXsBiyc
auV12r6xGpL2cGrev+bEv/Tulbgck0qv4R0hir9VJrifyP0UwBNzltW/A8WF
REkkVURsG+pbrRc4EeDaiDzbTT3mJLRlKebMwhfbUkFZQGLCTuwYpdaF67hB
+Nv8VrLnkWgYvowrOcXiGdhKDZD1bpyU+Lp1Q5jMJ/8vp44NkRKNdQS1IbJM
fb9xb8vB7PUKB50jZmoQgM4iuWK/Y72Xpzrbenv1QpcZCXnG+mz60LVZW0Uw
dbIEED1yA99rPwrT/vr8UBZZlyOA05xZ2DI1SHiPnEkgPb+See0LSEQDC9SB
MLRHKJASmi1u0HGqrDyt7uyCua1DNnr2zygrx0nPf2o2OR+svGwBr/xGEhDi
yJ2UXneu8xFS7hG59UUErMA0LpxlQmZO5JN580QW6LpLvumwCRlH3adwYGZ1
8AGIUVXrsOHwgu5ZXmfzE5E9d127vDGeyEKUU+y5hIT3rNOsHB0U6fS5CbbM
FCqQGaFvNgXyvZQvfKiDnkZN2V88OtldMjWggFr+vmLsz/iivf59Pn0JdoB8
B6mXjYUxpv9EZWbjT6lELDrDpAN3HVtskyR4SXCyB75poT7ghY6JkT2ny+2O
IkdXtKsBSER1gJs5pFnFbRvWjfVc64v8I7E4zIoi8LUW0VZluyKV9AkyZTca
eY5DIwwAjuBdZYCsWraZcqVz2UrW84tI4k+mXMSZKTq57p+s9lbbbQAXGOtw
iNhC+0f9ZyC6Y7r3KaaGnudm+wMFObpryKoRaUYCnVVFa55f9rLUCG0jC1xB
uxZpbbnslohYt20+05mxv9jHGZNZUa2f2VBjZzKVkFlwW7dR9MdDLGvfA4fP
hvHuoAxD2tyBpu7h6PvWsvMGPkeMV4xTxhOFhNKBP1X6mmofUw834wHacMVH
93dpQd6olUFqDgxtaCKwMq+oIHxtGit7sOjUXZrwMCTK/294Vych3le62cAZ
X7x6d0Snh+XIghNsMevdmsS9JhY8IF77cptbVR9JjuqQo0riY6YReof0I5Wj
WGbuknd8Ycr8SYukV4W1dG43gSKPjRxX7T7hFZ2Szhf3n8bagly31eGdWmuQ
2DuN9nIcD7KZUinEmV6eMJDW1fZqVD/ISyRl1QOs28aOCisxi9PFkj6Jsh2A
pxFlwQDO1KoHknjPfVNCZr5oM2N6OtwKZC5aueqw7U1Cotk/W2oAk155skTc
cPoPck25LqQJUCWw5b1r9xZFCXovdIfbgGXN2aylF70+QVLPjcUkXOe6hZ2+
5A69CDrBDzpNNRASXoB1J8KJl57brxaDIo3IBo6/Q5RXromb/WCSgnmFWvhf
zktvt0pyGNPUaFK0HAxjRqUAv+YiX7UvKfRxgrqAvinlvAD6B4rSK6wGiSD3
Bqo/6ECP/A/4LGDYdCY93z0A68ccCKr9uMM/U6lLHYCZP1CESaxw5WHQ/IhN
vBaLFAGmpPPQG5GXcQBfcOxwVT6sl5iZ7jQrznmKHbFO1RjHusY49HWD/2fo
PgYxcR1M8uEiVVv3r5hWPV5YgCGGV+RxsTFuClolfGQZD0nRggiP3rgWiy4c
YY7H09mY04FVVwMAo40oan0D6sAuKVu4KCohDlnfnKgP6XPhveBSNnUYY8jN
5KiSt8jWjkGLIkfS4ob18XskhTMajcRT00VfJANPO6UTN/rzlIvYu+WMWUmO
pOiAQygXurOz4Sec+7UKgq1CHCGYgDU7FP0wPmOPAUM8GS8dRiOPIhA2YDxn
t84W2XEKf+VTIbWFWujzT+QMwSspzd4JbKNALIrxt+J80mOX75yW6+u4fAGx
Xmq35HPdR6mmrl9wv/HWWESoWu+XFq/wXE1NDu6HndfJ+NEyMGj2Tek+zjqr
nb61UApOi7udNEvDS0Vm2oYC790Pjo8q8QqHa9LT6gAZpG4M5Rxb8gAU5xd2
S4RbMNM4+7Al7b7wZEpbMn0Av794VV1lJ4hqAadpu8GlvWETsuUJpMRpYHSi
zdPEt88Gp6NwdZ8QOcXlZMJ3VNS4QM9njLozisHBevkhJud79OfO9BB2bzzg
IZRWkiKnAkW/a6xI8s9jf9WeK+xgQ7aw9Tl9Ppnh2yzplOlJXAvqRjsvg4XN
L1g4LGU5Bc9cd8+Tlay4XjVlW+XRXZ9gu5goTEW6hb/87gGwdy3DKv2eT7Q+
yrOpY4a8t8PBSFUc+nsvxqLynjti+oo8PhU/U+++DYfb1g6cgg83Wu8+XIgD
6BlToJtTKBVBgNJqC1JFS25P3nPfJo8WCCHPYJehcGMAEDQI8Shsc6KflxBl
uE2YLOWI9G4MBx0ogQQfM3ttj3c/c1Us2pzy0BYEMikAfEhG7IG6bWfu7vca
L2tgcOQW2O8BRjPPPmwtToJYcbR4H2OcM8lEZkHaKQtfXim4rHdzmmecE0Wk
N6NBJzUqAbkWkZwX8FPpnbK6zivlwgTdd1bna0wsu49Wm4bPYgN5IeTo5z0d
Ecu9OEC+ewmCqjoUJbPBCn6T3l900AY0i2hGWahTFfMlb7AnsoiwInFXxhTr
1nv+dROfLMZHMQmfR9LKurAUwk3tcFJilTA0GiwzTYBfy47WcBCBhuYvHz9/
jiatnrTG4fHEmbyLbvyNcJ6DwQjFV7YQRBM46bvBujnZKFzJglPhq8naViGZ
nLo/OpmVaYtq0zoOIbA5bZPLXT7cb4wiUizwV14Zg7aCCRwnavoiZaAcVA+D
Krsq+SRGtR9N4d6+1Js0lrtfpzZwfLmJrhSv4zwwLbRAS6DlibEGVQLWlG/Z
KVYaWw9U2M7Iac5qAz/gK1txR5AKnhWXdI5K0iPlKUvePtpQGPaQ67bisoDH
a+2tjjyanEOC9GdZkl21UdRsOGepEx0VM88A6MdkxeAP6rxXauv8rq+fjujW
kGdKlPM3dCbGpVHeKuTTMR4KMhbSty+JPyYZzakzH7xvVfM38M7cjrmV2VO0
lonxICaidVWDjzTx5YyvlugapzNxNDzgLaE6LaYNo80hEg5hNLyp+ykRphOc
iJcAYxRNj885QdwJs//b+SILkcHTuwbKAORxGd0zATGCawKwDw6ojpVjUToC
GnILogekUbv1Y0FFgE2b5ccm1iGyi0LDVhg/qM3MZE24TR3x9lj+7cq/1TxY
JK8GTXEkHVA3qYa2A3k0pNJ4keKenkjFmMJexuSyGVENOSLkbC9QgOdpeFiK
P1nRhP99fx+3wFjFFyz7B/K8bomiL6xBq1VQMuzAwq9aK7wOnccCOYAi3hE6
sW3Q8pyf10jauKXtyYPgPlTIZQ70cduzq8UwvIQfFODAnKuMRnmzyzTKm9fB
7qu11bP6kfmi8AGXcxfXehAtxem6gMT43E/HE1g61UI4A/ceGklectRGnRw4
90SCqsar2m7icf57CwZFqi0sjxIM/X+tznAuh0DmqGtKkIUEZqPN16i2uehw
W5vLklspzKVy7PNvx99v9rLpiitC/bhY6PZmn4mnFFFRVby1wNqD6kh2KL3j
GSZkSXrsM0vIrFVw7LxS46OyBAQkWxP8bJ1rNm6nTqFQnejsD2GlXfJnTrsM
O7OuQoZgxg8YPbC6GTRrmjFDCS2Q0du2P3aCyCG9bgkFFRvy++dSs37F7wsr
Zu/ydv0s/l/z/alwiFyf++878eKq16f/br7YYS41ZG6wXStSza9NLVXzELRR
uOOOhbolIbnHWKmpNlNYzr5zQk4Tlj+uk0LYkUs3R6+WBDglEpmkHoCDZTNR
qAyDOujlUWItcTawohgORbrsK2kl1WtSPJGwr/co0wsCBh6MKP6W+nBNFtTw
a3AUR0qSQplR/bqSZzkKW/4g+bzSG/GvQVSyMFc7hngCKsHBkLn5aVdYzP9F
DHJcFP0GtfY2eJ2BUaeNeW+3V0PYbAP2B2Z7pN+nN+lEiGBQmVAT5ALJj58/
GouD2qvqm4etLEytcDl8SnZOi1HVe4zFuaRPMGsYCOWd5LelMStZ9GMetWFB
boXzEVqEO6FciHpLR73zJj6Xi6+AD2kseTkuhM6ZfbjjVwnvH6G0KB4ihak4
mMYPSqOwRA9mi+fRG2FFCja1onUIyMOgb4kXACbfLg2n0yr8Hv7fjEHowV4S
khf7NpEogrpVQc59FjkpYL4q5naP3wwQ36EvgBxjJHg4nIpmCBXAzjNfefID
c8iM65Nd29MYDabHedYqlXdKIzaov8ljQo3Oa55t3MrW+osC9Y/ZnRo1ucwf
zP1ygvBEAffLM0QjAg9pBCjH1qEwOFg3CJ9kQhYkEZruYGMCud2859EU+JHP
BoRq5gd5XZHSFV1YIL0Sz363epYFVHA68ijPEly0CDZ4LwKzJFaH2tn2UI8A
dbqP1Sgyz8FbBQB5BZpzq6Fi++0yMq8Y6j27vTMDWRN2xAaBHwQGX3QoMbaR
GrG+i4UzMNhZPo4TukXti2wV4xJYqgd10FLeKeR5rOqaE8Y8t6cF+XJmejw0
p2WszIGyz67enq5e3AUpQ2pb5P9bMMwaTmWdvWD8gMMMjd1X6fOf09kVDP0a
3QHOq+CW4ZafwbygBXhJOUhxKDvNgYhNgzUVCXZl6rmI8QADfBQa5tncBXPa
ldIN/4uXp0z9FwTEUIaO2AEFH1ijjazDEDmzfac+4/8sJLIkzS4gIgn5j9Ld
sFvVqM0R9KRcwBBZwwhNcYgoRhszjWqt7HILWdxMnidmo34D5TB7GfH4TWhF
fGX2VxqeyfVQGmv6yTdf2IVbJqwjv+ht9HdrNbnnYn8kcid7VetT4bWJbbrm
iQXDjrcUrVJCBDmaQdRmUVpbXE+siYctnfFDo1/njgnwk2kpTSHx0q/YoZBX
OGc4zm5RbUM4a4fig5OSRmbBpOd9JxaVWx+FQmDfaV38SElYU8806vWhZUi3
fH0cx27AWY4A7N8YMbDJgkyzKer6EQHiuax5kMQiTY6Mn9iTUcVxG0VW2IWa
FvZ0YFnfVfn6p4Cf7GUKW4qV90xDbAkjLVj9QIfD2VJkxQng2aeX9ghFNOmp
QQquFNckiLN4Zvxj67nZZPKM/yelzdoDGCovRSw/R8/NxSAcygkwVzsV/g6X
wvumhybpESFFC9mCICo49+J0LFnuPVSrYyvjJUBoSH1tmEuXf2stYPjlthZK
xY0get6mWJ3d1gnz0MUKJwGrrEMrKPpQw+kJ59OUZEVMkKVtMcok1cQjBrFj
Rwaab8CtydZqDgLdh9928ksXpL/3pqhrGfFUXpI2IJfhA1LnReAQOImaw/Wt
6dZ5z8/inccOqNzPe9lV4Hcsbb2IbsGHCyy0NqnxMJ/mDGaOb280Iq59wAfH
TtFry1wgL85ZnnxzCgocEd/3jTvEqGAk37D3tBBuV+mGaJvipm1gG6yZFwCm
tKre85NsvmSbRgMxj14obbHXVV9gEz+Sc9g/qexzhHSgtoiGTYu5o38WyDLy
i9YUTk6vfQVBXK3Erz1x1wvoLl2Fo74EjFNPMcAdLbdrsFKB0sAk49J7B8sO
Wt9WcK+eMaxsvmFurokRFRmy420+2wq6fw3O0vWo+bIlVx3ZX5wj0FV0ITnx
yAWZpF8L65uczsyPNc+NvSaO4fYRkR4e0sl3N3gMm5X1N42XlxD+kUQVqFHA
QVI2EGpowkhm4lZAK6CxM0vO9EsLa5dv29mZzwHpCl4TLeT4DNIS8R2Bp+P0
CLIn5i1674jT/EWVS9Yo1ScbcZj84VU1xte2aQ9Pb5YcYJ84fRBaZa7XtWIy
fvSKRJj8DuPYXGlAlrvrZXMBQfjoBHh2Wk8HRLflX8bBwtKHRtQ+a9tMQ8Nz
jJ8NxofB8C44u/k+S7GP5Sc26wZ+XCUM1gVBNnxqhUV0u6TuQtLZPDe6sMK0
PU8dyhIezuA35zUBfVHjlh5K/LjYp9f2pYl3hnvlR6SHL1VxYEfpwEPS/G/3
75FMQh4jdEPU5CY6W5ynUWtiPfXoW17XtCXwIRly2ZHvGNJ1gnNDzWsdbh6z
+fdh+XX2wtsz7iXNSteHOBYSrvZEpLpWbeZh8zwE4lftpTI4whrBV5eu1ths
H0KNhmquf7VKVMTL+1O6xtT8vqVOOEtpUBb/3Iocc5TenrcvzHjUgu3oyD2Q
v3TEU/gZILlUIu5rPXosIL9qiNr3NNJ4RgKOflfFtUuvGfhiEIwfOKPY31Dt
aPwVi+Gr+NEgCgvjtOoYoa5/WWa6RHh599QFXx/kaBW2FRXAD7ln0OZbJcpD
kBC9f5Yg7lSLBfmUz/w/3qo51QdLDHt4sQFJ+JBsvFPDoBPwrXKl4vSOCl3v
A56gREMR6H0ssIDWccXZdcwDQLRHAlkYmuTAkTP5TEPEOp04iiGMFmryUbEK
9mZ8B4UdZduAKQhtchEekHI4lnemkxjZYK8dXz/J+EVYXV1cvB8Bf5WZCVBB
QXXS7hdV9ksjvi7YHFDLEDeepyECCExCIOebHFpILsJEsxsfGM9CC+VTV6Qd
3XdNXXxdSaEUvwhaA2yGLJJD5MnpG5jszGXtBZulsw9l0eR87VxhQ8/ILKEj
qlEOzbbNz5ltUWHYS9YkzbIovzyeIACw1BIXe3P/ifovfI+ZRv0Ov0e/co57
NoOnnH3sy57BYcLTJaB0K1OsBjFfjnmBWrzhiVfTvWor+xJmivg3i5oDXnhF
NVaq5wIUMJRbe2wrl5eQ9d9Lvr+uSgaV91oZo9bcqPPFYBlFjpgiQxBPHc3U
N975vFal3iHEiesWJdtoBYc2TwTg2oEzz9zqGcE8usoi9qCsXW8ZeQbsMxl7
DpG97wv0vzMclIUUJO2r2EblQk+6+82TOQUEnqbP0rKYJ7QWBasAB0lBf5d7
mEyFvtEhmlcRZBCbD19LpSIONhwNpalL54JCVvwsL9HZDi0b3tA4YeeYCEwx
jpU14zeZ7zGffLsfm76pYgRA9ltIpt3ssygZbByDUjliNhf07OEsOMbVaI98
5ZAcpCLY8U0OL0MBjEJ+E93CSNFm/SoZVQIdGKaAz/RCRko8lcMZ07s2+bLW
Il7OghRkRHiUvxw9pueg8i7BKwwTnbOaputKrZh3VYd6zSPFJQlQGfNPKGQ1
rHYM+TrB2vZoJPx/rrz7pQhUz9Bxfg4UlJf3oH5JYnEY94J6Y83vinKIbGud
d0k+yod0SYU2jdDr05uPrryA90uNwpZdmCsdl7MBL7/jSpCUsX7trU2sDQGi
0IUNvl+KgUEz79kIsmwr2nRe7WDiaWGtpAuVz6567ujhlef8Zj5+yRqBWM6L
eZLMCmEDGCZvf7Ezk6f4VlQVcLhbwuDTUSjMrH+hROp3ELvIngE2fZtDHJ0+
Bp+2eTUgITWY/Kq/wx232VLl6uqzmb4AVBpdTZ8oDfv8kcaMlraAJehMyg/y
EMSZJBFJAmq2etXsBm9xofNvg6n9+IvO7GM7Jv7JxPyzxVSMBV15cUIRApGi
KYwuyCijIGcJDebkqbVsBl8JhavTKEcsRLx2NgBbEAflM45fl0i27nAuZs60
iPfWe4pdsfSoGova5vSvS1FdLuXRI31OMTMIM4mbBwLZhd+sqy4fM+BZRK9L
bh6rhWm5+02d7e7OV+CF3DqZXvczWpZYUzabMV8PblwGd64RJmROuscm/a+J
8Qge5wVkBSyEvft7kt6MuKmV6vHz3o0FHPrqrV5boV7ESXmAWDtuiq0c2W64
lrl6EZn5eXSA85LIYarV5qgV7HAiowrO2amuaQ+bYjqRpLD0A+WCSumSP19Y
ma2x6S5m2WWac1OMVlIwo/wKoHz+RSsFCW0YzJ/BrjvDhBJ5csQRfEElbkKy
T59D8wPAnuJv5Jz355gJQgfQs0UvNBtsynnzP7/fmFR3M/hV9dPS51a9vtDN
n/rTMmVHRJkgM2dJXpYwBAuVTKoNzfvTE5f3XwWDMOg+vKV6zIMBu2YWA0Mu
CDQhmXhruVgS3cMjL2wriZMy4VLeXWTyzEE4z5zSY/qjzkG239HiaAwme6sW
8F3Tr0pOfuucpq4IC6/UsP3eg0qB2YkNiVwy/4cDt8EuhUro/t1icIsGy5aY
SaQow+ViJpOjopJThzHgNmT3wc+1FIQGWdHtDB+2ik+Umjy7OD56Y4DKuW0a
4AmYCMawtNUjvMo8AHPzNbEVsv6BX5ZOMWXynFO9FhVyy8NyZl2Vw/quV1V/
6KB6ZdXMkUARZTQgoDgpugHInMfsYChgEgH1rTTaUuYkMnGI6qgO3Jfubm8i
/NpYVfCK6xMSbKZfbRC6Id2rg1arizac2p79EH3ok3/qwQRImP4ywAsviveF
ovqWGVQmvNaVi7mP8vd5O7djgp7I2DX1QHdWsupYJuGvABJZSKZl5eFsyr8y
Ds/NlzH7akTTLMDqqMYbWoiZxBPS/jHV8h2+kIC/LUe64iTZMdhxUMk46wOM
fKha7ve252UElCKJEptFq0/HLU1FQ8MHo3Eaq+8W609UHZWZaavmHTSFl5F2
1wK7hpAHthb5YdyFv2KZzjZZK8v19R4RCDZ8XLeWhsb0ocRaX0EkOXXRsn5z
1f2Yod95mNm7BTeYTNonnXVklCL+uOs6jWrAEftI3NEk1dM6LOiBgAHUdxBy
LBpL0DmKdbrqe83ovkqyVQoW8SHlcXCm6jF2puNuKyS/yoKEYxe5PXvF738X
oOK1PcY3GuHCg371y5HxJ5s66ah3Dv6cCDogyjwlSh07sBoyJyIS+U9Gfc3x
9oYzxbcs5Rgln2bPQB3m+oTCJkNvOtzIapUP8lAJa95zIR+EMEbP1C/zbRfi
XVG3jR+yK2Bxlqs4FAHfZCZ5cPxUJrZ6Nfle2PDHuQSnVVfEh6F89yaUaezD
pM3ABSSnn9cR32N19IRlvU22nO3b1qPf2Ohe+NqIAd0NXh1was+KyRcI87+J
qDsv3LkfwCoT/uODKduI0iBc1hAXA3pTF2OL9sasstn/qw0Wg7L0Q/kCm9JH
T6ruZ1dF8AIh8KiFFDvOY0/S3R3W2jaaYktkh2z3Z7OnFdY3h9gXfRQ0Xw/d
3WCMj43Hz421JbU7nohUvA6exQQn9qTRO+NCRBkZl4vAaF7zEg/grSvgo8jl
a6XIhSNNMhzrulF3xfsfA/WhCIgZWqxjf1U51evFZ46X+63EElLR5fGgwVXd
Ld6dyqZkEQnJb6cbrrEJNaDppBuD9z1mNfVMvz90eiUh4U7NvBcuPil7xF1q
mAdXU30HSzMyUQjP6xUzlvN4xUWyipqF6mnKdvTBY9+yKVIUHwExyNlRKGcc
7Jim5URoQT5z2JBzljHpzA4kwjiDzRSHgR8v8zE0ZdOdryg06Ugvmuw2DEwK
XyaQi1/O/9mhU7nVRsVPUUJvZHNQsfPvnA2jSHaC5GAZKkwE1VvCdoYeFI89
rpLglyP+4gPvrpXJXgehf+rPJk9W4N49ldR0+KT1CUvxncbYVpNHf0V6Xtsk
jrjU3HSxd1yUsnQDgVC040UL9CBfNR/SsgR55VaD0drsZTeAgHjjzwfGI3uM
/5Ht1sZEwX5uWdhwZ3iIXCjgyvir7OuZfjLywBRbRxh2v39ztTQlHB1kW2IA
7rnvvoWUMIHBJqlXPJLxA8tua0OO00cS8asue3VbG34278sVpBW2Z9NmUdSl
2wJm6ZxzA1qxDjNpUI3/68ZlX3oxYeb2Qcycx/vyvKXvOX3OStQdPi7p+ZSh
b7fi4d0yXFOfENjdF9pm2chCBpgRNwkaJgKB81trPL+86AeQSBP57PsaY80Z
UeY9qdOS7yrk9byv32mvBDRSRxKajNlEDvkjnqBcMRRfh3PvXKzsh3zEVNW7
JtJrLaed8HTu8jMTxJRBVB8xII07ZklBDOnEMcrBMCUXEg+6cUpW4C1VwMdI
gvuLq87Df6qiVVOZO9Dm0wH38Xq+VvMcowKtXrUzwzdqVe/Nf5eNtItGuYFU
p39n/Cpjtsni1omyzovKG19dDgRD4WzoFrovBrffDjWrBv6peVpG9iPQ9kkj
t9AzkVFwnFWvVpqNxBImLbDKeqc+p7MHZGYjU1jkO3hWR2BEQZ9WQkjQwF9Q
/PhY/h7g+Zeq0DTv72Xisda+znxj0a8r3ot2Fn5qIBs1yiBQvL4MOrrLMZ0z
LkNruwcySm3PTLF8QsssAGDJv5dUxgd7k/7nJPurbRvkHZAyG1NZf6BPkKMp
awhgv5kY5OtLyl0EP4m7Jm3SASlz7P+61TkrAcVjfry3iJavrJ4qinvLWWuy
Rm36/rYPhFZ8601xUEKszyvXh5mQN7NvLoq0TMqeJGoetDcDZoNNTzJKjatL
fDdRv0pB8/BLYcMLplRPxnqAKmOzSSh8F7d+4d8ZIkp8PTeL6hb++5+miX9J
XfjNA3fK+hf3NOWlvI3ek9WK9LQOhVcn+dt7XRGbSfkyxNmijik7tdhwEQJW
6nmpQT34zz8sHDNSdQgVBwaX5ew7cD5Ee8k+lsETk1IjcS8VpeDfBofPKgLc
bWU8kH2gYWDSdovHjdtSv5DEMyPXHA9boK3zDHwcR+t4XZqwbEEM/IPNwRG1
hHCeQwG1nri+X477fNiVVLaSu7GUELs0ikZ4kFEjrU1zdi/FvuhD14bVUwdV
BDG7sUiqhhhXAXLGnmwclhai6hLz0heqXRg1vslWRvcDHjXLg1pQEPeILfbh
2SGCKdO/eb+o5hrvFacJLiJHmTPAiy9puLwqY4LVpNq6ZVMGvUQIOka8650I
cT6WeJBr2eC9t2LpSDK9stRgRqAagburlc2kV+3Lgjfwi9CSXKcI/4kFLuAA
gbszojhoE817CnxLajyiYklBZl8OcnuB5RNmVRLcBJHsluPwETfKfmSz/XNq
k/12VreMJqnwMDdflTGw8XbnGuDvTWzS4ktcJQK8wr3SY85M0A7IJVD017tl
5R7YIS8A6AOR9EJtol5bung2FjOCCYI2K1VXJlEBAzwsuQTgivpSfCKrqRlR
uO8qjhCtjNxJlsqwQylg1SNBS3NPp4484Zx5ICW1UuC3TcvNd9RyvZBScAZB
7tZ6ad7KDKw5rynhZPlGLwb1AbhbrcoGtMsRsADoD2q2rcewo/ZgMun7tFvU
wNgA7YZy+HHexo4yGadFB06hiPrf+ctuCy8Bv/AGWbA+rbEWB0mfvMcM0WZp
qcP0pzgiMFyfY80Q15QEa3A6k6wFJ60vKOk7NwZSAWftkWwUe/pzeZrWfcvX
yRw3xxfs8mTZHcRInqwt47uhGfW4T5JGbDt3kWtlCxljuK4pvv2Pj8XixUIN
qjF1viuFKS7igJSVhLy/SsxcgMSCfB6KLOi5Bq0ZTI3cE9C0H6rRVxfSlguo
sumXUYjwswgLY+BYcOyfxoInFm/kYkejDdf+D5yUJfrKbOL0ehUo0fzV86mC
JOOn0/8e0Sfu708Cmv1N2gpx8PU3AsinjPh7PDu6MLEpA0prfaZemDu/UXRe
o+bD0qafxqteQWpupRhanDARCxGLlc5Pu8vaeYSVPPbhTyVD8NI5UjyeKIXe
fjS08juHw+OwRXpF6mcRdp799fGctR4QVJ+ZlbdOXxqMPk5swVy0DGLUOwGX
F3zptJO28QESHHFr60oAEwGyQrLp8EeRjf+1WDvSb78ad2Kucc2VHx3bRLdz
0BmyfWnedRf3YwS6zcODJ0FZEN1o9ciuqVyNv1GUXvJcntrFfKRmBIv+6AiY
X32EPsSr9yRdNyI/eC09G/0pYqkA3KsHxGqmJVwE5S13Ei1+j897Ent7Qg1+
Te3nOpPAcB439S73gHr8jBgMaRvsiDWJvsakiQOYfssPIQK+3VhAGy7RD9Zu
kZcZpVzCl9mphLoQ2mdyiMutQ4LNoPnMcV9pLFVH9uVujYbyaewOKJq2xJB3
pb85AeYtSiy07ssCpVrVTCSd/Q3qzDtJNnjCIYeCx1QCHO1mei/3sFMuEV2e
5UkbcVp+3qae2bPdBwEav7iZwz/rmwJ8ybM7I18hg1Vz6DoaipBPkdYe6eUX
t0+ma2FRqlqSOAYFmreuD72oPsI3KIslHZMI6SQ+65M9qfAQID1VeBh3SI6J
Rhk9L2i7XHc5jNxoDVZ8JMbTgNq0zkjlrKo5jUGXX7RPkaOabhH0mxcuAauo
9Fddbfd5LU1vulYPbDcLj7kSE6YhLr+reAj865b0ir3/3KIs1msiGcNaNu5c
YLLWzZeVWb7HLdgL7wwNyFSLnbxuPlNBwkZadFt8be8WMXntM1V3Gm1Y3Iav
8YpTg3h++zPaRmUkoCs1iDyYfwZpY28WerzJupRJPaPdFRS1OwqbDoFntBSC
PoCY6TK2/YbRU5zObCgYfa0QTnb54xa6Aotn9I/oUPCkDNPpaNjDDe6QmtJw
zJWhtA4n9GIHNnZkYUQ/0fbjEqeL8htFYX7yu84jcxO5HOmUVvsXYx33/7i7
bPpvlpml+sAy3yLa8e285nTNBnyXdnzEURiv7Sz6L9fRef1e44zsxWbLfWCO
wVrgDcc5m0yXKS3JL7O4ozBibdQQ9DrPqTkpuCkxw+Nxm8EO+UjYheKqFtjR
2ugHm0vOo1zWI+GjfkMACcjNoIobmoQVCK7AlSmgbWgIoPop1nyt/3FnjYd6
jcmsF47IBdb1LbasoQbwtzfarSzRUG+KNPgg7TBOvwu4lScSHkgVDJykFIbf
Cw7y+9UjlW2Bx9RjwaQtzPUQiqanPxBWe0PIRdLjTMjh7IZz4lT2A9QGJXea
a10TWjAhp/3ttALyPEI7bBUTr7HP4kZ/f0rj9PyJL/orOrX92gGb6nYrz123
/xNEtW5jGzb2TDiQEZytRKAW8dioSLX7vqvdKBEMso1edw9QENGgiIiF2+FZ
IJWU+oJGIH2kuFrqNfG9147sE1GPfYGHim94UAOyBkRWr5sItaHVbbS9yEoe
o9Sr3FUWMcDBQ7NXe39ZgUUHTd0Np2aRHUraTKXY++9cTeBw3woIRjLiXLef
LeJI4RZOdezCE7B9ifm1mD70C/HAjLInpEp8uEFIQg2ZypxrHJrw3gRqkjbL
Z87ImfZHk3dkjKryaP2ltGMAVHaqkORIrNfUF7ExYqKYfHKL9Qh92Dhe7LhY
NDVSaX3MLDzhXdZ5X2l+eWjY8GICQnLqV2JWSyzZXEXKB15FlzLyon6vXCp3
moCBgCLf3i4HydzaHwkCSkHmv0U5i44skYghzAXrruF0CLqYTAdXXYCqd9xP
3jfNo0fZ19l7nHD76+NyQwZ0A2O71KxpzCyyq8yplf/lCiQITV9Fc85mlZJa
Am1XEoc1SqADm++SnRirOUgkmsrqlGgVHEPcuWUjkE+V/mZRjitxo/YBJzb9
I3Icp3boyJT86buS1GkJLb1iFEj2y/MmkP0u6bv66eoH5jCmdo7eZSeZ83bk
6sPbZcNdv+/nNsOs2tySa3d9Dn0stMkc6+IF7o5w/a+y205k8lh5oKjLFKa9
OA77e4W9EiDn0EzgyQRjAPmdEg6K52vha9X8k47vK1WCRbgtCYjv3LEE8P0J
fTUvDbAY0F1O0gbi4L7Ly74UHL7Kuw7gsOfD8d1MyIXl59WMEj0UtG0cql5g
P/BWaDk6Iu8myirJUybZm4gA0Qcu77RbP2+ciNfGgT/NgX7140ajwCaa/g/x
b94h0ud0G4MimYWHm6z27t7BUCkNwMFZoQQDRSnc6vSz0KpU5bVYQ6kZA3Fg
e4lRWaCssbW3zwTtIDAHjz8ynkUfAoGpCbyN0S9suqaZe/jBHhqD7WwCGJrs
rhIh8TBWMjr+XjrCgWE1/VBzBkave+rIQl0eY1v3uOI6mZlwtTMHo3JXgQYu
WgirfrcDeJcWqa2vYcY8sbPOh6OTPXGSByHiCSTNyVpB/zxFDIhFPVKgKygo
658K78hRbbpe8TziUc4I7IDx7FzivwGz/cVLlwSLlqTxACLYeySoFJEv1tXb
L1Ozo9EDFZwvEpLBoNcUNDBbOLzkNDn3FWEr34NxB6YEF5FVyvMa7hW6heTU
ce+PHhQYWskSJD+iK8ZC08pTUbojZSn///9eKXIn9KgzQBeoSw20DLANcdgh
ILJ7Rqwj7C0dqs3HBMMHLtbJ/oZGVlsL7ip3JaKwbhMb1fnE8VMit0YMpQG9
grcTpqXeTNEADUIPWIibCK7we+FLb2oyx+hUCF0+Uo7FgKHmNlXii4H4RA/r
I23gi+cvOu0IXROEiQalr2EyGLwL24LOo93ykVd5iWkMJDDZh259TARotemb
yeAIfNXDV/OY+61oq7yDdZ53Er4auU0S6hWna2zMc9nw+YOSUjOlTi75o9ls
2lhdInaaCK0lPbdXqItQS8KNXykdd4qyVwhcxYDnnhmX0irQ1zbSB5IrBEkF
pkVym2la6TEGiwQCBvLmYGaexmTCR6neikaj2MckNvI8FgyRm27q1MrT5pn6
RqYcZNG2KIESgOVhN9lYylwdvJdNnL+OU8p9stK5MW6bgG9nbHiFg1c2Rnf7
rkIdpgx6NOSpN5ItQNoXekAbaz7/0rk/7XxrOaIVm6g0VeiYfQSSN9jQbGc9
oMFz2HNXz6gaerS3pZag2PYKSPqDn68UBBSk7Y45HdiZScNKFyvLlmC3OXxe
A0mY1uwFueo4et77pjAocfzGyIicw5B9bpAdn4OlxtfSo0MEh8tWzvbLtkGt
QgmXW9g8B2hZ/j/Mw7GxRudOsr5EzYhvpMkFS1dv8BhJEwwbsTWjvgyy9mQ9
TMZpcTBn3GemnG+bEc1CEKjIexhyRaMGmjyeEuuBpD1knd0SsqsdrWSFCaB2
2cd58jQRR+rMiAu+o9rYWgSNYjXLtWkCeQvUsT/SaQXoLpiCrqVBSF9c18MB
odhkZFq+/hqpT0BHQ6xZ8kBuE2vUN8zzWOprHHp9MOiuRbFU2omLx0DAmTAr
iT4w0xI007DrXjTK94KP9I+mOGS7NA3slhTGN5e5m9EgoKb5CzKcTGIJGb9h
PrpUwsmzLen6KkDzmp0y6LCcAyw+J3d3gxyZU9k00Qq46qbpklv51gaNfkko
qz+gtH/ZdDBcdCKk1nUU6jl7HT+j7676TYexbGKrBVxDXqKnIJtks+rlFpzA
kI+W3cjWWFWmR8M9cFeK8XRITRyJeRtL3zV9I+U0zQmq9D7R4up17D2BpVM0
dfCNrDdpKkIkaEf6zqFgB/heU0DqiZCGoiXTFiBR5txTtk7vjfi7CloPvTZ9
Rt5+g+dhfzwbEWaj/foRWlAcsbWkYAS38piESNmeVVIMhyBFFBz8SEsrDmfh
YzaXD28frMgS2Awk0k/s1XfQVwPq1WQ+Q+Urwqwj/T/Bu3XlL2OijUXSxGrY
XPiNy6C0J12kbpC9NvDxuh7isAJ/3Xv4gVDYXuZ3sdVr6lCOjYz8VlVhBpV6
x5h14BXSp7QkrelgrJqjUdiFBcAhUWL4QNKEJJtZyQ13owqAAECWy5PKo2TZ
zHXDbslUv75SDt18ZaG4T5lgX+qlEtLyvxmtpcsdmRUu3DICR5IxjfxdTP/W
8VFYcsszQH5FP2udqs7yoNSxmxywEqUyW3SMiF1iyBIXxQocLT8m05U6evEz
8ztBk9X9Hj2z8EOtJNMtD/jz2lqZM8BEgVx2N6A2ZNiRY7DSn1j1P5s1hpEb
rNp0E9eCmKkRX/eE0z3nnsZLdC5VgjCJwxNxBTzsg58/z+UfswIsZwJawBnl
psqLtM7XAxlAq1kVklCQgpEuFNDpxG+ULBk35KnPcnM4QPGlp+s9TlK7NQkC
I4J/BlMOU4G/nN6clcbT0MuhvdRtc9cAGO5ErAsk5axdzBQ/cW7B10Jl1yAT
Rg7rA38jVVfCvN/+lxFeH1jJZXuqqAjrf/zNpF4/GD9RgHG7ogZ8QXTuhlHl
xtjclQk+1oNf8UxouMZW9eM0KdMIQHbZTARQMraz81La0im6nT4IMurtlPRP
z+7Bln2Pgodbb1M08mJt2gryEa+lpsiIC5R1yeCtUJmLSkTpdOtp/mt+cp7p
kHrlXnGOzLMzW5DVXRF4vwzo/Drm+RjVyU2z2voe0dfQJvZCT3S3eoz4MV4h
Ma6gzvPAp6s0ZuqqP9zUbeb3RV4I+T+5LlayWRQFCYpFvWt8YoRdjx35cUUe
mAstDALgq9yDOdo+/X1TYLJl3u3IHxglQGPqOvF6X9qG9+zuZWOMcJrBwfqZ
2KmHCRoJcYnPd7ZKmPfQHRtM5Ws+CsmJiyuvPw7Wr/9LFYJZuz5CY6PMT/o2
a0LGzGJmrVKyasDMgh6dvaFYRTg4l1cXwydcGc8zKi/pcxnhk44lI9EmBty/
aMTlHV1yeJr4btImsCsxssgvqDtxdkqb3px7Dm5TkGszSuBkdGT4BYlXFTjB
OuywfoiGBjd6crSn8/XsHtqBH0KU81s3nJWCJ2ymnrCYuPfYM22Rv0xhttUa
UP7Skjmm0lhQ5kPDDyx+d//M/AwrUxGB2ix0ga4LuhnWYWjvhEyLo1sjJgDg
YcvV7cr7g6nPdzYIZtY+0yM+McXGl8poRdlpHB7lVmCOVBs0hwKo5JHzPLFm
dpgDMKFl5rYWXylrVgk49Y/9bsuBK2Mgi0leMti//gEsBkviAvhzyVgvNQY9
4s9Cf3l+aZwydk/Vr8+RGsvG8dmcZv3qBwCl3emarsNx1vTNjL3CGSBhoAKb
tEcJuvqT5pm9EZrldFUQyhxyL99TQRqoVySJnkZRY1NVqJqZzK3/vJH+D7VD
g6Z9fTnqx2oJEiAy/PcfGsTZbIKrXgfI17CvCuN0IlOihE2pZNuPj/oYWBmm
GBm9q/tejIaIwspBqSDXb6e7HxppMrWSTU2ABqKxdE/ZC/G+jWk+mvpXQtso
T1KumrujvbxErQT5PW/NDiANinR3GFDprvs0xvo+OJFYFJsWddYwTWQDy1sU
BnYZYiOBc1pGDDn8fhZdiDSIQrrGjYmSQ4Z/JFnkOoPpO0q6xGSkkovsGPRp
PXMt8tO1XyRJpre5n5TPL++E3ZnK1vhFfWiZKCyajYQ+e9vdetR0YjiUnUGO
grG/s64R2DldSFAj3Wk4UzhG4bkOV88dZX3cCQlMqlraKMk/ldhBV0BJJRI9
1SdSLWOwi6rr5AAqwDFzKxLH+HKKzMk9NfdFdK6MkAyVZAWKF8Mkod4nM6oT
uB1WcGo+UQGgHw91FJoeM18Mcsr4igPWfWcxPLajBhslC4jyMaz1duEjqq3G
SZOmG65s8r/04Jx3EklqqMPvfPqg0fHa85OtKBi4Cw92pg35tkNUtn7h8+4r
Y3jbgfWxV7bOfX/4k6v7hloZjcuMFD4fqGny4v/6aCdy6MhPAxrrF5NIvTIR
LwGGcD0p/360tL9jM8gF1NlfxQWJzD+17CD5dM7INP7XZnbJsmq9BxGk4sA0
L1JwJ/rDkM/SwFRlsXFaF2iKwuWTJEi8H7+CH3A58u3xfwbDa5J7R7FO4+JO
DpEa+l11WGXUFwt94OhPHp6En24kL/s4U2BUN/+M4o+KkL2VyFgrVRnmLgR0
B0G7hfZrkMxhk9Xo7BWHcQ3q0QpB+A+7W5Kds5X5I0daRgTRqUlyHgvjghdz
7g883tKu17BN8A+jWUrtWTEA0HGabtqog70ZZ0bByz8bEby74oBGOrPh2RTg
CHubfzHJ5PRltlCMhRg4gxZeRK7yX2/EMlPCRwOMlWC+ml5UrxCuYg+qA7Gc
ZenDvGFo99slu3YJ9AaR9MKtJrHe9DBX1/3imGuFP7/DluXcpw21kU75Se2+
+dytvZV969KOQVMS95OuFNFjBMVm8rWs8NS3thFS3Ocd+ZVRZH2/2C0TMKci
6gNZW5lzf3SGHvpYXXIbrfQcrETxqFviPca4Abyq3RmsbFZqZ64DLEAkY53u
HlV44HtDuA9GWObK5+ZsG/OHr3o7xSPCLeLEu9pwGSFIOmr1oZvnsl16OxuR
gJp7g+f1tr2714rNvWcNc1gLzDpsp2BBpQwehfXJIZvsbe4YWiFsoZY9X8dX
hwoB4jSfzPY9RDEMI6U7LMtPhD7MeINYXkzPUiHPeUZoWKjBVxP3UFiZHe3K
m6XtjQXllW+L3BLoYlr5zPJMiEvEsrKNpOnflLRJ2twgDGIRrJKxl2Sp92uJ
KrW9wnIbx+mM2Z72W2W05Jjw5YELxN1gqrPu5B6Las0TpcZwNhzba9pXBH0Q
AJcBJpNB4P+ou4qalLhbiRp7JIR6V6LVgxYCoE7Kw4iD+w8MeV3YoQjCH/gG
GbmJew61KbH2fOLgj7H11l9MHQKIBGcRMbFXtWhSS+Bpx5HqumGD1Mx9RXqu
wEnZ4v1MCljGkdQKPMSLCT1ASzgA50tUBLK8UMnzeqs04/A9IuDiUm8dc5pt
ojSUOcKHu/vJMYHoTBjx0dOrs2xrhpynRgWCl4q2uYbK85GePeECpB00rIey
lNs1TvwWgeLsLwuUKhfER4HX+0zg0P3U9rKhflU6yE7Pwkl481UqAy3gnvk4
bwm6uCQHg0kBWy3bh2Y4vwc1ypTXYr3hNxhV+cIC4HU5QQua2gDMyiA5vj8X
MPrHNquQTbMl9yOq3XW0kt2THtZm+7+UXbOHhHPmOWmrcDazH9U2vlu32Xli
0EKqEb+C6koEBE87nQqv7uwYooOBt4zZnNonwIKmruHoo196Nb9Y5ZDQDytL
c7BNbsroRF/slwZZ+A+BBzu0WYeXymd4oey8Npp11Oz+OTyMRakN7qeh0O7r
MTfgJj+GgUJAoYKzCusMKJ1fvK+WuyE9nnCtnbns/sclrqg0jIaqyPGokon8
4+AJh0zimu78vdLtpRKoHWXjQMKn2w79fNSlo7yYqttKDBXdnI0FKxLw0kzg
xMA0BfVrVAcUwWzm3WCL6WY9cmKQFzpTbmWsWkxyx7jhl5yjVTduZqZkGg27
D4DybWCJ8wmhnv7yHMl3azc0MbcvrKvimBNXT7iUIss3PKhpGJv387jl+l4W
cp+YQoVEHEBTCFMtZLUtoE/juClZQxtNDsGfZ/WOP5/eW10iX04PFn9akWCR
xDB0VyXSs6WMmZCNO/VSoXbvueBesH/8ybUAmXEd3kyy5lPnnLrJTDhbH58n
L/KFi+QlCAyJxwXNRNL56jQOD+mSQpVA321/5g283uaGJyeWZPAEMtteq8sT
toJ/W6K9nVfJoE7SkARDH5iAU8a6R1TK/aG95WXfJ4nZlY9a9VtwTeyFJhKm
sJOsn8HYfkdXHqN4vNzKrrTmqdXCB5alqMeeZ/Hrduokp+I/i+YFvj9Ukd72
AZxmIlm/qK/aTzi+/PUNWujFU8/6CfKyX5sDk8EW5Z7WbPtMl0bABwHPqki9
pvL1JMnMkm/kuUlhwPeOjXDVLadU1r7XNThs/P78Pg1lqX+vwYpvRfsh1zFz
lt0E0J79IzAbU23BQNuuiWbhtYy4HJqmPJG37iwRqmiCXlOjRp1zE17P3Sjg
Ya5aMaoGWzhjcJ7k8VlkaVrWYS9G3VLt2du6Dph5YKVLT1UYYttDxiHiO6ky
d2qXOyjbIP0k17V3vun+7f4bK3vzij6SoFcPYSrutBDie2zMmpTuWdgJJxLl
riV7VsJJCMOcCv/+jd0+j1zzTa0G5gMjUnYayfaI1bNrHdnu/bXYZQkbTZyW
CNYXNi897kv8u8vsNjhkFx8nHbDZi+vaG1/t9SeIoUbk+KbsLTwDKfOcdxsY
l2Og2R5CSaJICHr6jUMuB3CbdZ+25EdQXRQIVuNj+hTUIst01B1xG506vYkL
OL8eEzyQHvy1+CvuJq+s2IINUAMCKCnIpMJfU1j7JxoOXPfTrGa7OmSEh7nA
3bHTY+2l8uN+o3VO3IMIiUd5NL5Tx3vHvQOPKLTKYz/bcMUO3W5ZsfRzs1h0
xr26nsQq98//uPBP/A/1fhVF4kvIHSU0dOcp5EklPLUsGFHzfvBnRl1Sn+da
aytNsNW/Pry3DsXc+jJsIF07UpsEjCwKbKE+EpDWRRhtQmZyzLc2rlU2E35W
FTp70bOfG1GND+WyIda03J/gq/R2nx+X4jQWWkbqZSwWdgTmSM/9P0GCN4VZ
lNzfsulTowiMFs/6lIBfA8NO6lPhnrwlNgf4TwObwKx05ag1s6XkVo9QgApQ
cz0keDzVlGWz+bXkWlXc8JVx7349BrISCgUF7pha7zZs+ogP/8JtFJ7PVN6T
nzQb5IRKXn2qURAQoeuKL+vBkAelzRl0C5S7HLir8pI/usI6ppOlYqKI51Rz
yr0sIMCR0wk+49JzB8C1KVnT5PmK+digiIzYBnVlJKpbC5W01s4nASZmn/17
DYCivrBIrh6/fhWDVHIbJdnJ1xbTUdgw7TyNIjYUuzbQlWwLEWUGwpFno+bF
Fu1KH3FBuNS4yEQ/BX1qoqbt7INctn8lYZCES5+OCJg7hafbqEkBhqmgISSw
dWVTTR5+p1haONI46HaAMIRL/PNAkRjS8gfr6kRucdir7PveaPksf1sfx1Sj
z0mCSFYhMJ0z44uWeM90HYZxrdlVf9XtjJqt1HtHN3BGM5YdnVFbSmEb6Voq
m70yxHubs4N8b9JxnbmCcacAxkF/dzDs7TUgqvCHDjkO+tQBDEU04PhSCz9c
74GoGf/+oaOBXX9ASw9hcrTiFAJGafPOu3S0sO6t8O62zPMrhvTH+7x6+2Rm
H4lEgTyOcd1kPiQRKU79psyvRSI3EtZI8th2Ruj3XtdbzkT6feBxbKnrD77g
my0uSV+GXZzdNFNReBYbBWRueQxjzJQ1KMKjm0gtVvbOrbKZvSsnPuXx2oLF
agDYNfKhRE3N2oo+MnFI6HBWhwu2BKVfVrNg5ubSQysegUycic9fAe94YPYY
o7qCxAITCkgZQeCY6HM7Z5Ibt29z33dGPv2A+eyrOGhANDCrOPs2fALZos3+
ZcUzp3Gwds4G6IndSborGf60tQd9UyRLi53+RYw9EUljN7tGo3ShA+F73wyV
bjAHFByzfauLCrZh0fAGEXNujHh+XZY+uYn5MxlPn3b9KxFbjD7Q8cNN/W5r
5EgmDEcaHyntLfV6NTJtfY0XUMkD1x7diYEGUkc7BTGUrLxTKZjpqx6v6OjK
dM+tGclfONLlh8+d6f/w6dkzdJaOQtJfIA+4W62uOx9R7PQWQ9yULL5IGKlV
a6cDtMSz6fHz2uiHQbkxGQH1AO80dgPxz7RcuM17bFMjZsnasaldO0X4ZPeV
nDsQ3n+ojxBA4IcTJzYMnkQ2sx7iI3P/SNVfjXj7whbGHte9a/thyJReILsZ
BIvd+Y+ZaTHr1XiCvla5GSr/7CO2pmvYd2vy0z1JINFLuwfZ1ctnSo+twS3W
iVKjpE45BMHADcaMZkBUdhUVcwg0eI2iVafo+kIkyPxURZSswdukq7Mtm3/W
fwMhx7EPRoOmSyhyPAjqwKs5DnEA3hKRD+PwsZxsqIJ2gW6a50QDtbgEyP5j
Btv5RNjaXYlFO45h6GC3Q0eCKnXrPQICTkO65ZKiqVZjbj7P248OW1/iORZu
29vttUS2bwpd/akn3RbQoMhXQCq3oPyte3L+CjbcMlf/oWlicSTdltXiR6tM
vIrSWXg7GNK0FRrvy/W77QmfVGjQE4eyIG+PYZJVlyeH9llj9lK8AvI21IxC
vYSH7kqg12IFSvRTZfTe6LN4dDbhDpD1/zw1wEdH5YeBDbQnB7qqnWsthiXN
ayYlEII8MgDlOcvjdmfxdJRS/HdvGQTar8uTUkk27EkPdeyShS/dg53sc9zL
FCnA9rZo/Itdsft6IuWA2g+Xtq+wo9re0tkSYdqXweT7SVzYJtbOn9ZW8xua
abJOF8zmn3EjoLiWdTxyRbLemv/RBU4uPaXUSl+xdIjexbm27ZuLUNkQ7fC8
Twwa/2jja6dytE5tNMElsAghBIoiWEOO3F3G3VLQLFR/sggjdyl687f2SfuO
hRUuVVSa8hLW6udDS4hLlcKzy+bN4cie4p4dMjSdhvAHbr9kOxqafgzi7pwn
DcAV074c/qBXlWFQEOuRM49Gvw/XfN0x+d8WizI+4BkBG1hfR3fI2ZwGsNJ9
mucTVVoJb+EiRVvjo+6mnLylz/C+L5wNBcmJeLcp/MT1RGbe+Yq0fwPPE6Je
JrvCuOhAjr1WkrxGDyYpaQoKqMjmzxGh0rJuafLp0mlJOfgE5Ki8K9eVwDNk
49Hwu1ctAAHNG09mVWEv5elYgKb+dgXZfpThHFg04qXMmEI8DvaDEujXRISa
JMdVsL/i40d5D1NU8iy2FgQLvxycSfNphw4HFvaWGhJ0oS/o3MMMH+KYhk7N
ogM3j2rnfwnLZFcx2kzN3nTpqEmiDTojC0nXYc2JOUbFhpnwLXOG3j0sZhae
6BP3YHJalyqhaGntXz6C04vGVwTVZBbkN4qy3jlYkQpJLRvyFpmBy8s7ptGQ
kZbmvsRFzAS19Gkpvm2+7Y5fvZnv4Cytv2u9tjMWujWei8UBpHsSjyzrNjii
Wp8ZHgOr8AQ6LEJ98Q1Ih/WEfxM/8Oqiad8/LdjAq8HyLDf4RWIEQg4NcXTi
es7mG5thZ622PXsvU8EHTxyWLHI1ravBwozJ/ebnJPp05g9JpKcYNo+vHF/u
u19cX8q008WY7EfBYyqeWI55nu43uhya8cV9I7vxPTo2W8PyWCSQEer/hkc7
Shaud/+Ki61NDLqdqNQCnCx0or+m+oB9kIFGHEa6g2rVOjFXMme4Ha39rh9l
1Bwggng6uT4024oUwtHIgh6PcqTGcrbyxDQAaM9tLZvjpiUI7QsahF3KaV3n
jPKkaI9IUNdbDQA+krTetCZ0QX1VRxLyeZhRiwJ3HaTD4WIoAU5f11SS7mAT
6CkzsTUa9H8/lHMt8aWz84Oeadg8cw9qtXad/E3GY/a3K6PK6OXBV6Srvskr
OHDXhnvO4WPHW7N7lRba7S5hiwiGdMn4Lvgyau80+sTFcND71bnud+0sCi9M
bZ17CxS7Kh/GygHshef05lJJY+RtOYvrpLpl4NEm1Gt9XKQaeX2DrdG+x9qv
f9MMpWIm06tWFvim187vhwmlYV1XuLfpfOe6KC5UkYr7J3pJPUS0B/AlUYHF
ywLjGEKqVSSRh7W4XOC4lgkk2lli/RWRb3SdXOmwTqfLg9JVmEBeiu+P5EtV
gW9IG0/ivvEh8piCbiWGFRiiNJUwnzIK5mLeiugSV8Z1aPdGEqt4a4G9i7qX
NJ9ThWMFAMGokBTqdUJlOQDuQudw4yLWty3VDG577ZUuicbkyQn1ZPy5haqL
uOeuTLjaJdcjFQOtGxu2gO0eBpSPyc1v/XD1DWX/OJ60CO2OGb+P1dEnGA3k
WJ5PXGOe4JYvggKDmJc4APWsDIQry7UkpRUFmf7kv3RhMx3tw1+AjAvalNd5
A3TPQN6sCxfECzl4gwrI7iSXJxDY0vMEAIWOMs5zeHon/GcyGWRiwMqd65Ow
7RlzW955Q1ioJyRlNJLjE6FjH2iGGw6k2OLYs3lHvEyy6JGQwraKvCuvG4WV
qXR7DmQSy7LTZHLiueLoM3la9djHyWUtS+Hsf5N3cxNCz400xzAT+gi+qBNv
4W0t1Kh7mIOdKYLunIT+Dvhekz2MhklZcI+3fWZvixMfi4YE/Bx1GlxEtS/3
9/hgzBok5Phtvurju6D/rQVKKsjUflW93LxVuFoG2KBj8UfOSPW+f/KRs3cG
Ti6L1+sy5Xljpt8N1hZOfnWqBIK3wyf7q+jLeTU6FI9M1ArCoL9yLotbpI6r
+e8bPuN26MGPNyzLM11dOnxBAnDhMPPK0Yp/xcZSTzathJyKEtzHeVdzWjbQ
Ii5B4zh7fhT3WuOFw7ugP+01YcbFkOBa0i6/Ley5HIyqjk8jbjUaUe7sNiMm
FPSTt6WfVHn0vR4nJgZ2v22z8Rm9DBFtm17d7X17oHxkoVBM9pav0cp5ZnFF
czdrI+z+slz7u4QtVI46ra+SXktV+BIr0j/0CbiVOdEChg5ZI8XGGjI/ZMkX
v9BZych3W5XIInrrs2MqRCMKY490el5FZS50h+kmQM+Y5UaJ44wYgW1ePO6r
PYivRcv2Uo3x/KJHVdEMnvEzR9IBwtD/O/OY22Vc7RK4Rmfp+310kGHOZQI8
fSJYDols2gPdpBjWdwfxjwo2MoIpP7OjGTxkuz3E27vlppyih11r/Ej+duFc
t6WoH6BpFgmRjOcVt+twcsdym1UeeYVAJ6XwOTwY+5l3jPczAZoATYKOYLJO
6sG5OG+ENC3xZW0xZSTgA9V6KD6sozCBws5Jtb0tqCD67Sve8wq4gZuqJ7LM
68+ca7+9foH3HT2i96vYd2hBFD8X3+g8tShV4pqNMZCXzVBOXzT4h+DlZQZI
T2J0OE8USydC5OjvTGMD8mrnfj1S+aWpq01HIN9t6VcdiHaJfolHTEte+HEC
wFl78jkVbtrISXfua7WQkPLZChsPgpeLWQVG42dnrlmX/XsRhiEQfjJCn1uS
d5G3HYD/Ej8c3+Pho0SNVTJpxiiM8HCTfv1raYXUYU6sl2x1RlEh1NJYXMXM
ffdIAWnFdmASlkoKM5SYEL2NozlFoiTPuBmSjeK4NXQXVbE8Dox3pnfkS+iP
qNLpI7R1yICaHEP5+c1yGEE6lVPuJ4+ge3xmEY/8+NNXGAdHj89FylbrSQhH
DtJAQOhXG3I7yfw9Q8E+vgkIXjVlmqCmZvdROX0Ye8vvWIHr4fthy/lgHozr
HjZYpiaUMcroNeO5g+PHaEQEJ7wgfoH4JoS7k7aWl8lou1RpxERY+8yJdIWF
bsLC3fjlnNndp+fNnTVAmhRRh4pBd8x2gsYjPr5MqJjg47bYkAEbio0rhJjZ
BVSWRKz44rs9Jf/i3q46DyqjcEtKblk4TEaaih1go0cw7EbLz9/D9j+s4NYp
gSmb7XV9450qDAX9xXnOll2IO+PEYSOI6Lz0OU9nI4JM1wl7LRrwmjhO9geB
/tzNm7apY0fAOhbnQ5KicBneuv0oSirxmdZYVS4qgNeUWcYnm1DoP+upLtPl
zQAv2G4gUXeF3puDFjoJ/TynEnj5smYQw0CcKv8UJghSazsXjFuT7rGDeM/6
BLuaWgE6smduVu1O7kP5c/FhBeXzc14sYaTN80P7O2aek+qihq2j0esd4LF8
Deoow0b4jka2/NIzqmEETXvFjlUStxZDmVMD7X1YYf9nb4g+7hxfTV9V0T2t
J6CWCx6rkSsGl1hPIWo03pN0V9L7S1uB+rwo50rxyWp+TXQdkC7kOabJZ9Zj
nLgiDneFsQH3swpzHY2uXqjW5rL+G/1QUQYGFshDjx5URWa8OsuykcmVmVL7
RYaJ9Ykc+yvipb5xDid32vomNgr6y2zyN917jWVk/subpGrUgSioxv+qFluf
WuFPrbUyyWv7+ZKtLIgnX2WvKaybDJO9ta3CYr5hNo8gJEy9srWefGuk3B68
ITARfe2xugWMUlOx4ipt8hAdp2naGRgKHQ8h1CTD3NB825yCqSbfR3kxDO7Q
4fD1zP2qNwUZbR6WOA4LFWS8p3FybRPwaAl+mwUnlYIRPpjQ5b5PcxG4PQne
SnRGNO35NxXvipQY7sNhR2hQkKxuAUxYxSEYLhqnlIn8P21koB8i4+BWI9BE
1g4gmfb6+Cb6oI9c1q7WAqQ4nsyigdvNNkV9S+1ZKVbPDNUf+00CBjpIre/b
KqG3Vw7EUZPg+CgsvWXw+NAtlZfU/zvqd/pc0Pk9ZhEM3JtHi3FBVoeK0SQf
uKYylCwoVzZ2H6GxfRyshE30AvRG7qm0cp7EISDB7RFg0ktk5yUp5LzD7AHm
XI56lSopdHcpXThu4QFq+3XyMKZIfKhKbOZ2elyWtL0PI+6GrUsydXBFuehW
9Hx0Kbs1HLrif3QQ+wPRFXy3Zb6GeSyw2xCeH3oc0XmPUWvLWZFpR7req7I3
SJd5DWfbdd+LWlmf/sp1vmopTHLJdFxktSlB4KAHBTZyY4v6u+uQdyuT2Dtk
1m5VaL8kWL/PELLf3tUpSPl8Rq+RInSEXRmWd8q3zgPsNRa37zU6EpEzOk2f
Z1uDCrqWbRY+bQpIBphD4FV/Vri+7W2/vfZ0goEbjP+bdVarGHW0ICh1gen1
D5HXUskvaKSpIsl18rOCbCBtY2JnlVd2YMc8wTQvW5kPdQniQ4pigCKFAFk+
kyREQG6W6pniUTIWkj4yAdRb2wz3HokHgKl8ppOtSixC2U3eFBNkFYW46d+d
8BGOmtAeHh0FdOrofjKGf7sJAJQHPi6/swzoQnyzRJPrvgTSNLn3B5H68jAh
CpVqCDwbqFrAvYUXOnRYdo158CpW0NN58DwpnLNAp1DMh5pPxh8u56kB5uYz
GOEFbsCBJ3qN/dC8d7A3iTOhal5GKiJCmSPr3LyWjUa6nj8L/dN/L6NrT+//
yOKLIzwp9SRN6gf4vyG39Q052GDwmNw61dIz99S6HQMaMMaMsQmNFVSihVNM
X6H/QD+S/xC2ZV4mnU8Ia0Lpp20JKzMo/fXA8d18ZPfcnET0ZWVaj1iVsHKM
v80jzQ0riFARECgPi/AjVbr5bTZRaEqK/frMSC02+1kQLAbHYB+SGf/knik/
DrwTOx+7o/ilapjzKK50XXjy9TJSAf3RSV36aDj2GVtGvwIRcMb+yJuN4sUO
5/W4u8XxwpGWVQxyD28PprTNRK10t2VcSVXzMaWrwGEg3oYFEVWebEFC0Eh7
6QiJkJO3iFWEmL53esY8Fv8WQgUS0KVGD+YaKDQbIpEW9x0D0Ff9/Qm3ZTQA
Nl7ytF3+Gn1DYkdX9ojRbU5ynF/rPWwi/ZLdiluUqlvaDhx1+VxcG1NsZzEB
+jBNjGiFp8+sDFwdMGdgiQu2JxPbTVAa1Mw/SxqIJllU8yMvcXtXs5aOg0fl
RgsJ87Fl2SHnLHROFxJEvNLYrQF/1WSEqt4wznkcAKtMkvPx1Rmb8xfIYRgh
4Mzf67aktxEAyAuKvebFlWG0MRZw8tB32eSjbfCdNVDmr1j0mXMIUQxGhns9
Vkx6vdVs/o4cAEUu9GCaPOfYOcbLtafPk2SO8OUwC/6cY96gG6R5Q8MpHieO
Rg5KrEsmcBnKkVl8VKwYB2UnVTX1dTVUFEYZX4RjdrsmrbQ9QHngCr8DRV3d
c643YvsDdCgnY28qICay+ZE3RCnie+UNtZBiEhxRdW1OOoyKcT33EzK0wqoa
LP/jVoxdELIbvS1+1Lyz0cNRKVRS1Qs2XunQbXQPSrbjqoQC2WfpRUJ9lN/2
ZLb40Klq+I2oM51ogRwjCEHM1JhRCUgbYO0W/fD0cvSbDbTOfgRTbSy3Pjlg
U3c+qgZ+FtWtogGiFGioRy2fhBfLyyHjE88zgsYm3s6L7GaoKNvmFaxPNDpJ
I5W2nSiSD1CpnIcqjq/4TP2qT/Ixc/F8hq36Ncjav0i9sg2lifgiFAB3bQTX
mw628YFi/Lt5yt8FI1DGVXjE9vDuwJ13mj8OlB+JQNwV1vEip1yZSxGTsOHI
GBGOxtFJwyU+OJMJvyXxo3galjn1w3WLiIrFVt9zZxEvfC1Ce7youh1qV/GV
kwXHTI9cuvIsSPcLf9LeaxHOE+hIhRMD33382bKR5JLcpPtjURv5yt8X/IJU
OMsNzUky/ImLU77gbEiFVhvSzz0yEfVSr6cAm4myQGhUz011YiMa3GFc9sJV
FJiwgXPFziKMofY1L5dgrCKElUq0IEeQuJP0xtiG/A/wBlW696uK8BhejuE0
i10as40FchCTu60sgb3pnOFpTk4r/0Bwvq4/JC6Ffddj+9V39B1VvkvLllm3
frdzFPlSBpFM+3oWs9J37ZRfiydC22ugYpyl16x06RY0nkxmdIXeFTnTpvoy
7IEtS5PU5oCSiOcECpWC7o/w9fjyicR+cpmQTSZQtus5jKGWqdBabLowj2+u
IAl1gSszQmHs5J/VmP+9LsH8eRZJ5ONRvsT4yzXA+0YX6EM2tbL5fGcSAL+B
Cuyzj8vbyDY0UdXMuPFOMx8OdDa3e+l/WX5TrS68t3Ps4uRya3CWPIyvGeeW
ab0PVOJ3GvLvjw/OglxPkXRlmWNYgwaimY+edfuaDX/5wPMXXeQF8ejj4s+k
z004dxJ28MLxGbPmSLPKQBZmTXvzr4x6LydEmbRnO+pYIDLNIayX+KmcxqMp
c5kk6qdLl82qgrUR+QJOpqPFSGFfRE7ANtWbNBcFBEX0RBPCprAiD3OPuvmH
CrJs46d8xSwJCQPCyVj8njTltLxnl+3Vh4IsfQSFIzZVyZu1KUDrMccv/S9z
sOQ3DxVSPKLkimcn1/samtJo+f1YCZK6KRBArsWlg6cnoDbEdvG5W+bS2F9j
K7lkwz7HJKynTdO9GiudyLcYUXuCuTxRliiil9paSy+UcdiOy+XZEL9kcitJ
3tE0/WJGTf5+6OADYPjPte7HFavCK5MpbknuicPKE9fEGK6X+1DmmLRtQ539
q/qiTLk444POMwsDJSIqOx2pgNmTSceLKfqocbtGnbQBrJ9lL/UY0V6MkReq
U3CLuSoKnGxZLuB37mfr9QLdKqjkkrHI4j5UvXXyp+zdpPu/4BbUuV22ieWn
ENoB2FKIU9lywc8izlXVYeBUjyowObvxMlWLk1hqXHetBvIQtzUh3iWuwtyb
iuvRpIo+QdfTu+IF5wThjGY2kwsCrnG7QXha0H22llFDaiGuERbT8EmtjbaZ
Rs0A2H9J3RV+Y+GDNtdxQr0Ojb6Nlv2UoeDpC4gDif2e7QNStDEyuujv9949
IynZtNXxFU+Yfv5iJCm/eUlb0rsgRYiyzv0nDLiImvvNrg3/NrDqhaXQv2p5
eumgdLCwE8EL9Nag70UAlQuTTr2Y3TwfNsVw3T1UQ3MFNdN4KPaxvf6s+b+s
FRQ5iBFWtsDjfMz29M2GNmWmTN8rYU1Z7GhgQgJ9gYhNZVPVQYKDjY0W2uEp
SShBr1qQ+M2lNCxOoWgB7UUWwhkPc1qs9zYrNjJbohxXSi253kYWJB6N+5Ip
wHVIUpyfPNiyJ37GtwuFEaaIb530RbWkujuefO/JBhjDe/n4kj52pPjIWiB8
RjTSRwHqrNJwdtYM/Zi9yvLgFhueaSOzdkhV6sBr0H6C6i+NE4UwcFyBlmWZ
ySNjo6Nd0dGuuT1f7fmwnBGOETG9Q20Xmc4TXPQrmM756tN8Ge4jLiBU0Fjc
Cd8F7luuSQAZwOJGnGQag/2WM58VXcx4bhhP2x6a2cJq5mqfCHiGqc+J1sXO
qaXeeeLRIx6buu/w5OBXNHJ8iANW4xomtr2VMcC4Y4e0ZDHnshg8kOQrUBP6
madTiL8jEqBI1mOepaK5ejK62NXACgnRh7NAgsz7TjiCxPTrRr4DjutUb9Bq
Kx4xQal5WrXrQ9F7JA3XaS1WDUiDcPFyxKy8KzSgBkVW2FN5ULFfW5qV8QVs
Qh4NFhsiZhpNbkgKbZccoybpE1URHM5Eb4Ym2f9mQhvJmgOUz625Bq3vMPs8
DRnzjoClJw4eIo8Fs5lzVGGPok4ne21l0rqVGCYhXzP0RqVmGM+PUP+boI9r
wzqegBQ3s4DlFagnYmLWLUNIFzn1aRD92+G6APpSusIw17b+R9eFgRswFIbV
2IYgvnB2rR7PjOa0snUtH7cPDabzMrj4NhRONf2AYGJ+hfP4DuSjMOTxyRxs
XvnibiFff78ylod3c09bwYovFBpFBCxra8YjXG2pMwZJRUEJYoZF6zaddzVq
LsB1+fUviQdHbsh33PkJB+b8y5zvK04PwnnoWT0AiXmKESkSWFVSjM2IYMzL
jm97hw0wgU0Mq1WqSal83dCTPzwi5cS/w0fxY4klMfYagkHhhQqBRSssw7GE
/lmVENLTPTrZJnh5j3LPRKSGQMK0yu3PKhq3XycClToFqK8EGWWeq3v1t8qL
jkygq/LuD1mKS6nJifmsf+kAsLSRaihWbRG4Ph3AwGMtACKi1qUp9uKynaDd
fS8PrUQo614qhmwwulnPwiz5Ntfa3H5Drh8atxOwgLGnJsJEPFkcxKqLd+9V
lYSg0zskYV2Gh9RsB5nGSqYFylPCvSnW/PhQHMGraL/cMqcb6LdAiJYCbdGC
T+nWmHs/0Dc6KNP0K/C91g/MDRaxI/8LFkr6Xg5PfyCT3BIiLdBg/MTGGrkq
Kz90ZKEZi4Z9MoglhzkRoq7jKRp3loSKWKQwncfOnqZWlNcd7Mcu7lPXOKDH
hcyolWEoxKTQUQ3gLlzN8wgx+rejb4vBoWYOD7MPY5Q+SQ8gVUFqRLMLQDkM
BXrC9f8lFpbEJo3nTE87FODxhKeqzKTV/I3JZn/p536dEplyjEhz6qY7qjvI
7nVNixtuONS7BrDzKRlS92dMHRzwUxZB5rvPVeSrIcoi4tNgGCd+Lf+QrVpx
YwoUZ6omH5WQ0MPTnXkdJzUAjLpqPnBpXt9uE1CXKeL7tPe8nfMMKD21+26V
o69XB6+R3wjHcWYh98OVWDlxnvpuMboTq2/LZ1ipEsfjntr6hWDNw6egCmzI
pPyI0ZNhqC+h498pyRbR4sWZT3xOnEGWw+JQw5SUj7tc6uSI9+QmKLPlTQ/Y
781g2oD6CGwV5wGszrK8yeOtPC8YFwf1Bd74/2PPk/q+hvdJO+enZE0XJTKd
VkC7MSlfKHkZDgprkd5hFh2qkmPhhzuHiiqetppbChs7nm2jSRyhyTK/QlWy
SFL9N53SxsZE+UFvYorU9f3b1FcqpNmiOlXMaBnIdLyW8R2JtMnBE7jpcUG5
uxi6g8cghnvvKux2qKhI5YMuKlcJWVsUQrfFuHllocLDGPmdrzfV8CkjhhOx
Slk+8rRli/xqnf2rueB2yfd8CWy3Rkr+HudvmTEguXOKE3r2GF/Sj5f8s5EZ
e9Ipo7NBVlCihvHdYHdO3g3lcE7rKS8ny2z/WqdbsVDsw2PhSZE+RFhnvPIY
pZau54BBWZ7FNdVhGrCDOG2f3iYjgP12+ORgOwDw3DcUHp4hDBAGVKHtp8oO
LUg0ln1RpKFSWrBZwrCF9QdHUupJCMIMYVcOtNTrr+8zxsNiM7GOYCqM8xd1
yEpDnFuxdftziHju/dVLG1w2mZDobe46GqD8FqYFX2v8xVcoQRKlIqaLtSfB
Ee68XTRMaQRlSvJmh4UaKP+zTlx4t9D22XCLahx4EirsSgMM6Rqj2uJ4z9wz
IYLlxp7c6lXpzmNwTYB4dLBJ2iW6IV8h1TBc9N6lX3EOAHV3TGRMwSVZ67Ko
AU1pn5w92yw4mH/ASDz2+gB6HaKLjP7v4C1K64OmO5qc57H8wlnrqy3xLM7j
0985Hb6WC+d9OZXk6Ct0s+JwelyQE3cfdNdPsemXkMx+Vkvj7XRT1CugkKt5
UCuzyK730hP3YoffaM+EYJv4mOgq7DgshUExS2TkprZB1AQnblO8DKpfJmBW
zGWoErdBTAzkDOPzj5Mo9Gb+LNpfD3ZoRvWshC4rUSCLVHZUNL27OPwBQp6s
wX1cYN0Nh9B2qlp1it7V1mM+Ea1T2Nqkfnnu8U1zg+V/X6pXYvmsmbmcAs+M
wkIHWy9wE28nEaW0bP+1r8ug4t2UzNN3g/5AXIbnjfiuiY4Q+gSt/4qS8V8c
4V8Xj3vWEY0uPpAUPGAQTVkdXBZilye9eMsgr2MU3tDjPKvgv9JGFiYkKdJ5
WBxXjiGRYPrwgDpHdrf9wTrubPg9B5Mlbs+biW3m3CC+rpVYOsMM1+xmX43H
HhcBkMgtBBnsJ0l+pD0qLFk4HTFG03lIcQseqDu5Io4dTCloVf7R0VjOIGAm
pQlDRpTRSHpbKkwRHg+aOjnWyBOUA8Dw8mNynfBiwhg6I4XUkV+3ZLp6zhQe
ohHr57OTmLQHxSJkAl7/o6BLEh0yXkHgm26UmGM81i0YvJdwcB6VSFjNVtb1
tamMohW54UyKWen/vs8G26XWKXCbKn8ZQBVIJ+vLIBMUDvpkMIaeBHF+sxX+
PuJbfxHCAmIn6rK2RFAL666VAYw9Q3/k7TAaudvzhhehd8/vFd5uBLttIRNs
BVndsatLVCdlR8GnEI1v1EJogxaPxw90kTBrNGitDi7JJYpqSJXR6sAYyMS3
XukhIh/e2gHSiQn3g1Af9aWAukk1XG1E9muUCeK9sOUH0oMAigxfMioK8yYL
OwruHrcgXbbIk9+ilzG7dCPeq+HEVdb60FWnKh7JsTdaTBbTLsX3gOoyV2Ub
M3QsWmT2Ygl6nlj+y8kR/Kk9o+JBTwQT9V11gI99+meY1RJsrvlwQjFAObO6
yyfE/SsRYjsAH1e0U4Pq+2Mu4En/0GMZ1d/QYAhPHYJnJg1EUVXKbm6bqVIc
Ldr71YGsZLSizPzNP0lUVY8pzUgGXRKMyH8KkgHTYjudJs+TXxFLj7iObLzI
xyyUJt2dx7jMNWAuH43RwQSeBtZfRJzURHd9A0Xe7WeRtL75qHF84c+RD7Bq
yph4M47nxvR2IjGr84f4oXKJgOgCdaDKehgrm3qX1YrYqX391vhnuYruPjwk
LgG6cyztMic50HAXMRmjXokRV8RXAi4OYWtiasNCcNHLoW89jd7DCPjit6TX
OGbART4vYzefO+vZ55UaOY3UCs9nErCJicLfiHww50ulokOTP/bQh4LnoPEa
ESTQT+elgp6ruO+5v6thP2n+6aXdddBL3Vu+in809gl0jRiDNhADEuvy+PJX
vT2JtLwPXuFU9q8jlQ7iA5dgzYCGu6DNLnRapf0Iw4p/kaRfa0zdCzCCoMez
KTA5saBB2rUJf2OGhQtUt5eM91DCaVM/Yg8I2tyrQlYisIKi+WPQbsuTit+P
NZPortVD9SSs8xuoBDPZBYemLevfAfNpTIyeHURz0JTk0ktWmBa1P0G9UFm1
gLBRpD/v/BRyQumwQ1vLo7PpNcjChINl6g3OxQjXFTvhSu5vzpTqfLlLPMPa
6Gmc+KRl3q+0xUmSyyk4JSdyIEYmN+mVDKPBXrtK8ndHK3Y3zIcGYLco/1KC
pUf9BVYKhkq6vuraIKjizbDlD0DZZnIMIEPnIXZR6R6Op2gPxwKc7aoSz4Cq
QhVV1GL3hKE8ANyHg2W6I+EdhTbyAicoUtxZKVYLf6njNkdtkYnEIKbYqEvX
66DkJSW/P03QEZnCkIbX+8X/H/zKM1w3wd1RCmSwaaH1DVJC6BUf6WxxSSFJ
VgeJw987DsSpjonfcqLGJWxsbszRYtmV6mSdSR2YMVLr1s8o1OVio3b3lVcs
bor1TVgfjiLrQ0JUbZWDEZx278LmGfD7cn33Ln5EsZcglcTHqQTRxvggnj2U
4AL0LUvl0i6s2tORZmDiY65U+r2AyXWgtpjM8a22r5UJNLW0eozOHi8rJuTO
vTF3IUCVLEAAdDb8hX/W1hy7MGWon/H/eFwgd4SRwo1n10DG2+U4PyM3bCo0
IQl4+ubJ4HsnPevOaOBG5pPccTv3RYQPIfhu72JK2XBnFNzPs/4Y7I1nteLa
hKIJHouOy5dwWej2CloPzP+nQv3FRrMVn7wks7Pkm+MCu8LoDy8QvSEsateT
hQ0UZ3c8xPibrrc8D4WgsopJc/vIy0jaLFgPUjUTQlJSMBCM53Vgzbn0ZIvM
XGzm6u49t2DDLUBOVmzXCo6xmGqnLb6qmgX9gMsx7l0nQxyPJf+xtFdVchK/
K9SPiOYZb1zAK7Fjs5a8bMA5Xetcr5h4Zhl+t8t3EtGq55//7vUIFtVBA899
77w1tU9eAxerxnLXgzNuR88hnCx21u3xPxE788sErMqaVPKp7WtokmER350G
BzGBHGQivoSBOR/wa8KekJLk8hJMxK5+SBaerEzU2xtKXD8OJkvDdxk1ta3y
04A/4+rrCS4u5rG3Mb0Bpk8mnvNZHrS17FS403zDHJjzXNW1AaeuSAmyiJO6
Lcqh8xa/oe8jpiV8Y51PwkbN/r+oepFMa49WBayucMWWLspHLMiKVCyBl853
Ofny6o76qP2DDxBYUDTU4RgDkkSOv6LrtrztZyhnJzkJSRtbs9gH7Cu+M076
Gjpk4gqAaGMGIYptOUmhQpzbSmqyFch5aqQGfGct3zn1y3M5fzi0ICG/cAXM
UFVhujdz0nyIP2AONHQ9wuELd4S/5JMH2QvlRweXh47LpIuHa8H5goKjKw3F
HA3GFpD/QtXhMp1wghNNp1fERjow0WrNGJ39RbwUQEEdbTNQljbucTUl4WGW
mjDVFw8AeLxz/XAnUv81Xusim2sgOh3e7tkbz/nzWef+F/lmTbrhsm9bvdZK
N8/YKVeoijc43whDxKyUVRTAr7tFLmEjOuYJvLpXC/eooTPO3JcejAObUmFS
ruS9GQVEYS6UqP7p5TqpBsOVKIrk3VidJm/jyqBAF59EBPwqUS+ZSK7h62Y+
In9TgWjF0nc7hGXh+swq3a54nYmfa8nDEW+sa5jHxJlrA/ShMBvk1qG62ENe
Yi3z5Qldmhli1nl4djTFGSlBsBNRxPTjJmzyu9sSC6hSHG+hhOHDNWXFvXSW
zo3MzJ/XNnfToAqaFJC608HGmeC1IiZ8qWqqWv1rUwSOrSID9GW05GZ5T4/Y
WmAv/8TYnQw599+Ohr/lvApoZA7d2T8EN5qW/g8duGX+npJElFACo3VubWDV
boReK6PxIzA4rASMBgf36BUJmkWvUyxhug1g7zX4uEZ0k7FJsNgn+yqPAshf
0cqR1RizieyLqtT+piQ8Hrs7DKMNtkzYTNOLypGSzY3LIwEZYqKch95v9yaJ
78t4CYljyX9VKei2y3nAe3ljCkQkF4nj5dC1wvh/ydnAG7NauabSlMk/Hjgx
+yPz1k1PhkHPwXCvkjwynuWp+u8fFD82Tt2VrtcQBmWr88DYxddJaf1wYdeT
RE86UD5LzoAuBW+fjiXduIcNlVpwXBKqYR14EWzpquhfeKO47xuvQ3tLF0Zd
p3RiKyudsXZZ5dUjrUC4GACOxEJYj335tbRCjcDW2zbNPmyNsUd9hMEjvX3c
xhvuPQ7C4zt5gqZnrAfp/QMqTpHcuNRFqP8hIgEfxbVJbNk3Puw/WpY1g1f/
h/zHMfRRXgp8p9U2c2/7WyyzvUCKsaqNpGc2pKEZ+GNaqtu414xKfxaN0WSf
UyXL7vP0omcf833REqZWKawFcsrtywpVP8h3GeGBpbkvgNUBtR/1i0rOl7m5
HKkPSEuDISWPoJeS4RIsaMFVfO44rfAzfFo4Bausu3D2xCU5RzbsPOP5owG8
/HFhI54OaNuv/BUz5OFh6+8Ujf5nuemQ+PAFEG+CBSzRyzEpHqSu5w9q4XGZ
gQcnz1oc2GNGvRwTCm9BcQCTmS9rjrIJIIb7rdpj6lOA0u1+qcu+i5nb1Lah
KmxEGAQMiUeasLvBo7kGXuZ5Fwz61wHt2rKviw5GZM/C3yPfy45+wJ8ezFNS
l8YecZCQ7VF782xutX45Lf8M0s25ZPPGkEKhkLEYsLlTyq1kBzi+Bi7I5kO0
mGLZNYN0+DCVEpWR2LWPmP0aA+o0y7Gx3qHecSq09y4O8R3XWw8Wi4VredrE
lB8o5lvAvhMJgQz0v+vWF+HEXTQwRphu6jZyaXTEFV29EVVgkfCGoHEP7w0p
gTDttz9WCzENKCh3lgO9nGaa98E5mg687ZhoiVZrCAsHR8bIPPij84qtjN1s
00fpj5vMNnDwtH5xdP4ZoI7Zw2VtfE40twQkmMTP4j4JkGrrzFy6eXVyosQS
IN/XdXgAteIt6v5NfPFfpTWA4gJdNDybatA8q4KAyehZHOadCyFd1XXJEgmu
HGJ6dZh7WEcDkyWNoYQeSMA8Mw/obgTftS37aHbkbbPN0VYGKJ5W+aqUavuC
RlqidMIMW1cSd0aC7IFEWkg6Bni9pHx5p95VSo9C2g77WYlqxPvYNy0WUbmP
x5OArooKWiFZd2kTA5TjAl/U9Rg9zDJ0fGAjxbbWHn4fmXf+jGfeIbpolvNo
+AINnAqRFh51UpO9UO7LdvYqVzl/FzUsTot1FfyAqpF24pAUYSnI6t714+ye
d7jT8E3rk47zJKtuLm5/tM5Stvf9nBOn9i2/UJ1sG3pjlr6KoyOSTlEW8nUs
AMmUqYfS5uHFw9tm1cdzqlLRDu9e/fIdkR8n7VKylzhQubaov2yztP4Jj4hI
W6d9wLiYuMwrnpmvr/qriImck+XoG2+NrP2P7Yy6Qy/7VTMVdSAAjRfXvkoz
lHVm/h/H+Y2pftGfIfftLcLoXqqys1gsbx59+WMZv3M0rW89omaAgHebwGeT
8w1Jb6b8XvhJ49CftntvnFDa+l89RnMI8TLDXh5knbt3S1XwEv1O663YZfQS
lk2SUTbsvWDYJuWL8KR3HeAHOsw76+nXDojDRe16kmnFLNM58HpomS5MFyK1
apWfygf8r3uzDhLuvrf3+YJLU5z1QaCVJrnQs46o+eBw9w2VszL3QLmQpbb+
IqucoJAgJz3UmYAvAAu9ldF6qEwL8OjaIOejInFeuPctY8TmHjjlgJLevw/I
zKOGaEeBqtOsZwxYwuJbVyEF2Ye2fR8IAjl7wrdQnFJQLyq9y3oBuk35aGVC
rwHwWtVH8up6BOOtol9vgH6kmucVUOl1pFfSit3PGU+6G9mqXYeoGMMe9MsS
zjiOiHlQ38+TFxJXZqS9fBHabCLJM0DPjPiNeQpxSex5jWEgooa3ipmgSTsf
esmyg835IJv9mw0Xx5+YmZ/i9S5E2G6C0ZynXyjpDQF9JSjygaQ3cg0S5u29
xA+qrtb/J2I0Ak36HH84d8x8/FGnobkkQuBCibVBr82EhYEE/qFtnklDgrGj
rGnzbqdz941nv80f9wPy1Hvv7Vyxvn9k6ZnEUYy/7kRa3tQzUGcEb1m7dlYZ
LFtchIWS8Xpy4yGIP9L0UtbzvVZ43ImLk23beZ859YWOOYElU+NovzhGGmbu
J2nQJUOQRcUBmNaekRtMWqKSV4TSEE3mpbLJsSd5TQI+heQDnM+AawsxUEFV
cpwz+l2r74g94uKBoXYatjs/+zmlo/tVRPAaiZ0w5YB78t2oEzXmkMY0lc0K
V7Nzn4jn8od0U3vnFZirv4DrZJdrtA8dOnc1qnUgHSs2pyzr+ddLsh4RLE8u
N6Mzs6nzZ6AtI1mHOcikXeWwgaAc8BcGTZJOqmHznprOfBAXmkT6OK8PKOwq
Sk6J1Q6VUDn5/Us3fkJecooGYoIx1cIBN71Fvz8zzCoNofC2EAxV8JxWJHvL
COMdk6kxfDf2su3yNZL23iJgVoaDHcWWW7ibCvEGMduSF/nCrWH/LmgUWXaB
yi5KsPPSulXNgl7BjJanp9bsHTbaMQQ3uzx6xksB3ymSn66Djly7VRJG/CUo
74ZSqCsTEcFVYjusC5PbJkER1+c+du68Bd8ZwS3a6zrtyaqz+SmYfjTK2ffY
KdMLm/4DWLGk7IWGMCqzbYekJEj75oNpPULJ94PyHWGLc2REM2ELUEUgC6Rl
YBOqEaEo7RK7UoOIJ7DzLJ4LFvtXXN5gYv+St+sRx8mdKOH90wrGeX89xmhV
CEUGqmhfrVPSd6VGCZ/rhd3yKdrrcJbu1EQfDspdXK80SVB2uySCly8k3LTg
4wcRnncHcXwhLHFX9V/Ok2+S6bqdi3ayVS4/eU67PglV3uJriaef0MCm1Msn
+3pQ1vYdNeOuw6Z2x6j6m3BMiLqqPIXsTI9TNhwDO39LTI4Z+I/EaJnQ/Mxw
PL1gKcLbaD+4ZE/GrgnKOH4joydbnZ1xsEhH6Sn/WavhbISujmjmQridOKNm
BrNBt8RRW7YEfivghq0LxWy+OlIwAJ+Ce5h0dDkTxi4GgIk0PiAsSEpLY6UL
M9oJxsZfvqyx8ZEggngG6+v4veHqC5OKdsfGZ+JIDYLUpdrHxVI+94sOiKVF
HCqJFE1FnSi5/aiO43Cm9sYSYLtOeZHPTon821LFF2ZptfHnJNdcu2UyGDum
OyQZLGnQy9MUr7VGHnIvNSZV8eL3I/yVEt+8evW8iPuL8e0HZabgf5v1eJM5
Z2V2NaYuXpkZu+pFqWZAeoGUgLUfsakS/jNsFl+ToNwEkPQeV3R7ZQHNYIwm
W04Kdos1UHAamHEqtoADBvchyI0UrK6Lvji0PGQhO4ZIlZE1CZDHgf0gQ2pX
we+J54SAtITKU405Mkui5TNgzYPLOPhXUR+byal66lEq984DPBb1LhB+rpVS
tDoklX32rDzqEcMbVJ2j2FhEprPf29NAW6PODg2m0PUqJrkNm6tnSOZRqbH7
lI93zhmZeBz2HqRiHps/MqPlRuBibPgZOVnJC8QYQeCqpwxUwJAdLtdBadie
3d5cyOGUR1RRtgNYs93vztGc4gKZCPw9pJn6U8e70M3jWHZLJhdZEWZA4TiS
CQaSrpJTmid2HqTMhUr4DJ0QLMEH9F3q5x/70wZVJwCCvQsdGFm5whj9uhI1
PQ/dBx0bl/E0F27G1xbJT1L7mwAtywiDJDFbcDcP0OAi4LevqQAascv//JSz
q8n4swKYGDltJD0xQ+fz/RJmajbiX1s2dnI4KmYSVdlxawyvUyt9/tE5Jw+E
QLscOf1Y6sK7bkLWx56xMBgNfsI2BX63RjLJ7LjkDGr0D5uybNmoCGPaqUoa
ki2h66amR26phndha09eF5m7r5VBJVz3LALuvpXwsaEEfBKO5zlMmDeCoDaw
kdh3g0vwZFwsd0pixNDJBZMtWv7Iij5hAv2H6NzxaqZOd875B1Y9Fe7JpLMH
kyZqEjNHxhA3Cpo9m1dpkH5kuKLstkpp78fne7nP80km6HDI1HCjIRHcQKsv
cNSdNmZQebcGpC2zk67Z7kg8h05UAfDAXo3ryienCPT1sCjgnHqLO8WJPJSa
GNM9Z2u8NjzUYLg/nAUSgq/97URKc/iGLpwuibnrJtwlAVe8EfKIYopzpBur
Pb32RNDnCsM2FRbOQMzt9Mun0tRQbzs/NRuE8mjtPUK6io6Gnz69z0Qv9uPo
aG6MiluM22g+GfI7bH1mexp8EInYKQO55oaDiFShWb2rMuI3/tK/zshbq+hW
A0XcuJj6qgzWS5WqFnmDgHLOglaVoa0CABIxwSkpomA/Z4WspS2OJsVnML6n
S+eXai2rVUP44geEuQhUY5qGFJ0oHt089n+dUslqB8A40P4u9xKvdmcHXPOE
Rrr1rXWsNBlYa61cp5SklgN159MnfyYNV4rky9pI5HfaYJJaDjWB5rjag5iZ
4BvK0m1JwOYtw+WULgsZu18wlzjyKFbF+L4a/crnw8PuxfupJicBF99WlM3M
6Li4GgdKRpi9kMqntZkxCQE5f/Z3jgzOZmXFncDXbyffPhX5x26M3xhRPZ0m
cTBPxuCI+YAjjO1jm5vHF3s0hVdjXKAASOhvc0Yy0MmP4UZ8K6WMv+zqpA7R
osAIGc9/d5vO1rmo/DqZdGopPfux++iy1/25E/8EqLPn6KVNhAPrDiD4GclD
Ca607CMv3TnBmKOBs1CFruW0y8dBGgeYbverGtB/62Zje4iFXldhYXZhzZsU
oYtOWVCGrBaAgtNJWKDJ1aEl+Z0X8exU2IXHaIPTDlAYBHTW9rOYay8KWCdS
o6nneV6DHpiswYD2l/KzfzygZ08jaKQEAMXeWSqZ614NZJBJEvBdYLI/+8ly
MlXobbHBtHJKWJSNQhe3Cq290/AxJII2GQGOF2cCLvNa3+GPra3AWGpbRscW
nL8b2ASBt/WEHL3weA497vMJS1BI2EoxoVbeTcUcz7G0/G4yutygVt78a21H
6ziufDh2LI/9G6EeiNNq4F67HvCASnGGPJyGdXGdbmsA/vqsm6DuTiltxX8G
pmAaMPmtMgu+2kTqc/xftlsHLhR24qQcE3ILXvdiPBXlHyRb+bRbnFbahz/H
9p2trRPvTLOUaBOGSCcosiUU9pTB9q0HW35cJUbVxe1aAJXeMhXJvWv8SxX8
0mQq84xthHzruS5ixqUk6LlNB4XtdKhFKsE90rGRiAnKyktNiTsq/8Qwdqwd
KU9C/X0ZnKnIQ2N3HGQ3du+vkmW3rKLSTa8vvIvGsnRkQUEgpgSKDZzs+7r2
2vy/LBjbB84SPMWa7LmnsN/0feROAe3AuYEHITm/OyhfsPop9DHIKze/Dug8
z5SAO2ZOFC/5byiazZeLt8Q95yVfg1a/nZMgjYQ4OPbO8H10lRd2aWKqnCiT
NFsqu3lguxEI416Obs5be0ku/kaulRlO6FmhsPBVlNwJpUNXqFsnejRBVg01
mar09xFwkBwZ9oo6NlI5bx3tD8DSXyARSDybzmcahHzTtquELQKJ0n+m3NqF
iPkV7qv3/C5b7/vmtab2Qhzg+QHDszdbm8aAveuGLIBjc23xIzFIMnmb7o6A
pDhizHFiECPH9pCaV0+NVwMsGcFE5OOd7hccw56H9f1eHSfeZXfJp+fWsxVx
NX419ebcanGsJikLosirPg0A+Dh/xGPWoVrInv0YBboFn7fkWAAQRm3RIfuh
gqrCzsD3pjpoqc0yUnKhOjWItBGeBD1RxqmUc+UIj279K0o3wlTdRoAlmQ6B
mb8wyn0LieHyl0QlXpuMl/Y2+i3SjjONWtXaYyTj//ioNNV7JvB0O2/+2Nc5
QOIzbiADqYpG5jMYkzTZb9E/UTigChQkskecX1MTNW4NgSsPxGH97buOtGEP
S8C/qltXCHpWjHS3h1aMA9Ivgc7H5CqufFVkThQgC8AZM8syOhEyubKZRBuG
0N6IxfzT6p5H9CBCaJh7BnQyj7LornoMzgY4V20kgyC1J+PGZ/7RNaTvmhAn
yad2YECRAT4V+WK59M3yxc6w893nCk1DBg4eecxRwlz2rngZVWAnTy/9EwPf
3BTDYneLE5pZedmsTEf+S0tPsRBesgB3OOl/D0+c8+AWc9zuW6FHGc83I92d
GHljdepuIlnuP8QQUI3W1gTiZY7yfEXq75SF6bvRCF9/F2lDOXhWjWYgnFXU
Y4LEmom68zoS//gw1oJQKwrvACPOaQUPUoq45WPxA6F0sQFRs/dLSZoFLbKv
LrXc7HP4VKA5JxO2WMo1Ah8NgdpYT+ouYYk/TRNDtsWoy3hkeg1WFZnobXdo
8MfnJntevpPBzUbF+WuOXDIjC/EY/Nr/A5sbjLPuOkTBE9r1vGNj0CLKjHWW
7cE2rjl9KWypLFvYbr8dxr+QzH5EetTnOS7RxiaHRJ7ZpzcKjE3fAPH0nnjW
mdXP8EsE3sVO5UCd5MAqsi9Jgnke7C7HBZowujQWXqghpsEE3uVD/Qox/MWc
UdWAhKCWlz9sSj+9xtIH7+JZFiQoSETwyMxWgdLSbiSRrtqYPrW1afzT47+L
1GZ8Ftp61I/KOwm5n+pDmHoW9axLVtxeANp842huidy54LoC150M/cNW0Wf7
MpQKBYH1fieJTqmkBpuDQcGNrmvgcyTKDhu+y/Md16wkGQam0fz5GAYrGnuk
TqwXQ7wqUgPaVAReLdEnzmyeQEBHcgxwL8umalV2XSLPhgStUbjCIHMaTCv/
wJK6yvYE+0OgtIykC+uSd9V6B9fT7DYMHbpI59tHvp9fbgcOsLphilljVw1C
1mPEHuTZiAiYLRkaxvcBr7lfdeldnU9ZeGem45bKnLsqOIYGixH0M8WC+Dae
S9nKWqZV6jZlCL9Q/Qk1qqfjy+j4qOWuIXzcNUPavaXnT5EeFrqjp7KMCH79
gOFarQciK3ptd9PQ/ex7nqYvWjPVkvGAmzrNiqH1dEmPvp1mLIFFoVCQFvm6
ZVd4vf14xLLarSt7IJSOd7VHT2RS19wOn1/2HFgxW7LtEE43FcwaHm5Ckwq4
6ZaSMg9uyJJ/XeeClJc0R7y5FwEGkeJWuwQJQYncGcDW/gowq7wO5ql0GAeu
e04GFic5kTvsrAAJ81g25UcIhp5xMzTWm0esH4N78ljfyc5dHpuHeDxMXjHs
DIn4qDiWbuqMTPN5cxBGqcMq2Y/wJwoR1pHITqkHovkmvrcjwamF9vOU4B5g
Hri3RPi25ytnJjWv87JsHTtWQbSUVHe8E+kgdO2xnVwFYJuPIG/mPKKkFaC8
tVw/p9E4sIPXYyh/ReHNYqTDE9alBAy8nexIiuaJsB0fhoCT/9pWpTal6i6N
ECd7xnlZyqsxKrRmMCrCqa8NtUZ9y8HNk5mkpehBkqJIapGc/5TDBvJzRGkB
n4jBLTp4tVRK5pOIagiO/0zHuYZT2mlhda0PJfcxlEWJo1UQyUImCKmgyOrD
2gUsKOU2fmfFYb60MAXrUGyUdVswlTj6getTh2IMwxC5wHJoeuO1Rvd4TnPS
PmZJNsn+fpSUFI04W20/rjrubVoMglDvmlEMDwFQlx0RjSHv5HjcazlFaDBQ
Jn5crPeV07vJMX9o659zgCeJuc2c7d9QUbXYdfICespzbWJGxCL9IAfmjIDG
afyGfqUBZeNyROoflS+fL9FFM3x3Jv4+y5pnIkB5AWI2r6mHkdAmR9uYFEOO
JzRrWEnQG1pS+bLCJ38DSFNFY5laNrclk4zXOTJFbqqC3wfBEF0iaDgHYEgP
UoqJMmnTPYJ/pCFiZRpZqypR1Lxa3rzQbCxD2t8ya+/U5ylZXH0prUr7oSIw
rM03rIF4o1ETRi2MF5QTKmle9nBshOcXmRb+JsLZRtdk29uWtBFvddZT7XPF
cKIeLD/WAaSZ7j9pRIPEnJatC6AeSPWg3ytsaHUjEKKSRiKztnoqGgQFzkE4
2GLMnvysW7w2RzGMOGdX31OUwNa1nz12nev2XExVsrNpDWgEZkp7k3LhQMo6
bIjtZKVLqzKNb7tuOzI5CtK014Skr3CNw21BJjYCeK9TSi7iMtT8fBU1/deN
/VKmoGazkVy405rO6szXXVCi2w5NisBn1dMM0A+iqziTQzfOM1QKEA/KnPpF
cZ3RBsbU4zgvQm4j6TML26p45KvjwumvYwYQdoo8k4vH52KYQpUb0dplwB/C
233bEWq2bjhCoz2dQSvRw+JkBzrbaU5VWIxn0pHqpQZhgRUW+CKlvpy63vc9
C5ixT9e1tJHvKXiGVss79mGayyb9rJ1CXoMgSEIDFDfTCa068GlPcWvC60jl
TXxY9Y6n/pQ59UnXl4YFzIQciIB3cTqZikXlDrVIZFFXALwDvTspCdEcobHh
TCXGstbvyhiscWkJatql6Tf2nAUmHsfIEngedb2u5ZDLI1xA/TrE2XwgOoaY
gTabS0+/PpwL6Ap67JGpo+9CMDL6MWqus2GKPsmEz4elqm/ytllQPu1tA3Pw
95eroJ9E0q4f9/50N9u2lsUCA7DzK8hzuM2jwtvfmDGSOEiXEiwgEh2W5qpc
Ldp/TxiGukk9bUttySLW3U64Bt/ngvBSjIN2C0LNDkhTu3ObIMS+rYQnxsA5
ePk4UZ79Ryyvz7Pc1UHXbDu8CyJiid0cNvH7y8yVxO1Ye+G7adS6ZRYiGkYx
rKFs76M8H4ayfE4I5msD3b2oYM6mbC1CQ8UsYWl9IztjNwjuYZ5N0Gy/QZeW
sF9F09elZL8rO+hF1ViSuQH5mr8V5xCXtNWkwzlAAxVpOaLeXsGFXuCvATT2
TVob6w2tMXQMdXpkrhu6Q0ZvBU1Brw//gGdoQ3sNUv48U6ZPpnudLTuUa4NK
m9S1gis4kjebqd7zlTCumoRC7g+lKYHgF66RVDbsbhpH0fAQIOdQBMrs0NSN
MyJoBzNh8kFjUtP17ATgkmj4NFH5hS7zjJcnVkpL9r1Kc58aDqeLO/tIRHDe
sT1USEIFOaGxMyFr4BJxrKCMYTg8ueNQTAmSThmI6oXWwCJRrkOj7TnicIZr
NrPFYXIGBHt7nSTkwjPoCMVgcAonlXuV3DoTASpctLQ+2Xlx4C79sSBTvM9R
66FT75kDpfwLkxqQ24YLSH0aqvzcUom9Hy0vWbvUz49iG66PJCoMBoVXjDKC
juVcnB8qKi5fHnXbc0Fwo+0AYfGjBABEuN2zOcml97ONnKOTK2vdaHPK/iBg
iZ+pG0br+5dzZrEafFyzf+CmE71ezje3H9gYqgeUHsUbeTscGcIV/twOm40N
DCocXLi3y5xNPAgoSkg4yZP67NJQaZ1FY59ZGlo/utm2G+EDsxbUEh/S91Zx
8nygrHoDZraekl00skcOBf50L8uLst/j5nImj/mfnefcGbQDCAu5TPppi+/L
U/494yiO2RnVkLAhS/MtXB16uzLcFcdQX4BmnUbiKb/EVcfI732cq6AyDz50
VzYeKEqV3q1aOtCEG9nNEWwHsC6s4kB9L9NQv2a6KcSgMO973LPnPXOWknu5
77HLFxnM4vO4XbfV5fXlcumfhGvpf07oWh6vKCGutV1eynbA5VxFPSmNPlt5
Jw9JzCGNdBAJboDjD8bfb6U3gK9jWEFk4Uc4Pp8ld9ScJvX5qwCjpfxGJoSK
sBYRRPrL0rhH1FfPt8UVtjoeIwJ5L0z+vFXDrf9OJxgPXgPJ2GiDYo35Q6la
/0lP7tLzKabvWSOxJeUPtRA206emF6pko08/kYK6Vw9TZXpVlbLAJawVEzTV
3nBj1AkkAsOHb8NZRANnaXggrh9s2fUeHOeeCbdrgM9Yrv6n4sg1VBhg4zX/
I3FuwIdWN3A+dq2CI+SD6ObhPprgZTUzXNl2RY73Aqf3KweX0vyL8NXysEDm
nqCUZtckYNC7Lqaf7ovNFY5Z6JR8kKcqT2BeDkcY1dGyL2x0ST6dCl6Jyl/Q
wZIOtPGvAO+C3xnp4Bo6BxpMB52THO9NsZNlGBjTgnFGXrc0wmTnwYiZqTho
sUC53wudJ5cq6G72O7Z13M0+kfmp+9iJzfu8zaq1ZU6mo6y/SefUqe6TELY3
bEDOIJ+Z0xcYkbifN/vbshtzTAcJWimcNx1UC2xru2vITi/G90MmoZ3lUosr
eDEz/W0OZ/zjSbo1QdABZDgLp9m6iGHBiIQnIHz0Qn7bATJnAXwFI7o1h5ju
YnjcPhxwzCRLFSzqW689NLG/stKBlHc6ZUubhrapLfBk33q6AyhFYuvRlS4+
ZzCsOwNUSj1FJ8a+8d+EgpU4CTOQ6BgiLGENCqHT3uabZWDyZe275qy8wRvN
UIoZK37RGOroeEIiKhAdmPd6NEh5cmQ0Fvsh3bcz1haW6N8kusVNzRSFJIJo
7TvqN4fT80BzQp9jfbY7YQ5oSROGrcyAZr7Cd4SBPyBKRafel9xivNMGTqMl
/qBjzkWThfW30n3nxR05rlemSxdkotNpVtsnDhYTW/PL79G+hR9urhrlzKPQ
2tyMTiGXLQBqeIZiCJSVC0qqAQ0nfVVzwPuEiOEaHkPGtDTcX9QNQbOEAwOt
JC8wqPQyMNkXEhE98faihaabD6TsWJjlKZOmwekuHoTzESMPb1ocVGj4cQBz
7kMue6aXwHT67QgSYbilvPXEhc/UsvHk79P+tj8ChjnjayCVB9BGwz39HU6+
AiJVUCHcb4DkbcV1Ceaf6pSu/nWkbR9ZKEl1suZwupsCJgohiPDjCw6y71nB
uHf6g0uW7g0vtEyHj+rOYE4r8tpjxLI/0EJxmKULbl/ZqsTnA5QXEjSJBTXH
oDNkkTm6w3kE3wIAXeQwz/ex9gB6kgun4RzZL8J0IYOJ2o4POguAld7VxneE
HRdk+htlrcRHft0Y+WAX2J8oWWhsN13RJn1d12M6BscJMNCCK43+OnTnKrHj
N2Mt5b/34TEG5fxDEYEWMPaWarQicrDMWMIIvUP8skW7jRpc3GE8RpwbsW5U
xc7HWX+sYiqXqyelrJqJWoKTef7yWM9TRREvhlj5tvs51BRI5diAL3RwQhwf
MIt4oXbKKZGqiNrBvYbZN1xUJTsVOyNsuHqyzqTkYn/1kLma+OBS3QgN2XLI
MyZAFQWvC/JdHMGpVdwD4WvNHm5k1QS1ZSp8RlmoRv3extChEwrpLWIlA3+s
29pxPAeUf6wuxqkABMtS/YAQQ3GQVapkCQAe4yWZnRN5+iyZibVcOSiqKj9z
Mjc0mV2xiUclUDkd6tlRZCiNRebZIcRSjW5WrGW4E6zEUTl1g88RMaS8MEET
cofm9DuZ+OeWxvfu98FPrYC41YSFzg6HIpwfOfa2dtw9rOA3GmyQEt/IhFZV
fll+McDMnlmTcOfBAv9gU0+3ndnNNm1Co3nzcXZPELRCQFjheN88YO69FZRX
j01ak5a8U6HTGkl3rTLo+/Jzv3Ww+IWxRWzVUBilNLIHWnWOpm1jRN/8SXhp
59uDrnS308qsGe2Cgqv4qdrHv6LcJtLHiI3UXCOjBH/jCeKaFj0meHpBGbsu
AefF8N1myvksK04tWZTWdA+MZIBDXCD/4tz3vpP+eDQfk/FVkTltXUcrlq8P
SLhg0a2XzZKjdJejAKgBjsjrpxFNn30eQxFHHvL7LixRIBY3SR6yhYyWL3Xh
NLQra8Go/wfL8NKIV64Xd7dgBkpDhOSLLwa//siznVxW2ydzg76OGxLUJ21j
4w6dWgLd+G36SQseGI/bGLOCagGDipMmzHyA47iGmFGtlQmDEpq8PI1lbgCV
0l2CrChFgXPYWs2TXgUg2Nn18TiiyzWeusm9ydhBMDrzC7d+KJW99s2KNQM7
m1QLLJF5M/D15Z5+YmHN1aMk+kupGwpwDUFuAjYA9bLmRwc2pWu9H9Pq2Z3F
ME4oArlBEyoAzRvtrDyd/wnVbEGAnFIpiAyW7yEfDQd3ObUG1TvI2q0csG9a
qLVKhqQy7yGoW2rSPGsiGeeiV+yp7KJfzIeoS8yp0zkfk+9ZuJ+oQ5IBI7YC
wD4HcIFzkmHNaD3/NL0eEfBbwAVfTGw5KbISe/j/MM3ir6X2KakPwU1XXz40
wCLcnwSLx2LeTOc/4j+jwXeVnFjHZYVSdvoCrtZWGx20nI+yXKYlmGA39IRV
r2GNGfcWRDFPnmRK++q2/BHBNBQHabXPf/lx7C6Kn5gb+ybwxry/QQPzQgu2
i12xIT2jcvCrYUD8Y9tKh2f6AU2f68EK8ErJBgW88q0YyF1PpLPT6IkCX1fi
JcyYCXJYhLUFjjF1e9Op8b7Q3FH1zNP087IAy4lS4IHxqa5ArFGtbhFilLo4
4OLzlGIxxOViaNq2UjZsUFqb/ledhmKvIOWBGfnTK4qfVGwBhPZN9O9282og
ef9Y+RGAF4CA8E/hbrJyAoXddf61/4RLUjVb3Kbgf2ukFauKILVcDfC7YmmI
LVzYPe6LtqbQ1oAeIWrPv2rki3kOUOqUiptqxeLwMJQnskIkoKQ2NfP9wBdz
HsxS119mFGAV/NJt9vhcSskJMxuSIwC+Nafb18aajr0UJwrwbcSoHr1Si+xz
txkWRz1tyfpv2oeU6a0VcuQxDVX0OLokdGUELSuqrYfKzOkdg0plw9q0mdby
Aa8GKVV/mQPNZxZt/7pTDSCkrLezQrAGlZ0Z/EFGTg2kEwiuqAlSTPM3KdEc
ifne4CfcsFlJyL6QYxsUnQS+9v06wvofMz1P+lazWUZT59sURVzBX8VQj8g9
Yy4Hbl+CSbxI2/U9tQpnH+FOttZTn//FpKoGbMHFSxSNcf1Yj6J+Yl2vmLtu
MjKj6C/TBTa1/jP3trWExsmw6snPYIdu2oScb0JtqKFA2PtezPOXEIgwTugE
8nlPRmcqEW95v2Wto+KuKlbjoMoATBuOGd3pOY2GAwuvU0Ea2Bq4qjNnnRzw
5f/Z0Ad1GSSFjj9iv7rkkoB84cvKnQweeELO5PjN9tMRLWwumm32EzRU8uVy
c1ZwAPRIBVL8GBx9NE79oLpRFUgpN6Nep8hmqDlR+itYEWNEFP5ZuJv5TEsA
xfbaDhiJyZksne5mXjz/jXLOdqzRgZ1137i9cJ7ZRGMa1geIW7V1VsOL6UfG
dvqpKS3P6dXNd+Biu73HVQCNpY7AoqdOGbeG02paIGuPXNZIoPPLjNfdnKw+
n5CVEx5aWOaQ11XxmO+YUNjCIgL/k+GhaeM8J/gPEgVkFQgqqn5tFwR0Oqg7
WeCFHnzXxj1PsaEeG+BONkPGvUNBJRGTv8TO8NTGmi8FKdMy1bXA4DC3CG1E
LvflyTvUFxGop7H/LZ2W22jqpaQVrGm/WZRQzOk9pF5C71LbH7RDavz/iZDm
6r46cWmb5PbiExTqSDlhyxBjRH2lnXedEfcWZNyS3bPzNFsISgeBiWXimx8w
NSCHzk8pATvGOKvs4brnBi1CnJHvnT5yhfZ7h4MjVgZAPwkbjVlkMb0P77DK
LBJe5DVW8sJ/yYbEeO/SuRnEw7mGmvTqBoCvpkY3wYcZ3WHX+uMzZskuXghO
CNDbmR45FhUBKXVB/51HamAra3HarcR8BG3yvBXyF70hsh29ekhl4uV31CqR
TuNVOUZDYLo+iYIoBQAhRmpqkmbgvyE+9v6iM0rBpyzOGP0OcDzAjH/r8MUS
3Zf1EO6qDj6umiNysczyD+JI/ix0gbalQTQrxeYfXScFKJRfsQ0C8BLc5dA8
CK89Dg5VQU/zqE5NWifXtivRObiYWObIWaUOY/O6hzyw2BIbG9c77Gywd7Id
a9cLnRfU7yA8e5YVe/RVHkH/SlANNcOfDdCq9D+AW1+3WR4ubUcCaYyFwdgb
mfx/3xDOiXhSpjst3m/vU18V4SscfS5F6pmRr86N+GEW7jjC5L8IVxT7xCnV
+Etvp3cqdybH+x3nn01oQmIA+CEWxKAJxg0fFsyK/ZtC7nPyl6K4SS+iXvQd
cCwXdljnGgSfWjeAcIp+R332iJ4wwY83ReVJ4IfRyQsUsb2oOPDMtIM38iCr
ZQwV6qiyJzNbTojBvfiSv0S5M6CNsfFskyDBHfUf7zYtSUS7x4blHnp8FcX7
h03bCEstvxLIK7/gJF7iWHMwkHpenC9yV61eSh2lrIOwL+r81etPR6A9lGzk
HUvABkfiDjY15dCa5UGmB9Ji9jcKyf22EKZUg1oxRQUsZZXsz1uNk7/4lYUw
UQtt9UQS6v9l0RKVcxCl1HBZ9gcj5SOkXcZuJeZRA9sQBy2J9E7gCxgwqUpU
HtdRoxK75ba0S/F32uoPvAcGkWrFMoCoUp8rjHneubd2qXNG3326FTjZKmQJ
+PUrExQV9ulVafgcUxRek20rxm4gNjQI9HLqE2eU2M94enM8Z0rOYa0uYSCz
rcD65h+N3Rkr25OG6zz9hvIwvMgI0GdGx50GiVTqKKaWonAf9ViYAV/jOTK8
77xVg5xrwR/MonfhrNsibnawRCkA5mp3qwFgYjLE7OSPL444gNwJSS+wU5za
u/+pu1osIQqk3JtZCIloIVS7ngJrfY9TIc0haooGMbDmKYPrn4I5EaxDJxlc
AEvYu1gEqwjp7n19SsgtsAmcKXqlLfsFaeEEXsXBDMRqmzyg/4etnyEFBypW
Eh7qy5/7f/d0mo83V55i5a4KACeuDapgy2MZzI1hbEUtgGMQSDO9YIhD7FZe
yGyRjSeKMAjBba0qirZ3qPoppg1rxucE4s0MYOR9FRe42wjW2wGAER8+BWz1
P5xA7+SananWkVdOGLD5t3CzJ+Pnt5SxzjrRf4a/qneoCiAzIYexUjBRAS1O
6L4Mazpg0wr4y1hlQjiHepvzF78ycthEyou9+iz3UfS8Uz/c8hOuRIcKyjK0
lfG13UK7KOoC5sUPaKWVkusIZwcTnqcRLw489Unohc6ukbd7i0+enWR0pYCn
BHBHp21ihAE03lJ6Eg+XOZyggITlpTge2yd37UbKeGRvBFcwQXTKO1TMWlrZ
XaGo2TgPd2lH4SEJ+8g1dyn2nmB9N+eE9VZcevK7nzu2tdiLbIdxBEkfuGY6
nvltil7oaO0mselSTaXLa+08drWSXkSXnS9KqQyM+hZ3qYYU1Gv/ZHIXFbCI
rFQPddAhdh26MyoYJunkJUKEncn4Q6hxFGdrH+wXaUdgCR205zb3UQUzjuXr
ZZ9sMxhdWTTG+Pa2TJFEJzviuFDgVMO+9E4ErUBW59sLy17tJJsKVEB1fvrt
I1rJ7hHnCXNkvRMhVAfD2BytmjpiAiKJfmMG4MhpXDliM3pYr54EcS4G0jTx
Yg3leTR7U06srg5czfUVTrau9vXAKjGMpTu/csTF/aKmAWWHYkcryAD4CNhn
vH/0Kd0EVehbnWWnCadFQ92R+pQjgTo1Zfh6bzvvczEgB9czC8FbHs9EUP+W
WoWuySrZ00y1iYAVu1KvlFKbfQworBLRcuRH+EivyiORERy05vOmG4uX6ipN
szgLPbqZTUUAH75/jH1s968GCu/cIKs/MLw52BOy4nKl7v//OMQzSDZvRYjG
slkECy/tlWh+uIxXT4vn2BksWgKcfQqQF+xYNqkn8cV5mlGkbqs/26prAQ+y
io1EMO7CQIOZKWoy1Q32f3UVs0tw30cCq3wqKNSdNs5MXwiCna3h3YQTHOOj
PyW129G0tAffnCRZXYyvu4Z8Y9rAnnF70qWaY9+39HT/T914KBXqob7q2GHK
UM53oNqFwgA3Sb+lxIk4xeeeDhlYfpR1tIshJPEHvQWFDEXSNoSqPoHE7wGo
Z1HFdrlfQmW3uS9W699VfCmgNTrtNLQWCLoAMMDy1xxK45uax5Xvb8Onwuct
Ed8DGjgTe4mBqNTw4jQqEIT+w4doqyV9ry9CAnfFR4JlwSxtsG35+xFB92cR
SJ/yqaefcUxwZKp1MOO4KIuXRUl6bMHSrwKWKLrN40uLrWHsNIt3OEB0Ljun
eGObliGUKIsmddsrjNSi5HRuX48sArOQkVId9OPuYxg9NZ/bDmpem25RxKyk
aXlKf76/4+HerRZaQA4njxxoWfzSsIxBZFZo4Ogl6tHaaqYQhaTTpFfc8l+6
nBsaHU3Iwt87sPDimF2keMgJiYlSRQaAhCremMbf3vBBcfCtGGYNoxRWvQUW
MF0HQO+D6vl4mf8eWq9iygkCGApAP7Xd5vA4UiH+Z+KoMrGNWL3eUEkLiXe7
0HKVAAFqqXywCejQ5I/otKXRkv5B5PBwvV59UQ/SlTcVMO7N1boHPldh8feY
OE18jYeqdZ+RSR3fA3fmOyc0f1ab/gbqav3e8QTBNHDwUjErrlk3Fnp0aJVI
2TvFdRGyiBYlc8icMuioAGCiI9cxcGdV3ijiSlonbSVy5IeIMY2vK4A7IbKt
MLGG2/mmzi0t/NUtvSukdHF9j9TYl+M0usoDunKVCupHfsTnCs2qVz/imCiA
9oeOs+zKH/4EZZKM1afFkvPIc1wwwBGl6t7hbcmk+xoCpNf7Bwd3hE6WeKug
EQDLgOe31dLVSleAzu9UrDJKS2SHFrffrBhEKMEIOiQbZQz8cexyHzyI+JVt
ugq3nagkFjAx/haApy7Th/akhCOPjDrF4rrU6RmVFsSrbepuCPmNvMhygg7b
jjBgY/62xq9CCE9ovNsiwJoMHhdJvUfTXYepK3Q8gta2zABU2knja/KBRbll
qr/OyyzTi4O1DkLAeKIIaa8Yf2jtzlGMEENSlexRRjO/qFuhiLoLO+wxYS6J
Q1mp/WInNhfXlmskTwhEpX+NBQXzGok5Z2bfaggO089LG+onkrkLcNxRb3bG
29m/0f/P6QKT1crNFlnJoHGwXSfEx4DnFXG6Yht0OeCj+wD3BKmPqT21qpCF
DB9VF1AqxJoJDPCDyJq1fsAevroDr5VmbU90cjPQIqTRup53Aj8esPMjGh6G
U/70YhePwzaX5qas04m5rKH6m9ct7roQV27QI2rC7scnoxcfTSwQg7sKBWFV
kk9J/ow2vEwSpPk2862lmrtUoaC0ZTb6bmq8e9Tm5GoAvfKu0xI1CaD9Uyu5
TWqMbwmzfEp6eZ9yza38vqbE89Pgn+ZMnknF2dKW2NJXcZc64ctX/Epvy0Hx
rjWtj4L7c+3Ju7tdF3ozyEd7MojE87gvrocT9XL0S/og84FG4CDC9JH9TnlT
SvdYL5w81AWzqtzeIsJqlK/MI7dFyTpjWqCw+HBbBcAX+UD06egUZF8IKgty
irrNTCE0P0oqPeTxND7zF8KkjWhQ7dBr86UqSLfX2Gfu9LsOzd3ZrfjgzHci
jQxcjY4kjewEggFz3cVpkj/NvZtZnOlhUbwyjdRm1qdaDfW874iWUrcJ23+T
YD6gy5Sbi3JlGi9lgkM7OlJzyGzTrVssYGalS7bcpiuFpl1iepYtHtYFdys3
AIsIH2no6iFDf4mHD/1p3adE7AhKXgwWEckRwIqId4TLF+NzNdyfLaTavEqC
IJnSjspTlVnL5FtrANcLbwJCifZ7R+3LdlR6J6GfCus80qjfUab7lFbf+uTV
lxqykbus9RnXJcChb85qpATWyR1jtSz3+bra19ZvRMIQKlFGgs6oyyqA5k9n
520vtZ2dGhAI+x10nzJ4ALJXnVSLIS2PPVPML+b3/YK+kkico7hZxyVPb6aY
KQq0dlYJArlKppBnYTzrbIxzklULgHiUdBXfAI2CsjV4idy+QvSayPgGjNnQ
jv6b7BhHkLpYj20cpPQzPPy+QkNSL3bEc8NJPXaavfFp2d5NnGtotCTAtn4a
XJa/54fexPQjgPcrYCf3UdlkwaTcuiGEgBu4dnd0C0p1pFCwrfhx8A3J5cmJ
eUzwSIu7dZBwV63uAcJrctlpmgyRzF3Sp3iduMtcoZGYihHuUqgrOotSYd9F
ZLtdVr2TmgbVuABvbl+Q8ek7i4/eVz+wtHYkNqFBTJk51eR0hTW83R9UPl3R
l8XF4VgmQJPGLabEo7tAMsZ3ROIy/GmdX12NsKIdpsPRLhjIvkcG1Ei3gkdG
rBq03Qu/2ianHUkE0OTUW7Xo+tk72MiTaDpP+qwPRm5hMLc+QJsA1y5i/tw/
hhk/NWKhDiTAt2lby2/GP1bTq8T71haXRCa+r2Wbj4oQ4c5jMBtcPsDenHkl
llXbHzz2/iVbs/TcDr03hvgahoLX4q/7ssaT1Ae33Pb/NBPAmIpAoWnMLGMK
LdQ4O/c3tEaF+19zqh75Du/MIX+GP1I87x9glnP/gZCosNITIBHrIAAPxEnq
+9bLHXiIVgS9W8nEIIRfG3/rqdJ3TVSVdix6btisq0UN+LBlRagoU6WEL1bB
AVYfKWtCHwOf8U6K1eG6MG49ANiPcbC1vpke+WyepLhyr36VUIF/lf/DRyIH
i7V83P0X93okmOdDsAWjMNyI2qZSs1cqdtBWcFtUUJzQKU8yxezXsoaRMLFA
gg0/icYOqDXMgdVS+c7dj6N36DsiM3B1nHDTQuRIr/o/gnNEJm5xGegO423f
cOCzJm2wC+D1/8wUCeJSPHCv/FQDAAmf2BUtkZ2pB6Mve/YmW1paAE6fntcr
oo6iDXyxfNE12vlRclMvJRX0yYFKkfRcZ6T90w975N4pz1hdNALPPgV2SLHf
RyUmU+hmC7Lx5qwdyVP3dg9Ne0FvNU3FNuGv4i/E5kp+tAa4IGzGpby1+cYs
KSqfdlXq2K0uPcfMbk360h95PlqFG40BD+a9E5xPeC4S2d+XgKVGMPcG2/3q
bAo31bXdSI6X62uyCarIDrFVkdXOpkOlPIS9yOhhOUBvTmw28curqe6GtdRU
5owpDzSanDDmclpNY8xiCWi/JthS/qkqViP2UaOeNobHSF3CLs7I8NAd6PM6
ndjUlGOEjqdWyo/g9U9503H09SnjL1KD0FeixKOkOap45aq5Ue9Cduemzv/u
GWPJfk3mCP0sVwLEdgRVpp3OiHBvnr90Zrs+B+2jePD1LGN3IFEj+WgryVs+
DOxslHXDic/JDhFELglfdFVR+3RYBHYCb1gyyJs+kYtnOPLuW4OFLDsR8fr9
yrJs72m3L1UuP808Oj4RQpMKTVNm2C+WJpvrtgQR6c8QeADIehCQ3LTnShO3
R706erVzAsv3O4HGx0wTH0fdMPtUuXFDFULoZw10mpUXp++0osjhHX04HiB8
L2/Oy1JkqB51DckpZCt6G83yfz2sjmfYJdD1fI/ftN4i83pKayaUbDXjrJ4W
tLjs4JiXiBWelCqmvizi9y1j+kOJbCnNpgXhkmAGcnPnG9tJCXChZLx1Yfd0
Oj/MDp9mfGa1RAtxsvc+hW7Xn6aOuBWmTtEjweghNSL2QVz1AtdGZ8Rs85cL
zf7gwsp0sP3fKtiIuKfBxijPTl4TzRSA2bhRwkYYxBNXTsd4YgMJ0kY5GKM7
mg8iOSJOKhq/6aFm+7BU8hImyJPk+0eT3jbdXrrqRIqDMScElUovGWOmr/8O
m3zEGlaHGdezLj4I8VZ2CARfxKWpGfejwahTi9y8EEpcR/kk9VGPRtgPoMY4
rIK2afMxnYRtqKpZi79rerlu9Ww5jjDqdzzOESXpymK5c+LKSx6XR5N+XXRf
ZsQ2SMh2u3mzVlMIj9N3Qtgcqyoibug+PGMnxKLhtogK9ebRoD3LWcO04ha8
cghMoiEsPG00xRqGz9aQwZC4Yk+kAhpla2l7zTti9NxEJn1Qh8ceJTZoiuSe
zty91MT9+AdND7sEyo4npc1yYxXdCmqEC0sHVR0AGohX7POJI4BOcJgm7rJB
DWUb4YMU9MY53bJGPUA3Ytf8ZS7ldJT4mx3Kp99Hww+i6HYv6zMX9qoMJkmo
cbTqCeL1UyJHv+qK6unwTjIWtzptZNwxk4dSwFONB1i+nrw63wlOTp1mJVMy
mEjAy797JhZ0Cp50RgrZ98STb7sVHmLRXhYlSTRA4dz9R0NSC0kyDE3KQFrI
wkVxMxVPYn2hXRIBvOS9O4e81BeWHn54fAZnE7TwRzgRsIutXuOFo9IMn/Gm
89dCfL+GfVfa5xu+ar5Bmz+d0QrtpI/1KE+zInr2mxMJl5z45YZ8dSFAzzpC
cQddr4gIe5CXA7/vt3NitamSBWoBOnfYFT04zhLTgO6NFqn8l3eftG2afPMX
xh1LLxON2ILIWCSvaHNkAB99gPxGyzdjL8gfssJiPxXYO/m/0Wl8lwuvEY/9
xUDsmhGx03Muel35L+W+xOaiMjVpGRP+HXnBxnmNLgCqumE/h9facvmaTm92
MXeXfGK3DaMVNUXQNcy2CYbwHiCI98xRZ1nJyncvyfsgKMhSE66wRX68gcH7
MsN8VUyUbMpltEHqXVmGSYEY1wB/Ua67KOCJblCiIqH18ovaXzrPz1IdTnK/
StvwEvbbeujFF3l03rJe24KSm1kNNkOFr9iQQiDvYBPUkxus1tdDqp2B1fo8
U3Jx1vRvq7UFS08K+rvgLYAqdy3Gq4G9MJdVzyUdqxtrfnIL/hZeL3QRMSu5
C1Q9bIy6VjcTfEySLi5GOgMZkJ7GfFKp8ZYkid5UNw5yCdJ6oWamT01I3ZGk
ojB1r+Y6IvkVdakBDF4a9pV5KFmTtJi/kbdpdJUeNXye4x7nAFWM0aK5pYMh
VptSnrUa5fWMcZEfnXZodREFg6EKoskMIWoraAdRbB8Wcy2ZKsU5oQwIVF6R
nuIC19/18rYw4DnfrYUmzQ4JyWXuBySH9PLtaGDtKsLHPuSIo3zq6j/9KEDd
SZwb+6Ij9RmkA5A2q6DBhy8X60VapU3vI+LKIzUGRMS2YcPfIWkzwo3Cr2pM
/iXksgs11QvWdwhNiIxap4DI8jr56xkiZb60960Cs6yVT5uaX90orJpjReGV
CjuXkMy5YOAQOuo38O3x52+jK7yONuLJbwFeff5dO95VpQm0cZ47OpC7YalO
zNjpE59y7lwmy9W318YBsztQl8qCmBOAcwrPVWNeaIdiohNUiYZwH38lDU9P
1nU4sX/7ChUXTArh3RoML2+/j3TX58nqSdeYZvLt9jV7PGvAb4ZjvhzGR2ou
Z4xEHQWaWZ5v7R/7NrBSFQ/G/guPP9wRASqDN2NcFO+JykTkalHVwtr6nwfS
IaIfi1Ac70/Dh/ch7Mps61jKUVuw4wq53tBsCz7/gU/bjX1/qysDFhShMx2P
5InK2uKJgtkYrNnuPdct8GGNqHQ0OmTvf9XvD3ZNVBNk2T6cSvUEOJHrSSUm
FmsdiwpTRRFZa/n/HRehrfj/mtPKWd7pO+gXuzwlhR71DrbTsrHFqDZJy88h
LMxRKZB2KmnP7FRyIlITzD8hwVR6zRHLUEbpkomb7G+9GwhRYaFozL/U/ZNi
Jnal+YCCrdYkjHS8t4k1LZbe1ApDnlq4vNWWlhZq5Rkcr4YuVTWUT1qt5935
mPejAF+7IJMWgDPUV5D7c88DdErljJ/ANYnZwVuhTtL6Du4tW/rfWug7IPMp
R3tHCGYbVDeyb+yX5HX4Ew5HcTiolbSN4ShEaeYvrYh7yJsk3eGvQmaHdOrF
hVIEhTqHHOtHQ555zOSnzaX1zqCZNXM6UgUgy3GxTbj8koy4wTnn+g34lY9Z
ZG/bJvFFLCEjGRdYY8EGeqpLJzlynXnBaujVri8gotwZOOJZqCcUHPrW92ZM
9HwuCwYSQrfWj7pTB7p/+IPVjSdtcQdNzQQQs+4IFGaPCqi4JAuE4JC8zKYA
MhXPyV/thPHEwGcudh48iPjAAVP7jM8QbJyAweKw1hFYhCOY3T0XI9SVE6f1
szhQD+ZLZc07WOqKohxPJRfpNQCiDrK03Lg53ZhAzA39yDx3XfhoB/uE1XQ2
7FM0cWh4xd+BUBgK3qHzjswTwJM4RZiCzRbxbJ4JAUxEFwh3Wi//13OrbAdP
kwo3g9OuJKA0y4gVX3n24oRAszs7VIWQw9oLK2AUmaIP2r6cMh0v18HTu/eo
2qmqpQj39gn/us1zmbndIOvTXouvhTAVc3bMi869e42tNhesBiHQrm+uv7MU
mSz8tjD2jvvqYnWTU9S/tZn6JXUf+mXGiKDuFWGUVLLmDIR9QRhZq/c1N9wC
/bqjURzRifeznVSln+yCU0o7IzsTXlkx8wg5RUgFMepF/CMOLYxcBqgU254l
qFcZLufdT1R/20eezAmZSP2B5jPBQcuvgSb+117VYbyTGn90my1vM7VBwJNq
ODgef/9cmwXx1L+3WBdcZxLSeLurRxtjtGqxnB1hOkE7l9hplO89HH//V2mT
WELPX6KVsP9bfiG1mBboYBRKffJb3ODPZqumalygIm7gJNyuVzxSGWmRUktx
8esLLq4RaIU3Jd9E6TiGvuBj94P05hJcvpPRnqMRR+BE71kY4tiAOYc4XEla
oqSrCGhHhiV7loCelMPBKcVrqL6qSLCRz7TZ7YjqNR73VyUbGhVOEogTqBpP
JNUHFFnPWvq4cvldgFHsxgdlU4Yo8SGCblwjII6fliGaXuW7qZShetY6NZ6M
+Lna72C2zehVOVTfppIwbVtnC8q7yQSSnyp0cT0prk2/jmWURAadcgLb8XXb
p/S4RtqzdpAL/k97HElyzI48xz6KqD+EDJNBEpiayfrGson3dXmI2YQQ+/EP
cfgbyMWdvQWGLIufA1TtsImfgm/zmjmG+GQS7jd/kv8FPJ6/nLKGJYhpRA+W
o9Krml8aqn/kP6nRfYMTTQfplJHku4Bed7/D0WP765xPhh8nuf9P/RdwyVlF
ps14rIaVfqyrzUn8oOfSISUpuWH4CzLidU/GBGxm12Dvjtu85zB7LskPgIlN
ka9tCuJORWlXDq3ja+n5cyNS9RYAXtzUS+YxCxqL/wOIAGNOjX/6vqrJBOz/
CIyVtt45TdEtJEwRfBin5qPvSoPtoxdJ4LL/RFa4bzTpd7NrWd6T0a+h7nz4
pclUCmgJti4BZJ7RhtiKTaq6OtJoEWyJ26K7iJAaPeh2ZdsykMbmiUN6hS6a
g1XJhsigZBl3di99PFBogkbjwI1YoptUGWfdqRdhGaXb62cq7h+yknkvVEVA
EHSl7j71piHbICrabzuinW6an6/fpFzL5ldfPSxrVHBPEsuCPf0sl50zuOXA
Xzz1YMo33dsKHPpmyGcLV0TmkVJmiB40uGQ2PGf0Oj44rOWVQFkjSHKjm/L/
frusC6XKV37JNGqnALS1oAapv93r442iRGfEjqgF1sy+3zkN4BOobll5lnjs
7gK4XYnkCXnyYC+dM/GGPIgresPCiePI6WmLuN+OHaRZzZy4S5OfGQ8X3OqQ
xZ7yqHIW+cgu3lXqM929QDTO5mWmaVFYRbQkAu9/Hg4H4Tvy//xe+grMbNK0
DKJrDjPg45lLWcwZPOIVJhWYtg7VoZjqb+Hbzk26c08Ler/MsTfFvwtlPrrm
wgc04Wg0I94D0ezcgO58PZ/tPgDeB4wlpEZpQozP2s1WJootkBVq4/InqDFj
+tTs3xRbbgUabtHHd3egB0n+m0SVtJqliJPlXzGjZLCfW4EzM0FJ3yoPG2+k
SzLjEnceyxaUC5i71XP8id0rX3bzakNglZegMJKfEc2Wm+eEhAx0y2pdK6Y0
nQl2YV2u+0C+ZiIZOmTanF8VZuVjf0KdPVmgqsDcTxVVEr3H1EfWM4fJDal7
oI0G1hQPnnMfMsEU3Vnz3DzC7G21NyzlmbtbgCq1d+B/RUTsLmQOfB7lmNeQ
VRec/Z2rcSXsFU0IHwM+RPN60zcvPSt1lWaKSGYnq2CfzjbJwZScMOK5rk6M
iLlgXxTWmwBxWzn9jBDTwDmAKIj1Zq/UaNeg2Nam1WTFyhAgcXohmWTQSV7b
Mstvcin61PMEGpqlrmZq96EDbFaUQD8FmhC/w+c/PD7QRf3+ExgZJMElRLwo
owG3X55MA9IOEFa/9C0JaaE6DUg51fM2dXTXbAE3oamwk5ndeIsVI5A5pLVe
Lo6WokcFkPArJY6O4YOJiIoY9pSVuIznjSk2zv0ZJvi3qt/LQJ1t6KluIqIB
lr9UTF467IaPVwMkG4qNPgVIdHXeo35rIUQOv/F3T5Po1ooyAbEuq8rloch1
GsjFoD5YO8io4BwFowxNKbpcAcLTshGjpvZ0V+hGO+FTl4+490kfG2Lt6Met
NZ+MIKTUp69oHG3DNd3BDQNA8o9UQ6KdhtLW5U+vmbUpPrJYSHWtM9a7l49A
EwnEA0LVOzwgQJorkKRpci3LlVGm12+aRGXNwJ40TXheXXFzt+rqP+if6gz9
H2EJ8b8uorzC01uVsLanq9sHf23ST5ofsg5vI6HmBkNPZ1LxhjQ7igcl0GOv
o5MPYS4S8htvkKcrAHCn9vHDC+uZaSl8k1IYGYQyu1Ke8ERTIJmCQbB+z39b
eTBrVnL04TAfCWIjF89gNRe9pV6LAKFdXpe6ssUmVJ3yohy+w1/Ou3JwBhvt
e5A5pCZM38Sh/NaBCogBJ67933ITbYqTRjMyiXOYMaJZz3Z9lhDYBmBgBisr
G9cAKvnANnNy4ZLmd28d03SpKBWRQYAUrP4nVLQ49QdURcj/8LRt9BzTFDvN
+NWsPQsORqbzHz2sUUoNWS7hRV2sfe/8xYzidFXzOuRrc1TgD42QCqKN0tnB
EkvqMhbv+o30KBzW26q4CmUcn2YBreCndkSrVN/oXAVXl66AFSaFTR+xwVqR
WyRoyFhIsKbPcqOduJuvcoFZpAR9mVPkirBZq5j8ny15XstwCVIReQsffNyk
KAXTApy9izTCQpab6VI21NPc0GwhnAcCOfGeWZ0Y4e7RI4ZzqXm7i1JXwwAU
W9lkc7X+ZfusT6YlIUpTh6kbkanZvLMob9jAjKRkd3d4YDCNWJi2hYP+4tL8
nujG7mT86SDKZ7lCXa+Z6VAalimn7W3pRvxllnjlGoYcD1qCnuUmLq7PazQW
8fhM6naoa8KGNZyP4GgMiUrxLgEQW0PSCp+hbtsFO4VkI1RBbEUwUdLtD9n1
VNAehvgf/N8XCCGebFBknG797oqXcac1YeCcFGxTWrvdJkM2TsOPqT/PG8h0
4F9CHJu1qvKTpxty3bty6n0yPqn6fiknpmbyjJZXQc3/KjxIdTtOC60VE+Gv
Oq8QbxDPzr8eSa7fU5JbMINNArMxoznXCfGaxG/vSoVZvRPaW60VOiuJx0iQ
pArgNjXqHwT24ZR+Ss3rKeq2p3iDnXvONRFz5L3T22ZQ+FenYYg+MJjRx+eP
Sbztv7mamqaSRDTmg12qffG4NJm+aUOB+5/JPkyfQLDImwaReHDvekhn9MeZ
0yYN2CMDgITwlbXuvLj2pZbOIGdNotah3IpTyB+eTs3TqFA+wziPvy3Z0EfT
B6tggXECl5yDAfA+P5xfpwhBB3U2li5HLRi2yNZ5gled+1f+xbkpKWW3vqy3
ttNpHLe46wkZOReLrKA0lJcJ3s3yoj3oXwBUWq5Ra7xnpBbc0UeAqoueByNO
kHEcW180tpTqaFG264y/in/B6o5N3i+Qg8TEI4oLTDts1AGS1oiEMj6Gpb29
a/MAd9P6u8Fs0ZZzhKvK+Zii7/RoH3FSy1tcJSf7q1EgOpKeIyZw8p80rYPL
SvR6XFZgSDYYV9uHlFIbzxf+Oo9xCg66QPGo/77gYTcPgXOTp5kGK5unwaL5
q9rhPwFMu4rH11ZG6ye8ux+wlj9Fjw5ouD20+ei3d2JLzseQct73HL/gbBtZ
tbXnzIT7aXTIBPuvMzN9VHB3pAJXczVEbC5jJPOy11qvIJuMzol8kN+Np95V
MMbJIAZlZAPZ8HB6IXfwu5gUM4UFwUuwkBlbli6HqixYj+1dGiwr/vDas8rf
RrsvHo0DjfBok9jBLLn0d3j5NumriNNgSD/suLU3c8k5VpLkg+5Pgl7PsaUU
xoqRlgKZcNYtYcRkQBIzSmB4/PBCmWlsqt4GZv1z+40he+aSFPmxoL1YVVeA
SLJcmjwrf2erOg4V4Q+oL7lsQhtEn/By5HBs3gmhIZeVWV51NLxy5l7NRVQS
eFRi07aBgabCViCIjFzJDWulTAHdUUMrq4DMkTgp+FYB7Ybr5ysNZSIdXpmZ
ygC+2abnZTwMlC7uO+keV8GOTToY0WvOXnEN/laM+MTku7Ih+R7ZqLoyYjMs
a4ILNFDVlcqlWJyyxRb736Ezgv55wwX3r9fCKDkNKT5h0UwZ+srjn4AIazvd
Y4MRDIQwcvB+y8R1E4Udo9lsxbCCjNLr2m0tKAwYkyzxEjv2JYX2lsJc3c3e
MYbO2T057mftUdQcGIO/YYBkKn4ekWBZ4KJt8JNOUUaT6QgAgXY9i4mgJYlM
TynmyKMEV1znkuUqemYKU/+e2e7z3gNY1TZ4UhaYjOxGOw75I/cTuI32FBt8
rucUyR3bNlJCOVe9hwcvYJUAIFU+20KoYfiD4xtTjz7QrKkcZBqDlV9As00S
v1dM9aRWmKN0BP/GEuqBLvORVPQcrQrtZD5t1CvjqOlcWl5Tj5/FkhJbwmOP
OzMSRZuvlR9XoLRIazO1ZFed2KEyqWI9CI7ILrkjVV7OIS0gL/l9v4ivZYJj
xtUD6ykofhelfG1mPhqVGe/c1I5yM4j2Dlr3Ex0UzCD1rD/TLnOu4spP8Hf/
05+TmmobHjp6WYAdEZd7u0IpJWamRIPpIgYxS1s+gvg27nSeOBVDcU6LLY0P
igNTvOBzCLiVSdFL3Z2XEukPUq/w9SeD/4Ei2GYREj+h8YAIDf9OtjKfHAZz
aySloMS2tMQM9rj7lLH9dlU86I+leCG59IHgsSpW4kXbRz3OYbA1v02bAvMy
KMP65R4+0F+Af63Pdi9e+P6Jf4yw7NpY37HyZfa8PscVp9SbVzsEXcwv9AWP
wRot8Qi8R+vf21HQ8158OUpfRq/rskTQMPPaUIGwh0HpkamN0IK3bNAGmpvJ
xukR6NXoNYuXmFQYObYfIcQFL8mPGvj00kT7tjzkvSqGA4V93t5+WUun15Co
qLOZYE2RgXhfGluPJZn33CHKEWbTcihOrp2peOrXwa0CtDDzAtoU63hz23NN
lsEnmgt4d0Uav35lNPljRNz/kBJPChN0yxKe+dKqwR89f546RMvhTrC/Bqf0
ERFaALQvpkuhK82FkjoBsIyqDbNFkEi/4/RiRVD9kmRaEeK9fDwNsPJgRhXm
qq2ROkHlGatLNOcNKzCRVTaiJl6h/hqxcatUNkJdwnyD8aJE1XO3/gyeqssY
IN4B10KZml4oRsP8oof+3Fs2zMPqKwX/Upeez1ReEJsM/PzqQYKq+IGpw+uF
EtBfeNsA8cEF811RvWXqgwIeiXYW7csaArwCKCd+tR6x+Eg4ciZ5bMf8mVuo
cGVmb9Vwc90r7XTU3QGV9gPplZW7klBCjJczw7XZqI0aB2ff/c8o6qbzMQ4T
OG62I7GprS1IJkaJA+R6AxPKJpYqxXJh5pXmhk4kRXz+43uMFkt1OdLOMuVa
lhQ3/ZckujTxLI/DY6EjK/kTJOUJ1unXOnOWBU0H9ZmUP4G0e4T5PXZ0gscr
8EmIuowrWhzavdFe+a9WYIeIVo4QhHUp6LLaG1GYhce1WjZ3d26k+eoBQrb+
AEOJIrnBLTmj3NQPH5lVdMtC4vAXf5KEetgkpubJq1RcvAcyQTGfvaxx92Ci
WA28rtenB+NhYFYoO+DmThBEMgJJyIraDFeWvHSPNMZa5tW0aNPvAdP41eDT
51dlVocpzIv3HG0EzojIr9W748oY3F/rS1j3mcpNHcyM1B0FW9fxNsZhshqv
0cZo8ydKIJtEkeLVa1uqj4MmOgZIc098bW+1EAfWJiytuW6TaaBKR3cqJphI
1m0KShK8jPM5RE5xYo/cT5qwRZZoc3oqkFPuYVJOgVv8c5J+2LDoAkq1FiCQ
CDYxlsLdWr2aOKkI4OVT16gbVGKGEnA40nq3h6yvZj7xqYuSXHn5yyv7iKqE
fh1iKsXDBlyTup0b7hY0lWSFe2YmWumMk1jfb9YzCSM+Ek2bgIHRxlQKr7+z
9q5cHcsMR/MKnKup1s6fFreyEX8CviuKZxpj6ClFi1ojOAOEO6eGrfBYMqMF
O8cs6b8oEzN5pHh42UCbXzFKaW0mJtC9biAaFpq251gXgThxifB1SJ8M+p4c
LgKmoONJv9L4lQxQrataU/ySYhsnsWJlqFT29mG0g5zAyZYVpY6kHF3dEzK3
+rXNqC9LYVxIZBkdEu6eDnsed0RyrXT2jNnzXKNSHYbT+++bZQBowZOt6w7q
eOsT1FhURuEaGfPZIMMkwISABOMTApRZHZyvABhGAIkCeLG6FEra37eVh6rx
uPGFml/5pxcqkclHnL94aFAOrghIfMS/Qe7e4PNd+lnfcWw+SCfYMWnMCdys
wzq8cO2m82UpVTtti+jlP2MCPGkPTZdTW1/hGx7geI8c5rJtAuMZhuQUU2ML
eHOaRCOaOQO+XYgt7nHMToz6YCNtv54QtaFwcJSDYGWpcZSTAl3o7F9y0I5q
AMbhGoA6LG2+YOqEYFO36UCcgAYz5IxlGFBgJGBYMmV5+9SomKs3W+nJxRhG
8BPtUVR/HRHJ0nWftJOEFgr2KfJveHwyVBBPHQYofE53LJUOm2w4AP2RJH3I
IHl4XT2hRz4/W6RtgOOAWgDaIbbb31NclvllhGf7mJ+0brw8hW09g4jtDt3a
anQoozl/J+L6qAOnDYVafaVWe9+O0dr/ltRnMTiSfa7ovdztFh8j13ogsFLc
fEYGKxj89IiODW3ErFk5z4MQdGXlWDNgAFOR0cgM0jmoDZW+zhvwiZJ/CuGJ
09NVRb9IPnAZZTe7FBLdtgPB1mVsSJy2sqq1s+YggeJeUn21KVtC1OZ3WM9R
ZVttzdTWaMRYyqGHR9QygBZIPWQ4MfPzW5RilVwn3Z/ebRRl/GWMTg5BXCSU
88LmsYFCxWG4f2tpi3Gv+CBJAzQ7ENcat9wp7ye4QjsiSUalkEFmR5VVDxde
bfwD7kjtyWiImIhyk8j8BJwMTckQRZ0TePW0BpNa5BOsqXVgn1mxhglRm3a2
yXFrAk79YGDNJN9ZdniSz7009vaf8lXkWfFJwIPxeK95U8yb91BWnSaNSZ9o
b1s4//u8zIACJRMd0lBNTBUubn+zsDA4inYfELG0XwH4iG5BD4MGnhEyhULr
yGvREhefF3P2fEYMNuhxGpbavKV13pBP5b9L5W64Xz//cFUsfJWNG9JCHMIY
pnHyGMJoq0oLTB2XNQWzteyvIDMrK+QzHQ+12dYPaN6W3PsFFPxYBjB+nysO
eUvqUqVBkpChFoPVHjtqrCeVSQ3iZ6BZ7tLw2FX/QfJX0y8ePRcQu7kMrx1d
cXEBI/qXxWD7yg1UvnK12LSqiCVPK6bR0lGyboymuY1/GmOGKjGoJQXEF6aI
6RBWyWJ13C6VDDFDJ7WfP+FP/Tqtzm3B4zHuD2LNzp+Lko/W7xiReRkMuyjg
tlwaTfkf2+KgIv6ZdrO21XmC4S2xc/+j6+cyV/CvODT+H5wXUMBfXGFhs07r
Wnux2qZArxtWgnki72dPjdjSbUVhUcGOWUBauGlwNiOFBFqJg6OF72o+tTJ2
dkQM3xzPI/Bjp/gZ0lzPM6i1EDERRMz9TF9xAbZpKnP5Tf1aQhiGlrBPGAkI
H10KsmNYky/q8j48fDDQzPxbSGyRugFGChmqInXY6oc3sWB53DFj95yJhqRP
tO46UY/7H0m9hx/EuLpgTGqcp+he5/bOv/9wqnfGyDNxvqEDiBqIi5oJGvd3
99wEU64ecHxKnZIyH70xTa7Va6343EWWZICHmV49TeuFrD8JT73VrSI6GOM9
ohQJgr8M1tAswgrfldEF04AZy3dxHYyhQgXDNhxvnhM0R3i9mdPSkVV2SPNc
3llALDHdgKgYpaSMnAy1rsYQ511Mx9qkZ2eXino9axgHS114PtHHQDuQlqn0
qN6/KCO+i1Ytr2L49pOxc+EzUkp4ao6drdlaiR4ayK5WY5Gf8nvCX3xznwaV
lq4LE8wMXcY0nvy5QMLtDU20P6pqY1yDGwCXLjiR+JyEkwLdBXxhKlgrw7Wy
Ci8KBiqkKmhmt4dAL5690qpne6CF+zascS9kWUuRxsU+IZ30AW8iEGvYEWiT
q2qcOujornbRCADJd8d2cUfMzOSGcunB/7ZueBNbT2EnHD8Nlnur9HC04qtq
N6VPOw/23B8IvmtLk1RoUrKl6PMurNBRzf8NOC02nNNgikNHDqK7h25+JgZG
b7OJnv9DNVrc6uOOwfWtuzVx6udpfvrrtLXi3efmEnrhflZDwzFoXMfTZYRf
SsTRuKt0Q8PBTojz1yAwfVIkvZHJIh4tsJ/C0XWoE+Qhjn4ED5nbLp8PTqBG
FuZve6a19UhweGep/tZX/P0U59dakbFuh5dhi2YRN9PT9k/r6/k+6b+piygH
O30yL/neDdKdeHnpUyVmJEk0o4tA3Mvr19wvAdYORED+2MomDFg91N1WtEvv
hkRgky1X4vLawOJw7brEf180Bt73Ii10RoiVyhGNhjbAk9ZT9M+kS2oIj8EN
lU6uoknTPvhYqo4rA3u3ytEtLUUmm9wZWVeAtQqOIHpV67nO6WvrnRfqcfml
40rIYcV8gbc1g0s64EDX8S0K3gjGhh2B+oQUOE+lUBmF8Gl41reXDC8Frk+e
SEqeIHOFNGyawnZyETTHH5g3sDOhjbYXu/xLV2Lg8grvrvKcE6gVNCkTqx5y
eeourlwo6v2dEuKsFyV5b5337k5o1GgpjmyXy+xuLK80eT1ER+1qFA9CKNFS
Ny+cJJDSq66+KGjMd6GEtpJd64S6xIi1ggGRCL4WPQrYjpygWSymx5Jtn64D
niQ3JnRK24W4aHSk3TCdJVVz08caLjthiqo4cq5IO9FHLHFr68DaKdFOfirI
6jo0xaCwkoiqA90EeLyMMOpCi+o8CxPJLG32oM7VLHMyrQlRJvOFcSxeyOj8
v5dLlJPB+UgZMX7Rz7E0LPKNLtpanyTAee3gxSB3hYZcrZLpE1kZTvhBtafI
5eE911F5dHddB/6Og9tsMTRpyxozMh6ZwoRDVJws+LXsbAP3SrvU8tPega19
wUtiBJwpWhryTiujQITZWghOpR2NZXuZanc3oPJ7rcRUVKFrj5PakcVz4W8X
aDrruajxqal74fWlo0XVs7Ubg5X/eRpNrb+lzOzgBlTYBPwrIWA38gAiBq6o
gzub6sqyzLvVogBtk+u15oE9mSXS/7J15WAS8HDIKrlLRmg19Lspko6PuB2d
JNuhKFyhnL6G1zmhyokUj2LxFq4qc90Ds49y3zPIsBlWtPUqjAAJeo/5rxsf
rKOPI3Lb5taBd9pE4UK8eJ9aUTgsVHSWm0SU29Ynb7IjOxa2iJZNuDlcMwyo
LB6Z+tPy94dJF7fisA1Q/GLk/EccOd/j52xYuqpsRZE7y6Lg47gIPF7PyyXE
T9Jue8jz5IHXnkCY9m5z67xDbRIlZKw7wSj4TyNjw164epmlU27czjjM5SEp
W+/DUPssgX5ROBN9Ifh06dbYD5LJ3ZFNHjjI8aZHXQvsdv8vuQ5GHdbFjAxl
pl2dsFaVSW/2lxayt6J2LBEfKzRme8T3gRc4dx7ZnYMyiD6G8NnxPVbw8zsS
Q3X67s6Xh+I3uynMBJGFlFgxePxOY+ejvZQMaIfpC/QMtXszCLqX3ku3Jkg5
b9u/IJNl72qwdPGBlEgyvKpKuoxoyQwCG7WMsIG3D8t32UMhDuiAfgRRKM94
VT35lhNXLgUxYdvTtEo5syfFXA8uRCVALOAu7Y91qcOLzGIusq10mgr3DRK2
rHCAmkGqfBuNrWycLWeeFgU4BvYUWKeVtyuatg4Nopns0cknFhJ3635MxliI
9VyvdrqFKYS16Kc+mtXhS2r3co0h3TgeqWnHLCttcWwIiJFKztLK6xZ7OXA5
f6+znNIDV8LdRNyXK6OafJtiln1JG50nAMWk65STFMSlayqyB0iD3YpDh0l/
1n+5P+QgpNlAluwjSRC+yqUSwPUX3C1m+7V4mLaxMib9Sf5OYttTeMNX1NGe
DjZ6WCJU9IC+xVfaqCsVi8rVKcYXxLc6hQC5SoXUDkECLrKxXpsPytX837Yk
JhZQN4Lqyy0Bp/4RgWmUgI8HfVaCnuvI2EI7VzsA5iobhMS+5WF/lUPmLqWT
lEfc7+OxHR5fnIDuwK+HIQVHck/y7miJ+4I8BFxXch5uW7BwkYVw84MNQEY+
rCpvFwq520c9YAm/f9S/YRFenM2ecINiyC6sKunH/NxEIx8/lgf9/+gqUpTA
mtS74tX8Ol3Ba+i3YJSObRCzWQwVX+Gc9jqq6VYJLmNW18q/+sdWNHn6LoNW
ofP6GvN1mXjkozTttgW7fbGq2LNXPVL4R9opqJo3ru7JLBHf/kznJkn+0080
ZG+o5LrzpSCL6SvpPKbE74J4K02nQ3S33enn6uHLPSY15RuKhXstMjJCPWXB
PZlEAhivAv4yl3Afw0GqnHpMT1D/Ypan/wYB6Y7aGntIYsVmpcNYqpGEOz6U
yF32Mdo6iA5TIW/JBqkSRBSz8XZSJbYKGIRN3/Mtlwfx9yuK8gZZdaH+Xx/F
VsohqCggQwM3h+wmF90x+aVQr6lK6yYH9O0mTfzXQZiWf7xDclg6c8cGMPMK
Sl0vKc5dL2jrlfeINyibtSWgoKLSfELPTlcbiUHQsYSwvodoUYz0+zCCyk1z
j4FrpQ9Xu+WCq4NIVr7Se6kjF2cY7XHMM/Dl1PbFK0JgwnbX+dh57daTGFn0
IvFidKi00dOd7b0AaOkJespfMdNbSvOrCwtcHAVMTV9GZK/R28wNRu5c3CG+
ZSR3cuKf9fSIRtDMZAWRAlALovnvC4TrhZZAJG2Dl5GUUmWSEwkMSl3KtiRn
5v8a5x6P1BguOH9KiXpnn+d6RSSHJpnRb/nxLiWS/Lmp1sLjCiW26jrnNCbb
141z6K/ZPP3MxsK9y2xV/US8rxd84a8USmJHAA6t/WtDgyLjChHIzEQvm5m7
PHCfEhEGXq+hL14us5AJudlYZCDgehMTFZWgWI8P13G5+IycLBxHo17z4zXR
+AQD2I039csdSbhUnEEgA9HYEqh/Cudk26W8pOol+PeIXoRIV34ugy5yNGGc
1ZMnwvJZEBzyRy3Qok774q0EjdLBnZ9KRm4GXTV8JLYdkb9w6rj4fxSGVbPu
kMW5CV9e/L+reu56VBzH+xPFLoU4nWij7QmTMROBeZGFHJBdsLO5V4BPDa7K
TvYIskJu+I2UVts6NXpSQakBK0uZHaemzFfKt3L87TcJlXCa20PdLWiE2xlD
jpwr0uy4HrFObFU8MOeej5vl//nb+ShFKl0tM7Q6XLDPLB1nWj2uzL9KoFNq
w/xtB7x6CeEiJHcXxIsVQUDlZCDjEPQ+qT5gzAO0TjdnaqvOpvJafCnI1ljc
QHGhF4zsKImOx6p5A/xm609/Nmrj4Bfwi8+in9675Ay/HsSemgCC88tDryU2
tR4iyy8VrsxKSnTdJtGVhwswzAgqj1hhm13byq8rhbjbTGxaW+nmDa9OMJ9R
qJudApQZivu0Wvv5SJOn9hz0q7Q25OVvZk6b64ifpmRwEp+93T8ZYyyvTLVF
eteHu5FyN+7Io0amYS1CmdFXBOCoRqtJYGRjXQJf6/YcX+TbvaVDw96zVOht
rGnWnQxKTcrKLRdB2a6eEdcx7dVXWozBeJJUDwikBYoDSexS+s/Id0yuT3/u
Pd85ruwcbErAX99WMs4azhL0FELGOEJqfz41BpCqEkQnwTj5ADgxtHYtrqvQ
v1aasNP3Oni8lCRZrRbQMdnerRMKm0bq9KU4Y6PeapD5SY/MuWRcxe0BHW5o
h03ozvdEejTEZ2qhH+bUxXrylpSaoxG/mhfTWUBrRzPfo4qgQAY8EEYYt6mf
/yIu6+r1fLWXNK0kqxb4wFshf2GErgxDm8/O8CWCUw1SsSzXjNSC9WgYhIEp
1lmlSgheoXuXVhnho+Vjm23OZJ1aSE/0gv8Unjb6oIy5XEuo7J7TmDRkIJQk
LQpwje7yh0Gvh4FsYw1aRUdehRLd3JkKEBMmnRnmI3KsF0RbDFL/VcXI3xNd
HOt4Z/C+jqbErJCpZgztTKT8qEaH+w9YU1dcYNxtBEpjC1FYViRtqjzEnwD4
ZMcEgOrcDRw6sJIdFtCgPDp9wQA3a+b3cw9WXzLRCoRkFwm/qUKdHBo3cmiA
RswC61F42x2TAo/+mgwnYm8SXfdbZMthbzMhPTXCfVMhlTdNOh62YAZl7Txu
+cftNd0In2WGoky6IcqDtWOgESLpFMbblt0ZGyz5AvTNuECBqJjgee5h972U
Z7qZP0dW0jHjIM1Q/ZbXgVUh5jbMZuSU7tl/xvgmyDHM08MaRkjCrfyNQGCM
7HkBYkOkKt5FVmWSInrHQBvsSOuIcwXjk3ErSynlk2Q+uF6XFFFIYG2IqgC0
Z9Ego12lTpzV7ds4UTR4yjGEKWQ9DEDO9yii4jcCeYFb18oJcNekqvYqerYn
FFUwwqklvnIeUzk0jiCSxfayTPl1nQyFaxGklrM0gUXHZVIuxccFnFutgNvb
kJ52/+cy6SJiNePagO/1xCAkE6bb5uh65LXoZbnm+/tz8H6WGMVmv7mO5d/c
Y7MmAxe4aJZ90vQWBL1lfL+wnbCvbeXn8wLtjEg7bJmrQqwl2NWNWW8LbRZQ
D1bBfBr2WisNJk240Zw5intdX/MBliLDDEGzXe0TOSEejInJOJbBPY6XO1KA
AK2ZBWTd1OgHPl7+kMXfTEs8lj6fxZIRnM4atwftz5NI77Gk66L6MuYFLKWM
dzgtRkjbkDqhE3kRsMPDV8sjnkIaFccF2iwMybI4A2+0BMRky2pPlxfmogQo
zoRJo+JX7Y4h1ctjEMioWcRIxAkJHAf4GVL3iWBAD035VdYYARgd5M7siry3
eN2Iuy3WFWtpRisqQ0056TrJQLOBlSk+Tc3udo1DL70iBq3x1WwET/omN3q/
MQnbX/ZjfdV7rpnYOi/66gqr+8xzoCT20+l+Q+m5wAwxEc7rYo/0MCDyGu3p
Lu6ggJrh7th7RM8Se5DMdjpVi9I11/6fpO+zmn80zNuLqAbSCgyvgi0rmVCQ
lb9pbSwFXGI0xIy38hBzWlCGGnCNrOn8OGgrcQzNgTnXaO0W29aI4DeCDZTz
DgiTrWZ8QWLw3v90dZq1YHFZAYzQhWqF2T1ims7ikcu6bTBHZiHdwwNFlwlI
JN+2T0/LyAtnGSEwB+bvtL+XLXPPTyIrcAn6Uc81xOc1zmn/eoHhjLQqs4RM
obUvfqX0z77gBjos+o/PgD/JIc4riy0lqb0MOT6YFArhDHPe6EjMqUZL5gmc
kVv92m53HFOqKUj4QeqdPk5ASyyD8HwZx0dEf6bhAxudtOvqyNTFQzLdS/WR
tMp+EyPAfmXzDFrvSTxoLZLOL3pHuPlN2AprK0aaNxNwK3oH2gnPYVnemhg+
Q7CWIzuBSOovvMv+zMNKf5ZdEqOMQVbneMj9fWVKVpSTDnsR8+7OG02qdFi9
gePzVdhgSoMhFBEzIvkiMTIbgh4kl2A4dXV0LhujMp+EIZM4/LNCbk7k2MdT
IgisN1T0hzqrZpioFXZXO8cqWZ0jBs7lUwW17VsAMR6m3nMyUa9x9XiH10rm
m+63AslLNxWrqyGIqecfeNX4VIT6JGIRPADC+kj1eL6V6ts4cC7hwAiNDJ0d
gZHqW0ADcPgde6A+h58O0Y46CA8/svoWFYOlR3MhwDlUfEdNBpyAv7NJ6msd
XcXhfxmo3gNQ00Bd7FMobc9frTKbKKS2JtSf+TVyBIbzrsnosZTxo5LHgDhw
dMaitY63BHllACIbHwsLr9mc/hZhLlWNKfoUL78COo7nJkBNEXkL11cpGLEU
fSjGrMjhyQxwRzbZHdvPO7rK/rkWo10ru/vB43VjMnGszZe9jp1/8oLDe4kz
8cFwMthWSOrOVC1cBmCvn0FaY0kg64mdYhFvAfp44DqjiwiUb07ygT83fzQY
hfzn8DZWSKq0F6rgxkSmPFwf9ST+S3+OxX+HymvJAkNcSIHGP4ElIeEeSERR
RWKyytZpLDcqr6veIMAgLouzHZeFsTsqdnlJPsjVFz8o3ylZWYttiHAgfUiM
b1Y8XPVQ1mAAUkDyEeAUUGXFHm64+wYhkqTqLzpkU/okXRxqulKCHCOnaNWl
zUYpTPIZbV5UykkA8M6x0DHCq98pEC6eEV+EX8HKkcopUrnch5ljtwDVYYFz
UvqRAx0MkiV668y+fiSJBH/0MSpjJemHGuiGcj5Vff6xh+kbmue+LQbxtBGp
8+ZIZ3FFHFzsxEC9w8dFMdmNntbfgYrbu0D6olAvmE4Z1rovOkahmbqouHkT
uvY51YYp+B6Buc+mpM4eaAM6kmFlHZy6VUTIThruFrxpawX1Bzqx+/CO9+d9
WN13q9tr+ztW66DfGEKfmiP8MRQ3ZON/qmwqKRLqxX6pxH+AXJDWPQAtGQyk
LvjmgrsmhcMEahjXSSDmU8bhmlBcfjLJnS9KjSRQcTd8tz/rqFd5RB73wrAZ
7mmi79xI/wq+0MO2RV8HjkGljN7/Gfj5BsVDHA8eAIrpYF3sSUXBMO3re3qg
/D/2Qm6qJf8SU0W9CDACIEezS1GepMMa5wf1NWxXmqCyTBnsF89xogvEkl4U
vAVLymt7FmoaHkR1a66mvDvRLyDYdEXcS909Nz6j2Qr6kxaZXMFAoTE7/2wC
0x8Sp9ScL3scNuEs5cMNl2wi3nkBr7lWVaxEgQEp6H/wH5WbIe5QPeFWRnv5
X2T6LTI8ct1zYLHtFuxcNKiHNx7kdNm7w036V+03r7yDrmJQVwftDAl/LZhw
yiUlduFUEl2sIL/uGRFM7lDBMJvzZgvnlpNJ2ABk9T9+LDF65dF7qVQsoAXn
1Zpty4nR5tpJDG22PfH9fgpdiB0m85YyngMzNMwLAh8BtHxI8R761LoKPTfc
JOb/x/MVj3Evo2Ai4UKdoUhdPzGSJ+bkY5lM0w4+PQohF2E4/D35F4P/HwcC
0SGl8ULr05GAM6v2Kt2GkKT7TfO82AshJ1m8Y1MHZz7OhZx6kMk4r+0L8kMj
82kdDCkxwE9YXrsZ2WvIIOhEqH3pHOmb6bKrx5I06o7T8uMmhejmQgbKHF9x
+6AEeb9GljSzgG79ktm0Sn3wqtxJqDvs+MhD8UaZu5S2/H5d6S6oylRF5pb4
50yvvkHF9JnghuWUpjgQNSm6842ZG4L0HIV7CQNEolp5ngHLbmR5T4KYlBgh
Y4rmoVw7VDKEr4HKBRIysc/HWCvNqM7a11N9lZw0Sf2JbeBgca047bE/x/Lo
bvVUhbKV9igHJvwYYlW9lPp6wrDk+F5qG054DA4wYA3z9JB4OeRsgq00SsGd
3/VO2I5rTsOskYs0ACOmsz/MdtsJsIcV+/SgB+Y7SEeX76XdmY8SyHrnZE6K
B2Z3fsOPg/IHSECVaKRlRGSVe7MVLNBcXqFEBs/wuDD5m8lKBJkaeBcUsxbp
1VcnQmxGnFenyXfa8rjsjjHpuPCjJKas9lTADXkjrRjzvM/Ip1cfc8zJ5GVW
CbswL0VYO/TA3pVSGfv1EjfxA/CYFndQveP3RtX/nBOHyB25nZy5Nkhi89it
OW2kbOVgHP59SrUMDz2pqhBWnvuWjmbrI9/lcjyJybtnlB8ou/0ywZBVjvRK
fbZGT9QZiAU74uhbIZc2aEmZHTT2hizMe4nO7PxcJJ4BJ5RkF6atg58Y6mns
eEwS9+K85N4pxe5HKuHFlNh91xuWGQJIxRdYXc8fECTYIGSgs3buQvcx0tX6
4Gr/aRvD/0ObulCumOE7GrMUim2St9czmE7CJVw89jZvbPdzStaZn/1U0sAC
CCWJjDlhnT6wu8fFKhT9Ern6F126ALgtZAaqLKz7aNUp7qCH+D3Zpdykz0g8
zNCTNQJEZuAMKat06+JbxMSno7NgdDPHmJL1BXjJg+tHvXWBRSdJlhPCwwi+
o2pT0qk18jPz7Bv1iU/AfL2YdkPSPxZ8Qeboar06Y1frhFGjSWdQgRxCPHB6
iQ2oOoFywYfp7Edm55c5XoeJmb9JLfMB/hFy9gYv6azyyvlDrp0ZN5x2lQGy
ep1LhDXlbhE1wxGEEkeNJV6y0LjU6Df+e9qaIb7Ru6X3jA1XDxFnkWBSkGgY
MFPpSc+9w4qterDp53zyuK1vS4JSTU11xxoUWmleHA24OnLwGyyXiXvg90TT
/CaMN4GeA23wsMupP5Kv4VHM3+kApmKMr9yN3moEXZtkQpN0oR8hfILDjhjT
XzX6Q9BPa8nZPS43JwNAd+YaOO7HDNnMfCi/69WohRsuZsfKkSyFFXcZMdd7
xM7ghMHwQMcQRM9TsqVTq/Sv/nJSEeZUOaIUkTyW5hV2LAB/1rZ+QsL+mcWL
Ywe7ulOD9swqdFeeYl5GIZ5CiTE+UFrsjDCNKKdbxNzBmEGJG9bIyurWArDE
B6RUW5Pb1/zBpCXVBU8wi/HzxYvoqHMedanj8C5boyZr+38O0nWRMg++a/H0
jRDW0HB+dTZCYPF7wSEjYiJCWei642ojtXI7cmkTu6LKkSKoAbF8wZE+iIvb
j7KeQkvlx+1D+CCf8CIxLbQf0bIeJTcshRFzkr0uYztV6FWL2e9Kq0P6vR02
dGeuuQJOE+CTzHARznbvlFbRKn5RYwUx+5TFlTWjGo4NWUV8YbPu/Sv4YMhS
YhRuVYYczvqbKbVSG1vl5SKdcmUx0alLVUn2UZTW4qw5k96uwjvfgiJn40Gp
aQoMAT1bxff/vArJA6XG3a6W7uPyRkKs0814gSfKmbic77DQ0CL9wMUOznAQ
/N0PRgBNwjIEUYG+GNXIUYMCeaHIHDSpCUeCzCdzdqhVQiZhxwennBVvCqLq
uoXkS0snUokUgYM0r7w5kRDyFSqcDoXtQJdCrawFSJjZLKkUO0z3Yx0GejzP
MppR9+riX3k1+wZtY5qJWYDaaOnXuWz/R5A6J71C57TYGDlHtcB7hscbIUIH
GeHLjFgY1MN/fMc4puNtcWczJVkoJFJBvkVJou0Z6sd5wEcGTnrVyq1gwjqK
UjRjO5CXqHp0TRTRJ2RvBpVecHEJeXJGbpia+YWyxLn9BBe5l2w82bNW+eZv
4zH0CyzoIC8JECqN8VRsDPM9GcdLCgxKvPfTZ0hrLmYehX490AUZr+2pHasK
g4OB16waHTmQ2EXz9efvVhgD8a+PIsZEqTA/gNq1PHNdoWfSX8j4YfXTzTrg
vetzPzIUuaJ+h+BYvl+gPu9I17fA8c5ufjvp2afkoWjtVoQw1LIt9sG+lLrq
JG8zTAmCDsObybGSQX68etP6wUb6OeQlnPVfe+44EAJjFtU+QsGqaJ25HFrA
UV+mSOR70bQtCqfVo3GTom/hdMWn8EoMr59zEHYcqw0qbumK2Q83JLLuJBvF
nRjzrmYAqNYq6SNJP1vKPyt8+KE9xIj7lCRRMU3LObrxdCy0Fj/7nFB/HN+A
QHF8u2a9DYNUdDP7BYky+VKOJuYRh9pY9nGZ+hrm0kvCZUXDoAQdKw8ZMp6X
mHp78y1beUrFJTiEvGPT6SxR7P/gln3ttYQs7F+cjj+rss6VHEA4wHDIfESx
BMfZZNQVYpBn37MEgsW35pjdaisOWCEus9Es+lOLCR0/nXOD/yNkfAqOM/M4
ua9a6Gbrzn7YQIjZcp+T+ZWoeYqK6LqZ5tnD73suQoBzCo/JM6xTnnLjqemP
tc/J+YZ/bWfhpgTA91nvS4KPE9XcAXgn7EFWW36XH/7KWNWG8mGl8aMZ0eic
8rM0tIamFHSKxXYObsBBJTZ4os3oaIMd6RIi6H+nGn6ZiS4FVVTGxisiHNU0
4XgVCaXb5iYT0OETsZiF5SvL7XDHrFGmr21XUzF47Zo4xawXQa3dC31DyN/M
N+G+MIZY9PWds8N8W5yseie4s/1JMdc3ji465FcSpXofpYN9Lw27OHzI0cLu
DPowb8w/l5TI4hFHBNPqeKabWxtocco9h8Q5AlZypTmkgNbDdat72u789Lys
9uMNaj32vtCQPlMgfKuEww5mYxZH/tsQKeS8AJYRWOn4nHhRAyDoL7QtIQ3Q
H1VC9APUPr9Jz3OCaJLGg4eXgXFm2qnW1nR9jp+myUAucH4trybGXWolEJab
v3vwCIl7KPMYvSjUoDu2O07hxUq+/fAYYRMiFN3s2sF0qFn/gdrFUB0X1ejC
BCTERp6OsI8Hz9I5mnca4yFWGo1TUvXbnR9LbSoLsrUWpBJDuEvWUFhBWlOU
QXDnjnig2+GctMi/jAcY7kqMJ1f16ttv8xFGrZczI3T8ieZFoZS5JOyqlubk
LywSWz3gxyGhbSQqOH7RiizjEHiCg5JiRZPaU1bZd46R1Nbs0iYAogEM7Kfa
dvSkYpYdm9QNYltB90RmoR36Ce+GvUgelBxWEFhIMmRV+M8vAWCRLo2mtZYG
ObjTO2fZ3lBbZkKD1Hl7q6xtblyqc9b+rt5+xK9GZ92k32kQD0qLggBbm+BS
W1xJyTbCmNz29APQJDUBT8ldHy02tEBf1miL1QX3nsenLuwTysvNGj5T/q+g
c0mhbUQRGVi5yEoovsu4agG2ivMd+2oOlfgbnUIJRqvYi3nIZkbMBJ78Hx/C
tocQML2x43F8mO5GndrdOc074rLsmyejYBsRG+IDaZDK7x3vRn+/o5ZNtNl7
nTt0VJ7vIEhPzTiz5zT+SIiX3F7+huCwEDn9I/jqPAwxJE2GKTMudgQPeenA
fIKLnpb0vR9/1VcGUVilY1otiNGReE+emJ89z/eZV96Uuh1xBjuHrlazEWWt
6nkLMHucmrXuXElGdLJ3mUMwe3S6JG04m5MjcA+yjZJTPOspXGvI7ZPi1hba
lKzek8x7vyjFu1I+Ak05tnS1gn8eidh/pITxeKKh1MmyrM1QM018bqGz2RFu
qYeBUahjVIBrcIYivm7Msnwm6KwHAYX6im7JQjRWC5tVFlcvfn92aShpYykO
AnLfLc0yBEUzErNKPLz9oNICzD7x6V++GTDzwTCpp3jvFrt2OVOFxLzlh/Ln
HtNDFil6TM0izblr1Ek0WZWDpdG1km+wKUgxYZFRTczAP/E+wpx/f38dMso9
1Lrcgi8jx76SXpOk8N58fuCg/7bNAQ61B4p0lVYnXmxEVepYZwQHvG27oqE9
r4003ykbwcCNlXr9V4mecP9Of+rbg+EBRT3VOH61WdBgTLDxb+Mu9Z+IWEgb
0OK2Xbj0j/95nziccNPz88+bFYm+3az4nZhm71IfpyUJqSN7xVyoDMdip5Ii
RtY0/8f3ie7SPn0N6ZOgRX2qXafMkqVwreNRYbOM5FSD8HYk304ybLd1RzRa
AYO+HOffQIV3FUL/q9f61Z88vvYpakiz6bj5QUREPOwBu02jmhyTXc9uopGq
8NS6/eAba1qLfF4wwpGgPqF8Rn9Uh2wBNMcV2HDBG68qs1akR6cu5XUfvBkU
3GsCMSJs65uNBOW48T7wrmBRLGCffz+94lMjnmKQeD0ov0LGgKPsO2ix1cTR
HtblySwMhZzyoUtuF2qd5ik9qJUBRnPUYFYTzlbfaDU/1BqcMoTQ2FHsDS0s
uCfz21+IVeXsY8jmNb+v8k/QCIq/boZTPJfM1quLDXWt2ef71kAWai6LEvwC
hf8TkGQR02sZr+CVkfCz4HhpsfdnLeJ/QQboNNxD2saum7hZhiQ6cxLhkTb1
bgyMg2tqMVifAxnuoHepQWMHL/823jz5SY4nXQl289yqB0eb24jlPHiL3Pxl
YtKKzXhKMjtKZHblA6KF9aIR59D8kgcsEgQBmNKPhWlQyVQqA+utkyF4bI73
1EZFs5LuRLZ8ZRzvSQeZdJJcxMGxU9LnmHQ5owf6CKvmcBEsMfWDMAE2I0yJ
ZA/2hHuoGOKQ0KaOh61Qteux1n/s2DxZZbQkLB/JnCdao98A6c6w6zZYW8Pr
NSkbsD0egoR250++9MEB8u3bUwxb+7Y+JaGuwF1CPIMiAH35vy3VIvQ1lKj6
PCyhh1tF0MuCs4GKK8znJ8Yp3zOSWkoYDKq42eFVs7dohF1IaM/DiBCkzJrC
9HSimHg0wtaW+Rx9Iqh5KiIhnoOM1Apdhl23zG9XxctML/1xRI9EvprXNAjZ
u2lpG7qo8GKlExlQGiyLJNpRitEYyPYlfnzx/jdSISILSFDO02EuwknCPOg3
Sd5gTn8quWzd6rSxIQca+UY3DKgZymnDlLrahkd1rdi49f2cNAOCD6cheAjw
a7Bu9yMP8natipmoZWGCimmjaZ73ix6ywYTrfOsy6lFmMvIhxKTKCAi+PnOR
faPlqmXl/KMa0AldWKFNwhNzcLu6CJw1c/N/ktPXFIY1ZZHMC6mT4JmVQ+Bm
LO80PL5RPtZDjeKMYfHk+H+msYZlODSfQDoIZ2QmgZIDYru/0U494V0CTqUs
B6WFBPeH6GYNsaOHQdNhZBD3ift9DdsUG7WXOMC5MYjug3Ng50GGYWmCYYmn
GHCsaVIiw5GXU+xVoHXReWnKdbyhUx0qjREJf+plaTmczKGG1liTVVL9Rq3Z
cdJcxPtRXV8XUeooVMpdqTfHyxO1VV9oqucX9jHcyMBLjMmSgKMImv/bjX50
nsMD09AxF+6tHKjk+1TAh28azOHNkb5hbbeRsE17QLVIXjGOZdyxsDhU0oDh
60+Ko6r28aS8kTZlI2Rmu5rj1iGjzMBFXf0jk7qrCxZeuQ4343MjEG8/uxjE
DP2jya6GU13ZfFycMtFq5CnZWm/HofWHdscA2oKSBvV7VKuEDsiEkLCjAlx7
YEkoAjDDs4rgYhYnpjGItNNKC9MeltwAJOQsjH/WvT0Qp+mkAhMrLCvI1b1P
cg0PrtoIcaqvpBGYD5ZVPgbRXdwQBCBmreIOhwfAdERQrfahBwBGyfY3Elne
7ZxxzLIkvzN1eymFnn21ykK7iT6SxY5Xbny63NpJMHovvE6vkbuh8pCPrRzp
B6qYR0Zc6ag/PCfUs7k50H8sD6ftZ8En4rl9QI66dyBv93EyzHC5aUZIkRMl
TvBfLAIMi1gsAdmAFwsC5NLDlYICmJXcPWKky+v71vG7bzMi4vfvZq4A9b7C
FuGFb0Ina2qpaGELlzHCzzUdIfBjqxTWOrqdwPo7nCDA8qBNfXgusAmXqnt0
hgdZm4c47KJu7XEt4fhiLClJJ4CJiXqRqeoXhEXt5Dy+IaRadVwxyQI0NLs1
nPfPFQGDobSuYd2K37t3RrwBznaRhdUeO5n+8ClqlN2w7KKEq3ZCgLcQ+972
w37NVnsNxLdnCyQ59HIhflIHtYGnedOj02DpHHILm3hK1n2EqZ25ww+yme6K
AUcV06CxYMUgzQw7OZcI3znwPYc5vIPM879aPdlL4cqzaziYOoKB13j6kxhi
yRtM5d6io6fn4qNg5m3rkBJ1YYyXGi7CD8eIl77E3g7E0WWRiU7baFDdhu6G
6OyRNaUjMEJ7xrRJE1/7iK7UlnXEcrEuwilnBwwlgZAndH+ejGIBvGx2pJwT
Vn/MNw8YvFKQS9kdCG8KnEmnU965m0eBEDiwHvKTFh2Ud5MqSqV6wDiJCbmA
HyKybBS7dSpeGe0eCuBnfbYtFGhxNcUp8kVzDON34n/fPt1W4JjAJCiVJ3wE
IhDzx0BR2D+dYOlOCZi0bzNhz8/MF/aTks1QclupvEp9IGLAsvGtv4rHMEPp
5FQuWHcEtymkWv2yaeo8Jj4CCW0Zt3CndPemgskuGUeep1xD9ra4K9n5tLwa
9AE8WTsh0fa6Cny3m4/8D2HQ01WglSsH41+OcPr4ia0cDiDTElYmwDl/Gekk
ZEVG8HZdwCD80XY8GcnBLgDoVPRZwV3MlCdVSiLgAWtS29473nvA92PY3us8
RKWtrjFIyeAm0pdvZIQIxfUGow9kwrJKMV/TTi2XkTYSX7ZDhkgoihADCcfS
b5mOBAl4yLvej2fGKz/BFxCIRp5azKZo8YeHY1UuFrBh7/GWg7d4rR86zp8k
DpBORkco050z1Xrb4Oxqy1cxCABwuoRgnWO7AD5Zc7wWZrkLiXZkE5OCJbcV
7ZBnoXJ0RxExdDM8+E24phzNXAXEaSewVyq72S99sJ37dslsW7SjvpdweSzg
KYos2oeAunGghizq9z4aeq/eHodX8shfiuS6ygLRh3LozrIklhdjgVkjxdG4
sVKZLSMx3n7/FbUvY26ykVGz8uYfXd09JaijwLCiXr+k88srRgcKuLxTLJoA
HFRsdxh8Lru1eLknp5XK4i9B42I5PB0qWNcf5G/BwKaT8vZ/0d9V8U/JBbWY
rIljDg9Dlm8pP2Jhbx2yuoMOS22IdpyZeR5zIkxKrPYxtO3UYX0dQvghw8Oz
Kbzd09skpWZPkaVECoS35+9/N3On44hpBlC4HQptTkwX5mKR7dY2suNZCEqL
N5klnqepmydfcIUc7Xo4psgfZkNoKwFwGEFJS/+CHjgFL/1zo4xi8Zu7cH3F
HhZZDy/Xs++v97JBDopaFUZDSkCbXL9a1KctH4fiuBHMCql3NM8MqVQATikr
9LjAviygAGnnxRk0j6Pkdl6gUKAfFJ0vOd855mIeAid9NugRSxMHX7DQsPcK
nRGx16CDoTCnwBM1igFpAXh3p3hPEkfjUGiAfeMWJ1n5vZk/DkKyYNyTchOG
hHDVfLTGBSfDI7/e89+L47R2h6JXZbsy/C9XvdHtwo1LjArB0Dt9ac4KSgqD
Oj2D+MQ3bV/nhx507egctDdN2UTxsrBDByX7upA+647duafZtXS6wV80bKtV
O+R8pWMsgtDbXi6UvFXUaP2VIbKDa5Y+gVAbhyMTTBoX8ESJLUvX4Jhqnixp
PJqOXJK1ae7wzbR1kJgLRqjtWRp8sNZeMUTRz+uULLdaYFCUStVsdM7iNcXs
+9aN3Lokq4AzenAJOfN6Cim5jvql526lpYk6ByHMChkgwrld36ECi3497XaW
ebYyWMKuGvYTHQFX5G7TO7Bm/ilOnn5M0EIvYroFNY74Tjla9Tu+ZPJym2X2
phkzNmGo2agr/nvyaqT+oM1bbcg6lmJU0IBlXUxCWxfhGohScDua5maMH9Wq
d77XCqRrT8+KKdClalN+cG0ZUm+xCHf72Pc+Aq17NacgPFSiP9VkHpO6aE80
ZboVoKaleHBtkaDOutSicPeroEgD3b6eTf+6rjRwuYnSEXgjaRsX7DAYH4a4
z4aMyfGsCd0x5zJGjg4GJCl+2EsLmiskltAP19KR4RX1ye+xRGdC/IWumN9a
ocwlNgPc0+xJyIvGfn/pIaQXjIcL8yVfZjs2sm1EMTlo8oiyjM4xXfgHsAwM
UWhlcT5KtFb55P04N9BJjsqZimhPOifOeBaSNT6E0PCuHyIkqB6V0ZfutBLI
toO1etentNFiF6OpJH7qcUEACfuzSPB89j7KEsBCeSOdUHdczMx/zJOwHb2o
AtKjhXMEFx9nblmBitkLLIiZ0CpLa6Gi9Xqj1oC9dcFb2T0eKi9vk+2epw4m
yNCeiL5dc/3BSFvI3FOCCr3zEU+akF6VHIYFvTMrQqpjjeM0Sv/rzWDloSN+
NgJJRMiHA+OfI72MvxqZNo1spekdOC1dD70bWW0KpmouZ8Wf2Feu5AYooiHy
Adv82ao9+kPIeXiaGCrUoo++XauBXVcrpvyF0L71iFolqJGcyMNdF/sibvFd
ZnXnTgdN5LoZzCiI6LZsS6dUwEJ3HagH25OiiYTy4bW8hxDMTu2zR07sL4Ql
AAXlGGc7DWiHncFtthAzBGpSGh10dQW8S+RTCkoPjhUu/s4FcuRhH2k1DOFc
jCqK+UqubyTZHZlIAzhzw37PUPCpj7F+FdfAlmSAGQIHkTe+NwyLqS6R4gyh
x2jRmClR1HqvvjxCydFPDeFy8q2uYwDsUgvK6UHcPW3QOdC6DRuKSeNWcmc2
PtuO0cK3ALOwTuUJZnucvEdRAeQuk01fVGFQN/3ANhmoriVpRzkt3/LS2Kwk
F2bCettgD6jPGLVMP4IcUsvnLujQYzvMvNUNjwByAlBYHMdDIiMY3J3jajIN
S8kjhfdux/zJeUtSg1JL7nmgZlMHZ8iNqplOKn0ntEdtjtlJA8IqvPnh7V0p
MMTphbCwq1A17Fm2n44W6KpI7iS7tyUUWqCa0/eDiwhNdUWMwVQr/IKO1rkx
2DfK3svCdfjtZU7Qd9cdYkDSsh6QswCGWGe2UGfwzigRRppJ2nfLv/mz+oHB
K5d+A3048KPtBGc2xWQ1VCKFBpSQCdeqNUc+9PJlVCEa0uEWjVZatvY8KaTl
h48E+PZ+VhzT0xGvXrN0svMh6e4ricakJefCpUqbze8Jfon7nLRnwKXuewQo
fGBpGvFQ7VsUBvoYv/3Im8Vy3jlTrQNssNoOJFYIy7FFMQhwsy6MwW8ySCuT
Fyrq/S1NdTZa1WJ/xqnLDO++k93JQVX+FcJmUdGQBf6Oilt/PnroL2MRZEQ1
Juziimr4MHRl6FhPeKlOIl6BWoPYcUBcUL6akBxOVGhuyPduJ1EOw0r0bPbo
XzKoAxYtmHpEgdrJ9wx0cBqC0SUY+4lKA6BOLw/ocmZfPzQeAtqxS+bwYQJA
GQMPY4ciD1Ec5UNVRI1VdDMZQ2RgK+fYTp8CZ/1QF+A/4eAdd4bHUQrT7dt9
oGPH/a8DG9t0g9X1zlG0nwnob4WH4+zW3XPkLgMBNviEpwGu3D6ZqgblIUPT
3P5wdYcdLMNofVj62It/zIH8REszrZWrLLCMDsYGgJPvj/NoIJCegM535m0Y
W0EHN6DSBbupkQWQQ+7wZqFx9P2rNpgyYcO5YwqsPRyRcZNl2gRmAAp3iztS
ExiT82f3OIYMLB7CP+RnKDExVLRH3u4M5E2Sx15XLiyaZBTt7zUZZtxIOcgP
i+1zVAlj2N4T8jmBysUqisxEseoAQYjRCNjj5XA5Cw/KCw9E5V7HbmzfqI8k
QC/pREGs+Wv52EQWA3vukdtNRdBrZzTOMkzhOsTzvCkzk5hRTcJTL5ctc7uO
jq3SQCX4mKE0PixmBa42NZyt4oRMG6sNMYqkBN4HNvbuJxa2MYdTdmIP+62I
iFtJTZWWOjatAnGUxtFODOPZHP+d4bi3mcHeHYYl1lgUFvb8lLkGAPdbQ8X0
/gIynE5cGIF8Wop5W7saGQK/mnSwrzw4PUBhIskDhDQR9QRkMW+HcZC7hDuD
bRpHlkA5LKQl+TVxDYoZQdB/imDBJAX2GzTjBfKtW3ZW9U/X36PMXPskclcQ
psvBa8t76ueyzW1wYynBEGCmdkG0OW+JMKx/uzE2FkDpcrp2Kt3yp5F5ZUW7
VYQ20GHhiPoFY1EYOJS8HGL040o/Ba8L8B7JTCJ1AJrdm1DuSzUd/TUz/cSO
0boX9G12OuSSnO7wN8NZATihvNPRa7VYVQFLJE56YtTjsa+yscuu/T/Heyu4
N9tjG1Bo/BT6NvpTkphLw3OuwD76vKdAVHD3i5oqxNmvKLAnknpOwVZgoZru
T26MHUgg2HSA+o469Myj6W9E9ZDXIgpUlgRoPy1jtOzFUONNikPzDxfNdydv
3HYg9gqjmv3MfGEYy1C2yX2UApKvaGWosk3iVb7VJ0YVSCX6xYPBcchR+G2k
wq+71B8CqhqA9yTk7yDU8Ks1o5gUdmLdZlui5aPYmcDEnk4PSVfXm3zmPZjx
mbC/JftL1cEIdfdQbfWBdy+gnKHCzQOr/IIVVJtpGBvAWJ/P+8HtygN/M0Ww
XC+nAtebiyo3YtX4M1xIWl8rZStNzrfgrKjEK1Kdj3R36a0OdQJ9O/m78We+
keD6njTvSU3zr4kqyIwZejZ2rEcAd2t5nvkdZLJRyt4qfzDOs0whnGAX8wS1
VtfJZB69AXFcVIsBDPZa+nmm7IobYAon/7f/lLXsnxbwzBZWIh4TB+LBqWbB
iRec5WlD3ZQWH50DhYhBU25XJR6Ogv5owHcvf6dcOchp2SvNya7HynjoXXHJ
3Ij5HWwSaNy0a9RSTsicKBKqJhor9q7mlzkzCq9/lPcIBi3sgp1vgWujrYo/
VRt/CxCmSoXrFYlMwX3MXIEKLuwsH6/QNFCAwkJhM0YbReoWakWtE9K0jqtF
RhgzdoyYe7qmvZE1hQn3GlvGbxMD/4TfeiheAhIDOiLsuWnSwY60iCFia4cU
1ImCoSC8JbcVvozZxYFc157llHDJJmszI8xkeh2NdH9vz487BxHwjrNWmsbV
L/rQGjLdMGFxgxu+IAC3kisM5PDsY6XfxCoB6tQGFEswTKj5FoDuoQb6OZF/
FbbWCqCWyilFzY8Mdc0jBkhJ/PQl/5Z4Kf2P8wQ0xiPHcVCgt+t4bvvzgv/a
9geN8SVgqy9EB2D67sDC0jZlmT/YYY8WBSqoelmj6Ub2yEcA04mqlFzDeZts
1PFs5aES6FCvh7QqbXNWgiWdzykKuvAMYTgBgg0g+aJJ+jpbHFGtumoxCF9O
OI4DSLKGIqT9kGrG68ZBt1yilxJsDuGJJ4qlx6Qh0dWKrU9enOaMsH4LQ/2R
RJPq5u1V8rAYlfNt6HHu+U5ytzzLcR6KaSr1mI6hnCZXMl0Ccffn47ni5+HP
BCGSFH9THlFlQU6hziUsEbow5aWsKzHb1dt+5OUBuwKT1w24LLs/3p8E3pNx
qTobEJJ2XnqYuRv25Y9/pcy7JboR6EbNyAztdIM2c6aWzLJVlINmhUh8r63L
YHOcz+TbJJ9NHPMOKkkTVnwHPd5QPROCYRoa3uCq6geAts5crMtOkb4rKre0
YBJyRRJKFFwUGB9Evy73tMv/5DxRrxwI0ZsRxCSicGPcctWLgjdaxnpkdq8y
gbY5kTd8kIl9BxshRxAm2xw68M8eeX5lA3Se3ucNUBReFlSb5cnUjQHqd6Wp
8uyZp7tA/HOm2WLE8dhPvkONUyoRgtRa6wtQk3TPAGYdIPq2LlYJB3QfhCDF
p9PImOeCDBb0CLW38hEuzPIxI4ZyiP0wTqhZUz4EBie9eekgsawvhBSHaKIT
UPmu6zv769veIYxgu10jY6L1od0MjcPOkTugJIXeZ027W0OQ9xGtXQBSSE2P
iM8CndIy3XdL9YAYT5EGHP2cdonTbvZPFucWIJNE7dCTbzdqGmEaBpaY+xzn
X554e92z2fzJ/aahyOzwbfhkhVLs5mt+KijA4qH9GVAahtpHp0BMx4yJGghO
99UyHGEmDWkjzxUk2lD4wYE8DzMZJBQ7Rm5dkLEvaeeHFoh7jDUR/ZIm+Oat
l8vk0ctnhd1Rz3wOn/v7PKj6e4G4in+ReHIz9ldmWDCNZ4BoytkATHztKJYq
MR1Df920456634JiY9A3+tVljG9dpgLqjavGV5Xe2Ad6eftNZzeXTT1aq/SL
6glz0HrVnIo4PmMOlaf4G4BdyvU7E2+punq246AxXmVWJ6orYd38jWSiKQb6
Wk6W47qlLTuyfnUklxyIg/eNet1VBNtdqZFHLa9lGkk+NnUdY1kgSBmEkZSu
R7GGMmZx5rThXHCWoKZRczvC8P2zf+cR0pptG6Yfx1BW7/mawLb3fIVTB8tc
wXlt0aOUvNtkifIz+0xzNjK/Fc7b4Akq1kkCXJMrUaslOA6q9G0RLxWG5Bmj
sy98W0rxb2TlmjR6OCjGq7sSo1rIIkNtnRFrQyjCMFKdY65UUDl4zcV/Tcl9
UJRGIQigSgbp/Z/JiXL28ldV9R4RpOKuniOyx00nkC42ZiRbdia1O9Nkzzhg
pV58j/MPL2RA4M7MvZ/T2hLlQVaMvq/XKnRflOhDKln47R2+knsvYSl12p2+
xmUrdJT5IwPqfmwPLAjON5Qwb1FmudWXOHEKVvdQ8l2htErSxPE8+PNffNa7
0acBKyZuGyZ077Kn1p2obqdnRsl17r48RabmUnegQOh7hTj7DQVt2qmO1Y8+
iFvibgkkqUUfYhuoZ4Jo5n9/UH9Z5P0xTPd533HymlrCiBPdgXFQJx1IXjl0
aP5LOtGjF3zBtFx3ft6IccnBDXRnWyOVChjsSGHb7TAo1Fbzx/DYZvePu7Vv
WPV6JHrGMkGr72pBQ0f7JQlBv2Vi0oUt/Q2sNbiA/yVXFn7/6TMQfMTQdbKS
Xb6Y2egqm+wVR18rD6mmCKUaKWlJOhcsNHjnZaMnvbj37LoHDleKr3bb0Qa0
mXrXTcdNFJy2MmTTZ6nWcG1rx2gey5d8H825ufABbRG+EH/lOHmnytRif2Ho
HgwjkCZouyGaJcqr1Q8/5Q5b/jSFX5S5fMmG9Apr+bDzJWuyBHPTnvIoSOIM
aOoFoO5vYqkb9qSsVU3YYIfctvHTCswzJCh8nQEYGOnNpO4TlIVNaUpzhtEE
QDQqIXv5M+CEvIPmJkGZn72wViLbbeI1Zq2LjLSPwZTILuCQDC00vYLaxgrC
iNH2tRvt0yoG44vURrLBAIAu8Du7JnFlCxOAAoNB4zUuVldM90iq6JdbxnXT
EYPh+/VOcsHNeV6WCbiZeyjDPJjmkO0JJRPZ2e/beVgDFe56vfjl1wh+Zjcr
zC7b5LXwzqgbFSLWjz99kqAY0cGy+Zq8Fk2uN2iB1Rk3tD+5jxGf/lHpVDfC
o0XiQJm7rUVLD/RdksG6CPE9lzs7xRYOQLaLgczMSUkqO81F1SPMipGDDRKb
JyMxsFi1i52ua8SRNoCzyRfPHTLtCmIabz+btColIlhlhcj9hE/DGEKHM1fO
GvqAOl3/Zfw3s+waUwL+B7AKwVf5MiA+XnzmVQUhtiIsdWEXQkBASWOx5z3j
OhusrH2FWwCG+q1ppXFFUUqZmbeak+AtJhbddq8txEQAIvWqvgnUYjZXsn6+
vd6W5Gqaq3mWq9zAexSlLKASV89b6L5jt6r+zSaDJoJ06v8m2XaS0qfkQq33
cXHEBRlUsDS9PNmWeBVLykVCk9wCzeoWDDhTlRM6uS+5El5D15nzEUyvST93
aIjB3xWnkPFtMZVuGMeGqm8HpS6+MdENxY/YiSLdID69Y4lZRnzmvQjo8F0P
bh+zNTK/39vTJfd29Ud/lbnmt+5qoqq40yeOOy4NxhAUORBsVTiJR4/ib26C
oXppWyAWQ4UnoLpacPADMX/Z5Nobv+gLkDRBGPfGWqNGOdX0m7lzeQsKiBXi
lxQrCmW+1PCyWW9hoOn3Txx+todk630+LSRHbp+SMrAx/rraA0oGrR9wRsht
QELoLF8YaYgGpV8w0likn9q0y61vPViPtutVAe6y0QMZBKrgUDKG7wJcwsXi
uY6CtMUeUlhOEf/drDe+Ic7NirXeHIRppaVSPhxlfmIPTR1mhEGvRXmpRegG
vaITOU+vHpTzeDoht9RcHiQZ8zATZqrAqHgI3mg0+mUJxeLZFQh0u6V05LsO
qRHiC2UPI94QamDxzzqwQ6zJYHw9zNOfZ0WiynuKndnF1C8tAsKk1kcj7pmo
8kZunPX8qfw3jYdv4DEYQxR6YuX4SYtu81rX/+y7zJBfaQftuarRM6WlVXMG
bRnT5Upk/iELX2da0qFszxDNysGcn/kG/FGIL+a0HgIKeVOpDgIq+LO5D8va
NFsj5fQUYiQrkCMs2g2Ituib047STXqm+3P6VASdxcmvYVyaciHdWzuGSeH2
6viz/eeelyQAdrs3jiuFRtnqxYCqZxosVWsJbriwZVA+3tw/pIgAfDxdgksu
YVLBwASeoqe/T+/uhtmqDow3PKB0jmoHYqTxYtXz9PmLK6DS3/5sPo/uZM9m
DGT9BgUjmM+yEwPgxmdMLkUu780O93+9nlsvIGTLkMXHGqjSfbAdRSVmo/tm
BZ4HX050vjHaqikQzLSwr9YTnkfCypfJEyNABnA9huflbYKwi4yE5kR0BdOm
lEk67e43dxuVJgMPbc6I1qynCcHKVHRLUm2z1SzmvbSBxApPG9tt8k9aGrIy
er2M/Sa2IGoNZ5MQgaffEeUL5DdxV9/yjqtYM77pQL0RUJWGo8iC2dF8xN1B
Qni+LWwH7EH8NdEbz0TVD3TCNDZjG2HUY3zqflkg4HeTM8Og6Nsk56GTp29E
iErmQpJflv5+GiK99DRfILNVOrUvfxkC6PX1LkJSP5VZpMK2zUyo3+9Tiln7
EfbeGQ0h6MU7gU2U4c3WuZFpSH6Z/TpeayDB14yyHgBb4R8JN02Ga0sp9EnF
f7+g/M260a35KwCcXxQ13TJjtIPW3vLe2ogFjYdrU/zeR4l0Ir9quuasrVQl
cga38EqOof0fKQNVw1gvxlS7TNG2kAKVu2PwtSh65SbOXu3whpas/jiWlTK5
EN4zZYumYKggtSXb7ZQ9OEf7J3vVygSWDlnirFD1zUtUDrekoGHvP2X8RGIk
KpReYUYiR82K29oDVdGBMS1qRVSQWlMXvsxWohHgiGl+E0EYFGvAzUPlNt8O
OsWrPNMUyGy5edrDT9YIWU42bmogsFMTDk8gRWtUHsQVDJHiqk2oJXzdqEv4
5X/igFKUpsd0Cb54oM/QcTJX2jN3UKZvwUBeWnVml39lEwFZ/bdzBXN941U3
8xcIMMhH/lsWRoeRWJbgawqNsTOGJEntqyg0RynGUzh/ligZK7NOzTTe12T+
xs3CgOYs5wM/wBEMehJQvA5XBR7vQ8IBbj+uR71bhA+Fraz9sFY51shNhj8X
zxOIxV8lyaK57GSHf5BZrsLAnktMdknYB1A9hLxVbTC47C9vppf2H+1Zj8lN
gQEn3mI6n/RAoZM35z9OcGB6bW/fqah1vm8JokXPGDzgumQMhgemi5x9jXJZ
J7KdwZqqI4dXQhrs/t8bwYP0h00xU6RoBsj5Hgb2bdwHmpyshTHqVLO0FfZJ
TvtrNmkR65MCgVc4fJaO9d+XBo/hC6ZCwzY4PZNhGcRm/QpN86ZomJVh2t9d
ZI5Rv5sy6CX9ynf2GyYhD0FJyQhHDdhKpdqBT23etLXZ41D7y0HiopP/EaSg
lntNur2L1TokCz891zv/JHGQI7wuavATfa5gGuCzl52DfWGhId5DxU4T7E9L
ChFovzwFfDjQyVDsUrE+yL539R1Vi9+Vx5LrDSVC6jyo2HjEp50B9KnqgUsZ
aUlxoIWEmWS5cetDezs1ZWdK42cZkD/TC8lM1SPlNgRkC1FWh4XyyQZu58TC
QATz6p08wa8kf+fy4k+72Fz5rzTZ0ULv7qqgorlVSANZxNtdMPgxssrnKPkI
rwGp5YztfbDunn0Sp1NyDvwMt1CfNBai2HJaz8QQtAZ7J0OgQdINl7xYaiyg
kbSoauc2CamaEiJnXkRfpLN3LtLnZWamhJXCB7QKpolNxW6Skx2/wvnKX5QY
kKhWUJvPjY2ty51m/GyafLI0hYixsV59N7Np/nTbM79zSZm7WVHxKUesCH6V
HYYsIrldesDLoeeFvKgCmygp+S41iWF9BlbtkfGjXBFLrh7zgpWilJ0ZGkuv
H2Am3H4uHDLn8WIXX7OxrZbb82p/81BH/xJ4YJo2SkV4nvMGYscTAp0wyjCX
7Vl//Osj67c67jwXHu3KzosXMCqqTqfFkldzLfpjQ5hQDe9h2R2vbpLkhk/r
01YlycVMo09gILhPd7bRL9UkLqVmHJmB6zznXuiAbl46hj8Hivg/qX1loPiE
pENv+Gda1fbvNn4Z82Q63mY4Nb7+Pkk4q6MJ/plV1mFTHr+C5fG0SzRGhFEo
UxtQ8l4f+BkiXHF9e5d5tjyHkH1mV3//TF5dhG88aZHz09Jwohk6w3msqrx8
s/2zFZ4cNRwWbYr0ug+6xCfResPUHOL7liT6T3K/pC/tWFbfsfJT5qkibXtJ
L2JW5Lm+/H+DFMeEe2m1tXo2fqu6PUwnt2FwbFIzDClIvaF3ky+KFFlOy/d1
IimzOMA7TFuijgrYq38sNUKY0xzLdKgR+93Wfc8XFRIAIHAV+XiyucYdHTi0
Mb2wLDG0D76HNXkBJ68AnMTYplgwMsJDPNxZWkrpc+/9PAb0MA2Akjw41mmj
okdZwUcqAauXkaJtZii8XpKX78E5GpKLAIlH1crTwGePApS7L/6nI35Cp2CA
XuKlJ25OeZMQixQcT93tt0sXjNyByE55PvYdwVkbenWbkXw40M4pnQZQajDF
La4IXI22fFlrr6QxIjDBYrkAEYqt166hy5XEpHL3YTmwVl4QHTBozkdw1ySG
vb2GkYXi1CAjpFf8NcOGpnd+NN5eDhnYIRU5zSYl7lGRghoMpJjFoET4QozJ
nCwmesBEDnrzb1gJiG/G2nHeeGWMU3RbqZrCMSMiL9HNjXJphV9KaNinQFy3
1HWgRxlv875YDbgxvuDIrIqpjIas8XcXe0bXHtDuQthkiL1AhPjAUdiP3z0m
gzKMAeL98Tn3E9DHy48hHs7uWDPthxNg9EPP9Vi+mhLXDeUsRk00SzaX2xiY
nZ8YkKVO6pmn8aeS5dEwAdvjs42eqrCzO/7DG7k/Uq9l+JVH572pR4l8BRfx
O+iwwt1CjgDIIwTUKVLWrLYGGIJB3eyeZjR5wPG9j+DsfrpJaclsJVuDU+dq
6GOlKukspnnzDWjTcaapuVmI6nwrFiEF1F/oBgTv0AWgBSjR/Fi9xIEdQ7wj
41Hb2A1+GRtA29XoLNzpAKzhR+CrH5Hb4SrBAsHLC8o0ZKzXE7CqsraIW3Rq
qih96k5sSBz+Gwo/Sm6fZEb5x2EAU04iz/Q5TuQim3hhntt1qcioy1255wsq
N4dI5veU47cOqX7Qzy8vOov9xe9PvgkDr0nsHRtVbYsnGFu7fiAXqZ6XiuM/
DWCQ0S4T9XB7CGQKbzW1tFlS0WoeM64J/3ay+C9bdfgxg6fdb7cLsP3aodzp
82hAGSIfm19QysWkyvzLAwi4ENdFsvI/8K0n+zJhkoD5vLApqVn3WXbWXlx6
L1HOdJ9syvMrQ85aP0M4sQOTKw41h3mFDppZYFFSGb1uxNsW6HuD/fvgeQ+N
z6xudcXePU6zw2+nUjgGU7Ty1s5XhqlmUKdsmgSJe4a4NPcyNiGTDeBrwER1
cYsh56cTffwWpqp8K1xnsXUuJiaErTeYlvS8pwTdmIVoetmN17l3d83oOsWy
ShFPQPC1naHxVc8FcfcvqXKGEOx+QsQ8kWCLAHCeUmI39i8Qt4Z2D8qsxrLz
OUQhWJwGhz8zgGvF7ycKswEBUHP+vs1sdmOFas7dJo+oSc5eCHCOc2fpZxDq
zhM28OTyFdsSYAj4ZsnkwcvTA6HFW490E6GsTRDhj+0TfDQ/h6dLoVMEnuEi
UUWPg21MjTnCQ/OtKyCGtsRZG3fBmMNjo418Ymx/G8SlvnU3IHpOVuImnaSN
KihMbPZLhgaOMqvFytrUPgcWgyQH8tO+qLHyGaqygTKKwGo/WGlIzvKoXtsv
8MWmRiOH2LoiG5ZX8VMJDOAzQAIsFEeTGWN0pEZyHoQqYgxBgyBfRSqDNCXm
VHR76sFTGnErAFkMeVirU+2xTuycL9bZUuuScZ/BjRMBERBlG80s7cPw+gR8
IuOosvNNIJAfUeb3rYm0H9WzCTkejLt3xovgIes8wOQ46twJH0xZOrhfkVNS
HtkMker9uFaNB6GWrfJfkRFXbqLCpjm4d5Vwai5BxTnWQuIPQNKmAQJ1rZAT
gnLDuGkCrjbyMhvABOlWw6noc4gpi8UQm0Zth3mpJM8V9ygGOxha3gahqpPE
NflrKiXU6cpG5DqEwDlWmJH1UVxmLTVsKiLx1F00cZazOKZghkg/KXw/Neju
E0atlvFk/ZTtmxoOZ8wgS7XQfia/v7UdsdrUrCjGSaM6MXnTaJuwBGk6I/Ag
VdxzxYhrJIsOvArLjw6M6BtrMHQYo6kvO5zvt/B2oVQMu8hetkDN9lWvijND
ZkeJGD4j1D4/oSxZb/iYLZD+ztb67oZgOdYYjYlrAM4tpH7I1igJNo3QU1nx
WfIzbwRLpQdhTini2rgZ1oBcQTgjQogeRg+kDHDmB/6OKIF8HApH0tFP/xCS
Ru2TAfYmtLnFd22T5lh1txtn2FaQq6/ludZEQgFfek4Et1sQilPlRhgYRRh2
Kq5wDNPbmnOFlfZp4mg3EtvIxzPt5nJ9tU2Vc+mxB0o1ULW0AYFO3/znGQNc
75ggimVAY9uY1Jcgz5Oo3+tmmKHRvGGywQKM/SQHjyyi1Utv6iOUjqwXkm7l
N6zoXlvU3F1nehNPwOdULIwJ00RAH0w/XE3GpKQubsgDdxzUDUJrH+Ilcv1s
b+zuUemSmfNogGJ/tFsnF5j42kchxcRxSgM11XSNfJIGvquHp6zhKZkgnCpP
cO0XmlxWADLVytR7K0gaAOUTiFdo7AbFfR4Tbkp4vWQJ2j8nwFzPjKF/p9Ep
yUihHjGNcsgvfNDywkbAPMZUKkhVOw7uibyGb/gW80e2CFuOQcTrnzpGheTP
n+0nFqD3PSJ5vE0QhDBWY9XohM6oCkIbrFBQvwIem4Q0xhUyl2aBKNCEaikE
YXZ7EJUyARDYRiorsvTVT6jGs9yAPZzHY6IKvjGOAb4H+OQlX+L3bNG7Y+CZ
tHsd/8s9T6wJ2BPFzc0zQyZ4CZpSyj5hzeJp73qogr1G9aW81KJFU8vCbpXO
kuLg8+/EvuDEmILT/5MOqQeD3QX1c6THUqDc9dKH2NCpaPAXHICWx6+rqM7B
tB/MI/okbSRsxkOR2dld6pt4Vr2sDqEdnB/9tXTQgq/1VkLL+Z9IXpx7cPlX
i1qsRSlFHr3WqznNhfaJUta16hm1M/h2UL6iC2hI6AvsDbkgvDJWBbgvx187
CV95b2w6t8xxxUH6h/jG+pFAK8odDKJPuGksFdEYamTkPSGqMFHOOY0w4lNV
nXH5Z9v0ogmgFi59rPoizOUJAgh+Z+P0slBAQqMrm3oLIr0ii5wOtIYaGlE/
zVGvtqCysjklZPLnMgJ4wSMBMXYszbcwmGMzNCkpGtHTLXB848AGTUZFHCne
jboQ/UorAGbUuhvrtzHF/qxazZQkVqqwOzcdN3AkKHoQCP791M1O3gBGsGIc
rTXhUcjPpWR+gJfDqeBUG3qsTlMCo1hEJCNO03jHSGRMemnhEu3VTPcSz5kE
AfZTtbANRpjm0pG1qKgJTGtHjsKlOIp3aj8SefnpggyvGIeHVDapXSExsuR2
M9jHbFvgthSIfurMToaKE8ZZkTrz6qrePnIo+CvnaM7lbAwVQx7r1pXbfLXS
vRbyTuUERX+gUWFws3YbtqaMo2N7zChWlBMBG3Q54sKCLikCSjuSN+qtVzru
DuXQjSX9yWlw4SJlkkSBD4REHrT8LAxA4jVrF+tKuHAIt6Q99Sn4byBfEDJj
Pz5V0OL4umioqjix6jAnAObZ92b6MIVgMrvi/lF7loyF7PgIC2HYBu2jIKsE
5iJlu2KZ1+smyAzy5f5gfoB+jPzZG6KrgJra66yrPndabOpGWAENXJTseNo9
fepaAmzYO02kJRld8g7jeqMYRA9rYsS/VkHEBjS978cryLCadwSPte2W7si4
L/Jem0Q3aKByEvsjQjLAe8xfqnC4vJ7O+Cp9dnVLQw+8HEdz/oTZixGqsMrc
L23uxH9FFj/oKiYrnnO7KjXIxMt+CXiCTJ0E711zntIIk7vBxeb8iurrpHXT
/EygVzqlHaCYHhlsliALSryp9ffDOV4fLQINQ+P3qwYYOMLnwKENjnOxX5lU
xtATrDrp9oWeYAVe2OFyBMYDpnJWiAdOrh2ceEH4v2zM7J/Yd7JEkxVGQFmo
pHFE+fTvwg1vaalX1qSvwGhcF5DftNQaaxVL0kOf6D1Jio2TW6+saDk5/zFD
pHEEkdRGm5C36K30bbCKprKCwn0y4GI1wPz9Dw7XZVi2pgOqmO+q8m6786hQ
TNiBocmmddrsBWEbqf54oyg8euWjbRAbXITWoI3OBBtPLMSYloJdW0GTB3SO
yOReVSTqKgPtw4OH3XhBC2JOiHvljV5Pi5q7INiak1zvnA0QGeNhKibLlNhy
JpZmkEl28WMvAa0GhHLAgFboGFlksmT8QkbkL4Du0Y2HBuhnyzOzmEbHSA6q
hgXGVwkbPlIk1GAj/sqda6bwiwqpczd1raNrXtiE6lG1CFNL7VytV9fV2Jie
bPmbUrNedywHC8+uzsx7bwGt8FC6WIkGFdkhWEDFp0oFfoSi+jXLiDQNcLlX
A5PEArqf3wBrmClriyPB3AfqosA8sW7JwSCHsOpM8XY/T+aWN+2Hvx+FzDvr
3UIeS7atKLp+Q5dyaDy2jC7LSfzETIdnV5gWixs8pbB7TsPyH8zgtdSbt5cY
jkPQRpiGnxLe6e5Sy4SwU0ghwbBggVTuV7zPBIY3KmiTj3LM6byHarMCBcVW
XlfNEWWycKT5Qz+Gp9J8/UUk5LlaNtbIS42IrTh6zMswH2f0I+QcjlCJBfC/
+p+28Fi06FCyiUFijD/DEHSfhsBlF4r6+lcFRArlCoemTP97mBaTGzTDJVMP
JpeBMf0tZB1miN6A+eN4FfzuWfCeV/vWEVH4wyu7gjuJ1TRN2xOgy1UapETB
7aP2oMt+w3PGRgK4XQVBy6Sz03TzcQZ1ASHB3VQxj3B7zmMKLienvm+i9A8Q
juRcNctxrI5GnVr9wCq2Qv4yAWEhAYabKIiSvrLsNBMWyZk2AJdw5OWwr1+G
TKdUbIyaww5W4M+yGENcVW3hd0ad+02iYRAi0o4jfGS5BcxeaOEAsPC0qdUd
0yS4kZ1+1ZFTJ1Nv/5FHaOqg9LRzT+W4zY9ObmPm6iruhA0F3way53h1zdA8
qaRVgTRsqfDpUs3oscfB4OY92CiwyWfiA1yQi8UTzamzc9DW8w9o5AkQimiO
AG3Ha0+WVJYgv5pTCucQQyb6zLEw2JTtjrGhtnlVh1fUfE6He13+WXg0lMUP
RjcBQV//buPuMw1KP19x25Mr0WNJDEJQG7rz2ABWDhWLBRWLoW+r/8841qEt
8IXvj8b3u9er8Sid8pkOx+XrMsUQA5gzjbNTGeUQGpjfC+AdmCW8dJVjqfLL
KzzwByoPnR4OOv+6Vs+NKd+PuWGd94dN4C/zcOZR5sUtlsDWlghkuRjF/Jzk
Hn0CJW/P0P2lvt4JTn+UwR5kxlvAvAuCj40G/kORv46xKUh3wjlawCHqy7Ap
5TL5U+YtC1Q3dIOziE1Jytff5G0E1gQnlFUvh/j8oov34jsUUWA2Z3U6xxuX
/M2kq/qAYqH37bk2QqbRvbjPdwViJASrQXXi3GzaGSmsXISUaSAJBhrxRBep
mGsq2a8BZSuu5rg+a5ahdd0FCUhrLqpLIMcWYh86SaQCNj+A3p1tW2ZnepA9
1OvK00WeSpmRa0TmuqeHE3n0K+75q9qZGNr+PluKzg3BEYsSscOTHGKwFybV
byS4NEa+RhkdBgq6FOLPXYX67VZlgmuff9jhUe/PEcHFEdKxHgxepOadqFS9
IbSvQNgRbwCQeNJ7lpUqS9Feon0S4TRX7gqqsW5u2E4n/QncuzbeM8neMqN+
G2lFDqHJmn7kUPHHekNZ+/UOXD49WgOFBfkcrQStemmmQFY3WxSUuZtJTlPo
jzhvntMBAHLv1qrkdEdybDDmhspPzqu9JpCQSSuTvelrMY98cPOjEOnx1C+z
BVddOXEJqrL+x7fcixonJeVi/WBblGyg3tO9IH3kHAqKSZwFoh3Vvs7uwXWi
AamD8n9ckK/bWOYQCsT1v605mEbHts4oSO0gRHkz67HMi12BH6xsAKHXDrmP
30MDdFyZYTzlXuuVfSdLltTHH8pDsvAqAMYY1ZuTx3bEMtIImY5Orth6lzqC
DVrJDvCIB4v/Kg9w9nbTU3NTIzBFNPxmqbMUAqCV9LPNgMgTAwqxXDIFBx4F
yp4GvzvMBsa6YUMuTPtRmrYq/d8dlS1tHmgM/CJ68/fV2y8kA2jpoXzOJmPb
Q4EztK9V2ecvstmzWb0FoUz2GsZVMy0jWcGEEnOZgFs7XGz00Ayd6CZVJwqe
5n4M5YV1omdg50DszjRUOOV0pM/Q4f9Xb1D/YP6nLlICH+Fi7XyNNu1RGJeJ
u8adRTjMVpArDb5w9PhZrnNNBY6H4qe2ob453Sdf0LxY9icJ7evqyivOZFK9
KENdGkyQaCGMVgEoZpp/j1WGkUKNCarq5yxC5FcO9b0M7k/r2ejQGYQ5tVYv
80+De3L9/sQGIDzt577Y0Gi0MUxy8Q6g/YKpXU/2bTvIffI+GiXkgDDfS5c/
gYwp6wRNSi4HpRDD2KVzrwnoGAe6BYHmHzhi/Xe1ktjwq4zLSxgPlUY41GWS
gPg6HFCDZ4jeMgqPdo7NeqP7zcOe3mS065WP2ZzbADqGSBFwkGAyJs0n16UU
mfkslOiIMj3LGJaWxinJ8WLV8kE0xqVa4ASSxMg3d1dl9QFfSDFipRxU8STY
hfdVePqlwRaXSt4xfFAZdd5OU3hATS62cZTJqhWUpMfS38OwPGQl8JNlTL74
xl5sUwtEEMQaz4wXxCVnSiW9RmYxS7RClaIaXMFHBTzxsIzfnbdt6hmIZxWR
NCxxHLUcEElSwZ4md29dFVDFWG34ZwHfeMxYB+C9TUiXqP+8E9NqrCoUOuqe
/j3vx/DdqMici0tiNvylynyRU6FExyV+fBiZQ8TH+bJdwZSt5+JymzFG1smz
uQ88U79mDte2IdsyWN8NMQ3nXIZbaJPEfnZvFeZfGlJbzsyMF0oWxCs+rmQB
lrzit/oXNmm4AHRduJ/ODa+yy7qLNvRdUWJ1x0mEHe29z9j32jrs9mYUr+v+
ajsHGTYriQNHuT571APWvUw4zHn8F5F2NxH4YZxa/MXCDk4xh0TeSDLMJerF
2Y1BBUxJImug3MUT0qdHJdreUtZIh7yag3Z1+Xw8Tqsx+5a6JoAfJZ7leDKK
eFbQnP5T95cHEyk+INYxSlSfZxtp7+W4jZX6XiqEJS5G4hOHRqozTeR5QsSJ
iZFBNw4NFKXtF/GQptiIIv/eQ7JNlxEQ5k1bNd5ES6ScYQSGb00q+IHctOSQ
8geb1OSSBHPjnp/1VJyk+cuZtbkIxiOa04JXMWz9MLs3lPq8hMKOdDo5FNQn
AQsx0UVPXSsPD402R9Jy7RmPRph5UoAoDx1oylRXwJ4f/dBEnJ+YQ9w6U5QW
OrcpAdLCUWVR9fqbfasIGZ6rmsowt7ZW5WmfMvwogHyU01ME4nO73WCDBQNW
+3nuuYOy8Bi484T8STctIJX4s4uov9BlRXD351ePhik4OqZYTuwILYYgssd+
P286GkKC5aNXClQ+E48lBDzgUC8QUi6TiI+tIZVmIcd5NRsXAOvqNhOy2fiU
xpeKNN2sgD0Or1vQ83f2nSd1obzgvE1fnyNzY1uWnuL4nPqXPVeCqlxY+bCm
NIGdap+Ztc3ZH0vuV5tT1zKGDXxWIgcRmcmEoExeBOOWO1QENQ0M8sbNSin8
VnUWhl5gV3Sd6Pn+rxJEV/JtFWj1Gcot/sy8ceflmqle7Ht5RqB+0+ch2OaN
MT/YEhIRxVY8NnzzR9Qlm6lZvUmq3He0GAN7O8aISRs27V3baNHtbBo4BASM
Hrfa7DK9vd/sfr77+p187n6MPvkpfyYYyVQzKp2YYD3iWirxrduRnnB3KaE7
TrmR2kH/OL6YbIUlr3q0ycpXCsBmBtM2LvbwE15XIthQaXgZfm3OT6/yJs5I
77vU8g+lSwkreXwloaG724zKLkhoRarBaeeyzi8oFVWALB95RpkrA5kofoO9
Phdz5Vd8DZgadxhYK1Q7go5Kslz0hKDuqhRdkWQk93t7CN/OxMR/UFXQylg8
b1JTawcfyKkeeptMD4XlAsknGSapyKhsXHbv0+umHP/XwmAv3oP5mIRLo/vi
ZUX5oqC6Ebzt8F8qzzqPtq89LtHi2Ye8YBJ83LCUd7KpGqmMlWUHFx9QQ8VN
RdhyDHKIlNbXXStPv6l5dtHYz3ZQ4XIFG9uWcRGqh5d3o4Kv8ErsvzVJAxgf
tJ/EIF4D+xVPPGv5gV5HkilebXEKR2uxfN1Lj95NUXIxVrPoQvLOkK/VqaFM
w5Tq5Z4hxK8Mf8Rhu4Mypvdd9LPn7Jd0gbfXoxqnaU8xfMenX1YY7i5q9fJc
VzxXAtqvInGpqq2rwpe8YLfdiuOZ3PuS5b5kErT26a5NPPTlKWwrRpBIkn0A
5CIDyy0y9GfAyefwTw3qoyngasLBWu+xnAbGF/eGWAOjHC0mX7g2ZKYAPm0N
XCuDfM8r4hhEnwlixoOyVSh3PEYTOhQvaG7rUwgvxFsFBeSezyLR9NjtnXGA
2TfJ50zxPJYmK+AaUorxFcBgsGS7tFRwH/12iPY9ycTZGh/WwHmlJWYFsWgm
5JjUxx7SH709mqv524vky+WnaKtdwe43m9xtdjZdyqZVeiAmIikDrNZbTo8J
JmVHBqxWKc21/tXhClSx8KDcRXaE9WH+wkifDbdCP6tYXWwyqDDvyPNXJGJW
V3nk5Bo8XjDB0tkDJDFd1m4v/M5FS5qLk8pn7xcS3gglHerJ6SDf3yKDtcVZ
fYarxGcgUF2mHuYgREzkuzIJmlkj7Ah1gxA/HBRBOSln6ToZ6kcakFJOfY8n
F04uix/+mxJdkWntSzMRy0KtXDMynv8uFS5W3ChSW/z7XksQj9LY/850pzqv
lOSH6ES1vIuGwLW7VX3SdQe5vkdt0PH6JSFZDCi0/CwzZqkCMHvY/zDGSxts
uJZHgEwG/kCv0PhFGk6XL4YjrMtUPiiBoxQWfmQHdYSAatrt8eZAO/5Xik2B
bouS5Zflb6Oe0san88Ui2vSXFhhBoZ+Oyl2NcgyhZC6dXMH4HaFPQNShDWZ0
M2/UIkwYsqXRNBrl4Ce/5jdRMssfaz9mq0optphoT4xDfxM3SLsSKCiq4gjY
CKX5xhog71x7i2CKxqKHzBXT6CaanStnhNwtXj8YgW2w+umMNPcDxL5D6O3Z
AtBO7LwLlrISPj08mYT1TsuBGS3W+5oQmxppdyu275JuBuoUaHMyoUmG+AVu
qVzvDpPw0qczgPnKA1/3FaDZZ9aobRauwoIa9kEcbmYSU28YrBPXemTrb7wz
HEzgmzyyp2STJIUsuznSG3xbiKGr5ejdNDVvA2Crh3li39+Ct4ujvNmpAFl+
A4bbJAfK2cbFNykKx/tyzk6a9dk3gPYuj80TNYArYbFjTqDuEjv0b4P98slA
PyYsI45NpmBsLmdVZcuczri89fdEwPoNocg8v3XOdZ4TT4A38v9gB1HkcKYL
Va4PcnNViMdxXane/LmvhHdKXuvq6l3y4R90juHgZK1mziGrI7HSMQFuHWN7
4i1u5Armsyqc92qwft5IWQmoWnJGKWWR+zgM/4oiGAbRVHmK8+cFMQ5DejL1
dl8jE0ZWqU56O+KOl1Zd8Qks2uktQ/1/kCEW0DjouRjbOwqLbDw0gQ/L4EvX
OHL0B9igb1ilT78J2z8jh5z5FxSF2L3+V4Qn/KlL7Abcu+RsDxctfjJN7a31
miMDIdtRWJuReTrOQ0QqZOfTecykj78RMiPPG4Vs9YKPiku6RF2HqeRMvuiG
2dzDd9HTavP2EGeI6dcKigD2VdKYoNCglBXNYyOK8fYcgqtqldgBV3vbIpn3
K+DqPT95y2kLcIMWzrCWbNu00arIuOAgittRxlNTisZENRLuK+bEYYbEOuus
Ir1FJECFCBvFimAMPmHhs0KCeksJuMZEsYpEvbQybrW3FLpbtFtP/UejDAZ6
tub9RvFPcgZ1nV4g8IOclfOL6qQrGRfrsQN1h9RFzCU70hFKBe9+rjb3cwFv
lh6tZ9T1y1Y0SZxxQMJ5fRHRvjpqRs0fY0MRk1PN3Yaeze47G4C4ofaWbsHD
47CiLXCxSxmInGcPxdrPNeEdo1/52nsxph7BlxtR0dYa297pQphBA46e4pxE
1C8t6ghJWzWMfb7afresj3cH/YhdqkQoBkvR5GZSGHdRHHa0YFokzBEqd28J
4y2pqLfCA6gqtbEszpk3ui1VHe6HOosdQaWM1cBMYwMNWqWv7VCk941BQPdP
7ORtkgMOxX8Bd5/ztaHMZaBkket4e/7gr8czxe9xOc1bwXH9Z67Netat/06u
wdzlRDs1AX1itpo/lUWQ25mBZOR6ec6cREnOaRzPWJcTD5eBbH2VhBmGA1ZJ
BTlgzf2VIBO1cn0SboMZxgZv8tTdYo9CQmfEsZ05WaZ67wFno7e5BIA4TMyq
WBd/2AvAB0xkPSQ+i0JZtYPctGQ7VmOLDB1jw/2Iis8prxDsfy5srQqHXXSK
Oy4vjs0uaPt6K39oEiPvvj7jWhEnspJ7dP8VIB8TqGycG1yDzdqDhng/5PIR
74LLaiA3i0QpOeT1TWPXmnHVaWdYTca0PMFh9tbedD1SbFNwJs2UhG4EuWcr
KtfWwXz8rs8FBgnWH7j0fL1+dU2it0FhomUvNKq/A3q5DEyzn922p/bFej2q
kzuo6bMlA6lukXkDYsEk+t1lsF4LbVDSQoK7hPwEU2TACLeMO7FVP5dNe48u
cidFcch72N+O6EOgGFtgrL5bXhQyrc1FDzukFf86mkFJt/4IKt1li2Fe50fT
mCXH96yooY0hhcpp1SIPEvnDKufVTEEh0B9h+uJDPv13Vzkx1Rp+SiC1f3N7
dZ5wuijk7Wl/Rmh4LiFJkf85Z9nJYS35pUqjInAH2osJO5bPXxhyJ79kU14b
TsyMn3EbaQ4QVl5T7yE3PhIguNYZnFwYiUzzlfo0tJOzeBrFtC1yTpbjy0dS
bychENDnXj3cVIMw8MG5SgyJr+ZGmZyKEi6rEpq71BSWK7+DgsPuSO4Mml5l
7FTVBjJg5M6l0YwnIVZLp0J2v7xZSdTrhMn3kQ8oIPlta8tjJz01ABCfgnVt
yAxRvHH6G9FXAgjMFzXpV3UfGyDwKvwMS1LHfiNoKbEFPGFOafcLTCUMjvZE
vyYjCRAAU33rwPbECQ4AxPIgdbQws5gKcYqfeWyeTplKva/niR7Y2Jo/ynC+
nkttfPwFDv5GZfLLuWf1gxFOpBQLQf5CI2mIpED+SmMMdotcMNLwvFh1uPtM
npZ2jk+NnHgrqCBdIkJayb6P+DBLd7D7irRI0hgvVIL3RibtTghYMT5++T0c
qhjkeLXaCoJlZG2ZN1ZUe5LmoDx6dM1yNAwt/8WFjWBbmM8Ew1GFXKYneKGp
eA5rI5C9Uzy/gdpsg7X9s0qFSzaVbirqdL8t19eaK2K99gNR0EDdgc1HzURg
/qtJSNuNSDSr2YHYjE3ISwvxy9T4GoHGL1sndMHBmB2nw+VDT/qsAXJAq60G
QJ/lYv2XRcunU5CIQxAY98JjO5ksvXzBV4Ol22bKGgZ/icW+QpLYFyKjmLQX
1C+DUZ89G1ns6pr+QhQNu/6rj1wnWdfbyLCmcg9RUIGeGv7fF3EZhoqmXHyU
jbJNONz0+ZPRA9Cnz1p0PHQr/Aujpw0uj3XfvU+lG+kq6FTg3d7IBtFSqTDD
4hEkE3c+ePzo7BHtNhCPX95S9PzW0+fjsdtbenJzUS+Xz0/JWriyLoeFy9lY
vZSI3fFegzKdjGxY/r0IGlefXwfHseY7MJWQYRspDqcs1qTbgrc1BtnPey+K
VFK0H4YoNLGv7exU0b8tQ41fhAq96jIWYYEi60OIQbpkF3hV/yhkhJF+vNlU
n7Tb8nM81Q4vPsvToaiYcNFFT+d2kYqcZSwG4LpGYI1NYktmVQ755ju+SzsW
WvyOtAkt3YQDwGOfl6ZhXjpGTz7jsg6YbT3f3lWYG8nTtVpIBrLBym+8F2mb
V8DrxiUbMsVaQ0QoKwWvfWwEtf20l363l+PNxINJK6D22CmV2fbiwu9ycNe6
EtUYdFZ5fKYD1h9xRb4/ImelQnGVD1dc+LOLx61FwrcshVN1oigYZ+2nPj22
kIBP+BypSTJY5zTFuv9ZzMLdJn/U14XXBtqi0iMKylwTHd2z2Ilc5pUwfiHh
UFUVta9ED/vYz5HmSTZMgJkxKSWqIl7SW2BLHZh8Na65UQAYMeFhSH9yiFjr
D/2+PuD3pe+MwuukS+8LA5qApF1xnNe1xCrRV/+nHr58x68oeXzjV4oDByf7
sB5y1pSNzAIUF3bx8mdQymdJFIVEMBVipRTbp9yHonzBsyBwsKK+0XPL4OC9
Gg1tWsVIkt/EXTsNU35Bu37cdETs6BnnmHKbh9d7tVOd8dU/UQurcNHWYYbK
Wv09sPVjVEqaCdzimD279+yPRrNPbz9sgNMGpiG0BwFq0PXXgG4OhVbsDtw+
AJ4z1OB7g1qFc6RrIPUkbsGTu5VRORM9w5CpFwZdj/vdC7yxi0aucAU1Xobt
8/Icg6nzpeY8u5LOpWGiYy8Gsk57rH+Xg5ddXMJuYkOTU1VwELagGviIlz7m
K2xk0E3UBX+xG41sN3fXw+rJLiG9rn4dtHyMnesJhScBO8iNxrvXKh7O9hSl
jMunKYhoS4wqWUOUKR+BYtX4MNG3jkTWZNBskLAWSfSJnPGsNyLVTyuKyrUN
PyNaE8uPoKSTiuVofs3QlBwI6sEICfp7rhVKz74u6MN6YM0UAZsj4CTrgfq8
LcWcLEKe+BMCqIMR6S2Cy0E7Dwun+YN1PaK3dZEYHw4n7NOsTyWNNChB+C/X
34W5dP6BOWxbjv9EQpS29YTlzJSqoNFwthwe8NB1GgGnX5iLsDWAv6s0UyNC
4x/2MgvuGjzZInyl1/x5iukwX/m0xoKtWIFAzaXA87upbUMH2SLUefoSNCx0
JavgQDv/tOuiIAOnmstPs7BDB1uLxmCp5RAaBEPxETwm3F+ix4w8/dxAXw0c
fgNHg492SDHHM1wxr8LPdMG74Ksox1XWOXC6K+f/wJt/Wwjr6/EfFfsDlI+T
BNJW6OOlpPO9UQC5o7ArMW3SO5kFz1jrJgFCDLIxh7J+xryO4Jds2cj8+rHg
zkE0xgY16rFZiVDWGHXiZGT3ZE8/UQaEIXWSwNk5FgtorIP6ug6u9zdcTqin
ypZXIUR771JqEldMPPzqPxvDEtbK071fSiQ2DCUbAJ8iYJrHZe/cFzuf6zn/
NIOtTknrQB9hKlQl1+Sf2f7eG7+xAljGc+J+bFDKX6pXehLW85pyPSDadOkV
t7ANoHQMYoQCzG4uwB3cPuWiwndeM8RfWVYC79i8RlyIAu85P21ZZdL+EBWB
Dn2aRQEOCwLivsQlkybwocIkYWCcR1BPK5OsNPvt6ivRKF5YJcOOB5yYbphI
hQMJcAu04Cdd4zXPwaxJv8zSwvwIx6OVkNFSHMYFwisfRW4emx99THMOYcOo
mWdIkzXonzp8e0AvJr0BwjPR3KK3hcU7H1gkJR7h+h3+Zhq+sSB9ylpj/OR6
4KGnc2FUGRF8yg8l/C1nuaaOY1ZafWoB3yWl8NbEV7L7G2fEUdTgY5sbpDbP
naDQrsC7h1Y8RmFd7BU1u6O8UwtXy6ned5EJUw+AHouqIl+4apqzGT/vTyL5
Z4YzAFJXxBUh0v7ritOvV0QYRCaXLSqBhTVgH4L/t8jTEadyLzbFgBkVa+SN
BtqbyKw6nGHB4vGvIx/T2p3hp/5H248FhtpLSLUSrpTDm7/VpOTzx1H7I7T4
ZDPxYdE1FvpOxCowf+dw8MAYbT/95RrFRmRO80ZIGN8TFCq2pimlqa48jen7
Gur2hyfKfnyTLpLkIBDBDK6MlRMEg8nZEFS3kfODWnxR4urkf68+msI88roU
w4tFIzJQSxfj/FYUe3hyHiRfMgOi0PnoXMg1fm/1g1IRqt5Hss3b1B/vq2V7
5M65DKxP2venwsUklCgRCw3uRKVq2Hu+HISpbCOfdNJH4+WzZB7MhURjFfHh
8wyXecrB7mCSFkf9KashOnk2etiDCrPmujFUoyZdmLLr+GIvQpfpOrAr5qIV
dfRvux+Q9S5Msat9Etp07kBej+tzu9t0dtufJrRT0U3SoZlWiW8uoQr7CVvW
Qu187V1mzeO4GbtJhx5Auc8z6OusYsx7wlnuhzmWHsbXq4IjCZ014xWz1218
R0Z+VMGc77cD2dZrIqI73sexU/EoJtf8nbdPThX19heQA79Fl/E06M6gh/mf
xu59xoF4+PiAqUU1oECaLz8BPl1viXMlgppCYvJtWgOJP/YlyL6vwXGG42IA
38BKf0sNPFFPoqQ3pVrYMst96iKQPmk5KdlLyt5gzUI7oPvWdLM3cl3EJIf2
o2Fx/zKd1geLUcy5efvo38rhsIO5xtNKIlDrzmc2A8W9Mi6upRXzL4pWrwIc
cNB3nd+YNiGLZuYh5yLtfgQEVe/sEfzMrvTyQ+8opV3ZC0dnC1xt60Fb32aS
WfxyTmW4oMtZD/PGDDRIvExKXIPMsAOlEonokHe9JriBtHxFrF5152eM1qqM
YV2BJeM5/yd0rrsmpG9AovkoIwDGfmu+XQN3KWudz+umEmyrbVvWIDGGEQ88
tDGeXmG42U7cW2ryOKJbme3OuXQ4zzpD0+Yj0bxC2C7sroFzmRJXajBhhAfM
xxdyfivS9RXNtTPXZT5l2SmXu8ChJGH9ZLcqJSvKMZHxDGdW1COflRb7HTdf
6OPqeedGrHfzUaNY9UENnI/UKIdrMbVkVrv8MhjHpEvzNFO/KGXqj/1sXm6f
UmAsa4fQ/tShNFTiAPjOgtJkq3iOjjW3FjCyFw/9qgbqkLjLxze+4SXTaAn9
XPcnLJOkKaRJpJ+kR2XSwQMS7BD/nsIvAVFmimUW05SIw5NW9QmFLVAtqeOw
apGnATjVl66PtxnYP/K2JIz2OopkV8pI06OTD65EUTGweVd3BweIy4tiz8bm
NzdtzFCqYBJXrDoemmPyJJ0ascQ8W1hmy5QcxJeIHzLZbqw9j/QgxGe7nPAJ
NRvRuU5gkq0/7ytY0bFr+NcuuZk+Sfl/dNHFYJvWTmui+xQJCtDAm5lQb+0y
yieQ1OuX8n56hHJtnb5OiQqP5kLYAXIlJFZ2XKfAY7uro+JZGhnMhI+nBy6/
vNO2ZAzoEZgjnSIm6Z1h627jdTdiYoXLESeFiD8UP6Oen9J0cLJUceOQLN67
JHe8ds+EQikogr6tD6eDHsP2i2Lfw6M5cDTue+dZ01Om/aF6Wx797WRm9ciJ
rwUYe89idwj6wcpkOETWjjtby5WSDynoBCxrBOCNgKYkHjFfgH8mQ503QN0+
Tmdoecu0AmdUjxQReI4N8zhayrBOckjqv66nm/QpZ5m7KrOanrL6fDOGA4Uo
vP3fFEBWIuQBCnyM577cQtLsJoeFp3LbvKeNvgpR3VddFzyE8EekZAUhwJLI
JrcDzZvUjQYHQLr9Y2jn/Uu4a8+4oY0Higar9oDtvMhcGmbb48pElC5qxiVW
36eUD5ITucjNYepv6uWZGPuPCLlYjmkJdFlQMWswyeLruOsIksqACPV5pAoG
lXJJY8+2ex4Q6wduE8No7l8QoaSPo4eznwm46GxH0GmVT46F5/qRSyGHlRNQ
POqrtmECRV6v+NGYCWFC9EbRpjhPMGEcqp4B026dJNC7zGXU5kRPtP0BseaO
EH45xpje0o32q8NPKo+hcuvG5CsmgMNo17AfRsfHEoeo7gu2Xs4vAWzL3BbU
kSp7EALwtKtniUlKleN4iuXWF4KuPcFxgoSG7mUhdT26k8a1CGw+EfKxsRZ9
ZbUJhivsCBQmOyXndffSORtVxUkRGzvMk4zmFc1Q4QgG1msWnNr/Z57PkxkI
7cZPv/Ifp9fT51rFnY4ImE5hYznL7SljWEPgWw7T0oZ2/x7GszdqCpQojyCg
FLC7MUTf9EsSpcZcEwz0RxurjFa0Xu0RgbEo4alltzbue4R6HQlV/nin2+bX
5Lunw8MX2DUJ3y+l7hscJPvgmzeTAZF2Dre/4tdrZ/4pDBeftYZ3b4Bw5el1
biwepvk2E1MTnrMWMKwhF4Xyrtlbqm93rV+emxXm9se1w9b5tAwOHPRYgh8k
65JaiP5dtLuHU0cgG0kx+tZXeXxx7S4XV7tPts1HNctTnsnu/qgiXRPg/b8e
QEj/Lthpmq8NrF9Z3fxwZlWKL/7Xf401OwqtZLgJJYNjLvtZMO5zVPILNsg2
8bbOSlKem0oEwRve22uYE3UlyQziAqBLYX4RM4/O4A/28F2x5NzMnvR4hMKG
ipOMjnG69IcJihLrFBquDnR7cGFukB3oZH7uaMfj+I6dww7BnXK0zwMMoEOZ
qjZUSPr9QUWj+l1NUw0MJSOFEryhCsBXQUO0nDSKpkqvW1cO08/8ADGYmZau
id7NV+r0xq4KBkVjSwoqIa5MAXEM8iS0bBh9vczXTLq6zCawVM/aMyTI27Jd
hCjM3WqXOJqIGMXv8mGScdSiTKZWirgoqUHezQNucH/JXOyjbfqwnuZ0Uv5b
4yleEFBw7NiNioG+LXuSHVzn4ZrQShWuQnncVWV44Luu4mEOahTdB3vWZ45+
bKgYfyBplW5t0kAFDh/sDpUL8Qmdtvm+3V0iwQ/v2wY8Qy2L4XKnVBgKrQrQ
shseCggm/qPuNkA3vjVFXgkcgvdqyCvCyBURKO++Lk0Wv0Duq0iJNLW4mraF
P+DGRc+CRr5eh6DzOpiVxqbCBukmCsN8XcbJaFSzKCZeuPw+e+KIu6xfVtLu
gZ8/GfhbuzQZlyo/dADjxsQ3XBOvGJHWWIAdV5x9J5lmkEjzmPbg12gl87BK
zMBCfUYkn60stHoZofBWlp/5fKOj0dMYCJZoKfh2hUYwTFcGg9A1Ixp2UKjA
iqjtZxrbgzcMG3kdAhtY03flNlmwpgIXABJawdsSx7VMYtIjX8M1hyJM9yBG
7wJi0zVtKO3y4Jm9naRPrjUQLPjXadhYNHanJDv5xqSkR48Bb0/plVc0Euzq
EAKjzFpjrfd5mx/fZ39Nd70vI46fiiDozR4oMUt61xqsmnynQXRPor1fPfow
ZeCUZvGnz4v0tWphElzspaMwEuTEoT8YpL63/6GTl29ZQeS2u2tP7mzEMrQy
9fg7rN1YqNfEetcPS/t9gOLIuZ5+zuklFLUdvE3MRJjsmSLPFa0Z8k0nG1dD
t0zwTa7tkbjqhdHFLhGwGVMDsgSYjJo16y25rywRxfULCVmy5iwEa127n2LQ
JLMa6poiTgnzkQDxijT8/yEhPqjTIc1tGxF4ZjH8rZ0eSa79zW0BDLAxTNBF
3NAVuVVobZi2x1XelgNGPioAH/1Z+82YAKKXgA3fcfVYbjNiD/xD32cIKm8J
USVjQF/X3Ki0Cg65kDYFUROm1DpI0uEoFRtrzF4jZpcbq9JGqfrQiTet0H5y
7vl+fLqy5b6j8fpAwQx5wob38MtDk2vB08jBam9H7miwaHmsQlN/f5kKUqPU
zlYG5x2o57yeaHNc9jY8w12BMN7YPyxIdyVaPZ7KqpTHXeENSfyFpQ+4TOQI
YAVWup62jRHIbRQyYNGdTodUVPlTtivTWP9InKXqzVa9nNHSCUHj+5yDIKl6
Z4mM+G1iVOXLnqCiBDSYibr/f5VYywbfmZV1/+BT82p9M80TKqW1veGzUMsE
cSWH64s5uy+WvwlXNtAPXfke9CvkecHMhBvYgobIwZOBmNkgIq/US8lYBvkq
9dw2GH0cgY5ZKDNQtB1OyHBEV4yDL9SGK8ARUM4BL4eoPPBjd4CoRWbLJxCE
AaKWYek0+OnNK7drg5OHlhfAvrfxpyNJUOvnjnFMVjS+Kwa18P/W5sBIYr3v
9i53PXc12yuSalC4g4fsnL4OCOH3HEgF/KmYmoB0+D4E76MUtg36dYlCDl9c
M/+rSsb9jVn2i4ANDV6CIa88ts9DHMwYSW2nSu/u7PISrU5d50Fx4hoN95bU
UiQhv++DP9NNU05rI+63hsFkLCoCieR6y6G0wUzbXb1/wjiJT9h9rqQuqFHM
LZcqDRasHyLrAakZCA/DIinz7qIFefx1TmhrCXhlmFbqy3iPXWV8s+3oqzDb
dHAURiarnZ8JNy1MpEteznYYNNf4EBZMx18gR3klD9WjsN4ymhAjjTdSQyBl
PffWyQ5azl/pCHDfYNhm/pknD865Fx1D4I4tu4k8Po3Gl6LxdtryX/tsoZUp
6wOTMfQ1V+NigRVYdK/l5N3VzgisdULHNoj6ybAopx9ppZVRHS+BtmquowYO
MJYOUlchee+27AcIxrL6FqouYcJRuWTXa40B5jX8VSkpzCQcO+zH+TyedRkR
P5t7hYwJoVNIZIf3mFr/XrnTbd86x1OSXJ77f4xK0jPZhtHEX1u3y3Zk6z5n
gTqjDLWPOlkb/E2UI+MsaenbDoHxy7e7WuQ6DQFWP/TpuWhrbAzqbI0FCeer
hVGcFLxvD2EeraUYQoZgmj/RhbbG/xFMA94A6R2S0DZCddWJncYi4qx9der+
4qXz/7/cea28TfOqpUZXvLXwYhMGZ4GLCS01riNqwrVUqlV8Udflq3bTFor/
PFgZjKEHsKlz7lqmKAReiLggg9Hl5pBc0TWfe4lrITGsVWnBbhKRz5CwQlnp
cqn6cp4BtJ3BNpBk1CHpzM09wcQpeXRsk8U8De3K+N4WNU5Mz0bkuKMNdSw6
qeyWSnuUBQPVQrY7eg9Z34393jzYFlefaFSn7o2BXn25VAUHtR6knaOLbNXk
BQrR0aa0jTzgiyKwgw7IY83/WpDLuxqFWqXG5xgHzuiqoJWaLACCBsW1AUYa
G/rSHJsBSbTMfS+WcwaxZqNps+s9kANq7mzwsqAum+hU/HFXI7USqIYOd0rZ
Lkx6IktrNL8hFYtT/X1XVLuH3FKGSXDkzMMAR+1KQ6m3V5wRd1HIyM1QSkc5
i44o7fkk4GpGEEQ77X+e4LKkAz6wamZGQTb/vQC58G8uOnglSMZBSfpfMcUJ
2PN2cGTggmbHzaoYoQCeO2posQA+DBwBHI0BFIJvcnuUR3UzwTK7WERwDa9+
7m7EdSD6xH2jcARvM5l9k4YN7kUlqVjNIHBDG2FYPqZWb4bjjPnBw11eC99Q
ypnHrLNou8MrQs03L81dxjzhdldTl1qP+VLOs92pRJuRy0V8mnSIvFmbBB6w
ykRj9/FObsBot/DfXGaTBf5n8sjdLhA9+DBxUMsiAXRjpwkD7RvVEZzD7UPf
F848BlFP1/FWlWnPibvqt1DQIml38C1+nqFDZ5yCCwp0CEcVjWT7Mit/PrG0
S9FFTZvG8sq/IrF/Ce0a/nkQa/Cg7xzXiS6Ug/jf9lajlQUA13qmcsLbxwx4
deu+0p/idiIk+yolPll/r8ud8eJSsqTHdHD9XJ+f8oK+ir7ZACn1bEOs1taa
Con4M9hPY2BSSki5tyYQxwXTf2NtZiUXUKo3lnhVmVfzGt7/27Q1pWJiCEnz
MIrxqpQc5PXMLZzgg4o8+4EnaBhvPH8kC5ML3ap2AoiIjrWVdRsxpY0QnhM1
XqIyxab0sym6LE5wprAGafpSreHew2f627Q+PnxgVsxj2T4Q3/kq0PhKuIqV
y5QTUu+6PRfnxKPxOe6oNIYUz04hWH7CpArrAIohSFqdthbxUBAWblaLkNM1
tmkRI5mlBo/g4qL1SMVZWkf04xG/uY4dZetwGdVL2yjODeU/g35uw9NwrCNo
YEQ0964bIDb6ftvcZzhyx/fu/C82LB1vwGQDopapjcWsytx5ADBucDR+WON7
toxJ0fu/jx1mzrxwzZpovPVBt4+vEBqzeawQudYZedFs9Sk83vs3tY8MqSJO
SOBhLuwSDl5pTIx1KuNjZIF0CqJ6oAftGATq2XmGDmetywfeCHKaa1EC0K9U
DC9SCkIpNbWUsJjtqWT4k1UeAbUbwPII0r9uIbfEMJrP9Qy3Ngbe4pTi4PTI
Y5/wzUbizcBDFt7veCoZvQ1hwmSLKwiflSsVNyyGFBQnMQskfmpJbXKm3AVx
5I9jWeALAcblBGB8wuNb0HgF017hH9e0yLywUJ4E9orcpnJrf8cNCGHGNXtX
01fgyUlUSPidHx0QUo3AepecAdgTNGEjtPorMI8qgGzLZ/ZK6BV94Ib12YK2
2lFelR7kyzTa6Ip4+ta6fiTNt7L4WRuZ4iRuOh4ZrSEij+SfNzDMYGfR1MBT
fi4aa0SDyRRFWhb+dnGF53wYyaDUrMmW3sMIymOERZfCxLKK5k/8vCREbttr
IeUoo2LfwZeYABNCJfWmysZDFhRYbx3m78JkTWvdGOkRwRSFTPcBs24xYS6u
9Gc36SMVLZCOwhYqgImgG4tYQBlwsCTkSJj/Vq2uzH6FcIJh1EG8B+qeVzZV
gFeT3nP91OHM/71HmgGFd82Ryuzc6W0Xvfw9hA9Nb7MxUYe3RJlUtFXp7s0d
dEgQMsWxTkh5lW4Cw3zSBtgPrYoq+nfWmx0CV/p2dfLqNJnMijChllaRKFnH
8W2j3ZefkATiQHTVDhokFgKMJcbvdhsEXd+4EBxGKHQz1VT5CMRn9oh83dcn
TyQzDt+1UzOnWJZHB9ioWSS+rFMEilx0L6qVk6y1K+BpWfJnnEGwnStEmGMZ
h3TyQFBvt+YywHhCujpIPbPFKE9AU3CL2BhJ4MXsJe9X02Aaq0H6LWcnJYcw
uNqowKh8U21Bp5WuWLiQOI46zKcM20dPpZnhzwScSB6SOJf2+tQ4np0acur9
PXvTW6x5ld2DwU3Q4Q43i4fmsat4E8lvXFDsQtxRtNleAPPdPCzi2b2mDEhi
ROSMICmcJVgc2bcOQ+QJj82ABjXDfMctGTb5Fb+lL4yr/Ng4Huk71t/lEaWs
Gb4fPj/NcqHIc2Btv9lmdktxeyjdyd6Lrdgp4cm1uLHaDFCBjIVrR4vOpgXq
Ic2Sd8ugidAP96sWOEPVH4pWERShU3ljTieefqwRYVKI4DjuZp6LZ+YtWVXE
pjh49pzdOUWMhiqhcyeBr42kwLc/g9g1Irr2+tXZCwSJpnTAb2f1tCl89obi
e5tkA8awX5IAn/X00DpGP2zDf96hGqmbSV4cnGGyr8XCjBUPr2inQUsZgs4D
2u736wBHa3VCDpuBERGvueXKMOQzjavfeH3S9aZ5b+HPmnyM/xX4Zb5qXG5g
NHMo5AS8cDkKOOfkBeMd8/IZquELU9u0DcQPX1RZB9Bk3e8cI6LK9R/Tgzap
TNfcUGLHsu72QrY3ws2/2bCvt/5kmHIJV9ek0xUpEDrI2gIQoRCWhkrBqkdn
J7bReuZnOgpvH/Uh6or2Poh351LgrNko14cs7jnJjSjpqAPDgyk6Qa42r0m9
8JRw8hCcte0WtIlxUDUiqdnqkBT6QBmsENz5gzF/vGzwR76oVjgxzmUHzKFD
VmmYjMMQWHhpGoJ4KgZjA90K/obA46RN8JDHaXk9w88QQLbA/uqG1picyGWQ
Cdhk+aAwbY4j1NRfuAZFBzHzxtPYX8Pkbe+0NK29V8v3pW33cQ+l5POe6XG/
aYD9SjBUZukhyYOLjMECVeXcijpJbC0k+xXK8gRtz2U+05DFN89e9RwqbM5E
xXaJc3WC7W6EnL2NjQbZrMfWIgjcrWihUmuqQU+QBZT543TEQfevbLJxw53L
8hHBRhyggvL5lTYNuRImViVWVlRlGy24QwtInYV6/yUfvLbs2pSEMdT5+d1j
WDvuOon7UyQ2ZlQ0PqPZ4CBSW2CDPWW9/qRE3Bd5VVNEwM4bP+koGVpFrQbn
XHhglinsvsOxtS0krQsz59y0yXeOTDu9d5R9e2pmWz1sNHRu5YqyRWBvddjT
FZaQFsfTlVqDph4r4gGMqJ177eVjRvoonOSAFVSg4ZCezHUX7GvGQbXa0yhR
jSqaI1Ck1ChFP/LgbpMxk0SLLTcffrzECHFLczPSBvPG2lwNZXv72BdVSoDX
v1C+ovzm3U5Ek+RniKV+C82o9p8YpkOi28PnkPsMBqwt75bFlz5K3kpjaCrB
k9j/Z6H+3jdvUamTL7qaeugwg2F+x1aoeTAyT6GCbAzncyt66OlEEWrLvrPL
aSQ2tHVzTEpdDpJMY0po9tNK2J8nqnLu1x2EX0tnFe32uU449vIsYM1hcAIc
HmpnAkAb8bUFlwjS+kCqJ0RnkE2eq8ZBKUMIT4eF+tch7ktVtLBjfAzFURWC
2Qvoo2uAZjYw3TUHIo743m7uK1Dc+bbTC5ALkXD4lww7roRLyVUu7LR1iDXx
EZvtnbUV33reY/NoAbADptncgjw67x2RxyIoootHqP6XHSy+TUI9wKkYnnPP
uzl1fksTeqGYqy3MQVwNSYt/5p5SO40EOFjk4gG7Sxca9boFzjr74u9C06mK
GkyoM/7j1pdS/hh6D18BazF88BD0dayssaUaZIdgEZB67kFeqweQ4lgZC7Yx
eptTLQxXyL13K5oHOLJ+elkxlnB9B5GnEHikElBvtQyRenn+IdShNJxYNdKe
3lOJZ1jkvHsbLQSYC8bugZmYKpVm56oOSf41gcJJUmiGoS1mN0meZ49OODbo
oTfX3zWpwlJtL7cUSJmmshFLjVw6aUjd87E3bQzBkSH2QYNLma2839iXvLdM
DftfZwvATzjDM7sct+dHLSRmZtpsx7UN9xaCaX2TXipilIicqQpECHMDCPF9
ln3DcmjBO72VeyzeafEAvYmKfboPaUzfqwPnwMi/BXcbssDxDWVofwkkZEWu
XEYrNJdQtW7C2fzsaqxc6BaqslO03Bdo6PM2JNQ+pVO6MEjCJY33b0oEzE2X
BWBuix+rdplG3toxuQsLDdmwZCGTdb3kSUrzVWGIGrWVqXlQ+13YHDrye7wH
nBYLqnPaJFXUHLerhE9PnKnYTOkPtrR7jY7QHkgrQBlUCIq8QyhTCY+BBSye
pB8dMKNEyvKakskdsim7iSQq6e+Lh3ocXiDyMy4RVIir4pC9AZJlrjGiTVop
9USWlC8oUZkwti8COSIicIoVXMD3D5tkOeU4wpijldsubLJG6d0Lr9lfsinm
dYnjcV7Lp6N982cpFOUZsaX04HZGa3zo+s6IIuOPwmyh+KVnbuWsqelKEkdQ
FGEgMEP9iMjkT3otIfNeRVxPrh1sqMYi7xlQ6fvYfyqpYyHLDDIthxJccA9k
ry8r8K8keOAYY3fppjyU1jasF4SDyHah8pUz9U5jbXOCnTXjZgWO731lVU0c
f4LONB+qRlM0e2NCAFC/z/iZ44MT1JC39UY6UqvJMzbC12QrkPSjf8vKmtXi
4k5Tns7vcEWa/x13xQVvR3NnP/IPEiQR0EFl/F/xz/hq5XCDWX7tnIDC6xfN
8opVAhxfHaIy66l2mypjt64HJyFPr2gJIBdagN+wQumcrXn75Xwopr/PghXD
85NSQ9Hax6DMi06R4qRUCmRpTMjTX4GTMT9EJ6mY89GbK8Rs6HgSEQ9cSnTN
mY4/wQdsrZwIxAW1uVsu6LNxg/Y8NslB2SBUnz9mdE+pkmbSReVTJO8PGHTz
6Z0GDNb3b/riB2lsFkkksL7A4rvVENZ2KAN3MLckf3WIwJUpuOm+ds6YO1hS
vsoqKX22MB5GSeF57EdlNwXEazpUPFD0IQSJepYp8le2HgYrcfc51lzbbbM5
L0feVWudi1kEYEkp8TtFga6D1s3lAmp8H38y+as24hmRKYn6qt3TvLzkdMjX
tLkchTE9L/zeMS3Byq8ad/lvwS8xhmvT4/n/tkjmFFUfBQSZAMW+iygzwGp+
W2GlVuVVKviNZNO5tixlLyTFAmXxIiqkFCB8VRhyc1XUMvGKVnX5AvgW7beh
XCRgH9g9bE2viOoEw5qAyM/o/qNPDFPNbRNQM9lEbjFiUlitgaMR71JAV9BP
FQqX6hfAxKpLICigB9jycys8KdOYC0rBe4fSX03Z/85MmKxc1NG6lPlWR/bt
8RDDmLElULunobGG36z4Gn6Qvb8M2noEIEnjXY4gXGQhBxZpKPW1oTSN5lBi
yh9uHy/qJ3hHnKc4BEb/qvsNVmiKAeQNhwXUSKdclF+MmQSUGyRDqpyMlUfY
cr1zvMzkJsMLToaIJZUrY/jMhL3mY0nc6TozRyadrwzMXgDNa1tNpFEZnabp
zSQf+ju2hgUAHLeUh0iLlHGp8z3WxOZtCFr2VTEFZHwxMI/jQPjq6yDVjTrt
j32+31OwJB+p/vCAmRsLoEMH9Lx9TALjRtxnWVZYZ1Q3++qbimBw1aJnw/io
WOpce96sR5CSFo9AXNQmj7/KQ95muR/eaWeTdMdhcv8PLIzMkAemhEXio6Em
ne5Sv81gXfn/kfhCMFtqsqoTajQYWTnn/8nVDTPW/PgjXUAtI5WXn2Td+Mtz
M1cejV3oItYEQmzqAF5Ej5Bl1GK70fEJITVSbwbSBu8oh2IqKJ6utzNZPs0H
xm+peyDFLrGpJbDcycoPJV6UNQvASDECPyPxR/bXp0x4/JOg690+yqZqwVK5
topow4ILQaOco0Wj6CmPOCgGckZdDtq9Bw733quqExQfPLmCb4Fffh2O2B1U
NhHlQ5gOImF/BKi5Iz1rvccRmk5hRBAkozY216yTPaMQGFt4eNhCxnvaCnOA
lZV0qvi9i9AWx12+CBAqT/XSpUzoyquR8L0/gn0qwy0Ml3y/onfz2Xrc5hqj
qTuW2ClgNMc+bt83aFHGYyMlv2dHfjFh3bccZNLEwZdE591OSz8x4TnJ3Hv/
VcAEy0I3SjT96wpDO7DKwNiExbNiyDZgiUMRpbhGRIYRLPG0W6MU95ctBZvA
hi7+V2i+PBIUNVMeqsK56vw5LrEqquP+Sgs950WYWheEJOWDf/VsGxqvM4Mo
f746GpEtQ1yrNanNf/IJVHERhAZ5tb3W3YgcB//RbmYPiOCZaLN/oEmOyvmK
rpXU4FDmr91oUCgR8Gi7YL8vccG+XLQX+ES0HSAvyX+snaP6u0mTXYWdA3O7
q6Z8zXejPV/8VK6A6qiM744bJZi/PKe7vr9I+uLIE1CTa/FsloXgI/R9l7Zc
3q9fsrh6CyVsshO9cUBzTBcV/TSR/z+pvfiVH4EkVrjW9FzDlTZs4RQZwvkS
2KO9iVNyJPPD/MenyIQfb2v8Da3kwX4MdPgySvoMFDJ1RFENErMba84ZjLmR
X+86WxA572zIir54cMftpgsskmsdPIOD77HLzGy3gBrDIgtZZHTN0zS6tjwm
A7V7LEmCuAu6cZLXU2rfRCjlet1TPpWMemeTuu6UtcWvZKlhVS1WmijV5o1x
S0n27j3GW5X5jynuNTN9LJYtUiiUV7M/e7aLqQaK4xprvvmUmigWQsBzwzC9
7RVZL2L17dksvvEAw9dnC/jdIc2LhRKd9k8ckXfxx3CLQbQFO8UO4ikSQUHP
hTypN3VpXlH/m8zG3IWifcPIOPQErqfB+E+uMGp3lhV5XFH/P7pGV127Y2qz
owQ/6umzBNsDDedY2O0YZRBJjHh3tp7QZFaYzwdDoEmfjF4LC6ijAcAjaqTK
0GMRmGfHP2tk+nhgS/VX3J01g9BohHMCyDrwYrdZNqhIYfMb9Dv+CtuOpyUp
pdpgzmh//x/A+vXSysNefapkEyPmdYheTKm5PUJ2Ej5XtgYcw7EvXTAa5DOE
+lrEEDql2CMFqN3w4TaKLIY9ry3vqKt6gRh7CCfW09kGfwaJGJNTD+gsmb9g
fqPkCyT12Wf8TqZfeE3ejbzUD/ol/AIdLNpHFCEyD91i9awhQNy1D3EKAZC7
FwQjTHOC0IJD253/YwzIB8Dz1jrw4vTPqhbNo8UBj67PsgiWzljPkdURb9Ut
0SQtk0ZGJc5aQ0uG7TqoA8vswZuRZhvuGFhffYW1iHJwVIVpAGtPs6C/3por
0k9f7CgVzfqqk3NaT2FZaHca/rruBZWCXRuQRy1F75EDA/3iQNvF2imoT0Wq
A9p8OtHR5yaYyPKY5d5evu0LNnv+t2keSzA2EY/5hk7KuO17pKj901qxPYzU
fnX+NcVaxJvTmCDnA4G+LOmUmJuUA/cVFp1W0ijlByF2pCLEcMYSKRyCLIz3
LhRskRxsulZlfGogMRil69Sw6C3zq/unGODL5PSoO7r5ZXbh0mc/ifnBzmvF
3470IbvlDkyEL4V2Pmu5562iaaLuY9RqxUnIv1J25oFnrmtTSI77lK+A6YAG
xi+T5JOsvrSmEkAMcDnqJxWJnZ1IUhYhKhJuEbNwErXIF1Z3rBdBEQsBrLQf
640ck6u8E05Yf1fYAcSiwbuyfqA9LZBWUtcPyglTfKbH113icjMSL1GNYldx
xLBGzexdFuszVKuEPhPHBi6Xz8mvV+zbIi1aHHU/ES6tTDUVCrwhaedp/QQH
ka/w8WIVFCTRi0JiHFowzcoBEEeIHbP/A9hi4+7fLDjAXBYxJyNl93DAYoWd
2MrfOtjeVkd9xnl3/hPJr7U7gVK1hrpB/RaYjkf5sO7qD6MwWezdduU5ak4K
kUiBsv3UHUaIfgpigUPWhFN8RvB6vKH8zsX5P1hdfuepsg30unDoJ2MjVLYg
JY8gVQ5wbs6Duz5KfZf4LIGmNCoAC49UrV/MIwfLfdpvcjeoIWCf26+8FKiw
2NzzYZwI9QOp++mWJGh9vwiCN1mIZn/BcOhFqOhbiS1dwmejh3AR+T4Tijo3
yC6fmRx/6fi9jtV3avuuzZtFw2gPKpmYoFR4Z4Wu8M6jlj8oc+TsGYBbudWR
L1e49hagBNRhQbpJEvhw//loYkI7I74O+DgtjeqfFyud6tH/0xE6py+CfwVj
LyJ8rt+4dD6x08V+ijvlf/d2i4zEOavnanDnxqxriaoAQnvW6WbVv1u9B0vc
RmQTP5bcOmH555DyPZ0kerbCt0uH9wZd1FZ1oRof1BTHZ4lSLoSF+EJrt1p9
OA5uoworrkLqnrp0j/twFug8vzGgOKxSWn5+PERzB26uXJRVfxhpx6fbo2yu
Uf8Bvrug7/8g/n8OWJTOo7Bo8IZF5i8OjmZdYvpKjzd17GxKHvgGBYurM5TU
hR4AH/X4MLeq8vwlRR6C9wJUUKjxNcgLKD8mNsS3MEZW1N16/a6GtsnAsQkY
WdsND3aDHB33zzUcCvGdKtpLfUmEGZGzQC4jyEEDik67GBbDVvugyquwzTbE
/fN33C4Fug2fFsGL2+pf5LZQdVRSYn/WnSI2LJdYDVfHoR82nOLICHzL3Hzh
OTB1yF9bNLjKSosqqQk8GsS7G/rHPM7qindoTT1X6ViO52O97Jg2SCVjdn3e
WBC0C2oeOqJ1l5srh3fJvh6B1QgPDpqisSTCsPVqOUQu6m/+bORgnWybp/75
6HXj+p7+QG6FNLHHDTBiTlf0NqF+dAmZsKKAT0EFON/lrvm8D9AQfBDK3DM9
9KApZn9aKxfKaRO5CmykxmonjaKd9UURQWq6IM9UozCcmnOqycDRrXLzOjae
hw2F7cwf8wBcRbw8il+Yjwdby1OV2frumWmUf1c2TAJ7TOUQ/pLT91JNgxZW
lK1AUFBXOP7rfN5mo1lBTX3ep0dSd0XOE8aZLmZnCyxStkWYwLE+gmOh77+J
sloBoRhCeBDmIDh1mbqbtksUgKcr6/eU7+bz7/9GizaqWNJ03H8yh1I3B7aU
Zkb5RUZTCUuEjxubd0bsblIQNthNaNiAmb0N+IK1/XZ5nteMUnqH8BxvjNxh
Bxj5Vly423MbDhtdJLXsex5vU7Aloor+0vWM0uxAKoEihA2LvxK81EMY66rG
NpqgYt7q3PB63OQdf0U5RAEFABe50vKOPdhpDVQQvXQ1gHQk3CGJGG9MRdpu
R0ywWS9O/AtJuUbrbq8/ZA2EkZFZ6enIfPTVvLfRHxpNBenXWnB+iZpMotJv
dJ/m1PMp8Te/WY91U6vRSzf6vH04Qb4h9Nq0s5cWJPUuZ7hrtEF5ui2tPgHI
QKZmZ8HN+FJKJ2EMh+MZFrgZTu8w/qdN9RrM0UX0/RkF3H4WdMh2f72zZ3N1
xzm9XobnnODmgZoQcBK4cQn+QHqwmqTlLq2UFVt0tBWsH75A69cR1cR5vdW2
zezroiFiXbzuA1yYkVgBaLXDGXJph85Cyk4kKnmrE+6RhU1FylOg0o/mKcKr
YwXj5YrMG+0lAXI3QI0yzI4GfAoqsGi9y0Dz57UuUDNmCGULNwsvpjYCpMji
r64duAAyj2VfWnopMdVMzhXjiqJ2RtR+vtrRlsfY2QszOazM2U72XiQeZOsJ
Abpeal+OX7OHPtpKXuPBDRKFhzriGNEc+aczvO6fIPTyzfYJFv/adQOidksq
PzzlWIExucgq5mCGDBYL+GKpD9Grdun9hObAEHyxjGKW0nwMcrcoluO50jjV
4Tc9FRtfb6MUszINze8No0euZFWWsZNyMiyW5KaTBiDKGwk89qabgAxnw2Yw
SvwbuwbS0dacUWT8fU6rB4SNqlaW1oT5hB128XEN8R2OduAIwGarqKAZ3Z5j
ZlqVnvFK4ElRi0SIvKBPtKlpF7/eg1XLCEXb6v1s3nJPzCXUdyuA59diGqr2
dTnyW8uOLWqHYiN9/Ng79ZFtgm+Xe4xqXgWAt8WlHBkGrDSi11nt5jdCyzyV
pvWE9x5S369W4GZTbEdvijmswD1UYa8t9wnGgaaT4gc+BOUMhcxtP/HbTucV
vEzCF3GFZQHuBhnOX+nAIAVB1FTSF7gdp/ly8oepKkJEEzBMQoJaKfOt9fOY
Xm9sUnQt87rdo2tzht0Q0G+u5DiRr9do6zqPzQBEzMyu5Nc5NzRTwt8UcsNZ
C+exeCx/KGyALTigFlh/51203fKzLV4B+wsqonQMiOI8obaLb0AgHngNXvb7
sXmbZ+tkV2PwidfKi4n0pVJ3ssjnZ6EqaFIDIzTUwF46109XbIxdyHS8jIAd
czUqSB93XZd0LuYEbPHt739j0/RvTbLoFSocLRIBsS/GHwXYkUhapBuDcVjg
np2CeGPru7ekEVWH5poBRQ3OhH+wUTQFRTrZt5N4+H3OkJykgs69+tbVVdbG
u5CLJbzO/jV/f6872VlylzZlXu6Y7phhfThpsE1dymmMasw0GHxRn7iWwAbP
GSbBgM4gvgn9EQjngymM6zVkfZ/6cPJy+KDjZ76JmW8F2BBRfdob1N06u3+u
ry5XVFWhA2Nl9s3iVJrmxvn4P21beb5jvtYtpunmFgT/KV2HlUdDXAg32/5f
LO5PMxE5lyeFiLVmkZs7GC4VpCRY3y1nFG4tbJVfQ2GfCRtmTPKlugsydpQX
RXF4OG8FDZt/4+iAfGlla7dgxE/vn8JO/G209hq8JgipKi6AR2XLqlTe+ZiS
QkOsDuoDe7b3qkdPXcDDmirLqLm/7pKWOyVL2dRIUMaj8Gg7P2JminncC/LR
dhpXFPEumI94AYKoZY/tJYkWYY17ZMTY4TCKQBiqeIb3panwI+JXHBHcHDMh
lpiGxuXEI0LI3tRSuvf54kLvFaLqdOZIbRiW8gbCQUhBIJv8u47suFsNFN0l
nzBIdhf7ajehYao1E8e7hpMH5lJsCyIRQbYn9paxN2lmcpHiJzcUkJCkfpD1
gwQmvz2N2xfbloQpbZcYDfo2U285rbsu07ImaypTtRdVdiSjcMFXl2R1XorM
7gzBWd6WjhwAhuOaOxxiMugFrzCBZplDojuydOR/gfrhUp496C5gV3NFX/Vp
uSZ6ccI4a5HNmLsGQiRWscstdLEtnp76GmWccHZlcTbsR2Tj+wIUCn9q2CuP
lRmqHw/ZrmnqfJro8vg3ZZ+0oJ/ssmumimb8zkTK+iz0pxCIgn+zQm4lCLHx
LBlHhFqZiZcT0zW902+5EDkd417VbOpcVkgxbbwhLBTs5A1SQIY5jnM3KyEV
6Xr+NUeOsU/UepcFAlI+M2YeYlZf09ukP+TPXf9erYNEL3afq0r2fIhQrzEs
2wwPFzk0Mq0tDFw2+saB98Lv5JRuwdE5OVXO6gAbALyY/NPZNU+4MTJQfl7h
62p8PmE8s5J2M3nV9MxVb2LZ9GdcpH7Hsp+M0QaqT9kO754Pp6wHch5dBgKD
xtCIf1cD0EU1IEvqMawW+yJDuzssGTHZJzgVnHjKxPcdrsHdVVSDhODDekel
wI3UrEFUqlR2zmWPWhlV3UwDl8QtXSan7oQrPxA64Zuls2XyjJusUfcrMntp
L8HUYGyQR4RAT28272ucm3NLA3Kjpbq3InoMgXI4iRplyddc/ZoB8EtGgunQ
9gSbI4+dWvy6KQ7Z2RCBef7+ziWrPCBGNmxztzuivrJvEK5MnFm+uy7dWpz6
yeGbNeGrrkIC5y4IkDp6PFDLNfXbuZ3TZxVehHdudrICIBLMIKngnwup93Lu
VEfsk1OCzkkuemdIgK5gZ8mqKIAcO1lz3vTtTRMF2pRBqQJJOoT8YN8/TiDR
70Smh6gsyduwvlpjI9wyeHJujqm569U+5NbFKYwNewK0C1cO2j8ZkS4D7PfZ
ecLlraI1A1ubgr7n1+htSo46dCjvqhb6u86sLpFJuEhac7w61gvUi9BvPTO9
DlRlJn8f4dz2cxvlyZLyCVAwUEOh78vOL/3oUcGZ8XJT8f6LummJv1DyRiwq
P+ihKw7SNGqBGOXiTCWYHziHyWR192GX28N+l+UmqcorAJXz3LpAqkNHFK2m
5V/fCQiZeAwj69bmsqDWCdeeWNccpw6qp9SjAC0NinCDSqEAswugYGg4zh8f
RkQlcz8XWPjEeD9KIu6iGIIzhGywWF4qK5sEPMBDcQtZ+nFfkzdfLx1Xs5xp
PeIfSXeStHHz6DEueMn1GTottYVKPYqJWNT1epVr3bDabr9s89cZwtg6AQpZ
nAPzN2bCEPPE3DDD+WOL+FzOBHwN8kRxaodHGOLzRdF1mIsdaIXyvBaMb//7
difyZ23wskIQU9KKxU6M/hDVA/6C3nqf4wkReB753p/UEyEHrQXVtlhbVAkr
D2gYqPbEe1/6zszZ4AItLNbHspr8AZk+TcRDbUwcjMn+m1FQVys1eg4FU3mQ
LyWxNyNlIpQHvvqmY5XDHe88ASETS01YWaFpsLO8u2hhJmGRYBEpoZzKgSv3
fciqmaVC55bqTLolfN7HnwVoq+G3cslRbN365NCYGPB8/qtSDZiONBjbIo1D
F3Wlj17ONISTz69b71rpsLJkyfCnXfGAB7KHGU5F8+77lz7wEeNjN8XWCl8l
LzANe40MUFyl8GUnfsij3ywGu06qOp3N9qw2m6aTNo6GDqRO55P1CMwsnVFD
U9qM9NPK+oa93ZH1NVXnkCWsHKC5FHB05qrg20RfWouOs0c7d7C1z9A7T7Uz
xoLioQ9yO5fRHbPxTIZVkE48VmYDaGOpMTcDBzMhllbRSVbFcvTLpVfV745v
xkl93xNgp1/83249G0xmzOWiytl77wP/xYyItaZoKU4J5yLDpapIFbNThE5r
Dv74yYpKAD3UBl+3xUNXaLmO53Yyw5+Jsgy13bbYKlAKzh3vS0XBOoQoaFUs
ij5Tmcnbkcw4Z/pvwNMheIvN/GcBB5Sghoh9iOMQD5VpF8/r4swEfBINpyi/
ZVrPv7t4w49ao2Kb4ROx1DdpwIlTCNwXNu364o7F1vjaJEGQSyPlkOrwwXbj
t/4XhfsQe5GC5CYf7ngHMdBX7/9vbWZnmEKCd7ELrWeO2Rb770QhHCDNToFf
TNxX03xGejc/394ZbhAKZCk9qBV3SLLxqe3xwg1n6d/VB+V3Z75szjoskWY+
tYWvvVlt+7G2CR4x+jAH90FzkZhSzHlj6ysfWT9+y3E+KDFFx5VQndUYzLND
/6UHXMG2CG7w8x+D+84hvDaeU5s89wmLl00/IiMTmrAbJVEtfOBiThztB7JZ
qEVhYgMQCqrKjMR3W05QmWYpBYtxxVY1VOE5tNAFzqx/WQ1UMqsOnkR/0eCL
nA6UKjANjy9of8o6KeHDmI8dVUQzYWyyTD6kmK6XIxF2on0nRTbrtWDNTgwz
C+SWRetLaaay9CsKZHyQtHZFrauNDNkkT7jtrP2keorQqplRr2g6oXgP44im
XaLLliFJ4jBkjZQLNmbrX8eYsgEQGmNEb3F0+rKgC9ZSzOarZIh77ARkYapO
w4LaL2GKatJ062oSH6nIL2CRucWPUlgkOELNClmY494SCUa3FaYqREAIRs2g
83i1xHSWUWN4lZ5epm/JJmnw/2wIMUofTVSE11W2mH+MH9q19v7B5CAQG27F
zhmXWYTPNKJetgVne0B3clqqAsxgLU9K1bMZU2xwXznv3tn3SS9+n47DaUfM
5C2O/rzkHZXTfk1BwMCuRYQJU+lzH8RRRPx79he4bQYde4fNy0XVicwgiwhr
LesL6SiTJujW+o6lNx6LkXY3qxw3d5CZet/zJ1YXxiLSeY12rpb7qKpsfUdJ
kI6ZhJq+ZxSY3BbT0i5kg2/ZiTmWyNdT9aL9WINrdVU/dQ3KFyn5PBmLj9Fa
rZBesmzdyJLnLBkFtqZ227rkAh4OyW2M4nTAaRGP7Bj8RDK2i6TQ5IPTUgZO
Y7P6V8tyxxklr8qhv7E9vFTOTligSj9CSGCWLqHES/sPeT41lc3BiAHXcgOD
xhxp4AfGhHzYJjMd3XkHzbSGcTh8UkzFuoD0fayeT0u5sS34SO3Cr/R+UmZX
vBBPK7/dZlaVsDBdBlKem3tq+u20yR6DeKPD7KJAHgXHDq3GPh9MXBbR5oOR
2Ka1bTUF5vGk2rMiLO6DLNIvvaW7YIzDCnKWCYA3ToilVxDWa4Yxi7Bdzm5K
CVhC76UV3NepFVBn4Ztx6wAhzV0ApGVnZYGGiOxenkBOdZhwM/Bk2FrD8DaP
TFWM2SmXTbvVzeCP74dhieVYKiB9wMlexha/35T9fFmtY6O++QwZsFChBDpk
iICGz5L+d34l/uqdV5wPif0vK5tN9GZJ25Ar+dlVMwkGMTEsVBeLNTvyrrZo
yRfARCxcJJKjbeZIgB46ZcM7PYBwGQOaFAbFZ60MmQ08esXPyK2nL7l+b9Nw
fbqcr8qdCHN5CZx3lP5+JLF4bIRsYuWwRS85yKeq+1AMm91dqqqF0NwHPqPY
h1SpZgZ28p6BIBUkYXv+hHNrcDBwB1WWUvqs/lE/rjAv6gPLrtPEVCDSX+ur
poXjJWCU6h9v0QOngh92DzGXK6LDo1fuQmuh2Zwll7rJGqlhdH7HINqJs3XE
GExM8fgbsuzorSm1skdfrtlcIF71LMeGUqqsFQYhnTctKzgA8WmCtyFOZshl
oITu3NnHATdmUv0K+rE9Ta1KtiJnFm3l+6fIZbfSgGcHmoqIjtrCyKWrOR5J
1KZBMM6lbEtcPQcEuFSDz+1Dak5y7fy8KSwdCzq1vbdYecXx0mTgqG1ajtGP
o7CbaXuCELVsks8CP8V6xoT89DxS4eB0txFwApfXcnEIG9GSh1szfeiwts+x
sMo86qgtLQzr3x6Flmc1nAr24wqjCngkc0A1vsneAQJTXvcZVpHePXXosp3v
7dTLIWUp2ORnJCXkyGzE15Q9H4gJqkWNIN0Crz/Z07u2Hmj7XwSZooF6e17n
1j6XcasJ/1aGUx6VgOR3OAT7nJJnPiD+v+lUMo9tx35F891NYGpZBaIg0D6b
gLkYGe91/4nd6DG/rcyxly8EZRJKjsRYOAhHFFI2J8m6tL9UgRXsQnusJMUf
jGjamBgpG54lOVnyJEZJR9AOfXc4D9L8oQ2VQY/99Xxi78s6VTdMQhk2lxCh
xx0XWq/XndQhnlQ6NgZrLhK66U2ON/0IHHKNNDTo9wG6iRFcfh/yPWovUx7g
fbdrO3rt9d4YCPlQLwL2ZWTmx//ItrtwUbMdQVV3hCTye2dDVu84bju+C0ks
suKATHX2pXljVtN8kKg1Z4PG+CjIWBEDdMJH1bfDjX3hiLjCZi0c6i4O2mBR
JWpSqDMgv6Wp7A6/M0CQQDhj7JG9h3ENuVnqhCNy6dfOD93p1ZlBI//uTr0D
adN7/CnjmuDICjQtDlTwMch/WckTIyr6G8UMBh5AZDKJeI40zBUQaKPbnfPb
S+UKKMHmh1XehlxyZTTDUK0G+Ld47Lx++iM3PQFzgdCNcIHn0KkoS1lZYjV5
FiGYZCE/rsLDkGWSVyQ13Mxt8KB53cQ8yPI85z08oZoRivgHQaCOBpxak2mR
FyzTLCe3sP7QqCaeXS/T85UkjDz4fjhX45xnu6YMTMvNifReX4Ex4aOvLmpn
hXtqao8NNEM9BUPDsmFVX7C2/zYNNw80lYxHmFVdJCKl0gnvPDFSEB03vkdG
23C6YKjTL5Q66uWVXg6/gnG87uTtUKVgMZ3WfIN8Wn7V2exEDH/pW2vutuuO
w8pzhhU2eCW4nqCUDy0AVABhhRpLMhQSQli9+Ybczr7bVe1h1N2+zU6sHHHc
1CvToBlbBxagmc+N43llMVIllxolwxr3662GJ+8duGJD1X8vZf/V8uBLH2sD
oNg1WV0vuKlrf7iphpDohROQeh/raD6cNX5yzQXinCdMyPh0X979tzyDdk/K
qohlVEM6EO/S09LcfShcfSJwJOUoN/EUhdSrM27IreuGaYssvF+1cMxnBXgt
39M6LkqENWDU5h2VJZUcXrX1L06cFfnFw43SxtkYl/swG4wFhFDji4gVkO6O
YTMvs0GbIVIU5wciD3uQtEwUqce2lGCP11EnzUJQAHS3E+7Bk5bjcm8BLHzv
J86cY52wbhexFpwjMYXYYGA4rXmFe81H9BdVzeceHE9/aDnA/kviuUZzYEuU
Zhj/HTU4h+0plV91xhLg4EXXjhO3d0GLTG725ZhvWm784uVdnIv8YSAD2q9I
/7DVDkArF7AMau8+/8QJvrqbccw4+4hT2a+hS4tSmVp9OjX0WprJFPHorH6o
co6WxcF9j6xoWWqUUSU3EGTCyKtwnV963INrmWbjVhQmoDQiGEXehaVbj8R+
D20co9pqCVLMAkDQ2ONeXE7BIZ3q+68VenMEMnJuCZygGvvCER05ssEfkjhX
HNeb3P2ChDgQgV9kf5MUeTtr4t1b3Oi6vakR+feH+OD88bwO4HSkfmbQyCT2
SQS4fjxWgVGVvIapxEOe/GZfkNyK+de9fgw3rdit0B84B/dwLYPEaR3bU860
FffSFeN5E0fn1CLB+gvCoh4PTb4EXy3Frbnn2+BQbwzI0OYo/Xgz6G0XejfF
wSVVlsOuJCMtLquQfjHbVquSdSb7O487eGHb+z2+jP9s535OqYIHQxJLWbQX
/0zkkAroJcM0zLk1FzLNF+u2N94+wMv3R4Bi9HGT0PafzxfRtLLvv5CULx/K
jg7dhjqGXQnYqotiRdtoByJsgzSG1jhWWOcAh3Gyy6ep8/NC7R8pv1BBFddQ
10RWny1hPayLxgMReKQzhp0+eB7SnbhFt9veOCy10IMdvUDui8Yohpcm3ZC3
wSbt6t3tdSkwP4nanfc4Ak9b6KhLeJNV5v7DbOJnGE4rRW54eGowE14tpnkR
kv78eymv2YugiIRs+emMwyzvD1E0nSnd+/CmtEUEKR2Ep8TKLAx+SAekEtyl
ydSARHCvGC5Nsl2pcqNY1rxMT/nBoUTFulxznxqBQPT/Kb4bLxSnacSG/Sq4
E6Gl1kbU2UycUZu47RV4iASHK+zZIMWeuRn9x3OZMI0iNX2AlY7EmS6SIFtB
KpKdiHkUbG20HxFDjMnM50OPbKA4QhQ45iyDd9tpZC28WyUBJyvpVcc2LaL8
wW2qPkAOtan3e/esCP67MZms+x23SvZywq/XdTFoN2t8s6TLHTqscK63NymI
blv4rB/1MJ81iNt9aZiy+slQD1FNtWlSihLpqEt/2se1x4Tm681LJfQywtoO
0RLaNG7uIfef0nnZa8piv9l9JEjRkoiIi+oPf5snOaEFNZVGGCU2dSpCKeJX
DJfq2leMHvvR17JGpMevJBjqzEhN6o0TjY5ksZ9lwUTGX2WyiKrEIUg0tgUj
6kXMtW5HxTxEOe3qqAgywFPHBb1Wagwj7gcY2t/MFS1tCEA4L2OL0okB4NPZ
+K3RlOt8ttf+QumnAe28zBnCcae0HGpf9LFwl0tBBRNLs3w8ns4r05ekRRe/
9zOWMYnNU6Wwdx3Kwa48RocC9TjO1RdPhKX07VMjhrDlkQZWPpv5iovHPUF0
U4lPDdy05Wd5hhgzdsztXoABt387x49Yw8k6iXp3//CFErF1pXXChepXmbhM
wnkrr7SGgoco6UGgziC2u/WJbTmF1BpnOCK6Dqcq0nLZUBju8hNhNBNQBDM7
E0d9jYXMzWBsCnZk/kisBD9C7QwSWkezY0Rl4wiPkEYrrU/x6ikMTG6pgyLe
QsTOcpDUL9aICP7oeH9L3V0zL2k7t78AKfEAdXMz41+e5jZfS2q3YSuEQ1wI
OBxZE9zG33K3zMaubgdhBNwLuADvPyDY0Bn3JvP+Gy/X+8KWt7GDFMR6cyGh
qNdq0jVF/M6TUoSMOxn0QFW81XTREjkycQ1YXzUplaLSv3YXdpkMk4LYH/EV
Fwu3/Okrh43v0mTHC6G4l1lmqGoxEksh5Li9nQv6GImcF1uR2Qfw7mfL19WJ
Q/wHn5Us2oAkQyC7fLuESn/YN4zwkspdV16fbROpgzbU5SlLWW/UVhzfJtJm
MCKCgINKRzmkzlzsjDjnYwophboJV6nLE3I4AZRmKvsyhTL10FXKe8Fqb2/u
gQvF5Mnn9TNVHpZgMc/RtyZb3W0uS3QjrVhQ73pcytVL3v/K+AvmCkt6PvID
xKxh6t0rxNW45yB5Fu1slGQY18mvkS71avZJkzYLogEXGd0Ua3SX624KVY8C
hFpaJm6bO0kxTbVh17UhovwSSp0/xL191e3i7xgzzWrnT4VeWZQPJcqrCf46
1XHyfou3jjP741mIQIoJcz0fHtBTKYpFEHg5lgboIP57xRmIQz9zzV2YiNyR
59djeaf5Glr5TYXHX/yh8LNNb/WkL6SaDfpUAQ7aTE2ny/xsOtgAZrdB0I5X
T36F4NXd/1vm8EKuFjxm0vt/VEzLyJWrjpwWXtMHUV40TpA1XAhuUNwOmt/G
gistBFoRgwwm6kAmGBjkFFe7xae6xehUx/w8Cll4Q/XrzYCMVTaE9dduQM5X
t8yCQ48nfBVtTRG85L8R+9U5OT8wu6SFNm3kqyfPqg2XmVC7pHKU6X+JTPGv
oZCSlQ9qD+rT0yx6Xf0kouPzAsg2lE5n2QE7EVo0FJepLBiW4oCt7UXvXQC6
6wLcPD3VMrdDBtUSTMvmin7QDuWf6wdBXzwdJvahG1dDZrs13IwzOdj/p8Sr
3eolIDFP1ziRk3fBoPA0hfq7/4Inir5d+NzEnHtznoudpHd09fH+0RIfFfMx
U3/C4KhW8vSW3AWGBDNfOmeIBSD18iM3djuVavTb+H7oGkXdu1P4J9/4x6+p
OBLaxLwuWes+6Ya+YJjZqLnbP1Njg+fu+oDcK7xOGf6ugUCup5bxykU0h7UZ
4m3VdvnjCWuU+CV8i4BbYYXCqS2wClLnbaeElH+A6VQT+0D40TdGIR87ujiy
GmXABJ9/XKdJovPLDgCSdB5KX/hGEPS7UL94ooHGurBPn+zO9O7RlCEf2gXv
jLuJ6kInt7Gcb2zKLuo4BnQKApWdSeVJbjuYp7QEMsl25lZeaLjLy6tw+2MY
1NX5bO5Io4HGSfmUIv1CJIdKI5yntYHVtDBqRANc1QPwM8IX6iP2Wwqwzk5i
MG/rpZyZe/bQjZLMc+CM38eSLsuh4aPxme8TDw6gEx5yyCgxwoyZG1t+EGkK
2BPncihrDGbTyE+U0of5kEA+AkehYLfmIQQuUEQe0sUUb/lUORifAfGi73Aa
ewIeFYpVOiLtb+ghQGLpQgXqL1/uaLiP4Lr1ptbBNG/x6h0WoFr0J0rQ4woq
E1GRqLFAsB2Gkz5VSx0sBV4VJdD5ZMXjDpaCFdp/EKBvBNHaqdPjf4VLSJQL
Hx+GckMqgVsVVEKMItwLxHR9GGrVTqzUvWFaxP1c8nFjeAiAQkHRKuD+YNxq
G0j/5byUas0dQFTmYfCuZ3yxxz4pqFqI7riwfY1oAyR8RjcQvtaWRGrUT7fj
TEwiSiy1gM8GJyEeXJS7suD8gzDy/SLhwcS67GTZgljM5Ff4I1tbr7IpbFhV
8ccSevlRIHkadQbGP0TvbqMWrWGBZstVEbAnfpvNRwuzC0LVAqY1jtxRh8+p
43XEQ3AfvN/v1N00kUlhqKjGxDV9qreIMnvDua0X/9idMSlE7laTGauWzruB
tjlkdY1CoQexUM+mMUSWysu9/8VXJxnpY8Bcrl1fcDGHfiLPA/q/cvY5a3hL
ckmTpQZJdmGbWu++NhjOKeo9D3HagXdYsBFIKVaD+W5L4j5rVp39AunNwehv
dO00g08NEH0cxDsViL0XfIzjifw6D9WYVPu6MH8aUOIKe7CxHQ7B63yLYtjO
ponyjBaM4M1STNj1OBmuboRe7WADeKd6daXziTU6hM4x4CbqC4Lxm5VYl6us
bVejNR4lx66ph0YcCo4T47vFX3W6/dHP/QE9btEaMcSpIIOSoCbFoc1yxK0z
lHjAMjuJbOe4hH3vTbIKG8MKiXQphWvtZ2gXN9rVnmTGy+kfpgnrkQBYWleN
8B65XaXHu7VodkjnfQZLewjynb4KuJ+q+ZgahhczWcNP40x0zv5W5oIDEeY8
XPRuPheNes66GZ3LypJP+KqT6KOp2xk7Q0doBAfWGeoBz+ZEdgZD/1ANhJIK
nPKVDb7kSxbNvquqwVskQc3B8M2aL8FrOpHKe6jzumC1A23H4+gwr/Yw3WpH
+AawVxqBQOTKLVaFPbuT2hHk/0860Np3s7NCZZDVScRqqRPmhWOwyds3riuf
YLENr7dcEef1eeSSCkDkxLKOkK3FTYNoyEmTYz+gafiLvxRPGygB2iB2Jp3m
kzoUlHwzXgtw86gzb1RkBShj3ALKxLnYzFJUufVw6Gn9Qs3Uf1ssvnRjyLne
uT5hltWH9osnSjoewjW8xLBZLq9SE1dZ8jIDF4nPgkYILaM5dJHDkP6WlLCi
6bOp2GkS5FYRkgVmoqQQs3wswVYS/uqTr/KGeLvIkiV306l0Ev7kiJMrpIgf
77n5QExQ/66dgRx0LY3MJGHa444UiABNwB2pxf1EKbNN5/Q7dDd6MuTiSM8x
T0Qj88krRwGYE8NdI5e9qVrmHgon1bbl8tW7mwPhq2tfoAjCmLJ6Ip71T1ZO
btkPt06R0oiN8a6iZE5KKmQBGgmNq9irGcwIEJYKgW4oNMiM3dNEOQ5kq/C6
8MZ7LyAjc9Mn1QdRAc0B1nUGAwgT5EJnq5YoV3hZTK4pS6uPMqM/DSSjRzh1
6TGXp5bhPf8TpgVBl21v1+/Y/gsJhEFRcOVJDOsZ+aNRuyc6FbvT25smw8L9
9MDoNjUQfOsxYDxX0M8J8JJBImhwGVbTQwIrTQfBran6zBtUMH4JPf4wiBeI
PBRLzzKLYUm9wPsWhrp+27CwiU4fZ1j72lqzRctQtb7etG7btPbX8ziUg6B+
8QfiOoiNLdvdXAiqHJA/5rjB6KJ89dBWvrrf4Fxq5qV5kZ+40wxKr6Ry1i+K
pfndGkt/2W9suiGo3aKgEsG4qpTCccfxFBKQNqyBf0/11r5uXr14oS9lXoXd
0y6zJpuyknfWwlPPQDIs9WW1nEFYC8lVCEXrxZkIbr0Qhtf/wpwvwUp0H98z
cft2ALy2xmaLX7/Sz1yLUFtc0H5vIJs6UXPrsBtnaVaVozQIFke96xgZvNZH
ibwTEpRdrFgYHKBPhKfILz9lLZ7l13gpJW1sBSIxwYdTU4LL/SJrcYqycVSE
6yYHaEZ7ycxsg6YbC1aCwF+2ajbV/eJANtxBEyCTpQurt0W1V/dD7ugDmQfv
CslmUbJN1GRhGotQKSoIewbljD1ctQ/peR9ga/8VVik4NLLqb1Q/OjyO5Sek
2Q5dFdd4XfHYcFi4F6rnX30Wm5iDDMcLJatfpedpGVO4urVVRvgZUFe9Tolk
Aezf2Mf8jOmf8+syXCJKNwt9B2kMGxmUwebzT9hKbpyiBq4v7Kl8659pVyrr
eCjIldL0FeeWDKR556opM4Q7wEcpX7PHhau8Y0valtfCI4ecF9K/R1zy+zuk
2yDa/VUY6Kg07omSB2tGMAQTI2S0WzAnHHua23uP2n2Gh+pOdKXPHAWHDt5K
496KVgw72Kwn0wYwtm2UZNQwCKuomx0+jcrqRwPerbAiTGnnRql7MwJv4VR3
E/66dlKLsseX1YfI4237x/mZsAPPki+FAQwXw4nxk8QVFRqn8HXLaKuWgBpu
xwjrUYnCs/KyfZxBmkWC4tr8QshsOq0vl+3E37NFaEPbGLnQ21jdcYRW22am
WMHMZTmxGMF9BIgjQZBarhjjmnfP7fL5hkNQYtlqana7M4WYhqUxg+ljmoQ8
1FXK5h1I8jtC2JnRr6tGSFumh0rq67fBtfGSte53y0pc+8Tm2OVZ70ZvUTwK
Q18VuUY7af7XvlFQC4LHjghu8gNCgXFuZ1i5Ts3F0BeiemygE/Wi8vn0GoUZ
xoAlcuGYcAOT+Pd+2SkNIYhZmMWv1ApsYs3oDsmCuiEoUhzdoQGUX7vRo1e5
eANieJZWe9XHILn/OhUsAbDS3vFdsecpZXGl4UTJny8LV3vQePX3NV4GHsj9
SsqYAsNpoZHa7yEdSSzaOzsrbKJQ0qsuHL2fUNbpC7PDpnKdvnBmFT9F3A6k
F2ugDRGO45W1trjQYUwT9g2B4SRdQhfOiDU9vY6fZMrNaOJUbqaf831P3+Qv
8Rmj5dS8v+pcaOuCxqrJ53rT4KV+4A4IINRp7SiDAf6paQ1T8aPPancAJj3c
wp5xa2WR1AEAoBdPEntFUv0IFx1zNfFqPahqVhhN6ozCpzzDjXYOLjJHCcuA
aQA+YLnveG0TRqQodR0SIP59CRtiTB1HLikLAMbwc29em9BI/gSiRK5UzWuX
ot9oSQZujZT/ziBlXBiw6c4ZvDjkFFygbSfdnadUIYUbMOvnFCfgoCsqnJNw
rbW4bXmK16Eux156+6XgHsSe6kmSwHiNaCechhCS0eihJ2AEXhA7Lpr7x1E5
zfskqCcwvKio8NLaPhxEFxVf58nnwCxLwvoDGLC8RtQMtTI5RLJRae7xARK/
QR3DSuzLj/t/ernoM/30iK4FzdOmjUloz8ruU4I5kqC7Bh+MlVJ9bXmYJkEs
byVSJkP+dxwOnD5syyC7ByxdQq8svmqv1JNMc9hFzoG4JN2fgPOTp5NRpdt1
M/t9gJE2YqCf+P9TqnNzopxXSj6SrFxfiF+4N4/VAD9KijBTg00B6jKBW4X5
dge7ns7OGxtiEIrp5Q11ZwIIkpK9sIkloJi+/tkJLewxII6xoCVVNX08haez
khxfaaksgd0Z5jv1A7Y6yYFSVSZZkHWuLoXSrxQNeqz4Kpdcg1BqWDGjDMyg
HGfXh2QbDmUPlS1Jhtsi40AidQ03Sa+AiNiFQFT9YRZX6O5B+ablil9LdO7P
kBmL1dd/VEAqqzqwqUOHz9twmg+kS7kGKDJrtZHSmvQtC0/DyGp6kiTPSdJy
Gu65vfsGcmfzpOIEh9tc4s47RmZYKfexSUho6wfKu4fdizEypKV8imnr9F+e
liR1istQI1619g2vmN12XrjfQxoVZAJLmBaPCvMsG5jrJP2+ETDsMysxsYIq
h9Ocs7N7EHRlArjeUi+H8hWv7Gf76lUXqJgbLStYu4FA70Q5zCfDz11si7NL
x/9HF8h0cTY7v0b2TidNry6MqC0VZBSjvoQ12vxGwVcs876QaezKfO0/1yQX
1U+/dEjKSdzE90cI+YzCC85KnSpHNvK2OIfSfMWlXiW8znDP5Fnb0KV+7MEd
UunQc1WwQ+grXgxKs8yNib0naHIj7LizdrLAn1JG3nHpzT8qWiUGb1CMI//e
g0d4pIE6HIeUKXtSJ0yINuEvZjt75cyQ0iVOIjdSGVjs8i7zYxLdJL7IJohC
XMBUi1ELRXgbvsQRnoWi+VpmUBLl+9u0rDqd/EgMWGzRKWuI7hRrm+faMbYB
BwkiCnhhqA4IcxolFXisgzkfH/E7OAEcaD+S9Esfyx3FpNoEpG0t3Gt3y8Tk
INajMawWSmqjtmyv3vAZ0YWRBID7hro97VLPb45vbj5xaCGId8H6jJPWD5IM
lKo78RBbNxq8RtRG5DLU1xE44cYQFb0b284/gpgBzs65DW7urToD6BLNy4Lz
DbSUQMrxy2twxQV9s6NnKalSl/ocYc+3TZZ+IrZenC7K5ebi5y5rWa+XfWMC
q+SEYHZbeLM5Mj/fVDLJ8+4jv2AEeqHxPhBZHKzjg6WYbCmQh7DiEhrC7PU8
DOlc90DMKb5NcHG3Ep0R7rkxdpZol5QWUaonW5fxeaFnmywiWYfvQcEmh5bY
V4YIFCQJ2aLvAKikJgVi95KFEUosrIlZmBNcyPpFQQ5EZpg62tQzArCXaQ3d
LU9JuxKiWTcifTTDrs64AZdQIE74Hw6dpokHv5nrZB6MAwX4mU01QYV3E51N
QOg/3CsuA5pyuPGf16yvCDudDOyY5cC1f661GmnQ6XeJcP4i5Z4kvnSsDvQY
2hpHEaYMnQk0+GU2zz4AnEsKOSdBrobw9IKhNoCvUipatnGJxj/g5V2gpqEl
mHldVhvY+1DKSgSA2I6mNfk+9RVhhosbCMXhKq/yT3OGRuk0m+ZACkagKp3R
eSn0L1zftd821yRQ9DCJKRt6iaCCmaQDv1IS8rPTClYchEJGS2hH5QL670Au
tJnQHzo9whe+DU/q6wJ4GLqnVLtwB+fYj/pslFCDZiorFiQ5flAkE2gDNdog
b9qGIX3jYt45rk0bwQySIfkWHMEa03W+ZDQyaWZrRwWe3/itBz40MZHp+/mT
gEElhwyoZqf7vpkRuYyBLRrAcvY4+juEjDQDrZAtImhmGkuJECBzliLzJpll
GCeb5ylg2HYImpX/5S1bacG1wArktKnp0V3elVaOVCAd4ogWBKOx48Y/TNFK
r6bCOl42dnmmifRhivDk6L/TPdVkYdCtaJPvllZ23RE/1ZcqGHmHmCs1z43Q
NcXSWHNtveQIODsZtbSYVIojipS5OlIAzDUR9fBc5pWFRujgXIZhEMUd6hAA
8if5RxUymlLz7jFCUNAdRMtbRsK6vr13mOJBiyYIs3SvSStMRJRchnjmjJcx
fdn3p+K/PC5qvAJmbqnC6SUyfdMy2zECSFEJxu7jEPUJyyEYUHm7WNLAy0ql
Yf9zsW+yXyzet7GCCIp/eZhR7lySW6Nd4Gjs4RUZHWDIuuV/hr1SVFvYcMU8
CQTMw597hCYdys9P4MNSJW6/tifxyd5dqGMUdf/Sxf+KiZFnN4jemlJbLvHt
VX5Nk4HfpW05Ee86pGW78dfaLc+eL65ImlsAx8ZD0xSivO9BaPE+d+Rjo/cf
K8H6ltgLjbEliPSxLeT1PtNn70P6H6utuhEbZQ/DKl5pMRWBYU3Mh/Op1Tbi
xY5U9NW6FOqyLwszLbA3okU8veSFvfn3GSjo4XuJcEQRYzdAWUMjcnfDkOs8
baFbqeTWj8LemaW9LHnGGBdKDZwn4I9arBdntnt+1cRP4Qqbu9td1vr14i4n
WqcnRjn7N/UeXLJIGkSB2x07YsiJirm7oVX/0c9a7EFzlzm2MlK5eFipIZxP
9c0sIuLYtbhXxR2FXftulid1RvWgnl4cy1kLOzwtQ4d6nVxzcjMB1T6jt3k0
Ix0XHwL4VmGva2TSh0GQ40kNYq1BXFitbeHOAxwNc4dE8hIBzhQJvRPaKU4w
oihBgjjIg1guPpqDkNJyGM8KmWu7cPg9gyF/kH0y8tXY3Bv21g5L8i4xbywm
+HpPChDfk1x48SVfGHlIq+zkqQ7AqPAcmmeeJD+ZQT3ST+B5w4z8R1Ptndw/
8wotsh06aBVrJVnkpVoFmUZnIzftPKySNGlBCn+g986K/crMVUTa0So+LC8B
2DYHwo4DhgHCM7LQoGBTPEHQLb5vcGwRKpeaJtVfJFURtRVwc3YYqpuDmZgF
X7g3ZHmgUTw/q4TkZG65aWiKkPBSmTHgGK8Rj6GtCwbyoAjEedcfycjxRWZ3
Y9MydLS1T6cy1Sd0/Tmu/rPFGpiMU+mF3Y2iBOR9ARGDLKrfQNAyR55QFNCV
FevZo6pxyefzxVeXdIlVWBdT5qyU6IwuiUHwGqeJDgC2SoInQEh6F2z9UYrm
99osCQ2f457tV8pELMb6a726z8aWZQYnBIfS8IPQmdidKElF+JGHln51Zb2x
la1uWzacTaJd3QCB9LGvyUR/W0bA5vByNkH7yD5sSnUV2Kg9buGg7WgkkQwc
T/ApvZPtelr8Ciw0/Tgns6JXdCuTdY36eDMjIACdp8ms+k4Q54qJOzGcSryG
g7PN8Vqv5U3tQsr6AQv5Is2Z860dRcLuLFKJTpOeL793sheP9n8tEK7UHQBX
zdkPM7/K41ge1W/mGE2qrUBQfLCfhiN0EgjQGzDQkEImVsP1RU2LL8hLJ8G7
Pa2C3g9UcUHR8I6J2oEq98t6r6kLlfgP7CsihYtI2LBc6ToSYR5Jm9vXoIBY
W0PnjidKjoBKvUHyGRmVtOn6VLAEcGHJt+dLku4dfatXwaHrKCrs57vWPCTS
XLYjhrf6VGo1e1bjBbt5FblrpxQEefovNd6fYfXrO4OaIeF16UiYXLw0VdSf
oS8QbNWp4yALr1jU2pN3KVdBJfvmLJ94/oGKnDnUIecEZ+RPCOfMCeDTDkvB
91TiyayvE9EgnCx89PzzzpiZy9RHpVlszcmkXloErnCiPZf4fG8M66AO+Hi9
mTg6y5to9bfrmwIKqsEa2eIK82wtdkNI1BDPe3dKGyDijmECZ4bAQlWZscJA
4DpjrjCGM6ZtpIXSgKrH9guVifENIu4881xyqhw7AbDUlWJHH2W1d9kJRcpq
Toj0z5zKyDdvSN4OfJ/pvzx4cvuwy36pWTAxFO+U2+yJYdJSPAMCkdguho6H
LtDWsg6t2oJEZ2IB4J8ARjPAzC5iNdW2SOgnByJgGo6htRmikCO9no7/Youp
qd5wLkjHA3iF8iDFcRNiendfhTMwMZNTybykaD+o6npD5iD4pCsucduiF2Cn
VzIW3nYOtby4bkc6SbDEtrIcayrqWbuWqThvjR5G6lvD2WguKA7uvMgYlPGP
UkJz9XlOuTMtt3yNXO/iJfB60Qs0SC8/5Pe4vjRqJ0AOO+RRj00Z1AR/wTCw
pyS4jyCKH8zEkl/u42zJFItcWhDpzJHop6Of7U+nwd8zfV6L0rAQvK3BD7BJ
ZOlqfiF2ZdG4P0NtUQR0Zxy9mDl+Ce8R1Y4oRcl9QNqtCBfFReXYUz8cGmS8
CV9/ZuT/UBf2yurxLp1s6qWBJB4CLypdQQD6nB6Gdqs4FiuZqpG5RXj+obQJ
1spiuBRiW2b/i2/4tahemG5DsFpUHn4pPlO3CVkM3uzyfs/xQ1JfcpPSjuHW
2+En3X/GnJlG6F7wQJEkPlzXKJhhBlHXD3/Ksj0sCqk6yhtkY+KLiF/9Grp9
UjbTWYq+a3ee0pES0PWQZ8SmkOJbGGvWf7sBPTSf9gTk4Nazxbsff8wMIdqz
/eh9F1dgMRPx3VEiWjw1ITFIzccHv70Yjuy8lvEt6SGZ0GzUCdgelCvXCv3i
Vs2M8uetR89vR4Z5fjt0wYfFAmoRjX2XIiCNN7tPke9g2yfdf3WrOkjDntbh
ZzgnDI5CmnZJTJVaiTfIQSBOF300UlG1d7a02SOhRPRagE6hOrz0QKdt75ae
DzI2aGqY2Hn/Gbawgaj31aIASi+17Yl5AaU74xDWRaJzf0LHr2d3aXB4NTmz
rlUepRuDA+ea7vmoNnIh33HPlSCi1z6stuGCT33WZ8MYp1wvqu+VD8yd075I
ildfpDdoTySC/oqs0N0XFB+l6zY7yB+f2QhCBwTn+CNrMFvEY8IxI6pahfkn
rEbndSBLk6du8k5qawTGvc9QjZtUtgIRcm0ue1uwwYqmfn8CGf6Anwe6PDpS
pAGfIGAnohEaYn3Rjf0A8WBnI5j84cWKntwMGNm2ApFSkvvOZw7gC7hVWdsn
1+oHqhe+I1KkKyBkOkufJFF6JqEqR09b1woW0+2m0tjOVUsHuGb/O7JWlTyO
TZhRFqPmAi6oXzWtrjdCxD2KFXAemudDVFVXeoaPVazZI5pGP6DLDhtblduI
yqx6qb7EaomgAI6sfSemO9vd/A8sQfHLe3WVUMqqCfwf6ZQiH38VUaw8q/yi
7dy5Tr+1wPYNWxxeNrTkB7PpHCXHOzdcZ5xJc/+wCB18shnsmC3rY6ZpFIYZ
5NKsBFV8jWBkcHxVZvOT1fUFnV8DbusxAVGWWPsR61kAJt2m1wIRsyT9d9MF
hbdcs/dvYnZ1mlIz7tEaka/HMw/5Kdq7NHBFpFWD8JloR/FQYxIa8zsGPd9m
kxkCLasifAyGJ/KNRhVxGsenCXVfQgSzhPw5xvt7j3eHryPjcnpDNvDhlVgA
Qt/hs/Ag5yXxwvWlk0RHNsKokSC9g7Oixy4WhZ/qaTL4Q+iRxJwIltxstkAx
Aw9y77ORNA7mzxmX9dsamzz3Y3Gkwy1iQCsSHqaDEmjMzQCfhzarlHVqWoRD
dMBxJp0/5NhNhjorny5JCFUAKsJHqTJHeLvP8jSW4YzOQYKXClgFd1ZskhjU
DA0ecLze0AgHzZiXRjeNWsUil2uwbjM2AG/8ruh4TFNGqAB3oJV9nJXLQDnE
G34IkIcYSQy5M8sWaSJyilc9JXgq9PLUUrmXGHLagKq2tYqhpjtflRpIa6lB
ri4eM38AVk9PH9LBcTS1c+LsJ/yZo1+qmxPqf1AlvIBfvH6cYe9IIcFFwBKf
1BOrpmrE4g5GuTSBz6N34LK7QizZJomPssb8Y51HKF4RY4FPoCeQQ7yEEaxa
7sOBFb33kkLme7r125C5hAm6RgQRcDufZNMvgrZ1AEA77Sb2iBokZ3Es/g3r
TzMbSeX/KhaaZcynAFlWE+uR1/8coe2hbgHmF4kzo+L78J6EwA5OAoLbTqTv
yO/LlTCDLOKux0D3eTNpSLGs8JWFiVLap66LjvDYkColJgGRRkGIj7AUdKqH
4CBVPE8jRGUWgr7QbL70DXQ/Pw377xffMnnyi+hA7xlzic+1tpEnYZr6CV46
C55efGK235ySrWOMyZ4J4npcVd1rrWooOBhmH5EZK+PydsA1qhKthiJto/9P
XEFvfRFKteguxjjBBhiWPtyJ3gHhxu1TsvLXJVpNJOhJnRw9fYDoWx39w5dI
BK+HS8INHLtBkuqoqLrs1Ndg3oWt3xhFAO0J4OqiJiw36QUhx6S6gjbl/Exf
M7NlzF074G42Gd0rPHVOqPLMWgXJQicpalT7OPXUw5OO2k3oPn+WPfp56Slu
NNKHApqVEpvCFXWeD3omZFkov/CbmBrHfMbl/4/iAXmZZdeWQrcdR2C1nW3r
jrTxXmQk5qQtvIkE+I5gtCTol/w2BWAHVp26z18b0gIWiEeswQmXJQDbM0Sk
PNcOS+I+pFSfszDG0yyk3Ky7DK7JOqnC0eEMgC8Wn++qedkvyfOGX24d0Sqe
uo5uYZ74enuZvMYB6Ndw/zziR9bdPgb531G+lL92NyhAmxb069CEnuJ1PKAF
9ZG6u2PWTSG8Gfre2KbITDdapE4QME6xiF7McrKGAPnSC3hiYW2ws29hWabg
Nnh3qA3aq692HbAO+zU8Bw4CywDu/s8rT/TMCIXNEw71VHv6VSGdsZsQRnLZ
0bQMuFcSztZQIMeMG0LCVvCEiipG0rheiqNnmIDlb6g4Oqv1YsPQ7ZShwSvo
e1fAZUOOYS/JER+glNCbvLNSn+YxODHRpPw4a2ca1Ozm9BYo/lvGMnG0AMxh
+xF7A6koEL7Egi5if1Agiqk7ZJjv9glJtX5KHCZt1t0D8B4OVm75r4fjSiSa
rwGVMzmD4jZqUmek/fEq/K1/71TrgUchydDOYdR6nnRemikqhGzb94Q99K/D
qNqINFQCCitrYiRY0GZpI/XGT1CHlfAzeUeiSsarVLYqn33qgpA+6K9iL3Zz
lqabC4l201C29Xks/KcMxbWeaf79DkbQjaP6lMJyik2Sp0DwtbAjSxKWo5Ft
hfG2RRG//uENS2L7FxetpjypN/zU2AeyULQo8FAE0xaFgwxwhZPudi4tpiCC
HGZmJCjQEW1+92+G7wYSVN8NTYQHA3ij8I0lF2NgW1IBnvxDYl8zpvEZHf7V
LcE6iN5BfexjwrTRXvF2OP0B/wYS9QoB01rhp25mx5jPyEMzlgBoCvcUx8jH
piaz4HMI4rp212ToDh4zfVr4ujk5QPZkYdFXoGZCy+df/Bts86KKBhpSDzUW
GQbDEsLD2CZlk45GX6YFzYsX2834IQDOuzpPrsD4iCmgqLW7wAOXcSeUITS9
QwyotfckGOqK63S5//Xk/RIEb7Te1qvz/jZdIBJYlaezW+T6mAMUrpbYnwXi
MMlK3K9hsBwbhEUjSypR7Cj8VV/yB2BRs4B8mGBmTure0I0it6JAB1BZbP2S
WZxsDy/HLKAuMlt8UxyauYkTpqHrqMcdhyvyZpgaAAwDc6JJ2COstQeUtoMo
Uh9EP97ipM/EuqxqRi6UqNgLItRmEafelQmHpVGwO8VIDEU8y6EZXbiej2XQ
p0JrXAR/3fWH1UspQ4ChwvG3nOoCW6i+R97FzuqaoaVFQItViv8hJiD2BHw6
BUvbNTcAEcjYiYQ9vgdvjGhh6TmQyvhnBfz6d+2ojrrqcJs4q/qpJztSPvgG
CLvgnkv3zQKCyMKjjXh3zeGjb0xKrTny07YjzSawmLmaRcDrUZPAKCxiH/SV
Jkf4JIw/ywyzSZxSeLKfchoHx+ZpGwMc0RuMHPZ5TaPRsdhlgBeEXbe65HdR
WDVyN0fRqTAVwKkHRJalSvoqz4MNw96kQqqvVG5STmfipMlPXB4sDQ9EYJG+
aQN1FoVXVCw/rq7mWosknydgQ8M6sAOR6vPy4wEsKJei5rQ08pWsFc6dyWPz
7cDFauDhDocYCYC1Go0CnCRxoJCpHyiHOdEcBT3ucPN43lhLe6/xd9rfELoP
wPDNpzysYhNAQBijEAyWS7waT9tE2OuygZ0E8+LV5a+R23SC/bRWbaFxFmtv
MtL+fAh365kVPbjmMa91OnZ04TRTKfPNgXxYPUNJWAXVEpMd5zdeAkEaCFbA
wFTjNnBdDsOOcu+D68ZjhKghecsiit9IhT7IeBWiy0CU5vnXiQW2mYjKoGtk
NLDIYw+13cNZQTfStbXvWZnlziiqwnS+raXdjRs8n5n4o+Q/svqVoWgcCoV2
SY49135h8Flq0X9WBkmFEAoqC3wr9VuuqKhR9tSWsKxlNHOfcL3hYR4Gabss
LTuP//tiYCM3DigGzvbwVHO3w9V/Bo22Y2lQM+omeEGUkh0fffFb1W8vCn1p
XhIvq/5olJjHIFGj4YY/r1frG2cUmdsJxKkW2Ya8Cu8+bNrZ7t6QcmeQZzMP
pKJmMTN0+3p89qlnWJdpc45Yi6p53ihBFRYeT7iVvx9K5liFNWdDAqiwcMjd
0X372JMzUvocLuWfAXrOuXurUZzUz8ZgzbvvVuelwvO7C+QXWsHLkeNUv3ha
iJY8H8/7opyBTZWj7Sg4yOqR7zcDW9kq8obcJlx6796k6hXU0EPllc3avWOl
a/lCIEx/hxGv2Ow2X2CPyq6Wt9PxEggO1F/YX43d2YkwZHxenxyCA1UyQWPq
BTMrUTScTFq33+G3Ksy5eviOwOJYB92LRUa+MuKgMkdezP6d47FAGVDogDmG
cQVivqfgPdiOvbJQ5IMe9AjSeAso8apQnBRKXRLq4nKtraCWepY/8SEDhXQA
vcN5HQLMvKYFK7xin2pZxtU/8Ye6MNS0Mv27Ym5BzgwtfLDXtemMj+tTGHr7
fpeHF2ij8Db2fvQO10fhhczsrlgq+ucZV00Uk/hP7Vc23Vch8RYW8/iEWo7e
3OSOhn/VtFZZG0sytT4seRSV+zM0wTFC2Ej/cOBu1+1v2HKs2/1ys4g9esOi
+3c7yE/loZA6pLpfLNmVXpgJANOKC9KwB6It1vUK8dByfnnAjMlMkXe8NwXH
n1s/5fZCteZHbsB0vNe8GqKcxlIXnIn1tlwFl5bg3H8texgsJX/GTzwdGrzH
5K0G9JsggFs5mPOaLbpJXrC8iTcaTblaQGxKyPklOIFLvA45tmu7d1vagb8Z
9Kq413ixSyRwE9TGzJxObrOO/7JjLWw1IHIp5D2xVRYmg/GjZrgo8d9WCyR/
aAVGs+OyQ4yb6lYJ9Co7aA/RwzJBwLbL6yD+Awy2UhJ9sCswlRcWCf0YwLz4
GF7UfoBciuhtU3V43XQuA5yxm+1x/aFwlMZGk+MXgCHAiaAOMhh94r+YR/tl
6PtT3P7Xor9MJEmkfcAelP6/aaguhChazIbOfLPUYH+24EJ+lrAuU/QwahX5
ERF/stLgYCpiOzR6QYR9G5VBXIeHsg/KkxbRi8J0xRpmLBd9bWu2LRHPlP+n
9Xqzdt7udnr8+n1oiKNTidXmzhsDll8+Xw4KpqXgaNYj1QC4yqFYKB1oly4x
O3h/NRgzfJJPARsN93hU0rZnaobEdR38cTJ2aI9Lq/ob3GCzJpgqFpuGb0LY
998EyJMhqCryTexmPocTXY7teETnI8aAoI3VL8R/J7WwhoPfvO/ZZ+DS1C4Q
RwZJEDYDQHHwMXnMQ6WJpanf2u8nqcKrrQNihlJ1SbFxeoiFZWi5rFeJfJ+Q
yB/IzRT+faOuZnWaXbEKvKV9R7GBhWWrCALJF3m9oZVkAVwGUo74jklXRLJw
ADB7qKiLuYb9FUPVq8nRD/M25jh1GZGg4Ww9lyFdpmR6BnfiKluUZbpQ7R+d
2y6M8AOFCEAX0qmHKzU2q0AfFz5pCNK0qAZt/IEk9g3MOc5nLjOoRsQ2rboE
4OFTYMCvJEgWPapcXPcTa53i+1Ak/7OU9NZq/64uyaDzoqLC97LRdBS9rtEn
+yI2QAg7UTQmEvK6Z5vpfjwp3xFNbR965xIYG0gOEukiVhGFydcowdviptjO
rdatI3yQS8oWgpJHLAjWgAzogkuNlpuhqKTcIJsl2k7iScTlDWomHDWgitEj
5ZebtnE5BVmRQ+NfmZ12D2CYwtRwsanhlKjH549E0qA38OD+Uamvo+B929oH
BsaEgaXaGCOZc8QNQZ64ODsX1dGDg9ysFQsLoeG2inAmsnOkTkOBqrial1qR
fLLgTtx4t1qlLAebZzcifwZ7gJl3bHK4kmIl0ykvM8QFEU3x21jUnCP5chvl
rOwLKh4JohmbRZAhILCGiHkQ+0hshWoaMypg3AL142SNERmBUexXSKiI7INQ
19EHo/5B1WoY18WYBxApW/YssfD6DmMt73Er1NKgOPbsN/Hrq9f0RWqgRnd+
e/k6ysWgB2KdAUBZ07jtnYxeB5N4eYzjO2zqjeQgxeSS2mZiou0lna/7smX2
weeUtLfU1sNhr7z4Y5+P5qmXeIPp6t6cuHDH9Fy6upb5l8DhtxzCRzB1Hs0N
nNUNSWNIHGzZec8n63LznbF9de9dEBoNyNQCkCwGyR+hUKOdlZfbWwtwlN6p
fWWYF7e1F/WownoZB59I8Wp9/bjUw8tD5s4EVljiCC42QSlWUM6AFn8FSEjb
FRGNXJUhZ00livy24kH0roa4bmJtF4Uf6bmyERoiKb6aqFJL1FzqKJgklhLT
kpafAixOGKsW620yRZdwKgmVfxNs1rjIvYhm/4ZKURE49q8Ly5i2p8k9gGAL
0UGFqNOfX/Ku22XcztrB45xCfE7ClUhRn+x+x046UGAr+4BR4+uVDA04AIPH
fpPk6yjS0QLP7rQglEebzaqGzJLgaP5Z4AEmeQnvB0Q8KrfwH8yMDR6qXWn5
lgH6ALd2eeQHdiIpKRC7xc/xQDkGXK4qv7tBJdDKQ6UtVBBstWylx4OA0nk5
1KbG6L7bFf+Kdv9Q5kuIXIlp0EK/ykVtSpe0oDlSuKEELrus52HMCn0h8XRh
9WGlrw+iwDnnBnMIteRZvo3Tl3bLrhvYurCEHQrX0wfdIzDdsx8CgWrhrSCZ
R0CoFebBNRcXvBE5ydM51Xqt1FqrGHL2Dn70G1D5XjAvZdyj7t3omxT51Z1I
1C74Gn+rEZFPE971aisvsn83mkUHl1ePAr6ZqwirhyKFGGAkMTqC9j8Fp07o
vilZvwKQVcJ7pc+ezGgz631kEU61UBfCLUfRIl4NcpQuRxbfSoGgSv86FSeX
Lica+Md9S1UHBMXIgnH3GVx0+npWRG+WDZbeB6W+t99/BcO9cwdIox1JhjRb
RmZyB1cUCdIJ+HyhlCl8WhdPW8bTqQrMeey53WaY+2c4rksVKLK4/4Om3AgH
b2p1cvPsPSbXS0OVVZBQjouYU1fQK3vdqDKryGBHz9s8TWq6Lk3xg0Fpte0h
RS8H1o0MjlR/rRXGL/EbpeIwrd2XgziKF9pYWOICwpyfHun/3REZSc99fz3n
zyVgrmN5b+8fEJcGJCeeynbsazdUvZ+mp6cRMPRSdhAsSIzAb2UASYHLNf5c
mL7duOKCGUS8KgB0SppSY3yYqE1WHR8fEOfTmFWKbh7J+E0fYQx/478zqHPQ
pnL4NXLNp/NpLWq/GvL9R9qxCc0w5cz/8lcQaO4trrur9fh85n8Uzd6dAElq
w7PJ+3sfHVUMF6ln9pYrfuC7y5FJeS33zOJ7mmtPN/6RnAMZeVARwUHE9gjZ
mwxF3/sDtfvbr/065NODbFrblFiKRznPMu2leACYotJtJxvqwhP033dhAep0
WWwtIMTFFX8wg8KzfnKA0xELWSR0GAiMAkEHJdN6UCdg25UQCDweVcy/waKP
SnKWuBhj9wimnQ6bUbuN8pL5fMJn9iy9fIOqbOImY4UfiWMyKzRZu10ZVgou
RAu+yGQP6hu5RuZLZ1xoBhbEXfO7ZCIZ25z8z/DHO03SKbEBMXOWG+kjsQSg
Osa6nWfq37+asTETn/7KWuivw22B3aBLvkJ/GJt2b3IdJzclxy1hrVrcac51
TL+Fe4+lXVeSBYHybV7OQkSl8yRWFPd2jv5PGfjG6KTb19/+XdZFG0M6Wtkg
aOmR+KEq9dgBvubeZnL0SbCuMiGKPWOUJvSNsvaW7fRhvwO4+W7sOnqwqUYY
SZ/GXnMPjLD9nbA4yq4SmwodiLbuv9AmuRLi0gJsaNshNjRzi3ou78WtGEzh
sCgzydYBGD3X1rqk7+U6hgGK4HTRHbAcBJEh7vH4/tu2q4nXuE2p9Lsx9bTL
a2sH8mFgl/FfTrcxthwnXMCTpKy3H2dj6Q0nwQkpEclV3xIHlmV3lurrXlKy
8Dgiso1fWhuqGUOyESQE2qIEHROaa+hsgRy7zf5S2CIcIATOLeqbpXV7lZHh
XbEY9mZav35FwQ1DJQf14KbkYXNodWuxgKxlesdunC88tmp+D5XJBRlSYT8n
GRWCDlm17JNWAcISQFurcJgZ8pSmZ9jWSy9yjF5qJZVCp+ggMucswqkNWyCy
bdftPibAY2WOpNEt5xKf4Q1/Hnmhqm1i46Vbl/U/lTzkIK8fjkLvEkGCqkuw
RsAJpWUDxdNTf06YQBlAaJJxTxEO/tTWWrduPzcwhWrCSVn1BPc/Xnud8qQv
W9ZtJHD0U4MXzsfqMSxr1Ni26wxtjxPOVlRV3ME3EY1rpCOAZhNDGNexfHI5
cjaM9hKTcD+laYdFjSfVMRCp9VZKW/Q1Y/wFnU2NVCSni7w55+JCTskiAqeV
oK9IksVl6qJsOUpy9/rt7Deij92XYWKjLx33hJDmxKfS0gU/DO5i+d82l281
DyKgQ3gYQKxQa2yNxidcFUIrm987GR1qEf9nPxF80pqTCqMACdY2k44p9VVa
AwrAvfDL+H3xuJSZVrlKEucbTgH/fZzO985ZEV5nSlI4+wiA9snf++t4dHp1
1z3yblN+frWfRWeW8KZT+vrHGlO8SGI2ZA2U1n3JyojJ/2AFFu+Pus3HTXy5
eCRihC+L22TMQ4itcSKFhKc4TWeinS41YtPhFVmuE589Ezd0zbRzLguFgvEc
wwnXSNnKJZSCUqwTgNZQvMtGlhgN4sB0L266dwXnRrqSq7DeTM5gCet8j5NH
rEz1HYDbFsYQFW+QO7nfYFZygA9arlffztKcDIBRR8yYsPNtKdaJfgDfu6Cn
arKk544C8mjDJB6XlgtWARP5Ge+wUnOR7UQ6CRVi4ubW7P1OMGQck4tsTBsg
MjRS1Ka3hk83dyIeovIPSKIC/+iP+DQuGXLbKByCfzReT5PspxjaNwEYCLLa
XwH/ZpzaxUEUslB4+W4nms7yMjW0auYiEoXU7divZERzZ4Yc6+6Np69r+vw1
gA70CD/uicxoPP0tZrIrNO2Du73DTnI/eKIjIG07tHFTBoU4/B7EfXU8/4w6
OFyyblSTl36PMLko+OTe/NyFqYPaST1VaQ6PYfRgWjRTm6kS6jNjrfuY9Iro
TCaO+q1eZkWI+GtjBdtlWSbS4acuLgGis7DU5qWSCiKJyXGHptUzC9gn/8zg
O0QzhhH0UDkTwHkZENIrl/8kcIj3bsewsVmwJdAm4issZUPU8mXuh5RtaHsh
QP2vlImYXrJHat5mwhr3bn4VFX+CUzaQh+xGM4f1bl8dvBJ7k5MuSBaQAGEZ
nAx+YUocR06jqHNnJjIRuvx9AXN7VYH4cWYzpHpHrMbYJHsP3GSfRMJmfhYt
kg/ebqMYBzsZ4hNfuXgprPgQZ9FMNj5nybWALUilRm+flhJ1AAWvHQCsjKGM
I7QasMAQIpsaSajsfcyGCTQxzk4KAMO/P1qCqOTm8YfRTtSXUTlRl9XgBvhA
FcgQmKert5qQzapg9/Bo1lvCUMlTzKmIDQ80WXaMNRChtjjtNilrQFr+L99M
OU5T0u0B6DqimAhGLeTvL3iMg3bDeUo7p4cigYMb7eQ2GSRjZz5muTLNP8vB
0MjeXqbh8INjSUmPtFFTmRolhk1zOJSd8oh2LeoWVq+Dn95w81wYfMvdcMJL
XEuQGW3lm8iqxJFcHVonhSF+0ud8Vab9ji8ZxLzkPTY3K1vHztIePFwu3qk9
7mxN1aCUYvlgpcdKtk2KTMOCNaZvI/VtXichbgb0/+ga0+yVPSGTctGrogTj
7NkeFSn7L/BlAk07DfWL66ycf+tCDkbooDtcjLhrcaIw8JP8o9bHCHFiGmrH
26y/gCoEj/eqnPlOh9onU0ZQ4dIJS5F2ht8iDfnSrKd0ON2SU5k2U6ijuGFN
CG6VZhCaWUgAOm+BUuxbPQ/c29ZzbBETRRy1WbFBSWf7Ze9BvJpM9n5PZuC4
QJGyFw4nuRrwE98/6JY7+NWHsuRSOZmWOYmGEpMBe773Bg7LrLrsPa8xJWE3
CIR/81w2mdnXEhabYSvsGStvYt6dCLGtM8LotL5/AY4DMgRmOA03NeAq8jDR
Mls/7lKLfsSd4eOxaWpadHbekuwqpn/flVSS3QD49pLiKbripEIT//SAESLR
higdSRws9tAV+CHdpWRfb7bIRmvgrMlUgWat3rR4so7nstlI6w4TY+0wNEAD
B/1SUyzHwSezIFGmkbPhRL8KDUc3AIjgDWuRTR9i87y1DAY/GyKYoaHfTsOU
eUkoVuXeK+D1vUyHMTiEukdJoSmIClKsWnRcbvX8mWJXpC3E8FlHR/F6NOkN
4hjWJgV4oGDfZhaDFNly/zXsGpJnz5BDCLLoEU/6nY/9WWXcTrrZ8LQHNYk/
QgUNrmSBfLOz+RWfE7h0NRpGxXftI0hVZUYQk8cwQVv4LZ9U+Lrnt4A6iyYr
ajdZQaj6St4/SJ5HOudLIY6a4auhLHLhR4zfh+EHyTxRvoFB83PtAbl7qhLi
zsesf34r2JrScAJiHJS6cpkB6uAJDn8srvejyV3cFVlPuQJAMr/OKqKyMgHH
g+QRY5WZQjAWaDjMHvGw35g2SU66kyCEBZYAme7oj1CKrEhhp5QeknriUeUa
Ns+PF4SGPZUo5T46DQF7oDNQoEFH0VAElgtrrb2ocFysbDgGeGN1hxKVcJWT
e/deGkWT0GHL9lF8AQF8ot+MLFGY0LHlgiLDWHDv+udzi51ttEP1MZQP/IB0
hq6e9vRArTrTxzogLhmCYXXIDr2flsBV0F6BMA02UFgVtgKxdyG/E2vPLGI9
rqhgd4myrDoBlzehGUo2G4OYjMblr4dZYKsRAQmK294GfrCqlN56rAHwjjRQ
dWa5Qh3Pb0khq5qvRbeRZPJZt8bKV2GuVKrLnvSf4EsefYv6Ab6g4eAoG2I/
ceO5xCAel5FTFLMMWaL2RJ2v8Ia/uXttkX2BQShLXY9L8po3Y52EfrgLow6n
PEWcnU4sEc7CGXSvbf2iMlTyB9/2c06dlzMQrtvK/6BlPQ9TQ1psOBYmaRd/
FwJ8PeHUpgA3p+RBCJoShjQ2tZb2aWqPdFss/YDqB7o0A/E59Ypi/E4hC/bq
4gkOtkhyfvfKTbqvO2CEzGobZBsfTC8SsKW79J/f7YIjaSmhMka948tGUpcY
kjDWT2HxHRW4hS0s+uU4pyDmsoqlbRsuzjl9OEc8A1mgjfv00xX5X98N227A
lRXf9NaiurvmNvo0lDR4wmEvYxeZG06ypxgTs5byvcgLXSWnGuTygJS0voGF
bmhCnSL2WWVLx4exyj6wAD3uN6lBMlyFCC7+Gknf6DUZu+EJhIOSG0Jr23F2
0XmEPk9Dac/PDSaJcRdM1Qb+Zzfzv7SXGlQH6ILerZirRn9sSaUTr1HV1t7x
0P/Wgk7qT02mktp4/qhuJz3AFGliU8JhWsPeOwsGhMxcX9fyCPV2+1sH8sRZ
BAIriwxN7l6oUYYKOlsOwgl5/LtSv+hbqBoEWLM6RBt0YCTaUw2wzMlOLOIv
+CqE5diIfQ6J1q4mSB5+mej9TW0LMQQx1BStOMSPX7wUcLgesp+Rz+1Gu9oz
DR4ekxtLVfFYy4eVXD9y/DX2sB0zGBr6r8s1c+gZ/B++aqw4NN1mVlPMC/Mp
zhmpmldfDVWvfwVDQwBB8jMaqTvzPDovcgioOnbjgniHokivy3bFFFCkanj+
pZL27z9bvEUdUuYd4d4OIflEff20L757ZhLJD7Z7t206iY65dQcyNwkjhSFE
kE534t6u1ShmtZbDsWdn1JhIflYYsUqoFWn4RPg23zQGi7elDlBZ5iNOOUWS
dXxDSvISy3AqEmhcdq7h4PP7Vv3ycVrxn7B/LXcggFoKcbR+gWt5r0+D/gc1
fP2ZV4G8byblVdEGaNA3mfLYhdF7BdIOtwGzMQYsH4QcCiqyA7rmm37ey/lk
OUTAzn1De6jfe9dHWeWxPV3ObcdmSVdXPp41yAFTVYxCNoWk5ZQbWdp4C/N2
y3OQgemn6OQwMTvfB9fRizxphUfGxBMr92A1g83U9wE9jm/TaeTO4NvrLhF0
QeUKSYuFjzGXo4qPXk5122aONzrJ07RwpBQh3LRHITReY20I9GN1SHe9rcqh
ukMkgK3Fd2/82qvSEktTatXNOUY0R6EJXpQdJcVF5tTk1ZxB0iEhHQNq+HiA
diZj3HoxiOpRKk8EB4jKN3lIhrRuZ3DtEvSBMj4ibabqrED0ZnFaRwPW4+tK
GUZPNgreXcfL35Qedt6RgmcejYFk2XeduriqmKAxL9yPcOVbzrlIuIiZYenM
fS9ZK5lQmFOHgcCFT9lFm/RyQnF8TL9BXBM+f2WNQ6+BDeld6enRYW4WWK1I
blIC7CGwb5Ac9awhvHoONJDEhfP2jxcHln0fOgYGBGGKvP5FTFweE1lgu4Qg
yApOSbJ8bV6StrQVDbJP2eigfQARff2U2o4KC/9zN0XQYVW5akDNlhzvyl0z
I9flvqkFon+CtUpGaWXvlbMCQRe4qNQ7sJGMfifxsxQVyr2ri4kP8OdWjitr
xqYfA4WYbcr9Kn86Le630NLkxv7bqcgw4QWJ33IiOu7U5tux3GE3fv1aEC+U
5KVUb69IQ96mojpCvwBO6wYTAAwOtcRJxTqqhXNz/Xq8DoPOysnG7WXgPAMe
zWc0/3VLKT/zVU15+WcUSlV/bYAOW/NIeJBoZWDgev14xCQGvvXSgAgZLJvM
M/pKZ5surVhSXX1C6nDwoaziblpMAnMFai3NCb62BNFtWSeael+gc51ruM6B
isTDoPNxNxMWclUqPYf5n4CF0CJlVl8lptYLGMJ3yeUEN+zAVpRdUe/FId+F
WVPbXWqybpdmqDFh2YhZHE8gbGas7Do9Z2pEqi4AWkDBl9Dgw+KJ6Ill5RFk
hwjXaegtPZBwOklw8UFbLnZbMHSrzpETWfVm2ZQNUmbJ6+fDcdgfNY5/nMuA
RSI8wEX+6mNOqVkkaIL8IIMljpKDJzw6Etm/44p8YbWS3SYroHBNSBpUgmTz
0uAdlZp4bDzHwRiMeaMjQ7XqS4rPzNA0Ccc0trMTkcWqgj35AGuIcBEvtlLv
9nkDL8gJpDTaJdOjqSRDSJ8dhqg4o9cnr5Kle0SE0182o0v5FugfnGqwgJLT
+wiZsFNi45wNT7BnjfqIGYdrmCPLdV7oVSghgWAMYrnWQ8MGaVDzbMf0xklb
aV2cKYFxNz3DnvZ9ereu9v47yYZKj6WBNyzr0pH/g+cBNR2hA8Yp9HMboUDd
rbGZ/bzCTi7RO76bSmccZZS85Hb+zW16uASqHtWuwEoZRnyjwpfXeDTb74dL
vxWdEZTmvMRRuUZNAma8yTw3+wm37PdBrVrDGI+fhjUI0XiHsHHr1fbYoQYC
cD2CMuf1zf+1vunfJL+xk7b3MEFZFAdoliW7SazQsNQfJmXcHcIWcruaV1Ds
3wwyCs+dsLgVJy4vdEqdwHLLMSCYsJtDHV1rkqve1Tm9UDvP8qaCB+EkfmEo
OY0C0squhPocRlnqCUzybDXTsMsPiIhVeErFJAKZVPozgteBm3pOqOGguDYi
tk/EocoFoVUnPAcMp4v4+sOK0/d03n+oklFdlklT8DxKifqyTeaEbPM0fhMQ
2akqgYmDeZwRcAjqyJBmPss0WPn0A+EMkEp74rLTF/ta2b6aXaddgM9UV7Rl
K8f/KhNMBUP3vdynfJKBCXThOObCykWVbv5VKowzO0BSAfoHtuqIkBDcLZE1
1SBPcq0gH0UcPTfI+8zIHu+QuCKRvvuw5+J82M3J7gEDG2Zi8g2/iQ0gBGXr
aBkEEiXBBH7VGGBPWKe6r+XHlObaLFlJHNhnRSKSoUnc9E8zvukSJQ4NihtE
Bxvi/0eVLyTAomDcX5Jm/976ZudjBHjuApOkUQ0O2iLOGxEiFaXL6MjpUI4j
+coh6Wwy9Uc4CpEIr0lvUpzSwFoPHNotJLy5S/FPuO+uxHqJicxfAjUTUwC3
G5bN0D9jqalnk4R/Z1aylp37lvnsgfjaD2fImQrYSHLhfPyDq/2FoNxAMnXp
GhCroxAI2pzL9H36NH7fLGN5tm5OQP/SRynN7VbMFW9F8/K4DQra84/1d+Iu
tvPKSHIt75BdhS0TCl1TQlbshO5y0KQ2KGXIpFu/twK47y6sA3zcgJOTlxtO
dVtnpxsgaZwhNeBwIwHdbgX0U50oTDPUUZjkmpkeD0bMnzLM+99UW0WA0Bqp
PLLogUEXf5Igual9piQaW3uwv0z0KjMYV1HOjy1OcUdM/gH5J75X26I3rwvH
y8/QPf+5im/cRSgPWuo5TDNBokfdzlqEkNeP5uXa758WpROkbrxowH+VQ75m
upKB1YjcdsnpYJSISQKm/7HrN78T4K0P5rKmInmctZF5ORSIADZtgm90IXhG
lbOHVK+yNJc7PhiFGs5jp4HnWdccts8DDNac07IXnYy4p8StWNeh4I0ocNWk
aaozbIL2iPjBn/yfc3lNBXeZ0taAWjyFj5PxNk/P9tB9DPMCUQvsHtfAW83i
TohRKkOI0vm3RhmzaFsX57ozBaTXkxsCLTGeyvyDoDcx65onsdsJ+cWbAxRm
aJmoSPoSkUoHSSobDQzCugJX+eYFkvKURCkmB/qeSwiUPc8uzjKeLDVx/8+O
ao2+PvXghJsfkV59838OiedCjJ2RCpbtCK7qkpSuym1Z4MbQ4lWFHQRmRy8e
0SolkkRk175PsSiJwVhiZBjcH1Qwjq16ovCNWgfIW/o/espqwHVzvXNSHZ2D
3k8er/SOYWUZmJkGXMqfdCGaC6hBRqZz8pqA1fmMcyGpe++uWJM+52M5XXgu
ZfRP7N9jOV4UBhr/YDq5+SqR7wRCGoe1tpxXzjUIs5U74ejHjAOAtu9GXw4P
f2onNKkm1f9nc48qt1Mw+Qhb0piESyz9oJKMn0QrwnBTXgwRzMmoyABsivxC
3XSSsWMrHcCTEIMRAwiGK509bBcfgMFzOyZeYtxZO/XBDd4aQbNWkuiZev+w
mbcBNbJnV/kxR+J3ZFZUuXPuiJJ41NUKWObjY81fs3TLk4GnQMPJZXV/9svE
5kHnTTS327rw/v4eqH3fzujvN5P2PnBUV5sNpRDUzwm3soLwyWQU9nXPfsJn
FEyojfRX+olPZ5IkbUs3TeZgDciQOwt06N8i3uj0UtSytZZV92taeDOXf5j+
O+TxOBD5QPQ9q97qfYrQEmQOLAGMgDnoUMJQB29AZpVQV0UYMZkxHlsSYUhd
JhbXUJd+2BD2hXwDgrutBPAix1fHvASDAMs5DhvoZa+zim+QZI8O87HK1dtY
J1amq0MAcjgwqJ/xvbPOiuZ7edCJQ6Bb6NpNHUMGL8kqJpvSrrfjD/d2t9lx
bhMl/DqHIQrNJ8tcvDgOljXgDaEMEEgQY2CG1EpyruT3otHh7gnxK7MXk0ne
xQUdqO22P9QODT9jnvyUz1th1VllrIi/wij0Q2AQgVDO9VZYZgLJLgPhWxL6
5T8ccalVEa3hqfDIYVXQ0Stof+ecAv+qvRg1VO8ZYg+Qal5Xr3G1Dr5JJpWW
uGhzQLWeCs89azle0y3ksmewuIjwKxbQbSZA5LX6u+qZh67ir0XITousyiWQ
F9pjqcscn4FI1POqk9tjx/i3toX/USo2fZIe3o4AiTsiONWMojucoOJ1U00Q
f4PLvgZZfyUBa+4wvVd6QILFmDUbK0dvwLG6hr2QAd7YSLNHzo+YkTOtkmJR
pcrVWohh9LARdcr49a9e6dPClNZhQeNMuN6ZsF3RnHHxM5pL6P8aT2gC2RJ4
YJy7IsSAbXO0ArY8xzA5PSDTe56EUd3Hb70chVO5Pyvy7FGMr5SODh/s60yi
bjJ6XLmTaXGx4x3QVrjumxrkr7PQCmoQf7hUFIVEFsZH7IFZMJf4jp1wBlQe
Ms6YDSW2PD5QLh3N21ul7r3e+GAXIZZDPOYjwKhw/c56FwVf6GIfjPEJGv+O
WAdd9JG1yAjwKM5yDQpN/6EHYQSzJH7OCZZKhmcDnb/vau4ea1YYRuWOOAip
EtyxHxhdNRn9oXgt1wgqEjsNy20OPnTqOXV4bPextIp8uaMMqTGKyrtDOvoC
puRqMOL2S9QLMkIOLTGqUeIoXfdAipifVCSi/FUuPkS5lcyyuWiYMqAVl0PU
NtfxaXWXy1UMVsR0fxcIRONg3C+IcLFxowAnGDPj0AEDJo1peqMv1TmHrSdS
HIIWGookfngMOZeqQYe3TAqbCfIqg1Wb2c4Cwb7NN44/1TiM9nQhZg2j+FsX
8y2sxpYNZEF6ekdKJfO9afIxaIIulqgG2E/acS8I7jggisx0KOENOxQ0oadZ
jzyaOhobZFnz+uTKCsQU7tbVERYtC7E+LEXR5ZTZ0PfeZZujUhPxjCpkB+Ho
mJQbobeh5FALy9OIX+HSCL2yDB98HII9Z2Uk8qnQcwZqnQOJ8JcrPmgYAYRq
R9/sBkxCdvpXZdlL1P/Fbaf5iwHC/et3Jsmd94kN/JxvOgZnhbFaQj5TrGUi
6tR3d/ljA90CxGsc0/b26SUDs70we0E3IvrzMGXcay2xHD3ULOXSD9C1bIAY
F9VtdVMCxvfKV0VENj21sAg25GwR60+sjsXW6By7jeHIEKvfWSeiVuwUi2SU
s7hv8zH6pEKcqfDVBR1lAfaBs4QFxOX7h6ODdgHQCu9V14MXPM/B7HE6M4Fv
VPxr4pbplq1xjM1oQFJjO54oTLaWIUe51rCLth7mwMJoTaK67Lo3nU7UxxS0
f+vPZGHjdtiOhQSs3LvbuD2A6v89MyBnAmR/XOFMVBvlodO4tccjpz4JD9Ma
7H6lp4vQJVYZZYzD0JiCIcpSOhwr+Vob4j6JhTb4mEx/jFcg/WA+45jYUJZG
0FgcfyCzf3TFsB+ULoe92qupDJwWaRtTMaHC9fxenx9sg0K9cw7V053Nufxe
Hmm8Y6xKovEA0xOoHslssH2Sl6maxc7NLTAzqaJ4fyDNWGuz3U/HXMlhRtpd
10Zj620JMmVKrSANMtTb2s1Bl13C2ij+Q8Wdj7vvHa1vx6bK2gkLwF8mr29H
HwRN0HMLNfiUiY55aMl6awQif/FoRyueZjWf9zpdjejvHMuAKHXqQVoPNh18
me9+volhtk0w/If1ykIYelMtetbJ26VMJnBFLFrcrHxY2otKd1JXeVbThoik
OpwCbcpJBEl9z90XxEWGxZAMweOVAiRqDKdw9V0kQqh5LJIG+o5a3xJu+FjM
+fpGZfce56VXn5+nLD4hHhfp2VwAd59gebY+alK/CRZULxajPHH+rWF55DaN
s5hVbn+uC54yslLv65QYIGhJVzw5tIabhLg3iRS5Z3/WXCuIJ/GJGB6lK5IK
yWd/WoQ4xxq53ORLo6fA4GTBtcjKG6U4kihlZb519W5CLq5kuKG/xARoQKrz
3VKygoUWAc7FMzveCCUzw3Fy0u4JwILtDenOTh+l692ui6gYbH43TVEAhEsU
phfzI1qAUr9GjSawmoYcAmO8JYX/5qDYArqD3+q+F7br0isvgoh0E4gCb5iD
brjNnuC1rfnn6OqLX+aV5B5ofTmT67Qp0N6OM6JAtNi5QfgI/s5uU3s2PDiT
ysMAdrqqMKv0r1wmGzW347QlaKhoXAY1BliY0HTNaS+T89c3MU6gl0+p/XOs
Ga4qywuzi/X/Th/zZ00F5OOoDJZ7zOJYYLXWEArj/3/W/GGGgj6AR0DAizLO
7oGLaB2kFUEOLf/HQWpdxCADi7t/ZLTTCRRpBGRCXkKxhXRUC/XSFPzFzu2Q
9CstfvHfD//Z8Xj/MIKpPUrncWeEV4EIfharB44tEH7+7lMz5N9rOigrOaRi
a5TE1E/NFfq06r3B/t9OV5VOS5v39Opms/ik0ClQTD9BgOTHqPSoREli33ni
5BP/XEjVyyJdfVxLYgJDZFnpmj8pxJ0k5YAQF7Y+SvyBqQk3l1SN889LgITU
yjSbx5RCsljfF5sPwe5Oiran2Vhos9KKjm22UPdxLAVVPCHsv3/Sbg+6OKQN
hj9DaofwYHVpueLhFCAJ+UcNpnvNjx4bVgMW0JP2GrPwxnrfPGugdiaV8gvd
2EQvhNAE5J7okYZPe4eTLqaARvDq82YDK+iXU/rPAM+8jYVexDPQEC51fx/s
rqt/v46PJb9R+mjO+j0xzzVb5NTZNC17Dp9RpQdjq2hxt18Wz9tHLe8V8Ari
2j1d5qE442Na4nGnOrmIVl2zPEvqzOQL24733F3sjOJ9RQlL/ukz4RQnRz9W
Mmg3wzsw5SJwohuuPOsaTYWJp9eFMChHuRS6cqCPIDCGoFtTR39Q0kkU1i89
kUdqSsWy8cgBG6d3Krf3VoXnnWNHkiiZMEG9+C1wX1vZMlWs6ni3udUjnXas
ezGtTLp2mavtxEjFo8ul88t6a5PPmgoID7OwjSRS8EZyt9/ETbejbYMnXq0Q
kpLvGpqV1hF1CeWuvLw2+s2k18UE5bJs6Lj9mD4Bzo6NU+butQ2A6y3fXHOc
clVGTz8t5w2wDMwL+HdSqQfpv7HCHQALFXeRspp0A0GOS5OeQMa6JX4f6Hl3
jaKlpQYnpO+UMQwabHTqcwt0C/jbbX+bch9DMyO8OWUo34msZe8W9YlNezK6
EcKSNHdPae96o3yuEUUz8J9sSOAcL7f7g7AZ1CZNwFGbZqDUWgl9lyGwx3de
DDlnIGJfGDxxGLJXlyb8vFQ7wvYDBWLW809dnpMXJEi+B6gSnK4tx1A/iAMA
ENMKyeAw2WEpNmlm7e4GdzqkY7opAjivRgbZ0OL8vTFROG85+L14GSUPRWDp
XXttnpaf+/VVoiN96SK3Oq2YihTIRovpMC+nfQQuCQr0nuO8enQB7tQMdMkA
WujdQQDidNDscCljB3H15LQFgFfDSHEZCK8Zb41pbo/nM+As3dCrvFf5koFn
rbvZ3Mq7U8f0vEqjXMZkZYPA/9eRjmhvQhyutTTVNC5fQNDLWuvVQVu9XrMU
3ZnvZG1ISEVoduSLXfVEFRsLkSXHsm8sITf5C+jAfHslvPXdRm4l5xz5+YF1
4mRNhlvHqBxISrgoAYhnw3mMXwCGfqwnbxY3TwKYnCqFaO2R/S33mHRXy0MJ
eVbkGfH3+XBzxiRPjDthOS17Q5XGgx3OoNfzRa/39+La43r/p6vY0HCOeqFi
07K20sABsZc12hn+koVDHPuzDCzIKLDJ0uScWz7O3Ch6Ig9SHNlY+kpNE9DR
cPVQOiBXBnOIde4j8GeXzQLuLUORzZb0kK6Aw7yax2mOAsyaECEDoia6YT80
yo3XhHzito0bPtStHd9EnW6qaMutZ1vFGR4BM0eGvpZ6y41J3flAMtesyhX6
WoxSbaaMbRj+TjigdHSfFixIytRV9Zc24BVQWnsypZCxWa4hAAjSMXEdDjrk
6gJgdgawsCAOzfhqvu7dtJ9gVm8tLsuiIPAW/cjzt3nxNXvuUXA2zbPDzs4C
m5tkTf6bLznHgc0j0uQ/WS3czLqxX3INFqzjOWec+Shv0XsK0fyM52VyvDMY
4Aj0Hswb4T59Epw+4vD+6sJqTRCAuxg25AuXtZEjN1YjOIs5NPfzbCn8E3r9
S5Nn25MSyjEwTFsemV/rNh2mhuW6uY2BZEMfmlhkJX03LhDON3xRqQY1W6Qi
5ySOgrpWx9WRYmSsMjC5GkOfeKzsVLR5dlBfmqH1w8DdcBJd510zS6gmXV8/
nyB6kEgmKxZ+rBeNOJYZ/b2KnyWQxAHEYktDkO7iKrzLoLEONNENAH8mwtvi
Jyy3CqemSAMuBFwtQmkFctx3+KHv6qU9CSRGswYfiQV2AdEeL0mpHU73bYLa
kLr/rSrb6wDD7Xh9L0ARRBKxgiUnn58HYYTiqW3Il6aSXwsvSBYSXrubWut1
yPlSr2RDiIed/sMYYe5ZMy/I6d3lRkkWzxtfr/o7y/mznFZsEGKXgbB/TwSy
zcF7Vq5Dmr7xmZ+RwLs/CXMMED7YZgzwSxebEefa0p82gD7yUlWDNGDfFFAl
P6n9huCzMBgqM/YfwgQfxDVEezOV+n4wkH25LVD509Ja/9pfW4akCkNBHLd0
8xrQ0Xjnj99Rh/mpNTderQdHPkdYUSdqgskAi1BOxW4xdbV95AsWeyDFfLvb
uOJt7F9ORzBUXHBejIni34JnLxK9MmYUzZ317hlNtK35/n2bmtDnNk6JeT6G
fnUKtJarAkzZ5ZG1W/gJqYb5I0VnX6jGvLFsipiAPRx1gZuH8dLOndW/bv/H
73R6TGhg8G/TEACwsGnT4+AqbPJ09aq3KSbmNd73mD0FTe0srOCu6ywCYdtW
DYHtn32HxNX1LYn2aVT6r/ZOSeFoLD/yZe77ipi9JlrYt+J/EnrutT4ERKuS
kLPGUoXDkJlXBctdORyhXVIA0dJLPMrVkeKKSJndi6rq8w0p026+aV+EVkvs
bODT06afyjh+l0PqcPgbX0RU0H1t28gvmHwmgg9AwDtPn+HMvRygof/aROBk
nGljO2p0n+jgQjKBpRVpYlFGJPj08pWnpjCXIc+ruJQT3XRBIy7pB65gjnS0
bzL0Wuzi/8tQaMhE7Kiv3rSIZZDusHBEO6IpQvryDIgFdMQ4WUvcQwH10pDw
3n59j13AlyG1jWyrld4ChKMu0flS8k6nel0lZk21pDk3whn29PEuME8cYukf
fX5/soNPqkbi6axqiQ2Kb2C1ZEb4RRCh3R3tFsMnB/Njak+IDucfxrR0EIwP
0aHY/gMSvfMc155WFcoqWi8EcUM2uqXOQfXfIz6xW3Iwh4JDVlfGDretZJvn
hzHbrTFqPb72wwrXA4Qw3wHvHCx9pK92WBgKYuRXNCVF4UKx6IanRee7YXze
63Cfn5g8YRlfqsbd13PpDIoCrcGLJ3sKAeAL0c0OL+G+sxBcflWSVECFAaVo
jmPdNTyYTkk6Pu+DMKnXfozNjDkMOycgy+T1aUkXE+s4yRsjJ7G0qOeDQ+Qh
y35mm/777cFCpnhCjrNqsysh9DtiHU+38C7QRYBS9zX3HEsLR9kb3Vb6EN9W
cVVIyuA4Ed+r0FxhfAn/pGMiy3xTaWx3rM3eQ1Ij2TfE9nvrsbtBYnJnYrBy
1gy9qsg6G3//UZsm029LkC5G+75bmU/Sr0o/L4aanvaQLxfmMOLMAbVuPCiv
jDOj3UadyFc4hDzUPbl87MVVEFsUA3JNzWJK7ldu+3FQ0K/xGJ3NI9x2/DsY
Uhx3sSorZT0qcjQPX/iwEYAYuFGKEF7lpjyVMANBbFTF/V0W1Zh2Ek/uAWp8
elgAmcndHk0e9n+EoZ72LHztlWFGen3BUT6yzZL2sCxzxyNkoedRSgGnYAZX
TDA721vN9ToFd/85w9zG106/NMjtbjsy2WXoA45rHsZ7vRcd7bRkzDG6Xyff
eJRyHahdje1/Gfft3a/JT8/O30N4/fG98MVEZkZ1WVOo4Ihaj0duWd3fRern
UWoEEX45tLEfvvcVAymjzhmSjzktRexXZxGcPDdvPRycm2vrI1icRmsidhgA
tXy7ce8dHHByE2tfYgxs4LpepooPxZh1sJR+snJqvPKKCVCSY8UhryUkwoYW
8oifn3No5vCqXdG22dPpV9lsuUtgeHdfw7Jpa+Vpf654pKJiVT4vz+oteHzE
AuKTOeGxtBdc5HLXCc54RPBdjS7BOPetqWAciyeTo81dDws0jchwzC+2aQmH
tqv/pvluh3g50sDXYBxPf3+L4KEpZNU0G0Xv7wrB7NbxKWqLvaetyV5Uyc7O
j4JCjAkBOwITDN2sYhHlfdRQGt5vJ63mgmIq6hRgFAN40xgnZ2sLHzVrU5zJ
C/gvGfw+SXDmPcX6kkq3mlJtb7ZvmIto4Xae7viD1XXLCbsdCGQeSAlbRek9
coJdHwsPderDTnAlmTRAZBZICNviSeStH0COYoGp3ITnT//RSG2UpNodMXnu
tM26znws+1p55XR2qdex1NtQQr570ehw+msmw4Vgh/25alB2/W9hrZKfZ0VP
5QIdJpVMgnc2Z98OH3SH/rMFgOxkh5oB1qC2YruN4sLmwTWLsT4hy3igOgL4
WHeMWdlSwW3+8swLuEAL2Fm144BTHQb+if61vx8Shu53EORiVqbDAoyFB7un
CUnFmdMkEOwqHUqkKlEXR2s1tJcpfisuv+od6eHBWlH2Mh/INOQjeTv+VvyY
aNeEhDOOk8FgsM8mTutzCRav3hndCujOPG71yATvb/7L1ea4l9v0GklUEQkY
dPWAeTcbgIIm1LA825W4jlIYTtkCs738V2imh+0aiYFvxJmw4aH+lU+TCBkY
sX7iJetRtJoknCmbuo8RSds7QuiCO+DtIkdA+720hD2mmLhsvA+owGr892nA
0HYyoeJosIkdWAJ0ewUUAhxUbLKmbW9bVQQvF7sl/94aq8WbbPhCipv4qz/r
czM5wBv9hYfeHrdPQ7U9oYpANnm3eXHgSl41mcrdZp4ldokPlSj3WTlEnsmO
8tjh66ajIkDSCEAzUW86Q6dBLLVtg5LJKDHt0jzLTxpR6DZ54w0gMPu04ra9
sarKUrnQiu1b1zESJYes/DsBxPwCkCL3r6t8104o698k/fXoraIpjtEjmnoE
dQXAsayFX+gWyRMAWQwe8m5DDmZEpEqDGaABwDoPhZ9Q3iIQ0Gz7W6lxkj0L
ueK8QE4gaARRg8G5TINhArHloZ+AE/FHxDbzaYYQwwEmpLQnR7uDh+hgkf5n
VdKTyAaLJRpuoJa0UOFPk0Vq/k48Wx2Pm0n1WL/CqGVVU7uKtxSlLrmPC83j
QrXj06P8RnJGzvsdSvIGS7sKBo0RbGOaufp7TSDrMK1kuJ9bf7D6qkbqT0SF
T+R89bIz9ZTsVVfnxEBhMqYGgygKf4MwsyIyb85qKJEqkbzxRYTjutmvuPRw
oPLRalLiuEDpSRiRVTW6msCU2xaxvIk3fSvnZoJlmL8oBn1oZHXczhHorfz1
d1YelrCdEvSQeTpHNDPjr59LuN97QmiILnB1eYizjTzWzyjkQSIZMhxcx8ID
PhOTdSmccvOmHz2J4tQy5y8f7f0kMnLUQqL54HUcAqVE33VBQvvljlrrTh7G
i5YqQ8DaEk0D0oEFq7bP9nKH7cCuZVEgLfjYRBqLMugw1dvdLEVbtVFAW/3N
fONdeYuNct/MLbGYpPNYpGZOXkQqOucW1kzYo1iPn4H3jo5BHBCyeYz1xQTr
np+iS0ZP6RCuCH+jxQriYw/+P1SsVx+9K5Ow16r4eyo+xqjRPYcw9YM4qeCq
A7v22xaH/1gHRibpiD09cigjhekDCEpsNCQ2CbpZUaELVkhvbrYEYTTHWj2n
wlFGWlPGeERR3z7FTpZI0FYAupvclAo5Qypi5XlvrghVab0Iny/sl/Opwby+
DvhC1OFBzq0Zg6YWhsbOTuA8ABSBquZEt6zh2f6dq2n7dp0guEGkA6k9JA82
V9oy3jIyej8Bki28plFZ5plKzYWgszlHupCjYMgh4WE55lSjPXL5IbUS+avp
EQawy0mea77H222JWTHSPL1uVdNjVbYYSdCmwke4+tjGTJ2us0aN2sBWSpNK
S8ghtg6UcPTnGIPCF37hF0Gwt7ZqPw63dAULK6zOomIme4pZZz/p8std2N2O
EIkPghCXscdg1yhKhvRCuSoVkAWzrjXfigLqjFhClvH5x66dGRCHRNaJPMFS
ayYyp+qC9/K9BI2l07KyC7KwCRv+ONnvf8zglUpHNhZFgj6dWFvnaeqvFYIv
fKcjNamDT6yM1pACAVnq9Y5wWLTrOodMo/9QtTnkSDQBXILFzE/EGSiR5o0L
T8OqbH2tyZxEvr9YlqsqPnbKl+rEKL3luAa36unn7Prs4n1QrY+e0Xo3bZ0+
/nV4w6rrUugz14yjHq+2EFbAHJ6KB+GxQEA2yf3jo324VmvrFA6MEMswcxn2
q4SucfdnanIu6RCcAolC/e2KcCO9tjnjjytZJyrP4VxHBxEezXLSUoVdPwON
g6q5KKuDjcMGyUcnvJXANzOJ+JJXEoFgoa3kNdd5cgOZTnKCN7g7CkvfAlvY
6kWbi1XITSJR9P1p0lgPnKmDBb3p5FhlQAwYKugyMMmJpY11v6iMcxAfQINf
IPHLiiN1O19DRaS6LBjAXhdO7qqjK7msPYGTSIYUN0Xm8RMdOSZKotVSIHb0
Ph0imtRkzyBeCHFghXOPL7N/S41OYDneOMWtOp1MsQNJUUzRTareHwAuKXyg
xXSNeHK6L/EpgiVxVlhgCh0JE3aH6Mqn43A6TbUn1xNaM8U8d2HI8POuyxWE
MySaLSlts1vhaRCkBbD1Jy9XocJbZO8pgYKuHirkL7L7AhqdUHqCGhHE3qvd
HFPrM0rfyqF7crWNw91gdf1gMN4Sd/iACURYrtiq695A3AlGlf+ueu94q7T6
bzFgZ4Zr8Oc1DaXwHeU7LaBLGu5Odg+KN6eD27kPShZKiPxI2I6ukixgWpRJ
n9wzLoFHPZOZOCiKzKJkhPr+1Crz26xNfoyRHJXJPTrT+QVCV4R82zk7F/EK
YC5oWQc8BgSUWmQt+9+066hEVObXdcxzBE1A8IwMeKHquj8XujSVJKoZu7d4
i6uyWxNKMkov+DS/qP+A3UZqgTK6Z5tiA+OkAY6zrovyytBN7gmcev8O0VTl
DyM2mj6bf+2AGDk3IB/f6/FuIR1TXgReAFEVGeH7LcfLdIh4V5tOPlLSxgem
CIkoW4FIYxHQjVDpoMiR0pUa72sy0UykJCM5VHq/0ysmLO3hT7bu90gAdDff
NGv8OjZYk1kifmT9HTyxyWNbDWP+shEFsoaQGT/cI24I0sVy6XoLbZdKThXJ
ZMKI6hFmMCIj+C93FIZTHbwpch13dIrQmxXwYM1DKjUpaNUzsvhvzl4NTp0g
kl3IijkhpbVNW7xoTGsRuTLBDtECOh8Qyd572TPNCgTL5aiJdJdWJwQHn9ZY
D/c/ZD/tnsHrO+/Vz2WLYJn6xseHPYkDy3QhqNgr2gNoh/zZ0uRflmw/zdj7
BM6ckVAuKMtKDyHiWRSpM0qtd5FZ/gNvE6fO7sVVTvYU1RbwsElxCEvr93cC
veK2AhxOH3msXiE0ksS8I9wpzUEN2520XRYzbniBM+0tWNfCpa8eOvfuYk7y
1htWKkZVPV0Qv/gDtzA0tyHl4cdveqgRkuxvwbb1qwxJsbXSTE1rc3VmqBzI
lkm4NdxSfRUNM5/gN8gQ0FZ383SOTFusGb0HfZcEkNTDv6/y6cUj54B1gSjU
cH1L7UwKQqy4IJ0ffQ9xL3sVzRS+atms06vsSvs3bv2Yta7s4xYbc43aHBoo
rFA4iRnvWt3Q4u1/sz2wSGRp8/8d0qmQQUA0qak1RULk6Hybtpm3evrHenIr
D/gCZajw0uXJHO9ca5rQIgSbQ0W0/ljiDc7fjyGYsR6k0ajlXUmgvROVp6Od
z0ozaU6ohDFPJtkJebMlE2bQ997Y1tsqaR2HoASKOZANQUZfbYoJO9FSz5Ix
LyFRHkyk8SJSGlPNdbaD1uODxts3OmUn+QLCulq1TeZOj3gXmySe0TGNFxQ8
ZaMjXZlPkK17IvQpmlWYIxbkOIO7Ve9Wm/FJzhKw5FE+eutn5QH44pKkX7pl
NLKNbxaCfEs7dGk7kGyabz7PgJ+edSVLOhSaFzOz+1yhWnJIilDzh8V7okNR
TU7FVLso/Sg1HW/9uSKREARg8L4AeQAghPeLEWLr7B+rmeePmlBFRWrZzszU
XR3an6GeD9ONMB3LJvvpnjH0rpVciGPD8K7UJRHAF8AKuVLfKyqZxYxVtUUZ
1fWCT0IYFGr70gDsFXLVOYbVjjg2vqWH8QkukWfNMxlZksfBHisa/7eVRqEg
lve62AEVxunFdTA71JfLvAi1CbidMu6Z8JiK1cMyTPg24Hwr5uuHVbXnxPu3
ohinLyo+1kM2MgPNtVVJjQGj7VPfq0Qm3qX08UMWUizpWChZVzp1tOoMqD65
5MHPYgWhj8VeKnZmUH84oWmmPPCiWA/Wx2iN6RaWQTu5FpqD/3cvw/DmqgaN
WhAFkEUrV2DzQoigBwlNN8FpWmgcBFofG5yRxFDNcIw9NhUG21XUWn4umUAr
J1QuOOY54C7F4byzpl3rhsa5vJTr9Sh71oVB2QPStJpOnx9db/XHS9MbpTx3
gTaQ/Vku9Ndvcds/GJpBo9fzxZRqboepz9K9y7+gZVALG/aITCXIEcYOP3KZ
Hgf6NMFqy1LDLzQ4m6Ckcf2/MKTScyuo2pwk8xLHkvIurVh6jjZWix07rLGh
OlUMNC7sCtCMhPP0Xzkzu9DxLElsCgW6Vrl716u3vOV0EwpDtKcA9vvDr+A9
s+hASWENO1JSQxitkKB42AVGvm7+TQqUnzlLoZ4uBl9ZhTb0gfxXS9pZOpNM
E8uC4bu7Tj3cJNmfy4bmLk42hSk/Ksq6kUbhgFaqVUNysRV8TY3PcB3lBWmz
zdM3OIZuB7LUHIRoOKLN5VeYbui/GYz6GE3U9dflqU05O5xNzn5ahkjoYBDn
TisZswhpxHdwFnDLQLEpOz84V6yRnHQ1xjSUIGLknC1/csUbw9uttF14ky1/
//2N0F8j3ccI/G/rk5sD9ntVPv1+Yam2faaxoP3e/xRGP6OlYRUBZI01wtAj
nXn+VzjdY28FDKEZMDnlHmqS5wXxecXn6fiinYooOv2AjAFA6FM2efi9T6FA
h6FwoU1zX2ofIOO2g2bv5LHIK6U85Wc2ktQd5h+97mhV3epin1PXUzR8lCQd
GqRhQketyolY5bZlCZ1WJSbVF2PxCh8Vm5o2muucc5DXRaZEBZyCGvho2/vY
/5ki/5Gz9qDRczj/fDvdBSCafL2z0cXElzDQ1BuqrTGBjqdGWI4UppKBWR9R
uwbGh7a6KgNt3eSYuXRl8h/DMtRefIGo37CUwRV9icHK+xQytV/fj17+Qc5g
FPD/jetE/aw6qzCZdXiDlYSbNtziJ6YGjrCDy2F0lsB0BghlWY3ekaRXFM5m
J7kuIxSwEEiIL3xA6vWlP0oUDMwpFTG5Vl5+L8UjkGodwGzavdSk+dMA8uLF
9YM0YErfJDYC5hDM+SPOVjpABkLyzUGofvVeMe73A6ZG6W4vGfma4yh+P6fH
JU24kbXaEskS6wFL3Pv+5ySTrc6XERaGkJCwmnpA4ByAcDMayyOo0u0nPoQV
tR690mfewJroAfoMbl25gKb1c7YwidoC/WA1yuk1Yi2CqNggFeqIyjNnq1EY
hVEpuDfAdsKbievoM22HHqE+LaD5JMA1EYOHjyLrbNmQq2LBN/t/VQYeVAZ0
uM/ePjPhk6gz09reyDtgz4tyu442btoH1ERH1WfqUIMHzLPic+6ZepifSJI2
Ok4cJZje4ehrTakeG7WXSRMYdSvbHn1MOgfi9M+A8n/G6TcVwugY3Y/rLpbb
oXBzSbnfhhSYGbVgDc3VACL3bIG89mAKc54qPj00XmJW9ZzcK+sRfPFXOd8C
4KISAnmulJvjTSQAGPK4IZ9aC/Gjgglje2gx2keX44w89sBZmV0trV165BAU
egpHMprFSvkx5d1WOXnJvqPdoQg0mdZNBk/y8u2QOBZgiRYaIgcJqdH40/Dd
ytiCVEpGmsH88YfPNqE4wbuwHNE+hNSmYrqHWHxPgC3GTfHg8YdyqO7pOjA0
XVnvTR07BD/K1qCvy0JXe1yJJJ22v+GQ9/Rv7NNodTr7SghNMTaiRtxSTdiW
rPIwn/s9drYhVG9BF12M1WNCXh3+PMiW+KUge9CmagPIURnjyt3sQcd+wGZB
lFNtcv8b4xepzTouov8V0tFNXmTkbka4cLxuBu0vI5Uzkd5M2iKBrO3JDm4u
3Y0nn1ueBn8kjBboWEUkriF0MBeW3VWY1n83QzDWJmVEwA8eZNrjSSdmx3f3
s+PIP1uK6dvIpaQzlPRvVGr+f2WMQ/1OKR+xOdMnG/2vPQ2y6ZTmAWqyzAiZ
gdwIkaxk4CFV171zQCJ5uYOJ1+UVjbYkNIZc+Gg1LbY4sAlzbXNIKpwYjH9k
ruouh+ETKwC9lE+SXWamKR5hWUT6om1xbUO0KK3Qqh/mjtHxooytMKeGbZs2
3MwQ0g0Cl5kq1V+1K3CjiKMx0IwjKr62He66ZwA/Uq7XMVY92yGbahZh9Ac9
jr/k+lSv7b+onJc3D1tbZUjxsv9cz+xzq9PRwS3pZb3h1b7ds0EuO8vz5RXK
v1ReDc0/S3XAzQdlkgzb3QJD02oFDudy9Ysz3Ent5thjZD4Y7FlvL+DBfyPz
ESIXcBXPIUtIqBU1uhObAUJwpM1xW3mQNJ/+qKfMKP7nrEtlEtrdQg4XYJHP
rwjUW9XSZxRloJbxQar36NUo4YwAa8qhlbydB3afivU8l7nZqZzIkgYeqD1B
gPg5A+0NqYWfH1DPaxIuLI0BqO6qh7hXlbXwUizQxp0CJ5lKKOQfaq8syy3j
hLD9Db4LLG+azfgX3Dg0UHd5nwvuq5NEr5TGAErkhDYByx4OhbW29+yd7GTJ
6/Uqzv+PDuUxA81/BuZpaol4lslk/2WlmIdimvSyu+LcKosx7FWy5W6Dm/YV
vRvbWxdAV373cWayFBzklVuL+/4XAD3RBn8AtU33qFJm24eKOCJ2LmJqCZnA
OdB71P+nVLqm+g966pjVzlqWh44R6lrCPD56P348+0axmS6FcDtPp0GaRK5F
LW50d45XOn49ViWxHS+t2pPwIPlRHScYhNquRrS6hFWKV3HaTo8U9maufRmj
eF8Yb+EJ0MOfAyEd1D9rkiWa7RCdl9p5CO2JMaiQizdoPNVvZ4zZaReW711l
sWk8fFrH+2vwoB2BA0uaAf200geFk6tnXMUuyZBgw2GjzoRUAffmmm0NGymn
nhAUMg0P1NlRdkQxAZQUiWuIk0jKMl3Tquk1ecX5QReZg1quGfWkLgGSRtU6
7Te8yJtdpAva/TkLXnSKhHYVrfbQKE9MD8gQwD51D8aY531N7SvuxJNKyw5a
yPW1FNjzml0Tl9+8BYLcDJas85OTn6K1vXUM+mqVcNNurOyGcKvQy8s4LOCx
D40Q5i2mlarEFQ7k/Vtfz960fmInfP+xQIarkXhSebasWi32gdcJ/XsZuAnK
ypHAKFUaT1XZMbTWsZ5WJQvcgM4Nb/eQWJZScuVGkMKOQvU+tmr0FyNvyCYa
6pvq8SMGCL+dXRTCu5HBQwpRuAPG1EiSRM5dM8mFPvwF+VxZGV1QUOb10ZWO
rVT4Lvh2r6OCzpE1yCtCWq56SBPfAzbFcFCViFgin2vGb3VP8IxOiTV891Ks
Wi/96OLasaWcxPq/BnYdV35tsX7JN/UuRBJfIp72UpQoYrwAfH8RL/hI1I5f
Rx1uDZpUlZbbaKIqQetmFeY8eZKLwUbwnEiiejBaF7Ay82hMNBr9MXURtQMS
PtsRASgss2kqEG/MDSrfTc3DHSaE12L0vLc7eXFRArcImzWA/lMzlZspUoHF
CWBU1w9CqIiuc/bVsuAbUglJrvz3Z05R02ho9ONmh9pFVjcWqYqZjWcN4RGK
SNostfFgonlP/pLjmi3x99Gu1mqGsr2jp5hJZArCZRF9SjMuwMjrwDhXxEuS
piubND5V4yBKT51oZcnPKTcZOvLe5hMNexI3IIvSxehNPtVWYsLn9sqWYWb0
4ZmY+X2/fdyJhSFySsU9eyRWcoDIb7DlwjN8LtznpTQ7J11Tmu++V5M7xzPh
EBirb5kzXjpHWpxmFAjIOcbiXiELMp5DJD5ZB6TELmvUpjQkfu5Zm4L2vTQB
gIDkCBDEVoXd4fEtyqs1um/VeXjfiDsNd319JjdDfVoyml1rZY+xt1l+7r2A
3b6oVVWYmKtOFqld8LAG6gM/KN/4hVavhI5MI82HcAwRQ2hI/JvEI+Z3cN3f
uOfK8/obmJl8jW8UeFuU1sS78f0OCBdQuT8+g0c0z7GkV+ceuquWZhvfV7Rh
mSeH5E4gWj4kt8GxjdbVLGb2hi13DiU2lpgm4eI3QL8TiLpCSw3H3dMyPjkO
QZ7xx4nla8EvZboOuajONqaOIo1iwvUVIaWGQ7V6exV/8vY2uT8/fMeZUj4j
0gbLyo3VsuohBPaMM81QiM6QooY/SY2dOtRTEg7R2yANOplFw+dHGpyX0+VY
MlJzvoPTxkViGE2Ez3BZ4t//tmtG4GCZmaF2ndlZSwcwLjoIWfUdlMvA+wL/
V7yOO2eiR3xJU8pfwcxFz8unA9Rk0E0UmMzdzMwpoI2qHEU/o5nBIZyoSxYC
pfXCKK6KaGtbKl0pwK+7P8FHitfyqfrF3SuUV/myuD7t49R8AxNrYrLr88ed
zzAvNvEOYfAVklQ8qLP2lLjKV//pA6mWSZMeceFJ6Q0zuczAJXsYM+lltYho
ql/hsrOz1B9QJhJv8z+io7eXJ8BarBzJJm56znA+0PwFzEaJjAJWWOC35gIJ
KGxlZrYksUNQ2SxTT4gC2xU8H30ljIuAEpSdBdB2IoSqny5wjVccrUqm4sl5
H1vcJDAadtZARa5Xdl3p7Zar9yXw43l4xwN3Mj+eTHIlMW27Gp+9ndWblazf
Msgl6gCn5zznMXREGAoy1tC78O7CDwVOnuK5ku3Jsat1dZ1diKzqnyST7ES/
TaGOX6cxigZbh4CfPY1p2oSoDRylAeiJ99kEfY1bo1Avh3Z3TJBJU++RPUrw
hRbKFmqE2YvX1Y2+PTpvWWcmodSmVjIK8A5TKdrpWuu4/c0Y//0HENSeTeYL
uKCY2PXcM2GPoNAtMwaw61m26D7dH2HElJNVp30Srk3F8IzvbU+JGToGpcGS
oE4ZW8DpJ3FVaHvw8KgfxbtZXA5pK38F6Toi0vIgwIDkGykf/ED0cNWmf1yO
dWiD8xE3As/oK4RmxFCgj99cyHl36dXgcnucYiP9NFRZnQOU/R9p9icklXIJ
ZR6Ubjc5d+wB7AbO+zZxsFont5Ytn1QTAGQPD1mM/5lqLjdKwGTcO3XiraeA
jN1N1U+NnfnIie+vCm7J6jkz/nIxUZ2He36HyzMe47j38v+C/K3PpkCjNS1g
JAI4hUSbWkhZ93JCQFjPq3V+EFjEsLlWnP6XHnLMMAka1eOXS+RiYHfYqjYP
FeoNo/NQ6IfIyCsD6b3CDznFtu4S7dQy5QFHv/malYexbeXWcjFZwx/FNTb3
3PVtGfK+CI8iSz0nlR6tQ7Qk2JTubgjETEu19S4hLNSzYz1HvOG5e/bDkB7A
zGLzIORxIP5LrtniQUAjytYH+JQYspcDF45klcPEfnOxaHPCsV16Am3Px7+3
UDWM+Bc012BOhrOTmYruSot+8XdI2ZQ+SVY0NFUr3I3bBPDY1lTts4rkfufv
rkEtsi+ud8ELkqlKtJbrvVQMam+polikLrTsIKrQlrGl033jKK7M5CMkwbUB
dB2NOHUPwQUIpw1uvv3KrHFapyHRldRS9vV6q8fxAGvxoGxtWvZA+czDo5Ez
uKNmBHNFocf3ds+t6KQ1wERc4U9HP0q9pWfp1KMqehn3RkTcbLqzuISise/j
GhTsfr0JiEmNA+v/Uz+Eiod9uARe7iet+aOlQHM68C0tZQAOCLl/SLaPkzy8
VMujjG2DNEKXWQHTT3HtLragWlK82Lt+eqXsCBuObF7Jgw6QB97MluHKUOWe
gv+kUPobI03TSwJ7Uv8m3WqY4gGNk1Fi18pLAsw8qZm2mPC33mN8eUf3M+dr
GX4X6gvvmKSL4kSbmaBbBefpbopGVU6Mc2q+tQ/nlMGWUosbCCnXJdkRoKV4
jhBo4DTT+YyhW8e0v5iVjgNqk83xmBlyakgcFAIloyr1nJtS7tDmG7JG7kIz
oLY4Vs8yczapZ2sG57lAsoTihyRLypOToqtkku2RoR/e9ym7qNgIt0XoqWqU
VaBbXb/Ihy9/mltJK7154Iq6P+h6OeQ2hNP/NrBIo5BQ1WillYQQ93lyMOgH
VkcIbabkedU1AIvuEMEagR8HDbFAjgaQ8GEHwPh0PROcYjlCLjd+zlnB/Tgi
RM7AW7jv9YLAqFIwpWo2QPZawOa1IUHekbTt/P5jyksy1sOMZ9Xqujb1sXMN
VMVPoz4CJDTYnxlBo54BGI6scl5AT7jIjfmKSacjRCHivGQ9ZY+8uv+HdWjs
rVP/t6nBeJnxsNUKiuiO+dJIvdqPOBBgNlcRtfNm3JlSte0HgH8VILsoBfFh
SOAuBu2EsmZZVjvzhB4mbH93YlktM9j+gIQrUeq5oYGdgsc7IA6GvCIODEDD
XePE6siLVXqse/GwSDPFX+UP5gR+2f7dvBtOvBSF2XWwNlTr51c/tAbSLO5l
kmcDDPtBN4sNnfqgi/di0Uob28rgqnRAM9Ow1NWg2LtrGUd0L/4McVd0BNqz
CAZNhfgSd2FRtGh5ht8oOJ4cFm3faJeStS3pobhZmwliBTwRYu7r5slz7yDr
Vuf4tH/rNM7fIZ+1gIXJqQ5P09J6RAacCK9y1HL9MaKttMTue6nOph+DsfnE
UcbYxscif376Z6d3BZwgZja+juTYonM4J3naprxu5ddVV6epLfCvxYUw1lRq
osR8Mu1upksrhvYo6Ki6koMYWEbk86OMPfAtAoj2cA+f8ud8TwqjabqQmIp3
u6jeHYgUKX+ZJuQchE7pCaXSks8Ip5TLIuBwjjLhKv4/tW2eJQFp63TqB7jv
cj+pYp0F7XcKsZ/KhAsdttRFmqfVcaI8NOWCzkUUK2Djyhjoi39a/ogMp3hd
u12F6MHzF0X01PWX4rqccEzfW+faE28cJrQ3VS5IsMIblK1ZSFaxdsmh9Rkq
YNsLeqWZ1YoaBM1EyyctXARBXW08Hir398Ev32VQBp8Om/bn/meVFglRRe+z
68z1o3pr/sxnOOq3565U2LPRacKCVwFiWggW/vK/pZ5hXCr+P/dQIrE6XvYp
77BMhPQLaMhexzKF349s3rAzNMAH3gsrj884ATt5uU/58pDh9hOZ/eW37key
7H1XgzqjZ+TxuA0yrvVDw5RIvP3c0Et/F5dvnaFIKoS5w56Y00YnrgoXjZLd
saJyaRIp09urF/byp4qXPWQEeillsAO5X712HvMy9E/EcutHFwfe3iW3EYE/
o8IlRdZ+Ck59rI/zaLhKf4sph20Wnd0y1jHNWNqOwjfNMiMpW0XpdndOoLjU
fUgymtrNCT/rSGnwo/0GZb0C1jDZeRw2Mt8hja+Xc1Q9yIvndn+ncs1YAGqj
6qX431xhzvg5QLzo9+ZLiQzARR3h9c3mtEF50+W7AQ+qyha/Qsm1NPbthtBO
cYSq4gPPxWcWoMfxYk4/ToHpNe7pSViSE9cLvCY74z6CW+gv6NCmS5Y3EP7A
isW4cY6mTVdHFEl6v2tUoBHdmxSqD2FT2VdPEfkOAkrn+weQdPE50AK3fnXR
zYefYVYEbEDry/LKHiifAakEoZwjl67UmNlvlsr1BJqykXsc8zW7dWeSUoih
x6COs3BC+VC7wgpXrOCkpZ5y8SGhmaNjSommy2HOiA1aJGOxs+JWZF3T6NKR
tAm27hVWKV3naLniskW09KIcfLtCTi0tL2ErhyYHodjM1TRuiM52aYYfBzz+
+/lJtWPdty3M8eQE1MZKBN1xAkr6rSeCsqfWXo5TkBzN7NgOfG66XKCtyYlD
CiY6Kh80Qsq+HhADIfCUmwTLRUB67x05CUaV02HkEPpHlmgDiSfAN/m9Tb2f
5uFKS/WPcEh70kbEDgeNpxRPvFCZiRwoh9RKOcQ24ggil8Y5G62KIc+xnGSy
CxVa2B9pYSm6p3TQiGbGKVRA0mlaC+xXcR3qcZNiMQwjh3dt10F/RoywhC6N
uKRv1jdS0ae23QAVnPpfpDRh7198RLpPW0L54uNW9wKrmTUcSxFonn/qNp1T
az1vBveq8DfSg3T1aDizeoOZlOsT82BANg60t0UoS8D1f+CYvxUbkuSS161B
kQAFDrLQhvEawnAoCWu3QRXmXlKO/xUB9oACN0x1t+llYxG7CSIFNjN1hSdx
DNoFDhI70cEejc4IAwhSl4hWTyfJ8Lr09mfiIhfHpfCA78qBWb7eaduzjca2
MgmCnqOnqyFL5PP0k4YO4v5e+gKmBbG6lRG1nm5jNZo8pBpwg04FU4URw3EB
X6Xpf/ojfG4cTdvNV6khPsUHCqb2ihwnqe5liTRDbJYE9pwUdD0eHrNRZRC/
RaUd2qkFPyCGDVdoROcBQRgca2LyGHH/6TC4hCZqzsBJfrxxa6lzCinfGr0J
/SR3LwqTnTE6O66CLOi3vT3ksgyG5JdcitRtec6CpMe6age1I9bhALQ1ZO6I
vD2H9tE6X7RkPboNptNHF5tbGAmFE0Hmc2LYyvz5UuDAJ60qLj9xWEqyHZx8
lnT1142kkmgemnLBdFGIWDZsIevpbjEOIySExNFkBnDvecPFz1R7dazYyhqM
wWGzmp6bU2H+B47TGWsoUfKUP7hv/QDALO6r6Vc3HYpxWqnNEOxa9kMavZzN
23Ibv7yOFohzcnxp8VXPUj4cu2S766Cz9zCdN42S3GnGXRQemYCdk5bmbss1
vnT/kFd3rT29BwBuHH4oF/VccboFf9kQA0uXqlkUmSmRb5BLy+Lkao9BimGv
PVYNYteyVnz0082n6QxD9tD1Mh6kshYBFMbbdslSYHBc/21A/TXBnT1qEHD2
V/qLoQ497a0tlPHJkMgT/igIdmYuDLriycfyqvWnDZsDfhC4mIoDfmj80jT2
nQfwnJO0e9MYV0/A5aqfDS9V6ZwcrQC5JJ0hF8PwnOj7x9cc6vdZNSOthhRD
Tx8hkcej9k/MP9yn+g61jqkKwVSFZwx9Zo7kbhG1i46lEx+GfvJhFMffZvZy
8y03m26BNv/dQ2iH20c1KTp2CPKBvJuJi4D2oE/qBRaRSyUPQFQiaHN1Y96n
St+iA2QZn/d+VryqLXn/ulrOQekKs5MengghqgkiQS0gA68Q53td6rZatR9h
vHxNQ2KroQOIQbEptFzUv/nqzUfSMGEV0k3bP/wR8cSbG3RzqK7r4Qryon5q
bPBxiqT9Vb5gp/6ZWn5YqVrh2/eL/2cXIv2KUYDm3gBPqmy+JFJazscNOcPk
gB8FNX05ZE0OSHNIGHc3k8hxzJUNCOeBWq7886AgxHfBp4H1ShmHP9gwNFyv
kwGEMy3Vt0JdwdJeNn9B86PUslo1cm41TC7ew0URCGWIBmrVob/giXZGPLBx
/I8TR7L7AKMsFiSlKLzdPGDnOe3BBYoaGfTlWiOeKg89QVYz/8dgaEe7qRtr
as3HLZ7la13WA3zMLccuNtDzmgwAAngwUXNnbkuQA/9OGq2JvaN1GizPSAFp
inkl/n6p1FWwDGsG0SxeN/H1vlOOVXlSnlfGjYt81898s38RCvWgxCtdf647
ZekMe18g6bP9Va4fmSt3+D38IGHGE4QS30Kl9gzKGVX+MthQVGpqvCZwGhm+
V/+tdx+lkB48CSU2Smn/xEWG1/AHIShpUAH/LfiLZMxmytVs2uq9iX7h9heq
eK8t3wQ+PiT2TNPrtQWS7M4dydtmbtVjQzyJYAommxayeU08ZnYfXjbTmwsP
umtuAnp4hP/XjIbi0uAixACy7BbcU5hi5iEDqbKWnreVEcytVQnrl9Ej0eJo
GxiUeZxIRS2aE4fHCxv+yZqwOid5nx7myzZdsQr5/KUAkxPa5cU7ZZrbzzEW
M71Gv+CIOw/a6/sk/b1sWK0pcdsFRpJq/xNUrFcMtnfuinvDUfoJypJXZT6J
IdcVFQR/aajb1nkfsifZPxpAEz05FetJ4rAjsRocXY6phs92eVhJgNYKAkdf
u+lf9Ell9MpWzCd/IcFcGS5AiKzjyBqZ3+xLrkevunQMj2/u+aWDoUlPuvdK
cXTHyTrZXCtdibICJCnEoHZOvTP/h8vndbPxrqrs4FuovFngQo8zrikbJmyo
Rk+EULiZ0APBmsi7IO7sZlExbKRuKMlw2rEDgrdLR9WlBYeNApI26J23prT1
7g7GtR5jn6jjqYY/ghHpYbcpA9Pr7CJznMYTrZFZGUTh2q0ipdD61Oqe2fM4
UaWRlB6nnA4xawTQAHQJih4OpGq0z5MQy6/9bluKA205qlLgBrEZG3R5dSaa
hlVW6VSk4xlrLJw73rIbxQvCRpOCS3QEfvsV9Zla9w7w/OLp/5v/w4VdJdJ5
TRs648dTxlLC5vMwzxLqdgGbwyHl5UeMYlKT49oKsi1qDksBBk8Sin1oTyAl
0azX/bjU98dBWXBlrfeOfPbR174teyHBmKoD7l7eaMk1ozupgxdDmgCTRNA4
Q/JDHkMyd6Fma+cZwkEtk4vHzqObBh2a0VwJ2DhGs8h2FjkuNCZ1XN/+Nz+I
o1X7C1+ZH4GUgxQwQImfeDoKeYCCyUun8WtcKTbIYQHMd85dEf0DfUKLdD78
Sa3gz9UsPqKT3IKd2bM1SQ7zwczRnl4ala7k+AJQEkcMdtvIElw1mXzHzXUo
hKpb1AzS2az9sdEKcj9DJZwZRLR3PglVe/LKXIH9B+QyagEBKYJQArQa9hhY
6IGBBHQ5oEnbP5d7s/jyVqPO8H+TvbnWuY0aPtObp7nVSniSgI+EyhLRJyfk
NLsx83C33sMCC27Fecvy/16SVdECaT5DdGDkGz3Eu2Dmh8QB4qaYZKXjX2Ti
IWLlOkcIm7ZH8zeTbFRifil7fLe9nJD/7ZjJiN9oZwW/S7eMyDiayc23Wm0O
yEdhu+amwtyzvpk5PwqnYbHgECB+i+9P6MqHx5r69fp208aqmj1gUfZ+BCH0
zYnOL3UubV6Yt2YQ5aTvTIm0+smOe/KzTUqzpfUP4KuSYGL5Bp9UZqXPQz25
E24avhIK6vcFF+LsADleDrlV0le3R9+rVmK0A4EWSbeYWrrWUYM2eYKCw4+m
s16HYLLHyffpgZMkYOAxCFEwt94C3G8SaoguwQEqXuimmLKqg6leaCqHQnUw
79cHwAMlIPNe66jqv/ZnNfgXXD5ZkeFfaGcyvoAvmGIFEtuiwEwGE+vUsOqP
KvMDfTzdQyMs6QbcGxSmMnr5nzlP4wKduRqSiIGurSBU7xw8JxLF3slUnzpO
yr7zzT1YPT1I1PWc4vIRvx2D+qyrKRz+B6x4QpDSLHTUHReEBkx0SHQ2Ao2F
L+Gc4z6bMVMyGfSVMzXXI+jfK6vvPNotIzqo5B0d0s25HMFPlThuylTCbC37
r2H52AgD/Khi4fstcExGk/e5JrE1S0gGUdnlTaBYKSu8rUtWJ3EaLIo+9gbt
ttiCOyt6gG0hOlFzzEP4QWS7yROaxUns62VD2viPG9h6KLcEPkMMqs6U0oYT
yw341929EcBiOByKy08v5Pfc2NevigwA3j8kwExcybGdYS6qYZtsLmh+Y0rU
pJGzpxAgnlmYtdcUcO/q82VtMHWtMIRsWYV9iActjwpIVymr0mxKHFrwBbsI
Zys9v9ZvCxj93+7IzU5r4k60lhYwhvLCADJwyDwLUQHzYdkPtcfJJRh1rE12
lTT0GpvupUnWBVJ1GxlxkrcbnPxk3eGBTKW/JVqcqLwJy1CbTyy47glNQ+YU
POUeliPWh84e5B8RRwlE4WUfKaraFpjZlAfDpd72l8MK2CnIpM5fvuhpH2Dw
7HoIzzzEoSlKwM5gGrWvt6+M9BAQFCvP5iLqnM+O686Ns5IYzNCugwV08AWe
S5pecuqoIkrxngqYJC2/F6dgPP2TbAlWOROc60Ufu4HiS3rLykq8T216+fyd
WHxGDoJ5IAgx9xEoh/FZuJl4wF61vXRVkRaNtjRDYVzVWTKL9MKVyrqZAc8G
0cV19IXWGqBf0BI0N9pnxDC1HBK6dEHzVhHBLubUUMYN4PbhpT9RHbMCCZwU
dMhTaTX6zMQ9hJ7eaPJPNij6hvjERxMkQqliW+hMI4lwk3tQd5o5r/pVj3qr
JVTyvilIdxgNBg+iPhBr0iH/9Tu8XecYOjnTjqIQidLkqplpCI462U02SJCz
VIOgb/eRz8ICXyg9jy/559sTzXaCwx3OBvpGzKWUmfTfDMckn2RbRPr37o25
Le+ldADp4UvSqlwWMC4UzvdSC/Ij10MR0SosdNg0yY7KVEc0F5AusPGa1Tau
ew1IUqqZHQczOmgFTf/K9V7RrsOdFJ4tLvkTBMdCSxq79cpPUfA4/7xBWlKP
x9o1eI+raBJBzL3zF7luHnROxBTiB3wm9a1jtgfhBDav/2xPI+5y1XfQ2zb/
cD4+aKJwrnEw8YrVkYrHzhREsnqS7fWie7vINYIG1wmL+gTxgbZCSNNK858J
STVBhuCT5yjejlATMQ+jFFpaykjiA3q18exjlshkxYGXmXLkn9zqqHUdRtkR
9scFNVLVDkScCiV/vkwsRgYb1W5cPZWpB25S3XpEKBaAA+X9dW1Exdo7sf42
EOlM3NBQrakXCb5CEuIhN/8JJqAJzlO3pfq9fujEQxt9TXBRoPZs+dfjmU8g
NkdWrk1+BjNzl+u9ug1Sz0NSMvp9lSls9nFmeLSjXSfGKr1wwKh2m/lZyWik
lZ8C2ox+Cx5N7gXkJuMWrcizn/rg2jlVbHr9s0jzcM/GcWwlUxaz/Abd5Ooo
UbGC50JaVZiU/ujLTz4pFgC4tsEz1cxi/tGd9CgVnY0YNO7YMpQ01nMJjipL
HpZimFtpaUlYwox+mW/6uxIX1MPyJ69IF4S5GJR64wQEYepqobH8PAxl0vs8
l7q+WBnEjltvWrBKMljae0kCN5ArlqJC/rECXyWUuP8Wwb5A+lMNf2XRHi6H
T0c7idT35HVKLFCcerhNbtnoOUhfdxUa2BWX2bVzL5g7pTkB6l5vqXoAHKWA
Tnrt8o7VhJ8kje7QiKpkOTiRpjGsDuLPkD0CnaaoCTjiTF6BNAS9eoerNwxF
uB4LHBFAoKE2OZxbegqKK6eHhO6Zi/eix55jV5ViSAFrqHLod4zcQ6PVWhHe
a08lqzB1cCIWb91+fvMJfsg3r4tlYRCX24AHs6g8F40qUHJozpZTx/BY3mVq
sYsWoHwaUD9m07YB7G49l1cV9pucb5PxLgnGxzsqEQ9fRz7DINb1zcfLt+Yx
OG8CHYYj9JanSul+AYaf9omgqh2UWcoWYdbPDvEHfyn9W35svBHdwttYQBKH
gdxqlxuFkCohJ/wyXPF3MSoYH2wWISvE9kR7ocozXlwFT4K03YzlW1LZyNX1
80mTgSkReu+Rw1CqcCtJIiEKqu6uNhuVCl77P2mLhGxYAyuUj5LhTgQYb6ND
HuyMVMK3yuRo9o3hQfDbUYwCnjU1w5EOYp9SsMkusBLRXr/sigA2zKwsJi0d
lL7FkiVyl8bfp2Ne2l/FW/sJiDO1v+IwZujxne3yHv/OJkQsBqiSlqWVH//f
QyL4+SMTHcWSdpf/31n5wgrEHw/tJM4jxXco4hsH6ZapJByadDG9sWKJI8GR
MMvc92RYWWJWA5DAO51onsSJd8eAbYc2OC98GVsWXA5D3ew50KOBfhXutTyV
7dlD8ieFYGf14i85Lg0Q7Qcu0dhgtcV27y+NrRI1z23vyWcBdexjDC2lE9EV
G/rT3QyqIZZRP4WnoFkZZaZ9BXob47Ne0iKW9U7KEK9pMFkJc+Zv7Zr9cKLw
D/7/o7+fJJduWepE3xJlbv6OQ8xoyhjtMYiRnF4gRfh6oyXnBDMf/norP11m
zbQ71905xcpGlSL6arDON71Bj11tSTmYQNu7UxCpT57a02hDBN+M86jpiFv3
CGUMSZ2FZbkuNFOW2H78pB0xoMCrVc3QrtEksLPDWiOVihfFfvv2O1uhdhy2
q3i6WAQU9FLzN/rCu5pe0DjQXUgAr1BGlnKf6OKz5h9MBOih4vwb3mLCCabE
NEmsAMXXsKBne28dHywqs+YcqrFeviymfG6CdCH1P6IL90aTfM1PXlXL6m0E
l5Sl9crdXNjQYJ+wcDBK+9UfDorbGTkXNb+BsHQzYzMyOhJaoe3MnZ69+CnI
kouUhOmYSUipYHPT3EVZywu87FwMfzxv4lV9/u2fCGYwrigiKn7Be0JUY2e3
l5hLfaxTzrN/k2bffTPqOE7U/L86N2Q9EtJCcKONjPJ98ifxLJ41V0RNlJWC
/EeuPNYC9J6vO7mvtWbdLmu6Qftkt9zCcA3aNiRepLWR9rbc9GQxqi2PdJVi
/7rTg8g8RiGC+HdIH+aPFywP9Zqr5D3ohzP5vPVyIv+uZERbLaDOf1C2k4fg
je1EWRebeCVPE8YDG+HIQH40BcYBgEBpc/GHKYFvmaNOi3kjkKgrpXykKdF9
xaLu2B/VZdFAGfKLwMafw+v3grPkUwhKWOeegBaf5KI/Gf/JNJEnDX4oAxdW
RdSurkk3bmn1kTLZysoBY/2/hEF+lckTvEmU8BbK4ZRum9087+M4nzEOGObd
0NBdSEQ8Pvhf/G1r95ngs5OVepENu4bijIv50OHzt8t3dPG+UfuNMp45tDY+
qUQMalfIe+zypMZ+XMw4O9ZqiHiH2XNzYMZAICqgBVnMDYB7cUKaCe8oGSH5
wo67YqsdQx+gUCvO3hrsHmJShY8t1hCMu/9W88GBt9uQcYGk4ruI9XsmzYra
C54cH0fkH+qUiS7wRz9Kcy3FdYFoucahB8z7WbE7S3BvkAWvOySam8Vkr0WF
CNDAOuJHqnDgUkPoV1HudXooXZFyq7wk0OsQpLg0qeyQJk/x/aLYBSYPr1Es
1PqdpjtST8DWIFaM5XCJ5rZETQ09+Tg1sKjvgHaTUwkbl2VjY2FNMHfltkvC
xEzDmabQskWryJyCxd2kdLxY7Qs7OI4xMicRug8H0ayaTJBzAGSi+PSBxX8Z
rdbOmYSdF+6LtfOhnMUpHIDF7cwWLmIbxLOeNiXMrrVyHN+B165zAIHfjBAa
kofJJKICNrw4o+WKgT/1WA8BN5/XfoeV9fOauX84FJD35oS2qSARS+cyxTgy
k72g8UCIZxoENfLaOXBtKGweqhODzw1nohD0dhPYHIQA5T1LU4MkzPyoCRiL
LTuO8s6PyeGfXQpQ7pijaCN9ipq/60UFnVeyVY0P0ZMieqniGa8YSqXLhmWj
9dhC5M27+JnxsMRK9vJQNfkfak7SIUEgP2W0pG/mJd7TlDbEoEMDL7mTTvvW
Am0KqFI0eWfr9DEAUkfVHqOmEyIQ8fYzVqCEYjqIN2ocz0Js/FNk2R60ew5D
6jSBS6w6ADch4GMLf0YP7dkkwmWGFLqR0qvQpIceTdoul1nkDZCNEOCaIUAJ
kF3DD2NcvvwSoMhuE2hB2IhLVXFCpSsMdphzFX9lZA9sakwNdD4vnBDP5AFX
wtYgUQkjX6dVOxOhrIq/mfQHE/hRn8xpE7ySRENR99lEOAAZTKLXkvJQ+ghj
Mw9O1sR85RbkO3rtqpWlmWmS9sbmHe0zY0V/O8Ef2nhkCyuvJBhuGAij0AOG
inJYYT2j/4jmkG5DYRjsklCWE0B98+ORkD5dK8cEH1xZ4KaCUQM3jYe79bzm
nH7wZ1wDp0+HcnYX5YECjmWIBOfp/TLanHKZsgYncRO/QBrbqtUu7YS0W33W
TvqTkzUFwkit5NtnXwoPCKEVx/FKE7QtUDZ7uA0B8LpRf2y3Q2QZu6nbgLHT
DUWvFW5FLssphnVf/Kku+libTM2tI0YAIwGb5Qd7a6zwt/zZdONxBPUndn6f
13Ofh4u3wTu2tOnAo0wFWM5Y/3kf7LZw6YWRqyZ0o2poG3+jqPluWCZF0I6G
RDKobWJly1NDvo83gY53gF//Egg6qap8AHBr/it20nD+qy38geOjJtARzImm
NBrbOCpVxNXlB1OPvY+2M3alIX9qn0bXQ1hW3NS7y3szq43W/YmuTgwNTn5N
0s+WE8AWqNlLFcAJ/1dl9aV1cdSM5MHWNJeS6CGyjdu5P4Na9NiG8CV+AWX5
kTscbU0C/Q3v+ALBmlTEvL83clfrsjrIZXmFMfaoBBKLp3HHTQNx0I5smbYH
vbYtP3a/ODYnqxzwjW/GCrmDuB6DHctOVpeLjNzCvm5y/w+GG8p5OaUcRTRp
iObMUOrKeGcm3PauGsnswkWbRaWieI56m47swZsT8W+GUK8sEo05ab9l6sOx
N2vAhJWRRdym5glIiVGL2E5rF2e1E8yx8otccJ/EpSGFEUBQ870wrncMzkrI
ERDeyNOPomEF3TQO8bIPMzMehx0doW1j3x1bZ5F4tSnyzixhiJ/0eeiC73bp
Q7UYcjbW++rTywC9QnqKCpR4lhRMb9MltuJ2VA8K8O/NuuCP0jxFHuPYU+NS
cJGtOY9eOMq902Y8g8EeAKZXt58VbfHvm6E+eOWrZ84qjE76Avht1mQNxJq8
9VQVGRbaAYN0RIx7cNJxIanMmQn4A2xR5uWKMNi8aDZM0T+mrsQY5Tu5dww3
LmzUMmxRVOzRAqVXhN8j1L3GEuAtZQ57ML182KwmDTvkBskCkpmt3HOw/E8r
UAZTJ4qeUc5y9GL1jwSLyBTnIGY9h+bIsMSeR6WlJ2VEl746dHoeYKiefFWq
LEktWeB57mI9yMK8+CrUIBUyVyFpQIF5nDS/onoedQ1kKOmWYmI1+fwoOnx0
aB1GqbpzSzj3TQIYD7rxNZ6ESn5fCx5XQLzGnD8rCpEnZqFdpla02h91JPOH
44yVRh3AbcRdjG/6IFfPOSmhGXE4+WNkQqAT9J2TPz1dylz8A2QPhwuavax/
1OugYpDUw/pu4HiiURlBpNpvi+vkJVD8nbGs71KgM7L6crY9/X4gIsNW8JI5
EYU/2TBiTkDB8zMCymK7+l2FnTk6D233XMzxQINS9eCd/mGvVUiCLhqnKiXv
SObasTnQLatqJldTD5PiLHX+HcXMPHHShgYe8Xwq2TpzZsicgglR4jSpjU/5
fHFCi0RIeGuabV8vVR/CUjCKJ0Al/U49XUzPZ/GD5JeQdA6xDoLOw646otwp
I83cLzHE9QJxn8/W7oijgMZfGFBJRFmlE59z0eBWYpKmn3jxRtQSLWCjGFtt
UqNdk7DtCVX4G4WDPEUPeDvIjDxBsnP8PEXpFwCZybW3/k1LCVx0A5bxc05s
VJeJI2XnH/68QnNZX48z3m/pDeMQVT7cmPJM9YNaCymbx+aDNpZSPsjRW8m+
ngNI+q0denPRyUcNeuHQ24rLT2nhPz13RmkL4T2UyFqXUJqKJS5eU5faesfI
JxExQbuakr79hnGDkPix1lg7iRpM9elCp8qr9SzkjuJ7kf399OjmUIWOrV3x
7AoZTbudAtx0EbMu9jc23vIvwGxmnA5baGnx4pfMMRPHC9x54LT/Oj6CpPkZ
/5w5A5dcOoEqPjN86vUWcADSN3Fbtr22MT8n6soWT3S+DcRBEUKXUNWvtz19
ba+73J97fjWSHiWFipT15Evb9+XuaQ2JqQpqjVZL3MwQVw7zeCgv1PJMKadL
l2R/s2+/HrNtitdsxBMybweYky+ouZEH7/aH3JAKWXqbkM/9GCmiyzA/nGoB
EgeZuVwASqrUc/h/FBxdnE8jEsuXZ4GuuymxPKqFsIbv+RRL0LhAJIM0adtq
pa8TGP3r9kUgy6KoCI/0CvYvDmTbY/pva16X9lLKlL8nD28pfQacyeO8/gfH
XD+3XnQcbAeLaOt3b6Qvz3gkEGczLYT035ZpJuRqn2VOVWWYJb/XpVerizgF
cT4COcD1fPW/yRMhF0yM8Cj79U5WHySYK9zzuK10tbkw3xi4VFGtNxPB3Xbc
zVCPpS8q6Vat4yVqUrfV9yYRi8EAMEbArVEki/fb+qOJmFuv1/85/anizrfN
LeQDF2LY0ZThrBPaDaCmG5/2jrK4+Ywsj1cwaaV2F3Ros89VMX0oobZko3Yv
1r4fI5hGNtBq7rris000y+kR9DhVCf3oCRweSzlKyURkiAlu8UtTQ8QsbrkS
mDuDhAckEinYmjle03wG+4/vKpqd/u7/OXDljfuoKmXFBLEgiwT2cUx6QK/X
NdZVta5obrXAxzE8d6OCAKzVgJObF0ffmV7B/p7v/IW8j/FSxTAfaDlV31I6
lVDY3fhTRNPAcYQStVifOVLxV8YRrQ3jkMRLyd59xVkLzkwPrRh/NPwvxy97
i34rfFrjHr8XSy+OG6f8Gfdso6BiwBLYJltEYm2Uj7sEpEWkX9GDR/gfTq63
WZJgxJ0wssaH9eCVGn2YLwhwgt48ZAs9EefGf2yhy8djMEQLa2uNCNgLMncN
5asGeE9GmDDJ6ZThGxOspItXyidkWpV7mcl8qu5laCYt1ble9et6/UixDoZE
euPorTbb612lNfdpvtF30dlgfc7hRaNdixFd6iwh0kKY2DJgpvvLXw12FCJM
OT9z1eSlgP1hE9lOT1skwCqVM9hxMUiJCfVpAR7lGLRNOLF+6z108UQOc8g8
dT7/72z52OVk/cQsalKRU6zs02LQd9pumI39pr5B+CwDNRVDkJW6R9YEmXoi
WxbFHapo8W5KTriiyJadE8cBZSvGh2CCfkTQWm1i1F3LZh9yDkvCNfTqS8jy
ORDXo0XUA7RkYeJJCQfk0do2owxGP6GtZ0vaPbLw6DloW8BzrW3f2UcPFUra
nfVDWCnexVd0gBiyqjKN/8N6VhtsIO4vLvXWulJfnprReU7Lt12xPIo51OSU
Y6CiXtQaBIqC3BW6gxBuIrvfOB775JQUtaAOYH8GCJv/N+LQqlyuZeQFQx2Z
9w7uF8HoR/d/6MO5v8pkP02KYnxW+Bawk/c69UdmUMBl7Za75tb338Rtz2BF
xJIBE/hKe49zG+i6lE+xBwFHfN/0sQFCfyrgm59hH5F+Iwz6k+J71tk81/f7
M9kHjD00yk4hHDLyak2AsdkA03LHIijWEOdPfBZdaWnV9Ebq3MEg1gdtJ+Wm
dYbfGBfWNu1P2BofwSWmzuKnsQeFpHZBzrMH8f87Z0LBth7SFvN83Dgn8tTB
t704Og6mIQi2tQvhK2W0Dw2YdQPdAraeur7vI+TVLEz4CXfdQReXhztZ2rhn
Fc3+ILcHN8R6/oSfep+1Tsggulb/bYzE3SOk/LR162TCFRNvVe6SeWpIuP4Q
9m6ZOOgP5gonS4a5VBHH8LN+b13+vlPisSq9QEWX8yL7qn/dfsvBTC16G95o
FT8kwbm8PaSf8i2x1HvxAZ53O5jGINwlHP5usaR2BTmusy/N9Tx77jwIhQ9u
Ju00N0ExZcRl8ac9nOtGTtYtRBTEC9smmgh6aWWNPlBmzhwQwZurQKVRnRHZ
Xc6yBEj6bacw6rWNSISj9VJRR4qQKt1aSRLUTUuifgi4jVCeorC7ANKL4Sq4
MDhk9j9DX58gbbj1VRVgOSnLdGc9CcWfC7D+RyJzQ8LW+cQPmdV09DV1vCYf
WzSt6s5PWrDLplBumrUAAY18mZb/6+/oK58YJZPuBcBxMsbR2GDmLuX7yvpM
EAKSYTs39Azh6TU89ZwdkQvfKejx11p8JEnfbIpGMtltfbcMu/e3XOHp3XCC
QgL2oWyn+76J8gCCVEKE9IPvmRB3Kq6fFZTS4sJjfMsvMW1CWZMZu2AdY5NM
76qGZ6KJcT9cplt9qkYxnhBwuZBO4Wlh2Mw4jXUPvd0v4MWst/RMZIVpEfVe
JjzIlnor+JmgNqG4meHU/cFFEUCmdWLUKJ4LGpyzB2afO1LubISNG6vn0WcV
4hrqEBGg7IPK/WtBWfHpjKxgiz9L14bE1omgPXTCbLeYoZI503/vDBqFkk9X
z+xtwb7ue3zphM/kFz2ldi/Cg+upQpyaUjn/rCqXPY+3apwNNQGGCPOwU0ys
MDgrINkPejIk/XJFr/bfEuk72CrCaSBJ/CL+i/QMdRyhTkadSUb+wRzZPCCJ
aCl76XAXGzw6qZCUcPbxrA4SJmBmjE0bEy6fkvPjTUpF8fypi/MWnmsFeVTm
CbzT2/OOwOgMYdhfpBaNQtF5jRRq9+xFZCpk1g3JhxRgMqw04by6V6y5lFr2
iQ02+FbQdnb3+IBLzcYQY5FHdVIvhbtbbeeC2MpzRb8UI3VVRBgIPe7wE0YO
mzLXm2i1E9fm5h/J5LtB7z+DXqyDV8t3jkghO1wFWSmr++yRdwQrgrZz7qQW
Hf7FCb1T4iLYcH1XLAomOrZy9lQ8MUNWH9qRoBn3lzFXMUOPS6tv3KxE9tzz
55+9XpvxUMuw+WTLXPBWHcUG27ksNi/tVQmvv+ClwAcSznIlNfOOI07JnT5x
fA+mBphNk/qXzG3XglQ5EPtq8QCaWTpi/t1Nx50qs57oysEt/mPSLqlOIx1O
ROMOQ5Za0gF/AZlnMxU2LZDsc45v5UHUvKRloEtumxNYLQoCeH7CC1sE0y68
O6NFA1gGQ2PESNomE8F/GZEenMi7bUBAGheD7+Exu9k/Yr4uTS45pHZL4vb5
A5gO2hrlhx6aWt1swYcSkwaG9e2OI4g7SBJODgMGFyDwf+L9ZmIXMZKnqN2n
/QGqw33HxJuKIxLUyMrVHDx8IlLeLPDPu6qe5NEnWABOPkoXVFE3++uiAAYD
klIkf217b5qqX9gxJWgCWX/OiUIeE9ENd6wxoud+yuQLsZ9ZvI19efTS7L8S
rggoUMUeHBrLMt1Ixb2zcCohxaOUvH5XKV6nngUBIUtYhX7Y83ApTrUbA84C
UQ5Ta9IwFm1RCpNV6GdqSSy05D8NBg0ej2aYVkp4StKPmuT5Ix76AlpXwQwE
2STNXRyC6tGwgQmp+P8R8uOgT1+iYRZk+6J30N6R6nXmzOuD+AHOIm34ad23
IYrLrbWtwxWRWDMFOivs5Adv/qjWJfjYIeo82epprdKTOzZ+ucitmftIKR4c
ZdYsYRn0Xkj3G2VsH6+hqhQtijBStkfGSx5vz/u7teggO20udhCJkvR1ZqKD
MfBzsOnrgCLF+Chu9zgVoFKCycgX4VwkQ2hyzIdjhC3IgAkM1zP6XoHWL2Pz
hwyNXA+CdGVguh3kf/oallqLJWzmusmQuHqwdjBDEhSQU9j9wotNWadmbyeX
2ZDN84yqxBmeIIeUIKPw/abpL6KMFXL6jp5cW0QI+LJy+HSZee1RyWRfG7kN
H7H4Q26JYjc2mOPwkG4Oi1U5vIG2/lL/naARdubAM5BeHW8kjY6yQCPDkd6K
6cN6sP1Gm20236eJ7upOBS0zpXBQ426qXJqy372RkuQggFvLykF4HDT+MEFf
UkI6vaxZnU8kSDQB9BhtgZ8uFbGADSTvzktyk02qH7MeufLGXVNoWCENqD69
xbqXLsl1ogHZIldW6jMKGt75buT8Cj/ZGmL/nclZc/fUBYIsN+I419KQJI9Y
/gX95jkpmpUgkaU7Jj+Vvgt/R/68J79cyLoAWN2LNP7QXp/GnV8by1T9zeA4
3Rnb2ZqnHNRri8Li5nbdhUT9FoIFFQINbFIVN3nFV2JUEjFwn2D3XgMrRPiw
tNfofNRaIdjSdk/8307Gq8R+6t+O2i1FpkdAFfGWjkYsAGkCCmXMVrgyvLpH
BJziU+2a5ETggEVjXpPYq32nJtOzBz+C4bsZE1NVOoAHtEGxHfm9rSAitxQe
WLOKBpnY67M4D/WRtodWC+5r5uFDp3ROlkOEAgvHIQNlVCJ9DW9NhponvTUH
P1hkYM3aGVg7GjteOr+ugXOVFeD1QZ0ijWh3fLca2q/ela9O0JzGjOf3117z
O94pBXz97KhdXkP6nKC1ww1DS3Z/vqo/64LTir3+9dbqleMGEfZafVJc8hyA
ZVkn6lz5LM5/75JQx3W2stq5xB9Z5eiA7Op/fPu0gdfDHNFxMXfWd1SYLM9a
0qUXdeCCfJtaTfZKchNXu/kjf1MAPEHwG5qIvJFEFCq0x5kTV8Cd1IxQx1ic
KTw1ojoFtcgJP7HdjTArqr4Q95W3fGxmcwZF4BcWmDRfcuQ081OttOzH7zTw
8/Gq5rRKmfm/Osue8pQ1oOtm5Vknzs15OgaQqOIm5FJm+O8+ePi9T7WGQ2R6
LHy8g12NlMJZj3l0NTs+2p0EAclEejTACSoGfdK0EeW0lsExl3fXmRrLiLba
l66QWikVHNtp4DFXY1FIGKKO36fJm7S58w3tXq1Mq5yhFvlInsYc3aBwKgID
y9q43WbIDTKhqfrNse5f79YEnGEC1+o1gUoiuB/2VHTbfJTW+ak+wd9+knsB
m/Eq+25OEZvODiSz88ELkiBbazwC7KzBd6Zyuhg8tKd90OvDa/umdjedV2SD
0qS3NIT1VVIRzcZCTYSY1IP27ZjAMG+PNqIevZaWIeiBvNMC4D9mdCUljrPK
ve32K+NwZR+rr5HKdxy112GZE2opPzUDGP/XNpNl06hLuHtl9jmfQNMioG9J
9p8Lqu2//l8zpg1ZsxjKquD7wwlXxQBr8APC7Nk5nIJH1HU1gmNomjCJTRG4
E250dOLHaUISJNAM+dn2nb7FQ7+Cqai4WYI+erpmBKuBPHPQbx3E7gXwmq00
utBVyPsQGGF1eA3VFK2+L1zXibbT7NUcYPPb15Sk289x3pYbcdvyJkZzxj25
MiGCvLsnL8zIXXyKbCagkpoFCB88nhDzhGPqHN/FrAi1g8ITXozEK9if9KT5
EYyMbiNlmuxf6zbOHvJtRYmkn2HIn/4latV/kh3+LQR5oWKEoAso2WmsJoGo
36zxLKMEHObMe/Uz5wtJTpC0rwn6HQm6+tbb8XKcaiJI0mNed4fG0ZVC4aAb
HXQdip0N7dmUzah5eb/vAC50/X2FQ6GUZd2RiyFlbAxTVbKauNUGczhPNfui
BjHSI57e2PkW/joVefZkkzhVOerZGqsdrSc0wfxeZ1YFFkrPTUcueqWovxjY
nti71HWZDs2mqk+dIMR16ad1up/9E4PHC+fPB9MBUcdPrI+9P4h6Yk+QRZ/M
BWCZ4qAse96ub8Kq/1IJw17IZyXrgUZ6FljoJcVwC6c4acpO9aIuRBJJiWRQ
EKQ1iqSeM1n1ncNPBV5iuqHrzCT/1uu82k8xX+5bRcYE4L7KTpYRUzEnFnqH
AdVsT7RShiPw8PUFn8yAJ7/XGN9/vFfh9Hl7hB4dVrJqMM/1JAm6RbjLroYf
GEXGECzlzCLIaOrZZmPb4xzo5AIOaClvxmBxZ49fl6KmYK+wFKsf6x0cY+C0
JkNQXRodjXsbsykevvQFvD7cDOtJkXxYIzinhxCgeeaFiXJZb2zOqGR/gC8N
vezhVk7l75ByW03gXMo+1Z4m1akp1Uf4MV8hWpIgk673dmYEXaK8YRk4l6CR
V9W21N+rRy4iBa+P6dS5PuaAK06jppqZ+v1D+v7bsEB3sDNuLuCk9YncHpw2
S8WoF0sCzAPVnrok5lqDHkCJlxHczQRnJH0hPNX7uXFQ8MorItmIJX908jOO
earH58LaqZ3wb1EbSh7ZgMc/TkQhASp3IK/0GElqDVH4J1Zv04kjtybUxA8G
e3ddoqmMh8Zc+op/AJPrTRce2rrFUh+FrfmvaoUaEkDTbmpCFDcRtT6Zn0Cf
0h+2Zyd9DibL4zGk4R6b+6fSMjyBMGcBpXewerHF3VQTR/vAfe/WRecH3xNv
MXw13v/+fxh7MjHkqH9Zkh4utpP3RnQLi7Q4BrmEz5yHOypWaZG+olaiYju3
jqfhGyo62oHko05pTTLIJY6YkH9iwolx2KQqDdGQ8Z//9Y/k+2cT0IiBrOo0
e8rypDT+r3Zqqli3byM44+77ejxZaoSFGpeXOQuJQWxBuYoCKY0XjI1BeGJ6
QyFzV0LyreQLRihhX7b+VU7YsZ3/qerNWjgngUdQlBABL/0+sVz3VNghrw7y
WU8orZuBRlca9De6iERBzwITsfb8zYF87IGzyWLy256KhD4b1cA2HHpo1SaN
1N09yv2socGCvs71bUaQA6ZKNavRc3JZPA6X7G5/sFzVixDzdNbdeXJcgbn0
ZD1x/U/lWm463ukBUVtar+9TUOlNVf0QGRKTZN/Nl986aMbXluUkvEy3DtYe
JNswlm2oUjdag2CyTPDSEr/mQOv3MxG2hmnroajFUFJdmVi8cVgV/EsF1pfP
9s7py/8xLT1g1PyKcap0GAOhV5rJaLFJbR5392N2tKsLr97P2zAkxdiQImGy
qISsleYf4qIW7vGQRqudzEVQd9jkDPuTw+2C0zzF06u0P/sO7oB09zSCIkAT
Ap2OqcJ2F2A/TDNVVZaNMjllUG7EhyAI3lmpvvhuDv37j8AsNs4BekrUvimc
74oNvJ+f2GFmwFgaO2K3yzrvoFb/y8cWos0UMwUdA5xEuRoycYV1NUfkyvJ4
JjQv5rSpZ3ZvKB1pkd5HQgQNkEqqEeKt7NYrGSeQilaaw8ydyS02NcBNcUlM
vZfcOCUom/3M/R4f9XWdK6CFBgoAYRav6lyxvNn32QB80WrNUreZ+HaMivVl
MFCpUp1kDEeCY62fMDA61YruuJ4ZfRuN1F9+4UAd3xTEXpKCZtcP0fMiMV77
LJAGhpyYLVDjB34wMgf+Cy4+JNxzkYuhJl3alZMyw5mih5+rXchC8u5Lxd3Z
gJwYXBWrszIr3ArfzEMiVew16UGYxIw804a5On0Uph0ppS5Ygo4SXhRSAAP1
lJJQRS0yY6J5KFKArVGt9VKTRfNUTX7ALE8KNh3CkcZU1a99gkUIxHK+2zmQ
CmOM+3Y3R2081Rn+oasJW+nO1DGBg99DEftZe4uvOCqhX9gEw0E5W/aHvagK
Mei/mgSVHV46XExlmcN+XFUrBVCra0O4VxSar2/cP528z+2VSHirjYKmOady
k362gNAtBFg8/J+WPgj7NM9H8D6HGKjWarPcR6tsK4WLBwEsxmW/txKP8wqG
H7vb9SKRWHoijrbBJO/d2j153eiOYVXilyix6+LZq7AiNsk04UNRMlF62raI
3dMj/lj6je4EgDgV5g83ysoFn5JykK0ri+oskA3yAhCN+vOFoBQhM32NOryq
LuvcR8fN9PjoQGG13q1W4n+rFtTJIzJVyafUBLlHinrQzokaICM9yhAPSgrQ
CnT6b9L2dcs+2KoIATLvqFd+z93QgLf+FZkMKY1P5BynE+BfwwDmW8uGiW6o
Yi+31GT0YglVpZlRiG4WX0wvg+csuwFlPK2oqh49k9TOVb6y/B+tmtBID/1Y
ryj2eGoDsnpJP26N4LcCbQOwPCvMREzShfL/jarrHIplYRYy0JAhvN/ACRXE
n7cOrTEJiH31n9RF1fVAU+Yz/kjbIPySkobxZH8KX52wJwIYEgEd7qUg0/Ac
6pNPrcK313Fyl9DivaozPU1JVbw34cNWChSOIUTgczEijEmiTjvSQ7Sy3gTq
GHX+yguW4xNi94MULWTiCKrks4R8eph91Uk+JYZ9QfNim+boYNdAUauLMjJ6
XiyGxPdM4fih7XesIKLQ1QpkLnDSIHAf8eimw2LxgGqAwtpl/76q8bczqifs
N7e2l3t2Sp4u19lllCVSB/nt4D8TCO1mm77d7KjwtbF/tiJ5dOrDBLe7F1sR
Mu25H+j+oWkVQpcsLMjV1X4/aNQOfxeGQTgZvWi0+jN/hMg1pdechyqqWi1J
D35UGljIsrxN+DF7vtM+9bHGlOD5gOQJRWNnrS3Xghf7WdwQgf53cXa2bEpQ
9bCfelvzATpgA7L/J1r8Q9UWwtzayd1gALv1FoedIjJ52HQxcG7s5MElPdXi
X2fGeJep9KGRpi86EuRlPZz/ScxoQNBOxmvr1Kh6P2MtOKlj6Y4QqtecE/vZ
NDHra4L7HxKl/cZnxuhPK5vYcEKs3QNoU5aIXNMoirEdjPKkGU8NieKwc0O5
ou8ap/ZHiAoM9M2ZmOcDeNGOFBArUWfCn8Vnu2fqOgAj0XzFaXiSMabDDjmE
5AtY1I/T2N5Kwl3V77IDKitxd7NUy7jXd/OuMKa+6B1JUPneS17xok1J2akj
PZTIk8i/obAKxvAMWomDR0NRjBfeaF5DEO+uqNsLqDNYf4nBDMdlEaGBIdyP
PWTR6lrg5jkbV5cr/5u2pL3a9etnlJ+bxlzrSKBS1a7wWAOhBQMwWy/NFi5j
13LPj9T4x1UR8ekyXVv9eYZ88FVn1mE/xk9ANSgDrf8JB0cxN/Y1SjUbLdMk
wA4q12U9sDmtsPEWr4wi44DBaY+Wsf8loAUcmfhBLqFt2/YFsh21EeVUP41X
e1yMDGbilG5v7m2A5NhgOMY1CgYnmv83DuS+068l+7HFNPv4Gk62zoF/XA3r
asUTAsFNThFuK3Hr8n1N+NnzYTZG6I0J+FVQPNGBp8DTTVoMPBEnvFoqkC4t
Bt00TcAZZ9RL4VYAslGLxO1zqQt498WIz22/KUT7UvWyjL2erO4X6SklL2mF
YZ2KM9ZcP3nOip5+eF9U9JoiMBNLaBUbUiSHClr4PylJWjlF8XvPsE+r76Lt
ypmk2Y9QLYL3zva8Cs11aE57AO7XaCruv5eWKozDm2mogxOxmfU31IWGpJDd
wXaTEzLe7wsWiWjGh0zu0/0sJAMvMZPJgSEEyNtDUd+lMbw9apsLB5TdBVfd
Lki6nRR9eBMd3sBep2+8YnSuJMNzcBIqIYsSWnOmzevMgJ6yfuNpQPkA8fxD
znjfQTkQaigdl1LhKa/JRWxi+k+KVagAps7JWjeom6qMVU6KYIZReG8G+w2a
Q4mgwrEh4+PtFtINVZolylHiIMuWNH1+x2JAoUA5IOnDt/1YPVEctX8nqP4W
6MffvC0rJ4IA+DHccBq/cPmRCiwn7Q7AJpmAuPDIZt+N/h1S+yTl+N594PRz
V2Py2v1WieLO2HZ9pTcfi+GHU9WGQe1+4Ck6V6edRk3Qe8891kIm8gajg91b
e2TOcv9aC4VkCNAcnyBASFYAeXw1oDdrjdY9c0n+9IhleZBxIyagmoxNJkji
wab7XoFY9FWQ6A3nOVLKDNlK5LtYvgkza3iGbZYR5pVnxobXd1Iu8FDgrH/W
7Cl/faUDstPWlL/phIlV2r6vy8gnBn6WeNnEKDgFkJDBOQ21q/o1r5f7Vzi4
LSnNN2PLAN990uNoxsnqIyMFbvPRF7zkYOjMhJ2BBKmcFSmXMXANBO2a+iFL
N/r6EMD34TI2Of5OOfTOly9ChGLibqYiBC1hRDDPxdodkpHtPfsJKa9fqGEQ
Y2TMU0IXvnzerbIe+cVK9O1ls2CVRR4obO9KwYt2XfR9PxZP/joi8s6HDJnw
XeDkKqVzJ64kjRl4AJNlicdpnwunx1LaVT/pQrrfWfmkvW1rqGLr3R7Od21u
ZNVFmbx7Ex5HP8GB8B4HArL5G3caplpxf8e4lZuAIyxtLldZUjyUzwqQR9h+
jMIJqvnF18VDdRJi7ibA2DJeMlK81NVtLizeA/duoFTzAUAkohjaoLmk3bVZ
9SoyqoJtQgVONCyhsXJME4Mk25V3WqghJsdBdTTU5aWt3wDmz/lBMQhStnUs
AFPNpZb/lm5EVm5+ou7E9aMynIaip1IQhx57hfWkSsrIR0yUS1wqdAWkYGVT
LEjr6Lgz2bEzzzb5ZUbcMdvE1L6lENoV4DYZE4zqIwWHJDWYi6vT2s5AExmM
ExH1YvE+uhxnC/GvCzrMxoqO/uKvx3/a20vhR4cJf/3uxt5Ut8S3Ph+2f5Gb
NPZNDz9RAQMMssmZyneuTjXVQlRlzamuWIDkm6yav5EGEeNJxDwIV4COB5sL
ueAv4S/vM0aB0kOswWhgCHglep1qncjmGaiDVv+sH92pBCftL6nC1523oCjn
yRoTjrFCc4N93iQ7ZWha+kSNccXA7HEPNPWWl6BMKrj+Di0MxIuT8MbaTTs7
fht+MsEEr8HEnuCSGXflZHdPci/sw0pdrQyAv7WS6xgHBkcmoIsQ4m8MkEV1
AJLyoWMaEfTzy2tSPlb5vhDvkMnbcvnGUFtmskIMLvkOrORGX511Gj4DC99U
PUmrYLc1RMUDKpgBeNr6X3MphhfHJF+79QC43UOiOSc4JJZKNcNU2IEGXo8V
J90Vd89JgViTV2TxSfHcZWDDktAZSzmMO8VP65Mr6DSRY2izP1DEnePDr+qM
H5yCoq1tZ8HYItysJmdKoegglhcIu/ybPWcntp6BfNwHi6ay4nWqLjeL4Y/K
DBVhON+viUDKoCMPKP9r+u/cq72VmD6x/wIW8kFvv3lN1WDhVzDOgn6dFb1Z
AxpFntssZ+GbyhlIoUuzUs7oCelzLghvCcmqefX5cL+MZUNYZ226nVJ21u3Z
14bLWc1sd/VtY/SfTKz5/E7CEYYVe4jopnEntoFvKN4s4w2kDVUL0Tyw5+KM
/WrjNcz84js00mb4boMZ+vu7Q1qhLbeTElYExqejMhXaRj3RdXEzGd/HI5TO
AttCosXjemNy4zLV+dxqMn0kyZQe07ppBwZmIqZEMvvJnyDontDYLyXcTKFB
7ysAiQBZ4yK2fE4cw1Q4yadkWV6mkabvJWJpg/H6yGBc23PwO//odFskfP+g
pTFabNX6bDHr1GLaUVqOIrCHeJ2ZbF2W57MuFic7R8PoPWYDfJUwMxyzjZ8Y
GVl82rYOcOPMlFb2ju4UmfEERIq1yj5eNmWgnJLH4qbKtYRHQU6fLb6JDX2K
BtbI/bQDVIEBJuvC+t/aFPUiTG1KEGvRSBOrm2aq0BAGHXNWAfbkgly2WaGB
fbASVPZ2uroc6XXzi0cNmG8gdRMp72BpB6dGzl/sVncfH5Fs7Rc9m3oxFiWu
9HCu1mZS9CNf2BuJ02yRN1DIOqbTn9Qxg5Fsi257LwTK/oAjPokatYAgy5DS
AnMIIb+F7uFSTNJQ/WbPQWomQIWj95cPFTZV0jq9btSOuTiH2Rt/8zCBQeO9
2VQTIz/o6nhgAZyBC7q7xao6HNiBPTcu5wTtXXVt9YuyQ+pkOyYMxJv7y/d/
H/W3XZPtRhhMTNMQziYZScjbQG1OvkzTSKpcxKkLv3pudYWnPUcXG8/gaBKB
x+nI4e+cssSN6bLi+1wCgpR/Yg2P6+rdXSKsJWPpkzdrLvO9YuDGbe++sOy4
qePuUsanmGZII3gVCeOAATu6xruh1TyxhPlzUSBkwoZOOuAcHXlEs0y0sz8f
4AE03vWn75C9fXlWTj51WK4EfxdBVBR0gJ3owRk9wzPUmUoRBlIceLo8CVMn
Z+iZrsOQdJv103xR/M0pqXmgibECgh2zNOIXROR1SaTvPBta9Vz+B9I+2fT1
E6jIBomxwvICMKLwpWmxEWzoH2eXIeNcHIc9EwAyyTAHo/wAO+6tWGRU365j
SarvqYysHu0ZzwNu5pLcUdd2O10N8voGWfnNmitMfAe2QmakGFDc7nkqsoVH
xggwtDncRfkfPi3kkiGqNriohBih4j/qTePtwm33mnTl8sJL6rwrEOwsT8Gr
CkdjC5X9WjvkHdmnNnapnIjX8II6f+ei26jNNr2tdm8iYNHm6RK/E3p8FndB
sTVGR8jELyrBhznq/hSFEmOE02c3JLRCKkZ0S8XkNxxM+zM1eubuGym9gX25
F4/06S//5nIhCfMRIFtPxeG/PV/7VjFqnFURfDjE8AKP0nia0iH6gZ3lV30x
z9q+Hjr9PgfW4hfTjBueI6HPVtNJyIqZJGJVjlXc1BAPmPWDG2xuFIyYf1Df
yWlB1rTGLGWbjR6Q2YUwlIg24fh3fle5ujrZoi02/08n0ec1q7thV97jP25V
RvUIMgu5wDphV47c8V0s9N/Vbw6nF0Z8vQV1mVBM7SEYBVZhLsVAbNAiDRHf
h0/wPTrcBLJ6M6Ebr8xJ57QMKOVNsAeXDa1SXClXOdddke3FWK8sLrfPm+av
Gbmd90zec+J1W16x/qQhQw6G16NhkbfZ480lmbOPTqsf13rFNYbsiht4jQrG
oNxg588AH8Nrr3PZYlX/HLgZJqwqqGlryIiawjE8vOzQw9LmyQ5Rs9w9U6vt
ehpwqgnrhZ/pjgV4yhen04YihDKLDHfuD0k68bgYPXvfvakndiy976wy57P4
P9tYP++ceLkeYNBxV6Ps4/nLRVIF9ksbuEheeFQJ72OSmrG58w3L0NV2wkUt
oHShimaZxTAmolf1gBlEa2NR5h/eOxYRYnN7GsyE/1wpaHUy+mvh5vShoAmd
BA+fW6+aOtrDmLvG9A8PdF7fdUJSkslX0ukHd6NLBFrp3SOG3h2+Ff3YBtcs
yA4T8rw5YrxkdxqE7ZLakjZIwJx/JdLsRQIcBBoN7Epsm/iQmpPBaFVTEZWR
jFJv8vF7RNbfP+UiPszwppm/Sz6Xd8/N239h/CxQ5Fdiad/TfMDkbmgRFleY
S73O2EINGi+rDgQ0J0wZd0wPsl1ASv1TiB8wWMo8Cz8Nqo8OLddYw7W3BA2O
pg2EJF5OEWLL4bYXGe0gNc2lSZDXSgi/Ywlg1yzJYJOQUFYvxsVAPtU5dG+0
3FO6GbCyeVGmWGYw1VWtzIYD3DegYT0eirPKHtnJlMvhGm2buyFUURgkww7t
rXLpdIem/zc+1QkFwCpy3Kpu2w+g65skLmJvyuBbZCuyBbgkZjiKHi8/lQxl
Uk+WSDsAgq4Pu1BlmANtQPmJlH9Q+cn5TX0IN0GzXloytqomUvkNd0gSpw66
a77GTWTloELEkbSKG4au/tO7N46jcrgi/ZCmMFerVGmjWzaHagg+KPse1BoK
go+xbbB9cRm+LGXnVndm4VarwCdZEUsjZes4rDdllNdxrRAAjRwk/4/jIYIX
NtyeMID3Kkf+X8dpquIj3HUZZo/9GkdFf0swmkjBrmvWIRUBQ54Ld94XL1Jx
KX0gH2Ab+Je2P2+jUul6w/BRgpCsAmQGuPt+3q1o5eA22EOjecscCmMXBE8j
hrC9LlmQDVxmGKH1dE55dQ+HxwVaDlH9kWLWGNjMzgMePtCso8enHLPkpvwv
7UbTohTJhGxuDeOWMvwEL/5pRmYh+mnSHRfXInrr89deF57ZubjqnMEJl5xG
ZTqBWvZM7zEPT+h04uMUQWBB4FS1RLFEPXhRJ/oWxMwJX//GKj+CX0oyD8SB
e9jmpgFHRpHZorLfWtfx+5T7JQeA6kh20Ouz02XaqfYO+ddPLeQuL7/MoJod
iykVPkTf9M54Jt1RdQ5DoEnBKw6t2hbjQkkc6t5Ecgou9Qt1WDYDF7lE/lW0
3zat6Z10dZ1lHa4uXk0SldjTd/VgwsubF4Y4NIp6enpRnwfn1wzAgT2NhNjx
cmCK5dMqC0jG0jZarYP0X+x4c1C2IAlX4xzvOssBhenSy9VcaU2CT6nMZS1k
V+jTLSWJ5TkNLArEhkPYKOZgjiY639aM5GVYdkB5udKebVJIebCERPdWqLAX
zomQjJujViNhBm/LJB5LekxmgGyCYJ7mSRTyQNUwPx65wKfUZzrFsZQDDu0L
SC4/Bd36yXjUDKNcctljhV6C/guMrWwMmVlc+KtRMrnpHkp24wq1hc/KQwFZ
a6N8E77viBS2wV2nUG128hkjhBwrJEELKK0Oh3alUbrLuReOe/F7Aa5Q43EL
LIIIyco5cs60Ll37DfhSlpazVKgTsWDFETB9V5FCp4fdVrCqR+8Tn3BzkjUt
HCfskeYvTtvPzgQ59ea1h6le0cvzKopPStfxwtegx8h+yGhgtN7wvOIeiBkd
TxfMsfyOI8NtEpYn3paEyQbbBmptkoXQjfcZnj5k/Jlx1WVbPYc+/xXVuOep
lZCCVnsZS98feE7VjPS9GFsHS7Z0IfF0SSLm6fUdLXqa23CD4FUYzvxFxxSZ
0rTVnfRU9oWdF4N7stoHpAvzMeBEtALsQosdy/FhAmygYUkia2Wgk5EBWyQR
au/utbMAhwmDl/JCscTPeJjRXWBOmROy2MjIU356AvKoCkcES8LnzBczqiER
JbnszpX262mpDWcNIhrlgmcMhiPs9BoGTGYFygOEmEB9//Y3/850LrBCyVfj
mksFcmP8xu0cZPQfpbxqYItApJCEG8dd/LOBd9T+i94xOzKD6BrHT/kW5ZJX
x/147mIrGwwDoQ4U7QLoskKOslEsVGGZB38p61rN1IskmlgcAd63rFvuP1/x
PIwFWg1L2qH9tK7uViTW79yOeIayc4QtZ9xocfGFr/Zt47mF/xre7IBQHUYj
L88LBvwDD6IOnqHnQr5Y+0jYzV0UbOb8XNM4Z54SIZapKHFZYBYNks9ZJwtw
XO2HIkmEjGyUYkLNE4wR6+vjqQJZOZRtGoFkpEc9tp+jqA/MfrUuS6NKM5se
6XAS4tkKQ6i610Fne7sv8mNjfV3DhaqtXxoDaCm3o/IswuEknESNwtCBJUDl
9pUcExK3Vy/OxK1u9OaUORM7k4VuEcaxcHKDTsLa851ZrEkLscCxkHew5w1p
uxEAaO9Mqn230lnGVIGAWl2uH5Yvsbe4Nms2JFYwLeht3qVh0rePYIqU6V3B
LEgAWXJuSSNlm4fr96CpAxboZVSJvYPAGfnJBDTx19BD1uyrAJYsLPfwRJQU
5QvpqaH8Y4lFQSxqUu/SneFySp92meHZSz3E9haeqLQuImzndtTdYfO1Nx5J
t29rgczZrxHfvojHGh6PO9OSoafWssj05RZ52fhZv3H736IsnHlC+s1p6ehb
GSPf7HOX6Ez2euTciAgkNxXJYUY5Bdm8LJ0iR3llrM9KP9uRFpAOLf1JsNBq
nR7nhWsbNB/96IYgmNICzp+zLym3X5D3uRLhN152JSRYAzzvbSXjybSyF+tS
gISKeBfAEshFJuaPwU/1bd42KlVImmb36xLYNvK3M2AzhBKEomk1UsPrHHZf
tR2aOdg9Wa4i+80tYSaM2IkfQBgr/51ZlhY9KZj3lUv85s0GdirkFr/kMtLm
YS25ejn1O7dUsORXqznU9R6kpKqDZesDi+2IBLK7M2fB8+4OFtjRJwxjM+3K
MV8IG7MX2/SnFztAoFnfDHrp2r+Hfl2W4cXhlWJZ2B1iYIkpRa8etkmqE9wW
ycH2cPbALq/71Z5qb6dG5ee7pu7r49vKCgRYQJUmsJhsEncyDCNypkXvnVHG
IWM/VHJF1xP8wNNRCWdSklqFdP5IhTSu3MLX+9ReLmuXNazO5ExIEFhhAAp3
w7Xl/1pd2/7XVMqZle9MFeKhycxrg1urr81UGlAwnUI9pZkqkmTZHzaeNIFn
X95J2lcrwTOWEudJzazTHF+ovD99kufF5Nxlz0qh8pyv8c5SQazXmVeBXQSQ
TLAdchfY3iblEkfkVjsPXigvVjTLzd7C29AUkKzTUSbsJksnvX0tlypj4oxK
ygSHJokVuE+t9opzoHykQP39l/uKEzT2HPFcXgspr9Mgz7Ex8/RHOV+bCf41
mpbEahkvkbxdWZX4b2xXCzuCf3jr6zDv2VddBgeCYGkbZuQtKs12Fysl7sTh
opS2yuSmvFA+EM6W8PHlFUPz+0Uay5K7kDYQ2suhY2UR8vblnzd89WsRagH6
sVbxZUVwyTyeQRhhENaC9tzfjSUEVeEiJ1CRctZ/3nMYALO/ZiNgmIyFfjq7
W8FD2hxXfnktavhNZTaNDqrpVJX/VCSFtCcrQup1kxNJOctrIunQaWB+1BJh
6IHLOk1DTXVHSO1H9i+48x3gNp8rRo3Z/8jqRAsD3F8+4VyM+X8WQtvCs4Nc
0Xm0eq8v91GKLkn581wO+jqaHZ8ehq95h6Wn9Z37K166K9CBaEiOB55wE8Bq
D9M0914eryasaznavLKyWC+hXVy2TgviB8/m815aBK66txFsfKZJwuoHEAUS
no2yNkeGb89ZFzyUcxKAy1GpWt1Wb5KhdiWnko8K9GK3AW0hFmF4STtcjn0+
GiMW8SoNjJUW2ievO1IugfzAfqGlg9boALEPpOfLlmWOsrizYwE4R2902Vo7
Z9W39rCRh+PPjLW87KwZmAV8HZY6zc+aTF0gjaZbX9Ih8k8wXcQFTIZ//Tj+
GjmCeSpmVecYB/9E6wFbymSECIS3G1pSe6brh52hy/uusWM/c2ZdsVuJR/KG
HNE7JVfyRgyBamPWMSQM08HcnolRNEVZmOtdPsvtc2gNF6atn6aofgqWKPU7
wC7nfaI5bRP34B34MtYl1FueW49JlFtUWr5A82ywEPT0f58xkNq+6SFU3n4Z
Sx+OA5FzvC8eZZ+0wtCDTUI13FQrYblqLVv+Et/UUBM8WV00tBkreLdTMVwV
5QPpLBMxgpWVo6rFQa3Ev2FXDr7hZ5L7NNwO0jxUjc6ijXL6vPN8juV9MCxp
G7vOZZjELUIq1z5mXb+2RynwMnw0tdJxpP9X1LSI6CfTa6cw6WILzU6VXBnn
f4KF3ztHqJy6TGENPRBoX2ls8UyDmwatwoL1sXsLK6fdDL/ojS7JeH9ADmLj
qnjB3hPPULpuRW2/iCEF2/qyuXcbV/kyEX0tcdKSOGcxEmect65Izo+mTRBa
qE82vJr3iHk9xn0HZV/e38Vg/Ke5d2FS2wa7BHvznUJ2q3kHh4Km+2JO9PYS
H2Gkb2yhElOcom16HaF5nnzL5KS41MLtkTuZJOroxyIVBwi5462yHDQowyXF
GYvEoQgxU6FVNGEGuZQaUFsuoXyZzz6UgFBTmEEWd+apPzlpj+R0VDNPYUZs
a8JwwxWkpCWCG3I91HnKlvtXxBr6ZbJyMBRA5IHlNyNyvYDIqJi6McR9X0hf
HJ6FfxCA//pODR7j49XWslowWOIYRTsshrdcTJnWMus7c6DclzyJZEWwoUhi
RKTIx0/z+nwmJhMZmCECDrSTlBcB7KdQqx5Qy19jGjvrHKH4ZMAkFxiDgmCF
KGamavkmvKlsRTjXYBu0qWdV0OFlIIykGC34dA+oF6/qP8fFDh9ed750aitS
dlzFT806Igcc5wzFDfuuCQBTLh7GvmixX5JaphWyP7OdYKIfgUIDUOHqI5Ke
MPCNpsLb9/nz0FBi3kek+uHoKQC5h7NFsJLfQM89RHT/8JoKBS9AyrJnlKiP
REhbzEl+q2wJLZsg+GfepWP2xbJiBPKhEV7/OMO7QXpYGiRlBlezdyynXRuv
CNNNwhjpxeTxIAXtYSSLMDNF9ZO6Xd33FEk6PMrlJIzGKMlUiO0EhiwynZMe
7bULNOiFOb2EEIyO/SQr0OA9fSms8KTOckr7XAmS7YoBIfBawyyHRFN8xNac
G7U9e1AkCBWwV3AHt5tAR74EKFbOXPw3Sby6jGcjZ7lwd6nmQor+iHAlW7Tj
K01SS12M6zUmXgA9QwqfiMw+35WErsCZItyZy2YKcCl6jQyitTmaTDFeBEs6
UntOLDwMUDrjY/7RPbS0LtZfSOOea+HKxOua1WW/IJO23zMOtDAWFzZLoSVf
MhIqHWzoEC6qvlmULF4npWzhSo8tG07ZwWmNcTpcg35w7oBJCgSlIDt2Ckgv
tALGXCrfJC3LeBpnf+/JlqrBkokIW4UTMrPTkXJNpa1FnD2Rq0YI/wqsgt67
hyZpT6Qkgr/qgo9R7lHMWGufy1zRo2nUWiuiFnxze4hFbxPTZtVscxGZlPLZ
Ezi4kizYWGVdRTufO+ETS3dQs5YnB889dYOPqlWvarxVctFohsU/YbOjRfce
GdNtvj8DLimTvkkC+ICKf8DVxrIaPvX2FDOEIcS+8SpHslK9pXK4FXB9xZ5W
UqMKp0rUnXd+4mYgwBWabGjrg4Pc8dwNX+Fu4cgbcZGeE1UcpBQJIxQ7lEK/
iiHeP9A4tFNkPlwmselQuZjJ7lVc1GcUP5DQNVSXnta9v65H+RcneVsmeko8
dLk8Vh3+7MF5gim19tr4NDGip4TnkSrP+EkRTey9obCSt8gu2YfQLEGRHi39
g1Vfj8gkeoO8q2a76uC19dR49iYad0N4NpZEalPaOWI/ox5dJeGslmfE1axA
ZS5zwh6xd+i3Br4DJ3hi/2a0zMOSppChQ7hQIGg4WhNg3Yk0TbKIkJthzfiG
DqV8NylyjPF8o/UXStJq9JL7ZMiCl0R+JvNoukOn37WkHhSzx7i5VuQ9WJ46
6XEEqHxy2jkFxzzKDia1QJVFUtLvro1DM87op3XVtT3ka9eBkiU6mubwrQCc
Zsvnehfc3xJ/Du96zMznzGszGRceVlvt+OYZOe0XkUbTRNnajq/eH37Igjjx
sMmqbzGZQYOFWExS8LFcQOlvXrLGsVSvmxjzPCGIXPLlsoLb0OE+38T1/B/g
POjoOao1RUyPOgxHU+uftbEd/Ra/CHGNagc3DJMoBx7w8S9WjS4aP2KinrD+
nFuNV1qR2cvK0juUWm2xZG3xenaheAKEeaMXo3hAdz5m4tBkUIXB7AYdlNbj
U0tDEDjSVai+8deeetAEjdhKZNNXezN+QY5r/S5J1I2s7Kqvi/TzNAkpkcTD
A7TlXe+ZLhENT1JIX4W4gYjmFQo0L5+gF9P2kmXamehwLxxVTq1zX63JQ4ku
CZMI7KxgDzHQ0T8mRYjqxU3z7ynF7SI8dMr125/GNqoqO2rHa2CF72C+AGhG
sdTdbuRewDj031xwz8DrCszmELlQEg8tszy1nAjU3IlRxpiZIZlvIOKoVM6o
OpxDx8+YLASXU+L32FSy9l+xIIn3TRu2mmSyxpr5Sb1oIx4E1ovQ3NQq3KJK
bz7a4UOjt7fQ8uystqhBIEUfamschneyqN4fWCiFmF+yVhIgtbDA11218pis
qG7jew4Pwl+NYRrUuwrFSA5pu6R2hfHs13+aMSO17gqcfmef+vt41JPg0pg0
jNLqDT93YVPbAKTJDLFY/9gvu5tLqe1u1gkn2yCqr3iiReXTYYGXTPrW6Ss3
e9zkK95G+W8fwoLPccCr6EZJjQ08wMtpiZOdeMqBb24xZhhXfGy1bC2VSCiU
0GYhOucR7yUBgoAO5RujPE3cHpkmwiidbO6H0R1zILr7wFuwdQ+HSRfM9ycD
qdlrUhiYj0gjZwOwR7qkl0eqw5bfbSmNwfDqIJ50C4zqXJnxOXe/zsbptEeg
9qIRVNLYmEY1t1ZoGkW/PinN7X/+al4NYtuugAL3YJWD4EQWyTo6etG2s7wq
8pxsArSet1K4KJqur1Fr6gZw5t+cBphvbq7xx6nWsJdvmLpp7dfkKKyAIIRr
IHPf9t1b6CSedA9nhydGg1nAErtG6vESlVE9AWxGa5pG0Qhx7Kd74r4EmFct
g+zIcLgtrwr9HVfzRnJID64/3q0YYLAxwV7ftNZKehCd8dqWfiw3XPGYuzep
IKfILmFz+6tHg54wHr/prkESEF+rQMh6Ge+XmKh0sJ00zzTb+Oamoum/nyNn
3sBWbX3qyBIoxvvIpgcVCgzXXJm8IhQdWsigHJIJqTUobiWV9k/dzSecRCTe
ygqbuCbtx7cDskSjUwEUloPIncUzYe0S/tmM47cSKab7Ac4jPLl/b53CbzD9
QlhoEfTJPwTl12qjmA8CpEIlJRQbUVediwHPDPNjZkxxjQrzAlHYliZ5iQAE
42/csJjs/IEX2xM3zxoaUh4msSUOoTQFYtE3WSjeNBsFKG2A+i+HcKIbBKJo
XosKwG9nQjULLW3HKpfL+csg8woYsg9JZ1UCfDj2+sPYAdKOY8JoOz0Hr00w
iSni1t1CSsWBKw6Zznxgd7XywWdc1HaQ0Ms79AxLUDdbR7c0pBoFcB/PmgJP
VH81qkJtroqDWzX3ObVpmX54Wz8DOOAsFeEdcKTT0EoJeBvj3pi43sAkqlvt
vN1u0tGN+NJrd4UkRWihlVnXn2E8TCa2zFIsAVHpj2lh3O52mAe5toyilaG0
trBd3kc+EhLQ6pgVjqiExH+deN708/2x5Bje8t9rjCOgA7AHgfU65RHwUlAk
kJlx9gPoLKZ9Wa0PIlYhSxvLedD3Gb4Lmhx59KqyuJ1FAK51GGJEMAkm7OCz
q9f9+XEcx2XyZmz1/srmrHDHkfPYC7qvPOm9q1QSOVuD4iRpBd6c5fm9yTMP
GpVPmd2Nx9PR30gIcUqHu5v7xaBtKzCndP6BNF9w7a9DPxB9eF/1c3sqDeXD
DJZ3/KFesYDymPrJPhYz6f7pXr+4nlO0BmG3iiHhoQRB5k6y2qaZ9QQzDK9p
5sg0uMSYackdDU1eOhBnyjMcv0D1O4Uf5LKiBWoUc/NAKM/er38X0NV7blQ7
cD/22PjxMoeOJOwSK2AUdNyqj++m7A+C8yjtfgwlmvzK682BYgvWejLdaQJi
Lwg7g0f6t0oBQv8IM9iMDeCKSxswwYuX27tDWw0QCuIx5rl8SK2xgs9Y80Ti
1bG8+/q/iRGTo+CHdgQwaK9gzd1kInzIrMsdGO9DMr/c+LOo9ri5T32jthMc
CNB3cRcxxwbhtpn/W9s0X+wheAHtda+/TL9+gYZ6ibQFsmPqW656bjibKOCI
+9c5pLF6MqGTpy0wadnysHf/fn2/uNb+fCbg8hcUmUVfAydIqkO9ok1MwbWD
mKRIcOnXzfyRw0ooY3KQuR7i2D85d3yzGtqOprgAweK5jOaF4NWeR8WBSako
97QmtjeIm2Ph+5QoUSkEVYvTRzbCzXBkAZP26Z0hG0D/wZPrToxmSbmCzSgo
JttTJ/2h7Y1QQKUWStWarPraGdp7v4FZWJz8AKnrsKjMtVUVFlHOlkA1Ga6q
EO9k1oVZ2EviQzAiiBWVHAoG/hhzH3SSGidlfEDcGz+966h2JYf/FpDg9+rT
DIT2+UdibEk4lW5vQoSFoUkm5UXRk4Nfe68u0kicLQ2WpiVnR9v5s33ZKL8z
Zph7dKvJJU0pKR6AICHgVD5dHWezQ8IsyBftO8QlSmO885iT2g8GrHiRzGqN
zT0om0l/CTxkVnYyQC3rR5flxXgYYXJubpj8b2Q3FtGWadNDxYp6qDK2Z8rq
/Jzqhg7mOMjMgW5Dol2CMOd8/QuGL39UeFNYSsSjUBADxLhjezuF62bNHtpj
5xLqP1WKBFaBWNXOReYy0QJcVdjrmAzk+W6owEvNFjU66LqUf3O58oZHhC/h
JRrJWq4uALrusA7lnQ9VoxS96AnoVDXU6kSKoAL0dPQDQkjScLToO2/MJclR
VnDMAavoHcJ7HdypqSqsv2ZPfb4iTRu9xvvM0jJrYchubDLOCReDnjqLH3Ko
jIYv4iV/gQN+nDPuR2nlTQOr41NiJbOhcOKa5CwoRNvpU+hpnezsCLrmgioe
UfNbevVJwFTDNC+8G8FpE7hh4ZCHP0hLYGaNY5f2BhE7aAmu8UY+ctWniEkQ
AvO6Rk6wjSvRKpR+ws9G1RK0my0TL6GmdOXhRJPBapIBvgW417Z1Fe0Wsd4G
Qr8IkZGZsH4PQkVzd4ZbplKLhbeXy2xdXYnEtq7uuM5xpIYN0+UtFS75+Hmx
7AJ1dbGFdGhnEZh/6G73fhe0yQ+DdMarIg/s3DR0eLDNNi1dh8koaXirKCQ4
KXHLr62MaBD+9a9kFIPz5JvmRquekmO5jb8lis7xRMj0HGCV6gi9i0k7gMs9
QoK/iof96D3PHq6ZyF5Kn7SwuPNXkuJkLfGl59S+jRJYZzPD24nwW1Ok0clT
9Oxyta7eCLdj+EOMrKJgx3Qj9eXHNDoCvUCjqCQ/jIdLSAYLbrNdVIRl206M
ZnbqudFFECS0T1SLxpeawdz9g61k4mTXRSv/uJz5RswdSOKO3947kICyzwjV
/7jYYITpiPvlCSw17z2sJFGoTgXV/heLMT09Il2N+veQ0kjl0DsiyZx5b1ns
JLh61sqmqz9BWyyPCNTFmDyYxvrqlBWgwIGN2FmyU+0zmFDc/ROryrgyJ5Pm
ySgyC/viTqKUnxo+esTiGrvu6E/qAXVGGoYWPkS+AF1s1N0nGEGpsvRAztl0
GXrWUC+LTV0JGT25NxiOjNpWOnyfozhTyVGZgSxz1R9hedD1/TpbmzDDwr35
TDpegb0YikkjK05uG06PBhEqO6ecRm/PElLnIO4l6avAbh6DNcWIzwg+b7zz
ljeJsy5FhLe1aWt2gm8ie4uVm2GR7BBMFWW7nPvKACNcflVcJnTmH31a3WSf
+G+DriI1b7NZT6Rtfd+RoqMG6hrBbbOlUq9/g97md6gwYteO/+mJIr8YDKK4
q/xZ2oieqJL7ZfNF9oCZg0L9ybKHdJEkBfuV+f+8UBLRemYYVJMpINFBXgJw
NL0g62IlgSZXqFjwVRfpGLOQpjdano0wkseymzQ9WuvC0lJkWnwDUPAg1WEi
d++cUUcNsXadj01JkSqdmY4fCZ859HD2y3KO0OwtJqam6t4RkT7CcKHKBB6R
APy8y8vKGuYlpuBAwCq6Kcki9UrstGyCz5TyV3xCOivo2rAI1eG8PSUngS3k
gtt8heeEiW743zeBhqMV1FKK9/Bfb/U28jnS5RXq370WU5lsVu1QLVqPyXho
ZvdPrDBAzBcmAlg1jNxoHqgztAN4mHK6Guk9TILF5BS4pO32nANMFhxrFxx7
AhY/FWO1JBnvztzh4xuBTqv5YtTcZoKlOujTjJHVcGK6X59jaq/bbio0/IUQ
yhocVQaZEtJyEUyeMdSgOmB3lJUf/JZbihVT90LAL9CaMScqcoO3WixokNKU
+cetn9SNJQOZl5Qr7s9xTeJnbRXsmZeWaM5UXuz7nf20P7FP+omHrN2IUgor
uI4KuiTcJaAlAqlVdpDWWiHi/rvSrWFuyN8j/M6oc5sXVxATGR8PsMTRpWzR
LUWaG8h2DCI16pXvkuO2bYGFZi1Au3i8KUCYcWdmJ/7fKMB9ugQwmHEIIqIG
nSS1kKywXRB9tEBSxXHc7fHvXFxBsU7tr7sO5QNoZeDAhAWL9CRD2rAF3y9b
aP2rrUQAx+rji5LWjBYoK7rWNKfVY304wA2hUbaUrq8VNdv7CGJpJ+jSYSfq
7Z0FDa5R326SzAf2hcZU2xzFLgS7hzs7M1A1b5SmTMRDdDEg1wXI7vUmEnUp
jKc+XvSYQsgL/ADZl7RBeXpGu2EVSyt1eWYr09nb7K3VZEgvuzQ1Aq2n90wv
Gl8povaWLBnq8UdpHbDXnZBwFCTpxHkqf1Intq4OVtJ8ginZvhwLiXBBWS3G
s4kfA80kP+grMrKPOd0ZD85ygoD5VewSG0tXntzihcSKLtgGQenIeQLK2Spt
p9/OPq9leqHPyYgeQOESCrSmr/ESZ5RqCg/z7LDPoVC77D+KKfxmwyh60PJN
jTgJTZ/uoumfaOIA8PjWAj5ztfrcU6VmUBC8F1I/qvhn4ZDe8qvgo1XJvQYV
RbDxvCYHFjI4zoF1tB93F5A7SI4DS/B/sPTOMRtkTaMv/RbUgIphQFQeCqjb
z0BYs7dgHZ93xgXjhlEp5o30RaL0PxAOzhTNjKw4OcoqcCZ+JUO8ZxPS/+Ac
4XS++kzjqiAEoF+tEW5f+8ZLoKgShaqGsAcBcFIQrvuTDD9MbAL/79m6GvEi
JbGPDjSsM2MdafdWuuPQ7IjvP9M/UR58tq+oloBleVYr4QNvikQnBDAwg13O
w8Rnafd9zs0bfJMkux4w3hshKGod/EHCYtgAN32ts+Slxes/bRBJU9MQfLIh
wGaemTR0qGFGt47vPVCFe0j89RfB9+VulJc5qkXiWMvdPJ+h+g8j7jPvUHVo
I51H0Pwn1fRxsh4qy8k8wRbCqVWK3SF5A87IVI9x+mZFafp9lxWYmXO4RiWU
Dun2kRh604Ij9INWPvp50ycSMOU4O6Eh0Cep9X1b1zTC5mSeVAhJWAhJWZV/
bA1xudVp0lYaGyMvCltdN8peOh2mEMDSOjIpbLTx9lS0sNQpnHg2pQAEOyHw
p1VNhMuAYgTs0lM9A7mvwIEJH52gzzJijJKtBvQchfh5dkdiBWnxW6iO0huS
BVqe+NMqlI9ekalt+prqQS3F5+cs8uDvajsRa8GzBuxJNMvFPGqDCpTtNXAC
X9KcbJOZkRSd4AyABaqME4wllr1igrIWZ1LwaNAQW+H6K/O8WqDdvJi4pD+W
JMpe0kgE/TVnFj0ZW569PGTd8HMJNJO2w0mZr34XMzxp0weYGomCLlAAM09I
3MhVxQ5BDd9UzxyovPZAr9woNGUOHOQNRFWXSM3fNUkD0tUGCm+yZoq7AXt6
j5Ik6S1jcEI9VQDFsYE2UURV78z6vXxIx397d+B0aFoxNciJG2WtsTwQpiuV
Wh2ETsLJRVQNPhfs94XUX+CDaTHYZDKmjsT20kIxR8/dxprfVRO6nzTfa8rE
jE3GkBibIWNoSQcH7Ygz+cFSG71uXSlHUCs7i8H21yea/UjXZAtx5q8uDzcM
S6whyEFGDl1myn3fUDNan7dCUgkD56wMj7K34/aA5s+txcpgGRMGTm19BF3R
8/xABcjgQ2FpRPyOUcry5IiHDjpplm/B2080N8X40Tt639km8Y67gBpVpU8U
V2fCBNAhNq5VXUS3cVp40E9VIyiZHbZl7OzJ9UEgGzGi8mHWkFZHfZarL1WB
DSALDJnDDqkyCjIX6qZ7oh/FJFyUWaPdag5zQ4878xDlPAX6GKVpFZdppdcm
Z4qTUHju/+9JYKe2mQkVo+FpGUonHD4bFq2hEc0fZ9PWHhEbyzHHQdrf5n8S
GSoRj74SYUNk3b7DZpJFkJyjCOAwWitZdx6L1NU5YvgayRgXtf9DdTsLtAZW
Ff8CBv4kJXAQARvmoMxTH8wJj101bsW8i6D/pPgJhi8n0bpckq4EGmucvS7p
5YLwZvtcX45C7V/mdSEhJmBxSNi2NkecWy9ajGZ8zcZzZxS+UynMOZgfNsn8
G7cOTYR4L1aiQbkW0ZtIYxlgXlgoqe13MahJ3L2Bd5MKdJIZlzl4EdZvB2mT
DXgqGidpZoaeFvrjMdW3q7qljyEo5kqiKHbVbssBTxYzQZwFHiPGlzdrXZC+
N58C5hL4rb13+s+cMoUpLfjELv/7BbCJ6cxlzXZddEfz9eaFxc+xxhhU06q/
Z5F+85BIxJWFUi1MCWf1oUuAKu3zw8Y6R6I1IMs4CXU0cYtNRVpRQQO0yz4l
V1mvKz0sCOVfCUtHni05gGwpp1nZl9y7VTpJ0bIgLXDo0Ekz6Nvymz11p5wc
tXUDcMYJrjyCJ+/CKvmyrhf7Jti7CXZA7dzX400ihglyxpl2LM8++exVXMeR
nYHiFV5vTrW6xRfB2iQcHvgUpBlT9SFOcJ5DZYS/WQkjX7++RK/2Um1e/hPS
f5lVetFaJdJsvKJeIryW/O3wxSrtr9kAMB+k68j09k+MUaG9l8PjChv7/y/+
HJwkS8FfHXsaMsH1333KY1U0wmjQgU43ZeogV7Zsv5P7C71cTIHJCs6JpdCY
CDmJc69YzZbZKpStohXf2ag8wb94nSC/qE/MXwBp298O0ZBMPsTBOoLstbzC
rKQkBdhuklk20j6lOKuWcGAH8yyXr45VU/S5CgV/jUeV6/8tXmXVcDMGygtZ
fs3UVcOxHJc70sYg5hMv2njNuu+krnhikegSXvBvI3ik++20/PEDF9Imy29o
5C4Mt9iDKBtmKu2RQfQ/xhOwNV5dp2eGPT7ibNNUSVDDFkefJ5/FXjU7UEx3
ztO0OajKvlDHeIwi9qP3EqPdCyk/awzThPYEyPVYuGqQ6d/HWJBKH0+gGUtZ
pbIQxcxSIm26GU3CkO5PKqK6viJeD9vXtA/Ve/78O+vS10oGZW+170rB2nuA
oSeSwA9COIvkDYYC8Jz4gtFPehHmPtF/pa4FiodxhK0Ob+bM6Xew27KyPkyy
ftlfRlPGUaLALN1dPOU3AVfhVsWeeJVI96Nad5Jy7auP1zvIbFCSSnm8NOj5
OFPT7Hkx6m3HA3ewF9nUVYY/ivHzs2OuNnHrW7Sh2ZWwL1gQHvn595hY6YIk
Or5ejJY4zNKNJ+Etu5wv5neflIqPiMkQU/OQ7MqfXrkFWR+5yFOLCyR57Haf
P6PZlEKmFBAq5BBADF8GBGKTWxrff2SC5pFDRUGByWL7QuiIlSDDRDQ5RY9t
J4JRzc+C+NIVwGY0q10OSIfATOyU4DpZyIeJqiHv8lq6zlEZiHd48/U46FXn
ipxvGSmhnvUTc6dcW7JbIGuyXtRiM91em2W6HyewZfhimERHjUVNwQNFuKU3
GiJgovBjbfu1KhvsjMbZtcey4uRd+6Kooj/fqF4a9fQjgYWYmwdVOUkSAchX
dvuIiwNI8ZtI3zCQb+PPcXrCDVyQ0yRdftHDWuIAi4KZ1IedhRZUpG4Q9oQX
Bb02M85PSZrOdjXXRywiQE9Gg2SUE9uq+Iw3klaGLD7ni/9QmaAiT1wxsaBJ
g6AsVjYtKCEKhESc3aVdd+8bRH/M1WwewjAVOnAvcmqjW9zJziSK693oJRBb
SNnx2irpo9BH4VTY29maB6x4GiuIFuIs22SU5xXspoRA53GHKiFAv0C2dQyr
sCekBOT1NxscHg23p1pzcIkakzu0siGDHrIM7ZzKvr/yrqyrCJlPzEB/Lp+6
fUdJC57zqfC3Gwru7LF3ZMj5L4HuddFn2oK+2cOU6PW7TMaFm3GyyBibuUGc
KJCQyC8dNRXB8uWADlHzKD7cWT7bAi9d+fUteO2XAPWg8O6AFPUzTXavf919
cI7wG3ThPDUHzVoHrXWjJoltwe35kKN2FO59gU/PZTg7j+6tp72Resr2QTUC
l+nzxUGSbq83lsyi5B2mNDDtzsDUd5t/Wsex5EkYMpZxYgtwlInqpeLhJSpk
KjSZzEk7hn8DxO7YQEOi8GTGjM0LWx5hBNUgACSIvn0fSfj21sZ6uexousoY
cTMiHW7c6VVMItCfGoENvAEJrA8xj94cS66LhpyaGLw2obaAZEvRshp4pEox
MOxi8AKeJ2hQ7YAF1OExfAcB7ebFBtmF5zTFuetroJN8oLFQt3AeSK5Mwfzi
UxYpwkvbyi6hSjQaLE+Gfz6JfdctcESO89dSeuuKLVG5u5NDUFe3oUwZagkQ
R0h2URhiYcUHi3zSGjlUD/D8njLXZVjtfbBjNOH3SwDE+h0ZQGOZg+zUVLd2
PPCVKA0bAq4h4pskh+F+m9AQQpXJZAQAYJRS8T+SDm3d3TPe8yKoL9fBOC/h
X+v6ToWeKWfkmXoRLhNmlcez/2ExeR1tmFE9f28aMsQ97fZCRUKsUZ0j1JBj
Obv2VQcPzIUdHHyVASAdvvKhw1yjVxLMSgQQ3Xsw/X6Q9GGRZP7Uv6DdGmDV
kzYuDT9KUIhg6OzkMyZiMJWKbPVxP0to/Tg9nbUvZlWSFW2DHCukiK/jQ+/o
gqWiL/1lTCKu+zNX7R3yVEoQa0CyzQ48c0x3IEj9QIoY8/p+uDdixQN+Qkm3
2VDHfHPQoY5vprQX5uQN05DKnFqFcF/WWzDEGauRLfnqNtSj7YhZgzLU+5C7
iS+xYurDD8vnLAkqzSLk7ItC/DP1CdIvQ3ZHfgIzo70xwohWGU23yAXGWWS3
ym/ptBNXwSHZ3VKhNAReh4axLQ+iE7ggKMBVn2QmhatR/L3VtY3G++mLgF2F
p8iEi6nfWTYs1l4W3zlPwIbE6pOUhkI7DjRNynVlcut8mW17XLWthywfjSi4
xW98+AvM8INiGYQSzyPRoDsdgb9PnITNZYvR7lyfMDPBP84+RLW7qcgD+1Pz
wGYUUqG8mwQee+uPThJ3Sp5tfvx9p7e782wvKMk31feJI2TLk4dZUKNMSTJ1
cdRGX+npQCiZItHb/7zswx/+zjtjKSYe8eT78pMzPqIbfOLoQSyKPydt1fCN
wBZofxXrOpP440V6JyNbQv3ulgWHcbi+l4KOfhSwVL1lHQfYt191WJuN8673
1k2tFF+HWRjM2unWdYRGDLmIn8qS96GW/+K6nU/NCCRhpGn0yiGfE+jFSFcI
t7/KU9DyBDWvLpWkVd8viTQ+BjKohuKEBG9eUtEoRi50MlmzK1urayliuguF
NPmbVT8KQd3CaCkr6DctkVmRjL524mBqE0vgI+c4Km6DSGrbQ5EgeNzTNozH
nJwZVvxO/xD680R9XF5AInTMOl/I1A1UxsJnrKbkzVNB12yx0SCKyI8l0nQ9
BW60TS+rCaZeb08VxxRuqjoaWcCgi5MfiNeRjClGLtl+2h4FcZoOw9Wt0xtJ
PgyrhlsDAdjvpmLOxQe2VRyjH0j/4tEdCjalsJO08nCW0Jm4A4h7iTy4ZrMN
L5dp8JBkUveFea540MrqrJyNv9P+1O3XkDslQFeQmo0ARDWB8F9JW07jANCi
/tSm6R0kX4ErEvx2NuNMdBz84HipQdTCdeRajJeYsRBmiSBZeI+QIWPBOhfq
ueIL9/61p6uz4bOsXh3y4yL+EbStKt+pWxD0vNOi7TIt83oIjVrewefsVZzC
RmdAaBozt8nHQVBYFLCW+Of5gHhsFf70hUGMEy48d52I86qn6nKUH+CpY4oT
ssFkJtw6pHcg016UY4PMOZn0yzxY4dYLNkzmbL6etb/d1Eqzm/EgaUfRxoQv
8vyhKUDgHk/RhvQvvkxfa2Nfk5tkiHDy1yf88jF+NEZrExl5hgbUD4JRCiZV
OmFEGdi3VHZeO5PoMQBj19sJZOZtH1K8Zg9qtEX8fbDHDlU7YAJ+2NUlhF8j
1+c4UP1T/Vq2GLGn7Z2wu9tIFMJvi3rBkBhcIrgkkeEW0rkubilZj+cfUCOt
zYKHpg/AmpUT7QjFREp05sxSpqK0J3/DeYhRDLNd1GdX7beV2v0drQDEvkq/
OU1Zsyzh/cDx3NTLmumcDymrE4wy1s4DAgKUioTbIPgEn+I0VsfDiRszlkrr
y/B8IypRuJ/ao45z089mo/fc6dWh5DmF/pcsknLVO6RYZ6Dg+c8KF8Mppw7R
cJ0bZdq9eHUg8QT5JEHfU6ULxJdTyqfKukOga1R1qysBCfh4SIcBXy66+ncv
HOGw3MfmBvWA+N0wVAEbby1OhzMm3HX8u/88wKxU2F3SSDhOXoIC/M9rktiK
0btDkNeA8K3qSJW1+AHbfhZuX0UsP31FxlqcjMmOdiEElWYEmL/ACdgxk+eZ
L3R6clWxGh0y+Zc8UZPix6RKoaGi+pnriekPOdulQ+S0945n02N8LzchVFYC
1xb7V0XzGCos3jgIMA5Au0bd8CaaEjjNfA4eQM/E3Vi4FsDqH4re4JTJ+9Vr
aUIWP6afAOOgjuRqJVPwCcT+BjL1CXtZzR2rg3TcGUqMfbyecEmwVFZ70y1f
yhV0ytXTa9bl+j8ORrnLL0vGn+qEFBi7VYdjNqFLMmziDC/+cA9RywaBZSSL
KQCZHocfcQM73M/zgWZPL+EQ1P0eRXiz55tdzUXEXqJE+2COjUoOpx8jK9jn
GoULKFXyiuX5H42XdUtCRDnHmbG2gwus8ILws1veUlyUxfcraQeoYXs/ipA4
e7gf8Vy+v+OXu+FciULS0jEEnqY9T2xcJK7Y/Ni3Mzcs4IHAfRA6mj3nbw19
xZqnC2HWmTPWpHHrOKzeki3rD7tKGy0OZ94T5k5Fsu8tlXyQFQM8NBntSTMn
1DqbAsxY411mqYG2K+9kPSHWsuRkoEVpJnDaz75RQ7qcYwzoSb5BsH4ntAFe
TQuCfCCU/4eKjjlH0kX3YDyBKm9uF3UZ6N86qGjVMVgXhRBS0dJcMPrsxYpk
gk4Xauu9iuAKooNdiydCMGAPy24jauFogpcAnWJGeX0WPb8Q8ongV+LXAa4U
yyCGckYTs+w++CCScjHmUIEbgEWTieJK3cqOK1edAxT+/ZiQUTh82xX0qL6n
R7J6lp2Fo15sXHuZ3ztEuhjHlunEnPfjtbwdVNHGt3Yfr3z9N5QDKLvCciZS
G5ZnD2cCBeRD94VaWFt7vbyV67SMofMdH7EJkwAnuhPGJ9B2fydHf8LrBg2J
KgA65uzcEJQLHM6ykWLNXx9BdyvcCw+bJvycNcVTsoegOfBmOI/PAmJTdl/t
WSv6WO9LUrzeh8zD6Xeq/qPoZtJiakw7MD0ISgTho44pWgACIb3Q5rZl6mvA
J5J8oEMdO2mFLhgy0C7QzbCHArHKrUiIn7UKb2rxj4kscQqWlOXrLEsJk9ZX
KnAGfYYVQT5YGH8TJxX+AfsWXPhmyCJh8UODRWWIuY7cI0lY+sF+mhbcX3lx
CdcXgpdUX+1AZUVgHP36jqk0Gg5J1juhBayTYKlzw4kcxwtZqgGUsji7VPOI
hf3ewJU7PId8rgytiwczLy0s0TAQkFhyGPox3XTe8kc3nPQeGc3NrovOspZX
mXDQXWfgLGK3hqHYq/jWXPNUGiv3T2FhVzpv3/ayCVEnco2/GqJPK9WdRCpr
olWODA/cDWYnhENZSY3Fof7U1dWtIaBlCehBO+ZwXF56r7AgYdmwmtiGt4Zd
jehwYB8CSD1TGVgB5U6sAW9Und2Llq/DHS1H331+Rv7hCWmQ9zbPrflDZrJn
un/u97W21lKUP1e25Bv9VWbVoJNEA6Wa4qt0I959mieTSYZLXXky8g0/wj1Q
jMhZEpwpfikVX5he7SrdLo1qFbRqHaIhtUz8tLSE43IhPM5TEEgrxgF/E3H6
RxSjyYx0mNGGOVcHh+3ODI1v+y6mqQovuOJPU5qn035db4M+BVhr90Uq3JCt
wELgEpJXAzjpy2+dwOZ1FUVVt0DSepFb3VNoRSxi+fEISJx0NDD2KRGLsuUz
o2Jfe6frinJ9OV9VSsNaxEPDZc18vVy0D/YdiszDKcrOYqioxr60U7VKJ4Yv
6A8UQ19VIXFvilIkxkByvg9vYOylnLw1jCLo0nPseLHCQ2wTv9X4vdBvcd1d
ziVWBlPdARFUsTWOUcY5bp/LeAbLr+ZPU/0nq963Pq19u+FJU+GNqZqOmj2C
Z+mxm21Qlc2PhWBekcQJWDVx+pPGdS9oy9K39CPdfAJiLbGNeJiA9Ob7edRY
MYFzJpHAgnDvHcxulDN8CCplOooMHA4ZnOgvCDNbToN5l21SZkOJmVIqfbQn
2kQiuPKcDtVPDoLGn/pi0eze2LbJ/++eSUOpR/j6bEG4uq2JT5wEsY4W/v9F
GfucmVI34eQmaLCf83D4K8Ru9eSpzAu2RVSkqEVTBBoYATpeIauBIHkAF2Lh
baRL1/SWyd2PH0NskmWLb8hlm5LSOmDU3rjXFkXLmpsU2RmqjUWQlkffxqxz
MAGbDEM2uOo6mWAMJ6OH0ymZ81kVBWW+SoZNb+tThFjJcRdSbMtnr90db8/f
AJwnJj67P0RILuhDlaTBoQl0WiIwpFM8BghTBysZvzgdYsQimH761xX/2Le6
IZevWjFYjZLR6CEnpmu99BVKb2F6BKU+SAwc6mmXh9q0hnWNBp0urJ56DnIl
qYdXSXEKoDKY2wJVgBm+e9oDqV6mv14WqxWwwYwb4uZrQOYDw82ytNEoTdlA
i571TOxYTnpHlQJWXFHc2cvSlzeWJnmxaPWvwdyiWLogxVEkce7AC7kRzhd5
FETpQsaT5mnn3Q0jwqXDBeUsaz2xpq4qCdd7FiaYN6qc8Qu+ONsaulCxbwHY
29GSZGAZRq+WPUq/5kKjomFOYSZ5/kns/Wqz7qQGJkimK+Au9CyJ3C8A71oK
MNFhC0nxwmbgO2BKzEF6Z2kCGFfxkTmx2H1Jb40gVFXGxxAwmjHUaVxwNEJs
h+O7Q7d8vA0B5j9DsdNWI2zrSAoJx3BI8qtcGk2i0/9HVrLWfUI9zaQ/t8t5
USoANHejpRgUmpZg1+UWCaHd5hMRUDBXG9G2eaRV5DYoBRyKP6A4ano/Hv6D
me8LWuaoJn5CBEbGOa+kH+fIm8VdRDEOiFmXFbxX8o9UkHf5n8ep2/XA80b+
fBPqdTcBwV5fOMEXLzt4JFnU2b2L9yDAdMohFlovJtsS63y42J1shZOoeYsH
/TldcToqI9QCMN/N30cqTk/Ea6Kw6BaMc5Dq5uq1QkE/qRLeToEDSDxmzNVq
rqSinTNegxqwrMEWDuM7NMsNaSv23Lc7SQFADwylm78Tm0FvZalMWOMpA99b
IdgQHY8HkjKsPcjjuEIYPYPzQS2QmsNn7w2QAgjMMCpKGsriV6LfOoxeztcZ
IU3U2slV5Mr07p9iL5aHEOffe2u6fq4uqVAk+XkXAt5+UNde80mgyG05/K1l
S1RK5Lu4f62Ch9JB+h7Rm55eBO/YaksvjpSS0ajs7eMMfOUkSXEvoj/D6DWK
KQGnVf4GQc96yB6D09H+riRnHUFSrFiw8qA2t9Ql1R8H1agdnkixvAFsnDu3
jCBfxb0wRAGt1T3yKxXNL5LSaq3LcQxGejO3OkPKlfDMitPHgJdByVT4oBLG
8uRo4XsMuHBphLJkI7xud9d9DrxPMBMnvlsMaTqYAy7Vy/rpXzgB7jug9fPO
/bvk/PKp1Hbfy6/uBj+EuG1UXkgf9E8JByPczhhAR03yuop8one07ztv2CVc
R4rW7ie6mzviIE1ZTBYBIduLyx/JPym2OMynZZaYQrHe8uh2Qa8PjYlD/vTC
vjsjtSLQbzwuB5ALBKZfRFsFi6LWCiHuFMeeYbB0XQPbu3oUmVsO24R5EZTC
PmmNYf20JqW5y/jUT32W1ZOiOpxK3u97Yx368hEw1sCeZYtdxdZ7MVeeulmM
42K6gn3tO0JTbbdIeOX/x76/p8/RwsvOGRdAVU9rIkrQ5OXfZTs7Cd0ZrX6b
xj+LM+Bcsok6ZZL4DyaHwpcOV5UIsVHwhZ+08G/CaTR3KY2NLwh07XVVxXcw
n0AjhAUuz821yFtocN3O6UiC3FhzdHZGmqGY5SMhsVU7FLXBNUNRF0AF6K/b
hnxfudJXyL8GrkZGKW42P4gcjHqp68EsKXQukn5lb6950UqIZfqnfJ+r9zh1
8oClqtXf6nrQiMsK8KWEj09Z58A0DV50Kf7oTc7Rtk0qlN50Nm35oUnsyRD3
KPWmELTj+6MOnvsG+c7Dhlvzj7UM4L8Q/Dz54c8f7a45ZZgI20leuGQ0pqhS
lR4uW2dFdVx3tupr2psojmqpZ9sKeE90LdbgCbZvntV2lbjesMTl5hWCEvTl
7yAQ82LPC2GgSU3j+jZZ2RTihOODc5Bht/TwRC0ykdYILGD9ojmPIGInxE4t
3S8nraGnhq9tv6csy18zuhpmYxpZXHVLLhvZmcuSIXoiWz8xNiX6GlV0og5m
eq0Fjj5A0BlOEZW2tkxq8Ym6CsUV8IYQP2MelVHbKpAugpyZZv4E5btN2IDn
nnaYYDNFlgRx+getgnS67dcRsRRivg+HdY6N/zWMb0jbFgDQ3ZQBjCSgLVz0
EGOZPY0Vr7SCm134sf69QLxw6sM3q32UEtn9la3rGhYKXfoCDfhzdCsjzDRz
3Avo15aHlCgmxX71/Plr3KoTmnU8cMAbtmDkZQ3EdMcyayvJSbTikSeSpuiB
iWwexuDwbY+N5OUUna8ObOYcHfv3vAoBNs0BKIkOMKY56SxP/xUPLHhuM2B5
X+4AClNOdy2X6JcJ/oCGY/MB3JYNMsVNoeBgYqNJJbm5wANkk0azfLQeR6VB
28Tb5zbFaE/AukzctzbHHS13mwzxA9KhV9lpivLLW/UAOJ9fp2he35yko45G
1BuyrI56cUTNEJ2rvVE3lmkV5XsJ1slrFKbqc4PttRA5YG2RisnLrOPw66n6
qIIiZWLv3pSRYDrcvXmlykBBpo13+Y7Qrpe76kcYQrkuviPJGGz+XmTn6gK9
AJnSAoXiB5nxzTKyFcC7IwgEC005cyenZbOgkyfc846dQ7cEEGL6IKY34xdS
xTZX1ManPt/aEacLMEuy5Z6mh62Gn5NbjhkfMJ6MnWJHincJvONv/uoPFlbG
KIzrXpfzqqygg5Vtt+QNOidZ4dB2IPYGc99wlv5awCgIUFT7oyASd6QO1gyY
6pduys2hOcenl+m6lTMfh0RXSoPg2SPtU9uTCRtAuch2diVzzpWzmu2ZDk3k
8/k3qhQBa82bOuY5ccEOeK4+Ldk8ybSe8dUqLShCMhsSTOPyffRyg0h1PZWg
mk/y1CAJvygW+akBqQGs19yDtZYfiYJGAvAnvwFYTSBYSa/M2aTv7aZW1ZOJ
jJ9hmKU2Bw0uNcqa+iRJNXgnu64/Nitbk9dcowdlbk43WWv4k6f23pHZBIT+
JCD0s1WztKPpF4xxgP2dDdJdd3oUGR7ShM4P6gy50yHlvkqFFyLeboAOe2h4
DpLSHcaFXJbOmiL0NSfLMiEodNSeLUjkQDt/YSyNzeq8Hs/iOsD3iizrbAn4
M7xddohvLuzFvXacBd3bNKZ5v35NyQ3yC2TkNr9rBuwAom5SkPr91PLx62eY
07pMG6OtjcfCfKvQsgtCkEhL+n80FbcYOHo220+Ni6qwXsrYdLbiID+bcahX
Ssq6ngn/utQXsTjRyh4rILrzAWjgWjnYUic7Y7W9IGk+0TsyqPcepuiody7R
VjqvjDuveE/yDULp4A2V177INdmkSZagmzYWqK+VQaovyy18hBw1Q8UYUvXS
f7PYoTL7ZCCwiuJgu1hOHHhOEXQ/q4NXfkZ5AqIk1rIquyHXpwJte8bDutY/
dc+0LBUO+y+GtncU7y3mylrAQCFDem8O6y6MbhkKYCrvFv5sdz+v9BhAQ789
ID2AiDIP8q805ExV21SY9e4kNti0U0zjt6nfE7J2XfVLK7TZT/mvL/N+Bfx+
3JR8NyMlzETRF4GI3s2cu3x7606dLLJ/2yxrHE5M3EbUSKRJim3/5FfxdY7P
dVvzUrwMperNnkIkWnahHU4CFWqJ2YxooR0lieQS7K9hD2gJyRtkbhSrWEZv
1n2ISqvs4b0Q5uWpUJHsmGTNz8ki0zr3Yhwdb41SPe3bLohnhX07eqTCHdOk
GOue3ELlO2FwbS8g0B/hL3GHazNe0KCto/HQ9Gg7ZUbodg8+Dq28xnXeHqoB
V0jKHFSE7ubat7cbYonI/OtbzNHNDvxSVewSKYiTyn+1HSAP7O8OHKj50RCo
nITBqvKYTflXymfZFljwePo2Qo9LKGbP54Czkx8nZhv0Yf0kmNPnv3wZkEXP
g/5UP23+84RL6pI7yJikB+53NNzPwgpZOr7ZJ+JkSKX6Ot/7pxTO83nGkDon
VpE8FZ3GvASPWqwPc/oiLNkqn/A3Mrsaxij57oiaiQZ1++mC/9mzbpSV88qL
OPpnVF2U/sPUlk0LsVXkv3LrNY62ybqabbR07IdA1iF4fFfzkv9PF99rsQeO
nZFWUZqETB4oPIP70h79gm0e6LwMWvKgqv85f0PB8hcx9fCB4pNJ0HGTAQp/
9ciwbtLf6JUZzjAIhwVFyjbmygNcPrU+0CAg6yKdKoNC8Z2lzLrVLMZIr51M
p0dG+1WVt7eqY4X4LBFUDFkZIXTFwYp+zfTIQYb8qgw8W95B9EmITR78h+4q
7pcDkf3o9XjRdToxeU4hz6GSlGNrceq5SuACzh1UaFeWBpcYgzbr8PA66PbB
k1h6EWlqmkpmeQr6agklEWeoHIhpNG5LMJT64YbjsAzCsuVMDKSXi+MIkotN
DLu50DfUBimbTwC/7GONVHfdK8RUXGX3q0ycQYL/cYuNoLYM+jhD6X0Ucd1I
qYlqWcDZR7xhy5pQFm498nNRbkhpwD1VxLS7fn629ZLsPcZ/JYYZXsLEJotl
ILEtWmKhtTa3HqWcLVYcavgeIJrdoyBcQceMgykrmGm7syYW9oIbevVO6yJ7
jRP087cxnB7PMsPNV9qhJINRRN8hCefgpJi7H6PyFqgNjt6mkCI5Zs3Jw+Bw
3he6W7tD+390q9LHIFrrNzxhYxgtaGf0OntNT/vYggWT0pNScIA/ZuzXmKNu
R3WFOYZc16hp9bO3WmCdNObahhJnALFJtNDokeR3S2lgNfyDJZcAvQHWx2le
Z5gxBh0duos6vgBTxiUIlfVUBENv1/PE04N4ZcuGU4StV6GN/E4LbZJRQY/A
0BQcF2wqWsafEdTGvMaXujKj+/ukYUFfFLhm0aKN6tpggUPvBtooif0qkNUh
xZ9gYXPbrLFhXyo8IQDwTQeXQ1eWdXlI0lluIZcXDS0NYQRJEwio7LmA99CK
gtPvntDLJAXZl9uH9a/JXnoVyy5RjOH2q7f5iQQWnc6XpvRIWsDN1IHbnF3p
FIeFibKkOEefehcsc0DIFyK0FSeRzYYt/IRMVIAmSJhIBC2RaCMC83CmKsWB
O2q0mh7I8JrpXzC2aMxuehlQ0QzN9JoC14pu8mo0tRO2TrquIIfgC3VmUADF
Rsd3vG5KnkBfWN28kT00cZBKq4Jts+iZ0G5NyJZA3HEALt/UeHaSSehBFujT
W6XC7Fzj9lG1q4y+J096LWSaQGpTqmqm/sIqiApDAaTLYeCfc/dGs96BReau
L8mT+5eOm/adRhxEra5QMrtWHsbk9aSPBsqPX+87G6/ROm3JGp/2y7D4isKv
ew1EtocCpBhNXmn++5Se7VindBDJtEN6n4MaHvqxLwFK4JOMOx8TRSTS0Cy+
6BEX05morM8Xym8+dvyxj1yscNVrpiVAYjbjyFvQnR3r+nielGBnZ0wasZ5Y
h5bLFGXJaE/TNk12EyYWIX1C+XA5ryzg1E2+9SZxpT3Ahef59PTiv+QapXFM
Iq/4vchd06fVdN/FswwP7ZkVlegk1ywmpAg3vfBDtdClbKPyoTgX8yPVZB3y
1HjHTkm2IaK5o1JOVQ5qvNZiqu74jZD9qZJRsbYPagp2mVII3KxrhqrFclU6
vfCREJiLiL0PIF3A4qPFYzJsk5ggd0For3ppX/Os+WLUipfNbrPFcBVYjXRE
vqkM4ULXm5/gtm81umzYihbZJ/edXZKQbnzblhdbp6/NcP2gdBx2tCcF9FVa
qwBGm73T4whTO10ddG5GoLV9CZCJTYvNsAsuX8ZaMs7VmzWAUfM1zv8AgLR8
YS01Y5sqSl6VvEyJO9lO1in8F+7Ij1Fq2Y3BrI7eMqLsM78jIaAkpjoX+bnB
FtVVzra0//pbpI6J/CqMCwKQUWMELy4khmFPKHA4JMZgiFeRqTL0SC5MtaQI
eyyPIpFRCNZeXyPASMp1w5hL84b71E4afKK3EF5J8VNN3956Hb8XB3WVQKBB
g0lmKErshD/y2EonLpw6reqG/I8E/F49UwVdWvbwuwnr4jTSu9906tU6zCQR
fLbl+azkfq5Oqo3FN1m6FWf8Ni0DlVzaW4tVe7giDbXz5Yx5vOH/N/aJdbaW
/T9YgfV6KQG9GVABiQeJvGYUEUOEH+6wWxyYSJu7tkfHyFqPPqIvKvg3TP70
jp3AJOVKDrkCbxIp87tR6plzrgGX5FIsKY4S0ZN0nPiJX7zN/7ZHI8Nz5k6O
0711ZlAtKwu8gJVRNhNllzkuzNCO877Woy5psHeBS17qpWd2FVXIZQGVclz8
eyA5UMp8GR6+D/DooM2cNx/evYAgkDNBNRf7Cnx98hXRD1sWzpKzYC/xZ9/k
NlzLMnJOSibuyJF9S01FoQUt60c1Dg52pRXaEa4JkDJpcdC3aIJANLHwMvfZ
ZjCa5NzHzDxAgnwtXERRFAezLnY3eKqytOWmJgRgHppePLhDjTq3rrNwKTng
r0U8jvVROKCjNn4KS3+LloombsrY/iYOX4lOw6Y2Gjstu2Z7vYxN8WVlGnoo
KyDeqffgnDk4kh+MH2aYOrHjWlSqOVfqYm/clswGw9Kbk9cRQIJKr0hSINhw
tefMSK4wu952tCmvzN2q2IEDsethriPzd6w5wo8FFkN2A8iX+kepsBUwt//p
8ZfedPS/U/uR6AjxGiYm3WX0GmfNUsQ9sWARLYrxh+SH0d52IMcjAuH1nsPD
dMFtfhg1nqwJG5oLgKD9FthSW3/EZdkUGrmkdNaOqu5xMQXRj+yxQjwCHj1A
UcSoHjZzocTAyaRZftHRYhgbt2GCEO6kc6wQAaCwpzfxb3hTdmPLFHoyEFgt
7TsQircrHXEAQXkFyu0UhxFgXaUfdScJh+jtM+x3ep0mhXAKHWhIYX+sV/5S
2cuNf/HgqISkGJ1hoyt89H9d4mcxSr0IdJI5C0eQnbaUOWRDeNmXpHg4e9FP
if8/nkRZiZs6ZSGGmYf1Ci01Asp1LF2Z4qwfgl7XWUZZNxrZdMU38xB3zn1o
LFzqP26B41vxccZWQQEGsgFphq41KKjwnGXzbgPVewPciwGC9XKaknEdyKzB
Qx1POXdJLkOXeku9QF7rss21xJanRv0B1gCTRUkHj5Y8iySoiqD5ub8G6JrM
5pMbFwOcCh/WULjvvmK/9y32eoIVIGYnnx6Y+J3mzQ28+dvwkObB4MzcrLS0
/fvJarcS+G2IovvVbri6ZUodxtOBDuRRlOXgjKWjJBw1tzpVzEWgS3ZOeY08
u3vq0mp/lKROHeLJHxrM+BNSDEHWr0lV66DryVMc8ScKpaSTz01yOz7bLHsr
4bw9j9K5/bpW/aQq/Jz32GeVTRIUwxH3qTX9XQj2mnYhfjp6c/tMO9viuBcB
eMHeSDvzD1ZFsa6W9kTShgmGb/zWAbxhddshBzoOFb78kyT/jP+FZgeig2F3
D4SDQ9/jHmcf4t3nkh1PnrSBRFY2mnaY2wQc1uOFjEqjk0EFNA9GwLqtRal6
0vTc/MikaB3iDaxd8o8C9VI/WQALnoQWyxa6ERRLIir1SINYMJw82nqeU5u/
0lYPyRed7+HCN5gimw4CZPitkg5bwDfpFyUZmY9LIxpTl5Y/0t3UcmagYDDJ
DW+wSvmcnP3wMAjfKOIqL8o+twJV7iI7hS10W+QqCQkDdmIZZvQMzT5Lzm5Q
WrFGl11+ySDAgjM605w0sF8rRp4tTm4QwzpfXcLh2Ts4Ctw7BvRp6n7VRhSk
uJgo3jUyHQshhww2qy7sKnX2Hjn4HGKMeUKD4grhyEr8b/4JQ4j2oYIQgB6A
EwKC0bSn6JGnChEPx8dMFFPNMfM42Q1b5FyAfPuFziftEKws74hnUOZM1i4i
BKNc9iwXEuD/AjGL6QiPGmk7aunUU5JPCLYykSq4fbIlS5c+ob2PVrHMn+jv
7xY2Re94Ly/4osNXQfX5yIu28mXylJInUzF0LOe59sh6A0q1KMCueS7t+6V6
h86Rv25n7vOVWXKjcyhBHF6rqjNvXYh7Lj5gxEHMrHef9gAoMeTW0IEakepZ
g5C2C8R4EcSSsVbzZA4hsz/1ssH9eaqS/PmNuHbOCEy1Dwq/kigkRShAFrUO
UTHfUo8nnM97mKq8k3szx33eV278ZF7E75E10sqL+28xIyCu/BNZiCnQ5MNR
edgO/WjmfZLaxCAmSiYri+11LxusF4HQoxr7rX1/C1SpkaVJD+t3/W4e/bRr
8PtU6r5E/Xlyb10gqLd4Y42i7Kh/4EZQrPJevP4GBp8DHDMVz69y83LeHjb6
t3IhozWVV2HOrGGE8eewTYB9gG903G+hfnGWABO1Rj1sqWLrk8Z04bhr4Y+N
dKfhac7vPIyXQsNLYyEG2obhUPPO7Ka6POJbU0/DiLiBlBd88I+CTggUi4mM
YLzXmgfHoJt76arhISuukYx1xITGt3rkCye8f3a4gF+4SXSnpd3RqDTIq4kC
xfwo2KEQ/SlYl9e818svj+Oag4EAaxNllu3cDnkqtPzOE3N+AwZXtj9+5p7x
zVSL7KoHgvRSBLpywmOPYya7U5l2bHRQS1Iemml08LCFxrZY5uuy1Nc8rJ7u
7/n1+yTSE8KVw3qEMhyuCXWPkLTR1Y4YYuepSbL7aSaJ0a5yMiGChtMp1F+m
M8L5XxQ/OLRGRghTelX65SBKHhZppUCabNUgesGtcMOfmen9SZ056LOXOnLB
GQUkCJVOjT5WfBvRI/xmrs80FFUmKWY88YN1NRI6RraqovNavAbWxsbHC2FG
eNz/0XZlE+oK8GVigICmHTQRS7XLoyBTqMVHDNI1glwiDx3njnlxU6ICDk0K
W1SMcnNC7SnWWsa0WOBsIvenuZV4nDI32K5BqTtvDfPIht2LAlSpnvQidbRk
thjwEo4627x1jwv5mqOasIyvh2kHQtVrsgQnt3HcX4q1DQvnU9H/y3fYmjYm
AvTovrmNt/Hpj/g/c+8s0euEnRiU+JVjVduj1II+Tk/gJJTg7eSk8TXbpn+j
Fyr5mHlRJ5JDUtWLg1xci4I8KcndebIH57HOy8Wn8h+RR8WCl47R4bAYh/ca
g5NmsHSC4hIoJWP8/PLGC9I0cCU98Hdg4kUJbsUaZuMEBKIJ8ag7A8ko2WaG
GajsRd9W1OMSk+Sar/hdYzASVOHhlQfanLBx7WrHfmAf1B9OqdXMzPhylm3t
0MBWRuBL61y507i3qTnXFhBm6sTn9F/NNMNzBnsGgD6rrSIBBBt8MRs2mjzd
sEikLzW9noE4xdCfBVA9R5548PRtR/Shs0VG8WOSdy1W3q2lEZlPtKRbzdBQ
0yDaneHqRfwYC0RECz2sV/jDT+QhDgv1+jGE+OTwgC7hXfR8lZp9fdAZPiz1
Emh/d4eEy/2xE1Wob+Ieroo9pt+x3hGUS4gCD2Ef2yvxMnxyWBnJxb8FyUlo
6yix8yZ+tg9XbXcnUDvPGD5ibGsZOCNfOIot4nktO6MZIW4w4FBak2zUrYdJ
7P6S4lyEgI/fKvirhQH+bbvqano/EQhU0275IK0jpSqCz4m1MmrnW5ofCL7O
5h0cYgSFeVN0cCCe/TRuRU8vrMY00nZzybBlSTLcnSizUEh8wCutSclAh2/G
eYV4ZhtGejKZ4ZuRQT7cgwb+a1sDnLdq2JQDCG9rYjKbQZlZAp4y7HkTAhUi
oH8gV3Lcqm8iUxwwMCx/EAUfSjFgBSs4PjvqizmEUNGZHNHZKPqpjnyB7J09
UUFnqtT9LKTf5joaU/TaQopG5rCqoJRsRVzVlLzN0N4DivkijDtF+YHFrkqd
AhHe3cMX3YsoVtOXyrdXD3csXuk+S+ilONwotCOZaeCTguIlrwyDDokoR8YS
edaEzcLIRVJX6+2hE6M4pUs8CKe0Nt023w2hDaH5w4oVWEopJezyc5PGIkIY
7vY+XKDOfS8fhImqZbI4AsO93//fM2Ipt+aAh0J/ICpF3pDad9K3nAY9vi0f
d35kxBAIo8yw9kxpEDSW/S9DwuAJhQjHK7oUNDLM3FPx2l0qJAz2TtJoQkrM
KXDoIHM+9YHlNpLjjrEwdFzmmE7G4ft6xbxLnp4pqQzAy/Rt1SFsF4I7p93Z
6wKKCbxlZ+CZ83CmpdmW0yZ3vprvaDoNILTSIIHUmcqnDFjhQriBrvYpgYyR
+26wztg+2H4tk9Q4J9RCA6jxRwBgTdJQQNgWl+16UjlXFglIfhte2+ic8pas
uI0TPhMpMpSXDo1i3l+cFWwLXAaq756EKbdfIAUIO8Coc5euA4bUHdhxjLg2
5/NSIKGSlz2Dwgm1cJijFzQwW7NKkWGgpmeBFfZa5poOmVq1YZkl/6csK/t4
Pnc8Ac7uhW9L3dx2dwNzHKBm7CeQ6y9raL3dBh6O6vcHD+MyK7DMtc6VKC2t
FPunEBZx3MtPLaWNXZI09fvoRWOVz/699p2Wx1OZPWbApDzbWiCQlo/vQTIp
71U2+C9XZGGzsD6TqMFfjYyccekPhaSpZY1rd6D7FrPceeg1qdtmqaQ/0UkU
sEEiSZ2tzIPmbeyAdyiFlefxV5Bxq4hCT4Kk57bKfB8On8BzHhfA91ynL2q8
DbsVw9f/AzOtl7RXwov9IxcQmg15gVjABsTNexk0Y9rWaRmu70Z4kQdhklgb
eyrRvtYtxHJ88dTD7CYOZmva8wh+MmJ1qyyLy4Y0h1fCkORVzfYBg3T8s28i
5iNJjzz7ud6sPjoCTolpzCapyzpi2nDT+v782MO9pw5K+EkPnBY3QD6vHWpN
kY09uHSe9H5LsXjoq/j4JJ/Pf9UUx6nIrccpJz4bKD2yo0Odb06x19LPCA6t
CV9kmIt/pTUy4StzqdH2fC2GsANDHcMjUQUAkYcqa+uLP6zOZLU7OBd9y9sA
AM+RE1Lf0erQ5RjZloE1aw3Jn1DLZjuWC2iN9LmbHzRpGdVAfEJglbyfV+dA
2ZvpFanZZcWhlXREow0nX9/ctH0HIRSItD15a8DVITOyTa5qSLeOkKhPWArO
8RHcSYyHDH/2prnQMQku88q6mnzgKM+1nP8BqvKa+jrfSAe4FKSFWkRsju1j
RO6WomQm1/ukNB1DE7UjRz7ZbDkaGuqXmUdpIbiByvLJoX5GsovzZs8vV9nx
J3srw60XyZuztOCWap3Bl8I8GNBZK7TIDyUV00o73f+vqoNpw+bJ68Oa6oxp
AA57Lp56IlF4qn8VkXHVGmkDR2MxAFkd+2cUh8E8fzkHFzWBF20PV+sLdO83
msbV9qiahVPz5qpc6FeKnERCSB8DeNsjnBE38rp0UXDT/UqDU/60dBTBTh2J
JYl6vK6YuFtDPWCCPJC2ivAgQkNGqVSprAdzPQfcOgmB5YR28VVkBuLs3WJu
4eIF3Pbipmg+1SxZaZLkK6j0OQgxhH1XXQ4yQu8Cd+/CULBOjLduWIX2CeOj
ryPdFsXOJs1ClpEbOOPOTWmQaihSf0qjXAv9EEQVuBeRDCTuoZLGrwDGxnB9
i3kFyHbHqeZ5XB9tOP+J95iTLxL71ErYWdurEwOuq0MYqB6evHS9sXeu21K5
u6gJDtVfwDUcBlzVxwqk+jhf24GLIiAMVSFjeNL7QwOsn68h2rOICPjVxTb9
RP7+zkzHFyd78xWixxy/mselxAEu9Nq9dTZKtPiPwfxlWKSazLSAMBtPF+xk
xHvsvUUXNXjEIaEqb8lad8Sv304wnYzQB93QmkbXbOWqSC8ExekDK2Nemmaw
1DGUXZ0nD7eZazz5721yciUR/8Px/lzDIFXE8O6sYSIx7Z+9z/gD9R1SqvBM
9y9yCqwqtUlsbF6wQ4hzXhKQVSpFG8KbJNF7l3CjCmlryECPYGD7RK4z8du8
HKpUPuP4141xJobsQdBMSkH2AdGy4vnTY6gbRxFCDIMrflswBouQZlpcFpGA
WDOhtebwYSFeuhfkAj1wZPRx0FBhYn0OdBpF4Jckyo1G8nGolCS7QpltqE/Z
SPBvGnrMjILHtPB7DRe0sW3SYFNUBu7HZWzGTtw/REU4d9OOB0Mr+Z+Hihwz
jssyngNy2RzfNjeYWS/v1sGAGQtr7rzJh+V5trO6uiuEazrDhHVvMYmvTOpV
z7Gjm2dKtNECTh/REtUuvLDkVqUFl50zpr0b8Lxgh9odUrIRGMO8NQcP3ZIa
G03jRybI23CsvWxsfwNH6OyxIXHekLLBWniAU7H/NvFvznMfcTFig/1Qnm4a
L47UEsZxduI2S/3/cNYl+RAxtFD4LD4xreexgBFp4xCes0WxTus8jt5IlPUT
q9fWT13TkEWg6bQ+Rmjx9HzQbIbbJjHDt0BM/XHxrThRyUM4oraaQMA176BI
4z28BsPKAgDPqUCAB+vtiQ/QF2XAemd2kqAMhlJP8gdAIpo6hb/Z+Em85xdo
yVRw00J1xXQF5zdF26X+wy8oR7mABGmBlZzqD2CJkIS4bgCQNxqW9pyWCq7m
Y2Oel2Pz6aUsfIl8iCf1L4aYPmPXXDbYBptQ9858j/hkV3Bxh//V0boMkZNJ
4p7Zyqy+H/YD431FgbvAWvmpXLyKTR6Phbc/kAx6V/PQCvJuVzrDTgjIoeo4
23r0lfobwB7nl5El71reypk++yLL0zrwvgVSFkwYK26JebfdH/tr+RucU/C7
WMg9ZIAgW22svfZTq/U+UGWWSdfUP3HLw/AZEq+ld9R3x2svAWsO/wJiowh+
xFrLLv5wIfGW1/sePAXfA98AomCAZeI+189aVFxhOKBKRx9fNR15wm0sd59b
Taf7ZU3K0+uJChK5RCdy+q/LUTHb7kbvPGd80pO5GOc/IXafXnSSGiad6UzB
m5xL8TE797ETgm+NezihwJNUtwNgKN9BazlDzcZK1ykQZ4aKBjScSJKwRECt
Lwq7pLxWIjAjR3RfC/UGt4Gijp6G+8ALF9UyJFQU/K0n1AgXr6nNdIGEmKd6
cond7W1bdorP4bct6RO9ZJOGzilJ2dTx4C9UnFx7/lnDCvaMMCwMfPXOH9HB
jWl2+65KWLz072KQ8sOn6hax1RmK5/hK2i6n3oH8hHPk59agHgLmjBdoR295
qIc8IxRRn2P+Ia848pSUNnzLbGTvE3kvycihh9SQnIzQ6H0tT8nz3/sUFxHC
pD0YSA10AaUXWwOFVfHMUC75QsANHwasn5RiH0IUhtRAUdKXN+FvA6AQdZpk
671QIJ4U4AMmwHuYjuXea1wlfcBzPDKkKpV6nSsWcr5ff2IGbaHlWGBp1EWc
Ygv3mYJD037lBlBYNsXYomE0BksdA9TWkv4Li0POWWm7QRUEnymPjm1RNv1d
NnZd80joy8WOAC10Opt9tL/4bY863VBkuoeiBGtN+kcnEgsZHbNd+eZSqSmG
t6TLuTO/wwgkVNwVJ0aNuwMoXax9y8cB0FVCRB9UxHOXj9VsNwtWOKkhOd08
UpS6c01OPFlUn4hiZez38vfD0zfS/JlwY5mDJZzsmaPuM2V6kXFt5sEu6hUb
KHSSwdrY0OnR2yaAS1CCpNnK70ddqmXx4IY/Sv6ikl3cMHu3NoPg9g57/ma/
UWA+eMxkumz41RlsLrXOxbB3UIk4HgWf8SvXYNEpxp8FcVFcnK9Qq6vQHZj1
bxsz0pJCHbxFLlkhXWtDAS2amqkb9Pq65x1cBzgIl4fHPqRhhfHVEOy8aFpI
YXIe3gwn41Y3J2xC8JVftsMk6P7PCyQfPldEibRBNudlSw8hkpl/XATqsONn
/YUIqvFUYbrqG2XCCis/4AxafduWTVM8kt3EvaYUhquqarB9gdrXzJEiRK2I
KnDEj0h2n/2e+MAzbzf5iBrtCsjNeyHn/4gtYGgel+QDL/qSHGdhYXy+rLRh
eAP8Jp25E+diC209+1ya2xS81Kiz32pnbIgcSeeNsOhXOLSbC29xcyKnvWnw
IwpjLDFSVKerNPV/QggMflFFpOPeR8NIv9pAR5p5pXoYT5hba8FM/cpVduDe
byHPQ2sOqxi1KSst7k21XzwVDfXDaL5G1O3jrSmWzLDdlJiTV7PAx/AsU7Fl
iESjwMpm2/509vUgom8xmrQC7IsAi74VA7mi0yW6Gg4WxfTyHyrao2f0pcuq
lvY3C0irmum+KY77HaQfh+4Uf14Rjc6kLnO8KrobRjGUXb/bd+6u0nv9SC6X
+pVjvQ4AZSmN1pYSHMY0+TwkHpivutqcjTuDhBklYcvdH7/xjcpWHf8huhyn
xiAMtys4gDLzLQNP+B06BiWeCjEfZlYxOETKwkJnOJjjQ9iHsut/Eol22o16
SkYsq39HUMRDjhJZ2yGvyE4FLPx8LzY5R+69qvCcip72Q5/gGui+2W4t+dlQ
k8kU78VzhTcqSOakGMJgA819kjrHk0prrgxN33eWeeSX6uGgSB73fuEsuu1A
MD8BpPfkXQKhfORLZ44eS71ZjyWYns85qPhEfxZ4FADOLtS49maY8FJA81UA
INaZxp+zdiFzEbwe/Nd/Z8pjqx5sNrKIMH2zVK8oG8ojpCmFoJk81/4puegh
DjAoaRtX8FQvTdZfB++kX7JsCAr7YEupATMEF7/+zTdVdxfbQs/cFpiWkwdU
1K159QjXpNBgssizLPGfdlaZCpCZuU+a/RdxcZxJbA9igxk4+81bdBBO7REL
NrO+UHLJ6vi8FhwYWZlfK1/HESE311rW6FyLNHa/DdtgV0gRqFj9gmgw8zwS
0OMEu3Y4wI7a0LBNiI/x8Xp+/oZ8dNqAtY6LIKNSrZ2wT/2z8mKiuQqMkB/t
ex/ORgSXYfpsPS3dRJ6PgcBdl/X/BIhEbFxadL034nXJ+EvK9M8KktelXnxB
BZx843TqLxFP2B84eBSpqLVw3pAsNsze16c9Akv/xfvIqezcmmE4SQgtdIKS
/XFpGJe/KeoLDR8DnrgG4lweyAWKuT3LRQCfv2VB3oItGb3eFCNFzchUNN/J
/9h5Q5y6KpDNHcIS39Ou6AzYED+oS797yie3PfiacK1JI+gdrBnONID+UKUp
79zut+hqo06CRETnfGAH/pRHjZqx5Rr9LnJn6ngPXS4+8i9UO0BrNIzpgjqb
/LgEI+AAVaq6/Jww05IkJ4/QHvQnHFSq6SqJ2AjGT8kAlWgBr2rVhS4ZgTaU
dZqKZZBqbhu9FYQA1uf1A5VG+wwfXRodwQfLg8gqj0bz73YA7yrGfkbGdEq8
QSkat2BHYPXD1h/lNjErLsWsKHhkl39HhEXuncod2YQfHdBUXqacHbd6RKxo
0G+yQ5rqK4zxgyrvE6O+VtOEj0iKoZPI3uI61XdpT8HUxgzXKSME04wgVBEb
j+9Y2Eyvl9bZfBXfvfmpBErwwK8eJNQ0rqqGeBPcgUbv+dqASiSs5TWC50x3
GNPgEoXqlxkeMnMQ8r543BUzU6z67RZmx6KYrRi+r1FIqhY0M01UhB6RJv/N
C3Jtn4cRama4zf/JyNxWTQHiNP4lM7vtFDgQlenXH/iips6ZBBE+iE6RmrJn
gAKlPKCPKrBtDCfvqy5wUDqdXJvKX1IjcrFst5rsgC3haYNZyadObjNeTwNu
TnqgdpUlGKuW2fTU3UQa7JT2Mg2Q9huOIpVjQcsFbvxUKPRyQ2ww0qQ0BwM7
pSiAn5X/Dlmt2TCDnM7wcvjnozXIWrXu8zhO69SbJ33KF52X/0Lz7Zo74BLo
iXf+8k+3Fua3o1kLdQ+Tlir3qFrFsOxorzf9KKnr7yGCyBVWjh8L2pYubOFB
F7ns/I6OAEV8tpDNsR14i0aSKnrkXU+2uNbNELFPPcvXzMD1FxyzorK/d7LV
SvoMWS4on75wGErqTsRBEJ5WVtzL3tTt+mEKDLV6mGJkKRfq3RgTaIHLzDIp
gHN3G3NTDCQmMMi8uKWmFFw24wSboTZhdL7QRdT3EIkqLSGcE8LM/jG8JORy
u/pNv1QEerMKe6L9Z+lJm1XhuNupP3gsrTatAzPXKA6Qh9wC2Z8rESSNcUpY
ihk6I75fj5CEE29XE1dGXhu+WTImso8oEonlUxMfWaaDNL2flMFyRbhRiUPF
gEatxjxV3JRcYdm3d6AjMUjVFkgRcNkfmTNnGWDksXTb75boShvHhB7GUSkU
TrpjCXd/SZ8464f5oJMBrNwSBxkKWyQJslt72HkCFbNo/i49SAMQxm08rCRa
RB6GBTu71N6fyP+mz1GXNmIG0qcy5VYaSwv1kRLdGJ7EUNCXZkm6imdIB93x
eugUfp9rieYoyvUPTPqmJl3B34OT2HaTcljIOeGLXV/RCBg/XpXOLYEjIEnq
DTbuQ/hP/UsAHzMkfScI3n7ABnBc8iu8D/CGI/HMHBhHx6NTY1N9c9/6EWIB
V+lMC47GIZuQ73Jw2d4QW944s87F7GEXhFVlYwNYUQp4+joHMid5EJqFOI6b
TnTjrwPcD1nx+aUIQuX46ip9bAFStdqaKDFMTyKen3fN2Ji+ibaE50M4NnPQ
/iPy29Lb0nPoQrZ0F55kdSg0YVUSHp0/avNrfI6LkJAol3bMjtcf/rZHgUcU
CvJ9VHiU/MFGs8pFIEqtmbkY6m1z8dDyU2BLLiBmXdfPbYEnsU0nC5irN+Ht
eEYV3Z+xwmh1vXaGVRVi145LoDgJcJO74eR9W2qkpxUVarARd4krzSW8mbdY
we5XYJcl3pkLmXP7CF+GLqikSKENEpCA4QoGQZ5nqsIMJaPJsSzrd9+2zDaC
qiTwkAzdDVUzId3cQ5n97RHA4Pqr+RaJk3kPpO0ItgYxKGweCWVfQYpk3hiG
DqsoaaXeayCS7d/+jM6/tMYL3PycethT1HcE3nTpXin2riIC6IwjYqce+LIH
xAnDAdH1riyCvuLJgK9tCMwUrkmzQrX1Vdm4L/MSpeE3lxadbVPqMUL2tJaW
XL8iVaJJleV4ubfrJ1BVpfEf03gfrjDZx/oY+9GWU1dYzKrbWzsKNObDPoPx
HI2OAj3hSyT5dXvjnglv4gkc4lEU84NGWiGL12JW56Frmyd6QTKnghqBUsN3
qaoy/98hObRCbA7fyJBKRr/1vWkcC6liLkmCh+bbPzE0AooFMl7re3hxjPiL
GlukEYsQ1uKN41Uj5S1lpyvd1UliO8i+d/mesIi/Bv3PSCeGoavouMLG9aHP
7r8jpAWUfgEQa+mLb6J6X5kkly5dOsS4Ce2pCQFprCLDInbnZT5SKHpESUWA
18YYWlog5Kv09IQpH1wEKQVQP9rTZhC/lYsuclY4qlp4S21802Ht0f1VHPoa
sED2P58E5OWEHcCBz9hBTbz211IBkFoFlena1gMycQu4YmlLyC6OZgxJjXHS
93qayT+Q9LN+Xr8wOemaDeqGFTrHO2ug9T1lqSJQQS8mEw3Xd5mvK57WiuQD
+2VH3XG6MmrgFmPrb8CPt6LQRoIL8qTosILxyhzUEJYGSD/M6EM3ndUDDF+k
oLfQLWrv3+SDUtMtb+b2of+KjaqmfEhwvUyfhfWxduNUAhT/kFljg6eapZR8
15zeCIHT83Thqa0iYgSDQhmrFuGB6n8OoMzes/nLIfEq3+toeuxab5fvD5qv
Z1a6Dx65pia+PKpctCQ15VW2HDyGmhFRnmfwQTD4h5HmLwMSFMTNLiJC0Vg5
MyN4kAMQbLQqJq/PApu7Fsn7PPLwaWdtG3q4sWvii6uCAlBQD7YcKLNSjx+p
kdCyTqfY/8iM3EOmID/5RVsrnMa0HJ7+CVyYNi+5uhKnT9X41dDTyMWW9ax/
dGAOmdP8zGmuow4JoNQeCuXWs/rklxmrkMI9ViFCJ+3PUXma+EZaWVXrQMvf
SqsEQCMaG743N8YDfExT/sJphniVBp8e6+lNYrPwB911SG9dg0YkqTajhF9n
HR6UuKWBc/CBNgLFxQ83oTIq4biLyg0UBPXJFoso/ccKN1xShGWY+CgjvKQH
x+eG5Opcm5eR9NiHWFgZL8uChsjW2CW9SYjdivboZ1OTHSn18452Tl+gpyVm
AfiicWpdiWdLeb3EEw7aFPO4i176gMywoEAxgN7M1vZEQo05jmr0pVNHqOt+
90gcOvh3uxlEtF7AQQw0Y5WGz044wu2o3lc+mvk4cs6RfxVOkJf1kAq7+oDD
BTM59+Z4MxaCXgk94PA5r+qPgLS0uyWjtn8iTDSuaDgc/R1S7xVN0dOGLaSz
syuQMTUYiHMN6ZrX2Qcc919qhgTIf2GizOqSqJf53XNdQ/YMsOJVXZr81DxK
9IY03nx6jkFTC+JeWT+qMdboe7rzsCMoEvixirOc8uRyM5C3hrYLVenB4zIM
oLOf4+x0Is0P47e7ll3KT5+22MY+dIAS0oIHTByQcHL/NagtWclL2zuJbngQ
xEQtaLfCxWK8kN299oUSSzfQVoEzVjOkhGsOLdDCHUKnrCAQeyvnQ5AlZzbk
sOEVZKzrxov78G5BOBDpnB+GckexVNKUIUVBVmB+vViLGn8WrH6VdQNAXN28
27mA1Jy96rBjuVcUscnrSZEy41yc5J1unlbyF5uRCCopw8thLUsXblFwVA84
vrGzDkavxp9U/gCW/TRiedXidTTwNfgTvuVznqWlPgcOS55v8b9Le2iHR334
ivND3pvDIMNP+E6hioGyX3nVmLuReQtvpJhaH4C7cOYuw4TVeU+yIVbg8qDe
IPM/ZJxdxBHgsdYfYgcngKw/A06lpJlQkfwEUUGwOgiI2qv67SJGLzFUKgAS
Uk57TkxJbjnbC4WWHmLSirE2QmAee1FzwRSUzypMa0tc5HfsQ/7d30W5svUa
r/PJk49DSUzDIp7SFVpe5Hjb1nzpRcObTuTT6CUR9O57fruoUcrw9M8eXE52
kOrwmwGXwU0QOI4hjgw2dgMHROJN/FR8QAdwlRWDti7d6FN7pWQrRGPeO2+A
P3q+RpUQjKRpCU14G518qpAXHEN9lEk4exUC4gxXBBwtrWWMr5RAFFR94gIr
J8BeQlZdiZF3/o/3h/DOLyk/th2UVvzJLdc+fz1Zuzch2Iwx96Lo6BLlA3HE
usrN+Wg+F98GaAjGklYRrstfWdzOU0+yCz3xfwuHK5iGZFdVoAyFmBz4EkP2
ZGTO4YV5//+fe3adkcTBZJlcJZe6iK306T8A6Xwh2sTyOrwB3FzSVDqXiXkW
5pdGtqI8Qx9Q+fj3nA3+0RBHYSvwiExC2iIxkdX8aykoCUeFmcqM9Rhp48cf
WgTNwsDs5YxTnYWdOb24axp6Z8nKP7zPbrGAINZhHdaOC1YYsyIpDqW0SQQ/
iZZmOojg9nPrFmymSYicA0SLN56+raKRIJpusyggO6U9M3IlrKQBH98y2fdL
Em68++xpZ6EKlRKc+rFLYMx03lYA5YQkqC/ACTM5gNBbMbPlEV+VV1pj4xoQ
HBl1vYphpTlxsQcFk948Uq6UqP1gSZVEEy084w4Q3x9kIDP2ePHpxOy06nMI
BMpX1396t1peHVN25d3PqoII7yPErRJRSuivVKfW3P6lYWHkGXmApPgVgN50
CigYZBf0Ws0G+shc3p/OPRXapwbHFiKm+alBBH0A/a/a8hLocNvqwTpR/H8M
lUzgcj1M+yIiyynRghtI1IxIst2NdW6D0wCsFlU7IFYJ8GMGmItSQZrdkeUz
kI0RxG94/WEEs3W4319NOqwqn4/TC/6LFkrVK3SgRqXvJoXR5+z9E1xS6zxv
lmj7GcbM0MO+ftviY9lmX/fRHGdD4S2Fs0PYX6LzmqcnUN7WiRhk9DEQpAEa
xWbge+yuyyNhQkXexGoNc2h4JNAflPabtQ6kQ5cmoAiIPXAAGln+LEjaf+ju
S/kb2sdQMChi+KdCEV/eCSGnaeXkw1q488TiJ/uD2Mt0UUF6NXcymgiHWqad
pWzNQhNwiJ6Hb314KLm+0nX8cJhhqT4bboC8qE9Xp6N2YFsTC6iiN7lw4dis
+ruVL659NenxsB2aOwr1vwzXiS/ruTVI1Ci4KHfimraPajKXyit4Ulyx6/AB
0BYyClDpZlhaT5IcQhykgzCaYn7a46LuHisuPO0BYe4PPJVGDYwMtpbGxDJN
oXLmy6TD2jrENGUWx1XASoJrfFrvfRKXLRJl9+uNGzsBN8+4mfGBCZXqpSMZ
Az/d48H7A9zfu/lW2+fDkMLzmWCw+9zHa241uE55BczTRMG8Loa1GL7aC2Zf
htPZ3DE9idGgVDurn8mNXpj8uGnnlszeCT6nGKz/kw10KW+TbSRUP9//ZXkC
mOYzt0xlin2g7EfIQRcUK71u/QphW8kb0IgCNoTk+BEzU9ZCT4Qi92J3JSxG
6XpyqKEMbX3e9AKcDCLltUtHxTEhNrpn+ebSGuahafKR3zcvkQIo1lOO9+oo
A8Fyn13gE0NDSJFCeq6g7na2N2dCtPxKSR+uQDD8gaCQUf7ATf4CMhh/4Qdi
6RXfddDONRsdp8wivWnFt4sjh5vQ8Ec0lnx7QphoXD+Xqif/aLKJCrO8R0+b
tdDvv9/IdVfcV5NnhwHGB6Ji2X/LQd/xtK+qRkNhAV2DqMBzjKbsk4VN04SU
fk0mP1x2eryVph6aTazBnbXyIr3w01SWO2egUhQ6U/ZfWmTjUjfLcbJy9L0T
d4Jjl1QXyd6jZS0vu1RxlYu/wucG/zZJmG4YF9nt4bE0wGck8B1EFgyAIG5f
IklMP9uXsko7Nu7nP/ybhn/EV9lCw4cZq2IIkQtQoY6dsGUH5UJR9NUAkoMN
pzeEMzaIbrK6r4QjDcxvq2FM8aRp82GjWkaYb0On/chj10waoEmgvQcJtjRl
vYAhFdzo51iQ4ugh4cDjPuoqBL3p6OqsB0sz4EiOwwA/MHgKyfFshqw67tY/
9LnuCW36dLn7NudxXa5v0iBdliJK256GepNehWldpsyt4ThJTKQ1lgNX+1Pa
r+UhF4hJLUOtC/L2QK77Dj0BGTKWZnmqOBgUC2qQcI0hzxyJjfb+VGhnCCHU
PGR6GqyyTJndwQsw6/LPY8nG5Sgh+we1vKgKbeYHr9Dyi92o2+hmq5iwf60b
HKepeip18krehJIIK9IDPXumqemiWAasp5FKJpY8oTJxI4YbQrBES9aRJpUq
WFfEPv5ML++F3ziqFewfYgV+bVB2TQFjVQfGK/tr42kWu8FHziCD6CrnezfM
/jipKnLEkuKzM3Lx//eCCupuQP91gUy/drzpwHqqGDluSaaSTV4mY1zQ6KzV
OvjfYQaIfC8QVfOyfuF1w4QWcTvAYrKl6JSIg5ZarHdcg4sTLvAXmq3k9A2m
aK4LC+p5eZeHjtRQFxe+SInihJ7FRG2Z2aCH2goFaHEIi51xRXNkFmUHnvOp
1cn43WxNAMJiRSeU1K8rCnjZ27F9/74+lg4NG5kdREOe8PAN/g0NlGPCGYZw
5x8OEvfmKIb4kDxMe2plxIVgk+6z71Z/LoKa9y5RQByjPvPy3f2SAEQvxCQ1
Dyc4diljilgiji20duFbuWPL4Z/V9vd2iKUvjwxIXmbABcPXOSHBt9hb4BPf
UliVvaD+vF/ctDUE0r2ImZrjKUwaspFRktSTPK5u+fbLDaLpFLER+eG4ewgo
WTH485KkbjNQWh+lIus9FKToalzPbf4rRU2pds9trtiCRsmjX8bCxdKMU5jQ
52nZs6uUaKGdlp2kRWkHCsQ8a3yR6zgSTCVWGuLR1pJHSVa1QDfqwgXryy9m
foIiY001UAP8JDLxJIYdaLCdQNkj+UQN9Luzh2idNWRv2SjaaHuaPv5eVvrM
tiwGa3n1xRgwg4f43Sc57f0m6jFlHfri+fee56x6fJ6m0YmJ89UAHJJE0Gha
q4P6F4Q6eUAlk7maZQbdTy3miurbjyrmZdA+Ng9B9lc227cALS3EUqo/3AQ0
6sIGXXniTZH9+KIAZvcFq6v6X6b1XZaX+RDyVMoVwWE3Np7PZE25rwTsj1oy
HcjdfbqoWfM90aa2yI+OS6IW5PUd2Wql091SdLQpH26T0+m6Ww/WDk9BQLoZ
eT1q6YPapf5YPksr1OGvo3kgPiImya/6qMImW/UXOC8hRk2VMc6omYT4ZDHR
oxeraWNqGAqPrmy/FNIM/VI0G6Bz5N6IIv8J+FZAYcnupXDpwtnQejFHFL49
6D46g85bey8oOeadxp7i2B2WesZN/m/SlKglE7dZ9yuJB5Xv/jDCFXGBgPF+
NuLwi2Qzifav1nEQpyuH+UGQwapyJ5S2GMa+WdjcfJIUIexI0l1INLbdwA7y
302kQbeoaLwN5kGwoUW+ueL9yZqeap5F4ki8MDU1mUnFyukz2KFGcrnKtarC
ogZ54fxbJ/F5CnVmeaisFsRSLiivCwfDE6RY969cYyiOmq8ptVkDJ3VrJ68v
2lfUjolJUgRWnjThf+ZqEIwIqcu1F1H1fv4rpW2jnCdBMNjOaqN4k1fFolKv
6Zb+2d3MvQLkpkLnkorJqvSbZUtTqFft/KHlSHSGF2dVXKkk1Dn1hYFL95L0
Y0lki6/2swN2vY7dJtLFj2pRccv1jyz6H67LO2YjiKow/gMBV8VCZygRJ39/
i0HpomUhutT7cTXyq1HxvgBRxywGLctoMw1l0WDDHWfUHh4Ls43iKn7KuFSW
KdyTJ/QU/U9PJVZNbdrQGh9772yRYgTk2zVaGvfYgALor3bm79xNWF4ohmb8
IXUJmkUFA7m8E5BFYpQKqc+woA2+SVtvaz+4FAOJVt3gg/8iUhDVs9gwPpwj
C57SEsjyN82bvR7PZnQ+BzAZPA2SedSMF5hdn37gNf/cINwIdxAK5Jk0X3BD
G+yh7+EFHte2F4PzM8HKd4/WH5XBUpTk3n7G5vE/oqO1IdunJtU4TnOyxudw
1Phs1jF+hyn6U2LidpAEnp03sEa5LPH659K9kZb9IhZopWRo4QoQg6hLwZRt
LM69zCqrFmxXRC8k5NGYsrdYskbp6hRe010Ob+oWr1nFqma3gHVXwQN2VsQJ
nzoha+2lxx0d05PeNb+KWahGG340tdeJMriZZTW3PhcIHmOLwkm8ms9eEvlF
SeMZdKXp9JukqtrBPQ7d8o8E2MjVZ4usrrK8Ugh2HX5EVOQTmKjTPZxEnqau
QQssigwg0k93ZoYrjl5EHo1C+rTudTURXGEkwChi9HYmR94a99urDdLTWhWF
yPaAO2juk9WxB67+RTopsAIiVvY/LOk0V2JMH1FsASK3KZBNn2c0rnaTPJFn
vHp8w4Ho3gthm2ZxAYynYMqqGjpAtVG0wkCGcMi5o8y/nIAf8OF69iwbgH+7
nyLWphw8GKcAoyD9wSRAdNcVy1H8GNnkw+E8gcXH16cxf0unHtYxaqtl+BEB
vqsDzmddougCoxS4gVUTVX1KTQHfhksM0D6hV4IlHrjc9N9PQGWjPU5npxjO
K7ItFohPq13rkZyDlw0bPoxQmf5j2EwfnMdVE2sQnrzZIuOVaah8ZqRvODN2
g3DcQIqear0xgHZMBKJ/SmkbASlJIf/SLcCqih+d0Xx1vBfXAckDdVhpzTJF
TYRjORKHWEUw2ceoGw+qcR2C8M0U6e/vEZ/G/siZsdicw+xxBJIePJHxQgEN
coX4UQi2laZbAQ4CEJHSy8eJIz4QmoNj/2dx/ZzmhaV2EgL1A8uYU9+rD/hf
VqigPnP6FxbjerdCCOeLDLRSnVokgxfgN3EljmIhp5XwxCwNQ5d7JUcR/XRq
CZCfqdpVe8N+mvRecdiMM77edWpqEbpf4BoXpVrnslcVxJdfodGDBeTddgOP
8AZm4nJja6c8dy/kJV/Vd2L7t48UiPxXaMuwVCmaf2ez0XSG8wKWcvQxZYqH
Q9FpuNfsHS19MlMEUdyv/JCWitXOWtNIAqnK7GcGC3Hj+M5T9iSpXJBNQ9XD
KgByWtnLxfF/uoxm/47NHsIdn2js47Qm3ypFcsy34KY/HQjKQ2/Sf7Z1ZpVf
SbPa5rko718OfchjiV15MIWvt/5LrK34FfMAC1uNKI7qs82nGlXRjYhj4alP
4djjwlzO5E7aLg9cdA2dPEq7TcmA2xa1DFVElmdL2Xbyqa5Jncn3sW+gEWRv
Kb6J53SGz70l03Cjyb+o5tV0/zcn8rt5pvrSk77BJFZZWpjAzKpkzWT8BL7v
2yHe/jeiFQvRV6b8GZ5I7D6UxWykdKZO204XpF0t4ymXMhF8LVxpphFpKZ8s
XM+sJJ+7G7sBroya7DoeCu2lkPeWrUbTw8nPKUSQbvy9BFQjRTck5U21u6p3
vZyUAuh8Wx4+cPAmwEbUXzMeTZJ4gsHxLK+uFvUYpjq/EoZvYL5UCX55y02N
oyp2HqQXMLGgRuPiR0dvbbEVlOstiZ1hcVNw3UDx/v8WHk2A6bjQgOhSJg48
717LIu96UDsA9vl5nJD4CFhEMEmtWdAyEdgtwYRGwpVwtN016crE9E6KeIbi
u+CAmx6LfHSB/tRYNwEwDgQrufJ0+dy7OfOmq+3GZPcF0AOEjaHSGT0mJIQx
pfKdadaqTqDnmw6giBHkqdCTlvdSDs1ToS5WHFmQmERuqIknu6B9RDiDs99G
M/RQNcWEuTwRCpvi8Om5+vK7I+IEAc0kpSBy1RKO3aTpjLsBO+FE0wQmvY0Q
zcEhl54hmD7u4tvIAs0kbw+tWhv2FfHxzIZ7T5GeJ3km5KZbA8e/p9Uwpn2b
s7ME4n/tZBWb5bdVWAr5K99ax6CfERvtq7eRkt5AOrSGf95rppEOVexVJ+32
He7aCyYoStSuHB9TGjhNZKiFW1DYv2TS8F9GXKAyIeUzr15P5BOXwBZtIR/L
4PrYm/hBDJrZvHUt84BdXHBGPS5fvQMdt0dMWE1QtNlFKHuZbfIIcMBupJSr
2IYVecve8w701H/lZh7qDEHqJiZztqT7ccesj6vMV5DPuh/rKTE0llZcyoIj
38OglYAoJVNOUlxg5KYYnwSjDJUNuu/B7m94hZwFDy1qn7tQ6rCd6TLGpj/R
Rt4K1kzt3369Q52NFN2IT2Q6lN78mcBWZkn9wYf+27uJcY2rK4l6wOjLYd1W
6FrmR7i6Nnh4y8qGTf1hOdSJM8Ybjwc6wMW+yxswcZs7RXpuvoNzMmKrKOFY
Rj9ExOYkoxiSd/7jZb2tlpwb/mFiClsazE4m5h9GUw0uJs+dy+VhSKQwMQ/t
VnMoWewcMsmmDBLPI8UgNUKAiuhoRSeHBXEcUATxLJhRD3J1I4NmktUKDOBa
2uQV3mkvWCAwQvuci8yCE7p5aiyIvxX+fG4GHaK7X/9HiygxB1h8zLjmhZOw
P9Q62WEmkGsbD730a9oy6LuRooXmPPSd+ryxIE2I8frwtshiFmqqWy2NKAp0
9oS8useA7iYLmVlRpFr6wlrKFkKWIlD9p9V1yNZbySFtmNmFoWQfMy50tFnh
5WDTsXQgJCp+Wg7u5ZAonrl25BuuNAfgEMpn0NWa+4EUrXcB+qCTyLfTQzjc
q96c2RsJ/3QLhlMbeBJVv9NbUhg7iExnRYOpeiUOraIWr6jFnMUx9/BpiUkJ
XwIuhPIS/YQLcJm1cIwnHhzKETMRWqEwJWXD0BRl+KGngaevT5AU+JV7ljlq
22iiJkApnDYimJ1jnI1apPlPABCGmpxgSvxhgehzWFav085Ypsw/by0G+x1q
IhXqkkDKsoStAXT8JCQvIyUDprXqzHp7fLr2FXd0GbgNvxnhzFZFSFj8NzIg
EGcx3FLfmf3qcejLryqLAdiSAWqPFPAa7PkaTr+VZU1BSNcwkDukOBFCi51w
goLIRvKtWnQrL2W8kD+TWw9yQiGVdZ402RZ3k9UP9WOea+/WbZISYqdj56Nv
Axkqm7r68aG1P+3ckZpPEf7i5YadCzg1KOQPoKvZadP8xVJtFkFmZRzfmmqX
MGBoPp+F+EyIBoPICA+foJgk8Mv8cDDNEP3CT5WWJBvKHuLj1bZtqaULYrfz
Ofj5yAyaKCVZa4/lDwRJ8dWyobFgCIvKMmtTkMdJUc8wU6POX11fLQvbDMaU
RNokOjipwnhpZJExNeyQhLH7HHBhmaKXWke/NjbPRcsLtW1/3+yba7zK1iHw
CQiii1quQ+AIi+Fd/IzhVWbH/CyyPJ3JWc4Nu/txNt8U0sZKE+l3IYC3laVL
aF7nwGaqA6xntO2/8LVDldauMQtgspmmHARry53F8Or7MnsEruZxAVpVxrzW
YLMDCu9W0q4Gea4FzUvTKttim4/ld01jUjjL+KdOUBSW6/YFM3E0N+dcPd8O
dcgZHdxj0m+BKQAytFV7WHZuvycPrQe3R3XT4nmNhl6BCtBEu//O5mE0aZt1
0WU4cxwjKVEbDG7ronEVkEfMO8K7+65tF+6Hs9tPmNH4mX+9PCZRf73rpdoE
AoIXAR3yFpcuoQ6HAgCkgLIhmDRhG3NCJ7IpIWRLlJDI9ymw+orrWIIE1iO5
x50V25v1PI/YCiJ9F65JRy01DjoZyFkA+UxwadWMCZqeEUzIyytdJWhanOq7
M617+MFW1MNQl+94Y72/D2HS+IixCjoGMKAl6dt2dnxS13Yzcyx9z1alQzZn
ydJB/HjioViObGboHBJTlceM7WyspMXWSMn8KMKFPsRZakEOztLIwf46X3D1
oReOlbTKseZ3Fdiv/UGzuePOO7XKm2vCCkXKFrDgCkra6VdmD+BmOn8fDPb2
baYPaYo7Ag6xs0a0lBy6TnGLnH0S8opG5uMOmpiwswCPYNtAlT/iEkZpP9+c
NKc61Z8CRZiLjEUbmJ2VnVQfL9cyfTr8LwHBDcs42j8Fnls9lUsh9HTqWiGi
W2U5DEmj+er/vL6h9+yL/q9Pmg3oV4VqtEKNXsZHBkBmorkaeoO0dkoqtEyG
7Pwq+acppygbpJe0gHAyW0p1UvyruTftb/W0QnI9tnyCLIFiO4oSb7UYaAP8
K9dRXUDVc5CisZN4XhLNesayhandO9V+ZTrCSLWp7MHKCmkObbYqRBr57pIG
aWwpsKw9D5waXXsm2aYOJ2IuJBJF3xAXOH3nhoywJYApH4LRa+WJCB7o6qeJ
6iQLsULVSfSWpcmIUkKWsge77IDyj/cmncgAJxoKSyaAPDZHHisTHuby7lkL
H9QMf/WcxQuOYADQwyjaSwM1od1KITlmDdoGWqOdFHS2ACB27AShekDuOu08
OiD+O8O/c9ya8SuywbKONg4NRPZVC4C/MH24IKV6rvpiIr/FomkxbWxfskqz
unNI3GgrF3PDdAGRPzbySD09qe4rL3rUoOO13p/7+YjruSJ0a5MLTYcCgf4b
wKowa68ZlsPvHf9lEqkP1V++3E86mcOWspvgUfmGpLDxO1RSB/P/OfSr9Luk
QoEDjZeCgUa7Xheqph/stb38vm/C6V4ycjSyUqd0QzqW9LwfU0o3NpJIYFI/
YN9NYcoL2YpaJJgOD62MxoeRIEXyYYIKwEA5OwJ8uWd3v7DYEhkZ0dCg35Ua
MvB58vkq/2FSaaFwG1Uo03NMePGdB/zDcFqeMrAX+aFnc7av6INNNuSA3Nsa
c/wIbQMGBOerD528TlgP91GFrcEBZ2Beknb4FH6g0h9KBN0s+JIU61TTo0Zc
eOAmnG7xtdltYWAhgoLrMsDWWIXZoZNiENJ2XDqhZj5KYrpedRxNy4A9XTV9
QXTsmHRI1U7CsuDLuZiXntH3iPEWy15Ii/V+KV7ZjobJfRuLaDlwieYFwNSg
GK3T0jlEDpV+tQuSOmeUCf3ZrxRtlIjIgs72agvACQ8q1BitPsdcrYVXT+kV
yGiksToc1JY6ImmS+VakBngatr6cz+gdwr1SksxbM1CI8/wtRwOkMfcKgPEu
KExsCGEM3OsdEsUxFTQVm63FjZMBKOtX4vYzRao1uaE/tC+tmzL7L5y72QG4
OBcMfCib1lZTQh7zrdFtDRuS/rf0thlUo+0FUOM6yjrutyoKeN6Akt0Of78R
2z7wkO/QofAoyEWJzD4+ats9eNriRMuyBLw465rvlaM6qhy+rz/d6EM7F+o0
UKV9ocv+GedlseI5t6Wsyizzp2vS0JblffnJT0nWvEC21hI8mc5E6x3tJrUL
lKADWQTZr4fFOSqvO0h61siIR8XXntQIVHzaIV6nALHJ75IO5bdHCtI86VKa
upgoljERR8d6oSOJp8cJZLaFVVQ64oP85RnKczS/cj3+Pu9faBrj8kkxONNU
/wIGQcg28gFCrn2GOMq4dEHixJ6HAFrLKAder/oXDXXizKNJE25FVx3/bLhR
jHrQr+Cmp1+ZUt1vkc8hQZvsqcJZYPn5e8cgbm+VXo4cnAme/lvjyaogZ5qh
N7o/F6yxPqwyuktpA/vQPRs1OwjNDOWQ5JA/aw64MrLMhLxpR9V6/5pqD5T0
o7z/Ry5rX2omcsLnndT60bP12rYr+oYS4O46cPxfxEyqcVOlS9AVLPyoHdCG
7LpagwZyYieI0p65KOCJoYBL9dlZODPNgfNRE4NwPUa3HLCElAeyg0kU3L0R
zXMCL0C0Ij1K6BqTpQDKn5VfeRWD4A/6OGBVkOmMFBlu2vxiWqxVDA/AIdej
x0SSTsw4U6wiqiaNTbUfaiDM2x/YTv7AbIsSKvafde3xc8RiF9WxE/6vE10r
ngg2vKeHSsEqhvPGVYND0p7tgP6pykPjmmoxVMlanplBCflmdqey3ZgfoOOc
Vt+N3lpMK2+MIrhJlyazAqee9myZ3qiepTEzlwbitiD2458yyjLzgNWYW5qG
gv95ARHP858/PUqGjxTMM2ICECUAqFs0OLeUQgR7TmvcdWroUu1i7DKUmTpT
QN5w7lPgAld64y+ou/yn1kRIPGBT3+1JkGBIE2zWF/SgGziyCGkcq1hr6VQ+
Mmxh1LQS0MicgQpTA5oizBeEVzPZ+nvqxEIGtr92b94wGYsFnby6XSDEfdGQ
EeXh6L0s8vVF8Ch/e6XBxIWbORqLcmdiAfnZbnKDdDiz3zymiLPDC+F3kH1e
2RDt/1fIJXZ5TD0zPSHwG5eHq5q9nGhDSNWyw+nfm2TnsHfAO8MxiJpLrwsq
Z92tu9DkX/ZKZoyX9kFV22+/CA9M30O9cGDZu4IpwAosPYDGzHcW3J9uf0Ax
5wZ2F6VJVPwbhMclZ6/6aLlhgEJaYwh5kaMSQRDlbQV2H0oO4wu6XuyKg0uF
fBtdb6wLH2CcTEKXxqpoxFUJ7i8HT3wYby3OvssBOyqO2vgxgGXq11IRAov2
2ZOqVJSg+BcrERAAVGN8Fj/WKRJimQbInMRdMVurGx/2E4qp+EAViDxGttoX
kmLlDqeBakemZEhNrSUyk7LhwwZPJ9fAXnuChsnke2nuFeB82wzvcfiYG1+W
AJCaYagzq/tXeE+Fo4FBqvOf7M0BRzltonKLKny6V2T7pohbMULBgsQCF6oZ
z70h5Bje5K+MR70vNDE9j4g2vOG4kibh411RWIdQq37ari5wtxALbnNjyzDb
xPTKK/pOXVczSGNCBYVy9tdr0kqE8bfOwcTd8FaBZXY2obnrobcP0q3U0//B
hGzkH8wlkf+p6zrpZxAnzGjiTejADX8zW29QnvpgVuaGTSvVlJimfLS6Uf+U
+FdjxKD8LW7+IPYZJZEPgh4aGRkYiHpqbeF72TV5cQZBEYEqpMDHQjtxSPY8
9P08XIg4l+zXilyVrK0Eqiwbbl5jfIeBFLiad9O81BuBV4DK8me4pIFUbjH7
82ITjzzYC0uPy3VnFpB4145fNM0jd1vG2FjgjT/pcnpYHerUcpU36zNiyU7j
pUlYnrHsl2t4aQ42PEMj2cCS+0gDi6yw8suQReBZRIJoh/UFeTU/tMz/9sIT
NUIDyElUUrrN3ted/G8esB1HdrCz2k2B8EQRuagjYgkLWpwV7HXfr2k38a5l
+e9EZA81HBIeX9SaEzDr6dhPOD44Na8Cj4sKfI93a1ukrJ708v2q0288rZj4
VHtUdB9Ywuex4VC+Y0htzT5skqHD3rS5bV+7yt1DX3B5qvvcwdy0nqlI7J5x
WHfx1cP25E1dhzWIN4G1DZaQXMXsgaEqXCQIu2QWLxsUAlnO7zF20GpYylgd
lfKIZC6hhk1f2L5L3C8wXDJejNmA+8CJcrR362f1SOW7gsf24pxc2+BhNaSW
WBYZf8LxfbgAfOt6KxSRs6CJ8kOLwItpBcFCRdPjRXrISlldlzmSitREBw5U
6092dLqbnopFCgQJgZb62aGBcmY9mlYNBPsvUgl0l3EjYe58R8romx0ayQjq
AfbZBUWDf0wtx7+Iyw5Ha4beQERQ27mITGC1Fpz+SEbp3n18zUZe++nCNSYe
Ud/rYyYbYOLiur1TArF9Dxmfk25qFZ/RjFYOwBA/ysHuX6TPXag+Hb1sow2t
2RAaj8/Rq2sed0IaeKRjq34WlN755SkkOjfjdiS9R48103Ff2IVRBn4xrgMU
I+Bl6weS88NkMmyRt7+AEk3KoK67MIxx0CpbQ10fY9jdQJsMbTJy3YJsDk9c
Xytch3yTvXbRovvBbL98VjyRBFW2uwYe0hongu03KGiRC2eBYhVPVZa2MTwo
MNlLEa+HETB81Zm2/cmAOSmIhsYEoKCWvD4xem6Ha9FwbgtCmDUSjeNP53Ps
ulW2pvcZaTac+IWvrNBDA7w31fIEkySEFA/6ZZnfMyDaYSAshNxmHWYjVCht
9VfLZ6B9BLSI4lHIYTudCQPfZsNFBjyqHvrHCvP/RZUaOAwLfpaDd71lOA++
mo+gNQm5pmA15WLiueh6nAluAODQk/9ESsiOIxI8mw6VNCA6KaZRocAwGj76
1iBnXYEcNkwElL2DHDhT6GZOMTRgd9r8Y2W86q91uMcvcysyG4p/3wDJHhcu
sL1oHLOJpcQlwPUCW3F5xTDQN3NqHAbQSTgajQHS6ffE6S8Gor75za08lEmQ
5Mhf+PN9dLVjNyGjSih9zPQG/aobuXgdURKqKaYCLKY0PihOHSEpbG0QbPbo
M81eSMco5T0YGt3yIh6uiSYvtckDUkv8YAzpHEag07ePeT6KFa3FsFfRzAgQ
ghMWlq/MDzWOWGqiQ9+bVssQxOQY6iRSAJFZtFWSPQsT5ff0YppPgOhA+4HS
4hMPjA0wvi/CHqnXibZko2qrG///3SJZGZXeUj0dx47zcn/W3n8MQR/BDx8p
hI7txyjFqAu0rVVvbVrDiAeHACGcIgXLyLprZg6aSXMw24kPTbyy2QhdQlm5
ZGgWEUg14ib34udIcwTNdzctOytm1HJbVl1JyJf9kx2+bQKaXyXgXhBwScBr
CXeeNhzSfeaUOjXneKHbV+DXk3iuyfvL4pSZQnurvrXPJzkTgeFbHyjGi3C7
ARtq6FW8epuGQCGPIMk2+kdJkq51wmkc+s7QjYEL2Dnbcso4ito8U9zVctJX
+Jcf4xlSpq+MF/LZCRtTk34To1fgy1j1aHHmN3wIVKUa4nzjlFH10gKh0f+S
ERsR/0CaALwCSrgpc/pT3ZV2dFQbiyTjD/dC0X4e7Gq6WgykmkZ+mBiPlhz1
dsVVbhoMnauLtRus7OHFUsp+8FgqB1BCwrepwMEa5lHX9A/84/6xIbWYjFur
y6Gy5Q0O8MC6iwRaaP/YsnlFyx40+YAh2A9j1uXYRSMvSggHZZFqluTBDuwh
5UQrqepi182+jw2dInQyiKL+CUwWWxpK0rUY5/YEK+jK2C2JxUV3DjPl4Vw/
i7jHL5k97OWpjWA/PwVQ9QoQcAKJ6TIqXuzcTEwjIbeu3AStoM8GjVtvviw9
ErwxsQB28px3LzNAFeTV1ACe6aeNgWVB++IpFcAcJB7qVxmfi6YxT0BisUJG
q1e6YNlpiFQtKNjYu1yLshsi/j8Pz548iFozgXQ5gfvCW+kRI52d4UR2Vo5u
yq5/g53dwOt/e6HOWwXCKrDpRf0AYWl9j7x9u62+ywOrZYga0E7U1FGVjC1z
xOWomJGlogSKSlCYY7ZEgF7b0au7yXSG3m1OMZpQHVF+sD9NhumQWrB648Z+
GHRQmz3o8b8UNYwDQq6XDX9xzOmjWronRid8fy7841Md7fF7EB4iCB3PDrFX
s87AOnYYC2Bq+uOjEH5932G/Ut/knky5rAvKv2UVWOkEyH2/bTfQ5htCC9CK
xuIHTnoqqz4F/7D/frIG77j8fVj2Rs9XPIQKtKJktlUONh14t9MOwcrOl72H
LfjB1T44RmQAXH14bTQ3TFMbAnp8diezCjrfWsl3DQLVKLrDTclGJn2ovATd
eMN4OJQnUzT571+r0MnplS9BztndwekteBQ2MzAxhstBRo9ipWwCfnHC3vQw
XEY3BxL5zedTZKhlHeQLaLAFoDZ2eUHq4IIzi2z5Nm2T1bT8zdF9nKoQthvF
+CYIYeryM/XXdEhDnRKufZuI916HMkiIpmY6U5BRvtuCutUfr39sX0TdUtU0
QcjVEUvB0mUpAstzfrtCzmWIY2jLpu6i1/Z+GQvYvByvPvtR3bXbf1lGtaZf
HwzjYLzziN6HMie2QUxoJBzynopa7GMKFTpHtthqmFFjHrIE8KpzSFwbgN9M
EGD5IqTB5yMa2pL+prpCSF2AdYhF5IESkNpJ2UdSJE/VTBd5ejcn0QwS4dFv
9hlWC8h2ZJ5qFvrsA9kgc1XyB9uqLCaweURK2KjC4xAal/pcT3y+Ko5ywQ9n
nHxKN/Db+9mRqCfPYAznkRDPjmRaH6kWvur0pGQ66fUkpLaykXkZ4BqqA1oq
1gJWDaZrD96FKNxfk4vhxmRlw7nfATt/VSym10AZSL3T366YQTOcKUVrpGYI
yx+3ovW5L8aesYN5enwfdQiO9rDZHs6zk2a1iRvGV3GSMGAqcxgHyjW+yacf
+w8tdqbs0R5TodmiDoEgRaBOXMd6HDhDx/I86tjCywA2EXcDmfz5reugixHX
uXrPISoqOON2zJ/5rfewvk0KyqXUeMF2QQM1OCDEe40g0sehyEGgvoFsb/C1
+r9tZ+iW8DQiN1+vwPKUKnMFQxpRWrHU6gMR1ORODpOAPMswB/KgV366bqvi
mtnSJHC6hZQcRFGcn9s32xiY56LrDCzNJmGjTKQEFnL0X7ho0YZHqgfFHceB
R5Cym/2PP2IuDrq8+d9s8LFglvV3Ua0MiMT1W0rS+s62NmAFdCSMvvY+TlNx
Gl2SoWwDOQAw0qM4XghAyxWTiNptsrju5KIAU4fSMoH5cb3QSqDna1bM3nl/
sUSLPTByOtpcAemzt/94kNgAl4e14cbkJpBgmkffQQxLPKO1qNlN691pkAi3
ttHRo4sWUBt2rfue6Ylr7KlxThI58lblhpFrcItytiQ7ESbh0ImVUL23CBBP
Qljum3R5FYS4NRjO35Q1JUyouVmaVOdQQCPC2fA/tP4zcNi9dAmrL643+VIs
MByJ4l0JLMgZy8QsE91P4shJHt1jVFLzkr3xcsr1t1caJc0vsUHzvSUe1oE/
ISqfYQ5htwqSkpF1lW7lhbJfeG/jQ4zcludCcYZF317wOR+Vl02JUMCJu6SO
z1FNeUQhq/PJhQmBiVpfPjed7aMuBo3Qs1vWXoCm7L6lvvuKnyYyXwaPCX/t
k36uHDRIS30xgA2pW0mkByJuP/Jarr5loE2OEsY2Ih1hE6ipIQD6zHiIZcHl
3oPsMSms9UuYOVLTxTl51HGtBrSN62l6t9WqiErNuZhe64qZUR4AFK9kPldD
Nm88kvlzNStAF3kzqDoI69nY+jawOcKbTAABGMcE8o8LDPxv49IbtdjBQCrx
6njtEL/2iAJOz7x5kggml8r8CKISWusn6g1k/mv0Qtx/hDy+TGIFC7ey7t+N
0jPHN8dDnmoIx2o+AIXwnbUsfjml/hZyX8DziQdt+nETT8nBGpym2qKKo7tJ
rvmVYyb6kufyHUAhrjslTHcILKWaYwzkVOsrIq9KWT0q85i78JKsqLTl2msg
vnFL6YaQjZw7V4q689T06kl+Mf+UnKhNiV+vSuBeN5g1KpUUFixHx678pnRW
a+4fEoT8QswUPg4T3juziBgmMHwXkJZQggJPPXwcRYrbcH4MX4wvqN+EjoIL
2TXeeVOAZRRdiUikLEY/4p357LmAoMRzFyHU90M+p0qwNiiQU4pem/GkVfLE
P3kk0ujDDMrtp780nT7pdWeRe3R1EHlZN/VfRPt0tOe1DFQqgrIRuLshwgPr
ifYFDqcEJTmoUfreFfQWZzlqcA3uk4sJz96J9Z3ulrqiqZg6ZWu1LamJgOTK
vW6BEE6X3YClhUK23JM6lFubRkkFAaJ+i8ZX2OOPk3s1w1BCuaN9njJxsCe5
DcI7kejLjTGaJp2pwnYQ5LWaDEm8BTHkRRV+Z8S3po0Qg3QUk8H1xZA5lzK0
avuSk/q4Gan7exeE/PwQGO/KeYaAJVrvA+MFBWEOVXKPjIZ8LctnqGRgZgpv
6rL2HaRKJ/G3EsUFdrCGtIh7JbkAYtusNzwsolo5Knomc8qIVUwBwi3JRv5u
8fiNXs2nDva8Pjs1qSapq02D+A+20QMt6IwIIhIFJhOrsx2ic5J5xiJnj/N4
9lUe2DBWGs4pVEaCvqeIlH87ZYcbM9Y+ArsXoyfJkVfUkr/YqjXbLhf7Zy0x
Nxwx6KFzg1cemVAUT5aosyhZ9oj6Is3MhM0VXUaV+b3ljncLSyclIwxJIb6p
Sqn9A1fAZ4NH2XRMYrYcSHC+i+7u1PxZY5W20c9FxZs2mQjy8rrddU40kR1l
Ac6/dQm1ms4+w/i+Nb/4j3DKpDLLxh0N6pmOuzHK0XCnr70gVnWilPLxoQLE
BumKIorfRGjbbC/d6ufHG2JMtIFzLPUZnOwewBDh6ML8pNdLv/PK/t8oPO97
b+t+GSVaF8C4OqMGphIrwgLhoEThH3VfOGGfyIkV1j3MGe3CrnfuI+kYzBgg
HwnKGo1DRA287zY1NCr59FpJcjaXrV493Wg4fNTZxiVtrCxf8auIXr9YdtUh
22YXouZbJCvAeHZaNCLS4fkQs7NDhRUAYA6uarB3X8V+ifQ+SbRh7H+PQaBW
XujAkKXy3Sv8j4gMzFAZsf5iv5OQfrcAkc0NF5jFUYGDQiSn1eNsluK4PfXt
hRsSzys76L30I0cX3kgqGKu3elR6RyYDy4kWLvN5HLoeAurD2MggppCOEYRh
GwDF3ugIF4QRnDmegXb/iq2yWb+0BnXLXwYLh4ryjUUDLpTMpRd2fZbZWZ5H
bFhmDfb5xWprR27SM6IvJOgr6QIcaJHeNHqjeMO9ohSvGK/wqh1f3cOZ1f80
Dus058a4hQgNQBOzA/OsqJuyojp5FLs+SRKUnu5y8307PAV9c2THEEzhft/z
ukjnnMz4iqXhraAGB0OB3PWyve5C4YUcRN5o5UDsHG384ki9mNJjtgjnWDpg
AAv0w7y+8j0gnz9qfngnaHuwzgpQcMZtFiqTPmukLOXp7xHp9dphES8V+ytm
AZeZLFRXGYpWhhmFz0W66u1ZBzHnqIccYXX+Emxorcj7e1we6bKezy5uYAX3
uYdXOjtk9whY8f6CYZEish2BaYVqNcdbAtAtAeA8dj5EhKtjEtswD/rrSClW
ZGiUP2IBqh0rSpFDLsLov65AK8GKyaLlL6udl72dUF9mJBg57j+wlMZ4o0Z3
nv9oXUvT8eECT93gc5gVRpGogkBtDxXziybqu7U3abKtctDctmaBCzrz+2/L
MrIDIqGwgee0rft0A5YLLmvLPGby2GOfKRl5TfyAHNEZFayp/utBXx+9F/jS
+bHCu8+AKP/cfvY0wMcB+yh7meZ8GzivfYDe232OQ5KH7r/mAt5EnmJksRNz
GopJcEyDmEWC2QWxInU9ybdYAFG3a70WiVtumx/D6L7LxLu4MPI2nBOKJdgr
vmyROYjrdTy6JCLvLjHyuY8h50uuFuqSxzYoAYUpnIzrZwb4ZNX0L2/0hmYj
gxEUK4y0AN36+hbj0Uuqzg3u0j9U40geM28CFfjBOxxGcsqoN7lzYW0+lHJx
z2Z9dObe1oIpw02Vdv+VZUpeLrBncrFdB2EC3hWUAeWDgdTERHxDtxWUcJY7
aYo7r/PzkfIlDvqHFqFHgC+keKqYAkwHGxaKkF3SG+PhjZtXDqFgVJIgW2Kq
2L/9WDMcehMQT/8PWb5P84t5KYZEuoB9sVCTmXxIwdwZwekEaJ2Lz4M6d4Nz
PVqqBjuXvGvWz2+4bAU0Nj7gS1kSWZUNDRCDWKHa4HmeXKAnUmC2qgRorA8M
mDjKlC0dxZMXTvLI88uCV2YDDuGu7QFwix0kO8LU3KSn1rHQHvVYc9snyaC9
nwnZu9ytgkgQ+IhTZOy10nC+uV630fNyri2CdEypjQtjyfQD6aAqPQf1FNJR
svcfECVOjqphHyKxbvcCUOUGDC+DpRTA3lr6vUO1jRq4A8jkM2DM0b8gqfMz
SoDgbCMPoDlUxEbbHxSi3tk3u5aacR9cAYV8gZhkWbCXS7t7skN2VzHOUjq3
azhuHZd1TNjdp95V1qsyzQLQ7GOZT4zMDSuWBnNWjd2duE6RC03+jLGCVBGq
NKOCjblwA5MBp20226YKckCxgNd8jXr94PVCSrdyu8bCm3lMov7/0c6FV3/g
eQRJz1fQKyBPnW+FL0fx9UIdZQguTU4kDpDCGA4aLROkMUnV8Zu/SrD3+UQ1
oFXpv78x8bjA8nL7L6asoCXUI1AANDHYsc5H6a2qY9bKdFW2dZJcz2N4jhYc
uZRgDr+4Ozdsmh4playqZnQbYWSifnz3/19LY0QpA4kOBEnEKpZBAR6EXdyb
J8FaJDgfDGJ43oP2COygfhy9b7dEX5Gu0ejcY0rRiNBou863/gkrvzZWfP6K
yofXqTTJm1c29hA+658eA9zfS2JtC22YcooJ+pTul83qNNdd6kh64hKcat0V
vZvW48z+vbV4HVbtaKriC/EMuZUsotP+RjzWJp+eTfnRRT/SHbod0+PLw6WY
/1HP+P0iZ8X+0cM8YuD+Rb+uqXdwWkRqBL9LnxtQARwf22I+xCGbYoqEQQMr
2g9Dz319myYVn0j1RfHpGngZ5lUkBsIif5vN34dNJY6WZ+tei0oY+dyKitq6
8wYSUCmzLSYfyfEoV2ahu9q1lyNSstKU3ORQlQ3Ak4OCnCO3Mt0b4ZrJHC6F
BiRw7l0eTmzBZhTt6gQrZFDncS9WWOiRwu5ayAMjZgw3ogiLeVr/KVC/q8Mo
qiFWD9t5tFXp0vfxA1C+mczkoQ9e1gu9+ZfamcTp68skNxKpjvgOmt0vabjk
rUHMF1FuTT2hmRGjL3GtxJmX2HlGp1vcQRGVB8ULGhhKZfz0WionUf3cCMn0
fJIJ9EHgaoLAXI2qgXHM0m/v22XgaxS3tnWZ0j4hjdrWRbetc+wyUTy+iAJm
6swdBgwNo/JD5pYcyYnaNs0fVigjmh5OO4ukIittVuLXBjS+l+iic7R8YJT4
DKzT73iR1odP0XOw+und/xVVlg1kT+3+FaA5k4ZMpSd6TxQIn1GujMUheigP
Ji0HsKT4zFpWhdfdgWAAVbQOw4QY6Wl2Evn3RFcqyVPlJXLLGoP/HDI0yJe6
feJ574TcIuPcfNOCGjnCSl+zJCxgG++tyJDswuC66JXLGiX82vDTmvyVWq9a
TtF5f9p7fYs2gBCl5DsgiFSExDfkG2GR9eBdi7vB4CBzE7p2lKfLNejOxx6q
RpjEItmC3faLuuBpaNgqwP97cOPPACwvGwzoOZMcYEXfeYQNsL+FdEP9OGHW
Isi27a9PwDx7OzCkdRNOO1d6Iex6ftBKcCVZfPerO0dI7L5c9WkMuZKRjVyp
ORJEG/064gwX6jzkUrp4VRvF8Q2NLUL7TdaDUzmtLVatkq586quB7zq3naDQ
hSPoND7DscSJwMligw5ggxPE24tRpe4eTgdVTqusRtf1M6/w2GdWbGskcRy2
Wej/kDXpSs2+LrHSW1o0ePrjMPzWrmb6RqDXXmHrdMbRFsQtHBuPcHzdsI5t
mOG8e8ACdGtGsHb+LuJ7jFthhFhdyWRFosoGR9jbY2xynO0m4VZtRdXuaIld
Y6Ak9Rucv4dPTAdx0rLZgE89kpbUW5wMJUnpNyv7cLmI0npph6TnoE6Jk3zp
cD7yHp3zxYa/R4fJNDhw0hdf3w13fuM4A2OECkXPLrvNpZONBHN8G1fcnm+i
2ZgrAA9c/UEQKiuFRC4NQyR8SNGiiRd0yxO7e2Zac/0f1Ioy7N5yHDpyZ0K5
3DmJEPtdV7tnyx8t53d2tPACpD1qHfncttq6XHn7g+sU8IXdcj9ayTUrGV/E
v2wa8JAk/iHZfIAh1XRTOx822vKT1v1POICVA9vJiv5+lmBC4Nx0mw9DArpY
a2HQ4lrFJQrKN6Uzskgw6/BfHADdBYSR0QkykkDNNVJ7EdBs3Oq/P5UMdpSP
foawEpZqok6pzYGnjbnpIEgPrDj/X8B4IqQgVjiWwCvDa6ilugD+1Jx7g7S7
V3MkcuPxfwmKZfZkuDqEDgMcwun7MAX9QjQKmUrSkWJkpLKCH/wSD7uMIOYG
TUygCYGR8yxIK3RVtzHExPOqdFISLTztLbbW9W3dlRrawNWAH1YRRAk6kg58
+kJcdvmJU2IXRIQg/ZL7w2mQc8JFJYhkcDrbl8nxqezphhFKOq4563pug6+0
kbiJTWtbkDZKoSDvflT9kY7/1A8kSJDroU4b1R79E4UTb/V1QB0+2g9qc6US
xRoyuLSkG6OSxaLNxabTU8lpM4Z09a28SSZ5MAFE7dCfxW/9ks4LnYLrGGhT
7hLlTIsV1B5fwp2DTvuigkvyYv6a48s04bn9sEM4mDYQeVGqJFgg9z1+MnVS
RKyXJ4Mt6/HET2kr4/onP4CjihEPmubsmFYIWJoIU4KOEBup6CKvDr1ZzpE8
vMVQdItETNchLn6GZWEKefoS3WRoIvqR5CM2ngSXqIYeRtGoiRrdKVoppKi5
knwM1H7TWEjkBixtVjLnQn4e6beXJ50JS1HwdoZPha1ZrGbKz/PGI2XDQwx7
c3N4lHzwk1GU88cYtP3rZIpjpLjJNH56/utEgT+Qo8Bo2aqAa4HSh65sjYgb
mSNlYg7vagVASLBAgH4RM3oLyLr7IaPvarmh01mVwe6ev0CJ9mMeS6UTm4Fc
hWxP/CKU90E4ABYYgXlr+5rg/zq/y5gO7FjRQE9I0muO63exA0R5ecr5Hyt/
aKluQ0YKJ5MWapSqWNRocI3C7qWYGJkrEKvuIKC2ldFaLWozl4NAzVo108ZV
0saDBEkVSsT2mH+oKFQ5sj8dnXJ579m0zivO/934vA5BmuMvo3tbf/KClEpq
FLkcYl0gPPhz189yQIUXsDfZWG4lUU9exhdtcskhOgE3tsS1/0rX3mCMa2UO
MYazThrBgcDH+7i+/+9DTScVfXnzlK2RLu/e96ITGI5gHUQSPmcaMpjq+QLP
cH+Y5CGyUrX5MFcz3P8tDCz/1wjOdHz2u2KDAU3Od1U2LgabIuK1MTXG7KwE
renbCOMk+2go3bRjbV3/h2KJs+abAMGUbs71slxmobigVPNDc/vuoIeOXoMV
I9KT+H/eMvl1yZd1jk1///YybXH7BsiTYsIAHLAxoRXuN7rSinyZ10181lxr
+3BDwRGUcMvKVZJwybGrdZUtjJNfInz3jbzzmNHOTeGSEX+e7rD1/GZb59b4
shVTHXrmwUhAaPyHsIfXx77lHnh9y6NtJD36gb8rq0hnlHBoyfZqFmKAzIok
eiN5GDoQPgNLoEngbaX5yb4GMKEqFw2sPb2tHE3voDwLUDSoQ+0DPGNbcHS3
TbRbqx/Iq+Yfhb9Q8byUgl59WlNzvqraQsHFqoylff3k20JcKqUyfZzRs2qF
ntbJQRs/GdE6HKzZhV1ZpxRqxHW4WHNso6AvFWfSN2SK0f53JV2O5oJDxOk0
InhO1dQnFYUcaFEB11IxjyxFZk9WOvhVqi3ah67E96ag0qjgAI2EQqK4ZWzo
t5VNzLZZ1sF1S8hsTQqVorc2Knf79w1swa7IMo/8g92u+WFrPedz9CPO7WB7
J5h6lFUC/FoTWSA3mzCYQ6hM8WXiNxDPjmOktqT/i3UyBsHUlcPpRhMdgamT
imyMrtSqrIZOqmAJJcTGk8PypDmf/F5sUiLafHO4F5vFJu/mleVai4jPRaVU
U3hQQ01uQj/exPwANEf4xRCeIla1q/tq5h8fRPr1tLWvDdH1DzdDokaunwQc
qFDCEUHal/XF83AKxeTMti+gKA98cPNFILiXS2xuKfFrZNVHORA2GOQK45Ez
0H94DjCV3tiDuyA960ltSElRxdY+d+M1e0MHVEIQY8TG9YQkI68TxRcZDxTd
xwFWNN90/yE4+/Sw4lLsVSM0MLPVwzTM2D53WT+zBHJgc33mKJdhrkDckMty
9CqrP6AKUQ4qK4PkkHuulryc75WWaoH3/asGZURwRyzPYiVyCRsblXarzbOP
VK4Y0zLYiUGZr3e79TeDKg71t80XTC5AmJpUtOzWEhG+hYZS132aIE9axoMq
3SAv82LTWp3+bR4Z5MbvAz9Fwx/pH40cpf5RHHyy6d6sfkKiRYQUJtH0ShOE
bSuHSQ3kP4xcK5hBuHMDqfUl7Kt/n+0BLADBzGgrAFQktS2NBaW3HV7cQkul
U5kyC/x/wNNpUeZKKhuv2CDj3DzvhvPnfjiHiMbsQu66CSm4O3J1CZcqavYk
23JI5TvSrOwrlQce1XQFTxX8pZI6OKVAP47gvghSg/exDHd9gmhTTE/STQKS
ImZmFNdv9EbM6M1Xv2pyzOPVmRce4L+5H3b1MoSMuL2nvsqBY0G7wliNQpXK
qih99vl/T2h1ItJTjgOIwRIdUWRIN+17CtM61yPYzIxhrxgTMOagQeyxajpc
nCpnnOD8oU1MCvmtl8l5bnRUMjqJhHfwE/ywrf71yUkR7TMClYw3IGAYOG2/
sPOSpa751oFOYv7FQS7HB+9HJGKiQrnTWPdPtYjhZTGSdfmbQJMZeiBou4YZ
unPmFkdcbw0QdWkSjSeGRRXBCvyUOsvD0GjcK5p7WexIXXhZDeEaJTfnxnLe
rmI2eea2jXvRHb+V0r4iOgKKvkfSKKVh8Ylprxzyoj/a7jxCyuCveKbLB3uf
yAxLM/pwjBnpEWAM6FHe2QfYKmiLB976OT9QZfp04MrjXDhV2RKuUtaV8fgm
V0iJSGd6Pj6vCxKtWmE1Er05XSETScPZm1r9e09D+xz1BHh9Ue1KOM3+Yhjr
7v42iOqwcOPEd07IYnox4CQvvh/ToBVu2+NCzj2AFk56CPcQC6shVE0L9EzB
sGlfQlsfBDy7sAIBJMWbTKd5+xo12pZjDXjkrn4mT9+QVtSLLosayRio4OEY
bt2SloUGEZKVVLVZazO1Xc+7gy7wKWTBGcBOhYJnUl+2F6z2EnakzjxPH6i3
/UnXt7mxmLPOJpvbUtAOO+0ph1lKu++B2gCkOfRAaaulDTSB9Rjzd+9ZGYTs
rGK9YZhL7uYirYWvG0cu6UShwSiVelCgLNJIU+mQ1VSSX3f0a54sJHmeVQ03
ww1LSNchuGtKDwfSpTjNsuI81rpnJ1pQcofNf6Rya70WoECCvwraoFtIP4HY
rp2JhN2xA50dfEyLRmuEVo4fBMFCvHYAiRF4D244HoTlvKsVJ94f8a0FXiin
Fh39ufGHEbsWxx9nnexi2cEw3l3P4swCPRDKHmMKYmxF+hiDjpUUwj26Zdhz
/jzJLDAzTHFb/6/BZWULKXtGJfn/uwAskcvkMaHyOmL/gkYUpQBsODZahDYd
8wc5TrFtBIxbLAe8GBi32iov+WCCjyUDJr9jAf+1IpWLxD3+lYTSkkw8sxsG
wEQcTV72dIhBODfAsD7OSs5YPRzJ8VYEj9IhOWkA/dsyS2zLWi8mLcK/chKb
Va2rQpcKQy1CxejmXrmv4MYsmflXurH9jViH5qVOKfuejTJeWfnw6+ZX7K4X
rsyTLIWKo8dxXWDQjmLpXCdxAL0uPsj5OK0KpIYZYdH+ubvvSG0PHjRsvP/D
6D7NA7tCjkFF7eYNRcGU5eATgust/gy5/3ElUGyK/Qq902whlUtFQ1yeUZ49
NnlDExkZgg3ko85wUrFab6kM6q5ToZgVSUWGt/5q4pv75z/bziWazCqekDEr
PxeOdnyg5MaiyMvooyzrmeYLd0ygRzOu+rWyxyzRtIfZfcw5RZISBEvk8OvE
H06k6bkcGfXDXWWKYlls5n1SyMtq3fZUHrxBGdzpqt9ffgzXgYR9SiLu/NrP
X+l0gTVMTHQbBF3mqcx/5KWTk83O9bRHt69UHwH0rOKh1qOe6PJ7lgAGSV0H
++YM+iOeBq4SoaCVwDCZQupQv41+gwZpESs5ulHgn2Or0e0V97y2zD+N/3sQ
wc8QSUO2hZW7rRo/LEgPDHlDEuJk8e6pVovUFa32YG9ZQHmuRru9JPmTftSL
+GLOLb+aQZFcOJNYARUjIAkMIBnAJOp299EIMfB4g+se+fJbOHO9RL2OWRXG
Bu9uhoW83w56WwGkIr45us+A9fK80y2H47Vqydm5OFNAiviAwv1PX8gzgArT
fexcKTls4u1V8MYICoJ70QjgGr3HtgWKdFARlNmYMtXN4L90qxFrYnNe4JPU
j3HRj4I1KAgmgeKkUYzBDXYgKEGD5cLSyd3iuTVHctbQIGwAf4a8sC/fKP99
cwuoE41Nt+qnunV7a1PcvIsNnckI1Y2F8NqU5A+a2OJ/mk1KABNuriQ4Im3w
21Ui92AMvpFCtSNAo+FtslkgxM+XehVuWbZkVerl0MNXGE3tkO+N7j5qIY8K
I5kBnyjEszfOE0L9T69xkx7YR1DRndnsrR/aUqkoB4rdg+FQGY1qTBI3K7ll
tk4VgtycEkyy/WF+vTUa0pB7qO09NGT3sw0wzjLrRjaKMFF0xeqfF8zN8oXD
UH7YxRYfXn6JZyB5UWaBRwu2A0Mz1gP8E0GXagvBJH2oSPpza3SoxJasbHBG
C2aQR7G8mNGbKNdjhxPjMI/mxt2/sVavkIS3QqVZsXiuhx2s6yqkybwqAe0l
6w33JG24UcEAjBd2ouPbcSlAoCVpHLKAvI7ZKQdIHmuNKT+NRnlk08o7JevY
3vPLydViHvWpcAcqXd349dMLDX9SCk6Sjsx7oe5HX8/hTcVga/WjpQlP97OM
/lGmPGbST9iQFYRq7jzoVBAe8Fp9WL9vJNXWMs1EQtYHFvqtIe56Q3ukVAN1
9C24rjKPsh9j0F79ZEbsWKNQz+bE/uv84XcNyaayL6dKTAfOt3zLR6nAYTNA
Cu1nUsaIAxnrcLi0E+rfS87O+1kuImub4uHzdeqQ6YM5qYQINDkSg27T2YaN
kEXFmuDkb42Ec3fYpUvD1tDJK4RlVIXOntGY22KKETq48PofbaTYynAGnMBi
PYbFSVCWDks7JAL7ouJQ3ARFurDnacemM9OrczdAqjobHbhORCdrDg/CoVU2
QvYhRXEEZB9ywk3gxcVKjlgZe3/lr+r75hxhx280X7EZM+mLkVeAsJNFtrok
gedGeNZQj3QF0/BN0AumV9FysMvgWCMYimlKbL9lFbM81MiBha22IfiQ0SlO
Nha+mRujdB89ma32vDyYOTzVk0nxEEwx6mhkUsBzuUIi+uV4ai7N6i9JRM6T
9mC+L8ek/CzXgiusb18Ihh1p08KevTDiYiZthP61gL9b+2VmDYjgqSXRknI4
RYbOkH9C9CgJqy+T9lPtL9pqYVIXY5U+J+WX1wK5KpIDMg/gserKhbuORn5x
7Mjkb/kkX7Ico25lKQo290amhaEB+vvQqgMdqZAVGq16JTg4NipNPjr1qRwB
FqbZ4FvCSGPHdNbGmu7mVed/wKEMIU0UIUao3z4oOY6iUUFm+M4hFOqsWJdm
MF1G/Zd7PXBUEue/ToNE2Kr38y0PERaWhkjq1LvyU4t3Lhc9t/vShvYWhvGJ
MOWfvOr3/wqMOnESyVNadOTD3PgrGR6pvfw9qX+7tNNbQzbsk9dQ4FTKm93R
IpWlPvkuRKyjYrxymmiZZTBVhzBDImJfKR6/ldusHRsgbrT/vU90kEDtPKuZ
XGmknQfjejmRwBFvv0SufuSducbZkYloxnuUtXOrMQEOZ8CgTRUqpGENxaQK
dyLoCb08zH6b4Ql35zpLz1pFc0fn6E++agEE7hvNWDhemVGSAuIirPSCvT38
eeKN5NEYWopLuMUciwoU4n0PLfPrZfozC9xEkhJoXDgW6SWSAfJ+cN8XNcK9
IGrEOoJ5j8m9Amn1LxDn//xeahOCa6Ln3d8PQA98/UXyDd823PJo4lk0uN4d
gFBZ+Bqzqu7/9jTayxnLoKpJDf7CeUcIZTY0/X5RWgxeyBVOMqHy4AgtgpKH
KAbyAjm1Uo4KiU2GY2uPo3VOfFmldD5lTgpqXma47Y3IrdEKiXOKuM6qYHZE
zlkK5DRK+eLiide5KUYWl+/3+YFz4qWz3VgZ6INFFRgRDvQWk4ws7i8U6O1b
5NKvCUJmw3CSWv4vjBas8q/PlHGiQ45wPO72eigjw7bP7snJnM+GVn+hqi8X
oIBnZA2Y3N17bLGgGsLs5/MbyO/6pM0yhaOGSx2OWX5avxRpztZLRTu1Mu0O
Wa0+CmGF1dSM19s6/G/FZMkNpf5iRlXuAWNzq8DslXN+XoYzAnta60bmtSyZ
i2QnH3RQt2no1GONJ5dEwgufBATtzKunej865COeSR/Zo+OwhrICPrIWeJO3
4aq3037NA3f0mXhYferOF9ZrgeMlJol3ZeAxgQeERyJfIdC61FmaFH0mgWBD
ww0CvfPm8uovHTMK8wPa6Z0jBPb+97IqZcgin/hIxCGey+cCzTwTH1Ocxs9i
iO8Mqh80LVDcfGy1302cO17OOdZrG848oLjzHnFosqrITwA3gAxmQOMP0aQt
vZnMZwLLwQMtMlFm20a3FkZXUSjcvAcSQYh3cOmCt6mOAe0DF4mafx0nsEh3
S7cP27q20UddlZHPxVtlKUYvdO/qbr9dGKazCII6KLT8kp1U/dNQNSqU7VoY
kgq11pdUcne46o/Kk2pYsM66LysZbACOvX/YTj9VL0tgBK1X5HTq3p7tEBC9
cUuKJVHl8fjprV1pAJ+8xU9g4cBNh3dRjw1Bh7t88a53v/U6BzR2codNArX1
Pm80MpgTFKVJjtwV/NrfNv0YyRPLDLd2xd12noKT3FprBysiKXZTFaEUd/tD
Zw3W926NJ5xawU/VYQ+Pe2GrmMOvfF3DkMRiE2cFyxbFNnzIDEivre9EH0wW
URf6RQ865P7veE8YSK9XimawNqFdBZtlWKhAKhdsm74ZgeTfUfdyP2ugOG1M
NQ04p/4RJR3K/GfdCvFvcuFYBNtkM8V3niSyWIytrh6pAMFm/affgLcz8x0l
OiL7XRYozqrrrDwurAKvpMXUOVV8hfo6DN8h/d4pNeeNTdzgMQarVDZ9IlVA
5GAPglMuAH8huKnWclACvaXwt3v9obFesPRXnt58UvuuXo8afwy+AZh1gEDv
fnXNdDSuRkoRFnytSaY5Lu0FmZL0+eFnxLkHdhhOWvFpV9H4uYpEx+R/m3ba
mwCKn97PQAoCYdbdNiSJlfpGC6Pmsey5dwbFRwboic4hRVtO3GbnNFIcXJW/
hHGud86jOkrsImuY2Bt1lp4aHuIVBY7GMMfEBXQExoKq3RhRY+Az8ge0AIUx
+UEYpyd9a9q2pjbM4Op6h6KzWwtCrcE+Hq7s9qxVoZGedEJgqzpd4Xvr8dpy
mcV8fQJkPZNpTsaV+i2szr5N+F0P6CyHg2uq16CbX4LJ0UdjuiBPuDjm8UWl
nNxu4hqteU5KqUdzOWzCPrwSP++VkzHqY++kZz1SF6sGo94wLxqO0umTF4vo
mMyJWjaTVIznbKJnKhDHyTQRhTDSgmLSdpFqsU959drcIXAT9Ooi/YUpc7/E
NU3ozovjJ+mh7tlBMA9xc6awgI1mRU6+U6ipI1omlNuWENlOw+592pjb3eFY
l0kG1MTvJlVMQoSNVwsQTnUKDTBO5g7pPhoibd23VeEKj3i/VhtQ2TWeprwU
E/cFuF4OjQtPD9JMBqP7M84/eDBqj5C528zV1jBFIEw2QMdqnEDdK7LgQok8
HmT3S9CdIhjuiBYFdCqy+yUkuDAP/4cSHIFCpDQ8kkIoz/XvP/oqzoM3GAEk
qWBu9k8Ukg/rl9xyWciv41Y+06tZACoatRUAlSS4s2VkKCnWeHEombbQa22a
J1AHx55ksxGSldsOdXI4HtkW5ooIIwWiJItvDPA0knu0TTvWh8hL90EeWO78
TGOteKm2lVzFgKkwD4NaFc9CYRRYR1E7HoBK2ZZ60Uokbsq9NJrHI5AmA8ya
wIx6Z7RtZCb/FRXmgatV7Phm/pddhTBcL6lIW0B8ZFqWRZUP+iB3jdiGuNEC
mYnM1zifZQOO9YWUpisLC46srG//dA0Rfqqz4uu7YWbaA5hQXQTKkt08SIUw
9fQob1cWbToYKC632Y/JDVpzZHewX1T/JCwO07QfHkrDOLVcxtm79+rpbbqL
QPMR7jB2SMme1PgYlqLtnOt8k2IdCdmxSWS2pYXOuIazFgi1cn61lDwdJvHs
mkssFW8vUk2qTlQ6yUKzmloxV3M+bCGiS0E90cLGRbyZMBYgmm0zKyt+0OwO
xGmSutQor5I0sFI0bk0cv1csg6zSeKxnmZ7I0LnK2t6ymYnUoN65t/lsFgc7
y0V3cgy5ghDp7X48cSvsdltuBm+YoeV11u/SUVwOvVdrBwc6wyKXB/m96qjL
Ca4K6D76rI1BbLyE28HOrXCSkt9yh3PC52V+Qz2Dy9H+e5CFG936E4QuUIS9
n0wqoyMZ84idGkVdvZO26fbGWIM0KJn81DKwht4m/9UMPbDWHwnQXxJNnJdS
2ylWsz3doGewnkwKwiesId5x/emLdMN+G+LWllptcLmIqN1S25FCh20ROk/S
9CpEEvuCtzpOc2PBWD4Ngd49dJU5cIEv8ZD1Vv0ObBfLCqF7pw/BEiiLRN7z
RHl3H68aYrL8naF97bip+07brJ5bFY2fFsLnXZDyxX8w34SnTcFYJ7Yuv99t
fa+LKkVUwMdxWDx6W87wFbfvkOMy72XkzBUOq67sTIKdL3BnM60rMfa3NPS7
sFlCnlgGPG0nvNmjzaGxOAMShiu7hOONB6uFbCO3/qwy1zV7lnF2eSqT0a1o
89KCNSjQ+OWEexyg+ioJNaVOJyxAR+XoY2Lb4HXX8Hb1WpujSvn8JqDF3IPk
lc34+K0PTOtbiHa4sIej1iUBXdYxNNbi4PVySUG1GtHjJpkwzbNXXdgp8IAz
RgDuRWXmDujVzfMe/NzEGRRh74nA2hdfdb3u+9q9Yt+TdSzH8fpUaqcvLiou
+/WyxHydsB9JsoP8ilVERjO0aQNbUBnU0VTIQfDKM2bUaK+aC3z6MXod1/kX
xp4CkV+N0DSuBRmHLK/1ICdHosYUqdfBhtzj5qgFZBpKvlie0z0isaxYnCWA
hXAU7YDvWnZ6D+mUwn7jsPVRJ+O5lLYWZDusZ1DoLJoV8jHM3H9C6/iWOZIq
f5cGzo+aWlfOE08cyBEwYF5C5qAf7M6x55TfbNxBcNAD5TQbpqKReSjp+gW7
7GrAE42D3C5x1Mq1hx7C9O5kptCJyLPNoeecSxCF/XDMwma7aArpD104jmZi
t6dhEJr+tDspwla2FUvDE8B2C3SzDLUm/Ko9rGeB4E5lzbekga+TVdbp75BV
JbXzHvbDDVcJ+rvxZBfoqDHaKX1KSjTn3n5AbT3Y6S7NQLtVMVOIG0FHvB1i
W+GRnjYuVyizv7arCID6t5MZGKX3skRNGP184Ex1OU09AMAhGqQaU6S4BN7Y
ttvHyLMvlZtsknGeteDOdyl1O8se330p2IpFbfDfBq8Bz7yEeK33wrlhfFQ+
rdKhKdg3NZmdKkaC/W7rfbSiGyfzzNlXPtuf+VtNnUwOCU4N1g8Z5bDx+v9P
5JMFROINOYVs3LbKl81nmlZMLaQaLVl6jmv/QsquLeH4FuUNjXc+5zijoIZf
Jf+hbSiMP9UdaQ3GeSz4Tekl8njrkqMuAnA6SVqcgqK2uBYI67PPadq+YjoV
du/+hQxAd5Xa4ad14NWJHQjwGJKmnJErFjxnC0ruXWcg1yXSHIJ0NIVxd+Wf
zT1ecq/+Ab1a6KTqgytcN7PyXyNEec4FWx77tJppnxg2hDgncR81aYYkFlON
p7nfYdtdbLetA0yfEbyna2ndQRJkFa6SSPtsy9IFSzXecYCU5MGyj4UiMq0g
Kda5ueZ9uRzZCYBXt4fNz73i4gov/yW337pGIe4LdS/hbePxjFgtzVuiLxvn
8D+XBpDbyKTqxy/XecfM+4XTv2jpPEOdtT5WWtVzRnJ0e1oYC1FEwj1XmqCV
p6M1diK+xcnikeCWG/mGu5Zx/I1J6YGfNG85RdxLHmcKlv9H9ekHSVa/+bnC
auBbH7VfDCiQ/0mVUaHNsIQZZMgJ0n9HhLliSNtfwKl5knx6ZVleLAUtVl2d
xa1YnHgejfSTJKKQyMwOVJUi/gL3SYArIW8XEy+ePyHw9og/UoVF/QrAyQwH
m16z6sP0aayOnNy6OM/Y2yYcFZ8w3ouH5ry201JRz5MDGp6Nu9PCjzfGttuo
AY6OrFr5iuJ31P1hRaI59eIMRPNt30Kqhq0HZ21tZ4/QxEC7yyEnVHgoOJ4D
t01RyYBgPJHnNYuNSsw3T17VGqWsjQeehun+mi5k+mt5CumNgnix9pzoN4UK
kq60HOZkks85m50vd7hDX+M/QJxb+FP+Xr2FiCtha+RN2R2gzPi8/rlKQdKh
1VXDhMYBeLrBC3Gvwg8IUG04PXEtuRd+lCb4BTfRRs3jODVebh4UcZaXbFAs
C7mjZVmL0unvNdrcgfzTVRwFve+Wp5JwUpp28KPcuxVy6O22OFgynFHdzjr9
DG/ajDopB0u1J40UHkUXt3saB8v+TaTOxX12xPSv4oyu++VoRKptVFxuSlGc
oSJ+8q0ELboY/J/KFIn0djgryup5HwH9X3N4W14fBNPs5QhCn0ziSijOZinq
oAD9vrKDwrgSZP5tcnws3WfsInhJ0g/uyL+V5AKU5gg6XQC8SLPux6BgCyk3
1uDEBKHx3E/li6C1eV3at/qbW5tpCty1uRah1x5qDgknaSgJnsAo6NpW+Ryy
XqrQxcrdSiEfK7bbcTHLVPCDaoATAptB8ObEh9UWZY4qc1KvAvcbd56rEr32
wtvbF9g7bVLCoEtffJEKaBG9Mwm+4XJ83dAWrO6tklRmAhW6iTdExhcubWBy
l5ptMPXRgd/1tdUSUQPIa7MI4p+nZXlIX/6w47qNc6k8xhAvaWaVf05yDbR1
gaz92MSRsJCzdr1ve9M7fch6qqCIS3IgYsLF9ISTyEsqFSjD7JYeORPm08+P
rFBryUEtLKO8Rm3D2QLWAYMjeVCL+ipVIs+1fy5RKtHOaT5NcQsfd6oZWqyA
3DoKEPTAHhAPWGevlNgcb9WaqzfOLheowr8NghW52w7KbdJnL2/gxnEYMrla
+iOIt5nydNQGiMW1R28pMud5mdzBjwqc3kyfvwdn0EOoh4rfzMGTCQkGadzw
dAgPX6Pv1zDuXmoavn9vlbyHVU00EF0Ub1vTiELpCLSx2CWy6xNemYWQDmUl
lQYokBKKNoq8CUR5A4iPid1t5VyEPbc97uXxQcCJsx0d+PFkKE/qKRETIct6
auaNKsUxkaVopjbVjYZGfENjdwOG+ujUulxP6rPaLNi+KfTfrQAPAr83PVNV
ONix4WTE1QunxaEF90vF3hlKNc2kshEbUp4ixe5B15in5mqpdYDCiUkp70oJ
lI6MdsY00lgvxGRaOYzGHQqnQwZC30+gEuYcjakP0KETggQin2WTfdTym7+q
d8yNpiBjT/1+nOjHJLWTDREkfJNZJC0j31fObgaFUCu3H16ztgOM1zmEUMrX
hNigMIYUobYZ8YoSox1UyXuQZNkvuvtTY2ju9mzYbobRR9s9ld2CR86Mel0D
cGY/np5rCBkSpY2uYiT7EwJYcAhCi0XqqkGjCS0eALSEIM6wt9Jbb7/d2GYU
WKfVqAKU/VwNO1Y/fOweqQGGBBgrNcbbp1kITZWc3h5e6zcoZOunIPyxVNNq
6dy09a6zrz7d03u8LICnvltepxy3Q7ImuthM7N4/fyQaKFhDg2THDaSK20ru
l2UeTEs4HeG/zOoA4h1yuuGVsagWvvQMaouYroqiM/AoNu8QGlnWS8TS5F99
/s7A+mkSL1JupKdgqxYFK9L8WUKQlW15ySBHXSpbgCsUe1dPXLUS5f5oC/Bk
LbL4To3Z2rcvW82T2I1m88b3I1mc+rLnFDHUAlDA3fBwtBKSfB/w9XIHLx+C
5nm7w2LUVsiKYgG3f33NjTpY6WBkmy8FJWWWcNiX9k4I6bMKems1F2qEobBA
kgn8GWTp0eaPhByTFQtm9o6vfIhho8J76TIEQyrphajcO9p73MJ9gN2+cqPh
h9mJ5K7Ic6Pzsde6XBUHvSU+mfBCGKTxkYpmHAAX7tv3pzEMmbkKCmwfKBws
Wsu401ZdUUulblv+wBHyENyHTFOSV9O/XkoRsXiZCqXfUIcvLV4pP3WW4uS3
AHqAEJSvcnYpDDz1dlYpj7bk4D+T/KSMysIPgUMQnFeiLCXls5Z75gNGYGIr
HZKpeiqRl4bnjKGpY1JERIjkOoIYP5s1Z9oroUoMcDy5p9kTASUUrYFqW3vV
AVYFG6osd+FSRDBPCsvar0MolKY69qMItbCjObN1P1H+M84WuSpD4gQTfgaH
63yDQG8e8rusJ/AfasRT5spv4iWTMQk3SW6xZ7zK1vZSZhxTGY3TgSbKpGVK
3+nP8Z7XQHr5uJtLgpqe/qagdXis7WOgxjts+3Tk9EzlK/sTrdF5kKda4t7D
SXodzSivm+WDqlIJMvaKy2WuoBRahiJGF92DsfZIzdaSVYOqFQmo43NW8BoJ
K6TSoJvAFOljApU4nJy5I3RxMGb3arYcxcLMv6H4ThWBFqNvhCb5Hm13WWhT
a4L+vCBc1FDZOqTUqYb/Rwyh19SkHqQsTUMs9FQ3y0k/KgOhQxLhDcEC6jkc
ISMplBe2r+6NiDc8h+vT/kOBrS9A06xu38QO373x/Uv2rmuy+2nfMe//if8y
rrxOm5TNRz7k65vG0AFl4vrjl8iKC0OoHb05r3MtdLi/1kK0nc/jcsrj0eTV
nkbzG7ThmnDtnqXVTk36ZGHLC5NTD5JHrpP1JiCovGbc11cLv/IJ5rqFhR/N
gqUl1hMwSDPtaXQ2EVA5PSTsGfVDSJn5sKn4lHusPPc7s+n4FBxTwnz2N6Gp
Vv1oYUIcA4PkRV9x/CXdI27uf4+J9o068GH+fbg0bfjbk7nTUYkEWIsSCZQS
izVFw3mf/oDeksltUvMuWn+HtQVEj3wMFBB8I8YSc+S8PY3+FfNAcrotKMNi
US8ev6yApEyVC5/E5ivDSrXUTA0/A8bp0ro3QdYOyubp4I/AKeaEE3KpgdNN
+9/khicykyDFMSBnaQ7Mi9NK+2k3EkP9gPQN5vE4q6qID+Ai316MzBVH2mz4
T20oJhcFjDiyVJWqxFENCi6Z850IgndbEuB7C2b7oz69ZlHkDXkxttPWOAAU
5GZw5Xx44hjAodYCOdh/KKkdSXZoq/47irI6CZc7oahi049aBKRUdWHj/F6K
LOd80JeduPKZRFPQ3t5Z6LOvE+WAgvQfIry+V5hlZM5eJ+lMIAyVveUdm0j+
0oVgF03iA9wcellU1i53dBCMtzAGut/BhRn3obneANlPENwxpZuQoycMaDRQ
AuJLTXucxfoS2XCbmwSU7bWfy3/rd5AzO0W54Bt9G/ZExYLRuZLbz6Lldvo+
6RuI6SIXTodxNpUmjvqL4GS/NBtX0orUjtWRYnwJBlqbI7oYUyiIza5EE4hZ
lZ1fa0XBdfT1sG4vCxQ32eS7xvevI5/FZ70inXz9qOgoSI9kxLM5wvPKVSmH
1OTnInqUM7TOlZlzhgwzFu52iordPjBTb2Nl3esxKQhE6GVcsupk9A4tC67G
iyAC9bUILi4qUL02VN7TMRLehE6+fBpcBXgIJGD7EEAoLQl8LOoYJWmn3xIh
4/v2EF3XZL6b++FLW0wY9nl/qrrfns6yk0nfrFQUJNAsFGARgnQhqEpgxq/3
PL584E9J3gnHzRxGpotmSm7XevDKz+YB4kQ7rQObG/d09wFIMC3X4yNQnMLW
M/Mk7c0AJQ3pXeE5gWqol/zSIbPylW6Aujy1yXChFHoehv5rxW2comYzCEmC
tzamZQMr6idGOZb/IBXswSXsiMD04hCSQXNi0F7Fi/EkPCyCehGy675g5Xic
oTUQ/zy066OCR7UEfrKtrVUm1XPFcijZdzaDAm/CKlS3C169hbHWOlG7MbYd
g7yZAjDZZNYkFQVtVDtGuSZvtn3S4tUaCf+HZfQYyLSTSYsYlwW8C3AH+eZj
UxuMOLWxHTMW0q574p20uN570e/5pWF2PwRJEg3EbqEz8FGMPm2TA2YF5Wbm
C2tVkyvlKhHw2JH+FvI6lgOChGGih2zgTh1syQMm2A2aq66n+FpFh5MP6SDM
YUu2OxtXkO+OmSNLjcMbsSlnGhIIX2hS3uRRzGSyioKaff5DNR7i0NaAOVSP
q1pkX2FPW1XmmEbxZlcMaDNLFd6vLnAW2wx2mw7a69L+R11WRBwVUi5J0fqt
YrFDtilAXOedU2itTrnnu4s0PlNotekCwn/z7Yzo/VluZe35axqBjcnOwgVt
IbzKH+gmZI2LVP0f//Iyd4kdEPRDHovaFsPqkOFEFf48CRuJ8Phz9I2IFd9h
I2fAYQeYZl2INH/BwysOTGueZmI9I+XBHnvF95GXOVt+ETmMow8td0kPVtWB
8nJlgZngZCraBfKzsp/h6rJNCH2js6x23xrtcVycpj7WIsTUJPdcJKGvdeT/
CRws2ov+dGIwBYvu6480pETHkhcUgrHndsH5+uMKzSg5ecc1/8ZlKKDa4iUM
kR9f/Y5P1u8VjZcu5A7QZTJIvW0kRShOpV2bHegoFc2cml+0BRX+ilWw5Y+I
RYNN7nurYbyI6eAJdniloCEoInUwTT+48nRQBblbcqpPQ8mvHEXRWTZTJJ87
LYvlz0ppccC2aP4k0lJOBj/03L8drxuJJRwzIsynO7fpVWjRGT/d5itFKX34
KlVWcQndljMtNR2LVid23JjAyFx9KSbt7ByI6BLwZ16GNCKkHt/XoRdSlSVJ
eGdqlHcwKK6eborCbXQEatEkf3sCGdr4lgbm/15hg65jt/+T1DgnY0ae3SF8
owrSwWgwmulwnv7RNrDkIw/F5Hsy/RVOKLa+P5OJi2jdPk1EuJWqO67HrOMa
dXItCLS70nf1A0/zPfuh6JUoyVCiafuwyVhaU8cOBQhvBqz+daYZaLuc7AKn
nc5vE2tFPs/kptgFZCuXbZ4avZw1XpgtBMs2nqOe8ZpbyRK367ftx6aqnbrX
m98p27UdzX9MI/Bh7Y7DULeSR2rMDkMSDgndXEd7fZ4doZKgIMIc38ZDL2WR
2ko/Yi4Quo5J9CkK+OHAa3mw7sCq7tbWV37FPV2jBRMlXfbaZMgf9NFNh5qv
431uOo6QriyOuRnYcBYNRp1m6uXO3J+1l7KoMytuQoywaNc46Q8PJ38GpVy0
fnAxZMG6UuxbNtfVLydD/6HK+sOu4GHZI5fl2DZ9mUqkKrDX7yORWxBkuiWg
WyJWBNwl8fVOcQ8AE2tCY0yl17/nmFhx7H11b6SuRYA4+fj518b5ebUH//H7
rMddUpDf0tTg71Rv0r+TbXGs0GsOEO/pEyiks/VoilYkcVf80gbxVZeJBB/7
X0HKxekIjEzC9rZ8RJU+5B5Y3gHufVKcBgQJ4ZFpVdg+3MFXMvnubaFfyZzm
ziIn6VCNzQZE+WnERE10u3j+qpZizUfmWC+sHcfsKfnAgr15TdeTyu7rVEsK
s+m0GWiwIlORz1oX6uS6YV9gYxDP/JAtbuksd/ce0KVD3KsZ8BiKfTivUdh7
i9nDw08Zh68hBAgiHIggjma69dXtKnPytBNY4CcXRNI05ZArSxYqMMQRAJm4
F2RYhh6eRW/2w5gXPhj/Lqqaa+6GZmFTWcYIfLhipvZ7gZ5zi/uQgRXxhOhW
NGrKU20PzyDN02h8fsP64nxFWxjUaXBkU361FLtvfrmjM6w3cavayodSTMIQ
Fg85YTVKUhAPp/MKx0gMWVvL6y26e9j0SSgyzZC9aE1kFaVIppLnK5Xfs6oF
2E1W+I1fSIpSaNC/AR2EB6IqjqtFmAD2oVdswheNYBKqglxQdrrYiWJPbrNy
tbufGJ4QCWuzouip8XOJmii2h4nPyDYTfSRjTQqgzAevcAV8AaBVj9vE8E++
72EX2MLl4sssk3dG8geyuZeviLitSzjlhPbMNSkG3U7mNr17eWHNriSjFZ+y
JmOUf6H2UszWrdUg9JpOfVQ7EdOuZ9xOCsQEtQRNtwGneGYWf4k1B9GfrY3v
mWk83cJS3tj4UQ5LICASsCTWC+aHLbyfCEmMCHrn/WA6e93KbalFSfiPxAuI
Sh7TR2BURd6Qf80Sh9SnbP29ECZO83HfRRQgPtitp//ghQa7Ffwb++xo59Sd
vhVC91JdT3Su8sWwJeK1hum15mWhgWTEjsvJ8iSMXcBoZEYLKkwAGL/MIjzk
Vn2mKXge378b4/OONO3L1LyJ9WCr3Oph323tCRKe+9IHhbvrf8f5+ue3TI2k
KSpHpwZhXbtYgRchiR85/1whFlLTSbXQxGeUwmfjPaCGqGjFSsTBJEw0Cz1X
cWLwDWY5Sa6sNHNj3BMN3no3sUYwcsVNoJASkgDgaPHh3wcXK9hSW7psn8me
GgWSB1HZjF0L9fh1fyYcg+wA0q57xT+zKVmuYMB7muY1FY7XkMLq48KsS/cM
D3k6eqjH5FGcRLAkusI6APym41MpTNYYw91Ow1PMAqbwjOu9Ev/JLlkT3085
dI5R0I839FrdfScy8V4IU2c2oKAG4LeWnH3cuOcWXwbrfYQ6P94F4XLdsyS3
+fI9/YWGeMJImXRfNAnFjPU1GumIPvE4unOGc1AJTZO1jAekzMKjHLQ6SD5l
UNhP2R4PfPyhYCk0EETax7i5CuYs37vyyBy2NtmEOX8V9cL50pMkGxEhPckL
Kr6JDJkpRD3s8a8ufLJkxnCuEslvu1Pv1oFLlVUoOy2gm7Q7e0BIT6hgZ43A
htjP0JXidlRvi48GFtoUXKTQEygOpAXCvA1iwJMPPb68tFnsMgz4WTB2DKrO
Q6qVAQp0zVSZjKoF3Ys1NJdEdnmPTzyewMplFlJzIhCVcWMkO5tGdxRcgUaF
RmtgH5PW+tG166t4U+ypAcEsOgS1L8LmIwEklpL6MhUDa8vrqzymoEU0Yki1
9N+VskELIzVSseWqTeTQZHHJru5FXXLX9nIHKdPaz6k8tXjheOusLCx5TddV
jeqejTqE/gm39y4oT+JHNRZUJJbEOuR/drbalvmjh161nTJxoAcE9l8Hhpl/
q9HKG6IHIcjSUgADa+0Tq9vfADw1kx7jTEx0P16JmCC0wkjc98bksTp4ykDl
RPigOkDQuII5rmG9tuvyrId6Ygeh/Bj2ZxCG2RfIzS/x3xBwixi+h7h6ExHF
QZJeLnifzLWzPozJpq3kGydGRj9ls+ySysam2t1NLo86XtU1G/rUNataIceZ
nF2gU+EBeDoyyWghnSsHQqncQjzrIGJtUzEotdU9QMToehIWpjBX8jaNUPpg
6LIO2r9kM+BJlE+U+Y0L30vG+Q4sJzawYYLCYlfIMj1kk89qArkoHZTuIH4F
+YYw01ufx0lnfWC+us9yWCCFTC0YgoDUxQlZSEwLJYQSB332jyQqp08bjXXG
INh4Qg5NrxFHSYfwi8AFVgGu6XxwHzIe3Eq5UVuPtwKQWaT8kQKlVEkBSiSV
ZKyN6mYQ6pVjlTQifyd/MfQL8eiAh6huc1hiM2LtKgQ586KFBHxtk0oiOHTa
o0bDXx8LZEKXhPgFF/bEyy9nJwHOnegiO2VsE9Fgy3nf4qhMf9fLOk/CFN8O
6LtSZr/2L7zkaJ++pcU0AFyOByn8dDbBQg4Aw1/CQwFEvg0AtGuY9emdoyP2
lryhaOeUb3yvJyUKk5Zcy4p+sy1li30laZwwosT5cX7xG/nydy1i26S4OglH
kqCKZYv3PBqQmd3eVU9vT4YqsjryDz8yJFbcvfDqFzczcGTuR/gvak62VhTQ
V+2mMz1J8tErLEfYgYQAYQS7FAT+El2jTqlJvrchy+DHgc2JzM7zXFPJNJ1E
NloO6Urd7qBvockNp2PZxhLZng10q/78IerbZipznGq19RY8lrOLOSOqZ0LH
NO92GNgec8ebyfSipIMLKomKodPOs5vgHScyM3dPEcneA9TzZ0cocvVXSw+l
xLCd0SkN0c/Dmuwv1InDKl2Qu2yOYTtjrb0NHXk/pu5Prqe6x9CVn+jHaXWw
6xREFr/xnH60AQRpBh0bOyPhyRtKlJERINT32JsjHzaTqYFiJV2l/lK39u7j
AruKoJyPPAJG69T1+HYAT8qaR7L76RCcT+vYwg+iu31YALXg3VeaqYghiQag
H4B2CrB57rCQRAb5sA4acNuJAASHEs/EIxcnx5KWB0WsXi03nulIlo5ouVXi
Z/qUy8XxcyqhXVQeVfbINHTW0sbUmW4BGRb6DB+XIsd34MO23MDiP7caw3ND
7eNJv4raFivP4ecbRUnLkWSjP2qek23n88LnQUe8/xoe+lHgJ4ex0ue4Crva
LGVIEjhR95AtpKQ23mfy8ClWH3Kw/RdIT/m0aLmoTWMoTDZXJRDURs+zMo53
B5i0wXlWy/BBwHla2xGDBScrARqi7IPfnCsUhMXT5jKSDpQEH9FyhVcF3Bde
XawIj98oaDwMRIOV6X5738u5AsJsyIa44HXTYTc0VB5ZtXoY3SpujZWkD1Ld
q6JiQXocD3Bkt/QRt5xA2We6kQCvjhHB8TjYu2+mBgajmrAGHmQ5r8w68FxC
P1yFU/1XSiqcuANm36/K+RUGOVEL/ZwVtAWJrIbwmOkUsFhpWbUYVx4afD4/
ydZk89e1eyaMzAZbyYW8sSBZLCCfKcSZV1SUjaHZTS3mmhlBS4D0K2l4OoJM
6inATJe/3nIuAtMHVmnLbwH5wINZI8oyUTQ5x2ziaF2Spq8fcLo40BKp3sly
7uwFL9LFL9uTW3U3v8G6DF2oTc8a+zuIV5rescHbmEV2IOByk3gbzZK6IB2w
n+Oa8bMaSI0T/FuprB5IPqc1Qv7dYKYBZ55A+dWs7WNjxXIy0nCtdvCRUtIn
mARQtX1GiWZXQAkgAdxaQwj0DsW9G0wPjvfIGrE4u94olvIUldtoHUdEuxEl
a7Pf9Y4UUUlhdq8B3Eq9rfXG9J74R1h9haZJlWLZkeiPLUeUa2m/ZHxLH0Ya
5bTkNqkwXqJzAzxGlNO3JeZ6peg0Mpma4JGEg08cetxYrF7r/LQbFlzjez6o
Li1KY7PLEEepi9u9IEPvaLOd1AwZ5zNl8dAwg7aU8HbEWSTp+kB5nIh9hSEs
Jv/+usA6tBntE6bdFhunbCghk0lzWDXBtybSJeQGXI97lbiTFKy4UTjIX1p3
grsSkU9Y9B3mon++ROBkfadr5BjxwkNkXoaSFLwYUoprvc29MoGKRMAhVQT2
dPWiyb3kPA9S3W/foru0By68xaO8LO1kBjpdTJdbHQckg994ZHJyMiPev2CD
Zhvc52PfhkuAWaWKGhGid8Tf8mc6tR0F3mSiDm17NDFSl2uWC2UvD7c03Z6E
gH0dFmodE5IepTHCaydSFYjz/ip/HFJrYmc9zFxfCHOi5z1rO1vLDWLcGugG
OmTolKpzMXRd+WVh020vMT/9vVd5RqHztEVsHvKgU43+0ja7xcymfDNZYMCR
z/UUC2fQhDzhrjwrm72w+QYjCmlmlgHnf6qgYXyBywulM5m5SCuGHhIQyg8E
OV+8NX8bTW2nbwHgPRzbXWvg2TAjCS95fSJcpM9zgLAcdJcK2VWpwCQDpoZI
KZyH7o93tP1FzD9AjBFNvaVdFWv1HSYDm6Umljgtzgs1hNacOotpiVvW5pEv
4MChI42ZNrEdrLZW4RwSU+i6kkxECEMAiariAnzGd8QPlRGQ1fYJX6eYT60p
6SkDZQFXpHHGtB/ssyB+xgWfHCO95ahypZMh5BW2PvrGq8OxD0biRj3IO5ZY
Iub3aoerKAQGh5inBTQh7PmnYXujJzew4OM3lE5RkSncuDPaAdTaaBZzNbxx
qvoYf86YiV6RVvueL6q9//qmhG/6lPHlAKIZgJh0rnoMnXU0WNFCs2GIXgqX
+G0SJ+SjrPcpq/+AjRFSucA5P4mpf5EiNDqkuC8ZtH2FNjvufSxgkNAmgIVC
TZuRgj4a8p23yzIQQhqdJtjAULBO8Czgrk1rZ5mraHV9dbREFT/xRpe+R4BN
kQ6h1FLQcnxSYXdaBjKAq2lFUzRr0hi2i3NqqMlL7n6NLhg3rsh8b+QWaMd3
xDEm5C7CRgZXRsRh7JttzveaPrtb/A3/YJhWf36qNsU6MPCrtlmyfkaT3jaC
ICiXBpeUx1H024a+9wpyuMYrvWeSR0AewhsfBq24xQZbugPIslGEFHT87S/j
LEd4kxow2OWpLNpldRSHhrFYrvBKvBF5ARXx5Pg8dy0QH6toejs4DdwMkFVz
9HBaJtH+VB7ns+T42cIDB9nApQQA9f9FvbYmrinUqtbz/5ov3TMkjlgT9gwi
JsP+Sv7/d6g3Z9zdLdkXa+YkzY1r4irmlbFn0F99IP6sDpthuQ1Q+n0sZkWt
jko5KwCFjAMaeK2mk+eBuzIhoGAH8DS7hoTcG1+c0ovhocBvR85gEaS/rkbM
SwLJg04gbYtltDOIjXV9xUnxkMp1R3c5CT/1jFCOTgodHpe+mTztSS1Qdsvi
Mttd9ge4A21/9nJfKUzLPibSXbkav1iLhXiFgFdM+jG+fk5JMFq0/XWYrC6d
C+d5PxArJ0yt5o9c+WmSIEsfCvR9W4wbQkAk6e89NvA/o3KW06bCQ4Bebn9H
B778ISRw+6cCv5O959hfeqShDbUM9bAw0niSoR0JsEoKT66+Mqyv04hQoXZs
9yir9ty56NbOukHhZh/AvbXPIonzgPmRZKDqiFzUENByA7/bd3odoLnjPiq3
Uvhifh9FlDVOuCIieR5zRVsDZNf4w7JSH2yOjZPbMbEympJ3pWQtxuFmtj9f
SDLaW3FpW448bgqA6rPQ8SApZD9K1n96luD9DW1kZpLYBxwlco+Y17gqHdGk
HCN5FCfRBvNxxBwyVxKBLPv/aZGYd5QQAY6GLdnf2p1yCiqk1tJOTSfvYr5P
l5R/G67PZ5mpMK5g4zCr+kYZrCX6KDw2+nXD/UU0kM+V0UQu4TNAL0WbWlSk
3f0tz2+GT4aB0QFtnEYtSY62yx87Ab0PhUz6sDKbaFxrnJ+rqOOY+ulUN6FF
YcPJBC62uEbqnE4f5IcE2a/DUxqFXLi+SLwzsLbA0qpopfHqhgSoKxuQZiJL
bYQJS/ir77diB5rWwbTbzoqPTy3s4nJLRyGlFhjztrXalJoLNzZJ+WqZruuJ
4G3UoctY0DqB1Ow0wctCC3klwbzD/twe1D7YA8KyZXl+9XU59579PS7PYOp1
fWRJ3Y5bUTsAT7GNqhdWSwBvBn2C2S7vy7AInTwiHpFpsbWjZk+oXg4C5U6z
cWmWjHYEdIQ9DZ40U8X2eTa6UgJu0CMY5h/cYC3Gz1GcSEK0Rrm965kGkJ/f
KfYb76blzs8mLDkkBBtEua7R6mU5V4RXAYfPdi8Qx9lXS2YA9LNIPGDtHXtJ
nTAfLBN7gmZC4qUXDqMSmLyp5AcFSrQ1tvxqwGb6uZXw3Qjv5whGSZPKe3ZY
fqvmknDWhZOssVc2iWK6Ya6rvRO5WzmG3I0q3+quVu4X401e0yLvh6BUbqiD
zBSIQn8DgHRs5Nrw40BxsBi88N/NNGq/GNnGSF+9I032cPkATGKnsFwS7Ndh
yFqqNL4Uz2aSSbwnfZuWTptREsTX0wO7agou1h7+LEcqTDKR8oEUpSARL7ud
xYfNrsVKOPtu3TjXul2erAMwGs8w+dQD7WDHH0SG5X8jHIyIxw4a8NXLs2rY
8uUhkFk083Zaw/R7t5D4tSVivhIjwQ1YOYFiQaInvCMy0nHBY/0+x6ZZuPNi
T5mstsq0aQ4vIt6lUmJlzCFXNpeun36aIBVZUWE4Z0Y3Exz71eXPzxuxlBTy
fFAG8YF9gUF7iM4M9g14zgNnrKUhYzZEbUnzdizhSCEPih9UmR7ONpb7N32X
2EOvn9/g4Ziuh0+CxN6ofUGv3T8F/41RFYghv946NajqrQPFxXFJ/gaymesE
g3xdL15pzKt6Ijjpl1LdASBXHIYGXWHvYNAy9duHcDQwfZy4716M/owdbQdD
8dmw7MAbSYS1lFxyYLKc3DXmKsLt5d8XEigDkJmEthICdiOoNDfLXvAgjIN1
xgaUz5Td81jT+b5Efdf7kMUfYjEC8NqqdLChT4LXRBgmORamHfHwtk18QilB
eiPLd2JZJcJ2un+diuhol8DYSkG0c0DHR5pM/MN3Wawm4pnNAtq98e13SiSD
Xaqa3mgetnSGElvgF56vkb/RfRAQ50RRK08t0DwKqJy5OYGc3MDhOPdruiBp
JSupB3qFBpLMxx4Jl67gnxSXKrL4mpyJ30mEmdZl169NldJQ76H0xYXWK+cC
PsrL17ReYlJBE5UmOGtv1oEPCDLQufd3lcAxa4CkUnrKBokRbmySgbxOaicD
Wy7fqMRYDciFmVu0BOF0mk7NgVoG7gW6umycpWjfjMQ+oadmQBBhbGd/498H
+v7v9cnzKMk3ZTCCDiA0rjS+0JYdMijnITVHn1EYdrj0BRefgZ7u3iphY6mb
aLNh9O6Ek0r0QTxe8aZBUl+vQM4O5ImBKIj668lkFRIiqnqOiK1l9nXXPTp6
9MoU2mHdGjAJIE25rpQdmCiNdjvfEuJvOYo3RHkWJ8Ncehpa2AitFsotdsxi
hYf+tdP5BCYGooZl0b9+j46kjnBI6PEVurBq7FuLLvqE6akeygQFVBpWQ7qL
j5hD6B4y7x5Govn2ixgMKPm84ZqULupx6S+U7Iu1ecVKbOV9jWVyEXa+ehXQ
2VaFjGOWavhWK04iiRs52jyrBc7SBSidUlp7tIMg2zFpbld3jEUujFy25BS1
/DFqWwaYBu+NODqgUVyd+6Cf1TJe1cWVQftlCLc1+IL3K1iK8K58yj6c33Ov
Rq6xMKsgy6iSLa42/b6iwJbCosz8pLnDJSdLBVD1KsIHgZXEcpGABxSR10t8
SP8DjW149w2BeM+lz0xwaXJERGj/XzhivpWCnjFInpTeoZafF/DNzhT95NHm
Xve+QaDgwK1BUMQD07sTqsUXbRDUxTIKywaOkcQ/JEmBNt1pWURBLn/Eouhj
keD374QzQSkIntnT4/k4ZEa3SIFgBL74KgjmUlyFwNGGPmqDcCftlTGnq10z
udjN0lmRpFIMW9W9abkzG1Z+YadCFzF9VdfflPcQT95CDCKoqy2VjAgqKNOe
axX0ypLQKBD55iF1Q5k74t46GbUADrqK18UL9C7VSzZqJrhQShR4/yhHlGes
TUUgLowu3OvDXZ3r1buJwVBkRKy3l2iqI5NfUZVnjIDhRiTDZgWEbErpAGpt
cWWW4KQp2mUKvZ8u7VQ8eZ16yX0toljquZm9Z3VmJjsfU1rrjFu1t9Knzp28
vNaNCYh5QPLFpZCWaEj8VUudZIKANDLfJCRlIoCnxF+VCgykqBMEwRgoBBCM
ofrwUhTl36tREqws+WpDbi73EcXiBlYs13wOjMiLAjNlqbxk/vnuQdae/2Qj
gjvckAu4vPeyBKM+Jw2OjqLKOSqrOX9ZHOSDQH5j6BbXpss3fR1aQndDi7RU
QRHbhQsBZYJHMPFzXdrcta/GhBuExTLV3n2iKaUIRmzDQ3k4WTU+jHdDTUQC
vMSQU/LNT2IHm9hc5lAqLAkEdbTpMVd8QcuuvTdiKhKkpLcKNPFyy1Fy0B1S
3YAxccr/916OVsCfETJX/bA7uAysRzKgc69GFX30A8BTe5tPQtAVAVgMLRJj
l7p37jh40xuCO6MjQuu1qWLUIRjGgk7IPLQs3kYEhhwbNvKR0iAQZqM0KOtF
mqdSxciKHhEze7D6F9vW/DBQPu/Uz4CffA2Z4ajDmcye75OXRuqJbmkXSMP+
mG4pijflrKSW7QidZ39Cibn1bmvLXG715PCT9K8nF1GA0aCvpxTmhA+T0Td7
JxQWaq4nH++VKldqnRGyEFajeCR7XO9jj1BBHYmKHnAaTkaLLOiCYGJNMNO6
TOSBS5bMv2G+DsQHz7kSj9t8PvRW9dM0gwzSM/ClFLBr1MBisypHNeIHOna5
9dvc1g2CFfxiiqwfoU+nJLYwoB1bxKdS5EB+z3ORdTug1ZrHytr8ZM1WWXDD
kOQTTJh0iCievIzbmiM/pyjUiLkoB6DZUBjYWDilJUykXloQOAb4Nx06Dv8m
Zkfc+UbnoeGYW9OjaZcv1coUg8PCumsYiWwo1UNmG9WSMoS9QRPO/WH+2nY9
94MMy+iaL49FNJxpJOlfBEaOcawtzP6k6ddPM0IF5dHIuDUMWd+HGOEyEnEx
qpWooRYPuXceD/+BUP6hkfSz0EBWPVHkCcCPZc0vGstNKs8knJ9Zeh+nKoCZ
YXnURBlkLYeqK/yLkKcwQJTW5fWHjcyzXMZ9uPsGiHmAwkY+0AGS181wCKYX
6yylfZnnoQ2oAnCMWvYuYp5MMndukEN0Gz2ZMPwLk3yyNHe4xd8OT+MFS2lU
7HiYaTo3SwxYe/1xZ+5p+HiLR3g3Y07KdNq2dNUHpEFKe8w8Qg47Jx7jh9Qg
dvM1TdUsiPbZB5UeLLPO68fs3I5NSXdrUENtMiwuKfXefJr6N77GBm1THzRh
LK9aYCYnE8BFN9kn1tRr7DvzUciHeUZ5Umnz2mt/MeDFOZ8gE6pKs3yp2Wol
h393hCeqULGavX4APMn8uQwPQXlMbucQwbUOU7d8pIDrE/mFcgmxzK9UzD/e
IK6czREJQA+rae4l8ZHYk/yjOj9pU6nGZS0dM738vvJP5//hlkl9sKt3hULi
GSbysAT0Ca2R/lmUHgg8+B5FNIXS3vsPLhEaxMqMHAQnajXYIplsGYUiMTwe
PkK7zn99eF7rblZ4gztE7uo2hAZt31SWEMgwp3xWTnmjPzw02jgOOrLF2lpo
BTxDAw/p5J/pOBJeOpf7zh3X5LGUZnMTyU3e1eSZxBsv2vE81gAAt4HBXjNc
G988poC78kychjzQuDNix4/B12zffzd7wldvULZf9v8Dx0O0xWYf3gr7+DTn
mrIEXN3Jal9N9pevodQNSYjVIJiuZyqMokzoMTS650leuVnZItZazMC5X3Rl
sAbZW/jpdRS7MErfbrsnTcvrikOnDFqHt2JYZbw04rx+aX6qMBxEYHp+TK6X
MN+KucV+mbmJie3V4V/DRRsvxbjckUHo6DEnhSLBXyt3kXYVZsBE8slK57ww
Tcuup0Fxg6FbiibZha1x+eYEjBAGDTD6lMLgbOfxMfOo/AlEnSXCOsjEGdjb
LYekwzfK64KORLkMdjETVkcnKH+l5gy4C/7Z6UGCjDQEzv/W43g6z0RzkNao
lhpQea2Z3lq4IvZ3+MzRalWjbkVXL/Ejiylfk/Fvr3flh9pRjrB72SoMXXKw
v6+7b69LdzwJSOl0gVUhKB+5TqF6AG6515GFpvyV8xX3kMuZTBlJFx8NNteX
FnDEOIJ2C04HtaOlMufOBmEttB2BJHcT/kL2xHkDo08yroVX/Ll8ZhqNeYG5
q/9vsVg+EpU9eTHJ7EiIZ9nciTaIdL9SbyqaUaKPaa3+EQt1fBSx0vNlDlUm
Zuu4UkulSRfU5dCmX7TU702Gu4chSuZ7i1VkOCTs2PAfhwAe7AmtKpGASNnI
hybInKifmt0WXitJ4rNc2LmasAKXD70XT6QE4xhbMJgvKpGkvKrGzA6EyRxc
e2gljopWFgQZ3Pmig1/Vh99DXO9fidMbm7TBGYMMD71wOg+BBS3TzVgdvNWP
QzWTj+K/yE+wJMZX4arM6GdrjJlawBFHHrdulMabTNXtjar1ZV3fTnDPN0ME
B+iJC1gvmE4Tz7QNyaG1u9S39dppM09loJSgVKDaFHqGP2F7GkY0fyunO6WE
7KG1NutiZvDQwq85mjQ0exhwCRSBh/3aBNHSv6a18v/hP/AH1sLYcWXzEg+R
efQSaiFCIkZHVj5AwFKBoi7OjzHL236v60DY5W+8dO+N2pvsXxgHTh+6MYGJ
1aIWmjZhoTrVyvU/FBnAUV63d88h/fOhtreCKsL4q0W9LP3tMOKrKzWvuJ9X
miIg+WIIfN7gKCFoFys/MJs5RYzxXaDtq0fFWsvd1vObh2/X4EX8YQtuNTZX
duYskPjaGU3Vc2vppw8fKtuAuZUnWfptKxT2QjiZRe72Uev4Ig/xv2214YBT
x0/tc9HLm1lBkPoy9E5sZnXBWehQpVm5EvS8rceKMpe3VdGWb9yChmmO/Kxn
b5nOo1Qvom6OBY1LWYqSXt+cG6b8kGiLt1Xvn2dbC3l59XI8iKVwOv47z6j2
N5P7yofM0NMuRH3wvkB9+e67OAjmDR175ZTXk34NZgwiVr8CMvVUtCAmoic1
ihXs/F4rwYbKkMsrQdPAS2hvv+0ymHiH1xgZ/XdypLiXZ8jfYCHuNuJxy/IK
oyCq9DCuKZNYwgzei/yypHOmgKWoMQ6tiIgArXM9bkFO+irYU590DNXRvNBZ
MYkmYAdgBvYQWGeHoVbyCuNm/TYF8yClIG/LYV023mQv4XI/N47x2wkvG1sj
W/31eUJkIc4QDCEjjOHyqNBB5Mxk9yst7YDbPvYB7gmAdewl0fUfLfls11vy
vzx3+rBrMNFN3ISDiPFZtVJFkPXn0FMJ7Bl7Lebsa5YNXXz5Gqr3JyWcPZNq
o/0FpJ7F42fsl1A1zi6MY8fppAAMpd7mbSQ92nh07cwkXeINqkghlhX9fFGa
V5N/2bylqYoYlkT2wQD+/WPUgOziCUmUs2bKdamN0U564HldCWow+pHNj4Bk
h9d21QD/935S++O3xJa98mT3kLGnVt/YOZ+UQ47/1mWpoNcjlVAfIuFlr5X1
A4QKTb8SDS+KtMYnkfwjjrMwl4k/bWILJuJE8ShQHflMJWIutC+5+QopyblG
fI/6aaPYJZn7ae0ikUwe4vCJsBUXegz963EWRhRcqD3rGmDIu6g8beAj9d/d
StcVpEY0+H96+tx/PJ9MgCRLhaV+BpuQlEVdTKb37kAe01xioDYXCMJS9WwO
/ah3aS+qAUSIpO3ExBxjXuK3zSNdZtuZGc8Qo4DtHpIUbzDh0oIOsLc/S1rw
hBjmiCFKTeK8T9XMoXAsxXj9/vKHJJJRE5ZdNhL/DEv6FKiDscAsTL3zHGIW
zITlFey6p0EhFqFe3L0IcZQtkcCtTma8V0WtWwSxpOnzxnTqcPKloifxx4Al
6o692Ba/R8jGkmpipsJELMvgzNZHpsBYmxtF/whNLAfkXWeq3Bo0AnVkPqxS
lrEulQlaX8zi9sum5a5FwbOFbi2vbhnk3dULirVHvPrl2BsCzCQAlkrX2q++
Es3119riov8FRf9a74Ra7846VNIKuVBgmo4IfZtQNmZnirLJgnklvRzPC/30
z98FN3Xr2Yv7zF5iUwogQwNfC2VkA8OAc7uptXXkkqyBIek6jgUyC85Wfi4O
Av/E3wNwNU7H9PMp+DuiME6WCym4TVp+MomIxl0szBNPHbPcAvOZqdBtclX/
+L0k0QsCzO4feaFwefUpjFvOMcT8K2Qs74JvKLc1rjt0Vrd9HCgK4vcUdkWe
HAa1Zv9lMVzGPtxGtu5QuTfSN1IsnAZFQvG/KEXGZGOZBLSvzInuA5lWn3OS
HRZW1Uq+EuH5rpkLBtfMKaxw2+Jr4+LYzv+RAbCFWeKDh9GF9Nc9zUMZqDNN
dWUMpX7ynTHI/BUA5vQxCWXQiEi//skq5rsdaG02UgJd5xseWE8YM/wtjM/0
cTXlgJqEPqP1c4YIewI4VUTHSAx2k+wcc9WklWTKPwlOHo5VUuCCGGbXk/Hl
f6rZ6W4h3aIo5YI5iO64poAsWdPOpQgWfn+zdw52wWpGN/D/a6ylPBk23qbg
vceCxJEbjqYdK7sc3T+wFli27GXZ5kCmPxmW9HWLrS/Zayq6S2tJnMijnsk6
k9XzmEh8px2gXQCfMtgzpl4o10gxDlJb1VbjPGAjD04vR7EA/bBtsjUkKr5V
wDy4qctcMWZpT0KoeAcEJRT3oJtzMhamV5LQAZ2fuLnGBTaBP6an9dkVmNrH
cDc8WfpuMRd4y7EzC8OuG6gAo/VHEtFH0JGcTpxdkh0ZlvryBPcLQ/DbvU3R
7NGl3BNS/DNJ4+56vafKpgOdm3wmCC4hohYDch6qyoD6pSAr8pPjzlOmVu2t
xIgpIZzzLI+SImfc+f7jrRE2mPBv7kzN57GMj8MSo4K6xIgZfufEhkXDf6fD
y67QbBzbKPSlmGooZZnWs0ve402OQoMDzjNXx71ru/TiwU2nIiLqVYT9xNCA
Qhvbemx6ZQRUjbFmwGZ5I/XetjOmhT01UZwzMRO/NmUQtxR9u6d9usf/Mraa
3LLLOkG64ml5P3rCe17Bz8R9hbSFGjbr930snm6uQ1J36mVbDY1XF3FtF5Nd
L256M/AZZCpEycZ1q+A11YwFSq7sulr9GTbpHvJgcOnd664TfDZ9AO7fOmgO
cJ/X8pmqwHfwPX77KE8YLK8gIozl9Wn9avvkL0lKvDpBjJYg0RN+W5vKt3ci
zB1RZD4sppp6+aZZ7Fbt6tIqPwL166qpk6odmoS38d9sZjjMaq2LLuk04et5
xIXcBD6JLrL34EClVGWN24Gwzz59cLcfDjTdKoTWDyaio+mUWpXdqippxEeV
nVjhfDO/bpHpVNJBw73PuUyme/6Z6jgaSmRNer7XdLixBjPxVlvKBRdusl8M
sfkpBAAFtP5p2zndaVYTT/wV7lYSOM4E2pEVwZxPru2VcBUU88I6bx1pynky
AxJ+eF+LG7gW3VpD30HAlhiF3BmT58yPu+iZNmFPjBUR3o8BZ9EzHodRH4N9
c0vvOaQYwO7L+IKTPAPCl56daeg9tzxCsm8+kWee5gYkM/7iWSdwcQzaNvTX
5zk+ewrNKXkBLWU2/MxcuxIe+S4ZH2PBSC/TpCHIMGvvXC5RYCJ7gLCwsvF2
+/mGsOfHzQlBbOZP0YlmA6jOXQWrHxzIG8Xi1Uz+BjE15nW6kGajardJyyF6
SLikUr8ZdjtmLjD/mfU/NbvmNZ3zqeFNoB9Aaf7e63lew68Amkyl2CQ8k3Tf
Opx5kDlBWXRYFCBZhNJ2mA6zbPM/96k6z1i+IiQZ5YR6tqV/6K9SMmocnK0X
eJpG0OvFqrDCUedQAxT8AUQXPtIEoj1Uq8Ar7nkAEfrfNFFbXxDLr7q+Z2Vo
LLrgaL/JqAph85raPq6zpW3OhsoXCm4AehHIPLFfjPx2w+J/FUjr3nUxpXfQ
nEZZLYSI16Ko20eVR38QnaDq0c6L5Kb9JdSKWHvShtGXQqNV+c/i2KKuba1M
eM5m3AOhRu/7UxbrNdj3b3U0XqVpQH8kU+WVzgbUC7YaVnRz9yA1f+7pGCqT
AIfSK6nK2+iBjKw9AQCDQdmOJVVR1TupCPvV0EZVzLh5cqX8IdssCvmufnmz
IjTTiSa86332POi/EupPROARcFtV99ThqqWuFTr3r/B+1/1BDllxqUtkl/q8
q1s2S4AL32X7s8vMsdnsWi38scJEZskAQOTbyZaBxqI+c/mIIlCAOqEbBT5E
lkJJh1X+ckyB0NWBnoAqDCUr63l0nd/z/JvHA6ut3GD4pL7JH3iHoFnK6fWO
tYNoxh54eGwMytr9GS1adFgd7EMJXPE1j0sYTTr53/sbeGfdesvO2uh4ggr5
0PRGrjkO3yfvA42N/Jd2jJNEOTFtDaOOhIEUkUKKZAn9NeA7WVgbcTdj3a7G
VyFN0zXwHELtaWOXQdo3hV9xlERmavbbTqMso3YdDmhf2MR3fKoMeMG/xayr
7cl8ufSWHzbNnrmpPf5cIkErU0gv1UF9npLaaRYc734pnug9cHV9uaCZn0rR
3z8cfUIBLU+a6FhsUw+EDMSwElQUeJVQWjrU3TKk3fIpzx+49HkcP+qoE1fQ
+0g9RosdH5KNW7jDPa1ucojMwTtndPcy3NTWJg0LTIWDQAntO6XzzNgia+0R
/vKYd1fKjYrXJg5l+UltP0rFPR1sbQracVEicY06DtBNgB/ufJrsAacByVd3
llK+GDqr4RwaAgtHRgRchqGsqaSXEmusAtcOJP2whRsJACYgTpJs2fQ4bGDP
QjPAyKTKpgA27EImI1/sEm7E8UlANZsk61Ol0JUJWq327yAy3MUIuYE6iR3j
ouFsH7JMMmNZbD21zFdrImO946Wi6sRa6deBiUzzUgUBn27Vs40KYIhfQ437
WWooVMQmDrCnpvsOLp/M6dfX/QN5e0qYmaREPokLmSXP7CJWn9cVkdOeJ6go
DvbQ36Ei/0NQc4tgPt03ZhAROTJpCXvDcmon1s5Gb9mhRBQaY1RtP970bqqX
ZEo2oGjU4eH1qeSGq1Any9AZenUAVYfPza5Hg1+UD4fPPfVfeBkqAzP3+jqh
Mh6Ye8hBtqKay2q5VkSDKLrc/Ng2JCstvaRW4/xgujG28lprYRvFKRvH2Lcm
l22tqiGHPDSp0trGrJmPuOo0GvD4C88Sq9iuYgTJ4Bjb7dehMHZ7HAaJ7+m/
1PAiEAVXbnvjqm6mnWBugmpmGhD4A67h0ECHUFQEcujMc0yV3BuQt6ULDI3B
npgRAEakDnfHoAZ3xfMaxwlXDM7oN3glzIZ+p4SLh5ha9Paer+O4JDWEIHkF
1u/jjGIO4bhuIik+gaftDbGzzhO/z2IPrw4MsYeQbjYiWZT6Fr4qukgpUR2/
5sH4TxRIAmmTbqfHTVS3ehXH4DEMFeb7sialPd4QMDC7TcfcZWWm8Ev6ZBbq
LAVRvoALjJ1KjP/23LtnYAZVFH42SnvtjiYEddy6jfBK4Q3F39gS+n+C/K4c
FqLkfp8g+hiA+uPECV9ytpwBzSuL7U7TH/RU5SnWw7D02ZsjDA+gsZxOjChJ
gyO2415wbvVvIXbBApbGnfk40bU/NA7XJBzArwl/ffdzVi0D+qLIrx3mGof8
Ww14W4m53liybYyWLsfKbbrOz6k/LNzXxVU3LVnPtc2WQTYWSSlXSiqAYoWU
ApVs9c7EODp7/fmEui+o+3Vh8ClT+1c7SkLzwHwJB9wAP1gAktePqWZ0gY4i
UfqUFwHojzfSKUivThmdRdYTvBdgxkAfdhn2hgESaHOK2dVlVL9InjKedWhf
pKE39q57ZaTICN341U5VkcN3Ock5GAeyJf/+2Ovs+kE7xB0m3zm2BLrV6tW+
EnGj7BJfa2EKD2ZbDv93SOj48Qd1c4We2LB/CwlxhvnINnNqH/gHBbSfzn6L
C2fLUTM9vXm1aAXi5QMZErE7O9zgYXkxyxd2JIuNk3K8QFOIMRgcADZd7toC
jUPMQrxRAz6xQGAFhBfjh8nco4lHvqU2PbyF4xH/Xox5J7I9GuyxRmwm0wDv
oj+JDeK44cz+d3rvcIyGTLN/KG8onkQ6C795kZ3v6qsvcKYL65h1OUbDloJM
hsERJcNRuLR5N6s1egE6HKgFgNda1+Jun5d1FwxvHbITNOgnfjG2bzXvneIt
rorQ6d6d1Ao3iGYwsIrutJuhX+rZ+cg2basJUAJW2OAUgl4+Pz1LF3gkC6dz
xzNJnGVToRlYs+89mF3VB2pr3SF2llMzNbxiPxQ1ajsoXl09smPM5rTtyneC
7iyDQUrkedn5AzjpOsPomvVCyYSmvaYl2/CwVfmSxEWTnkEKPd7kC4F9jUhQ
NK1n/NTROr4/EoIauPwqQcpuzOvmtvfEjz7PqCaxJX9XKgSQ8puPNlIY8f7f
yZAyhnS1JuF4YsV9bWw6W/lDLMfelmEsYBbgJLJa2m8OgwsIha/Tq5+Hwc+E
8/SX8zFHveW4zBDlIGhin/0dCsReF1r3IlZE5/QRm3yeRYUD63hBae+BXSvs
XGqCx1vk6+CAgJwglR2VyFYDtjHSKXDeuB1nIB7/kWPYwC0H9xoOX7KqVIRt
W17YI8A6C2ulZiy0CTcihFxmQEWeSCO8XP8lKQsZI3FOuhF91Yui0ZJUBb5h
ZdJQFivCFo3rUHRMTxVcXHO5ppVJKFYi1vtY2V7hs3z4yQ43u8J7zUy1erTl
lVajIExvpEj0Lri+zsGht9bO1f5AyMYNKqjm6hrSoxFjrVnZ/NJqy4P7qG18
Kp7bKum0ot3f6odbEdqJJWjEFFOr88/obo5Lue9T8FOgo0vR0rv7rPKS7cnJ
4N5+atgxSZeYFcL9aS5EuUQgm6PsS73P9o7N1Tt4Jr+TqLjl8Hyp3bGGemIb
Sk9rv7z+z58Qve6RBeQiw4P6MoxD4iXZjpQ3tHFFjpwvflxjT0YOKpco7QWE
XZne1ZGkKDsi+f+TwnAXsGOy3s3+FOI4U1CeZvJAezZaL75+P111dm0mGNEt
fFFWanPZv09Nrj5A8PNKO6Dr57YEeJZiGj6fxvrqyH+N2qS22w5WAH9S7emy
Ugkeqhvu9nvN+bxQ5ctIcKSo/U8glseGLjxuQhgs/PIK7BzwoblD2IkgPV73
1m/chlw4SVXDZI1QaRKNfRxAPyzKa8yxhXsuENht8Wp4eQqAcRvLX1XI+7kr
qfOiWbt2L0N+sCNNiT2BGtaToOT1qSacqMYqusuzaCLEaZq/ShvkX9Bd5ZUC
oiWI9S4lH/dDoLkmsrCwovgbJZ2jVbhB5zLG7KCrLR9mf+RKl4OLRFNqlNI8
M3IguwZPKTc41mzy/ZVq4uerwTKvrPdUvNSOozhbQ9GUMy4v6liOAcS9wFhm
aUkc7Im6mJhWtu6KC/T3RSP74+1Xkr4DUGNp5kCaZD26CbIS0/sUsZ/ilPAe
IzBH1+vqFf95GpNDzJOwfGf/qY8Gfl67f34u16EPhF6EtBXxsDNhoW9XBToG
5AFslbT9UMRGAE+PVjH+X9DGAVBg9YAiXHPvtk4546jlOOrIM3Sa+4EiCYuc
4upXxtg9Fin8GlnYiFRqDUY9XLATHxOQMWmYkwF/io09g9i/H72/woRrldYZ
MFi2NAHb0N8efpuyU0IP+CQKonpYH7EhJq2jK65NDe9wBOYyusc1V19xpxvq
i3u+w2qCWNaaJqqTyOSFNRJJpUnrazb9rvk4gA2YxL8ZmMQyBR68joKiduP5
5cqVG4ZuBVF2atUSuP9RQ/Z/AVP3loogjXKx2AoF8lmAKB5LpMNhkl586690
tZKEOTR7WjN3PoEh9e40X0kuEKEayZ2vztmvYfFjU9VTW6HP6GR0lf4V4k1B
pxRcZxnfCAJvADE4CZ/vPbSgzlDZspc173GbTlCoq4ZjXsYh41CB13OKDPuK
ZBGjy44eCq928uV8RKo0Me3iFWst5Bl3YcLSv80W5wlVDc3PU2pVTZ/X9U/e
UVr9eG6EU4p2NGzPn3G/bS14HLSIznZXq81WPGEaezMVHLR5yF7AjrrYji+K
b9rzsGWLDoX/RPoAG1fjXzMKTQivrw92oXjnBtLEuzpxObGknpiz/Ja9trvf
co27+JCl8MnMeXPlv9xKP3xg8eLyYYOFdJ6jxD1NG7I/6bNxc+Ujy++YPEwI
bPMmPLj7k6MrpBYI8psonrVI0OVG/zZhzrFQvPSQWGJspL9L9z5aZ60Shf2B
UoM49LDnTO+Ti+mgQ03n4IoDebuEm2EQrFyDbvKN1Pvxl39o6GldeWfwaV7j
P7WVkgjqhAyJWwfI5VyIgI+WSj7cKkNFXvclzAO935kL2ylGKlGN6w7rcc+E
CJfld9YQQftT5AxEMA47qsNA4kxHoLskcqbsZW1j0F0SXFgk++qldL/6aw/4
NzhbmNGOMjZB6J/sR5AQ6d+6WB/Vwq5fxhKWCJfj82Dij8AA4nuW7Y+WjZcr
+8m+zOmzsBRkl/u0R8wJmyV3Olzd5a1PwbdiLqkAvmzc+jakIzENPxnzxgoL
SorwNhEDhrXPvdp91FM0AySrKh9UvUMOWFbiPE9jfR+d2isY+35deFtpKz1H
46zfjmjZW+cits+9KAT+O6QF8Yx7Q8gDOpJUB68Q2rB2+8M3ed6BTVUvSlGH
2eLGFWqF1Xk7dd5Qr/2neeaf2CwsBmiKekgXsnCoThGOgFoRIA5ciSLNOtwR
LX1RsklSz8++YKAjcEtrmBrxRg6ewWcLM2+wG2LQz0cimNzRNSmzmlJlOaZA
14XmVwZ/6o2A+X2GSxsuABBsXv7yydr7HEv4NVhoGPJ9FM/OZ3qIlLb7wi/P
lWflqQ3tK7XX3yMybgYnvTK9yjSoXR1WvlhrpHRCo0bitD2tpVlCIlNfFUXE
GGqibmkEHTZ9YmwrQdmZGOlLC0GepMP0QKAacdLiRa+2mkDzt+7tLp7vXerO
7cP+fsmtrmlY8ZcpjZCgAuHQ5A/ZocLeTwBIrmAvt3egZJisX1OAOQpIUWhv
+Sjhw72fuTmOpux978jB9XAlUhnuXsfw1/+M7UhiLjzMAMgLzQH80CRk4NB9
Jck7rU+czBusBvcxnMUXfh+eaKpN8svYcpoGBVYb4cHaR10X82waZEy/3ikc
afZvwhT30tB+Xq49Zrd4WysFbQXmSIWdn5F7b1i3eRQ2JNQsJGJdJ+/SMyAA
8Nw4BzTUZMyxPrJCIovz1RHqBKQ9wz84H/4Np3qneclIectV6eE4tZygJHpY
R1Yp2rrIPrFzRmxciyfJ1yJc2oVSPbavNUN9dRW8mppSGQ280oa/5CnXjcKi
nUYtzBY2cOydGEZbLjKIz3XhUGyvgGH9mT3vAZriD+IKPWkZ6yCfqYp58rFR
z9ii0oIkucIkb6fJWjgfIwTAhk2irPQtUMeiQECldgPxiK8PhdcrqO7tvVEZ
Wb7zOCMepFvuFKwUUakCJ0tqC7Z5MkPmMVUMbcINBFXdkfP65gNjcJKb+Ahw
d3ptqaqFPqbDEJcxd/X+rG0c5pc9RXMfcNCIXyg7g4Own8pq5GFtAhafDtQI
VDxI6BBxrc62NnFOffe4ZzC5cSNdPFsKv0me578aBi3hVABZYh+BvsiXh8lt
+ckxi62VdU4VJqhK+T6jhzlBUBWFD9e1YEnBtSY0kaJSM1dKaSYIzT+Vo9K0
dEn7P8T7jbnO+5EH25hMIR+obOsIff6WMvzmAn8Z/HcQJ6oCGMVVXnCQZRlX
eRaOFQXlTEnwaRhDYFh+GEG56lDasRQOatO6zVC4Ziw9owqILOj1vAsHA9dx
kJyQyYp2wRl9X+Msjqa061UQ09cf5PTAY8qGTiiiguca/w6S8Umd6l6ij94o
BrTpzjrD1WnJZ75+nhlRwCM93F8qYeqiSom+eZ94iPfA2qg3J7LaAE6BT/ga
ZyB0bEFXhM1uCfUrAXOMQDt4JIFBuVKxyLjeVT61q2FQ7qhoGWDGl0V9ofuu
0bmcw8dzvv6N3hollG/piucGtudTkOMfdYDlmOK0PwM2xr3plBvfkjtfYZ2g
31tyWnHB3Fwg+YNZ3gbFLWoEgPR8y+256hLZfTBoV2SZyU+lwWXXKRypn69m
fiwFb2NUMz4uJVP9Y68X0Tekoa5y1n58Lvft9VVUAQCBSEqh2RcSRW5aByzs
NTNsyj3vbEalYIlQToytIMgeKqaEi3InbsCy5R8b7vNzoBvLBcBKyogBJ02A
mWnHwD6ebMp/9OGNiYUsvZzhW5zjl3x4vF8VmeQE1HhT5+0q5vFbcyvpDLu8
09QNazExteTOw1VIiiKlvwx3/gdrADbR6afSOvkQX/M9WoJ62qQIilP8Uj6b
ONPmcekc3L9HqM5oA1jafJmT3/sixYru/ykKXPuuIgPp3uY8+lBB9Y2Vc5yk
uIHA/ZmJ7a8hBqMm4CdF3piizaRfgjn4vRIv66S292Tgxa68DT23UoMdZ429
DrPW5Z1UlSd8h6GXaB9x2yTopihZZs+Rola4ltVXojiqsq3R3mJEmfprQ53A
8o/03BXHkRYl8FFFo3FiUrQRK6T2V46YU5RUrHbTFg9yLVkPmyaVbFGhPo4o
Bw3LlMNYcVlvbevYvFMeasaPprW+kaPNvIsX27ET9reVfQnvIc5zsClIFZFS
BPucIx/LVWdz3bqATtQtPq0i+eFPnfS1mRElq0VF8phLpmcSWkAWRQxrHYxl
8Qu4kBF/oYQIQtcC7vHIwQ/WE2T3zBXYCjLWo5MlTZDN8mCHhEQP3SMo2PLM
Hf1BEKKHPwo+o1D6LLfGrjh8uogQ7yIYKWTTIYNvaHn1j4fUxLM5BINjIzAX
S4BiVF7p0WtxJpaPrOOpLQwhzDfZ5SBV3DR54RloCW29zRXiAy92KQS88fOo
ZtAWHgmaksrOJM4oDLFaMFflhFLjeyDZIs3tVgUVbZnI7uqqN0q/W3JayYjy
g7ZMb8IBt83/ZD6nFIOPknG3sYe3153OJreHC0D+xhRpnsICu+TT6Z+F6iXv
wAgLXGEPkprevoS/iECRmLjjmxfPpl+hJl3zHw0h8BA71/ELCE6Bo+7ZJJSr
NZcYstKipuIYa8QcqCn9+t7hvVJAS/arEnpI4o3aESw5q78NuX7G8rBKXr2H
cu51gOJD7JsNjmUOwXoV1TJ5JK8jhyJyvsaPQEjr1p9z81VTv3QSkaItyJ/s
8/J6a4Dx/NeZM4FBwfoN0oOxIUFYkzio8wD/X0SS66QellHHoGp+StLAv1aM
hqVkhQ/ejP4RSSDToRzmayhs1iz65YlnqnLj8nX7RV7ZZPZBMRZA0tG8u75Y
B/qK5b1S8QD/yEa+FMDiFOcx7NBlGH1c6n3B3Bw1luRGxrBLTbNl+B2wU9PF
i5kS2M4LIB6f1qidQ6PKzD0p0fd2MtUow5Q5Ue/tSkN7IG/X1r5ErVQxq5uS
kBgQIwNgWn6gQDbg7aYbAMdzDGFNMl5Ph2e7/SzWpGEXKmpnSIe1NZDXPzAR
8XGA7p7MpPiuncHQPDurFyCYRPjm9Nlix0O5x/1USGb+n9TTEnVZPWhhuU49
A8M97mOZ8MV9Jl2DcIKRC4Qhr5qQAVBQZtZjPMm0F/IGxvAxgXatKF+c0obk
i1+O1iW9tHqcHStZoLhpkq+HUbrjiaRLokqgiM4QXVu9A6PzSn7HR4aNvaqm
Zay6aCx2roPhIxsz4+H8mQcT8Yy1+TtbWdN81/hZ91HnGLhggAeA7gdGxQH3
oKY1QGHBCrshQYqlFWm8cOU03VOD4TXOBAO4INcutZ4noYvdRe85ubivA0BV
II0mYl9doCDqbvoJ5Kub1oeZSOqIVIp8icsXAsYxlbeW54Ni+++TdwWfRpGi
FIWsmWvbX4uSk/UCTqxJQJNpwlTf84m6ZKQCoLL8KB3sNfNWibVrseFz2SUe
5+dPmoCq6RVxL9YXz6fn+MiZJ+fcyG7qGHR2oH28lsnoAGOsWjByj6LujDIw
Uu8fEo5WO0KcQ17N5aCdekpRFQ1lhqsunQJz5qliRofJk5xuW3UlZYFdQEZI
FsYhTLZ7WqTM4JdDt33bqwr4sRwXZ2eQC79ngJ8kMf74nNV9akxe8eCpR8gd
6OvQ50QxP/rHSNUxk0CuuVCpbIJ0dNQJrjvadsZb1NZMrrqgzagRgHL7ryMU
bRwDz1BWAQmMo/bJnZP3BM+VUyLqCFtfGwZKr2uQSp4jsIKXSSxA01dx1hFJ
6GEDRlzv8VyIRFjdtif4TwQkVJeyExD9lqk+E2yTwq9iBBWHbSDlfblxEvTu
qy+5l8vgNTpezEUCve2Fsr5TP+wWCvpFE2o6o+oVrukSZ7BSTAuOHAEhGBtk
B55wEZ/zAlGkSM1Cm66p9qsNhZQBctHaSjlbG5pGV/k28/jYNzWATdsV+b69
0XigldqbV3lwzHJT25CcBH3Csi8Ry2QxIvqKUJ/N1mygJZqfoSIF8PV+5tGr
95jBU0+jFGVpsj7Q22szVQLmZcPPm0YFtCFehaQRpeFXWWKTOgBh7FG4VTPF
1OJjMPYC1sbGyXmVA/G2edRD4Tls0Y8zU5HcvubGuKAz5Sz8kwEHMudlR8+s
abJB1Db84Dy/FGq3yIfzZ6jTfJ2Jh46S7fpGcnseNm3+cxVmYQnwwGdsVTkf
WmTngnkPYNwySzaJPBIsBy/aaglSSztWM1yfXgUxQvOMxGYoqoYxJ4YJjG+r
DlfDI2b4/Uulthz0xSK1xdx/J5tHJGjtOVrEYNkZzuvYlHRhDnF+3CEtot3S
VLttT1kuRvdysv5iKuprCmP3FJa/ydrTA+7YslENJXI1Zgxsc4XpKaBPS5Ey
SmUK5hWN2BsNdDrVjtugN5VthkWsuRv3/0TD/D6q2N+vKniKLdMiLr7zE4h+
R89Jv7M//RVl13Cm9A6Pr5ynL1s2W8yjlz/5xsxiLVkZU/wRYxqKvLeiCNNN
AwYQR3pr9MXkUuE8mDEAQXKYUepqLte1l7DLaFYSnsm26zJCuNEY6ZH7kPPt
DticYe1+f8knTNUxZGWBs4nuqaVy4y194eDIJgu0BjnTsRWuTZ46eQRgFeJv
OMufBDxFDCEeG1hB77O4FCaswIhhJY4tB+BFxgaqEkt08Ty4wh9y8z0eIX7+
jw7vvxa07OPhPh0r/D79aSRIbD74GgV/RI7DZr+CUrHBRwTUjrEi9X8firpr
uTTBIvR0qLSMvLp8JZCdGRBv+JgYBgOTF+kv5ylJwehj7qPFPsnZ7At/QIk0
Ig+m8bO6tH4/Cy9c7te6q0SWwhqDvrPuMwNK0ObWHrSV7dJIEBX1fYYzLP/o
fCr77YWBCILbH7+IbA7tzzkhucENj3pEgWWrqvwIGmObCCiw3HsYCyieTGrM
ZgcFIatxRcl3knLhimjM3aZg+qD1WcoquatyuIxP5ZBxU84DoTxGWFihB/H7
18TEYTbKeF60aofj67x0isJmVmS0MW8y0mUT+At/qaOJCYmGQ1W8vVpAObzZ
wJRUJZAE+XBOxnBTwaUbmYm8bFRjDrNFraTNe1GBEm9nltbunkkpBBeLhN+C
sfo78zdIYp0lyUXm25PH7Qf3oUHjrNDIUjX+Ye8dl8I01UoNp2O/ZSvvkHCu
TWvfT2xXzlAi5qZT0SSXsLwB4yMpj0SBEtolWI/s7iOmY0kjhTP9voA7zHuZ
895SEBE3ygpLmjtLhvk+Iu3sisZqFEytitmPZ8e3j3I53EkPTzv1nIbCJyyr
BUyEbQpZ7fuJzbQXZ/7cMbZ/YtqtId6dz6kgZ8jaYVumLpAnhcKdL7cERbUf
lJyBfw5nfHUIwlldhK2wmZ/s3bxuGhnLBkwihRkMpxjBmO4gcQCTU+VVlzNZ
Thq7m+kU0/4iDm4SrpHkYYurQDsUP+ZrpKO5BjplwOu2gqKDDhKDoaIKR5VI
rdNqZAnAINsOC6MxtLSlcbw+F8M6OTTncbWpZTz1+oNu4Qy1jMCFxzGs7qEn
eW23jOqibZNy2UshReQEU2fD6liz6mkU9EXBG/wX80tNldjoiC59bWPqHBFb
xRtDooDHCfIXaa/ioc2DnDsczb14SAmvrvBIYTuYEvUXhQMbsyvs8NvS816k
u6LZlBZ9mPFcuAicHQLHbvpSDTwM1qkjXBOsPMxV8Y+knqdmSCoqkSIgbtIW
UtivoH7NP5IsosrmV/oocMbSGV0Oc8RSokgrhWysk6yzVueWDlJwURx2/DYm
w/lk+OgZp0iszrQfAD3kDuX9qXgJNiUwzrHyl3aRMHUz1wlMPXLYWPuNVX5L
RwuEQltHnWTsRAxjo+A7SsjuWQtWOONiWz/iq0hcguYlF9IYHyU4KbHQU8Dy
RQlshBGE4hmkkgYabZJQAOjhAoC5+PpUoAZ7phc0mDc+HVyJ7bFFe0E9m/PK
ieS40fFHIWT94hOWVuITcPC1/gJJumDAFkjoWDafnh762adOlk3VIMr1xVIi
EstcEzSzeSvE4yGnnITec0K0NEacn+TjMUfnX5YIvUma6VvDzbHodMKdsYPW
1WnDMfNU/U3bMn1wspR0iHey20jfgm9sanS3ltR8nSaOXPPsa78/rs47cPtQ
s4ZQc0uwV4aQVsFLuIE6rM9RIjoC4dOg6dKveLNODIaXpdsitt1hqgSQgXqd
RPUZzTUKf0DrlVM4ydBLEnUi9v0wvqREU8hNcDbf+beFk3LHCgyWGC6A8nzr
SPiB4pzaZqtw7c9B1DNQ15CF3snCxF/qcCP/NQBixk7/jNY6J7iC4xZ0nvT0
oO8ot/qHw4tIQYcs/CvnthM7KEWYLxxbsEEG8DpfIXVnl3Y3Nynmd3jHMKfF
r4fokZwxZuJq+HWlyAuRGZO21TYCmlZZXh3rvVHKOvA4ThzfqXV3DkC1UHwJ
ZTyZOie5KowhQex9jNOIpgt7ELAVnvdPGmKucRKeQ9mYEIN1RkIcRp8TGFnU
TWQ68stxGKYO8Tzte0TTBuNJfFuaiviA9syFPCaaUGbG59ScOSrg6klbEcYD
GVhrFg4exD0pgu3eNNQiIKGZov8XRjNACs0ObOS31qRKiDk9c6XZafDjkfE8
VaYSykYyFeAFxVOxqdvGdu02yaw1czkhTvthPhZ3mqEhcexxW6ZE/dQQZEFi
egSHAo1+h46olO/3Dgu4VQJh3jWxU7J/5iGV21M3QN6oShTk/oYu8VinTFQQ
PD3q0B/9mWgo5XhBNergKGNkVaYETgbBOcILf2S4NxQKq3tFc0d6ax3MATQ9
LHiZpeX6v5TyeSfMGNs1LbaHRpI9JobPrOeO0M0iWl82xNwQjV6pAndCg2/P
2cfm3Wy7ZwTppHcOtG7P7WUnRgQzTRLEi3dOPNnXsctgU/5qjmoB8/+8C+Dk
jLAcpjk6ccAFQY4qIlOq3i0N3V+Sf7HobFhs5YcS094hYa7UbV4rf3H8eqU7
8ubCssDaDV/pb3787qg/R3CtCnwQYeaEU89j9ym0WC8koJYPwgbaSJpXHg48
bs1gx9nFml0RSuvk881pEnYQr8eQc6eMFpxYegOFLrn10f5g7OxiOx5OAAQn
2O8rUpf+wHPt07EQZxs0B/t9fhcSH7OUReDLTs8vgmWCY1iteSTArQ1w0FTU
ao/4PeiPM/1Mw4ADbaVdXGr7vfCaOfKYYIegPp47FWki/9sdZYhcgZ1xbYcm
9nFzWdA5SEtuNImaRUWTbb17xn/Wnr2Z6Q+VFwrJ/+PGkqn52BHwYrvhSjRv
LmSncxUs51MuswvloVyVr3wtb2/zlG3JDPScVsfTInwGGTW0RYnpWWr98JBL
uMG3QxUFDDisRRMAqtrvv7Qs1ZtGtep9r6ho/0+r0T7kcWyhEVL6z/SdWevu
b/yfYWlRzPG/TO0the5qFeJv+zXKjueqT/N6mcIs2m1VAmQWwJM1VMyoqwFM
3tm46LzMuZETQXUHeCxa7HXyQtfDMmnRiYXWzPGAdzcqbfe1qvaJlmkkJBte
WI1Gtsxn1i1VIyvBKJGrpc8ieOpJaKAQa8YwGLi9Id9o+Pz+uk/qEAIF1yo8
KfApZIIUo049n8NuUQ+aPReNK58L8cr8QHNcIOZwyoiScUnbrHByZLtcvdKM
RJUdmq3jnVbeKTcZIYWowQCYZzfuGkpNCwDAcEHciRnKtNYK4QQeHPz7p346
kd1quDWjHD6eG4i3apsrMrSOjkHN1ez95DerEsfj08Z8D5x/lM1QbyI/HBRX
AdigJk3QuvJob4R0soA2/UZLzePwJ4aqeW17X0C++mjGPK/Tvx7oL8Fg/mh4
KsHOQbdql7fMK1yk9WJmpoepO0qv+H9dZwoC6J2+LC9jujKY2ElcPesuqQXN
+9fjafooWgph8rdAYFQep0GDQ0zHtFM1HPH4frHOqX1kKP4S9vsvDmpj9Alg
VgjC3h83TgRfYci+D/XGetF8h2hJoiG1Svzr4zqxU5U+uRx8FAQsMzkD7lC8
BKFByKqxCSpr6G3NLy1UV3zaG1Q1PpKfmd59bc3aJ9477QKlFAGnByxS6XX9
cEykbSYhPiy30Wnq4+/wvYK8h3P+PZiBzXO5y6CaiI3aDv+MZGWzYNP+1BFC
GgRyVAqZyMq7sMc+dFfXCSGVQVp30Qtl15lny1CbVGzjqQGFzWge5owLIClk
1w/VlBWttH3Hya2061SYqHEkMAeFIS/49Ro6uBHG4gi/FttD9VCNIBtTY2uJ
1oVtuKA0xb1tELZNcgVbencd8nf8t4RgAeVLDN0vjY2uLkHNXYpK0lEIMA/c
O98w0Y9CO26HCySURdvFx4uj3dZT4bHRi9BGkzssbMyroNDrTifVLdFkHYeu
3s3dnEUPYJSW67OPnNo2F0pidNsLvcsecsXbiJqMzmovdxnmtxAP/oTBfDV/
FYqlAZp+WnC2ZTIdri+n4QO+RxaPqftDOJ4yCaBU7rgJlH3uNdHMB2j0vMzB
KvcmjVrpbyfaI0O9R9Tq3oL+xOAi98mNs4XwvJPYNNSCQ70ohErmk7jWQHD6
tIrezx4S5L9X6zoXKF5dd9XzyEbaOpTY6lIh24WFaPL01EF6vCCGkgskacsG
MwQSrAqBQzHdytMmLkrkem5drUysxNboplLmhhwqg+eZk/FnS8YYR+4oumdE
L+CEKC+4vKxep2A7DBb1wargFraZP9SAz0Jos5+BF4nnANtXeorIo5re0DKv
vyI+yro9SOtLr447KLBxEjlllF1SvCHnZ6e5zmRLrynElCdDUIX/x5XmkiIL
+izLcim3wc2nR7ZNi3sGshZP9Wsbu/OEPCMbSrfJOso9oLS7SgzsO5PyJbNY
wl02GWQxoNfu0ECea/pyPXalT0ccEydyBKb9MK8sPBjntVqJjMsGuBLsPbHj
C2oNMH+vJ4Q9DWUPOVAxYKUIe3aYu2SB/MZLNM737XScMJYW1OkZr0g6SURq
R5/QpI0rtW306xdxcuybzrkXUvfWd1Zmlmsu1K+P0oKJYmvOyvH5GUkVdWds
WGrKZ12LZc2kxoULVEjZAoFbm+TnSCloCQn/PR0FW2xxTRJsgpA39cE1u82H
UOxn/+d4OEVGdqCFSxRS2GpaxrrWfFtxSyV92hdunG/AsC/x+MV/SbkxAzBc
cK7iiVHLfb4BtnaE3Pd8BLnOCU4R2w3CNztmO/PmuWWORE/uEyhjGXrTRUoj
sxlWSAC9ITDFImiRCAh1PkZ0TBS55wFnc3jdDKSOEPZkwU3Ng592mg22uB1I
zGB4fZa1VFbK07jsTzahufK7wm+7DZ21sIOdAqLs7CPQD2c8agvpnYQkIK0C
Bq1HdE0BeXf+tbkk/v8NSjCWfcts0ZqfhXMIaHRQCazXGP5+9oBSEWyLaE+i
oYBQ39DMW64ndTgQNwIdrDLDDq47RSRSH3HEVisrrQCIr2MRHd45HTaunYh5
bbodO4Ru+7WIWSl1Y38zcNPHJTFIaLXbEWOwEQCmsMhZrj9HrTTJMLEcW8Xd
xVsW+7V9NWpO96L4hngCLN7MDrh5Cpe7PqZGb4SM74RSy2c4i74uhdf6uNDf
7F1Xw0ZEZBE/w2TBQxc+HdFB77C9gHAmD3ThWzYLj1R9WeJJ+qEiWEX+rPDd
8PTYuhQ51G2eLR6ubCGGGbEE5mhDr3L/4J8dV7VT8EFMSGjORtHyai6UwrUC
ApnJ/Lsyovkin1faAHveaoMUW5KRWQZSTqKwTIAVBhxdFDzGNAbcLKhM2veT
sxaX2MorCrjzZwOkodtv2FzAtrsUsZCAkln0Ojx8GXXilrLA0n6yxFRK7Pqr
UlHBaJjSr4oRR2AYWit+jpY4MS3YVF/G2Tn+PCIx4J25ciDFg1lDMnS7dFDZ
Wv9DftVk3PksGSz7RpEVxOPpuGDPzRfFZgB6WazOB4Qs1vqRZy20sD3F5yP3
aNUALpvlmvvqiEcXEpZWquZNQvCgQoko3mG4HQuDy+nGk897I5klLp3leGsK
G6LuPWnjGecjua22umt3BsW7LOu1njASOwV1mwIv1zeNclDGK274poncowJJ
4GgQ1PJHf/64p2q2MCPRy9hUKQ20tzy+QVtKjU1o+MFlWOSt5FLn9sNOUClp
nsHZsyGiojefmx5aHjEpcIb8AbkJiJUhrklXp4YHX86f/Ol/G5gNyqLocRUa
2rK/UQkOQzfO8rOZUXn0Bka8K1bnbPftAqZ4fnPhrguUqhUrOwrIo2WcnAYn
tyAFbNUSZl6KgOhdyBR43w4h7e8jI+NJi/X8YE3HXT0tKtm6sOhtlGtIyoEz
RGGrAcau2p6ayc5hfp7A2Uxdr+fSbOWt2uLTbmuNYZa14x7J+sngpYjqzyQl
npJEwc9Udq6bFD4QpwXlqvsm3C51gbXMfJTkyxYbbqLuweW3vaDjjESgCEqV
Xa2wt82/t8JuIxGj4o3LSx3Qx/AZr2OvDUjoJjN6I/2nB9vJr7npinFYgVhU
oq4cXXl7s1zhLMGipYrqGm0nKkOUCcmMvDhxYUBT2na2FHi+fm9VALJZU46/
hhvAzrjpIlvel1Z9/7dq5cRpNODeqhgrwTyRDjfFJRL54gQHVIg14tcZkcLv
b9MoqmXFurTWEK6QteTKRoA6Lj9LZQSsTjr02IEcRJfAIs3ID2OZuRmBUFKs
Mr5LoLYqHP1uOdbmaIiXFLIwTIPLsMRSjrSv1W1Zc/299dE8J9mUSwL5Kqrg
yshNNSh3V/bCUBH77A4fonnBhEKmECASV8UZy27pU8J7PC/OClaeAKzd67Pb
us7Gjq3648eKQbLR0iH2hEId9Xzlpc8hmJF59l9d02kcGpkrv0Zz3f1y55xS
06SoCGJLVC1IvJ8ESFKoyWJg7GFRFr5ScTHTwSI/UHe6B/B3VEpeMz6Wf9z+
u/VY1ozFhsaOYktzyAFUWZLm1+xVl4EH0TBNfPrj+OxirYIrxd039hMR3ARf
RHzpEamJPQ0ddcXVbwV5k/a7+W+1yBkmh6KbXV6GasZyvSl6jwbrf1eSenuH
3ZB6D9FN+h2P+G5NHNTt3yMyYpY3yf2q88TEuPrxr8/f4nJcJMQX4+ckFF+4
RFXIjQaJslbIuSKj4ieKX3l+8KFg4hk69THL6k5XaNjIkmQLBDDBxrmD8sQ/
vd1tE575HZHEFmxduUh5hdh1gL6CsYyIyqGp6gkantW+pzY7VBWILPInMbU/
SDCr8wFaXcIG3EOGywoImw9PvtuVGdBUnfNPnUPyOpYgf/FlqRsgo4Z8qCMH
moJA6LhmB3rV/gA0gitxKsiHGKyXMPqZa+WEbElQ8BJ/+7NA3cm4kwQYLTUO
YQUjjmUu1XQqSGEfeSdBO6N7+I0SLdhE1N0iHqkHqofsyC+lAd5cdg763lG7
iYZPIg42X0Kr5wNLWhw8UK5jmKmZIedC8+4HfAr9caVmNVPj6dymNWBRgYRU
/orVRzzfn/NEsROeBhS/gWC6meGjRMtQmtCgflsDmT3SnB4D4Za95CizHgk0
ZN/mBONcxli/5qyEJGyGaeHfA5KH0WWbu4Qa9Fhxy6DZAGfwQ2wf6SqEeFiQ
DsDDkLCeMDh3iNkfI6Ce9KSERRnsUVaBqofXcvQx8gWIFm3z73HO0pojj8QJ
16AtiNOVMXsGzS7EtUPkyG5vF9d8d6CrSc9LrY8hzwjtw/r7/4nVoJWe6jrS
n4QOVAuTZToW8fVqvJk8fQWnylOB3K9NajwjyRB0HmolM3d6HfoX4gT0loBu
d1aohTuDlBmDxNV9XBCd+pjw6N37bsd/8T3wgWpxG9HZ9nnmcMaBOsWzvSww
0hH7CKNNwFlUj2+DGnOWAjjQhEf5AUDQ5YfTMHRZUHj+dln/dgARr43aiSr+
Ghzs6v6ZB0sBfV+PpdOXgJBYTHiVOImGY03lpHFIKyK6Ikq5I3DdMC8WeCr1
1i9q4uXGfqJn2loDEWJ4KiC2kfclJ15DVwhmhgbpFUiO9iQntLtF10VnUjp9
r5DVortOp63mQa1823d63dgzntHbOrbaNpNGcQpBceRGEKCyfgulQjedmvPz
4rJpH9omJvxJJNlETokPzS+xvBF7ST/MVeawrLQ+y5weL1yUeivgD804TVj2
Nfstzp3ibSlviN00JPN2xyhVVO+BIuuDnJvzvTU977YDWhUKZt23zsDP/RyN
zhqnVnSYAWP71KpNkzLSJ6DUQTSd8y7cWGVNCfrenWjYxrxJvCbeicvmtNhY
/xs7qo7hgKtSbTqjBm2I9KedbmQTSR0Qhlv4ZEc5cdGumEE+mEy9MFhKhWok
vNnSNOLAuh2FyETwweR6NLCv5lz0mJwIQny4GuEoRDWy8crsnab+jr4H4htK
kGtMSjlgJMxEVO03gwzmIq9eTLNu+xbdau+awampBaTvy5eBEBZxR2DC0pHD
GlhCucz3dmkEK/bKXL9PbXaQky5AJ005DGClKoHmgHaLaAKkKBnulPk+Coqo
2MK05762SSI5ybZnbNt++omqlu0CbciNXWDlxp3EQUTTEYs3qRT5EFuuldFp
BXotXJVftCO0UvuV9gvqzysCeINUQfV8rdB2kOX9BQFTUsCWMvouy9D8gU6y
ya0mOqRGW5NgkfVF3xBqDDkkjP2tIXYcaB2XBJnXq1eDO+i0hkOi0st2bNmr
T4oMt5krGwkFe7rIkBX3Kucr19sBQ1WdUpvgMJbHv6tbLfWHjjRsJWNuVr/x
TqoEUyO2PQUPYoIa5hIoG29HytQi468f0AXtzRrAR1sDfWI9OqpZO/4+rDj3
chrg232X9BuYKasO+b82KrkHwOVISIofly3S7MI80JX3rvLEyCuNpk5jJOAb
DgWaj0AIyKtiToeqYNQHPJQEKp/GrzzfLWwCtti5TQpKioBJueaQfnn9Vquc
Tj4y9HZhsLY7IF6Mo8mDQL/96mrImvJNOEfU5Mjd+Qf3+T8SWqxgSqD0vsE9
e6aLWEyMRQpI+be//G4Dc8sOhWeM4zZo448Wmmg2NylMMv6hZKfJot7paPcl
61N5h8Uut0eBPQ1NljdjnYq3RLxypOcfZm0s3UxPiOBxFyaSm3nzPOpQZwoT
Wpddn/zu/lv8M3chmmJG3+niGUjzQ1Y5B05eX0TYAGDz5VWEm82FyIzyXagg
d8QnFUNOzYF6IwHtTa7vRxkFTeY9dE+dIWhxycfdHDt90zHvsf4HdibxUaQc
9CqiMnfzRMlGjOPrVolNjORFeXq5H0P9CRX/Ay1YX5+n1HaRcoKloO+p6EQ7
ZQE5jhEviw2QgOP7f2tN/uIgcnqbXYezF9/NBhTq4mFHvoyGHG4qWKuBGKtl
orUFpwNnvCrsA5zo/75C8I+8zsC2QJqnkmWERO5+dWTBSpusoJBjwEkzkaT0
PEEzmuRZRPVDWIbx27fTiuvSo/9hP4b7CIrXcm5UQ2iGi4yKM/4dYJ0cvnkO
x2mswCIczPfGy42nwiNa/niiOgVnz61wE0f4cs3ZduA643Zqc7Nbzl6qrYQs
/oqYgZ8lrC6QD39ELcJWqsw/WBqiWBqVdA7Km3mcOwBmsvg3Xf+rYGoAFyhw
2W0OgPMzx8k5STh8z4U794U5P000YFetRzW1BkpSZ+/eU5IC5A3P3ghL5V5P
vg9tEa/PegpDHbNq/zowVPszLP3uUAtGlQcglCPa89IAHS6d52Gnm5RQVCB5
6G+qS1ZbMCRLIuY5TOzw+EnUKvQuhuBB9qhrl9gWKUxcHIRrklOUjgLETFHl
AVSvqPIhLd6GICohfN7Utjibyl00NaTAuwp9/6SPQmupGPt/72g7TkJ0rZxf
Kke7j3k4oh6kWioc58HIboB21dMZxLcqw8fmgIBNAZjTsG889t8otaNLk80+
Ka7ogz5fR2ybKr46QAm055YNslMLWq9ang6LJ6QMaTX6W4KjcqNoHUb0LUDJ
hryjNcd8eoVSB6bMA53nafCbvMs18Kx2YnlzvbcHLqJY86Ug1BGDMbVyRSR0
RQzw+QE089l0QSECbz/0djomZ+9fFMIbyCsi1q+FKIyEgfIM02Ifr5FPrkcJ
cdfoLUyOYMXdw+BgywHP0tAbVNn7Ajf5LKwN0mWAoEMl2HTkjA/xCGUi2YxE
JpCccL726MfLavpU3mpW5X/3VGjog3ewg0FZcNPcb7KECTKV9f0HZ8WKu6xP
p/R515cwdO2D7BXijLZGKk8S3qFjUTrC9F/esGoW7ENWonlPnAWCXENvjorg
yLP+TQ1g89mZ7YJFr6YHfzW0ywx8zP+seUGWikC+kyd9gBpD/i808Oq59Emi
vO3RSNKoVFEnqE59i4Jdh5b2uPj2LxR2Fj7mZRcu0HVSooxKuQ0PTK6sBQAk
yqiBudhiP9ENj9RHIkLMkf3oub1aLN/4uPtCOxSkm3wGSFY4Szf3e7R2nON1
eN9qFbedgRy24Dq5R62l4HxNeJ1NHad7eoSTvcpmDgpvWxbVeJEkjoVhWJCT
Cg25jHJUDLsySANCcHRRzRKmqcB/+np3B8idAyRLX7B7MmMpTNEsvdBMfPd2
J7pm6j+trUcQ+N8fUKzindyIDjYuXpCn2aEtDfJHDEB5nf9VBg1kPlpgSxx1
wfZXNxYiugnh4NXYelozYmQmR8ux1vEMdKM4EWLUY4TrNPRDD/0E20IbYfEQ
EYaMbc1jhU0axonkpQBCR5yP2kXFGKxZ1YSZK4KN4XOXby3uU8zVe52MbCQG
Orn51BJINhyNBqYktWBcHJTJaqzXm6LcZa4gClLitIrRKku7sKHqQt6AZ33Q
1i/S5FaeIBj7fd4XnVnimq/ti/0dNH/tEgV01oka66xtv8b4hj1L7MSFUGcB
+jHSDPhgknbNgsTO6JvdHfAiGiVsrpOC5lFGDvsUMqvw52Wb7Y0dhpi7OWoO
jBUNx2qcMle2iwbfoF1vUkEXToNB6iivoLp1mReFj4KTO2gW+oh1NvolFksD
SXoC7azb+Qdm3EVdhsKWToJm/Fz70jG6mOmV8RaBEpoCm9ynoQJKqM0OnlQF
/3hqJUKP6raQvB6LAGmB3/R8rNuvTjFUlxj/JemAKtftvmuLQQriD8iAgTLg
fh3d0aH5i5DQ2iItxaFBQu0NgAOu7VhCxmil02diLMTYVmT3H+XSYvaAdIAg
2rik9iVNd0PE4DNu3E9AZeCeteZ74KGu/ZRr3PWfowe9PfpGNy9jOgZE+qtk
FWOF3yIVZtn5QU8fVTxmJqVhAaBIoW9A5eBHKimCaTIzZyIt4fns/oCHdq5b
WEjQpVond58zQ2iFS5TZcuIFDF8Dj/dPmmz3emn7qYdhzfVMEEKOd/OUL9M0
1bVmKb/nvazyc6EkGlWcvNvccVeM6Tyeivtcttowg/DmlvbJWIOs13vC/3D6
dT7lI1OM98JP45Gc/kgnx1jMlS9jDAu2v29kE3BClyf98yif567Tl26GDoVq
1z9CrZkxJQnEX9etTfePsajoY21nnzP1NhalpJ+0GdqLrGRUzixwJxe2gUra
h2fGBzT3ncNaGmTyJpTRy0dxn07fpJ8TsbkXXwoqf7t69xMPF8d6afWB19dg
dr+lju/kxoTX4Z/U7BudmrA8kLkldJngiVoWzUjyZ0xpKeOfZ923P15TgF6N
OxNoav6xRkvpDS86h4nkmpNSIBNHTJ/TVkVTTvgurGTlUzx53gg0h4NSFc8o
UjRBwPT+U4IP2DpCdKN1jPbLx4Vnn8Ks2Pkr/XOXX5PCHeHDSb7qy+a1APuj
Kx2Ktkl1lbAHEvklLO3g/YZezuyhEGj5ZvyadQ3L3cQVt/qTs63Na//8/GqA
sSnihoXLEca3SPJi+4hLInJqLwRbBC45nIpin+c6AYE1t8efgWoz5zyX4CeV
ZOeVRAysyglaoKwE2MVa+Rj2CY+emJHNh8/Tuwr+gVmhCrFl0/f7A5XyaOJ8
8ykwFX6MQzgHULVvJzlzY4tkxULIhTTy1GjDBupNfja6hbyx1Pra2tvz9MHW
A4kXWJM9PD13Hn6XErmZgczFYqS/4HdxfZLFwI6e9mm+1mo7B6+/Z2L68PxM
s+nsujCmx3KUzP0oKtTnC54C7agAfjrvgH8BpGEl14xbs4nS/KRFEM7FQcoS
UYehRCaYgM68XDsYfOpxc1bw7BqwN6uqPdG14hJxXoCQ9b4ZKUAMWs9FrZjX
oyLtqaoEliSVoZTgCEHrE34XcZHPaMkEmD/rO+UzIpBCCmWUVdXU8N8R9Gff
kq/OtCB2d36vkgCGXv+WjU6xufRSzM0ezMFW6AVHfAZrBjD/9uEvyD+66wAu
MMW+g+c/1GbFvgQ3sDIM2RG9vBLDeCMVeT3IznuskhSv4zWvAVO9MvKrqsuv
OQ5bNGs6+wNBoue/+ogXOWM4q+nK0GpAQmCEmqkf3ko85dlEDACD8Q/7ByPm
r1WjoAvALdbnmc2Bl4ESBpjZU3wSXxw3D99Lx9iaZ+G5+csDbgV/A9gMmrSz
o8E+6KvDSUilrp6k8hPtVKcwZPMPNcdNr3zdSAKfwm9v4VXios42s6JcPp2J
ZntmLnm5Y9M1Z2avAgblLMwmfTbBD8qycF8rkAPvPsceRQHamrZbWcbTKYOX
/FR8eS/zW0WN4juaAC19zpeupuG+3B/JC1blTbQLUb0ks6zptIVFDJ1VW2Iq
5u/028b/XOppweL575fC1YAN/mnysIwJri9kcq0bKB8w69F6BmL8rEn2fTcl
5wf9F7RkV07YuOkG11o35thku24khZ1Oc1YeCs9aglzJAuYGYM4E4MUA/eps
Ukgrz5jl8h5R12iUX3tnghtQINFk9liyd3JU3ZY/5orl06qMzfsQdndpDVNG
s49XAV/KyhkxMOg7UN+ruTprBPdjJpatE+FQlsKrvbYeZN+m+HYQ3YlPr+1I
/QJFq6dwT9O0sr/zo3LX/bhQVcWF3Ass99i0NPMAlLew3WT4EqRWA4OrxDLm
poJ2wCGTLNuqXAozyB5R89eMd1o8JvBE5jEQqBJfmPNixaXOj8i7ZKbDHPKJ
1I5fNdXA7GRP81m52C3GtdWALvRXPzFkAxVLvQzBzc8lI7tKuX573mQUju28
qXpNOdYcPwYBJ5qZgbsVqVYlDKCXhiAjNLvA6sI/tdkaKC2vGqCzCtCV+rx0
kQqMnhYUd9t3NOiVpt1oUbsoq9sifF7jKmd/772CRkYVW3Y6cOvvgzuT++R7
k+u4f2lsFIOvC0OWOrYnjHx5kS3MMHwNXhdcEySjRAMknYLapF1+hcPX+DWC
PUPxn10r08WLsF2X9A1UCPA60ERigvaiV8rNWoQAHvXuPWaSwX/SFXSvgwl2
4syzhMqWqAzasqw1GATusjI1y5Bgt+KoYndyMdYzTqYreEvaCwfNtHU2XrHU
k8Sj+cL6vT6CNbO3IM9Cf5EcOjTVdwMPYQ4RnFCcFLVGByZ6TNb2zKHXN2a6
e6qxAYydlQqCzf7AbqAO1MQoTmKKInsvRKBRMZoM7bE8v/vZ59Bct6GIQ/BA
VNErlxo4cERo8/DeTZf20rRHEJylGTl5XCCcXtrQgo89GqMJ9ymIuz9HS1gs
wVKe5bYFHkyJq7hsF0CX/5sRqIvHE3b5OgHrd+sXk5E8toRvkdZvZelLQerB
y//ZgK3MWxcd6ZqAMAx0wLrQGxMBZh32ewz5NSLjH6PEXJpRpU/74QSwBxgk
VBe05vRcjz2hBbr+WdbG5FdeSvIm0AzHXbA73yYFxYneyz2hAxXqjb3xGU+1
4tv96o14kgq3wtvQNjkAyP6Vm+0/lRgsfLRbZPkH+BmwV4Htgp8ShoX1RzJS
MYSmtFSBZEG/8rSq413h//yJ6OVnUzq1jTuYsizcWaVx7ukg4EjN9KiFvoo1
/poI2JmFDFX+Yfpw9zOGI9owT+TaKDWOAKpP0Iz37oxb5wHY8X3450tGeNxB
xUfQuZW0t5VbH5H9sVCaTNPqaWo/6V3ENyF50Z7Y6rORnHosjsXEuB4Y9xcz
N1RorG3jiEh7LIJEY2CcSh+pUCxOCXED05ODDcRWMurhm3LyOT8CjH+a2SO/
ey2s3ggE6V5MNX5wQvVhVRU5Z+zKQkVsutZlUgPbJbDbkFjc+7I40qlKD/gZ
II+kl2swPBEGCYsXMrOWeyp9BoSkSJwkt9H0VWM2uVAosih0kI9/yTcX+Nlu
YEIY6PvpS6H6tea+5EoEHAfPOe8gSmLlOdqK4uf8WqQgRVP+DXVzJ6vcsfZf
j++mq/Yy+fPiZtN7d+SGxUBxR1CIv27Jdj4TmgiKIWAVG1r6z6cSnTah3gsF
bsoT2GtKa/lVlLRI9IpO5pNgtHPXekzwED1P8wPnD8RfVDFpvxK3dvh0C5IA
1iU+/f0y3CREA2hSwpD5FYcifPpC4EG4LpAIZICJyouyL0dFYDDFdrfLApOE
C08JsHkYN1L4JvTcZOrS+DQlm8pqUBkbFizVoLGyogS6Bfg/aZOyrcHxiEBV
TSoFSItzmzFtdopZrIoMWQDqRGvV5a/IZ6vPzQCRC7ryhrlS+Vysdf/QIBmp
Zuv/BPjgxxwWsy8G01REfxdeJa0x+yIvHV46dM56mASue/lHlbUjHTzmtznE
72KnYiKkNqJ9KsiQNtecbOUQN/Xe8CqVmUCt7J6gzkD8wwPTIXnwABcH0TFp
PGqC5Qpz6FE8XKVqFO1c8lV5+FpfbOvb9e54BCh9dVQnfBlQtdIWqA8ySd49
XEvdgEkHixmsuyqznOc7t+N/ab0g6qHzBFFMgeBmy32UwvA7BL8ZlLYZFfOj
jrbAM5zMnoekgc4WRoYwi17iGgqHrY4slmg8Sbs3TFezcPzktVr/w3E2YyoL
T57ckKA3ekw3okVknP3hipbgAzqm2aXjljg1yJZmu9/sodegZSeq8nbirFM9
deFUHfdLUrwfrvGOWmxmIJM9D+j+utR/Fe1USTRwsWNAFycXNq/RoUIDnZS0
rcMLW4KCpKfZeeKnwqghWtzj76nkwH+5L6ZdJadinjYO4GClOBXan/WA/52q
qv5TJD0pbvA0ZmBba//TrQLjnq5viFpFLGh4U9e9KLV9zXkXnMe19Y5M1hkc
by8W5YNaHmQgk6oTsLr7BJHfytCK3OmE5ubgBObC03/MzxaJqXP6POR6GrwH
PiSCDtJfM874zUv6Mff1MkTWckrMeP7W/wL+qQ6NHYkGlLhjAE7Qhe6LsXqE
TEDOylCHPYPY2gp567al2MVjcadzvwCQQA6zEBYRUXahO+TkncK/z22RLuAt
mm3uYeAxZkunZ3sbhJdrPyBLrhGFrPCVzjZqT3FNxmXtzng/RrPDz3M0Yznm
3YhEUDCZBWUrhkXxLkww2TEdlTpWvKxrh7kDR50dKLUolt9wvbkDFTrDGxmn
qvgNlThyjuiEtJQ2QNnF1qtSYSDs2+sPEsi+UouG6/8xpKTE+dSEFS+fnmpP
Mipw2ixKWNtBfyXDBXlY4WQGzkIr5dPPtVTnjRC27bV9yzt0iVj339vZRC1f
vD4yX5fswA7QIgwFqolqzdnZ4OWBCXppGAegy6vDsGOl1Epg6TQQn3E5GFT+
K1dWNHGGp32nVn44kgRlUB4CHWK1XOObSyIl/D8Ug8Hr35YSS5SGsfZ5QPU8
3ZKzrWIdmMGiX7/MUbWQnn4T5NkQEGG36MFBTaP/EW/bK4VZSlh0x2skNOi8
aLSBNqLTNZN1xQuV9N0DjqyiNTpdPn8mR/m34D1YsBVeCNpEoykSBgtp0aAp
vgU8bvx2jLnvJTkRqUlPs63jOm33NKb8mEbwQN1y3WTmO9z8BtgMsg8J/2G6
ErkZumFKMJ51GFdHK6DYGjBSFK8D5pHRe3Tp7KOxL8YYVWUr/njay5bqZcXq
gSsKMDmDUeycyliRhjGFwn1WSqUGA0KAK090Dj8VhbMVgwHhagEXwKa5GVVC
kKFPVU3fzCD0sHfqTP7abHp8AQSl3p5z9Qz+Vrtd7aNQ6t9YgrpulL4oeBEV
4Kk5OGDeAAMCUCqjuP1q91qBe9emy59Q8G4DgJFSAm3D6hMalM0wCaAHJy2k
sArqDpcvVAIjVuHp/q6YHgsMcXJz64P1RmYehQlEpFAOgPmC3De+ZjMqkF4e
6J4X/pUmwaMnx6KFA/qFEZN1eiMaALH1EX+R/m1rKWLvA7MK87oraIalq5AJ
v435q7s3TK43CdtrDDC150KA5cgeOEWNdXafFDQOU9Pb8wuihAFBCdSCzxM3
UeD7fo3QWyQ5x4HJpcueDG75+HTejjLwnH9QiszHiUkQJAn0IExhMwmnExGs
3NYXvOTNw+BbXmO16X6SlZyY79RGTyi+sqKzrNLGfwiCKEN3JEvt4yPdIKWI
hnh9Bry1xNbb98GkFLLjzn3AspXQh8eaO8gJVdNoGtC4JCxfKnkheJgPq26P
Cs5Ovk1FEv/Xofp8c+AyzmGxw6X58Qcdt2dxtzfGcm46WloPzvmOEphDjc+u
YinYUp5cGCd01bscPfX0BRvlUCT29jWFHnasmznLW85OsjMTOKqr5iwTq4PJ
5MjEn0tyxh54cIOEDRdBeepoh+dAsMFP2fHX2kw4rjPBFk7Gu7d/Pd4+L2ur
lE9tG7RuKf9zbiMLlx8z9Z59McwHdFjfBTaqORydufgjoXm5OdGa/hoqW3j9
KuXf60mSyupvs1Bj90e01HWk/CiosSsQRdzLc9fTU7gvbWGOV8MREjnIvy35
D2YsE09DkoVTi1jQyTLANltHTzcI46F/AGH/lDsQPeKqQrLRqVNIoxZQMDpn
+Qn6iZ4uKlLbvE49GqwPEVINPufIUlysRigrbciOSpyUWIYpEB21B172kXCr
YUsrJRLA54aKj1UyXKwln1qaFAU+fXJA6S0X9cezTnd24Nfi82yzoy57RG3d
MVeXx9nbQmBp+XIBMpN9T3FaHB/roW6NHKf/RfUZx1NWGsGI82/voqIJRi0R
dajzr8/Mms7HkAgcWXxVb0EeVpdA/LM3xLLZVOXxm9WM01V/TinWQ/B1m/cv
XdnbkXR529Uhj4CT/TmO/vB0YE7LvbHrAcW7zyBhJJciqYZo/Tgt1Q/TO0Xw
dsRJYPjtSH3ZbkFjiG4cqh97sxDW5cM+KmqSPiuDLFFq4lErcecxZTkPlKEx
XQKFmDNSIIqMCeZ9tCMR6SjQK6PAzkz1+pcPJ1tST6ht/fI84uKRXNojfHi4
ofbeOm+RMtm5zYuYbdWepUSj2SkV22EICvw75BJ2UQ4hNXcfVhLyWfbsNYL0
rFVQ+si0L6SeWlY4oDV1fTl3nyr/Vr+AiZMICaU6MYBcnG70rp6ukNq0CILn
dbZFmuPOA4cOg7ywNpz8MFN9mX4w9Vt8v7MNODEFc61pJOv+zEEBpWotU56D
DMXbiDeR/oxR96aMS01cKRddUBMlpW3FLmNal511T+6zEBx+5zRy78Z4FMAA
uil6dmj6Fh8S65S1Fe8CAs/l4Z6y8t3GVahb9AFb7scYcFaj+UGM+zF9fYAx
h6DVCgbQ/2634XeqICRCEx3AQVhNWySyMsT12MxBeVjfN2RFRzoEh6jaQ/G4
nXK3YvZpqJTUFP0tFK6+lBYS0O3SQezPz5obneKuDLlAr4YFpsQRj7vDokDV
alqmm5ZQEhzCOqT7q5Ex44vSZPF64NjIg2xeq+rBXifMqrIwI1ierTC1SJJA
hiVm05zWvX900xcTz51uDUiFX3hQNmO3UoW9yv19ylXiM1DP4AucYBYIAT17
PkvZEjCj5CMZPro/zlV9Pk6vlZ+yYif92adf9awiPOtfZMDnzVro65O/U+QD
Ll62ATCuDgRPC1F8aUnrRAzRQIx0DHsrlZkllIIAnn5rh+BksC1RIdn47ye6
pthYN2lAW7+j85qPZM1sW8iU7Cxs4OsYsmzz2ScTMVfQ7GCh2D60IsJ/TjQR
/SE4wONLHuGwGIdImfb5oZ2nV/KIAMKRct8xEWeApzZGaafzFc8VLS9lRCMr
7IUjKPufbI7Rbh6tqhAsCaI8qWezEN5SBYevvy1KxNsDuUIssFmSpTsYVs3I
5e3a9uBKbh9UAyBf5XzgMCjPoxV9I7eCoYXg/YL+HPAD/je3rFzffi6ZAuUR
PlWMhFgUNHpt5GkdUabpCrcMSGCaKrcGlccJdIAi/5pb3ezs0WeWbD6EZDft
hamlb7PDpZB3H25704yrA58KW1M5krkRMIqhkuzQ7LGZ1YejoFwJ50jC2B0r
S5S159s6CSXAeWOQCMWQXFQFpqS+hwJ/WtWUBK8gVY5Zr7JIIOmgnr6NTg5B
GpebKzXh3KIsME3ZAe/lReoErUelQ/PbMiYH2IZXUBtDz3R6ecakNZMttcY/
vWM1WRSV97p8LrGZ1iJ6KgVBAqnyai5Mcs/v+/h0qfUHQx0Km/8uFp85lQdI
vMUJAH/esfSN2I08z+jPy/RTy/Cl3yBXoAXN2yUSJ1wzbSKa1cBRStfjlNjc
BWz1V5FyE5u7OO4qtc7M8gVUfdJe0/26T6VNGt/GTNfnxqKPfWWFi9DBSl/i
sCXJJ9ynDLWjH4zi/Ws/Bo7dBFBgLmc5+vuowf/Dr9GXG0CzeLZskoKZ7agg
W+oWX7oSWg0GtJG8Moc8MZHdNu04qxOpdyXIj4KOG2SCrTIvwh5qACFMWICX
QGJrr2AztKPiq0KQ69DphMSqik7SN1Uh09H8FNmnaGM18tpGDY65bR5OS6ar
FvW1bW/0bBx85qp2TKeAP3b/+Leb4IqVZMVQ0bYzeV412hQVq20bBaCFGJoC
nd2qjcl4tbEKZOib46S+C9sAqtxVHa6uBHmwAPPQeMB4TAWACofTcc9Qwhkh
eYQLC43laIJbfpiVM5+XxmTJXRsiEK6jYkLpqzMNI9aCAdwFiF5J11gZOMYT
JuemDyXXrRusF/mjUhrIAg09jIY60JCxn9slqdDOKDAr+4zlpjeKqxm1heMZ
ftbk1EXv0fEmws6ES+EeAvw2UJcMN5zwIJ3/m8dJNbw8inna40oe0BqrZ6a8
EpmANk5g3/FwaUzblTNctl56CCWL1ZIlRiZWi+zqmoWQ5xSexwdcXQ662y/M
CsJGlM6u15LgNy0RyDZdRj3UdH95YqjnICCHmLAOyzoXwNlJ/dXmdZINmMg6
UXV3uSHYMGEfuPyVyP20ohd6RctZo8wt6nQmWyZpb2kWET52OI1vcEgItj8U
rNtVEfvUBBIxT3vlkPQb6bkwcymGqVl990tq0g3atreIS+Z1ypuMaqmm4/NG
pIl0QcsKSjKvEY9pVDxSe4/sUltOsIokMf5eUc5mIJMVg4lMA/WbfHxZfH5G
lBIf4TtdaBUBa4ngQLod+2Jh5nAEmE3b6EtnuRku/f8zTNp1RLhJRIAxvzZg
8FxnCeKL8K2cYgSNk+vXykoZzHgSTqHPsks1Fj2g349r0l+TWeIWXVpch7PV
ggRMQnosn0aT+6vO/L866c8wtQh+QiH1Z7bmXAYTwkpg3L5w6eooYzw6kfUG
ssEEcy5qSbEqvwUFuYLslnxqYw4CeTxKat0Fk8WV/Yvyf+ShDPxL9wSOABdY
AvPS8Welq8gjy/1HTNSFEYZSZeUnZCPug3aNjTGf8xQHbn1P+rAXdytff4yI
6MNvXTQ3v9y94j17n790c5U+oMgRqn6+uC6Atbx8WhduupGvfBms3xuIFPXS
jdb//LYIvhit1kzrXwV6B+AVZLU8AWJ5jEgaqdwbQqT0M7rMBPAnvdILQ8a8
YzxEXoN0hUbt+2C/JUg/9UFu7QXDF6ZTInhNvE6+W62ouS4yYSmF6ouV23MZ
PR40HJuIVaEBHNQLJHB/3RSORrvonFneyV97jvnkoGhodAms/kiuPfDJ0DUL
cPmCwLefCqjrqGiH4/mf2YOFLIE+g96TdQayFjBro6rMU7AlyjvEMhXKbf3A
nRohPbZyN+vj9A3vXCc1/XxjQtHiomaWat22rYvGrCf5WmZoxz0Iq93NJotj
dp+QvKRlVuHtzxJdrT968Maw8lhQLuNkppSVUYh/N+e6vlx9kaWtFqlrvA3v
wf30QQlf8Twu/ErA2WxsEp8qXYFoAxikwMV9uKgGDg4uKzBEn3Z3pjVhDlnF
iPbdtoEZ63V+ftTa9xKYsNvSSnplhmtYXIgDQ7nJSt4poGC3/2V61m8ztvyJ
xvWbPGfLFPQCp7WcLJ286cR0+HnYQIFAFIuYwfvhM02y3DDr6+ojStHLMtcm
YDYm4C6GDexjWKn9ApENZXK1UMH8eUhCspyYOs8zgmB4JULudnkvb7zvxwQK
rG6lvEOs+FEZawO8h36p7BlfIVTxiTjnHwxGXpxj2WtnaZX4hDxiGFE7NM5a
l4d9MOjiehNNit7691P0NUTo1+YrgAm0bNO6ga+j3+H7AC1F71X1Eak+gz9r
mou02RR7/c5v3LnUTtnrlhARBk+9meIu0gr4dE5cNnYDBQS8cYvR3utIL1eN
DjYv9cfg/TnoVukrthVOza4gWdfXwGyOEyRoVwwcIMnKSsc3nHchY5lVL694
Hw9G0aktsYgK9miBiHg38dn4dQE4eRMmAMOht/aSiTaSweZ3hsJ9ASWN2Kli
MHSd44EELHJBm+1qjCfSPbQdh6NkpDlyiYqhnAqwAy1BjoJVjxt7UAKVu18o
BLzcQeoHWiUxPdj5mim7t1Ccs8FsfRKnVv4UHlJJPmyqTz+nkqKBMEDyIads
H9KmpoDzOzQjwdI77NxwV+XwSg5dwn2ZeeLIHvGKf0YxH+yOJ6imXPJhErCh
p2PssU1EfKCtDQZNwRp8dkwA8yHJZB4TdSHFqOWN3SS1Ognont+F2IM7zpBb
BrX5kKWjG4UFkk/a5RhXzr3iVTqXDguPRm6KFZDRBPHKGO/yGvJL5WVFf/le
xlJYH/NGkXTmwznfh/DfdGi2oMJbL8p2xQzkU93fv60GIQCV6jYd0m1OmfwO
RjPMqcK28I7RdQrA2oJv9aGS7F4vsaGZ8iTMbxiPNPPUJnyI7obVbA74ob1M
BIi7K0kV6HBo3cW5lF+1IOE3uUeMNiv0PIG0Oz40YhwWz8XccpcSbZl00N1Z
IhgXeCQ7fVpf9Hn8PBf44fq8Dtll4CY2v1z1tp0hv89AiWb2sVYUqZ0Rxlr2
Q0axON2349W6HzSsrDjMF5l/+tpbrrOqhRYcdIvl4lVWomyWDwCHQ/sSZUgj
Vg6k8A070Na6JFezi+8TyXOmhaz/cK/E4Kq7fNNPFiTLKmvQUUSAI79I9R6z
FEUxbeMIQq8eCuO3dllE1H5Lo6LNeDemZPplW+VMZibGTqit+YnzSYe+tgrC
YXg5frvW7CYUJQKjbx0gUMWVxetixNlRSw/DJHMggGa3zIst0XFZkiITjhLS
31QoT34WvjW2dhBJhxW4uqQ9s8LV3eiJhTPHrkU12fFI75cXUxMZtq6Y+X9T
IcytvXcw43OdyluAf+3czf6PvFOuK/qNbVQ+sArP5TZSZrTgDhWbyRjYXOzA
jfv8M5jDZErRFYNH9xDQO2IOhA5RJZFJNTVuoHy2H4nKk7WtcvtJRMe+Om2K
jnTR7Lzxt+viRGS/TTw2mjFqOsXnaBxcLxL4HX7qQpJk0+HBv9tITaQ1X47S
wZ3Did26Nn1mk1cEte0SRCMtNgIXvrKE0qdHtBx+c+opnnaNd5fKTdYMw/tn
QDsubMMWTQb7nXqHBQhcH36q2Tnz7R0eL6j+ry72qBWl56uI32qBYrnXbS1a
kTwJyD8nrnHJXPUljdHIWufixPCAGTf0RF984rxkGRSCF5ws4VCp8YZZogiL
CHGvEs5Z639XN76sKM7EMEolvi8WfPkQCuB1Mgx529QxxMX3N1ZA8Mm1s/ig
D3Y4VRoQFE/8HfBXT/mfnrwhS/0Xc1nKRut7f27SKjioV4OCJUJf2dRQ980u
+zX+yScJYf1PsgoJbM6S88R+S3jAx29pJuUedfkJshJaJ01oW+GyxnqN8XZy
KDRCgGhQ/t1HWvVEAoShkg3+dzmm9TlYCGUcLkAc3AR0+LAC+d86VZ02/yBn
fg4xrlS7O3wu00fyeumJlJWx50qdmwfHTeu4ox+kUXVLmZZ0RrLd8AnZT8fo
bAmjXrpEcOMDOssPwhurr0Nad4FswtlXHE0MMtcwXJVGVr2w1JInlo0QnBZO
C/aSHpoV5EqqG+zg6Ne8d2FrtXQDHbXHJYa9KwytLQymKOI0PESaUjtTf14d
LoNNHtSS0ajfoEUJ+moiKF9kA5qj0jFJHd5VBzd3pf/he4WKbAbNURpgDy6j
oZqHdK9Zcu38BIM3L7nr9tY7h3EyEEyv60P4dqkYyhVHd7YjxFEUF93txf/E
Hd1rhvJdqOxFejvmbW0auI60X4//q6LGvwLuTkDV8RLOTNcIx8GJLmAXEkBk
JlHgpkoRAXdy4L66Vowt+OYNuBW3CtuYWVupuWUOOAqyQIE9VSPcKUDC3fZ4
KeExAmqQgcKXh2nDtZC4dM8EvH1H899bg19q4zdhWhiLNCYYuV20VXS7w9Dt
PzLhcHAI+/sSUJK/YCE3sAgxlUpbbW8vSPy+/bEt9L60tHrvDG0augQQS8jU
qB1MB5O3FU9gf4dTOVjjWa9cg+KaJuKjBbngHmKsluwKdze8CniN1fGaRzAV
yw1SeFYzAJSfGnuUgOqd9N9wGCjRY/2VSlbaZiDXAmiTL0S8iqeJqmdRaAEE
tYRYbfYf8DMWjw6KFOnX/y8K+mp7fbsBqzwjEabdgEFTcwF0+51ayj4xk1WK
SkwTy2CyxE5vV+WHBIL/fqIYB3bnFz9rMEjQSkI8+aOoavaIfFRSXmMUL2x3
Ky5GhneV10I5XFYSKhIc7tkrfRj+lQLUw3kbiX/12B4xPKImCv78kInVTayp
Rox6Dbj/pp9uPayRhMYVyLOqxCPeIERrTw3XHlZlEyfGEOvP8x4nJCsTa5No
QpMLfriAC6af5AvqDt1uvq3HNhd/oqPlqSRxwErRIIwnHcejWKqesGohXck2
xtZchTeGH1ULx6pgGwAMM0ocZ4VS52Vo5GHkcsXSs5OOpwdxm5daPEjdVYLs
ZNKvBnDVQNf7ba2NjqjXqLhK8dMkuxUCX5AyT7OPiUm0kdLUHM8I/JIhDDnh
qy5c02Ub0lkK7tQzXKMeOmC15G8Mx/mZQ97DvAmoQnejkdHy9OrX5mSGurqf
BX+c+ti8uEJN3YqEOodyKb4/GJ8Atvnsu8bPnhzCW9ED1xVy333YE2W6Yecg
F36uanajsyM+R/C0IEsvi27KRwdpQ6ZEba7R3QGRLk4KQMgZ+uya6rjwkuPQ
ODi4/+w1xNjWK9f4bIjsEJtSrx4wBduPgdA2u6FfQeIMQ2PSE4wEsToU+JOm
koiWfrH67yUjSvavNvpKE+zS1eA832riLC3txt5AmlZd8Q+hVGU5GZ6a22gR
xYBsxM+000n9AAOJRLEIvgseuhCZkFNsPoctKBNCWHi17tbNruC0Pjmdwz8t
ZMsr8A9yQe4YCKm5ilvOzDrIQh9TFs0M7/sXrFiLzP0RS0knaTscfVSTglAv
1sQgFHXp3DMImW3Rjh/h0BxSLKqW5KA7Er+VH8OhzzSGe3/uHYYVx/1V1vl8
oHhs6gRJwFlYAnKkHzjEGZovM4Hfvta2xMxaXOYm/tLZKPeQBep/Op8MNV8I
Idy1D8WnruwT20eIARoeGnQVX3TlYy6wyRdOe/cCQRxd0buAYeijFFj3BGY9
Vcvj/swRmk9mx/lihwahUzdVHfl8Xfhu7k8XVrmZoEqWfvQ91jhceoSdp6sp
+tyb1vLOn2HjWRr5lUWjFMrNo/tApTfaUxBbtmQZImtWHMCemxGmkn43Sztk
ykNImcfWtHE7JlorhcRcEHAqLj4m0JdsXvn/FbxxwP7pF6KfyUPgqlcrJRd6
SnT9lJ1F5iMRNeknA8mhg8sm94woYAwv3dFjLNW7MkVEhiqI5qwhnuY+xYVe
lGiYfCeW3dLIwhPmV2X80JwJCvzVuFtodGr5dd7UeEY6PnNSqfI+t+0Fbh2D
v1B0+queXqHkcvIkOuWBPhJrYGFjRBfqVfKi/SKhec3e8s76S0QClzqKVOy3
Z+2e3NJqeSUpL1iajfKfkvNtJUsUaNSwlM2jXsz0RwdFcG0j7fqnuHK3SHrm
SnpQ4sd97eR8jYSkh7qv13sbxugpjvlPNxsohKqoT6Z7OkbdS6GkN4zR0YBn
BJGUx5ymSktL8RNwJwwhLvfv1ABZtDopJ3h01QVwkvsvRDBLkio/X+iUyvF7
OUkZPmXR6HNoeihiBTUxfc0Xqs76XVrEpkpeu8JwAceTLGAvZzHyFvWDckYC
3+vApgIM5yzlYMXwvQ+NFNbVrtaXSahy61s899QjC/J4KNHDb/ucn7cyKU03
7HkuYLicyfhZevpyUZenujZcAcQhWMfO1yE/8MUXGst5aB90jL3PFlubzGCD
C5gaz8O3lH7c318FNVGO2j8bRVwob8hlUJHiTz73aNoZosE5fu9E3KmqfhCw
a+Xa3HSCNPVTCpYTDqKck6W3rQRR2AhulgHQKGsz2FDb4buYfJJ+WLOjwFr7
gdoifz1csXpsLKFiHxc8N7pfA9epN0dhZCOHhBu+CJjb3ezdMrE/v0B6lTtD
jYKvWDj8gpZugD3OHu18GKrknLLSPMJr/UWI8cUd9DRK/B4YZMWs6NWQwoGf
1ZZv9qLUuT0tdd9Risp13P1t+O16KV1IG+OwMvtzl5oeke14A0QPdoUSCIWw
BIV8yHlJzrEVam6LPpYoWZ/Z3yicvFQaoOz16NNhluuRNrFEc5cDs5FeVvPq
3krnE4/vyuil31TPFrsRLCNuZ3uF7MdezZcxHcAP47OAttukcnBVo+Sytki6
7hZfVBNGpfQGlyT4mpn3UlOD83Egi/nmBuoyBeHptBjys7JlduRUAYFrgsZJ
wt6/4GmDuhymsWinfT1hxfy5aZG0sZ92rJeeEHUCmWXdUcjSi51ZM+agi1/N
GrF1urq9ETgn6/sbTwuOG5osuFVPE67AIAeLVPiLuqf1DFhCI5SwjRIWFCkN
umMD3StirdLt7kvpOEtR0O6liWOX+VBqhdTMs3LYcoGNjzuUptsO216QhhYQ
L8beCvqRcWxTerigsu6Zs6BLbSyR47hL/5KrRVbj3+Sa7bmzpBu0GNX142Vl
voeHfDjmK2ikB/d5FFjDU7cwXqbzPofaDsiI5Hi1HDR99Kz/9faFoamYUSEi
fu1lCntlVa4IDQaBLSjEFy3Jc7T7JbXx6jaMOAi8FR8lBHfB3fBUySh0VclI
Y/R85ZEtsH/j7thaRmWSOFlCU9aDB+DyrAbZncMj8pLBa8KbxlNfdvOYM/8E
WG3Fkux20xWH4sLFy41w6c4ESwMKS/hmCXjqm+iaqRhK7IKJLye0EuD54LFD
EAsoSl/tEyfYClyb/pGGzZPUj5Rl4r0VBclzpd/8kxmeVMfR69YZdkUv/qbk
pktG0b95uCaYZ+jiJ6u7C3gQoQgLS56di+6ka3DClHBd2Hmw0bKBFWVn/99W
BnA3shY/bVJ7Bvm6F1uYGp2ViMInRhZiFk/ebP9/wyHbfLpkXJWGl9fB7i8E
VoGn711rurSJZsNokw/St7q0v4IHyMcTlCIX4A4MzYSgUsCrWMEWlW0NmgJr
oMlrVwnAXR1BVet3Pcdr8G9wS10cqtZhZuSfVpgbt5SOgqJ1B4xz/RX26WPv
3ix1dRXq+Q9+B3Fa7HobwPc906bTSm+rDSXOkivNcljr9yZnmr54EazCpU3a
TuWp4J92lfsOelKaJ88PWRBzS+zHvrl1KrKeCJ10hsCSvL0D+3O7nAprZtV4
9WDs9UVTVJ5myqSI7brf+yh9JK3KU5I4legarqdoLH4Af2db/4lbtEk5dERg
PEYH4UGiETheQ4gVJo/t6Ian4u4/XjQ9D47nHMlQYWReujIzLJuWTniOIXWR
7U9jYiWhjqQrowF15T2MdxCqPl27GfkL8W2CjzeXtj6koD139xjPz8DL8OoS
c6G4SxuNbrWma0OjEl7QRo9kSBfW0dEXxPhfFdUnc5T9IcChns1wEM9Td1lN
rL8dL/pYb5U+l3/pUgfKWJgyBpPc7Kr8y/4OTGDn6r7snMcq9BvWm0SGj0Jp
aKPBSg3lRjJlVA8nGuGiMuBbXDk7+nYdPWK0fEWQo8QKsW4nTB7l0WmyaeaA
WciCxvrFzXVUOWh65zrCeqx9LunoDsjBIPt+GWbTlZThHj1BTcWXysHfpAKM
7ZQhIed+5vJ9thF6sQvEj3L289VcKljoAvLxhjMFVTvk/POx1VSTpchv4J4/
F7JM5xUcGnfoDIVJQLiW8qZxsTMVJ8clQxxdw2LUdYaw2hDOt40sxTqbOXik
qTvEOKQspXa2roODzwVtf1sy6F9cNo5qexL2WbiqpfqmeHRw7UxeMZn9jUbT
/wDObnasTz+E/hXx1ExHzkzSK+M/Nm974A5BBLTI0cTkVZfsjx7sH05BaTIG
J4LHeR4F1WO4miC4+XbSCFat92Bk+WxmdMmp6fiYEomF/N5JYos9NAOdx5z8
dQtEg/w7xT7E9w/ufixH4MqxjTHvhSUDQZafqQbt0k99HxqrgSmrufXftLf4
MO5KhOiUKlXkRTD7N8ee7M59QDdNv1/l50D5WvDktmug784gg0igm/nlrXjV
EA6RgMSwIq28okYc1eyA08YSsU88k7GNJNPZ2tH9pttuNWO9w/u+E9RuncBD
tRGQwDt1UkEwJ6I2A+A5KwWtxspzBxQJL37zuTYqwVQ0RrextAnrW6l6dduu
riY6HyXenD1kXOOGzSNUm3EzkHcSYIsH0M9V8RXeccQnWbNdaApD6PtjJUOi
ZgiOpKeMaU381F6tTnapb53i+nLFhCou0pC+5Sii8YhUx+O3rBcagvbzeaHH
HxKFyEeH5CoUfSgApWwQ7WUAaCPJcusqqvzmoSF4iPWDHVSX1cHv+lxnrt7L
+JSqMLJADgSRxEAQe0je1ODuuKwshMHwAtacTGxJeWX75oLFLnp1pYK+s+Qs
go+yG/vUKQqbwuduJppk7T8lyR4ajeNR0c7rUlWfdGrp22K02iimhnrCQkQA
XPAcJuq1ZCdFqLzPGQscpv7cS1Us6tncPBcztTozj8VvoAD0TITh/eTqTgAh
cC2orEAbNLxOFS1NmFeRgFEyhRR7NllVnonStNwAB8jDot/O6ZyCXfeai6Oo
xCNySf68bLuWjPXfAifxj81mukTcCoVCguD3LeVDJzldzA0qJPlUffz++uOv
d65xCFvbm/GijAjxEqTC9ohbMK+ff0VBEMvFwd1W67OSfaIdgoTRnDdp6acq
UaFtvgfhPn5hRov5JWhEvpWNhIKxfkMgKQ32f6gPLgaVhIFL0cMXItHqhcH5
ncZ/XjTyVg00Zm3snKLytTfS1RVap/me55K5x0ILibc0VM0yQCq72abcrZxA
SPOIg7OAIl3wd1LbcVnsRrkQL9PvmGpom09JGp431MoaDiwB8ddzQ5sl0+/l
lLpQhJLOOsWqUYSVuKlDs9a53cBCgsmxekXmMAlhOfPx87FUT7q5B9GPiba2
KiF+ow/yhBtBLlBNJcASSpLdH09vQWsUpxBEkebY53fhceHfNlJ9/2l4ZM1l
I7DbrK9MrUf57QNxgIcycSqnus5und9k/Efcbs7nNJnvMdNF+/lEjiDzPtNG
ngBlHVRnMXlaxspvOe8NYwzgXA5FNR6smcvLk3mzyxYB6F8I/X/e59hJcJhf
EqJN9TRqkrNvnSjFEXPTSHAn9hsBLicQNPdRNF43/vF2vsIwn16+L3i7Wnv7
XFImaFqlORWaT4JaAxnWEdKjGdIvV8/qEiwpZ6ol1r7D+H9IMxg59R2RTTTj
vfuux5K4uWXZa0HfAUBIEsZ+mMshg2wCRjOnNHzMgoU5oGHFzabqm52VYRVp
LJ+PeOq8jvIvJruGeZdpXplbHDlHbHdZ89r1Fj5zo2TeQjeEPGoKhjS/Q9d8
wqiPXBhEFEUTUw6ttObUPTNxBk89w3gWnx8jH1O9aKKruMpplIYx0s8oR3zt
mZ/wiQxji8156e9prd0hslLNzvze7+D+BitrmSInyM4zQNoIwt8jx+JjuNLr
9dZciJn0/bo1JVXJaNDSHw16k+veb5YtW8BEDErZACTA0vayFC2ify0XZ0Ba
HeEZSQYYoifIBezbZQouSXDg8UXU/rzZTM54nWNfhIUPsConZV7oQ+ijLghx
7i542MkEtIz25M/9hd/8yNSgxbTMLpXIlPincftt8CvTWNHdFTrpMaJBtUtB
99Wc3I9I5EdnQwN/QJYEhiHomuZbn8ZhcbGfE6gElF3CagOBPFrCvMXoCEqF
1TMRMucv+JmPvod1e0L/w4GwGKzfO9i9yo+p5mwBtxXibSil2bwMOa3jtTUK
72yIZMitrXGIQSKLHjynEr9/A23AJevPvJwLfoi21jRQe8IcvDgGUKuM05kK
Z2ns97WGV60JjXHupf+D3ETCGrTR2tWhLpuTfC2pKcwf/L2NRPh6HWxbAiWt
6FzafCO3zknoO/cClGi1liUWDIuzIGE6/G0PE1rQazesx496CwJzN6EL0188
NxWkFYQaS9d5tSB0/ZQ76emulw8qQnA4DnTRJ1+PSSX8StyNbkqaWmfjU4Sg
m0RNi7PKwssN58g9akINwKXDb01blNTWNDrEmKOt0x7+anpv2zsmzaqJ2Uxs
si0uM8KtYsd+2gknok/ijQvvnQgH1UFmZT/NjJbj2NF1JPsH/+URkxpdEB4O
mU9SC9Kx4KDRQctRiOmTcm+jUHYz70xCgOPMsy9i7RuCkzqz1OqM8eWQJ92p
6LwPUFQ03nZTX53+/w7IK5kuf54dOJdG5A3S92d6KBZWIT64NvLuCOdhgPCQ
HJy8ZxAy8MDei33biICSkAufcCmmlEE2OiALuKDSNVoz8TAycWQsjoVL5UYv
e1kNULFzqhwVM2muyzxzaNUbdQtHO9myghiWznYqbzMczTsOZrwa0Opr4wyz
7eSL8enyh3tQYjZb9UrG2ZiNSKj97+1azRB4IGYSuvirruHBzs+Jsl9OZL9t
9hU+hoKyfv5k7yDCdXTHRP//R9msrvBlf+P/LyF6fhRkr/0OOZnfKvJK9xJD
h2iW5FDV79sC/8CHneO/G+hnCeu4KFeu0d8wjy081BZPGmk/N55Dtg7KV4PB
BDMlMk6SQOOOEPo+367EEoAE+hU/V9fRZlLJnpzxt9+DzwpvB9vKO19fjcL+
Oua0hGwqKuiwyKiW8RdlqvQtHo2Tuh7odQe5Ve204JUk7VVV9/+gWS3N/PBE
1tg+mutG7p2pOQ0ZYkGKiHFP+0yCJrpfoLtmVCl2E7otxszP+kC2iP0hdKJx
g8kQVeP8lUnuzKTPbaA0gjSHnzDT/ZgmbK3OZ53mpU1lLXmz6qRcOePAhkTy
I8fB4yOnu9qBL0TNgPdw0X28PiTlsGVf4zkcGubKbulqGzkffQWQJKImwgg3
4Iza4nyurw7ct1q50ohsf8OKu25jxS1J+3Vlk8buoS2LqMPVY7r1bVF4JFg2
neYgaH67ic8MAa+n8zJ/PVDnuJ8FhVGXE9/0+oYq7kC3a3L5TkxWuwD6uckf
Mf04lW//pC3aWmMJPwx4naU+QIgocStYL6PYl9dl2U8aQCzXrKHoAqk7CHdU
uY6sB8d2Gu2hEYhJj/33DTakXykoYUPQJnzomxk5OiN6FidSFG6et6h55/nF
AEUNJFHdN5/47+0vKzzbcWmfEnzX76fYG4cpXX4HsSzU3uDt+DJE1dhtHyFf
KD1AEAU+Ael2UOpaAunQWnae48BgPp2R9t5k8Nmq6UiFxDuWPPfw83vRqfDs
cGzmecugh5uViE7OR/yU+SpOkdwKrnVEHGHGChAIXt13o0hpWKRivTkKzVFI
M4+9+1qMKTgWOyavazlcuyL8D36LApXiaevbe9ZOaikTmiDm8NyCGE42Stjv
pJSMOzo9a6vvYnlwbkcmgxgteqHT+sdaC4TffFu14gufcg0tnt6eauyBd3j0
NeuDHYghK7zdXOUxVn/dmkLIZ8u9NqphaTlviLHaIK3LkVYYWIuL4xcAibLo
k0r1esGm8PxjCm5ishiMrceHQcy9ilWtzyM7C2PMwAVSw5H51/9Q3NveQgqH
LF/gcwjgamjSxJxxWcbidCMvGxGeXTxqrmzCXYBUYUqD1ePxAwWsWX+60tHu
XnhwJkm6iPr0f311UBjNTB2+PMSdswDq/GhH4ctVTxfSNCFfVuzoOv7J4kmS
PdcD7NRwjQz1WDDd0BahGd6Aebl9ty59Xa4xPefWNSW3Dzmr0fC5mVcreaCD
pDbRW+zaa4h0kk5PjR9DzuLkGQPF1QO33xB/JYlupKeJ7kLV4GTHTQjOgE7w
yRJXRitK4GNMwam/R4/5aliLfyyT/efeKt+3TDYZBWbXgld5AX/5OPxKoJmE
8ntPwuIytGS123NGoLGZlZUHgHobD+lN3lwDzo73E0X53/s/FcNRAcD3DvjI
Wim/0a0gKNzb4ZvLjpeFDW2FSm3kL7NCRtCY7dT6J6rh/f5QAbaxjyjbBDrx
LufW/vLJ7Md/hOvlHlbjEZ22DaZRzAb5ZX4DbB6p5W3pl6zgMlOOfZZdHcsy
AVjn6IMpTl2g/JGnsB9/54poYY4vTRzRvXNXyqXg3B1kRjskMBMl0IlRuOix
HD3sfTYLevDz4Hc0UcF517HQ4ZsUZEa5AHwrZZJOGzGyAzbQFAlEDToAs9XM
tiIu6IgtlP4Kt8VMrUr0nynbD/1kFtlPGy7vQN1HPYlFNk8UjlE+YdviDGx/
SveASx+vXZSyGduR9hCGDnScVkJf+rPivjAdxT9rOVI1cUJKAPP9XlszJhi7
mh+SzulDl0phrLxHKvUKD7XhUb9rKTgj0029YQ97y2lHj6cN8ahXwEH9C197
nKUSRstoZ9lYvHKDYyVDK+5PiVKKTuasXJFw7pyDudYK2IWeTewXgtlouLSN
a+TXIL2iXQ3srzNIPSUrMc0skVlZlvuEkyoKJE2WnucKR47d1RU27yIr1z+b
TeGzpNT609TwYEyOPRYBGvJncjg9XV7KEn34M/lpdnWpiOGDiJJvv+aZTzNo
SkWbDB8XGml5EB1UvjTGSSO3TLjcXH2Qn3Acc4qIRH+Xhnhwi6ODH1uUWvl6
eFxBLGrTJuBrfONxCNqM1M8ZC0YagY5blyZi+MSkvXlDnLGflaPEv0L6k8bA
B3EkKV7MPRLGNaoMqlOYPAvMMzYdu6jTWgRAqkmQ+IoJ2zOytp1EBSzpTPYW
ZJA54DIm7KI/E3FJzcxfXS48OlqkLmBIg4qWhbnvkABc7OUMLUh4vQTyEDkI
v/0PYtWKcKhCaDC8g7Tl4BTQvjNtDGjWd5n6hVwje167Dj6btoULofIbkCuS
3BSXsA4T49liWWyrEVBfKCH/IojR8D69zkFxVhZotwFCJFAm4fjkeKCze0Hz
P+qChDevY4bJ4k15xLKqV4YlDoTdgB3qGUGzLsCpNdq65gKFGpgMwb2uWaqW
ypbNQKGx3GaXtVdTGCjzNgWilAH7UJ08bmsuqyOi9FMQQ+5pkGeTAtbZ7YK6
OMmzqXNSyw88ZDq2EbhQ7rPcycYgvCLlmyImUSciHeKbRtGpLj5qIrQVB7/J
SdvbSmGfzbFDB7/c1DXVr6EFL1w2X00gDD+0s01D6BUuw1kXRVtF589PYGWr
zVibQgnbdL8dOQmlonUR4hIFE7PHKO9tzITNzKP4HqhKFprPItfZDMJTWiIF
d5AW+LqeaX/CB2JgSEmg9F23q29YjKSh7xMM7etXcuE801i5edDtuseCnMqr
Fhk5NHf3hdSbAhtO3uhaIv3qPHUbgWdWbtnhkkNVJojyAEM1zIBTUnHvI7D0
czRT8Hr7KCjatCqIfKw8s3mTk1wg5bR8KWlQVTUYpYpvovpdIROFY1YAqXX/
CXiUEV7x5mnKN70DChIOc2HeqRdqLQuNoFkwP4QppsEwYrNP+0XSmUDhcMbO
q6H3NQX1Z4313JxfdZKYZZcDBaL/GP9AZAfcJ8c/FJ6vsCXwV5ZtpYUGnXmb
J3cnLXo/Y9j9UYcLLG7IA1Y/xbh7xIBJb8gXyOzemHGUWr+yRqObBOH3hQ79
P8qAXTIv5ueNe6AzSAIUqK3gnY+LWQ46R9jKfVkZ9dzJn7689JMK6/lF0FFH
Q8RMkRwYW9mppEI/VWKyn97TRZEFGZrUVEm9ULecR91vUwHcS98+LbaJSSPp
e0NDsX8DqMhu6zZVojM0NOPySuebokgqTxABYY4dkG3m8ys0OxDdUIQxAoZX
r+wtEiRfu48ySgZ7KpsS2+UoyVDM/tbPOA+hn4bzG5ieJmJrDgRg4NtoWfHh
42wBS2sl3q2UzCG6sRPE3buDDCBjFFLCGIKsEUSaRo/29/tpH/QcMjIa82TG
fWQT2tDTXtBLQPFtSgO8P+VNr3aCyBJJ5drsU2KzNg/Ld7wCW0VFUqgr+Wna
z93Tyt1H18AomVaUOFK51RyqRVRGtf+I4jgaLHeuxcWLKOLQ/J7PXU+NuStK
eDKwCjHk8KMGKGdKyVgIuAUxqTWfcfL7vqv1yW9AVIJAG+AZtmFlDPX5nmDy
z5F4Eib6DaMNfkBZbfOU4rc/KvDoAHhjzJKOqU1y8s5g6myoklsAHUNNpZy7
O45qal5A/jKLcIQyQN0+4AC0JzmO60SsumeNSpZLjcPxnZbHwm3gtIoisZSt
fLUagPxdfr9iFYfisP2yQ2AC/XqFRTMcXvVj3vWvnoiU1U/MDiHAFpaCwTBo
5goMh9nRzXiFOObjUwo51klP3mIqZPY7Z5HRVsWCmRyG+FQt9MAapehzmACz
F8v7MLLgnPVhHNWX6mjcz8YS5JpeVmY2/YaG+IvfooZuJUd5nq/+eeqcfs9c
fW1U7WzKDVg58PAxlniW0P2pp8cCctEwIKhuUrlhtbuh5BWfPdPNj/ED8FQ9
hotnGXRCfgkm4VeVqI5rnkNHlNyz9HBLdrsSSbaQguAsiCXwpRNrKS1Dwejy
DI8qLY1MBycp6REMOZ0gvJNwyDr4d017y6y/xMi9viKOlGFlrAsJkBoPWDVw
ddd4qX9BV9X/X0kRAypVyOSdxYqNVggMfWoP/8C0Nae3gF9pRVx4zOFZJi1V
0VItpeO6yV48pM2rV+BvDJ02Q6mreDspZyJyvNoMTD3wXaAOHkZv0+gho/fA
mzkzP+ZrfI4is6m+VomhGPXoAtRoX1oH1njH7P8GCAisPemQKeypdVO02jCY
7DFHKrBqFVel6W+1fus0VL9u/9o8GKT7lx8i3AAwzaEMoQkJ8D5zygX7/cVs
NQ1lIe8R/nvSrT6CXqjgo3FAp2OJJt8EYTAsntobtO1ydrpvqgjZBRe/fQk/
sTzl56ZpUXa/BXdELXHCQOwZoUfikM2XPyRUesTzMF7fLmUi3OrllUJQ5R4Z
SFbmIBokohfufhCMUeiyDsNu8eXZGk1qmTmpkmcerqtIeZIbenSd7c3ACWOW
xbujO6k7DsdOGH44a/k8tzab4oXuyZ28RWA/36Bn+Mx9Jl8BfRENlAZCdL55
kHdu3pOSNgupAsBim6Up3rYtMvS57RtMMhDoCgIMVTkv6j3K3VhrGobC5W5w
YLCpJQMNXmeJZ40WdOvpp9ZI2dt9w0OE2UgmcBYOssU/RXDk6sHL6eMH/ayz
JPL1SkYIi3aXff4qoFaYIwla3wb/dJej1x4Hz9gkMD5kN8pzqs1BeqpvE+UA
9jzL7BkTw3oe5Vl7O5h7LN2XFRDque1cPfAB9tIhiP800zPoYPG3IrUd7t2Y
tO6ajTCb3Yf6AH0rDUj16En+4joHNwWzFuZrlYfA0+SZaJAInf3AmsZ++vWi
zxFfgab2hxbHbeRWbEogNewTrWYhozRgSiXe65dj9y82Q9C+ow8zXz7QWFkV
MSQwA2ne/e2XdQtx8W1bHUDMgngwE+Lk0gObxRHaofZA5cpm72Amu4A5QZDP
7t1qPLxk5MYPwE+gGILSMnJ94dr1NKBOEuzkjCcT0kaTAA8iBIWY08AyWCWF
uqn91ck7h0dFisSDHkSBZz052Q//TJFHA3i5lF/bpxVsvbAUk8Yl/hqgZUqX
N5a/Sqm+pQc8hYaQ8sEAqJizl/FsVNAUHhJtxN1gojkHZ3UpEfkqT1zdnkHN
r1tbH2RnzX7kzgW9hRRHuOVwf3YXhi3Pef3GJJ8DQ8kQ3duZoXQCF0/vo764
bNvAsmAbESupb17HeXVdNDu8kNm3bjCaDaSjIRNXs2XIbVcrvabolHLN6cNh
onlUPZU/u3gnFqlQvG2VrUVWF7wT1J7dPvfLx4JeFidOPP0y3RR0gWSpc0o9
w1ZnraJNL0al/XaszrTakF3wTRYc4FxbQ0Qnh6NcfzRDqRzZOpaLkQWio7KL
ldc3CTZvyVkIcSFYltbzC7qOazM/qkm5LIaVlbMK+v1J6OQiVHvqZoIl8rtW
rdA8xrNUdZcUpGa43oJ9FLwNIqqd23UbDfMW9LnlY9UsguIDqptRYf9jI1cu
Gk0rAEJDkdR/QE0p5ktc+9SNMTwIvNgab83lokdMFmBqEJ/zrDmlFAm8Iij1
EFMYX4SswbPiehNcVt8BdnXh0i4fqirFD5gpXjAsMWvjzOsyXJIRVw44u02I
8u5uvMV2lp61lvVK+CvfqAab2tutd74g7L/b3cfPwHD0QLqhz58l+1iy6Ggb
V40YX4A7i6FPfnNJAnLtRjcGjMGftySz5QAWTkOjUxFfS0STQwTYVOsoLrNP
IDfrg7LgPrxLc30JrNs28dTxfn+HYTQ6d3pfcKg2Eopco1AfUvkCP/BtuRfi
+T6ckyfer8JX6teCx/buxxDHDniG/6WR3HAyxWsRhHkw8lARKS6WMRrT6fu+
jhG4N7/n6T4mQe+rd/0KthUTfhPig0dMeUfdvGpdu4XCaBmQKAg4V7yRFAwG
/s3zUPm65MOEzQvt8MEhU0uxnUAkjzEJmKOC8WrVOcJogYrZJvEjD65u1N1X
wIU8gY58JGPKzJkNgYfC+T5zi3RzBg695dy5/m3/Z/VK0uSrWOkklDcvvipI
8y1XG6VxFOkMLVUkLfXDLfFCCqSe5foz1aRqRdbzFIxJHIs2spfvLCzOHlj9
DQ6ULTMBMhUiyFcZzVs7uu9aMKcpNMD0xM5dEKe26FgKkoDQc1Gs4baPC3dm
IRje7b6V4CLCvo80wzRiAZ0hLxgOH8JKnNSNr4Cm0EVHhVLgBJlPAzyvYPKf
wq7H3NVF2JiVEqZSl0HjKnWCoGUSkMApvXC6soKe2fUpqKNToyzvK9s/lJpp
aZ93tjXvyB6jY2bODrJKICqOYRBA7wYPfYA8YKTVk02/IhoPmqQwLwqV+h6j
6B8Wir9G+OyOWXWE9M27Ty1V1RyFLnhLuvpfHHJAckNTX4IJ3ujj6mrcK70D
4qSFxuRgwEGslz9cXXN9WJsOaGk/wth45UOW1E8LSX3BjT/ahtMjbwKaDTwx
E4aD3p/cypaHbs3nMlflfoFkBogF/alx37TEqJ8qmc8H7HAgrKIDuKHcCs+x
Cz/z/P5um5BEYoks6+YuFB10Wfv5iGRavcmq7zP9sKZZMlWnviZn4WKmYRNR
VSvphNsW9HBUo3bTV5g05YpscDX/5JrovC68N4T/ZoP88buZv969ZLsJIO8g
MsjsrexqWx9kfxhMfaJhLLX4sPbPgXgg9m0TLu2tHl50lmxMEjCYrLCk8VCh
iFfjkfiMPgiUxHky99/Bi9t2aGrUpizb6tZgZk+O7zn9mr5uCeR3C3H4i0Kb
yQ4ffKBWIeMSXvP0tZO8ganUCrUgLthY1oFGxCW1jOnChYngpYgnzWCTBOIr
uQYyaJY9BPXHV6crA/Oraxn77sXptf6a+Wj5IRNnQtSENOnNekAug+mCM48D
NL3rHgQK6eVkww4QnP9G96NWQJezS2zNmYW/SxyK9eCyF17mw004Ec9w0WC/
YlWfnI10UpJj/dfv9yUFA5flUzHWQkSvN2kUB0PVOZvHoDrXoCeUNrcoXf45
DqD+dCwlz27R5dkhzQVkdfJlatHlkoP7H86kUsQYuz6gyhTSNAPn9vtUL4Kg
4hMLrey5QWoonCO8ewudBi++Y4tWxkHuM5/9KXB4YbIZNxd68K+7PrFitw0t
khqcRD5g0iGD5iuHfLATo7GcVtHkYoZPF70AqOS4+1rL2qsHGZEqlKQJMy+y
xkdqx8mZLloPnw22c+0d8eHUoblCdMOEYVsEuPxk4RlSvSUzqigatU/3bxY4
3vjgpHLwt67GMl1eZ2kcMn/CovtZIRblcXkVlLnu9bg6loVolLObkHwIv2XX
DyHKYhFeJl6Mx1xdwMoOJe4nctkeGFkGWrSo7tZPzAamc25qF2JHid0Tn6cK
5v3Qb0UH2xB4JKxAHfJOYuz5gXBis9+CReAz1WMaVPdcGNb+ZcCPohMr3PW2
6XZWo85ftv5Ygs0juhNsMYhtF2SJiNQIrBbR3MJ+IydG6RbsL+wBVhAOPtXa
fCbRd9FuCAXq6N3mC4mm21iZVPTLBXgewxE05jdNNaaIzO9Guku+veF/vthN
Olc3cz8RdbldzX8QMZ6MGy8MEs+IskjMyi0l7j1lT3aTPVlyaLrZUdR9Mtkp
1D9DFQs87zqJhabD0Pak6mwJvq+sfUZV4gL5l1C1TmJQ9ESxsN3INmRW5nSL
pvdP+Ctf0diEautlTawv0ZUmuMqq8FhAutObVVFm/+PDp63K+pm9UATWv3+o
beUNorRcC7a6HEA8B9MVzSMI782NIAg+CtNe+lZAVZDaUClHJ53jbkUVKWp4
ZvxXnhYvgUsnZUAZMfxXrNS52aLDJLcHeSUeCKzZxoI+rS9gOF3rlp1Wr5KY
YeRZV4cqSCiAZonR3sbupPczorlcnwNnEd+f3S27LkspSp4crU3B7sY8HUG5
2LS8fjirTlJBwIOeeUdEm/TAS9R0Nzy6GwZ4pdd7shKFuc3nll1WXClBymIj
qZeR5vvz4dNTrzeHfpS6eoFrFKbdQT6mmy6tsQx3BZTCqjykvAltbBcMd6Os
x5fYhQ0OEU7dqoV0YCVxDDoPqgd0rvzzRqnCacSLub16I4wGERKdWdaMGb/b
USYpJfwBo7ZCFbyG1crDC01jqVIbK7t30Vz1vhZrgjRDXQMPDSTk6qjRtCjF
18X6RQPf1UapSWpC+6GiYWvnZCiMX//Tm2Vulgvz9IRMq9cBVe3PshHuZnNL
8dcl+WYXENMt5m7hP+BH+bj6psrU6FBp3Ixg6SocK7h2EHsewuOkQ9AQ5Dqb
S4uQ+cRUBxyUrJgrOtwBWTJQWYZc2GG6RiVbhrms01tKPUVyUVO4Noml+9Sn
1fPfBkZtzsxHhTqzq8KiEikFlrRioZ61Gv5DP4pxhQ68xnjp5fO5CI7uUPva
8euGKLzu91jAZ3P3CEp11yJi0TYMnqNQ3ptno4F8Z7G8z7Zz/z69iDcl8FBp
u3IcFvG/L5XnyaQZp8mwO7NbeU/EIAmzScmuB9W+F5bf1QArfoCcO4ZpBBOj
GjAGt7wUYB2B6HT7h+1oyJhrKIU18U35d6XLrFGjn1GhlzkCks9XhFzyaQK9
DPXRHzh5w7t0F/jlYh/TPzG++XUOCKDgxSq+7edldtQqvB5HCanWKkRm+w8u
X96DM3V15cqo5SeCMdBKP1AC/wUumzzaovA95+gu6Tzk7YcgrZgO5GErLS01
T8WmzUpXrLkebDeWLeVgyrIzvGkXeSvTFvCz/TL0txqQ0trk6/xcimQA4P+q
OYSbjsTWKpMZwMDjt3NiO60x7ldVUfdjwjfFSCiVnQrprROCLhR+auLpYfIl
tQqHp/cgiBxPmwWYnKO0p+qa74OJEnGBXoPpx+s8fdUjJm5WNibkhKiWESs2
EiHt9A/a6gOZ0f8TWKa7madNB+Aw0nr1owsTObT5ZpEglJCTx3ZPznfjomq1
iZm9wEgpSCMAMOH5ndINSPd/grTWNKS7gwvXVEoG9ZcbDSGjaA0EXVWxFW5/
HUXWv0Zb5Ni4eNa+FG2+I54uO7ELvfEjG/x7O5Ap3Xh8fvbQ35XKfxVCHiB0
llR0l2frdZlq7c5MiOtihiVS4aM8xi22TM4tb8ESFJ74PItPeaamapfEOEWy
H4ysrYNrkuR3LoYUti8ofkuJntgpIm6RpVGZTa6SLgtNWekWcvRnA70CtWex
6OX2uSyA+coVgofvOCzgr0OO1JD1guUsTZ/0L8E8a9I5ZHJ/p9dfGYdSI72l
cabUkoo0eZLEQzveCvrsKZjliobsPYJTvruXi9QmQvWlVG2JWa+0SEgnkzyM
u3OfGSb99WxBVzPuX5BI4wktxfdjXNILMaX4G+5ScmS/x0e5o7064yQ4ZE2X
fIWYi0WVzpDxtpDG4zAMiDJg1rT+1WWBpGY3CF58RgokhdaHMQzGrFnaTIxF
1jnJa2hwIIAoKqNdYcLTEjimNh737801ANzHOUiom1HT0fKhVa6nwsh4wqzd
nFUiInJRiIU52r3Mn49K4ljoJ3+RZ4Sw5ftzGSG/yy1dL8E2NWTsE3ucwUkS
C+Ct+j6bwO6NoylGNuds77YAq4rGkwkJn8c95KZg2nhLIDM/dobViFAJPoHY
dfVqV9vYf+t/P81lqnvRcVJN09U6khPYI2YhV5jfuVQO5iqQfKKB6j0T/rQl
59FPUNltzNKWDYEm3wDmAv7rICq+9UxFVGBsmWi0IG71t68ha580KcgT0gM0
ailI5qsAMP2oPPlhrLGyPmCgr41IUMXXp687tiWdOKcBWNYIrfxSbLjz/Ksc
Qn/BbuLxHM6CZxo6SNqZdd6BTwVIXVP8c1+p9CXLNBh1Ds1H5yn3OsNDGHEq
O1RNmnySBD7KZTzd0UVKWg4l+ZG9ocveoZi3lrzoM8u+LvoYaX1meZOWujjH
qhcZyUY1vY5H0AiYvL6j8Gy+29XVWAYQ1+/HqmkwgKkF6QqJWeADGh7+bKy1
fTZbof6ZIDVMX2a080i+N/h8UiLQElipMnDbwUuLkxqTM8mq+yuwD+t3/UZK
9l+igX1aehS8v6JXnNz0RiTtJqgvK2IXCTjbYAjAr7gfS9l54ay8icDkNo0Q
ZXsRtAydbkHsH9pvHx+u8e0/QvmYhHLgR8yMuJPXwVM/wi8NdxWPe9NmVlwm
LfAZWyV2EYK4G1baXyG2D6eYoPSaRMqMzUZF2klSjp/jupyfjiyDWuGAX1Fa
8RKpuUy41j3aCe7S/HBLyzFCgS7cCt6kc7gc+CfJrP1z0es5tGAQ7Cub7knY
0ZAzuX8WzICeLMlL6wlwGDj9eUqD3B4vI1M2cRT8rR9ipVFo90m+IRRSFWMc
EnrcByQM9tvu9dXaoq4vpcZLYjBEdTAPDSIN6DAD8sBkld7or/fOwbs1STCK
xJUD1XgewzVT3EJ0uAUuvPjf7YoU7YJ5/EE7XA4xdUsMyZU2etTd6u8L+m/x
FEUBkcdH8Dp47zPjIV3L1YmuPcuT01YeAkahOnne5uyR8k44c8eyTiZkXMVk
KVxSCUWzQQ/dndCGnOltiDTz4LX+ipxEWU9QglJLGwdB5AUGetwvHw92/z9J
7736yECrLIB1NZ9rmOD44CC/XI8m8RK3A1aibCqVu34KwpUqwYzrk88nFzsc
lSA4hDD3PNwnyLCb8Ek4sHLWv3uGsq4UuN3YD2QLUwqNeyXWdF+U3h3k2YIx
sAoo5vzZ0EbDOD5pB9EfUcvdHwRdH1aRFbrs3X7yUD3FqryaPseCnSKuMhwL
Gp1ou5WdGT3uQGTRB1Ph7Juy+9f55HA0Xw+d5pfv1sHZ7uLyytVIBHpEpBD5
PiizNOCOhbF9tKpVIZ3DK0+A4aCmZKA9TvhMU9PP8zVW4uRX1gE9uLpnbHQG
KW6ayD8mQdIM/gCBqgJSnEfW6yu9XsIpTu0tPpZR+nhS22kfLqe7ZwptCRwa
/gN8hBd3/l2fMajaU/AybpXqPH2L+RNAoZthtMZ7A7nl74ooYfNgRK7k2esi
7vRZPB+NJ5jZnHT83zS2NYDuZIhkfwwNZsD6uV0LgMkiMWo0MdpdEYGAQoar
BhAViQTrohtiU/3E1+c+usKFNitMrxGy4ib0Y6sgYc//FNDOHLJNqoWpjxmR
kLfA+ZGI4i56+EmQ57RF4dc+uYtx9ipuMiw7iSJG2dt4kD8/c+ZmVDiVYu9D
QzOdcf4C6RdFZ5bvzKBs+Nd2qEwAJJKJL7dx5Lf2wajMUErFqw5LWiCn2rfU
TLYwxjD2VE8QrkhPZP1IeBj3gs27V/JqJfNb0uGy/tlS9AG6sg4OGEvfnLML
po/XwY6MfePc1bI2mz2tiZOscDCRzqaA1JlKuSun/ahMfhGQmK7HKT9fgTUV
TwjQYbzgeYBhVOOyDjAkvDY5CDVHmqkk3+CzaznoxyZmI98T2D9faK3JIsSN
QSlnOp3NnO5gU586WoaqtLNhwd0bZPcmNQHLrlP3pOMw/e4kJ9JKL7lZEKHP
zTcuD4JZVAI3j11Kd3VAndA9PAFF2LDqE5fTJ20Y3R32i9YMWpXdvqA8UC0A
QGesML+PDG3g47b09p4YD+iO1LOYAHVf9CBvHMNxNoz3c8kwpBZlCFQdpxc6
WeGXQGgXL0hFWXNLk606BdC13b+vkf4TJIGanZy3LOv5WyRO0KAWSo7ZVxQ/
u1zWau1meqM7GZOpXNm4Avg8HzzrJynF7uGbhHwCdUel1qeAabIrGsNiRED8
BnUomy06nFAfe6Qkd9IZ+LnDTq7k8mieYoWLJOYxCTK99YLODPULWZ9yB1KM
pBxDgQz+liTz9DSe3r403dFikvEzdN6mXqbO0FvwNWnaihY3Oq6kX/BnPmMj
0bZfyiEByS8IPtMO9KcMjrcbldjEjSVsOwAS90yXuEHj0gVO7vBysUg17CxX
KE/15WdKpPTDPgCX+cPNmxxse7kz4nhzWCxDhfp0z9ChGo+JOiBMoKYwxzeo
lrYJp6pI0bpPa/o/7F4UYvr9VDhF66ZAZd9C6nukzVb9YxoagOA0A8N619Jd
LSLC/WCxx/KxpAS9JTqzODHWFzWLQme7v5HyG52yXdDfDVBXowxkTB/jUPkZ
HtQs4sZpoaoUW3W49tJllB0V/NBVXFa+MN4RK2nv8Z7TjvEj4jaxAYSWEz2J
2ylnDKRHO3YUkY+J1LhUc2mptZE/szYmeW8wJWuzrTe1h1ePh2vAHHHNm4+y
UI1/qACxWwLtsh+yBXdzRIbSvWV/wmNsVClZ7DkZeb66ghZeBUJqgPD1lMtW
/jbD0V7WKNf0DL6cuiMPAPWQ60tgjvv6KPrn+8m+BMSW8ZhRqyzrQqw7sKna
XweDuONhTVPPRoS6AH+obHsBuiyMP7GsKzarrEa0jTDLkq0qvhjAVhr1MQzv
gr71//orzqBUBzCKZrJPPC1jsZY7FIUR7xPuTmoyCohGOediLm9fZ6+ZMWL9
A9SqDbQ5QeHC4fIM0SyedTa1WUP6EF23blvRveSMEiF5+mifVQAvQ35as8xb
OwcDKXnuon+1RhLaZdVjb+oK+KD5j7C/0Br0wH6TWEXWZaSQbADfYe82+SsC
jhCyndFNMAdOHoR6q6/nOJP561CMtCevC2S15p7+sJqryQe0gqpEfuPDPhnX
PyvN1TbNXsZiUZ29qkojCw8XAtSvBq+qhmhGIKU9m5igcDtR5sCcS/3DSCwe
ELFTyraM5Yt/mWSE+o2V68vkd24udQY4dCb+pF1J4Essw37mNmEuhCadvazs
3c1oIgd+dbYdgecZikZMRLYZgd8lXZ8Yl9dUtwzTgyzKb9TRA96IoBX9yEju
biFILauDtDBETkPWqr4YcCJJKd0PI1VmTwpWSbGUZV+gmJMi4UqXpXU38r0K
i5/JZuUDKK2GSj6wO/74LMCPayvQnjyDK2RpYaNCa0ThHNWfWSfMMwepCsX4
OJHMwVoBH3hsrojBEMhKvFDCBWpYeJqsHdrB9A0Yz0mH6qtou4z5MOwnNYM3
r9S4WwP4soDygasr+FRLO12YDbfi/TE5wQN5PdWY47dE9qkHt2MqdIs4/fHO
PfucOHM9NwuEzERPrEC9mjhxC2Py5290nG64DsaHhBgWA49O0cxSTDrGBiKM
vua5eirjBC38D/kJYiVxS3vbK6/JRaPImmXguL8Ikb0BgCyN2XGF3M2gzWOP
IUu0b74DO0t0loD+Hfa+lwcs77ooaJ1/WtDFHZJL2GUHIStSSYNTN2XLJWIF
Qt6KCa43hOc7BYK7X5rvFW2ZIsaBH9s9P9NCclGj/I3gM+DqjgZyHOrsKpyA
ED0GXaAJt6UKi9jMNRaSInHCqJtnx1zlFzcDZDxjf7kiy/FJo6btfioNf0jo
j9IpPlxEfim06P+OkKDzehfjE7kI/7SvdNI/2qW1rmk7l/no2AQHs1I/PA0d
RGwKEYT7uiL4MR16pRq0k/eN82xJRMbOEKvNaAOpP6q7MrEyUr7tzthkEalw
oaHPa9TIgxEDDuEIPOVqE/T99L9ufACkIbpf+s6ewd/vd72kI+3j+LZdWYwD
o3T8uZzP9VEQGCmvy0/Q+ke2quYmFGzWNvf6jeBq2cQ/Dru8f7mL/aSPL92s
GFRggIwdz0JRIN8YC/l8L9BjBdD2jiBvepKP+EJT9LeIuCwrHAt6U9l0q8rf
CU2/K4q2N7CPD8FW5bnn+eybVA1IgYVPG94QYcODiap5ES2Gs31RonCoFQtU
6uNZU+ftKQ0cHVfvLIy21Pbto+Dv5spXV6yS6QOkNVenvCxsaQ3NUY7MD3Ek
M15Q7id+Cpml/YGsk5+nwjcsNQgeYcynCV5Z/gSBYbajoQ83/wXRVWkhV1mK
cTBD6Lf0NCB5xcPWFoM1EaUCYPFxbvpVKCcw9S+4eBvnjwS3jyXES5iOqaBi
NaGX75RfHNXImkaUeS63KPw0XCBW2LJXaMmLyDFf45zdTwLZn6PbWbeB5wDd
B8R/oVie91BvX8ALffbmP/t4tQ2daZx9XwPqSdwzeNRXQQDT8VhJ965yO1oL
mfdIs+b+1ezaGqCCLaZudG2lJ6KyFszpowVMut9Ie0qgNoonpPC3/pPA+0eH
daVBHmZsekgK8pcUN2wGhU4Bam83w7Nxzn6E/URe/1YDBNWO2H6j7IwEBhur
lqFnx4uOymYH18v38PAyJlPPv8Q8gIEeF8PqStVFO2NaKHeaLzKjCAMRlEDV
LYBZRkgTDcMXN97epOuAdBrVstqH3xVpazxaGgd8RrqtX1EpiUo8sguXgejm
kTPcn2DGJqo/BRfOFqDMVqs6zfARIo2YhYBZJxvJCKvBoPyc/x5+1O8/bs8I
vKza2cM85itGkXKS6chJZRZq0m1hCZHa3RUQaVuekWs0zJQh0nYuoVBm06aV
jG3KPKcoqITC7PEp41FpMN/AUX8gyoF2yfoIg+dNplXXU3C/h9yLtyhx9JDM
UYLyqVTCNjQOwVwRoKlwDSqiJRVvYD8HFH2m8z377KSeb33k6PGRptzuOdgf
QznLKCJZoDn2nJn7+ULPFnlE7mVVGgVfQcQVQkRcuNyL9opoY0qDxgQ+Emp6
LY8h1iURyoWl63w6hCBCBhvDRA5YbndbU9TVjT68Xc5X4kXe0zaM4zs1cxWS
QCJJF55pDHtKMf15E45+bFov2l4T1okvK7O06PbCnpMcS1V/shTyyEzEm3Z+
+EzaVL0+sWC04gQ0ZHxo8Xkus+HpH6QUqt1hn50CtM5go5gFfusK8zBNaqkC
OD3RRFKoZBnFh7ivpZdGk9JNMcjGwfGIjwwsAo2/d0JgtdykoFzpSkuqazD5
iNXy+RMRCL++znqAExWEn7kV4UXiPVVBsuv95LQ3oC7KUgKRZzM2Xy1FemV4
RScaKqWfdlZCYnUiBz7lhTeO9q2n2/1+wqEcuteDPK5U5p1YnUdIOpQ1QMu1
sV+DYygR9HcCokMhuuBfIb/lCku7DE3Fc64y5p8A/Uzf68ZPPDubl4ZDaADa
WcZ/KAcLir3p+Su8V5B93sPEQqSy1gu36tLrw3w4LQG9t5h+qWyJ3heWxh8c
FateZcHelBlzZAOpnGMIq85OVE5BEb5UuO1lZsxNm0jrc+LplD3l2TC+CxdU
vLGCG2CYPIZ4S9O5SCGnlS/LasUMD2CN3hVuO5IYuMjz95NhdPG6rYPyEpmN
ya+pD1w8hW2AHXRi1/vGuGQxdbEmIt5sQ4ArYq/TAHdpUykuOZeCRyDAk2QK
Xt2BMeD1q/jLzVb2vvudNPgn6ZMNHEwzpaOMGF4EAubZI8g1NwQj3JMF7HDZ
FWMO07pMknrVagNCZBf1nfShti0yV7vXstOPpEBBHqdVOb5WZ2DJHDJ1D38e
UPyJnHezyeNWKgxQ3Dq4SqquHaXYOcclE7AZ/CLmIBMh+yIX7csT82rcFbvC
hLg1LMXkPewhG6zjmGymzFhMp8fiAG0pl8ako01fG9nG/ls+LtJGyOca3u5R
jfz7ZpDR0m2S8JRa422L6WdqMnDVw3CyVfANq+SrY0+WtlHWU0R3piRA2hOT
mnvgaBlacF5fXMWZncBkHIdS23T3NTXAMEzxiVKF0LL+1+cJ/Gg9JauK5mt5
6hvVQBQXTr52ux3y9GWPaQ9GEh0b2rwNaitdjUJQGjvzCU26D+DBQ5DB3+n6
Np7xEpHu2odFhcQsdEHvlk4jlCDYtDivk9hIa04oEHr3ppGMdyVYJByaZttF
B8JaEE/HzY38Ufxz2Mbg4rrGDL5aZzKguQkgdPezos3mIqtJ5LJ/dHj/Q4Di
2GWAiHQAvTSOnRdFAa8zQ9dQ3Ndit9QqmNMx2X44uvfq1RLN96drTr5Alt4O
WtHUeM6gkP911eIaPxFI/6fj7t9qm8t4WgpfxG9IBmc120V+68nVifKa2pgK
vh+jKEf3dJOCrz67AxNqbzxKFKKD5o+Jdta0PMxpjLR+Ddn6wj7CokAx6/QM
kRibhTQvir1QfI2jtUd77of2ZW8fognamSNfANH5fAuXuOsyPrOKqmLt2NQR
Sz0SW+xjQFPY51WB2tsFWbbGSyLd12pHoade0GuM0DMBSehTlxZff666PSZi
FSJH69FgC4pF4Be1oDVP8IR41OpphAwM1gUsIRCqzY8i+fe7E6MZJ9oltI6s
9uWRsOK/IWXDOd7iHsypUsQbFcnmkNXmOQKfQ9FFaPdX8vYthW1oFlQTrOwk
ObkFjNcobaVbzK3H5jhVrShoXE635QEb384c+YRnTSxTmQgqOx58ep+T65+z
hnOCayLMoOtkcYuIvq/lygPnbzKDulruFnEQpLI87pN6D6VeuJ9cWXYxXSkt
tFZC8w1Vl301poMyXDGGQxhdxPo63SvwmP8xNUlPvJnv2zs3bSeZ070VBy3y
O7EgNXpokhAkvoknuXxEWryCTXIjxinfTJvtY3l+9kWpHQAVMdV6TuZp0r5h
7Qia8GI9lHCyvI0+e6C8zEB3t9pWYKpz3M4gZeNEKLedUNB9ccHJ8Jb/oQBA
V92VQ0+3fzCMeinc7koZvTiFmwcRJSEHqzeYxoegqvFKXEPNu1nd3VuP4PRo
CqSJ0IfSpX3lYrZNU/Mji+8QYq4onprtCeP+UkEEfLF2fDqB/JcA7CDD1Q3E
tJ86BMgVdZpty51SHxT41ULHL6aAu1WlWF//pj9CHfn8dE3mkTgCwBbzYcns
2gQQRZBhpgzyL0JwTO82NSoEOxU3PoBbYBMB07pjNgs8zOwPhNyZGMrPUKyM
aCwHVjPiUwaoDtrN0AE6H16j4fR7QXKHgwR+9/cViblyZ6eUucPBYnJd4KUN
YiBw/Ndfi+WRwL/P/2F8JEN1k0k8z11ldOZV88xMw6SNdVtvb+9uRtPEWUb3
ws70fcYWohmP2CQ2aNXSbvdZtJYeMcnMXWR1I8puDS5NY1/mOho+BjwKhG5S
euBQbB0fp/IkAZViaKhSfkVFIuTJnhzHtFDYxOP3tOQR/LU5mLZOclD3gWxh
fe1wLrS5NFmbsfRKl5TTt1/xGq8f8dtN2YVeIx+oUUrYccTbNoQ1qQjcOL7o
9FAa9DMD0Tm2AqsTh6pL/c0xQxng6y21njOQYHzmvz6pHCaRDgj9uXqMxFHQ
/Lo7apk+CQVKJujW/ZnN0XuN9g60HFvySYGD9hIlTHXdL7Yj9eoB6P6ejlUS
wvpwWKbfHTg8Oi5rOuxUVeECwVk4nxrQWRW8gBFKAd0bUXpp2aUOx3f4xWK1
0sAoUpnZPfbopNAfkLCQ9jTLgcymVnq3kHtksMuxK92OqQn12uQGXxLQxgHT
T2vVfkqlePEQczjzgAi0wiC4Cwxb03gIxRM8gH24I3Q2bPahAfyY5iEk/1Zh
tyNMmLk9QumYrvDuoRoj96PyJuyAaWDNY6RShXpTF1d7xP/sto3yl7f8nOUO
mFyhsjnq44w1cUBd465mUzoLUHI/YkJV7Z6cPY4XVGM2vNwJFVUiDkh+6EUk
XOPQbA1UJHuOUjvkdCaXWjy3u0fRbfb/eT+em/K0K6IPnQhiD6V8liLie0n2
KyROvQMedKX+CXVI8wWemcUrj0hy1UPVRMNpOO/OF+sEk02tdP4qvV+cOGXV
oD0awJbY0mIaVZmj89qY1tCemTGYPSioPHa59tza29rrQNg5q5D399gWEZGI
VuTQHhj6EaT8Yhf5+3yI88/Xk1Z9xI4k2ZYmC/Ha0IXcsPB7kmqU+/oyb1ML
EfXs02Otg0Y87CiBvOWIZfuko9p4bnkE2cpzJSBji+zD89y3Ct6GZHupyzQx
rC1e6KYlpt+vqtoNsveY2u6UQWQH9SM8FEV0ui/Xlvln98HANVkQXksv0vJ9
kERU1+Y/TRLehFFIHBVfHfro0Gy5f6auB8ydhv0J5g2d1DClatA3qZy0DWPp
2ovZWex7rXFYrINAf7pAteiS3aJoMTExfKJIbQDPZnAMFxRv6O5KH03MgdNE
Ef1yNwvnN0qyKYQsdeYKhjejoi+9f6TG94wTWhUViZCpUk/mAMaa7YfeMzpE
3DCcuZj6fW5mtOGstk6hYiOFiAYEriSp3abkRWZEf9gtmBWPO+AaXoJI5jbl
HPUgysOU7otb22h4R1k90VoiknSU1bnIx8meTxsuU/WFHm/nlNXhn6oo3T4l
c5coL1pJOK69gwq5roFQKTkgqbt2fa9jXi4MUeQN/ufAIYpfj7eDtnlETyUd
TKsMS2QNNjcYvhdM0lDsvHnxWICAftPb+Pgm4BOzreF+4msWvfqnmLSBvAoU
jx9JTdCby1OGCPMVLUiqOmnhqQFoTTmZ1Oy77lLqw0qHCU66aTQliDtIc8BE
7XVJVLmt4nfjSNXCqNZi0A3jllMp0gE7pMV/6B4OxJO9NlaGar+BLqYxR8lG
6BdOUA1I/slhdB51nC2MhPXAVpFu3fsV8YjLCg3TyLg7Zmq15Wa7sZm01eAF
R9Asq9uDc7uqg2563sB2+UaXbQh2W1FqneLLWAma+b5Ev5WPVG3G2XEMOO9o
VzjUHd1vUZ7AFLbP67aB1ylOuzQyXEVbmNPokvJA1wq8JCVyG/kPCzTSuZ8w
AA7/BQsedtiugVN2M9anyrbtzhvP5cX2Dog9rVl3OddHyMdKruja22vR0T5C
m7Iicxjc57YnQzSxUz/ZqlX9qgPMScfPo5wVd79jWKx5+zRp9sPcEYBBhmPW
jZDAwQ7w2wYd/Dfb4JtL3KDg1rwa7zasuHf3dUQLekYzZnBXqiiFutVR14fO
fMh6rX4fLTXFRjkw/oimplV6Z1VD4hmOp3vufSb+rhayLfV07mT3cCdzFhOT
p42Fc2YZb1e+Eq/Yxu7IgLB6KZbF6Ado7UNlJnoKqmSJ2j5NtlBLI61miF23
kPuHtVkO9G0k1s3BEjXD6QisdubCulc3E9mNJt5Trg5NwTKfuFwBS9EYhpNX
WcfxahuNsX23Hu8cW+9Ez1F1vN0ooyw5i3BSpezFe7JGtHT4i+fxNAA6ku/N
6Q7vxtQip2r5qL38QLux8I6NlRkC5GYI9vsOaRQR6eFrCuBPY+/nx8+VlyoQ
CPa5s9Zg2NBGz3GkEMQrww/7L149ugOGnYUd0scz3FXYku/MVuGpt+PesEy9
gqZ6ZV0hlu8EfiI+ovvTaE+Y3Xksqa/XOeJLwBoUdDUKQmuoujn0aDHDeHqR
m5UaYxwz8WOZEU8BJ7L8jPLUJCoufr2Tv0hW0aetkqKZuQVEVl7zFUrq5xAN
u9mvFrOXVIFPGU/9smbtyjQ1O2SpBmCnJaFJzELnBDENreqM8X1om67/nKTt
i4S/GYHoP0lmIbY5BJ0JXFyiFnPCMbmpxG2uUKNSJ3Gyfu+kz3qDjqnuB0Us
sg54kNvmIk/BBqmunbfQmE/sIEqv9VhfgRDX+0y8NiKORxoqwmacbsAdQ9Fo
/SjT3DA8exJc0X0d6iZ66pMBdXkLNjY+m3x7/03n9fKrl8+3O3Ntsf81h8CU
NseCLemXY7iTzz1HRaaeB8aDBjSR9uBsuPRiAp4RhH8U4/qYzdWO0/yBTtta
1XCovf8W8xzZcSbX3Oz5sIvqW89Ez+Q2B3CXPqiuqiXmoqPYynIr10hrPg+s
ID3BUgVldIb1AQ3/RHOODZOqZK4u4G82ZbIqGs7UftOQyuP5q+cooRfSRdI9
RrMuv1DI6VUOszym4v+pvoDfy0yutVCTSv3gWA87YGlsqth2F6XWusSjQWp4
KHZRAZLHqEhx22K6Fq67R3RBkIJZw17wfXfmYN3D4i5PeW2NWeY1Xtbf8Bdo
b3/G0ROFPQCv5Kkh0qtgIfQKYACnMJmEH/ao0QMq6Qm4Dh3VFUVAhK21Dn+h
9VQUKScldH+bu2pPvsGjkZkGdaML1XO/vuHKQf2shjNA8f5clWjHg92jIzN6
/R9EwJ78mTVtgGyi8wl1q1abMa9lnXFi1HQ5RfNcMQgsRCDetHVaqY8SkxLV
u4s/4ayhJmvLYWs32PJViEKX6HJFiA7cy7+A3ns0EAP4xYwf7z1Q+7+EIM6G
I/cggcIN6a24TBUXFfuC00VqG4wMLwNINTAiwbmohcCgWIQ4Hm6PcWaTmtje
a5hJngTdVNZpyuXvXXyP/3HOeRPDahT9RjiVkLtTfmHVspdsiTUFpxCkWUnU
h2zyFJMiHZt5Ia2rOBb+VvrnAgKPz5PUA/r/jAmgo0FLS3I0dhc8/qrqhICS
pX9z+j+phzcwubGh7umt1l011f8KZ9N3SuRIaCHMdg9IwTZ8chp7Kwl3cpxd
S5LNDXWb257XFvaOPcFGL/z+C1la41edhRYe7cCHmZ306+mkWOZcMICo2guX
O1dNI4mM9on2iZlyTvw+dHOdTEGzEk7TP48fkBSm80R73QPiY25qF6cOLmyF
tgsNSQd8R0EuSMET12vWJzMJAT1nynhLQLm4ZTEg6Q5KK17+zM8RkeRW+fY1
sVT8OzhrwFhRAjEdyO6/5NkhIgkP6gGMPFk+svX6iA24CM0UlReVPyHlJNqX
Jtpo70Q6WZIRs9XyP7VygoX2PC921ORTeOBBlFvVSOJxAG/a0Br533wuHdJ+
smUfR5NPq0Nk5trshoyOsp56YiDX74tBHT/40YqIqbYMKFXxSHBG3P0VfGHJ
M3xmIYAHq8eQKhYle0UWBHG/kQ6ExnrYi6QH+ev2zS2A8etkMl7Ul6tjJh5u
k3TTG62vqe8nmcZMKZzeksYJzEMI/WD4EpxtfD4AA4t2kS4CAnt80bSgJe5d
QVMmE7HP/Dg+Au2HSyZM6egdVegr8RsS6lJsUztHamdOiGk6FVXJ2RZBSgt5
2tUBkaLKBzmupT74BY95vV5D1Iv0a4QjNQgAEWAvReRy7sIRiHrwL/T2bjyi
wNA9zd3RrDjf5AdcKxSu+h42kyFRpNZeEFqJiiQgcJg/D0EELdr/zsQGmBNW
Bak4pLMp6nPlzruVYIxcfMVK1NwMixztsDTBvGKeQYwYSZGTnBmbU6bUJ/Y/
h/lMYEsJ4dTppqHIvFuQhh1w4pj120tDjelU5POYjjPYHeivYbqR4C7PKe10
lO/69yJQUR3nA/6UM/jjz1KwhYnyVb1ixlEqYHvMSzQ4mMKGOYiPImBEkoYH
iwa4F9sMFs4nti/R4HNKxy2CR036FBL0ZGVy6sh7DZeXzo5PNh9UYrgfIGQx
wOHrH/Q8Vn22FV1evoPz3tJLCa6ZTrYk7w+z6Uql3GV1xXCpBJI4+TEOJgE2
CED1vMqOxzlMRZmV0SZIqEE89KnMVAMsO09nOCpGnBIjhrJYf3qPbgwzgJ4p
DX1+DzgsO8KMvRc97o1w2/cR9H26NbO0Nny8rlz2rFmwmvh6ZrQFkMKPhj4F
tHNzF3K+yLKi8afLKAVyoDEPFZSVxZ9xT0uIgX8sFxuOVW3x8G7a6lSC6j2I
zztlfE3rVuWDsxgsgmcchjFJNTYf+LG6EPn4ByLhAFGtIj4Pq3xNdrP20tdj
XfgPhuQ+wygyXeAPIOIz7BTwu3pMETpL8vZuLhpEw1ca3fDcJm4OOSEFDecT
OATBs3ugUvHd5m/eXbrhoSVypJekb60hBOVl+DmOB6Pgb/3Im55NzDEoxtz8
GcvnHSZDY1psfjyvGDLPql8xOIYpZXvEZwynRuALxC5UCgCXNjSqOAiV6/dT
/C4T9Vla/BpTqHb4K1FdSvPd0P7MttJjg+yAzvkI73FMi9DRn9OwCK2nPyql
f4njFLoV8C+48IFoSLfpLqQY5H8RKWre8EeTviY3e1/u1wJhzSDgItCXKFxj
8YrqHGcHJuZzPHSCt4KnBDTWAurV+/2W18Sz6a83W05xhZgE7gnwHFwcBzsk
UfbjkStPXlVxRAC58y59J8FdLcSdL3ZzYIcKV23vnF0zrzzZjPgJRZUm2TqO
4UrCWI7Y3qpQE1iizjnxh4SK6YENHYgFqNfJU9qCkw/Rsm1zD/q1igdq08b9
6w4N3a2Bzi/pbR30MHq7Nvfx0PGwAa4CYmK93kB7wZMg+F5NGNrn3uw20gRR
3C1NzqF1oEFuOuNgpTzJ9kymcC50c0FIRMsKe/D53fRLfHrUcUJeMRRaxV9C
Orkw1P3wEwSDtYmlYnWWCsI+A+iQmkDWCAg0CkZDXpJQh8r4vMPDKr/1sa1W
OkkSO809r8MKuqRayoUMeLMjRLQKfR19fvr1M6j7hAdjTtdk11O1tIFCH49D
WqcrP7d9P/CjnVJcE0fyYQiR6e5r+zMdUgl/ml2OLm3z2SS1tXi07VwVcRKI
fEZbpPcOa4efKC2yAnOiv+aeLYZiMHY0P+PBy0qZuVqk4T4dXk+zQHvZbmIB
1aGIbbYlh8jqp5MEEzEvsq5AU7l4jLXnJSsas5m87NTLfIiPJwUmE4Qy++5e
l6fNZ5w1PPZjbc3H/q/rxMluc8FnyoHZvHaEF/5vkDD+WM3Yefzzwy2kiqGg
gdmLZCcaszJ/zXnIjB0JtDipOQHfJJncj1yTx7G9O9jnfCHAVK5hha7a0X8y
8o6qhbzDmSIoJ7/0YPixQe3lUn0CEVWCEJ2qqfyrwgxQPpV+65er/JUDEeQ8
ZwLhLl+SPvkgsGO5GVxJd9/ir2iRuxhuKm9wJbDMFo2wqTrfQpeHXCquv9pV
dWHusdKOhbVf4UW3pufzfllDAoGuHhRumkdq84FzF0agKgAlo/WViKAOJ5ww
7Y1B1eo3p4zKGIKu5tup6gHhCvGY086TcFcRcwkogfE5RJ2/izedjovZa+0g
3TM8KvKBri03P3oG9EOZFRpJtLb/IGoyZWi1G4fG/zCENmdpl/X3/j5f8lwe
gwTchgcek8rJONorbjYgmFFsu30NxUb4rswrBTlWptXkXbx+ccOa7vKILWI+
AGT4Yr8lyWvWD6xA7rjSfPozpscnPZwNQUP4AFxosQ9gRL6MNfoItlFddkBN
jEf3CUXoCd/nwNuoRAfbaSKf77DjaH1fJN7rbWrpSvgQWPmYN9+907n0TS/t
9DMcrlbxYo0tD2g3mXhsF/PYV4f9vLDdpbshHEinZhxz0clUi+v9eM14jZHU
DJC1NNLTEfJ1BKZYhjT130z7zG9QEFUa4jJqs8rxAjTExCV4vhA+XhE0XfoC
4sLhbE4yXTVbvmrzGeBo/PCfYWQB+8tcKTQ7POa+NfrwGGwtDin8ktzhxIVj
OVAFSxMquhq7uFnTiWfEpDIucI8QZMdPBSa1/7G5dzixt88xo/+TZlJ5JKad
uK9zh88ZO7GoHXszs7ljlxMZI5IqibRdg4Sp5EZ9GWYkxDpYABj7F93+OdJ+
KfRmzXJiOWrQqIF2BzTOzwpNKzg5gvV1tABaK3AMOMLqQCLW/8r0JN0wBE9f
jgkE5B4CbJcMycx93FrdPEcmcXIyyMZ3gfEbyOzkyIXw5+35pTcnlkYOcRr4
Zc7yAdfrxPjK5EpIZmGB7M6PwavKkCxMbSsHwdeylp7W+lWjpZtiIlX+QISZ
tNwDINSScetMPLfq2MxvOej/h7pYD1PA1vB5lk8Ul4y6NW1Dd063CbrJXiBd
SecZgw+oVZ+oQKlwv4asGHaYL/EsIuoIRaPR3/BO0CdYxWfaV4SjE5Db59Ec
huNo9vCILlniP49XBDNuVFDa6YNdBNj2XuRPGnzxvDdoPMeZrAn+n9si+y6R
GXgXqSw++01RzU50/p5frRqpLWM4W37FopEPtcrSkTQpgnLlMXXyWa49tsY9
4JD5SV+NGH0y4088z1iht9IalWyCMBL1Bi0hk4OkODjCTHI1CVZX2yr92YGD
vaGUe9iKgNlWgJWHT9CJpR3U1u6ZHrgK2jKeDlemFgHwWoz7KIZm/u00gO0z
Ma/DhNK7zngCX1mTML4ZZUMSScTJTjBQ7y392RBw/ojk8c99pOV4d517/+Vk
l8HGlUlAG9QUYKu5pyd3mhK8bnJHQfiXai9+sznxg2fZWmOKnxvgNpviHdUp
aD6TFhmW80fAz406TKvg/fD9WIFi6+irc10zYvcGylmCT+Wql7tLOeYV8pZd
7q51ExZPBaLftBiYNeweOoLFCuiQPXp4exVLWDOI+1mKTwCM85sEXlCV7DlS
EEYpBIXpLntyPBJXfcG8n4UFCYbBOnDA9cRtsYPOYjuKe3GIGP0aXyG491Gl
MjZQ0nz9fIndbQm9vMHZEZ8KqN7Z9ZFx2cJixY6DB1X4Vf5u5rORS4AhZxeN
vU5hDrEdgo1ZeTO92CTsgrAFDtJveya9zMuewy1vzLaENEcwpM4f9u9LbZct
npOUCu91FIAIuZwoVFvdHYff+Sz8RW3o9Mlxh+Bq5lcDW8JB68nDGs732CCV
+SO747KppwXNm1kKVEQSFL+xenrIYmfMOTVeo55a8YjjRxdY9GW3OlXfvy9T
GB3PlJVxRoxv8xsXp91P2rc6iUFECkj08RNi6HpiIFOko8QIAZJ7Uvxlkroj
YT00VnMnozSTIvuUvhUTkiV8/RppScUVgQC4McvmIVva59CuNlNbjaOaiA0n
J4qiT/8MyLK3K7IusVAIs9DfNURKQ5xEJlblXBiOUcxZmD+Z7AWADuZFhvAS
M4xHD6cGrisrokm+4+j3ytsSq4BmtH7hd0G2aZ5WJVCqv5tp/nLhwMVIDg53
wGkFMJg3cMgdO6g0RnOZ8wicGz+k8pvOWgUVoWk2YIssXpiVGur1eb02iD3U
60f0SGZoThsXw4BD/PPwNojbs805AeoDhzy+97RMZTKoTAxBjOunwW80n2Oz
bCoUfWqQ7c11E/siM3YFExV2J4bWFjAxOHE6u2r918BmcXUN2zun4jB0nLSH
MqFF9CXHsaBRfyIuQeE5iflP3HTs8hRD17kg9OsVWxu8hHBP6CBgrevLvafl
73dTWBPG7JY5ThzZDfwDhZNGIqYUusgY/TScXgw4q0WhlVRgmEYEDUtz59kd
D2hTNWwBPbVuo5ZTsCeEQ8H4dv/SmMGkPyUUhoFtdhcTp71qe3B3iW6iM/Sh
umlZAVq/iZwYNmjtIww92+HLei1MYXRzhHZmJG9s1XFLua923+xC27uUsTyI
cPev5FUqYwaHrl6dbauu7br+dI+LPPCoAZVKkuqmdG0fhdizqnl/O3EKFarn
/qgCaiPWBYlzk5bkVzto1Y5ypCpTvhmuPb9fO6S6c8qnRxTTwvFYq3xMAzwv
uppzPt6koeCbHh9J/Oc+VDZCRxf9LXrnEhal/a6yAgxRubLbVkzmwl3Qv+nr
7oy8pqDeNy4RIeKzvkapMFTGqxWjRTITkzB+W7k31aldCzOqsrlEkgwNe1Nt
RhtXJqL/b1E6x4Nz5EiJdqWlkL4eHvqByOUa7go2S06yHDFoA61C/ZFaxbOW
i/Bb8YqkA21481La0/uG4PVZbjwD3Bf5d7TBpzhmSfPeAQotuihRCHzo4xHJ
65cj6xLjr6dZxbZhW3TwsOITwKAcI9/9Gdy989B9xG1OVTjd2HBiBx7OUp52
FuTyCFZOYYRuEaxdSGEPFlFmIOHE8rlUsTcqyVfVU3Fs+u6vomVkc15d11Is
y4gDVcalo8WT164WQFMk5mDErx1VH1CtIaY4BppnGE0kzsTwH7a/f/6f57Wa
L7xI20e4OPmYpxPWj5kgR/meQvcw8MuU/+Ph0i3/7qJFZBYLTCfZJDFt4UNT
SDPJLSrcgJMhe/YVaC8s7DotELlQSE9QlIk3McP0zmL2rz89lfx7B/BY7PWt
qjRUuL+SAqO6cXu/aaXsUFiB+x7O9d0xbuz20ZeLhNUUN+khMprqjdzgAS8R
+d6KrLeM6vnF+E5ptGPweKyv85S0ZQ/cUArpmB96rWd6dGJkHqQ6axK5x9X8
JAJ2S+VpIwdw/uemAFiI1ETmPyr1jeItru1djdH8KIOfZRs7iAouNUNF1PHd
yPD58k8yXq/9c3qw/nLqbh70YGmiJZqThTeLb3ugo7jgWbbcD9OgUqKsLH2q
bQ738QP6Jk4oSWoIZTkv0NcFchK13UepU/DHvdi4ktojw7j7xWJhep8vFavL
Flqxb+l9mVn2qPGfPdxnXh4YxroLulJEWoBkA68cEsoOCAXXCM46k4VwBRoj
ZItEp7rrwc6SFl4gaNmshkbUT0mYucJAOeJBAQLhecHBNu1KkQsXSqsOlzDY
4KPBEZzUKltVfzUskAJKUhNCpOg1FqfsB9cfyIN8iffVWXUMO15wUIesuqDp
FGGaaVFhT3fzsszup6ni08FuuDDCFAMwwqMgZb+cueOXs/ugy4CTIw+pp91+
SQX3TgTlRNaFmEsAs91+INUfVE++Nr8HMTsxXHwUI4Pyso4mDxxN9YCgQjKP
jM4g9YPv7k7S2HGuUIYIcJ/0ibCay9ub5ohD/xa85Q6iSI6ZpKbOLV4mTbV8
CP3438LmROolsOxo7xGmscssY/Rrhu7rbtGXx2Rl7ADe13CUcYg3+NmGX5GS
DkW3PZdw+w7iZxIm8jp84Mm299RvUfyyjJ8ReDGzvu1vhKwuolQb2fY9SOe8
DZleAkS12mUkESAvkZ9s0ugrzLd009z8dbiMQJyoBRsUp1LaRDtzaZRtYr+q
aWwsf4P+ap9Na/koRVOO93y0Zpbg2tixkqJwgOce7FJeea9EsNCHGsq113F2
OpdapzRoNlx8qHcEoIi/R/quAa7TKHyFkOX2EswkQakmq7t3hgJ2YPl7321w
XMf9+RNozScimTxmoZaulppQhPuyon6Jp1qDPmEPAApS4dlh3Vyw6Q4YG/ix
i0DtCL7HjONFLNT7mFcjeXF8C0EKjGLhCAJd85p+dDZ+GghmvqATp/47Hh0H
g91HIb4keYeuDldFQJoauzdS1MJS6wnV7yruyfb9iZDwv7wS/PM8ozcrn0Rz
dF4HOkwZtAjNYxEUXnOgzTIS07uqdxKgyx0ah5LudFj4gSmszf2lakqQET+N
//JK00BhNUQ2KipbAbz+ELhRgFJOUvIh0BJIRjSyVtIOtts9jHxYgQqfScxe
cwuV7i5z9876pWEHjjQ9RPG86qwmbqZlFb3wajktbx4Wzbwx+6MxRcjo+MLO
tTtaskoRepi+gMoPovvdE8ofwNWxKDIY1Fiy/Fg10BLAOcoo+fqGj2SJVpio
K7e2fglXP7VfOWKH7gA6XhGitie1ER/5XO0emA9dH+kWzB7qqDIqm3gVGPZ5
qB02e8umVu8ls0lTMkcLBQfmJ2pWXuRnaXAHVMV2ALFI3Fj3ml4u0RF4GWTs
z6lCf3ok1ZgjJKR9Jeb8eb30939ZQpuP0iTh3F0KSLVI63DzHeAMe+u7f2Lz
9UWkXI9/7+lXH3r2Nl6HDASoFdt4D/hyGk6UtS78Xidm4FLx8Hrc/MY2+rsI
YWUGLJjy+q3f+qfJa3AZucn2y/d8a7gyAhUNVkAfok8hFK3alnNwuv/ehGTF
M3onSEQb+g7rtpcKfxlPfV444sflbhH2WjM5vdkNS1Y5f00n/eWzZOUN6xAf
r+JPvJoeKZTVEM2OsaUn4bfFMlRd0cjmkQ4CimKDa5pL2dNlAXSwBQSL1EAZ
RcYlCwf6ukH+3yDLCjZ4UxX76FdGla75Nz5Ylaa8g3XinBXxLQZ1duOwaEvQ
fO0pCQWwsf5L6YASlvASfFizgaRMGn8O9iN9w1mV1wvR9yfGufFL6B82AZJR
Z/hbLAKIARKvrz2RsPEQAj+u4XmiYHix9pMLxNQhe9Wi8Te8hFIDC76H6JMO
KYEqect1+Q7dH9mrpubS5SxTeVkGmgfyqyiCPK47qo03r0o3roBA23BVeDNm
OlFb6Wtxc3OsGgzXkLqcJV51xQKj8fsY/5DHkSBQg3un7xV+4YFCy09FZdal
liiy/D3ZydUc973oZBO1ilD/34QLrobT4qAJH5WmsTrciSIwBg+fXdClN8XN
wfl1OvkIailtuxsl3Ov21n9GEB8xpj6gwsnLJ0H8A1GRa4FlEcMxuuSiWk9N
a5cGQwziFQAPzimjZ3thcpdx3O1DvwpFAvxBHtDrFRBu8RtL0ockteulI6/I
yLdZzE+SeASV/VDE2oBpjN1IR0zYXKLwIV+GhV/RVxOJ6603C4Ul3hUncHcn
nhzXxeeB6oD50c79weAxDBFDGpGla8ICGNiT+BF7t1bPBdm1b5CtyoHy92yn
VbH/CgHdJPMIN9ycp/XK8fyQHL9d7U86OIJ+F98k79+xG4gPRQNbZ8cEEHNJ
NLAIlxXi/l8ZD+gXV7vUkMf4r84dbPEmO24NUaxWp6uPJ00PDVGURee1ffFM
rtszZRGRu+0lDQfQPCfQyv9RMth9Q+/+j/9A6vtu8xlLSEPxJkN18zUvo8a8
BswD7yAoZ7f2NHUpU9i+d2eYohpTawsgCz/pHXb6GeDxjYE9AxfXFfnxuJZ5
f2aAbaTD515MXMWbRm57xD6QEOOymhbGYDGMUOn/4/5qGZxJ24TNmr+PXD4b
Q9lMWVu4yPMXrwFPaUDVQZjzfifclum4OlhHkshto4xNtZKRLrQJwh4ibvSP
SxLYT5d/k3Jgl5Yx85tx/JO82hIwHhSVy7sCFg43GbelMV0afuSTddGSEcqI
bzMOYzszMBrTNfZn2oInOyUaKYeElXIV1PzTWO0wezyISQrp0Ygf2bHJVFvT
kGu/V3rlKl+7huoYI1gZCNDV+QHcDG75RN2/XPEg7VFzS9UVWSgMRdnPmQ2R
FvhvMk+moN0LpGIqKdRWFayxaUCsWZ+SaJkHlqDSazalJhfA+el2AsD+6jl5
FZInj+OyW/s7uqfR8oSL37+b9R1Afccy9zuFgAJzRFMUut9Z+fImrac9kiGL
WaBjvANfB47C0i0OZOoTI0gyqY7gD6NR2+DysEYQsAylDhwqxdrJFnjc4C7E
rabZnfhETRcChS/b3qKjxcIZxWDX0rzh8gHE20KMjWkR8hRUiwAgjN/tnrsx
OEnZN+UFrXyCQ8jeLUsAklwID7WXEY15kPbtgC0tmBAowAQc3JdD2nouo/90
LPV35o9LlZdvIO7HRX5VctyR5typmvsnMATvRYUOXVA1Tqoe5ydgM5IeGP0i
S4ko9M+UUvwB92ovv9pRrtiwLIIhcgLnkHXNgfkHn0ekOgJUPyIDuijBts6/
ZexzjsLfDZd/dQxYp5GRt4cD+FiH+HZCIj97QqSoDqTNF2lN4qlmk6au95V0
ZYMu79Znuc/XW5t8hlghona2b62Ci8YSpVVAZr1HZgflfzb5xxyAwiwYO9wm
HUAvTq760NMCePSv5kJ8ZaBisHp9QuhS5qc3tXs0M4UsYNuC6o5mblU0YZSx
smXOjHOgFyh7p/EsMDPCASZ9B8H9cxNzT7yGDOBnmmlexiriXR6MdyL25CtV
4tomXEqCToslNqBD22l/huJrookVXS1aw4LkuL1j12NvVosuAD6RmimQ4k42
Fn5Z9eXNUNb7bY4D/ZtlWgE9Kwmx0AnrJL/eoDo4hddgb+bl0B8Kdr54k1Et
Vur36++vjIDamxEIxVT4FHC3pdx44YEhWuE2YeyPQbm2+mHIYAVOzCJE3huV
ThD0Q3jFjN3amYeOoJIoMQl21W9lCkV0uI1CpfLhW5rzdszfqBpA0pUvXIhD
IQkx4wX8QUWAqMwcByLe2HJsGYzkzGLe54hdbba6OZunzojM/+NCzfubi5Tw
Z7X/HjAdlxvxp31GOJrjnrgS0DVw5D/mwdbmJghx3XoHIAyc7sQGB9KCGhsP
DwGgnLtRHdpBZ4e17Y9N2LfCZAm2b1cRyqu0XTVTJK5b8uDstmQwN+SWYynF
5iw0aOCO350yN645MbACvgTMY4vUCGK2cm8ZOleJyPWs9CrwRZUHnba1qNeV
CB7ygsZxG9ABvmUn71XsBd5xiH1iGsPL8ro48jhXpzLIJcabehkBdinlPZMJ
ejKHbvpy6nDqP9xVWJFjqrdmxMY5MJdOZ8ifzGR+ymhJF/QAzVTpxjRaZll3
LCV5bQF8t/WOW2iddaDqorZhOGr7xhDFwpMUz4RMB49PMiSxyaAhNw+73BSS
8kq9lS61vCh8Ipz7Udfj8tpdIzETaz2u+hWkgJoBUmFtCQLfp7RGaICsh5y/
HYgzIgXgxPR0H40V7S9KvDUsGltcNckF2yDYA4ZzJlQUNsHjEn5cjFupXOot
U5laOoWte/fI9LALy6gwU7Yvni+mLQQFnh9KnVPzJ3PtUDvQKvebp9RZmcUI
maIcfYDuDukFnF2CBrf03eBwKiCfYqv3EYyZhhdcBGKFa4UdawFt96YNso2d
TX102P5O/J0ipcT4c2tRinDD4HyuehrKIh4q9+xV1q5y3c6NcPsCDszMsG4U
ELia5ToQ+PgFcNuhk7O2mhLfr9Eus8EKhdmCwUEUd7UA2R9dpxv8kt3ltVa4
98rubsJBJuIiWG/kkEyNTGP+dGh6jXlO7e51OWfgGpqbJfH+KiVvUNaN+tHA
3RCEwRRhxO+1VwDNoXaap9oeJcTlK20oQWQJoh2AFS7i2nV/ZuWkUWCmFFr7
53l/R/JsIgydcyfdd2xOvdMZ6VcmheI2doe4quQwxjOcb9F2azJg9WYahdJg
4+XMmBL6qLBt9UzK72KIBtM3XjvRx+nCE1+4wRGd2A1lpuvnYxcDtSJ0bvex
NyIAkt6ohBnVcqGb1WaK0MucblFQyiykWqMpG49g+h5aFC3TkK2qjA7T0vrP
H4LoBK5yAGvxHRcQpmCKo+ULbuDzgoH1MzBdxu1u8GkdYn7tym/J+INzdCTe
MVVvCWtp2SJR5kB5rtOahJR9bOsn81dCAYUD/plf0JADY3rSor7yYH/9/V4p
514exsI/qml9xjc6bNRJhNZ3wwjNK35P1ho6LSRhR/mAbnFL7geFq0D+4JN0
ztYvbUQT0E4kcZfyIBxugmjkJvCwcnM8peRKO2imIQiq8tYo/d8uPi2LdoVx
hwEKYkh9lypyopTb4l7gV9z18Yll2zvtbFgd7XtDmrFKYnlaKic3rmc30yVA
sNX0J2li/M87cjzMVTmpEuf1BL/bU9fCnGfBKQeCMFqjDUFjwuuxACAbX5pk
+SwI1GIbFXGiQZLzY78lLEp6GlxiIMYgwNOfrCkqkgl4v825Ogi4L96v3NrR
zr7SS6YLCUl0qEpbQ3iidJSFPkxwj9BFV0vgSLA6/tqA9QUrLuYd/3h8KKox
cBt9hX6BzbD2Gsn5gRX43nmnXf3mhIl4cj8qdCHknOVN802Bnayvul++zQ8C
7jc65iB61JaVZ1VOZ0ame5zyztJADWlHVJgewrghXTH1b8rN9WsGiy2N49eX
oAOaSA3EWA40gPHu1rjBG55EQzWb0fEd5367//3ufvhor6CsqEf+jVNCs/b4
ElJN+8sPcNB+H7fseDdhHMaoYzntOlXNxgoA045AiIGgpcxwCn+2F784bfVL
SoMGXsDiHizEuTp87LAnvCfpzIqsLcA9kPKvfeTM/PfYt71Djxu5jAizZ39+
pGa/DTShET1AigjyWz5Hk/hsMjlQe7XjSd4b9a40fYKVhWxR9RKobCkiFo8u
xvVH7TxM0l/agHTI6evcHMBRmntJxrhrVNU+6q54qciKyWkOmIKyHIwuWCYi
Xtg89rWKDO1jALIzFnpIcBhiNEv0NFQfTGQCppzqAMBUUwb0zUqG7sB4YEgh
baejTjdOeGQl2wmJoi+X1/d20J036fIwxsLhqIxiaqxrz1u88LxSN4McamSC
tO/7KTtGppygYMTwqakIPj70xx3epoVpfJZMi4FD6gBYXLSfDu+pTJNEmMoc
r1lUKRE8/rnMEGly5bPOGFjYSHsM5pSjduBve4KvpKe8CCZRTGbuICfKItyR
F9qGmEPBt2E8t+IYBaqpELRsM1xlIaKdAgPJ79nrWy1zds8BcZcPd6oHs+ww
ooZeDEwQij0wixs2wSB4CiirI0dSO7XpaUIXVaj+her85GPzems1pkInG7gv
fn7iABfYzv64F3MY5QP48uW/HLzKcGYnV2yGUFlQ4yNWt2wj5bdg9eG3dPBn
i3mlV6B5hHJMqQp2dkhVlasDrlFZTps5VERPKQ8uk2WICaRmtIFIyx0aFI7r
e79WkCum+oT5jrS2dQ/Phb6BXWRe3NmwM1tuqSV6qZq7EQdiXFfH7DKes9FT
YuMpwifWKFhIogOa1RkBAI3T19E5EQzsGDA1mGwSrXJgv3a44rWOoaFJ6BjL
Vpy+yOxDG0TY1hzn6y/mOdxpBQnJDETJG/mXjAERznwKnm60lDebPa3EI2A2
8/F3Mc5QT4GoODzVCxOrEge8wM321UBVKoD/SKkjYM8/okvxs5d+Qr1322Iz
ezacADCL+riR4/XyImrm7jDbGqJ+t6Ts0nWm21EC/KOUjlSmjxtls/RgSQne
AZXEN8mOU+jRmlZkq820QR0De/E9WoDr02D7uI8GRsvr6QpfiKFd1t66jzmb
RhiA9xkZILL/Qp77CKTW5Q3aR8AtfGWEkpjrLFiM8kBbrIHtD/nk/BV9zfD4
u3Dfiq8IBEH/ksmkbQVNPD87ZujD38Z8PB7on8Ptp/+oOoX8jIsa1yLVm7o1
J74YNGuj6O1IamTlIRqxF56+3m/kzEiSCojPmaZWzHdtvqUsY6moHzkdlXCG
k7NURd836Un+zFSEugPz1zSitOqlOnsAgEed4AvUxkMnG3YzlJMgDFSKu7eM
93S6Yk5Nfd/Gk5VEMQdvMVzLTB6NsFe7ArObHOFAdVzQQRDHClHc4nqilE3P
2xypggSzTRiTicf7n/fl+Yk0MmLyijTiqImElXYIEDOLOiIpQAZJjiBx/Atr
0M4+Tp8sn7ez+Gk7gXf+i7zuYU9Omv342LQMh6YjvRlv1e6gXD+P3a4R1Js5
VYMRb3Kh5Dxg7bovNngu9jNb1JR2CXQCaeID3W7XIsgIFTd55FEM4AqZLU/9
Ta7bzGbt+7GqrNLCqrLDwgHO7DDHSyx1htNmXeUlq5VMxPY/pgP2gsusFAwQ
RyFPgQpFtkLlCanggFiPTU9mE0sIOjK4y8LqNTtDH4mDQwnDXhrfJekB31Jw
PSjeXptlKhtLUxlFf9kZDJAOcKFoLEAhS6ekyt25ZMGJFHkoWi0zhC6g3McG
Cw5Noy9TprJBNb5W2qG6xFCrHdO7vRt3PEwF7fipJN7j4JZVUYjHBIn2W8O2
oSKcuS0tC4DMWdTDnOgSlViDPGfC/SBHbHG5Hnv5nFHd3iAjYXC3TwdrRD4T
yuJ2xvO3b180Vilf0wEiR4EO2DkKiCwnzSb74FwlcFIuBTf3kqb5O396UaeM
zezC3522Pn6bDrFPAf2+zcHpzgiN4RJPzRwJYGKuXMtpywiCW6PjaUtyaETf
O0hC2epXOyUH/dNUwixhJxS02V++YoserTvQqGU+DIyBOFbux7UWYcBqSYhX
Tg7tVY7bLuo+qvwB1Novx3Nexla5BctkxECb5ecbnL6iuZcc98ZcTScCBLdC
NtDDzm256lLSpZdKSmlVmg6RrfglnaCPF6uIiIBfvRQPlklL/CzVQubONkXa
tCESWjSwKIOVgPOXHu7GgtKU/6/Z2byWX7eS3/iVQm6t6xlk0ORyqNYzMAMU
hloIG0RSzswTl3B0hva1PdvHjDQRn9SwLqPSeKM973Hwo59uuaHPb7gogxJ1
6xOzgqOJZIQ+YQakdXN2kYp2ww0+mFy6shZ8gWPYbMcDMO8r3h9gm7mlX0S1
4r/gY5dgVY++C4Lwa1gjvijSHfV5pdBlt69RDLIByPw78TM9mtQJzwyXSt2k
xRX7XGsZGmbZq++o7uPxkHclLlj7eFnC9Pdoi3KcCUKhWA8iucnRTELojj0s
qU9QJVYlVTw8o/je0KEo7WapkRzdnLRUrinIKzQwZxHWxGPMUtLpnYOfgmZu
vbX13vRbQv/0kIiOG8rndjgs76uCM8uJv/HBBtpVdlxcMoc/2INvfbUTqduG
KQOFFnTf5FO3YQ9xjTMZyyJJGEEF4rJrKNTnfv3Djl3cjVzPYdYUSBbTG7xe
5fD9rlKhQ9/a2NhM6QWJRQenlibjUb54N/MhgD+CttRZiu9LPlIrnNGwf9bD
NTa2QSkLJj9ituhykGCJuVT32kE4se54oyE/FYHgb90/O/fTkrpmr6DYlQFZ
MMtkYoGZ4njSTd0vpvB7aB8f/up3KDjQYmRiJBJzR64Uqp9Dk55K7u4rHVNG
mo4/bfzH/3KbqPjNUigwlqUCfNWLhIMN4PoCd1T96EwRp79uAuV07kub/GD9
zaLvMd7ESN8XWEzjQzM0Lin76AXXBFJXw1f0pVwgngbimTL+ONch+O+tfrSy
tPQOFUsLfCjst8FMc8pxT4RBTp9jF48I1TnV0SuVhsO4TNpI1seCTXlekoSa
6Zw/ZZowwjR3b97Qf3gVSAKl8Y84xii4lOpNTPrZYaNx8KVhK308P6UbQnRj
GjWmKQb+1Mue1p8U/49v/GZfzhuOo3DV1cIF2emzPG9gEMQ1v8RZeuOVhUtL
vqQ2uFJ4Nc/CFVBeeZ8H8CNgsroHwPNR3gerqyqCc6W9DIlWUcrNaYI01f3M
IuIDrlS3cs2WHWy9J0wE0wD5EsB0NS4W7rwK1Rp8Ta06Lem2VraphXhZjgd2
x79CWJF2BW/72TUN0Jw7HxyXjfSx1wdYK8yKBhQYKORUNZPDARLIWA27RfMt
tnR03KPRP//7dSax+pO2FL1vTZIBsponCwFfEvNyABQtmMXcu3xtjSmKK5Fi
75YLACM9SMvBu8gMlFcOR8FZCFoHrMHtBmvHzsRD8cbVXB+GzZVXNvNT/DLl
8BOKp1Q4MyGnZPi9ACGoP4RJV112bTsnj/4Om+Xi3jHN5zHrKUJKVXMJ/sO+
cuSR6WWg2jBxl2l7eOJOa7Qq2qYtQGqYWxH8wJTByAHsEDSOFDZ8F6miKHBV
FkLvQHM9vYel4L0JI1IvM+bTHI+CN7Vw3+sRfAsrT+vTtLlefp8O/IgLuQvT
boMDLqj3sSwk5ScnuaB0iejbFO1jBEW3I9sRdX5uWCF2fxWgGW6J99ZLvcYP
PzNKwwzseAufVzsfmEBryynAttX4wnt5gey+k+MjOFvGdbKFCIuIx4BHhBxx
CX2pMPtsCewlmpGLS38gAxraHVSkmWzv4UdzChrY7x4NqjKjOxvjekHEQuKZ
6fk6l8dzOiMBYShfVPFPooFVY6KVnBcYPFRR0WiSjWA5wwXyGvG152fkeQRt
sa6UXmztpfxP/MIerq196S/NrxzaBvMQyLW7Nl1fViVYxkA4s66avE1NB2kH
phaEiRaYDgtLdEn2LEqFrrYLAa3CdpJYYrSmluYZygdmhQxY01a6RJZC2DaW
J/loheky17KB66ofF4YPrcBYJhqaJ7/lEGU2yy/T/4wa+QAMMkPvRCXJzNCG
q9Epp4MSJd/MDJo+SHb08711wVB0n64yMVZinNqccywd18V3KW5JVstfcyNu
SfiROx6TQU74Fu5lfeb96qOOwzjRQdT8o2tdnm0wmWFJ84n6hKCtECheTIoQ
HYUQ0Lv1QN12NM1MT/ZzHa8CvrumjIoNYmCa6u5omsDNuudKtoxJxxaqYmte
emZjmmzKhuI24v9b7bAPuovKYYpUBNJE4xSYzxkqW0OO4ZYEIMOnvMr1seyh
4Bx2V5cJZJjnDfuavKHugh2V5YNGfPqtKuNJzTVXWHLo2A2n7ig/OW1B2ZaZ
mgOtv8xiGBros9zllsUnP+21vnvhRGmHvYjLJzTVmi6KmMioVs8fdr4kTqIS
DIwQoFRni4P8Jh09cbXmH19UAC56h2SOufyxegZOJjpnM/RkSLTku4I3Hdy9
qltTAx2pz7ALEnld6UmlYL1HHrVSHrvUo0SZs3mwvPryoWx5xPqWhLWmz/So
MKQ2eqgvhy/ytBjhlh4vEJ7fDmIkxS/Dp3VVf37DV1L6FOMQczJsVEx5d2Ox
qlyWRVE7cE+RqrlmM7NBdnyYG8I2Fe787aRiprYEvaaFUwysB6p/Q0noU7Yc
kzeQ+8zVG4TSV7CIhLXDWw88kOyZMI097oCcU5C94sJH6fI5GxKx/sVT2D7Z
XnO42zfAXRM2DzCMTjqhm/LXyVqGf6V0ZXWIOMbsRuUM98ZiASUNWlKLnRP/
mh4qmc4adcmJg8/qHXabmMJA+xuMcURgTG+SkjozgKiJA7BUMgRgcqLzY2kH
WbGzTIS8+gACYqiyDQlwKaVMkB7A7VPe2jQXy5w8jDVee66e059sUsIlq4h+
hs8jgNyTWLDB9aWxRWf8vBESvJZz/MaP2BA/eQiQeApwUjG9MbK3pIpvISqe
4dINLUlCK7xs1DDGbKdPdCrYiA/hjNLl8sYidjwT06e40v4TyUxsu9M/LplM
G7Cl4wZp99jgHMiMjwQP6NLL61re0rlcgJCnCh9T+LdnALjm61PGsujFBhKx
vIepQQK3E5dMxK5S65/pzoKIGuBmv4w/8G3c/IM9SeqkdeniwPPuk+1/KouA
JUdHDVm16q+M/JFsBx5qKrYQPEFnkeVDFTS2WiX6apBjElAaY7wogOkLzOUa
5AFr4Q4MJtRg/8Hmd656dy1KqIEJgwhs6bGxHNpHmVhaYGc9v2cLQSZJC7L6
PXHOx/tq+wPsmmqcskNkXOVPQeC91YEu77e1jklY5HZIqSUkCwMsDxwnmePe
RMechVVbyqvOiJHPZlCPz8Z4B4Ehqfrbp28fNAz7OP/hvrwsQo7MDEBmWFWH
AULZlXUkKNGco4Ir5qhNMZ+UhKFmN9VVg1fSh0Qylaq9aApU+nPhQbUh5GwL
BuSvpWDx63Ks83uWhxc7oGycGhKlG9AQX/Nruo4GGR/6G8R+c0Rq/hiIL85q
tIfG2ALhbhxXhRtQ+dQNQV2wrCrtWIuDymkQDqc4oQOR4CwPf3OQb0QKAZOC
DYeWAq70vDtCne0992T1oASwngqRgSSDQVt1UZf5PSNiPA+JLhhxMdUWk5y2
J31lca69TkeIqG1VEcVmFTHbF8hOH6EuUkTr+GZALTmgclz48PgHiIDDD6kN
lko44cnfQVyBAQeCOEMyCMrQV0p1Dy48KEhe22QXf9qh10ZrVxcJ1c1PeaUJ
5QglDDL9DOiy+F1FUVnXRFg3Nfnx7+1Nk8a7ibOW5nQL2oQTaJqhOcgjoFDn
0TVKMswhFACT0nb8HdaS8QAJeJT5wCwbFXwFFGFrnfaEqF1EHOHKV6EhMw0E
taJaJjMk1Z+iFNUBPQoTGBrlPa0CFM/tmDpRwoUMYlhAxYhghnPQD+pmaGi0
V7Jws8/fMv7tX42DUDMx5tRwC8CUyq+KRLscSxgu4CueArZeHU0eYrxiGZib
bcKzjovPxr4zJPTM8T0tDlEKfzhjyiLzvANQx40YL8CnZxvqQsSp0e2fEzHw
jiO3zPahUu66Jg1snKUQYGpSazveqsZLzHpYYj/filZnVvwb6s4qkxqa1Bps
S8MLif9OTFh5G6kV/PAHetNM+zQAdQpY6lLyNuQ5vyRxdakxNFZD4q4FOl3b
NBeGN+As5S2ch3M7X1V5omqQDI9Zcnh2jLUviLu4crRRC6A6HvebHA0rV3/3
Cwsutbw7VsVTxbgn/64YmmDmthqDaFxxoWruZXRwso/MVE2U0ew2/mh+j+Ht
mPl2Tdwkjc4zqT/044wBMLu3QX/+p9s0+W+qMlHJuImgANt0JR1JB6UCMAZ8
3aJlZN9BhPSdfxHazA28N7VZh4o80bc/mij/menaLAJJKhvZMa/U1bZTeWLb
ssb8UoomHBRJItwhnWD2OUKaslJ0ZqsLFhzq4BHwv1ikxOKiacAYUaWd7Ki0
3qCcwgT+o527BBsLaNznnaoz9tgSsPVGSeGpe217ncDEl+9ZwnYK/2eWd3aU
N5B4SziifGg7H+FTCnutyuPIOcDbpucGoUdYJeOktebvwU7Q5Ob5kpnKKEFy
7ObRhwDOl8jHngoDFO2ksJM8k3EbZvZiSJCXlkg6m5dyQw3QGyNyNiBJW4UC
bxOd8SlxfOJFvMgImLJ1dva6LGyK3+onPkVKm75ES1bfF8ipThK7UYlUEKOv
DdyJmhaoJmNOxBZbF2cEKlgnk6ZOpvrFB8gAIXU8SZ2teyZkR7TuHdKTdzs3
O9X5hc0k34o7kxMyUW6z9p/h6nvXnc3P7sSEqaQSfTfDzKFxe9MmjbYOybYF
BxmaLHTMwB038YRIkafWrdWwNiY5flxIzprg4OE5DSLNrG4LR5vlgx+OkBrU
EBSiYfH/JHEpixVHURXBj1I771J791XFzV5o/pZDrjvkGI7CEGOoS0oNCMTa
4nocUZA5yA2A67AKgsu848FZ5IvlpHwUBOXn44dzpJzrEkw/HuSLbbyiqN8M
X9xe6RCOMp6w200Gaw2grsneAtQhe68sE/JL2JkbpnAXK1cFWFa4boa/oVdY
ek6AFa9mk2vZl8IRFvxe+KQjEDBp3bT1O8GkC0jBSCdEktQJiARyM+7VPfUC
tH/oPqUy3j4ZCb4LFurLY8NWw6VP56K/mEK1DcRo4nFHt7eAyr87GZJnoHkC
4HlgKFoWPIgmFPivpyZ+I2xrOhj6WN+MR6rnvzdpNty/34CiI7PsfCf+kVWJ
o0dHXffhHTVUtBaRfc+3rMMtmk8+xmElU2XfQa2REQtVhiB41OnRJ2bpMBxL
MlG7i/0TUA8gdkpyTd8TKXwP6SNfa6zxKKf/dOIZPtRGxmo/Alg0H3LUaBA7
RZHdQH9p4m7803ygzxiF8AcdNaUqv9cZ6wU3JKqo8Xa+GyvgWJtW4vV6RKdg
/dOkjKiB98IZEyISCG6yuKva6oPaZhwcMJHU2t29kN967gv0K1tY/hnE2BAe
/H9dImP3w9ebtqWROJZg9u/2y5vTfemJmGYY7qHsVV77WDZSZvdMr5i1zX8a
CFAuhrVztvKbwhRKJq1QQkpSlbTAjF49vx5N+GmNPpSbRhP4vJD5TMM3QeDX
pu3x0H85Rd4RAIRQfILN1anY7/CGLeoJcIvaQe/0siES59vpIPP8Le9pXuFk
dRV6TTTJrPvubo6RVciHp92RJhsomJFiezCqwS77hFdxNJkIF79y/JPc4jGv
nPFs63qt/gqUhBLKWAZqcx9p9O2SPKyt4cV45+tPsEiKuefcV5B3iLRdlqiO
q0e2p87d9AV+sEIvVvctdgnqs9NRFK4WlDqWPOgZg7Es0ORFX8/PwZSnFZQ8
RL85FBcpLnomYHrNLxuDU8ESetivryepiM+54Oy0WDLAH01B0eHuBaPi9LVr
2HVce8KVkO2HEESfNHRQQEwlcVZSAz1Y7c81Qw49cqlVZSEEuclitwFzTl43
ZmvzYmZOTX8QNGg/sPM7jtDBaIVKzeuNMBt0/GItPpA2//wGff7OE8314m+v
6rBw0PlWSWbsMApNqEwwDx7SK9mgtjrB7qrIIVQMWkyTXEjvVOmiAfVAQ2je
E3n0SjPXEEWEAK0+10WsthypZPSUmAj6HlN6mVuj4j5dBLhPJ/L4qDeKOPhm
ePBrB9ma6M8YhJVe20NWmp7J4eACYl4b4GUsxJwjp+liFhNM0pVZ6gXs/a+A
VeOurRWs804cZfQT9G/r9ElKoizjyHKXYej3S+1r1mjZvwbfcNc7/EdQ7T1F
du+Pg85XUHqVyU5kI8U6DoDWCm8Tf6W1ltb1UcMhPBOKPXHHlVMJxM3iBI/l
cZl9cW5kt8250peWjfTujDw96UOmOcoA9SuwfBiD9MQzw8X8R8mwla5y6f3j
SwUcWbSNEX5DYWo8ACDaLxyRoMVPbd7wwUR7VQzVe8kgxINII/2ssDY7ju5k
KScetAHOM3DzvXW3PdNnMMFiauIylDzFNylZH/K684pBjRkXPnRvTXAxu153
XtYY6F8xuYQpz6Szw9eKgSbcTpAYK0mnJ6ZJgHBK5zbTgK7i3RLdF7kmfD2N
Qyk4f6MjolHS/Pg4lULnR72aM3/4UbD0/Z74Mc9z1uZ/NzOvhBhMvDibRz9X
UzeoUytdY9EHGDAomzoptXTEhjS1k5GxQffkToHXTdlS1OPThYKAomiHLgsU
+JJSFpsaJizH4UxjXWEWcZyk0vyLx9v275JZ+tIe5obqnFYlu+cAc2mJp91A
NgEnbf1NARoiKQ6pPrucC8aJJXiHcPr8wl/YChZqfjloEIsVj+/A1gEXKlmL
oTj5KewftWCV3R4FAjtoz8UQgTHH/4NAbX2i3+qWzf+yPNrY86DSwJqTg/gb
zNuiNjcCb0dS/AqPKazFWrKdfi8ZeU0djBtltGLjqjExlFMvc5/ytZtuetRf
pr0hsfI5R1dld5lGGQPBuimYBrMUBlvgKStoscTgI2DtE/gUj6YSIazCMNE3
ZEFvF12HQzwlF7K9KiVNhfr1ciVT/Nkyf6EUAPxbAwkZvVpfk5RygiZyjQ3v
41KgYsy9FkaZozZyi/h85I/JxlptaBMR6Su0srcOTu8d+83rlMtqqsN9xxSt
4bkF6LhFOor52Vz8G5A1FDgBeeF4M5i69gqvenxcrVsnwTf1r6HeoP2LqjSt
sACahT9wUk9nOkWQ4h4asr5udGoyCLJtF4R9BRXnmrcnFpyCGYaRL5nPwuEs
y2BTaJdpS7pcKRNnYLXV/wG/WuMEKZxF0SYTSZNorl90VXBVKOoRX+d0JfdQ
c6BZ6bg1Tbu7zrNI0uz7A4TSpdzoBy4NMVSSAAB6U2t+YF+gbDKyrJm2+q9g
n1OGZtWi3Z006rnFNnupfZIuu+KLF8Jd85AHdfLT+VCTwF76CtOrDwRCv4kf
E4sITqerOivlm6yBz01AVDIDdqgtVFTB3Mw9clRK1fyx3eH0NpjVykNGx2tj
nmkXaZR/G16hKl4849YwG47YxusG2ScI7zuSad6Z4mvQZAbjC2sb/HYKCX6U
HPYkC6rRnCasVsPBxgnTkaSwXZjeI2yocg21gJqmS+HasVsyDnoJyPh3f1Tu
knbDw6cWpp/MqhxdT1mMjBb37zSsYJ+/b6lPXB50L9WAm1ob3q6Pu/2a0Fku
y/oppymg3aQr5QOy5zcy/Ocn9v5KmaV3pwyDmftCv/9m5+CxMahgEwWV0nJ9
wt5BaU9UKCtbESQPSM+fcVBFUuzY3Hwswy2sxcy2pzaCgzXT0+RVjSqC0F7k
jt5wDuTb31D/MxObkRUd4yMTW2hr9ejMIpMQSYoOWtK+0md9euwd66VdOevu
5xkmtlE3U/UH0XZhIiMud9TEIU46NVJYivHLBM1Nvks+IfToJ/iVSWI62iX4
5v3dto8B1PW+FIP35WnxuVtPUgpJFrcXh5esuMco57tqcgK2JtMWK8FvmY9n
jVTdQJEdKPS/YfiJUpWGG9rbU81PdcwBmLmy7MM6hM7Gw47UQ9r1vb1Iseh5
zltcPYD6k0qQ+DdD+kq9H+GoMdvmW5vPFYATxqPMZpT26zD5BZM50oO5UVQb
0CTYvdlXSkCJbPZ+NJZ5vP9oO02kO4gQIJ++saxk+zOFL4HzjzEWu8JOn/tb
Ft+5BoEYjNRbD8ATtC3rCGsn5zMYK2835xwuyDaOpzMH3tZLHWa/ln3L7HXP
KErbtA7kmP6Xl2DN4ZYrCT16xCy7k/TNfR+rvd8PWgSdyqKKH+T1jpqj/PYB
W0vGrUU8otvmw9TMlBx6v5ppipzuU55pwssMkB8Dm9xurV+SHgCWJ0BzNLOj
C/2VWkhCWy9SE6f9XoJEw/E745ywWqo4ANl6SGhdYgNo4QN8SZq16LWMCWHE
WrJ3fHSoLS3Dq1GhtdTok5gq2EXPHnSeUEvP9g7HdIGoLqDlZAIngEApbfQI
Waq1CgFo/XIHgVrQqCrteMv1R3li7jAUjEWyiKqCnXlj/k4L3o5w46PrU2WN
nEpOG+1a1JV/up6yCqXjBGldB8apvbd/QZ5wwbrKoc9e27RQ8iGykyDuZojv
9jrdRTNx3XkQGLKUrVqj97DeFM+7sP0338Nypy8g388F3LlZhXbgoHiQtNXP
PB+qQLJRjNqH9TNYyMPHNX8eZJe/jEcfi9nEI6qX4D3THwh/qSG1Q71mzUFg
IVvNJkATKxakV2xP6V0Y1OMc43PQZTRfrN1IG277bm9+loZnDkRIGbh4qz23
TO6fck8LkH+L2zRjqeejad4lSoTMFglcVlGe85rIRnIwpdHNRB5YzcMpMi+0
wEuzHqdBWmwJ/4SAl/q+qIF/5p+9WoXDwNIQG2Q/00KAT/OQHkYGrWRM0vD6
9vpP7zoiWMN+Q45BqHzZZex7PdIFieGv1ZP01A9zbF1ZVWyuE4YHmHTZRkK+
414T1ZIDU3letlj4Rq76cCBu9JJLdJx7V3CbLkYWT+weMuomSm1/wZYIYA+I
LJS227uYvlW1TWxalTBvaKyTcyVZqP/xHFB501UR0jkNEQLadTO7DG90zdMc
sqKGV95cle5AoWHcsq0jANfRKSkEzLGGhc3dbN5SvtFNzlYNIRzgeIBekKK9
8qJ/MCDmayyXrpJUgjz0cikBBK4lMlj0osyq9H9vjUt6gJ60e08FfSM62dyp
sp/3lMZhaZDz29UTC8sHSUamdNrnFLFwbCATlqU1X3cbS/1FGmkdTTh3reE7
dZmcob4/J0fF9d0/jGrsbcnIvIwlwiTRpOvRl/pN33+7ZftatC2LXQjBbtCg
WMuzac6JyM0TU0u0GmPtsVTXMEwIntPIjOzWRcjzAZyMNM432ZihoTT7bHwY
6fKuczLTPSLTq1o+6FzjmbyMmTyLrt7Iro6UuDW9JQrrO70NuVbmyeyo/L8T
BXRJHy5G7B3VfewNRKygOo2t6X0Ta/N78V4jI7pb13jrLbgn/GO8kjH6oU7e
mgLkj5dSlRWBdhfgWPNXBRi8ibeb7j3DLrorefqmJR28GnwLex0S7A2Llk7t
XxEvVuvoXDXf7fw9l0fw8KJT5L6uqyG5amIl8gH8YFrX8JVpkO0L5EsWT6oS
KAUAeitP91pgQyRvldW4AN0b4sRy6BKy1FuFBX9j3+T3rjgXjN7q50nagfSZ
gvQBvf6T+KUay05o/fAy4T4vsJNzeKlZHnbt8PjQl1x1v+mVi2QMZ3I1Achn
RhUkHTpNeCrPM7X7vtSpAqTg6GwQr7f32qY7axaVosli7jqrR6f4OaP8MU8V
/ywPVqUgyO6+BfWbrDlvzdCIq+e9cVcB/Y+wagNqL4Irg/jCMtDEMoiiBHAL
qRKvkWusj097UmfNgDHIvBg1bHwN6Ri0JrcoOXA+XanhEkQd8W69FdvF+g7F
MbSzRPTwDMd/5D3RMLgB705kWWWzyZXGHRkfquer0UzqKvhe7/PRXJ7ILd4K
2dO0QQFiUiCa/bZPQ6BRZKzd9wfdQKqC3uxbZQcqwA88PJMZc0LAbjC4ire0
XOW8IFJ/OP3aNe4fbdCTduIPdzEVGuBn7P5LOe8WcsPstP0uCJ/d+RMXWBbd
J0dIhDauQkSebUVtMzMP612Lur29W2QWlC5EY6EMlr6R9zlGtjeZ0LuLnz0T
6GAEzzyN2ziSSFDjMvtto/XU028PBk6PHOmtjBGbG+lZrazWWVVjkZ4l2+el
uySbK/DUuiufrgL7UBSeS5gumYdcKmRIbhBuTCz9F/uLl6gyfz/AQa+mZY1P
jYGP2w1mkNqG3t1gTsj2zt4of4rgTnGzFuKM5yRBBCNLLBMB4wW/FOy++lYr
qYJ5PvdswAG5jA6ROvMpjzNbyqLm9BdV6Ah9k3MFnOLePa7Pc20ziGmWA3d6
JYiVTK9AiSl0P6zQC/6xInTHTyrfFFeV2Rb8Dbf867H8E+gLJQQI9cjRcpQh
n65UMLbBzcepe6vAHRXD9zmUuNO5s7VOwvb+x5YrhljZf9RlwF3Ynixpdo42
ciZHH9FjKF6b9aAXDZGhcoggr6KISm1+pavz+aZK9KnWLjwLEydMDrFJfqkV
yTFgIrcMqiv3VSowgbJ2SY5mEh8jFu+rW8POaLWG97s0uX14XiLfkTkrMsW4
PlYoiFLj0oh4RdEMmVBTqLociVSdGdFmuhERASbsfx9t2Xwkq0h8m0dZcuKS
h00hU9qjqBEVNHC8u6Z+2GNgca9KeM+QZzjKMaLWIw7k1Ag8XaIqn5Wmg5tu
ULpj2Tf54BWEfBhi6e23mRZG4VSa/pfXaXoBwu33eAeVhjUOcs7JGwypkxYo
DezNbN+YmpCCyl39GIaURdfxb0KYsO/OKKSh/6HItciIAHWlPixsUp080IiP
+0VxujXcvylJ1ka6XusOVB/md030JzmrYax2Cmu4brgZOqxXQI+Kx1we2lbf
9JOXBtwYpr7FaZjj/0jqJ82I4IYEjfCP0RzeWyaVS8Au2yjPUyUsGa90grm9
47RYuURv5ZbCFjlYp0CbZI/i3pWysvqfcli3hZReYnJO1cqwhuBPDYQkE42K
pXDcNOESTyQG2UyBjm3EwAfYx73D5YkHf6pWChz5Z0oDNpfSeNtaFnEBF7XJ
Igfl83pzTkBHlr0mqR/jZ6OjB/IKDQig9x5LzuUmVyXCIvq8GrwWw9WJL+Bj
mJcBe9Yn7dyxJBMcabTM12K/o/G3iNbIQbTeaJKcypATUpxb/eLLg/DydIRT
6wszdzUnsHg/vlEZW2dgL4DtwdyAn17lEXugTwOO1x7cVBGEC482s9fd8bEb
vP1yHm6fs201yXGSE3gQtsTCF/6ww1SwjMm4kTNQrcXI5jH0c6ORqs0RkdwH
HeCy+ysU8M7P/34AYK3ktITLaEzKoHMHSZhWBli0orCB39UY++K4UzDCMGZZ
HGDGBAUkohXEgDycXM8pgQEQkP+goFzXHQahVGb4E8syALRG+KqbHaBhdyUw
vqEkDgMVjuwRx6k9W36GB5476qhWob8a1dbrcVjv3ER7juS0k+ZF8CtrEPIG
SK/Mnrj/Tsxmh3EnGSdKpEfvk7xBPr/pXbfiir67UZ6On0wadsRu383m/Igi
Vzlo9QEcgr0EEQYTa5pWOhHVsia74IVRt5kOB6seNeMUKb5VbZVhDjDrltND
D19evDNGqNvj46Nfjn8XK5GL2TRIYxy1YdcOawrUKMz2Up0j/vzqbiJ3foxI
kJZBF4EpFn2f7/Z2UN5re966be3RyltWm13vRLavwTAqL8TCW4DdahEGVDOx
aZzwz0mJZQokxGwHSccTV8h85sn16J9S1QkVeNHiZ0uxGknj0KgGd3f2vEO6
fick9RqkHCfvGmKbbDzEhEimr1vJkIScPVQw8ldTQY3YAnwNMzcBGYw/ueiM
bHkE7nXaJYuxPwfXaEmGQa0bS7iJZxvxIiexGvGv8BZZArEJI2z0uWBUsPYp
Ub1jV2oKZjhebvKuKn3Ywkbcs6HB2WJxbuubuOo7bF9D8IieOkYn5CE2wJU/
VyRsKEmmLfxR3JQcQQa5anl0hZVc7DOUY2jIG0P/ZcOyy1Zq1lBtw2ZW/T0C
S/DRvL7mPQPjnUtOcbTQlYjsLeI3yO5qqMHZN6HieXD1/MUxsHpxc/KAnWJK
b4shSHhO96bjM0M/SLjPbd/KveImMQE8henT4LCtBD47d9ea2i889gxBXzmJ
jqFDqymNxDhkIdeDX7huX+QbIlXTGSxztij+c5Un+MHVMyv5xipyFU146wnd
Vc989EIpF0eb+w2bStz8X4ZrugOwk75/Tk/IY+EsrPW6B0F1R82A1Pnd8t8m
hRYeu+yliSsT1dIjWUxxLGs/VrhA0aJACAxcIWNHi2t81s+JtGkG/zG1j5lQ
utb8ehmXb9rU2Ir6hlfW7B+XGelwD20RxF7bUgx6NRkZ0UXDj9Xh5qhw9lJ5
zgmNre9nuHz2gETXILuHcaz+wONqX+6xaZe+8wQUB9b2GTue3sXgLjYPOzu1
3UYgy5QlvnjPXsYCrVb46Mz8SLJFSUpxQQp7vGlYsrbXBhwkc9Mvp+DkSusp
67SN6E9BtJ5FVKNjOEO/rRQaqNUIDPeU76eIIkxA6w0PIWlRLKNd4N/jycOW
meHq6eLlmSBYvmD9HGx+3mamocRSmqIxMvaGJOmf0EsEvnNrzgdzNLNgEmMf
b4VO+3toC6puTvGxThEtspZIWDYuo3UnFqe359LfsZGVlEOA6cHne54xTylA
EXt5T/pib3MZU/VthIZp7oRc5pcL/xfJCBcZMPjUf3OVHyKk5/Kx3JJWHejf
PRHZKOxsLbE1vM2ytFJ90n/iriBKj0tsNisDDq3QY11TbUSvZfFjWt6NIjrC
kbIZm8t5VNfAKGSURy6HyWzAiUxy9EG9gsUDLsZ3QQ0Knj4C5nYOvjdS8G2f
VYoUU14JmG+tLzQcjQbYl1R35fdmKJ0mYz3mRN4QAbXrmp+mXS4goYpj/4IR
dQ5xcYRLKKXRNGGbxvA57UkTDw48l8NksIaHvEp1jcdnyorMmerEA3wHUoZD
X+U0Vvd9UbllF6GyRaau16Fp3gNdhXXbXzTVCm5Zk5dGXGX4woTJWTtlwOok
aIwUei+sxG8l1rGjNYhizsjWBfRIkk2KNJIuclxXVgyv+OAdLJmYI4+8py+Y
C0Sh0+v7QSePIQ1SnThh3s2QkoPYcbPRRnzaYftHy/MJnyWRFXYTNYsuWioV
PQzsqB9g0ehRH8rlfGbD5ouAwLgv80K6TL0gyS2VF5HEYnoNRn+WDkNHiWXP
5lLuGbqjNuZWNAiiqnLdWtDxVmbYWtuEcty41gbHVqyMS+5whye/5S1/119f
NnF+5ZPTgdF9cPEX2nkpHMbfjV5h2feJjKpIPEYusGPsxmIvEBqbvi5eJpM8
dwCzl75RP9Z11X9UMnwaJmC8Ys2JgibPEK59d7umtB3r/OrOck6Cd5G9kIUt
cUycaT8JCX7X1WiT/lBFiQB6yrtuTCsaHNBeP/bk570NMr9Vp6IwvTEyyqK/
+CfNH+5WKGd96eAuZ+sBgnBgOoGsWdSoAeCk/M7KlDzpJg1nyEJScg9wqWZr
Iglh1PXvNEO1BooB80+4pq0oTLM/iMp2pPlvakuIWk9XLDLy1bYdyky6bJnv
1Di9DU4ubI3RIrCkaduLDNyufL74a9dkeOSgilY2PU17M9Y63AmMRMfAYhfT
TJvoSWYrXvjzmVNNZuKENZdrzKXxEdIWm4vrj0wGhNBgasLEsTxYguB7SSov
LSsVx3qGsxf/fDp8Lqu614nTgYEBefVmPKWimzmHNEOhn4EB30bxZ5cjW88K
7RTCXEaY2IpJnuo5D0H5iJWs9gJezsmth/rlCpto0Lqv2g4HkVQBz/OhFZSq
bs6agHlwCzGt/ggYl+asAD3hRYv/20w1pN2cAX/+/lUnLB3K+A69ngYrgOq5
8OlWJM6BmnlVUW2y4HskWjf4+/vqubYRJAjedF7oKLhTUlQVocSpng2g6Klk
acUwUQ62eCpk2ngoc5bcEjpSkSYa5YBbwOwUtDSfRqY6LrkugC1J5mc3z4Rx
eXClt2pl2ne9ER6ImekpHCwDpMrbeMW2imMEHfmZw9y2ao9X4kntSt2JjTbV
Ve3Fbz7UVIXEYi7dtQlYmwWC8uaEusliLczEit+RNg9aOUK3myW8C0S1VlN9
NXR7rYCxINAePn+fLmqgrr7+oL/ZIWeey8jE9jClm4vtMM70h1O2SeNrUlfs
Xyva++Mw4ZA6yeFMxFgU5gYJsCl+tPvPJSFzUPIuDbgj6Xb7bqUZBME4d8n7
Hr0ym5tIw/GSU0ZEftj99SMnrICQfFsfkA8c5suiYmr+kPASs6VjX8RXIEzd
1zy3qflauX4z2uZTDcBePX6tViES4DDw3Hzj54zunZ3IUAQ37DXKtBpAMGKj
StlrgZdp/pmLqX/ttQiSLaPCEwsBtscO5qjJOPKeugCS5AD4o0mtuKErf5JS
Q978k59qNQ5Ib9gdpD9sNMd3YJwvnd9/miHjbS6LNMYOSNbVCun89oLEORc/
1zrJ+l4K72aCbP+vSzz5aoUy7Aoq4P+KGS3N+d3NTe1wrzapXIgUgXm2DQmp
bFpwfN0NWUu/5+dUayzWZISi5x0oqcFo65+OISdfq5Rm023NXhXG7E44Kk+f
iopzki0lLigk51EnqYvU/SC19qEzKCrRwqwl4lE028b/tCZhDiWQIndbH/1R
LyzUmESKdkYr4pW/L7LNsB3hhg67/LcInueYJCzKpreB/je47cbZ4C5A80wm
d/EpXe2UYxrSyoeZY3iWBI5SNYLQbKdcGfcRZO4llTEqV+BeNCl+28+3n6o6
FE1ocl6zKBhPgpXnSMDbrn3RAB28e0rpx6sePXBlJCreSuEeqgI8WvIcN5WP
7y2tFj7+zezRgxNyX9TexFmk/V/TXcfD9+Itxhq1YJiwZ0AQnA7GEG0nH0NK
4jlUPjzxNuDUQWS0QxOChM/4Wu9c2jzFB7NFzRI6i4EK3W5YyOauWpbhccie
WP4ZsrvFBJnz08Gm1Lrcym6OHVsGH51u8ySBcmJE2uCVVCZTXPjVlzB6r1pj
O6HR1n3d16fJJL4MDEjaPV45NUJQGam4t4mLlhfpTIKI1T9+6wUeA0XSMDA+
IDT2k35kIlA5GQcQGLxMzXLXBMcv01OutPZQ6l8BCkA6b1CbqGzyR11ZPs+E
7wYGAbpTkc3NFG9Sdq6gsjtsRvf6Ry045JuYMdi5ql5H0G6fJrcwX3vofT3J
YYAE6CPaLrGfLWN5mbno0lqxwIhMIj1arkggpvVGSIHqQUBIqNp6g6RLZgLQ
nzRx93POSPIgCCY1wgy+Q0qtIFc+PJR18a1SuCwC02gfCktGVCDWdI727g17
Fx9IZMaECfy+NXV5z7CaX0V0q5Q+mIKgzx8+vmgrQ0Tvv/gG34vKGFgfVmLT
DBU2/TX+LUHN7tORId/7I5OaK8i6YsxUccnF9ujKpwJyRIMUxOXfTCuGUtNg
1I/xhzU4kNIUseJoKNB4x5d6djcHRvBUnJFiPddpr0eQgYkCbgkejCM1mW66
/dpuu9l77lFzHGoyyjRRcx5YPkcfXqMOvjYiwCYhwZmCGCvD9nUEe61VyQ/Z
PabBRyMNt4v/0j+1w6Oo1JuwpQMVNgfAF++woNQOR/+RXinMEHTSyKMV3qL1
UkoCglKf7amdjB1F6+AyOFsFoRAsn4As0bvPCDzADkplMiZUgV8zsYLQoRNc
/BNVP6mpz42AsEnvokT7XmajGwIBJRgZHI3zx6VFbqzKXdbMusBP9qUWB+q4
ca2St9eu4mRC3ZZPwUjcY207Ly0mE1AMdsrY+IxHJvCptDxLFHOCyiqNCfmd
kAGh/gdFq11vvLLlaHdtpOjZUULcdAE2NM5oNQGuYHg4t/MEKGwbKKARzSRp
Ldv0U8Q4p/14gGcAYmx1UNn/b27PSfHr4tMIc544nEqaoxy4fLLZXRtZPt8S
PhBe1vUEGbb2N/8RBSnVblSUAlW4hIwaf5e39YK2zhNxxnStG4QiaJebkSfG
a2/CbJ/lQ8BxqxUwgizfiivel7MkLxvp+r+sG8JbK9CpbFl5oKmjwGA4GzV9
b/XkG2R3n0P5ggwnTyicGBZ+2+tn3o3IMeCFRl7N8Z0DBUrd17MsQBdG8K3j
1rgZ+hON13jXdf7xo42Ee/ZUH3cUjRB4FtHI0IndUJV8wthoDWMhbJAfI9Lc
lbjZ2NT+D0Do6gZoRo03yuG0idwIVmDwQgfinMpYdGyuKPUuwmJSObph1q4B
ZJTGkhKWU6gWls3rXANEOKwDivPKkx+dqzCos6ndnKcFvOaXGAJ5d8r1rYXK
2FaEWFCYGgqS3Xrwo02Q02q1XbfWZvTKilMu/7Byqm13qHdPo5WGaQKiFoTg
rH5De8u98Ddd/BS+EUTyOqw1dQSQKK0yi7u/axG1WeW6URXVmSs3e/uE6PUx
r12bg26rG6v1J/kHDYxcvFeK+cJSOgUrNgLAUrM5OzGJKByJL8HwIbHffcEV
7hSrBUaLllHsQk4+RL1xxqIg6lW/YZNj51lV1jmstB4bDxzacE+BMli1QOn9
IidxklEEfm1LXhJ1KLEUMMaCAMs/vHiIs8iqEcQ9B4zZR+wljs8QpJvBHoXr
EixrpGXv5qyB127PkNa0fHTsmsAOD1nL/3ev3+zspx8ieXNzOJ9x+n1vR2ma
5lb53dPuN/JXqBXcA2XMFc1WWRriRQVPEfG7WewAVqlusWvOSuegTXJFe8+5
uil3wGiqXb4FlE3XkTPWclh1kvGZ1T6ij4MBAdVLaQEYljSoGyzYAN/sK+Al
JTitQ4RW/xzHsYOJ2SWLalslMJwaqq1LQd9ohS06eu18l4I6j8J6R/u+1ANn
djnPpQ7omYXs+sCSa6npOpwdSHPKLvM4yGqQILie0eyQNJvshfJeH7ctnRuP
pHCE8cDx7FYKE3ZEtSIOj3aesk2HIiFegP73wmdBdQD5eiSri9OY5v1JPdjS
06XAs2w/g0R484uVwM41ZkKhJErx1BbHu921f5yZie/PckDC9+hXRHh9HFTR
a7SNZNlM0QrnWnzBD04mF1II0byrpC5ZsEcLHXM+D4tr5+jNQ4S70TQml+NN
ngxCTSYJxCeiYCgy6l1aA3xwb/jaO0NhXprAwTVcJ7a+uUh6difWN0LFdvQv
b++IVtx6dfO4kXemWXn1pzhCSNUWUpXkCWTLvz7SeZcdMKOkpan9IwVqbVKi
jTBYYS4DOAtJxp+Xg9RR2zu9de97IHTlBnmBydZXbcl0Kh5jr48qET/YnsC1
N0Om02/zMtJIRPH2gu06eEoV0/ez+JPeguYcEsdGNeSnCoPfn8cdWzOJXPoV
vhLw0QL303yDoO26XbVKdjQhpk1fLDK2I862BEgr83DPKpEhMXXgzfAnNlRr
AnLEhfTY4KLQBPbEN7xCIn8JraQ0uFM4743Tasd11ArEKUxrzkactBivyvkL
GvoaxflD3rtj+JaLMIt19dYdLsbspb+pYBB9n5iGcSFpD7f8SraKCyDu4R1U
qxYW5hKqfmOamFsF26KLra8r2648SDWrYL2+nMK1+tPijT8vd3/9vmHEKCza
eoQjpR+6suHM3NUx+gVEgQmJ3DL9TmiXlm1OvfKq7pVlWf9tG+RzX0bFAYvH
hm8FInZn2cTw1Sh0f9TIiNvAqUV11jZIdap8tWRNOY5S/2aPOotzrqSgzIWJ
sP+37/Y/z0Zv4AzPne37kENdtJK6yFoQMKP/ekCemZx0AI3eHvYn388kgpRC
nvUOY29/T7/YrtfFDmueeHahQYjWFKb/2J3EHtQPQQFz9ogS/HxToOqV3/h9
YNWOIvVYUzmEi4pgaN47fIuA/TKXCR4f7natsib+TCkIcj0rhGRpcAJx5iae
lfK0oPUosTsQY8x5TjjgOa3+jfrJi5B4wGDZhsi+nyLxabD9TJjnZJK4HjXt
ox58mqlPm7086AwulgshNP0/TeAQ4eeYijSns8VOaaYcWPEIjuTDNTwAy0TS
h8UEHSgQV+Ur+7uNgmMskIQifUrgQT77rT9GV6UtzbvOV3bVEyeNPM4A6wfz
pUV+/ck1l9iDdnuvHWuBve0gj1i/yttG5Kq14O76rmB2f7RQZquYlvHWz717
THZvydIh9AXBgrohRo9dFbF0oeYbKHaCz2mx/YcsbaXDd2G2mgef34Sgna7q
VacNYclfeljx7LfcuwywZPllCpYMUEqIfvO/uBdOgYVfBZt7Teheqb+91Nv8
OVCFIY6QTq3OSH/rMEE+OXhll58j0m7JIbcTvC3OR/mycn6R98VD380fxZX2
nhqVPqnPxN4JdYODC8zE5rfL7Sh3E2123nC5L5Nk+vFiZ3NYkXnofcNj2t/k
OiYVbjhCfkGjy+c3NLStYztqEBEctORY4BZyHw+C3K1vav0Xiev86X00tJv3
sMq26MZyD5Ky73k9/+pvUbLFYBaoxQigB4TqzcpFvW/6kvytUlst7D59xA9p
cPQswm2C7LBQFXd43YMbs0wgmrrxboe2LFlITdfkdZ5otOdIcMbMGg6VUfeq
RHKPrfnVIYx12DVkMHIje2QTxwwXBiwSHDqvpdrlm3dPKk8hf3EtsaGAV5AE
uAXS1T1yT8YlTxZkiZ69wsgI6+2BoetM96Ogcr2wz/wbR/rmUivm6rU8EOvG
s6ZtpEuj1cuOP7zTT9pq1nfB9FmzgelPquMGBxw1qIU4cNtccOklg6LI+kvz
vZTomW9mpvmN85oa2BYiaCWH33zPR4N5wZqCiu5a/Q+PCqpTO0yudq2F7PRu
nMPsKX8MOoqwxfDF3GVoGIwVQOmJglQIJ8hqWJGsEaE5p6FWfhlGvH6NSYaw
b3qgU0c+k6xsGqOQbwXiylER04D3M00Z+oOvfrmaPQnIo3/XRyGjKOK2Zvo4
fVc+mLcMsaMdI869i9k+qHBfa0hinaSs/jwcdfEE3600e4MpFit1CyD4mHNO
hhW6pZjhmpBs+KrdXOSE6hO2e0+KrZG8EmL1PD7F3dbXNAm3YwVHj/4n/f+i
m4+8WXTj3Az/yV2XRkJEz4vdbxV3ecPm/rAOdkoDxel/y85LF0hUZ9QwU1q1
tDq6F/hndzK3t9WCD2xqDZSBo7C7MpCeaMpPMwjgCaetA+Da+oU3RCUc05CI
3KEOz9fbzROOddv3hzVUn17gk/2Fw9pB+W2ULZ1EP/Wgq0wJPQYNxMnebkom
e4uidaGtrNekTm4v9MRQxs7e0nyTIUZlDEI1okIE7mvHkyizmlX0eM5bMaQ3
Da0Zd2twRyfkLBrWpF9QtTxi6DArP/nZYNvq8jej2KfDBmFhCqPvdzjthgBb
wW7WjaYoRzu5s1vui8sVNnnEJnZ8fX8x16sqZEQtHlxDjiNxIeO8263BO4Um
QqyEQRNvyd8248NmQNv6X/IBq0OsntF88KBC//uDYQAxK+o5KZw6InRzXwLv
DXwdO29ksPIMbveMrkjujkgQpwjEuKS88jgU8b3qXOWacRllUPRmfgRXWmWW
BDzGc5ppiMQEqJ8jSFNc6bSHGdLCjf14n8F16fX6VEwpHB7I/TebrfJAHwW6
Idkmp/ZmtAydtPMl9CNIy5g9PTQxuTm63AGQ14Vu5uLYpbJ21Xzn/mvXD+H2
8vqRfsXG4oGvJ2ddoeZsJNCYo4DuA1/fzvkDLwda0F1WPJODg63BNn/XYZYK
NbHU14IPxc7NuGKCTmB5Q1QEBEMVrnqj/oevoURB+p/pIkqQmzNQCXngvY7u
fWOkB68irmzljoqcx0Hocb/epTZoxHGJzBZJOBOhpuk00Oyuu53XeI5UbHO9
yjralm8uK0kXjZOv2DE5oVycXiCXix+i78sPVqQrRnz8qC+YQxJgb8fWCl2J
kJL0IjwugWTGIqBKnb1AVADy7C94mw6wmVbM1mpYNJm9WCvIHQEXmN6OF6To
sG6Gfl49dvwNjmvcjyEFWVy0Rtt9VvC3FSX5XD7m4KM7mdmilB7QXZzCpxqN
xLv4/Bli9p2Ukx4rcSuU4zQqGiFoIeH2CB9p2GCXe8eCxvucXXZ8yGWP9YzW
4N+ZeyqXyzxzh6KSpXNb5BIWr2NSWm3WKUjJoXTazc9Ayg3c+H7F2kD/7hVx
VQczXaSE2q24bU92mCXKVhJ9HEBhuFP1yWnxn7g+3RooTJFlQZ+JPUAeEyeI
9WArNba8zuqfOrVWd5jaj3AaRkAPU34FqEcp/ATnuekNJvU606EjtVcdioYA
g2Y4Xv+s7MBvulqTBxO6wWDAX+2r6CRs64/fg59rZX4chKoj+gQ3EKmWBMNr
ytgORHwJRrDwquTpaAqZWSAquB9AB8hJBULXDXicZAjgyaiqZRo82K1MvT6u
UjL48EPo1ZzavqAwwHTmLqpSKTijr0k6d6C4AiF6ywxDKgA9RU0UB1Jhg2Mp
djzy3Gz9mxqnrTABjRiaE9D71TT0XLnCry3Esjz744obinVfcWXeqEyC81AD
grmkAzPJuedVHQTv8MbkCMWjFW8q6BtU2lUqhBPCNHJKjS7fMWjeCAgxw4QN
N1iExQFjvbQbKFQVX6K9LxzwCM6NnnlLb7SDThMDURf5q2bzKIHQGuZVgpFw
oKfn9gQkAL6lvECBa/cDX3nG6vUgGlyYl+LPIfJ3vBxDe9A7MBwKJSEw7/AB
IxevRiUtjzUB894peTzeDN8kYAToLzaXTT2JenJDolDV3+uCaTKDPIAcRBKk
HuB5Ex5lsMWhExMfavTy29i+feHAJdMGM2INCmbE1aLwdKuJWqjXSjBvYIzv
RPK4v40oSWObKSuFP6RTtQFI6dAk8B5ylmSb2NRnWiLEI8WIqwUspueDLRFs
t+ieGXQztn/16GomQcCMxGzm35Z/1Tc684aQldTqf6VLlq47RXw2hoaUhP2S
u8qPoWCfpH/K1PCVgypMVDvsFQXPs6F60m8lhl8UTqi6ytscPutfb8mNQMfi
JG+MniaUlAqO81T56XhQ3ZQcKr7ItQeATkQJcAnDSCEXipI+ghWIkAa7/3ps
05EtkC4h9MjhA2lSnVktsDauq3HJj96j4HmNf/a3osuUXiQCCLmyLqSIf7Bb
yIpmhbsCcrWy5oyWHmNxCvwfVVIcRPBssPxqspQiNroxRsPd3y12Pf6AfyuK
cQXRPZfeHUNeTXi9XRN4s593eD/OqH+gWiQD5BA50omXjlvozRJrQaYP9J3h
ljEbCirjEsj7gdCy5I+ry4G9P2XkQAmf6nURYic83Lc/1j6oqegYsj8rkZsI
xXLoSbWUCYlTtj7qbEm438R4Ot5ympYdTd6YKM7DbU5b1IvvOV7SMkXIat8g
RyTcp/qQqK8NpoXAzBx1ipNSEtnVGJmBDdh6pS3RyDInwopvVDxiHqJDXYcC
B8CvGo3bXT6OJ18IT6Zxy0n7SOQcCyI5PYNOHpTxOmvIdnSfu3FrLCQIOIMD
KsDUm8dYMtwQnLC9wV9hfOZqL89Xj+5Haonvq72NBa9i5NqpX2RMcx1T1tZ9
76slFdi7zkQG5N4/NMlRNlTD84ggkOvTgWStTEbiMGy1wMfu+V4ys3JdWsGk
ERqVRINQRpcFkTXZvyge2Gxd2uBefQwcLEIq8vGgSDlMWl0Kctpi7b8CuRVX
s73q4dwj7/qcrZydYrXtKPsu6BnQ64InZ1qh1PoKCHdXLLwDQLsuivi9Lj0u
4Vjf9MO8JtOGxOYcrKg5AmHhjNxWRwO9cfh7hlRkSfPnW/YcMQ8XJ/yL8TS2
AVGoPNHKgFqTI7AbkEqE9zS9wiGnpVCS+36uRMbmk//TwNCV4XVwxyy0Lrve
EachDQQXhzpab/tGnEcRabW2Op7Fxu5qIgWcfroIke3QAofv4GDtuFu6tpKi
yJJfN5UE5dmqklCc7IJj+kjTpvKoHMgOBusPRZNKNf2wezWhdFq9roJCPvV2
5t/60jrzv8UqEvaVly92o4h6ji3FSkHuXI02IOqmkc7/wySaTZd5mkxFp/S7
ct1gSdHpqb2HXCFv94AyqeuK+xO6bMg62KfhsRiwbYMmud1uw/B7fxamGDqM
Ra7ZAq4bZb7pVbRCibD4N/NZIKkFXNlaJJif8KmeBu+2XoI0iGJS/9IX2VLr
zV0fxRRWti/55QhDOYCKpEykq/KrxvU3WJ9bWZ9bVwqy9awQaSzYDri4qqz6
Hs4mJ8szr1fBqZKH+EzhuR4p/xfqqe1ixZqzroQ4ElIiRcjTwjPE876et5nM
Ym/6Yw65FLq9nOZfU1rBTjHy8dMZcD364ipDtD/UDeXu0tfW2vLnOn2vETwS
u9dunJEehMfjoR0pHQuR7AklCo1VnMub2jpD3cK0IY64WQ/78bH0xiA4k8G4
SP2z6K58zu8AFqtfh1yra3P0DNXgSorRHlw+u2tPJo0zVw6Q43tsdBFfpTCa
B9/fnBsAAqL9HEX/JMV5gv2BogaQOpb9Q2ju0GzAYxy7cRFaiaEaEFrHCcMe
Hf15oBySZ7CTyHLbZGq71U8g+6TUbIuKM2U1mWpxO6tHEpK402qZR7dyd7h2
/nAwJ7EIPO7DSZxnXdEXdCdx9t5uFMTMntdk5m1UpPYgbyFcK96oR8otWTO1
ct6iGi0lX5AOyrIUGmJbRogV5bCyl8nK+pxRQIbrBecuKyLYA9NejorTGA/y
KtpftXGRsYALDdS+VeOBXk+x1/nnWW8G2eQpEMLX1tr4E6YSfHdW/7fV0crY
v4oY6o/s0AjONGJ0MbNKivgAFG/Atpi+XUXosqBQ5jIWjszuD2Ra3oMtPMdF
6DoLV3CIWQPeVJ7Oc2gjn6jTHujunJUyQTFgz2+iuCA8ozGZgQHGNnin5uEh
g0i7C6LyfgUIaneIPMaG0rwEdsgQAtHj01wK6Lc9I8MmdAVjPiprSdh1Ttdp
t8M6oOuVHUQeDHGtqrG/sKPubbRjo3welNesjWWuMIUz94r0sJBcxbbnk6uz
GqwQ4Tj3yqpp70usc9Enpic2SdCTxRA7QqyBXvfZH26EO5bUXweT7GMAqWef
zI3ZUCqG4IMvqI15hcOURAseR/vn2YGZ98jMV1fidmhhEOqz0lIBu8LLPPpK
3d3PNWn1Mtvma9JuLhEJ2Gcqw8iH4DfzTsQ+Oq3S0DR4wWr/bNrvoaG2jXLf
JkI+t14GAs/wF6bt7KirtIqRhayK6TwDE0ObnjiTvih/4e058Nr9MBSSpshv
Lc7cSuo9DCx5iEe+EnXNCf5uhzV95phFo2iMtE3fSklt8HlgCzWGNp28OhwN
Ki7WqT1hJcTUOLezYuv5O4y+Omn+XXNYRMJcgPJprmBSps7nUcPLNqlamFeZ
XM9aK00/NDwnu8loD2+jXGAoe64zawNPq55FkoPliC0OieSgQuvP1YW9HW57
oqp8QZiTtpefjehiuIitbN8S+cfcj579GgAxvOTOlpzJF0WQ4DFCE/H1To5L
abmowZ/XHtQSIvWHcBnG1DuZ+trxxygsK02XjFaRr7/XQNMxqdnaxKgLisdc
wuO/pKULBFYrNfpn+EdbhLfwqErT8TSFtLOXwqFyKh0sgV2TVv5JvQ6EcYF0
VNGtShWMPwbQBt8Y6jbYovX6UOn0qitTFDjmaZcZRgFcwL5SmHGeeQv6wv14
6wxKbAHIBG8oXCXdhBIZFfm6mCA36wb1Q/DOfX0Kg9h19Ymv+uoaKaFpKomG
ZdfeAeftyar1LorEC2nr80sMVpalu6jvjFd3R4kxzRj+e+94qKJEd56cC8Cq
i6k1Y+pwci6PRXljgOkYTTI0dpfi50GThS/EeA20Rs27DGD5nIURfKeyMcEj
eF7FSgXss8BXtFzh097heLk54Nd4kxP3J+T0JoySVzuYTT+S1rnmNnn+fPVn
ut3SGAosrS4w6XuHPDUpEJJwtrAPMAmEzlixDV5h+9Iq1fBxXKkFF8YnLUYW
R1zC1I5dMqO4GJxkqeEkmxdk36j981Tv8KmqJrZajbyTrl7iT0tzckSSo5Qo
qFK8hflmC9ARFK4aeVpJ4amkrgNO9efMaJSlz6kJnmRtp42LV9b+6Hvg+XW8
Y8ou0R3XwzqK6lbB/cIxSxb/ABlRalZGKvoTmSNXeK3i5yq9YZxqMsKS2VxM
kmBDfHfNF8IvgW6vukdlGToHql7nZ89ayCQVVAdKFE262Ythykzql9mnW8R2
MkAqxyGZ7NDtSV8d9Gp/ZV7MJE0o3yQvIhXk6w2eD92wexeiWAspBcdXHmUu
e+0LlyW8A4OsFzwhWm+t63M3/LvcsqzpY+ZK2JCuRpxlH6OJkpR9aQPyLAxa
SPnO7AikuxL3C79UHUkVu9a+knhpQp72AViRNDyVUNlHRqU23s06FEvhMEp7
xmrFw3UXNCi1X+RM6igTfrt9XS6lnhuyqoMccEG6vCdMBsyLezld8mwQCoW3
j/5sow8+JdvBXOD1iXdo1KbJV1y/nEiu4GEC5qfEfCsJpDrixzvM5py4RXrN
zc8NdgZfAuSF1KC9J+5biAnh6j2Iok0kBVRZO5Cxq9/D0hZIYpCluRE5SVkM
E0Wa5lO54W4ZGEtCyxSyLwx6f2ZR5GO9lTEZPsjFfpp8KBkLLlhTEIylCYVw
yxRJ4V4p5RxP5/o7V/AfKIUKo53QzDOPAvxaymDuCNuVAij/odMAir0Kbc5j
nV0S9lpBs7q5ztBVKVIqqCCH+ITcDcXV9Iw7mwHblqHV7pOpF3wltRAPdjGB
MJckevjfWo2rwX1067aq91FHKIZfb8t1FAOho7UKRmgxJYRGuhBkf64WKePn
nRSQQek4yNGaZwp3eYQzn6fSlfmEMiKwDa5Pb35TPk/1BKzxmkddMX277U/O
pPBz6NalXFl+SnbpcC73IaQRmrTvuh+YA4tRCLl39IgJEeXnRUxmkDTyj6EV
iAhQRYW2CM7WUdXP6pBOHSxXlb5NwkpaIidRu0czX0Qutse2gTmOWemS+q9U
ZvTwH5l3a9dHLatB7PiQNG+vFcIh7gIZdr++UKvxoDYE4qPyUmBvw7RkpJtE
fXHdQTrjf7Rx7MB6j/D0omzSjUQrfZQbO5P0rbh66isxkPRfGEMb98qbXqSO
gBH/XKLaFE1n5EfodnwQmmxHKaYogbkmS7jnb09kl3YH5sbSc/+PNqxtueAM
mciqV8RJlSrH9NFkgvDdV+jg4LrDHrnXkrnDvZDCqP5Nw4lGnBvP2dDB1stY
n7XdENJ9Am22qJpDchQ9W3C+a48hf/dk77T25oh9s2jcmxzTw6fWQS2c8FdY
lqBSkrqysQdkBjLvD4RCLK1kV/HKvUX0Xn2QSYfF98RkzfwVXA/3D6aQK/vO
ulfFxBhkhawdoPjtjluNMqoxNvegjiIBuDJVGJPF0PD8655GF7Rl93V0aAmT
8jsNzEoX5KSoT2JMtFCFrL90uTznmO6spJpPXqrz4MI65IX5ZB+ZIZGHUhzl
FqTxOQSVkfmyoCRwWa0HG5JDugagjX7xnusIbHkrurfWYhLmlrP2po3ajBo2
S5AiH6z06S6WX5ERSTiucr2m+M6RGJG7sjW/vKTKMVt9dAKSSgiFMdUFNKh2
B5Mf+dwH1s/vHWRKxjZJF1i7SlN0LOvEAkdv72OBHJvjUsJEMG4gJa5/G20y
GaQ4J+h1Zh9qEHPi3R0DBpofonKQy4JHKPcH8r8DgKTyZyJwvXEQY1EmZg4n
1xcjDsYqWaEQH4Z8b2jfm7MLPTeBAhOzUGa2hivNsWJc99YRPCVKWc/e48qY
fr9ks6wIv5/hdTjufVRT0iw+j6Z/vMAJGtgkvi+kekuSrjgpKJ6dPJvcM6ql
8LjkyyxgE2NUGK0CDk3enDmoXCc1YJqznAAWVwXz51FCf+Qq0IjB/ThLESDk
1f+ielapRsWTxvupdhqNVwfJa+ewsrdPnHMo43rSek4XM2AutANGTVCnCWIH
MlucXRvqb8V13VflyQwOJA5hAt5diIFwSWdiG3RubC1udfVy6aLedRk3bqbm
uOLsaG1EWHuGqr4aM66tLATbnqGoB/+U0LCh1DZ6lCbPqGC6tnpF6x4VMpnC
xnvkFaRhlsazvV8voCseO5dMA2gpB2IEGZExvtU79GVr3RKbSWKRNwQzw7DV
yqDRRFczd2DxNL4z/PzlbafYDZlEPR//ZHPA7MMuWctv4gHjFEJFcbeHrqYj
WHJVvtZlM3vI6RD7hhIZEj3MbWkUZUsL5fwOh412cqbm74xpATxcNv8tG5bB
ATuhaTSnMxcn82ut11buBq+kmruec/tiu4wvW1jCOIZoaj4TgmhAlQ+B6JOQ
Pg57+73YvBxHekFLi2Va8ydcV+5k7pTc/qkNMjWf+Jscee9TSkQLRZSnI9R3
W/FXWkG3gfR87QzllY2i3YYt2s0SI24Q/1hqs95YWJodGs2VGM5sdxEQdf8M
r4g21lV9PBLKiEVKYRB4/iwJRp/jEDaTGsb6Sc2dw9RtvlkvkGpzXiv0my+e
Fo/x7eALsXVZ1SLeYqBCqDOGTZzczUYgGc0IVvjicUMkAdNMYOAi8+mg8Adp
+QFyLTP86cd7Xs5J+BTNjiJxuXfmqiJ1mJws3TvdNEoBi3L2pVtpeDm8CcNB
bx5YnRD+JHwLWhfKdol9VqcPRjfXxP4P7gbG2SLnBuOfM+0Utv+SNS3yk57z
EEmSH1PSBkO+aPUhjeiXVcu2jK+32tKmOqwQsBHhiDm3d3DcmGPWmwbzQZsc
feP0UpnlqGAM5t0TPxlDk0rRPhqvlEmAgsWe26LVevKGjibWSN2UPGkk41Kz
rtzA13nUdGx406es2j8Ei9ZcqlFhq1hGSE1jmjTcgJ5uVhqy0X9LhoCqMDUE
reYMmgwA6Aut/5X1UFHckYFf1GukvTeLY+6MyIGeMgwOIxDIGKtybo4SfjzA
enQ9D7Oo2GCTrfeokNv9sbyM82rnaYxzn/GQUlDftGao7DfFZPhBkxvMZNZy
G4JL/q+a/lg+Qkd4a269W1l2JuooBwathbC/77fUHFS0bopBoblL82ldeV9+
0nMUFSbmZabpE3DXK8AQTBcZvzEzCDlwj5MRqld0Tv2P9DZxBqln8xcEVfKI
7BRpPsm+xCW5RUUqdAL3+wexvPlIyGluKWHCnUGBAbKS8zP84zRz2laeNvg8
8P7f76Y3xwHXi/mJ8MjUVlCRMJkzV0stUMspo9giAPc0+g8vP218Cejm//a8
2S3AnEgOQmpxW4H9ellBllm9x2AxpIZa6uxIEyOrw31Abu680hc7RZVbcqf1
2F/DncpKx7nHty/t7ODGAAZE3pB3KE1awXWkiSvqzIZ6lCTb2FaubpkupTqP
OeY3J1QGFQ36scb886MPSmere5p8pXU++KJwaZqJijkh2SpwqaiaInWT5i3q
mUO05wtkc0M1kxyzFKtNLpNOqv88pDcUiDUlZiuhYSKpqBVl7vhXVKfShEAr
ZeoK8zEQia1PfzijuiuznqZV1a/HAv8JrTmt2yiZMPqLu61pLqCNAElwtvTM
8oLtaePZg2h+Fl/Eg8tEUX00Oiywjf1q4R52Clff/nu3AxAroSRCabeOD+7m
FuTD+n+ezJtENIOkpBosM/SN3aYx3YcjjAH4v7lMyylz8qqBTKFv4/mMh2T1
WI1QJodr/WuH3WY1kyJcbAs+oeI7vw3W6/9jEb3bgquu6RXJPIit4OYRt+UE
PaDG0SIg9PKikyhM4IJtSQHnz94BfAjeorq2fZ8Hx0g+JVE1KUEkwt4LTj4l
Bszl2dQheZGNCvhL2h3quJ62jRU0sj8ZSpHPCIWNzT+j9cMt598Y/yShegq8
Nj2dCxus2wTFvv2oqkIjo5OXP9WXt2DHc9hrY0P5b+q0ScboKz9gyjWSWAXH
aexcK63/qifdMKZ20m6BQZJ6MYCKzRDhEaz1OciI5VNRLNQWB4Ebi1lW96Jx
AxUD5zXYrUgaAxi0ymYIU3o0HkG6VynDmdndPyaUWXnAXSsBaIRUYmRYOcAE
wX249eleJnlNXuh2JBRC19wFC4W7ADopr9TU9czExANBDWgmsOJvV+P7OqiY
9vF10l/v1RVGTIuvvwxqE1M7dpOPsG4BpYG7W2HrpaOvU1I5IovSrnqj9q3m
YNrHY5G+bntwcoj156uje6Jfa8DxJTw7zFtFgYpj6Gd4It8shr4AnyRjCKez
jKgqVXUO+xoaOlPnQxJ21ir0wnPcsoJV8OOZWWT78YBKwBUHSZNO+u49X4eL
5FjxJnU2AdVfcBcIYVmdmWew4krVWFq+c7kCaro0J+7z7ACyFNDD8hUGcmOR
IYuE+egZlsRAXMGIJkoNDz14XYDfLMJD0gNWlFfOED8ToOQeZ175BoagrW7+
D+dR70FwD0GyXBARSv0urdjC62Jd7oqB/08DwCGPB3vCp/ATPnCkk6PDXgRz
2StYj9Wz1i5r7Jv75bef3OVVu4ETomQpwfDrvq80KwaTKWfBT9KKdAgi4bfI
P6fbcQsJt6oWAxj6T6K1kN9q7V4Q3TDpJRsSXXLFI8TKv0ly+G51vTsGV+ef
i34EB4MXLaXjnrXPIruU6sgVRyp0EMTK8+zTJfJtBjqKgLdbRs0b3mazS6lt
bO35sfEeVE+gmbSTHZeY3Hw0pd5sdtsjVP699Zg3f8IjYjl3Alpvb2rg/qCE
TlUR8A1fPAdQIhQLiJAGrdBWgqsCCLMJtawiYE2pD51Zcq01vNx7BDK5+dae
3BjHofe6/rvIrVdcxKJSczEc5OgtEp8+EqkE1prjNbfx7mHkV5KvoNIfIqgH
KXJnKj7WneNZB6I9IvYlj0e4gUDUzLSA9WwByWyvlGlpkj4G8+MyROThIycf
sh3zW/+Dq++sgRfLElro137vuwmG5HkhjVJaR9m+Jpz+e5J7hT8WYnbAfX4o
Uf5dlaEHPlhmFAQYcSXameGNxmcam1zl7/lqZpKdWBVfZIdLvU2UpIkMqIT1
PQ8dfJeT2c67XUNCRonG/3Jk/NAdaGtoRwSeSKx2f16+/aa8VfdLCumDIY4/
OI17izwnh8iDeYqOFRM7AxRo5agJXzl6qCAFJykZqowdKsMDZCKdt4f4ysLw
h52SgwP2DRr/PrEVP8EVBg3EwFvdoApSZpBgCfhycUnNkrQSH5xwIkqlCKc8
M5t/Tp1If5DpMp7G76F4ff0Th5a9GyQAtYq1vTKpbhQLAYxGGhhoRWbbs4vm
4FbTQSHmok5ikJ6/b2sFnHShwacdM7tQltO3Ba3rdhGUpgSCU86EQXSx4Ckf
5XfvX2n3utWZ6wm4Tg8HSTJ7bFv8PC/YANyVwfUDZ8F18gG5W035PLSIiiKQ
JVEee6mIZunXtPxEqCnvFCZY3+hTM39fSuO63BEg0EopEEElLyHMO7oWqlX/
syyj4djDawYE6vPIW9dTpMVCMLGZhtiBYupp4xlRJqVK595Mq42jDRYR/3J8
xV0fM/RFlJT/oZOJNxkkJC1yqYS6JU/nwaXvJGbkjfJ9uveJugCaAxgxAcGG
msvRT6wF8LijCl3v7XVg2HCCFhfHKzXloEYautFOda1SUQkXF1XzP6HIYM8z
nvx4OWT/Nt+CRKp42tJAEK81/wEj3eSqLfWPO1i2Qq7B9phO/ogKrCa1ev6K
7n4ciCWBH8O0ws4anYpIfHIzEdONU+fnhrA6roJSiZUbLfU0HyFFY/wJOE3c
YjFCTCklwtr3lL79Z4KNc93pbHFb8SBajxl0UoIvUoQLbNW3GEpDK+OJAFl4
1z+zGI5RIWVXA1nDV+Goec0lY656dgeYl0RThoq2vejrXMZzJzbOMQJDeMDc
HmynpAeiJaYkXo74sw2PWv5jKrqJKxoZ2OGzZXX5NKnrJ9iKQf3GPHUOYw7x
eAP/T4r6X68rmmmNC7OSJ7pQ5aWmvbS3EorqbkfTTtZ3k4xDvKrB278LAKoV
cH6s/2WCAqGriXkcQJLpMwQBepLP1MmVe3lTMfp3LT7qSnln0z20yC5yLIDJ
Jj7HCCv9cR8EenOKlU/AMYLHImrzijO5xGgp0uI3XiZhQmqshNYH7ofU90HO
ovX0RiJ73Cje9JtApnOiF2qJ6DiUzpeTf/X3sJmYj17Wk0cM257Yb4VgUtMc
Q/1kjVANH2OpRksUEw0sNOcvvxlZmRsjKy5+eueh5a03y+jF2IFT+00h3E3z
0/HU5k+DdkX7DPPZFdEmns2VPoJApQMCmAvAFhiy9d7VUdGD57/sCBJ3B7cw
YqcczXlifWc0OFYfoIcCWpzDgjVl4bwt4c48stn+8eZBBIaQPcMzQCx23/6P
JGgInltXy1F6UMhYeh+YFE4qH1vpwrLy3Do0fe2W2ORz4xaWY4pk4/WVAebv
pZjypm0Xnz1h5xcDrsbe9OFhalMZgotHiuUkzGhCIUyGA0+9wfs1DQrjbhL6
N2n7lGQ7+Rb0e5GmZhGZeW01xeTPSlP+Q2DgX5ncDvOyRoCGQENkeheUFBZ+
Atl2K1hLwH1oYzvmF8I0XRlv9sTjvL5PBiDdD6yhTGL5gT5zcSXTkzjIb8rb
VrPY1hYmY9eLOIBaTwdcHwPEe7JfVAoTasyik5mQ3wmwuZAD+7xLuBEh/pJh
BWmp2bZG64eKKAj9QNF1e2nPKFAus2sAcisrhzLWqEENproPkktZlxbM8lbL
JaAOb2/u6W9GcqBQ9rDCmYwnGZC1u+P7eFZ+UmxrQ/uIVjZPEIRYOc77KbXC
W17pkezkBbhMgQaz9MunlYJrvtYsX+zZuq8b3xqhlBEhs1XUFPMB4aYbP44K
kyfqDMbst12tMaapXV9XLI0TTN4gXoI86naoFECEGu9PXZ1W2eAjVaDrRYO8
N2JspX+czpw7Rk2tVNPxhyFdP6biCehFnSQ74p7iQM5j9Gu1/XnJc1yTlu+9
CDDFHwJQdUK5iPac9wh4sQu2y/+N+TIz93VolHTjPgkW46eAyIxmNyyXbtPj
sCF0XYk+MtbPrmy/VP4JbUmuffPTjNAMCz85Z+KRPcuCgoZQwWGg/w/aQ2aB
q1DhkiptUlBZWzCZ+Xa/f5OlYF7bxRX9dvIQIARkuvr1fWCzw7WkU1MxEN9p
3ewwYfyp/mx6lbW7sY1ZlnJA9dUBoI9Kprx4bs+uClkhLSn1WIpKmIVhFtXF
+RSBMVoOwr0dKO4u61DgWjYPXjROQH9zgex3RDvI4h6Iz2y1bcypI9uIRAQ2
nQniiPVsdzVCj4b1hr+7a6Cz7yjolXgdGK2oy1sM/vzEuUG7nPL8LND//KPb
+MimIkqHk3/V/y68IPoMnaRLXRHzOAGWzU4sCvFhaG62gLMhebb9tVsSm/X6
fC5gE+44PskKTC/fK+wAaPnChRIT/27wQIjii23/hvwvY9CIUQw3w1tISwTo
56RDkVzCg7HkoT31yZc6KLN0lP5ppIhvvSTH5juNm2eral99s+9bm6hLZZWs
WfVW/rfY2LUXzQVaCpF5vwFj9k2AtFFyPifB3pNP1GQ+x8o5PVBm9OwCtGJn
0Vu3l8VYMENCfIdXlVl+x3X5QdgY3QwjIjq8Qx5te8vz88hIxz59HRG4REXg
cmKJcPMGir+meMO/JLGLiDSzqV3TM11EECdUGsHx9MBE44eHm2Ry732KW6G0
NPbRY4MoOQHDZSJdnXZ/SxkW2MiYnNEQbsRuLbIP6F6Zc9vfoK4MqaiDaWyw
J2SVRq9ntRA1XJEFQnu65V3Cl1SDvjJXDrMI5VlUE12P1W6Q+EPfuZF0hO/j
SsJM2XVJJT6DNVwAA2DKi4jt+6pD2sqbIx9jXMZS5nndkLLcrwsI3O8LFhIX
eKwTQZmSjo6Nr65f+wg+taqaZXNuZVNBnqMCEsZq1CICLk+YUCv4Yk00OYMi
pfAkhG2UQeE0DuDfFJhCZ7fjHA6452iFvmFbNftVr1i2pORFRgjjfNIaci6P
AE4f7PSJPbmzHnPsHgKN/WCgZIfZ9f5rEOPTLPYPYG4+TIa0iHF0ErxVGF3h
dAsFAWgFIhCgQP9bTZtWKPs6pT/+HmNrWcD19fbV8CdX92kGUeL6VSwlZAHb
KvCrGCeEMgTu4YZ5BLQC6P0jJ4+7YnF0o5jAPIqysFQK2riOryftuC+74t9+
pSMmioVIkzHwxh1X6hIPr0kqnf/JD2oCAwQACoH6auz5lFpie09VslHVzilN
3qK7MztbWHQ6/tmwdKXkEk/rXFWNIOEmDawpGqhjOC9IUMlc3rvXY5LGKCb5
H6cx7Nr32bkV175tU39qJZJ35Jm2D9eIzHbloMoDJoXJbOAazNmb6G1c4p5A
xlxsNy7R6IjyOt7hIRrTumiiUT/cFPuWYPmM7EmUazJhLYMQCzZv9x8JWdA5
YIa31qQnlAf6+t4NoVO65Fv5+wqI3zrvXZqB3hUqhgx/JGdoYxSfO7wOyZNU
OVElT6KZZzdcUIv459rlk2X4dGdYySNy0lINPkDZ3q6aRKjugTIzTZ9n0SAD
k1HznxoOvxEhftZfnqSU0518a5BKZ7d3BOwQYJfFXVXxts1yClz2pBu9EvvU
5JINhUAGSRoA2x7VPD2+XbnWUrlVdSMVEV92dTS2v6T0pihLTyUYBpWwSp8K
IrQAmonF+f5wv0O3obupb2OgNxk7E4YRzRLTwONweWi4RHJo3JM5EafN6X3F
RIeE2lNiPuQwpJphNwUl8kK/ClsdW5hKM0hDq9gtPQ0lUGnu68nAigBcWGES
u1qhf9LfjW2uP55NRj8IF4Kg4kQ11sOChLwfeqm2tJ2vgi8UOjsfAgVOJOw5
ctvzsZmIHnSMOlNVnGDbTZzK/WbIVQSk4QbDod3nGg9aUuuHc5+HauEeu+cU
aOlXmm9x1YdHQI2Bp0gbF5KIZHTk/2KSlyZudj7hTEhi9J62aDzaO7HGcnqI
oLySSZdxZv3vhFS7dY7zlq06jfLnw0XaOCsaODPVMAgOuGTs1VTja3fXvFfk
yamgQw0Nxtw6qSc055vHx7TtGX18/PjT8pqXRSTUjbAU6FsXJDjYd8emoz5c
7YkQpNl8P8gIFurEqNhCs75LrG1ujP/fPYHvebJL5q4h52r7HVk0HKqKcDCj
FIaB860f0SL0Whb+mQW2VBkgG2S8L6IeyVwINe3ZvN6nnqEUSZsR/uMCBLxP
Pln6IXV/nbI8OxOx7iOA5AV1S9AQyqVnHyMJix+yUm7+L4HmyPpiWEtiZBGL
zlUo6edfrjTCh1DjoMpNA9deg4nOq0vaYIIgMtXLmFq/8phi6knmaYyztfDi
f2Cw3GrWJN5rZg0ea+v/HwNpgPKrzwYdfl+dw9wfyum/HPZOjh0mKsDEE4GX
iFsDORpOQz4xY6337LaaeWolzKjn+pOck3hXqP1VnUA3dw6+wOK48R94FQ9Z
zjUz8HwBZp2WLElJCrXCt/Jp/4UvC6fBdnnZcwjhQJgN4nc/TUEkWoO2c4OT
hD17Vqsu4NsLg8Ptr1JgZo2zYgNlap8anOicLQEwgJdkSpJi7pjThWr+h20N
cThzDVlYZdg7glW7zKRRZDpt9qd8AVOO1iYyFUiJIfTGkLwuclOwl1Oor/Vi
KQDQfzB/tss4+C1VE/sdFaYTiBOVUE6KJujYwASxog9b7d7+6Io8BEK3RMr0
OhxRA2ES3kiulBrOF/DtFACNNjxOMSeGp1Ef0x/D1WFOF3PnUBCvCkGQt5WG
axUy/CCmeiFVPwsRrZcedIaWzDrqj6xhAdR+y3XNLYuj8h9DrMGczQky2kTK
qdikNS9cVY4rfOui/QLKda6L+/X8Wj3DqVOm3enhY4Gc1dZVQ4e7yzNcavni
7kfYF/8JmBUaJ97lhEFsrM8z/zfC/2MQoyy3OnBRUd7NoHW+h0nGmtN7LmnC
qakdOEyLGWMKN0KF2XKFNcFWXp1QNa2iAPon292MPYygDv2Lf0w1sSMSvpO1
PGO/UT/ZDw1RalVMuJIp0fujJ7MhMTbgagKMoJSyxXQtMkTshPP8ttmjeR2w
+Bph6v+W9N5yiALq9UbARDoyoQFFTgpEopMxzW5/DepQSJfC78EdBUBcgFm/
3ljx6yFvMQebYBkRcEprGoYMCaWeLe90lcQHfj5UHS/fVNq2UcuPyyL96SwB
99gcfM+vEYhG1ldaTipXNyr9gbVDKIEICRLMkPGNI/gUhXv/sjs4HhdO+omH
HPFVGgdFUqYqH59MAzUFzr/AEeSqrNxnFcCG9pqie+nn4RSQ9Iap11ICofPg
3KJNDOLnOltMltS7x3lcS4hfSUSMshxFU5Bx/iK+ncSWUJzjYzXD4SlWmgRB
46JCYiIWQMyAC6ku9q1gUjR19So0y1xfOBdxNQzqcMFo9ZWhFo8PPjudy+ib
h80FpdpQXY/igcB6V7r6NzFONY3DV5p6AWv5QPJwJLfF8k9/mEPjGLrzFjAE
1PX8xak+J3h+tadcqaU4vVm4HWe/t3bx727qLcGd/8tnXPn7kPzyGTAFIW9u
S2E3wA3mV8gPGYtFh+f/V5/ux81CJu3uSSXIBzm2q4i0JDjgt4BkvqXMK/ix
1PvVUUN+H56vaCSs5DiuIaUJMLPdbwWyykAu4gutmtjChSKe01ez2nOxIg7o
+WOKsElvVUFuxOOK3x7mrIVS1vsG88RsNmtSv7/QhmzNnEv6iOWrlYQG1JNq
MsNSRsQElU7QaHQtGX1xc0PJydOIAc1x8J13K0Xhu6ey0vpnNu0sKNAzKUzK
uenKsHPb2p7WDOdHS70FqffiZrS8roCw5CEf8xfGxmd+WQ8/SkJBwNf6WLqo
uTaU42SUgUnprEYyvuTIl/ENDxm9ITpcyNgi2Z93cE+UogLVsvaDltS5ghiX
MbdK4om/3juabx8O/brIakL2P6DIBXtE68SElS1YxHGn/r8s3oDL6qbwowKf
YLUfX1YCTBsyoOKr3/33wY7RZscZpw7/7Z7o/GDfV1wgAwvsXWDLfRuJBXL/
IhpJQVlKAiGmWEGjKwxo1OBASgQKM3k0wdT+dKeSJAgsWrunaxhxLwYZ5Fnu
co7wj+aEQ5x/EtY7arNifQAf9N59G1j1GkwEnWyVR3MIvsEPvPuP9aqoP2/S
w4CHLYKHeysnBX+CNCj+UjmcXVs/XPKk8Rrld8GuvwtjfYaKh3r9x1NHLICf
Mdv1hTfyEmE6VVyRtVePSMYV8rN6fnsw1fVGPRseUWfZr1e1H01lIB5JiKBu
HkB3kWiOBp9zMzmTfcpWDT3rAM2vZZtu62D/+1cjsxBE3DfGam/pXR4K4476
GneQw/qUHN0dHWLrv8G5PQRZjzpxhq3pRTxop7alG4QBY04dEgNGW+tBbyHE
IELVyB15i5MzW4nfgdYKReb+acccnuYC1zlmwpFYNjntm4zF4LV3DKbOOC4e
tGGRQCnynBdAY/Bsxx1dcXx91cXFKlVQsRqo3u77al93XApJ/ibQeuEaqn/k
dCWA2aHV4mRlt8AbWinWILoFo5dOv4xQEyKbJ3J/wb8qmQOyT2qTJ/O4hOOy
l3M7PS0ZX7CjrqRp3NeOaK4LTy5tLdHBQUwcUAduPAjQsBfa3LBjgRd2X0s5
w7pEvXAocOAj+m0WrEuddC8LmdqZHZY+V5bQKNFQ6xrdjWMIqLSl/5NjQPtu
fOXGBIiXm3AWlpjnMx6fDnuKWEE7+Fi/zoTDoWBikC/QnaOFxe/YjStvg9Cy
aVxcozU0otuCUfftDOrfN/8yvpS7RqOogO5JbsU6Og7LIVRbja4LT02hpz20
ZintIT9oAFDKbPevWlePxvxyMttoFjEXZ+5LVfTDjPooo2u7GX9de6+kuU9+
6cehg+zAdnl5zRyYl8L8+zIhF+fCrQqX5Y+0RaZQkenZbGTTQlosuTxiKgoQ
4F+G0zt2HRYhe5RD+3wA0gdDURQmrZb+dCFYRNjeMPG157dGU7JGnCNlmTT1
Y2y9CEX0qGiWtSgWsqGcbb9Stf/ER3iDKRgOH0WhweQl3f1ZSpIGiFZxaxuj
PO48XmcnJlH5AjnFJcMskvpC2nmH8SZnqC/N6UUxvmDxGE273rXo/pqd+j1l
gng25gp68oiPF8DfEtX9VhyWNEg2YA8IXTTXrm8dxSCX1o43BvM7IZg2zFMI
bmluJoW9MYsZkieg7xsjJsNyaUCb+ljVH8gQdY0I/8f7MnyHDkDtzUGgSJLF
He7q/H+jjPMX70osZHXkWVlJUqSuVl+S/y2fthib4HimWUzKmEghFEG7dmP6
O+HG3wbvkL1zpaUGPRoUluhPbNXol95uS0CqbTt5OAproTE6ih0yuXpQ3Trw
ZmpgVSxfhRyC2nqmv6CgWvXx9L3ZOj3BURQFCeIUsHdh9QyXcKiPliG8WBZU
1hDO67Bs0ADQLC+dbp2rdHjFpc+NVYlxZMZla4U8/1eCKXhfj4iOtlClTRbA
qa8168nqLwnsvusO+Oyel6FokCr+vrxQ61GFPSuPuS9mpz73pynMfkPHIGkv
Tp8+l22S67jGL6lM5QXmzglvzandgEv/PubL9NN5/WwZDqR/9GOJ8k0u5irW
99B9gR2cNu0N5hGwfzKP/yy4KiTS/Z79QlGgkQvTFvLyd8sOC4IAfo5DC+Xy
vCXOM+21qfzIMAyRdBFSlpWr7g/JoK68Z0M6gy3zhU7b89V+vFSnNDvSYBS+
DjxQg9zXAVDtdOk5IzNpxs0qHPzFspw02q0P2LNSNFcVDLKBP498Xg+g2cU/
2/tO644HzJ7ySogDMcj1ZZfBuq/EW3SZZKddjFI2xMHmktA2/TRjM2PF8psb
ECg6FERD/9H7rAZD6NnVoK/V11l/eI/2kxGBM12MfX+qFHZtzJvdLJKhCsTm
E49uFTXkjgf6F+agQ7x+kS+BSHW4r0xZgaU+hAnaopPDNhB6hWbisGhcJ7B4
cy4MkBzZvknED88NwiyiI5o6cW7FpLa5jHUbK1oIQg2HO0rOBycOclHxA7Fq
96oOSytXz3YNFv0g98m0XDtlmeaBjsWTCnzioQw4etPIZTnqXFpiAmmmGtvg
I9qlRLQHED1UOBvqqzgQQ1+9mdCO/LqJJ4CjBZPYWJLtUkI41ddin54aL76Y
xPgrXKd/RNhOHHZ+az5QISNOsirEziF3AD9UtC1rUM1F1JvnySoQ64bF9ifi
Na653K3yjgod0Bf8Yg0H1WdqKPHtQEZjZYZRCvdJcE5CTUXtOMG/JleL44+B
mgHfp08X19IWP5guiTytrW20BxPhIItHnDmiKmbl4yL5jitCGYbxuA3cx8qt
FBlvsZvNfyJEsVRAELXuDJrTzoAwXSSShjoc39vaAbsT5rpyXvMBp/goamLq
aALodY4G3KwvJRwgAZokYU9umngzPdJxjqUFRdbNR5NG5tSCEcVIP1Eni3Sk
EAS7vlCpMrxQKNmxIuEMHorQIYIAdG2eLgE26RLvnUaNZZWlZ3w2lIqjVSEJ
0+ZaT88f9nFjs2GNMcVXOTWRGjRT3NQDn7jLei2rBic5cSMWlJ3WAHaUDBuU
xcEtsn0COl5abnsP+w5FdJLX7WY+iZw1GBOuEvIzy9D2tMEZW4KlCcM/Dw/2
4CHoRYJmPlV1Pp6BbpK0v/nUJMMkvFIuzDtlDAYM0mbUifeqNfZ3ZP0BEcMo
kkEgF9sT1JIrtnb435LPppU5F78pm335o4MHuUh+17jpPbmoeJU11UfBpIwP
h0xim5N6E6bxFhWHvLh0o8Fv7ay7COXHusdE98Lh/KdyB6+8thYPeJn77zms
KU/q4mbij4jsq6DCNuILWiOm6+qclDthkh1YmDK3c0tO4Z54TampY9q7wYIf
G0Gc7VC775DmeladKaYjOSGCxicUkgQX1iBgYi6HbxI+msebzvaEVqNQsOOL
6NIUTvdiYE9X3cDFj/bIbAL+4yz/qxZvc7xgzMpNpU1Dj4Vqej138xXEjM+P
SboTvQKByLQ33h5GsuZINadoCbLhWtmo1n/qJEafLxkcO2Y4jueNaS38hTvI
lQ6jb+myCsKR5pegsIx1ALglI/ohKnJWs2fhvdRPKlT2+aQbG0Cwv0DYfyqK
efAYac/AAPmps9H5YnfuGeGlX5cE4ZGDZdVRb7e8lZAXLGC+QECNNqPsbwx8
IDQkZQV/rHW/nQTtTY058NBo3fMMDZy2x7yNjaUqlnXzXlJ4GhxVFjVyVg0T
qzucZ9w5VYcE0nbCFLtoaGIxFbUciZvnhM4K4rmUno7xhtyjxp7B5si88a0h
U07ns9/JQujIUAEdkZZdsWAf9DPfavViGWZJcaxi1hfnxqeDugW8UMZpdLNP
XxZqtIma3OFSCq+kziHPBmA5NZ3I+i2M/1CoGsZylIVq0j3LMgMCs+kDGEyG
vIqMLj+D1dmeC1pgDH9mQzhIYrgxD6AYUWJjYJeBdvM04G++blrAueatChwV
bVuDYS7chiOKcU/09d78BiE1NUP5ErE3we2HLcHkSB2Un3oFlJMt3lbokyAD
AtmW+PWPfmeWx1Qf0NTOsx5k6++0EZM8U/H2nv1cTjVu1sJEISjUrQz16j7R
Z2MhhcPl50jW33gZdNBj2KZn+xVX42uDG+AY+2FXKSEbGbw78jba7WpvMv+I
ocZnPi/8tUOMQi7CHAic0cp6hxcPuU67eQN37waplq1MmVtXv9rqCOrp5kq8
u1rsk2mlT5Cix5Fe9PD3D9RtTh8bpoiSTZafHEN5NIbClCnN8ndY27L9NO2w
a2McyDAWK1xcy5SbwT+K1gkBj5PFsoq5brOtNKvyVayAVG2L5QqHh4JjDhCN
Qg+NWZFzMdocOTQjmR3g1wtBofYy7G1HSHr8dJ+qMxMIrmiogVo+E1Wjiasx
Gn1FRXtueCEmk05dUhDbbetn1RpLRxNPdSEMSrtBjGcOl2O9qjIbr4Uuxw0o
ZEKG4W2ZkltWGJNYSYhYTolhEFEfxq/HSzxZGCgsjs2qoiffk/aKb0ZUHzrk
VHzEccyjHEK7MQYftnx9VWoW/wzcnGOjaX0motwdjd9f7yS2hlceJrEh2qhF
qbcRJ0LQWoiDPYcZhgELr6sRYR29Y2rFGrrcSwwpI+BENK4LtZKBsTY59mRk
2QpcFhhfO+aDKXRFno3qcwjS46m8Kzi6kg/InVOBEQT2+zCq9gROESTWFd1v
s2WtH3QtDCwMMtpyOiE7G+kTQKBCEQt6ObqW87+DlYhpDEBJmT3DnFNq+mzb
444dU8MyzJnt1AhPjTKyDwbtY7Jh/PIpVOAxTEBsCZGCPZ7nfAxNrgl6sfei
H4Aew3CM2ElQFgpNr4KSwow5SoLbQhrw1iFoeea1+rL2zVBFBRYzcW0RYsSr
iLj5QwlBrsfzTdCc/5qrKKPduggKyWICAIv6Bg6mC9FSCzwHG57YBtFCCzxs
wYkWLtwpb1hri+chDLKvBJMmfd3txyP6gH/EtL0ixHWmnTprl+kp96DfSYqo
1ewn2Jkg51jgM8Y4IRROkqTJNb1gy2vFtTTdGLfmLnALIACzSEcvO9W5HXxM
82rvGGfDKwu5R22D4a4DWSUu07i29gC7jye8kKU7exQ+rF2LWqALqK93yVEn
GRAMjYwYbHfI9uBr/Va8fs5Emvo/Dy1/qxCEnxKtufMwhTGEHEDysChWfvkf
rNt+knI7/KCqlbDWw+YpyAxhAlaUsSN76Vr97zqA7Ap3HYwecboHLsiyim0D
66lgzY6hSBWKkj/U0g4ZIn4kjkNfW0aRoT6R6rTPNLUKdhNXQkTysEs7k4VL
ZDKfcWEm/JfoBfpbqNzOH+KoXvE+1yv1aOu6VxF8mYTtTtDjfZ8lVU4ypbSR
Cf0VNn5ofhFnzSPxRmFDmp4XptF3PHFD19EnBc5ahGfRF3VEGvvD/NTKl6SL
YLUMtZ6JbWUTIsB6Xr3/mqMkW+DhECwxxK09sJf24CbGWTArU8QD6SvWVLxd
AnH6tFkr8j79JhthaZP53aNGfWh9OHg5cnZtUy+l6kpo+P0cyEJYEnzVbiGX
P9CMl8omA9xtiV3n6Wz4o60VcGQcrxSmg5RHWesS13pCEwmcJJ4Six1rtKGu
YWRXbMZs9IvPKqFILFeBuLi6haoKnr2WfVpghv8Ie2rZ7Z1906iOerVLQVP/
Quac2s4CSqPxYR+ELblH3G7G0InjcWfQRE79wAEW/ERGaMZVMc/ZnUlp3XSt
DTeehLNUEMl3vi8cMCdW4PK/JPjTlL+o1g/IvhJwR99EQ1BZk0rlEszbx+NW
RI5Xy1QIPrPBd/dFEgEHeS0PLl0oMLO8xMxgSRWDDL+dNBz4DkcfUKlautRf
i0L3ziUI1adYVoh/v9ubw+PyligajcFAPQwL9xlLDBvDFRtjYJSiEzptVBbO
JGRNWDu0u0/S834xhqdbnPe1vt3J+Y378V/upe8kh1ogbh/9bGidu++oa51w
82wUHtvuBYB3/MP7z96gr2NxOZryl/TaQyiwU0rxpOsj5tadzuSMhQqhcXWW
LEy+DLODYTYjxWcHS3grbMuPRgPV3cI/2JuLxZNgfYPZ1aHblrAh9N6HOa/R
dgqa+7Nqncu46K/Tg6edN9HJIKH9zJmWxZGaZWqobchrVhdya+mIytkitWDA
iil1BhRn1KFnoW1zWUshycvfLLAOkW1qA5b6RKrB9QGyUuaesL9+g0CHkgIS
1NOmD98vTd5lwSNu12LQZ5Sbf8xkafr8/EvKJIJeom1Sa32CFyoSb9kndAwQ
ZlZKoASDI5Jzr6P9YEV4Sq3OGN/U5bx4NzX6A4DxFz1IRVUqGgQY7w6gz1Du
O54dXvbBNk2fIm4/yEB9zDosL1gpE43gMVo54dgdRhN/B5zD2S5//C/RJbtH
g+hiNLq8XYo5T7LfeLfBcgKd7qr6p80x5LjtZOjndqkQne6YVq8KSAMNdmxn
2tp/B9+Qt2iDFTUO05CwPIm/0ptbSRW4HbYFvt2kn/XgvNQjBifixIRSTeII
K4kalhYBsbDLo3DeoDamc/iikSDgNZcz8nYjKL2Uu0ykNl9s9zUXFt1VA30t
lMIvekPxNTdLpZxavsb/wL7VHHaB0nVP9y9R2d2j2iLzf8KjnR3fmbnDUr74
gWJD5ss7E86Tbl+DKz+IJUtlBkCAOrLlmRlACa7c9maQkSPh9XaKQqjCcZCD
YEcNx7mhJyXzikdICe0GDkmWBrva7sDvQ4WtOJURQpj5My8gJ3+/CF84ASC2
u1p4OMC+3eVHlmN2VXF65o28Vns0Qp+30hJVMAuiDfNxx0/h+4KzxRvIIk9U
HGU5Bg7dzq3E6PY50i0Fdjm6osm13tdYTvS6Iwfwulvdpb7zLK1bQVpha8Ol
eF/fjS3QCoGiO6t816MuYmzBLWoJIxVGZDGyG71u+Y14ztaA/483td9hysk9
ar/gR3bQEcaA+YRdOTxVo2i9VWeD2TPdc/VSxmMw4C1+lEHfWFKNuF5A5kGL
NAt+GQijISTKD60HMAvjr6S9Pt7TNShbyy1y5cU9iwfu4/xfkooBw3TFnAf4
c3+JJc0eTDAP49Y+nWQFZdUJQuQfRUeezs0EaeOZ1j4MoOa0OA0+DgXhCSjC
2TEu41j0ZpqPRRvfNE7EWaumfLITHuz4Qg3JL3n4Anob/tvll+Q4crXswWFx
TxEPuPiA2Cohsbn81J8PiWPjOgckIZgU4hTb6ZDP1M6mOjC+aecEReX5f9k4
79Z0HE+uO9L5Nls7eqjzpDyGSMyH6QwA2r/DJ5sWE9zuU5l12obUa+5u4RD5
P7QxOVr/E7I1EpS7grGYvs9OdPnGQAn8dUt/vQOt8hsQtPRSYhusDQLRGbU6
k9cIklY/IpIW2lbg0Ks959Jwmebls2JwjK73xPaVc9/zdesdLDUalKNkfUyK
5dC5UiY40CDinWC51fL2tTX6rZ80G4Tr3943ixIsT6tXA7H0DCWeuvgVZmyd
FjamsaMaaIgR3TSjPpeVdefbAC6HQF1JS52zXzUvEZeMumc04mVe+XWgMVbC
IpULSuzAosx2UACo7tyUCobzXsd1obXEm8VCyjBKy+khii0KhmDPlg+nbvBx
EM3VIFXBCUjzsw7XQGaoTfrQkEl7zt5cycDUC8E5FDvqIExy6av/980nSR1F
V1/WV6WKVXtc3CbNBk/9bg6K5Zh86PXh2WpDBZBJE85WGKCthwXSlAhXZcjU
OcwtYgOhIbQW12j/1D88FU8wIpfzhecF9lTj14lEZ6ghbMoQ+YA8E/RilURb
Tf6CvQrmsHclxAnPuMlly8DlJ5UOTlxST0eo0ClOW1YW24NIUteQy+VaPxIw
wnpdR4O7drDDK90sJlXA4/eZNfDbFFESXvKG08/H0M/u5DoUVVOfJIgoCnBc
T34+nFKPyAv4AEgYO/vn57XRM8hsufZ2mNhjxoWsuKE7i3fIu5zFtIC4AuxF
g7iMH7T2zog1AgxCncegZvNoyjk5yNYK1JwGDbnK2KKcWpff7i9KTMzZK/Ea
UJymZh3tN9p8KPKUmDod3fQYLl7HnOjt3A/V3bqb6aDi9kIILTeBSpCEfqAt
BJwEfgBTwNV2TcaqilOpqO3sNYmBddYe7VROAQDjugt91Z3CwPbxNVV8fC3r
RiMJcNrjNiuznRVXWijFyJt3dLIwInN8pvBgf2IjcksC+TLk5+IsL4LwHjw7
1/qcCip25nbQ6LgBa8EwUtzPBD5iVVetYzHHisfC9VL2NUyNzkPEU+cgo57u
aghMyAzCpIV/4PFl8/6vguZA3blXHYVun1gbcx6iKC2n/+qm4dpFGwQ7EMw0
FrfEH2xOGy+PYHaC+p9aDUDS3a6tTmQdz3MXAaTT62cUTXXqfcTAhUANDfTn
gdiyGtWyFlFphsIYqHY3WpiuZbHJ2PXOUryoP2ymTbHwTbP91lcca174Ntd1
FU3WqwkTYDK0w7lfoB0q/LJtA0blPSMKuUeZoh1Td7BQNGTR1ARRbkGrEHIn
vsU0Kv6hIr8St2WD4i1JanUXoE9NDHpkAgcxp4UIrMcsoiOdkLRRWsY7ppKo
UQSwCSmpfrLFy5JBNUEqp+k7fmV5MpHNu8FarGUmDYTkJ67utZKCVaI93IKc
X3HQTOId8DixbGpBCjo1fpH0wc8JN4h3wN8nouX1/HUoy0dOlJWpCN60454N
dFSTPCqZdfw2gG97WsueAMutsGdT+MI55xIlM+wWX9M8fF1OMz+vWb3hGD97
R5nPJfuV+uvyy0shwkrJgwpUQIzihcizkmFZFekphlfzBomTdokxlBy5fIXu
rbW5XrArdr2yT1xLgpKuVc1UBPgU+TBfBTfzS8iTfX5+WrSYW9IIIc/h0W3j
vczxWcMPKtuVRJb8P09KMLBIinn5KgC2lrqQP/NwsEG3645d1u4CmllP6c5o
cvxJVjogL2gxfnOPI5/LDvKmHpt/3Hxv7y8rK2qZd/JuUEobtTKqfme0LUDW
Min1i2lQwyQcnXURk9nguyG6XqGPT3Ysgv4ao1C4AM1b7cB9Rn2D1KhG/hYt
SFGJ6iinH5KknRS2a7rBGE3f3lnPgFP21Ky7BS27E6e3TxdFwhdhbG3910Uo
QtjHvTBYHkCEAkGH/RMLz9wSac/HfseOXukxWofcW54wn0hWhLY5gG5N8Aq6
5sT4Qk0GnTA1MOM63efrx3ZI7oAGqKe1mRP7IfJr4lnBbWcrs1mKYoMZXZcC
oesS2g6YwF63Kmckmz34OdhICrd0M2SezgP+Cn54EGBVSyw6aTASXc4FzBq3
sP+4ftBWTJZ/BuMeSjMeLFPta1uHJoB1wUojPPBeVfZexXgcq9eBDOhX2RrZ
zsrl0BWyElj76HxtwggvJCSPZuGn9xZBzBg68Z76swB+pNq3O9EO/UJAFNDY
aXTyDBEY+J73Z0uhEFEBpEoR0jtqhoNRiszhcxORF3q6Vb9200kTqqQmGe0e
EYhqyv68p+IcTxCmFZiJKfRxP+vvL2Nwh70ibXuowEYWZR/LcPUUTJstL45g
2O2MAhYzWn8i4xJYDwkucYl/gddGd27Ab9bC9du9DnnDwacyLLA8HGsCM+vu
QqkSzhLawiTDxrzwiBZ/AW/N7dea0LwsfSbORiB0dQgSOyytUcH+SOWI9VyG
Fa0DMhnvOWR+qTXula0im0ZDP31TCppSG7u15Oe9WpZKC10AMTxn7JnSdjLT
R/AOKMLoEJj4EguUgGExrfuTqCXoVAzrFGGsog9bOzPblle2QNco1Ib83XyT
NKsGeOrE9ZGz5+tLZx4GpR4VfwwZIwQOwBveHoLl44k4BdI5wRctz6NG0lQ/
z6IKomG7I/P1ZOacrpWH9UYZYH+1ip9k5l77sIaw3vcB/mDEZdexQDud0CIj
2TYJ5s/UXDXPkQ29WpEbNiRZYdLCdGDmsFbDMAPbcrjoUT9NB0doLPaLnWHX
5WDdnAhg8T4/ve/McXjYSNp3QbHmoXfZOjX6hPAZNDV+4uce1SSPBxBEJiCx
OfgpcWas3STazrmlT4MUT6Lax/ntkToNmFL0yJhEU2c9xU76gvX/CM9L+Gou
K9RDD/3r64xw2qZrn2XTnWsKfZzdZXNYyzCq3T+CvPg47W2PUGHwz1ukcMQs
wwVsSbKCJefUccjFCo3iBmMnUohwxdXkHSC9dPd3Ofq7s9+K4Xz6BmK/DZTh
Sf3Vkuy5RRskSB221fqAGjHpG2yPVfxdw7YcjWsxkEvjA6OxFjoBfMv/UcaW
1jaEkZDVf9FQZnWslnK7HC86oLvtSGaIEmpVkYwyemFe6NY/wJA8OaPoyC4O
qDBPnY5XImx9qTaI/MahAPBdjX0MncBCGyNgsUz8Qffb5LB9OE5fFrXg7joR
cLIuhlb3CuD9MW7KImCK7ZHVvIenANC3PcCwDm0cLopx/x9NWhtKp0vX0Nfd
GXmEBIKyysX2MpxLqDHq84sJNTCZ33aD3c7WShX7fjmht81LSedsWT3SpXy+
1GuUok0sUjert1zqlv52FahSpwEsvmgXK2lKeoUPgCpVsyl8jj9t9Qodtj1m
mZeh8f/thdImTbcLvYAHM0OLJHK8MzV8t4lsZYS0CpDeKPFi5qSJy32SbM3i
ZibahKhsSU4nWyeYgZq2hl+ybBEBAfuh8lotDbmB82Ws0EcvtoVgq0SsTMc8
QC/LmXygJg5Z1HiblX3hVZTnHD1N82vh2I0h8n+1F0ChvWmJrDNm7x4cIlJc
LadrwaoboZFb9iUdDk9hVwZxk8rvIsxkLCwgg4CDhY0+D8gxgAGyyucmZDof
c7XXDT8J5gZC5406VAwEDOkl4yYJiedebnSac3r+iVNaY9TSL76UI8/p7ciO
XSK8LLGxy9rdqMHU3ZmF9ulDCzFaeBrlwcWOtxICxoZDv10uptNyZzorFDFi
HHhRRLtiDcwKgTepX8tXHMdr/VNbdQwTzHumULczZMJXxG2QOTMi2xKU66Y9
s+v1tJqrBH/DctVL9v85E5YnpsOsxeqmVLhy9NmzDExQB3QMRz/qdsmVmYEA
uwfTeumfQnlHNabxSC90UGsZ1Dq2jZ0Z26B/lW8kWg3qp2zYFifRzyrKWEO4
Q6tt5HM4TzqW83X0TwjBzTmFyF+QwpKSpiQEllSdAlYK6t++6cBTRpUsNs0N
CVUou6E3WPyKXb3/h1apDXW/vXKcSr/0f6W4scKDA/X1LQKROz0+CPL2QZAR
bicCef6+evNStKX5qMMwPBWA99kQdk2r/nk0/mlt3Bc6pKxPjk5S4gwcxCVl
SrY/hW3metB+0hEPK6lCcWWDXzDOsQyTQgQQE3k28FhkTzLPaEKuvJgNn9jO
aPMPSX/EtoBWEycuFKC3c68G3Yhx+7Ym+IN4ji/Ar7T/31qy5dQSarZ3tOfR
eozny6S4+AgwJ/quHcvAJEY4rtJkko0VYUr4G6NipkM/58xs0MtvySk1PNe5
PVFEKc18tpB2CppL2V5X56aRkXr00IO0cRAjcWhO6LG4oFTWz45CO+mSL1HD
LqkEvowPhg5nO6MR4hsyG3RYxwMijkwI5kY5dyd9FUowm+dzcdciU+kqh5b+
qrmsxPdxzP5eWOPvz5/VHtJdD2dwMPR48QnfQXxsfEkxcHB9NOhTDo/Rxg/s
sm/e0aY7XQj0rvvs1dAcV11+siBAV5esFqvXqFiO6IwvxSVkw5hypk/BbuTc
T90jYIQsTKbtvzPpMhHRetN8W/xVXbwAVAtioy1uwOvMfrHhoEoUDGCShh49
NWsMaFcUmtSiYZQjCj1YzRiT4+nG55Ejxl9hnwJvAIzStOgMcpwEW6a+Vjrl
BDf/zzfPRIdf2sJFgVGQCzYpQIyukaXAXIoNFsTWCQ1wzksJwLuPhgBVlceZ
R10G/j3GAxgbKG2tGsgGKhI5+xB5mE74bF3EA1vui5sVNEejAYGQZO9Gu+4C
NS5BrufaBJaL+QIw+rMiWqKHM/nbKUajBSWSYw/+FZd2+hc36cktgSWROLdY
xkGLacetVerj13TVhXDE+1sBoJu4xlI9NYrgy+nj0gosuMvKMQTKL8de8jwp
YH2QqTioNV5M6a+g/fTUjiDBJDbWb7lnIeaHpbYpWpeHJ62t6AorpA3rUDsf
JDMjcLd6kDGob5vlVtBgN0VOaSgKha1G2B60/8lLhNFX3rj4CKEd7Yx1MI5c
gQAezeTFUTKikSlqZoFIttduho7SN+e4rcPmzcMxLk8UpIBeqMKNsQrFzfzb
mqx8FGMzGUXWv8UZcdV2OC8vc+G2rspbipntrkD+Yh73UuYzuwQ6QKN36LQu
5zEnILubSYFs6h2lwwClQNteEbYFQ1uEl32vgZ4n30Hkam4Vm/Yb/K0P2eDF
rpcjjE9CaXG3zYzu2VCI92u/ghzzXFkOMuwZGGqQ4+4/WIJFwS0TObrTFNBN
1tQbjP2oeCJgwSG36oG2ownCFFBQBy5BCcbmnSTy1b4AlCAgVZeLIzuTQJnn
Bs0+En4UG8CvjIwlzofYFtKpebua6U0fOL3tRFAlb+kaAi+JuQKjCTJ4g80B
y+LHrXmM8t7Hw9Axsp2kLutzjlB3v5dApd3aXeiu+WeTAVG3y1w+stjOZh75
upR65oaBmhiX0svDQO1bmyfZvnMqdCMW7wvyv8kdm/nUHseyW2BySYqvJWvu
OomN1GwRz86TsFSevHGbK6Joh1eqyP72MlRK6Bq22tS0CwZ3Jw9sMJVK9UBA
PRdx1cCItTnoP7JR34G+c2Hl0TlFfeFGLEB7aiLawewnSesk8wg1P8tkUFYt
xJRKGrHmBbDhf5YgTOKcq9FhH7LfmhD7sFXCNxVWuRKwmIxDPaEwc4PLumDS
JeD0ibO02+LGdZWrgyl/JI5ZNgqwv/huHoIdB/9s34unKVXBEiwO1FnDg2bW
L234rpeBwlBBSvO9srSt2kM9tEgWx8v+7uuZghonBb5hNeoux7NItZ/Gkic7
vR1LXFcAyHsxgsValMrGpSWlRoVeimeRTXm4GtL2jOlP0j+BgWwUundAfSBh
556kUsfkRzkPtENjkmyMHI4ifAuUHwuN4ePjg/CLbf82peXRffsqLPU0DCDa
ICfXNU/DKqTNKn+D+mjTOfbfHCFsdgUjiFohhzeEY6tm/YS6W6jf/4O9dHN5
Gk1xAskbGv98zabnOwYpuHZTfmgKTBkXULVTftfkJEIAwsoUoUr7Lc9UCKLI
sGJ5keaQkviom1aML8o+ZEl1JSwt+JJgca0vQO5LUAlTST/X9PLfPxhVcPsJ
n7h+0/qFzKYv0ZSJIkstOM+haWYvZhq8rILCvwUIlxGMSbXV39eJEV+oStdy
0zv6xWQHscqqH+GXtxhFMuNzImJVL4Y37JmaF2nu3+w4dyv7PVpTbrATrbGL
ktvzj9qJFjB6PsVL9uW8FQh3/50eZ5u+1CSz7QQkLa75up8cuUnuDDi2XgT8
2UsdCQaq5pTCjmlkVTQMAW0EbaUFSB1ew0vu58i7z5ys5nESJawwitt8ROyr
/QE0bp8mF1wgHglIDbtXf6/9qchESCl9MmOr3sOxlD2wrkXl+8yaKPt4vmQT
OelZMFGVoR8stE6NvW6kbeJ8KnwzuUln1vskbj2ylATgrs8VLZj1H3easeBs
5MuwsemircV0OYub4jrzUigZFJCh9eRbxbxJ0fostly/xdB9JwmQl2nFuFtz
rCH4Hq6YY3CZ1GIa09l+gD8PAL5YHg5qEgDUxQbc27NX8zCnJSBLcovoRLBT
qUvEhiqXbayIMmELOhGVLwhihPlRcp9bOoakIVfYbXjWfcDkn+LdJsby42kX
w+nsX8uBQihkX+JUniddtw6/TLaAzDfzuXCKYeo0UUoQ3PiaIJXIMxVYBYYs
4BYiBSjDMUMd0xSkdrMvEguh1sVQgnnOt+b/LIfmid7Td0kBaPH4A0sbGZVs
4Nor5Eqn2wYjMgeu9tjVe9c+gRnshIwgosPZ9bAg1AZ7xIBUKQDuA4RxTFmZ
6NHTf6HqZJWQPbRDCodcyAIh2M26vqqV7T68nNtCfbzFMIJwVpW5c1TvaiuE
k741WK3Uwq40P+dFw1DX4KyRniUwdml4zKvMDOMXnhyOfqq21CwbR1j8zOBD
y9debqWP1gzFG+UJnwO3A4sql7eG8R8qoPSewadMsMzAXhFoD9bRp3gVqYck
DY8D1BKWKzB3fVnPxOD23zEaLFlAWscBkro1DYm4amWhOEGa0R2JqotDjR32
SVS/MwNqLzPWfeAXTDIi6RAkfbA9V5C/HYloF1mh9lFMFit5CQENGwcwBc/F
3O0+59jTSodiJCoqWb1VEx+N7/SDls/lcUYQFOHSZ61hQVMjvbgUDvsTYa/4
EXbXRRvRJhLKcD2LBx7UILlUh4jyYka3+0gWuv59A1k8YLMyT0+6H7oNZNle
42rD3T+1Be+RXCixBl+yaRMhq7JZ2VE9aHDNnw+FHxW5y3qiykZmTLsKbs2D
0lNAXkjEoaWsz+2OxMjZmM9/Ol1mRftFCBwdoox+kTZCZ2loTg+qbnBq2gyU
/K7hkT9yY7jFhr0ujfUK2ugMQfdY2wBn5wTh9a/x5I+SzDhWkiyzfUNgKYkO
76vA9+8zxwpuDq/UtqNcGuRJTw2Iw9LMpmFVh7IVy+78PQbpOovkllwyRhRa
bccLMhwQ20yKXWXR7lhBlM8ttOYuzB5mZ7CyBkI9K4eBUMU9UT4paqg7QGw7
DynuC0C2NMDXc0bAU8CqNkPR5d1PzMpHMn4/EBIaz+IgNgx42oTlTTqUpN+P
3cMzzXL7ctjtDiU8bAl3DwApW1QQ2/fhE9DIiTGrG0djtBFDaydI92RGux/p
Sytc4cREcxrYsWfdJjDiLDo1sEgw5YWR2aLC/f0khrPuWsV+YivXoHBVUp2/
zxoXxx3hJoB/V8Xvfc0C+FnsBNlfnrcktL7CV2PefYkuLMtkjyjf2iMpy+u0
SW2G1WDtFC+FSflDIzprcEIEFNq04ke3zMPzyzsZ0ztYYct7mbvsP+tJ3fS5
NKnqs7xpNuMZLddQw1Hm2qigxnmqv2dAXR5d0gq1Ly0cBeGcHCf7RWf1z6Mi
ZZN0Pduj1TQlNnRlAnsQI7CtksGwAvM5bXSoaMQxtQ3Isx8T3zMHITB5DMMB
yJMhbYTEcsHBF9Q8LadgRwfvnKZD3Bf2dDTLAMR1flfvPzxHu5AxMVreYM2a
9gVEsXvLXL0VMEcb4X9JY0noVNPDmlQiQHIL9hcvLSKyJI+SjHjSaTmdPxpW
XnKRJF0r2ytsSK2ZgXlQmm9vapBv1W3aOc6CcE+QGn/2yf7wNRs3YctM+4rz
atuP68Vx3hArI1rpoWiIadHEzKag2XNnTxsAl6REq+gme3jgqv1QWTR6r9XX
d4Bw5A8BrDcz4FdDidiQ5rUsdWUY3hyoTJ3zV8ZFe8H/48UfvC9Uf3cTdasG
2MHoqTfKgmYMaSifQPKtrOYZjR4123quQPQmi80b6crO63obDLAmjlLkszBo
fLZCJENt7WcsugNVQ+mf6ZhcqAfqQR8BIYYOfKho5gJ0dOo0vYDn6kbfXUeM
mBXWlskmSHdX8LZM+0MIkjPpvJdFz4D3ghkdTNC8B5LeB6yKnHz72kCJj2CS
mjjQSvRyFdl6qXVan/a6AWrJGtbLdhja7DQv1gYODyl2URVf+g9B0gsyd1ut
kwKnhaSLEE+Fb90KFDUjy5dCFCrYya4YF/TbQGMkpBQpXmt3os/KIM1ialGX
VQwpo0KmrwIqtK9S3c3HpfouGoldn4H2dpG+rDdcd/SbXEobx4s7zvYmAXnm
v8iHr4ysEzxEx5yjB7nLZHX/xho8enOLDqSpy+nCMbbSW7WzSjO3kih+3u2j
I6ijfDV0G9U0iUSAX3mfEHYLI8tAIcybNBhvMmzX9dKxgBHoHLsOXizjNaeT
mqz7Dfz7Hpcfpv6UM+S0eLNK3yumgXBamvhc78OgeU+1PXLgz6J2/z56coNE
hbv8pbdeT8MGSwk5ATMxoZm1eU76FMQ1oA5BGIwvY9qqzOw1PPpUeoE/jhz+
v0ieWVWlLexiq9UmNi2tIOp4BGbg0oDnFnJVJm+U8WxX4o6NGUjcm87h7Zxh
sUteoGDyOJrnihFiWEIo2dxGK0k8NDEUJP5Sz5R2XzrZFS/WRLonLV1QBUwe
fF/3lM1AJu3INlNCuH6MOBFlY5l9skTFp8XSGXGdjksuQFyOogvY87o5K6Ld
Qr+ICmXCazsJxeeWch0OCP4kWa+ktYrlJh0tpqUZPr17JGvf3Zh4xJ6oDwYL
FSlI/hXggFYVJH3r0MysLX58Y377fKvy6WeD1UtK5azlD2V+pvd7/dRaqQ+C
MPLRFRNW1b6BSFOoPL8zE3p4px6mZeEb0TfN7J8fc73dldHUYGhipNXfSzuY
vqz/CfsJej+Uvn7tgasEOj34yRCKLvuBjNtRmtgzMX79EAldhkz0TJskHKR7
gDt/t26YfTZh5qNFay9Q4bwzZtqGF8OiF3c+1qdUFp2Z4rhQca5vbWl4SKW3
4rnmVbNMVypDBq/yoHrAMZuZpMzVK453R0BuxZ1AkzeIUTC42k48POr7q9Xj
Rsq2m1WuftjSe/+Z41tToHykyJcem1oXrOwtuMCCCWvdrnhgTFafq9ugDbb0
fLJB2A9Jn0+4of1XPcpEoDt1OJPBRnwC1Qq+Yv4Igo8YEzHPmuIQ+2iazpde
ZGjHaa1z9dlyKawldBVrT8OgbZiu/KScyZ3MdGoqGAOywCvFP9cnM8L6vhFX
4zuNpgV7uC+Tr1zVco7C+NDcyhUNQt/mRcjwB5Z7/dbof47xVYcQeZbaXgGK
6DSmq1cuaAuO0xQsQNACdp4pOOoxyRujWUlVDQhMUwtY8EKyh5FjWB7KY6qP
GbkIG2gf0ubNk2H5YCblS86CFHrWawz23G/LNRTOaPQzj/0fWzS+GZUDSK6R
uxfR9SL3EIbXS7T3YMMIkDFMgKOdtj/A7E7YhprgMhuB+nIQoT0aFSzQZv09
8kvNYJP+GkIaF5NBj5IITqKyznlMr8VS0/gmFGymvGpfVz/syfFhpv13y4ta
SRRZA7YFfy+Am8pPUBSDfRvyi4OdiiHavhRkDCFmzmEdH8lb9Qs50LQXKYYo
EK1AAwY/5EDs+IaKJnN3uqhvdJC5DwrtD3+f6xPDB3GQBGD4ozGaQEfRiKx4
1F3NMdKcL/7SHBZqnOd8OzYxTmRMb+MJJXGCyVHQBEYbz23pwn64SzLlGkYA
odrbxl7S6pR6U/4RYp84J1cRa2FJttCrSU4OESOXiSkChQ28X7k2AAhxuwox
Rx3mqzcbiA1yhtCo9as+wFvmPoa6k3JsYbRGcwt8sqlP77pOS/+pdE2BjpAl
TwPYoVGoH10dBeEWVgoyT0Z5KTzU7XZs65k7IPG4lV14DWgcJbcD41XQptoI
owBUbeRXXX1Z7VzVDCOCCYO0IOzbr/TIj8IPumgsBuusd7NF8wtQ9UwqOevy
LkM+xGSFSZbgcsxp3/VcXQmg7TqVLUthAub1233gPe3I1hnY9Xv5/dxdEHeX
T1YwteA2GVe+X7/43Yxb+VFfIsq6blre67WHs2+Qf6w1YKyEjUVE6uxiu0dV
BTQeM8LGeLQPlCXFycCV7zPQyJczRb8COde4XOWbAejIOTwNN4Gt8pQNfg0Z
IpFNYRr1/MLi4d/ZWdW3rOQA+wcmat48Fc6uy00KekK65QYnjffTaQlqKL92
PLJ4zViR7wDwagGCqz/BGke+jU9mq481uPgLFGBIbRcESCS3AoECsh6JNB9z
brv++PR7nwE4euEVuGSEOD7XZFrvL20uPIaVgsOEwd7PLLpc2o4bg4EY0pvi
gaPKRpqfp3FfTF0BPVr83i3v6F5hP3e5dqbSmET+mllmS9OMjClpORzwGDeJ
djyX/lZL4hR8SSvUvuGbxCa6Myo4wApRpiw85OopnjKCpG3Y+2RKEhBZ9+tY
vD/0qC+n/ua+eetg+Sv73gEs3URXu28gUy6J14LZ5NfC0ys5HhvBFNGBoO7U
tBUyVA/BleNSeHkFkkxGXtjp01fEpNLKLR+3YwegAcQ8fIhXSdD3dRIlZy3j
2R0gva+QmvaUjuraLgz20AA6hxQNGAckGshEPWPzrVNjACD6V14BSCPSxjk0
ilLCK73fy6r/hixhImZwXLGNPJ743hDwOd22LbfemdcycAEXhBLToCcbDPtU
50+jBVTlsAxt/OuVb7L8KB3NkQnYcbPgHz3bhTIaj08gr8P4w9wS1+NTSRyC
CVQz43wlysOR4/DB/9O8aPYjsqsWzQi/y7ZxaiOAGNtlad54fMFvPBrvb6NF
LwDJs357c204BvGKhI5FERoV7wAY3GsFYW1HWVes6abVDSrT5vzAw/iCNnno
9toNU5VDO7ppCHguWtyt5wU7pdHSMVnZpnUYJ6mTfd/ZVoVXTrZlSzEU2J40
kmOgoejeAVZt47qeUWhZoCcnsui/lEXTiwI1QfYli9ZDYWp0oUk6rOOeI73w
TZvJxMNQsNkOpJKnBI8iewxP+eakL3+m0fiRAM77Vda7DBHKskpmaUJrGNyN
vtUaWi+kY2OvtDnbYfIQQYW9oSNfhXAGgvix8uynXViPrEYERtk2PdZeeGD7
aBMCZ+aXWnTqvkUbjL0yITir+5zmP5ExOBSJrQtbxg5Uo4qpvPXB/IdLnIxq
2pi5wSmYNTFxNDMPlGiyLNJmO1zrX8zJgfZIiVoQggZ6bNAO5f2b6gtD2vED
FPM0V+Q03MMVOGVHBbxdeEPNLzTkfCQwqp3nWfbIIWWjssIh92ZJUQYXgXKE
ZpJR4EK9RkBTgo/T9aw4rXlry9PhIObAQlwfnGfMMBThw712Qj/2lX1b6E0l
8RCvCg4+h/cU6jiJlod3rOEvkSHrMqDjPpgy0lUC6OGhmEUtW5t67HN7AnAJ
w2YyMLBANhirI/xBr/9cV6oWVD1dmjH1rgm6YhCjCtR8uZp13xykCgw1Iprg
8Km8XlhsVoBweXSJccjsvex0Hsg6DNO8Dgnj/cf17O70wfCs9IeDDyTHmaW0
IjVJgONr67858INyew5jvCvIaEFEwTxnwfzeaStA/oYBJvBI+F++fGFPgJs2
j8qq6EuJoNMLjtzy8kywX/Jzdvy+WqcT7bj3RvjWmhgha0ZRh4O1XuigtU7V
34eQoTCbq/InNXObc+AoHcNgAOUHD9Ys6FU1VzZqRX0nPeVkNd8laIvkF9Te
z19vAZ2zQ1haxD0KKhBoS2NIgZtfDJgP2ZbctHwnln47Jbf3M8M6GhWMkH7f
8ZSBv6cJnfbKCDVbVaDpGHTAQ9TqFGN6u3z2YLq+EXvq71n5J9tODFU8ayda
B4dFFf1Km+SMNjzp7arKc6cO3OAVuWnX2TdCqNuiNbB5ri/7UnZ1J8LYNMJY
l6WO5yS9qd4YGy1haI4RpDL4brece3EKDhY536wgB88GFmvh3o6Qgkmzh8/v
ib25Zb4knzXVxwOHOBjQ8Ck13gwTW+pPShjhqTpgFoZ6yzCQeTvvH6hcNO3U
lShqiyKB+mKl34OzNk4/0Xo0ovRgWhbvRPD6AYySPUiN+DrvQqvg6on/UruX
elJUooxyvxemgcuqF3bLUmyF5mpkrizBBOIZyWKo6ne6VLpfoYWB6GgFbZiF
z10CDBIHZqJKka7OtJeN5X0muTGgRI4iupGGTwUxOijs/mETXupqIO/Va7Tr
sycAD2aJ6M7o59AFakvjfVLfiXvsHDQgpJx36jTVpOla4qA7KbDx/Ou/r5Y3
Llyi5c9C9mBGbV7pFxt9YQxyjA1eazcIdFWgMGwYiWpYaKSNpSTiZQb80o8E
7PSIJVkZflO6WaBv5Uhh0WRzQeI5AFSkGzxaC9aVUyDyZXpuH3ThMYucouJf
j9Lt+3zuoUjMIDFnGCWMfKgQWdVolytb6SNckkU+gfbwPqvmODiiI5SLh2AD
1K7MdhwoOd3UVaaEqaIrDpWlZz4Hwglr3efYRcjozGnfYmGkHU6os8GXT7zX
08K/ZtH1dYX88x8ikerFkZc6LhGAl5Mv8sH4beHbtD+R2UTvA4v5A3t7/2S0
dRZrlUsrAScPl9WH6v+HDCD/+eGVAiGALhgAv9HLNK8zIHy5uINuBCCbCAZ4
Pf2Gvsqtg6g1s6fMcUfDnqtF77fycjjXxVbexB3DEcnOp+Tmlunio3AAYVc0
fi0m7PCu1EYNiXT9OJKAHi3Jz7OnOOKLlvlk6CsdeZ11I4XZrHbhBC0DPNLQ
ZaHQT3eBBxa9/mgpGO1Iw3e1l8Ar/SvBw92MdJXhTVpLJIAvXJTWGdAOlGah
6ZdfdDzYsH99oqcQTnf+SsuXoxzAnoQSj4dOG/K9t9RW7cdCQd3LMkYfENKN
itbdoXHXDnVgKC79W2gGGl5QuvIyPtiUpdCB2/Pw/46zLTCT/dPbEfkHF2xW
tn2Ugl7hyN2WvpX2vQNaH9vhgNkSvRw1Wxzmc8j+urU70NSMha6PJgcrjPAE
eAjF9AnfWunficaL5ELdLgROqxFVpNM00T6vEoVGOYN6tKC7d+unxay2vUA/
Qv9YiDgtnyrmtq/jEXYbXYwBUYCzs+MM9qj58+TCFrsOu5EVm3wbUttRCmfV
I+5yPmDPCaIO7EcVIKuvqvg9D0zdH85n/G64LxQIVlkeP/EWUXeoDvFzpWRM
KqmnhGejFOZiuuV+YtAkt7OWyHYMOvkNp5KhTSuLuB8Myo2pjC9LZamX0WCv
3RSUSEeuusAE7iUz5UmO8Fc49LOguATQgPo81zy+tVJu/xwpcmRF7XmfuL/p
xiB9W/CnQrCG0jPJI3xbJpjx+2AUoAiUdQTUiq7v9d18WYv099W496vCkGx4
6+OkddxNDXeDqOmXzihWyFWgyvgp57PEBlvcjuLJVNP5ZhYNu1zHjQxUR1Wc
XbaY9vIYu0RrlFDYpkbQo6C+kjynrDRdEtff/KS8A8363Fcn6jNwOO4HHWx/
G/7rppAwlUdFcftbURlez706jibjPQcnTAp5riWojb2pL6m0QhcCZmRJvrbg
txBmDgGBNx67CpY9scsRXmw56GBnv00Eg53SC6DVpxa4PJfB2Oh5ERNBAlOP
1KysBBHyb+vw6FLEgkbP2jQjjrwbaSWASIWphw9lw+ZGDkAQOmdNSGmqbAuO
YR8xaPzVP6iqHpPq1Er8ZX32cKTkUhQFBNgyrTT0ZbdVwhxsAT2PSxsX7N1v
fo4kEgZLa0SMVcW11krQ0sInRMTjuvs7HE3p6DONl0qCGwPp4s4fiPHSFrMX
KlCOaUGDPjZg24XlfwkdqpQiiyPzsGRgZc292URuuHigQB5JW4rUZ6xIeWP0
rDgyDovVTGAirfrF4qoYLRKcUjhvumsYVFHxlpjVmF5HjAOhuMVUuiOSjt+3
Yeujrjeh2IkEsNq5ghtm9aXGRwPJ8+vIqhOYwayU2bEGtvpmSBEuBmEFyMf3
Im0GBBDpsFq5jN8Er/bZDbeqCvyhntCJ+5j3UNoyXhu0arC2NA4kib/v/KM3
Vkq/+3hZIv1FlwS2TiFllopQloBEEIMLk2DoT5pzvNLhG/tKYQVD8RmzzeSD
v8EJ+R5NZC011I0QktHC5W+37T3fbdS6rza6pFf5Kg4NCEl9gYMErNxwS4Xk
FJcFhfZKOSWh5FTJ7OdyOMgp3KBhI0KOcl4icvFyA8k57Y42IK83Db8MpwOO
4SRpZugNYF29LVxqVqrCDm5UlZNpXfCXmXXpN3Tr/Emyqv98IHAQ4wPVg1wk
M28yqI6hTR47r6pj0CnqK7OSRB5mH8nQZwLyDtgZh6M61wgEeDF2PTfTPu90
jGlLiKzezZIaxBcZaIe9nqSGgZR2g/rxx0Y67VSRRmsN44Io8+/BY5ekx79Q
LmclHPeQR8FXjOdiTI5IE4948tF207LN09bGBCXTTm51dlPm3SHNiQEFlslu
OKdePSkNs7ypNeAf+EcVm75IKuR/J0gXfJI0UtEysemsN++LJjUaH3C3MjbO
3iJWz+1dOxMss8hI1/U6c1nh/ozjdxFCK0EFj1UQ54N0Mn1/mW3wQVQJLqxj
svK36L+bmGe9dX+0Iuhy8hkZ2AGLZN1vNljwGP0wiIbRi22zO+nELBgqxFbY
I1RDlCGwLup5unbIJXXRH0ZGXGC/33gu5hU3I0obrKcsS56mHvDEeV0NBjrr
xjEh7jRExKC58b9PuarXe7HDlfhV9nusY+Qhzqq08vgfEW0D301EjK+4aMQw
5WdWeQq6hLV7DrQxnHTB0XI9unDEuD5DePLaJZGkmHQmE2j3mtgFy7vXZ+WY
8sLCTa7fR9z2ja/jQT3TRrm5MlMLNT1SECiNNtezvKNQUJu4K+fIwGRqfYvx
68Dylq++LvAzHTja/mJGphU3I3D8hUc059Q+PwCI4Bm5PFF9eWfl8w/6pyV+
zsQSQJilAJXq3yBemmO8PYwscwn6awUHjHN0/q8qfmw2Sq7FgVu6Bn8tQJzk
uPjCQ5cCIfGz+Kxck8JRTM9xkrSbAUTDWHtG2GjQevabQhbsbZDEvz/gZB7N
L12gjjoN78Su+CfKdXti/3qoBlRrylQ+3zyvGZ0j0/JkYo1WLvgzTvh3cGRr
TXHx8Y9ypi+2sev+cveBYg9JYL/9qHHC8yqMF2WVoHCKiqi0BKXGr1hrP/OG
TYzl60fQHGZYzWOwsM+QNbHJlfRCxFBCstJLxunNjG8Gn4xxR9Jqut0F3DMt
h0gyCUTkmN2rar9+KBNytgkNi7ckYhAcfNhWnXZrGveG+G6mbLVztcf/fcfk
hBV5Gr1OTUKVDzHqkw7HRF9+NJqHE6Js1NJ/zyIIRkZz5Kfhd5vQPc83ojwc
pjc8PFqkxRjGKOZyrxZME5Cnszi4JgdWzm490kuePIr0hfj6zk5zbjEfeMFt
r7eNNxSx+QIicUsi4UAImDvRA6i4TE01IT5kSM9nz95psoH6JUZ+bZVBfnSh
ZMn15BQN5/1Qjq8vg8RqxbYvTcqBt+i2hdAA7YYlNwqV2Rqd11kq/KY2tiBZ
PktCvHAb1VUPHKO3f1+JVu07kpOWnOKX/RF4PghLjoT52EfrD2HscgLksh7o
jDzXH5L63icmxcUhPGwaKUoz+R37uoA1ln4TyssrgoMcpSpPgHer4RSe2tUm
Pf6B9cSI4CZaYgVwfyDejRUpaVhZPgcLr9JSmgdiFTvNKB1/nrf/xAUbCfbM
x8I0aS4jimye8TBSYNTEzAxzkFrUrIXOtXtDoroGhQhkN/9OqaQWN7pL+pqU
yeIpslEyhv6Gxb+HejQgRgcclqpPYOnDZlAf3AMSNdQKXfq9c6ZFmIuXwmGG
MxH4PPPCObO5+1LHPCQWauf6XO0hq/jC3HJrQcyIg+XJ/rs3cZxlSqusAtu9
r7hEwqDqN83zyLO18Sk4tRCYnvn7poKuLxNxSX3wpweEZA8BhbTm2ZYk3EcU
q2lukmHMlyAw3dCw2uvpyaDArq5WI4b405Tz7r2ghdjSW1SmRlPAd1T6w/U1
ef8zsH8wPAvnmqeQgs8BF0KyGvTZe5EWEX0V7lz0gEEhJO8s8M8eosZweOt+
QFHNxFAC3b/MCWdpJTR2KxfXXFC124emOvsbJN85BeKeBK5UmWwYk2EzfIEo
GyNA/eGFa0KdsSJiEBcyBj9N2eMKl9cr2RvxVFOijmoWcUmhpJmRGN7oOGjx
oGAJhsHpz3+QnXJvEHslouswoeAQvyLr1HSeZu0rYRKqciqB4S00USirOLBr
vtUNxQt3wzK4grm6WB8a7Dk6DqFy12+PHUoujwPciu+d2Amh/fHUC4oaOpue
76ciwsAShpcH6Sjv8yPtFckJGL33y/qJL5VbDU7vkMzIM8RN+zQMush6cnhO
NTNEQ7VoWbcY6qomzYxKgNBcQ4wpKwjfVg0Q4iCRDyMnetnP4jEqDrL0Ik16
IZK7Z8PjzsFZ/bqEbXWpHxHY0GaRTWkhJoheZII0XwF83k+ITJ574FBDd5LZ
rDi0HSBj0DH1TxWp06g6a7c7qu1UE9qMTbd5iPQhYpwQCirazb2lSjT0GExC
1XChgy93CjiGZrwUBBrcoLC0pRqJSQNi+HaLXip8CkvqW7n5be0YUbZXwFGO
18jUFtoCO4cwtkFDPy7g3wO424DC2yOnpFU9Eg1/xbsQFXzLOFF17ox18eEM
rza1QiAJG4Pco4YMD0s/ZpHnBdQ36rXikJwidKPs9ZkKvC6yhSOad0YGkrjj
GhP13MMga/qsvh5WrPQNLOgRiITaQ2gZC297VT/wEK/996FjSbpQMeuKagYM
qIH2h6p38YuuQKMn4jyA3p2DielDr4cImJRQDfnFmVm7r1tbz12tvSJnOz0k
knTpVZVGxaI7MFEm+fcbEuxolQeHBwCpQzJTirVK8ofRFV5No1pAJMoPQUjf
aGMdYShGy5NVIg1X7Mc9XWFX7wPIC7yqfcpgG8vF7UKJuWouq2FN0OyKHP90
Zak/0P7C0fuC92AtNwbLxEo5HlzoHdSI7gMjfIBa0BFPL062b+2AiExdrr7b
/NST3wBWdOE+pJPZnc9z5+c9N4ZJ1FnXMvh+9JJmYuzLNrMquLDrOJnp76Sx
J1CCKtHhe0+1lavhaZ9po7LiEahGPRgFJtkECiIHSI0g+Cn8m10qRdghc1hQ
bwvXHuAWUm6WZYdc7HWKvqwQUdoYENk/iTeP8dJVWQfYOEUSRSkgwD42Ow3K
YCe8Gxgh9klENElLzT/F2TPXFXp6Hrx1fgzURJ4S0DgZOHNQcAaYM5J7L2Zm
fB5ztqYDPyNUdET86I84UCdhFrP4siAWkJj14uENmkOTAPipks/oF2B/FiWT
AgppMSNcDhPCN1vFVf36Lfxalr2dhh8feRXtKpWWNsGDb/dgQ4NCKk3gFKMk
HXHBdSeu8js3n7PJYrr7yj4bmQT1aC8vYxKlWc/z2zirbiROMjVJq1BsArex
oC7fk1sb5Wa9UrukXQ0fnU5k31yAijtx83i8fVGeTZw65cLVBn1hUQ65kfQA
gEJtat3JTTVKo2slBp/jTY02MsOGWmiCoIcPOl7V6O0h/CHNo/dTsWyzQRxw
aefp+kv2ZTL+I+yTX3v0ZijhjwAdEZGCx2B5PPDRctpylVsVh9b0i2ttlMIS
6UbBtfvf/QTEjY83zrzMCK3+ER2kOyg+asDQCdJE5PlCNnSkZZITk4pKwmIi
bq2iv5uGSvvUU8Eh/paexozqOdNLOValrxnZG1i3XNixlGAMcOYGbOva1grv
GXJrZPoXXt6NpweNUUkh/H67gSA5i+xUpvsh0XoZbhUXH26VHHv9zhnS3EJ8
UX1ty9JjDIDwczag75fkOKwOeGXfcU0VZHVTPikNBznbNdHnkadM+VupoEaO
1MSGB2k0GJ8/LFHoVrSpbsMu0TgIFJltebIn+xT3vv19stXf7275c7By3Bb4
QvFdQFfabd+KCr28VvkuvSrdPx2NjRv3+tNbJ+W9hVqXNyBLXk4KTkXq+73N
p2zoPoJp+zx/xgas4emZxH4YHrnShySbpXRsV6/0MpVlKzVO6ijHXaMw9tTt
pycp9tFmB2gg+F+QJ40q4G70wHcIj04c3qncaB1dmBRMA57CZgUOxdLNBRiG
0KBpykNFvvhStX//K08h0X0r2E9Yp4bWmN5lq5fovkNF2bx82RorZ2/tOp49
HhxyR6+7YRRgsR7qlXViPaLmVjBsxWw9dEPGxVT+rdrcpl+JRHAi193QVg/U
l1m7xnuOdBnHr1Lij1XG1vtno+64c14wUGnwJEpmgVI+LwqP7FGicKcda5dr
anODpNeNFjUmL5dV02yBH5DV/mpn3KkQ9ZDvrzWuXMLAhxgYU3xcnt3sd67k
atx5zwSY/zGyMz89MaNaJh0qkohb2JNHxDDIgCIvkA+USPUFk9exgSMX21Fl
e8dgiDYAr3qZkd0EHSNvgw1LOVmmFTjCxlNqjLrWpTwakgtHxpS2L1Lwq2QU
3V6q3MSqYbSzojRfUv8H2AfX6LhE7JEUjkIh5Fy1TOhOWul7yptBKRerq1Q2
LXp34Gn2dJ0Wc8hP+Rofg7+3uzCYwJDUj5f/4nvbV/r9ZfGu52QSscFL7s4Q
BdclUZ/EbNZlTGw5AMVPIcEyzcJvrA8hUlPYYFebti37/DZcVoctXvRK8NVH
KVzKQt+uwX5seRz2qZPJITDo5QKZ8PyynqXxpmMfRyYJBVEsGy5gFaYFjYSH
gk3tisPUaw5ypcUJ2V49W9LPqduIradcEjv4/eQEmDF5vbRtCa7Q2mdNAzsk
UjpHspqCtNnpmDzlNYspVCFnUSYNZYBPnZz0ClhuLdy53WVpg1GOv1pHL+L8
zovbZS2gP3DZCAaA+d5mT2mQyxaKB2Zomt7AfXeFuGvyn529dHgn5vE7cSGi
rV8zbu8QuvGyuRfZowI8JqFLahHf1/ieyQp/pt1TKgSBTfvv3xJgPEUo5C7o
JZgVqR07tUZB9qM4jV9JPx+ZZYZ5A+cu0bqZ9W9syb4d/WwQ8N9zEEt5F41o
+j36CyXMA/K1/XL+Xhowm8dPwOqeEEqShyZb+NmGLOS+zPVhIWsWim5LXNw3
0wKIovt3wSq3zZ/4BIsKixlV8xdJDP6owIXeykMZytgKR8ldN/pLtMIaPqc5
tFt6dLaKmhvB/Wc3InaVHMvWcM/A2CGj+q+FbWwPPpODa2mljgWmCGfQPdcw
6K8CAODF+U64s43pQMbu/3XtBrb4YL5gzNBtXqhbZnNC4YhIDEfCfLZ6Uglp
oCDJX0sM+KH7+iBLWErev8FcPmvn6gOClFWtIhYSW6ZZrvtLdXGsppT55OAS
9LTzR+k/1YG3fuH5gXTi7ti2caqjKlbQmw7gObJlAyYKofglvfGsMsSQJG5Y
O1pjZLrufGObT98iAq7xptjVx2j3NiwofUxmrMpfjk8rM9aR/F3ANiIb1iO2
RHrV0qDJHx3jNd9uCy5Ql3TkI+bLvhrsiAFIRs62OK2TmhSrM9O8yMQdtHLs
v6BMfpQdrHyeCyhCx6riI5N23QnUHQtkpcW8K1KCeCKTd+/yshRFtU0G8sFW
gLsh9U2jWrJiNPpKp27fQXZoFTkaqRrUWlOhp/GLAQJA1KFjbM3rl4yoptwz
Wecz1huSOLXrVraWMEuW2RZ5hkAfjgtfC4Xocin5sqgEIvwVVFLICRluqRtj
bHGSbXeILA/ou2KK/WNMO9wz4nwCf9h5xzGvDMg8KD55pqa+T7S08z5XxlVE
uSPICG2iydPwCdbPXmwuuNXC8to2WTo/qfG2LPh5gRLn9Z1O/KpXqDcMtTEW
aGPHML2FW4YNyzMMg1jIngSwo0AciFhbrZKndT8XH42zm61MgMJhl2atTrxk
0TQmuBocMJKzJF8pkitKzGwpujhOS8OaHs34iSzmNeKXTvZessjXra6KgBGi
gsDrtdAw5VtSn0vKzYvZm+/wQ0ngWBzqX82j6Si18RDvEdcSf9pDZRgydhWA
mURYARdpeosUc2dVcl2Y3HKBeAecqauqAN/KsTVb6DHP7s81yw4ivW5u0YnB
R/AK+mN2Earlx3xcOtyuK/qzK2COUsdX1KYT4N9ptV4/R3UBJ7DIje7o/Blf
TAf3TJWNLO0u8Ir2mN+BJZk43m2JZgwuNmBdV6hvnSyfD8/aXnvW0jOAT4S0
ODw1NpnGtoccczO1GU0slDrn5gjIZGDpKZ1KbR0Mrq8GXymNwTexayZNM2o0
7YW6NayHn1DTFF7FvlVwqHaNLkgqyJDASvDmCuLIFoHDihivl+WAQWD3mI8r
ZVerp5kqQCnOzl5Kp0G7tjUvAhgdrBPUBNo3Va4wxCo0KbLu4k/86rJisJu1
si/qVcgU25QXDY0kIP70ctAEl1DXja7QIHPSI1i2MWjOn6RB3orJNCpvWgQs
CVdEowtc4H9naojWiY2K8kTzoPPvQXC0fIi/q4FQkovRfUU2SBML3Rdh9GK1
55uSZ2zmC0Ialx0jdQXRTv9vnXMr2wQK18+T0LGOM6bcq2A17aqLgeC7TG/i
+zAvaBKoLhSymMkH5p6IKGifxrv+JqnY4vtfoJKgV2eL+Q0weV/UOXln6RbN
EmO0d1lCy9Cbbxq1BnxcFJPFKTlQ/UV6EmiPheoIJAmUtzBcAyf55QoOhZNK
M+yazLczoBmaOYKJo/DCgS6wAT6LsZANvT0muPeX1p6KweKSGoj4v7funAM9
tm/ysQGDSaEH1OvMyqqW5g3Pitd4sVr050zOXAcpV3DL6v98lscsM0sqbscT
RMPP0X2jDDpW7mPfS/QYCstW3i5tkJ/46f7KcAPfndkj/3QgTpsGpmYOEDoD
BZ4mEPqQ+eXjxxBRFOXItM7CYV8CHmu1ta86XSdPhMUOBYsoxjWmAcmFMNpk
iXCVEL7Z91OiNW/ge9H9nbbw9Xr9lYIu7EUSbLQnqp0ZLXjyM4qwtOpKfu9P
HNRTGvxAH+HJ0ohDQ1c6nNNzXQw00p2rtDQf1wQk0zbmKV7Bc3l6TozseUkc
T8eguzHKvE67x8Ij6UiyEetvtbxp5jvAaQcgJ4tzJvdwa9Q7B7oF9/46M3Ox
p1kkPpK2GoZoQhwc5jNBm9rKrrGF1TN/H6DbqQ9qKrJFeRHjWizacSruvpQB
B8nljH2xDzxNKFk8j0ljYFDlvzpGuThIfZT2GH5OD9fR+VuLavgesCmpKtQp
fqBiqtEaw0628AZov02o5cD4TYDUU3KLb+pX66X5juA7e+QZbwPhSFCsv8nA
dlJiBWz/WuFJk1V79xV+Y71FmNn5oxnBwmvI3JF1v+nE7ZBhThLDY58zUn5C
XZ09rbYfssg0dQVgTg2Orhmr2G90XDBYIgFP1vkUbC3HIEONTrmA7Q9l7YMv
bspjYD2Q+y9qDzH4O5Fg7EfPThZyjKKgyfyzdtMwWpJkbizRJaLNSwwVUvPk
xFjmKgusGHzM9aGTSEQ36JeFGlK6BFKqJQM9yid1ewI2BF2KxR/jeKxEBXD2
f+NcN+dh9S8hFw13Gt4EfVE4XMFTmKdicsPpSPfGXuMasA30H/s9W5RhVac5
vxVjjldx17hhlk586k4Ff1DIYi+UMEgZR/elHXj+bQZZsRBnUJYIW2oCWnPv
7giHIz7GTzFEleud2PEvAd7WsTL+IU3ySXMKR+Qd4gcWHod3Cb2D7YXirR1x
ajX8SEMP4NcBjMH1qO36iFg0k8zrKnA8H1KC1tC379auzu6He6YMSvb8aAcX
Lc5e2q0p4Korr92OfdhauYx7qPYRx17xRHsfBr2dPBR6jqTy0ZGondOWRu2N
MtKitxoGpy4sHMUlMTdcmy8QMrDek2tF/SMdvxdATaxjVSRN56IAYqB7X0vn
4hgYrgj05ZygV41viejw7vVPqaxWn9RFdvuZQQAKPxkAhxPTiLbE4/vBMJ/c
X27R72lc6uTMNbEmO376J039y+QRAEocMcbxJPqmyjtlzauoLhmrcWPBh1DO
0QXnnY7q1G5W+KS1k5A4mcxUE+pxiW/UPd7SyETFxVIhu118BiB1ue0Yhxpt
5EN6RicWpex2l3QmloogVDU1YQYajabXYX4/In4o2tWGdI2NrGbdbLGFxNvz
5puLfwQ6J+bHk8oaZub/00nteSdOp9UU+hR4ai/kcHWWBhTEmkLbqTWP5UYR
V8a84e4WYurQut/lmGFis/g/eDZtFsXsMsqpif+rpkIlT97naqjxIgh6F/LW
jhU4E7+4vzTmu2gpyayNGyvViVr9K1cYruA392UKSmdG/eRxD7N8zzmfWho+
bcTh9cCS0/F/EBuXDzCe3b/tJiitbn1bzv7FW2UdZ8sBK0ryh2Vo4YpEFMGR
mm/DKpFxhPSMZXeEuIDM+bXzRgrlH7/umxvn5QteOwhM8pCgQubRyFdjusnT
R9b0SnQvm14EIODINr1tYzh6hyekcHTqjZU7Od6DdkdYN3RYGJINsPogKFBa
now4LXLe4BvHjaQUzX5yWr37GmLa3hkpHffCB3QE5J76wFOgJ4szVm6OUwu6
GnYAOgNKJaCA1r6ANkH8biW2fC2ViZi869RuABq6E9B+JdZ52fgXGXzUujke
P/3v+BFZv2Rd42bLHS75Z858dCuY9wtsmzpxyQp/NpF9JOGjhISFEJPZO6TE
dukuKZc5ALmTKit19aUkAujxWb2KyC6duJp5p3eKLLxxvkfuLbpQAyG5etYk
0bbX/mPYSQJ9fa9p4WOU3d8dzEwoDWuZ0ef/ixJZZCoEbjf7MfjljYCs7pFM
No98zNP5aQ+gCmtqtbc+RTpdB9yM/yny+JxuAYcWhLCNiV4Vcq1dep5kBR+c
NXlo1i4ZENLezXoU2Wl9Wxr3VkhmTKQa/otKsexqtcCc/vGQwvI4tZ7pINRP
stoRLy6u62/blgTwfXfPjTnZQsLYWOPx8E4IijY6VzGswoAaOpPUpvobT89n
cZ47RjV4fwFa7yiS7dJtto1kYlWlNL60SSbw/G/U2vfJUdoeWOUBet0n2ine
ysbK3nyUhksOEnBhldkyWUb0fq4sAnOhAPkIN59mt7OM5/9URsWn/PcJflEV
/GsBQSKyqAqcP9rGHuroCt6qyo6MOSiGIR7smTxWOeU1gBkuMxRCTLUWU++t
D485EUTiB4r1n3oCdZNEl0XQ5/6AHo7fBtrLL+R2F7XLflIoivfsET+qnAxT
BK9GK31W05ebn0sBkTKAel06V4J1jR3oI3Kle7F6l24stE0r1n6/XAtLV+sM
NPCU0i8C2qt/ez1iHEkcUTwI4swunkm1iTnn8NBIgETbiaSw86y9tj+f2Ve+
O8F4fgCMDJ7mcL4g/4iv9WeP2LI8JI6ZlvsW2tUzw+pvltzrh1EDiH4dcl4h
2lHWJV2FH8YQD1evkbWHXSFfdaIfOhrqqcAv6DvzRrxhlyq2khGOlUUeLhub
5ZeMHMOsMy+Y6Ez9pdLvmrar6ZY/c1wP11DA+LugyRw/wF3n880Dpv5fat6B
La3mjSnPIVkYpSjTv+D82lESDLvc1T98/0CcP6GXwu0lKG7vW2a8MPr9X74V
rvmBjd3NeCO1ur0mDmPQ7TFun5ZbmTHE7I7b8FhjEJe4DE9oWidJ25RsS2rc
btkPikLFwCsHV1Ng9wb4yrDH5bhsCKwHwoD/AjGf1lGqZTfHkOVPjqmCRlrY
hcR+MGq4l4AoCxCdLzVs4R8Ajav8xv+YglWuTG3jRwJXJskW4zt+fGSOrr8A
ststEMA7sQ6q7JxUwdcgO8KNNkLNzaaJiZsgWbNhRfbkCTS6Y7jj6npnyseg
xw98pgz8W/BksVMTmMOlJbvBQXM4MceCDZkaDuRem76Rw3hT573hciPC/1gQ
71lppoWbRw+V7pR5Cs23HVsRCRs7U1LHUD8zr87HoKuFLgsWN+bX3zCFvFJQ
dv+OdgPLkMH8HAeVFlB1XRVsv6NyG2koTCEavbqTzmyGjAhcwkWQYvMq59JT
lodAX/bguw/UbhG0LhlgOJgfitJFABNmmvHIFKBO6gP1qvwGRt0MnsntPUCc
N27iitne65E4p5XgMghOzg0QHKW5nr9vJmIzWrle6Q2Gx0Oj3lmfb2oW3GV3
UFCha93ky40JRgBJ3Z9Vivqagh6i/+LEg7LzVC+2Sd+/liKz6OVMLp9jIOdQ
z2YL/5580EZ0Me1Zi+yVmm1/ekSANYKjv+nXDGt+ciVwOJodH3i4whNDWKqn
16jNvdTzviy17UXY+KE5NEFyzfBjsLRKtotbX3WBoSFlDXY9TeyeU+Qw/lOD
wIQgoCTagGy51FPzlU1Y2Hou5W57RL5lb7ZCqRjdnxHyz0q32w11uB5gTbqe
0f8EC5XGJmBB6RHAFCZaVXsVTK3eTMr3pXbZibMN0LWPG/rASsWBWHc77FCH
WhcvsvSQtHNB7o04NMIvwHNkSotGpv+R5EuSa2c4Sr5JzM/uZUXoV2cTMNCe
Sdqbb5RTTpO8aG5hc3XmuUPk14af47eCuKgyaBnb8YRMpr+V2D9V7VPRtVaD
zfAZBsssD3sgEg9n8hJjJoEFmZ6emrIKpjaHukZaVB8nysL3GXfHP3BkNtEd
zQEyK4Zw2uvFRB6EKCmFDMyHSojBRV7HevLyBXYuN++OTA+LUqpcQjii+7tm
8ilNQboA0JebWaEZG0OyLlD3sgVewNp7WdnWkG7j3VM2R5RAe1KtvHtCxORN
7lvMMjHQe3CPrDMIIWx9H7aWT3t+qw+9UcIg0Ux7h3IIsGRT22HtBoN+vSWd
+WphsOu8R6ypOGS3olB9eUbi+XHLE4RUJzyZ/jFhK7Ptq4AukitEdH08obSt
qYUB6s9fOk4TVstEG+is3M/tnHu69XYIpVD4i9uqCk5sy1Q7GgUSr+NB0D42
rLJ4THUA5AAWD0RJdZWNgW/UA/DM+8Woh6SwypIdXOigxemOHEYVS0lDajQW
1OgZeod3ai0oOWZ2O8jOp7SXhTxOeIAUKKM77nTWvrMC6AnN/SHtyEKS5T0S
5btrrJRVh0QPy0cn7AtpbZqwXjkfRNIncylOHv9Hwfy4fLmmFFoxtDd99jZT
oYR6w79hHxJWHycBc48g2mddSJOhZGhgXMhOrmsGGJjaBr3xpHbt93nPM5dh
aZ7FC3y5m4XGb5RVeVAbLcimovVWY4kLV2KzIuLSpB0qsmiK6HgTPPSyuyZX
o973/+Df6N+vc0jWaVx33FyT9A4N2+kkhpTcJ90ReRZ0pMm5zuUg/ZKsvk4I
DccwYCp3tSix8cXMd5ATcOctHbH2XML0AVmrx+IM3Owu7tee1++2PQwqblxn
QNikHthtccONVoApLfQ5k8xSFirV57gOnAHJ3ae6sKBYTB+yyuHF1ci51YgR
ZIDFRHk6p5wcT2TNq+UkIgXITrmjIU4pr5ufYKoG3QmRAoe0BWOB+1xzZJqr
OVmT1kYMTuKsWqqsUpCDNbLg7beEfGCIKVnDKliVIcysp4UytSRYLQ7AnTJ3
FuQKftle1otvpAdsCfc4WKNtxW+54sgqMNaI0d21GfdXDAItHcRd/HvYgh8v
yGyQt3CtY6Y4B9Rah6JqsE4Qba1zutB5iUCip6bTH/n7MdC4C9/KcdB57uE8
YnYYAANZeYlx5Ts+8ROsBtPnGQSe9FMsdIKqlcqIx/eeBuDnhF3g2QLVSLM5
o1KcHGq9sD6CbweI+3Y9VkY8Zzc0haTZJJHnYZiii02XXFu9r/8WpFb8mf5S
Uhu19UYE1BGX0KNIqtRR1UuRHZtydNxiXf00JrtGkuLLE+n67GM4F4sJErjB
+SgQJQ4AGfFO5DB4f/H2rD7R+5qFb0wuKGIrAImvw7MUyNCp/jMxMAGpHU0v
lx3EPQlo61Fue8m+W8MgCjzfBsy0/AlP1UhrOfu9dnXa6yAeO+zkT/XDnRqb
IZMhvWjK7AND4+sRMbetr/vvT1AiK4+Ld2KaqPeywx5qh6oJyTbGCdZ9GXU/
7JBrdI9HkguAlzXK2bM1jez5WcnEYlCoV9+tfnSmWFKySdAxTNuWCYvFqNu2
DXz07il2DWqUEWexfX0s7/A1lkLImEljb8uvFk2We1IKBAXSCjnyyNwf0Uhq
H5+NVqU6k+7F7brRv5+Mw25cQo4tpGc+sylRueaKDMIdcxnULya8Dmnn+jTH
ZPbB8Nmt3W7oXX2DaU30hTseYfm/ogXopwCJcDOhRu1MDdRYfLV9zq5x7hVL
gdu3G9yGmJwrsBLY6L4DpchMO+lR0Fv8T1xDxD6zDoQgA3Y3wAZXf1c2u1cP
3AhpskG7LdC0gOxaJqSyzmMgxXpU9tO92l0GWu2Q0Z2ed/Kp5W7SGfeAOOtj
ZuU0DuEPj1VHorUd2x/nd0s71aq6mKUWZ2vWVwLf460eHUyUseNWPfiSdcXy
Wym7KKFswXe9IMZegVoR3OYD//nnUdB4f/sRr6rd3eHnMqKQJK2aSItcHw/F
gNMJ9YzCc+Z0NQXcvuwyxEDFe2DlcsSavFVbcGeZ8ZRE+GhXt+u2AxEM/9Cz
b2vJP6r2ntCLzHiOmOSgQrKYfyBkGmQyIrFAgoT/hqXOkpK6v9mYp4214Amr
n6/hA5711Qis1FZWKkPxgsYVXWqdgBsWjUcY3qgBzrBXl5TLsd31EDB1D1Q8
EOYd/syDadVIgTs+rSFWpA3wzjpRNh54X+M6vA5Eo7LalJF3b/eIgZSC078i
LOHp9j5pVDwdWaFGtVuU45+oo9h1AKUkRj1iEnSMJxtGUJtixFJn5I9qQN2R
g46shPqhmHlmYsahKr0MGhhPx9q7U72+EUtFjNlC0Ew6GcPf6SAuu/OPRrRI
QR8NqYhN+Wn6lwP1bPpWULfYv6LZvu/nr54583LWLAtFPWlPjIU4uCmJJei/
Ptim4+4OIHgftT8s3p8P6jWCCe/EUesRS8j2xqTV5HyZitKYiyRqR/+CQMX0
Ni2rM5dZzVPmgVT88cI0lhKgJ7y0f7XEG6Djkv1u0Nbcp870sL0daLkDbQYl
QLG7MadeYcHsFuwnoEEap2QZZ0nX+x/T+SNo40LqkfGAsZfCxI+ctU9pJRts
pBln/eSpCkJtNbjIpj4gmVqNz71LH5Ju/e6kF2TPlgt0Qvpa477Vo07yaoAU
Hzui7NupmCKnsf+R1gW7D955MwUcByFgW20C8FUVoFSk3eXebRA/iALm9Ljw
fkGTkaaCQPIWYtvQqkEAfaYY307tvZ17gw+pyRHL3yLxV8losLmySiqQ35vZ
aQaiB+S6Zsa7fgPmbNJh/UuW8zSj3ZAfLpIah8H8pn9B0Vn+keuLP5vRfldc
xq28pIzgVhqvhvc+3BkqIhGKXb1y6m3bpZGPYFv6w/cZ7ST6XDIhHfrz+pqE
Qo1QGrHDXOoAbSJimBg6OTI3xgJ0ZDLZ3H9QB2cpJirhKjstOl9AF2UtoGM6
ZZ8kQ/alzSTSJf7C7oOjHrYS77nA3Hexu/eZ90zDkYq+vPH5ye9tK27VxOYO
i9JWWg+AFY7j6iEn8bQM4lMppIzxp9nkiGWY3lTEHBQR5tuv/Cs97O0fZ2IR
mi9nhsAun96x00/ofR82H0fEuVNNpfb1WWlMiS80tgx0/PGa/43M2rh8pV8m
RL9SQzC/rr41BA64Belt2cYRs5m7BFGP8UeE13MjRp01DP4l3UMiRHyhae0B
dqLSE+pym1alJbPxuuXBIm74snvTj5/sWu9Y+TTBP7PtFtkbRRn0CK5OK/Kn
pXDqVKhm578rrAF+1rb8dZeihh1Y8NnIcTYF8k2klT0dol+2F2L3WNyIj+Sj
vWPEm6yaZ3gc/VFMskjt0DTPGAspNc/AUsflYX+EsMUxmjkuzRPLRCnF2l97
A5a8qlRpR+BDeZb7CkLqnwme/xjOHVE55xgdio6Hi3e8TVtxX5jGvgwBcojv
vBlhj8hQYjF5uxZvg7GpKoMqOrNB1a+Qzrqnzm36VIYsyeUsQYux+EIav2q0
9hfQ0BZ35+nARnXPDmcI3o2LbKwH1zmOBg/MBchwLU1tjdYOThZNsaWXuXf9
rWJ+4krQp79bIwEUKMLIUbvqcl6Gq63N1uZmTuI6GO+ho4ohJNtFKieqn+Dq
YTQrAnmdRiTv3qlnOOk4o4m5Mb3LwZ8nqaPUmw9BaY29rsRaq2cohb7IYYmN
XH/EfjkL8yZ7smQy0CLQsE7j8oIYowghndl4vH7PvSw+ctpKd0WQzvysuzk7
67TfrfUa5+oYuJR2I34jiPeaPP1cyt1khowTP82o7CcFN3phCwI5XPCNDuH0
W8ciAod0uNeBtn6Dx3nbEpYN8Gjp/4dTQ8jIIR8COwdNIz+k7+Vm0Y0aecm3
y2fqST4ilF18E9qtOTh45KgjTPT3YtQXeXMIWVibkQ3IJxkHtlO97la9cF9A
cC+uX1yeFLJW246KhQ8CHdc8vihOK4iVbX5SZUkdGMg9B/NJxFKbWu8AiagH
7YycZAQ4PnMOqKNq5HDHG8jeuTxJ/lVfqQnopMDTq1YBSBsPOwwktC9tR6dU
x04dfi881vXZ71ADiyqkhMoO0LitFNAX4jQlKmWkjovMR9UnKkOOrDIIlNPw
56snLvoUhS7Dff7A94g+YNeaBm35K2U9eYEL36y5SSoqiDEn4eou1E+ZgK/A
nm/zUvE+SmWYnMgnn7U1sZ2RJQDhlAMvfuUg94CpAiatBOIEFxB34yCzu7ok
CABwe/cwSGAHXJHCcRGS1jCcaadCzF/WJU2ues1xdr4BfGpofIUm+Uu3qPGX
ZWw5v0JDIrz21J5qE3+ltuS29X5Kr/M5fQa29bUGq61C8royed9TJMgNeBmU
fZgILpHK6ZGeNKLC8T+Cwp3/dMbK4GHu/iVk0S8Z8P23m/PGJOW+fVpJHBVr
Y+O8J1/p71u27sSvYX8Coil/Tx6RJryS3BCWI5iYNyGBX+v7dqAmiuGJqLio
TZIn086NYSTrfKQSWzXGQZLGzmeeMJwiq++etCud0aWtXvz+BSvEf7RJdsXc
S1jAXIxUi0ob1UZ0BWSbkZot4gQ9PbMMc8m5E6Rrz4Zn0K/Y7avLFdUFe5SX
7u7BAlssuCyUZaDlDGoy+79y33Lwae7Uf86/iyhK8AcBUNIWgdrGSSnKUkk5
7SrVBaQjKSZHA5ruPSsuBDft0rKHQgn0tBQmvk+vVPO0Fr76kHyKYlxhKlSh
UscadfHgpsDlVKa795ApoaZsw7/nbJvJw0h1s8oTP+sVAEc4s/ZKvIyEj6wH
DGLzEdvXQDm16GxEDt69xnhv/P6MSobA973qZqdwTHO5zlKWIGvl7P2dikZw
kbc7jg8p94ui1X8zRA8dHDl+JLWqWQfrtrZIxeUggYsaj95AXhpjmx0HUh37
cw9b/3GXnAE8v5KJFRyED3s3eUGtPZlO6up/o/HmejBA/RVegUPK2yCdvFBd
ncYgZZTQFkWntD7mw9MW3w/qAjktatWemfpXdLrnBTRPUr/pvznCPJv79ll/
kAK1uL9MolCHu2llr4w2shfQWBYAqzdoBAc+X8yR/1cWGCdnTITU/A7Zv58M
hvJs0J1nW1bRFTENL41VVvFWbDXMx82gonou8jxQwvxjOUvY8xaCZH0A82lK
Ti7DWdFSaHca4wDZxFzTwEl9yMnQ9S03GxPkyNjaCTJk79cGsfqlOwT0zSJ5
sVdgGPb9CbAGqSxrmVyUfX/l7airCfig7koxmgaaE0TghVbdLjtVO+7YSyDw
xU1v1hDkrBc4hyWLO/X+2t+3YAOqEphBCzv1oDAtobXwOXTJlxa0pwQyF56J
mI2deFfYA4n2DO+CLaGoyu3AqjSfGgSBaVuMcX6+rxyOiM1XGVepsBEZVmdn
ta7f6cOvgQaf/Gaf5+k+3B77fJiGuFe9xeYcIMZp8PhS47hrjZb5HNLKA5JI
U62m2zz1Ad7ajFy+k0dhOjfNjgmfohTJHIjPyVppFoXpX2/0DOkmEGAr77ot
83MVWNAjTavjhUmFA7BaBeHNrl63vkIT3m4zU/PKNJnbOFLY0djEG2X+7pNT
WuB9uE6xvrnJ79/65HSHCpDtParXoUTJuVC15c0stQPIM61GqihHgFMyC/Q0
myV2NKj6qX90IyrU0jwXvZQ1AGQgUwNQIc8z3zRP/VwNPeeSmPL5x++h5CQf
jx2lqukR984Ca0zLXPafl533Ncf3ze97EuuOLNR5Y5u2003mymgHclnbAf9V
2EzMVK+6SKP9a3+hE0MoyJrcyRKCFomJsq4Ucl/DMiKBlo5aytNOnrQ/Pha9
2r6jw78a0w42gWSPgBNST9e8A+1PnEOPAuMSqo0XxD//ZuuOjrHs3cmI9SAn
qWL4QU/WmMtKEyCKcSoUt0UYj8pTNz6wnqYhRMzvvBurWGUFP0vthLq4A1od
HBYDCtbpPcSy331qR6Ivzf4u5f4QBl1C/nLXizl/AImeI1XIPS1UsSQ1BtOS
xhfWxRwO6t0086sLvRgRn4Ksyj/viheOe1bCprLLuHFmMU7lZUDE6z3A3nGG
+oJZZ0MCJImf9GvU0n0jARG8ZHEt6szKJO0jC4gIh/GeX40cP2XSrTxzFZWv
qYRN42UDmLUc/GHnkSPaiDQi7Cbn6eCTS5L8tJxzZnw0hB8Na4+gH37859V6
+O/QknaBy2ZORjfwAMic93E+3WZ45A4q5OnYG7dhLPoCegMfsoOcgfrAo6R1
/IhvNpin9tRThEOy9KitD6M2ZebWpqOt1LA2C5YLufj6O4HOfgJ25H2KGb/n
nevzMTG/w5OYtiqcteJ0Ck17sv2mQMvc7F/oayJL6IenFZx9e6KD+7/RwQPl
lflN80LY18JCkx/RW3LFAnsRxR3hgXPDEqgLlHmwHBCBwpRtvfIXFjM0jUvu
EgOd2Mzez6/OoQjjji9Fz+xAIefOKtf6+MrApr4bsM+nMTSXdQz/840VbrqR
+eMNK7Axww7Eo62h4ZXDXH3KBY4QvnrLazzOOwtz/WnXmhoCWpUS077Ir5jE
zOE/u9f/BfHZCsmqDr2WmwJY77TaZP6Lw9HuYvuRayNpEp839pqwRW/7hCDU
bJlWJ7G7UbiTSS2Mlw/VXp+0ww8U+JCSAbUsQtrNEgu9lFUJX0i8horSZ7ep
f01dXXzGKDDmvYpnBhnkSlMtVfANKpxcPmqtuYotCkDaw9kStw+yvI+W4g1K
PNshyscE1SzGyfGtYi6i4DSFhKlS9MfUYPzph2RqdSeqDp5pZnw/98vury6z
gV+0+R3qDA70B+cFzyR6ljBaaX1c/hmXBNNhhDiykpAdVTjT5jjJbD7b/4//
Kmc2ELmBY441EXANlCvpTkogxG3pGh2L0GrWn4EOI0vGa68cnRVaVLCT/14X
cImTBfRI92ioUx/vAZk5ZuETYt8JSqhL7xbHX8lLGIjmhuXTPf6obgR76PAh
Z2NDicmQLa/QX58kFYXejUyXDbGfv7W50slVSpGa72kFOx5tEoouz04XruJc
RmSr0JiR0diLsmU7f1zsUZf4FsaJ2t0H4pSSBNFKAXOIhcl6nH+kIffNW59d
j3UWTrh6W5DgVH0VCddB8APZ9//xaqVgzX+BN77KbU1cxKA6aUaB9Forybzh
Spv1Rq4B72PC84omr5ug1VCMOPrI+Wvz1SwFAixDPsKVoeUx/UH2CXJLeRfP
1y0AOz5xsPr62KDDmkOalIBNc7dcz0AN2TKjB7xWFVwEECzKiTrnd+s2UmVI
mExyCtTczUvstDjpxm9CJ0zW4FElHYaFr48+6FCaewxI6IB3J7aW9GF91MjV
01SINXyKkt9ougzsEcHCLxZNFIjTMu62wUKToV+Lq0KFm4SddacfQYJFhMIa
wCAywjRfuQQUl0IEZWcIvV/WwmLTeRzQoeaf+h8HZ4dmK4I+KCCGRVui1FD4
BcziqeAEKxzsj/qa/sVVlc/+nyi7XZO6iPuh4nlO9S/SAxoqLoENGLyCuqIa
WC3VAQLXGhiFu1uM7WeknBb/sg8vVweP5ERtuF7ulXveQcukuyslmXC42OOD
47qCpeEzVQMJwMavmieFJRLKW5u5rB6CyiAXI9y9hq2rdQtaahgf9QGzrBwz
qTYrGeJZ6K96uaScNbgnP3DEiyOHSF/TrzDkD/Oy2YNIDymHvTLHAqaAuH4Q
lwxr6xX1KM8sU5UVcRLPqCe8YUxaBjTxC/RtTLCmZPmeDQpr2MhlgZ1hC8wo
Tjb5KR3cQRdmxLC0EEAKyoP32G6zzyhd9xluB1HrlAwDg7slDdkjFBcCWG45
LSY6H+vGC39/34edYO4ysf/HnjJ8cRC3nIN7VvAS3N/Z/eG9/k8f3CSFkiwd
dl7lZmE6jB1t2Px5JhNGRX1Ussl490Zw3KB8okf/XbQAwtjLMypV23RNdjo/
dTnuKYSU6wjCaJWmobTEr0DOrpTw8b3E5legGOSXfK5upbCfU2xwuo8/vlWM
opeZp2MXx7rjlD2R8habfB4i4eB5CNUysZntoiN8w7Fj0RkE7NlmaUaZ0V2z
m1SEQY79UjCijIMOp73EJJe7gWLIYCDf+57OpAV9e/qALzlAilIYXWUtg2XU
ab/CWPYXnLDrdBN/ccaRB2MrvTYc2qTclAwBd1Lu35IemU0P5kwGLEauZLGB
FE1P6exRl24CJG5JmYBV2BNj4ZisSXWkaKOxWuLLxc7oeFcWBTQAuqdtDWrj
E2h9sVdU6+poWLdjIdxDihSemXkfPg8erQmiuHTQSgxxbQqAVtpRScD3jn1l
sAjaG1yk/lPbg3G/+JRERRuAxxwYQp5d5MLIH+Io14xxbHQYoMZwJuEYsxuy
h8upF3nql3WwlxE50vnxTmWrT+oVY/I9Ynv+HNeaLJ67e4HbjryBKVlFdVzO
FQP7rYjYr90nRUwnOtRN4en5U8JFTlsTjALnlXW6Mm2FzzVD6J0yiDB74NXY
jtoem/FZ3goBFTTRsKEiDb6PR6LtB3NkAYbGrvb9guKFt4Od/n0GJRPJhZYL
nwB0CbFPW1ibVZ7rG0WJTfBSlB3W/kl002Ey+2V4jC6wI4b0PLZR8EcbCduE
H+pjJnYHEOR22Xm2LCF8Jrrci6bGwI3/e0hrAXqXaT05mklE6QGA+2C+cpV1
/fQCk2W/6jKAuWUUx/yrI+GoDeeXJlWaIs447xU4GBtzgDujn8Xf9YaSjssI
J05fcdMTRHDZjtV7hDqQxa7tp2hZsopOgg0cHC325xtmk5VZKuj8GwYjnwFd
sU0d3If2nuVnw4J98opYpb4eId5vQ6c5BWhilwB+/9D29jhaaBU93Lq3U1m7
BwwVEUAyRMD/sodc8n5VoudArrjScgPtgnRCmYGZdeC0hUJfJCdhDrZW1U/K
mOOyIvzSqbAxiy1icTMyTwM2fd/qy4Rs+e0jtUCJmg6BwBtiJEiXRNf1pvkj
uMnmAAAwvXvRd+WAwAJe9ztDV6tc8NncjRFITX5do1qMB34hLPnobSZUWJk5
aFazRJRCt9tJS1OWtkvoxcOhAxY/zneskS1Cgj37WcIRZJ7ek3Vtz2ztuDyX
IfvIkdVcxmzYvDTjOMmY4Xzbz82NQzCsl4OMJlP5zC/59prWDgXnhSsuqzjy
2SxqBbMc0qF9SLlrmGKNRnVEW286yxzP+4cPz8fIKWuESDSD14rXaZoTVl0H
oFhImuPs+VRcDfb7Tp/UIueCLQ1k/Dbt59ZOr7823o6Y0PXcTLQeTOMOxlGU
gVBnhBZ9vSKMKaEHHWect5PeQzQAJEIq+4AdbMzM98Vx/Irhs82bIuRyCyVU
g8xrptgyo0brECwmX/TVrP/CUNWjSBg3phh/QhGEjv7XXfU4EbPjke/8eXXO
filOBnhDvv+byEJ09Z6zAYz7GhBJmr4sNfRScPJSUKlGUUEkppXExwo9RF9N
1BdKQ4JsdTZiSEezusJtzlh2BJBD7iCIsR7+oiM6Yt8DMDrgwHTGlZL+xgPN
r5LEw7uAVfnwz2CypyywrScKvsF0HFrl4SzQlfSLEEyK1Ci6mYAqly03bTZM
ZSKVMiRYLyme/hvY+Qeu+aeFwyqwOOanmyWTxTQ/LLaU7fjYk/4daDJ0hK/i
gbd46PTlS1RTY1HJ5C1Zo68Bm4cJVJmZx6hoUJoPVin9TGzwqXBaVSvdPblw
37koRe4v11H79rLd7OyQ9TAuCdJP22/YgwITpLV8UIC/LK/lLr5d/y7H8Eje
AKqVcQHHwVqSkkTJed8HDEVqzd+VQNAHUaSjU9g/sDSxpE9vADLUAUmaYQ7g
sVwsRinyj9gC4yvwARyRTD6UnsetVfEOQRjJP8SpY+C+3vbBxwr286cqjq30
lJ6g5Oa/XABNi0MW6SBBy6rA1zz1LA1sWIXEhR/TJC32jWdnVFWF4aoBFefw
IkI+owW2tSE5sMWhduBAfSD2VUvtSLhkUyFh6kOQ+aHTG9HF6jTjzU/drctO
U9JRSOt7w9mHfGIN3cVWpNrkQLMG3HEYXe2s5iBvnm1816x0D2byI74uNQkR
tQk0mNa1cX3tHizvinMZ4o33y+zeg/cxPDNVeQP0YDAp5J1KOLTOyrR79E5u
t99YqfWqtBLzQMa8ZgwiXQ/6MqO/95/gEDVs3r0pDqBNl8oIzClDo9G9Sujm
v8/Npac8x+EjjZ6/l06AHagfVn83RnF6BI32tZBJkwOzZVXQ5gZwrFWiLuRP
4XXU3flJ47JHe7VUOJ4/3jArf7L+/gyxn1YQPEwIDTZmAzACjY0O0l9hDcJe
8VgLQzsEbixuQ7Z0DLUHXShRgMehFbB0e4+io4CSpFFF5bdtfQPPlzl7mDL+
HYS0a0qZ92GFlA7woU5WnBQfLv3/6Vh/sa+pWqykmsNRR/GA3sdrrzcatHfP
DLMwjTxlezRM86EGfwj0R+sYFR4EMDedsJt8l0mILgLTnyD1kNd5/40DHn21
0tFmitRkrOQ07KJ5zAz8beGjjG1tuRT5A/hhu1l7eMQcOecK4gWsO4/uNirC
bmW/Ht27ISfyhQepS5/vFQHqmkTcy5BZgfM7sMlkHYd4IBodbIKXqMmCUHHk
M+W+gOupy2i9FxUd0RUBsKhWL3e/hBpe0Yzkxaji9PvIjgWEJ2SDWz6oNr7Y
gssO7s6Ih2LXl+QlkOgRrLMYpWZ9Zq0u8Bs8E6cI6lO4clglXegFUi532ueX
ZNOLsziv6661N+ddafQeILdp6WEcrTU47RMCj4LzQrpE7u3StnSj8unMuYvF
2UgTEYOW3DFJKuvTTwgLx8giuV0Fklu4k6EzeC5hPeSFIOH11mBE+5XcWxjI
2nKmYoOGue2HT6DugO72yCiQOei1x6eqnNzpufCYYvCbkBlCb8yqFGVIZjrK
QuvUPQTRwheMRz1BFcxLd6euxWRB/9BjI/HRO1cGcwRB0KdK5DEB5cHpShZO
/mOPTwTfdmd3Kpc4GXXxlKbvQFDz8Hfb+sMGXk5zDxLA4pZ1+ybIQXIic5f6
AlJfL6VqkYGN/OXBaK7s20Jz5eraubxF954MQae3D4vt/NJnoGHmBUx9h5nM
HrJSkA7pkEJ9Rg7FM14ZU7vo9M3tEJscyFTSKdtT0oKoCh2oMK0O8LcAH8KC
DQfMzKUwKmGrTt0KlMxAmLFEU1/mQdAaucG6pfx6BT2uwee1u/glHwgkb2LW
JekK8GUtez5x2D9mWzL0nmdqfiHaGOOheIaHnUzHmzQPZF0noTt8tQXZJ1WH
HNdsxwwVz/y6oygqGSkp6kIs5LAH8RTUgESpdefC3D2yILJ8OdSDp0o+0kOX
7dfRHysRH0EmUZs6uOWDUIH8/9RDOfn4FHj3pU5gfQpe5oX4nlL/7weHk6Lj
XgzrNndM6L9N5jeBGIKfip4JfuhdI2PxtPPOrGk8eBKebCbe9iKXIAflmrbX
wOdgrmT8OQPAZ0nG84pNMlOMtviUMUM+GR2YifyJUrUsu/hsJo5clNJkrKWX
pkjn4bldrLPokW0+guRycY9EOlJvpXXUr7AmlMAor4xXsLYNAPtFkSNpby57
EzpLDypZckRswZGj4rN/3oRaimVWu2fGCeTMnlYz52o8yw1cTkuROpV/Y4HK
SeoY3xjG+dbekfse4xjUlce43xUP8cmVaE8uXYuD1rUoxhn/AWoWPmWw7l9T
F652K3Ns6sQtAim9ervAHC1S/hyANDKO5sD4xgt26kcCPQa7xvMzVBD+OInp
dEM8XhceLo5FMHWsydXxXfaWAgirJp9hemABXkeMdOOJL2RkvF7K4Z+oQcyX
gu9zN+QKhgiEZkZOlamqwVw+McHtWNiymdHdti5c8L249FFaqYfV/JGPD6TX
2Lshgz6PVnaRdEKIWWeYwjUirLK4vXjz4OEFTqFWoUj9GFS8jLbyNNdElEVE
WWmevHKd1Mj515x/ophwlxR1fEmmJ9dWCUI5bRlxdpgVm9VE4SAWL7js+eeq
0jkXHs1iO5obAerTrZAgjCSLjyBpqbaAkorcalpum1njYy3+UOA6ME7ACkk1
F6JMf4lmgzw7QUmPkkPUxVmkhgZAx4h4r3+9bNv+HyQOgLbOeKp7wozfMBos
UUsfmh//MPaN9r+w3WWr4XU8Vgpfuov1rHDJ6EWMFWo5fYYYwrVIPszJcaKD
VYJcIF8IkObmKCLwZjhwYnxxhBCFnWTQiSaCP/7YetzzEkHOtWHNl9l/+pIZ
qelVpHiqdsFNzu6AfYkozj0FpUGKuf/0VcYsi3DXH+TpSI76MpujbxCJED/2
4v1qAykF0IE7MqA53kwQKDplSD2vzhfD3j0CVjVazGbMcRJQKl0NLEPNxKGc
4/wM+wSVifX/vP6/KZ5Wlg4b9m/U03chCBfdmVFZyKNeyz18/0dZm0hNBLlu
z/OWBbVM5qPF4S9/2/rCV2iD2c14WI09L89cxta3Ul+HqG1yWaN8bh6gzM6L
A9NTh6mH81XL4AzCOWWcWBqGCJhK8rVCESBB8bBmr4MfHxoNg2QmnYaEDAF7
ME7vS9Zoh4rXspSDI4poK4kReD3I2ZfF5kfeW40xZaidgAPbktVU6gYk7w1+
YIeFgd2qJHJhruuTZZ2E4+VeppFYmQKuwt0hSGjcRlnbAJEBLnuMd72LyBz9
aE/36ff0dUv0k7B/b/cemNrR4Uxovh9kDQSMzZePo9Nr5IkyMlx2CxrTZvw7
dLMIzig2EW33u3Ikkf+JuzR2Fz0uVModkEohBJmx6wkDMHu3UwuLy67JRaro
5GHTkEyxpknZzudfzQo4S3JV70CZiVXJbauKlhDBfO0R/C0bA06jUevE/tA7
NTwzCwYNRq6X1GyJkDlsLpRtQdCjYbVDcS6spJgOppR3NUkPRJS8w8619FXM
QIBDUhGf6UAv9+faBLreD2Xit6wxGY+0HFwMBiqF1UDspXsA+XpsRib8ssXR
zOmsTTGHf048cHQDcwCvL35aK/vmN5EEhEmg5k1C0SZQ5tqqhlQH6/QN7O8O
YAZBMHWgAfT8cJsag1Ng9YlT/5ansbXEgxqDuIwOPwQHaED5ljm34krc3mRq
sRZ53GzzAURlTF9Xa/+gF2LttbB8SUCnxSZ/rBwIi0aHhNSh2a/WfiO1mZcd
Oif0N4Uh3FSkNwybmfAGv9lOK3iybzCx18dG8OJeWbt4KgcXFfTDnLKMSeI7
vovM2IGdikdEHtaoZCWXUmHlyLYMRt1SFw7x2+lOnCiK/yIRPfupbdp5ruyr
9/E+kdNg/wpUo1wX6GvwYAw0xZjCt9/2vxauCPFWyb2bklttfOVb/12samOo
GQrjF2dGDjeuLDDZHT/kio7zxkzwYhhB3FzAG3sIg1nGbsb3bfxP4ovYz/Dx
oAKOF/3XJkrfnOXv6xy/8H/pnDucYkWzWWSuB9uCcEOLuSEhZff6Z31SNwQ2
rcjbVdLcAz9n0A3CGRz9A+zmXS6x4h6cID+2ZOOiQa42fpjjVE/JY9Hdt+sR
Pmio4xj0C1poJq3EfaoD8MDmrlFKo8guGtUrVpuv4LunjbOLwZ4hmQpjXNYC
7sNV9NlXP07Xa99GTHNVW/7zZUTPU45TfxfZS+jFU0LwCwPB+7gUgBz8eTfw
mB3BEltemxVKK3FirdZSfcSraeV05UBliqjGBzyikNnZCCltFI1xB7V5Kcxx
VyrQeqvqLJYBlvJ2rpH1L/TUWjlhY5gsL7Zy73KOn4W1OSsYnnTvlDJWbjuO
LvS/fgZ0cqCX++MrVB/Sz1zb53Kq+Tt50ZCOZLswNQtpfvzhsTsCBMQBVqjd
/IZ1tmncMQQHAWWjDTqnyL5qp0jtSCoaesSqk1vbbJHsBKL8/XbP0OBuQ4hy
VJlruDML5/LVhnzE4T7l2oW4rZBFFcgtOHCIWr1HdtC9zT/1UA1gXwerU9bk
anG6VNhjlv5Q6pAUyUAl0nQ+x/m+SriZOdVo1qTWFeKHdPU6ta+WeholkwGR
U84XXSt9miF0uXjzqZqFHv6xZmmuIPMLASFwC0adhd15nW/Fv2wiB42meqN7
Kwazej23LIogjHJ+VVNcgCYOfkW2Mg7TfD0SELtOPlJPOPGY4+tkbVugvtMX
kRuhnxDrEnZcqVWfuhUtmMhqkyES3hSukvWawXPsRAM6764xmjUdnxI9La1i
XKBsS/pA9f191qkiU6WPPVUqhRbPICic8om9i0D9komFTeVyuFktJD9WUu6+
TKDHGFeZURyksoWoiIGz3QDQpLLiVuPzolp/+5Z4cYIUtMKw5OBIbtbbZaSa
at5fT7p9fdguECp3WuHe6ahZYw3+VW0hMC8WuHQtAYkPbbSMmQNPNXcbDmrR
KAf86G5q8JF3CDl4Vpz4JgfDj2yfwDpT503o16iQKj60RQc/Mogc4Hre6HxC
/v73vGwwXtYQWuJ2FQ6qSQxYP7trlV6K87oOrrYRNEtqmZNtP/5/oP96BS/A
kvQa6jRrkScsak7Afe1X7ouVAj5LAeOPWL0IdyEaXJiwm2Mb6P7qjMsNKWba
zGyaxYG3U5YPFrAQUcIHgUv4tn/WpKfUDKPgXApc/SG/fKhH0sE4Vu/Z798h
gyuDoUO0+zbrsDRJiD3YSPc2QypK+PKNI71hnk/11Y4NykccCUNA/FECVr1n
gi1FMF31wcWKmMI6LlViSqbSv/xrrDcAKwsbxiJhD+HcZ2yI6rXJs7JiJrO2
QVhzISQG6FqP+VLcxCUS+0WKAXbCmhjORkeXMW/xjAX4Kk68gmE5F7ZOO1Ez
I7GPHHtraBGVEcJaQaoBW1GSY6yh2VMh51K0V6zfO0IXq9Er0Vik+dnfZ/GY
gpEINDJ0Rxvxde/e6eY2NupylTGx/RObvroHvbHLiHFB/CiFtLhWd/eiYZZL
zwwrs1x0vcyAJ5vCEYo0Aes235xexDQkJTlkkMvCJ0sqg43RTR9ug2XYnfHF
NJtwfQcb7u80s17b8NjYuFAjvXqSbcOSBmP0QBi2hhh77dbb4R5iakqxAWAm
SIExVzn0m51DBigtoYhDoDw4D2BM3iB9EjjDzFDv+lv2TqZjbpd31L8UnT5J
vGG/28JhDeCf572s6h4UUDwjEg7EZhY80p664HZlvw19fztRKNTaSrGdFMuR
iUjONTaLo6D6lJUmSQwqidkaR+DCr2SF3dnKynwGke4VuTlWO6wD7vvjfHVP
W5Op9uTj7WbfWI7sNV3bQmYWjR83+dMOjy/26tRHmD3bzKUPNj58PEbxRSVa
8CF+WSiKf0Z789jMX4DFWV20t8OdqYX5WpOoSficNfd2PjOUNhEqgK8PDnGv
aVicBCFRFofhGyJ5bB46nIohTb/vVrE10DbT/5qloRNVwdEgNrE2LuAHRw4v
ljTJA4N2zKkcl6nrdl6AlGbLow7Xxqu/OIW4eVwm7CvgmMnJPeuQYbbYy576
c+OlTHvl06bbJE5j2S3MxrNTWcviUkg93eAuV7Y5Z0sYIQ3zJG/8ubNajIMY
7oTXmSZWsHCPpU8kYmCvZBHZdvZ5owsLKoWzLloLSKLSKFXhRIzZGU59khuI
7LkOTWXwoRtDmsZ/eWNSnW6ZcFz4hZkm6r3mobKYG01JQQB1WHH85XQPXxnF
8DXKcxooEVnXWZW+Qtdy0maz4kUm37jKFRkl83TzudvpG1+TZ4M9agEQ9uyg
HLHvn2Uicccqbad7BgEZa+aJRIC99TatbC/8qU+ImNCyTKO2awhaBEcUikvV
teu1qNLIDC7YD2yKQv4v0EaktKzMawpViEeHacBIN6uMsPcJymlEGCYjHbsk
fJqG8ZBdxD/5tYNv96xj0dXl/lahtes8V9tlZSeMLRAu0w7i9X8dJkATGgYw
Qu1z/AfepHrDXGUcrwPvDJUMjL5a5+/wv9SCYUUxGXtYv5azxv4IAMjF1b4e
mlw1lSAj+06apueZL449SLzgQ0pXwUlEuClzo/2qEriYPVaPkimawfJeqoub
tjpSJJVEt6ynwDbNUAYJVrjDdjJNAkkCWgqpDVWyTvFqVBTz28HHA7DtfU7f
mHV+xmUC3VBDTfN7Tgi+N2efvUtLWhiTtorrF2yQH+bL92BBhx6SJnQTdYo3
AVkYgDJ12Lz5271Ltx5hk7j6PfQiwAtClR0dkRopOwlgjQqGLm8FWRVoB9N/
t204rZUITmixfbX+nOyG7u8IzAqCmi7efgIdqVMmNACp8y0PJ14TGHBg0bl4
U21yytYmnwPz9tvdch2evm2lkdzP0V/K0qIqGYpQkZhKmFQ4I9HhiAD+uxdQ
DOOKay0YyuDeuPtiD/rVZaATdmhzE86FtbY6z68jKOVlhGK7k1/Yj2o4JUn4
uSFSZ8uD2SXFxIFAhyGJLnrGvtpctKjPZxWbV2p7L9qPgNUfzBL3eWccEUW1
GpEsfuRSr81xo8B3ZazN0g4dMt4O/QOF+bz3nani8B0hChRgSO2PjHgX+sgt
TgEVxdcZD2zFzywO3WsynOJQowC2TNvvQ3Cr9Gvw72Fs3A8VXVhUd8fDfiIf
bTB8jQnQKxuHBVn1ROfA02EY2tj2E/Rax4CHTE87ht83aKwFd4rm8nx4Ymvh
sT8I6ZDKayeByBT4OscGWHehwATMUljkZAeSCmXmjwP02xItbTBsLTEbSsNM
l+fkZ9IGGM8P1GaQ3jAxt1aOI9KCk9+hJ2SQF15ioXF3C5ELYJXt1EeumJtG
4BpaJ31tqSLXewHbuZ19A0ZmmtztdXKdeyvQogfaZHT/37bJVCN3UoMXjnQp
BTHhw0opPtF7Hy9OBF9b1OMM2/MsGRuEd2te0GrU75jYsXjCekFiRRqWx0T0
dQAzS7DFXYOh9k6piUGWn5qwy72NAPhkSDjmNjtn+gtQC0aIlZvLgMcEBvk5
VCQJ9vU+S6bd4kZBYyP6SNgL+8j1QXvg38jujZUVkT86lRJBPD1ebxxqLz6P
ZWGrWZwqV8mdC4kSmcXg8WtOl50rVh5zijqu9Ml8XmeelNpjGstkN24qzKGy
isGAOIjLMmBvdyEeOC4/gKsujS8NVhS9i+HdiAP3VCaZ1b6f4LPtdrj6AYSI
YEU+jEdky3gEtqusN2BHNti4inVoL5t0vzWU92zGo8FmbJ4QnH1Lb9gGRR9m
BffNTkp94DCE1n4Bgkc51SvrW4k62jp3e1/HQ/bAHVa1mw778lXcYLugI4Z2
rEMmAOnjIU14SpVplK4vgvAlRLaLX6XUdoKqFlKQCCXKBt78RbtlJMoaUYKY
gTgfR/SPJwfrTHGf1yssWaWUheR5+RbzZSiYDIK77pyEnEU2s1b/qgj+jqvR
Kek9YBFsJvzcb60N07WOSCSDV9tLAIcNZ6G3Ax/Vxq+wjl5PjjLP9cn3TX9m
lxZeqJ58YERiQvU74zW0qSgOroiRGDGx0wR0/9nxyQf+Z7RhgEbJNWrMQfrf
oQqGOQ6Hq9IDZUK6st39Amc4LyMYPCg6H51nnpxKJKTsDqJtxbzM9N1UPUYC
CCRjJoNTcFH7lN2vum11LhI1MfFBSbllG6g8SaCx/LIYd+DC7oHfUegS7PjG
M3rzpfRZ/0geSw9vnNpOcTImCRCpVbTe06WoZvyjBoMkMaXTD9EE29i6VgV1
FoqShRlZ2T/Gd9Hdie7F6T++EhAA1hw4OTQmxFkup9LrLV3KhsYWdsk2gD7h
WZucSvhfSEifmX1MpVjy2xM84eOkdmcXXyUOacX5lK6B25KA3QTBad0+ZIUn
PW2Ier8fs/vE8IrgkmipZXmmVG0UHNst1jpu0jZvavLCz4YqDUDAZ0NPzxZt
a8qyDFMODP/kcVVswZAO0khF8cFyrsOXnTi0rGxreqjpCedQYflJcjN8Gc45
DC3EZCsXogsu5OG/1eFN31isUC8kqiG9F0/D5fM2sjQKV8CLEnxI2U8gCx37
8IaTWpEpMMAyovNpKdmOZbKCqOkFe9+TrFib2Ga1I98snjhH0aZ0GC7WJqv6
kryqxMR94cDZng5FM1s0W1JBD/6bEDEUULQxW8OACLf9P3+ECDEWdPpB0itA
nqjGTbT++avbMqGZKG4GU20+rtCesWIRusrH6QJtFWK5q2soTCN9gkRppTR4
oLelFWx+QzAY5/aU+vMVnPttLuNfoPfG42WtdK7aVQoTy6IxenGXCW7gzreF
ioGXzsCNkVtBzTbcMBvlKPUuZMdGBBj9mppVfTTaikflpqOClmUJoxT/jY3l
xFNhEI0dEl0kekzLy3xpyH2CqnvQMHgS+I5zHvlOoa57Uo6lKqu9VUl7F6Ix
qEmdmZ/fbINPJ1eoMY8HGjqO9Z03Cn+ar8Gry9nk5eB+2fT+M4FhU7WXpnWN
cSy/v2fPue1kPPwE7iB047bP1dVWlygdfXBI2a8Vd3yr6vYNx9FJQNaJ1xuc
BNLQQavM0xp4KIxMgwF0/AACd5GuZ5CLJlIeZyc313znI1YwwRc4uuadtMdM
vZd5nMlrAb/mby+a3HkusmDYKo143TB4BoQwX9rSSL5pnSGvDEkBBNup9W+3
+WXOSUXXt+EEJ5KMKo6EryB6PDQ1TIQu52OFWpmyo725z2wWBenlASMODBV3
mAESCcYF97wAsheWg3s3X/tdq8mNHH7OdqiEAqGrpiG6HSeHmhITvq8j5Uxk
rXFBy6mOBw+wrAPeSY0jzwx5Zl9yW45unBS0Ouhc1y6IcCeEqdRFxCdI0eie
+l2xvprdepdCqOTn6TUy5notv/Ia5mIxD1ZkSJ58keOt6Xi68xIBg5efGED9
nSx7pu0Z07TeHzso+kPkCuipfycW+UIUpSBf9nxloVb5S4xk4aYbjyD4ESj8
DKab2b2jzDdwE6dyJ6apm4HWN/n/QTHpk50gfZ9TuYgS+yvXx/qOu+/yqjmn
YDa9ZQbMglh6JBAYRnKZLRLrid+T8Btw82bOMUIdceQkPUQp3iyKZec1BTwY
/UzZ3LxJJ5oq9ZAhg04uHv36cciTMTIkXPguID8laZ0RImIn0Io575w0h+gZ
1/TpyjTYcYndStpr1Xx5WRQ78TVKkjreO5Y+ioUPK59/l3wIKrYIF/QRfqhQ
m2pzP2zkydGXSrhLGBTwv5LBCZTputZikt+od0CV6L90Bhf6jJNhtBRklfBi
mS1e13qMMlwAV7BS6veoYT771aojXQdaBEE5SYH7vCLwQI2FI44/KiOZsGv1
eFJ1pCGKUXdc+nKaI8sxNXQShZQFpfcE+qN2g5fzgmSdNchy7vKJyo6F0Y7+
mOPvgj6dckUO31jiaQim3gTg25NzXuuG6XaX4lbeTG2HmvRy7JM33YxRMamK
iLqZMrsODVAX5c/eJGmHgGJlaDDcBLnh2c8fnHHi1L0/0uhw1OvNzu4hg2ZU
lirxwqYsOdBLMgixIjkArNReKPyvxOda00W0/cDQfjIeDk49Pal92D18kdzs
+BlCP9oBZFfnC0tkmPS0NhWnuFHT11GYtqS4j9qYX+4iVxA+zGxbylaAuitT
wI8rnZ3CQa/uaY1Q4IHzkABN8EUW35zGlDcfhtvY6o8NDNb4LAce2KqLRhYC
fgYAyEA9wF55nC/kJ9RNHpiYWkZTCjNODYzjKE8QAOlFo9x5q+4PxkQifQoa
T3GIOs5EI8oA6t9DPiIZh9/5aYzEhO+Y4VIKr00ZRPxBX+jpu74WEWAImGPG
yWqw63YZ2AqVlHUAXAqDeijdS6rjzUQ055o/WJUhm8AQXo260/2sViDTNxd6
H0zUgMz7vg5ktUdEF99xkL4TPiv6MIVFcqAInI2MWWHIjKVJ7nVjqxP4lQfF
+SWAs2/vJaSVlaPddgvq6D2gMNb/x8MAqY62ttA3sBM648suCNcX46wzmZPN
zm1gZ2Ezol2IjzuI5lKzvxb+LJStgVyHkWhqOcIcHIXI4Xc3Pxq4au6vQ1GU
DuIUGTrDncgAwSDdZBFV7eStNFvt2OofKDgpu/ICktUPNy3qNI2QYdObIVrj
4bDVqHdBbX151Lq/ZZ568XcI49yIz0JOywejSVkM4/E4bxAuqUaztQeQzDNj
CdxZOYW4KS2io2ljNkMi+ypVL39jD9B0IDHeo2ZsNbVGK/VZSyZ8fUU/gT+H
pilnk0LVHps22OAg0tPWQ8t51iRCK1bIS9ldPk3y40tPzJCcUncllsZ3J9Ld
U6WWcFyNFdEgt9HOB+akv0+IaoCezPNMuCSmMYRg4k8zntIaL/AezGZZjn1A
dszCbWEdnWaa3bj3gr6ezk5GxHDXmDlNifbzHvVi9pfEP2RSnLd+x/9LZeZc
+jQBjNoQFSn8LlkM27cs4+bSDBLP/mR3ZP4PfZZ/fMAj0zRX5A6yQUyb7jWW
IOXuBuqHRVgOo4Kfxil/rUMkcTSfIthxYEKGnn02VgZxbI8mRh3VLQ9zm1Nw
BTuNGZud21hmMrEgAldXZv4Zx6oreAgDHc2jwx1xJMfrU8e/uEsco4frKq5t
xxC55BvQHzFr5klEd+cwtvJB5fl1qjWiA6/WRUjWiBgJ6FHMJP2KczTvsvv2
/Icxj58JCeYoiZRCrdKFlvCpUiz0Z9lIzSJeiwieeuhxNhw0lXM+BSMr5fTJ
shl/k4kC0GO+bMmADLtf6M5gTxz4ks5y+AUzfQQZpn/a99vUfWzAwUkLArVL
oZPjtbrlHc+Vh0aaFf1zjwVihAJgLhuQtaIEWnaLVegw5shL4vJeHnR74XHz
G+blNQhzNfurAYj9JLpNE2vgm60MmIjf5IDMkTZwOpI3TBBriaY50JEdIDWQ
CyNfS8GQP3p4+RAoyshtiqyLbdiwuidtVcZh8sZpPkBC47EZX24A3RSYvCkZ
2fvAVUE06y5NN+DUt4ksy72zDg8YtNiQv4HaJnGGutsRUA8e2zA1FZCDmwMM
V0aJF0u43grBzYkMU4qmGQLGW2XkJ0BGzrYTEG52A9MhwSqtC1m3KsvQjRup
TfXmA+EJrBZHzelI/nLpctuGDDjWNyQ/UqKbIDEu6X+ZIaKGByRpaM+ZsS8R
i+4Tpp6qeKeWGx3i8QUZza/z6rhYMjWfQoTIHx3GmPDOEPpkF2X1WijFyjaz
NNoe6DfqAb7I2pTD33O0HmXBjUXoyuy0kE5aEg7mZI8rrlUB1QddK8pL2fe7
rY0efC1HI03pybgsUqEuGRHHpbyW0AU3YJ/an6Fm5ydDq0qTQqkPI+J9ws5w
kQJvf8MrqPePpV1m3yYUsq0kl0skRvFqOzJd/f7x4JE6mBBJblqPjXjFKIBp
ewwS5d4GkBZOn93oekWqRaIfdMEhWtKRnLVhSGJNFpiUZ9fm+jbbBCVoFxU4
Z5R9a8Ygf15xr0ZzLNF259VPuuTr32wKxQhhq2S1TC8D72xsZQ50vKT71+c0
uPkw4SngepsOPwSji/h1ias3gZot8Rkw1rXCQ0QkILMTZQoeduPnemiHCFVb
rv97dOX777BD6SZDuTaCTb57Zbstvn95uLH4QZ7PDUiqD5dxSIe5FPEtTDqI
vzUyNj2FGD2dfgba/WGzw9pY1gSvheaekZwJ8yWPdFgvM58YA5FLBVPh80RI
Q3yrESVd7TF8mvUW2GwFgCfrXOcDoBlmyAcMZYW7Z5VmnRh82d3F2MrSlQor
Cd4hMjG/CKhB6QE8E/Zgxay7FZuVyiXF+5vuCTycaKlhT46VW/OSsyuXFHzc
BfEuMPn77cQr8PaSa7csewf8OVtKmqZUdcAf+38EF8ZQPV4e26ASK1BkRXOn
+aKiqb2hvM80Ax349qsPGENC+vWJ9LeYZE00F0Cqio6I58sLPKxdHAPdpciY
ekpYXM/nTdpVp8q+zEqA6lFZqbzCJApJo1tYObs2H0pn1ShEMJyTziyqY8Uv
+NPSy7zKkO7l7oV6g4V1UeluUhItqGEkWILm+F0Tytx32xtxIW0OkUi7x04l
0m6V6VEF6n0n1vT+oKHDHQFkiElsaioRg98RsEXlC0f4E6yj03NA8s5X4whe
Qkq7P0qnmGqGsvetySGES4Cc8+Ltj+YY+10oPP7tHUURQLvmbRwMAr6N65al
gfAWUlXuO6r916AgmJa5lb4SzHeGU8gYu7VPakAWBeynlaWSWlpQoKc1GDP7
6kBw86mi3bZJYx3+iujFw6augvm4eZjl+2YUFn+IDAjW/Z+8vBh9XqX3T7IS
rq/g7KvUrz1v6zo+xhq4VNpXOxB7HFOsu36cp0e16gaKioHhXZmxcv6E2CZ8
ydIPV2CZF24MJluqkgndsDNjgoc7dfQasZMwd+YjHEt1/m/IA6zkWhCFLdjX
z0MqJGvfDbI9U5qGoLDMT59Vqf7AfzsmWx9GURi8x84DcRGSRuuEsXJaym6a
gSwEuLnQNvt9PBmAA+2icV0P5dzLIeD1LNy8gJAmpJ1H4eMvrvkUiqBaoa6z
OjkKJGmgf3x9MtYbUqcety5GV9/zKCkMnfur8lbnwkW1pnFUmBpW2TAqrodr
dvyAZ/1mhFlSTU+mcBZeY0IEXXMAZeeFQnjTBiNco5Mbmz3vlHlbVcPqbytZ
0fKFwlZim8+5XxpkACFABWiqo1wOpmAyfAL6qQLWBqMD3GYg9UkBiF6i332X
9xsXMsli3V0mNuKCz1Rc2S8nnwqSdflzOwNyG9/qCNk1XCfFKQWVNn4AoBUl
5h/jpTYe/b8LOt1kBGaJ2S1kaGJwa4/GLSZdoNzBhbwg0YLG9tL78UNlMXvy
wulm3eYqwCsEOyvmHPwxrd6sNAeX5xSe37lvI+uVQtkRvyFMsHO0RCA/+HYY
PNaAXBuWPVZPsDdOieed2WR9XB2VNOZv53A6BKWwhZtBrGkqkj7VGbWBxE8m
eatFqKUXlwU5nXuxHYhu5iB64tdCjFExY/LlePqDNM625zkD0L41IlyM3tlA
Th8qIRepQKCxCLxY8XlvX1g7PZDzB+DhYRhIxW5bGY/APs/brI8i7hJHVc9O
htdVXAdGzpQexx3NdALYuFUkZYwV0BKCPLEY+cH5/D8a9zumIyJ8BRdpA8Ft
WE0LcfO8Go1Socp1afvuWdgI9d8zfKaXivvvQffu2Y0Dzo/uf0vlFzkVYzSH
PQ8tkHJJ6/+B6eq7RWN1oHD62Of7pTGYwX7372V+GJrNT6dW1YmelV2aPGCS
A2u9gz1fKmW7YZJOx6ZH5sTP7ITX+iPfGNcw+rVW4aiNakWU+urm5vr4tXV6
3HHLJ305jPJ4W5CoMdN5e9Fs9mpSd0zhbg8uYdHfY0xrNfy4yM16QKyZrRRB
E+v7mxJnXAEtKXltESC4v5/9ZXyRFW0GOUisrt/7waF9ZNtdMuNHOwc6FsDG
gJFu0q2Q6oiNOyNdDXEorFMjY3+U2zd9vcXRHokAsJzxufvl9pA12WuIWQwQ
pNIWKBNos86sQ2ff+FmWNqaHVMsnsjezk260hmySitIEm3MpTh3o6Aw/eXDD
fjKGs6U5m+TD4Z4oNSmMYr4X936OEFKNVZpXIPUv1gpuvHKdxjhH10SebsLV
HIy8Qk+5FUo4MGCIiRfMYnLYOnl8DZESFSpVX3399ixF85HGM6Q6S4tVSN++
GPBucrLJDTHGKmyfhfFFQH+x339KqvlS1FmhywH4n3SXQ1ikz2V8ZWyRh/m1
P1hqSQKgSlPFrPk/OLmdRn2EMClOC446aOfjAzZLCSPIvPtyzNKTCgqdZswP
36SwBLK1fAJxJu7Cucg8nzDV9pH68zGK0Iq31M3aHVby8mOSW1j72TmjPWoA
9CilsukA/srQiuorBjWa1Bfm/iVXUeJ0Ujxv5N2K/orZaXo8AeoEjqTJLNq6
zl/atYaA8C42Wyl90cJiUqGtoZwi/Cr0vm5+nmg4a+WHrH4loyOWDTXIUawf
VGTaphYtxPSAD1J6he53ZqIWT4Swq7Eaml4CxqKOCw6yUvl21l5dHLZFnCaQ
xnvPCENvIR+YvixbRXKEfKOmk+2BEma9w32bnY9+8A831MeT+HKl31BTh9ec
7oE1KS+5jFNhONMkJanAavzshf75jWS5fffXPa2ecdAKecIEPN1zPVzJXJkW
oBr8Av68vHJCyKubMKamhh8gG3cSQuMJLi84Iq9/bASdoOSIQoOw2Dd7TSZB
Jr4hYScoMSk+OAx/E68a/aayZufrU0+IL4xEswXsBvSVUoVAlzbWL7s0GONG
cBXd4SH4TZGyQW5F6WMTXg/Ez5jlhwzuQaW27FKKkWrSnOG0/96GiCuubuzj
5/uh/jIULf/3roQP03gVcHvBkfR3UWghfYjllNaOws/CrR/IIdZMqtAo/BL2
bfweD+mtPSo3U13TAW1AELmrzMjkMS+7HE0nTwyxMnAdxUIp68HKE2fDtl16
2uAasJCBR1wSPfPop+LoI/X7qscJ7v+L/Elw+kBuOq/1r/x8eWm+nR2nVCin
zn9fEXcw/y8gUHcs/WGxxffhfpGAZmoBK4stV1e6kxZldYHm7MRZK0lqp3nh
bWFUXWtkrvZdcftW8tag6AFvEGB2VTzifukMMmglZgmwmP+ngu7FF4Nadhl/
QAxQEP1/ko2ON7vNB63kE6PELd5liWmCYEP4b81FRxHCa95FYrFzdzYQ04H/
kU4b6zoSDzUdwQxtPKbe+iyRZMFqqNc7q5bNF4am0IiFvx0RdqSO0HzU0qIi
OfPV4jn271uVn/UqfB2KvItb3Ec4mc/iwGguoWdY+PCc8Ih7cWMO+4cv9eVq
ciYVrpQ88gV15hU73F0iM5DSUF3FMiBzETWtqcidKghMVnqUAe4ZeZ8kvAO1
5syvmDqxlDkYekd2LS18GNsUBirC4regZDv1PEPvIvUpCexZFTlsAifK6fig
PwHI337V91+3tDKEtxZ4eszuczu6GIzZg+mfsAaoiBt2ZQ4slrnQNpuXq15Z
t450VqCnMvUFFBTLSef1XT5GCnCjc7c7vF0ohd6jVGkqc4WZFJ1fg1QNDuej
Rg3ja5+XlJT3zGtn0wZa7SjEZoBpyQ2w+bRMeiMmMJ3gUBYLxQZxdmjQSie+
NV31RyWn+V7YEvcsS9e9u/bgqett9eHjJSPdtWxuSiEbqv/MFruhrN8yyq86
HrLlCiDw8FXWgIytNZf2wGItMN2Vd/0i5ekRIFsUhKlBapbap3BPPfZFesq5
VHSD5iTsn3RI5B48Xuq8/I2NvMPTLoDvLciviguKj+koRp81e65upncr7IWt
llAzbQchudtuYfb4SsgszCw6wYyJPIu/yMgjiEi626AUlHbPl/WHCZoJkFiD
McI1qJ/tmHFJxZsY4A9546DUPWzmXwNrL9i1c8bUKCb7We6OMQpIvkAPIHV6
OJU/eCZSZBAGevOixs6q0n/zUJdfP7K1sb4tZksYhKWbNnvXU7LLd+PAwqeK
3f30OF2lun2HjLky1RrEGQHGoDreYciy5kD3LE0QuInnL2m+QLPQjo9LmgJo
ABbaXzaiv6es4oxm90h1qqSH7CV3apUhfiO1exEpa4P/tlLyB9LvP0IrHpJp
RIlqTC9PtBHF7OKvsPt3cKF3loX/Pi8/R5gDk8bwg3Eou6wI0dTGWHMMsEuG
7KSIJ0zkX7fhas8xcMCsAJodFQVLR2STrOV7OzNmN4ot+7Z1g4KNzwAfly++
VcxZM9rWRcV8EA4vVgLa2tYa+lOxtXnypF5/q93m9eLvzu4qxW6+TJhTUCDR
CJjyTJ0cO09vF3owday6yLArdgj/c0uw/aikCWMo/nRxX0tRolpRHUB1WmEx
carrtj639kSTgmSmNuisNW9G+iRMr+sWcYaoLT3wGbvsWWKQf0GvkoUV5T/A
U+AMoNBkAV3tHneGp2UKkMsbbT0UitIlZejhJtnxfdIyuMo+/+dEsxB8JtX4
Cp+blF1m/3KBCvPDT8clZDT96iD7ugUxDmSRHJxGyn330tSpTZcxzfm0KWTn
7rLK+awcJQvsxTaGhzdPMOlel8QSUpoO/2Ni4WVXYN4eA+FxP+EPHPemk+0Z
nlPwofI6Z8xnSvmgZA0yJt3ASOGs2XSb6rgXtZx80RZ74xjftJJrsiV93Yuy
Wx9T8d2l9VpjB0E54/ks1XIGYR5BWfDsbOMbnDY4EiMgt1eSvgM8dCQgLYkY
dFxJP00vkXRuIDrMfp5Znk+9/7OAUUtplz0W49aRJLOn4pi0dIb2JN+GNHTb
Fv1yqBlOYwQJmU08fKWNbh8LMV1Q2PIPdIhkwESIkctskeCMPBWSLq62kYDz
SyP33CKBFHAQ5xkuQCtCpUGibXZ2m7Xkq0PxN4URYbfA7zTgiG0UDYJoZ/eb
LN1NzIRvDBLdBPV4w5oAl5026NS/7+sdLjAJFgLrdK3lmhsPmX3iSI2YVclA
Rdx7vaxKIINF90IMHqS725EoF9eCppxFiN0QN6q2acYt/PwmsJn5O8aAWoAq
pNiF6m0UmHzJ7Cdrx+snoQ5CPMLWgtRO/c4+vszBWWxVjzACQykXk/6TSqBS
CpEt9HWG5Vfl8YEnKrG7ROGylv3oz3UCgppsVoGvCZyWlAHosClcrJu6XUvg
by+XlB4juikDE3bbOF+XYsJAsxBSROAFBbCRcaSJKlkjGV+UkRBYxWi95Glx
61FXZnfXfNvQ6ChMTCv8cFeUAetqrBMjswBcLQW3y8P61K8DnuGBOMgclUTJ
8B+vN95TVJ38N0LLWEAaukTMvbsMaI8+T0B7aa36lSHAwVY6dCYIVygheCVI
Ctn/dhBdqI6hT8+9WFRnNrgujeKaqV9DE0SFT+UopbNf3CFxnjWM7vF6J5j9
idRxUHH8l1ZGMSOWodgtuc0gU+R8Xly7fW6wFK7AdZlIKsS/yz7VHqUKU6V6
zoqjsy5EpIqIR0IuaApMbMPdX1J/vgEN8cNSv5jFJ/20Ob190fZ0tZ9Dz9Z2
YAQRV/YuuaVTcZwiAnH8nyvDrQb/uA4d7pMN3foXrxTPiuNtEx5nBhCJoGN4
tAxa/jplxOTYSGgVyHbN6GQz+zGH165mkkxWJRrBHrd4q6YCrH0iO1NAChZk
67D3Pexp7iEiCZ+VV2/8CBrZotVRZJGCeYQclvAjHg3fwUAftGTglWBaRcZw
VhjBhT4QQp3hOgvze+guHsd/nPf3pP84tu68pfgMRkal05IrsSOQmNOaFNtZ
w+T46jWvSoukbW1CNGXDEMA4Ecfb8PdnIByflECp8BILgrrSVwq0cgglbcQP
o4FfcFOSdwvWGGAYizmA9tWaFSwGmRdZ8MKEEwgaaEP4O8Ai3LhtTr1CyIeW
pTmA+ekP9EDZtyTQBohaBxL3NM48KobynFMXhNn5bdz4oONpn2seJCC6f3xm
oGWJ3vknXJJ//WGRulRZx/PPU4YC6zn3fLz42AjG3vCA2vICh+p8+57VfV9A
ySPL+FsUJP6X/1w2AgqVAtVLfQJfjKO3/xRxd5XGQUnR0kmbl5RZhdmSu3kE
sVKCoYuHVqwilFUTSBWghCAOcrWUUEd8eWFp21WRxSBDxyXpLJ20f1tnGLa/
u04gJBpxBRiIP71goFMiwK+14FPgfcKvEKw+0qzHClvb7fW643PJsdEN6PtA
7/ILw/edSmXXwu/qIrHmF/bJCc6cY/L74Ian258rgmi1x9tfs/UAfkIsw3Lk
hiZD8KZjgMJjgeqEWNN4ldcGMCeI9R9lCTXhhR7yHk0/ChoNJXZ7PgPOuUSz
x6tSvPJLVs/IRy/7NfxWhaij2H8ZLyYQ2SC25O7x6NvVAtOo6YwrugnjPgCG
N3PB9mrpHWB0MvUoTjUGZvAqTymz5ILwuNsc6ZNiF3vdDQluFmECveDLeQMm
Kopu0nlV6DqkkMjPt7NtWnOL7rC7twIv8NmfbQ9aogMe7yB3gP9iYx5E0/Tq
6T0NM0xaOSxLdROSkrhlCd3YgqCCD3QScB9R3klJQrSzwhZanyqdjr+Ki5cn
ExLxupBv9UPeWHpdMe0PUx9QV7NoOEiem/xW3AXl/T54vsO5eh03yL9ul4qj
+UahCBvFuJcXyisIdV9moknD4lAcakizOjUh1SewY7/gwqXteDJAoDtYzj7d
nKblK3Xb+eIKiFXGdUOdhxMzaNEqK5LYGNJHy3nAXJptt2ZoZrJl+SqF6J7M
mgB5CrzKP7A/j/ZDJdu+0XylSJaXmq7JcQ3giSTAkJhzfD4jQ4gsKD6Ttz20
Q14DqZHlq2IRtW8+zYGKzrFGuD2BwbR2N3tIjjq6F9MpfysUswRsW2RmQWhm
pv6SA/UU6BQAKMF56SMOcnOPK/LygcZovR/vcjER7DhzZ4VaBDsFRJOg2/aj
W6chv0lzydkPo7Eu4Kb431aydbgxc1omDVjJapvhShgw4DI/jsuJOrpiPsFT
nY2uUkENZHbE0YErROSGYZOQdLL9FvEO8gy69CUJ+iDm31tOYkAEZE98mf9N
zQGOEmQrZDB52jhCuPOwZaBskzj0OBBzUu4DhEiixeHSmts5TsJXPN8IJR/y
hZM6dPmw/GfwjswxVZcS3eek4TcE9tMPRNj58D5Guxh8qwa2ZAfQabDyHr/e
lVc+V6lRAn4Azf47hiS4G6ugR2fmV036hVH1S1d0oUeq4xPQo5pkz8IwYsQG
aPP1g5cpQahHECuQK18cMkhlqo8O42DKlIdOIRBjjR4t+iqKfbt7Zei8fbp5
qaXAJeIM67Q0T2L0b2Yj5tvAsHGr6jsaIPPNS2/QjcQvhdlJtuB/UbIzipGO
odYE+pWqNi/s0/hIq9VT1ifKuHaayIqRMSkl6gRdR98mvxGdjPLsI9R4I/y9
S2+YLC6qjJQzjEdkdqTaJtlHLu5XLEjzPVJE1l3/FSqUAPuaM68Ovspg05Q+
IvT18cBNgJPWNexmJh3RhZWeRZfaW65x8R7hjmnJlMkq/XPhDOz9nuK4RP23
6GWtsWrX3vHfhNPz7P1QI8jzmLT5Ben62HUnOw08I62p1d3aqUAU5aANB2X/
i13gWUi4IoT/l3X+ehIAaPmumXN2IKFRNiIglde03vVFNeGiLKbA30P6DdcC
0TgENkhjEXh3+K9cIdu5U5J9rUB+mU3xKe+tzbsw7TYRuLSa5p/S3Wd/NEK6
uqqVB2coDxc2XbcFYsnxLxtwrs6XttDAOIlc89GcomqaGNK7FyT73XLLr087
1k1TD/8hALWBVN0mgInzb+aAPORzV5bD66iRSyi0vEe1des2ViejWV6epCdO
6E0pG+9r1ZiryaEh6VSaiUIZR9X0m3ZvwxHCApdK1G/j80bbQ6EG5l9dylgG
Fj6uaGt9T/s+/DTo22oTRUb6AQZVlz22asy8NSJBTFRusmTxZAOoCCePNbUZ
frsmRNgNQ7sQBn3Gn5gVoZ7wft2jYxPPwg2AjxF5wB8D/8HyceGILrxhtwVj
uFbLpq/FrIFPJcGWzHLe9S+wKbFO2WzOygSQkRyt/RCaL1KvHBcaHLwCBTRd
SavH4mP3kI4eN6EL5rNVgrxjX8b0ZZ9F6XtfJ0KVhf2ThV9YU0I01nuiw2XB
y0VJk2VQdVwrNdIANjpt0+fdNGtkI7netgNdIH32Drx8FJjYFs7UiPSSUeH4
7w0gyqYJ0f7/BQoLWPJ92D1m2m2ztoafHRB20ZVJgqRHFphsNEQ5izBK0MUK
hoS+UoJyugHBO6NO5+POS1gdcB02pYAL+Hk9Kf/lXB8BO2TlsysMg3viLmcx
KwA6GMXMHssvLg6AWUmuRDrq7FVwsxcCnJQsu8aNyOR5OrPWh7YBgdNTJguo
LZQWUXfROV7J63oKqmPCgTWopmc9SuXwLbmr4YiqIq0pSghWkT0A00GX4Siz
3i6S24C9A+9RbXMrs/Rvf34FBorXYFhSWXMAdDLLLQEcK2/BH1fkmNf3fxx0
VAu8+SZ6pvT1991YjFr8RCiJtD9HSJNuyHZTeTMYbNXhDbN83AXcnrjfDBCZ
oQJmSVoe0nr5AUYKvS4p5cU0J0XBkKxODz3Gj0gc73LitXxmaZALsLMZR/Gl
+qzIHZu3jTYGRiayqhykekTib3zKviJCV+0vXS+FXBSB5Wk7Cmf5g3v3jNn7
/ptHS4sXZZs7OE1iFBHgIU7AG3xOL74Ryp56fUlluUxOYu2w5cHGhysxGJxl
1m9vXUlcuH14nCLQReBColZ+8y0RpDFucgZwGOn7EfZMdCIEP0ajnvIW3bGD
1Wlw9AMn2Xwb7aQKm1/MFKwCniFuudyZzi4lEPHWtsLzL+7c+y9QyDK+2Fj6
m/REbLUc/wqjv9fjzR+ZxMTnnhkC79TtAFzAnlgOMARHcm9GCbL7rVCFxWDP
h+YII2h4pzeNdRHW9W+vb6EN0J/zogCEoaRtVeMmWT3k+n3H7eIW+CZXjb8Y
fFZzrIY6fbmB4e5bjIxA3cigRZ8v/vhj2a/FTZz+TZAL7ocqh6/kvc6gXF5x
YYDY4rnvuUA4LNZL0u+3sll9LkAJhIAUP3+sbSEvSuW1Fj/FKcdr/ytRGSh0
9A20rG0mumbGfWeIdwB+KD6pgUD57kQZHvuIQ+sY58l0XQmWaKJdbGuxRKdT
ugmhwyBD8VvDtY0Rp5oQhUy9U7yGJfJta3bgzncB2J78nSOKlsFA+Jzh5JEl
+vi/T0uk2l7KlehK1zs03hxeeEDlXLIrehOUOs/XvwAFxNJdbxQauE9wb/6T
GIN9IqehbvBs0yKwxcFA76SVpyzOYWXQFOdU4GxAKXdKGuQdrCOC6ZmUnXHg
3sujZB3D56wOhU83/+dSMDcCm2Zt4bUAuZ08rzPHtI68PHWEJ5jUGxF5JN6U
i6IJ6LtSuEDRFcQZrz4Vdjk71fl5VFPcFF+TmX5ptSGGgPlRlFhxMfKVaa5g
ZPT7pPBDW3/JNoyd5XxkEBPWbIoYw8B2aQ00vutAoIXp+N1eOw8Id8EOItTP
qW/D5aY6knj9UKHTj+1V2HR+GDXd9muLP96zMDXgChVCJpDSbC5SxlOuZwwS
dY2KcC4U7FKtbpqSDsHa6ne4mRSR8M62ZiIcefOpXHOA5UBXkeGFhZV5/0vj
K6GsBsd8qrDrIIhFJig3o4ccZW/sZoHOnIu2XbXPigXC4dYU0a6MrJF3743L
TQzRVRxYkfN+DuyX9bHGf7eq2dyZlVAVarx1pqDyq4JFfl5RTHMGKq/nZUwI
eDLStBi8TtIQ6ZEcIBST2vmDp77QF/uOxFI0czVzZChTzi9FACpulHXCpufq
uKbMiQ5oZRk6b0kQERvzP8SHwnZ6vTt2S3VuektzCzBKtHWsFJ1/4vkcGNYG
BsGlqy491Hb4IO4GDB22O9sJyry72xm6tkxCWc9vHZeaxRTlsbkfYrwp2ElF
fe7NQYBABBjrM+s6lF5cw7zuqZ+kvVW6xe0JQ4SVeOJVRmiE4QinKYfFPYvG
buqGiQwgl03FsS499NRUg73IEM9pEPD4WTkcDpphfI0p1kO+kgCyk4Lnc7gS
prGe7hFVrpkhVM00NafPxpn/W+kuUTqdslzOKQuijR/hkEPBqxyNCsYaBkVq
6rTYuyS4l72KPK2qj5zTHF2BGC8G6ajULacQe7Y4W8snjx7uM3fC/NHMCo+T
1WJnc7Hr24QkocKIpz1XTjNxt19ysE3dRGGFWfS61O87ptgREfMISGVyrG8l
fhdxxC3wtZlnsaLGNXw1Dqj+jvpQX0ZXECNBYXZkl5HsfLLknPhaLHgscPXK
fYHLUd0a2fMQL+IvxtVP589driKg2+JXGXNsfUaSVBB/2BhOkycdODHWy8nS
mkJw1FO9GtGkXhWtJsnHaruweR6DxUAy+AUtdivr9oM5GDpTDk8HVwOIAS3G
IVfAVOnD/cIQpLLEHjZo7+qpVh0yMKGumHAiBAgZ3gx/dM9bgJQpqB9Wb3ng
QSFid1fePat8nSPsLOUwH3x5q+eCm7OwdafQoSNMF45tHZFh++Ho5ajcsKZ7
VtbU0ttB9zI42f4+p0Yrl8q4UCssY6Uul67BQ5+fpKdE0uWLRRqmmfuF49tq
jtqlLPqwvgoQxQZxEV7Wq57mmEx7db0VEKy+bsw+dcoGW8+PYAbibtIS/32w
V6rsujsvYEWYFCIEoTYrC08XjAknCATBblLZrkiywTBBhnRvTtkOR6inwRvd
OQWLyvUlQ6TV6UcdfVN4gtOYErG2/9dnmUDwJqBAQRirhO8+loUdkWEZq23a
R9ObrHczXDXRZGoyfEXvn+d+QKUC5GGsd84YUtLh9WtO/a/SqVOdn3gXBu4O
4ty46ARmlotZLqoCYoonWY9Cuc5OWDW8eFJBjzhFUGun5TwRj4vxoXri3IKJ
AWgcLcSocTW8yqHeJwO+aI+pQsX6qNKS7v1w2mqoZcJXpEQ6QN72puRibOg5
NQbG/31BarMmwzk9lZPUzo0Onk2pLVMGW2kXgHuss/5aUw368zycGPxoqdHG
3/+ndZmCTg6WDhN3Q+eW1XRUq8bXkq6L7si56JPP/TeZPMdI3R0S0U0X8BM8
BYouRfcIeGDA3gk7Z0P9GGA86utsefZIzPGN0dWK8aFjPhxWDIe9NEElX+Lm
9iquTB6cQU69pH6xcXr8Pgg/H4P2RT6oMFeD1N6VK/dXtD/eUkDk85+GZm88
dF/7B1OqnWF3GnbfduiVtF/KRE8Ms+Fa6vqLIYaCoowwl7SynlFmv6Aw2wQ6
1+Wi7qbLmJycGTOQ1slobmkRZRbfPforUAMhiIBBxZDRQ59Uqbmv1o43+DZs
cMl2X7f/w+ZXv/jLGEiySigjhoYoLQ9W4nX05IN9xMuAsZye8CKIgYxH1dLN
qDUqiCn1KsIkDqYbGliTzdjSNy6LJBTm8S1jUAU9JkZt9MPg+cgVMKIOGstl
8apG4tAqgHD7E0ZFncltls2EVi7ovBbfqnVnBftRvsRDoOWs0Hm6oVivNAEM
V8Kl/Ao44dQKZtO31g5W45PWq2bK9ZKG0EFBqR7ZPtozhw5Pg4ivJ07aE6iE
w1npRLOWyFIjYKG7BtthPv3KQpbcTC9Ap2+g/ik5zuBRnOSCR8fpSPivv9px
TTm03xyM/GaoBbJPXiD51PFf5dG5wcXBH9J+ts+OiLCoUzU6TsU71dq3DIfe
pKGeBBBYDG2s9Kx4FHmoLZgLTywBNJmbYK+tF6XVQpojmWxyy9XBR3vthHox
Oixyp6qYw3XiF7L0LKaBve4LXxBx8Gi9+WETtYGf5aXjYTuE2JHO/otnY/MU
szP+C9dUJDj/X/PAFa7ewFv8gWM1D3tukeBSfwFAJJtyF2HKvOeOrwoQgYlR
xvEYqrcabYc571cGQymb0Tkfk9kcXNU5ach8ZaP2aO6LDi0PzJ3W6gQ/pGz9
mDgzjWIk1i8Bc4czSVF9cQae4CnF9DtyiPOKhARTPzFDuZ74kRNrPLnfzNCU
rMn8vyn0ncJUu8yzteQgFaD+oPOGoottK34YTvQN/F+oNBzRaRwK1Qy7SnOb
EqvVnS4AbpSjuxOi95r3rTcWJt0Lf5hiNxI7uTxi8Lj38EItHtxbxvZF0aAs
O8qVqZzDtQMAoLgFU87Wyls9qzcNwX794pUv7aljPhb7Y0RpU7cFOwueLTLn
8aT8Rxcr9uBoaT6R+3+vEegXrZ2BP2fJFjqVbGDCOP3PTcTSPnInqU3u/Bm6
gT71V31dmGZUprUxZxEwPdw9Ltw25xe8/0ivykWDY7yTUDxrxNbExYQb8ic7
EYfDtvaI/7NoehQKo6zqHXMLWrMnJQ9WzoxSzRPwRUt2OREY1Hfb03AQwBwK
gfmgyhgJT0mVdVq1caoBO5B2zTZE8t0GEzIWfwKEU90qNOIaugFAhL5djbiO
wfVrZawLTidDzpGuvnkvL7pkNxEr9VQT4Gnf/donM3224i6pNC4dVxqTRipR
hGz88HMNvh6sTw1Q+5sON+PrxTOThHJHFj3TatELL9gsrGERwj4d7w8QDTwW
9Kw5bmRdxSiF1g2wern1Cb9T01heyqNOPfvKkAKmfIN+aCcp50Brj/EJr/7r
NRneJ5ZSbowQketFQbXHZpVoQSvSdyw76MGSPB+UnyMS+GNTnHYt3D/0r/iW
oPEb8mxunY9rcBvdh76MLFnX3auvd+ELhsXQ3VqpqrldgB7q+lPSP15nV5rs
fbIzx75pNIHxulowr558F43kkMk+g+5oey/m9BJmjjUaEsOTrttfZuEKmPGm
BlAMFVUJG5z3jWV9P8jwSV9M3UFibK/qIizGEc0Z8ZCwsw9E7DOFXFhRxnpO
6Xl+tmZaNHgC/qvbL8CmsbqAe4A67dX4bst3NTQ9+3XIprN9/9ZlRGCdLa3t
Hy/ykY9egh4U5GGnRQNHRr1IvnI2ZHFz6BmnP+w5FEUWuj2Aaqlyj16pimwI
ooiqBC1O7l3Zv2eBOOrRC00WzGo74Mfx4datpLGBMZw5osR8fbAnginNTV+h
HXeRC2dNVQbTz+oCb/7HbOzldyij+M8xTDF0AdlFj+5sy3GmAJLXrlpXOJAA
rmIW51MrtMy2tUqjt3gYARPwdMhLJHnJZy7yfzSVrltQEdA88/Xv52j4yLoh
Jq8foC6wYrJmbwPJye/zQfUfDXIITifg0dhti8pugBnFuVvG/V6qpxQkVSve
MoRrgtuy96aMGHSKwMJkBZIDTHZbv2VtBf8PnyJkeF+VULi2y4zGdBvw+v8p
fSuJTS/B3MtPVM+u7naBpKHhQdyLA3j0/jLt4ciXq3xAcfbJbM7DuG6so43j
VXF0LBCBtYCUt5uQ/leK0rzhjIXPHy6ULrm6oUMhjzpcZmK8Busyu5APA6Og
tycTQUs8UnLElRudF8eNTbv4RMzO8Ebvs4oTaf5s9vCpBPqj0bhRb9O5ZDo5
kpDm0csSSe58fsJfywoSAfqFicOXxGDg4YZhSH32eFyaRVFlpbuVOuOK1fg6
OqWAdhYPnuqqLJOg0RZ8VXBB+GKiZdG3LwB30juX/CfolanCbrSwoFvxvWb2
a7X4jvfdn4NFLSJF0E6E5xst5q+6gW9Can3yW0KwipijkJ865MBo3EpulekC
lwJMKl0AMbNUf2RQFUnx7pnlSfGWBd33UQLtG3eBXsWS6aC6uesV0Q/OSfxD
M+RnNsRgwdKikvTTe8HtxbitvgMWF2MGHbP2hoiWbr52UjHooCtZ9S6bxAy/
B3htAcqIwkRKlCOmban+VkNFWQtEzKIRc8VSsu87gTm5tZUWEi3RWGUlY+QU
hicabDGKp3QHnoF0CLQnw4C8N44EwqUp8ScDBqRaFv3ASPX7ce2VKa/XLuRC
5UG3eCH2dwuN2DPpFNkEAFfL4yiqNKFDN9Jc6lr7FaBpvTZsyIC4pyusceZE
MYl0Zr7aCi0oueCcXITpJQPHXPQQporAjBB4GXTmWPhr9P8HXqNLXm0fzeAg
Xg7RqzE87Kq3SZkMyzbdz1U2xnacDG7s3jIqk74mFIPR2YjB3ZbAEnhU8M4H
OTMFgugaCyDiNLvcNLnLKxTN0ZKn86PO+lUsJbYnSpeGrNQjAGYddm76CBmT
bCiV+htTvH7Hnn0sVYBdqBlNT2XlnYaRh14MnVhjeP2zKF7+S90CLyVr+gJ6
UnyS9dKFvai0PpkGSWVntYlWxNjKm+D7b2JKCNIT5jZ9xX4TYmZNLVrZGxzJ
4CrUSuewq4jcXf6iB2ILuMQe+oHyu5IbaayuJ/AImg1YfbVlvKpDreElBJ2d
vdzwsM/mkGLEdXg06ZF/GSP0UZiCcNRuDaerrzx5SKEiqzHL8cV7mbRaI8CS
iTxBv3ZN9d496lcmcNAj9DJ+6tuwwgs0JcL3UmmKv1QhziG/F/DoJtdnRNEX
Ho3h/wiBulQuKDPhnOHVCyJfw2Y1OOyLjuTL0J7LONBLeJ6hctJ7CLNKeEMg
tkFpXqC7VfnMg5HvNbhLKGnRmsaQ+BDZFuxbpeYxeJdLs507JXAuO6PHI4Jd
UGdmDcXPH0k/mqefXRZAB/KNqmPYbbbV+NhoJvCtTXuGszbDptXygD23ShHh
/7SEGj30nSZ1oCwV24wsDUjW7OsB2yTrdRxa9wz8fMxx2qr5LGUSIGyS64Er
Jj1p0giWy9BZO40zNiyN24KbKDcPjxNwi7j0X9p/Emy4ZAMCwa3Lf7S/j8dM
zLdOFIV8JNZNfuvdZznA3cfHXzDYHAhi++gF53bFurCxznLSbVS/xXLdvroy
0A9zV63nhMc8FF61TyYXeNMD0QyE7sB+RcGlMsg7kI3UEKVCGbLT/ELpuKLu
0iAC4K4fgy3lBfAY3tI/v6ejUHdbmjJpLmWl9DVt2cNN5JoT6JSsKLxcRs67
CgBUa6yAOhmm64UvHOs782TYrQe51vLQ9IUN3K+kE0I16D/zlM5F1+ZLLZHh
NWLhhXZlWwoDKYvqg/zgbrK7nEFQI8/3A9Yqy7Z85CyR4LkacbFCu/VGedeL
23B1PHIGy7s3daxksa3O/6EK/odEHz12kyGGT/DXUqGxBXIG+kZFM2eYbWBT
ddhcAQIfl3HpFxNJU6POMztRfswOcXHLArzA5Ah06naPtAunU5yCewO0VQ0q
Rn8Y4aV6oS3HUTSgfqLPdYuNG4hUHUK6yJLODALLwr8j+nFZJ3eGIB44TNN6
wLgU1f0Dt05RNpZ4yLhgsQRYMFOSM+xlziBUnS9fuM2LTFS2vcq46WYmoBFW
LYjX8u/TWHfSFXhbe3/Hlo8YEDX7808NWv/ebITrY5w++73XCCrdxesNfz4w
6qvmIRVKm0thfglsMdi05xMkmMUjYEcxUfz/9q41Q/2J++spz5tcwGwrm/Tt
xUSywQjhz9I5T+GnqhW62Oy2mJMrWcllncfVFbcmofenZ1MA9u4AikhC89Jg
b0SsO08I+KwV025gSE0lRTpD9Fq/BWI0Sdc16gi6afSWRHytMykffcJdnAFG
KDEpI+SEn3C2125C0Vdnc0zPOyfxuPlQprs+hK56wm68MxVxpkAhdFQxsqJ4
PsYq80EV1icP69ixVIgMXwxKB9jg6kvakqtMOjecBuLvaO1qNhEtmgzd/+cs
Nb0FkhprsLBI2SsYge6640ujNu9hfVMiiuJaoHg+6p7M8w9eHCembnlQ+P1x
PajcKcZivNbSXlIZey6trMqmY8fvHN3zEd476HWfLVZ6zZPsT+3uktF+RI2a
iYmrHYy63wvGB4FROG5IQdixeztkxCWWfoc2cwGBb4nFPj2FPVur7xOf4Yzl
hyn19QkfDsW+Wgj1s98ZPt4gaI7Erv3HErBqHUXdyv4OvCJuA06UCkH8vTPU
v0vgkZ/Evp6jHOyBbivHfa4Edm1sNlxmyo5bmzL4AYZ3mchagACIu1BhYcp1
BwxKAVF4Of/xpglDoPG5N+ucMXDDWCvgecjvMS4ryzQGWWYUm+JWuySWsVoI
nGcEoxGG1L7kBZpWMlKQ7+cl3sqlNiixKIOECMXZiy5NwcG2BCHCsSqHhGxE
tU/ayu9cQFzXAUIXR0eykyUTmq83B/V2FS9rMEpQNceX7Hp70hsCJncVt9xk
4mFvtOukOrwyNsw4t4ZGfJRkLUWRNcaujir74pLzCelCHrJmkV+Z3Enp6IYT
6iIF/V+qKJNZxmkgKEQIpL9szPAPqnV7jnGCmjbyhp49yYj0tXF5tRW2tXby
OCuf/zQBhfuKzEYq9muE0RulLtGRnYdBNgS7DRJ86kBL2hPPbnoP50cOxvKJ
/NB+JjaP2cqZy9xXPVWMBnHobIQgEN/6+Oi8vIuXsODO0DB9Gu9jJXi4/OjZ
hy7ofa4/ZzZu2x6EBV05wSYTcJuszhKlAq/0wJtvtQlgvOqY8TjCfhgaeCad
4T1XMd95/m26lIuFgmdKlE2f6Xm3UTmtnN44hk+O960ki8p7e4WO0VB1AI0l
4SB/C0kML1s6cFYsCE7PGVZHHAf4+xEaJ4TI+NcYKdt8WsSwcwvXV9AZKRzW
ESAjAEICQbed6zlhwiEgfbSMWOAFYRpY6+eKh2ssJ9TseTlaZ87Bk492LOPt
hIPSlqj1xMNkM4ml1ygz626UgJxTkcqOmN3NmluQLlK0y7ijIr8J7QrQlZDr
w/ezuZlU/grKjRs7QYIpN7PB/VzwFq8ouqP/UM9PHPCijlxQvdwdVaIOgTLe
SQ7x1AsKEbJ77MwPEC7XJCZDO8mrUA8ezXRrKPKp8y29T01scVmgGna9WTlT
IbHrxe1cjUYs3BMWr3Rq7ZQEvKOUJjjArdxQ0N+m4MTivt8ldo3c+M9ZiXcR
oirKnYOoNwTIsJ7LW2NiVDSP9EKPxsakpittjzYYoxqtUd99WAGCM3Hv2PzW
EaQ5WqO7SOUHS+WV/yp9z5FAuIlDjiDjrYMIsDLpgZNkHLsVvuloB8CoC8xR
W7c/gzHoMgDneB/InDWIQ4hpzK1w3C9QgZYDJ2MjZ8bos+sK2K2zzRgg7pwX
67iwj3xBV9nmZVmVrvZDBay2grZYtTa1VlcEcAGVe4RLYXSM7T1NtIZObXyY
YtiOUyt07Nim4PTEjgGjVJsYipnTIX13IW39SaMAMjd+Y3hBn30cJodo3IAe
ke8hVk6xS8UT0lCwTTbr/tjja9h2t7oSLYnuJgy2Vr9hxNsMj9sTPEMw80qk
pNp0n6o3JjNKjHTtv5xuv9ugC6OXeBvbANzagzb69M5mR2NdFumePZRF6R2F
wwErTzwDt7z6QsoIsLhTzrbpphMoDLcubSHs/mg4W5NKXq1OIIzoq3o3CJTm
cLMbmsMOnQYuEW+nl9VSEqDH/5ZhluqBEw7MozYr384DTAHG27XhmXiCyRKd
jCtDtQsDsL78aHNr1/9rUIsZhH7Fio7ClifGYVr5Uz6TqFZ8z+3vpUXPwIiI
X9i5NRiyTHRhFxoCQfnlXLxyCr0Wd4Zizmv4wDw0IFRCPG0TpcxMOHW5f4zB
GS4/3iEhsk7r5jwcF2qxuw+6EGGpNS9r7wqQG+ML3PKWDCDtJ8UrD+1b/Qyc
nQjNdtdrDi0jJf0SeE2vsMGiw08U89uD+5iYsR/o0X7zpzq/TD8fNTAn4uow
F+p6W1bjRwFMaoIqT04B/vVggmf6pnAPMtiNspWi1FquH4lliOLFgeYnkHb7
6SE6HAlZrv4H/+F46DdF3vv+atd0WcCbrLVSZH8627e0sXYyAX+y2xGpge0F
3/d0QWTx+a+ubS6r0lmtHyHl95AOAmsNl8GO9xHDBhy0pL+9yfsJBPYXCVgs
Ru/gTNYEobwGCkF6JtLJmeu4kVkLOnwxx1yEPyTtVimfFl9CmH9G08EXjuDF
8RseVH5U2LSZR/GbHsqi5yCAyC9ihENClzUKN8AVDCnnyWPu1hksIU9iGnR/
GgOd/e2l/WEybBu9/dp/zSmOLt/Z8mQpKw28nBATQDz+lPsfElBSazRGLZ4g
iFI3Kky4DCYyvlTbnab4sZ6HrCfOXFQHT6ommllaoSQ8HWMfuS3Y6aH0e6GU
9d0nP708Wu+siWQ4yPUAGVHfVvR8Zm6KGE8xOs8z9G8KbSHkc/hKFmLYc91t
RxWMDKPqXf6u6ffnyX1e2Lq5lYtAc+GEGVedeMKRIsuqSKGJZMqqQOWw1suB
rHsBIilpZWNL6904na4MjoiVAOS1lF1c8b09x+GZkqIsW9v/douwFPKKHLGE
VFyfpeY+TaZHOtbJ/NjGAKvKNahtTzN5YE6ZMZAXxml31N9bkw24JjQQl4PR
3oL695AJbmG9Ugm6Bd7uRnh0KAKtk5iHHXOMHlH4VJay1dc/zPDgF2hxjITR
GNbF5yZK1gUigyuBYbghMy4BRlZqMXRDbDgTk34w6btH+AYcnzYFu+LtJBpT
neceQrh2GV8HG3na75TyOamyRTrBhJCKuRV59eHIzviBT9ZkY/txzwB+d7kc
kJeBQVC4G+oAxtgdKmAW6eps8VEuKsgRKpgkQKqFbBblqsdniXPX/8b6oJJ5
CxQ3bO4asC2dpou6ZnF+DhVq5QcnrvrkXG2h4Y4m435lYPf4SJUmFZ8IaP/q
Q/5nwKUsd4Du9I1It+WqMHzp9dv1bfS/6FZgKPaWZ71V5rB2Iz+ToSTPq2a2
jFUg6K3yUwOfG/ObGoTalmpzga3F0HDGDyBqOLQGbD+ugNbdG3cIk1CL22hj
p1AR7nA12JtsSULDrlxmpzZJk2X296OsuibKA/bt0xDHkwdZuiHpvrUdKx0g
Pqd9FFGWEfLCOdP1fme/ps/VD2HMlXfHwSNWfR+om569N85UPPN2jZ22KKtE
Oo4/IO6Z9rrr0VTxbHlQaotVHHcF1Ci/lolkq+oiKouCXU8/4bLk88xr5MLC
k6mN1Uyr1QNdOkMcTJ7brGrh+twACrlDATo0RLGRpTS2VwNyrOv6+BHUHoZg
Jawi+OY0Vw7EOdMqaaPy1MXu3FyJyIT3ETHqqIvlE8/uXGxY5/fZhT7piTfi
ynxiBDVhcGygmJBZlXkUw/NnvQXevIrQjoYCdbSnxV+gZqu8USbdO5GNlQYx
bj63yM7rUfeZR+vlqO26kMHlTBTg2s/i59YceZ5ietC80KP31gGLc/xK2KAO
aeQQs18OTf7fuab6V5BCpm+7s58Gzese86WRX+iHxjZhoSjf3QSHNuMlDOd7
X0LjCfi4zoyMArsQ4GgLe5gSI4A1YUi6gf2lYa+2XUnKfNhqI0v9CCFJS+cu
A2CDEFhngsP0WuPAjvuynntuKaVGCDtddfqYmzo+woV9GPP6qTukaBAcWOhK
jOubTUR4VSG6AbAWB90Z/sCNzHcYaxIBbwXO78XUYDwFHsdVQFfMRKrq+9yU
5EqoM62+0Gg+EX1p94XDxq2LpxZtuHterodymrqcRaKEXdqXeWuJsgmvSbqP
MIqTC6D2BQj1U/6D5d/S0DICLCEmXr91oiACBaDUN7jcrYaaYEvNNmfdmnO0
ogsbXOTvtN9YScCHvkF/PSiHZPbjWNnAlWx5WcPE3pbwgyfENIMfk9sxvdVD
HfC6aIWM7lioSE16LyxQY6tjasRMZps5ZgYhdGzmsjIahdAkoWMRbcEGRE4q
y5dQ5gnTaoR+/fI8GEkhz/KOHhL3Yor6y8CJgQOfY01eUtXJx1PCm/35Bobd
PaN/QTG589sucAMY+454t+WZs2h2P9nwVrLpBNBmT0YaGvftsTAywjW9u+fn
e2v8xnhML+V+i25HZAWcFaauf/vDSh5xYp15LWeByyFe4P+vBV/Qz0cqvyay
li5QBQS1+gevrCbxoIb4AZjO4tz0aTE1XwLqknFB5WDUy5rAjwbE+JoCK1sD
4W/hkJaaLwXaAgWQXgXB98eCMzQ1lnH5DRsd+n6QUqbkRLEOLrvyaRXrr3oj
kokE0uAioDSA7HIH1+j/g+MF+hF23R+ednnIjPJjHl8Ka2x+j6+f5gpDGdcV
ffaQG2VW3gRxRlzI5OHh0BrR1ZEQzh92RHXW8b6OFNNDTLJqV/qvh4TqmWaz
6GD+n77RaEAAtJqSE5Ar2vsGTc71PkuI7aXYvr9UNjpOE3o8gFuDcDMxmNrY
K3R6R0cawLq1RjltdrcbMVpSkyrp1JJ7Zwj1rJo1dFAPJ2XzEhOevI6CXmbE
IlASYgCqNsz8w0dQMQhjF4BTZnriq26fpL1mPtp8tr/fAPCWafWzWXs9pJUd
z/o8LXpM5H0IUMnot3Ev7pwMgslM/i5/DKK1EXzU5gv6wEVh4NwGIu85OWgv
56KHNMOH6bczrHFQOSEZkMP54NWALSPIXT4043cd4X4+Q0JgNw4YvD08xSFn
eX7s1m5RYjvdyCswabGUTESj4xJ+PaH6SebOR3Wq+/K6zZujeknEO55rbnGt
gZh2/lwU0MN5jhnGBQX+CCp9b+BysPKZUZwSx2ebdSd8aOF/sPbUB4moNF+z
yantRF4UuPwrAn+902IksrCXcLuSj3BRaU8wY0ehwmbzGFo7UX08mgzU6IIH
vYpgcIg/SgBVOfbAxCfwE7r/Wn7uI/4xpxHmO0qYbXQhT9KWrM5C7eUubRhr
H1NUIfHXbLzb23oaRScsQAw48+cMJi/Octyne4R3jsaUj559rpIbOU8bmAvj
oiZqjAC4oiC395R+glNZY3t2B/ulM3POQU9IXu9SODNrrKCT+SBY+KBqZp0H
RcZ+PuTnDj3FWk+C/V8h/ShuBQgBWnbtTB4agjSeSEaWNeeVXYeIlakyAjX8
FWBuczIERIsYeZScHLp+US1y6eDFcLZvpIwGHcg9TwKdh4aS40lNHdTqm7EQ
e1BlJQpjTFQjJ+QRHjvyOxCaZvJUdvfSA9pKYpDNkeRkPRbDvcE52p0Pg7/D
CmvvP3ZCXgSd0HXLPOUr+CewItvL3y+KPJexXRjqVW32LAQlEaK4ewF4H/Yd
nlmX37XgZLV1LspkXkEytvoPL/36nzAF6gUASG8xMzm7tD9/m046f5c+TSUz
0UR11vhcz33ddrac/30cxxufxjlK/N1foHSZECm2hvcg6/QzCuQBq21Uqw6F
SdOeonpkOpRL9KmG1SLn1KQh2jkuFqbfyRtt658Z8KwtJPuTstMxUs/BXbHp
1mFJ3Vy/a+apKA+VNu7wZxIkiG7kP90Jrmvx/gzc/BCskebLYptf0eofl1qj
pFDCAsU8zCJLwoQGlc2FMeRJPeTMzF5FcbOZkWlluPidyoiHNvOlYqec27ix
kxtSBd82JKit5YYqqhR6FrA1CVcA9GXPfki0xRXY1HbeisZsXOZsg9Jz4QUC
OGprBi496AK54m0SxWX+BlOJxKwNzRKkqqrVeZFS4ekrsQ9NFW9LxTjlEwfV
Ou8NmxchULQKQReyg7a0irrmkAsPPn4rc+g/OJS6yTXDPs9ClhB4Z2MAsWVp
Z9EHVYPgD8txPuFg8vK5/ju4cP8esNecx2wq++iQyg+r4w2Yfa5OIff4LJ7m
E/wZ7Dg76pJEnc+7znOKlkHFpXcZtmhRo3W2JnWoxuGBIfEgrcj31n+IB4lF
2zy7wDO1dZaVVFNU8YfKUne/TvoO921aaA6y5syI1BsHjNYJTJuwGugZEkJD
2wkDLj/iztOx0I803wDNHlIlO6szHaXWxxNDZX8lIFuKkd6CzI6LlEIIKCm3
Sl+yHIPwp+lcMTUJ6uFCk+PsrWsWYusBh9vJyB5SsoSNs6AgXQWMCwLlo6T5
wg7zr4fhvnd5kgl4U4sefgwTWnwvydrg3H2mTjvA0yMbE9mwjWxlre3mBxUD
dhYE7FJrNyX2ksqGBSexCq7W/gl8HMt9DXufsU770P2zuo1MtI4Os3eZJ/Zq
OwxMBNe1FyOq4LRUP+5hTwfOANBZt19Mz19YMeXmhYMyw8A8wroUO5NNriCy
FrO5O9lWm0tTzeniQpkB6+p4KlOOaCe1he1hXrg49pUFnpt/BjB4UA6WlWYf
2VuAQWCeugkoBDmVKxhgSixm6PlFQ54WR8xuUey8BN4UC8CaL4Tg2mcVkLmz
kJj37RbIvAmeMaudYB85vOfCpecVGdNAZyO1UObwlgAvRMFzfoAqYN7J+hvD
RuG7EdLSfulL9tFjKsKSqa4BGFmHcmcpQTAMroEiG+KLtKUJGQacM3Nn4vvW
P/7J0fJ0/LxE1EQYrbLOSR1Um787WKFmW1dxWFMt94WqGMtQO1vil4Y5UIdY
LDb9L6wYyFyCG1K75clhI1obb1tFTs8eBAFwMfQBaMKAooZfAQpEX/EAphI5
I6FfP98mHrXx18CbGpbwvXcazRX3mYDF3qgMO91tjgy96Ar+/rPC1r6k0ANF
aGciPxxsblZNNMXztzc5FsmH4Ld5SUHqRzQoMacjkWIK3yMV8Q48a/HjZzU0
ICrZqOP5Q/JB0wA4QN0HyikUccSFUPvEhZsojAwpx9tKmnzQ34lKliwAM/UG
qiuy6ezXrxe4EOvLwCpCK2cI/To8++xHTuyczJ/yCWQiJWc7+EPsY+r2umvx
4Wh0ULjXZ/UmN0SkenD012rnX3+b5+YcCJ2OQyyyH90YTZT7zOXlcXYrijm/
j1dQA52qS2GrXDJNEWCDWsokGvf94lI1zhc6vJdpjQ07DUL9Ms4HrhoaUc1N
gdrpYu4YId2JRWYhPddUtACCtnrFgO3R327ebTgG9He6JHXfdpX9Wdld7REA
m8BkjwgZ6z1dmd8IdXZTUrg74How2mwBkbSMBG1Qszpu59dSJ8g/BlRYTpB3
j23WN5lOLBNIqbcglKnI1NSagWH8PdQjE+grVR3Eb+C3N15RuFUumHUx0zuH
vsl5s4n7L+kkJWR0jDFQak6hyj9nQPh4BkjUS4hjaO8PeEtrfheUx8kn8Bia
p3EdxM69U3EEpWmAScPvCRq3wuQpfWaLb9JFryQr3KYixKaCU62nSoOgnLd6
ckfR2zvMwxW2fy+mC8+EPvSNXx4DOe17gfiP99GYavA2z1f6ZH1OlhjB3vYj
OZJe+x3u+JRpkX+J4s9ECiRiqFkAEDRRiP4KCFi4ne0Nf1WxzqXekvCnUCRS
Gn8cFcZU9rz5r4XvpIFXY/oBI9wi/ysLvSv7TFNvh+9ew6aylSDpzemxSFMt
tSBgh30MSw38P0Bx0AA32tM2X5aIBr8WpABqXPstl6Ntp87y81FwejM0JPCk
zdJgY0k7yUekxzOX0nmHzQ597fpNoUuTyI6e/kghuS+Q9hgm1u5lTbaNQZJp
/0JHcuBzRhB5UhArTiR6ixdeGOLl1kuoY5lOhrj+baKYjpITbHqFjxw1bzx/
m5nvLxKLtQo9MdQ5O7eK5u4r+JbuNExrhM12jk/5l2nvDEd60EcKCHwYma1r
KPOZJ3bIRbmr+TC6PjAwO5xNXvPhx8dEbsfQsGOm0hHv4wrjJwtGWwwuquFj
/dtRfynhkmAKiCXidVpZFSQBZyicq8RYSWh5/JbsiaWx2g4o/Y5OPKaew8Qk
1qcz/f6KVkbA6MOatlciux8J1S009b1RkHza49gzXlj8B+TyyF2roN7unCIP
TE5WFoWDY2+ZMYyUuBbhorPvpfn74CRapAmymUkgxtrKWrtttI3WYwn0kNlg
3EFsip51tUmSzg8dI2wNI8bzZsEXL2+dvHirZ9P0dtXoooUD/10nee60FsDj
9VNHn9G2BilMxMSMwNhkfMeLl9wKZ4dR4X6A4773GqapFzxNAhV66HbQ7z11
NxVqwunuO3HovqLlA+/Fz+dI3/SnFH8cG9+pDZXmz6/OlRfHMvS6SVk3n/Xj
U/CMjv+7fe0FLbxNcp7Gd4M3uU8776Ynv+vJ+fT8uijqijx9+r+J+HCt3C4n
HBFJR+24YwB0mM2enYu7l/X/LSDFPQPAUgoVE6DOS34s5q2jgiyN5+7BAEi/
Ncnpst6gwWzp6AwHLbDwChKA4OuHKa2SHqHLQQ8rm9gLMqMsHr1LMxTG8qeV
EkI/QBiVCfBhK/bBCgF6UoRYjT3k/4aJF9mPM109pln2s1gu5lIyGZONGZKH
kiQc05WhRs97KZyjtLgDQOTi0U/s4W4D0AC1zlgZg5Q1QbyLVvUxzyE6nxAN
a2HVm3HyOXJeYG9KgQyQFHxRTDTvxAMVth08eLCvIXDUqHGCbTHa1TpYtBnZ
NlokIBS8FT1yUF1qjg+nmntrpbt9SyHVE6478DaSFgg9Qs3xD/uaUBOVBxwc
vk42e+kXutbLIZ35AF5QrU9dzMBFtCvfEX9ctHRrWRe88nqBya7TtyLhCv07
jlK8keZey9enJAJGqEhdhUb3g4Gse+ZkYXNAosJhtMpBAc9qzAhAzJYiLvcC
melxdbuhlTAoN2JdThFJFA9ohWMrdD8ZNgRHhZ99RK976USZ2CSZUo19sQJ/
anLMA2NRgaBn3aSUxAh8G9iU/5nqtAXJHEF6ZEr6xSoGa+ddU6MWAwMlGmmU
CpYN0zwNx2zl6ifKcG+CVK1TMRnKrL5M+swAELchp5+Xl2udD5gF+aQVQW0a
4A/HVvRM4A3s95NhcJaaYDyIOGBs7P4tcznvksQy77k4PM/+M4GEvDpK7NR1
SJg7/AqCIvgF7eY+dJn20O2RiAc7K9DLzvtclLxqCBKZPsX6Evhmzuqb4IUB
8iGc6aflnLgxtjJ4cx3oEC68zy/WyI3x6MeRUGke6NYtrXglVVToqDjKzMgl
EBTSi0C1Pidncdsw1ZQeU1tiqmtoHms9qe9nzq3eMZppRc+VSaxaOFYEPIcN
2fY0JtVqnj+yiwDvf2ftpl2xoPDX6TTJhGIffsUMRjDrJ9eKqDl/2TdE2htG
CFBE+V/p1+3sMnpzwcACxGchhy8iWpyLziGOO6baXv5OoN6Jy5wrsEF7+nq2
weyNMshgsv2ac+IbMSJ3RS59ub19ts4NkbuppRUM0hqHtLFI0J+KwPGTmoY+
MGpePuPN90NtcRicobCAE0SGJYQCPJCfP92EWMNwrmi4O2PHI1A64a3YcrH6
Df4E6pmgAsJ16UGQXl8954bcogpcwsaGpaoGT3BtUEHENFSjqmXBcgiXjIai
BA4BQs9D2H1ekTgJv71+HHPCoIc9IqdEPvsRc26AJ/+HfTahv+nnZiw7deoX
8RVLrSv0OP0YMLGXXAmsLRRcjojvsk3sd/ZjC13CpQe6LchjOsOWdl4jyqNq
mohDGMafAEUGzfSjHCw8NEREstWXWHfcXCoOE4JEbynR60qksSIdtgQEtcu5
4GovNBttnjbTlchWK7y1yiR73+oYcQYSbMZTZvpX3FoLqr7LVRvmHNEJEWx+
c5XN1Q4b0FtWoUqR2ULPKF3w1xP9OtM1Do9W3e9pVM9c+Ft8c2Ztk5yLfNFn
vgSDg1Y2rIxyLiVCus0j+IgY2hUVm8HPSGOuQbm9LQkmLNnSBfIAgAXuWcJ4
A00RwKLkNhHw1Y7mfO2Q+M+u5WXWRg+EZRSAxZJ2mG0P7RU6bBV2wZjKLXKO
g8Cd20wpJNNPayPPTzNZZmLzeU9nz3kpG7uNgmZPLVvYkHH839vKYbje+kmD
qVsY5nQCZDbd5ADVyl/zUMoBCbi1dT+Tgtq2/LSd+FgDdc3rrz5gghkxrD3X
tB75LQwIyaHuTHfPFlYYohj+MaRCfv5uNyuskE40C4UBpzZkML74ESNDIs+D
kUcaeLQMFcY2ITOBPgHOVmWqy9UcYbVsNkrzRQWB+yEY3rrUTj36P5pg+os2
J5LIQ7QKhSh7bMUCtygwpfowLLpYY66rvMSKqaq3e0SmkLWxUWUapBPkUZZi
2n7A/kqzG4PCnl6mA3lep0kP+l4b1nx+Wi+KGwQ0k77vwgYcZPAnE2Law+Gs
UdvvB7Wf8RoJJp0o8AVKhtVYhqgmvxAw5DkqLZKogLQyQ245GIcfpQUwFHmN
yMz4+p1Mx4AGwTfXssU+6VibNdkuEbSy+n6E41BUMMicJJ0ArL+JWKUPV8UC
VG6n6/2AO5iTlIEbNu/nyqfJMeXO4DnPAKcet3NTwvF3nPIMs+NWEUKf5Hsr
X4MZy/IsHeDsHqIwpgpuaZCUVkz25uKbEnhlbptyWi6yxIggckXsASAyypQb
6oQp6I7I5PmdTUYdwDBINwb5Sj/wCb/jG13/avpDoifbe7JyAdt5Azco42Gm
ne7dyCdm3ZBPS5VsR/APHlm/iq+XmWeNSG+6xtDcboJNPBssBgUB+I51zSK3
w+OUDE76+g02ApdX0CAGyWwk/wMt2x/fclfINs/7aEhUnDnwrA8sOhKlcx90
eht5qQsknbkgJsY/0NkZyz4KQjhykwvnRSIelMW15raAdep4lFLyEeNN5YGi
pPKQCev/3ZSJL03HUomkcl68VG+5h8GWv0QSNsRGk66gHr29RZ54FPHzq17Y
GNejYuw57U0eTJNHUHE4EaZdGdYnwWFitGdxe+4gMyGy1V5KNl7tkc5szHAI
7UbN2VM/4kcW0HSVurPGP5hCSYEn5BNpIO6+8VhL2OE71Pw4NUEpLMwRDI5q
8fh9n0HMy4BrfgyeCrUYu5Rt9mwmOQYraVry8lyGgHTE1320OiNAb8zu7cMp
+LqRgvhijWS/+84x57Rce/SuI367lr2cfv/EMJXkihDplHXlxideTJl+VVNk
bbUQBoh2cBm7DGTrfHiDwf6usMbNcIZXvwH0x/JqYlUsEV56jEOlZj6p3OO3
qm9x72LupcO8xGrZxKcjhHE3xtdWpWWt3s4JuuXpnh0NCKpl5IFmax5G4yrE
J+UrgA3BdNWm2iUDhwLInufcYV8z5tCKk28LbF4/NdjN/BRXXRIIzWwfK+SX
4f/9sImElc4E4ZXq1ZI43C9kxYgWtZ2qCY6DtKyxaBG+LWIy+Q2nmmKdBu3E
i0SlJKX05hBkE6zWWJ5rzPx3jQ1CTCYk1qTu2ZtW1y8FRk8amSykXsL5GTWJ
7PGLORlNNJsGbbKRFKrZXSNHINGNDoUAqZVT6BQD2WkwrxWBhT0F6hNnB7DL
ROA51dHcXqULUWB+bLqQWkyDOOXOYj66IV2CJZWN2BH1QjxELJlS+rvoeIEI
7I6RhNCLicPhhxrFBDkmJU3gvgCRSnzojzGFQkzPnGRjgNui6eCxIzTH6Bv2
TW6ZLuToDEwbVy9kw6KruQhiXXHZc5If6XzxHfsJxw4k78EJiSe+Y6m4LBIY
FJO+QNOVnPU5Z6eARYsLMDMifv21ozHWX58fnpB4ApHH52ChHyT+2NSkanm2
CYyVGD76QsFruTkP4FZ+MF02Jznm5GgRjgsYABxbAwL0TKtCt3wEeI776mKg
H2W4nWn9tMbQW80mV3eJhTXeMfVW2NPSeMQWG/Ot67z2UVndSzKuk5J/D/9D
jrT83gxREydpgrWLTReDdqDTOplziZiaJtwtUPkV0gFTB5Qqi28VOcHsNInV
2L9EMEZW399vcBVriTiGZ/L46ggSi3czRSv+ofRMrk6NB/+yGe1HUgM9u6KT
pw7rz3YeDcCw8k3XlwUbn3bf6umFxYQ3dGLlP40CqlgfxhNFt7ESZneK98wN
dMdZoOA3pM5qpll6PPKaurEPEu/kGebH8tTMXCV3NBt1BetC5KUN5y+T5cZ+
7OJutlsoqUtoQrTApkXUly2sF+isy48Cz+wzcujJzFSOO0b8VyTP+/cFwUQV
xPwEVQdnHr8Cc5BXhhqsWGrxrjELHyrSYt0E/OZfgseDtLlbPV8tQZutdzuU
R5onAcdaNORaciTTKouPTjqPRcns72EdgWHN2Qw/lUEEakkfSff9gIb6VMcq
lPf65CtplyvHKpncVNeIa5R1QCf78KfcxJSlMnCSSuCFofVuYMPM2q397EKw
oRld28rSOjWlvkQEaauqbQyKcwzGWl9P5/Q4YjUzhNJGaxJ6YXTt+iYQV3ut
A8VkUI3DAW5tz6fkfFBNebu7YAXQzY1JZ9pzcjTM4pCIwnmEPzuCmg19QCmG
zVD+dAdejPBFkg//CReODNHhWDMHovRd44MlJtpoqI75N6dPEFpuzBs1AJqR
hC2Fhag6GE2o8xwQxsW18FBDMgGk+8bXko8Y1vfG81IO/JfxynYuu/tbcdD1
1D4oH1T5MH925jl7V/GUMZGBq9eyYF+9kEYjZUYOTcweoM4z9FzHfDNwzcRW
dDzjcEMemhg3rNvPA+K4t9L8XRQpseYzVQ2GobFvRU+lt9exlLhm+hk4cGfR
TiiTNGf61sRjQLTqlpLuYh7UXg+VzXQ6JjlKPbkb3ue+acr06O5uToUPgFCy
JkAY1GbC1QdBKoodjCJJXD86Mg5QCKjD6kiERsufrRMOQVxES7r0caNSIPe1
CWibIi7DrIhLaC55cpfPQdmYOGtnUfLs8XBN37JX6CMXWzgHJgf5mIqZfEAx
i5xUW8TI8er5gprCtXQJKWePqmtfgOWwUjqN07H3NT02ROOat3PQdnxd+G0C
igE43GUekjB2R2vRiUGpHqQvr/XlPBN9qEFVlfRW3fo01O1N4ZGuexETz/+I
B76xIK+/c1QSfOjK/z4xqGuH/ZJJwzQOKYkVQFOqvmlJ09fBrKN2u3ioiBz+
0l/SaaWq/0/VkF3t8nAUAb9tSN5m9dBk+KCSYsojriE0FzMk8VZAcmY8k35A
T7ozTm8OrYqlbsyGhsWfGgvB3NibJdnMy+z2wQmCWMG1ZWugXHOJGVznNpq6
fIbhg1w2HkudhWakiHuZIttFEsuBQD4DfcHiE89IFN6uujrrUZ/3XSA5JkkH
sdH63NvfzbP49UP1bHbSAOhhuBj0GsRf0ykWiBirtBoSCelYqOJ2ibosg/Qu
Wmq41FnA5CcNPbIIR2JVRPG8CgRDGSZXaxuwli5kl4m2fAImOqKCK2h/h6ZB
GFoOK2e1OSOYS8vmB98arLYls4MYlJAGmk3F156K+2NN+vu8Z7hi0hdM/J41
UUUZvO61Ar2/6xMxH1Ossx1kx/vJ3+DtP9TTILmh4DSdPbqJ1+RP+BhMtonO
2REvCdj2wbFhWU2IVHkIl1wQjoBZeBAWlwEnlsWpD6edlOqAvb3HbDnqXfxm
8wnlDD1wJpo7KOsfEnqmcP1fQbLJCN65HcCjc3VNYcFNMMW9N9N9xF2gHmwT
6PXjxMPefaxSUCZyxuu8CLKBAqooS7Cr2AxXkUQx1e3Szol25mz6Aw9rw+FK
pJWtX4DINSEdwVoc+CN9/AGXn6JPuKrD4soCgJ8ydBaBc0ucG7GwhzHONOyh
E8lmjkPIl3s266mm4tc+hRRKafCGwk4XLuJHpbjbKc7+gDehkKqXADawYU0F
A2fbCCBt2kbhm1uGp4sOtZmUytWTsU5RkdN8A9Jry3OUqDj2YudXNKmoRH4m
YWeucCT5Z7lxphGwy8S1ymUmthua2WRKM7cq/8VbSiaZtCR4MkB7teALd0Pe
C358XPLtegICc/hOtcdgemdloZdTODtQfoPNtgF7r42TKjxfY1vqkdgCvSMr
upD9ApODP+xlZyAqkXkYZ1/w+ccXEJGc91REBeOT2b9oKXF2HnXXEDohvQ7E
IINAjWHUHI6DR9exeatohy7YWr+Du3djGwoYqwbaVMt3EipuMEU9sOOKj1fx
LsKCeLVSncvcSJLhQX9Aywjm1PESYTTZNch5TkgP2v0yKI6EwOIzlH/b0nFs
VKvWuR96Lj4eMCCpKTtXx4irHbJ1isTHtW7iBaOyEpsfYy7pTawyaVbloETo
Gmy9U1d/Toi1vMPiggsZ3BH4HIRDBj76D4Z5ZC9AFejFbShuGWK2frF3H6KI
YSYnB3Dkpa6/WNZ5zx7fvouFx2dQwc2ogxY2MDarx/WVLWbxhBEvzHiyE8ps
iC9ifYCfJrhMGIMDS7Q+fMhc5HWHFTyGAvQe15zLS1NzN8xtjlJmFcwriNAk
0McC4Q1XItHHDNlDwFG24T7l0HHHp3xI/5DGMUhdThY5ozApJBVVNLXg+Vfo
93iGPcq9W0l0HfGRQyL7Pqd0auidxGoyzDR2kPmbYpzCV5GBviU2cX3VldtH
LxZiuDaWDouGPKtsrYQAk0zRuLecILiJKl+HqVYKJoEnntsFYgaJMvSHk5ON
OOitgXsKZlLgM/pX+uhDYCg/pv4KteEzIdAM9XZRPulXermcejwduCs8wBLk
So7KHOf38ovZyq/SCFqaCMWEokmdK/o1HxOhXyVF4Ghv3zgXKEfCSHKdBRjZ
39Hw7EBISDnCrRuWASY9PRnRXG6hCUBAdycobtuho7YzvCjWO1iWetmEd27V
GqxNAfUCUDdMQYvVgEOPo3DirxBk+V+ocjBUsMCQtVJkbKxCHoT3IL7+xz1Y
3gKVzOm3A3vJRnTW27gKSrBH31Iu1LwZ+dt0UV4WAvvJCV7OAMhmm4r6YKQh
2Exb3CoXqdHYlsjtYH+ymrsdt97g/q1My386RKCtIJk4sEInbN7aSPfyKTF9
LqSzMd+XhmIalFCpsbzTBJENJoZZDT/y+I0U7HxH02aSdD4rpIbqJcFkQhsM
yAb6XcqbokszEcOcp8jdqElXNkn1RNlNbNG7G8VWIUzgyxFugXKXv4iaGo3N
Q4f6EUQWoiQWCD+vPymijkUFoWui+lugVZJssSXRShqVt3OFvp/XnaWXUlRC
7kgT+0yLC9eFKQOhqOI04LKGleJ9qL2toff5zrtnKJr67XK3IRoRiLy9F4ei
tc2KeQ1d62VLMj32xxtvTG/BuE0WkJexiqPg3xDZq1yrrUTsXTwRruTbOB+e
I0PYpjvCHiwogot7qFeAubblazgWbpuZW+vGX8JTrdRRHasbGD3oN/RofNBw
bOzwndwnRwVQjL4MyqpSMqkrsamEuA92W80Aps0A/aKOpKc/ewwHaHAWEchq
DblBoKhy3aD9enRhZnqu5mM16nrucu2zUV+m+8ndrNiooXHBYlQ6WImkXOWX
6lLbNCyXRaXDJ+HII0PVeMWJVIRFJia760We7eJ/UkyZfBH+Xle2EqK/plpF
qWOeYLNH4mjlUJh7gDrj7ZA1/LTAk9w5FtYVVwz+zCeoT/IzxfLFvF7LFiST
Z/iCHw4viTn81uv9Y/WB6jYLo95nmOWXQhMovI1SbTSDyo/rwiEfXsXztBAQ
0Z8mJEJDTGVsb5Cz/Z2IlsrCvl5+cc+gLRZXzJvwL205ddeXDYAiyFKCniNf
Nco+NVW7xCaQM4YTuGwX/Cdb/83fuRy/fXmhLjnLf/izW9sP6cWV1jrWjlCx
IyEQ2HaKHxbaFjwuC6BSUx/bMM0lQpvcvZ3iDseKj5wk83hGjUL7gddNoRe5
2EwCsCfJB8qWWI2BchMs3YtF9eRJ1OUQ2f/mb+QFJc44djoJM81vZaxHNIqh
6NIfF5IZ++qnDervexWlsVJvUQi58ax7nezxsss5XeDZVfhUXq90byEvcu7X
jgZZbF135ixvkl/0rmB86EY1yneP7nLHlh5EicDlbzp/Dt+dTkHnXejWuifB
EaBJEZUY4ythWqHV6EvIciArLWPKWK531KZjK6m8tyv3bpLjcJyk/CiUSgqn
OCKzPgFcTIg9o1aIv+CtWF/8qfckhUQRCj866/ElcmWIWloVWDn/+rAgIpWK
rrXwpgi/1/A+vv0lHfAnJ2KOZWydvkYImKsOdfB2N6u5fNoaLOgShbELGNxI
8pebIESgTKwKp34YAzYJ1SvwboFjmLYfj2uUwEhCV0QfgpXBQfTf9BXZhkdR
TKH3ebGghS9JJArv4A/qCbpX7en0IFpWXc0h2gqzzqW9YtLv2/Eeo4S4cOun
h5Q1Xzk/fESV8Sew8fRQJu9eiE4BC+PIPh4R3FODNWOrfYNTXv4E0PEPQGg3
hf0VVS/IWJovzCGXYIBr6laEgDJVrfihzMlAQiUck83lR7fpLIDY3Suzwf68
s882S1oeVXXs34XHaadQQRo8HK45bA/VtVbCIzT6FLWlcA52mEIlTCD7ogw+
s7C8z5HZt4geXhvRcinWS4fJasIu5xxjozwA0azfmuavDmHg1HPzR6ShhvN/
VAJPjFOG3HzFqhYZk6FvhpiuVm17eRi5BxIVd70h+NyGGNP/bweOTDeskbgM
prOIdRnGazef+pGCFP/5dYHu244gAmYX0tgnVerTxa+41lgv32sylqSsr7dx
pUsNInSnJtXIUaSUJxUI0qhTpGQTFb2UlgeB+Na0eis6PCTfaXq9ep+rEh9m
66FAtycB/0e6qldsgNsRZ77sq+AimZsVqDSWCcGVf4isKTkwOOTiHltRejp+
JyqDT3+ZDTA8Y+SJcezqLTXhICgoxqbHfrtScwy6yMC5XqJmTGmFL+/gGBWk
oUmqC4OIHyfiEOZFDhMTp+6RqJZ4f+yxKaa7A1Zj/AzBiw0co5n1WrZ3yPUH
saHz1GUyZt7pM9tNr10z6V/xj7NpJ5GBQpTAvTKRc40m9aQz558fcEne98zm
nSOUANREwzyiKJ4W6TDJ76Oz2gX7uXglQsSbhczRYzkh2Oss3iHjURYO0t70
eq9ZS3d4uc3PtIPvUhW+h9QpGR0CuemrLzNFe0Yb74c9RUn/kexQBS52zvnD
GDazVZ2KrzOrlnCj00Szmy2fqdGj/qEUDMiMWbnSyYB3/Wvt0+mDzZYr55fY
L63tz6bmeBzrApSfPNPwW6eojctkvHYOfuKxvUqPPeTzczJfwtjeTL4EQr9b
6DkgV44HsP4JkFFxnEem/ROT+iut4PVHc6IH0EQYfrWK9p3Jcvhdf7u1ls4y
xKiMNKCMNdNqVAAfFKPRrF/ZliUK/oW5tYyGilAZk17TCIn96xNnl0B4rkgZ
wWEfmP39MJDx2wpeYM+VQBlPa5F8ffh2GjeGV8phXCq7LvFUiORNS0lyqxiN
bwdiAmf4FlE9ip1qQoHEZ1vzqDPKcH6sNdjRGN9MNwePCYuPLljBKTXung3M
9crV5L+EUzIKsunYThSyWWKjlvEA3lMmVjcuj538NY+uS+fLlNxcDSTqgbfC
eq4Uq5ThLe9daTGVnDCFQ4ckBo4QHWpOw28/Ec1OIo7Nab9DPc4e5m8htrab
UsiHNrOncJdpFtYecWfOZNFzHEHsAbxg2prA4kqtW5ldL5lSA9kc7CtC6t0M
X+YurhTougoR8zE+iDxSoZZ6mJYJKoZvKZ0nOWSXxo+d0yfbcIGkYSK2rL6i
V3G4YDC+/h6AMfL0ZBRzs/glc84WAqVna+kIUZ+aVIzNBdQ1j3oFC2GuEOFQ
U1QotWNRbdXfM/sxlgVmj0kdkgIf3tbTT8Q/OIBJ3wlxwT7HZ2ZpMXiY23TP
4+fDG3wMbtit5vKL6CAdyWpRdbpuTrgBvn6dNVl0oxi6OD4qCowk49Z+eD8u
FG3M+O8pkEFRH4nXFB+IqfvDgZ7UP18ljtbR5cJr9+KlUnZv4hTARzo7sJYI
Knmy3c9Sd5DpoSCLaH1Qnn14WS/1t6UChWr4qAQnRF6Hiv8quLV0o3fxH3NH
eT6AldaT7hWisDQoaIwOVbyKLzl8crNHRm3WB1TOQpPVsFWDZC35lX8SJBJs
7eKFiJRYdq9JXrIqcxY3nNQblyJW39vCkyvQjdAb/+af6bcsGcOwRs8sqZ1J
bgXzXqjj8LrU9HPYRLbtNJ97L8exKBi3l7NT9aARy6YNnWq8yJqT5bHR4tdq
+YH0hO4Zj7dt9qu+OkZ1GF27q98SDL+LDY5qGEWm2GS3puu4jdMRG2f0S+vp
+6kYrVQzjAXtqd7ZCa9hVdYtKTJueFd886d4RRvvwy3ZhdzGcKl09VEn4wqD
1p53MyZRr6ZljdALCXTCLj0q0VFmPu5lE/mKO+/XAelPswJ53ilJL8IQzWPR
Ww+vCoyNyRjE/7vX3QpZeNgMNDURRW9ST7yIyyXGA8fMpteImCXX+NROnwWF
SUWJH8MQY45MhuXMxRTq/LET5IVkBi87Gl2N4C9n5LY89vlsv9T6M48BTjqp
WF4tPktggTu3dPPt3irHqpW8skolQXP6uMVcoa8nZ4OQTNF1Bka5vlY/LImB
lToSkPRVx0vhq46qif0n25spSSQngLaOOlT92NeQ0WuFth5ZA3bLP9NP0c05
+KW89LS/V1F5874r2zwLFLFOJ6K3tnsUq2XlkhjW/KrBfN15OdXoLhtyLRpc
HPJnAT1qS9kqM9wL30l/zXHeorHzLWM+pRU8vq9ION5rwFvqfbFM1aUXWgfg
s+iMrwstljPQhGk43wiM0sT0Xs6fmlsnwCdQq5AKuZwirUmym3DO0nVptE0/
jqPAqNRx2ZYsNHMYp9LTPTzx+T3NgN7REiLayeL+AsgmHpj40xM8eDstBrKa
9uIb9GolxEjFr0SBocdA/UuRka7ZboTkvkJ8bGLEQGdjxN+QGQE98xxQehKE
fVPdXQOmhfgGrF8FhCyA3SwdMxOvFAFUyO6Y1AwMIReJJ55ejPRc5b4hdWuq
dPJEIH7WvMrz3pzv21S8VTAOPXoMBYqNw3EqkSZeRH6pu7YQ1WuoywNyfb10
nqICSINhiejn/hvQ6zpTcw7vQRBUyR/qbVIm3SuCp5oIGgjDR/k9N7Lh5noc
9SIHGjEgEtRgyvNSDQhGOqELjd/xYSw+xe/bJUuBj1++1MURy6EMib72beq2
nGQSpcp37vTCvxStE15krPn55Juy8G7aZ6NtKscKcvHeqmizNNJivI2rWMJ5
s5Xtx2t4myXeXS6xIEWSJ3ixfIQCxl5psuQz8p02UKsAm2nxmhvoVhfxVb93
7O0UzryAVYcRHDV3vCAION7DIkzVNWt+giIxsoxyQMXeitQenZEe17HpmCz8
v+is5vnqdA6ltR/Ai/IE1J9FahGHiP89KtOZtnFdRoTu34Su7b9JcEx3qaHp
ryC3mGoaCrz5JDfk6muhkDXMmVmUBZFKBUp5pE7MauOEuutlXKzlmOFymLwb
/+eZ5LSI58jFsp5TFkpCDp+OGBqyHqmJatnLFYVLD2nnPrZmA1s2Wkjc+8fC
o87dbowMICMBFROq6jJ5hr7i5Q+RrO7dx+GK0jutfjyUZZ0V34GFHdj8xPEr
wEhRc+LLorDRjhCaljDx3BZj0aBq26Yfwag8EILS9Rmd61W8YO1cDTd2mw5F
UPyBvcXMzlJLX2rep7XuZx2SggkXA7T64HXk5nVJPMrXPYzbxs3iiNKdb5SJ
MKkt6VsmF25RXTa87RgoiVCaYHsMd5theEtSiKITUqesmtlCLUJlFTrL1M+/
RrNjtbos2UOUnX+A/OE1K6nKxgduaY9GCRm9hIrRoa8G8LEfFfnvZHM7znvV
MpwbH9h6D5nimQqs5FLFFXnyw3fg4tfNDDvd7zOspEB58gb7/D0L2Dx5kjcZ
oqedhrKwaT1VxSSA7KeNqIzdYo+um5K05cl2fpZGnu3apNGCA2OuabJTnkjF
XJ/fFwhO9opOUMbgMiyxXO59ZwbgCVAl/tq1J6bHBOXI6FB1huLUPr/Hi25S
Biu+ak/noUsY2aDBOW0jMnhQbpVGfAU4K67/Sh9y6/bC/Zot0MN/tCf9tOCf
uc6FW8ui6z7zKPSpiWfyo0My/ikU/lgfEYugeuWb3iE51vzrIT6buXO+bTWB
cfi/7z6tsPySkn4NE2MFBjZJyxubL31mKgwDlWpbiNd9nzP41zjMEiC3CFLi
tf1HWjELwh4rlRMbcXRAlB0es8gCnCsXzNwIfypWOFljr9n9BiesZTlM7kLZ
KxR74jBZ2j3W9l7mjj9x0kxmOPNyP5wcyxyrP0qR53g5W4V3AZakQ4M8hMfa
WTouL9udBIqLszGlR/yt5h/uf7VYkOUx0fuDdHAZc/J7hb1mSwtofshtFFS0
aluqsmNCuGYNKJxdGAPLMgZTUhOfLsyUQJdp7KWdGG31xcHQA2bP9m/OyZwq
FCq24iV9vjRzEsb9k/DxQAFesRF6IEgykDVrCgdHX9Qf8sNzj+FcCoZka534
h127PKZUVxPWla9bKa9Ko3LkvX0+c0IBubyMJq5uWK0QM0yitvDEOlAWHnIF
7pPPkw0reRuU1F7uZn+nz2z7E1D49xdXd8o3YT/VBlDaj85O/3zh4wBIirO9
YCVXQFxtMqmsW3l7/OgBzRIrY2mTfqntRuIYC4YdTCCieLuPAQVRUQvA9D22
DVgxmC2DDndVl65G76XoXv1qU6cfR+7rSll0x2cy6ficsSJVmJ+fDzR1aXAa
zRbf8Eh6Hs/8G3dDN86GOIdIz0ZcXZ9yV3Cgg+UdoydGdFONf/dU3ju+6+PM
GeQhFuSH7UYtTOkUrJ9CV9+vt4/7lERYjR9z9dC4sH6v8A/p/gC2nTtSFHFw
Wmmacib5ze1mzKkyETnqhG+RQCsV8+Tz7wJHAqqwUC6H3nVxqEp9Q0yzA92n
FcQ/ygolAIV41ucr2MHJkXcVnlkx9C7lw8sxsmfKNn2ozc2a+tQP9ZimTsYV
f83v4uZO6XtgRYpYZtYO5TDB7uLNV8lDQXBRM6ii0CJLqwfZWB5xUpi1ZLXg
GKIMOeikXAycGcXZnPlkx4gvNR3qPbkQFX9V3+SnWQuYLEhcPa9i+QvFVZt9
pb3B0jBgwC+mh2/+g930rY7TuknF7ViZl7jO5+w4mxZ5Rnp+dZXvWyPdJQwH
rK7Y6y0WHCSFFAfFmKvr5/K8hqWcDmz5s7w3jB+MXX/JRikU94u3mngGcf84
s5Gqctaq0JB2i9GekLto5LvhyiTaBl5AZ8mmwmFRCDMvgFNM22DITJu7dS9/
dh7cSCI3IVwMByQvfRqRjsv9KSXXlgEOE5kpuLUwXIdRhcco1+ZiCIUDChB6
6rn4AlF09bATfukzWmT7L00cVhV7E1nNpmm8Xl/2hJyRbrbwGiagKDLj/8Cb
OAEllhLeA4F5H8/JbpbFhkmPoGoTxbu0YkeDR97FGPvXHmcATbYTuYJXs1e0
qi+MXKyG7zICR9gFSIdBroVwBBJkSj2essK9SvhtlbN/cNCzRn9OwAIRUlSH
mnqQrcZOOsDGZn2EmjdTIdhJP/msTmyASQMfqEqtjfW+mGCPWyBn3cAdACha
+VR1R9Kd/EPDX9/9WXS/OJ57eZgV1k2ype4TMyvWbLZjBUYtbcvbxeinYzj4
l/S4Puar+kPxS0EBvQCb903TmJfyjOyPNNBdyBBV1Yp5xoY3V/a7JLWStZ3f
RKP0d9TplB++ne+kJX4smU79Tn4St7bu9HWSnpT9Kj33rxPaNWdTKIoezcvY
hXL+IP/foz9s84VibDztC6WCzuod1Psmf2BP8D86Kq9H1Y5Z+1OAK3tLjtEn
nlrRi6dGTDRqibftyWkQ/iWcJrjhnLuKXkt81JmpEAWBLgwLImmrvWVLLkj+
z/hswTBsde1QN8SbYzc+t94pv8W/GufKvGFwds6gTtSurN7US4Q0OQaBmube
cFxsnf55uzHGgHEE628NjltkklkYUoLxNsZU6KQQkPAwX8JCyQWeHGlxP1sE
zxSEUPg7r5l5Rh3p4w24pNWHuSvKOUtFAZKnb2Qdzx1D4mH0lCr0sZKFRgCg
6Fv3SBesVc/lcnQEYeKdwLFnxCdIT1MhnKboumSmOy1Ti9mwHF32QGf9Zb+1
KxvUH8xCxehMS8Up+A1OUAVU1KZ7JAKc9CcEXsSOHVFoGHxzL3HdBCgPiRN4
JQeu8/jT3kCdJXItM7iAOtDGFrYvCU974qWdTcLYtO+3q8NkuQ5Rtf8TYlbF
Z7RMeq0N5maJ3g7+pymaSaUKlP/xM6kxaAP1mykoJm7WHSDI8lSy2nUYnBSd
GvriHp2wa2U0HVWOR9GlQMYPrGLCiv9J7w67kRrOhEN1d26tXRmWDaxwkMiA
8I7fnlzG201AK0GMTmZAJdq1dVlUPJGlrzF52MAf7HKsBESGr4UPO6bUWFNx
HXwmbfqmQYC0JUmYS+VDgsus6pOw93tnDDDlGrXVnSDvkJiqfHlk793AVHJj
jpWanhTIUcJ+FNrTwdZCez+d1YG1IROhdiJhg7xRx5WjCyPbis6S7LiNK2++
VIxDnAmVf4PkPvPp/aQ49oqUPewDPg3b0b06bNaIZj1tHVjsAr+s9G6GWQvf
gBam8tc6ZvGM8451YkN1A01eHV33XjZWRq4eEfQAS0xSE22yCRQchC+HCxB9
AjPGG6n3rRaOfrrl1YzNe1Mv5b1gFsrZm/QCCE28W17e1DzUHA+5z5l5xIty
GTcELwOlnASQU6kUlNZK92x69uAulsWZJ5PURxBfBl+OnIioljqrl/OdN3kH
jk4HGb/9h9SpbuU+Me9D04xYViw4hE1wbbALrhRVu4ZKZpoQb6R1Yvt5U60x
hGaRwbDa3s4EdK9Cg8sOVIDeLNlaXaMAd4QPnTWhI/MibZlsnFZ/KLzp3R5h
QbZIvEr2ikCFA4QjP4g/2xDr4dZaUDIiynQShMw4ZHCqpikloi6sKn2/cnPW
dP5O/OrH3HZKYVvguG7O+MNpKWyT4Ouz42OKGtjEtGoesGmk9XTq3WPS1PG7
jsO/thbm83xBszABL3iy8IEHBpTcqhGc/1zY1V+pX0qM50ztGRFhjwvxSWkC
sTUwO4LeO+0GDDoXF89fouK+0VQtIZlqrltFfMam8+/ciUjOQtUTKYwa1bHJ
aYzceC6xrP/rO6uueQ/vlSOrVU4+eM5BfWNURNnLSzU0jSLwW/z6lbJEaPbm
3ukGoeWvvl2GSlrhmnXjTJBeGXlUbLue2AgyxKdXVXKC0eyqFOo5ge+ykbIf
kNlvAG0SfVg8Di4A6nM36rRqvE97yZ40GXImdmkSkm+BeGNpD35gOCBkaDwZ
jkbhweBVlot5DbT6Q/34bSqXY6mKWk8sIhbdXHkxGylVge+ksulCVgt0ceSK
xiKkG8ZBoe3ty2s+9EUjtH484uLTkW27uU0L6m2hYtdrqU1WGzzKQAfj8HB+
LV5ikdKvz2Ckp5yTnmaq1xqWZSve3lql+ATGrmlYRUSbPd/RkATv2K82Y2Yn
iw7zVqIMwjB0SMOvYigJhRwsVD2J+/kvNwQVSn7a1esJ+YYXgMRJ8H4cCirr
JlP9ipJfuI8XJmghoFN8tT/g3Ydv1ODBCQinaPSpQy/vDvyksFGmQXn+ZrST
MSTD/61DKJ1csfj+OOUFWyULlroWcXX4v9KrCwmEpeKD47tyvfKx/niJiQmF
bk+9yPbxK/VbkZsL6mGlRe6nqFrHym0LacP+S5CZnJulSRME+UyKWn5S0j/e
MC4INujD0WCun2aZ6ozdIWeXaip9ehQF3igNqjkjLAJMxffJkeTMmiFK3hOF
3EK0sX84qZ/bAqsCvc7ATy2oHL8kxWarElr8hfLGCfoiOkHRpXgLSaJCytGw
m8gKHPAkj1PlKXQcosGU9xUF3rmucdUk+FCHoeKeBsOAR5yuG18QDVJCbAyl
19lWHPQHc4jRR1ST1SRq36qxvcLztQxx7uciIvXRROGofTCEl3iDjb8lsyHI
1+DsZPQqHYPcBzY53QZdmzNK2C2iTfaKP8ShswIX7/dXHRKH0HpLuzw1iuwa
9YGps/Vfz9qsyjo9ZSCnv95F0QiKx/xCFWz0SzU74cHmqpGmKqIr/dk3BVRx
9fMLO9c5V3hqXVmRwTU2aUHBnLLlEZIgX6wxDkbxq4WM8UzgwelGFQgyPSxs
dr2Y/WIb984C1UTaKjGPlItjpmfNFGuGMrHoV7zccqxS4ZNfm/a79CgNuYlB
Q2XGv8/PaYsJ6gZDRkGY00Yv93R4yQAfub+b5ix1yNdPUhq0/7i9S+HPmNkF
Jiwx0Wa+R2quMsq1yyhYouuut9RkMS8J+H7VODHRiGfqPrgGM2KKVoaB2Myg
aVOZP2m6dZmxP1Pd+IvOiBhxMaO+HJPlgkrlcIFEh7NbZO6BgrDiOUx4imHQ
nD2y5gpKZP5Kpyy3MHVZ6eKcbJlhLvthBmV9oAw2YdCmUqq29yEvmA7IdPqJ
Vz5QfvWLPJ1D0PvjOkjg3F2J0zJcJUyOMIYZLadDVDOZyDCRWrrEoOWbflbr
yTi+YLcphDqGnxiT1My946gUlS/tt5m89b2j5blJlqr8SqIHb5IVrPREqVAm
90kFE0THZuvsOaJskDv5xrzRzzbdFRIYGhEDbCoTXPNbQyxyeAhJt59wcVcw
KFRSlCf0L3aeUYCqtWXDKW+NWH5+vHZ5XCyz7yUOfQADgIIe9nGp99sQJQ6y
ywovdHwzUgn2K7cCol4nKoXpTUStxwO5cV81xkjgWvXY27QVoy7iYb3TRr3X
WVSfWocR/atSKA0m0zQNkkyA0vD79oq9fkzsb9muN6wMTYmkS7eW/kbhLRJU
0/p9GftxC7EqncG5hs1bFBuw0Jr77mi54sFxYmpkITFeTawe4+npwvhAikDk
co6uzHQvL5VwtT4UVNxPVDOyNR67wsX0k5bk9BxBMT39lr4L4flp/xOdnG5g
UoxxMg8KTnGY4sjjJ3kC+6+/NWhGWcGc9iS3HbQsOTVuGIASMxF5lPWUI9w5
oI4BO8LjkozTb6Vmb3bsNNJXizWMX2KB9ROW8L+tbNja7UK5VpHQy+VN8iPR
hMek25JXz6OGzt4luiLph+pcMus9iteW8h9tv46t7GjJYXfe6bBx9nREfqzL
bhSQR0zqzLWAaG92usb2mcjOiIX4YNSILAFfOp/hfXBVrp8b475ZUmSFvenS
GAZZvuy+RCgoGnWoAJVTylkx888c5Vx9DCDB7W25vxYcPu4Fr7qLmT/nISAx
Pi/7N1CLxSN0HxD9W42Cv20Fbf81tCbdMT4go88MVfzZWF56oo4KjqhctJDS
3pyEYUzNzjl0ps0kS/TnDvkz/ftMdh6ADknD+PzkRmw/ZWy25Lq8WLUb4z5W
XBohHdBDcGiRgIu7r/9U/zE22PlMgXLfnXSwlQnbfHnmS2dwwC1SYl8D/TGp
7HEw40zirXMgjDxftXQgwv4uaka4AaIf4kihEF9AY8/63dKPAHCx66YVJmQ/
spKVHFftthetTRrJ7dufncgez5LSibZyyxINoffvPuEMwjlnfb+SQaJ0Eg1f
wIxvtHAImm/iMpQSC24lxVoEi5BScFZKUGs9suqgpph+6H1clLQCJPEU62nR
L5HtjL/RP+dSJuzX/9O4tZ8NAzn4CNQcCQk9078IlxrIwn1D4f/UichL1vNq
8kaE0h2W35kReucmUf64avFiCRt0cJTFPTx0obzP+WFUwedkfn0etsTCH//y
Uv57P5wdP+1oxUaRJEULqly+n4TbjRi+lOTvcfOgEkxSzFUsDT+72X9wwqkk
TgQNc00InJGpHgJtr+5IPZ3Whi8yG7VhUz+3gUjtVy4cfxarokilDkwzInOn
Evc6YOlNWwp6Pf8FYIl3UhisePRi7G8KEU3xFJdDU53H0/MJgr7fmNuYKMvG
KL9coGqKZWG7QYTuASskYPsA/ebQGxmSsg7UCu22HuMfOgddVJNKJpqa3jll
LIYvWd5yvs1KtAeyyugoLIjO8vtcBMzzrRrK9SmaYT9Fv01DFHV8Q3n0bv9V
rWmaA0ync4VyX9EtVvy9buogec8SQYDyzG4hSXkj75ob8EEHNl1dJCBtHf+1
XUTS8hwFYvxA4RzP5Vt0/2ILWoQ46nbUKC3V5ea8fXVDsYd+/SICROdL5Bzp
n1dJ19HLygJbX9Rne+xViTTxNezMSk/QfxeA45xZAzIoXOEcIuIRfbTvYiDv
duZ0KAEqsWlrXWfb4O26FDukf/B9/N5SACe0rdl1Q+Ezt8De9qrcudaeVgQ3
Jl5OQiFNYe1XbQlL2yUNBmkhQXvUd03XWhk+1rFwbm/n8G+x9eEGGXU4C9RC
p1+8b+xVTeIxS8GptW/yB563ikYJPRmHpCbFxBNGu+zhdVMphsIfoNDXebTt
NTIOMqR68Mw1p3RV6luFkey+kCbVawtjcOWqGteQDG8KHSwyBRa95xW1dY8B
ermDNGGiIOWGeILyt8HkZl0kxt7S7lTE9I9frJki6oqsDLLCiOt1aHJ+Xvmy
l1UppXA/w7evnsPwpf1QN7kLrypKrQkPx4mFcinPRJA2UTBSf5bb+gConG1u
vG+cVSgRa6yyYn201734VGWijIB45NWLQQpd4GqtLhjjzVwhzyScrYHBIM6U
/7TpmTC3K9ffD5Jt3RhJL8kwfsndE2Ico6161NjA9QUEVZCHiOV+MDNTUeU6
2av/U8xY6IQ786gw6q04xf15ZlPDgjpRT4dItUV7GtHf/bLdoKzIkZoeQlOl
Iq5clttUICFlzAWjAs5p4JH5nnJ0AykD9T9KI0866/UiRzI5xu8rmxf4i5cl
HYzsbaV5lzhNraQOgHHjUJdh0b7XRSHhet1cMpyqPDzfTSQctB1EnIUTu6wr
Q6PdW/gS8HT9Vmm5O1aRe2tXDpgKHdShchvjjOBpPuphz8oBfda+QLREPjJ5
7nUO7l1GWjgESSsjAd2S3cmPb+8XnU/9f1n+M9nn+nbANXvUOV8Y+QAC7SZG
vyhPs1yUmFtu/vhE5ltmWJyM+ppeyhssYU4k6E5TomPFcDxUqqSsxBuBp8g2
fUgsplSrq3Gd8soWdtYh4Rfed9QlHqB9NUYB3jdD3zwn0iYNQgbNpCPuxpsH
UTqe0kkl/5JCXzQFVP9fySVjyJaV7jTuyzmOhgILNS4Jb0YuE8o+/Pgk48RD
7TIu61Ihff6rk+KBWNKwNE31CGF4OeYzK2L3gZr3DDAGX6SzLBNvszh6e8to
1NWyFvsUOAaYYsRHoMngDQQb3VZrEhEYPcFY0jtFk47exc9om1//8B5Vmpk1
4zIsYkMZE7WD6PUdEeERWEqKFXeYewQt7SJc4/DZGQDBUfuWxbUxz+IeXrKj
aJqnfqB0aRgMzYwUR8GNUWSepJfcyXs3Y7pr7k5B3nLtr5kUurPYKtUydGLf
m9xYGxAM/pKlHAn1aBKo2Ogrwz1ybqfWMmvu0h0SyNrUJZAJLw71/Z9Gm8LA
SlEyvZZyelzf5W6RP5arcJScAtzrgq2oEknh2w02uPhuH3dpkUxOQJz0eOZi
fg8APwg84tIp4xtiAtRFO4FbJ/m2zIoHGAzm7aQmTcHZuV95LtRAsjkhD3hF
Xzl3Uqbz4UISzlZJFJyRgHJM4WNXnvM48QXZghho5dJeCj0FYz08Kq2VnIUq
r3SsmXtdKBt6S0XmmyA+D08zuGPTO8rYpM+drVBYqbBIkxMsTof37zi1UvlA
uFq9KXWAjxVrYmNFRyA+1YO+Nv0cHXavXqrIKl9s+n3i/PzDjEjjR6dHxJa6
bntmNqgqyF6b1bNTcNvs5No2KnNDelJE9tm6NmMkh7s0eTwSMQ4orxXt1Yzd
rbffb5fct8oB5+rAXJmiThV8hIUFAX2VQNGLArnwpYgWvCiE8pFh1c0uMrDk
JwJBIW0JQECtBukC5mgubIWIRmBdZpeyBqYYjT+3aja3Wnd+BSi2OGUaWrvZ
lcBcgEw2K7rf6WcmVBXbNwrBFCKRK2p7eclypAZv30O+iogFx3cz0UlE/tzH
Lol6fZDR6BDrOJooktPNGcd8AXdNij5uCa3S3hw2OHhn5RwL53QH3cfn8CaV
VwDQVjC66iwz6sYskiSMi8aKJm7ypI2SVOVZwZSKTmcgF25M1TSjIQChnExs
/5lH9DuHlyKqPOjd/6SuXYRu44icPyycr5VFkIv5pNkgoIV7TshIEM60srtJ
jhU8XF1sYnyrcA+khcwTS4ukGaYAf6crMh7bHjV2kFlD9pZS3Z9+rtUZZ4Y1
bNsgiyzbhpt+Vm8qEdSQ0ZOsrWlEz0AKY5lmXCQ1aq2CRUmQN8L5BEzCToj8
sLXMwET1ShI3vnYsoGYjGDZT8Ki5yB/bsvX+mqkrPgjlPfyt/twNRLB+mgDX
m4A07o67SqpPzN8IbDBN9qUbGPn9ULEljRGFlks9HlWozFxnrE6kuFFK4F1+
re9GtG/TPMhKmfja6z4BkOf3sNh13i2KRf0yfiWtQ9+92+frdPo505bVpzH8
W/gTKZDe2hZazgIMt+yEbKR9fxYjTrFElOipsZQiMZtf5pJwwOOmebZW+Wjw
nlM+JbalMeHTHu02eOyW1kFT7r6Rzl3SvEBj86TXFeA6HqWMwUkWo/NUMEnX
t0w8u5oFGqGn4NPged3YmLeHtvvr8G9xeWVt5qccJMKI/1a28tUAqMWzr//t
QpHN4Jvt9o9g5Pl/T9RoVHkJQY5Y5WjmVdzcMluGtwJNySCzxtCQ4/j3codx
97m/XbxnrNmAKz7vGe6JXlTibmOjZB4ZEEQ/1GTu4u7j8rjCWfynKbdR9CAX
+Ht5C+cs5K4jY1Lq9DV3KE4mBVEN8Q++/yx1F4ZEjBTE3xw8Ixi+4i7Fasxi
mZEQdRMCA6zYSURmKtDOM4io7KewNEj8M4BzAXrxsADduu5RgXAxu7j1XE9Z
T+BzdVDYUWTGANjLjwpCvJSO0ln4mSbr4UXB2a+iQfPWQZQbMFZwKTuOZxnl
eI0T5kbIC9a5u7XbQ5f75nPRw5ysJ85emMHJEbyKQUMYgzydnW/Xo4gEpHWy
HFe1n6Ox1RyLaVOXjy/+idDX/3/AJJitCxrwlqzObEWdUhsRo4kTbU0yGMB5
yhUiIhJCqZ8DFusczC4thvLqyAHTHFR3JGAYNw1Mu2Ho86sg1hL5fpotEQJd
9vvYo4moyZWrTA8dbzirBK/mAruHeyM+FJv6r/yBUN+0EOublbDGB2hef5hy
J77hkD/haMzc9LK7WcLLbRdSkKyI9r7aFhZIUEqk2iPlIGiCVdMms5JJ/TEK
EdpRdNLOTJCIxkHphv94rqJHj2OAElYi9trk5YmAZFK/zGomxyLhy2nMXpsk
uvHFv3G0lt3BWLlTlHRT9T7RN1meBj/mcze9DuE61IPZ37IiItTL8oM0k20B
vIlRBI57ScVXBWBmGfZENlbMV4EJK+dILyTAnoN/tPKTsOd0iwUHwwNXe5jL
JSfZQHiFFq1rcm9rN4UuMIlG/v3/Df/qs7TTZykSnS63H8oxyjOLtin9qhHn
8gthchcdLL7ACb1oUD99D9gko08AwPRjcKWZjHrPEUvfjxwC2LG+6hpnqcuL
wOtd0WUZzHLa3TOBLX9BQASZwR84hTeOvcifRecETu3s3b2OUqe+tqCc7FCc
pTrvyshsZLcWGXwSxRTWvbvz5rZHpwk/jZ3rmGdueRaKsfU3c824JV3A1xx+
+t4K3DdxkGb5LpDdSaqTTdvbzF93t9gzM9dwOqG4RLdS/dIEzit4s/O790bC
Iwh18IfQf+QXVeKEBAE0g9JOVCF0GadsIYcgJuC1rxJvGIw9c7FUQlsZBvDt
X6G/qRdvfjjM1O5nUsRtNLQtBfMM74VcCxqQOhfnOoLc5kVxVIlbThQRAi92
s4UC5GZeIff0NQhaebVH/Q4CQeVmSkDvDQ7IhtBZ+vZwru/yePJAvP6t2S9l
Aue52/9w5pLOdytCWoxaDP5sMS+/l3k6/MnGyh8XTgtEOUeFS+QghynBzPr6
LDi4sjMdTBr4RsNjXPBR+4hl9F3YPB/2wSzFBivSG7d0WIwfR2kXYwU11AEE
uoc/Nx6Y8ErCe2sA7SmrFnXYCvOqPFrNy4KADTvLlB2n/H8Pd37Bgva1PkyW
io7953ISVUkMt5XJxUzb+7q3zjO/CC4djRRq11EPIiixbAssUiSGB/ldk1/9
qxeqMbonl8DhLov+w0GAupAP0sCBHry6sWho97FSAwAMU4fLRg8TUM5FUXrl
kqA6daCJ6SAUxDD/RrgUtR4utjZ4JJSIefkcBruJiz+gDyn4zwH2aQ2fyxXb
SP2KhwVubXLPFJhe8C0IoREFfY2/QR7pJBwpkNT21LFIS1r+ASR3zDFDvcD2
0suleDZHb4062D7mnqOfWhLmH+p3EPeOjPxbyF9IdZacKlXYmPvCHRXZumai
nmb/wKjVfpDiLhPDjDDZ1g5bEd1VVcvvjK/mJvqiip6k0tMdlF9by/2C5hQX
RvwmGrsROZ6FVTFgdY8HvaXdnIb29iRR1nSi0eZcov0u8+lmsHtxDih9MN8n
FVuMHBOJDFyr2VY0GtuvsmdBl+5Ku2luE8/GJ2idOH4DYzVTY3Eiixu7SBXw
fm02+rJaoHnJVcwBjgDiH7mjWTnR7ZXUjxbLkprZi0j6Z24JlkFwew767t4S
4R5rEMClI2ZDlAGsgiRHLwj0fCR+X21o0LmicRAHyanH1fKeMdrY5Op2K+Tz
hsp83/CMglLYIlkfOxfvrph09nc72GSCBzAG9FeocDx5trLHgISFYlkgZsZT
zdNGdP7UBogHN57pD0smLwWbBrnfZuykhN41Uy8cAiv9r4QRMzr/kDHuT9MY
HLkDI+m9nl1wSHqO4cHSX6MQsCCp4zM13vdAh9kj/GwOLBg3r5TTO15ImMfF
vsIOoXMx6x7A8c2krfo2TRgTmrpVnZ7rdQlI28zXW+FNd8ANNiv+107XSHUn
9//H5XEClS0qS2TY5IGFvAeZ6KTj1DdMMoOhSVoLQq67b4T5rryvARaZ2JCl
7WgjyAoyfjexnbWoMJkQc/sbVUlo5Jr8X+ip6KQ2WyxssaeNj7UOrTU0ZvD3
UizpYPUGogLuLuG6aJJBFWMo990XcTliVa9dy/s+ZzIvfvydvAjH7j07fDxu
LUiGy9dw/6TcOU7bfkZvkVKbe07Z/bNHFADh5xv1/Huqr8QLrbOSkfJG+DtU
D9crJ6AtzzsJQGF3Ea5SzZV6PN9kNF2/e1J6gsRCE1GHud9wiaY6mUe+8Gpb
+ECkXpozoPolxwUG4BL1d0W2al4tAGapdGkcixZYtym1NYsHmGkT5Hv+wd2R
FSlbkpdMkbusGaO1o5gfg03kJUhLvoYqBLO/mGaIIdrjCWj4wuSyF5YZ6MAk
sLZzWWEVEAOii4qpkDW4EcleLafA3cJCbS2M5yE6aJlLtVI4J1cEa+9NUvtd
mQhgafcPXa6OoTSILuYUpvfj3k0QurlOBLx6GR+j3ydpcs1Bd2tzzi5Np7L8
LcoDSXB+7RnwEuw9ZqinPg0mYFaY9K0u5UDUsxwVt+SD7LfbZbyqFh86QcOg
LhY4TMYTeN1/yMa/NNAEVLJN4fjIl5lYkjZHiyhJpBs6/hJFYOCVkHsypdBM
de8V7axBsyM6W1jRtwJROsByrwiCy8gPH0L7td8e4RHl5qGQ8kU0O5K+00VK
Wa2Tvku7AVHiS810lODE35P91By4xnxRgmI0AHHH6nn4fUg/6yq+vD+GmT6z
r9c3jeOdRiC//8it3zn+TuM444w0Vs7RbleAe+m6tkuGqsPhYAYP3SfsXfK+
eiSD2d2LKQ/PbH2KGeeX5dGIoG+DlPTNonwYh79ZYIEXDINaZuDLCm9PJVga
INTGD6Jld+OWAw7KxyHJDtiYzmmjAetXGhgGb35wmQ+vg3TI0Ll8iM9Ndo4o
4LgmV+P2ryHUZ2ZFYxGC/I3youFdhOfOKnRoDcZxuEZhJrHG355KX1K/SWKk
hky0DFo9RZnPN9FOT8ni3QihtDIMluJ0C7ivNn2O9ZzUYH+U2B/BQ758KyW0
4RRx7qiyQ5Dw+j8tTJ/SauIzwCiDjn4fMvsaquzOL/tg3R9GWp+ATS7xiKpg
Q7rU1IoDFTfQgeq4ovf1PZQaOSOaYCR8PWQI9ujEc7tK64Yp5l+ddvCpntID
ms1GUjVcMOlINdvOb/DpWYbZ2VrH2k239IW5YEINB268OyQP0ZYeBKvG43lm
xWaf4q4pqn3q7Jo9DGJjVQcPMY4v1NtfyI/OYphkYk+lJvhh1dVDBfDkP1LR
Z1HvybSLsjy2ELyGNhIIRPn8eXR0oYkNXBTB/5x0YZ5u1g/PfXYLQFFIxPNk
fWCGEvUa307kfo1SLg5TdElann40HQYx6zwv7DR6LkcXZRku/5iBaw+u6ZDF
TrMyOZMHG3t9XmN42uYWIa9b3kjRVziH/r2lOvp17qP+R0gg1KBUBTg5Oq0w
s+8QcqCZBHDQGXVconw+99rSqrfYC0XKaeTjZfRnntEfOE7lVAa+WVFvvoy+
b/KHie40wHuGSKrkeo9hUb0nzvm1k2PIbcZ/dGNUOePFoNkJtHqLfNREp+GA
3gZjCteffJf+2D83n7bv0yF3iOjQ7JeaSD8EvC7bwWPbBz6FTY2dAPZbQ5o5
xhSwTgJdP9d67YsI6j2gTPOspAtbIajRuIBqaIrf6tYH47i3zhhIl8gKgOXt
lR1zOOFr0RwlKS2RXFBYzW1K78gkcyO/ThQVBpc7DrI53HnAzQW6+RuYjzKG
q0/6HmUZh/kWc9Yab4up8HtYzbFBlz1H8oq+IAGu5RHnwz3EjCFDsu3QbjpR
an9CsO9ZnaCpg2GqnELTWdcJzPl5SEkrJ9rClBGz5rF8Vid7hlDYKfd58/bm
+cdWOLZMsnj+rTTbbIswomppuTrgbcm0r/P5zw+74ljUsGDmIWYD9Yr36w+d
CI1GnBtLsU2mBXohbJGDgmtEjLurKxc/us7waQQFISra0nSzhPHkAW+tGJrS
RiOhSypaCKsa3S/D6Xw30i/9AdGDG74lLYquSPOffmY2a2Qw8JTD+iAk1icU
A097ZG8+P3/rpxR6O+Q/9K4TaHKSy018qyt4BG7x+AgXKz+wboRz5PkzeatF
w7MQqeX17DfhBn4TEkFBvv/lloEy821/GMD9ZO37W1qxuC3HuDPN/E+fXR2U
4NLxRiBe4ZN6JaoWiSmVloHqd6GBmL7TevApDfqnD0u4TB+P31lxEsfetrzw
oBbKsXIsIf4B4/ayl/c0MbNQMEsHN6JxGKZeh/AOBK/dkOTiU60TPYNzJY7E
xjrSdJ9stgeSHU9MK0hjN7TOnlgeIuQ3w/KA3QNbSum8NiGVqF3S1apqZQPR
lLvkVBxlns8JKK3D02UDYKXSAcBlQfYrfrZNnkjr2yjVbzlC3Zut5Gc7JBZo
McesLH3pjaULzZnWEbkiNCq0b+VYDnxnskLiwcc41gMbnqDNbC3c24llWNYd
5Dr2Q/RU/AhO9ljcoosQgp3YKAuBqQZfk2lB4Tk90b0TSUEQgYjRGUxzNSqz
/qwBcD2NTZQd4yF317BHcEgDXaK1iEP0yi+WNCvvs45lNY511OCNHsAcFhsS
wEV/Oky6d5SJ/92josjt/r3y9eZIL8KH30MmoAhuxcqupB9Zx5LJDmxWZ8wM
sD8ETHk4TmJRiScmuFBlU4Ny9ZzQPEZuvQHCRECAJo2UqmmRDCyUaXaOR02G
7l3U4PdBLpDbjVPxv+qi1JO9m/iaLydM6Z3GGprwj0pjyFJ4WMGrFSxjqT3K
B46rtRO3yvjxXj2mraTY+cg1xW9F54a8e950PEnqQP1XsgWlfB01Y35M1wDh
RvhBXPPoAFAxCz3yAQwqBRryONqsSW96UeFHCf/+SyuYYjnq/6vx/oJtkONd
j4nvswXjBNUUKDrN91AwEYP+qF5fQKCH/HGPfAg/AGmI/IVoKkLSYZmAj8da
/NhsbFK7RyhX8h+j9j5d5rz06Y3Cnp2X0ORdeRcloeUCQq8v8St0cf7jFnd3
GuZJvcDB3o7Ir8eyNvHz9+Sysy/zdtdCQgLEHKkxIn70WsS8/yeozqIvge59
pkgdCXclRsXGPjhIk6rclXai/yM1L+AVGwe3cjFM7QqZRthMrUxT+UOCMI5c
CjCZ9dEvm4yZxLSAnpGgz1rs1PAEM1xr5B3FJxTeBMLoa8TstQfTOT8qfDOD
9b1DebQcfr1eA25l5mZ8jLsn5lSRxv+2xk/tqpZLvvyo752G5DxxAf91FICI
Pm2fHpMuI834qA/Yu6Q7H3W/A+FIC3bJA8fGuC6JpjSvvQZ3N/s2nJljLYxu
0vhHyPfgkhIbP985OerL4p898Vm08XhogYmPbyd+W+0x5H+vUlcgL1Fv+8bE
ddCXy76g5BA32XHZDGb0yvrpQz8awJA3tpuyWtiK0j36/FcOKAnfOtx6VU7O
yfMryKnp4FkPyN1ctzaCXWTrFScszw8bHmaoyT4JVplyKM6d9AnPK94kyRlW
9b5x+m2dlMNOURdkw+wat7fFzUay07W9VE5XO4dr0W4VF0ojgJKLA1FsUzos
6p/hluxZJ8LZnyY9N3q1030GFNCUj+2NU0Tuzsyf39uJ1umofebwebFGwzm7
JBh2XbSEjCPCxlDVFMhfV+fYiyuGgWF8TejIa/aCiu3HaHL1hJqEIFpWRa7n
mbAKlT094Ma4/SaqMIAOwRK1DrI91/S0DhxzbEgX075DdDaDosI9Db5mvDzd
maP42bF+xhnRb+dG39V6/4RvuK+GL57aTQntsulFc99dc/h/78ZiAYZ1KDqj
Ky0S20obecXrYyNhYlB+pdSVasM3+2mxS5HkqnYZwBkdZNVoeA0cGOTih/jO
0qNy/cy7aH6hkuyWBKZiyLXfmecwpBUYAr/ZYekewR5o+ATqpzPXsuvfNIwk
LKnpT1j3XWL4YKZbFuxFml8QfSZaJ538Z1rPpG5Ou94Rni48tTo+7al3AL0y
+WZFja4Gkwp3YGcpC7kFnb5AzHImZMLOXdC9k+2xdyulBYASTSkdhmqVvUmv
wGoPvw4FzO2XT/im+l2vc6s2MALbE/ACB5/GG6O9eFBQrOMHfDwvPT7xkhjN
5v7HMdTW+Ze2Fx8q7yWu/NpyYTBlek+ypIVK7cX+dvk64YCHtvJ8qq3xEFOL
dpeSJjPo1BXsNo3akJCS4uQ9c3zb1NNzBEvlGsIFKvWMhPoz8ZisiBXXGY6h
mch+FJ2m9MtU2JBk/fP7+0Z/+HokERFpl6u55iRnQwkr5t5NStnfoRss8L+r
sE4l64kRZKmytcR62IOTfBJMr8b6GBHRPgsSJLBpynJxl4dcoM0co9ArgECc
/dglWGtur5HNfzDTSjYVuV+S+gKNjT7GQDj8OB17oYginlpxf8heC6UMi34U
Ma6X4rfTLN5Y476u2BHwySAxVKikl4Q2ONp9PcE32mbGaeTfWEXq9Q9H3R3h
HGq+y4OLDR6vwRBdL+eObEzj3/DP/HRDm2QXTCxTHJNo5Ogfk4ihdqlNEN18
PFDqhSxXPOW/7GsVzoWwsbKm5uDQmzS46tkeMCdmkUNeRq5qTwRg2b73hpLp
FDk5f0qaIeqpOvswftKVT5IzvRCpKfOiOMAygUJIYNdOPESmysHPW+uXGOgi
zEEp7T1fkCXoPZM8rdJKG7JvZL7JQSgoNuZj9+y7DifdvvyWpSxMnknGMTh5
268wqdkfYptHYdK0bLnDaO3VuJ8FwdrEpYoyTVbNKMhoQhSzMEc4jM3pPEoR
YWYY6I0VxaYmUs38w6ylLucscJa0NmX416apLjHpP29Ob31mUAHClVWTun1g
yeURtUCpSDsBtztwYHSb++IR/sM9Cb+dx1BiNNtKU4MOalhKKQW1Xj0hNbcP
Cz8DSNOsWOlbngepJsNDX+TKnU1Mo4Tl00vUb8M6dIiPnjriA+LHSspIlkdI
6cKV1GAmFQirIBEi52SsN3f1zYSDzyo5ZPp3TW2d/DtK75ypISM8vGff2ISb
Jtt4JF7ihrh2SDXZJdmfxJpuqitw9DP4oJjTNa+FiZf4asUl2IaPTQGMXDTC
VeOditwo9KLuJd0ur2ThdFtfTFAB5VQqFASswXXOxCqXPj/uAABtk3otO3h2
q/JTz+oldMdW0UnuM1ed290B8a71BwTjIwMoWb/dXxgpFOXAldSQ/zp9LcGZ
m4cmct8xpqkrh2lWFbNUSxT5zxtNnJzLPloJ8PWuMQ0Zw3wabU11YILXf+Qx
WIQDSQ8ftev2H+YBRZIZE6MfLu1wgfXbAWxeeU608d8GDbErLANhF113dR8c
zZimxJg0FXTD10f4v97jDmJKp4tvdUgbUE18YAdxJcHBDC4gtI1w39nAV9A+
IBSBR9ozifOXD0vd30dIYIoCysim7NCD8NDt1y1e+zh+dgJXGFCfMbwMsIYm
1JyyK2Zjlu/1vyoDPlZvJupJ5qUv/0cbTXiuQ/Qsnz2YW11bGUWrURziMAFB
8vkQFhyynCilEsJVKAjBh7RT280e9zsO9lG6C7QNAK+rK5YsXV+zRbXKuciF
b6+L7GPrpL/kP0H+ocnjA860AV+QcViWfz1Rj0HCpGZkX7b773rWXu8d0xwu
nVZKgBSszrDGLD4/twVy1w/ycKtZo3tCiIhlRuO6fxUlxFlw9/sNUVmOCon2
HCv+kEne/ApGAHQTFuRjcgID+ojHlhSyUFjWChZW44qlnA7ethRrAJ1sBIJb
BsqqUINQd+NpHV7J0+wXuZMavLKuxwfR2HKfirksQorHpK0lXBvHJZDXdf12
01GyUlXIdc4JD0tRYxAPfuElUCgWYMLwIsYxNQ8D5yGYxEFu90bQlKKB6008
wWT1bRoWZqbf/8x2PdDgXDXNDlWs4JLyFVdkSz4Af3HFktR7Psj8J++4V7xm
iIt0q/IImE3J/XySImpGsf/1LBtvihVTeGIIbmkJfyADyM0Hhfn9ntMs9PsM
LD61ewu8pnnHqvGqoHGdurFpOEgwOWuhmao5HsnvngwNm49kk8EYxRaxMtlO
QWsERPszXK9CBVN00MoP30TnMHXxjMEflS7iubH54M6H5Jly1XhNh0hl6Yuw
KDmND8yt+ve+QOgX5C+VnilW5rkRqaiD4WFHnYjrYs7yDL7u33hyx5Ao+zji
VahadVkAiICPDmf1LlEQUmx5fC71zG7U7MfF2/WiRr+nGr5i/yO/MBgSG7TS
/DvoKfoZvwqQHxH9lrAzEeFeg1nrBfF7vFtQIvogkY+SrDgeAefBh2APCPq2
kFf22MvQj0/eHX082MKs3e8arFDHzrEDEWGl0RLWIO/9QI7l29u1kb88ZOKL
DfxR5VOSCrOxWErscn6Gpwo/coz85lYX55pPAKim0KvBURaTa+8hjxWYXde9
z3OX8WUJM7r8BuSH8+iHLeuWOOD20pg7VEhypBh9T9tAZHf4YppberH36Uen
7nwBepcJzOhyS9j94O6jxyy1FVAbxvgmWq+VPu4dAGLCJl3c6EU+qcvz9uOJ
29PfmWhubiPneM6Eub6QwLFlOXH/kxZBHJyexLPihDL7gjwpTYKSG2SZ/Nwi
WUEer+7M+A/YIXLpK89zU38NhMDH9rGq8Q/Nrcu+iH4v70iN6eVL7ayHwudq
aaKEnfAJD1NyaLExdKs6sdgOs/o0IyPz3qdpxIhJExMJznFnOT6ge7gPNeVC
8lHHBJa9CQjsrgLfim+lh3T0BaXchX3fY7XanxbKLMW9QKzKWKBagg7fPdZL
z/T+d3jKCqazKEh9d5mtsrFEMGkn2LfU+1TDLAluAr0CzQ4kCN2E4R0xSQNb
MOSe2WeXXjBwJeqigF/U93KswAE8LeL04C5cqVhCFVy/FP2B+Aj5IDOhegVM
M/8bonXvJVGjoaUBWlkfMO6FHyPRvfLcwiAo9NtrzJEMP+A6QauiHbBubU0t
vLshiVLvAc01AeGFr6sW8aDFRDnyRXrKEW05NR6x2AqO/h9UdbJmsCQGS6sw
JpGQxdBVlBkXOIysvtgo38rVsDjbBB4WfV77aoogYlEvN5GXVMsY3KtSKBTr
tqKWQPFA7XI11qOQOGhlGiinL2KCLMAcCVexifqcXYJ/P3ggUU8aTjto06Ag
rSSVluutTezkZxa3R2/uv5PcdNGqDFN5YVJM4bjxsP1ukrAwveixjIKB2rTY
9YuAuT6KseVtuNRDPOazXzUi7kK+freB9oHLuGF4bXlra3SmyY8xg5T9VdAc
FsvoyzVwhK9BBgLHbXQ8x4sjw3eT67J06uthd/y2jbCbYuClasOMn6FGrvoI
GH9NrIL9NMEgC07Y/oXVGuZZp3C/NPxfvEbApVdeWpopV0B/4F1dgr5LAkvL
Za5UBfo7R2PgjR2HBV6FQpNqesQOYZyNYC9HdXxvqg8gN3BKaHLnmFlLEbst
EB8Ci3/+IP0xJEwzZPxjfQOmv3ih54riKBcMjhpVa2ZXRAyPiFyAhk4tXjXK
U0vYBhkAFr6NcIbKeGmxy4uWWOTa3vunYn6aj16XefW2iSXd2fOPN3chtUc0
etnRvrRVWYtwIDaY0ccWAcphdUOf+KwyL+o10+Me+sJflaUJ8w9yuNZs8Vrd
Wiuqw4niQ3MSrEFL0riAxVft+jWhPDpKMjtFBmBnXXf2j9fFNdqrMTFZo0wA
2kX4gmRyroKtmogEJjac6FPlNeIOAAQmKzW/IwCMS6u2CeVTRoglMGFbOZAx
8Vod2vJLawIvD9IBp5aDRb/z7Du9Ti2e7SZTNJIbiH+Q54/flrMSPvikwIvb
teD2lqMZqwqspDxB1b/gFVeJV+t0AO3Z5r2cHifhjFEBPQkq/4RccZYvBKta
d1vMOdDl1OUFkvf8+wvnD2Xunbm3lBLNJcOj2mjLzoF+TTr+Domu/eOUi3H/
x2AB2TofeU+tqt/9qEl96O6wAmS6io/QcX5FtB1+bLOjYq29Fep522y4LIO6
5Vu1CTb3AZ6K5YkjtzZ+eeMJ21Yugg/43LakEoKkg6Rr2Y6He2gnhHX6gX0w
WAn67PhrdiOP0fcpdjnq44vEmnCBN8egcS6vc5Ito7e5mY+QJR7QowNLkaly
ANNrcOizmSky/rdLSfL2RPQ2I+FxpzI9WtI5YXbQ+CqhVjgYsJFTqXs1+oyI
atU5uUDgjVgXR/vW8jLlQkOsWmkuoZ4aJu5Nce99nFGlJBQEc7v+uN8MCDxL
trNnnHwxzH67K9HDNmTNx7/Pet8nmwsKi+xQB07IUq9GNgstZ5HIJgm/Dj21
HTriOIwNNKJnjVFwjYKmOGOwYtGZsYt7KZm0qQY8bhjhh1JBGcZWLcLikjAW
+/kos/tao/NZFd5eNz0wOS0d/UHypBM1Wjg0sy/kvBPsx3cToovZQUg7g0jL
Dj8zgn1dLOKQ+piOVMk89v9DSRKe+avr3/jL/j9HOTuY/S3foaUcmQqoXzX/
lg0syXewZmEzLPFojx+4suCnO1stuj+oD4mtLPzBwHtkFF8pPoYH2NNFZp+V
XaClAjQQCOvIV7KCZmLT6lnvO6iRCXZZfUaJlIlL0Rq15b7UL7kQ8W+zlR8v
AmfR4gMkTUe1xbdFozaEo4unVPI8LY0aW4ONJxgLf15IGw/s8yMFO6CKQPjQ
b2FKmex/LqtI9BYki8zq04tCsa55Z768xvn8GkRfVDm3U8IS4C7Eql0QezsU
1LucVdApUSXdnC3cX+kiPlq4aEAhfm7knm8mxmXH2mlNapIwnhiJYaqCvat+
p4u5Ib7N6v8e3OUAFNLuGQfdzXoUwU9rEgCaEgUvuRZxMvca3b81DGuXcFE9
VgHBL+DfXyQOrQBhgZLLxCqhuG6pVUmTf86Z8jltw/6ojNXeYT3qYgVV0Ax9
KmDkXuingVgDo5ulJy0ijs53UNY+efMyYpdwQyxCB62mRTYpteHVysfC5jcP
5KiyvBC0Xg8qNtpJkmbL3RVJVipbwLGq2MvvxI14ymrvw4ACE0ksZaOnUe1k
ur3B0nBbSv3ZT7zO/eewKiDJtAVX6Rnb3Aoz9oarJlG4kFeXz8MeAkhzlrvq
Ot9JnpCmBLasP0iCQH6etA8G5PPCDcwGzLe8LtHTA5XkiioyOhM0BF+oDRDW
YDF5+NrbdqBwIBOnpGdNDHAgLLogvVJ9666C5bw25u14BDgQ9eokOsfws/vz
719a7LcAkcdmAqZHjmgxtAwYw7QxL11I40T6QNKHOsucz2RFawi2StZuTgaw
G/ir/2inaHpfDau4PlP7ZXBkJJG1DJsxerik2brB4v6EVGf8UYquvs815n+w
wwo96eueIFuG3PlHpITazIYlFUpXt75T+1pbAf/csnxJb3HrIhO3rlNxAIAn
Jgw9DingC0FWK5mtEi/yeQomGjjzSCHd9Gt/hu0vGM5z/9w/dZjZMh0REHQN
pRnWwuYq4bISlJufPRbPIqxEC51JNYLHANmJHmMKbbpXBITRrOC8YUl8moG/
MSvOAhRqmN37SqgfnPpmlOZMmHsTY1tw8tDBC5iRjLl/T8l6P405GcN9Vi/r
O3iF6areTI37XiIVjKzzvNysUlq5imyIOhAuFZnz9m7AjWcysxgopfBnGZgC
wUpNRdLuLDxlOdPIXHI1DTHE6VYIP3qssmK6Gj2twrSonYqw7Us3gSW1Xq6n
6GKUoqLfvsYWwdvjkkiPVrwQHfvx/qFZ+rvzbKeHS+0HrCMQ2mo5trC1gszV
Q0OmA70SzjhhtXmgJjGX0BeIK/gUJvuWx5ZL0cfuX/V3C7hyyv+7bUryH71D
ZACXwy1NfZHoA0qVhRK8Sx3UKKcv8ddkQNppcFWm19Tdt4fIoJomoNkDLzXw
tGQYwrNQOOPuRpVqYnOfDv/hKSeRw8XKSsTayH0FEY5DMr+k+Zx7+4AWTpGF
E4T13etNPQC+p36KSNj3HtKQtOXNJD8gMbUafZ6PdCzL28DjvNdNf1PpXj9g
xPC/BkXShh9iKMVR01jQLaGS83yMmYVtoznQBslzFay8hEOlOTEF0ldreZvK
/SjPX0Iaevt/kI5dXRgPidgu2sv6Jqe9054HI/KvAh8ljF2XY7gCcRVIp4vH
SS6xtJPLHRyAZ6ohOCZrP83TuK79ly9X2P5zHOlJQDPS+rVvVbBhm/quGVwp
sUA9syVd6kDj5A93dwAxOEJF3ZDmYXMS4rOqNa+R6zOghsfv4OGAa5pJykjz
kL8OKtIbFqRGtbdRWpHn0h5UJSojfNnrTjlgdqat9NBrjauU61j22NbAXfDK
OfLZIbFkTIGzolY804jLj8p5Mf30AvssDaOr3gb9UiZTyp7VQCFhwFCMtiLY
08lpudV94ZfoFZULjzo+uzIzn551x3lfHqgpRtn+I6q2CQPWv8w34gQ9ORfX
0yrzmhQdOqN3mmvBkT0lJWfCo8UmZy3nMp/D4p4I+NVI8hy2Edgip/H5etmP
4y77FNZrId7tSLyFIImrVGsRGE0HkZRfLD0f0jR0THrrMzqewoXxeDALRUJT
eCh0c9eBJYSN0LypU9ElLAK05NCIWQTufKyeKxI0d/3GjehJX7PMsc4e424w
3cMy1DP35M0moCzVL3Egxa9Km11f2WP44yYpZLiucnUm4DiKxhq6MJP8G1O3
dpVz0pwsmyYno0gpbetqrtexNDThnZMfEUZGD7dpAdIQt7mu43C1tIfEeKHa
q8Du2NgzEEA02XNRV48iZSFE3LOSTQJuSdx2AHX9hwPwwbW1m7xPZNysT/27
Ym+3PbEP6t0TNOiy55LeKl6jBA/znPGs/j2VvHKjEghjuTnSudXmt3U+iE/e
AmyCrypTujbusf3zhuHd6hL27e4O2mX+d9PzmmBoZAQAYNDGGfV/LZZe4d8/
ZNhTIEGmc3GitVKvk6SYu54yyr8cKbvxMo/ptFbHvNvm+yDbtmZBK8KK3Dyi
zD9D8CYXvecyWB9HMYjz+r5C0mRTcHqhNuNEcgR5aot2uDU76NeJS3+xJkxb
JPMgZOzbKylwSoTaHpZ8Ap8u+mE1GVJp4311NULyE5R/3LBdViNtou099wtY
jceDLH6La4jHhYBVTW2lIqjGwVDCqHZksCjIEqPO938VbdmDmQuujVXNWVoi
TYrVxWyXtNxcYtStrUfFbb3a6KURwtV5v7cNUeMS5OTOLNakv/jmXFPgB5FA
M90SxMnrLEG60vvCNhUag4pCEj3EbNY9aqMRV8KO/1vUKc2gfgd89eKV8QW2
UV9jdOYgYvjBLP8LAW9f+tL75sGz8vu+N+ipZrI3pvnu0dENHdlo+40L1xfD
zCN4TNuUgUSk9JtmDfLX1Ujng/z+G+wTA/KeUVUZ0HS3qEg86uV7PjYY2LnN
qL3ZT0zI8fEBpAmWR3Fz8H8SOxaROlbaSW/d0+hEjKOK+QxlmuNcnDgWiAjl
ZGHOjcvGdE4zKDtxP3gMTzydEbFVf16O/Yq+1BDWCSujR6rYHI0PdO8DWBSi
nSEtsFESTklO9RakIi6os2WHtidc8MhHYwGaDj3uX7eN6esCp8t8LFc4i6/D
4qSLP1U0WHjct5HdALbWsxsIT+/7aqQ0ZmThnCjcrIxKIRTd5t5UZuqKT/iP
XYPd+AI9uRZTjDhKqy8AJwtj71bFFCqNlfaXvtWe0SIZObUnqoovhmc6rkFc
zSIjH5mnmx6qUAPhjas3wlGPTFQLknGdkSAXQu9nbB0cN1zYw5/nAic0Aaey
AyQiqCTvOPXhZfkp5uPQ8OEXbl0tSjh82G5HKZNtfDuQyrlVO4r2C0Kp1ijw
KE5CtCix+rYNQSLafFG+kOsRjjlxBUQq+s0wc+Ux2ps8w7WO8ezS1f/IYhnl
V/FZaLGiIq13uSF/F/ObDa1qwTVR/ZitYchAul9xkfB9vycw9PwUtlnxNYM4
uVRSyYC7fdb+Rm53Wl1zOPxKjQv9vcMnz7mtc9MDaqLJ3qWNMER5RkcCUuoZ
aQqLG2Y9wgA/6BajD7cgxhHfosaMQnxiVhj6g4l5O46iDIhhCc+IhbDC8V8O
sxoe+h/SECZGJAjTVqA+3KMgOocPgdfguhHf/tK6/7a3R2/kdmY1AN7yVYDE
NAalh6wJuYPGC42IHVJy52Bz2l61MqhHRvKsfBJ0R5d1ae8xRnaV48c0e51X
QguIuGh0foImlYTLR49OIRAU4Wppb7j47lwFozirFXgkEszM/buIp3FPYLgT
JWXxamwfsTUHOajuQkSDEF9Vv3kBcOG4CWH7YZQ8Z6tJvBV6eGbRNRMNVVQX
DLTqKJJhEDbnBNhAst1Moxlf6cHzcg5Q8JN0wN+FBf6FWM5cf0Z6aK9vFWe2
o9cUgmrUmuhBrvuZsZRuXxCvIYRM+MgMKoq8/VlpoptJfKYVW4Ku0vsLj3aw
/bBmVUvFLIRzMd3Ka1j5c0LXXBG+Z1xqnhGJnXfe7kv3ij/kK2DAD4iySnvU
ijZ5frZjwuWdwsQEI1t9VRv/b8Ey5R84XdKS4lVrFUJ/XLQkNdh0fZV9dL0A
C+wBOLL5CukAt7C/SjnSAmsTPS2tZ56NMPZ+rWxP2hLSJherff7kF7FWhKaC
im+RNWgCkFKNyUOgvQwyHPiwcgIGrppKCecUC3AuuSn11Um/+xldYEUOfOIJ
JRJHyEqhj2qz+8jpGnz9RJF7SmTh0LXASg0vQOM5LAkiepCjXe8m7lf03EvF
gGxjjuVQE4DOAE0rT8+13sBBj5rGs/2wPNjcu8qikqciMrRMvwpEXUOC2vrQ
Tbu3A97Ws1PWh7jvJZze9riP4NeVfXyC5SEirK342lwhLO+MjsVZxHSI5Yh4
nuB6fFYHNLvUAmEs3EmY5rpXEn1mOmpN2IvvrSbSNy3Mr7Y1JqamrDJoCljr
vR/nf64ajC0+Y8lshbQg/X/P9OyoDtAqDKYQLCDoB7VWBksWOBnWxQHykZA5
fy+aHF5lcvNwWF8I6W9KW38LssTnw4XtWCFj9PfPdfF3/fYM/jsWNeV5x0VS
74RcS9LcBZpILHg2Cvkymb7eo2kshUmZM0OPBT5lBMQulkmGjqeawiNnXc1d
gXZ0PgWpYne1wRjjkxa/hpI82clF3g2Mj8133ryk6QFJ5YRLZBEDoqi+3kwE
z6YyRVXXMbf8WanxxAUCpcny0S1CZtO03Hd5redDKGF3OxDJwBDQQl1nXQFr
xzJy8AYTKdACUMJ/skZHJCouw/Bh3QV15rd8ze2hgvyVPt/4SW2OEedRLAYK
cFIyliEkeSV8pfVPd0BIwtaYv6Ye+ZoPDt7C5rTyLCRBipgUlb9qd2SfUtXA
FMyI5esXLRIzeBwSfNRb8xIHJSBgFY9NEvIuvnh5fH39pE+aEp4OblgHqHnZ
1oqXfderuG63WZ9lNY+XDpjFt/T/E6VRh48uMDAIZqbIRUW+z8bQe7nSanjL
BJRLFDxMfglq3xGJjKPzK5ntaWtxDXimyD5H4kuCPjZTHho3tKFNvKetBmUu
puFdS7L2wBcrfG+VtjL1h6wYMVFo2cGVhb4WTOm0ANR5BFTrEVVsB/BiuV8R
Zeultn40+nk7J2o2f+NqVuO3e6ANkD4u/AgAT0RVL0K1hFfxSAAJm9m1XevG
Ys8dp5EuJYmjZj7bSvVeeIlPzxw5IHiVhx5eJ670Vkx904oTew3BpgTTZcbs
iWM6z6pKw25D5y3d5Pj3+RePh32mqiJgnANvnBeYztLXUneX96OX4Y4rT6GU
8BF76+uxXMKxQ0zilzOb3aZJLxrsUF0z8CsckINWnMlfis5BS7hSq0iczpqA
fqQEGukPRSMNRswS25DEe4ex+Aqd0YavQPfzK/Pd+aS6qikHwKLxe8EoroGe
S3KAKpuMfhWi6mfx+JxlATqvVXPBSBE8uD0kvD7kbmw6j0In8zyAavW84SAM
3uBtzu5kpo/4YGGm/T1OrSN/h+5svi8WuQSE9KDDFb06MKgptGNqnqY73eCr
eZe8+WAG9CaHbIi24H6BGB1CSHu7oRe5XbdvwfhYf2BgYusAUYwDU6PeZKoE
hNd/7rkrRN0GOEjNwlTH5Sgpj+qdSvfqD2EvyYQlomlby6GvtTOBl5ehSIA6
gBo2IgY2/2nC3kckAQCGisfh43Zjaig78pNVkYW1vqkChglXUEosHCszLkk1
W4sF2SNbO0pSFp058iayn5HSHcDNx8LIiWiQyFqmxYjCEAVNy2NFfSLgo7Up
phqj1n4DdDm14wwVNPticpinCqf8VzpUu2HsQDzykDc3BEXOhTx9jrD3KpPd
qbxi/tUGJm0/vU8qQHQbOGsJWPNFTD494uWJwP2b7qyOu3ULUyB0YiWtH/Qf
fA/tU6WtfSOw4yJZ73FA+k+I+BUYu0ozN2qJDbGyn3sUwA/58trHjw5/4d94
ivTrJxphSBS8Y7vY1TmFYFHi0//8MSdt2UXmYSz/217ogDgLF0zLtZuLp40I
E94KPE5NGmqg0ta5WilNIhMoTqyERKAwL5QIEjVuzqhzONd/jlCRGmXWq7M8
5Zc7koJdXXIy7NN2guqPUMPosdk2JpDAZhFnMcQSTKwWRvhjPkztqLTcfm1j
cpQ+QE0lS0M6Pstk5DdlB/Dnp2B5ioH+ANLPVlWrVBrzSC78zv0DzOjQZm3z
/rOftZj71LPxL9sP7wrGcEoRGkUbAq13Yok4IEj1Jwwvqc+WhqcULKXqep6b
aPfblHocqo6FVXy8cdHRmKXgJ7PIVlTQChuwpHNlSCAuBhCX5Z1AaRIDd/dO
NMupubguPBVi1gYhnP8DJ3Y74VniwwNwBWJU9jsvCTCDFYKLPZ3IYmHkCRyX
7HRiK+tL6m6BJ3wwm/BFwE56ZIR2dq4J/bZCo8wZAv46VCt4w373hESqRoMj
0tLOQ0vljGM4PaHCi0CpVqA3PIg/PS2CNHzhQbRVFwV04nsPbd9P+LNGOmyl
nzPP8m288e5kfs3CWgC4pnmJ3ZdIyNKd9aYsqOufhJ9+ZOcQJVfeaiIY8P6G
c9HzLXff8RWnCpYCzLxYtnzLiTKysPztgZTyDA4tB6zq6R8U5t1H9ZE0blX0
tqCxxQgIvQFH1ifOH3XD49KVJy6LF4mYW5NUi7aKvwmiFT4jJbpysORGQDmg
2z/QyZw+revkS6jd98wtEF9OE30yOKfoj73pBVsjbCUvgVMfFNteArE+6vmL
eL11KbZbmqfFcWVhCHnSz9suxTlDKCN2NAIevoAtthm5dQ2SnpoFUv1K34Ji
qYp1vauySLsgOip0XkyrCStpW02LICcGbMzYx6HIgjfMTLdyzDvaU+IaPEwQ
PcVgwNXqp3/nNiv0OrNvnYXwD19cPxvOdCkvVnkCZ6tr9n6hy4NnLzWQF9Y1
KJUoEL5NOVI4U9LlW4xD2hrCh2ygz/Jpr3CH5b9oQrqpPJvR0nn86Tw8GjhB
/AMdQxtD9pltsDCysiBUzwgeTW6K5kHvQQ3hhEJp9FIfEK/A+qP354LgKNDB
Ka65CvZpn9Fjmy93QNoHksbzBBDxmCMXl82BBktoimh1OsLjkDGNcpBJdVoh
JzyL/ClWfK98ha2Zsc6mjLwR3Su2SACkSFe/PnIt6LDvdQGzUAT4ftCOyZM1
FEZIsmrQmzqVFcfB99yGMuGC741aTsn9+KI49uCxHZ/XJVk4gw0v0EZlUQm3
bqv9mVdv38IxBvWVEGs+SLtQY+tohf0e5K8crFTgMjfau/O0TaY7AkTuU1hT
bj5Nreh15X1XEsExK5idvwxeuyJbiOC7wyWotEWZRpxoALf5Sq+HfxF6mSU4
XTqQz15VqZcG5RSYSTJDwXLE5n59Xti/0SrExAbOGfiXgnQemSYoQ1/08OZh
Iqhw9Mdicp3sf/PyXaQMqia5XyIjXdg41hHFP/FSzKOfiHv+J/CLk3MyeGV8
UiTXJZZiLDZqL9XHL/YKQhpeQZzFORjSyFl9YDCO+n6zk+TU/4xnFyFmZ2a/
HBqpm81rhQfxCtjr3wR6Aa+GFa+G+My8VTgY12TYTINYgb8syeLg+hXjE+ou
vwN8f3jIhsSaVhCLS0DsHRVMNc/XkgS2NSFhm1dSVcjK+nFs2O0tpjALtgd8
K5wxSKrC8oZ3aYR4Q1zicCY6q0Xc5FWN52e7EwyEthUZ+kBjzectRNjBRlIx
XBgHMxqb0lDC9f5HGFnKGpIjxBbEfuY3FCbLyJrM+/LDY7IJ1SizYPMRN3Kr
KG3PE7WJn/te/eAqKg+D0jH5gVTy4WxqNXIbKRccOUmKW+z+2anQmpfR/+Ma
zKbk/vjtSidE4+XlHBju2eF2VX8Hs4GE0+GlzXiGR0Wkv+hiIckuyP7jGh8y
dClwN54z+bzQ4vPISE1nhMtCiynTGNSnwLxpZdZG04eogtoJmWkkXec7GrCt
Hni8JBoUMnxfFV9iZh0NG8LwrO0L1deGwnmXnQ8k9fVVvcEu/Ff8xuHfuJU2
Hj3iY0YgQgzbtfJ0iFh44lTqqadUoJGlGzmjHES5DbWYDl+nEv3qfDsy7WW6
ja2EoiJdPLZJlUaEBkHxnu4L/QGWV0ebZG6SE+8EUXDQNti2ARQm/Tq1foD0
riyEyDIx23Wn/vuFKXfM8A9JSHJB/Ci3W6iVWsq5ICn5pIzY4AN668b63AhU
sXw5ZglC6gT155c7taQoLUWwjMVOL+OdReFg6eTP/9AHKPdiwKfiSx3twyxy
g3S1ZEFc0CZ7YyZK6gnNOwEZMBoBSORNtZ5/Bj1DRuzcJ4UxbdG8GTCeqXPJ
rOmtJkpKST4G1AQNjxwkBbUOMqV5APc4RZx2HQTTNP8VqTCaWScaK29LhkAS
i03mjKdxdFxqenp0xn/Naj4rkri+J1SrPIFFxzXpi0ECSArq7+G6zxhWdopS
3rAzBuyBCJJRAn7LDFKIJRW12G6/lEZZMaoRCWVtF5z5FWiFp0SnCNBSYXV4
i/4S+KZHfl5KGkd59jhN6/h377GyGeOw1uWQVw1M5nmGFtKH8ERTIfefMy2A
evDLyZhwMi2Ws5sW6guLkc8g7+m82pt/6kgK05QKbOgJUwt9D9T7FaKKeYhu
z4dWTWqMB7AQdLA7j5y9OiGkLa8jnkTs+/xTLUeM4ICY6TZ4tWGIcoL+FuIP
/YOuSt9B/q1oKK0DubxMQ/w0tNfHm55N1FUbXnr1nx8ou0RcBEV5MnbA3a/D
mR2ffxJsDH2ZicDuF4U7j27y7Wb53Z5JW53Y3i7CF5MIpyN8eOVNZrIowxj9
NIa7/WXWtM8DnEL6E3sHkBEYa5WpaM0OTpPzOo6JvX1hLkmeeOK2tQcHsWOk
jkXDdpuKUZQjMamaES9rGM72Zb8tma9FV9T4VaxNTD0wouovgGeebkCE0fAt
JCA4KCRC7K+wn/gDLmbIpbXDJuKwEhnlW+HusYNdZfJ8IJXcA8SL64sLJ4g/
Ii+TGuMgiw6SropOuI9Vo4lZFf1Orj2DnMly9TqDufZYRH/8gy9urrRGi1ek
KeGhcVHmUm43QBQLRHsCpBDXHhJk+7E0l4rNEESbOLJzoA/KzyzAmNgaMqsI
iaptZPo9gEOdJiIZICpWJENKxMHRhxqxxhvlTRRWmqiE1HOqBDFQKSGh34BX
gTW/5mo0Fy62ObMF3jLEFln5GQK0uzVutwR9sW3ReQWc1QimohTpbHKqH5Mu
t1uOpU9kUz6Qo0BkF/Kgnno1/JY188TtK5POLwzkiBIg11kZnSUh2IsqKQAo
s0klebcMSZcK1DfQGDRtqGGMQTzjXa39k6Kgy6R0/ztv6faEBi4RRNROlZl6
kCKfLvbsrvGs69lHmP6Oj/GUgSDW8+jTJOIAMmM0A3cq5MxcQl4tOgdPZwu2
e/pq+dDcrR+pKiutTl5RrYI5vh+AYW129slK1o1dHpSD6FSID1MuceYzP/Cq
7j88xIq+DtfmpBVqbcHAjJP5+Cnful23gsidFHmGXNqWvHNtLyI7jrC/XsCI
lO6cxlfiEp5YGdH3fpXNCjBielQ2pKEdIXpc/T3Mmgw53UXC+upEvfxDXIPl
2ggBqSwFVKXv2nxihN8Aud3jQpfJzPZr0F3Vv/6SqKte8CtmFn+3N5edo4Rx
U9xtuvCSAwTzOhPGd/RVxSToda9KKXl8VopZLaekOkutyLoylup/psiLtxsR
sGOBPBc9iNCeD3CVx4KQC7d16YhDSUZPF1Ou33kxnFRkYpCKkS8mbbHsanOh
kOUYK3T0x11DdeSzPZO1uARWGpawpqlyRb78RXpDHBXrCR7vKbF5uxcF7/YR
v28pSGFMBIWZJHCPQAHqercDdgkLfKIKASo+EDeDGyQvHp8B7CMNsN2FKo4D
gMl6dgN7HdaElI/Sb0LYbAHhGG/UAQfufTtjVURPck06wVWTZn8atQJrz4Rt
nzbWKvGwPtxthRCSrKTsJ+3Ubcx1g/y3WaQ65cch83WO+3013gHi+BguPLB1
rwDbyNgUT+bcKHBSGaxmj+P1yniQMdRheydz/BjYnyuEEAbJayN1BaWGAyzP
3dnaMcFO73lYs9HOu8/Qx0kfudlgClKI+MssSYgZrE4rteCPJ4d2quJ+1l6D
vEusduW8VcTO6sy7Ba3rsgVzbAggOKJOgPpMaL3j/ecnk9FyDazSB+A34B4A
CNI/rB/mc7vqyLN7JM3qguaLhQgGraAfvoi1qUgLZ4H8+Y72V8YCu8G67ls0
Zzn8Q3+fZqHPTJSGxjA8+WWAmC+DIzXI9Qsu/T0oqdGKElLdCXh4MK2lsBP7
FCxp14TDVMlR+QHYZ0Cf6UQW0/ivxffWPTJVeOgTB2ObrMZdaNiFzNvhKVRN
d64TEAQnmITVMe8EwusJ8Z79YT8amsV+Ro1m5OO0oaEjsyxLJt+9qoLr1HtR
mA+jLCiGtnsrHnkkwtYwcsfWlMAvgTbx2VPxwTMV2fK1+h+/Io+kZAtKtIkc
D819IIH6g/212UB7w+391vC/O5npEqkUY9NDihfKb+pb2+86eGDOH7sXDVt9
AysdZH9Jc3pihyKrXMHykjPlA0ZTJclrk1bbZ76XqGoDlrJnPMMkWt2xXpwj
3KWPPE50xajxH1HNPi0qIisl+89vwlynEvRdbRpgXBvctxakaF1UdfI5AW3o
lFKunKvJUOfV43uytNYBtUPrASPqJz9wuYbDRC+LBqScMbrl4UzfmdD4uiXB
Vaw8uHNLm3sus695uy4ZV+X4s3QH1nZMzZNFWn+EPf+6ixFSVDqEqkEzrIWf
tLf2RThFTP5sizkghXuafCtEEZmrXG9ExeZb4MgKdGlTXcojw7tAh6P7+XzN
jf9GhgN3DzHN+gNRX6TPh1GDIF2UbXBFMNPVqF97VGVuPtro3Xjw61H4aamk
ownCaGLu33yuehWUc5dzPF4mdvix35nKwYLb6BfZbbwP02mdl75dALjAmuXs
8/5fRJf5NkB/Juer3O/xLv6BpXVf5Q+MSuvFEfJahYBitwKFS5SZ9PMdF/Sn
iUPB+yci8+pmlSxOCTR/bZuUPmNNUtcx+kgV8hSe/ICLnEq5g6ZakLriUDyn
FAnWfgqTopTue5kp8yQbWFiOF6/Y/2uSRHn4ixiBrdU0/SH0e8knuuzY3JJK
mFlpsPwIkJBN2LFhoF/rl6vfEyUUzqVICmtuBa9bpMRms9J4EmNyN9odkdJk
QIKqrdkYuizfbU0S1t2Gnviy/h/18PPzHOkqHgkQhOHmZOjvdzdpz3vw8NVj
e4iuivQi2LLCIj+7/TV30+zyEKq/uQUo55lhWUb4DWIKamMhcDIKI+ydD6Qm
TOfHyB9iTnSfkXa1AWIeBEx7TL/4KaBYpQEO7TOVYl5XnotGm+jqRGiayr/9
Zjd4YOMZ79gXeSomucKPQLj8baQsx37BoAABgECEebQW2DZ8jjRC052zQG9K
wx/Ks4Ge5B7DVzSLrB/LqLNsUjPz7JoPC8L2+N50ri0VNL8UlmZ5hBNNQpLY
YBPgduCsLzQpY9MVboDeq1QPfYmS/llY/tpgRPDjelW8Dl7ynynGejrxQILy
94EA8fPH14Vp+H9PmrOtkvFELegzS1u8OG5oo4SrJzkuhtwJMhFDm6TtiODq
h1LIsH8cwUVa4u6+ZuHK+uLOZM9lomn7R59N/gyyRwFJWc3RjrB0bSuQ0hza
kySeCsodqRYcgxiV3YB3Ol5BmWToXKe/Kjwi5+bm3hifwkEUo0eXOni4yT/g
GsWsquOXtM80nGQi5Ihx8n2dRtqUnQYOaRCXN9nMUc5p3qDY/nbkOXhT7G4m
vBYTyg4h5sBkiQtzXdcoHP98k5kOkTDWHzeh8ncfNhbfnVttzihvn0jxeGYv
x8MPmvDW+0WIT2hTSOt/pkgQw9NyqKD3VN94pJeGlt3OHWUr6Ajn7HiZbAHc
AtPfEjQGRTc72bjoV9mftUHyK7S5yPaLdlF5ynAbn8ujLubRZqFvfJe6Iscb
9diX4pdjOL2hfloIwZz7CTOh3Dbh9rKxvBDuklLuQJ2/4LtI5kCXn2apKfwL
ccTbYFsxdTb6QkyQmUKPtYKKKgG6hPae4pDsL9hkqfg/Z9r9wBNJIQUrEoqR
vVmMOMxsK+tZT7agK/8tb27HjRrGgo6dujBn0X9ggVWTTiy380uooyQK1AP1
R47VOemAH5PUfbYz3RL/r1VIviBtpDEIjSKZB1hIrCm4ODc9NQb0iS5oyARp
Na8mY5zsWmu07BOM/4zCt2whrJMWe2osK+o8oG8ONADDfaYO4IUCRp7vOKu+
zL2hzomrPBfo2XHqcGx22HGrtvAhuYG0S7i37Nebad5flsnWzNfTVpikVZjw
3J8EJnOL8dgjXEpfqeUuBwVIQQICx6Y56QW96MjMbcCA6bVjNoTc8AXBICkX
81udgzmevIMRadldh1unC6ZSJsowhORV6kIyp6e/NMZk9P9UBwJqwUeUprgu
RkInUm6WZWUjQK0IS5W0kvv3swXUT5J2F/1OVE7nJDuVoBSFLJTHXyspjmJy
qFCv9xzH0G1IratZagQNmVVGsFjz268DYd6v0KdiEd6y9SrAlg9eqY2szYnG
TnNGh/fyvaq45ccNOnqU3c0woX9AzMKcbvsVjktbH2QjO6t4377mV2XPShmL
7IC+M8ZAZQei9npZYP3kWYlJxiT+JeEhmpsVG0skyq+97St4GQU43Cs7fM3/
NlLGE8Qd28BhYTNlrHWEpqViQfejOKJtOZqohb9p1SgQn020BRIYDlz9Ti/H
G7a6IxNPBthP4jH5uNWjmoPtxpZSPk4yIzd93G8jc0khybguAkDF5eXmjzNV
W+0GuwzOgJOC+CbSVoOr2JGsLJKjvzIfPC1Afm7f+pNDH1UTrif074BqoU52
8Ds5U+IUpeafUPIpPkmtoEIKZPwm86+wf/OLdxC7my1otn4ZsRRP/jyUCGyR
15KRMx0gmQVbL3XGHg7GUVgsu5z5Y9ZNXMRFv2Ml1H75tFf2B4Uej1K0/bJF
70z6JwozMTtvu2x5cRugvnEjMcJH1PkT9+hMZoRCi5b64OeFvsJe4PMz6W+J
BBUk/mG3ZwqMvbj++G9eq0VCiTrRhArmalRSmfhDv/hTSukUw4O4PUpqrxuK
Z+R1BOCo4lH7tOdk2kIF81qYwJVlw1XnGpPjJcaeFvTNPXfduWdYL1fzPDe0
uRLpzqX0nUajQLOiTyUtJ/yvjD6vlMw/mat7HbUyoxXUgv2Pb9kZu0aI8E/H
A8LzujUS4uI7yQfE33LFHdN/QWqZyDdUQ8fUiPKcfJTSlxkQGI7CKQkMwYrC
BefsYKxqQ2IGA9IVtxhskV607ZwcNTS0cLFvCVVISUrY9gH/olMc32Jr+cCe
ktJ3riyl+eFNdLeMN4/CrjUWKaoUwFl1FRIRZr0FBzc0DUlRF39P7w3FS/ur
xg+/4yX56uZ6dEeJimIgXJDkMTk0Hr+cDDnCZm9rxC6KhBP9mUTjxOBYLi9n
/k9Idlro2FM+kdQpbZVlU5PYN+1iVSgVlWPNeFfGvViFhZq2ZaElu0ayb2VS
fmWxjpNKbglXngUs2v6GcrBAV9sC27bqRT9+AS6lAghnNEs3gkLSIVUUpjkQ
khgTICnFT+PsKzUQ0PfC4afQd8895aRWEXhhhgVCSeo2xrMEX0zb+hJPe1RF
nbvdfVt0LKWAZ+4o1Nn+T7AfsVoCj4OHJcSTT46OrS4LExa8rHfLn9U9ybQV
ROoYdYZ0e++WktkncPR9rZx0wh0/AZN66hQAD6se0h7Gtn+2+WZj0OupagvF
17HWxhizGm5rvhwUrs898UYJIuMiFGSa3Z6AaCPOisQVFHgHhZrcVHzbPEkT
W4IB6ZsjTMt/a7lljkJCbcwV5V5fALklPXgDd/1k34v1gBXsbW6b+NM/bOGG
Ss/k0npowEcx5cM2JHguoJk1AJDLuWKv32Lz7Xi64cvii8CwVf/6fKK6Oy87
bAyzxcRqpQo9mF8C91kJboDIcHuDYjWXYBG7+dsRPTpRNcYjWYTXhcfDuhUH
QdYRCu1uoiHeUkqd1AGiP55aXarHQEL32el29QeMfiy+mlGAGeU+xxqeHWDM
BgFAOivooYrN27J54qpqXkwA6CnNWHbniajnJ/HyPhRvR1Fx20SlZlgFtrmG
54cNCfQBidyvBLKNwJu8spJmcECq7w2ukFmiHSzowedozDCmuU6IkQBi5Bcd
9TyYlnbehA0L/dJYSY3C7k6EyAVl+673zzd5gkyautIXN7RUFlASW4qAsd/v
duZYdHbcg3lIwmLDNhXhaxRzfSqq4266z8SifW/YvdkHI6apycwDZSsx4P/m
pXMXoeWW5QaqkIa7Jum9cGYit1Bk1WgbTfCxQb8ccDMsGawwhHYu6mF0wROZ
oGhJxigwSNHNIuFUtWuZwPajz6KXCFb/UAfEJ2ngG3NrRLMjyMH+ScHRc0lF
i+hqHtNCfTk4wGgjV4ChqVT1vKP7V6K7rjEFBhQD4wMjEVxGv/W6qSzsnm6g
deVuO6d/GsbuZrNJ0RXc+TzNCsLNx5s3q94B+aJerFPeT9gJOBB0WU0Wt+xj
RmjCAMXcgTIideipfEDBKViOH/LNnW0zGZHr+xeAOwFOtFlhNLsTSRG+qOQb
SRSn8Kpg9X6CEd7X+uSy+C5gWQaZFjLZteNhl2rb/dkr8xXNz5Q9BKnMO9/E
fRwfaYrDD/9Zil6veulKrJlysZz3c1RihGaPgexJJUONsk8xyVBhFrusGywM
XH9QdCxU9+cOpnlOZENv/97RHIMW4OHR6C2V4RKTsOldCJrhMNepGNadVl3Z
MKBJ7Ln/Io7RPbJgYMPQq49a84igIHM/REzpdiDWD9FQKP2HhBlMwYlUVSpn
8uRD9yQX3skiQmLBZo6itgYSy7Pw8Tl/YGkchI6a6NRAoyPcDx9z+z8GYVTy
+CoW+TMeZRANh3cQnTlVEBR+o7jtAD6tvy/NrIPBCSCLm/t0eFpc0604PcD1
MpaUJRt8Cd3/bnfMojKpY1LKqFfb+DCSurSvdHt0oq3iO6j8QKoVBOLQWuhL
I9S+6loPCsSaTLan4SSZh5mNoqBbHv/90IijxLeejIUKGiF513c7msBXJo4M
VwEteTxagc/uWMQLQzJeA9R6q7aGg3QC0GTOb4537ag9fuHE7nwMJ0IMOMWP
FCgLJiI9LnkhfIqBHI0iIPNzAbyPV8svJloshB0AaK+lebpTgDZZSXkTVDKr
sjuNasApsqUgRGH9biCiLJLL+19uxtfMUyW/IxfntVvSlyxcLj8M/vdlsDnN
iqKLJAGIQxs2b8yQK6oWUPtPpGZtxJoxl8YKculObUHiKk6t7Pxj+XarCrmL
Td8FiJ3o255RGdMdHQJg3q5hjLs3mOKIIr2n2bZgn6Lnv3F0CtBU2RC71Vbl
2rE32m+nkZ7p5RQ2KakDPpdXd2qK09c5wNaOiDN7i3Vk7ofK4FhWn+soQmsj
lJBW1LlA27AFQv7nP05tdN3RCeNNgkCm0RxICn9/FRd87mQdqel3h3rS2wWX
7tu0274nwhHdrdwbMa/YsyXocs9ydHDn5R+awH90bUviUYjQYBTvy4UXU1RH
nDfwWqVjPZc2yTE6kwaVbPuIXD3B4v0XrY80su4ePoxeNUAIGoADO93KryoD
OX+qCi5ZXwDB6LrVaYfnpJvnhsQu8ruBhYjmxnA6ZdRwV6Gj4+nxQWOj25JD
veTQWKCnQxv+H0uerIh745JrlzVij4mt0Xs8jY03YwJsx3I7xxKstoYwWqsH
vDpVECDqGHAUpWvIUToMvNtAkS5He79gBihav/ltQ4+ELvEIgLbIkMtr7kZ2
bAkDfvggAoKoio9RN/VMdtXLazpAeAdFT8QEW9ztaYRfgecYN9ba4GWTuJM1
jJA6+StUR2e3HFmridlNX4EN5U+Tm+AO8MrKMALHIRXNLoJ1MYi8/WqYkdbH
FYNCQvHXOgMSU0irDEkjwbzwi4IHOfkc2b5Y/ASpxyrEyE6EmKqRd00NYL3+
/UVLCaX44FH24saVc8cYTqNOXcmvPmS3VYDoXZG6r1By8RVXoYLsYB4drNLb
uLp+ING3MlHM43hlFZWC/XeON+gbSIIUXdGQunG2EYTQkNtqGp4iKNFoJ9VY
DjzWW0hQ8QM1upF+ek6fR/I9dzw6u1wUfDA7b3VL9wvpg6OnxLcBQBNITXXO
fEXrBFgptsn9oe+ANXytGSHrDXPmzZQFJ/OgUwjLRR8KuGtEtEyip7UreZWb
MPvz34Qof5rSDBrvMFE2SyYKVtGqQCQTnd8tIM5cvI9TgNfiTJ/yB1yIAa7S
SEl1JG6whlpWZFiE+Nc7/YJFb5xBv3C/E0NMBi6g1L8EAE43UUnsa2l5Lb46
BwLroeFlYE0mXulFFE/EuS46RpJxrfVM2ZdjtxMaZhFjhGKrVuLfjsKALtq1
Npgjl57W8TAlSOdGzamJVXjiuy2/g4+20RX/01WPh0WpT8AQa6CB45dSAWKy
Cc3U8/Cd/YZHPhi+bcQ+jD8E0UcHE5SB6kuSLkO67h64Yd50suGRcV0ZWOVi
YhzPQAzIFI5RHV2bRCdCXWE6Yk11hOeIrhanGqZZbRKjKJEm2cSGGAzo1QXp
cfvvP/5ZIk/sERy7Y1/0tIS+xdY4hwiGBTf69H3LgEWW8NVmgBRIYxTm83Zj
Y8KWxDCgEsnvOLmQYKYmz818FN7TZxeUGC86v18WggEK0xB1FxpFh2R7BLAH
DTHrNkwAHrbCovZWdfbZbcO4IkhDd4pd3yB10AqGJgxcGdnE0MRlbfcWpDZS
MYBgZTuEQGi/RuevXv/7rrHoTdDvqHPobru3QQii2qmyIOfmCw7Y9yTH9CgU
kFS5LgOOaHxJx9udrWMvBNUVw8O1heN/QjAgPiQg0lf3ap18CivPnZzCzsNI
Bx9ezF5goItXgOwm5dhSLgWZWYHxPdyQTlmshJNX90Kd2uXx7aEdtiOgF9/X
rwIshdalvW6lFu1OGnH/+21ioysOS3khl/mRZz5/erC3dvdW/lMQ+SKhNhuS
calGqmiNSBXeZAcLSOi0q3Zr1rtStkIluyH3svw06FKu6gnfw85dWR4kBsbh
vveyA3CDS7dtngYEfs9PLf1k9Z0fVyJWYXY8GDDihAJH/aQdMh1e2sa+nJzf
DNaRyyfPbS1GwFAmncOgeDx+hvH+E62E7poFHv+d0abys+GuI/ydzqbAw7rd
l21G5BRAg3p/dRdo3GKfzla6hpZXD3vR7WO/GP2tZ5bYHiBdDqnF4GPU5blq
SgKo7LQ/RN10VEzE9LRkRixNL+unlWFt3jQaldJ+hrIt5vxpGk8G2igopZhz
5eCZc/9b4CYRX/EvYwBY6JyY/gar5KbqxJBbzao6ndY3du94u59l+n52W0t6
KizkonvWSwHduoAJ7pPsGfqNssIjMQwRqFh5ekRZEKq/6Upc7AMD/aZj8r6L
oJS2iY0Mdham8KFW2k0zGUWLTHFiXNAv2O3KqL5vlKVvlZHkmeQpg8qrjq1C
BFtFSZve6fwBf72OLp54h2oaTnmvb1ofG0mICbY5tky0oXBPdvWHLI2noszq
KRTOcIsQCIqeFZpzzgd0FTZO+lmWglzi2zY+Gz/jrZNxSPZKefFzlhHXcyKm
7PRGJzbxxfMgsFjgnIKz9P5LNYtjOWEKToLLxrjnN9Sjw2XId+v7pJpjfeb2
XPmKtlh+xJetwRU6x/fCWWOB4ZrwWbmWq8KVwMzYrWibNSnh6Pa5astlK2bd
qYzHGf0ipUDmoxjQ7ItrsmU0XiO9hvDr954+2Sgj+Wbu2RMNStoHqTbKjL4m
AO7hcGT3oFB/lSDHzvPa3ZWPPR2EtMUWKw30vYmLTAi9DbrP8KDh452IXoXG
bSUYzA7gS/+Gu0k4rHszJLX2MfOywptTmfXjyc4cVby4MNhI6c69wXqeVsNG
hDFWQQYMICXFrYovDq8WK5HaeaOjGcVdNaP5HK7gGzRO5CKBFdCSV2V8kuyo
dntF49818YjVAvsZZk5sXAau16XP3FShVjllaUS9xhkPVIGhNSpTVS4ykEU0
OASt9asZvhiVbWd/XvFDJ+LYWDlofxipASLiX1lG1QyjAA9ovn/sSv4dcUB2
+VJ0i/jnrbHNX+f3qZTjQNTH8PwwY49K3KN5+9KowT7z/Baa4u3WxMeQWkoB
hyS2YiYXtAGNEMyXaBkEBbsrtn7Uuth+7PfbKO1oA/jhPrUWynsNYZTQytaM
Gqy9VMnSh7ND+Fl6RorL7ygBh0tlJNYUapflgr6VooG0P4SANXGIDUUJUG7i
PqYVYXdyxBaUZ4Ud0d3jhrG8lAbBMNK5O8eLStUqHgYQtMUQsPyw3gS8Xzcm
lpgFDYHODMwWquqR4NoyX8ZR6/XYO0BqdUL5x2qquXk1DDhbQzDyIiNl5oYY
ZAtBwlzKgRZ03Meh1UwT7wS8Khz9fxP81f8mHicLz6Ax7gDnAiq4q867vTP2
TgBtWiu4ouIZfPgUyRGzpPoIzXDLJqJkQPGbyICE7FzazyG2XEtfG1/keOZL
y3fkPvjpfZ8+DUi9eihr9hgjsCUE1ycghY5gcYHnE0TBV4DaYjakiu40Me/c
IdUaOUh3sMAUDohyk+qKYc1G/eK7ESmG7rNJwH53Xa8dqpxTO4CnuRZsOBQP
C/0CylBP1EFNPnmpX7xD/ciSlkchG9MeT67Dc6/C6o/kO0MILGPlO3uUTdHl
wrOuuvu1ca5IK15jfvKTAcG+PSQ3J1uOw+/Jf8sKWSFyNqRpl01+hdIqHWCz
SD7uUvhvLrWWbPYxIFVAycTpSqKj4IVygubcVEBx3aSF3ktMVNPDWB8MApbS
E+6Nek76V9cXYwfytQmpkopD9KUFJbm+VCx+8QtTWHUz2EEixGEA8HnSNCCT
o1eY+2/NBCsXEtKdJOi3rti5QCTLYVMOo1K7iTm7/XwFSdaMk3M2YYgiOWjG
F1lH5zltFZqqK5A951Hhp41j5uN3c6Yvaxf2D/bTQfKBlP07genK5+staw3I
x3S44eHx45tXhI6yBi6QBbyH3CEHZiFFGZREcGRvvoiOLrBRcWOwTtddWzb3
3UZlo4B64dXQAfDVJYoGRvrZ30L8ceWiprVMDCGo/w0tEQ9h9q43yZsn1TfM
UFquUzmRn37eVvibFZDmaMU8HwjxnnbWvJJ31bz2ba7JHIxIIVCqs/MlhFnd
3J+QMytQlJpVdn1dk39Zfdf6yuc91VW/wO46RNlkc0ZVYGtGNYQud++LbFfR
Mhicrrvd4jB3D8ZeTYmvEPUxN1vDVomPb0yf4YZP9QijhVZiqlHkXHpugeix
nSsTs/McoErAITYbLBMsJEBA4vwZrp5zpTKRx7Lc3NV4P/eet4k/+D/5lCZ5
UUvs2IkLBVqjkF2eAfDRH/SovV2vO68yRhJYTl/07la8nEGlIE/afzhDsJnd
vQ33UE3z7lJ05xRr4gUddg3F9b6to0nujwTFZRNwoUnvsvQCc98NNjOUgQX4
MG0ncS4i+4Ya0thCFnU0uwNB+smII2kqi+E4pd4oOcy2mG67iwtthSjSVmxV
AMkrf7KSj550IK5oqL8nt6dVVf3vzVlCXa8f50J14wPN6Tp91/FC0kcfSaVq
qipxaSt91CdbZ9aDamnfM6azXaD+/DVkpJu1wCOFwdCdupcZgiFxeURiYmiL
TY4mRKqNOYURAKqpDCc/K1MzXfXyzpLckok+jOt2KgtDzdb5NEjRpz95GgQV
4ddzNHC3DJkg98J4CpDVVvf/NwK0xLbybJTpmxjReKvXqkhMG3iARhKHythT
jCDSBHJM2AiBjj37Bj0u2EEmyEPBQxSuYTn8oa7zRahCjut4280bmSVFTzv5
5omENyv7g8jyyu//h8loJcdZT1KlWtg+l1qMquxsV0cDSPCdnREOx+jim+FO
+8zHUCrVqLvI+rxwlyAg8Ptsw+jPIUyN0mgUiu+D7+1VoB8oAGtjgu1gsqcw
Hf1t6tpZiR4yT/LltOJ17V7UyMdn03c+adRQnRDjqn1s09bJWiKxYYXYRKnR
AnSo1CvK+0jBOVZF0V664XxtmUtLjkCJcy760J79ZYH3BAEnVKS8XRTmvGHK
NgjQGZcnhWqOrOx5uvoUNR3JcixisyA2Eq8/vhve9M3BtbJFQB1O5XoJJ4JB
OGoxITMsPnLOLqoHeTJ4NpUMIjKDTTyG44YlqgYkUZf/6KDp0FKqKdJ+nLW3
usbIYdmS9F02mz+gOF/HF/HvggwKJo2nHKtPWcN39JYzUrOTmfOhhZav+ZWc
k+axVdVXpAoyGll0jfjV+J0sHYMEDkEFoQHspLUCNgfqqh7SN697MM2jPPBK
EF4jfCZUMr56UnqMySFNiuLXXYCToTA5Pg6l2KGkBXAEQ/H9QENiEwh4ISJc
dnzHWq6csL1A84zvK/gla2seZ9OIfWzMstwFj+R0734g+LvuV6ByHn7uH4Td
47yq9m6x3ph9bpkXZrBCbx6sPRvsH4y24snAJzVHP1tcY6u5Ms3m8u23oo4Z
YOpgWqJMgfIAor7Kx5ZTNpXdbG6jNNgFy9pxyI5ERyimvP6HAM2737MOHSJ+
TuxbjisEccb6RAy58GPpLtZPSXJzPGC//+8ZY37nbYC/lYxyFOgnJ7PFBBaA
gvcL5ZVEGmtgFa/quSF7u5JDA8Xf2TgqZOfLLsmpU9s0ETRVJ7oiZXSsT39u
GyqjsaOS+VUClU3dsz4Ezos4sUQyZAiZlo8nrlsbe5Ez+wXUUYj/jyvzPqXx
YIflsSd43TBYBP24vgb7tHFKmDlhNe2R4To+2xD+qG99uz4ARZR6t0zHeuHa
SWJU568jVQjqGcDyCUgg1qEOIuu3KrQq1zdXXok7vuao95zCYK5AAfdNvVyi
GV3SQFi7YCKX0lAKOuOxKHWtGL6QIYIsB9AqMXlfOlvdrgzHlt0nZBdxvBoL
5eNZalZCjIqaT2dPM6Uga1Xaqycu2Ojc8/DpkFxRFOCldK5gvYYKCCRxtzRG
ZsrmkNLEV+sS2Gf24g94SeeXk26WtNQXt+90XLG4HWnYXhW+TihNXOssNeUJ
T+6tNxueiGVcDeDA4+ndMOuTZXRCv6juLzc3k+00ae4yUZ63Tlt3Kpjc/GNc
KtQDKHYuwfHcwZJ1xFUZDBTN4BIUnCVDczW2pc0nnJINTJPlrBxdE8lLNK0j
976tOwAg9KB7kcFGBRWcHRGIqwN+IESJSqgsJnnpDLHkYwGaopU7b4G5rmoI
5zXAgLal8zUGVjO4xCwJxF/Oh8s+VgjBtvWg3TIt9W1YoVsIuWZDKvG8B5we
nSE8VwXycOEyUZ93Pw9i/NBOx0M3xzoFbtC0LD75gOmUybBMkip5V/djxd2X
DAVSpmMRxWVjFQprfhlhxz4uHWpuaUpH1wILVwIORgbR/tw9t/W1hi1KHswG
K8q6uo5fSFqCgbxCbtKD5ku+sKMSigGQwJhWK4oy9WE0jZkBzoGoPPez/qc+
KQkvi8b0O1dTf1UduGSBzzJumbDnZb7bWMRJyvBUNJSm92ytev+umoPQ3Efg
p2krrcwWFJiLstZhpV/pDpe1ctKjgHoaxoVT06wA593RD9/0x71LqN5qCkwi
PV0r6AKJ9l4bVZXevcW5fp9mXxAmGToRKxbaqWH8se+QDXEVl31iTtmW4Tnj
Y9B4CLStsekBNtsTfSWjmUoRrkKoxYCi6BVetzEzcRlLf+fRhCTbg4vpeu2C
HOv4J+53RuBlwv6Cug4J3P6cbDVl0/fwgHVWaCStTkMgocxyd2JIYJXkxToE
KR1IPw7s7LDgxo75bmaXjjkfUnB2N1auUSmQdi60Dxd3MDA42iwZKlVccQcA
qG/jkAHl/jlLomP1J4iP6lYFbJp05Aezn14Ey/3Y8XgxAQPWMGXx+6ctcOUz
ucelDpd/jmsT/IlFK+wDIxTA5K8t3/0pHQpTLIVanpC9NJ0gp741rFuE47r6
Yop6SXfEOsg+Wup/g5sbuFuI70M5fG7CZuOB9l/0UZuUW099qMX0DsftYUno
ENYy1OqEaYLk7+cOSt7uWbmNK+AEm7gTajvEZxpq7mTs+Ikf+z91hIVBH0yX
+r3VDv5UdRPKmF/0TRtlK5kdL2QjlK+TqLfjLdeE+/jUsPT2RDgxTvyurTrr
xog1GgCQsCjISg/2bC99l95KQcr2U2iqOgPkWaUINujuuiRmAFqlGGrIE79C
ZVODV4v74shKTfhaFjd/aAWaqms8EEESPQy8y32Dr0l4upJIk3dX0GnA9h7T
utApzeOBg0uz4Q4HE7CnhNNH00VUuUWRt5i6uesN+j7m92+K72bg/AXOK7xw
kODIfD245YoVDjINLNUVU2VERnS2HMr4Sbe/H1sbeFmgHkJQCTE2dPYFqPD3
ZitRZqIVwJEw99+NnXV8TV1zIeaO8+cGxUj1RsxJc2LWop0v55VqBHDn9/0G
aTC2YKdl55LgkfsN870yX5DUy3wposKwwV92c5UauGARUZ5zDDTtldR27f8+
pc77ulS77pEiRJoG1zuBvbcS1JFQlqmidisl7i80tdSqmnbK221c4JUspFpV
HQueFL3KOTyRcexC3CuCIxQcygQo8F9NbsR0IbDdT2U72owNcpOpESwevL32
Gh7nL7H39N9ym190mVOuSkZadtIPMzMtlb7QjFAFZ6rX1xiLHRR2K96OaPzB
A/ictwuSOIIDuPOH5OPgoNeKKzCfBKpwliaXMyYfU+5xttXXtgI3jo6b4Z4A
xni5RDCCph3PA/KSNhq08BZ1eMNXETpyD/qFBsOuKdYFGqiO6SBFdOpJ2UQ0
WqiUwUK+AaP0529zLo8U1EltVG7sy1JX9P5V/qIL2VanwzJCfoKpRf+bwefZ
MHzj9KGoRa+sfVDaxB6RAilVpQLPDLoAYZ/Qtmz8mAa5OyQ1+47Kh68TeAv9
VY5bSF2P+xnqC2R9F4DAskegFz+jQQK9cs6ufNfgT5j7W8dE/qa4p6VzEpnD
PX5sxqi5TB0IRIhcv72lxt/GZVeTFlg1EzGTuu/bvLKnk4r9rOd0WKHNrHwx
Isokqoo56jo3fQMHxvNFKdBYsRHd35NsEND4fgrU2M92bgTFNzhPw+o9pSri
OLOszdIUgK3N7NcAm6EW8aQFwf2bN0gK3Z4Mk7EYc5w1iE/Vcg09f9Nw5C7G
R4+VmcwhYwK+QDmnfKxgEGBXSqKmLeiI1q1EW0gDmmrj//Iv0WLUvCoRERLB
q8uKYiv/E9bLhdbMSbN98cEcAloLQr+es2QNlRXWX70jptkR93kiNMTHXgdH
A1lppgG5NDOAp9NSzIay+r6E4QKawZZLaYQkyO4q2K4wUnl5yti3GcdDON2z
4T3rdxNbhOWQmkwtrIMvUSqmCR5Qt/AzIe0Zy3A2OFCudzhyiqYvLBpF15nj
Bgt4TaAaJxznBAas1Ef6DZDVLNEidId6ziBo67h7+8MEm0hrwGFCYdXqP3R7
VBVqzdyfXtNh/+Z6SxnlhSid6zbsvKHeZt491nl/uRB68M/lSQTGTlVfloih
TIz/Qw6V6flaqLKf3zBGfohEPFRQjYglclOR8LAud57X9A/c05UDvWVJu9Ud
PMR2h1tX1KrjRe0XRuwOUe0nr4rrl0yeZ6L+hwNQ+sHi0lSIz5obJH3f04qt
y0lH0/YE055LHtkbT/N7PrJX9HkaIMTGgruzmkw/ECRoCbylXg7UA+QqKgKX
Q7e1CvytW6T3fRkKC45bMuWPA4K/71bywf3K2sfelpnijBMBXKYW2cU5gze4
Go+LG05if5IsfE9lI3uh2JbHM3OUdx5HurfrPtDCZ7zjpxDEAJhZhq6A0GzZ
TlmF0RDEe6b/cQXyZv+xp8p6nnnUR5lrHfUso6RC+9Hs3cGXC78QNx7qf23k
zlJCA5Rv80wNVd2g0VIdm0hw5xG/U3Pik26ayYep2UN/bAf+9IppaiKlIYFc
11OJRwTJBB3GZr2Q2mR2YmSTg+6KwkKVJPubKlK3ZVgedYcYWa3IxPzSq6bH
dNF+hkzcheKlmLg9S+V5MQpoS6jVaVMr2H3RnxRX6o+aynieBiImbTLGhcAb
hFsap76KCIYmF5S98MxLerlkaxNKxtWGIr1+0sIKef94n69ZIQCg1hvPdLtH
DRIvgPFJhrtOwn1BQw2peA6TbLE81OziSjO+zDGXv1pXHZLC3HsQKFzdXvvF
bSBdZPsIyAFRe+6uuuOlXbkmVT/OmaAH2GKGwoaUzYnanefCh6vNfF2/e8g5
wBWKimmzQWCbH4StJXF7S5SAK+DDFW+fWN62PMmcVzxf7W49mdC2diudlcJ8
ki3z/Kfga1pY892FtGUIgRIfx7gOWbtkuIv82vN66D3LKha6pr4wnCbbIRHq
v4dcR8c21E4r9p8TMT3lhQAWFwiXaprgAUitYDULyhDR+h0DoTkJpcjUyLsQ
EQCGzF763+8ruq47gD2te7+8xGTiZNYveyqIMo9/ZcQiaMro1ztJrmmSGwMO
C9vPm4F2JA4+WToEx33tVNSbOTWse1jV1/PmTAYHunyy7rTJlzmKEjFe+Rac
VtZZg7tNx73OLH4QLMMzRucNUXPrgMy3HSiSUI5M8ktx+85EzfqUnMRFhVSW
bZvvQrgwA+t0geViTm5/OMA1rZOV3kPAlfJQKl3PIs6XqNDPk2SSgl0x9Ih1
E3yXGMunenCtNKW4kJWKrT30gTOdR2d6ob9jIcIDzFedtvYBlabVWSe+CSvF
op9p3UXW09J9LU9sPcMIwVioTT0A0DayYTEaoAd9RNe850cXrVWSdKkC8F21
f/KmpgD/n4svcpIqoNtEuxTZEm6uCcD5w68kJuXpPgZ/a16HW7gWfTJydIrx
xAC1gfiQlp7uey+NGzpu8C+UBODPtBhFR1sz9p3/aGI4DvebXKqa2rdhtXjd
jGNu4aKYXZPeSv8HFFtIChQrN+Tvq0STg+JRJ1RE5vTplQThuFI9zJQh7164
JouWzs9u4RbjYkdjC7aaTFLZRLxRhgHHAxnC97gGdFyKlcT5fGAO4NAWHjsZ
daDhBezchDWmUHRyaa1O9xjBviM80c5bM/fChM78c216+PT/oo8X44T8hMu7
p8TBNjjRzwhgykPrnV/eIz1QlcfEvmXOV9GSS9syH3jDPYo/Me3HWvGN2PzS
wKnDmvRM99y2al7Kb7coBmT+Ls77n9pcM8tJk5U328lfeSR4lC5omaw6P+h0
+VTEsmz1YwJdhm4YFB5BMvOYaQ8s/2XViL8a/3rZmwPIHxo/Vdp1PV2+dnz0
5r5PviOrehj+BO2pJSpRUjr5mkf4jM5Kp/5RoX4AagKQRhtLTFVdWjd6cn8A
2VSfQBZudEHPju5WRN5BAgpFaqy7b5DVDvrlnajb5IZ/HkrnTf8jbvdgQfOv
LZEb9F7T7zogeT9hZd1jUSz/OIR0RbXngOtYizDu4e0j8e0lBUugud25Jt39
dn9cHatpQVg+unqadsFXHK7j/tuleiF/8mVhwK4mttUN7hv1RuGL/4pVjP1k
DRGTHjNy42f5/BNymJGd0YWFti5LebFYQDE+jouocvfQUTt81uHvHC+5MJ8v
7/4RjckD0LSDr3OwQE12pKlPDWvO9YpoVd9g6ZOBvxsELEvI+rJSD2BNlejT
muiwvAodSis4lgf1oqjtO2DMk0myx4fV2IaE1OyZG5c86mMOO/DBEQF+3cAe
yp6H0qjVCFUB3qytiu8pgUiNQbNoEw54anQnXyyriPEX5CTi+t9IG1Qb513L
nq9CZ7SstPSEDJmUcV8kCf8D2IW8rJtxi7pTsJYoLoofi+M08GfwvoR99Z/K
EQZsO7/S7aavY8eI0buAQWi7+M+m5myEKWwnbosTv93Ls8s5OsDFIMxv76E4
kZNpuzs/9Oe3I01A9aG9a2nCofsp62rNhOoP7tTgwxtvwp+iA4vDPoW6DcMW
VB61Lkgos/jRqOhBIdfZAyGQZU9zJkx1qD3wn9DmF7siwC9m0cPH+Yipgclk
bG20Rt0DnRoGCfbO1Rlz0IxLcmwCuXeHwQT+rce9GmxUVZkRSTaz//hjQnbr
u4a5BMkvf9e5b96+T9LOOxHb6gIfwwjuv3z1dsBbXMLwEXBGEWnk/cN6rSNE
C0pQvAayMdUPu7Q8z/jxh7lO3P6wEd7h+KTB8ZnQqbAPTLdnOr73tdrzETlL
5ymSZ9TFEx4kIE7WFFKpG6amyta0HpZFGRq7RoJJSfW9t51X9VkpCFZFip+6
GRyNi7SK5FXtwRrywccEa4sHvFWRgCVpbnPgr9aPXPWIaop4VqcFG9t+r9Ju
5S/sNwoYw47r8xgR37s6xNscm25Mnpj3mRU+AiNJW1XR6OrAA+zQmbBhS55j
LlU/Aa5yszp5gpeszvNvxTfwr9Cvl8ko0IP9tNj7f8mKqgSqfevmBcjmn5g+
Qjha5HdPDyvKCnIfbT8dEifcRKVVa7kLSYsCiOANIakKB4YQ7M1NzaqF4rh8
NpQok1bT/ydXwIYVyAlQSBZRidYW0RM8AmC8244TcwvWM+C/YaSliEvRCfFr
To/TO/zCIKzdHoQWl6VpfHwnbmmDFTgf5pXcuKhsqezc24XyxyojyqYz/HLI
Mxkb2cKM5pr4QUVuShnhteDZ1iT+ivTNFrFh8fP0/U4rEGL+H3lt9+oordgN
JkyyuY596tGK2Mb8gTo1W3YLkYxXzOFB5M6Un7qxo8VWTFKaYhQIXYSu7ugT
LQno4ny1mWDHvmVeGO9jsL9Yb36q0n6oF1t1mTJCJB7Ajh+yw9/ISnCrhk0i
JA3JPENf3vHA9uwJTmoiIvEXZ5KGh0Lhwtv/Vcr/4zK7x4mG1yHlfPolWo2j
uJTJ1jWx2hbdYWmgsj6T4HyodhPOgUbDTd3QwSU8SHQHUG3FqEcByMFd6Aw8
kcpU4/A1hc7AotyF02eTXSlvvPdF2qjtJnJPlb8s9aJb0aquIG9ZuGQRxa2Q
ep3aDqafCxai8qZrz36Pm2pMuR68+Any2Pkd0+zxQgFouDrVTrJbf+Ri4ydk
4JHWFm1QpmOCD/4OWSkHI3MTXvmj9zQhipdhwJ4d6q7AQTvbN2gwV76dVHGG
oowsCSW3dJbC1INTSj1/rhdIQTh5AlEAbk6RjsrA70AwTy9S0vrbD0qsgcWz
blsLLDsEFHjhVmjqI18eun7SE72qcHPDOuC/9lfRmsnBGGrUdsp/7pZflC5B
jfYxLC9jp6VCpAyKgrSbszcAlsgUkc2o/snVArl1HaTN/ES6OnMJYtk2IPy/
aap9ZY9DXhxyT+OjsueDenGjRLBcf8rv1TPNL0urQUUPSlxPc6TOUOk4AW8l
gVwe2eYEgTK08U2Dc1Lif824Ouyuay6XVIItQEX0LDhNClFzNfIBM5Uvbkki
WTb4nrJL9Pl1piRrV0lnI7eitl4c1OOcWo6DHhIHAste6sdVmqaIqCwTVOOu
xTsYLx41obsL44FyTzsYjUGBZaHcQ2Atb5c2YU/+kuho772EATY+ZBS88ldX
4ISJtsu2+wFkPPBdxWI1Wjf6JtlcA22iAz7hjHVn/MRHJTK1/I3ryH3YaGAv
hQJcKO0Wp5uOhwK8vkshCmGgHNKdzhIknFWAl/by2hV1Bx0AzVFpSv2JsTNs
cgvGyqfsFv/bxNXnlj0f2L7xBaCO94ZKHwG7zAop11blybtm17sGre6XFMdp
JTgOE45AVHh52zmXQusZGGsIqhGNU5CvX87czG/e1of7XPaEQUlgHjuRx2/v
EXzAYL+1hiW1nMEfMju7X2PeU4MbQ+pykZ7J6UBxd5lyPJQTLuruDdl/I5bp
fjtcqUxy2anaHdS6L7NPHGNwG0qo/qxti7VgwpabH5CXzpbQ/5mWjruanoZy
W3/pkzZr/8/S8xDU/DEDuaUsuHqbWFLDQI3Mefp6V99hTWqwh2u2iQ6x1HdT
EhXdWVjxIsZ01MSeTXqxtlVxSftzsct3YH2UN3GDQCyFfDtMXnXOdWj1rU5D
1yfl1tsNF8wpdDuNq0Ic2Rc6baOWVo8zqq1eUb+Al+s8cxVt45hbUq8FRNml
rmizfqiuM91liktK9OSsKZJQ9uDyxTd1If9fF527pq00R3fqK97PrXG5FpCR
Zz1gNsqwqhH5v/uKOTnYFhUkwvNzeBMDySpowJyK/xBFmovsXyYOquIhGb94
EV9xKlhTNxfmCJqCnOuZ4WDaH/o2+wPD/Es/KWv7p/svCBk0KkxNzQtYovHa
W0kt4zbMuUVb+QY70Vr9EYB8+/VGFFFimorusHCDUoEvnOzBlCj2sLAFCuz9
cm9HWizbKUMRZOPAV3km9BpUd7Gk2hT/RuK02S7RSrf8yroUzxkOQC3UU841
4buMFR1pheHeyftkqUkC2o5Pf8oTCmduDaITCgW7ZivFsxNDCwxUxBm2wwHR
CNlkEs8LbYTBC+PqT2XTLxh3KyOiKUmcocd9mfmJZ66FjPZo30sMncKhWVDV
//eZHBeWkDGeWmpJB+I9hqLSm29qthPMqOygUm8ePvZZuVJFgPBoC52oIlTt
kOrGDldfyAJFl1+pjih+9mxgaibEiOv1FnqlQgTFbRyzEV2A3dKKz3pRQmce
FoO3y/RjAvg2WfUcxNFfmfmdG+kTtyE+QGhgfvuWXzckc5Y3RCXAuUahsktt
SS4w1ByUEq3mJGiPUMjJIMeJrflmmvKbYnZdcSZB2Tls9+Bxnm/vHC6zLSPJ
c8s+WxYGu4I5uOUblL39p8VPd8nfII0uaNbvzc4PF21HcwM5m8DMECo3yN6k
NSnCRC+aTEltxkt5cxVXhHXVMZjbQGajleavAiImQ11ZXLo1CypDOsf9EYYz
BU9Z1EramWPAAuQykooj7qp0q+yooXqLJF/QkzEkj/tahhWI03bC0cS4UVHr
XrtJMfWP8aH5QOd3wWePD5OoIbTjGaV6DZcnQ9Ft44yhb30S7JqnQFQB4MGH
08Gv0RBwRwDRcOdYGtTYsrH5kNMxXFQV1Mga1R4G7J6iebuE9YSvwVX58BKH
Tv2fcfrFH6P6OoxEIuV+MLkydw1dSMO++qmX6cLsM6/75UF5SPVpRUvGzdVi
OrJlkI+N1zil76GiGHwyGcow6GfTuYaYPg47XSkuYf6fJ6fMhbzOmDboLe2V
w9raLjga5V1ej8Ngdur7dWx/4ydlScoRs+hTHeYm4coTKlAMrHcgjzQxDrJ6
gcrt+D1KdRqEYyaKNnYYAQXbbdrvLXsZ0j4bxfgtFqt84YHphJ1bIsXfvHDY
EYKvxLY56juicCPyCtYvk9dZyxHM+nlOv685TqeL3ISz4qj0uovRAY1mDMvO
SPjDCXBF9Cb77rCXJ0p/ljPaqUosgBZlo1TwCNbRGEoiONBnx25+TN78tBT/
ip3nhCMflGAmXYnKHjsHoXZTlhCchvXbX+7tXwam4qGhOT1cLt1oQreKzpSx
RJmY8/tu2KND/ryOHKYI9ZYR9V326IOAX1qOeXKu9AXxQS2M9rTq0d4vXrv1
zibhkx5HrSGd+FUXigFoeKvhB0QhV6Bg20a/WEs6Q5IChzHwdRadZFkJcNq+
qmF5I3vpzkPgLHVKuDBXAk1Sc4XlaLDg+cap9H0jFLGzLGSUAfWn8s58Iu7X
502siI3OZ2fdHG2CBOC7jxUwYt3+vYvAi2CA5Dgs5b9EvKvSr7K0JMEd/0TH
A1McLG7iS/e814TwrvPWDYr/cpSlKKlR8w8J017Q1NseyvXqAJ2OOwinfi+P
yIRtF9ZcaPo66EH3UMRyydTQT1eSF8G+jrktn9itgQ9bqJKt8niT3WsyXA42
0WWmY1My6xUR69bjLaS+URl6mnwb1lIDuuHpJ1Er5YyBHaq0FS7vAaGalLi0
tOuewLGZ+UkU4ZMT+4v+Vq3ODF8RoTQCOM6CSPZIpKjsLDSVUXxVFyg8fu/9
O5TzuY25GCCOiKh/GzcMMpZVfGOR4PG2Q/PU3F0cuRe9rpXyTVH74zAUTuJX
7DsgT4CWZ+8YW4jhPH1s7bivD4bRrjFuko+YUIvQWY0C4kHOV80Wvnv8Aaar
0zeJuUnLlufXWosYWRYvZgXmf+zrRaijCWU8sOsMnRrZYOrsi2cmSC84wHOV
MPzjEtmjfcemkbhHhVygvybPOyBSi0jWjmDHGmsrY1pL1Fr6Gv7hm7WwOCfx
Dzx9Rl9omLJwIHej9dVgQIKCIVWPptf70az/6aP/tdyNLLgckTXMVVbLu6Cg
Qoz3zg3onC8J2eSpRsJP+/uml0ZaUcnPQ4behH4pxS+hXjTeYhU3iZ7qRm55
QdIitdQ3BzqCvKGDnTxteSfS+6w+PhLQLtzDBiesCUR7vUlqugw3J2Yg7UUW
zFXymxSykPi7FAhRwuDaCnyRqEfdPq27TyBCHFqwhR0W2tI4vjomOKlWZxSM
5QeNVPMByv8/zsxCj9BoUOXJ9MNAoZ/2Af2VK7w7hkgL/UlqacewuA2O/aXt
yWkW1tcUIwpPo8Wgjnzo3XyTIf4cUgIkVC2XhxJxizGi6CEdE4Q26DzWGvVW
sden5FLuE8vC3FcSCoOFUb8rs/ACrZ0KJgQVqxpxrsYxgR3BsX6EO89l328N
HB3XBtBXNypPBm3XKwdMtCuwEGaMbHDJzpyCVziL8TNTjTreES0QGo/cKJuk
2MwXQQi3PG1bTLgIYfuSqZLMTYYmit/FbtBjlw2ND2J9niyqkIi2DznFZpGt
srTScSuGAqG82Ag1v2+WB9w0Y3iNgk+5R0xgm9zswBbZAb9Xx5n/u4ZFmKct
wxP6wadGZm/hh0YpWagf6ssT36REHoJDD5qLjVum2jzDgolLjCVaGVtENpBi
jqESpS6fffyeeNcfyamG6oXidt07iBUykbDjkEQvnjvUX4jsT0pCZEfcH99p
jO2h6XP9Fyp+dnAQeOOYRNdQWa3J2cw5XuZW4viD7XKs7GsIZoX+VBzKt0Kc
kikMxMBiQIU0611fbtu1ScaaclrhLdI/K9hnqfZSs6dwXJ7UTA3yUv0p2l5/
ixpNAD95PUA6dmTeF3GqdSkL3PpgZ4VH5DxQtt2Hh8HPaDTYZkqMH29Hj/I8
BCMkrFF9G/xq55vgoAjbbptSeOSimCOhkJKshBk1n0VK94ZfnNbopKi2lTbj
ZpC1dsRv1wEUINNfE8QSgAwwhq3vzVEapXLeGyy3rNN9bq0hTzOzghLaamjs
VHuApbbv+fgMgTJReag7uoIKspSGFvmk9JTLhqOXXeI0G4iOFDLm4DtCiAP7
WzmyuoaXEZ5ghR9Z+GRzNT4X0UNrOapvAbo3q4+K9rJOr5ho24OOfzzzz9n2
DlLALlV8ZjBL2Qsq08lZZu/URvXfPfJDwCKyKfKLs8hVrlzV2Z3OWfcI4OL/
vDGW3UthQvFLYPT14fUvYFNSX+runPXHQFt+3h5EVMaMdbjfy13Ba6r4Fuoo
Mzmmd/LJxgphFfO/d8BpCFKTul+RU1R/+6rtbwUIYTcV3jh0KT0JCMj9mgwT
wf2suzY3Iw2LpNVBH9n/vqDwb1fgYojV3VpLfK32lr3a02fDmFuY+Csv8/Yu
er5VAhH63I8z68izqIie1HduXNe38P9iVgs6zGDNOLbhGfdbeKIAuoJHRVkp
L1nwmftePJfd/ulUCkHvz9+md0OUelhq9hwdQbSHIRyiCSTCuD8Oacz59y4k
Yj7mqsRxGNaEaeyCzSJ74OAzI8OBMbNi4stBnuUIale6K5mM66rmuPRq8O+L
hzWcyaClxqBIrf8DtNorY+5WiEMNlVHcWH80hNP9pIKLc5PVmlCN4Z3Q9xcj
vxFKcJtS0L140aL4f+iefKQbELcqGx4zkzMy0SH2rPO9Rgi1uje+nYYnhA1v
vWZmbS9D7HwW1l81O1n7Pe3ckVWGlOTlDj2JODiLGExp02dS8yS1OC7dI9ii
dmJTg4aVCDXw+zs23D1/NxEb27xIjFZgyKfe0GrkkE+rhQH1mQCEtExmz1z6
4qT6dYWv8o/f0/n+/nNwtgm0LRDu6bsAzlaZikNBH7bMoKJ+glo+33bmX4Zc
6tYbeMHhRQcnCQ1pvM/ASU365SwmWo4CdN2nvGh89bDTeiHen7QyqtOXBVE1
3lHpZxAk/BmaE14WJi3skQXSYxScxFIbr4A1bqQC0UyoVxuGttUTT8K4LEXu
9TDR/c6p80f7RR0vwUq/IP057fPgAO1IOYI5e/mqKQadMDq+XlG7m7ZViYNA
wi7FGLxLvLyTZsliCtLoQNZCXYriPotditlVgPLPhWPc/k2oJlcGCd9iLXQK
TFEhibF4Fvk1QKdU/x4CKXPmpopVhTCCqjTXNIyuPyciui0mJ0XXkNOU4xvo
WS7lS2+8kcIg/nPX+61Avd86kTEe6eyumoILPp8WtHV9Z37vGkcdmGD9b8Hj
xw0MOgqtDhLxZc1safhiBQ9yVer1X5XFKBLTRI9jNIUHAWF3VO/45k4QxU4j
XwrUhLeNYFsyr66XpYmu3Pa/c4aV3cCxkuht0qoX03MemKd8cLabwP1H1HZ7
NA7A120G7piTL8Aa1g3x6xRG8l1glNkWZ++mBDBdiR4D/x5OzM2wmB6ghiKJ
+f30U5B6fbqlNUz31JnBv6sdEqiKL1xY1wDx0Gp7zZSF7ueDayql67NDIpMs
QON0IXrUJvS5+g7Ke1nAw3Y1foUsgfBuB1ZOXubFR+UJvoftOmVsgcU6k9bO
Se3wCQynwf4hBba8GI4GgxlvkTcYB1PSHzDvL5teV/fK8nWezvry8xPft/be
zyrTV1BGsT0zOExJsHSZvlkB8t2THDLUkcThW18jeGyf+t+cKAU1kqv79G1U
1Fz/IZb1zMJMQE9wnlDG2ts1sQ3Gyb/xlnb/TpP5TC5fdX12eL7rmMUjHTUF
os2FVW6Zy9OlaQn9Y1+0Id1qvxqfrYTeGUVSQZFOVmQyobFRVx3yCUQl72VQ
HG2055N2yH9RJIFVkzhZGLU6vK8wBruFFmlbR9eQjcPW0BaSs3jsv7ySI0Z4
dpWEUJvoWskstM/gXrBdfZSuBLqrUY7JkGp92+mlF7UCk7ILpAaxCaAFqA0W
bVAVT+MnN6IwWP9qKtdTGFdnnR6Jqj4Zsj03gAwUrj/hsDGLCnlmZB8snqfJ
nhBx3IOUn2s9wms2XMKqzcuF92r53VMHRmPAlFH7FXP+F8NVU1kZwXgghTjN
J0lA6DP0mjMCarK/lq8kYHypZEz1HlIvq5R90Fl5eREJD35NeVtLIaDRo8Om
5CGqQPZGIrbD/s9mbannDscgK+7XinBRVR0oMLscjziolpHqWzd0gYpD+yei
lGOA8UkxDeUpVlMdmk2YC7kfDSzgBoYgyyQvQVGi0/aWQ2YJ9PcwKs3zfx7F
ZcFe07WUDQ43hPDUq20wyk9t5q1KC46gdzGf9MvKpmPuE2obsO4FvuW2vhpd
1qqzm7NUkstY5PxVWJmVi6N75b1ptxfnfbg4yZzJOk4MqCmdR+DkYj+kEl9a
smKUkHHVTpnIQubLZb/qZbTeq/amSrcPZqb+s/DEyH+PbYU45sYrgMqGgRps
1RWQAMcNf6UrReUXlFQzkgHzEnIyrRe8cYi+32wYylwSOQiDt/J544UWAl0E
d6IAZiGF20RJwnyCrsg3A+5g3C6aXgy6F2ha8Nb4xxDUDgxLQrya+c9nM/ZP
Fg82S54g/3HyPH3LJD1lG0xGw5N3uwuKMrJ4FXYx78V8pD1PDpcYxLHxwlwf
mKGjolaO6+gePy5OynONOEBkLZY2ryGjjSdMaA7zL6TwvhCXnlE51eIlDB9X
kh0qnag/b949qL7ZFAtVcnEDiMYdgNYMkisn8u4FN04v00pYtAcQY0YQKYhc
uB2b6ggwD46W8zgJ5tNcvaJCKDHtIZiek8Q6HSWqre411Fp+IgQYoBAxaXcA
kqLq2nwOdxVsbR5iHoiHmXq4JYSLTL1phJ1CDbTEpF6Y0tDwzunVRlHxIa+k
IoelkeNdfP8TcbBBkJpxxWLLbG6xksngVQ1VaURhsfT3A3C1ztXtNwVDrryb
WeWJ4KqSzarEXOsta4P0+dCp4825O677aHDnHi3rUpz/8bK6NaMX/JNkAi2Q
CXj0A4FSsTxPBzXAZQxeel5l3UCTNo0IB/58NiXCqpHXHMs+7VdmlvfzDG27
HXzTRu/yXy7xIJMW7u3vvdgLRZ0iSDmqSFc6b3Z5avU+TozqWcKyCuaRrBoj
h5J+Yu0WlZwMZmsZyygqyEDeljXYtM5QwpPpdnTZvLnSQau996XGQmPG/Hdv
k3BaBOAfv04R3xeanhcU/loDFJfFfVXK1L1+7bvmwTBi6KgI5qm7uCSKm2fF
U96uQgv4lu2ElUphvuLlLowggysPhTn9a58RTmJteN1q9GvKMlhu8jpZJhEW
cZ3Dyocyc44KgJj6p0nwyQhgRUDo0XFqV5RhTaA2ftEQMmFuMy6w7xZAFkuc
fY7G3PREhsdpFYW7+PGri9ztvhcj00HpJUm64WoipPUVRqXRsYrCQysutonf
JnjiKRacLVBM93Iqf5uJphILFIuiIaROuVs7pKmNX/iqu2nZXhcGwL4XBxBk
r44FPnTtRZNxQVpHj8QIYddPS8rPj8VVW9F+pLlOKzyUZrmQ7enXhK3zOW9r
BVRRAsqXWmuXHI+PFKuRKT7BQY1FlUyBudZ3UGiS1OiM8qE1RFg5W6samtIk
kFaueSYpGTh1frPOx+7hCjDVAjcs37pcFt1lPFNbr2RBx5wT+ix9hRsWLxcz
cDFlPRsieiHRqXvkHW6nAbCv980/aBjwEgUcHDTYqqOtWrc5OCbFXJOvKlRZ
A6fducym2zZ2LbMnn5sAf6d4S31FdqTHg7NXkB99fSFCz34r54LyNWXsimJ4
vp87/Hv/UftinYiCvaJvobbPBKTRLmWOaTauX/IrDVf744Yo63ZhH1GmOm+y
gCkpk8tNsQ0Fwl820FLL2Fk8yc/EHtDJKWnC4sSiVb6/3XylKo1LT/XJk/p6
gH4R9iy8rfUcVlDdS5z/3jQ4mYih7tft0t34FxSz1csuJejBbvdRemC9mtYJ
SO18A+ZYfPIwqwsGcDn02V5gK3ZXu9xzzaXTVXtXsCFxFlqeNl2xUjX19vLK
ZNaCMJQkX8iivoXepcJ6Rw9JcoLgOdwxmysrSKYqiKa/gv4/6GFTouzu8rXr
CXPjr3ovKU6zw0xy8+prgIbTWc7mH6aLnD+YC20tMwdudgNwQLC9x2B+nN0C
GKlkEPzzoy00vYizP30zZwrIGAoefJg1gQ1B/KuSwNhrk5Vtlc8Td0ZTL70B
LL8iD9BijL2Z0QFruJaRVtJOWbj6GfiLqLzAmxAjwwnRw5Uys30M4RbYyd+D
iEmYk7QYmX8cFDXE+S7Lybe0CDoRbbLXxuZQLQxn1rUbbt0JrHWmyqsutPYl
gM8jq2OxrSReYWebySw/Vp1/5a8mroP/fvrOqWjIo18r5/bZWIz/VvZur4Tv
psnSzQpT236SBh7ms9zNZFRPSy+XA+HI7d/YAXoOYlVMWrHtaJ2SedYDJYEx
p3zdoTmbY7d8yxtfinVkvE6QTzkMb8twXuEeu4MvHIm20YaMfG8T6RakZWI4
IQOdNOcAopwD8MXwV9GiWUV44318opXec4/xQ/YQ3M34+5Nr8apAyQ9HiV/p
M6e35wo42VvRwzP+g7RSB0AvHJinL9C7N99N8hdvKnRqebsIXE6aO7pqCBMa
ojVFYXW7HOuLVMHoHE1sHob6d+TfI/SpEA5mdACCcjc9nhf1eDPpOiXMaBDU
1mRA6RmSBqONsrpKOumpXMJGBAiikfoTBZVwJTLno9aHBo9ZO6mVpN87vfoG
VfV23TuMw6KKUYGBGc+akGpddEknn1g/sNzCPw5yHCuYvaeHlWSxqhEukfa8
6N4AnG+dxAu5zS/GAr7lk7/ry8yFBxUIzWbyXHFQrl87wDiXkEjCFaO80GX/
5tTeTS48yloFebVjfPtyHAlK6+N7limUcfkJ9V3FY5bBZj3l2PdHO4AZIWQi
q+o/bpEi+SP93YhiexwVOhJjzKGFATS+xGQUnfEC15/NQD2LTNuQgXHy5ZDd
8GOCmGLXaZtRg33/P+zBMVMKwnQx9WbGlbhPLJZkrOtyAtfi3u1zMFnm0/qz
y4PCkOc0qADOgnhafQIiyPdk5tVaDXd+3mvh4PivVRzPIqXw2m6r5i+mt8tM
Ajqfv+wUytUWXqvIO+YrIJPJJwTqhCxKOBtzuaunB12SxFy1EpO+CHkxxiqg
H8srlmlfr0dfEs1Gvo/ZpPXp2fRKVPuf2qoVqcnoly7p/TIyoHO2UXkkEL5q
LF1mCqmrhWsAzj/Ra4LqsyvYmc17hwAi5JdUQY/MzvT0ASiA4us84mt8lqRa
IvbqDqdPox9UbA9jiRNEu98ELMI7MQwx45yfkM3k4k+2EVw89Rd9+bxYx/7A
Qeh+m9mBQKeVSpDj/OTq2Y6eTI/XBUPjyj7sumehbAxUqUuqxo+/hB03UzwO
KAaMV3s43Pv8VdeamRIzuWn1SRiQ1z2W3gX23wjX+owdWmLArqPbCgjLs9g5
pk8GGq6kf+UZ+WwwX9mhoW2Z2iFb8kHY9U9j98XqBScouanC9K2SAWxYSFnr
4h6rqGGKTp7M/+RQN30H0GpH5hbKxMV3iH0OcWdubqj/VEGRPNH9zuSTmf6l
hlU7V4sY767idouQt+WQS5WCQwC7mEPD0CrXv+dAJt33qRTcVFNYRv94Ze2J
2to4I03/Pd0fJLhyIh605axdihyJJ8iuMQOtDUBH6/saUWmor/kduK91WpYF
7dcoRv0lMTIXt8llPLzVO9v+BK3RuT5pozwtmzhnxB+MoRnr3KeAJ4IaSdev
ykXMM8Y1x1y3sGlkO7UDrVJbHk3CqkrqcL9bT6d6KRw6OXsMpGugY2fPyzPS
fnH9yLzF5B4RUQK9/v72+afRkcQcN4ksyoPmlZsAugScoaCbu7+PGPBujBUM
IgXQvH5nkpiCrMIiO+AbTz4BPQOz7DwkGAxucIgxkRx8uM5BlvEkJ15LDYHv
xymJ4RPKELzBsquM3Tm++rgk/Un7S8VNSEe7VZ6alUXq2t++z8mJ6sEjMTj7
r4rOFFDqHW7LEk5RcOBOr2UeMHT+lhJCDIIYXF6xwgSgKncCHDHyHOHApuFB
b4MXgI9d+RJ+91k/WPuUePXdUq3YFgEj6V7nGCc0OTGxQXfLV6S6YVXhYgVg
ultesQ2tV6CPM1DJErf8mN7sG4dSzd9OXKtLIpgM8IE7gaz4CXTtSGWoUSXx
lB/vjlrcSRDxRUX7Tg2V/Qhz5dapNqHc+BroqYnMlEmsvC8lSnh8J6I3N/z1
WDZq0NZfgNlXFnJlG9BiDRSAZsixiQZI0EcRCGnJNgCfHZoofP1a8XlZOduU
66CuI1pgimUSoWbSapG3dBSfs1w59zJX9xBxWsu76V93Dm3dCvhObT0N2R21
jamm/ll7hu6/z2Y7GvoV8Ddi9B5o02zu8Lza+CqR+3oiE+F2SfeQuZMKsJHs
u4CxUeTn5Tpgg27bbL66f6uCI0D57Mzypag8M4mYEzK4eww37xYdGv+80bRy
+0IAMnJLh4Jm3/mU1mVV0SeI7DDami2tGWwjG2znqolXwDrGyXE49Q//nC0A
zyyqkGqxR+hDRQt19aSPBD/80FkbhM69lfYZY0OVWYdDjDKemtX5qXLnbmoz
V1bYFLfZur7/rjYsTnSV8XzPAm1y0x70v/q4LNgs3aCunNw9MoOMI12ONmWJ
xJHjgx8lMFlCDllZ9aiFd39Lj3TPbhbaIvSZyzUsUqfjmJCCKOeC3ZP1cp9H
aYA2TDMiP4irQJrOX3IDecagrmgKCAGFFHCHgrI5u4yZsBECP0ki9F0m9Qoi
MncbIBlFuEFcby2nsG3og24KBE46Kyh3x2DWPww8nwXFa9MvA99gG16vfL8Z
d5Jg0MvesTVeajP761y65wgWj/ZSgI6bcAHmKxVsIpQXVYbJakZi8QKd8PB3
Nrz4Fr19Fj75vZm/7glFNH0ft8Gh83zUjXjxVp/NxJKpoRGjvfyDD0Y/xwV0
eHaMZ5yoan+3EuuBersodrXFHa7TXq5+6ar6+cnsAjdEbKWSN0k02twUDXWe
eSJYpEdTNTt/CmSmkVy0ckJcYHobEnk0znVcIJX4LTTkBFkNGN3ALZvkOvMn
Xn8aFOITyJbsdO7soYvMbdI8G9ey3aRJZEgaeMFp+QRoIOkdJ+BfFosjlT5w
v0SD9NEq6491GJTiP3xhjk3m16Q0YuZuKc8LF3cfkKv2OV3AZxlU8/GfZkFj
f5FticWBL+XBERW41a2TR40ou2dQK2qr/cJxh+memwRlkTGTXaXq6wwquf76
m2me8MfEvCVQO6XmygBIquhG0QPGF84uD89uq7i5v7P8poxdLz7jAhDjMLfx
BsYXIXQF8My+qipmkTzp/GTmr9y2i7B3g16JHlZXHLWDsz8x7iXDFxvbLWVY
7nwugkmO/iZiToZ9mK3BClcjiEyvs/bWgO66WldHkK4879/O+o78Gr6N25Gv
yAlGAv/Kbkj6mKnKoMw4Ls4phY6j0nJPMDaZPvtt/pL9iQOXDulQM9EkgxL/
6kgitgl5mKZ0XEk/9EnoMFNW4yoCKLRfpRuHRSo97VntPZcTcL/osftsqF8c
c7Q+E9KThytDvQARRxahGePBR/dbAiBg/73K76FvQZXpjouMVkfh9u18EYLH
tw+QotOy19+pDmdjflXukic1bqJLOdrPiifIfWnci7rP/S3nlIFPOqGt5wq9
Lk898nMPKWRWQGO0vwiir/BVaaHhPLYa3z0/YEyOWdoOl5C0oZVrojTYRPaf
NSW5gAPtLAZNmBIIzX8ece4KnR8ITX9RZTHcgO3d01p8HHyPoMzWzkAVFFsB
fuCunE6jxoNdl5uiussX0ZwA7be4Wxa+xNe8knlXZ2qOTZZ8UzEZjBofkWGE
QOup6YexuUXjGMMkENAGYp8c7Hu/NssbJXox1HUP0v+3ffQEBDBGL/zTtTrU
jA2FXypwFcV2ur6HBE/trFvl+574shcvOGuW8eluwSTRxl4/C2WIgnxBlr/4
oCfdg60mCXwNNcPJ985vsZMHsVH+/7DX0l/5umYzi0e/tOLLqt2XQvNNIKSA
3P+7ADn5vgsu90Vo3TtmLINvhK8LHw8EWjPNPI5Ru62gAWWlzrpkyKVvISMf
Vx4EegoSagCVHa+NySZ/ol9yMcJoHV//2ib1MeBtstn867cgvW5VSDuDo4BW
BX+rATlliIccU+n+2f1HntQMWJgai+V1dNj5CDTmItvMdTl0h/OhCpNwNshB
cm298VowIcbau0ipV+6XpkKnzwiZ4xhJjvV5VvbBETzbARWGDNR7TbdYHwzD
/p6OXYnTTZrDXKK0HI0m3ChWBkobrWJZE7cz3M9HYI5QGzJwn/RysfRWGq11
W6gUJD+91f5mqJI6oQGyEkXc8a6lGjEH5SrcxQR6buapCoOR8mS7RocSESN8
AX9pUp7ziEkJj+wcbPWihKgw7v47aLturg3LpCgXZqi0XoZglb7IHnIkhCWt
gx74Y0uWT7PwEuthbvnIqpocLVoABWpn239BAqPhUDP3uBTEKAYDil+J7Hjv
QyBdXEN0Qovhiv2E3dWFJ+SXmXsf2HDUddonqObVeB25ZGbmKVlfqUIqw7m4
cw1lRXEPOEwlIrRRNbGRAGoty95IHtSTtPuaLgFq6i6H2yrv+Nx8pE5oClak
/x+bqU/E4KtjWqT/X4PAp2WAi0nicWMGWkzjIdHTU5zPFTQxvuL6LUfzLfRU
lBoI9XAhVZaJXk8ZkchutqGiXjutQot2OcyRTOMZQjKtLK5/5u8FdPcOuSuL
qcceRZrjBHacOKqr3CKtxSmVtwANRUp+r9tgh3B2LhwtktAFGOTffZkWCcpK
AnrHc3adgIp4G3fGDF1ftLByhQ5knZt/CWLJOwrsOrlaefqyaIc4GyCraCGl
B0+wTdOmbT0tn3uHlD7eBXJpAPpUp0HR7Ovrnu01xuHS5dT8OsZZrhZsJz6c
MMde1IfsKINLo0ZujKkJFZ7DHonYpzlILqtpZZxms744MGdtssNiCRgPa2Di
zWzE/bo7Bdvc9AgBy1kVj197i+ksCtJoIQakJzyPdOO65VxOVm67p6w8KAAT
cFxqddf6L5e3Dy3B1QEKIGwb9Fiaw1L7YxypUL4MAHrHha4O3PAsey4SN/Re
rzRTvJdSTgIa2OclcElkCC6nDuuCOzhxiNQ3LMUXzYY/soGtJMPtcHey5klZ
W0F6Zgy97rDc1jOBxpKxjc/kIkNd97wguD5ndyt9ko/cXDR+fN7TZyDsRMXP
1tgEYkd76N8IM9QYH5Y1ximz4fStASZoqsLJln2uybxZYgDtSbeYT4GGXrWQ
/Ldb1q4S6Dp1DjTbA7YJKsq5wPKcdWaHENbuR1UvFCyJR5wAfB9VJ1/w4VsI
QgbX3cVYclslOUmOGctQ+9M4PkA8SL7g95sCzQOTzbq4LlkujgUIsaM47x1I
evjikaQS2VC56zLIzT3oKvpDCfBudTpN5kuQ5q+AORiM53rzuRNj3kfI1rGy
EArcGVvV24skYT9OnXSaAriweSiWbBRRTsVhhN//k8gR/pCsXy247YYN6koi
oe2KJYP4lmekh/DIsQHMoojUYXmTA/HAtC7+7Ma4DPf5LaE3yJKFMEX+HQyE
WjvjKTNmoQPotKc1J+rIoyqwL4wq222VNXTO1S+VuNWgm1nGIlZUph8G+NnJ
9EMjaRoaeBk6UWllrp5+PN7sDGIOOsyMdTVx/GAxCJasv/Zfe/bHCHxnEXPz
j0tfwOeGtS6PUF5ldDxFbcwpHBqse9XUECk7VrfDAPbpe+yxwraAG5vzrPvQ
UeqB8U5sOYbdDFmNRFI/OiTyBaNsMwAyWlRimVe0OS7bZyz1hXJtCL3JK9dE
ZPzvVZsLpku6P4y6BkVHckRNR3SaoFzg3Xtd8I5CjaoDeNylGcxRQyL2xQ/R
Gvnc+vrLsRw0tNX1DzGG87iFciaPUC6L82eBYnvY119ahs9UgRwHFVyYjy0M
8v0J+TLoZX00J36jTjL9pIeNbQ3TRcXdbdB7wxM26pjCPHDvz5RkgRH7Pbvq
vbi4Fpk0QC/B91h0tSbHQmCIST1AdxBDJv72+NwhPG5b0q2pZ5me7sF9k1Wl
8hjTao/GwzkTmw167cSLhd40fY4q4epP7PoH5AjhIdt3OJjtXnn4okZ6w3Sm
apxN+sHzAeP2x52oXvGnGz5cwpenQ2HzjCE9RKr/ePBDJX+Ftv/ti6luzZ/F
xaTrOH0at7q1+mbxeptrrApSA0EdixC6uLrYNSayfqAO5Pei81q22k3V0jnd
klQE0lcvK+C9dan0jSeM1N22VhXCvfP9xvBz5f4uHBHZRMtDh8hmq3mW0+vz
H3FDr003fVRLOKv4LYCyokg12iT5F5KmF52JcaPa1/FfrE3rkU7mKfgjodXs
vhcNlq0Q6VPSweH+j0AgSjCiBTaDtA+3VuOoVVJgxdwyUu+e7TPDiDU5cOj8
lOB8O7qRt/cA91BUU/5qaR+ElzJO9s9WaXeHSzkUe2L5S6ANblQEwZ+nVu1J
dfM9PASM092h0HVCsU4kyTVmFyt22URs6vIxD3UM8IcggPa4dgosGlguXnvI
EeXICI4230iYton40ZPIzlgOzexrEeHveJOwrvGA5aD525Xuk0WUluDiBtao
ubDcsBqQcTP6xLwfc3ToBGVDfzodb+ZaD7vUdTDk9azW8T1MsX/qVMLfhIrb
EtJfj4XXRNTvE6SUagM+7UGuYU80QQWZVXnwYpoVS97N+z2nYaNfyNTvDRO3
E40Rd6dJM7kI9bIP/myLSQfaJ2Y5ITDOV80SvwjrBAzR8l6fLcs3SLppQTGC
iusL+U862UqzeOY1RNVd8gbtn+Q6Gs4o6P9SaSb30hpofEaVRjx5D5UuJ9IY
ry0DMFL4f7TbaGcf/Pz3a4wWecA/7NgG3LWqrO17urZPlRNY4GDPbnVwdMpo
z+SYEiLg2yNmmFNI2tYR1CJg2sGn+Kd260m0M730SQ7cOSdJRfTefYkpQQGR
0IFjqxYPRjPCHp5MUrN1CsmznbRPnmthSl9zE2EbYTAOOgKpX7P5u+PiRb9/
lA0siCMgQmC6kiNLV1RLql4rgB4l56nIVnSyWV9Uj0qPag6uRiaXLly3ECgj
h22DFM90sM7poxgmqY0dl4Zn10CtQ96VKzymhjpQrZwB1yTxTDW+zDfZ7BOE
r3gympQjf20nfvmeZACrXd4wKRccI6W4TuFvSf2iSQ6gWyDHQ12d6G5AgK+2
7Ijiv4CNGHDTnS/ry3qHAf6d1elb5ZboNhtfMC11JvuYJf9IKCKWUU7VGfWS
mEaNloPMja9nOgzUge2IYf7VW0hWUQvPghOKwua3xGpQtwbJ05sHP6HZatOU
XQDs5AN/5efoA68Xi3zGgqJlBvtASIkduiDdy2j3cHX4LaBeQGLkzPniQ1W0
4yOAQ5KL2ckDzs2LS6Mi8cqObIqrpnHhpC7uyzZkZJCL305kCnDoSgCHjBTB
v3hNpe0PEcigS5idOtSGwm4NkSi/J/HPTD0qeO/5rSoMLdeqZr2bRNCtYa5y
fUBqqqYac7/tSD5bd3XXfbMBaVGw0sIsjLsd+l+Lx39duGqgMSy5nRfzCJ6j
1qL6Xc/dp69QyJGK4ukXhMSQZ96PUpgRC+y1sVmivkNi9OJpCwr7NGEy3O+t
LZ6NV8iudU4NgzGIPR/3/ACltfB+ptlkGFnFYWIgH6MiAzqcpC335o8nOcjW
N105CNCgxMBKJCfc6HCgL3ymMGvRaL+oq28oe5AelkuZOOdQXWVhMsVFSgoo
QgaOa7kqCH7C90f/1bOrxcxz4LhW5UMV5IOw3Gh02lHmVxTm6miz4AYFgaKO
P6h47CpksUNBkGYzUEjx+eATYzCFMg3zKDw62A3JaaJTy5kCLD/iaitqZYyB
K281q9v/9wZhbvb+afmhjaqV+ytTOraAFBfWh5abERau6M6MPm3xZuOsYBLx
c8szJMoa0o5BKkaAYsNilCd/8zdN/Er/Sg56ZU9SSZCfqb0dK281h16VnFyi
sDlL58wOppj9LIPolJIYIzHg6sJn/wh6jEHsgDtw1ERw35oyiZ8dj3qKr2lt
sA2KhpCuPfW9BrKa1JTttzAOM6JA9LrFeJJkI/XFNbZPuufKh2N20xG3j77W
wxbVfECdfH/t1EpCwBMWncDVVs8QXrh5sIlQZVQY/BYqCekI7A47njQiatEu
31m5Vez9xyjc95XmYFwg6yPFhHsluCLMgMQw0pGSqzf8B7v8P7xBPMeObQHh
p+qaA5LGX8dgD4wb+RdwXlmtOW4S9xbRONRO+d+f05mg+TelnpIG2r0q6cwU
bTUIoPSBm3Yh/2jZeucL4VPck5sHbrwDlhr4TYFvFCnWI4/VLUqaL4FHW++q
DBLz4tZaSS9xkSkKMCHB2BaeABM7y7yFrrHRpExEmRFWHw05lNGNCfHDkQ79
2eeMEEMkBrSkeui8UHSKgbeXT4hO7avbhcfO7rw4jPscwukIs9nzLnQCxu00
eMzQiJaLJ0u/lp2vuolmhP9aZeAYzEu9zhYzvRrAaucDApX0cE43BmywQoCo
iEyVlMALgjENkvZpds01Px9GyT+i8yFtCqZ9IrDcsX1Xj5LuP5M/yn7xnvzD
SuxNlUCS2vFHRIrUoJ69jQ3/FZ95d+FwYq510rliYRGdUrEJ/OsOUv5BcGeE
HQ2Woan8rHIrQfn4j8o3oAAj4c3LxZfOAas+sw6gCS8Y2intdgCm6dkCmNAr
um5z3LJBn1Is41dwqrjjxGZmcRb7Ev2GFwceZX2+sIpFj6FFVNKEaSermEbQ
nMz7VizGRda76MvxOvWfq31HTiFkYNzrOm8ayBRv8LoXUxd3IQNFOPzcBfm8
JwEc4BlbEjAZORjlHGfosk/arfhw0Lt+fGc4iJnH+xYHwhnshkcLa3n6GA3E
GDZAj7E77N8NNVhea+N/p/WoALYPDzkuQlMqFnLt+AZz08Os7C4IP1JahBhs
O1ugy0eDfflfHIOnVWe3IMx1lJd0ZNcAPq/MaWwPnL/M1AlwEwUxMhpQnVeS
z9nrRgUWje2bi28koUikGiBdjbPyg7G3i6yi7/87tFY+uNxCSKb8Lr7pt71D
hm+dzxaiUVr63piV0c+Zaxioq90GUzsGymi+qj1AkmR4pp8GPLfMGJDw5PhZ
2wJyZ929zpex8ApUzh1oRrv88KwNVIJDq3o/L9Dkgba+btUyP8IlJhlAfvqv
7vJ/gfwJTLWmD7pm4udqkfDv7PttKDRVGqR9qvCHsPHNNaGembZm5T9GhCs3
RkJEkBzHl3HAKEr804Y9LvtyC1gxADa7ZQQEcaSpIG81DTNv6578iTA9ECQD
PCLJPotxPR5VWz8RAXgyg6uYPmDwrlfFnLdEQ+ypgod7O+3RlNyuLbtOy8Nm
AOWsm28nMFdaQS56ANb++AEdqjXhWtA0CGl8Au+KCm7cgKdljadFQIuXYUrE
ASnbqqT2wH7xNRiqTAPCifLBNXpBcNrUwbpVQPa20XkgNpwqsuvlTP+s5mKx
bGF9jzLs+EC0XBh41/1422OjtdQZIqu3EPuiYsOPInKwMgjeX/RsXZWA6MhD
b4MzPL+kvUmtO+UQCI+VTqzEpGioVRxh1+AMuW5rBMN3TkZq4uDSvzlpmOW2
7XBaVVnl4z4ILj5qAhT0XD/XDoP6NdKtKvkPlY1OhGJNUdbdZ8iPujVPzGsV
MCZ2EXqvAaQIkB3mQNPB/TgGdBUXah+mCAqPh0jKEPkoV+wIcyMfsR8PPWqV
OPNrxgRABUoy+YaNawp9wMYy9LeJh5M4NzFnXQb2A6RtClD22QikS85yjqnt
ODqW/6Vm1sihaIHYCEhYHXq93ivTGH/cfv5nAZZHPBATOTrHO+KEal4chpwb
ALieK+Eus6ejEYAy/M/eNh7vByBtlYtTJ5zqFh9OQf0cVP1bQ9+ZmUCIthAF
37/u6AzucNT47Q3oX+K+XvVdBDGFsjNl+5erkChaRZlei3M3EpvuUx8BZiFh
5punPVdKA4UVmgmYCiUvKOD59NU3t2vl1qtXuIlMafoHagvk1YbYHoq/j6sL
ioxD0EwGwo93Ren0jHuTfCguhAwFhATDa3q6Ri84OQSBT/qdrgrN+sg0s5+2
FjOyvjgKBUlycDzdjT0QMTL0faqCL8/3gogN6R+ADdLcEm0xjcUJSggGAraz
Yj5U8Ukfmbdfx9PxxeqpWP1QH5Abb6k3Kx9u4mzTyaNU8p3GlhiGWLMOWEGY
J4rb3X/RF8/CjeDtWtVQkFQ8aAkO/80clPEXgLnFrDx1kLC0zV+1Ji9zEaRn
IMu5zIw+dM1qo6v/WwDmwyZNnp3jTX4r09sO7K3ldBmOxTs0ZgVKanIXwgef
y4+LIIwvbA+4TBzPIbbZLBqict0nFG29v8iflFMk7NadYdJv4D9jU8gdXRcB
vzMCGOnjKWDRSJD8XcmMQAMvAIfnC0grPvvjFvO4UAnSCwC9dgZ7RE3fdJ6k
5yVYpeqclIXf8yljt8uzY6uK7lhyYwBR/mfzjxcdUgPp6khj2PovEXRpYcZv
5xPgfYOKQ+3WWAys2IGpSnCzBc3Y5NNiYdbKG/hufBf6FRYN1z/BAtWP+A4K
xsj5gh1pWHBzPteXoIGb0cj2Qdb2fGu/Jq0z38x87TScrQFZoHLnQiiZ6zUB
9dUOu2GBECDZgaWGfUIMVBZH6wgAlp44OUKYWxzYCG4iequKAmG+g6dRtpMx
1Dqz6bny+r7qJRjB6+RyXt+rRGWH6uaoDVkxprgxTA2wEAe7kAz4q8dZ49fJ
4I4qvOWrnZXU02cJwhdGMYzY0v9VNK2F7MYP/kTPWOEu0IIYgOr59G45HIsa
fuAurJa7xlqOWOaW9xOYD/m37GEUI+GoT0CpPs92bIieL9j07sDSYvzSZoKn
fMoHjfC94u9Si84Vf1DKZpXfa9GYtGmDTQF829JJfOObbN4jrv3vaB+oU8LL
CTJP4TGAH1Bf4evcQm1BkikQjKAxg+nVevHF/QPswD337S8DWkeu2mMcpOiY
6RYLxJts7c/VNSO21iWXuPCzBIT9cyfQrxmjm2zXwZ1E+n5fYdDOgJ14c+bi
WU+xgBE9AHXiQwJGneafQ7kbcQU3dhNesmGYBj04g7QVYUX37lDdg9E3KQVX
S1JjJX+tn7zan5wlb57CyMtPAlZBmphhk4SW9y9/dzcf3JjjD+xtLWdnkE0V
jHpEBoNcHn0BmlduBhs0sy0dWONFci2mcInwqyPEnFDLoLzwN0ltgPzCBpDU
6lVNqk/dYYD55XbZ9vd/wum6e5bEIP9Ts2tCQFqTg7H3g3uCHbkONKV4szii
Ra4r5vYCiprhENlK6sAHenrk4L5tMLsucBubhAuHgm6VDM31YklE/KXCLU1g
62sYsS38Kjek2aDKe5W5F3CEzv0J0cC34tk5dY6a56qAuLLjTinZKqtrZcFq
CCgomHGRG+suhVE7rtqBVfY89zEPxic5K2hP/rGvP3mupKUVRclPJzfAyfnc
s069O3j9vN3FB3UcBz7/pYcTHyELoxZh76x+itYoMpJRazJsoBWxXgjAkcb+
neGhEVyLyO/GKm7cNBQCirztJOX/KFeUiMq9WXdGr1tmXbuNGsNNFsKR2Poi
q8ItO/O+ScFgEvPmKA6/oECS7P4In5SCq2kQCys5MMUKC0Q+v9JCod13HgTP
aaznBuPsEcY02aWWj3jA7yAvk12/0RbnAKCE2OERZXTWyvsW5pzlANfecr/a
iSziSRs9qaT3TtylYOgdF0eSKQgMlqWLyT0r4hu0DuBfWKcV7zkz/gfJB0BK
hyOt/dqCeYZCoTLjQaTpN9+ZuDw9Wm68pTxR4U9UsBN+ScvoGlI0KcwT4DU/
hT1H+szFz9HyRiVZg7q7Jiy25aPSpmwH69Rscp9QDUgED0b+4kbOOvOI+rBR
Y6iKYgPn3OcLJq3r+2GWWyFQiYWGF+aDZnmBiiYndFzbWsm80kLiOhAuP+Wn
NB9/44rfpjv0B0197dfTbT6M45xQG+COrrVRBwOjd0BREeDbNZmACysCSnkp
UXReDzcoaZf6qPSyBTGR69f1TvSV9KxHhUVQBdzxWQ1GEvv6H/RUyAtbrQMb
pZmIEG9M9nW1eidHpSi8kiIpDG/MnMcT8uxo3fvYR8tAa0riVFESllBWE5Sa
AOwvHtSw9JS9CU8hfbM1UeoaoibQD5P74dVowKRbkRRPfoKLXRb65iEJqWIH
fa3F61VQei9csfFaXRK2q2aRhNlZVuzgYR/tlHIKm0EeXzKLlgVgMYLLSFk9
qgmtHnPAVywVITdS2SXDwDTphry4MHu9OaZkP7Mq5N7SGRCQwuck7agAIZCP
WbHDYiJgSLydS+kfAok22QNIP+MKce/CqvL41AAbD7kJ7WFgeJM4rrSGwE8X
YyRT2igXcEb6OM6aZGzs8RJADXkJETWgn6/c+B6AJEunvyFSd3pJrmqsShvh
nkb4/4sUOEF98dFg0fhCri5z2HX+hsdRez/RIsk0WU4Ip5PFST394IwN1fwY
Ms4VrPLutzSJNAF2P/yv6JdWU200p6m4feFS8y0ZzPU7NmR6bSVAE3rWBZLp
gDm+1UbooIZmGNuvq1L3RwImDyVKwZFYdMYUVJoUA9POS8wxR3qjQrCXFMzk
g00sh2TbmyjpU+F9hbTK9loQQNutwtUHJDvkVu3P6/SD//s6cq672eR8OzRm
ylMlqG6OZshq+ERXPqwMUAFnvgn3EMTdgDcb/xPKipVFLg//3UDC1y6fJUKP
SAUFx+pX2yuzC3q0vQjVGVVAtpYN1DcOZCftKTkvmNkhcl/79qsaZ/mTuBCA
zw7w2TYLJwaT1GxrtJehGfZIAquTNZzN6uj+4Df9KipWL8B7gBTzjou3hMVw
B57FTtL0LEPhJ5l9w7n+IVQMrfdZoc6O/UES+CiOYBa/QNtZHMHN4PzKOk0a
k7QB7iyzM75Sl4OMlaVilG7yF9syX5FGxseV0/zfiR7GCPj/3NLO3MVTHBgP
h6hwdJAWgVw0oK5xwDflAbG2PDMsIwqh+wJpxUlW9aagO/eU2+GFNMQTHaHs
M28VBeetAlvZ8TrPnGpyOGwRSVPu7TLexnl4QQJYx929nfLuA9yeRbJTF/tF
7J600hpbQZzYIT4yrmrUMnDOjP/qkFM9Lo5gb8AD8YNIWdrgWoSd/N53ZXtb
hQPAELDiGVlGktEG0foA07NzT8Mw+ZzgBIYvwIOybk5QuSfA3/fxlY03Gzmp
Up93jdM+hBD5qvugEB5P6NJFAauGEM1+t8e4B1VaMCkxh1USYc+iwVOcSaPP
UziaIAqHhV15u51ftFpwQHsFCmadMSDkRlXeQs5o+GB1SBsnRDCLJ5JbWNo1
2bX+hsY6VwzhsuohnVUXUBNQCH9LJo5sa7l91396MB+9CQkzYxDntN4Jwyso
4MT11znV5nH2RjZfcBgBJzztDCN7YoUab/kiVwR8SQb116iAIQsvDiO1EEug
NpF+sig52euervxFWdSTk5VVV5/nEypi5+b9oAMOYBApj0wNt09RlMsMVADt
l8xctSvdhdqQnOfybvm7YycSzdvjwm/AQ2wxVqLCKEFtSSxNFWW/IA+kFlw/
dSRKVOl/jPF0RcZMUQ7KF9LfIT/CXAadASWH9eyCD3JTW6JEJamy7iEyymQZ
HDLalwx6h+dOL8ePtF4v4uA84f+V0T5VpO2j5xIhxxnz1/A1vHCLqHpSOPF4
cS54NZ8KVXAmOzJYlkLK2NsQcctgOm0F837j/ly5iGoXfTu27I1aMDkgJ/0/
3qRqWs3EIdjCFGM3Kmve5zP4dVjENYdJj9tP2/9oHBQBrWNl8mkZntintqbA
1eJOWR682rQiBfcezXcc97dAWuZe1IAJ/ApwJ9R/YFPGsDIFAXwOL48usdDa
/ePdDQqu+XZYLcTVrI3N2GAN3nSHgfXNIcC5NkLzNC/xlgoozP8zQ/EAHZAK
0wPr2shHdPkGwXYM57JCSsXdZKa5Eh/SDoQI1SgkkaU8xWFFWtIlyNFCXnkl
0znbi17zfwSH93KDlQG8UU52LW/dB5rYBWdb/mnb9GaTuBMWjZaOTfmKrOS6
pn9+uMDQUtd0JmPyyoJG5tMWu8AmzuNRj3AmHu4vPlJUtjdslDB3s5iTMPy6
VNe0lom4/ksBhmuw/27d9lFdH26qJfF/B72fDwxqh7yIXYHrj8GXS0UIGUUM
CZcPULRrd3fzJcgr2RJyKOgV+L5BTCxsWGjw07FlwhYKmjkoVGAFKJ1lDNZQ
VjUchiAp9+pThO//gpWQ9Wv9v+qgTIrBYaR6QopcSJxGi754alETRRGZBfuH
u8IvJkKjJDKhMPobAyXx3kJVx3kj2wqZwjMm9FXYDdaoAAWcHRvvU5z874ZT
LHvfrbXUTLE3CubnzcLwuKHu7V1nhXBuKCCvMbxdWeZOxDu/atU9yQhBIRtG
A2kzPXLdJ+BfQw4y5Ce8i4uKVitPB+NrqXaZOm/sUbRL/f+uvssLiDJl8f+C
B5IfEn0BT5QldPWV4UpYa8c3FVRKfOlG0EYx1BXdiYeYfDW31VcsdfU1JBa6
es6ok1fGnQNGxozYNYGfH3peNxmuEzIQ9IHkox8rmgkdSdtq7JAtWnfeL7qy
EUH//Ec2wmWVM4Z5gPf1uMb0JKyxcH3rou9QYNWQD6mdlLoetuGlyuMCrwaG
MoRQJr+mab1pVOktZN0Amu83Kvj1yDLccix1bYO9xFbtpx7AmeNqQ5/Emdzp
qTZRTkYnHkWkhmBk+eWy8t+On+6x/NpHVQO3P/nVRh94X9K2FUlNzl7Tqf43
Ix6yWdrWMm5ds7bnNXpHPnInu4ozlIb6ewht9sIl2idFk+dH1oTKLWeoBmh0
HZsaL88Tk9fzSzRrAFgf6PnRH4LYsqYEnbBRzNFLptwDeiNeob1c+JNQFBXk
NTtLFX3zM+a/HQbZxTWts0QJHhweuaVX8IiYtx8KpfJ5zReK0pODIVJw/Vfl
SrkjQUrmtMMIyVcAqrNaBmKjvT1V04uRvK+gGp+koH5jeVdqMdnM7y4G/Q7o
Cuj6ix7EosBKsxTEEgzi1CuQIVGSAQTPlbdx7KAPZEDOZkhNNai6+5HSNf7b
ENDPpPKjicppGYdjM0cPmXolktGLQQVKV72VYYmfUCc01Lkv2QKpw5IyRag7
UdZvtYX7blAn3D5b9ryAWFZcAjlZqzuTlffGK8jTofCF/EOFVYzcWEE7J2Xx
j3TRcrbcvRLw6GYN9DyEbYxqZDOavNI0ZXZq9oEveRXZau5IlECLBPfnPunn
UCaSEiZRXgmtCM13zTjQkGJGBtJ8qdjn4/MQL4soG3ylY2ftB35tOTe5wGK4
55wgFFpn4uP8kk3RMj6MKFpKzdR+VhcNGWrHedgrfFQj7Bb+ylcIs+2GWFQv
v+P9S6UlZkfemgYbHDW6pcqqDeIWe3WwBv9Fok9e7GN/NaMxA3cwLNpJxJRG
SjQZz63ChEe+xJsq9wxVVxAQ1PXhBFd1JDQKaPIuciWSlwFxe/ePIkeKYImv
JDrxlkLPGZvlITsi/9OXRzIB4AtLIyhs5+JbfzatAUGjIdUJiwoOMZUIYQXP
SMt6tvP+ByEe90TPADBO3zvTMmgJvjJCnYznnBsrKwFQiakKIzT9yMtEUjhU
eEwbAbqRWXnMX7msJZt9xRO25ZIGGGs3zE0UJXBEzMT+ITHm07vN90jr4dqj
q1Q+sHwQTnnfi+RvfZ6z4h4qvJ+1okCIcS6XwQYw4qSQ8VS03ksKaEyFbG9O
4VU/GFec9xIsEmHuCxsywxiywGoQB/IAewxd0hNIACoXGxQFv8Qre5fnJIQA
6xA84aZOy3zx+RCgOBPcAXlnh9UkWKj3El7LA6p9LpLCaDfW8H3JFaKRdWFN
o+Pma2DWCVmtfvtHn1MC863t57LkhFzebBA4l4VdPsem/OxqBo+Q/nT5ZioC
pdkEw6yqLazCV2Y1mGKMq8TBA5Dk2sbqFkjrjjYHknlX4W0HsOwvgIdlJRvV
CNg11mcsfXVg9m0sr8EBecD+f2YM8I3sjPwFbh7kVUj+l07+FvVu/TvuVrob
rWoq6JCnGvnW1yFtZEDWzWOacfh5sS63laNjkUXfjHqRP/nCkeJpF/7HuhKR
ZCBVbQwOzLlE/n8yujoPPPSa/DYSlogcEk3Y8ejDRzC02Rb27ljSiQjN2CYa
If5cq1HwB+BDITaTBZ1ZUBOl2vWCgtgvYahXdXZWD2MbwVqVyN6geDFIVaJv
yEjgzA3DF2QUL7ge9ULp3m9gE0gdsJywEV/nf7dFIvAkA2MAmwH70q0z+PBS
9Dti8MAsKLgVrck7TtcsEWPUFv58yHUylBIhMoeWqYdBFr4c3wIO8IUcoQLl
qE5kQ1OqJXZrNSaTIX2PGBhGZB27i0EychGA9oG2qUKSqVITU3Fh8qZwR1IH
+BX7acfXIpEJ7FmDhciQve5KXsTRwIdBc77QjO19+gRpxI2e0auMH0Wj02Gl
jLk8YGRm56HTHtsXi1ha0qOTDBskZEGb+dJRVre2iU+g0D3WMjy3rX+3nCB3
eyDreWLSJ+4eI8BctcfJXT4E1BRXkMUqc64jCig4sz5rXb8XMB7A80YJC8Pb
xWqJTkyHbGflEm5SSEvMFglb0JQ/TzpLwzxfFWxtS0A/P3R559t8y1++Ja2L
fsrIS01ojxHow0PBk0PgRwFoLbqbbG63/xC5kAYxR5wO9UW4b3xGLfhQb2fG
x5egQAOzwuqjF44KBJG0aVvhUhQdtpjuwo/mhxG+yPIbMX26iA0J+4eSKCVZ
0qMWxhdrQEOqUDORfuuCbmS839snUASaWfvmtGYlpyleY7BwiEgR3jrVHwOF
zhC17Ggk8fDmYLqupriBbXGaC9So/BFAqCCsmr6DwL+3KoSEz3H6FsGyQUM5
kwwTJAYTb+R4wxeH5KOw+qFZ3dF/wp9B6xb37yvxfv3SelsYZwyM7bdsgIFq
vVaJsBwayTbsUaMlFpCG72/+415GCcPzUknc4RsWhiAzOCTKPj3k58EAYLsX
RNmh+AN0nz8YNVKDA3LAnBsV0EX1gdx1ZzAYjI0l0tT+ZJtzlXDiX4uF1mKn
3PLvYAiohyDRAqWw4OtWWxIz6piaIYqIfDm1ee4N8padhWYVZs/Yyj7qHYAz
/7uzo+4LthaKMVodEAsgL3DAN62B1k/LdctTkSQAIZUUa4+SmkUr5sHE292q
wK8NWo2tOchpLqmGKP9we1GlaydUt+UZZFp5XBF7VXPRZiKN2CjXcxyLxv0h
hFGH7Ce/JRYXKZNvjNqoLnptB8ZxNFzgbohnE9cpEoplSju0zW829asAEPgO
fpog5G7/1K7Ufugh9uLsPjr/76tX1GJusNmMH61O0sCaBv1WW3l7xrtpsl3m
KMSbzky/2VBIRO59w883nEi3tf+cb+Jk4JkAM21/8W6dc0lPxdVGlHgdzC4w
aWHC2HkTmfoqD7VNshgsstcJmyPLlZ0WdeJ0wk4YYAMJJaFSjVH41yRM88tF
Ukg5IfXSg/fZ6c9AwQDchmnBwlyT/drvEU+RN1Cef7DQZvEmHrbkwKBylOyY
b/qzGcG6yyNhskyI6dI8PcFCJ3QudsU8aTr6zcnMvNF6NOl1NRB4NonbJbFT
4kJ0cHfLL1ZhMfPdZD7gg+yx/IM3xA/z7huZpZJFBE+vvMQ+vhtq6GyDDzDU
oMbt2c9BbkM8bhv2UcHjEV5tShtQ/an9Vy2o5w2wkrD7ehsYWiPajSokOt9g
lYI4Bd68gspcL26g7Z96PBFyfDMV6z86c/Ui/juJmyfSZdZiG8fBMCn/P/le
jOILGzLiyy0uO4hvdITtM7Yn0Z73aF9n64YIdOdyAyOkw1F62OxBEiXYepTw
f2/AfetYpDw0nNCVwYwExt4iv3z+MlxZJHg7CYaiRbRXIPQmDcd8r6WSG2UH
sbX27isM6LGcJB5g/KXSa75yey6ur83w7qxqnzI99MIjQIwnv05YlStFejt7
ATB0SoPsKcDqZSreWSqztRbZRFv1Ey6vATcVfUL9FpoTiU6yCjdMAe+Y37aM
ZoqKLSqYHlc+xwlOcGDGk/vY5s5uaaZepiCnU9B9zaxw4VB1KknAhc35F6su
/1S6prYFjG+dRCTHFJsY96LLholKXOF33eykdUunugsOO/g4Y32YfogOtnCI
+HIY21sjtXDolcde6o2hQcRmywz7r02k6rfXII9gfx+3XIdsPWYA6cuENitp
Kbso9VGWMRMAjVGJOahINDpojUxNLGP5TsXpFm07jpSsJWBHwwrjbelvS+I9
CQz0UzER6ifR7B40GUKjsVIaaQtdEabb2JemCtzX+ffUp9hjN9CdsmajChY5
SmACXptbGW8e3ClezW/waOZEWYu5yBW1gHpurZon675bnD7BAMP8nort97if
udscTNoZhwr5pGPyYp4w3+j7s/iH5DZq3WMPv//Dr/mMFQuxr+JLuM2NOIT3
JkDjTVwoZ9EmvvuHOucLZ/ZNTmHkMaVameZm4EWBajPfNs1fS3I9c/cWp05L
eQaQo/kl8YpO+Hj+Tk+nKX/4vfKf6RO2/kYxMBqHH5MIKf/0DC10uFqKt0Tb
r1j43nP96HIsNRIVyNPzo+ZeU9h/7NBj5WUOf1JMEN0SyKwV6RNEtweCdte8
luxS3Ukfof5T8BQs/DuYMHlpOrFowjJ2YHDgz4otzhwir3QlwBCxDe9p9joM
UTEfP0FmXuHwGOymf0NNS+4it8pW0CQxsw788mEpSEn6MvbpeopT3jEdliCY
FS3O51s0R95wxbfLL0MZleBLEXkk01h3goS1c1TlUClABF3yHpUjPIzTbDjK
oA44xDtaM9D3UNaAC8fDcNUyXRUtN5ENGrgs2UIapAp6gcV/dWh/Oa8Ej+q3
hsnxR+YidvP0/QD01NyBwr0wmRa97Kt6p3aTSAWTLPKwMvyy/uVPa/CkePj/
eGJacovd+QGuPaxlLN0+J/k0l/11osC4aaNymYcJs2YsDg4tjoFiD5rPNFwn
zDWjshaoX1ov+tju4/rTi4DlCZ34XgRixBk8R/pmhpXZBI+n9+D3Lu4Vbyns
thZTXHo+HpAgPb2sasJx3cGnUlr/5zh/FtxBhP1Sz6jvrOqiyqTGnTTDegIs
P9dlw2GWz76reqdnGL+fEpDjmHt8Y1DW3OVnnhXeItGp9oJqy8/W7W7/8ci8
bdovCB/6fPBkditjudq7M4oieFBGUlJ3EXndW7pNdscIVSJGgrfzNKDkSDtL
abgQ38NKKAr0aIcndS9FqbpQO/ZAk5/G7lH3Hn03bDdnlAedF2HSmTh1Fcz5
Anm+KEaEyN5HZRQxrbm4P1fWjHA3yJNbRAwxZpeDcMGW4qVmXDLJFeS6NzDU
hhex8CDfNPhpYuAXWx1hyyLi9XTitGSPkTb36XsmeTRR4wrnbijUgrXhk3jX
BKHX2HSXDGKuVrV5FCiqvQJAaGhyskc+oElbEFuAhYgdHx+tahsmtmnKzxvG
btpoMDQUyTWR1WDqhdo4LTkS7KUOhLDh1plkHRYTVn0AosoRwtdP+AHqVvlW
4bBv4G1vrywK7BcpLQxr1TizucuBMwwOEaOv3ynlaR9GBuWP1wp2Q+RPnb34
qok8M+9x3A6WjB3fXUzuudn9lGu89OC+CHnrD+RFTYf6Kw2Cj4mVwhy0UtHB
hBOW8adJUE0kqIYwCVTDFYKfnCuCiYcVehavzzsEi4hp9IlBWttmAqYOcr7V
pGruOoJ79QSHkFLPZ+xC5fC+h9wMO+2iPt9bTZYxw9JFxJ3Iu9Xgz6W4NAuo
Y5nBNq2VvpVfFPs4R+3S24umL/tzoVnbEbtTPlp4IekMnJ9JW1yMlBx58HCM
kmQ2zkTdRcv2VigY2KcMCBs8W38UiVOa51o1LeS7TrknHjKcN53MSlZfvyUQ
5+tOxmq8gBEOjB+MjUOUGAuxxXinkiNABHEHcmsFMAGwWq2heSfRDdO72qW3
d1Kgdh3Yfpvd9o+eN5MwwlPrpJwm7tCag3kIILkhBi7NEkIpA8KsJ4S4gGAR
/kWgqUMB/SINbjZICR2Y58Lx87KwnnFFnMqRIHo6D3aG7zlWuWC3vrjq7nDw
zKxvBvbKN/ssQyWilLBWrI6nbnVROZPWxzQIYq5R36IMgQPSKNXC3i+/8xuu
6OBXDXqBBO0gr4QQnxBskpuAH19HDJ2lWXY61daHvJ0Kwa3bXmAXaRHtdhY4
Pm8YvShgK0KUwf0WyzGw7Dm106hKwg8tF/rvRlh6+xf914YA8/xK+w22jihL
uB/O4/OTj3ZVlKn2Cv5RZoQszvLOcVDdf1b3Bk2H7zcFrM0nSTxBtrcnD2OZ
Po0h6XchjU37wTq49D/xTA7LbqXl6e5OTm2+aoLgfFOjnAteW5UKTigtaPde
FDrNqZDTIzySrxEiNy03ldBTA2qFYMk4n4xtsTn11pDoVGodrRnlgYg0Du9P
StgNu0eeewDhBPlrFlBm8kSHbjvAA2UcpSpBMlUmiX9xo2vca1mEpw3uf2bA
4TjcMU3cN8DUDgnmojIaUTsq5YdbfmMtPRDdcRsb+3seUWhF0vRjYm3yNFxo
YM1lTjDEiNOHrAfEtRTP4pHzZefvT4t7abiZmwUdxPhekft3DThxGMCVANWq
fjC9k2jkXqWUKLyWfNtomKIAM3n0tbf8ZwUyrRhdPlhu/rFUIGJ78k6n8XG4
Y6iPotMek16rOqyim70oLGGa/KsEU3TMXHsZ4KnpG2zUphDtY1kf9/TFPTFX
yUvEzh+vZFiQjLHIgQK2fG3IhxBprYl4qQ4rdYTRTJNEr9thIdtxXeY6EG1X
pUB69o9NExLr7OMbdUyJx40uTtw728+fTioDyln5TRt1Ff/tbgs8QPEAVahv
HZN4ZMqPlLgi808WQHh5A4pBbeAwk2VNfvgnLEWkMftUA0jir9qcvL4AgB43
RawRpXJDXC3mArKuPDtauzjGOAWvFs1HfblBDi9BPV7wHruWNdbnUnixTfjK
nMU4n5BnISZAix0mE1Dhjg29xNfl2IGA0lF5hjeCaQ31P/o4iGLNfva+CcDv
fw17q6Ruv/U5kfCisLwXApbB04f3BkvUA3IUQr5VK+P1tXV1ZKcRThJNcghK
oQeyxUzU385j/fJwDEf0BIhYLLzbQwSOtb5lbiEya6lumgLIvMz4OyzzeoHu
tp7j6ju/DerWgs86t8ouJXGfABgBUyj9+FYyodZdxpW+DLjjP52Dgx9fD87W
wk6m5ghQ4SYL27MP0ZTWBKq/TdN8ysnh3BeZUQDhJqO0YZthNTGGIkFNbRlD
Qd/zzdzmvNBdiBDVvYP4B/NC+VS2pF8HP50SivdNHhwe/YhEuyTBOL83afkK
EGQq8qFfZoohAPGn4XDqoyg7+wwJA6e8CysxeO0xk+oTscUQ/99kyDxTyKAr
T/+7rWTQU5TkVewg9fzuAXXvxgqfQGd8QOXbvNziVlq20pFNvkjUbuvxQMpm
U5PZ8cPs9Z0GMPOwJGis0VdtGTUr1Sx6MjTL5haglmc7SrYsDJR80tUgCjDl
7vphFj/TAB9W2C3JjR5d9XS1+vUn3hISI4e/Wc7gikNXZ9gIRwA0f3Pe0D3H
zqwuITleNrVHZNkhubhcFtg7XPOxqNp/bEbndBRJVIX9+McKi9cp73isdCLV
mitkPF5K7OAwb/YWvBbepdnwwIXfbFgDVVh45TcXM+p1bI9vy7OeHzRCCGsm
anqtv9yl5ll9ppng8TjfJ0gSGTQU/lAGvPORghjPV3r7EMvSdbQQh2Ec2MOr
IxAdObGbZrqG0Jry8d936lvGDQZqt0WUtfH0alHc4Dm5vSAaoARHi5UluVOy
2DJOnjLpnzM36CP7TLVPPywfNTqyhg3ckGWzJ1f3oeeDb7V7GyAyvuu7iHkh
djkpVX8E/Tb+wt/odXf7wwBWWquO+rQgQbzkFm0sDhRlGKKj7HmrX+2ZvT6H
H8ro2WuZiqQ1sOiEvVGO6qx9ClFJ/+U/kxWajL0zwnGqSVLMuUt9GfundyFZ
bAMHvw/l6v5yXogac9Q1/hNczdEi70yZSOIMFdisvfb/Bd1qaPSAQ1X0rMT0
fpiEZ1y/JciIfizsdIwemyOqkDivTPRx+pNFIJNai6oE2Yb4uVUC/bh7glr7
ybBxVNCUCqo7WX1y4Qd2RuBW2747VtMz6tp2JqARVK0/wa6cc1jI/VS/Aqrp
81yugEBrU+UI3KDe4axVSN4QN+YZrLt88OJBRhfQEv5g0L4t7mqPZF490sqI
6FqRANz289d6ArlT9/W9H8FTMyEFH6kQVGaXru1aiBW9Wtkv6LOmBSUrFhUz
44OwV0vSjglMGIvnRQy/+20RCm6fNFvjwXD0Ce1xDI7FU0HHpSPWwQySm5II
LlLABoaZXcZu2n23Br6MbALqFZ0XH3brnMQJ3Rn7Djx1V7CSauJrPooUcBmS
iog0MOOnuBLc1PVne9/Tg3Sef92FYl2JDBTK7iQN4WmFt0+YFXV6jFrknSbL
RWMSzaYk2KOED6Ke64EiVXIlEO4TLrh4RUsCkr82+nFaWh4KQf9iSDCT4Ly+
GKI9//bM9znjsZtJeZOs6SGc6lvc92VlBmqPti3DBnkGMo5ExVB2R6xLxySa
5ysXYkIsdjEq/59uTNvhYQCntwPaXrUGgk7WES1V8czoIHKd9tI5JQp6kd0t
WCbNj0zpoSLSBQHLNJV6flTwneg/T3Jg3IvyLjUzmOG4XbTOEkyouCh2xAmt
0G2/Vmz3K2oo4vobS5B9HOyWvG4qYwYWc7qJgMSmTUlcoHbtNcJTm7SHxML9
wkXrMWL9o0GpyQSGZF6fZ85tFqMOS8nYVLLbweEWazqam0aLIb0+4MRrpKOq
IbnlALyLfS+7EVUbqjgJ6AcZw19Jvuid5ikyvJo7dg+GCXWXXGydQ2iv7pSF
4dPf9KtyWIfYFIuls6ddty/KXK268+QZY3NK3B8m9KJD3d0fhlEz87gC/g1o
PlNIlQsPTeF3L4s6ejD4BMONM9sI4roXakLPJakxCDw97WqVSTOXthMvccSE
VXuIJIfoxlIvhJMZNpINWe9Wn2K5gxmv2du4xNkIHlFBQlAlFr9b00Eg8Hrb
OCPpx3AeABHI/91E5C7Zo8aDI7wkWQ2q7WMuGGoFCWWBQpgoqL7Xe4+rDkWT
/DUs7RYWTWritKuwqnkU2RBEYGHkmEiURzUG7Hw3/1sNBXhvCJl5z0zs4khs
bg9zOWmZduj0TT7JFk2D9aSaouy4TRSd1Q0H5f6XXzgftCNNOO3lWtWA4wzB
7+tijHqA/o/RnyEuvVkgXGcxfWwAZ/nwxy2DuHNaZzsWygKEYMDOIz6FFbZl
l3QL7E5Rb5EKT6pGq/nro0sHlM9X/YsNqImh2SxtoU2u5mpLOhRI3tz6s0gc
oCC7X+ecN3pTM1e+CuUWynU8FiAqUaFsKShRmizB4oAicaY2EliMKX8TtVt5
K0nL+QQ2tlcflIXP2Dozz7bJS+V8LtoyKlGnCD8FN4yTNheDiSZvrT9AeyVS
tH1Szha8UoqEzTw1qyrmxJuhxlb+sCW/xIWHNIvOSocDKPpE5tRRZiHBxzzb
x4zTAwcL3zpH7MeiBqMuu7qLUQ7Up2WIG7bw6O3D5eymrsyvbR5rWX7DOHJk
KgmEKIDLBfGeIv9R/oqow9v9f+v6EAecdR1TZ6gCUaJmhA+opX3U2wpOGRGQ
ZO0Qn8xvW8aDF458sdqC3z9mbFwpnrsRD6UMNBTqrfRUd8FSxxeKDwTL8ZR5
65jbdQZZV8ioj2xCqBXgLhe40v+INu7jZdBrIp2nQCGH09LZ/lEm0VXCW3xm
WA/HPQljcQHd/PhsdMhRy9bMf3sOvsN6rHeZQ3amVe1BF8RSn3G69nwWGZfv
5mishF5gZRVujj8JQyb2OzGQnv5KAzlMuZtprj9KwtiqYcbkJBQJ6rfly76h
PN53u6wbLnn3eLug5u5ZS2u0tSiTEusgTMhY1UYDN9rl/YPk5eJRXRAuoEoP
Rm7bdkC5WUciQEmlasi2xmDME+HwpCrBniK8shBtWtkcbcM/SXKIlV8QgSzK
2d7mDyFVyd1vxdKJOW+QQerfN6GANt2SBB2RwqZDXox5c1kC716YSEvfw9/O
82OQXRoksx9/ooTH8xfgy7GNP6+xUiyD///NeB198qDCDA1TgafEXNwnwnE8
ObJatZ43uJnH+20OdsDkHu7Khceqn/JlkE7QaAbBsTdLpNASB2UHmYfGTXge
LpbnkKQv8tw0xNyb9U3zVaaNjqvSZXY8DHgmv71AiqeeWH7zaF2H23pXfKPD
2q9CW54NZymyeBMV5cs0xOs3L7wPNQ/ox7rhistlwQQq/GvtWOlaN9VSqtQK
XVDYKEE8myWOOtRorR8ng/bD52tI70FllQTNLFWxZ/pKNLUo5l2QDI8BR9Ff
Q2FtI8rkimj4xBYtcLMAa7QxVARS8327mvjqxcc7FgOxdzD6tMtG1Zc0rsDK
YwrZsmhzjwxWwHsetKuMSq1dZJS/1I+kNu0IRyW+oYkVtduGwkWwM+rr1nxr
VEJtxMAEBIIhw4Cwh1wX0Pnm6u2KY/e+ALnSEr13OXEjlyZ2SEpl7g3HAzQ5
2Z6DuAHTWGqdrCYRbfuQdEZdJLhN5R0WKc1IQaddUtCP34QOhQR5g9OCDMfW
ExOUWCcp1pS/Eh4y2mDErxLzqRvd5tYw+rzi30rFnL+h4yH4jY4rLnJeRS8o
Cr0k1y4ar3VarCM4SglKOb9XybJttL2RNFlStPhyG5lyr5/h2Y/wlO/SgGuY
2c49VvcWhSbTCeqxq2uogzQQMcO36bhOvpKaj8KVid4s5bQ1BWkBfRGu92Cc
WEe4jJnrpTMmt/XAnc5AIqiW22t6maBEKSo2y/SSxTXnbyT6UsRk+HLPe6YT
EpRj1SOwy3I2RjzzX+YtWq6rxxrCqjd/7uFBPHO2lPrlfbWjyyeYDQEcNALk
Ay5OUkdRcayS0O9M7OGaLGLgEHWjceDaRrWO46EN7jGx/4NcgDVuTTQsl+O2
dTHSS8FrXCxpHqk3vq0eHUXBXUxsYX83F35T/Q51TvbK55itAxKwgsaUaZxv
G1VvhV9D1SUh+G8xlXY+6wm1XMvUjxjXERKLOuRGxpPIEl8ObLaqokGxXCWi
yxw/tUwvFdnMN4PRyurk4KspmUPz7EN+A6JYQoJQAkitJgSElv17U6CMUivb
NhvDcExFGUOmqkgrpi2/r8tMpykboM70xXCr8bUv4PuWSeFV9gqbX/WK5gdU
Xg2E3lMHF+hLDsXBpuRufmFsYNxfeU68Rb63CD2VfgzpnVcGamRmIT8eSu1H
TA+u4aHdl6q0+YwKImTRty+98t5i0WYIa7+Az/ieG8uUF7dFdViFa38+TCU8
TM/W9rb2O4yta8cnyR6SSIjtn3wgHAyW/9zil9H8jE29tNhL5gU6vysGoCCV
oRbkyRL397YzvwOXGkTuS+dkgNq/Q1o6UEIswz9pQTWdGPZYu+i1x9gqlA/p
Q9FX2CtyxQ9scRX35rQeFcVMpmbsLVbKDCVVf3+uFl07hrsTJNUdhfOu2rg3
369XO86aqyF7Pk60MhCRT8ru1wNLFaBFgs24upIL9h3yIbAgnMNESQo3UW6o
TXmY0z2TFbJ5DDfiA4aifnrNA/t2byTsNhYMeg/MEHyAlX+TNAIKLjXOnThg
xd152whMQ+fXBg1zC4s9z77fPYgIp9Up3xr+m6o0lebFM+VKStqFKaxYmir0
V//gKMi+jUs8TL7w0Ty+R1hAkBOEcU4TH/g9j+Ey9ZGwAdzY3jKe6Zq7Zufj
kUxfeK1GQD+wWqB4nxZ/txuBEt3jSI80UDDYXrieBT6cIjaRchpuIblkocix
hXykId1QpkdfJ5Xtld8+adJHOOVp0eYem0iUgZR+pd2xTKx6n0ALQmEern4+
STkMz3bnKbB79gaY65FoCvBLgVNZZudCoIR980aK2k+8Sf6QnJ025jY+h9qD
4OoUy/rhXscvynRwUd8zzXQTswsmy5rJO4aDYzzAVSGxUBnTT7s9ClraeLDn
4uxjFbD6yY+hwAbS3VgerlQzFMfPOQkAs6qImjA+ZES5LC3OSPwPYbKxj9uI
Q0rR85AJCB3z04/BdMeTxjq8p6ZoAqtKjlUftJquHE+4cYN+RW2wjryBqCue
1Nb/QMmtks6MYDB1Iflz2k77O2OnAzNLZZI6lo0biMtHYlIH++nQnsEPCQ+Q
Tg0umaWxn826OqTiIzEJInbHBfgQWKWAhd0LYuH7h+i7LH0cUB2VW+NY0lVu
70wx8dYyyMyhasY8qN1ePb0zJ9Xecj8tUWmi1+oX4mznQvmUESJvTHWApkwB
3WIJKc2WKV1kq7vCacKuJ2ZxUd1WGzfe5EQDn96aap2Wj7YVLFTheKVYaEe7
7muL2aO2K5/5tPWE/zBmcWKLe7e+EMQ7RshE8QCJCAmF/iTYqp+h+DoUR8PH
TZ5VC9TCz05QWZuccgr9lhZvJCcUx1PRSgM+KQu+n+M1eOWJ4v6MfsYoGTRn
F58sUc2sgsX/DQX3sh6dD1WDwiziebMR4PwGGopTyzJpDXmfNSz89RC8WP6u
dzsVZzzrUhci95uJbeMRQV8LdpEcqsH7seig2DA4oW7vLmodarbp1CBDazGe
veDHgRwa8QYfTG7WyBMe3IYXLwrU3dsXJ1CemCk248VIgQockTFhnC5WkQOR
y0mT9uAZzfdtXbfZzEqL1pUPGzMl3vbZj9BlbfoDB5LreW6ST17HKk81ywLr
k6ZtcTl2CJDAY3Aiu2k6wviHjIOrzpLxKmk8AyUwa18L5EWQ43WWqMDUye1o
khn2I9lCok5c7sAPhZLVYb+qkbwrc7dT+42tYc3q2GF9gnjs9BExurXjZxe4
lyk7v2FfHeV6tbySEc/ZAnlNw7iX+sZWzF+HHbCS4hK2VaMERK98JFowlB7V
ezK9QhLmLtNHoo0qkPsEYtbJVjngleCImf49EiCsLxPmIwhf3F/lSYz7aqw1
TkUbkztiIz85r8NszcGIw5H0xgohKSAc1FqZ+J+PrfyziTRy8IiA0/wwRy8j
cFt55YylSUttgenKDyiPH5cuBO59w2XS4Rl6Gl4BGicjMFlLkEd0YoPmdeme
8HbQkqzKiBeAZCjDCEQlYE/41zGcBySERfasUtfpcTnDzzIzFjXuDWbXLmZu
kQvKlS/p4huzt88XSm0sKhO2yL+vB7ftmADsqi7o6fIAZSZ5ds/8tnBDRz7B
48gh+9YkyEx5ip9Fwau94/ZtoJ+aOG3RL8TELCsy3UO2EUsmzPLyJXRJhdH4
+iBp3TNOoMx+znlQUshjspNYeM75TLuWggqpnYiCyUOXerRZAx0PsBNA1K73
y1tjR66dyJXb6DeACj5MJQNgvF1jgIICmnADlsodNa6cmUemN4DPchVgLlNv
eT1CFdv6bnIzYhG6GoDGYS/NDJpm9DKvXIvNrJo+MrUZ6XArITU++JtpDdSH
jwrY4tZpyobbKwveZQYhdFihSb56PXzmfu7fvIMHOyR+VlJECDuWru17yjgk
LVtJiZylWlleAQR5r6tMuf3icty9PeW63pth02xkS6e1sMwcrOB+sALuOCKR
x0zUV8RO5odGtDdJ6Nq/Jbl4GYS2pEo+6wz4oDMZxVWDQ6Xi9XFF5sbJtJzH
LOJcUTTEEVfwmrT/boSbDbtDJc+7vf9NlZBik6cYMhy1SjPC8en23E1hebca
11HoxGxTJjeMTwjwwJEp90AbP1IqI2vs58nuUOzYDwT/NLUPWk7fxFQDfUMV
E4NhOsnGjdVFKQqCOGAh4uH9r9f2BJY2/4hFte5FFAPeibTgBXR9EvxIg9fL
Gwrs6/zCGyALW8paIX+//zffjgDKbXG5JQhnpNAbhiIswvcvqp0Lv5vWeqGB
7dNeOuzYWYyRS9sgry9rcfcWXGeI7oqG0wDz58g6Ku6HZP8B4RgLlxPrsBNj
1V8eHyUyej6XtcdRRRFcRDc4JMIHapMC5yvNx1/pP7SgEm6hDP7xxPQa+sec
3Elax2WSd8xcPywqsCXMHG2lERycTu4Ofw56R5o9cvIqcUvbPjKw1FrFWgrw
QQvcLjuIh/TXWR7B5BYOexVbV8cOA4/Yn0aI1HwY7ycXFQ9CNi+U1MfVLHL4
sEmE4YqOGt/dI1Sm+X6y72j4cWc2rNMuXKwDpd10ZsUGuoYUU9RMAhphAS+C
484/wu0ZF9HumAyUVAYt44XU3sQx0QZqD4zRoVis4g94G8fdpyRSzJZluHO9
hg9Pvr8FxO8GEcyERhylgWPveQXvKo7msUwlqa5prppIu84lci34ESzONiEW
ng/xq3XkFnbEIUiLSb7CMH5iJnTXQsFbZDZd5BIqqM1ICM7PatVVWumS08AX
JG5US7u+nzzFxAIYgkWA2OVAqwGx87iwplautO1+xr41AP6eY2gHFVXuKo1L
+5PUw4b/US7B6g1FdYq59Uii+W1vdvWD+tvh8RIntdmKrqKyHgvU1UlTFVW0
83MZxFIpzx9j0FCalZdXkaJIkVmlxNalYee1vt4uQEUMFAwaUdIB1k7qeN8U
gGwxV6BUchk8QcJHd1tPcrRz/aw6vRh0jN3+DbFusf+PFG2QqgIuPasGttu8
Hg5sA8Pw5Ee7Y+U+2IdFSSEN52rFIUEqEB/UERT52LKlVgP1p73+bF4sY+6b
6jPTvaG6ejlnN+J+hGk0VVh11tPF0GsObArmb/AEOMwG7OnCUVhKdWbjB4I1
0r2n8FhplP6DKj8nprN62LTHKFZLXDGcL6YAZppuuhb47GoeJLvQeX8TWPdT
8TnLR050wY9jSQC8NIkYIcGUWZcjYFp0dXSW3arsrC8QFP+ZxyHa1u0jr/8L
VRIKwGJpVOnctpgjedSgEiZHi4UXTIDf4Htg+AYPesup8+9AEgACElt10y8j
d4O2NNH3LrAoRz+JNEgco6wVXKSBJveStkeh8X8LST1HeHRD5P2enYX3a6KT
z1kLUzyPbTcHv5NtwV4p0VkinxiK2IM4A8xOTzhDtqRz9QbXNdb3rCf6edNQ
/c1K2MNoXkQHGEbDLG2KXi2auTwarB3qwc9ZxLB0gVHvH3I92paAEIxLQ2j4
R2f4m1R+qKMp1yhLAdgVI3IxdajVaSOsxsEht/51cP9RR+fBLXHuc+EpICYP
+PnsddPJpdMyCHsVXLHt0MK9uDiTiQY45DuYksR+GAA7N2dKP688cKJ5T6LM
epxXKaZLO7YD9cShW/vdeIXKOaHo3OxAf1nwsXy8z94wMK2/9wMlLoZ1wEw+
j3nTQ15suZQMNOsqWUyiKjT6x2d6u5AcYYACfOjp8rW3x/PNFxsT7QmuF8gB
ZYukTAGOVqJgNwoVmPae1mBIYEnUFlSxwhnsSwLalmPYa2RMh77pW37/RCww
V0IIv7eFZqotNHmnA25DbP68rXvUhSphAKvEiuEMwjufrkjEixdKl7HiVnct
W97+qNGiVHNQtao+5dLdD3Na2pEzpnIN0eq+pbh+BSXgvL4gJc5yAqHKEHQC
s8DnIIyamT3DSdrv0tzR3dukFxynq54uS1PEzT7Hwy0rzrkip/QcCwF4uecT
dXFIuVk91ts+WmTEgKDwRpJq8taE8depHGao2l8GOQFWknhmEHVU98n8zcA3
yf1q3XkRuv56eE4eDMaXgw89FH7ynA2gl11Av93GU6g9M0lQHkEU4sFjeaHm
tRBgpR+Aaa9zJ0Ar3Zne9k3MhGKuDa3JQKp6W4Y91CI6uHORfpHWYnEGt4Qz
uyUYMyWP2alsjhgOfDW4xlAw5IXd52rLacFe+Qk0CyXQDmeRb9cjLuv6X8Nr
d7OoRGVTC7YnDgMdqJmnOq4xX4K8GqZVhvKta6iYuVZr6+jDH4gN6/GbuxF8
psD7YjpXHuhxHlgNMMcoTO1e4kszMO/CzTmfLR+df39oy9Keo0bmJTFsS3ok
Hq90+9VdGfEp4JLwqu3J3opRWkItMq/nIx5d3OsiPOwVeyyxgnBoZ067S+gq
RU8OKoRh7ElEaUqczhmvVau7+/iHscsgxhbLqIUNsi2oiNYNFIZOK29zB6JG
AjySpt+YPQs6IzVAzM3oiz/wQw+ZT7LsUdGM04+0TO6+HCY7UNxmcUWeWIeH
YmrRHdLyfHrTRdg9fpvkmxeo5RWUgMZ1o9+3lX3h8uYQyN3U7FwzJ0t7FJjx
Ul1CJtrsfT/perpCa7QEaild6dEFD52y+O77ZMVn0a3pNx/5j308M1cYrFvx
iHsiMw3cHLg5pFbYRSHO/CJRIaicyvR1pT2aKIrfqhoKcPXddO4ELE844QCb
lgJ4ggM+xcI1biakX6Nbs2x+DDYGWE6x81yM0C56vFvfp/pe2s2/VOo2LiTQ
e6V6goFafM0HqE6rnZBIUa0kPY7MRMXbRf6t9ssWWe9q9UAABw4kxZM0rfIB
8nT7gPXHH4IlekVlBoQ48qMUSVJqx1YKDrUMu9ia4DCciqtbvI70nDPMoE75
x924UUAS8oinWq5ByRNl1+x08jkx1VcGufcrSPLl4uqrCLN7nOKV5NCdzxtO
/au+9poPNsTRQo+ySyFpllCC3YulBcpzixbi1PBgMhQw8xB1QoeFx9MFJcBP
M1IswMgnoktimIcNLdFmqENNE2meZv5V+KE5OF71NE8y2wOw+5h/fzheDHVS
2xZohgnyL+wgStCc5rZ8jF9s9AEsLpAFUomOw6kDoSIBl6VrHZKA1WkRDhck
iiGf751MiG3nBoGiftulab/GC6oztmN5uoY6ua+Ev3+Kp4qbhqOOT28X4XDq
jawC/A/XaTTuYCaf19WbsT4qt0uSdDT25a+NGR77tiHri+V2RemLrXiJlNHf
/1Rzrko5s9blcQVkkbXDtwyJzOLeTjiL3jHMlzKedssWZHk/pjrkHS4n68Dg
iIYtXvKIunIdhx9Ua0OqrqQxN9HIj1LYjnQG/QXBV27mybJjsCmn0faiMmrH
FxTLbBJzXafHKJ+lKDrO6MMuELU/OXPw63IclF4eSQuIWTZnpaw5cLxu8KIg
lYqoJ688pWwaGpXn8ek2l+CugdsM4XA41T8c3g+w+4myTrIX23+Djk0QaauL
v4GPmFZA2G0PUjQ7xZYQN5xKublTjsiRVFA/TRB240qeBDV0FgBt0lxt9naS
nQanByM9isIpdVTRc5dOzidDYCAe77PdyWhr5bfohifOOYgk88u+1g6JqHqW
G2wyPrYLEYD30ySN7+ZHKFBPXmL3ClkxoAULLnCOrPUMKd3cvnNH/wO97409
pYsB/ICGDQW4/pmh/SxWKyv9YzAd//6atH0QJ+XXtJRG12DFfLMIImuUq5h5
GTZwH5Lxanr5VzMF0RVzr84eqqZPXOoyFIzwH2e2MI8QUvdbtAJU1xz9sdsP
uEfFW1yHhPlNyzSURP+/sTb/qJAXXatX02XtH/REr9ETaFxBZGkbaIbb4jOB
8MECQ8FfHxB4fXhOmK0D9CAoS868xhME2xhbPbsPrRDa3JW0DLZ/5M6cOzdg
gjWl66NSL3XfIKQGCJbGKNJmysNPG5EyUbQUJqxzzne94w63nS9QrhNAIe75
q4qTaN1+/dktxJWdzT6nc7DCy/qRFgLSTWnAqyMUyffjLypChbeVK70Z21nI
hiuL0t7pP1/QPjU+4KXkCVV+ieHCAFnqnaCk61s4DXCETQXiavjfeSjO4vUx
Z756XYBU1fi6UDtYhKOCtVu97YXg1M0XM1dMy+fIcHV2GhPCqyiLy2PsnSMV
Te83E8oBenZjk8/xsDEtpoy5qiH+/Y8pC3G9G6al3i0tNpg11fMr7WnYsxew
Nl4sBWUFTXPpg6Ar1np4c5LeZ7svWfDSuYhepd12mFqg8YChjq3iBb9xFfKa
V1CkW5nKUXl9ghUfDj7HHhFBqcuJM3PI2+rhX+tYeHDiWwun11YuGtdhXMeo
290JXhIxT/jn1t8LrfJ5CRhxZrpviJTbhrfDOkrkEOi9v1lqySMiMfxLATbq
S2A/WYKHOB1xMaVAUKVdPtxloxUNsdIm97nIssFf5Aubk7kGSV1l0ehlQ5QL
fHyk2dc2OYrvsSrHrNiQAHRI0NTCocP7nMvk+mJM9fUS3epAuD+NhxqV8xHP
hWf+iz0bUDTflsrooz3dEp4NPUf148et3+/uVhqboPNNU8xMHYZicODGrZJq
BEBoRMf8d51oTzxY59+X7/ee0fGyS5m+NRSPBoFV1bAwgVt0bNn9OKpMzsZH
1kiPYNsiYqOcMznqfw8mqxfn/qcHjGsoJJbHf8CgdntgQEfBp9RMXCNDx819
AL1DyD/DXfv7NCqxKOWW2pkDpvpGJH3O1zzKOgJohJkwTgcb9fvnyn4MpM0A
5LEH95r5IgGYOclK81dT2lEfeCp6ngZIvRmQBkwjdjMHd/0Q4m/HhQ2BZXCN
Y12Bh9nj6c2Du4bxbeN+zJj81VB1sP7fTFiYEpBBxq0zavUqdGaF+t3h1e+L
ZYLIuPbDl3Qy8ieqehhjEF+hHGsx8qoqXJxSaNMI9UR7IkO9FjrR1AL9vLEu
C5UjtSVvBi/Xb6ry/raWx8kP6vuAsj8MBd4IFevuAozl+oSPaGXyy3ltYPpm
tiVbqJAfL8H8fmQKsPkrx3i547oQe5IIDr3yqBxnfAZxWAitAU1IbqrQ9ZqE
YuXvUPZC5H1d2UG4hktG9XTfbqf1huvxwHFsXSHQmt/YXTFX90z0FCNPQCLB
74iN6KQbjYHY5sX53EJk4IdJbZR7dRojKfU3IPMs3Pku+1x583sd+OBzUBsn
n95SyR7urprr2a/2rdcQo4ibmzrKAD+uZeZMpwkKDJl2NPf3VezLOuwm18mD
ngC1UDVYWPLVok7IrPoW7d8kQ1dFNWLNd6aOH6UfRsIP7mQiownmqcG0g9ey
3Lwk7i3Tu/7Uz5wBLvaWyQwt+h2/B2CqDzq3CLiAyjcdJf65TYbIt9rXexAE
Z0JNAzyLmwD6qTx4dqcwzu6rnqkTuORmYQ2j0xL/NqdJdjJ9gKxCNGuCirH4
YrmlbDjQD9a+7zzwR1FP1yltlcoC7hEj18cjYMrLP1z+iZ32a/wa/igU1rj6
nuLzs8zdJ0CSH3kVhIY4IF7xxtpEl+G9zKFajlw2F4fhi6T1VEaUdm6nXu+p
5AZBAFBraQP6xajZ9Pj1eV0AL7sQqfQQ6KXVe1uGMc0X+L7fRNOoqsGeCbb+
m2akFbtZYbJYnHc5oFJ9uKAmEuSf6CEFltyAwNYb5pz43DhHsHCqEZr8D2ov
4k4EuhgZnN9iS9PXJmRynNQqDyYA3Vi4BMh4wQi1coW9ukqUUufUh0+FgtYA
rC/9dPbnaO7prtqeIcHV3RGFQMPlEsgbLnR76NbEjoGiq9zlvsLgbQZ131go
mpGyP6LKZxG91B39V6FMfpGwoKJL+cS/wzK7BjlVL18BPuakO+PekOW3QyYP
pfq2dgHgOyXW7Wm2SRBFwMuT159juu/zWPZ6VMZMCRTYix0lPzoqPVfP1JdJ
0EEfx5Z5GJYnmg/8sGDjsYTe7xMW29eA/hkz8h3qk252IpVd2WR/McNVT4ls
Jn0xGUfG4NZaLFAXY39H+dDAx9RGrvloyUcWCcQGCn+87hCLGvKdPsnBt1Mc
f/rLqPSAep51DNW+PheeIOBLi1lywYEAgQoXZOrKcVjTi14w7NjZ2XnDc5SZ
+4rEFRfYLUFgRWLwJm4mg4xM4N2AwZgFFGXVw25VTn7qYPKl4pwnraRuTAjH
c2qHr0cKqPNdQgbR4rbN1Qi4wQeiWa9bFuWJ1eS5XE2m2gdFDaOtngMMwKdU
Nfjit6RY/yH0CxKyP69kgowN/3mrEdXkAOg52hxLgOEGBrXJrBW99F8/HNPf
qavqAR3deCijQdKbYva5PpQpeJ4E7Y/Je7Oc9iL4caIXcHZ/a9sZlq31v4KP
ka3DPqZOmBMBQ11+RGx4D9kneWyR1ucvybfoVm0WD/v5U7fzT0Yxf5Mlb0Mq
5GDJ8ThgTeKcx1L1TvCoJiiYrIsKpMWV1WOeWWL9GoFr4Jl/avxUOwfq1QV+
K9X+HMDSGMKF9/Pp88uDkDFVqcdL8dwKzONn5Xi8eBbUCJ7PT8VfcV1EZkIv
s8dd3uEWog2EzBqL7ffpfySz3sTR1mEtDmYWQJIvlOTgjS3Je44U3Ob6WXLk
uPFMjkZiVyUIMlbWrZhdzgGxwL25M5nnEGCHE2PWvAmpGCTsfvwV7JNPgvzI
IrFj9xsehYdEYuTR9iI76fPxxr3eHqK2jAUf6JtZvYKXI6jspJ3RPVgRzhC5
X1FvWIPFWXyKF2BcXbOi/SQr721RoeGlqHKhzX0BwkUX9jIME1r/X+9Qx1pL
aoypTV++/llk3ljQQlP/oXEO+9ZcgYfT6kanQ/F/zVC/3QaToJc3dWbxJPKB
6gLBwJnQwzqU+PynWvEYc07k5dHazXF3oMwcz7cP1Ku+lKV8Cb2MypiHtKMi
JZ2DckTM72XICE+RwIOUIuAPM7t3Bqp8lVKCHCan5wRDA4Zr3g1ZAIPCvjpv
bGqXXXHA5Q3ipbU8pAe2XsGkqBAhwktkbKQF5+f3gjOEAFDrsIOT1p+iel+K
LzU1RSTkTiRyX3H9eMoEejCt3XCJcS0+edvZFPo1gSxiHYp8vRm9lIgd7xmB
3qXITssn1wZVTmgg21Qycx1yE5M0MrjHbGnINWpPh5uOvhwDpvMYGgul3v+4
vtkCI4FX+mh51RGk7neHQdPljiGIlVfKV7fx6V3m1nNQNyjME2LNRea5BC0J
5tjhk76HMa3Rk8uFQ+sxPH9C6hC/TnVFv+vsyrBddohgXbVWIfgvf6nVknco
ruDtuAj25WHkVh1xH2C2i/VpQXb3kb2ZR1T0LQe6T+GPYDZkfvlDe6vSd/1e
fWDbJR+2nBlJ6bXG6mAM+j1zVHIS/ZqpWm0pIIFNgOGUZKFuX2JcJtcp1MBW
Xz7lauKZuPjR2CVJfJw6vmLj0mB11LXEDMHI/wBGkHNjDa0Wax9oktKF9qgA
lEHbQEBB3rzMVmOXy3f7ApnuVGtOBQ7/WeL5DEQEOWOnRaR+w5JOgxngcgSu
8b4xr13j4BNq5Dl5ZxDKSAKlmqNcexfv8ZFxUsQkQ3VT4thBJnwCpKP8N6bw
SW/7YsNZ5bnSpgMOMJWmpq2uH+JFUukhxQL+kwCzxQTLZnjtqMW1ujfh/zBc
p8T/tmH47DJ1XicPV+/4WxDWy07PEzMYZyzKKL0ejEAuZ9VI7nE5RcR8Xhni
bC54a0IuH1ZpGTy4DW43amanQGr1+cBX2OUTPy36TYl48cGZYRnTfJZIHMkS
43TD+SYiH9Bfr63JQkjqsf2t1P/RI+lhrDVxQfmsIpWcFwA34Y2BzjNDHPak
6fd3kUaDvLdteU+xjYIdU7VVaQIaQAXmWv00xcf/kmtzAyWqawqTHB8JhSXF
boQvhM15gXPVfaAhEhswy8wqrpmCg1n2peiKbPTVA09zbkvAphN1ZQazRchw
qIff7IVpDG5UBZAd32O5r9/da5wdMW6lPLVYs5aiZxOm6WPUmSr13OIab7iJ
YEOpTSDN7NQhXez8YPT00YoDkvf9XE5ceCUDYIYZ+u2zIg/FJNmmnadcCuEb
9tVfmgEyURZXKb28L2SxmneUfNLScwI7R88mvD2BpFQbaRj0im1zMysng/7a
Rs2XnwarHJtZR1D9CGaSx3W4paFk3Jp7mPb/uVymEnEiLfd6PJX4sBU5oirO
NxHl3XRbRj60YWeF6j33uRrXEP8jV7EgxNAQ8VSZ0vcR2/g6At0/6cLJGeER
XNj9wmj8IEkRiRVKFQcvS0J3LE9huWI82IaQhDJUl3kXU4U1Uy469gHg7pjg
sDyMrRC0Un1StKqq71kMMNDG/ryU2ckcFJ1DmR0AChMotCqtAhX9S5b0SJCX
J5rP5nrP5PeN0CBTntqyP7tva1YGrITrU9lcfJ1CasBb3fj7t7SARZp8J7q7
rHerQEoC737sm3ertPHjZqzixZKR3xBQvd2tWPg3tUag1j4Us7lvCFTnaNw4
6pE566vM1dm6lS7BDTlxHsnFdqt4WSQSL6roihdlJou2GScqRTGoNt85sZD6
8H0FAU7QatVJRuit54gFOORHJQjJfYYroeGprfy6pHz5GSwIydACQmBsK2D4
ZCSlUCPFDRHgsw/cAcEimLRyyyOpITpMpkFm0AfrqCtpZ8TU2aAiZW42w5wU
XhD+/zWL8rW5HV/9+4ymgtclbmMZpv9n0KB25r9V7+/MMEzx9tSY4xoM+AGu
rKtccN5GoDwzdy+ju6XeEF4+QxsbSQ8BISHBLliZSH1RjypyppgYsZiuwHkH
eJQAZA/6tAfi6TSa1qfoF8vVYqweGBSQk8b/KSZit9MLqghZ/Mp3PK653av/
/AgSOrlRQODHTfYTjd4quSsLpC+pPdaRKknxwJcffY3OJ75C6LYe5HZZFjLz
rLev2YXljxbF9QbfhQegG9+X/WNfn5cRAUntaOwjSyFqZ+d6glOV0PVgckVA
deFNuTqy65BB5EYxEXUcNjPNMbKEpHzKHGAwmjfmcvDYsp6oNLapoSpqcUTm
2a02M2bgYv2fxcCy1MolK2hy+AXYfFMiYPszjvyfAiZCnVRz8FJyenqKKPeQ
Q2aDBc04b8FfQSgEF2O8glMGcUP7sjLG9Q8JJI9jl/E736lijOZaPurqLHdS
N8KgSV611dTXRF1sy2khEOwtibPOcaMzyzw27kIaAwptyYeq+2IUjdZFro3S
zjq5dFRDumXchFXog0qf+fiPY9RjITwL5hXFkJ1ZGKjfVSrN5MKN5ENkOWNf
9gpV65ZtWO3BpRanLT3gOlDGiFxA7gdngAMMWMOnKk5+LSJGBZwJSqhq2Esc
pmIGGvYmHxlPBPyiSARDGCIntmQqOuxrdN5i9wxEb6XyPXypv4YkBxnkR/+A
Fs08tpwUk5gNGZjmOjElGOFo5WGx7xZb5kY/AzlCeq3rvRuMVy4yckFJM87e
GeJilYHoX80lsZL4EzIfQW8KMe4ovgSUbRKPMWJfkrme/PG2htu0EmTN2wxz
Pel6K3USs62893t9MFd6bBOZYeDmWebInar+Ogb/CJ4jFT51xTwoG5Y1vAvN
Ssj4yWcx0iskajcw0rP7L5/cRLQw7UeYLwvN8tLOD62H+6vKZmgn8MsWBQMZ
hY4K5gJ2hTsM0sA1FY0oexGfWFW9HJ7XzRNUPooCiCNmU2KhCJWnmMurgavt
O2HuRPLHn6Yn3RQGAkM+SYGa0oU2YffxpYau1vO9GtR3cIRDbOu2kvFDF5Lh
sWh9CedKpq/hCZfCTTA/ia8ZRhEq+3kuHTQzHHiaOoQAwBedAHzIBVhUvhui
hIyeSJWBkiQRNt83TDXgIuIlKguxGjntMmBNMPp9VgXOariPXeIJTaGePs0e
8L75U6wZ0u39uWlPcrACwuO/ph1H/dFrRQM9Y2BQCBPlN6BByyWkucKE3dEI
vI3NpwDiDnYRpWy+rv2zw2wu8Ms8MYV9d25v5Gt/9Ky5/foh4S7jtxi8MhZy
i55rnT5+iNbpplFl/+Dl8zsK/Y/KHASXvTZWa6b0yJkT3G8hI6SZxU5xTp9N
Xy93CYaPtaAJGQQc39tgUZI/gEA6s4xFvvArlR/gs+MHb+s6dT3WCrjthd9E
X3PooMm7kX7knQaIfFU8C0+grSocDJq8xJkmrfuDD95UP4PV6BcF9oaevueD
w9mGe7xwcVjlcyHXBFKjYHdYs6+knzWyL6Z642tyxLtGe3AMe+abaQ0ryoR5
Lm4BmyAnPEMFQXuWlGU91iOhiPqan1sYygugJgxFBqolwTGgcQQWtsUxua9f
H0Q86PtFXrhP63jn0RwmTA4p+gFooAiNdgiv1yMgStmCCu3gpnW8YTukmtLL
Yp0Qop+kriCt27mYguIcGRS93bHWt5Fz9Wetk8eHJ/zxsFznB8D+OLG2mUvx
D2rCAXDjiJngHTmvSisXTVjzEy0xdgvX5lrK7AThEYna1VNUv78xAz4n542Y
1uZiXBO1MpalB5rFmj3A/XWTEwOw+5aRsyelVvHsv1K5x489VawYP12EFwZv
w4kMdokDMLBgDtbYJQIMFOo03X6woGRWmSvhY/YUcxjYYOZ5Nxnww6p2i/3x
y9HkVxVykkkWWNHb55OPONTQ4P6uR4iPuPMUbugg4UxEX188Z1w9pLP6riDl
+QbXIS4fF6jKTZ+eqB9vsK+WJNWBWJpQipRpMiPOT3LTElUpbDZ8Y7O2UpH6
kjN9jZP0yW8dHoGcpzfr3j42ztE32raE8b5ddn7XEPytMza8Je0cLC3NZH/O
vH+GzLQz5OCWL2inC394koXoMyKEGfi6JT5LabSQK6eV16QyLpHWjClOS7n6
uH2DQr1iFjvobeoJOYmu2E+Gg+nAkZJBMBHSyD1WuVaW9YNC/+QYHDx/ytNw
4LmcoTNv2uZx6QfdcrIjZPypqLQWNPV3QUEMFoZ+brXiB7NrKgmoLKLGLCLF
qMqL+hETo20gq2qzc7DLt0P5O1SlrrgW/hd8Bx3ysD7demyabiGNHQepWO4H
TW1gMUZqd5BsvNz8XBSktw1GTc9Nw+8i+Ty+LOA86yifM9YV6E8TPbYWpEVz
hl06eLvmoZ2xij8BCoBLw8JykfzdTCxAJNnktFSATx8/E4H7paeLt7sPNTAC
gDaMX1O/o1XNtt4O8Ddlf+3Bfy+SLJ0vSQ5rdZVLAgkfBs5XiVCMfjspieiX
QRZbvZBP4YEeLejwXvRVuU4GwJMV+VKsHB5lijqwpNjL/Q8LeT8NYSO+LgYn
p/15V7gY2HirdGtnBD5NiR5S99TtGzSj6OxqmKK8J1+cM/eGTkMS+crDhjbl
sKF840vuy/n85ANpVkOyYuMa5SIGRv5qF1vk1AQ4k5T3EbtaS8kb3FysEVv1
4GCU4V0ZYRCONTlMSvhmHeVFv8ChH141nP1bPlVQF5LrXfAnzpLRP9xTOAU3
10UlhfV0eF/ka2oGoxQvATCPB5HU+MMpDllQ2dmxaPiIdq6Op495DFsQJcSQ
VOmgzIILpPD9hr2ZY7DKiGmemyEr62rNFmNYUfMvNEAnk32EIqmIC1nQqnh7
cmwYyV1HUS0vgbRk10StT7PHxSLrO0ne9YfdSXbcFyX4LXDZbg13ztpbM0E5
ONkwcKJIqQX4RNVUWXgoP//rlX6wDPZb6jSePNLk7Z+AUoYCmaFQRkG7LSe+
anW+E9OWS7QH3gBWsWdTLbZPC8btGPvbMifSNhKS0jCxiNKy222u+yvFf1BV
O0HKGGRIR3uAgEBuAscXefUon6WRqzBi/CDRQ2RHU5lzrtqX141+zC7Jk7vB
+EcW6Kx2c3IK9IQS4xPirwDFcqLeOtg/MfLvtMQYqLcv/1snF1JdOx3ryx33
SH4Nf9bcFyTBreBrBkaXkzr+Yw0eOF2mRc7RsDXABLQbcWs/FQcMvn7vIFUl
AbXqdiqWReVEfp09Q5YCurCRttGm0A2VzoIIs3EXQRss156izwpV2mk41Zou
hFtGwo1zO2yg9bnbjoqsJ1Ahg8kiCheinSjDh7eE4JUqNZv3ef9nVSxgfEcZ
O2gUUVowkBdNLJRexOn5JTe+GX6mCxTlneo46yx74x0IcpsLgRcyEEhFqrN+
ihEKzJK818MqnXm0VCvWU5i63yinHj0wxtpRrdoSZW7cIKl6i5v5j+9wFOz4
SJ7StNQcJxzeMKl6mpZJuahH9820XePnTwiI8SYb7yWSs+9fyQGE7GYMPxsk
EgXgw75uV0c0swYukWDQe9jh+J07XX8xCl1PNaVZ4jl6TEbV2dXpYxOpojDW
aahpk6XDlwLL4f3KaeX0nv2v4aypvk2xhkyXPC9FoLhzBhfQSLSVPy5BoNco
icBRhk8Gdn9hbDBnixHkG/okPeEz3NgMTBGWBQv1K/4Nnzs7zPH0/umdlmda
WlT6vgvNlpASdcAwgomOH4x0naYqavz22ReIquK6w+/ligU1thS9xBDDjPsG
7Vg8Dwi+IkgBnUKQgyGWCMvgM/lLjPyVCh/2J5Dk6PHH6SMqdc7wUn3Gmb8o
030VzGvPq+GFlSlELXkPqhyviInc3bf3tCEi4hK1A9dOJwJ6rff33s3QANPZ
mm3wX8hPo3fvqfU92LWbJpvG9gYYMVoZhmnMpW3EcbqoVJpHkuRds0Ua99L6
7iMouwynX6tZT0tzkGe+yh1RN+GVIImwEKZ4r7vxptPdL087P/EeQsnEeiCj
wP7oOcFLUiur2FnmSQ/w/YDZbyTnVEKRqp5/g+tOkSmd10F44fHUdiw8HkDd
A6AnsgIHhMl7SrrS4FqLu5X1bieKIqFKxad9Lk+orO3GKxSq+g7+4wKO/JWt
Sc7mC2Jmm2uLURVYZ3Jf7obKpVZ4SdZysZmqC6eleDV4pdKFAQXADpt0VTUV
TTwJzUiGNFlkJTPRIg9+rGS8wsDS2mCedRei8zNMNdX55CyTxvvjmZUPm4az
NhGMmaJ6mY5KAnyy3zgaYqkC2/iO1loQ4n5UbL621jQY407FZ5Fxq+r+MrGj
l1uJa0xTHb+owlfqNMV2LGTM9XUkeB8yTTjBVTiwgLziAXtVqcSIGanBdpBn
GNRXZAuWlfZeBj845Ye5hV2RJ4H/UzSWeI+xOoyRrAqkw1KSdXn7BuJlsBFo
AhYPtIvxUTw7A7nUjIjVT6y5wIuJJzwVYrnBwbF0Jhd8nStqy+p/ET9fdMIU
vbmZbTzuetb/qSa4/zJkUQuUm/9Pm46zVMSX3WqZmRkOZEdhl5nzghDA5cbi
zkBZXCjVTeeaJMNBGuTk1yGErlxVe42Ile/LIGg8Cgtqircl686QDRSX9ajb
GZ5JI1oJUMpsL4oSAx3hr3NTKhECJr9TX38AVSbDDqm6HOFP6psc+hk8TSir
j77IIrH+weaRZOjfkkzodAMiX/zg/rHX1NJEOZX4uFzwYfL1jmqKDYL/YQ5U
SCJzHpOmciANLIlBQmGHK5SoZHrrWy9Dgt/O+9xSdN79CT8ffIc/4luK1zG4
IlVw7hTvu8TGDVAcoE635ZQ1WqwOGNKFCg/9/qzRTAACnGudMkzzeEzkFcrH
sCLhn/2ObTcQFIW0G8dT81feSZZr8FqRkrXkHfvsj854EyeX5xbLDclL9aAt
UubMn3mWCoef+7YfdhOWh0Z1nCiuUp+Cf47jWDQrEbzcL4oJsHBRWOWZzFEi
m+JQx8IYdfWhLR3fNJZ7ZX0YmZ71DbeFjVI5mLeSfohpO8WlpKdNKoOC4Q87
VG9KuDqguTs8i7Z6CRXUJJtqoL8Cja+M4LiTri3A7RRUNe6KJTybGIa08k9M
ymIQUV515mZ9tDr7h2C1QkN38w7zOkZRAcud3eGk+nmADEOkebc7uayURZyY
H/rV3tKlF2hS9ZUTCIqdddZeaoOn1yzn84w+p+veo38hx6vax0r1Oa6HqqnI
A7qfEeniTlEi5SniXUV1QJ9+Ow4EexC0CqmN4jlZGKiylH+mx8Qr9ADjAHu0
9h2WuRfnrb0oKo9PJIZ1VlMPlr5Lu2aGOakWZ5Nms+zxrdRHV2AriuGMKG7j
gYEInQO/JkJJ2tyaepnXj44tVB44VL78HZHncYbLed4empRi1g2UinHq2W8i
s3JlGW9JZZiafC9i0wLoo3bXAdSQJb2nLKcuCHbwF4YgzuuA2jk/NyK8BdXj
eq9RzEW2xuW0BixrumhT8aghVfB1Y3bPplp3Jeiz8DXVTy2gnr6O4D/9h3p3
yoQrZZJGPJ8c0Sp03EJ65Mm1bgZesZmOHguoFB111aebH/1q/TAQwlUZLcQ9
UKeDl0NoQTuM+o4NiCFqk54ajTITrI22treGXP07ntCQg6mwzac+MAxGf2GX
2evg9+Wt6kuCsvyWRWyDA2SNsJFeIFJTZvROwpwyRCW3YCma+XtFUqgfGrIM
4vr7w29bshbtM3zUi6IonNSR90n3wgZ37c3b6ch7dQFeC5IaC0TaW9Qr+H1w
53NBbCJiDVF6ddZoi4mpqTApVylygSvzpi6LsT1lXIVWjk41d31lHLhObO0a
FoRZA1UmxEvpxLa5OC8LOun/ssGyjkcoeXsXX1cc80+XFy+nxWajgl9CPPpH
wgsjXEkfUMTSf1Bu3ezNV/DFisVdfJ9qQIOyMy+hr5kwweYyFsZb4gMmbMcf
U9wD8S/j+SaJEp5wHUiFdULoP6m3dmyzUDG5qr76Y4mTb6wo/H+7dMD2pd9e
Smpt5Pnc9GWbhSDDWNPAkTLOjh9Tt5hAMCuJa6Gl3M76UtpUAxnfBZyw2y6d
0olcLwUuYt5nVSRQ7jY7DfNJEvVJzFVxzLeYdnb74faWC2Dqd+khAdVi5SQs
xo126SD8smI/ilsIrrkcdYMK+UhPB+zgmTE1qKFCrsT+Jp+K6DNlpeoGa93I
NzD4mBg7H10uDSHqd1NeXT5OvbELftM77abDY3RPtKGtko1xrT1aSB+XJ9jy
I9H/rmHbG80/lezyvn7dF0bxqXSQtlG18OgIy4waeCZH1m2MDr6nRhOu/lBu
Peb9Ifupts5AxD8SFMOuI4xXxOqB5u8z9bvJ8ulNBT8Qk7Yx3xB3St0xBboI
xjkjEJUrVGCDQt/el/eQeaiabjsHKfj2U8Vdc3LwA1I7ARXv8z8lIE5SRLOV
S64umO6kb5CrhEjCJGleZLB6icf9eWvH9hbD5hfwNt8hy88YIEJdtg5pDu86
Gm0zmAzAunoiqVIj2YEMqti8ARsluwcwWdwbR7DW9ZH+K8nMaCE8tva3/ReW
cgu7f9HDD8wm91Jr+iOKTpP6IdUA6sQPlVBrymKr0T4/NMjra7l95SlLspyy
bUakQpEc8rRAlLCozk4ZpSMM7hYRXhSsSRmVB3gK/88ykZV69Gks3xBw1Bsn
w8+LmENXoQaLJCMz5rdyYVIi0lNpxRnFuZB/NQ06oBPX/Sgyrbukwv/rDwNA
poXdbUXuZ+ESdAtw9OeyPJbrCFNmUNVBNRSDlq/PwIh41keneU5B8pPolyrY
X++YE71Q9Z7909+WWHHOax6DNhE2YwAts0kiAFo/7K9nJaPc7WYCFIJyyyDK
ldxz3wJsTYmWluiy3A67eDFj/wcTGmujwPO5sox2rKX6Ls4xNadGYWP+X+Mf
/AhSbPtBSpQ1tm39M47mejfBwLh39WLh1urQtlkbsgiVfPN3S7BIkIuSGqvY
Z1r1kqK4y+w0BrpXiI7etJJ0shDqaSKjv60j57/WYM6H295dJGOYUSc/JqSM
suwkcY3sdNyIgD51IfT/gQ4JzYDIcJjzDVzjgMNdDhWLoGrLxJJmyefLO8uv
DEAIvTTjXUFFWSxDEnpYu4VngQSIW6AY65wQIlNkW6YoUw14TOsdlFxzfof+
irPlLi/OkpxaCEJSJ/3c+Aip9hZxqEQ+SrEx4iE2mMLNugg+6fSCsPdGCSSN
VVxqtQkfFwq6RlQplozhrQCOX0hoCtX8TWXqD/MaaMUqnccEWKo5Fwu51W33
Hxp7DDSgaVctSr19H5e9AfnHuqSH6umktdDPBSzoaSlAZBTB+f7q+2V+1XDe
/jBTZfenzDnOhKEqXJlj3bqscK2rgTKu0Gb/Vi8h7JY6Km5SqZKu9GFzENzW
CX/Eo0Pc01PjWGXKXK7Dz/aVJCefjpSUHrF3CcjLcDR2uciK/nDPAGljgZhI
02sfLuc5p1fpi0TH/u5onRPX3sJ7JbC1MSuEMIc8VcUyRab/BDS/M/JxO1uF
Tid2qfjr7dGEMzJ3pj2dcVg5RZTHRQHXmZ2PTwGUhqDN7LJnDmsw72HaPsNO
L7hUmt+2jxBI3zmBJ+4nHmLPNmnuYJ3B4Nh/tPjYh5e1Qh9Bun+i4ty+Ohoq
ggsmrn7KxU3aIiXLZa6qPt6wU07fM1xKc94AUFWyMkal5DaQcTz31EqGa3kJ
ZXHJ5dXYYulkRFGPAe6biSkXBq8O6mDygbC/a28IzSvKXnHwmKvGZxXbRkqA
1/QTd+PzNxGs02WKNAoOYbevc1qKY+MomQDsjYTlBdICBpG5iMSGlkX1B4nr
9u3mLb7naazuvgOBdYAa758yjrZblJX8BDIoHZPdegnymDD3U/glODLvxK6I
XeValDc1S3VZi4DdpHMq8wN9qw+V+Q7HW2x1KkNz1nBFOoc5+HoLvau3846N
Cmw155op70VAp5P4joxLBQbCYwGoarmuPvk3y1F0vFnCJPK+MlBhiBG/rtEA
lOffCExe8xQ6PNa9eIhQrtsKUGlX6WenK0XrbY9XzjrbRK8rp3dNcD9WHRRa
IKwQkOYP1YtU+8K5JIdk6+t1BGAbwEDrslGUcywbE7xJJui2UQkWCoGVsw8K
FsOVGlouChIoe0QqrFNfX/y5RoNOJi/IEYPTxjOsqRuHE2wz4kYwickJ6xO4
C3kMp/demMQpZh+HvE3oB61ZDJiotHbO9PoUz6cOA/o3uYFjPu8PXu59wCh5
qyQUbHk7upAZq96ZK6UqsMUG9VudM/He2v7c6WlkbtYoGzYAJSFrfazvKC1B
JCbLydroZvWt5tWZ6DaMS8PsorOP9op52GN6JKha42+zB42k3xDkwvNq6NRt
oy++VEI4PBA4SATLVdoH7wqjDfP+7zhr2OM8vxfHBUzUx71oOtnBk0dw99Ux
LWJ1yheA54DZ3KKybsITvyOgPIpzZM3H3XYsoRLVp54y0S9lTLqUOJVzR8XI
N05efr0aAwAldYsaOKV5tfXWredCIbPsx3h39CkRwaWHrQw1bumcK89jY3J3
MYaBtrRHRVpJDKRNUAHeOPwgt3P3EB01AXbcC/ipjsd6Eup4s4UI+w1Qp/DG
sAKjByyzvER18/N342qwIWUxGCLgFkI5k27rT8jxoZ5tqn8AHD4LAAqau/Ha
EOYXMe6J+u5FlQRjF7RZocmPyzi4NCTG77HYBbpImJpQz9+BsR6PpQr77sz3
QLfkNoVIWne0IZqckHjQVYq63IbZhQi3fV9P/7j2IwLuZcP4ryCgk5tTNoUT
VZ5xjn0OKHK7/qDvSqdlD7c9Q0qCjJx4Hz1vuioCB/OVTma1SXM0Tr+oJqpB
H77s5flmCWon0+a3OXkTstBCD+IhrvGBVLHzNDwoN1Z5gq/o0PO6qDC/GbR7
d4TgukF2YV9bNoQ+Ywqg3jrfFzUO8S4IX8KkDCLT20oP+G3Bf3EJogZaGFtT
2JrRbbF1NesOj0RlY70JmEsbxKHE8VixlDjeYIVK16CuRkN2ALf/oyxqD5n4
rFiCRhJdvNAUrvT4TaJfduV4Ax6qlIfiaPa0R60uiZdRUAjNWNbVE6iHFvay
YeTfUkeJMqAdBNbKk48Qm1A+AZX/J0d8j1QTjI2B/c6LfFCa5vEdrhBqzYCA
OgnNuze+OsSc5HkXCtVHjRjultRV3I7gvMJ+rO5c1GEMugwemncOeckCowos
/Kk+fKwfJucwMBXev3jEMGkJG/xnTf1MxLOwYgC69+eqPNIftvDOsguQWFrU
56zaBRA62g21vQkcpqdCN0+4l3rFzgrfgLPQyExx0doUU+qvdY/H5h1gX4Yq
Yq1Ct0XYWh+sowDClXZOwy0CjCfknVHeHG6ITNtY0tDSXg2+lqtfhbpDgAKD
ZKy1DV9hYSGMeQOb4FFw2kJzYn5gZOChgDgqUENkWkhWF9JZVhaDO3nqay6a
tu21qn1TbTjoRFNcD5oASmmfeGX8Uq7zVxMaJ7i7ZZB3BsE+wjCUBBs5VMiw
hPALdE+82eJja5m6abdu8iQoM+w7GkDln2WQsp2x+EXLPkdwD++24AyrbysA
I6bgpiJLTTMXDTvCk2CYveUlfdrohKgIHpFBVM/0TUQ1mNvIXKXY12T/hebq
ztH+ChzwijJp71Rnr1o4HOk1t+GSNYfRWPW3HbhVLpJ/tLZnnkAnuLfOeM/H
yLgLvUv/EPuQh+eTfUtRFqy+FPxbrYLZAiqITnfWsBq2e9/DrcKlQ9iKkrGg
M6doxjRFwlDZYinJ2JLG+kTbtWlOIZ/OieXVbiQf92Af5OOT8wN+DhOYYIhh
blFCqIfmf6ZV6cV+gekjgCXbFHc6971mDJ0g5SHuPX/UPVFFRS8ivnLEEJTb
DvAFB3B8wOVY/4uyuD8LzuYNyGyUW9fMOapr+saBuE4JVUh+BzjQ6x7dW7OE
PpIwaOS8K6W7H/Clq4yOkQ5YdYrbcGJYi/lD04Ag4gpD8rTQBX392JoAndqK
dGK+HsZOnke/NQYhWZR1RDC3L/+JPsj8fVuQQQXt1PaybqtIbLANqx0M9uCu
GazCjWfdrR4qCyD/KOvZzA0njmZrDgCjzW7KL50WR8GZlnnfUun+P4NDsGZ/
S0l9ar+Cve6yy9+E2V+J38jIKUGIrYPGRtjCI2cgJsfoLPTOqAh3CpCkoDco
e/GlnDgNjYzBhjtncdR0sUsJmO10lD6xy8l1HEBHaJlujnh3avvWu3b034T2
xwiHnkF7LQ6Kd34k7RVVk5TrUY497m6XcZlvxvXJD0nq/HkjsBoKEhgP/zlQ
BMx0x5J8KJQ1BEEXo7fHK71tQUzFAQjwp/45WGzzy4tXRgpUZpBmtMpyyGeL
3i9LvmdGgXuUGxjQeSbpps8uYRiu7Kk4Qswb3hbTbL7QJnJd9tMw8GRx0L56
pRih2XcmPYizunwWYI31dMsy26cWR3oBQenEtGLelU73a4Ur4oQELsfZYwo7
vVI2yicYWkR22FKMiu+8Li+IMOP6pUjiYD7fCdwgB+O1/kukiqo6XQwTMlpf
+J4n1YnQzr3SVI+ifjccRgOxdWSIQYzumv78RkaaQUuJhllgNrmp1bx9rx/j
r4uYxWMeND47Ynm1Jg7HHpc93bhCV9tG2DSOjgDTTL+7bQBgMyCydpmspiny
DHuDKE/MyBGSxNHr1FWAo+EsMqPgKEgfiKK5nomf1d0a65398vkSdP1Nve5H
H6hZtO00xBiJuCgCyLTUDPLVaI24lh/W+O23IV2Z21WF1xD/47cYru0YB1Qh
8mO3qmo/pGZMsNvycwn7ygxigb8CyNaSjjJzAaqDcfvrywPcAHr2etnQqK6N
LHLo18Lbp9A1b9nSnh9bw0KJdn5CfDwjTl5aRnO/wcb2OGSBBJ9deX/aNTH7
M7A9PDPwf4id3yKcnov4jottjFqffdHP4q1obLeRr9WjvwyusmfD+bAjct46
0VpNUeIGvxHCbF0J8LkvMF7SidQNIEkmmCOjXTtJrp1NSP6GuLXpEQgwyKXC
1fB8l/QFoi2z+wbwcWK/QFB3sQ0EI3RqHrYBjDAxJFNi8e1J0GEqex//3ss8
+DTXjm8Gg4tefBF2g57lb7zZIt6eLQ15wy85L0Qv+3ESVmcHSgoHOUFi6xJt
cGLPjvyuGIdb4r1B6odEqeA2f93Oxsa75XagSmWjEFq++VwMy++wJYs12kQQ
oD1YDPmhPmR2sw8qL7kFPCip0ZUt/iXv2+TzeAHWjItb4Eq2Eh4fhe1sflGC
YEsn3fwvTRLogdsJm2Y9W95pK94qo8RN1A7s9VQiqhFd1uB/f8PO7Bf5JQPN
m3IIddWZj6RUht7AZqOGJSJ0fa7hT54NYcqXrZo4xkizqO6HvJSTK6ZjgIvX
FFUZNmyeSb8vmPG5CyuZ/KFKIN2K03qNnmEvoupAnzbt5PejmerOP6WmoiGQ
IwqUWtouRsn3BObYmkwVtfHSA4MF47JtEm636LfG1wKBJC1fbwiNPfB146qU
sWy5gLwOFCDBy6cEreenoLNCfUpSizkyFLUwZf/4OWs62AV6TTAhuCc+n+bR
6FiBAu96BsugvajZ/pFXr+cF7/LOXYTn7DDEDA2dUPwH9Aff892rJe5MTwVP
qtFwk5WIExUQeqzAOBoJ4o5M2jxvXzN67OXhz558gFDM/ZoZ1bn4TCSPrWiH
qeto6Wtag4dwWutNFuP2I683tUFKar9hdQvqTcdPn+UUlgyoEIMClbythuuf
NGiRnZOVEq1rrQD+L0Ho80lzInnQD/FiSulDYRN/Ym1Mgm5Tmi2Keu2DQBg8
sfcYBwI9D6ha/kHJ82UAhuU5P1Rvq54tNpZ7IGSeC2x2df6hK9reKUAtSVY9
pseAobhjROL+7qRRTbR4RiExNIv1QR62o6cZffAm4wHp+bHt/6UmgVCyAKoV
LKZjZFsMiH89Q/NNH8hbNojiE+QV0yKMQErQhdIDL0gt+npUv6FewZ8sjl2K
aqPLSZ4+GFQN4UkR8ctr0sRnYE9ErlRoY+NKEiQMqtGdK1hp/+eZT7MBD7XX
ZkrOPeBzOzf3oCjYItdhCyK223WOKqzajSKwzXRgpuKfjM+zNvD/47lMOuPL
NNg24TB0wyHi1MuMGjKIDN+/9d2Bn4BcfxySwECwk/LUyNckiMq/psgH1Bie
AoAVUrunq7ccZ64YG4QSyt0YO7/mGNUWWxJ3G2EiRZ/Q5tuP4MlQpwiqcb0i
fcbsz1NFhIANi5PZhF2/7Bj0mkJmVJkuxi6rh9FnsUOPqM6R7tTf7OSwpa2K
n+FCsDnmgGuzwTQKxnrdcE/kTDClWHlglpiyPJayXvX/+miMajLaRns5zzZY
21n5+CeDrPXvUB8ghE+WM+URxRYBN+XQ09GOQTAFn9PMRmpRX4s+Lk1nro0B
yFKAoL/kmn+w6SeEMuXGWCelSyUQLZ9FGx/V+/PHN5Azjd66xvdW1zUCFkJQ
9/IT0nNRyneMwI1Z5liM+RqwkbXjk7ExrUceIQiX7+q7zgGrNKFf/EZhIjbn
LJGCVazSsyBFW34QoBMsjkdMPUIGXGkvH7C/jgScK55/OuMoSuB2LCS55Hqx
AWBQom/EsKa2rc4XpAj+i6FMXLgcZTF58hjpcmEDNhyOvYAL7Auu4WBE/BY0
fVuFDPuipPotyyxqMz5nfDq1fUp32HbWm/53Ej/8oyHggoCzcNZEf1kg5SpL
u3/DoHBkmoK1+saU+6tJW8ls+2rruuIMjyOf0PtJvE/JAJM3EYJ4IVtTpjCs
qx9Bq9DvCZ82Q1dIKB3EmuX3JeH8rHCM4KIOICCiykWHN9Du31jeqq6qwKJx
rzsdRKvZSHTG8xd6LV4SaBhC+1pi6vS1lrzQGODnS6g0Ivpec4qAyMamE0Zz
EXFOKkO0G5fXLAzyPzvQq29BHHRVZBns032jYwIrMB9unbyO/UlEzfqr654J
IOGP1YiLqOchEQADbjeSJQJ8kNfs/GCCa9A6HpKslZalswbZyC6dAW6DfaGB
YNtDGF6dCCdsO7jAgnxGJjBxxRSo7dI3fZFvHMzXOxjwWnHlvSekCjW/ARjX
PUsiioaV0M38v2YqqQJ0CzZZyQgr45j4yf0AtDRrwFkFZeRsYdbpXY+Qy5Tp
wO6gxKhDJYrh2lTo+Vt5LgfYbzyhqaq/kRnPOEQvvyldh9z6D2/9UhZ3df8b
SO5vKhRh40m6dqNKgpSPCVzW0p+TkC24a/DT4yaH1fM9Nq+Of4nGLAjcSA68
l7XvJsYQpfKaOO7QbP5OHe6oNtTbHp+QWiAi941ZDhIEs0c0kPoBLxGbuf37
HsDGZ0L6yTXwgwpGmn26iob2k92s65imq6XPXLj8NLLuhZyixwiRVPw+sIrq
mYgVEbI0LtF8Pi0hLYe96nX41FX0VSy8tDaw0eVKh9SFzWJhualhqlupKYEe
/3rtQU4U/5aev4t+e/DsLISw/8Hz0VcfSIij/5ZnHIDEzKPei9z56yRn43wF
4ZFHkwzde3MQGCesY54WwZ7tzaC4liWrY3vjRllZAMlJJFoQV2l6Ut1zCUJm
Dq/3JCrRiTj7vwhJRPfJ2po489aWw5mqnEikCaIOyqS+BflmvpzA4D2hHfi0
ugTR8UVGriTtG6l6ZhF/6pgX873DpJhxjEtmHbSNaWQu5/+geAwJA/qnEZ2M
TBgjRJXyys6hG4XQqppVM64qOqyhAPuRrdJ4CD2TjQ+76DjhsPVdKInNlAxr
F8H6mbwr134EbHiDCS5polAQY9ao7t6P7VGTbg6uIoFJQdf2gQBOKfK8brKz
khCRD4JVN8b5WC347daz5t70S+TiKmjOUZlKNjssZBAdzPqKuN9vXwH6F3bq
H6WOpcnl3V2RtRviJONgbT8sEccEfU41WfHvbvu+zqNFquRLCP6QB9dJrMrc
AyXZQlZ3rt1ldcIIP8XxPTUTKTVN+yGhnNe/xmJzZVpREhCzbLS9R2GgxA/A
Ps26J8cU+UqRGkBuhWX17iZ88JtfHb1SoCV4kaVgPKFj3R63LjhdEDSGA7fD
sC0+39LOMU1ft4YnIvl6PchyZTHypdeU0S7IEKG7tNFLN4q68a4YLSg0qzdJ
Bn4a48XLWKaRYyR2IixRc94+c8p/g8fSow+b1fcUn1ypmv6VkQ2rlO2kwMEo
odC0pzvTZwsY72Mon7X0K1S73kEcEk8Rv6QFBH1t4mri3px2zP6t24RFNAyT
9Ee6+w2MPmEQMfU1LMdKrTt+X7lAeQiAnzrWqCtMu/cPEDPS9OUH2VB+wDDJ
oRijVIXU5Mb/Bb2OMPKr1xPZyAS6QazFxjbi+t8lvIOzeecT7W2OyDj18bDt
Ud7Q/hjdXXiyaj5evGM3ZFdYYhUPqEEM9jIPBE7oPEN8vglNWxBO6F+0StAh
NAFapkX3KNG8Ord7xthiiFHcagJaOdqexLXSuy/QeH0iYczvFH5Kebl1sWnn
GHPz/rPVJfb50sybjxuqDM7m0//6hxeCQInh0lp2JevCIFX+ecn1ZvFR3UEO
M1uxcIpbFjyEffskhrl+2CMEA4NEWvy6G6DVmog+Ig+bd7OsD/gwnuINv9u9
JriuQYhnz90c4eyb5MC4fznK1jL0WzpE1qZNwv8M0AOPDSi6xMqMyqO1Qi4T
qCCb/CyIGvnF0v3D8pzHsLJWlho2RZ8Gem7lSKHueTH22tRqThgNxfnLvHbP
nOOuwWyhoypgLVd/ZGqn7PJjZ5V1TMNJkvtkmsq1hEljTy7ZxmuaU1A/P8cG
PC9okS+k8B2xlkrKvblZaQecggRa/35/eEwkJHiJywO2Oh2zGkTcpJC7FDez
vb5IPzdQwtCE/XwS2acoTjUR+cOYgx/G50qO1pdnJkYuKnl6livBBbuiAMi0
yFWz18790w/oWISv5z5QCq6Y/oAkLbXo8auFxUfArOwl5D0BqO4F30I1KOi7
weEg0A+IDnKOq7uIaFjzKsMVWx7kahOAS5YhTtTXsytRrRftpWrnrLP8Vjjg
AInZtkgj+ghvGESLkgxXzHTFwrKg4nn1eWHcxl0D79ih4611iuhd9Hb40FnV
/tt4HhCt3GAd7FRRCc5MaMkTBCgoZ63cIPLs42Zkjpxx5LA3YK1ksbHtlsOg
OGTgqb857hJNxdqLMVIg1Fzj303VGyLyKqYPxPVq9bzZz0NjkmhSXmajrVbp
WR9KaRIbhFOQJeVG0PhtNFaZEN7BHHzRP3akJ5GKyi/hrfnFwOXzMg5x+CgJ
eM2TXPSRBMqOYnyH6IdgH21dS5C3Dz8V3NxGE1HYlunQEsyk5Cv+D+ahuGI9
mJTOJi9VOnFLnQBu+yV5/88/JifWvRlu7HTeoCjH2QEdx0Or5P6f19/OLVXj
/43/2roYE4Vi4/Qdz8jxxNTzbwDWP5l9tECLo0CMkCjIi/GQvPh2lbaaabBF
avWny4hTexgAFdnDJLuTVDzL+Iq/SHPTCNiNz7ZKkvTD9ORJ5UmEfGJlZH49
9zNck04/VqWZoQZWQD3sd+p96/ap16K1dddcWltGQgi8XM9uC9le+TR+CbMH
EcJnxVSy1ZarxtlbajMTfqTvLbFsvBSmb1e6biTCzw5Eem2jdZLlUkPy3IH7
aRFzo9/UA/Ln03f5oG+TEfzPS4H4NSIfT4ZuPHzT0pldNm1bKKgfkU9ZQlHI
zJvuciEd/6GhsPsXb4Sj3KT0kv/mvuygdfcHsIEGM0ZkGT0dzx4IXPBAT6R5
/OUI6M1Usuv8ihzh84kJ2QqDy1AQwdRdiDhgvPWPL8KImei9KrpbYZDJngcJ
GGNDAXzRKwOuwnNZgRflFk5bBnz8QIUmUHz5sfkliFApgcyXkkmFhxudmPdn
P6XPbLeB0d4uGR5sLi9gwg0xn0oKwz4yB0R5CIqLp+jM2krUW2CAmE/YoHRO
sDnb/4ECR6lA5YX4OTxIthubBq0mayje6jx6jmcV4TrQm1gKB20RSNKy6Fyx
tEQz9IoaOo/4ZmEpjtK/9MnHIud15TBOfLNIBLooPm9uVILIB/7gjcEOvXBp
BZeQQYZ/XeVHUaF4Ss3sXc5GX+uN342i6Dt2Ict+9WQBUQjfH6ZwS1C97Q+F
E7mMFsyMJ8M4ErLmppGoiwYNBhAa2S73TYnOnVCx/nsBgjeNjO+ka6E0tZdu
HKjqkPy/ZWr7A+IzoAKdgl5NoMoJ8ihmz1HuCFjzTCoNgIz9/RN3zFPktGkd
NU5fxrrFbL/n/q/pvARG4ZWkY8W/qDqHe6E0eevzr5W2mAA8cw9jPYFjlZx7
0Qb4cDAMwI1f2lZBEKfQR1W232lJ3icHj8Ufju/StEEYpTSeXpiCG/HZAkHA
YwSUXzfcZvMU4AXbIpxHDCEFVbUCR4gzrumAsYoqPLN/uLrmB/P8hN9cz1sG
RfZvzVTFiMSyVbVjIqT0W12UcNvd1YliRv0HZ+L/0uKrVuunr8DMIAoZSgY7
DewnSJuOtLikHdqdPZw3OWOC24jjfjN9bWmVVjWSPOvvyk3tu2xzDyYb9Da6
jnTkT0n2EEut5IHb24ucdHzxXRBlYG5tetdc0QoltJqo6RuizXH/2EQqDzLk
LG+4NhtabkuHm6hAA/gr03jkckhU/yJGRnGQ7A45z7bJbVgZUSG+x8nySETx
G+vQVNJ/MvUeT4bwmCRPs+lkdzvafc09JnV4FSwYqTl4oCX5Y2XVR82mTiNx
8fLP4KLXu0CzAZKW2VwVDsdbJrSMeNSgJJ8hV6L0f2Rvv3MMkPM3wEPQBaOU
JrJ/xkjSQC4wx2PlP5qp+qPawkBGdjC3r2k18qEFKplD3gl10BVAkzeio9+3
Xqw7/s0IYUBlQ6hkGdOWh3sxnsuKMRWcRFN7I1e/k6mbkhT4Ip09uqbTzQZg
gnX8E7ImtJAmgsAotrjrTWvVi6k31nqPqwx49btrn6ffR2IqEUh2P6iKnK/T
rymfZWhxOKVrd+8k2EfwPLrwSn9SzPeR62ODFD362SAmQRNseJPUWAKw8Ga3
8a0/Y4bzdv0Zn3zF4UdCTxhBC/FzZNaEwnqNO1V4BSGmX3LMR0AdzlxiKJdn
JeqYIY+0euMMRneg1XubHUwoojHfHLTHdfVR0Y8v/wYnQzHDgTUaDyowfpHA
Y2LJlSyhiZysmjOLks3L/GEDFvXyqQBIferUgt+M03RKCBWUM1yPflZAGq1H
I3NFPb4HfTwrfUx4HMKpIQFsefd5Kuu6rKg5UYyJXvRgBct/CwnlfZWyvt5P
lz0FUKuWZ1g5/Rj57TibVi90icWzNAlj1AtdpfzBe1tjkcicSESYrdva5Cjb
pJNtN5Kel/va+rwS0mMCg420UEo40AemRPDLGumKuid2v75qkteOm0mfUVj2
a6MN6VRj03/vd6C7WfEchyRBUJdZrlOkc23m4zykNqx1lRNtz417hgjtwSS3
7/H29/4L7966499KDag8LcCbpoxUoT8/cHpn/emvA82sESzehT8riLtwQS+e
MxIjxipmL4UIzmUnhhhmq6VhuHD0TPwpfHpiarkajJVKrnB34UzNoaUDpr2x
NhPQe+PXutnTFtbwfM4s2oGxt/ZrS7jtkaZDCsqyOYLRxj0SbMuNmQXlGzmm
GpwCOxBNSm9oRfcu5kODrqv1c6aMk5bGb2NFTxOHWhUuDVDL+FvgiuD6tzcY
JotgOJo6WhB9fObpcUyuiSIzQwMe/neDcOSiGm/NJQe+Ch8ogFXv62dI4HlJ
U33/k8fS6kjR1JmN0RMJYeX0OPDIexzuTanhNdZMuCcdbYB6KPMOZRaLTv/0
KX4ijnonRhCTx4Nm0uO6lAAoXth1Te4/TvWPReS3ZF3wh1z1j8HGLT+PmH9k
LINOt+pydxgXDhfdtwDQUFJSHHrO2kVhS9zK5V0rF5mSZsMbhJgxvNrrOxpY
Ur06f+kXn6UbWrobO6pRQeIWijYR86jjP+cFxlVka+L6CRriwZAxkEhcdIon
IRYbRXavyb2XvDSwrdhXtb3v3YdzPRsjIrKpisM/To6I6U6iv+aN9lc7GQQs
6IfMnIGuIDA2A6RyWUayPbxTVDbfw6cnkXXbO2imscHGH/oyYgg+NZcI82eV
MRBbKJbuDXXVgzpDKp9QKY7scWXHyNE+55M1Q1i+r7h8PBn33hYIExQkpMvr
lOZGx+cAxgNp3a+u+kubbzzAbH6zZfUIMUVUba0V4imlZEmvRyIXwGy13tzG
YY7RQzbY5YgSW5G8kA120sTWGVnmnVva9d4+u7LloW8xDjRyRoj/2GPNTumc
zaryAr/DNYyZiNBZBJ89w3lnFcp3JAu3CwCblwlCYKn4jo/QJTOnsz0Ktrwq
AM6sq5jRGWeTW2MDxlgE2rpsJN0N6HuvgGrKORJ7eBeSbF34A5qY6x4n/hqN
xu/vDljLjmTVjlWWNiWAamtqbD/QN32PU/p/jxdqBFRp8Dy1uJ37RRiRuSRW
+932V+ZsPsvKRRS17nt/RcdIhAJmgmLz6tXLCzXnZUIzc+Vr/ulAHOQFt9BJ
9xpTCZCzhGE726E6j2cAwNqJmVLLdi2OnYneQ14TP3C+Mscmfse7eu9iJkFd
WJ9PKw3VAs6K7COWo9qVdCaIxm1uwb9WlCq7epa6dsy+5Q3Sn6d6N17+amfj
fqR62QwuWD8xYU2g1dzow0ksnJO/6b9GmuyrBqKsHNhdi/x82VpH1JPhqcjj
o0TqDewCSA9pvqezzjuwcGgO9pugSWFQMy3VWhoelzaJiUYLYTd606WsslmQ
BhO3A1vISy9q3cqMELBXxqbBFZ6NGrCwQR7IgpeeWdioTWdMDnRzSaNo9qaf
t2lGyBh5JJsR6xI5/oeyary7L2mwyN+xoxwVCWZoaKCcVVXSrvgIh5a2nE06
DW/5AHs3cqMNfoRHFKo/eJt+v+XK3JOIHyK//r+K+3L1N8hBJXv94Wt6Nv6r
BTI0hTOj0U4Br54xLncN3axytQdAuY3t6MYIk2KdLG//tPZpUkGoU7QM1vCD
/V3Uh3oL0olNxTU240NNGDvwGHX/p44QnhGxO3RnapytpdEeyZkhT+WGa43g
NDrynCTDibN1k0TxB1eeSIh17ya9OSKyoR5TBh01+LofZBbx+oUMLp8BOXOQ
XUrfw0jBCAa9LevHTDoq+JL8lKZ+e+xsc8asWwpzVWPAk2gnmbCHC7elHj/U
3KFUn9emaoJBh/cFTU+uu1P/NmSc1m+mfSmBYjjcXwnHb62bSJ/hziZFDTXv
9sz+2mJBgOEWNGiualCM/6p5uyFSR9f05xkUdGjZfDx+uxR7H4h7xtZ2UYzm
dwtdM3ZrMUEisKTn57tBQHeoJTpx6xoyXoelyzLmsculvuWjL/IlrIRmuZzd
kXZVoUjMDo0hnA7O2TFdFbe9Bqnw5KfMle9I3WMjUMOVQwgnWrEJwZBfaj5e
9yBzdSTW9q2AhLQDcVHUYy5FYD3n+cxQjIK8eZBCvh9nXqT9JAbhGml+ZtAP
iu4z5L5ghluvbI+dEAMtb6RmLhqoOOnFno35fmpI4nEZIizK68iBpNwfcDw4
4+2+SVou6zhNnbOfgFInEcaSxBhJvdRX/G4NArZtd3gxhgjLrd1o4DJMw9qK
VxKyK1F4LqrlMNBUH4kpxjy0ohXInciujSIWJZ5ULTF4nYcl9Gg5ES5EX+9g
WetGqbVBnU/l7y0WDJdskEbdXWrS+yrDEwleZ8POVPRRXte8URWg9Fwbd4t3
jrq/8z29SzfvET/vUvz9XAHTWiLZa+bh/TA4FNzKPqLo2PYcvNasbbn2ub3H
4yGdV1c5SXncgWliepS/Dkp4JeS4npLjOkbMocs4h2TLCSyS1Bjmg+7fw6Vo
SlmKYrtTANLGpmJZYzIF3syhBS9Nkb0ocUOQP6FEts6LTij7AGazjMlNdUKz
A+ZCvKMqn0G/Jpa4fdE5mbbZnJ0O1AjmPWMNCOYMrYdKpF5lk8FXb+xJa2LQ
hEpuo3TRvYUq8R+MF4Og2lXrARtOyEnAmF0QQtgjkumWYyqskDB2ZoIza3wY
AoC29qZMVUlXWNI8pkHnKTqjCI5W/02gRlaO7KxBzkIuSxKhPafXNaFCunkT
6ppVDDtUuTdzkcUHPOkpWthWVzoLn1vL3kKDGOopt851Z0qzJ0WjGklc5IRx
tHbmmK7XpsBG1OuUnMLy/JmfbMLxN7m+QCYaP0sA3MGPRazHmjS7Qq5iyZW6
lj7Yrp2NGR4rpcdM3KscFon1q6Mk+oLmYQR5llW1vFbh79PlQ+mIqjJtcYyK
eSrXqX3WdWJ3t2hyf/hTG4mkIGNtSrBqUr2OrhnQEpUBhndzF0u8JacR+aWy
daYVvrOJcYo+qkjEXEc4gKXQ01+OyjWbVH2AVAYdhfnKgZITo+d2opEtNnpV
dROItsKZR7R4ZBEZlEV8E+rW8p7FNinQl6ZHLN5NVlSpyiSG+6y1z+1mjQxJ
4nOXfWHhCH8cAXet4qdrsgp123D7/YbGsnaphw+TQ3u5whJC/jq8bYvnq4Dq
mGN/mN5El6bX2PG7AEOXT+KIEORmljYPw4GXLHGJZNvljKITI/QrpcG7y2Sc
DSPjt0FbyHglhqJ4/gDvldUEhftR9mOvkRw59JfV5WcfZ435QyozlbQm/SaJ
Y78SIxyr+/GgfiS4N49DXWOLwQMcMaUIR1eBGkzL6fQIYaGwSClKFVILUswc
SAwY/B/WQ4XQRj8T24h0GY4pcs32lUId6RXG/aBPEF1ZY+btG7j8xiIPEr1/
0TuDFBA1JSedeGRA22nTQOAnLL3O4Eza31EVoHcC46NUsQl4S9p9+FfTDqHc
5xmEJ4Wq352G2lrIxD6l8b7C+zXHyV3irNF+muIxB+UYGJpUwywe1/NE8v7P
5FVxCeU/PQ8j3UV0acQsa0Bc1OZSQ+lSu/ZSF3WZsq+BbyHD10S/BQ/1pFbm
UGUDb/kpRv6Wlgo6505es1KOocxHbJqKeYHeIMGrhBUavki76W7styQ6WJo1
BrydnFgJkeEaoT72Weng2gq3/ITGm6ZD5mColA/XO544FPXKDJth9/nXitrJ
bJdg/HRkat186adovsGHVX5cHw+8JJFbPbqJnsk/zWFNhPPSwUfIFC+MqnFI
ALhx76D/Y8jM+2SlW7XZQDzlmY4C09DA9bGXT1/Sv6Sp5huVdUdmqLwbO7VF
wqaQilWUpoYw6Adl/5Y4AuapKQIPZ48mx6nz5VFivl2OZkpNQW2Tqpi0UeLQ
qc23NMh0HXYZ5eJkQdNYj3tZUce2ygBpddZW9Rs+jxiqnEQChY02XLT77tpw
4wsYwngDbgMt76jSiVyjEJEsLMhbTh2D/laY7H3jENZ4Q2FnubZlEZFhe8h1
qe/qqoNTshXZ/a+U0kd/Au/6CCCP9LpG8da6XynIFG1pmrVdVazVbiyz/d9Z
l6CPgAbkhu3cnt5LwiATlBjSA4zPAqGM3ae6GuOYS/2azYHOTC7BfGLZFZ/u
SzwmBjwbR5AKvbyvmG3hqkdRaVXc0lLYMQTkR59h0NEs3mTlZU0u0v09wD5c
dZ84l2mVLeWkVr08kty7YI//y+2/j/uoS1LRctuucPzIn4KQ0qs9BMOdMTnm
HSOISle9V+CNg+hBQYo1xHc/hmqDSYkBjd/ScVRhkwgAks2Ig6d4OW1aMjnO
ef0EbVzgU8VdwczM/vTCW8X6Scv9IRAL8vtw9A+53OgHu/LTbEmrtXHcz+un
UTMl8cIsDyCPVm9D1KEzPK2u0RjNRi5Rn23kp87M1+sIgLsozcODnkZoJbNJ
lwQqQDORhIWUwfXRjkc7jG//l5+xCi+ixMT+iBoaJ1JzTfQPsa6Cg9Y2d8PQ
svrLY3y5k8Kt+j4/EWRY88Ind+Z1d8TMR6D3w7RRKN/wLe1ACEPPpIJ2/opU
UnOXVFoT73kWhHXh8Z9nX2H5hTDA8DmKtO65B9Lx6dIGvQla/IVynEr0y/LZ
PTej7hUDvk8GF9OMfTMU5nxUkh1HwDkLgjFWe2qaMfca5N13/P5QaR8BnaRA
3uSynpuq1Q21fE2UxvcbKL0Dj8CPvlu0BZMMDC2WUFWInbxorppap7qtHDW4
ybUoP6x/2+ZgPAg5n18o1PgA2wfib5UJ4e5A2iTAGfmYmjGsfwtVzPZRbVtc
SOG/PLbAIZVeeFC9IqlwiBsgG+giJgcSF53l37z4DFqNAlNU6GGZIx0PPrfY
IZvbX8lM4EnnOJ33Gy8vHGGZpYqxujS8Gz7ngj0LwpECFe5k+gIKrM80Y5aI
cMBgLuqAogIp24uA2Z8VX/sx0Gx5mPciXBbh4uaCmpm9p0UwvMdpEySg3arj
m/iJzKaGyeaBiygrNMkP1TJ4l7lJGUJbT5kfg/tY8en7ejP3h03HrvoYd4BR
L5YnfCYseceXmAP8Q0BAnPcFFpSts6jEIV6wIIycNyTL3xFNPO/zKCSdIkF2
6HHpz6OZYt26JY2lKX2nhzz38I30tHU1ydcPyXSRvj2YBexRExb0YC8Id5o5
PsaJggdy+6ZBuL8//BVHK2/C10yXc9/Ncss3t9cr/CPzDGyfwARZELREvWjE
amgQBYZDZF31GA5y59EDUF6lFogctMjCsLHLQg/v09HbRpqPIFF/Of4e0tTh
PJiB3jmMyWq311NmdeKxDvQmlwxl2OE97LPLBTTyvVoaBwLbsLGDHQjlnsaR
00/25VbrDsEZwBr8N8Sit7JopoiXWfuPQIkAKHNvKVf0mUNshEpo/9NASozJ
JyZWun4Ati5io8GVmlVY7phMjB0hZ8xH8t2EmCm5Spb8KvgeCGfNbzcI5Pc/
XWpB+CKZNA/k1njFsNqQpq7AOcQ3ZiBk+OWtPBaTUfppK6bCCCwnhhERFC0g
9y5D9xJy7awO8d2RDHzCTSLVOKiSvQ2UR9/JNS94D1T+oOQeLrHXI3ZvYp3r
BGiBVgscyYdo8aCojqvVnBf0Rth+r7f+KQLHf3BPcyzVDPw+XIFCXH7hpAxj
J2VUn5awMVxUxGVpzk30iqO4EUp8wwhD5A5NTBVBUrX2BKtlZJ3V4K4yWyuE
/i/vRmPxdLBrfBnZOznHGpNH3idtnpwtIUcbFlBRcOulITBrg1gaIw4xVCRz
+MZtdGdj5tlWQPGGjQlnoUup5fpmwiajzNm7g5z2GJDLCpMMwWEo3ItEhieY
pR1QOK17+RlDCyJLs4dsrI+DZmyaK5BUlPxCm94ilKAPXZOPt8/EhKMnFcFn
NGUtqEGbFBAePWQlId7CpO6PgJkNcWOHUvfGW80HUVNOh6wIH3+5/6lhdFg/
iHblSlW5L5D4t1a0q3KdFe6NMUJByQyXqOfTiMy8XKqHG1c3h8IsqsE1wUpl
5GSvynO8X2+zTY2S0e381avsqlDGdsbiQ1zydb2WSmaHmAZGZTOnfvF5oFdM
TczsZr8fLsCpzGIXI3nuuHkHQKAi3ZDoLa5cybZMEcarhPxYhFXCAh9He7fr
ULCYXImDs02CfYPhJp5ghM9cxPrvFB3edlx1Xs9v62YN4E/DMP3i4WhjU9Rh
1mICgjea9BjHwXrOttRO+liYc2WM1ywsYYAgL168rmDL+f17jktLp1SqgBP2
rGHXxSpyzJiEPXI+bBgEpqhGb+U7tgDxd48N7k6I4bGPq0BEXDjYKpK7tvJ/
fQ7WFg7cyUPGPqCLhX+89VmckIOvZOqz5lFjdgsOxYME3VcCLyCHzDcy8Nbv
gLz+BUpTJ396DaFVPlLuDTopFGVWHkjVHu4vOOciZPCxPvSkL9ieVBS4WEtR
m7wq+T8JmSn6CPP51sN7d4tmmtvyc7TtNGk0ivJR6tbvGVmqQR9HJgHXu9M/
8W7GGoX9nw5hSNDyx1ZylMcHb1SVvS1mc5JcLTpMPT2Nfx4cuRbjQQSUwucG
vk0kM1EzBUdHreYrfcjwPUQonnu3vLngw6uVwwsPEFsRcGNRLn10OOGWvCwM
59ewB2NvK9fiF+wr/ne0SCiCEUIehU43AcuHaVRyCum23W/cKwOuL3vc2aRn
oD1EA1Xed7KHRizaguWH8+mVVOrsYfHmK0YWzaK/DF0I/hxmJNDdNUDHQr5+
AOTHLzv/Jrl/faYhNH7XA1znyHzQfcniDTeKh0tAAoOi50+8i1zWQXRI2fwR
TUYASgFIMAtoggPCRd+8NTeUTGdXXI6wnOWjiGAp/jivDp1lze/o9+totYAI
Dgp/X3MWMstJDNAWEUjlXqUezUhzLUfaeuIOebbY1Hib90MtPKnP9uha6XLe
BvpyBaFg3NqVtM1OKtBa1ym9ufbKc5v4CBFByADkKd6cSjGltWCRSCl93c1+
F7+fL1slvjsXPyZ3cPLrWKaE7akW1KY63LJKz2yhWZ4I8uc32zUj0i9XtRCj
TmIZhGCHPiAb7DuE3CQhU6IyQl9optNPn9G9Q466BuY4ydOD1c8HTx4gv9fh
E8UdwG4o1qGjOicjuqZiTVbuBr+YF0PKT5TpQ0qp0LiDXWz48xfWMdBoLBXy
G1chHrDxRHgaEfxxCNfB3Vu0rwKWa+JtwRe/H9IRIFPRe2vYT1SnnqdIQA6F
MnxnDNro9LPuViZFyKlU8G5TrJ8JUk1uaNwYBXSod0l23dDmhRxHeKi/k5lT
dKJsHcxeofXoI3gVNKxuGgtmvTjLv+bOs9k/3vm/gac4mvPeNQzFNRoOqXDT
y49UdvjRZU5KImY3NPUGGfqUGGom8crfSExtz3MUslUyaoSlpv1mILTmSsPU
kVNDlSAfcKIZenytYSldayeDNAHTB2w2LjvKTBtyPQa+S3vZ1qOffWaPsBbR
7vBtjj88W/AAXrWjlxebxtBlcVm20Xm25A2byjoiF2QL5saZdRiHFIUL+7/x
hQpkCBYryjq5E66F/8+12ZSHPJRuTPZndvP8xiTxsJC+VBXDiWt5F1x5WLVT
mr2lhuCaeEcjKpUdL3hSCqmhhomCXQjexsB/CpRDbktxqh+XGfMtgCwdydWa
Op5wOlimUbUeeeSeouXroceuFL4+Tkkt4L7kvUhWX4gIm5xBMFaYx4KbeC0U
BRDgwUgvHbllEAxHKAtA2YI9GoHmsukyMoThor+lHnRmtLvg+x2Mld26Bhhe
LDwQqB0hZ/gbNDTFE2XCVhl64oUZUwbF/vHT5NM/cbx/8ZubvoyzbRB3jERX
ZuYWq2NpQabI6uEbTlCzvSkpDduqqa8SSJvSkFsQY6+27CViaxP+sIPROHtU
uTcr2tkjKzPZChYB8YrNipCBLj0AgQ2swis4cZNYi7KoOxOsKMzvZM4MdfeW
XJRJoGkXVhqyoq3bft6m+cFbXLdun43zQCixFM7FTXdU1fic1goJjHyTQdye
8VKrdOuyPMUJyYy6KbXrno/X/7Nvl1h4Aje7WMa3wYO7Q5mSaKv7mF5WzAgt
5Q/xHtxXUisbKD7CZwd4KUIRUEusl3zDMG45sSFhNAEThVj5NJQkYp+Vgm0S
qkRbYDoSxBwR8iBPCJEqCrnB7RD80Eu/Edl3g3qa8ddAooNADvOm+mB6nPmN
DPEgbknxQwCUe4pysXwUiJIFj0iWAXhIztlRwCl5ZqJ2c0zKRhokuSu3jTLT
MnhqWc6P5ouK+vKQuKGl5+UM6CilvAepreWVNvefanitpUsJ1FLs9ZOH9RFB
spA6RA3V6i0cuZYkEh0bfeurgKkBklisOV4lNZSQWVxcCKjr6pN0lVCKLIun
PoRU4zv1LvzQ10pV9uOC2TNpydz8JSEx5YJJ7qjDz5GlYA1GJnSFMn5VWVFZ
YoXOrdYuxzCj8ADIAgdUgstDQlR5jE1qW/uOZLKhSvUe9BL1W0WLZu2TZELl
cD6iLYSzDk3YpQWS+9qJKPNSJ4Lw2E6miaI0kvy3VJatQrALrHIfiZzr3xT8
3zHipgBlTnHYJ/gWQ/Yp0UFwHqSal25qPAPtH7aNCyEBDDpdTapJtjOKSXzQ
h2phvyuqiTefgLyEl27OUY306HKSc1UFm9AfmWAFBRnOXTsQL/r30bAtlwyV
RRuxKTVouyIbHa5JgOulg31pT8v82iNnrnoPfbg5dDzs7XQxUIb5eIuRgzaC
M+l9dfAwz83sPNtXLVu5wyX/ag/sykRDbrn6uNf/SmXpU1x5u8ErbfhvkcUx
DLUQpqL2LsHkpVjBkHuk3yl6H01r/WSjlWqUe9rgo6OThzx5g9yRoyHriOrQ
kXkZdOsFJh2P+RdTg+8V2DmQm05HRthLMR49sD7QsutRoetuqYY6tVG9MPSA
fa0qR2WGJYWcXNyn4VOFtbXJOyBoE4b2orsVydlLbWHMfVm2I3O9AVuISeBq
mRoWORmf7dL1uVaXfcC1mWLMQeUIwqHax4EwtfecFCcMC8z7hOlpd/RZ6hR5
Czw8a/I5wsXXUJyCv43AnG0H2/rmKVoi2LlyLAJs1uNS+hptWVCxjdzfKXKQ
32A3PKZlRWNvECAKiAlmDcN45UL3CCHyPr6li2D+P2A2NXPxWcZXunqoudBM
8zvUXZB72kJ9oPuKfuNydf69NXmWp/AJbGp9vcKAvZQHq0JO3D5RxeNhaPn+
3n1oxroZo99N3x+0odNrQKBrvH1MQNyMTjrg8ZGMhCVHaQHT1Hxz2ThXSxMV
GdD0ylJCYUJ2qlgGxpP/1ZwYw8kGcvcLYw31OD0IrRtliRqmbhUCXT/aIrrx
ClayRcirDX4N+7JH2MXnjfyf8QcJFCAKCSH/o7fd6hjIYZEAYc6aGZOgQe6s
YTYXZ8HQQjbYrZNMc7om4xrP34TJbt81eQhaXD0ewdjgcZf8nE+NBvwwAOF6
ymzc6gFebBGkFodpCGPO6+NTlYqIw56Ng+sz0d+YEHiMT3cSMPzKLMtYhy20
FEBpTzzmAy5zfJwNdF/SU/WUrZIgAfPjLd74BbEUqAw6oxIKZaxzBBwy1NHy
7nTs12rvU2NPfrxSP9qD6NkQovapLKkvN1MiIB4NO9EQ15JAFtZvVVH7u8Aw
quzd5bl3tgjWvlL7yUdG1SsL2p74SYcHYAeZC55cVGF8PRkPximPf7j/tIuM
qQNP2u7lmp/VEsa57adU5L9DaTuLf4c2xC7R7qpOTocouZyoWiX9omYb9rrX
wFs90moowy2p2oGIEZpUwebolqry91XRww1aDleSetmYxr8k1OOzN7b0VQNf
eix5AWkzKrv3xFcHv/IkuRzds6O1MXZYC/+CVbC3Y+SxqQf97DVjitLsBQxa
Vg3HGl0Djg++5yxsdwSDSjMFryHSzDUuoF8I75EcVFczGe0b7qlzd9Ilhcqx
Lyh4akVIR/w9Rno9bmGM/URJZp0Rl5Ov33nlUdryK7KFfiejQI8xSYgabr6G
uzKvqiDdQ+CoTNT8JiK24hAa01hVsdio1RVJUFXdFb7Spf9gy0+XNudaEIoq
daEsF2w5rRFkTr8wbJPILpzV2FbjuRChb7vzM8JteG9M6GHWoCyMnQzzZW01
bLFohmTm54YFWL3ykrLqkEXTUpb5AHfxshzAZrwnIkrj3+bOpUZxrl6JAfgX
zZGq39ERKnuFhCzwwsh65Os191glnkzLDfkdglOq7K6+KKDoVkbc22FC5WdF
YdWKghU6a+H5e/U1q/fIygHddjApbtL2vSWnoNzolZ/lRXKpSugl0SP3Nqzi
B8w3G6JKdjElQeA7NHwPwVmk2ikD+eWDr34/BZXCfE75vS8vkn9NIjWyFgq9
39SpHF1zbooZlh848f79y7j/AevuhghonKlujPmXmuCjIzwv96NMq1ug8gXO
EIBrWKMfPzRAKFsV7L5CE0PwQW5AKAdrIFQSPDJpNDJAtpolApNdl2Ek80DA
GMnu63d5m6XTiyUBNa24uvlY9aROWSujKuydLGwW+2522umv7MlXprT7w29a
+nmAFEWHvWlH080R6rTDGN5Ujp2xQ5/b9K2e8f8XSlwskwVDqte7MA6lPd1R
i/720TmYnOVzLD8S1kaBim9AoMTj3/k390Rla8rqk94VVOEeSIpy53e64hMn
8URRx7xEP3GxJhPL3b/SRSkD8p3vYsYwZWG7ahe7dG03Ltough4JZw3Z/Mfd
2MVi+vV4xc5jIL90sz6pdgx1glqEZILLOlu66/x2euRWv79ccXkzV1HVGFKi
BWcLDLaVx2T/RBX6WO6YGFvrI+kSiDfs02bm/lXPxQxbcNOq+0TnZjWonh75
49f+Vcz9NsJN7O3+bNgw09vq312IeyaJAI/IFs8cDhuu+7egn7i4kKgOL3QY
aYVEYteMsfQgkkZ9HSw8fdanSZw/MejBG/8dm4vNmLhsNOEKCfjIyuko3dO4
I2SFkQWo7PwLp8m9IhPSeMHqTMTgqvv25c/6DFa5dQcYnPbq5XL58vlVA/Hn
bNeS38fDWVUIb55CwoMlCTG5Z8qF6jqa7ZwsJJ871YA+MHFKhDuThHB6WVsw
SG+SD+kPzZTsku3jku0RpDPGDZK0Lj7yoVuMe3iPF/8eXaN8RDZUNFN1qre6
zD0XMLRcxEPQ9Xw4HVS1S/U3RKniYoeb02MIpnymRIowNWJmYWTxwLZPmNpV
l02zJKFlaAq6orrpSC21EBkc1AbaYI1rbEkuSkE8kERGLpjG4z6n+UEVyls7
znnVH2vygGjZOiDT1333R76Bh4zwtAB/w+cefk8ZazmnVwVt5UJMmL0UPVO6
9UQPR4KcrdVwAmwvbbJUy0IuBtT4ywDJ1SDLUPpmegTxr8BlNu3SHo4eT0Hp
zX8ODjlsmVUEA170OoRTK59WYsWpjbmzEbrHf1i0+A8yDXG5XH8Ue6oLbGIy
QH1KkjRV8qtBK9dfz0x9HX9pjeRnoaXodEuUjLsfD8wjAJek37x0zb6v9b0r
2w2dJrfWuY/IipelTWa7jGb7kWTXbX8RJxWRfOZnDkCoFxW9PptZUdTcrx2R
+PEMAmPUK+QipJIAW+nbf2y1fcatB95m+5cPJ+2wlDkSBZX3HQjpvSIzAmkd
nk2YlqbXFa4X5pUc+BNyOxLu1vhaOUHAo1ioMbsFYvEDMHh6iB6KMGsavgxN
qv/n+B/mvFPbPOSnWbQ/Q0xeBNcKOF/lej2cVhoCPiapRIEmpZTXznXYTVlN
BxDWCyoQHw8MKwSMwhacKibtcRiYY9dpso70eoQ9IVbD1TpQk1kzeuDet7B/
K9/S9PXVBzJrMSOONySC7pV0hUC22mwVmHz5t8/6M9b0HdwpVDt0/9F7SOUN
3oq6xgs9FAVM0SI9vxBnOn6IYqOBhNlKUYpwHVO3Jx7/kfHJUbF6EVmqCq29
qAMWFJm71yrIcuI0FvQil+LQIhUxcn7SH2oxQjL4NRFLWB8fjFfY4LCGqN9b
is8bwvfZJfFLVXfcKC83vT01hqIbjp1Da4yT/FhyP6QN/wcW7wY6rraJYdwO
K4rpuzdXW1MDOYi+kDIKRXvNaBSXmOh0btO/w3h7nMKuVZbEyDag0M+7dK6l
mF02UiEF403K9N0NwCJnrtVD0hlIpDA21kBdbKmXsgm/xZW/Ob92zhXOmBMj
6RInw8rJULlBbPpozPFUQ57GdTqtfGwwop+FfoGqNgyqJirh3+PbX5VNYC/G
dVAhL7p0aVPRijmBwDcXoSfLNQf9BZLSZsfqvUc/4eKkO4kPh/+oebGMC8Ny
jB4DjISSSOzyoYMUl53vX0j9yRCJRQIC9KEcfIeMpXGGBNsq+qAtqLiXU/sf
RyyHFjhgGshfOejoYRYPiSyMyQ1XGjn5o8dKYaRD96sq+1uI1SoqiFhYH+Gb
2Gna4xF/zRA/vVo34+BGKownLVTLljysvVXqrJEaDHLrvkim29gr0E/qGc0Z
nqmt91mNL1K5rbOq0+iuY80l22IOLD7LW5E/4wqQlOzxhgE9PCr2vbTjPR90
0l9RC6OK3eKrFWdUzAgTh2m0VYrqxJb120fmz3HfF8RvY5132LuycIJB7f14
zjDgch7jSe3v5tdOd9+4QHGVGspFZQb3Ul3dxRnQt5nrvn5HS/jtKq4JvHO9
ef2kLNTGbRo//khd+6CXMmhifEluHPRPdNAAM5ROhKlW3W/EusEO+8PDMQlZ
XGXJQxLFEEE63RNHhLXHp1X/Wysy0DB4tvUvyTZkH+0HQmsj6o6B8MC4nZkj
Zy7K/AI5gL1Bggd8v0EvpaWSZFIlqIjO5S2UTdUn8YTvT+BT19AIC6j3HHJ/
aK4Bsl1QkoIx8aCdjgudKCPljL37jbvQrRTETegDdU2iGTNWJCYx7NM1eEgf
RSfgNZMtnMwu9Sy53zNfHPRgo5GsjG5HEBurvPaFxB91qDJNAEN4+tLRNp40
arV7qyEUDxM5/zr/AQVu4vpmCp6nuB9WdkRDXzAfNXr9f6toFZgeaSkVkoUs
qpkA6shmIpCYjWXPZwrf0dF0NAxWCQTRx2cPtwjuwjtkgn7LyrYg2+h1eVGx
Sw0Twf7uM+qBJ/qBaGgGl7A340wy9EkEy45ng6wtXGXaO99h3vMmC5UrPTqE
IFy0YQpF03SiGLTuW8+mjbbJS0IFczRTvnqzgegR4FPdjwL/nEjzlH1Q7tvj
6ySm9uYDKXKyb3WrMyW9By3UsA3PXoDPLlA4WPtr/wcpfGvQfLXNMYkWeQq+
HDT5JB1VOrRoBIaJ5yn55NZrUMY7f1J4IVqH6L2EkVe6IdGhDcOpl9dkHEqU
5j/f3Rw8sujFEGvw2S2hPbC49I2HiiAapJX2iA/sXLKn+NZkNvrgeLK3nHWp
8eXioRycDT4j4IFJUcjW7GPBW4aYU2pSeIknJLtp4OZij2RSXL+isOe5mCUD
erf8MH4ihq7sWw2m5bO3W9rs7Wuh8BFH3LTTqgL+uGNmi1xgkZOhye4hpBMq
bpyAKIZ5yk42pjj8kr67Bfu0zSSKAoDF++O+lgHQgOuGd60EtUlrzDgQ4ufI
vZw2z61PVQhJZ3kuJFb0wgJPTAF5Y+ZTfy+Jr9EDWcjH+AAIaDoHPUt4jjOk
wOkcNsDBAlYVljYEL8mT1qP2Ao2jnHeDxqpM9Olb3TWGQc4fKc60pxF12l8k
oKLnv9SH6+TmYHIxX/E8ZD/zEFbp7Lmy6xkGhrqQnYRh2bvDT8+pVEm7+AKA
LQTQITEVww57eecxZLObcauZkDGxpxcbn5TQSJjfdutd7rO7YjefHl13ueq8
1qhNf56AMLpLXyslNdqHSVmb9rfX0PeeS+xUpM8Qu0V1dcMa2BV6XpICLh3E
Xnw4vWNTsG0c2EArpoFQUEwFbctgNcrv25xBeKvKoG4RTbCoXzrugJboBxqc
HCm+2zN8f+lSWFNgIZkAArgkPzgTx+pJrAHFIywbcn3qzaI4KTQClM7C1e9Z
RawwCYvB2Btzu8p052wDJ88ShQMCD73kJ1VgtHA9qVq/7PxMLsL62Yy4O3Qp
3GhM7FGGKE6bzokFenQRAQbh+N1oMAnqGYgia2vQHMrXqZ0I9NiSGUGeBHvy
j7jDJGo6m8h7PeIZMnzEBNrQF1y3BiHc7sUSHBN5U5KwgfavV6nIzQ1MX4lm
XvZqib8KIlECFH/oWLRzOjpjIpzMgpMI60mR6TXo/frkwT7MTVmYvZ6OVm3o
B/RlGEjsfRDtNU0hZ4slXQ21/LtclVTmGtO/mEQtvJeQr/5ac13tFIYetUAq
6VPBwpsiyPiE36REvSxMWJkyXeHP056Cvws97VUil9Whobzg0g6LBu9ZPt5q
tnrtD5Sbmr9BukeOR4H7d5WTgMX0ibf578zKP2TGYt0bht3g2Qa9Irk8OH47
/VDDX+wYtheDbI++OmUORyZfQP8pORrwlXfZTg3TsXuJxDjj0xh5H6Ja3J0Q
44SoN1gjXOWkZvl/tUwJsJfK532BgguqQKvOMQJaj8BqiDMrwUR2RH+6c776
rA3p/wlMK9gaLLOT3kdY1njEasUfXMtlbLk4MbGqd+1DHcpKx7xv2JmZ4eIG
Eo4CYy2vZs4EWP920orJdFP/S09hqViK+FvDJgEnTUGiYnrfo7JGvASxfTtd
WIa+HlWXI6Ykbx2au/gQMatp62EbUxWgYqjBfvrEgnFKmXvZV1H3KGUHSLza
W1HqAHAzxCX82KPKWojKOwsS/9Sr2lHek+DyJCWY6BbiSSbHIkrx7oWUamMl
+CW0ssw7CZrXfHmUUvxV66aV2cokWkeDnGIq71oVJNJBkWAjQ3NgcwC8xnhj
jqjRD5MBk+oeES/z5i88fCXNCeUB6Vyg66f0V3ce3xShPl5fPrykuzqJVFfb
akA3sZFCnil+82WATm7htZptlOSnaTxz8X3EC0PXDqf2lm+kgA3Yrbxrn9Oe
sngvCJO0zr/j5Ydx7WdOZdRP+mUAK28EjJn9N9hgNrnPmIv9HmAKrPO+NNsL
4z8c9zwPMsXogwi4czcyYN0T8oYNzZF5E4pxKtY6p9b8sx+Puq+iyfNUgbs3
QqBttPGpmyCjdwrLh2QCIqQU45MfRIAnJwPOkeLLxl05lfPmFzPWqGchQqxB
ohKbGEjWA6xz5BYKF6+Jh/laQTPXiUgt7yvzlNeKvIzlVxxITT4QCtVikprU
CV0LZJ2HcEuPtXDa0BP9glnnrAldxjrWHRzE6FiIUgMhqS9Nop6XepBpBXDa
5Q+6IGTUEpP4/zfbTjjx4XkW/MG1MElTWiPmub/Ly6XAqJNPSqhrQh6+WlJ5
/JLgbKWSO9nkubnGKh2JOsNndSF7HyFLHllsYzCWIvKntSjAxIzIpryQvAdy
C01BWVVs8b/t8FRhoHK9u3uZbBVXc1D9my202zwzUdkQiZHZ0EfLsn3sM0ZU
kaQDSVlvaPN3L7qXK8nBFTHmWn85LsxlDnfeD2AxM0RYj7XmyCB+UAZOvnXJ
ZJ2CLkI6HlydEboAoKYYFMuaGhXbLUiKcMKXtuoCUJWVgHFj6bwyrOducihG
SdjFHh0z8kNrqIVK4+P3Z5LrExUaBOkPxMEd3jA9DRYfJiaxegnkxjtyoZlS
Ii+UCCD1ApkqDXUKbtdWpqFYci1TR7z8rxgUWdm6wqRWK4tBrhPygTuPB/S2
CTXGhgPu0R+VYmV055Ylap2ZghczH5bTyobgMeAgQJHHhmQss2PcO810u4P2
EVDv1vOKa6dqeF7A64bCGVitFsYbJhTEDEKtwojeu1Z26bNE40LxNHswA6gd
oZnQmdcGdVf7HbceAbk6w6s6t2Rx0MOmm6GBWMAtemNzSLILrr93Wjrt3uzk
1nkmlJili5KYGQQh9NmOI73Is8jprP7dzVYDrtfRGTPAI7ytSt4xAcfy7Oim
GIPBJauytu+dwVj4ReSOpfT94ChUbWjHZ2E7yqdGBexVyJ3ZAhDdhziKeGf5
0Vx+QzvOLLtoKQFeFZWUfBiSoH7UrWNEcuhmaMxl+gKfTtZ4fytE3KEk8p/A
1+M1SAPqvyCvwVeZ2rzXIjEgaeU/1G+bCPI5wRchEFN4VTJNOPeRDUuX7Lwa
rSVhHeFxx7Eti3QrUKtxRWvAdxaiaYyPGWk2qyS1CEiF2s2pqFMgVyf/Hd+V
5pALxNi33U7gME8Km1m6KBpMaPv0fdYKZPrv+QrGbka5oq9XM0exDdTv4BnO
LbugiledfWBnfE2Ta+rWfOMOrkBCVgdW2dUFWPVhA4r9ZQo/rHlxWfPX96tp
vtwPyE7ca3m9sT70vQE5N6IEkRtKFzMLz2y3d95Wevra40qe/LOSSt+rdpb5
yl5apP4UziKspYHgsqUh+hAyLw/Sl1g5lrYPbGLIVCXG7MznhWnEVLWxV5gu
1vou2MQfG8Kngu71e1rYPx5PVCgxkDsRddn7Nwl+2slllDO2nHSbXiuBHi7l
9QWvm98Yz75BYniUzuJeI5orHZpU4cci6d+AeHGZQtgeN7RGUMMb2dV8dE3t
nNA0XpuPxSBfecP/WfnhU2hh+32+V25JUCfQLVe53W1BSOT2/ho3sZETg3VF
tbOg31mFTzTo/MbKkqZmQCW/twaewSM3vsu5rf+xDQtqbYKgLNQhW/CY11B/
AvVjEk4OGtT2z9ZVTu+mK2615Rd8rKfRuJXxcEH+gPYULOf8S+OTgd1j2pdd
UZ8W1qhdPToVfNUMca93G+fZK/2UNdTziTdUHsy0UCUe8AFZFdyRMgLYmQvx
+UFUCGAsBeUZxP5mB3EjNvxMuFOlTl6cs6FgrwGVhFBnyKOHu3d1aSFDmUv3
bLfybmJeZGzlM+42E5/ak8ywxd0jOjLIAQD90v2ETeZL0FB69Gerb9nCphy+
zt4k0AiSlkeJQLDZe8Vct9YOGVg0zdyyEdsY+CtwKGpiDFQyNtAEwlrHY1VR
ao5ke7d8dXq3E/yhQ4K4gxVgzqLc+jYPdy0OvfaQ3eEU49fQVnTsxDIS7N20
T6/z6agQ02NxnAIpBiTM+wAHX2f0dZQil0HDHReUtrXslZTWinah71SPasNU
JXJmn7rca8QYjsiVtrwmAaBnI3sK2PhvwpDXIfbKJgdDMwAICzrxrazLBQ3s
EqTqAbRRp5on6aQ0FlrVaKwGDH/0ouHwRrFU8NNnNbuj1hKmxbupsuntbrKA
rpUlWRrrPy+OoB8IMzSC/zjoml25ZUCyYWO830C6IQ0bM91JANveRqYz8ovz
qMsVAvP83yZyC+hJyNiu3J+bdQlQhzhR4H9zzxe6t0UP6iw+JMrJY60qP/0W
oEzldE4G6r4GISbJgy9aSd5h+CRK65QDHFaVJTkyMGkyBvRoYhA9AzwoJ2J8
x0rLk+5crUwuVQMADLTfNpnov0ldkrrc2dqN7hZitfl3FjamkPYY0/Af36lf
GBBCqdwFHgDttsrtvXFB0SNssnxcKvxLDS5hGgPq3pg3jWRsfz18p+FXKFjN
/j1u5bZXckjajTCwv+a24K81Uj53OYx5ouDiha/0yMCAnPhLZb7v90buB3tg
jezOLEBkKsRHwiQPg/savaFDLVT/yfoVb1Kmu8bBgIfkIob1gpl0UWkHQEQY
JsBpiME58T7R384ZcON+G2AzmTY23hyxYkinKD1Z1Gp3RVDVjnDzw03NljML
FOfCP+WXWgZ8K3Nz6aVUtAJdeZRR5I8WWldq9txOeRiGV7D4RZ2ndNLRo2AS
8Bc/bkZUeHmyI1KZd2ld2kHK05NKW9tFcA7lmC/91uMwoYGQ0qg8pg4CaaCa
l7pAvOCCz34R4iSctxPX2fkiu8GR9B504448sRPkC+2CPmD/iZQ6xraVlzne
IZxk07AOhGpHftD5B8eRiAGUQn4n1pyoshf4ZpdjLQ1ANMLJF5ZvEeI+PDq4
kXexjl0s8nXLMSgnPOfVE7Mgoi06XHyUBFl1iKsyiVecnPlsH2xYlWGexSzh
1OFi3Xd7v+RJWr5aHFfz8Qn6f+MllAp6MkyQuHiMxTyy8HnZSUCuZuC1ihXh
KCsIcB4BxNvPFc+CgNrl832OLxWP79JXfZJ/kSn9Mruuk7naDEOuIIPHoYdO
xaKNxyv4SH+GTtLVi6M4MVECnATSzXq4q8eZVyTjqowDY/zSH+wKZX6wLwcr
JobNxzDcoR5B8AbmgM8AZ9DVcYVOVuzF6GfgVLh42DXOso+RHXF89AVXcjgi
5EN1OlFGO3J8y+ZPVEc7gzfNgxcsGGmOhpc1nWKIPdAjWaK1AQ33aq3WqiJz
/UtHwWY5GBV6KiTODgGONv55APLB03gEaVvIdkucpCDjRvvZzL+QAoEKEXcK
rJBaZ2wENRzqDrXTR5JwoxgSqiK9iESHMhSZ79yMEeeY2a6GV97vEpj3jgjq
uN0dG5n08X0Ju5dlSVZzxYh8n1mGLaqZ9DGcmQqJ6qDwGJlmtN3j9PmUB1vA
YY0ZO6KcGPMJEzYnCpPmf4R1T7q2Poo8uxMV0yvKh9GQnjZqaPf74/jSGq8y
JLu9FssnPSdLomyzpk/VA4xZg5vhjKF79G5RUlGtXndXczeJk0dmXnZcmFoe
pqrPc4pZw3nMphDM6X9X1Med1Q69JdRN3baDmRFSoudo7RdN9IoLhi94Ly2y
Z5Mws+mftZUicfvVkp3JOPeMN4OBtEOaA9jPEO2vSwafrJkEMKKEMX57gUZo
fEvmiwQ9GbcSuFwo1DDoeB9H8fD/zZpB64ssUvcs2v3PUbNBvPssxsImcYUG
AaUMA7gIpcI4ZcLHEeVR2QUwLVId5hCgK6Kpm5JlpUugoUcok5ATBFhr5H2W
3dil3jHSqWHb2pZlhnU3ffhNj5tDJrj/RpDokF1VLdzGw0fOZLJDHL3P2WxM
PuBQXzBea1DxN0hkqWv2BZSzv+owRNwv7JZqepE+rKomWfW8ecRYEACjzgxK
y9PuFJa/gu7Eg5Kw2LawVvRy8PUE2B10G4ZTXfx4Q3h0z3qdC/p9/hw5dpDQ
vnDhQ489LexalFzHiU+UyXlxihVG2AQiM2/d1Se05V6TzusN5pjLbCfo8bEy
YAstKRWfT5zyP3RW4NmTrDTc98mWzCJTz+mE8Sm3zPNXTohNRw4iBVnpHJXp
KwVwAcx2CHwh/F4HnMDSH7sOF/iDrn1MjTNRZhEVF/9LtNvLxfUMZgsm6UjK
xpSeeyegM0rvnLfucpMSEnlEAaSnXjLq0tri9iPDB3bBnFXDZjV79JDVELwD
snOK9Whgw8RKrgs59juXK71cuenLiQlSsfsIjGqUsUJh/nI9iiyr4x+jFf+L
ioWxe1OcOfi8gQOWIsFo1J986QnRiyjq2u6nqicH4lZVFxh9G+TwvvTDuG8t
rhaofKe2ru3cONn+By4CSjJm5YAu55BSdn6wMrIzz6fqwWiqHum0H+JRcvFS
5EKubCfjklrs/zN+CtOncvM0MlBoVA0Ztqq91ZxbeGgp5KdtmBLs3mspRjXg
qceXIw+BkNaA+J0lwfqxvar0jbcXj9SVTULFm2ZDhJSxtoVS6Q1YVvPbWisn
rQivnNw/gxSrLzj8Ou8ABHz6ROSisCDHmo4Z6W6MWKnvGBvYUmcklZhvZ0wM
BPccqnHTaLfUxdtStSxx222gFTFJ+BvYibte5AyiBHbLeJ5+maocSVf7DG4p
QBxVNUBkOInnO0XAK+UKJlDgfdiC5aSgVz8WMmgsRm7/k3B3eHFUYPi+8hez
9IhuGcP6S+vLBFziePtklIMzsB4JdKs0oJCnIvJKlbX4/pW6CAqgH2yGbOnz
scbC5Xk5awJX/GG2z1XoExets/8teMAA7SdvK4qtHsR7MQmnOHCJfzRwxIdB
za5ixCz3x+QCSK+FHI0CdVD4gDxyXQzrPXxx8eTJRL8I6Vi45c8UH37mEok3
BA0A4zY+kIQ2LHHx04wmzu8lwzCiaZecpidi4P3J3zVuYDvOp5mMAaX3Puvw
VhdrXRfEsmSXbQl5YsNGFSGnpo0A3Y+dHokiJZYR/aL1tPMKna6T3+5S6yRG
6jZM0xrnnQ7fKbQ/M/Hq8Y8K4Qcm3uou21ad9+vIkHcbnRlUdGzM0+eANKPB
xq6mA/HcBLOvulETufWbTmNTi6ICuG2h0rJnFIyWuHD0kISormuom8VL+hiF
gklDcn/14LZQok1+1VKQu8UtYHao07v24CQOSewCzj/jD8uWg2/xQw5k3q7X
EX8FV/dcaqbPeGj04vD/WG/+6ACPr/VtiK+5+Wf3m1vkwVJUGloEXCWu/uBz
wSGNecYoIrwMGM6AsI/zD/mx/7u6SpXRu544W7JDkthplFkozKOX0343utoc
NiK21cYieF470XDc9b1lfLIVc35rP74a6/qOfJxE9+kLtgX7QKe+Tl1AQuy6
XZAEnv0LD++v21Ajsfa4RTf3ODTscLoYXmjPDCjIjcTG6jOQ7WDTMIYjgNwx
dytIGrbN4HhN3Js6AzGDOjItAZltblNJSi96kPt4Y2Fc5/Fq3k3R2T6RS8IH
UodHQxWxZ6R0qU92UoyzH2yg3nsDc8oW21hx7NsaNBIeWfFNgJN+ePKShy59
exsNQayPZvQGjIhjz4uuaQ5Xysfv/y909Hb9Eufz5DLrmiHDQpRx7JzgLeGG
8ZWOnUw/0UDjM3Vl1P7lLiE/7waiXK2h3fuW68rxVsejfP5fQ3MrUSew79DH
7eYiBUl+5LEjaPPCqUx8GZKWD9Co43FDYO/Ix2vRCw+fbFSk9a+ppDsyJdrg
BcZZcizfPfbZlh0Yn4b6DQt6Wphnq5jdRxdzAz2xM/mcBEfE++qQlpwmSjbW
opW58wq3T05v4z1hPkrLMnshkaPTCuZ1MZvCzUnMD6tmacRRi4b7Aqa++afu
Lmg6ZlkmNRTAUiUFLBZqWwWw6D3KD2HyTPl8dc2/8DiCvb0u26fYyfeXcj7n
KWbXwdKQjzkyf9idpP+vjplsqwB79veIriwOzVpvm6ItN3mBpVJHpyoMyrRJ
Y8UB3pNGFMkxZznLFq1dxdg7K3bHGEoeGR/6VBJZ5441YMMVl8Ylhcb/8/6n
2aBLz4yraCjT+iOZqHbfXiE8QRRiWt7vbEnER2u77nc3K7SPX9gZ5cM19Leo
osTBYdVj9LLgBUNIgdMwlhsIEtaT7/HgjyNwzkv/b1oxMwiCgCpDGIBvEXCO
js+7nqN4cJTPx5L/MzWJhHcoqYK6iv+fWS3XHT+JqvrS2C3hhLzNd78CsiUm
lQTHnmiCIAgNN8QCN2RprIVrxJjTNWdgDlY9BqYSmUySBlRmRplq+73/OscY
RbOcsDDnlgeUuywV3mqwGFOO8uaje3DUBH0idUfifuTeaHISnuSCcTsmmwhC
/jYPBYouRLiUOeUCPYf3wDk0gmyeZJTmFYPCc6gRxMYEt/YB/Xdwu4JZcY64
iCNNBkpZV8NkDYxrnDKkSMdMm2I5vFh+/uYhyp8pw/dG/wwujuxdj8mCkGV2
yszgq7N0DyOi0W2uNcrVI5S3fbQXHXMKy029OAcHKkeilKhf2QO2uZSUqhRX
qjXk3aSRj5g1giiB4zX/zA7MJjVYVT95HHDTkISMxIJRFZ6cxzYr/N4FGsea
Gmws9l+wC/9k0P5Vsm/UzKDb235tr7B+8KeiazNPzRdhqfzlAKR7noOHTV+O
poliwgiN7OLQ3b8bxh7hKWhWUBwcu6AaPfIyLJKVROq+xI5ti74SnwCN40qi
V5WYdG9W5bmbKvApggDi6Xw2jylk6OMOI1+yRoU0wQqgCbFGbrG13XKbLnGt
s8PJI8OzVLehjWjel700pMrxnazgofJvBa67ZTk+QHuaO91LoqV3+nNo95mS
E4fi6NcJtZjAw/+bHKmMoA8ilV6KqMpGFA3QjYcu53212JWWHMom2oQCe7lc
ZEwgLWCWPgKopLtD5o8HTT9AAgNSDHWe9Pb1Q8/9jvNWehKQRT1B8aMVL3rf
j9EtfNebx2eSYSRlZvPX6fNrpd8L7K51qMx8R61Axtvw/mgWeuaMAdI9fQ7p
ZjjlxTeOr1AgliYOBYtCUQKm34NX/lQnEo7inFbplAT8CyjSP4xkMgOst6fj
4s2dnvh6E1l6lodIl1vpqAvHz5yoB2vuc6+dS73iZzB7VFL+tDsrVajXrewA
PFAEMg6ZUceSf5xt0saiph/234/J+KD4v/WffJInCWo39ZRh/4gnttGVrFqL
/8aKVXMMCTwjJXhf4A03hAsz4+EZj2n1yY6Lp8nLwuikMC2Z7im+GKVcAb9w
cLvU8xk8fMbj/PQiTKr5/POCh9xeoM2TZ5OCDomENg0Ui/LzB48e6eDfAeZN
OTsO5qztS7aE7LKGfndqyAkd0At61hWaotCCOxcNhDCWQZmlCAlECvQMTQQj
0WR2hWsCCSgEcGUDhUWnhhX9btDqWY0DaBERnxdZZUD9+5lmXstchN87rYVa
qD9VY6tYz0UpErbFkH9VLujdgvEvZw00Fhz4HwwzvZB/qgklHwVWNSGvo+E6
mrdpEZZurthza8JY7chyGfwrYNtDMrGvulUvY0MkuLKzkNOMi/A8lzISpe4K
PJHOtECZ90N5SRCm1xP81uIXuI28dnTpq1jYZFpYdvmVG6TURIptzFau3b5X
6C4Me7bXksgHL1QTdEH497TT3KyB8wVb5NIU87X/UpOQwgefGTcI3X6g+Vdx
WdeG5sgrBwPX5lfCM+4nqb/7U2tb+F7R8DNBnr7mDZ8TMJ3qY54SX7xIh9MY
wqd1uT4ZNxVLbsSzv91yTKAGbJjwqCKa1xEMDxk/WnPQmb6InX8Qi8V6L5qq
0ZxcyNvwF5MqS3BqSbMdXf8+9uH4rS52Mby6IYNByBoadlGur6RZ3MEJxy5O
/nBTvQTcQa9oVG5M+xFQCfArwYYbZ+tslp6H6yIc5pP6EXwShU2ewDiyQXAW
dunP8GWFRFQGKZ5pfrzynqqIJ6VSX3dYiZvcfbtMhKpy09m9Py+uZ1wfRWE8
hguBfNv0qzfQMf3Tg+pZTP27RL3+doiHFiWUt+JR9GC7GmkETvvN7R/+GRLu
e+nu6sVk8OslRDcpl4LAWZNMAI3Lz1rW+Cprh+eFRnx5tiIhoSbwfhRGj4Qu
yWx2KgUuX9f52BnY7jsPpPkVuHikKOWyXC0PyNeReqZkYg6q+B/OQM+j7PmA
IPqeSb3GMiWHbWWEcx5pq2pCOs9cpSyjNqr/WRkBXGXsUVUVHXI4BK/b3XSf
ewv84DRdgnQFcUX/WmFQ+WvmXWj+9cOayf/4CoVWimnv0LdKLHLcK0mjw8PF
CLARr1woTHZ480tCFlLvzeJWkAa52PG2xhomEH+DAcYRsk2RSA+9sO4EAjrr
0yUesB7v/5GWQhuyi3+V5BR9pWvFqkqRsNg+tTfF8dCY7ZJYLiiad/97NQDR
y0L8AT9yXyUGEaBAz0Jm80OEvs5a1SyQu46pwfAhxr3r3LmQJ5ygiYJvUaA/
oH5r+3Zi7d6NrPhDYJdTFjN8KRVBzMamanwUHuOPCVFti4Bynrd0w9HCEmeI
eNWHwXQJPCCLEMrhdzYbPP6RDU5ttTOxbI2OtX0i1RBvjb3AH1tpp5BzhS6C
xuqa29XZp3ToLqYaFp6HeUCiVYtF4PudYYkWz/UdMwrC/Qu+QWwydQcGJnCc
f6yZ+0e2fnqlatQDzr3/hcY3g3w8xiIkgmQHN1VnKHswqHEmAzKVsRc6uJZ2
m+vi8dsaiSQS2iSMuIjINSWDUDpIzTDMOhzt+wzy/QqhfzxbnFHWtnZhEekk
9wuuU/4NyTifxrqScwHW33RQU3TRK1wfhWwYiexSyKz8IfOBlkfajRzKRrmV
ARpic4X7sPihosRqI1euxCAn58DGbw0jajYXPi9lcIWJBIJLUxOggQzKqC3V
I6826NoBgBdQwJYO8tV47STh2kIfR4Q2IQKTjp6LpPSrLcRGeb9S81KHjmaP
MebLgI5aQfUTRm7QlF3EViSJGGxmM8s5x3tsQCynfxQ00TyvLCDxYTrGKiEH
lhwLrTIy4gcjtUTdZ0rJWTQomZnRviDv11O8PWH8yKV7RmINENvl+CxxaOAy
AJpLIIJiVUdk74O9hNkShr7/mdDtpU0hA4Stn9xX14Fb/UfPKBSAz4WUYbd1
9em1osPfecUE0jUw5tJnYUAjpjiF7jFNnf4NRROdo3YqXNBBro3ONrwkX54S
AC/gHJoXH7wUFl9NuvZE3RMTI5iFMJESX3WvIdVXKJxRJvm45UWGXuWAV6Ny
fD/c42nZRjyAk6gKllYUzsvSite+cVSJZrdYvvhoYqgjYBw42J1+AuJNru1y
q8NZSzVNTagOzz/a4JRqOr78+Vx9urKS8EwZVbtAvqXQ0U6Q3KqY3PcoEmjO
pqsMd/Vq/B5dRMVSQ021efsEcRbFCc+lbO0XJjAf2MNo+xaEm0fiUOZvNEQ2
eNaOsqtaHHrbqvbzEyUnUdeGeKuITAiv9ykJHBZuGeQFyR3ReUNHIJ9AEHni
SD8iU2xU22NRiKHtzyVAgqB2pZ7tBZmwU8Vy+Vp9D7b+b71xd/Cn6qELV8sd
0vrTBvxb5yk03baI5NkAJZwUDmbOOzTtYfw8UN09izr+XIuv/SDSwwBBc+MB
G+lQQoxNvNqRudt+cNm+H3G5NypFdS5pNbgyNbZpmSO78SPM/HamBFP7rEa/
lLNlWetdEeh44bj7IZR6d+xQ2ZkKcw6Bgv04j4fIm2CxSsiYzekscMYVtmy+
75cbvyUzF2ZMTuCAhIIQwDoc3UgPXmyRxJuPGEX4OOaX5mDj+SNIP3OgQgBB
Ki8aNvljTZs1Ah1v6HKWZXjuG0jI2OHFdmwXKsOgyDZfES00Jr2cf1VFF8Un
iEXHvJ/V4xp1bGdMEg87J3fzVWsla5Hj2boPSIwj+AHAcXJgtMZLRSnrEWei
UPp7awufL3+pceBe4s8z+XNv7mgPdGkk82EK7Tej1A7FGFNT23QRdAWJhXIt
ToCwMwvLB9zY19KPng4jnNvkpFTmGdKB8wSFoEJrSNgF0xHw5gOx16l1RPmr
14s+dIt2pTJwf2oZFcUSIXs0GN6qt8MNTuqTk1bfazNP9MghskKUxVsfA944
JuJ90KJ4K5EZPGzF/pOBGHI5Wc8lfGFrrV4NgRPL9DikNnBVwnzOihgT5Z5P
lGXesGNqAmA8QuiRCrs3Mh8XJjl+GlDnQWuPexJiYJzs1nyqRSks4vQRnrhP
0GPzr48k2Lv472T0z6S4k5NTP7WBWUjLbXpzMOxBZ3wNIe0HzjpQYHz74nch
SQGl/1tI40t0Qj2JSQNVzHDXttgnc+erYEvqP2wNdBmnvPuk8U/tKY0cm3Jm
T4FvBATNIX3UldpBJ62Rbf3XvJLCm6U8XCjBO3PJDhKcEDAzohxYns54H2yd
RHdgzcC1T0m9g5y1TFWgIyERuQS3Rj6ifcO/Bp4lNMsKC9a2y803lRVJG8wZ
l2fMLmH/NsmkVTIBmu3fJ6Hj5W0mjJMXaVpL6NUNwEVurdRNYYuQPEf1NH+m
IjolHk7HZjsz6g/67wmwus7h3HIusr9MXttPPq/yg5r8goikVNp8mmDjS7Pd
hOAgSGxiRJhBkzkRe3kn7MpekI6J79iW6LEbECaf4/fCh72kIT8d0A9bf08E
j9Kjq+QGT5Sl1vsz/rJ5NXok0jD3KUlf9Lw9CPB+oq9Gg3DqbOq9EqRUaYVg
VWVyWZFolHppHPotu0sLr+Rd4TVbqrrh3cyp6vihsXFsaE++wzcszLzNqY1A
dsox7GbHuiVuLbm84OaDomwD96RkLTXjb1+Gtt8rGuzLNiwHtnw0x6JP6idz
S0kiY28YTfvhcLRU2wCcLT3lGkQ26PMdXmF1DMhqgbllqyXydvdWrGcsME4p
1/6qxoik0+9/i7ia6FHyccKVm2ujfP2wgbgvT8x81zBmMXlf3xs8/GRYQCfu
49VSiUokqzuvjUkwW1L/xvmO9mL6vFZsvNW2GlYqw/Q0tkyUniB6KLYgjxDe
MJtEcOBuos+LGS2EY0xzs0iLSUfo6WPsQPQbf/gZJMPgHxurql6XHvUTPmIu
14GieUu51i3V8/23uRNORULY0YOJlcSJHYImyLYch/lh5bJ/640KVWy0oAkF
0vxIiAhpkWPpL7p5Btb95sVZ8pUhUNM7IMx+dptN+UwMkHBTVoEzVFwPIoVf
E3tES61C/ecOhP89B9XAOZJSzLyWaOSVSDL1jxkJ9tPrkKMX+8yU8xUw8Cb5
H+vJq/TVGr0S4lvg9/31iZLzFaOgY8eN8MxK1adSlkZd6xpEUPuwR5ti1UcY
Rkxj1r3SN6VTZbxUKcU+Pc5kHTV0y1vEBRy8c0gfuBRraVdAAaecgcpRLbVc
mGB0ayI7PEtSYvlHiUJZkYxLOg18+d78N1RUx7QgGkKKv/4VQSEduy6HJ1I3
MI17u/KV60pJkrQYrcbz5BBrfCbU9IAs5MAP9GajFgR/M+lDJXUUwnlVte6T
09lT7CnIPqHs2+EQ8knmlf4RPdg1KfzBWdHennRstTIIYhp6ZC/mMpnYeXwS
SsdjtPlIU+wVMsLOs9zUw0WOTEzwNSNEx5W4UiuzWleFKaoY2qOaJKF5fPee
hqyy9aBcPM1Ge1/R/k4nVtXbkeJp+FFJ/blUow8AVhyHu/e+VXsHDTG3zG+h
VOBtd0tmnGAwTnwPqZ2oKM7jbLaqD5KZYTgy3lGWHfTnN9U1dlTfMdHYI+y6
p2l62w2vqu9HY4izXK5Sp7JVX/jynyUdD+8w09TtigUPgVqcBJVVYpfy4Gq/
qRT7f97zJsL3LG19ILOdTWc+fuutY8rkBStLCCPR+uCMkVbN5xbBXPD9GQ8v
knh54WavHrIWrqJuRdHUdZROsOCqWlYrBLwrtFHI/Si4QMxGYWg/Os1FP8B0
UYVICN8pVxiyzYqm8RBPnPn2bO8jO0K96zVBzPuw+IPVXLUNOsH9gR7iMZmc
2DIIRcXX4EqKk54WQ0v0izqUkm4bnhBaJ1znni07wE8MlIKlwER7wSIga/sI
+EJF1H93pRT5oL4X3zLowZYRGxp1QuUDEFyY+U7tqbFXTqPN0fzgrYLj6DWG
SDX8bIqk/5Vp2nd43moBbG+f/9b7i4uoXgWlfzhZvzaNTUz6Q9K8RHAd7zAx
UBq2csiWPHrBi9a0fAtjyzvYBXYvWxWmlW1mFTpDfTRwbzCbDvxVipSjezTA
py0gMCVewnvkbi9K4AI6KGwHDPwoAPPDtu0elgmnYnw0c+1QL6VvYy9Mn3Y2
fF8AN2nx7sbmpkuWcXmszlM6Ig3k/Jo0wF/WNgbX1BjAlY0qT+YRgzx1JKFK
hGRQlQAQfUKdaWCumypqz2j0qssRHCw001M3KljtYPt2XFK2NysDZ1CaG5/y
ep5X4qK2t3N6Y//c0IbHyzWBd1nSSgD0Da5jgMTlkiUdBJU3Xr+6bIR00s8p
mRhhlNmB9AoPo0GIwQtNwkCt1dgHMYoS1llH6Q1kk8XqRvLQmln9Hz7MK18b
dvO5yH1LxtnxTxt3b6xj1ou2QsgZ1nK5E1r0QuxslMvS2/KF6C0urf4BTn4X
U1vccA/EaRuWfjgGizPknr3kGlrv3uZasGoEqo8fGMlO0UQfHNyTokzFffAW
EBRVNuX1qF1MSOXymRZZunn/h9P8nWE3N/FszRpwKsdyA29SQIzEDSjYGNAH
OVOM9A5c993S0GLBolUCyIBt49doUz/pUB2z7u5TtoNcDq1ISCfZT5epsDjd
O3IkZXzqkimUT/ecI9cjW9hRcpJVmboP47VoPqKFqlIq3ZWL0itGdN2uZfiX
XpVPysJBieRqFb5EWS28qeD/h9/pjleJMC0S+EDEShS6ePLvIh7qgQNvrEHW
Z5cUBoKlvbWDx+rDZXwa9L2BZLJMNiB5VVku4ANRerCw7x/RHtX0eMAEHFEE
CpkebhMdNAtFMNYRRzN1T4YMQ/aeBBUZcl1kvnoG8l2gQ8c3Ti4M2Kyxcrj1
+fG/vxH9jNGzlGGzG/jlKNPGyFWBSNumSlyrykvnBP0EdKgEGQiog5VPslHc
YBYF3P3buasazvCb/oSB2EdW9svIGzD7iRA9Zts29n3FzZDzzt/OPpEpby+0
39/mVk1SHv6H3gZagH5DdGffIL08HRR4zjHXaAXHWf5Dx7xHDnbWSszbpqzL
tH+/lHEwQtdxKopcavCMGxJgUV4e7QscjZ31p5757KMK6aBHxFCiBmxbPPVE
lJKFvI8x15XL5ifpvQAtnlaRXEUkgyDWXCgGepnKLCIwyBCr3ptIep+YXFS1
8XKNvBp1pJtmrYP3BlCY+zTqIr9UK91q1ZnBF5vMGKABFE5TW9WTO/9CIGK5
ougyOm5TemZeufn5T5IYzHvu1j/nWdOMP7peER7B4t67zIZ8oKDUru3pNvA9
kn01Akvabsmnarnu/LSYYritWNxBLom2L6Z8NPyEJUrz2iPmpvWXW+ByBn48
VgIlm3p69DWhDiAi0bHsTUtuyyN1X6DqjqlZ9HvYPfv/E46oBQBaOBioijGQ
YS6Ih1ELjAkQQc9Z/HPMdrFTj4WNLU8K+FSkczWRpCVSVK59iwE15VfUEZDp
Dj6ByffaaYoz6i3rARWezt+8vXhxIPtBGrKkY3LM/a5aahITfKXplM+3JkUj
Wmcf0mrC7Wb+wAuEUkWPtqyg3mcmv9BcpcZPIn6qf2YNnDVtYaOwXtkK/IKf
ve2eIvlsH5O0k0c/yPYP3JhFceVyQvQoKmCGiOmKJia8vK7exxhT0s9PSZk7
lKwqG7v22tDsxRDOcRFVoTO0T/z/2Dnp1ZBV7i/eBeMbvMaVQmQTY8Hn5AW2
Ck+AeoAbCFAlhU4mqQwwuGMOLQVRhRsbyq+nW5rINJhPAf6JCkpjz8M97jPQ
2hDubiNHQfHA/mUUUvsrkF+9/oCr88l80YYzzJlhTk4K+n8iPtwsZTNP/z9W
4GJ3v/AIGQ2AVSK4ksLdRhyA2SXVZuCcVaKSRknMZNnC1n7OnQT3R4c48HvW
gF0QcV1EChPN9+ci/PKPehAFoTSf6An+MLUcDvVpelI65Tk3MJOKgFwdfbrt
MAHqU3olmNE/oGHuAqBBE/OxVdcQr/QuUDMy7RCwb+4XjwrHBQdfsvp3LkTh
X+S/K6QbYX8vbxbGmu9QnZ+OkxOCpzd3X1tUhzad2x68IrIJQDvmVJeR9YEe
7UwBAlLEKHbUnBjTXor3dW+BENWGdAD3Y4QBJpUgRXf42eeOn8OZ37MEb3XO
icMu1+5qpPD38KFR84mEqiAP7AXPdhtakLk5Tz2lb7PG/uizirHtubyNlydH
51JHk3UGD6TDA1M26wpDFhnLGBK1i/Rt3fcdT4PXuS+p/8Ij2pgz+zoQ2ATW
GluksYqOyJgQ8XhoyNqnUObPbEmY+gG06+bj5QMq18XsFMiaW81LLVRtQzvB
guqd8GChRydXz5WC5h/pQvwNIovfgIJAk72SFP1i30rIQCFaAXyEZXjkgmhg
vpZ1BBfEKkL+cj1bCY9MkNhwSwoukwud8GzlpaZTrKraB5LUcq5wqcWr7sOY
vFuK6veI/j9hPnUxuVRn2X4lRtHOZLSTinNJ83cyHNqTgFTouiGcwIssWcDc
SUcDkfA7HmS+ElKUCm8UuqXXuS/8sCewRc81EsgzttY105yNxc9Dt9b7VlhD
v+5u6+5aBSdjgVT4VdNLi+MnHuxtofeQ6+gdUKpYECVlfEeRHbjLKqpjLiac
kA6ROJqH493SzMm+bQyTMTMqWbrRvebNoSzoGEWPKHNrGzsvkhqDUVJuGScY
CQFVNMLffK4FwOkeN00C9D350tO/vhimEzF8oSpcxGC7r1NM+bDsVCRqQQsb
INaFTy2xSPXf+O5XSfLPy9tJpqlxbmVwID6w7WsLG7NTQbH3l/gI3AGSkRaf
5fTEmhzW0HDK+sRYXd36USca6rCMTiUKRa5NIeqn/9ZKKyqEBYDGmhpKudqi
3m+67Mw7BaOQ+1qUTlWz8FsAu2gCZTzbRaujlzkW8KHYEr6zMNVlrMLqiE41
FdbNB9YXGno70uzJCven3ZhZkXN60wLFmOmVVe5novRaA27eQaDpRhYQQ0Ks
laG6bPqlEUuQi6iZ1jG6CBG8xCZkSgLiraT/KenEbXEnG8r1+VX4bAL7AJ49
BO7IRH7gTcVO9OPq6vGi8CV1WzxI3WKY7+2FpdhrE33zWB/a2R0rt1hd/Nmq
dVivAh3gfK+HoFf/dW/77OEojWlURR0y6rQYSthwNOxkusP0dmXUpLPYm+W8
C+WM6+7ndeU4FiOC+0p+AGNLZ9wf3K6KdSa7abZpMnRtBqj5YHPToMtfZTQi
zQB0Dt4Wer4ZYH4vnbrLY/Qc5irTlfbWbI2vAk4ceVrkx4IT9nKfHhDfOFvc
c0NGhx/vxqdO/1SCTisCBa3n/iZbYLItv9S5h8cGxNm1QTWmGw/h1M66Gwnr
7C8dFN1oA+l9Ntcl9eLFS9Zuj41ivMqnA09eM0up4Vd9SWDwzdUDTFYzRGhe
erLcr0S0JHF7Q6XhDYliIfbFLcQhq6pvs+D3l5NEMJqJLoVqLe+7NxDFN0uc
Nc3GutMzT9tCNdkQCtk6TUY5qTjS1rbWHl5NomtUL8lINZxxyjXGlFo1e6Zc
6sk7/vQE7pxU3rawbHyHJisDgRAa75cyKaBkZ3G8yHgl+ZzJdMOJl7fqxJFV
ZzgELiLYT/9Sumy00AUx9+Lz5hnAuMXji3dlTeUVIxSMP8TefZpOzNBw4jbh
xK91T7d4jwP9X8LCdaqoleSKrktDAI8mA6Ua8cQvhEv2pM/IxdUWzKruJKGI
ON55U6ZMh4vxKgN8lt4RtlepxwMXd7K9ogk3NKSFqn/rCQ+C+0b7h2UjBMZg
RWJOGS7ag/J9wyGQZck4LCYK6rSpDUKNf4noZxhvC4G8UdWlpt37AiiqS7Dq
4oFTYX7iEhxiMFw+NIYb3KX6pSXyp3K7H5Kr/CjOxMk8DA/zDdDKLiuZx44C
i2kU40lHoc+EWufmD2a+VKZo3Xqn8NCDgo0fBD7q7Mcx28IJreaIibScGT2l
ZBI22qqTXhxrcB8oi8mUiaAwciHdIOdpHhf4TdKBbomZ8hmC3CXsyUc5P7HK
5jFuGdixAtT0iUfXR01uxUlxnmeo4M2XmDKW/VB6K7qowJBOTxEBeHWqnGg8
gtkE8zN5p+XqUCfcRbmDxYJyaqkhzLw2rEKsaM/4cMuClVTT6M0ooZNlPI6L
aDLjEpX149G9Dcr3pQyAA2Ft25TvPWCnSSBqHC1pJSGLctk3zU6qt6KJ79qQ
auCe5VuFH0zt9xqKir+SDRQ0j9+Zz1u+hXb5uSOTzN1rsSpk0Js7FU97eh7e
nhA+5afMbUJHmTARCnnpJDLowVdOhQr8/bjbLYyHA+SIHrhzGVH5JQuz8DaS
HwZMzerTMmhUA74cYK+DM9h+XB0oQLIiwsAN9IRhBHc479RYBn+bUUKZgxj2
0JOaHQ/eg/iIx7SIUWCEVWts17F2lEWV7Q8nCUNsZs7/QYrPYz4xltvGa6bI
XrmYhRHt96M9iha6U1fN4Yh//OBo7g1TrfdlxV5OBlci0K6Ivw9dN8qU3s6N
v4OrzcyV4cpfih5etLpnpesgiSFN2y/Bj2gQ0aQBIgIq7UeXkLcUrNRULT4Z
6DXrDKISV9g5cISuw/HpojiLKbRsx8xDzdYmtg9ixlkQqmTEjpGxaCtJW51f
D+G6iFzugxQDrfaEL0PGFAXP86xwOIMUexfX+s9cIjpzlQOBbxwWoLZo/aKv
JhUzXTbPVKmXyhTStVXliPmUum0pGycP4MklFaEl87VPortMOh2c8lCmVwJ3
1KCdtDwAVwUqiDHGJvy49b1Mpnzs67ep3iCSiSxYLA/FjUf5SPi84oVeevA4
eHKJx1jjT0tv+32hvuwm6SWMWz1+owmt3Rj9tLTfKGZLhHQHenNqOFrfN/Xc
v8r6z5ArQbH1Aez6F0/pSdz3/zdaW6t4okz0xEjUxz8kmiHCQ92nM6lXPWym
PzSgnDTRkWjYs1/AvotHXZrUrn2oXTPfk4GxtpCb31iHNezk4nruf/VyM3aT
AlH0vSjjZnbWtLwiUqIEd1z7fdlRF0qudEj+KsPnMvvt2w+fc3eRkUhXjh/G
5Hf/+GVXLoYhHi+SbK8W6ZqNi8TKboBjvJJE2kTH+NRRW9+fiKybwf123jtg
ZSmWMbFR/WAtzhsD7GF5EmGsj3qktmdIXjlVUEobTTepCknkT9QXTFrVZVGH
+LvrPZkixuNdcqNrA4/NKLbzzaec4Lb0jZX/OXZ2IMCRWS7f2pbXKxzm2gBF
Zusk6wb7r9juEj21xIIlTCdaMTxszLOE3YFPZ+n9JVA4JghfEP2ld1FWeWLP
M3ZBSbPU95Zs5eHuqX4QB3C1QyTKD9DfkDELMYfSzbW3zCByP7TEzEXjJztc
aQbACgxM/XvI+6R9T8y27F0jYHv2XMf1uH4uwRFyYB0CEmmum/0U5DKsPhBj
RJMTYYC1Na1jfq8JgfLCU41E0Q6a0pzGe8lQJmhi7xjvKMlIk9fCw9sLS+ut
4Xd1xs5x2ZU8iJc76/Mw1ucOKj+7kwhKSStcTg7cRhoBdBLwYDsRchDJE+nv
YgKxvoAlXwrVH1yYyNpF0r28aNwoHfrDLROuXOotkh5f0+ZDoWn16PkIh4Ul
X58VZut0L014IdlxloOBS1dvNnuKOUeM2Ck6Xy7PsS0ZNS2xvByvV77n/1Fh
ChZxiF2QgD2U0CDfH0dRgt9kJMDLkv7D8JdpYApUzbX1EanAKKIgUk+lPGau
xZ/jcb3i1ozyxWnaSg7i+sxaJYmmZObbyuzuzXWQP8N4Ziz8clHvTREzXclq
v1xCwK9KPjplh4NI9ZEVKg972gTIZau3dNyGO7uF5n0I0ypWtUbJJO/akwD6
ZhC8MvIg2Dbw7e64j/f30VYVrl2IZVrrOHVivtlOLnc/h8eedKnJ0Go3lDe0
mLTfRbfyDNMzrplmya5Pg0A6rK5lI8WiznFEw5bfqDWvAswzQiQOHugW8soW
dC8Kp6y8gOdf4+3ZUuUzA0NST+8TSk89RV1fW/KtU+cE9vvDrObXH36E/Ztt
FhD4Kptuf+Mu56CawKf3HbvRVGDPpi76ptCbe/8B54D0Fd9i4MlNH1Xb0Wet
P6DhF8ReJiveE1DuC85Ywvq0vlH4MTaSr2a5BTeDd3cozTRWRL7YxlSKJX11
MM4Qgg0L+MYKXxplw8/KUso5FhJCqdkO289Cp/mgVVDFbUXWUrke+kbxussn
xh33HxSxod8VWWDm9zh/C6APNXbFqo3yG/zoKqI/gmk1qd1V7h2RnW79h3XG
Y++zHF/nblHFWExcmFiieGC4P05vqJEEftHZjyeFbvSSWGwe+F0zAAj4oqzf
c3vzyttD+8KBTQ8BmkcFMxgk6jNIGFGGQGJKD4bMrnNstHUGMJE5exPv6ebY
ZwjiNJ/bGHYZNQzX+YPJk9SkCl9LmY9PrF59AROEu53OFSrZMxJwrBDQmXDN
xLW09cqBdAKB96eQFRDCPWTFSRX/evl9NfB3CnQgM+rAKbr9FaT7MI9BGlEt
OZBRbmg4erDUtWhdwYP9phReJ580066vzCLfffML55UqWcSjE0TfL3Chnuqb
wz2FSOvq2EziGBFWAMgwBtE3cMJ3UK0bD5QY2wMTwW4x1MCRI91A1fGwKQnJ
OSc4yqsUOnLhiUfPwqzEggZXSHxqcxqn2dL4N4ZlosQ9Epx7LMwd9rfN3IuF
EengS9FSQT+b8kdvhnDzJ+vXivjiWQXR3hiNESOIDRilcOWRiu21gzRqVc1w
GZL7EikfKGVL6kIN4908WhpytiyJPCy92/5TQ6Yez2U4Z8MdOUq6wDxkAnZ6
8Ym35rhRaJTb4QF0m85rsx9O3ozp50x4pEGE2C1cfuyXRAJ9qhfHqXIokESI
fPn3OjrOneFJaVLfEpI9cQ6ql+4/qx7xWqa+PR2f0fzs4VH3OnEl7Q5LMwzL
9qRYhRGIVlLyF0UChT7mgarBBUGB/NFBP6Sj7mZsee9a1teYzVJOurf9NM9P
jpyAQEvJ2ByFH/kpuPpC+t1I6F65k3LSMAy0qYMJ/kvnC9OTYW/g7DgPkfo1
8yQDvE67EG9HlcdjOdY3rPg+2HgW+SK2yaFCDZ3dxGYurFfwJ496UXEM0tUp
tMKFv3ONFbwlr9CSXhmXp36OvSrd314/cDYIeRHXv/TVwSQdL5TX4UIKNlLi
tAqchYXck12hPS+XyDKP29PeI3wU6EF8c6Kh1t8Ox7SdW6XY5sQqykeSkr7J
Y/ugiLiKmi/7J3BZMREdRlM4efL3nRXtMSw0SUeW28wdc1/wMPnfGutFOAAZ
sQiRn5C9iS1UXvxyqFgTars1nlWTR4gKrByOeEmkNg0bBP1LK5I0rcEhiB57
tOO11LkXiL7of+1Mm+C0R38QXV8L3K9gVop2QCPTGs2raWqktJPvBLB61BYk
5V1qYODH1iAjLwRKv8kvL1dCOw9Fp7xTplnDg+OJAvSLBt1KPZ9gAsBNmanQ
cR+v+3rRHMMD6DcWm3jSNTqOcIwXwufqd5HbSeyATDML3QH5z/9q0c0ZtcCc
4J+fyoZ91tvjBmD/QZm8fTJXwZeSOx2FAha0fmdMan4BnUdqnxDmZrzdYyE9
Xcci5/xNfqsRnrm6mJZyTN12tD83uXfPE8qqVbCD6ZxTE1/vmCezgIyLTs5c
LxHzVPTaXuDT2XcP7ijZOzACDI4fuXWUAyaY6A4ujwFinnwESyKO3v5Zzd1o
nAWBhXfNTFwGy3N3EYLjkwynqGRzc8JzKaTT0qxTq6p9xoEW8yx894dyGOfu
1mChylLTP0s1WidbdOTm5W9ba68jquJlMNgd4kJWOXC2+B4XaoFv18DRSrTF
OttbKP7sT4P6GK8LfQmWsNI/ufl9exa4GG9HOtEuIvP5m+i+iIm1rhtjzE04
iunn09zjTVs+aJNgAVNFAlZigr0jDT8XAFaPZuQGUAnWp4xn03niJfAJI1xz
lyc3b9jTNowM/kXfvDv0ou7KWVohJmxHTI0n4SnNA61Bi17qPkI7rtnqh7LT
tNTHjR10sogyxuHTiGdq2Mf1Yp6n6P3fPW5TcYomQyte7zogKF6LZzVzQky6
+lefU7Oc3IEW+80ViHmj8NmNDUNgNK0KWoCftgBPPbVF6odQC7aHwAbHX3hS
sX76LrPJF9zm4eOjknj4WEtmnb00FFHvbbY2/abhb3x8pKfcRRR/5+QBmMny
eAb0aoyyWL1J0WHo6x47v3CNy6Vdjw552jO0vhCHlhz80cLxmop5nxrLzPi1
KE7uPsOUZTLgI7JSMJscQkM4gVsX3kKKeWcL4DsIXKSXjFJj8uar1gi0mOO1
fzMLHSmz6wPeLO1oac2NYgebiDCxTMX7iEUJxr96aocihbm5Ic2ozYjBcvPE
ojO0g3n+6Y971rwM5/60M672GtWBYlrLhMKdiXiGHIMN1hqZaXgqfE3+fwQz
s8vqNvbZHx1kO3Q4CNH+R0SeZz9pss7TWfygzA8GS4cpUMmrR1QEaIr+KKL6
KM4m/RyjPG3CwH+oE2THXH7htpg8zc9GiAC/ZdrCeFJ9Unxoe60zlUwH/iXh
jYQZVU+1qu8DDZaa5hlE7D4pq4mTnDDUP1qD+SwRDYTqv4OPhKTpADoDG9nt
kWWP2V+ggL54JoY+WZR1uyLvIsKXxFSx57LLhOR935nM3vs+IiImGnEf7Hok
aC+5NCQTO7rr+e8liP5pLXBzImAFfnEc1KJi1m0uUrIQQ8I2kyHvCwtvjFI3
m16sFuHddOS8g/HBIBTHnbTpzmNUjujOgsZfev+r36XWigNKj7M17GVmBGxk
0XOBdbmn/GUBBbPCx1DiazWhsQfMnT1mHHUX3BAmuOrEv09rlAa6DdyhshAL
ANhuwA+m78gW4TjwsW3L/uIwbBGEa3J7nioUhKaAuQ828ipaiUfpTxEDwsML
y33rEoThvWcbr/Yu8dHrkQlO640zRGIC5XzNaRFQ5s4/7nQWCgX/LkiG2LU4
s8ZhIW0UYNtsQxDVqQNONkgE5OlvlZiS5006WGzdlYCygPa2f99JRgzpph2O
CLu5V4vlUX6IHV6xpPd3peFZQOak338cm/P9it+Yu5xdHTBgZYBgcD6+gG4o
5z7MD8Sppl6iGTzJ+IIiznLBGAONsB4LZts7WBSSYaYImCm+M93zQeoGEp3P
xACunOPHYBZeR8eILl6c+G47Fn/P4v8bbyi8ieYcmJjhUZSOfZFXV+EPbHiy
jPSC2O/vkWW+dIQgTT+TaEmUEutPMJUCX5eJ9WbPhCq3j6udhKSeGA0oQItQ
YZbgkNCDH8nUh4zCxuUgH2irhVSSEYjsLXnrWYu0yFErzMzGxyQXvwDY43eB
olc8hNH3Zd1sMRigExzFzUeo/JoDPXqT/QFIiJn+4oUlK1tTlPuDkgpJFivS
KSyNihAaV0qrx7F1seH2znIiP1Z7TjKNmhxTbLkB1tTWM6puEQC2O6zVVVtf
8uTiWYPP/tVbGf2gdzTbEZUW5lrxMXWJoXEbgNk5G6WS363VG/mirL828l0w
ILvx91oCQvqxLyUogZVEn3vYbn2j0/EMK9+Gfdv009hiGPxY+Hy4EoCUUspC
64OQDP5hyg8A0nyBbsvEqziJjuPq7zMDgaTQXyx4kAiF/LY6nokjKLKYzkFq
tgxe0UhA5KITfccoy3DIFmeRiiFmPSZkyjaeMTahBGtFF/KbAb4DvP1PFj+c
5eZFc/Iyx/IsFOtE5s0UsjzJdeIIAwdWXZuQ+9mocZgcXdvNPzpFlpfdeH7Z
Om0nyrb2WhBe0eWdgGgugcBEWzvUnVG/O2E5v380ohor/Qn/MUu/XALwalFj
X3qvlZV6IzbpsfSFBswCuiAwXdvh0ucOqU12WYHNphjYwklsJo4cpot7mqPi
UvaGJin/F0jkzr1JMA/L9VTxMx90ysCwNuZ7Hn2dRbQiEzMRygF64uupz0GP
8+pxBKtxFGZRrZS8A13r0Ewmzq1zuygSSlk2J+jvOIeuLmrYaUscCkopFbyM
Pelb/w0L7JYTbxE9AJUXMnjVlm+FqeKghqKmG6Rs7wf5Y6Qr/rPFgHnSJyij
k1DyLxdYvXt2HEMu7d3ySThVWx5W1U9vnYPsS/GGti3LMVP5m9WjXv64Mq8/
Ps4qQ3l425o+A9kFWXIuyV6yp6FzJgav64BD+mBbSx1kYtzbJzuOYIU3794c
3B7VjoGWTUnBHm9ZyNoAVeGclJMy7twBDD0jCuXh7tpBhLzjibClJeM0vtUr
EGZ5I9yIn39BRpSsxgr1uswHe0uF6AWBdpTo90O1Cc3+eZ6wqnBiRud9xkwx
l7HmwB2dpn9u+0OUx8EzMiZNs9MN5+VF4h8Dc5TkeJRqF6rWzyZP7JzNB1GD
RaMq3GNqnn30ALoly1Z0UnzX2BkD5tW7pnEtrwZFIQtmQcay1cVlq3NT9ywK
M694XthJZfbB6RLYecpggxpAtp4BbII83iJCJ9eZ2dJJIxPgERRkoJX+gqLX
GThXpRTjEPoFM61uVfJNgVxXiF8DcqYi1DU0ZxD7YvAk3PWi1KnrqAiIPGEy
WU6BCJ0gpPDtXXJOnGN1pDJCFtsrjbAACuCMympaCx31eUKk7AFIZ2Rv1KB5
vzjBcemllX/AWVVJCHDdB8kUeQDwJLNFKiFXKmDHwWke0BHz4CHlOGwPmftI
UVj7AMDh35j0SZ32UY5YQqMDiedbYWT/wc+HSlh+AOB86wH8YkQBusgxhjWQ
eqQ48qaFy/kpqBP/nD8KnSFb3f2/Pd94L8QjiS65gCkkICQcwhNPpNj/H0Qc
2z4NCrnbQjEQmPuTmVcYEmCL7nTfcDwHSk3yvmuw73Abccsn39V+reOLjKMe
712fvxf2W56WWHnnripmxIZg93zTb3JDdOc7UxxTetTJKWmZofZvbPfnLirV
tTJgPYyb3R0LXGOWUtD2ESyPyoqFGdCl4jQWnmLIxtcFkqbrCCAk2MbrpVCN
86WA0HvV3gmce6Ra8veze1Gr2ytRKLW7+SxkP7Y924sN7vMn2fAElgKh4sWy
dS5BIlMzNkQYOb4POQnMwrxYXv+6A/Lpi/E+KmFt3wa0JGgCXNLOoAR8gEO0
7moRBTWu65CU0nJpf4KrfzWLL6tM6wScm50658US6P6M738XgVyQIG78bVJZ
GS9gj/dSPMTsQTXMlXQQtO9eU4pAsoxdnS2jWRfEy20fIKlWueLMkS+OZSTp
5LUIz8Mdeg/vmx2jzZod+pnsbz3WJPJ0F4ioXu+GOSaxCj2HJpXATpVG/vel
L5r9bLW9rZMGQHrpmWAuo0k0RsN9/iokba/AK7nHN2z/P/S2GU9xSyGA0wgM
L53MFGDTf67MNOi10vfk1nCWoDuRk1GGjbAeNY4R21TV3q9YgdibAC2FbSAD
Nu9uFpPde+mxwsr2aEacEPSB+WFfoCv74iPQP8q+kEPtx1yAQrENWF6wDSFj
lJoPYuobGfaHlZshXiudWsiGMtZ9hLmg4UVYSlpymdOlupLr1gK8GWX49PDk
VjtULXyTdOJtt455cGEbTlIfHIGi9CGQD+5XKrEs9ZzY85Zs5O1NxN/It7eW
Hwil/IdTqC7lAd9pM8a9WO+/eRWnqeBU3KoXuRdq4h9T3k6wRnF980Ol/Mwm
gwhI94r6cmzBRL6kWj3d0Rgmy4/HeR/hYanVyuvw8Tq62EBvUvEGHL2nh2A7
HvBXahPoHh6KjyRavFsRH8u5zJB+cGT2bUqtAjwc2gmAZm5pTe53XjWFwvo2
sSvHoB2avpcQ2E3p9JNiYkR3VvKVC16qZNz2OqjST7T6Q5ogKiCGlu3wweXa
q87YZEih+efVtnlxT6dUna/N0QGz4A6Hj4rxYx739Jwf/VC/vvN24UTvYnMo
4weV3Da2no4XFvFWA0cBxurl+mvkA3ueeidFcydbtS8ArmzBlpaE4n6D3kQt
jlkPW/JxQVPIQZHAYOKkMT02Ag2n+DRW2G48UYujIpaJLXzm6L1M6bvOvgzW
i8ejoEUhtp2KQGDw9AyyMBnkWS2KZ5MiA0keZ+rtmFPZIKtDBuqYm5nCAGxL
rFshlyzlVKo182mbr1ifjq6boEJLDXEQSU92EHI2vS7GVZFVanj7SzKSynYr
CERdqW63sQeGbcm+dj/Xm+2+r1BUS3jrdywb2ZXPZ3XE6WECYyVo5TY3V1pA
Jw7w+d87yiOlN/R1A6jFPOKfS1o7ol3N6ohVChHv60CO1UB7UnWhVteZoCOg
eaatpDR0fu5b+zgZxr/NSPY+PYPDaufuEBgJBtvOW5/oWMSO/v2BT/GnUhvi
Lp2OwNkWdd2F2VEhpNsepZDpOo2tb1SNRQX9iGlA88WT68iHLzw548ieRp0n
Mjn1F+quLfOpFmrOq2CfnGGcNcmHSTsR4v0GR7eqw+nFyMlRcAPRtpuynVvn
D+6k9tNAFSK9J3Pt3Lcdf7eXbdHfZvYt77wQhF++neTtj4TAzPDYoQHPa5+d
w3b9W2edNeJogxFdoI5JPs82fEoql/V3VA4McHu62BmD+eoOmZ3c5JEEit5W
qEq7RH0jvy0wEei18vImxwY8RYCIblAA2mfpa8yNAhcU1KYlBreYqcvFxyI0
mDLKboVUGJMhXBNQczRwkj9vbStJfW3RkhvwMGW+4wet4U0SUCTlqwhpZn/L
prZ1hKkvTUEGiUDbnyrg0cAuIwwLBvyLZ/QtFb6dQxtnzu64oXauXBwscIJr
jlndB9ux5XKQlzMi4MM6n5z5iCVPJbtb1YW9fAY30rYPqkGU1llv0YOG5uah
NHGxaUwA9STC2Rc0M0H9utABQx79n51VOIL0MRe3H/L5C5GcNyBy1Ah+Fjls
jB+nhUGbpfMHTwha0aXynTeDyywmTfQzo2g5qm7T7KneyEEsUdT8Jn/bbkTv
7OV8THYhpJcVnGbJCeqTVHslhEN0CTqHJ4AZtXokxSZJmaps/llbDuf0OJ7V
GHAXpDc7DXKn/Vjw7JjQ2n6wOxIn/As0nLdtBANRzl9k2dMnk5DNKo9iEArS
LJIkD9B63aqfZDJdVE9G8W+Z48bv6w4A2DbiiWj3elnUvO70213Z1ChkK24J
LWk3eoeOViPZw1Bl6h2xS6Mh9cEtLjNIGlXp54IhN6blqf6k9tmL9LbZnMYp
Yh7rdiUkeDDxkyXmfovZ7vDun2GNYVJZFabRL8vg2I/G8btRDpyt2hohYiO/
JKYQvD+Ui3msXgW3ZkS8bhNptBl0tp27Tvw90X1S93g7TCq6iKD3ZwBc9xpA
BbIxPQx0xaFlUiXvTxLUOP/0SUyHMg+Ux/LDOS7Z8N+TEoJZfao3kojbRgS7
UAkhWI7/e/lsfw910E2xw/es8mKKktUHmNwnAvTa7S33a84vAlyXxviM1vKj
4E1CICxF+AOMPhGD755fhzdbZc+uXj9IO6AR7TFTdpi21NuIUrUvAjr76P4Z
WzENdZPDAkcbZEr5xhEDCQhLL+sApCe9VE3MVXywTvEFQcdb3dzM0d8vzXbR
gdZ3JA12C+n5cUqqP7ZBAld74yjGVnELGe3ivFqCuaNiRqMxsc04jQIUouFy
1IvUyjOOrrJ3cEn9c6RoT+32j0dbcg/Sc/k41OAjO/TU6b4bhLoYmQVgIxl4
SCp5bvpTJwmRWkQ+0zNXmtmGp9d7CSW8+9T1t23PcuvSUGcmxh6byZ5SdOEd
yjH3GfrfoD6ZfakKxX+7Z5L+yfgBOWtknvZOvrZ2EumcQNk4SNSeVSumJXh3
GFnIZQS/sxDMXLyLQcZLBmsWvM8Nw1IoskgqSmjV47HF97oJ77s5H3vVXKFe
yvegpt2M6Bl/HOwPIX/tmNVn44qB8MqsAhedsDFqMNu6gnT/tmyoh5CgyMAy
4ffCHFGXertZ5bzEbn86lVO/5K+VMgg5ObYkIB5KcOkOXge4ksqc8P+MHBk6
SXwiLY8AGiG6ATFc8HfIW6ABfdwZ0cJw8n86Fo57twmXHUJHZRAi3qaqrGnq
vvAkAZlC1KYzzsRi/BMeXvxvvCbs5KqElMrPm0yPDr/kcOpICTPCSsBk597C
lmdn815MRsqYXHBfsxG2FqJf5G3HUWcpKsDwWSlVXFKCETM3kG4Za1owgwt9
LOYMb8fsTkE7apzhX8D/r4Vklf/gx5tV92s0ecdQaPnds0rZTajvdSb7APVv
FWHUtvEY1dapPricFqfQg2jde07Qf/dVKsCIr3qcuPOB6O8z+GiSaLucfQBi
dSjvMPHYzT8mY4UCC17XbDJe5EpyRLQQEuNhKIrzG4DQ+0fRnyQJAbtxLUzB
zUjT+zEK2kfsTw0HDFNHUi+z74cBeUDVP5rTz57hWQbjBlZ9ytqXSnINBHpe
pa5KRo0arFFOV7Cp3kqtlyQjraev40GLpDs37diwwUGMbtfAtCRasoiKLB15
cNnV7buEJUV1cfsPn9MlawC5vdVgUJwUBOqEs8nD4iQMgUimzqvdiv+hw14L
FR+yL2qKJOuCjnkSmdpUtI5tYr3ZI/snB9jsbqF7oTtz6jYCJql/X9UvPlar
Ypiwzo1hKKA78ziMnKRYwM+9zc1UPnwckHjpEVS/K5l9VCcllow7HtnhFWlK
wL+UEFuh1GgKpk169Tw28QP29l7X7BU7QUE2G7KrQG4ytxhQ6ewUa5e1a/ZR
aPMY5vdvU+2IAnJwqevGFD+vzIjQHwZtydNJTPaVCSg1Nqpj1Wk5SjSq8n+f
gW7XEV+6PYQPHyUUxhMpHQR45inzLeo5Su+s5QPPza7SOYRKf/gsvF5v+1L9
KHatlmnQ4XyT6ofB10lIW5v0fCv8jIgAcjhsJ9Btp13rMQvpN/dkPfFFGW0t
rCvX0VJGRhHtk7x1wSIDT23QhQGE87t81kyJxriwo98J1JHq2xvvp5mYy2iZ
n1AQZ5k7eBllFAyX3T68+v0BqLma9+vyk17r9RDApM9EDS0oa5nIxmzFgkg7
zU3lh7m/JA2T3gZjBUdMwmfaOOJWasggoZ27jrozxkFg3DN+Um4hQR2vA3k+
yoqbh9+b2nTTQgsGPZJ4wOQfy6vFc95ZeALDTLrb5pUIaJsyE9fw4aQ53+W9
g0pb4pDy8l3T8Ie7XVeqk0YIv5LL/tyM5zdgmp8hFAaf07eB9bGnCiovvtLj
ZmjqRduevIjbamoFI6IfUAQ5swghfwyePICT3ntNFICan7e0mexO+21iEf0g
ds422xus56LobQYAmqHqUNAYf3Ik5mcGUGAhp+zrl883cYRAG+FCrhh/2HSU
vvPA76HElO464Zir4Q62+hGnwtnumXMWXNc+anIgNqJJMNOta7JEevd619gN
o/SVHxa8e3P1QJcmx3UvLqKyqfGeoUfAurRsDKXcFMSKQqKub12441fAHgV0
6Ppywc2sQuLVZh/8pzXlp3AFHqxKgYpweJdUmVZ3w1orDmwNUOWkUdFLR5To
YuBNBenvM6+gD/bOX0hUUuxd/kdpuwGg5XReXJUZo8oK6IkHwqFQsbj46yTz
0KoGhLEuuGo0yRlUJFZhzlK4Dgg/guRZV7pmk0Q/GDpjlq9Rjj7QULuDyIfJ
CpnPhIU9gxS0evv9ov4y0RjW4WcGqiKffFdLa26ZvDx4XWZaOvK8GpJGYunP
BZqQK5WN+BiKW+I/k3WIXGDFBgsZkMGniUXfvKYJJzKlUFXxqPdNEneUjMX2
aGZsEPpx7U7OrD1WU472EjXVrwa9OwKXarwZqgEBRkoTXM8BX3blqPxaleV5
rc6Px8m0ZtfeOuLv0GdeYXbp+CXliUH4Acks7rLawYVkGuY6OKji3rm+v5Ek
YLA+XMF4uBDeTQWAA4U9iHyn//OOVvb9JQU3hQogFs0nMFR0aBeQcoj6bOzI
DEhqt1piiTNC3FTfcCeO78YOPI5a6d5ZcjyjpA70rmo1DPxaKWUcEuWU1POF
9tlFAATiDVQF9trr/drKdin3bwUAltDRlIlJJgWl1b7mPf5GJ9TL17XUuRJd
BjM5quSK2HI8krBT+5yDGHn41b4ZXB/kqBKRZvlQaLSEc9Vk656t0vRdUxwK
zQFmPe/rOr3k7nm+FJUbI2x7TK7IjWSZCCbbhIp2TOX8gHefBuBHomloH2GY
eHq9QQdtATz25Uk2i4JdMBIwVIiIzBu2vJS3O+XtqqgtcwGWcemKde67QinZ
xrQNg+PapbY+tu72BU2JD+hycop5VlpilBn1U0UlAiwhX2a2uqEWwzhOJflz
pIHm3C1m2+6V6syP3JQD1jRxWIGAZ9e9AJ4gosV7q9yUqNH3FtCFI//tt+v5
XdLJbDR78zfYzCEHb4LU7M+gsGqq9pvlrtS4LogBpCIIETpEt2n1e3QRcTH0
lc+4UD3wIZy7Qd1gB2Z4P9dK5Sd3LDYNnRVD0mkgzGWGcJPumiuZhKopCRIK
VIaWQluRodJRT38brV07R1zQ1FoV3mPmou7cnCJkW0F+i/fZP03zI91Ca1r+
/iqoK6tFP507MFWAlqbJ4DJ+y7VgjA2NPRK0Ul0B1Phq3TVFAt6wyqf0FNpM
kvyxxa5t7NYlZJ9W/QSOASC2URsmRZkXN7wirY35hcIolkJfkZoLhkaVP9pR
xG+gK1YHMvg0dFrBn7Kf3zDyWBTFOlOG5C++m7PTbSokRJIqET1F15hFZfYA
id0CtyVIEgy8+wezIY8c21JMMp8en0U+aaW0ptS1TFu2Z5Nomq0o8nMqTvZx
+hJpnq4DSDk2D7gaOnTOldk8VJejro62dwlTNFodHuheory1rSghVOhLrwki
KMK8V69HvsmiN0BxpEqbYfKOBjT+XhWVIGyZTahVjibOMqJzcc6HzS2dftmQ
1pEG3je/fg6HG4pNEndJSpI/+lVQEbSr5PjGCFetzxCwvRfFlfzXg/UBxmRj
G6ZIIqNtyYC8iQw/2GLt4vf0mG6B2FllI4Uq4yacFKCPyI06SBfSvV0TgcB5
mGR0Gsqj+ppe/hsFpBPoK0RUwnhrjOVhEaT3T2vyOChH/46d/Ymp4mDh7C1B
dGyOEZ+LvL4wp2Z6y7o9maap/oK9c7bIqDj3NiXJVli5y7OdeVoQG+qu5dfA
+2/6tl12gko98bBCQ9qGMY+PW5OIrb/GVRnsap5PP0pjxXMKzjSDUGW8nac1
UGzm+xHP3uvmg6+Do4sinWOW3qTvfYfCl/xNRc4z8E+Z+tuHfGuBRxPKSQRf
wenx8Y9rK+HSkSIPKOclNHr/Ur8hAhCJhnTOFZyTMABwESHUBBoh34o30CWh
YPPLZdWOt0rrU4xpPDryX+N0/YDkEfRUXm8AJ8f40EkCdWciwexAtWq3u1qZ
sOtE7NoEI97GOFudt1sCgiL9HrhiQvtefYbJ6bx4+a56T4xk8kFvdd7XGV8I
hlo3KrVzogCZDS8yxu/vzMZgk7ws/1bi55AVHheH2lLznnGKxqJi3ZonwQPk
hKNspHwaZxd8Tu3pNrd8hMtavJ3KlUZke6l/zkTa4lcUyqW0PFEqH8wgJw7a
mjMtnZW92pBrIiCOl0LmW5YWnbscKrrw5l1+UrWa12VeHHXLtTepE3ImpCYZ
8B/o7mrrwqIZkG0Q4+G6SDVFHBaURRDN/qldGkMg4frAWZrXbKHEhy4VrwfW
puDw+Gv8CGnMnnLEzsIew9ej4jGP/cRP/y8ypm5xObiaCoVHlffU5jhsM0ez
2LQr03aPVglDeaL0/ARPjW0DW8en20ujyfsWdKngTMFmumIgg2+6ErWEEYfW
uZCQM4ofBvpt4CMagmBd8yWozTLRl+gpwZhkjRdMTeUPhRMV1r9BJ44/kkSc
8rK/THCXf4w6lTzONkMNOAClEcmx3nA7mkdESXnISNAaaZHbGzlCchwvx6PN
gO31JfBb1nagKn43XsiLBp8Ht1YZp+Exfr3nCqEISEH+NRIaMxWY8SRZLjt9
gfIhUJaVjRu/+kSam7tC1DuLyg3xXUztyz4ROex+FtfFrofW6uwQ7cdFOK2/
hKZtrqIgO+2Ln1Dr+kPEDVFtMyyJdLmMR6omwa80+3d/TmVLPPx/OiDqX3/+
tIB0vGWMEEr5iiWLHYqSmwD3JODld7FqGk//4qCeAje6cba7r8vlCcuomRea
wPgVZQ48MuX63bY69nEBmeTcdEeg8e+mCGnz6heQqrv8QD/S/TlqhLIJDR+Y
r+4oZwroeayiBnMI6ligqb6CNBsZ0DVaziJW99/fsSh6B0Lvy27133JoJd3X
uGUvUNdz4rno14K0d8NTWHP3F4KKNHTYTEgLDXKYmEAWfpXJXMsHDjcnMJl5
mp1Gm635BwtCocMEpPe9HeWOzSzzFCn7O9/Z04IeP53zqO5Q6XFMKHqTvySG
e1L5YsNVNwOcfcTK/oRUwQQQIyOWkMMT3MTm43he8tM8POsocWnobhA70otj
4WmRKz7nujOAEzaztsKu9/RJX8eT3cpiojHBDd81R7H8yl8Qx8UzGzeAP76I
mqsPnYirqivX9pzx5gdgmM3RwJFuvXvERvhQSo/V++7Ydv+O7DyB6Q+4dMVm
ySvfiqHOUMPBGHm6BHUhLru9PD/7knfE4LQxWof6Aj9v9+vfWEOyVSDSd6E1
cvL0lAAyv13J+vbbelRyImbzmxD7B2J7REj1gOa166rHY/8/DPl+t3vcO4Ql
+Id95JpLHSp1hA7lkUQZ5vjmKhdyYofCqlTOnT2Cu4Vvecj8y0muVLlz/Asw
utG+b7oQsh10EuS2hm72PuW8J9I1AHe2pG3XUbYWOeDJuFrz042wzIYoUUuW
VWyivt6sHaPQuPygqDT3UxzsUM4ZMi0Hf8UgfKsZSRc/rC8pH3Q4ABovbpuE
dYAMvNMO7GQaZcV5qWejp7r8CTA6O7RYosKtaUNJhQ0JfDrcNx28QlpNLu70
/ASBj8D8qn4GjxJSNR/T0HXqkwGfQvHNg+dDAp+T/UW6ozSNjpbXi/tbxDEr
W8Kh+Y30leYXAz4NMMllDLBuzhBgme+fVwCY8ksAv8t5OZU5gPYwH+KBWNmd
7hLssyGO+f4VORUfJV16TSWSkRpqNjrnirTpKlSgCwLhecbxFwEJry/OYp26
mwpkbRnOaWBvDNUOf0uFKYPVp3ItYicj0W+tZ+I9J9537Di4kyLcWTfvhN2N
3es35wOrqV5jhw43YoFRtLGPdERbO9+WitGgeD7PqoCTseJUdxg7a/ZwVCgW
1gGx4givrgZmlwcV6nx/ixhBmqZWHC4ZflnElfdMpBJTmVjACk3TEibfMRxS
4767bwmIegK1zZ+vYY2xFXQ++ox9jTF4Ca2R0ue/N4sji1/shpgoJcAfvBOc
H0YFqBoF+VkwTlWs3eHgnz+BZSqG3MoUeYMrNPj2pFAqZtCAuw51mDXP7cJA
CM4M6DWHbk1f4SkX/D7X4QyNttFVRGjLoRiHxeu8lZk407IgOgtg8wsuA4W2
0Vtj0ImP+A+EKpWCMDvZf1ABxjCfKezHZD4BHPY0Thpo6Sl1euIkXb1oLbe2
8snHuuvEB2oGaiwOivgz5c4bHOiurl5SSej2agGJRjEBFCCNAVb0lF9yFb47
uHXapKBc4gDDNs+fvjiivcYuimp207FIhU431qEA+Dy/isLUmmUpVQR6JYgA
jvSP9AijtgbAuPkt9iWbtSfiCgtxIGgfT8TwQ4Ss/nGO0ZMpBI2b1gKw5sFb
tIEu0LXw3q6DDPlNhNT/JZDUb4ip8UwKvuu7nhcMakqlBqZbkoDexfd9OTXr
BIWOCJs2bB2NCOIFVfNj7ASu4DX4j9tlj79RMvIqcBecLTzZ/MBE40deHp9T
PvX/bXrDGiQa8Ia7vashR4zTQGIffP6buDab3vHV49n/q+KUdladk7H/hUl0
0FoW02fsbDOJ4ALpbA8WT3tuqD26dBIAmjQdpt4Eejfo7m0t2mix2WKxtgcU
BNItYiVhkyVXe6tuy6DVHw5Pu9HxkXjnebQDG/uEP0WqD/2RrK3Lkeq3qFsc
Ng2YanuCRoyHiXroK65fmvKRNVTUBOZ1oJEkxVl5hePdIPXReidigAtP0ezf
eQRUzg68lU6qf5F4RJ/Kvej1d/4V3XgXDOesHv++TbWYQnLYokXDiuiNBZhe
V3RpflO4kf1iAiEhMJvTNSRBCsSuv6eXIQyecM7EA4XLOjlZEI3U28jq2SMH
P/nutsFjNIptLWuOGyxaKkYlyhuOZMglilGMhE93YP2ec2yg5g1vnC0xKFQF
iFTSxr1SYUbRlZ/iHfUTxaTUfa8iPspoNPMcC0fNp17MyNuq1NOXfeOF7tlJ
t/oitPv8glDMVw7ZFuNbooexWl6eMH4bHMed4GbUHkkIHnkWIiAPc4xLaE/e
9sWudsNd0jE8C0Uvcu6q5O0uRs3oSAi3zna5mPtAM0NzOHz0J2deIpxXpN6Y
mjqy7ZehiK3Oamp8M3GI7dsG2a4kbHpO35OE6RRVOksj4+/aH+TGOgyg8vGA
Q3EImeCJ5++1V1rfrpwElLIyU4Qa8wvOGRKKfVeQ9nSX6bJASbdUuirWJFx5
gODZe9Z7dzHRKFDfB2dW1xJ7PxhdaAXcmlnmvXzxXJ2HGfz7dMlKYnzo3x3y
NySCWvqBC0EYVp7FvtW86di/nyBfC1Ap3lKbSThThanA1IENTvpB2yso3CZl
i9ma3jxC2tyDQTnNqY7fANFxb/2ZMCvar8PBNhskeT3KJ3sE7rSQmhtz7dfE
xJq74UZNrXlLmm5C6a5OCx9HEMjNaby2SUIIr7iBtcUYfg/LPY5Ck1s1KY5i
VANYX2E7huO1st5CxJj+KJFA1Tnzl+77Zd+fM2j5jAsh81O+S5ohHU9akgOS
85dQqksklaYin8+nrHDga+v3z0BYWspOm4t1XTvwTeYWeB82IsyddnTt+LUd
OwndG4A2qT16NBB3Dl9ZDfNzbvzWxFIEbb7hdrTn/2vNkujkk2TQzD1hUW1o
VRV+r2MUFVSQBz+TPFujPZrcDASY0/WWH/qu8Rc46Sp03gE9rSyK+bSDxlZF
OAx95rEaGhSi9v+YdseOAikZiWs3R9M+sHveXKJr6Ifny5+Y5rTAQaa9HUHn
Z7HBr6WegklaTPREoCydzO8Fh4v0bn+EIfLoA04Wo5oGMMWTDk9OrHCWdd7R
eMrat6tMucpeY67E1wVBUQ5SX+kqeZparFzDfhVuVqTNp1sjslqin5HdsIJo
o/eh5nPG/oygtgqTLEEfWeWuyHUapOrbOnx8bugDmU7AA8Ty/1bXGzqQDmr3
BEXyukOvq2cdMfqI3IHsVIqBtRk64ItIva0Sa6jqe3n7qFu2RnH2ZWnFDO4l
cXgbCODHrRTCupy7f0srM1cyDCqkI8Zfw6oKINVJ7cG9L+Mmizp7VT4qYtQN
HEVuft6Nh3A1MoIZZbJ0Shlsf+DUj6ButT+RU1N3GRqLTpRlyWH69S34s9AD
KaidTb7CblqQDzKlYWLPkblsO3d3mIASLhWmDxx+ydjFTbxdUhOSCppcG+SG
OY6Whzm09Ri/u4EG/hNnqazI2R3dSv0rJmR2kI2F4TP4NYY9PRsa88XIvB4e
1sKVFSFXA+rptYme5N37ysSc7BsPPdo8TKMAeGh/wntZlGg9w9zlrym5moPo
sLHigeph/PkFfyJ3cVdruL1lt65avJifO/7NfHLgiLLVHAASONL+Sjb6iGv8
UXf2P8a8Uy5x0O8X+pUrh2yXLjey31ccK5JAl8WG+6RyMHEry8l+btf70Wry
v0pIaNkJkeNkZjSXZj3lfuLxECkCysV2ph8ZW9wUHt4Kx8/vOc+B68ZXtpWH
gXe/n4RLTx5XxlZN0uxA9RsdsgsqznBksvPk423ptcqPEqhxBOLSIor1TZjU
x33WWJYoZGFoRwDjttfpXrnH1QCSurvHjch3vLiUS+M0y4cohbA0wwa2MkoC
QtpU2hg+f1XRKU5NWt0VdVgBMh6NOUvBxASrULkt9hkF8g2GaglRnwuwy4QE
+Kjzwu3NxSkvIau1/b+W2bjd3PAcc/J9hCeCRnVbtwuNdrY8mfNhh3ye9pfE
IoHSaSvle6b6GoD+TiOB/4ZoExF+swimf+YuEEdUdYy6SEhl8mESHpFFsVyR
AM38O5IhpSPlmuWXszbpqs+FDA6HDzH5lrEoG4dtKmHvuolIeq2yk77iTa1u
cKwnHTtYqc/bw9PQl1I59pH0YtEDd9pyJ0VZBWkqoxXn+Mx97AdaEKNG+pKk
Zk2vel6dcCjw0QTuvLBiv7APQWKS4cWPrtaYXm6Rus14LIf4jnP+Tv7AFlmN
S01Wu2YqRzqvI8mSeISIfh5LZnak/IoAUY2Lx/ht8PU9SvSpu1WW48DANhJr
13qDiQZPrcU4hh+Y1AqvuWyj9bymqj/k3nhe4JuN07sLALACdInrISd4+evI
+WJ0G528wKwioZXH5Gn6WBqN6zlfulmUof7vJ71dSumSBH1kve6UEuJ6vZY4
VVVwd7cgUFBFt1H90xDulbkxD2UC5saMYoYrPR6X8Eocup1saV/T5ImljyoH
RGRUpJutI7Zc3w42PpyVnDAIFNNGdCTLNURanF7zx6DtKtEL9ATCPj4w2fp7
iQNaUG0ozfEpmVt9exgIOC8KkMp5lg18g94r3KdOWrMjOM4FNsNZC5k1+cGS
+pHf6ZxVkC1VhGwrv5LwPCkejXO4eyiM7ruffet19L76tlKdsEcxIIDoRtar
ZH/SKyg3Gbu8X8vEg4CDon64XS7jCWbP5HaSx9io21OpwZF3gXu5y4Iytjyj
JZhcA8w6KVJE2AzOAElJd/7Yks0pNAzXlOpnYJuLhWQ/uyEOdKDnTWBPpli8
9T7baRpDJmPSBmZ9bP8zG4q6JOIh+l15GHgYcy6rkoHqnMbiQ9m3J3FZussT
ipITL4PZvHq33rm84XL46yho4CzH3cIfiz6A9h72KSL9d1Si8g3s2Cof9Z5a
DxLxSfPrgsXWUt5lUS5pfhY68MzXTZCv7yhM5vrCNQW9DgD0PHoY48PdiwWm
s/rxZF/LKTi+fV8u1nHjOLzLGmqQhG/EXthgrXKUJ5CyeFgOI3WzyRBLHLEy
EUuqKptqtwCHWVHXFWO6hpawBUZP6uCEJ6jxbXRrhaDlD8qbC3sxNx5EJvhl
/4dXV8v6rc2WJTFE/8gewjhYaNjjP2eN8wzOd/JsGmMXKu5gczhxohFQy3oC
Plth9sSKqcw1+fLsVPmCipcQ4IuS5oLL9S/W7pwqiO1GoFOL98EUGypie8OP
ZWdwf4W6Wg0TDZcP0iJiVKln2vknCgaxdsjCB1Mi8imkeGs9MhYqiauuI/c9
sZjYeJn5iS0gyny7l6ebOAxwnlkQX/Sd+5sOpJ/5HF0WdFGGK+y0j5K034lP
Y9JPq1+u1vgvv37J9IKudZG5axWGNXd0nAlp1gQXPOnUxlgv9C9vwdpRdSGJ
kRDOP3AsH3UgViai/xuY0lN20b792eeu4ppGHxJPYEXHHq0uLoeRIs7/tUwV
vievLL/kZfYxoEuUV+xbiXOabfeWpv2OO8xPqGjqf0nt6IdtTDf7QghEOwbX
mdS+0YEW/5WH0+PERTcHac4b4zXy2StlSXnMDzmmxMlqGWk1qQuYc7kyHCe3
ZLZB3ycHSVdcu9gXXNyWckhaI0HPzX2RyC3A7JkLjwNCJbZfdgWs+E5KHcgm
LU/MOklqpUK2/L/vKsDbu+rybGXbDfVWtfnbnDne5G43JcnzRQvUUpfgEls/
Ix9m/ZtiqQYMjD97f3RaJhxMBnEGmi25EZ71hSU+fD6djznTAWLdYAfGvFGS
uVRyGfN64WFhiILUBVGy20NOZ/QV10XA19hJLbs0bQSLTwgXwzV0mGYJUflW
ULXiVPekP6G1uKpoy6OdN01+OxgrvBi8f3Q0DXkXpGFifvNVPPKUMBdoxjjM
uPukHtnspwMndS/fw7+LQ/1wGBZcfqzrz1S51Q9C5FXCO1ae0Rnp2hx34D2l
YoN4v1TtK2CngN5yRH4me8R/1D1338CUvvowJRP1X59JAOmlx5ia5mCE+s6k
VusZEw7DW4sbzCCr33dLTM3TwpypMgeO1EWf1lKoapWrlcFVa5yMcbMXhtTe
yPTwkfkZGnH5VHDJ3kpAw8GGgydLNv1PHUKxZ/NQqKIsnQnkENuBX8OSQdf2
9mYrDCqjNMj5xMYyi5dV+tFOx7yPHYl7uEuafZtncCjd/pF3R+uCYCpbscdx
5QhW4d//wxce1vfXzkLFjgZ3A0P8xyiJW6C20vOa0KqE/BOckRfDjVxtvvKG
/FZ9tmBMKW0KFQyMMaLdJvPXUsmhvlNuVo1n+Zunypf0aHgvhWroRphsL+pG
Cw25Iw47H3V1ORQzDXEj/UyhuMQShSJMvwPtZ3kt+lxQsjerczUSBBdIyVbl
4sdHDX8Eni5ktTSo97jMhF48QChaPHfJ+9ZxIxJwPKsgwMXaIzBOruoIaS7u
cHHHMr8NaJoEIYUZwXXzdG2GdmfBn94UAoA5BQSCVKxfGUD47JP7DL+ZQyRj
OqSDRjIXJL2aTlJVp3pDIAMgUcIM4fDGI280J833HAUqWn6nr/FqGLg2fJJf
nCi4ep8w6NJuXiS0qaMEgBF8Pdf0VxwBai6moTNo6u5OqTnr93Gxrg1Kd5IE
84uubLwvWtzlXmnLSjtLpyYUl/CIfj8+tsmxXNTrZmuoOyNuOWoL4jeANigA
h+YzJTWynfbr0B54IUBHNhn+H4/+JmzbEoSnhfsNE68b+zTm+O691MgSX6M1
6WRgvaIJmznXQH8eB8QbEoV2s0gwoPE8y+TxwcG+tz5fle+V1DpaMVlVW0fs
Hjovp80Be0pKW4sC5Q8eiQKkDpPod/kuOjqTQN116WrhjrnLvXOcJ7ishxty
yJmGlY5r1kxwzbfJXG/vCdthDIU1iAoCOkk6hUTSZGev1eG6jgdtdzbucr0F
RT5JqaiTm25NHPVmDP+gDEhgopoIa5l+kuPiKJitmAk/wbbs0507NBDo6Zld
iAacU2JDq/KtzV0I3KjSsWdxCkpBzcmJjuzxv+jMOif89rkjx77Q6wyXaK4I
1YbJTzTXd5iWQkxAy0TdWjz+XnZVjGnSYfE+QXuhyc/ZBIQrfUgHF2ihuqjc
KqU0a0Gf2ZcN4HKZwtuDOEq6ZGXNnDKiXfRjuaHmvZ9nMPZ6lmQuyPdl4jqF
kmbtZA4toDU0J0QrUa1nktYkcZtomhueE/8JwUnFkMQRHJ9qwetwrsTmTjLS
7xEtmkh4Ro00GSm3igmvedZ/7Wef1h7y1elzkuDEUZNAYtK21iKmUK4oOoxu
vrzw9EJNig/g+hJLaBnCv1fdoidq4UFQsrYJslmcwBG3VmjY/UsM8I5HQy4G
5X2LjEhSCULEm7IVnly7wLGZlIb8KDz1Ac4VVC83oT3Ba/4F/AKwHwdXTt2f
stIDR0RaDUgEp5aj/psMrf4SREWqtEYMdUZMlTSiEvb+whtTEOJRH2L7Il1q
FpmV6650GqZT9zuFyXwKdog1QPs+23YvM9XOb44Sgj7BTlk1vn8akrNf+Jsp
WW0wKOQNMn+y5kg3AgojVjGXwMv92Eymn9boks+5kaaBaEa/njuTvpo6zDcf
vAYcfufXsUx8mjlrwx2W6J/qCqCv85mBMDzgPmFvu8g3vGFJOM/N9Y0dXPTH
/N41lf2ZDK2JuV3+SH9n+/EI17ENzkaM2cx9AoX6QTrx2whoMkFfwlNBqTuC
911oPl9IqBWGKrlYlxexugws02G476T9UkagW6eV4f5HInyCxpkpRTj9sMbg
2BPOn1yLhyk/QS1EMT9otro8jT4InxWvsT/2rfxn2mPl+/V+d9rvcOZq2aez
I9AyxJ/7OIOHrFgr6WYVwSFzaVYi0Ku8Q3kMKe6jISSIYj+nf9eJlFsAq0DT
KqkmAyCuof7is9sdg9sb7g2PW9BGOaEAaxZGHSFYM6qAWaTt6NRBJ1hPqQyw
SHUd3s41LD9Sv6mUobMikj5Yx09nQQNojUMPdb16MrmR2cMo/T8CflJ8SI7L
WVddleolt1/3RJNwFgU4PcGg9C7W1xt3Lp0Co2WEt0ctnQo8c8g94r8qxDc+
JTuNiiwtXiFQRdVbh/sK8WhVLYYPXPOGeRhovzUiLf63iqW5YQBkdO0feKNf
c8laCPznHIz/a/5RIVyH26EDjnYE6hqrB6xzcd4C8AzEvMp6UgUO3ZJnHrE0
HzQ2WyX8L8V9+Vm97+88hCu9KjWDupkB8NsY/fkRx6nlc9/d2AY9AhTxgXFL
xPybLPNPKRp2QfpLw8SIQuXkghfdf4g8JSYNWWA+0EW3Atv1vt3uuZxZeUM1
72WcXfhiKwpTCHnBjMdm2gT/TG135A2/Nd6cgH5tUeaeef8NrUJdL6+EMecD
WyG5DnOmVodhd9KWi7LhgYubIvsaLqm2+A82yTW+VJ20TH14rgThGoj344xc
KadBAKiEVBlYY7mWWYA9cM5iQQAjICKhHpueMPP5HXHmRc2jnEkA+wklUtIG
JV98S2Soh+66hzG7JnrK3Gfpq5TurypLgPM0MuIe61L4+0AuC0/bTGFB5AM9
aZvyOgy51c6zrmmVvReFaJqpJDZxMvtAYBfgWgppPZtlSEuhi5bXEq+cnrOy
d+UyfUUkygl4ULWEh0LlnjZEn6p4zoIYskxwD45IXwEQHGAJwDccfiUfhFh3
+LA2mYP4h0ipG2ib62urbg1QxyK4F5a3MYswImEbVSyU+J8+HXdZxzuYZqJq
o26pp+cs8RnyxC8Dwixemb1sgmqKkTdkBy3jvYgsE4rZdxslAGQwX0q1l+j6
4llJ5kMsIi4WXG42lhKUyaE5tQIYpavBayk+38E3Z9e2WBrWHaHRzCCGjT3a
vWWnHYXBFWdvpnh3CIMUxHnTx6Cwr4Vvzn4F5GkisrV7Ufn3kfDhUkCP7NNo
GnK89GoxXKM/nY2AS2qT+Hj28RAHQw3xnS/11ndFnMljHe5z8x0GVl8T006Z
0txYxjfcH1jMCh/JASx1IDN3aBj1xj0rWLIeP6HfaMfomVHp/rlWqEh9DgBH
vnGZLeR5sbnsPRZBeHF1UWEEweIf/b/oKaqSt9qwu6B63EQ0+5osamPNbTlo
3jBNooarFhuM27wlRXAfK74JjgdnvcOQh9wJIyRVnnh7WtCL+EJmeMC7G13E
VJpzwkkYYy47LOYiB2zS9uRPOZNrJql7Aw+edGgqk0d9Xxs/A9VJVmDBPeKB
1zu7Zfql/6PEsWw2JX/QrBZIyyNqSdMpQg32D4FMInNVKRdVBx4KJvZUMc8h
fucuN88j5qWQ93kOzZqs6A97F9NB8SzwrlASOqxTVGU4J5rWFSlpLCF9jjkQ
/yrKnk3++1k6mh+B99meM6aqYSWy1xuT0FwPkTZgK8HS42wa+zbPpFv/+urS
gsZD4dmWOMMXiKq9MC5CQcwGpWUbg4rY6dHqKCddqyDnHoeS8OXL52ODAKB9
tBV6jhK7d8UwHfwHbqUKYWeiw56+atY3nplEMP75+vdWp2ys9jBF/b4Z+gii
fgITVYb57vyeBvPWk36sCJMmuhOkPPCnieshfL25SjOu7qrqt/myph1qJgm2
qar1yrx+yWk21kOSdgW1Z1mWeHhJEsijB8zda995+6KxaML6SO2cDPXwCc7u
njEL0yR60RkbdV2xgvOyzGkp1ty4atqpfDGQL7fL3BjZd5yQmf05ZuJ7Vruy
pT6W7prHW4FjeD3aMjygxHswG3iIcHW3H/mWpp1ip1Py2vQRSkLpBF3IYDqQ
N6xlOfIPPd5Ew2wgwADT7phho3DnSNdkzkAGANDVjplVC7Kmr3XqJsY7cjpU
x/lBblKWD4Ag2ZZ/VQFicjIJ5CDkTKpiPLuGipjbM7H3mnV3H3MXAUbUxu3O
aui1jUnfJyRZnHIEtINantZDFXam62erFSLaP6ssb89Oq4ftU4N+pt0GACHl
PJ1SsAJb0FhMYFS+cXJ/YE9KgilNQ84pwT4/sntguZDK471os+oo4LmYXRPP
L9ULwMAu6xOoFSwuTeGcNOi+xG5hSV7MG3HOcVomQbcPBW4p9z6PuCr9qFre
k/KOXKMoxxn+EMBQ6rbXhSCyJST/QIM7TI2zWTjts4KuED2BKaVxFqkSHB88
XH2C2y9ErZLyU42FU4LKQPqGvSdNOd/8thKFZhib1hgPh3nSlPNqf5pdTfqs
68TZlkg21FnP1Qznha1CxWnOsjb42tM9P8wBaLG4WOjn7mwE1EZ7SgMLvst+
suhA/S6SdJ0TQEcfOYgpuQ9kvMHDUBYFq61Hb0AWI4c1v9Rt8c6cFMnH92NX
1QLtQ6oVUOEywV7B405hTCRb89+ig2Ij+g9sfJJezSr0ISRLMfCvByEL2CKN
CyWBTOwmgmmPd7q9mrVzhodyvXvAUA8LHbbrcoKF0lQLc+3P23sRvUMOQb9A
dRhiU8FzgI9RZ6TccurTNXWuhS0qQit6MevvxSzQAw/TZePtlIk1hDiqCJBO
qxUwpaR5YgTsee4kqkAlJq4fyuPsTI1rcHFV5wxQOiuLlwrjHy4wgWKRgoAj
nIUJp6n8fYX5iIRYmPjckJtrASbzDx6SSqetNdsoUu1LMVK8JIqjRwfFMDon
I6G1mPvYYkfXLY2iIaN9AEDrUCIimfQC4uRXAYanq47vOKFhs8kCCBMCM03A
zOPXMwG1Ivi3rwk5jsRhOmLBmx+MMUkUC0nhoyEiyENtnScvKdMz4uIiY2b9
dupWO0pKnb6ihtKl2SqmLt0OV9xR/J0H156W1320dWDyo3qTwE/8mfpWTO4Z
fqkNjs+UrxqnZuD0iZ+aoqWZdiPQ3qDVySBdIBGDJal6mWhXw+wCICVeWbT/
6nKa+OvSOIi32UaLKlh+oSbwJtlmRjesAPrn058UyqrygX3YaEx3KJtwWw+q
07e3YYsheSG8r1MxQwagg+e7f+iczB/Gw/Zk2jF65baR11mk9bo8UTpaLCbF
O/RnuLfo9BZ2vJlxTc6c0N+jqQ8c0P7H5gzfQajC9G4Of71G1aXgY/xdehrN
yctsWA1hreQUQ5hkRGt5X1k/0BTqkasz3z5ENl1JFaghg7Wfz9xNFIeESVMP
fXEYz0Cf3Ibi8UepJ9s6xw07EyMb5RYmutZBYV3pOxeGzrnooudMp1fA619a
aH7d0+63XESacVnOCRPlEvMcICTtPI6Pan2RbXwtlzfx8JQI76TdKEh5NQdh
JfBpkYA392NNiz4PEQR5hEEcmbIRL3yqZVsv3qAt4d27jBGTdbJMTqu4jby1
aPQkp04NZ4wZXZoF1xdRUs/K/Nd2YK1u3mWO24Ib5WdByHy6Z5eB3xTqdf3E
tNFGerY5a7clCS2J83r6Yr7jI8ML43KcUcxdY7smE6cqlaNI0JsfHpV7m59p
1cBgxvjA9Em4SdxuMXA00k/uk0+MuvL7rAeAddlEXbhR66EfDVkQYC/4kQFa
AEIHUC5dN7ofsupvYNox0cjm0fzCnOIxq967w57D4WCbuRbGfI4rh4sIafSZ
Gu5U9DVXkQk8m3r1xuV0mMDqtQsK+mLW5G7lUCvQoKWigXAebksr+ZVhCrzU
UN8CexcNNa2VIl4uvx7OujrsAFtn5MJU6ejTgSbvY5IwikwGsx0DMbnzG/QH
DnuxFnjfxJq3AU6J2TVIRZlOt2Dt9pDFlcpuMgwYygu+I5slIvgldw9I8vC5
SrJhqdSIYysrZrwAJna117hbNCDky/AtRd0EzWxsvzTOeWvsqkaWcAGZ9uwK
1DmD53qg5MU/g1AfFZ02pbZwmQDH5OukJzLNbiAr0uIuswowr3PT6J51M/6r
zdmw4/gF8+JfvGVN0nT3WhEjj2wLIJG+T/lxotdTRBn6KobuLrDbNYS//gtY
ReXS7KdPNcpdEV9nf5PUzeSCjicEvMWhovqc47KakisO/cKdQx1w4ccBuGFT
mwB8QTmJaEy1oA5qqdT/obgZYk4jF6SGgNpy9AUy+TigQH/+SMQGyJd4geIw
PB+Lz2zyyYKm2IaG/PjdCQ7s85FweGjfrwP+l9gVyV+2sjLsaqINUQxszEC5
KDYJfhONTSMOcMUblpLGplDq4560n9qT1q6ofBIjK3+b3W+ypOzYidhkL9+s
rXAsnLHKr5KU58y80GMKHN+J41jstlDMl9RyXtKXrHlFe7d4gPRz7yFZMJFx
z9WBYkoJIqDu+3WD7vpscolOlQL0jMFV3REXLM7jWkwmPx7dYrzQWLCNAJVh
3fGxRpXFt1WcDtd0qpMOpyEMeSFNvIwSuErsaIdpMgIPDTdztqAvOhZa46CY
wqIk9hQG6UQyrDKTcJKmRhy2VO2/CIzZMr4P3/ymRky310PjirqSlWjm3joU
z/4dn3Q8Macq9ZXSvhRwdmzgauKwDHlYimgInyyR3vgyaBlZNoaNeZN6W4Iz
dAnV1YAcNmrd7UZOfcj8CJtyrzt4eALGJ4yTD8gCNNGx8v5S4ukJ11obPZHK
S7D/N9wRj5VcDCo8PXBtil7njJFvatSjbHJc8D7C1wsLrTwoJYBIQUEHidoC
+iHMNoRm6pSauCAHR0Np6tGeofni1CJMKGbAlCzmTs5L6Ozx/s/ull4jkTzZ
Y+/MRPa/fh1lsbDFalbtu17gnHFw1WStyqroVlUX0yC7NGEW3OTWYSI6dlmi
19u8rJwUzPIUOVVx4OBXkb/JpEeVm1UAGlLKAFfGbZlg1+QQiBYpoxwvUEHo
nJe74DgW1gp1CcsXWnKl+DntSXA/jWoBi23Gm4tgATRN858BoWvvTdAAZZQX
cHL1pmYxYtogMfHtDQBd/57hVDLdyX0Go+xUr8gLEnjDxOzamHmKZ43piszS
2trxiVzU3VFPYFyDjblaS7iGDY7x93bsMECIVGjb7UwjP2GfAZcEgzxlOEor
gmFzFBUqxCL+tsKEdTXLCVz0WxMwmkUtsL14mZH9tyXbfW8dvSArKpKfEVua
I5DiTPIEa6jteEftmF1FB/AFf4sUNBZnIebY26bEy2srZQ8z+6XlzI32aVIg
jAUt9NPH33++aK+H7hXW8DTNi69jxbDPvus9flAio/sFHbmIcPxwu8RaSjiz
3MnG/4Rq6tAL+1Pc2GNi1ix4P7s8D6HnB1I1doTVmxsvO8H9eknJXTeCYIV8
bT07fVlwcZLaV8FugB0mpCFcm3V1n6Ei6ksriVMz4bkd3ClrDzuguoidFZ7/
lr//RnfD0X/NPnvsOxqkM40vmX3sLI5AxSuKfNNhSvXgzRtTczj6KMw0Hz3y
oJ2yKxJLkHdy3eYAXJV9vjCtBHIw2i3KRaoSO678uys5eZORQMJtqhPZDFLd
25mEDq2qrFCH+O99kHlU/GyP56dfdDJJxpiIa53FbfBW1AOgp6Gb03gUY3Zz
b9rRHpJ3F2G8X2Kt5As76reNoEO6vUdLH8dMKnV01Sw1iDEFCJeX348viu75
lSBD6Ghqx5n0719mgNcfbJCBnovQMpRi0+1yxl6NBZwJQ5s1n6aSfqMfx1cO
0x3iiqZvuRY3hk9gvia7RvhcXiHotnVFtJnQtzVBuN3d6L6/PKiNycpzUBnS
5pZOCiPc4vh9RD2sMUALqRY1GX/Ewxrc3r/0RgqDCPm7/G5V3EjP4hA5JQGx
XIvBbrzvgfBow5XBCXubqHuzgF51Mpi6iap9kTWNz2YqGg5qoqfGJYVHdadL
yWx1h3DK4usuhWTjG6Fnumpfu7IfCt/Z6SfS24pJ3wYIIQ6AYt1qvMQ6x+gg
nouRZFRYEjX9/uCVVBW0VXl9pEn6ja1dyI9acx8Z/0oCvJxqdv0a9p4d4ekm
gt3+RKpWFclSQwE54MKR13ifRbAH81Wi5dDRmF0XqR1jCSnv7gUW2Tu2YXgX
kJfSmt5r07VXPwwZtpTLxHp2uTwurph7OyL7vEe5STeGx62h3eatWBgiZlhh
K1T99gl2QSdaJkJrlpGMH9tB7f8zh1wcZCnd5QRvzi54sm93C6PIhNe57yzv
L4vOBtTIQM/fMa+dA/fZR755PKGdNgwT8jKN7JI1ZBlocMTSKx3tbsOv74Xt
7xMdVYagaCjU5NFmp9EwwFMOVsY4A1t2noozWHojil0O68V0IUMObsSGLZ6F
nfuJpAQLon1MrITVZ/CWhpRi+Y6wMAWiTH1sDf2T4NAOk2hvs9I3LyWspcIh
EHKFnPlfa5IKQZ2bDIb9kJ0xlrlpMlGv3Ooxm0V4KJiSRLK5IUCU9ZCLLlU6
KaBsuVpUIe/gCCdggC8uUDo4E0tFyQDtIRQh8cpfQ0dsVWPBUeU9Q175TOOv
HbGvq3UjxvrBrIY1mORF4BFEKkdvuQxS/zUoASZ1eSs1M1zhC5mH8Ovdd+JO
hFf4pTum7EH5qvm6hUyaDUzythcU/QtMHoLatFjqyK9SBQ9LTDLLt42GmY/c
EwOaJvPHr8nThp2oSaw/jhP3U9YyKnxjChy5gOq5VVfMhWEqMLt6kwzMSoYB
dzJ+Xu58lFUrK0EF9cYULcQ4wfCbGdfv1RYxeyYQfHUYHh+coYwcVhGfTkNw
CuhDRZve33ym5PaGB6s1to9qLNA73GgGkU6eWbLhCG4LVu2huzw0c/P7xbqA
lybmSdJ0RiquFr+2Pj8GH91RRHZ3/quliH1/erzR2rbZW2VNH1oMsyNvvDEv
xDRZLKFfN5lG0+YLtGTBWf37kbWAPg4YdF4lms66+mYIVwdSkgULG6RkXJB9
KlTqWVev+J/ulE9cuofxvyys8ipvEpu/Ay0SQJjWVoeJFmBMnr8JIN8MsxNt
GIxuYjbT/MGlcBwDikuKNofvuZ5+7HbfVV2805UC0NK+F1aL158WaPzrYrh5
mUrWe2avYhSVaK4SqPjPB4NOfazHzNYO6+PUkI+veBnxFWTpDXYAJ4WI5Fnc
pvsnqADziai/1qEO/3COwU/RLWFUUee/oBjy64oqkhS9wfaJnj5hl7kLIxWG
zliEFyEQJMq7fTdctSeiuMREih1o6imwYV2cQn//lCGYZKrlII/h6e/803a4
EIGtIJTJ4BFjgudF2ysFec+X+hOAcVsbXnxYlE7nHqgMyjdvWQBe3iurGiMr
LRjhpywHt6nV9YrtcrxYS6/vB2IsttimyDeUp0TDeYtd3+vMdX075qyzp+gb
8SZ7KLA9H8iUEZ60oVREYysCQFg3pFVQqQV0ZVvC4pqZ1npeJslFj1ZX5LDx
+btIMzIUjZFoG4lS5qSPyx22ftLirGDbAJzzsJmVYGcERpk90p0k60oTTrIG
CuRdqcf77MJ9Rm8SfCE3QQbOV/rDOiFYGaAsh9LFPoDUkXEq6fKGj8Xy5qes
ReLd2JPR66sRs6BkOn0DfE6Lv0lDiqc1aC5EEgMg2JJglzPFVRvOifxdv4J4
1woJiU5dzdlfqhv3fQ3hmeNpPsnnvHKr1xsMVx4DWMCaIMNJNqW7IWd09sES
ibanftrnN6qTf0Ub+eJ7tYSpJxShNF6oCN1vtgW56FaAw+yhEi8lhiN1j00C
M7K3CBTIh2wbVfKVJpwonkestBPkKc426c8mXjZTPbYvLD//UXf0P6E2goh8
7KL1TvMZHxy87ZZP9By6MuD3eXKHoPX0ShqmFwsbXZ2JonfZYNtHWolkisHX
JDoxaqs4cNy9SMvG6HFfKfOn2bemb1TpG6ALngI7dIlbMFUQNA+QVmqnnfuz
6831gykk9eOIp2OlZ+XPUju0cHY0l/l9qHmNZ51GRbrtW2O7CfNxeNzaUdb6
VSSaNHfTHKlsnJG9vaFMif8dxkY7m16Qf6YmPHs2X6TzgBk7RQvGy4WleWMU
PqtOphhET0gdI9GlW2/k5QLXBAl8BnYS9B+IRma/eYFuOqN57uC4/nByW/NW
YHAZo9q83YSnAOl0i9kWBdlryuR9/4st+VWquBwjp59Kcdk5oWYQI4twezby
RVQKQ7Pz5DfeeH/dEoUXsi4vVi++LjsrSnM34kptovaom62LKznjRdOt/SO9
W2TKt4nilGPTjV1o126KGK6qjHEN4H9tG66bS0B8824PzBQmbkQw9luMzoEf
cN/nDzVta8noZyf0wlBBtzEE6JAhDISPfB0cthqhEq8z+BLXA5q9rs3hiR2I
6WUo8NcIk8qcmf5CG+zcAZ0mCJWoyCiOV0IfyvR0OGe1PUDxi2v5rdFydHbE
nTO6M7Iv+mrbMJ9JTz/L9LVpgBOYCsANEgrsbKgNCocY7Rxlz9aVjvsJ3Obq
fkl0PahtJw7PFhVfNxj2b8P49VF3hB/zyYF7vfpufuieX0+YiuoTcP96kR0H
/lTe73UyP0xBiZ3whR91dz4I9+vSjJnzfAnCQVY+iDubIroO2cM8ryK2Nd1j
ZX6Z5ekOP+z24a0Xz2BoSKgAOxGJKVYsW0DnSEgaFeijWp1q/C2u4Ohz5GVV
b0Ks6NNAijhgMF/sIAepQk0hTBmDZk9jQuMGIeT+pNKLoKIsZvpmrw2Wv/mV
vMsEcOL/skcODpMIDqG6nIxOiv3Jn7XXFirpmC5kG3CHzOZzP9MermVt9onM
OJZqG1E58eJARukvD3LEMZ81ZepMTmWsMx4VD+5L6HOyErnCxxyVmuAyWFgo
F0NYRTZ30uNNf0VXYvd7leJkAw/6qxIgUx0Th9oWZjsTNgFgwBkuxJlSal1+
1udJlVLD1OpX4m/hW6cvXUZFrj7niIcQrkxRsxiUM6pS/+Gys3YVBbwPuZ89
/teQ1ASs1TZG6DGuZZ1fjCRskYFNyBqA/YNhAwgAFSeThzOCfaYuqMpyyo+G
/hQi9YK1uxtlxX2+B7LKwFz2yowgft6q0g2OLLpQS4SbK1W6ZY5BeHhQ4y8S
GSPY0sD6G8Nv3VYQtgzVw8dqJea33/Q0uChLJ9m/afMzXfvQ1gYAoq3A06KP
cQJcd6/F8V+sNzc0q561xqHYrOKpUM1mwFag9SoYL7HbWj+egbOqAM5YM0b8
zgD3KZpZ7QmgilV4yZn/pkuxURPOJ9ChGrMIRlefBedKyFlmNv9E37O8M4qX
v8bk2L9McbmTX+pZFMwna+oVBiN3Hivqnh+3fKV7FKedWAD1lueDEKhLJWKx
/j3TyU1xZcxMgBfAN+vdn7DXCIDgEVM9YbYEN8o6HyTo01O5dCnQiVDxBfY8
fa9ppYusBZm79O7glHqlVh1wIX+bhmHUfwKwq2kU5DUP6f651qAB/VXDd7va
Ww3vz/fOzIg508sTOb0/LyKjBQ8HelO7ubeFNlgsTEpd1+XnHcb+hVD/GtKl
xbuYPzlDSZUK+3RkqjSZstmcSqwo3zROZzTo9PvP1zW80EpaM10ho3X8pnY/
OhQHY1rc66sHWLXGopQhE29R6vF/DIA1l8oCE3YCl3YcSvQIk3bSz5pdnEq4
Qvf+u18GoARCLIgknT8jhUWWY5bp8j1GdDAJKXKabStuSRd53DBbhZZ2v6+C
IaVxutBT00rC31g0WxqSFhXnBQ/7+mFQpqIzDdhaETV82P8DSPHBZGoJwqWn
RQZLfBwZ4+PlIIpuIK/NMBlNzbK0ePEdEA4RjTaSIdPQID+ZtVPk+V2NRYQz
NW741OInA5bXTNLA5szN6U3GhxCWHB+faNk/18vof9MEwagZSdYFLytshaXm
K0BbuzpwIRR98b2Z3Heu3/ljHVt7jndNlOO21lf1pKO/ouME+QSyITV0TvGs
i8MeiUWlVXQSQfoTbKftmBV9CczeXkVocRvjG+N62Jf7oWsqVNBLpfRxFe8M
7nNJv72NAWFq8Ac6g2qrirnOr07xQarnYq/m08qr20OT2HtA4pxdW5XbYCuP
Stc5NcgYJQkzC98iepP4ah20FdYqsYBOiDr9SvWTpZmAuW0Zz2QbjZu4VWOK
GR8VZpOVprAHNLgeNNpPiI+8UD/148dzo0iFFTiWjvOL2QLECTPfw2FtQd7s
9+w2ud8+jlt7qhB5SCvOgAQqtjv5rUNG1fksDpugvqpretvoJfYHt1kkwhUZ
n+b8KH272rsgi71QeE3KvMcFrD7O4x+nAtC3+PtrkD9Wj54EOmy/c1lROABl
pAZ+yWQuvb6CxdSWpCMdAy1YUOU0ojuTowd33RxKCNCkcVn28n4ZmjxIe36T
M1FcQnjS2/nCEntExzjBvlhHAcf3KJXoQebfPRJ3WxTa7VGckHpIP+g+y7fJ
+83tulYRqRQCqofzVL534Zdf5d4Np8x5ojxVo1th3nRHqDRoxVVaHjJu5qM4
LwQORsD2Nkv60pjb8+ThO2byIJJXqkKkcTFRgrG+hj8NCiw4Vy7n9xTFM9p8
EiwX70+Tvd9y/hRcXYNuc870fLdFzmjXidhu4XX4Hk86JNUEHXx1nvzovAVN
HEomzrPVpeyU34H2XR8ZZOjkdac81dXQ7Jm+6GExjdYEN/U9vSehIdjKHzBU
iOrHM8skv20yfUeyeKvSWcg18e1MQNr2fRAHlKq1vwj4/Ia2Gp6mFon2cswU
RlYHitiFlqqEbRU6dwiwYhbxDZjtex62Z9K0j0KDRodj4KD4CVX2K/Y0oGlj
JFuP3LFplKLhlIkqNDfMKR9WW6WHMBc5RT4tGpfd8U+XhHdNdj9t7wczwwMv
6q0QFgWn+XG2BnBa8fM78oif4Ih2SJ67fDARDoRuF5k8yWYFTyuofqmEFBaa
wPT73GPBNNkH0eOnLnbKjaYzqmrSO6n2fGmkoISWmQbi2RBxoeq2+vEzMtFD
1H+2a3KybjpiJd4RpgGNh30qK7bkiN1U8jZhJiCddARo2BIyPiFH5apEJNmD
7wV4bsoFBPfm0rNTE93BTM+SV1ERNkqIiAgJvF52dGe71Seo67raHzSlYT4o
xyjemZSMQ9L6oAOiIkPTwWol7+Oa8RuiI1sZVxhr957osNOxETzuA0xg3z8S
x79oNvXQ0NrBM48T6gBF8umWr+o601NcLnHOI4Qh+Qe7xSLiac0YbEP4a+Nl
NsniesbWoO6c5/X3gb4Pzd4bimH2HxH+QoqOfBpz2qcVsZe0l+1wLzhMb689
m7NFxw/mpJfzcaBFxRNHHA/0cHDr43tFBT4QgxLo/Z6p12XCla+4/Y9JqAl6
V79ixBpWeFFS8xmCbzq7nyMvr6mb0djYqoCCec1weCN8ve9sH599Yy+efauj
++XS6AryB71tgAsz3FmqDmgJabjlhZz7zo3tK07lH21BC6aUvMl/f368uXmm
tgatNuRUV0a6IMKNOlaZQ4WROrHHZxzbmUxlIFuw5IJAznEyTjIhsb7jzB5U
RKtVXGBoTBb3YBSZ4vOz2QkhpBP3V4NDjAtYzBcscdVxvQxSojj6q5tIqS2N
c1em60NpXCIFtKX/e9yDRJvdnMaz6dhtKi9AHOULi8Vk8JSdk0wXBExjmyQg
E5AbI98McHn2FhQBU7NwdxZLjk9TlcmOKhEn2Z2XER3qo1o/papz3+yL3Sec
B7lAzlNYn/HqU8Qb1Wd3KlQGCH9G8K3dvYYU7OJdxbQHeSi76Wj76wVHpGSV
btULSjpmwchPRu1HLOv4jB8X+vZ2QCjXrC1vrgwKBO0TT/VjYdw90+QfIwrV
Dz8bmWFuMlCnUAk7B/WkMgOtVcMpcfYPZEraSGhxe7rpVg0RVvZ1sAcMPKRt
FRLYtFjCVtotZ5jnqRPJZ/6MWBctHb+qq0bMrGR21qgsUiurXqNhZtLu4f6O
5ogi5p7LBB6kPaMtA8GRPPPkO/wga9rFbYyP7Rp0AIVcBzvdYl1p5agbo6Vm
xLQ9/VHmyFrnApqCisRiiI0rqzGXQSVv15qkNmIyopjOrCHyBkUuGjeRygVn
c4OvgF2jjs6AUlDbeEqloZcg9e/reC7EuR5HNBFqFjYvzqIql6/2XqPCTl7l
NmQgr5a1qYz76twBUjUZjgug+KalvO85pLd9TiXm9WrnWBUNfoqLU7H6L6fH
FodFDBoC5SurskHmgfnHs/vFvtTI/BuuYNgdAARPkYShyaI7JzRWng4xDdi1
vMm3XTfspvxT3XNTKMHuwmNl0QN0MxbLQXAyhmomhJkrTg+IBKZ/gDkhw23X
WtyxoOStTxq8gtigS31zQgT4pVVNm9JgS/8usEmPvf9oJSLF7lYE0GDRtIEw
Fk6uoGaYNhnIoJa3eDQc+saMeTLQUDPmt1PBP12Vqq1fz+iSbLUDK+d73sXP
SkkdXPgjpCH8G/6tVUIdtGQfp70G593146Nnhh53Z2DjyjbRDL4LsUl74xyw
0vVN/eR9muoes4Q7/uuknRutY5AzTK6jQrZRIgiCerKq2WHWgbxoi2IuBdef
k/UajuV880MwrrwWE4GnclgydXV4BmYPzXIptGzqhNOKKZdnK7A+Htqb7kkz
H06PfedeR2KabmvYag8SaPCEv63wY+6lvmoC7/SBF+sBXhNAVb1sdZK80rI/
tsku2Ogp1HGCq2EvLFcxYE2WJx8uYMOwlXjPt8pTNpXY2YJ66MN//NQpu8dN
ppFEF/Wo3Qa7qbfU6/qkWms9fJHdAK3d7GG74RammQXDfnh15/6kcECTbrEi
s9DMY0xhm4Q/TjuJ/xADmzL9WTkEFtfIf0FtofjuCudg6psa0ReniGNU1zNZ
WBvN5of5PhGDjrzEq7g49VZiU+DRKFGwvWY8Lh+V06rDZAvTjRhaVrMUQze6
OwMmSVZoUt9+eu3xVuhgHFzFeCq7gO4R3vfrMnYGYlcQcOAL3BqI0mxWUyDV
K0TXYzt6eOgwZGJ5YEmdVFlxkT1NBYigboiZxyjP0A3hnhExgIjsNtuNVlJj
V5k7zJMK29+W0S4/J0IysU2uTDNpqtz39PETElDJNA7jCX9sOmAIgt1oUEaa
1NeaL+uHrnuVfCV8inv99ryZ0cPLj1fvk6AWxPDDxvybKXMJbRhIWRg9G62b
ArYc8TalGQrFmMgjmvVGOFPHpNr7C2kGkOpaZ59rFLB5w02T7kH8bsoSEdOr
iFGCq0yjq0BqvSzqjn6AdgHbQWM0neER37kPi3AIFc+ynQA+k8ZiJumxMe51
WahnpdZXRUthGkwR90YYhBh5IQhxuYhwveI3ODove5mMmrA5mpbH/ziNvjFJ
JT9IOCEs48bh/r6F2ABksS+JGva0tl7+T9/rz6SPW2EmYL3mlDReLvy+tGkS
TaBP50GM2zeVYxRvZEWhg6XsMRpg9zyLOWObp8T4ZmE6J4ZMNyh8RWQT5oJ6
dhMb1ZCrwiGZnwx8nCMqspA2X0d2MVuDOHi2YpiV+UojyI+uSIHgPsv3HGi+
V7g1od7+8/JUgfWjCq37iMuJbZU3ehamRajW3mSwhfSz8XzvZFdOs8IaNl2n
K3fsIshZYN2xcOTw9UNHwFaA8L05FZxzFQ0YmDUIFyFYN5e5rjJ1dUIFxn9k
RWkcYQ4wqjIX2QywWc5QEXUoc6+f6Jy1/9pfC071mV8ggU6gBSQzkjpUOahW
Zs88ItSe6oqwQGAHjhmcb08NLmuAzY7YzdMVYvX5zbtsKMSYKInXZg7cyiBQ
UDgHSWjXiRcvhL5ER+nZdhc9jIL2lv2p5/5Z2uLHIXSQ+0u1/mzNEsHbgyXt
zcofqNZd3u8dfAAid7zipsMTNYb00WTQ9i0mR/iT/wgEdXpFvCHDVHz4bOJt
3tWw6K9VjYPBfStpcDAR2yeqM40P2ZN2sHS37VHsfG5OjrMcYJoi8kcJonFZ
cyGOgkrIdGgoMCoa96zZrfnx0tCFhHbR3SRQap67RZ/1PEDfd+DyCvh9eFiX
hURFeikMpxiG+0k9Xqvz29FYht8nF7qrqRz6dBXl1srB/v59u32zv0bY3vjl
MA22TGb+FAgaKehEzwGk6weyGNefJuB6gkBLqaTfUa5hyQ/ohujfXUHJgcii
55ZRqxRWbD8xnMZ4OpO2OUt3tF/r8koskxBMLZ6pngSsXqiPtBXxATWxxDwS
ZabPWR78/muwHc/Ox7cb4W5+mmiSZ/urZVoOjgICEL+7jn0RXEPwsQZlB023
GQtbEhgOVRlBtQxm51zTNp8oDb3ClPvJVmFjfslQUSqiq0n0cB8x9cIejGqK
KU+qItdtF68iyM3ydBnmO/0LhztVMhZZLCO/CFOQNKAGInDyaka/bCYOnwOd
wNT06R1djOkigGxdp0gMPYEdHqIpWN+Ey9N9RkJK+3erV0I/oIAKF3FlWVZB
Ev4YchXv6Bo1mP2+nNs8gf1TJgStgcNYBK1oVjVujVzHQkUV+MpT642q48d3
Za2pAi04MVfD88NA0vJ4BIT7mQgxHZDHAAKhgxcl3rZDXJWwgSpx4zectPyO
Ov7vrV94CxlNo7J03r7v0kN73/XxElvEEvldbOFMCIfioeQQf+oO+OrtGZKg
BmvWpCtb4T+ZQrHCQjF3ImBay9FaDPZNs8AFiv61ksYuG8IZtDifOznUp4YN
Oh+AesITUA5eO/g29x4EJ/TbTqv9ZyuAzQT0AoM6KC0iVPYuNGtX7NZ5HL0z
+yFoJgmC1winMgVgFTzUy7mRXQm9oOCaWmdgPc3+pfm2mXLauumtle/Tm22Z
klqZCU1FdRYfAghg6hqaskHb2wqmpE+KnD+6dYR7I7kZYJYfrKKIKaSr4u/j
+bdFBEgaT2rXWYJz4KAL8WVg+/7j8g3v2bjwxeU8CtX3NoxQtT4F29F6zaMs
QNUSW3n2PUGS3PbkzxgIL/raKAsE33xWsWWf5KzzKZOOr4RXUC86B72To9hr
wijJcgr0JZgpFi7ap/b+Si9Nn9XUKrxSCocOMxXLhppa0lP/JB6lv0PkwDyT
kE8IDCARombcdg0FdqyidQQsb7pvDBPv5I+p0qRWUF0bdyi/NRfXtMiGLn88
Sct+Dxkwo76Hlbog4nS1O1BLa3O+eIj+DryHl5QeIUKXTbA9aogW5UssFbw2
qkCUwAiWX5KDxU1hzL620zpMjkDuTXavuKjjLsbsJi8LM1BqRHUY9nSIHFNp
K4LyJ43ZUTDHIgJdD+6/QWZohqrINs7cUqJ/AcI0LqZeuvmhixHN4OvUAbIM
TB08cONxYFLidr+b1UqETU11Dm5UeIFJXq//7pwV+RGNpeGgWZr9K0YKoORP
wL3SIDAxlIv3YGL7L/eKEniKQL6HKjY+IbtO+lcoiDBiaCOK+VFfd2L6rO8R
jVvpRYMHn36wZvCB6mb1Vk6f8sOkQeyzik5uU4MRiUQhOC1G/vfX5z0QtNsi
txkK+YjZOK7Gd2Wy+l5hUpPYt5m5RexZnHVxyuRcC9Zxz2RdajoprzSNGqdz
/4GyqnQeIvsjY/HqjsRAMi9L9q2uUAybk9YY/SQFm3DJMQBji9xRJiYKSBuo
KnxsI2NE1rSO3TREWojxTsDIOZoMIV9+UGu46vP4VbWjpw23Lt5s3Li/xyub
s4qhjp97o47ECjUC29W3jLmy/p9V7kZQumhua9wRZsMx0fsooUkR5eb/cG4v
l2CJLz9ftSEeUEKYar6n9fGJmwADYJ9bnqiAM9DM9KhfUefKkqavz0Zc1LCE
hejxnxHDdJYXiEdl4xtAe/TjNBtYm9J9cPyJwDHei9hen4OFTwC44XQXjpWU
cl8kOjF+p4vNAUveKG7nHw9Z2MjigMQYqcr6XIGQL8qiQoULC6i6Ck69ZCcT
QgzCeFKJEfIBit2uGOArNjBVz0qUQXNTrSLtVLZH5hEIfGmwJukGvXkOX2mX
N2ZLu5j0w9zqZBEOt9Q4WCHIoAMvoBuBxyp4kNkggHKq3uZdBf7BzdXNsFPu
EuQxDmRz+GJvJI40PMYFVbEkFGAwxiRtZYuTHO2XOgpVrz3snZHFhclErosh
3X6IKE6OIUcRDw2v7zhLJ3Mb/pdezlFga8OMEC1ZWOOsTibjhF5GTEWZy/4G
eNZFMioFU/msZEWtYz0JDAg2MRuDNxKYj1HERkFluteYzzpJ0o79q7TstZlk
+wKKwwA3r+RTjCZQUQ0acA1Kbh6yQxtt4s/MG9qq8ASVt6rHx4ok6Iey35HS
Xx4oUN3tauPrQIpvyx7cw7Ro21u9wRNZ2kisdSN/hpK7emN3BBt8mFwxpZkG
F2s1Hc0a0Uio6GsHRwC2jSDTsNLp/EdWtRzM63K4Gxxn4dCAayUF4iXpIung
yXd69VdTLbs7FwucmajrN9qbC5xbevRKB0UjJKiqJFmGvQTJjwcLaDfTT3dO
PGdezfiR6YZczK/3fSN/DPydPHGE3CmWlZ6GWm+/Vozh/K88AYtdcuqYH/d5
I7pSiSfiAlf3vtAn85TCoZq/EKxTV61Y462YxE9znxjP9hTZm2+WioMFahz8
VFQKDQPmxVrswrYF2nM9rMSCjXyb0mz+73YNvXlvoUaMo61Yna5+TGxfCT0D
xiSrpWivnZaY0ARj1e4K/+U43H2Hudzhc7eQxQ15jmkkOQYT6zolkg4L2pV4
CbN6V0QhTBRgoolGpjdinU/SMuCezUho7zNwxRlSq/muombUK34lQD20B1YT
9DMaS77EiFz9WhwoRFK3AxkhJSBpBdUzdGU0UvXs/VIXP3yRBkO9qPc+/5tM
hNthNBjY8IlUnLPhbdRpe7Q+ydGAg5XvqQT8S4WcEoL8LXsBOQSwBJG/4eCL
DMv1V9JbZYobkd+Au4VOWQCCKc4GjKovX+JO3DyvA9l6R2ezEUxNEmxPrhzs
0hOHCS+KaUXj7lSgMXinnoGDqzU816SpY14AFAtf1kXk7Eio/AjRUYKCBSYS
6C3ukgMNP6vjGb3/kU9Gpxf4CplGKLTS4C8A0yWWgjFF+inzdi7PSlNv5Vro
f5QUr+tEDt+d9D/JpW7NRvgfvZEpODDrSwmschMheCeTO821lPI53XJMLve7
xhq6bbrh8LLmGsVnxEvKoDxLCdKF1mYk3D74wvF/Vs2PHc90BsjMWDIKkRTJ
uRIicNEzq1TMum5XL5s6aBL8I5m3k/WWkv6YbubOBVsk/V+L8w5k2i+awhRb
dCD70QW04EIP0om+Dnj7lcj6OqNSPWHD1siBVwNWfAm5zjaB6gKO/7UgHati
TtotP8uuzodEM1tNtgmFVdA25vxLes2GKsOf4x84pMigdCwBo2NSlR6DLgwG
fnCQ/ZGVgIPUt64pkjV56AjfWU1VlxkPsJcbeu1h/uYBHzD6xj38t0afhSOD
tmQ40OUQ+80G8/Ad8E/Ccf4wPEpwGyzOeHT2p8YXA0XZvWDSciJkFIHCgXRS
nzUMjP++yTekvispsssz/j+1/RCJA3LKhtb8q3y+EBdJcFRgTsXitLzl+BLd
vwsrx39vLdRF5NCx7uksg+thsFiyN0U4PiEpAmV1gR+IBuRZN51EssTk7kg9
l2P79JDYGFYF3t//4CT2qnDsnUDR2AKzhBJ46SSE02+sSVZjXHdlkuMG26pz
JVMj6sKDD5YzaG35VwEjBHGvINeGUCCEladWI7tmBv5eFdvytZKbvyEKkQye
aMEiYs3c+To3jxa6bfeVas+CM6HDwqh8pWC09H5c25vydEX3gsSSHmI4Awt8
0+3P1jymVtcpZInvwwbBqa0Gzkom5ziMgcOaJXI7/UT684wBYR5Wz3v843T4
CnL0ky2omo5G9Yla2yVXQdWQXXgZMjwOo8WSVSC27r9h/NLMU1iE12yFpZvp
V8tTuonLHNRXKC/oPitOyYwZhvpzLN2JdCagac3eHV+aPa18fmrmTUdos9Fy
aSjXQ8XJw0WT7tP/OfdQ9PtoOfgAlST9a9LX2OBMq4ie/PVnJoqfIT/irZay
SzLNWUxkIB8998bjrr9WdpjWL3fc6NHMGrvdwXmCbMAWT4zu4xST9vlHZgp9
t3BMbfxtl/LwZkcExWGHLwS4Wm7NmxDo5ew+1c3XrFd7nzhRVusz166A3g4u
aMIq7vsVH/otzr6AsyI1I6kQQ+FBmiZ4tVdLuDsfIVS6eIn+gp3aJSO2hDVt
1M+DGEJfwypRsk445TGZY7R4OUNSiT1IPTUYj8Ip96xR1IKYgnGeGMIuJVs+
vF7z0ztiiyz/1VvS7xkAauIJ/x8eB7q16MIc+gsh9sWC0Cf44lfag9sNijOW
ueRQSlWUevGNaJOYgx7m4q3TYyiXdV+UFZPp8FKpxa/Lt6TYlNdWKoiKHxkB
jTZvna59ApBmCDeuvjyiKwKn2nFVhQsvm1Y0mqWaDV4Sk/FBO1WIETxoJVXr
tUDUVLL79cXOnOVNNoVDypsBwU9ZjubjkENKxP0jysBqSFntRjPWVs2y5d+M
llWHV4TNQe5no4pJYfAGcODrJorVtH/78BheOn+EOuCtsMobhAFPjiovj3w5
MpFunYdobSc9Ht/A7CYdiyKAp89WoDJ6EVHD0Pdmc5Cn/p3OJ4xOE2NFrSaD
i32jD+w0BqZ0eFNDw9PEu2rp2t2TBFPfXVWTeOKTtFl9UReon98P01E+3rHe
xlZ6plurDiJPwZ8ktOl1HiVoGlDpCgF2G4f4iPMOBIGdEats+RipI7Rtn8k9
nS1ctiQQwK5GJkCmZ70Gs/OQkKhhmc0N2S0vAbpIPiPXQ4EvxHSvhLJCQIzB
wKVxWYVHbxJFj3AS74Uk9AL9snnnzHzLbd1JeWVuaQ5yRET7vYnYXQ/o+spK
AULmHvqKbz9kkEzkWGThAqbGWn7CWbN0E82FR7V9QDC/SffAXhWrXSlaKxqi
9L9PDEoYeuA9yD4OK+a9Fqqz/lSbFNq+dJ27ZKE+S4ASKpoA/RvshNZJqj+w
COf3gE+PLpjRosoeiEQVlp1y7ny06Ya5Tk7pUEYjCB8GkcBJJ7ZQtug6gXcN
IYVueLoBfqkwcObunyL+mTp8Hmt0K7IpZcdHyBdkEw0OvZAkS/naFWh8CXl4
90RPYjCCljMbtNmVg3GY8noEiPy8XNMZ/ozJ8BR7WdhL0Gy4s+cKOkPJoE27
rnzbqmQz6fxQ+SjahXqehEfKdjpYX/GgcH9hdae+ks5EuRJ2mkHbvKQmyaB9
hE6RPcaDouCzJi30x1LnG+TPhtjW0lPev/b5qnFEUdQqiFzeYhLUHImEt9CX
+u8RixpROnHbJBH1GVuJxLAbbDQ3EhZK5msjn3lVDb7n4I2F+LeDsBbp6n3p
6sQ2nqW8Sy490PEmCd/5dTRkd244Xt7/tT6eitCGMqg5j7Ns7wMhLc8dDXEA
fQ7bOJk/0gsaAkQ7tbnFclENMtKPevqYDPBctEWccgrwz+3IPCGeSJzx7EGi
4BzIKkcHLafMhkuDrVN1xVbYh6gLy9lOS+MuIvbwSEKpDb+xb4OHRQUq1jDz
vTzcfhiA9kO+dOpJZ2X0QGQvV4D61ZoZfInBrY2VOLYUO+iWcmeo7YRPjcOO
+rp8GuYQ+5t6MveEQ/3wV47afY17uyHLkFCpdNthcJJ7BXqdRhV6cMbyV0KN
pFO3M27XvTlt7+urZw3yBwQ6tuW9WoxrFqH18k9WGiY7xLaYtRrlf1JTQP5Q
uqhV4yrT2pO4/vTM2NvZsGrOtKnUx7KcqBu6fRdG53tgaTocXtp8CY13Id2p
L8E7z9FX6l1DlIrvTIhihvc36NmKfZLPZOUkoGsQv8MFZkexF7SxkH9EqOWN
OMmwnIM5VvSlxry8OUpC3ptwZZepnh8bYaSd6tP/+myOSK3JyN81stAVw0S1
AH2HEtKTzwTbLGrw/IhJp7ZErv0Hkl724f7FrbqtPkeOLzR9Cb0WbIlftziX
nnkQzmKVNpx5ewiLb2CyaZ1KAWy8Ip6Bo8F5m+SrJIy+2SSknHbg1gKa2nmm
gGZNCyPH8cSPnSSMciTQhu9kAIJcK18qh3CAh5YUpJ64lmhGvkpscpmjIKIS
ZwY7RZAQgSFGfC7wMt+yAQEGYd4haSvKcJySFqDUrwaLGkaFStcrQ/lKWxRR
/zvijkiTd2QlX0WgnEj6BHxfbewIPQuAkWWljQtqbTJgtB65ActkMGcpLTEB
IeRHnOsXMwEOtbOBS6YqoqRa3IovCtiKOe/xZ/5/TqYtXG/EytgkBeTzXkWU
Ch8Ssuswkg34Wca8cmCo2eRBBgNoTx/v1MxpPVoFZgVe9ZsrDrL4xMROBV14
C0hIfNQ+ZObIiVDDmZTR7Mn42M/xXL+V+75DUJKsyEml/xF0mlEO/rsrwSWP
fj0E6j7ggaU2HYnRYKd30JawrxPsAQE91irl2nuY+4jHALbuy1yUdDiS6N32
nFbkMRccK4mkrfwTwmG6Els8fcKSSPvkKqBD8/TtbIu5+wezVhLoqLx5oTTt
SpfuTWemhq9O7T/ZtBU8fXtr4Yiopak3P5jGvjKuSsML9kqRmDEXTivmKgmL
HO009m+I/RXUg9bD4iv9052uV+JwkjLlJMU9PuD0IgBVqyxx/cAfU6GFutOY
FX2QNd7jgt/2Jozp02RK1jFRPkYJvreAvwvWiI8yUMFeePhIlUIyk875+rBZ
OfeDZU4Ty7GmIyRMrY8UZoLaq9SkNYH311lPCqiWmnktxPiqIg1BtJ+v1tyT
BAUFcKd9mHd8ydwe9om7Fh+21ipSYOhV2HmDNn5wVTCZ9hcGo0XhZTh8ImJw
XBbNaAOO4/STNTEyvOz9N8G2rM5rXQD8tM3Iqh6UrtTbnTGWdBVUYJqUCnac
GDrdF5YyHqZ/jnfTaKq5ZdZT4ydypytBIQm0JEEhpPwJzqGd3wUgDwUoMsAA
CqIUA5quQ2Y/aJLHPXwk/75HcJE63xSRFY5okLfgnXYVPFuF/j/wm2EHmT1y
tB6tG/ENZS4qKpEeNWP0tQncqI7q8R90AjvbN1yAwTjh12+lxaUWUUXcdLoU
jKT415mVRj+3sq3bN+8uk/VgsUbv6Vfc66BZk56rKVBCBEWilK7F2xr0vTKW
VjzAi6QaVh+uQHlCJp/VIWq5pXbMlghblXiKaKI9r5Cuo7YTcekrLaxQ5sAC
p9LnrZvQe8nBXIIqKGesf+chqss8asOz7pdRqNvcAiSHIFMHnX3ko+lZUv9P
VkAnHPe2/B1z7TkFYbh74YJMeho5M0zQr9kxJABOn+TYXpuysgOip6hnMX6t
nijzWc5sAxpdCOWsrOGrN990oehKvwkA4lKTLb/N9bxI9D7jcqw4IS2fOWwP
uif7F1aadQ+dy7H5bVavCcRUjYm7jtdFEt+BqoQHzEt2UAuvTPI5g1HqlGdC
SbzAHBo9LZJZfanzN1ZLbuiLsvz7fgrRM5Fln1m+iPSmDdLCaCHv3NGDRXkJ
NZx60hfg62PpVYYZyoiP45wD+wmNYDQFPocmufbL+x1JvMxAM3Cbo5iJJaud
cZEkYY9EY+inSZHEVb1lpDTETljyx9SOv1GtfboN7qFWWn1+kjcZeYCLO5Kn
oBVE/Km7muvaVhl19xAhpbWBr3I5QvqDjtpD43/Qstk0+zv0tyAi+fY37KB0
dDLRt0xdOZg+V0X9sTE+SAvxXsUX8VKfsNcDCgDqCbd4WHAw61ordX0iyGll
Abx/KAZAJv6G1iR67WjV9x4VEjSOoIK9l9/cY3wRodKt07T370+DXLcSjim8
yRoG+3o0D93YtcOtkme6p07KyKlsajPOanTbPFiMoQYnRexmNUV1K+eaBCWs
Kt6YoiiA80276EVNIitWRD8TOZxiOmIA1d6xBpWK8F9bUIsmiPRf6rYxa1Y2
AIKrYvGxIsLhiYn8HJtTjjhse8VjAmkBve0WefUlzD+wJND3VRTWvcGy/YBF
FRlleYIz5U1mnFjZQB3NzYRlmv77Rj2cqDLgrg3AZUD2nLBvU6T6VY5J0hMg
oRqmPgfUm0RmySDICytPV605gAKDpShL77zfUFtRy4AUgAsId+SGx18eJJlk
Dy8+LDX8T9D2YL2Q2RiOIzNhua16OCPeKd07kpQZjhUy09Mhi8Adg3e/WOag
9ouTAdTKZmTYBJxEf6v/3oBBZw/aYq5aviQ3q0+fnjKrbmhOj4iDa/dJTf8W
5acCkd1o9QMgEZQ3Y+zcPm5Ay8MT368I7HpBVyLuyUIlfvgfE7rrOPUED6gF
C3ELrY2StEYsOcBXj03tGE0MprbXoEYyP+BB2ofWGyzxTL/gcD5A2ljQZ8f6
c6Pw69RUVM7IJtLXzneUEbcEogmoNIeYKP/gR7sG5Bju9BYPIkS53AOZtjwq
BUO/0qlvPSdelqVato0wjUHIV9Pxfi/lxcn66ppymlWRBu8kSGcHQEhQynh3
ZxvYJBMcEmsDRW+jEjQRrEgcnpsmkwABrY1ncFo7Ftf0Tto9JwP1GI2zCQh+
UzWbbCx/6KeAkX/cplrjLD79+eJ5jfKJbEhJeqO3MPq8h1XxSAOB0Nk9A4r5
rVUzWl0xnER+zl8Jkqs8UfR5pjkO5o0qFi2Pi5NL1TNmR4K0cTshMIzdualE
1scIyEZf99VJ0TBW4GKYdrYeqCvtq2+hYW1Yfqu11oIGKoVjkrG/sORuebzO
/bgI5uzEbkJ6Qe3fpaV18CcBhPu6tFhEdjNQ1M1tsGGybe4/YoozGNWwjvuR
SBaA6vgM74QHRJwaEV8VXKD7cdkt3bay+niGTyyzmWjZkUNiIT5CBMQQkjf/
b1LNir4178iRS7wEvmbg4hqllBMqaSdhVJXKIuCzntssGh25LzmmeVG9FP0W
m/BuwIPclndW7TWm34DDa47whuYW6Ux/w4sEalVRG2oSfY7bNm73TnIJR9Z2
F5E4BsaJBO4XtaMKf7WWfJieXIbkaWTebBkS3IiO4PwBPovh5+ym5IbJq4HO
YE3rzZ8vX/kuC44uf2qqBdc2XyE0NyOEclGn/PnwFtG0cTDRlnb6QwYW0uvJ
ljk/XOEcBD0IcXKTfsCGa/9xp9bDUgAvxgyLsDpsWMs7D+Q1YeFAKrVAQhQC
/5z4PFOFmEYuGuqMkbDpj0GSWbS14L7RtvH6Sr4ODkFzlnoxSxbuswKeKWsM
InT3WXrqC7J2NYXkp9kHK2JQrAXozrm6v5/BvLWg6HCrokIcvpvo8DKXPbGp
qlNICH2Uz4Ug0nDOp4F++E6TC8ebyYf2/Q+p4KKUTyY4njw1YiTZDpdnU3iZ
6mOQBeY0FCjvcKrkP6C7yf89vf0u+nTG1kGnWV37BbzQWKvk/CiCuODMHNWR
LheKb25acw5hqdu50M8FADX+c0x8FWhANIYy3HH5gPxHeWu0ShqvNwcVOWt+
KVHwvsOfXR29JRY5EfLOXRmTnYoTUnMGBv3WiKfehKODks+7g+WKQCgd374Z
Ek8rOENZbsFzT5QVSLRXrmnFgF0vF7ygE+nkFnUxpAA+5nxpbTbT7yNi6dJY
ooGLtz3vn9GJvNdRLczO/wG89YR6Gpi2k8nW/GI4/g9SjiPL7gdyBUu2Da3V
5OuCWNGFVafG7LTVOsJfiAOEFGobrSvCh2fnJkoGHMAV8+oR8kpU6DRTbMNB
9xxs3mHNDhCeDjpUJ0l7WqZJxl31RQnsn0pgB0xyWt6qcd8iEDT2lyd3Z6hC
86dN5+xCC0lOLbalEL0EoohHKcDZ2/tTi32B9LsWgayXn4TJKyo0oIygaF5v
Q3lt55P/uIAGWIgmehiCN5PX8MqqighT8C0KU4iE6qAzxnooimeHUU3RwDci
ewVdqRW5/SDUwlaa25cKuTFmdmB57sld/oGaLQTWA8vwITBLNJmxOYspWx83
XGw3CO3dFSrAjDR1Hh35EEShiaEteCpFplC0eQdVNmWahxWD+n4Jq2sFIjZy
7kNB8BsHqpIX5r4aohKPta1iWxxfrE2yxdWx2TgKtg/w5gXPbr0M3fWuuIRC
PPVVposjKANsxMqovJwBY+9Tre30kbm90JmR9jyAAscZogBam8UE7Fr0ThKx
ztZn8hUJvQacdVmqK6xtVQfgiwzP0qnYLQqJ5oEgtaP4bRtegrntkgTI9QsC
MmC3yJmd7On/ZAe8pMMs5DDji/y7Ti3B7Hii+obHmYWV5ZCZg0oGPLdbra/V
D1qH6EYYUI7kPvnhnwLpW/fHidDQ7gNdbHKL0KYS2VOrunokMhNuBqVff1c7
68NHXtO871t7XyIjPMQpSgsHHCUFbVJFReAR/jbfpGnTv61P5KB2GURBBVBO
Kbw40nnAPKMWA5hC5Vn5Uig7G2VYr6i/HTFYr+HSNqeOSiSFKYXJitgrh+ZA
FLDEnffOO3ozRtbDGZZ4psg5VpJEZB/TAYnL84P2IZsi6Jk+CgIt2qNmTolP
SmNoxkcZAqknUKnWCbrFIU8gE+N6OFiW6CY1h+QvgaF0IFFI5Mxg5jRtpbzm
lAsWUjAaG+6HeDsJOAwOM30n7Cwf2wY9APjyzqQx2tsyIl9Tev/DbViOnMeA
PrMmgTNV/CmFWPEsCg8BNv9szFlJhkhNi6kK8Qc2OeP9AWXlJ3v8OBZU4Um8
V/EsIzDqFAt0QWKsMKSdcK61aARGCm+L7xrDxbFOLgKWNjQScYD/BYFlNjKp
NdsbWS0Q3FpePhVllzfmg+UIMcworZxVkZmPpO8in/PChsPDjzH9uxwmjBxp
pRi1wsJfXRsztlGsQHr04InKYruNyG3C6rGTRJ3MwnUGN0lNW9E9hXuNS8zj
sGP8n1+1AGWWjokFOvQcQiUlUZY2CrKNCkmKRV5PiNZvV7AP2QjFHX7KLM9c
AbIy+ogwGSE117Ar4rhUMLQzZwPNYQed5EfjZmKTCjAdNah7u6e9WibvNvbS
B1fH4FbyXVnISdyZsqm6jeYGukUrVwfJbYuAzWllOcJogGdBjFjWdcrZJthP
lZn1GJw4LPo3PvoCIDoWO3fkVdhRGB0m+dCINR6A/I44vaUEq2wYsXE5aujo
fNZsnZeddetA7upl5/0OZxIjtNMk/adriOtFcEyZ9f6tdEHoMFhlsMhI5QW0
PABBYsPSz7EEggfFQmLqqojG2iMDhfGY7csdaYhMlLMigSoZYwrBsltdV4LN
O5jFuH+Lbh93oDYM6XF8VyKEKjtukARqkpbPawfvORXLXUrqiCF4HfV1R0iR
mro3JVu5dEIksd8aQdQDBazicSlKiYJqEsBch7uB0SLlG3ygtR/KYb1tbnLP
DuAfS0ITIrpyLRuzFCOGVOA24q2SzwVSiZhncgm6adcrHdglDFOmKPihxoFU
cs7SC0Fv4RDfIU+5c8kM/lN9ij9nK+ONagJhsDxOCWBXy5sd2eCywP3IJN+U
Jaj9N8TSC1NKUCN0jBTvo9Oa6L0VlrSaAChYFTEU4IQQUMcBfo6aBEJeBZQW
ga3aeZT/jWBmL0YOQTkPro3jzcqKv0He4L/bfLaSXXE2sGXrJt9J4MFP2n9U
Ecq2si2/5JqVx4cHu3hcvvKxtrt9vHNylYJ11gNbzc6czTgcRW5zEQOeo/pQ
acMs6HRD5K+YUqpoGmZpIuL5fuC/Ekl6x7PmsIUyJ6bw3FOUUIstk/AsQaGF
1ITpZJ9aDT5ioaoJIEeP4bLC77die2OTM7oElIwXyvmxLoPesmbL0ZjjwPtD
bmB0yF834ZP9DYe7URxDYpT6gke2QbA41Lh/mNuRCuLFeiKcDY9seTEvRQf3
kj5tI0JOWEzN27vcNqFP/B5u2xjbO2n8blGwbny7dou1E8qnqnfUjj3ZoJLc
X7hiFX/bUoSX60cMLIvf+w+E8W9EotcLK9iUX6+KqG1gbCsssGxsUYsX/AT6
/GtAFe6TTKD6YmPt217Ni2b67xLRjGPfUAzD2ItUafjQN/1z1Z/8azABluT5
gm/VZerLaMly9cnCvOAj4hEdKcJpCTCOTPu5N5wvoHTdZTtPo9xU+kt4gwUp
i2pzAPjtZdQfIoSFX/54voqjZOwlFd0ezTa1sSahcUzbKx8Rx4HBjDl51mw5
F2SzQT3JlMngy7NWfParFKjZwONy5b5dtx9dM75uvrZCAKaoyJr9cv5lZfkF
LxWzvqDMU5yJvDOdV9eTFTUKt7C//NWjUOqUJ0OrjO1OFlCqJ7ui8iI3hd4f
PXlZZIidxEwLQKcuS/1nyPnf7w2YoyHxZiwPQ4HgzZhnNpLPwtsNEEKVwglX
6aD1UUkCI6LA7K/1vWPB6+Bqr/HBjq1V98VvJN6eTG2p+Zs1mmB6hLm6EGyp
cln/lIis2ydgKtl9StAd5wVV736ei6ZGd9WvZc57nc7SzLQrk3nZL8sntzHh
lvOR4OXe26ebnSng27WRIUpr2PN0ODFIshQnuFzrfyq0XpkTm4eGx19KkB3p
ZCql+LScJqTAx/IWpjQqLck7C3mDXtJN9zPQ6dSSMw/qtYLKQ/c0ASWMF2Nk
Sbybo55iuAXi6Y1UUn2ttgALW2OmA9wBn+ECHXvJrPXqxf4VDFzql/8qXg5c
uDL0da86A/KQP+K9AK51kXPp3eboIo2lEqawAVwTI70BQaApPKxkKV4yhzwi
WgmhpvqrrN9xiCA9Ip66VjmjKKP1ZVDFhpaYCjLZH3P0U5oAobfnb1D+jfzl
AKwhNQ5QEG1IVYvpdgD/owLTp5TdGURRVXC53ogMa1aBb6Dc+ueYllqX8u9/
/oJ8WBxBmkL/ZcpCoEWBwyLR3HKo93BVyWYnvP01vye723FtPIc3p3JuEATp
09jss0P8sdNJWQf8fzPNvEcup6F97Sd5iO2/vELsg/YNRcNpI32LHPI7Jf9z
gQ3bsM8weKfN+yJtoUiOnV33fu8bgmDncHlayNFpU6QCm95K5OhPO8L57YAz
2b6LA45CM1AicbXz49pZuUljEGfW0BZ74Q+9/1dmIUphtCBH8z+JphphW8TD
2w55bY6BTv4hyv4gaPNe8vzPlQZqofVFpbgexBCxJGXYNUTW9SRzvqDU/zlw
MKKjoPWt/+yXgXrT9bn6oxseByo1h00xYKTrTZgHkOyNC5zR5NI3blLFp3CQ
ixUm+T45P7/NMcVAjaYr6kc3qHdGPpI6KT4YPzhzI3gIcuH/dvdu02cIQo+0
P3i3CdUFJ6Ere0qRI8T2gVD8DUWy35vz17k4wLu781ICVMbI5hYp8FKfDDiz
DlQPNMKZa30TYX3ZzJ31r8a9mBlzAWKVY9yJOjRnXGYDPd3B20VNMvNW1dhd
TbvP4ZS8iVTxFWoSYrD77QZV+Cr+AVKpFcU+Y8GelKorNqlQldEKjewnwzz0
nmpBcFtK2XvgB0xa6/0VCHTAtJ3s6ZUD8uET5MNRcLvVY4E2+b7pGtvWJkd3
r5j0Yzf5xYIDLnzJ2p5Co8ppULzCJSsZNcstf30SxlZNmpHdMdaL9YOgFyEh
dTe1SbvcDzd0gcrvielGy9u19Jv9CFsJF+UFd8YNgMfIxGy2PnMW6c/zlrjb
Hy4YaLgCh+Cit1Tr3YJku/HehRsYa+Peo0Z2gSBWpdf7FcbJM2tZrXGt5wxK
Ftr/0ZZMvGs6V1aOKrOoU9ZnRlKs9mqCnNyJPRwU1IOyFETztMoh0xdmFyO3
RDkfpUJxK/MChjUj/a/POEmJWDWHmi/ENuZbW+vaSpLFI0d3n28uMpCNhKh0
w6gK/EhwJ8KiVZ0HCH9u7KLdjPQvhVztwLEDBWOp9TH27GLhnfmItmhMqCMH
8Mqqlnu7QT/yeOdwdu6obGHjF1D3+oQkMHIMwZ2J+jiYJ2TlEV+44kn1Vq4h
RDwXmLB+XrsGrCiolKf+WajG9k3sWt7sMYyHgusZubk1xIcoIt1+/9dU7ya+
58Gvkj9YXZ82D3PFB3PUin21IIUWKx+VQOf10YanX6/QTRQ1WFzGtRAe69JD
+IkWwB/G5ay8Dd8uxq0K5FMvwEnO1AQSpa2gpF/n5ugbqQS5K3ZSnpdo/pov
YXYoglhXRpjQ9QekR2XlzKpaa3K6hNCMAo1hJji49ICkEPOq93p3kCzGCosR
cn/rg1gNxBu+pivg28OwSrxlJc7UvMNBVAx6TYzQb1GdboXSwyRo5nH3K7YR
zwQ22KtsITJAtNh5S+Mt3lrWdb47fqiNhQiNDDk/Qzl7HlNGsbRtzRU9uMx8
z4cSqan7V6HNkt3+GNi3a2GlspOIknSFvnmIlIooaV/WKRP40UbBgagQA6U6
Ng/bREU0xW5HxNnXOBdHzh6uDVX+IcAplu8wNVonddl2pfA//Lv9TKpcqoqF
Z/EO60pddirtuOlwLt+ah0DBvPWqN0xHax07xrJsxBnlP7AeqgOv5dVIgmuX
wvK631idH8sspc6DR4mpSBh8njYbLw2q2r4zCoBMGmZ/USauopjRtB1LwsPd
m0ddnAhGnL8qIPoD3dSPvPy0ltKrTPqReTQ+5n1g8JqOYPQZRUraoXODQN3q
ABVlXMoim0gsVxzNwed88XAsAZL1a4arnR/GBbjHvvaqyQvgPDHNZtLFLJt9
fH6bbf2XI8JH+QJ2x6MPcWOeocV/HMK3egLgwEZg5rNB6RU3/1NYHrSUZvJ+
8VNm+Uw3n6dMUv30yetPQNxyjoQULnq5injSJjeMCrbU4+QqfEj2zWmwAutQ
3NMkl2+GBV8niaylkfqhRZ1SsI2FQbW3+HXMzww6NNCn99nqDk85t+ByyTrl
LQOAFpan72xsENdGgG4J61QYjB62bHO51omvtbUCDJE3f5a/AlzQkpkmIJYG
jgNoAlbQVj3XRh73nn+3mOjFznldNThAOscp4g5DMcIlyE8G2y2QA0STeSdZ
qiRxXGfiDcPz2ANVRrDQ8IYdxn/HNrj8zuSfymUAn1odcqFppIUqYd/cxccQ
pToH+WHF14VGv1Wd6l82JRGhJNbNfsP3XQhvJ1RtNZIFdF9yfxOW2AWtKPxD
scjOy/vSNoRiAfdfGAKJoBhIfoaspRf0V8f328EFFF7dcFse9JprUQDojVEA
iRNwn/wpwPom4Zrqup0Z7zELv8CPdRI6o+j6E+/uWmP//STP6tPa9nr/J6Lq
bcSPLCj4HCnqAYWRmsZSjopKGT+J1yzMXVvzK2EcCJqFs+exE4L7YRPJwvOP
BhGhkDMCJ8m+yktmI87vAq2NEJY5EihiTP8t//EM6U5+0hN9iKUmYwIw324p
Gl9dqJzQA+Ab8hHS+xAD+DJtUfJ8QIupJE0L0vaWdOEnJJm8/f7xKJryoPpK
Z6ct5gmm5F1awRFGTbLGGotgTUqVAmGz1JO6znLnu7Kbjs9xBDENnubct7qr
O4oAp+uW6qJHqToM9aTgPxN2T9YK1cDtoHOeT5GQ6p9X6P1aQ4DjiwKOG85Z
29N4t7h459y8b22U0u4pPzZHcFJzeDJbf3inQ0gZ5lCYRrdMyL/ff5bYn1mh
ERslBqH9P8Ls8jNpdlLmQsATToCErRryf4AkJ389vNaPbnEERJQ3YO2TD380
03HUiLSMpGvG6gVEOxNZPjIV9YbtOoSPvLLDNbzUwie5zQc9IEvGfgtrAK6q
BlFa3UGuoY/eXfpC7ENSANePqYNofOaTgpLtITUwZJJwXqIYZgPQmDopUNcd
O3AqwqEdZsFAUMAiqLuTbUFnOWcXAjNK+0XhBSpvq6J+N/QeROmtI1e/cooI
OILfrWPq8kMP3VQhNk2pMmo3ot6/l7dX9vUmdWxZFapq3UQ45Ed5Qw0MSADV
S0DPdwMEf21Z+bPZshBjCS5lujXxvm/pjD+uvjK3s+YPdtcf5Lhs1BcfUH++
KpW/HGTD3kPG092prBLhT3QcxWa31/zTyv3vmA/4oQR0uNuqBYvH7fecCu5Z
edsVxmGGXWcupA/78BdCud8pPmKhQrKT5ogc4vg+Y4FHnchIeXpLuQoRTrpa
KE98AhI+wis2bPVcXeujNZAfHBBLBxkkxm8f6o/0wQ4zYnu+h0xYAZZYCGGw
Cw0ksm4jYH0V9pBCSkO6GgA5EPuBH+4yOcUQC1buq7ICzm00jhtAeN9mxga3
NzF4m3+J7zkoPWdl5h9fBOlvv8PcG9AY/AVJdF7kmUS2aJHONco/TEdAuNGB
/CkptbVHpJ+8MU73rAgEFXJRIpDh6JUz5rTVt+Rauhu6tWYMKw0wxEJvvlrb
anv7IKtlF1vWWsCF/m8siJsiPGCQ4GS6in/5uyBgP8504UwaOd4cOcG3ZQbn
KmGRB5jGuoKf+/+EDpRyb+QeEyYPc1/deWK6qwj6/c04br8mBSwiCCjzNGmD
+w+M8TsPiF6oQb2IBIgoCoKxsSSu4o9GX9PdkrFTt6Rhp8teYIO0/e0IJpa6
qBU/T4NPf162RNEWWL1sv1vx4yuKYIGjjZb/vSeuIUc/BZOgfhE/gKnow12j
TwxwSEGXaPZ2WF+i3jjrpDNh69s3x4RE393HA2NFHNWJHTb6myztPY+gGubi
R6+OLEPlokSWL62KRtTApUhPPHUpV2FtN1X1ub/35OKiltzT03WSS+e8ifBZ
0K0ksmZtbWJJyGtwg805Fl5AHm7kITqloyMOEFpP0S1MuKOp9NokUdPpttZB
LijaUgMtA+IQ3tE01ha32x5ingCaCxXdKoBPYQk3tGCLXOlgs0zTdKIaktk2
qJpGYyD/A60jii/c6z8VJrgorjPXyIdbjtjr2u+YcOntOoWz7vxt1bKeP0tr
bnrm5N3+qTHB4agwSiklC7p10nvRenBcN28hSoRNkmWYP/EgZJ6d9+HpXZLX
thC8ads2BkiGFQAMpnCmFQCg8gjDr2V5ze6EsPekzeTbyCIcmaLxTMX9iKmU
pcvEZXtQaCYSH3CqUfWxhg8tQNjc0gZtVRZZxUPCGY36EhdEvpsMW+WQP7K5
Pbk4toTSivAWUs0MTscLAdlvW3MjzpUGMXvK+GfMOB44KHb5YnQpxLlnwOVb
/sPnRGIKi9PDIs7o3Qm9hJ9KGfG9u8uEFEtsjXq6XCEhxP0GKT4A5WFKHFmx
rsV5fspxmU11cB7tKAu+K1Thqo9BPyubfbTQYN2PAdCDnAHQCNM8YMZrwo55
k/k+zLb8VbpyoRjNtx+kZ8KpRdSQqDfnM4Yvs3HLm2PCuBVbtsm1xW1BvyR4
1tnLsw3Csc9c+i3hXihVxVKtGcTIjj71qDK4oTNsOZWnexp64hH716KHiIDr
a/ehZZP9LblosqGJTO027Vn/ajEkADX5ZNWPZoRPkRCRk9RMAIw/tvXY1YoQ
3Yko1htvpjaeECh3FdxejRjcIFsHXdDMxLZVEBH0cn967WpPRR2BwaKmek6Q
4uF8TxaTWcYP+8txau4aBMJHxA6ukqlhyABIDunHyVTOS0/CPrzlo3ao3X6a
E/qbudOaKjLPTsRLgmD1nd4XJgEl6jLy/pPSKazMGvTIV7Tv1leOlEqO+Viz
kX11W8fdhPLh26i8+JnIZXR8guJgVwX9jEywKY9AGi6W3y8bk4vkO6wxW1de
Uhu+Ju4Tagz4Z5jA+n8rVVP1MvB8+qcJpPfAS2rkMFhKoRYFkFypXLP+Qj2I
kPRtFkaLOavFobaBwq28gzTgyYtheqXlL7BSZBqaJW2U6Q9K1nhaF2RKWLqF
Oc7vSwTlhskdDQMk6v7t0L3eS5YmvJaj2hqV9XSbOKI/T5o0KTukS+AwapSb
/qYMCQmUqsBFfDwTY0OUVlrfIJg0/rqRxY1XubYCY2bEFAK4u4bwqCGNZQ9B
9gB5ETMCchaADLDJkm4AfZ9OGPWuLbqwx4Mkq4BbMXPWq/GvZE9lZ/wfdxut
4WRc1wUYrjU/1QXr8WIbozliEovjBUaJ17d8c6EAPzkSUkLh0rtkNwBN/cnw
g577OmXLcds3JW76sfGFE6KUq0rGTzl8sSKTvIkcgnrpAT6OpKMipT6sSP17
ASVWJNhio4Qyp5gzGkEG5KUEPRBsVcuELwm9vhnaAImp+m4T/Ns0XCRWu1KB
q0t/5eP4a9lBJihs6ONssclhomvrvHqQA2+hjvaFMPiLihs7W4OVdtA5jdZO
D0ql6R+VP2Epod8HjIojp14otKP2NHSd+ZseYQ7OnLt5lvVeuQAC8ObxT9hc
4EB4C2LZ4jsOT4E0U8ma1xIMfvedEybAGIwkdCX7HpNecsgV2xjvDu37CTbW
o8ZEpVTCYt4pGcol+Oy5jMz81eIlNhlssmHC/fUEXtYO0teIR6q5axwBAWqg
xR4XQQjN9SU0ebIyN2znoh9y3nXBV78R0SMZh2I6QqeykmhBbEhmUdO8Dtg2
br9ITdpeI6m+7Pqd+3OxSmXIIHdwWhFOeqZlT8BbuDapWLRNzxEluSn6I3Nh
pa4kE2fQ4OvXlpiPHazHCcgIspS2ridXGPrDqhBA+1OEMHGQq7XTUD3DYMDH
0Eyexx3wCPYl0ApV6bpt/AB1XJxwIFDm+IBeJYRebvvr5w4thaBnOjb9GHEn
9LaSA2i/AGWLhOdgdYAjw74veZgss3Yig2u/vIVD4wKGnMWLZ9+Zeo7JadF/
gQ8s2NE2pesi9RkzkpkFEKDqWKTOkl5PpURIZB8oB7/mggbDyql2q96uxA4X
N3m+uacyL9NC/xC4VtjPrxtRfc/UtHphWnlHfUWcyEl8gdNS2P8P7lbL9rmx
VVrkHEIDAmCkbqhfykAB3kgXfXh6DhK2QPBMtohn/HAgD9d5W/tWelbS1c8S
mNlhTzSpMSwSIw9QoP67T5XRoo36GAEjXsKAF9kKY0Kv9KrW0GVukfwBxZMf
jap5iEVR+aVJem9udBTw84/nUKNXc3CfszguJVNXcqYJ+bWT0m5romJpfGjC
V6EO5kSgQM6kHGKdyetCwcwRmyBnGDaOd97moprBsz6UNA7/r8v58h4Uv2oR
htWm4jGqBUVQUtl3FBMU/zykOPgIJNs8F6JKwAXVnorWJdoWMOrp7NSmCf5s
uNs1eo/NQjxveJs4SYuAhuUuQc+7Q4UNE134zJM4MPYfrQAYf57XrZcI5iaN
S30pVATBKig6UPLnvlSlSLLIh/buVCX0yAg4QqsQIrYI0RrVWRgRQ1ILPXMo
eSEktub73IfsXtU598b/gBuVqFTpzxq4q6LAREj0T84fN2E7mK6ZImXXmL/o
dELk4aStzBITLiQ2H/Mfqw/RYQOuSCsqHhVFnio5vmUy1xFEv6j/hDhogBRr
wiA0MH5HVZdMpqMhEVJ/qwNOfnyimn2L8gMXUyHXRmCrPpe+8b7Rtm8TaKAq
sjrYgwqlpetesV3Fg3VpyudbVSWrD1YB+HJff6mT9N1B3KB/NxtBK4/URcb4
6O1UQXcqYwq4iLZJ0p+Mt/X0X4t3lebuILrFHpNnAilwOAJoTy7oa4UGjd/S
ivRae1byboaQd9gQ1ah+nMBIGD9XYdVx5pqsydZOT7+j8DRvz5MvlnerqvVX
wUectTcL4h+7Bs7PJ/La0mU1KnQxqRKOVzTx+aulwxUEvX5lMe+5dC7N7xDI
+lcM9AavNsjNuzwGhRclGQt0TFdkjJqwiOQ6b9IvqoPZkL24xvDoEldeD927
T0Sj6NDR0VZYkvIRkIBjrc3XKV5jwA3BJxyNHYGT2Z/hXPJ7EJHKfIF4vo/R
pzFD3CTw/BA2p/BLCDkiX39XP0Ks3xdtx69dvF2yfzetTXEzP+V5HSa6TING
DCsZLasbGkigXlQEObf/FnKgCK7N8f3KunNTCKIhIXbb8Vy1m7v+HR76ZPnW
2iotvsVb78BEy+ZfNFO1O6j80NRTyPVt7CjCG3BQXkOhFzHuE3LMQWYwvJuQ
zWRTVjs+EWgfTpc94cLrTDVXwo4XmYNNiaV/Tv/9jMvVZnlqVomvVHCRFLwh
vcx2QMfoLM/I2Acc7lbyVYXqjnI97mThTNgXI3/9gyq/nba/eUi6gdRrH+nP
3qw/I7sv7q+mrAC+hPPC87HPzw/3OLv6Dmdc4sskRADBFf3WDXyogRsb8zi8
OYff28iUm367FSWIF/QcwCdJQyCxVyxh2Ae4NkC2Ee783VUoWDzoP4BkDvZQ
q94dI7SOpJew4VbdrYropc8nLXVm2XfsEn9havAoeszcFbmoyUt0dJAYWQ4r
VoynY4yhfPHrfnZjfTRoE/Bqdr2SezmQDzNQTvbAvUAzEpnXW+fxrTTDJUKh
PcXseFqmhAdprK+yKZFspl/PjhZH/nDTmeDSfWvzQ9BxbIUSwcesvNYl4Iv7
6n1A/YJAEFqDhdESAmxsVdz+aXDFiehap/AEBrnWFkHPnakBHufHm9oUyHuy
10rqChfXsVIv3MJF4SP/jlGjcvOi7tHRmpOX6qlA4ImV9Qxg9LgE1i4Phdw+
JQOFVQbsuG0dBWPJ7uzod8wsWiwpqqynd3+to41Zk6GPxD7WJ0r4rtiCgKZQ
y7NiJ2kMQKs4hMDBLixt4VHzRXgETw5dhhDa9/60cPgkBNBFXjvRpuFVyJzd
jLR6leOI6Oe26cKJeD+t8ahQUZ47599UbHcrs2/0HC6802tQZthZMgKG9HyT
P67cv1lnnWuNKfvZ20IOgHT1P/n6I6A9pFRROM7Y0VJnUuFh1sT4fH+2xTmq
jPFo94esZgpFSTrtrRUxkHtVOkFAYukfPtlUlwa+ioyTXqz5XDD7Bl9JcXNS
cf3ckSH2Sc3TGzwu3nRWo+WpTf7v+s8ehYc/VweKA9caWI+tU1cb60X0oO7z
BLmdsuyCnbi2E5Fc+pPHuq3iQQ1+re/ycBBNE9gavC8YtmH9TQfQ50U1neuu
CPIjSDulW2OPUMoq6WWXCFggXVIgCqA465Kapc34i8wYIfZ6uNWCWrlCKiaU
qmctJ5jfWA1pYACjcsyjtdl4EAEhKwUmYO84Ylqik0fBZYdJjcSf1yWbx4aR
GF/QyN79PIChDhRBWl9HWe5S/qlDBJtRTyri+MCv+Ty6EFjhlF2hNTts8nva
IU9rOiPidNHY+1yjWxOfwgHauDwFbV0sWMbc+HNlLai9hLJegPF+XP+KZlwr
xnJ3Gzp9Pr0WS3YjJWpJvqwIDak8QVTOwtJuq3niGgl6Z+zHb2N/4nUzsg39
66SG4LFRbvxVL19alrlbOS7iGGM5qAyKCCoteQsQMzyV8H8/nZXi5i5YIsaB
l0A+iR/FIDWS5A2y5Vh8ZcybhUcMCnI9yCggmCOIKNLDob0MasdjFpgYY95a
pPKNVrETY7l5diMQbElrF+LF4+qYOCpH+D1vpmMU+1E7VruMYLcDusXj4FGF
+poepSPG85dQqEbuHiFM8tVBtou4V9HkqjNnhN+4eJlKtBgl3XFZzyAdwkjh
hbueUQS8GULxvhQRAxm3xaf6+nDspTGoW9xLNEKIaytN6XdpR3sit55ziVIA
ew1sSnlYQZ5gmFgyVMsdE5M6ygHef6BD7nJS4tXdvYjE3agJMMwWZeMpwRDt
M2ZzlQUOcdAZdj/Adrt49H863e9Oyg68Wt21qo3x9k73K5m0DTSOU2DGV6Bg
Ipiadx7XZ6lLhWS1HiDXSDc5AFi+fepdYV+oNIuY4eQ7IXWDzYrwBcXoddus
8zXQtSoorIpPkI2hpgkS+WnPSG4AyJ2twaEVsuUNe9mTLLWZYHxIpS4QissI
FNLJv8laJ3t0mlhDeovQIEgbbehAAdUd7NQ28XucuqZOnHTph3YCCuQTpoen
M/yjDyfLL7YSuz3NDDCtEetGyS7MsNysHKBq19k8eNaob5NcY1ZIRxvuzlhy
qD7SNZXcpOvk3SrPFDwN2gtdygkEaENNQxl2//Q7CzJ0i5AuFM26xK+PniIg
0u3Ao1fHqv/G1b8WreryG0blVvXv1oHw3CR5SBfnbUutZ+GeAo4e7/4K9+Px
NFxiqR5v1VguOElodA6sxMy+sREcWfoIWWx4tVNn9jafYjd4Sp+SsWz7zwkN
pyo7ExVvECQOxEzZNoxJBZOLXC86iWxaQMM6ZpcvWFeYFnXLUvPUtxs+Aozk
K9PMm7y3nBzY+mlSMmVyIQfx505H8+YhqV8FYf1vUhyTkDM6P7rxHECuv1Ye
TYN1Kz9WdJCx/RkoDaKiEo/4ijFGOsTz3ji23X51EjtRmQMsLPTBXoBi6CaD
qnwzfbNJz8HGmzFUAE6L95MhpV4l7no1GoxjZ0IAkQ4SRZa7D91wQ3Ak4aul
Ie2aXaaHou+9BYAy7TS0mxJJ7xdE/0HA6ktoDzZlQSr4sJxgCG2sg5lRl/et
U6SVRTtDgieTKRs5nbMkydmtTjG8DNGRVAY9SGH0EWC/YZcotglJdlavP+ny
vYTDlIst8d+3JBVNyATyGgGPcQdtos3yLrrrvG/SgwAA4WNmg78AvLpnCQtI
3bLqExFjHoB1qulO6l136fdhwR9OEVwbV6yAYRM7+MwoDky+ub1u58smovCz
BJQP60otBFKTRTTFoJpy2MUyGdoWPUUzD9/pQV0uFW5a3uh8iZ1TFV3rWQ5+
UJDIUsDToMDl4mYfSItO7zfgmCz4SS0aZ6O7CIHJhS5m9M1bwAyjev+M/EMe
krJZWtcJCrdzOCeZS1H9lJxQX41wi64oVwE+ju2Qgrua3WtYtjHUGrh8qPRP
LfGLlnehE8csEydxNs0aE4gWjxnIZelLLEUhBp8H8wZWULwlejeO5Qv5P/DL
0sabS0vzt29gbjdKbSIyckM2TNI2i74O8VDw1yszqORjc+lCSRZ2HpP3njMQ
2n+18LT3Odp7ejOyoyb4XF1Gf2u8WzcoXis4Zz0H8MtmQiXPQcuH+Y3r8vae
jXcxp2M0Fx7tyWguNQPKjb2kHoweTA5EA0GyU460l7dY1J9MEK5bpt87TNr1
EDDBGhMs3djMoXJv4x9va3dVHpf2u19wErbTIL2DR3xn7xAfaW+N2r4N7+UB
RF/TR7R6yXPN65gkGCG5+QG4WY3sFs1qt6pCH+g9TBTa85i0U5f/TrJrzQP3
T0DybWmWeHfFj3VC7OZuEcY/2OnWfDyWAI4e4BMCdZSlPUvZzIj/l4uHdP4r
5k8uM+MXJKLBVIFHOjIiYMcY4paqnVKzLuZknm0ZhCbsxE1rzxSmfndzwpf5
yvlizPFdYIVQTT8X8YTsFJsymHn3D88K+Lyeh3bMkH87K5ZNOq9tMxqDCqBT
QfGjrHFUhKg2F2WwyFxnBWtwKB0NqiPeBntT/OPnlFb+rYz2LRPdAdtVCl3M
Y54VWMWEaUTYemP+cf6aOZTKi8KWEjbmTiwNhigfULIjG4BlmYKM10KTBbJF
K5LXeNcH+2HfjLf0EbxoqmHQdnymEw/TLLmoZFLTBQkm2RJuBDDZQ5m0mRgF
vLlqKi0dXFYMAwhaSaX7bg6QCIQD1G8jwpXm5lJRkfqeK6+3/i0h7ICnAlKu
nZUAgdlig+g90LXSVPsdIEEeGXHRNM1xAODo3FRzQk5FGbwPP6JomXu2iIib
dtoK8XCiePQE+jpkM6IAa8Nv1dcDiim0hXO+WVZp2iGM0+a8VlHhHgDJ4DA0
ilOZa8erHhrCxA+ajA8BTZNa08UofFo8sAGPgGqTDPz2POFIsPBL7gJep+7I
PsGW9jS927tn1ej8v3Ll2S8Oj+Z3H129sfcrmI3tGVVZrTvW+wIPQkR/VlLR
CbI0wE4GT+aud4qZ+yMV66YjkBeMw9odUc5ZogLeEDZV0ExHHLaB50v/mFdm
q+O0CCZ1eNFXLUTrV4nvQ3VNqRjjTQiQbu+Lqjjdm2KAjx9KpUGaqNTPBh5P
HV96+FNy4LweCEHeKe9hcSTLycEBYxUpwT+uhtZJ8W0BKyIM1eLvMfHo0aSN
JIu3pv1/eKhNs5Ongligs5cd+r3iNsdfgqi+u+rHN4nttPUlgyYu7y+ZKNGZ
i84r3E/aXmqvH6J4lmjkqpra2O21AQv4vAPdDFrvP7uH145lH8jzSpO45OYi
TwJ6d81OU8JieXT1/5r84SkgPaCLGJWFUwCrmzi/4E819pfPNdjB45Bq3iWU
dv+ozm29GJGjTHSy16IDdY10BhrE0HVKkgj3VFWuvEoHgw4lQst/TIix9+QD
a4uQih/F14MadTLtr6XzlEhtp2TNWnUfk/HQfHjOShsLXah7ObbTC55rU/iS
TGnKE0LvOS4lrqigu7Q5Qgoh2W9MeBzunUHFJr3d1mxG/LvzKlxT8WiWtezJ
4n1CHlrDLss6d8PYmrYiLzLAu/vdMv/Rei8tJypGCPbow4GjE2httF3byT58
kcHz+6ukqoztkXHYshoP+vDyXo3dC6wETSkd0iVUyt+WSUGk6tFEpGVPL0bn
0xc6owUI4kvsunrSjV4VKn10oNBf1Hx3QeocvooOwn/k9EnEy+gb+SGMMJnI
UNYF2Bi7umiAgL9sAcrPd5gZ4+8UbE8JxzuUJAVraaqrBw1fX9GvsTIfdTOO
AIc2stenORGHlLD/+DGt4m/ZqO8geeUfHZefnTKSGyYxZACKsZNJcjahxwRC
9y1NJiU6b8YOt6nPlcLsDXrDELrGUjy1ssyresEfnAtx+vm45T/M7MivwzZ7
evbyDQ+xtEA3yjkraJ8sprvAIicZdo9vBwv9DiSqz/CcTjl1/rFv2MlqZgx0
LYKgiOuWvvrZFyXRTNV3E/PvktgttobPf1MO157h11adYZNBJQ51BJeeAS4s
EVDx2h/BjjoXHJ73d5ocAvb5fVPt3wmt6xkTJf03cVeuIE4jkVWIPXj96WQC
XUSrx9toPM/KlWHoQq7gvPbglFsTIMPzsOfxyfJjxxropzN0GO/uUea7toZa
6Gx/hQA8cj5jekmhnNOJboUnwqHGWu5FAsnVRSivwuCcZsvlEbT35WGEmoom
H+8neEyhJJKGNe+TA2Rw1GxKXHOtO9UPaBrrpGYMLiR4MElLD9oeiJYWafSs
h142vhIyNqRvZ9HGA+30DKVTOJ1FCSXfHzrVcKAuXRAKe4rT2EclOg5/45yu
urxT5+WEVEWkEU797vXxez7KJpkdN6Y6NsYS+1jxsyPYHUGIpqGXK1cCNuuD
ThymKTWE6qBOvyxDDIQ4NklTeOg+hqeEb0jOs3hVXK3wxQCk2DGMwAlePTIn
7SZiKF4tl1b4r9tX4o80MLXOmxLb/SCWpJO+15/W7+B3zjG1LW9Z9+jf+n12
1QkWC8ToWeHm1j304PMA4m5I1Ry6Q4G21vi8bCasva8wjZ66ZZPR7IazQZ2+
A52RMOkk7Hb7Dbma+7hXsuNNuj9jVp+8ZAQnX5WzL9UP5luHAna+Y4g9vseR
OXPZyBKFnca8rCrF8CxpdWj/1HysERIIqwG5QM3T+4YVFzshohHsR5WPvYUG
mvIUKajI4iMHJdh5VWG+/FXA6iBjiXS+mR3L7uTwTaeAI5aSoljTSIn7p0LP
Kyb1tSlgjFmXUjsuEEQmJs+PA3PSpcv2pSgvHxlV+AEX32wo9M7pzIcuwfhE
fL+eGMBUMVhBZd/SKc20Of1uxCZbg5KnGFiGhLFTXpieMNcj788FcDU8oVFy
KMxzeZPHvg0+elBon8ILGfbcQ+EUleDhsIrHzKX5v9kN/imOBrxy4xGopl1v
pkegUHvxCvptuWtlm2Dc/x/0RylYbSKRFC0Pcjs04hyRPCDw3rcScFKPrz3U
t3DNLrSjjHXINLvYFqJx0PHBCU6Oj1UlSkbJ9AnCzGu4P44S9ivI6OQmN1tS
KirAE84rsSeBiviHZmzp/l02DKfyFoudFw0tOtaxazlrZmj+GYawlvNasy62
eQBW5SXvcKHQhIOCyv4RE9npSzK8gt4EXP+AzfCFGwKQvyt2qbo95F8x4jPG
KaKWSx6pDXoeZ1tC5eYFI9nEgV+m7DVDC/UHjVh5mEiXDY/uVaEQWK3LqOIc
ug5U8YGcfDY9WlS7ZkCiqbzZwM9/gMqkB/Z3nug4dX/cB/1nddNdA+nJFAoc
+QMi7IFcMbiytnr6qrjsmxkt05kLdq3HROQTgWm+8ahaitQBdovw17Yr01tK
QVe9lm9b8bH8os1SfmaoOEVHJoOyKEAGCDa2V4H8J4tr4ssjpIpIod3RcpBE
K3VxpU1dewOqykCmQtRdtdT0zBzVbDHWJ7Bjeg5EHDM9zgdOY9ecflFiIeX7
CzfEMomdu/Uyz54x4Ui9wGJ2TOtdTzF6BaHoUsokimh1yBt4XRhnl4wR3qK5
eP1NB+uZXZ8/y1sMolp8qqgR45Y9dJbiPmEabUD7NqCG9uQnKL5Ov9K+lQCE
W+4x9lf9Yb9L8BNR9qZ7Y0ZPkxttqL20EUzIJSunKK6aAGQ6fJ2fuVr4GTdq
9P9ewEUByVI3b6t9diBMtAVy9LhMAI9t2pDXE+4F2qx24EGRpAo3RbsGEKTY
RbEQ4lkrYumlWg5xpElXBVB3DZw+iu99FNVHbUbqMqMfCLE4C3D3WXfiookm
i9Jy7NgwMh4Iq6cDCUlVB6fzWA9O1m2bZ2Z54oUWX38JahZpK2UKAryZvOTk
YwWZJW8z/2O4b3jPQhLly3YCdCLhL6Yu0JAapFn7MbzOQdOOGskuuGQZd6bx
lojBjL61rqL3BHJ9ka54pEieOIHAOmoRdWgRUpJGpTGrfn+nrokpdZTWQ8x3
FdQgaVHmpZbkLBXQcdmak/wySshA3ZOW4AqdP2arRpon03bLxuRk/Z5ikdBA
uuTAVdAg3sp1evm579zMbGtBL9K2wQYE38Nz6orVDFknYIMXqkBCU4pyNG7Q
885X/msfM5YouDjfn46l4qn+nA1QSDlI3PLd2xhG2dWkavk8zh+BHhtQF2Vs
whjfqttLkmAiITNHIuGaRIJMs7YHbuIkYZAV1NKushlpuPdjF9q1maL70FX2
I80aknFiEueOEcsc0V3g/7cqPsXmLPhX0VmuEzmq/ZRBuVXiMnoEJW9sw+4I
oE9Nj71wDxmM9kXnpGTGoZPj19dF7TcupqrxLwKVZT2iezC97k1Lpej5gB//
Cpfa6gQPlLHDOs1hqfTK4WWrVNAKOiqWICniK2YBxWdqFSsUNWHihHBZtafd
ddrCwjGUB9xsLi+gmUOnYHI/86d3cOIrY4nU/uFSMU7meWQvqSxeLrn0voXi
SjZZcXRHbNUcBJuZ3W95hJxbR2lUeeiQWYouGJencF5woylTlZR0lm6O05Cz
LSzC9BxqX7409mH2GPgcZ6yt+V4rtPPCfW9Dk71+R7psMoz2bv16Ga+5SEer
Mwsv+Azc80drAalon5ibOQrg1860t/EqJejRm2/QaLoj/JnhBWHu2PlIyqK5
KAZbmifplkFXiEweZmFxPnOrQC8jZbWNy5Zp15splJB6EEeXMoRkijEeOH8a
3a9vKF1pUlFQo4M6ytp+XN8vaj6w4laelonAltkalJ3QRyp6+fJpw/hH+N5N
1M4i+12Ew5DiEXIBHcFSB3pnsKKeqdKsQ1CIaGg2KyXkiAi6RuBxd5bNxvLb
6/Ys+C0dMJKKuFzJ6WrNF3GRD3gcrsBhHVNvbwBpQ02ecJBKqOMMxgDxvyhR
EtyUu9weuYVNFzzkkL91SvukTIx3r5MI73vP/2SWwcuQb6wY9O6Orl264sIS
D43BHch5Nmw2ukWejxH2vwFdiVWFYT6dVozFh5hHvW73z7VM4q4yOUQjhFTo
i1r+3tgw/+Cmfj9R2NWuMhYVGivk0rQB5C99wAvET76I8BR0vN34A4buzJuR
H/jc8pUotp7s7HVYONwZvMNqBJcfqDXHhdONeMUzEVWdjnazjldn1u3vhn9M
ZDV7Cm4uqqywvC80LgO6T9m4uDZtn25quHaFZmQw9bKeiePYiTA1+mzZphon
vJrFLv22c04/HeEKhUHHqqfK3G6dycfyZviV4uzmWvr3a1VwXI1zzGxWbcs+
hi6c3eVHz5OBOo6Jc1dGavFqPCMUYhYiNMGC9smoa8cPgBcBvneDol8T76Zx
+4Wb8z5UuKDifs9N/8HrCN/ZKzUSs9u9HPehRHIz06Ww2SkZNKioR3EJ/XRI
L021mUFNSnSoDcuGh7I5iaJ0HsKqrkAkOKQcSKgmhsL2P+KkpAwChjVulhem
aL/DxCYtqu4e/Wx4b6F+vkH7oSIDwFIKYknCo1lfJQxEAn8CdZ1AL1zxR0Ts
98bf8FUtdOD6QJFJmQoC2vHQ2G8dhqkKvn/XIWG4VGXncf99xzwsiInMBr9s
2VeY24t0u4rqtOslVPrrM9M60M7USMqHN3ESmMQAdIuLWWh6d38/8fOtbjCc
0yMlUxscGeBv/Ysamdj9ve9YIMuLXKxH+jsddXaE9qQSAvBRyEkB90FojTeM
2oxaV4gXHcFLlc7bZI9Url9wQVxR5YJcchICULhlG2WJWw08s5quUr3m5mnc
3QfmdMpp+vMGUyLoxo2LaWwjcw/WQwXZsurj6MJJG5jXEYBiKtAlorBR0ldZ
OwANXeSUqoUa3yER/bpNe8UEoAZW9R6iawLw9JXSu183BlN9t0vPUOgn7HwA
GBf3lFlRk+sFfjOoWs2etkdbYF6A4zsO3KigfrTteJOIx0BQTbQrvQSvUz7H
F4QZXxHlUnLLa/rhbeXvN6p2++Z02nOtUy91pKVB5hIGRpCy6UoBr79RnjxR
SsHVwnRfy/FoQ3yAmaEGHrEDevNjBWtW4f/j+9LmD24cPsJDq0p3nnEHjnt+
ecxmnD/0hNHtz3dQtgA9i10wfimzAL+1QhkSN3/lvvLjiQ95vmaTJqnK98sr
8/rl+bGgupEoPJEYITD6iR063DHUs7j0jNAhuaFhDbYdRlVMfsFLyl+liWpK
gK5vacrAQn8Fqm09FldanFKI5OT05fjhqNXiqlR/xdM7BK9HE3oQmoIH5Xpk
xb34Ps8rWEtIGWtUfpJ3Q6H4FwrtuqFmbB8pwjY6eue2HsEw2WG+s/lErfIH
wMB6Om/uRV+U2ygVW7tfgn1LwD470OLRDRf0laNDdEvlrtJF+KPTRGRkujKW
8eRwMlhtyy4h6XSU2Mng//1N3Ek9YKKNJL7PIGr4/FaO9M129Wk96+aV1sci
DefAQzD2ZTdasPQp3qsCkhVUO7RzKjdeHb3uTpACLJ0yfAFVQWB322xcqRPW
TY4odeL/lNRPn7KNi82O6IXBwHMUhMyfbCnaPdRdTsgTKJtLcfWmtW8z2+L7
vhFGYghVpYi00EXLYkQb7jMpMoI42MgPlc0JvUoiO28H360HmLaGcQizuVa+
1w3sDoWS970TH06QmKUGTlR0VeUTN2QOuKAoDlkpxb3Mfns9V9khLeQhlFtu
UiGmswZyzaYLutGv6cJzjdx6PsLM/uzBHv9m0Ywq/+F+2sVX7aiUmUgcUNFl
hlA5F5RiwAsdYaol2BLikGzALeFdgUbaJzx0Bj7Bo7fS7RcFTDCxhzlJ27aF
mfQJW+0d+vnbI6YRrRjnVE4N34wDuGnfKKNlr+3AvpwOa7aRZN54YfEeXVLR
+/R8purfVGnLUoYDlfa27kN3+velCguE/antPaR23hZd4ePzJnnhl2LOx9+h
hpta17UsZDgDBRsaIUiajz5mjhz1BKsKibQVxVpPT1K8ZSUGXGfLx3ZpDfiu
rskluW3m1GhP1DAojAmQMFkAhJNCh+ySyU2hImCdP71n207+iTQ+o4ivf/3O
AeJM+xCriJ4H8ONDaAGAKjaY7qTVpQe3tjDTuGPnbSQl/VPRfsJQbhXv/JM+
ApVQexlmuN0ygIMTjHZjzJY1F/O4Xe9oH3S9aQi7lM/DYL0U4WaLsJoLWVyO
KKspPT6z/6Gql/MbUf5hItZe4Z2trs29ejiyKhKzcupAAkiwOWKrteRe05o6
y1pKw6C/loHjZSjhl/94yq8MwZ0zhT5D8jIh1PFYeFt6iun5+4/jSxHZqX9z
K7xKNhd0zHWky1IFfaxzb6+aeZYx1yEAyHkxguhh+LqwX7g7EVA+dPew5NSs
MKltYxE9mk41AMnVaPQdMvwed/rda6yFgmXYvPsJMC/miL6WdYlL6w+t7q//
kB7UrtuEwt4g3AqU4X1W+Cf+eM31cK7L1E7n5AYjhFv70cowF2kTBoMEa2jw
PHjAtSHzXAiIgmcr2gXRF+s3TReMYq0P81lXiXzcRLvG4swHBLSbMaeN5vTW
BwZP48r5U+O4bsx6+hnOxnQfo6udN3J8H1fjRpZ27WjZqzTcSJn5eUpwMGXM
SVp1VCXzasxGL14/tvomYTACgny2E+0hi3r6mgCbgsxV/WH3Y7q0pAAlEhql
608Wbel22YoqW10uQQKj1Y/PrWvkLfM88AWoxl3vgQfCbaDCR1Du7kJT7S8L
/iMc+XqjlBcaqy6IMs4ExQsr4ArTyMDF0U7mBqlRY7wIwziutUJb039NM8L0
YomKJ7F1aAR+PfcZBVNw9rxIb1NjrsvC5tqCis1skv5wx4Lui3GyquyUtFzA
F86LJO1ojsU7XsC4p/crj4SXWckiVPBhaW9eq18xFCU6uzN3/1GCNLI0Mhv7
C+HoRtMy9dKORpsF+1qW9XGPSZTNskWnOJyy+tPkZ5hj8fz+0U21Kzew7LMM
uNs9EvF77WiZYF1z44nI/XbRqA15AafUq1PXP9UaNODqWfpyypYVGeUVqihx
9mRPWSL9AyhCBBFHaA4PRr6dEbyWf2e6bjd0t4s2rPrQ1cXYJkKM/6thOdtc
anQulogpNkx66/m+cPiG63utQlWS0SouLAXGA7IXBVqizi+GKQdxr3WXSaoH
z2eHIDg73J87BZyBwhymUqXhA8gw7CyG+O1LrJb84Ui59nQJ3mz4hObyIh2k
kx39eiGtaDszSThXqf3U3A3erkB/0qOVVG7rOs5VxbUzyO4M/n4/V0ibZV8z
ZofBSkD9ENfV4aaRb6IWNWKT4xKXRdBYZ3OkIRhY2JKNTUwN9vRafcIpPgXf
9Jipb0yF0edMsRD0y8esAWAHrmThdcm9AP8Mg7mrVwM1ZrwBZY5x8kl0/QjW
RH8S+W09nlbJ+8CVkeebp4HSH8Bi5tjtj+gOlKbB4GN4A/8LjMOIAQcAhqAo
u6Fzzj8vBoVoLTUPa3EhjeoWZh5zNjC1TJ/KLzs78hkriCbz1BDsEnoX+CS2
IKlSydfB3DTs2MxvAMGVPoF2hWY8RI6cquIOIfLWCLZf6gjnOSU7worxcNus
g+Ncr3Oyd0bDsz4cbXWnb7R6w/UMxMtKR6h9ib23naqF42Peg8sU3j9c6ekV
48h+Os6IB1a6iUdRp+Ep69yEEP4A4jDxZQX4m1q0Ksk36VDeKZk3zC6T/bF+
C2z7684Q+NqWUJfCIgDYriYwCKX9x72dpmUhMOm0ApYEsTEnWSgqLoKDbLmi
iWhS/XHvdEjwH+HCxf7UMl9Cu1SRvhrQfGt1J5poNDrdbeAhci1qbBKNgVcm
NsEuGJchvCIyVjAUEAd2xjx0jTXnYEZ/G86KRciNz6qXvR6TH9GDTLF0VoN3
06srGLiOBBC7P6AAU7d+GFsZmsX8zjXvtz5gozBe0stdcME+lNtWAHoaKuIC
Go2HcV3Bcu/Etqysnp23x/89DwaQ92pE/XeVE/DK53qptjKwmfxJIUNcEi0i
wsTVk464SCY/3mipOBelFD2l//zaYBWkb/30wEWRMhfGoT3kxc9Ld+uXhdFj
/cmUxjcDOhAQmbF4afgI3o9k+2Bk53nTlCsVeR6C5ItAHBauvWoQo7KKOjdk
lwXwYh0yxwptabYNlj2GzP9tZIWSIReMx3yp1nFqDFtpggKwxJIGWlvmwERc
DQgI5CznsqHj0FHP3ac3H3JRLb5PK3hF6sRmwSx2yLqJwjVo3AsNzev9E1+s
yLi+uy3N4dA6LqqKtdCLgqElTJ9Fb8BbpDmkw05QZUqT//erOkYrBBCq9BP+
gKvnLE2Bl5rf9aw5iG20wPh679W6wrT9YrtQBlXt4bYUC9P+0JHRiaLNk/Uv
o79VgUYeYc3PApOUn6ikGyHpYUB4MA1MdQn69BVPNr/dMsgrlQdCSss6+ehV
9DIMKKASCBdnGyJIS+wBSpOlIbZbCyFdkbTciVmi6l6OomAS70VfALc/S5Wi
rx/feE2V78fXUEhHZFc8QiTsKTgnbJ54VpBc5lxNKizwFDcjQarXNtzZIKXk
0ojus8RU5CDC0DpvXUBawEDnsbArHRcAW+c5GK9jDVGtBNTM0wt0wfExAttT
J9ozBDzU+tZrkPDguqvpXhrkNZBgMoue/h4nJAcGF/fHQDIkyAzZoA4AWXlS
tzY8iZgWvm7ax8RKo/nVG35a2DOYKZtgSAeIb2NsRqtmzWFQY68n/8Y7898s
Z6LqkvOpqGSe7IqbEykKrLeU7j0WDXYu7ZqpijuemHQimvWtBRtyhFU1Om0w
FrBw6nSECIWOgVMljIxIsoxBMa4oWzJm85S1yCE6ZTUwc/faNqGySiG1qAn1
DFVn/40P4oO/51AWt/zJr0auFhKIlg9Kva92Mf3um37AKH4xYMsB5eGIpdkM
yAUmP7dW2jDqFTS98KMTuC0ledVeYT92NM6kc6rG0t+DmYMj64Xtq8XV8eVZ
toETWEozt3pK/bNj6R3CwW60nNPdFjZPPKtLqNS8tBnlnDBDPzMGuXdWruul
tnRSRj2wUFAZBE3JyMCiFb56vu54JmsK65qU6G85AOMcf37AKW6gAlyPj5F0
7KNZ70b2WGyMaBpSpO86nu5bofEnlJJqLHT/fGgsLGeFbn7G5HUfDGJxEp6i
9VYAwAUThtH2uYh5aadnanz+LoK81N6zkbZ+Wewy1ZV4s7RpfafqJbdGex1p
Df02GVGsxonJw94/yhmTzjLpEJ/ozZO9X0U0OccnpyLIDlgBH+XbSiliMh9J
eqcVQGl9P+yxLrvTT97E/ZO0cWFO17SQkQrWKhl+UEZP/kqwbzHu8kFwD2b0
E+KfHnQfJ2MpGRW9WR/GHnKBot4rDKfv1IBg0NaYg7j46swQNxu/eS8sB1m8
agT+ySUIAQ9CZQUPL3YRSL9j1Ui1ZVVBYV78xPzYtTfqIsGCHx6miCXIvFg8
SVV/zTc6WVI78cxCSnAmd+c/eC9UVfsZFamoXovbz+M5FPI/XsrpxSYyShIT
bJudTXBwOzJgTaK1z8qBJONdCZTvtsgbb8zJyIGLk/dmvFriuRpEeUKe7JOU
XPkjhxzVEPn2KVQIS6xkWZ5k2BFgqCCr1EP8IcdnAPRn9S//n7spslh+/s1g
1fF6K3HvdiRcPSqU2k5i7ZCJXN9aKY1Kg0Yhvj5aYrw6u2n3yn/Dq/XkTwmG
hFHxCkwFaycVnB+fB6s6dDZnPesSTHY22H4XxhIzpuxUEZG3zlom7qEtCUNe
hRc6ZfGIIXv0YjdxU3sZkWGe9ALP6um1xmwcI63lvU4EzAs39IAj1IFCPuZl
UWDMAL1pZ65RH2DxPYz0OLahIWcGzrmcq4XLhBczOmYIZqiGJXXsoCIQfvB4
mIDYC7ZvNd+xXWCEkOFA0gZkk8J/8VyDpmkVxLLl7SPkz1hqoka8epVzfXM7
J8Q5fbwzdnkN3s69qsyxwOBMtJ7yGFWS+Nw94v32GmARWtS4MQNA8yAJWkBg
Z1PSzDZyYmK2oBFD9o0mk3d2MfRyO5yeFp71ar3LZqOfc8QBoRtFfrLmm6D/
HHbMt1k+NTzZvdPS5DHEr7OhBco9dCZ/f2IQ32fZ6pHM/RYxKTjLjvVnooFB
3LV5t6tNmxIE4wwnQFKqfr0pGl1BrJP6/3TH/KFxEi5i1vsTZyFkz76gxLon
atm97Ht66uEKqBXfqN9qMxO9eT4X0zOynSd/XpqniD3MZOYuKLD6TwuxMwsw
oSlb4aEdfoAEyvRpcssKwp+51ECyGSupDaWAe4zYNAPBgWX9HqBGF+xQiPt/
tkMZi0GUUmXnctluk00eUs0a5ovjtbdE1MKDWFbHhgacnX4alWJnFdNmMPO9
xxg4zATT5TfxHoxTy59BUyrDy8KFkOMtaN9SX83WVsByQRqkmb3V3eefzPKI
UfR9qsKA8aUTWLyHhbZrgbRB/px/5pL+EJe8sy5dRunAJVmMd/M4ChKFdOU8
sdfh34gb4TpfadFSVFuFTj6KAii5n272p9tPZF1YZKm2KSH3kAAW0/CPXIn8
Xhv5oje9UWzsdwFGj4Xva37gIej7hIcdxgUhi6o/8DmhWgubOEPcljkLjYVW
nspaX6gbGRHzksLF5PXCiA7lJ1pCtNpJdSkOfWWXhpoGaciO0GGEJQInJghJ
9vKX7wRHAp1N2TR5vmOO+3rdrOD0n9Y3+sYpFZA+M4L7u8nLKDThbkYa1P47
+vQLDgDDX3Tc6H+4t3nW9kht6/R/TDlAW3L1Z38crxLqCEPRuQlsdbWb32KK
IgayUFBNToMyqMOByyrosB/PhqzvugiT5Bsqqfnm7pOBCL7X0bIfwdrOsc3X
VklgevjUJkwchHrfBZPDEtZJUpYcsD0ajmyPNg0Aqt08Ytdb0+JamlJMFL0y
Zvf1HCpVPQPxzUAPAGCXFzFyzIDuunfs/kN9ZZ093x6JMzxj8t5GtEgublOW
oyFCGkh1eoJ/HScfRCWmoCsz3NiJLnuNsT33CX4oloRgAzJoZQOBtUAhGb0h
N51VcZTS8slwaTR9fANY5xhVqVxA79iqE+RtBA5Zw9XTOyc0MB+qv/UR5Jr6
1T2bKypseeWYnXDKCx6e3YQ7KekPLbk42D0jas43hDEKmmGwHPtErQYeKFeP
dmER6dlWobKBo9MmIfwSFTZ9e72EPiUrwR7YEdt3HjJNrRLKqyemZm15jX+A
Vj5xIKZ/j4PoAWwbZVHIkovwbkHwvzIx9KclBlkK6LWae4AceNNa7cdTqvGk
Dyla380JUcWiD+QGwAT2p6EfVROkRCzLii5f6+DrSxdm+NdJG9z/HrPbfXHh
GW2upYS3uCMAK+VoING2tteNye3ukdSgSfxcP18rwoSLZO5+ttJyl37KixAX
yHsdXazSWUZKE4BOoEPRiY/U4GMH1S21eegOhstnzBf5Tkw51IHdembLugys
1gQx4+llb3Ybb3Neoyh9O/T9dATKrL5vHJAAaGac8tAWNseJKLdqUPAtKSes
dZdSSMz7Dn+pRhDSk4GC7/aC+up4ILUmirjv+b7ulW68mVXTUYzeyhA0hGlX
JlAG+ai+2BRwaLFFjOAXlyKVsjJVBlEKwHOxNoQpyoxSAUMZ9X9H7i8QX1pk
Jq7ICk2gWxqgB/mFpDsO3rbTIeMu4Meqsxnodg/Mv2zZLegyDEU6mHC3VWBh
ZnzxDUbTvoQQsxWLwaUTuKCyGwfgbGmMpKGQpJexrnLKxzaohssM8curew6w
QtNqBcK7qK3aAfSjOtlcHlPAmC3zR/y5rGcvfuF9qIAjY6rZWcXZeQIm1+n3
1e4VLZdmYngno/Wys8qguj9mtSYUMqMjzzYpnsq7z1iIxbKz41FG46R7CIwh
BUPS+kb2BWSvSNlpXtnWmeLnTFsXlPK6v3Mf39mrr2nQ9MAsHJqfshGU7mst
JxF01xX1FHDFqZYkfPoThHoRebS5EyYle9nvxQVcsyVFDJxu85/fmDq/UIuz
4LvR3nzlDhQnr2cxhQPlCPDC3AA+Ezz99GXPiXgJBjvHOMH/H4Ja3kwY4uOd
pFQzSc91eUL+37eFXULTi4LvOiZkRbPDcz107wvFPq/sQwkYB64Dc/FCvnbr
AYCfComQgolPI0SRzBpq8cvfAB5LfO0zcvU+ctMsB97NeKbxitoWxvoh0GGs
xKSq998NIQciA7IhjLYk2JIe1xF/ZCATrmUv2kWxGxMOJSfh5wc4p7Nm0vDu
1dWHDP+p1dpro3qCXMpJv5SkBB2Aix+k72o3hzdOZet/chqysgHHvrdP0ryo
bcxNx4QZHuadZPggN1XcIPmP7DPi5qITwsHyQp4cK1Z+zUoOBZvfNKDNDmRC
oasVAOrnrXhq3PXnREkr5ILxZBzNbNPcBtKSe/hX37LQhGkCzzswIh06V+Q6
3NrW8YzwcEKGeFTB8Fz6Qo3g5qfy8ZpEowheDqB5RXDZmwcnm2Vsh2lLJDqi
11EC9Ou2l4JPBM2MK/a9ak+f+/ZsYOsTajrif7q4WBYMT2C4GIs/u24uVGQN
VmXlPziCkGAAlz6MueNs3jUggxMhD/mZg4A1VW/nCenTe34KtulOSG027NtY
8r2W8t2V141D/LTqT1Wo2UY5KoFuZiO5Ma0vNOYSCAvfRJRjDm9hkoGTwd2t
w7x2luOOCIX7vAz1fi8cNBCkLuUw658gGBWBvrunwV2moXKSzCUfubCjRhXW
3StEpm9irhqAEzgO6iGoTyUl+fOUBozK9Gpks5y/SWupnr/OOh9iz2/0Irs4
u8zTbKk9T1Pq+Q3dIfX6o+evkUOyXvd+97PzGeFwBTSW3uynT1nkv8l+jl8z
mbGcd2SjzO83bRz9tFY5ZZDcCHMgpf4ZeCenPq8GQdbSogMc5ebJnYL4eXMI
FXy4/15XBXaVIP4nmTI0bQdmWtlgVhxgXcoSHwk/qK94JqjB0R5JX1Q06hA0
4RF57tD4LcOD1NHbKmFDxxpZB6SjkwlKyN38qSwCU/ByA5Pwek42G+EmwWo6
GaYk5pXmSJcK+fJWEhXX/gdcjRCUO8u80EWr1Ld6LOwMvKCS+kHffPgou2AA
+AomOt9bi1Cq/0OtEUgurqkwSRjq86nkKEwQE6wGe9HyVAH8+4PY7ToBFYU8
/S5aHVn81Zc/TJf5U4MZQoCxugXd9ofbWPTUiKpWRUiZX+wymDENC3M+FU9x
ij5rI33XJfpBzwunb9P0FOKvfmhBmafE2ruspB4ZHHU+U0ytwfwnjOTNM96P
gNJnRpJtnBR4rCkGsyHUacVwLbltMs6dn9PfnTN1ZW7aLRmLGW4jiSuWN+lT
hGhilLa2vXIgNmaoN6VE6tpdBhHy8uFSTQuIEb4Qh+rCyWEO6bPjGzuzerUm
05uqoFMFqWQodCeUYFRKu2I7i/nd2/qsWgxNLSuQT0p5rQdHxv8Upz/tjaGq
NY03u+H/LPhQIFeuSPsDUw1r+Z7Osy6Btvpen954zsWqkN8sDkuAw3/pXl1S
bmcWih7PdEtJE/T8NRbnieMa1buoEAV+C5c75o58JfDhcs2YbRfZMmDYzZEv
57wgXP6cOlm4f19/Kip8vxV2uAglMxP3b6MmFNj0s9OdnLt01zLI6j7tvEWZ
upnFXnzs9Vky/jUjGxzbObdyRZWhMYkx5cyN1wmBKfhnXld5rqD7spkpJCtQ
JPoEQ7EYL8ipOr1x9vwGRrGH9n4NdGFgepAPXkkLP3VWCiNGfJGKfOtOTscn
Xq3qoy1e57ts47jWkRfRMcZY3WfYNGkNI3aktlc8uWZzo89w/wvHIPFhBFiZ
qU2nfHBtUa0hB7HovrQJrmQ016Cvvuis9p+WgojDMFo4z67dgvhAZYkhJ6RF
c4N7cbFYVUISdGGfXBWLthBKH/po8EMDI3FjExi/WGvZHKZqgfLwVdn2GRcy
dnqs3+pDkPf9QzEaSFbbnMJOsMXgniZssNrt5qqSclQ+PmAPIl6xnrvDOV3R
Em5VNjZumwhuxSdQS/YGEVZsM96bTGCfUcncYvAqmaxmd7jcWnevUUgDJQzl
kyGcTlDbr8gIDihzg0UWOtV+tCS/HT+izQ/TaGFksLCtHnvIvVAYijtLDl7/
jbtxUQr7tD+9Fetc/jdpAUdDuFCJEfzXTx7lIkyAMqMO29CirS/9s/agoCYB
nIvV7u5lWNew2MAs491x3puMUB1juJwC7C1Wph1zsmHa50oBlQLxmog943zG
SVUM77xOe/+1m7Wa7t43hs5onvOqc0WG4kupJAELYaWPaiJqlMBwQIR1nADr
BPaEjkWOGTubxl8IIhHp920SOmIdYF+ZfaoGcJMKja0RzLSS3w1+opS2fSUy
+XyK8JpnhIHO7aHfH2cUdQAPqB5jpAt8D8UCntwK/sdkH+3A7y1NXonS3CPC
CqWI5DSJzOaDagW8/jmCagVy8k+PBgI4r9yDHSfXuQvsbAi6+sbzNJui1tKY
MdU+bCZmclI3LzFpFjtNbmE4ZO3NMHFAYhHfa61WbgQjSRe2Oj+erYfAtZI2
A5szyCJkLDV3cwPELKfbI5zmuI4XcVNhHBfkYXDz5BeV5Z/c6KqqB3gVDiYy
nu3X6znpJ4CSMer6pHahRmjwzzjqRPN8yKyDpwVqS5EXLkDLTnYB41es1rFA
epYWfHcYoTuRm6x2qsaO8sgPg84YMJJjwVl8jLK4g1g5X1/6zonXcKMOeCYY
/HBZKasigHxLwkys11uOpoRA6Z925GYdsrt4PBIPX95ZDOPjRWweVEqdYNAf
sy/w2yekRdDInqWr4dezFrknZqM2MorILTHUWJBWihFZmbkt0xmI2BOJ24pg
/go53Qn1ssPYHe4tA0FZQW9confDG2rwiI6nO9KZM34sEaVvRH7iTlmt0Sz/
b3sANVHD7jlznZYy6p/khNqCtpWeI9D5PINQKXWxYKHRk0qkp5YAjcz7lkET
iXhUib6mj5a3/F5zPgdlson5KlH/Dq2/YHfs5p7Oqz9qJjhEHlz1mKxG8OQk
gmE5IvQkWfAmc9LSXWGolm/uojQQqbWGTsTOV2okkHiPMf1B3GPMw90S9Z2E
M8JtD9nV+5lGTGgxg2RvWobOd39LXc/SS0jElh5YRhBkLbbtsiLiTA/X3vji
aT8V54xh99AXc56qYnAk57uloeWZUUYFqaCZJIosD05e+6iofE/LW51tuJ9M
kh98Py6+nbD8/yA94Ly7LAJbcYtqZffYJVQEJKp7KjFFwxeO0KaV8VQ6hXoB
+XrRH48Kpf6UeoPBWczC86GFVnjv0uQciWTiPzQVIuefLgGb3P3r/73M2PIi
zFBbmCtWEg7diZtUfb13XXewhWN+dALtGDAHEg8+nw1HpWeQK4OZfKk7sec4
PvyK78X3kqix6PDg1p4s1auSZk0EZlsS2NdzDraEjgpakfTT4uMLnjdKioNH
pONc1e+WgWDZ3pxhEgwZ11XVEjhd+U7GZLF2U2KRzEwYD4zDIgDUmK9zUliP
bn1obW6y7kAmNmRqbPO7mKUdECNunwa1OZlTPaB1K7LXGQx7XbgciiMWHrDz
nAKRFIUws/FW+RP/zYqvRS7zbeRhqnvXTjHvDcuN4cI3VlMtVoDa/7+G8WQ8
cHd4Pw75j2lUR2dsXpT7BiMM6zvii9j0zbMNzH26eMWY0LXdthwGp92yLgUb
6TazJ9ktiA6UGVqmCLKHk4xT7IWoqJH5vRUNKReAN6H4OgwkSrZKLhlQWSE/
VIlT59dufPUvA2HRABe94YJnQxs48ieTbxmzwEcSAwqSdi/z5u/M+GyODgp4
2GNuAZA1FzfsjDSmvNPnvVLO1h0Sl/SijwKg6NzwNZuCmtDRv0ilH0lBMBjT
AWLPsl5DqWF4YJvrv8W79GC5ttAMOHvFA6xkjqKDn3CI3GRhLYRrsD752rAL
L7lrV2nV2O3tEmUp9KJt9uTJdC2T1tDN8xYu65of/1koPf/a+U9pDQIlCGoi
dZ0NkJFAGE0dO75WZaG52M5HvG+g9dT6uTCuYY0llLVyC96uITjqTzk9ANrV
9xpQ09ZT6SZJugAwpDOhWx+NeLoS92jmwfUXhigXfpdiSZhIx/ccMeqd2Xlx
UM7bR4WkcWy5zM283Py/tbnzXyRchgTXERTUa5Yj5YV2yq0iqaXlANz09wNh
rthgE5NX7poHH+EjD44nFJkDj7I/iYQukO1J/bO3jHdJdiATIgaCwory75U4
oaG1oH4F9F5Yu9aoF8eFsJI9Co92/9G525HWBscLVlLYQAo85M+VtpEXtNBe
rRONLmCpWZhSZbML58S7CKczvWN4gZJ7M1eZA8si1GKl+g1/YXzsCExksqn8
elifyTHrfV/5UVKo1fTvp76jFWGnjlpFTut5kGUMeDtGSjLBUPF17Pz+Irqj
n0McsI5JrVh0iJbCAebdtMKNht+lEGOjEqaNARfoRkrXbmhT1WF9kASw7zw6
zm6pg2s7eCIxp2abH5Wm1xGV6tE+hMwhuvjJVqprSCEOXaNTD5+P1mqFj0W0
8Uxf0VLsQ7ItNSnyLP5RGCDCE4ttESv7NFeDx3eALmxel8pvdd5kj7pXyvjv
KvCU7Vel27A8WV7wpLao6YyHWTLX3qZNBFJB7fm9iKoqJA7Jjjfx6K9+sz1Y
+uXHSwKMtWIvo2bjYkXCUg89jWMdNvzHvypQYmPhr28IXcI5mGCvmGRUCkIY
NXaiDdI6SxaX6ZG9pup9PUK4SjH5ZFFe2doY2JgSRCzdzdmlbjLMwl3+MHXv
7bHBGLYhMJQdMY2UWOmzzzuObrsEL8M3LzAQ/s+RigRkhlfCya8/y2TiT8uS
f9pmeLFbRf3RM0DTIER7dcLdVDflU0klh6w7oy9YEuyXcGn4U3RXAaAOWdYh
v0sOJ5AVkNPuWRIL82tsUr5V9Mp9apFAEbgrDGVBPc7aBRoAIzH//1Arv/RD
xEN1H/jezBMt5SrccFMK19w0dTuEHoUSq3BNerBpg+jBVj0lTRJitNWFLtTz
vKAR4pVx+akigYthIb3W/J3147PAsgm2LvqrH/cKUeRPidzm9e34rqxVk3wq
5nkpMjDd3zhUwPqemdXoj1F4wHklvZrN1iVgSAiFFIHcUyXXiJzvQ82R20Ds
fd1iMs59sMQPKzmoYS2L2OqJUMMD5OX190hzuH045NFsf+T95QsbXejw3s3Z
h9YikUNBOAzXY26iTBYC0I/SKR9nqWwxFVzwWKmdl57YLfkWlTgBqdH2xVHt
4PtbmR508Y9oMglfa0xkOYN9jl1AmD01Xd0aImNOV50zLVBbX34XfZfIvYtS
pGHcehHMJAtJN8gLosWrF3LRc79wqfGrFEzR68gU9DqGBcw9s1oeHxEsHVdC
5vs0RLDr/Pe9zCrSsotpKYwHJUA68qTWWLBz5tyE+pkbpCtyxJNfK0quubRd
cx2amXDCGHnSRWOdTS2hyHFlEhwLMeD6sBipLzPStvuSKOKDdniI0Um6IMFu
gUE3y40FF8HW7lN7TpklA8UQxtpEXL1gNL73t/IRocoRF13pvo4Ny89EUx2x
Fyn9NtDuYhowKGBHdHfGDO0+7C3zuJ4nEmHh4/jgkjoYAtp3OKBG3D1fb+D8
emUEGfK31D/BcQCBO9kQwsqeRc7W+85XCexCasY8gUvQqyzZKRwZnP78l6BZ
juy94ilVbAdTYZK46Bn2jlf2n2CCbDC4me98NmH+aXI0BT837/XK/yXMRp0z
5Fl3IOKcXRDezyTYRtRI/7FWHBE0F5wMcSZmssC4oFinCL+1545cWysoUtEM
yIJhBK7Xur2fEbE1KhW6yenYXhinf0YgQXH2t1poSKdxVJWYPcg5duJCl9pW
789U1jD5wL9zzMZS6ZB8Ki+8F476QF6VHJA+gsWM5OD5YjxOIZrnh1gGz2kO
oIcxLVCsD2WMb4Ze5gpZNJaLGNm+d99Pd2UbBW2Il7zfGN6k6fT+GhjoeY0F
F6VFTEc7qK2uM+A5P8tYzneLI3V/t2M3K2KWfCNWNImAD0knVhgNUI2s100o
FlN6jOBqs2q63ESWZJJJkDcNMx1waNMgcGxtunX3GV869ZhQjHZv3XdX+NFy
b80Cs8JdV24SHhTUafpWUmEkEnjxd8te02M8tt7x+WjrooI/QrIV4zIS1sJ8
n7fbqXJiJuhjznoATeUMB8NgZnqYSRrtd0XwQPL+QaLSssz+pT8TZmu/ae3k
ZQgCNfiUy+MiGJA5USyhqRR1PWXlLQBDS4LOffiQrxhprePtAk8/1IgyIrJu
Iq3pEOhu/voE3O4/ZTfG1Kzt6phONYGTVEiaQ8YvPNlRY7x6/BfDiaAY6iUv
BzrjnMHA2s3NxRX4zETJAkQGNMugb0H0sgyRFLE/s4CVswHMZln8Ldb+EJaj
AfjY0ogmjkkELaTIztSl6r8CV6hz/2q5KT5hXV4jIE/rmc4Ux69gNuLVzuNh
2JT248IofCrkbBSOqMLUy6pDILxlfwZYXH8DPJ3/lM7nXF2gN2BfL1CMRg1g
vloIQsagQ18xMwVovO4japmnCEPqvfUeEFrl0Dh6SoU8kcFWKEE7lM8HWiob
rgsTRJnO23mWcxvf6uiaUif7oy4LcAJis9rrclFgKm296Cf+AfbjfgA4OBi+
+KenuDOdHrKPxfQjgig0GpDBXKrmyAw89e2gWmA9c/OYe9rgQA5tTsbQXEc8
ivbmgPLo7n1wRWKcIdXCSkBuIdWzTkGNB1jfhalruN9YkZX1/ER4DcFJV7fk
JZg+zBqeBunsOJJfBQ+JNugmZ3yW8bxP+U4GhRWl1m3kiRdfrgPKsBvyShSx
1Z4Wqs403fxjufz09m3Lp/nq0z/EEqS4LebNxdzUDoW3Icpx3S2cv0AJnOOB
gycDqSnrVCpzj3pIa/9z2Q5AGZziUmZF1f2x7az+P6yHz2V1U2sAcPdB5Gxd
D1tpW9a50EtCkhXr9U4ysT1n4fOQpZy9NKsG0umIM3zgahiSmqM5AWUR/1Jk
FaqmWpjZaHimOzr38l1YCOUHDEHwjFEnlBhqtIxWlHkx8DZyJD8W5mJcoR8w
qD+FVohoV+CBujV7+aBkAsK5MJ0cTPoTAqCuCxvfxTvhccQ+5ap+3eLy8M/1
y4qpziXk3oGtBjHvdcOwTKRv32PFHXaSSdbMtmwNcGJr7GTlRkCP+/CrevMM
p/5FzHRVOo3j91SQA8h362s0lPthTXlCqEzo9NJ2LVy56Qyidq2nV/4sg2AJ
gDl4ZgGe7BZeAXpUKb1o8vm19R0sBjZ5CSDNeInS33e82swbF72YXxIV4BYk
A1uleNzPnj11GRUe25/D5UdzCL/BybKIGE+X1bitdooSdHnPAaIeUa+65n2x
SBHmhqkmCb60GvSz3nb0NoLToo/MnI3eWDGgitti5FbOhVqJk4JbmhHX19R2
dgmGUiVxc5Mp7579NXNQ1z4nMCDASjscPSOczX6RH5pWd3FSHBr3jtRNgoWT
S7XkBRP5t/z9y/eQlHh3dmfj2R+uRFRe7yPM2DqtUh58XuqYQc6LyAb2MJpZ
iPCnOV0X5u2g9YiuYkLE8+JdvNG1i/NElA3V7nr/RLqBpPPUhko7WVBZjJaB
3OHkwbn2kFFw7+dagnVEsDuY8fJ7AY+9aIRrl6XMXvTh6gMeKs9vKrwsv3TV
agAzJtbGrRSZecjLhXsmbLef9H1vNboUSIR2FJ0uY5jNgDG81kSZcwfyrmzB
EmK4OsX7mhOQK3nojFIJQ7kWh8RaTc1zIhYzASLb6eiqMLTWXvldERMwR5jr
eh/UcmxYX7gM1ztTzsC//5RT6fX4aaUK8FMNSDYbxXLl6bRlt3PMvCDQEm9q
CX1rLHZ0MMDyGPffgxf8TLlrK7NsKtr8zHIFMsViSiTQkKHoUCo1J9w63lyq
7mKUSZVT8hKpWHZVhNZhpAkgI63mGDagcIPR5hV7hurIXSsmTswdHk7h9118
9y8nOSMepOfUvli1eMr8y7juvc/Ye6+hDUwsvSZNpKcIPMgHrIv24OCxYQvf
horsLq/alBMS5/4yENEGiiqxYYylyPSetihGnrJdakOjlX432JrJA+MDb94V
F8kP00M5bGuHdYMO1jTYvMwfHJXanAZ1WX4cDq7u5t+QL9bsBrPteptoluQ/
zWJEfWIVVd1w49nlMfi1eVx4mwC8DawUBhBSwTLx1FlxwYn09UNVK6366VI7
SpxyVTFo4KW5gudDa1+FfBM+AM3Jfj/sEpa74R51KwiTnhmC1zUd56XwITBu
r24/zqNLjWfgJq6gf9kVQdHGGhHzXYNVabN8ly6xwZxDiHO+ga3r/Sj2daol
/WQPrDTQCSACmZok0OYalFq1Ui10LvOgKNSOYUqBYtLK+9PNf4CAA/tShaCw
0f1hah3Xjn+GneWGglTo5Dm4SPYtcWv4+eM0jVGOa2Akg3L3vzgTJq5oW7fK
uupinFczPdJxU9UheJ6X51iVz7xyZ0kA4VqgHjNagUSrknxtnWJ5OifYACUa
tWGM1nHTlui1Oz9rl1YmUXkBPRzbClNmBB8mRiBSJITtqXzukSW80TV6VWoL
v5vIMofmMiSx67a5zGY6dQyWsIIpJq828NY5CPuE6M3cLzqdSKkFDWtfmIVL
dxgmIDcTYIkZeQIJQkBygj0r0e81iLDCoopSC7hIrfKKhnC7/jZRD7Dp9MTI
iyBFcw3yQHoUuADQJVAyo4UeZUEp7YK/aPJHpSQpfENInWmE0JSk6WC3WBPZ
KLd2kc3Ltz3hw1E1WKXF51eSE+y/LjSmVa1cNT+Mb8bGT50PIm4+IW9gQfkL
CUO/1/FP/F8LiPk6tuiwvFmeb670ysJ6rt9VYWjqk7aV8ToAVTwyXc//gzgS
1FPnCj4CrxbuY1r3hzRAyShArjcNL9Ou/lAqwco3eyeih+So9/0afuq1wBKu
w7o4zcRzCyHQSIFH3Xh7w4VN7vjmxIJyHlh9zWuxXyMDMlleq7ZojnYcUXef
VMe9mY6NXfraOdXOMuiaaHI6K8yNAxDn/naUvq+31+DJsRQXSxEe2NetFa5J
fqG7XmkKdqqqg24Xn5wdwohj90LvOy9FJ/J0OHMwKZ8B6RKxXx2+3AYLn7y1
Nlx6iLi5lp3m1y9hxNAQ9swpLCu+tD1s0Bql3yK2a1VSRROWeAaM0OZsd5yq
nqScmcVqHvIm2s0Ytz/F/WK1NoyxwFmDqT7mRdIEzPD+pV5Cyp+N5IeeGduR
zZpRMbjaYdnzDvbvSQHU63/HHpxDL2V+5crxIR21eZFFbksk7RyhcCGYdEaH
/+wCUlfrrbKz6lJhkgftTLflPtY+8q8qHUoS1kJolO4EL3ajr35G61gv3Teq
SC7cgiuOz3JuipNmwwrvzyAxxjbKDP5jZLRYKH2scOQ+4fgWlpw6TSdzYyH1
iZM6zY1G9KrklCwydYy9ip3Fa3wB0r2hyk+r0jxYt9xOsFX7UatKEGZpfXs8
nnN0EX5KeeEAxTvCduy2SU17Qi1hj5xTdrzD2SJ2P0bI+N6emvaMCQd8v05J
mhDlQi3RK27QotD/y8wHPsqHP55nLGxTCT56Xv65alRP0A4Mh0ONqIfw4GoT
jqTLrj3xRAa2A0Pobq7lggr6cWc0NRFLcVOUZ6I91WzOADZ3RSgIjf5/Wa7T
6h8tcCdQcXtznLOjpUkkNaJ0zGV4z4w8JuOZ/kWR6ltrTbcRtovGzCiKnVHM
w0939NTJZY8Oy2MLg3oEkdIYGqAbHifUEEOZtSmbpHciIlPmKsgd04gHxLwl
wEvF/6uYJ0TY+7kK8G8QE+He47UuoF8oF4JXzAmxTmzlb1KP79K2M49g6IHX
4Zr1N2GieBhdcwyMrl8RqBgu2ag395pE0RnReaf2SRq6MBFZkPoKuP1Kw6Np
zAD+Gf9O61MOk2kPtjm+64aCv5RMmq0z2PZfzuwx2wKeCg15MUJ0YRBqy2le
l5cjqB6xcYLFS9GdBbBeFJCJtSmC+6fQKXzeessnlQK0baG00fSDm27iTPtn
QKaruBguX712jVxAwzMNdnvzjrOHEWAUCKnxmdD04iDzlcIO60R8yyDrI8dG
2UKYvCFwvg8CVi6t5NcIhpG1To+eNvDf9CPadQfIbgHhdiOCm//IX5VpQU8e
xkMtvOoXeHfoPQ5D/h8nyg5/f0VvMeK8+dp54KhreycMoUBORDHBIB6WEkxq
GW5C84Qal7VNvg0bSmfU+GxRNGffaGDidsd7uKDdDdWzMhaRbWvrurKC/cZ1
8fE3NQyYv9Xvzcy3S5T9xdAZAD+7yg+6OdODvYpCxWEPTZQzNuuorJWdQH5A
yXb9uvAeaTz8GFOT+pm5CmN6QsODYv8nq3k5CzkQQq33jVjbBfVMvNRfYH/w
ELlKa7KZp5QZwy78DIpI4im7r/iTfuZ2At3H0OfLJpLK6yjcIuhTt9pZ5h5t
MpzkozTYUHEp5rdQ+c3gUgOdMtM4/Z02c7ouK6v6GORnmLmQ2fS1tVPD3R4g
SdMEpQ7//FZlqHAEtbbI58hXI0RgTX1DsjbU/QkIssZgfz4Vr+VOW1/znC0Q
W3xi45Psz6dEnLzWaFq1byhDfFATeTko3BRhdtRNTRWhu1+klbTII5mnuOsu
AamlwaYFLPaOuSEmhiMYCaNi4XsKGMKXQzxztyovF/lqSB1G+iK2wjMMznqb
uhBxyN5EnH7OtZZNXBlf2Q4hEpEmqNV4Iofm+NQHMkUorTsHruQc+H1tmLb0
LrqYpCQj4p3CvM/sPt8I2j0BPJhKgk+tdqXpl5gn07kVnxfmnKI2Lb81sNuL
KZizLHXzxiSI2dQRwe/N50mOKWFOn7tY0R8onzIsIHzGPPTI3suuczTKv7mo
qIS3+dwDju8lMBX/6hdKPgUemldL/uY2csaGYlqf+8oImMEIm2VPSfdR4zok
iWEkXFkSRHiTrkdxRp8DPOX3Fu0S2W4T+NIruaxApxGfznMwsHtnI+tMXeWG
WcbjaT7WBkFHgs2x+HSaT74C5saGfKUJzr6gTcvB1KXNrGAHSO6U+DK4tDBi
zhMljWyaX2qcNgkaYr0SlNvMdJDQgok3gohjACVYAeJR9alq9xxDmehe8EAw
YDmsNKPlUgtI4ESWyM8bObDmtQwuqwvVP1dX3Yt5d6MlCTYevq/sFt9akBfa
zZLUUI0rsCS2/bQnaNX9BSJb/pHg8py2PTp9aRFDuhk1FDyA4VsY0SZyN+Gr
ncmlbVlwEyMiPqFDHo4XGYEdZyVTF8n75M4lwsYBq0KgM0n/ALqYLX6cYGqX
+8XDrWmyra0UGOOsfshkj9D+/rSOLYFN0D/1K7gOt+/TXEhGsII6PXQH85tH
kgeCSMmiFEcNmj1cEGmu+x5UKhbYMDpMF6lknGUk7QKXpZkPItW+cY+/xr7Z
KEn31FsHTMWRE9SxG3OBhe6rLhFQ/teiFhMPDCuocjHb1UNnjKQGJvhDiq6z
StBbA9PxYbWI5Un84EdpICIzBurbuqzctuX4WLcbppxjK3pHwLBj2LQ6NQrQ
goQR7x6xO2Qofa4Ku1F/8pV6nKgMNtZ7Ds585iz73GqdhIJ2wbOe3LTOhUR1
K2H2GJgI97IT+OV7Oje4mZSYlE5+OhDITVljntbyBDJwE1P+ZsYVbOzlRMfw
rL0C4UR+OMobcfEj1PG46NDLYKaROUt8p2r0oZ0YrDfc861UeCx9py1Ha0Ry
sjmElEOF2pzz2TGn9vhEx+0+bcKpfBv56nsGz6x/LYeDaxH5AHM7/EeKB7i0
cYFcZl6xdezSSK8t7DdQ4aFHFtwIPJiJ6Aq3hAHjtpNvLH0+g1XZHZMb70YS
bSklpzV5NqOvyWhGu1mRSPz1Ibh21bsjsK1SejtTKsdjOzBLXx+LxAZ46c8t
x2Fm7h+HUk4s7hPCAEjEBE5BgFM6XH7GQLYPZwomnLxCXBngGVXa53YZ1hBq
IgWm95nwgR27avqfQJmRUuz37I7iD4bdEf4i5AdY65xPS92tPhhr/Vs5Xuue
2PyuK+ST/RT58xxCOKT/XeIhVBomAj4sDkCAstzki2T6/Om/i/Lb7N33Hw5q
kYd/T0cC+dCE2DJGO5+VT6eUal0JWUZSSbyfM3erM9g8N5FTav5M0kfNV0oW
RosIIThCjaz/okFv5+sHD+LxJlagjdj3sNlrykX7Z5jut3YaFk6F8kc9SkR5
XpV3cIExIl3HmcGyjirhrae9P6bJ1KFQfh4PyWIcZ66eRkPMjV+rkalNaLID
acTTYpSUmx9sbHNVC+Xusvwzff7NrhsJmxZvwF9cQgOWbRmIdn3cgpTMAF/1
o6jtk6sAkqgnT+pv2+j1jmOdDmcDJ1FdQl3rs8YAvIqPFy+ZPdtZ5EXk6Bzu
oaehCi/TdHtZY3AZ//fgi+BAuXZqsbo58rTf6LLkxVE8NFr63dM+24Vm4ZAa
2Bw08YcbZYFd9jD29WxZEFJoKzoxcCT4IJ5phHvk+bBYWiCN8ZOIYmgIkk/Q
z/AMmp/75Inzs6drrWgfymH6iOq076x5nIin1wRgyVwueF5wijiIkq52grRU
6SKJynHANnxdcSW5oSqC6Ln8xR9CHJitNwajxBqVnlQMlW9i1G55Yd9wz8ak
fRl2clc3iPc/vh8nfZOaykgDcH6HOZn7XdXcFKye/saTr2xQl3Toi4t+nGQz
3JN+F0d2n49u3+N5crEWlZhCYmqtx6/WCNw2qUx4mw98DWUyXb0r+j41Mkv/
h+TkdKcFFGqkOyEckDkwc8fVukPNzr6C98Uih4uswwDiVeMQGOlX6vRtmRA+
YArSmpbdJNijY/b8D9T+lK6jbmHBTFUXTpsrY2j/n0A47UpYFf8yzH7tZkF0
PSslbDzHMg7kc3/pDgyEFzlHWLMhwLgvYRG6puNibAWjnjrcxIbWr0xSzrDp
p8k1YLh94w/zi/LUY6mFUL+7DFz9zrUe2xoKPVKlLnDNsfmcmHjwGkvhF6IE
lD+4qicGel79k+4Iu/kZUHfxRX2KnsP82bFxmuqvzRKnRZnuKKJDWoq11RD2
ao5x8xqJF3+KNHM0AXgaBnvw+VRIeJbSvIO63F19CC1ghGxCJns1l2RlwX4W
07Vv/6U2g7okz3IjDI9IddKO0n8BjbErVXBM6k64+Mt975HAGtOJhVznhDfw
yHCGoUNf0qMKcwByofBdQbaCIUu+zjuwnlkQjEAk9WJ2Apwk8Sff5Duka6VV
e/+G1OLkN2glNIMp1J0zVO3gEyOZNvpwX3DMYdwxY8/lpsiro5Yotfx1Xbeu
U1WvOD3VEOMhflkDFPIK6Z9DZjEWdruI1GgJfb93/5L8QbKAPDM/4AeOrEjB
Di4PzhGKT1oqBcBUY8nEBf8Blybfzd+ABVt7/DHb95HroxBm3bYWzI42fftf
jMqfKzoNkVL0iUI0RauxrfsactcaAl4ffMLMXqO/wt8lE6PahfhShJ1pFMM0
5RKKkdaGHUKULDL5t/bDx3KxbOIqvxz00Yyyi89KryVSlUbYlfBmxrF8brAC
5le10YGHpW02nl+ElDxTL3xUXUQU2MjBWVfu+6vIWMa4gK6PPM9lSCCtDh+R
65yqbn03/Fbao2s3Zla6hIyfpFioQqBH2DTJga/Ggg5D3CJkQNHECucBa0hj
64AnVxtRRCvxvtN+RyVoCUIQME3DYqKRCHpOHyC4zcGkY9DqCtLuzrNI9hFI
clNguI2G1C1kF4TRIMXn0G4Xj9T+9eKMG0tYwv3bLw4ir+YfeSI57zyAhatR
L3w18I40ixwa1AnmyLSPktTfod9tGSqlhxoh89SZwa/a2WxYatFNhKMdz4el
5/tgKHp6WA9jIirrrWav/VTom+1VRgZtzUfpEVo/EKJ5T2f7x49AqWdtLpLW
xRe+6i4le0ahenBDievH5nXWFIY3rR9JwPl3fJYNsWzOj0pFwBkag60m7LQn
Jp0sNn1cBkB2uXZvi/93srYNbBKKbICgNbP6tMMRP7OPqr4wUh0PUGqa6MAw
0Fgv9u6o5o8gD9RwPllAZ4u1oX+ADz6qOiKcQB/I/MxgjEnFVZaAu7bOC7iR
gZpTzuwgmu2fZAd0cFZ/MulTGGrTgOn6hQnA4Zx66X0OaPj24zqMtSeSLh8u
26uka7yS/7ZA5/QL7Z4k+kU+OlNXpfCrmgkOrQ/ZtMPQGW7PbEeZF3c0jGR1
Pb6eFqD09Gxyr/YyHDWtV3K5yZOQ/GTvils/m57AoaUhVhE5Aqwe8T/hieyx
WtSJPXxOyRtZECr9RJ0MhP4SsVc0V00HRW+Ri27mSA953Ur2Wvr3Kf8rZvRN
tUgNi0t33m8xk+uk9sO4EUDxP1B8d9lmfVvt2c7Lm/AXjR2XCBei0YNXRP6v
NXnAE7jdZLPhPZOxj0mN52fgBwkqOdvpua2UPoq+SlOjDjAWP5hmguJ7vEie
UofLTYs/+bYPRNvPyhWS3UGwOzvqqOTYm6II4QwOiJRXY4ovKC7hy5sByWTl
F+758/qiHJZkaGtcszmEh4ZnZ4EUy9HQ2DHcxP93Rng0G4Mqd8vzAXLuPhbs
kAaP2HLGVrvLlFGlGBwF5IjN53C2uH9GSGoY6BlczSmHviNxKNsvAqeVhqUQ
O8u4p9g1Vh/rs5Qpm+E0SSYNdNA2W/ZKGA5NQ4ulrVBMoK5c2veF20vzqiVX
fiFOrdJuZTSaIOUE5XXyG8/R48l1wJhTS7CJ2/x0799YIuYzZCDH/knrIsOC
fDh7VDyWMCP+p1hlJ8Ir+hEf3XAHOL6L+nt3ED5IXeM4v5HtS+iYyPLRaX8O
c2Mr6xvVvv5Adn3QQvuWOtTPbUeRX/vRiOYFkTFLVAR5gS2huzh/onWTB9JJ
xP1FmMlvKL1hI6I99ri9dM0hJutW9PpGYLrGmwKn+N0pRxOLDtJ36FTgEceX
1r4kSMT25yaCtOIfUqQaZuFulc+T2h6UiEymRMHMmKYQ8hF5s6Px5yvLEMhK
47aUNP3UrCNufgnfa5b57aLB460SWQtJ8DgWxo7zFnosnytQH5dpeyg5p/cJ
Ldh9AH7kZ/2srpp0gtsTEn9VCPZdCNghZAxulxRpgwwxuCgj7uk6Qyu2du0I
fp7SF6t57sR6R3AXnSQYcKY1PKycyOCNQwcc4DHlMwwouWfJag3WwyjeMF8u
gzO3t6mPTTHGVB+J9sObdVW/7OnowCvox3ZWaPQ5n3GmSm7UoQ4OJ9dJT+Y6
QKuJ1gmukTT2nQZLHqyfI9CbA/E8MxO+gtEXMKJ1OH5kN62Ve2ENSOhdo59E
laF9VQo7QU3/GcsAK8gqkAtyQWEGrlkM6wpzp9z0CP9S9rXZ/dP/8C8bDqQH
OkbAw1yYlTvZvCZlb1JQIZovtFmIbm0lTVNH83ONowhEAGG1q9zEyjeNzTE1
ws9Tp6uEUP0+CQ9tdJufgWZCNhZgnC7hUvfzrv7k8XadG1GPC9Lj6TYoXcvP
GA+cwfaDq8UrdU6laXmJep3RisdxrNsSPr+vrFWkxgqkTdGCHhhrB+uW+b0f
9ow2mpJUjUvO7L+Z0Pxq5AOXELVVCB2tDwc3HfmlG5rkMkbDfXXytEhupYTh
/NMnzYqcmEPEjvcewFzzaSnkWqXnvc5LHuh85zOTEN7IyrhpYFeY8InA0sUF
BN/Syn0mREtW3Ui265oFpCWmrVKkbnakRB3PeYlR+Ydp8VyB0B9De/5bu2t/
GQGQqoaDgy3F3Q+myd7yoACt3fpDWN6fC0GrwZq+FvVErprqD8vrYyYquH8I
yy9/IOxz4yy+VcvN7SqHPQTRHg+zNTk6/WK/yzyUJjq8tnZhrCICHO2Kr4tK
Jgy2VPe3k6UN+HiNdFRgdJvMF/IIU7ZknGcLmLV6BXh3AZ0aKfWqG5+omf2t
Qb3kCyKkEPLVOq/Z9EWIhTiqbqEuhHJWqOQZkzSlmp2EfQ80jOqzuoraeVnC
dFG34faeU8FgdeyykJ6ewLB8jz2Rvph7JlmIBGS05cW8G7ia34wvri4uOUG8
E08D9dZtnkBRkt9XqIUMC2SwC5Sq34XCEsSGPAw/pTm0ZvDpIEZhi9XobCUt
fZpO8k6bATBhgXNwdqgaMFbIVKZ3V9R+DDA15qXecHjrqnbXpHuC+6VFpvh8
hF8/EmlNLD6beOFSmaFw7ZxGLY4ltQt+TE1SkseF19TIn+5owZffv1FYYl4E
X6dYoazNguiNecVkTgIPEdd9MsXnvP3coODave3ufMahCyV9sV04ePphgDop
zNoJ73RGAamUlMrtFAsSa1HzjN9AA1C/qIrKbQZXGhUwvYx+7rIQbKivfD6y
PL1U73D3xYxMRKVfQrK08RB9qlTLoKs1OqN6+xgqdwmGgEaVW5zZDL15KJ0t
+hNOFk92RWUxXIVomHZQ0jIlQIOzzyBavCCBwFR16pSUcEP816OtVg4f+1/y
97A6CD7faw1rk86CkbB0Cx47uaJjY7uAazzZKacumo824CVGze0sks7N9BdE
GrGpBS0aRvTDHwPyd2QNiX5jkhAa8cKmWO+7vnvH13Y9xfylLW8j2pv4t9Zp
pqiepmilIHhMiKOwUoPvbRHGHpGIvDFdlXj+a0f/lsiuT/rwWnOdjf+FlgJZ
vLz1ZWy4xumi2rWGTpZYfh65ljXQ1nKoHpT30j07DP9G2nNsWMuTWAcU4C2E
qZhAGg2SQZG9KV4ePiXyxi3Grl8JybGD0Wqc2Ddy72st3ANbA7YzmNlAGY51
egUKZrkWLov+eIIf5SC8Aj54YsHvOPnK6idQxRhpP1V6cOb06pOJAKqzhP/n
+PUH4c1vYphiEwkP2SzsdPLKU/q1edJkFtAIMNEf8aZXx9gujIptKtW5HDcp
pOVg2SZ9N6HR3FzepTnaOeheJsQkLgjFe5D6vRmI/qxrqPGFTFk5Id9ATUvK
+dc2681rN7DR0XIW+A9M8VNC52SGHHwiUqJRRQ32ewuhwqB1ghqER+EEaoNo
bjfwHgRjDYzq1AnbOdIkXN/qtGtDX+UztSNOOoUYP05YHnwgM/SsuRztBJJS
vx4DOAHv+S8GXitCr1bViJvcyahW1ZU3JarpBmefxGeM+u4dSdgJ9zD3y5g0
PNFZ1qLTZg10JlI2tKkyeSxg4qjXjPg09VB7+Q8/ejPAqO2a0D5IxOLf+W+R
h4OS5n/NHslmoPx3uOxNl9N+KzXNkz/y4F9Q6spa59ZnCpo5rncmST29hw5G
hANMU9xe5UbsuoeBIo5015kXBkRS182kRuPHfgPPl5bhQycUUiuJUhG1I/cI
MYolFpb+N3nFQ+8Lpq75e4Mn50sOt6a7CcA3QQ/vY6gXc7OMuaiKzUwhT4FX
DOvtRIZ5RY4P/VexvN6juTBv6+DIZUACzO+ANTO4oOXwTwZA4XzbrF+RKFWz
e/CJT5jGLo6uExLdRX1V/eDjijbsZu4xpUgwK5DBC0gXmuSB3mHXjLUlvY8l
K+vYYCz3DSrP5Is7RGOA5PwTtnLyX8rqlxEHvcGl7I4h288PVlFHBgjQUXSU
qfLGgsl+nlJGg6QrUH/i8n5WUsYG6CzxhbrNsocdqvaXUbjpB/e9G0LeZSrN
+0fs3BUNn/xhkRzNF7Q70cbyaCLKtfXMGqiz0xHG1BRcR7/q7/Wdz/8qdY2o
MvMkQoYmfsViZM1gXqWG5s1VOhMY/RJyIkHOXPF1tE5uM49x8C2tffNIBt62
lgaEro3ur6dV9N2rSMFI57BmjkqdMuCGo8QRF2Tv6cev2zdd6GtiABkK+cQL
PkqO+QI0WVixKn9HuxvRGEoDRv81ze5bLSpqP5ZrqCuvMzrUbRumY69JabU7
lor6NBUgLJmK97kQdWdflukXlxsjK9lxM+BMW+t0lbKjDy9/+x+MAFk1h098
3rw4HkLXMs+mHb9riAvxp34YaPkh0HuQ9mTQYQ6/CyofzW74XDdvN3GY9K8D
3VbpMLtxRYmHJojUsItok8VwDhPqwu69c67c/4238PpP7Dr4tVDR3iJQ8bPL
vhfMHD60Yx62fogB2GoQUR7Jy0jUqfjd72+3fomvn1LJ4tsMANeU80jIGOlS
bMnyESifSWgu7etVk+bRaZR4yx+yYUTmWMjtCPpgR5XdSmFbWYLYuPIBbFFA
Fx8fWw0jFw8sAKXoZGBhOPfSDf2JODUkIINTChjhckXbnMUMX3VVlQ6LbxEU
viy6hlDDo9JOcFwlkXIfOrwiz13NdLffPkq1mwkkgDVqybhQq5qhsmEvzAgW
ZRwEDGwxSyjPK7mBK79cJyrHZ8m8/fUDIOroIbmVoyAsVARWwHXC6z0RTZvO
RnnetN0mnwObT/3Pz664hDeoH8fYGrl8gahIqZThhzAqMP70O29E5ZoWVete
k1m1sutIJeogmKTYxW4SYJPSAP1b4sxCBPBBh5iotsuGBVyuecMWrrgIgVHv
kaJslZ+m+dAdzJrVgi3NYgh89kUV09Pc+tSNQbtzPSL//lsDkrV9CDVv1Z1a
oqtMxW4GzroPUP3brU0iE6aBCu1V2Bv3imTT8ncSN6Y28LMoA0pUyD42S4kc
bVK/YbrN03jhZIf1t4R+d6Umr6BlL/exeANj8Wm/6kTG+G8vgT7crZ9HS91v
4f2DQqC+cKu6R2DL8W0vQlwUO5enZnK1iAArGYVA+uF7/7wkX4V/7uDOuL/k
bBxjnLh0jQWyiJpFBY4xuikF+5nDjuZ3Jw7QUbE1h7PmAM+RszV29SHFnI5W
j/h7kG0uSkI02k3cCgJLaiHLAnTvDNT4srQ5j61ivEiJnDmoGq/NEKlq78gI
gVMknjZV97Cxf2eYu0lSaCprZ7VSvc3d59Y9b2YQhfl+h/r8+epmidUrhhXS
MEbxq0k/JjSUqItF+wbsUUHBStYuHLwQWp4MrJyEF/Y8dC+fe85t4Px5QaSR
gigTRZDyTFZFbYUzoClH/AZTbKtW1atacPyP9UifCt81vQPxQPSRIkZA6mL/
cA3AgjBDGP+qwNoZCFm+oAetpSaTMfqK9JxY2MlFBqyV6ac2rZNXFU2glJ0t
YmMBW0WusSdXWhPxM65P2843/YfriaOg7O7O/oqoHtvhBa5nb9JRf72cKw32
rs9kHcixKGnKHDSXz9z79kJcAyMf81hGAolvQSTw5dr4shWSq9jD5I5jCQhV
oVv5EUoiF/vWchS9jOVmtpPoppm7SnJ476YMQCdc66zR5W7Jb0rgaLNSQNxD
mzsBxjp5eamUSf4ngg8OfW+sjvHdQrztEPjIvjeAqwUdYuj/BoV9mKLoYoRT
vu+aOqM9S9B5BrJ1pMLJ8A8XNqsyBJIoe7TIMW0oPwnRRE3IlJu+i9KycL5C
yllmu/c1ZjHwayxisXI8KzLnYhXf+ceQLlisusaR3VYbYlDlJVOBE3pYbgCb
NXON0qr2SuQHwHuRLiQiTKarazjWrqwikMcKI3n4BkH6gun2RS1odgxagkXw
kSoqh84K8E7J03356i6u/EkZXNy/x6A9+Sx8hREN95A2jMt9hearVFjGODAB
VRttRXYvwETVmtb5cON46eaI9jkNp39VJcoB6FIp26g5pfrKI6J4RzJnLxKa
+kEGclzTdVamepN/mZQ6vNeWoDPJT+9izWvX7KcNrBdMnZMXkFw8jLbYCtNs
mINBpBxKQdtW1pRTiXg4SnaeU0YQAAVuT1JHryor34/t6DO6+qSG4mS238Do
jj4GoFAfajCZefOqby4jJnnplBpF7KElEX3fVjTbslM4ICzGoTrHyPDwazq1
8NYLvSGBYq0EvsLC7roKcSrDdFmh06VpoSJGQMguyYRiziuXcPSvhp1aSeZb
yM1v6JAdaMEy1J5t0MejJWWjNHykLyl25N5M+jBenrxC7OAajYlvtDu4jhDV
A/8HILeRuEtLDnAU2U7ouxed30Mas5LLutnY/HRAFFVP6SDpVrVjBNobZkOv
sW/AVIXx+2UyjD087VLHfDOe0/y/ErxYx42DCNa7vhYH3d+IQHf2pkmvBFeA
tBkFuW1v1qA9bLCoKCZpkW9x3yH+VWD3IBpk5iAsqfoD8Lw6j3SZEVGWMFXW
zc1svp8ZHZj5Y5mdXNePVvlewfuGQ+N7Pb6OfTwTmUDZR8UnJhydnjatGYdG
cvUv9bSA0CjNkMKKsgmVLZWqmk/qjPxkU6vdE2gqBCA9Zau6RbVkhCBkKIA4
Kv0PSUGL03P0+z1QJeJDc/K9nTuzoaL9Trj5FudcI0BWuKLmOH1ZGezievTf
ndXaFvtz/xMzAZ3eFkIL1acgPh8GACBSS74COjfEWtfVD4NsoxyhPmkNKtR0
5/XYo3YyvpfSeFjp9Mr8gEDBJ0zh4SFaCbwn5mWHMvQ/QF1Z5Z2QJ4Bo3PoA
7eaBqe218GL/MMt5Waqo6kcyYhXGQsiNoEJdvIi7xCtIbLyVtYzdDaP/AaMw
l4oumA+UV4Il4AZUEu7Nz39gtfKYnrXOD6gFl1sgNf4WfDYENHiDBT0ESnon
Lk7D1a5dpTanOi65fBIVUEuu9NvkCTVRqXXFRU/OGDrHEZ9vqS4myqA64/gJ
l8o0ALEsMFWHREwKHHo5ojytCfaf+wG3+HLs9fWIh3YMo004phHVA8VH1J2r
0QwSQtyUYm5LRRW7IeVB5+94Q3YQJCERHyhPfZVI8pdl+onrprFqMxRc7+vz
7pV+tEXdoaRB2/Sy3WL+Dxe2wHSj7DkOx8tJqITgL5svX+wfz9LoyQHvtes5
oDOGAAQQ583x3oDbTnPTLI+zhfk0FvQ1iGjnZ9W35HGBrAXYduqtwTGqa5UN
8mRQFcWoy7JBnGCZtoVF22z1cD/TFuBoS6X8vu3ZVtM/qZWDdA+T7ltqC8eT
rAiscitNNl5ecFfnWADE/URHh3pZUQRPpLjS+jeAiB+JhJFk98s73EaR2CxC
M9cWGNO9uMfy1ZXd3AFLR+JtvML7xOBspxbt5DTiYAz/JEhy6MS2M733UoT8
BbrdyTuAa0jmaXJNrPxAtVBQDqzRQ5QC31QwwIkAlzsjossrUtN0zrLIULMz
5ZlF3cwp7zt3hE1xtLt3ubJ+xF5imgb1K+QA3Pzhz3yLw0va42jlZLNcKphZ
reaPAjUZNR+hgr0tcrFXdY9tjM96g4/qpg50Z08Z8EC0R+JiQSAxkurFchV2
yzFuhu6eJbkllFFGOV0Toj7T0hCxcNdVDFRSDHRzll1bAhhaCAlaVHMoIXQQ
gatqkTJJnULsS4msEUTB0r6kJPXMBC6DZ06lEg3jLcafUTKlau2V0ZHhpQNR
tai3MGBIk54xvAlR879jI29oXIcGlQBcATUSBosOapdnBLpmB5bRnp58VsUy
DIlwDCF4MauhXXKeBfzJAjsPO9HYBPf6mkidZFwlhmDPjPiuG7ZH7aykfKp2
XWr12og/67J37yysS7f+Rm0z1PqoX9mfRPsfrdS8OoDyv5JZVsOGHav5JDlT
evGnoqZxa15Y/GBifPERHmwNYxF4O1BdTognG1zVzcNXGP7KLIhSh+aqDKK+
OYKo4hv00IxmKjZYy6/njD5IqHYOt+xfFn5dWgENDL1PAcypPmoa+xGZVg93
pG9OcXZst5qLKO8PUr49E2V4djC0P1sIaWoX4LHb1gbejdSH8hKn91WFY6j3
jVbx0pzrU5PMkvkointuCRGe2I0/XQ3mxzHGZgGCx2Mu+YSDooAY69/PUgkC
+xoGkvfwCN6Exv+wvH7O1GRh/3RuAAgIo0RrUN6+Nr4+WaVPfd0O66HNWvmK
2HV5xwFq1lArrnJ5gP+kiB3AqippjkRJBNUc6/O/IlAIL4d6Z99AXXbG8k/n
Kbglg4w/9i6n7FXrDZsv0DdvDT3cYkdqwRkuTKtcpKZZ+sCUBQIZ5DwzUWh/
dpcx9Yhugz6p55p+FDyu6yx8W8tuCPM2ziIAKcW6zJ70CSbu9Y8N8M+sjlhI
Otx+2KrwtZ8R5qqvYuN/3Yi6/8ZbkmeyzH0dzyDqgF92je4yoDg12SzbVpRz
O9NJFYdHwyghm4mR63+uxqr/OHboLxTaPROR2O4vYRiiMZ+bz/i8w3pLYSIt
ah/XlEKVBzqP8akqMsM6szHps3m+9sOw913Ks2NjpJtCophtrWEQJ3migpoP
c7HJRAwMgXYQsPuRUf8zSTouj8PUSIT5LNkeMZ1xsxl0aWVNhSBUqSzh0Jhf
gVtAilLcSeyhpap438di4LPdLUSdi02KT+97A2WMU1AMkxS1fyq6rmnGSsXt
bnoBl2Xh9AtoR4w4va0iNsHNoLW54CEVFo3aZJvKUHMwjdkFoB2ILiW4fTC/
36gPwLOvD/JYCTQPKTabg0z6DEIzfCDTKeKw9G9aSXxabM4QOPOK/AsXdZ/3
aesBTdkTSwK6GKayPNZAaQy2eH9i7CIDJEYJpWLmjXAmOCvjHZynR8Hwo7e+
YiU/ylErvqoLJVeINiVwEbqVwgABeozRi+Yb0U3fUXVgJIkZI4gD1q5KSN78
NkGbRQupHtF0nsdqOo6Pv6a8CYVrZuiymxuQJ+h3TsSvwQXAbDBrei7XzJK6
BFraxWUZR9+dRjCSqTtvWZ6D1HWw56BnURA07/CyHHxcJSbOys9UqI1QUOwf
pgusrYMIKOBIPSPIPMbh2N19Fgp1zlmpmmSw1n1y0B2qYAPG8Z30viedC97t
EVIW3Cd9y75LwM7OaRBzR3yWUccX0g/rRUh3F0N2cuGxLogJ1axzso0OXtHC
5RwLecWvzeyRIuYIIO6IluOpivjNF/EBODQZP0H2LDFVBMOCjYe3971Tkp1Z
7SSrIHTwiZ1O0KPIQz7ieZ9UKabQI/kYOEd6wwsE4Y2YvCW3Dks59TAReNCJ
s8MjzopDcajBwOejjJlCCRiyj+8UT0apxpfaozF6DL2WLgYlOC3b5sBn5yoC
/JuUP3bkIJelVMs5OJ6YGrlLoIuNMglbMcLyRFU+tsKOl2UZOmz1HhugZgbW
pWGWO6BsQWTB4W0pRi42vhgWUcTO+fLXJPuxOoqsJNEmAeqmeiJM1btEFOI0
1YHywnB6+3jckq/i+kzhCRbxbaeERkvveWVULtF+DN0mXkOPenuQOvfLoWIa
Xb4qtwIeqvxSb+z6JZ4ij4e+AJ8p3NaI0gMQ/nMbTbLM8qt5yL4wRGL7hhAZ
PLtgoQkAcON99D6uW3sDP8Uew6qXXaWo6MVBsI1nXTsarsujjwwYER7RG8JU
DmxzzZEBX/esDa6e49/eDgER6io8tfHd4b2VFWyKjXcmYa9nSADMlCmnOAW6
gLGUpesdzolqFvz6BfMHLHXSBxWVxH3x2JmcFWUCqtJMeOyjDWf6hhKp0lCB
rT9LeYiHSdRdfWVfe52593OJZ7O558V7pD6PaTXD1r9ZPISR0lhFXD0tSerK
3lgwN+A3uZNA6VllFVRaM0xQ+M3uw3WXVApzA7utVFNkFCYuLGES6EPidWIE
CBjfAqTVuaYxJli/6IrHf4+DAX3gwUU7iBNLXqXn2+4ujYBnymx+p5fV/rwW
5gVcl/isl0G9VxWiibGKsnMdRpMtCbr3Dk99zYPJElWeXVy+uulJUbH5wgYL
4oThcvMW8MYEooKX7w1KSW6+fJhVZCF6HeT2a8yLD9Eg4AW4/4byJON4l96U
zNLEtL7cLTLyUAYfOxR0qdkthseAxNGC+O/UPaKktoZ1lgK8Pvi5jFoqSoav
O4eo6dzsJoggozlncDbBcvy2ic6ZNv4w/UOHOPkIPimsFYlbuA6dT1C7YTGc
6uDuamEAxWg0DpZIrVyWwIr3gGQlw9o2kLnDtz+gXEfz5UzGtP0J6deLxP19
PufH/jxyzq47ETthC2PRQPU4PA4KCQNAt/4Cqtu9FYn1offMSGKCrdbd6Nd2
eirXzi5HtCk4z5h62U/RAHT5Q9NAamir1SOGbjOnFz9W1AOl+HmhsHKOHohW
rZ6dkiXwQ/2T53KpYtgePEjSrgM1QziAP6JEqDjVlc4PkUBf73Mz0t8IIBgS
bly5YgFPrUT/XH0KoxrrWbto7sQE8rHQfic+jnZAg3W4tb9I+LRlihIm60Zj
njfNoPs5BtkwbdKNdYsZkM2pU460tTTUViJg6MRTebDrd99V6bcQ2Y7q1arl
/nIYcHzNsiaiw1U/jpt8GLJD59Es2ahzZ2n1RL4+hde1BpYisU+vuptuapmL
yIn0o+qkMWgz797DUvX/tN9wSk1Y7hi+tWNb87yw9/1YGQa6NV9XHblVhP/5
D92dwFs8TPev+BQroLAlMazR2+3lBUuDAWhNJLErJcNE/n3i324EsxQkTQGR
fjlWsDKcXpb4Od0fkEIxp+Dwl7vOuzwZDz9fahFOPoT5cUyhJpXx6L/5Obvf
PcO227q5BB7RfHjtNVBY7HQFuk6CKapLCOOc43Zx8nYnQ7t+DWg4gBJQgzP3
+gaYtv/1IgSnWLvYmIkAdtQMq8jIIoo4+B4nDcjoPKytUGm/tmiQ1uufJZy2
SJumk2rGNqll1oGsx8OD73xdbjXTrRUDH+fLfopiRg2EyCd92BiEwA9/fvUA
GrPXU9JI58TW5YoZMGWD7pDBkKSOo/7Tx33VUYH39lhvNcRSc84VDL4BreYB
ceC++qkGswaaHzOleBTM/kxex6IF6ugWCnDyTlyE4q6ygry1L+ahtwHNY679
AZ/hIywYNs4Fceh4FD5jRWDQbTtrCcFkN27AZIkQAD2lsJMHdsiFwX7XnJxr
W+Y1zcS9zOmA3lW72q52xqDjEV49TqwGqhCl+NnAz9UUc1/rkdN9sOKmoaEs
DHZ4BYv5evXu3+ShQ+foWk1NqLU7aUv6XIRWg8WQIRc7GLAOnAoz2SXhKR3L
tALlXiSeTrJgSyB/wgKAwz3Of/hxzGcW03OsBIpbp8oq3PAQoTJL7CB/LJxQ
ZWXj1y7LPOOjWoHKXZwIveChMyc9Kzskg9N94rr7TKdslqXo6G4KgF7p7XU1
9jbMz9vxJKJgOYIuYeYEg4C/5WigpxjxpThARLzq8sRlJKzjyksKCD9udQ8n
aYuF6voBoi9oyeHT5QBWMnSGPKgJQoSfSuvI/BtLYPzRYtbaqLfHCFCz7JPZ
xJF16sMIMb6YA3oTKwgBNm88+8mO1GlJMefAC+4/6nAIHHxt2tfUK4mGXPcY
vEkSWMILigHhWG5DaEDnaRC7ZRAthNWUgAM6sb1yYPaFBk/uAzIuCc3+lrPw
er23bBYBhnYE5iN2/ywYPjK4xXarTTVlPnYFH+lvBYhdGlT+aUKOvCrBKxaX
BMVIwWEUpBg6+r3a6H2I5gqT+C1CJzjFrtaRK0CNm5CfIlK9r+DzZIKeK3VC
szNoND3SJQagWkeecBj69gKpBtmjbcyhvxbQ5U7QcBDspokMVLJnsKuDk1R7
3VWPU68J9oq5RJbi8Zlpzux8xub5kK0mNxBNE+Wnc0X3RKTkVnYzcDXruahO
hLuOVUQ8zeGVf+RRkGgInQFKmuVaXLMxWgYHiChIG2DIDA6SvSX9NSFusvoE
KVQ4hp/MY6AxroqF/xDf49/m6GOlvVqdjTfWwNc504ffYSK2UsoD71Min7FJ
Md27UqKFu2gf6NfD16Z7FBBaqZt9aqoxdGafjF/X4cV3Gjggu8a+8hYk/s2F
2H61TG8lSZXmjO8HJNe/yppCfrX5LOnMwOUd8vmK6xkHUEhjZcEpM7qHftQc
CMikxEe5jkFb1k0GL3ACboHxnLk7wDXGuPURUsujv8CJ28KOjXroL7ydgX/3
Cv1kCG9m47A1Zc37qIzQlDWWtmL07HYaoD4FtbpH0x5WuBSQ3pHQEC+ZUzcR
xFsqP02aAjOKc+f32kunprvFxoW+VA4u0NJF5R8+7U88gT/LuMYj0ZbuEvxE
Ia7ZL7IDvKtT5EivDCfop2markoJzvwYaOHBpgFxLFNFhYk1AhMBqqTfePKb
8tG6j03/9jx8z1EeDeRlJ0OSvac3nLCb/Y4UcGQ7lcwjJPiMT+RhrV2hMiNy
Iv3A7KILfME8iMoUxXkHh73B3YXu24aUWY99cD2KqeKfnRdo0YAV5kyfOfLM
NvTw5cszqvf9k1P9W0VuNSJfhnRLPYf9z9vsaTZ4q07kKKMSX1nyHRfa9/fT
EFsk6MJQ/gIcJsk0cEiHSGlVIKGtQzxaydXYWO9qewfGMaW/7tytxRfUZm1U
vzbb7qFMoMDFDAu/rpjxiSDSSBj4Q8w5m9zeGFG6USzjV4QkloQk7gwT0nH2
mFNrQYPdr93d/HaUPBP+zasetd6n5d6Rmfa7Pvai2EMg1dZFGXu87O2naFBT
Vh6PTt2x1pmyavA3BkaL3yZfzZ2q32YrzH3mBd2ryNzRDrRTvIBmZUzlDwbK
PnBUh6nZtMns3S6a4vaRdV1FxxXBbOQDUBI1W3PboHZzw/cFsaQMx2Rbo2Ww
KbWNWiQjUzDTw70y5RlAfwbwokHEtgPml8+ZUCfnfdcTKskJ/89qdiwW4oD7
L0wnSwcyMjreqQGg1DAqodXgqi2HJz0aN7PVYgLLUZS2bNxRVpG4fTxIrWPm
Yx1bPlID+aDUBA17qDOS4gzaSkkPmUA6AfD6T5pewz3frhAunDhhOhUyHAy/
rEi3NeuBVNNVBLPbpdjcmzbNC8FYX4m1n4npQPyNvOuVU7OJZUjYbX8LD6tP
vo8yxfwwIozWeViQfMgC3/hckR+D6+hgwpE4Cnnyb2UjFgy71bk8+RyOwZwF
VdLrkonB4uVVkk/zsiy8vX76uHT62FvLfBsyMltyT7lzwr2hTmSJw5Qb/KlJ
flY4sMPiCIhSum5K8kPIQXQycJgWJe+gNu3ETSwp9v6mBcyySriy/DUUynLn
jp/8X8/WBaFMWAfFw6JFKciHUD7fu2F9wUmfaOeCIIxFVWfFOYLVBbR47baP
G6gJn5l1kX5/tIQBh00s5FH4KnOWHaobcW9Ryoku4lLaWLNhtTekUzWBdtVo
58WjFkE6qkpU0q1fDYRxeeDJjAGE6YZmU+utcf236W+NtzUkJfhmH0z1Q6Ef
ZVcsvAddmqKIDL2olboWgt7sZVgUiApkZ0lAXgI+4Dp4CAwEAgkYxNqkMruv
tZufi+2Y/Mv+V1J12xRPD7g4AFjn6JbqXF1RBdxyjxJ2hrFOd4BpPcBxCIRp
eFmO5X8v9mOntHpPjTiaAHlPdNdnIRxspVyD3W5adNOI7uY7nJAfsWuQI9TX
8/VLweu2/CVrqgBQ4HiI+MRyFj3yxYMcoKfZc8WJTtXmP0L7q484hHnut/aP
Bt5ZrIaozDEHxQZ0XfhW925Pj//LSot1N+/gUYjsbOnMlL9npC7Ogh6EOM/c
OyV8WKz7JGV6ecj0ubp3qczUm+S5Hl9CESdqhQOzRKaQmbDYqBbQdAGiHj8F
iOnnlFBQ20QR3EZFjoV5t00vqkSO9lS+ekDzXALyv5HBPX/Gnk6qVnGfIbE0
JTiZfb2HB7ZcR7TXw9+SWe5QAnv77FnIosZiegAPMEBO4QjJLhCvN8qVtZNc
SbcUzJUcrZwHAJI6VYQDghqQyVPoFg0C0sA2mxbYBmsz3zz2vI+dGmHdbqba
1ZEdkyp8di9gIGYc3Sk2ZoaJSFOBz+JppvObj8WQ/Y5Lq+0yjcDt03COJrbx
F7mL/l4ORiKt3dnrExb6+J1FWkFCshYcjHk8qL4BITmrvDlB6jY5G768rpIr
ZRsD2SfkdP+jmbBK3Yf57jvEmFM6iXBSrb31kvGzJF9o8LKp71FQ0nK8JutK
T4pId22Rzv7bth6OK2sKp4ibUtV60u2oXK3LI4TEbVy9hWGsKu9U1/aYQyCF
VLpAvSJvd8bEt4pcZFBukUS5716Nn4JI4vJevdSauNYG0rmJ92EwuiryS4xv
E9RytCRl2ZoXxMmbWKofCLb3MG0DI2cacLb/dtWe6O0sU5Cvj+Zb8ZbVzzxN
vLmV3AyOCtSlJP1Yk32kttPVC/suoRv0fzjsPPyx0YxBz/2dap9qTzyclk3q
DSlwbJFkXu5/UhekL2VZCDC1OekpEeGUEFpaIbZI0uSBbjPM29EXRk4LHrA4
l88ayG+yvSujZzQlUShu2EaluyflTwt4w6IwUf7pnE2p3EJkESm3nJPb5iWu
AIH3oy7RyFwGqnOSU5+uDSLjeKXUhdOQByPnHDCJ89W9VdYgsuhhsQl7PPvD
midt5ew3EDHlvZPlIIqMVO6YHMZ7exsqom4P2oZWvjkb1qMo3kK62owbZ+a1
+1hdeeF3DtAYn6jQEJN2b0OhNUcpQkaeHjKIxNTnjChG51yvfhm2uIA8T23r
Gc9j5KU503l9f0KpjSnhyF91v1zva9lmF5DGvpF0DjOHecgU5HId6oT8c0K+
c5KKMMq1FpGn3AkjEkxSSNj9Hn0pIijzsgfYbZBH7rMkKUZ9A8UAHvZdOT73
IHk75Jv3ST8X/TDa2Wbr7SA0An71QXeuDRhj3WiLK00l7vQhIq/p/8da03Hk
yIdGJNzGL8y3f2hu4FkpZ1YMw+SIalXVgmfwht8mUPS9Sk46JwpDhb+7QOsy
dYLD2eV1GZX7nFdNF+ORSfm3zvh2t/cedTGaF9R4x2G248iGJ00k2Fxi8kCp
5YoKL/52hjV/hrm/coFN74DqsFU/aLLEAN7OWuF7T6kn6o3sGLoXug2P/G79
q2TP2+EHklCDqeL4+esHdzmHAxUnZPKzWaefsyZShY6OTuYpKMcWUQWx5yfO
09rYpuouLSsZuqqCjeBFNs6cttnEKSbC20nDLUjxrby0D8H7TefIvYV2GFSH
XHutIUoRi1nSkpXWGXYPhrP1NRbCNnlKS6NXY9pFbShIWehYrWeFpeCkkrhI
jDEJau5qTp0d1wtP9egLnuDdledl/PcqA9q49tB9NoOHeoTtMaiANyp0OV0R
HXEviy8lsHb8uTTgN+s0VynrnC7vu6H9zVbUBK0LKsHwqLfeQahMyZylSWLZ
c1bBecnYts7oqvzLeXcyCUjdI5krZ2vZnBSU0+AgGgFuZ0PqFBAXGL2kWFKF
4smsvHrHpL6c/Q+TE36Hlv7jnQhovhYw203uAZGtfXFsUBfvU4Yon0E2mc2u
TzRTVJlbuqVW2mPHu60lsqHckTUb4W5Yfjg94n2mLuaVLbddMSMxyEEkd80d
6GjejA4SjdLDEZU74RYUBqfGaP/1tfP5IZsHhjAhz2IayBoJ7hj6lzucrMFD
v1oOSURrD3B9xLxOiF6+DoLml3OLNKd6Mh7JNGO8C7cTDjVkg35r/0Y81gCm
Lqv8b7f4PMLx/txa8cPVbOWXP4g1bsIfbJWITpr4qcauKFCk4pCdlRL7dzo/
Pnv65iq+LS9y2JV1o+5PHMxQqRLTXSCgWZhNBr+JbGsYdUPTNe5DuzecVCYE
ZhLcw5PaSu9lHH6l+aNF5rjS3Z+GFk2Iuk341gQWoy/5Rr5gQDlc71brJsWE
fGLyC7TlswHAN/NFeZ5s0G79GQb2DTCu9LnpRfLV/fFDbXwSVGsJEGHmmDtS
pdInvmVRf9Z9nn68VyvND/re3da3D03zN69dPBiLMGmNGvYusmqIbR6yA5t0
ARMJd703eNdIeAu6pLboGjtnH6Vkp2RmcHs9o7RKQLgjc9rNp54M/7UEemIC
d04ieihq5KzaMsO9CGeDZ+V5hIRI9grE5XvtbFfReDt6Hntw+cIP/1IZAbgg
vamzbyEwKl8Az0PBX8e6pInVeows9S+hCbivfztfVZMxG+V2u3ZgqqYtFENn
I3G0oOOfvHB6451NBlqL8ND39NqfrMnrlj7DWTJpjGkjMy7b+QyC15wYpYFu
XWELhrISn8sXUYrxHBDEzPZFtaQGlQZHJEdQxvo053aSrmAuy+EKvfyrMxns
CNboGb8GGpKcX+oE4Q6Yvg5xX4/xh3uFFwtAryEJwVn92nkyF+sLrpRlEFFY
OeBqQ0V094l3LIoHluTQeGqE1lNUU7p8DYCryRdJ4KV7YBXUEuzKzUCITTXU
VLqrp5dIJc+R4jHQBRgRCxsj2RTx2BGB5fqgLaeCPWbJW5Lr7Xn0U7rIcPNa
LLEfslPgVfqYSorG0UMTqClt1oeZbLMtFdRWJyILCbNqDmHo89Qi8mH6GE6X
eVNPrSYFKHLbVmuu5aOO2MbREJa+njDPHoeFJ63cE3SvZWOo0B4Es8YaU0+9
q/0tMW3imLBWVcBPxoR99izYs0MnAm3E9pm5dfYz72/Ch3QdhgLziyXFdrCM
M40GLq82zrWpXc+lr2gmxEqf+6c/IqTZliub6H7/dJWCO/3pHI4DQoyrjarH
GEXGxINxXY5QMZeRMOD1M5zJZ40zpBy58EoSeecVe1zehHMWnw82SX1Cb0k8
YYqeqEXAKkXSsObv+6M+ABR0hSZEUHoheYJQxRmXSQO4jVEN0XDKkcuL1+ec
5GqQTRXIETQBj/DPB/PVM7Wn4WZwhvdfCpZDwG/dR/hCry69Gsw9t/PgW3bx
0mvI8L/wGlCAsVwWxBqmGV8Rvwtmz6ueXpDTYSPw4KGl2DGG9gpGpnaFyxxn
AF9koefSYJPgxGgc7t7VynXPMYsa4hDpHzzZkkjkwMJcpPOuwE2xEDiyA7Jg
4T3IyCeYZgO+Z0xPIwm0MR2Trxj6cN5HMocYu3CygU+3YW3Nu1TbbaeSXcQi
zLPR12WqXOjil/+7dT7eykfe3kUeeYuVEik45Avn3fYSIfD5szkqp5+CMU8C
qvujNItmzIWCsSAnYGuJi6uyobqDhEPaCBuPV+/qEuTj2x7qD/aDSjmj5EX4
VMSmCb/JhILEtMu2+0mEFhdVsPbdeRdfbVfUQiKOY72aV3PVfB0XUFlI2kMr
AFfVqokxBzs52hrnJOMjas72RsHf5LV1S5h+ieQIk2yWVwH88lNQqeWqzekK
l9o59MoxDmoVPdZ5LGLK4ZeDnuFKtAdAVgGMBJTngLuNv+l9LZehGTpso/j4
mMGJHOFqKJCRGxfD0oLNPCOgISbPczsdbsPLFDV5S3hzZHKnbxmtIVzTeuvf
JJ2lctRcDG0fpq5qTCOiC0r4p1gORoAdKHoINS0aW+e9X6lBD3qnLUNcCn2N
Cntl+lUOCleHlVfRITJHuRZ+G+hhHDueuVc9Hmf8SVIESACSmhSwUOPNmoXj
duFgzeJpEAlRgBIT2X03y9XXjtiXtfoYkV9+tYcfSVEbYoShRI2MH/pkDyA/
o0HAf6hVtMb2kC2/6njDpbGwo09K24kzo82KvZPeIc8LVHA1lQFWhjhLO6CD
Pi6Apu2b8Gb/16cb4PGVJcK5v1i+XEf0E5oYwzsOIV1rNJW1uwnybqSzxDnV
mFmly+6pEISvzRHaqF0ih4MdOY5tNgWwgVj/31bfNnFO+FNifUgtMJLhTCFb
uISEKaJiikRRvxHwq14qafpjmlzCueVRAUwC1LjFBJ/iHLagsIOc3qYMuj5W
GKDuQAaPD0XPr56KuxMGVQtqZ64HehPZ4VC4bmkY9OCTFcmDrl4EbPuUONr+
RRJDZhvHe73kG/5X8ibElM3q9O4r4Q3+qOHTLDXEt2UM2MEGoySkC42miSao
yM7IYZHt8zs1isMfuZvor54EfIbz37LKdadn4uxznK5Z2l7H7NPhI51pvarA
SLn8rSoqztWqY5sCrx/D7BaUYssuGQrfU0/6GSK1usK97qaQiK1lKc5Rwu1U
Wdu3ODuLdz+XQGt1KwyquPPK6xJlJ2w9e1BTn+hdLT7EnR5F6EKI35HOR3EI
RooaEx4sVHlfvwQ/xXquygeuLH3S23HdUPtu0USEFnB3D+G3Q9z/1h06gX4b
2uFYgAfB8gXhYrhOOGpoRAOxRTMWOfejGTAcD063DxWG8ETnS/qQFYI7i5J5
TKTZW4vtnk2yv6AXvmpaGcs5cOaMNzLkB/QXkt7psOCdo7rzNUHG1ZFHi1dp
xPn1tvKb+qviqCvVWL5CYSbDhkp/29HcSjJeBuWhxnTQrxrq+/ddTzmiR58r
UifG8N6QBjQerXxfxgsftvt+9Xy8gSCgMxIP0OiCIRaV5DwaKj2dLbQFRqiY
1KCA+eTxb9TUOwmAHyppsb0ZigiXoc2ugrTuEUHmVxGJMCPskDP/CzjtMSzD
6A0HvhVRajGk7ai/GYFDRs+BVzTndnfQ/krTUdYuKkr3p5IZsMg9vjYraLRo
IZn1uSTCBGIF17UhOfglP3Gfm6fFyTcOm7lWb8TuOZzU80L4Y6YqYJ/q78Lb
AIsgbNHRNLesjZAiRuyWNRLYAT6Lq7hZ0RO38o/vkRQbmEm/xUJTIYSgk+y4
tc3aVg6FvIP6Xm9lktCKlwSoSCOCywylI+U+B4OQpHL4QQMhlXQzrm5/8sHn
ixSfkNVpAodOhyJMsaYb7TvEVnTbeNCPZaCLK8/LqW05f/dfBEbDnby8gJAz
aggPTsthSLt/KlT9YGLzPCnH2sIy4h7ne9odQbQN2r8GASVOECN1ThW3XwK9
k60I8k5pifAw9cTECKRTWRAO4qSUyDvAkZvXeK/ImwobEzTt4mCxZW5RRqpR
A8UI4eX9c4XV//BmQ6QIT14to4yHtUaPBninA9w/iS2JYm2DVPjDITQT5yJ/
cSbxGXo+BkHCl5bcHdF+kMv7YhB5Hb95ZkdV6znExTaPSLf2w/feNoYwqFKN
2NRJbvU9p4XHXg4MAiA5h1fx3zzkARjNlU+fkZ3bJ+x3cFAaTuIf4c82EGtx
YEFoWuLWxckVYCrzX7KmLrbcG3Kiy3xWK07D65CM4ITM7r4/bk47xRbmH7Bf
1pxKTl6IpLMhbxOF17uZ5kMo0+JX1DKKWi8QUp7qXjWeJJzxO0tImPn3QYsX
7B90Y4NYeu9khB/7/lmvO4iVw4WAoD1c0ZT4nwKhleUiOIO/tcVeaneuoZzf
aI1Mrs+wp3Qln8b03pgfcEtE1XRu1gQYNjGNoIZTPT6YmHtM2uVnS6FGVKLq
okytds9ThSv4AYbiuLGUddg8dRpN1AQiRmF5xs7irF+vU+nuCERQ0qZe5Ty1
5i2QkwR7SUBXf4g74PI/PNZe5n/P4oJLhsMoug8nboV8Sh9tlnHq2G3KBxfU
olGReoZHfSd/dEpQgDIZZyGHlU34mWmN0wPnMltkApYNJoYXR4P2bAnEN4M0
OBWucNFhMgtf7IoC7QXw89vK+NqyuB2kUSmZxA5t/SVe0r+mdUFPXw8zlDSR
f3+nJ1d9Axz0bIuctn2WMWhSxdF2NDqHdy2Cmy2bQtB5VLd1oBGKL0fYZwmf
2RVHWAN8nnGHzRu6pC+Mq7ODE+Md5283v2iiBjXNTmWLFhcrkNgpnFYLQZvb
NId3h+cOq5jqGpN1PwF0ZBSjNJtnp2XOQ7v6iIE2AuDRH3zWAlupDA2lxvGV
qk8qt0wEKRR0ckeWFyMo/1bK74f+yz7bJqF+xT0en+qdKv5OKJQfU6as2pqh
DUfGGtXcoGvE3ELxmMuHBR35JehDEd6F5+hWLOl0BenItwbn6L7yLJe47cN4
+9uNbN+l36EW3wGkaDQwz6Vb+ocEn9VzY35pmaRqoPysiV/vfRfeq70/QGnx
2Rlm9NdwjB1Q22JoThGQaBf79o4M5BM2UgSchRpOrZRINXesCs4crKK3dnMP
smNnsoSRxMLWSIoWkGdAmYiqKTX7Q4Dh4TiSVsiorwlbIXnRR2XTygUmJ1Wv
efzyBqhewh8vPOxC+SdVah7k5zi95JJSVF8bDIrP8ZJZ294eAr/X89CESXNa
MVlkNoMfP+JAUME0x60LKuTu+loKgjZxQ6QPFNtp9TFDUJlj5MIOUMPmHQZo
bRGn+R0NGQ8TaJM6iCTSLUyMlnTt29PrgZ5D03N2dItH6ppT5FM74ikyF10x
bc3orVbq9OnP4XcNprXqy1vUIPt95BybnwXiYyeDc76ufJCwuQh9wp6G6okz
o5EOotJrpc2gUy7YZQwHJNgczu+ygko2l+EbkKizHtJ98fpqynwb9cCPD4LE
3yDARRtcbcb2yKE4cpFGZRQBLsuieq0yyLFPLdOI4vPTmMMgGXhgdmgP0Efn
Cus9k47tcK071swxukEwJC6+afXHPwekVF/OgcqD1JoepTyRuJM2AFa37zc8
y1gOXSq1h8bE0wCV0LK2MKCbIUorUOe21rJL3Eiy2y9uBAOq/PVThDZXRsev
GBuZLOxEp/1j8kr2Lo/8ic5T2KocZ4mnIUCSKXxX9C6DdRdM8lbky9eyi0R5
zSDfugIfX+lNnpM7FdlWcoPjMiAWF73grw3AgHK7KweRflG0b3FINipHj14o
T4HFamwBE48QxPpIAvnO4iBJbn8emBYfVquhQvBQQjYSOrYlL3WREniAUYBu
P05Z9gLDG9hqT92VfPbCBGLmCr43L63x0x+rnKpCd3I4XZUM3o8dqHI7qZB6
ujYb3cYUppHosrPtefxuVKwBSUR+rGk/aPJLAkuxZtLg4MOUSLzo5t6x13bg
gT+OK84sRkgxSTB3tff5WPxJN2PcD//hk0nVwuHS2gyo+oSqjmPIUmX8cB1a
VpaTk5cfdNwlFuh8sFs5/EDquFbsapZbs4mJuAEqhElIdisBLLilo8c4hs6C
Te0RqeL1aJCpxFk6kctBznh8LdaCpF9CjvdXGeg9ORw0WOsLxl+xFvDdw68y
/4HafN0ZMPrj8QKI/8wDZ0Bgn4H/9mKxq0Vv2Rymn1pjN0l6l8SLOwCGGyLn
+0eXLsp+ZpU5owRgO9JjMeSGAhUGs6QoZ2xh1/LfKDU8ZxgNvwduyIlBAqv2
7pEoYKSy4EQOwpcA3hbGMGWQriYqFT0gcLR3irGctUT0qvJXSxkw1ZRF6c42
4wWsgCdY0LRnvtOwliaH2QHKx2iyNs7f8ipQrPTtoJpu1p7ohmDiyOZoiXOY
UfHSzdgnEKXvWNYFEwTRF+NK9XpMx8UvBW2IJwvwaaO/3bCT22WrmnOts0nL
04oUSBdpP/YRehfX0sea/iw1HbXr0kOW0xtBgkUbbznvAnotrquv32dUKLcg
zd3ZDI36VF3WFaNCOEFrDz9QumVskTzNSZtY2VeGau9WS6+CEmsnvB49I/H3
Yllu2e0z86ztW0rs1Krs6H4/Nz8meGvivjFjEuuzlKUOl+P+BE4hCmUp8Nph
Sb5HTzLf87XXgxsTNOc918rFBrwcar9VMh084Qa5b81xTmStd4qzLvHOLk3y
2Z9FY0giWYhK2sGoAn3RrDx00vtcPK/7JBZJ9l7WzBVx5Kz2fnDuXiVS2Rvt
CuYaVp9jowT/lE2Sfyok9q6/+eVzad/MwHI30Nk0kHtJU8FvJTetUEQefk4Z
niEHTzUonvQeUykX2m00Ug/Io1N3yPzEvFRoYNgXMa9rW7MlHKRl3pIYlEXt
WwASeXmd2VrS9J7gWC1JRlusoe0gdeSgWjy98iN65zzH8/cvgAo5NsDfh7ut
TkYmXh3zPI98RDDQIcFOLhUS8hvWY1a16MrIX0INMXNpdbzQ1IM+p2zFujeu
qlSu2jfj/20VYmpNGICh7HVA1X7iBeY+qsxXIpPRM9ayk1HXPgekYoH5in4S
sWJRnMfFl0+6KrXZ7+h8oOl5aDRe2+3TlXVP9gGHoSqFlolwkZKEgs31Nko1
DyozG11MC+4tfp2kIMZfl4Rl5eaoYqASJkB7mHe+q18AyYnIhNaXS/qbXv3V
idB6FBaioDbOzD6BQqOwzns9+oby1/XQPvCcm8TkfYuprcJyfOMg2NwaCrT1
o9YJPuGPiZPH3vC19o40z6GRh8VTUQgfQH/XbvPb4L0S6EvbqpUXrql0H+w2
XyqsWc4Tp479ier+eElQa2fiLf1gmHhdAqRyy5BePqCuxbEo0LxVCk00KKxF
MMqTlYpr8FaAV6srB/tuLUfURiMbLkl/evE/PfiAn/mAuYhwBEre1F9BbAxq
wsjUKGLpFVwenkUvgdoxmdEDcrUbMkVtGKXFvwA/7PIBwKiF8Zw1qDKszlZ+
k+mz+LFDNSsvSfpUk68hUrQKwKi/uRbsLYfWEH4xp8UgmIHiw2V7vafDEqQD
mwZliUPDgHMFj+4RONMtrgtXcOYGDLUtqt+mTCqJpLmi0d+FY8Fcko1+m4Lj
jmwMG7ira2vVcvz8keSt+S/2heNAyZMiUZleXI7v355zv76WvuqFzU2/KtWc
9CTXDuKHAhp7aC1FcGrzlYGoku2Vda0jl8mAZfhg8/++nlwAtD2mHtmJftcX
tZQXZJpQOY868us12KvdN7VQDE9dbAbfhbyUBiQTyBINpw2E+6gksxS/bqht
VYl3VeKqsiiYso3rbWSi0Mrovno67GyR0dUFZOQy2upven1gCTJ532BDV/I+
9a80k+mcmnrFNXHYq7BvpwtNGAIIfHUWo42O9o9+ExpJ2oFnjluJCPZn1Hip
Khz+fDHSl0EsjAS8YY48GTrGCbzjwDrJtAFhbHsM72Q6LvCTC3JE5chXJOBE
Lqo29I8vGxrPP3DHnu6si2VW0VZakJnvAe3wxqJETUhDlH4WLp+K7m70mpOs
qdJyZ9VEqaWbjTNOjs36lIrkCPNtplY7AjhA0lIo8qEQRPsRTBnnbOZ04Ls9
ZAg9WsAwlz0XmIqgLEkmsgeT9rUZdft9nYLCPeFjmQZKWkZraFhx1qlqyIFM
TZyU+KingKCslX6Jd0Vrp08mZwWNgDM8EI8WvgIuvbhe+fgkn4nzCazGavJD
Zlh0JrCqWlH5fopkdKrT7bNOMvF4MSx9Ymh5flkT4oRE4AqRU3ltZqzy5Ul1
UNvJ1k/9X3Mw5GYE5lnmJ2izdavGyQWkLFyNz/FWJOBkZ1wrIhBQBwVgGu/o
yRCODNK5Qmxzlh6lGA6hLzLdR+U83ZPJrxOml16HOuQQIQzyz0BeTfqXsv5m
vOTELKhAQLA0kuCOKUYi84bxbSsaU/M2yPa6PGXWyk6yHCsxpHT+NBGNr/l/
hosDHImTCZ+MaDutGq+7eroFG0+yC0XNm6NAupoetjbxHSxCaYWKWqKg5TDO
Gp27uuPCDl282YnH7dG20rvWkqixNydQ+0hZf2m81B11zn1z4N1M+3X6NBxg
UDxZ4u5A43uKsgRXCGzEEFGz87kszv+dcSQsJloRFgI7NK4hfLhHZ09cJQzB
YiQRdzt0BI/LsdEdRrH5Q8PhWQCOM1V1hlx2jg8eyaDyrxfuf+FyJyKFLsTI
NpyJBcCRnXV3aUXGQbtFECIdfGZPVhVejksef+oQcQyJjjPTya8BBgn/8Dlt
b5kI2yiPU1yzx61z3WUzp36VNAfTfgzvvoHmIGzUeFcsnZR5T0TQx44eqYR5
uTraKfy1vIsjJZt0Ph7lKkjRVBO0ug137aQI7BnXa7n/E8cWN88kMEZ3fxnT
TbvNOv7BmRprmQnaiVpifu0YBN6VUDbCxFWsBdw6+Ggp7ILnl7zimlgGLzqi
4X6ug1Ya8D5RG5Cg/GSofR+cNPnHf1Uz115MP6924HbFmOvgL67wX3BLC9Sq
MzjNJd3v1w6NooQhLiqYDMmANtF6vNhVwaGZZ0RjlvYKwmEp6WL7uUzYy+7N
o9XguD/AQS9xu+GDN4VWDWjdyjQiUjAuYZt2IoZLYSzVdINzXfz66Xi+P+ko
yQ5NiS4dLLA1BQsKyoO445qQ5rNRdr4qR3ho2u17NhHA6awP/0gPXyWR5oAs
TN2twl67EkkF468O0R++LcvVoNFYnz3xC/f76v1hncX7SnFf1ZBRB98YMTzk
SjJCXUZVZOflFvu3j9yMOuUfj56XmcVJZ7iRvPGEG00H0ZnjG/+/qnM2uStR
Gb3l1JnVcM+bjUratwyuE5Lwzw0Hu7W1aU2+ugRKzVhfHbaCQZCd+kGBG51y
bwtLdorUTe2CrxtcKSmskDdeHPxJhHU/lnIv2BxheTTdvnGxVHxLLBPVs8sQ
6Khrk8O8i+EQYQESRWSUS9SldpYi14D4Jyc0Sou4i7hyIZeW9BAA0FVcSpLw
7dtvi44yCT52+DZ2okBWCISoHzERAnoWAwE/wwtxbgqHJozT34HXPFZHNarv
LZxaBAaE0wSOfi9WpQO+21vrccuTJ0ifj3jE3rkmKIWs/wFiQ120RN+GW6E0
849M5SqtFGoPkpF7ESgx1hTihxAUx+c8eIjSQU+PEXHGIhu+OX4EOjA2ZVAH
Xpgg1/FOVQXcGQLQl7wzU/MZIXi9h39OF8BT8omTQKNDRuqGje93nWvLTNMy
i0PpE2B7GUJ8xhFairtk1tHXWs1bRbS46bMWqmlNl9ra81baiCsplKvoc1iq
COaMTNlgfG7sg2b3rt6SGAM+Y3L5MyLH5Qci68KryQXxmqc0zXQnuziBZAju
/IKC0pYyFJzbry0SfAw5SdzpVB7POpBtCX4OuJvd4s0nEOo2xEO6RFBHKmUF
O6bbU6CgeZLD1zYm0HUiB04Iii4kLtIqc0M4qYlszzajPgQL2tsK/8hUXJUo
eImqJrP6mmuAH5Ah+teVUsQoOnLCFNA5CwIn2Dcord2loI/n1IzAXvzJ0SXT
pnrc8tuhRBTwcccx869gMDj/4UOfaDczL7u+CBKqM0S/WCiub+q49g59Cgua
j4gsuyDR4gSXuRq1ux1aBRVOhhkv9RyBbjHe3mHzey46X1uWNloI6Ygz5iML
D7BBC2GcFE2qO/OHqTovNUIwEqtusYw1TNSSeAhFDPNY0dT2Txy2q2Imw8kD
QPV4Pl82YQRQcPqJaYiHh1pzX7c/Xk34vPLXtiT8m0NTnLqWE5QHnxYfRJmo
jKl67Xq2a+MOwvLEcSr3fIVs3cjV8W1RXJKLhZJNRqAt9nRoGDbhLsulD2D7
pDUPcrthLd3m9Jcp9GnRonyh5EHjsSAq6NBdIq/xjnL4xSMlotnKKBhAQQpZ
Wpozpf9CKET1Li8Ahgp+pdJ+5VmTYtoqSyLfB3O1gOPEDlXl0qCxDvNcUti4
wwLKBC89qU6e5A422pa+A+CtoKpTVDB18pKFFBRsotF8NvPhjJeWtsWzIzOR
bqOhYxYpkpLGAkAoK2+UmCuDFU5QVQa2tsVheQ8rLM5qGoYfrbp5QBRWtkli
GuI755oCDp4eNf4SH1aH69l4cKJtBke535mkhsQwd9B0EPO6hPnuxzx3YaBQ
7nKBC7//YRKHZXGe+s2koqyyjRbx9dPbt2DsTGZoPo+EF0ypt9Ve8NSSwdxh
azn8DANGhymu6Y1BgZr6r9cf8AQrZutlV0F6GUNKH3c1FO9OyYtUeGTqaH4F
VjDyKAobMOaBwHmgTDaLuBcYUOpR2DRtx1QR4l0dXYrY62I5nWeD6udewN7q
wEHnUFK5i+gu9iG5rNjfha3BVf1EX0A0HBXntWxiTT7+YG8rJOylfh9KuCJB
bb71nJuEul4YAaKfYuVnzDWtiF1NoAWLS+nc9ibvJfhA96ugRRfRQqevpWRr
T5vI2otzKzaO5nFFM3TjNsyvCXcHtA0W+X+/odKiYOtDEeom+KiJJWCjSpRv
ZdMt2JbVC+eOn7TJRQZP+MvlpGNl7ta1PV1cdBXPOvrsTCFaXWWpBTpcvROh
uLDyQh8eomrh0W7Vr76pU0JOVGKEvmBeP+uCO6N8Xb8wY+PKWyxbjT+MR/y+
WeM9QFBpbk3ZRl67Q2c0J5f+eyhKZ2uLwT63Jxe1peCIGK66PVsdI0STuwIf
2qtMcW1iAYrvd96hEu/cpaHx13FhwqWfB4At1+jbS+137TJty08ntD9TzCAO
k3AYdGU+6nth5vayQ/1PTFOFTcn4O/iLCIWHRUiaphlGVMy6h2xaeHOmJtDW
//egbMniJ6l03I+QSDV+J1ZA68sBh/fdy8DkByBa8n1MDhrPBnWxzbeU1gVT
e8WiwUX40ntHn9vIw3LVZzij9teIHcFG092z2gVl+T9C2zE8Y0PhvAR6nOhn
/ceiqunoGSHC6E0cjSOl8ddlxehZJ0LkiEHvkl5sdyx6VXbzITKmkGFdto5Z
zHkrPVPOrdUrEbezY3cS3JlyfsPK28Qj2pjEB7/Gj7VDxcG2VrP99nNwyiow
6ggHrmwOPiWip+rEvB5xnIkcglw0QzLd4daTeawNlft1fmkz58Z7fsr7DmuO
QN7m5bJNgRU+0/xtFuMKlD9vIboKuRdrVRJ7zs1H4pGA44bBWh4BQU4lQJBv
X5FxmJ23rbXVzajcolOU6rOOIvCKKHDKPyyXcBf1VCLZt2Y2qpgtREOAQ5dC
L+3C5YJ3v/GlCfnu9jd1rsh36d0M7Lw7olv+V8H2WnFOlOl2WfMVKlH+lYfO
GwMvXihbQNxF4OTZuGHnCKhXGTG0C2wG5F+pBUKsNLq9Wl/hbu28G46A91l2
dyVDyPJci7R2iUFEsYtRH3OIrweVNNk27aUIrCy46eF+/6rbalAKQoVbY/yb
sgzeKBC17PDtUzRxP63vZBVCGpwwUUlJJsYhoPA85peOBMQRdR2JhSt+6I6X
Ukw41+YmfFqpFE8j4pcfG8616LFy7Kcs59hfITqzGIPfY0rbWMRXt6BVFGnM
sCCZDkGX0Vik14juQVOfjdOG+nxoNXkYaYZZIYUKfjQj0Ox9rm7Y5JEmVJG/
bmCnGf7SkPS2yDrQ0P+D3/jixaLjdNbhdsf+8Njxar9m8bv3TTtF9pYa0K2x
eFqvZp30vFcAV1dndVRv+5gicETHpBzfl1J56XOixU8cHUYWLq8prHB2DPyj
TY4RR5+sjqX6MIj/SvDAgsqLvb6blbEHHas35vZfsRGD3MnEK7wMnABXqK/r
6pqN1XMFKnVcl8y7LEebDdJDgw7tqccY7kocDxn3XRiE3ycnDZQs576830ip
HNjZkl1+D2DJyvccyx6oRHQJ+BaF5MVW5ziFJ/pkpr9WOgOU2VBs8Xqk7Mp+
nfDTGLcel65zwyBuMQsIG64IS7mAZjyH41WoVlKCZVqAFBf585kXjKe2mLtt
WD23sVS5XSsdMmNeIkOvMo73aQYCREC/+iLOZkW1xc9+N1ZbpplArbVjfSCk
qHFgKJDMXB53BP6zPcTzkZgI+o79pojycVi3aBeAbYc9lP978I7iaGqUXs7I
4pMPepb0w/NOOMuh9e9tPi9eUJi2k2EkCV4OYoIWfNCB+uS5yV2kI+wqx2R5
K110bKzlwFsSm0LKh8eXT5YA8Taro1j5hPTLgUq9MjEUR12Wbz5i4hZwkJ0j
EIRJRlPQ72Uj7b7EkKT3jvPDW1KHO4ic/eBBq2M+iaB/ZrCIGVGZQGIulIIl
KZNytBjV5BQv+bRxYmPw3IF/MTrsM0d8orQcLp1HsyWz8MQjQBkM5w66gzl9
G/CjxoDQueUTfN1EOrefcx0n209tlsLEkryu/gtEENepFRJrBnzCoUh/q1DA
wq5Y+i3cfKf7ljhcIk476jIRneu2M93F9mYofrvKp2+l+JTeWYm6La21/3EJ
ui1WgBv/QM3onYX4WG+/WEXlkue4HfA9nvhd79kHtO3Qc9ApNcxFZaf0dKxf
Mu5PsILfIuxD36a2FbgjIdB6qPJ5cou1hb9i/cSoA1N4r5K43Sg6tYE6PP96
yNYt0I5IEvB/TzIk7EeESpXff7V0gR7MXdhFlxAVgm6IdTbRw+fR4jVBCdKO
hs7kqejxE0i6Gi+rmxQ2JhJNHsrGJBzIoaf/AbISklzE52VcQqjFMMHSZRrX
wQd6Aov0rPwKNUbTnrjQcLjnTHMR2y6j7aOhCEbCNDdSwrN0c/3fd9hSt4Of
/pjije2uLwioOIU6u5iikUlu3XZ8SOJn0WSZPiM8lJVcLlvonqzsFQUYey9c
6ExDQZ7yjgYFv6qUFzExBi5/UiuLVPwoUt1oPRvpIxCiYSFeByWT9/wyj6/1
wj5ZxDbG1LcQgNm0gCS3cN8tFzvjrY2ZvBYeM+RCNljfyB4BmOKkfMcFCTXo
VSqEK3KeJmlQYMdayYcCWcQTMYhIwwDAiyfwrfrqzBksSbEbibytflNt4fbm
aN2UyZ61hfe13s8lZV3bPPvZBOPK6URADvirX/zgQ6Aw5D2NGAdTkiHlWwia
nkp84GHWkpy5r4br/k6uj9A9gg1eJEwpjIKr1jElwpAZVJPTMFpsr5omvQ/l
3fHeSLwVOzOrBdUzdupNGuDDxdQtyhxzdBR6hkYYU3WXgsSZb8FJHtThP7lR
1iqZPHJh1s8ydJaUOk0IMdcJg0fPhy/LfzcWRykaCm13YizwWA7/OeaDkSoF
eUgxuSBxAdQ5H7uDTNtSoN0babKQ3lyf2yfFbsDttM71a2AV/l2JWHXD1qUI
H8oCsZQoZPr/sAhn9Aym14PnCkQiwFcsaM24XdOFPmv7v+4YYqA91jZTSpJW
yKdUFV1yfhjce14SC9MwXhKXtJhnKHrjeg6spcRJ2ff+jCQecrmhnkWf+QMq
ruXH20OATdHzdaz2zPdXB9MSRi3ChUgtJ8xQFp2L9hdNCPlG7ePTayMsG87v
GfLVQ96nxNHRFd6TBy7SJqivFVUMSi0tGNi5We5wcfsWFsq2fiyoErZKagho
ZojdVWEiVAnecr68Mp1rRe0TAtD5T6sFd1VSuzJwWydP58oo6bqhx1AlK9wy
BvDfIOKFNtMZ+W46AYRX2ZxaKpnXHBskVqcKCnJy04OIV9GoT9PWamwM4JLI
n1w/PdmH5JHkiZ2f8hf9X2TaenfQnY/aOVKlsX/kzPifqrAXH3OjXCxG2Aer
3QsijkWwI+UOdwdF98Mb6d2iXxGzxvhiYCy58z94EZX9WicknCHlCwF5Krd6
6+YVPtiFHbvtmQyCp/2FsOuG/3+UH3V8BeHi71ow/7H9L+mPRMDjajkfOMN1
1PK3rzBmoMopYPqhf6lT2m5p0aPf4QkD/6V/KGVneCpC+K1FVO2qmmnm3jur
uoL/2vsDyQKXelwULzLlRzTlZN1ewR52nB//t1qRCBT8hXsXS8uOqjjNd9pI
VIknaavgy0IM8eLjd5OumP6sL0OFchIOHOVB/hCTh2x/VsAtCKnTZtK9X1FO
tU98twYBJ8oyq33l6iNGEJFM/xmTkj4vjvrgfsyWuveh2ItPjXm649MYYPU1
MatYG5jE+NI8gdClzBt0v3aaIxcooZAYjTxQDNJgts/ii+kNIrnjBG0X1SUc
Wz4jzTooP23FuXOmA8e+R7Ujg03tQWvJSQJWG5N+vCIl2Vcr4/ULLiTbwTUl
URC9Zvru8QY9Pm5Jfgd4Tw1jcE4/ztjCT4CuwX9TBAabsJVUQnAma+mzHfeF
MxzxXV4SDwPw64VHHpnrc68xX1EZxffokgfzIi21e/s37wMDyEpgixRJvXtV
ZXNesqjoCOloZ2agjrgkLgOsEd+z8DMAHrpmQxYE7k6xg9sthG3lgCPuRIHm
8p60s+putZtPp9/ghD7ghjCT7whd1iPbNKaHNBq0dcJBppt1MS0kQSAY8jCz
g2ziPqH2RupRvBLjhRDtDY5CJ4v5LCoVx7BpaCZRJwT2S/1oN9PiHLUwDGet
Srt42cS3V0ST5gLsaKW1w/WKdjTNMq9GmFqp1ovrc8ac9TBLSTGL1z2GlZnp
0GN13lV95srHphcltO19HoWVfLcn/VscGK1OfIbG/7NfFL43dr91Sl5+5tyU
SHAClYGj/XPUyU5krVKdOs/92EDLfpSyFzQES6dbXWxj2+QKUMK9u0AwC9rc
Xw/rOQnp9y1kWWQ0HMe3qf0X5Y5ZCtZ3QZYhNACoXlPSgeSUR33VDhptWiaM
PUyWlV4EiKJOD+54i920/1hTNpsj8zCVkUalnSlecnyNGJp3YVc/37Ouyctz
yK5qiuKwr8nqGDCDp2SIb5inHEwCZggLSdeMLGOy0E8Qg+y4ReBismncFvfA
c52ObDhPwQmHd8Vab3fd72Iju2Bisw1Kex+mRci+2zJp4iZXQJCFlxHxd/KV
/AEmmRJgr+njn9DAl8xC4KlfL4xqwFK+uvh/fvsdjzCOlHlsiY/oguseIoDn
OmPKPpoFueAogDKm/+aXhJqJ6jRSxXRq5eIo7qN5BSoYftdUYN/Tk+Opcevs
AJOPAwaFUJG1gkMdZkYxiyc6Cdt56xNRAo11OSI2+bjKMKcMHZve9sQLM+pj
8ERUu1cDcK/huS8tcsXZGqaIhxQG79UM2a/7ZAhlTJomwsSiS83o3IlkUYpa
/xlTrFt03UzVlt/LMOOfYTquS30W1cJAtweH/JZ3LL4JARqBjIPO/KU/6/Ze
M8uOCWOC3bXMVNmvOfRxiM1lZh9IhXbGDLkU44E0SGBOvJZJ+Mu6fMGtYn+2
7vLiAy+8jKed4KQj+e9iH8jqYfEQ8fqgZRtGmtMUly3UabFXmEMHwqh0Zjnp
k8Qqx/SyOnK1sQUjukFGLOaGl14rKXYiBZNBZHWKJmXGZWhHuZYwodsS+ctU
1KU2QK28C2vlgvQ/H0vHFNli9OVtpk5L5fSqcUY+WjNMohC+UdvEtp7sLf5U
c/MCmoB3c5MFdsS/T5byAKcIQeXtUOw4wUAEiExgCDS+76vLid4Kkr+SI+Lq
szmJSbSECzytW50ktoXGMf0DUFeVc+zKXhaHaW4VAE2CgeBU2KSVrOc99zrp
h/eG5nbNdg1a8X04Jdf66IktX6nVqMryKVgjv4UAp9OuiaGXh6oleiP4YX+a
xkk5FPYPRY6GiKtdtK+QueL+tNHjDgUx3rUeMruGfN9BGxOld4w7z1d6O1RB
jJKAm3C23ssWq5GooiO/21qAyrGznwotHbdUtt2qo8to5l4afu/4Oc3Nus82
rBmqsBmuaZKbnU7Egv7WAQvqJlBaXtGVMirJM2sPdArujz7yQTAkt02CSc7p
2/MP32iZqp582hX92uuGQO3gkwkvIlfsr5dM9EiYMjJpHwDooZjnv4UGq6uG
WeRFWVsWT+uSqCpQ23gjo1e2AoQguH7qwkZwlTW5yxYTgfpbH8uBwKvFGl1F
zhwSLcZwrl4egenFhXbWds8fT7mjE4/xVMyo2zXezGWfpSI7/mm3SJhXgBH0
/rzwojU1eXPB0P9UOnCJpmbWfK8gt297HXUkIp1wKP01SyyZKXUVdOMFSIOP
k+l0NHVRA+b152NPbOY/NktMq+RNsVERRssO5evLoZ6VScxxQnpT1eEOx33k
w5u9pKQVQwWCyDyUPBohbc9v/dUCXiRM34ODV5NIOYenSHUw28TCw1vx5GT+
sFW82Su+xyKrxayznjQRTXgFdN6Wa+wU6VBDUQCbzWsSMcaVY8N38gMDvRWS
2RJxnnuf+63pGHfJh86hQ4L+Gd2O/c/Wa05Y4zjBHfX7LdX7+tBuVivTa+yb
KjbMfgCJwFeyFEwmaQKUpbyyLGAKQmDVh2cvCabuGZnRGd+mziBQ6D7CyTej
Wi/QskRddJtcXMfLSMqaeHheGj5usv/RHh+eusAqQXQLV5umKiOnMzJoWEqj
5NWkiVoVRv8Rg5VdG+7CAU+cOka5PVCj70eat6wmVxoa8Gu02Tv9xbCRt5x5
RSMeA2v8g4Y2DwWaIXGWEprES3E8GTEBwzjHuXeRo5U+0O5C8qXd16euucJI
wpkyn1jyFwEe1tZ0mE/SC4vJzPO/6bzus4Pc8/SgkHplNbwLumJ6TopMksii
nMGip3niwfcvdiiWz7wtMjOmzWsIXdei/7N45JRRIIcpyu3xCozNeBsBx/SY
m2TjqTy30xTcWx+T8UX4EFO7kGNGVfyc1cD2PvvvsjWUfEGOTTFMXWQL4HCw
KOAmOewnxZCuihzkCy2OE9Z/uFSSYNBDZWElhh534nI3bl0Lr0GgsymTVFOZ
RMeqGgxFpvBOyysPgx7b8uhLum1kjlvfDAG+0rseQ5QyOCJMPpQ0i2quZSz6
PPEpqIjdVDaJo24iseDGAzYTb8lstiGU9eoc61ZGQlg9PZyL1Z3A/vKSM37t
DD7YQcVisRZebq8cTQu7Zh1XJnYew8ITYRgWn9Cu+HsQHClu/frIiu/SVYbZ
Y8rilQoiZkXsnShw3MffGPgBcty0xHjgsrJb5NLjHlOSLaOTcwzG4qPvGMAt
l1vJL2c+upZ4O1vqff02l35dsmAoM61XZVsrSXlR9uWdwrx1Mi2XFvV2IZae
5wbLA7ep7PHqnLtRX3nQ36Z778YPA55gdufw3UAFiNCbXqObB5QaUssP0oti
s0WJGtaoitb6ISPtaANg2a30vvKCtG2xqv0TMfaZkAZvsAYS1viGbSdA83nA
iKSNZK/MtnCQyeNiorHRHvKIg6EpGiRlDIMND3+/pDD3//aHBBmG7Biro7t3
tAY0O7f0FfgczEXuS5G5wX1fGGDNZNUQ75jgCu8mt5XhOD6xYHVmhTTUrOAI
5YpTVKtdzTu5aIp1Wb6I0fLtdoi0DeDeZ/xpqmE8mFuq5LJXhISYg5F9STe5
fAHZn6jSNM530GuL9MYife5ivTGq5gnoaNCXJymsflswZ7AdCahzzPC9vNZg
3ofQ7WwTFVJpdcgWRKGMv5kmGDQmR30HCB8PCZdk+txRtLReeatYHga2/JCJ
p8ZyZFezAVcwl0ebEcp4Ap48kbv+jN7gV0iHM4tKqnTSLY1BYGHHkEvXcSTt
/M2VkahxFCgOdkE7eWrgX1u2iLM7aclgzbspY0QXlrMNJlpWko2JSxKgaVRd
xEtX0nXSYWfWNTjKMQ3E5YVmyRy4T0tSgOn124XyXyMHTJdWdbtztUKkEPM6
ZpaDJPqDpDmrOvuqlTQeXnZgViO0QUPQ66JKjKIQY1GgPItaszVByo1MJIo2
67Mredjb6BxbQaVibfq2nyLGWZjcnalQj5nZgLEbtxwIpCSyk7B+Jm35OZbB
Kv0mrUAk/LEF0ykvsZpj7bJjCxkeKEoQJW8HHmbc91bXxTARpwt/JhCqJ3EY
oRsZchZRsK4TT0I1UmpV/S62XW4kT6tSLi3jREZKUolDca8iUHfWf0qQLYV+
IDQQkZ9VuPsTJ82hCh37bVsSq61aQ4KBRSG/FQ5dSh+1ZdsrGfug8X1cfpG5
mWyMeAv0P7aEyhKK/C41dFd4U6tZKEJuaM10PoZJ81ZYcWd0oMvTAAwboVia
KvrN0K1mPHiKowQ8LD+F6ugc9mIPim2/2zHwC3tJ3ai6EBQPAEsZTXlRF4au
xlsiImQgEoVpfOkElg8+48FE9MVmztSwrYyVDzpndnNyQ3hPZ4e7bJh9vPgB
6z1xyEj1UWL2+FXKCzf5v1F/lgz1Xko0hkWU26H056r5GEBAQwCSjL5dpPws
Wzoi39+bb3PN9fiS2bYxQqJ1JyoLtcgTDigYMvfXPXrBed1X8Y2dhzFnB+pc
Y1Hotu6lCzAv3U/jFqWcVz3BOSxidIeRShnAFwj3oBsJFeXuV/EHehFdsJVk
WOB7GNiVE/WhCYyxSrvyqEustxCIFPhOwwMy6ryASCegAL6RGTX5L4GYesNt
GAM47hfrXT72miaapDM7Ff+CyT7DViX1oc1+z0D5kOFtW2yH121pQxLDmYxA
CWgKUlmDOPO3nfXgYjxJxrEfCsiepz83tDpgQOvbPuE2W89MpEf8Uafu82vF
L64MuqgBWZZHs0kVOMegPI6pyiTfwgSrQSfTh2P1mXRl7opHIodaTm8AnVir
zSk1paIsEg2xY3gNaq8x+cKeKusnf6TAt1ES6jbprxGYbLgF7x5X9Tk6bO1R
vEKQ/Fto8d9i3rnQyFrI25vlmC+kef1kYTOr1Hou0QgnvFUKTMi3sfOtW2Oq
4lPoW9nCvV3qeP0MzIe7GhRDNyVeIHzyJ5fJUO/s36WY3j0LjOqPEIBzMPf4
Du6Tqttu78/efdwC+Hh9gDZqiULp09z46w3Afja9YpNIrFKcAt1nqhbf2f1j
wggg3h38T+wHR2srB2bmPin918e2UFAUULcWkl8zqX7OuX6fojgSJ+85JcxC
aV2dt9H1IYo2Hm7f1XsANGX/lmR3q+cC5/ElWdJ0VMFjFsuMvlOg/pDplzEB
wZLjVRryVdc1qGQCDi4Rvkr2kD2MgsduifJBH3SFBMna6glFhqSNXC81+gft
tidLVyj1RwuVTutcjrnc542MidLk4ykze43iYhLPSem21JpCbwcw2v3tHTwc
RU5y9zwrConAR3RgssH2Gt+jo1HCg1n/mqJQr9kzrmx4o5vDbgsBwM/UkU3+
0ryax8Ne9XcqpIeO6cd6dkD0nQALJr/r73qbtBT/ZfbggQ6NN9C5G3Lgrg1L
5Ns/qa8YAMXJQI2XC61HQQstXK9Wwyh4/MqwLyi1kVTCsQXyut6W0QZ3vDC3
XaEUTxbtYJn96tMM+AFdV+r5ogE2CmLFXW++P7Kpi7cQfGQjlStt+JQe0HCl
3VHOYHfqc9h2qIJzafKqLst4E7Ylz1RguDWFBCMyKyV/1wVQGpASQUTYx4Nm
z7b7rCyrlkIbugvjOSL9mpxViyNXXWiUj7zmxh7eTy42t0DkCAmC6MaolRfz
xV9txzQtvFIJU4QijUOlgPOpNrwvSC5Nd4S+YGbmATw2IOD2iyPx2H04jd0I
5nPej8xw85Kepv40ndnuKmjnup8zkJHQwt/OvFxEpZxCkOsPv2fEyJTGMvt+
2BZLLlmdQDt2nPEouFR28CH3Nfwsd63XnkrAIxi11W2zu5NM+E4rfKs23+qj
hVQy15EeNrjYGId7EDMTVJPhTV5xa1yNSEKkqkYeVTDfFB3W6G3SRhjs+b1I
Wq/RzKIRtrT+umxDi+nVDwNKfKyOrBHTU0dbxfA/x8W2Yl41kmm87GHsPrBG
f/kT99YN9+7H4mqWHgksHuqjoQaoqHDxtedc2Uk9O8V34iEy5QiMLI0O7yxy
PVqdB0NSN9f9aunWM9sPACNfZ23ZXTTMiWbRdgu20ap39aBflmii52j6vKfj
bVOTRk7w/Z+E0jo560KNoYl9Ucc/OmbecaSYcwzOhlx1x//ced/cGYlyNSoZ
iVj/d3DHaAH7NSIUnaj3MSHuPybAofEp8l+GakE+wIN+YOOnNZ9ZzykKEvgj
pTL41eFW7mTyi9uIn+By+jneKhMNH1nudxnlztMcYufN2yHrcwa8w1dpi6Ce
f0w+8fmSEmcckpM8SSgKu53wsNYWkGdXE2zv68+4z1uYmRm3EHMRlPKrvegP
0w9hBa4GWTaxDLSxgGwuAxG5xi2NBiUwRr3ovtXTuDQChuw/jMfAtLeIB9gX
GoA+aPZpomfuvaTLl+wKsUDwN5LXVuM7YrNCb1tkv71JqcTlC+7yk1R+N59t
r3Muwmi9z9j/OZmvO2lc+70RJetIlO6D5JQMvtKKRrLxVXNW2KtY/iucwNKN
sk80n5mNIJU3/VMfdmtCag6K9C+YBwI5rJsoZstyZx7NaFvoz4t8PdLi/Gfu
WOxaZDh3fJOAgYTgQx9s5aw49anBpTYUDnRJ7AQ/XgKLvzOiLQPIBKWqf//L
s9tqbB/03neRR/+jgXVt71nJViNl8Xyf4fosGgzvA0jy2DFcJCAILrv4+udE
2s6p0vpM11afm2B3mMFWkF6afiTI1E611xR02iala8CYSGPUBE+dVWTV5HBE
6/U/HV0VBLLmuZRC+JOMo9jJjWV4MZ+utb75BAR99oiqq+65Uq8izg9OQbqW
yqBZmF7GBioVrSuHQMHOJT/CWA53yEMFAjl97kTTnjFsOuknUzg/VUKjd3b7
GdyFqXr89OYTERkg+vbqH93FO0hjglPiAdH01KixuaVH8vcFp1hG5RhDtVsS
HG7TWZ6k4fB10JOi/V/EtbwmjdaV2OV1Cz3RbfIhJters3jw87BBSfIFHzZy
qqGOAVKHsLyuaROSKuBgRAkBizLKL8Qpcgjs2HcovN7E1ukw1ABBwVJi3KUU
6ias/QmOWVJY03Eaay6feZb4cN8GmbmB9y5IgpA8xQetbsrnMz1Xw0iNvz4i
xij0wxlUBUJDoASJuE2j5vkM9DRO4F/gD0tJ5SQJD9FwNv7L23e6LeNfY80Y
HK//30zGlF6afKJw6q0lYEGgRPUmFymnSoRJGkOo9OPrRag9wjPnfCgVG4gG
5nyg+CEbMKAd31pgwIf3NC5xu/VoziRX9d7JbtuqGIxq+oCFYbJ7v5gV6vHg
LL1oiJQjaUh17BiKG/DUqBzbYtSyZwkwSNlgGXGIa3aM3Bi0C6dBj12m2RCW
R4lT3djX7B//W3IJ7uYooBD2yHGRw2dz14z3E4UA+0I7b1Fgg5ew5bT54eCR
44uFrwVys24BTPcLVpU+bYFWtdz7rY4t6NMAG9y7aiyfgeAUMrT/zt9pPj2f
O+9jVxY0d7pH6OSJ3D5diXNowtrojp8EKkflXhos38ytw4qa8ciTSsupxXhU
wxDNKo+sLpFhccdHQQXvlQ5SfYj1Ois807e2wqNFIQmIKJcynzCZD5ijVsYa
T5K90ExgqfwHAKsvvn6T+hses6Fj69qYXVq1xX2kK9Fc2K1vvYSESbQmwi5N
EZkHh3ZTYsCnf2Kft13zj/hsPYC5dCIsaHW44/JgIunMmjzYrtJwEDEc3CuL
sKA1cl2048pqjSP0xEU5FEmwUaKZrxRmExaRvCmaoMHIrOiESdKVbF/wKYnf
S5ias3q6YB5SBhSghn2MZ98knJ3kw8si7Ggl6QjB3kvP0XiiABRiKk5IuSg7
8yp0n6gQ1LlR7IF1ZVl05EtpFlxpvvdTV9LTXqRWKx9pdMrn6SuIzz8gJrfL
iviPsHmcd4vNbpgfOOijGDVry11tuShmNl5i++fsOYc4Y7M65yl52jH3R88D
0pUvgBU3yK0HpQW8Z3lXfNroisWjuRoccMvg1rJqu7Mw5f6HeENeU8tnbt//
Mk9sQdpEA9aNrq/eBW/p6wogn/nSztU8INaxgtKHDTrv68dSF9NRDys2HpJN
9aawhdIicLr6p0syTWWnbVl1911StRxvnXkGyzIRdtm1yZG+6AD+qouN7hCR
5aXmZVHJ6nuc8gyzsM8+Uua55ha8Jxp0dh0pB/Ujc98rlfYL1GL/GUs+ehhx
PgVKbDDt0K5lBJMZIJcS5TlFo1O1B2zM2HL73uBc9nRRpIm+1pkFGdeVC/k/
sB9HINhVG4vYOaTIzoALZWQUIOwkGi8VgKl5cF838Fxg038RImlGhQN3nZZC
MeKFEs0SbJ1cNNpXGDGy5XC856CxGADrsOW9s/n+0CrzqKzvzrg+MkXuFWpy
iQOXgujvsCshxwM5ooYIHmm8YdQGIvWAyG0NFRAQJoaLqWyPANLB3zXRYpa4
lfyXCt6lliyK4h9RGwyhevQ/pWEaxmGtk1jq9xJmKKhmCyhAbT41P4m88IgB
wlU77F+A1SBFGZyTVXiczG2/lJ8qGqNxjAkSBSpJ1ELvyak9juvLzwcziQ2r
cf0axDmbfV5FyJZhkl/Ag8mSqlXRInYszJ9w16xAVmzgpswvBNFgWdETy1EH
1raEwyH93xFtxzhviLGc/XEPxeRDqCJNKr2Je/YFkg//KCSKPrFxjpdmN/22
MWNkloaBrMASJLHPGlaRbq3ZfBqXLGlezXiWNSxn1SKxIWuil93mkoI9wjAb
cg9O7muQcZnvScCrlihN928VPfAvUmAxhrNu9UOW+dimf9ynMx4wAgcgNjVC
omzx/n6dRhSL87VzjYXvHTD1D1+oe/wRUjccRG1rzv3lhDConcQTW+cOe01R
n6lKAfWx6jW56tO1LOaVJy2I38UcQO1smYWenQHQNImoVDE/Rusq6o/iuWQ+
3eN96kJhxR43SUAeMgMc3IKjXnuiBXIBMuZebbddzszqR4pUiFPTmTLvhBBH
j4Zb24Oay9GVZLC1W115HPguhU51GuN+kk1IvNDeEPxkJT551C1EXsqgcMlD
rmA327+mScHznabzt4Rc0XA8201iG7rc0Lbr6oGt+Hyz4jcsR0cIOBIKVckw
udu1mScRt55A5ZEtht8ZbrAcHZ6Vir49K2HZaHaxrNA/VG4UXr/4FcdfsGMy
/7aykVCiZozwDunz6G0jVOgh7XVSQD4u5Y6Xgzr5YZuoVVzsfoSidI977jfa
6OZcxS0MkKtm2KpbhDz3thVmPvA08QRbFFoiR5tl5KhWKYpP9ktaTsmrFuQ6
t5gV85FvDgYDoQny1kmOwJWrckSYLlbdKhgUPmysN39/HvWNZ9pA54FDQYdh
z+6IquOWkfFGHHu8sdJCQHiJ57cH2jJwshwsVEkB5s6tekFAQ10+HtSadYJQ
5crE1aqHEB3WrSLQhcFm8NcJYKno36Qbd7G/I4Whr4DekZrryORZ0j1MhJel
jFaXmHgZVM1g7HI8jUdPY0/GvYNBHLh9eJtwOYz1pA46rzzSkQWquv4CTasy
Jl6itHWP3mJx5ra6dqboh54l7KlE2Xj789UWryvXkn7z7ymbI7H+zYyLycei
MbiOwhO7wbZsBv2yU2D42LPcsbDpHHuXG34FbWEAAkDrvnjM90QTLwA1srGj
FwgNFA0NZwEvGnAg5Ky8oF3oo1xGuYKdcdr9BzMoLWVWM8Lgd15bKfDnGUky
2ZudFjQkic8FZxQFRnDohQ7TsUt+mA7RO2jTCS1LDlmUlgUUQlGRwNUXbdmx
EXY95NBS1Ls7yeU7IUrfrVkamHgPOOAEzMmMPedm6tz+kzlcbPsXzDJkzult
OIlnRqIzKtCGRN4lEIrMlIemD88VwB4hvICflDIwDuzfnoKsIATLAz64pKWq
m/SUxzofifQIM3p3enr6ErmUhtlaQnxnk382sgqybktBV6rO5v5KGoPm51PX
48/qDicFtrTNV7V5iKNIKeEHOFJ4D2HSv4JqxHAoICPKEChUHdMTP0C1IX6L
4BI5M3iQ52UcNALyDBX9VMtAbIQk65wpEtpuRkfepeeB+9N3wlGac1gRA1AB
6R/B8Vsu6wumM+1HjQBKbblSU+e4jvi6bWTVLVFdTIPBWyl12VnfeQbfZW7F
HiurtQzip0pJEvYJv7ENX64mVw98cDfvwT3HrEx4hj6YAtKg5LR2lY2+rhOr
O6nYqRxXfMvf/nrBx3/SrsMBCYQoWE/kbhF4JlVxNHmQcxQhhw4oSislH8xE
Tyoxbcp3OYcPFGKiPNC2fIj9M6q/tmF2fLdFP6tc4MpEWt/NIsJXzWpAlbz5
iGfZRLq35Rv4q+NDAsrehhWh9Ckill5XJ2my1MPdabA2pbx/1UO/pdPGAOCG
30w8l2ZaOLk1zXKPiqZ/aQFH0dxVpzT8vHp7vC1z6fbKAUbrV96PMyxaCFMR
OmkUhWzyEw1ZjBRN5DBGo8sT7bzIBZ0ZZrKe4FyR7kzXZOuBWvdROVx3637Z
HmHAHGjHFurBAxF7oqUC/AqCfYLQNJvZ61eJAhtA79OQEhbnFNXmzZypHj83
fsagooGxs+9iF4Cr0UX+ux7MZienJGXjUiifTcmXZqnVUm1MkhACp3bkRohh
Cl+QIw3QjaYq9JQ57yFt6tQ95LkPyA8jPmbgP5KapqH8hNa8WZjzM8QKnV2A
zvAoT0GC0YwfvI62iPaoNENV5YAkZlGTd1SgdvM/SZBpCtHMH1c6ccdwB/8x
92CGRLsxkyN2ydfAwK4BjaLFq5cPhCsQszUI/7rG495iX3y+efjF49jxvhlr
mClvQ04s0HEh3VZYmYswzN1qcvBh+aDrJtaZ8KSEaDpv2/JjpkwzgDjQD6dy
LuCOHOygObUKN/rWBAaDR7VeKwaUzUzzt3zIHwDwGXIxSgzKLWpL+Ivlp2Pk
0h/vX9GJPsCZ+WftksExFsMc/h32NoCidm8GdMCw+bN6NTMoH6/FRObhhkaG
QqDrXXzbYYp61JqYgnGXZtSiGGibvVwNAZlZ7wgcKhC22R7stZmBsW+6ser/
rzd7iqM//gpEZi/YczXKFyKwBy6r5CIxt6kGhyX6a9FYMOxBj6K6UopWHH0F
amn6JSvlQYEEHGqvdu6lXR+h9boRjn+jtxj2wyBNx0rUmA6dInLqwM6LAjKj
cYXJwnRVjOeCIy/iiwwwmtJC/PDZ47RGWitf9JDj4lUiQsPZep7TiGfry7LK
oKOnsPPXOHF/cVaBowubP0mjIALaBPO9H2IWcQKVh3ZdJnpIZDP3awKGzZb9
BnngdJ1VI05AsqhgPsbR43y1kKNNJg1/jANQF3tBpVRyVr1GVcjLi0d1kLNk
z9qMD6FVxasyrmDqc2JzybTD1X+b6LLmfR/bSvC/tE3HjtWYuSeaS/fFT94M
GBo6YBZyJ2y6EJxSXgCwtdA8hPHijU1tOmni88y4dUpLw7oyCvIE3ocMcuKg
P3iy0Q5bNAQslM8TAiqvSjDINoLGR3Isdh7+xq2dDnf0tJ5USZkcO1RW1U0x
J8PxyRguLjKHuTYwN5f1rt9J2dC342b6B09L9TUDdoPEWgQGeLKHYWXVim34
7HTJ+KhxpF6rAYUJrgxwN5/CdxLOzjSb2/FuibphTngZ4/fgAqSZlrzCMImU
duKie4u8OV/8gWHdp8mKnoC8HoLD3Q5W3P/Oale6gCWHmEO9A3eBKngpE9H9
wxlJ63izaVFy/UTprfJQ7eToIGnQaKpiVp1I8HTxwx8xQCYwe+wpDxO5UHo4
nspBU5QqU0EgXpWEE24+pr8t2OONjFPbvk69si4iChhNtDlEBWX8FCyyUOkL
1lpM0jeJ5+Fr1L1OsJknxyWIOlGg2MKRxhkCNzZLOFDMBxApRDXfHtk5Ynlw
4asgOBubs0R+UziqIyE0XkUx1LNcyEdFmqtoFAuQ/d/WnYnPxYWY0IBrckwJ
9KsSQCKByJCMTlBGPRP7nfiHhlrYhoBt9544+hLv3rhhJ1nuVuuY6UG0TVw7
5pyVfw9xKEiNTwPiWYvBCGh+j3XPkakAC3L0l7my5dFwsuj9mjRektWLdAyi
BOuo7WYm4LKEx/xB/rlt+C0E3IA7TxsfIA3dsKjyVZhZR85QY2tiG5g1zU+z
XFSWVWVGYa+TNUr6wqvXDOZ2tv29AXupVhbrL6YF8XbtZl2gJUf7Lz+rNNbJ
DqmgGGSbolU/BgvLpJpadqVoRzOTarTwkqY44wh2VM1PxlB4EOZAw5PaM1Nu
5M70Y1za3b+ZI0pYlaE7gLjCN5pbdC0dSEBJ3KPM4gLoXByL5FXpwzlPh83l
c3ZGN5UY2wCa3qwUWNFy7qpSaGKNPoLWoKg6dMv1oJrc3SN2clRoxEsM1tSx
kFHRTMVngPQiFyG9zGYyp4+98UJavc+y0PeT8MGGfHAfjniv+BSWQMO6/8Kl
0bEAthxBRa8vc7w7TQj4IxuGoJNkj9uWYj/mTw2U5Dlm+s11lieMv1BsCIR2
X1oQlnUT6zlTiUoZ+BSHDxc2BE6g9dSlmQ11trooh3NyWOvlVkm9GEwjB6Mh
TDtMfPuYtUb2QR0YhC15LOlU4kK1dmS4Sd/34P0Mlr+v6XCLyyUmtKNsa9vR
2wjyCQqZch+kpZ81ZPDAT7rPamknJkPvrU8wYn00OPfCefZJ722io4tU0ArP
dnVGJN8kFq1KKfepZpLf+/ko/azV1vs8vNAsj3vMkC1a+dusA++Q6tNFsyc9
OEKugQm0yIzXtiFEVLQHQec8dUKWPQtXxbLrlvlA7nqh37wR0GeRLQjs7YEj
wEEYIdiwGcl1PuvpTlSp2WREAH6CoSJW6TNA++sjTLVcQu/F1CHfHTsNgQS3
ksOussTYzgMuNSmvkazD+sBGLjJkN6uX+RldGqtDh/6Af7mxMW00ufOr5B74
YyKriF1DEvQdyQH6lpybvo0X+yLDj/mwooe04L1QZpErej3Mfd+9vFSXdowP
LCDf9n4gJujq38jF9T/vIeTr2nzwXa6w2gYcO88+HDbu7xqtW5sqAQa4bJ2A
qOI/7KH8Ri0k+DUkG074ee5wiGx60FFVUrs3SzXi76NOUGOPisP0EaMLQGr/
Ug0Cvct9AGUMHJ0i+NVvfEMmMRHF4SYQ1W4H2pYZlEd9YEAuQnV9dx3UDnyL
DR0S+9ZJoeo1CNM0UA73iyQMt9lkRAeAdv3tt4FpqW3urmDMn1C3N2Sh7Nus
zjPXVZGcd+LqKC8berT/IDYATKvUsirvDri7cpo+pv5QYbYbrNtXyGAY7I6G
83dLUzxDQTGAdamICuQ59ddTS3u+eO6ze35+1hLMwdQHgaRx6HybUTmfiPwS
ugheVIufwm0NmEi1CeYYm7pyHDFSygDYPTulJJ9nSBQ7vXGjV3FtxEZllOnL
Xf8tEjlfyJayo1Feh/A8khmFE7e1IB30ILLpjG4Wb3hJpPnekUBM2LL77IeC
1EiFzHvYTYd0r+OWWnCBv1WaRWLW66XwNy8BeNpFKGGb6TG1i4L8gGXKPxoL
lkqtQya9hCBCG55wYqb7xi/Byd/Xe+JSoDXCQacaEAWdbW1tN0msPl+acr/4
GPpP+aR7wAwYHt5aI93xmvWRLp12Yan4NKy+EceRxpFfEGJh5BCc9z2AttTZ
CoS2Tp1HEEkIug5XcYdAxmUaFbierQNErucP5IVje8x3MSw9YFFE3CQaxHZH
Y4pziXh6eRvn1tsw2JRi9GE34lxlB+5utAbtfx0H0SrdaX9qjKsTmxwLchbG
jz8Ir05bP2ne1Oj48B66goo0OV8hFf7TTI0R0GL1kO6L+tpC02C3Hm3bC8I1
oOn9sU5YSDVfoB5ByCqVlW/PUdw3CKpDTSc1KfnXzZdVz5721YriJTzqBFJW
sza69jis9syrl3+oICVb6oSDr8UK9TksuZ2jpKjKeNATMWfq1PjFmuut9hhk
j81BAXty9RPFgWx/gei91eFKCAICDg7S+x1W45yVDGatONyg8/4mY25UUlPy
7XrxjARdJwoO7ZsRCtHkYIE++ROPLFATT2dZxqisBYOlxSXAoEhoGMRLtyF+
0Y3TRuGeZKDsfqU8Z4XkZVcrI7EkuKhhzJpeCCzrOw3cFV7Fi0kyRUquSfz3
Egb3BDJjHgAxQrBwRWBIUEjgV9L5g7W8ZCe0uVwmj5HgHihTUWE0Kh1gMwn2
abTWp1pM9GmxuiBjZe6vcKKqbxBP6/QCCyjipLJUxsJw7taBfF1FuCWpj+Kx
7sGR/1oqkErY3wArbfZ5OfvA98nT7hGWWL1wuLaffr35NHCclLZ6U7sKACrX
8d+yn/Ppfbvw+GWfC8szHqCv75hZ4zTiMJKxlGJLNPDvVtT3GTnAENZbqRhZ
KVsOKTSz4qAj5vwADBW/uzbMhj2gqKvsnqXy/X1Lsm/tDdA5iVMUcpGoWWAP
lrnl1S3kdg+ugEzDrGFxhCGAInROjtX7kSynp8AWeX9eM0qRz7ll6W975Mtc
wHjzkf553NwEuwzErJvvwuyk080+COW+0cZkw89wqrdNxXtAhuYwSbs+ZLAo
dTNcbQ6e7KshPskpTQ7Fn3RDD+VQ8HxFmWv6UrQ28LsYvyLHJ7gZpce80RTN
amflccJTy2fFzLs6Le+bIG25FpELq4SWPpd2bCv0+x4rQtH1VBzwFAbvjlqq
WM0FVgAI/bu+KMUsjso09Z3EpHmnqYYQksqC4bIR2myS2M/mzJB2Wm5qW8wQ
chtUxJScwTb4uQTbl0byh2pe8odGvaVnXD/OiapCyOzMErnsp8CDPiqSlMY0
MLYFIgmKkyWFhAR+ri3Jut3EgKwCrIUr5T1IeC0H7YfXUM+GEgkzWWz2HL52
2neQ/INPw4eWmsdwqDZH+3CbO2bWN//OqFfojvWg80GV+lBYwlujywHKhOwe
rLBRw23BxuTcpm6dB5kBsMfOPZfcW/Re1YnxnhCIUPb8t5jelbX+FVwJ2mL8
8H4EUT9+jDQutWZheS2HpuKOSsBxQlz8++kqgD6F9115uQ8eNr5FnDtckD6L
/28D0lVs2uvGDcs5YIQdqvPt4FQhE/0E9p5DO9KoAkb1veHUhAVPH+XJXoV5
SmLGJ4bKxzGuUbmm3sbr4VQNNIoVA9wfxRNZwy3sWxXj+XvVTBKYVrqHjBEF
URIaqPedxhSB7SjIrGREwK8PifX8mP9DBAlT91h8aUuarnG2cEkRJ+iZjAab
QliLsrAIXbnRqLniilBpENP8hguNP+xZcq/kAO3g5IBaLvvXakR2mFAvUmp+
FcG5MP/bR4XZIhlIdPOvluhqIonyscGq6gBF99yitFN/0myaU5IMrO9pU+d6
kFuMfck5Dvd3NpXOVq/Ii65UYyxDz9fiMbq6smK3VmJHX7pHgNve6WBQg5Mc
tv2ziJfbBRWgIhA0A+Z5AfLtTQm7nrduMb0a7P8XGF/plFJjchjELwAZIepM
oyZ9IK7ULPVS+hyvFGSmrXyjVdabKl0AgBVPZTJFrjR79vOBBwxSJTMCap4Y
oFPtwC8qoom+4bqvLUlxHhpCC4I9U6bATLyz4agy28GJlGOxCP0sxGmEvcDx
J6318QBAyMku+NYBIln9tesQMRecJqfj1t6XjNo9raH1tux5DCple0tGL7aX
0zIPojpP7L7p7Lyco0/KPHuYsAL81PIvkXrWVs43Gj63ijSX1pJnYaRl+qG4
TcnV7znxr5G6TXaaS8lkRoLKZ7ZtjUw3qMkZxbfoQ92Ncd+3f3bmz9vTkVpE
j53F2hMhk7M9a9pgN/SZY4EG6VdDVnZYu/6PFmZ6KQbbk1LgujqKfNlvcP56
2KWoZ6yGxAkoqj8lfcrslPUD2sMiCsfzLlCZClHWm7TJsOXJBacXbHPl3jZa
w/VrKxeNxD/D+JisHcnNVy/Wgj0h7eyBuDd4KWTMjeyGrbRoAgTksXMxaJoB
bCketaYAAB8xC2rD3HYMB30ZQHBDgcn4twTV/NxakNZ0wAu4BnzseKKlTrMO
UK/DD2WL63MssLqjH5fURLpBZ8+qRbgVmdkbLRdCsjzhvSKEmRMuNSESg5R/
WhwQ27Xgicsa926ZWGMXPUF+JEH8wFA3H+KVy9shvzF6wJljwNoc8cif4Fiz
Aw4KjiB6QfsNbq5u9KvV2nH4sIl5Ex50jiXj9u1+6ExIJSPV7OybltO7uVGp
z9Niit03OvLSRDPuEj+cCpvCVkYoWyO2x5PI6cu0V9rHUantBsP9MmS8v8ee
zp3Awvqq8rnwfjFi2iZbBWwjdCnbbVkaCtsZsVDL+pGoa8II7C3x9+9cjd7J
AYVga97zPTWxHKsvTIhaWs0mrpZxp7hmVkt4pBzsCFdeTWtWYT/Pir5O6kUR
ebZ0metsHNF7oIGH1WnFf42BRUe+ELaGRqsq6HtwUN7HVdFizhJy53vbS2mC
eM+McqvGydUja66fXwjuuHTvVsZ/jT5PW/y72X/k/pPcJW1vDf4JiQYvQNhZ
3s3+PFobfcErFeiWThwagMxil+O0s3uEnxXiEyk0c09VVoBo2V+VJs2V4M5i
2XnMiq+5vegvZNQ9i1LLxgQeO4wRnRtsLsd/7DnkPBeLUuZKZwcTFM4IjrYr
Zln16+4pqzwpgqIfEPHrs6WsgWSQSaJ+tQRsVA/qjs3QVAgo80fPkefSswAD
XAp0vQSvEpgqMn6DVWAleN3sArn/5tDgC0WqdKIj+pIVmt5V0HDMHD38C6rH
r0rT46o7CN4OW5zwf2R2+nb9HX/olallBAhBISxEncvP1UjeNjdV42mj7e1Y
mCfbShOYKSJ87Xx+qPeQZe2l5bmHxP3j/LpWycsQdzZ0cXny4d0cNfuu5ztP
hWicFm0Yt7QP8YoW8Odqpr2h9fY6CASMsRgcKKuFP75fBm+MU88BRfBa4eUN
EkecIX17mm1LXVkDrUqeryOWE6qn1TxTq5hpw8hAdyDaVTjW8y+zBrPO+KKD
+Si2tZA+GQWpP+RTiq4T4f/4z5anFOU4Mvp4Th480ovPzhC96WG8ipw7JjZ4
bNYBE6/sju5FgIeSRbnYlFrUvjt+LO9jTq8jwMvZ1oPdl3FanvyY/Iqe2YrY
adYckZHIhGt4+k2LUlHYXta18LHr/rLjZu6W6KCqvqavUD2qnj2lSwm5QhRL
DsgsOG+lLQ/8Z2TTnM3jvmqszILdOGxrQZMo4wA0+87efMlvT0sDkVXcRH9F
n68J59T9v4UrMK+kTAwRxduV2oSNzw+uMya/pzxcioxl0/knJKuVmBGkHU8C
A4l8aVYbORbhoDf7RzKDrW3AOpcnViZVHV3DY9enD0pEanKcEGywC3SOh04D
6hfDAu7sQkhH0bEq4jenr5Q88zRXAf30Y8pblBpoxJ8RSPufdUEj5/yB6uNx
eEaeImPQtC2qpP06grLAPccgQXa1geSc8VDssxAYXvVoLVs0lTxBEfikZX5v
qCL8zGCnQ4pGkwbkIueC3Am1O2nxqiI7wr83NQ+hGUa6E4CJWsQUYjMYpaWG
hRyzUnMzk2X0vIxRZ5y0QiBgQa42s1UZLK+t35kS6ViFfX2rM8OzkySVnX/Q
noBHeEpU8WJwkC+W6dqx2/LiGAG9m1sTc4pSE3UcZm1HtZu6CoS1UlQI9VU3
nZcMJqnr5AzsOp6tod1MwZspbZapQcA4RS+Re1gM5Kj5VUNOlNE/y5uBWo7p
xDGW+5N7WGezsDRjaGY0IRROocPHN/xlM/AEgLreLM60YPTttEwyzKfUjSYg
7xEl/zeQuzllcT4j2GoJQ0fhlKoCAhvolHu+3yMf4M7d0iK6Baq3zXcc9yFx
ABFTz2V2ApFxWLLgsnSJD0DJ+UVuxxunESGbf5eD3CWvkypSptNpjdbGSKK8
gXKvpi/ImUmiFvVGpCQNhLR3C+B3yZhKjarvMSGOzUOmT2P0EchPNT4u0oj/
uFNOy/szhvHo8mK0CwPCG59OZnLpJYaYdnRlBo5RjuAWFxIqB2Z4bOf0VanN
/Y7iFyHqDzEGvpZgalZBZqT2cdzH8YUHoBC0c6P0971Tk6NPRjXq3ND0lU0v
sUTRvngHCwg5HntouEV3fFdPd2QmYo2BalXzX2PDRvp4HD3KfuGYgyirY3UN
jZLhxy0gSoXBzzxGR+3kMGeqT/kb04Ymr+chIGJwqkzeVo3IqeIMD6rCIXIl
g5k/LxWiWdQhZoLLHEkL8W+i8oVBG/EGmGbfsGpvKcSj+aRk68umlnnen/DG
spbXw+BmTlf0ao1kkK0Otzl4Y3bksqb7p8i9CfSfTM2kN6mE5lij05inFiHB
QIWeh8CIcPy2sf4HOzxXsJAsTHNOjRLPmsHe4KbY/ac5CebUxOIm4bbxXOED
vGSc0I6DONK4y2oC65VPkyHJfEUzP7hpifqVlgqEZmVndWjlf+Jr9NeGSJAD
WdlHkzI1B7k5F3eZ+OuCK9kWwotdRdyav1zq7vjpLp+DvDYzfvcOeuBk8XKg
GXb8vVuQNVeZqyPx87kJt7zM1YPS+tC4qV3C903UDmDqppKu7zxq3GuzXdCs
UYowlQOn538bXGl/Z0eHz39cCZ8+vzkwVmwVGNATO3/JwloJ+LcxaF0HAccZ
c89cVtqrNjqdOMtnANYgvfl9fh5zXSg2jVu+h0AE9uRUdnbZy+6Pvqk4ha9e
GRBx5PuCY9AA8ooj3rJ3eItVWOS703leS9tFZFuEcb0fyoGtR1COuffzxZ7f
BSQAZSw/Cu1Wu0PP6wRpu+gmZrV9uO9CDkk2aC910WgO5OH+jPWI0bECDkGg
2RL4ElryekUIq97EYZ4HGta4pWdKdB2VJfccBAg+2SC04Tv+NEYcngpEoQ7I
WG17i6l2V191avjZM4jR40P7jhIFY1nC7cEXct23ptXNMLFw+64NdRdl8sVu
mkF88Yw3qcv0k7AnTN39oAL0CtFApHTGIAdqPoXY9lNyIwhi7X9kofB7Z661
pqgkdQo0kWJeSiglFjs3XQYSMzXB7upl0bwrouU7ZqQFTSYu/48uyRJevndM
UiHn/masIWNM1FZxbEBLoXNJUM6eFak1ZhG19xu3AlPxRfy5hcuNWjc1idG2
pWCkn7RvV0DyTEaGpy573K1Nr4B27vUihpAEYnYYacp1VZzNdM7WCRg0DIPd
H442fwVoeu02AXYD11vo86Advz/OQoSb+dKNd/P4Vyp04XD1FW4YI1SzusTf
ZRMSEwzsuJAyMJz7DPwvg52Ud4mJ9p8lt4eZCjapfDzwd/+rZNY0rc+jjxkV
FmztDnoqbkcgzpSvQ9Ad3dTidPwfbw8hbT/+fCh5Xpm+tYkLIcsyfoYSllPK
42aexoULpd+Mg9NlVOqWbKsBnr60D8kMlbQ4nALbo8xNWjcaODpnwG1PsW9T
4ftuB+TZma4HKgN00x6Z7haqpTe6UerN64mYuSONRhu2m83t+nO07UnnqloY
MxFTpRpM0iEpU2/NHIB2JfNCyDLRSzpXOgtCzksXtyXM9dnBU3/ICJQ+lXTv
/YwyBGOD8x46Xcy9FIBo1PDyP1COwhFPESkq5Uybs95xXLE74MbVW8YOBeDX
HgYwlTij2qK6XmfGMhn0ajnj+/22qK95qEbwl3F8NfFA7NwEeOfigp+6QmCA
fU2LOV0nuZZB/V3Ttx8glGsIb4FbFkrVeE+qma3IlISUpFL8XTa+VNDkvbXn
zbnAZSs7KXiw9nugBreW9QHOZNrrnI2DTScQXDH3aDfLdLpb8MnKwxOKcgaz
Y4tjyAph/3+HXR4J0Eb4ZZWbHKOUWKOqyA37IjIb2g+NimeuN6qtlVdBWJ8l
EL20ZPqB5HLX5J2cZhU6mcYtr+Uo7jA6L839pqPDGyITKgFXjzrqswVQ6E9O
PxxWDZQFdZZED9xP/W37Kz7LK1pokyf8I79z8pxenVT7l22JQyU4S4bA27Mb
W3amY8UcNWl1V64Ur90u/rzil5vd5Ir7Q2f6w4Z/YRX1JLBOcg3o43++3z4f
rPW+BIkHlzzkZ040QY2um0Y9fsQD90/CksvAlr7CRnfFns0sru0h5PSOG92f
VwqDZUUCKCN7psgA1WWvXK8r1w+3szy+VIgdfMURBLM79whbEQZiFOgnS/mh
rL7fKJEoTBsN6tMnqCydQTAC9PCXYWz7x+HmBiWRPJ7R5OjknQ3CriWIe3s0
z6ccWcNXygCcxtLfy/cwrsLeU6gF0Y/tAoocErq5V7FNXIc1Ofy7NYILwQJS
vGzfJmhuYg8CdGmrVXzIKYJplORdV1uC85Bdz2ByDQ8ZbwnhQKFqdPbY2rwN
BtjOX4X7+mMHKBTHL4d35m8QZ4PXcLcaWoXTLLyT9ufzDFQTVubjsKrmXILm
xTHI3KpRXagu6kSiqIKTii3ItSXWHmaMvrfScZxQTBMY6R1VKx3aedkdp881
7KkxOHB6R7bAUf6r+kgjt3jLLkQCbUmRBPVazy3nqtCU1iz+ErRblE2leNu8
kD/sp5Nied/HAfUCOELHi+7gB15dC6YjkVdn+5FcdH0PAJ537AtZZnWXnjss
S7Ph7PcmpXcQcqGuG0IwCsn5VD0DV8rajibWwMuK2wZQoPIWpyUpLVi+CiAu
ccqBzY5yhYL3zGxyIQr0cv6XhNJhsQ+B+zFXudPD2x7u8v97uJB53nc6RcUb
ogjEpVh7v+eXxjafE57BbvhfmLRlHnBsNafy+6kx0O622zzVn5wfA2gI6tSC
zj69cbY9vJDLW51Ubmj5UaNmZTMIzMMThyFcbAfMmy4aFwRSYN0dWSHl+eoR
r1OpjHm/eKX+5Wm8GNW1oYrBAYiII6QEI2QAQQz33igaarzbUw9nZb0WyR1S
D9N/pTiBNBTVFZ2DMO4PNQMEn1iV2gbvY0MHtwGqjoyL7fjXNblSrxRKMwbS
llflvvs8boNVTyqhO0Rjts80ueAaYJEXU9o2E36NFlz9xFWWfNNgvYTnPnEf
Ba7JtAWvCSGOCBm0JZfrGMtSYLXDNWEv1jXEGaSttrxnMTHW4VBCfTddKa4S
h/s/AFz7dUoYF6kUwXZaYlwmqyAWtfBYWZJAdU0jt6+O3HoJZXZj4f1ZUB+2
vbt3rf76ScCeG8IAvcmwjNRzuUqjYRBYWEsvLlkUo9jpTlXWnO8u9XBcu1uj
CDH6aSEGNeGpUsE7jJeOwC06xg2oaFnL/F6doEW4uPZMFWVGMeb6bykiREGo
5abx+kIqnLdTzHLvET+Oo+rFDo3RDYjA3Yz/pDXKeUK9AQmNUI58DDcPTZde
j9Pl95qOQB4vzJFR3usqidpj6CSfmrl+SUyzMD0NR4Q4XUtOe0/Ycedrnbw9
9Sm3gnnaBKILIbIuXAEtZ/Li0rfb/uK4j5tjLzUvnkeMSyh94V4UarBu6lgp
gTYccmRMPYD7eW5KiWMdTXLF9DkUs33/ZPaZatoHKA0oDXyXWiZmlb/X84cM
pCgfvUaqPDAct/TDFMAbGkUrr3Q5adHMXI+VKPa6DrbPe4nCrOHWlMwW69cs
ubES5RDeWbSuYHSVKrBgxoenPQv53wOgvTmGeoSWWHVDvQ0FVVKBW0NrlDUq
DyU8UhrfYuP4+Pei2iDgyIJTFTvpcTsCeVUsDiu6K6shkZq5WHJ88Gs62iVl
akK9fn5Tsfurn4kLEOPX5Sk3pOmFFJMJbRCL1Ut1HxEL+TnyDQaFO7tqyrDq
t+i/DtVq7Y4gxGQIyB9DCzpC8YavIFpFw/8veu12xzdiFMlr1pnXqNqCUiWx
MpalXgMuHLDMRJPekuhP+rKRKJxrxFxzvqAhFQYvYjd64SRHdf5Hrli3RhDk
JPf7I0s+00W2sqpO7cj4ED8HoC+zQT8ohxHd5GX0Sgkoh+D2QERXfdPno3Ac
wNg65u5F1T90tY5U+6hFlpwKbbYaRvt9NY0eCxBmR4I3OCDNv3GzdNU8sCuI
a+W5ACZEDSGJOkkC9QP1B82KeP78E0gLf90K+mOrq025UuUhWMClB04tIadt
GVUH5NydJRWTkz9o0RAcx0M/ROxiwkuG6SPIT7PUl4w0ADfSoBwyDTdxi3TS
V+AYeA2lHqMvxV894snfcce3XfVa4oAVoHqstxKKS3WUAY1pK95u8GN/wMG4
35olSm2kjYEmTVXXSW4vDN+FpTYsKaVgMifE60WcJwOg7u7ulMEHhuRFo2A8
iqZRWU+3A9shyfgGhFfzkEVMPG0fhD5tR3swGT7/20E/zoyijLxYs54z8/N5
56Cr1GgA8QX+r1ay+tvQU+ivtmEzVLDom8Ptjm3eTqOLAcEWxQj0Pyerayh0
JvPrfJZ4chLtZ8M7VfMp+y+h+hzaaBLsq6Xjim2fSRn/rNbI9d26XIqO2+k4
FImlrHXFBLifLMWUDJ9Q8UZ2yynPw4pTUsTOvyz7XdFF1hXpvEDv+/k/W9NZ
9jdaCQxLeLdWROwocyyIY0tYucOtC73E9gEcH4H0UtvOnxnntgdu12Epa/TH
H5fUhMzTq2F1oJVDnZ+16HZD0JIM5ju8ua9IRrgqfVkMuObmh8wMF7Lhjd0b
hknOx2wvjrFnzH1maj5tNDptaBAAiTd587RmYU5ds2jtlzRk+7xuLWrJCzA6
JN6kxqEyieqn61olTRbHQQXaaLhUGHNWGYtcAnfHfsq8cB0V7d5Nf7kMKLrX
oncG9vAQEMq+EdZfp4op/UXBYYitdbqNLFh7UuhsmDd25j3uuXUe0G1IEhRw
7wEDL67JvhAgDjqRG+6uDnLDwf7JpDy2QfsEeVNbMjBARMbHoFuBoEnly7+Z
lRXOWI2BDMfj1P2M/MqX/7fCdpF4swftrYluO+c6m4Y1jVnwYF5J32UjT46o
NN8Hqz8vCzUNCNL0w2hcBZfl6G3OPaLveUaNnka8bH1bUSoFcZ9KbSe4IHip
tO/3DoVnhvzNl+fjE5wu1M7fGBGJZOLnBudofgsL2WegfUZBj+SW7+rfeCWw
3XS9I0QCstFlGV153vmCVhK6PHs5O+8fsJHUPIwP/11s0i+ytcZf3H9syQeQ
ixDt29uxbzqzybSKdcZejZWk4hzME3qtyXCy7JLK5guhxaGzw2TG7c6sv6cC
WfEXlIj8OviZJF2WJ6x2wPEkNgy4TOCDEdUvlbwgU3IlRjDEM+6ZPrdrmCHY
Z/waW5pqMVX1BehmXResbJZarqskcMNmJvYzdS7W2XZ/1PbPdzFuPV6aX8QE
QcKuLra963p9hVjSwJ/Cn9/DXDxpEVUpo0BlwbRz1arGO4Exr+8e8FQr4gWZ
EezqmURgowfWJQRGF3cIwT+BQk1ZfBbE/gdfXbppCvrmkCQbz7tq4DEURdYR
UcrWxxW6/OCGYqawuNyuYRtUOH1XKFP6EFQ9KXb0uuaD3minTNEDVjer6igk
+qehj9S9y79HrAPn8jYyiBOoFMlAEZSlPcov62fhPftlsMAsC9hqGRsVpUJh
IBZ3c5yCFSVDS1+7cPrN5sTH43QVkSVZkGJje1fjtfDmOEFrhocnWAhd8VHI
n49jnZ/MPi1vN3CVxrxPi6QYOkgrXqXa+DUYKWCg7NoyFUcUE/Ef40VOo04l
3t1tAXRCN86SY4XNkiNogNWlNSLOjEmsePJgTUVBstlXqFVRL0vUGhazYq0M
6FLCWlLWEwocbmb1R4o8OWjRyHkdfnT8kafMVPNuN2gbGi9zfVtq713dw512
fHtO1VL/r76CXoMoJ9hTW3DRmPyZt6SjuyDD9DBOA/bHfuExW8mks3hwoZRw
exOmxj+mSjxnionjHM7PrqrqTgfOT69AR2dmJDMm2IEgouuwfH8JtZHwDTli
r3D3tfvZWk+FaVaCMDzT/AXW4FvFoK7qyzmgHReKh4J6XPC2fbDZSue4NQZ9
VpZ4JiaBavLfehGv/U2OJ01ctLexylSUzRkTuPbCX9Se8cHVfxU8p2EQWc3N
cJXLe0NUOPyoxumulv7E4oF/EKtDWhhQw2rcZjUpy7WPsRWYtBfzONf0ZPRO
4uTi4G9zupL8UiOfmHsbWng9DVVrA4uUOo6KW6qob3PNBiHy9IsuL2411RpO
mlwNlVwR8pr1lQNKo7+jUpp4VfIJ9P8OPv5Nfg7IDIQUPwLbCmT4+6pGp+Ah
q17/Abp4KfeR0bGkn4FBw4cd3Auq0O2KWquufql3NBdCQekf0tdcCcxaIg6M
WEuxPwPJSe/6R3/0W4VCkHsIilSxRnTduFnHrWWXUDJ7E4BssLURVEl7nmcZ
gfzlYq8R/kaU3gXX41u1Pbxm6NZOe81/FKz32IsJgGhCJAlr7WsXBP6aFsGW
7w1tuIk2b3XXOzoBYMDZKwjT/n2jk2NZ3deAZebEp1tWDrSEnlj9EZroSPAU
z46MicdIpa7BhpXi6FKNovO7To2stiw87jJ0skwxKgeRil5LX2MRePCla8wG
Sacxwy2o2zZJjG8Xn5BnGmU+sR/Hb8MWd1Rq4NfawC9S0kS/oENDHLfDSFbQ
yhv6Z8OU3FIIWH3iEi7G49mLIXPft6tS/7gPFkkDEvF/hDb9JtQZX5IvDPTY
RlO2XkTVCL9NfOoTzkFReKTdv9izoGO8/+R0YbgX8R7zcytcrXZG9463IFBM
UnI9JrwYf/+zgjTtX3izly0cgZUXVabKPDx495MvLVQH3W6J49RhAMJ1O5We
KQA8h4YK1WVQvQ2LKrQJJsi/FSShI6jMztcNgvpGsmJUQD+a3mia6y+s/mOe
3Be09o7KNVBgEdCJhby3eb09wiNXNJF+yUtHznquk1jMcxTyklzeNQLYr1fe
WPjmgIpNdzYQYj8O6qttt5+ITbz2624Cf3i3/G09YBrs4Ssi51djruTcA4/9
I7FklU504m2PSRu5NP8GDCr5N2Hb+vHUt798dCPJOzbcfqNqFO59TM1fb/jU
+SlMnQEDrWPCTIviUYG2F7xShuImtVE2RjPOwJDmK6XDDsKnUhJtNcoqanuE
JY5jcmHSEeE/x9LKbJ9IGPtH693kHxRALWDgsTb53nO3NLjWmHyswjTpL67n
N4DdVQgbt/rzBUObyptviOJQKKxuAQIbZZ3vCCmP/mmtu4FwY1tMPwygzmY6
i9nnxQ0zjIlCTnQL5LHRBRg82XGiNJ3+xQra54U33lhaJPYRLROTJaL6n7eo
GoJAbz19+Yc9TXP4mQfMt/lDhbSGyyke76BLEnOjG9Md08DS9DhREJQ1GXf9
cxGtqCZwouhjc9ge+GZ4DPHevPL8eNfmKQWtl/3AJKh7sVXyUCvpgFaEfCmQ
oLh97JfEDbuVpDHyo6WXUIBAz1a468qkfvqis492Fn8iME/Ukl84+Z4rs5rn
EKxFpZRn3M7WodwNs9FkbFeFI+2AjLWp+hB/iaU6FXgva+oGUlwwNHhAkB57
+fVp96NfUN1x0y6fKj0tLsa3HjGivts8riQguaMyXbQXUMb6Ucd2kdyZ2A8G
0S+lqonFlhkT+0rNpkisVKfmplH3xGBgHEY3+ND+lsfFAtHGNJ1Uyfw+ZU/D
h25y8xZVXmdAcD5/En6t2kt1prWyuihJkV/860Xt7GB43OaVbf/oaYxGf8Xw
IxGcdKGKiJiC0IObx3+hj0AuIaXdETEVd5QzWgTNPuWSAFdU/Wkd/4OvX/E8
FLv7cJp2vKmtPXfnYDyUpX4BNjQS0tyTplTQsyCgyDPKJ8xiZBah/5efgUp0
tSS+t2p7BImwb5zHoFfTyBGKkaJwiYWQDvZ85wAfPOM6IRuzZWzV/nJsTdkh
DId6MpMKWIe5COI4US9D1J0mm+leJCGJ8F05LyVdayARB1ApWLMHBHexIIjS
acr/vtPEGxdSNrbYxDtv0eNEvYzj0LrpyqAErrCaYcTrxDnk5BbcxC136kgA
rEu8WLJL9BsOrEuoaqTM1O8TY9ZnIu841Xmwo6DFpBv+kO+mp6aAUVwMsE+z
MsSD4XfGV+ieZ2f46xHCBHnClN9Ftjwbos3lb+TdyEMUD8fMmhqW98WKBxdL
lVX+gm8WdEu7l4sXaGdGXDbfxvpeu0kq2XGQAwUJ8+cMCoaiEoLiakSQqcLr
/dUDucdJuiuIt+TcISWwGsOy3reITMsMKE1XuD/HD0Lg8Azr76FSAmhFs/jf
sCpiYpY8o87wbVkK/XUQ4DG65C6UGonxpuJTvnXOdIdrT6rnfTjONIgiTAJ9
wCX40MetOyt/Ls23WMwCZQQWvNPhVsF8DhIl6ciSIvjAQ8ZBugtjofbEEm/W
pVwwFdKjpEd87YKF4I1L3kqwlx5oUf3dm2SWnUSqb6+NsRP7EeF+iP7Vokxr
qGQQXygrIMfI6GSE8S/F+j7HkLewzNbUgF7sW8aew02oMcDkaCBlmFxNtpV9
Cr1IsQtogwTYoG5uu82pED550zIhtrcEJN1AIjJVGVRTF7z0127y6heS+YCJ
Y9JhelE9FpytXSQsfOHkBn88rfHRngEXZJ8d9L2b1kTCa8E0/Muylj3r4dg8
gCakFLivEQJLd/o23f4RmgtCSa+U2Ma/dxA+bAfF5x+U/gsaIXlwrIdOzFE6
97JLJ9H3xCk6JHeDfeS36ZvWZ4l63oGdEcsHtQQMlxCSgqhElvq2vvt4vbiV
+pSR5uwTwuzooDXHwmIZWJhkSj+onvQcBetfev7X8+YaTRhx+jGSs4z8OkZi
YuHkI5uLupA6tEwInHtNOWmwaw2gTVNr1sd0hnXAhreBn8TB5nIt2bG07RBB
ZY+gDR9FyWDDubzx2d72jNDTdCiAgpD3pZMNPLxFxV7XQAdACHyUH6mCvZVa
+tUmCqDlyYTD4pja+1FIUyjIQQYDNU6ZPp0FrGt4NA3GcqAtHMhFe1eShlm1
VNYtbqacKukGck7pxhA2u6wuK9mLOEYo6Jtgo64TW9IEas+fnNG5fV4tzktE
xJ4ciKEQ794TH+eZPpMHnoIx13J7yPTARLu2axEyFDO3lZetm+MHyp5nwQlR
D7sXLhZsZg8essXZdTx//1TMdlj0L0McdfZHiqtAWwFA5DRmu09xWpGOMG5Z
c5ungW2NXH5F8/xvk1BZ4SlWpScKfF26MH/U/6JiNvhpQltbh8S5hHeSbkhX
C16ifMzJtcc4crqliAng6996Ijwb/s+74EBEY9lgVGU+cn++RXbq5pV2EX8R
kz+pSDdILudIVqSt4TUDjLJfihIttaxzJazWImg+Qg0usd9bTvwxOPBrHdYU
4gDuuyasmkX/gLiaOaugYMIuuhqca/0lWcClqTF5JfzFulQF4vGIsyubO8nh
FgGZFWuGva7SmYB2XW4amyNmkGiI4PGn0vdGJl0swo71oNRHj20zjC2oJ7E8
S+ta90lvBnYJ6/8Ies6AfOfGpLU33wwUHBHZ7MQ9DUMOq4Fpk2bUAvZfGl4C
nHIc1cS28GfAXrGeZ74c8qFPkEs13hzxfPT6QLIInUmdfoPNImqXtgApp9wN
zxEtDwILYEgLwGLLRcLmxiY8Vk+6kgzPs582IQWt/gMUr4L8MQ532DyJf02W
jZUL8PAudwLiaGBifVm2tSO5za6eW0NB9/w+1ByjNUMulpkqdk/GU37rY0Gl
YMaFPQeSpRiod/0nYj2xLx3d8FjrvD9Jwar8m8zm8KFXPQAeSBaHlALSMFjy
VKn9pfvKEWCXnU0AJBlmAyvvKqtnyavl/2cRoEYvNPSVPGLaXJ4MZaoQO4uS
RMYwFQ2VBLKb4+JXtkrV4tV3IyfjNB6fjj6VF5IxgVaM+SaxjZfeptHTEUTf
9AN3YarbBhrKc47dlwhhxH1e1HBexl+r7Hypod7TWkiPV6/rLto+nw9HEU8s
6ZKB369H/EwcTS7WXvfr+YikxmK7+sILFz1gPL6RC4YERA0AUdoT/Gh9LRJg
kpWPGpjEaH+kwv95boQHpDlaljU26ZBoCL5zj8Kj8amsgLaCN6GSNhC7zbHZ
g+iMn1iy2mQ3UIJDuPHhgA5jNGRAQBh/7zzcDe2a3d73gPOgcETXRzdFC0Qp
ubImbdM3rcwncyjMwIZ/VI6AaiW3591N+vIbqXoDJG/Is/CV+7XS5BUSWiMT
jNnb7SivGtfESGQ5IB9lpV1XnhVm3zWUdCfFtN888xiGavl3u+ZadLPJ4UB2
/awVYPeDU7/vxvsWCae7pg0hlOOgMcnn4IYXGCb9xGEO8CJqYX1kGVltlER6
05tC6WJphvHeTqOiwEkESEjsqkhtXihjkzR+PXpn+LZ/coNumfy3tzI1gvZF
vlMMcZ3FnmWkZ5ciox2i4OTZJNeYhpLRkkIW/yHmyue+Hcfn89pKiAdwrPEr
lui9lYwPhiRg8ffayz50JspmpHG+OUL9HnuKkgQMlWeMsHXT+LzPEsxweeJ+
ETNp8hZUeQwBsPpUP1/EZQiJ3ScmP1wemF/ZL8ZkeVVimoBS6sr38gA7vAig
yIeC+JTMIdpATVBq3eIPqv1/wMAxZc4hzo0q+tQhOocZuUOT3FhFT8n9CY2N
/vJHCc3gG9Y4Sahje1n2ZHuigzSXf/zQGsNO3cOxF4jGFnDF3xp4Fc1UBbCX
ZC5Pg0v5CkjzkEoGsdZNqYCbRsJK0SjdzwDomjP5LbYfuXq+Dy8GsG4ZMP/e
VLL+c/K2O10i9AbanuNash621HfvFHu8egsGJbQSVqP43hrS4kVeXzIzmvAU
JoiP14+eYMWF+UUquvX355lNcjYHlrvY5n1GRkqix8/iCmnDlPfx1e+8arQl
mAkmg6RV61fvrX9HBTOgJXaUDLog0SidoY9VJEYffG9pfkUtiKCBG6qcelv/
tD/T/KdryAF6MJjuDoTc6qJPSkGk016slRB2TIX/rIIySJGGessPDCkbbmvc
edj0rZbqJmNMImJcshXSZi8FDB9M42NZaAdhLVvcjBnlr46Sxal32VRYI+5o
wB23UuKZRMDLPcykzFfxBlHjtEign3lcP7nSnTptVgV3ETOkJygPxK3rPc+q
edY9omByStEDs4/0qGPAQfYfwVaTvctCvLykCeoClWCg5h+mJE3a8ylp2MjX
ZDgySMMuCHVMm1Y+40Avj2Mqvo39JHrP6HY2jozXPaEy3nId+fFOZ+uFtsS8
9ijLFcm16bWDfPULKbbwNgSmGd0QqjBc/yQ4rSPIeT77f276tHNW+uxzZ4Ce
D8lTKjg9CnwDeqq028ozSspaVzE2Pz+2KPlWpo2xtl3XeW8l3b15aYmq188w
2TuWpGsFfJ+JF9FvbnY84ko/IqxP3VxB2rxzPCfYexoeyaqRfPtZdcnxObeP
/pqmmdSxcX3f4HajzQuiBfEc3NCj7wPpFO/41DBYxFTD7cz2iDfEcXMrSguJ
eKmVLOXeWXigG8zNLe6uSnq7k/qtxQ6vSkKc4QDSwbztmOu2ZK+Oe3JPTu2M
jgpnJRAfDQqDQIJEKABfZYJXavhy0P2ixXmHsri/U/kt5TxrrFDnX0UgXlhz
/DYug92JZg+ITDyYx0Dsr2tuGIiGK2B21XOlFsNgXPOiOPS162c39Um4duuU
jJBs5/Y7fq54nBQO6EV58VV2W42tngIWdfxvZso8ChMsryb57dSBjVx80ITq
KHkdbyJ4fl4pkKg/60HOyGKq5SknHc1RS4FU1qETlzW0A1PmHv+VKMt4nxDL
fX/p9BuUvgxoJp1TZ4x2KO+XK6pxGq9i0I7nfLDItimjgSsLGn6TZLF6Sxjd
3kcK6RLaIMGqY8SasbQhfC0kwQXuDJVsj2NswRgA5kzyviGrMBkrXl4XsxCy
KQssv9hiLFi+d/0wDZjfbNMr8B11cvl/M4WS3sJNcrMLNh+S+YXEzOrxZypp
J1eo2FCAuPueRRKoy2Cot0TGqaLn2gPfr7jFeGQQ1EsUwPr9j3t3NAql2rFu
VgZ8d+FQ1GqPZ5jV0Z1nJ7SqYj2aSMiLOl5cvuex+K7g0t3b/OxEL51P7VTY
aD953k0nbGFgE1q0EtLguEv02nXf+16rgiNyCf+AyBR1eLeVvXPuj6R6x4OF
F36c/FcVd5XR/nYFKHIML9ucs3bgKFnw8LEkOMbzhBZ+UtLz6mPHgOowXqxR
aIN5itriIgqyt1LjmAhkXc5suueS9Ay5G3qEoYab0SV5NsOtUBBNTAkd9zVG
aUliE7f70vrxOFA6rxmkTcgDfJmRBRQeD/KEur32vpulMfKPgSaAZ6rTExd8
QpThfq19oxFGjXhuG+JdnGWSyaTlERAUor4qIx+YSStGvCrtlQKyaLWzaf8w
Vpjgpuri1jyq1ur9wtZWstq6936viEZ6aH7MeGcFN5ehAkJKAFLuuE6qObZf
H/7H6ch+n08JzfcwE5abIWj5zhpJsN+Ar96OJuknzMw2FyPf6IIaM6oZb/Rg
v3zqjaLnWCHTswUl2+fiRswao3FZ0HvzLkdovUoG9MjQ71qip/4TBwXnshX+
QdGlCB5OtiuUPHYq7UctddpROQS3LhvS9jbx6WL4e6jC1Hu13rJf0Ur9envt
JSDSr11uwNvRiedrkUZgo92HcvI186C71JVhp/s4eok67gmUWiCX5fdimeOF
rluH6RSRUrdcoPAL2fyRWvgHSFo1mdNEaCuZqhthk4QgD+mtNDO9W1PJWjqb
PpKA2VTT42KAEA0cBB4Wt3PHeYfoRLfNJhcmJUeO4z6AH1wBmsWl0AS1dwKu
1IhU31bI45jELTCbjreZ9I3VIPvtVHjkFerz9GO8YT0vfi/jnVQ6tXLYVc7M
jjJVg21eFAYVOtJjRftDSFIfEgkCtCw2vU/welEMUu65pPzhm1DrTJfQj73B
3jKGAdM5Rdr3JEgudpJIEvi0C525SN6NGwzrmhbJ9F3XOpI2cSCCTmomypgs
uKEMpbkTlPLp3W8rdw9N63818X8xT68BqKaPNNaTRV3r6qm9dtQ5s1qqvxD2
nprVwLCAFLyaY3fUUFunkqfBYbSCUM2mMSEyZYeDU/HsOIHhQBgG7/v0rsC5
3k4obf61XPrGcn6cceS9OvqgWI6bNzKTbjosiRXRuni8ugzkEemDSuqiL//L
BRjesLKjqnQz5Y21P3SGDfnoEkm65UHekJ1DE+8WLkQWcib4gJt77sjnQJma
GeAw5SnXZmnxrZzPNfZHZhdPqzM1NFxF+ebCoTnwL6dlmnzPg4Ve4zNtzVa+
JJb0YVmsmSGt8v7YeYVy+Jx2hsy3aks7t14HwUswwwpaVGcx3XdY2PnVqODp
9N1tLq08X2RVMORYitupibdYZ+hgVx1/SFCgpIcD4tTl0zXgfajw3kviVnGP
9km+iglQ3zi+7om3KlGuf2jOcl3OrejFCBStdQjlF9IPcP/GF16BDb+tMGzB
eMP5lKs1Z9li6iIrSk1ybYZI8/r5kEmPeNr62LL7xmWK8GY8RzNWKpMlNXZd
eJ7PVrE33meQifOhFUlyay3ShlGhjATYIygHwCmHU/nLnxkuK/IEQ8fDMjn2
Wnk501+5uI3Ql8XwPxZejWUgYeP10DPWeBA3GNKX/NqxJQa/gjN8HWAGKsJy
O4n5BNhVAXXXETmi+LjES4KN3S7mJw0rLWG8PAD+P/rG64juenukbUAGSfX9
f9O+WOmekGzFjUPOtw/LSoOOOx+UQO7uevzaIcjMhVuNrGzAXLjeM0To1mJ6
KRYiOm/zuX91cdquf9JRwzfMtl+giYyOakqCm47XGVIhndzxyqaKBG+ulgL1
B8yJAqLL6RTsY5FXuoQwwfD3JF156o5z6w6Qtmonbg20ixpszx1o/MeWCNG8
DLKX4ZDdf4OYjNpqJOubgwsppy48Q0MlW9ZXvcX+LUNz/VzGLWekoFsoPhiv
ylCr8JZzZwYFQIPNQIVraOSsBtGeSQF5kzUANrmKlOTdFz9LZD5Igi1B+UZ4
dxGS/+Eauiv+2LA2leAmtk99ng6Fgjnu8W68qpM91xoTqfb00HXMqno3bOjI
yBmRjkHYHxl+xdnrScsBQyjFY7ta4Rki5fRhF7hmMZCxevh21bBy0hNFI0YR
CYcX0W4Y6FF5ZFmFjFbyusX2CL08WBsZMPVOqXyIrTdL85Yuq0rbW5YlyLXH
E9UQRbhlZtL+YcJ/19RxKu/eE2vFip14duTk6B6fiTpcZ2UnRyy3UTkKh26S
lKudD+qFtqtpL6co+RHin50nRYB28ve4psfw328nARKuQvIDmeVNPYFmwXyv
8Ns/5P+j6IBME9gA3b6TERSczpwLvKxGY0kft7Snz5y7rli8Dlc9QaflmK42
o5ram29/OmFdzJbqqLFtCysOB+kUngZfs/V9K+7nIQNuxJYw1ToR2NJW32z6
hczJDqmjcefG2fo5lGaJseH1T30fWneqSoxZtI3TzpQwHdgenRWSPDFzBBga
mQU5DcxLxBE0uVMRccNI7JE83fPOBCMN1chyVs/vnlB6h5V4qVYh1gyttrAq
Pzgv93VaYezuur5QKPAkagainaOUpDN61wuNTW+1uZGwgEFI7L86Hdd92Jtz
6A9whrnnbEg0SHAz772zTyCcyKbJTC2/0cywHM5SLCevx3InmkIWTkHWrvKX
d8r7Eysh+0ziDtT2RxZmEypAkPMZ5zJJI/8/zy5cMqWE8I6eUROdnKYaGoC7
RZbHt8vGIW0ad5Ws1uB8ANaOltRh3osH9yIZ7x5m8XxTUbbnES6cn4wrDIle
h2azQ5fqidamxoLirwTbA5r7cVFrmYeFni37GVUPp4DUQj4BeDx58y7a6aOj
+A5GQjxYMyxs+nuPyuWIEVJRKi22xOfjhprkeA1khVSUebs6OfsLeIZ/AEzx
74IFIlE3sq7rXEv3mrQ7T64d1hXs6u4Ywcq9BhO9RJpVJiDIV6iOy/SY1iIa
haPFy1zUMcqtHSGmo0kad6B/rSa1CVLxfolPQ90yfYFGlFj+0thgknlaagUf
HZZt4eBCdYkRHnlOqwbZrzZMyXtV/iw9zeoMwP9c3cmadzq0OEI8X7A6bs99
7TOAa4ayAxQb+AnQ0eo132fI61SwWZvorFJqlgnAEjKGS3zVg75CdigZKZKS
I0UVm8/geNCDIdHq/adgF7/IlUUrq95nWzqGHy8DpDwbuujrdNOOr1sw9m8g
un3Df1QlwYIdELLIys8jx6eh4GN9jcLmnItalasjOIf8kQtTIDoym8n7fCfJ
nc6LJE8OF2ty1jRY8Mn5KbiW+fpmetshOe2NFEMkFsvK0qutRVdD5uFQr40K
jhVsaP7P6cXPNpDOodCPUazNDft4SXJlpoRNKQgyMsNkxihGZX/gqtAtCJsC
6DYQIx3EGDfPD9AyStKCFTsT8EZeWfE9MXmAICk8HKmSfTK1tAo6DpjJeltw
mHaehPq35Y0nSGWOezNSg2SjuRo1ufwwdmwKfTKntc5kIefOrxjZ0zIUV1/C
paLxHoHQ4tWMUH0CDuv4/uN2p5DTRxbLvsilzYOIJnNUwcqcfSC8iV9bJcnV
XKg0wbY+GsEDeZG30oCgi9YAtUNnHJmqv4JcEISZBnDV2BJXZvWO+YOvsjNs
f84xR3/UfMn7G97WgOtgxZIAsTEaDezYSU7TMI4BWTNEW7EOykDRjMiy4MCb
+KRHd6RXbBkKYfEk1g6V2MAvKaEErX4f8aourgRq9t0v9I2F0Bk6XpMHTFi4
6+IED1U9mlHE/f4aU3mODQ0OEFcz8tXFN0wCSYRxVnefwgG4MN1fPWtCwHo5
wGxCecnmj8QppcqhFm41kuXO/XdBtj9DCiZP0y4s0rUH6EVOrMeBixVQnmx6
C8QC8NJQm0UDhaeB/aGQerK2UtMYquYz1FUxeOI79kRbxbHLu8bfI+dUbXDP
fkIUfgYyjCL9ZsVKajneFIjYe8cOjc4YjnqVfs4/aD1m9OrkDHbOh9Dd0mci
JYCJk1uXaZ/uU9GWwd01/EiS4oSW3Tj+JjQab+F8Rf9EHakYpddoh6RYjRw4
+vXwYYOU9LnmRmZLCxFKtHULAw8Jdep76r04N9TOeNwlvB6NgCTYU8vwAtoN
Vq6XW3AbHynIesqBKqH4lx/hwXWl9tvvBSzy8FLs+OcF6Jz1oI3nKuiMxYTz
bahDjq1q+BDyqHig6ritughpSZy1SdSzrMEyioQH2eOVsVaxKcQj6O7utwkQ
ili0FBPO73ZPiOGEcDy5t2kJ6FWj/LiWXbaeYVhThTOOhFr9beITRBnfmlWf
2z8yooF4g4xIB6VYsVfUEhL9nsfU69WbD8+T2YJT3Hk0uW+V7gaf8p90utq8
E8sfNdCffBph0IBSRvZfs08/hRSM1JCMLGsKX1mEIn2RlUjHaHBwMLYIGB6C
AxuQWR01vPfDlpDilMM9KiSk/mHRpPjFdxvPC9XJbFtp5tA5xWz+ykO8s5UB
qOqroXTu8DMKPIuItLEFSXZPWCEoNLqeMyEHD3OvJqI9gdYq7b8bXbsGT+Eq
01WO3V1Iu8rNMf9fyEa87fzCDOY025Y8zK8VNPieutNDrc04J9XvLVov35jn
dLeuUePBMY19kJVjtLLr6sG0YyJrzTHBMgXTHMEAZ973+cvztOmrcb8HJcvy
mBBAu6z0QkEf9ciTqssAbwDZFWWd/NF/yhaSqS7R688U2GZwkkTT1crLF40B
8VFXBuUFnOThD6CfUzX+iPf5JZotaz3IZlgX4+jQuvhzWc9JCnXTsNL4pn5G
Xh4aKdQ9ADipcdlvsBQIa5FI+GWUp1w6gPI61lKOGVu6jt7+QpjTigBZyyQT
Ca48U7R/snPB11oZ1npVsu0Mf2TyFPK2rDXFkiKS8z/r1sdTfkySNqj9UJpR
9uXvblvSxig0MkgNMGILhFNi7eQXlfEYVrYzsOEWPZ97i+P6cuFi7CyeyZWh
ju6z23nxBa0ccUSlyYt3F94sO/DDN+9Xrjc3gqJntUw0xZuKguYywcm03Ot8
RfL41kzvUge6DFZs5vQvRiSXJML0/1NFAfSokjPvTkPQ+DYAfdNW+2cZ+yti
BZhKs9jfsAhmtBJanAwwTTnGQKx4pDmZKBmVjFYcX/0J9SxE5slWZzE64wUO
jOSjLYPsmqcphUMIOrECflJnAChBZIZqj1rtohu1cB9zi16TSWYq8UOmjbQR
nUqPjElucLBYLk3rAugZ916X50H9HsvcA/DMHZxskrptZ2AfrTERNJD+DVVr
+NP3c4z5Us8cjMUY4olwpeg/p5BxDGuHqB+O8rJjHdxg0ef8gRg2psXqgGHB
xk4hWJoZSoMyXovfsIG5IHek+LNnt4UmLaV8l4ilRWCVWBs323irrRPo9awT
vmCAzkMx8OV9DKnREiJztzKWZqSTTV+F36sEHD2rMIUbhjOcboIrW3VysoF0
zp5s37FicfhrgZRvfCiXEQqwCS4Tdhi1WUI1Qu/PPST9vdraYzrcRH0exqdg
YwZMKqcwtqb0MKzM5ReItC5DGw+EWX038cHkKyDdjVUGTO7JYYIkXvg+MVbV
R2M48mqsJx/UPMn+9Q2YT4niJlXhEUYj0zWeeqBT0bul6iWk5tDg+i2ey9ke
J5Wu3R5PgOMQMsMsLnLy9wlwdpEFWgB0LjoyR3bbIq5zZQ0UXU0GiFMYRZx2
Yobp9vlWhxak3aO67If1HzM4EC/epbveTBsCWi5b9M3+HFfbTAtt47dYF55N
ssOdJDkXrMP2JAKP8pmiHJrDhMRaLJwcBz3qkX110ixZA/bTV2XInkD9uWB9
vGkie1bkWuXUA6tEhkQ01J9sm4tNq7xlOLRpe+7SCDeIeiMpa+MaBf+jO3Uj
wdXiX4eM6IM03WMdYF31Ycwi+cS/UJB4lqSAiNm43BpEsKpuCuugibEt2EVG
BWL+p++TxqWD4f2mnhMuq/CU+Z7mPuXjF+6RcI8yQjRtdBVrblRZWgewV7oZ
SCkIFs/uKk7GhTRW9/dFI81YteugfKhOym3S6keoNRFyOGM7pft/8HT/00Bo
BPQtSn2SULHGQb8eMXjLT1+4NrSsQ+oas/m6gtNKKjdLDe3Cq3jOzWf2Pz9o
ECW9DUlUyuwmCM6k9CwUGPvSCiSv8H/IU35ZkThKCe6Y2jbPFtr9+qahMh9q
8bmoqKduwjXeLYdB8WUikdmxJhxqD0O6U1S9QdccKME8kpFTMynJFry3907h
yWV5mTE18mmrfV+NjWACQbaGzLs2Rr0Nsp3zXsZw0FnvoKuOVbohDKT3JaAh
VgM/QgHf+9yzL361zc2H+dCtCSvNotO469EpqZorUR5BvFtTMSzo3CLqTAfn
Z7BbY5dlonBYDXSFGIY4rsqV6hMdQqVj+obEzKKxgWaHaN3r9YrjfnWinHbm
2oxAKz2zxzo3nDyu/9z+auOkzMwBzxEX2q3V1l45m+qihuDJJywRIM+zUZss
hr+Yw8DQb8y/GX7w4D44MRzz+pEQdkvjAvYj+fpTH2MgvYoBL/eXRVqvKk0V
euz2b30u7I8z2dsFoHfI0NC4FsH4XKXlhOgu9oo6WC+m/Au1ARA/A8RXDoga
JKqfphYM5RIhc/6LXNPChlIdad9cB/8E1bDGEXWux1xhbaHVUuSvaXg0OOAa
ncxJTx5/cf1iyM5QvT9ftNIoUvnwfahgfiQjCzEDfiF/dMD4yMrOx9hkvQKH
7t3cfuvXK7tC90x2OYu9XHg/ftIkCj02S26OFCXgkBdOvNh5R3AmplREZL5O
uauT3oO1TugbNaa+4ii5i8wWCIHTVj22QVrL0Xd46VJm06ZAd5dPNkLWs/op
fhRCzG1c+zfmHG1/vt+ml9XQZ9CsUBMV1EXdXuCErvXXNOtl0W0LKzcrm47U
Mmfp6W0rDUeTBOcHxCyQ397OV2bLhN/lGPYfJK0dVBBoHk/s0a1EmVRQRe/q
+/fFPIVibghZfxFgKjH2xnFY/B3NBCp4zK9r4T9zMtAi+lVBG12/RgXxE+NQ
N36zf1tKgP+kNRejQcvvVHULfPrEuoTk9cK4KcUfTRr9hDIAPIfAU5BnoC4M
P/3jJn3ZQnSEK9nwUa5Sf2dhQ90oAYvZxUa46cxDI/TmaPqRlbrzdAOeVd+8
1pmbrxdhlc62mZN72zGZoGZxaSqZpMf9ei24RMsYBRMI6MB069q+DmO1MAC9
chhen8ku9tkcNs1//ykhGkmJucgMaxBeYiB3IUbrODpTOfh67Jkgq6I2vWxB
WzUk2mJHVgRbcgu19/yylefU9/qnt57e5+dhHMVJDMierRvA9csfOA21YXf0
ugC0qe08O+uXFb4T4S+je0epwQixF4ABIsv0663l1B8J6sk26Yjm5s9TW2dG
6vM1edp3NOgiiTpuJVsf7EA+sZ4NagtDkfwJwUSiu3MCpOMuAmdWx0fEkO83
0+AduOVcFT9winjrBaQFm8Z7TLAvpXxq5GJs6IeNAEPhHwT5Wi8kJ7N4SY/n
sL1sws2qxlNqYBhxRVS3wCHZtmJk613NC1gNy2Lly88kFj9zHKc+gc6vX2qe
CXAQp6gPabUn7bWyS6JBHffJDPbfx/bduTozBGJdiXxsJhxYbZwHy69fSDRx
ZMM77dbodFw5qsZbXkwHN/veE+umgukYj2zTmRBHniRaYCzAqTC1eIgwhIRm
ye90gzt6Q4WrdEVe02qjzi+51TwDu0Guf0QUA9XxKTDMft0R5fcPMkSrXP3e
18gxLUSmBgKMfr3N2vg8m/69PY3HksYVydcycop82p9e186ZIx7FWHyCflhM
rIvyaUw8F2bTNZESyDdXCnYtwH3HyllR4SqFuPyX23UNodYKce0FFLyJd73l
V0ySsVRwN7utwt7gn/vqvQ8VNBSCZcNx7Oe55QUSlV7JB0D9SCCkhay7j+dg
k2USgHs1C3OaqjRBUEJ1fx902szls95UQtfKjZ/lBmEGK5fezxxtXd/5cpTy
oOxEIz0Em7DOPDHNzgvcj9r+nV3f6L5dbs4d8AeK5Uzq0u5lia/dT3Wzqn/a
VS6Hhq/7AHwwSdRrJ7IlqZeT878nyRcrOLCXjKDpRUayT2nQDCh6RJIglJOC
QwlS1ovqsOOa7BEn75uegKZ8MBWqaWUXCJmTsegwB+8u1raeK4svM2YQJSx5
d6GmEi07kyA8RjjJuD9n5yQResuLgIcCxiQPondha/Nhol6e0oZWZX6w93V6
R2dHXsGDJSxDwPIsrGvO+RL8LvbxmqE21iczTcxYtQRgVy8bE5T9KtSc4Ugs
rDLuXVmak0kPL+5yLxUHhK4Je62PEbO5VW0JAwCghmpLvluzqFB73WXSqcvt
KHB17FFzQ2aFsjbb5p9Weh37+dy0z2VqTivuF9vT6ONLiDrBdXuW2fiP6Xvm
hzr5I3IgC2iG20sc/SvhEfkSHobifTfwrOqxXAZjgjmubknmNyVl8/7qkIl8
w8rEG7TojCYd56FQxyqELtpeJ6yIEjJsHe+0VMr2rWQaH6r+yQzSG1o4I4vQ
NgvaIwUhyhx5baNJICg+ME8mpCWk/55ytgJ0xrpagl/aDjoH4ez2h4jTvYKM
p85ENm602RpmAZfAYS+xipa+V2RbzI+hQbB+dallFRPjNrgXR8urrgkcSKrT
c6K3W8Ph9++bd5SYOsEbUr+j4BeXC6snxNCTaiKdcrruhtoZ4mLeCrbPVO9v
Pu0AdKXX2sCIUi1IErDO0p/TNHx44HphrcIfRt5Ru2w4XEGfdxgEuj7b/7EM
0/jOtZgxVvAs9lDNNn+Np2ThKiU4QKeIySktzrl7RFc9fEDrrlDXSUp3QanQ
ZEO+mdvR99SR0PogpAUUu4uHchYJr7wIvg8+sNFkLfYxzI8nVgO8R2nXuq+u
eY+4ANyLWP3d3qCZFevq02zXki8CTp9CDXeLHa/lrGwtkJSCnWqt3aMQnOqh
NRwQaqP3mTH/15EA7plHe7r6oEegys7DsvSOZfx5qbSXCSzPU8vR0KtndOIw
MR0xJ56ahcwva1E8k6SLx6UMCcc6Hje07FLVmbWQad2j8i0E3lJJQ9H3mkVm
7oCghVyhxz3gXVuP1nO0XCij0tffO77qgR06+VSskEy+XR4BKv6TMbCLMSWo
DDEKBw7BkrDGaam8TtHi2AA33Jcj0Htih1qBlc9U3mZv0jMaHUGVhEpBTaQH
1qRVmDx2MvgGHcKR8j9AYpERq3B38Snt5kWf3wBUFxPQK2ZQTcE7oInHN9oa
zp+xT/nISye1IL+60P9TqE+WGyZEd6cYAdU5QaVTGNMrHU4/HzGWajOzeMQ0
Cxjgz72YTJgP9gVzqFB7fdNipXDq2khLvUEht7U23suyBFa6wil/LPnNXIYs
otam0RsUbJtqskfmqil0uNJo0KJjgPiO93Y0pI4t4rnqpjrpTEEMSSrc/Emc
opDelUJWQivaQo8a71m5xBlZ0EGMBwHxz6VVcJP40SPMr53uwrUi4fllgaHw
hCzRAXmiojaFflLnOotayE1PsSZ35AGiZFygpKltABdCaA0BlYpKScaEkmlf
AIdDPBJxCbAOj9chkx+4U8IU1A+aAB75aGKI2tkZDujDdJcgWe8CQSf0Olc4
y0kWEDpXpb7oDG6ME3EOEdfP7gBGoyCOCxaaJJyBga53pELoBm+gXQY+rJI9
usAIWCBWKZ6RTbdJgKwg4TgpFAqzofRKjCdQ0C3vfIhRAY0FMYMlYmmA3CJm
JEQysxAq8H4P1w4R2mDfe3BwcKrZLt5YurZynou7DFw84/bDRmHsTyaoDR6b
SdFlFqsHxCtZQFtLC8uPkKFKkwgVCO5tv7W46taDhZCfCDT/H3rA7Qe7Zw3I
dBXjeRKochfTu8bxqpkmYagKvbN9+3suWQIQP8Nk/dy9k1GRSdZELdqKTYtt
NUEyNudRPUA+pVjCpFFMR5ovMQ02MPqKsfm494+w7NEglqpVktZLkdDsVG+2
kIP1sLXf8mqtENupn1uVQPtETAmB2jV08fT9sFdm1T7MPdFJy+CJ6OrtdbQK
7Icpk0TkOUDrUncrt2bWa+HT9LIb8a2jDwF8XK1XgPtjlcKich8mazaHXidC
wbTJxPD3JHpCc5iZ60ySfgM/OvSufrunwKCMyq/XS3YuczVcGtu6ACbTqZSm
3mMt/XBfku4RMbO1oE6HVkihO/EsFLwpMx1XHGY8/0KXlkqQ9cPlFboKfIcE
rMqZYqHhwMKSMZmOzeKmh+nhoVXYmEoa4Hxs+f7PtSAZ2q5Jn8wRq8UfWBhW
Ez5E0rTSfsf7RQxzX5ekUdj1Milk5/c6KfmlZksC/CjDIl6eHszVUtbj5eFI
y/MCrkkjptllhR3JnIAgwqov8wyCd8Fe0mzDAcjg9ShWKEfCK3wcOWE46spZ
Y2jGPArEk+jSux02OlCElqjM2lFX5FvZHgvepSE7/o2UuZl7GaXUTlVxkg4i
pJt07ren1NWN2+37y8mnl2RDXXi9bHv5gwsikOIogYa+27imofHd5qqhdUtq
lH3B4Tw2JSIZ5i+FNMFmcea/EZBuruQVBpurg+I+y697N9O2uHNlCncRXaY6
WIyrSS6PJcOS3VOwVg3y3d1ncsrxqlZx1BChfVElcpUiRonEBlIgNZUk9mTf
pur8MMHDhRwoYnwoThw0f5+3UVby6Nlp9juX2XqvZTUJ6Wf1NDuY4qAIZtaG
ddWnrTXLWttHq6MwP5l7ZcCucOgDC++qrIPtSwCHDBCKZ/s1NDM1gVaQxP/X
YNJAUuQuawxPcE0SwB1m4Mghw6QkZhreQN6HrMnL9Rj9DjmTraYG692f9O8f
RXIi+krrrUEgBErc9mduNpTp2Teb5CPFXc/2baYKOjWTyYK9LxZknL9B+eqg
28ynbDoROXrYKlHgTGpRZ7Yir/JJzy06Ak4hEiaJi6OL0iBFEKJC8m3Hn6YI
rGuO9KHG5AyeVneebRdmNYv4aTHN6jJVpRZhXYftcU9d+NEyzo5tvZ2uhwUp
Me3VmMp0NoYWFSofMaJ0rw9KscJWl79VTgx1zz4Xaz7tW0GulpT8Ra3tz8Xa
w565MRAOv+IGYNV2Kw6nJfnDciDOJMbxYx+3PqZy5ob6YMBEHAKWelFGgNzR
2BFmjruh3fhMkTTQS/KGuCqYONLlRNQ7DL3p1E7gXWZiH7gybZEdwiXppN1Q
5t/b0PoQezRbvT03yc082VfX32nkiLfok9bcrQbHvnGklNaoVlQChu9Z7w5y
OTiEF0wcOij1MClaM6nWeO9zm35Ve2NGGCAdqzgCB0Z2Vg0ofAKtnUCdv2qA
LgCcOghYPgThwpaNAeMmd+hHs+5gARHkISm7XxYaK0vLTG7C1T8596fdpi7r
Z5LtkbetGLFWG0hkoGSEbtYK8dMhPzl12/Bm9LUFtpRXrjlnnfRxmVlP6exy
1wj0zag6CxgzNRrIVphpc4H/hfpV0KClrW5xJN1Gbpb1pRsWb81s2k/b+/Mv
uq9xu8tkbQsx3J4n1MHWwgnalFKEBw1ra/CW9b/mltSLYjVfXc15EihnhPHH
+uE9n6A9ItGqNserip7UkTucDqiorkbdSCeTdkEeVFT4cdDw6IqMwMOZPmBm
8rygaSPXy4nrwwsszaDxoYTugyD2hQcYjyxYDv5BKYS5L3HWccmphLp0qWeT
5QtVZCtPPnt5c6AD+2o13+HRT5hmhGns4lYJ8YJCRMTcHA14k8/6z1Wn+eLW
WpsAkl3sbDUIYE7DHFTqgrSnhirFgvyqhcXQEmamVe0bUlnO5RLNXTG3kXH2
TI26exK13/LCJDW3xmsCSMc9b20lK5meH7SighDjeyNdcTPa1htTHlKgdOyH
B4OCMapycGdVWV/C4CTjx2iGZWx2SrebY4He6CpC+ne0bM2VCDW9qYhYDMcx
4FUvPcA/yJDJfDUnNPHLzcVCHDhbx3s0t78dl7mvjPWKm4rO7sQcVEhM1yEK
MCUVJOpJczo36pgzgHanYsCcZ7GJAiS2fSk35OHUPJo/y1RKkSIzX9t9UQRU
VvEG23ZbgfsvCrIp3zgeF0ob8xFNmDaAAAVjcFlSux1hs7J5xaQ5CYiCS0Vc
M3zGSpmhkGPV5k60i6Kaz4AIXFLbNS8M8iqeGIGTf5MaAVr8w8ACf0UpjRhi
ZYGNQs+IPJXpA5bFSPMZ+a36wZh9iIR/XB1mfzH3GDljRudiYxZPPEtE1S+j
qqSLP9JgNoMTrpeUWXc4VSU54QlHOfEUlH2U65xwUUqPTFKWry5w43YpEDuu
cJKm/J1f2BdKdwz7leb+7BJmLN8As5VR0FiUSJ9ZZeTSm9jx2LepfkQCCu5H
Dfl1+RLVQtutEbr88xf0FjQMz26pIUogNHy5zENh/fnpiHI5h4aBHAqwI+DO
y/Ltl6XNYX1MdfjLikXh5NhBJcasc6qYVu8DMFqLzgfycn9HRWTTiPAZnRLl
hjzjtSco/ewtqy3vCqTjzd97iWiKTMqWuqhlQeTMuQBkvKOg6HpZ5LcJ1BIG
LG3xjf25BKFLKywnDTNjBwBQsGk732CkiqLdnL/2l+uE12q+nfHFdfUEBo99
cQ2N7ujuPkANEwkQWh1d4L9JCM4T349MsAqRJ+qA7yLmBFJwHWQ3tXa7q0Tm
RqTltkNKnGG1sovj0bxU9+T1udFM7JznJKliGrweTJx+W6ZIoqlQhEMmK1VH
F4AycXZO+A2mUCcXWDUBYR3RfkXHI3XxkDb9ibuePWFaGa+aPUnrhg2WPili
jNmzARWudfqiwbsmWzn+l3KtpA9R5Zs1Ak6ULMWbcL6ZmON+0UQcdLL44eri
NTMQ/qvLKlMAaSgasrPRjcnSbxloXZuCBFN+SHriCdSD3HFPtJ9nlJh1aO1z
vUHGNAqHv0oZ1fThtNBa+aJ1zC/SGpbJIsvx4X3prHEgfdxbkAWprJ53jW2O
+BhM6NZK+JyEjpchtGPzs3lYFAmmZqrDMw5Qm0DCIwhgsZ83z8wYJXkOo9pD
zlQ2V8ZxQeRhDqqjNDg7B7DpUTY7m7pD9qc7r7L5zANrgW6+tWnvE3Hb1hA3
JwzmRQ6l9KEAwu9HMo+4djyZBltJ7Vkc02mnIoWj3N3U2qNh0fzUuETMJ3aa
r6ZSgPLm8R4VDWESo+mrJbtbdc+3XgvRJXdwxOhDp4+QMO9s3HW8PeGY2zEG
rTeDM+b9FrhhRJaZ5+nTinJZt9Es5lXuMhaPL8XgPeurJkf0Un1SZ8Bhcmga
T4Rpwq1EnNuN+DPy/JfLRMHMqmQif0joCBBRDLhKX/19qhcH/8d92SBCqVLc
4W/R47NjozjBZKtG8Lfis9RZGtoMU3LLb2VeXCdYA+uV4kb5I1pW9x9wDWkQ
BQMe7MP+ZeuejPy/UjRUNHf6W35sP21t6Hhk9lmH587NvSiM72wPb5DX0LeR
Sq23g0/PJBtX5fvr3hrVBEXO5EdjiSk6gvgFMbF5p7fq4PkaAVmbg5PQMxSP
xH4eVfqeW8//O8UFRzRNdDTiUpBnYSIgeRg3JaQijL0wTWBTL+Ve/rKffRkD
E2hhmQRCQm3aljZ1Gv7XOcHnDo+uW4q+LxZ2rVAd83G3h4/au8/xGLlXW9LB
z35LaqCu/TFG1CPkoPwSklKV+O/2VrLg7/r8Nl7h3u+7IfjdZCxYOZqs7HF4
J2xPpVcCEHohHgYBVpwBmILuAiLSod0k1B2/Qp7rMNomqI+TmemylYMwCXlq
n32LZSuQo+fAH1KKe+9jPmeTLbuEX2PgOsMrpPx6hy+ZAqSIxeUVU78YWtHF
degE6CX3GTLn381q4N28s0EeDrRlowVIJxDEVKWtahRH/ew0zU8mu5mNOzof
Y1/cVbhQTogP28mSkJyk8zPAxFkvVSe3AW5q4kqtPQsI3+je77NOFbu1t1jm
UqND9Db+FlBJnVYPeX8MdiGmPc+/E+5mSBCFxJ4woPhKN2aJtvQLu/AmlhsT
kzw8k+RZPMX7VccSJnhEXAnD6TgIg2VfRCRCqIzTem3dIlRM3b+uI6CVUIkN
xJw6ZVWk8DCzGb3sKmxE691dreBbf13+wJ8b9eaZtyZH1hj/N6Bof40LS1ZZ
2Ss4Y182JXs0aJ51084hs/qSGoXnEvc2SdxThnXDlSMyLK93pJCQgteZwr7D
xdS0crneLSOHh4Ih3vTTAUhym9Vh0TgV5AYmzTacPbuTlfKDNkaPpUveVwnH
2LZHSoeUReNP7D/hZtSdXJAkzWra+nwKEKQtdwFq93/CZdhFzHeMgM2dRGDz
2JC7K6mLgEmDkTk1zQhAekSYY9wu5/2Is68Z3PRwjOUtTGz0BXmja0TrZKsx
sT+vOyzQWnaC1rtXGuFObG72NURqMREFPe8S0Jh7YpV5mSsNGLD8YSbrFEQ2
LgcMqpvm8eqo3y2M/isMCNx3mg4MpDKa8jtLwKgf62uCQ29z5YpUkMjoEmen
kXl1MU5IkohFy2094bpb+fdfBhNteKewlRDJuflO2wCK3le275yvPnh+McBj
yW6tPhy8XrkJQFEAwyXQjCtKH7jb4iLQ8d2sx4Cr4B8i79LLvtaU+tC+uRQ2
pzE6Dwuk3DK+jeIN8rFVsKJ/8X1cqoYL2bDrexGFHRQO8ioKkd2h8FB9U7+s
1QTyNXyyLcx+54D2MF10GRMaXOxQ9NOR3v1FuF8+uC5WIn3pfTAP+DEL0put
VohJTANh5J49f2sOW/xCPgTQq8iQ5Xq6nJhrxxR8GMZjETXaLoBo82mX35jv
hNK8v0VHr9sKsmLHJ5vTr5pwyZLAlUiPRURnif4K448XYoZacYDzEJMoUYKl
TK87Ct7hfxsXHdY54p1NWxzdCROTOw18AkrFO2Qx/ltH9+sORg3p1swVlBtu
FvSdJblNcIJFlNxE6rA3NzLxc5GuXX6SqE34Oi6sQsCNCROTxX3oZjRZQpd7
eGIfFDkiPRlZzOxGLXAPWH532chbeh+9pFBsaYe2ns+mpfSP9Rv5Pu65dFEy
1KQRfYIElI7iXvkT7kFuj6LodIW+d2qEK9TRs6NEwiuQDNsAxcM5M8vYDcg4
e/On9YNTrlsjOZ4O8OW4r/NEQ9/+Y4TAR/5PuSrms4YAZtPy/NfV2UOrG89I
VSC6ZWLxwulc0vwgAvINSKGFX6S2WDjtByuO4y/7wc+MvEJ1kgcOp+RFnHRU
w3T6q/sH69562JknEHvCvoe452lcr8opsxCOCiqdVZ254CV7uJPNxaK8HPVd
J//XZ3zgKzB1J40L2r182Li0v9XmnE3/PXxmTMAUoEboyxtDVNxjlaSceJqS
2KnMg0g3A4zsh8QnOGVIgnTIntU2abwdvCDzW3kwIEHwQ/P32emBeoh1GJIj
GpGbt9YUvhkRXhsRPV+RTi0MAQEJgmhnN8lGrNKSHtJo63pWS68mZNmpLNm0
mM/4nerw+oXFRFvhAHlhbX05OLIDWRocjA55a5rW9oPZqHHiiprcCrM8vCf8
WoEs4uY2DjqqsxQZryMFfsVziqpmt2YUOnugHxU+f7EsA8LkHWtAd038Mq3Z
BTk+CqHvIHjlfNwHFhSd8jyayKkOdwEDnI4qB4QvY5ZParJOKgcYEapKQeZY
cDn1BRYsfgRCae/DbNM1FNGA7BSsKlQBw2yy9QDSEG1ni8TbclNUt3mu9tsf
O5vjGMl4hLaDiZCEE7onYdsSSvjve8lSQzB7eXtz29bpMquywWQTvOFWiBXp
8NYT60ZuFw/5+DPuvQpHS+AJ3gP+//BCuWV6Fqan/DTNfsGkifJcS4ONP6ZL
aL40wvDqwTYqYhnqtqbHk4j4n463mV9KYUZRfqXjfKhXur/TJfSh6V85AYt/
oGzsy0+dpyjiLIGNa19Ujp3gSNHAod/EQ0Rsya1deQflHB5LN/ffRG+hUVjr
8jtDfVlWFejsAH6XiVVfjgl2uUA8p6CHD7oNigS62CceyXCqhp01cF/VeIqt
+kU1N7qLfNVZumdfdhinKZfXXi/n0ftcYdvsfnCYXrNq3xGxOOwHu9rUN/Fi
8Q+DSS8hIRkOowa7YhHJAYlfRVo9DVv7vnVtvAT4HePAv2rnwZ5L1hSFUmE8
GD7dVYxB3cgqVu+OHMW6iT1gPwjY1FDphfayX7wFYz0NbM2sAlDpyjavQT5l
8bdRWlkn4lMRNvJ7A2MDfkmnHx4bs5nokwlh/F0/wVWS8y6L7S911JtuK2Pa
Jq0Bq6NEGKUM3l1h1mvqH82AZqHw3sGbY4NeKxY8DtG9UehxycLCyrrNqBNk
nD9AbIpIoaoD6lUtDRGceEP06KwScCI20dmfp/RaQzlHsXByDitaaYeka/Wj
b48OPSRcbSwh6qcrRpQLNwSXNgUpXnmSMGOabu8J2KbU6JmxE6qu2wdKiwzQ
0pJ/M81Z3E8yQyly8lgUACxZCRR/wb3UoI9b1iWmYpBFa3q6UzVNOSLF07ZI
hgIPXmniAwBgTkByy6NK7Y8Vho+nfefw+hy30HsckY4MWS8qu6BuRlnWs83l
z4p+OXkQjt//RJxWEsSu9HNiEKIBWJmF+jTJjZwdIbPRIxVAoSF1P/GAEQ9A
9adUG1ZkNu/8lso9F171Fz7hLDJ40GoLuugK4voF0ZM+RKGcueVb+Fi1NBH0
SIDS+Wctc/ft51loX5gES8puoa20obraPzFND3OqHgqIpoc4dr50Niygzoy8
Fu32m8m2zWOe8VZneGDrK6VDGIk/oxtYmwkjGh7eUwS6oSuVLIxdnDtI0ODp
3PONe6QVCHJ0rl+Z7hpaHmwThvAltY5DtXitbpswBLJMu3wEAKoiONN/dscn
saM7edDNwmF9fWwon8TaOJb0LRn2V45mpgdripBS0KpA1KbiTUVMUVnQ1EKX
ttwa8vT6wh2YO3Cra40iLpidcSXxxwMRcYobIJPmZ7SZlS9O02kj+98Fm3Mg
6fh3oaxO3U2bj32z0kwsvH21g5Nw1n85CRcBczcK73g4Rwz4kC6+JIANqIek
kBvoqDX3czoSWcwhRgYaRQN6pwyXcOM6WhLqy0/vZ023GyxqOdgRXd2KLYOD
+YukLgHh4U1f8jQrCrDeBd8Z6eLiKYwyhVoZeNHcs9O195I1hvJegd9szO/9
O7dE5iS0MqTf9FjwRfCDKKQ/K+eZKiIC5fs/FGWxFxB2sR2il5jfD6Z2vDBq
TqJJot+U2VqjY4K7XvL1heLg0dVSsjKLXI2e1Vrniq3YrAJvo4LoygEBWge/
7cl2tR+pPFM8b6N/3oWZya/C8L7IrLPPelBQinsase+lYnHXrQaUTfyhslnH
fZdJZ2VeZb74m1u0oTSu8QjO+BHR2KcEcxzmwrnCm9OD1diP+AfSSzoQpf7G
9C3v9DNYm5c9HMYWwYzQyVuceGtWZpYmG8y0B3USYHHU31s3don4n0sdpM2d
+8+aY9ItiDjyzwGkZq+Pbbr6qTZvczEynmzUNxUb67wuBuV8knOlTGMIBUgH
My+wrIGuqJXpREOe4FF3hMbnDLEeyS9+PQImTiAvJN5LAbZjy8IHZ5ryqqBg
uA0Q8QCX2kmb/B88Lo7JOVqFCL48fGq2Lh7437UAixWLPXq1z35psAEuvCiG
jBid0AaLmc9bY64pwok+mtOIXseVgeBq+hEXHA3etUX025hHm+uVidzZB0+O
HP4CBc7TIPSntRdVUIByTq+xjiEpJObNFtDOBDn+jQJn36cLJ8BTXC06TFqo
i4w7eu+yYAVSSDHNDlG+f2BKkuI7TgGfo8GaBC33Wbs7Ikhv6cAnWSFNKZZe
AWDCx7pKEJkBuJs5/V+7/RwqYBxwvTyLPR92cGCVeREtpwc5NBLGvcAfAkJN
+DrRNsPH1bZZtlxY13kVpU0owYYkcmeTRZaa747+p4MpJzQdAlja43a6UVe1
eSLaPrlQhXi/knX8LA+OiuWteGkVLmG1w98iDl9Zp+LewYVyFGlQagmNeBAs
7v4+ZSZaAkWYVne14JHNKiQUJOaiJubPBUFsT80XBajDjIXuHno7pH1lAbai
EJE6Cvb+dFnPTulosThEPSGn1R5LQ/NcdMv/gQgdOauuX5MOtCR49jTzDf3r
9pIv+DTQXbHjp33zz6+nl9GhosNv9RNlAZGF5TAWIM4RUwzz5UhBU1ZTV54f
i5qI1cnjESrm33ObAMdrcnYxUkBwbPzayUtE46cs1U6V6LQYuY2RVisS76th
INfaxZA5Qyhjet6Vn4IHBoXSmdZC2Cfy8+i3fvp7BsXOwhjhEzRrtj6Fr/+6
toySrHEr5R8qsn0suSVuQ5p2WlYlWsZIHqsyn+B8QFZF8G9361kyNjeJvT+c
sayvbkd41iWThKDHQqvEe9sEELChcaB2SOQESsxZOfoWLqgWynsmggxmyBHX
Vcoqepp5FdrNKJHyllXA3bQSqHl5OY15qkGq3S+lC/Qw2H4Q0lOYbwebKSVc
zHVB3IamhZjcKxT5dhQWMtyG3zAyDBPNx+sY0ZMrolVRrNXBDEnc0VfhBIO6
PSxfJthfa7jG0ZdVSXyftfMOck+E+5GkBMRviz1q30F69iZCtwrZGUy0d2ZR
rKGJnlIKzt3a+LVoxw5XpJ/omUmJjDc8XSBe49gspAX0tgxmAIwQm3pRnsFO
GK5fa0HzZZtqqqw3XKNPgJh5fft84A2oCT2q0k+XteZSxLGY99zYrqFCRIa3
m2ow7M7ByEVh1YGFXHI2sMBg82xFxK96z6N22XAWaD3qNfm7Vtay1szzIPLp
mhdnGB0e5g0utjJinlmuKHgl79JhhwFj7r7gs3v4atKorGS/gzUBHoF0QyZu
iyWMPwZ2HxOAi7HVKdgp4KZnOvfQw3PsgsKtsWew1EzlOiiNaeBqp8X8PmBa
Xhg3wtlfvnC5jBQ2J4BUxuQ820rq4w+KLjAsgAlVRCMboGi+IKscq9w6G/pG
T4X3lpLLRkD+u/BQF5xxmrff62HMIV3P4DtxOUuw46rZJZw4xusVhcO3MeK6
oiJ0VJxg25cAZHPTX9RwGV+ZmmPPaQ/EiONNGvqpAgQcIEWYvV2p75Dx5afB
xqlwP2vU5RW3wbT49JABN1ET2n3DXQzPDr3bkOPrm/NcrLFMFl1DEUQpKk9D
P+0F1eYD6txfBdr8eqjBaEQyOFGTrRBBqa4s18yPdYUOqDP4rXIvGXiL4pby
bDMZ10PJFb9JfD0Fhv13sNePGhlgeL4FLW4rrN3kPFnNMWJAyOF28reAMMZN
zSG+j8LL5MiASQ/cBR287LhJdkfE65FrvYKg1NjurIJ2AVMEWETVQ8uKjOZm
SiUad4dt1kytcos85geBM9MxRowy/0JIgp0DhvLUiQ5Se3zbtz10vtp7WavM
/9rcc6Q8dLp3apUcMKkXHDfFg8HdCbwBl0BzLroU6GmC/uLpjoWxjRNFazjz
/UKTtjPkcCA0np2zg6VJGQYc4cyHfDoOo3yXI8REod5SHVDYjqtaWlvHPy8V
qYgM869P4y/noXl2gNnrWZ5dJTXTRVFYlmwK1FllEPHzSK8gxSiXfjS9k/QQ
ux9t+Jmy3j0Miob/xQy9qCi/Gq+1MjqrBBOS3Fw+dIWwiFZVz8baGdE7/VIz
o+PgWLu5u/Tz4qc2uLO+8E/cz0MRmxcpNPqRg+WpKrYYAaBZbek6y8ApzRXP
1Wqt/YCU9HJ1CHrnKjK6K1aM/+utLPpQNkyuaOqj/RKMRLuw8BeWb6h+aKOk
B8gVcfDP31/5Xt2Q4wm/VFWXRdghogmym/M3uDVt2yfoieen1dspE+diKquE
qnOvoB3k9zUY1qUyLpek3bZ+bGqAn73Tziwo3G9AqK4hnXr05bhDa4ecYCAF
dsR9DwFsfIohgHQWWaX0sublqGXjwTaBi8HExkLA8C7ZeeA6BYQ/z8PzbxSp
dy1yFJ7sXAaB9HJkHl38ySByq5lXeU6414wsBeOp+RfRRN30Zdqn0hkhE4QF
XRMfAiLF8b+LW1D7+aEgcsNa9ifXdPe792cgfIk3hIeLlIqnDNlqfuLVYH6b
m3bLCa/yknAlt0ExeZbYMndXbzA7I0xLw7QdwVD38YQ3AFZtsM3g5Go4p950
Xw1jsiOLiTXUe+Rm2vfaTD7sPxycgAE+dGVBYI31DSpVw0HXAUCLw/8LvN2H
d9+a/BSiNis/E9Rfz3flYy4Pn9IB402HjoZ7ylR8CSzvu1ZgkC4c1lHYXWYi
0f2lRTmyKMf+fsGGIDSV8twz0VGPgnsvXn46ocP5FqKI2t7BnY18KoB9Vnby
ycYGGdXfUYOLr+Nnn/n6pmSdf85D2GfLCGk0hJroemOOAmrahgvSC5jPyiXF
kpxSC6t+nSeTFYq67+bTKO95Pnb08aAxyzBWyd9tkqkNYzR4cDlFlUzKKyYa
AgwrSYOimvKBD1+DWbIeW22OKYYCyXJwb5CjSV5cZdN9E0V2Vpw9ToJpLC6u
ZKQUjp/6SQY7kwMpdnkEqfevdxWLsSbiYipVPQ2GJvCLd7N9/VlmQzKOW9PE
YRlpNQ8xrLSEw5pENky3fNT6qn9AIOOFd5lm9hKxg5mNaASkiztZmWjojLsJ
73LJhavIeeU1wnLKjJPYt3kzAwMczu1/NVUkpaoG3Sos3kOatYthJ5TLbAoF
UEt7V+AwDMck+bxfsoFTE5V5xAJOL6Y0eCqjbXxIfned89Oh9h816fgOxc8O
ZgkpEeINF1drJa4w0zijPMxLo5mStDNhfjMHEULLsdVw8vODXy9t8vqx9KL0
4kn4xMPZOLIh0rDfIzAvn2JS6kSbIUPriXj+oi2x3mvkPi3og7QMIzjt8De9
X28pMo4OcyTDSXH2lBIpV0VitbJGtgxhfPY5ja/Lm05MUg0jiHjoSxjBMhYk
JfZaZvR3aVTmOinCIpB+fqdvYV7KC9Vk33D6l/UymB+j9qrHF484MiUZ4X2I
l8UzaKaqlZNa1uCPFmkdbpO7882IsnuuTvBXoGRO7yn1T4JfSlpM5Wa9OwE/
HRa+9mwcOO/8vB7xEJ8UfRZJYaAfoP+DuLxrw66b2BU/pF4jm/9cpMad2udw
yKzxLaf9JVs4kMke0aPoRwUa2RjIcFDptqBq0ZdqcXFVHcGc9eJwKuRmjnlo
pz9eiw7embgWa+KuTDB1l0vFr3/ho03LNwJ+wSC9UjfeIUlXP6wpK4ChN66g
nOu3TeyKmN8KhcG3sfqgPAgYIgCO5G63zehroWUrIlh6j8wfZXbPF1OJXvkE
kVRZus8xJwH8Qu3JM9daN/9SPNQ+AINOf1mL2JTUkgaiHIpIaPnytGEbrBKw
k7FbMZkhp6Fs0by8291Q5oHuVQKVNjnQlySspQRKiLuNHnkwVB2WRGHOFfL8
cJIpa88jsLW+t/OPBDXSw6lrMCQkdmqj3y7JTtzh9q9IZAgCNNcvawslfLh+
i48mWuZijGLBNDDbuysrlkOEVaUFxbEojz5bxugZyydhNlFK2xukX6tzsxv3
WqStsiWyQKu3WJCTw0/KUx37AkMpNI9aLBVCCu2qrMkIxPCRI4Bj4g8y9wqd
1xho/BRZvSHGtI++PjU89ns4fR6erkNAw9i81aKKMwgo7yD08io5jQ1Mvebn
Qz/JxsuQWqyZmlZA7Twyui+lSfPff3Vyw2cYd5shta7II7kSuL4IrVZvguZt
PKvto1uMIymCJk29gW5fpDoWQPx9o+kgfVq3kvKn4v1v9YdCgQ9uUt4fbghO
YkJUZsWiMoKGzix/S983kmXnr8LiKpAtnz8rLyxM45IjwEFkY+5TJ0K9Vfol
vXQnFVz5wsVAWSKqOohY/DmfoN/G5aZy2WkqoijUpq4wBrll0Npuz8bVZAqE
3eIzEtveKeiBv8oS7YR7mf03PiKI5wgTfLNlPeyo9lnBiOars+K2EZ56jWUr
OnWBM2s3uua66TET9bm0PHmkDscmeZNrfPMlNGZz/udhpVnWG8XMk328HxGy
KudOsIv5nanMIU9Wtv8+mUBK61uA0Ab9O6JnXvu97P4THdNYlvjDl9GQ1fz5
geyAFGW4gXGFJlwWvCv0lJARCQ5q22+5PprbGIOhXAnsKeK/XaQjQuDAJIg4
iSEDm76dPAsyE06ZTlunwsrcuG5jNkhQVxr6kMoVH5kViL9N/q+Q9BUzYmFJ
/fphCAzKLrEsVgq+SMCDsENNtkm4trkiNE0oUD0reFoYOeFqpHlij5nfNBbS
W76VMOSjomFcY6fT7otMHahUXCrQGBGv31cmwa3Y2ebaO8blgY98vS/Str3q
280R4+y78XdWlIOwO0Ruijg9x0e1+E9dDqMARhaBGW5xsI2CQqMuzlLKbnCC
dimRbISB4YEZXxShA0u9uWkIr5LXi8EiSdhAIOC097koO0hwzNd9DbJ9DNCf
oRiMijkACHKwEhki/dlFtgSzHwIR65YfSsWOdJPw/PPx7Cn4A/bxTQQbwyzM
ohZVb+x4eu7N7XxFzWjlYVdDxHWrZfiNiMghs0yBtsZkC9ZVapbRabtnk0uM
WqsbQCE28omKT57BQ/Ie6tvoM9+af5CFJO6rCbhnHvqmgkZ0p1/5KEr7Pd68
tkv33MpqiMWMNETwKs4sKE14TaSTzrWlN81ty1T7/W24PkZTzyPMZI56nUT0
L0IDfQtGu73YAMKvhQnnIc4yy6+KhXP0vPwlKqXD3tgh2ivNHIG/+id2P1N2
BPOu286ewONNUlcG7MD7Ou/8l74kNTTYdiHMmkR46I/dAaJ3UbTZxMYWeYM5
ev/w26g2U9sqhKllvfVYDqsRYI/s67Rn+508VKY+YGEKdz3kzy+iST/GNi9H
SslbMNpJ/WMwIoneFYid58M9oU/weeKLBZ+tB5lk8SeCmf0gsFNQp2/4EI82
qIA6rleELSh/btRA4eQFS7ESmRtWTqhlr1AYX1um+vcLWhIGaQghswEk9LMQ
N8ak5MhOs6TfH7nMk/lSwUq+iB9vgZxZICvyc/VxZ2D6+hqzsVVq0b/j9w3X
M7iA6CfBq3ygxRAPZshhnuOIMfZa7DhiNW91xAo5Ggqidy4vKcCUz5hl42aY
Xw8nEX5ezdpF2D9ecXV7AQXiePg7RKwlhPOyTW6MOkaeACY4X2YvJMnnikpr
8ETxCro/IqFA3fBH1jFP++XUBSW9g+1j63bbkeXsOjpk2dkl73CnEgWSa1fj
Fl0CpHr5gCGa5ENLabkxbk1NqUhutDnsDEVN1M+00JAAC7V+SSupKybaBglH
jF1dXMIOgYMnz2nbCSd24kfmzXiivEHY5G4RCfV9T1Hzl56n+6UomNdmk+9n
1ZjFD1OEJe5EkNssWSlp7VFo0Xfo6Ht6jKinokIcn23nk1jqFXVz4Vcu4OfB
Zpr3+SqzMNwzPEsHmZL0lYZJey5rMNuNYOtMgbF4wSCTptn1FDe5/6HGbcis
NhMAF9h9VL/+zCl3hx198evLBUzd/Yvm/4Jlm+ORFHl6GsVzHdvdWhKrV/zS
cPliQzL9PsmFs0ss3HTIHU96qhN5nIz3PJIAFaEQkbwWzHhCwK4Zq2fYhBF3
M5RWOcn7fTDG/DtArdmURU6LNEDyjijwqNcM0M4EhF99D+dUj8xEn1DufsPb
5Oi/bDuBvCf4BbrvKF6/uVGEr8I01jPNJU5Y8o5cO7iPbA5hG0KOxA0Wj8ub
KOZWUEWu7xWe7W3jW6/0ZRoD7454UUnNXJqcqo+SRzagiXKcmVUL+udom27G
UWCd5aewqfvqgPYEh/XTfZiZfDECLcLGlvHQKNxTsV1gDiM3Pn6LSfrE6scG
gpEnw+NNJzn5WavkGpxZsXp5SFs2WFZvqyv/XqJkDII16KB9iZNC4J8haCk4
FHNI20WnYCPQggc3XYaypDBH4xsS4ALRjEGGqxnVG5PQkjxXUGo6dfqpyF2I
bz5yLHq07UqyCRNMolGADGZk1i60GfieVmlg0AARRhG5Cbr3nxeTXbFUWUDi
nHTEmqkWJ9RruCamsuufFKNndgWjiJR6fhzlEsJ3Zl2SAQ1yYG82o71s3dhy
czh2rm9Z31BPbeOSv3Khhm48a5+9ckbNcQ6FvxJb1uaVrIwIJWb5J3MaT/YI
m0Xfhvb8PiGYJ97Fs4h807/x3hlPzVcOLzowV8idxWu3AWy+TeOnr5Ap2Db3
CsAWsSaOqajG0oEdGDgw+h8V1lLDOP0ovxSJAdFt88jSVOHII3us+C3Yti8i
74XtMyuKFANJFSyfNREu5XWvXUaZ9KAsoFic6U8gTAvrFr/rDHn4mmPUlrEP
n0C9nQPa3DR9rGS4DIPpNGCAg0uQ6Jt25saabSG2EVnZfhUlfY4sJHBxijL4
kNG/KqCtdmErq0EN6yLgIqV1wGghqdTNzZxxP6/XYRnSjY0ERHFWFR5Xfy4E
VeljccCpe7hK9fdfJFvPyxdm6XCuxz+zJfZI1S0XpwiHX9KpoMevBwOEbz8U
51zzKq3PFyNp9R1HoqpEfRJuTEdoN7rUOBLu8MzPWfiYV7h9rfWGEAu/4G6/
pHeyyMv8nr/9/97QBfIp0ANTMtVJuO5NJCAPn+4VUlSxwsJl0StyKKdgG/CK
Db6pQ1BxJ/pXBWjZ9splaFIWSjOT1BgM3xcWNzmu3LY1E/Seo5OmFskyrI9Z
/XN4zCeTam14OUuMVm3UUV6aBvUIsO5WQoOb9jihI3nz9fY2xoUBRXB8AmsC
nvbYDtV7cDgTcboIFUrljSI1sSpbIoDtS+/ralCyaoUZPG/pVR9QmkQhuec9
2vDM2mhF5j3CVIrNrN+nI2h4+fRlith8FmtNw7UnZ5REljgHs4NVInyJZA4o
K6vtRL6E7ZttT8yOChAwRNTB6FFI8gHxLRzamOpzkDwjyAf4C/uNLwGlDBiH
XSklxAGiVQqDxDz5UnB+V5mKK7uOTo2NYYskqQXpOvHs2/ikgt4rCeND1idf
R2Ksjx1orh6c1zKV2VqupAPWgkgrjt2KVoA7dtDvLQ/J/91La0jVSP6TUrtb
Ycif/twBBju6bdsFvmWg90/fwb/6852ChveCqTVroZxnZo47cCHWt1e15dkk
g7d/m6qNDbNRRCp7gkpqkEQkpftSxv9xzdI+E8v+v89n7170XLinxOmVmKl3
rcLulidrhxGYdwqv86jC17MH6OimJvd4x68Ipejr1/H67/jq+jhGKGyifuAC
MC773k4wvC5PTaDsZLan0Y9ZglvZ8vuAg2k7fbaVoe9EDEsTM6yEYqxnEMO4
Wp+F5CJn27vZwpTzShMpIe5P0FlAKrob9nxr6m5Skbfh+A9h2oH3rWYtxvt1
4+2Bi+7k+A2Rt5aUIHJl+7UmtAYgJQ0cIcspyf9jpLvscMiZlfrSRdW84TeW
XKq5EfuduTEMw/zb3G5rlyv0VL5vxvny5v2QEHtesGwhGhLzz0ZFQCSCwoMa
OXnlps1yaTvWRDqIOCUtJYIJKarokm7aRU1dZdNz82m9UbjgY7G5OL6iKoP7
UQqlco/JU9pnMzrlZcKS3k5PF5M+HvFQqn1IvRT0WyLRVl+5Y8QSXyQ+haLF
mzdG8SQc/C/8vAqgAaEcghvvDOcAR0W0Go1MUPN8tL28NhbbK+VG6DTsm+HS
CsNSQyew7+iTRiHskyXD0tN2DdRujyXm3kfW3AYs9T4Ce+/T2IJodTN6QwFN
zTndVMPaydKH8lw7YK9pqnLo8RPUuutH7s23IUMVkv4oVBhMuI90c4S0ZxT6
Brnfdf+FyLfErSPRrQOz0NyrxPwA9pwomo/9/GXKS3PU2ZISP8LhzW9QGcVZ
ysFrPi4uvZX0nDPvNunxGDoOLP/zxj68fxxRqXqVBeH6C/dp2XDPdYVIv6KS
znuPfIiPyb3UTxRIglGSuoIQdSv+E4dqFyQsIDtIm6kp/ffCfNsb+FL7wE8z
BQV1Wl4RkD1abreW79zOUXC0wTztOD83q/bpOYQJ8cwN9GQkjuagHoC9+rVp
QUTwUvi7xzLSrtSqsvSBbWakkk2V+CJVm4aj/EcSG5q6i5tnLAfJIgF9n6lN
WI79ubmBFL3zGAlX4MT0Vr2zlQQqlGhIx6BrJzlsshWkSEQF8x2BEYMLBLiS
45ri5OY0BGyRME5DRg74qkG/q/LEaEQYznagrRGlOTagvwZNA0sMQmOgE2AD
AR2NsOb3kFvpjnwwqJqmVPNLjdCFxQ77BCgtm7YHt/WvewlYfKPowmFMKjXg
J+sQMtML/tvuu+0nDCgv6b9y74qhFJ6zbtv5ccZa8rvLO3gURVTF6D4Zykb3
eZc+eztDnep57UulU9oTAtRnvrMrj6EtMaTHtwc39yAfS0tpRzuETZcb5tkS
H8iCi9apDaNOecFsq80i4PqMjwOtyGc7ws+Fh8Yro0DiWup4JpOcGsPx5MGE
RhKmRn177lLr/C4msDWTk3umqVTdSi5L3g2ISx73BVO8LXXLnN3UU+OH4pK1
11XCUllxuhVdbhZ8IxIsbVmM28Hnx7aq3bXBGJ8zILvRfK7mAyt6ucvTc0Ix
j/zB2a/M8GPy6aNoU1u8b6O1aqN96pxyXy61VLzm9bfzinhwsB3hJtYccElP
Vp+3ekM86zlHjmfbZe5sjf1poXSHF9svqpEcvNFWuAG4L5JaI0v3yt+EEJmW
rffUrAULsFr1JnotyWECVQVrfR3E9jwJRyeS3AwqhhF9Vwc3unnFQeMk7Y7c
N4rwqhcmbMliiSARBs1v9Pajv4Cy+Vnb/Bh23SF7lIvzha7U68saq5OExgBP
H1oc3ZCHGR+rbLTNO36Ufxix1Gue62OGrOZxjoK72POqOqMeoALBQBDwPq6/
3faaXBHznYodQveztrIZqOMn/X+jgjH1IBbKz4/+V9N9vzJSuopa/Azlqxgw
MdmNq8IJsYnHAniBIn6BsIwb87BAZcvqY8yVVWKBzicSerJi9a4g4pASmX0W
xSIUPYcnoKywraFAcByED3kKz5dK2cY9usbY63TYj8MeWXPbd5w8hELfPqCh
xZwzq4kMkMtFYUJkuP6hBuWJIntGwvqR99x4zwVpObiK5nxftzgNrjuCeR6d
RnCUZnT9IjKVw1+fVaiTeKf80STyoIaTTrSzMXCb4h54ozpkS0c1ix/3+YSj
ZVJMRlzDWEOuhQ1k81IPGLS/sKWXjyshNZDXo76EqQNAhajsCyUkEITrHzcz
LW9qTocBTAZQSGp+g762kRl8V1b+Awbqj0y8lzxicdPS9xIe3XZdy3576gdA
FUh4oQmNakb+8oG+WoCa5jUX9jGSoexcwSrk06h+YpUiiXVkvAHzFgNulz/Y
cQ1T9ZRe3B7tG3PLZjMQjLSJa59CQhXuvB/ekHjOYuZmLg7+TexVl1hHeJJw
6Lxtld1zIMHFrFn0AxFWqscs2QBltI+3qe+oZvyCjyT88EJW0K5yCWMbwcE4
4P2zUSa+/fKSCj8PXNL8QTvtEsVNlNzr+OgIel0OsYKvt2+nEJBjjuvCIDhl
3gZ6m5KnuGLBPmITKh+KILYlmgq6WTZyGsC4oitfcDfV7vBHnJ8xTst3NflN
aHonQMDYO9Pq0XOO+QAcbFoaK99JhqC0XUnhJzjskrI1WMYE8a0cr7fwlf+o
XrSfJzSmJV+wfIlGmWJKxQlTucaVCy1Eyf9MJfMWCsD+A+KxrFLpIaFaI6bj
6eor5jhJoMgoV1n1CL7Gz+Hvlns6A77cmdrO0WKNIQb4MBQxlqYRva70ifCC
e3RLif74qdvKSfPC2WDn7NAzTa9RyvGG6JIVbF9qy4XN5mi0HvgLqp2U6hGp
S+EXkv3HU6xG+Bh0fiiZz7xmxTbSpLsVWQJTfDkmYlnWqfVD/vnvu0O0W+PN
tp44r130LivhYMjG+WEtQaTmRYwwae9r4jyz3WSHZiy+4HRZHoj4hbIIcB16
XCVumtQEnhqM+QVfoxN7pt5wI5sqb0Y5GuiLbzeYRozHtodOvG+LvKHh6JWe
1hDutO80wbnCHNSp4YvsAow6hqqsVjztl1zMnyFqfUzKephiBIL09tXVI6v+
OHSbTwIzM5Lc9gY8CoFZ+EREc64bUp52zi1Dp4uYNCS/IFm5pjKZK88yPQbD
HOrEykEI8JjkF+JH+atSvAukIJs6gvCE2fi8UbbzXf3gzaEox+JwZG4vaz7v
mIcJuex/XFDGfcUzgl074ofTUfCpQ0hcEkrXeEAqzsiJIBZ+U8QUAB0IEiSv
oHMQsuDaHkQZLEDE4TDVyYwDR5oPVOPKIiyZOMKs/BiZFRObxOwaaRPKyBNl
WK6+uYANg6gGo3wxWuyjXj8tFL2OxP7fjUW8EH823i7ucp5PCEpxQT4T9/8n
yM4p8cPev7CIcRWKSaj8og+1SnQNY/82Gdt42VPly02Gf3VBh4+0QSzEOwyB
eld85xrlqYxKqwNOxwZCs7lPoJcDO8V2aX/TkoDW4nzj1kqQuB3lBtlHKVnI
hum2AeUH8zalv+S52pxX9Q81NoEFNuaTWzoMHQ2op8je6rzwRS02mLH/bPzD
287ZhDGzfAgBcpj83rvaJqmF2DQ8kXDwcdDNapH53LGpWxxGbU1dWYXr0k1F
RDlu3/hf6WGP2x/glnhjeyx97DIGkT+UvoZ6eyAqianOd3HDqfU8vfJhLAda
qPNhmIyfARHKvfBvhDQ348enKkMtoaxw1WWXeTcXc4gpixlJSRoCUcJ0WA+R
+ecTmMi+EbGpWr7J1j39QLJRUxovMR1tVHfWSLGqGkZGNl8wHUhXbIaAotYm
XNp0wQtXrfcd1eA3Wy0QYnQyGlx8r2xu9MQXYYhggbtb85eZDLS+JYplCx79
A40ZV8JT2J2S9wgLAIvfM0YIMy0tR8rHx5plp2QlHPQrU38vyvJaZ9/GvDLl
tq3d3wNVhAbpfc0MWh8lJCLUVW8gxU+xZ5tsQl9aU5xTRS1IzHAlOLIfkISY
/PfUd6MAmaLeSgsDl9yXrrMK4mET/g7X7EZAmClhFNXCjmXas6RSTLpvSrpG
zTDdjdfbn5McF5GtxnAgFfzm7MAn24gt9hR3JicQ1qWH+M3PTvvLVwoCQkf7
1MY0EVhiSsiKHqPP8BF7BwA0H4SJ5/77EIl0wy+ZxcY62fTzpvCWo4u4DHPg
qXzJOEDkepRAIr2aRLA8G3z/vAeu0dJfadH8TTcXzhJAsmSkyivn5ZdfIVZD
obBb+d+/t+QK1deFrPSXUyL73mF8wE5tXav9Whd97hKRZ1UlNpb98Mgb0UTH
hw+JexeAtSLll0+PHah1xvqJtRNm07K9vgP9QCPp0H+tU8TM7/ImTi5HxcqP
Sisp+AUCz3mb/NA7yHMwXK/V7KaRW0ZVk1hFOFKt19oGNQC9sMWgfH70ECG7
XxDo5puKRFT2Z7b9RcyCQBztJ4uBQQhmiQZ5G8p3nO8FRHmHghmcIWdGraOp
AjyKc2kO2X9pkkTXddGriO4tzgnIEFpHxnbYgB2xjgp/flJ1RVICgwCAUduF
8nw+Vc672N/o/vvLtS48dBmTWmNIsd3L/wi9cQSuFNLSQuJBfCD/LXbl3GP6
/m2Cg7+f4PziFjXyc+iydxRwd5nWK7X3yQWKJ8B1QmPp/cFc+MG1dwW3NMA6
UJ4f2lI+0d4qP9bWaq8/6HhLXwLn3jt+EvhDsQarPAZyUccnodPGzQ9vbzxw
Dih5kuu3DZr+3xOr9YAz4AdnNfdw6KgMsHgyrIUf1dbRpTXROJ8/euqM664l
CF1bDe6Du1IVur37vFTl36Pw+624AQfuPF/fWjANwLuRI22oGFaoEP+SMEFK
HTiB854aJY63Qc9X225vp7ehTAPLo6SJAXTnAHKxM1GptO3vp29FxhfKCEFf
lRgkH726GYwduGseWHCkj19+QoGJdxdgim9li07RiytJqEjG4bI9uwzmVcH9
RUeolzoobekgSkTFDbNbX6j5asl+px4o5us1feBqunS5AlvKv+HK27IVxYSK
sW2LwkP0Q6KwvQhiDVR9Q9zo4qEELmDeCbNjV6fvMirQaxSzZkHbcCWzAXWf
/yCAabCZ0PQqK1l42HgyMDUkWrL/cG/bsoFl7CqRqpyv942lkNry/oqvdzCH
qV/Z/eXmBE8nNoZ8GxEos2JyWFqiOf0WjHPQD3xFtTPDfrC8gOHVFMqlbPqU
HPvLgkBQFBwb3135EdR0Ixa+3FrXFoC/8afNrgeAmkoJrP03/ckwwB9ZuH+B
ga4+BjwUNGEqpniAnJU0LfI+8SkSHh/PUzLK6kKUdEtPTNCceLP82xuTMfxf
FA7+2IafKuMbayt7DU4Z44EXG3Emm5rKlj+88/yOA4mi0dzsWmQ4fJdUkAan
uggvCILXVA1YBedAjQBycAdnorr3cjZ0Zdx3+p8jTtpOWLexxjGzDqR1S+zM
xnHUuHffoyzWW1cnaMjtP0RZHzWJBtiilYjxTrgZcTPrr9EcXy14E1fBG4Ic
ok/MWQAubtC2vV8mfhdjbl6kneJ6haFzrj35AO60eK/oJh3gGSpgGitnwwxP
iUHvhDCiQ/a9MbSfJUNeMHHeny6urAiZr0Us+7Y27Pa7eyDXMCQIq8BDfY+M
hBoBq0bEoqeBIpj/5l7gYoFoz3yEj8uLj31eYIm6AnedGSFl6jhAPDcFqh2o
YbqJUlNxu40oJxvDjDNv+m41xyoXHUdh6MBSuhcCW8W5BucpD0+Kg0lXxqly
yTQjlRKa22PV/ikHVgsoiKRuPZ+tl3wg+a6Ktr01A8pPZTGuwmuYewvhUfK6
jcb6DiA3pfAPQoh8nl16w3q8Yh9A79W1DTLnBZBhjfwzMVVU096u19sofMLC
/IBHYE7HNuFcP18r62FtqT52tARZoPVB+gmqRJqctmzvX8NkLa9ozqIw/RT5
8MkybcHX+SmiS1rhgJq2jZL0v9VAaaEp2k3d60PDrF8te1uV38wiMXsMR+5F
CudGXt1co91XamAYb49CBNPHipK97ssnEE+LCrjcaj7foYl30yMG00yhefUk
xyZ1FVxeXzkELHtpegdCu3F7ocEYArL3awSN5j203UsTqEUn8EQ4wB5YQVE4
UaDel8NpRKBZ594CMlB9q8peFu1AlnQTe+9n49rYNv0e47Txd/WV+Y5rjybe
TSZ6KP+XLfJr/WnqhWMkvVxoQtxNidmCL0i9dTbWlhzl7RDiEe5ScRkCGls5
K0b1Qjc8rfWyU/pLlZnL7a9OvVQUk0rV16Mz27iTKljPdfHVy2xo8MV1BwxE
gpzVl+dosmSJv8l/PURmH+ZTCeaplot5kjjY8oGabDFqUdhIgDe0dvOP8BBc
myVqJDkEhUnpzAnkTu7hgceLjjCxA6K/+yLGc8SzC0/xd1y5RyZIQbsT5Bye
jMo20YGCoxnR/witCAdYvGlhwOpp/QFoUamSGm8f7S+lniwevgAP/LMPWi1q
aoxrA4KWnTITsbHmInTTcW73DvUSwkQ+7wW4uOeyDBZHyp9tdLKLGfDx55gN
9CduFw0stkhhQJ01MYyhoRxmLgD+NCuN1ctpAQKQ7a4/+DmLEabiz4CKShS6
d9hVtzZ8eDp6zl8Bk3J92SCLqfq7ltxnOOe9PNhNoJONtCe4PGC7+xAI3UHS
Rvk4X8AJLefyJXpOmkRreQAuqiDIbuQ1M/6TSae1KW+IVO8h/hUmxntn2/mF
RC8o2D3a+iZ4yF8omfoeoZt6gG0J5rmCRwGd/usJvD++oafXPQ3hUZ8gPlJx
oM2aHpfwAtze24bA1UIhLieSbTYtsTi/ja/yt6AoWARO0R0fvLB8kHCMSxTl
GcRVpEj/CdM5fAUjLAA2DQ5ZjBjbnGNB5mtJlBdglXZES8B7VmARVrzp9yNa
IEZEZiXVKGrdma8DgGWDin9+B5WawyutP3lXIa3Ikm9x0GnrKcLSNTyTlBGB
b5LwuYm8WfF1KSHI0Ygskd9d295Dzqgsgxgg4qJTUD7VyOrfaEBT8jIIC37x
a6+OBtRefxcc53kFMSthMLTIdH7+BI0qTwERgnWh7j0dGrCoIdyqUswff6hI
Rc8GYIeJiMroGhNMrmV8tOuxxTtyZAjJPbRQ+fE1JtfFej/X8mgpoX3EIrQJ
8NE35Rv6UTRSSk+4/C+u+CdcICivivsWK8q2kB+haX5ljgLZdXVfnqoBzXjf
TK/qa6QIqIJiPiP7ItTZwRcqobHKxFSXqd8EauS7fBbpeL6UAcYQCM+5ivrC
HW4UoIRRlwFdTjpRzfsZk9Wz50u1QkChcCNfQJ07gRnzm26ka97AUIAa6rSF
gNz8j6kfXSk/Tg6Dg0qww3C9CQZwFi8sp7JJ1LqQAJQxU3JzwiOsg36QIDk2
WT5RX8AYbg0P2rSnjcvbi1+3Y6Xz8fd1oCKhMcm15mn9v0m6dwpgLxtIthaB
vNsV29kY1OffAI94G5N+QcAckWFgWJTk4BGtKS8mHebNn2Wos/mD3B69OxJ/
JeMKQBVmTbJr0N2ouQPreErjWLshvMGY/XWEsvc3LNjVthkd7MxcNpHBG11m
w/MmHzSOp8UWZa0XEsVc66Eo4z0lCqQaWJsGasgknGdT8Pk7vCOgzTvVl7+6
wOK4fWhfcoCnaJkSWhkkaC8NRjGxUpVYYTX/mdXCHDHsyqCP2Q0GYpeqm0st
8y8lAGIOtpQqAMG+89Qa6bIz/cI8gI+lU0m73fKU5XTVeizgHjVWXykhDTiQ
2rBhBUDAG5YrOOqCS1ijljBY9uUK56KQccMzHxUKc/dvfUjEd3WvQqo2Jmtb
+mDTIkCtZuxFKRPA1LQgHZX2ieFTHdpP+YG01zQrD+srT7deO+BVWLDEEzZL
3SZXiBXbDqNcyJnJlB1fPngWIFrugj21fdnWiuK91KMbAPaHEPM7af40cFhh
nCckqrozSgvFFkZUIK7aeiS7z+hLbHr1+nt4s7S8t/j5+cCdlvjqULyM/SY2
n5IsDlyKtnxhUF+kC/lyxzlnz7CsgISlYCRMYGizAd8f9eFjq4JJwy9rVFSk
bvFEgeFzo3wLxQPziouXPVJsWKLdd9q5unNPQWW7bJ0L8gbtcY6YhhBwi16r
+cVYOhC5xrIVjF9oq9UmV9NrBP4XYZ+3dtkItxh6tpVcBMi9b2VbZX3q4wMS
YPQQp6E/ClbKMc2QlTHZBQDf6fludI9AsUVpi4+DtBbhhddzaMd5z0H6Xkjw
i0welqLAGq6yOgqLzrQv1WpU9LRehBJdtAcDIfe3HVLyG9NKSVkAOTDxcFfV
X+aCvb1aJoma6qDgMlVhFmf8jmyo/v+nKUWhc3M1Lb6UvYcLhLXZXpLzE7hL
DOiZo1YSbC87dc7x11YzKfyW/AqTLQRHNuZiVf7YGdMexXHKnpNihoE94TLm
7IL4m9TM+vCPWHs2JWtXwq9YpKm5uqP97XdI4ZjVc94Ioy0saIiA3SNDWRWg
JycQ6AYEt3bV+BQ1D59nXMIFK0s3oykQFRtRUIYfCe/oatwyxpu/hpU/YKJL
Tg8F9D9YTAf/v0GDDpT2Hz4Xj1X3Ifin42UGgOOB1ggrv26FMxsW1qCYKets
Qh99ZhKpeZ9uEZTRphQC5fHtuHUIT8Ypzj8P2if3pYy31MUlCo0Uql3gV5Qu
bI9Uq8taV7EvGW0/eYVyscd4tDZ9gfsS9IsninfKecli8ILtpmRKsv0+Mwa3
nhDCqR6XhWEC3YE4TM4qexYz7yyHj0xtVQgGqXj0schY9QSYoVc0HTBAYmxv
iqXBpSxooVjSbMad/dUAL6DLyMVBWS7Q5xrpdhxYqDMtmNVs1FiNDUGb1NT9
6bIrMx6ztI/xHOShtxfmgaeJ+cvKkSdpt6eNVWPDILHKb8tkQpPE7XUWX9vR
AbKgFuBHfYA1EXffGsr4+rMT0VpzaSPFEJo0FzousLEaOQoMLeReWigl/zZU
oQ8gg1AQK4ukPN1uDN+e0xUzoeZR+KWyj5Z/D9LtpRVXsZFVbiZSw4eeBjYh
ekO7JOneLPmRvTa3z/K+p5kVEXvjHZaP4Tb1Z+2ue8+GD3ZaEOL06IsSCoDN
A3bVal1RjxjNut7wnK2OpRMLoP/J5NpOfmcOdQoxlu3D3vU4+4iSx2e2sUuj
udId49zDRhVzY+wu3bOwf8XSrPab7NjhWRsdGKxcsgQLeJa6WXiICez0XQSe
R0X44WmSQ3O1/Wb9H4Fgas0PgTGFOC5xl1zQI5Rt690xMdekbHUSBQaWsAuV
oprnbR3sFqWjRlx2Rh41JX09V59SNqekyk1R88fSasjpvMcc6jyPOrR3YvDN
5KltONqElMNLmguQZhPsSgWl5H0Bs3Vgs3JjExT1B2vCHGwEuJkU3LwJP9F2
1CwXAeE1wu3srEy9l+1mfCl+yHPIKoVaj6v0BFhG9jkPdToXBHZ2Yi7QLSOQ
Nj8a/nTAcA6bADISsumGxCp/YGA0CjNU/vskIybVi3bJvDTmdIqU1hd0X/90
Xr/2NiCnLSLJq5G/linHfIgdAC3ia7OsRZX1XNq6HfMFd79Gwe6leQTyHJNy
90p9/zHDkUX4R7EoSpQtjfuROTmwk8uhHWmy8PrYXvWfdwQYfxeZHtciBnJ1
y5sCXCf2nZip8eQtNvhduHU0CC/lfEBf3U+bd7w78Ij04jXrxv/taGxl/0ko
pIiRDX6uUryfyYBFAmIJ+bzNIgd4gFCSPvM44XO5gSmpysmyqCNyiBCdTxjH
YdagfrfwgSsozzqXe7zHrcqkI/PlmzQzXzxCYd1xFngqV7AsqWRkn2RudAvk
bWS31AlxtLFiIV6eSWIiR8WR3X9EcM7a1SRLO54Snzpisu9heCfRuOmPCKrJ
4X6QSXPENrORDj47wLv1gfGeVC7pWKKTKQoVdruHkxR0SjUVOFIEiJq1luts
GHJvp/CDU1iQHuqDzpYq5SysVWUPzxbKrcTGQyOvsCYlMhAaAYylDeDhMBj4
bvma21HOWMEweiPMhaq//Cp5uj6M2CIB2jcVNSazE9Pe/erWB8HQuzcFT95p
tJYTb2wUwGJBUatTe+68VP/7qCXvNmEGcQSNZ/5oL1r4o9mBcAwR9SZBMBPe
gqpRWaAOZmlPoEKFEJERb/sFAqVP4lgyOReZdJ7jq/g/8nC7tWnn4lQs7mSg
uHUv2QazDrSMiC93Z4Z5HQu021a6ar7cPWIXLNnHQBu5mHO5yogkmDVxPMjj
R0DERsEoFU/8XHJbs4PnT1Zl7sfJinZlCpCQ5hSRc4j8+VTztD4grjYdGRG3
txa6cYrdSoWDlqXmqBl90b2NWmb6pPhZdy+iUS27OqvYxpF1rJ/DLUsVdXLc
kGCJVSNmSEUCJyx+LpRDk7kPmcxL2kJ97+X1uLHNaCdIeXc2ysRfwIZILI7b
BzJ8zUhvZdh+Ps2S+a8/ZM7d8DxlbFEnvRERUgsZlpazRtfUVHGAoWrG/zin
+72FmDyI9pFtvNUJ2wdLczDle94vwvpxe8mtLQkHUcbNgXL3jZr62i6S9HQW
OuSJASvmcL6Wfj8Uc1dVmoF1zDWNCm0shBwZyRygw6zHgIq5fCia3B83OcON
io9L8QqSDspZSEui+Zj0XxPzgkhDCMbNAykhBnoyTEITNK7QD1dt/qKlG8m+
qMR52VwfiDzCW4fAPezUESDfkfsYDIRD13qEvsyr/AF/2z/tCaq2+V/VD56I
ClAu6YwKL7KWQtooPP0GGAGctCX8yx+ffbc+DQDytqxetPnhXh+FvbakZj/S
YU+SU06NPZAqUpqplCNWeWeY7XFcgIsoOlvAh2pDA6/acg7qK5zy8fzH7xSk
ybR5T51M2LauklHa8iwgb18lmupnPoJs0CQOVnUQpzuvXvWWRlgunNwyTK+X
6wTjSjFWAnuqKcRdpGbZPuIlQ3rAKA0Qdsx4BVbhiRYrJnc0p7VCYDcAcZ03
Pqh2JAcWm4Rz/RW0k+zIzAIZ3Kv3wPfzhztbGmMqFfbHaESPRcQeaSY3w6zl
Wju2hMiC0AEsssLBTa5+XYQZBPOgKZV4zKovfaZTrFtTOITn6zjPUlOYRPET
6/aJvO/m3zEB/G69s1u/fyW2Me9dp67p+Uv3cevjvghd3si5zeUIFKcTLV0G
+HkxPfKVS14fxexwzWlnNdxj85yDMtlTQatndefnryzrL6Goou1alekidqM2
5T6GvrzNIzCBcTDI/9qGynb40iuOFJdTIOhnjrVONTp2mDTtpWAidrNkMVmz
qVNyBJa0wOw/vRCuX+sYaR5WZeXTrYebF9XGz0JCdDrVoj4wwu28iluu5lU5
eg2Dwehgzku9lui1z0ZBJMT1tyMxE09ZJa8JamSsxrzHjo5gXyQNhvs0/hKt
44pHGszRlq3xdCDNzgj61V8suBYd596APNoqefFi28RfsBHQ6K9uzRcJ691c
QCsJFpbHKMlDb1k8EXa6RqVCQGe32UjG17U47o7vm0Tu/hmPqV/KOouiQmxS
v2PZjF7zP5MeiKTXK1YIIY/9zzz+Lc5V2EDZoZDmh9QhiKLaEBvZCnT4LAHO
h0U2kD7ikJK43pbqnyW6bNB6qJjzJP6SaEP6iD2oB056m3Nl6NdVU5INZAOY
56VPLD5Z4hO4w3NCC/RCLwbpFinbJHHjQtStisFKCV3iOgGr77vVSCe6QLKb
GaQfIx/8bvxjIWEvyCoSYuganp//5f3PJ5d+gThaca4kP0KBResp11NHFicH
C4ulvvtgWMz2IteuJZBf66o2HWGegshggLhT88JCHuyXIY1sfEHfx8lyBJPd
i1nixw7Zf2KvUl87k6dF6Uma3ZQUSgwvqGVWnTsl6rwatfDRUyo14+O4OoZ0
Dm887NDu+PUqWS4YDVEwJL95gFJPsXOly9+cmUBrXgEqKeoZZdduAct13idM
tXrQU/mAldsdZ2P0fMG6Xhnpu7WNHzHJxT+WKQOs86HwPprWbGPFVzmpuDVr
HpZMvdgcC9vQM3Yy94DDqb8uTsHmyA3+n15YA8sgEm4HfSELDwLYu3ewDJfv
wi1K5QxNFjiQh/pYEFC6IgwiIauTqRALRdI8LfOZ6L263eNJMty7e0b+amff
8pUAsX2umBh8Tj7Msawkwosd+suxJBNuWJeh9GcrRLxZH8ILU5bMDxsgACi2
6HUnHb+MnPWrvzEuO59cUBaH1XUvVgZgRbVpssRKFPw/SuFOVaYVdFdZVyyJ
86wf/9cMXMWDL7bKdmHo/s66NuTyFevoLqQf0p8xLX1O3k9Pz49acNSb50zq
BmXj2tmelLtB8WHnqeGe1w7PuYtJGShInillfK9p1nEYbASmzi34xksMHHrD
hWpd2MMcAi5nW2sni+Vyf5nQKydm+ScSsBUkx4ZnldRPeaSHjPXGVooCQNMw
JDr4qjvgqrXYmSYDUUY4uz0rIXOfGuyJ22rMcxCMVUBkWq8Ab+/2z+t244zf
ao9J8YHCuN6af6H2mEhDdYiaNoR4JRagBTV9sp4FSEHAxeNAqdDyTrlWTw9R
1c+pp1qU7mzaAFUw9hT2kkSKwPQbXUsMZYMPLEIkc62DWvHZ/BIq+/vGczOl
wPkNK2DkP69NJopvdXEMkUoDMRkgN4kGL37NaIqupTeOdk+gwOBmQvh0VrBl
ySZzUGuir6DEplbVT+/brUv8l649WAIoxPAgG060IVUKrZS5ZXd2oVtfjFSH
TzODBQmL5BiPmqq9O69jaokUXuvibHuvr3pJa4Jy3IfUD5a40iwwIFZnuPUi
un0M7H8YCKC1pGZ/dwZZ4fSeEuZLY2JA0de2hJ0LLXH6YFeRw5SLTASCU821
QH3QjHzwuVyBb8snjgMgdMtmOfWAtVDhlQHV3Tht5RaGUlFDFQyNLFECmLr2
K0iE3gDrTCqaMTHlI4+QxODt0WvBwTm6VYoCt6A7JGo+iUMJN/snInMnUHMd
sNPRj7St4daTsiL5eeW0/OEILNTcNUz7+cEj6h0Wo6z2XaSK6fbPpfcCXoy0
EAcZjIhldAA7+SI8wGdCi1pgP9JkE5ukgdaXMDHCpFFjzAxbQqobM3SPiLab
m44PHKIfcemJ/xrIEVmdY1BPTAEJcsKzU00hRbhNVyOoXtyNijNdznCmGbgO
ECm4nteNyZYJrcqgXe9i0mDMgnzo/PJO+p1rWYJyiJSEDTTsnOPfcN11fyF3
F5wFSKlIg1ZAW45J02y74SsbLGKqYht9UNSTZ8EhpT/KNJH/mABSgRu/Sv3X
yz2goh7Fb7o9S9lWmJF045ky03GQiqMMMcj2/F+O8SV1LMo4Jbhs5FYG2OGP
PSTi7HCyOVIaPHic+bp44IBhC1e1LBQNbQPhnTDaGyxLbu2lyc/UC/5OI2UD
BUvS1fxifYwqalAV5ppJuOzHpB4uICeE+Up2lFUo+4q7OiAmN4gyqS6+6n/c
qhOwU33IVjaqpW1tHaFkA6EBg8po5/SKymKx/Hb6MvcuoRX+mg0DQvpCRvX6
ohENV/Dsd7+65bsoAel7goZ+9xjVUe5IVKLftQ4FYynkS8t5vP1ZqfMQarmX
qBV2DNXKq4LsGEGEWEKANIL1uoA5FJi2/noBcq0p1gOojrX4ATE/QN35JNOx
/yH1t0mbJSTQ3YqAgKFe89pQzQBqNcxYIBXfy5eIq9YjDi69I6TWNuuopFZ4
LgwnHW15+6wNK35KwH/7vXjoDg/EasXoAFfcAP5dSy12xc7uAvhmIJ+TsPQb
CpeDo8XeGwMEMUsMfL3nr0rQvz0sNTlsf95Yqokdw6XBtpLQj4sIQZdXABh1
46iON4e17ya6Mv7EAklu3hjm80TL9MAJ2+Cnas3ZRkMDHnWyQv5E7ghNUVB/
8smWLc58/AjU5XuJh8N7ZqYMbwUZ8H3EB1eXd4/viHCGmFS3VePN9u0w2JR3
b+HMXqgeFvyW+TwLGTHFxsfNYIf73QM4E3LSaM+213JyrrYGQyphAMvN/jnS
Apb61cuFdLIQm8c+rYDIHmK5aZHS/1twHIZlbsItjxx+bq1m7XsdUkkd4qg1
UMZnmjNp+AxOrD1SGBu/68YEWsMPwlVfpJ2r4hNuwKfi1/BTGdeSODLaqluj
CG6BMmtbB8WbWgajQEAOUqJ/QANN8//+7RnOjE7bQCVuArYKug4nIR9AiHr8
d1ll9un592iVG5s4S9O0Wjvmgf+of41/URJIVcNtYCjoAh14FTFwXWwpRn/C
7y58pfPZYZ6YHnxUdRu66xDd3nc07XRGwcZuFTwf3kDZffjbJTtWeiXaayT5
yK1TNcQL/G7bLUKAItYfOC3zhsa3AtrkJ4dY2fRPVpnTRLSIB92DPDongrKr
/OagTN/PSTyYrNMFNBUCLe/CUtugfY4DUphwVPhmDydRoXSose2gH0ro0ywD
oGp9tZE7D6jY5DnEadxYNv3M5R5XooenLjzvADzLt4RlJdrxh0AHxv9fIMWW
368SgXvjFEwzsA7ic7updxLIfoPukrOreXd7RrFRVVn6I7CFBkn/R+SJhhin
phYCbTUCgwjXVqS26WevNmLwNJIi9awh7bW2lCSjinu7hG6Oo7XldtO1rM4c
NSeTBnq1c9DOvjG+5uN+e7mjLU3+Nkf0UXBKqyFjXyz8vEIhbZa2/Rl5fgWc
imuCcCfHGJlLgM+NeDp1gaww9ohA+NJj6jJYnOOf4ZrhvSPxw6k4dh+LWCtN
iTJ9XalWu8irGqX1UBzDtmL2ylsYqKczOqeryx8/Uipz/A7u5EROBYSzfdml
53vzNNxGILf5Rc3kCOHjMa2B/wx3kW5cHhx+eMVx40Mga+W0jMfwUfUktZyj
JK/UJJcMEkZkTYGXB6IXEAlJvw2qsMBHm98DSvLWTy4KXCMdlmA/5qd7SsKf
oTv1bFyCTPEIbFMm+r5ddwbwlVs8/df9e4H3trqzDbIIFFHDkbFx7FNr+/Rc
Ky0Ub7ZXTamxQ7WpasLMdXwBO8wXWkuj5pjA4zIHLoTvQw5m4I2wK43+SjSb
L00iqcY/KjBrp83Eibz9myzEG8g/3Y+nNMeCXWuLHiMqnXhnTvRgKvUzca8R
YyjULuW2mVoqr8ea0Z0qMQ7U3y020FySAkSs5CCNGMuW9j9ldWreJqExxGv9
00b385DQVDSzCfLjuiQQ53Wq2qFbW0oiLhZXzXSaY1FnY/NWGYgugx4DpNqB
dC6jBs2JEVG1K4uRN4ZwivZ9lMES7cKvIUj46GWWYN915zz9m+nZPGFo62fA
ImPrzP7iR/aEJjvAQuIr4+QECrDw6eXbN0LUJYY23LDxVdM0Q9jn97EFvh2A
kJPmguU0+HJiMQ1nmzjyPdcRY50DbA3btO5e9ktki/AqsUl8eQeEo2lwVh1p
ox+pUEBLjU+0GwDAbu8HahNpH/Ff8x2gP103bACuQZbAIFzJrOqGO6qBIT7x
PtVt0Mam5Ps6tGmjYiQR6mzOsUVK2cyLtlwRL3a8VH1eysXSgVkXRZTBDQuZ
rgsehxx5szdH5iqQs3LRR3yPMX4F6PvOByX4UUgLyuyJnClUcCWcMJgPPLAL
mrTagyuWJqZfdjjh571nljqYQOl7aXvt+dnQJNa/Cy3YkKKZNkv5kPTvnllK
eJwtD1EVLTjH3tddEG+pGtxAVhO5HxCOeCFPZm17A2bTMJoWlwtPQ7tHTxi4
wyPslK72gbrrKFMarJrMkyZ6leoAH/rI3HZqjksCx5ip4v5gN7KaNF4t4RbJ
peapZdkB33QT+suEbXejxH6Rwp4DyuL2UFoIebNfhI6NRLq8/3b9LJin/HqK
o1FxHEXrEss1pqnCriRGMAZVYox9mX6mA+jawZwAZsIvuccUpjdemSxghHfv
TfdKLFobnN7/EjcEKQFWx3ZPZHzj4a0ALy0yHKV/5U/P6SEJFbOqLDIm9lHS
u4XtpOWeCuwB8ApVLV7tWM3J6pqqCAH0y0YwsNKIcGUgGHt/8AorHSw32MjL
VYTyDArwrVxmVwEsoBnCpgKBrP1wRT2FDXKtKOzLD0ESyR9dxVqSopqk2fb7
PRfMrQ1/QLYy8NbplwgYoeQRW8n+FXF8aqWLbVQzmyeSOFObuPkmplgO8HyB
2AunhFUSq0rbjOkn0tqNA/qYTg73PmsJmNFwh0SNiiMxeKzG591uy6mQlWu5
vT5Rr4qUm18kBI7P/cr6NoXUpM3d2jwInAWWMJvbiX9ay1nnIzg5qZuzsBoR
vyZ+wbvB502fdCVjukPDD5kOMGCSVbryHJHmF/5r1kIuhZYM1fVRH9bqlhNL
GRmn5Jl74JnDvCLsMPobiIisVkBKcQhsbyU8KK+aWU0meCtPb+KF3C55YUlx
/uN0106TCdxwuF/3NRbdclSNI3ihKyY9hJMdH/eMQUZ8/L7U3wxTyjJknksi
n5UF6W+yvfl4rRR9PeB1usKQONWvh26J4wGIHq2dshSf+huCOLq0ADY4/mX+
pshtNIiHusXdCd9tifEYA56URFfVyY5kuMm35f4H8kQSKeG5DjTy6FhGx72K
GsXEp8b4oOYG8HwULm7YCFwxoNLHymLVuR+1XEs0ns2lGHVPp+G+Djb/phSl
DJyR1C3fgYG9s/KvrDhQNQLPUkEisjatAC/pAW56BuLIUcdEgYwtTqnWFQ+i
M3gB+g6n0ldsK13yb8wHXZiwknu2deOyOhtdSSYHjRUVpojzkRT/eKpKpnfb
YPoJVVhmt5YAE+KB1YUAsMYGAMoDeoet5B0LYM/KnuC2AZvHewOwG6s1rRf7
veCk5RzoAsCqMzddoG1ZeVZ6lpmQS1X6ILhjhQtYqOAT0sPharSoj1unljxi
Tj9t2Ei+RIa1pFP0qhJIoo+n82N90BCc0rnzOekFMuXxF04CrJWJP2CjV/0j
fX1OgNFzpfdbzWBJgLjdzlm0qDTcicv6FYE+bRLgE2h+7CRDO1lSPXGbzNF0
tM289+Jv18y8OUtwuQz8IyHaqo7sY5pYJNr5wmC8HidRsiLRPYpL6hFatUGZ
m6a/6l/PV283FK+eKpQkreRlRWBPCjD55U+uFVY1IzyKvGQJT6Q1F1Vm8jTm
EYLpv7z2sIXQXeHHXkWeOC+Ce+A1iw73qb74EIvBYdbSOOZAg5owTdQ3GZ8z
glrcCc7ldr/xTKupTPV3w94+4QH01p6fde8PcdWswGInjNVXncoRt3QheYNF
zDyztwkTBgv99HbzHDJHhmARGTj3ewC3QJWuxb+39UVfPxBer/UKJd/qei53
h/rPLAWLQ8uDWKuQcSGAnlIZEnxSgjc9WIRgNelekIJ2zBKdOFzmtusxsHKc
FATNn5TBrE8Ha6noAi2w0eK0lg1CokbVUy30UZdygfXo85P450Ey1SzRfxVX
TTdovH+WS9IrmUKk03hHNhWJC6zjxK6YeE/jJg4d91cN0hYr/5RQat88hPWB
XpQw2JAFwWeuyq9gj0Y/MQrvatsP8ktnCqIl6+PLVJvgkpYzYy0IKtzwOlG4
WfcnrCqWtQX1Exw0YdqJ7c2KP/+AVGriWItc7Sd6wIPZ3YFepnlHirqCuNVg
bIsnO7K3eDybpQSTujhca7gZhOD0td+VYJR9qQgx8P+LaQo/83XZW6C4qSSZ
IwmKgjMxISiO2eXHlc6yAC7GKKxku9XYQC3oxuJ8MdaZfjClBhCFyhflIWNZ
1G2zVbR2S/R1FA6dCJ9UjuNR+6Petl1M+8deOhr8DQtpCzXx4e1aecKp7Mr0
hGAeamyxdn53X69x83GlkM1I5H9sD5OKsGHokeKiEZRSAIIXbWg8AbY0g8u9
GtPUJ0qJ+NzIsXyboMycPHIB0WgUFPNF/9pzeMdJvjhNo3JlIV+QZ21WEYWl
Tx4UGAL7GjhydWG45w6vu8b6rQewpeUIyl3jaZbwiaMj0ZT4tIbbDjmJkbl/
K24+xfdm25zr0yD8O1iHCWBh6MyBooA41RcK8PuWPJUMCQoYoOTE4lToRRyx
KSBlYZD81vpUx/9yb8RvQ3EbxhBunKBTSOZlwThIn4rE1iFfOYMSc+30icza
ScKy8sXu/Rmkk2Q15KaR6x97kSRK7eWp6ZvnEFr3MbJQZON6WrNhyLyQpm1u
1i/U0DWiMiL5/pQXKDyFSykU3zPq2EALLWQGieNtnBeP1b3l8fjLNtTNpVKn
2+CqG2V5gs2qK/6/V7zuVNwu6TM40OA/jL7vMVqJepl1dundp+FVa+cEjGkx
qeo0fkgBkfcAJmkuQV/r17asZkpyyvERYZjxZasgeeZFpir7fhlNvp3klInU
VhiQJww5RtmprpW1iKdGsE5MQfde04iaOtEIeIYG0Q9MLRlri9pDE7J6iphs
IMk5aQR7Aq8ZaSCzYBT3ZCekMdaCgOOH9bAhrhJHOFzrF/3nelWlL+rCe+lY
581ID1zTpWoNYbXFKidrrcPAbHwkPzR4gvZvAdeBfrOhUvzREmeHUdfa6fza
Z7HhqcAvlZVqeuNd0NbVuD/2WMRvKTFBndBp0I5RZlICqO7bXWARdnxAzs1x
zEMkpqyrAB+xbWIRomUvsoleUL3N2r79aEUM8cUV1ooXP9Ck+zvSbiigr9VS
+Db5SgORh4Oug+XmQNmcKue6ZgV5vObor9UtS3GQOFHCQW96GXkA8QLQpvy1
/Ed1aWCjPNiyTdT68K2YmlBzmmWolmQ3K4ndqodiZI8ocrvzMfpniOSUgnEh
C+GnnmLoFqKLb5A4ET16bAbQ3HDU2ICJSxwSVl2blly6wiALbF9TyKtn3RSR
ZOmwnsJewTLuxj0fWGSP4cruq3y/ZrRHl3t0TWxHV2Xosx9xZJzYIjB3XebR
pmm+pRJO1hFZXe3Dx0XaaMMoDfLqNXjK1O+Z5+sXzx6dZV5oW44dqaHAleeN
g8AWyCxua1hZU9msTOUom35Jfnl+eFzxLYPHRYtI8B82ts83jTllcrqHj2vD
k/elSQ33O5OBKwB7NQZI52YFhs5/cLTm+iUmrwF5Zpp5W4iGA9pqSS4kzcCM
9I9A1PooIugGGrDGzsOT9ByUivHeIVz+2Ciwb9CiW03pM5L84wYEVt0EoI5D
kAcF4dVzqXmdxIK3kj4XZIo4a6glfs9FjiL4L6KnLqWYMBAK58scbmxh1At1
aCJ3a2XhH0T9i8DVihC6Hz2V3Rdoul6q4U/Iwn7Gv3hEj4MbXZj22DwMixUg
qxxrYDh7pDBfNKCRAZKV0htqifVsb6mLJp9hpGFKxRBbHv3fWCvKOCpHMac/
QrOe2bqtLPUCaS3OL1UpC/QCSaAfxCGw0c+UU+5UkcF/ByQJohW0gtsvGOdJ
raD6V3qZmYy+StC3+cAoa+pqBtg89Zw30icywCdi403wIN006jHr5HLJ6BKA
uVPe8BPVUWyjNw2/UQXc8Eu7rS8FCfArn6YU6ku/G5JxayodrrhMHaJV94Gu
SQc/Mc8PorJ5Vtl2VlpK3mq1tbBgTkV4X+axDrZm29zRHXiwr4DKTszntwjE
4MIqHCdL0JlT4f3nnxYiWhhfZPb1d0tNNSHQTf+Lmu9ycaV7Jvg3ReU/TOm9
4hM2wmVbYAuUAhAxFSodRb+FMWg1GEKRhl8XnBnJtfTPTOqoF7MlLWEZfw5m
CFINRz9NNy7gU+UNY+ZjW33t4IkkfkO76bYeirwbMkqYvaVWtAMY6/eEgIG7
gSJc8oX1G012s+63cdq8grBTxRr8IJEk3MG//zrJXb7BHvhPy7T/GbSExps1
mQH/ftwkqQyyWuZMLnAldm+5tFHVxUONxhxgCwxQm5HhhKQSWhF9k2VYWXX6
2aa4lqh3asyIrL+Hzl5LgNdYptQM5edh5rnep/sTXL2TByveOMjZVCnO7mX5
51GkIPvpyxJ+UiscYMkPGfi53FfKVea2ziFqWG6L1+vsWIg9Hm9dD/56Ed+d
IbNRnUA7+egJTJSS3pNC/Ji0xaUSy1BnJjd3UI/NwgHDSXP6zSPhXm9NFSYf
6NsVxqKyJLyYmsnJH4qTkin7Gn1s2qxLH5Wdeve9URsQfk3leQ6AcWe7hdC8
2R454gZYLqK/fa8bA/KcWtpIfCmnJO1wwjAhRmQW/jDyULSkP2FZ/WCYqRlA
Cm6QDqBYKJLufk7EF9P26W3C7vp3jg7uEA2p1tlna5WHXg8aZa0rrLdCbiFr
pVQCwwfBjFSzirgsF5FUnWmUoPMRtDFtOFJl5qp+yFJuXEMGAYJUUYqyPaja
PNpwlG1CkfHJ9tQg5JaS8QwbUixPDVPC03S+Jin2MQpuVBQ9EVHuFELF0khs
vA732+nMNgZWspT4E62FFIqymCZyVwzMW8LU91FtT1JCSpl7EmifqJLIkzat
LVWv04FtXP4M9u2ri/a3nURSjEds8kwSvz7+HA8tvgghZJn+WparjXFailvq
ewBUuS/pZyeMhEQw+1iR5id/4H8jqLPZTbuHFhnDD5TjLXvNErLm4Yz00dFM
ymkedZdE985Ut7MlZtuhm2/nyOiBo408Zvp1rt2xTgxUYrH3hAohCNGa/Fmp
Ryf6OFMPaNS2oFRYQ/TZ7N9ttQ7dJenIkB1wA/aUPit/L9Q67hq63+8NFMd2
QPM92TcZy30HdvxtZkBZVJlwL+IYMi5PKk9lQuQAVJ4DE3lBc5z+PL+fb+Je
tQPR3PPF0BJjem2wp1oG7eEhWSU/Tok/Nghp9eI0bs+tKEb0ebBF/0ve0PkJ
7Val7d9Pw4v3UbfBxy4fMs+Q0UCjmEVqOUgW5vEoNXwRiCwsh7zfE3kUqsqk
lFwu5Rk17q05ys6qSooZuXw23fMOmty5MAt4ZpGo893CGBJwnd+TvCy/Azyu
BdjltKqY/5Q3Zf+M8ODPtMBcklOLOeBiqg8cjji680tEi+lZG5H/yzrmUIpx
YiKK8usjW2+xo6DAEZmBowAInZFYBwK7pqTaaZRpZgWykyFXSqbHFtJkImnz
1NLZMlNLzUGcFU6NJWL4O1PDGTXpMOAMkbtJmv5X3YhaQMqwn4BOawqF8F2u
U7MvvWnOciabIlYmHlGdyC6GA737tntY22RFOUkui9lqkO70B1ZW7O7dGq4C
GMwVVrT7a5FIoFhrxSMN3Sdxs4GlciwN3WNGe4yciwTA0E2x06qymyKK3c7n
5NwVyLU95rTM0e4yKv1Y81AGOQ9FdJjk5RdQntJDs5kszzP3y+nGDusgqHpM
xrHYGxpVslDvpHmSRBCHgfq3x1sUd+pT4VJqUgOjGEadKQ0I0oTVZoAyE3XC
mzYmqt9loai013AlXBeEyiANg6y4vZiPzkRHms2sUsb4IBPWrdDZJ3WKvaid
9NfG3Awe3FLW2gsrspdZim8jopIXv+mpVQQTn9Qqxkm5cDacxS2CWk8E4v8K
RrEuU6nTNVWhWJ8yjC2O1Ig4f6R1gA32lv9EOThoyyH1AcZPeLAwuGVnk3sg
je7LpDSL+Hdz4zbMMhsZDhO951rKx1VZnW+X3zh+/im+VTU2XbjxZ+OM7Hxh
c8b+DyoB4pfiWofCgQIN4T4TNBd/mU07xkAucCd4lvDCd/qh9OMMvf+n2r6u
JQB99Lx/sQRnomQBq2vvEaly7tfceI+BJuqZ4XPfYZ4/sZBImCgpajRAwsTI
7xdBOMd2ZfJpwda4E40geYifX7+273HgpOYJgraUk71runZUf5rlasQNfxBJ
FNgZReC30oDiYy/obSrJwsUCTEBWPXnImlAV9jkn0y+NSqadtKDAzu2fdvHA
YNIuR0v+1LbZjb08H7lWaaa2a3eWr70eOGXm/DfOKLU+U4W+GvMDv3lFLzF0
9x+/+6GVMe/n+eaMXs4PJs6IlMKMyp4rcVLla/OXuN3eYz49YfTuEnSO0Tvg
24e8XKy8D29Hl/V7iD66xA310ZUK7AO0RDsgpFTq70GHoVbptuZFRSOTiTHQ
ozkZgbFZINMJGEeqD9i+9t2V1QlHI/2GgpnxNid11BVj0s9JkeekJRLoqRxY
6XOGXfJdt+u/REF4e9Heqcs+j/JN2q2y0Xv5nhs36W6OqEW+WMuMrS/WNhsx
BmfvRRj1jbTCmyMxtYWOyCyZ75FiHFjiK1xG+P81Kr4o6Udzxx2ynYvjM7T5
5Cj8u/HRKT2hOqPardeQ1JHve7Ccawe95n/HhIF2KHJaD72WXKUqTvNpdSGf
tcw8AC+98FGc8Z6Ot9eJeoz1LL1UoWPr56nKMTLjmzRzzHCXxfF4NPQfaSzq
FP76jPTuG5UBTGcDgfcAj02M88wUw75dk4AVEI9FyPWXqeNPhi/Ey2BcEQAN
NENPGjYdN5PpZaGDJA3vHUoudPpq+BAmhX6lIExE4yvvaoMtez6uAN6egmKw
UylcVU6lDzL0FPwHDYEFnFFIe8m8i8sBvXAuBuuA/o+QdwdVlEDXpgR5Ebq/
cfy/yTDBcRs8S0hvj4pXGFYINvoTwr/TmYel0VXeIQa3sR2lXeo/vQtwYKqH
hNxYITqmkW7xsH7IB95qxGEEEI6kxBly6EWsHwYeOdAQ2APDdSvQwstUz/MK
tu4f7VuU3TskfWfH8awRHQr+VBo8aDQ6OtVU90XQ6mmQ3CFbLg7ysvUox8fi
UeFU0gZU+epgxhpdpH2/YCN/E9Xvz+DkG8qkcXPeelBukw+Xf5siVp/LeJbj
s147PtZ25Bs+riuZRJ3vZX6FZ5Ncan1gKKv15Fd4WM0gNE+9WV0JerV4wxSq
mNdf+UlWii1UildSg47hnDQN1Kb4HhaXOWQ3zCtyj9rQbALZ+9BiRQsvI6IJ
+JVWjJUoYGNrCiokbTg4QzfaBS15YzsAlMb1Ekgq0lEHuMvCw+NIFZWiUYzF
2ztjAfyzMcCAKat5fM/p/UG5Asdq7kk+ZSkOLIDqqmojRgj4fLQOmroidbk+
+dnNgYkB+Xmn19OEHaAKaG1OgXFPzEdoof7L/YE3HVeDwvOFvBTj44gHZqO9
24cH2/3vaWrUWN9DJqL2zhq7/JqHdPGaJZ60NwN4LPk9f0eEVlCrCT4vYRSL
zA86aaSZgunxYpMI/xW3at+oRgNA33S6qtQb65srnZFYxPLfxFb4TJsldujP
k3KILeLXoQJudBkNrULNScZ2zvOsMrp+2tg4kq9dV0tkeuliaswfvK/vTwUn
P8aY0Ke+4geIJjzmr+0M3LA25FxA9N9hUqEfStT3Z+wKNCneabGQH+lWdnKG
sVFHYSsbd4vxJxVFL0OdA0VLzN6fYx/6bRVk627s7qqVqaYK92gcxGB9OuyO
Q4bvH6t4mNWO929mkYBufEtU1DrjYHLPIE2Vi42wRhppcipBxu52xNADgW4g
AC9espMhl80VJpv6AS7/nIbHEkqPw/BZFqBfx31Noig6WoUm26KEhDXskalP
0pH/f7eiCuu8eToH4rA4cmU+V77klrpEO0cUwDuPtYBk5dwpM8a1LE9JLCUy
0bfZzdv5PbHrImmB8tOa4P8cfW8UVCxc8DURwbd7NypkzJt3UGBoqAT8UVZU
uEtMdusOQiCiEgWvbWgCbNsJH0opPyIEJzYCwQQOC2lb896FacVbU9Ll7F+U
XmXCTK0brHat8o1RSU2j+/Wffjd9MtP70zo2bnKEq+Yf5dxVokQHLGeUFzBd
l0dje0FwftZlh/wc7l8DFLgVRP0TRmdCrlMdDnYIkNRqJwtqm9XCfiMfPCFQ
Z8jgo0P/SV9PJdkWKOsQX1Zd0zP9wuozr79GBUSNxzSTL2uNdXI5BmzLXwDY
oHopBhcb4Pg0bn/arzBo+45dCeEgMnijMXlc26YtqWtKZ2srUE122XR9pDbd
8dRIfx/mZ0tbmdJI6LAcMRAH6qV7CRatX5QbWdGBTb1JLOsVEiojvqRKdfzy
Ia4xDnX1bNBMgdhXWlM0DYUMOeuc3Ei+4sm/CG3lH7krvP+2jcENpgfmOjVj
YZP12X4WSXheAornCIkweXXW85vVef83vizYbmiNXXO09BSXAkRqwmrz3iKf
0C7ZFQFeuJf6+/6S4oPc5V0ujrB26CdigHfuifX7c0RL50v+sjBkOiqMM+Yi
wkO2GAfN+GEAPrRYyhxC3Owkgk/06dL9A9hO97KGP8HqokBzTlKYe/kWloi+
80hYt3i9QrbVPqHv2Bb3F88XyOBA3BtAOmeEJeM6zm+C2Mr4GfiFstKqSXis
1XzfiQgh9GFGsd6CBtck7Ms38Cku+QxwN0AyrTeX6jkwBmTcYLjBBOJmWsTA
grSRXmnLTdSDn4qL43ObFa33olVVG4bCgJd4TSg4jjOEtv0u4peKlMCwTMOC
0fqE/qicvkHadGjgi/LZUfMYxJ2HOevW/GeOYWZgyZe4b1yWzChXmNX7ajwq
3tD+0Hi70cjm9ykLLBgdkoYPwLB9na0xXLumoiHHTHnhwfJpGwdDowN0rufn
zQYuUzS/kzlGaRa1OHy4dYbpMsojLE2gFnB89RXKUEcvZBwk7eUqSaXNRtND
FTG45aYAN6+FDKGgr4J8Ge10TmSVSAnKOokeTBwjzQr5CaAMKroz5ACw81z0
Hzupy+VIX7ev0yVs1qgc/p0nGWva+cQ2bpN6iMSB2Hhm0N0OS9TSUuYnjsiF
B9JWDHOcBlL/M1X6+ndKSooQ4wYCHuok+ik/3Y8/WX2wV6cYBmlLuz0Jj1Bx
ehAWc4ov2+QBWGy6ysitqo1x/vX5ZT/s9yhGcxwkXCkFjS/QkW8o5G1cZT8Y
IzNVCAX8rSYvO8JdyUSHu6qPuZPteh6+B5myOk5t5MeSNuSafe8tspfhkhDR
wv9oW4ia+3O48B7awHZi9+Ihe+ZdBfJRqsPcOYtJ2HwmpOn+N1d0Qf0rA43M
I9hD/Oga8TeznPD1gGyuLHRMpF9AtJ42q4BGKc1qzqMo95GH8y+NGo63nSXC
Aw6nEfTkU4cjmv+XigJBUrDW9HngKXKuc0WyLgn3uN+ccXTkvXV/Bg7IULoD
E2oblGqAsvK9X/Vee6G6F1PtrGM1KdyY88kM57q/qzgE7aXAQxVFdUCow9hZ
9eBENn3ek63vnEeTR/tIZfF/ghlXRRh4NySfnjYdyq53zE1xxSctfTFqeB91
ZgDs8/ZjWsi3ZW+vFbjfWB38MDIUUkeosu3StSe2Dhlz8m9ZDlnoLdBrQq9Q
5oK0lWQZkDLjBP5NPk32FSxQWFrZPaNNKqu58/t/BbKKY8g/vr2y8n/zOwmP
ntKM8NecucW2/pk8r7AQBO0XdlIR9Xy7Jo+WjAAQvaozELV8nnMXtff8phLx
FMbRP4wCcn+K7Ld4k20jph/mGv1QJ43iO0daVSckVUIqXzL7fK32ZclX7Ylk
+W0jLB7099YsjWniS0ymfcrvpBR5Zv8eC+lPh2HM+c5O4ZE/QzKqr0GRcveD
ND2+FCLl/njsCLjcBZPFfPyCt4MaObBdIb7iG+VpX7bQ/XMxCbc/wQBGfYO6
W3prAtzqaSqq/MwxYa7HcMx+O8HCAPT+LBG91bhOeU92t/Q9Tqm79e0M7owV
rfyvnfR05KxjsYioqNesadAIP2JBp5DbK3XxyXZNNm9QkNgJvmZQ6JLXgaG6
c2fjnRcBfJbuqc6ZEuPAu4cEhUEI5NoPHP1rED52BLw5v9p9MjLUHvog07sU
OJaXSnlPFskO+Nsxwb75pfUf8XfZRtmWvv4Mcxz2eqem4Q0Cxtb4f+1XHULm
ZqxHIBudOUhyHkOOHOngUC8Pjz9nGYf8t9bT0Xp+7SVCzt/csZwUQtlLLFYu
cHqQmLYtavZtXERYm4yXY9wYdi308ehjel7vcMCHEx0nGWLmkxY/HMDAiO7w
FKiDqkItCBV3lnb3um7xN4Fo6kkL/lofvwcb5zOUXxwsL1DVbbtpk0dx4RHS
MUXeIDrUtSw2AIQLT3fY62F1LwCyDWQjrB36rZJusM2cawT0tBxQlq/GL5xM
Lt8E4rjzO5y0CaA04+ayrB7JOUwRDZwp56Rh2CSRMwnRAl+eXp+ClscV40tC
5Q61S9XcdYzoeMHb09oz/0+ABUsFS1TeKLlFb5e3/0Cl+FjNbuhVl81L8qLX
GYRKt1g/jscRkjojL+Le7IcedYI/61arBKS1NVGmDTQ4T9CY5Al80I8S+n4J
3eahdolfOdywgg8KjhE0k6r9zlKK1qY1jWWfmq0YiWea1lhdHCTpF+nky/Vi
tsIk68Fkru0XO+8lehHDX9H+JQ7Bwxbql21GZ0hc/7ON4txbAvyvsr3YSDny
cIeFhgU+Q1h+8nQ06Q1BqTpUt4WuK6vQxgFlsiPYlCD1A9Cfl7Z0Y4ahk37b
9ttKWRLBtIB28yTZS96LKTwd8qM8jZ/2cXiDI32eMAVq05F2fBCJ6zOfjseg
7RJSRiHlTHuuPTjYJdmXRVCtfeSAf1Y4rBao+sOJWe04sZh424tXnt/ap+p4
6y4kcx+lWhcnDJHQwp0d5VsMohVY2EHx+EHZMv72spzsDowniXHz5wqqUng6
6BXvxcQcGg2NCHbS9DPfCwxDc23pIUXp0JQqqVS69riSVZ92P6kK+W+HMZrB
ZYh8AYkEHuTVybODSFK3srsYmEW86fmItt2UAzurkXue37xM7bUPMnI5C6TN
HDOtMQQK3uYU9AjXxF15uWZCTSpgkhBLwzjhKTDwxmCe0QVKflta8KPmVZft
6CXKXvaRQMXdF3sLKF93tOJTmprUqKCv6Ytjmavz59SLkVQS+4hFEzxDXWf3
7vC0QKelOOyL1eZqeMNmdV1w6IlZe7UoQATSzIhBojMkKXfTIzZZQ+3I/bBT
ZLzK42m/UtrhS1MDlgHDEvgHcv2oDJ2pbMyQL9BAaIFcNJdPC5JUa0asywth
jqFqvx2FG3UGdD70Kmkoj5c3EVtg/xStVXVW12QXF0x6Xm9OLqwd1bkcxuEX
gk7TvBKFG0VeP8DhYcwB4A/ag6k4ExtteblQq2w0Lj00iue8Rl0/qQH0dNtK
e8FQ2jq6a/90th5Ar+ZVq8/87gAreSytxReTJL0V7QIvFmvix9hWGfL51DY7
mc1/AEHlZgREt0cNCiJX/E31qtEqQACL6tWls38b+F4zfmuGhdAfM91kJ0kp
bLsOTRzuGdfs+bEnJn8GsDVEm6l1Lcd58QsjaAFlGELnS1gBP26oj0QPbIv2
VlqFLZLcE2r9b7gACvLXwAC+RkwO97EbrdZa5iaETlEHG8FRbAyrqJbYsCdj
9LfaUyOy6RYitOa/kLruuNu/noG6Fi7sUjAgn2D6blx/XYLhvuOvbCwsA7b2
xhIsSYhY0/wCALZRC+5MXpzOYd/NjDUXedvWZ5yY77QvUOSqkfZNfr2wt3/E
rwgMhbYvJHLINtIaA4BhGAEgPNsF9gl/RJMWDAIzT2ZsiQCimzGPonb/w4NC
MUZZDYj2D7hNZTL001ZvOZVk1B3NHT0mhT3iKy9Nf4ZL+sXrjudPDCQw5abc
iQooszgbX7JkRlb1WoDo5k1ouKKksdBUr9BklvnXOsRHoFK4Jm8E3//pzuNo
jcwqx8r/m9Rc2J5ZWb0TDgViXyqZlco7xXaPf4DxeAlUSR2yOB/vkeAIimKM
oruYm2rRVEAMASB7R0coWZT2MHVNWyw7SBHOzWPys3Qq8zZANtvFXeqj2zU8
v0pf36hJ8/i8OpN0/XZAJeVHLBkSrfC5/JcKiqaHxRJ2XTJa4pZeEXUkOfqq
L9yO9rjsgOVoju8bDS/Nf+IhdsMZ8M/XZs4fiEvHvYG+oQcgFi6uuNlp8e8u
Elcvj+Pd3ztWFsyleN51kTBcky9ZtdhYS0OA+mguaslLmDymqwnqbfvuJGog
ktEAr7MGCiLsRebahMah+JUPndXqRRCuyrUDJBudnd7RI3uIeQGeUmJhZIRU
JHhdCCP8aZWEwJtVLr1eLxW5QjBG2yx5o9xVp5s1wVuCsmvKFJczKkVJ45Ub
Ge0bkA8RjCHzDFm83HPpC2xNEAYzKXr/aTYHM7nY7i/bhEfG40x7HsMZnoRR
JhZZhTvpA2cCz5ANoLQMJc7U/kBwrSFrUg3jwih4lT9VDLMW8F5Jiq0obOYR
GJxGLm44yEYE2XOe0ul9Zcq6KIBIAeovT+PupBHAkPjE6hDx2oW99rXGNgtr
z6jKMwEZXC7MwIkkPG4InvkKWBNWOg2Ua81Zob6hRhy/RIBwJINLMwY6hGO8
5bplgMJKhf7z8ndSWR8PtjK2HVC2gO1mmu1P+AspXuN+qwRGjpjCmYwgWVDr
GeJ0PLqYjZehCSh4+UFtG88W1VVCchjfporHurlwXgQ+WfMWnauXYfUahsf0
qpvvEc/3MC9ZTqrlFFFh5w/FRK3ePiI3YlrKAOlAzw7nt6olY7BGNympFnuE
SPjecU1vtYyCmpczsHFoFows4W6/yvDHfb0zud9ZQylhm7YB8DpiDjnDsrDG
RdAyl3xacoImwUYPgmjG0IOoBwKOSpTs51Ks2l0eXF8og1oGZXGwj7FS1KSM
aMF8lxvXdknSI4GWBkGWByX31rdrcQ7WEpUEwcWpsmKYPEWBYMhSVJVk//hD
x2JAo/cS8P5OIs9TfdFAbm3WGB3Sk2TodFR/mfFIgIer+yLyTXUtjCfFzlJh
diykP8oyQKSnL6r4rPj/IfKQsXqvggN4GypA+KN2aa0etZUuuzJWzdp92a9F
NVGfYXiIhJgThozNOQKC/hvHwto0sRlwSsPKAHwoCVeUP+lqbdNYA9+IbmlI
v1y8+XVePdoIohDiP4wYxSLxoHLGRA8lNkHjQR6nIQvuKSFLh9Rp49X2kEff
rV3p5M7QCGdWju1qRZO9L31PhaiCK5TVokaWOzohL+OzO4AgiyYDFiGiWqTR
fd+trihO/3IhkoGqVgf8Gjxv0Awq0I+5qQNrHopZRjXSvNz//J90x7dudtK0
DtuWpisvVMBQE7il2vijX6O+Omc+N1wz/WJScT959duRxu358D6GvVOS+gJS
w+ZyeTlYZbWSZncTLK7TdmwZbGJPkwJSGbnePzS/o2jfmp4S+TA+hW/5XJlf
/bgvbNtD8Z03rgEqaaFsvFme1cN9S4ysZz8hez81TyFa328zJGdZARkvHy4G
L8davEg2/rTKPeIUy0lGh3cxkSQCK1HlF49kP5h+JtGTMVZ3vAy2LQZoReMp
4Z0i0bz5TwxgAtau9UITkWcShSqH76G0sO9bq7PFcvW/cL9EAfFC1Du0/VQ8
e/RgH/bsv1l6jjjlsqrIgdlQPm7HWIva7KryL8SVZ+5h4ib8jjmZY4Z5t9UL
aUHJTzlGvo3TGKVsQWSl9w4EuL6cgj0KH/bU+ZzF6ovjPThfXRd5PuFrf+HM
W0/Gtxx2I/A54/Meq6uj9nkhLWcBeNIflveES2UIr/0bdlK2nkpUB86HP1aZ
UoNs1lqmxnS5fCBstkitvrJVn1D15JCSi6E40lqYYlsGuPIuN5JQhf8RRTGn
+Fs12Ko71EIH35p9521FyhtCWq+DHqvEyIXcGofmripuMpxIPp+JhJSBZuy2
EkUoyr/Pc6+IfHMPZtbpEZ8cwUWMaYuucc/4N5QiewU+l1zQ2cA/DGeVpIsi
X32QLw+6xhdMULy3z8vm94ARZ0EVxwZ9TWKHYiB0dTeUZSnGXY8dJ9iMmzBS
Sozmg6kdr0t7dzxcaZ/8Vz/W5aM0SJVtYihuA9OT6Z6yg+QJ2lJ7xyyyEmRT
q2yAxivzZMYTPoTucBRTS5Q7nzDuZAlAoYDQsP7Xr7Or46mrA+Nh5cIioAOW
FpSjRFXHHt1mvgE9KFl5RqNJPerjFvaa5TdVJxGcrVPe5/gc1Ghj0kmGGze/
W1udEnWCEr/3rDeS3rNG8Y5W2cVCWU8/HNa4taFiCPlEvpHE3tD/Dtmt8ej4
haYmA3JXE8iYYTWvXT9oHJAzY1zLHL1pGAeeSU6jGU9wL9mz3HMAVgsjZYKP
V3NFDjAxZGyxZ9tSRzaC5I61Dv2i3o8iwBsU3JW2prk1y9tKVHZsjrzNneHj
D2kzm+IrCdEQSy+4hJGdo22HesrY0E5CIQOQMbs12oLYbv9OcCwb1xBu6a2h
Sm2QHX7XooX9pHqac3I6pvqIjzTK30hI7M3o1LYb+hkQcJgBkhd7qoLnZ/Pq
vQ09Oz8b0S5/mxew7EqF7QMq3NUsV+sla+yOVg/fpZ4cYgOkQoT0zufmVex5
xExxs7i3H1FlaEiaxnrIPnTFeXBi3iALWdPpCPAPxVLjkOvbn50mRfcBqsYE
oBe7WhcFbIzCIz1gmE/XBuuBk9IsPeGuGF/Z9wNkasa/2c5lMYdaO7d85kBf
6czHNyZoREZlr4RsynNCAM7e0Ul2Ht/RL+XJTFUx/wc+puYGx9fJ7QPeM1V3
UQw9CHqTz2uKNCkqfFboBGNYwwWMWKc0+g1/XMwaVVHBugsdeFAqVVure21t
uQA6IT3RKuJh3VJBEvW+OrzbrIPP9l6Dg2HYC6GoLxda5DfogX3ywdI1Gws0
abz0Yv4FW7AJ80E7SXmZd4ODuSgFervI9hWm3vzgtQ4x6LilQF2Of9e9SBke
qKgBKCoGJfDdeZk3g3vxIP2r8Q7OUDGPRha/Ro5iFPIzjeVWHh1bQrJ8thzi
7aXQv+ChtQHWLsJnUjJuLtlUzEMKP1fCd2uGMI74ZvOjcyJw3SvILPJ0Qfx0
ASOP8+16ZDWtPnprXB7YUybe4OereBFj2f8W0J6AB/saqFQTTiNDGdY9sSWC
xuPbQ/Vh1AxaPIkpKhYzGk1+TvKEcXT41U5bGYzJkL/nJzdYzXeFh1X0Bi/X
2P1bBsn8JG58f2OmRZgMoS7bN58FBtM+actjI7zvOv21At+Pef7lYw1Tl4rA
WMV61uQwzswkp73oNd+0T9ebrukihDaxNa1HccamM4RIuSxKyzCj7wlZ3P/u
YfiBIhhCUop+DB7zOkNQZPNlxaNuZap9zK5+333Y8VsovZyAs6wDM+nioJvX
wLa45FwIs6zWfsMNDUSpAl5vANi8Fe2+ZVQcdqwsXzPpHuQVG3Srfuf0KCyP
9SWUedSWdPpAM9e/cy9vZz7/1FilgcSq2Lj3bNS4zPe4JChANjfoTTwEmgbV
Zi+Rk2W8uMtIJvZ9yRad7fWBQpTP5jALXStIG2YwFuMRBeRwBIg6GwpB0Neg
/WuhCpLMP8lWJwJmu5vadoNtJqv6GBK17H3u3YNwGoOoe8MAegqA8xiZkdEV
Sn4RjsnabYo0k88rpXhzGXRhzIRXSBTnz+VX8S2nuAcsn2jGLei1GWThtsB3
fQmJWWrtPhYGFdAGZCBau3c3VZ5/VyRisVL9XKJvUcCsPvbD9Lgs5nVHt7GK
JHDi5vKKMniLLo4FubklvWqeUcbuiSss7jT+wqnubH1O5c8U0/uHbsKYihPc
UEf+mOj+1qxREZIoHgn6zuOnVKC/O6DadvHIP2hHg0kUSLFR9YDIPNQ3AthK
7RZdbwtOjSWyMUXUci8VAdXJR0bNm5Jxvy+tKZ66GozoJg4JY+IbfVh8n6F0
e6yOCgO+NwGQqL4PliBpNSudYEA+K4uM46XIUxV+Jt5rinIomt6XC6JUD5u/
Vv0UK+/s2v2lezufybI7lrqTuXrKI6kXuBjosmSsu0I2DYVOW5xCdikFmOpd
q0Rw0HSrZSZDrD/JruHF6Ni1oZ0PcFa2FksVw0tud56btvXKEl8FMeFh2ELD
tQoD81+oRIUlJRRLYTcJYhTm7lnGvalA8e9quL5NHEVQejkhRnxAkG+jzCt/
kk4CsEXFazBIwtwn8FNUlux1zlEyKiuhxs4n5djqTZPNVPy0AaWRjOhT724v
o5qqUsactWD//0YWkVRJdp/ccggnIpucxWg7NUindf/O7YsSrBTMyddT0hca
G0f9/AmnWHhZLeh9tmQFlbLr+vt0uD/jX7oX1Z42c8ltnak8zUrTpewdLexE
Le7bNY8nZH7T2KVR1U2i5OmmwTOKvsxSnqgl19vxVdOCi9eMS3TuJWhh/M6n
5Q2k7Zf5r4oQ7vuG6+/pGS4xDpRi38Pu2Fwta9YeJa7x9oS/t8PIwSNmsr25
05WpkO87HiVnzLVKubRayiYbLwoYN/JhTV/pSpwf/U4U3oB72Bsnp1mwxjjo
tC0tNU+Q40m/P6fbpdI2E/Z5frIKAYu5OG5RGpzb3KRphovLgvVFBnZjByJK
ThnpeQ8cPa4SJVx2KYCb0IRmOGLYJEgMkIwV07SiW98E2cbJZHfGMjN6BMlz
3DdT5J8O0goLxl7+9FlPBXJ8yC+hdg1SNkDMQQdkyN8FHeRzJe/a6ayGK3OF
ghS78bwFeukmA5DHpeZr8/bHQDXPGNDMbwXBIy982/0ylylDgjPSS5pgGV54
3LF01PzfZlhVsaCfZNCQcILYKmjLfxE3D8uS+Lg72mR52Lc4l483khXh5x0O
sdeZbDa/Ai4qmxk0ejOc/pFAuA7E3pTh5FpC1wuiOjG39+lxWH9+XOWD4Og9
FCfqBL25iFDpFSrw4RjYg/sbyhkcnGWuQvNuMYo1gBUELp1OmJcnxq42Hfvx
JLHdWXGaSKm9bGHZMIgnohSptF0eLbrNGvOVN+OCA7qJl0+w5LBJNdfy0qHV
uEhbhjDcKaCSQPl+F6x0pefCzzC2Lec0mG17NmGO1PWQrjRJGPbGgic/LIBC
7ADm6FyFRrPYa1jUfFQXSRhU1pUzt9wKt0tY3YJ62jY3UVKqvDA+OjzTwhi9
YZWmGaMOjPnZQIKoBgx+YnwOJErubZ01sdNz6s3+4wV4oVCnzaMF/2i7X79r
nlMbsJanm1CfWGyFgbb9B3Xj88VMbed56EtqBz2Q9yj9GZaYHggEXfTU+wG2
OKfBLQQXA6JW84kv2mhsykiinBiCFzLAA8LYC9SEcBMSy6fgOdlZA4YC1RWN
rKxnHUFzUDVJKCdwzT4LPThzYIhfdwyFHjrkchmYEtaSdyX2h78cK0bkA5mR
F3th79GnPF2eotFYztcBjPcH+s+ynVd+YvmwVZO4t6eJn/cFbCz6dnpINcyH
lMN5inDKpr10O6eesF9rS7xAm1R0hoY5HSw5u0mBIt77Bbb1xMCWoSgfOz61
jrESy/vYsqQZQmDouXBmqDGoYW9L+CcCD2Poytkcuxgat+olMy/dy+szL3vg
LWkU7HzhZ9MBtBkGU8tkzurQ4Dcfhki7aJqImo7l4G6OsrJkhJJfm8lFhz4t
Lew3GdI1+9Usstwz32brdot2bJ8ZG9fPs6e6tUx1hJwqINKGFzSO47Cqu2zu
rNH/DQ8a7bCG91+BhF8wzTUGA1qlFfgDBlbQxAht23BQo4P78RtJyU7YoEn4
C94XgUdfEZdRbHlUyGIl03+2m2SCA+1X6Ho/ZJPZ+aJXxtcSWUdWaTuMHVVg
ImSpk9t3l84GNQqfl6KRcsaDch5MW5+OOFvFIpINVtNQ9aj0QFyxUZn56fqr
pnlOghCuY0Le7PFCX+Sk8Plgr288ShgXAggU2w6ga3BWxRSCb2142KGgKdVf
jD9J+TNrPEkB5ZQ9wwneEcsNINKZnVqrmu8J33PyWEmN9VIOLjQVlzRU09KQ
Azujkxff868yVyQR1I4xCeqnzx9GkA7TaKhafTgirogJ3FgPQUESt09iA137
6zqK418OpgdbvqZZRZWsqnXOBRDFU8niBx1wuEqgVLKU/QgrtzUNhZtLkqPL
ImUsxp0E0JbPS44symHTthlDryVQ0idq5u+hGE7jtg/QrTY+HS4zkvA0hxLu
bxCpv9i/nFaRsavJ0N63odsBfrJzCK/vLv4JoXvBssu3KoF63pwtLgClU0se
Ze07svzGvX1umyiBDc/4DSOIp9N3Ca/7L6RHGhvJHFQjhOO+ifnHJQl/rmxM
HRq1eay2Hwmky6bVu2Yl8+oiAShmrr8quY2dlu/oMB+5M0yv/99gJIOHH5ZN
Z5uIVCgEsnEhMDUZChLnTk/asY6b2cAfINn7TS3MhW8zfuaMNcqtChTn3pPK
0IFPpBeqAMjryZUamYJe7GNdy2TCmRtKjx1wJbS6Se8DiAvqcXP4c4Ja5Z0O
MrZRtWicGRDe0bKv4odfMG0Xls7t6XV0MbXIFvbCdWcpZ5ayukh6/nwVD6+f
TlzNzV67RP8RGhuj6VZB1pdcCNs3TPw86pSt6z/ylgzARq+OTXaTW/6Ipwnq
Jim1FUxcOzIVbgbn5i2GuHccJ9Bi9Gp3RurBhBRzfyJAPS3kIXXhsxE2EsSm
WtXLh/RnMrjSFxFYhl4MKN4gXAnB4zXBdUkPhN0D2gC31R6FhnfJGUjaMgh9
/g+J4KJrIBtY/TmIf7Ia/lhffMHNbAw56PnkBLjPOFJvqJe4Mj1E/87fIsGj
48qvNaxCVoKyknfsjKugkSL7rlHeGelqfki4LeQF8DNxVoGp1qSpX6UkfzvV
piBTMdi2ixBDT/Rm3NEBGdkpCoKWjs7m0jAAN9shRCRsHSq6wU9cRRj3CA9G
qhDykKxflz03rw4tX/mEhJi6VKqTk4dA5tXIMRm4Rk1Y2nRdDw0FuDSqyISP
kgZdWx0kOHoscLtzj5d3DeS0wBr6kSt6KCjte8x+H6eiDZJXEwZOb6Kn57Ks
N4PWFbcGWSQm2G81mu0TDahIKTCisEzVCjNPpGD+J5vKjtky5Yb3kSaGgh0W
lHw3k5dNuzyFLPQzIgBaAzdB37tU2f1V/OTLzmscfV7G0e4FWeqLT/pqpbK5
ZnItycU4mwgBUXy/v5m8idXqTpeB3uoyRkBkSg6uNds55E+nFrbvMzHV+D/P
/RR3O8GnYGWWpOVE79T/z9K/g1sLF6dYHVVnBbevrnEW0xwXhuKy3K+UBUCb
StYpGnC0t+RYLTurr9FQnRNEP6szmOgxV75brz7KfdlyRdkCcyA3vQyw+3b5
LtiyiSyiK5c9dKXfikUxNUj7ygp/PPqufYdz4mK5fY3iwV0l6BwyMcGCXyYs
VQpJxwkC53CIhCL5LQdqRmA0MGveTEiJI/TcIrGLeavxk3bxDwO0sp4sqxkL
Qh7H1tmsEq371/1Lr61LT41g41t+gSfFYACtj9/CU5bVJu7eO30HM+prOcKV
hFpWFXS9ubI1twkC70mmGShudhkJKta6YH3WV1sCVFuz9YDDosDd2mNPDiwf
YmowVmLks8SjJm8vhvmNKF/RzksebaCviJDuhorHNENINwwBAiXJTAlT4vVN
CRyTPSI3nLcEE5fWhA4t96mcj75+J8lmLDw/W3mhGrfddhOV29DTHwVUEqRj
u0ZC4KZsAern9i+C3PCq57LQcMXhhSHCXZCxYpPXg5p+XGClOvOQ9eB9IWQe
hkymsRNSbW3G88lwMSOHa3/mPa8uBuWRhecRsSiZonhYerpAkN4xVdAJOYeK
JXhhTljZUkosldY86ikJffIklFyFvueHw4aYiA86WsB4x6V6srsCBC+x/DyY
X71I1UBeJMLdy0kSaeWUrmJ4fczsGN1Jc6IaHaUULqwavuivq1nPt7GW4Ius
a7WHBFUC/L33sYl74lN5ZKA5QP8QnKP75PqS4x3LjayP0w5TLVjdgNuQ8PY+
FAcswYScRwlyQwvXwJvEjLCOzMY2YebwWYjaSEkPtZtredMFKHzKIB5A24PR
j/zZXQQGgJP9yd/SfDC0O3RYtHEQ+TQSo/iRA/sgPUuijIxjAi/DMe0fNd37
Wb444wVTtEfStQaNXO3ZMTIvdD/CuLFiBgTVGLR0YfRSG0ToUqfUjLJzJhIK
NdrtvHmwbMBm8dZtiVeYmy1sqrT5Gfv63SYAxGqurH24AFxhQLk4vrcxBPT5
QfS38WkSwvMLNJOLQ426OL6e/+MqxKyA8Zdh6QSsc7Lzxf05uur67jfQiDoc
WJcekXfr+HFLt2jZ0ocpQuulRsYclfaGPrIleXSrOVGYy/makfk+KYKZ2/4n
FQ7K9ewNzPRvujRWyWH+78YFCh82RNu8POnYW7YZi+t11VIGBbFxWC03p9vc
yROC5SZKivIDWOiPHSfy0V96K66FclFTjQjB3uE/QsDFhwnB3K+mGNyEQk+7
tvV1kktELmv/LXUf47BPZpKqiztGc+B7cLiRuAAYub5jBI7O1GR3KDs4e9cH
8ygfih+evc+oTdGze40lyDCy+9GKUc8WpEhXdrH3eIRz2puOU8AKxDkWHw/b
/RfrPkV0PrC1tEEwI9fB21oOyLlhNc3x9E0zE6JkBaAWOWJEmzoTz+3ovszk
eSjwo54umuHQ6qklOwaTjz5FBWxmUgdcferexuI31kg2cBZEbwzhqo5564EO
1NQ+97TPNQ9tNQI6qL/RqiK5h3O8lykloF2s5Kft4iNZHvsI0qWFeW0j/w0H
jxw4G0nXchGQBs26r/Tb7fiAwS+2E5oGHyVoF0QBlN9EGp55zRqX2Wx64Dsw
h/IgFfvD1sOfnQS2Q4HXHC4eo04gROMOtTxmY5tQfG3VdFxfeK/24YuHeIkt
x4OwzUNTvh+OuLgKdJ67dBfqOxxtx6MLAzBHn/Nlu5tpCrlx6SrYmY39jYnD
KVpTE6ai65fzu6p6VEaklfDHdMbY38D0rxnx3UPM80cdh8VnVbZW1MOn+LYC
sa2Ot7Gm8zkMhbUZ4fLoW6GTdBVZ0Zbmcj/N55yLvKE3PxYeqFV4o6GpZKlX
F7y9fKJq1kqEOF8eWWM+XQ3zG/HKy1uqCFx7oN36VsNRJMcNKWA1jnDBbKn7
kBm7ECBrFaCvAmCz24oq4HQa9WVHAzwCXa+MSOw1WwBZf+lmgMCACp4SRU6q
RjazIEE6XCRnVIVsJ3jMa0CLxzJosCZ99RR6kh+lJmVa8YaIQNwfjgvHQwh2
drCS08caN7sM0BPokfqzfCvBVQanMHvnjO6xMlEHUw1c6Gdpk/mptIyPPt9n
fh+l0NePx/D0wwTxBnQ/5IIhqOK7uU8v2XZoe+NHlmXG5j6kFZTD/qOLiClp
eRRWg18uqP+nc50OqT9VX3QO1HveXpyUD/G+VDGK41bfs8bLWV8bZmighfjS
Fdo24xi5zqSNyB46Up0Y8QmZLdYjQN8kmAKykY17w/U8Ouo2AmbukO80zn06
09egmY4aycGL9XsBECni//ebVfBeDPAJcf5GBq3Q1bPRb/mESoyDB5+GqG9q
GRF4/Y2Q1Psi8n/gYGEOKX4Le85PhDCxPgLccYV9HmnIajF/M4zSMRdGV/Ik
r/6skaenmntLLxJ2DJRb5jRyepVs/yyKzAkHgN6h/su67bRnGJNoyglH4vwc
Vbs6PlS5y5IRMJvzd8zuSr/rYxNIdVzcl2j/M9wzm10A7hsEId9QW7JcLQ2L
y9v7RAlH4JymeZaUQspNbcPwRTgwhh6JV8xRC7pGm2c5aKNaofRkWX0OqIa5
huBREcZxJ28XRj/sEDklM9IihMBO2MyfdZMygNvXQvxUzIt9fgxA2buHY9om
aaJSoRILgi71ddY2Oami8ZOMye9UTg+i37N3/VOa6Y+zXV26psXjhyoMAwTX
fkY03OXHDUrojnPVliFYbyqhxEXovxJBDtldl8TeGFi2PhyJpCNwFpNIYVhf
ImldtU5uhqPp8DmMXlxc2Iz/5HgfofpkdGwh+2dvfDFTWJ3z1rg6BWwj++7/
KPof4bwU2WOeK9fFq32/jUsoAomhadoLQ+sI7Yo767Mt/kizn4eHOr6URgXY
RzE8SaQbbOAsscXX93PUyX/hmqcFChv/UMU6u+u8frAKtDCa3k5Fc3ABooUn
0wiHuFvxzbQpDCnzpX9BP/gIH39r5ocsILkhu08d5x22CnXcu5vV+RGaRR3c
t+B4ZgGQZNRi9S68ALzvLrO6RSMtIBYPU6zXXak9QaEfoE++mQ1FCcqxdQW0
KiE7A7uVy4FN/Qtl/8Tu2C/Q1LuUFH6RVTPcKx8d8Og+nQyYXq5qpXvIt+rg
jnXzEcuMfnhapbJ3ZIQeRdjMiEfYtu+lUe7OQUtag/Z3CsK0bol0Xvohv1VH
Q2WgMyG4ttAwySXuOadZZ4GFNABTlmn3qgFKfinFTwN+wBWSVgBtDglY5dVS
knkN9DrQE0XamcviP/1uMltouJL9HryXMj4uOOfQ0ySRGh6SczHpXG0rRMHe
smk13DM/KCIgKTE0sNmSi+R1rXM8+kaOm0K1ZtGc7xamC5sEvAeHYmeUnQVo
GzcElKpqZQvnqppVX7jbDT+Ayb5zdQ715OEuR9EcR6Cxxhw3pL0+QI4Ak7QN
T/4VJ2okSmaxLmG8+/iIzFa6kome5zRju1YQaQd8KfKCKD7TDSTfXp3gXpiE
5WvG4v5chvRxkQV3g6oXvIPj2XMcHXo7vbWBmYu6FpxllxFt3UBoPi2tt2KW
d1oFMcc5n7dsw4NMmhJvbwSBM9yiK0KUAhCVKzv82Ljxxm1oawnfWkgCv1lE
KCLsiMQHSYLfczREj1soEIxjiSS4eMVOjdn3qmMgKq/3Fkhg0rzm6V+vU5KN
jlUeejvAk3s4s6WLWN390JiQVUCsEytGV8MiNH85Plym7KYNGbe3Cg/RF26O
UIIT4TSBRSjS5+iEsciHT2OPBvVoyWhsBKDVDltfde0fy/XO4Ydix9Ox9pQH
46Bvp8wUIlcjakT75p4lxb3GLWvMXOAPr78tNMePNdoo/sLI774MpGHpquzx
GUZg3JVTvHasqYFJRue6R8ZOFQ+NpzjLDvK09X50IATdFnVfTVd4MvWd7Is3
DbgBEknyRctMnOGIvDHh8umJgreyN/Xpedve5c6FeQqILOWYnkhFnndLVp+y
PYv/1wNMa+JZ//DGrkYQj15Vqp7aVuZulckz1Tu/XyaidM/cZH1AAGhi/wW3
MviV1fuvDVicybXTLLCX97KipHpsBy7V5/oRJWp/SDWafQqa1szdOnwDkz4w
6XyWXz1+xmtZsBzP6TOS5OiG9Q6O3maArvR2o9YGHN1VZyYd4hPYiPgCl4Vb
lF5WFF7FToKES7I1AMeTYlxI6MLb+dn0EQC1aKle+2CYI95a4Zp7rw2IrcAg
s+RggzrrEpFdSU5wvPz7ynz2dD1qiF8AofizZNXI0HmMZjPwxm3zj07ZPaRC
Ds4ixjx1ybL3/IbEK8VmtM7kg8KF5ER+Z2ZimFFBSnOSOvqdSM8tRbs/rpns
RE8MOGUjpclmaRm5hFUtRfXkziYUWLXZ++mgt8RGZ9pZ4T1De1Y+6W7O//Dk
idsVWhd93ogM+lVBc61eTy0mN72hzR97cGHJBbhdJN59UoKnvF/KIV0Z5eUn
gYXDP5IWnYfsmP4USCeW9Vn/H8KGzV9EnEfLxBuJ0m9/mg0oRLwEhpNbr8vh
/pkE/5PXFbqKQ/c8mmE31Q0suLbUm5V/zWpu54bC42dKuxU+QprFP2CA0Hke
OfGaRBagZMfwFaaf3qDwnTDWH6oH0B4wTzCLdVoMuoNIWQtVYS1KrweNtc2s
LyMctR+PIZ9StuRfIMQbRs3juEb0OYte8Qm8GLUetBuovYzCz6OwQJzyEDhv
f2ydckNlcjfcd51Br7IQOqAZGnCEcrfz8KAKf0WjmaRomnn+HH8J37GwJ3+k
HZfzK+CFJrTU9UK/Rwq7EgbHi8h0mZeczejN88HiyEBfirb2dv5djH38cRGJ
wYXpjarBhGnxOgPxfJWaVCgQ2LrlymPDAYODkYqyh3gSvizJfAZWbTeRZm8t
6piiHyTIyXFbAEeTlwEq4A0YWhPUu2IszHpaVVfPEkwW0SQ+q59gJVPQ6JXd
XOl8wsdUQ5dzXdx+SZ9c98h4zpjldVRi4kNL4t5tdZneAO9isgwvVXiapCYq
0nsJJ20TO3Aqty4LQsGk+9Ff3RXWhkxmkYgK7S3+CjqCY1QgN7BeP96qKH0F
dUc2C/EkPE18QV4mD6Fgm7Wpd7QR1BsEY4+6Mtdaw5m4PEuvyKEGrCOhXzaU
Y54xC/PCAhbGgT+67da5Ylj74uj7suXPbWUnkYjdrmJc/OYY5RzclcFH02Nb
XIgndtBsEykhbX3Ffb7lOztXj4HP3lxUWHwxFPTzUE8Nb/+w9euCvXNsYncC
MFEDCI5PlsOPLy9hIth5JThNepGisWzxC51+pvjRS8R+y/Sys0qiSJR5knk8
2XM9Je55Mpnxze4n4tulPKnnzIcVjJ9NUPZxHpsAvonXF375hADY7EvDbw75
7JiRkHy0meZyq1NbvzBdvExlEnmC9VMhEhkxyhbPvqpBkYUtgWbxaCn3ibv7
NM6KjNbw/Q8V4WHZRBLinchmvYcH8uUa3q0eAQCThOpm+7V81K0fMHgoh3i5
6iVImXs1FMClv+NmpqI9w6OaSQvW6wG3EoSNthbMQx/CPxyxd4j2hdkEqcIv
59xQ6XgvF7pHllpXGxYSXZW4nnz6SW2Jmlz/p3xcfcdWYCBwR/HDFuZXYcdz
CWEy+/VprTQb+aeZFzRtWV7dQJuVegMCq8FRLffO8KEBP5/4bJzIxvcdZ7So
PTtSJxY9h6URe8NNyJG5YIAwRHyG5AvDeOFs7BK0Sy/mFwQBLmAM5/jfU4iP
XUZnqsigJkQUj7ytSfLmUUEzec4NcnVLpprLEqXoCsItN0sg8msfig0XemPn
/p7GmVi1COHRiEPhuREIOcaJTdhCIBdZVuMW6jNIT27/eyAMwejXt7zeEmuX
bmhAJVWFYkS2NhZXiXjDN9ZszymA6fuj53nFPVrAfEMSLrWeNiUDQgTUWTQL
Emec75LCRjt8+XlrUQUBtFbZ88p7ASk2Ri5TSp/mPsLrkilUWVhK8BtTHGQt
+H91rL0v0+0ub89IEU90OFxJ6w0KGyWjjOgmmcnoV0cRxxGq1QFR+Sccj/30
tbY+ODraitrBISE78/14V5veH34TQl+JTcGZ/Mi7ytjTSPwfqevHHQGJH2RJ
5tCFjSvjSY3em7qVtHhjYe36yGwEI+RqYCcBDtQdCofwAGmaxf9z39yHBkyW
AEcYQPpo8YkYIQNQwnKF6+ZlkQkdOG5ICMJo8d14Cn6fUKOZYn2MROZduVgM
q3giPYjQCOZDF8xjfKxI8C5dGFpQOCKJrLgiMxu76RFTCpgH3KItuaQY+Jpc
OUCpyBxzM6zDOxi4097ly6qypbS1yBUga+9H+2x0000Q9Lzyh6AC5hkLt4sp
yyRWrDJmhxvCX9+s+XFG8MkNk2zHEZCiSjvu5yfjUPbLf/zvREtQ3nxnrrR0
+Xi5wAg6+qP7Bg77C8f5AFyPeYV+7FMS0NglP73csoPE8ljoFrZQAgmwTEMn
0FRiKLp9EYnSXY2+MkPwvfYt/KRh0BuyQXa8YfJdNqnUXLGUzkSQuTCFLCIH
KepSxHLqNDKarzzQvq4G00TsFJ0/ONrlD0hP4c93FoUbe+b3+riDDzJzYiL7
j3mTVLLK9q4ZA2do18YzYJ1wrm1tGiAg6+qqYbp69dfpie1CSd1n58l6A/lq
DtkKB+Xv066NI/aNcc6b2emZSUIyawY6uaUArblnauJ2Ze1Gf4mOC/WZCoWx
o19fZsbS9YMuja8uVcq+sY0ZgJ3j40ksjTEHvYgQE4aDflbeT3HjN/OaVQPh
emPHMPgnMUWL+JWYLoamJcDFU+vLdZKgm6KKIpnajeL1gpK1TBMoUvBN8Z/2
optJ+2MhNvKxZunOuhyLVlsLvI20RFCH/Ugu9YYMWeZZQ7WwgATNQXMAXEB6
Ttcn/bGyfhn+CiNPUMi4WW4vh0gTx9tpQbiqa+fx00Y1IYv+tKBXMmj8rzAp
eTXmTL9DwqjHQjWAe8Pmwu7+8ldNzNgmL//1zS//IakGY7c2UFeq4RgGNGl2
ChT9eTh3W+WskC4TSVnzqy0oFONQxgd+qYAR5PxT7XU9Wr1LvQDN8QCYYSb7
KKirB1vtFrf8LMNrdZtTVd+b3NCnBDt9BmTIs1sOtAbU0MpZ1f1puQ7SXooM
r+Y3TIghlM+fPGc4L8zq1F1lmKMNT7Ukxo1EBms2Bk4IMDQ6BLvHRcZwJZKZ
sMx2RJaySngws0HNIzZC27F80rDaZmxzDwBhxHRLc78loWRXaU30Tg9InAAt
pRYyWjDaIFHeZyOpHmkk6JwRkZeDKYGn6izmNP0TwU2TuRbchQZG0qUeNYvI
7TD+kpMbp35lrtDuHijU9aNIlgClIDJATaDW3KufciSt0dxoJq1TkhR1H1Kp
p7hIUBDxHGi5uamI9bn88upAuOsGnNypQLtaGkaAc6pNhrHv8sft8fxh+Ikd
grfOc7NjduhR9GqR2H3HcAuU5G5QRJ+W4OjFfBK+ALdNl2M5HQuBnyuLsaZR
lABWISaDTX7LKiYu/tjzSirkCDeoQ6m5hDWkrpDrC633uyeiVaRley9l0jOE
C1KL2luG8qs4h7OFlq7VEOv++V0kGN0DXh+esiUix1h52TEvytSqU/0FhIrR
Xy7DZho6DxFUMa4jJBzVp0PzmY9KmPF/RscFXxESx2kWV/6Y9l6uo5HeXfav
+LvWvd2hfVYLnxqSWC8e2PlDzyROmcDgAIC3GCivEa9H+iE+VzjTF7NPwiV9
fzeoXh83LwqJgvMXRmb5+9SXKr1Z2Bl44LbZJEK9ckdHAJzyZF1T/nNnSBAM
z3vQREG8B1r6CDffImzX8F7yNtuxUd6jqFuzFeRTapNwF1ls/TIRdSIFHtiG
Zeq+0zks2y6YvP/d5Of5tbXD8Tr68RLYhzoXN/ZhdZBxi0LNJI6PQV45Ygw8
lzUcNEmhhtrUUVkUkS8xLGLSP35VGN5qFL4Hq4XUySDm3v2p+3GzFCDxkZBe
EJU8613ImG3CRJVhaB4mCgWhfVqOC2aYqsH4XSp2J1XtMHkqcwgkUiP0gNBE
Qta2qED8815KZ/YkzYFgiVpykZGTBkRdKumsSpAfMrrCik6TULZCXI6YLDMD
83ENqrO/yY/u8oVj8RFBTGy4U6UdEZBjh5JxVVpniiN3YZf5z4dqb7u8gObJ
lyW0sorAkSODuqhi1nUtwtJjrfB24dDicevK1E+Qyk5rgGukOYzifptKNrG5
KpnkaL5a8d71JUS5cWgpl9dPBjRbFx0W1Tu2baGVE8vtj5c0gZ2HHuaaCryl
HlgijjRnqQhh92XNfSLvq4/aJJnQIlF2lug8NVbNLssm+jZnsSeqgJT9jYxE
zneDCst8E7DYdEAKTMHRTOBqVR+z6a2pChA8enFKu7RRtiIf9BH8g8GVjpvu
sX4U+7gY2DufJTrCAivjFRk7+2FJU+DbldK7s8N3WwQ0tRdzMfiTjGrwVJ9L
lZPFZ6cyLhg3qICL+FgpYp/4NXt1aWcPjRWf32Sg3oH9Mn2LmCL91s0vJkTQ
6RI9ZUTaO12yNQVcDR5TS+BZQqSuTJPjK9itjqwgET8qGm+Tj7hp85GJOVtz
0p+Enu/l65w+5Yq7Nf8QhPdOhiLcQ5ifUphyC07sEKdmtS1ssJf07QpfD3XK
28dQW21SvUmGd1aBKPUrnnDlvExW8dCqjjirNhhpwsphewxfjmaSHS7iWhR5
Q1PBy9PGQENuFIHsqPzvjs/dYXk8CRdvgqvW16XF+EFs6b5q1WJ6KJCChHp3
uXStH0U4uIHBXpfg5nuO+mMZBuUchUYZrNEYvVyTrmq7epqetmlJKqWT1KvF
CocNETwDlgRtNLayU6gLgbrCo/7jROmCiMZgw+9aNGzmwaFj0V/GsIIF74+I
8d3KSB3IqGtJx27qLAVXwSqjo0nEAGSTKaZBb8+G9Un8BY48TplAdksJ7nrc
SPK8Tn6OHFtGkT6PD7ZAAKMQDgT7TLB9oAzn0IGu3SIcLr/U18nsRprpvhvG
MRJu4pYfx6BxnTRG+MaSCZ0A0nvAb3ATm8Byjf6E5kE5VP0WlKcudt/zUTe3
v+/Pf/AC2Dk30HYmditEJWVrVYLzuoWX/CVlNhdWVoFQH3Mn2PUeGKqIWdMT
ft702i37NBzZn+3lqJxfdz+o4ObYmdzJeQfSjav2uGJqKi92luI9w3nD6Bul
cqnb2hFlSs4TMOMg88srxB34FiaPqDM7n45jrG16rjzYAgi+Oh2Je0drksAl
rt5HzUgQ2xiZ3atJsnu9EU6DvygmEPPfGuG7UTMCyErbh7ZIoVNN0I2SHv+s
ba3WnKVokGMvN8tRkO10dlImxC+fDKQBR3zH2DQC6kWgj+8s59lvIC4mRuaY
nQezkmYXYlSiMQ8K5EoU4RFG3mqOxYAr3sMPJezstwm6+6C1CEZ+6nVK7J4J
CBOxtARKeN/5aVRtxlvb186eQZjPJqRKCf+FsJvybwcn/66JthSCnwi5BORL
b9RZCHR1GK5tmV6IZS2B/c6aOsJSGH/fvmlLJHzdFLLzP3bqNFwUay8gTqBD
y01YOUj/WeByMoZtsMrvNBWO2F/ovdgESeAGQJffz7bpKISPTG7vIhf3/k6n
6MPkVK1pnjWB62381fyMBiCv/7Wwh8MhNEVhCSo1uM1AYkMx1Efz/FwUjFc9
PsTdJvhvzbZCp0q/NRKnO/4OmlHVgiC2PbujWfZokULL1ozWpaUMxZKR6ov/
AhwkPkRgkVZGu4/8UGm3SCmUb4G/IxXHS0n5whmo7kqb6QQdZ9ehEPfBUn1y
DgnaoV9eU9gOXFLRL8kXWS/FtEww86RCBJPbEADNE6NxvEphQc0osEZMC9cx
QHcgnxQRn1Vae+IRYWxwYaODk+zPESGKR9vKBPY9XCfurgBF3UzDFWG3T2QO
vK9Vkd17Ar8+15co36U3TQTAFdovLh6iQdwTZ++3Ea0kKwfYxjJZc3OC64LL
7+jGS/EE6k65+fHBiUeHBRiyuSHOdKl3o8EeK14Wwf0pV761UHfSW66BuV6E
DNCSYP0D0BtZBRsLFz/4ewSrcgKCQFzlfRop03Z6Nt9xZWb9N5fudKg/HfNw
HgTJx+kFYBco2tiif8UvFjEnwXZXjKSylalP93wHGIhf+PgVGX4IZ7rebGdy
jToJcRC2W7HFsolBXG4G18pWFR/k6JtgwiEcIXZxZ7DF+ILT6vj3I3F/Avt0
KhPaowBzvHrpU2ugRYcwncOC3p3isZVokA7meORdzEynGpkNfY0rBFck4S34
nfMitwrg3+9BXLyVgmhU/pFfBR6yNsFDbp57KcWCI7/rcWXTdDfsiYILKmr0
sR6s39s26jQPWnafjXzctmNz9FSV3ZBaKHaLfu5zrQFskk/maQc7UAqUYkqj
1LdGCwY4vzbX3j2Ta1GLHdF1WFlcsBUDEiw60h28VUiFgllFfYKzEwiy0sjt
WtIXTVE6zg+oYzO7nNfyUnXR5NXGSWbdSiGwR9WthnDbQkEuqfmKAxCThJ0V
dHtKPXKdu8K2ER0FbrGGMLhlwxVYRM7gFYvgCj04T+OsFFHgLIiJ8/940jNy
sAHf9iTwZ04nJXDNTnyWyI+r7VBh+miukNFFnKEUVBeszTb1srA5GmKr95wu
qeVKX0WdXcop0DQBeJR3pmauL7t/AXUBb9ErHwr6F7fl3nSQJrWzvf/GqJNH
qFkE9SPm/CEHwAu3w1LXluZ+mJ6lIgwZFvTJGoxViusTNoUDBNDn5olzIcvQ
qV0yQAaj9ygDI+IV2HhEvIzSGxixdObFa5GYu3VDYBmokpmcNsBm/fKx5MGO
LMqAHjwK7ghdF258QB7xNcR4s1NsX049V+yb58DcErNICCHHJ9OjUndheWQd
/4m5zIcEXoWmqmjAL0xdIS91Cl4wgVqjePk/sjxl8Isn4ccPq0rTLu4hnxEp
XOZwjAziZ/aBtWHYhqAUJ0QiHQWHK83XQVzNEqAp6jDxxzmGkLzGSry2BWBZ
Wlp6+M2QlhKKV761zlKuc/toLlNnnvLlDBfwHfMXSAtiDTsoRVYY/jcW1gYq
Y9ZnWmWF72axwf9Su5ecVvf6QH0G5VGVG4qy4pfW5d4hTRwthYT7X8NN9eQf
KXGHv2fDwGFuqwV9414/mX55TczAdCWUiB0hMYqiANts7u4WLHGEpiJgwKQt
C3yv9XUsGNLcyn/R6RfL369vBbPkXqb5LU8zEGtw8vXlJ6AqLTAIgBCaEi4F
Q/ZyiWimbW2cZ1yiwaPFkGtpVJoqTwAoES2Ji26GgFuEbX3NOAFcR8baiL+b
Rq8bN7NeBEBKL60ZzDvqk+GQ/6d78/doWcuBb2MgCLgL10oYYXem/4TifcEv
wZuqVEYToVQSV5lFXKMheIJoB/DTQOQ3TuOYcI9LCKdMM3845p7PP5FxYsHi
DQfEHsRhX4jpcRFYYazbAa+a6ud2Hj6uvW0Vk20RnOQWTpGHYj/lW7OmEqw/
4ZZfeJE1KWswgoFOXkeAOYECmM7dXh/96P1tEHgfdxNcGg+TvNzvtVGayxGn
yL2xQrsrOxilh9FZP31Yf7vQ+eH5SIf0Ge4Z+OFOXQg2iNMTYV1Sl1fqxDQd
yIRr2ITi0/AkZ6S3yHhBp1VaC8gzTVtiI3Ukm5GOGDfJEPitGHp6rHFJjMcC
DJbRvq7xwfb1vi79GK2AfDXtBYawZN4VVZyXvzKbe4k3B4DZ9KaOLOyItRm2
DFr+K+a343N6vhHpTCeSlysoMcA1hBKGHpncGc4tmgyBbii0ITMB2fvwru5c
qkcAy0kcPiz2djIvCtVRu3MLaHxcaoJYA7VLjRQLnMSLNinHYHv2gg2KI4Ov
zgGKQuENuXaMgV0zg1RQd8WGLuhqRnybK/am+9vFDPeZyMzIynd/xl1vnvC4
H6MU2IK8Ty8e5/p8cN1wTIMf6FNhscxOMkKO63UsGgAnWF+UpxIapQ6ZYWd3
UkUmOsBIXp56hD6IAAiQ4gqHFstRN/OdT95Gs3GfJW24dHSWlK/z8pMyjZZc
BPfbc3ltwOSb3xg/+RcqKkwVF7vQ607e1Syp3HJ66bkXZ388Chn82zsMmA8J
s/qIdRSW5ZG6AZ7LyROHJ4jU0plapWq5QvMYdoFE8+3nB9tKFPsdOCzOYWip
gdlEGJ7SJ/7GVzsnnNz8Atfiss/xkLUsd8dxpHlxKk7x+ysXv1XoZoKCCuIp
TT0H00dBTkzMJltyJovKSoYZWD9bzbMa4y26CDEMGnFt3lSFlNYF++AE/Twb
pPJoBDg/K8S6u27X1rd1AocImMQ036du9kFPze55sl//E6sOftlUENMofowr
IJTdRCkOtkZSYh4W4KJc1GT3vKQJHqeypn6uAdrBlf8sXuHcp6UQ+WdLlFmk
eNrv5zvDFK1pBBxTWEskAGsySQloYTXanyRoNxDcICObYXE9U+jevS0DzD0+
7ro3NVyKzTzmIv+AFIOGogD6IY/xGNdlfJDaCZZ4egJEh/4yoFD5+hPvEfl8
G5EJdlOcQZM1GHgUvJyNsN0KvV3i4c7Np0+EYeo8lkHFRLWcJioreoIWnsmk
0uDP5NrANSxkSXdFhoXd2jFzFHAusglV6utz1PoqMK83EL6otaY41UZ61mSi
zxR6V35pvhjWtNJ9NEsPbKT5IPGdJ+H6q/rZThtxd+FZYbtel64ss0WR50Fm
0Erl+HIxEctEHyaJRDvxicf8S76y+RR3XRFngWxoVCXILbuMRBzr3pqhIs/3
LkMS+6kWkGWc+SKkEpzrgyWz7v+AEY3Mln58fuXQfWhp59+4x2a1L9pu94M9
M5zp0JpmxqDlCM+qFaQoJS7vXm+gADglk0ndfMNHB1oYDoGdx58lIBb6wO9s
8dtVHLNBpvxvEbqWp0OYDlnD9slUK888/Ou3Q4MwIBz7jMRxbTHLbqfuUclK
oUO2OEuRsUdf2yihPDojOtVz3ivD3JuWNykL+fYJnrKPVpy/Zy1cxameb9s4
1WYfoR+L73/yT9Rtz7IHo8XWwbeq4peJXT93yA35w6CvQ7oeOLsex2DhD/no
t+bM6u+upWEuqYcY/+km17fDHGiZke/opVcqeeXx1N+8TKsNxqLEbIuMBkoQ
aqMfBEoU9IHGwgblISyqy42L3HWlYGnk5hFoiDRmMAa+W1V8z7PlFk3ULs9S
pi+FI1o5zwxHxB/4AD/c2S80gKJTSuUPCUuV4JrMl7/BDO+noCs/22Mmzbo6
ihFvoLkfreCsqTafu7afy6oGuGrtEE/eSrcLo1ahRV8sgeRRXvFRabzbxyXu
2db9BvWkw8xUixLBVoGWw25WYICj2n0HnA6qfTTG4UGW/VJNOuxkvF9kjlGK
nxPSvslcOfI0OqyV/WopE7O3GpuXvNExKmy0hZxr0BPcUZumWauLo2jAyYRL
yCOqFvxUyHrcOXWnuz7NAwaaEOBipRvGzTRE50mxkzoQlTQdvF5vkpDBr1pD
P1L4A5ggz+FoP3xs9rfE5rxQm1O25/Ow3AMNmTH8z07V7y4EenuZuB00RY58
Bu6/eO9yTSSEapC8fhfa3K0v9l4SQyIHLVQizrIJSRbHlZ4kmFOakrWFUQQq
gR/oXuma7z9yaXjScMu7WaaMcmGfL/beDMcHayo9aUDHRqhqNOKqko6o0ZrT
CuTwSGcpkLIbXRasIoU9EWdeZ8QIdSrTjMOvIbYFQAohqJdh3301M7aHcfjg
bKTvy6L/MasOUuXiasTPjR6J1rv9GTHDJTmrsEY6Glno20EuVmD2k0BbuzKF
krkbED5HBeGo7cCVIfww3A4dRAMSp136QZCesi9O0sHbzq9D0o1QUSa69FVc
zpEb+OT8aA8dfVXdEBaXP4jBCyXSxVU7/vSoLy1X2TqyI4R4UrP87fyH9Wqo
dxWJGueP32VIw3emYvRUkn4Yw9ENqdRyNIXklUN6flvD3PeC1uasXkHIkK5Z
eupUxQunLwzBwwv5s1cGE3zU3PJT6d93N8wJO91ORkme7SoUA0ww3Xus61s7
YBU3+wj99sl9F6C+58r6IenlYImaGSdGr+oLJrIFY324ggksQr6x3/eeCHnD
N/ABmUtRVYsC2FLzkmBzr7jrBfQi2LJvT5eWb13GFBqfRHC5w18w0Y0NyMO3
gZm15zhT+U0iznVYALUGI05DvmSXfabR4mvNSPsR9+lr3thVSfc1cbyTdudF
DNFQljLZdOdkLtwR8BXq0M575Tt1RMOVJIEvqMr2A9IRw/hDHvHl0vvY5TCJ
ZqJpn9y4K1m/wFpksRG4HcEKgjZ9xp2YRy0TlQtFCQc0xYgJ3kWkQcCinfYs
++C03Mxki/SaDg5QCDBZ8omqymRYLRDQH2kd9N2nOvxIPVPNDZQpCrmajlaA
Y1YfL6YKyKQRjhBrf8XwDVLS6CNahjZecVV6Jrxy9GHNEcU2otERQT8Jldty
k/EEnLfooLMPjRaQsi4+pkjEaF45Wgip+bYlAGpEZWS0ECbxT0l1STEDdxVp
k39lI5YY4ihvcKPmUOaBI4yxdtwTeAs937LBm7qNcEo7lEQT+I8rtOpyAjkF
nMZCr8RGuSwhf29vhilY+dkOK8eeuWq3K0mrqNUqqrOoCRbfYYTUJCMncA+D
GjGXDNNbvM5Jh2QAolaUE4S68WU78UpcdyB9JN2Ix6231usU5hNMGtmlbpQw
qok2f3BZ+CzjGipGkbZSfY5nqqhzG83uDHxFtzF1eAB6UMT44xUOyNzXLhTb
3GsrGhsmsp9bRUo1enYZbV8xsWfGQ27WX6LmOFsFR92eFJMgo3/HFFIELoJJ
R2k/ACTThl/XcMWEXrL9zzFfaE9hscoSiyNRlk4fP23KbMas9qypvDQGSKOK
i0DsmUk8/MAkKAmdDDXgG+iRwq+MFGwH+Y2MLAdmrIfQcOBYxvnf5un/0JGP
etMufvEwunJiC0bid41mCZ0FBV7MTL/09FbiH4rMamMvM7I46GMl8hPkKVCL
Ln3w9LL1ZcOBrgeJXI39wNQwtMrTfR5nPm1sB6mgSeFGoVSzJ8exztFPQNLW
jf9vEH2xIlxrKMXDQqHXzoI5vyqNXCloVGm/1UjiffiNzvL+LmoD/beQ0Oha
dkZ9fbJcyZXivr4LdZ8/iCsGAvYn4BteYK0lxTXUM8g8OsnfAAKb5iTtLnvQ
bNLQ3BRE+zEK96fvhf9026d3YDtgNk63O9Y5BzueFEOkqnHgBO7B+YiVZ3I0
7JmzAAohZkEtwS81T3smC/ShIyoqfA6A0Iy0cq5GSfia2IPYI8aYnskG2YUs
KFavEwXAAkrI8cLClsEfwzPsrjlucrekM6pnyrN6urfasNWuEkV/vt3a+ZCQ
7sLyOa7bjJwZBVdQE9JbwNxuTvNMbS6xZRlDvDZe5cUE3mwKbqShI3sPryOd
vViX4Fd73y0BWlcDsld2U+/6esXB+e4F/r1uNHT9v/UZXhFToNlkFBicwbQt
6M1Gj4YABAHX/a5Sn+vvR0yaDzSi77fjCHSciYTqEl5kSTNt9h8I0z97rkgu
G/eaWTiIA08mzftLTiQNnmBH6GmLUjSXpQY9I8t9ds6QaQ0kQKWuY4FapgFZ
rwz5ph6F7WH1a3YPt9SaR/NRf2H2k8Qp9KtyQeplD5xxaMlpsOw7sJw5oOBa
xO4pUCQ6oit8KXb+hOy8F/g6AsINCeznAX9FrozcG4RH7a6u5iZ/0U8qURTF
yCR35g3bFhstZ5dZ7lobMI9QTjAIFxK8mDXbzE+Zuza65EcP1OjSRW4VJ0X1
sYfpDvh8zPYpjmtsuH9CLUYa7jdrFHNeA47+JfvPYttDrPFPLyMQqj+aMTr7
838CkpOg50KTA6QqbQxpSe9/mGEyNNYSKKuvfAEV2kUF1Uxo0qlY+SPOQFyg
CTivqRJvZv0m+KxadeLUBnNe5W+9uVabVZjgEll1RDjdk1UQd+9jezCPon4n
/ATxTtSB6zWCIlN1hAgmZKrC3x45mzoEBcIYCd+nOypc4WpahfRG5RaZo8fp
OXfyuWuQJlRccQBfAvHwOEErzP02jKCUZy5hqg2gbZqVudyr9BFcfurfgRbW
XRU9eXHHhKHnW2nq0a+qlay6T6xwIDQK8NAEmj1szsNUS0wiNYJoqTBMLRr+
ji/+TIw2G6lLNFt344/U+ebX3ZUa+b9MUoNyFf4yHSLmccBxMkuElFa+FprG
EmJgSuBEDsg5J30gko6pS/O70EngnwJMY9Ja4PQTkpyUPmASPyZwJ/W8Bvww
YvkO/6p2HxF3GAD7GY+NB1Qsh+bGnMFeFR03elnJzyGSxxG9JxiK8W/DRxZX
k0xosM1mRZEzx4LClZnKs8IbKv8Pesf8IalXP8dvLL1+i77A9Pe15oRiyv8g
w1lUBbc2B9kArXfiMOKFmByXVygWaybvh6aj0odMVM1MzolW3WOOQZfGmK3q
cSWwrUB/w1dd1i/WbO7V5vA0cATLkEx3/BUtF6Px+5TNVxXDavD+rC06CqEV
tdxnkvG00N92J/gFgpjXghJlQRpvHBS4qIdOiSC1edF92pIyEf+SPuWcETD7
iRVb9EQaN+VTUtI8vpJOQg7TjglsXETw0rdAKYOZafAJr3i4ZRVo3w9AP1LD
Uu7sJ7CbSjXFjrNKDo1ryqEiGbM3uosoPIGGYSdqRGy1UYuG2fAl1elNVnlO
9NDovoURmhzLZKmrKJsgHqCTKpfJnYKspxXhLwY5EI2Tu7p1PFYxBPgbZX1D
NsC73/s0bxo04rvJoFVGnJvSiD/AOUvKV1dji2MywoUwqY3fs0Thv4ECJYLQ
HHcNizmYm8usWuVe0G36x8VL+ttFru3HbkUUH14NSY4CQlR5gn33I7Q/gDlc
7/pD+d2XUZAps9R1+QkiDEIkqC+IPZH6osJ09btemWuYgc2agI4r0ObPPCKE
vEAzxoUWymYMH/49MsdkNq2ZbWJZr3lGoRVZ+UPzMQ4ThlfQckBrqTJ01IF2
qP7GJwjNqa7Rvq0mHo3mpgK4UCUHy7D9Ub/uzGs60ytsLK181dZk6xT7FdFt
kEor+HcFbucAulIvaeJIoY0DU8t2cOCh5D2KU54LnAXnB3YWZ2vtlfJCbJMv
qv+rqVxMRzEKZ5DyW3kQYoS2F7CWSYQfwrN7HOtbxTP+8672xhBc/vSartNh
cErngzu8oDFHGhl4lllf6GCqWOGDg+9LZ/bXJPCasC6iJzeoe73/V4d/15Aw
evIC/b2XSwzGHHYKl60eMdaqr2700P6ukoVkRCyl2DPCV9jAfVQnq/o/AsxW
PFdQA+NCDmn3A7J75eXeqyWMMuWJVtwemNetzgr+wg4DSIfl6nyl98z7iOZb
VJ603Y3PU9PLZDMrUnj5FjHSSgD/kzd1wsNhnkmJEjarBaW1JY22S9uNjxwN
qi+f5jnYmVfmoy+IRmGMb7aE6bMncqMhfCEYCL2Vx74MCTm9lSHC8EOZvsgi
sgifpMhlc64XZlt8/je+g2nhZ71vHj/GOVOpZbDc8I5AsVhXdSB6GKQKI7HG
UnDJQdY+h0L4AaT48cLuW8dNZVS+JN1NX3gg5cUXjHjnmZyzRs+a+78z+fly
D9XaDoytZKZdmLewRILPzLRt7P8Nm4Gd+Jn7XUBcgyjx6AOlALcFlLCKMykC
7JoVGYR2AX6svB2hbyY+BNGhp37gwqEEbvM8aAe5to0ZRb1NvqXxxxtoAmni
M1/xa1VwiR9W/bHMHiUwXlj6NnMnYectSkXjivSWqORMjkq+7p1hOKDeMcog
4eNqqRtjjJvOnKlFuakalF/xEASA7906kRR3u9AV5EAzXWzIc8H2/9oVWxfN
iJPBqKGTjCPWmqi7OdAjFTFVVRLBf52N3Ydi5wZQ9zEKhsvb4zA+xJb+T0yp
sUrtiWsf9dkQ9woc7XLMeXmtM+KN3iDQ5RspPIK3d3iSGrMJhg/+MomStF7A
9YdG1GFQmjHYNVoXoJKcblazHoJ8NlQdQ82RVhoy/OQBvI1p5AQ28/+6aaRC
TNbexitcJur8JBhggzhiJzxlC38M2ZSZwjVOJClH1nVk23fExH4P+RDxhAUR
8BMBsF67snS4/P9d/oupg+KtOOa31cDvaNhNRF1g3HvRbzUu0WcDTnfY1PUi
epjn6TP0GqDWVFEYIZ7AYuGrPlRy+kiO7NoLbqe6XL3SK6WTe9RQvhmLms+o
/VMf1hJtidQWU+mJ8NBAxE29PJvLOvyUzYdP/nT8yaJ9T+k1lG8uvuZDgUfD
z0kpuZcPr5Vt8uuz+ReLqpLb1QqucM9rmQxK7yRt7+ENnPEc+a0blJ7PqGQB
52BOn1GtVd+yMdJ3XilROQs72wojugw7O2nbEDw2hR1hvmPN+XUGrIGD/vWb
RZmCEYN/fe2k8JRLsNXlnB7Fpae8aKQ3w6VsKYUfYDtnvU/meD2/gJSFoSF0
wWNzicNsjQBdaHGS0+FHfYSqVgTkH4g7VExydKPhjsa6XRJzPU37EaXVedDu
CoFXQVXKEAykdFq3EIgHj9WI1jRNTxPXSuq9NMDyZZ471plOR6O41nkVR5kv
KuX56QH2jvOvD5J1EwpOsg6xopdepQifpVLd4J14wtyr1q13TKJ8MeycnkFz
nM0LW/6UwdrII6ODXkJpkp6BYJX3pGVuQWNDnKLA93UlyvLO9zlsxiyWsPN2
YBJ+qZJB+WlnY8FOS7WkvzHrqVw/Hu1pqjDyBdc+VLDSWchr030aNmgk2+un
MoIWGrNCckrbT10yQ8nDAi1XId5hfiz1upVcg8jMqJLrB/61A7+CcHGXGOkY
dCbhy5qcgcQgY5lJ9nWl5SPVQG4c420UD6L75UGlGcDFrWxU97pNE1wIGLXz
yjdPqH1K4wopGcfeuxTwRAMtWj59eM3cXi6pWEEvzWo2B6BcoOi/iJ5oYLKa
xJozGPdM8BztNOiDoWofcRwYcEsccvrPsIbAsQMfYVZxAtWM5XhjAS39IE6S
NwKEypgBeFJ4deLLT1w9TJ/BiqLaU5PT6OpNxFvSGWz7OFnxSvnp3plHVdmm
VUZFvxFbDM/VtmmZfYGvQUbSDh19Hp/mcz9hFVRwXO9AxA3a9qKg9mqulJtm
si/1JFReu/HwlCdsBDISgjBxukdc9nRs+OKyp69CIoY2TZrySYB/fwD+adhP
ylT3AQ+RWbL3SriE6Z+aL1lasz9kSFV7/QMez4cqbNMioymjF+G9UhXQ+5TM
EFWeeC67s/96OyjolYFHW/VlPaxW4kqSVOk7EgJPsPDsZw3aXEYoUsnvDnfN
LXz/TK8DJO6/RJKbmfsgCqpB+4lHARwHEvmvaWpvM8n+PJwY+cRkan8sDHME
5xAXXlQJ52iOWDPGzkpVHMkYZADtUNeVXSWBsofWwrhE0X9D6toHsBrZwK1s
uQ1XNQ7ibF+V17ZM2oZyu0X1L15+a1mQNgBwdbcJEo2vT3SDzP3p4MdI8MA7
uHqj+y8ujADE9zWxE+6Q5PRKIFlRV4Yb/2VLVItD6tr6tNFdS5pqwjqdZh7p
jQInhkHH8oWWbba0oxSy3aNleEq80Elp+7WwYSAZ8JKcS1SMgkRMKFGaHdaR
n46aB8sTroJSYJ/QbHvP2NCjmNyBgv81XulZvfaJVLEnFvpoYjuoEqaPYxyG
MxOs/W6/+exZWVyEBPqmQlHzEeHYFVzKhpiqF6sOjBMNxdigxehMng04OV+h
RKl9IZqLgybeN6cvFP+wiEgOJg+KGGO0lXHUNv1yj3uov7RJpKSEF+Snvgwt
70H9ljNP+xMh471LKKgNzqzYLUD43ypudmXMzQ93d4O0xAvRf3HiGID9MeH5
BwA7F/7DgckwaaYBvc8r3uuqIFYwzz8p04iIsQjangFS8PtkNaZGM3m1e1df
pkxNC075JghvCJ3+MIAyqe9gGs7zv7zWe0f1ml5Mknxbj5AwBVxcaPhlTBrB
bU4OBvsbRzRoYxbhh1Cecq2Ts5XrHdsODkmaihFqQcNgyBkHtK64fulLDtUQ
nAK1KFiuhOVl4rH2sOnSnE6Dkq6XvSA9xoJ3MPk5sqByhStXK4Cxsc3Ls61t
qLokvunR5DbmCi9j5Qgq7jbxjYHGvnmx18a8cBxTgEu1SzHtmdTpvU2kzXOA
Kd5twRNsh8fKBJJxWU3FoWRC75AtE4BTPcnwceUtbs4QzZacgn639TLdAuDt
aDt1peH2cH9PSzIlvIRMwgTiB/4EbvputMgweIn7zWiPt6rAqvwmSXycuA0q
KHEmYbkHkrfBPUj/71EOBaWmCasm9w09pfSdXFybn36G65Q5AsSBbI3ZNJAX
F6frb5QeHlwLMklkwXzShqxzLh8B072FpVzR+458gXbHTpB1piW5r61u+Zb+
xvQkXHeAN/9hEhTo2jyZWg70r3m50pzD7UegzAGzneEaOK/5Hn+DEnYW3D9H
LpaAjzU9COFccVCgS+nQskNDAYDevP19pT6twRg+fsiGbCGfoBn+HFwAXn2C
3fT7Tbi4su1TiY/xzi3vufjb0R703M6zLSSVpfGuUCRDzjlr9YM1LOMPWKGa
rK4A5Hnaq1BpnwtrIltL2bpBr4huSVNndSqHT+L4kgmd0LIliwA3rFElRuR3
nu8hDVgXKEzsHa6HoHFDxCyJzcjLjnZTaZshyl0Btfpd8dJvW+PcCLGggZFk
6yk8MTEo2Z7mO+Quq0IIVIQYLAdppA6xsRQ32TkoCXEjcYsBT7XI5pmhEhQ7
/l1Oyc/nkh5S9LyEW0C5qPddpAaoGvbxsDfnUaMFiID84UX4sj3x58afgIrR
Os2YHMj+qh8UWabWErqShaNv67mDDvdpYBOQBomPAyyo9K35vi94GSFuIfEF
NrM6hk+m90RbzpxsF33YkQZ21OSXIloirjXTQuwwi+jZAbG4s9ReYX1y8Xt/
BRPLTAeAEp+/I4n9rHZa7Zk1UlXWI4bBkjTiR+EvA1WeMwi3CholLvuTYp+F
YTKw5Y3LxiJ2mz6p9xPZRV+hN5HpRVODxacjPxnHoKClPSB8l72xOJ/NZDzK
H0noXzJN3mtZTCQugDjnd7ISfYLRreYxtlyaMJ2qSVdmtzhtMZSFvE0H9zsv
7KkPoYgu/k37n2Qlh6bJCqCu1AKOqYjv+xNmL7tJRnnLFA9CC2hGRD1CLFQk
SqdUf9WX5V4ycJw9Kp543ZX+RH+t10CtVgG0mLQEouuJEM5kgu7RC/waY+wV
cHU5UXC/2PgF1EjcGx/jgQ+CFkBVdhelvm6R8IbDX/10k9kmHWqCqxJm7Adr
mauyrFCzuz+7xPRlTz7zITy1BsrNt/y0B6Pl8s9tqjkqZ53Z+r+O4mKRZGSq
zYGB0Hmc0euyBhF1xDjOCfUUg5hLttqimmR3doJKWn7XoW2TPJaAve6JKGPD
WOTnnLdg+CDnU1v/WabJG+CyI6QwhY6EXwjfg61ynK9e+ZGFuo7w5IF977BQ
OQmZBocRuRFZfFEnPd0gZfTBC8hUZUWFgW32ycedbQEnP0r21wqO8+e8v1TJ
RuoABG7t21vYIujbybL9I4lbmvNIqnLWL0MzdU0TDIkw2HiHOp7mZ5az2xZQ
JnQyp6DiBXm/gn3Mh63I1nZdmDw+jjYD1+a3AWTUIZIqjTXAyzWTUEG8JVNZ
kTV+a1ozjAIQOeUXZRd/YR87T9ZCfgcxNcFvBTSn6zvr54y8/nKjW9DuEsku
QUlt3MJAjgqJJ6XicqfpHPUA/ux6dKyGF7xzJhVPd+80BIZslJtTgqPVtaCS
9XzrJKnBC3DnGDeXQv4FCPQYB+6kKL+fzBN9gFee4UgQpO3/NP+45Izg45bW
IV6Pkv0d0loGSYsSlIw1hbm8e4BNBCcBM4BZAFBzvOWJZmA1nVT0lEIMQz8n
wTzRUI+8kq9dqnZRWgd98kA0a1fKSvOOdwqpT9dKXPOSDEEguJb/KY+4R6xv
tLRn0o36FJ2R9cYsHSkjDOMezj7oCOqGESJ/FINrwqqYv2la2phrpmXTVRDD
x/NoGo1IC/0DHokEfRVYU8v+GkoxMigNnv+U6XXnC2a1horNUEwd7ZELvr5M
cG71BNdgCiopVCZyuqEhRkfzrPQC7COXT+2ez1KiysHu4s+/yOX90lbez4oZ
oPuNrvtg5syiVPZKU7zNoi92EZK8q268JIVD6MRi3zG0MmeC2mv5JwuMK+Su
BcXyOO4JsdLIu9Pxtx6u5aRz4omg+g505KLHH9OgoWUf09Xm670Uwwq6SKUc
G8qcY3RaQbnn/e2igFzBZyWRXQXVPSgWHXbXua+AoFIbeBC54UJ1EWXyuP/s
habTPmjMCte/x8glpUS/mo/4TgJqZBvTNrLeh0ME87gJpHhKzwTkv8e9VWzY
pTzfnfM5TIkFm6SUYfD+cq/VJtse9715d1NYj8o52/sA+yijPD8lrAKUQEZQ
vGA64+R7k0dVt17TkSGlzcM3Si/ETO4UAPl8rGwa7IFuKasSX30bFxR24EaZ
Ui9XUHua1N3v5L5xtyZ2NMXpyH88w6T8aNx9CUdlFSQMByXQgrDynL2ZPYCq
Q/TsgGVY0ozqel7Qs1JVRCg+PVkBruWCmDEgVcP+D/EWtSOkkz17uVBTlzAr
7IZ1DxqnXMKZXgOg1SY9+gbiILDKCFoX/oWjga5eqikzvPRla87yJmWlvU14
LjD6COGxAmuo/reoMCu7JMoTjfg77kvfHa4hg0bZmfLL7gX0J9gJ2zzC9Kzz
9dqck3aukH3A+l8bWy77HCrXhCccleoNNtLmY0HwRC6CGgJUc76027UmQ0GJ
sw6+t2LXZnVF/ntOhHzLccoC7MHbgkPf6aNLMvCii35nhdtUBt6XrPn2ZMGn
ihpwKkfcBvq3kL6XssqZh0if6FmVvSc6Rtb8sVQ4PotWaCg2RmW7LpPk93g2
7foJvKkVJYIEj/JYHb+0V5Jtm/12uPbHB/XD3+IBzsalxE8BwNgwD49H9J2+
45ASq2wSOACl5RHTt0nZVUOc+n96eIBK0da7j1PLwbus4Ex7H6R+MRXXj/cT
8oeXjaCp/EeprmNu4bOJkTFvyjcvgGiCOMQz+Uabq6wmUU30KbU5GQY5DopJ
psn6JzhVTvmPskMsIz0ckH5IFC52KdF79nGs45uJHDkZ8cAaLAR1MO4G/m/+
IOaVaAhzD29jj2la2T9rCMDj7T7cvdxVIpzXrnkhzxP1Ex29n+8gFoAuLmWw
yuvjVBN0UQXaWRy6+xlIbll0Zo6fuaprez28Hb040fWR4mSWtYvCwkDK0dvI
xVbyxb9prNfzh6X1HCcp7HI0PSGr746qGSizl4ZtGew1mYm/gCNgbL1MrF+A
GAnG6EEWyWVRKkAA3i68pI3bWSvrCktsXEd24+W/QMZT2ZyZCjbqZskgD7ng
CjBZymIrJiyqlWMvenZekl2jUoPzed5nqWWEOd6SBqjAGYQv6P9GWFVjfSM+
y/sMKuB5QlXVwFY9hQ2jix+3W6AqmUzqKxKh+TdNkQfXgOiRG2eOa9pfTVFk
2kyMlbbACGyxJo15mxMkt3dRxo2VRpSbr+ozgGg9KMUUcmNlzrt9c280wkq9
wfkP3QcoEle6cMNi5ZoJyLvt6GWDpU4KCiBNHwbRj8w7SpwlEYnc4K6zld2A
uuB/+3CaJNIcK7XKnS2lejfWUFGhO/z7hJBIwGacl+sM+az8+GNy9X6aMpM8
gL+I9RU5XDtm9NTMSvt9fZ1mx572oFYPFbY9uxjiLtV1uxM0qW/WLyXHM9gf
qi4TyrwwfC8h0XQzZuaZH6zvxowP+TLNrPpg9o2SK1JDyoKIzJYKLT5EvMOW
4zpqP4cVTTVPYKa+2f6Ebn3hwx6gkCWJxjbm6EcgzrFzZu/H+JF7wYK34nW1
rcmjZG/DOhugdXpOKwmHfgXM2cTnExXWJgPlaU+RziAoK/S8l37yaZFBXRSq
prb8swPLBFFv7K0gFHUV/uvXPqKg0eToVzgFlBQKH3Ddo7u9/+tkUzqQoTAH
Lle/jcEin8yyVReamStEjbbr4uYCiBpEyQHyTphc9ONdWaRir6xkY/TyT0gy
gsnPytgBD/rznGBNIEkPGcCP/UzJ+JkNHyNnjLQToAMQycHjNIu72fpb6WlL
BVywZ8wIJ0RqC+cpfoDOrqSc2LnQfXYoUlmagRXKbx8DNDS0s1Vt0qdzuAJ+
ZI88X1WE8zi15Ky0dYuYR995o2jO6gFcZkF7kC+D5pKgfZbfSt2GG1hSBc+H
/JSDo3L/1al+uuuczMpvGFKbff4zoRFzCJJ5bnXwBlLRkQ+zoUuUkeGgKS17
zF1jBWU4eNyh63CUWwpmtsyB8oHTkiX7Rs4k/F3SCA07+no/oIN7pRotuRaT
UMJZViCHOvGPSEjITBYmJcXEIIegjmCZiGQUBh6bOSWLXkwjTIBVUvjYU54X
moRNHfm6jzNGLGGKl6zb3YXuPw0DGtp5ToE4W23+H12B4iLYPexjgVmzgJDU
tB6w5KcIYVaxTG/PGaUOOBhRDV5S2xObGUUJc6Vg2ztSFOBugmUOuVExOQr3
Rl0dEl/RA3FHAq+rTVbuKi1nGFTBs4lUyF70e9ilqzG2EmWFX2u/MQBr8nIf
bU4LStxbF6pMsBCbVaV3WdrJAA+LhBYNzHtravMS3CteWQjx8V9J7Et5LosG
0D4lFboMdGLLaj6kIBXhCXh4e99ZvtaIxF57JTJXk8m5tJl6AsJRQ12aFOkb
TT0h0nOmP8gPmYU5b6eCUqGO1rDjvCjx0fJU9b6nHX/GZubnRyckr88Iwe3D
qSJx2SeQxc+QzGlNjUCC0dzGTs8qaqEsY2qgQmYvdq9KKcsB9BY2ggYmvAee
UKu0Xvclm2gtUP0MaQYYVdyfAD7ZNZxAOf6JtC+vB5GDuY87H1Y9c6Tswcbp
vxIiwEg84uT3AGmguwQQCB2pGPXMlbpZFcc87iqz0ijFWpYGZRZ3RAaZvViU
0Q4CE7Y+3x8XPl6erg2i2eIyZv3rfUSFd+WRFNIz8LGNABXEYY1c+2r1WI5R
U/6SCu+4hmK6XClThlSzsDj/hpdqEPTpcBDF5gaV78oDmSQxCt+NCHCE4IdU
pJ09wFLl9Ioo7LwbUfSwHmnh1FU5sPt4TJ2+TQvSEWcVBG6i3bzZblFAbkYP
bCe1BN+v5zKrC27BHRCU0HT+zPkZOTtF13C1PtwMp+zASeAG5WpJkj1nFJCy
yqKozBc18UWw8elz3eHeW/Aul1rGaS9ENdEU7fMO9cdemb1vf0ViBg/Bs+cG
QP9C4P5sOpxaW77hENQ78kkx4qS6lKKNH0Cakt19CMWqHHwwBAUlg8D4LLN6
MAqJzRcGTTumNL08pHzuyynP7WQZUMYmNEjLWexq4c8KcpJ1AaRHGL8WR3I8
yOCatLRibBWxx/k1TqtQA4EZr4a7k+/fB/WTkoRTAQwfrcnpLkklyko2W5Pt
NSAsZQhjZzw3BgTHbhtXIyGAOvDkjPCf3uCT6o8nJOCyV8fWVurEwDOIuWA+
/ys9MZFta+bwR0Q6VNNKLUzBTgmL6nLEBAWvwS7/bRVcB27BvsB61o7L0MFE
vLgQrkSLQgJMJo2DGJzGW2cDuNcKkj9RjZu1A+mRdCa8xNimkd7PQTgBzXXj
FD6SUoHm9bBxlQaLSXj7X4A/vXFORj2eZK9DzZL77V4eAQ+6s3XHaKJ6K6o5
hz8XELuurNZmDnooYAe4+BrTySUlCjqGyNk8suRHNHhIZNNDXzoSEyHCkQrM
mszNz1t5qJCgGS+5dpRDR/eU1WHw5tPhiODNJxfHIY2qg6A+EqysN+RDCZib
vmWysA9zytn+ZfkBl/A3ZIHjwXjUMgWI4Dgh1HNLkmnR0LDi9HQKRoLcoQ1o
Tf0y24RwRDsMNrde4ph0ig/3ImFmg7VTdi8yU6egaaQAhaKawbyfpjFH1VQe
E1KdYyqxNhmB8pnLpABUA/LfQlQ020ZzatBQz+3GPOTr2TRbSIHKmlhlsyvO
4P7WHq2lNPk9jH8tFijJLWxHQHlI2vcnAoo5h2ht0aVSsw0NmYnQgTIA6nrg
M9+Y/QlQ9TduVB3Kef8khGHzVgNtEhaZSJUhfpRBeXnI83OlE32qAJ18AC4R
bwoYf7ZTCp164JBk9QkQgq6j5hSqIeshnwfBzL/lW+6WHPVbfbm8n0Xgo0oB
6K9TOi50+zfxLEGHQl+/PwwhHov6MUrQAU2cnPxz33w3PwwREEpHb6o+z0nu
l5EcX7TnLHiz72NlhG1Acgfyu/+KD6L3X39aww2AedKckG9fn3ub9BZtBFIG
hZ9Guy/ZCw8wsZmaEknm8VUMX8iGGASQFmiegoRxWNEmZ+ecLLXuJtiqg2MM
Eh8rTwxEuibYn39AVW59LshGiRYK1erH8yMJ0TY5w2lEEPKZVmq3k9M/knIv
Vacl9l076Glk42oNz+FqDc1nOY24T5cm0sqr80BEvE5NtZDjZA4QrMEm7cnR
bdICQZ1fiiNYqfz6qhWNalQ0DQHQ84d3xo8O7x80u6oBgfSfY/reLFNlSAvd
EWljapGTp8stATOKF2v5E/5VycDIn3Bq4WMzTZ2PJiC/zvhBqEstVPb/F/7n
u89MDz+yg/TwhbmSg04/CfCc3Rf/TuJb4OCKncBYCiYlSOivzj2YiRHtMu0t
5ktKQ+/+jTV4VC93As2TKZUMBe1V2G/hYQyeGlQeNlFXnamxaOa/idmP2++j
LBICwo3QHtPuceBm7NJJjTJdTTkx4V2rCGZcO3dOjg7R4yrp2vPVpb6Z5zMD
RgTiU5WXxT+Pb5wgniRYxDSibgOiyBgJBv8bMnPzLhRqvMYusPZOWfj9MOPv
n1sBcu5biPbYYSmVbsnLycoo19gick1qX2s+XJ19kxsM7Bh2ob2Nq4J7QSgu
bnXaIgLn7Luqyl/xl8o3tSlfP9xdYpKtx5PjOmY7wvMGKhqrObUsS99cl/iJ
Dp+frucTnSY6M/qQu6UJqK8JqrVnY4AJAKbKFq5SBqu7OBestcA1/4H1jQtw
F2E6sXl8AEiqMvgR27HW/NPKQbdbkAVG+k4TrE3G3EiJAf0Yj83rjd/0QWTZ
JecWLdCMK++6UlmVDbMSZmtn6UM9f3Xq9FoT2xm26RCbiu+jangbvNHvg5Vm
xwxtHsxVxI9zvlnlsYetAusuGyWZGmuSKdA2jQQC27Dm40TL8Ir8Gih/EV4H
eWPN8AiEIeEzOC0uJFYV2t/vemJzW8obC03qx5nHdB0nNLjT3mPrELCmveqX
q0Q3pVMF9LBAL47Xr/KT6QozyOC4bZ5CZEV/lLDOoD4dnEVlVCfZYPznKSY/
n1/yl2bEjyOWvSj6PevLPcwbwPl+u77KAf15UDGQqmc8mf1bLIF69eIxWHHX
+LTFtlIsEUSaKpcLGvSXauEoc/j/UZbT1YZessQ2YaGCEMk87S6zdwwz8A1g
4ZyGuJzK2xeS0I4e90mp/w9g24Je0iA09+OkQ1n62SYBl5/o3tbFmu8Unv9b
VaToJuQRJyp6q2nPZnUHewVQNhrnorjUfyHVfWA82T0eApTcZ1pTioU+VmJD
8WC6+pkKrFsAvx5ZEvj/TtB6s7oyjQ+Exn7Lm9Hp3pzeiBy9Xnq1DvDRfBtY
5zEeC97FvdwZi8tPJZsDxpwfm5XTZTTGWE7m216MqQORFU5c8/NFP1P71P1K
GsuCie5hj4ERXHSznmiRzzwRKNCfoql1sCxK2mhZ9ddTQRcG0Yfmc85sz1Rz
0LAM/23UlkYJhnZ3LQh7x6GrZQc2Xm3OgJV7JiAAoOTa0NTx/sJDSXnVZkYD
QZ/dOEWRD0JBIZNOXw1/kuZj1635ndRk6a9QJjsRsOHD4bkddzZcCtnmhqvr
8+GdMV9BHwk1mLVZGsvCkJ44Nz9osEf+kHAJ3tSD3ndBe3CJNDLu7m8bxkuO
4gToUeWJYzLIJ4YDGiM+seUdw7Q+k0owETyf5JBoWEGzVPSBRzesaDoLH6ps
4mXxdc704EH3M2ABwhE9Tyn8vTJCZtb7dK6KpbwCjuzcpZeOwxQHWV8EGgTC
kkO+tWY9nn805vzjoy0FfJezkvs9xHTbDUkrXiKhYvW4ib8hRwUjQzPfv21+
LXaow2/N9C8ZmhzNyzZF+yOb/0KdkaWzGVB7HtRSefHdz+glYQo7oOqesIDe
Sk2G5u/h5PPnN7yimSXJRMG1ACIhkWyJr9ZRegHLlznlvvgBssT586F4Komk
opEHCDL0+pbPOminT+buu84Qw/eJLlFAWCXdhHrY76ryxvP329+kJJwHVQi/
uq9sHHgoIun1F4K7lXWPnZPri0YGXy9+Rw1QFIXCFbQq9GaYaG2cabF237t1
diUyEMunSP/3CZjy8rhDSjSXiGj+7nk9Dnb/w0PaLr8E83LdDBIXjLaqqISB
wNrtW+oZzg64f9vQWAU6ihUAXJEayXfRkC+twf8w6DBWwOM7jngy5I5vqIG3
8X+TIUXcRkAitmBgVm0FRfZ1/NY0YioAktGfLl79MHE+kFcbZZcf0SJvr3ab
Yy1q3/drqbpKRLfZqcvIwC/86Z5UtkSb+wiZ1HnVKaHXJA4tOBhV/5XVLRUF
zoqmqQ+/T4QbDv5/sAveLQgK0zY8nUM6BhOtrG9QkvU03vLWlFjpLxogOezK
FP7Z++LIWyMVBPJOe6uO7Z0HWp2Uf1aW+1Qra7xH0ZB1wZW9t0SRnlQv2mlB
pqkt21wnyd52OBfkzlsIG410UbW52516pvEfk8ilsfhfS6YDgt0MK2NsAyz8
bjcAkXJPtL0QqPzLfHMStc8GLqd7Bf0bz6RfpM4S+wOEXXAX1LQ9m6w89tmy
LU0GDWdrqvsvfed6sQ3h7nO4NZTDvtq4GMj3j1s3O5S4rucli3WyFS7nSFN3
hWxXSchuvuYBjWuTYdlBiR/PC/92B93a1j3PB5K/HhqSJcP+CKnUK/CQoZ3K
g2QqRHCFksnhKrlKXB2bFccn3uqQiZ+F44cCtmjh1PLsVkylamsGGQ50tkgj
fx9ylII9/DhDR+M05GUjw6Pq3FnUEWmFhdpkINPGALnu76o2gzI2szUWJ4L6
z4kmjDnjoIfXRjBsrVSTvktOS4OixnPZjHIXR4k3Bui07LevEIjePFYXGlSV
RrQMnwXvSdUmkPAyXfhKx2JcqOdi95yXSLbHUwqKB4I8tIF3wFECeeXTLU04
E3MPbfhfoK2Ey0CaXPuKAsGl4q0Mu00dn8TT6TKbudS+5qU8k9b/9YsacI0Y
m2AXopaL9kgjWB3VBW1KBAiZH0PRO0EykxcElxAz06J6oRbSUDdHKbPRRx9L
zMH4NRW5lqcWD/fDRohQvgh9yerQjeaQFJ7jtUBJU0kqsOt8nGFW4cFxVnXK
jF2QFzy+nQ6roFKWMbUbR2q81Z5Z4WxKKyXuRNmBonj99/hNvZ2wgjJfAP2q
jYucxZ3z/GiSEOB99kWt2PnPlGpeynhStrhKM9yZqP5nbVxp3s0qDeQa1mbD
fV6VWwfkYQuwhwF9iq3yDmdCY3Hm/FMvfHxKaJrd8sHZ1Rj3Fq52PpzKeTta
Jp/vF8rGkdgiOkPMx280VEdWl2fIWs7o31A9hPnZ5CPBrA3oTXLnEcYVvz/F
Jwl+g6Po3FcTOOu7H75wHs1+fAwzqRgEgk1cPNisB420eBgmraMO382WNbjD
XnaRS0zNqvo7whCvjssLudZgPD6bzjatmxlI59nM4TNr6NVH1fHTlO535AEK
DCtgM2gdDJVe7ZgProupq1v7KPYNT2Gyp6YsadJf4cbvSYwU8dvIbJdMJ+yM
5cv/vpKiL4xm8H4nyhhsAs+F0jzI/uMIl40nijLQLgeL8gqqSkO8RmPMoxbD
UmNtdNrnpevbpFPZsQos0zT3b9hKwbvRq/WvUkqrMKH2pWrE6ZVAR/9L26+g
4XczIDfQc8K5a9zmUXDCyuH9dWCyWXeGDZ9nM0e3+CMx8fs5xKv/dp6Jk4Oj
F0egtI7StTQzqVR2s/Vk7fgh5SUoGGNyvlEiIXZ/eq1iUUzaLx7pKpxazbzz
D95yEjL2rIOmvhxedbjNCuDYqlLySs8JuJrYHGjtkdTFxWSY7Qd0smgakfiC
XQBHOO+b2PzapldRQ4upiHafOmuNxEiVkPDBY/T0EUNX/+W0yy6qVG++gapB
0HY82tRUrj82Ueq33QmzD3TACAcZiFiWo3alebY0M5IDETAcMJKGWJeyma1i
CsV0K6KH+EL34I8fuqG0aIGdr+Yde8LeDLSMjDC6gl903A+vO5IAzQGbKpfl
z1NMIeMd8Tv01Hwx83s7DuGw+tg2R3w1ZoLSaD9dcpooLHo38npKQpOxb+hW
CaJwAwksgxGyPptkjc85PrDlAkg3+Des7idUR6T8I1X6SYOlA9Vj3AQDZ7zQ
EXwqSf4AoMNjPIJhiunL8Q5EY0MxRyc8Pk3dMLf753ndPeWYocCNAB8WDYY1
86CG3WkGTjCmo21jDESOnXmmom5AB2gNuBG2QdFAg71lzLD51XdDq/D9jWYA
qGuqL8d6MMlROO9lQt2k8kWDoV0c5c71nlAOXZo5xBRW7l1T02xzMvwonFYL
DNPbr6r+5o9O9NV8FmPguYP+un8Z7HdJxHCOJ1c26llBUJcE50Aao/iPbmb5
hSM0HTCnlmfG316Ckm56jomlCAOoAXpu4NIQteWOv6VcL+hXfHiyzMoN6Os2
mKROGa9DGlBcORqNAnLQBak1muIVzupQhkoAHMdtagZPgNW1oqwRMmxfoNPs
5utjr09rjYWy3sxzjaXtM3e6Tb0K0z0RfMy3UYBKpXVZDmh5tZAhhfTBLjnt
kQrX4jaQWfm5+mjuC4T2Jvo7cxhyxzEBNZmfpqi++eMcK4ACIuVkDHMRtDzh
RytdUdHfoBxZUbJeFKz3WkMq0eDZdQ7WqJN5gT5ZqhzbsPKFObxNzI/U3E2P
NkWY2yFl2GZmUmTW14qZpW/llZyfYxaZg4A9lLByUNRQfYtOUz0OU/Erb8AC
2PJtK33cUlCfBA+7V4Qt1YsiJv6b7L4f1NdUFlMDmlEVQUFpYKblSWsKdgrD
1eKcuzav35PV2h5rQ9i1UEWulm4p2X686AKywK4dey5jksyG5pbzuQvMFDqw
r9JmUkV7Ift718Z1MBJ496tnBEGVMtcQhW0Rwaxsn/S91OXAIo0bomICLpPA
BUYrpDg0i2hbOttE44k/qFpRKs8Bi4aY4vPDCG/nRkjD/AAiaTbh1AbMauQw
2lbSqy0sWR64KkWIDkjTDB+keIezmoOxzNfXebbcLi6Fo/kKl0AQ8r+nLNXy
8TkSyBNXsZK7koL/qjDmVuOSKwZAAAPAzazjlHhUWy8BhsTt8rDsPemoA0HI
dVveAWw0YzEIznJh+TXarvMTNBmYUphwby6IdFn6h12xGmizP1rBBlmggqTb
qrzUuyQGzyFmgoBc5+OnhenoJkjHgMkE7kSaXj48sLw0Y9buuhBxcqfGAWrT
vK5s669acisF7g7Hexa/o5OnIu3lB4k6RZZGDg5OYE9rUBfeHyjadqSbwdbP
cN2R8VokyP02rScDJ/c9ZCIroYr9CLR3xunO074wm1T3CYrWWH4cE1N/lpnX
/sJ86MhseMeaHPTyLD5p2DgLgL9McjxIyyzUuqY/Qd9FKVfzMWY2a4W5lyYX
WjTPFJ7BjWbwQ3HPdccCEZGm0z6GQ1h4Eilpz2Icul0xyYEmZzxV9dlnNDes
N31aWqkUgZYcinbRGKJVpedbI76HbYDCBrG/WWSA0IGMu8rh0wR8uZdLfJn8
lKt6Wxb/UM1oLrF+VGbcUBX4ozIaQ+dulM/f9vgoGrQ0fNJv+V/amys6swEK
NKPZu5j9r8cy51jYvA0CAmCFjp208UwN/OY3v8Vjpw9xg8eoI6v+2DinEEZL
DR2I7dKwuNjBYKtyWUOZLpOnsZ+NPSY2AICuZQI1xoI/xbjMEgDuEclKhS0R
FfbF6E2DWM/ZTo0HnyjTUIIZBdD+YskXI2ZxSst/H9US7vrPrIBMJqo4WKmQ
2veYCLe3kpzJ6QOmnXYZB3kBHPPGfT0lgszuVIMvZBWlAsgtJcNR8YoJvKKE
VNEH78oolYbpEn2bCw5iCJ5rV55FBhpz6XdlQyhM2rZtOjVfrUWiKYPdxo/n
UyrdZycRVBn2wWFHGjiSaew3UQDKp44p2ueRT0f+7ZUuxiiiKpmhfgvauPEf
CB3IX7eT8JkoRY/VJmO2M+fwJiCPtUZWwTt/ZjdcdB9afVKI1AS3x8Fm03NA
7a+hXFXYY7nj7edOC2dDOlBDnYsH/Qnxd9USUNDFrLsmu3J8Eky0FY5TxfYm
xtYYn4JPTjhlcvUJfFbNiCM+Cz+sgB0n6285NP/O9BHyM4AdYSaU9Wyn5RxD
u+CcbC9lwfPwRpFwnxJsuqQsEj6o9CyCl66mhdMGA/XjwVBkfcgRIJlqKxel
sTTPKyoACMGtEFZEkfgUaTnvkN2UBI42oa/itmYYZfpriWH/GesioF/k+VRF
xwhU07/PpfIhJcc8n8SjoTjd3v+GhVoaRn3kTL8oZKbjWnhzdvGYwWDBdGJH
Nj9250gjsR7ymTPp10QWE1Y4est5/+UKAjxJ8B638ztbZVu0WZkT8I4hchTz
2YmvnpXbO1GdG6wGIjQV5P950odTL8dqqu8g3Jc0VKUmwqjB16ihfsnn/ss4
DW++5d/tVPkSjvJkfxBdb2xA4Iz6TPGGpriNB+Edfi1eezhgQXmzYxGsEI7q
Av737NAspYgIAfjfmggOSxMhbWBuyIyD8NBC7vApVrkgvCIq+sZhyW07+Few
ae0VfW3/StDqe8NKNwsPMd2mtt4FRH3f5sDoD2sQRK1h6o+UGkmvldU6A7ci
J98uuvwEM13gyMlVOTgtirs7/ouvqSoxkNdhSMEiIcZF8AKUIRdCCqeFa259
OnG93HKsUiabgfb+crFGOefRmllV1k7kjnDJ0+spf9EZ0pjHBimh/i9SJqTv
r2SU6JN8HjArZuodXIMIOVv6mKdgL4ZiKNBiU43zFAzqa3WC1jZvY0APTRaf
7yqpdBBVHHhhgUROjYoja2u34vMgMFLvh6bAaLDPw4SBY0W5eE8a01cjZNu2
Zvx0cE4ApOopeJaCFhXIYez1dSKSd/HYSMH7+KV7jYj/FJ2I1zisg3VBpEdl
Ftuz1ln2ANrgKeDz0YDdrKlZXf/PxAb4EAhNJbpzYFyczvPrMCubdYDqnwAQ
crXDesj4ZB5xrTGP9VOitIHq7xCmAXjF/XsUyJ58a51l6FbsARSKya5uR3ol
0/nT9UiSHnND6rR70oMGCZ6mtocrqmFGBEosR+hC7QSJFxq8Ds5+z6a3t5hl
A0tn8wjFHShvR0tdWj4IogRJOl8J+8zV77RpGsZ92vFPV105QGilNV/4cXxv
rbTjQdgJVUljCB0AK5F10sOsF4zITcZTj12ktePrnIsbBF8lsvZuioTDtPDw
y51Q45wa/3ZyScpHanz+Mvw+vQknhh6G+2JdPJ2jQOYnSPC3D5Qgl4C4941P
WIVs4iL8t7Ps5yJyPzbJimZNcwCnZODTSh3VCzuiruwvStBGBbe6rtRki7BN
j38L2WL1QPwuvp/gkbWKpjaHJk0p28Pr8BpUJl3e5qCbr8lRKpBatNhxTXFF
avc2AUscCbZ/MNBc+OpG4mOb+GFiJKrk5n4MBtdphhwFgYc/YcefJE6oYDyD
C9fTTpUB/D2Yo4+og3CbGvi8m1QdMd8nwgOsER9InaX+9XhvUTATtlHF2s7c
fhWC4Qk64GiHmOhvI/aRGRosofaxs5bdbTCucSczmNBPBulYc9LqThWfdJDy
4orhTyNSxnK1kJtkJV4RVS2I1BFJUJW0z09g+SgUkt8fkEBKx+22byviFab8
cx9vUdUlck6ACkqAwJXWAU/k03s+W/d01LR9cQ9ank0jLyHEtkACIhe7PG6y
4CLk6nCPCnockix4y4Vxn8pVuoB1pX2lFern9oRBNakfBr1GYcZQ1MyzwPNs
q2Mv8sBOx7Z0R0Ly9XJrdsiIVtYZzaI49BUYfZcDRxifmnjrmDTy0YTknKGa
60HFJbuzYo9QNVYT68cWPI6hKWJ7fKOl4XipcFGDhU9raCdZFrHRZr1aTLur
+6oeYqHjQBFI1vHdhzJNPGPYVw76xVh2kNUfLIoe5QtuDPxIzlb1yG+UbCVg
hMRBC5VaagFqBzm0xAmcbKSTQf3RM6oaeGEGL9PTv5bndBuztQR48lB9fSWG
dxrTPgP9tYZB9X+qcvL4wAUVexzi1SQAUaXVbE8j3QLAnZ2W6LZmP++vVBgg
noiYnC7C1iaO1VPRhrCkcDWFrVOTUwUoUZHUdC2nn/walnHYW9Uq1En+F9Bp
FQBqF1Zr+NB/TJQQDNZjzFSteO0PwejJL2xd+bY4rmG9Ev5c6L5aH8IDr5Nu
BwSubzK8JDX/WSfIvfFIt/YZUEsz1TeEARJZhyZAbaUybDHq19bGcVanbKwB
uADr6hBdognA/BA9w6xlUwUOmAWjZAgvfcI+EWCWwowfU8rD/1i4vzTHhuoR
jMiNxmm73N9y7jDhRT9+h6LwN819eDzooIncqzw+f3LTuvJ/o7B8unJrDBu/
ssjNGLJBw3wwI+iOh9dymm/iXb0waZXCMNONsWZGNQ4K+GO7Pzcrmvds8PLt
pe/eAKpPYg2gXj+wdS97uYDcUqIJaFDT3/4+Q75RlUctoIGVWiYihSm4Wowx
ynxOFn05+k0u9GPVGO2arRGhnma5S6t7MHZC23Z6Qd143fl0sJ5Zu3++RD1h
Soz854Hnybftn3WUWmJNy2pqRQbsEoFastaEJHhA0Iiblz3AfYJiJBXngLwn
Dq7jaUP+ATyOjYo+tOwnMge27Jxp2YiIVQmD/dlBtW/Nvks0hmPC5ZKVSHry
AAwqT1WFGJWhfbzVNo1HY8jZ5h/m6sLRKkCtqvsrGUv88VqwzFDQIybsV7s1
QCTJsKrx/slFTDaLvJjwZFgLlxAvV6KASx8zJmGXvdhnOkwDUtuMGIjE1mfS
fSsu5K2TCJluDdshe5l0EWWV2b6pZMb+YVGvoie2fo4v4QvmoHiRtqZ7ofzp
ApxgM2RhmtqB810ShxhpeMUFpa5z6Hdl80Pu8Nw1h3J0fj0vWihyRqygW8iW
lRD10/Ynusphxe1DFvUUlFohToVRDt/mGWIFRDJokRhoLIGASJ65L087Hrg1
5mUGI28GG+NRdzRM79zaZiwHVYefo0wpmNvag0cz60PddJU42HdzAQr27Gcp
IoAwayExmGwFj2j3JLVZAHz9OuKpdksbuJEeuX+2epUU/saOwH8tthSLdN/g
mUUq87uJ+ZlyHfWE2IJADknzlmwK8e4qIkWSqY7iW7LPrpZP+tOdb62Ht2oT
GB4Y6nxVrHTivSUV34MEppwVjx3Wq+lQ1nMH/PiQnyq7JtUWxMz5QMoq0DbP
bYG6U4BOHQhPUpQWCoQN1QY7GJ5dkMtgVg+FGTnvuDT45UdU+HBDg84QOMoo
N61H3ciHrRrm2Tr4ORqO7KS8F4WAbWt5kAPlhLIM1Xd5vZm7oo3ra+GBUg1A
WIqTPGL+dDw3SXXmG+itZnK7l3Ixa9yzso2HFZaT/mdEiD26vy+cgTJUt/nD
DKMnIX1/VLvRcglfXCyNViuABOMLdDhlnQDcrwCrfUU4Us/+z1m+ONfq6lk4
d5tOoZXyHwLcWfP9NfomMquQY3kWT04z+0LMkCpf+VUrYve7nIGPCPCFuqqo
zep7liQKkXFW8MUbNSYD4sPxz+EiPMVuWwFu+u5djO5b95J5qUJYTQxwQPgH
qUt2uR/dRvW6tDqrTpX1RrqejmkJeDSMoONGi6THRRiHVhjG05lVgp+iHIvT
2DMwMkTaz1SggaFUm0KKP8XQs5EDzsGcvs/evfT2reSh+scK43Xadygk3vdi
wdJVI/5ML4V2Fkh2KHaoQyanrTsBlNNgWqSUAOqNTsnAYYsRybpMZ5hGOToK
OSapkaFtfp3oFcKp3YxWRDwF5HZa6Fy2WXVPxKrhbrEFoaB59QRWVnroGj4T
8s/FPcmMI7ycFYRtRtalAEWZAMae7+dc1QBOeX4FxYYsTeyYFHi6Iosc5uIv
zecCl8z9lFBj+Tyyptc7wHS9uOzJlmPOpZ1ISB2g7Xf3RwJjiGP7yccUCj8q
9bSbAQ/klcqpuTcgPy8Im9KLBz6mm9O6Bh/OsWDsTF9OmRjEncKkhyzNXQI+
OQjStp+rJ+q42Tx5QPin9GwBJbM30RKZmzyjqmhy4AsLPm9LurEozZWtFwzB
k+DyqnKHSl6EvNVHdXhfCjUFXfHgC/uO0ItbnhB51NfM2dMYinyXV80GhYve
3Yv3Dr/KSUUEeBOY7/8NstEjf5x3KbKT+5Ma0CtA27WyccD62HOu109OYoDg
5OG6nGivXfEvUHEM7/+Hp98SNNsh4Fs3JDeyBQoKa2kViykEaBAd57oeYrHA
3nSF0MSKI9owYKKgsE9jzvV6igwgD5Y26GLkxrlKD30jqHtjtrKOACXXo2I2
0a6VUW+qlx6njdJiji2fTEffW4AZioh3dOQpn4/vIyfd5wcFZ4UWIFKIrtu6
YvL91hguiAJurqqloLHfvvtJQfPUqvXuFUGIb/eRkdg67/uxbLW353T99UzL
IdixS7UpBCp2+miUxHeNg7y9aUL5Ud/W5ZvR9sZLS51Rtcfm9QMF/VBb+2uu
zpagd7SZ4wUbwJ4fokrR4VVdqVzN40lUhqie3kSMkSM0LklpK4uWEPd2D3f2
VNCSXRriBSX6r9dxldokpYAryFaQpXbU8zLsX8quVMfgwlvuKcCx8eQOOlyv
F77W7dFFZUW0qg50eYfG2ZldPawqxa3c4w5qLTFDYH/KioietDV13bFWEQaq
94ruLOdbj4sVFB1gex4kjMuZ6T8WEAGzsCbFH2nhOqQ6+00GhmVYQDtCC2Fb
uS52IfEIjfMzE9sirf/vengC2qpEInUPK/Zl4FLyPLzv/3jJsz/LaLfqF1Cf
z9UzjEcUsD9Vt4PE95C6Ff5ZHnZIyq2DF1TGwfEYEyNA/WIdcl863ES8HQQo
O0ucSL2Bysf9I4xfgZsLrAcnTM4REfGXdI5N264W6Yh517QL7in0JkVNagUc
M2Bkb5lPQasbSts7W3MBLL1WM6UUqfMH8t+UpcLR3PvQ6bI2UVfLL5nwzdJU
Hv9L8vk8V95Utl2HHEVYU8J3eFKFv+2lhcOZWhpoKCnauY4xez0l2F8jmvnp
wZJkZlMiSH4irj+57xUrltD+pfa9K8w+pWXzHJCtbsb+z7ARrcnxDo0aI3H/
dbJG12kDFaXi/5h8nDVVA9/1lMn6sWnvI7hQPfnqOCy1fuPrCtkDhvCx+c6L
lheOcGBDUwtJrQ/9Xu7YxE5p4cIBw2cQY3yvT7e6g7NIvE0j9H5iTHJA/Dw5
+qBKg8bTK8KQfb7yLZdktBT0xnjSGuTbT+1ab1aSY7PTlNC5R7/2Qokc55Tq
lao705gI5ExpRj3vY+XaKCuFEdL4XYLf1sdYDkz1JJn4NsrXn1i5C6B0Rn+2
Lb1bGGEg+NKKeGvMwBtNENp3nWQ8bmTn4MNkRgH9G2XYsxlRMZX5tUf4x1CA
6/GG7HhzEF4cXm5o1lDX0SwgHDH9cxgJBfBBYfh5dArchJB3cRUn4CUG9DrO
wrhrU0QkJUau/6xGTPp6cP9ZYZAnRhDDfKoGmWSEFNUkVPvZ+l2pCtsW8R+e
awo+BQqWyYOy1KaKEwqYYA1lY3OOTSkIN3sxWtStXGp3rz5dGdpqu468uZkK
lfrvITAVepFQlCp/+4oZJb+EnkuALsYmL7V0n48/0Arhh09e9kD2Y0Ep71oE
HnwhLdrp326xHD8mXaUo6MihV1ytBj5LLqIuLhPj2TfTo6rNSuqJhEOt/e53
tBDJn8hReTfpgSXD+4AstQrVHKZnEw+vUHsYisRKIfqtX+F96CZxoWJpvDW/
7fEJVL6oVfkxVIdbehtE6SjIaKHhXKbcIKNegff256Me5NuyLpyrkzoRD+cP
QTDfN6anOdYwTx55gqxf0r4aH2hl5GNvwqoMAcEiXROIXMMU5elFdCh9ze02
LUKRntxX5+0GFfjI9maQFTWW4tfFdJWStqrgA/G4vxERcHGptfrOE3mmXZjc
77a91hKzYNUOHl1fiRgIMFfgR44YAO2d7hMUVHlfB4A20uYAIyOujPVL1Sp1
LBCGDHfxbUOuNiD3WginnELi05+QpRFlSakDc5/ZVDhBeA6F+qxXS+Rp7uhx
hhVnDvrpcYG0QL4k/ZiEZtiIPt/GANt5XKO3k3HtIuNU2hN7XDFzwG0tzZdd
Moyn5wmHydUtueor2vZw4fSTfhiGP1xtiKozrB9yJWhxkdgKOUy/JrRvPUzK
Y0GPAbB1t4dPXhrvqlDa1jT+s6g1v15sV169EpJVqM/Jt67yT16N/oIOicZM
DOHrEF8GNpNiWg83yVQJXjegfp8/ouOhed47OhBpzZcKHRHO5u8W/t+EKUFL
6b8HG/S1YCCV+I/ZfQprH3TokR5gPji3W/HluHWGJ7lxmpUz2IevDGN5ePgx
QjKpaC+aRrlyjiBBYjC+d2XumN5XLHaeDam/3r2Q5SzcfkzxOLULvvqGaViL
wS90EBkhecmIkBgPlYgRAauvv0MtKsNPx30K+/c/GA0r7ZravfjWxEcl5WWJ
glAhmHaYudXwNoOFH34M1EEFJ/D9tm+Df4xn0zraxyC9JMxG+6Vk1P+G2v86
FJqEMGq7W0aEij9EARJpZ3oMfstTJ2OgtqKwtv75ggMnyIHXvzxr9aHtilUy
BRgFer1AcWoxJ2yYAMuvPoDa2KqMjuVcHKYut+Z4CjtT4grFkjUzJNq+KnU4
IGYXHDT6wxAhFZoN4CBWmBU/eHKi65OkY9gr4grgSHhkSqNKgnzuddsaiFTO
iCp90GuG812Idq90kWX8jzuWiX+xEeFw1iMZRS+9MeQdfo1TuPfcSp+huZTh
G2Vupo0x8b4Nrx+d7pW3MfYdTjfyRDB6dez+mC3SEicpHceWkhpeNSQZ5HHb
6Up4M7Jv76leiwVA8dPVxEeMhe+do7vIzvJ3tVPEk91h1T5XdIDRQ4B34jVt
izGZ0E0CFKvTkFkQO+hXTKeCP6exJ9QS9ID0QHX9ssp6ZBS7AnB/3OmMI0GM
4z3yqcBZlHKBjJSEX3bOnpOcHTGGbpzgOTgCWx/PoV6O4j9VF1WkAa6c+IGn
clBy3M/sEg5kyA/KFWvrWFAR/xSSEo0T43V4KkAscouaOipYyB9d1JjME3BY
dHGuwJSTZqpF4CBN1HRlJvbvKH6cHmyIECV5DqQoDEAF8rE58WfEas150QRg
XbJlX6p0GFb6AIKmUZaV1y4YxOpg8ZZOjc0NpTaKKA4q+K2PdQb9bWWj/hl7
V4LChhKXb5RqGw7E7ZcWuHGEJEIBb9HW+5GAw5zXQj5cMt5Npiu2erONS34U
G+A4pjT32Pv73KisQsIEfoDUMKrbhT0gYhAkmUzk6z/SkYN9oSDi0CauHneN
DpudaHfchOs9gUCFqEbN/62K6NLwkkVBLHuYzax9G0a/DSMOgAiN+su9fTK2
aBOFAx5mKnzFOAhLLaeWwQ29DflzrfRemq3d2mx1ZCRWZletipPoKJw1qS6+
BxTJayurfn9eR3WahzEkkpGrBUtMJC1M/KGxx3EfB7DS4r/zM5AraTN2N7ww
SKNKwBP13M6pp/P4A2qAvkjQXs1rXkVKJC0b6nppsAqid8yypd9ZfTllBVSP
3OayqA8+VmNUxLLds5yUaPPB+lI7jmEwFrkHhcfa2qLnuKwAIB9dm/BvUCqC
QT+yYbqfTDJ2zqAmWwMidaAyt75Mu/o2DCUF4KBJp/OtXWT2USYETMASURg9
MUImt4LfgH5bn0f17+4rUdNoB7M3cA96xLA3R8WQ3+cJxQURPcgCIb8ghLSd
ggOg41Jlcq9+FPYcjiwaKlCS88yIKWNG4ivLzmMK0eGdPCvn4crUG4MzHIWL
/kypxTLzsIvVxNg0G7pp7N8k+gw2Wj9SNIE//uhn/GQCfsmUc5pFYClwvajQ
sDNJbtnvwFVbe25KT/Sg44NrqTXl5/OJqQuTEl3F/q/Cxvu7f268+T40gf8G
e6v3PG07v/2NkVaOWqcdd7EyYz/VCtvSaWGzWGRnwc2VBZ9F47c/AXQaMiZj
pFG3MIK7jO5PgtlpdAMCVynm8cAwB76pTpd2OaDgSs4oujBN7O1yz/FR/BLY
ezEBwsmHRgh1AMidEiz0+VkSeaas8Ooa2PyfOi1PimVVuojRoDe71nv4fXju
kmYObwfHAA+rYBtLMRmKSqkRn+celIw5tgN6vJoT6EOWjpkr0KkIinbPyD11
MXkq+pqFvdsXigZ+4cF2KmhPZSnZMT1R4Uzsh0qX4Y3QFPLv3zyvR8g9MKWv
MdlChbr7kZmqj+AIw5XE8Y6NY2tYh0nM6G4szy0Ahyy56H1wb9XiMUlcHkPO
WKtKPKhqboRD/M9CkEB56G9nK1amaV/4DLIn1mp/cURXa1R116uHsOy0NY2H
vsuBY+L5LrvwL6FLzfEDd9MtZ7BEijhvZUahkVDbENm5HzJugzf/+tgu4oNF
xFcoJe5fVEwiqpmmEjc51SCJxfKdBXTX/ZcHw9q+UB1Y/h5vBY+oXKuuAbV2
sM5e7B/evU7tkOmrItxsEDMI5Nos4V416tauzTz4VTh9y7xxLtw8Vc1bzIql
qJPdnaM2N3FvWrtw3m+LvSqjk0BtkmEt8DrtRpnUjBRdpP8LgGJYaxCR4U33
2ylkdtfsCvIKkI8exJVFurUbWOknRrMjgpo6XtmOF/magwyFZjxCwfk+1p4R
Yd7u6MnA5blfyLu8Sf7L6nCth5E+yGku2T3IePWRiyNU2mia7anmPPEmpxD/
uDTtfmW/quqk4YeOFnDHUKYwTxE++OIgiuxaDuCR0mVFxqZ6p9UUS+2/r15H
OtY4eUPHoygYeMXSAf/R3oZKfkfrLCIrDYOJpa8UJg2Nnj6XVrE2fGXvYUvB
dR5BawQZOZgiiiyPdXaKLrYSnLNQajFQ95GLD0xNOylQrgJx7Arqm2kwEFaf
ZJxiFBqsCWtepvKoGonLbNO6IpjMg0vg81ika3amKi6G+4g/7o5OaNSATNN4
tWTBuZp5ZnHgT+4Pt+Cg3Mta7VT7gVH1fUD8dL+m4d7cD8jo6aKVSQlC6UEL
XZR0fGGdtn5ju+fuZYrksegE8/vT41xK0Irr8B3OLgr6/1g0qQ5N0L2r3AgH
fdyrEp3BLuEqtMZL6zLWiJzd73F+wj8nXC4jmYhatyx91Ugs/cV1iG5YqP9Q
+bZBRZUwjJj9O265c2Se0Te8T4eU9V8cJMKmh7wsdadZeOuQ2BJRfppU33Lp
cYCHuLTAnQOPXWM9uVOJZ5HurgbVc+6VMIJoDgCsSFPuKynfQZ8FNg/OSlYB
7e3R43wsg/D1WTWJXZimxbeE4pw99Kiv0sZITRp+foSERaDQ7AbY2ZSgHp++
X2gJgd94hRv5Xm8JGnWagQnpZ7zOadvG50vPbYXcGhREnA7xemL4RMdDnFT7
E+Em7VMCba5h6DvzqTD8UDU993eC7dbPseoR1jK3B9B+eyCTwktGVuIYrgP9
yogiN1WgOLcidvgQhUQjsFab7vs6Cz47lWQMdSNF2AuNZIRdTNNwLaBxLek/
M8B7bV3WCJl46dgM34LRoj8zEl5gkC5rRIwFm6MVfDnNYl7F8/vM0zYxwH7H
fQqhR+vp5iGheQ1seyhlOF+4UNAtkVId8KQwJBNJ4tbquSp1ImRu2jW9cXRd
X8Rp3qK5E70ERDuVm6qOzdXfYqvGZi2cKI63pRV3VVz5joFha/qNSwecbpS4
OYd4tFoN+KksBMKFFMjFK8wzCteNVg76XT+MaXmat0B0gqzpQCHmW67zdWnA
cugo4iVx3qHMfNaXIFwgQ392+rKzPQSpxiFJmQnrBjRQw4tk9pjl9jozDwxL
W/ertDrlhTl0GFBKrgaCOxih5jKt5sz/eGbciD6ToVsMMqmODUEjHUGyr0ag
HFTK+3Jr5yWeYa3od/ZdUeCbLqUVJVy+X1IaA1j2GtyVeeX0wVEu72ZsdXrN
ULMgmTsa2fc1L4+vTtqvLlPHyKY13XD16qsRFrc9AZq7Y/GTE0+8v8iC2OiX
TfLI5yLmfY3RsZUgUKCX2sUCNM8U0f7njJQAzfGCx9G2HcoNweGb1k/XMHM3
Q5taWXEP9rE9aeFI4ydpYCr1ALypXB1CRAsqMdvcaM/GfVTPsZSxmhGcZsKR
Vcu9Iua+15xZh1EP3R2UwGtSD30+jvF/+5pC+Iak2dsGAbEmeo01ie7n0fak
d7qbBNIK+HyLrfuPNwxkwVKn7sLI9bbGBfcaaAxZ/LkpLvtmwr9pkRba6sv6
0XsyaVuemAwrAe/LSJ5WHbd8Ax4dVmV5WGA/Ol/nmtFZbw/hGAJPVqTz3OSn
w9hU/1S7yuNqNs+jCPWkYTABPDwP6ewFdJalxrUaBDjVH22Nx7rdM1znIdYw
nvRpLeztuRU8f+KTzGM4XH+MlhJO1WR82gGBwVsD4Obync1etioN/D55tUG2
x8asavLRyEkTuwdmlcykcR9ALXkh88sx/NEoof8sJ6m7Evh3gOCpdlTycpJM
OzEB8BsqSeY0qlDAX96LpPEUhhWN4JG8F3jPiIUrVmgD9cR3yuoHWf3jQ/n/
9lcLn7zfxjA7BvCB77C/qMgCKdpwnXK6OIBqMKWwjRNbTrS3ZxR7/9kZ3C8q
SHmygE00JsyI6gqstdMq05uCCV+KXN02UobWoXgl4lo3cUwJKAq9G5R7SrZ2
Zf/AAFpa7Ofyt00Q8QYaYNNojWL7U7WuH2hZoAHxmxiWPFNF7jPsk10UJbGP
EF5jrsuqMnA5D2fMKDty/Uw8drzp6I0xPT87aDldk7ZmRoPBjuL6FVg4YV4A
0sTJaVbf4oK6Yi6NwjRfkYGhxu9ar6IMadqbks1+mnFYY+0SWEyMTZNSHdgn
jlB0ieb7T+uwg8/djGhtyscQ/bcRzzrJ0iMn9XvLDsi1zfYiYPng86k+2Tvr
qp8CXH7pFXEVYoou4SeVCJTPbJhLnj6A9Z0BWyvy9ppFUjP+/d9D1MI/9c0U
+a5ZFDQt+RH+8xxZNjulwAUcxtJAiZ+RM4Z2/Z3nFyUiJTTuorVYeT1TsU96
5V6mORXcxn+YKY24+NKVL+RHVwNrh5KjZHoa5QAN41QA9TucCIC/luHbiW10
E7GGJK4ACsZogqtLrLZh7PDXfSnYH4mBkOqNS69buXY/S14gevt1dMxHFGit
Y1et3scKP7VssJ4PHK5wWINAjVXC0U50EP8NpqbWoQbvFarRBIokESoL27VN
hNNz7jVXYZmiDUo6WpRSGEHVZ54FD0y08/uRtznL6w0AQBDpbax1THLLTGHn
Bm5W8Htvxl8KzOlQ6bTIIIMOyG2kPZ88MM6qBnqc16LqhfWOOrcw+Ru+AECp
qK44Y9Udg+8JReTPHwNdCpOBzqAF6bgqUzajLdiw80nSSBuoGOgINxcEwelc
ABWg15J4S81OXEG3q2YshOe1TR9f8igUvX8nESKbUDtIQy3fJLAHPnV+BZYH
y9WpkYUJmuVsVOIzCd4HjHjwcBP9cgaW837U+F0Ml8wIX+f3VoYcfN5WYnAc
DkOON5d97Z7YAiulxe1eTLh3KLe9aukWSOgSz44d97fypqMUSubkyfgOlUaX
EjnlkRUsO+k18dJQQSjKXXH8obSdFPIAFl1r+nrydgAcGV9vVIq6ye7n/ntx
xFYnGlG3SfBJDq2rKCBWL526UmCgHFgBkWdfNpQDGJUjJ0MlcXCk4juKW4SE
tstcbnOGP/e5j20E5Tituj8VFNiq+NY0UtQ1Pl7iBnKT6f64MIhT5t6JI+XR
2nlCw/5Z7lv15iH5JCthpJ16TP1qBwXnnipLHeII+W0EgX6Kt1ikxeLtcxrz
+Ye4u8rXYT9UQ7VTqFuPCtbEwVoJ+rGrMpOmCMnXC81XPT5Rj87txxHMB0CV
6V7t+fNdQuCU9OIEpUiNBuKmFdjvxR+w0+2c3BiVhYGVg/K+UXdmhF+s9n08
YQ68CKYmKIFmPT0AktzJWu14taeWHemE0l0zAat28o4PvPbIA0v8WxdqtmvZ
qJ73meoUj6MGDV5oYQuO+jrKc5KnUDEMbgpA4u9HzkOmtKNT8wqZ+r8YVb2b
DLOvzCRhN3QQsL3lc70oAnpCVtUKu+xV+N6Q6kbqPjh/qub2FPwpoAz+aZDI
FRQAfZ35OiMAuziuJbsx1yJnrE/PV2t1sCsEdU8Lt+sF4rwz/2I3/oRtplPc
wTclOnAnlT6fAanflC70s2ybyrFqaoCea3L6nr2E39jmBsYAI1FaUF2/eKAQ
l51JetPYCnkvbUrB06CSapfR5gtIF9Tykw7yQ+FofxEh3iK0nfbE2L58AiWo
+JHHJNH8FbNKYcediU4IoTCYDAfUYREo54Q0NaxN5qZkjVQzHtmcSp9BYWMX
S2JnyQOFzjAz2Smii/tb04PhrI9PHqw4kS22/TYdmV8hpQDRXl1u45ZjVAVN
bEpBsjjbHDQCpqdjKYxlTsegO8r/O9gAMNsyKidVHtv5r/am/ZKz8maSBuW8
v056+YpNwFgQcnrUjEdqF0HEO/zwReSdGxnJd2ddkLq0VkrMWWO2/FJuxH/n
6REmTD5Xr+QTvP3QXwKJFH0smXvOBvcfOvE5JLJpqRfW6b7c8xU09ifA9SyE
hPVe9xaDkfzdTO+U8lhGtzx5AJ5Un+wP+he40H5WK/UTy2gldDxjSMxL58MA
mjjZ08nav8tkNvl7MuTYe1ypvbHGpNiMY/ykfVzYAlb/ts3z9aVb1WYPFtts
lKWwmymzscyccXs8iImJZ4AmpxupNKbnJo7jMHnHCUO/LyVXvxg0nDo/Wthd
f4eiTVwZsu/c0idK5ZJ+qgT0yBWaiwOW+2uX8GOj1EKftO5Ay49ltoyTpc1H
6ktITd2a0fo3TUWnd37qwHyMJlA2MLRQKiIJQu1AeVJJkFrEMPfoGQPxSgMB
F4VGJuHXM7ELm7tu0yaMrVxE8LAlpejfsdAggyrBf7bOPMPphFygKV8pEi3F
06mF2XEqxNgTWrPMYG5Q33tkx61/kI+8Zn2yJDysifYTJX/849GZTd4IuO5N
Pn36uufO+D0kY9iy+fLoI4QDPJqKzONw9cmVd3La7tpxOMgx1mGUbdRcwdRZ
5wYmGKs9f2HFznkpnR8hVUVXUwMp4bvJPr/R/eomlrOn2LKYAbAJBeH7uwep
bVszOrgKemgJOA+OMDch70XzvVe+19AgtZ8dllORf5HDlU7wP5DhmT+zI3+G
VwwyALLghBZWOAcFYh6Zgk1TMJqO6zZSf6bQLmD0SiNsXq0ex8cveGjP5mHy
ZoFY1Ju2uSgpaBQJNLVSt1+pIl/jdci5HaxSevBRT/u8/RUne0nU336rAwIi
5Z/2zWZuBLNv4P3LKMtB0UmJOlyEyPULIxwczIqFmGOqI4x4IssjHtBFMuyJ
g1SWWrQtLBxpXXY/FJzr6NuJhzrPnfFhWK4qzohj+kOkPoIlymIE91DvE3iV
zefFUthHOWAwMy3UkOepYEB2Yz93IGDLRViBfeIvUPlhAuHvyZRUBfoGIgUo
roRxnMr9T3d1/huSzMGgot9dKia3SXw9lh9MmAeKCQ3vjbOvhwgsPQa+OLFR
F1TZ6pfT3WIPvoNPxX472kTFHMT6MN/qZdZg/qP/GlIuP2pf5GXUF1dSqW7f
ueU4BhYzXetdA+Sy0z0bv1S9dNsBfaJb374m/Vhl2aEs9rRznjaigMM3HVge
yp7RxC8M+TcZb1y4tMnEEe0+XU8wjyHlO28cQ7ozSbHXCdCPIL/glC7/4JkL
UQIOJHr6dugbdvai8142KUAvCvCse7G5y5NIovsnRa3CO4zxjlufACD4Ty7X
KpNq4tLHQzlFY4jFTRQUIOdgmQee1cHO0w7ziFp5rbocbnWcOnHw8rmyke4m
4hltJuuLJk6bMbznTWPNha0LCk6MbY34yeLzrwodBuxXlkl6Blcvc4hhlGch
Jms8iIY61tUEiEZ6rLiHix9zxu5bN8wAIQooQpETHtL8YwhbmcGbWBumwHQU
kGHB1ZR/RY9yDngLDGMcqjyfWZQgG9oP7/UwJWetacuJBOHoFnf2r4Cr/ZNi
4DXPogQrGx0WbuIPm0QT6iLqeMuqFiBy32vXijrJTjlF1aKxZoI1TOTZnw+3
+la5csvD4xuc7joPKUQaj5W5lTmOJVhB0UBynw41bPzPcQ/1RcN4YXmq8JpE
Fx8PmLHmLKh+XEk67ncHEzgp9jfPyV0eA8ohT1mx9uiIIA3UCKP2hQpiLHcu
PB1nhBfr8QR8DgXH8VprOYfKiThxDLplRw1PUkCykNV2pOVZx9vXubePa5Yo
JnO+ygiI3NjMATZEkZwwwOBCiOems4P3NdmICmvRzVuQZFFNX20FTqtNYPAB
Tc3sivlFWc6EjGdy35dquMQdORpETI1l5otV/cjnSkUa/89oR73Yw5nIztsf
GZ+E2LRISOlU5VFYrwA64Cje3ISjlUKAkEA6d6cNKqOv9pbrlj+Y6yZiuaOb
4niqUVeBTnQJ3l9yxa0SsfKIGNN+1Ght7JejftosRmtnrtzhcxGDmEF2I77t
vrF2JZR2oHP7Dt55RgvOvq7MHThsMohBmK8JXZqrRjGju3zlq4wfJGgx85av
qd1HKnUAQp4e8V0tXzkc14n9UZsFRNxo1eMTsmvRwx/V87gezhmBQtSuoW6R
vmROWuEl3isYf0aG0JkLsYM5pXo4sWWDbzY8/C3laekgSUMLDoZBcpjRBIN5
utUyetk81Qw1O/JB0L0LKFRyM/ct401cNmqh4bJgJAUun0J+3MmzKScraTkv
2JXl0XcPvMHGumAqKZGiln1hnBo+8OmqB371mouYwvBbeZ9dwyurZHlrSmlB
3NUKFhDEGHYGrkuC2gvG2Uhvicp54XaybuKinDwX4yaMghBCNmAb6kyOCrp1
+caILHl+p1xjkalzyr3FLWIFaVsKVbVe7UitA8M7HIbae8CqEO8K52bFVp6k
a44oLmIBVj5zpuwY6z72q3dWHK3Iqr29zMJUeBcqJIAX0lbLbyjGrwG7F3Cy
077U9hgqF6fXPapDcVtw2kDi0+mv9kr8H+o5r1sImUAy4itFsYCOKKuXdYDR
MRlqMKE3EV5M8QFE4hiw4vFmwOpeSPL4LHd4IafgvaDya2whg7FvBQ7cvn82
e1YR1Ag1CyUnXPAbCRZMP7xc4NEW34qrHJLfcuryIWTLdWOjMmi5HeoME3B6
EuOsWyiMYvwjVe0J+lwHGFUxbX/6GAkafEvVQKQ94a68BgqnAEuX588CdFMI
UmJ4RPAhjN5xPe9ohXQfGtVGMaRARZGF22trbpA9YYrTnB15uiHqlJuBSn+N
J2OCC9YQ1Z7Mof+yWivZeHULOPQy+nKHKcTtnWfPS8gXYbkYDkChJhpicUtA
De73AOB/PFZJfsUExL8UXIj+yjHgp/FGvqt2EI1ZN8Ho+E48yav0YlUx767H
gI0ypJjepIa+egMHcsnmKwuwlJe5Z7MEvqqRd9A6Znr+rabv8/RmogUfYeHJ
aDq1krTxfJJTURKGPgXqaU8+QgEKoM8+JsdBpawai1d1+JbODkojhfG1rn9o
nxeyNQg2CknL1dR+eI2PHXY+rjgbgpn6J7E1utoocT76cCld4oKW+2C4fulX
R0mm3T0h2aDZYOuJDrclSGowtSTT/HTZoqiiMW2aZcqw7tNOVjDORrgV4dcw
6rH/WTVeh2jSm+h0SpDvtCOdT/lnCLYmBJEksfkXpPkvsRcWSpHE4AKI95pV
RwdiN+9PvVwNWmIlsljprxLLvt5DUkIm7b87nGjC++T8y9uMHAh9b9PN5yUk
HDnmas/GI1unk/1U/a+LwDDr5v6HwiCHJC0V3foanjfk8hXuagumHXp3+OEF
sszw2G98frciUUk4/3f8UE4kJJh/wfzRmGuFy+iOJV7G8hyTXHQFBAui09Ml
ssGl0oRyoEySOWJSF1fovFht9LDzgwaGFK3qVq4vLTL1fxaV/BXwqrR/J51g
scxNTsOpQIPU+3RuJP2FU5Hzd+OWOBKUhxLrhLORnhE3fg/+nGQrOBUkcQUq
KzGqpaALBcDJzlGXxICbrt0V6zlg/dpa6TiJvFOS/9qGYBCB7J2nu3xfG5S5
7JBwyFRYhVy0N3gmy7d0Xcskye79QvWqMSpaKmVW/9vaA8f9dgV3EZRtRwmz
kp+s7SePphUZ5DhO2hMUP8Yd7f5O6BOa8e/TjLytkVetsG0O5gM7pRH6MgIf
dTdlGadjmX39fsi3bFZ6qiFmxgS9Z/G8EdsmXjkqGgW+qXKAKpcAAMyg+mwP
2yfHh3P0FPCfz4JM0NCzwKpJc33RQbFPnOygegfiBZ6ywshJ5V9EKldwJ/MH
Gsv91rYR8rrjHk3HRhJEf2cV6PJxZFIXlZ1Y+UXOuIIBDIztytKBFarfM2qp
ba9/4GlezGepWkt5HN5nt3cWLIpSu6jyMh9b1w5A55/SMEjk8k44y/pbBDkr
BtrLJ0/QwQOGGbym2kq8XJOsR7WYBoCVQ40/d8uwpLLZobaxty5ocT4aQxos
3z6wYQnSTQMIOphRUwENYEjPFbRz9K9rBX6v39DXF1CIAwYtLqHn+In9Rhp8
g3de5ShzbiCUyjwdck//CEz/3Xdpeh4Ue7JhiGsrKhHyjPEA9HvenVnTr3MH
7Mk1Opc/vBvywDG5oVlwyp6DETSuRN6uaglHc2JnXplqBozrOi3Toikxb0o2
uvrBSy5NVMm+cYZF6Ct76p7tJR9lmT9mkEIrrI+Fd1VNsgbY2rGz7VlWlseJ
p6GngXQrOD6BvByN11aumdrnecADTNfMypQkGLKbkKGdHTBvJlyYZ3axmm+h
3T8QWxd+2X6uvxf1+LfPaV2Cw4e4cu4X4kKzS3LfQnlSXSSuHHaCQt4VmdkY
Svt0iw8TkgpAb0p2pOav3KqOrfAh9TEHYp8DpxwxZ+IKD3DlZwAg9jpPWcLY
5fEPLUGO9gHRi/u7LD0/k3GYPiTRtYVeq1sg8fQTHBhZ7LKCDvk9upnbX+Bo
QYgNVImnB0e4Sj6JXkEPkQFgQVbrAK1LgtCe36OqLQbM/r+r+UPWSRL/uPhM
OwW8pdF46T9pfxJjeReUscu065QSiQdcYxB9JBvjKCfrPH0MRDaF7lMGqVAT
oGiD0hsT+zWVEYGk611OUWxewTt/rYoJdiDQC1MKY1UV1+/8FGZQqwXcc+cr
4VeE3ABf0CkMMgrl5nTp+s2IUchJznLr89cAIXihtC+2i82H9cm7G+RmPs4Z
HeT8rm+g6L0K03MUByB93MFLn4dTMcPoPhAh+Yl91FChmyyff0ID12JY8jqU
7c5G1+9VDCqgnBltXHDeukY86NfmnpzRH2Byk8QZhNppjNNevjGjkS5fPOYZ
QJZt0L7/kg2nNGlslA5rtdJ5A6JCtif2ps6jgXuDip+HuCdMmwFbyXdiaBwl
RHmtigc0hjhlHVIfZb+uSoA5cRP9qhsNIeKen5vS+lPJEGaRmcbW8bWm2Ww3
C7XIoIe1nezbjoRocPbLKVr5WZzTL7Cla8goXLKlf+8IMw+ZK0FZSnj0hFEF
ZRk55EeoxPx4Gfsm4xWXsZ0lnkvVkxhv/3uIdSqQJFwbWPbrBeOkjGFuOQT9
67a0OKwr/yUOLBXMdh2sBJmRIL3VTJE/Y9gN6w3AJijK75NzfU2Szces9CLW
49BpKQf63OthqJJzPRD16Z9N8J1ckS+yvRYbvIZ/ksX4vx3f6AvVEVSNkvd1
YHanmyM33xVJNjy7QMbWjLTchXiXba8bLpKSF0pfv7IhvSTj1LsjCsJ2LgJR
kJVgFbOAgLt8MGchMS54xm6VuXdkzoNHu8IsITaKDseTaXXGv5brBYxfXyjn
t0mggwt6Rsm185/XyPoqGwnu8wp8clh9QDh2x7w/MfasTfw78i9EjDWTd8Zv
I4/RU/R9zP0cVmUKe6pkHMpjsi48UG+4xYv0O8DghcLAQe2xReFaD9/FT4lE
mFBZx92NGHKkRCjS7rFjIWglbRpJhjEvorMpgQxTHF/Vsh388GLuDrzqryTj
AhBSqhMT++RUE1XSfbKJQ7iRgSMnbWsalrxjf8nEFGB0Qmr2lhBadkpvqro6
LsZuGPzz9yzG1A8VYqnUGfdkrwVmcbV6IqydFWdxTcoXs6RnZrEv0Z8OYd2f
N9epTyegK1IXLXUbdNRcnfnKRgPjFwyO0NUY3+4kkqwDnx3nT/b9brxQfyyS
I3Lvj53KsJxxBY61vH5UB/p+hBfUnT1pREsnjZRT7XLgWY9LVpcJj/mNAU7n
mOxF1M4F1GvYX62fB5cCprwa1kCbR9eRtu3X0yhHAdyyztk7zC659O0FhWiS
G3sxX07BGUQ6/bWFxY8PT0qELrN2htOYAller9CvbJ3lu+zA7LyVhckCRvTv
NqX0PCA4LUulNVavX2f5N9Le3lwJ3WoTjmhpHgpxR+bQNW7zwfGxbu9PPsFS
UGWcqIQTaBIch5w0cBr58i73W1VyvIU95zkoj6fXhUe4du30hZU2M2oVd/vx
jfZ7e26s+304E4/P+uCKzud6Il7vFLTE2KIhNiIr4Fjz9rgHxn0Hdcoi1k4Q
uqbD5Ezna2VAf5RayKc7+y5TL7laX4chrZz4RSmpq9bP/s+MZHXsdv1uf2M8
rIcfQ6iYM21TLGC57P2lodneBiks+WcY4NLjR3ZnpoDPNbEiARbxM+hlXVR7
Mqq5u3uk9nNsbrTKHUV3oeEHiZVZ6LtbCrQf4rHju/hbIALEcO/rOZcG0yzV
PviDdpgd1fCczQ/FGGcNdxpcIyBROumal/yn0LlvcNqUsge1den9pSm5gkxF
K1GzYzigh+IXIr+cL27QjRiNatAKMyVZo4bfo0kPTp6BQu1ts9jt6Z+5EyaH
Nv8wmc5c1HWBxy3iVsTqo77W9l4uK+pyEDHXlXUIWwg2llIgCuYCBqdV7E+r
/8YONzOq1T2LrtO5pr3biYsvoOb9iU4+kG4IxoJ8O3aTZfM8WpbQArxD0u+A
juiWmADRFFXtq6U2bw09FRajjjKDojsPiXkLaKVP4VIqwWXuhfS+utfb4lL1
6y/hnhn7VtfOq2OeVFfyvyGO+f66eon+QAx6z4XmIanAQLGzolHc1ns9Zrin
asCFycQ+a2i/k4hB0ZMsYTnur2howLr0AsKdEtpJtATrf50nYcw5KW+00/Cp
zWj9a3Oye5k8bnas7tAby75vPm4cYgLv2gdZLwTo/6D2CLK4mJJtQOiHZnoj
AZCJiBfPbjlziHARpwe2Bpn5ayA4ASptVdrb2vUrWoGM65MIOUsRL8+xZLOS
XFz2/zG32EgqVJCan8HDLC39dJ3KeTDC3XWf0U7iED1mdqYRqtV3+y125tRU
5tZeNPyBvl8uJ0+h62TssaOAErBV/KFTQxOx3aLZiMFgf59I7z33VNZ1tYdi
23JsM+af3DqRFp5wJVNNEJ4tiTtC/znzo0iMWzPEMprtMvR5Y6Acnj7jwuVB
Vny8kSJsNXJFTnWk+3ujxKHtdG7ZEaWBVD7jlPfiIU2r2pBeXm8lMtq/bbXm
QXl5nks8uUZ0xkRLYAaWJ387vZsNFvCLL3wCJzSvLqX/bFCWJbA8CeGSeFeE
a0Xs+47oKVPoi4iS3c/nXe0Xp+ftMlrPM2d6wwGfJ4lQY6hgRetckyPFJlpG
Hmto9oagxNN4E6TDHmwYIe21lUlMTLq63xoR0B9qIZJKahsLqRK1W297aGJc
64EZCNQtUhS+BoqpPXQqZlESdtfm2ESyFpSsyKQgAvTSXofrADla+RYBKzEO
FlSAC28r0h7ksPgdBkQmNtTUwDysHIQYegKMFC/I+6Oh+vtFNlBZJCOQtrRz
sNowXMB5p89DTTQJFzhpsXZy6f18/8Ffvi6ZP87AvUErDkWRQSBTCPXnyDpL
kohDgM4T3X+SdMGCTQFGGMywhneGCDhjzLxMubHjW3UHh7uTAnCE1UVk1utt
AbOcQxnlN6dzB/LzcAQ/aeeiikEkRPhe3giDD6iTRC+Ev+95UtEhAAxAnd4o
m17CpkDQVbb7LDTMnRKbHLeshgL/uPXUz9+Vo9bKtYOTutxH40MZXV1CSXPA
8ttHy/kkETX73kom0dFoEU8h7J2slAkg+j4aJR1I2PaQ/Ry9EaI/yEEU67hv
Mc6tU23prU/2IgWVKCBcgb/hKt1ks2yrFVVb89q5qSzZjKHyT1yeOYgaFRNT
iQmHEYO/AnfB6zY7NWI7lp4vdV/gaqPgmJZVZrEmBNcTl49G90BJTDm6gDyt
zMoCwnPWPecI8wHXdG9FP8nHvRwvIPl4PKAPlzcEoE0AL7uw6xJfKCC3Kz+V
BtGhJ7Tiw8FWNqFn6LZC7RLku+OuBHjL9HesncgEc4TO9sPE812zXD7yOud5
ZxSXE2u5PfB5Xp25OZLDhEfdfxQLXRuFhGR/sTrNzxpX2exSIodTxeEtMkjb
bi8DJ1pOX+mxG83ivSAKOCj5eWKppxXNYepmLhHLkwwDsVXVQYiH795vvdRH
nvRW+Lau+LUEVuXcKOO2e5hB9hQv135SNcH8x5BRLU+keskHbxCqWrGCkMB+
y1lSVhc/o/Vrw6/FtsPa9b+VGeTsqXSY0RqMfXHv5D7BFRPOfBdeOoIKXWR8
q/YFfpgRnAvgFdmz0nBGE0HgWTPxIVko2ZiXbzUJkCCUsK20VcpCdcFAvfRo
NWw8JPNsZnsrftLAuZAP/Y8KeC+vLuZM8FS84UMMou21aC6EpEypMaOqUZXG
8igK+XKeUZpLzO5t1v/hXooBGoHHNmA7qzE6KiNUPCsRMcKTFznU393rNJHL
UJ6O5IsTEJwZkAt1lm+IDdH/wJR+F8n+awq/meRz7maCqy3cNcaDFKBhoOXn
upfSSiaOtJNrzJ3Tvy+uWhATYM2yzIk06dpDzuNSbqzk/cdMnqu2Paw9Pm8M
sMkGqy48do4wT4pYm4BCl6EZWMlGhu/dVu2wht72KIiv4N7Ywv4eVQK4AqGS
cnaZ2tmDpYQJ5qaCOuG+0CI/o7XosbVCAyGX/5uYwL6AD2lQWaVA3iwKfZrf
xblzAYff/y/Khsk92EJwl9qYJXWUjG6fYEG5e/5IsvQDjLApYJacAbTXOvlz
47LjqdGAtGlMCrKm+a/p1r1Lh616cMePGjVp6VIj0T4qy6rfFQbosNtQ7ARo
s/vdJ/zNirxMRFPac11/LEAIKmP30s7BlLr53e/Z6WML0DwEN3j/3hrHxzn+
aMQ9ah/+M0+RsWm7lgF4JXNPa1/Oa2KKSnm7Q3SQwhgh8j6eimHDcQK4wNFc
JPMhic9YuhrsN9cA3VThELr3XBpNgre3ggR2O6lOTG1MFd8pukII8H1cSyLh
/EG3Hm6k7pRqkzZnIA/UVoWq8PQ/uLKAp04uBwsgPnCVcvgysF0oa/Ir1JUb
NJfBwxT5lAyVKiBNzosI8gjK+L5FLhdwABB8vD7JixgtsLL8aSlcFMq7G8/S
qC6HE3FmPBWKmQU47qniDWgECy5KB0Zwqdfn7xaiojH6V6k0yQbZUJLb2vrd
F+HcnWMIcY2oZWepg74tE4uaDjmqkwtjDIfA/eEaG1FGbyfVBqg/STmbnWTe
xn5RDZ0hbDSPgo1ARaytvtHUkXlsl4Y3g2gr1xSCzkPubLhks3xSg+muvNTb
fYvxjTPtE+YuNMvQzcYsWHEaPycO69dzmQwMOidLhPgqmbaXsp2GrB1zOPxL
CxFU7leOMG3rR+THqG+NnH283kM2X/yu+aH9bt9muNbCJnVtPcrm3KIXWkfR
e4ueWF/ceUjyAS2xqYRlByFnkvXhcx8HgIi0SrkkZeBZOE2KExN8iy7bXjOW
oC0AUDmWNd3iUYrlneBLcNLjFdWhVEM6U0GQrTJP/NOjj64rxrzL4Q8GmmGB
KfQZNI+OPtxUoYGGWW4G52nuzjUrJM62RiMONg+a4rCxVb1H80OYTF9xLHvQ
T6x+yGF3BOiTFdC2IDOUIH9FxZkoDypI+xuKifdTuCaC/dnXHDOlvr5oLUdw
CnotcBTp8mV9hQ7Gm4+G9CiIXrGeL0C4aXK6zKklyTPD9u8MxFiOM3zzQAhd
bYT29zPm5InW45WCZv6FshHlF21LPTxGjOCN7YdyPqZi7EBWCu03E5m2Rnt0
EYo6HC/B9XeENprAlRqlgzWfw9TwZDbd29ZMiQ8lhn8blCJ+ACyJJlvFd+zM
WIDLa0BJ9NvgNhLyhDxMRWY14c0T+8MI9evm+Lnq8xV6DezNqxXG/KCOIKki
qkcdmV819x2fxWoicsyj+nDjYQw09vATYj5E7ja/mmz1aZHrhPm2ytkotqhD
c2uoflT0EsZ66bKZOmxk376nRyLFf8KPT9/+N7y5mFxzvEFHMCj5C1rnjGgh
gqfYaxX8qCnr5qWCwYJKnjdXk2SfLONMkBrSlsK4ZO66NclWg7st4tLCsEW9
RRBw7j66n09MGFu6sc4QWWdjhsMTeJLWg8gSpm9rx8xElGPg3gaRNN+5tpUE
W/smLQUuWV0ysPgNfb9HMUtOlLMH0d5FxFOmf+nQwWmO7S1VmTxImjrPlLcf
CO7OgNoTOobx196xgbsTl66z4l/5i5ih/qEdVz9RZjQC41A2NchRo1mU8T/0
odGvB+lhnzH0j3UntaHBIqwJSmbwB+cO8viGJpen+N4i4W1TiRH3Pidkq9ZC
7oaLF5ClVdTCEgLXEZHWmESLl5afzGRjjR9Qi6hh2ckMpEOgA4gVXdvUJ0JM
ZLsmUwablwlPXVZc3ttVv4DZZIjn2nWoBFVyN2RJOn4rEeV1NY/gGb/8ts+e
buXjb4rLFYmdrP2cWcw62WxsaMHhKaNdMD0cYmXr+yV7fAP63gPcAtcxRP40
/LmAgN6sQH1G+8XwtSi80fMa9Tm29S0OZljaSOqlmslAl0uNROYgPfrBwrOn
yEiJtRCVFC3DcyUZjO4JECBW1e5QqN6+01EA4esjH3didvaeQw/TIUy/DSHm
HZ6OpgBnxbGNZim6uaB0TDVl3bjl3G9s4JHejJUI46daqW1axXKrZeSAfa9y
H8NeF5mFyioXXBemRh+MDoVyi6ZJ2fQfDLa+ghLVWkryxXZrXbiPAF6rsROj
rd/lqXbt7PHa6Wi4eSncMol4yGGChvd27rp1mXwDd2mW26yNUqDCSnc0VfS/
MwFEMmWMAKgMDoNDje1d69BAOUi7wpeyh4cXOUAE2mxgbDyzhLgWjgNtBgOu
FZ0YQ6tpZkmKsZ/qdKdQ4hNdpqcj0Xur5mnrZsbp7p6Ic7iQZ64rrnFLksPu
8LxNluIzr0Z3ZWDupyhS0hY63+JCLCEJv86x5ITwWqVuQ2VXc6EWM/SWEhPB
gXP9tg35dQlIOBRecBZQRNv9hN+hOAZfA6YaHtwV7HKEdq/sDCDzDU6uUcls
r2wiA18EahL5

`pragma protect end_protected
