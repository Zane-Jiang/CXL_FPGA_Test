// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
G9zTHCJiTvg8d1nga8U18QRlWsmYPl99Y6z5Zfy1T9waWJu2k2ggceqM350k3Hs7I1cjPd55z6tr
j0cc5LZ/6rQPJtnfcu0XoPZilYe2IWMWlk/UG/8+BHK1Ch8k6tb02MkEjDvP96LQNRQ9Bxk272eV
rH2D8Fkn3va5bOlUqPu/k3sDD6JVNuqrbh89LbWsTwmPHfnddKbusjytu1HaGJgAopjjMPH2Hl09
bxfbmILU48D8+ZCbRRquO+IBL8v2NswLcN6xQZZCh0XJ8B+GtN8tT2BoCHbAvpIqqFXXEkvkgiWG
hYSGlGZevKXk1Sk+lWZTO3drECsZQCVs0S2kkQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
+YhzF9gP9ag5L6HKKwE73QSF2wwYFjYnwGVf/eJgyNZ3s6HEr9vITfwlazWNJusHYS9X06xQCglU
L45UzxAey9JPh9DVV7VWcw6en69BQ7Cxewmsm1DMVfrW9agvGaX4Vazn0LD1zn0q8tr8STdNpVri
EF0iYyEZ2qSjXn5vz/dyhf6lUo0L2rWah9JOPD+SBkmNPqA+m5GEQBPjGk4gTC8XXEIFXxKmVukD
NGSM1gRYEAOqcFQmxsL6EIFQaSlC+iIiJXF0ROsdL6Iwpe3xbieino30FqZ8ab/9iB2qtvI3Dt1p
Gp7x+cpezJNvrZ0VdJUIqVh+3QshfGQL2A3oi8jEzNd+WHgBm3wFnvQ+T/bljIsJWh7foGUIvyo0
W9dzUJNukhRFo/xYQb8KgMPT5vPwU1cjOm4G1HNp1UDyB1Wz112D5LsgKfbXRjnk2Ctk9mYBtoGa
QGEFxloNaGu+AyO56jDv0lJejOAg8Zf4NwIJEPz1RyfQDxM0APUZqdUQdiz+UBm+moawMa27Gfi4
olZH+MNSNqm8wPVfHJc34io6sZODQKa2WIAXdhN9NKkdtrzAESja3OVEcB+OTN1LrWhHNNLug/OD
qkO56pwtYxJ1/X+a48YE8IjTRwUwqUApSobduas/RuYydl9k4PCLOPQG6tH9dAZiCQZrG+6nWA5U
vLEZ/S3Vna9GzKkpaJ0OuSaEWWus+mva+NGsijmgybqki+3o/NDTCckHjJacKps1+vwdRpYa3RIq
wdqMjFhMdcvGDVboCILa1SjPvodzUmyqRCebCMb9BQD+9SSrmGykMLy0FeOUaWjfr3YGZj8Qb5W4
CdKRSgKkFNfIbEMn4iixqsSzmOyLJp+bJ5XoQHlrXfrKqfXpmmQQ1JJbwHd4JUbN1MeuiMasMV9o
zmLB8M/sn8WOviUKbcdePjaoXqDqoObuxGsV+VFSW3ALZxU3u1pRkK7//1D9UxYMwpAY9AmGJbT4
JrcSbI3WDAhmOZjZuM/veYFwnJB63keAaPGggGDVx7KgpYpzywjIjD3ffwlsKEVdQkpXNvbyOYVa
S1phUXIukTancAOJZQAIsogGh3KQ9f0kGVkk/GMGVG9c6HYTQ3ctltJPUu0MDFHbbv/t2Ag4SaRo
/Z87TfLEnC3jwNXj35bl/ohOVKQ1Z2ZfgvMCtcV2stCDsyCK+aSA5eMQwyX0bJiFDCeqMitdZ+z3
gEBk/2HmeI5E5G9c6YJ9G2xljsp4jnFqQbPsLH20QlJGJSTLh1YHoK2vSqqfIf8EaNBTi32odRKj
AFqRLOqGYXEzXiObVibIPkAyI8hjp3uBHYShNnjd4pGO06647kWE2d3faTMdX8OwNNum5E/UnCyM
TmNpWu20LaOeIxem/jieWsPyluV09qXBGuUtJzdSyO8RTMJw01n9rOE50AwzZzyOpwMlYQSJc02Q
D2JNzZUFukOmp0wc1ppktSkKBJD5muIWLV++cKjX2BX/BlDcivzb7JxZj5KsNsTs3FCgaybC8KZo
9a8SHiw8EDEqwKz8JPTrY9q1zp6Y5L9+SqJRHg7lzP8FGvMrwoHn+2xhoqpoCfZkibiinxsL1Ceh
B+lVqijD5aKbK03k1hzQID/uLfnh6ZSl78qexldaz0JzcPvFT9JZRBxgvUzzokWwa8AiUKEG2GSI
4lht/h2eKU/f4R4VJx1cUWyO4Uca8z133P5E3NQ7ZX4SkYv/EpVPfmcZC+YKLG4No6qTsr8EDMtT
lXHTMMj8pg1nFun2hAHkNhnJL6YmbBUwga9jlxg81rueASKB3e4nTTBK70K14I9B+U7M0aeR3E5u
M5aS8yeLt329+lHN1a2+F+5m8JaKIUDwQ9bNYQ1Z4mSfIjnw/fM61rmO8TKtzXPDzV6hrFpjxt87
MqZBniHVW8Ve+yYHNrpYCBF/03N2pT+UqwDv4SrL5IYCWYZ5hdmHGQELrS22xtvczPSF+T93blWu
zTRaxFFYYVUcnOV4W3Z3rXSf1nc3T+afcnIHK2Ltm80D/2jHdByg4mWARgZmzkiN0P0iItDn0tyT
Zbhkge2O4MyZEEgXlNZvq/CiTacc6Rv9ob7Cs/bGx/GzbJgwYJ1YpA2xsQ5XzjKHEcBdN70JAeMp
SQR934BvroF331SiFmqUFu2jjMreOoXyFLbgaR7mq8CAFqkMkcY4pM6ka3prwgrTPPUh7oIoiOpE
2kYnRKErR086hc2LNbUY8lghdmNyo3l9FGLyIrluHZUDdxqKQ6YDbY5Wpyzal8Q+KwGMHils4tNA
ZTiq1yIZqmmLyxOXdR0WSSEWX6LvHGd/OqP+kJ/pFEXGf1yk8JQW3oiFfw2ht4JFImwJR1msPosD
qZ/p9MiNQ6LF66tEbkA1cNE4BPPsZWdYQ/AApHVFdKXqiYq77f/XthO69LAGuCM2n1A4kEbJh3UZ
gLypCZpolwtC0v8NlDNYoFRebQbEb4KJ+gT3Qreb9GZmPYWHtVtBWIOc+BFq0GFBHcK2xj+vEYmr
PxRkH2Y4ElKXJu3kO43PmIi9NXr4sCbWpJ4Mo3bzYpUSKhrtwkamV+vJqnuYhMu0WOqo2UWdf/Hy
UWU28tmxBwqgqXb4a9CNGuKjYagPM6FXd7ktMrXV8B/3ZWb6AnvaLlkNgMefu0/m1NMHSvT1HH5Z
hHwP3zVW+1ACi/7FBet2IgReURyM2mVxild10ofsL61zBDdWtB6updlX1D6IA+Zx5U/8PTXfiuJE
rzHdHRU3PkkEs0y6u9i8yGvWkkXHl1LSDOYhBJ6PSfLfuzwyAdRAtbcWuxlfyqXaJ45rX8IVEF2n
wWWily4wiulK4MXO8PRMcHwxIMOAIoSIc0LSzu9AY3PeOjBOF3x+3WRH+oPakQaGC0pwTlNffkg7
iFd+c/a+X5o6egV/1RH+GvLnz26VLOsgU1SdeePCIso+rd6acGKkV37lthC7bWp78ufiXZ63ybpp
VYannVaa+LcWHVikTXlECVTJqYbCy9x4KdtATHfXsNXDCRZhSgzB8xR4nCjWDm47pLE8cD9Nlg3I
6HuVrea0f7XyfwYJ9GZVo0tlTOgyNqIGclRzEoDzf47W8rkaLApyN7CPzVgTtPK6gLkgdcGetbC0
EVMpY7uJyjOCUwNdAyRzqaqnu88fy41pxq6N+p9rJi1eA5L5aYCXL2zlVq+6GrT3YU7Eaj3J/lIX
UBlYam8HXOJOnb6VDY3jGK1k0FW9znf/lCuXmRk37Jq9yqER7FHmSpDLWzafEtxE6uZZK8A8ILWj
ZmtKEii2oOcYw2X/f6uw8Pe5hRE5QV2MfpWuFcPfu6c845dbJIjPNkR2U3lZ8RoZMBtKPCh7aIsc
K++2sY4FFfBSl9MyRehV9KmFTHnSLeYVW3gZLRexciDUzCW3nb033yV0hriDDrwf1CqU0n+hiOLK
rJPIBsBNE94lBQ9OJNArCYPHtyZu/YAEY8QAxHjRGRDjG7dbAXoxIDAowhNH+nhjrm5EnlIuq0Dd
/mIx4ATq8GiPskV8osUxtxwuuzazffiji3kc/m/J1kASShHJYuEGR9EhBFUi6Gt6u4mPtyixDN0T
CbQrXWFmTenWFn86Pal+ASnylu9CmxBm9D87AK7/GsJ3/cmxP/rlmhzpXJPjvPkIFgOyb4wq2A4R
DG3xajQ6oiXiXnv5TXVbAYA9qFPfDhshkeTrL2jDcx2Jqr9I0Ek3OEDyJrMyrRJlg4AfYLDUWJTX
+gTJhcR22JGPTRiqa3DSWhNol+K0e03MId3ikXQo2RwtQ+03Mwgkn8+jUDAdLhMqrRaYsYlaKTfC
wYXmhb6dkXlgRa/1Z4ihEmBcQsMQhxNe8QIipYG2MIUAJZ3aihnD0PzagvyaSZ5YMJ4YrqUcXQ/e
QzPsY/Y+JJ18PkqxXsQa47oYFrUEUBV08Vqtq0yL2VCrm/2XyFpmql6vdVjFDLBz63KBXC79o7Xl
epzzswDCJDnJTIBuWEORzyXOulrVNKbpW9uiUUfxzjhKVXgrhxlcht+UvZLox6zNFMasRIYK2sRo
2+2/lt3NeL9NleDb1PibRhbIbwYq5EZkt41rC/3uoUZ4qlR7NuA4Ly+fffpEF0SZiSNLEp12uvtu
u7dEoTsE5UVJAfdqgeETXR1rb0pgDhei6GZBFlwJoZ2itewAE12iA1oxJD8ci9Fk2IsZj8KNm8Tq
xIbKjSZajLtz0FidnhxlJLVaLluEAtO+N30mYGPRWZcKrtgaYudA+8dDWkEYwSvX2+XBqPmYSRni
01SbA3uND1d1b6MVMiEUs/WAcc4TOPInQTIEQ1HvP8FwCgZJdc7lBk/Em78daq6lbfCXVKHQV53X
iqEbwdjbeTVkYQM3Sp3qmCjf2AgEIEyElNDEw/hGy/YPFNmxrCc7n04mjx7SwProbo8S53+VKASN
MjHy2s4O3S42u6sb/qrCFdlV948hVvKnKWrKxMUSWZGZyM6C7TPtGO+Akr1tkeNVV6rkN6ZvSjPk
+40M2JyF+Aolnm84NwymOkmR6M24KUj47lBHmtXgPgegcF+8iX4mtu76wKvbQ8RbC6V5zdj05Lma
OT0Vi8k0qY7w4MEx6jrW6MDERPoQ+VbPlPw6VIRd8cgw9lq+yY6r22RnDVXVj59ZOqlpiFxj0t0m
mp8HJ5CigAla1zVOAlJcXN+p7e27yOboIgCchmztZARLty17dhS/m1kvYKVFfWeQt7BE/fE66JVn
GBSQG1iBz5rNWhLsaCTfP0UT5MzGRoVJBH/96tljCg7DAgh3fO39qMiCrwfwxfYsTgU2Sq5A9qUD
e5h4H0P98OU+QCiUFkrRhU8ynm9ROGO8er1UAEj23zf7HLZ+W/SEceg0C0uTegDTsxxzCmxMO+42
1XxAottMGPYZqpcd5Z92bLeUnKQWVbHyB2F31heAUTIs52SHfpBJ2xihitnJgeih0Onltj4qK4tF
hoe/+M44oM8eBof148E8hmN8LYrWLW4BecrdWtb0ihtDvnXI+f4iPOJNDRma5rIknlCs4khu6Ies
oHrre672NVNqIY6Stn5jTU9yXzIf6e2nB02YlaXjZtUopYiUITffCeHmpL85pAALSPlwVmceD3U7
oWJIi61f/Wx3cn6SdcJnVJP/cYIaq2jFqxma1VGKUmWXHgsxRTEC4ItsJSweMxPMbtOl3yWjyoGa
nfEYoO50lnnrLsZLJaVPyyOYxjeTBOScfQuEa/cfHN+F4jqwUAj+m1uT0hEbqyoW6jAlDEr7xSSk
mlQd++LWzYmSoAqXBaOEDtOZPJByWrLzzNPU8r110mXer2Ir7Y2adLaSr4rN0Wu+VhlvTjMGFOOy
zDagV7m48BwUla3dsJgtLDPfHR5eWpzV6lnv7j3xYLQlr3ESpybHRtbs6Q7bkSassS7Y6FYQ7AVG
criGct8ORhC7LR4nh+Wd1R6rBt5oT+6Xc+H06TUF0U8fePKb2xINufCENySlHbsrpyaFSkPk1JPR
R8tEHRQuM96QZqyufdNQC8cAQD1aIQOvj9CARab5i3i6GrK7EsqdNINT1VNXtpxlojmJ6UKuUlqN
O8fsxGY7noKITP7msTYj62dV94t2Jrtb6LkmhCzfFXUfbuztrr55eKZstRwnYJDSh4UyCms/jgwF
54gs9blXifAS96ngYyv4nnXTlo+K9EKO4Irplqe8N4LWHqCEfLE5WpIZl3zZCD8xHSzGGboZttrI
DowKs+Mc8BCwFRpnFKci+xRmdRQn2gAE8yb+8dA/mJ++DheEg8qAgg/ifJf0xk4z/KSHGlfPZ7LJ
F5DOvzBoW8wK1Fce8zlvHHmFbtaphMKcyL1AxLNjJW0sGLMxw90BfOQglxnc12uLPICwpD1ecpuz
gioOnEMWhw+8/JrV3A80HhgekxO4z5Q7HdvGCq2owzgnqbQkh+tc9R/A49F6g9LRtWkh/u4OPf8v
PJ8dsV5E76vpgoaGfgfny+wFjec1iJNg8iB6sHBAnfBQc3+V/IRQ5RS5TkJv04l1YSUAXfevzJYC
BJPkRMXTyp/8qdhKphVBk58NJJlrI7ELjYYD/+MnVzVOYyvxS8UJVqI4yXfyTfU+Chpkg7saNRBx
W+rij/gaYjWcp3veHcpdrHGIcqbPzrHTduyFficrhlOx3D3YSyoHclPOEo2rvUhaLSwabpkfrceD
i7s+5L+wYQm/tLBN9Ts4NyghtBolh+TGP8eIm7oah/tuvCRjzMtuJyE+B0u82qoM6BIyjNBWupcu
TPIpLrbBuFnDmYA0J3iFxjyajvIoj5EeMUuYA2dea/phJq1m8tBlfxRJBqPb4+wK0op9T1BDgaCi
PX0dJj0qznRN+wTQ485KulzUIVC+CpCfTNXN9T1K3atpWItOLf6cVczgQV9iRHbh8nPE9u8CxL7P
UP4bYg+8EoPfBpD7bFsCg8EEe7oiSyQyhnBAqkW4CWVylUnF0iASPfGs015tiY8D87oJEbhE+PIB
BTsSjLIxDFen/5mTs8sp3K/2+oJ9tbHTABfxAmiTcM463BfB9kZhsGpywRGXUR6VsIjDi/COpwYX
qn4quv3RnyzT+9wyvbboFYDMCLtVm60y7LtDuVbPJAXLGPzrTCZ0yBgUSNZDV3eUQtcJZca7T8nh
sCekHXk9VfcNZSQkpZIA69MPFwLeODN3AODmG1n/F0RNQ+kNTHWsiCS6FwSoYQIYdcEPExAAU3ms
PM6cDCvgmtyvHilHf8lkaZPJCeAoU007w9fh+cfvkQTvqhCIkXugdtaIXaa1kUsTSBbkAe0QHhc6
bXMP+w9HHP2JlITb7Zl7/3b6wLIOnZtZ949VTuKtWiWz1DFr1Kem2AGnXhLtfA3yioSo8QCQ4Db3
oPxs/ZhpOhXJFUSMcGqBqU6/CZ30UL5nLGAUZp+rf97npSlEEswSoha+sXXJQNp1xOs7xaW/qM4i
nCNo7qSRKaxr1HniFMXsZ8/cVONp39Z176teOOidegE3mvsSXffAayhEUNFI8PIQ8Rx4ZpBM2gKQ
1sLHT6x/gT9SB4ycVNykt7X7lwuW1ABURIblz35Xi3O29KRUcGOEWnWFxaxK4nTgpKpzGVajngZs
+YSospB+rRLDAj2goG/mlsdJAO3PK7JYw16GUKg3r4hNQVDyP3vkpDKApsAOZ2FCBg2gj0XKaDFG
Gt/bqI0MXLGzR35Wl36jcfnL8/BlK1wgs7Pytp8u7ripsgEwNgQ5A8ymEjK7GXSlo9p2NDxbdF1i
B2mQTFrGicvVj7cVfOrhgdelpH69oLvo4IuLddzXkrD8GyZwXbC7zVPqKDxOcJ5Ag8v90/Wzne3K
8kxtqzY2tXJnLwlnKG6pTXj9UDMP0LMpBy5ilAsNaVG25MR1/L5FWf6l5ERvn7VTOpilhnzZo8XX
0pWE6MY4oc7GAhiVVJxlqtTh9RiulBT2tqst+FD4q81a6DIFJyGpen83sEvRx3QBlLoNocbycJQA
MRvCMn2KMlZuLtu+fg4TkEVPTEGyZyHPIyza/bQwf1SJPljTr/ZNTQk1/mUk6k/OyWMOpYf5wPDG
9IxQgLUYUWDfV1xl1T/h7omLqPUp1A/+ZMakZNur1CbEpl8gn3xK3vaqwTHjlzEJz9xbuj0P3ZkB
hsAl0KLCvBW3aVpGxs7ArKKF8F17se/TwA7KB6uQ1qYudm6PoRL3SBU5h7fEn/fU3LBV2Xbnfr9F
xyjWDBtkUbD5rnHa1ZAM+rhDT9b91Uw30PzOExYcw/zazRcFf9dTnT00snAQhXDym3RwkY1C4uel
fzmoA6oyo4MU/ywHrS22TMkqyTyQz6LmbP53E9VAJ01I0uW9Day2m3GAtg7/OK5MJa7dTgubbKo2
NgHSmvhl2yS/MvKpBJQZ8nCkpODpqGMsg6ZqFYNSCE7U/3XxMLluwsutk5LpgcJEJThU0Six+cw2
Owor5CmO3jWPaodxHQ0b7vstkm7bIomqFhiDNaMV5TN/+XmAtcuHhVBci+He+ZZaGX4oe7Qsudyh
EbUANTfm9df0Fn7fKXXPI4N0Owx5SBwmng5zwzR86mP/81wsOjEgmzITxnJVDf/olpZao0txMQKO
WeN+Twhdu/cXkpcIFbMJx3osTjq5wGWfORlUWZ1ZqeFYCrSU736ZMowGGZsC+Rn3jywkS3s8GB+D
+p+6qeKK5H0KK3XYJ+fA5aW5s/UqHZA/qozxkUynuYTLVKNlx6mao7OXd6Sjk7qTFaQI+p0WRh0q
63AVIrSSPBlE+0J4UBpRBIxB8Q6r0PcKYn9lduaNr5flB/+3bHEXfq2+rvWm+HY97godEVLAelgk
odG1lCGmCiz148uq4+UwLrZvFjFkiwRXTottW4xMiSn3QSRUQlIqiU95g0apM8pnyCKjZMnS4mTl
Ow2/a/hqv2TaZ/jqZEZEJR3fqPpfyplPWWbc0u+95WPa70SNS4tbJSFiEXQOxlK0M4zCvjLHjJBC
vvQ21GGurDVH02ZZ2oDiAe34VsM7wY3/H+ndmjuusuq3My/n5pWCR0dI4g9slPzvYhccEEsLRemT
dkhXuwJH9AGC2Yfyk8oAvthWSGAqKv0gWOGInOUed2Byu55CGl1xZkXiuJ75Ed1XdMqrS9/eNkK6
QU9ZvtGPQ5FYbepRdc6Oy5UaNEoSnIMlncG4Zu/VBdsVSc7ypwCELjTHHGFKCNrrZdQNKCpNjoHD
4hVEKvJW/KCJiKlICD25IuH5PofWHMYLqspZ63WX+HhASlWpzEJrYOLoLmPbu3ITVeVA1y6DvBwb
asg+b8TV+T+g5g6WCzY6hIm6XE7CsUyw+Qz73rTjad9j7fp6dxieMzMBHGuxIbt675HtOlrBrehG
/ceDd4MSeUDqbhxfJm6AJWPvAZqy/+bk0foFuJHFCWc3cyKfqjrhqKUQ9wOMmq4uAMwlEVCGrc4m
Fx6dRTDxuUmLfu9vDBp5ubl2nBlEGWAyFVJQH9LkrwiGmtUXVw0mVt+gSRmCNMjCE1Cjc7Xnwe7z
2djVYcOcyXYyRM+NGjtOMFDT/yTo9zBJl5+0QZ/C912fmKytKK5W/M+kuCQS+KhnfJLAvuny2Aeu
2jcLFYGG8/YHDkr0lOkY/y+GDohqUTO3Q3z/qEfLCpAxxDf6UfSaCb+6hf2uVSus2OfVZ/9w6bm/
CbkVM5W2aRZkLeQCgKJTbYE9aIJ2zSTEy/ErujSuKt/Fe7RCsFbKy/eC53qQsC56zpbY3j0nRJ3a
b7v4hTdsr24ktF1OyoSBVyra9AvOKn0SnZk8SiazcP29ODRplnNZfovvmuopSXMAbqpuN8odLW6N
FpMewTwEPKZxFvjUHQPnJ6J/q5buPCz0Fr/bWTp3GXVmXtRR2CUOng1AHPufrDYJ+MBOK9TdmrKc
gIHttXV6iTw5SRnm4VUGeXBuZ1Lqu0eiWQgcAkNpoDG+fwBL6Ibk2m/ECd2XaS39gdVNIH2OjeeR
CRrmJu3uKSoKSO4PO+o8u5D1j1kB/QdVdeQhsokdUp43MXgkQl5eA1dgPOmyWBAb53S0v6rpl/vL
6/hdKUhbetRjzqFEziw0RNDK5lQObqb+WOo7dQFhF3qgGyxzd0KlXmoVJw0yHPUEJD6DAYRlopJT
TLwmtg7+lkPYunRW8/4I34z0YEmz63lTY8+mXVxUyBXMYAzXegdYrL/4LHtL8qVqz0sqnY0EUGbh
TKe+xuxClegS9QemqnfCx1JO/frV9ogZpHnsNoNutPF1SMnDZ4kVtpv1Up0FEXuNFEHjEGdJKopQ
0YFNvBTJfWR7lbH71buFJOqOUoMmtjokp33nozno2q64n/KYiaO7QwbEow9Ev/ff2ECEjpljkD5h
t+7K7hduKPNIHCfCPGsiztcWiEQgjXuMBPQJMAnVgTALc5jNK62mQ3L73dysK0P+uMp6wNXY+gm4
Z28dHSF/4m/tSABiFF6zDlcWHsc04lt22CKQfGSuUf5O/Uk+H/H/L+PBYNjv02mEpwTQ4ZwB5T90
6OIEWwFcjkGxALAdpnXVBQz3UQ29d8gvUzLNvHWjcXV5/Iy8F9w51pD3Jff+tay453MN/oSODWNY
OTnCHysRyOZv1AY61flIY33QL/NHzOnShl9A+BUtqL8rlXBM2mGqNbuQJ3vB/a6lAQEAmf1JKVal
cvOOPPZvnJstS4IaUfZJPUde28sR/wbDGVdS4ALvCR/hYe3P1MqSrcMxU69GgY34LpvRBCvwhy77
Klb7om1UcqHiqrU/aCRaqBW17nZ+o8aH9Gd/B6C2y1+k3wsm32Hogh2/FRodHWUya3/IhkhODK87
x+NuqXPwH0HJtTJPx4XoPKjk/pJaRkDrSOQ6lxLGwTaxVIc+HPIXNaScw9kgTChTDHprUU7+PnZH
DP00PwmhhhVkLi/it/jz85vXosF/hvq0tULPi29FueahYpMscL0os6dM+M+xsHCFS0+lRZHg9sLP
vMhzyDilzphOMWYm0Xe2aHiBIDbOZUsNEQN+8iOQ/FPLWokRCm3MT5pt6V9rhcc57qVCDhaTY5xI
hVTTkAEzU6iVtSOzEK2NnWZmqyAg9qfUBsSXnZuWJGw/uKxsoViDm6yxto6w+1j9/mGcKR/X9+N1
a6XFMOTBq42EYChpFdmqU/4pg7D2/pSxCxsH+FSzV7xnZBV4ONOJI0Kh6cM0fpCBxKTEKv6pCu7Z
zgdrAasMZ8OxWwie3D/8zVZzpF+PmB2cmCr3m8x+EDgS5Cj/Adf+tJvUTBek7aXpKW/xxE5de3O1
XntJ6P8w7bwry6vPH4ykbgSvk28XSFtw+kIuHOuhsbJFuANBuqRooWP6tcqZoKRALaH/AV8QeHRD
c5pHx5L1z2thhfwArEpXIZ5ABfOMB0O+iRfxhvDDPSPsFK+ssvXuBvQWxu13M0vMsu57s5RTrBug
IhmboYnueiMe8Jhp5ktDYEivhQPhhKDlvg2Y4Nw5q4tILUJi18NNo1VB8KstG1BZXJCwUqR7qjls
54sj5tjbxNZUywu24w2SB/0lvHnGHrCpuuf6qJ5H39J4x4NlQjPvpCy1MU0QB0P21yQreEcDedRo
cIkbn4LxBesUw7Fj6wQEQnvoFvfiY86dBKo/1VsBIoZvmTHr3wm5Gugb445EAuzuF7oquWpHkuDi
UuFiAs6EtD0A0VBiClNBxW5hBb+HhfQip9kvjOO/4v+rGzaeB5oHwLjpKTAh71rFuZwBE73cB4uy
1AAW2oaTcMO6Xr9eb2ZxgZE/F+G2oQhdhos4PSNdgbewzWI9XWSL33gn9cQ1oeMrWcCOi/By9I9f
gawJvB9wyza1MBuQfdBStVJHebYV52WkGEqWqbmf2oIrQa86hQw8O7T8cxX+5k3HZs8ieURDTVic
GrTf
`pragma protect end_protected
