// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HuEdowXIT5OERCYomI5nh0P878OMJlXSJo5vjT8Rv5VUYCl7vVso6ZFt7Wdm
IborbwYk9WTpJmKHania9YjL6DJkAGlH+9PuYc94/Oz97PViHn74+0gh2aBl
izl7RcNaZv/+hg6gY4SSqKjOKZmSslUdgrrg7TjaK3rORdcNxmnyL4A0QTvb
PiTkFIG9rLHemnr4o1wPBmJpyphpgFSPck5WXgndnefO+aIBE0EpTek2+uPg
Pq7dHTPHEQ5ShL4Y1pQQSefJFYvKjcwnxLJ9j3vWq7qkKF7qT5AOxRiBY7DX
u0HI5bCmneUpXLo4aUAMWqhFiyJ/dETTwM37yPK+ug==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FBStPwWCzIT55JxnebyLIsO+AL3cE/hVOoR+xih/am/rReK/g8vZhL6ARGRn
xmYM/gHi+LPTo14qB6z0o19s4VTFSkKFze+azXcVduq3Di242d/TE1WLc0+v
Uy1ljk/SLkkmCVAWPBsik3o1mkYLe0qHGc3vtl0I44m1CDpJSp0g8AlVD7h0
nE66Hs/X4LNYGgEj4oqWiFlvGiD3HFAAzJz0nB5Iq0fy0Xgpdl51xGsvaBE7
dmyC/KZjya8OJ5gItRztHoxcufQ5RotEmH9fpvwSBm0mKYsw1rya1TW71747
xEvOCxAVBFrgXkMAgY3RkNMDShBb7uFLAHDi7+frpg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TVxebM76cQA0TrKpMjo98ScKEKMsnnaplfqLdz3I2CER3HaHtSypSwotIWwr
qePGJIg9LHTB3yNabsfRGzDjF0wmHAitqXegKqa8ZCNpfVdDEc2Z6YU6aX6a
6hBJS3Ut2WwAYMnrObkZNzefXzYI7NiXEfM7ZrHke5XXciSVKLVnx4M0tWAM
6x1kGORpJBKL4VlaKobE8O6phcThZzVof8SYm5YiVCSuQRen8IotxLlO7llf
ePUA/JR6VtxQWv+myPs/XEiW70G2sXz+j8Ra468KrglyEXLSqPscqhrjGWVG
VF73aiO6+4TpjjzrJC/55SpwFrD0I0aixJRrt3Waig==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qdkPk09PfeuboVZ2nfpzUHECe7fa6jY+ccU/pUS4bfrCy2VJbli8F+uLrVph
oN5Z1pmROKAAVhX62oMtjzMidv8kZ73AiNsKXV8Uyq3jqjz/JeoFcOZCG/HU
mkWFBzjGr6SMe/icblQNP5UruCsgQ7fnTLVCKkz6Fd60Uwf38TA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Y2dgas4VOQad0NaakDxqwf5wFlMiqPNJpGyzeAj6inLE7KbB5hWVqdEHzrSs
XV+77O9lXtup6LgmhpGoAR/je47QREpKDkQf40Bcozi37olN751z7n+gajLz
ZIPgM58ATx+vHfNeW9xbAOVU06tzUR3pA1IVFk3LX/YcGpBaacF88/0PVAZj
GHq/wZ3yd1DQDO5ruQdNujcezLAGgZDQLPVqPdVkRLiAkjZtujGuAMwCtSDT
SvJ3RjHk8LGPsTBedJT8aEwIpBiLD0SiM00WDn73m0vsLP3jerbMYGs8pUet
MQwHf54WaCFExvebasvv1WxpGKhN8uhqMKx2h/8Qx1gP78qKNrfOGoEYtjdR
F3qZIMcThX6dBgpexLuLfHhYb4WRmXMOBhp5zjDOEyONVs1Yhof0IgSoO+Od
ERK3qXRuer6aFjvgAcyoZumdyl5Btgg4yZ+niqVPmNq3zhMHw6VuoiB/Ae4y
gMd2aK8/PNisBa8kICCgoyC/7cUsBBDE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hmI2U83tIo1DR50QFH6ra/Jcd7OJ2t0RgtwBzYWq+5reEcx4WWYgGLWimtpS
WCk4H4/qXYV4n+0Ph5lq6nuXBwpppvdThzZWyjizBy5Ky6BaUhCuGH3T9s9K
xM9mWb+VmdXIQanHyYR+rjxGECfLMQZPrgdpkwvAvgpUcmMYj7s=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IVSQ5SYyHIVFJ6BhNwNqYJLjyzIjOvuF4expDqz1dC9hBbdRGHbS4yl9Dzw5
a/wfyGCbIHg7ZqaObE+iX7R8C6ke6wOXKDO+yPGkm40RgDsaYd0XJ2AnFs+c
vsmoKsJG/BZiL1q+K0DP2cugLriAtmQBpSqsZqwRf3V0HCRHaEw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7360)
`pragma protect data_block
/mbZ0qwb7A38bnB0AKz/N1zFCZdMSLcn3x7oANx9wtAzGPm2XPySx7NDPbxe
3TBERSf96icakkP2u2UG1ZNNuZDHsS8zjw4ZUZl0Je4MmtZlDzY2C9jpCy5W
wSTRnuQkxkWWcmBHDlbvzuyZ5dVqAFLG6b58GpD92WCpZCI0fXUT805aTcDx
P44I/kqCS9Q21lbKXq94Oe9lu1bxzQUksXLa1UZ+Qh7kGViQKko9pX7rtL5d
L385Qhi5o1rhyP/KKYf6KjfLqD/JYNiJNpJEt8LwBfv1uUKW5kBjwvQ/KEji
+NmC0MC8yxuTDatNibmSJW1F64aZDUcuiMQxRrLhuHroP6KZg5xnXKyAtiJ8
RjaTWdk0psTMILvN+z93Jx03T5kMjfKCTwmjAxLKQfVG1/bA2w0nf6R8K6nc
zCS3DARVZa/mRKTLWmHdqAggtT+Oi+SfPOhBh5ajHge1BwU75resoPe9OuYr
5hMLtanRdbGiMwvL/OhC1HKPFaUf72qaITHIfCt/0LF85zVB7xpccTde7hZE
iHBlnIqvqh4uU8zxbYZy6Sm9QzL5nLC6J9tSSPVVKr5jNemrmGmHx/DRhAHR
9E+5XCCNw9sgXpI/xwQGz62TkTkxaplil3FiOhbwu7xO1d/CD7vjTu97upn9
CQWvf1qFXybmKwNteQXgieioJWsGxyhy2gzCd4kXy7aXFoIzy/aX2pDNhEf0
17xAkAz46WkE7lURL6vUaQwBLS0E+IiXF9qN3K/q1nyo7b8+TGELvAKiYOtt
lLRIYo/Ap1Io0lHXNA2tnfo0UoRskz2hlSFTQ1NyoC2hnBBedsBcHxp9TukQ
CYmHxjkH/FZZdC6q2lp0+pNa6q/QIH8hnXXmn+LpsOy0knIQy8bND9RQMKaG
pTGsP4V+AfXyjIipBN34C2Hlw/cFoFK4dJ0+aAejN8E44amfuj47t1JH3Vfp
o59RFX2Bk+0Nr3sktUH5q7zuZ4u+d6JBsBDSdjVo7akYUqw/3HGNCZlnu7dr
UD5qzzIGqi1pSSMs9JOCz7rcs65+h8GU/cuYn47AX7dPW6bSjnvaUPs7vs1S
fdHX+VUibQPHKwQEOl802ara0vLLgaRCZVMQJoogsdW8XL7LsEoms98BBFYm
+FBfghoMpKmLA7mCNH1Uk2v1h5dcMH3+CHiRtZPTdqkuzvgZo14cvhG9uXaB
P6Sz6b1pWliTUb87pV2eefjXtFtAMWDSHOaVQgCFOlhxOWpS7KXhFjDVLuNa
lFmKqDFOw94pRxdeM64AVJhvvRqAXQvs1+9Lp3/4vtxgZPlBqMiLDA8x0pQB
i2lnDMU1fbj6bqq4Ktevu/C/DtjIk+wT2TDlDT9WIuMz1zipvuH3pHpEXvdZ
G6WSa+wrlvIbq4AZBANYdicmMedbis7VMa7u9Xhlj5e4OdrxdOPG3R2zY+qy
xQMX8OWTC6QYVb5qHtse6Eay51hj98X4CGIzIR9MgKzlFuutgX76rwFATw0M
CqkDd/qsyYikhHrI6GJqO8xxnoBDDHNgmU82z5FrZvBQYteoj8TnzB5NL5rT
Lpr0CrEgil0X6u3UckUA6oKrRWuCls6QeJYOREYEQV0zyB8osJjfVf/+aOqw
XoUii4Dc7tfa1BO5FJ8W+S0xbgILbS9G4ageSYqsNAjPw7cVo3NQQMqTsWVo
27wXWBXtNS2Wgbve9Ol2QEo4La7lBw1sjeSEy989l65R1PB7N5iyW88gXHRS
wfoy0+09VQWF8+B5JYO48mM/9ml462Zd8V8Du5VgGOevH5K1K26qP9+VnKHj
miTLovsQfmaiR0oK0i4Y630b+xqe11khUkckO1LL21q0pkUeo9RU5clllSbW
p/7yco5AuUIz96TLhEqlz2uDYhIPpn8Npu6T192R80GCOjxMw37p0aUSeL+v
v7xGw7XC8NaIcy+grmBl2x/4NCyNdVhZ5Pe7Xq5IWotmL9IO+vmGu9UX0PLk
Thbppjhw9xqc0zIA5A/2v/2exhome9a+9II4HMBVabjLGHpQi8RJHvItwf+/
onuIbiHg7B8GBtSUKYVfQQGYDxSXWsKaYtOrCW3jk39CVm1CdfffIGJm3cnj
D1ujT5wW804Tel1ct7qpyawuG9TpMwEkqaPki8jTomeymiY8CKiof7RfEkaG
KVdn3lPTKByTy3ByW4XBQKj/ubgrs6BHKF7yZd6J/AAxsVGvV8aVpYChsU/M
ZaywF00VJPYt85tJTA/YykDnPLK22D9qoZyFvcfdtD1KyR0/bylak/iSGnvt
Ug9ldzWrF5wKKscAW/cgXcqkPQVcFgqOp/mTEUiL1d7gkRW1SZWYta6r1joe
iZTBySExsAy2M29eird21CqzWnN6njTHm1lfGcjh6PTZcFLmFCM4l6qOk9lT
Gh4/9PZ03kC3Ul1Q29PQtV2jxOsV/oSXJwtM+6Jn7/SI2seYUe5KbS7jyBfA
DDZuf1JaMl8ACC65G1rx9SQHhtKxOI2Ntq3LjT+9g1IxhGpn7MB/bWMfNmU6
u2zLGh4WOhqqk0SirYxUXI8xFIhv471k+XmEF248lCOcO24yvUhhwwbXDpwj
eKoB9rPpym9amSrI46j1RNodaVWFBA1J883pog92EO8CAjYPyygT6bpHe8rB
DhQYFwam7+R/2Jl3WnjpE2/+4IHkO1MNng8XdgTQFJXNOHi+cJQ9XyUefhmt
d+Om4CzJaWC5ZqRZm/8rNCdc5EZnVqQz7Y3mHQdwSdB0XJiIA34apMsMVdND
lx13s73faUWPN1nAl7Uu1myeuCmhuTdVvzN7+hd/ZZL9B/r2n4Mz59lP2ZEG
HIYf/zTIoGg7uZJtPt7YQWh+S6BpBJqxjqM/5RdrLRwczbmnJp3r35EJbXRH
S1KC1ScNI0RAB9yK1kq4KkkJ3o3Yyir1qO7lIBzNOW3oGm5jEtso+UVTIsvQ
OsweS5hF6Hb2iX3j3KzziLQrJ1uRxtWCGgRBv8l35zqJh6aWNAqaAdD0dK4n
2jwQlVhSAQLRX1EYeeC9n6zQ5olCbO7beitfpxfP6b7cVdLykvPcR7GjJdVC
cTvRXne3tLmaAvpqDTj39tAaYefaYMj947dmYvlqbsTWlgnR6413+uoR066R
smDSMQOPczY+7kxTBZGrhfcb7UEoxIfj5E5BMBAAqMmVXhmBBByp4ywTRwRh
ycAXTriSgAbmxgnuClgveIyaEv5/dhEwIeh3ria5cpp5jm+X+qoGfsWaVX84
M6VrM+KS4Kft/CAoEKYyvxQW1r1/7CAq9Id6Y/QatiDkLso6PPsAC3JaAvLY
q2ebZQHChfMrTPd2Qtiday3lT0DQiWC7OiLmsQTgCrg7WDARAnl2DCUV+5bH
4h1uKGOgLPH15KkdGIW+d2iPHlvDMHEYzHK7Aubh1UQBxmPoupdkfNbFYMAl
skvflmaPfBBfTB7VEVONMsjvJ772vtAX/ESrhtA/rdBjgZOtAo0r7+q2o4kF
Hjspu7Dzgk7O3eewisB0l2UgpQMOpfbvDnREVJ33mWEV7wHo3SPgBeuO4DUz
iXi0vcKBFc6cgS0v+pp3jSMcydRVs7ncQ/m6RCbClQ8VjjqunCOEGjbp4C6E
IC/A5+PYlsO3RTzbTlBzC/hZ0XElEo5QBJaMvXZCZ04wA9gDR1ew7c13Xy9M
GxbyKazwLd0GnH3UzraA0M+n3TmMWz7mNvzGiUu716cMOLD8jcqQ0afv4hcp
16r0ACM6Qa09DDbBvPCuFXGCGk89dUludaB+LvlgczkFOVkE7jHBOFPbqNc6
JOPAx8L5DMtLu4TrtIVGnHmlDZNIY1suuZKPDbE73pMpytORsj4qMB1Jx6cy
HAOai34FQvScmIIyo0abHGMQbI/XU4gX+DHCWFGbwfO9dfAVsT5sqjIoE7Kn
jQ5YhlSWGjH5Nda0utvpdhMmpQCLHiaeW4ZoeqDfCfyPmRx0S3W4foMeiLBY
gRToncSg1yAhnBwcvys5Dyx2KgHYC/ZrtPQYtHs2EwSD2S4mx3IihRWyoPs6
SDokYDzyZOuIdd3F2a0jjAiepHYQa/hceIrHCKWn+EA5Kt5rKBQFoTO8zsuD
vSMlzeIrLa16fHepFrJjvdqM0I7fwZG7k/oXYor0mDGFzc9nW/fSPu+J48Oi
4t5WyUqezWabGHS9Jb9SnxSGdY+w8L6nGftmcrS9X871BB+jw+CZnX5bdG5a
SRpRGs7Z+YSk1zu72EPE5n0H/eeQwy6tLZ+zCRYrZHTRYGGxKGqRf3Y18YAn
Tgxty0/1FC5JMPqG1OAhcwHTgJ017JKaImJO7UAx2CoXgJPBahPsrZYEzqxy
r1eZGD0q4quRfU0W+IZBdrJjvRhhzt0JpB/oXraMHM5YQ3XY8/9KPTWba7TZ
Tnq17QYy87UK6xGhPoaOQ+jsmHvbomVQO+iaIWkaeBq2h0nqaRcxz59e1U9n
fZz/yGzJNZrwzjfacTJVrIa/UufjqkxeXaFsaDpjKa+IkolmurxBtO7P531K
xQtUkrdgB+QwdKidBi173gFETrTuu20dwc7uo1Xq8f9bnsE1BTcIqo5u3jdy
fBTKC4RtT+ywFiYTeX1QLFDkH+VLNWvxX0AWOVDZvaNZbgVMZSOVNdY5v6Yq
Ku6ac88g8pu0KDeoP5Ujt4vYf1xAZYSkUFZRjIA0J6hNQy1bDOQWOQuBvAMt
KVdQRHbnUG7ciOWOenzgImrq/CAs+cwpxx2HDpnpeJqmloM0vUJcRloxH7nk
wpy0lnP6Ub7eevF7z60qfIM2AfNQEDoAOZ/Kmc6JvDXs99N4YaMIbWYjDg2l
jbDGWSDBKzTxiZuir7Tl+236AYvDik6wYjnqep//cBP6ChBGivukpmYwRQVZ
VpefF6QEtIfTdXVEutln1OPTwrmmHw9NKLivxFLy7zl+wEcABus/0jHnRy3u
kBKi8XasfPBWF7hLFLjtUY52DxppASR3G1JkMZtZCAIAzJI2TTU9n44ogcsu
PcEqmwuNBUhavMw67df79xKBfbiJiGKX4AIUI2nXrHfdXM2awg9WLVbZmNFa
1y9NcDPFd2Ekdqu9ds24i8A/MPeyGEZ5fA/vJ/Fz5vaKJCa+eG/Lni77K6SQ
dIHEXtUbtZB5xvwlhRmxhlGJVHB9iKQrmmCfFY/oh8oZr/Clv3jtd8FGAfrI
/v8s1QZChns4KS7xUnD1AuL7yzM7OrsR3TFKrqf9GY/8Nu7ZqkXrTffhxJgX
m33OqB/6MSk9OkwWDXh3c6YCefUz0XaMK8xwT0prrhqa8QypPlioJRslBE4o
rxQJR4NAcr8iUO/ZKlnJr/NL7oRCj1C14g8Gy0m5iwuyuEpcjHoQb03ce8HJ
WYuHXEQqro1n5832IqDfQ7FgiK0xfy4SVzdPy4Csvxm/J1L+jufkv9SKA8PF
OHcc82v0KsyEcal3BChA4jI+n3HtdW06kXq80Exu2Csvf9stQEUX3wzYgy44
p3YQKzsJxOAnZvoiPkMSR92rWEBFnY+cvj5qUlbsvhbv/l1+ty8ZOGQGVu7a
RklKCjh5Kfgx1v1Ba8fuhXdTj+FuKLjUKJMsyMZV9TPmWhFQM0v+Cap48aLG
2q6BCxIfQgCe/dgA2xjs55Ykv5bCtaH1k+DPkunU5e2maicVdCWOP8X3xNCM
WFpTr4yK6r3rcgWxKWhd9G9GYWbozAfIUmyvwGWbFaLPi9TcX2StjnIQyTwp
WkNCt189lRZpeGqOtZEjqWt5iB84gG0ttBoZ5eFRDxcWALi1yKoJUdrMZ5G0
uUiVHv5WZSQxEx+FyoVUjDEKgCLe1nj48fXkNk8Qxzky16mfV0mN3H8jaESB
LKy+Sdneu+KDc0e5oBr+kYplR6VGWLSBTu2fKuIfAnikwku79sgCb+8HVjTq
BJM2xUivA7X1iQRrK/lhhrr/hg/Vp0SqsipM3Kerg/iuL2Y4WbtnoPuT5OYs
/386uB+++hfXOtWufPm7ShNB0QG+ix1HkdmaFEAp5ktUw/fwhqsHDim9Z9lr
XXKfjpVdD9ri3RuS/eSddQjM4aQoaqH2fEgbZnBkVO1vZOBE891MsDeb/LFi
k2bW1aXn5ppTsHFaQLJCz0Dj0kSZKjJir/CKN0OwD2h0aUX8WtcO45TxPzXP
8C3LhlJapjGPWNft0/umcsUh2cT+3bQaudiPuBwmIMFHgo1DkbbDwUkWd/lk
GpcO3VKIj8+5kqadxAAldAlAeQ0jdSleb8Hx/h3cloxpAQ8rtoAUBAbtyYkj
Dl1AiUCoEy7OIiTMpQbbxBmW27SZeiwpVaaM3+crzjacyxgApmf9EwVauA+s
nlF4cfsqdUgwvL2w5O1xylIZq6f1ShQWQ1Y7116ZIOoiQw3Vrh3yEgFc2Yfw
RDryV2BY6hczJSsDehq9MgrELIzPuiYtZvcORDSNIYbiSWn3rtMOrFW93yfB
H+WdBRXapMPiU0Hs/IlgPt2Cl37HlYm5APagcv5nXkoKhhszviFs4n/lmyT5
2ilStOfQDeqo4nC14KHgIlMsBTQYwjxaxZR3w3B48KPKdT6x0+6/uEdmNgOH
3czSJF4PyCpi0BoE8Jro9MIsbJjxMjal0Z++Y2j6jXyUPT7Z6EENJiHj9ca5
ihbwpya/mWMEUMl54Bpf3BJdQuhPcjCHzowzh1aYfOkhWQX+TUuGZPNaTM2L
FhaSZC/rRNpzyy/EAKCYOQv4neOzTEJaeomr64VY0yRo+Z+5xlkpBhw/Rhy6
YG4BCT6IKAyJEvXDUs7lYpGQMz1mtSXVA187G/QWKM2U7FpElFRUusGtQRJA
88f3RqD+5C5egdMDTW+a++Rt0MCTwXo+eboEF2GGJPDS+Ze4FuvNZei9+gw+
ThYe5B75A6pDADGCQ6I7X0pT5CbfsWZ0BTqHb3mQRHKKlcOg+0gnEqZbhLLW
aJWqAtfZAOYV0Cs4FhRMvVxMxNXYctt+DedHEjKB7StKTYIvNqHmJSP2xUUQ
ytjX1JXee9MIaQqKnRXwaka9X463gB+hNBkazmJ/laElNTVr8r4XgL4rekK7
o6sClv50Mj7IxGGsDN7GueD2zkA5TXy4M6ax2AOy1bXFxFgpqVrJg0ptDxub
G7dy5PITXOmiuqSCUGYxfjd5F1qY4EyLFD+Q2H2sJ5gFIsMeRorR09JS9ujV
H9ijgHEZdBLa/1f/sJJvh7mKEkDGHQwz2l/eKh0qjMcJmI1chOf+TB9EsgOz
wDOY3WQlfKM5Xw8jnMO8gjyCGeA71HBpayTLa6kVbg1/L4iLtKqYoMnm1GQS
z7J46FDyT1DJDuerAy2wv76q6OoUXJKif7fxWHfNYK7WJfDLjG2uwMWcDM6U
gnJ0amKV1XUuQJXNWwK3zamBymRBwZ36mcTfsUXoo4/KNF4VtXWH7HmXq/rg
QZnSTGpjp3e8iSmgrykROyHusqnXZ4dYZf2lI0t61osZB8gPtoYl9n/zu2bo
b/jFeEdHB7nzH5E6oVX83wZ+DJvtJnTloEV1nz/hMkpqmmB36zQMNOhOTZ5G
QgPBCD5G9Ku+SwC5NAh6BZBrN9d3j1Y2Un1aUGIZ5OQfMwjU5YR86tLh46J3
Qq8TE51KgIvD1+LN1p/cGLSaZH5SsxneckI2x9DDMWTkJd3kcayOI31FeeYq
Q9hP7VQRaneXYCvbd2+S8n9PtegvQGumEWv3CBn9hiwuMkDO7Nb4TLi/PNeM
dxrekznPx5eoYnyG3HoTYhqTX5d/SgR8fbtz2V8dKCa1q7MY7Mbr2QCXLSRY
Wlf3cSZryFL5ON58KINQfN5TFuaOZug7qTD/TErh/DqxAOYsWCKaqko9/+RY
NgjjBbW/vlIqM6OmkzJ9m/qBT1FnrX8FYx24P9B/h3eIxz15zan/Gy57dXQ9
XMCBOuC56ymk7uAO1OJdgU0pCgZvUzNotIhyZ2/V9msDtOf9M24+Lw8FAicU
QIC3zE4e8l4nSE6tlP2GuBUwfEHhfGL+fCIUYaxENnccKMQS0wSPSdKNYUGB
R4MonfFlwuahNRBGICkxrkFJjHL10yu6mapuxXc+8UXFBFdQiE7gym5v1z5J
X1P6QAq/VDGGz4nZqVmXWX1SnmlgR2wH0HIaL1ds2GXykBs8TMOy9vBDmhLA
VysuAI7/pnIoJpeWs7P3w1CcPiI5T6no2X1dtjp6IwlgMmJk25xK2Zc6hsZP
c+gZAPhuvmSc3cL3V2osffMoFfTSG6b/IsOcUNRPplSwZ+pzeZbjPEqyJ6Ic
4odI8xm9vgBiMozCnuxd5S9ZC1xAaaMj0MPlcZxlGEewZtSxmtr8L7/ZGq14
me82KcD6fhSKX+sg+7AyHGKkzccWofTAFntCa2f+1j6W7rxJGUsiWyOgDeSo
CWOPoCeEqdMhQvAwTR/V2MRPO/InH3XcXiaKOmH2570D09HEyrDG1+eAnzUh
68wyPtsOGH1iNj/9SD6babwZmbDz0Lvnkd6JXCfjXWjlzQakASf0/dRdpx8w
hRQ66mL1W321TkJCvY6OQJtoP93qakJ7J51dRKlPMv4vq2GYkEmknuAafBmG
3+OLgfDJ7RXJOXqHJeYP+t5RCwWqnh1rFXakjj8vN2to0Xm9BogX/AgGcioI
iBE/gP/IzmBmczR2BnSsd6NhVd+YM7nifSYtIKwItanT6A/ZgH9oQKY+eyOX
KHm9o0OFU3xbm1uK2ME1PsKdysng1eTs8Yoj2WZ4V1AgDgb7zrORfRSIpJUH
N4LPJWVUujGK2uSfsz99x/9RC53/0NEUKmcG8TIaD5DwJrh57pNUbuzPtYt2
X0C03dMGh0tTfmppF1BEOiL+MYAHJ8JxvsITXeyfduEnJB5VtbGc2qK/WTgV
aVggxp3yUa9CL+vxsgAZmWWiQ1fWv7GVabhhIQv8v8D7MNXz5GGF2lG2fsq/
cTiismAgiI9Bm9oIEM83vn3ag0+xQxrnrn4EIzc6soiWY8yJN7qk7R5PWuq1
4ZL9ncJYEUwUavzQ5P+Z2CUhCRAWgSY3gRzEHSukTt8JBniWdOXuvUYpCteW
xwkRo1ueOLlFl+Jkm0B10WuOj1OiBfFFv39615vEbHOTAklLpEaEneb8yJ7T
Jk1TS2yrTzr484MorfKuiDU+LMkUpKjZbN9xGlI8k4bpF89etxRlMno4TQuB
qHAJkU539w5ErR/b5LPW/2a/C0JQyK8kHqbSB1lLn/I7G7Vc+yo7B4Tcbs1Y
R7n+y/KyIFNd9nr4ACiNTOI69IJP4O6MJrCNXQJY5kz1fXA31PVyOT6jp0qA
xtvNS/YcaHb0N087wpM6CDuDLLA+jcH5Ox8l/NbFjjJq24JFdp/bhDSP7iky
IDRgODT9AGEGdVXZjo2drSGo+7+uixZ3oJ2g7t/pyZxwW3wF/oNLPQPOZB/q
MsEUwOChvgse7jKxb8LLWxOTyfSduzI8wtE2BxrpsB+WmcPFXgiWiPXlD8vv
rJe+HzKCmGQRFh8sg95jcMkt9pm4rmqXbNI+vtjzUI0UHEjblvp49qKVFcVx
wJ+oJP3vogphwMN59K20Viu5TwqHOwxVzc3A+MZ9e3eRybcoE9N2kwW+UXn7
A8ULBbpLGaKYS8MEvwiUuYYbmbTDDcqfCHOGaByr4ufX3rxCrsmc7yQf5eD5
3fcb1Ke7BioZWntxUyhOeO+KiepY5cuoQGHxDelhXRqLrabnAuVwn79Je47n
6ZZ1lhLojzxpJsYg4g/SP/ZntZDsbBENWgTWMKBaD+Aj0V5vtQLm1WMKoorq
PC+/NCJKBJxTi6uSMac60+AN/Y5vFQ040i2RCG0ZaXw7ZY9vVl9krBAgDbpC
esw9MbU5tSxy4iWwG0wAl3k9unYogOmFbw==

`pragma protect end_protected
