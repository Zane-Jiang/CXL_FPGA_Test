// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S0R7GZUG4Eg7O69m1KygT6bMC43s9hD+KhACKFxMatpfIcOLyLLuw96Gqls8
7QGNmRrx/zNUeT+E/PO7DOa6uPN9t5kzlqIEM7E6HV/AvMLd6ZZ0D1eHpCvg
7WQhUq9vSWZi4oliqWB2WwbwdhLvJkCFlaYAuAZ0tCjZE8SpVj5951eo18lB
WUAthDXjYxopkcyuE9ehPbdsK4xjROhnuqMWDrBo4G81bOatI+8bD8L5dt7P
nzRT2ngCPF0Yxw910wdkiEQOjf59KicfzA5vngWkXbBMAwq8m1Z6a3foJyu5
XaYIG875WIIoAoNfrGTxsbbUTugLpag2QpNJkWuXnQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VpQpjwS9N65R6leSNgeQ5fEzcH0PJCtlXh79f8u6VW5oGp+/OjmRKr8U1Bjv
MiGhF59pzLIwEbK/y7se0PgzqlZtxBbGVBKI4iFlFnS0+JMfYLhvDF8tOn3V
iUoYu4rYeHgITcudHCjy50Eq5JEMaHpL4v2iTSVOvykHO16TypSefRqZZosJ
toI1D8OKRAgQRVKCGVZ3Hy8wOUFs9K90Q10Bfh1xrZxWrKIogaLQRcGzvDnB
9va8v1Kxx9axSaagaTHWtI+HBJ0lqzvc62MGMtNLiJJHrHKG68AomQmePR3z
GFmgsq2cWNR3D9BQjux4gIEGZG+dEOJD1qsPo/hisA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TgArQ5rTyqxzxFdUEBoP2Pe0taQmuWCCAsJ26fDW2g/CeVGhXtuYsXtCJj6y
qLGTJBdMwL7grpTWkEV82feaTC0hnjzDV4K/neM0XWw7pOGjXsFJTC58pM5Q
a9BRdp7yHhroLoGcfEHZ4hYP3qqIJzXADvMa9Vdsn9sxwhTPpgk73IqFxwzd
bc4wTHijgmZLNshSYPXhKOwYxqXmKHWenjBANMaSreIpG0TNDzrRIVMbNCiH
nWR0/Eip1hGzJ9PvUFs9O+nxKMKHNpY6BpNCPsEjbP4tGphCugocZ249xXRS
ujpUYjDK+gPHAqFeaFLToVhopqMgzniZc3ZxBlcI/w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
C9jrOv3zzLXOSfZPZPqPf4uMd3bGmPiTe+Hrac4lpKMC+D8W2wEVli9P+O+0
JuM+fVTy36BjuR6gxaqPaYWS051viewB0vfnkrBrALdT1fHkHrTNvTRxevyG
ISF0YApEmyiIlCI/ou7mef3G/fh7WgcF0y/fbzzCnWTIh6rj/PE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NkmZz6FCtB9ts85N7pd78IaM+AL+3k9R6knJOMxcAx9UkaNDKL8PcT+2pXug
x9a7bRp3GJa83XSEezveb6SW+Neng98GVE6B8zfXHhWFa7KMxaGUfsjJTE7y
u33WJQ6XNVlHACTIZ3BW93nlHuqCpiY+/tGmVFWxyvmoyvKEkf0QVjzEI9Q8
bmfASb6zBBUiu+m2eSlUsaxhuKW3PnkKAqNVOjeZYrCwkl7A0Z/7kYVn1Mm5
o6b5WmvuZ0PXeYekX2QsCNzGUEi/VpYNj8+FRBrLY2aGKJiQDDirLO8hw+G6
EmpR2T3eWZ2eTROJXPaREXtfdID8+yK9JuxSxSjV9WD/b4Y+xO1Y/PE7vPsr
ylfp/KawoB1MbUc5oGDZCiQI/YTgHj+utgcRuA/oW+ZfLHlPx2+1jiUxj+ok
KAifkXZmT6JgpTOYAs9aFh6paJnu5jHiDYYIFm/OtRzt4BdIflEgA1cLU87C
xLYv9feqQIq9LHoGkryJdhT1aDD1BePE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kyNg08tWg28f6AeVCfX8lAKwB/AlXi+57zUE69/45DQbwDpvMGJ3LpIfH5Y4
tjAU0v21EsspiWkWPdLonf5f8y/2p6g0mQnvXGTQ+0wO+JmhaGTuZ9IHHKnH
5f3MnNxgN7UmWdg35o1YL2qBuFNIdFyqx8ymX5z//RauJnmsZFE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TlW+8YlcaCXq7TH5Mh0g6UQw5qNQsbCmqDsiloUsMETKXPVlpRgRINaWoy3S
wz7Ns+mePZeroofoAoL8XfxEsvKZSDqNfTL5OX/75boWzd0dQEqQCOby8s7Z
4CwzSTmElBo6sDmPg++3YqwkN9lB9yHUTLkPEkry3BVmlBBtfYo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14960)
`pragma protect data_block
EK8dadq2MXWMCZt8KCTHmxGALNSzN8csWM3s62SVXcT5ccQPFtRl3r6bqVj9
QQwxAmFxB7PsckfVo/37OCkiek9dZ0/bm4Qw8I0Wa4Tdndq0euUzB256R9w/
XFaGckivVRFJqQOszIgkFf7H6lQmzAhoc+4ofXRb66AKeNKYnDl0OTuy0wFv
vt5w0wP3HE0rtS6k/El2rBlUAa+ar3A1Jicm4cMOMIwWDwtRAt+wCoYWwhJ2
ZwetQPpOhAt8SMDKNiTdLvRpeYv3Bs0s5BiqPnznm8HHdWxuHKxTP0x7MyLs
l/6iLQfoNzPyacgf+JvOKig1T0AfViIHh0DdL2cw20K2jr3LPqlDtkoomD7G
ZoNoNHkWmxWyhuEd6XghsBBxE0yan/pkMsRAeGGc6YUDBuFUATZDDJtxqvCB
gEv14XKK2wO8Op5I2F6PPWO4lZPj/ssZbPVsCmONz/5j2Wpw+c5hAJWkCjFo
fTqENQwBaEZ3IUr0+mUeQD3jECOuQ4CtyiRPt1kTJp1ExnRZF5P7T573XIjx
Z5Tmf+UW0scP34leIrmpFncAIolK7L2pvknWM3XBcqZN5uTPyY0TX12/muPH
G5FG6AISFguZmwzNan5Fr0CWnXLu5DzVE/IX3z2uLXLs7m4SL2xZIlQDNq6C
dvQJHnJ2LhP/1JnVEowRblCsBnb4X3Cpu0KGpkPGWTphNLuai2/xc4U8xovX
9E+4Fl3plrwH2NRKbxvVGGFLtLRidwyuGeV1t4mHpvtFgf7omv+Br526n2Oc
X7LAByUUhKmTljV1ro74OBv+pWkQkzM7LQeNohLf3oIBp0T2QvLWSQmLC0ow
AA975xdbXYD6IL+7WhmN85dPlfpyLMt9WRENUyBH2KgqVXvxOg6Yko8Z2QsS
F2Q5pdq6M+qp/KU7QZ4ETMXk4D8rU7MMsJ1aSi1+87BdxkCLVbTQizDGoLxz
MSMmLc/24c0AT5MibpZ+dnswmcvysDzbirkkYbHfl6eHGJdxo0qRcE4AfLZz
xA5ActkFbzEQJRw0vgfzVXAd7rNSo+sGv/ZLvuK31++AnqONm5zJw+1mnFkt
HI+w4QH1smcf/aWeXy0ouHSdaNVOznuV/5DJv3dGlh7V0yrBqvBqvQKPu1BD
SxtP2U6dBwdAEEjU3b84FzZbuWgKldEr+CpRsmLglbG0f3/e+hKiQDi9Tfly
gNHQuZA5uT/2XdZ7qqQiqK4JSVFreyJnmT5VvTrSyPXegllFHN2pW/O4DJfY
dcWqI3vkjitHlDhS4aYFYnMjn70/a/BnlgY15XMTaVQB5Jvv71ipKD8IKdRl
fzyZSJy1JHdXFJKg6Q2Uy/RjvFqTzlnD7Wbh4NiVbFoCzrZ3dx7HdJyyihHb
rsDtzO7hOLcELr1+esNu2CkbWW5hbI4bq4NisSMEnJgT920K5QaaGlAzAkcn
hZLjUf5fhJLYeCxVCb0klTfCSyu5eHE0Yi6Gw8Q4C9wBsSQ9YqOTqRhLbg6T
dhDym2LWsVr4BI8mVP/2JB5ADmtz88EpMWJN4SDqQbNtXKZyAKege8tkINOE
SuFos5gJwUN0PojdnJ4VKWTqqC9GRAmy1Fu5DLXOqE24p1KKubTLSWDAJQN1
Nqb1/CVMYZ8qKEVNdYfYyDx0VyV10KUW/HeFuETrYmIJfby6am3TpGm+7419
0zk3ZP3aWL+22Ck+FMNV4hAvQB6mWiQW5YDbvxZzmsDTazIyxMRTuTxLaZqw
RcihEeVqP+iexmldEyaZjCECOUQddRbXPZ4WQ9XQ3AEJ0VyaynVivY+4QXAS
P9BQDaQigSUVMIE9P4mMHfSsyQYGAGpj2haVUPS02faZXMNFqqN52xSzoC/t
fHBlJ4BFRH8Pq6xR0Uv1twyKZW9TwrA7mgPYl7gOt8ypy+D++ywsHqo2jCH5
m6RvMaiBcT8IvRMT95jLqX+rOxaS5ZbsPj2K3IkBUmjVrWqnXLuoGnGvhlRP
ssl4y/cFGyg8lmHtIqVxRjvKNcO+p5amf4lS1Ntm7G1OKTMO9IChayU9C/1T
vcr9l4I95XZ5Jwqk/iLpiRMjWc88ryQnaLyEdsTy3cpYwFAEVuBck8wLDOoh
r9sf/wsr3XQFbAcSPak9B6Gh0gsrgeyWR5JWxzliG6yukliY1CAwtb2WNNv2
VQd+YfZRVEdO4vwHxe69/HHerdn7Hp803qQvFHzOTxMaO+yUAvKZlZ0t4t2L
6LW0ieAMoNQ0VgWFtDdVWBla6pM00aWF3t+YgTXmlETkSn1fmco/5wuCZ6q+
uvCkP2cN/O6jDfjzLUNhEXbXQrTlw14DSGhkqL/NjT5L1utDFUNsGlV4xR7g
B0RCIMgjlttTZqX9sJ6x7Ks5hCNQ974GuZJ1Iv5RG0X+BLmiIdNdm9g5AOSr
j1wlnt/JWerAZK1MTmuP4HUdChbd/BQhveGABq5qucv9ht2dz3EsE8eLfQKx
SiASNhCHqyby7DeuIlVYN8Suf2QpzZE2FswIMgp9j8ps/KL1WmvmmyLIu06F
jz2Xlib3C/2xIcA94A42S8fP11Lb5F34yX/pNFwOWpEPUPPgaO7t+f/81OJH
DN8lAl1hWP2rbgOPCYR20Ek1mEJ2kLusPYKMaLZQkyZjvnNm5cGXJWxWTCnQ
S7cJ6/1fefSQ7tvaSJCpNGITrJcfc6Of6IKL1zliMUrM/T1HNecCN8wlF9ag
2idlVtHu9B35ZC1Hup8kQmFfyGGlvy5g/VhrW9p1nN/dx+Qc6Ql2PUgZxXQO
NvV6VYwaxlSQEfRzePle2SC1DKg7rDX1jpMjehJ5K+8ByWqJRYej0pob6STn
F9nuCq4/q82Dc9IGGlmkB9gMYULvB2sd2D6sJYuCwoItHP5rO9NB9e+0B2q9
hMDmgTTDv9mpcqIwZ3qryaFBqQrVxhDwQr0oeTP+nyKfaeHglBMgVt95+sGz
dhSgxwq7pVGExlI4mvzv/MuyoNOaAsnBvqgi3OUJt1v0Q4MdJkXsikneRQhz
34ABTavK2fk1La0x6vpO2bdCORvbHPi80idG4HdqZQCUtXcj5v/GB1gvUlfQ
oV+mr8C2CBSTpMaItWLXmFLOUduaouYdIfQPSs2OoIfsvY4Om60EWNeaX8+2
Vki6MQhSbhk/0+X6EznSgEcavHEY5wWuSPs0kyRVIaAe5sOgsSokZO/zGklV
HeLuFYdyrwW7rer44kbrz4+vCqn6UEAkK4BCm1zz3dIPzCB/y9WKeWJn7s7M
hMFvFj6THMW/5yaEkJYvt4ndbcMPSiNd8Rei5XLGWFqCRM5S/zxEvj8eeV3K
HqSz7hB3mf3tw9w4qGzDqQi6I5XQB9BMdi17hguiOLb9bazYApXQEx1UGbSd
L0/BHtHmoKFTcu5JJWgQepZIcA/obtAS5x4jN0VT2FoP90Xpkv7m3MSTQ4w7
trf7HYE7tlA1JO4dlsU3voqkn+xGvvT3Er+1ajMdU0MMHqtAe0jr9EmRGLXF
IxVDj/D65g256GxrWAU7X7CduXdC+Z178fWtPf5SIMPNhXq2OOrJBqPUrAnR
Gi6OXtxK52u9z/1jMNR+L5uhoDNsbNPJnZYYpcZgiXj2Qrne80NHvq6/5Xbs
wZiSDeldGsIxDrtEK+TBOlLeva6vOz8rU7v2t0K2y8jC0hnC8chxLBx7j3ys
9klNjzuBVo2vuqWB07Dv5vArUxvMu5ZJBw3J5jFXwxzS3IDmiY2gqPoXDouy
OBXkqwqYTZaUHNWWEVYZj9E7fXwKTA572S068UP3BQ6Ej0iMbpIBTZU+Wi0x
64kcasUXK77DNdHu4/o3QTZJYaRwCZV9hoTXkYMfeo4c9PBpTmhub9ku5vFe
U05nwE2LoQpFLkJSGkqmcOo7Bxu3dd1PeUNAQ7F5i6cKMBAUU4IcTKOKT1eq
1kZnFdH5qBtfy2hPP+VX7bCktQmG2Sdv9tFnRnB0GzC7UoW7AfuiOoempXiW
zhBG38/PIa1uOpmBAnNFravUQ+Tps8ldTFX3o9Ea12W5oJbUmM3nLNjSgG/A
VZ0Ev5UnbMOFhUkc9B+/eh0L7fbXCRhxLdmFT/EDVneO8Sr3ZsUei2h995CU
dKgV0zKXfDsDtehAOwLJHMje8veTi9ZF4XDuGbeak8QSub1dFKXLP/E41Wk4
i387WUTp3myZoI2Pzn8TSo0iRHEwRY5ABMRWSOfpde69qQ2VAmoFeHeweBlP
s3F8wnj6gc1r6RbLQH4L0km4x2eAkRay3mi4z7hCWjfz7fpfP91ubh132FQY
xZKD3O7O2iXBI5vKzi7/uBalo2O6xDZB0Ob8YzkK2yHcwOHcjbBoxAKX4ewm
uGWeqXIfiY6MuCASu8Civ2mZfI5J8TbtWXihluxWqoyngmmx+HeedStWbF/o
VKcltrq8Y5Lk/7m+UxNTl9P0ZPfwueLUqhOB9F3MBEBQvD7ClXqxfwMBFxfw
ZnDf0G8mSbcuJz1HGwNYB/exOR0hFwKMy5z0njCychHhz0AaOdB4ooe+Al2t
5rS3ZgQKyWH3DKFUYmU9mGOWHSU1Gb/Gk5/p19NRddXKn+wKs4vVMBRrLS6p
kGhV0fYu2gfSOHNwRwxNHBqZ1En9c8uv3M02V8FJX3kybHqN1OsIhxaQ7o4Y
uO7VnNRJA84ZmXV/CsOGAwyu8geTJtcHANmJM0b64/FnqLgPAu/VmfYPyl7h
Upqn4d4GGHpOOvu92pJGSGbHHTk24Lsbq0JatMSR+VEvRaAcEARerpn0dZNW
w0d7Ag0ua6zT8WA4iOzr7CdoG/JnoB71apTUAMR5Sx3XM2boocyzxspUMW5H
46mgJ5KS05vVcl+sDrY+JKoY8EzQOhWzbU0ChwKGXErvH2pt3vU3QYkRyUuQ
mtdqhsZLeTQMXA8GaKua/a6kycrRU2TkZV2zzew2uIbAPJglq73dNvAsO4JX
aU3igKdDknYjplbOmkh6vBqva3uisfWfCVAOwE0XrTS9ddUhiF80SnnnUlih
jBjrbCtY1JgC4f5+W2HRT1bj8Br+RZOu0yXCHmR8Xrruhmo9x9fAAvsGni1u
vqsrdH3tRsHYkq9nKK2E+9ZroB+hoKT/uaNUFy8oWV07NY8flb2pfWw2TwRT
6pdeKmWAwX4xtTcV46AhcW5AD7nPNw4yQ7VPMbxYVL4CjrDhUfZcF8qHeEUg
Y3/gIszKuo0NGkT9+3GXte9IrgybvQn2gpiihzHtBGzco86KALNXWMDZTs3v
43PYeOQpGwJbJFOa6Dy79U5GjiW5Xok4TRN3QbfhbJglZcCKqYE4+rjQxv63
W6YhMHI23wbKCpWrMnk/cge+B+soiztD0CrBUETwHsy8o+PRYM4+ZNrQYaYS
lza4jpMGicx0JTpz5gnyBPvP6PQcxEOpX6BLyi1Vvqe+ixORPnYXIGXUUa5N
aFQQeyzCXr0OuiqJ5za3+44wgv5hsVp9OVIFPIKIRgqmqQ3VHVzBOvMX/Smn
hWsqhB5n9cgYN6f0EcUV79416HBI7UMMoXHQKIrU03koGf+LI7/HifLNtAJU
9vl8UO9aXDGO34xwYso5H+PCrPLQZ2POCRsLfH+cbP3fx9b004NZLrKYve5a
1Bvvv7p8+2/pXT2857yewaNlMqaTGmkY9gC+cskvTun49uI3AC8E0DW0VW6i
YAxtWcXEbEa6gTPaGdmLqhGZYKi56oYTdIGCxDPpHPPF2Gl+ixtOvJZ9bW98
xqB06jfirn0OlcqEPR/10NCS1wY6cGSdJlNyv4pdleZu/KYKHfHkJtxzFTr+
fcFRn2UmwwkOsRds3AWarQ+HWz/XcY3cpxAkvMpF0a+SmqpkRkzl0iQxndZ8
GR9jFc1E9a9T5aXKKl+tvWUWQCEK0qoID/ALBRLbA0zNrT5anCTlhJzRLrIb
oCdm6sigSaMlVg7Pgy6H7+nkR7BthQAD1N6SRCXszHf6Jf9CPP0HXdlWQY8C
G+CxZC6YAUAwD68j5zBe9NHfhpzasHf3npN3TkKzhlbfCEoXfPWuUo52GF2B
2YzZysiWxOj0Sl5zaqj6bKMJSbWHvby/V2A2JR0v1iFLmOjKEufqCcrtNBpS
MnA9OUwo2JxCL4VeflJULKXSSZVnYVc5ZuYJcAP2cOspYcy1W0avvJkXKqLd
882+Yp2FKSg5rwoD4BC8EAbjBGnqlc0iIeeng5TmgQHxP1ZWVTBgIqcUzj+e
QDE94wEPzjbhYDzEBN0G05ToUwpbTnX6RIgJNDu1rOuYJd/IDHB0/ueQtdvN
8efNRZWrrF95W5B3OskM2f4lB5DqMZ6xIpmaH3A0xEcNPAqPQZmcgLGaRKtL
pwS6MVYkSjNLgzWTJLolkb2Mo3a+3faQyoOuLH7lB5asM/a6tPzZvsacqmhO
TRpiFXYuqdPEF3Rp7l8g1Q+xGK6rCrsjBS/wQhfKJAdblQXXAUkKQQf5QgYl
01LUEE76toSlgAucoN+rOX+yscTj1iPwkeYk2riabRn9EirkNAyyRgUJ1riw
NA2rajOib2XPFKwriileJ1eIvftLsxMo7AEiRKeKndOVTbyLOMIz1X8hKAWQ
3OljuWxn81KOUt3WS+5g7XsUEgG9aM4VMXiQskIeZyYmT+41BrL23FZayBuS
+DZBxzDgqx7YSD0K7u2ZwjMJdFQ551VbmPLdQ5heDzyATZV2vWOaP5AZkp7f
A8xjoG+cjtWsOowV5PsxsXP0KGWPsA0J4kqjzBH0uUGBx2+SVD+uWYl39Fi7
OC7vA+oQkeT4Tifk+ff04OD49wxMyd4fmou5nnMr3a45unqlyfdWoADMk4jN
Q8gwzv6r5jX3OV9mqX5+kCQu76lZkVd3dDW9yv6DKeBGev8XVN5GgERbf0cc
sq43m6OR0Uj4ShhW/IBC5OjF7i6qY76ku3RxXCIh9HnE4G9gIVuadCIoO96K
dqFVdDM4izzZzNtm/TTH1bpNFGUC9DE7kFPfZVMai/JUlymILP1FAiF7fYV0
wyl5ZtX8aHkoEKYc4ML+PAWK7Ef53wZcCLIREki0zOmr0kzNOy+1ZpiuPa1H
KxHCshckCN6HM9hFubjrvdowfBXMcM8SCn/26YS0aW/V9Q6dZz9rYc4vz7Hh
NSfmc4J+jXVJNbczXUXYDWLqbixbiW3ilmNe3g002VlCJgQPy6Km1r9cCr+y
HcqpLQYKa9k2hsqkJTBMda76A/dcjrqruqw2nGtt264+bLLpIBxD8lfBcByi
dSvkzfm7L2gXGjUU9+Zw6NgEYuZQKQ02sVx3iSho5gYLACB7ssz34V3Nj8Qn
QvJIA9WJ8VKiY4kZvBM2nZyTCppzk/NKfFlKXnoPgl1+DYdQEInAIki1zKEo
fJCZ121OY8uKt89toNTaX0rdC7jLJVuvXuOBo8tSO7cKoclnTr2MC13z7l/T
ktkEedFELtdq7GNsLM/ULPlQkFQb6ot/Gwh3fgLHt1fHr0gLmtSRZrR2Ji/E
jHNUsOUgCngdJzK36YcSdGjZ1Av35isKDwXQKTEFJpexcK86a2lW71wl1ct7
Ol8A75QycbS1ovz8mXaDOTSuth0LzBeKDPzjHa4VSLDa4+esx+oStORM9lgv
VeUS1RNYRFndI4D/4pYo1dT7RceJOrUpUeGpBZLVMQWn/y6ESZafxRxqVX5o
rVwTwdySq2Leexr+ctJRe50pfAf/X2qD8jkxHUDKvw7Lr0fc9lsnezjcp/ih
4dPN44ms6bZTiyqFssBAEqSgRw1ChdD48c7/KwMS9D1P0u8bxkwMzFPNBz2B
sJODCFrjjCEnif+BHQEqHnTKEXQeHhUKsqIQ8/o5mGctQ7GBm4JnTKmcnByF
EM5w+0hvJw1mrMCeX29etdXwFDDPHxJ7f7DaIevEgqr5mqMwR0CeOO8Wmqsb
ArPVmcXO9SMRF8JDyrJqvn6TWa6JBpGdVvMhTntpxISU+zPr8Vov755Pg9JF
jUe6zAC2+hARyg1wPYtJ3C/muXahFmbPgtZQ86a6txVfwYZRQFNtcpZchbFm
0JCwyTB+yx+5tQjhuWMJFUeuMnlEp0q60HaKgJQmAm3RDECWijLRBxWSqdnP
JhJvBaBAUEfR3dYkVjnkmPNqWq75UhRTw6deviPrqPkUDYSGZFZJcSg4bRhH
PmO4bBZ7DeKtKPT2Rnup5+7y0Ox0vIqRF9scd9BLNlc77eir61k5WVnyXKcM
NDQkXQY9/w1ySJ5guSdikoQg/zrrXvrQihARH2lYqMb8Pvnzy0cLa3ExyVUf
dcb4gN0+uGu4BVfOTP6uQYfHhTJjQYb2qz6hv5pWE7EeMNPMkeYopoega71K
3/PXL90j2pJTcXAI1PcNBQdeLmQh4EOSu+T9uUbej56u9R7tDp6hieXIWFC4
JzLCCcFcuhhdmsQafNIsLOUUbJ5Rcbxp2CSuuFd0lGTucDZGoguh3p2HHZgg
L076ry96z/tjHZUvt+QLgaOvvXgsT6n9mM/GVkMzoBZ83mSM9ZkKFxxTcBOc
vSGSlFFHHNOejklg3A83xUWRL9QkztffoAzsoQAklLTISwhPBbOx4whQvjxH
aw3XlkKA9yvq7k9KIZVtxwK3U8skytT/fIrtIrcBMxEbADJj2toX+AtotElO
4dC3NIvgelylugojnoOFpjN3vpiGcGkkTIhIbvk4qVdvDJRDM9XUbwnaxeKe
ZAN2X2/NwsyvuvkbcpMIMl7XCcxymFGtm5cPRl5vV/z4LUFgqhT/LudDYu8x
2rP9qFuAIsqYlcqWSfXyYT87QyrvLb8pkCi1e69vfUHaoCZN+MHMHA/9b1H8
XqZH1YVqTGseM1XXcCugsaNcktoSkbawOih4enzP1e+jOx3zT1xCy34jbZ3f
I/eWLYriLJ1rIDWJPS/ghCYF+rBZqZyiY1heMDMtFvCtrip9Gzd4KYclYJXy
AQbfvilkpa0xn0pQqpIxNViyG5VKKBobTjDL7rzrJtiXZajI/zjLKMfW8wnu
D/yFfyj3+UCGr34WNUo2jxu6TJ3iHUssDNFgpO0b1vARgoJuvyypcqDc967K
/lAy4MgVdrhELohNPUZjuBRTBWkLp3tvmAFCG6mCXKa63DEOYE9SpnhGM/Wz
AvbEKl6do3G7PLcyz8qoH89a+P+QQvoyUt4zNzxzzkYiQ5ncxu/vwu63DMqN
i2HCUZAQse6+dE2T4UB8BeJzcBc+JHTWTXVjGIsUOUToX15AZ6LHQhXbkxAK
PJCUwAsufFe7NKc5oyK3ejARVg+UVkzFxjewTll4gHMCDlOtBDkf3+QvJmA2
9LGyP0cz6nP0048DR18qKIhRjbTuuHu9qqoT5ZlZNTBYfgrAAjeh9T6KEozy
/rziP5OYIeZtYQJTPIn1moZCPZtEfcn4zSgb+TB8pI8kJp0IL0C0xmwkgVBQ
wQjuE5oQ0lmKx736gYKwZGAc2L2cLNGX/pA78TY821HqzCdLy74mFTX9+q+s
w2yBPlAJZ3j7Pnp+TozkkwSiWDIj8JrnpJkDer0XsiMvDFND8PwqrceRd5WA
UhI55XIwFbOFphmNdrzHt7rk3NW77j1MGcpj6r7VJ0X3vgBsN8OelEvpAwfQ
4tk/6mWKgVePHWqBw8MlHQuA+QlbMQTnFgStkx+9SgmaBqrmPuoJfO6soUI3
zN+N2hEE/Kon+k3N264QpXnm1gCGP0bNJ8UXnO5ME+fSOdOsaN3LO5B9vVnf
C0VYInDKTiosPmRwOEtSDsJzpd+zGpAV+w2NfRJYDCIH2w+jnA8gdPn0/dCU
NzPjg8nNL+xNXihDGjHuIFxyTM3tEauFzvxinFv4XYBD+PkGTNHLl1AEwzZw
/6yQwCQl9LEs11LZEdtki8emBJZEz6xzzQnLRxQ/OKhirVtAFAnCcdj3h3Vx
SJFmzY05Ai1vh/uExZQDb+3MmBSeyQ9maUOspeUQgIAalWVAoAxT5G3r7YzF
xwv3bbkTE4/bcq5+i9kKvSqWLa/vwLt+ONJjS+cyeahLo8pNCgjJN7Q0FZgN
hyT+eTntX0XWhrBbHe/8EyDgYzdbBl3bKtTQYR7ual6uBIith7WyryeM8jcB
zJgSCAsUjStI9T5YHWK5y5o/V4vSzbQhz1q9T/+2GEeXf4hwM3bY4DvH9Fpo
P4ZTQmQf1ft6v1SuqsWIA/xfEcaPzJJKh4M7JzIaRnsos4/ACkZbHzisq55X
Gq26S1gBAodB68ggU79ZH/7WsK5SLnbdcCLzDERJ9oiZOi6ge2S/j+p4cFL8
26iYMcZGVprxDXdGCGIgClU7BhzWdzXBhwdYGwuQK+yZuhQhYMMlRhzRT0Bk
TAAWOZtKINud0e2SWjln7Li6Vu5TWMnzlqlbpG6LBGSccyk77LaWriOd0q2q
IMaSqLtxxMZgKoLFbvd9UFz3bVZ8NGc95KN72VLazHk61MYurPBy8JbbQntZ
IZvnb2ukglUfUhBBV7D06aLoUt5W8o/SxGadG5OYT1xJHY0d6eeOLYtU5yQN
KSA31mLQq04w5yhYJ/x5i3izBj/PFb3V4m+kV1Z/M/BMXUSEtE8g9yFA758a
f0GWq5A93HRyjkBPki2iZD4trC6Npj59BFUNoCZBXKcsOWmoHCgqX84RnTF4
5DDoCyAUEOu5GC10xyNw8SRxaNJH8d//zY0if3iM/jY2IcW2cpVljEfzqtVF
IpuroK7gXes7K9r5l8VRO3XlBIDdJfmeQs+LaAmco4Qqa4wQsjwWVqmf52A9
RwXPouiqdSaC8p+6AOdIndWcDFl532OMsb0OD7nElWNeZZBAlPtLocukZAfc
n7Cj64Qq4bylHwPM/N3rKCDRm+K602DoLL11ZWpJJapYMMIrL0mdMqlHDvsV
0hjAuzMayaTw9s/qZ3vrHl6F+eS/a+5tb3snDGQJhH52aCMznWswNPlw5LNW
zzidAwkSjvHU0DauclAM9Ua9QnAbiyiXodDRi7OSc+I8JkFbqnC5B8KRMbUU
fJRbh8K+wKTNb9G83w2GjgYuKqw6E3ukzNEUe+/5AQPSGTQFIPb6j9BHX+66
roS+ByPumjyL6mF3Xk/ksNwqR+pPxkcWGuqhkBca/ihbODLKdE3/5S9pHv+l
OjgV6L3ez2ged4xF91SH19X+DveUaxZOk2ndmXH2wveLxKZtYiy334URP5qP
lQNBK0xA8JhRTgOH16iqkH7/opPahp+ScSmZ2Eb/wteJ9upk+1DoZVDTkSfn
IYXHDt6PAfx5ZfOgQAL4lYftrns8543PzlT6p2xlNehZAuX5TFaEpuWnLrkH
ZBeGbQy8PsMYSb2TVf+uTQINk4+TzXIyy6t+vnbGJw0zdPWhdNaP8JNvUUJ9
M7OMtOTU7Zyct3we03l/n5V+aaYhKaEu56WXE66R1Zya0f9UOxbY5J/k66Cw
DKi2hHWnaFjMD343iMSLg6XkO8A+BGSwHFyzH3nRNpjR1F0HJNGXvvMFhSjV
sYiIy9oPG2vvGsMbH56R0Gn8b7TocdnLKwLl7MuToiFisLJ6EpQgGpQHDUW6
uxCrPVwilmTz2t1zQqWq7YJbgALjDb3nkjuwgLA4syl2lt6dInfRhHXbR3wr
li3xS1GfEcpEq7dDOIeIuuiQwWdTLK0CotT1gzXMBheELJ3Nv7uAzFCCk6TC
cAAn22CTj79KMakb0tlUHKVypnXM6KL2iPog0/7/tU2dn+yi4OlXtNNU0Tre
ZmuBpivbl38aQFM89JaEZb7F/wWR3XME653DpM7WXGGYMCWzIIBELans4HKE
Wq3Kv1PKNf/ZRBfRytte3VkGOyqXgNLiXk1SAe+bCN15EG7ygIesdEGh41ef
3dqnpi9It/H+2w6VA1y2WIDNZiAGiFeOTuHUx53bVYg0VdvBRifm+bLuKOD2
8v05SqUvsOYFMHOLQQpsLzJr8daMSB54Aqi9eZrINB1kTBls2HeO8IiAV1Ni
GS0O8XZW/ewXBZcMVyNbSvv3J8QDGXvGViVV0wMMumfD4d+lni1DCKTMCJhV
nXyRbYZTq26rmbmW0/uAedZ/Hckhf2rHjmhlD9IxzMsrsvSfMO1d8qif6nyM
9LoPXOCyJxkXt77z1JoV/sYO4vOkRPmdQvFTTSxwBLC6qDrijxzSsn35W7lh
iAO06oo/4I2uFG4JxKcbxEcdJb1pA2cmiPil5OfpXuAZl8O/a2v4GLf/2+UT
NtAJ4l1sErgMZ19JFOxbh67PQNB9KT45LE2uGhXzCxnOulTJEUGlGS7xq/Qz
57qRURyh/uq8rpWruT7BUwYWgiUOK2hsiDy6+PLu4a3jxTFPLcoQKJENRA74
xe5/WYDNYwgwiKzxmKx/BeiFMcXH6O+sZiy0TAsN0iH5hBcnvnrMY8NOlNjL
wtbFPDYkI2f015yjptUQKPBXr+Z4xYRnBhwzzVXPv8SlNOlfcyo3aIp469a9
gL6C7ZuhWuwW6WDCVXwlwXQqcLa+EN3lmMfFRUNXeqkXg0RbZdsQN+uenrG1
PMLAYQZUz2gIMf6AGaJJuV1XgqM+LnzhxDWDza73ttFHgd9PPkE+sLlNSDI/
DKKBf0k5tGytMV/foEMyfqchZSAgSJXhACZGrlu74QniHddAA5sHj/qm0EcN
ayf4fp0ihRW7OmWObR8l+z4NzZQenwQL1XBSN8122RpP5vrwrbk6mLkSl9fb
1tsWk6oUK1F029c8ibB5tB8gv23qivhNpc6wFC+nqPJBCvIpATpEfduyhy5N
8pHR9qZPCuebbvK2DR6yyEhgmScZpaQjnD3nEMb+uHfn1MpM8winBVMB0GKj
LVCjtieXT038Wp/YJFEhYeZqG/TTkBb6B6jkZsfE9C6GszIUa96/yhyCNDxS
LFSMkq3xojZLyqsSBdwS7YtGjkj/GvifWJ8NiUI3fanzJycFQHuta6HSS1dg
az42b5IxTNfB99PS94CBsG1JynvQ47DUJrpEhcYrOrqjkcjlQUaoP2f3pY7+
ksDLVa95QdNP42IBHDKoo/HmXjyxeYJUEanaKJqyjwTiTtI53k7/5XaUZwt1
5SFfMKLKEk9+ae6EJ69y28U4EgGiB5XW9W8Y5YQIF7KDjmfZISBteBzVzp2e
7V+7IoxrR7adehqt1W6WpvchqXOVNADGs1mT3CBkHNKcvLy7sZq41apzIWWc
prr3Zdfl5aWf8T5VuzPUC6GryWzFCmEFvG7iOm9USEcy2SbIodd+z9Y7GQgE
QoXP6t0IZABlaBVQxHwvcaJ/4kRPSc0kZbIEp4fJQB116M9/GE0Gh4aN2HIX
9HxhieOiO1wBdE+L+C7sm25w+4cnThL8uCkraY7bXYqE52YIGcqfEbyv17sC
PN3CeaCntC6WcT57bf5WV9EtEkbYC002dTPmQ9KwWTKhfwfeSLTACnxn6nQJ
UKBP5QO4z5l4wZfc3AnYdl6muE7ajLYh38GnF3us8p4UfSA+bZCMdQ3knaeM
fN4SVfWGuSc83Rz9uFfNw+bR7mXBj8x6Uz+GzNZlSS98kTtVwRyU84yNpNQ4
myRa1DpIscWmTsMQphK3fRDR6wBuQJFE73zCxZ861ZQwHnQXaRv6zLYamZHd
zt/rmfi1WdB7gpOTWC7JYkE89sXc/U0uwVV1M0SFGwzrubhaK9x2/noUidGb
5vno2kAECDOl+Z/JorCyKtX5gXXEyrSFw7//xjOST4tTqRBX+hnYSJ4Uope3
DOA8OxkWIilwhrezenM0dMscL2YaBxn/cC8nAG5Ri8EXg5QpNg82QLXQyT3W
qUQiy92NMJ4vNvmU42dqwmUJ6Mx3z9AqHMoBg0enH/8RW8uIZrG9PZNG95VH
izU7EVZ+2NDaTV0E9wSkaY2hjEiEQICtjVsxWQYPSy4wDTR5dwStzOGn5C78
OJRNyYsIxA/T2H4lQCDdM6wz7LGC2V3HU/vW4+JaCvBD9tK9CkdoVcQ49Bmn
OzVcbqZA4IXD5UMWe2IxAPHh4tl+v5JsTFkBT1b1dvV2zXdxLm3sMCm9gnzo
XrnAvAZlndMblu+NsR8FMvzEzOByD4SKGeXIR1KnPSKDvzyl1r9zK9+Ct2/u
08NSi+mCrF6eXziCAAALqGY+PlvSj8v04mPtjsrMOZV1kSqhTyPgiGa5M4Ny
asEiJEpvSlgWvg9wqDcUrNOjamrqvyS4boLb9e/iluvdXQESFwzqeKKfGLxW
E0J2H8v48VNI8bAP3fvlGlTcEy2exUDajkAoUYIrY07htuH7wvqDgKeteTXQ
jEqud7ca5mZPIKkdjbNFOqicQbLc2RC9b2p5GxwitALx4qspF2vSk+cFhtQ7
ZNTLcYUZ+83haTid+D+zTvFpnLlBA8Cp3g1ikOmx9ej/wLqOo+KNbjvr3qm7
UevdRk8XvjOuf+C0toOG+cj1AvCZr9DETZtt3rw7rRAkXwizcKjrsWqz+AT9
BTz8HtfV/Isn3/w+snVGe6M+AS8e8JtvQf1win0pTtRnUAJrUyuV2NCge6Wg
vOxrRdfJk6tU/ZdE2f53sGo8rG1qnnEAnrVYYL+kujsojjtd+6Qcue+VcgkK
yyV6k57SaUCRpjDZroLdSNYBBhPgzMzYwc6e2lgQAuH6NYCvPuCHXOgXXvoS
PIw7D1BXI13uN/+6LbqWDFcWZr+bsqnNYuYKZkPyRLDb04ENTKXYXoQtAq9S
1OcFyShgzeXAK8kgq9jNPlobCsphKEG61hOQcsT+PRU3X/xSJkuLACE/DQTT
pGe3nVBHRnzKW83wvWDHbrGa3bVzsHLXt2LUGLKpc3jlHIrK1x9FCGAvMGwu
oCZXxpgHEs4UPzuNR0bEjMkz5QpvpDRLrfqXiaklmoYrZopRE79kpYZx321B
PJjrK2EDSiNgYz0G749+m7du+t1Hmuj1r8SvRWNTUai/hQI3TDMxBccYbxZc
g2bpSlJ6PGxsxUJMgzDTmGTikGSQJvOumwo1L48A2TojLqwLdHMPf190pPW+
btIOaMs9fkQleq1vjxpIJ27V9o9Z8Wr6vIqCwsrl73uyNFDo26M7GG11wMeJ
NltNPNt98v1vK+SP3ceRMGrZEFtsgS1IEM2fPpqHr9QoFEhDjMUuFrU8HjTk
BYzP2uttPe23u49WqZjhZHoqxR71UtVs5l1LDN30YqUOwLQndykJi090/QA2
e2s5uqMfBfWsveuFiO8M7HSKR48Yosjz8O3xHKEFHAkyYGgMo3BHYTiQ7pOd
izCxSLuz6eyvmBpHp0L+YGcUgJx5zSKg6NE/tRNiDVB4hT2B5NsfCeANIG3x
oEXVIfM2ggTTnNlRBuRHX1sCp0//c+bPYwW0UuYqFAxeE8rYGypXFzbM15D8
WtQhrx1HDwwAWBJNl8uII9wY2vZ74V69+1z1X/kJvPRWHMauBXUV3Q52Hew8
dWC2B47r16hWLOyOP/XPs5rdZGCD2bZxcPmnNPZns7rOmuMGo7L4AeBw6Q0f
nP1SvwXjdTD06Xb/oiS5fd8PpEUeYTzAtTW7GH/XBC1a/LO/bFUZiq6zwFlm
wDXiA2jnT3ZEXP3uy4H0HqmpHcdNtT0QRXPW7M9Jdt/xZs25ziNbh5rlz4zn
raAHrRfZ2PPv5BRWUSTdkFqHJtJ1+2BjC9HGqGwye1UkCuIBYZ+be2TirMFg
qtB//+ohxzdFv4lSIujFTy/bjEfzYyegwN5gx7smoOE+WCIO0rhT/WYwiAhu
mxxOEvoWVEG5QMVUVzjaZU2XgqFfoKn/+hyXeefpFfqnBBOw2VuDcUA5bUXZ
HgCTio6c7dH9R3Er7W9hMta00hlbbjPbNPtFzBUi+Q4osM7Atp39CuGJu2WR
6N2YvFtcBNWqFpSRYed/Cx1LhvQPp7kORo15kh/xglzzNpuzhdiLueIilgmH
znjvnSQZfp330SJ7R5ciZQoN0tEHdkat8usLuErzX//INtxZfrY4DxShxidT
chQ+dTgl144ozcsib/yYFA5NEpKMgT0/zPWIIoNRXe0Dc9HusxYj8B8OSoYU
9RxPqowsfFDYlTp8+ShhakgnXqb7tPvg4omCTRxQCLJYBTfNBojNHqZqVYoQ
wY8U3LSGunJY/3QihkibewH+xCjgNuizgKL2zUJVaQifQzOj8o8xJLeUlUx5
VGkRgBaHC9FSHsihIGUgbVS2J28SBX22/tgnbbTzwUvlXdxRj6jotP0TOGkx
AyTg9UqkvLcq3YDJmC8R0SNfe1xp33wg4LFALHcmQ+dmDnTW4kW4FQpWUWjU
BJcvRWzsMijuw7Ts9EBoqNf7q1CDn17RezV4PSsBAV5f3wUsD4G+wi33RGD7
+TgJhPJfahTCVrKm0fLkr6vcvYW9JPYKN7eAeqHUbmNwR2FlYiE1G/dXcTZa
Sm5FCLL2Ag2kH0h+a0eesuyH6/wkHpxgmCOiq6MUnzOe9DqrdowS+biAkJLt
ameavMv7WXxQPFQ9blceo/CdD2UYtlY3FkCyKlZxnad+T95zOFwugAExYH76
T8dS5XAhp88SmF5Uu8lPay+KXthBPmNkaJeXW1snBcnDyJjnPo24HTZVR+SG
MSVAdVVgHEBh+JKCqczq3UGjIhGnIVpdPqIc5Sj6QVZ83HeUwTmh3tI5qtHE
qC0YTstop0bFIWi5/6ABQymTrv1i0yWLnLvTC4Wmv4OfNfj+GG1tO8A+Jymc
ou0ONPFw8mGlr1FHXPfPGgy4t1kivMvoLPYcOgpH/gwj+ZMDxid+iF7pnXaG
VrDVHVDznmFzj4NJOEzEnjPCv8OARujjxPb8JOF2RDEKne8BoujvElJF+5nQ
8YHJmdvzZvKZ+gPw4TCnkxLZfJZ5ZahD1W1zfuMYrsS2VQO9dBylfJgT6zsE
NP2oPsDQKyElDySoeQIV4yRpDt96pEPbDmWkO7matEQGZdnCOgWNLym6rw98
Mji5ctNLmOMZclFDMfdptDO1Yy5tU6bzwrTZpWJpnhyk3cbToaiUbPVU+BBE
qXQEyc2sN3FLJHaeVoBFhDmyNoSLKE89mYnU8qylBhQDo4iwzU1HSuaNR4WR
kf5qGcERNefLz+EkKezLVK07P3tp2rXHj/0PS1/gjn08HwErOyGfNXpmn4Ob
fPjRFQYfdTbvKRSLD/q/AtGL6i/uF2cR8ky5SsYlvO7Dqxx6EZJL8jnrw7gf
83jn9p8ZiJMxWFIs6xnPC3rquU+KWSU54yJulRuzfH2nROGNkEVk6j/pPef+
fqteSPsDTPWlRqvGmRUs8CPoPXwOjH6IEu/i7DBvzCfUQpjy/E7jerXDRyKs
L2qJx5WmrZxaZVmhE+2GzoZ+DT+1wfM77GavucDDn3BT06ETx+omwQr6d950
poVvCU5MaG7gSgCVnAaRUvdyazOGMO2UGAm4LsLVx+7jkcue+aeccqkVhIng
H6A5Ob1rSDDV5svi1D0X49QTqUtTEUv2rzLsyU0iHEnFmD308al8qmKpySkB
FlfRSFVV5IXCPygMpD7oG1YzlgyvmgzdMS+YVsg83usJfeNkS4hwSCn6xKuH
Oe6sQ0Mq772QOH4shvBC2P4mefP11SMnV/zv5IqDJNKVDUNaf/9TQ7N/slWi
ZjrTs5Loa2+S0FfPrR/NsAllOH5b2pD6/yV0eT/nug66a4jTDb3BwDJqtr8P
J2yNTQCjpSE6kR+deMWL+8VQnP4Kf1YraQ0PusGALBB9sC7Hv996PoWdYYci
6TQRdpMY8o1sEa4JRaA/viE2lBvN9S0gb0Nx+asrMM5a46mLw9QlWlQfHuH1
KM5Mz/8wNn5Q66y8tltLzE004LHQc1Ag2lldHd/8t8K/vZcJQVAjiuuEzctm
AF3WXkXlu63zI8lmdkXHHEt5QlLY85g8iYc8l6Cmz3ARyO3qwDHSZiD49xkB
Mi5T0lhAdH8I8oloJ2QuWVV+NiT6TEjregCPCdsHNp4TM0JaXu1DNvaloXHH
5rwatF9mEfJ896LG8QOQf/LDlGfALjXhFQ6o6gB5h5XLfC2hQWwM95FF+Pln
sIhPhcLAT+Tokirn22Ld5kNLlpENxQc9cFjYtfmd26lDPFE25KvvAqtOm5G+
cEH0ghOatTLFmkOFgw2wHjrW7c5Nx4Cfz3h9yF6JuLkDG6tbJFRVgBNFiaYl
6pf0oq6QqoUa8AnXuMyyUatz6o3cu88yoUTtqdhkBY4hXnaCpq//n1+F7gGo
JM/6ssLNwP52QlxW0LmF7owtFJn6cmO+2b9mmwwJWAQzrg8bAQufEFIagqJR
krFJL7298yxrZF14IjnJaIOCyzTQrLPleXUeph9x8Qc2Mb/LIJg/WymAoYZY
aRpJgajxRS6SbAmU17x0dJaHuWRRdtZ3+ciEjoVB2OWlVNVKJt/EqPTCekfK
j6QjMhUAbaT18j5HeADKNQk8VJYmnMJ8jCw66b/Ss/8chFsozhReWexc4d6n
rPN/aIF9KYFXZSdZccOuDP3vd+/7yKA4gF2IBfjmMARyKUtq7NQHI+Kja54b
PCvP/i096JjQJpdqGZqsMNbiTGIXldJV5zHJw7bXK56abChx39aWKOk3N0Z+
j0x9KZBX+IyVQE24VnMvDD2J6MGWnd+vLm+IHHRNOlx+143xdTsYNh5foeLS
6xQEW+3S6l9F0LzCdpHOfwUKC7yNZile1EU/T2Pn9gGD2e/hhHcuf18r7NP/
rKHh2PgcVsvsomr/oNc/5Fb0KZ9M1JB8XO+HRa5ExV0pDWnztFgasfj++nxG
1a/HzH3EUZM0QdhaYf0+zdJ/ReQr3JslsHbF8AyxlKKd4x4KnXPIle/NtBjL
U6GYEUNm96eeyabsGZ4nS/HqvWhZwZ4bt7/X1l9YFisQAz17QexHhAxclv0W
gDNMjsIaIlTyQ9wvBvyDmo6OQTUcLqWFC/6OHpinCVzP63/XNPrIXwD7FXie
ge4M6DUFJE/l8JHSS/d0GOnbKllhq4QQM+mSkh1cIbad4O1B3UGdP7b6IyFR
gB3Xncx5T0/C+IV6fw4YVQr/avNRSeKAgKX4RAR6uCfUPd0exc4Wa3OvA9AF
+HzXlCTI6NTE5Vq+NVrg1vbk1VHXphsKKufYaBJcFeXfCvSWhV1zcHc7B7+b
f0Guw2SIinBzCfQ39B9XfqjNu66CrvkVxi23nuEd9JotLfKZK/KuS/BStCoQ
xy9ngwu7bZjm9xq4fffO5EdXVbMPklwsuBfQhzuNhlMv4sbdsoLe20KVYNnI
kXkCGpDcu/u1QvqQh10Ktrg9mLcWUStyQqIeymMy135lssUMic2eeNnFAEjc
g2a1pzd662y3my4xPCENpRnA6I7qLoklzBj5lqnWrlsjmfm4r0hQ7AbtXwb3
Q2QctiaoONHSFvRwLkj132ipVwZ6IbXF2AzyvStzvMY/7FKpAWszZnhmZYDK
Sozjod3b2O20f2VSuVPTk9crO+G/e+4Z23bvFzchF/HvHboMEyF9uL7AjYuj
K3AtAFd2OY795iQwmZeAAi6/P8nKxeJuytLM1JS3jgPn3TSDqVDxhar7VHlT
NbtT6nbEu3IomKZ+h4ky/xbuRgmDU9cJoeU8nHPj2T8voi13a0uI0Ik8PSCH
sEIRL1V36GYh6iJXpR1twSNrkNSh18rRLZS2I+GiRttwZJeJET3im2oKNvvq
O5MVEfTSgTcKpOU0gVUq/5hl0SM9yUhG9KSw5eFDEVU5m6j8zl3GL/DyvfP4
ldxsjuEAbRqMjYF14ilz6Tx3V1R0OI9kjI0xahA44wP6YcKavKw/NRBfbDbG
ca4Xst+FB5uK85iK6/FyDvdPO3SHCVTzE2F601rlhkF1rA2ax2+PuKdL5Aop
/mSoqwBnsy0OjBbztLx1tTKWsSDWFJCIiRKaybnD9yDSt1eQ1vc4bUA3ema9
56rYrtLBlKtFfC/DVio4Pj80Iwd8glUeGbkTm+0YHHfk25Cozy/jRHUMDdOZ
dVuPKRGn2LvEreWMXyonBLqjN8VB9sxofbPboozZ3VtOi6Oz6bmlDcfMWK1t
NKgbVqA6zzbJqlBvUaS+sqCKFHst+8I1Tb3YNtTc86xDPzESoNT6W6BlOM6+
XV6hkBlPRifOdTHk592mcWgOiGg=

`pragma protect end_protected
