// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
6tilW8nnkVHjiVAPn9/+AybJj2VhoPFe5EMFoSMcy1C1RhkPrwUeoIsW4PJsbmBp
5KDTZwCVI7Oj8ynzdl6i1eHLfCrtg6doqe1RP9UXGcPQ84nGZjcg+mFS1fnuFjhq
CFePkCQWWnoLnkVYps+Q97h84e+iOwHDexZFzlyEjamFTnM0QqiS6A==
//pragma protect end_key_block
//pragma protect digest_block
lh7M5TT3Tw4RiRl5zgW9ZeqbxKE=
//pragma protect end_digest_block
//pragma protect data_block
rHFr6FoI5seAc9rdIq6NGIpuKxK1gVV++H/NGx++58oA1ayQOQRLXmB7WrqayPkb
5R6+vt5xBGF8L2A+UwkqRHMSMMhpBBImq92ptGmCcQ8NiPwsiNVkJBFTCO6eMG8/
0AdFg84WxoYFWgxtpc4NPvzb3FdaK4GX7EZO2yi1IGJuLowGzW/TM88E28VZBkFy
Wb5IPvJb+GfFNQJiyuuHMavSnD8C7L6vZLrIDKKZp6XD3FzfKSuhA+xsuM0m7kCN
COLRb+UXKJuE93mV0F9f7UauUtTmj/ZYDihAMwaFPjfh5BRAmQG1hQ6FH8hfHX/0
U5aGdxnrrC+wJTucngGxD3YxTXhxLnfUQvNeEO+bfjaZK1ev6BINnaTu75xSQpjE
+G4ele0nXCmGamS9413OZ18AIz8gscnQ1gEUwT7wFDZ6u6fYCOebewdYEd7oN8/o
elEJE66DfOMdMIMzy/GxnDOBtBYdm76jMe7BFX0kg3sOVTxNdRBfNgNaqRJIyJvM
vF0Lq4USXlqIvmgnWG9262lMOdW67hUvR9HJ0h+AbmMJEOGunCV8kxGtfUjVYdNX
50KCVurxubE7gOfDIKVvvEQgxQki3NClr82JgFnefUY9lDs73/r4bVHav19Q/XPU
nxVhtbNbcVxQPUBLgZsMDf0M2Ld0kuJcQD08jlxKudN0h6q1yf3JqydSJK9UFcE3
UISkgEmpw8Ba/m2qaHcMwd0rrnH9Tog6RUaDKBSStbS5KvNC9dEmZDSC/8AOUzxu
g3XE3i1rSr2Wj3BJNEgD9XGI26yTMfBTNyiverEbPCyO/cCoHNfMwvHLyNRi5gFU
4HQEo4/nf45p5UB7uNQTPNYyYKCSk7/lXD2mQL9SjXM4k4Qp0Tp9obhwGfsDmPfh
BS8sGd/5K11o9SsU9k3vyH9r76kLgwZF9hCgScblPj701re2Iz2A3ZPnKp/ZLrxV
YAHysbqYvqC64IhW76OsttFkuvsHHSI5DRsQx6+S5xwGZeEI4UN68CEgv/OzK6iL
L32EbibA3Q723dR0KqvsezeJvt+5qPxYlYsXX43mgmgx1Nf3I7MesLukv+NhLBb2
tHhsRoGlRm+iub7qAwcjISseI5xcVj36aFwnUc3GmIzTCqRyNL1sX8JCbwnikIFz
xEIYbyj2owUND975t/4yGToGjl8NOMCSpK/fY52jRM/gvJCsim7thKXJYiryPFOs
A5QfI4Jhzs2g4Affiq8fIWoZGWYXfGo95Ux1Dk2kCM1RCGpicoeoQB6/T8/7lpjR
BiIXmBhug1xWfzGOKkQYpwM30XCqSXOwLgHMbbQ9IgvE9ZdqImskpplgFxRbby08
p6A4KB+kexG71/m03vyRlaeZ5wI41MAD3ogtTGMahIa0GEnnN6HB9lPF5uw5tVSn
4Hcr7krusQLQycdB9vVC3VWcrep9zYFySiOhDwpVxrl4pFoMKW6xSjvYpFcvs8bT
cNRf39/lt2AifjpHaGXWyGESfF74nwANHTv7O1W+aTWJTqjcdBNj1SU9Z5AVKQOX
5zZcD7HGwpF6qvX1I0xTC02XszzNdp+sbplVeBV102K1IkCXwrWDeH0dHaymLmLS
QqQS/IfG9jccCT1Wc0l6Q8j8YUMUWjm0AQBbYmZo117mzM21UZOOwJNueFHjIhaU
1MzhqCb7D2tLqInPOrjJvoOB1OASkVQqLPHlrYElDHYx266+XcbHWfryMKy5J2Yr
qBYFhSE++c8lmJf/I5cMMgL27AmzzW3myJcs/IBFN26EXOOrrHcI06RmCVLw2Pe4
b2h7YlwNP54JlAChCofQJw8Eldj0K6Oa0ceuE1ECMwktC5GV+5V5xiT2GFhcLa0O
32DK555xt1/x8AUpv3jhESb2W9siB7Pwf/U8QsEJ0iqcrZ5sPCPfr5/uZ8qPZQGz
h2ZoQ02qtWEDc3zloARxZZbo164jKkrwzZBh5ZjaQOgpbczXrYAAb+Rvnj+hmzau
iWfxc+s/Sn4ILSsGch7do5FaEMlEQ7PEMspmWX4ejPMa9ceEIGJHRpagJw9P+dz3
pDSIOHIgsOEzyQfdyAwwWejKXe6yEktJNBXbfxPvzfNMFiL02O1QSlueWvJcNsNZ
xDQsjLMApi1lD9QZmVH5FJ8wbvwkwmepnm6oh8KgUpYRThjN6TVjZ5S2CfIAN9xp
tE/rMbkAimlujqve77QeYR2m3o23VfHf5LeLrPwVZu917aMJ9W6Y3BzeF9ciIBI0
FIw+vhGn3FkqHZXQ7j3U5X8GW9GcehFGOssmJ2mpE4AXOktsGtpNkdZlTkC1WlCD
Ul5BHGYoFBQjtYacRMf/doCRc2staiA8rhnLeEpjHqyDGDXg2befVHRmzyQuLX0d
IsnKgPm58+aSdrtHafkmuv1JBA/RVAQ5U70eju/T2tZNFQTUmegDhBCkCz4FNpqr
C5d2YPwfFQzS07Ny8y377oUMSpDeHGJuOXNbjX9yZXjMq11ZZMU2HsE3UzOcZw8b
XU759RbrueWU+NYOWQN4/AzUz3zuff0WgrJhRoDf5V+QGBZlwubU/8z/AB/DvQYG
L+hynT5CP6P7zAvvE6nQp5PlJNsuzEuMRRxLG+GOYB2EtcNkdlFDh+89z1E7vlxn
rrYTzOtGaLsjzzNVnoOY+aOptM3Y8sEzkxzbHZuE3FbMUAON+Fv+pha9N4lspqXt
IOVfmSL3U30Q21Ocb7ckVzaJdd8aS8CX1yc+rj5Cgmgznxv03E6f3YV5UXpczYSr
iFDY+22cYr1Yyqm0ptpDpP2c8J59oQ44PaFeVM6ZZvall+O2l7pdVoFnZkJYyjnL
pte7Bxjyy+PhvLHDUh1wA0+LGbMOApqCBx78m7fhI4Em66zBW8hG5ZPWWkxAN5bY
qCDFnXgla3xYpON+mJuaQJGINE3lNreFfUfr+p950Sgc3YsHZdLgpKGBXfu1hwjw
2D40NWXKg2fsF9A1s6JM4g1xf6Wpk+0FBqhQ5DSZJn5I+kXtzwTypjs0r54PSP1U
lt06PogaN9A70+wQXdXrDVpeOA9sOi3aR0IklcLUAgcQMl+5Btshija326tdgHcA
HLwvqPN8uncL9sVRTUh14ghrKwivRpapXqwgGAgMzuzPek9GE3W0LfiopLoVNsJj
PGvSRnEmO2KjGZXEdKdggqggCRzN5rN4X3bivFQf8jaUc4QLtQg6oD0ZFtgwvOXk
AEp7AksIkUmafdFm3RIoHrAfHqxegZ9wyY5xvkX/j6+PjCUBeqSRHXxPNRGnzGXd
6Zw3iAP6M+S5JjwD09oQqu+nSBWc26H4fwg+pW4gDQCJ+w/C+sRTtyXQEPabDkkc
9f1cxdDlKbkTdLSrxySEiIVCQMvTC+MwOvTKOd5xGKwlj8J+X9HYEB2QDt4cwcDi
+LA71OYttsjnbm90XKqVsOdueP8bUASlRaYyE+2PSVoOWGgbWALRu41ysRZ1czWX
yO71P36gYR9csstZA2JWt/Q+QUs/E/odQmlq2eWczaRPocxGmR95UdzcYh845PiT
rA/kt3iwM+DiID2I8jeulxICawxEDQylqe4B6tVuAvUMckw/utCv5pNRh1SljlzS
ylCUGS69FoW+BRgCHEsWgweFGIdJq2zuvWJtQCJPpGL3ggvx4enpL4H86du6onsK
iQRRB4pnVVCk1nS9kXpaBhSHBlrMc4/fP21gHyzOkJTtLMJIqHAn3iwBdLxp4FJO
yYJJ0bJMeL7u8Qg1L/HudGVugVRTvFPwMObEHQxlpJQLjXnP5iVZQiIf3fl+HEDC
BRE1GvAJHGH9P7xp4QEGCVaQjxZO9Irkz0iPmboCV5g2ASzN49D3YBbsweguqyeC
ugfS9hGDhrbLWqcHTZSV8t2zrBu+mQBZNv76z+YOAO2r/gVgN0lluiyUTfNcq0xo
9d8vOljoetfGqPoWXC26KpzAdv48TAQTifYeSLnC/iPsl/Cg2MoxFyusEeJX/RfC
ZFR4WD/d2ptzQecq3LnlZXj9iaw7DKBNIyYLiXkOtZpD7NCDOZREhatYvzWEzR8H
HiZZo3VxnEkjH+Ze+p8IcFEN+jJjJbjmIDiC77kRNw1TdnznyUpll5nd9H/Z+vQg
sfAr+275FWk/WAcUD08iT97mpgoCi96Q9jmrScs7GqbIyOVMtbLoY2/PwvK5YQpJ
y8OZiz5SnJ0dTkKTLnddlHFBCmhE95TwYz7GqP4sJuIpI14paTUM6QyjBZYInbHe
iDTd597rehqH+Gk6BvZJ9jHq0jsvp7wWjF6VGEW8LQRd8DQjLSQcr86d96j1LAxn
HqKV2o7rfPXNFM0OhkrhvfjOF7OFkZJyT7SRCq9f97BvtjJ9ExRAEVTbvAF5Y1ES
qCrBGSBWoBV7eNpoH+8Ut1KECvoYLaXMa4fypAqDnnT9QeTupWMvQn0TQLwMCHjk
A/4WJE8blyR3eeD8mlG7UGkkdld2ggggKQHrF4Pm+W3dvOgCDp9/AiG5uzRqojKG
kE/CxhaYNQ6kKQaAV1gbyQ587WKVRETPmViW1VeDuilfrgaSUb2txvMhq8eq7YBj
qqu1HjcUkClmI+rjEP0wtDGqod3EYFix1/PYytYz0Xupq8XuZf/zs/4vjAlNrzDN
FsFBDWz2x2oFOGQ1O4yETy06tN1MNvWYBKnm6wep7AK9xOB0PWANM+qz0OA7D48+
DkiDCg7EwFmqbqQPao41oCvJszW0afkjloZ4bwu+u8R07SP+iifYbGHLdLESeU6Q
uas1nBS3tNY/RCtERCEBKoOX8q0+VOUdHnLVqVwYLVXya+GW+SS8EK/7XBVJAH1u
k9N5Gf6OfhyUkm7rn1p9rSlP/KmFqAaS0w8hJBtVwV8igbzb9QqmjxLDdT0Wghsd
6J0S8Z52KcbyxSSR9zaBlYlfvNuuDRhYHmoHUfF78/x+o/QjGOgO45rAmeYJ1wGW
dxiEElmPV5YBsWulnXaCy3chyVGmXipymbwXYSvAacFnVOax7fp0KNw29rh2/MEB
LHttI5gUJMQ13W7PV30SnoovmmOK3A2pPVn9uxdmF72uruYM9ms6utNmxIiN9oqE
zyAoGz5oAncj9vSQou6tFCBauaiC9Yf0kXSZBiVWALSpw1ZU0ZsLWSD1s7gsHnS+
ch335+U7NTE+xkxbyAuLEQCIdwY6QDyAcJskFn+LS8oxxzsjYfILGAMpVUGqtXco
Qe1/RzkSpUAIox+2oT16jXiXFoRTYWxLHvolnO4U8mu42KF7wrOVX+6aTbTvXasq
i6wxDoxbzK2aLvf3FI+Bf1X8YJPpfMr8uVLn+wUEb/19WT3CCzhIt8pIlalIQwhX
fVYXIKV3uBa2s2YROzPlPTzULSiz1F+TwcdNpCg9tSFHb1RrTZRkotWY9QKCUt1w
scJEiiTnU2Xb+36kpBk18QZkf3KJer+IOYr4m/VWoFBtCrMLlbz6QhWDrwWg/IAr
y9NwFAlt4AZ3syTTz0KsQyHeNinjXDOoSO/oUoCdeJQCO8Fpbq3ML0wapyr/PQuQ
YwI3Cniq9I7HCHD2hwDdCwdrJwT0QWmCxmjrmF+TYPDm1Swl9xW0i6O5SWSHFH5H
4iJjGfwRvwWnWOyDbGR3uIQF36tFUozfDFAu9V/13Y1jOAbLlmQdJSL+V14kbEf9
VH7riXg1XhUa8uiRxU305qHnDP9ewt2Xza8OVTS8zq4jeMwtaNTpIW3yvOkc5Uay
SzagNC9mFF/cJcM0Zr7E0DS59wBQpTiiE37HfknhsgOvR+3CV5dNgjhETFhyVXBt
5leWtw7xFw9+VerrVWchZsPMzmkpet3A3VDQwFoyISuUvQfzhSnJ78E5R3/wlZWY
rHAxQLkgPqGJwmDLAt5NdIQKoaVLKY6EGYXe5Ahlqg4LCJI8osQvGs2VoGG+kqdO
ikpHmlfmwvoid9jTPUJy4olfZkIibDTIJLa+AWSEz//bzlpjmRlEkkP9rNuN9DAv
SU/TXJQEWmBIO0zTA8PS5NLXLAZeHSK0I7s4nOvZZjZSdSvZBprC63vGOeMUSDh0
+7NOBkqn8RpxrV1PFz8PqpMWDubBes5w6JPQgp5wTeQnapUOn+uotTRcVrQtQY+e
f7cz2NW5l6nSlzZuC3DMmqIXrF3T8SWV6gxIaWlvhIgJdAOPK36Hu12miKjBDF23
izAhkJguerWuFzzVIfYn4YpLFPAbA4wBKf0Iy3iTIrcMMXPS71p0K+U7p6t+QI0f
d4WJ83NPgBZRUB2/J2JHTAEsGQROrFcM42XsCFg76cZlmHX0i89sQFsyORpN/GnD
1NJxPm2XzSs/mOz2P6rov7eCoSI0eX3B5GUsVpoGENkZN0aImrI6ug3eXPsxZXtA
Rlcleg6BcOEKiekk4A02hAYgAMpaO8tGqo6A7X+5jG8D1lni7uyLHr9ZQvjVgaSy
+b+ZCSF7GF+6kBmi4bqjKckR0hsvNBpStP3e066hZodBb73mh8g2ffQ55ph1mqJf
NXpJdmxGWV1Z/bxpu8AVGGNU/aTxNN3pvL5tGB0kRUIDDHL7MjyuP3WQetCJYSHG
8E1TwVnTprnC0h3sQnrvmxCHymMZmT/BKmUf+GlWZ1Mhec01Nh7mfAOn9CaZu9KU
rg6hLNDTTariqzBRVC/DFsE56+vtMzkIDYzldDNkOYz9IT9z/t9XhQW63dtyEWWK
W/OUlXvsQ4WVzp8KWD+X31qYNpgZkCfLNhToYrDo04mQUFM/4Vpy9ByP8XDUonTe
boJMLdILi7aQ2n7CnBlw4U7THCSPukLmF8FJuO1YStWjt/41bv+UvxShekeXcBLg
KwGEliTGUCrFE9TlUyfJSLwck7dImerOfMsNXFxNtny0ycx0il4x4R4UAj5wvS5y
3z8SrNm8wI3lThLDz31J+E7P271x83a2PoAksRGg4TQrmwA+rNVdvAh9D3VwLA1R
UfdBjBi2KB0lRe0XkY8W2lOJXK+2aQNn4x2UOUMSIC5jMDuYj9BQl16byKmRiS/m
1J6DIDgZ9TUji4vwWgKKqnjJbcrpE6XzafxngFWPTJ0tzqiJkiNH8UpVEZ/77lnP
Fe9H3ApY2DqDZSDBYumLxCXnhehqFPZ43zax6oEYCqJGSiMUWb7s59/bJOg0ZAXZ
TzyKjIfVpH6OYoaK1KuQESFyyWKt4zFNBXzAjJoKBij2gtHfRrXiKzYgFhA7nE3x
AnCMmNaTlL6weBRjUKoWMOc8LAyHM0w5LQgZm8h91ZaNmHYpXdntwrFW94s4MR0o
LLUNJiJBr0O1lwU/tdlUtCA2dyaaXChkVGyBh65eUwe/sZ7ZmycP4DZT4a/8sW1S
T5hRPa6c76xlD6h/6Zhj7fhaLXvyaQFCHL2dV/1t/W3amhV/xtirtrJlaW6Ri3ig
zbqJF18mWFqR5073vwbBwwLdcS3ailvWMQllDCi/LrE8zDW0llsbWnPw5jf7V6GR
c4RPCnfSPQeDGyePSWWmUASEkXjNQF5YxPn1v7yONq0XCuEpaGiroMLBXCWWDjGm
A1o825XY6y5IdeLmM/hNeW6HyxQtF28PDYGwL0uNmRJtHnKr9KgRggYIZVIm1fAJ
MOalelIYhAhuOk+xAUA0PEExZZbN7POOEYze02iUE+oWPd1KHHYGRpMUV4nwGnwk
PiyTrmhC+244H4VSjoyrosU+qsnDA+XeRUFp+ofvJ7ZWAPMkOFdQqR2vni2yi1h7
ajeJstIK92A5xorZZbNb1CXGyDGOl/Ro1eYyLRhtscuZfniaJA2Ra51uZT0b59wK
kKD6QuEeXu5/Wb+aIIjyAUbxB05ylP2WUeQApWBz1jA70YPM/Op2AwYp0g/n8gU7
v1HmRHPkrJSVznv/s28AGzkT1+2dSfW4eY3yrx6X2foCQ741C5xRDNnQccxVmd8j
42rFVuNbMIsd/r641QLCeRw0KcQ/NG3MaYvRpD43H/sQ/SQKfSx+LMDk8rTcXFSt
sHnFSBKx/px3rse9RQrEpkeZ5qqNcTO0uJsMi0gB9y6XJPl6QJWVcd6Z1qvQMVIX
jD+jEiYLP+rUojIPLKf10Rb2gkGR45SeB+90hz2ztx+GyFuSTCz5fkJWGiLRCXDK
2edmM021gStM7azPOjrsZyFwP0TznPw7U0dScmN3lTlO9Ux+65pbw/0dH4tOYBKv
3qMixtTzCTE6UuziN949aXSD3085PFiCKAiL/H2eWspNKwJPOqMDD2NndIorijUF
NnujhnGFcQNjnsiXA0ylMO7cWA2iwjdvuDu5yusyh4Hb/fs0/WoBzQ9oAEwyZJsx
XneHd7JH2tfgn+qIa8/nOd8/YXdS0p+NoBz9aTlbKNUSTw2z7Q7XvON3U/eHDlI4
vNHw4JN5YEgjkS74TALuzVtyqnLBm7E9oswEqHcZDOYPF+0f5UfBxOS/Nz95te33
bzCtRSsUh4iRu+wMnCYen64n1+lPMjubjG23gdloYMs/YcpKhXo92E4OVDVS7SSp
Laj4yFDTA7DRdQMte6EAXWY5nTS2iqlvDo9Sjis3BFMa6k+kikAAfXpklkwpJGP2
HLbJ+YyNWyf1rfWDfNAeeXeQpvnI0rFJdlI5zNdbU+Xy0DAR8ohvrQas1/wFHnLL
B6L2CTZnH8lYH4M/o+j0H7DU7L93jAVQGzuurDwS+KGEzEL7/4RQQ4113N8jOpPi
cIu3Cq+jGYCjPLB5+zg1GEJbk8gqdMgMNarCS+9VIdLh02fNAx8Bm1+PyBOzuonJ
QKNPQQXNubM/Do1I7/Lu5EDqWCv12zGZgzG9bjlkVwQVmeAlgwtxkSAcP6iYMir4
t+LWqODkzZHvUpOid2AuWh4y2jF9Bpap8YTfZ3aveo4rEmhkxJTG3vag/aDyE7XH
0b34OJGjw67jnLssujKh8ycimTtVoHxIixtf9N9F9NTNBvEpoaFLh53z+pjDA+Gx
fFgDpN1UpiI88BU7wShUclVx9KIx3VTKP907rVwOSnpblkoo2O5BO0EdafLxoJBZ
rFMjY+sKn5mrFeKwSzKjdOeH4zfCzXDsh0CGuHvo6YAIazAGu1YhsI/bzF5bWR4Q
Hmb0k1yc0eveNl+LLrEACcSKXFrsDsR1AymOLKfLpaZ5waz6F4yPp5V7bI7WGU64
kslOQ14rd1DN1vOA67vZhdS9rjh2I0YeJq/oXLIZVbfybX18pzDoMBU4oTieByxH
wO+NOJvvSNN/Xao4yO2+qrDZzDi2q21Stp6yl4I8WVtpxb0tOlQZt8bPlPGWXchs
NJ+sBNpiXLdp+iQvf+I8G+3tOA1ZcOmGLwG56nKhZKaonU85CAPByQksZA5QEtHN
R/qDPWkWuDNpJiS9P5mHdhrVtBx566CYZCXnAc0zvoazENGL1Q7pQlLUxMtHEAJl
OAPrTQLl/vlZoi+1bDwerXaJ4Z4fZl/i9ak6ogEELjln75k0aCLsfIcQTjhx3wkc
yrJVT33iISc80FRPDwguDMlb7d0p2TJ0K96DE2wnzrElI9A96sBs5IL5LFmN/qUn
RjPcjlxWZ+w10av24RnPMa2XNEeoReEqeWdtbeG2qhN7wviOFspnsPnCoNDRHrev
NH+AnlF70Ibiy3VnlrDbTN0orkKNB2331xqeqzUGy5hTbOgy15mICEpzi2JHduzI
YSaN2si0Oa9wCaKCpE7cOGp9jq5BxNgpe0CTlNd03+l1gCdU24yKg+Hcydp+JCaz
N7cDpZhfQH3+AsOBp7vdBGgOI9+PRhjZ4P/qcexWvNly7D9Xvv3nougV640dOuDO
BwvFqCGkt+Xq5tbFdpAg+vcRiPloq+6eHuiMRiRvyFyDohnUDnhI2PqDkTrtAplS
fW4vccK8i6WOJJnSj1jaJ8uNOJEuL4SW0BVa1qehnUUU31nKtoyfpogAf1weX5pM
jrFVEp6vaI9yd7TUZA55LyOKM84UiLz0LfjQ+yOCpkPSEC4ShuRX6EhJfc7R4gzf
LEls7PBfiFSZTl4w0EjeymMTiOO+wG0hn8sBG3OpT7GRquf7vREre0dmlLDSd5BE
rDN1AO2IYBpjD+Nq0M3Mulkpc8eRlxOjDAIs5a0eNy8J8vVmYb8vCNnVRM3sADo7
49XUu1MFJhvv9uJLa4tlRojsNWYBzDxoUK4T43M2vDjVWTTaCaxtZp438hedhHDu
jQ1VisQ1lXvu2Xb3cIS4WE81p469OQCkY5eD31KAjld1MjDtCQSX4re+BrkjAWWg
c6Psg4lpCrcA4ienr43RazHR83Gefbs001khoqOnzRwaW8JKDhOU9kannUdUqzOo
v8KU3p/MdbW6WmhDVYcezXhgW0t4A7iIXMqzSGd4zeAu2izxTAdeVlEH51bjimM9
PeWMqYqbGRRVpkrAGg+zBkKhGZHwa4mtxZ56zsPdKRw9QDGUa6OBTY7cmRBEjPsj
mWc8leoMGvGVsfc2Svk/FwllEmaupqEPtgG2hacQFJPMQDweBmQLWvuV9EWeM6Wx
iT4jMUH3rAPzo489Zo/6xLbtzwIEeozTsCsjbgUCwki/47FxUxfICabVMm4ezmLh
eBGF0Gd56tM6ID1r8Cg0Aa6OCK/kEUQfPRwkYqtQP+gxxFYNg+USIXl9kaESAtrw
KXbtcE5chhJ8VqWK6QbWsX8asosV07zxcdeFsyni2O+kQXajrx8KqdraI3oAiBah
+k5VlRfRs8H55BCyYCVqefJMiv892vKtLDtSDAIwUP3OdGlJW4bwULvSrDxwzHbx
8eBjZzPavzvNh2Fdh9w2z8Vq2e4ZB7vce4oU5YtBs34sxHHIvSaLCHWmpMNDKoSC
bSTDouOr7qbSVdVQsA7Ma6k7ifM1OegvMNAEqDK2CxEc0bl0agfpDMeTR0WgaguW
v6jU4SSOae23h90kcV0o2Jk2Us5JAtajHmtIrC6PvR4iIVan3ksXxYgRuV+S/7i7
BwwWhq6sWmZUglIY65CTKHGQ4G5R0N6FNL0DeP+smUzGsJS/8i5RYzL5WPJNcrZY
SPJQpCAWUF1IYpRUtykDLXjnC8sVwhvDiSYbft/r3SxbUCtn8i9QH2OlgCf/Lw9H
2QZk8E8yYhX2e1leLkXFuXxpYaHop8AOkue7KWLE6avuAdb/EQl4AhYryQc2+oGW
q9lkyW7w6JQLCzrVWSRLRu1ntZ3OqMTO7gyBOv7/+UaYn2keaTQn9AhW6eyd1GSM
qTKcwfJSGykJKtjJGmOrDKgeGcUnuzW34LPpjNax44Q9vU5ZnKPUtzsJbpBNFAE+
xUmw8g6S24sb6EXHCZO45ZgoJer/AJ+LXxLwAnMEO3IrV+kkir5GFjmYZ2D+b3Ho
H0VQNe6ldhhEOYQTqMIb7K8In0Zk1IOU9EmCfhKfYFis+symAiPUTZRv3M0ph7LP
WgG62TkMVQQ+vi2R2yPEfTi2jtABqb0Z97HLUfpB1k6Vl+Z54pEh2cYj/ZC0fWMO
Ov5Z/t9Meww6aHu4KFVXvdC3kIJ/pNYvDOkkpxYaOoMRl1JeF7Z9W/dupN63c2MZ
iMlNRXhOlGGF/h3J728ZYatYSYGebz0pd03DFnFVF9LWY43vtqneAYSsCgVON7pz
zzfzaLE/6wTT49L+FsdrUrkYtc1ES4meBkjIDsAvF4HykYwkLw5cFAJRD/yAYJTv
P8kUK8dT1W279r2kb5xM0EyLPvbwmYXhhKgMTqgHleFcrbEtZGIdMhW28yveuJze

//pragma protect end_data_block
//pragma protect digest_block
JBT4sCnDJOaVDy0unC4mf7bLU1c=
//pragma protect end_digest_block
//pragma protect end_protected
