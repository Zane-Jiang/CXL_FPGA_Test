// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n4o/Jz5kC69wvkXx91VDBLd/T3czmjiJidVyg4w8kX6o1Znz4Kur68MvwddB
JUnxA7G7fE4sqCs20qkbadVOiY9UqNto/1TV11gdYQMyEQ65Yfy0PBrudEWd
npp2y8J00tz62vrfYNKN7ce1dQ1je/BZ/vjUAJk7/NCI46ZOfqlCjC7GeY1T
rrRUFe/sEdeO7/YX7BXCtkmRU32N8ijRGAGUQU5KAYeJpPZlgqdUI9E15N8I
+ohf5fCvA7Q2PzSrCczRmD65mLmieXoh3AdhrOPjl7e2XALBFkK2mPamY6LR
75/C2379SMXOJx1bS0Iz3sPjdI2YHer0vFKcEw15xA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eehYu3pDiyrv4sxf/O5pWj3Jt7fWCn+uPl45+r8cIekD4Ie9JoQnzcDym+Cc
ONPcWw1G7vyNMP4ed9UKa5vdCeiqNIi960vjNbms3FPzEzZIoNwmVraWgzh4
OwTQmfdFJt6ov1dIJXzIJIzC0OOUpZSL8hlBADxPFPBLpiLFU1ekHKWdHvcx
6iMuWCWjSgpcUpzE3UnWIwvPRbw01gCJpO/X1vGBRDu0V55R2I3qikoGsm7O
ZMdRMR5lr4q/8GHvIl05krcJ5Zz0kFcN+psfVORnDDd3MzA7EvKOk1jZYtq6
dY9u28yvIs+xuSVV0EpqoiM1Jr0AB8DIzi3bB/hshg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lbIAQK8vKBjefXY/WfEa58cScYqPtuYzzPZqEvmd2ydn4FWBFmXkYdoRxZsW
hU42F+1eatiPgpXI00wajY30JSv1CzsmAia0409Z/j1TrxQ48XT1QvFmpmk+
T1DgSPrU7CxC/ooBw+z6jtaX0xhRCN8kehLmTHOOOG5vTqs2BRbc4hXy9iSu
N/A6Zfh6dS/gQqbLncksChlBjNu/LrWbQMmyK1UuHNSZrv5c8jWXZsjRpAUr
dE/nVYR9e3dtxpeCB6GCHrfYp9kJHx2tC4SrZffH17ayka0R6OudSPkpV4Cu
8LhWCPSba37fGD5umaYEvY94h45D68bRR+aDzVsfrw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sMGpzrHyt75Fa29CNx/iS21SUmTnuivRp97WylZLY4o2kHaIXLG73lmavwWj
662fkOSmY/HU0QF6qik//UYhEhg8FDV8RylqLEO61UYi2+UzURVUSfztU7DN
nk88BWZLgFbFr9/Zs2YFrfmBvYXSOEtSGEVALpov8h3+2iMWhg8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZdHhpCHSvZ9r/jSCITRyEx4KyX7Wt1M8bjTyYCfSM1NCyaoS2+xM0Pt9lnQz
rdU0M8fy4EGTx8Wtwn7Yzey6S7zV8/bLwoWrqqE0IMLWhNfWkQXp5AvnieO2
G6D0RFbmuZfG3aYVOrO2RjKHHaXRNJK3AZPn4weH00T+sFQllc3x8PNr+C9B
rhLOgiKjQ1GTm6ASl0ckuGPutjpm4InPSKxvZOLS/GSvJWbrvlJxJqsodVx/
MQ6Udg5zrSe2ZVv6TJIcFFNU4H3TceIG6PRoJFJkvX0cRWU7/GTulnY4Z4vZ
e6skRdfiwBGukORo8u7GXryvDDPdalKhToCpV8dc0K70E6OhqBird73L+WAH
Pojuo9yaXU7nTVWMHwcA2hWXOUQFDYib8Te0pnNuYYUSyNt6nq4QYkfnpi2W
oSoes8EAvJFImTLUGufER0A0rOGPVt/Ga0VNQqOmsUQK8X86ojhl3V8TFI/k
ntc1987q+FRilW8aGBS9zlvzPDu+GDkE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dRdv2NjAqolXxdKPOPOVLciL8jbx5c0Yp5hvAHfU2RXOKgVXF0sp/146GyYZ
d4Emv0gEMCZsZd1CJJKc0u8sj8uWOY+ymBcZuh7LC/d5++ECsAH7PpUvzZ7w
T3v8x4KuQsJL+fQR4vutHSQDQxahFiTTBnHNXh5PzwZUQqRxSro=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rapVlnbS9rN11rysHp5rmAL4O3v24CORRJR9qv4HDDhUZXWDVP1E8/pO/IV2
DLGBpJudmn0rR9tmdqfRyCWSbM40lMTeS6LGBixyGYRwTa/ELnxbrTh3wIO8
3uEynqdICBIgKkv5+lp0APe1SbMgEgDtSfX4TtOis+4CVJ25xCc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 72288)
`pragma protect data_block
PExGlXz7zuJSA2B6tGvt0JJh3mKGOGWHcNa0Cc1Vsvzmqb2WwdrAf3BgFBMI
ISigPK0rs9uzxuJ9c2w17P2e08t3/zsnxDZ3hpZQqPFkWI+MpJH25u37rUfI
LnZ+fcrf5IBQZZVaM43NWd7WrnSdH46kmtH0bn3QI5KvbKLGGHAE/fuB9Ghh
XmEgGRq3sPtecNdM/ROAQDsRdlIwjDK7JiIHOUKY7+Jj47gc7sS3SUF1RKSf
JKKLslW0caOZJm/9PpuZmI73EmyzKBdmSc+fndaVZxzcVt8i91KnuQMQxdpu
WAXZuGa0i3DeeU4OmXqZB0nvlNtW/vVT5N/GuPiuA/x6Qlzu5wVi7zYpoGNG
sUy6Q8OzSx+vjf3kRx0ik3h5w+2Qk9DW0e2OzJ+juXVuG3U1+pfbHJxq2e+2
cSKOk3dmF/CO9yYOUpR2/lgq3Aa0Uai9gFZhFndU4o9GNc/2DW2fQgzNjyTo
TAjTRrzng6gWovmPum/QBHXR0tF8VIQBsdgDcjraGds4EePLUCJbb6ZNKdkO
Wn3bHIFBGIwL6DHH6e8EEEtofaGV3kHL02Guiz7B6WXUhaOulR4WNShst4Gr
76nfC9XbT3cjzBeO/S3pB3RdKZZ4ZK6lo48pRoj4qFuxePdHPGL05kfI99FC
+i0O3DraFMzEYHFJp9ytBOZjuet56xDXC6v9D0ibdgF/absb3qOD2ds+gagf
iHW/RYX5ItveJsqGdUjHV5h6wtNGja8bTtozBt49pNiJwhIwWj75FdRFg0qb
hksJlvFdRXtKEYV7EH4giLRXuFLqrVFeQAmZn9CZOB2ME17LWeSNIsGcmf5w
7RwF+xA+7lB15EkrspxRLP3CNcZPzpIbb8qVCJpOm9d4G8yllPZcX/RLf+kv
FoQL9LZJW8Gxm6A3C4jweQauYAdfaZnuBrk4jAdgria8R2tR6Xlg+L3RR8lm
6Vm3UxBx5BnZaXepmcGXDDNRaWKX2OheGlJpTpKJ61aqsN/0YrJGW7hr2Dmd
GoniBBV6lJdGcah4YKj2Dd7weVA6h+FnFeAxymDTzeNJyfYYE3ZOJzKQwLlD
EDl3fU/NW5+BuYdU7LF9EfxIK9JJyJP/UFn0B2gyTUzpkkfrEQUWqlL+Bc/A
KdjE4oFzHJZzzeCiybwAfNbVG5hinoXm2VHsOEFOv0/BJGilKpXrYJoBLA+2
1z/P7AFSXQFJJiYIrvHhsvaMGIB4mq+iaLU1boDhyoUG8/zWK9s2tUQmvy5j
Ka5ykn9pZYL7lS6uSUjBUdLE0okh5djUcOb+LY/yTCSFZMd++Jv5AgKWfVGU
zC7aQyjNK6HNn3pWpgxh1ywcRqGPn/pJ7B86I6JbAQ8Mi+S6vbF9nHiG+tcy
wCOvERG1HesuXDckKV913bg7tJ/ampq4L6CO1QZBwvsj6vtuvllwZUri//pF
jaIsrHDdWOgQGgm8jOhipK4Jdzhkfz7NJf7qif5L/pqE7JMyMpeU4bCmcnPQ
Pe2jQvb4Qc+7eBx8PKhPTd2pgQXNjSuWRLh4q6CvP6qOzP1LXuUge/Ch44iG
zF49Y4gJTu3aZMNQQ+j+XFMYkXg2IBPl/flzXslqdn7/ba3je66eQ+k/oYX8
e/7LYW2d0k5pyW01AE9DimiqNZZT7R4619nLHe6wPxDqfcFk+Bz0iQ/tcSd5
O8Ap/oEpnT8TD6z2SErH6/G6YirWfr0x4AWRH9/Tg2ug93uqTKgJ7Srob0MF
UcJHpDJGwDg6jKJFN2bi7x8nKuOWE9L0JitWKtyvveBqevjTJQxNw9F3Qi39
4Pw6rDunf0FDKJ+fgQgjahVL2VIeHe7c81GVUgIGy0QUVk+y9aSTOuNvY6R7
TPRN8J0L1RsEAEjAYnlDowS3cHRV1irUDUxnUgIB3JNLTywXh9MUE+cDdLmW
5yO+0PxwWnBEZuObm95l0VW78ow2GCQKuuIORpRgARwqO/0aGxxILcuoo9Qu
HrAcEZnaEEEUQdOMC1t6u5dcunfKisGt6Wjv8bhdVX//zw2zax61Tlh4gi+r
lGo6tKhItEEgmLW2CrTrHKyC/dtJNL/OTOhmXCAhH9nnMutU0SBrC70sNAms
ysFEGvDaLQX8TEcqow6SPrBeTcCkEu5sJ98PeqDotZFMivz/bpsxKib422Lu
lEI/QdFiYtYqmIHNwfE5ZnwAG2XqvIb82lpuHsfGHSN3nFhkGNFeJV7upFrm
QTSklrasK0VPZdDtnCFA7szF/Kcw4JamQZRxdO5AlrrFU6sx2yO1IlCJ5/fR
5Hoqd9YUOKHl9LK99EwT9061TZIh0t6OZ1K/MsEzhgbLn3FxjcZJFQ/ZXGnb
GyftBH5aqPN5Etyz9GfbwZFfbmZjmUa1ZYBpnJvHL+H80i+eLcSbhofDX/ev
YfOGyl1+dcTDS3EC/0/WuS6VCGzTa+buXoGJjh44yn/qzDeFw22HhudefjzQ
8obiWp1UXQVi9cQSKe7BI0WeNaDy4Ak1f4zq7+IAPj70vFmBaNoGTCkQLEiX
8ft2SlNMK8aPyW2HPMfvPjhOj/57alCStrSny0ZVkU6Lo0kVWnDDdKnWzblV
X3zQi0Ea8MpZMGBrqv33WGv0+bEWXAPxLudx+CZGVcoIJ4z/TaSzTKrtF3mH
x4znkqGrGSq627/STOAvR5BLDcdP+GJgqvdSmLMQ4rGmjXTtvQukAT9j1C7K
a4kWMrc6OhMXg3EnmJ1MbmcgnNb5btCcWlDZtf1lbY6NLjCyg7ynm8N/C3KH
hJsa41lvKdfp5nFv7Jbt53LUq3AFAFNQ4A6LjEBJzvyx3D2Al6Ue+5RCRymq
5IUkEFwdOvxDnpfiYQ98IRHkhF8vz4rHd46fUsbJJZzhr3t2ioXZdydvFgcd
GKkPH7lOAoKbqjcbDN2sNBS1HVsSBYVFf4CYvb8dGin+cZfVjMu3eet9jedb
7lF4N+fLdjDsUZGB8z+ttYJKqQPqvfARJrq5PmSP2H28XoW/JL1X/kZfjwFx
PAACZHDe+SddkJhL8LpHhe+0/+x13GfPyAteC3VoTk2aTz9Lb7YPMxVVekTd
QZXMlb7BCJtERwB+HTQH7TXe/uPLXrnYU6rfU9OxOtwRPeCvA7BHk5FNPHeY
jRCyH95s48mo9JZx551hgCJKoE9Iag3sPUu9GM8DcPNWQYjfd20o8CE4Pjf3
1/VWXBm3LVl/eLe2h34tP9eutK0iieYbpC1gHYJNaL2POygaqUdqVyDaw63k
QJHXRxlpcU88ho68G+SWQAtZIjr4sc7W8gLAYN44Pbcwh8LwTAaRmkB5ajC4
Bn/ttnT5Gd16lclQF00zaMqj22TLK7ZMNZa3JTRxhQByV/bcqiJwOk6m8855
UfTk8PMuTftVuTN8PrKI5uK6yW4T4/KcqKxSrL0Y8beLugfirUw512BRvg5k
z8fjct/TPRI9DkuLImczgN0HKItGmR5QqTFypTGE5VlhkBwTGtS5LYFT8fH5
mfnUKRVPNR+kd16LRqiu2tb+ht/bTO198hl2DNg83tIGZ8nIww30by74tKJD
CQw0ctXzg40e/cI+BhNYmWii6PHvcgPcqk1CA86xewCaXuUD4WdcBFlUa2XP
75VC6BO89vF0Qh5wh7ZH7g40x+ePujVZJycHPRzBuYXeAbP2y5ybwIPAUM6b
8YQavrysYAgidVIwmPdFR8CdMRDjPYE80/ujAFMFzvTrOuVTbqoSpbV0Nvz6
SE2OcSDh8Iw1JQHzNOtBusGJ7x6ejZ1DZzs4D+WXrKxgRBHQGCDTUFeUDzxm
lVhDkcSlfY5VqA+IF/y3YiMgZF6fINITpYN7S8Flh1JNiN6+rvFBPVZJQrYG
44AQqBo2raby6BSbAnwgbH1T3bHZfzEGRBZymJQyKHvUmyrnqdoJXXz8C7i4
R9o/wWuDWKjQISbRRtK+8YA2pfteKchgXQAL6GYIJMkyLP3GlUEgJ28OEC2h
QxhGEmglNGxLP41HP+1sCrfkdgC9YkBA8ivzxToAgf+pwmArhzBb9ay83o7X
6hAiF26rh2ZEPXqSbEYdA640CpsX+2aWfO+hPRqBiQ2GP+Ib4+7BpxDB+VyI
CTKqF6x0354rppJ5JIdOTiXzqdohC3H6ifQPdlUyZGQ5BdELf/OCu+pe+3jN
qQnvqvfj7HW+bAYnVn9eXqf53H6EYn+5WAbSnP7TnYsumK0rv4DmPRoOxXc9
0isOU9ruPaRwyI6w4+His5X0O5flj1UlPVtStZlT+u2zyFis3Dznpjv6Eioo
JxMzuCTS5Ok4EdL2zXdDXro5dTM8Yk/X36VxXa8Py4wOHHuNSVAkQfiH+Tae
wdXmZcf/L7bCnzBSTpEmO6XaIyCQkexYumQ/AmIj3b+2G/j0dPtimyRvhMCP
pY+6RwlihOH2eSYbObp9wq1KcxPrATKXb5PUy8k8nCQA6kxoXeBgiOl1hXbE
Q+tEpfVKy7kzPLbFlBgxBea8S82cb0oLScI9/iqE0OKiy5/hnMWyRG1Y1qVa
TqY3AzeI53u5A7ooiY2nS3sFA0pM37ODbb30ZYqvJR80Qw4/xJAQvotGNSq1
d/nu88qRH8K3ie9ZiNbYI/sApIPvjjt7Izem8r+Aa5BadvWw3osoDqOBQ6oJ
XUBtEmSRFOzvxIXv88AWV+gbXzZ29Us0fJroHJ1lG0jX3cJGxIHlVSBv9b68
AgS5B9ibMUmHN1Onh2BQgw9nNqOvf1SkwMiP1XYLl8trqTyt5oXQgVJVmM3b
6JBoDGqhkID5WxFZSJUx+vJ7sJ829ehpbsVxv+FxYTJYgktfWofCnFoKHXvf
RN3ZquQlItXIRzaN5Nzm6tUOmW6ygMCEWoyPTblEuY1XSTBDiPVwUCRUDxed
2sdv00cZ3O5vhLpOyfZyvfI7GgbLHstwwacTKlQVgH8F2U3lJOFMpWB9zVYK
fL/3iEiu+UKc35i4H6x6osrKDrHX19Fg94/TvrehuYyp4SDJ7KpCcb5bJ/2t
wnDQfFJzrggOk/lCN9OUaNb2WLEWpnlBVC0qiqMiRH018ULrehMb7vMTtZZK
tlL8wo340kw0obFO+jxdEux6+IkM0nTQOQ0OgeLfecr7K3otal7Bbpi+KuXt
B10ceP2wYNYQAlGgdky15T8X+eN5gfzfYXp4MY4Hk0yueFMU7aZj43UYKbnL
oljmg7IYzFmrPYerEdMk+Z5sZrxRUKqcJsa4HZuNUmGg8gov+QX1yvduMdQu
bXC+PfC/4SiMJxw8wncieTPerGPSvtsJXCudEzDWURIU0KoG51gu2X9zRRDa
hjA8s42HmylruF5036AheMbVwqYG6zTROCFcweyDOeSYkapfqdfHR7jSrd6Y
0W7vCixxWm/6dTvz83M4KDRWh72fWT9HAWWCtzYH52sUQYASFLUrSXj6XxdH
OPFkoIruCK7u+HABdMvNqx3jHWDuCE94kn5x11N50f+Y13Y9amPsNmwAOfwu
aWSF7qVkPCcbghGx4ytiFJqQTToXNW90/y/gB0Th4espcKtH70xJ2B/PeFK5
Qn6pqAIfqkbt3Uvr81+n/guWmMt5Ol9PAVxztmUfLiQ40897OhXbpeVZF5uu
9cHcxjqACY4G9dLTMnFuisg6GEy8F+9Al8+GK+LHbf6Wlo2mQHLOKZNecrEF
ktSyq10/l/vmSHyRjzTy4DkP9eLjYrX15wxsiJ7U88LJi4n7tGjzcBdQj5rV
yxd7qmvE9v3MrQcFQI3BXG+zsEWQsmRc4zzrWsSKwWY9lVvtEVZUAc5TMRYE
3Srb9R3+LQeEdD7mOxhbUQ65vDbFkmM6PTKZ7kQt/o63qMMMKFttO9KV9l3V
AVpKdGUOuSno5JgS9de2vcagt2/g/4TmkZYVm7VrF5i4kKMitFsKEBEZjmnW
VjDeqyD4lFIgtZQx2wpygcz1DlwWYTRHx/rIcQIVLslE8RvbObGOoY61NakS
vmpewX8FjxWzSHsZiM5he6I5r5WJp/SZoORFHrnlTGw3DiL8/KRaLkiUEJNJ
LneRdMRDa4pbekyi5IolyUEeV0Jzs/LWLRvlipoNC0d8eTdTH+z7Qy9DUYMM
EXGDlT+f0+C+cVHUdWCAxwb2xnabNWho5+jYfkAw8h8RVYy/e2pq0QTgz6+M
nIu+OUQ8Ud4gheXR7VefAN+SDzHOyaK/w7vO5AMErfqa6edUtIhqEEcINFx7
V90AvLi6lrhNf3Us+MV8gP8Sj14I2j+lIVVKgoXg6AbpCVOo7L0sFKzJNN+v
Kv7S74fVW3tTDCbXsq55a4fmKjcDT0KM1yZzgycqs+7nkmnBkPSMIIzNNbav
ppIVY2kWx9b/u5fiqsk0ge67rgRmeBd0g8P/of66Biss19ipGN52mlOkIxgu
HRX1k6akKdiv9Cn/W8i6MJUHTv3gjn22mdlpsOSoCKO17DneePw+Wi4r1YHw
hDVJUULLWhhyvwgw/VVewar9C5IMN3UEmYcl0qWpRXHNrGYPv+WPYJ2kWxCC
qYi7DTQOznZMWtk81a8GZGyie35SzaBDKXva70P4wQubmcYWoiRQ5hi3JW3P
q6zgD3TVtP9fwmMfsxQcpDq9gwb09cdbsbsePT/5v3S9yBceC41cbjOKICtY
XB5c8gXqtm2ykTxWt9EqQ/H4ZGQm+U9Q9+A/vwYsEMPcgMHd5EW8oxPCjfMk
XFpD7tMtKaJVLtgpgAxB9FNN5bsQEo4dOnD4rZoxbDujrO0bdjjUtPz0+giP
BeQBEMkQ2Uf0jvvhyuzrFSSSNFUgtzSzFUegdKVc3wndySN4YrYl4yanTwcp
QUESCwwagIP7ZTCY0aa0MAPyWWbzcyb/vOVIhNSbo0dG81qkvs9zljpo/JGJ
CkU7l6Cmcqj1hi98p90UrD8H0Yz9ntl/DmGwi81DHjUdYCADvW1vNCTYaJuS
2yPqifJqUHNJkTjFsMqDfhTCSoPJQAr76P4twSH8eKYC6zeQOVKQsNWcZAH+
BNr7NJTjaXoJzuBP7yvvtpYbrnmp0mGC3FfsYrIVjES+xUcomz7EqLnkNbX6
F0GL6lRuXm7xPuMhIvOGmrezUZ/dHROK4+uN6LWXlgXv6ZDcBeo9lLRktv4Q
2Zi0Vk6RFrPrgRcWLAp726PHEuwwrFvHrgDfl5A5ivY3iAJ97q+RRwsGfrKZ
0z+f0JiI9sjvsmbc2xlOZnBYlxfjsvQNtg3B9FvS8QxRaRxCNzupIdWU/yMC
SV9M9P6Gn4Q5x2PBU9Aw/KMhNvSGH199QeG4a+/nmYgyShNI6NxBW+tUcbWU
ZI5eJce/scz2kFZkiD4XnPpdbqlOXM8bjM5WKuDPzxD3niPNh3nHOFokS81E
yLn+ehs9h3sKmFF2kfAZIIwLcVhoXXHcrKI91RJU4xEe+sfXM8Bf9g9mf8wu
QqbYe7FCO2+C3U3Tk5BKPiGAsoG6+2ue3SN37ouMKaHVjVDPPhbWxOEtc957
CdkXK6+vT1vBSSUWs1AqRk99zF9e5hWHGBN93ZUiqYqGFelGQnfV+u2G9+p8
z++m6u5/EB6Mi75Gsgs9UmJkSs+YrQmxyTcxzH2LEAd7IUxxxgysu7QiFQwS
8imM+kaGI7I3AADPpHNGwqA2+BI95RXiIpZUrnkY3HlTo80cE70La1A05qFj
oIYAHntjPI2MVM9i/nCECECilkbx+sNq7U4CP1smZXHeAO9ftHfXrzFTIDKb
3/O97mdtJqUNBdeudVDk/W/WOgRXTOavztWx0j3OXwrM3OXh6rNAHIfUETHp
j2unE00zJMCaecccBOxRfq4TR+H8GIMfI28imuk8CPOOzZg1xmKbldn6Rkrg
9C3wFGMNHh1OoW+GVG0v9XlLvIDp9E6Y2cHKZn4Q5eYbWd/jNBElKWbav8tn
ZVeMp9nhxoWuSoUrY+nnjp9J4OFPpGzPQ6Tsg3dYJEbg4LCvIX8A50fsGVqi
cRaOn8Z+m1ZgLDz9I3zUBulUuKXwdFncndvar7QQPTqop2Kqs9P0buntXWfD
54OcKd37sDozlmYlKbVsD/S6uxHSXxq16tmF+2t5HIdfqevTFF0hEPjZH6DZ
MgNkTGAxD7VyzE2Q9O3Pgm9TgO2QikJDn10NSdzukWepxu4YJRnDLdxXax8P
hqxksEZdQWUJ2G1OgXJI6z0mmfH2wu54cHTgTws76gbRwyYKU6NYVd2f5tfE
nnq4amdst4nDEMNO3sBD2P1dMmh5Quq4rTNlnaFXgBgyksoDjO4r5N3tlY2w
K3hZ8FkBHkfKaGX36/QAiC4jp6IgeXsEsmvLPCNRz7+LXbvkDjehwrZhn7Dh
SKBlJkY8Te8W/Wndo8oaDvOMJxZ9cGhUvDZtutTRdIAUcMzBnDUoy0Scy0zS
nOvBqZw1oCT1s81JeeA02DgFdl4rYOUKZPAXur66wx7pzqteIbmn8PEQ2oez
Lo9LXgyQkhAfYag1/nYEGoR/KyGk+Gmd4/0Qtx00FzU772SlehGYYLgmtk9M
/GfreG5lZf2bnNX5dHtF2AYn3QB1e3mXHI4cBkgHNhUPivmvDc4a3E38uVQW
Guu0o1G04yK1b/ipxrulS0yob/x78QC/2/bfg+bUlF4c0LPG4x/tVszwEtCS
GeSC/O+xYnEjzIErGlxiQpKTufSGzR6j/qbACStv2Us4F5cb6wFB7dvDP6v/
Bc0g2bQUZtBZbiC/OQ9krch5Td+Ucd/eL7orPLujisLOp8bOOZrWuClbdNTM
AWwhsvZMGIU1Ypl9B2LgvmLFgHfuqCA/WV8C4am3oOAmDT5nQ5lLrVsuxoAF
8j88HWKDYFO7vFRV6/sb3oRtz1n0UHmTAqvj/GLsEN2aU7BZ0BBAdZr56h2V
k4wCZRw7E3QBMjU44ZB6Vd8X/Q98knkh5kVia3w71UHZ/8JzJuYhA1ea+fKw
hpj+J6jo5QUSbCh5wtDADMRCscEHW2nxs7kLer5pW9ekjxpENb04ftra/p+P
5GysfMnbZn7wZtcUwlRoYW4fDE8KNOD/lreYX7tAyLkdurh87HZfIou4xZ8k
eV8b7q5tQ/P5qVJ3UPr1P0D3uz2a8VdVnfGriIHU8Lo35pZG4IsGfTq59+WI
vvyT+woFVPQFTO1+7d6URD+DM+CamY47hDf8pV6E1CSpmljowK478IkWmO4S
0mCvGj1PbOYECvtPZB9jkdfNNgr42odBZOMg+2De5BSwbJeKihTl1qQm9HdR
GWulnRZnw2zWuSpasW6/nq8RzW49Pasly1JwgZI0PrkRpPTH52EMuZu8ShDo
90MKNzsgR/MxOw8fqKJJjOyaEaJVtuabA8obIcs//e7VQ9ObRuopXQQWfKYK
gxoYWePY0cfVu2SbV7wUHCTxnlo/PXtezygv+lnlfpxJSndBQVMjqa0v7bEI
hSz9Gf3q/ZE0+LCIUuejUBnS71oPWWLLe+pfqM70JLjiPifPO9Qtvj7tnIm/
PrNKAqYnP9YC8tqxOR1hv/oV7+zhe+7aBQ0msOpyCmUEZOcSfPNDGdlgG0uJ
Npy4DvirKqCQ44ruXI7ohCjf1DBS6WuHVS+73EAXpRVhtvQobdty/zGzIu4w
BOQ+fzLfpajgXQZIrcIVy+BNjTHY4Nm6Vc01trdpAhPvRr+dYszEqnboo9wt
bPHzRfYrf5zk4nmAMj9RNDoGYUgQqAMtmlou7PwNjyy/DvzV1l5Hq1UHGFPg
PLFmSBUEJY7JBzSvup2OUkqtlaNt2PamsN5GQg1IKQi1rfdTmrCCVwtMPY7h
XaEtxbNTPxZEmp+3rybTpjd+P6EVAiMNmyp2SBuZKq87URCSrJp4cqqauTZL
INDdLiCqa0Rj4C7Bp7IznAhuZB2m0EKxs/otxRMH9ZjJmYfYo7hQ5LulYz4/
SUa+pDlLsuBIhiEGmnVUM/7dfIgMAePbB9KJ6ziNOhEu7cBEF0ce8bXLf3Cd
yQNPvaB3Oe7W4Adb0yvuWsobN62NTVU69bLknhaedUWjfY824YdQc1KUd/YZ
aCJqL5YRUIpOBsfhpgAkVq3/WHVfEAJSYOsWNM4m3qqJB0L/fOuh/7/agv0P
QKCYjecfiF4OY4hSmlK3NkhFqUoUIrM4jDr83iAL7SvRhvtlVxK2SezJBA/X
n3PhrrKKsVJEvUbuOUjisuYugOuLILys45R3HC7yPp+aioNO52MUQpRnMAoH
tDMCgl1Uqd1Ew8DCwpThjFBLxUEUfX3KGdoGrx0qUIrTd176V2o/byCH1jB/
YEycV4udYFcQAeyvaPgY7xzMsDhKtyq7PNM7C+sjjYBeehayiupZuKvTZ8dl
VIdGzAqAnCogcGsJWPCxIg1KYyasCq1bJ6NwacvRpzZs2lewX8Y90jT95EHg
HSnGQcQ+yMHPxAPhsK8aa/HVb8fcWM7NVKABZX24hXqmQJJfOK9OFgc1NHMv
KFcbPS0J/zp+0TfufK19UCq01qqJcmP9Z88pz/bs1nRULyukYba08k+SvMQk
Hx46/nqNSTxdqvyNk4ShvdkiNvaW17rVAvon+N8ldkUrgjc0OwPZC75vViUE
qv6zua81+Sz1cCCGdcGdSIeYSOY1379LOCvw4qVPs4zaI6xwJ2FJEUO0KlSH
g2z3GtsbYBxhfBXT0hP2AJKKYO+4L/cdWAyW/QKtk3++cIGOhRmOjOkritGi
oslNfl2PkrOqrzorfHjh0BX/cgAicuBA4LFUbY8bV5lZA4yN0Hjj9BqE0H3g
VH3pFt9gQMJ21mBl39BUNI+SEPDzyZNPby5fLLU69dkX1RcitibRYPiAuVsV
qYoTg7s+R9Yq1u6SX3QP+vebkRQisomOvTQDw4WvfjpS7Z5S9jtIpobNtaPs
l4mu/IEMOTkJoOd89Q85N+YCOfUAkSq4exjYpUr6Bswzbxat3tD6PpEQh/qN
NfRMxGd9SmpY4bXdXE4ohRUKGk7cFkS3WnM1tu5TsOw/RaKLkqeKsPEz0nJq
w4zVFVBBNitWFHbvNqy7SAswmcDF/AsJP1xMMDTYidZFQIvDD8hHKD2nXP8r
WVGFI9JRxB0qmmVTdd3NOYXyGZf2pqut9NI2Nyh2dPwaIiyhTNUiHJJ3I9/p
x2CzX3agpMpSMhnS/jAMpmmRn0LHVu8kJoLsg9ZYb6O0dmFSjT3fj1ZAEFgX
rm/+wDRCteAiSuFODKE6vNyPxEPa6CVUz2iZWZ3XsScrxDk+v4GRpZeEe4UV
0kTldd9HJ0aLOt5eIwA2JM3zVQwo3bXoKORuAZomEzZbOEq5QhnWei/A0sWj
q8aS9gpz8O4o9LAv0nD3pv5sR96FNDElnfG+3TP1ezbqYeYAHdoJnG+jN1cF
SQGIzTdHrDlki2EjTDNOc2yabmuxtPcCBFSKo2QbiEaiX9i1O7qhxj7JTKlw
JCAwEkJjjplymQOztP/+CB2YONBOV2QzXF5wd+iVvwGNpTcQzCddJLaSzdzb
BRjJYAkRQR81Nhqi5/CVe7qx7AYg/1pFWC/EQux56M+BeEbe4OEFX7WNyju2
AV9wu409MIs8kWPPwHNslRVqq4K8cFISiviule6nLNCHqyZF9jE1ftdmMW6+
Kf26kYhm8kY2s8yjJu2Dt4O27E+Iy2gf4HXkqo4pSFBwXtxNMuQExkmeh9MT
+qAWkSXXf67+i+3ojHXT5fToMzAfz7qsCkoG+wEIFk+uT9TO/yCpkv7B1Fnh
0qhTtkw3EbHjm8ijvHIZh0ZuGG6wJVwLezCyirCepUEXCbjn/48fV7xxXNop
eXmvqrmYExhzECGysi5UoYQau/CKglWkvVtJa0mH0SZko9C16YKAeHhyCD+v
c27pZKSv9cOwUWU+vWlctVxhctULfA01TuMRyeYm8C/xXG21C56myNTgBsxN
QkP0Y2g5caSyuxj7c+WzOXLw5nl/I6jskARy+z8vlbEUYRPU4TEwmY2tkGu+
yeno+Xfv6schKYCJavU5PwWLH7HAIlX36baQyvE7nXhDa/HTyes/Fhw6+vlo
RBN8QY83IAccOESX28J/Bi5Fg7i6A1xbDr6Buvd7BeBbRVReiwRPQpl+pzvX
1jTPVmDWTCG8BvWjt+ziu5xNGKNdPZy0+Yr10ALpqfKFCNRzhrucZznLa9e/
j0iHOmHtzZINU9R2AbBROczc1UOhbW+ONTjW7b2i78YD3BObWs7QbHkdgiC8
fVJeXtPP8Ld43Mmm/750J96HL7Cd5Zj+0jDKyCkoaUy1Oq/rEtzJSZOC6qGg
UYhyg9xs2opQbH+Pve/Cfruw0VjQCiAvsvs6PynOAdAqBVA7KNTNXs7g6A44
2ABO1VG3+wRNYjlfpXLm0WsBd4o+tmc61mhKOCOUEJNdMiV8cmIWkErCLm7x
qZSP8IDLg0NlN54CcWOaVyLfEqTS057RioNigb42YWbBRcpjAyOEEXOZbuZE
4JsOEXGo1MMopiyccB1g77PZfgvvWrC39JUqT7lohSlrVNw7SlupRMTPhFQz
+VHYoUpaFBuHyxHGz1me339dB9g/s4HyLWuUT0tiDeoGwd1lshBF3myvQLjY
NWGA/38uXRo5y9WjnjVDz1pAlZVo7FxVC3vj3SsffZDWeWJxfY0PvwI22tnu
Aj5Azk1RzB6TYekNFtMKBGIoILFUFTTR+6SxSLOGVRiaXn5tyCwYjWImqGy/
XCin6aA82WkUd/w7ghwzWd1wWNnXOQ873p4DmOZd5aMuqxO9JKJjozu4fff2
KsUrqeNFhHW2qYiKybtHy11HTA1Gn/EM1tUHiermtXOuMaGwVkv5AZ0B7deq
G51zP8KXCP+PtTDSglHJ1N+KhxkjvlaWDPjCDdhq+1CL2PZQPON9MUD4rO9f
moOBqqJK/jw7t8o/wYZgOMIRC0rWG3GYa+qCeZZIIuKsu+b1vraUTxqVmP53
3R+2lVsLIZpubMF/legX1UCPfDx3LHL3L5U1BjJrzNpH9rq5jnkqYHS986VN
spMIleAYH0vfEVZsQmM34ODv+zn5fa98ybom2+Wqi2dqGHlKXWnhVcu4LNh7
D8SgLqIhlWk5Y3FDUVN8Zw9twzhFROFYxGe6eTTxcsYccM1VMSU7jTSO9Jg1
cGmH5XcBI3GaO+I1hmfV0YJaEz3S85Tluuz2gK3yKf4eF+jM+hz42DL282LF
hQj0ldwv8LKGUX8rKH982Zm0K5Q5203HnzUpKIKZT2cX/sfVT5ZCZvEMBJUO
1w5OI6oV5ONt/gIFprtbCcUQhnUVGmcQDPu8ZOcVN7xFKLv3cp7uhaQb8ZiQ
xqeB376NMGkkImbWbT3ntNrKP16fdJO4EtJfoUjVy1y89HwSNUo1a4xr47FD
BfU1mTeh4ELu/0q12/sHI14IMZYvqXYfiquG154iWTIK+hFWFcydAtRryQxl
ar8vWPDORckzorfDrhTu8L8AB/OcQhBBID7pr/fJ14U9eHJh9eR2uWnjBgwM
ZIjshfufBcSmbTTQ6Db0h/JH6zDz+gKRkPk2693DGBAu84iR58Mr2oKUF56X
67yG86fBsH4eR2iEdYTHMBE7GT8hgeFrrlDdVLWWy+Vjv0WUjBQyJBXYHxXZ
MmxiuYXb5VkhEcjY85J8hKi54bkJwXEUmSaljtLJMuYVbmRDWjcdg6/aeuMm
znjvLHnRcMxI0036I3EYcHH4zHn6RKAhAcUZ5or0f0D1fKQiO9Q/UIv1Imyw
S4J2LlwHAbIKLbZYBLsxaZZ+XCFmx5HAK/0Rm8ud/MAP6XEZ6EatD8dj83Pz
gKRuSGoNlpn443FZnA8U5GiGnYbvso1XullXErjSj4TGUFSaqy693j1JYGkV
GPY70w8d8ySNIW4h9cccLFCdH4GziNlSnprJyhdsbLK0aNO+hBGtSnsluZpD
rFytlZAD2uZaHf3AFHpB4SSWmsYDfgkZ4EAm+RDzH122xB91ZH0OjRqGWkiZ
MkmhVaPNmjgkSYTu6E7lLaiB3QvWhEROktWMDMUj57N35KeO/+PPndeSps/l
YAPea+LjOJgCRbajb6psaCnglWn+xhM0jAT/BmBS+XAlJv+vPjXOoV4dzwSi
gOBZj9qXWKvGrAFkhh9Wh08w3aAQe6lM91kxll0I/CVvtpP7+gZi3SH85L2r
a42+Y++fkrx0EKsq+1jQ+bO27MUKpGw8RIngcTWrs5c6nnzWapcLy2RezOGD
HSgsHQL4iDdyHF4mYu3YDwwa0DHcV5jmC/4+1m7eGscQZWwWa/7BYrPZlbvh
wW4/mXlshDoA8bc0j6goOiElF290P5o1PNMkEtK4eh0Wm1LU+ishuMWoMcAY
COXPOi4pl/ensdN3L22GyiX7lopmnLVagoC429S0YWtdh/iC2dd6E8ys0wID
2OKgWaA6F/b59aLVRw3LcENbruAhxZIqQ+i2K256BGs6pXgdFq0voRPtBog0
CpJ8BrOs0N5UTzE/hWrE9OBC+IAu4no6eRx/n4qGLFIJ0Bu/4AI0fmzV5kUS
zYodocJskr+8NdDbDoi8PvT25XJw7cm2s97ydLuFJNo5iRTE23VSLUpVEzRx
rLyiZq6sE0zH5TOwVpyG9RvoMVWy7lnbsKCnT0JXrQttoIn+PlYJWZ7BrRSY
RXT2odZOKLziQmjVjMFj8BZ7hCu8XdwQYvH/b5wN17KvKft4SSu5vmfnM7Xd
u5Zgmki/hYoQWya+LO2Uk8WHn+/6Zq5EOTv4gn3PViFUzvW62rKxN4QCyjz5
MnS0axVSYKvunWISAgKuzTxZA9cAuXViP2qoh73DFLNmL44N0v/M14zn8PmG
IFoQJM7f4Ksx2UxGef5+OAIaKfPz2y04Hw4obh4Rw16JUuLQhYC8VTmZDtYU
ahAkwW8QyQIjneI1TKtxEXr7hCHiZck/o93C6djm06bUAf+uPehy9At78n5Y
G3mlakSExIigvGOd+pyjM3Yc1wSobMQwVMUbOhMrYefAFaoUQB5ZGXZvMLWW
9cFGnL6W79Ibfdh0jVqqQrT6lXZX0KynGcMxD2FWNLxPKHefH4yMo9tlEo65
gN7mODOIYJAYa/U/eRXRuYdrUXJrknFGI3p3qRoDurssFeIuI5/wiUPMNPpe
fznEIRkcuGZvsSchHJGDo11QtRuHOh94mJEVjspcTyxLvW1wdpi7LRItYPr+
+p+iPbevq0kNV3li/swFasuIdN0iTnstqW+h/C4Fqm16tUKiLrjwyIIJgcVZ
Tt/u1jXd9s5L4BYobTnZ32CLzYZXpX9CKEJDs324GN/x3z9GJoU69yAveTft
fiUn+UF2QStgm2XL/B1tNu9NF5eoOuB/UjxYPBDqt69I/xslY+lPMaC9b6/J
+lrtF5qMNcUmQxRNatt307mf4OUs8QY5l5ziKGcI+Mupy9SREJ0/lbQ4dr3L
+d1cno8GIEATmMjonsB+5NKeSMfFrp7YExuLY6BpWMCgaEdxzIzbAGWzl9JM
8CMaO7j1aUVtdceWM7VYK4hq9hw9ZVF1rOjVvaWnlrx0g4eT5nRMo4NQmWji
YmpWJdYn8rgVHy7OsJOMLzxSTAEQHyotCZJ8DL/X62q1obwclbJorCswARgM
SpBALj1eMajYp76F9fASF/AfRTzMOEpsc3ssHUC/u6RkjaJJJk4v3Ti6N+le
seHTDQE4WiSRcge0oxnTSqiRldvjEWMDiHQBgan10B4yLbqusavBRdJv9soX
uzP9VCoCAZ1zmers2QedVvt5iL8ZFh+DBL4b5VLod8YKLcD0h3ANjzeGAcoB
8enfoJok9Fpt9D+Ea05OzZ6kvhUue1FcRfXYZpIfhFQfa2GWeVJ9f2dW91E8
G6G7oJVoKs6dzsYv5QwJVgGThfXdn7Odi9y6jufetcMzHsvBk8BLpvNPFTFm
nb0W8LITOXnyJBOotSvMcUPq0UL64prIvwN/U4M396aF8jT5Qe7lCb9WaEow
/6P6cXmWKrLwk5+LotUHJbUvEJQOfnGA8Lzz7C3bxI+y2+GT8dQs2dE12ZpF
QdJ2v4RHLLGftFrLDiMJMCSigddm5sYtpYUAeLO9PfOHy+9gI02zAxnI8EoL
GEiIg4+d5xR5rVkhlPVpm49XsAMOttxrWHBpGOs+Qn0bAceO4ETPXUs+13tl
I9/RA8A38EgQ1zsUZOANKAi/9xKxDKzJ/LP0AVaZxXEJyBI6yMmeBEQHOTIS
4Z49wYQRR2VS4uf791ETcXszSGQqC8z1rn1kljO4XRH1SbabuP7FS8jnGzok
yQP3PPpDex5ER6GsiDyazY4Ih+E9HcqVhWkD3NySX8ZokrA8JqdXWcPtTqqx
Q5/myCyOgG98rHGjC/dOHFREosiXDRPV2TGs/pipUdK0ephyzB1mnRsLh/Mi
v5zSUdeJu5ZO3q5wCQ15ZOa62dD4S4YpUYKR7Ug+/CNHyvnzHnJc6b52DdGS
QOC9Xf65tm70Uao04dlQO9zRXb7whW1mkHVNvI/ApRkRdr2GfTiLoWD2MAYS
YpDqqav7W3Cd3s+e/X5BbWzfLWclm6yNDAxi9d3HE7ndnL3PteyYMjpWaT7t
1fBDJEiwWlrr49V8oWyh8v4woTNvDW2yfsWyUDNpNObjZ1yReHGSmocUjtsx
mIzfj7PrIxeLyHx0m8h2jd2e63yZhopBbSrNADHxizajkUNxWsrP33YFcfia
h0PnfBQx7QvQTr3MgthlOAdhM/vhic1g5QvpCKDNBQrOjm2TilFlQ9S+zLfp
GM59sZ4sXyjBcTjOT8xejGgV3MRDY3ApoPYhnGFjgEfyP/aohMb/BUiJptx5
F1R3fIbTuHx+pr/5IhlgtjqaaqD12fqUB/6L80PxADq2i6LhMJsIVS9WVDtP
Pe0wMou2kLWas72gcrHSDXgRm2bhVOpTTn9WaRqBY7zDKOrBEaQy4a+VPDFy
jum4KeQKymWre9a3R3Zpqv2fggJsCW8cgl7qpINdUq3etQxYRo6caOSzV48J
Aoap+b2NMvJ7y1UZTgIcKDR+3ck634429kegpRY4CX+wMyfUG6chPVzJEsiI
J7IosAoQUncM6CP3T2OGRJ2wk+U8h383jKTsAYHWC16+HBXtWK+Uzt6DFGqB
k3pm+mx29CVwD6X8E96YbEqy6QdSaEuX7qmagpg/KTUUhAuydSm28GklzQ4j
dI2oqVv3RhW3EHdvs8citEH9w22/UmhiJ9RFfRj6uFW3Uy5gnTZqGch/HyWo
tkbS5N7AYf/IKKxqYHWV9iwhsi4bm1SEEmf0+QLMi/LJ73aUndy6coHQciWt
d8AzYBZXWnva7AzihJBeQ/8m0eM6U0Xu8KVak7QK/gVaMDGZgDZB4cOn3tRN
UzfuHYnsWac+/tXTOhNZfqOrbmWlCUgiqpoG5uC+nazLtOJMXNQGRMdVH/z5
fbZpLbwo/p+5bJEL88PuyyNtA8sa2t97V2tY+CqvJyHy81Uhda+wvyopKL7o
zQGgXWW9J1IFAhasjwKYxOwDOtfB2tSF/qnEtOmaDJctLvNyHLEe1zYXXCEo
YIvxYpB/qEhxxX4mtdMFBnXszmOLnwLsu/lAKTdqwb8nrKwIdd5tXRvJ65SL
8kPVYpCci9M2gVg/pMxObeeM3WJ1iG1fNJQ3TNbtN83hfnNI8Dp6dCpcpPFN
q7DLWao8qZwGdxHt7ZgNIVPhc/wDzAB9ypa8BXTkipn52ZSwK1O2+6mSM8nN
W1y0/Gt15THbesN6zFoAJlPrJrLGdo5/UNkoSORF6y2GYmj+Q6EnvwQJQib+
vvYxNhcnYITJ9NDK0MqI1+s17+SCQlFDrUAFAxzsx323JRhYOkV2EI2+lXKl
ZAx12e/ICR1YW+w7REwhJtP1Jza/J93oh9+vXt+omDAohQei311MlKkVYmfw
89hybHCEmi2fTkXB+fjXeHl3fgciqAtaBn9U5+3kncJnFcJwmKQJHwNQns48
yCtD16GRcBIO7eWvajUZnGpEbMPElgKxHPv8ooWcv3UK/qbzK95IQ9zwjm7l
Ny57SyFb+m3nGTm3iXGv8edZ/wTTUET7bGiHEsMYbVXGT+SUYb2OtllwLBJT
FR44qzRlt4Hwi6TVcd3qs0qEZSyp1p80kxKcO7KLbMKCl0faE3u0XDAb7xCv
MeA4MnlMZtAhWlBB4eIIdHL1NKzQ91FwZ0jRnbPrdgbC6nYlfSLKGNkx4Cxl
lHy9n9Ci7jOdQ12VRiCTcmJ/WupPY912UOIvfrcr7tNKnCK/kxCx8+OJiNBO
9oYO52oTtYofZ19cjBvi2EegvmacN1KyUOHwfks9474tYL1uM1+yvTW4rgsM
ndiMKW0TzgSBBlXn8dT8w9cN6WBfQPdZwo29R0vqpkqAtCK/CtwjZIqM4FnW
l5/0WNReDtjETHHPY/3C9NukgBGwh3pEixxPR8Ok4Q5w0umEF+d9hnzBXNHA
aVkC3JhoXckhUSIZvBalChaVuxx+TrcS5oxfXGG89bgE4gE80jwoZuZtNFud
1dgCN60hkxcrh9Y6KOihOXuDbHqB8P1MhrEy2ExASlv+TyQ72sV8TFqfZH3x
SVevUU4uajK+L9c0Wd2OKT2PR9bff4DenDrDZs4fj1kWLtXw70FVe5bD700T
AK5dQneG9pxYqffDMpmvZNp14oTN1C9u0ztYhg65ixXo8s92ns8xBJ3Ittzp
KUUjmGH74WFpBWIYvfboO9MQF7uWIqM7EdAgmwUgh8CYUZun2CMYk6Mk9KKP
fCP2hTul/r6pP67DMgJudC7GzZmKxwxW+GdXxUSvFAJO+yfrCtMbY+q9s3a2
OYnIqJnRK2WxtRrXNkkYKWj2MgmrOeQeU5QHVcrdbjFNBSsho3ZLXrq+ykA9
dg8tg3K6Hne4gIPa92ft3P7FnQ6W/1OpBXfYuIUa45G1O0wMqHISrNoSvHud
XR+ShVKrI7d2teBMZ5/U+aWpkyifl2M+HQyRgbB2si+enJPcgbiqLqBUiPIz
GmHChyvr/wESEN7TnJCEwe4Klbtvdtj8dt2IT2lhsFUX7KLe1J7z1Sj2k9E/
bD3ZWH2Z4sP8k2hhzmlqLI4YaF41SroaXkIrTC7MAVT9E+M7V7Z41IJjYzl5
Bv59PKowZiE/EdRVs9JfMDPQL84M0DROqFpIhgOk0SuM+sydILCqowyvY1kz
Lkl4TfsopdwJ+4oN1g9EbBZMdSHdphhmJIIOvFy3x378xLuF8SrqGdamwDfI
O7eCzGOWJGquTwLFGvfX6MfLfPxNaGsXZQkY3kLc8+TJAz5D0Par8RD632h8
ZivR/qrU9Sk+7Ns6nHsLI+bCl2cdX2nuWwbbgNjxndWqguT9G7Ly1QLKhjoM
3gwqD+mosS6KhOdNea8uINSfufCItt9iYmjI45N8BzD1+xSYEKs9vcO6TbTj
Qk2Xar6HVZjz0A9pQpvwolIRoj1ki/9ezsXl4tF7/7P7hZ3Lr9x93Tr+CHTp
sy8U8htrB+v6sAUDgDaCFJXERuc/1/FghHXocjcLShvPIsPBquCxJSgyJUci
1s9xGyVb4TuQeO/RiesR1ECQtFDLr2gWkN9ZJxEr+xPtAjY5o7JGRy74GflV
8/FKiEWYkhZgM7dxJd49K2/Y6LUDeL63JJ8lxMsNpEcjN3LITOaGtxeTB8h7
0l8l5YLjODJ9mL2oUbkQqgRVqDgniSNL/Jk+OcA9jMy4DkfYkCy67OCSaczz
FGCniaYzr4r1KR9ws4bjbzwfIpSW9ix0dV93PEQSimoOF1k07l+yPSl/7MV0
K13ycaKYWjITUCfprwf22xdnZXqUU0cIHWkJ7WAqTqu6m2M5be/16WLNWl+Y
zr7knwdfIM2CGudch8AvLgyO3R/1wljFh6JuTjPBbFXBzaL7iOJE1gkqVoqG
SLyDX3F+PC6mrzuhmDAQF5W0YTfu87HSvqjvvww3J3gBi7/wCbnceJK1jKRg
Aa3uVEa/SBtXRWqZaGOLTHoJADPT2VS1FD/zxkECU6fuT5c8a7hmnfiuVPb7
KY4zAjVaDNNkhqRVKMz3Bi1ax73HDaVC73PY+RrKXk3B7PMRQL7urAYGHny0
p3kJ0VfeEDV3zmbQIQXmx9o5A3vmSK4zFNdE8WMM3B1rnS5D2rkMjGewe7wv
IqqpZEY0Vr4hrbsT8rHeoFNocLUz9yBfZb+OaQqVsjqbdufNytqZEU780oJs
/S+ZWIwsIUC59PB/J7qVs9LV7sgISnllZO02lN5BFKIwy4ItET6pRHIGB8z5
fL/R8t1dle/JKySko4LtGEO9wMDZ5yIc2O79lqZBTO952zxsEJH1+aq0SN7h
cby2xiqUetN+ZV2q+UUqZXfG51XCJNljx97osjL3FehZJZrQ/75yzCopeFzF
Iwr/5aAwaeLYZvSL9JtXnyh19LJ8bUhtBhI2zqfde40sd/JzYdwZb5ptJtbT
gDNl2l4R4KcrGnxLNfPypfKv/d81WunwfRKn1H55reC2xWpE5vsGgAuHo0G1
mhDIR1h3xkBQ6r4kCVVKN/UOOICAajrq+ljS/gaxq1WzZdrzLQVqrxVIQFsB
LhMvFEwsZYlhv9kGbpagb/zzLW8pA4f6YqmNTD16ELnRSQGxtx7LTUpZkFgA
mRIWDzGqfatseIF1d+on3yFxKnPFe6A2/NVoiRGQU+kGtyDfG0h+dr03woGE
nymJoa92+0DmGt69BuP54wAdiElwZeUKFCbo0n5v+FKyvXHgs/A76pZwbHsp
wKKNqEovLV8LNmm4N/4BQh9PAJIYmFU+4VD03QFtdmKF9+ykmU43Ybbt2CsM
/hhNgwb0DQpsydCO0u6ZvfjHz3U2kP/I1x8LfaFoiFsLKQkjL5xwWNAxgsHT
8UIcf5zH941gmFJYKvIGBp/+ypGjMgTX0yJPqcVp4Y7jDi2DfrdgeDImfR7b
9lgbt7YqxMj9gkOuef4fGJHC5c687Y/anck7Dv3ZFrWmp0+jzTvJu+QeC/MX
Jv0jo2JfU4hWBsdqSjcXjJFj9qPmJus0bx6ZIrJ7a3KK04G5+6UXYkiq2qGD
wcK0xuOIxuruLEMkQ8r1RK4ztU8tAFz8KVaqc9Hq7h4KOeI1CbeA4ROs7oCK
LKt/xLJs7u79HyaGrLhdpr3PPC86OtvMrIBtaDQcMPKxTVeGhT3UlU9QuvY9
Ji5uoOAkCAcnM3eU9ChCfEVPE8E+L19S/VQ6txW4nNXLvQAQ/U/0+EBxZK2g
k7ev7bXYathOLryLeO2Vm/FlBjiqWLRoT++x+6Nz56f6P20i3fOIE0gXYI9Z
4UthLD5LO7wVN2/6LgTNCwzOJG0Ax0JeM72SqenbJdPhDLjaAMYSVn95mYj6
87bcj7hCCOv0CnRhtjcgS+gTEWO5CpJQFCUt0aOtZkTFwaHYTazZPPLkQCu8
qOgE/zJ4Izc/HOXFYA05oRskwj/0/Bzwhp26JWEFoz/mgtE2FNmPk67a8Hdp
O4E57S5xxowGiAqueEBZzhLAC4LVeo/m+yGhBShINVdKZQhNRaegP/Fu07Ar
z3UcbBn+7JVVN1tA3S2h8wkbkn2fkC6/P9S0rLG/6KjrY+wVVRfW+TLs2pEr
htphc1bzxg+GMtqXlKK9FhNAVyEeZXQzLP2ShMh0k2v92MVI1GATwBAokYA5
T0QoNbd1LkiLiKcabF433hdfTHsAV2xO/ZaNHb8nZJYHrOd35xsvYa1bgaTl
qjuDF30Xrivj2MEnCc/MzNbyMztKrG2RdAR1sQNowVUFttWpM4umWRIRpRc3
ZB2Pqzo1hvnCyM8TJfShN6kPgwGVsN5+mvMHUVe0krEt7tWEEpxTqu/wYxIn
sKPCUaC1w7jLKAXRhavbaSdWoBd8W2/vX9/Ju2EyEkdS6MYnGzlKkUzy0awE
TTmDnn2icIrHhIbuU9cxqeCCAixY2oM5wSz5eEzwiec3mj+icVMl4X1hNx9U
i8H2Aekbyn1JnpPyaSeXSJ8XDp8RaKLMKwYrumaAwnZUF9KtXUgBasvK4HRy
7NUe8WjdYqyBNwZ6D5w5HoqCUHZflqalA64b19s6VfcJOMQ8diGe9OvP/8Me
I6MxOGc1GJ2J0PNBu5npBfsd2CP/HRY8JPcrW9mDT/BTIBSwv1J6wPYzKV/i
j6RswGYqC2T1iwRGNmNpKPsxTBgvJmjSXmkjN9/kmERtgvYCMOSRygiJBmk5
cqvS6Ezb9dFUWHVfo7EKkKKZ9Kde4Ori/Pv1Szah/ngkXBYaU01JTaJ3+wyK
FuqJbOuWDPKbwlvcddU4fkVjOcKniMGQyFPuuHX5FoYkPoaXwWaii/HQpbt2
pRK2cYG3+OJTTPOtDx0Nl0sT3cDitJ+/lLMiH44QD0ey7ER2Bhwpv25YuTp1
zQjNLOF3tvpGbQhHor6lOWduQHh2CUpuyhIr5GaN46JecN2cmNQoPAAwP8OR
VlPPOtTway4c+b9Fcowy4MWyR16wX/3LdCoopvyJsl89hPjRi48BwPX6KQrQ
a9XUnWjZ6Ccg5nckUush3Bk3IbaNPWxxT3/QBIkVG8KCp3QUAi4bSfwRAAwg
7C5MOXKw0aPQsEKZxondMvXXc0tX+fr1qY/gs1PcHAc3/Tmj5O5L18qWjJDp
LmrY0AAPJ5fjWTE6F0FhgBZRM5Y4wGAI2+DrX5xMvvZlZzuSuUfVM76E54QU
U3+iFdtKizQVtzml7jPa8N2JQfl69otBaXDB+IlguxK3ggriBppM+Z22WaCP
+R201qXEHv9xHBWbX0WvtOv8Uypw078FDIurADQSuD2imHxB4puYfNU8nnjC
VPWxat8NrT/saxj0Jgil62alP+/Ud1ByjxlL75K6l+0R8UCSr8UMe3J8Vjsz
cg3EXQFqYnMX2YMvEQlmjY7p2i8gYz32hT/oyjNqOI5KlrVLqeYE+uWslyUO
Q6woPfuqboSih/pCR3T9/xORi0nP6Dh0fIH6A3HES/jIJEBSRDmLTknzoI+g
7H1i5zQDXyigzEBCj4iBHfkiJ8VthhZuF1J2+3HueROS9uXRvi1h/AvSSmbk
uCitBIyYcUMV/+pF9golNyHUYVr4T4tHjWv2akrPz0zSMU+OUYvY3mYqZlmH
I9/1fjj4GmTqiThkkR2xShCDGFgrLQiPGJjS3rZVMJK+/+Ysktq4wLw2b8zg
sKsKcpFIX9WnewQqI2/5ZxRtlxfUSTZ8gAOmRE79SVunMfKIWw5WBZoG3bVk
maMOOGZ8iIev/HHnJMXHH8LbHnOS1W1QKwQJZKWUnu4Sh6HKe0KnjqTFy9s5
oyhBP41PrGFlolcmgACYK4p4UMLyq8uK4GJ+QVNUV5q+rGxrkxqqv9qXa554
l9lT1PS+z5Ja0yDl6CflVwbZJi+/hM2H2++GV4JHORfPSF6MppgAFbGzPHmY
3cYKMoe76UF4bQYxK4D0pdrHAjOg8FnCwkoDrv5Brczm7ImiUlzlbuGhJYEk
oc8BmJJmm4MHRcUUCOLTp4XPNyhl8YH7EJgpT+x28CjavpPeYURpYi3c7Blo
RTws4Fhx5+kl57KXASn5EMjkpsouD8wXmiJkGjHqxUptuUv/UD0b6ijK9b13
/GKwLNB9Bz5W7vPlzfn7WWGMOqB4RiJVTwJ1eqhKiA2PmR9liKHhiA9pyCX3
BwV5N7izoLNPgQZE3Qaf2kwz7nBYL2K8rbiSmb1DEWXyQ+7MxXNa11kVwCm+
helwXOxeYEe6KNuzsrJgv8k1nqWg6jHbY8qEQkgWQa+lCNY2mR/cDIxEpQzo
S64KXcBBpE2FNRsqyfGOH/rNMeEFLlE/nDCqaWyg+3Bzczcq1MyH6+Ol1mHS
E5oTXUIeAIT7F+2gdxA5iJBJpAJLqqjtECK7AKm7esEwNCeT/Xu5DulcHx7Q
1hd0G6ELb0pkx3TTizjQ7LJ/hwQ/W4G6SkcChcajHTd5VJ33cu/9kcLsg8Up
dM2tOBcP+jbn3tlA5ULTh3xBLZTkMRubfzZ1CxXaeuc/bYUIp0YKsLeqRJA7
w6rN0G1y4CLIqbU5lrhJ1KHAdQdO+x/t5WEFftKtehBMdq+mczWgDccwgAB+
XWdPFJEUni3KpGg8fCP98e4DWAt8aLds2RjnF2qZ85TUnOEZ9bc+XWQ/RluM
7pUdDlbaxz1SGMAYJPqDe5zGGGk4yxxBk/PmUljXP3ap4rkG4vPSj3+nRtbd
qO0A+Xp4UbokIAlsXnV9XZHFKiXV6jn1nS0IrYdHKYMGXhPm8Ps5IVuwOINU
OaTBkRdRVgWP4lSlL7955WhvtNhphHYhN8HInH32XshQq8pJVaEEpaL/eML0
AYGSxStf5YL09g6lLT5UHIpFCR0hITph2gBE3DMbbdLndmtcFzWZVI7qmgfe
8ps3lsQHXTb8kNYM4efUw7d2VtUa+mWkd6XbpJc1xCdw+mUmBYU+Ogppoww0
oDuzpXxuSMB4XQAO4t5IBJPIMpxxeWO3WdUn6beTj7bGaL38f0xCJjtwoeVE
nDh5CyKkCN1VPvVCO3cFNChqHwI5IOvxmr0LeIfPPYMaTniV8aorRiDtctv2
7Fxo6wRrn2IYgbIa0LlP84SARNlDBcMiXLyzmQE/9TvRgAbdsoPSq/Q137pa
A7fGxAUZkHUWnUTrm6SXekrSBjY3DxflumPSvc+s0JF4XMtt8sanUOvjKFmA
rKQg5cq/zTnGKvPqJ//rEOFWOEHZfFUraBs42MaqASci0swSrJWQaFUFmwUx
KyBagM1MUhCZk5a6mg6By4iQHfjFG8IwRvrs030y2ZQ9FPBoIQu5U39hCqBS
YEIerK9l+Ry3JHy4KkFd84FYf9SKoJQvgpkeX54FwU5Pl2Z7auWF+l8QHNRW
gIbj80e0CH1zZ3XcIiOKYaMcZ6bxgNAOzNXBXbv9fSRX9Ojt+k7Dc1DB+Fu4
WaAZSkIvaVr+RqWMA8xQJZlIy9bJLA3Zkg0i9DYyQESeLeKpIuI6Pf9R9ZR5
m/xswIHsqnx3HyTty9qu95gbaaN/lptiyMvsio2Oy8BfsRd8BaeWs2feDooL
nBl1075QAFCbrjxva+er+ChBBcsZ/GzI88TYa+lRpCwwEIjovEFrlvp/JyLQ
tv9rmGLfmVExHwj2k803hw9hl9J7MBOA3Lyrm79xbLAmLFTxyYLtXko/o0WF
2A9hZjHSZqq7t7FND3fwUSMjjqN0q96UttQON6Qy47IPcg0n+H+LD36+yUA/
nE+RrcB8t2tuX26a5L20ADC4TRhfvStFrfmxbTdfW+TrTMOxyOXfEZEkt0LG
jE9OBV6G70BXyJ//Kh11+TF34B7akpoFlpIiVsyUZSy1TuDpWYkFYbthBMDk
1RgQ2NmhATN3wyYX7C0HLjlBkChGbj2YHfILfXyMs0ZP3GBgZIR0vDblpvO0
yBbv2FHqRW2csJ3nCQphexY+PcBaWXzCCx6Bqj9MLx829JbXwyYcGsSUsZPI
M019Tglm1Xfm8u7zlPyeOf8SOUrbc0mUPZhBS5j8EkUiThmqjIEPdF8qswMN
XoYHTxpmpA9zmoq/rtuwS3MoQEig8257A7MGaK+o4JNfVyDgk/amPfnedsr8
/G/SYNNk+aVHHpxu/VE/C8ho1VVsG0PRs/XItBXIYh9WYag5zx+eMD4xfH7U
O9hGEZ80a83YmN8Tq3TeIg3q5vDksUb2NAQepNd6bbmCUxgqC7DeAQlS4/mD
Pm2Klv+B8NF4zHu2xaqB8SuTaiQxsDKSXMI/XZIErbcAO7VbsZeeVbD5kbUK
TJ4PJfGYSw+gFO3YYpdUKDtXz/Obpfk/UVXTJHZCm+zuKCPCcJhfhlrbMndY
0LOnMMZOe95FwKR9hKtraHLkHX+T7QTwppatl/gN6un4CJf6n4PaGMxk7Ysz
SCrEZIuu5tHmEn26XJHxSNd/YccdCTguG2SCrQitKNMU5BG9rDFgHr2Hwv+b
Q8QHir75r5VUqesXpH9NfVy/kDhWlXqprzYoJRK8SBxgFXq5OtJ8kM7MdNYz
nFOTvFLLZV10xmURr2dBhQUJGRUdLWY2b5UNpxRR1YoCMJ9KW0FWpNWUCDc/
tEQ6DaD82/4xAek4lkm//hcylHeBNZGjNI/RkZMQqt7VEsAHeA/q4G8MJUTg
EO6vMwaP+uNDSPFmDN6jz0zK6V6zivETJde/Z0p4o5IGX/SeDp0/31WuFUY3
Lk9mcNdilUXDGjjb+3Md0qB9ptk3n3khUfwkmjwONHbGp0p2dBbzR15vVzm8
e12jX7kvxYjVEX5UIvUh0OvzdaCz7AJSEMF+YkQ4YKUazNyaU8aVZEWIf8qI
kTSYUf5Llh0OPJ+kyKEP2RMhPgfGF8dK9aLNdaWIklVEUglGWTiD30WFuDRM
7XKXV623jbeyMyOQ2F6NL/MKf5y3VjRCkv8MZC7ODzvxeLQjwgtVxR1FuBu8
fAgH9iPTIOe2AWZz9wioPbORs5tbdu/+K5WT7iZsiU0QKR4ASHKj2WwVOm7k
Csj2+MRr4J76t//ONP3sKR7WQu2/GAhPn62cu4p/ab+YJc0rFoWb80S2sPU0
J5kT85gk8Gy88SOTFwHKJLK+VjcDtlYuY55HTG1012NRPHNFSxjy/LpT76z0
LPpaWVLm1ZVswm04vTLdY70zF9sUBEG/U+yISqyaCqxJihKHVHfUoTANRwdt
2+m8PMPZ5Jc/+51241C6qvtkqmLFtiKaruiOxaYGT11ApA+LfLpUSeO8aDhd
JH8ifDPhf8uwbwQ5tF40vilsjvRGmrTVylo+OErE2nMqTVASgxVe91LonWeq
IbpJUTfMQXM9bjY9jwh6wPyXbvvPgvdPGHlme7EUcy7+GIx6cAPXsmSvNPBI
JwWRhm+hcesqulDyRfkHnQ7YjtX0SQJRDcTqXuRQcS03UTb1zkjiB98COxF/
f8ynWGB+85XsSYvivAegBjkZnOCRKj0G5vJmiBaFUhByFW6sLdc43cA8Ovrc
CXS/2PtI0kt4oM0hZ7/ko5nfuyZveVLDmwPu1JmL0dDea8+6gC8lVZzqpetk
AZZu7WbZuvzA2MC+BBCsp4iLl1kExOTomQmAM5KtBydPR3fDpJi2+LZj3+Pe
I4DNyTvByyh0VIXW9gLVyiCpILPVAZg2bVfa5BXP4OrpQlLzv21tXSN9l22c
N/A561s4ss+wSv/OFWOmLJSihKFx0Bi7rTsq532rY3AzSJnsGtHyQlNWjyC5
XayV7EGt6RKljYGyyzex57ewW6Lc8n6SQKRlKB+sLuOzzy6K3JyRYuXIW/bf
9ThtTlWn4JHAJtIzBnf9cMogAOBIMo3iLNt/yO8nw8MY1zyAdBGGQFomnLmO
dJQb1e7LFxlDK96tjwNKvCE8wkTmLzjgxWTBkfAPc9w9mJFm54djM7V852o9
+Vm6vw4YNNy2MQ1aRvLpt/cYClZ+thHvmawkXnMAu6aq6XLQ6Z0wV640r1PS
HkV1OTSPV6JaJ9c+3xT6HbRp1G9sNmHNqUg2vQKtbW8IkRLj+zKL639b/69a
CzA8LiShA1lHcHBjs5cFNIYf8pk7Cy2QmmAcFQyw6C6RVpo+Wcnxw+2V9dje
Q1JXmm+S24Ydkpb0qgXAcVBEJ5Sb5OaEE7D+m4Id1PDMAIZQTg+40G9xiZff
rbG6sGueBM5+m8E/ZnvrSGsAimy662bjDXPtVFKV+o+poJItG1LCOknQDOgb
0YUFX4DFKkqadR8e7uGAczHRgrFSs+ESwUJ3vIZXTjULYsdEV+40VX/C2dXW
59WoCtY2L6zgEubR2t/OZ8tjJdFajetIEnaIrYHiMn0kkAaafJQff4XPwbq5
SAAsZX5kYrwoB2MA79a3+hfDYpqVK+quf9AccAFfBPfQquMY80TvEdl1i9+J
lWbcLazg0ltSNqcLIx4jt+bhhWZcX8Bh5lCluesEqbw2mogEMjVVnDJJsGAh
hUMxp3SnydV7vTKHQc90ouuq/31MEWsOOKfU4NIMQSehDJeZcZW3eoJP0KT4
pA3ULUYZMstuFd6mTw92sBoocsViXKygO+79vPSTT+rdOn5REhvdHujAsXLW
ZqEhaClAfp6wFnRZF4xmgOAf1BpMxY/sYnQUDapcWLCIcGkNQv6TVU+4iVVr
Qz3jAzaSC6atGVS5pzZxgir0O25tKKVjo0KUxOlNA6tRgdvhGVuNRdvZlfRg
+B4mEnplkSt95Md4SsRnDHFHbbwxCsz0BU+zvykLwi1ukGtriFHkEFvSECJu
jy7I/388ZN59lmtW56f0C/JRs2wJzaHWEKWD3MNwhH3FPlL+gYyN9yNZUDMN
+iWwFvJdj7JtjzveR4qQZ+mPnc0ehNc2VfvZg4IEFmWv6YYzqy9fOvFERM0g
l9X5ymRPPVV8JY9Ipm12e+7ToSENiGJzZdzczDOD4FZy2oKwSljs7jo03h9t
WSNil2R0Zg0rrTzu9pM1RJU21NuyZTrmtU+ktUQ0bEzDTYl7/PeUP38++h6x
XmPGurMOK4AtbKpi2cxZSHIA2smi+yHE2sW16h2q25MLBPmnr5UTpPsYVICK
3XIbVOiszBJRgMtUgYaTu9MJZYeF3tcmtiCzTuM2Dg1a3UyHOCbD3pnlDV3v
+6C9rxWdIndcL4AXrYcVzj0fOox9cOyP4AW59kyLqiIuVttcnliSoRp1MhT+
sVn+QXe+9BruLwtaHEQbcgd1f8eoS/1tBxCPaqrKVU8Pp+MKR8cROeT6KLLd
QaHpyTWjLR7Es5X2SetJ6C+XPDYKLZIJ0pCSLdVxHm3wRDHqPzX0xpHllr4g
nk/gdHdQcS118iWvFK4sy86tF9NxXc0q5phf7J/6qDHkezXEQ04Rxm5qa/Ij
A4OlQXUtom0MnbDa1n/powX37iO3KGNMKy8wi8NlPfc22efjOhPTC26ywuhk
5k5wAH9abWN3Ux28rzIasLgINqsJul6f/iOoqCYmsxaa0z8ogbcZa88cByU4
VhO7L3nYZVMLlMXtlN8EGAtymBGM4PumuAv15NV5ckHF+tCqPjqeqc0s+Iqj
xYc5mEYEOMPCMyQZLhDn4ucXZJ/mcH8/lo9hBzLoYCsy3D1/SGFItnUVI3Qn
YBJ5FO8OdE0A6l7oqaet+bqd3IZCSbxdvmW/6qd2diRw+1LSTGZlOqJm/1M+
chNgPXMjDw5H6QrTS4Q/QFTLl+tvg1NRdSv8Wc5nq7i8ZQPqo4c53VzFKEl2
WE+SewNPgYj3qcxQIMLBbxhSRoRIQ3fW+r0TvYubdK1ecdqpe0xbeC+uxDLp
49TRquNsYAxv69tyimjiiLgA/pZ7Tx5rN/oj/fg7utyHZO+J/VUqRPgRiGo3
BjI2FaGPjvwG5Naa/01c9n1Xg7apeFoBa2gafNkWRZhqj/VJYQPrQvkCcbcu
J4iRDvIJvXNtlRHhf5QbLoCDyir355zyWMHqabvT80Hwv+JNCPLRUktiQ7dG
DbW+ewNvg+Xz0G4wQF6mXhXF1k484GQjtfcyWOIFuqlR/W69dl+7GHQI6RQB
pD6NTjcRO985PBlJU9EtIbHLdCLXwMR5HYVtuKl5VG94lvrHTpO5tKqH6+Qc
393D6TA1APXuDfcq0XIxHZRpE9+oIKWPlDiLAaEtVyeoM5XiG0x9pvvAgvbm
dCvr49BnhzwW5HfW1TilycJJyfkS2zZNm6eJwlmP6cHIk+2GrojfmiPMtZ3S
wEJYDMVTeHM51WVJVTZnsv0dx1ZaFDbnt+1fflZQ+w6a4A7f1DSYUznf6hrQ
zsv4f+sgLaK3LubJnFju0faMU1SrI441wlztoJMUQPIvw1fqmBWM2VR7jGyr
+LEJRJz5LX/z6/0i1JLGJylHLy0vEN0KBV1EenhcIqpyZ3Pj+1Uc7odUKfRY
bnHA1vaEq7WJnur2KXGDTLz2xJ5bUQ3+t4QlYbuIHfc1YvaPkj+U11o74yUW
HPOTrmoEWvve86cmiW4CgobyhzHq0XXwJy8GrFBbVRZDT5bLHZOUqN37uAZJ
ngr167CEhYBmNkuDdrlbDwsrMIPjv4RumsOjDyE3Eiz6+AaV3T4LcJ9xC62o
wQ0L98cV2IT8DDyVJeLj9C8xOvXxMi535ISc+/bhYhdm56o6A2/5OuTvEDcc
eNviJOmGb+zDF5v0XWsk1JxfZvWQKn5Dgb74eTLy6daiDXGJw7idaU/2QdBx
ARVr5kR5u9fjjtbHQcsDuIq8qAmehruV0whQz2NJO5BEXcozLbRa5nW1guVI
2GBfqlpHK3jfdTV0ylBTLR4q0+NeufXxeoszExAR8TmxqeeROEXkMdDLm2qh
Cg8pAS0WLULjaFmVTVRS9ITK4CJZBahHPEH2+4rVq1nIpH/Q0UVC4slcW43p
W3NanwqKQrMYk1IdUf9a84dynYenLVvAyuEQN7fNwgBcdXqQJJmFfsKcOzQ6
ruxmLEZn+IGrMD79i1+XntPKVGYvcfCuGaahzLNohVG2E40Bm05JS8fIMsYq
ZXpYITtySLH5OaSiN2aLcqL9CiQQ9NqcHNcCK6FL13s4M/TqP4gPu6rqDQu8
RkWT7SHvqIX8V5apvxn+l1hXcWQhXmMdsjbDIVtu+umSdVvBaU27X0Kx2sp1
Gkw/VBVquAWJbQZz/tKTN/Qbs+Mv3Ghu/zbHbQEcC3i4WN9j4+QUuttiZ/MX
OSravjAu/zq/btmWsBxEkzG1RuhGYUZGOn95ny0LdVYSS/Fib9w0izLlaF4f
eOKb6orJgt/ifoojCDYbet+DkmowUZouA+h2rsjjKXaK3Kk+GLnejuNfOguU
yNsLc3jsDsLvpLJUP+J6YkZv+q7MX+mgehK1XYSxuTuvXuAbvL/z+h131D1n
rAf2V3mioSA/esap3+px3Zw1trRoXr4z7D/QrBOYFtA5hOOrY0tChPy1pomh
HndjW3exKOSp2kv2g2dijGuv75jMuqsPWp0cpitJpDI+6NKqpeO8I4qpjTNF
rlcxMk7xYjqJu+JxhcPWmCjPpfKwHfqRaBFS2DnxIUX6/cy73VZwLyIzOT7h
1iStCtJEO8D5hVYAumrFu0G4KvM6e2HeM2LOVvlmcUN8lzRvviij7lkfSzH6
IZWsaHYdTsntW04DCF3VijvNzEIG/wTFfhYbap0sCi1aaXQgGvHrdx2XZGRO
W2o77JZHw/gSO3Q0cGXBy8J34iE+woM/VlqttoahOT9bxavHLf+sCTIgi9Cr
QQIgst4D7RNyPwKEgF8aDTdvYeo3A4vhU+9t8udbCUyKX46iOUrQBVTn1LL8
MRl/q4U0nzrx2/9YPcuymjEPMdrUol5O1xDo2A8RTK4fgv1QCYLU1jjPW6hN
tf9BsySSu+Gwjty47jwfSDkRFo8Ci0GTo+RmOqmlJXJW1kL4VbvjU6YRc4CM
zKlxLGMHkdZ8a+elglbLDBuky1QwgLydPkZcUTkwz7I5WhjCT6wLgv9VjsxA
W2BUANRXQaIfm113qSQE2cafNtuEhi9xuuddsGBzxHqExYKsYXZFP38bc4Lr
o706+0rMptuqtJATXjMsMWmpKTDJMopPoE+9xcWNdK0L/Mw8rBvMV/e3qEpx
mh/rf6dTzmFP6XcClLzBH+2i0TXlPUEgJ6MGUEpvN9Rt6rOlq9ZCmaFvTioh
YjDdWRH5m8QZBSjxZfJPjRY+hloJEoUw19+FggmSfOVUXP7uqrBeLmcnoUzS
WRKr8QjD9YTjG/z1sCXWpO4f27/Xqb9D3OGe0Nd3sasYQhDDKwysiXSde8wv
DWIhODlnbm95G4Y+HGjZZR3ybFo6+2BcvyZ+GJhSkFEACzY7FsfJfawwMiLz
HMGI9w4tZsmgB+IBVUv1pxPWDwo+tGFChHKbKDoRf80XaegWLTdSro+3CDCa
egaAwfr9rDAiqavhh+lbCQIdpwLDAe37CEeOniYYsykTuP4Ka41rT8dDxDS+
AOWOVoA8EGpzFOXUJ2IhWlCBo95rmBmeHuSdN07Df2UvCLhw7D+vXK9sr+Ng
pBtxpVO9KvUobOomwxO1Bp7vAy3AHY6Ebj3yB35lMS2XUKZlPNb9nSEdZxgh
rMv8aHutyDfeOxxw41/acBlrC1ZYGMuB2shWHr1F8fBhi5ENqZy4SkZfqB8/
oOjpqXvzXwyaCDeNuxYe96JFkwOjI0RIMrQMUYXZH4xIINQhI2NAeBKcShr3
Dct9HWujnggSKJzqRK8PrPEQeHOQ/6DAMHnm4QgjOtmvvqSMgUQOx36Whhns
oegSZb6iDcqxGscOTIZozNFR4oCesOOTixAkEw9xXCNpE6enni1FIAwIqwG5
NzSBFGCVrnsiPR9UckA3ZDcSiR76zfsDWx7b6FjpzmViCq4ZSrzGZPo2ivpu
Ig5Xr4EzSVQTka2VpYW1/ueDmQ+JQnYmxw7/n+XTz/MX46zVqlPnWgOA7J6z
tTvxDz47AEydvOjBmHv2N9IP+N0Wf52F90JIYNWH+KJ/K2X4zmaV1Bu8MQMn
oYDsJwalh1XfNKMQPd+Rscr03QZ6Od393gn5EWeaaeHwMaF+FAn3jpp27BKG
f4MfSkHgQzK68ewKFT4ad6tPlT8FwYoRCCkleqvzsIDKGHAss3kqcJGmW+AR
3VKVvQ/x+Ey1CJPDvB9dynkN1Xd5jx6obLChakPkB5ZiCneheyASA6uP84nA
O0UsMIfNkz9qrNxNil/H7gLvKGAgwQT7pHZiBUtxjBDgBGWalp/SKO9SBpho
xsP4jAs8w170abQ4ljngAFfE9Gg3N710OVqX8b/Nw+RnYu4wlKHl3vpKbfZC
w5SXjv9Hpwj6GdfLQo0sWpTYOAOSlVvbD8U4FdBqCqJUEUMA6+I0Vc6e24Z7
mDOlxsrN+wVr2h7meUlN4soed/3ilU+xHHBMiHR/dEo8pW6kBwU4RPWrCBWs
5oTNJVM6fMelMUA4w7qGUrvIBrbUg7Tc0FMIVp2kQV+cKqbCy8kCiupi5w+T
1QoLxW7YD6IZei/7wMmAIs6e41H/SS9TPNs4ygCfWwIXxD1cUmRYKdApSa5d
5aRvY+3HnPpDluY3+l2nI1grdAzgbxGtV4kKUb903aC2tE185bscNmEctmCT
hq1dbZ6yHStr+FW4f0rmA3FVep6pR8+okFFISkyMxqTQk0qgrKrDB1FaNP7q
dH3i443Wo2Am/1DCL39HCSLg1yd4ZjDH5YQsr/zixx1sUdVKW9elvUEgZI3Z
rXWTMT1f3Gf7Z/gbUj+aSpBPDpc4myHx7X0qOIDV0wXeqgjtVlEBOnCmfzdp
KODo188zPnTXYnzXQUCVkHQnEuJ75gjNTsdXqdDWrj3rH6vduxWEGh+BT0uV
I9Xd12TXCVPwkUNaF6uXR55hbWfgJmi+BddLUwnqC/PeTDpcmmb0fUzhXZI6
YPXHBAsogUOSlVJnBKB16v8YhkuwykHZMr6OS4X9iXCwlX6MUj+ua8HZc2w7
xBVxXHz/mQgynKRyLmaq2Yz1Q8ZEUXwzpJcwIpz0xOEajS+MgeIUVnISfx7O
Y4LA2c3dtythGyxcl5+CnuSRrNoquG18IsZwlqSM66JBWbH6MA3FZwb4chey
+pca9lIytHTK7Lnb7jyBVqQdm7PIuxiMT8RcoRp0hUfOX9O/VbZwsQmfTDKJ
KPOcEvvqemFvY4ebkMEkiFV/DjbMA80QwWpLARjFgk/ZQwzFmt961bv0HvjH
wHnfMzWiM+bZyVMOrxmWIPRS/+gb72/XDruTSelinwSKQfvMwg0DkygTyr+r
3JLuMrLwDplMevh13HQ5A1BaiTL6l6daKMOT4jkuhBoSUY8BzyqFpDr9VzIG
GoH4/b12YmOi1oyMAjA31zpH2sCaFT7yjfwHhBn7O0deZn5/T1wqKvB8+m6q
17xlEkHYaOUk3F27+TStgjGAVyX9cHcFbAcwJJcrJ6i0pS1Lzaod3pxq6qZk
ThPNbRhUzJmmGpAgbWEvfZOeTOeLnEIJhmx+F57QyS8Wn+L4NWFLREj4AUVH
s1xnE2+TFb/7OBlX0dFVTsR6EA7L9ttj+BHLXVx9lS9LeD1U37XdMiIiVxkn
8oo4a6peE3SKz8AxCIz8gl4kwOqQROv1TyEzelNLw4H9ZUQqFAR7G8CRn4cf
Jex0V41CW6ew1XFf+zi0MtAN6qDMuBZdLiMoY7ks5bXCbIGhaHdcF8NZ3ZXH
K6GUZfewZciVm9+Zm16ZnPYJKFdgp7BLHAcPVRSm10I1WI6Wq84mMGUsDIjx
q13c59CC36gonRWF8K8jvxu2FIlxMW3VDONkpPlNr5cULFQ2uggjo1ttZpK7
r54iKUO49uipl4tDAto1lp5WoVMYy8ijFgFnFsqgAjFNaoXqwFpajuRHRlBq
X0nXQ9JtbwvBJHWOzWQI4O/T3DjZJuiu7XnXyGPeWecuAZoScrBWFTqQcWbY
q9ETfi31tmhglYzcZ/itrlRGn/QJ9tcHy+SjltSlYVka6qVgEMlncMJd3I99
RYD8SkBYaSwnkUap7qn38jsHD80q5cVmHuxd7P5EdaIKF1G2tdWpwNWx3ACm
lz6bzCG5lDzUN61yzvF5qxv0B0GE+0kUcvKUXSAX9EfKVvOHscAXOjxD25uT
6gd9Kv+JEeIBDrE4XfRycf2/C9MzEww7IONKkjZs/f0SlNP1gdCjBOvLJs8L
MhtXSQfW0cxakAASwgldDJiJHCxYRbuue9+5Ev+c3/UkzSwaI4NWLjlmFTAr
LcvRST6VKgw1NwWmGiS+S0c+2E+nt7ZcqKyCvsiXDaCp0RJXslvb+n6UUY1b
6JQypzCrGQ0CfIYoBenVBIs0cTZ2/49WPS2vNwmlOYpPHAgueL7awDOCW76m
Aty8QuuP1jfusgGsVH/IJPlHMd9+Kdi4r5bjL85ZhEoMOuMMbb72cyVTjrOd
2SWgCx/6I6EthxtTNu53XoVwF8datC2klXhi/zvP+ApREs4qd5/NdpSOWJkz
GARdBuq21l3Rhud21Qa+/j/xpeq/l1QDorna9LQqCqkAClPEdLEQ5cQKELb0
on6Uoqo3MJX3QwxsNX1OIgGKStNueUCs6DcQcq2pjPpx4nJjCtZ7iYGlaBUp
ad8flKgTX9Jfe/0UnJoT/HsPd+vClJQlDvqxIxb78oAUmvfh6FbAZpqw2VYN
M9CpASZyBIcFVPk3oP44wCH1nlfloltpqypLg3Z3rOyZpU1AkTosWWUnREcI
mlVDmBGu3LroTA+nJVfrI1VTz2QgjBgCLe9As6/eK3ioKVyFB+5GXPS4Mgo5
dzcz2u/Zo6eNbc9aGiC6RYMpIxlhzjjLna3aw7lHvTMZf8HAJEGWnR7IN/eF
nuIKbgXyM15f0zvRA/fWBE9MH190Lb4o5bMKqabsVC2bEg0qeqlGXVNSo+4S
eooRlXmu+FPVrXenevEYO8/Uak/bpX1VIMlm/1lg0Ihscf+NA6i8I5vktp6i
HaW6Bg8NYR2MWuntFqAUlM+VoXBDXMtI9/NCzQzA856S+bceAyOqBzc0htiq
2Zv9m3wAjtMraHI4UKkuwmQK8+8/WFxbAiTDLiJ9LppkVg+yJhHWOjsBSqBJ
7B/g5m97Q1VHS6l6kzwjuG8EjOrSJeydWgpaQruQipJ/xGG9+J8bVJV0kMB3
+GEP169DrZ04DD5fGJxGqJ/4YKM/OtkujKcPpn5rfsmfB57I5KaWnv0ERdxO
Mc1dHlwL2oQo+9pIM5wbp938trOHu5PjzKPNPu+rzq8JF9bZ8H4hO5MTvDmV
MDLGK5xSZgO89muWFVTkMjUljnKvZdzwj4cHEZs21NfiIYzVdyn79zngXIFz
vqPhNz/6LScJBofUV1012T2INgj0zpBgX+NwcqgTncZZ+NGKlftHyarl2BsE
7HnfEvjLQz6boXDTVz+U7hXesa8ZrnxX2BxnATJ0LQxZZV7uyf5Zp9Nw4nX8
n/yeR/uIY1+LbDmKjsxYQbEGP5WwOvmjoMgceE0DEUvEUU3CFjJeT2Wpzyhw
XAtOz46tJo2rTi99mpV6mgKdhBxaCyCg1LpU2G10S0uVtDZDBkdhdHOmTgDB
2TECExm3blkiM2EPHHYjyE+oNB72IfDSH1dveZwfaAPlVzHJVMLGe//jrFMJ
wTyQa8KY/syEo0pTZhXTsl2xKBXjCXPWjcTy4oj/m7b4QS05VuhkAOrwJncV
/qOj8n0noUr+PxvbSusSMcxQgHN6c8X6F3cV6W59fZ1GVlaUsgQbh+kp+Q2q
6x+PspFY1LdETWfGAMwR1QZAdMtMJJ02TXdhKWUKAHeH4bZXaFv9EBuNBWSB
1aCFtUyE25bO1DoM2BzRtxKHSetz25A+tml/a7a3a3VjGHW8BAAQBUtXR5QC
0WB5EDdT4S7c434OWW665kMxF3KROqZWjiRk1SnkKPiJtx1E62cdgzZQEIbk
JsAtKXuhX++l4y8y4Za9B4XMfWueUJW4+C1csQV5hqncjQlQcbPaJrIg+XxF
kxsg/3wWzNufKKBKhdBN5HsbYN4A4/SSLKyyu3vuneRhxMu9RKycaKQQK1M8
dz2NUdJ8QLHIkGP9MmVTnqOGI7lOIVb67z2jTQpFAGNh4eoYOU4HhScKpP/d
Sri6UBP/1/AlR8Tj0bthOfHexpwKv2ZTFiKsYTxw3ADBTFSKeqLzM2y0wK3d
h5pl372JPNGF+yLxbV8HWxQYLVKqaaEMH7UfW5YDpQZmw8OVwUDUou8ZgxuR
ja8pWJ3NMqln10Mgj0RghsqZgEhEGWk6eDHthvkEsI4gYFmyB40ID8nQSR1X
AAmQc3NdAtedjfuP7zQ99aie28/UUFDkYAJ8Q9mRvUDuaEYClCszrH0t97l1
biEi75YPgUyrtvuX8FPITzW3F2Lqd7GXyRHHxkcDd3nWS18PQQKR6prpE+bG
DWmxAWtvtA7jOMxAOzYvwVIRTRf60ol7KQLo1wyk672KSwq6ycAIjwmwtuGK
R3NWF2sRWUrJ2+bIyhnlmxwikDeBNW+//yJVguEDF60krybuS2ajNrsla+xG
/0pm4POCiy5JdHK4eQftStKEErXLm9YkMymiaWoJdNgQib3e/5TZ4Nr7qSxM
9kQF+h3NWyYbW/KZFwa1MGy+8CpBMUhs2/UgwmeeqaVMURtgiV2h7tIRbZpC
diRihQG9KBVcIC0mbVewGVq3nnSxHfmRrcQrGeKkHyT3jU4Ysun/tPUdEt+Y
ZVjM7D3zPDIUqkJ7DSLEM4caaFjskE6uXViobLqYR4ksGuwZ4AWRSmuG0XtU
/adaAOhDBNbzAEoy30LFWsJsCMRdbmeX/hCHpNloirRrhpudxpYPt93HY6Hs
A9QunertRmrGCswwZmKTMMZ6s6wUdAbtF7kbRpIvq58899WKntBXGZ1XYqcY
2d8JoWpSMzoNlPEr8JOQZMRe45xfHU+kh29cQCcVvGklNmJJzxtPyRS+OVYO
wPn50uG661ybrXjRsKEdr2tWzsvBLbFwoahCvFbdxZugdmppLMuMdV1WRwWH
ah52WIwJj2fGlEdpZCgYL+VPp5mzzsAfz+5CjJ8i9Sq0nq7t4siM6R9VPmsf
8vN504kfE69OaFTUaLllUHkdwtUqQ2zoDYjGEvPr8CpfKSXBMd52HAip2gxW
KNTQhHZshPM2GE+5t4ppF8HdllJvx2BBlHhgoYnOZK1Jg/JlIosY3UCyMH+3
qMlOE1SlqscwNVTs+Z7+SGqwUXYWjdBB8gSDoMZqVznU4JUfWyRSzHv8YmFj
Z39Sr9sy3ZnaCCm6U86Fp+r5FREWuCVgKeWAYKKqzLKPtiKP+e+jlqhpNp8+
EgTkiB8guHSNnVwnJNMFtPkxOHHULMa9hvHAUw75rscu0gG2gisu5/R23tfH
m5FzgkvLo9f4KGi/Limcrjy00C5PZnys8mpIeah1ymycbC1cZxY7UMyc82Rh
9JygeKOEH2CIWukA2/Z7FlzXkfl3yGdSFffnkEl51/XaznldSYK3q1+fyNeF
BY2tV3pIh/IGewEgE2ixHT2yKZLWB+xPX6O8/YdU2472993op+LTCGVseYez
KANd3oJwhpeiTIE+xn6YbHdJd7FNkda3dAjFEKTyyYfIAUCro8LUHj93S8qa
gMcw+MlzwhU53BtJjcooPiloYDW3zdnld1G493bka9t7TZFEr3t6AB2R/u7/
SNHHcthHc0K3G/tv8EPHbbwLDMBg+s8vRU3WixF94v0L+XQRWG+vELK5UM1J
jC7TECmUol0E/tRDYIVYVrCJKa4wN7w88sj6133qG4fs6BImwgbBJqRizSu9
x47cbRzjJdV9y9FvtODwVPgU+GHuzWX8Jma7TxuqufNZBpDSBX3O6sfLVAim
qeK58ka1Vj39C0y7rgQl8Bp57knzHrfZf3dCIJIBqx+4vCqFugnNWkHxbhQ8
Woln1+BOUtOuYVuNPCMWsLiJ6CG/RTFFugS7OI39T16PsTf07BY05YuMGqy+
7H+nVoGFoyJ4pELKYeWOmw0HqNDN47EOilZIjIcNvBwaUXy/nrnwb+nv/JrN
i7x5CUIsjvdKpa1FdHmLhioyZuhDhnfvZjkm3REgXikCcXyBeLVoMu2Mc5xD
Y7oRAGb63bvHinxCJoIZIRELeVAu/cTz4U7EspC8z6v0R7xYR5GE0XVZdGmU
aIKr+baIp0c92L92ezpyuY6ZeSXm+utk0tdiN8cjgZo6yUb2n2UnYsD5f1V/
tLYVmvcXO12/Wv1DhNzUExSxjRekJFf/nSMmy1Xy8gCj5TYmV4JC6/cxkter
M0FLelH/eiF6cZk/CYSn79/T4X5qv6Dkac+I0phk67kFQbGEUHCSLqBMIRSO
tB613gGu68bmgD7IfKEj2vkRWulNFGB0T1pFXwJ+2N2ii4MR5Mz+6kmZj/mK
CXw4M4JJEpNBwe6dz7Uj6ZdNqvrORhsYhrvWDK/flAkRiGqpkklZ90K4e+O4
+GfwcQb25a5C3D0eQWLgxVQfSsJnrQudiE44RaVyOSmmkRoPBvyoxic6AA2p
4u7wflCv+h/S8or11mpigznjCZrZQag03vRy3EFpOgedLIjUP9jCe8B0VDlj
mH+nd4lWrmR8MQgL8dkDTjLY2xFVZc0oGU/ouyO8Zjh/5yq+HhPqaBSn/uBK
ijm0JMgJY1JY3DiLnJwugnGHmm3zTaBdCC1Sr6WnQkK1guTrlDwHYM8jGpdU
VBgEx6c9FNLHeUIvM4L48cMCSpbiub6AK4khfN4keYgHbpRYKiPPIlz7qSCb
jGkhB7ZTXlUFTJH99NgW349vsYQfQ2/Efp/GJIR1B5oEq40J54jRLEhHhhWZ
k2QtJ0tf9+Y00+adXVYcTUiG3SjjEQAWdoqTUv8S4WM3qAIiycXGqj+I+r8r
pImaikfrSgnnyqCN7oWiufCAcwcLJ6IVPOHCH5eNWmambGuqzDT1WhzWCymM
BeW4phGWC0YmU0S52BJ7RC+HZHU0hWD2VfuQO9XdA6Q9eFzAgijZhclsVA7J
4IrHgYmVzo5u0TTsmsdtj3hXqfL6ySgULv5cAjB8BSfwx2SRxqacVWEUi4V9
d4F8wD/VyID+CiAVEArXDywK7W4Zar4OGs1pBqlmDI8SaHjNzU49mZS/BXir
8inK3WxdU29bSE6DHRDJ/mXQ5sDsAGjetv/6n5Slhr0QmTVgqn47ojkIeaHg
nIXgvoAnQRjoX8p8lS/UbKyV7xQTG7jHtJTPYppcM2PqMHPht3UNmBtrGWSk
THeuK4tuKxpvtCDRH1l6Jvw+qMnZsCcLyTYdjEtFR9tw6Kf1geKeH2pxXwOa
gm28Fw9JcrWFwQfVzUTMinPkAonPzqDDBK3ivzTaBdFmHLa7jMKknRj3KCJV
YfMLOOISBc0U9xAr3habT9XVQ5zP2eLTP8ohBw+ehP/V4a9s2wGHa5QRawk7
V7XbLnlStDBjo4mIwTGCrvv+R6nlgjxAOuskH1b03ZuR163eA8nT9XefHZs8
XttYG4zXVDV6CL4OMWrXOr5+f+FeIPBnzGOsOKWRZi3rXKlKbTnRklM3ykp4
1tG28oJ3L5oDnIkXdIVl58C6BQ3cvDNyTdkV78sVozp6omzWrGH6V8ynviTJ
7yv1Y3a04kG1p7Zy1eQ0vjyTxFGyrTrxrN0Mgequwb/KbYiKh+W06I7YnDtg
TZ2Kni13N5y+dLhrPJV0cLympAyIlDS+vXhWy3NvltR305B97P4BC1txZm5a
OZneZARzVm8GNnf3CLLzHpXfo6grCM4pU2UjICgExyltG5ZY3AEUCAQtJSza
+mNjARZ/FYeACpu4U7dKx9dSeitQnf+gz0KPi69b6WwuSav2xj0A/iMEnSJP
3tVWkd+rIiEUyqYIJeLJrjUOk7tW4Q8U2Jsh2xBOiLKMvVLFocL75jYU/hhi
GX3bJg6zVdCqD3kzWnkliFBGcKnYVmI8jQS8WlV69tL9FeXEceseDnXfGqWa
G7WCU7Pkad/bvpd7FRTJACyKXLlhccEmB7urRf4RnJjNb3gU5YuHb+WW5ge8
QqV1BlW835uiQ75DIjEWFP57FDiYBGlYZIZpTKFQns+rwrDRezJA65y53ZVE
Db4Ih1JAW6Rss72evKmOgj04HurRif//kIvWHWyxUGKsj5jrM6ZlPxpEncjS
7nMqbSjCHX6LlZX9677jDBejRVckW0fuSDs/3OgJa4GydPVDMwFr4erpup1q
zlX9A12x0iqa08TOKHmbJeB6tAR6gnEqdCQoJW4OD/PUQ0/a1g5ot4Jnbmi4
L3SAALope9K2X2blNtyva6+0UtCvRpPa59Js5WnBC0xTDbz3TzQL+XidvXF5
VOs1yMctSYHR96z1K1qabYuYjlgbILJea3FgpAAHd4adyl70WLIuN/wklsmP
T9acSoIzv0snokAdfOnZMaRdq29aIU5RknwhCTTE3amV8SfMyXPYE28K8G1n
LAzevy7KB0z2Ncf/uaWfosmaVWgX22vrO6m9yt6/9sI97rtgJYtgTnOK16jv
7UR2S6eiAiyw9z/cuyee+5x39YXLpqJDFs2mZrZbCGjJtyT/u5ZYBM23fHkj
EWOYTsFB95GHnu59Rs1EwtLnI40+6kBceLZ6D1hrsi4bXLS/2zF9AZXENukq
7xUgxTmQCRwIaSfCkD9IVNexG3O5QUmzNdDKJTwhCVOEqozoc/CUf1m0jSmC
SfkkHi3SE2VlvMomDwnBaqRe3wDuWXcoz78l0VlM0/Ht/dWdeL5uNNhfUqS1
NaGJV7m9e84BwNcg8dHn+slDDuxq2hxopx1RQTsj6cuyqNj9rJKljrgQhqOo
hLbVZQsOV3zLXac5p9VPgk1/gS8R1u46fhrda4rLqwUz9/X+FiDbQuC1WoTo
2GJB66XeEmX0SRQI6gCNV+bzHS4g5eCilf8OplyF1ZcTnWpD5V8+3yQkD1qg
lZ4FltlT+ovOJysbCbMVTisuPUKo6WKSdU2y1oe/ClfopV40XY4MYIgxeba2
ZGeEyXYHCLRJKZgamEPY8yzRh03iTnJQh64XaJQXyrrHxBN05SU0Wsb73TKa
YzgS/3dQUflrh6oUSdKYfh9bDaQ5jRmIzvmYGu+AyV2r2gsR1MU0NQk/xGQ1
pgQvN3l1sEGm8tVnl8+/nAvZtd9WWYjK8g/C9KovpFtXotoKYbGYgkp/DsZ5
hYV4ufrpMcarbnr4Fkq7dTnXmWjqpHnnqilA5r/BJ0DHRB9PF4Z4Q2SEOzm/
xYhkfDG0OBUDcUAilyNr2SctgOZwohSlL2FThRAvuA0qN22yC7Ya9gFcTJwy
uLKVfUg5thVnKS6HRKiB2D95Z/8n7pMQkq/7EbFXMHQrzEvC9mvTPt6FSvW+
r17bcJWUdjGzHsreE3FXXMp1B5zorCsdxyJtEMkTsbsWpc3f3/uTQ03bjDsW
zVyIBV+ratzmlSE4EyvVNwFqnnx7+IpBOlvfxDCvTqeyFp/6diu117qU19JS
PdgPKU8yatWqq5gGGUPXN0vUfuCQjtzMHHBhfx6/UpfLjnJd68ENc9invERN
M52WAfZ3OzIWK0snUqY7lbmvXJMQMrOix342oDlaE43FBDYhVHsEyO+EBtyZ
m5qKuS1mEoowV9BkRjC8TlAeT5iBpydRPN8/cIjaOwxlZ2dDVQzukHPbUycd
NjAJxDVda9edbIFYbKIcwJiyvB+KjnJ6eZzTTGzIkqdLfZaHXt0mL3IkHJZt
QYDIIOM+lct0JavZI++zLHnS32lKw/7P1+cJ4GcWu6rd9r9SlNWxwAwsqjKL
dZBYHW+fGuRKeJGovSbJOQ4NiIDfjg5H9DjWuuI5lBL94bQPLIVOUpvJslUk
zGb+4tOrTQhVQSq7Uulhss6Gawc8b4k6q0DgP6WhqDzIPYs+FrKv1JQ9wCL9
esMh0Q3E8Q5ihrvX+Pp4INSJmZz+u5UusBXaREl5bLwbEOzdZcOPdC/gvOLD
cMVhp1nYzbCf09BWfyGg1S8b3F4smlKKX70emJGrFFHfmFaS/3ZdC5taildZ
A5lv5stgiUwrfIiYss+MAcyy0iGsrVVuiXNonl6V5QObvDAJgcMkoteyaHCk
+u9YoaRtRqRTtRbUXqAXoR/iEUyN8yw+1up0uiNJ+BaFMcm7wUnew/Jb5gQz
xE3DB9fUcmNJRMjdRW0NoqHb64R/PdLiCTiK+zksDV+iBNwQWBBwBAsbyAgB
DIUl11SnGr4e51OBipYQzrOyz8irinwXkn1dxNo2HlkFZCRfPI7rmW5I2dlM
rbiILuhyqVFU2+X8EXvWtUUXTihUsQiAYQcRt75m2YEpU/dSIxKmh0vvYyVB
lRzvTZXxXw0sbVfaHh3Dt7SaMBavgHW4OgAQ7NO1XDsL0MHNF5qvBWQMSAxj
SJzG/Vn602p75plThj9N9cIUlmhKIFL4Ap6qW0gjFXJ1SAqWg7wJLJrDdIZi
MouVc+XIOiwGVVSsE0TIkHfC9qY6ETZJr3vcP8K5hfjMwXp4b5pF6vKo7viX
2hopgRCa8YKRVF91A/5VdX9WbkEZOhxkLkueSzwZ0R8hUYV73C/cWPzszmlT
XHFTsXvOw/F+3UOnwuS3GMRddn78jg+3GqSlK2Vo78WVni2KvxTaSkJw9vIx
+ZZWH0LbESf8khsgbZSFifME9m4hDAKSn6+SuBM9dlExCLNTSNklfCS22O5S
s0l3NbDSKsMy18Esd3L6GYHJyT2/LNMWlTf0I5PYZJrPnZdq38wjuZifcGuL
PuuVU1D+ylxgALsJUhaamlpcn6qDcz+JtOwhjCK6/z9ZF5gj3mguo0J+syp+
cJI0rK3Y/wTbqAWCqLtpnSYpQJvy8/yYgPBy6PbDQQ+okTDxOBN1yl1EX+0U
sK5txoYi0eo5lMamliuKP9a8zgB/02veZdtfwG1zWLKVScg93YoRIL/mQuB8
btZVY5tRp/xL8ly0hzfCCSHHU4zUnlkd28nJl48O0mQAZ6VL/Pu875CD797z
+uZnN0hl1fBCOzt0sYws1yGPkGnMA50v9sBhllyuuz4xnrKcjeUMYuBHz5EO
E8WvswDxSbZFFQHzRDOPcVDDL4Sg+exKAXZy3vG6/+qO0h8PPBhBXvp+0a0k
3yuMdLQssmd9FCGQvt4l4hjdcATX2opQHhz0U7RZcmJ4vajtZq9954t4a96j
2siz39xk7YN1AxB1sx57QElMcn9oG8GuTSPuoQHhlD7ly5vphBRaN5d/ZOyB
W21XZi4PIdQXCTd03B7NGzc/IySH0cUspbLYH9nS1YsPcOLexPnUAaL1hRrQ
ussnVH0BSkJci2NMVpXg8yYrW6LZdzMSqUlAxeWEyixV3mGyuVwzAi7oTW8n
jAFtorN05KGjE8H6Ttq2hPRdmDDXBTmK0XQbNcB5cnOyzZLmnywgO2xTDhTp
DSFZiDd9hswDfs25rT/xb2JFj5OPr6CSmIxRVrgMeozGYOOmbRJ/D86wt/mx
Fh56m6t8e94xoPRarSQCGJ6/cc17H2h/MzszOMWM0QNVGOHTiUOaqaYTsjk7
IajNAta8EJNWSJi01k6DaRjwyLHrGb6Ke6du3E/vXWEQMalUejAWx87EFmFy
KJ9Zho2CZAYot/shc1hORBpP/nAthuQFwHVGJrw9qg9nW1kx17yrbuKwXfoH
C3LgS/XCAdzEhfpeMt3IAqkjQwG+98Wj6BQ4C1GkHO45uFDa/bBa6n80+Ny+
rnYSNAuveMe1W+O3vVgLjSqPKh4504EKQOSAljtqKAQbF+r7g4gvYtQu8m0q
A8oPOjBfGNqlS2Kr8026vz6jG0vJXMdHVaHNHd5kw8UV2Cm0c/2Wh0U2rJ80
QQuvGMdhlQdGU3tzFdJYPAu9DnNSkYKfTMvi9PT1+s8vViSUa59HMl3okvwQ
R005U5u1DPrgFf4Jy9TGOKZWFALmj8mhsepvNNULhekelrdhhla7yr3mDiLo
fDTHlyvCdgOMEYN8GYujWXebg2xEO3invRY4HIHqbmos310IxOp+qnfJiXhn
eZZc73FbRffnztGgd2dSFIQp4+vDewsNU+XrH7WcAzxQztD6ghXAH6NiUICe
JOCk3mxm5AjbkMXc13dV2woY19wmQa7/ff4TFm/A7gKaQWLeqjEkxkvvO7z5
Rps/0KEH5OV1U2fIkaFZ+jn9++nno2RE4N8WskRtfHGnhhGvfpa1MGTjvxQf
td6TODrJqVkrKcwM6/08xysEULjsUsw5cwsRhOX7c9QcAb92uiEgKVBWa89l
LM+YNzHxImS9xMG2YPeVO5dM1ndh9IKx+/WxxSRpbNEHaTjmMcBmB2snq32a
0veFRLx4k+DmfdgORJ8dt5knk6l99E3lSTCvwRM1aS8BuzV54BSkdj9TYhZ2
tN17Vyy4WQ1Lc7OuXRE16tFQsksE0pCAjgMrjYTUuiAkAekP+fdkrXpQpjz7
VuUNsAkz9R/+m6hX22jLLbQKsi/D5D15IxFAyGfOuSe9yZBAyQAeNuSQ9mxb
k+Nwyh4zV1894oiqi0cbGUM1fHp6+4os4M9AKuHcLc2qJewQWP5/SY8fejgl
oSwNcJ0YgU6rWF5lLwXffmX4KeD+TQ9gnMENa2mqSbwJainE7iolkW4Kj9gJ
fxR/nmcqyj/1ebakpY7EB3ndws//CKfMMhFFWSjkNIJd2/mM/J8LGc3HzDSp
iYyijdKkRWoh2zHkv/wbv9Lv3bE+of28QUOIJv5gNpbKDhClrV/Gc178nmvr
Ac2XaBjj4NKvAFZFn5SYZfVhTxmOtepYAU6nuaG6qyXIEDxjq6IpJcG6hYQB
Z+oT8cU7omfDWSc/C6OSddVEul2givXdWfmEY7FZO3xxEU+U/080H2KUkwwD
rkt7mYKlH/r7B+OeEY1twAh7+vPG0X2A3epKIP5s/94h1FmQz/Vd/RDWK/py
FM5yHoGR7/WRaEwkPC98CHAMqrPApAL8+jr+nQc9zgGlB6PZpAnC0h7ClvRC
/Wa7E4KZ2RObHHBh/Jm2jvX+p6FQ2P+ro1E+hOhg7vydj0m56cTO3DiwdufK
xHn//xSP4j5RwzAzFvc4Kvk8PGbAn+uppjt4XWv0WUMJz5eCRH/b7Jl3vqO3
H43RyXnKsbRpKzogfLeiWokNHprdSu8Bc0iqvAAfIWPZi+8jYK6p9C+inH0F
q27n0D2JIITJDPuT5K8TlbQdaodMJEu8Il/Zqqj4So5v2bWSDxS6/1Vd/aWL
VCFJ8W8tHBopRAhFybRBGmjbvpE429V994I4aIaT5veGcIpOmYPVUKRl6wiz
rNYQSVmE7YZvM/sPX7P+nasd1lyHUJvfGgRe8RcYY/De/OOZG1/rp3k74oiR
57rK07xt50hYGg8zglXzUDbZxLGYfpJ5dXFpF4I5a9wq2dCyZf9cqZEqQl6u
gHEt4O5UYrNB0slau3ARsw3zZMyvWUV36p9LNrqoKHSzRf07m6/b968g1D+L
zuyJOhg2LvaAdHYHokrF/addVTHShvVao2potkB44mCANSiiGd+KxV+Vn1+K
9MWaJIs8aqMkQe5KEFVgrQ8tGnCjR8Vagr2U80PiKlJbyoHXTzHt9oZfRVMb
mxXp0YKUGxbmUuzjtKYTUTRhN5yZUREoauF04jkSID+GRkNf+0BZOPa7aHCc
5WCsSoscPmQLpc/hDZfdMLjfkdCkJfcEr3KjaGpRurgNMCY/4Kkm7kCRvaFR
0QO9JJzYcGSd7wL2TBV0Ariou905oHHvhjLci6QYEP7wPfXzvBEqOfDrNUaf
q3wsV/EJfkSsX/BbDKLY1ha5kWMA1xzD27Z0WxAO6kwEVHFvoApbYXhcS8W0
xWDQH/6WPrP8YpeRp/dPddyO4iYNdl4AMd2AzOQLHDvulZTg7FS8sWzmIbcY
mER8XomOziY48VxukT0U+rwuRr0kAD69dLCQ+WjNqnPsf3niAMdbl2nIPbKi
Zo3CIHEt5yKS/o5o/Iqk79K1PEBDwjLIIXqYNugWeEoHclGtVWJYg0pbb8zZ
W7LlxE5XISUPaCEmfw5tAWQUSre4/A8Fs/lET0HIyurHW7ItyFHTDXZ5IrKE
OeTloD5v1Dx4Bk+diRkUMblMli3+z5DZazXTptxtSOOm5BS8/yGkTEn/2CVU
rHYIbhIZLK5dC6uWiofDGyGkTqsKqfLu7UESTXfuj7LJiohBkNDulMqVszDX
LF6sB9FkmzJtAAFuoUASz8B6t7wZpOzMy/VVsDRuUjL0yJ4Qy1iX0jlT148F
4z6bNZ5K8h4RzM6IlMSduBd4iNMvE7nY7cr7aJTRz29Y5zeKh9hN/uEG4j61
SnC6c+imDrsGN3aHGXrquyVd2Qhjes5ZczRRw2mqexc9MXNDai22aQoPcuMr
nV2+zCYrfoe7x8PNg9at5v8cZpvATeH+rpdLqiXoaRo73XPaoQ0S/dfMbApw
jsYBgqeeQZq9Mg5anddnuZzb6jIgZVpPRlEj//KKM3yqfWqEv+TVjGzr3d2U
0vxSPqtbrMs/adaJVUBgCyOe0v3fPfG5hWujI9EDPmiWJY4cpX2Ma5Tt8M20
nmmGPKaGgmYa+eGwRLskj38fOxLJv6uqP+E94jF/lFlMMkpAubjNbyZMCC9n
fPEdl0x2KMXs+R1xoA4XrzKTAgcIxc5nGHElyuIn2eLaEYu3dYnI19T90viX
ZWUhtHLMx2XCA8tTgoD1z/I/XmA3zpvGk1eb9Esn0tN7yhQ/V/LKfgWR46wu
w/hpdo576bbFk9eSFJTl3hqm6GLO6OTYCGIKrallIc1x9FGOGR7Phu3Awp2E
nZb1qLDcTcBYuJAL6/7AVjp7YA2NaShzv72MXL+w1a1mBx9dsRwuohVpSFaW
aaCdtxZuFgHPTvNzUcDvuJtb6RzUE1xekPghEoMTiFpChLkA4UWJDFJt1/QL
O0Gj/cZbZwHdtbfJHsD14kn6pYSLlAoJkZOAgqZVZlswD1fT/cYaZqXiJYa4
JK7aLUMu8rIMK3UzTMTle4ZVGfoTD9J5sokpMWbPQA0cqw6GbbpbDmmymnbo
3/mbp0PtLqRzWu342n1jwuXB1wselja3WuL5jD0mKqB2KCpVvdSJ4es8CmJX
gZY844cW2/Gq0M/ZZU1q9TBMGhEZaug6eDkCh0vkPf/tChe/xPbSgXVVMa4B
zKBPfaGXCxErce9/QY5WKr4sBPO9cEw/pYz4zInT6xw7w7oOD0YxKsDmMhYi
EXWAfKzir63847kpdRX4VU4LfCZb1e9SXjQhKecG0DVZQLafQgTC9r7iZ87s
1TWz4GGigUGLLZ6BRB5qhREhDkQ/VcAGjzpSwYiycLoEiicXTaFuU8pyTiSB
wfvDnlQDDCWcNQGX+pu1d+hvy/ZaIxnR/IhoNGZzNaKE0LOm8jQ3jcbxDC7B
ZnaZamykfCYsgbxV866jiAW8I28AmQfkaeTiac0l+WBqC0hg854C6F8I43dL
NAOnHUi5kABtWaLhTcu2dJd8LbihilqFChKTMWx8mcooGP/FcivkRM8YsW9z
u5RXmw4KYoj6CzfvGD1YeMIIGjyfcQU/vBxOno1dbsknnicVbh+b77LZhhw9
Ui8bVdwl3jhlhGAnL96adOGRCBqEcu1sNkBFCBezodPOIH+TG86RWQoKEdjc
ivM6ugJHklYVNmLxu/llaUmaSJgnResQCZeUA5Z9qFAE7iRsLGuZDN0d6BJa
+z90Uc64d0toYera4HHZuyy3ey/jId1gOzH0JYjh8aVBQJayrWwqCe7JMiyj
EuXpxWZvkB6S6XquERXoJdYXa1PnMO4kOtAoqCKBOLezmPr1UE7zDORIvPO0
tRbASNFcYCac/Apq+f2orxOqwzNNLh5iiVIRfz9Bw/NOo6NNM/F766KOOzNA
pr8urWERz1Mmp7cqKeu1BzNJXTlIEYiKHtRdydO4aWIG4Njw+f+UQ87oRHWX
ly0S3MYZTA0w6axqrSInbLzW65fShPjD/0mUSy05uD/+AKhtG+Ucl0Zuo3ds
8uQrrMMju/3NH1FKB2dtmHDRKMw7bP60Q5EnHKD6UUYe/XMHuTSQX5rDC9cx
XeBYdAVfkPL0sKME8CkYCGpKOQjKPyZ+FngF2eDIUYtGDRahG7R7LdrQxYPR
kwktqFb2Ugxl1UwU1vaR2VO2vTNVqXa0AjgPkajIEho9a4WE4iM5XLdSysyW
pIjWNCIBIu7b11F/2A0u3drCSz25lSCC4KxQ5s3QMQExHPlI4xcJqEzhL1iW
5vC3yadHJrLRdFF4x7ZFM8V+3EeF+eXZAEtjgHuhud16/bpifop0OuDvDJX1
pZ8LCJENr08BsfwGzMq9eoIKvc8HmI7p0jFrW8+58yFSOp8Gu5fvNrl9GrOj
3IMYtY8vIEYoYOeQRUzL3/Majfn1fEH3CLjm49+Hf/W2Kf5BXEM+/CvNuX/x
1hxIzlk6jehg0SGJqZ5Bmh1eOBVwaBdBL5vSqGQ36HHDDsRmT8Yf5W/byU9I
v3575FLjz6gYRn0UtNLA4EG2wywIR1wKWXTBTNBw/0K5wNER/IW2QY1VNozs
8/ZYJR/uvnk+PO3T6C2G9oAek9sA5YlS7K7FhiQyG86oq0vp6GUdrxrPX1aB
4D0DSLMQEoiHGF7fqADDp4+9y+Zwt6ZAAbKBGfRMdyIokX5w0HiDF6g+oHBs
BlOftKuTa9CyALMaUPu8Mk+5drcHF+1iD1x2qN84bPPp2IKXBzdm6aRYVmSV
N+/8TWuvkb/U3e34MMRbT5Y6jNtDboUePARhLE1pk3MDWzuZFlTjoCLP4LIl
8wh4Ci4CCWcOjaZBOILWpZdYXAJOEKaWEiY/VLydPurJ5TD34GXyg9acoKPu
hFFbcAFYWQBECERDsPfChL5re99zfN6es59sjLALFPX5RDCEEow8F2klmzf8
5qAHeg4MrBHzHc9lDXr+0MKkuaG+GtEHm7Ad6ES2bpCVNqFK8lQ0DPAQmNA5
UJecycpCwqgrNU+wnvFtnMg/Qub64A9Ll9yozPM1vS0VqvghUWUssRW7V2r2
Gv100PseMT5x1RET0gzJphi6n50OuJzJ9QBPiRb0zubmNiKPTxR6Kt3lpaG9
8ucSbfhTdxcQ7KmXxVy57lvmhuzwH+f5RFovRaznEgSem/lt2TtC4pQaYmsP
d9GzyEN44hp8+D6GcuSEqsxlk6be9/5kSB2FoqmPyd/TZPHFhloA8xrCYHgy
vH8AD1g3Xw/IWzv/Geu8FL2/z86r2cx2CU5TknXNb+lVS4QuI9NZXQujujwp
wJlFt1UPzD8tZxaG9STLdQKfrhHXrxu43t+o05RVjv2JLhCt6hSxqisTi2Y2
VOKOFyKa0anSDTGhWuQhcWxmMf3rURb4FlMKeB3Nva53FmgqHVRJKNMlYgLe
h1Umv8w6+kaEzh0fawnWEzkmOG0RJBbx66CqZRejzyT/J6S46iC49cqKT3c5
v1WxH8FIWjaXnx3Gj0pxMaTyfc77dChDs4lLsfC3LFUV3g1EBFs5p8/h88EB
m1/C4arZCL8zPiJk1+BmRcdP5BKVX+2UtSEijqtr/0P8hnLuIoeHT7f+fcVE
HsMNxw+w4DYY3Syg1Jqb2lrjtFzsEk6ZKm0cPTCkoDHJHrpcoORJjC2dMC83
wuAtC60ndwNs2k/AjYUa4yhl9y+rvJ5HwveVZAg6vrUW2ssvFx2jKFGSFsqF
5fdcbn7555gRJHWE/C2Y9Gd5a/Qta0TEim8IHvta92GjhnvdNba/CbK0X6NI
L9FoHkqCDQmjShWIlDthPJApk0EgOck5bZFdoODoGYM4CxTerO169JQ8zwXk
V1pWCT/xt9oenYFQrcicTtGMXC/SG0ZyhNiSTkZab0W7qVAXHKtltSQQwkuD
hFyfShQpyW7hOIJ8fp556GlFeR/obXXSUyFzLD5023VQZcgtyplEQLX+rvQb
50EWi5B98UOyP3SU8b6rSWNg4JS1UZQ5ElPElo6WGic8ls/Wa/rATbXRYS0J
FFQbnU4wF1sIl7ZIBBKauVS7d+eMG1DQ68fVZ1eeetAQ6dlJc9OHL+etq/84
81ZWjd2eJgVTj7ThtlgG1klK4eDf0d9T71INb4S+AtoMmXgivo3UuxB4XAEh
qftz+VfrihOjWFR+hBSxAIuzd8SWHVoEHyawTgI00lYMYsbfSUvfovDV0WKA
f3LoyaI6znBJR9zA/Th8sRJIfxGoa7U12qnBdb7DVeK9ipi8QBwQz8V1nPA9
UgqBL+glrKboHGmOiZcjLPcHFoyEXaxUsoStAtNCospNT9o1/WkpAk3AzB4r
vGXI4kuQU60ZVwCUBJ27pPFoECMhlcY9yZpkn6zONhUTdO7N+Krfc5qgCIYp
iAQetHv3HcYrxmQ7629OGZzSoPduQPgHL3P4mLF62XZteYhNxvDEumzFxTYq
oBaHoGfyoe45RlAVCFqa1O2vg5YjoS4IwlyXguCEBgdBFVuJPEAtrb1lcXLe
P6IQcSyeq75P0CXubGHPiUJl1KPabi1XSUeFTvqm7pPa0AlIrA1zpN5uJGzY
gDcLseJFKCJMdwQPh107Q9cZ0F3YN3rGLXrOMmUhEs7Te+IdiR+wwTVBGv+x
eLLFFU5gEoatqjJ1QZ8f03alyleCK7ZF1MmMYcQzfRqF26GHdnJfdtZx7cMZ
VnaVcCqLAzjo4ZCuCV+2Lkys+dsZBztsOfhiYWxHvVWvjRZk0IzzXma8UPw2
sirQBFNDb79BjeXR7EUgJdZd7joeOAUzsWWfLCutH6XBeP9xVT62JbrUtTLX
yQqeRHwEnsN8thSPES539mki7ky3lCkXvE6LhtEoKuLNAvDlM93GpJdnsrSz
AYzKlCJ9lH5L291cAzGBmAUuJ6/ua27xSigFR0FpHnmQ2ZLGvH0LP1RzrFMO
bsC0I29diSbn47EMLM+4M6Kz12eG8y9toC00boREkQHTVFb2xmMROAci29Pv
JoTJy3BSTAh2jl8tn5adQ4qjiQH/UKZhAhJ6q25Wb7tZdowO+LU4iNGScaqg
KCmW8fgRVWnMsmVBpMze3X4+tjj+dPkQbD9hh7kXznGf+6pKHMpBdhJN+Yjw
GYfBxIRz3Oa5R4pvhFmVjpVisHjI2RjlUy9DGGeJ/3prff1vL8bxjpD0ZtS8
ks8SM1WEdsO6Pt0Fh84BQ/FpSws0eLS65U19+oeFyITb+I6i2jT7QSdenvSs
PHd0TqQgW31+jJvzdNo97lKt6/vel5117cr4enwZpHiVJKMiwJhf+4+Wgjt5
JisOynjGTegUM0YPLcL6Vj3nyQuGcstfCq+MbVK4v1VL8qPGqdZRvta3KEXp
iMGPKf/4HdYsUCLkoNf2sXV2SEPxJM0c9hEO3QLhGbOQoUnwHb7qvaMtxemn
Ml6FOx/DEwwuoIJ880Lz180WZwmePlJNVlmet2mgMRM2wk6Z00vC+azc+8qa
4fE5UT2aw4VBoQlfPCkMQI/i9fKoBbI0PEu6BX2RcZRA4brDtX9G5Po8geXA
g/vRvAqkNUys3RdQXzmqd2MBCeupoalbO5h52pNvqcC2XkG4ka41uxC2Rfhp
yaZR6GmwVBHBsS3SYL6Z2nJQWuTx3IFas1M0MRonAFb2AV2XhJTHOeWKhp2k
oK36DQGWbTzCKsX6PIFXA+6HNAg4iE+EbyXmPIB8PRuTRoBiFO6O6DlBb19b
WhbmK0ft4vlHHyStSrAKvfBocMPkvkic6GPiHMg+ZsdQYW2eYACz2tynRrs0
QcUjUK/7G+iJeZFdi0VSzdicRh8cxMBY55j7XxECydiw1D6ZfVUvO8M/3vY3
046j2vssh0ISAljo5wnTWlqlJIXSby0IjURO4AAIDBaMWZTceNaeRThEBfGI
EPHZmUmDodaOxzkKf9BP6LLxzSsw2c9b4Gca/l/2GHlb1UyOeN/NNwWzumF7
CYP+3bBUg2nHqIyOpP26FJEHRys8sgfW6duGzZJa/vME8Nr7hFn0GfATUoNL
WEe81Va0+eEzl+GFsX4pDulD8HcJdSTkiaPumK5dSmddBFsMHcWRRnEvPqJZ
zMoN9d08pEIcajFlp4UbEhgrrgh2ssqfuZKQ/unyuwMdcDrCPmrBOZyQtK1z
9SzjxPxnis/FqB7dXooUq8pdfWD5uy6RCVPQa6REOBIlLx9auXyHaTwDzJI+
iu7HoL98bMKRBty0NZQ/rHKFbCSmO6r1Xy8h2hsUSX0aLeowU9b3YY29iLRf
/K0roohq5lGkMkAE1odpc68ufOT+AivycNsJRqQ0+8cMF+tp2ZHc7LR9/FdO
sOqr9jITWZoMdBJBjcAwztIMh74xDP39RCV3DQSqF2J0yCphT3aKdRkMDltm
ANUSTc3xh1bIHz10iEvLznd6KfAmtJtWNhkB1ZNcXzqzl7xfP2GA4tBQfHl/
yGHuo01NqXNw614+4YbMsgDYDAyzrqlxD0hRYB7k5e8oX+blUK9E5/Vt5/ay
njzSe+hbU0zChMUEQEruLMQSC1fHqKgpmh+0f6HkQlRHFWORE7NsyLEgyx3I
1x6nfNDWOIZwrXpXcSQrJ8aZp+lDG8A90z82TQfe0pWbRARsy4oD9WAQVKY1
E8T7+wePoqdaJdtfGD/OA3NmuE77WdW2WGE/KqNvgPoGCp/ZEFq4xlmjpxD4
WtQXAShN+D9SP0ifSo/U53RK8jjTH59du9GVWcN2+9/BfyuCs7A3e66l6JH6
9K0cnhErGdfKp4jHryfUrKVGSofgEskM5T5WwV9GD87wMcfvUK43dEH9K50R
AwdNiJgHtIEAzlQ30eydxIz8qywMwAnEc0aFu8b9I+8AZMsImWd54WBYhOcf
zEDD1mR3AcPm81qhC49K51B63hdFZ/LjFZ5d5znMNIbcYcTui4QW/iZ0HBbM
w9XAZCw0Cy28TFQfxvN/5SPqFaU/bzqgN8DujarR1/bBW1LvLsmwAByZm89+
YGpWpwXng5Ua3PJSPO7+ou44qA3IPXLxZ9FjgSX3XC3ZaoPXIa+wtL1s2pcP
8xYcewLrPB69dHB8949ouccCekCK6Ot+RPiL+KOwybmj0lHt7GilIQdPvf1k
9AqkzdeXO66BjWjAYi8AUAh+bRbMqFxnOWS0h93wzJwNCY2GPd5aPY7XiGaF
MTbbTbAhFqe0TeRE7bBzLJ2C1QIUBYHWoTzjb5Bt4+UMZvYon4IyDzONMHh6
C2ei3Jxng0y//Fzraru4a2f0O1IkkY3KRXFtzKToKkJMAVPoWPTA/lc7qEQK
jEhxUFsijzg7/sPoDkXc3ncHup2uVjzOOvC4BX8LXSSW2gHE6YM7bUB3VYUq
v+jMxh7tOOJa1HFVXOLrK94j4Ut1pkehnBdXAPqedyVbR0/TZSdsQm0Mdptq
iZkc5kzCJS/tZYJ/fbPrRHD7cg1uVzCMJKlBx0572JKhS+uACryCZQ2cCyh+
1+efIEZ9c7K6xq4SBKCZDTbMSIHnMzGkfzUtjnsMK4+ndovif2NKhT3JFZRB
21zCrXhEBNUzs+jIBKP1aE5uXlcTs28NdiVIkiBf3z8vEXwyMdEvfO/RYCWV
j4WoiMPUOlbk7MKlGX82n6R2AQMC4z00kg0MN96nWQUkdk48pFHAqKSokq8L
w1+AwlpCiD1+yfzWiRr57fSsMU10O4k2e/DmtDfh9TwVD+Vl/dgAvlRopHMw
CZQXVqvEFKiF+b/JaTezs0WunBs4JnTfYhww4N/YlLfNhT5oAONTrdjiKKi4
aMw/sHwuK7Seb/oYn7sTmQ3tUqFEO69xi5/YlzQn5FfFAP+5R25QeLLP9irQ
d8q+f/IfHn8jmt5+97wZSOKxsmrKd+wfVvsxyElI/IQk7EUssXH3pa92aXL1
vRwWaN76WTp5iRrHQP3pGyPBpOpXS+8sk8H9cc5YnMF9xGZoTSIX2JDBTOTV
9vQ2tEZ3agrdTnXlLQGtjutHvjh9sbDST8gogr+BemyI6oA4n9FEj/28vomh
ALZ+9m1LkV7BGTYvlyCZsxww8EsytG3k3WU8pmSQgaMQkpGCQdlsCAvisoop
gBtQKBxhLG3ghlcbqyaN4J0lfACxxzI2IAwvp9RQNILzXhRc03vn9YMjD6sm
gxB+mz0i8e9W7CpPdi+spAMfAxve040Ohsv4hhKIJ9tIWasl8/OZg2/CM5sl
Z22jQNsc0oZSO8qTEHdc0eDQLIEuF0wODpplN1HJf3FxuMkfb2fepjIiG43a
aF0YfkvX65gjOt1JeIaU5cN6duxwU0N3gVi+lK+rwh3mYIjycuvgFemOA2C4
Fhu9HERa3DR4mqZQ/GcZf1XE1qVZzmtcomruR0xjFcbSt3iHq538w6cTYMny
J01UMM5ZNzHJnwZIYc5AZwb97Ryn7Y0H68XOHrpKXmvbJzJDN3APdQPu1nZ4
rInKhLcSmj9D4VtM9/O4SzpxMM3gfJ4Gn/1GH5MjFs3PUurWw/+0lnUiygn/
vSUkwCbvjscJux4YzvBUuip3LPQ5GGxupq0YDlTQ7DcMurO0qDPQe3hx98AG
CfRCkZxlL/Zelojch3YS3N2QgD7drglcUwQqHNh63vU7Q22GysUuGkqwjaWd
jiUiocA/C/1KK9Tx14pm6Q4PzwAs48jW88IYQgot0pcBMFdfjSpT3/mVIFWv
IVTjfcvIzxQOLueIGXWR6NIAyKb8eFtRllWHDbQ24nfPPvACQyiPu4NmCMAO
8pn+UEgQBPzkEULqYb+DK2kJ0LoWSG8c8xt5RxYeJV2DFHqxKsEMOqwgWfFU
n7ercet+kYJFvpqt+vWnQCSDHcsYwKtpPkonk/NEh67C/hjWHTH7Jb2qUyw1
2ZX/R6Y337EaysGEH/nhPOYAsobCMwySns8yO4op+FJdjShD6T5LlVjy88KQ
f/5CJiws1C63M5L0bm1ceJBc9XWOcm0De9/Qamm1kNw9TAEjkCFZZD4to9dn
Q+SAo+tc7CmquHoYCtaEHuq6MzucoJejjvErhrBSTjxscFSZQC9i9WvnfS54
rE0HytRaXhabnnDKgv2dYplNQmWfhikn1zCmakcc/ni3XcMKGj46VTMkj9WZ
oB0U/sy46EioSMw+RetEr0OlQv3ve66l1lRc78L15DnY2KgAoWGmg9ZFpYIl
zPMr+uYqX24lynKpQ8Wo3pxas9BFv5ObTaojUQbsDODEyamylP0ggNIsO9WK
o1fpHFTrUFdLT/nYQWreuVWbiSPvlyYv4QLE9asBzuXY69lY+bJ88EMJrbhq
3ANiLzb/QT8/DoHOX/GxUUnasTk2sR4eq+eeOZzv/cfUTQL3auiV1E4Ga8G/
1SW5M7Jbu642/VSpDHmO5UNjEDnGZG/jrgq9+8tUDjmtS7z5IBJHE9W39JQc
F3OE9oBbZ6urWPB8gQyVJmkEAoEHX0QjY9lWQ17D+HYf0Pl4VZX5IjeukpW5
HaLFoD15jzz2NJAW0N/hjrdRPmNwD66SvpqSAdKH5i9VMwKxIq+Gvb5HhpD7
QsFc+DM2GZaty2g0k7fuXHJhEIh0nwGNrs61vABcEqIYftNSQwEMEv0roiRO
ej3j9UtvXvNdN74Ff8gdUJcubINkeiuYnYbbFtvdTlINVPKxwN+HxX/zHgYe
afmD4cIbxe+cdiqQ0lLmcdjOJuHjK4C+xguG0gDyxzRM+yIJARhoYYbnS0Ir
iUclekSpyMnuF47hMrnBlnfbAjEuwTfFCHtqzdSW9mVkTaAb55HHlY5teNxX
eFEfJ7bDbHX9+NgCRJ0LynlQIWENJIumwMj6S47/xDar+kGx8dfSNoTQMG4v
meQLIpapRNQ3TODgZnFkppLQNk2yGZvReMwl5tVw8UQIJC1f5MF103a5RFrq
mAj09V9u/g2bGOxQuls4VK2LKZpmP7sgMZRBafab+kB6D8Haf7bHGyl47uE2
VUQS6KEy7UNvjuYCot2jO0+WNv3PtA9jLZybUi7eQH5s3tJWBnuxlhT/1O1+
RDGooar9IOicxNo3kOd2ZWPOyLEtXRYCv66ZuLVXTbYGPuYSMq0yEoLtksc3
AC2tMjKSAMyNapc+827My4kFTeMDvIW/VHrT1kpW0+AR730XK21AN5eyqbw7
ZX+pf1YKsNXQrV0Y0rUle/yIDLX75pAQM16uUNJbfEvsA1hPCfKci9Py+Ecr
OzwY3UAY55P/WRKsfdujqN64Ma3QP+9BHwfkUFz28KysJpHJl3aUoU2k00hA
k8xRTBc9aWpWDqQmrJMt/YaHPC4if+nyEAGDZDMRnIJ9YaCzwaLlO6dYEAht
a8qm3Er4gEEeYVg56CTJaOjTFVQd/S9kN5DKqc3GDL+TrD9j8tjesA4/JWxT
8me0M4znE9SPt9w0ErOR0/v69tjjyHHA5nQe4qRmrMsuk7CpDbZcp5nMx2py
WDfxErPfP7Qa4QyHKGQt00j5GWIut3ZjwIbiMMG3mKuCfbYGZVzHNoJP1Ihz
+Y80ANNZq0bGUNjuJylZzE8ekG6BoUaaV0DF32I0YPIyeCF4I2VwQW9hi7wi
hy0u/Co/6c3pL26gYHqDGbNQTaZARMsD6L8Y+75CWEiUc6PhWj8Q2RnhnJRl
k5gUGybn2gpqjEzW4ZqKeNw3LmiD3daAwXCOPh8M/Lx6hdh9t+FkpwgCi6+w
qojMLANSWYkb9+su+COOzZiX+yzuyeFQMZv79kPS163FF2HuYI6mdoBMcI0n
muveNnPA55ybUYed2kw6RG4t+Y/hPqnvCEvDkex2WvRIO+w6O4VTPFwC1D0a
IfKpbrDO2TB2KmJd+/dkYo+D5aMNOWucxjdj6v1+Bl3zH/DrowxdBla6VYbI
k6AC2XhTCzn29j6YVZQJE9LNoqXzZO+1+99XCrdmGgJ8+UaAxAy95ez4+Z6B
4GddiR1xMt20vmHHGGeGoJOPmaIJYvgUPU3I7IFe4AhqqkzwA0ptH5zpwJ7g
Pc/VGuPFrAUVtTjKxKQYm2fEvl+3mUR5h9v6VL9dF184k9Lew+0Uwkc038FC
VONLBozUX9l3V/ErnKH4fKd4KG4BoBtdCj8NEM+FsZ/5IHtZDelaID9gSTH7
ap3m5RpDz946pzca6wzUZ9TsNHKWP8udw1/w8D3xSR4M4tnykVBClzZPiCPO
V14tA0I8jYYkiSIJqA4EmkgP2ioC6KqRvAbbeRlMkNFSPUZS46YsMGchy64a
e5HRBtv5pKgKPU/2RNic2Om3F/MXxFvfd8ohyiwL9UkcHRpz8je28j8guBGC
C/DtiA8VFNv77GI2oZCOfxZsUv08wumIlGWMbIyz7GLFOfjQzo2HWPWmI3f0
ODrKASu46uZUtYobJgSvByCdqUqz9TV3xHiEMRKFET22D17TbNeJrvzlmsdT
HKm9VL3UnGQi4B65P/wtH1uu4n2GCZLMPVsKrKKpKuVJ+7x23x78CwH/6uMn
2YAQPH9KLycZsCjtK2rOgXQkDk3KucjOjHyV26hcR3wJENdHzULBCFToG4lo
VWxE03fLPARhLOUMRZUAIH58BYQRIQ8NpOxN4kixz9TXzZkQv2EyqiS96+Xc
SkkdsSna0mvgnbp0MQFOVyn0AK+eS4upm7qibEuDk1wSIYFRQnf95jlYuzyn
dJ68eLqa4PknGU9kvm25aF2IXkpCnC9LEFtymLGWGTYS6JCbdIXoYk28B3ii
l0tKMMzsAdPUBCcpemmk81+hjve6PxzKvBxdkKzxbOltn5vvUaEHPLkK08D6
tSZTgesbl43a7x9YQnSA2gj9aCzOBaqd/MlGZHd2dt2XCFJ4Y9zSOB0JKSsX
cnbD0HJeRFUVMofbBaFRRnJ5Hjv/DlDYfZQsMEwaUVAd99eaW02GV8X17K9R
Wm26k9rgNSw8fmFtU8q3bQtuiTDZp/yuFUYkd+gxUsaLT2gnMusD7+pwR9pH
3Rtp6CxG1y1dbYGBRMRIbgGrWEK6D5m1LTMODHVnF5FsY88OSpmcZQ5tJ0b+
hKyU3xAs58Gnio53zjwEWaVbBt3D+wv9qjDaYnuNlkvUjXhspLYdd0sfrZs1
2J2S6+Jf8I3WNGc42Pj0S9mD5VF+gp0rSXF05x128bDw5zS7BsDg2BZHt6mO
iDEqXY/SIOeh3lKj2N+XpzXTqDfe14MIHaBVmWCgdDFUAH5+arK4jmheYY1d
y6BR6i8ZldcoNGJK8o+AVS76DMRWHPPgpZ+AmjKntx+hoMJUaC6lwFqNgilL
W04ICqyFGqTxin9wwtX/TwdQ7ObnoHQMxNnITUnFo8vty462H9EmPIFUVzqB
EcWuBTDSyVgmryIuCVg76MUjDVOM+wMtCjoaCevAHvgu87FoxoCTFD2rETY8
CqdnVhx3FQRXVfQTmrZoJ7Al3ODne+6QuP7R9BseF6a6iKi8ZtGQ/x2AFQaY
JvulebSDJqaUCUfJMWf/fu+BvIgCB927AuGyl0hNNkHobeFLhe99WX1bId2x
n9QYqSErYm4+TyxuK8qa/tbF4gljEPjMa1pNlhfNcyWFl+rKyXlez2FIuTBI
xTzuexOgR3I9Vr7sSLEwN97GewqVv4ybHNoIQeqnknepAT2OQqiFuv0P4qrs
dMGNn23v2a5SQuM/1Oo46us4m/m71Q4rm2RE54L90pvVLSdUgI9z3gqSco74
GTD7Jx0tA3CwihGaa+cqixv4sR4GkqhCGVEsYS6M7NexTJuLtmR70U2+6X3h
ZMKSIqjD9Z5nFMZIELKhRBbiWNKLsY96EKhGbxSF3gpPtusA6EoVa6foaOyx
MJrtyIgbZtWhUr8UsITWSxQpDFEkcKlHeymF6+7ncTWqgyaMEj1PI9QyQRJl
2rpPjX/fxrB83ASlqUiiUu18VfJiYLwnl6OTYFYOa3PF+MpS/Q6pm6hd8OxM
SkcwAVFDC2nZgRutO8UTl5XjiOQhqTDCgXRnde6u8jxfLOXkrjULK1zAD9Zw
dD/7kO6NDxotc34d0Y3aZ7AGq76oYRE9kcspkn070figlBZ3liX4ewx5mpbX
UdHiUlPiiX8bDprtIuXZsj4/Ris1CUu2N9t+h1sVF38QiCEw5ib2SEyQbSMg
iAQixdKb5JDS0e3A18k5K9KqI9DDnTeX1AJ4Ynoo9mooMVIxcE9gxC9J9mEq
TYf1HaiRo/xjo0FzY3UlNEhNnCURp4WcTMvMAeWQ55J2Igu0aTP1mbZx1qdY
6G1U0H2y2u7WGSTYF9YMhaKe1/XNbaeEMjWVcoKHlOXdnSvs5YDd5hT1D/Wk
cdqFidF9iBoNXqizuwCrdgnGGX0vWhcQT+dwrwBkJbeEPRD1CnPOikLbM2t8
15BN5WPA/SPV8omYeS2CJ7uDSyh7e+rmCFs16pbAgxw8cwRbF1/kecGwJrQB
s4z6DfgHVd/o+FDr8j9GkPztYjMlm99Z0KnNDuDqZjad3DOvJOimWQFqv3bU
b0CB1rfLrmwMN+LLeM78OUhsCQBCNOrbUQFW/0OgKj+c5SzFWzntaZ/aK2IF
7kjrO1VlIHsyqd8p8TShe8bWRsHI6Ty4y5Id9pd6gaadf72V6TUSe/HkXwp2
yNxGiIwthLt/8p7rNejMhuw5+5zTxyynSosqu/tpRe3WrMyf7SUR99OFm8rg
pFknGK/jK1BqpTrJvqqAhIbOijKh8Csl7MqhZJvzFGJzndUu+pXiQ/6p7vfn
aWnqjtJIeVMryB3SgM3gQ3/montngQtuKlh6CYVGHn+oIVpnp4DsNl6dgDHV
L+IGG/yODjf52TdNCVLi/T0WdqSE9h1qWc9HXfIQz3UdLXQsbFqLhmG65CXw
/bCxUnBBXRijPWrUJtOVeXFeJjTmWrDKZW+ui5kgwOPGdnXWPMN26oAi0CM8
8olD0xV4ylH3ElNZGPcgsJy0kn44EOqyQzbd7IS7P3Nodl/HJX7oh0ZD4fWt
pmFVZRE/CU3/20LnlJLzH+x8/mLpErNeyRd1LfjTGFKAFy/gngYBmgGmJafa
YkSYOOD/Bqotc6LC7hh70v/qR64VPPM78cGR4zn1PL5ZCp8R5fbowCkQi+fY
ZMhq+q7emo6gl/8GFyYhEZ3oGXkaP9cF4mW9UyFqvBQ48FBcxWTXH7EyOdoI
NP+ds8Vmx6qn50U0ttC4MoNCJvzCwTjgGpB8Osm4z/JzPwV+mvle6OK2FcOV
RxgoifS6TlJrKp3nj1qF+ZYlte2pk3BHDwJ1NrF5ENd8UnffA+FMxjy4t8tJ
IfkkrE2PE5EeKBNlQEk7lXvIqMhaUJFHD9hKzpSugfFKfFjgMSCO1mLtIQp8
xaUzvdaqwOs5TdS+rb9hhOCrkRqx10mQ7GHLLoXxg8gBi8Lww2i95Hyo9qP1
pEpKObVMymNc/tVeJVuAGRmXu0CJSJQgX5Mf/a1mvBhOV1pvY1Tc1GgGsQ1G
gDAzd0JyZHrV5T9gCn4Vvr0eh5ftkm61G1rx4PITwnLRWNme329dvvsSthAg
MXH8iw+qC2bHO1UVZNshuutly++EKYpUcb2o02AWSx+fGyb0lN+XAETwSV1Z
xDS2fNLOlC8w7A7Cz/JNaFveaIKFGYZXZIYbXAjoGBT5hszbX9MTVkKTSlWk
Oqpgz6dTXUQmRcaDZ7VCWnmXzbJwrtqc+Pex3oy3/QLZNfX8MGP7809qOwju
heYzvaTDV+JDd6xG6jaBCA3+fIhCywWjiDWPvMzM1LnpRdtW6821Xwz6A7ws
QnXPH1nO5CEuQRxMCBqZ4uZAH/RIaaKKu396iM2kOuSFoSb1rYZzUrzmk9h7
tQXEE0mtnRyRxJqCOcvEq4+l31wk7zXwIRQYWm2dr6Zy6G+zOLWYyo6WEQPL
RIvB344l1uVqN+RAxZGF46e5QSptdVJCDu+wDSuycIZt3iwfycF4yQzXvMg4
Sjo0WHmrrLRPFqDl7YVacwL8UPdOSJQ9Ove5r8dPX5E9xmrwqYBtmh4L6RBf
wGEzQLHdgm7Jf+C9Fp0vzdqNs+Plkk29N6MaZ2z8yJMdDOp/4O8zy6bWN/Q1
fwB2EHYQa9V6Fn0ElvNf+hijjW/WL3GNbPf4dm0kT6Q/8a7nEwhA22C7jsYn
nk97qCkUOJQdi5tZNLoESAQzdbpEICa54NKvozbS3xbtE3aOYUlnZpuKCB2M
fxuaI52eSsk6AIqoPHF4lEA0ot09hriBdYWxP6toDmqMWiPgowkulyzsqLSd
6+kwx8CD0RZqxL7wb0cixt+qy2JnxbzhHzpt7h85z+xLISnEPMEAyZsuA0RI
pL6C5rNOlFeMmgfoh3u7SiRPNMJZh5n7d9fGHuO/TmgdHcY5NmcS+Fcjk3NI
1jXt7QhYosMMfaPlwgDZBNuyiVHeW2b5AcAhVOh8uYwbT+2yQZ7d4pJtpkhk
nwm8JXXEAtJrd0w4+9B7jhQXaAX6+OGdFRRYjYyPhq9GSC+Y33MvbX1+Vy5Y
16BSl8PO/1awaU0BMB6xU58RCLiVecPN1pdddaDtty7DruA8amq83wQKT5pn
PhZCQfjABQ2EjHitw7FN0sqqXydGeWwFmg8wI7dUkyL6I01UhRdfNIIlfbfm
7Gi/enlF3KvxJM1j66SOAOZUu9QWg2xOPNia0nn4xrGWKhxm6wcTL6gJvcIZ
T8bNegjK7uCtQMLTyHiWz3O0OXBfVEI27s8Sv+ukGw6UNo6CWMwtaaaRnGOF
E8hHkFlmKVo9m9a3xgCB0ZrpQWNTmVXvgiPQbai7gpeUzLmdtCZ/WdcuruGm
q7360OwKTBsKLO8kMtD9yGPRAxSUeEm8VLAo436xUrTdXdUCf5z0Ix8lkWok
5ROMz7k1ca+KzTFfp+mDrY5MNA+kPbuxDMJ0W5g1Irwcn6p6loljTooHi2Pv
JHQEZzMoaaePfuEqR7ns5l/1AgmlBWy2+iPl+8+c22PFjfXu/n9/Ib8e9F92
VYvzB7JPAYd8XxQn1j728MpzXKUfTc8awzkTVcx1jnXhm+CJx2i6+WCqdKik
BEXCJn/TQo+IBrj13RmWCbnCDtQDUX8TPExy2asJUukK9gywrI0ItXHKCLFh
kVsUTYMikZk+xH/+jVHOpIey16Lo2tM18lN4tEQebHVT0M8EPZtqCLdOnukp
2d5oQUUQcegMwKk0al6TRbsjP3Byc+pJsSLvL+37mCDzhYiSeOowWLLpyIRd
nLCbtaTOApiUVFm9gjz8oe2cVSeTT+kLfDSAqKwsSegvDLb7GpJdNEc49+Pn
gWmFdY++93eAsH/Kk3FaN8TEZ1TYd9KE8iUJ1lGWO413je70zVruzvBZ8JRs
nrS4AuDvrrQgBmrtqSbrBI7RJXCEf9V3Y2/gLP1b7PbRTSRJwmRtsYCtvTSH
/VyYb51zsa8go5rzUErLC5/vIL/0VcFyWKaB+IxkNlJ24Td9j29UaWzufHX0
mWIidtQzHckh2bLqrgpVepk9wk2ovBtEt5O6A3xlBp2YCo+Z1CIrKGWZnhB2
53HxWc7DPHvAAnGrhcJdbvSnK9CnUTcLCwYKHSpPQKoPo/rgS/IRL1OwzX0Y
WF5nn1gbwXk1wHdsvNMOKhM0WQ/h8mLFZAsGVNyTjO4Xc230pDa2lMxYNJNd
g4k4rO5Smxr3PYd1ePUzWkn/N87/s2Ap6ypY4ZWF8MyNv1tI2WaHMmupdgxd
wNpBq4XLJb1aTph71Cpmv29+8lF0DIdxGyDARGKog3gqjRJ9/NnpZEZ6OSt/
rgeTUic7ssCHlaTxolVfnfShF5cEUdru3d+1+EgVteVIWBS1L1RCiL5l/ba/
6F/8VCDSH5/wDKU7eROramuRUgr+ZOlue0RWYPDCTfYPc+raOQCUjMVGzJJe
jO3ymOb1a4DhmzVJp2iPIqFL42bZUZXqsxoeFkNBTh6p18zyyB9lCiempf1y
tmzGoFWQIAqzN8THd6Kg+jjlPMxTtzBblfMD5MnmNU1sjLcopUQr5alDWRCV
ZoyKnMf8d1JM9Ld4PCfdCqTJ2zu/QeBB+sxOZk8WlzzNJGPuSgxg92YQp5nA
dAA5hE5YmdvRtzEwinL0exSHnMovKR6AVdro/79XsT2IWW/u8x0Xouq05VQf
6860x9Hoy2KFLG5BxUDcwAVbkho9gr8oYraU9RvTOJ0m3x4TXGlRQa7cl0LV
6oljDnMUgHDy1+FLGbl8DtizdskcvNQ/wEU0o0vSwGXl/6Iffq98CwvoG3Q8
A4dpL35M/2QoWYsNmPgskGzxWC382q8b/Yyhbr68T+QrTpfc8BfDRqbIW+HK
lXS0WVwWPY2mpAepiOKhP4DHxLJ6BNABek85K1LThAPWyGF2bK6plvuiNqRl
/oBFIDq9TPcCVORoH3Hi2BbU9YZY3lmWxzmaKPTu6DgrlMQUVTTGrbRMhXSa
gLcztrrfMsfA4gevR3a3TDquR4ErM7ra1FOMhXFmRW5zGmaPrpK6c6mlnomj
mrtP+ldaIsK8+ydjAoSmCRY6j7wScm9eQRmPjQKo52wED5Jw/2OkX5IfwuCn
9z9Bj3JlG4hJxUVBSgn0k8QYe8Sw+d/23eH7YbVKnZrXbn19ZxVxqQSTgjs5
ZP/L2NXLEHkU3kIl7pJqENuN56ERpNDY8Dlm4AJZCsb8RJcyGP+Kx44cnPZ4
8Qwmye7eCEA4GiU/giaZSa+CveAJsXLm+NDtXN6Nv4x9pfp9ZkiHHJLzJPeB
eiIrr19fKzcq1VytHS9xPpvBeFTIjIkjJnSmtbRsZVZ7N/zKnRmb0oxNeIS3
Tag2Z/88eE7fQNu6xjPcFocOMs2y5wXxvc5rKy4M8X3nYhkxE2fjY3gUDvIH
wjqWIVC6c3LDp3QsMklOjLGsNEoXV0p2+D7dUR57KVL1sjXbtWhJ29fZC45q
tyx8ZiukaiwNdx4tNvH7jon0IhfIfKcmCM7FkiYKnMYqOf40OtVB25G2uOqR
JIWAR1l29pmrYFlZDj7pjIyYvjaTA+7MeM3ULe2WwtJTM7p+Yu6htAfeVrlY
0eMz/eLlsyp840CpAMGQRjISDdIKRYFdzezZ4C10g2w9A/kBi4OweD3fsoSe
5VHlHqnnszynxoUiGL9ADDqh/pTJ5E8ov/KPOhkDp68Oh1GKLajNNMKKHhvk
cIg6Jx2iNJkTz5irdswlAyEMA+0/gvj0er1n8cigCTj0LsPjIw3EN9v78sdm
Z1Alx7pUxOeIYM3r9W2DYR+e8yECRYhTxSNWdmnUd54pIyjSvDpsvYFrLhr7
FnQ3aKdt/6g5nhd6nnloOkMH4OXinPm6/cPM1ekJmvhH7QtpIpOj5T8PUsr4
9nR9XQ8g7/dQT7klDQVinGeBMe4WYT7X0fW5n3lD6pAIyDRFCSl7rq37NeC5
XvjSz/B+IZX0D7r65rUnN+/7pj8H4vHhL1PUu4QDBRN9QiiVuLAe1j1JdBRi
lOhnEsPIfYuN/Ez941AqLCHr0mJ/nZR2HcOq110s2kJ5TRVPP6juT1NFPF7v
dCg3JhZPw+KhLSAvkeVXNXiwcmFvRErE9ivJovIEKB8gYgCSD5yiS/3OUnV2
fsl/e6AMNNsEINnYsoGt/kN2VfAXvz0UYDFSRyC+68RGLdIWNlx3jwyKFBmw
84d75BK51o8yxuWYLdK5rCuccqpAGkQgjmePKbV8Q9dIpjMYaVhMvwzYwrqM
Mg8siLInn74Le1MjHaC63NXVpH8pfhRBTRBmAM7qUkPt22TUs5pUYm5u0OA0
1LLG7OnbbcBFbzMFex2SdKIHo16991tWjjaFJQgKWFf0miFsO0bsmis4HSil
vMfZq73QJ0QqSHGoq2Xvwk6oxf6tXzS1AfF83rxgJ7fvxLy7h/ElypKYtPjn
j0fyBQ4Y1N8AvHNwUhqYFw5NcAXBDFbxXSvFFBCtn4klZ2Pm4y+UiXtqMxUJ
7+gGjA9+ENL11COozLOKr9UG6hLpsp1tK+AD7Tt31TFs0lnd5LCqdjIbBjO7
SopLaN6lq3HAegRqj78gJypHJ8owW6wpCqj5IxVPvQYaPlBevZYMoUbyfYDA
ORuyYq6qWgS/Qb7WnSgDO63u+tIqCwYXm3dYs9fKGF/lZO8j/myF7UzoE8Zd
etPFvkGQBy3AI6vmM907YNq7qpwFFmYfJMaYFsPBoSeaqI9WAZiHzmhNr5TG
q8b0ngoA0SF59h/Zl8OpmlDIrHsxaMdFu9YdoUNBZpY+QGd9go+kQWjY+w34
RaIWQY8rtLBqQwYnTAJfKq9hIbbeEbK4r/J2aXOyGgqOzzNeK8NR345yAAo9
UTqY8VBSFwvhxORCTt6pt0J/5335JLLNC5ix2JO4ySbWsYMfts//Gj5Im0jT
7hy4/LjTjOaTDI9u1VzWq8bbV/XzXrylhRh7Qy7M5yycg0MzCa1hx7BQacJt
Vc2Q84nai2SabvVQUtJQSnsWXfq2XK0s2oBMrpCGA1/lsPjY7O+bxzh+RNin
3NvMoa/yq8Ohecul66YWSO1tcfEqhsYmB1kCq2rYaUSFlgDoimrF4nybLrRz
sNhGjxJbQi/ZTPLG89YeSaX9++AqcSh3hQVNGt4njtS0xffnnklwq8+cuhLp
qSNOT/Ms5NzwPGjUEv/AYeLu3NmfIrMcR0T/mBG7+1nruHmdVOmAtYQ9JxPR
sM4P86COiWC9BO9TrHSuhe8sioROwUPs1LNFHpnmOaxYPev+8+KrO4EurGyB
xTXXhOsHs7IpyLq1834VE1TK4ZrbXkIiXs8PiAgIT2FYRoiWLXUn/TH6WHQF
5plgXtXvdZzg4WYIomTCgG4qQ+v/1vFB5BTTzjqm4qxRFIijaqf+mh58VXPq
veHkDgZ6OfXEZY4hA51iXomM+rG1JzQM6Nd/mAazg9/pubYtpCPPM+0SnAoV
FAPHuVO3yf7K2PkhOhO6QeeJYMOWSvYLhMDQIIh1gAqpn5ojAuZMRGvzwD1j
dz+FkChd87QFcJW81T9/HsrhkUF2BLOPuSKR/gI7toFg144ntPmsG+cVlvRX
3InORg4dK82UV8qpNUSROYS2GO4uF8id69bqKf3Zm3wx7jedOkzVD0C90tO9
16fTG+ZBegzc3znfh+HvUnH9TBT9ekEF4vjN6UhVhCt63aHY8zPg6lZl+R5V
eB0zGcBPziu7tDbBy6DQpOEOZdxl2zv+secSOxwZHxqQdXb3B1fM1+haIvh0
bW9JKqdJn38aPdg90gl9BVYHuhJa9d/BNwZ1LMSbdowo94kAY3j49W7LnMS9
CPiHKmfrEpCGM7wib+qQPChu/5Tlw9xcD4qN4Yx4OnN68Ou8p1nz7/y/PCAA
chqZGI1g3RDdH1q4ILmiCaL/a/dp95sIXgRBwz6InvmCZohO2PJaem55GW7z
7LthBsXKXVEvncSlEPOtS6Fj7qxpZUyi5tNAWH/Q0grKxZw0OJW+2F+udH/G
vuZSji1oahtbsOZbHzK4LHW4cLmnZtOMZBeVL5t4aA3NRHCgfiHWj9Gjvg6J
5atlixV3PIqIuewN0VXiKAGvW5WGx3bI/vt07KtYH2FY4QsG7/5a8iRggE3+
LDKfXr2Gm9iKuEp4g26hi5b7rHSKsoaJXVibfi9Opq0dlgKDACSF0+GgxG2D
lavh+yzzJcu8u5E/qqz0DKckq28HNpQxijZZpiJEoWz9mnGY7emxX28Pcc18
2RL4lleBFP5vcJNexr4DxjMfEfzKya6QfRGelSgrsz/Lq6nZtUOJVjmY4sR7
LmpqVNGuMR8ma6w+U56W/76cJnIixRpjZnUvQfpP946fIwG8fiHOO101LeB2
w4Bzj63GmEmqn9pBr1zxb8s+VpYnD/iLGghvN3GTY35fesBmOnarfcu8VQUP
GoVonapXyz1fBExIE/C03jaFzm66Y9kPJbft5qKdJc4Vqil8qSrolC/BHslR
Q/5MIXo5JFzfKPZVjPv3PiYP9QMMP8wPpvFfmgoze2zNh8KkTcjtWnZGVZ1z
UMh4ylGecvaKTrhsXf9gnNaqBdjrDrPl+Ew/27qEfwE8begmWfGr4gYZNHPh
FfDAT/krYZFc/KeMzk5DcWp7WlGbr8evnp/7l6h2IXhjY4ymkN3CNItSPW4t
i86+o2DOI6WU+KMoEkRnw7GiruBK/cIjlA3p0zYE3vSajIBnLzOiQkpRXJFO
W6JzpTnhH+MlGCrGwessF5Zrp3fkDsp8QMUel8h7oUbudPxShXQ/EtlxuhIc
W+DQXFBw7BQ1Gl+0MKlbRJFut/wcSUotXfKP4lP6f1/y/Z9Zw16dQNSRRWPe
uyjcOz1s4nEkJEWKMuFFw18lD6N6Y4aFn+Y5sHwkbKP+xNwcMjjO2du3Ngxg
CXZhGtwijrSXwmKWmHTFIODdm5Z/AYmFxgPdEjRBoBf4rsTVOsjyDyPuxIGM
8RRc28hzo+UyzyhsiMSkIXEy6jRAp0x8xdP219P2Ym8BZ3LRktwDiWJ+zg7Q
7DEC/o7DImXefeosnhBvZhojHPMLjO3AYthYh3CuA9HoPaywfdVyDBkCJctA
j9kzVQkpW5pFCgcSiID7D23+XH6ABqKXky5JiNSuvIpgvAIuEYAzscsN7/xB
8DGSGstOBOGVYfgd5ygKAthZH2q5tW7R1aqIzRJUAYhFoKk8OrcWIGy4ZZfk
mgOesJzfyyAPUQcAt0SNqQGn6n51YmIbTbOzZzKn7b4HcyMDLyoJslZtwKBu
UhyCSWaJK2k9VBp4WzDlSwCmd+zS/qF0u/PKANfCMrYyc1M36QynUAnS7H/K
rg0FFQCV09A6Gv3n8ujwA9suzZASNK6paRhgxgqtISQdQWZL9csvEhhX6uRZ
veZjIzTazvZ3a557/9Qr9Vig84i2UW71c8lenC6fliQ32AaogGmLD4KCleml
pNc/bmUDsX6aGu3lT2ROCxsa/HS41LY9HDUREiH2DOXhg+KT/NHRWq5XSrq0
xbTOuGr/Kl8J3AsLQuPeXeuWacCD5ajOc+g3ClzyJ2X4eWHoFU40vdx+5cji
G0IQTmQYH9+WmP2+gB4Ngn6DNPXZZPwpwbQj1nIPPCcioEkTmwhnJwwnrmhC
E/dnioLSJXmw3hiuVgNytq2utK1nFfjq81v7vqQ+dchWFDxbYty7eTNc3Hsv
M/aWyswriD6oTONqAXYm1cJj/7iTPYHW/MENSNKD94kQ6p3ctIus7tQVNdA9
te0Hc7wlvJrijnyGtpsWYZ0fcyjT6gwoVUb4gi/6eouRxODHGSnazZv2Sl+W
JsTR93ej31GiAwnyh99UkImxhLnw4biq3IjinwckJqFxFIjaetybVvFj8xk0
Nly5p8C4lNVJpDTl0rqZwdi6SzVDvOy3gwG8/mhuhoeUqTS8SZgsNLqebe3C
i26yWNAr7+g262g8IDYZhOuLEblRw5HI5RwEMUt5dzHTPvDnJTHGF2Imf3h/
LxqRL9ox7mQ5emst9obgTKWfZPQDO9AAHxTLCi1Aub03cUeiJ9T6toYZvMwg
/K9sXmRlE+c9hpK8HU2a8PpVGmH63x/rIxG2YQKzwGyz+pmlzun4axkXpKk7
uj2H++EbLRogWmqTw9DSqU9nnvARkZ331jk3UxqqXDBcYlQUNmfMfX2hzomY
urhSzkh8J5RyABX9ahvjZovleYKJCMafuqrPtBnzWJslYUyWU/jMX11M7tls
6EtjPOYPV/7dud68KwKP8e0j0elJQi5kbgH1AdCjqtW04AylmW+1FgDMsoVS
c8/YVBj5jnZoi/p7Jim2OkZholYIynjq3k2a9qsv8mepVgT6DowvsE2stvCv
Uy6oRnx5ugjuWAwPlMcKyL7LDUq5rHkVkU9c5yEhNSqohVIQfa98OOBQNXpF
oBov/LkXXHUyr3BnvUvwCn8dBbaMPyQIfIucvKXUsKEinWt9Teq91UAV4O4v
2fjb1CqiEgZe+SSygrgPGemoJnbA3idEUQrrpAkVJataPNzBDapaLdNBxiNR
5qBJPyiaP8VaWVFmJMvFcWQaBIiFEDhshUYTkXJDupp1uKMdymndO1mCZmNq
B84Q1dHYjtf8WAybSagYFgPARfQvp775JE1juaiD0MjzC9N8F/MIOfBTIDNX
tV8vumAgW5MyxcXCMCnWAWu+37SvJKQHDIjNm2u2C2ovQXFZ3y3qv8RSgynD
4EE9B4ET5G9kWiQZXcLvX6hjGUIcZWGNZYsQXH3mtqGhjpEmqTD0SAeIYQBu
LTdiIfTWOeVtK5MeKSef0aYJ/v/Fypb7oxG5qEqYxqXZ6rjWPkevge4l0BnO
oHW/A3udKMqOdin3nJWZ4cvzLzba6Y3DHDBCzZqYUtPgin44dBpEm9GMNwIJ
cl3R2z4b9JGI+cEFxcRN//E/ohzp9dYjyzEwjHB4JRt3qQujsLBDWpM3sMs2
FSis2OTZXYKOvAUfm1eQJHj0Y0fATJmWp+etZKztcR5MRK46Nim3G6SjiCMo
3pw1zjMxoDB8ckslaM7ZIfV9fbYGjYRHUNwsbYRVPhlMK2YYuQWeCWJisoqo
lW176T1qll0mTTwz3RZ/pGQL+YeEKrGMTcyS0TcQ7FeAdxxSe0ODRjDUpLZG
eb8YuFBqvF5BbD5/2lL6MTVFF6D0icVWkprXfRwzHLt+4OH+fAd6GcHAimEx
/Qdzsp5KsNP1IS7OUTTLRdMOf1WsEArXdq4ZOV5jDAC2MAwwFh/n1ckXbnPO
WI+iCQcmtvwJrZ6uh6XEc+Q56Enqd551OHEMcpnpbba2cvjUukJZzQZkYVSf
n5GN+Wkp+cd6pejlbrWVB/KYv0m4moHIy9mH3rjudiUhW8IUFQz1JuSjc+VH
ZdT6Y4PDjQk7c+ajulZnQYbA23SmUvoAAzvIV/GZrJn8nCVFB7alLchz2v+N
9yA0DzjiuZ4v0RiONZXyYGPPX/XyVbLbw4C7adW7Jcl62u6rz89i5LraVQw1
BRB+jVnpTKlBX2PpIz7wUFAzYXXgXoHgc2bHnOnn7RYXXY6lw9DrmPC2lK11
bTzbfl2gj1HmZ61/nn366akXV6MveenN26px2O5Zd4oiTAM7xoXoLM7FI06F
WnPBBPFBFgYpRZbZhYDEBbYz9Suv47PuCx1Lx0xEPfQlEUxnPPSGFkFSa8gV
pN65I24uKglK6Gz9NBRpv79EATTzbdLIHhr3b/uuSWb7DI0Q5tBuqJFAnkHG
JFT+akdSo3xv9/G6gwuqukz8V9ypIHuPunZkDaW3E6ax3D8ddDFN6t4A8B/F
ws4T/jmBbS+1d81mQvsZQqFIzKh2tNCbkcQRTXGJTljAvGWA/DLyDk4jjkx+
yT62bXw+t0S+fFXWYir+ZRqmlw40TviS6UdJscuPvs+Im2/xvc/6cVucXiyQ
RuTUKU8YEs4FFPoS/3LPu6daJY+eFgn2Cl+aLitLimrLelzH56HmfM3nNlbQ
NK/xQCCQQyn+aTtqEBPYzTy/ISn9SMj+v+p5kEhK6dDylpgoiX2ja1xVQQYl
hxVRsOh72701hDlJWK8pyCN0N/W1yY9l16Vjb6d6cemA/rDhPjOHw7nPQZBC
bd+A/HBD9Gi94sLgvNWOUZFlo6DYeHSnm5LwGfLPxfjEX5o3JYrskInA6qjC
8yT04KvJLsbKl8hOLWC0dOQ+Xgg7jxVl1DFP1wmwqlTpdN42yK+ejGxDLYes
SfWOtVCiqbK/PpW9GZjucoZwJxjjWTpgoZ/zPRvZqZI10xxsbl5EZbrb7+wu
s6ApXS+Abibg24SJ989MiZx91aIDoFgHGGdeXWGa+QGK6i6Ebr1rUTsZ3c+r
7okgF9JzjnMEW3PKHgqJ1hWQLOpVL/XoB034LgEVl1pEhUDkdOrUpl5Xkgir
DJ8VAeAlnlT4uywfEQWx43Ki94+tHL3vdY6OOlxxPDeDKDaXc6fZO2pOnCVC
riL8VuNJz9igv3nVeQyP6Voc07T9kyIci8X/cii4FhKJGIzzNgLoK0o6/afI
CcCnNzEgZxO0Ztu1zXJ5urOyzsrhmNuKBpUt6rOI1KyQGCwglhPDDJoNI/6E
F1rY3Pfw/BVxqnjQJ3fXqD0ZhH+HSNVq5t03ajvTOhnCHMn33dQh6F/Dt6jk
Y4/mKhtojkfmNqMK75aazaGnK/FF9cjwysm+XFGvZFBlUnVs4eZLXLBvYGdO
Rc2vzXMImpMjL8lgRIzUCVcT9/Mf23dwaktGgAJXsNmZ2nV+TDPFhOyoIU6M
nRaWr6U3sKIUDeDrbuKNntjqL0XwZcdLj3Z8A7c2JM3sVuMIYhQayMhnU8yM
J8AaAqRralxkFzNkdu3jTRx9DfQy1YSID4JNi9/NabBevKw79B0LKFGbqyKV
UvpQ2KUM4KIuqV2Oo2OfBWugbS/8F5e/Mv7/8khXUS6KFmrHmGDrnHS9i1n3
w19aVFuYweVGPBrOXRPvoLlB5FTuwAryvpA8dQEBbWboB5d6FeqRtfvklcbf
Oq+BNJNTCzBFYkSljtBdXzH67P2Zwyf7laq0AnYpajd/wwl2yppxi1C0BBad
3gW/DfPiOzB/pSELSFhm1cIRJwi8kbF3sVP9BhNBzT0OlApQxktGzjkPlwbQ
O4/IAw82P+WSu6ywIB2cGk0jwF5E4mMA9xjuWl3x/dCHFtHL+kk0PiNiAPLf
qvsNswK7URiqLCurVYDd4q2zEKkSHPZ2nHSZjT9OHFQqANWt1Fm3MHBgZa8j
SfTR1BHA+F21bW81ob+NtjW3wfwiDyqi8Ap/SKizlarHyVSxxNXS7QVmw/Kr
fEPBII+SVfBloZpJZPwLPNP6cc8dP0yLcGqNc4ovwjJO+/6LVNdCtVkv/xzq
jDZkSMx6uEIIqgRUjWRRiQ41i7pbjDIn0Ts1gjqUvfIdSelp1kCBq9rpLowD
g4abIrtVGnKDA8DiNVltLbPV3hSDv1GxsMzcTJN4xaEApWiWLysk4Rh3kmda
tImCEBsZpTkY2jmfxHjKx5S6ogxO105q44/glBX2JU9aYvwXiLQdCOy38Gep
8SO6IWIMyjiqdc+TX/+fo+Cgts4Ridn2LI53JXbv43uGXkFXqD3oJcJ5in8w
1QJzjBYLFhkPJHvlMueHObdTZp4b2667j7jKvRRAndURtJ9Vlnev+Sj5Hoc5
5KL/hJFrssNcuMErXwOKGEtWT9JrxZoKP0FJVq2ume1207r1LldS4Z8Izk7C
rBUtNVH0TQZ4O7KMNtBlZd5IANoMeyRjl2zWIftDN8bUJkMDAhfkFTtUkDIR
WLRF4uYQLy5WrO4i6aShYCUVkCMi/7V1bLWQglDEgbWxaSWYfOeh+FYGnnM1
gmmViUsskI0+xVwBjg2KafM08KDOsAShWrjpOUmphOyNc89BNXEg0vobYq5b
ElDJDFUmWlqmGDLTA3QiSgXN1YHk0JIrTvxGS5MCiDG09Gl2zHNzvezWQ/Tv
IDvIjN8A08HCmpHTvLoY7GV1iqAEJR7U5gdNv5MP/zYD9hzv0ApvER5lkfP9
zE9gOnAQd2iNW72e1uKIDF0POt+76e1JHiZ4kYzt77xqxuvx0LzSvNtIZ1yk
ltDM/nW+Ng0QcZrDrkEWBGupoOVYmELoKKELhpOgy6GKUOscAEKb/D/41s8q
qFznAOZGZ9graOFG7iWOKKh0zjdc1rHvdvBk8nI8AKExGKXQbbNSRUxp7RYK
nB7fHGhZ9jBTVBAxIH+Tj4aQgvLk3JlRBqn/ST/t7Gk1tvverydt9vlMTgft
Ym8bBtxA8Z6CWmjuJbS4f0Qu6Jph+g+nDKOWa/RCH5Nkb7F9mprdmEAh4UqF
cgCQCM2ROUSN09sSce6G15Sp/Zk9o6VUtkhoYQTI54L+Ta0KkoO/vxHClJ5U
VOkwms5N9kjJWlx2NrRPGfCNVjhsj5u/I6BGW4R9h9VhWVF8/8b2a5gT8+Oy
Wa3dHOomj3GBCb0w+xBH/58NHZBLrUJvcB1sDvt45cCd+0GdjAi9yETWPsHf
J+iKamgkxXuGoDR0vRTmKr9OMbO+I1DZrGHBBJCb+zSafbUlMiotiQww+1MT
WtYkyZzYxVfU5oinAMSIpC7c96DWnyMtoP6Vo00KLFjhsqQBhBK58uH2QQU1
oFEqqEEMMWWxPvbTbTZBSHOEpUoCGr9wyuUw4OjqxeCwT8IIQ/KtIBgQfvoX
O4t9FQQLiemvWvyJvhks3x9VcthWLOeseuR7S9MDyNyKBghL1afyx17C4L6H
FYzoOB/awa0LobiT+PPomzdbwub8HrzkLfJXcLYaGf/EWVuCVnZ3sR5wt8sU
JB0jd6wht98Xvz4gb4+5EOHiNdCUzNYhWc5VOOkbSzLdNDU4vRiCdRc0qUio
6GYWMqx4WRykovrx3pdYcPEUPZec9suWWJoVBzoVBmRp6fRgsczuyNGz3K4G
e94/h9HFF8j9xCsbCRXFejpQMAAw6/wQsWDNexNL8TwoUvcLnxnn/IMXo8Rt
jxui42SAHI+PfqQKeRRpFXFt01Nt3r1lQqVZoLx6EF7EXDXQwkH/PJRATWfy
UBwAohYg22Oi6ZzDePmltCj+C4th1NPjFFYE3aW05ob2PmRW+dJ1bOTXv4B3
JlvvW5K9FUsM6cca/GUAYUVEZl2/5jCZE/PMpAt31v2cEg8B/OpkPZYjsqcF
vB+AgtHtNwXJ5KjbJWgVRyHo0ky7aYET4HfE497qYOM80BjLMoA8tl1YuwF2
X2Qb8kToYwTbsSlMMSgpQyUznY6tnvKezPxsXosjP7jbYclvlYL/DEnDCZW+
wW0me02iZ3nB8RW9ZUoggeVWEZmBaJW8wl+u3jiHPVe3vMuI4Aory0KCdFxf
R6NfbH6wTLfnuPOyxO4JkLgQxXz+HXlQS46oDD4cLlFIFKgs0vpXDtxy28jq
OCMd3/+IpG7snhhgfwWl5lIS4q6/I5zc/R52dIUz4hv+NFj3zY0uWk1F4hks
swLcsHrF2AVvVu82wRMKzh3GjSqsOlDSlVWtsd33cQKSmEfVPnVzDUkkKLbX
2lMCEjbum/OFzlrTp93k4wr3hWHCOf87l/duJY+Cio6Y9EBgV7udY5e8Jifp
1j9GdVsuppSprnphVgfojV0BDLGUyk6OGThU7UDWiij6aVShQG0TSESfWwaT
6pUETOmLWUlBWDkyjp4lizoe3EHoHlS4+6KKLwYEkOofc5eyKr9EsrBGGm5K
yw2Eu4EYccrieL6bR2Qy33nO0oKCpAKDNzKZ2mqWRku45EK0Qwb5hkf8Tynj
4BLIeZQSjBaP5FcEUCYAVAS5zlU1cNJxgmGBCtgBa5iffwje9ewrDe1N31Tf
uPKRUDqMMg4HqOiJEO+fNn+7vWYvKtGsnitJ0XNUpdJzMpaaqfeOTkOBneRH
ErtU+PQgbDilGsn2LwgxA2Vi5/hHYaXv1etNPg0e7YuOslNpmW6Ormx22zAU
iTpTfsdM9pyAjD3qB9f2ngu1wqQpNdQOIDpt657JZWs2FPIYpGBdkIDP2t6S
GSTUWPFI3VSeS2drM1UaR5A05NxVh6sdBbFi2/qBsWQvXLEKiZ1SOCN+neoz
0FaTX7jhDMrbJV3CYWMOk0DmTcScW6RfvpWhqznewlnlSMCWgAPVAWKgCkEk
/8j2UUClKssj3AejwhrocH3HYW8g4gDKatBL1p8QGft5ODO563Dlc+Q8NScw
Arz9AAu8KK+RiV4lCdfcCQhh1Yi1OUgm6WSauvwYeKsqiM+ByfmnpuaiwibC
z7ydmLjG77uPJevunA2v87EKyjqQpbTz3AeIFzSazRfROr0qeFoKevkRxymA
6ik/BOJf8SWJDaPBaWLtv/N187UxIhY3/SQwJaBJSaRglcYAvCrp97itM9KJ
zBo8jBPV2/RIrRO28zBHV2iCmyZKTPcwmCF0xCwAJ2icoe77yzhF+HtZ6tcr
nbUgq8ENHVMhJQcaMAP7lb3R20JKRCAtCnac7pDanoV9DrkMwSP8DxSF7khi
tMh1R/0zhErEFy6Frwnae3DAmiijG81H9nSltY5Mp6YG1Lspeu5wYWeVWfUh
akz6+pdYlrmYOD+dENTyaXl5MmtOUjymCbVv0XZYhU0017cLK6F3M2HNe/Of
nHdLwmWT8JxGOXCsvmPu2Uz1bcqEoX0dxDXrOj8zVGERX3Wii2HDIbPdstKS
9FmRcdVi+8j4OwBOqgUwkMD8jnVngOesIMs2BHGPem+giJMejM82hSOW6coO
OTALmlI5E54Eq9kbyJYm+xw8+gPnbdELXt9EcuQPg9qBNqIe7N/DzNAGiBH+
1u0ruW/Ik997Zoyqw/QMUlqVTuW94H56laasEPiSAJYezfCYkpcEhERw/aZx
xciKFJ3s7mugOD9u8ORRJnptN3PNxXpzxfWBpQQ0LD+vhmD7SRBWw65MKRxj
/folF/LpOxzBaMrpUQJ232Ol43uzKLz41ac7jY7nCYTmgzNtFXD9HZjIVdvw
8c7XG3mRhGNF4kNQiFImP52OV+ir3/X5/KeSuyqrj3CbTQFUPnrPlpu2/jNr
S6fNZOEcBmskS3+7MWsK5q4tZn7pjtNfsDzTAO5fXBWlPjsIEW2NTkxiKRsg
nRvKrfZAWC/1U3voOa+xn6ERr/rpY5XHUfRfieaeHUIqNTapTPoMaYFyJ18I
5onvvoi9En+wQmDHEU8DG4xauUj/BWRhwnFsF/gYzOw71tZ9uHPMyY97nbH4
gPKQlQQ2epnPl2UwuCPv/NfDbO5nPaMr4tVkdyU5JDM9QUiLg1XrHvsfWyad
kGE2VRscxC+HwQVCY2m+Ah/6LqNKuQsZgU2vIgHkAmYuKuzUkBRUDSCmuhwz
gJWfR331fKev36DSamI1068IM9wDg9ICj4i7QutNRr7TRTowUriSg+RLRgPH
rswB48HmMGiqrvlY6MZtoR66LSlyIPnzcEKdJJwqWBsU2xbObbHTa28/BQtM
v+jD3l2lBSNsIMjus9dUkqVIOZofyc5AMrp6s7lVhDItg2SM6YlXT/TM6RSl
tnaj7r0hxwKvmxIawdBl3svyAjcJWOcOotr70tlNY9H3fPeO46jMv1LxDnu3
GzSfH9CzKkSQp8BTrYTJpK12iUt9kT8jNbAMx+bNuiz50hyQpT/nxoWI20Ht
j568MQbE0RwWmosYZdOXgIOCDBaRo94n2hFOwgFUlfFVBGFwKKvkxhfnqAgR
KvdBEiiHiKifJ90nq+NXg/rrs7WtbkFdxE6rDJFlSNLzaDo+JiDZBaHzcDMr
9pjdISrcg0ePbVAiyVPhaHkVFFOh0t5vhrtaexkeODCVsJMOdL+Z0DIDBbmF
NbqFcTMvr4ce0YimRfDxoQGa3Ap531G0ySOrDuly0lrpMaSwLAyQ8DholO4O
vcxWOLxI2UioXC5b3hyX4K8EfoQJJ9tiLz0Sl4z0MgtsmywJOeZRDcPgR2Ch
eG0IuDhDKwrBxgCfyhBEPavsmdjcMpGO+rnOKJ2qzC7Ut53OsXjyA8Ri8Bai
cm1ecuHkaGJrHuJ84FOVTPNoyjwtzt0Zcw95WKzqiJ0uetUPSypXEXA70U7h
9xFEUjSWNOsZANjvQtgFwTLOpwRZrz+6A8PFxw1l++ai/19kmkxNlFW6Fy4F
OHVf0bxOfvyix2hom76DR2XAAL2FBjZbACNRioH4iAty+Yd16pH2JN9Z5PRW
8SaI1TrL7k4RQXF2RisPq0fIC04VxS2K4YcxfbkfP0obyxmL6+ty96o7m7pR
0inxV+8t5AXF5so/k1+w+U83f9CJZ5fYcca2gc/33ssd6VdXcbuprGosGcJD
66RBoSxHa/7g34PWaG2wW6ltsDeQEU1XzF4421ZSgaC6FEaDHy5UKGlQHruS
/nwiy/9u/xSkP4QU1+d4haVaBieii+HLGenOuEU2BUXNn+9m5KqePyo9ULK+
PWd85vOlgCt1RSYfinKs1VOSYQ4cwYVy8/JUu77XwEJGk139MU+VUvVpKkBd
yBvc0FXg3Q31Q2leOdti0rBT/l2I+3nvmckpdj2bkwjbD61echSBY5XVlNgj
nGl0qIxahwbEF3yYG3he1oL5em63/YVOXKRnw313V4umF1XuNA/Nh+P0Kzrc
tmf3zvcsaByB4Hw4OxtNp8x5nKm4pPcTvKyp64KfJk57U+kn9+pSUKe8C9tC
8r9HjTCjHQ4v5IFUfz6SXlAWt47vEe4UurY8MLLbztXnuFFWFRSwG+K2uTRn
dAIRSL5RwnIXnvSQfqzrmE+6spYOk4EBv0CrCUfjEQxR69JnOp1Unhuxbh6U
SDPdG5LPqDm+T0XLY4Er7iZMkkw0VicAW7jfw+OX2377kiy5HwKIaMKVA5KP
8KjKhsuOm4LZ+SOejBdGJcNYgAYyuQ61brKuW0K3FJT8RjFSdSenIA2rAtRA
Ba3n04TSID2ku7eu1urSVZ6P7lfO0JqLDaN0aC5FD4lK7/InisSd3YMvA7Ai
YJEkTJWwABV/H5LVWtDunsSPWIb8dBayvvNUGGqId1N2bX4242lK8IzS8SDP
CfyOeTOJuIPSoK8oluhjVM3Nvdhg5owfCIJT9dm3JWBPfnwY9YU1UB+IZ0aC
e61kwTfEqC+B5s5JbRtzUfJQA0nO/tRN6D3wezagEKc8sdME12T1WecGB4Cr
3rRVWl59HQz8oY4meIVpIuc/ReQcuPQKekt6HyvqTsDSB5ifYvIlgzE8uriQ
FzPCfZUsNmw2pIa4ky4Mg0NhtXbpnVv8/i7FE2DuLkcJJuKRM/szpiri5Sf9
8jSgnyv8BhHXpuPScJ3Q/WBmyEFxJq0pd7Zfcl8itHK6yQNwNKy85wWGbZgX
pKl+nY7qTee/3XYu73NlB+Pab3LewWArcxMMawSKVxmkKzqOjKAir79m/T92
6bOu7EtrtLGkBpMPaCNT9ugen6kz9jGeDXl782dn5XJfbJ3ntWPAPZQIZ8FH
W/Lj5mP7D28N5aT9I+OJS6TiJ0zKph7JbJhEVz4/ZwtfCK6uW8hKKDX5feMy
u0HkWuSfBNwZvejwxONQDISMWujeSIQlTv3OjDrku+IxsgNdFGP589V6RUIM
CaahfmuIRVlh4QnQJLPvcfROkUrx/zvmcj8v2IsBcMvSDq/WsG5LyAYVvTSd
C83+GYlB3kDlELeKlnLNnrZ8+rKibW0GIqbkzcC0bA7yufNc2r1kHINeQBBc
G3JRDcE/hzIsFvwaLPsBXjDlDsyq18etyvT+hGQ5HLGF4lnu/Vg6Iu692amU
plJFB22Agdo4Nn1tXQpW+O5DTk4m88byBuvZJUULrP6mNOpMR1WvE4PtbsfO
3rtz6sWMRLDE0FUz8GUMpxCQKulF5q2sAhhf1wHhw/GrZRatMGBBJuuqb2j3
mDX9jpWXsMg1E5+aeNjmigwt8haK2HHRkZpDixEdFl9Mk7VpvhRur1D6R83y
d+a1jcC6gEDzWZpS492jeB0qpsYc7goGrec6Viyg3HvRstJnobn4FT9zNiuq
doP7xcYUlKFLGqCFFIMYOgaf7eUhgqVK0WBADFpq5yUKdP6A1LRS1pip+sy6
8hnWgjFz8qlRvmaXgOGq3MrkOtlOybgB9x4awnqjEJGNW+DYz/tsztl3guXz
CAA02SuWGCd1JS/yZcF2Vw+mJFWf/3Emt4U03L9BypUu+6l/xheTe7b56djz
ew2sQ+e5ZLmvtGEw4R4LAMhbk2P+V9sp3IdjnZPuHrVxUSCPwHET8CdCSPQT
aQJw0CQr4urIqd/vc7YGVBvymXaA3kmwsbDb2y/AQBbbGZhGoCq92yDEGGqF
f4qxr3oHCHzQn8flp+iJB1cFaISvK1gUrVS9J3V89knLaFWxSMaIEehzSRpE
wh0u8mKcn8K4FqdB87L0M8co6JcxYXBPS8S/y3g5sOfKW2e4OqMmv0roZ04k
J+0ZwsNS6orVdU+oADsmqEMFEk1RGRzugDGW8Xp32H2NZ7+m/nzTIJDpMABA
zbHkf4yvwTSDjqybuZcVMIIOHwLjhH2xOyciS46t0P0LxVKwOidzszhBZSYu
RJg5msvyaQ1dMpsjS/6PBLJ5mgJD3NOrp7lNaSpHsBuvwYLaKbB0Ga0bZE88
t3AHCsz+F/8Z9xxvlJ4UpD3PipRSBftj2QcMmEqV8Wrk/DbewZNgJcGzTT31
+7gyncxUQfSROWdA1JAYlpvGOGfwVt7nR2RzHgXGch1/Uu3IKd75usHHmP9z
9/Oe/g8+qf0w2N7WZtJNTX9ntmlIXXdZ+imzyYh/ddyeHCRifBBy9lFcLJVo
5h+9jXVcH8PyKpQ34HtaC7OuEmTKeYdpW6kGnLyPjEtqkDvRjEvhYqOA+whm
+xbsBw0+v2zQ2HzgkLvC20pA/rHguz7pio0YcJKVcfm6vgpFIRRzo0Alg+6b
4orwBKktjhyh6CTd0WHV8XwmWVyge1mgLj2QJbrcTGW3FVf1yPvD/1VfUuWz
63QHWnK3BtemWDH1MGiAbblNONeTCmdEKcmYf67gs7fCCxqfvjQYzof1qaqY
gEpk56PJzKGY9Vsk/VEOiWMU0iLEUPbElvjRw9pxxHagRSE8J3uRPNQx2awX
lWBr3zR9e8R8neoMNz7PDQI8rGQbwXC5YJArhr0qT+eenM8HkO+FN4aJGihM
Y1S8ZzTqRUosyUI0+u6arnfRrKprQdu3NaS5UJF3Mp098/gETLmohD7iww5W
b9I+zGdUD9tvsqY9FrZu1q8SwKhi+OW+SmZlZ8H91DxfPrqAVkuZdf2hJzCP
JOzImweYFLITLmN3PeF9qwxtkGw+nJJHcnI9t+g3A/LzXQjXN2nw7BWaxEUI
audrr9j6qCJc1ZvHcYf1eNcZFA30y712x2S3qu+awIz3Rt7475HJ309w3BZa
ZAdhAf8lsELNvyPUrZsoVsLPpBDnHAEzAsyCe/E+lA9voIobsB4P61pKqMML
8QN1GPFdZiHsHPGy7KkugYGsU8d0EBc66p5TLH5EhfoGCXVO4Q79dVdoNGmq
zPog/cCWONgUpthq46jmqCabe/3DJaft1SQz+bsnuk9L6wj7SMV1YS5G6S4b
WW9J7F0ejKDONqy9KmrAIBgHSBcYMnT0CrQoVcu1CT2x8KPsGsDrGH+YmpH0
wA8lmwmrWrN0eggOyKW977IaNq5cXLR+LS6asRhLGUMPZpl6bewS9WkadXak
BIDSLsKjiQ88znuPFgfuwGPk0FZn1JDHUmA05tmOx6DQqxNbm2q/e0Fbbw0X
zIzWpTPnPsq8HHUVIMi7jWwVIQbEz8Rp62be5cuWRAOS+0978Ht2FBsqxNm9
2YjgXhLjTiLACBK4DDGjA1S8JljIjuC64bm1rDqvGMh+H3zROanOYeXO5esg
PzZX/7PfkV+meGD0wrkSBVbtICK7zl7hwHxao54XGWd21EeLfcyAUKXVj29Y
X30s2xXr7S0zrH7HqvgdP6jcD00GG5BUI0Piu4WadMJ0pXq2eOXqPk41sO0/
p6oTcMpRh+G2GA5actHbhn7Fq8BgRSxwWnOqJ6CKkEPxfR/8t+f5D5Tb9psH
2i3H0oNSxwflVWAk+pOlTaAvYkoaz5kw5iaS178gGWwzJNSKKj6Yb3E5QdTB
jKz4LpmPxuHA22YiZo8kIJo7DZ3AJiuzqto7OzxSMvaZ00cnsRxS/jSOXopF
/otqygH2sZmOiHxMD8uRLUgt3q9Ung/n1uS1/v/cEoMuWi47lsaqQSrfs25o
cJm19meHO7++tIkBcBG/SvZFYyYlPaaTu70SBBJznutrcEX03/PSsm2fhkkV
8c5Hq2eACJELn5foClDQKG8qOovKOOOCmr0fBW1KKQXoBi59Bjm0s9vMJpSR
5oAlB0VLlC1IJTA1nNV9accCc2TVWwF4KvKQefOBRHOSzp+oT/1Czs23YQxX
0yYC035rBzhm2caThko4a1XlX1OHTpiZQ5NeVvgpPuigj6+sUukI/+PwP4eA
92nXY3Ocx9eUXuWHLUcL/Lzmz10EpFgORFRY3MbNEgLhMZVCRDsZugYWtIVM
cyVbeINNbXC5MuSHhMn2MiC6dyjRtNIDPEtQXoBt5v3eH8X8LOCIwLqGqAGK
9LHGr16mJACmchbfmn/3NT61EVksOQiIIAzQdENPajij0imrnufmKufXJYjj
a+CXYrxW7J/PgV2usAkbwnn2ueK4CZAVV0ckltVB9M9xuu3GgIgoiXLSyu5S
Of3Qtb5NoX00z4WZJHss/e0e7r4DYRN/jAUTZpNH4WN9b5C7JaZnlW7UBVq5
XUHUXIXBiQOb037u+iP8wlIwzuTIj+BmbsPj3dpUx9TYzMwPuTS//11zV4cr
R9OgniT2dhMGysnZhrb5dKD59iaBVdmzb55N3xQ9NBc5u2FZ8P+HbdFNqGXU
3J4VfktTTWgn6kp9OXOsP6ScUEFhrBGaFLlqGlS9hUF4UoQdqajfnJrUMs1c
/HlMh5O5UjWnztZP4Ph4G+xWAb1LVMRvqeHXgYy0kUF9SukZ5UmiL+8p/YSQ
taq82sXou0ecsyL4yzZP9aaLY6Q7JhAoF6uCsZ1h6ehU68muOcozK0RBPKgM
WEVtlfrMa5ZbcBwJByyOj6a9Q9cPKNkaRnE9Km/IMNWtWUCNOZjr+3zJuMWR
ZpRf88gPHkODQnSvPiMq0/sErrXMYtA2Y8XozL8gWMRDXc0GkJRBs0pLchSh
NvwDov/OYjzDx/lT/lG8+Z+jIAr4UAldu+3fEaHVmF/XXPRcYUly0Fn+xf4f
iGWwpeoMhNFS79G3MQF2s2MqcJFBzhdKrAapU7awDLy19o0BrTEUD5wzgrQ/
ESOigSylTwYr3pQDUxO/PVS3zsUYSRpK50VbMBp8MlMriFbAVzHYvfGKPmrh
7+zsKTM6Kix89C6vlm/iJRhyki/VXx8MB+z4lEtJ/jhbEc3UuecVhcf8puaq
oub6j7zgCE+YQ0C2BSpWtYWJKwGSBWRbe7a6JD0emmmNaWjTzmt7SFH1Nzla
enc8ybBp6ork90dsrI6a8kfIiyflV7VcHD4YLQWKR5Cdrt3MmdLNSbhyRDeP
Ld/Dwva8alY0+Z6e6xGHCX5icY6uDIw95ZAo8UoTwCm8tIpSDI+kDA+MyF21
Qdu44SqBmDw3J7UqokWYye8kLsSGpxI2eNpy0ycTbQvFkPZakYbQUA5+za42
57okOsPk+3mkdlUdz5duzaKqu6F9460lJzLxccFQt9Il7l/Ej9+gWMzA3fOm
/x3HByMh9yg3DDbsWr/MB4YT/MUeJrBLG8664ft8iRUommiHTG3PMCJmhz4Y
KXdL7lmoFwIE2ybYmt+oSKaldr464pUkt595Lfb1KVS6r9rbW7Injexqn47O
6sAmfjMZSn4GLObr50HCvriJYF55SjFgRrBOq8FgLuXLVS+N2vEkar48pSFJ
hmMYE1Icsw1MKv51QefkOi36UKJuIY7uZe6Ixk21bXguJ1JkNSdXVfnxhUzs
YOHpfYEenmngipUxqrw5i6sYLL3e9QOVNc65k++wCFRk9eqU8gByNmZzcwBx
MfSC02TcGndyOJPqvNbEKq3KTOHHhIpljCu6/3BICcqihdHa378jBwD6goaG
1yGL8iXz4po2OEoNM317uha/uGNQjI4k5jjdpA60gIzbOS5fUrp3zSwMUE7j
wGGgcijNwru6l4Ul8IZc5H4mw0KVW5nzDqI8O/CdEWYQ4Ep6iRhEhq6j0abU
QyMOThHyMHO3q4ngN0d2uGXPI+/GqxpmsuEA6z8L6c/9BiZUxcl9shbHliA3
Piv0eAec7SkjRl5OoF5ujqkZW6J4GaM8rnoTTFY3mE+tgtmgHLnbJXgO+Jd6
v3Z10CbMT0srT2DOCQis8WFRytSmfQhUVP0yq/ygsbshC1AnCNl+jI07jPUo
av4fsf5AuashO0IdB8oo2ojsGVtZCPqferakVWRt4mVDFMn4z3x1RH1ReJiQ
m++T07qU5vZTIVqW/ivTWj0XbVkmnMSxqoLEZgXOtx4huf8BEZpT26m9SYn6
GFKoubbpKuRvDz25+shMBmPpKTTw8+4BANY7oKS5rfJWFVwn0mVUFo5s3/34
Cy67v+TGN1k9ZCBiV7uVDiidA+2LtOXrNnXORYB8c2CxD1tNa1UDnjJrNc2s
dO4eBJkRLpK1UqR+/7FeoUZyc93FgFdrnNR0+bE84vljCOv8pb5e/WrMjZ8s
+BNONiXhAxHwEesEJKIw+vdVE3Wbr42/IErmFUoCqlN79Z1uBHexU2jgvDaB
2rfFY+f2xT5+V8/E83eoRvf3qBDCgH1c5TsOJVtMCKFhxwY7qucb1BGYdGe4
IOUVNB7sUnnGR1oJ/6ZTuH/fkw8Qb6mr8OKSH1jL3L56hzAJE6Ruzmvoimbw
qVLKYtvYWlTH2YMW5SCbC2F3ck6MinMMcHqAWAnjuofaX+5XMQW7fQvJrNoj
7lZAjDfvtyWIQDafyIwvq6cPbsgddeHxWQlTAPCi5M4UE1RL7G0gnc3rs801
TqBA+DZJFad9U8lVW2p4pkIaCVVjCzVRdJq60PkFBPuS9l6UoRjdFSywfU/d
axL/xLk90PmccDxYKFyhRcFJF6/c1IRccDAeB86OY3Su+mJXggQRpbsc6r7c
hXT428gYSP5HCHSo9BOiryn61z+Xlgj3stKk2faN+hGk5/Qwb52GPBLZVxeW
dB6yWKthzBTEKD3tWbPylxKDj+r492KjMdgLHvAXrUd+3OaplyokG7+zCTob
tTwXomrBnV7FXNX81TXgHKu1/kWpkvIq335e4iZasbo56fCBHevkxo8g01dh
Xo6idtcT2CjFGR/z/u3+kiYpYDuwc0m1i8M4RJKUviQnkkxz1mQC1U3B14GA
dQSxVvQl9mj2V+9dkOqc503PdKWFYFPmSER68Svdh7/8D5AHExnK/1RKG6UX
Bd+QVes5yz2cYO5novt7Iv3wUOr5mavSkU1y7OIvP62u1+gZeW+h3aW6Lzah
H0Rh18GmEBvGAZZTzou3OPM93C9UAaVn4ohgcrXOQDNfF8toRomrNu/KGZwW
FnnpvnPIhRfAHAYPfw8NtmQYHaQOdKAlbQ/UNVUwJfUeQifKzcQ6d+ELM+v2
sAcKaZrpeSmrx9A0zET7s7et7TRCV9Y39qIQ1fYaptnUTJ6vCzeH8DOLPw3n
SZONwAA9BkvlvxOxhAyIXqKT7UT4e6x/G1g+KSQvAB1Rbx2gTFKOntrT6Bv2
YweK2R5T83eBkuXarDfuxWWEyERCMCICwcoQ6gk2gDsJwZMA8dUcpZob8nIS
+nnkWG+Ye9M+OGllszJ6Dyfv9N9Ur1lhutUnnS0mG9dY7fLsctAOBhLox2r9
Ms1xBUfqthmE5pFZEsKeh2QCS3IO3B3LzzX7umtmVbSU5OP/xYyUnRcnbJlo
zkjbqyC/BbXCkeErqDGE9iG+qAuj3W64TW5CFAmwRIDVE21xCu7cqpL9/ewu
DoFSRvZtus56FIc/OV2bQfh6nC8iWNTs/WgV6hgoi3OtkMF14Bim9UjpPL7h
XJTj7Nef9TCkhnq503e1tCFaNfKsL3F5mKl6wzS/PS2UdkOW2a/YpxU14kQB
cFFqT0DWt2z1tKi+nxjgaTtpazHfteX9M64n+lZWxF22q5jeikHoHTWJuVlz
ac7rozePETuucLcfy5nmjoyM7nEaX2ffk2KPZKLlwOar2WbRLNt7juCgpw3x
ilcObKGs9WVk3Db6LnJBm8idpmXbTelsHQFYu1BTKJK8ZjNX4N6d9LOPA33K
zrYxgvbM21ka0VK9WDaJnG5UXdDJCCX5nvxrmHY8fp8aouLE8QNC7i4sXSBB
koTF77SsKteAf78VlC4QZYpDFFVcB3OgFG3+NS4bkwo3rgPtAKWAMSyw7nhV
v0rq1XAhLtR6uzAR43I+zrh33m4rO1UcDHOcY03Nhxp7RQzRedLbZz/MB7tH
QuhH1Ox2yExTDrnrzXOH7SPK3RW4f+cGbpmL80zTsLapaECBe+Ak7NvMPuJE
JeRWMX0Nag/24SGcNuDUppyXzqdugA9gN6zvV9E00AP6l2q2VWoMuCm9HaOy
2c3zdwRPqn/AWTcBdDQhKMzzsFe/ZBWwhyHNjOoUV258WxALZBauoFOHKW/X
+e4VY3ZA3bTi9jZ1gAsjrtZv3Q0oodHuu4huYYXKp7o03CcxplR9Kmfsq59m
aN5cZkXIkc0GjIISmeCJS07RUen+BCBfN4PbhU4lv49qEPV2rHgN3zb3N49q
Xy+ODpJG/Udqx13fjq34r2PEVEPcvKFcBboT+mX4Der4kz30RAIjl2JmFFbI
pqlnC6O0WQys3fCF4X2hSzUOleNsVThVtyCiyY9lS5OHO4BVRfFyIllhfkIs
OR4yUYh/9IiZD8zd8OC9DtS61lRGdgmDCa/GpmCaPbSV3AyJTsAGJjXbpttP
KlwgbJN6wY5t0B+ilXIHUwrZ2wuXFVz8R5OqGAh8EENh8Scb+/AITfvoU5ya
itDBvt8653jqFAlFVs8VMUNPz52N32cWo5vK/Zq7oTiZLc4fdnG+EwGnRXzd
xl7fIKSVMsMZgtjeDRiqpK1z0nSKxcinNcIExSMmOqx2mb/a9kxSI2A7cAs7
plGARREf83uupjufc/YlrF/+TQnbUyWR2V/pzId0QJcMKgb1IfhGxn4cAghj
ZH/0zoHtguXHtmRWlwNFk8+R2ZF0w2FJoC4UewT6cr6O9U5pILxEJw9i0Wf5
FzFhVRqrKBfdJpUZodlB8VhKxucknNyLai6IgxUY9IZ5ccS/iAFwO+c7yoL7
478noH6JBd4cyUVvHi0z2T89hT5Jkaedya06lfmRXjYvKJpG4PJ001ub4XQH
kUSQOLRC0SA02LzE0X6TFm2y06hjNqDWMlWTGeUr1RlMj+sFjUe0JYntBnjQ
hKnLa56q2wPJDtvJRbAnqCI20qC2tHUngTdUDchsjpW14UIJCCYQWKnUMZEV
7e7YYwJpPcWoVB+O2FHzfjdkIcC/7PlDXPPjfBemaYzZKUGHGQYKi3d+0m+S
2CHtJBRtCLEq185LVF/zszJ5kMjMHdzjoXNa2tFRYvbt/DeC7iSRwR6NtJ/F
qus2+ryGf7ju9GYMfIfLZT662VBxx0xmXV5rWn0duxsGNaG/Ba/NmMjI1Mk7
v2axR/8Nwc62+WWipzOJL7UIDSGqpFsIbvw/rcrrsR/2iGss81awXfRAm/hF
p0JYBc84GlS70I9S6fAdlJ4yzmSpEvgU0DDM8VRQavYBPEz+LF+Ho9wBrhO6
DMvMYBISP23VqHSw0P1C0uE7dYBD6eySCTqcGbiyqlq5A/VzYKAjXaQtDTCM
S7mAcZcnG5bZJO9pef4rslibCeWxdzCwqwdFnsQyP7E6IWbpGpMRcKJAwikK
3/oTTnim/5oTX6sMP95xPRsyVJr7SYcus8CvKOTKTtF33pZIcgGL0TS/ql1K
wt7D8qxCzL2+2v5BlncNJMQYnOl6ga+UyXlqWN13z0CoT+JzvDsoazwy9o9M
QurgKuaC9PX4Vy388oZHxaEaSDlEBBJgnETE4Ta5sSjv2W5GtBPEeJ5KGgZt
HdO2ui4XG4l/fwtslbSIu4yb1qubJw9zqgjocOCwYD3SBdZANsUSPt+X/9q0
36w6SpElgNQqcJM70n4I6+vaTU5gPwuHOB9A0iZPrKVxSBW5hxuj6tjRbE7b
hZLAJDSAeRoiKmOremRnsAx2s9dZSVxXCBLvhzveAt7jUNdkiafqoxZbd6gB
6J5r9uAtgrGtosXs8lQ++PQLJGaKnyRUg2OpT3BvupxC0BxEFvZFjq1Pvk0Z
ruJ5tIQ+h0mabEGo1ZnIZb0VBbNsgQQLRBubJG05LUoaUrgVFPGZ23DVS1nn
DBdhZ52Erm1Lzz+Ztn5odVpvOUO798cx54vWsp/33gfc1a4MyEshpzX2dBUc
BZxU+YMHqwShFyBN/wA0nFleA8+j2hgsHnssWlsaeBSe7JZ5+i9Oc9eSP6Ce
U6kommuYHOIYo2/lLFFejGGBenFaPIuP9V20Zp0alvkX8adjzk4Ydg2TaXl+
Jpb4O7FHztt3x5SQ1a5Oz449glWujRsGCLLKS4Wuaw30e33edBtCghU0+Wch
PkcUCCYEJp6BRKJGXduCJ/W3qK6jCD/4g7eL0SomUmxCivsUV5jRnqrWvrH/
3EgRE+/gWTRbkwPI4uBXCNRLNb9e0YuyzIZmMWxn9rcxvziJPUAk9/PnZ8Lu
qO9eSbHXU1nElsTk0ETHSRE9ya9InMGSn0iXVj8WIG69xSYL1g+rSj0guHLw
14TojTqSEaxF+971YTtnAWQnAhUxwxyauDCi0f/+GGUPdwrqfDKBi7Ax0nyH
G5iSCznWMVV/OdGJbtaat6nAJYPXuYFQs4TZqYQqhE8W19XUiUJmfE1EwCM+
8PDXjZIWySgrXI1MbkvKKuzPSC1wpXmAneHp+xISgonjzuernB4N9L5FDfwX
a7CJIXECQ3+O6CYvSAiWyjh1iEfn2PxxnZr644unzkcYnZkHc5Gvn0o36TkE
1//Yw7Kmu0Ww2AEcRCMvwaXDtLOQHaehWzBFHM7xzdH7oxM/R7T6f2ckB1Iu
cDxDaowMOkltvMEXnzLmXRVg2Gw8Wd5grI7ABiFxFvrkbfInUwjW0qeWbHQf
qEM7w+mqG3a2YKIW+X9vr7smlZVckVH0IdlHsiXlp8zYm/cqaMwuTPexQ5Tk
gShVr955QruSixLInl5HucmuPajasPQhneLn0yH36QYv+sLe/HFikBTT7c//
4BWFUWPRfwx34+J7FoeeFgYS9SnoEPmyQLWyqFI+s+9aZr+NcCcr8fgIZtYZ
8FS14wJAcPytz8gluKruEwK9kPiBHbobnhWcPfZ33Npz+qMHwP2tV8hHGQKJ
uHwKmnOrN8sh4QtMOXPaxMWv6jte4bgG8N6o5tj7VOTZH5ciuW45+yeVRX3v
YRMW8ox5b8WU/Erlmd/9EzEs8WHda9aG8ItPKot0p6Hb1Mzkde5dzuDCunox
4WHHOSWmftBaSOeBx6sV0xpuA5+zZuhTo1hWxOZMOVnJT92ptopbj22PGYw1
gHp9vQmc08k6KFZ50gIULgeiS+jtyZyeOnrzehh4Hm2AVvuERA/fj1Qf8hUx
sfX4BN2148Z3aQQ3kYrtX7F6NwnvZGNE+tNt7Q/6pXSGHyNfS18SnZEC8H68
tX0yQqm255jsWmqjONe1xCbkD4JF6fgb/gFW1pnfYJmzJ7mFacQhCHPm09/Y
PlinQGhOXmp2/lXPMv4NG2tbsSyPmmdTShM4wS4MIvTjNSbwAs3Ryi9Gj/RB
NCf9PrjIX5qurzmic6wWjVeqvUDqrLrth5bPSU0sz5s1ZvioBZbEP2bRWMX9
Z8zGUmjkzl1aPk7nuhsK/wyBGipVUNRLmvgifYeiciQOwi+QQLdba30PBsTd
sXNSf7XWO0uRiOsU+WJuXfGbXADES/FnzPXKGIJZsMX7k6E77Nm+kTeAbTAt
lI1nXvDxpa3Tb+C9ZtUY9v3mrXvf5kE3Z4z1dwYo9bgwT+Z0rHvYVGTuibFf
f/AqC+qAjUWvi7J4b5OgAgP9Yzt986TmqcQKPy6OlssOmKAM7EMxajfZOKOV
AfGW6vueIWmrICxsSeOFP8adNmbHlTvj2d8mcT8S4kcy/7t3mge6ZIt65ufQ
3PGbwInJVHsqCU6GltyuCBvoLUgtYAER6t3+P0zx1lPpZh0FkRgn7FyyrP77
kBOXWV8Amln525XjC/c0qleJokaAqKsPUTsT3iAKxW/8QSTaJgGHbzrB3oPg
Qmi+1NRBFXNM9yWy3VkGLcBX2dJwWh5dTK2rOo63qcP+Fh//pDoDvWkr8T3v
eWWyHwR2khVDUmYy1CzZobN4G2mnheCf7YsziiFGc52/iBDB9tk3qGs0xorp
PR2MPJ9zp46Tu/f2fR4pKIfOLBykvkoo27gsV1NEMQf2ZgReuuTD+li0IhAR
Hgzl+7C5QR1mD1r5ukiFBBxCuUG7Bz/6DvEUUF7qYKoEMveu1LNKNE6MSwbo
bvPRBYoWv62uF77W71ccMsKuga6VHJ6w+1CUrdwNlPLxel+sjjrue1BePfbx
pCeCunw2dRr8Uoy68M4Fxic51xWFGs5oReapaJd18+bQbgfke32c8aGtVdR5
vU3kaf5pGBqaqEYCQDaFXN0KI+0CHSIE6E9xVuIoOHIFgRuOB4hgxWG/7taQ
djWQkT69Z9Tl+YMGSQsAQwFd3O2jPdunGZSxGzGQwnP50sDquvDDIKqTC0hh
8p6gQKhhdYS8uroXZ5RYrynUcv0WJh8JUjG+qP7sJnPVpRIimMFeN41iOq9v
Cn8jWLO24CZvkBHBhcUeDvPp1pMgVDZLTgj4XEMct3EESST4qCTcevAX7HlV
wZkwrvipla4OWcZSKB7zZ+KRtNIyVAFprpVLMZJkDS3Jemao0tc3UFFpqKKd
icOhiSJhrnlWLm5ivyBrwbPkJAvRVyAfbaqGfl1ZNftmeeabiAEVeWuva3Cw
01n/GqUZx17rOhtZvhziPu+9Vy27sADFN3wKCqbh7mC2q+y6L9FD1eMBO8I0
3uKBkn2tlOsud1KGRsnHkz2PvqPMywyWCVBuXMFyOMyrJDPWvt7kwUlyDDHR
x4mpI33VG2o+71JdeTloYHMEzti+cMKTqD0iWfMRctVcRdB9xCfjfpBxxgHi
xrnw3U44LQ2gw02aKYYquWfAj1zvzkP3lMy2P4z3rUBe7t2u68gkNXREj5Ra
rKYQrIVGzXe03hBhZUg9Zf0RrPmfkVfkzRAXBlsRWRH76oRcpMpARjOQbKLb
bgON8z+YNz5JBwnFc8MpIY4vcAsQRYewZNsnLZzQU8aucCW3G1Npd6m4O4Yj
BPCYR1BR2ifQqa2f/ZoHr/DVP/iqezbQAIMoiOsAaDc3Y5B7d+hRV03C7UF5
EQxikG042QZn/c4ejbArleFfxULOZVmVczw6zdp7+Yca49Z0IfnXdNTNT5T6
3dJ9fSxWr3Ji/uPtkF1FRuRXWN2I9cle9v6aEyqj8pt8YLd/XZPU11aH7Fxt
WceULZuHKdJ5y66ki0L5YyDiG8ZAFJQoGDJQ209ZIzYA7cPSQytWx7J2/pXK
XggxLAuwkG2QAcBKzDY279+WzKW+3GM7620mme3K1Din9SYDoYpfnKxdqIZC
QvrV1JIQymsRNywA/OFTFYxjRU2tnyTQKIAxx+Vvr/Bz4gPYD6Yf8cZF9/zr
s9fi/7Px4e/iOOriQ4EFeAFC3iHlfPWgtZLc113vavGQKi7eVAfJ5E4DE8jM
+kn4yeEXMFwq6p/n3IoXTDinqQrIeAS9T1J+Pep+GU9VvsarsIBZRqXK73KM
yY1SCOMTjMxgqB+hNsiexWdnU1MGxN4/BXTv+Xsup97TsZb6KOQ9J+yEsD/z
GvLv6qcHYfQKR21LdmNQsp06i7XbsnvCOGT4Fhw1PLTON9mvTVBQiSzDRaAI
HlroJVpUMxBUea/pgXKFBTjNl2+bbg2HDGDdBKeVHHaSHORXUp8eIqssBcdn
p7Ss48bq1S3uyM19dA3AjmW+NyKT2gM0YJ9SvtpjhsJFa+t8VNSOTdWKpNu9
bxpXqkoW79UTaQczEbqYZ8zFeAw4y3gCzBYtK2LkLQACw3sl4wunLFwSN53u
JaDbd17cwEdpDFKlWiVj0VtGKVmAQ0sFsdZYnRZEcs5/nlcmUNe6jOdqBeSk
2qQw2KTyjR16HPk5mxMa2upQhKrsknMzJjVZDMU9nchT98Vqf7vQXgAHnZH3
1ATY1yD31R1EsqQbxRvHi1vo5e9wk4J0dGrlW+RhW7zp7eWmCWVWBCx1L3Gy
NmyWrDxhTWoo20i6uBsMaG3MQ28hIP+1ECQJ7VcoJ9f7FnI5+pi1Rfqafa4e
QOqECg1uC/SDdxvEqTh5NSAO1zJtH2W9T3NlzvyDPAzQq0GuR/viElUtd6pp
DcKZ9ArJKfLR21+JaPDC/0aAQG/KXXlGGg508hEUdKNGhGXeqO+t1IPVudhW
hBgEJ96cNxqXmTqa65+ZyWVQH6ggu/3AB/7Jj0nHwjZ+hmwWgd4LFL0zyPf9
KYjfSqxVtcSEuBC0s78vds0uk5CrscMGZSHoYzoZuNeha04HG14BUqbzqCp0
le7UQTtrZSZ+P6omTEX4pQuqJt1ttJu5JyKeTlds41rNkM0o2am12/vhXCuP
4aPfKYbXhTjt8HS+dDW5qXW6MQFku9GpnfQ0LaGHB03xhrDaqJ5tgt7ZShid
8sHfJPIszLTgy0TdOksVfVvnMfgOY84HJJ1ecliuRTyiPuOUQg+YxUBkF7Ed
ZJUYK2YGCyzdgbmwj2kkoxb8sbP6u/WwVQDodZXfYgEC5woo6vZuMp3hPU1N
MRuwoi4WFza6Mc65MqhLe5iNY9pvfj9F3U8qB4JGCDzvdFOYwt+Yb8YI1CYR
SYtFnE61bYOEv0lSqY6whsTvczOB0Y+I1U4vXJOS2iOC488oTyQYXloHCJua
pwZ8pBMPDLLJKvxxlE9gALklwBh2mvdoBlAu2SstJWnxqDlj+rOy8cHXxxWm
ZgwXZaLXw6Lh0dGKSQlbhPoQFbdd0Maqy9y+galreyJqVpbqkbx8YanPLtzl
P/u5IHPnym48sLYiTxhcT33uGxMfk6TwjjQcyY8Uo0vb41f4OtkH971vFCUs
2kQVI7+9DI9aPTpE/uex5C1PtAPEreUNYFuL8deUw4aejVpBKsjNnUEKktX6
TZTpl5ajDeHxjVK4pJRJYQrngXYPzJRjtlS0BlQADe9iYP+hBTLrFfvLXoPA
6KVmucJ/LeIFKOihcFCDYOndQ5zI3u52jSWfCF/y/Cum2FSVBEq3qY6W18id
ESS7+ZGtsBswNMLNy4GX01UawMNM+GPEey+XpFzpcSoXy8N0k7om/LyoLNZY
iGs24BhJWndVwNzbRPUvqZUiFLFkg2hoCRxOGnLa8CTktr1PTJuuPtqMccHc
YoPE8JJq3gbj5HympbbQUm4VblIVPg7oYT7d1+O8CN3QbWn6wXC2Txb098oD
0f5972kkkRh9B4+A8sYu9zydQnozi5tascZZczRRUu9/Ez1D/mkzX4mNHJyH
+3Wc3Z7ANgeOzWNdnmtzp1BMxZKUQO+SBFKaXjewlXzHVrCY2fzOTwQiNoEB
cNW1nzCQkRDdvj6CHPOWbHi9HrXTvxZh8cFvZSDEfpiHd6RX5OI9G84PbF6c
PdnOKZkFdnr8b1oWPLmofPFYAo/m8VGolulGheRBWht8ZyFWnt+EWdB6Lf/0
0bBUp0or0mxonnJ7c701COgbENY45xO2xEBZEa3lchlxnOuXPzEkTC7/vKuU
uSp+oCgOG0SnTjxxZaNvIQiwMFFQYTZyLxTF8tckkRu5QY9rix+fntqEKnFr
TBiTgedrXY5tQN+5gz+Ck0x7Ni1tMefE4kNjgN1UCOpgm7Tds3wDptWte8Bf
yu1eHSqoKTwBSE1CeaEL53HTNV7rs9Tct2oTVkcwbL+lw8GywYQkAH0odvCt
HYu5kzFLXR5GvWyIbagk2q5Y6Pm9vM3aofI7hknYY3lJu/BeRF5exZiJqkVl
BAlTfVqv+cL/J+KHPjtdkCld+8E3RmAR1ElBMFggagJ45yuzpl1dJXwsdlli
40JpCb/Nqt1gqnHzfk06TdzNVqCQC/w5FX+45rTt4VCJTxrD+7XntnbOJAr0
fEQkuBBl35vdqGyo3NDLVLUspPFy0dNpRtPhdNFARWQRU/wOeRB8o8IkzciP
EgoDkLKYdJz4m3ysJiCnmlnuJhnODKR+NCKSUvoO973Brr6KqHOFCX3JwBp9
Ir3grorX8QMqaL4/zEx5zzX5oeS0nHTs+pqEdrfhH1mjc9qbGvk5CY0dRTUR
yjYXYfW2gaUYvLWQt78MtLOwZ2Vdwbeorw/7Mk5JqxKSuPJbHmkqTzEE1pLx
QmeUfuaiwS0A4d+4+6oFndwqUop574yA2ur6lv62GBAzKSu6uv09IAOzrRU5
FJjl3bVYCPYd/bwc5/VRAw7jY5rAxQiA9+nGZsEtsOGoaPao2sGR7CkoUnol
R5Q+BNqqBA9547nqGfgpFYYf3RUvQJmZgYs7LZA20GqLphh0q0cAOQmysahC
fQAlRXxZbXLJzEdKHDzL2AuEApTUc4QTA6XOxFZ8omMFdme5SS9xq+joDSDg
qYtwmsEMONXAOLidbpnpMrl8SadMG1BkarEDC/Cgomijv8Cn1xNyIFRAtEIX
zUMRSYZLdU3XPhXrDEEYugHpNCNC1jwfbqOarzlIwf8dm2mPXReqnHhw8dNy
tStagLEzm2+KoecTb+je7ZU2kfAY1BHi5XQwk5dfqEJJRRlS+5WcxLdGy7wy
gz7QTZE36rpZzr+2vV8TOGv40KplwUuezrb8vL+K5xOQgGMY7vkhBYjEADJn
7S5hohcMzsakoXm1wyab9I8bS4FjiBhgNSYnbqLjjtVDgax27kak3zD50W9D
J8F+MW6nW4RbcKN7BWfkNmUeDzjSvyTBGmOWI4KrG4MOvQg5IIOrDdHhrMIv
EHlzcL0FTx1ciXVKYsQdtTNMHp5PVHuqTu9L+kGplj2CRcEKCvsdQpQf23QH
F268YgWpHs3BIehnc0N7+uOaYpwYYlWKt5nEoyXh8pea61SjJozf4jAjvh2f
Ellen2jY9/eVqD4/KOLCC0SGclqe6ACGy5Pc6V4nLiVPzZrC3VzqFqz+8tXh
bAtLTVFAyGQbZ8zZayatBcrWNJKiB+NTDVYPHMnJjX8TU2WQsa+O2qnd6GeV
1CFK5IfQfda0VYe6876givywFJvjc/w5mWF2b5iBKVa5FxH82isB6UBqucL0
FX7X9dT47TUMNen4PHygG/BjZtApqXxdUI8mal8ODJcDg6rSEQyESil7iZbf
zhoRjdCTgV9T3WsFBMyVjuHUSSL0YzRFr86FjzLE6vFm+/cJvcQba+fSGmFz
XnhNzjgaVlnP33PdlfnT78BI1soYVlOGiZuczPPNw0QMgXKTZToVIsRKk0ez
2U0r8BJOKINSirnpTkhaVzXJmTptFYgdBFZIb19eIXYFtOfY/QnKFyKYnPOB
qHHH0FVP464N8jq1G3ZZABPVPXdFe68bQAGiW/JHE3Ue5/G4iETV1K+d6Dpp
zsMsCqbwi3a7yS/6XK6QqDmb6bqzGY8b5wQDYki0YqbH2zS/qYR4cboiJ/lv
dNjZvkRp3NvlVlrq0lbFgNrdBGURCH0GmPPy2jae5Co4kMg3KU72qw9swKnZ
fv8Vp5zPaPpdQet8jkHZo+Zxih28CfE1iB+Fe6JmSJmXgiEmtlxutuvHz7zQ
egHbov8655BWlRBkzxgU/oa6R+MKzP8CFMxJWUAPPrjLSrxkfbVwqrR65+N5
1MShiXbSRwgrr4yfraczSJvnl8N3R3PAmsppFEXYaviaKxecj8uBcKBewZJH
YmmkFSJkfjoOaTAoncvzoP/xCNaFyeormj6ucfcaqkFlo6rYR46FTgiWOXrU
U8qCh2NsuW1JaR0YBfa2ETc3Qi9GxzGRn0Dxi0LQzbXSZ8mqwAidQTD17z1/
0RGTQlaDlIr5WugN9OGdsM39q2/f8CKSIpIiTNt4L/GmvdYp2u/KYUWrr/8u
hF7W7kPddHRZmjVkIuiGCDdp+aoVRho3D+10mFutSrDd1iM3r2IBR12MmI43
5dssOhFEzwDoEE0+4MeAzxoLxJ1skAZGQnbyvmv4F+qq7c8PDlWEtHLgPiOb
PGqDkr5fWkoF+Ht9sFeBdSk7XED26oCqxt29xTBoznDJNyr2k2XDDv1+YXkx
MWSqtpJ4Rvjxpzs8JHea6TQGMC7daqV7ZEQbzVtUrXZ4yzpuYvFB14cNidBi
BCtSf1ozZqv6XLTTCwQtEz4LxZ24MLatmOjElLE3rm4j1WCn1QvMLqMsoyNm
P+Zqytvw2K1LZnkmRFktWB0l4LOX1gbrM6gr2zg9P0ultzSKLyqHvZ8BtyRB
M7hK50aXkyGTkHTx/ArML0pLqphLTJUZzVVRFp+FTFkiabCc/XKqkEsTGsSb
1937MPmsaYdcItefLy3y7eQTqc1Xc34c5VG3En49MA92+Em+/+XE5DaURg/I
R+/Uk8uI4g25Fg6fZZZCvgKZDoQNoDFsfLtmbh4b4PdwWr834+3vRlJgTGML
PKEB4nryuOU8OTShoq9hIIbycyCnFEUilFR2JU0jMYSAk9y3nNStqlO3qCnh
3BEnePZ6yxFFcCKsoXWYYBQtS08RQJe3dC2nM1gv4oXY8lCBWLZhZGY66bcr
ipNJaWeU+3JNnaK13MbTA1pUsMwWJVBhvxiotEbkH5aakR8OGohYeXoY/yNE
rQh2gB+/dKHq8vQ10NE1TDwyZNFOJxGuw4ZJCxHvSMpsxdWR+8zAo4t2xf12
0yZBrTpthjTVQbRQOeerrlj2dPmA9FnV8ziWiFBkYBWxl9tjmVdRc62QDtES
cj2HVNIx/HpqehS6uEl1d0Uwbe/4wV0gREx/1TzkidZQ+xTs8/IQofJIl214
XM/EVEI7n9AWKbl5x+5LMJVOmIy9962yyrSMpLyvTNqBJ6caPuMgW0hvez+Z
E9TODLemAvXg/ZQjbZ40EShz7YcHauOs0EEE9gVy4UInQAJQ9Qngfq8L2ABh
ef0u5xSng/x+jy+iqRmXuow2W5X3gEJDrkoM1zZBps6zdyL7ussSYCo9Lmnv
RjfdvXC0GB/qKedOMQpxAeGwulhVeA0cqG8XA61nVWrunlOzkAimHdVIaSnC
jTgik/Aq9VrGD3bbO4jZdMqhRPBME7A0KsSsaqliUciLqJKlt0kC2awT0Twb
QQ2ImYnAO8RpgV3TC8KYybJS0VURj9pME6lgi8kACrJGGsPOK9q8+bEavAa0
Sfl5olv3M1nXvazHapG6zxCYsMVWbvlbRGSJRH4c7GMTIqImkJv5qxL3+z79
UQ/O1jgqqGuNwUvAb/PI8vKxYCme3pYO0A42WJ09Sd65NUwwJtfbZCq/WFPl
XD0QqtPKOMzprhcnGgPoEKuUBedsP2vuMkXmIQAKRkziaSZNEol78kKeOvud
SVLIGksbbsA1ztXOJRkxVSJkAT8yNCsaNesI08pnCO7g08nJL0SV1HLDONGB
irzN/l5ekmVv2TOcls6i4eMtfEimS/llGIW9UrqQ5qR041JiLrTBxfLN+ACW
frYK8KXFafUdLqnJHEk3MYu54qjyRmhSa3kPFg9zg52Srum+bGdC1PbfGyf8
ho5T0aT4lrfxoe1+aP7TxwvSBQSSnDrdVa2ImIXILoeuqQmYxCxwLOL0equH
SzK0rLqs+KGHmjZ3pFQfuOAXBMsuA3yAoA9Y7EumZvd/PutrRVR01qTVWtCr
xktHZ+JzEruDSoLBHuXCCmS5UXgADwx8MxC0O0fF232L08UdGIgTIP/4ReKz
pINtAi0cfkczRF3pzYKqEOAOsJ1AD2yV3EkX7pRU/sH+FtZh7oEXgq7LRGDg
iB9qZdqjP+2ilXGvtNzQDwNafbMyDMzB/5YaK+McoNa9Ovh1dpJJmmdBBDle
t4Ws1nRs7+u8NFIGgi+DDV1sPPQcNzv8hDVmmGBYOMTkRC42ECHaqiKCQN6S
4p36iF061YUPq1ub/VtLcZ6e

`pragma protect end_protected
