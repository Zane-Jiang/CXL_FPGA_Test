// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
aInOFsuvMkuP0EeS32/oMlQWbXWRAb6YWkqHQ//6Rvho3sz7mC0qhQ2TxwZbEOlY
AdSF0Rh4dcZbXM+by2WziWOjdAi/JpaMzlxQHd+etmiA3gp6GiJYnNmJkz7IIksh
HwsSXlHiePPr04ZblLjCzd+BF3XK6BCMWpBNHBZZvRc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22160 )
`pragma protect data_block
TZO9X6XL47+lMVBRI0jqIt4BvRc5Jb81fgf+/pO1Oh2DqxhngKbDLrh5c4PObx0U
IOQ4HY1uEpbqpo7faGUNcv/JMeLB6Lw/Cd5vJr9fxwNDEQoBupR4V728/passQi4
Y1RI4wqiDsYVSIjkUFf5WT2ur7UV6ofatHAiKksYBdoOyq1AMl51GrMCqr8hE/DJ
AAj+6DWKiCGTDRJ5tJlm3cjSf5TrCxDngDBBiHFrqNRObGubYNbnWckRFbJ1WZlo
DeqVjTdsmMNE3r8VWGzJ5tv4jE8Ma2rsrMga34zIK/L9xKy9OfxRb7px3q1VbYus
uUwwPpS07kQRzeTOm0moUXQj82iLQ27TEjIuIfQdl80q6GIkbCAmG/rikNFwiIjp
2uO368oxztjNIb/SFgR7EQsuKiNpPgOrKj2i2RJhkZNIbCvCsSMZXcTVW0YsGhrl
qWXRLDK56bQSvTLyy8/zuNjjgbQ4LfRMKXvTHA6hLs6judyxlHONqHM9DHj+/QD8
4KkJJFDx0FqvmX9XLuK+Qa2wRhVvX9QM1H5hGxKxkcjvIzINZKhKMHHHzCXEn+b2
NFqWJqx3rdhhHverEs4uwQBY1KpTZzZuFoniIowSmnY54AZw/jcsGjynIt5fDmlw
N8eBFVjU639AgUa0ERbv6ZPOIJLBvZseRcQWk6srGcdo89sfCdKBLmnBxH6dsnRa
wI/UI3Hwp2tqIE2u11SOR1RtAkLM7gLQCdOsoLPLQnej9kB3p75U1uyCOwjUOFpI
cHJdX8EzyiFdg/5SWOEx4MTcFcMeP1lLVIFDbvY38F4lgx27zVUEWXhUQ43nfGQA
H61DMcbjDK6MBS5lO/R2MI5Dj8lCQ3C6eGDjGCE9ziywNeseZJWy9IV+mC4Lpv5H
Z/hKruAbOmRRr6IXawN503z5V3bT42dww0T7Tq3nETsMONbsjKXuKaMqPs22msdJ
qgnAiMWWts64Dwo5afTyC59CJlJEM6f/mBdCfGxVnKxomrHpWziiopsH8kaQK8jr
yN0s+utX+Iff0QnGmAbq9qSZj3L0db/cngTo/tcKUd8whsmZd5CeL4JN7nFO1rrx
Ls7Wt0+Wy8C7AS7I3cSul/xCHv/bUtkD1S+DNarXpaCqd2zJYq1eSVNrGzgoF1pR
ItjCfnmDOtur0gYKq0tYcOa1kMD7tZES5Xf5exf1kMEtrC8L613QkxAVRUW5dATK
pD6xSiCD/g5+8Gf8dsFOl0UrdCEc7DN5d8bI0hNzhHfh2JdedcpdelCCFjqvG6JL
5PFILJ23qvm4NyJUvT/HMfVG5kTI2sKbbg6gxHVcDxdtoSeBS5zbjlrnA8KqpWeR
y4sPpg01OWpVquCxb7/jzn/dQ4BiAnKw0yZI7obgPH3p3kPr/uUAzrchwLoxae11
rNwe8aJjwEIaf1QKnBH0qX2Oj1Z8sCgfujf4jP1r22BBH5/waXhjq7nQOE0MYcin
i4PAsTDFBon7FX1m10ty/AFPXbUEc+2pOE+YaTZ3NVZv1GGQo63qenRiwgzcvXtD
6j6cZLDBLvicRfO5N3+uBHhH0s2EJsEgzxhlGCEE0sUHxpyWrD78CfHl18j62Do3
I8juubn+Xju9lYtt2uStXE6ri2LubPwjK+xGkgSovk3AMaa5rQca9KlfNpfj/+J6
G/HzWtOIEp3P0vjDer5gPoOMuEl+UNIqGtEbQ40pPaewLlvCZav4onWmvWbHR+aO
LQdMjoJ/kEd3TlVZlxFZPNO77GfjD7aeDo1161UmQvIPcqUbMiILXPn6cR8tVALs
L+NtNQVnCwEm2DP56hmh5GMrzEhhExUT9fw6EuikXV2aGiLzLEFGufSiem2iuayO
6SlLaNXj6X3HLBYKU/8XR+QXVzV2/bnbu77IjiGaffEah2w5a5L9rnJUu3ia10Qn
RqJyhE3JI7HNU7GkRah5VP2doF6swepUffDmDLsy5JbKGppdmK7+8yKHzAeaGPgr
bDZLpOAof2w4miwymKqZzoomU4dXGdAXZnb2gBkZF8T6CkH/skxuyZj4ICmqWjlP
1/p2NpYWFHjNTgs6x9rMqh6hxws39l01GDil3mYbwKeG9QhvdFDr4tBHPtUbNl5+
/KHT4A82SP9iY5i8fHfTWQUhwiZ7LvMhOYmiJFuPWTrW5im4f/T9yft8D55XXnWT
pt+f2DdYEeNcZL09puANpFdN1lor/4stJxOlzNskFThKHJuvFH8J3v1xusVAWfIp
U7hnejM2kgUbKaY9+e19CNBHoRb866ieHS2FVS2Gsk3ZXdciP1q5q+8VlarjLEc6
Be1Ma2A8/m6EOBYLy0QXohbcvUfXvdMIjLKkkMgYWtfNMCM6H18iIZO7J53FsvJG
f0FWGJuPy06PRMwUxq9nXSV1f9++xbDcvoWd/0EDPeuBWytwFb/2JS+4HpLfvHZZ
1RQIoH/HBUgePtu2NjZP3H5No+71kMex+7TNL2surNSDAqFocraVKvxBNUpPMUR8
76RbGxKd0/RSxcnBUSZZNwEQLI3Ms3vKJbOR9NyLq+gOlYziWWxOnjQSEEK4xT2T
ot4zwH8ESnT8pvrX+X1j4MXdSOSFitbLeS/WoLDec/PuXKFuWuapxv+qnYSHPmaN
sdaQL4IcpvXnLMwndsQGjkECejWqoQP1cgOvAJl499sKCzCA/gbKJ+1x3x0XcMUY
MkdoGP80VW0Mh3aU+RHkDsR3uoRxuWd3Z9f10KM8cdE1EagsmsaMd8A1CC6Dh4lq
tHkPJg0r2RSh0V2C2bcW993J8AerZPTNRv4AZXR4AOE0pN3DJc18sgsJMfIw+C7E
qfnJT9WPZ82YWSJJkhpTHqbTt5BG0Tu1cn3cjdD+4BDky2Ym4Kyu8h5H3Ruyj/Vd
FsMrSzjlVTGLnf160rS7yktLGHmIRyVqHNq3Jt1mk788kTVg51e3JYxY4y1v94Sp
r84s8xQLnAaZOZF4h0E+P01p9V3LRwq7KeRYDVbZ3Wf/3YPSX2XpQKyQEH7hCnQK
nQ/nLTF4aa1ixZjFiCaj+wCAIsXjikUmkJfTEZT7LZl0DIhgB4qrjbACBLmZ9Jh7
OlphZjBWCRbKjX6XFfVp8hi+A/FLA4C4vbRA/60GfZGU9pgFiGb/jt+JnU9w/9Rt
8RspXhNJt1SRlJirhDWKJ47ueDx9GhYA3DnfIkCyZJu3sW5+qex+4Aza/B5RQ/pw
E1/UvyKiXl3HkAWkOhvnGx2Uv8PcFWT1bBYMPnBZf3WesQy/uf7qrLl0Ode3/GHh
6zxdzxpjsYQ3bnvSdVLnJMRF8lVESQ55RvotdsNTwol+KrcI23P6u9ka5uUdDxgh
6a8flGVGAC7R9OykvogQAg1qmGIL1XVsgERziPdk1YCBmNFiVrstgnfHRvvLjNiR
V8Iu7HqImN8D9PhfRsnrNkFE1ALsvdcQUQ3qIle6nxNU69IaMq9RvgyLE44uzc28
0KTGb20K1mUGDGVZgabgGiT8xkJ6mbPVEK1yrffuk8tLxPNgNEHPP5JCZ8Whjwzg
CLavuUMOLbktgZpRyYtVxcXWnF56qH6kAVHCAD2SZuDGqVS3CgiJTWBYl23WHeDo
/ZvrwVR2XmtDibMnlZFc8UMsZu4ed95dZDKzZhh6z/0SFSRq49v7szOmkX4OkLLX
wWTkiR1pZtzOM/6u+kmUQg95RLqqGXMjbjAeGq5gCUMjHkBotpGCo8ENYR5tPz7o
dHZupsyHFHbNDm7RjNr5ShKIqUzyiXCUVHW/sb+SJS+4L9VeifHHEoYJckXej29m
paBs7cl/rsuI5X2z62MI0fI5OS9j+I/fB4zEGj2MMDImoeT+eDqw19dz/dswTVNn
CeNJl9pvXKX3WSZTCtSpKU3nB4qfvQkRtakcYvy8hC7g/AXOx2IuU+fw9P1eps3b
tRm02NJcgOxDHmrrYijOt7VxvAb4o7hjFaWGHoqDHQAC1CVXXzCyJ4bSqNDeFt+Q
9BWaextd9Rldo81dmMH01wfFi6pqzweC2+uEgAVJGM5NIhP6Kzd2rFyedYmJOl8q
0ldWuJGupJXkefuxoSZNHOJfgR/ij7sETkd/Qpt3CqbzESkRVUPi8+HXnBMGVF9t
8KJAgomZHFA3UhRME4F9m7PFqWvR/bZVJK1ozk0F3Uvx3Q/WvVjfsqVDi/i+vKQC
yG/1rdqkN+C8Oa7jPA49YLzxJtw3SlhnUxalrQasvw2DGEC2i0BhaavkQ//c9z26
P4h9GSXY60qzpYH2uSXMjiLBNR2wbQVT99i8Pqm59NmBz5Xxf6A+PxhKK+6HUFyM
MdIOajSB3tqNbj5/SPVg0o6IgltmWhkklFPXD290+omWAYvERt3vqL40lmAwhPTV
gI3QtqFbFDODLsWBa62E3hR1MqEgrCeI/oHWIiMcJYQtufnuz/k1L2r6jmxpfXSG
ast8VIATTX3Fio5taDc8mJnN6zh5ajBg1m0jTXXE8F3EfZMS/6CrUCVDl0/21M2b
xZo1aOyrkPIvupzFOWjCgL3KTmWpd8Pgwq52mYoSjCaaWXoRrNWR5amZrojFFRnc
gv0Ra0hrlaWLO7tS7KibG7ruPL7B05m2Ef+m3eczKZdY69mZYVN6fatRzfx0KJFO
aZ6fPhMN+mP7eDIdDR5LAuc61gkq/fKR9OMVo8fLAk6qhD2M1GsFO1CIQWMma3n4
vDO+CSEoHNtqYKM5eqnrNcYKy+HTZBjWI4Z3h+rbXBxcnoBTE+8JBsZF5Tzrv1AM
9fwQub4uD8sdEs8SBrmTGr1y0xh0FW0ZPMIXkcnxlzY9D7kei7qnNiX6T+fQS8MJ
kRq+6H2x1xoOwxQp70+fP6QSAcPBRz9cI5KgOeEV+/5FxEEohXqAyJ++paQkE/E8
d7cukTlcVEAy+niPpCw9TX9qXzqrLtJrtTeY5zslxwKz2mQm6KJZOmS3UT3RPwPB
kfutO4Nk0f2/ZBaZkVh2788SkjXUo/vWNo4jubkx/rH8ixMUhnGnWMiUneA1oF+9
fn6qLmyyBL0XtRSDEK6U76Jkfp/RG3kcXNLaKHNVDaA1qVwP6EoY61du9pLlBUVP
pBCvsPFDvZJrDcNCm7LpKtpEUnr3S1oYrYbfS/c7ZFHkPuMOLFCYpY68Gr/D3han
jNbakQU7TQg4xL+L03Y/AWUqRxGfGRt5kq4BELsDY7xNe38+J7Ew2cHw/8oemq2q
Q9TjlU/4+j2k+Mm7WsPPKSXbd4gL4IKRakanCkpsnNQnR6ZpzBJOYtZjq8Gip68c
MF6hu1r21WlarcPETGcaZ8vAqX0pmKMyklF5sEwICErgCkN1uBHbQy5hEsVStJTy
oXpS8mB5OQknEu2kWxAjNe72dnv8rMjk7TKeCeGkaWnfpPte8nOIqub+gqBBTNiW
3KHKfTCXyOKuugAG4zvbbkFhImqHRcGggsHo4JWZIwfwO07K0mbvsK/AysvNjI/2
gaAqkubqodUb2N95+C5Y42WGFWljhojDI5MWRBwxq271Q5BNiy4uNQyDDYRsdD2S
LwaLPjlTIxqvV/oObvwI9qYved6p0n7h/qnb96396EhKn5N9Urw8zhVP0ZkV5UTT
yBiIpz1yxvbAAG6jk8HDzdZtAzITZqOJSY9qNbWnrBjoTQos4UvYaGkYoU9b3dvv
wMQAcaf+zX7hAjscds3p8e6bkgS3CtOql04ojokYlz3F9GdRl761G7WrM3MOexZ/
KlBwzep3WZT5C0+MgOLo/nbmB0xrHClwKuEj3JwChVtMJkJUdFh6Sxw5is3dt/xX
fd25UJ6VcG5UfWxgO+gHExdBgrg7xhNhRTh4OCvAaF31Uglcc2KKUch72rmqxaHC
POiI6lbRyegAKS2a6To/ryGfaN7cbtQmu57F4XLjuKa3qzTg3DWuBU8G94sWOWFX
YXgh8/8l9qErSbvZlttlVFzNdziHk763eoJyPodcMJdEmNaDNckqD3768swwOdve
sCG6B2jwt7aSh7p9lObFp/713AjmjtltAIklX/7ZDb1LsjgdRi/cXX4mYR8ZIkvs
S86C0QiMnKiKcHypAEoYvVRM1lbifGnv/XO+ibYciJWzaK7dWgxWf/EcDb4pjGGI
J8HnhunKOdz94c9hy/WifzMwcvARZ8LN3XYn9W4eyFPNCoZjTkqMPHLxUTp4PeBR
Z4aauGhItyHgcptUpnkwIUgUmpjj6KJQsx7G1Kjh6t4WbDOdeOQwjVANyk4rgPer
4fVuXRm5vaPS+O/2sGkKeosKOofTsW6wbBrNq5/c2zoFMoEDwXv01AXcPfoX4rTb
EbVOcIxF6s15mMa6v585uomQ2Mo/Kj3mCoesZaLa1IIlNxpkALqNrKt/OjopUAar
Jg5fHiBQREoJ7im5aZiJIJEWKR6Yvstkj84EcjAJndYlPu45jgrwk5PEmkhrpwx8
h5Ao43D6XSeHJIBimGmOD5FxND/6fiZNiyEgrQcOOTgk3bnCd1qPx+fGo1Lapulb
oIwZnWWGYj3m4paYHLrQootjJyp/lyp+sULyqwWnIbIjmSA/10u4aKh+3MCzPL32
apKaBY3eWU3DKT9LJim4OJnZCYGdq5A1YBeHK0Z1C2o3jBFHrfn13WXZpqJkiM1e
F07ZeJfOYodjW4J14wUFh6vMO4XCZCSQhmNg3YJtuRUjZWrln/GJ13LaaaONZFrh
D7L0bgPHdkAGOm1QDEOYkY0sm+xZKM6Tviua/x0JtTkR3MB9vXPnqz3JzFRZqAuT
7dK80dKJK7LjkrDJW4o77ubQBEV48jmfSGIzfN2kIvkj8MJpQBHBDXQTJB8kyQJ6
MqAUQk3qQYgSUPXeVB1QtCxZTt1WeG3sHLfJYpOSOlyG7y6gwPmpzqqeYeWGonHG
QMrSiQn9n/w5ErdvYVcoBQkXAYAX1xBRJnMkBjyDoNZEetwhQnRqVNHnm0EOD/4v
x/MCgE0SfMpSdGpyjQoR2DdoipSRNhlrSXNRyNKkLhrpM/7AeC72s2/1sJzPIvqJ
KDMcHrXbROwKLlDVBd7hHCIF8LfOrVIQHcfML7yK2LxtYVLvOcpbwFaoyLjpPDvm
rVyY380mUc27Dc2J92pm2B3l76N4EZnT41SAEadOua8YTQBXHVabE8BB3icCF6k0
hHn3tZ20fX/IR3p67ec2wig69GWxwMRewtaYTuo90wF9W6FraynQ6Wr/8wt2OMaL
Izckvah6i4v9juubOroCwCYYZ5f+ZwtK0JgOd+AqVqfC2jFPvBPxNdKl5gWMei3G
ILq0gh16Cw95pTqArxfohWYA9c6IcUgCiXjXXqwa/TVqd6UXhGm97357IlZcvGDC
ELNC4GDNJkJeKaV9NjM6ZtlxgrZvxTv5XDmUgs6c7fI7l6dlvYm3uXYEH+mrJYKm
LUUu/K/xWi76t4iHRB3lAsBF34tJXM8PyVMnb5egqDTuTQ1A+Mf8QGQBtNUY3wew
B6XH++EQuQLK2UZxnwoUI4erDmsZ3PcL9SX0kDv3lF2/pJ8po7r8nzpsXlSox2fQ
L1IY8V5q/1s5cBvXw/4anZPbDi0T86eCleziIjafdHfrtRpAzm/WjHRbT6m4XykZ
mmFCfX2U4mgBRYoV99v7lJQKcK7K9rwPbuov0HsuLOINuyRoQGxg5Y+cNxBuj8Ed
TlX/33qYmpwpB2OxEXkqhxMpwto9CVdG9fQWEVfR9/iIp9WcveEjWIqo4vN232jt
0ikb6LAh8Jt+o9ZRRfSnOtQuFFYEKrAMmrNi6yOFxuH5IWlUk7v2fJpP0NHy6wU4
nRBO6+yhMR8IRUXiIALT387l/3a84lvD5ssUc5oWiIiR8aJMYuvtw1S6lSFBQq22
0AT4ebBfanRbjWbtqy346ZiwkU6MwWkKPpODLYt9EIN7pnz7VizNb0+TO/1JSYS2
umwjVKmzs58ZX8pvqzN/wJhl5OF4+2gHCKYyaQGV7Btcu9WgBpNlHm9uedkV0Sfx
klQEIIVmN4AyKoW9dhuB4M345UKuXFnp79KoBJ4HkGNPx+Ouu4+Yn16eGx348vAI
aej6e8HMYz0TzeGxzKFWU54goxIlD6qX05+Ryq4Y3ASyobWx2gDsR1L7yuNghq6J
XtWGkigAKYhngpA1Wk11AZWjqz6cZaFQVF9BklJKBDPS2f+jOlbifcyI59zFsQGx
0Z18cjU9vk5bgAE77XkU5Pd2S3X3oJUhFac+MbiTKN5r/Nup9TfjgbY2YyOjSS++
ocQlT/Ddx/SWEFBGSn71R7v5eWGLKabRsHQBpwMgxwn1YHTfYACGSoVB5oIckuDU
Kjg+/5dwgWXpjpmd3n3QPm+eQXc0whEBy1VGE8RkRr3gG5FAgmuPxiufzVrW/be4
9mBeGYXaYOuq0OpEmQ579OXLpqhfA2t6lKLX7Grdb4kVgAK2zTpdkOCES0PyOeaw
+Dl91cSP4pAteABg+crePqtBtRnHtqWsD4yjpC7e0LA4awc0mkrI7Wm+zO7UFq0S
3PBA8/X/t1LU6zszurStSL9U51xlCERiB2nlM5HwgQJswcCOsXvmAv4/QlXwgWeM
guFQ5hCgEp8uX5li5rFc02pflmtHRGG5c/ZRhclE5dok5owMQKePmk9+hgfSw0/6
HkrEKdwG3mHE7QfgwTxFPSOfxRB2CsMTsPiQ+sQ/JocamXNkWqLNwGyLs+LxPqFp
3HVvsjtbxbiOUNZDzXypLjpHSmMamylpVPqcfRuqorMX80ArZyRpbSAQt1rTzZmY
XO4XBuI1+0x4LFjFwwwjquqRlSj4mM9Tv9t9IpldDsuhnlDiYoNtODzetZJnV4Ow
Zbni5GWgLnbEPIR5hbQy26K3j+Boie1jm7AgWXaV9pzBq+dfENt2iP/KWfsI8Dpe
O8Zu8+eJcyRc3zec40+6/bLe39o3kMo2dkmyTrObB8cK/Cme10ifCmw+eUk/9f49
zW3ROA4qJGlhPXGwcEMTwl9cbsUNszZuvVLgjrdw7P2xOIpw4sYtm6HKXIu6zqGl
qQIlIKv9a7pfZwXM7YJQAXXq9pZhAzCqYl78dFw7a//TamwcnXfWN4Igl++q+T9q
ohUs77sKO0MQ4r680BI0prL83WaT4+HXs89jSiAX5JbQS1k61aR//BuKQnAwW6DS
IsBQWPPyBD+lX2zOkUX8R29t1o20It1CW3nNtwKKy8hif+14wc4em/dT9zsb7tZx
+hzbMMCu/8OwnG8wnxd+kwEsztqF6zTbv26zoLFroyP9WubgvvxavBFYAHKqDXlh
nfNyRzwyNCi1c4p1AH+8KuVA2v8fw8BBza1tXqOHsYeMsfTbzSotYtbWY3wESgBi
phAkvSSpbLGYmYbr0+dHb/1vJzeGYnWXNWgzNv4pH63CqFDoycGPtXjyjUIMDnzd
x/7eQIUzuT7rKBcjbVHcXliF2x78uiwademUnF0Ly0AQpSCJ6xH6IRlcsnqjePeS
w7L3ZlLBIGlNi+YgsFTSgXbf7J6iWDywou10I+VnrXFGe5UJO+iGOdwBrmw07+a5
clMdThrL1IMOBaDk3WBFSqKt4ht6pgAvhN9A2GP6BLSGh9sxzxkmDzBtZ7EtNhv0
xXOmIw/L/LTQmGh+KxUwuUpnqZ6UcrNqz2dmQaj6bxytR2U+u93iHOYUW38/fbqS
mMiEetL1UVukjc6+3Ccqp9Blk4AgLYCq0m8kwS2BH64DkYMHwlPLLRufv+JWSvuQ
aN01S82gieAyGwcYcC4t9H1hWwrCWA/6Vqo6FGV0SNQa/tXkJuLUjw2tCpNtInoa
9QO+bADFtoSPR6+bgvFzWBs07/ekAx0Tz6OLPWl6m5zqCEV3/bYlcQ65mgnBqaEQ
wecy3wYjimcBmaQgGCVhyDUJvmvbiCyYtuGH4xgp30GLdpG/YCYkOy9T+eiyh4sY
Hdv17gAi0evQgl6Nc/oLhdCdCbqj8BqIMci6i02V++zbNsyYMkYmdI5OvGSlOWDJ
Y29lCZhRkplN9ZESkmIQbrOVerQ1nWxKJ6mj8fQBxFZdxnf6PAtoxlLgYKRerw//
hpDWWyAWF0WgwuSbN0utt50IpLQq/0BeKrECJ20v/XUvBTH2vRV9RTzck+3mV/x2
2xOVer6FgwhoI829Bn+3LoKf7CUk/7cnwZ+xxc40iSXi1AhyG4qtyC3Mku34b8GA
5mgiE+kieZxGDes+bHbiwaQ8mzcnl3+xG1XqzvcgkWgWRd5nfVafK7LkMRWiulRB
FCf/wbWHcgva0vWgI2nTSI/ZBBR7NHDhRRsviNB+tISvZ2qQIm8KadgU2fDvloJJ
QIMAOzY0FtrFfHgPWHw+0OJcOSfSrQiHO9MrdMqVJCfOhigAk4jmDwyBveeUHLIp
SVC63cWN+j8StggYJSVZarlP5ul4AwhY7iMi7RFyoK+xJmvDnOZ1et+EHKxxQ/2t
QSxiqzaU9K6MTi0l8p7p44FsSzIjZeEWfriB6tZit5m1PI+YrZEzxscXg0NeBBzN
sMh0//oRXOTOLT4MYTOcmqgblW+NxySdDL1hBBELFLh1K0pLqtOqjVnNHDPwqs7E
cw1FaRVIXG3l5flTIwkIsePvCV8qkXxGfa6kl7Uuu6DvowmqZDZoiSuEXT3dRBkt
ZKZ8XoCFibnzh6jp9KLnTXHIKqiwxAL5qNkqGAiLaHJqs0Csp6zPN1NWybw9QJPe
CVJOonIH1fBrs2YmbMtud0uG2suQI4hkgrh7P2Hw8lcB/AIwyOCFU0sCEIH2YoZB
0l+oxSKbJ4y2z9ZR4wJ7+AHbbhKRDOZ3lJj2mOZ8fR6515UAp7jBoUwNVccSBgBS
A8ulW3bwkWrUYgFeC5VKumQXwbLMMO4ywA2dblrragu/LP/gyBx4sWKC0zJOuWtC
G5HWQ+VRc+gfYyTT2Or6mrNbcSQXIkxYLRPfCTKSeyDYuWx/1moQ0FcbP57Rr1LH
996xlChknJkr4SOUYhaSwTWIs99ekj6GTtBtEQLwtLa4qjZxXE5hQIuxWbU64ZhL
UQIgd9bmB5mpOXbarhgISxLiV3B2p7z10gnVUtjUJ26Lyegeiku1NdxiwJyKMOTp
6pgEgBeClbJHtvHtM1dFn9vrL4kt9LdNsQKE0OsqgQr1NXMZqFyr0jQjeAA5Aa90
0wTJS1i10o7HGOuhNX03cSWHcWHLeOv7Ikz6QzMfP3K4PigAGbp4QXPDwz88uNYU
WDOVHCRx3voKd8gs2/ZOvwq4Ie4tKDoUcoaoRuwnBRg6lMK/SgbgBic1FXa7lnZQ
9Sq0KX9aO/xEJqi2YEaYyM2aicHfFyGkkSef7e8mpLnGMg1/pahJKJ+IJA/VDUKq
uwbIOPzkF5NcQSWPYpudTPsffS9WMGyB16MOPPTKJh1zibZhfamnjRcfW+pwS4eH
/803RJrN0VK3nVfMxqvk/lJk4PhBWB56P8CX9OXzVATz661CFPkrzh/DynarDSqZ
AI1muN59iM1K/jLEMagktZbfwGzrb1hIolfv/Ugf7rh3SIKGXXWtEyr82COS0fDt
JXa/t4BWk2lfKYln8nmDi7Tsu4/9HTWnoiXxqbxUvn9um6TKa9hgyfMFd3wjndd4
Qq5Kj8VE/7AGZVRVEOdLGZkYbEn6VQzt2igiU5r0GYvUxf6xGZU0e+NBewZ94RdZ
oT2/JX340l9/ycHyfcxSpJIseZWw3IKQm6koy+wiXWSIt4tU3gOVtUvvG3DWT4Qi
dwPP17BQfvlW0zFeXHLPmlBReiYUbcVfY1F0M4C0NdZvD06YQSehNg4eMwuPp69h
hMm52h4bUrXa7CJ1RIhGjA46ggu76sBDBNOH6mLfDn0djAZNV5vFNjGVioxnwpV+
vzeCjAsidvZC3XA8SyzdV9GhzuIMlYTfsHSd7CEdnlU/+LUl5HAsi/PGIkxdZX+x
P+OvoUa3CF8HpKuItIGnxipgIs3IKOUNsChiYB+kTlSV3KAsFWpB4NhNDkQx5o5F
S6lwj/ObQ6d2sMJQ826sfSK+SoReAQueyM7HCHJlEiaSK+U+5dqP/pkGpBJz+NoA
7xNi0ASPRCGssHazSg/3YTJkITEk2wXZJng63ikh7/odHyObclOHkgt8TZwKYCez
dPktygal+3DQzYXJ+jEgV2CKpS4OizMF7NPJtWemM/W3HRyTi6jylol73FVLpioH
fOE9osFN0ktrH1/oiuU57Z4XZWSrxWJDNAuItkPiGOXeSJbFhhioU1qcLmW2OIuK
KksxGH6MkV3h6uG2yRea3ejU3Zjt2q3EwJxlVFRCiFp++BT32xD2SzG4z7xSv2yd
x1A1MlegMAi6+RWPWo2OewGhjX4Y58h4zZGuHo8c4jLTwzhgKh2cHMqXNpcigINt
55vZ6AVSeWy7rTehmuwTTPtL+iVWfhBK3XogWynmSzQYzza16hFC23HC99pq9HWH
8DkbkqpnCKTEE9khaeCUjgzIpmVkp7oMH9rSFZIeSx9K2edr8yFglYaWjrbBKmzb
PG/us4mgap3dcmA7kgg7vwbLfDvCmEc/C8od3PStgfmUMV5q9AkDRySnQr7cFs7B
a2bnGSjCUzFFSPEFa0owuZdkr7eQhG7fd8fL3qT9Wl1LxbLVesibUrPsNW9xngN/
4/fnHcxGE5mZMn4vNM+L1KQh6PUdhTbi06p4WBR4mtKxE4rjr9Xx6TgX9GsIYaGt
eA7cTM47SS7TXWkx7nJucYtH+wsrB0laoVZuAnPmaMCUxJPIRn/OHtuBOqd/qT7u
DR0xJ05imc5FZFI/e8oPnf1Dvb/SGS0EpDU0lQZhLy0dNhD3A9l9oY4lg0OCsG31
kVhzEDUqO603QnAZIoDkNzJgiVHeB9qXMMrV69Tl4Dr+ou+jLTP36nfL9JnV3ltN
59fO7CqXsEAXCu8IBubcLNjZxZAdxtZwYIIAqnWFibjAkvWn0rg4X+e+GktLRLvE
vJ/Nbazh2GblgiunGm+r6akh5NKcNQ2cjqmTUQQcPKv11aHIFE9ROsU5Mq/fCVw1
qokvsZlWn3jAnPUud4g4CjzZrqGIRWkfr2DHgGrt4XtfH9PZua31liDF5g3jJ//0
puEo99X3d4jUY0sYpf3ly+CHM/yJWebpzGwM+fN4iuqwX3pLoV1YpyjNBsXe7vS5
JDfG4HGBJx1+NcFgqPzQYbLRciwgG1ljSv+Y2ia1JpChPwwmmASEM/eo2iaTNs06
xK1kxTUT/erW7ypJU97nfZaJ6OMKj/UpnUzQefc26eC6cHfR01jJnLN6GOxeHK8L
eEnlVOMcytl+cHYErDFsaXzjsEVkkS/Z8wKOxVt61L/fBKyL81NwizKjDL5M0o3G
G1NKAC4/RFX4bVKMU696ZI5LDOg+cutk3yd+Lne3YOZveWzEgOOt2YEC6qkF4vz8
CLyh9aJ/vC1n76tKxcvNUgeBNzIeQf2Nfem3ZEaL+FEZbCPEYQcSv/Ar4oaZpMLV
a7YXUX1aBe6mNGhjtPlHc2ulkobPAn+NLW/yLkbyGfkQEqOXJnfe+I1K0rtsJ0Uf
bZ3Tfur/4g9WWbKkMRTuDkF9z+8d7ZSP3Y0tFFJUkrz6NFPiwbhjQLS7hdH6VxqW
zfzRFStVo0isXsh514OQ5o5v1T3c/6/aOxWCGpebaCKy7HB0TfD3E0M6hqIEgZbZ
QqBUATwgK7krBzwEvbVeZrLRoqWIeLPS+kTiGJD4t6NFLA06ou2WjI9yWKjmGuWX
k0U+28nqM6m4vrZ79PuzqEx1rU5WfJ10Qj9OBYEkgVLmRJv7N4uY+XBs/bS7To/s
RVEuIUMLz/vDijC5ieTAu/mO/AMh2iJQ/UcY9guK5uXPtOlzuh1eeDmOtc0UGZjE
q3J8rAtl+wJ9w3ZVd5T5420InW8IYZhjxaej+Vu4uV90PLEVTnU9jAvSSVV5na4f
4ox1b6Ev54M6RPGSZZCRAop0EBszSUo1+iNFTHNUMlfadYs/AdYqjNrd63pk8rfz
AyxjH0MX1nO/TIdSLeA19tsKa22enFw0z2lE4B6vHrJbmVbaBrPk3SHnI2DFridO
5AZFF6UNlAF4dxRkQHy2yqFi4Pr/KuyGn1vI/lD6UYveTjkTplCiYMn0lU5ouXty
4mYQ1yvZe4ID43vyvqI7d++d+xlbXj0r4QRRrgs5ClhmA3dV1CSyvrzzNpvtO30P
zyU0481zU5v6cjx950ZeSxVKfzxAiWH57uYgc85rzY6bxcjy0XKqGLfO8N4rdGWv
L1sVDVB1uu8MkJzi7a+/A4o20gm7BPPmOScC+uLrTHF62eNZLIH6pHACjI58fYQU
ZC5PNwNSlgEbCBtAW9/LgyV2XcrPyWQoq+h+Q8XFZfXC1mdkNjtMldB38OekidNI
4Bhih/XxNxAicQgpAGKXjicvcQfEh+RnINXhon5dzBVI6gG1k0kRsC8kfSLaM1GJ
HrDmSmymooINKgcooLY3A2sPvkQd4WVfm96BhtFDaZyaZ38f9naZZ5BlwTiVuQ6v
u1VsLsA6gX4v9GllqNRNoteIjhlGJ4juCWnb7l5UepzMmMDvipr099AZQPAac5nc
um0XGtt+R071oxHIO6m55I3K6/6jQGsbArxVxOoHT9LEu5tH/1YUSg8Glry2sm9M
64FhacfL/FJYNVc+WUfJhQMYxqytAeH8PY9Uz7/tP28H2REX5FXhM0T8Ex7dWIvN
85iIpn6zfdIWBFtLj6ltDk3fxxYa6KTdN6gm3LjjhGm04ttL8Qcy73HPWa8866iZ
oEqy2KmUaEwqdCLtLTp43s3rXs2AmjoelpzUA/xJip9rMVr315X8rElXryWpliQN
io7hTAY0MMYgmi+47FYAFL4SMvu5oTsdhpypF/uTCY/pZ4Vguj6xDz7OW3C9wssh
i5NaeCn0AYw2uiemnxzVkvydSgUmMFPcdOGt4+cF1QYBGI6Oi29aYp8Qt3Zx/3u6
zk8AjufZihEVlD9HzgtEfyJcoMSu1C3scgciurwFhLun962yYxpabqxy/odEbYhA
b3Ag5FhmPcQR5+EzWJzfck2z9pwI06Pkdoa2eQZKmUEl0DnSmpQaGq41cYZGEfCY
RDB7t71sVe4pEO7qg74g0idMTbhaC+eGyGQwGtTKqnqdanf/Ya6JzDD6ZQ9jswze
Ddnd45cEDO1NPkI5q09RHb4j3imAgGEArvnUsQ5ug+/U/+yBIrHBN9MNN1edVw6H
IlMjG1o1xAW/0tuHjSCbODEQP2PYGf4ghWNYqZsoowDrjRTRWGxtwYXzPiK98LGu
etkeG5+SzqNCL5udsORlci6b5t79BRKqzEA8qQPeic2bM7x/les/hOumwSEsqbGq
8QAIYobP7C4fvbxaJWKVgKagN3IZ/3sV1wDSp38FI/C0IWzgh6KIp+GF+Jux1D3c
b8VTbsZr1IpbDBwHOC3VtoXTFOPCMZvzkP4CFk+0oTPHDXk3Bdg+YRXCsuCSZaJy
40BenOs129iolFF8mywIHXuvWqwSSTvGNqZDXMLQ0WwkScEE0GqKxi+Ddjd3BUEt
T5BxyLpWLDYDZx7u+48qvG6hEvgXxX4nyQzpzZF+ZIxWWcELJW8ZE5MS4NBTQCiQ
N83uaz0iWXjc8yXpQxNb9mw7UEpiAk/63Zw4H3qngYIzqO1yOrKHoxOb1DT7S6Ja
yWd0D4fTNG/nMeWixZk3wekqRPlAJbepCmxGSyp4vsjxL1LAiYeH8aEE1IC+tgvI
TyMRdltZd+COoHXn/q8jhBqvvNyZ80l7SNnPs7h9S4xR6vJhLABEgEuCBd7PRG/j
V5KR0vrufpF9QG62cZb2GcNF7XAVb41IB0MnvO7WYkezoN4lB7yupBY4OD7kT7T+
aVYPKQYVLAbeTHnWjxNLfNu+w//89f36P2UFmxNTy9qabBVl0ONOBSrdsNbC0qjF
HWqiPQ8Nsxf3B4Rthn3/7HBEjYNjfI3X6gUbjHHoO9QRvjJVz5GbgdkF6MX6yd99
iYI/KOYSiNiY5kpvzBsFAYuh2xMp10C0KVqHWpVryXzWV2wBoMNbElkpmBQaAIbw
X5MvXh19DVJckL+BfshorsX6TsvIWkiJaB2+cosLI942CePJm5CfsDZ+j2CYaPuH
9WpaIL9di4VsWtlTlf5Avr6Nvp2G7AYCZuMAuv41hIzoX6OZZ2bZpGLATZBk40Rk
L60mY7Pbf4F/CuubA1kClIcCyC2H79/fFvfNs7jIVkKC9iSG9GLOAZDPP5HXSsA4
oQQIEjIITOeimWwUWadduzVMaRSWC/0B0BFxvzd4IMbicNtXG2lPusY7SpL7yPlD
3pIpUzC5bp9iBhYAHK8usR3Tj/QjsZuQkCTr0tUfA2o9X8wTqzdMkOXKEHUxQGx9
oXz5KkCR1GBeubeKPXzgL36g6cRFE3dDoE2/R1afVcHNbAjhTmWjCqybyx4fCMl3
YJulW1LJOXCNMCtR8k84YOllBzZpnWB8fvuA7fR7X/FabuOrCI7WTIR3Z4us8jCh
FNe07IcH2yVcmMSPYFaFQsg2QH+zGk7OnFAP7xqr5pmUXPV24VqmGll7GXidt8/K
qJDRNka3rtDQgKN4WGfc0Xcu6ffJYvWklKDOtihUL2YO86Wo2WYq1CMUjsmO6HCU
Pjx4mcbHYhCldwLOEV0oo9kIjCaa350DJKzipttgXN2SyD23w5ps8gCFS+PxvIhq
42Vao+jSWkNDJnNKU0zzkDRWrUU/tq3O92NfninYtmsU+xvaEcZhRV3xGlNAekfP
ZWGT5lyJ6uOcd6YMWiYJ732y5lmgxtQxtRnUCc0oCqEpbxigB8vGT0toN0njF74b
EW4kDMhTH6k8EyPxMrG5d5HHJQr8+grhAgvQwrp8oWEj98OdCDB78PjMoxI66Gu0
ztkQu6dWDw+pdOHP26rtDx7xiDne7ZKlnuXD8kUpEmAO3vwAdvs8lE+arrrjNKJU
8P9k/vm3HQzzrErK7thylw7aVb8p83dew0eqFpAJMzPx2oVPJUetGltMFGUMigBL
AJmdZ7EwOEz8Tn55SeSheUIv//4wliH7B6dQsDgDyyBAaHOIYCK8qxkDPOJ6iMYY
uzDCi0MM76YwjeU6RyjfrPgtKfPEJtDtHBIQNAUtWvuJr+XeEeB+3EKiSiAfiTr/
TdVZUhrcxidbTw42bA/Ut2Iy6doRB8mix4szzHWVbhv/WP2i3MUEMvSFaGfiDTh9
Na3vIe1iV6/n3ez5ejcTKmz7KzowmaHdy3YWSOd4m1e5718ipI4wZ7T+s/CJPUC9
44Yieeo9EqWWCcUxHJfsql6rsVpKBbzl7wpIacUHv4b2F1webFuMrK1cONSzk3r9
aAWoBke9XdBD9L0MgO4c1FhwbfIdlqeLT5fPj49BfhoBuZjyQdn72lKRrvItjFNo
lsGrgCh2C+pL7c5Xh1oLJZxtRRrxa52cDxmdcKG2NZlWhVR5PBq5ecY4V34vw4vi
7GbhLbz1Tjp2A7awfs8tKuCf+gA1IbtoXMpqbw79yvNMrEuou19XtMVIpDl7UYoo
fx8ljo6kRrVrbk/fIphq8X8RWwEobqmsosziVQ9EgJjd9zsPHu5BoN+LWogH/b0r
ug+4IMBWbtykegCGcY7iieKUPj1cawrSw4UumA5y9+s+h0O+ambttY9fhYLdlqjT
0KFjReqP/Zu0/8QgseI+LjwaYgeFftAaImL1kU5sVrIVuURy8E5J/y3k6dIMscee
o+feLm/XJxOzCsBVVcLlJO81sTMvTVhUBgpPDMcuI2LkL7IVxyc2xF2HadFhzEYs
FKVxKAsypKc6vamZF6F4J64u4jQj3JezyjIfq6YZTDevz1P7qlvtjc8Q3NbNfeWq
t9A6nAzlHeiMjNZRziozAOyvzLUfjZ3mi5M+pTyOLfjlKg67o7iHezPfPKUDWuK8
Hi/uBkPO0JsMZVbfTXnEwmfdXXx83PhIaOGgbeBepdrKvPpdtxFgHakh2As4WjZs
4JDuQ/ciHLcUh6A21QRLTMOZZL9CrRHsDQgPsaCV3JHy9PJwi2bLWYWjC4aT2x16
ceoKPYgD5OAXe74FDs32I7INgwGC6w5u2g+9aG0l3PT0gLu7V4zSMfWT4obMthiy
twW/ogBWWUd3TlBu7C0ym3f3Bk/D/eTP1YC0c6OSwXyIq9GJl9YQmJsQj6nP6wEZ
iaLX4+MxtJjfp1byGYk9NRsWNttJLXxlF5ua0l1fKlnJa3J4XGVJ0dw2Kqs9eBd+
V+0j/BroglLL+qzjXDNhnSK1KfXRWLd9/PHHAJHQ0ykr4pw/gAckZoyGdjBff4YI
lVULo4yxvTrappgmgTLMNeMcsNaf3qfO2S2AYEC9Uqc1s4xyFHxyxZs/nU0iXAKS
wCwvaiZ11TwB+lSx0k5VqXGZ8L/eLCcO2WBWf6kBcEf1oNxxnGw/p23iPu00h2s5
k8z4h/yTRrc9CAg0+BzP+DM2mqhVzO5fKBsFXg3yFm0COnhQu2gG+fL2YxV5IP/C
opn7XKZzEsMrI99YE4WSJ2XrkjfJ+kuo/3H7+9gO485cBa8+4yTuKCOX3jHStptk
ZaeKbJGyFLiyGHLWq3nW/rZOKQxXVsLjYDEs3ed9NCp+j6vmhgdNa5Y8bIHYpviz
eIx+y+Jg946VEsJQt4WzuZDC0lhZDvMa4MVdL7Eb+sz7wWKF8o5JquVKf8uxkT0O
bROB5oNQrpKBwZrN3VRGUvNiL/GBHwtIWIgLgliOigrBumxdlLgaUp1PtkW6Jaie
EDwz5COj4uhuBEfr49xdiGa4tDYDUlP483VwFr8Li8fxiNHtDqJljqwEq43tQFoL
yJsQbBgS+Kp0jfmOPtAylBH2E3YCUmM7ZykDXZ3lpOypES25lAIGIiPnG7jko3ss
NHPNMr5XFIONtt7tujzOb9+lrRyqdOgwe8zuyGDnpWpb8oLXXUNtYxbE+IP0eYvF
3KqVhYizPrvAt0YsGndTCgh/qB2+GvnVyI5oNAPrJS66GMEozgUcpTVoTiSWf0gT
rzzdIf05xUU6M78dD+gnXFf8LvxsWxcgw7HKinjr5iXiCKkiO4Z2bHsl3vNOUTa4
rOtiTY2J07ahmu8ek7QuX3Dy08CkX2gfWldE6z8RnqE7PdaaFP5gQJHgpUzgBoIZ
OROuANtx//rmSYUnmOTO0mLq0wQ6oGabma6qhzcMvTe+jJsGrxLJwYciBdawr+7N
v9o0xZq7RdjyLKFrofz28dRzO22uwlfLC5kBOMrHHyl5l1iedTHw9z0//Y/e7S7s
aMw0EvTZsU1DcXdtv+PR+lKcXFzDY8Zm9soosSOMUIzAXqWlr8Yt8LkRnyLiyRGf
dU7t2N2+w3rh3CEM9chQc6bMI9ElA+2hBlMDj4B3fZs+fv2uZ9YAAbxObq+SKYfp
GSHrn4GSIGh8uXQRdiOCTl5SEkw/jWmGniIAyFbH5d9MX7MtARnc4hDifjsUXlgV
fJD6rfcoZKNxF2P4xNrHzcwWokHNUqou7lN3HCYZnMDpNAXM1C1zAu0nfuSsjuT+
AO8EJB43CNY2CrtQJ+y/oMM64slpljkJK2oACPJquGf5QIm32SNThsVLR4RpYAQi
coVMBIy4Y1MI8L+kt+xHa3DYYm98HVG/pO2W0mTDIZd+nu7q8bKjZEG0iyc20Ku1
VJMHZwHyL0uI/oijuP93PhnxxWONcp15lT3b1V76mKDVj6M4CnMQZ/s/ky/R87He
0BUSow8jp0edB4v8oYQ0ggzCEHHKgu3pTi/BDpkBRYQ+xgTTCqNV77fBwdz8uuxs
BdT/ICXrIw5yQRrFd5jGC5o8ArXdcAhE9AxhSdaoSzDN2kIrotr7Ssxpb6dGj9e9
vrwzFLGbLo9+pS8z9ebWwwRpEHUu2wsykCBRkSPYnosPEUlcjU0OgrNDDRqlklPU
ERGQ0r72YHToafhYW0PYtukvbsXmP8KySVr9ZBKsmCmqRRtw3iCFjl4PApICCsV+
wd0kRAI7w97pEDY9Qf/kVGtoDM/hhREPnFMDC6I8qXtCTdahY7FUqGFiQWIwoOAT
o3uzQpqittXGXWhzkaiSDCRDOxzU7IifWI9yjgUvGOdZDWPpMp8edjbs32xAqpQr
klEoq9pV+yVURSqqhID6Gyg1LJFk4crQqxm8DCEYAQkz9yNbqqQL3SVoeQ3UBPPq
jemNh+w8nbw7E051rJbhmtLAyiu4BnkmG88iSqw5HBTIwdNuIxB6z5ChY/KoMwtt
o537jiMp64NPwfOfHI6Kd9PmHu/dHsHLdfc4fN658tDwOlkhAFJGvDd2waDUtlGf
a1wrQJseXodEOVF3h/x/WdVCMgVUnCypRpyV8oM+d2g0h1nAMyAFSN4c87ZnlvI8
plhyr3dBCxamzMiZjCtGAyHgH/Mt4mbdE3cjSrcbuFGW/0xlwgjCPx3WKu/1wCKk
02Hs72r9Cgmu8JDrkra99FjRWq3BN0SKVtmPWmFGKveYcvYyvAcHkvCtF7241reU
e2Uy3PyNiYQu1r0GKkDAqEslKL6tDJkWWhccLxH0eNdmI7aFy4Z3SyU7jB0BbCYY
Gc94ZzSE5TuWFEpkeJ2TWK8udGEbG4Vbb9LZb0oAy0N1DHsB4oPMOqtpNwIDkFaE
91GYoRYsEpXP29XflEdDGP681AGkaU/T0YZg2KmIHoqfkEzAL7vUj3xu2Shh3Xt4
HZjNnHrvxy/nnqF5zU3JHjxcsVBRr74FSF5S/BNocoJd95lfgsBHdR9eSff0iFQP
nsF2yB1Wbr6ALSOjYqX3aV7R/FEHxKxa88H+AXYcu4mJCPncbY2awEgZJ14MncJu
DWUN3Te2U1c2gWal+JVq/uLkf5SKhvVJFJplpazTRCAPkKC6gb4KoFrjKEuhVifg
GUNajL9syUMPjBNhfzN1V3vKBm4rq0yeGbPjORPSz7O0cd9GrrrQGHiIAxvBIJgK
T61ml813wiLE+1qzs4MnEnlTTFgD0qpiVOkaL4YNOSbU2FkVkIvtDbkzl+QMAURX
hK4Pbd0fhJ1Jmjc1QTk1dVBswAtF6SZNud80414ELIawS4ZazZlyH2ijKjCrokQN
a+S53SHVPo2ltV+5WuRM4yuKpDSUSbUq+rg3yIqkTfwQkmb5sdiaAwOgQ7Q43E8H
QJA3KjBDTzYTqprWIrm5TbJCCaOczBYxaR8u7Rz9yRzioggmLhonmZsd2YV17D06
hNH1xs+YAcJSaSEiCvbpa0yqUNoKt9ylqXDVGQuhMiB4ROhxkMqMo6oZ8sf57BDa
eQjzXc65CdQ6QXXu6EucCUryLNkHz5GA6JBjXj5ypekhfyyCFKFCzM70i6tFqfNK
pqBSb0DDDvyZkqFcBOydx42T6SZilTIQbP8n9Cd/beOB/cl1KC3CGHDcez87eSeG
gA1nytaEq7XqBS2q9kKkU7KfSETEmeTnfrJbIveG126RanZmh4uAZX1XQMumxNls
3uHVmB5tyibOWyaIYp9pbAvqsvhHf9AjU713hLElslQQbJ8mejsZWKRP3a+HFPIA
3IvQTlHAXCbN6+kplaS8DxGVCAZItjOwUT8She+OCf3t2dpeoqs1aL/j3vtGgJ/r
Y08hSCcy7uqte4dN2PdEm7zY4wgGJALOQpBoKvskja0ON6QPTfHBUddUDFj3Yeu0
vrxVmjOGUnJ3TOSjb0fUPEuG2/rfA3u7UHMtxMW+vQWTJRKrznJXfN2Kh4nF94ky
igVdYVYJHIxFK2gIVVTgNw9cUpEV1evgOwGyexcXtY4UY7OVMd6lg8qDrQ1JTr0a
T/hroH6ayn9KIfPxJwGUjTfC5JkerErIryqVPItfHAe/XhId9hT6xbp7dtVA82A+
3mVulHZUMFOYLYbiceHX4VZfsxhi2CDM3uPix+uhvBmbzd52O75tF8tEDKdaQPOd
D6r81A28kyL7XblWS2VKIEhbi8QIgZvDYEOjKKxwGj1ZlEkk0BbM1z71b87gA48A
jE3/drQ72WhbcvEhbryuDdfKHqmI+CWwJVZ0+/I6CfImR+wJh1zSyx+SkU/esKmI
hfh6Qh8UMGRfwUE8wtsWjmmMA0l/35a1UHCt+wylPD5i0nLxoHYGmcAlwkWvbb49
0Geum7u3oXdHBBr7C7WkRcu/VSs1TWzdLrXA5b1cMVf9v9DkOinP6nbiaAFL9iGh
FFLpCJ1tt+alnEu0t4mRnmB2aDweQ/ypESeac7CdLWQvrT3+qzAgAgTbVFF87NC8
zPCbmll6yaydz4jbZ3z80xcTdNBFdlv7USN2kL3887qD2x9g29AoYYcFFFbfPehc
K/imRK5qjXESTEhZiVaPtmx9sCecbuYxyWwSeuTiXvVqmfa9ArYg9rmhhLW3Rzko
V3UXk9h69yIPdzffSXX0uFX/hVKpoTPmML2qEvGYHDHkqjkIGRpeUsIiGZFLE/Wk
aAygzkpbrmgBKkWoSSSVn0NGm0jd6sUJSk3yO4/EMIVYorPXaDfKY6/yAk/cHCQT
iTD2AWj2X+OfXE9xLsCcRtHshffNizkW2xnKW4G+rPNVmRbbnth9zpUMZfbQNrjH
Q1ZQXA7BQceLKp3CFi+n9avGikpzKo5pvmNHM8AUQSfwX8u6Fj7fvpT099TCsZCK
bpHbYHoZqZx74SPEbs8o/lqJw18qEMKZBhQz3FWd8qWABpyoKoG3nNL/zWviR3bt
TDfihG3Sxu0EMuYl1fkMlVdvaxX+twH1zoB3ZpJkFgJCTCkCyk0t+OD1e+1wfFL4
PtMPtSs8rFryPsE1z//2d+LkoCYwsfFe3heTmsQcs2Mk/EyGYVo3Cycq/qSpqejO
7WPWqyo6eXiG+u7ttV4kTKaRavE8etytddg1wA+34/JLhDqWYOVVMCHehNojJVbx
6zS9TOG6yp6pON+9SMTq5pvSeZMMVYcUkQP6CuUpRv5695E/5isx3TecSXFlC7xM
QeYUP4qkCxmxX/9y4Vr0BozLyUXMsF0DyHc4PKWGOtuTYMMlU2E31AS5aQKnweqs
HUnFzIp+Oi0JgdoVoJgo5iY2hGHWefcKX+b1uWz8/Bezfc1rxuHM6+wcEucsk31B
s5tCaGWlhiii108Aw6SykcgpgtJZi3pXD6Ml+ltb+Df3SGcCRUkKCuFg9RCPU5T3
JztkTU+X6PFTz0G1Q/HbACdktL2GNJJF8xunITuYrBDYsrladnZR5ygUsKswxPX1
Trzpxz51l/h34I+K+tAKKaYDn/7caCmRZ1Qz8nq2x3+zJvBukoFR1iXQedzihgUS
CsfLg/3o8SvnhVmKjx+F6eclLtESu+2o+6qk92R0DcBMkKKH/JmM0XA7k+toln0a
wWjEH+WauWeoSrnTmGqPExhEmeT9mJ4Q4Lmh+ZAo/obXkwVgEgBGZxMKyqH0crba
wvRhJVPo8Q/XPCanzHBQid2CD8E4ZXVAb7p71i+Opna0tLuz3RWl06k9OFlA1RYM
QIr8F83RyjHVc674whoIcv96lDoi7cVkhM8YDRZO/ZztQ7g8Za5bQK17jtY97Voz
XQpc4hUW5CZ2o16cLTAXkKatP7WItaz+ikNOK/vgF7Yv2y/bhHIzqSy8+oJ3SCnH
8hLrPZ0e8xBMYb6CBM8fjsbEzGU2HdP876jzU+itBXzlwihPD8x8q8QnvkkJ7hOL
kANrOTmWCmrZ90MjjMxKkRjisrnXXMoOr3yqyHGwsoz5So6YSIVKyMrcjqNqvsbd
2akL0Y2Qkpuybgmuu6yZyhEQwOOJQDx5Xu2XznsLWPYdtP5q0ZxUiV6T/T8x7+RU
x8nT/2MszikM2c0X7s4OBuuy8NpXfGXCpjyceUfPVc/7SFTvBtHm+b7l8Rt7z+dQ
I8/0Uvi7hC3Ppcyw2HwRfjsKwAwHC5oQb0UMLzTQq54CV4xM7EOG1f/8cKtc2VQW
8xlcgn3qHqh53ozLYTOhyB0FGXjRlM6n+5dvUh03DiEPo0+0uPNZWalafIfz/Cxm
LbSfZJUL7HCnXIHtbQb/JmlKk4fKV4LQ8mauoe3A8CULMz1t2gg+2qQXhYsGSFz5
pf76Ma5kKD+PoXX78preSkxH0VbJK5Z3E3aJCLMMGcu06PfoB+Q4JneeX5YIdBly
EyXmmo9lBmQapAzJkwryXpcVyQZmbcNvZDQAyRTw8adnTEy9dHbg8fR7Xuhqn8B5
nmf0BEFI5IC8U7wEiOL4MzSlXfkEnR8ncicp5PFsQ/Mspamh6U9eDQmLm8V4oQ2J
fNWdAv+aAvls3/i782J9JyETBK4OoO1t+i2mHL5v/U4nmenhmvBNdYYNhIYVnem8
I1ilCHOXVZXIoX7fMlhTZzckRkgaoaUGZdhMKd9o7yPL534haOl8vxclG8lSZfOW
0iTKbBdJADwkpb2WorQMjBt1qQD6Do3ITccUyktfYBfHe2otYTuGYE+5vnKSGMzY
2xGDhA1ymESDCAWDjUQ9/Ie0WvX/IUlkV6W/RZQQRY8bxUwTXSUgj61B7GTusP7g
0xv2u90vWzqGObSHr9fNR75qtV2g8G5q2ovTURjR/yjlR4nNYoeR7Cewm27rYNKe
vKAljV3Gl9Bez/KS/NbqMhVdxmAdxIzE6BtKazW8RSx8ghnJzrzjE6eyW41Axnc1
VHt2b6pv+DC/d4CeiSLakKsbhTHRrWPvj1WlxJ7rb2IKKz/0r//BDH/FahF2NdG+
WKnizjMXl5yhhqGtWH15pL7FHrqcOJh+kxSDfRIZ1uX6yCp26abP22Fb0tShmOm0
qVa+C2z0BB88Mqnpv5vNtZs77frQv0SY+u7giiB3sVbjO7yUCYO23iA8WEffeT2e
DsW9uNYiquSM4tpH9nmWNaxU7JnROy4PigWIH8zD/9C74WRpzY2i3ugrvVucunsy
cEVqSvReOvOsuNPAodjSfkI7X3GiiRxM3dayKpNCx7LQNouMtaJ9mUYNle9Ececy
f6oGCeW0JFvDOxsEtwvULxgShPZjq7ikQfTRyLD+CrQQRoyP0eFKZ3OQljr1P/a6
OTOUorBrjZHKgMmV0HMzXYK1Md4L6NzfI4uHA5UM4s6/YoNByG80Dbuqn/VVrFpJ
os3zmLrUFwbep0u66wLdLkenRVYlqlxSe/BEujk4SQjaSXCZPsI/2c9MJN6JHH+E
3CMiMWpzl5S+5xMX9ZjAeGlhCQGm6EQyjhu/UU9zbz16CIxaxoj5wnazMcrsvix4
vTVw/GppRsUfF9OrkmizqZSiJ3ZgMo2v2LHs1e1nVz0tSCzP8+gcPKVuJKmzHomW
4kfbxLw5BV03/IIz9L2P9DoZ6lC3IDrFgM3m5ojRjYZQ2Td/Rj7M8K2iIabc070M
7YJztbDTgehGdTMxafoZweRoY+MRBz8Bie/a4BbcddDlfOTnnWknJXhf/O6PEuJm
UoPcmILPa3MJYUnCCYKiUvhYWE8kVD3WOowHELTCJDJdxWLuzLBTREAZsza60Gpt
HuQyCcm7yT/2bm9TQ9QCVJbvM/Qf4bSEUfgUKjSF0yFN+Z/jWfSBRWVyzua82ip1
9vmYFJN9DiRgJKM1jCkbzLcDDgjCPLj/AowkqMQm/slWcD1Mebml1uFTAS/5mXdT
bNXIakPRU1hdfILQa24x+SNdBlWzIar2ODVgCKIiwAXJcsIRaCux1Tex7HAas+Dp
E6XIqDly3KoOYZCfQUiLJduaZIsJhr+ekg5yNxs0WlQIOTvhwzr5/bri9ZmSScZo
+Pqx7Y7N+1xUx5dHk/H20Rr5nMJfMOe83IzIoG2JUyZwsUE+kI+nUOYmBS1qnFxu
+gUzcKr7IQRzTNjYToYldX655ehP30wnl8Ss0HgTXAy967F+bvkqj+29V+CaHB4B
WAdcvw5bF9QotjOcgE07Zm/nNZZQnEG/327eKlIoHLwRE1XfFWKQKBTyTpskyCMi
gOczyHHRiWDZ/Evb2XKEYBdMRst7CrMz0WfcrGMoK9DSa52ZzMdwzaP39Lf9+uNe
gVnO1Ps9y/dQ5RF28Ylx7XWJjlv7YSI1H4tdGEfl2FeV7+cjVMn9bhWpKv9p0cfs
SaxaecdlpWvWblPjIjRBH1wZjFJ5GgA+J+oHPg0VuuMCo1qqLJaK1ZzuUYzE7D/s
jEG69Ec6L6KpnCs7mFYYJJOVcAFzzV9zXRmS4rXg9h1D51NSX72m53fbSTyAxej/
x2VKO/mp0amr3zHFp/livippf00bKieKcR9q3wDuS5LTA/96KP+K4FnB6xVIIe5i
+InaAYGbH9XM43WOJLsH073PI/Auh7OhJL0VRu/pMJHLzR7oZtaJPKi6yE26pl3W
Gla8VcfWFe0FXtVV18XadoAZUu5qmQribdAEg9qh0I/UdaQmGonuoM3Pfe2+8JKg
iHUbIdxSKuj4t/tyOPH9N94qOHZbxH5ZJ2Mx2AjqDLh2N7ttDeUtFsuRzetDHfck
HRSQmsMhDFfD5zSKUaAuwNtsctRKMyeYH453VIN9gAMLrGB8fSsQedn3RM1PJsMV
561DmEmHIP0mWdFDLFbXbgBkUZbGKigXqPIQroPJm5h6GWssBBpVEJ7p7tGzU6FR
J9yC4I1Ed8nbMEOYNMh+1EynfoaoaS/McKsXswVXXbdEPOpZ71WrH08k9DLQEdyl
NRtmPb3GECWNo+LABvXeas7YXMYBo+Ks7Xn7r/ka1Cd4Ia8dnL7oUQ0tTP1Rxpqf
V1BPm6O2MtoCo7qvKFtYncVlEG5yifIdOkBJrX2CTP+pGJiXC56tb2B/JHv1T2S5
5fxmLKP19etp5U9yudJrMXOSflwDWpo7Fw6KNFQQ3QWG+YglR8r+i8t2Bzx5kWZa
nCJg0WEAtWcuNYxXSBfcK/0UiNWoR1w/WIFMDL8Ef4yHuxHJqfDgBhRb/OcBL5VX
DwigEhv9ojCzBpeKirlZne6zVkwV1zQCPCRTosuuyYPT0JpXUVQgGFMLjfr/Fkl7
LfLFNxmjLyEwJCSX08kJiRf0uB6oGdWioR2xEKAElixhHflMa0Rc+ZdSIbGNSE+8
FoM9DSZo8aZzGWoLVWQAguReSjZNVuSqXftozfI7u0TCchuvhD8VMlbTUkB7rnB8
DZJEHuoEJr7eu8z5RP29ZSaWNMxKnVBx0GlhUD0srKwEsh3OFzPKtQQGpsM10/T3
3Kfd649Dsx7EysdyupyJUORGdPkfblvtj1ECYiz4rchdfSWtAAxdtcRLotLaEcBn
mC9JYlfD8zVPHR0gCHFAxqd3McCKdmJ1rU4LWK5DAv4uE/+xcsGP5YhAsv34n5id
CQw/DP/t/3J4HFIJZxDXiZrmIXhGs3YgZxXB+H37mlo8KP4/TuOBIRXmhwzTsRgv
Eq8jnoSPhbqpEtJkeiRz3gIQ1eu2eb+GtP55+hMKxVKeaqBn3vdzn6EVOLVrkVCG
k22xIy+BzKEpgwEtkGAl70g2PcmEFtc8dUd/pI2KzmxdeKJL3c/SNmZyTtlQ3s5+
BqNVw+K/8fUbPlQD8hEn+R+/V9tmDKrIZa4vnAXLj47mp1L1J6U5FQ3R3SEVOQVc
8CaR9QrQq0SEyDOWDkSL9FxLt3tq7JIVLNr2UyK9OAU0aka7cbfYWlKYQ3tb/6fq
r0X3F7wiqddiOJeK8P4A0C5k+m7/HDiI1xK80mtzAtC30xr3/hDKSxYUsxcSUe6i
7y8vVQb3oej0B2T+ziqVqLqbrea5rk2IWibczQzwL7GlnA4b59fVkWyeyQVg/9MJ
HdMAPGFN8JuZIWAHjqOrxSvc+t/ggkbgQl6eCY+JJrkymIjt9uP9+/pN+DVAZS/K
39EJGuuY34lsdt8HvvNw52aO3qUusnflMlI2t9qG2uL2SSCNpBcg6TJFZ0V0qtnN
CPtJrXkrSHbfEnunR3LkdE74TKGRJJK8xGXziUhjCkrnK0yLTr3NV5/MgTT+ShnP
Yz3G8i3YyLU+36sfS1hj3BbDJywwtbX9zX4NubwJHa+IiZ++qPkY2KhQJUvQ01bK
1DuJwxWPrwq8Xdq5EuT7CVN+YuoADJMRC7A4ZCtXTcdFCnPEx0Pl+nRAvjE1ewd2
PYHJEOq/9r2gj+WeJVzvw1UXXwVSIEH4YITG8xgC649hZxEF/FhAEdnU2cHG2m7t
Cddl165cKBbDfz94/P+vCfHkkdnVaGiNjiDF2uCFmw/lbCey+N3+wrDUJLxM55KD
1+UNm330iE42r0p0wE8ZRwYZq52rqsFmyv71aw/AfjY9DZoc1XtHZVczYnmo1nn0
mAycMyEzwrM3/pNQ7yElrHU9zYbswifyEepOo85sY7X5rvm/NRTrcywO7XwGZcxZ
2ycWxqvFzq2DY0Q+zPoPZzGsvuLJDHmcLF9UAu+sVS4LgW//qaOEj0m6+mJZZ024
1nrmLedegIN+q+PA/thxQkPshYrqb9EUkRyarjonSeA/w16P3hPdZc5EG87grtqn
7Zj7ycMPsIDsreBciZDA5nSF2kMVquFUXcQ+bI8cXJv735kdQ8bVPx8CqLhsqcR2
Qj83Khdyshh3T6yeK9NCsMbEdXFBjvfL1ZMHdcKLWE9jJ3ALFjZA52ETb4CL2gKB
7wWa3ENllhJb/OUJt723GPqQ4r1OzJrY/QLxKgYrtg+rPFDWcv34GplgRQPgW8L/
NFwZSx6+qgzi6pj65+MiK7JwW48qpTrcbVxQwTqGIegNPZ4MMADRtv+3OE284Wxi
mjjoDhlUYqUcN+I9e+pjssnjydRIn1kDdLmNMFsohtzk2Vp7FXEVyAjT/YiEN/ze
mXmLGap0Yng+RJ9JZ8EVSUsL/qGNh2PFn7OHmAGzKE6Aa6oWVhjhHsI5+CIPsOCO
G+MR613VOVHCw+mY/sVIZL4Gyti419N/wJ5SsXM8EwDLsib8/OgbXxOH+6bCY7De
XXsBp9JV+tpwDBKJagGpnlajgwB0Uq3fDihn22f9YlIgF4/PTjdcmxPPJTtkZ7Kl
xI41zDNWrKxCuRtJLIUYxcVKnjLvd0JRPMWQNgyniLy8vUMhPlw6RiR27o+t9o9x
pmudK3rKuZj9eRCLxS/w/6fridGWXwruLUykGHHYRDfJsu2O3Fv4Qj73wCbvb0RF
1EHcDuoPEy7Y3tsnD1xxAEbAQlBvyhQn2EJTfjsh2k08MmGArL+4iwhI3EJPpsHw
fwTEhcaheBY45BmxlpTfRmKh5MDlkbAq9h5YaxbtlWuoLKANj9KTP7N4SZRM1mA6
aJfCMXrK3ok3oztDZ6SRypjYjYMlXl5vTXPkbZpD+gXeRxnMC6ESAOdK7DtJQQdC
uCXEPr/cwu6EbnL+VF8MCHyKDHnGECQCK+uMSQR/SduUdac7/m7roKtZL+qWoJjf
u/6LAi3T/D31ybmJtARFGshJO3wmh5gsdkxs+Pb1SpBeAaKn89nrzB9mcBEec5uN
CdxzZCweEds5iSxW9LEsot07NC5Ej4Yqywdu2xiBF2HSAKMcBO0F15mQl4GbU1Fj
WXqQaGxjTF3+3ZtIJ+wlXBVTzu8RpGhkX2h3A6PNNcwiyL8SxGQPFFdxpnlMDgIB
USoaYcIsNAcpNtZ28Nx5tnazV0s9xxdxmLnLMhKZUsKnDpN/exJNYrPFUm5kqtGd
ts5QQ0HouBuu00a3scGxDo4t3qJLfS7jd0J0aCHF4iF6BytXrBtylmhCmtupzeIX
jZWktYJGioMV3JYL9OE8Fiy9ynYWig8PRbD9Uwgj//1Z7ncpYKEVVTKEBaqtPZqH
Eq742lyyIl7YNWlWmbbtukoOhTBOSnY6xaEdKRCq+UY=

`pragma protect end_protected
