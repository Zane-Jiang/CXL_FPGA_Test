// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wclurTnIoZjN0lU9vuvA1RH9th9alvBFc+0m1GXNec5VO/m+mZP+AdSLS+/g
mwNiBEp7li4HEXMIfMNgJKD0bU+hv7V1eJ8W0U2UO3DqXHSW9qzvaYIydNpn
CVlxJVR9/AShbAYwpdUBrCV6DQZ8uT2VebQQT4NFrzOxS9mOkkBRuLfFjKt9
Y2Thm/Yyu9zeiEVf8VvCW6im/4garPHeB89LLRBUMta6+/XNx7Ey4GVImvxj
O0qo9oa0CcRA9KHr+NIDzs7w9Gyqa+Uqalo6IbUnFIX9DnmT0wdi6NXpOCX8
ShyjCAC0xc7iKLnTllDK4DYHpf0YnIMd6kRrdjHEsw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MIP4TkQoq444BLpg9abWJCnn5rPGMTFwgB+AlrshR4R3H3JGAe+f48CxKUjQ
VjJu1FyLHJUbPPHCoEBeFTWlcAcdh7/R87O7y64MVWKoXnQH1FKVuDUnxu+7
9BTpdOFgazwef6PdaEVGwe4x5YVKv/xEw+t/zk+kzBAuQhdUk/RMMGvZV+io
zlVZMZxKJvpxJXA97dqaLinolzIYq3MSzNCaBn+2NgE2vwIHueEYyoPS4U30
4xVyQjoNJix7QQJaCWvveXm/hSYgamrenxjopKNJajRAxgqXmGasE/JWayD7
X2ReBrMZSTrXSwu6+2tceyY2stdrcrB+ULTmvjMbuw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n/GYIRNjFJZ9adZr0gw5EJ62t5nPCZ03DDkIiaVlXQuzt7uVdyJGIqTYnuAS
LhXMqNNbD32ZyFpFvGCZGh9133St+IgLO9jd2jqPad0scYmHnHBUwYS8JN5B
Cy97ozeGbq9Yz6pIl3QTFZatAXJrGBRzb5sSwDs7z1yVjkhxJhMvc3dRyCJ8
mRUGdvC6fpKXyzjJes9CulLSPljtFOFphOyWbzkBAkcQSnnCw6g7TMIEqcmL
4KmOJyQiSJhgDzy9+gSR8qh7l0jfnejuxQ8izXwkbsHt8Nx4XuE4T8vrtXyD
d4+ZsyGdx1vza/dpKh7kVNe0drhrzJ9D9h22dhXbeQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
p6T+/9UOsC+ZNTJCLEkcMhaBlO6MUzzzMcCo78PqnbdD5gXVI3yVEPU0Dxhc
jy46D3vWH0Xc4l3nA9w9/AOJUMFzC+VqK1573DMq7xMoWH+YCDqxK7N89w9+
iISN03z0SCeY0spG5Bc19Ak4qknZlZg4rQjGq/1kUOR947SuLRY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
v2htPUzHSAvvcg//Agl2Jz23AOhoJuJ6QuHFlsY0HBJHP6rF6qcAD1OYOSoG
j2IZYxijxKST9OJLwcs+99bftsW/Wk0BK4F8nu0mKNGJEljr3JmFdea9SVTW
kCoYdLuQaebWMuayQmpvtdIRce/2v57tuoWRpr0DyJBfBrLCVLMqFWeu+UtL
lkvM1H3f9ANX+pW3gfIhWkk/JHTzcC3+73eteNKMZ7YW0XsfO+HssFs7+9oD
fEGGph/+Nt6vxO32M72AQaMYAZbzuiE644moFajwcOW54KLpRKSWCDTsNfN1
qgktv8ISIfwKix9PPyI7iUdJOBewPp6z13doUs2IMxOqvEkh+XNuj1AT2+Mn
oRrpcRjV8KBkTqJLF3zr43mvdyXrTnMm0EmTKUcEJRlnSjKpVbV05GExS8cm
2X5aDu+IFSVv9jHvQFzHAHwt8tTGN5hJAPuIn4JD47U7jy2qC78GelSzQrh7
Ne80AKpaxdST3eJZpy6U/EaiLBbVcDS8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NwFKY01F+864MtABAL4NcxH5tTjRgD4ba5t4LJF4HmHAAXpgnVVc3SiyxxtA
ScRjUNKhsoCItQs5/CwevO73HrbYcQGMMO7LRKv35Z+xfXfImukuWQ0ZW2Xe
8s1hxSftPlP8+KxpRJAJfKCRMwa+Vz/S6u8Db638IfqOKwrRNw0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pHJdAaQyi8QYXwLalaBoc7BbfRgkPY+7f1LDjAts7aGgHrraxbVNNH//+Xf4
ZRLkkE+JNWXwM8OM/79SZTC4eVqiAOaaORcfSv2IROlWgdYvWlgwp+OoT3v+
OCiuHxMuZzGcYqxjIDoNrF1/d7fJpYq3zEHXpZDR1EdExQAC8ss=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1280)
`pragma protect data_block
5RFaOur3nHqYHU7yTCEHdN+OC8tRyh+F6s4WZ7+cki2H6jH2+CP6Kvrl31pq
ghZEXfL356n4jICecO2abqMwEWdVrnzsInPe2TO655s8z4J7mq/6xNf2vTwS
5wyjUWcniwvxZcW3yI1PniMPU5FueOAZNwlyWTFGd5H6hdDSSky4zP6DEGdh
A4q2xdHPPsMdVyld7ovhgdZkaORQdP+faY0byi/lcYnM46kcu9LurNNJE10u
LA+pS4M5hPeN5CDm4dCSRiRKCY05uVEov3aWtIavMEhh3E/UDM9r8hp1KefP
y242/wl+fsxTiOU9KS82eNQehgOzo9DJQa0241tK6Ra0ChodYUMRnLY6GEL7
p7OPwIzpdLVSiuw6rogkS5M12wQ+p6GzrjhZ2qE9Uovbll5CNevnp5USvPk1
hagZWebpsFZPmdzL8WsGw5Db9jSmXP7aQyL7/A+zOvTgwLD1N3GLPLsRp+Un
GLeZNd29keifjHvEIN+cTdoyt0SBU7tB/ku7qbJfd5ZYYCO36/sCDzNqJt6E
TTEwlojr9/5VEEOO7zdtr6/WO6k5QApqXeFXp3cGn+Xm9bZKi1X7F9Ks/UzD
oelTuLRD0SEMIe/NG67tuDtMsmNfE/0D9zYkkQCoMYM6NkaD6QWNiJ3d5A/W
nzDLi5j/YFhO8BIEeFQ91TiLx4PaDsZfBvOKoMZ/TUCUUrU/HVn30NJI+eds
KUgSr76b/yyPiH+OjcFO2k6Fkd+JPswWOg2WbNms0ARs/Q0Gkq47hIls3GaB
AMlI9gzyCXXT7qIigjqSUG3HBqsQvzhXdU94uS3axzZ82KwfAFtRvtV8GkOa
9nZtF7l9wehdhE8wu02NQZVnJ53nhddxtr4PDb4OEnI5CisXCxNB0q1x4DCK
TC22jGbRFu9WzXaSESoyZ6i+wi+30ycS55LlE85LGwv6PL30E82IfHaJxdNe
j7WgOg9PpDVpVazcHAEqV5AeMkm7MpCALGQOJcN8b51WgAQ+OhuGyhLWGLAs
ohwn2+BXe7TSYD8RSV4vtQ80B8Qh7tiK+KWiA9ZR0PqGrSOHuQDj4BnorahY
wCh4OHWJRokds+cVkwlAHwmjlGVqOtGwDOwZ2KQSYiumT5CAds7QUZ3L4yIc
PgcHsirEGz1sThejNApHWkbs7CNC36RebRoSxQEZ7KJocm0dxag4NqSdVMqI
MxuYYiovtks8wU02iaOD1T750/ESjnBdQ0V5SMKqabNIkmThuiUfCTolRdqb
ValrX1Hrppu1oISkhsg3z3knXF0w1BVj24AjBCP77L1vG6dNjHVLxQ3sCecw
PPSSBMwMR9tOz1tHdXmWech9SqZkvhBXmK1whsvGLzVGORu50qw2O8lIZyMZ
AG3NdZ7+IWZQGmPgQR0/v1tc8z23i/Dokx4MRFhhwTQdmJwb8Qt9X2QeOryw
r4ctm2cIBzBQ8FY8s0HT7tNoCQPtrSqdyNzYTiBK8KiEcojZfHfMIDzGgUAP
/2yAUHuIFZB0QevTJQnpTS6zF2RYBzKU057DJvg6dlsLE2kSYn34eskCvO7P
L9DPoySJWxH2cMWVVCfyTPxHwfAPmm+9kwEKK7gLl30tsMVIWKVP5GtHLRk/
7EUFgBOJh2YfNKEkLvTCjRI8km4ccsJJZYQIi7yGWk+qdJrdPfNp6yM5YQQm
Oish132TU083jtDs2lz0ncJhfmk=

`pragma protect end_protected
