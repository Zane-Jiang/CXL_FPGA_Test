// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rS7CLgdiXlWCZKsxKavnNFjIs1IVhwPfItSqJvJLLbwnRrZ6uFn/8AP/skDew3pLVI4tQ1V8xrL3
5W42sYYB/BGaWMAYsFd4Gd8ZgXIjGR1VrU8hydKHxWny1q21C7P2rkONJ69/tw6n52CzTyKQprvU
OzxtyerTcKykJrpLmF6hyumcQVz4t2VbPmJ/rGB50Ga7sJ+7tbuhowZX+xhdk/wp/Dwrygc/QGDG
EJ6HYqw2q6w05QMKDvJLZaAhTB8Q3887M2EfrT4Npmmx0+1D87aIKsXVj2NEWq/mJlrEtrxWBrPf
waRYvaFadCxeVNOQ0baVkMlCbYC13EZROHaLdw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
2bZWfRn3ATLUCE9Ym2Yp96hrtQZ0VyBUx2TOrFtuHB/Wm+SYq93ZQDKVQKOu9H4b8hx2kEK2PJtr
mrq5q0osOOU9tZLbekX/2wAFvzPQ0nDVh6kW/WbaA56QZ1/CaqfsQXhq9dnswgNmLI+VuA0YgfMl
+cZg6ZDFDpEuU38tPpsSxBwbGMTVlzdNMxww8Ms781T+DXgueeWjaN2fl1Y0sWObaaITqnpCSawG
KX9Tvz43uU/iTnoIb0U/WTstuu4exspJ/feQaxOU/6MAQrecZel3ko8Vmw29vafs+IupGCeQ2q+u
U7HBmyy0xvkQbF/gdAYM0U69e8WYhuM4kjtG/0VQyrSn8/HFqvnVpd7Z4VMqORelTAjlKRgN/rGA
0STiRfeWhUlRI7rqVo7LkBsA4zERpIWcC5LswwyllZGkNApZiHswHNu3rV5mGUwYpp4G7fZsIvX8
HjeN2s64x9/g2OZZaYMtoB0ODw/B5myf7hRJi0QNbE0b/RqfAmtO7fdZ2iDB5YUedmRSeAhsf8EH
eP/pK2eTkKxl00ZttyCmYWP9BJNwvCWZ0amM/XV+x6YVsyfE6YfA/67X1cWu660HkfQnedpObVOY
CyT7tYS06QCm+jCF1CtaD0GeXNt0JZbTAt+H3Et8F4SAj+vXOU1wpic4xC8WjObY8Nx4iQLTqn68
Cxf+KxRKQpKKY8Dl4qQcHJfpZHqUuHKKS0YyIYUgPs0d+/nPt+ayx9ygBKU55bwudDZR2os8h0Uv
JeAH6YAW2r0jbV1CV+NcmaU+hTytrp7HRmcu61PXmVYyknOVo1ZmIF+pljqdawc09uLlbY6qr/rF
+8x+XG/nVxlA3j2epAbJWBeui3BZFdXnJGvcrxXil4LMev2Ijv8rnYR06L3dBvRtnx/cNSAtSXV2
KQZSxzEYzDvXGSfsn76KF24ykAWmUTJ+vHEuSHhpmkk/6X337h43g/zQh7GE7SEmfvqZ5SWF9/BX
rxtpkh5WsWOJFYmcYCbtwpCnaGVJ5TCRLEVfCqnzEp95A1A/QW+PIEgFkAgpe4Jdr2JqGM4YB7Rj
0k2XUQUlW6wRTHXkYSdRgQKM/+gzG9L95oHuquVDbxzPbYULogtbvwMOlJ/uneERhmmi+WQBiuJq
T4WwvHLxZ4FHWSQvDSIkKXSKYGbw6VTGeKLOZrXK0RL25WNkgIeMV+qAGgXN8Hn1K6xyibtSd13K
6wbieWx3UXg4L49c8XVpCA8frUiuvYBk+WypgdPclPmhodITETj0yXqpo33adz+GVNVbrdpbyzZ8
7M0tY4cxu6NMxeOY0NB2wevoKTQdUJEX+JEY1+T0PHpF57VOw8cYXSFXsUzZaY6r28vdPkrMtgfG
09xIzGBIAnN2fbnDx1aI8CPttvrTUoJjw6YScFtMgE92etSox8qPhpMMLKq91YBtFocRYpMEg3ec
pXEa1InFe+jfVpsS7J1fPDD69zjF2alA3VbX0lKOLg4dQp22LPT2yD4Wfz7wfCim87+QsYV5cdqR
KMMUKf26JJ7Wb9pUj1mjQSZE9m1USFsZK9L9zUnIvpi9/M3bTy1rzqJSIt+I/hCK5SC1OIAHjRsU
MMf7ClE1Z7iUlKGR7nzv0F6juye2oNyDLNR+EBBKgStzbesmdPtO0QgZCIsyBkHh/f6HE4IjRoZn
4udI150sjARMyYxhlHW0vImTRBOyUsLQfDdsjA778iCo6fLvcfeUGylK8ktQoPs5Zszupq88Om0g
ISEUbVWTTT0ZbxV1f3uumFGOfXwDsg+KlMP9ilx7sOc1S4lo5h2LNnmrKUc4EM2uAZPucojrknnu
l31qcDjIWyacMGIss0NgarJ7WnH/h22tlM0dEQYdgE0gbr/T4Ff1nJfxcRichtsa6a6gHTLT4MAD
fl5eX1xqNMaogrL4SHt5ViueS1q3JmaL6ZA98C8g3VQn2q8QOtlksL58CwbO55KeNq9VGRjTfux9
2rnFiCApLVUrMYi2tKwWr3d3vFrnD2m2nUKSsd0bu6aBOtiJ51zi6tml2ZGfvTOIbvtojy2Mluc/
5t0vl0gLsgD9CcQ1HUE1qTE4SaSUFd8cSBla3GOIK4TdU89bPcB77kRqct3Nms8OFxfOGDfAMeHd
IcsCZjpp2GKh6Qhb/5Viwvf5PQMbFnRgpP7HTC2p99Maz5gZ6l1x7Ox9i9/b6hHthomS+Z5BehdO
+RBs4DxpDw/4tYXRPAKaQHVf+7c+rTO9xa40Hwq2tnck4oGcNYE5gdqF59RsrsLCVBkIMiW9D7Hu
RlPLU4r11cywRAHQHUKSZAO5La7ZFfmBSMIbVYUCkh/LBqLI1YZasrUBsbQvj5QO6MIbc2La2wsU
4r4v1Wikc1QgiY4iQQoKhePNyrxyBtc/8aSQFL0wrbNS7dzdzudWAC4QvYJDAjxh2JHiprGkKYKa
+TeWEZXbLF9RFpPoe3A9v82cDP5Ias9OWCHQiJREVsPhWR+Od0/ZUOvnr/RpROEONL+5+8TlRM4X
8l+fhjAIhw80qfzGELRPCe2O+EHJF3J6/nZJ7MZXSJW6zmATs7kxjcLDJwcdK5sWZrmVOoNAER9N
BpNmd44hdLd6u9TYjzXuaDU1sehPbuiBcpfR9KKr1hsekCZ0olfeZjhMo7VIfaiWFP9jmoGF0sR1
O6saIsO5CJUparFyEgH8TwYXB9FsUdjOV/M31tJ3nWMbOVtikPTCdgbSgNG5gxOP83EcQBOQG4WG
CFeibM765OX/01BUniA7hkjalTGhGWSoqn6T2+Iyr4oqVdrKo/LJGBqHaFJ7nxQ4NmFp/usbwO1G
eHZrYJaZR2Os8VkYZRUspxDkXzNJ98qzJohuiOdkcFA9fdBHfX3pOcVCtFtJyCWN1fSUguKAyevW
NaNHUt5X/o5hWCRn7G/oiTCfowt5C35rWChyC6FHEeMiIZ0z3+n8Xz784mYoxyTojalO7g53PUKB
ROpKCFvf9CIdyzDmEQ9JiB8u2cGG8c2YenBkEOWfXp+wY7EnZ3/cbiPjN9qz6A23HGlZjKBKX+4Y
ZXZfxgKy+2juLv8kd7HWDu5ApGRZi3FObf5vp6yRubd9MW5+GTxmRBTo6iLhrPN0xMg4KO0Vsm7A
7DX0CITcOJgVuPlmcNZo4+CoAyfQUWmRB2tVL5CuMqzmKiqDw68jVvoB322Y88mRzhe7FkDnQU6I
qLG6242pJovsHYMxAO6rNLYUXOrudHnsx9MpSruu1eNRYzOu3sAEvdDfifk+Dfqu4xlDhEpF/ayn
pU8/dyA1kwBDhUBH9BfLOE7j4GD5/NX0QlJha6e8SO4uZvlKBmEG2B/oj3DuloXsLkmiRiVugXMp
wvlwgDofvjqdPBMV8PKs53siMT7dYUMIoAvvpgZ7mluFNAJN9ZzHau/ssKsRrMpTLYUw7O44faEq
ByDbvdWWl/2M/lrOyzSPX0ZAP+xQOHt1/PzADxY8kVq+AtD/YSYvIuItpCYsMolHFkBlHqSQaApU
xcjJfIJyYxibZfR2Xn3caBj2f+2cmZH0o9us3rh0UzZF9lJ7xEKtEcwc+Kb2opTal4fvoz4Yx0EF
qiqXNY+LJfEcubXphUfoQT/eESRPpOKhKyYXr/UwMlIjViv43mzcGDCIH19izkvoh3uvUJ8gZqf8
VXHAZ+f+sOI8NUHCbndpLAJigJhsHsxZwjUGMiQZKAgboPdEpDZb07FcoIotjxirhFQvU6R/VAjJ
ZN5zmp/QCL+u5zCc2iCMJWSNGcVAnbmZwjrEKxVQGpIaY21lu93OBTsTt3g9e+xhfT4zp9qsLpdz
5O/aX5k4ANEZU2ZVbmm11y/tciGQN47lawTpjp+XE7BQVGRj/GlP+nqoGx/XjGkf43gqWYMkk6tV
8IBsNdNAsdZ0xKDvZ0iGJQtSIYJb4SIH1B8HBwBqFfZcHwI+ZjTZ9UjmXrOH7gi0ibReDIbhar4g
TeOGL9uwxbfcr748CGg/+Lyu8LDLi1L0scaRO+nL7DhpqqcV0BoEO7PbhkjuGY3IRLvzyh8GANYt
9v4FTWDGFOgfIP7rJji9UBKrLg5Czo2KusmyD9K6b1JmedyWpRcRNsQKHEuxqyChZvHprafksJR6
XjBwqR7P93YNJTF0RzWpq9PzZdrFLt4UCvipwOqH7AnIAdeGW7r+HZQfKv9so+2UTZNltP1x50S/
sAszeNKfP91UMERNRcWaIULGEJmWQx4z5dWK8NP5CTN6iMzo7IeFkSN3RhTekF5010srJJWy9VyX
Zw08pFdbt7tFUwQ0KOyXhAxcGmktpQ8duyRtOoXIGXuz1bq3Lf0bPe7bTA0iMtpe9nNtJzVoDviQ
jMTzjmXNJWcUYEoyUY9rQZDT3gMH20getMCLWwnyvhB3ljcc3yQugOI4QRZ5jIzZ/3e19UHYGClk
VdAn+DJC4wfeHCp4umlW0FYOvIhjnH72iYTXhYyOQz0o8XY0Y8SopWe/8ZvYYYR6TsTNz1j0OhT9
IfNLjjdrAjpA8MlGZQujBLqW3OHH6++Dk5IBN3BcgLo9UlriDRkio5ddGBGyM5RpoG2Q4d9/MWXX
Um0EoXG+rcVGRys1qbVfRV9VGWe3abhrss8vai5ldVf6jaKkpozJcl9A3ZJaNmqoDmfA/gNDkMdy
7kSegzqpqBk16RJ+mFCNdafnIi7WnIXLf3+cU2zrF6Hvolx/srlu3GomPorVtAu3oC1oKRHga9kz
ImL7d8dKyOrAqiQAGix6tV4yBWwJXSlC2H6H5QdoitDV1yNzW7bZG38YPBvU6EEhULGDlNDwO46e
ITg+hrFhVBluiWQYQOyzGa9Ggv3wWYu/XOePTavTfjrYJ3074Apl0YRgT9b/sk33/9K+Ri+hbzvb
tnxMGYzEodSSU/t3rXYMgYwVF6xhQW3zEBoWvdYGv/rPOrsFe7gg3l1LBqCu9E0X9+LJ8NSEaKai
qo5ejMWScuoMA21TgHvv4U/ZCz8h7+CcvvRsUYOA0ZRUhjTk5dCgbfL07yd2V0ezRqPY5iiGKQYM
fy3Zxnl+wVHPAJUSgOD+0s7npRnFiEMA5Ibooh4ScvtrQ+w1OuGZUI+3QIUXU5E/9mu19YPBGW4O
MjXZmv3Yt25ofeY7RFGnpCHkRsr+1vfvy97LLZttkrMGMOXrBjIFsXuAJu4ZrNyl3ShgnwO3ZBYB
IF6jbfuz7E3hZERMfsuI7qv+vFZ85KdnrJDwJPa2nLA/vDknkK3ls5IMn56Axd9SA4fbd6niEVjm
fQh1gXKAm48keSnuO36fhjmvewLB7nbUvqreFS5pq0vtxqTKeC7PeMSrGh5CSXAmFpS4bo98wWvU
tY7pFDuz3vLvAu8a1xOBXCirmw8ZjWDU3Ndp0hbj3lT97AGkc7ZouAAoECLzpxoWss/QIm46Bw28
bb/4qWJ/ujVGffk/MDg1GB60Z1lW3L23VH5Zg4xukpRKTw8l06kifw1IIU6BHgJbLHyR9sODgFJp
IVzoXyaneT6PMdVzvdINFWPB1KsgLtwHUJkVDIEEc2Sb9BjnC4ZZiWZ8GRMUzGnY7Mgbg875fn+e
07VOCwlvZk6ntqedhmCLW1AHk1tV0px8y4yjoCVDd8VrvvKLJwv5FE71TIIvSv8n9NMxUYjzULOs
I7WSXOOMu19Iv4eIV8FtUWeXzLZEdeK06HYsbYWuDL78gCJtoXrqlFFWsw4Soo6mn/uP6ZD35fwr
FhRkCUCitBxKwdiYVg0xy34wnY5hzJTUzHnclGj1bUT9jt5wx+c8tt39tvS40nMxmMuezojmcuz5
oZ/SNyNmi1aS1l0kx8QgmTJFQyyV4B4PH3HFna8VYJX9U79h9DDpsdt/S1ReqaePa3BK7XRt1BUe
Ds/T09axhSmu/+4M2Ca4rwjKAAQJoiyl2My+xqsfAWGVYajW1RlVtb9139mMb1rySm7GKvxaaOa0
mD9NRCZoW6qKIuDckQq2Ysnaoa9OewP7sAbuXtGjIzxxvvHPQjzYbcHZ1wWDitTY1l34ua3hIMZ5
5oOBCwSFFH/WIyZEgf97WgjVEBwK+YCLUFwtUl0aNEuPK+bttdrlhPy204vhOR6vYyAW9MQHry12
ItQ26zMInkOBxfNBTJIBQKWDvwo4U6Q6Bk2hj7IYTeviA99HrzZCxm2MMl3tGZ5h8F40YUrOvsE0
BrekDSpQ4U2FN8964Yl2d/R28UN1WfqRldF0J85RBP5pxDte7xEt1BHq+HyC1QA+2PTElJi8fUjA
Mvj7ZqxBLtooWjUswHBhLAf1t8s+giGlINFUdxNdmDemc9/GHyft0r9Z3fFSACFrabFAW/pKk+uO
nhEOzNShXeuicj/AkaLbTE1XsJNuSPoY+x/vHpIH5qhTlGpTL0H2vYekylP1r5zLu7w41a3lYKWP
WtQVnwNVML8bEh9Z472kO8ptwTX3VCOPZo1J/KtVBfvjSZ2mNdnI+Lmp5wCluH6ZEUFX24etUXcS
uPzpqFdnVsz60OdlMlIkxBywdaanx8kl6Zr7cjiOWuyAJKMJzdfuOfavtwEydDcC9wLbh6r3uUgG
fkxski18qAdNadqW79ZEHUbQqvmdvT048dXC8T7JVOtBXB9YlltsEGb7xtKSMOq79A5fkVDlyh3n
g5N/bylXlqxQ4h9c9ql42u4SZgRzxTRsOtqqUK0fW6Cx3Ga7TbfWthqE1h4zAqam9Zvh9tTKXouH
E/hqkaxtHQtQwkZTgekfRRH/2srcqyCMuyhb/0NkLth5JL+8Zb1OLER5b4mxsDBftFmrvvUvsiHm
AGPiO14NjA/LNazejzingi/VBMzzIWN83LywoERic5Ls+EZXkWEZDIXt7/Huj633V7n0qDLBoOr7
LLtdsTodSwwTyh+98LZO9caOsHuhp4cfTakE5NWpJWnb/VSUnjjK+7omkQwECaowKkoJwu7x6UeZ
OXeJkwVEx9RrClj/snuU/k20qe5dTjVhSU+o8l+5x6en6np2RsH+1fCJwrqCdthnF3Na0uLvdysy
DhdhFwGNgl3y8G2F7wT2i43RUZMN4/bS36oR18bIHgElN8O+Jf1sMv0wJ4vqAEC65VIWi4sYFvs2
qjnTL4C90pCDgjLSltZJVXgqtHJs5sd20V2lrp/FJS0/0TFOlP+dl+C3K+J22Mal4PSYAkzB4Zvk
K3J9cBWvnhq3TQuieOsizDI6E9Uq1J4Di2LTaq8EagnPj4dDfPCckSwvsqo9e8Vo26fwHwt6XTs9
4b7/QWHMaf9EIslYyc9gfAnuHIlP5ab1LDby8WuPE4a1jqAV6sIg9KucKs35uuIRxBXlQ2fVY4xJ
A48MBu+Gkuj4OUpmya5XQzyqDkWGOQmwjVZtxJWSChPdo20T2fvo4ilxg18XV82ln5BiKvk1gtXz
593DansrqZ5GflejiqaS3/kEAP0VJDXR4gzrEp731p8TtYy9vq0dwUOEbu46e1wrebDpHXkmRYPe
DLfMgT/bbv5nigTpBSEhOpmyn1J7j9V1qtrBgAjAO7T+j/WSoeH9RTP75kJZmtUPCqJHM+Gz0Xo7
DLbS/dZ+DCDKpDS9jnBysJ7a7XpUWoEGPmozM2RoGemzLlllygIGuvCU7FYOp4NYP7EBRxhd0UAC
Ys5LqmgCyGjPQAilI3kvXQ9huzJpQ3z29H140R75uAhtawtfpH2bgZwppXjhLsNbu0SRgds0QT3I
dLSaGaXSkcqvmaJzrI6wIHwzGUQJCxuBD/xWOZWekedg3IBtevXictjEYiphzpKizHmMr6AMPK3G
FEGoQeEjUtGTCuVF/5afpBbs/orPOdwSayIv4wiCDxtZfDAM9hgnBCzfXs6mygu/0ZVPBS2cvVge
mdUe94yMIOrjByFYk77PNfrvuzIyHsK7wuMK4Dg0CvK3I4OLWNSXZaKBAapVuuAJsp+XRQIbrt3n
67ORH73xeTgyOS2+wOnhQEWYgqeYqfX3qPIYZkxdzrIjkCDsnHNflVZuL6FvWeADngYY1X6buXaC
wz3wsqemgP4SRM8fjUoGIhfoZSGnvh+i8kyEPWOGKJfHUYatKoYNwyeDy+1Les414MpmlVgeZFd+
mWtQmrmw7jF5igXI6wivgogbdBVJG3Eu5t46etxwCIxFdXm6tq1YwpevgxWa9c190fOrWHWxjvzT
FsMyvVg0uKJpoQtp2IOUcw2FVH2lLS1JHaQVwGq+CsrDQPvqVhrYwk4NSNANJDAVrn6W3/j4Y94U
ozGAS0/EAvVYN/L6B249RYzA6UI2yXFWnnMMo6cQVPKKQIVBWJOOCkHU98XMqsRyVIq1R1t7NeJO
NsoMUezQhcwDtFBUtMMF2IFJsubhwkDY8/BXQlYfytDKyvzC/XpBN/JhyiMzS2ZEOI75sz2/ZF4L
uUT4FqElPpHu1/gIdJOdMrjj272Y0f5nYmUFWq1GIRBaPRm98heEMgYIBmcRjCw+mx0O0MNMs0CP
ww4UMNXwxLhZunmYQ8QiYj2CRC+xgYNkDOYiCpFjd68G+Wkw2VqiAX+iFdGb6neIQbfW61gujepD
mqKsk8ioqtI16lAokQWaCBGnUHyjBJYFZtqvcD8FmCgq6n1+NtYGnzvBYGe2EH/Ls7t0yOPuDQqu
vRwdLQm3UDwCKq9DqsP/P1frProOJUD5Rk0gIbJAC21pbR8NHPjiqH1TjDNgz0T4QE97FhGdqSqR
tssbxbCdtxELKwmmWNhiLxl8VJIAbKbhwaDdz1wF8082w39Ps6YKkTOy3jZwjqO8lTrK+qT/fLOm
bIc/ga7BlhJtHCIZWlwWnq5xcNtYZxEWSurzekxcpY1mRXG96Mh9x6coBKv4uFmSTi0TC76FuyQb
tSigQUTAllrzHGdv7MSXNFmZMgA5U1HIHSXYOxNMTaVl7jyKhxWczKhvRHP0W6EeJ4uwWVLOL6rX
n65eVKeXLrojopM2dpXRV3f6CYq3MppOdVKpvpEbEm2CoQvR56TeM13zTi/yMoN/UwT0KDH0Vq4J
KJ9MD7uPO9dqJprlY6FSgy7lNbrM07zhR7IlOvABNTUiDYofZljAPny3xxBzUw0bPbCB9BHAhuTZ
Ek01ycIPirO+4482t9ODLi+37TRAsoHUlykqXlP83jJSRrldcwh7jvCj6ziVCm0Qw8ej3YVQmxtf
dGgoKm2YCrUlBksaZLr2cmJFVpjsKaAQywF8ZefXPwUv/Ef4j+L6s/rMpQ6KGM6DIq3cXaNuf1HW
Qyn8A3RvyKk9qCuK7RXM/d08OInbNNPRFVK3G3TH5AZfA2rB/AqLINilE+EhlWTVcB6fCuSSAsNm
OzSmaZRyXyPrlTErJCKp6CojLOTAMC3wKOMmNT7BpgFf/QkmbzC4ZEYczpOLm8mj5ZnrN3GJTETX
H8xzb55Y0GeSK+WtueSp3F9n6MlHdeqVwDo67gdkRR3gt2LRgIHWj5+/ElAAnX9ZX4vmCi5AUr6p
/pKwhvFrF1+SpCPyNZi1t21229HFZ4DyKQ436kVfuIspzv1KSGQRV15n87ZgVNacHQWvwZ35X1jo
Y6uJ78XSk4yMQ2Xdz8XdIKo3aiTn1duO58EBx9p0bmViqMKDOSuClsxdgzcszlcIaQnej6Cg/Y+p
WKZZGQI4WLwNyQYv0LpqIX0nMBpEMJcISgrjJeLVgnPDElTLT+3SJntx76xtraCjThmdUuOxNZX9
cINWfHVg+a2wOxFXi/130BcMEs2aTlYXPNit6Zg38smzuKYqidSv5Y50vyojfDuiPJJ6+uao/Phh
QAJJqv6sCBSeTxPikqbC2Gnh9J8fLu6g29PjG8foozGvQmzmoRfP60Af7df33gBrENeZXX8UEWGN
/qxqA2Ki5NRGqLpmmSwaMWj/ZGwgzA0sZFuHbNPgj8AF3kZ5xTPksQGUBGYI7YBdzT1vohSuJila
z4b/C4HnVWFvpro/UfQ5zookhF6SVeyw+nY8g/vpRPvUUhy68ChAnZ+j1t9N+yu+6F7FNNxKZO3v
oAMBrg0DhsxSndhjJmwUgweGy4MsSPcxTgjWvG3tJkpodNGx04k74v3L9UckSsDK8aU4HZazMH7o
m0Chl5CH2OyLUf9jU5GiKLyOCZ+rN8IXtPek51OEmhNmurMxftBxGRbh/BzaAya6rp3I0fV/G1YB
CkfwQ7WClh4fZK37IP3xXtCuBd611wWcX2BAHnVH2iGUMQjS3xI7P9s3VObM9zre137RoOZlsOef
Kgai4IO2Tt0xHVT1YwcLeTyBchTkkLeWG+ylGlwErgcwruvLdn/CEL51o6sUFBFgYq2fKNNwJJ+W
b6D9cq44d5bnBm27V4XYYZYmy0guVA4MalAEU9DzaS+etGvcIgYp1uB2UYGSDRTzcXZXWbew8yyT
HYjX/g93fIcUg4rs7xSn02D4jVakiXxxfYU1j/FjyaKpefwBMvkYPOAyWbfHQCrD3WP/gq1OiiVU
4xx+bsmVIszQlyesV91Y5AwmeEQgKZd2jx4+wtbBXpbJ450jC1M2EUZypuKPMk1x0bXbD/qUslk8
tQmfD56sVHeISUsI5ehJkSKDozNotyyp7sL0PyG95Bvu9BrRenbn5N0SS2FgsjTo6GBWZ2VifkPG
ubNWE6X9CBXGyOkSl2fJyD7Zh98rI+/WFNxA9BJpwxLNzSabhQmY9LcR6voE6vSO8dxvUljv8Gm/
P/Xhcvf0lv/qfcsNhThGiagw9QWR92031hlJL2N8qIWw+Waa+UMP+SF0T0kpBQBplZO7DmoqVD8i
zrXUN5HQrviZJqs5Hqb4+nDSG/2ZyLZ7i41H26eXr9LLi0sAHz5VeO6K0sJN1KyJtNaod2cWrlrh
oXOUZKUyYNFONiBQUgljIi+1BzJRp+lV+4T+zs2OuSjOtTrUKRR1jKHnUj9Kh0MkNPA9HlboekVF
yfLxgHyCbJ61IrFmvziD2frcdGaWrGlMenvWrGewQBkFSVq4RA7+yY1fza+/xt/LVlV/wjYtOwYb
1oJtxVfQEhlwP9RCHSXopiykr8juUQAgGbZO1eyRcgn1YtMoVROOnwGWIuHJbeUH8PVfSjKp69d6
Kpz83Yf4E1Hx/aj19BSxe+xs3FsOuGT79TIvwdXDXbpfKOfqvJJ7DFHfJCAcizeU8Fl4zS35Y+zn
Gn8lf/Xasbrr0XbRdZ4NlYX+GnwKIteO7bgZYNb7GbrTctvijuOAWCXkpcz1IpZ9VnlPYLFHge+P
nU0l94/85ZH/xENqrSKSaxECDiUosiRcZvn0izkf9pKTRUMShNQDaTdH2UYXueunmYJrpVihFykm
qi6s3rJCTFUcXdbmictiLHE762HkVsqOy8zD6p4xatTaKKaRQe432x/AZKCzmXVG9MxgFE1JF4ne
+j6l
`pragma protect end_protected
