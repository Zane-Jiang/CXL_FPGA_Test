// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
su1ZPzONMBiT+YYwK4qPtZXZsDhrG60aCxANVqr6iMmMX0Fpz+vfH/T6IfTLKwaN
a0+cjh3BgxIrnlUXusrauP3O+sYzx84b/X8l2NMDN1uGeNJ4OhJUuRWGHCTgO24h
NPox/NbXB/RcqNvl+5ZS9kMGRt4nAfYySgeJVch/vb0jpNOcPH54IA==
//pragma protect end_key_block
//pragma protect digest_block
kd/S16IgkI4w3m6JB34Cu1BifHw=
//pragma protect end_digest_block
//pragma protect data_block
RGh7PXOvHh8brDr/LE9RNiVkEyHMRq7GFnqo6MfKvmVVuKVWF8mA3Xkm3JlddLHa
EsiY4GA5F5d5b+ZrZ5RlBrA8zR6N1lDmFdVAFo9+Z6qZXPhFlMdFR6jm01mBWkaV
sMl7MdeYvpYb9Hog1Sny7sHDTq9H3ryfBgMnAbizVuNlUWv1tWGBXJYOSQ/xfDPw
AeGlE8hIcOkB9j9uti+wzzTR7yCJdvjzBll8Yrlj5LaFwWE4rGRBE07+2q1HITit
hnjyaEQy2tk5LMwpH5ONey625wQDKj3ioJBzpqXHrYur+5v0uniWXycr9ROaQAfn
IJOaCuJ+16Vo1JDel0gkCsjPuGib5Ggy66H11+B0Cn3d83Aac8tW5l789lp2bbdo
tTzOaoXiJ9kMu0GhBUB64gnYWoxDRZr+pgcDX7xxZwMLTWog6co7M5lF6AshTSdC
hcIUtulMxVuztUc5RTYzNZbaTH+3CzE49udxp30nu7R1uQFi4ZLd+pXjVbGpfX4D
2To+tNp202YlvVQVKupqC4+826QbGbl3/+QKn1mdvCfdPCuVZ2HU9hBY4ZIa+GlC
2oPUP7wTkJk2hYzLJTI2qArosi6/vBQZaLlWzaALLhor1/FnNi9eGvNuGrrx1uX8
jEbzsgLn/f9iedwB/7ZVbMyW60fH9IH9jpCYTa5CNPuhgKAEL39khHtOmGNJc8GU
SD2/bW7wDKruQZyBpLLGoufOqYWIWM840z8wkvMzwKxGE/Zz5SDXNIF5XtI7BD9e
3qW2zAa6ENTdG2ZGeG3rA3vGf75KFZ0ZMTZdtwjxCnpJRf0PMVhNzHfEHFT1be0d
VKnLdljWDrdklKT/VIWcJbKvGRwga021MHgX4sMFqHec5VeWP4EG2INjwl28ejte
AUgRaDUA9/5e61M0pDlgYUWhzM3q+7YD3qkAfpCXSg3P0oHdNWhqAIeEQ0yWT7zo
97L38AERugcitOotNTWHcqyZpTY19BAkPDWUthWrf9VgnsibbuDzteFwyXqQg1CO
rACV3Fiem5e3XmdSDXO836j2Xngty2G3+JJYMgd9uKQ9JM2SfAhZ1MxN1tzRv9OK
Fa3aTxjk8LpJENbz7AujBBgc6KY7GUCbAenXKCthmjt8QICM6ndXMeO9JzI7KUcX
0rQS1yzSObHpSkR9qvw/M93Gorw8TGPw+bT3dvvf2kPxIhYkEx+QDwf+KLL7DcGC
8+x3kht6lDpnUvD6hkADljAe67eOnKhp6BNZbk618hVm5fNfURTsQsrXA0LwsicU
PEDk1DqrEIxMLM4T3dYS2jj9QoZYDw5R/qf+rUg8XYEvaFkHLStR7hR+e4PSDSCE
CG2/occuvkcWhQLJXO40N9ZzJ+mQVIJxu6UGaUc0+DBmdfWFdp0oY/7lnhtTHzLK
t+Kz+k+/G83jD8ndLd/CSXcMs+cXWQXKc5kSrYLgD/RONHQny5YWWcVHYpPMA+F2
QIAocxf9bnXXIZGKli3GS5mdiNkAD9hCWNOZJoosP0wNibFwVFcQFf0Li0+TZEDX
q4UD06MLb2ZrRHvZ3CMfZQCDX9FeEiK/VituuhXbEZLqfNkkYolSXzuLBvunGAHu
Dpj7vQ5dWiQucVj1EsAckVbrBhvNM06TtQdibnw+KtkqeyxXJrC04tAFdtaljE1I
o/KZWCNcyO5EIxNb/Sy0VgW6VWm/b4pmmONUqBNJdyo6GC4RfHwFXxsVqxTX1ngm
XqIHRx0S5hZVm/JM9jHquHZ5FRf6EL+1QQdQ4CMFAzlCSJXezR1uIwmt6Gwiv/Jp
YWDWqQB95Vrn+3ji3POUjIfESt2mJMMtXwtnwI0npnR/320qoskmaWiEGRhWKgNW
GFi3JTwF7FWVpQWM6dzvy/vvFLTEKMov260mXta/y9KlNFvNfvJzQr5455X5ukHu
BrbDokf0XlkEaRQEvL2XfwcMsSFCDAM4usc8t4DoYj/Q/AqwGj/IxWqpvechFgO1
d5MUEi+BLLFBkdTarkYPaOXTkWlJv0QROgYNW9lWDzDJDi2LpqG7xKfar2kaI1OC
RIPTWPZ6964+Xp2marThH/yn5LTzgIctp+jDi7nPeXcb4SHjQbL0kGkGHDwdAjhG
HTkgT9g4AWPH8txVoLVY5xe2ddZP9dPrFv+I7aqe6qmKTzukecM6+x69Hwh/5tta
zrvvHEf0P9jmysVpZY8Ttpx/kUY/U3Wu2vqrcC8jLXAPS+jJQN1dakMXziaYUKDB
+Nscd4GafS5gXCfbd6/XZXK3mw9Y5x6qbM+nFoBz1cccAzUtJSPn9H+9Ppx9Mlfh
N5E/hn/97p6Fo5UICBb+eaqJ0xvi9k6tuwflmtH+hN9pk82GuXUWGsTVQGzJ1Bx9
fxtC5gPapRqxNFQcRc40UXhz2/Et/VB9smG1GDPGuOnAFleumeXUy9Keh1io4eiS
nVHPHk1sEEOR4YNIbiPKqz5+ioxKmyMrwNgxqqNgwFJsHrVG5iFDZ4e03sAjuWDw
RNDZ/BXZkMIgQLqFVoitQG1Tk+f2hUpaGAa3a4ETBD+U+hOIBHBeSa+DI/JtDj9b
geWb7201/vcnUgnQtLetmyiw3o9MR5esPhynAaiztIQi9ji9W/GDpYjfBMF1DxXV
gi1/LFg0N6PL+9WmXDfhiYH6XpzZnMZ8ky0RWRMOpRLpZ1XSK0OiAJMmCflKXuwN
ZdD09ehCK6tHwRc7YyOv1eK4ERyput6vjZeoTVCCXTDDFPrwzLRLesFFG6vljckJ
CVtyMorAvkJnXLsNEvn1iVopTBWVW3sSP2ZnHzPG7WowlpQ2n19Yj1k8F+RfgXY+
OidP9KQ2tXYKD1c80zlf7X3hvjJmztc1mm6901J1yiTy48nGGBlk/LYk1C6HG/5E
n7p4Rc17BSSQ13O2K6+tLANXa9U/yNZFAhwy92DbHhH+toe83Q2YTWqnvWRTTBBS
D5fqbFPQt/humOn/U600TJVJ5vmqyVqTXUBsw9tSCGBvEp+meEJKHhG04RX7tjRD
E8gbR7ubXnaAEuRX6qXa+Clg2IUr5P4tqGneAxDyMfsRdAkuee5jQSQbPWnyFPna
4B4Ycnb8mIpGg/yKOMSptxWC8gF6C5EbSuQgQdfkfQs89tmCSYsO+C0a6bC2YBoq
4iawk64N4N/kvISsb7DeH6djaeZCWTPzzST+1o0OAT4oui9aMdGm/pvrYR7bdaqK
vtmfqFI8rU8m9nOIUwDtXhR/WaljUNPMuTOcjLha+LD62UnEWGcaWhImH4JgiR9w
x4ShH1tR5I5moyEBFec7ewQydS6j9kzQYlwDShBj8WcfsgK6AvsIEG70i9cLxGXx
r447CwufWwk5mzMXYgaj/fHe3LLQh5j3RFPH4SfAJUO5FPLJa53ecziyoSVpS81z
ovkv+pW54l/Q5c/VwMSf3D4DuJ1iGv3ZCrU0rtMri5xNJFUJOn3gAH2d4GazDsYd
HSmQmRGXfE+N4oqzrTuzu+UoGq0SDtdMz2+0ijt91lXbmzZ8NOmkMjcEOMBs7qBN
sB/C26cM+bQTyqr/r43rWXCZqqlrrxRjdINNlBhFQIFLLx0lWnhTixeBjfL1Di6L
n3YxhUCkcpyOtLBn9xeV4npmvZtscUKeaHmfSVh8KQ4ryL9gAQn3VaID4lUdA8W1
Ta9GJhwmrWL/ENwcBg6Dysj6VTcwlrZtFJAv7h9dTwTPBSUcPleJ5rZqdPK858X3
T2p3Dgai8e5WxZQ60QhzIM4c8IiSnhNxQE8mRVKJozmMIumDL5WlsNIINdNuxtZd
5+pqzmJ/q17ahg0QaPHUyVnFYLGasOre1z9iMt3T5qON4FDg5KOeGJXCD30ByDsG
NENMo0S4zgwwmpIC2j3va7qEaF41Bki3xy0UIz5jtp1PhiQs7EbUFklMHwcFb2kW
znSCdU6y7k/xiAOl/9ir5+j6nHCr6hd7GV0nO7Ef8cSdhj7i19k/nsT8i2YE7Gqo
ZmetDp1Zbjh9pOvNh16HeRFrwmOdSboRaBvMI7FiHOLKhKGQZisQsFs4Tgw1TptE
3sWGMj7RQdz+ofEVO7L9pUSTHzkaKTeXtaG59uIfcKWzZO0whxxquFYKxeW2MrYy
joYi8VFIDEaSfYGHD7Sc3buuXnxzuvDt+rqfn6ice05XbDcUzyKGK1WfwdqQkjYs
eJCeisWmQIjmaxa3Y4EVHgG0TF416ccz1D/WnIm8t5Vy9RuhOLu2rQJ8aaoOw+dk
JJH8J0u0rfqkf+wpmClwxM7nJ4xTO+3mbBM7y3b9PXid/gGehEasQ3OffD09lC53
F6AKF3GerrYZz7hrvIxZ6BkHJK/Zo6oGhFlBxIKpJvjyTRP1nKC3dZtuq4ldZ+KS
q6wvNw4J4DKzYNA/VF2KzXAzIvblbotERMR3HV9YiOvCzkhs3d6ab04rJar7Af8l
CiRM+rJkMEIfXiMK4wOhPEcdduTiFXTAMhRjK2HrvcmnteXI1L0MU0ekuip6DE0n
ieHbuihOt06ZsvOTbi2cOH/9YxLrzqL4WmbJvDI4xN0zUkGEmYMi23hdHVZzvry0
YRXLQvBtwr0TyVnErY3AyDKGx5woZeoI/T5z/+UU9Jbd7GhZngFwoTvr4RmQIfLC
BuofYPjojiUNKQGo2UZymONzVlieQcoVqGLkyKFLDYno7qMbozwb86juMqG9JTtM
4mCoAxnvRUy5sruRNH47cmKMm5xjH6qIg+1LoIrLePxSFCOI6TCNJfWHdlECPuMZ
xz6RXPArKO2orOXQXHy908stVoipCeeSgldLP69QuVdB7Z67HGIhRSzFgNaeCLXF
Js+nhmOWAlCltlVtVGERigvWTw8nwbWz1WV1ukAV/OPU23zjwzmXoZ5lH15nICMe
xqhD6kWc4Lbm5OWuRP/Xa5gcU1u0iQlMLyzlYscg6SNyd47weOPu9cVS5EfWq8F+
4v9E6ZkiL3fr554Ny5dy+ohE3qHuNLuxQNnOHhdkEasFWTajjqxWNgf+yT7vV4m8
Jyc25wsZhwGKcTl48WzE2I0w3uUgk22CFktA6QlFNpWuns3czSnUR9C24m24LO6O
UkTvb0HNdsECql+cM9l8TatBFKCY3vEdZ+xyRag9jYitVM1IUQkyTGZAgbFexmLv
XrNUqmPLWdyz6JCvNQzMA/qgBkWW7wgpgLrmpQ+D6ZlnLM/7j9QA37PyhWwbUc83
C2ctbGQ6IYJctaRHGHoJaGekav8yzjfyQHh2gC4RoSmRBm7EBOsd+5Nmy+a77sO7
VSzexiUrkT8iJibobgxDJrvKbp2si8VKP6FWY93ti9mpRzlWx8FD1FL+sHRMsphg
6Op/V4KVeszk0A9IV35k1NN76IzhE7H2V8Fity7IIsHeNYfiBMU24u+fXA2T4lJf
6jyvi8IfSUFtyR2RIXQOpuUTnQxkXtmEUy0+AIYz9+XygvGCk7AI44aMgIW3kObJ
jcb6dIcJynI3rxCE3JDlmUf89NU43NvnAFpSbHyzXxOfMWd6CFNa8e2MloScZd34
TTQqQBn4QJQ1QEojWjyuksvmnrr03pUBIGC5SEYq4Q9tjuDHvjn37hh4++5YF2yI
t5t4XCzDhVuPM23bNstUqwmceBG1tig3qjUQaWq2is3NpXNOBydc840C/63gVthk
tVOfOZcwTo2pKqksqXauJzCPplW/uQXAuKFrNhDnrGnU0AY2X497UYN+LPVDYHMl
UiU2zOh8A7kywtHkhjhxm20AJ96Ixb5de5DsFwKSy4uuH86hdIWnQWBGLShuH35m
YCyVW8Vzvgi4B83A55Bb5fNidR7vt+teRyKddFOsvxbsGJQ6eKYJH+VsIy55yHO4
Glz/T0ohIWY+0iQzEz7dG+XI8sXjk1XVL8HEAVC23RJOupDrhzwlBhTiJTjbI8ZJ
QiPu75psi0w3r91MlETf/bkqgcN5G6R5YLq7a3G7Ow7PporbfSIOFnJyyn6DQG6p
w5RjljPc6Ut3PmxadqsrDStpjkR0MdETUhfIjfvs4oiHadPIc2zGcA6qqqycKuea
ZoeqDIS/0y1vDt0qsbypDVvwEWu2FvW9Spmklml/IwXvlUbeqEkTLsf01TbLaw9G
yI/xKhGf+ku9R9ONlnAn5GzT87VhxRphJa4wdrQai72hwpLdTct2y2M0uRQFudoq
W0kYFdbHldyW+KAPwtvd7ibHM+sblbAJr9NiEvGyn/Si0zgbSxGoB8Iq5HgMidCx
ceR0WufbGp0h3CaGG1Zcs3oR+ZN7zaRSGOFukdWJj/Q7G6wIxEZfRRkVCvsxGB97
3z9qu9mxb3E+FWy5DfYW0Qr+NeOTuP1/eHeQE7S21+iJgMDbqm36oFTjObqzc1Kz
UZdAUYXPzMB/W+hEGH+84Q/ecW2pSD2l3Sl0ougyb/EiPCsGcZNsCthv6l7xk24F
0W0w3Wi1dHE7oBVKq56RW3ZjHGtBvpsTDqZj9v4XYnEhoI6bj3yeUYt43KTIzBJ/
JEGPY0wnkFBvwvpN/Z8ayMOtix7OgxCaYKgLHN4XDy/4a04oThldsfrEWsaPSum8
6KG6dh/viknexauaZI08qiHFjOvNOYUChPu8VC8BBY+a+zGhrHLcZii1JDkPTIfW
IiDRw9EItPq1Oi8r0x2ZB9gVU+hhJILMJq5xs43iyz6+DugRYjSapGb2/7ke1ZLA
eiKG4reoIJ2+FQ7KGFw0JJK2DgStQiU7y9kgVdiJGY6MgDzjuqW1zxlfHY0oWn0E
OHb7WChYfsYdMJb1o5oIR1Vu9+juq3oROKLbeSYcvp8eLfmemvQSJRsD6MZEGq9b
isLSEgmcEs0m1cu6UC/jvBHwNlNVuHF6GNweEWXIN2zRuldj9m5dsTUJcW3VQXc7
tlEemCqR0YnMFet54eb5wNGJvVTG1EbXt/viHQaZbsyKSYY5EOm35H+Mxxizb/rK
/g/1Ru8x0Dhp49ml+KvXsIZzKuImmlTajz1GnIkD+xu1QwsUboFwBxwCrg2/rTXr
sGw0x4gTIWuQD/5XOOcWdIbURtEsRYNTXMnkIo+i7YX3ydGCqhPrbp2EatiCYNPI
ZFb+6mprBqH3pg/nI6FzAejf8sqA0AB/0vaDUvRcy+XVPSmoBCTaaWcNF81syQb9
Qe+Y65zgi8QvX5La77vVt0yWCz8DyRBbkFq2m08U6PwCu4sMppyqa4phuVRJeSi6
L+rxYFRdstwT2dMWKcy8O1Ai4q+if34o+9JmHLFZ3TtSX0W0vykfRjAfXs8iEeBl
R6qcnVsZojFD6SF2A+AqmJVdNzsoPyBAbFDvvTk//w/Wss8kD0Xl4rPWEvNay9Bz
7nhTY71dAyBDHXfegcrg4Tq0sdkLdSo8ZepD5xGRqKSoFl/mbAzuihqKy2YZITpA
mMvFT42vPSKgKUj5LMFShW6uh9mSadZkvZfXAY4rjb7JPspx5b8UQPQ6b8dMWKLh
+HXhV/8LFgwaUQ4MvPlqoSif50eokA0uopdhXYUrEo8d4C1FQJkTI81LI5feiyWN
5pmBhoT2XWHHzy3+jEtEAg0shoh2dQPNts6JJg9c0qfB7H3rLVZ9YmQv+UwDaY3Q
uiLawe2/8cD8amHOlxgQC9hyquypbTEfjkppAp4jHXjnmyj43vAI8PWF0LLprz7V
74DGkGenO9YXVsgtrkDJ5wayOLZrTXoRpSjLZ8tZ/WFxx5ajC94i9Q7+sFUuTyp2
XyxrEze+eGA8m6iYq9OavdyLYwn5dCFRcT5lSIcziABo7dyHoImoL469y84/o5EL
R5JzuMFG+GpWrsFyim8wv7tvDXL1Frwhwgx27yRej6N05NDG/w4JwNKtSfVEMsso
IF2rl7m9gmQYxBYpyj/0HfxnuE5XcKa/fo51O/S5bEI2OkHFeBxMOpaWn8IqJJ2+
XB4shbyXPyofy/T51E6Ic/1SB1Pzva0cF9A02jFb3WxIn+o5cOlg7ZEZt0O5w017
5yZzpoS2odbwEzlmo+TV98ohljeBg/t42OWYtfEiTQufiADPK1yuLRIjhOyyQFzh
9YN2kkLWwdly5GfMxCBnv4era+oeNk08YAC+TTM9opNZnk5EiilmhCYtuF3ids/Z
iAw+h/CDEWi5o90QeLVm4SOYJydAva4UjzcG7yFEonavEGhcDuCYCWRPR02fLSBN
FlGeZ9mT1ddf/d1m9FF6h8mmUg5DDX2jIWjVZYAetxocMZah0dqo1si+pEWiuhK/
giUFrPLyCaXZuGHu20H1TiOETnB8egA0C2XcnpS8U9dngYlbObwl8br8soiO180t
n92HgGoWLqiu9W5GK9o58Zfv4qSr7ugi0PFlpeb6+kRsl8NMak69YGge8yjCioIj
QMBstsyYxquPpWUMuiUTkZodb3Pedfx99ApCFOHwvE5etvKCGpl21kCa7hSWksz5
Ymzsg3YrhNF6FJSa6u/LpVakqRlzuT5UuSn6YT1urZiB5p5kyGFzpQ1Y2YyQYsha
MZfR3iYg2vPbdZjc2CWZLaqziayzeq3e6v0USeg7u9thB5JauEMGU3hvjZHLRzUN
AWEdWefi+80OK01g6s8xACyWmUnu5ALyE0Hn9oVKNU/XRsXLT9rycZoarOoma4GT
4KkVdJr4UKheCcdRbPFz5+pTnghQ9d4JPeJ6f52kUd9f6W0dy/ig3b88JVisBKr+
87v7EVe9102irRaa2CxH6c3MJGUSDJ9nHL2RJcPcVeng2h5c9afnbmJiCgfD07sg
1xzqv+LM+R8ecs88g5YYDpot6gh+RNnGXXil8xkjBDHgwzMjQRPJStSovojnN/5f
vdE+jQ2N3lFyNLZp1XqmpqBUXTa8jydbY7lKNIBarSnABYBLIxHoiDucIanSBZS+
+s9Mh0NuFffQRYavZr++JMVNqERxYku5Ysu0QBRQHZvkub5WMJMpfTpx1sDqV3E2
h/vuse1dgyNh9SS+dBQaAfl4AphumrATt64g2Ax5xaD1rwqq4nllSzk7eQ5s3Sdo
+uTEJpwpfRhmyY/QroruW+0ZE5oTF96v8pYbz3OCqXnW6qiQsJ7zfqw7NA1uvhfP
p4T8QUkUx7xXMLp+afqfXUGGBvywwVAGckQcc5N2hO6MD3LEA8rGQIEYxqMXH3Vf
DafCjKe24VhiE1xcxGss4AM6DdpiuVa9FgcagAL07GkDateZ9HV7iuwC3w1wruzX
WnCrbn7vLAfZCMK5LvYV6XMzv9s/kcvFSszVsLat1rOy4JOMZDxaDKeXtZbUleZI
J6yA36WUz/R5K5DRA3DbgUc7PeORk9L1HJ3YJpc8jCLvNCsNMTmuQHmwqok3K8FY
38Wq4oJ0fs3mi4/l2l+zaNQElVx1V+XGE5h1qre1Rmht6IRSzawWTFTVK9og/DoJ
yRWkia5rFGqleSGsuCmp69KNQKh+sHKDRnaCr3pKxVPEmHXe8u1jKtbBRaUoOJS6
fUgRkkyTNN1aVmvqGjIN9z0/7EjHcmAd/HixY0mRzPpVxrCyKlQpPHAav8r8epOr
pt0nnoMzjfHxs1N66v9C41+zqDGHwvhzniu2/QxqmhYTbrSvv/FpSPABj4QTrN35
kjJbnBTNMIJIhSnk7W6rZH9NORrqeVPjFVndE8PttAwsI7nVxHCQwGl9qUb+jZ9i
sHvPA0rnhJT2M9YqB0m8oh0lWvIzVrTz7LUIxxs5TuoEfVN1Ae6smP7m/fUd35f+
b0LOfRX//yMGGQlY09VIe9gVAfGBHCq2BdnomTnko5EELvJOdnOeyQCUeeLrf8BK
YBjlrWV0r2Gason+YA9rHwDDVXfsrQYP5xUxiMKtQaIbH0BIhXIEqSL0Wa/jhE7I
TFs/VgUIKz0h1t8cNXMuzDduEBcaXhUVHgVqERHmQFCmnI4Bl2Mx2Eo0VoyGeSmU
3oCfDLxZU5IgezGFQ64KmrqcArn6hOBp8eKCtWCX0QHSp6J+aR1Rrc/cLmelBWJX
l1PTK5dtQT5qiQDKqLx+1S1yBFEz+ogZUttTryK+Xsun1pYJnJzHQa/UfBhtA3iY
fXknUBtgZg3TIVVaUkEyE/DiBaSGr7C4SYU0QktyF2s2WE8STJ+FB00zdP84Zcqz
oIJMkdEAGXXufJqMm4yPeb8AX/Ph9QABxf/blm6WQ1RQJcLbCP1PSJSweklA7RkV
Of2rakn4xlUP1e0MzOMYDzyiN/cSYhaw0ULF1S7bViozzRvp+MXjNa2AtLY0nNk6
3zmOJ4osSq3SoRUisQS1bCxrEvd2K520vOmsLleBQ6AHSRktV8UMgFTAespkyThc
HHtLn9EUWQOtBq+LSrJ/BtbUSWRI/rMh2eUKm5KwWEjupbBvXpPTVrcRl0i06VJO
T+n5rEQvQzhAbrMaP3qihAZkeX2p9r+snWcRnH5El2tSJ8h671oHbMxsgxqR8G7d
x0Nk1cNjp7IJGwT8K62ANhSgVZzOzUOik6CyFCVGMdOV6SsC0aUMqmyPCCFGXMKY
/0KVId4YJrqgGQiDbD5IHounALBvY7F91EPIpZfxPmYoPvzyognDNmTyMjpbB9Hz
k+2s1lNBcIIdPCSB3orslvSiDPQDcDEkCfhJ970a0jIAFDbq4MxbqppPr1/b93uG
Gmbr4fjMRtVG2B/PxCVTKU8Bnexy/ylH6wN9iRVxd5n84gbIwpyBXbru5CVhu5W1
IPdqUBVcw1YOusDjkUKSB/1w0vOqLdNMNhR2Tz6SSDM4RMyx9fV68yrJk2BRNNq/
ZbacNq9JSvbLcZZxIlkKvRRBNfMB2Ccc9OD2kNrjbWmeHkddGmWacLgXype5WmjO
L8asQz0UDvjP2FfHFFZmHXyKR3a/Fk3z/4GkSPMK6iJTiy/l+XB3vjD9rE4BYFC6
DbnsTmK7qIkJ78bCnBc+ot+QaT3UblwJdJ/JqqXuGo5FQWiUNQRZ3RzGzn19HA8P
xCVNgq0GLWDO6umWl5lvaLGuDGO+MqXEQ9y7PvUKk2j4c4edeHJRlDdUWfk/8FZr
zCKserBoAIw0PWE8BhX0BgserNh4ezBjvGYN3QvgldywpipEurnqOVKpvwnZgHPT
rBuCbk3VfFlinnu/9D5RE1kVAAxITP9T3W4pX+h1jcMdaNb1PPzUH2wF6B49w9tM
YSuFcI2iRS4SInyNmFFhBrJ8dytOIxYVbLVhkCFcoKlxMjkS4S9oyqESz6SwkbuF
dd6WIjOVLlXMVEfVjEtueIWQjuA9YeGt8HdF4Bp45H73s2qy8wiPu4LwcKyJww1D
irHDNtXhGf772AeeCQO3NNGBaOxnl7vdIusny0YKOsP3rVLI5mvVlk7l6VEFPn6I
48DZe+tPI4fVuluRwRwxFPgJNJMFmJvSRh4jubS6GVXKR0VwMpFdGNtf7AKiVjvc
RrvSzArwIU89QUms/6t5Ctt3cKQ1bRjyz2QR2cRTC8zvQunYXhelU4PiHFqevolP
kflKjaq4jdRCvjC2EsKCjyaq2rHHRiFeEHFgfF1x0CrCbd1Q5F5Grig6sJjFQq31
+MpdxIccXLlxi9sywze10endlqXOfa9LNF6ifscZ1nSKATrCHIbDH3WSA1s+iLGi
bPaPvKHAWRLdw/H0J+PrwVKBUg914cJofY8pWhCCcclKCaIvmaCZpcCCkewsmEGX
ENI83SruPd7WncWdgui5GDnkYSdPojdM0JtzBwlhjyVzrXqzOSyYYhGkxrNs6yNi
C4lJSLdBpyR3ZsmR7LA7x7W5bHPLtoeNfowa+Jjrl/0=
//pragma protect end_data_block
//pragma protect digest_block
MlksiaC+z1L9s3kdgzpodUq/WbE=
//pragma protect end_digest_block
//pragma protect end_protected
