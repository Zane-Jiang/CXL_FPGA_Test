// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Y+RtKOfJ9h8W9r6bXhtOLFs+YNdealtKffRbjOl1UA1ErMtGv4ca7lMCy7f+lVEv
GHAs/Md8RBl5bOOehoO85ou9MK9W4Hd0zk9Y7kFBZd+oZ89DFDL8ySl2ZSxtTkGM
lZ6/R6IRBLrVhFr0cPmqq7N/hqCzL0s94U1WsxIRwGk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 44848 )
`pragma protect data_block
QPMkbb58FDfZmckHfg7yPBMQoXkaKFhdmF3B++jXs+svkWo/K7LpNePhW6KV/4sK
Ya1m/XidbbwVes+7FnAFYFopNrxiBYzBH/JPs78xlPXhiYAhcatnQ2GKFea1Xze9
fZKZLYgZ3oiXzixitIw2ule9I4xOicYtOT3b3vbTF+iHEFc3RaPD51qtkAG5cpNf
RDOJgg+tEJb85s+zdJ7I6OD73f+6n1qQBC68HerkoUcehZ/p6t+rAbg9N/jooKnc
V+5BifrDYZHmUvnW/nylNyIhjdX5YMb16M2vAM+b79EF0bYWtSurGkn3El4u7FwD
0uZUDCwGiXe/4defisNQt1QUhbdqEbAXj45dhMr4z7Rj/gfnz0JJlZCoM5fMmUsT
mcRJvn8rmXQVrSkEiSdtEn+88UYZ/bXNtMsme1aF3pPLdLAC+PV0xYyXB1KU6HPw
frAYjiFDJkczcAIVZ7xkHghxQ9yr8yGVICUUhbM45w8LG1TSqSwzSAMcwwaPdjLB
+mhiFyl1Rz3vE4TOBF+xY5uRhvWHcGUfza1IRWH8Kc3H7hjhE9seO04jCcOZA79P
w7OoTqfngA4NrCkoxO5wjV58C8qZzL4AMvbOko8+9sank7Q7/CvDsAb6TnLrRZ9t
kx1kxZ0PA4vYFa9wjqJLWWeFd5fU2RgqGUFmOBZiCqf+f0bnI22M3QXoUDMCW3vV
/HkQILpCLdfszVksRaTr5g/rWk/aZeQwUykTlLdn7N3IQjDAfL90V34qcYNNl9UB
BUxOby3OtresjjzHyJGFMgwS8K4CTYtrYOOG9wtiR9NNi2c9yR/HyLiIN9H7iJ8C
jEcWhC3socQ+QXir6sEWRAWbfw2qA8KaMWM8VJKkCudCWWWz1Kib01zTeuqO95w2
6h579VBSzpS8LPNOC2CdY8fNSLlwbrddOOVMjAK7vEp8HZNCkaoGtcIBylYBrCiQ
HvafSLt19nb4eEQkV8oak0E5gOPDZcVlTLa32uwuqaWAAx92/lFasIBkij2cn/dP
FnKKYLWduNtbExvhfURdpYSWUK230zeOQA93gqt5fkREQyG9bV6QtRoe6nn2z39e
KEpavXi5Aq1lt2LT/K74sLaMPm1fYmP7wNjrcFQ7jLSw2xlZXm1WYfpFVwQLlqTa
3eNqRSGeICfOlWwk3kYUw+skdvrZwBzfbu9FzoBxsJ3xRb+FfZf5UIHIh17juEnH
HjqTowzDi6hZmfUB7cqGMV1I6Tp9gFdaE6OCx6lrz9wwSUcxfCpuo838ByvLvF5F
YGvV6s8jbKgmTQtjbVIi0kG6sk9JgYEJkcYQcJq5PNO/2OtkJ05ldr0k4qYKUcfG
b3gszFFyuv7lr7MGkSgmL76rntCcjqp8T2UyNKqkkxxd87+BJjlfrM7t2CEDBgxq
qE22TwVyeOOubCRugkiztuomYWUAHl9BFsgZdU1DdIiRe/bMuK+rsTlLOwTIw2Jv
7gbDf5ExHRr5tpH1Lh8a2IhLb0o0P72Tf5AIVMKtGeL/teCpDebCSoikcSa7Mhl+
+j4cOtGV7kfDUgzTAybTZ6GvMEDyl8HT2tbUfOkPtfP0lcgCqdhs+h9UT80C8IpD
47kW/WDWSrvOmlOtxpyuwFVrXgA5z4KigTwK0IdN0niLzaF02NQFWvrt5i1+L/Cw
B9yUjbHlm5wSJ/S5VNDHBBY4xhRzQ5ThF2yzuBO0hdEO9KEoUkXITOaWLxf/KP/G
ykd1pnTk5d2If96jj2++W7Yfxd+XxWograGQqP/p66MfE3xpaBG7O2aWyqw+tXXj
B1VKuYgT7kwkWgADUDwVZP9Z1257E2rLPk2I/os2wZwWQA0K4cVnu41qkCf7hPQE
P2z8AAqZabQDXNysOe3IYEhdYMor4FVCzmFs+VuvHiyk+AtVByDSqO+gXvHZmatp
Xh55YNxEf6UdRjcHJbCqIriTsPf0J2WrxYrfyRMnNf74ERadKyMMq2ZMK+wsm2wB
wnLgkaAkZcsL9GjoR/epOhWS/yhR+x+YzQZdSwxGT9pujOTEAd87vQSuTfDZo6j5
OuYp+H7RCnO47Ovz4w+2nQSvkkaNWDRo29YdPU5B0iyxEfqQavWG01ee7N0EJneU
iciIerKs/DMTn9zoccA2TQtpjq72BSZWY79LTsvo6CwD1YCRv5dFL627k1+h6PxI
L6FObmI6W+AKtNLlpchs75QZLo+MGbFOwtCT65+huL6vivCfuBvdDTTvcPq7ZLTf
MZ/vu7kKbVwVXKTZHgzMdONDUmR9D87pg/kXrrOWGlcMxQ/aWuJXvvY1rp7eZEMf
DO/NdsSBwrbh05kPVe8+JMg/JQEdGx+/ibwIqHAj9n04om3mSECOJak3jq98TqHz
2HFVaXOW94OQx5OBFgWvesfXM9VAMASFjD4o9j/5Cj/D9Y6nSqpAsg8lmt8KeVi4
EtsBL2IeL7VbpNrQacFszyIEjGKgQmaIu1M6z/VofRv6zEx1GiOL8lsTyFzlniRM
vavSZQqvT3SVbLIFxIpGDMZ8dd0e56js3VAHQ0b7K4iJ1cLl5nBiFvV2IzgaR0Un
RZzsf200KfIkfa1VmAVbiJLWhNTJwy01Gd9P4gfDGO6+zoySkYjVWwAc62fpBKZv
tuM9iBOXi3Kgyu8TCtgW2C6vWB2YKCsKXZHcISTMTwwAORFA36LUNTYXqv7jjTJh
JNBYNjauJBsxVvHKs1apvtjidFQ/Azbbxeq6Mh/A3Tz4nm8HnJBeG2QGWOwkcx9x
XhWYBvM/aqOfsVAXEIcbHYSYeBxSi6c4PhuAQM0b0DHSzMO9ajND0UE68Foap6Lp
2coKyQcpZpA7B5lnuVUQc/0hHnjNTdBFEyp4wXsk92zFO2REGklsWOHb3p5i7IHM
xzSxuV+V4Su74R7EUnn+2kAHNgTAEq4mrD3pgztgMNodZl5+zeElXdsuXRlLZmJg
6OPVnoePVBGhsQD62XhsNK17i+f9j5F6g8iuocchIvNW2nbTDE+nyZGeLfZWaFK9
qy7+QibzmYQ/a2TLpXDWMAsBn+n2uC2mRDK8ZiCiGF0JDIAQi4AyfL6I355g9+ql
BfU2Hb+MVb99uFJKO+JOxRS0nB25OFahBAaNBh43ESFQX2B8Bh6w7WhaUmLP0h7j
6G49xrATD0uet0nYD4oEnSDFziFgerw2qI4kJByt883UwYsfUjSHPt5WsxN5uIuS
SnSbFUwWNCw8cURwOaEyYqSLfCdKsNbnPnAAPRGMJmq0qOpd+cCUY1oRQeIUk/UI
jml3Tx6pkGBGgoNvVtkJ8sNaDj4qbJotZVPrY5DDUCu0ADMLmhRDD/vcBLjSNqFs
CnGSta7kGOtG84fITYp1+eYlQAX3nQa2JgnTrtcJ9KFHr5oEZtN3HHR1LZntJJ53
7VfcKsVi7AE0aDYYs1hoJYRlk9VF+F2eSV3fYX92zKY8OWCNRsCdPt4v2k9F0U9H
yn/ReEjrig9xGeREQfLFB/grxeatoMS5MAa6YOHvYa8onae8tixlm11g6rz66ghO
scizZRa4OuDijobzqAuw+WsvUZX+986Se0zbCOZ3m1Aux23Rfr2TvnK9QaX+mrGA
1FoE9vsLnMi+JtRUZDvBQTJlNXbu0LSSlBeGyo7Hvrcf50WpEfHSqDvbRivp1Q0z
K5EGtRH+xhu6QJSTf1ryOCZlLAgWUsHxl+z0mNhCtna/YEeBwk1hExLYI9hB5bOz
WrJagr68vLBW9FjH24hka+K90TnY/+OYgwdaVPesZg4jgS18oj8cuZBwejvenqPk
sIaDYpkcYtn+HXqRpQc5SZlVG4RdKPkiWifeV7y9z2L0LJgdFyTol62zm8qWdhsx
8EM9UemfFV7Rko3DH0AXCZXeXMcaAf6x9ZiFEk1BnyLPZFpvLfluVxocdBy1u4TV
LJbhE2Z3jD7fhbA30tLJ4s/LxXpgMaOZ2DJZvgGmUADI3HyL34XWhv8Sywl6YbVs
AqvsLumkhHqcDWWFEdH8tR1V/+qIn2Q4uiDKlJ4WwbkG2ddJ0wMcBxcspsCoeR0d
2IQTSbDqFPgttbgAFf9hnGotiWH9srX8kFmlVdJ7k9R30W3akYgsWh0cLDv47jz/
NKA63hjgNJxhnotSrvk4d/Y+kKPq337zGdyTTKxdA77uaZM++J6/mrbXSuOCkMoF
SF5J674697hZIVRmtezKl0V186I2ZXa2NJuY7xMXIz/JsM3IvppE5KjV++OQSsSB
Va6vPghaXs3gCeFTDNdcmIx+4jmABwedUjBSljy5NTcxZSf8h3Vyns/sL8WYQQAp
VdSMjOPyc86r9DOJJH4G8gytdfGQUrg8qqjNtFMthQzo8nUF1LDMLMvxHzpBI4hN
Gt4cz7PiwgHw2wWM4MYINJokojus1BFKhDmfs8+RDV2JKpWiZFrmr+Edmyxqn1kY
90XSr4MAfvO8qsVbQDWsYmu79e5vMdi1zVaVWcQB+ueXSbe/UvGyc53BeIZV/ufP
Ls7wnXWpEV+8vejlLEdDwLZiQIEbqaD/tQQ7APjfkST0n9DoqYzM9eM5norazia5
HNZ2xzRSDh0WOgEM4SVqtIocsg+Z8g0L52WWts7QGQBIGlAw1rfmJ9RfC8kegY4j
1MkVaGYOcTR514PUxzpFhOei254gV1xHvt4+BqAvOzvZOmIEvNbcX0Lh1BhpIqfv
iW4UVNdiJ0khXThfhPgtEB15Z6KeV2V00KgeVwRCFnwqZmQSD/x2iblLy8OaLGjV
V3jHO/B/lAlzKR8z8Xbl7b0kB5mo0JpOv7xB0oc5wvIdlLrdVANBPTIjTLdo6Coc
bOICXv1CqG59HFFx+vygbcNAUC8r4JrDywm8XmhEpDhIJGnNAAKLjLpRsdlJgrCz
7P2Y6WwnAPaps//w3LB1u+Ete2Q2uaEuGFgGpYlkTRmcQUCCFek+/jNb65myqTVZ
wgeQPuUGQG1XvYq7/A6aFOSDLWB7MCe0OOtJmuWO5AW4M/nGmHZ02iqR3dRXoO/P
KtKv2MvVxAnTzuuixpf/AhkplcpN04FRG79CeWDV5s0SRBzytnO6c9RcEnvjEQOs
tazYn4TqkcuKGA+vS4Docqqblk8rYEDEnPPmpxckCMS5L2Yq6lolxJvGtyI4cdFJ
K63AC8/julvm0W3nkb7eM90JCntbc8ynZhw2IaFBebIRg1pNUmhwVgshdpE70y5U
+8xnC5bnvs/5dcpju+n404GW5AQaYF7WuL/LNtzGcN0Mtevt5IrHTpAKOc6D9Lpy
9UOU7B9uZcRqNmCKeI3bJeRysRnKD9iFUugK8MP4XZ3OQua+FLrV12oRo/cuJrV4
81U+mAlrKKHixMBCJNoHXLVvWoKgQjQ/+dUH6rHISQ6B0VIrI+EGbRcOCD48vt50
6eOWZdRzHjt8jMT45E+LVpJJ5TKDRZzK6qI+OBbW6ok4bTpVZaSL7zr5jANcESlP
Fvlm6U4mYDIeX85NLnMFbQYn5oQqb/ZrI5Nl7aPbDB+VroMBYIpfPkNpjJgJj2Iy
vcXdeDHKY8Q8iBsrt+xCh+JlEhtQnkEgTbE/8DO9bpYjYaLUDol5m0POV8jgYGgQ
7TwMBsXZ3fqbSpHiW8lp9wwTYws1zU/yknQ/tUcnpywi9stgU7EoAA3bi4jW8O+p
ZJEHZdVCqG6crVG+CqRTPHfCLXIKjOTv9PNivwVB1gvM7Ib1NzjnCe25nPU/HFru
KLnZAIdBhUa/L6kknRFRJLKbDub+LWGIFVAdTYwt6oN9pyEzqDLskSlBk+Rx1DlK
B6EapXxMi/clg8nDcKHHH9eoNtnuYIAA4q1JY41DBeXL/MJLqjIL6jbYQXWYZxjf
s9PXP1jMSLXP8CU15PUzHG4r4P1S7vwq5vHMkZXiMTZNYEp0icD7PvirkIxmcjwX
JIvNdah1NwhpTAwL5FqF0Wj7DIHy/ywvZwsWphxpLNvF9IhjwZMp7+jKHrGR7M5s
2WOuT+Ddu+Nx2s08sSeJ8ZZ9GdShd86Mq7rJTbFLVdgFr8tu3Ub2u3Do5H/4bGrb
UTD4Zo5ODBNkQWrlCiOSfylzP6+hy2Q5RYoje5DAHLujpMURegMLD+wkpwtOeqDw
takjIC2J/AGKCbSB99r/SwXuQAAcFTJ4dPmSOXj7KdRj45kCrBRapHbyaMYJaHst
cbfeugX7Mi7rQDHVEE0+vSTF7U9F8STpvDYmpvOtpF09mxd6WTgFYTyEFMAP4Qtw
g/y8454WJHwJ5bgUNLdfy4KPRWC5W7zPTPAX95XoFO/JAD9d2Gcf1PC0qvlpQlg7
zJ0fWuNxOhEoTasA+kMytYEM0eVSsLLjThao4FQBWiCcxu+PEnM+uSSRqxQyKEWm
0Va4JZXLFmhRGLaHQrF2sCl/Zzv+HAU5qnQG4+eh4G3yEjpkS7wbapYBowC231dZ
Jn5etL13JP+Okaoqku38w2GNIROM3ZC0EOAdBF7ZYGp5D0q++CS8XUAjF13L70hK
lwKVv1cn3tUxbhHMYjI3ch65iCIAUZtNQAf3dZoCr3j8YoAvYhkrQDeIAEHYAbQj
NqbCvBr2HWlB6g+/+YIEmUqQBtDo7C+VtSsDejY2eUQB/USqEI2y/nwhvFz3OrlG
H90MMI8d08L54pGtLhqOV9NIqQoi+PMBkERoHJvoWnLhmouEg+hdPuKIu4phh7SA
fWj+tp0L1MYlSTTnocThM/ttTtCUkydqw/0ZSKAf1wwD3HgkMfO3CppYoXj+DnEY
xeyXU8CPCoH/gqTvy13kEXn5+40FRKGa6WF3EVz3JSCQorZxELzetcnNKzrS8RQ8
+3ovltKRQCFpUcSjFNsCUdFI65Q7XjxxQ1H4qHujnKlALbdfvYMZAuKg5hmFOjIA
wKRLZHzmqacyBESm+7+5A5SGg3XaTRk0nBOkCatNoTjXukknaehdnKYRLybqQzVI
3BmiMMib4y+zM1qMXTK2aKF2wSkKPVv/kimXlbLuCaQPfgLSUEAT+gkXUtXxd4gK
MEDWxzy6NtRfkraRJbPaQVOiV+Gt9HPgSAMlxrpWX9g/5KbWuuyRgOnfaxooQyuP
xJQGKdEHV9GW3eraRHqFPwMF51TKO+nIJ/8wab0zz5/42rfieYjjsUIubLN/2Qeq
hECTZ0kADxCgVE529UhDjnYz+tOrOOYTnl+sT9FpwwDFMV33HsnL9nRMFWn++p1B
09eIzlW6spb5T6iQ2nQqkiVCsK84aQQ/PHsZips9jynodgwe86gTYR/+YTGKfh0f
YnrjOkwowXxRBli0uRNiggbK1wfOM51gckWA6eOa370adC2Ejj3/wEBLT33VP8yB
/bKdUYm7zcbuCebtFRgfWT1O1YYmD8vc4k2YX8kumoophgp4oEd4CpXyC6jGR0wE
RkbBrPB+USHHL5sMM9H3DkwTzFiQgTJxXM1DqvWcE0ZD6de0mgZGDQHdlGqH2bEb
JVd8PtJNU08TOH1leYXIJgXpDwIXnwJmKGDnGZDR0vaRptDGTD2vLImsLBJF+w5p
7qVIjdijSjTD+CaOKM/rMoB/XI98v5liavP9HivPZNipQ+z5shMSFsOblL2ZMhq/
ASV0jkBjEXYMYZJ5s2YeyH3sOWM0M09/GPSTEr85KlHEdMggm2taryl0ctRGj3Zn
libYfcAE/HZBFDu2i6sS1diJyt/0cNLcka8GE66TXO44IrJyy06inkm6FrQI6pBU
NgPfg9aavv8hAwqrQLEyJh5hhKZLFrRnJSxpK+5MbF8aPzi4PgwHePPE1GmV+3qC
TRPJsyqvFy+wI52kiETCaSxKTXwmhL+eGLKD6ctl54yS8Cj+1r8fTcnK6s/cuZ7s
U7zjS/N6ZHtgfvMMDwXRZOQCw5flfoU3Dvj31jvka6nwR+fBxHxWRnyVgB1OMmUq
5lY+XEcg/2uLqJw3iRKqZ8gNmroFhNHfy6pVDRRi+PSFQTwvzaJZjcjQEqpIOzbb
pIB1/vMh56sGg5T+JCle2hiPYpdAyPQHTFUyH1zjOnnePL6cEEqe8rUrfeF3HBUl
UWi+CTNKXEV5AWgJrqXxkGX0YVsxQIfrVXnajQCpfeFi6upJd7gvYB29Vh7LJSV3
1NvXayWqjJopodual8UuG2K5xY+PNwfscQx/fKUWCmFstfXSI+/FYDt9DDojZAUR
YFxCX0c8aF5xBWips0G5Uk9RiKUl/7NP/Jv1eTI1j4yxu3G94d2d5eYOeQ/+ZBcY
aA4P9kBt9/nvoxj+cxae1ZwcRJ42EyxJc9Q9ZdyLopSEEbkPOz51POGTRIYgivNk
6ZyACRHD8rWIRrngszm3NSf150atloF0Pmup7LJUzQMo30yX7FhNzboD87kv955F
veSo0gdWe6q/BNAZ/KA2f/Zkk0wMbApVrqPgyUQ6gfxDiq+PPG/1iGsrrjRdIcZJ
mEYAe676dsSbC5ci6Y1x9iY7veqSrpwgmYibUUC04TTLi0a9x3h3dTmSNL+2rzTX
+5Jm+WddhYjprXejQi8HP65WOtSqA96vOuy9qSwRZ62XxAvLaPcvQ6Oj12JTpJ60
mJXfmf3Xf/qXe37OmXL3lO/PSkozXRIeXDk+NwA1QQll1rXffhNz0Ksir6h1ke4h
byMJzv+RgoNHxXmzWnzrx6fEEVlp7B9s47wtVnU35FzqT/Bk49s/vIahJANRt9Qs
GOKcDReHRnSh9EmlaksMDF8wum+jatILDWRE0RXDJg3CUVNUcotBxSaEUpU9jL/B
G76pQPCtUAimm/EgmYb51UXlLUa5k/IEbSEwJxrihOxtdNiKGSa1n5Fj2Z0FrN7k
okaXdOYfNl5ebSIpt+UHuzGDiFmWB/gOHysPUkqWxltHP3QydqqtDZ3gE6t8VtWc
8dXLDFeO47JJJIZwp3cvageRXpy56puK+/ocD3paWON+ciXCr5sMF5qiX677CUEH
/INQfbiOS+t2MX5yb0Tbn9siT64EiqrYiVDQbPWrdq6SXTeQVOWqmZyVRx9/Bq4r
PVnpCU0Y7gvbAqDuwoY9FpinxLq542f8EBSz0P5dbzwJ8wQhvhXJmLCV4HTlO91g
7zPH1jPspERyMgFTfK4fJtP1Lp5kbdnlaOaIefftsL1+kI2l4vF/U4AbZw5EQfTT
nhDJ3JzeS1B7/cIyJoBlG3I9uptQLWqYSFsXpLTd7/26TDKk0o2148+vcAjF7lbA
E68hBR0gpJtsmsJOVxPP+kb6vog56McXfogU9WKp5RrARaTsRNbSAj1ORYIHqQy5
V4vqPoFRWzciRCq02rg3agCr+Uhy6W2cs20KhhRfbqoSWgIzBiEu3qjWZMECjQNK
Flvuq6g1w78sFrhSYkvcblwZAy2174oubBl8s1wzxIS49rWFGYlYwOEViUcSsREh
SLdMX4nVbOK6fqZH5YBgbWBOjNmy6yK4Ot3WD6YA/JNRUbtSrubW88AqVFpf1Z/y
D2x0xeDmL8o97BVbfWIr+wUp7lMo6/tf7c+FpyKTdr2CRqT/vqQKGVbOTAqSBJTe
vuWH0LtA4UEUDq3B4ogT6OHPyHma7NAyW4lYKZhLlnISV567oi76YdD5ZVlf3GtL
LeKl2TP2EKCeb02UuP0VEAQExvWeq02WrdlOceJGkhAmH8G++q9AnRndSFQRQR5d
4G2oePZFGrnzsNbMUaZYZhZoeCZxb503OsJ5OJQcM+2/4lP3fBkK/K2t/+/lunpy
Di1WT2T5cFp+Z7iNvjkrhwZKNuRfvSato57R07Bd+gdE0D1DQ7ivyE/KjbKz0ac/
74spS3mMZvUKPqctAXIehoP3hs+adA2sgkxjhjSRViHnUUDFSiIVJAkFP30/mpQY
ztw+457K0Kex7i0jQ0sbTFRtGgvUoz9VGRm+rgJT4cd/dMAQlPFgMvZ6SOYFKCea
+xq8DLd2FqM9cpKgPke+KVb7qM6aAgBTVZ0kIZNspBGUXLCgOGOJQT5jnEn+aRSr
YePDALA1d+1mr1hp3uEDj9FtUTz5b1MrIPF+8CdyJiNodqWbRQoLkesbfafqwnOw
dukU6aHFmRPToeIhd1/MaPSunQWOLlhCeiaCBsvtpsmlk/BaDtnouasrkZsqAMnb
ZNnrEh9BT+vFebgb3ICOKcdQEMQv4aIP/16nqVoCwKjpKaCcX4DIhywlCqRizRwf
K661nK6QMA0E7LOHHRs20kZfrysi4ENqrB8olCwUVbsM+iAjxEWKR+8H1hEjO5w4
dO7al/c3/j53umJV0aFOsVmoLvJw/xaGUBbm5wwmkmsLPFMmwDyPhtTCchdYRf6P
WiYpo97f2EpHCah5dTGpVKY+GDhujb/n7am8t5NkESV2BJGjOQEMmgBroRAG61cE
DmkUsP0Aj5JppVQYoYulLfxx16I2fapCOaFaTIBrZfKbftl+g1lJmEscsgItwDa9
vpxbAZLLOvhFts+/V+BKtkaEdrPl3V4/S6MMnyaD2zWXWiEnmOxiVg9iLfzt+6qq
YSGoPDmOhWK9G2OdI0vwONyCg4g4XR9VxDPsq47nqmH6X5e7q2aNppBcaibo/+gM
rmvvoLQHsciJlJMUEMWgqVkn1g/RVxRsQx52DZc9NIVob6JjmY1kOO7NgpphhzAa
olsLPxgM+2VPs96Q12+KwF6OIeXhL6RT33kQ1u28Y0krmdMGHmGBKd4Da9hl0UEU
cHHcoscMsiUYx3brr5ckbogq116+OC2pY1+XqWSxj/tAGXr5muZR2WmxgGJmH33x
xkqc5OqyqBLG7Sb3pUSholkK4xUIRh4+e5KwtPTSPJa0QzR3CzuppKuS8gXqhhbC
pb0KGaFHaqRcXVgpYLZiRPjGYMNpAb8A0oh95IRMJwfzmr07ou4KVqVi3HKD+sPF
Gwz0gJfWJwVKHUqJ+VuYAaCSrsQsDfFpQuatD+tyop+vfBZEwsdNFICDFhVaL3C5
HJzHBKSyXXfBXCY/+OnRGjaHOHGe8HyTbm1J6BKRdTQK1Z2idIQXtwAAuWQ7AzQI
V8+dfAyeC1ZByqA2eu3WylqmrnsIFw1sDFede+cZJeWLxGhDbz0/2o3vdj2XpDcQ
OeJAbLwdmiL1JZwwVn6j6xGkmg/4/VZgmetphnBdSbOjmqHh7JvIvC1mbnkeHik1
j7er4k+mpfaXYVdCVkhPbMuKavsKCHgMPfh1kmsggcqKXWxu5+V2+eXjYE/ypVQt
hohrgLBr79XJ/7787gxKChUJX2ulFkaHylwdGrxrcFjhbOIRLceE8PQ6eCo7NDN5
nrItrpNFCrVm/IiHDmObYwriyU9aQ2qZKGgumXfZbX1B0BQ4JlV3UPPEYWnTYBum
ktW/xz/+ZVhzruhUniHq9fChU5e7uCcmFPTsNNVYCVe5QlZ08AduuWWF9xbMWdAP
vJ+JNGwT3yNNZ62QOy4AW/kA3aG24IljFMrv8QXsg+tKtr7zaF/Mrd/5OjXEDVho
IRL0YKP9odSxh3OyQXDW1vfJ48MqJWkJHt0Kg5gCLVKBRL2Zrsi8lO9k8M5katuf
qdhnCVqd6pCHarv+lN1CjCMHk3pbk4we0LK14yRsNrMOHwuxkAF2l5eEHhhvHDMR
Z3BTEuhcwI1wEt3l5UkJlpND1reDSqlGJ7plcEMwloIsQZDOZzuXUuCQ6csvpnTn
UtVy4SJsNJdbDBko6wIDmhsRO7XS4A1BFY66wKtolesoY/ryMjw5VvyQZE+t/jYU
RWDclioNpzWNNjUrA6Px14AN/W/zLQ7GL89WUTt978kvNHc0AJFif1iOBfS29lsk
Ridn4SE7RY+finfa9hHmGojPRYmXd20itAol0h6zzjAWonpLnlJ5SefnhzUIPBHr
ViRGzJKhRlq0by8GCciBb7z9mI2zhrRxMJAd5BqFz15oONAhyFelprm6aO+Lf4TG
AVqPb0798zR2eHewksX8Rw0J6CGayKiIWgA88iGrwhaFfTecRo3hblNXfLHSsUOO
trQJ9q8Zj/Bqi0jtM5TwFKrKKqSa2F5lIabffHJb5nkBmifG2CWv6TGqbM78hEGo
+wTUuF3LEBhkk1EcVpnfpeffasw4Lyug84EDVrGmKQMZAZDv/BQ6Z0rVMFrzz91L
Nme0acuCEZ6ZWH05zRAWA/JeBBIhUjPZBKd7EkLo0EMi9N/ZeX1Upr/trl2HPDZT
HkTOdrIuTuGT5hOIlYTgW2Y896b7kx1MKZ5wvH0iokZej8OgEHFwVawwjtVXD8x/
olWdnmhnY4/MCwXp5Vdf+x0NtESGf1e9/BC+V5OhVk8Ety3gADygJLeZlQyzh/7H
fR9ULjSbXhtHPaP361j7/krRoKZfLZWDSqBhCRSZpU2GwTuRS5ojf/4wd6ZgPVYT
6Tt9hQ5lAiLg20l6/PvUqSg7zf7Xw9TmTMX5y32CUaxSc8o1PkI9hAfbU6zJTOXL
XX43Ut6nXuCVM/LsnjbGB2qcMyqDN2+XxJut/wOQk7KLaDChwV1a/V/1T1yPgGKq
eiWP4wvh6C/ugGG6qqu42h59Z65ZJCVP9P8yEKxjCCKDrx9rlceI19QITNYaflXi
OBRgzfbFfytss3lBGnvVswc0FONWVkCkOUR0P/lym5tsZjWHA8evZephyBr5x1K/
cMvc2mBIg0YO03SZfxYH0RtACzR8xC9qwKACIv7bQ8mdmQJzphJamQoNhM7PfBHi
3AvRWEcJo2a3AysijtHAzV3IZRkhP4eCP75hY2sfXLsSnAacx6Pn7AvYuzWVGtHZ
hcHGORrtUaGNP8y15Pd+Z8GXcxNT2Oy7yQvfbtkT1UUXynWRU7xrilOxTpMdfF1a
FCj3IwaLBy6Q4ZTnB2n5xS9UJ8Hj7L5SbUyPlLx58I1r5081rsgg87aVM4q3NL0n
bsxg+WdqKwiLfC1Q85lKrzWwc4O0uK8pJERQLOd5FMKuYDZlVnpoc0nUg6wCTklu
bTmfWygp6o8Ro45WU6ShRpj7PHE8HESXB11suCi6wMAGNkCPJAfml2Sd7Cq6yZjW
2RLquMqQlEIUJIPViNIvuyBR5BKlFM6Pu6rdZQjtyslQ1X6c/BmWhF919tZddtoO
z9+mOrg7mKvTFWJqI3FBkVhlRU147BMUWCCx2jj9EgDPDHHUrdK6oqVj04gjxCb+
6l7Rg5EIGLWjphTAyYy1ed2D4M9LNowgrh8fAupfWuT+xX087lbqnj+0tbRsUz1j
rWQp1/tfSg/eLRuL2/KBOqulJwt3WXNB3gatbn/WR20Tf5k3qis3Uk5xzWl2sSzE
urEjSOvmjSJYS00/wEArNAkfgWtmJJEl4AbtQEQuWuhPriPfyeMC/VkRL8nSNOlU
Ees44KqR4nhSMYVw/pOK8p3oGvG5NU9Z1YquFi8RED4y3ik3tHBRNcwkYKFj7Xle
DT1UwSPxB4oXGLoa+BgNH4msHGlBYQdEMZt2NJn30vh6bRAk6OLDPdLHKtUx9j0W
0Fv8trt1zJDU7b1kmWAsGvhMSp1IpDy7iXtQ0OsURYbuaYKw1DZngsWEm71JFINf
uPcaSNwkci0NwqIidsBIX3zaXh70p1ZjzPzCjSPpH7BxPoTZlbuxJoGTh4GvrgU3
it/NHWunGn+EluVnqAfjjklsKCGx8Kj4EVEN0k55G4YCvms8oxU41oVjvzvgXncZ
z6XjMU7TGo3gJTKYz2kjljEFiXhp76xJ1dYR6lQB1oGwtXkj29fVfDglliujyrMm
I2smO1quKDWpUdhp9AfGR5aoecDcB+cutPcQP/ZrxcJIv/iL2KoBsXOsZ4773MsV
RWnbrLGI3OL3zSVRTBPHL2TfRzWiJGlkmB2//IgLtI4YZc7pb/nDPrRZ+YdIUI+5
VH3kN2tamjw9rZhBTrYODFMfYiv0SOjWAtSLncYkS61ZtG+OfnKRsxOgZnpyclr7
3tbFtqBZhyiz6MSu9XqJeNWvws5QBw9Pwtz/K0IO6sX+AMeJAl3Gy0Wz+WvZxv8u
Zh9HHXxzM8Axa1C1/v0Fg8k14fs3A/xV5GQmVLaBmKSQliFy9f/QSr2RJf5UBw87
5tQT/8Wih0TrdhD+zKW5bzqHlmTcr8TqXSWBJkACE1hDcGFCEl1v/bXBnV0zJKw2
UZUPaLS9HtKatT3FWx3gKTdYFDCqoLsP8UQrxQAjW1/cZfp5jThKIsyReA8oQW7m
hbRA204nCfl6W1yY4FbAWdOYnbNiAIo8kSxThhVPCEFvHNh3xx+c8Ix18smL50MA
daKqfmE9CWjF42E7ZsdaD+ofJkmATKdlswn4oxfYOzUUAbtatxSUKZ0K98PREOFh
r3YDZ3MKG8S/p80BGzZoPbfWtp781H98ioW2+/Ftphxg3pOxAkWjFKOWluFQFsVr
mHWF85PACz36pr+x6cB97K6rkTaMSkkttnDqXfpJZgkHmoOhCpKDxIYO53EOt4k9
Ay0hClPi9Ptmsz/xABx0nRicCqSiRA6JVOPzD3gKXK8A4OHZu0zrqZk6UzsZ1cYo
mkkzjzaUCtKoKZ9CwOgcGu1OPeJOXzhLxwpCDlHHHiWpBhYzKYHB0Qf+obJaDk7h
6IBJRUVzNm0iKDBxT/v/PXiqGAOApWDcdBVIcNPoBXR6Mkn+0tTg+inbHPGdmz1L
gveLPDoEKr/6j3ml1akbqfVQJRxlkQbywZg5D4L34yhGkmTfjuaLbJSW7n57EFkC
s/jQJEZ2nBSa1e3xfZq254gL5rGotlLrpl6jnmLWIhYWyaaf6aN1L65naDnfvuWc
fbP9k6qh4j9Y4jfEksP6qH7n2OejE6cbOMQpEPsW61EIlDDWSLowIO7xel7hC1MZ
tmA2ORgEOtU5Mf/pEZ33Ad7SOg/BpBVZGilF3Ad1lG94WkB+4i1KcmqDF1E0Xl3P
pwtdE8IiBEqlZ3EmMKWGRXK8xobU2CiQ8XlKm/AsU3ou9GP2GJrbUrGlWGj2uORH
4qat/zTmXUrVp6NYQDVgNn/JndwiikJh5a8YhER/yRpUSxDQajj4abDlnCoFdYR0
Dz7MKYNnaTSqnn/i6RqkIZ4bBoTCisBH5GOc1pUu9n+NKTYm2Jj/j6BDO/7vKwK0
VVYgKZ0NwX1SZIeJQq5dXJsw1ZYYkV+z1/9fqtBNaXWvsyTpjbADVYs/fMGLi9V8
UWf4HZa6we6MONEc2h1y+WnwY/A98BVUwgpRig+5S7/5+37tF7DdNR0BDa2GFdWT
bJsL5/k+BgdDwS0tAzYCjm+f463dxMxX43p/ujHaLxX0NbJeb5ebzizcAqJaMzde
scolMlRmQwLt3Xb8QgnCdSEZaVnh8RJZcAE4Wqwy+pQYD4KeHywrEjQsq6aHJyUU
y9Safx688N6LzsNwLZ0bDh0bRe1ZBsP9IZElUqtu4P+AB0lkjF7CysldQC5N+IwR
OBHNBnp26WHX+t5U0av8RjrR/OT/QtOoYkiKZ/3+jVgdhthBduGSYDXLmfy52/y3
vUCvWNKjP53gc0N5aMuYEqOTgHDnGCtY4EQX0zncmPj2vn7d5a5+es+d1I7SqEsd
f82mC3K95QJ5Boamtud7kqZXDHz9dGbLokYKwuZgGwjvhnz400VIGJIvVAzp1Mkx
bJuDEVTn4HUmA5zjViC3lcXofgyybqlsl40Gt7E43ZBObrsngRgNvBzhjokzPLZ7
E+S9djjD2lxvhEEznM+pWkh6+GBBQE704nm2LmcbEKiLWXtZPCC/02qjdYtR/HeI
tP+P8cxQxa9wIIjFFU2hr8/GfYz113Z1VHLt7yK1n2G1WL0ibe7MnVnyXksFR1M3
FETY2W3CoIw5mktiBBvsik5Vhqk3YWMx8qUtlLU3kaoz7V/DHZnwc4y5Gzlgvje4
rM8Ha+j7G0NDRn5njtT7agJTLpx3HX7MZRwIoJK12SllFxIX2O4/rnC1mIw35zAy
8iWjdNsu9uDjAoKDrTHPxC+e0D3VsLelFrEJqqMiwX+++x2mI3pQDKDreQ5cLmi8
Qjm498Lqxya4lE0uVEYDU/B7DxkKHd33WuCbENga1J+4AeyfraNJFIpRtLn5nO3a
ocDgdKTj4gPDULkjfpb/hKVgjd6/W1padweMlSiiSdXCJVwUVWuET9o0psnKopea
mOF3zfSTBmJP0eECLx5+LHCffzQeA4sGp5PEnN5csk2H7H4g4Pk240NFgVe86MDg
lvKBCVMbwzPSu+zHfBIYPIWi6eIk3G/eqq6rsXYPywMcIm1dl+YjD6ZaJat/6YJN
WDCwBC//REiswklG5ynu6zFMVKZFN36SMbJv5I/4XfSJOHV16BgfrAYDUUYpT8dY
JnIIfExKIoz9U5hIBtzAAOjOswIr1PcHZD33Bupdx6qRXQhfIOPLy71I7F5s1BvO
YinX6hf0vK+3exIcM/OwymdPjt61MLSwbgmw8AMxHrmE81yyYO19x9jwEMo6ohVX
GuZ8hLkUqcbTUINat6gCabh1m84QzNYA7imnU5H9awH4vecgd7Zhy6naP+sAjHNe
XjRegqFsaMSQmgfXqYOYtH2IUMcDR8H66GIdJ+IQQECJmOGyh27/eXrXsUl5aO50
OPqymAeaw727L59JrTzTNTi3ov2kGVaYqQWu5KXT0CACCpRcz8UbRCQc5kbFVJfG
fqWUGSeKjEcc+QAjhDqQzM64x0JDJgfxs10cbrT5xdSQUpAkkQmLDdiPWN1fDExM
hljeCvCdGgMf+p36SJC8+H6dFFEmv45xdKwIg6h966tu0SX9WqUSz594QdS+jnld
N7R6GlUat4/KXnw9OqiVoR06epsGu3QaIe5ghadYB036qARh0889Hvs4Edd/jX9n
EEuEoqW9DxBXSh4g31gusqvWwmC5ql0F/c/HS4WTqG1XXX4++E87ajKhbMubPIJh
kIxdXaIyQsQtkezX+4o9wQXIsQGfy/bUL0M/XkC7Gqjn1v4xxRfOits+WlBeQcEB
M0IpEJQwlSss+B+U6J1EsLOwailx6Dt9F96vFruuc1eoVUaqtxIW1twZW18KHbvf
CCHY2TbjjrEeAwLBx5OcQElijqvyuHf7hMmS8j+XLlZ/hgCDNWsjdDqQai6eyjg5
h9jTzXPt9uLA1yHaUJcB05JN3kINSEwA9YsKZ1bLDagCtJfEKoU9uncI5pr9FCtq
Ofpkks+A6H8xwevnsVb7t0sYphAB2icwqATTEx5oUhG2CLuLx/2uPLOHcx9lOHPF
IMISH+prt0QD6dcpcY0jpXx0HQKc6/d7MpPRVv1iM4l+ZtC1+HRf9eaJNZPp4mxO
u8SPJZlCnu93qq1O1fNmI3cxWAXYZBCqD9yl2+hqBO3LKBGzhedYlz4FQdVUoxlU
6E+/uiBj6YBwaNscYSI9AImeInXPmrePlfqzurNUKKb2cfa/OmcHvCxUgyBJ9uPz
/dohP0ZOezxYL/QQ+/ZNEZJWdeZN1APLh7OUHjhLHIJ+kcRYn4kspEyryP1v7d08
tqupE9WymvM0SMVf6WoIbmJNL3a8nD88niimg266SHKcow/Xo6y2sfHo5wtImlcO
d3utUIKHb41V1SN5yjdy3VEEeho8VLfxpESQ2Wgcfn99ljFMUQHuyQ/Di7ensqtC
k5ynFssXhWmN91xXx2xU8OZGHKzWmu/s4gSBr/YbdaVgGoWI0WB2z4ChFmxZ1V1D
COxel6lO5+OKrbRP3cF0LJWX5o3Es56JbBzRFnD88XZSGBysc3KOJ64eA7lsEfzx
HSFo9D2bRGz4EAYEISNUTTp7yBEMX1R+AW3M8m0Q7+Ikayu5tGPxyV2Aw5iWf3ro
oHgwbhh8kpwW8IphOQKxPljLEDU4Sh3l+0HvFZiCXoGXpWDeKBs1TkuZ11Tno7pS
RGTualpyPMJXLPiEhrd09zArZ/NLq5HHZOy5Zu4w7nQWeYKHMum457k6lYTqFM9b
w13L3nCzJawJFPr8Q0CVczMbVlPvKeclkYQgHeS/tdTbqHdUAaOrrv4amx+P0QbV
Hu1JwY6uoNmufsB+z/0fKKRtY6CQCjuxp0IgtZSTpSjpPi/5ZmRgu8wsA+d8ITdp
6rFaVkWbTcYCE7uUt5IhG9aZuo/KkX5TMxGNDRjqbTa+Xg0fQTvoSxbk8sQNRBew
x+3+cwom4PgkB23+Qq8U1ud4Frw63VVoU7agYqFulIalsRE/03nKNzt8Uw1KmeUq
TRMw1FERvvbUOAKyXXxfyHSDsigb46UoHYWvnNeJHZ1NbQh/YxuisoDx0pfF+Ftu
3R2Xdfffw26AbOJY7MD4UgigCS9GYJaNxHwDIzVXYozhrFSSMek383USnHWp+RYD
JTatasJVCs6KLzGsXknuIaWtq0P1JocHK4yhBPrAa/J4Ptox8rqEbk+ZA0WoYrZw
+7yW9Qcwm6HLAhnxWM5DT4rTSBeULtykoCMKgRGsDo5p1EXTv6uwXZBASdU7X6MV
DjoIk4XineqWdEJO7Zosdva3FqmNgvZQzK9dKnrO7qMdDEigaIkjQvnSNlj1IYpN
CI4epatQlX3FTb0i4U9flETex+gP75+DZhp8WUtkCc1ucXU9CcHBQaEc3427zB8V
tGo804SkU4z80uxH3M/beplCJqU0Z8GIPnOAjmf8ngiZ+BpHz7GsOu1TkyYI0BLq
6wZZTfc+95tyYrWjtN2FrVYlWwuKAbprcYi6P3r7He3Q5RV/b6VIxxZ43Lp29rd5
OdRQ3BMiNuOSof1M1gGlkuVscrBQLzXOT4WIY4eH7yEkHO8XzIka55LR00t3NoPw
TRdbAyhrR59kVtHwMA3x6fDK0TpH87IKEoWDN+7JJGq9peoz1Bwj9nRtE2DJD0MW
AI1XTH4vieTumt1SX/qwVMPruo8ETppLMjBHow87b6CUs6UNJIvy8QU3AFwvA3oY
esAOPu8BsYG2TfVtFV0zSfsVMZmbeAFUbi/nr6+CttVZxbfxOsrY15aGSthOWJeZ
UyhiiFP5dijeOVSPIUNFMaGV2EaEAU8bLR8C2JhH7OYYMKTNs+t4IanYQx9LMLLr
MWmom/sL86DERSFyc3VQ8BcMFhxooGjMCH8Yzdq8GdJs1/4FsluRe1SKV2oDofHW
8F9yGOO3pfOUnxGONVjvy3JEdjHS4Pk5jg8GlPS3WiPJv4O+vQTiRocY1uN91QzR
PeTAdbFA1HbvC+3rSN3kQLU/1TcWzgo7vlii62vl0T4IyfMACI/Pe5e7445zTsLV
6f5cI8U/onHlCD58ilh4p6/8pfO/39Af1dyFxnivtIO0zaISqQ3N7GvcI9GRCNSG
FEXQnJMA0mG8b5wgCtXUArw7W33qCwdK5stA1gs1R6DsPD4CxklnADPpW08VN4gO
hl01Udrl9fcqfCF/1pc+KT5QPhTxdKFvB8Rqh7VWSF57qChHywn2jQTzf45BbdUu
+jbzK4SUPGVAg9Q7v5+380Dxk4SPp4WAtn+jEWupZA/dstC5pQNVBB89tQAwu5Qg
+jmWTIwjMoDxFCoWWGqlzRA8vru5bNUDDFm5XcyO/FaSXN4Ud4gbnH/ESFwTWiyE
/PMwrwMkG3Fjv6csu+P8ZQr53FmAY95YGdQZG1G0A1VNBtn/netqNB1HbSkbqi+3
4XnotVQ2Cf4YH1hW/XjCcVPiMR5irgu9ow+GKtql9qiMXgwuqUzsNndWh9jom0jI
3k2SyZRCzDbQRKg/7vxGHazcYsKRiiO3mJXcoyNxoJRmB+ELv1fZFSAjXrJxd+du
0///GLor5OB1qYUTxvMhQJ7TQYDhbtqcFg51zB/IBfHcNGbylUjQvqKqpbaYKbNe
2gwFQAa9iPmTMarQX2WOPixWgBj/qWfw3X/QGtryqOv6k1Uw4/TwryRMJwZXGq7J
mzWkzRKfYVXI1VRcz7xrUj5noZbYwH3mZyos3q5yLlt4S8qO/MonAG8KlTZcOH7/
i1I984KVzcIPLfOBsJIPo5qGSESwG2hIl/+19Anav1pCoyVcbD9KRYjUK+3YETwc
U5Qaj9XZBIkrw4DA31lXWDPAVFq2RS9tKVp4HX5MEw0rwYY9Ts8L0Hmb9O5CGFGi
2K/LRZwsPTAZk6PnYf1gJm1jV0pZ2Y4CeH+aPU3T8HbXpjWEda3XGrJJtyHQJ75G
9wxaMS1G/3ZUSBOv5EXSq0ntZYJ+E6lUXR4EDuReXJJ/dzTTp5pB2fmqhPz7xmer
ellUu/zCl9H72Qw838L02lhZtTNAWnLUPABQWgEty3lMlNxslR4BgMpmcae+17fn
paa2tKUsJ6vFuEUKkUG/pnmVEEZuYjI1zon4rae3eEEUXH/TmFTTL7gzziurMLFo
EtXIHdihpfXp9mzQGfWUh9w+IYLp1TGVgOBl2oHntxpoPuzlgYvN91fOU8In6RxW
ojFGarqEow5JntqDLmUCu5tSXPg2xahkM/Zt4AG+Mg4zo+GZVD42Nee3zZIhKgS2
0f21XbTvAAs4lapZn8MeVX9D+YpH/MDM3PugbMvnWnvE4MqMaqJZEYIchnTw6e94
l3bod5p4HTTfhjYCki4hy4pFI19hV1mnXC21QAf36MeqkwUQ6iOdbTsj0xWD9Spw
8e+630ciEa4aY3q39LDfnoAcmv5yvBErsUxPk21MCMBe4T9UfQEXN0A3fQqiXkfr
0W+2UdPSmhgFWa0meTTNNbNjZ1+oYbMVjALVg3UHh7EHA6ZD6obRof36vapF+jHI
BIdzAyl5oCHbTL88lgzmzyLDizUENE1ycqKc26X3JAwhQJb1hamC29LeACIYpf0l
snMMITGcYVVtcyqb5mlmQOBp7rHUnRXeHzsOFC/FyDTGdEr0n7sayGoMXdCy0pod
d7jA7wwAu9n8qm8oLalghxgZn/U3M66EFbR/7m1cyL5z2p4TuG4STXa63hwrWZ8f
fo16mOj3ARStViEGswyl8eXv62bEW8HUwtBNnLE5xlP6RzD7+NWRB/X4Rx1dVA4a
gYSo1e4HTRHfh4SvDWmW+ilig0Rko3q3jWWIv4bMCCATgOYKuIfwY6X6R5TFS6kA
Yl6sy3uDu/GsFIIwNtEGOMJauQrGo7sDZSm09/aXkpADJYRKuAxfeVE6VAcKtVVl
+kmjR6OAmEJsj9iDUIez5vg9U37sLUpHQGC4D4GMsTIdcgG/HcKTXfTamI6PWVm0
xZlEVozbam5WKvnZyWnRZT3eVq2baCGyR/peUOJv//fS7COqpn2riTJ5+gggvuBU
4gNJUG5zFbksGkH+ljS5ZcQ1KbuBME5HWs73w3D6syNlo80oCAtL9xiS/oAd8Hej
lvsDBnDIyRgKU4S/C9IWgAFeIa3Nmxzpp9s0VAHJCfQJ4xGsBs+vAgYgx7bpxnmK
lfs4udhQNT+I7Y0VVgz53q9h0pWCMHOlFNbXvCs3FKvaCyELZ/C8RLOnnnbCSDPd
iChM2csW0vtGAmb6KMaUmYknfeKuILo0uGlwdzQJNZrbbRpfLFvA5DflEN9FbkbO
vOtSWOnG7swlUiMwaspBryy4VYzaPESl6ihMU/CUPAOcKQVQDkTWbXXkNazPVeSe
PWSMefodZ0mDLAxGle1OBXT0DA2DkYMpCEG3bC4irTNAZg9GbVfBFJW0DGEzBf/n
MX4MaKuxfPy4F9xo0O5tN0mXBgH07gRQoIbjh9y6c9BWEYuzGjdXxBrau/BhMiIl
Hb7p+AJmeFoyegduni8SRoErHGz/EVnCBESG9VAjKQk8WsGV/tzM9tqIukVSUpJX
Kwqe+3weB+mbwlI45mh2mQmMA6+qgaVTsPuNFIcv3MSz74aJO0YfWZLbckBkAx+X
ysNXYCPXmtuyYo6ffoesn5xUjnpahtea/t5hcFl1H6iWOSYyi1EA4iFL8Vc4pfMz
4Xpj4aE5q6zwjip3S1KC81fRP6+4I+h6cVnTJ1nV6igivZv0qzFlHFUePOui2sZt
R1D+eu4x3cuwMy4k6q+i+shD9sscg3OPryjsRUWh4Np5/7eDvGimBydCDl6wIN/r
1sJEunfiWIKEUd41Y//m+SRggT32QGDyn+FhwcD+sjcHcrswM21u2EZJSycJ1iYt
TH7qtwxWpD2/9A+w6N2/gRXsRqUF2kVDs3m60qv0h2AtVP/bwGN4aVHVbJp4Cwe+
bb64yegxwCoNcPOQR0kHN7gE6Sw0kcj9RT3yYWE7N3iqoYREN4lCpOLEhZTsWsB/
IkN+RQWqpsYmL7bsdCS04zULF5g1DKLS34rMUFcTXOOswU0XXOeuURFmQ9LWxtMd
khCZUWl6CNA/vfl3wuuLxCK+TmQpy+dNY/fDf4vsVag4AJX44Tv05vIjwe2jslxR
j1b0i5+qn9ELfeGTNVwnrvgGkyv6haCgGXBWZwX+4k9cczK26S55AcUkLtN3GW4z
KFjxKLZSnWbk3lV3cgSSyyPGiiswKjvyyj5RXIWU4FAQ122TDsaxe7dwuaLqDN/+
Qu7jRveH2i/Lu2RI/s+Osyo8OzaHlNBRAWlwQShjpWwqCcSAudM8pAKVvPhKu/O5
v/unzBLPNkAxFJh/CDY83z01gfENl6VeaBQUqTdiKn1MjW08m9BXB7wqmI5y7usQ
cEBvbMU75URugpjot2hKc91UgiO2uWC5VCyEzdBKjrQY+bNZww97WLQDdrRJkeWo
BoEYx6hrpMvkd/JZsIzz0tcVOQL6MXDJpV+7W2KPKTpg95KgR/dyNc1pyYzSxBaz
uNeCVwG+Q8EMRQZcD0YTkkQtWs2h1rUz4n6ErKpjHxSrEq3AK2SB0fBk5CeACoQu
OIO0aEi90S2CuqRKemjoFbDjtyZPoA0VwRxgQIPPFzfIMD8zFajB5lDhsMI+RcLu
aIauTNK7v6XY5XkRHVOKzI8xmdw2YHAfux8feBBSAM+spLb3AHpXLedvBq0OD78K
nu8p7rx5ek1ngq0dtnFwoNBHwMSgzeO+MdWpRONwXjVoZiI4PCvfzWDSXqL9v4xN
UvT2uGtyz4ajOoGr+N3X4g+IPtVuE00+hIf49zkY0OuMSOhJKTZ2grurK4O1Kfxc
r2hnQqQuB3uaQwKA8a+l06Ob4Gmy+1IXySXWZwamotbNLdKVh9r0W8vFoV/Twqqf
URjznBe6voAgHeHOg6kZ/qSFKXWYVoGLtEHuzdC2iWxuBx6IGq5oq/imqIEFn6Ep
05c0pu9JFdqqzgDJIqBLgPoKvHEj9sUrL2WptRzg/cBkTw9evLaHOem2ppDYd6h7
1GxjzHGjFK/93kKUWpXnkua+64hpPxa3PC6wUzncsS9C6rfzunCbZ0B7V60Y23lC
5H332Sen4APtV7NV2jxeIxC4HfPxw7Xjw5mjv/IK3yO0CQTacU03zbavr2s2vKDt
CDYZTrDWNLshRzvBKTYtcn/CW03u+2VkCUOUf5qEdY9kNYxWvWVbonKUvPn32JZ1
hJBXI2vuvuqzzaCRqtkaPrPHa/M+fcv/VC5AGS0xSCilK+QdLFgDQBjIGNYUfodl
Nb/hRr73qKoSP7gtJ4TKX0bkoumRGpRUh+VwEEyOZ5NMXhEJUbU1V+lYzZig2SUT
Pu0KXx1uuXsg6gUcHI7+uEkju8CPpNSMhSyrI5g7lWtwjnJkhyMv3jcztu47BXZS
Sex1ooYgnvUVFI4NuFs5UmvnTcTe4O8wIqVffkoa8+5hNQEljo3aUDyTOOyWblrf
0sq1NDw/iD0d5gRAzYL7lqBvVnCY0fzDySRCEwdyas/n43NklCpieg17s3fyAnkj
ezkdk5yX4qZstWWQTiPenAIjNYWYJGDyMH10LWDvXQBo8xx00SW8WpPbItOvqfAP
2tCxnGSaHQRqFaXzIFwTPw2rlZuYbecohOU7PBuf9YEwIhqb8Px44xzMfjnhBW0L
Gj8JLIWU1bSh1yv6DdwXoR7Y3rbk5ZfhwVAy5b1GDASzpBHGvqqQbYAUrkFdQLi4
PaSZ/ittPmfDc1Vopj/4eTg+JfKqU22EtH0eAg+tQ8tQlGbFM/o4uiMer1uOTkOt
KKu/wL4xZwAa2Ez4Zqoiz1AOnlgH1Qyk8BUe22T7GOsNYetCuPQTjIg6nDSS++og
PK1MVy8OTCv+w+Dq2asoJpwIks+oZVPiKGoaWHvChQLzgwJ7op/Et2KqjWPqVNrR
YBJBCNCjDw4mfjKFfMhvZ3wtoPC6huG52iRmIzgNGE7JWmiXaUuvb0c93vNPvzHA
Lxjb5nFGXMoR2Iuv+XzerVC5UXsjBCofM6ulJBpaLjfcztf2reBOVYN8BTnDY/Rj
hbSNFupG56WJftfmOf4lyQWPpH2SpTYrJ3pZimK4+wy/gtLJgIiarIOc0Lz0VyyG
tMgk6CWjYQoVLfCILlKNuY/odw6/nlwVfQ2t69aIYw2e+v4oLq/RcddDpvOUGHo2
uqCbqxmW3A7dv6Bkr+ZfAWsjiysre4PfUQpG4r6GDSgTL1F4xcRgnu+Cnn2rwkUO
PlLTx6p9/QT2CaRnTWGfUExN9lSQhRIobN/mva2mVuqPSStW2s4EYT0PgmVAkc8/
dbRPhWb57GNHLpcSkMxUOHynZeM4HqYbi9Fc5Flst8qGpDaQyLAtljNheYv10FVS
s1cR4EqWIchmJIvdo2Bc+8TcRa6qlxfe+i7Rd6cGY4gHGYtZLPKX3FTbS+PFdzL+
23Z8nfSpHDuOO531zkKDBaDF+00drMahkxQfDuUncR7ZvdeoMiqPNm4ic10BEXvL
MpcrKlSLi8OUFAWc40aWhjwX5oJnb06pqgllPLuZ5gJQEEZ526ZVsYzY7wb4SCrZ
Xlk5q5giTkiRSRnOKge+ws6mKhYR5ftZb9uuO2FRu9o2ebbzq+Zp+JvR4Ak4yoXS
7TiXwcTZvOrqIoENyk/s7523+PqzeVaeOGIvqq4hqn7Ak2g9yVBg8gWbuSMQxoaU
PQ4rL1KBLU1Nspf5VB3I8ZLxiCiBFa7bUenQHmkahUJBd6hR8eAGave15Nt1cBNK
tQweWr1LIH8G13/f9Yqqy64NYY8NKbi8ZhD7BJY0mbbOq4UTU0A2iP1V45jRBkCO
ZxCAsGKbIwBWsS9XeEfAKjIyzgP7HdI2M59B27Wef0t46hk0XkATHlgCR/H3RUv0
WasGdRBFqaY9gW4fTFGQfpILp+XQ/BmOtgG6UqzubPkGxiYPQ8D6ln8yiPUIIJxO
4MK0XIfuvYagsXq8KudhO6Rjxe6O8FlVhqjqe1BrXjL2nCWNvyi+0VdybbTkhW9C
8f6xMP8uj4vjrZMnNHzhy5aUobXqkxHnqugqRG/pdNr9bsozCY3XjBqtcETHieRf
q7qRpslvLCoHdmL0tj4cxfS+ZfQkO6F1aeLgjU7rnSlM3yuvzHdIIdgMK5SggB+D
zB5a9tVeNRXLdQgFln4TQaE/YTTpRCskmR4nyM/CR4sibUixmR0q6A+cIyaaqEuf
k0nyXoFPiGa6JKTMx2oK2YJzr1CCpiaj62BZgyaU/eO9GX2MeerD82/AFjhEtxV3
J8dDesh2Q2eGSE5GWq72J9WXPXGovE1ikH7Qm3pvE00f5vEHprZQZhanjCKUPgH2
pvRM+2/aitDUYt0ZufTWp6F6DGOzWNbVhsKqhDRcGZzSVlAuEbbrSaAo5AO1hrIc
Famc6Y7HL5uh6QvpGHiFwvMLooz/ehqeBrTGvx6IGl0/+TBznhIeYhmgzWyEWzF4
Qpnl1f+fKsqchZLSH5ouO4HbFIzOSmut5jnuxx9J/ZRXgZrB2jsC9US/YZKkUQkf
fB9o30FX/r7xf93RW8zWfi+2orPD2oR/MrHpNBaZE+oLvU1BB4OYen1xpgE9u/ag
6Vh9AGrK9Ax62UClrD0xY/eGKG2bOKLksWZuDrHmZXmI1u29rXuN/vSzwtbCGC3Z
WD0lz7z765xZaznTs9rqtVwIdurKjkaEscStCAehEmJTYLRkX21DgCXxsKCUaxSB
SzjqF57zT8BX8lSrmldbmoDFjF0OZ1sI7XJSQTBNTS+hFQDNePhLYs87tOEGbUQb
Uw3Q1/jknpIF9wacrSx4bQGYBEqTbfrg0dofbQvoOTzc6Twg1mHuKStodYR7BbjI
IQaNZ874Ku1vs/YrPb0vPO7zPRBpGFQTM1b+5FUPrutoEA57ZYDnbA865l05htcP
B7VwX4/Au5N3i/V5Wsg9W+qWmmhANJa8JqkPF5BOGgIJuP7YtrzppD4I1bBMPnRj
yeHDb+IIs02wrPGLShsyzCfHUEWxBMN61NlJw4qHU3Hl8u16jGRAm7ChEny6X4ft
PNPmuY/kf+a7N9uE1PXUSA4o5sCQSwdcE9eWSsnfz7zo4OPLu4KvMFOrHVmqnczc
z0pdvmnzxHxwkP7wCYYvD12efkUST1SlnZyjLTW7C5uT8E/O79O4x3dNfGZg9IDo
7GYdp4QHVqobFNRnj9FtNBxaFaUiY1oEueoR7nj0Y4jkFeYY+gNGzD8TG9gni/9R
BN5d9m0+XbGtkjWjYNRvFvqrszrLTQhnEbqv9tzPIsAisgmY0V8OEqopWecH13f2
OjeJA5HjLBZiP5cygF/pcq5zLZOFmGLDTFH5OVQv8M/0ihvbzEhlFy4zmwTGyf9L
m22r5Dc7iLBuGl8HWWDugIymQEGC57YqhkZPp0CoDMrbOOVmM+xuF5lQ3KcyBJBC
3fjFF+6VB9XpyvyODZL9ge/CMVQAgl6RO2HTvdlH9hzV8VhkD68o4PuU7uETmB/r
eEDZir4JqKc7XumzrfBj8YhW6CkRp89+530s91lXLw5liox+i593aFNiW2pkgI06
SiODRnuY3rlshCE8alUkiLb6ygn8OnT19jbUAfgxkToxDqy3FaICOi8T9tzaNo4p
SBz/eQAzsfZSmWzighez4jv6Wu7ZVOg3prBWUFC5z42wQBh0Z/GGCGe14LKUSt4f
wx78qV0jZy2sLTCPSEjffH7RgUxGYu6sguyllPI1R020SIeW/FaAcDD6SHKLzSuv
rMFVahkAcezzYc42Q2XqDYxrch3FjvBuccWGgz3P7imHitLTmzmzQnc43+RzvC0W
qUuzAo067JjJJ2zzEsaDmwLUftAu3XePg8nkscqYsa2FXW07hKy39EpV/pLCsgTN
EpYDfUp/Hlb/PoRb3680yw7f9cWIxtRDiSRznSktq48LNxGSl0wGM/0K5Z84fKMN
XhQRDcGTBgsQdYFCJdoUgH78fEJuPS2DVBoD+LERr0OyOkyiCE83qMSmTlumZSCC
Ce3t1IwYnZ5H8BjURL+xjYtZK/WNZkhUPLzq4muiiFvdaHuciGoapZjQTigSzbCm
Qq341Q4DTGrcvna5ddIaLgcmwrrTOGZH81cJoz/R37sOBcI3Fj/NZ248Ui3i/gk0
ec/zp10dfOyzZVEt0PdT6jorqKReIoms5u60YLAHyErya7xhA24hMnrceSR96XtX
Ehvzjchib9+2UaQblyfkMmMVonzNAzhPsP3bYVr2oJ2B7pNDI30xqyHBhzOr2xSy
yL8nBekZM5WGq2PfyFWW2hJ0OW07DXovPM9RXece7+Usf+zlz+E39zEuC0/dfBpe
mVcbt9LoppFV1/EWSBNXyK9ZkIUSRRG5a45N0LU6kWQK2Lr9vNlAQ5MT9gENp4pX
kLLEgMrFKU6rvvJRrvn+yuMSguPFvceehUEs3XXkyx+szpECUZV07gIzZ/nlqd5l
Y0/0IfleYzRpx4bknqi7xCOsWMClN+hErD6C2B8BDNd3ADAlfoJCCQsMrAkLNkZx
m8MLa6UKcTwzGaFBf6Fal0aE1iuKreQEUzs7uW+dM2QRUaXDftNradIHXXHmRKXu
D1htfLEhdVN7Bg/rOkLjQ2dx2+zpAQ3yaxWl4EAxXYwW8+hXUpelfMk6ZUJ35HqN
7c3P74Urg+y71HgMO4oEEwaUJKZxnaXI6vDicfoMHQnqMJ52sTceammAQvwMCH9p
P0ymCqbMNNcHiXxdOQxqkwo1Qqa1/ZxaEvOoovxg/EqWvMqJGvBGiGZ0/VJ8C8LN
qGUFFVjzhLAJpBhEB5rjsEjntiFRA/g3zVfGXAQs0oQsJBLgCSMoB8K2vglhNeQv
VtKAyVmN8in4cqRbXc/BDs/M4qDVxabJtbxWc2tgp17VjEHc+kYr0e/GuuRHLhvW
9Qc4ui1ZEG0y87wG6eTNphHQPZDBKMFTNSxgAdiDZBzikEpMRsP2AcGIvz5VvaBj
Zdn8xPygU1iyuULAnXtm+vrzdjt7Fltw/81rqCAxGGjh3yWytHiHySwQx8WNv1Of
eazYCB5AYAEhPK/wXQEPWajOcZwLpy9mYkt9WiggNlcC+N19sMxYeJOEJViknCoz
MN2vPxqibWKlbAc01ASN5g4syz3hoS+5SNv4pkzhg79+EPXweXzp9TeOlL5v7uND
Y/31X70YpUdUXlB0yRwGAnPDb94XkPI5jnorw+UDaHpI+1SSyrmu1BcrhzaGvWq3
2TQR3ALUKG/m7xnO3STmv8erA9KYq6EyaH6ZE8Gk1GLbbzQ6KM8CDkGOh78Laj3R
sXfxiLVv4lp4d2acasx0BjUkAzTb9hq+36Wy8XH3mDtQV3Xo8HoFKT1RfcWE1znN
VGyeMoB3Aoc3aMBOBD0KgKmGf8dUKzecd1Zs0qpOkO//hHjxckxMdveIiV+vNBTi
mAdSc2YweRLVZTe4Je9NxCvHB8oh0p0XI4ta1NdbcA+vGOIUJWY0AquD28ruJdSB
pljIBqxR6gauB8oTtqM6azIxYrqKSXthUM0T2KPjnA0btQwxZzOTdHJtJ+baeQ31
f34kqEg93YWMdPFbcrmC7SOqUBsLw/YE9oUAuwhYM9F/gfgdynB85pPdiFj+PAcL
S7ql9jvOE10OdwndmvCeLr/XYHV6S2vzFYlmW38HvCbW9+jOjUJm2rl3tRdzyq3o
lH/YX4eTAe0KILnOf6VJ9QapqBYOY3fMHP43oy78we0sq8Q4dWZTdzEErljGai06
dRO5cdcG3GLN8V5DPysZgCDplaAyyOL2ZvSNk7GgesQGQmYlf5aRlgI21/mliIVA
OGbI8lCpoj2Mi4EeYvR2oNObDTou9Uurp0WgdLOz0Y5bcmlPIZ07dRHTi00DAJlG
WRSN26mc2/nnny6jOvx/p12/yJc0hV/OCwQyrOTuUiLFIvyQx4PItmexQ1dADPF3
JZHsC1IVmKwBVvwUlm+9G5IEd2veURlkxsvYysgl57J6yX1LHJxidlbOnFzjbN+U
QaKtMpJ5dXs4Ykuv4lL+8K0hbELwZAUUXAps+m+GquaDam2bN730EFu2GlNE7Vjg
AMDwjuASmaphm3kKwGR8SdpsGj+sLdYzSz4V6GIznOfIaYGzmOa/Aoytqx/0UUmr
p0cUVr324m/BgbpjEeVS/eLZ3PpkbXeFgO1sPCmuHHk5FBg5URNLTMMgjcDLwsfN
E32isvcK7rBnf6xYzC6o6yMj75MvzN73MrCpiUXO/Xzjez6OCuzbfJYw/tgbE8L5
3SNOAZMOFDzeFv8TNC+rdnBbBL2kh1fHaNsp+zFb7gDRZpRYsVTUD4iNR607T3EW
eA5SmcGTRvmCRVkLcUyg8w3aXNq7CvnlfyaYrHbifyujqhjdyxMG2ECRL3gpROJQ
LX3tNh6xdM+dZrWMeWTKePn1pmtyGETxZ7JKl/P/x+3YajNzWf0eCnPPMG8XLOAV
Kcn/hNTueNvGaBbQnERyOC2wAiQTjvfm11X4TZiqXJpw2mTd1xsMDVjDG4uq77dB
OgIxj+a7EPoto/xwmQqB8fRgqg0cYxhVUGn8+yfYS91WTfOqCA8pIa2sFg5UkmSX
vyESwsHCt4ZCeqQg3yI4ONcu9TKNcP4VLrpqDy+/YzRhg8dp914C6YWuxqNaAcDF
jlY8RBJCJ6e3TeglpisHEYbxkBIsdbsvRx0nZmoeCKNkN/gXNpxC/eS8T9Lf7ZaD
Ds7KI9ka1140AVf/bGOl4Z+BnHppCZqKXTc4g4Bj7wVDnAIGK4smFANB+OE76W/u
adDSBRiT85GtPdl4gYf2URkmQvkzE+CjEity2fN/pHE2sv3HFki5gAZWiKJTznG2
gsCrju8Qq0Ux0VzzAQay68OSPL3dpxI25MvDod03u4TEZU/biJR6KD6GcW1GoQGy
R+3DdhHJwFKve1s6mK9wTnZHvdTNX70AauHPPmVC5lLl+UzzZAa3dNC9tUUvUSnc
L4INEUI9bCaRu7Vb2Ii58Meim3YxShfHeo0Q/BKZ8lWjnEhGbU+/A0GdU+P93HCO
YDkMjH60IMJlYSVhjpazQ2h/BntGbVNUlYuc9LQR9gtPsNc4g5yzt/iSStrEVL+5
84jYc+mRZzGYMkBWBjWTIBJLCVRhAOEWa3tiEwLT4FWP/MD+c4yoVpyzkvtJt4Jh
r64JCmdLRiTmEKlkMD+6SwjdukcVZFohQEQsKxe342je8Iapt1YxNPfDBdt/RMx9
VxCDRSHhXmjBzD/1VHZz9gFASeJzmS5NQU5mGSRLgRdCDhEerFDhWgWrgKBPE+C2
+Gbv1aHLUIppnY8ZvzCjquWqwBsU9KJsrEfn709uXEC215VvMLoXdeyEvXb4K6/T
vZJ//U0UsDyWqJtEAtr6v48k7mCBLR4tTAdX+wlDNia4nl3aDvmPlnF7kOUmH3UC
ivJ69/1mx5qqWK7Q0+gPhQ7E9IUFb8IJ6mTqELVO8MZMhHJWiOhk5LvFzQHRbPGD
ZeODMBX4dHANITJrmlGQBEa2hlaBm6+i1lS87SjPwa7KTugfNHw0BVfLXFdJwZCL
oOOr/1n8ZxrnXrepf19+/r8qUpkk4zpqvrJ5UuwrueAXY0+WIH0zCObZFEGyZi+d
cCH1fMC2ab9YiAn90iWXCjWpM2NJWYqeWrcJPRVta+JZoNVzTxBsvA/l1d65Dncj
4KO8yMnYMecKFB2eXO0rzspzboElBJfnspzHh+x8rrorWqzprW70aSmNgfXaHtzf
ahX5khd/XdjpriQZXzqwv6zF+/dbTbGuTZ9MNuKqlImmxuAW9oqOp+buDbtB7yxE
4vQBIhE6PyssISEIlX/JtvRbllYUuKGbuhuTDhvpnPjos8ibaFrdHuMy8ZqSlyzX
8pq6WdRsxNJV22ZP4hRSpuyyI393SLRvcVJbAflZL5pQtVtXz++GsBFJU7UlEdNb
TYdzR4YH6F2coSd0xss00kSmYL362p7z6jJ61zQNUlRIlCVqYRsPsggDOjOwsrtS
PJ0xr1VNq8hNXXzspQRizWjk7cBqGGFc4jQa3GNL4Dv74gbOfomN9whjc1MwT//9
X3Jj6cUPIdE2uQr+HyEinDEdGMReuYjCwAlz/dTlpGyrbx0T59H0v/sVsngUrNMW
8muK8wLXdj3AF6kvBwXSKr4wTin8RTegmoXPd1MZPnhQEIunBTYma+aORctE01On
o8jBVMbeJdHf0t2KGkojApNqhWUvkhCm2UJUCRAKZDuhH6Hdjjox+9KNtVZNGfIe
UCAk+LWl05TcNKpqLHFMnpo2iPikZyq2U/16gzxLPqEcpV8DFCGWZQNd1ashWNzM
NPQPRqMb4SHQ0rlHlwcJIDySG1MOzfGiVelOXesKeICj9/SaD/u/PX+GwpfYHWg2
BmXTeJLIy3tk1OYcclJsTx+uyuwxFQhXDMtgTTN/Nu7sid3acUgjPehmMYAMwTLl
v9kcnloyLspmBHiaxybNhnY1pJJiPTLTFWIZYbWorrwp0HLt6IBE7G0mzBnM6+IZ
y04WGuefAsSh+/IUODtu4s9PoXSye9pVvzCVyE4fAQmhZYOuZKcF/0WL1d7T7+X8
fjHDsKfq8TCUDNDE2tC98Un9kd6vxUScUKSn9SVVPwAIELqcEJ43vzgBVlG/kv5S
Lb7OEju1nVuHvzCVNT10TQETmtG2ypmvJS7Oa9TQDpzrUd8zzouXEHgcxKBVfY7D
/yESwvKlIeuFkxJKMD4NMrhc8+UImfR01eKXZ4RsfGSKv/tQM/5i9uwcbXjaf499
ltgN6tBI5V/P+XX7bCgJFsLmhodGzM2lTqChDisUklmYx1W75cFyEFIJLXx8kMKJ
tjC0e06ONjHu6CNI54Y2IAbcVkYa7KnZ6WvY8vfYIsy4uRs5gKkvEgpPGZAJF4fY
j6pYYuCrHxJAPONW7497aMxd24xnslVXYkUYv0UBuZfjan0sdhw9EIQYlCvWtvtz
7IvZl3nSxbvOhA0uSzm5bxXtLBKfOmq+b2pvOG8sRg0F3XC4YGvPHUMRMyZ9znvB
rmMEtE7R9WpAFL546IXgSSavG/XsVSJoX9EC/7negI7ILtrV1xYtbFaNaDbyjabx
V/taQbktjG12uY4/OY1TFXlUqXJOFDc/dk7E6vujkJ6VrjUctS9f9s9FHfhxZR0M
94tyqZ918dc2OZ191ju0y8RlGqabUBGXFQ+4Y/WyacY4kAx6WGy3ELgDccoL1/Tf
ZvNg/A2RgSaei36IsDyEsM0eavM4qdTjset3TiZXACz9lAIK9rzzXkL1Tvn/PKOl
ZESvTICWTuQOvDCFHTImDGdgSExPf/Yd0rSEgKA4aZO1VTArC0WhCIwbuMDmr58X
JLmEZJEyCkZzkcwjRfJz2Id2L2N177RJXElY/p2edYbV8ci0BYxCE4PMTAOdx+Ss
Pt4Cypj7dmAwSwBKnSTJiYApx9/Iemp3KncwcCKv9O3STY5AIqwnhj89P3TAQLBw
qV0zw7PPPm0NVAzkjde4gyFGfo8hZ6BQ5SetbsFxCcbX97r4HbUmdfTSSsR1ghB/
88SgJhktZtf81Q0TdQbyHmsZyQjUQHGie3iXfFHyyE5ZIRYDoYngbS3PMxnvrFOT
DTlrXdVhqkSvs79una/2khe4BgTV4FF0igHmblUMOmYLEiQdao/mdoQo8niZ9phI
GtfeDE7GrEVJ7k4KLMCVu48hsU3JuQNWtoa3mHO3szHruRwYfEolDSVshjXJ5HGW
bMu3/mcgDJp/wSg7fGF7rvwgAU1H4lJIMt+8he6J//mNazlgV0cPMsFmdIN98Oek
wVKprHWU2qLZUmlocYT5Ps1vn0n/Z2ZDdUC1IjTmNHNV3yuy+VdcnFL2qhgzQn4H
pHoQcJGU/AKUsUYVa0gbUQr3Cji/LUKPJ6aeTmJrkiDuZ4FG+/KSTcJJ8pPYF7ui
KcBWKP46UFhBndR/gd8XsAbMHJbYTrybeBDesofO2rOPj49S/rt4GVX5YIHt/R1I
LFh9OC8KK7k2ghkdPmIA6s6zjKAwJpAKmdiebULhPJXzAbKPQJbnCEf4naVC/qNQ
0wbwBRJJcf3x9Bp83dllExP6dwp4hZdtT6k7vwDYLbVMUDk/z4iP9EUmV7A0r3o8
4G/VWvc2hTOpUUIWsoYHaekwZ6oD8VKgBTg2Zw4DRR86WUpIVvoFuYuip2zKESro
FDiy12YOJiA26yFThGKjsT1vkE5tCupCSCnKBYvJ87cc9MsGXADEvOJvvD2EnFtr
zYfVqLc60TQ1FohVMCwpjCsKFwGMAq95LX9KZo2MTlQt13qwy6ws4h4zFKLwaEQi
uFzX9Yeno4SNZ5kGwQ3Wt970Q0X3Q8OwbnlWOgJ+yU9c+bAu/Z1Mz22/pMtrDwh3
qTS/b0inhM4SnFQ+8z8IXlPQZxFqQ2ueXQmPbGMLu26QORyrashGJtKED5WDLCVX
odWvOLE6EaWyCaPzvbXMkuIm4/Uy/7dij9Ug1ybuA58sS4T5TArkfu8QtvNZpiAT
ZWa+OKB4i7iBMH4Vnjwa7aQf/Ot17N+rrtWlM7QGwppDfj0lIs0rwFIWOnCObfwi
MCwGPfGQMztdolV9hc1UDCXsh34mVAbfJ+w0vYsyRrIOqULwBJjgQwY4anytah8p
D3N3M1VCDZ3O8xN4sZFWgEjO/luCb3lzN29cBpG20AYptWuRXR8RJndENgM+/vs1
eRO7CwwBRlIrZCzvJccErviu070reWbk2GJ16l8kMRGPLEVAcbbgDZyIyu7ulF9l
bZy2HcVtMMRrdRpxBNw8rN9eYH1gRbkJng7uQYT3AmK3lLbQlAVFodkKUaYtrPAN
3Um/oZGF+MUZyvIN0vWNuC5LLlIZEEqARK2jPgQorwXe22kW0yj6s0mKWZobTfhc
wFb+IvlnJMwtzgnIrGt4GjfQcWRxLRLUW7Bx17PQKEn1zHN8Rx/EePy4Ug6D9/JN
ws69yc5c/MTOLIuSmGZ3nQIuMrJClzNpVs1S2J4rWUTLD5PL4Jx7Q2yhL/6fVUhn
Rsc0WukoAKvEPSYNHUzzS/gi8sPYxWhsga0qxmXp6349zPAuSf0sdQlEDDOu7zUd
8U1xW+Ef+wa+vmvH3x86m1Rbb0+h5D2Cwsjeu6+HSwlmM2+DYSIdthhNaGp4D4j6
ltdHDaHirR5CCWNakZSpvCpuk1ZZUNh23wguKeGP0kJ8JryqDLKHZIX7DwNJ6uZU
7e+K9qPcyqAc/DpVAEFJxubwRN1T1Lw6+z6wNAu1eSh3Gqqh5iJ1djb+83ffNWPW
gKAn5aLW21Oa5djgsKpSxLcFtWcMy24lAnWGPljBPYNUC6NZMZQbefQXA6W72wMJ
dHx1Y5xYk4Dip5icr3BKu7nndJl4Q9IfmCKU59PBjM53seMcYP5Go+BJSb0bt0hl
lJq/qdoukHEoHo3VASOHQi1xjLM5gTuK35nP/GLaEaFEYR5sTPykg3RIIDnBtC0B
gx885aRbIXvR9246xK+Uy/oj+OqMDClNqCm14d5kV652GUIWqitUrqG8XyyretiJ
XxXQQFJgqI6KUk5q/zh139Gk5xsmyxAv426rX7WTsn1EI7Nq+vgIOI9dt5Pmc8u8
o52h27xWcF055eGB8I8+3DKUsk/whT+Fmd75UUGIflyuDxLXIdnQL9YpWulthD4w
qCc2WGZbQOfzAeQbP3pr0O4UmrIrMot6liDR2VXOpMajxji3x1cR3EGBTdIfT2md
yonD2FVBMZ+eNOK2N0Gsk8Zj3eC/Y3a409ECT9BqzO5y/AkgPwJlxqe0uPkX9tps
bqKMDenzUZbnxodyYumIp+UwDqbqa3RavRBMzBas0TAlVGF4tyQ7aAeG0dRTr8wy
K0eeo/8bBYadoZSMfiFndq9WDqUOV/kwFBAZa9LSSloGeA6rh2aKZqk6vRTELZZT
8LlWpBa6iQE7/ssemanOiO8NDQqUd7m44ndt3q2tZeZYbmZvaR+zgM+oI59LPkQr
1B2/w7JaqKJaejjeC/82jvIFVYU0+y1tq0gJrRsOHj3bOAqDN84QyON6u34v2HZJ
3CqnIcHJ6TsVVLhzrsS+Sf7WIrbVONtscT0TRXLZ3Yis6IbK+xOJE6B8GlBeKD5G
0ZI29qhAfOzPOGK7Qa7ZWAEielAb0T3C2W1IftY3jhNdB8yAySjPZflXWx45GJ4c
Jd9LMJfv9WhFm2CqF8akwAg/QAIriFVzBAAASVaJoZCHrsoOqpEsWCx5nEblyj0I
JjMwtY6gznhmJEmj7pOWYi7uOnVjfKt3OwOz2FC9cjPO4VunPpy48iDdvmDpOVql
m3hn/1TbgVSkYF2Y7PXWcSAM5eKprsmFc5PXoprsu+qLz1cQ15xqu8kP8DRb4ok4
TaVoLkCvgERmPxbdnUQEt44XTx9st4657FHvQTsA7D5HX7ZdOFM5JTsk55bvL/cl
u8+8+rUyL7X2dSThhn2IbatN4DR7FJb95XF6N1FBUBHClPLq0EqNEh5WD9t84RCf
8UPXXo2T9ZNycVUFWKYvPwn5T29f18gpvN3+LQ5eAeEu5MRb93/zPsPuFw6MLlL1
zCTR40wGsEPIGS1rtU7Kc71l0G6cWAeTQXGvR8wlCI5nS96vPQD1nj7kTj8hHeb1
mIpwLgEtMdf2rI2nxR1fIfePE1JUNy6zzuoY2LsA8eL27llZrtsHoO2+W9h5MLas
R8iW+hEj22ggm1UKdRq/vq/lCMoElnw3I5RZfa8stxqGT/mcAbfxtP2UkOmdYVRB
Y0dSbc0YAiJyrj0Uqiyt3liJQ2a4inecdMxi2qKf6ZdyVOq//1xp4OtXYeEjGcbg
2Xrlx2VlQkVVX2vxprLtaCzV6fKesu4pEFkS2rMn/TuNdrU1r7gNx8fvxqaqt9nk
0HK6BVdwhox/ZRWjOAKItLQ4kZIb635hgVLodqXEH5NWhINnE4rwGfeO0vlKf3vP
4XEUvc6EN0Z4gtDBe6OC8x9bREhepTBBTG9PT+SJPz2cARTDIT9FtdI7TOTwb6IB
sEy4HL4S7IJfqyWv9tK30/e1zu8yP/JVbDpgKNOKxaOm5x9SrZt/3OKd8dXlqqYn
h9Hr2N/FW6hhP77c93BeaGy5HxwfSHmsZ/AW5wRxIUDDXLuoNjVS4N6y/7VSYeAB
6PkNqo/gwAvfY0spUSuZ9zWfB29oAVgbWbvKjjfVHprMYsqzcyN4wIeWLtzc4obk
WxaZne1so8xZJ0wMi1UIcvyZhnYwlSde045CVC4GwuTiAwiQwDvMKkEw1i8Tlf2N
rusBD/AtHWrjrCpL/hGd7fhXyZVSSuLAaFpZzbgrIoaagnv5+zDlC+qRKupbDN4V
xLVKbWzhfRIabQPU+GfD9gMhXT+wZr8nr7PleCQxL1JOjRIL/Spyh1st2Ozz+xiH
jHaFxsMEOZA/FsnVWSqT8KS9kQV5GAZTK/OQXS5Q5cqMcYTB4+yD3Z88Ph+hLmMY
YArUGhzUvHzAmWQ4JE6+FOgc2NUnRitVGNGb8IfQgEYcJnQpx54Thh5rOWaqS1Iu
ukxBYPq4k4PiCEbPQRT+zvJ3CpB8wxdbYhKfhtiRNfkdLRlEWDK2idOd5X9/JLRc
6TGgGY9Ws1KIxKCMCPV06bEgNDe5vkwLWLPACYGQ+NrAlu4hj4+hud5cB6vJkX+X
b2S/LRXswol6fy/IAlt9/CQlvJedWuwVWxQRsPPjN4BtNb8jAjJkhqG58hBK+5Vm
YEo8xcCKkPNib1k9eIqQS9ShxYLEDRmkoubJSTNQg6RCjNLJwTHWiU/O9Rz3xdMl
AXkZUQeDfmYRIKfSR1+iQ00WiaLyih1tFysxwBSoh8nCdUKzj0Q8Y058lYSTrOu/
jDaZTw8HRBa4azq03OoKHolOVhblAcWjV/07FYNJbHE/49PKK4wS40JQB+ML3Giq
Tkk5GyVaeIkkuVIMJ24mkJ7AfwI5Ks0jXwpn6bzDd69ZuJMmHKeJTJthpepqdKUZ
xq/LtWEM3pevWhBFjReUK2MfOoZuSdSaosZvpMlgn8Ufthhl+xuY6DTbRpYHst77
DcL3zGXADBsx0a8nzALcE7MZBLB4K+1zfhZLbZF1orM64f4EaI6Op7EKI3/4+F6b
5Aq8elQXAOzfHio9FRCLVe81AyykinaUHA1F+waduqQfQh1McYzr3oj9umriVuSI
P4uujEdZuDs7faoAzNDKqzUPshgEuEXxLy1aPZeNGCi5MAtZLWXgXLffbeRNRELx
VeD2rPzfMmSnaqtkWtj/gfc5ae2fuquCI85GE69gm8KZ42xc/EY6ZCCNbYmYJuiX
bueb7DUcj1wobqHB/M4V11v3YQFIxBhd+Meay0qG3S1xo4X8DlSw2KzE12QaEprQ
7Czv0jm8EftJZhBmJm8IFmIDUySStrV06DCxH2csQ4vTcgp056BhWgXiD+tYm6td
1fOVNz8K//BcEuUyhP32yOIbhELpGLYkTpeFZCQwXEhfSVdq21ijtsOqYuusHL49
L0xDL1xQTsHp49kIGD1c5ahgbpxCaFwix9M6Lx+DiVNSDoNL7oE3nKUWdvuw8ie1
zyErwLP+NDqjbgKMg7c9suxavcYzypYpwaCpyX705UeDzyEBdQ7N5UCBGYQLcuoA
roEPWU2w+sfKIecR/YuxV4eOA0z5m19/bvRhFRBaannhWFbPcSz3AbtmyAJAU5ff
ODifu62oqjuIUAYBloJA+8e62sG77qjNtNpCVjJWNS5veJ1wztrUTJnRjXpPnDTB
EO5IcBT78oyLIPEO9ltrJLAdtq0kk6/Qs/kDQY41V3dwC/nVFNv0D29FUyxSpLsS
tV9JsKJ4ir0VUrGZxslDCU/BNHrhW54XDlzPcclXJNcndxlCdrJN2cEWn1B/GEE+
Sy4CqMHg9kmmhDGnUV695xJLQ2erERI2GIYid5ioYSGo/JDlzZRtkSM8tie9adOB
BuD1RstW4Q7y1ZYA9/phB/0XS7C5ioM2SFJyst+oRw6KpR68pfeTnhvYahIBcdBQ
JBjr84vT77rEoweDFo8wb5r3ZSA6acPyF5wY5rsDbi5OwI8AXbhBcveR1HPN/PAS
yQzBI79ziJ5/CeZa8xjJG0myp7yNA+9AXLUJHQQTUGesApY5xa0k5O/PF0UZSmMs
s0nVQG6Mt1er0dSBGwJyaiw+AR8DiyYmJBITti/WXPUTH0Id7zoHJkL2hJVRV067
qSzhNMJalh4EVDXbrTrhOicgKc5/01IIsGMd6fCnftCfmVMzzuxhuWzQ/KC/hEO/
lycLO2ILYb9Skpt2UvIM1DEyde84WKDTqv5xvcJP9D4RjVePsWSjgN86y8E2Quwr
Rt9w6eGRK6ylPrlUmtrQR8sf87rthVMXo7GURzbt/PUov41Obm6GHPqYzJAnOxbA
YoiTN+LUZoubtqsO+wJX7ovjeKaKiJF/hqHfb2/nKBfuukBA8EXqwrhaad8IypRP
eR567eFPylDZzOtuyIYu590ti3x0l3DViSR+YLWdg4PrJT2PM3I7my3Ttqf4zRqc
5pqt6nVXOOqTGrPzbCHR3/VBLK/4EwLpMkBb2dxpEadr1En3qXeIUmDGDH4QNgjk
C587E/K/Wye4McmJ7IxR1D6ksFHcSyTldO0aIqpZOCzum9jqFGIsOEi1b1UqUr7H
wUdlzXal6lMLpGqCNQgEPhylk3ESmTLCzarVUW/ouYVfH9YhbdgFKP3b3852UbwF
zAU+oWzJgMVm2efkaTsi0Yfb8ArGbdB0Xc7vPzmhP10lwcHGuhDbMq6rgpvvy/af
NEcSlEDUEXcCaXSxQP+GGnOV9TRnsDO4loXfO2gIqRXaXlUvHDOtDpUtM+GdPWwX
vzbDw0zl/4p0Co/PFm6jD+/LPlKfj0z5BzinR6hfjhZqDtcX8P+jufm+uc0578c3
3Hh7aGAmYdnGV1l8PMrLb3p4VRb2JkpI5WGQNsUfM3AdB4gB6SsBw3sYxRkQKT4A
5xFdbG4/ZCJZdpSei6ljG1DoQJYJhq9nd3FNX2DP+zKz990d0xsqkN9+ig8fuOjj
OMEtbH826O+2eEuZ/dyux8nt/sAqYZyKPnN3S0Qp4ivPe4XiPVEEQq83hlpsWXvx
bd/tdeVFuOUifhJz1oi+xqiRJYNqbhVXu9Q785MHFPXv73gGMla9Kse0K2VQEO9+
zpojnVlx/Bvr7hJLiPfJkaYRK+4xawibJ4vpVyofZc4ICmF9iJce01or0JwBrCuD
Oab0AMX8rWLhQSfkwjqgP5gNi0/ykALS3ox6OfQS/2pCaRjj68YZZOApoHov0mlD
SgkoidyC1EHjnqGUkfM9v5SmXAFncGJtYoYIlOinAS5Zjb+S+pc4U2vRC4hD2WXT
x572AQXIE0WfdN1g7efMt3vyvzQl1nLjf9xBw5E2TwANGgUyTF60ONSfUkueGBPN
ScM+GECtVW3DPQ87552JYRws5FNawvdySbhg8Y7SOXcIsXy83vud1wV4XiDSzTkU
5cbzsgA7XtolrmgQta0Ob7Hx0EvdN0VWdzo/WcgGnFGtnX43vlub2ioOwEoz/IKy
ARgvJ3rRPrI7qWYtfQCq3HpW2FIGSZ5RgJ807esZuq2800QFI1ZzgNq+wxYMhzLU
mmenT7MD6vv/EEd3+AIkaBHpqL0B8o67N74n47u1IBmLtvRji9mRc/4hiUy3kz+G
0aKgfM6woiYy5coVBOxCAN+pUM6NHn0z+EXcvSE+zuwgI8pHBPQveXlCVeeHIBPt
GR3yQrFTxaZh7elOvo/TAIXaXX1QJz9q9T6VDIwmBAvMOCqLpUhx+esZKJR9cFDR
BRKRpoZgKD53mu/TBGUZXB3iYi3xKjfPjnPhiimGnAFRt/gY26OSid6ihDqe3Ird
g05yVIG6lX8/SCwRpryBYb+tDLEZWdNY5PoqVrKR6eQpeQTgTFrbvQvukXi+JBRQ
j+DAuwYDwr6JHys2FfBKwmbOJrRQvF8zdASy6g91L//Muv+qBQS8H4hiZaUBbUDo
vSDwZFbHTcaBCtasTVA862FoNvHJp09DLZGM+0LPcju1U5nxGXPxowokStt6+Vsr
l0iqIL3mLQFIa0YeC9Jno+SmN5+8YDierZW73iGwxePoSFrlwZkfNnbykUgmPs+m
StpO0YwpX0kwCC5koIPpBM//q9nXbEWe2/szqStMy7LmEriOE08Fq4ZamTafLgyo
iCeCQJTJeY03u8YN0eR/kq7H84H2P2P67KAHcSpwBqDVGo1qlM1J2u1YywcM0NoH
QU1LbS7rOmJSQUqC5NqUxJM+a3zUFiFLzMJR2b7U6mXAK/uXCCYbBnKKYuMKUrQg
FHuqtgxNCUNfb+HkOgongBTbkCdmO2hc22GjQSLXaIlE/j91MXlWFxUr1hkJAVkt
mHEsYkq/5oOzprMtbLRVHybBItygdeBzjoYPp62dBjXy6Fx/T0WF8Si3JlzOwDw7
fVBSsmr3VXOgFUGq2AHjTNAjp+eUN6BEc+ApDeOP4Bjdo7DJ0ZntrzCMu+lvBJsG
a0MvB3xIXIi/edqwzz/qh6Vya/NGLKLy8OOPi5aGi/INQBU/OQWA0Z22ZZE6o8IM
rnF0PC5S/rH3Ow36t2FxB3CBZdxIRD2EjGQ6yOFilLzVYEh0Rq+Lo4jQpnUeC7Sc
rzYpgjBpq4d45Po3u+v1tB5RrOgdmqk273vrx1bSngdev8R5tbu3UG1hSZ7AN6UD
N/p1UfIu2rASUFuCWZufDvrYebboE85pS4LqUHgX/v/8r5qgC0Lw6ADHzq6TijiD
UikJZ6ONOAvzBir0nlwfVNYFgf/RuGdZaZ2uvUQB/Qhja/zAA5znuB3Q4azcCmBs
Mv+JkAlYUE6DvfgonBnMXxD0x2aEneTpB6i+xs4hkqJlSmN62cs1Rmm5LlFxunnS
cH43Oh2WW5Rn1lYBDM3Y2yy2kCieckuA4lstfbrjVyCQD29pc8OSkdibDFQox4KU
OV45yBu5gSlB1YKQTV28vFtQIQO+tTKUYhYZkMtbQse9yW+mJ3dofSwOS+Mp5hSi
VNUT2hMuol8T8yyPySZ+lN71vYboNs//oCS9l5Npw2dFCo/R7kph77LxcfFqPd2Q
0755IuBlCJ2c/a6nMPesQnGcqdEsawlH6d7QhphfYusnJH/Z8WSkmKs8ftZ+Giue
JlrHbZoGg6EJuq4oEPqVPbA3lZeLa/ueEXhKz0KIp1+lAXmSO7CRdCglFAgdnw3U
kRsflIYdoOdec84tcpfkd+jQD2tWgxmFbgQBgVSr7Lg1SKLuoI5Ig7pX2CCC/07e
oE7FGml1WMzoc/c1cUq8AyOERKliauNYjkhG0CvqwsoHAu9Gjkyusk2irwjECXWw
s1jZDkyVHSR9/zdvQ89kMsKyrBoPjz8Q8/b6rRPUm7mKhYuxJFfo7Nj3olJnMptd
ZF/dfzwJZcL9Bk/PO+05aKQzFDEzQ3dvqO9OCaJoIJaheQXcA9Xgs3BzPo+4H3yy
8BvaSpFxA1rzomZoH+Pn2iq5n3EYdRsjTOs0qEuu9S6eAXIWazh7MDb8lj68WGl8
66PEY7GcOmA4z/2fabKEMonl8d+eVrJTnnzta+CJVS6UZSj3P74ZUSV/xMD970wj
Vgr80KojDsYYaUo2II0UTH7bQ7p7XSidcuqoQ+7AXeJWGzZ7CbnVIjTqWe39baVS
MvOHkdsXRjGkYTq0gJsMs3OxBFdoNCGGjYmCLYBfsrs+R1lTBstB1OIRIHkYOrGy
2pejVVQf05yBW+vMmzKu4bXldiQmBwQbpfQcEe2pKjnWv9+RlU7SgN6QvPaSlYZy
FcN4CmBGnEWpvkQyDLsRQ5yIYSium3P5qu//Y2uU0cLMNZ2PylKIfxecCoJ208iK
es2IL+Ply0yWn/YK5ZXO4rliL5pJ2sCffhmU+Q53+kSfP6/mQWsSs1wdAdwlaSFE
snM2V7xxouK2YzJq6LiD3/kTdLtDsnd4r7SiDIcj5VWFqWq+G8fmGmtiv9tuIWon
56rXpcRMC6Qpxd3vcg8OO/T9qSgZg5oZqGPcJ3HvaVrN79n5co7d2oDRjVFdhXRs
vBD2FOl1XGQ9oDwvnYzjBs8Am0Bi1fHxYYSe7ZxBAmLKmo6wm0f1o0A3W6NCL8mW
3pl2rxSDkioInPKMAq4IBSH8WkZ15ufNgVN/9Ol05VgOOc/xIyG94Q1z0oMwmSh3
C1bGRhQRqzCp2xnOGZYFY42Tc+J0Moc8N2xmfr++YcU4/nPybL+8AdwqO8vcxtzz
HbdJVyeIEsK4rS14zg53BV/i3uFWHOOKx5ao+jaJBkjd9h+nhFpbreR0dhlEg/e8
cZoquNcOeup1blgm9ebn80wzHUCeoElwT6gw4mipPatQIg83NKNjClccHMdJFzvB
SQ+g2W6/DyY3NCqjoKimio4tiG2EMwvBRK0ycmtF7exJw076Tb4kOeKFvA7uuoVe
nOqRM0JDM4zKFCSeqNu3shgTl7+kzujs28q73//3dISdQyO6OTh26i4Z8VvmLbfO
fyH4MWqa974ErZFqzLBvr3J7hEuUbN8C+PCWs2TE3ZkHbKEvlubG1tI6iK/3iTyx
4EyGZaZ+e3Edgc5BPf1AyxGTqEh/wWRPd7PnP3Q+GSyQYD4h2nvhLj13wT4YRoQ8
a+Tv6zcRC5M90HKYFOPtd6v1KxVW0//lkR5lpYsSkJvcADhq+cdPA+lzjqFEk6jX
2ll+c8khhQD5mmJyRtrQNYWOFnVILAguo6pBXAN5j/rudYNCPnHgpN2ouHmQwu5I
j5Jpg1zPRIhW/bGxdtSid5oqzeHY4oDJOwQt9E5fMfGaftXlJtXcQSZgLa7suNad
jKAZwABZW9Xyo7vykEcFIsbGgFRvyDzxc64AnVfHWOshaWtCJ2SMwD3GRhUPvfGM
TZMl9TMPHhJB/LMUNiCCf2t0vct+PMCMJkv1CzsNY/TiIcrAli++UvNveNIN3jYK
DVDQipqol9q/q/kwBYngMTLODJ7mn9usFaktcvEMmdHa9fBP/KNhoRffx+wRo129
vAPfDxVK+Q9wrw4uXSuTkcqPV8Xmbd0t1AYeJW9Ss+2rOTdEY8kPW6k5KU4NL/Ta
M/IbjrlGK9lfVSmdTYjOjpCUBh/J+3J0JsecrLOBsAWzB7f4fhThPErUom5aU+0n
T2AE/kB8dGzz0Xk+wmCCN+OXEPNTggo9g4JJ0PEnJu/l/Aqu4C8Wcg3axzeVBY/1
FEWJmcuJZN5YSS8Vc1MfAcwYOl2jM6OY2wIGF4pvSPGwHJxdA19TybhtwzLN2Fpe
dcqChw9J4Gumu7XkGiFh707x7GMjnyVP3vJlieG7ae6ZJU7YQSKr7EsuPD9UKFM+
DaJhO87u8quE49Crp9+z6aNEVtFkMxa4LyFl9c1oMsH1b27SqCjFPi50ZDftRYeV
XCq7zcEMyyaaVcrb9AdCnNA6ugRWFOwF7No8tBdhfpfl7jmV8t/j9bV4ZqFUyJVm
MGYg2V9qzlr+yaLCLUJkvqus0WdYrIfICJHDMrQpig7ebdiTZeBjZx7Vfj57c83z
6W5eXl2QOtF6j/+EeYl4ARFu2uO/iaxW0VPjJrjVGIvT9u/EX4kedRY+0T3xz1wx
H/7oFpzVMn+kKrC+L9g+fi6gztuGGxw4ax1jOCS3fRldR5POVPjot6DCKC1XfGYE
qgH90wbiukbYe1ljNOa88ACk0/rDkr7SwacIun9zXUS8rlIl3puBEvRh2t8Q03x9
VQT3M39iObzrQWoCI74VG3ici5uj3a5Y5KHnTv8kf+pFwy1XpthxOBgrrz9jsWuW
wRfCYfl9O8F1UYr2FobTPO6RfI2cke95JMxx5wgAVFafKHGck7JWAjq1n2bDLJ4o
v6NuxWBhVy2Zc188OTNMpVdswbkHZE79ywC4ANSiC5gVBQd+57Cm/ql/RSROwONC
PTzVuw4gV6C3haRYJEVSS9lFQokmHJzlIwBHqzZtVqeHS1ggcT9vfyGd7wgVZrWs
KVBr63sVKopL3jI0JsublXgNqJmiXvUVpYLEqMHvmYTzy+5kM9/Eu8ZlbV6nNVis
7ZLv3y2Nhe3k6GjISUgtrxoEq9OrwiPS5Pj9axQg1/g2fjCeR4WCtsN+skc5Cis3
g9v7AWrDxrKFflmaa7udjSNQLZCzJpTV78iNpWsCHp9DsQQ5tar2Q6jBL0WpNsvQ
G6nedXwQ/ueLMf9+HlX1sr6FKHeNyc0vukSS656x2nJmnGSPZOt+QzEIdv44jwf/
QNJfSLtVW8RfdMwua8Zc08fwDuPFEDvKEcnzAU73gbwOzlyygbaHns5a69jMA6mL
TWG9s2P2v1QaxeQuT4oOIln0zAal0VQWNgF4emn4IWKbM/CrAaUu3yUSj1UE4V5J
rE02lp31ssmTKyxXDuKd2DnCdfO3G8gbPVSDgRUpdlUd4MFy0ksjmT8t+swXbElF
MGhz3uS31Rvu8jk5QuTWUW+jJWdkmfjrtWWn1RUDqqYNRwd0piKWvqBEvevi/nMk
5r/XHm94mYmqK6PPUerUmPYTnDpW3f9D9E+DRUytz2grnr3AWRaN0B9I9Ie+Nwkp
ORxj/Wdfc8xiXBiA3BPLjq16+z3gi7fjGCTVtQWwbCs9z6IhOc5JiYTVfV5qiHRk
9+U7U6IekyXgdRnOuL+Yr+eXPNoa9AXz1Fc0SklTwWdUBMcGZQt4GYSSJWVFbsCn
he4FKq6P0ZiTprWKM+2xddvPXAERy0qFGvi/FPbxJ/7XjBD1LXpbD4AniVdmcLeO
iYyCv6GnvPsSTwNvXGuMu/2SRmrFxGNuVjQZlO/D5cm++Kcmn/b68OKg2dniS9MX
OEBZuHK26pfJfHwz05deA7zU7nKiUbaUedsU068rHlbhMZF5ZSCVKfie+has/nFY
HLkf1l1tp1pF5w3pjLKNgROYQRIBOAgjrkE4C55m7ckC29ziatTySCfmvWk6Psed
zcOFbLeuRqTCuOEz/bAEYvRATMROAufV5bLNOvPYK6/AN+V26fYaZFQKVMwuqwr4
9r+qgYbGVFDmrvE001e5SSRRmBWp2VBPJKz+NIRzVdrgoYF9qRhWoUMWD/YNXrd0
V8OzfuCKyWYBW8CQamiUmezIAEvVa8iBf7jxMM4L3O7H6/TewFFr/SX7f2JzkiT7
Jn3i+OaSFWaEIYj+kxsbBqfaqZ8J6yfKE03d8nt2yuKDRA/L2D4di9aD8GszIaMZ
tqADURPQ/fRz7cVl3zbBFwjKHzXdi1GJHxAFDdiyMZ5+WFIZr+1KGFx6V1+8NU6P
RTJPEED/EkNwAtAr7zVl8PVhB8ODPStZ75pqRtqj8UL5utHNs/0nQKFyIS7+XN80
VJqm0lErt4nWxIsjKLEPAc0qskth3SifyvfCPfNisGrkwGUk2X/3YR3+4Icu/Jfe
Md4VpUEDMILhtUIFrN1FrSBKI6ZXbP3Mdr0FmebJMkZ7zIyj5Mk6lR50NqISh3Vp
x19tq9oc2VkpGLWJ/2+p1+1Ut3sYm/gfBMyxa+u0VLD0HgbAyaZxvmBgKjZUukxF
ifdjkPFvH2FUMpXekJ01Rd4jNKUbX+hSQ/YK7Cr8ElHhl5ZaIvJrMtyBTnYBTOOy
z6e+T0k5RYspQT3I+Zoo6Q1HZqnLzIx8c4168yeCtbwFYRaOf3P7lkibNkNkkI1W
98PVZHFIAhoMb+ikryh7GCCiEFnolEKI1TRPHnrWt/OKrJrdgzZcWxAn7pa899uq
RR6/EG54+Y29a/RBpSvaQqnjFSkLAz3aSLIkBSHkCYc8xtCeH5V8W7l+vy5l99oH
P+JRppl7m1F4y4jRczkTtq2dgkRwWsnsgnBbV0QfItsVMxEWhYdj0wLnfr3+OIPR
+PiBVdLk1Cfh7ThowrSRmK8Et7YjxDOpfrTdhVbFk3eyRwvHAx61G73IVnc91FGQ
xTCHIjgFSO0ZYrALDHECg2b0SztlVr8sotGgtEE92W1mylqrCXauoNrqQuj7DDYX
hmHZrtOTFqogwO3z0vBe2WqG3EGzdJnzClBIIv1nYwFrOj3XfsN34BzhZQ9kCbkp
1dDBvb8VCxxRd6xmrff6U7xScZOKZnx1aJ0MYpLTQwOsh2/N+XbhzHYTYvq1QtCH
e2up7EkzoBsvz2he0GEaYHuy3+xWVJThjqzOxYF6TuQoVuoDfeHmACWeOS1CcU9T
kSlu1oRiquz6GAPbOwmW6e8B+Pd3K1DsQbF7lCVaQmlsbEq42V7v6adqBFnEzjco
bG8SejymQlo3Rn4vlROBYULaRaZsYoRar+qGwRS4185RoLiqWtvT+MVS1yWYpUui
pE3VDqL39yJXEfRjDf0NoiT/nlFaWVFIaQKsTxic6BPrqO+WOy1QFCF6rsnkV/VG
/79kkqRWn+8g8Z976u7wXkr/4Bykfa0kw4KnGNOb6f2MnkZ72Im2/RzNitskbBok
NMqcCkvdr5aO/dRXFZUb57EppvOzo0I1GSO+AbkITL7/Ba70ZRIJ43CwnuGCEOae
R+tsvQdpaya0DWhceDQgto4GopXExqAhQ97lg/xprMeLSgFynTQmow7lSqIMYKh5
9PBgPjxh4v9N2n+yuVAWbwiqPGCpqmQFuWZI42n8c2u0OAFktGp/9//jFZkooSDJ
LeyfbdwdvLij8eGOB1GVr8CSmKYR5uha5Ntjpf+L9xDsJrBhAUmp0Xjm9Rgs5+sJ
AC0vbXA4kmRSEHqur8VREdOtAUWkgoNCTZdIpmQZRO8YqR0xKBY+f3ubRYDBvr1h
ULizpgDYvpJk35BeS9sknd+5Zl2afY/eDa1TVut7GaQ0+YaUkUHA2ifkf8AeQAKb
OVuE4QnqT5bG7q/6wqnvA8vGiFhp5jFsX/RmB/FxEhr1JzxuevTcUWRId2ze32+/
xZdZevyH1VKlxu9+uC8JqgM9M2QlbPydg2sZwY94azVlyjYFcQwgHM8oMA6fDcRj
h0wfEJwhyaW+6jM9l+a1ZRsABCdr8GMSsT58JWwEun+kQ90IqcQWnFOxuySMe2dd
KgGB08gYuw6MnnLKTsutzRMCP1CwxTaqRN4q/pWSeKHWyFC13BEJkoie28+mKGsl
IjPmfODtylbWWNmhb4J/lApFQgpMXQs9UcSJzKMNR0sN1Hovg5lLwfb0C2ZenuFL
MKM/jZjDRDIGe6mSAPyAB7yr0zDFtF8ghaGYdqYI7HBrfbmC7NN+P1TEeHj1badm
RnnygZUPG0w28z1jvQgy+94EoNHjMAwEb9oPHxopwbMfqZFf2lrFYBgGufyMv+1b
25dnsdD7/cli4LzrIiq7l3ZA/ITcjomofOy3BCT2Htl9K1Xfpkqx/kmu/vRJ2g4f
sbRvRHmZowDj/ij7d+0ST59BlWGKAbaJjVNEcc8VwvV3hcX/AkNpsUYt76jCqdaY
4QYcYg43q8ljDm1TrVb/GnaOL1fuDLrlPEdk3t+DqX5wUXc614OoC1J/w4fi4JaA
jXdmMGMRH8+SqaGcwD1LtSA5/UOdPVcXZKkwqB0oR3iqZxeIcfYwU0Y7jkxST6TF
nlbljxTTAciQkSm352u1E/NqmF4GZE6xS2Nv3XuUZ4LoNqYeUGdECJd2cFHS5Fpc
WFUbbiLAuF7dFIRmSAFY/hQ3YohthPBg+moct51wtsIoAQIE2fCgXqA7cDvOHomX
BuxJj6OBr24RH7lani6wFedtBZDHeRCu89JExS0pi990ZoSRTpaAugInRTIKuy0l
7v1jERDdipxGAIHTOOqvadcp3PN3WhCCs/jsYGlgXXX5k/m6rT2zZwJOJWkpVHke
gJy6Wf9SiQvAjovHfmvMGfLfcmNJsTrkpMr6VWjLowWLsZayI4agFzFC4XhHwpYF
trSIg+YZ1bhl5J0AUC3nrJnzYXgutAlbK+Zfau4cFSLPaRqLyirCGsmhWN3nknSR
HoWFmrTxunFZVXQ7ptSuuJsqA9YKCX6tjkEJJKfs6RawqhhpgbRJNjzS1x5WVIcw
qhFPgthI5dL847n9BXwWWeMTlage0oXR1eKksdkdCl7u1yRrCQMHtLGAliSavsio
etaqHqrNSGe/NlpytBcFHnQyyErmomGklUKl/m9hmZgpDPrA5C26yuUkJKddTj9O
nUHIT8QsLZgQ3I6ulp/59o8XeqmwtvDpdbNHk12PW2z7NEZgHL7Cif0ho/yW5IRn
omIs+1f/AQ1RRt+Y/Y1HXc5hFxV5Nn1hjCftn8haeXvkFiN4VhbqmaMk1RK+292g
rW4B3XKNPyRPDhlQnrMddUJtJNPTe482a5AXpZYBdv7yRVSi54zbcTNmH+xRTZ73
iLFqcpsAdqHQTNtzMz1fYwOaNZBw3/VU2nH95Pu60igjpehMDCdozjsjl1jO044H
wEfhvCS01AMohn8VSiAFUsVyMo9rdJkvph52DbXOQGwvthHwBmHqBBYXdM22XHus
Tu0qkYgVNGY77IbvGpemdnPJK36m58W31iHVRkUcwmXQj77kEE5XyHeBeTh5KrOY
mEsVBz2T0DVmb6ioxxvK9B382eVojc/uXlDcrfjBQrIn85sXpETASZ2RrPmjn9RF
OG+0Sd3RQuQ+MI/o+DcriufVdlHxbNOExLZTqFKcg1iNYNEW0SNUDBUb2PdvDZrh
iMtbWSKWrvYcB8mWgMk1J/JixW8KEJNZ5kKkhj++j4Y34FEHc8Xj2kHsAu2miWMu
8KQTh28YeEHw6n3zf1mH9QrvC9aSCPgn9y4UaC9zy1qaCF0ojeEcIOVVs6hOIgKj
QZEKd8gjyl3LP3o6LEDmymMYCaCI8OnPC7rLaKVQ56++JWBFi6wuXlMuIuewKOSM
94wY0Tin67SC8tmmB5iO/ydNEO50lVqDMJytdR4ZboZoPjdQRYkwRuZj2SEwbwXP
PMV8Wu8b+cQyMQN98HUzRJB99ErizoZuol/F8gY/f1FlzDKLvZ4I+cnW2w1yTEkm
mb/iaEOFgQkzvbh/2ZUBpU4LMbERS5mnkUkeiWy63bMvvVdNvwxaNGNE0ckFTp0k
TJKLWaWdiODHWqEQu7BM0EljDDccDMXVjqElXppxCUuvwYdHQXW9XMEJ56QqKq6F
4m+8BeTO2ePjo5OGbsDQaMFy/8r3zdnT3YZIYuaHwVeADPIUPSq5di49Mg51ckQM
G7B5BOdFOaJbeo4R/zSrOzKWPuObz72Gj9U4UmamS1RdYSaJKAZI3QmCfHeSqE9K
0WGMK4NSYFb6fmRwY9ic6DSC+yYoQ/Ypr6P+xPvOhn/tIqcB+O70S3cIyR9wFObB
eZVRjUMJU8UWW0QimjXqNZSs+Wh4IOGAgWz8lp9cmcVuyNSeaAhwkDoSOcycGx+b
cr7L4nOiOcVGiNIdhKlr2el1E2MI4pigNgOqpP1c2EjPH/6wBMr2p7VD8GLIwjAP
1WEK0aPNqFMgayIi9MgOFgfxKD1IZouwZfPPLKJKwrdxPZgFiGnVTLqhCgTKXA8D
BD1r02ltZitNZyzM/pT+I6srK+jyskwRNwoDyBeA2flN02VsRD7bUhjzf6lkOXAZ
RmXDEk0+MLuy7z/2qVgfHx1BTScDOrrAOU9qKumVQE/4P5yAJTPJCt9rdLYAbEPu
0mWoKqciVgvjFD4bSm+83oe8nbe2C2uXQEJ/z18NVEH3ujzdST4EXlAQH6xX5PLx
l4TWQd4q2laO7m0+yv26jjtqrguu3UAQmHC1M1BSCZTnqDBrW94ZVFNEZgbLiS+R
yqLb0RuZC4zemQSWFIbw9IPVhb9wNeFQlVMVh7z31s71zGKQaOW4iEfmpnve1gWo
4mhTMs2i7T9fXaH12VqIprepcTu81STWMfPL5JSeadOZ9CMjhiMHmJEB47pGyypo
lVt0b5+C2p6+c7S8Id6tB8LfqCyNAzttDJ+kCsNSrpihuEkNhkxd59dpyLn+KaG/
S+VGyerCkfCPLbx2Ey6ylnbO+8/4Nx3ROuUOtHEx9TOvCR1D/ObzJN+T94MB+aX+
VM2TkJr+JnfHpe2rzOIg7J0XBzmPmh/kyz6hNuPCVsrjvDiOGdxm9uPAh482+gqp
5n0JpNicOXCFZd36P6qR1/E6tI1FC+gHwJ22+5MaiaAp378LS4OxULjIc5/VK0yA
cL3oXtHAlOickdm/4Yms3tqC86w5hRD4JCfQyu+K781SZDUdYsN37QhFApvQMsLe
C0+foPWnqe1jMfpKfYUZLswPiO6Itgv2/kRyhRYEeIBAo5kiLRGj8b/snmNZxnp0
hnrh0Dc4T4FrdO4L90m7L3dhHOD7ZjPLJe373nTjCM+Ltr7EBeEs+Cr35MNIzN7k
iPYS508szBjUS4wS770Wo5bg6rXw4NemASI2w7jgfL5comuGNnOQpQGN9x60eSDA
SH/gNik9xYk9Tl44ji23ovscwgIHdjhY61vqFm2q9wUnwq5Ddn6lqFyzuuE7krXw
mwe6j5RDgeADETEJYbsrYtZNUambBG2RRityt3vPlT9EAVVbMMgk4PFi3fWtFlFt
fem4hFUzmSTSbd+6EH5ejWn7LyYLQoJZBVLxv/f+9gnaxr7GJ/js8krCuO0NS9J2
dKV8DjLcB6h8DvUAYjmQX64CMuihQRtCIhGW8UhU8N3Qbnn+rK/duv4+GvykA156
HSyn4iWHF8e77PDgP7X4SWzideL5rGKmLUsJDCZbAPUsfPxKK+yU3oMxCLlGcHQl
Q1Y3nyPRieWKRVL7pbxTMiMImKrAcA/CCBDY6lsehmsb2wwhf+uokc0RxCUc2dGt
BTng0Si55x14oMzkxZMpzH66ZiXLBk7LLjSNO6hfjZSrzyxoq4+mu7YkMi7Mc0nQ
zDYcDMYt4ITw606q10df0S/vyPaqiyciGX/BuYDUpQ4w0C9g79jjOkZKAuePe9i1
5YvuTkfH/o9ofjRYluavR2MDtbfxwwdTrFhN4ckrsuSwEnTM+k3gTmZszwgtNoXG
sKifYWJYKdBRuEmg6Je9Ul1zXpQAVanWW3P38rKPx/vqpSLd6R9ga6KEd5SpS41f
jBC6d1TLQR1ZF5WsYlGETvdzyW7/bqGQB7klFp9ncyaW8YkqMM6UfZKrxOesOo66
a9UyvHnVOiOt3jZ5HoBNrxSgkLHIsSfQeIsjuHjzKvi4i2pSWIFRcG9j/iKqd+L7
qy8htJrM1iOELFLVIHurYOECqMs5aim5TMRyVP1fHk8MFS9r90BdeS2ieSs5LqhB
IRjqeCpASyomN9+6wHpdSrW2Pwzb2iGgPlTzZNJ79plZxiGa64xV6cFIUiT7aDiz
nxyl4LCsrmTWXEzwuiNpT/KJvodDhlchfXkYnK733V8VO+yWpmQBKibjdDmkyq6+
g0KFMCx2zaMVoXMfirWujsy4xbssQm/TQppZ5PiTvVp5HPL336L0HfNSKKx4YekN
t3wPWhIQb6ekfRndQaktVYrSO+3+d0MB76/MryygRKGhUD6ZPl5IBpXEdOY1ShNz
dhHaFOzieT0yuN17ityurwDDaqA2ciBbiyolYK5seUiMJaXco5PtX7lLUsgMdXyf
W97Dcw6s9YupXoXS/iBQSr9IEAe3xUVgHEaX883BVfshtOwxhhZD9IbX1FhIlEbu
8mORLl9RlN32BePwnczYijsN0+r//prU9ogJSWi7fGWKTxKGjX2jF8vYP7mXQvIE
HiUGILJ2kvmDBr8si0lNHWsQTMMBTniUdZl4rU36JKnzX3sFPohZOimTtMNNxjs7
xZ2/S3pR5+yKbQy8gPzGAGU3hzSWZSTL1gKrx4+VF8NT1m5v8Z2AVsjV7gHqdMuS
zgGI4XfMb7asp53dTkJ2nNFyNONh/3e0UAJb7n+GA+HtqNi6qXMh0H2JXN58kesR
rBf8e/djqBrKZL7C4z0Cy7GOR0JN3Mfja0c03t0t+hXiQ82K+5iFS6Uf7RizvIKy
A2WfDVj1+ffcFm7ri3XPj1/CCDOESNJJ2NIw80mZAjz+kI7qpIOno4GaCkqvC8sn
OY1zRCV33bqkY0lZpeHy233l1fOf3wOZIAarofy0Vl1vYLdxJaGrlfbeoPg2MtRc
m/fDrl4ErPheQAjsQ/jQdGzaAiws3v4AO8y7k9JsuV7x+iJUjy+T9WlNrawHNb9E
dDki5eFml17buq3eiOOZRtXDsR4pOMbod8UhgzB3Ri3ggdP6IRwwZ1UNMpg/AxYv
gAK+toIRHj5A8vaBkLLKHiK9X4uwLcvxSmA4ys/8Lpb4ibaWDs6n4nTQ9+r7tnG4
nn+JDmLivUFkUeG7yPnTk0tpMRCawrmbjcLubDbaiuyKXFzIqaFSbg7WaBzWsWo9
I6bRt/vJZDZXeRltQcNvdQCqQrKDbbIrJ/Wn+v6mcZ51UL8Ng1XJC839tQx6rgtp
0lRTMMH5DX91X9/gaHq8zTA92i16TU2Oyx0brnEUO02NG9nuSI9Ty2BOYW++fEgF
2pxvuIE4b+SPvCUqpYtVZhUo0p0kPOjAqMkEZ2IGMNDLjYZb5TdejEy6IX9Lw/AO
nebDRjm8l5yxHntO7ba+PHyxc75mkJ6EdXTNnV+qSjWCKASycY71syI5g9SxxWD5
PCmAPIXd8Tezin/9QFQ8gaNNRNfc13cxqBFST282p1khn3xc3l3O3ePj8nXnrUGq
AsfDnl1zFz1UxvqCuNDa/S7VykPPtTO271HwYFtbt4DwCwTqd3f5upn0UqbL/J9f
zfCvQO0MkWMibNw0pvx8P5DFUccMKL5uf+CqmHWoFNkJVHNDaXyc3nIkefRG5Kby
v66ZroDF1Ht0jRfjDeulSXs7FcXF/y6z6TdMSoX3csAHeR17iBLPaux8PYJgJ6l2
/ODbUrXogz+7RR4gS8Bh4t6npelgEI5sWk9plLV2FYlJMNjJlBgnl5v7opzAx5Tg
BWPT/+RexJydL/UgJt0JqIq61vxE0/ToVUOvJZDOwJmUhGOvX/Bkm5IS5lHkxLvq
+7c36cQif2Ll21i+dB4y8LDW/xuyOlfnID9FM9lNaVikvOQivdb4vJL7pkiE4H+S
S+rQCQR/vKLxtyG/Tkn8dhIo+MHvl/jcSgd2EjfNsbcE6Ew9opP9tRGGiUTQsXyY
iwvPQRtYsP6NKQCvqIchvMINQhs0zIg+lNYOoZPERlDkvA/ygM+AIQos++yXge9I
a6MlDl9GCJo7Z6RQn9kup6GvO0QRbigF/Vneh1UrnZbvsiHxXBxw+HKpIb5hGUa6
ZzqTpox2+CSufB8ZqfpOzeLSlYLako53TmcQFbFpnmTq54o+vFSHcmW7BZMCG8bn
EszUk9j67bEGiWIIv+i6ESLIAfaJ5j/eSo9I5zv4M59UCStIQxJkEW8S+KcuhODh
eJw9MaEEki+qBa8sElWB800Bz8dqFCeDu8UkFnLBNPzo6eTH6f2TuwsqruJuRPMn
vsVRyV4CH0K/E1OEC9WHRB9dewANhav+S6a8+o+fpH8YYlYKAaYNCt4CHcnPvZ11
kn/8OxCPwA4AsOKnmtt/FH/nN2Sy6wFE7wRypw7nhQr62ezTV8i8a+NAQyYbUCWI
WAckxE6sWYBinbtpI1lXDk2JvSNcOCZAmWf9/MoR0/MjEXn2noyBqF+E96NZN625
+EvAoYNIlxkVL8M3THQcrms4fOlWloHqSmVZsm3z76xbTJFRpltJ0uWtYo7nJ1XD
eH3XOQJtbk/Vn3mzJ7yAOvRhvPxpStea7gj6rKS1l5CI2JOk7R6R2Hu3U73oSnKV
O5AiS2hdc2ZSzIHNvyoDAtwVhf3cWDd/eB4QVTEtz/mV4YEGBxiNd7ps9mCO1y5Y
N3FzCj+XrEtkaPNAAZltLRI/GYRjwuIJVG7uwzrj2uumVR3DFIMRWIgouzmZAmHU
P+qmT44I2dc9TxG2qVfwtMEYgAD7YTFoFlwO2cnIRnSEAl2dbbEPXbw3U5Fe/v2M
HmWaRCk1IGH8akggUKAxZTGza8Wo08YL/sNuwajMBBm9zJeXxAMQmhniUwOpp+0J
TA7qkA0+jdLZ5lQsl7vxrH+QudLsFRMFWmo5liMs2YCQLbpELmql/fs35w8l9SSs
l1zUdf3B4qk6ui7+c5QBuPnzVnG2MpKnRenR5NqTBbgspbjUysVDZFhMTynLVKKf
Kr8PMoAgv0u2+4YNCaL7eit8TVhkeWG5+7EnRCIhFEklclKTP+qVf7b8/RxUXrJP
a2xVNAsHTA1KUslsnTY7EIEL8Qjp6FvhVyCsw8TCTDdP4QK5NUBgQ0w74dYSpaAA
HdhO5KzhlBHEIhGX+hlhgZBVMg0ySZfEswl6GspNymAgIQ5T1gcQInCgylE2h1Ts
MNKur4Kl9DMZW9Rfv1xqJKog2mEE8OB0pRSyfPevi+MdMXjgBtD9i9pMLFzsKm1l
WFDSh8o0dQlFD1qiPT2gzzOleIXjPxjrH+JY7jHsePPeK4OyxiHfFuphhhqgdSMy
RtFqwTxCYC7T1482f86lk4Oqq52VC2Q6q4om91SYFoh5r1RvQqMWMDq888qZtdZm
sb4duvYMwNorbWomYtqDTDhrQdaeXf4/cVj3rgto8YlZU+S1ObwyMaBcYVGu7Xwi
IJsGtSomuuGTnqAsvzKPz4qfhAzrbHBiv9cYhOkDEuxEisjq1TUisJaHQFZ/zy1y
8V0S7fWevFrydp5DfRqKLOvIPGMw1x+R73nCy+6hl0J+Sw9ckVWIACYp4R46o/Sd
bdvhMiObBRrVC9Iym3gGVDDRQ4tiMwTmub8tj46W3EqB/xm8aztLtkL9xdRlO9/R
PS8+dJCJM9jb5/f9LLtTteg8jZdKLoDCNLuWwjWD+FC0tZr7pUZt9VvauuL365E5
+ppDpwbyrBVieQxD3BBoUWHHuIC0EkbHRaSP7SLiywWMcLBGTsU/FMzqcpl2dXdo
A01lXAhqB7l/BvUuj/KwMAF3smWE86VN6+1XvYKt1gT1tF4auaf4e4OoOsdpZwis
//OOM5U5UL5uz0+Q/TtFiFwmgoZz/wJJDOXH5fqpFhSAeAZDlwVwpMZWWtJqYI/2
8IqVPzdbB3koVE/Yd5QxSo3oxFiU4m4N1Uj2oE3YogE8NqBS6QTqypUMPVcXfteU
WjYY1INJZSXRwUrKSvXlcdpAj/i8Xru6D9EtyQUBVVjmDkgGkKDN81y6szk+TnKO
IsWRuKAXlAMPt6mUV6tL4Z+y6B2/BGM9T0EMgr1apniSdsohBIOAEKXDz7DhB8cn
+CKUY5zkmx01nh/EDH16Q/cDttkkLrN1Mq6ijNHBV9GlI/Zibp3sSdWLhFDA7+XR
b9O2ideNFMykOjeHRNBGLzLf909iNXm2T4YfoClLPfDo5RUfDCtVPByBqJaY79tU
socf3TBqTii4kIfEb8+fF7bJDrghD3Z0fh4aMNVS/Tl5I/jhkABxNcBFBjHeFdx+
qrJQZUAkoFczaYxgakVZJO6P+6hwiNuycew+az2IL8asU/oy/cOk+BzXFwErYSdv
IX+C+ue2a7ZAF1cLgx6/iriZINK4g/2MgnuVCiHl9bUSnqSE3eNupdMKsK01LZps
Fm8NJE09zvHuwZYjc2gmG/HTtZ7KIo/czdziNtOlMBoGcdD3ukcOzcbOnNplSZUK
ss2NsukLBPE/8LKvd3uq7QWwooZQcOiIpNTVtxD6TvmaZt1xZvW26OfPg324ajP0
fmhk8Z2WoJ8u4zheNU+4kF08it0WjW10ClpHvyoTlIO4nET3CSXun8cipmkbcdsR
teDAz2EBbDPZ4TBdt1yeh5mQEpFwL8gb7YEQJnBwpalTTwIGnDSPCtdmvwSaUK4N
fUl7JFurWFvL7mO/sBbgTOtou26bv6ex+IP//+12IXM9N6L4iu3kTdoGbahq+O0q
1z1EEZGqIS93Z7pBaE7oXUJ0/weRQF8SS9UUCI6JsO275007F8HkxDEYlzn14/lF
KCiY6Dtc7pWjl7GiL9jwD8KKwJNGW2qreOMcQk0wUWceby3VJPcRtwKtabJAlgZi
wkIyC188q7p6/5Ndaf9uRmqzs0W+QSUpcw85UfXjHBNgi2ioe5ys34+VO9lD2G2x
FlGyybFgWA1nX8xQeb0ivdTO33exguy9EHxEZDMg6g7Fmq4G3YOvUwPftpBU+wxr
Et+qEGx8WNcbEVe2uWJYzp+CkX923olq45Jv3X9cYlu2lMD5emohDk6zuR6FpoBa
3MMwi0ouL0r0JU1o2mTwW/9ujlJyV//ycaMAsMwal/i1xyKdQQJmPggODEH11Jca
lAtKWRheKLFiIzFQENTAxg5BBnvlZYh9To4jcUOpUVzbgFuhtL8ZPrsX/JB6c9j7
n4gX8FY+zCH0Ib8+IT6VWl1gda80iHFBYNUZE++HHu22gSbSUv7b8AD/63NKdv6V
/wYafD7A1GACpHxDYJ7a1Y/iO4c5sdIz1bpM7mQriLXcMCiWE0tH/a7x1QOmRImU
07iwmeAbCVDD5xx71btN5n6eXanOPdmRMv0ZS+ss4f+OOqzRSqKxA0HwgSJvotLJ
pbGJkejZ/T4/TvQsEE4VaEZ3zYLX6/CjktcC+zjzYasKErL11EqxKKiVZyFKKD+W
XzsLkHoAYbZaROzf1WjSHKtHbNIqFheC9iyuI0BhTquy/gwvV+YEI2YgIF2N6hom
ViiPY/Hc3q4w8CkZrLTNOpys/3xkv6kiQTRbhjmjjybzrlu3OtCIL+oDKYFTk7+T
lbaB4J5m3yfkkTxAM4A91H8Z3X9Nc38CtlzxxU1oTO0+M1oCNGOzDhpjPu8J0afW
ZgefWLFfcn8zrYskaI5NNm8LvQl6hVPCnbz+LtlY2RwfzmJkmSIURnDKzIjWzuTe
VridVhG1J5lofi4yrb21bn+eP7/JGiShehb6kFksmUPiTwNU2hUTOLxkHU6ip/Up
w/E+ewEbvGONXLhkAFDzxRDGmBEQIws7VHlzlOIaMi5mHx+l7P0/pPONfgO5R8Ly
cWM/FuXU009VLbb3PH0CAB+B4CokJgIy+5Am3EgKxGAkOLy9WSpOEDYIemkkuD4I
6tvWK+EGsyZefFiP9BqO+ojEuPG9adGAhPoHkGT4fO/y+j0uBycaBxnVJuqfGh+J
AQQ2JIsY6kAk7aTEDBPAWPl4f1+Aw7d9CgOjK89bhnNhJCoVLGr1CZACaUL9L7JQ
tZrifkXzgtc68gO2eWZVt+ml2VjTcQDM+yJd2PR/kBNQXYsroDlo4x55cnbqj/bx
4/gTwHxd94UIElGLRFebfFaeRIUWae43N9WkZogCcepP7URec/lCQ3A3iF0wpi6k
7nkFxzQm3zGzpJcQZSfhAgoZ37q0/CC/cXQ38E4Jx8RudE9jk+PDd2cWKjsHXTkn
1ot+xYFG/pqmTh10BJ6ljuK9KjcV9mK5/I+xa0ycAq8OIKKOpqWn5KiPdTs/LCVD
KgozNUB0B6ZQDVGkhsFLc+nnh+MZlRn3y65G2rVs6Jp379jA+oy3RW9VU/HStTm9
rlYSibRoFo+kSP5+uGNUlRPIIEWvOjk9kVN9oL9cxWxTSsNsRzNXbAWqchNlrWvG
GohsNfPfqMUvXD9dfeKS5fNNA+EXruPnHRxwkK24ksYzvEWUh0wmzELM8rc9y+NG
EqLJttdLwd1XtvvIN5TqizQTicbP3rNgPL7dqveKAk0WEq0WifePvIn2rdxENIGi
ZlRvMb3bFStDfkYOa85BpcKTN3eC2KRm0OzL+OonlB77FUmGjorrxlRi8iRINiS2
yzOgM1o3NPN2yZERmNiYR0kA+I37mD2D80v7WF5IrJ4ExDoSXcKCA4tbJ7IsXPEt
ShOoWWlkEG602lCcX5zfain+g06+vA0mxDtNEVe0aAamsF2/4/h927lP/3wWze3J
npZjiaXDAWdu0AiXD5Ov+Dk8VHaeHedCcaqmIle9s8R7PN7UCIs09y5Njd2LtIjj
eLXRmhIR7i8ZbT9OAWpqLhymjWh0DXZVjQkwRD9ObBEzSgkQLpE1OljbMdlVaDju
p8ykcU1LOIXqYXH4UzjuT17rG3cQdnuMlAPPIqxNE8sgssvaAJ3ClmisEsdvTJmU
8E/7C0vm8jfU51f4XYCFRjokF3qp1kaa3CwomPMqZl1EgAELuacoF95DJieMOkW/
mZo7yOGd3PcMZMQxQepxda3DwmkweAJk5ZtEUq2vzBHfZjSNkvTnSHT0uZlZ0LcW
xvj6T+ouPcjiuTxdoARQQATeG/8YHU6bYMWy8seQLvCAUyr1oQ3C8gbu4Pcbkmek
mmkDpidlpANqNfu4eSxXf8S5kIIHDVu4h2ra221zuEwR4sqefM2kgRerYEsGZ0K2
+VX9Kcr/bDTuqu9bZcdGtnI178/eGon+OFSzvliEB+/WaX0LuI+Iv09NIZ0X8QWj
VoyZJiLZsR1g6dCy2rwZhJnSY1ypgZRdSlB6cPxuIvlZH2D4a1DECKP+mlq5gURP
9Jd/bPvMZ63tF+P1A069Wnuk6z6GvjtFQ032YW36NPAHL43hSoT2qEKNhb/ReYuv
y2Vxx56KU9vInFl1GjtX6ayg2342eRP2S4PuWu54VlCM6TSlxEYVRUNlFj5c+j/D
2x/NGN3CENzMwrP8jv1iij6mTV6Fz9/U/9V6WBuOZop1YMf2olVrn73p7iObWUNQ
8N//s/WmIQ66sANHUoVS809JcmtNZE4AF6Bitq/Tmos6kcUdURgEfpG0MO3kUG8I
mxRSbFeboW9rLX8MK8bgbpS8rib3CgUIq0y/ZV6lfie3t5qhwedZVK/jLo2RvLxm
431r31XyMCA07WPHPgH3mCm5xxtdsUAxs6mjxc7KHxZGKIgTq3SB4Wo2wWd36ypu
3DKeXsmg0mHP1HZTAGaZYq5fKkTlwgrAd4Oc69tf970X9FfuYht7Q3rAzcCvUXaa
6Zc2gYWgLBpo6DIGQJMfrTHFWH9NGvz8B5SyNYi5+QmpV3a60Yf5lfwbUJWBKzCj
zR38FYdStAF+9KZEcet1Ky+xNMcUbkXWGGH7zwdFJ8UALF3+hG7IipBSWay0RHE+
3Nyet3Un7TFnHL1PeJYWAlOy0k2+1MNlylChbzAaQE5Sw4xliCUBYO6X/89cS0Hp
4cv8H1M8O4QbX1tel45eIOIhZ/NCQleBWzNZur5yPUc083tVZhwpNVW/T+XfmDzP
p7sNQWs8Rqw1ONtHw2Y/dtG6u17QkccTXk9EFmuilWEOuCHpEIRK8DfGY9jDNmzk
+fICx+IpclhTJ5eCl4O3BO8Kw06LQZRLC6pCJqCPNfhWYs4Uk+i630qnP5IfgynQ
5ApDPs94005D8HUhLO/CXX6cldGz12Z8C5eS+v5gvtwRGgd5PI0v6nnaGWq/V+7m
xI/CAk1gF710Z2CMKBiEaiMdoRON9MX6bwpKEQJUoPO168J8cD4K7vzwXIcHg8p9
D0Xi3yejB2Qo6TpPry9Bhyclr9YTKaELl22TF37Bxm5vJ8jlVrNAkkXhmCXUIZWN
RHEQVTpBAOLm2uje6RXJx7zQan1kuKgUty2e0R3HFeGcYWfcmwME43WSI9og8qvV
AJb1No9qZ2Hxig+bEVSyOFAkGLfGMErr4h0lzls/gnSLOrGQbSTO8MWIqMQMevwY
9le5Fx86VHzcTyGyXpHt2vrEQNcOV/2Ka8/GzlCe4kBjGgPPfu+KVs6fy4uqGnS+
dwi0n/PR4nPkWUW4rmxVbh2aaNAOUV3IUb4mGBDRXgRqDkBL70N0t0gXqbr5VsW3
KmSFzFGb6U+O5QfbdIw5q361JEvkqEOhqXQJ6P3StmlmL9Dfh73WmxgwUaesn3Dr
YBdGOSx0NYHLWCv2EN2OsB/LqgEqet/T1JVaTO6jj1g46lMCvpd8D6xjBEHdbtif
9tvm+Udr9JjhWneXugLnBDF/+ieDHUrxKW0uoszzOdMip8LwHkk2V0jAAeY98bYX
9nxjJYiGG5nq/g7+tUIgL1Egd7LPIeJ+dAJaS+WDBqFzZBtr4Yhj6Lx60vzjGUrO
LkGZcbEFmsY4SUvbdO2/jQ==

`pragma protect end_protected
