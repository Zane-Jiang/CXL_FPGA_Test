`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
mIr2aIxl1r9dZPpTZ9x8u3J/Pgun+0h4EfUUp2x1NK22+0zbiDf2Mwyqpqn5ItPv
f3vg0lYmBf4avfY+hRX5ROODQkMYO9w3DeIFUv7c0h3R1p1FMzAmw7duAtlZX5kU
AhpvlCZu9sqQHtX4wpBPS9mKxf4DrAoTuWYVmyUNw1Q=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 81536), data_block
4x+GS9o2ks0xQZ44MY4djc2NkP5+2Vm9bLpEkVenZYaEEZBjvUvlDqAU7G43ezVj
+eDQp1BzpoPS+ipYxxBl7nWAuCLohrD8AjFxgwbocxtwIbDWvDOu6oJciO0Y8fI1
NGiepLnxo/1wmYCS9MNho9kU2hVbEN3viPCYf0EhwdRc9dzvXSgWkB5VEPFKRU8y
18T53M90Y1gBCR1H7oNGhj2yCa9vC89U8b4r2LrMAPW7HfSzK9QXrIF9aDKbkijW
MGkYDVeTzNYFViOoNM6PAulSkRVk1dEkOAKt1fZE0RjKp3PmXnIsH2ATU2ERhvYK
D/kXBYXjqUBBgrmIXNyBgQH0aZOL+W3xPoiBuoRIuxc7Fiwaat02rDxSv0DjSQK8
zlxdLy2V2krA8pTwuwG3dG8Cpxx8uO5Uf7fxYX34bxwXHZ4xgLEzA5RnqIGLHpO9
5a7La58nr3oUDEiz+LO8IMCfO+Thdk1pBSyL+Tz2Jh82yLUWZtG4946ZohMDxnmv
D8O6msFCcu6CwR701TInU3lDZvlP4++qyxTEO1GNwx143/ck+hczEY5c44HcCJOg
g9Oa4HwUu9d+qmf8VOnWL8MJx/P32xOiwXgngEwuuflz28Fxd4Gdo82uGyO2Ia9B
Ygis87Y4k2ly1+qMWEqhHUftOZOWf0mr0mEZRY2CqVTN3C9DLBIms4IGmateJIa3
gDwJG5b5ycQjGJhI24QYF6lwnO29Dde54ir4FQPm/tNRA6Awyg88KezbKY1NjysW
/zvOGv6c9Do6XocVdzEi6OHsBfojo4z/q7h2S2Pl4Ia/4vRmmtiWXuO3wwBkOdFL
VVFsyQHDXqC2m6UWPlM0yjHubb6rA773UvgMttUOfa2QFKp1Nv4PwZaCZIeVmbs5
cUR48iwrks++nc17fJiYWvUsuOcl5i5mXk/3Bv9H4Hpj6CHrDoth1HU98gY88SAz
zn91cqSwmcr0xjtSEAu9oeCXGPq9UuigphSO1tO5/9z5emiDKqIQ8WDGPSkYGV3p
gPrNWgfvP/sNZCBo66eQ37CQHVtJ53Pr5IQITmr2kOzn1sTVNKNb0ifr5xMjCsYF
vFDJvBbzJLcrbB4PlWbfEAD22AmMTpB4aRdlkuiajdHMH/qiKXCJSMDPnrn9VOfc
gyQHwxnubfjSnWLUH0sllwEkFQ/guoih8YR5f3LilHbQM/ucFSK6e/2fpNSRhlwT
ysCvXCq8GqYq2auXJF1+TSkVCktyNfm3lhLxmjZ6ETG6psmwDVBlbxnHwYgoOOun
xWIqWfbbS0nkbCKLVdGoK/Hw6DHX2DZkp215dn4U+8oVRSjj9M803yA1FhII69JL
T1l1ChNhBxgPXTpSblOoxh/wpTVGjh+lOPsDnM/yuTg8k3Ag19qQ4puljmM+gwpl
4I7aPj4jRqvb5Xfm95+YcbSFhJWDdVN0BbrC3wzoVjVpbUbPB+33HEcO+sjtVvNk
FZVR5ApKFR3DL/QE/4UMI6njrGB3gnlbJjZx4myiHi3/FepZAEcljFcRVDs4OZ/D
hCXFMZ0Ha0U1kUPnLO//SxxwxmT1luWfI62T0yfa8bBcSPJ5l1CUb/zTFFB7bIMQ
J5e/KUO6w24QjRtisCOa6vbOwuJ1fvY9T3GZlNwTuCA+BxUurWpmAatNHyrJ8K3S
T/N3ImM8x5WksYUHYJHA51h7p18z+SAvW0kyG0235V3O/eFNnsToNybQIne+kavW
kE1qEHail8TOHjU5MYNbYWHG9acypHLQsXrGhdn5Mo3xDZ0xKVfBNJw3meT3Urxx
avcfNNskWsky5wlKD3RolAwej2tE0jVfjTLDZKr+xYHoKfgOpkHwf7DeVszGjYun
2vmcih8rSrrd3jcCpmjqehTDWkL6da7dDa1A5+NlL/BoH6PjcYJ8R8+q4PujuM0H
Ay3GNmziYOcAnCZ+KnG78pUWUDXTo+ioSxCvdJ2ymhoxehXCT9FqLXnedrbHHdhH
Fn7YlNaYG8O7EEeq9JhgzLQDAFvWXiLYaYSGpxpHVRawcNKE5Yjde9F35IhZmaVH
0rA8nN2QJxd7jw8Tsjh0eVGFwYNOjcKHp3E+lRg0OK3t25IEaMnWGT5kYKVYJmIZ
sM1v8MPU8vHBkC5g9kYIQTGANkuY2aGrb0vAxKRGntMnEkDnvodU04ZKwvNZcGVJ
1NbbLX9Gw+uk0yULBwfDmV++1Z2qD+IN2/4G6Yr5tf9x+67r6Ji/pe9f56ye/Wj9
8uKWmMPVge3UT7SF19aqRWB50w9XJZhGajzCQDpU564JFQFgKl0kTD0QuDZDEqnD
dBGMWSzY+JN5Bf7GUZaU1j1i36T7Tqq5oS4UOETh7H1s5jesZBaiuy0R9OB4u/On
4jLjwcOwetNTcqhVrRCBMyxPbwNvlC6fW6NqHuAHnNeJOm0rcYk+F/wfsfY2WyDl
1MGxZjBxilSDKr8dvk9AfaV3J9ccP4b8U+pEpsAfumDT+Fd1bgpoIGLHwr5eX2UG
+OVoIhN2TCpqqmezBMt0IuU/9RuVnpyhy/W1tiwXLB+C6+LsmKagckMBCr6qugas
vSU4cXsmVaeG2mGDZ/7BtCkF5fQPfUYQ5exeNCVTFA4o7tSWshLSn8xWidKM0WBD
OotiU8Wlln5Qsc3aoIEOHa1FltMd3CnbjVPZ2o7xinYewbkf08TKV94LUPbGzHfU
6jnwRYYnPt0hAykFeYcgyU0zn0nObdqHinKS2oUgLBvoiZttFT8i2s66K6N/L0zu
x90rdhKL5J3YEI3xQi8XV7R4+aFT4Tmce1Oh0rAWLYqrrbns+k27vljct0C/ggQv
wrn20A8IWMJQvJbQ1hO+esdAA5titTz76Hg4nQIsDqBs+CqTGkdocnBurwSQeU3b
XCuQvh6ZiJXurzWCIn0SpB00MWGEvsxYUfuvjCzRwkDKCTIStczOfL+38sOQNW9t
++mHXKsokFZjmXbzulmZMDlQSt1ncQSu6Fch905tKH+VyKx7S4JLaK+htQ5SfKrL
LDppPKufXcTxwkykahCVvm17Ncd6Dsq+gdg5vZxBdRJlt/HvYYbXa18M1Ztir7B8
8vusjTGUeyOTK5sasqa9SgEoxocfZIV0Ml6SrNM9Vpim/lbQREdrSHpfKBtiG5MI
/U3aQQLAs+mTuY++whrZUiFSFrL1x8H/RqK6bbX/cH+YmNcHblF+xbQpwTmzl1GZ
yE7fCeiyt5+4bkyoE/90pYwh76srgn95K4MHJCegT+lvz+xWxN4gVfYg2B/bvPfg
eKoCcQKJDyL8UR4fT4b7e3JJOqAPaZhbZhaus0sqvGTOYm+5n0E/wLLtPQefz0zq
7f9+raH33CcHg8Hb0La9yOc5BbTExHIwpN1sXCAxcebK4Gaf7BOQEUdeg9S1Fx5b
K9FJCKP+H+hS/1kNLHuljEwE2bg7tenx5gFP17DoekZIn8xJ3Fjj7Y2Gqp+GnfBF
aOefEbUWnjmbZsd691KTaOtUX4KwzaON4ixPRA8zZ41h7HSFg699dk6UWwz4ugf2
fLyvbgfm/U4Spawmmad/Wv/RAMtp2Rof9nQLSESJV90xVunepBtBO6KZyrEL3M7o
9CzLc2QA7zmBxi4FHS64hMV0uodKgdjmg91/ATF23jOv44LKziH31kXZBjnmLqHQ
Odv64Oc8IyEZgERTuo5UPmBUyktopPmziVTgwnEZzbJEd7ETyN4paInpw85avVS7
7kjW/220id5MGG/Zc1/2lEotkOrofK56Kv0QcjAwR0bdUUE/F+0+xMZ7ssn45UDv
4i8UJzivSkTu03PpkF4uK51xp3seWhUp83Qog1NAeM8Xya/f6uOgQNQ3JRcE20xK
1TuDna49dE5zAed0B/+F2/Gv3ypeqEiRECwZzIIx26uSSZvh4Y1LGDcDOTdTQj7r
y0fKaJxa+WiuF5FUc+f0iZPukAvQkCNarLGhKVQs+7UR17Q3E0uVPzM8H1Au+jnF
eUlqbJ9QSB4Z0G460BtV+Bya/FIxjWnAhq+dLKHkKpoRYsACg/Zn7J2yDVpoGOs1
oNyd+I41O4gK3geowMWPdbjVGNU3wMtr5NPoQ4NhFRx9OIMlC4/lKqNwUs2TwpfP
7E4vSnt+c82/H+pXGXD+Q1JG0IghQorjaO57o8IR4UsswUCmqE1pb0YnK2G1R5AT
tgx42Lq3rWYdAX1W0HM3zAmUVUgtB2Cdq2qki8eqDjU4nHNXN4X1aLYia38dkjGi
mRWqp7qj6xufVdzQRCzCEDjNppOFhQqlN6F4YqfBkC/AlZjVdKiGBFzv9VIgLPdG
3XMxzSBEKnCzDVm+wtkIZowf83sIBEKpddljk/fql99hTAmhq/UhT/JdmRt7Wt3k
LZCG0wyWxjcYvxuJFiGIng/XTfJJlgVF7Fnojk+5rR8Zg8fbhQgGFUusXt8W/FX9
Byt5jsNoZalIIUH27E1SLJkBYsXDACgMCrsdiwj5NAJ5JdyXham1UIei3LLNGQw/
Q7lsaorQT3OZXqiBG7CQC4AqV+sJwj4NrJUwH8LQq7pbHpUzLjoyYPUoQwUh5WdA
PDk+wr/IVWMRZu9RAxiTHKSw8YN8QKHsAo6+hWWxT4osi8slsx5cet/stm9xGWIL
iBSkol3rpjTjLq+jQwC2pVBvbLiItEgx07HddNFYO0ocs0ox6d12nmVcld1LTOjp
IXTpUYTsEI+KHytEG0ZpR9qkiku6FddpCQwUqwF8Vb09usIp6W4bjYvSU41vUea9
I03D4lzFX3EE5gGMdDfPA5gA38dX1gN5forgqA9cxxVJu2cuXgNretIj7j6yZyg4
0dCxQT1xwJMjcvegIA1JQfM2XsZYeFkB1ztFmYCAKe1W/Q0466yzCqsIZvms9UzG
PtQMg/EsUv6S5jLzHAlwa+4lGdmJ1Vhd06LEGYpjlrTxp6H/V+AN4nDBlw2qRpUb
IBHyRjqI3NNiyoUEk1f0nyWAzAY+wBJHUGx0Ts3FaGeu6Ui6Q+uHinvLF6Ert40o
WtSDVVOfoWbK9zoLLsMtQFYXzgizsjwlXx86cZBEh96cTe5Chis5PBBraMHZpH45
KUsLjIXhF8nGHA3n01uRG3WOGQdZ2bRPYmnENu0w7/SPdxh9D3gyDtQrUDqh+k/s
3GiJG9F0U6/XZ986fVhNy3dFmjzwJWL3oDgLBe2m/nt3dW1p5wZxy+RReMTaoCsV
OKi2a/nnlwErJ1HodSH/qSPWuZUdA3EOvtHkeu1F1Ca02/pmW8GcsWlMvUnA25qz
PLrnSO3NGSjqj2YZG+hn/7sJjsYb1KLTLcF+xEwW2F5HdD/Mi8d0z2SNZJRM2rbS
mrYW3FIG/mJic/pl7weqHWQqinVGotZpQQkn2LqrSaeFTTraq3fFJkHiSGt/UN4O
Iha6ACITR2MmgoWkQSlfbL8c0w5HqqajdBBPXk+0rI2ULKKJQuNBJq7H14qXH/0z
j0dbC1RZ5Rnwdr/pN94kK8gWYN6VBm6flT4xa4MbMjdKM2Z1JBiLHbU3/kCNVuk6
3IbOcq9vlsYSAesUVmFTLhVls8YCDX0+Gq/KcXW7gP17X+VWRtGfDX8+BTtdc8V8
viy657mNjEbBRJfqUly7ZxqJgw8xaNrIOtiJtTCQD5eH1k+xW/DMZmVWYC3IsfEa
CEMrfhQl+ZQsF/Isa+Ppq8QCMeg4NXkyf4q77mMCDpF79Zo8oTN8Cb/pUa5MKSy/
wOxuRYmie7/rjnEqzbCJ7qKSBgN9WprSDcgKQEjRNFanI03e3fQc6uh3+Cc48mPR
wrqaX6911NFxM/mcLd2ZTKaLwHoEfPgqjvOvKD3uJ7fz0ZlX1xR8bSnsICPTA/fL
FX7mO4AbpX99l/dTziJ5/IyxDdWd0fETLmMLN1q0Aj0Im9jlE5b6bXQKsvuXHn3l
TUVKrT2Zug656RLa3Q9ifP1WSfqEKGfSwlhD+GXJ4hLqPWH7mSI2log1Ycqh40bD
SFXUZ64wixjNIeuF3FN+9WpZK/tEKf34305w1lmex9kp5Y3IH1jIoz3nTO6VTCHh
mSLZYqWNp/z72va79BrwMPXQ751rOksoMsqCJ4ePdC9xvaNMCKtV1sWdN1lfREkv
237ki9wU584OSPpEFsS7sIAiTq1Fut8Sx0yW6jFEYqObj2GxmW/MfQ4JqrA2kCMo
Un09VNZDCIAQ1LNbFcBTbnDSS8IpibeOHT3+x/vyOLOeQ059Z1CH70Nbv3/Hcm5G
/HNsUaDUrFMKKD7Y9QaXWUQRhYzjsVptnj0fV6MKq+md2xT/6d/XO52O8snjLEFE
dYe1c9kWhi2oAhfAqNjJlBeQXQFK1vfcCT0/5RvdvkXqtf8EI3XrWMQ2Up5s/kXh
5gdsqttoue6cm7crYTz6QgZ0BiTPQrjsRNKqKI+vKXYBqOY18HfPTSRLpMH352+U
3o9R6oLh0k31G3fO/57YlHLmw/TZC7PZcwb2+UA2n6cxZahEgh7veEBCkhHxG4mO
UMA5M/s4XQnlGqrvlKLYlYpnHgfGciopYjEbDRj3No/nsfpHQ74Vzmv8v4XIEt8t
utXqZIdyY9AoV8/UsJVy52QZlhZT2ayllec1me2ZSmIr620xmL5pITff2Obo9MM9
H8N5m5uXjTQfZkxu7MEOGc+OzPo7wypswm6UEI6g8u+ayiC9wpMnKI9yV7kCu3NY
eUDz0rfGt9aUTbwnmCZt/NmdhIKB3KFCvOH8n8mnNLJkhCWDlvPFKt3Z5HeQN0Ga
idFnPX1SPYec9VClhupzlEpfFOUiEPdha/GFhL+RSyNwCV/5nuGKvS741FrkcGDj
ttSLmqsfVu0bj1qfsTo4skan+kVNEV9xHITY/O1th51zrpZEPRyIRr+OxEZ90UQr
Nn61UfPXaqkrEzsMQUTq1UYsEaFA5cSU70WlH8+QfsgB22XhtbmV6Lo5ZP5nWGqJ
hasqKaXj0byv4PS3rJWyWgnNNbNArW1DtAq0gDHIpDMEqjvzxUmnqfcO+0n5ehlh
cI0i5lsfg9z+rx1mFudWBVYq9zWtmsI95fg34SlvnpmubZE5ofH27NxPpBh/dm1o
AtjmS/Ivwz8c3Fj/avBzUoCRppPEbZcBCBFahyzq/hJ8PTQZPlHFvtQF2Z841JdI
c+foVv3EieELlWjHsbX57+nFcGm8jMVJ9Yt63b2rKWqBqzLcgL9Z8jgeWXACw9o9
HGKLlph9p6kcll7B/GXloe7zozbfzkSIwwybL9KGDZINkXlSEB3hiONpoX89/5N1
tGm7aXm5XWTzCzjD85GcSCcI6DKJgY2LoTId2XS6ESwHwjo4lII4M4mmDBxctPts
yNbVYqSA8gFJzgf9mBLP5g8rEjf+v7EAsOkcxHvidraaEopdCQhqeVe6uAffOMUr
ogkHr+c/3TD7ztlO30kP2M+Xpbnzmh0L0nU6UkjiyF9riQkw7U10lKrN8dT/vfwX
5AR6BhwNo56TeqFZllyfxYitm5k65lbfwF9IjsIRFTzH7JqQi0kB/rv6l7MiiwIU
bf6QOPIXL23CByATSK8S9dwtZ7hs9pINN16WfA2jd0Ec/YKP080GlQZ+PpPGWFtP
NUImaNYPS16nfN04ORewkxwSiOY03xVbQ2uxmlw4jExuR6hbNoclUqBukpgG5prJ
2+R4K8djTevTY3TUaIANuTM8dC3UkkR3D4hblaQGFPB7Gwuccdpijzj+1ZjoVObF
wuAkv+JHxyh161ylDlLHhevE5ePpm3YrOk0lk9KH7kI/YxJuDvx32VoHEqrKTuPc
CLFJLQePvM1Tv673TkOAWKUUxd+ycXMRQ3IUCz2uT8F9Fh2eP3D6QMoCOMV+hsq1
0SUDpwYkEERGy58AUXg/UUw9cJ4ALLFZlOhPlmu9DzbKun6PAco5awDgTpDXf/cP
lD0wklAw1u1owk2xL3kimVIFb+vQ0AcqK+z5g2BUVzwcMOvErNVLZyrEdzEvWmhU
MSiZpM7Ns7C89N6ySi8li5qDpOSuosU4cDFy3aFlhWl7k5d/I91xlJs9kXbSDgy8
PraEyAKQoFg6XZnvxMi9sVH1cRMEG2ktkX4MishhgnGALWAnDSFeJOo/erhuOj7b
K4oaWVM4mQ6+7rPKSmgXhq+iCkebGMxaZmxrtRe2leuPnOOIcM+7R+3xjDF46wQ/
x0W3qYQYKI/OuulvUNhVSXbUzzUJGlG6GbYdCHa1NQejF0WIQvbMI5FZcSxTlZk6
kKFmQEybwoBfAEWhT+oKH15ANVyIz43l0jAOfjPcGpP/TaBVVWxe36xpCoDMQyuO
1wj/bdo/CELWsc7fO10ZWxp/hl7DdDFNn11kndgAPaSIcDXaB2N/0otyTzGUSL4y
i4eLSjbHpBIGY2uthNJL1hbvPmkaJNLXI3yDqsR4kseEvKvacA9xwzJmnFlEb/ik
k1K8yocEKO3PM/wJsYS/RIlwfWR55VWFDI7JDnsJWSfmy6Oz7A3PMMqzpn1NhomJ
D2z23av3330kxsPS5EEC84ZaRy9aYWAyf6+q5iOqVc0Nw/kF765uLZCW7xzsAA2v
UfjDUbupLAtkhGPgUqLNbupgIUPpllJKCTKtC+EEVYrQEWJ6xFHo+yuLVX2FQ4RY
YaNbfv+r88r2gec9WLCeNWRv9RG1yI4Xpz9GRRYnVjQLu8CyHj1kQg+f5z3/9O+v
bSE9DjGiO4HDndFo58MXf50Bb3tf5sswbRz0Wg4oaoLmxs+124/t6d+wCDMmuS6G
172sm8UcjPNVKFdvvvjpc+P6VVzHJh3rcnw4jIMRw0irXEK/1JXDUpJtiaHu2Ctp
j7uPC7mraJgkkoHYkg+d3abvrBDiZXA8d9zHj5JgqQfYUxLS3/tyIT40mBvWqga4
1PjTRQYNRxGEW7mlxY/pIGmjDi0p19SIYbPYseY1ouL6YdqyVeV6GLn54PsuQjkI
iyc2es6MTMjAwDv+Q55nfSJjUvUiOP9nCLNhrV74JUZS1PA7xoR8nfstK6DNeyxu
CteljO4aiS7eBmyitBP4H4caBMeD2rFXS8TN9jcoA2yNZJepDM2BEmua1SGZIdlu
oraqOl588R+opinDahpovbbFkCiN30c0RLkJuWbx6cMmUiKsZZso7oSCKbkDSGiv
ZHDGPxxj8426bELsf1UK7IwZiYvBi5ERLIN38H8zXjn6jq1bl7Q9gF9V4Njo7PJ0
UgkRj4G7ax5JfxTu/kQIBn5FuL8wAgxSCz5dBQUPz6Me1ibPlX6z2fj9R1VL4IX5
1E561sLjYI1r+cfTnO5+d6Kc93uRejzfvbF/F1u5pES5K8EAcv0pnJEOcnPNOUyG
KQP3tUW9W0+IrUCGVw/I94KMUfc0A1DVwOvORf4Flg7J+0eemO5NpM3u1+IdG/kK
6KEMhqKV1b6uglCzdokifWofFCrTBdhty7U0dyle86BxqIRFeqv99UXyyvpnxaAv
UFt+D3QqFY4XGdtXPRvFWCkFEsE3IcxjACXXMXey0qaFQF3Xyd+VRkRoquvoB6jF
JZYxUyX6kgrqUpYdKAd8UowC8EBAXiJaBEpfFvc8BPVyISX3MHC4lMbRfi4NbTsh
cWl3orve54alHyU2PZKmeSCPrlZGZNp1lCaxXSkCMqM3kOPYOUjZJfw9j5PKSVQx
7SK6p5oVL4TNdXc4PJjQ5/U8cmav3dYp7PBgsm+l1n5bs/7+9QH4uKIm8BItVGhC
YKvH2J0l8g2a9OO1OiFB4s9jN0QEnL3SQwFjZQUcf2ovVB/oL+9qJv2M/iqg0cCF
vis1TtVBSCp/b3xK1Z9xbqcXAgXR76arZgwEG0JlNq9rICVyiJEoPRWas12WQdon
fqY4SpXwSemN9hbYA0x+NTAskB2JVo4QZJsy2NncduKQ9b8T8xNZk/SDnu8FeJIH
UVp6rYGT1+KoRBHbW/RwK26cnno5Ygz5rdN++HnDAfA3fIFBuO1lHzD4spnNw5uK
hCdK8V6ENsUiANMxLJeTJfH+Uvt76i5667PU93y7F7zuxelS8/2VefWOVkvzcDVY
KWAAaZTPlbV2vAfZBUn2ZjVqknG3CDMpfTHK8cfVK+B4JuKhTfzI+jdVBiojhTEY
/PDTk9fQlR49JNvi5h36Ahjm8+SkdWloXxc7lAixTckG8NGeA+MQNCAbKIfgYVOF
AiiKshC6VBx0Wz23/PxsSu35zPU6o9g+GuiAZaJF3v5GC2wK4VsS0xECl0QqKHQq
ou6E6zA3E7s1YiW6/z4iRINysdyW3v4Kh6LFfWET9B+SlYcNp7u1gS/oQItUiTxA
ogokVnCiKQSwleFTJo5wQdyH/VLGUuY+bl7ROGtmEpOwdnwlxJIHOSBHQ2uffJcI
Nhw7qe3e/BDKtVKp/agKHGu+59RN3CicHHzoNUSGWME3uUpMEg91Co0eF6uUbciw
xieW9BXgNa++qFZxakQKOeXfxQVN5d2KdtVE8trzDhID4d+uwuu428nvPqIn7QX9
EAYBnT30It0ESqsEQb9kHa++k8aWY3bGima1Yypu6TM4sJmBbGA9swuuFCwY525m
plolgH4b2wCXLisik2mrOQwbUptA5DaWGgpDW+gmBhASXH8sjSAvS37rjLebvmX5
KIM368wgfRbtX3/tzihAbC6j+34roOAwXcWkbwKC2co7H6Mq/ehvSqzINtDBWwOQ
CFEfN4yjE6pWtEtiZ/3sjZ1FOIBUZHtJQnKMKBFsAIyBnwfUdSfzxUqBmk64OUYl
5ShUCA5kWySskgjLsCnkggfH4ctEwhRCsiZco7s0fwBBn7c9ORnmI+z1358Gt+T0
L+igyrWDIiCn8XxAV2/JsNEIHbrP9Q4VCfWi41YHGUnXkhrH9q0wi5YYfsMZizzw
I5mPERiMy37BPjHCWlucYLvE8PD7X85Rl/uwyMEtadG6V+x/8CSzXwHgDk1B/ZFa
Rb2+GtriJRoHjfIq0DSUbZvetslFykpvexEPUMotVJMk2/HRrJSVbbkbEIdbjyvX
Ym0NX4TRtmK7VugcmQq7mD/1YEZoMvOKxvw7Vv01dMU/uFvknCWhqdrjG9X55b5u
8PiHiPNVzOq7E2vrQO8/o3ghm3aFN9X+SbIMKBAdNXTCLqB29+GVT6dXqgZ810M9
vO6H49xG3CYb2+NvOtUhDFvS5ipqsN93qaDaKLlX4v6/vopUwEeJtLJ6qbsDMJF9
lGZp1UXo7fCanhbsdbGXxcBFg1DVrLYZ08y/EzpBo/2Sq6wFwXyfZbekkUPKoWs8
Qu8b7KJQQ/TDmktFzz1gEcVopxe+BnYJKbSHZxqA4bF+c5DdT1MNFRv3YPX98eO2
l443ubO0I51zRdo9mSSuzt9kOVGjlkcJQ322hn6WqLkWoGjqo7sEJfaNm8ORzOiM
+rRNt++qQIseb+XRmf/245ZuT4X4Nhaardg4IQ77EwHTJoLwNUuKUwSh5CkvGWS6
eN4gMKv4vhHB+ZflibqFLQtlOQ75rBNY2F3oJpD60OWZqu2fbY4m2nHHA8D+kjm6
QNq/jBBlGE35ZiIlSon4pneW+n3JVsoIveIKSHVFYUpZs+BTcBb/C4MIIROYp1Z5
UoA0Esea/FL4XrhVYEiEhT4tdtkXuWwZK4m59cLw2wDxuf9vss4qx25+CYBbpcnx
ir5mdohqYHQv/TFKjtFNwNPEdhNWqu/SiuzBNEIfRW7LPMaakOM+r3oDPM73hi9+
J8iKZnw3jpGh9BdW+fDJgpLxKLlf2I0m+foBvFmRQj//jpBGDV2alxe8vxayjedR
JsyawWUtQTTPSPXmDwaMtsUk73BSY+17ytJ7iM0DnhfCI3xjdLF5JwtsFN4Xp1Lr
aHdsZvaxa91FFZtC1ooDq5oEpmXE2aGAo3rDUC0HM+UFTqKP5+1rKUYvjhxxtxh7
1UEHVWGVczNzJCp8P7WGoQMEPlaW45ajBD0bVNMFicdEDp5y5NvApvl6W6VW/ahu
i/jr26ewiED+++SCEOFwBF5tuacBIZa9MREUf85TKmsGlK7y+5QnVcSedNeUI3UI
Oh1rjr03nBJDfwslpTL+JYmrhwyRPhMjUySG0qXinHBIZDOcRF3hhZCbmCzIMWTk
ctFHq8JU8Ek5MHsZ2dhGfQ3F96ow1cDCOkfVIO7WtJS+vkTwn3ONkWTcnmE8Mdd9
yeBCnkHXbyVq/nZmItQi0Kj30qFsSOQeVw0JzoCW7rb/MfWBa3FghWx3Fz7QvplF
RHp40DJWu/UeB1w4MkhFiAUVylYIBlHbh/eN4np5RVS/d+c/PSjF2feDfg/9VWTf
+KkCg++sX7LU/NF7MbTo+vwCeWCf9L0ChhvURnTtOvIfNZIweaesg9YiAs2LTWFH
z8w4es/IaJSbYumXqcuvJiMVdMxab29M+oF7PCFfFBBj0MSfo5wXfCE+j7Wwl1db
QCIn3eizCplE+fdJiiyxVlRqJw6dk8DLCXsBXJK3Uvj5vbJLAjDtkZsDu10nD19A
D/eLsP4GpYGpcZxteQepg/QEsQp7bZRwzf/p7LGbViF6t6W6eyQUTPSRO4mvfNYF
SHjVHOfM18Zha7jXG/5ymwI0oo/zgbximRr9gcIedprKttU6OaVGWvqIbu6wGySJ
hDqgt4NnRBb3X40AUTXXzCpLKfdqPlxZ5wq2A+VGmfdteMNJQmpXlbu9LL/9/moz
aPDfwHdcOwhE5KMP5NC8VCVH3mcAYSV8j9JIBIqJktyrx87DYih4wSuS1qxLT/1+
ghSdVy2eT4lpoqELBrWORdaT/DykGm2zepctCUp69BNhuUIx523R7dBAuDloy8S7
6IO3i8qE1DNIRS5vxNe2pFfeG1w9SjwLtyBckpSSLBL2/UyQnYb0Dfr7XL8cu23E
rBx6IF0gITU/pSMMkRfvWDQwlHfBGqtGJfgOhhK5huPpuBfR4vuFptoqp+X3g/90
JPTzdTSv2FwQw0hQYUlICUs19u2GQRjjlI/9jxBza+N9HdKT4GJse6r5dRpE0APj
En7nXBC/FToMMBf+2d3Vog14s+m+iL/ZekmLKoPhhq42sd0civ4VYsPWen/UZN1N
y3f0MTyjI5B/N9Kxtk7PfNslKmvnopsGqouG1XxTlCmKkJpE4ILe0IEzGh76LHl+
FtX4MDEoOQnAjodtcUCT4FxR7GgjZsP+nfzJZzHGWOe/AmrdG/vlgTYkO4Y4sdvu
zi+4x9095zxzvQ/oHRhLVfDPKiEhv9tbwgaNn/syAq+pyfF9Ndn+EmqaGMwqsIQP
vxi3qH68nx5TZZXKV5btTyo1FRB/4wAleHZY2ypxtRI06VxblEblTjvzAg4b32iX
AVJ+PONNFjICB82Lc4cL05beJEVowkDtUqg3kQVT8tB6gYM926QxzXj2khR78Syz
2YdK2AW6pGLlLny5X+VeBMP8/FgOlOlWjuSOWV2ANxm7F86Cyh1/BtRGV2mOnS+F
jPCyvQnCHqIXBCz7xbnJm1qw5GYfcwjEuOp09UxOWXbyUWi3HzQ1mHv6Z2NJmkw0
SEm4Kpv/OlmmAXGrXkjnA7bej4i/Rbpll+pqru8KiTEsJ9Z6E7FBkFq4l9O4bghZ
2KQH6Vr7Zhx6iwP75s3Zlsq5bs6J9KTncYX/rytk6ac04WD24q39JXbXLM6YM2fZ
s9e/3/nzNwaBYqMxaCqY2qXQuuRMpXWukmgUg3C9KmBOkBV8hS/algtN7jejir6u
Jm1imVXP62WvFY9viKpG0yFuOjPOPUIRhygKSou/b9/NcDFVdpg/8BdSS/DX6SRv
VmjEeTOreLGZDsd4PfDoMueLrqh2j6cTunR6+I2IUziLDXexVgXem+e9+cb+/vfj
caKcpdhh9s/fD4LDWGMTFJ4mqlNEMy0k0UisF3vzDClcWWcPzwTACRqOmfb8SkcV
z+axDnnRCilCRuC5OmdVIuPAvmkeCrOMam/rxduXXCn0cTOFt5CLTmMsOoYoB3R1
GMwB+Yc9rjbv04botR+Gcgf02SOk4zn35/IMYiBqGHxDwZUFA5436UdTO1UUd4+c
+pNwIhjkU+eVQ9fpMpFqqiutr1W0teM8XOZe/znb+H3iYMBpScHtezZo4Hot51HE
kU2gUK1UxSuUV55dDkATQIiU8wQ+BxCmdtZnKgxCueEwXznXlzG5nXV3ksJFMOSW
zxEZnLZwGZeTh7Co0CWIkQomdjLm78jg8QHs4VY73A+iur9ZsK7B+lA2tTeXlrjA
ny/ke3M2Rp3tnKWx8gc3nOmhin/dkLhlQjVdEzgSYB796knGYCgXG2WatzCPM6JI
nhvRnva95utRDU9OScuKdMgMhiBYvFEDEvMYDt8OSqNdgRZzEDLd8NU+hMxvQcFw
cpSqL2iT+ruMZPoDj7RldyA3tkRIFmmys5V24q6YctDW75CYaqs8OOQaHhGmfYe2
zAFzNbELUJNxUM9wje3z+jiB2kZwO2FTbDpQf9K9blL580Mhe4KMmv+4YFaICyUg
8HTusqdbI1c/gvuvIyS4eaZ32X9hZobUpNRK83XnwJfK4kgGprOME76Ti5mc8+FH
k6dhEutJht0+KyWN/PwU8OLqMgTLmg4IXhvcOBDx2mMrsNBrLO8TqGjXlum+CIfu
8s8sDEFtpmp1iHORBaPYUc6H1hKvUFzoblh6U4PCLx/Ky3NSbj3ye551tBINCPgG
XyXi348q6Wh8wAOGSUDr5tgnwKNdr+cSxdLnka9MUrJPjV38PxPOI7AkehIkmZ2U
fH3o6kSEh9COuijlDXEBOL8IDaAx7avGeh+n4SdRIyfFhvoe5ofYPMbAgsLCxkX/
gEc2g6SO/Ahk1xkfWs2UGF+sIHt/SV19Gt7sTI1c31m5g0EMJyZzp0gHgGEpq3Ed
H9iC8Mch1uRx5OuszcvP4ZUrhI3joFa0G9DylVpo+BSAddiwiFd+LlH4ZJFgZG6P
NyLcTYN+y5KU8Jq0Qx6CtJHirsfxhdb/a4N5oFbffmH9dEG9iMlTERZZBUy7yOam
1hDULPW6NF6KzKZ8uuBa+oI0Zp4BA9wBd4IG1bcNpxJ1fIPevLVXgJDMG74mJIe6
zUQDRZfviQ0Bsdrbwa+n72UrSgdMP4iv0C7qZpeFXykB8ufXCykJ2GEAJjuY4/kR
h90TvkUV11ClASA411tY5G+FRWCgiwv5zLmdnhetTMLCog8V30crbXS96+Mh5sWD
z+Cu/jLBj1TYaweYhnVCX6w+fXHyKv/ai5QKXX5dTH1OejBCRqBdmJUj0m6vn0WC
3QyKdGT+3fU9yGzceeQaY4upIzzM1S2mMFYYk+qd53neW6PV60dY3zkjb0pKM1xV
JA/r07Zn9fistUg6d3J7nUMep0ODPeMCNnmqTKXZjEOEXBkIeqKgbgbp8tnWYQxB
4v1dtXL4XAkc/5x8WStEl2AqhYQv2PnSn40mBrdmShYM9rvOTCClWAzAQa8Y1ImC
+dSAom9/iIXErB+3EQE3y8U4T/SmlXsK0pAPLdY00FZdchgoo6507p19Rgc8SxiR
HlVDanVVbYF+i4Ed1BbYsrixeTFeKPaT+EwmXOKBn0Nrn0c8ySHFXvF6QiEyqyO1
IjJwFziV/KRVNynJojlCh4cmH3wxW1/8UtDMCif3UWcVErYSaZfw4z3Hwt3kbZFj
Qo6yIlPyA0ecAfbltSUqM0NIjrcXB81P5HzzVpD2pOYH3UtCbLAqnJC7OYeVFd9+
LXKD5/Ymwa/TbmKk9mQQ1zMHQw5qJWQi+Pd0kSLVzHqbemjzESvyk7LUdfc/eBJY
xRuuF4KPeyQi3ofvwPY2xTR4V+xxftMBFbVCAswbUfPWXz1sN2T6t7PSGDD+S2ni
a8LsheUaPrcZOADwVgO6pp2Oh2ng/7MeepAeL40IQCcUR9Y9M72guBiXZ8kLn9MX
aDckKwHapnCl7f3nwBqdZsiIL9t1IRh7AC6le7rEaqm0Yz3WmXikaKBCB2BcfM+W
zoNl4aWn0TlD6GkZm96v+X+SiGLxmxIXUmLolvhzAlRkGzEsx5CyR7q/DSf2gxb/
zKm7F3Z1AWNwVnVCdJjNMBbn7vcl0eQfy0um9gvh6qQt4c1DBHBBhWVpUT827n7y
5s8Z5EJXMefdmExTpzsxv3NUTgEDj0WYgt87UehKUdNfv7p3BZxNOcXViO3Nl5cU
W790/lxF0I6s1A9wCZ7ko3f0eO4Pod9nsFEJU1V/wROGlDhv6fB5U8maJuGDdbpM
tcMwnT1DDWeYkkgfeXFFtFSJjjjJ2SVjOVXNASgvDXDCZO4qT9zC6E2Znko0Wzg4
FmdOrAPcCEfVzMrRhDNQYCiMwEr0C1Wc7XzMaIgAzw1Bkbc/Z1i/VK0tyyjpF8Lx
64/LZ1jvO4/mdT8w6sglSj54DIAj/6ducch/JEMUoGBxiyMtBWRaHkDUq4KagOYu
sr95wE/z7U8qWfnPHN9hblvFPXVTlWcg4YaG8gDybpjBr6Rend5j/7AT7gSz1hAo
Frxx7N6R77u269JnTUfbJLgxOm/YBof/8qcW4jn2qqwBnL5QlSBoaN2V41UOofPE
AdtsqcNN1k7QIbhgcaH0y3EE5D2DA7lZDoyuMty4spgAxpS0lzM9LuAlCLjVggEM
YA+1WIewNvnKpM8XW7awjQV3GCfQMbNnE8WJG1rzhW0WbiEPSchrY8pQybFQgP6c
oIg9WQZXALRWRMPsLYCAflQdOB3mYBXu3IFwdzFhvUaldy1xFuUIechQ9smqCw9t
oyp9HqGvCoMQQ0onRmY8NIjgi24vvwg3dm0DXYsmnZbDdCddDhJsB8WPMaelQoJo
Xzej3Iz4DRZ7kyeNR7casED0BZpq4yapmkC7Q/bPgXKpsiP2D7uf2A50p0KRtJHS
p1XjQ0Vx5vkl5LpuNgkXA+4uc7nf90fBpiEqEu3FbDzKkJ7tcT/jJqOmt5Y2Km9k
L8JsnKyUjueNNNRxhVtnBa8Hg9xRXtetT4BtvHi5MaGHCSkVnwE0D87eFMk3dkJp
tV+dPuWxseNXw1289NznrUuGIEll0QD9oBBc4gqRPwVLFBzW0mhoskwZjVgha+ay
7uHbYL9y7drk2dKP4bPLVv5e+afM2W8TyR3SGxKN5A+DDi/x0NAGs3jrc56K0bBV
yXH043vOOAFHZwa1WrAhQ95HEyV/q+BnSLsSpMUR4p0uhkdvZdU5fCFtsortVKQ2
02ebI98oP2nJeCsTLS6avycvr1+BRJgsPhwwMtbIqGHt2jttw+sH8KLq/nxxTOcz
V2/+AJtbmQ9Dtmi9zrqd2QyM9qzKChgLBbKkbhRr3TGiUsgEpguqEiupASXzPbwH
vxeIvEFNC2MgF1ohP4SrRpKJGXpaqkWWHa9zlCTeJSetgCeO/1jXcYdrbm2DJ8xe
i4ajXS5maxTIIbCQ8EKKIiRgiNsyrJp8hOIRaIdUhgFMjNImuNhO29gdpzVhKryJ
RuDfNpX2rATi6ijQvdhlXidDlVRVdULjzQMp8rAeWeZ+FBWl8UkTD7bac9IVQPDT
huYcIGInwL5uguTGUuCg4qlCQltP3V6B8aVA8brSGePp+F66GVawv58sKPV1wMb4
eL7+BmzlovyDhXxPmggfdygT1kXdCQ1GDH9WNbnqGYx0dFvAms3+2NLwsbn07ZUz
94GVYy8dMNcsFF/gRXcO+8q8ffTcHN+OS7bGaZx739wIrI4tfT/pqjRAEz3rDbcw
OMEHYuuWGQZBvK29B/gJo26OmTMZ3SgRul4XCvjIq2AV/Ovp8WHcXI9GeMHycItI
0+bsT+dlzn3jM91RG7WOBB7V3TzQGrX+KaSRhXLVVpxWdY5a8ysYrNQaHVGjPlZ8
EUC58Mja5RzXT86tfrwFMwoB5vJO/Pp2GQlh+moeKqrhwIOMgsNmSAmalcoQXBJz
Rlhxpi7Q7KyBinlHWi5/QQCCRqulgWs3R+7PnX3Szvw84zkSvuKWaa5nHFs6S0UR
X/Hc2vvt0K6/WfvzbCb8nc2tfq8eKuO9up7VC1N2BNhCIE9k4EtIh7CCa6dBHMQQ
EhJE6VxJ9sF9GYvrlmW3VwALdCTDVrWJNz4hJT2qIIYatlyS9QH8/q+Bkg7IhSPe
RQjQioo0ddC+E188hlAF3VSL3aOP2F3OQ9jARZSwnZFap+IGLXgOhqsnbG5CGpOL
86fyyjd3rI+Kxbprvq6VsQ6fkX9c4Bn6QDl9bRFYSNi9/zRbgzTBhDScbJZmSgPa
/MiT5KoOvemCOPV3MVU3ZCKvkpo33qqnTvNCoHOxUAGmXgfM6UG0FyQLveNC4MJD
sscSuKoJzCZxqGqlY0+pJwAbJYK4LEY1TqnonvsYJ3tvv3ZnX293lycUhW61HLYS
BOV+RR16lOmcsQuxrSGTioqZMnR2oCoXmln/GoUbPGggOdjZxibbwqMedgmTmXew
JNOeZPWZdWN61JYSq6CtxylH/jQzlvKx6OGLHEhhxe1/AsQSbD5fXfDcJfqFihAs
sUt2GmuiTE5wRaGzKx5+CNa4Tv/kAvKXvxnfvJi9uVT09IHqteD4RZEFeUTSJMNO
NbCiB4V6jugvmC+E4AqLIDhUeOV7w1908D7ceCQoPx/1eTr/IWKs75yJNBCWthP0
9YstdFSRz6AFboDvSjtbr3xvZSbvgvcfCUF8HXXB4Ez+BVbGjELFvIcYFvfdQxnp
6VE5yKDMRt7TIYAAV3vzp/sHsUQgDES5raQLBtv0vzi7wzHgsiP0MYF/JzCZV/q/
JhTnUPR698m1knLiv7wwrW2lWv/8WBlaB0EvZgBV9YfuMhQub4hC9am84YJdp1rb
Ic9TrTcQYjtRtTy4kh5y5papt/1un+1tttpBkOqrgDHoLfSC5GDWYvBDuE0vX3Db
mW5qsaQWNobQGMhnr5LDk7ptNLGE4KFZWWh4Lr1C2wmDtLFuwE/iAXOdU+aT3D2K
QMdIQxY8U5ZGNWrXlRHcC+uIbzOnSwm1Ei5VUGMcd08vj9KsPInu0h4JhhK93oop
fY2CjwvoFZymEvMHbF/S8cvgGsECWEYo3WbyLEA9EKQPiQT6Qa+v2mvQA6wgmlmo
V1xHbPxmAS6ySaaj3DF4zu/UnJSHaEWMU4q4VuL5uCfEWKS6Gu4gGAEXDucIJDEy
XF/WdfPmCIM/4hD5k+6VxUGh5AksH2oKq0j3+DLcEtNai/lpFLBGYhr3iXoPyBGP
GqAqu+mTs0JCsi+U62kTc36aXfTI06EGGUHxA3bmLDfVs+RNsp+VnWZydbHHdJLd
ggQHmPv0oUBwpFfNqc278fpS/oksdxMfkkooZ9kGgs3KvHw4S0ksakcDj/Utez8I
TcsbgfKuKjMXuQjd0Lf6UIKu36d5WnErZtDuuupUcdgeDDktvv6NndD2xKpSPsNK
aQWS2qaJsbsUyuqYdENdrDEKaH/R+usZW3InGSE6BODWazSVh4v9BQofGrulzIHb
aTTWWoMQvZ3tDzxufucq+PQwjwSR7X9Hnm1bMRp0tL2dq0EglTHHzAhaxGI2vlWi
8pbMmemmv6f1qQlKvSQYQEH1soMReKXDDPbF2VE/at8ZPoLfb0LwQGj2PMZa51lU
NC3rovMsWKheMbphYciBIX0d9wOTb2m3r9y9NKe5NDuy+VWodJHPGC8a8NQScnti
Sb/HndGbazGQPFk2vhFHBQAWNWGOF1y/QjoQQkms2ymJMiJ1cgu87HuReu6U1CKA
dZA+9qXdKu3exZFbpYUuXkyrt97DJnUZyBY33heQveQKD/XauumruvNbe7AvZ5aq
KidVVZRNTGZdGM/EFxzfP+5WGRrp0L42bB7kuMPuhy7fEmxtcIaPh/eveKDNCScU
6S4ZQUAHGQCWB0s4MTLEFJzSvxCjhNBZWVQH8CgOsH5fadrQ2fmL+9AeajNeLXTt
fIwMr3EA5dJ3fQTH00Pnm9dtgIJHqtmn+A0cAk97qwHcNffv6jbti/f6TXw8BOEs
vrP+oHQjWWuo1MMPFn0UUd8A7kAfLgYyzstC7Lf/B3OPDnbVZOoLmwdW0p6XEIgy
1jQ29BWCgk+IXHpXxQHp/qcC8owU4kEn7Vt2/ut21/3UZoOmyyo3MYwu/ixQktNo
6CM1OVcrnwB6P2gKZvAJfppH0U8UXfNAD4Of841aVSzPi98A62RzzHjn7xDFPN8D
ZfIxdP+81WxUmyFSE2XL/34cWA0ZwYbkDdgD7VtcVHV53tTY4ZK3J1kR5LueKyYW
jkKfto/3+TOk2VOYG+WwA0desqZXjAtrPA0zwTIDQg14YLEhrlW+8X6aFIosCDuO
adKvG+h4hh4IajhVRMcCfZxh2VNBy3aqbWc/gGdWd0UrLcjjl6LaaesglcmYgYq8
4B8dsI9JSObFIJE0artz4DnQIjB7JLiwWvjaigzNk1v7Cf87PGSIZbrqjz7joSvM
1c7fvOGOJtIDhgaV6Mev79fumP3PezR3Z6x/0uBzGWUsZ8pP5CU7l2GpQ/fYTdA3
NeDZIznKw1b/b7dlMyTakVMhA59+rf8rdjafEEmljtGCgc73pIMb6HaRcWEl2PaU
IcTLbes7VKzWTt6tCN0JmAOHOKNYj2VPanJq6bR/+1Aj1t/UCHGiLQZ+Kh5//KNT
BaL4/GXa8oMEXLAiVMHn0j8Y4j7wXudLkS6TbDhNKFgFggXxvi0OPehksEWCJDhw
eXK00IJx9c963IdYQI43i+MhzSwT7llDU4Nn0K+OH2KYmIDZlG0ihyvr6+BHBKCd
sVsDevmKWGZpufMptlHJEyb8moNH+fbWYwM6rNv0J/LlkN3kapyEahh7IRi4+TyW
yUuKChNPFPbN6BnUF1KdJegoSL03huDDQWle12RZKxwbPw2dmMMZXfjY3xvNQr+b
k/1DoHJ1dv3j3asdzTEFbcOkUi/4pe/KyeIFChSe5PWjQCnmo+LGWW7+UNZuVGJe
7rGjKx8iy93DVefj2Qn1D6tYp3Xc7sRweh3VecWbKnTpH+bwdVr6j9bKTe9x4og7
Iq1PHMFYJzL40yi0jt1718ZN2J6VYQaCplL78jf9TRGeTP3SgfOWmUd7YokBadp+
kbltDwmAg10V1WYvQlaK8YQtg48yqVkA6vD7K/XQToVcTY7BTEI8Tbn9ttPbIWzz
OVPURQll4KEaWRrnpX1+V6gDz4MzCeqakM/QbI3+G/MSTm48gTkI2e8cSMCsncs0
sQnKMqRlMw993wgIB5TxCOwgxCMSUH1dl8wvxGUVm7OfxiMKZud3HdXkikifTU4v
KAUlYvb4Gyh2T2dsdrv0PKm17il55QcgWYKj0HRxCuWn/7BghLQTTv6zKFNXXDzu
uAYOHLNiakWJ+5nixy69qhMqUDq/jeupwIqoC9MItFjzNEVNjlu0R5m85grH3tSp
tX5/FNFmYE1HK9CXdLOMDXPS4BDEqA+0GNZIXS2wdr6nVytdd1vRwtcfbFnmo+br
R3bM6qdCrcoFimja6MjAJkJxw7oJ5YaMLvVThMMVXz41pxuRc31sSpFKMvtaxpON
kw4NUUhf/ERmTi4D017vhpsDVQ4q/4vfizD6rLv1YGFzwLVfQKmbxRrmSmvHPPPY
dfOTl7Hn1SHOH89KbC8sAhtM8MesD8bEkSuqi3tcXH2JnEc/TVTvBWAxxdTFEtvB
7+/IkAX7xoflLaGZAbcLGFAx5oMi/nHKvjzglB8S2gTnsO0jKoYfH3V6TU5wspQg
oDD+Mdr/PjekjuGPYxm9OVeGlUNcIUKM9ZCA9cJAS2SwIQO9jjtpBMBfbHFdT4BM
rsRPFDgwtuOn9LZlaRl3ThIaabs84fCh5JehNiLzoDgSlGMzqgUnVWvrxIefrfpD
YFzpvziVCAuWee/3IQF24SAuH9iDVwEWRu9RxjY8jNJ14hb5nLuPgIMLysCpWsmI
+f/fiT2IMYNpUcINaa6uxcAE74uZitQbFjB0+YULYvRtV3DVZryC/LBWxXNB1nT0
y7aRnQ/OAE/N95mygd7a335CzVIHlwd4soCuQbNhlqJGfgG2+0ABTHb0j/E6dMnN
m8AcJQ3qnZlDaC4pYv3QCrtjzY4a4Q3jFNlEFu0GAKf4ZpSQty0QydW2EBaU4XWf
WeVx/RQiwSOWvWetRRiiuXMiAYWwZcJwwp6o0/JWNpxV+LWXtWdOuB9zIhQExcER
iyLhF4bLJwZpxb9TfE7hTNU0x4fCzljIHMVPC+yEycICLl0ylSlyd7nobTcBIUgs
BPsLMxclbacL5Qj8sa3kbY82Ml3adZh3WWbcJkultFycRpHGmimKtO0A1TSytksL
JyE36pqmQULYI5jx1brrO8flIniMg4peTIDl7UbbEFRpG+kxz4yqGlRWxtyd18kM
0je5zWdlaEcN1UT8eZCGfVrbY8mZ5WR5ySG11Q2TgaFKq/3Ha4LS4Ysr/g3r/rA+
eQMdXltkQI8DDEcE8LumCBSdi5e+CsyIKYom89YqvHb1I2+dd4fGGTneRa3aNeIO
5t9rPNQQw/ZSE1QkaC9EbhskmmBSOSPGNi8fBfkhvt/kq0qlgLzlRvLawDMSv1+8
88/J1Gq09zC5wUHvtzsprI3ql49YB8HxdA16Bc50CpsvVPBHBO2T5NQwK0l7O0aU
Qv2A6rfj3WBtL2ICHOuoxYhEk2CkMKHHm5hhuFGBTILQcXIt/Q433U96aykV5Ds6
b+fzi7gJI0ypx23aHMXbqqnZpAgNn7pmJaCqoX0UsMUc4JN0S4iaR5SCvRHZE9AH
RIQ1lLWs2ze1K2EzOrppaDigUu4S1B3aieTEo7OV0yAX0FtSEsdRn1dVFW5TLKg+
KZxLBVrpwbquIxPnpbWpf+m877SqRAm73j0Kc6D7js7vKH7hRxfHGPNBp6tGFczO
Ic+L+TF3zIgXyNsAV24p/OTUsA/cFYjzLosLQs1l4sqoWpgxuAf66SBnzGVEHzzr
ankbapU3b56rhzLIa3wVAkC5TI8JbVCnFP8AkISPa0Vy0MAe8OVZA9iPuRS2WHnp
VqQILjn5mR6sYa01VNf5Io4DJVsvOMMENOjkgg/q4cCXi1tho2hqlKoFFbmfuHa8
aJbQaeywT13fu+jkfmAm5RYNTCmsipnQftsI7hc56vgAX0bF0J3xs4BpWXVQvcrc
C1WqtMlShOzc6YzA2ivx0OKS4F4buVQZ+aaRBRueqRgU5yaazuFHPSdOoxCP22/r
K6UjbMBTXJy+xun+T1jDLKT3kODRimMkkF/GQoRRjCN+M33NYgV5a1D9lczUJiIF
Ox9DuccLWtAaXTwW4b4LLgewXVIiw5TFqL5MARsM3AaLVOt/d2D5qnkZvupFrYhy
cy56kncGEAoTrsEpqx0EceIlxWgcyYB9p9UER68j1Vip5r9ueI/UMmWPzq8w8SoV
a4O/3Zx4B/WYox+OlMmCzfAo/4/07XEKtiNv6RVgDL9CXl95j5ZeuYNwrXLidbx4
dQ1NuYTDiBEnUb7oJHiSWF0+mz99ncQgEMGdktMpz4+vS2v04RC1KPhLuN8duQM5
2U27lnJMc7qLnpD6GhySlc/zYk51rSK38MJi1tz5sFP6FzrgFbaIcSioSDFqfxvx
DLwH2uYPQMbFDkmZBIwX3ZlBBhIFqv+RczR0kkx6Kodk/beZ/9cLO919JbvwGiAv
vZqgynU+DB/9CHvMmMMXn4PkEb+sAY8so4eFmjP65Wg3K2vVq6hFDgLgglvZGf5I
Ds/7mZhvB7RlZbgF1ba1EFSXVPghCMQgeM3F4R8j1pQGgllzU93WhKVtjDvUrzXi
I2RE+6cgOo2HBGK7HRabBGO+h2xF79UHMnWwtnTHYpNcEtEkftn7kOU74WPMGAM5
awLZlSYKHsqEA4ireD4MWLN9jJ9+H6+VRgK7LHzJg458K8kW1FQPWH/flwhpHMY1
jXmPJiWfhdcaKDt+xPtoKmdNa211xpGHCrPunasxr+DqiQYWdUKlqjF5eqHCdw0I
bXGiUGqHytl53D/3LdMITGuvgMaXuXQcxY9yPnslp6VdNmc3n7F/lTGpDVxdcyqx
ipZgJiONvEc5m4dtduPE/tFnFwM4v/qOmcW3wQtyl2KffZxeQv/xTmcrL3tJjMlQ
0wFBhh3JzHYyFw0LKTCUkYwdEdCCcTSX7pPHogEsQvxC7eYlpAF/AkmOYjMc7vEh
JZdx0f8Awr2NH7GdoQUWP9XJyiSBwpQ05apgRu5jWdyQtytpuAXzlwP1h4dxnxfH
Fj52CkNmYbzTo/czY5MUk2f8Mh0CjoYWSU4zW+NstzqTZ69I48EEHgKJ1S04YySt
+AVy8M+i5TaYANkVsF0LlPxG2+psZwAiFFFEf2d/UIHDnxmydYLD9K4EdbTYpgEP
S9dpSjc76PMZyFNpZbr1zLmG/0PhSOlIBOnclaMeNvRrWRc3CyZ4Y2G/l12nUnvC
s8hrGzJtqM6sZyxcVJI5asbO65HHmn2PpQkMOxbNxKwy1MpWKoycNQjQD1qR2wlq
1OnlN6XOCA73G5NXRUAALDpFVUsuDvbtmJf29aORaaEKAFfZBgUpBlpWNAYgFua+
ppJx4q7vQJB4ePytYk0mIRU0FmJtgsiEswNxw1Tp3H6QNu1KCulB6+CzxoXU1HtI
HnIBqptin/8XnjExugfr+i89HMvGBqzyR94njdcfShhsrum1pgRlf5lrqUuJ+Sne
MmDg1+v/CAMx9+SE1ngKDENK3+Tb8+5WDIw68LNwt6SEqObWYrLznX9Z0ei1UgAG
HwyhjI2luNadHXOaGGCWQp5yhLW4fgD50uOhpSlsJS/KapX088E8oTVCtg4A0O1t
k3ZvKJGMzqrP+LxGZhXLMM/LrPI3vVO6CiZApRQ8w6XFqZvlWa94xvZFR2tYne96
Dob+aFllhYUJ/JhUSO3qzEtxc5E2oqdLNmyhJXhm4pvhb4Bei4ggGbA8hrhXrtAw
7OrQrFfxrNFWML7gbGq8SlAZj99t08BFF96j+MMbc+PnWt3/5yk/PBMRMwiosRxF
YqjVetYrwbxEKrdPIlzbDPmli5FK3ANiGaNuCtOlN70EOsPwCHJ7mYUW2DNfGkA/
35SKmx1XqwrcpkY44bnozDbU3tGMJLWpP2TvxceLIZ3IlQrLfYvxFOVz1kA5zT15
L/pLKWIVqiJVp8Eh3mUBlfsD6tLAwgdQSHECdCFnO8dXUek4QlSHnzcp1HQWBu+O
tbn8U7FcbvXveizMrGo1XlaqrgVTtXEc3zdQ0hIhQVJWRP0/MUJZL+A9suTPhDmN
xqYfJXaj2Cu3v3o/i21zZCkwW2ZrhUXw/p1Wmbsxb+6I+1nywjObEcqqi3pwmLfa
Axk9sQZ0Zid10Bb6dMhB+p1OutAurX1xnhT9khib+pECMxZ5V4z83pn+J+fmu2tg
QN73w27xHocg284dE3dtUSasiA1VCCAAXgfxMWPYNE0ZvjvXXO5Qj6+dfX5Cvl1b
7pl88wBycZUSuKaWzoQ/O5c4x3vMXCXjVB1Giw3Wu4Dqs43zAemoCD/632ue6D9j
CDl50V4KfGNhwE+nLqzWQHfBkVJFgiKIcpwfHiUtPxnLt90jWOul/79qGdstz6WP
xLVX4gNKGPPwnhewSoL6xhekV2/Yeo2Qh3i7X9LMFDd9MNEtSe+GgbYovYDvpxmn
R85h/eQT+vMXwUDyBxdqHwzdFd6F20KIwUw2njMUfD6Fb2Jrcjy+IH41EwR6HUQR
yFcPReZSuTMEE1FduP41U0520rS8nydY/7TqrvWnTtvCDMRNHsqRubPrCw4bGsoL
2+S/vBbV4OAm3BkOYAlkZYyKRAdLVVd4zXDlh+mp/QaL3XJYEoynjfDU5FBZm8p2
uiCpAYve8QcNkTz1fGEOSYMU/tqjDyR6AQ5LwLeFW7/e46/o6X5mKplUZ/h1zWm9
xJpJr+OESm7sW9IKj7Mag1ddpKf3nzouJnpqhAM3e0kvDPSheYc5iQ6LpsGpwfUo
vUV64DXqbnzHPra8jnCniRiIBatxYDjnpIJOihCxMeajZoAyZi/e03CgC+JKKQFr
8M6q2J9oUp8wC1CckWK+uXXmzyNOLZXGetIeAjjy5TFqpDO7K7STOhVv+vkZ0UJx
Ng04V/f8egfkmJbJ1ZON/DIbiFzeWxMlYww5nsOBc4wSC2gXsw44MYk8hAFrPGCT
dOEU9UjKSnRYniSgMQdns9160D9dXAERLLEq4S5Pw7k+eKzTXLGipjLV/gtUl3Zf
tOk+T42mOt3fPTiZ+Z6b98spyC79QTNJ2ZE4Soq8qqDdZ4APxQhaugeVC24zuIhq
GTmevZZbegqvCe44Hsh1pKZYtdpU1z6MuPAf4Su3FrksZLhL8ZcZELw+SfMK3cuk
GaTY7Hrq0srRqz85F98+EtdwT2xFs+Fi8apS3IJWTRD+2GWT8PEhFTIjC38b9/ps
JRNnxHRCOUfOPCQgjuqhyqERSZl+ZvjOzft8wkyZNVHTejDkSqcJTX9vYh1U3Ao0
yasL8RQp6uR+F86YV+b+FnIix7F6IWJiu5hB88392nDCv7/ZZT1D39Hh0SlyIev1
5KJS/dq9r7Rw3Ju2bd5jygsGx1fqyAffePP0S5QJU3jqrKRXxHXnLfa5yGkOBEJI
Q28Kt/ThnL4smMk0q9pOHzZpGSAkkyinnR5OhR+BBAwQEycEo9a3FitqkS9/EZqj
dOn0Z7l5XTpPa4x2L61gvkoY+cSU4UTVM0ZvXhj8+CxJ7RR++VZe/8+sMgml1gUn
tyMbcmI77pMdNkzKMiF321oIKKNJSw29nS0TvNKeF5110iSei7DX4Jg0nnJLkoYF
pXKNEhxVX8MoxYNtz3l6vhMULCJ9Ijjv6mTyz2LNcedg5halALKcci92FrhQn7oa
cWapzZ9aHfn1bzT19kbegyg9kXM14hFeJQnJV2zVFn82cF1JJS7tdIbe/Vwhu+2Z
pJAaXx1mScot7aeVU39835GOY9yfjW5M3CxRwTRG91BmvhHmTH6IJCEq4FOxxhCi
yCw6sEF75eN8KLNt8qpjeg65orFOIupQFBkIUgV3ZoI3MpfuY0w4OY+r3r/gGgoJ
Sb9sCU35lAUvc2ltB6uq/DkxlM31Q8wljD26HBIZL/nPA59oddqeozbYWYROO6gL
k/h/HkBm/ChBeGgjxi3SkZenjQE/E1kvkeobWx3hM2rihbYoQYBkCGb7MikRTfW/
kLW7VgiSD057CubiUNt3vrwb3H5y2l5K8CKE94PNgBqsRtUw15PiZ0S7jpxvZqlB
mmYru3WIOXS7qSsAttN5s+eTOl/LihsGibSGVONYv7baaVq8ByBYLUZXpEks+mUI
Sh0n9KHTsbw2tVe0Iit3J3pVF7rTsJnwAeGBJXxQO5XWLOWt7lA2rL7L17bF+6NZ
iM5fvDYuEm2yfh8fjZQr1kcZd5mFo8Pm/VXnW1AEOt5x421IWB+tGfCQPjP9uh5f
iGsJKnsQ25Ur0p4JDT7OZTCZpsacoE4JDo73/dJDwaTyzD1mDCYz28QFzU4po3KY
WQRzNXtsCqqyyEvJTHZKjo16AQp7ZVzQ00B13cLFCvEh+Gi+ObSEKtqwDjuniqLp
wPoAiheKatpnP51urIE4Mtp5nSHyExsI608onzeC0OMu3a7bM1NJDbVt/qNMlk+T
PVouMSbb6Ce4NgAgXDa7fBQPmrfHxIIUW6HFF/vmpgjUJunRxR/IFOTOfnEz/Wbi
fmqJVlIQOK1n3UdTI/3e86M8zwMng6nBph+XGz/cQXzG4WGcag0xX3BnK8iUOg74
AnVUN0K9DoQB80g4eDrBX3tzm8t5/9S1q3dLqC+z1D1TwTAYCyxtUNDdO7mCA7e2
LmkvJMWuTQvotpZ71j8sZiwzYQOMlOt9Ix+d6LUY/s65HNhfIpPOAarGIVStLHTQ
ZMh3B+oqot0tX1ba6wPFx88/14qnPO9kNBqRt785zr7LH1UPNFwfV9ft0x11P/ST
OOdYKZDN+mNXw3WgotXofrGCFJLrCvm9HGriT20H4VmW9vhBljlJIpE+EXt2OPBn
MbLlA+JFcup7pmGTV3T8EIqtNjn30n5XV+/wFKVFm2aBQEhC7lQ+WbnoG9FWFeF3
1qZMteJVi/B64/nmaQrWcHZ14h/r3fqvrdvyGmHXq8arRByt41KtufU117yAbBL1
powl2GABgVsA81v5xMU90uYSidHX+GyxGTQYqM3PZ2ZSoqE3Ow9hpZVrMUBfbGRq
m27gz4mtGBsPmAE/6WLcrgBWhlCF2zPGKbbLzWAVTkZk9oNc7Fvm7FjCKQ9Lo7A9
Dlds7PiLg2D280qb+KFajhFChlsy4avakYHPK4uW2rprboWzh5vf6PLyN8UkeL5J
zRSd4mh3SkJv8LzIIbV1E2UajYGKaqlqTdm583pA6BAhzeT2m1YkIOo6ynAMHTFl
cPiYgkpzUyUMx3JH4kEWi+ty/WoQdLX0l7eEFsO8+YC7NLOjwbtJHLPSQ0JxxNV4
1QNWFWkxUdXY20Qcw2ws6qzCWHmSY3b8ALL8EQJyHLPhYoteM3KxrPN8LLYorkmK
BX0Cth54g/FKu8vjm/pT6DDaAJEx9jtfoRqDBVl9d4AvhX8ZaWMlYfKbE85hBpL0
vROBQ0sL2NHDgF4heh3/Gj1PKJSGioWxxACnGKt4Kp7ztCWZmOyoH0NbAqtu5eDF
R3rJ8hWAu+NLf+rOEPcq8brzDXKEtM8Z0AK3J/g9YaFubfefG1uIMWkQMdzGyQ6J
JpeicXt4H06yetaRVGe/a1GmI5jKf5xC5B/a9Sxcg8Ezioofpv7F/q5Ma28kiGAO
ta9NXIK4RHucHUCbJ7vvTJSsY/Nk/+exzUz/FLjlKMzryJ5p6LQS2VO8b0SAjjNe
aA93piGjP/zBt1F1tDD650oh8QxH438By9hLEOFn6nT5GoIN0Rr9hxZ532vsYHCn
tnT1ST2Cj1R/h8RiNP9nN4QoBdYKgpk3E0sj1AaOjkr0BOtwCotRcNS4lb1UQqzY
zaJk267WdaLMF9YYmEuvvdJKk1cavNXumHK6McNZWB6hz3WUNTTjvJHopJJBVwCz
AUyMxAAVPl57QNQVfw4qPyxWtNtu2MZp27yYHPW3MKmFycyPkZ2IDG9YJn3IuPbx
GEA2uic2zqYg6gWrLJhqMH7wnozG66H10hAT/itoWddlKSyNq6aMS00UYBm9ep6u
m3HOX0akzCAGLPH5/NEuhBiIOtPX37birc6ymXuNdG958Nd2oSGxGjGCgXXhVaLz
qIm6iL2JniDFXBCIjFnkQJTUHluREclC8C9ZyF0MKczxgXSfUvI4ZzF4XAU6ksEF
Y7W/0n87TA9Wm/MH6CCRzTfxI6XVkE3nhqpoeQ2gIRt62Zb8YEsqmLLulS0h8eGW
LsCX+XRAP3WK/vjiqcORkvu+oJIeOlEWqWxVHl/pL0CUS1dH04aKfUE8DOc/YrBM
VzQT15TpDnKqwW1aY0hP7vr3ddCsLl/VsCuwOjS2xkiCXzXZqM1x2sRZKh7XWoBO
XkVzVBfFqHVHQOde4ZDSLg70i31jPgJWrj9YPg9VPbSrXx/L4Ajx318PZgyasv32
Ws4NlE/t3UIY+yRUfOpeBM3IGjO/yT+nDgAAQHSvZ39mnO68941i7fMv/z7aGNrh
IDa9IooZd81/6Z5Gapezn2+EKxRN3006jlbRbDDtiTY+G5O79o0dmL2853IJw4J1
emTqgBrq8cjXSjbN6SukhqTTs7OZV/17sy0XYqbQtwdKqSl74lAYSlbauBuDIFVs
ZLuEE5IXO+aIb+tA2r6RjzIE/iSx/xF0Zk3rZwUdXnBluykvg3kaslHIWosmorz0
d7JAFwM0/4sdF1jD9QcDe+da216FBuJd2q6X+QVaeq4gLa6N1qyi+Tl2iCEobiJ0
MY0YxsYDE+zSWE1wrizkEFw0FkVFB1z9kJbCE+tApz4sL43zWaw73UnLSL+YOurz
myZgc3GBJ/gKEgZeWspDzLiYF4xzQZDpJ6rSSolLQ8Fe5GeZYcWoyjayshC+U67m
nVi8EvJUw4m74AF36b17Oy+NoeZfraR1pROQrdHbv/z+hXMIaezoIx1imKszzHvg
zJMOIUtzwMlCX9InREKPvReBn/zPhpWx2/P+2w6Ij44ZQRPcENO/uEZecWatRr6Y
2kEPT+/zGsYCJjb3fetkG9XlOXlDhh/22Wx7+Fd/GKwCaZU/8Dy3b4iKFVv653mF
TDE/7J6XqtyyaIqeZAnzLlYqxZIqQP455+nK68GFkb0dD4/ULqf/jjqL+FBjUJl7
esccYjDh4DvGrxRVwEo9Rh4ZFkj2uLCV/cAaVwpu+agTk4NKws4IgsSCZ1huDRck
vB/pWMdn8uKseRMNivL9D707oeAhNXHDPDpX1iT2gjqVqe5QXR9EhVmcp7rtQ4eT
+CsHksKwFrJZoR2z0jDXRJTWcbxLKllaVGV/elLkhWfyvbEWg50+AIzPzEX+/W1y
9KhOTrB/GcirG63jgu0Z25c497AGR8U2o+POAugAEedkWILwqFcHOaguDzf3pOmt
MxsEjVOO03sUYlUyJlHtqwY0kHokUOWZwkZv9ITDIk3br1kobjG56ebDdXdMQqbs
kPG//O3ny2SVo47qUUnJBR2WyH6i74pjtYXdaeQ+c000kDFPwa3aTpfmusuAEvFV
SlnMOhgfqfAoh54cc7TlJLtRJkm7vsPRc7I7zJZa4dg4xPJ+EXopDX8FsME2MiRm
Fj9iZ1Zr5JAmDKb6NHoyj108xLBw7mMLJ9T+TADuw375OsELLMySeVDBrTdktQ+u
ZqNUl3e6LN/g3PkOnnIeFCBtRYsHG7Ynwb5l981NxHPElxIyaPl2q0OCXdZkCgw+
Htz/w9otBaZKS322qA11AOx2IAVZoXTw3IvI34f7HD6YGpPyP6BVNJy9VhXi7Na/
jl1mooYMOZw8K5f2pU5pe/J5QzYdOQp+x4bLQsT2rUmna9C9X91Odjr8ccRQ1MHO
ISnMo07XbisIXcumhOR4/xeg6XAEr25d2QAMU1ffRJjJUb5nv9QfcE9mqAvenIV+
uiT7CXhGT7h0qUkd2xlSs0+jYdZ0HXia2kiZ6p3vlHr1epM5iSDsFBKmWB7vX6Ha
HnKoVtbTl8vx6kgKgA3hQoD9qySlBUvgLz1PwyEVn3xiqU4U8Un/Ca96O9zNR/lC
wCLXb6HwptCcpdUOPQK2VuDehLPsik22pNIIjSboJUUaEG9oz8p3OFV+7KFeOX4V
KJcrj/449PXv/K0joeLpa+5AJytPxLBVVtJxxnaLp+0/Sw1ICI3vHL1JYKMXC1pB
xBuqcxjsf1HSZOURZQQglxHDmaYJwnSzz7RxyyPbkF1tCkCJ1gILw7Bm/mK6YwOy
bsAn6C6V+s+QBjq7FrhZkxPPGOuMfRBbsXxyflnFBrioNxlaC2xenoXTLfKBNGWr
dfW8OZ/ecUmpzczdL37NT9P3gt7TB4b8vP2eWcN2L6vlBuEnpH1rMAXly7wmLPbG
alPsAg1LVZMZtMkhqIUYHnGdkwv/JHmu9BcfYu8ijvjb/GPelKabD05PpXmly2CP
XfhCYv6TEfxAXK2+4YY/AtsuUEka98fHo/hxEY1qUsFyl3PHLAgqUez4dx1XR3ZM
yHrKyy8p4+1b4mXjWPMs+3vvySOoHbg6Yh8uI7EWgkFuL2UKEBLA5N3bdg9XQP39
7QVsdyDQ3Yq3M299zrUuRDetPqX4DR5K3ityz2ACQtmqz9kqFMcKqQ5ezE/aNp4F
PdjaTh5tEZEwb2qxf9ftY9c5K9YovvHFvH+ztpMsuonAIa5Tpwv3xm66S8HeBUD0
X2u7+f/KqSkMRYYsFCCg95xnb3b+GTPRquYOmaDFef4EP0/+d2A8RznOtF79LLeJ
pOCY+DbQH2HY4MHpSH4HgM2dIJAUW0wCoKsCrdv6GpUDpC3esgjO9kvmLXOBKEw3
84LWwltkiC9ykbHp9QCUZWm3R05L37g1Ejvc6go1dw4ZHRDaoC5ttfwhMgUR1sC1
RRg+G62zMddBOOss0SUXVepvxUoCsahQfvxaVktXUlNlMfitb5zGo5bDObnyfLtO
K+4zCDG14M9N0CqihcoR0HE5Y8sj6dl5HHFWwNrdqwv0zWJ6+MSfLUJDUf14aSY3
bnyiAdf+prChtKJCjwfpj3QVpWx5O2v97EOSEFHPBya0eJIaHK243k9v4UHo4cZQ
n3lNW1SHCTeeZhFNKRGHZ9lIXImBkPaY3/kHAnkvVheHbdvfOWaYjL31hEgtgVdI
cSlBpdKgCQn+MtPtPI3SquJWg3VCo2xrllkfJMSp0uGXESM4GWaSQg+0J+Gx3onz
okuXvUlaQbC5NMJz9ldGiDr4I32uPN5zrRPY0FDdCA4dF5pcEBZV2ubVr7EZtoGb
SE8FVNkfA0gHu/sKdWJ3mdC7kw7+OEesEBOkHLPiiJc18nHsabEhrn/3D2FM1wSf
AXqcy5gSDY8m7fL+Guq7JwrLQw+B1Acyy5PHUMT/WhAj1ih+kkZQ51pdQrahpDo4
7Oilo61GQSculeFMHYIlqaOXtlGm2Fd/BuK7DTwMLa9cl+o4TVbT68Zswnxjm1g6
Hxo+pVV+0ULFPs3KkcxHbhYTDOmck2UAceqAz1yKGekMxgeS0OZaGHnfaRaSquoO
umRTr5RPauSBkici5ikP3Suy9NZj751hEU/c3b7qCuf0BhWnq07wLw9SbpPSqjP/
81NaaEY1GFZoQlcGkUT/+KfHVjPtceCMMJ0pPrDKjcaOhwZCBYFvfx22uwuyMKlq
d6Y4BB9xwMlDqLDCHM6l49bntJUdrj/T+0ydZ8YedDXTmSqNBce6+bByhNZ0IuMP
q78RTYA05dzfBQpFswSzOj6D519+9FgV+IIj9A6eIw8Gx5wRVQ/ZBx+GWKj8FUay
OlyEKSPbzdCWgFr4BvkvPHTSSOtFrBp636Ug8L0L3AAFhOear3AsW8oX2xzhK+pJ
zqAkWE68AHIT6voVRYG7eaCh3z9q3CIbtraorOaZlbrfP8w5Of0TIRbfkkk6avlI
0oFS5b4d4x7qg5cF4k27rCzexpMwSu/81UMgg2vEUrwhWu+5swHCnpP4qA8FpDzg
l/PllgYCxw0y9emFXpMANzycZFuWMMVdOujWezQrX4W46gYbakgBpRiSEk4ieCYZ
iXddUHT+p5LkOXoS6OGaHU6pIDCglWA5U32pnJ3btt7sfzPiU2oH4Bh/2pFJPs8m
W/FGGM2XtS87McUbnQYfi+MX8M2EsvrDWK+LiGSWRz3bpaWPwufwXigIjcoHWs6n
0h78JECyzlfshCavzqpDQdCM6NalP1RbffiiaBcTkJwGXeBZ/sKKy9Uvm4SrmUIP
KZGF6RDUse9/MfM2UFzaD0AlpldiCQCnqKqNKzIYiAC72bpOuWLMOIJtiw30If43
LOBI2bhzT+E8LRNxLbDkjhJmLLdefxPjIxEDCeovo7ldOOqRQjx4LGSIb3t7juEm
ZmUj/6U7q1rxKQN6fcvrBpdRY59iD1D1S9TOA6mBFMD/E4YygZ2ipa14OAL6sJF+
/jm2oHrY+PDpBXowocQ9vbgcV4ZlDaoGEmhgbxj/6Z1msA2eYyFeyiTayrNkVvlk
eoST9DXnz+yY3MJYepmJIapzu+BSfHNUZNiOhcyre4EpMVnom3zPtf6ptafix+ii
3ZYSpYmwzvQo6NR6SiTFR8zufB5O1o4lE9xthRsVbEJIbq6hGLC1eQE5MlhRaHfu
buYZkD9Bw4lv9ARJFNVf3+/0naO4neLMx9Tn4ZWSCaA+9ulftyrybhdjq8FQqSBV
xcZqLL1YdzRiP2POUm24mvRjBjJO65ZUIM58ztEKTKTpZllW4xVwkdTVGNFsqszT
0wyttvTsm75Q1HE9LtumVjnMlPGVxyECYcOUVWRQivE10oJN9h9Jdny7CUXWkWHp
V8OadRDREXixPwK7OisaH8KJmjn7O0gAh/Nxb0dENQBhUVRxjBbcF/XuC1Tj0SF8
i7LQkhVTdP9U2M9id/p05iNz6RQrcRYbkxkdSBIDR8V3mygSYUXoQf9f+m8eKIqj
oIYmP/TJBrIBqgGUrxhmJIPkKjr9LLogTL05rRc3qQNZXnYAOx6MTmCWwbASXPTs
UiG8UhOPYIa4Ye9B4jGxTQVoStz/Ky8yB2hF7ao6Uvbo+sego234Wj84wos8ijOV
hkwaa1pncCYKh0T4ngmeMWtWT17hmrfnPwIGREsWY5LDuAlUbWE2gzvBjeOiRrql
MSSs4/ndDYwIl3lvCOrlQ/3k4F2S+aQzuZfm59OoMC3MZMs+lc+N7E96d5bjThGb
oLqJ4t6tznIGmhY6GnE4NxZBgVRQROYLtVvQHrWPPgHQj5w0cGC9dAYoibEsScjO
vEBmtc1UwJBXb47/74AwOxeTq0wvQ+eEvc4x8sMKSD5POUDn7TS+yPuo4SyCpIr0
zhI8UzmdZBOer25pxt/xW0sUAbmj4F1Ctq6divqj5WYeB8CD7gTKU2jjI6BoRJ9N
Mi+dTDnsF1ZblfD2XQrV/xkot4fXLtGjeOJIAISpEOa3+LY0RU/jjCcxbqiyf52b
kuBZzsQnvUVGicw8nezIdJDjS8uMRJSwCXdoFSDgagIZBDMuO9XIMq7kWP9D+N7M
0z/giXR8DaD9cQyhbeqG9kLEp3GJurBK5hWdo38utbsC/cl4B7oSLzfPHpQoREJR
p1G3gbjKfcyoXx2hvffkprcPt1qJI0CoXaXoYhhuJ1MzmIdHBBdmEksKqZap3hZd
egHLUCeomVuxu9wMioLgzMewWIzn5/YXzFueEwivfyQUVIB0Ik6hr1lQ8U//hykL
zwA/yAMQ2DAzB4ccFq2jvoxcmsFBQxcYZa5nxEPEaQ/PNGuUwhR3uyIv7vDRbFad
Khuaq71qSQQEuuvarWOJljpPSDQfkbMxHyUiQksXbjICi9O4NEU2fSLDNpX0kv5G
gegbM9reIL51s7PLcqbu0xNDrkvkSP+8UAJteQNh0pGAvjwDl4wEQU/qp8j+dYwR
hfRjIKUyKh8KvTiwBMuarNQesglcmLB2tnSskypWuMO3Yu8OsN6WWoJTNst507+0
7LjzDT4+oV8WWWocOtAlFpyksG+zAt6bUv6/68ruUTJzjwFSSc85LzikgMzOYfMJ
LkZGs/cgPps1ej683r1MUPIEGoPmuKtGw1iqoEhNOmraexpnjDSn2o0PZeaREO0a
2eMsS2Gx/e3KlhATICk0689acdpxIIzlwChTriW6ht3p0GDjod7eFyP95SoTMAj7
n1DRBj2IdolEq6lpuR/aNd71+ONZE1aRmyYGRsOSXq8DwaZs5Cdl1LzmWtGKvYdj
a06P2jMq83bHbq0rlhAdSHvzYKGVcZMyUFnV0CUsgN355g5HIQTtrackFOMVjc4k
xGxjuAUj9p4HX+oq7ssxGjsa4NQZJ/yvmi+ifm0+C9EFUeuNsg0nSXJM/lMlFAPm
ZjM3sqAz5H/QlweV5ajykMn71emC+U6yWVpDZrG3w801z6Q7LoRBdWqJNE5jxcOv
GmNyzBXESL/cBTNl1JJ0v8MuCITwtaI/dGdGyjq6skeBkbshUfI4IRW44jJgCxRM
lhvH1tEV8shPuFFuY1idlEMensCUiZ5DIu9VlkNmtsvcnDpayHLgjiTfkSlTbCxA
tyxRSij+T001qnBDAZNwsH9eJAxwOY7OaDeAtHZFHTdj9NJXdFzT8d+3WQaS2xgF
GrRrXsDyNpt0JT9LlkKwGX6JpS8hyHIzffQklU/pFCYuWHJBoFMsHEHFScZ9hcWF
bf0b3fJgJQYMWyqxuHbKa6lwzwlun7B/JigVAeSIutEsHPM2GSEtXDznRD3efnH8
3I/DFTF7jRLoL0M4lr2MLHkbsY1hkWTl7Nv96gsQ7jkG0cur2UAkxlx9meVnQujB
HKsusSlR3EXGwTIUrvgP5yxsA4zGgq2suuoibEYqMIfxArROmU1s2xXLB3scz2I8
48OVmKAVlVYu9jodHR3Qc2nEpEjKFOWw/C9ZJcuCmTXybhRWmrFSjKMmEQG2lmEn
4RDxiw4GVGR5Q21UC0y/QHzervRn9ijHF5KebB8enPqVtMhZpXhHza7GdHc8nt6C
DMYkefxgc3174H/NIOsVkMVq1mum9rqfiagGtC7aEAIf25F0jmmjYX+iL2Q2Uyub
K7t8mC5BC9oBHaWaGPuiSlVrAZ0EZt0oGL5Wr1MN+TXRopcP7M2u6hFt03xk0btq
+SUO7lBlL32fsa1YdRXg4JN3pXmogEXj4bfWYlVdN9qgDHTtdv7fO9j++Bp2s30Q
PzX1AQVXeLNYsjGD4fUfvejV/v52kyAS9vmZ3SLoRaS/1//k9Q6twF+n77VaWM+a
54XQOh4RXMtHQUk2994YYowvCbTayMj60Hiwb/rMYE1K4NbezPMZvyLe8Y/ogvfr
QzyLxgqlSI8eg1azlwVezUfdIjlE2vln2O9O4ZaGlxbAg/GWc5Way+wtzQplva+5
uWl5C0Ms7/IO4fNFgajh8MCeU7cAFcgtCowG+dZMvuDYnllWctHD+NbSchLcInSv
pi/STuMQQYq8KJqEG+eMPksEIK3/xftP1OQgCCUbfv0Oj92nI43Zjja75EZ2bhxU
570j+Z6S/v8bQR7trzPNLYuqWgWWgv1D6Te4Qud7Vy3FdZOnOjhJnG7Jy/bwugzC
YpyOThR9nuFxMxEbVdgKtvBEoADYftkPUMJHwADGX4Tyt0v9mphhHHlWYfi9qtvn
xsvAenuX3pVXnqUvTaEJXBPuwje4Cih59dUAbDbfOoL6pXkMRDOahJEg3O11p2A6
2jgIhW5EBBYrPcGtBjU0tCXWjE8G36Qbi5ZSx8PzEiFRgn9i142FUEgYw53nqAMI
ZDlqisimlvluosa6xVK4/cg7hHYRaKowfhLIw6OMOcrFcLIC7teV8Qze0T/pkjnP
cFGP4+vM0FP7vAq7TpyiGlRHokEvJGLLfRr4dWovovgfm7KYVrY47HF2RCCivXa0
V9fnm2GRHN8URvOH1jR5qC6FjLgz5PVR9tFbiQnnaeXEn0Z2G9XYw5q4tSa/9I4U
EmhUJvAcxa6M1mMDnrrhlFp4DmdV+aZg0rpuh8I2f9PD+z4//TrcDNAbKLUjwhW6
HxADPXpAJSK1dluhJiaUPLQ8OpDyByE9/G65FiLChV6NxteJIZiogvIV2kOHOEiC
WK6B1nCBAkF50HGPjVNefTZimF/jrtgUEOR9n9jzJVOoO5rQT/kAcjhYOuDXvqqN
Uy3L2pMgsAZ7Gky979DVHQt96FhdNccoY8z+EoaY9L4gH3yqfK1RM4WLVPgl4P7r
PDJ4HIA8P3eapereHROFQBOYtlmAo8aLELlB2kZYnPCzmglzkCluBnzFA5luJeO9
JiW33/YEXWyJWK9LG8VUtCJRaz1HUnqMSu0+JtCA2vavEIa0oEGztPq3j+AVMKqQ
2ibJYhxfKZe6XJC8Lt5zm47AICO7zfSIWwhMjsRxNt/1xQZxq660akE78RGgqSPM
LG3LdJAvqum/vgcSoOZM0uMEn5VV9vd8OQFsBGYSeQ6OdmuMCbRI1Vt+5lz0PA2h
WoKgz+usPPvDyBoaRmiAt3bb6bZx5XTY2IXL42PuxR8OPUjldbGg7gJDPg8ZDOr2
5RSAUR4ITDCRuLu58PDbL2qZjjhARsC+XsyEFwIH/M/mVeHawga44XkwpqC7TpE6
rOsqh16lV4e0PjL2k0T1Fj06i72feykBNLOPHq90S5+rB4iFpv7C4KCUeL1bC03z
OTTXWKD6lKYTeD9grdevbcUYCeDEdp31M4vCjCT5Y8KlNRfJy2/rSw64zFGnuuLT
FitVi3J8C6kau0VfZX8KFZlbFfx0iJrmN7pQkuOFjnqViruMOzWpRl1SBUxk/mRu
T9nLjTWXTC9lT7mr0QfZHRivAwJ2Q5Z3bejrP9f3oNaixPXb6hT1d+vee181rp2B
gubjDgIuwHycufcwlY4YyUI/HAMIHvH91DiQioO5UUGQOXlBd+Ae6VqW4zCi5lR+
h9f9+R97LfO5ZeXWW5JEysBubKg57OGcfH0FyoqXXJxNliaYViQSzYty3bm0ucUA
ewU3m37r6ujcT2NYH3HfusMpTv7xaYkcaiXdlM8wS0TrMSYqrM1IC33b1M0fKiSj
juWt4c5jnPs8wVPyiyGErlR1Zd7tKxSxAAVHDDA1yFI2p0mgd0cT4uDbpdk9vboT
uuLxA5F+rj65yV8/9XQ2KOvLVjdtl8KG6YR1/PmuVGkZs48KH3Sw9l08UcXiSyUB
ZY+kyakiB0FcGRT7lDzKdml7X7RbWsp/dga86rZh69KwW3HTfgHEKTicX8u8mN5o
oCjTwZwrEfTWdptSu/5vfk2MmsLj2Eo52OeHWYKaOa6XXyJ1mkMFW5OL46oqX75a
4KJ5p4g6fYsMi53vM1JTscOAQcFRF7V2wAuXjNqLoa9G15H4BZMJ+aCR9gB1Ssvo
6OF+1hMdSYPhmsFoNn1DTehrDSXDCV8PBoJCtQD5KwSkAt3fXNC5yp6op1gAkuNA
h5VKB11eYgiad3gT+DAPyb8JaBtmwFvMChxpFVBI2o7PlGhni3c+V20/J+/wDZER
2IL74P2kndsqwWP+l/mqCv2DmRagwCVtIduaUomibDKMj9InPaLevstA+DHpghp7
499GZbNO3Z8ydfH5SGECi73103tF6eXa9LCjU+UKhsy2UVAgYUYH+8Lg6Xk/QogZ
Pn3Z8bvY6w0sQ2Sbr163ZCizC8X84O8BGNS7GeSluxxqBfWXcNDTrr1TwwMHM62S
9hNVFElONBBk9H4liz3yGZQAsRfO/isecbJLIwZNFOmrEQi9CpzarcXQciAAT8Bn
t5AFbFbOgjhJAHaY7o+lhzU0k4mto1X3aXo72icw5FJiBa4eyQMRs1SB1ZGJAMRR
o6F9zo8tCP+RhlXN90L2mEd8dcjG8gx8iykEwOVq/PS0IzQSnAhHBkYs8QUSNMgG
7/PBWepfii438cZW1XacaHlvQvd4TKoxZWWQfIlEYjP2NkNk9PreNLQGOvXTkOl+
6WhEJ+2YK17E9ESAyIzcvHogFbdpaUCJKVYlKU9YGkRHb36K6bAVpYLOR2fK/Rg/
BE40NMMb5oZzvfDpvDqdy8B7ZGSowGTCcsUNwRulMQlfdlc1tMBg80Zk8qhlyigb
Li5KrydJPw0o1rHzf2fjSexncXKU7uYW9h/NMA4TgLBWO2Eyn5tMFLh3xEf1sYmG
lcVIE5Vz59Fbvp3PdGqP1ySU2IPSh7Ei+gyljDPZCCBT10yb6BWgX/LDVI18vvGW
wK/V4QZ3cJ4y41CkD834V1qtkhZ5wltYON6GhZVWOgb2wRkwJRmP8yr6pUg6L8rI
io7URjfqzN69n8VBnL69DkUFxDLInYY43r16+1gHI5aCLTZPVJA1q488lhhU7Gd2
RL1cE3+ZPJCpobeB4+lnpUiGt+MzuNw+Gnp6s7/B6xQ78Go/lfG2tHSkld5Tjhyq
vkyaUeU2ttLz821Z4P6J88dHdsPi1OfohyZ0rmvz5DyG7D9WetPKdJXjXPodq7de
9UBpJ/1Yc3fk8NQE7Zt6Y8sOSALhcuLBba4fnYlzYre6nwItIK8oSrqVOQ7OSuSm
DMJq0WTvadHxwzJdLED7fBIgtc8UVeVYk3H2O10kWkMeXlnZZIKupdJ2IdT0V0hD
z+oWxeQQiFz6selhBP3fpNhEaPQ3E7gVApFl7bjN9Va6WxyNUf6rywhABZ6coVUs
9Uq1cXxnZ6ELCIcYgoRWNQBFRuWSiUQGkOYKX18kElF3HrCBnq54Qi4spu540j0n
jRlFfSr3+PZef/ujlyhXxRHqLbVoJjCK5Dp9OUL93kduTQuj3vd0+zfHB0KajR79
LOnfHBRZpyc23ig++MDZcJe281TOU1/tAAT89bvP4OyCw1otSEBlz7M4KmmAw0Zn
8E0Q+PxtRUucvma2iyOEB7PMLR/gHlaF9Ekh2hnzFzgCDndBZBsXrctT+YgBBjkI
gp0Np5xMWSodDga36cHJJW/nWJSnAKbSm5O4i1s7QDqRlqBk5aM2XAdGFiE6y76r
p8Cs8MM2gadWvDpCrgsg3B/r7r7Alb7QK7m7z31ds2+q66jRYBkt4PUYkQDKn4PP
yfVZ4Dd23Pn0a9vq1Ah0D/i5HB8XGhdC6FJJOJGcl67n1AzjTr8HDvcZ9YYUzHHw
TwHNMotQPQzJ1Ec39GPO8OyDoxhS510lfg9nXxhEDnsEJ9LgM2WDdr6CwQb6pshs
eLFx1YNTxY097omuvvQPi7lsDmQ7v01chjQWMVTsvaLHnJzOX5plj0ZmbpS5B2Nm
0nou0VG53Uu1hf6HK3BRiQhEeY7hvNrLtDC8wzcImUfcP8AysplPGqUIKdS3nUYb
XnhLiyUU9FCVlFrYqXD2PN3F/3SmWMEQAYv0Kv4TxOMLJ7RNZFRVHLUqzlyPTBei
TFpLXK/aR5aIVvu9OLAKgTwSirHjp8MOgF7ZVjQRcIAZysczChStKNyLU1Yrxoeb
fQ8uqZ2GKVcDk/dGJf7U9EC9W0boLyjSdRICfy4jqm7UAOJKevW7NA4oFKMJJ1xu
Y4aQ0j+8oZeaMAC5PVaDPTjODrtGqpdjk8ubzPZyonAFE436zLIY6hLUl1G7cAoj
FSCkU1KufjFwhBXdF+Sxbbr+zVL6BAq9O2lln3Q1vYbf+wtGHwldNL2TLENxenS1
D9Eh5WH6Izn7sn7UXfq07O7lDfEo+1gIPuYvl0xo8ZyimtE3AXNKNBYpOkwFfazB
GOppGaQ88lcxTZL/22VIQxVlJehvUxmaA56Jn8AtqTu1nu556f3WIRsn/GeyXJM9
b6rzuyPnesCCwB4tJMrMobz65TBmXAsy/8YI/DY31YEHjdjVtYYV8Sft9PYOvdEj
JbyfIQ1rdJ5FIR5cZS21lAujrvZ2aHDOeioZZLXG0A48BOTEzbGkUjIKH4ZSGZZ5
oSorfusB042cHWGfNkrY0zezVQyF3wuObhKo1abpzOLZgzyJAekkwaZczFYiqnwD
5v8Flnt6HYseT3Vsnhzfpcfd7nJZKGotaYiWsbhvt9UW49W6g7C+2NBUmBrcoq0l
C/UaSf69QDlIv1iUJ9dCTbMDjL+6yGv70O5PNHL0VgtD/7pj5xnjg1TU1eamgGLE
5pKxIvaKNNeJbfnXy+IgsVYAb9sawgWx0+QllBf3ILQNo1pb9q+yqie8J7HfB0XR
a2l4nsg/7iyzXXn8JITFw6QF4vv4VNTSyWwvRQeqZ7M2t4HMBgt9947LJmseQLLj
VJbrs3Bdh7zru7YNz+INhdvHjyLag2UAXB7bOqO1/4kpiEPXLfLY2rBLoqmr4aHB
SlhzstVK5BoqGnXlq4ZKHrxvunnCBRq93NdQKvqJL9wum8Lk+Ea9qf7EMiTYe/SX
XDNW1osmBZMaNg72/hbTIrDaBDVT5Oyp3EEEs59js3DLzorelIYsIW6v9dIXNmS1
5peBb06PXtf1qZYb9LOGAnbJrRiqGERHQvkoq6grgHOJ2qHD9J9PZG/EdD5t1rJb
MFylHCi+4T8yAIaN+CFl6qAxiKoerZBudilXIDw5WY5vfohqtVONVcEJoBZhkMyt
fKoejBIjQSFSwXDKqfW3vC384+wHJTFXEdXkV840y/jmgrKM4We5Z/E4kyUOlCdA
eLDViLPGiFPYn4sUH1fQOV9gdZfiocW4fScft8jeTzrY9FXZ/OCAnaloEdcq6I6a
0EMurgJ4GD7Wx/N5aAYpS401oJyl65i3KwA6CdOCJxPEQoIZ01VKoqJc5N1gsEwa
DGqP4p8ZmOCreBpkvBBRpQp0d820sccC+tafYoq+r4AeQw/YZHwujPhZ8wugbeY4
6O7X9ZrQUiLD9zUmQsT5xPehXrEgRPsS5w/6W+tHglE8VLhj5g7e1BOx9gvMQAZ4
EFlIX3t1HltgMowP66IglrxwxJzqU/+9a/UFJD2YnbfSFxaY7nzZiqYAW4ygj0Yg
dJV92A+H1HYdZ6HIIzJDXzPlVlJ8aZMNysnboq/+H1x0bxUGh6lSv6FvPdU5yZTQ
a08S+Rz5vxXRbRwJatH3u2liOS+5tot4P+/gJe/S4oKW4x+jB3x6qMkX9R7nK5Dp
X48Vvs+U2qQOY1kEuMTEuyCqJ0KO6ltv9DkXmUagbNO2p15pcG1tPaYzf5ZO3F4r
B2a3vRoWFW/nGaGX28ILHnrw+Bk1L3a9X6uB07bg0W4j6KCFXpfEN5JRYuKNMbiG
8kPmtcfhA0ULRYps8GQxEU/nd4Thj5LTzULbaajBQXRUSdxBd1S3mOlzYCpFozdX
g2EQffzPeoLMLDW4LdH91jEN8lrv7fX8lI3+j+H7F1BDHYZKED6xOgpxaAa/OFXG
n1tVdKdDxacBuarfX0ubSEgN235G/v9eBRvODIXozUCVX++Llzm+AlbuK00XEoAY
oTZb9VQJF7YxV7lRNlMUKVYn92lCPAQR+hBd21VuGJJrV2rCZyEcVOlsOPdupVuv
lMk9izdbJ4meeaxgMiIlyJIWnyO/SVdcmQ4kyfzBUfnri6Qx563f3dc2yzzrWIRP
cFw33ej2foxAbg06xG6H13+KkOpC/kGIFCtrniJwJHshWaqHhdSWoRZLFUXNSo+Y
EEXPfNVS3MsMlgvXUZLgMgW5sc64pmH8Qb4pOvXdR6gAnHC5iNerk1wBfoeagQqE
e0wbQxqs0yqefNdlLLSnNJFhmGe5IrCyIbNGAaNeW+o9vu4s3Nrtp5wSIFybqVCd
+mHrwICuXSWVLBgR6cTixNdgUdM4amg83qYDm3PLGIIKnzLHRhCY4q3nsNXfFFAb
9BEYr8hllmXHFMIo16cAx1LO/EOOqYWuUXPBAJPou2B3wRCDmefSUik4acpA/g+1
q89VrpXI+s6z76cpu80yhCnYXIeDvmSYlKQXBsQhe0uqM39eWMUNKzlmXMjzY/QN
AUhb7uchCtSFaQ+H26+gd7Cy5curbmINpfG9IE/ww6bWrZ0Zgs+sv7LwfX/ne25T
3eUHK3lDdbnF0qUjiroJfkV9zPFj4vrxElm2PknhEQ/nMKQLPvG8irKG63GMnoBO
A+MzSr84D3HzDICmvspnbX9KJW+mnshpacE+xmkJWd0p7UFmGGDqzTs7/zuCCapz
XkataOY/nJMw4KwvBFXE8IHYdNdE4iZxmFc55Sxa6jaw0CMXQPfKsMCie6jSEWDY
7x6OB5LefhEBdTVmkkgPHImoDzTRYG7p9HzPyYTfFHC8FuQLFK6makwdAqMVaE2r
I5NbvdKFOD1prw/1+VI5F6M1DhAq5Q6rnb7IF8KppfLqUfZmKZBoZtlzoXOjdHHV
uGXNx/Rvunh5f2kMvhmXF2Y/e+WQYZpszp0rOzo0S9BiHXl2ePH8k/o8SdFrrnkM
hJEbt1l/upFfGZxbkm5xcmqCqUISinUbcmX31LcjxRDl7dzB9hKiXYNwJoGGZuAM
Ka0ODKz32pXEEItgfORLQH/5ckebHw6P37t//aL8zsx0JjPBGE4BOrQMJlDKsL8x
VQ3A2A2jz+804OFYqYISSlU25uxZXJ/hTz8hEv/I29Dm9TVfH7Y7NAT6ULYE8oky
WXmKBO6p1PF5VCcs63CJetQiHG1UTez6DHvnulV2wMT7Ikegz+Lee7WZieXV2pKm
avH3M6NInpcklB16YeHvcl2tdTUyCUV59mBuWxRqqKm8K2BTzTvM+0zJUhbLnP91
9BEszakbjQ4XI+05E9MVRFoR3lHXCZoQpt1vYgodqzldXQaepZg2dyeiO+AoX2Tt
O4SDOcJ8F8z3F0H/vw+n9RORR8yXy/IohnvhrLBlv0IzjTGrJz0qiH4/JfkPcad1
wq98O4Voxe4t1V542ZJ4dYLbEC974KwP27FABEejIlJF/5ofaTXIhkRuA5yjoN2C
/kxH0oj9M7IXnXG3qcnUpkJwMSriYsh4uXgMXBspMT0sP6KR1JK7RX69od2kOyfr
OIcBbZSxxGfZleOr7X06reZ/ulffFDVXpi4eUiycjh/4YIOaxjRQE6yYNZ1UzNhi
tNI2Y+OXlSwKlQSmr8i6UIYNJJRIpu7Fpm7HiP+AdTWPqBB97OZrCgiJjMXAvvYU
/ZxeA3xoaolgnrLXrjxbj2cJoHN4wK9XFXtmF98PxL39u8FGJDp0+6RJepdtn+Wd
rxGyGG1QbW7+DerpKgp+0oKjl3BO7acZOUGkIrnKSnLSG5wI/CSIFzWNX3Nrh7zc
qpkonezse9FMOgya/oDPt2EmkpB3KLemLFRtRp/ydbyZT/dYB1uKrPVhUF8QgxOs
X+tgWh/b48UWgXO0YxXw8G8J4+kkbfsdTENXqdp8M6/Mw3SASWQIZAdtoejQU1xt
LuGtvo+aXOJyBbjpTyMmMut+iuqZqU3mYGoAu14S0WG5J5dJ1Xo+RnyF4VtuAJUU
K/xlP5WMhjcuGe5gKQxQTKze9ss+PKyq8cRe3lbnYbg6d/foZPyAvqJzX6gKHwaG
FiCzZAaxzBtCJ65X1bIlU0lYMh1glRQ03nECyCw7neWWLLjRlPmLvuKemo2dXQuq
B8a5QVu4MEkL6hx7eBOTgonyLpCXORY7M+aivQvSFod/kUc+mMZWLwwWIhZIoniB
x+ybSaqXn8MwhRIhAmni5evwagxSmoCGEkjAsT0oAZmG/upHG0H/6mvIztAjRbn7
0TGDviaxBA5GuLXYUUkrKkB2jzrZz2Z6b33NuGZuTaePqFu2yVC4/OJy9SvqyPmd
Pj2hBx3IbvxquK2VwZLsEN9/S+CbEInOUxH+hzVUbgOSsZVNvm3XWANcmh1b7JAX
L3OTq1xUwwTqk8SlurAlMBcpUAbIk7+0eeYOSLPfPQg/RijZoG0Rhd/nvaoy6wjF
npt3nGCjX6QpJGQ/HJ3ziZzGK1V2CBRldNbDaAd9Vse50Ulf5WfOrZpJoUIX81+l
TnJIY317ZKXM8TxhoI8bkMjZAXaNltmmJvWqBSzd6LqxlV6uFUamM78eXUNieSQb
snHBZp4CF67Vh4xAak0HXKKQOK8yj8lXGU2pUgMO2KoXgKnZdrqiInQ1zdFYXNpN
Q/IH62G/k/sIMW+byydT8cZ9Dcs0sbIbqmKnW5irPxVOgtn8TohubSEDW0ibS1n+
eQqtP1B/qIaQ3aZsnX2mg/8Q//FpRMycT2/rpTAxp0tqI9S5TqUcKbW6tM88zi0e
A8PLp27bFXhAL75pQDzVZfGAMSCVqYS04jIu1AmmMzajLi6HgaVO+M0nwLjOD00Z
e6heLeyTR1A//6zSFunyxNDckrX/pB9Oir0TlQvZ71CMYDTCAVz1cQ0PngIIFWym
El5VJKL0BukfYz0aQLE/N6q76xvhUck07tvwDcyrFHZa8VMuH6wG5uPCggvJvzhs
ttUPOkU82IcnbyJeC5JZtwIQx6+1RnHtojrT8bW55rXkPpHFy80BCu+yFY1HXQsV
E+DYsQhwgzrJdfThFURYIeKMtJmBK1AEyDPMhzu4kaFsNmDkCtjnFe9ihe7KG488
4xCsMMQmkxyGv9XV3PTCX+eEjkeuuL5OqCT27hq6sXmEpY/MQzR0RXxYf4IFvi9U
EvK4pDyv7BCCQ90TF58zfe2IpfXMGtA421skyXZCUp7+3OhQ/XOGCTPa+zQNvbJM
xkkDJnyIIoLYqGKxY/DQi2hp23GQ1yP/zbxTginRdKLJgK4Wc/sg0Z7Sbu6phPYf
y1h/fpdhx5QrHlHNSdJDqJWrDNdytYOKiVyKKFjab17SGoOnjxNu36/Ygc3MbPGi
LAFtqH/QgBNf3vrnP79oMDX3225w8w+Ae9TlVDYaZaQ9QTJ3p4PTWHMA0Z8JMthi
VuOujvZNzWGayLak2kSNYo5yH6bCKWKmP4GqOdfGmX/YGauGh/GXqhVDLKgRaNwn
jsCJp205pWoyqWnLFHDQLt0KJ/P5cKGj24AuSnkXcgKfxJUkYXbZZHrfzoXt9CW1
QCPiowOB0xNyi0oT7h2PSfxv52KBvJ64laVKPD67DthrXwzgkNZQkuZD2QRPjZOX
un34XJezlp2wjpmUINXepaj9gqUW85uaLkfQGZt0/61XU5omBAwS2P8E2UwMnHLB
fBpusa1gl3YqwJul46B2Ww9MtCdhD5gTtwc6trmLRny58YwA/ZkvFumIvE1vi427
Bx0HbWf4H71cJSbJNHY9t9zXZwsM0qQXKyxCmaeCuB84kOcI9VKSpySwyh3YEcRe
Y/JuDy3/VcVcf8svRsqtu4M5qV/2GqhPcsIeNLi5oAv/awyybp2HaR5IHL0oyiiZ
FW8cp637NiWFtPNXqvDwBm22Lu1dVzXzPpo5IbAlsfyBBwQeDmReKQV9bkbWoVWs
OKVVr+gb9zEi54SUZm0Z/gWWWMiMeoJQl63wRZs8G4Jeu5z86nxnM+9Opwo7wSMC
9lTK78PKN3xqHqZTtQQsDU0sEiOjVsPNDeQvYEg4+Et9S4eMIaUvrnEQ2f7LG8uT
mOrWCTTswl7RX8VbEhDFGEozXXAUSUNQnkbZLh4QHO7RWl6jAyBIezBXbag0/bXI
cciKud/CGDocZWH3caN/+vzLfZl5CIHHMbeFr9JQJPrEJ8asLtiDCUDcOIxvsUmO
ufO8qMse8LaHPynSaHdYBqRfsL9ryML0fhdiNqZBJGd4e8Chi6urNYPdPnDuKYaG
GLT9HblEm9gc49uHy/xu5OlNdh0ABZTUUm28vC8NOTUmw/ht67h8qGQoDQ2u9rH/
0Ovp6dmWb5d6iGapOo3tJeLsEjHCluJho9spuizYKCnzkWg6XADmExG7uo+ed4Eq
ynpNd9k7u2KBvtxcBeu8V8DMZBVr/sZmXAy6snTh23V4lhhtPKxA5Z/bcJ6PB03I
Fdkg8fKNh+dIOIct8UdoJPSWYH8QFOi1gniG05p+W5Q++ZN0uQb1NTD/njo2HM9h
nUti9CKBWbOYI2bip2I4whtE2sABydG81YKm5f/+NQm1IZZhdNRwSKh4sqOoRNUi
sA9/4Fuy2kn6UDjKSQCU7+nBf8f9536Zz/lDDkZ7RsxbOH/+IHlllyBuwmuunCP+
FY1vlsPGnjAybLmdi3oBNRFRYOJGZZhUqri5Gw2uO+QUuRsTHiMUW5S9clXUUA4s
uki2J9UtavFl3eW2nNT5nE0eQ/isELR8Gec6NnG2eiGcq/VArtDYoA2CFGxcJUZQ
B64jFWwP/mDk1NjbOvCXTFgGb2887QIRC8kxfj+qLHaHM4Z1dAVM03MFJUldPWzb
+wh5EioP4j9gcJJ2Rq7a6mlilf/HyYZsaeVPxIsZ7j7FqdwhTbbkw00R15wZmJFF
taIZ4YMpSWQM20HGwLm1rNCgrGyOJztoMIkYBgNqf/eU4rfwBXO3bPBbF/8VmZES
E4GwfajFAO0xSdTS61sW1xkxdjWpSlZsbfuA9zT/GKY/3rl+uVuSsrHavztzoKGc
Nh8+0J6DQi6DAMK6B2HZuZqIDuMf0ALSDz5W1neb0/kWv8IMxxsu5PeIZFwxZmAC
LsZzrGVUdl62oLdxyqu2fJBYtPezTi6YSLKSmxrBjtQJDh0soSeZ+TfENhqxdygi
10U359GroelfY4rDUSpoz3YGiGt9BTXRv1AtGMHNhseEEDSmtLl5AT+yI/40DikV
FyPCH8f0COU1d/BYrBC9YIGrm8GJiR1AkGio9ksfmEIb8ubcPb9w+mhEdtNLdw9/
3Wqp70O2d159F48ZQ//CbF4pz8+fmuAxbq6HNCnPyJFgN9fpMviH8dPSLChCZB1p
oMwHcuunmWmn+9iIsReI4tCpvb84YbrHxaKGquvl/wA63x7qxnuy1eDx3lERC5RG
KIAQMUW8QvWeb1zy/CgfSUp5N6onN/hCRX4xZ2VV3SQke7RzUYui/SyBSVKfR/AT
LnxssSE2Ud54RQWLEVpHxrOuf1DoRfTsROxM4IMnOsCz+lAPbBt/aod9QPXJ3daO
817QDl6uFKjdV484RRbFWgya/DAGk4w7A09fAGYDgZ1dceytEbjLRJD4F6ynBj+N
mKK/JoaCwCRLMEKPYAQTh2wvfLWWbOGM+JKLPvLNBl9wCVu39z/TKBNPHsX5Npd8
PGoYkmc/2Zef2zQOTO87emoY/0lqeF0UU8520e24zmUDxN2CIhi+yrqCJ++2lxdR
Z0/pBGEaOq1uEAuv+Jc+ALafcfduY7LRlWv4kHgkcqEDCItCf/KMiV0B9K1Mi4gn
lUVc5yxxVv7ewwHrgZn/gekkfuYN4HqdoW+sd1svVqEhiebisCzigRnYUbEnG/bj
FHGf6QRdxY58+W0gmocDxvRD7fV4XkzpcrURmkry/VtUqpZJ3IpFWZQgr2KPxsi1
yR4MtibCBw2jXzzy/kiSWIanU81z591rq+9qpi/EkVsICqNpe/VkIoTvP6euraKJ
I81ZGcywlmg1a8DzL+nQmcKF3eB6I5dWnCurTv0RvBgXVZprNOXE9uSEr7TzJ2+R
xck+Ws7zhqXDO+KlWdQYBwgMCk5v60UXuTyswQnFFyVI0mkgLSOuSvdgFHAmIoEP
1x2G/42ScQMSWXmA7gH+vDEFNO+zQkYKKdnmuW6Rh6hmhUjhbFyOlQYdAwdJ6xcR
8O2SYy4SGt3RGSjNI/NgtqhQCTq50IhqDH6TMM+HCjN3/d2ePuYLtAvqHeLP4w4I
gSzzoofGudmZtJQCwOaFrqLkbtr7yhXaz7XX9O9KShhriAgXY6IMrlPi+jZJ801b
B8vJMIpZ185dGyX0L4VEX4SGzGJ5un/d6+dmOSWvj5dgTt9x/pSHQaeSMc4EstRv
UzlcKWyJMI4K8xd3tOSofaap9w+Pp3Jq5aTBz0f+xLcTwqVxDUQSG/CZXfjfu/zj
j1dcHOS8wdyGN5Lo3b+PpxfXKkg0HBaC0b+L1Da+9yZz3Rg7u9+4Su01MzXTfY7q
NnkW+r2mMv38PMRTFpofo6avqr8s7A05nppaGEyJpzS9jP5UaEZriSZ0WvCrkdfl
gahHR6prmZqMwmIgzLPeJdr2D1Pz5P8qRau2swew6qnbDcUq6Qb4tBDxofiDzsKH
odnMiyJpIdZCSFvBC2jZqUQXdri/tzmZoPoqxaADSePziwv/Eq9iewWzYeNfTv1N
BXfRwHXIx3tXa7qJfolf7ZlrvSQYOZnEmfIVUCRw58IG/HKh7XsEDji0yW0mKmmw
B6+euLE6b4V+DwFbD2HCshLsRamzNG3FwjmL4C6fPLG4mLkpgKEfzOonpgl2XUzk
9Vgnsnqv+QybF/fhq6RpKJQALvr72OTmUu4lPhgt4mamCefo1Y21eKqbwjSHA2uS
ddQWQCE7qtASfMtDw2XqX3qU5qZYrwo9PFZ4/b6GdaQEN8edyv/c5ykBMLhwd6cN
VAzydNGQVPKgcpQqNwMup2Myyvr0o/rRlczdwc0aqMzm0mXiXf+K8tNTDXUq19df
zKVs1Hq1HKRsTfDCZB5R5Kor8yPUHDikzWBo3oCIArVGIZB+Rwm1mR/sb6AqMolv
QzZJ4JzkcZY7W73mFFVIjsjQOYhR+KH1cJ36By1fFUAYxzfyo8QzJ9DBDnDyx/hV
jDcd1l6keQZ+CDQZOKqL1F9ue99wyAAG0VUBQwCAcxvi8YSLwZIqpEeYO6BDgBrK
jNqmxl47Z7TI7vJ7OyzxhyOU4DcTSzVJ68big4LxhNKKpEtb3RreuSpjTwrIvePw
ybB5s8Z434P6k2WJX77un+1YhMkAnn0F6KKoKhVlx7Re6W5IlaD9P76w54JS0OI3
okjGRsCEic3y7ENT3ToIH/XEfR6Bt5jxFVyD46UiQ7B9PExs0iRargu2NTBlNunC
Ks39QRqgFEoUDQEMb2AEEcN51xON7Vdrm04VyX/J2H74bVfy26paQw/8yUtjgyhN
+olJTEr8PONclmQLUObz5b/xPegH5jlRYZrjLMq/O+8P5nQkRs67DlKSv/DUvabt
/yi5bgqbWc+g0hJgJn0x4pvCKDX+6EZOIqYdGOqeS9TS3sIAXW6kWlhVRRiR17Du
n9o1fuP+MzFw2eFtPg/XzpjaKHSS/M/LswizB2WOGYNPIdyuS8QsuiwZI/hKoQmN
S4nj+vWabQumUi2X+5a6lRqvyPx5IPourCcN6TcN4dNPwtldvOC20YFAitzY6xnu
TAqgYkdLBx2qmxDdBL/Vk3MUTbSk4QLQgfL1GDm6MB1sbAGzyvAc3PN82JBjVObQ
c5t4xJLEQ07DeQwftUUNU7IoI2s21nY6ASv0h7IVw0eQER1pZcw+fF+QEu7nEPk4
OuhS45dNZ8CiTqhiKiSQEEjfLiMw1XmP4eWjnWudqJksTJjApEo9OtFduty4KYnW
89OG2REhM1BnAjONlA9uWExK4NGqLLgCFkOO6h0o+raymoigjkwwmYf93Qh1gTt/
IzR1u2Lqe2QSaHiJvNyPqkk9sk2NWNgKlgEeVVuWNYqWTWBfY6naQqbvisV2JwWE
WHesyIC96DJgV0tKGjtExqy4gxrTN1UYN+bJUHsJrjNshToQjeal4p/69c8+2mvI
x6nU8x4KQ+S6WDoy4h0whjMFV1Ib5xkzPEG0PiuYhnXkte7V3ul+OmFm0BqqDIXJ
t5jlqo8cbqatj+qcl1u6JqhVxJGuH2+siqozxnVMSEtlXeR7Nj6kPDyC8A6W6tBw
bEviCGRotn0LTwgtAkN6lWveGzHOK9ues6CyT6JN7/ndqQOhgly7a7JRNUrwz6rC
9c1X7l4Vu3v429ccUONX+AAKc2nlV6ahc5rl3G6lR9fQXhNT1RNGAMOF0B2f35QR
U9KMeHnoJJO4z4igO0WzY/vDDrmgbOVEXSrbqz0gb/7Q3w5dMMGcvpNaHftaUyRv
B7HIxHnmA34JM1FQVhz20c6k2vyvoClJK9ErDSncpZZcd0lsV8tlWcYF5cadVlmY
GElWYUobfgw2dGQxQV2SvN1OP6KwQTrgeL2c/lp9fKgUh43P569fnNTANdHAB6xy
JEdSlWX3Nbs8rjKBcCUeE5MSIIzOc2PDmHE/mfleDp5WJBzD+x+JWOepDFFH52jk
RPVS1A87AhJOOVJkjIgh8/xy1cdk6IiNrUcacFq3CTJkYIQR8qRVp0hwsV6Dif3N
XZ1Jj+dD5nNTV4O0gpDB51xlx7ekfUs84vh+MR/7HHABwGy9zmYi3eOtR8+oifDG
ZYR9Nc35xcy3awqJhSzag2yqOprhRQLjy4LxGMc5tqXkNtLvLtWnRRdq6GswZ1T/
W/Rkqkyukqmh0GZaB0sBdtbT3zPzFX16Mj1xRYZF230A7+eaVWn/QJMh3nbBO1Fg
er3Kg0ic6pbKqgtOQ5nLvuSD3/JSeHO+3BIEjpH+B6p2baT+bMdRWIzNtj3C+Ya4
dwM76DyY1IyASfRbr/Y2sp63ACspYuTX6OCvEz/OtyYw4csWAuDLQLqsWesv6zXQ
0cCsqIeDK5P2dM4Y7f6WofdGrmRIL4o1nIy1icXjvUZ9Xlj17KN0cGabdlQu/bJA
S/xsizGy3eiNh1Q5EscbCVhR7ORV21+xa7biUxKMU4YWz9Glxoc2a1NUyQ6n5aOY
QiSoX+iYhJJRt4ReQ943X1oBgF/xJh4ZvOdG/1dAcARRKcNDskXLfiy/d4dkseff
69zP+jpCProZNtnG9VeZkKrep3lCNAOHoStmLxMEj1/KPFG07D3c0YFgiKdgN4Bt
ZFAt/w8KAo+v1YR5AJLypRljCRu0P3mFD3KXVii8i7BaamdhEyK1zhHi25H7xzxr
eusR1+FqylhEIQsncRIxEo7L55YrEDr1bMaIdED++qahmG4e4PlbLRTzPQCFWRA5
7IewyxkH7WtFHb1Zxsj7tLBFUgZpcZouiXEmDsDFbRZm3cOXKHzPERmc4mMrqjtz
vlZXVPyfv/WiHkTssAB4vb1jbN4mQqoQNRGQLpxq/++TUWjnT67uNIMZzbPNf/1d
PubvqXNAfEgC1GdD1D+Ti4T0Q8Z3d9b6CwCF5kZRg034mC9sMB+uLbThTYgxzP0T
fcXhvoDw2Q5zQONI0wBNha624fNwkAxFL+b63JpNHNqkPT8UrFoAMVmatJ7BO3dL
rSd//yk4vtz5jQ6WMZAHYyJl99Oi7jLunjEoe8oZGhxnUginqrxhPb7H/cJHapuG
cdk/QwbimKf1FqhSO1igScgW6baeuM0vYueQI9P3j/Z+tU8onMRhPy6mqu9WVUC6
l7FE1FDE60F65Ip2qD0KK4JfepQmXqMN2ZYTNEfpVLhD/VjxXtyQH7+2q+v+yUVG
9dRNuibnhXSqtUBt4wL/nGfYU6WDOs+lYlMk3tXf46EJmZJNeeRbV6ScIgaP7aNw
bO9/zmYq+YRtW9szCzqO+Qwf7+oKEoWmclVzGLs+ty3Kb2KMNMv5W5/cvvV0CGsm
c2zXVKB3S4AZOLnql4l8oNajSfgJYkbMmNRRepFyivY8wf0qn79kmS7HI36Ibz1s
cMjfpvzYxtfa6dyMA4VNMH3IbAb6hIW7YqQisswRMMApKckyNKaf4nci1nTcELhG
bpX853AECbj3RFQD1PWe9YWWKUBUCdqJ0zMxk7pAHoR55iX5toCG9jWh51BSzXXw
sfSRlv6t5AevkeB+7dMY4kpcmRYFg08DE4swECnaO4KVl87903ThWr34RIOVPem1
rrzoQd2GtWYxLpGsGlRxF8mfG4Yk8lL7X5A+8f6TpllOERglJ3M0cIhMUK7IkNks
QJ0rSl3y3V+rdZNwHW4V/UJh8Qen7rNqYGjn3LS7dCntdp/RXV/eg/2FdQ9lo+wl
jQbcXAoZWROcF/0slFAxrYjSLNjF7GH4cAng5DQ5DGWIrMyge/B1WRTD5UZIRdCE
Q2pi3eYyb29yjJmnlepy+pYuqfR4E+K99TFiqytLCkMWF4WTbbDztMo6FkQxclwc
9U2wv0CTOwJu0fgTULGDo4HXPM4vlaPhqF/u6EH14cawzhtb8oQE46s2IpjSTz8N
sstZiI975dp4ItZUkENC2jRDi/oQmJmq4lXlTPADNvDb/iEj8/1/BwmI+U/Hvilm
+fcmYjpT0hAsYtQB9CiU73/XSrfkZ+JCJEF+x4d5Xkbk1GqJDJUYI92dyZalwhRO
+f8Dj230rXZ0K1Dr//liHGhVXTBjS0OjmceUCm1R1gEbHZvbx+R66rxV7gacmsnf
7kW/zg7ZvFIm2V0jRwBGNEaO5Tl7CxGXT/YqUkdlCEjixueU3Goxfn7zUDAPcydr
TZBJBrQ6ZJQD42dWTvU8pXUG/eAtwGbnWrrHFcuRAaoQzI3TQaJ5qxPUkpK7WD6o
Ftr/sAKzqUjxkfuODt5di3imOTnVGERzMsCHWtLd7LUHE1ClI4FAsAWq0rYzqFBl
g596Tn+gyE1n4hyL6523HHhv4hdLl0+DLzWgLjdk9wSVLelB73T3sHSWx5B11Trc
e2mQxkwd7w9ccAArwuY3XdnYqeGErGHHLavMFO+7/XhHTtOfzjQBrQGjXU0OFPv1
v5ER4dg5voi+4GIQ4HPUAXz31yg/sLBi1W6GFUEScdzA7h+9mGabb+sW8+bLDsIo
fryU2Am+NtJjCp18cmf+lgTZBKuvXtmuKOFMdLiIzRZ4ZhBQ3tURV5jtDArjB84O
JMzMhtz6Ki94W1wHUb8KXd/KhDlcXvu6OPpxQcAc1mQAatLVzIdp1XGfbWTqoyoa
a1Z32Rn2HXqDOKcs4czz+Lts4/9da4AWft6IwaSLn2cfEW0DrtRTudkFm7WAX8Lu
IDVR5gnysgAuMnvWy+lkHqXBQjNHaCeU8WD+6kKtfROqnBISumDA6CLIEVR9d8um
jXWzb4mUyfy4Gf1QQkSpJwuMMUesoM/leaO75g8Zn0w44ktH86Z8m9I46erxGHP0
hCQFufWglXf3WsJLTeWv/zAWZkEqk2FCvxLPLXNZqj4bATYGiJqHOQ5V8IG3oVGC
AuIcbpmdZH76mk1pRtIlCSdXnI8WEK4fIRFSHrvlFBtMmic6c646MPJopPF2LUjF
OL2XFOikhfUkdMP8HXJIa/0JwuviWARVEFfdXWAFA7Y8vUtwnA8/P/IF507n501y
zJJU7FUSv9g+BdojHo6p0zFrTKlMPqRQUbUOwdl3ysrZRo92wnNClKdoDEX3JUp1
cFHVCxXdWEwNveP9vrpM2CvhzjXjWetlac8yz6aYQoiEX2YhlOSW4A/h3ExHmVW/
YsUwT/VeCvBStuN7hhefegKooDvElGmg+5dj9b3pancHZ3/6EZv7QYXDvn6dxP46
70rZHHBqV3tEAD7dUm8Ucou+sS6Luo9P+mBu1WS1th5+1IhRpjTpU8Jqg2XJ1AmL
YMpNgkeof1C1L9pTwUa96UtIMtvzgSv83y69XHOXt08MjZeTNwagKmzkw4eynwNT
avI5fiKsW5uQOwEEkrXk3yeE3nOdKCB6qst6VYxP3XmBw5F5dro0GKCQphPgU/D/
4zBbuxP5WDWEX52iSZeYNQVkPjKlDTq+4bKJQ6bfZMeIbaMIBnPI5pfo4yUatgQ8
dm07XuF+kM6YgdsTSSwiW4Nbe3GhwSlh7E8ia8byFRoU+S6R+xq2qgHYzQTd1Zne
voNkKX37BA1WUAOA57ye8twk7ODBr7zIWzXiusccpvz5IzeqVnWFSQTRKo+Gm7NO
+TPR/N0EOUqMhUZcokNt4Q+5LrAo8iObEY8pbMP93JzHF6P1S3e3G3i2DNcURKnX
/jvt5JUWITmyDBwfNMiqvjaPX1+iuEnrrsUR5KJzT6Cm3Au3hd1Sz9sq+BkG/WDd
0PIL2cVAoMD6XCG8kAysZEB5RLFprQuiKzVQrPVIx0ifTJXyJw/dU7KBg7AjSoUs
vmAIobQ4Sw242EGqOUl8K8zxhV8RpYDiAiTvgu+XQxdiV1/dvtHnYY3K7gDPsWFh
Lp30wTiJYlblDtmZpCh/LSInpmniYF6efQ6XmvAJKHFnSRPh42t3wWPmzjtMKI8b
HcZiVw+q+iiRs59qZXLX2NM2q48qlPXx3EKd/eGf29LGac19tajCDW9P3MyNE1xE
CCAxQyMpzFmuvd6vWHLgcitzpnnppLldW6hLNY7UY/6GXl80T/YPlcs8jJpo9pf4
i55Jl36QxXkMxQ7yKgenStBxNhYtKEHJmpcRc8KWZl34jhM/1ctNgU/x1OD700jP
mkfcGbMKRXJ1Wjaz/IdtbbahtC9vSCR84SFZTmGUr8C/VHwI3ti7g5G971vcG2/Z
qvTVuoobZVROMfkOSlIVaZTeYBuZliJodOd4aEJSuXxcxqwXeQnflxlR+2MmxyoV
auJnFPL09Kg3Ckm5t2ycgwONgrPKXB/LifoXqIRocW35jQxOURefzNn7XbkiK45i
I9bcuLiO7BqvBhc1/P4QCWzjqjzw2o0mutJ7EntYvvLZ1/BzwjqWdXC3ppUxej17
qcMHEmZjUxTSWQY9qyY3tZfzD4BIAzHqU1/dyQGd7x5gwZH7Hs1uhGiYN6CF/555
kMukyfRMAJ7YZ44SR9ktCAdKvdtW7Zb5kmLBczGudNYocGNfi1XXTNQTdD4NGXI5
MdvIGHGotlD3eMojtEs1I1EfHJpwwQSvEfuqFB3o3UDV6NnQm/zH8Jo0ueaDdJY5
lmDdG7dEajf3FNFscekP9an6BN6Ds3wdkgWTfMKDmUj2FMsnCzcPh2h+sKxfoNGg
IfjIpQWrdBtD/O3FYJeR6F/KGYO4O70GAtqR/a3D/+2YnBFZkwBvYVF1wGmQtK/W
FdeS5b7Pfo5qhQa0gpA5EV9a+RhD2wJGi18l4kKuqcJtCsRoYldJx5TtT2uaZwhg
YIy8XxqKoLb7ijqWpYUhYmexeiwwBgjh68wMik2OqVsOLYmFs5MGuDMCKo/fAfOr
T78TSwM831mFv2CLs6n3Fl2IEsKc7B8Cor+Tl7KwTPOxO/waEjzYehqpJ+NZg3AJ
vGtIWVOfz/SJBjGXXkAjF6h+/0k4AJFsCNin7IMRaDXEhbu5PausWV4z4+ORT/9s
p53oZYEOVPLFVCq/w2D6tia+tUU85ZccP3cFOQCe/72P33k/EE55XhOtCPmgH6On
pIE2tKtqt8/Gn2/ocyCmhUX9DrgskGdcgagxu/1/pKFlTDQ/7XdjydZXvxCf0ven
+vaDkt/8eC/6BP0ju6Cou4wrGqs/cTSoIHsvsAx9MTnZ0Yyd8e0ezDosZ0bgO2yI
WMAP0nq84ZKt0ljknZlwb/TjlWRUsaZxQh+dx0GdIpcF6x2Opm51g5NUKyAFqfXe
Ila8u1142fiMlAstopt5xCZK0d3T0eRs+xQ59+z+0FyfE2a2y/aCYdWur3CgrtLs
+B9ehrMDWWYcnPBkUohVF8nByd/gi6x4IuTUaumcmUN9jJlOz7AvCjMlVOIAeFia
1VBnqAMpF+1J8mUCoibLRaOgBu6Q7ElSZNv4Y+nf80Dlv+YvKXsfI/DdaFidP8L+
xFdjH7PmLQm/TZ0YG+/lZLj0+lIQ1XvQIkkJhuSjQxA6TYRLeBJA3c27OFV0xS5K
Ar9gNOpfdnAVmRz9PVjVdwTJyp4/ePdsNa9enY3hXX9t9tprdvMiO4liaufK1Z49
jCIU6vm9ouuqj4EjDyqfbF9W6Mk7Uu5KxYU988mnqjJjR1oMjkGBccrMyLodd+St
OaaSAFJZEHw61kgX91nCBW8NSKuOf+erqXyuYtgc+8vp5otx3L5Tpfa1X8KcFshu
fzKnjkrRPKuz1gesfpA4bFkxqRfvKwerU7um5F9q8TqC3n9y30VvrjExalLCHxFd
JMtCWidHAiklguProeVwjJFPJ3ceZhSZwn7OZ8ZIa74uljmvxVXflkZzfMbO891n
HownrW3LKhQ857L/WC3DXSar1jREfhQIYV/NeCH9OvamOz4k0PxLrIj9Ka+VLS1R
R+IF5tthBoZkf7YmNeFGY/owQcei0k48OAkjhpod0V9vgTQaFxw3vKLJO3q8pIRC
oV6v2jAz9LNm/R7thfnLCghDMh37LjFW/wZn2yUh4M6TQa50kvLnBTgTlerbq533
YX0xXCUfBvxUKf20+i88RNpesjcSC6owAGwmWj8cdI26X0IOZRd+/NM+7Sc0vhIb
Tc1wsqjwHYkqbxr6vYmjFf2YqDiByEeT9llm85qB4Tj0cYi0x/cHbyq+dOS9tzf0
QzwfY84jPi0OQv2XWMg3eAXmf8I/jABj5StjfAbHCTeuS0hPSHqBGCV76umgk7Tu
FWGKYvZRPXEU6pAPSYgy4S2Yxy6/FdNgoKSdBefoWYHVLD/QL8twHv7HS3E/nYxX
lwJgcEJO4PfJoY5meJQdthpCHLwewZS5UM4aFII2vVTORdYnhF+86Tu1GLRA5GWz
DbrCSf+1exlM+izPVnFHC0PvC4My7xR2GS9fPZ9muImWjgMLGvEOn2PRm304BDH0
M7HIIaaS9w3yzM7Dvf41rriiZxsmjZotUz/hhXRNwOZtrr2F6sO7F52DQoMzElMC
ZZgPXyeQw/W8RRzJKtuy9jkB/e3x1JaAO4SSGQ8XpyIcTI4sBO5wP3l9Sa9HlBYq
mBP9Z3BLwgU+FHFBD6Sbfc8y2jv5plDEK6lBy6RuHRCzStrEud/mrahCal8fAbyB
jDPeNJw2/NPLle7bWdeAZhXm9GWHwZmXCTFi1j3jGd1RGDG0fVxqWk/d/dmvsk2T
H/FiOIqq0m1PVP4NuZH2L95KFNg4PszU89w+SarFkJJv0hbopfIZYfRV99xQMOoa
gT+Ty1/X9FH9uepxgL0/FZakU8McmyRU4odK+8Th7Q3vCfqHlTeNBD6wqyozmiaU
lZ3U1iNkbg2dsXhvklOAbR1AAd/ZH/nKt2HAkDY+NDyGQAQDm0IhRXXUFW0oApzG
dZY+tYjmGVZ8+fUks7dDG6xm61aAbo+xRYxlGw3DPHsIM8mtZbUuYU7i6J8l3cjz
Aw5gzGY/QkeWDBEbcEyr/5++mcTVqjk7GC7yaa8hVP6MtEKsTXLcalZNm1kxJCyT
u9GuRdbdztsyuX9fW1OToD6X7+H/i7RBkdAMQR9g2FJABnc/olxRFdS+WvoPGHAb
oeRioXPB/14rgUznZAL+EfamXhXya8ofZh/vDyAQsvslZt0qF1Wr4Oo5tQdN6tNv
zf9wmFguScu7OT0P17l6mz3njvOWUl16naVEQ7EAbEsJgWp/oYRISRJlyVvz3iCG
UL7ijJ6iLzVD/FkIEtIqNv8sxsrh32+QylIk7Tjh17z6VqUKU0cw4eiJgFUWARdN
WyuZFiseoEKi0kLBQjR0xqtvBOabmNjBCwvSt7VJyKN9qSL90qHOLX/RN7s3Vp4m
BRRR4RL710lb0E5R3/H/Rg8k21X76n+cWL9Y6pWuFrd2BDl7P0d8epDZ4njTfJ6n
eemGWzxHC+83sdh8A7qMXamGJWmmUOO5TY2SFrZCHh3ueItjG9o5JrVN4lK+i3SY
+jvb01Ula+WjpibmBwmPJZ/lSAu+pq+nVEQVp19SroApwCLKcwruHTngtkR+ajZa
4y6o/LrVz/+5p3MnOQwRhIFaAwRFBOo9Txksu6R0CQ4gx4fsJhW24BjxwMkbraUf
/qZ4XlEH/ou7hH8SjMNWklqqQoYCJx+mRkXot6nRXNJmWSECWrQTX72vLRGgumHY
TgkbUEzg0O/G3VJhK+90Ci55LtROLTJbl5wBwdiC22Kto6X4lekBDSGhgbOIW1fb
hbmR2pwkzjUU7le/qfUTnO63Y63wXnZXGjbsvlt9yDjM+2PN2i2dK0iktrKTh61P
MTbW0DdC4+mT17+ABB3B+mkPvkZeoWLlQTQ7vsdjbsutHpXTnYlFPlMWeBBlqOGd
5aSd2RwfZO0N2Wyzn+9EHZCSuzdV87faz/GJ+RE6uUA4E/cRWUU62YFp00Tcjx3n
IhWeq2HrAJtBQoPGr7078Ylro9G1qjT0iW6fqqd7WHjEnJoyFSKKoN3J+bU0pI5R
B5WObjxYoEaL7y+k+fYyWBuZVEfaGmuqXkac0nzdkAJyhGoVUwgyHdqap9Yujn9p
HkpQ51wDLKWRXYYunpBOU7cFMVzdnltsUgR0HP6bFZyWZ4lGYSweZuAFAYTcmmDy
/PQVCZ/1AhqF7iVP30lULBr+ZHEX9/n7Mgl2atRuwRWjkh3khusem48Tm5xEMmvh
BSU6CUeHd4THo1rVch15xXW1/ijMLd6fOkabJJL/xBUvP71KD3bnH2cBNOqOp/eW
bB4wUr83CRskgnWY+Nm0D1yWbGGpXf8MqUtVNQL6uE8ULBP0XRGaU4xN2U3Ev5i4
dak8WIk/ys9uSpaYsktpIffgZ8Cmr+RYjB2iTNKXwVry8XJy092IEgO/Vsge58l1
lg8fjzuAisRRYtxuVzz46XrV4VlYv1TcsMFT4Fb4hvxfKS2kf56kVEadrChEePKe
v30f5Jq05wtZ7MYyT5zXbVpbZuVQTpPduoqs4Doq5MnF6k+kwv2/etXcILZdQUr3
tBbat/+UHad+04PNFIz2SE/GK2CJWakjGyjJHSNOIRg/m8cjVyoNxJBt5002IhwY
vydbtwWJlUQVVbLQsUSGwrqZXYJOpPehebiJ0GhPBWJznE4PRIlTPLSDKVpgnvlt
lTx9XaKBVRRt6J9WNtn0gD+GCPE+hRGoH4uNFr42fNOUYTfRVLkOOso5iFcJRUEP
eLjNPaZOwtTrfY769JeDdNyYoaCjsfuCdTznU0i1T5NwrH2rJFGBg4h0Vs93tohh
OZ9erGV2Y7iCLj5zrRh/fPSdDKdA2UUJW5zUGZUWrEv2O9aAwjDu4mvjpuKaxqbs
ABMPub3SKQ/jYZA58d2u/japULTwiPwkIDinvk0+AUNy13Y4VTKSm1NOOwgrcXqX
RGFhs0gcQPsuMpFuxGO6Wi6txk0W5Vb6PVkDgewvxm1o078L5pQNIkHKde/1D/8V
eVw7CKgjSf4ZYaeIjpQNNxwT2tgr4VJ++hI9U6xEYmw3G7Z194yD2uwWRXsDoNqZ
dMhiaQl4Ud/mVQUdSQt6mBUgGVi/wTgxSv4QTGm72uhIfxJdaNfsoO5X4VhuglTa
QWfIFNXUt58yPdnZUT7sVASe5CGzhn0Fbp4oIpxmofyImmD+wXO35usBHpUKiRcN
CIHZNgOhK6szY3plh4rUoRxs8RzMk1Gt4wuaazLghWWuCrCglRN1/E1z0Sje4UVq
iqgvDHC1bYzCDRlj4v4Pad+i1CFa1iS7R/yERVTb/o2K9hGeZKPoFuzFPS6kaJxH
Qvv5UhVuEI2iBvxktRssamdsL6kDvV/Sy3n/Em9XqeR0ETD4+r9CU0Z6NeLuq9Z0
+04CJsaDHdNlcVrZ9trZEZz9HoM4wZ1eJZPMKGVU9pFuEFsm8djkOk54+a+oq12P
IPMmM31g0/bcMT9TL4GYDzZ/8LuTTVr6+ahvJsi2sqdEnqMtauK0DPMcSyuuNOZZ
LalzGRVdYnKddKdEmHG0bpsV37QZZNW3Ny/l7h71IIV0BocN1osV95wFWA5tBSvY
XlPRWfUWcdzdSpey5KCLfqeYhekNWfTx3L3ZZ8PfqmcNpiN4xUrOF+dqoDraGcNq
2gq0MWRiZzncCeXOkF2YPr/Yqfq9N7hHHmnQpsEDpA+LIesQfu0+03j2p7TgwzqL
5I+8LblBjczX7qg6I50gxod5GTVTSgeINMLDMg6aBQ7zrLTX0CVzL1cQ1JsKqEUH
CdEqizTr25fOt60fJhywIprXU57IIXJekEdAw61URsczY2SnlZmoZzG4MMO3RMNr
dQe8BzNJLKEjLyX80Myr57hQem9BAzTfPiaiWQFrAc/rSFjgSrgPlTCSBvcEP2fC
i5lpNayqTLI94h1yEkObF3ES+uhCIlv4QWWYe5RvSJ9TM6mlF53/0H/OD9yobSO9
+VQD+lV9BfUQdTFsTWizOLNI9oExeE2bfSDs9bnwVlaYo1/7/1lnBGxYYUy2WmSF
4uRqPTJavTOBFWxOSUuu7okrM/x+mPHdfSDORc7b4h6LUv3yOateScy+6tmHoMIh
qUgSJ7EDKaXf7oE+z8fresbfHOqPgBAmjl9T0Xbssa0td9q3YQvGRHyMJAJW20QJ
04lTobK30IAooU2eq5nZJv528qYlyGiEw4jDZeiQa7xWr+XsjTZsibZFREvj50eV
goFvIjYfXOF7BZW5vgohKB9uL+n4JyFnmsuWgNP4AVqdTyd3rXfiwKeY0Bd8BD6D
dZUUZBBHaFhXiwVLLKMYvEBM6RNLQ49hx76NSLdSgw4MlxwSR6+XR4mwwObNIJBA
4BtxB/fhNifsAM/8FaDl1LC70yfhw7eJw97M8adzCDZ516hP5nBXlW/MQ4M1iJLp
5fm1GGrEQjrGzrrzcDXlIz97zVY4qv+ExbQh1P9hX4pxBgqqdlFsmQbytYlz+Nln
9c9qUlR65Rv+2hALAl0KHe1wnZxOQy4ueyO0GAzop6HX+2I5AURjYt4dPwKx+I2S
PxCWlZg3iTpYLTYXyBYnFPViWQm7xTilU+ob6xBO5s5MUQ7Q3/xKfK66EjlawosT
mRF+65hJezml/r0XXh1tBC9/+sTm+7NnR7EAlP5sbuy1vZ8XuoxPYHC2gpNia6k1
8uU043eS4ZM9irnQibAoTJj1+QxZ3pxGn6hMEnXRoDVpor0qB6WCld/pSW6OobYU
ppIm6XWwNu5ABPJbpA91wx2V14TJrM2mFPlm8d/AJtf45lobxuiayQhUSBIfb9qM
pNYAxCZf7hyWcscsKBkHIkb/6qX2FFjFEdLp7tt9Vqh2x9Rj5emQ39+8d4kOq9mf
fGWVAx2nxAzQUMyw0QWZnVKcTFxVirC/MYUOfKfX+u1S/RC5i8wPcprZDTUxHPI7
FT3WJ0CajUp4J/vTs2lUgXkJd9KG0Stv3NVDLHMd9IBrO82AHg6Jps3vT3mrL+OX
UFuuZzT6HDYLm5kDo5bwjPkTzKTJMT7jmgWCGFHBho1mqWMekWCWoKbScFQU0F/7
zvlCS6W1hKGAe6/CZ2KkuwMrzU2ux8kvlS4Mr74Xawglmm3BeBKslLcXG9C/Qjss
Td7x7vDZNVQMfqhFeHGFHsM488Cz/Cbl2mitcm3E+JjrDODKvtjG8kLWsqDwD6Gb
dTbGWirYI88nDU3Ii6zHETDxW6pbzr3Cve+LcmR0vGteLUKI5zXfHIq1fj3uCrdR
BgIR1mUoZYBF0HyMyHYYY3lWWnyA0xSlZNhEtUKwxQg3WExb9AEyBYXm2hWAAzpA
GAp/QUwDWnH0Q5sa9RSudtn5xCx/1HNKUnTlKUuA0PGEtGFtbnGYCayzlvj5xnQk
mOO/Zsj9Ukt+nMX0n1TF5Qn/+JBn7MCtHNWhDYeXlMLI2s8KfbECPvPAbygotoW4
ZgrTKJg+5Lo02g7xRR+mTh7rajhBbw8ZHTuzmBMqU1axh38Er6VLTt554fVzuaP0
SYveum1Vo89BHsvgXlw1FX4OylsT1/vvXMZnuZXwsnUEfZ5YOCwvGpYIajy6OBV1
MF6iRQbny6S+8epjBfzlUPj8Is5n8x8QrCM5pwIdbXUvOybvJ5HNgXMzNIcRH8nG
ijfXnEFGIKXBa2c/L+MM0TEoMioiHBYe0p0AtzYnZLlxQh7H33qcEwhItbYzrXrr
4YV/2U/EAF7sJJeZ60ygnxGyuQr6kGvxiDw1L10dCIkLw9YxRK+2dS7vNNEdbjKt
RC0wGIAOemnnnPTYdbKoYOU3QrPDBZ9xGXHg35viefTJaOg/xw8L6FvmILRFj3Jr
9fabXMS4fDQK5eUsM4k+yh7Vi9dZRHj6f63ljjN3GhfpR0GAysdS0IpSpcLYKFnL
r0oEADi5VE69entMid2QXbHbiFCexIHE2hWHiJqr9RAoABRg0n8oHpX1QSFraPyL
1mSUADrIFXhl0O3Iy26a6muWSe/g0sY6dIpGR5v1EcjZi9j8C/UT6aG90/Bt3oYF
jzopAZchejjQ5fr6JhR4a5oTkQpGsrNxsZrWvEfo2ShIBIUGvbR/+M6qTReGbgQl
DRihhRhDxqrvrFSJ5qregujGYNYQ181XJh/BX5DK9LgRnKfR1hbOCfwheL3bhFRC
cSasa1kgy05+b0EsQtWgnVT8pAjvIFyjY9zriaLRmCM9TlF3C6BcdnyRtBUTf8iv
PPstGst5uNkLiBKdpkgXpeXgPdYsod3WXgptrD4mfoCVZe5814BUHFDTTnhGAtep
N6ehMGcjGZF5OpExaThKAa+Z1gpmuIMoTI2xDtPUGcG1ZpOZufD2p9gRIPWYgULY
yUK4R/NnuXeI4K1l63dLCLnZrEOoGMKbMxw7QrdLsiEe9LE6h0mbhi/+VTJ9N8bX
CRlD7kvMrRI3SL6MNex+m3gXN2Pt15ZtLLg9Q0LGqPT0Wo8DIU/XS0uLRE+g4y3d
U6eKIgVo20EtiVLjwH4G2O+xQZ3BX+X6pNZnSUFwcKT6G7j7hOufVVbF5oQdACil
cwl/8E2+cQ/pfAyLt1H2/NTbcdQQXeIcbXjuXzeiFI60WQ5y80XJCfwksYmY+iU+
n9K4+RA/P7aqz1EIkqvlt9JOqclHyOyxIKJh9N7y6C3KbX4zrHhYvUm2wOu3eSxV
PiJRrg/F8w/f24Uv8wj3//WsIVHZl6cXr/MMaz1jtM/pP3LfG1ZWvgNgQBpHZ9fn
981f9BwMCsrnicOkpDDFsswKs1AIWbqyT0plhEbgdQUogeDgk0s4kOdjK0Onl3Yy
QG8pRUNz1AL9RAG8ucjH0/4drOOtfn4LuNoNg8U6Pd08KHDDavr20j7RDFiwE8lU
0lyQRDiyvoeJ9M5MjXJJpgtUXnPGXPwMAxCCPcKMW8+Fj5w/D0zenGcVG6Yr48ts
h94mVPFHrnbHOWh+dnRFAE5SC0dWHwyzVARHCMW/buBX+oOgXqIhC/w6sQtH/v7c
GCNtFWqSEXBoYvMjA1veK1d+mgwOnPfBm5hh8/buePcHjUd/s6Cgcf7wcfTbDiVG
/7XfCRV0ldOtmkxfygRNZrLhtAK+a3IOljQW+2e6pdtsexMFSGxkJZ0NTxry3+pt
c3bBU2YjFrim+fmXfhKWjaUGf0j643WqOsA2tQZsTzoO96jzL21FR2xOAIDqc2Q0
DBsIxmwqQs+cb9O4YGUY5x7UL8gy7Qj7C36z8GAwQOiZJ9DzILdveA8y6r8bB3zy
KxRvp6CrPfryhl2LKKJF8sskGO7XBOl10gVzIH3X//C/WCcRDay03H5HXdyLYi+h
nsWAdhrbyXqGeYr4uNZG7NSPZsVLWkp+WV9m4FOxfFhE/dpZ5mnfcqdwl05EpyR0
PXMDhwwtVx0iSzqt3xyAxfLO1HiDQz3xRJcoXY8MRto0XejRbrrHbVUPqPGqfNM5
OnzROSf+mxAQiGMnqkfBopbzfzHiFBe9m8S5yawlNZ09+/sEs42GpAoPQrhvcHTd
QlMc0OBDchu65AJ+Umy1XpYlZlZGXvj2GxhR51w1eWyYFZQXwXiq21Di0SqXJ5p9
J13qL0PU/lSWsV6xWz/fQeW57hYzr+VmuctrKD0rPalduaCyyvmxzOBMC6qcx9od
hN/HmunN8QwsIg4ROfrJOGk+sb5rFQZTYOBqmY7kowMZRplr3m8Vz72kCPXP/SEN
77/l3iPtJn28/jcwnXF9zTPXj5uyv/eXZzxZ33a1mLdUKHczgeWgf3cQpf/UBtoZ
Mm/fjiwe081+oblQOKi4tBbPKGY2zCnkBFpWWGm3M8YFMwqqc0daigpyx5DGOGwq
qw4xQpzVfrYCf96qwVirP45DoiQGX0j23I/ZWfCIHlIoeHB2BJutvEtALjmfW5EW
2mJOQ1jfjtz+OpNLFG85Xh64fLSp6li5YV4oCiGTgTvIPDD1DRjQoc7iwfcXnc0d
72OqRVO/TRJKrr3tTs/bkTCwAYDadd5m8APrBf8l4gkXXnGl/d6PP2dHyAV427Ok
cQQVh6D5O839byhZZchOzEPS53nTh2CqO+41yloTraG2U6KiuWJQ1yte+gvPdOWW
f6658ICGMApt1rCT4DccNT0FfR0wUDSWZhF+kPpbXsrKMnn7phAEEwHja8kicUet
lq5ooRlGbXBEE0Coie2PhpmQImyuUUcUpRpvaw/SwJu9dF7DCw6ipy0xDHNTAWYA
gmdJ1RMledWHfOhSaiRhLRxzk15h32cQSqCUL326RCy9y0PpIgdyBp2+TgP0vMCO
KDMLt+Dhrw/YOEViuk1NMfnMos1gRQizufPzayK6ymuLkghib6jw7ADObGyOVhGJ
ZZaj0baB8ebXbnSFoAkB/P3xJdccUgQKzTt1rIAgK9v1OJhGA3PARp15YDGiRhY5
Y+yeXeGKWNdf4kuPXdIwYqmUIdY6idYqYPFWceinivujNuSBbNmjDPcVCTVMQQWz
TnLsO9FiWmXaq6EnAeAWM9Z861thLl8/9d0AYUX627dO15xXAuB6mtgCJl3wbrMW
SoyNZmAW2lt6wEb++u0NQP9//8uQyMSEk3iMlcHnYRENBFoKp0io0CdNh4aWcXAk
QTRMpAIqY+JDQiUnMxuWxba7Lffp7nPS8sBLgbXfCSli1W4GQAsILNxiMMu6lbjz
ibBNpXCQo5+bY7cttC4+Q6TG299q/X+I1pO6ohWlNpC3+Y0jm4FNGVyim37bIkPo
Xtmbcv13JKksK/ZVkgFF/QrufkPxbcsRz8RPfFl/Xa4/SexRE5y2DEfQWapFTXsv
LA6NSaW1oNiWC8mgdQbBGU2jdPu8nNKp5CKnjQVcwIhAo8u5BE2VxpCKnvvkgvFo
Pp//FaUjo45L1xEsLUTpBUDMyV0fyGVtxtBONBAtb+TR9L7hirA3j2rtYYur1n2t
gPhtTe/aQ6tMHFicnyolxPpUSHptzqZ2dbYzqvRR+YqrToaOngOrRsXh7vOHilkI
MhFVg45dh18xIOifDoMcQk3uJIA/+mmebiutcfF+pqMSirkCdfCWXbBC3Zh6v74y
/e66/QscquJEyjfvOIw6F3VG6TecAvuA8uSljwxp4+KY2D+jylhK2pdrzGcfarLA
POEdIEBoVXK3CEwHSweCoEfSq8zFqigzAbTfUwUI5amIYY0agMxCpTJujGQlJb0I
qnM5A6QmmUsIUbTuLkOBzy9R7p0swM3FnnzD+cRSCQ4mBeBDiIf191biA87jUb24
9mn5bwpnPVgxfRBO7i0VSL7SzIPQaM+jHgRynYIsaPhiz18zrj+mBGrFPwI/G15v
fpqnEzo/lAKw2vbhH80SP3Ic4SX6B33wRIOyVf5jyao1+qxeqUkCzhEBWuxnWZQS
mc7JTtGfnpBkHMll34gDtUkSCUn/CDO5Z8YvCAA/ta+rw0nv7cdoGAh4maTqc3hK
qqFlEvdOBX7wJ0eET6AEXzj4TDJnDjRHSYaUlC9zdLeQo5quOU+5SyEvkswT40NP
QfGY93R5MqOwmVhPWPwuX3/Q+Zrd5ifqVxlPN461CiN2RpiEzuGuBEeg2OTuEOk3
HSTmOOv4WRt4Y1A3STEpc3XNUC1lLlakxvb+a8xqZo54mugBKbs640fT528JKczt
7s2P5b0AiHf1TZFndC2C57DExfbtgw6/+FyTDcOFrSEYysYRZGA/v6jJwMXX2HgQ
aiWrxbI/yeIIyJzpMomYMIw091VAY2zYlYV/LFM/ho8pMNwrKbQYuCnRRnYk5prS
FdLAytD8TDAvhUxWo+fwZyF6dQe5DR64wjF+2XsqcwbmQXyUrcZIVbE5a2SNlOpj
1wZmrN366YAvt0Bp6G1G0mjACaIeox5mwfxMHV6ZDpKnmtCzc7O1bXnS6vmo2AjN
uC6Q1zMGsQFAMz3YaXSvhVYP002xyaNQpgZzBhRKS9Ae9cJu5ElcNmoieYzhLkTP
feFP8pMy9eSFFEZCX/tWpPrghzH5+3FpIiQwsHBRvXEpNm5wdqDkQF6rUAtJ0Vn5
TzFBXTqIN7GmIYQ+xJpzAK2hE16c3W9a79n36MMqU6kibg3WB1mxFSyV6Fc6olJ+
qwR6+on8P0ebV0Uqk+SGJD1LAC5mK9g5yyg9xSVgxKbjQiSx+bp3ka2EaPnTl3Yb
5SV4sVRYpx8KKXSotPi9CsiTfute2rUKJ19AXPp9pYmzpICbRaJHGWPwMDracxvZ
3RBPIdny20t5O6VkSBAO1hKdpLrmpQT+5EMsltlueF9OZgLmbBlr0YfIG+fAVbBh
T9dw+BplaG7kgdfSALYfiwqZfrBRp4l6SzTMV0DEJGmzIlj4KZvEEs1Qyh3Vq7KF
X1ZlBaFXkBksRvau2S1p2NKQFMtWUMMlouJRd9Kc5ymEZMi+mnaeybNL/6tqfZ47
M6f+/8PpGUMHoo4RHHZ7ogEjSxRu3CrMpUc7VvavLbvAtEE92+hJ0SkeOlfeCVMx
S3zVq7ddtemjeQVhaq3voPbPkusMDcIS5OIEK/AQGTarX8SYLn5710olUo/wZrDJ
7VbYP9KZcysuDMJUwYGgKi7hk8iCQyplD3Qo/aEG/5o5s4J1u0wbSFIlG0x0dwPo
S9cWu9XZku6ReGvLoTx1Nh2u0Pv9bCGy+dguWT73UeEFPlkYFaGB3pWtyOEitO65
l5sUBqVgx2H3tyP4FArhUA8jUZviOYnnZkjR09liN5qGPIpJoM51KWZVsr4Xs7gT
D33zBaXD11iZzeiuxcUk3Zv1Nq2MupB6BtMPLO+zfd9FSYOpTt6H6MkLMfhzGIf+
rEFkNqfbK0PXV4/hs1sT4LSqVcgkL3YXpgzHj0EoM1tJha8ulaV8N1L+aKt1Cf1q
Qzs5LNyJ/Qc0bDeFbFaV6WXkAaiMpz4GqdKIRVXIlnPjXDJFldjIvTqSmpnxM6Ht
O9b9bn4DmY02JznbKQu8neAZm6WIuU6+PNqPRDuXUI0Q9DP7ha5UR+nKmau1jryS
o71KJrWxYnpcdJEL9U7F0BiHfDTDXU+AJ2Bq2ve/MJoMJ8olG1fNstwlksP/zrxK
rgtXWPsYX292jbIlqbqUtOogtBcuMd2enMAxT69rLNWJR0xW8lKioMF07ilOEdnn
vbylfxAPsanFuweiZ+HlV+dMko9gnFHkAKCZnhj6EFQeHzNQOj259uFwMlL96cpQ
7x8kqbGa6FYYGEPQiLyvYyZjjWxkn6oobstO0vqvEkv1el8F3K6vwOSs+oBv9Yes
Q1MpEf/kyAlw3qWubtnnGoJ7lvaQUz33wggxWqG7gepGQPjwBj2qJ7zFwk9OJMrv
tLIX0iB8qEUdT8+3S3nkDUbZV+TClsu475lhTWLqpxZvkhruHEXDqO5KuAdEN8bi
z+zPRUMP2a9pUSCN5wsZkjHW9ECeOdvwUhf8ktTCw8FukHKwOc2d/HUga47di9ll
RWlPy0D2ahccub7FaR8bLk56LjHW7JN7aST0Ev9p8xaDkT7tVOAjfU7UnFbNvPYk
RkhcoQkytXIocUnLs5nxh17EWPMw0Vb7qOhlG0ecmpXpNiaUAmGinfrkJdvxbNv9
uQT+P+oBvDGaMNPxUmlwAiwt6ZErWGAJfuPdta2aQwzjAYTM54xEFdynAoSiL0mp
Kf8OQe3PhNZM+sfSFhBAWTgzRe3L7C1EAb8LQUirEHSXrhpgrhPxcXgJOgnAuRqf
dSxmmlQMHNnl5zl6fCGObFbpUmiGCNdbGmxNUUqOFu1l6pp6lVDW3YiqzpYo1UYC
MVUMC5QWZ/RKjXGlBApkOXf+kNciZaS0MxzOBhFvFYD2oAYqc6GfsXkefXex+8tC
o8H9a/Hy3zZJMQ0sfyyg0Od1O0vAWNSnesjm6FAMSzxNdLxQIp8V6AqiCw7V9c1p
W5apxtBzE5Pa9Tz3/1CxNvb0sKZS3QowlTgDmz7gBKMtmP8c4g5NJoQds2Ew3/B2
OWV1Y96tsn7qOCfsB2r0K/JJoR1fz0hBUf+3lZZ41wZETpBFtSXEiqF2aJ2yUpOw
op6LZuWxSB3s4GsDhEAHaT/af5hNBcqLZ7eF4JEHeQ0ZqzE+0ZuJGuW6dUS6HgAC
Q+aLgwogo0pWiW5I+u6Ih8OX+421LPurwXnyoHqLW7cRNG49mGteSL4DVigM35ki
z4L3qOPHNyZab311Aba5YllIOlKxvCREAN2c53xvjqChMAw2qYnQHSmmtdRvWAxw
c+apcAfvl0F8+35uNThBtqml4NcQ0PhotjZ5O+UCiTrlCS0a/KLPNbx6Z5WJ3S6/
qhh7hNv3uMRpuScEitptEEm96LfbRTEE+DxkoSqZzbaICyTu4PMIV9tZKnAjLRwl
lBf3gC2KOfqLgjdpnE85jSUn6BVcNV5/skMULZkqB+bXKA8zRU/9Y0TopeQ7MST4
QGssxUV8MXCsrV2KsffGEC9Y7HTujjS8W4K4qs/ogcxYN8aD5hif56vaDT+G2+/i
HMzUrnZv9+4Co7AP17jfsE6UDuWAoncPHOHVw/Nqy8o1QHhI1PwyQMriD3qxLVpp
vvMkRoK3K1GAExn/wZ0xebTgdTfkbIOJVEr4Z43x4MkMFUyzBgsvRBgVUzquXW3l
4qB+56JVq5eRKB76b7iETK2mX48IJQB9UCbWS5RZh+yeXGhQKPpp8YunmPAsAD5j
W5Al64gVGcNLs5BAwTi1eCSM0QwmzzdsmSulXlxgvfha4/62mf63fP7VO+hzAUik
o6uXrJBiSlrdUY5d4wWV5a4haFFChf8OAUwHVCoGYAyllq8iG0IEuFEWmxOk+KMD
ddVXYCsZlPCg2m339dnXXViGeCtA2EmDBqT83jWc6QPT4fbSG6zR+fwDXWtt7WRj
evInT6IyEE9KHlv2hhlaw0RBFygb8LHsY7/NHSCsYatnZgTce1lzyhn9iwS2X5iB
yq0rMysG3f1478MfqmFGKSEda26EYldedTBQUqpsjGa4fbLNoEr4yVGkdM0YxB34
ZIHaPb5vMEf9SYxzytyl+UL+G2bCa6QQMfcE0tueCT7wmCmu5WE/Bax2+ch0/Auw
fU3dyGvu1pOAMJUfhLM5FV0ILFaCfRzdl9RzB9aXrqC46fczyoeLMFFNpb6cDp2J
pdGa+/ErNjWHEgnRQnw2g66x22ovtDErDg8yXR81Y4H49idFzf5JyfQPBsU0ftiW
NuvETXM/Sn0Rgh6FJI+hetUlzZ56kSvlD3QyGewUzsqHGOAZQNTZyrPnKre3O7Tc
kzNxmmAAOoUHj83WM+UjrF46e4bolH7dkgF+adTSXYbtRWhTB/4Wo0q00lL5VXF/
YhVyRC3jwlxJxWvyb2yaxj2lFjaW68tpNCEzxp7P/Z10mtVe72VGYIAWR8/B0wFm
MxVh5KnLLVVAJkKiqW8/sTp5c/qpUsNurMiu1pz+mKsWqDzGo8edMT5BoegPUlY8
bvU5j2CxxVUORO5ALtzd2Xd44uLTv2OVcWieXaTOSo82BjL0+WhpCJiodCaWldCr
X3Rd4v4RKIeXKA76pV0+dQoDdFHBd48FLZd169j+PSDA73vrZGeuVekoYH1Fto3C
nc1pstG9XJGAKp63HQfqnRoBNyR183S1gEdxgY1zfPN8OOgtTls8a2AzAbDZaJcE
x5aYeojOWyRW1qpjV/0WmH/ZvaYS8TknFpLSfThT8a6y5UBCv+kNzcH98W0zv5Nx
gjuoLGD4+pSm5ZRaDCGgadr4vy7YbRHAMZheTA0UuWeLpnUHfATYexD5JcqKATuj
vELgUhYrVzl9cWaYoutxpzMO7eeAvBK7TRH9uTIFOTlpoCr0U0exmlM8O7rzgP2v
IL4cMXtKX/CXxCV4zbMZhObN9Q/MtcbrC3XOUp9KGaAB4kFvDTlyt6tSjPyMLa57
Owwsv/eLO0v4J21K57w0K1FazTDx+3ThgjgFhnVQpLuShXG5fyHooamVepO9eL04
ZTrXTIUb7SZJMr/uoATbVmIzio6rAqQbVouWzrtHycDryDsZBTEM9JFkiA9kIHZF
Rr0rL6a2JIi2bkzBnSMUsnblk7sk/LPRNuih+Ab3AIc+rJJncgAmbo/jvTc+TYsR
+naTlo6M1bN7w7UImqSpFCzCZvSQVhZWJwzMg5O5hna7h6idmZK8F46kc/8DG5ZN
dWTgZWLilxpHZEOrWV8jQnD4iipRr5HTfRc5q1jBPCusn3A52mENT9gcBUxpYqml
aytRE+L2lOoHs38ILzPeMU/HYFWsGPILknQ/S0cDp4uaStKi1RXJqKsX6xjafK3X
0KiH70PhmAIKAskvAPymswnlRnwKE/v42I0XvnxhUXEeRdfeG+itTrXmKTyGFPrn
QlABm+M4J30blfKOrkWpSrW7lQHfnr8uSqvioB1it5C7yI7RkkbK9AoewsREm46q
8hjFqKosUF1j4otpic25OOZ6KVQAM4NRPqvmVWLWR9MfAaMOs70/SQ66xIUsphw1
1yrJd4YV2RtIn0yuIgf2BWH2yNi4TY3Y8Epi+Kn+D/oKKF4/C2hHKjxWPjS7V/QY
F9tnY7G/UNs+9vqCWWkgGnc8n0HV5VrKlUfmQ3hnyDSalQcuoLBDJCU6tgzV+0Q4
5LpxZ9Jq6Hevfp5HuJYVdcqTixdBkTYgli8clDADJeDVRaBkCNMVnfxJ2mtbN+Dv
UgKhOrGMHK77eB4E/frlLfsgta2YW1sTWvnpK7mvMQNpCdLiQN6zzY3C8rRuwHsj
cPb9w9iRminOiAZijueU92peyq8OmqyZGQnrbGHeByQovMgll34DInFQHUXSS2ih
kYG193Vn6KPR3Pms15jbbOWBlHX4XGC0SL5AROmmbeThuHGpahcmLHHEAYDGLNxk
ObkqeXOTbgSQarLUsooLyMNogsuexT3nUp97NX0qMw4JgCUs6M1+vbOSnoAiLEC3
AtkDvTQZdmai8nCmbR4a5WYo/q0DIVJqPtkWmiP3A7PS2zo7OGdykc+ZQmgIoTvv
c7eJli8rPBcw6JtOzRo3xJBBtMjTkuRe3G0aggHPUkY9SDgpF5C1Ini6P6A432VW
sFzeLdcKQTrnzxH1cCvIXiqNjeyck3ORScBm9eKOMHQ9CrgRC2tfDyltpm13q7VY
V3HHDaOoYeY44DDZ1RLSK23rCge5wDg5StKVI+vfNPV5ZfS+J2kEzVjX6XqcBu/6
yZag8toGbBp0Ffw4l+//8ER0tGHu3Z0CgxJEFU6bOjO43acx+bMUW8DTwi7CS1/X
unSX7m4pNL1LoC2uFS4JoIknHcnGUbch0Z/GVX0Pa6WXS5a5POF+n+VR5ip3rDXi
jqxb4jXEeP2bmuqbW2Bxnr4OSdHMhBkECGy5woV0btwSNqCFsbajbUViMqL8xye4
A1T4GCBUYZoLRfPxtczaiBFdGD9U82YMDVFcRL0+gl+/SjlFjXg0mMc0QGSn1TXG
eNRRq/a8/AknzeEy22N0Jo+UDQO3PhMe9qcV911yeqFQqzdXL1K2q9x9rCEkav6u
Lrb3y++m7ADDt9MOFaqHERv0LAjQBTF3jfF6HU53kdfOu9K6pq+8U3JEvBxaLXw4
on5mxv6fTy99TccJjLPURN2WHsz1CBHwgRMyf5gIaF53yNNvsvE3q+tdFNN/cpfn
Pz1OZBeTEpOwrmS8m1KD2eyuIawhOcrdHnHmXhZRzd4CkdchsYLZGKG6mjLG/jgH
zGGyLTicmEwwzBrT/OGmPIHDSHhJ3qTaJAojYIWPtyiMUXsnPqQIUpO1hwLcjhyN
BH9KhRF0rXn5cb8WDeKpa8b+o+NA8I8iLvlL5LdUYRCxqEf5s4cpnTE9bYN6eNUq
cvUlEZ8VUQdJw+6dkpcuYVsIPgeCi+SM1lfOmZa2koHseoCRXGYPhWrAdmm7QswG
h15Irk2y0zMytyp5W+iiuRsrMdI3RlzSwb4/sb97bvQf0CBWzq3R5bt6YX2Wnd7S
X2XbTSKbVsoqEFaChwY5IKK0MfCiOHg6DYQpGXyniAY9HRjBl8HJ3ULw0KTQXO5Z
ENcK6j2avSKGvZQvrcvDLYT/E7/i2KfBSvEtyL6lgTJwffKK4QrCFzYq9Y2E61K/
dx9+A7A5gRYXSElyRJ04PpP9GiIokOwhUJIgBgregEW3v5+NkmkSOlKI6ziqjY4O
7+vSGraQSFcAUiPe6PJKH88conSVsxCRFc9BpFeABHqHv2+QyiqBtvNJyFkFrKYw
zbse93r4UUFc3Ej1zpuRMZGfNRjeHbdnW8ekxW+wI+MxGYcppCSuKnTpPptvk8J0
LBtb7SgVbrfJeJWIq0nkbN9ONeNkG5u5OduknZwwntPrXmRuSEmKw4Fle4vrEUum
zhudiJB0iMPhbu96SB0o88afOfFd2QyjTV4yopW+SM2C1gpMIEMgR0zt0E5yVD7l
jqYh0i4QlVK4mgY3dC/S1i+PO2kOyUIzcHxotdobLnCurtSlFSZVmoRePRodO7TK
/4MhPGOsHn6VqkVCY2YWJ4QZh5pTxtb5z7kNWPAXyjqMkzQib5+tHqHk/NmB//oA
wGT28LKkw6AZV1Tdnnk2ksrnU4X1gXEYBU1sPUwy78gC+zB2ogv0KxzNhtFPfQ1e
3okTZf2T/6wLiEn2Q4XB9IhBPdDFFAlTPExilrJJyEHjTk7RSb+mQzf2B1dvSzXC
w90O2X7ptU8xH+m+oEt83WmZAr71MB2QfBqZWiwGIvYBqFWK+xJnTJac2KUIG6Ho
sgO4SJ8w3iBZIVKzEiZ4d4Tv7J1yVzUjWrVvuH6dJ4sy2MlS9gE76nz9N3Rog8rT
0fBGXd95GyGpcvAfyMBsLgQvEO1FwL98k3Wa8z1xsViospkkCK8RMinaBcuYp/J3
/bzU0i836waZRCZVAjBHRJ5V6kAD/vbcZA/YJFAsx0eHqye3lMpN/RYpb6tMGO6r
bhJakUx+4IWmsLIom0Ivx00itlhC3U/yM3oZm1dXmdUFcPuLrzawo4txgNayOwQs
446GAItcNNv7GEPc9CCT7ajAkEy56dVQQVHV6Fo/tzZiPXFG8Wtp1N+WW0h2y+6E
mXI/E3gHxbT1RRj01P7m2ynSwddmItmEA1YtnEPY9ojjLb8SxAAcB7Y3F2Z7wW3r
OAPBolZsd/riJuifCb1eSekZTI8ECbOVBWqf64AsWqjaZXD0dEcFvG0mgcEOpjd8
G5cvSGFKsS/sfVSsuLW2ZRl/ErTlQpKX1Jg21dFZ+I//449PMgrGvW7ESOpuZ5Pz
ZcSXbGgVTKW5Xzan44LBjt31oQqBZFdFamNb50kvSZCW8OpLwx0t+Taw9YTRwdmY
wArEN5MAMuH4K4P2gWEkpRBZnHVlZaoRH8TZueOLr0eoPFeFyv0MUYLZXP4TTNwX
gys2AysXCoV6M5jgZ6OXco9XdRssoGA5dpi+xUTtNqnOKn2LIwbPG8cgv3+sAuBl
wY50z91Ye9bOEjYAoQ4GxBJJcESAh7774DOagOxgsuxHY7K3/C+kJJ98U5FtCr50
BqXK+cP5zYtgF6A+sbH2zWppB+9yjb3U+tr3Q8vM4Qx1zlL0bR6Eipl9fdwzzQvX
2ORlaQ+UI3xlpyScE0t45d4tXjYh6W3Vtk60ziKga2CQhAoT66MBfAUre6nkzJiK
0ZgtvSuJVAHVP5j1nCq8842vYDnmBrAT/HOGV0GHwuF8YzQg8rjGzvEC2oT8yT92
0UXPqJnlzzzfJ5L6YaVMW4tD+elgnrXF5qGUOBeC1l4HBWXmQ//jlrJIF4G6aywK
gpHRAA7rs3lnu+XSRos9uKooN5NXxOi4BCXwv0KTMmXc2tPZxDd75p57bYyokqbC
GdpJrUDwllsfuw3z0Utj6QVoiTbK6Ow4DyIKSUpyPPMbwEnEmele04lGuWLHCFjQ
kzkKiyqikOfjjm8u71AiBxD42RngBo8b06b47Hk15LtkBg0JHZ+D7mGJINBxQ/Ov
87+8zHgF6XjtBFfRYMhzVNUbx1T4TmK1J8hhHyoGv8X3HLxVNK73FlAEvk3GbiTH
90GijGGMsml1iu0+zPtfDaaG/FqEpnGEvuJW9XKbHtTChCw9vPO6kC3NQpmx9CiA
rz997Xz9pRG2VEGyB5U4eXmMgMx9dmySQ/rjw7TDOMKAxgv/lCYap0zsatVcZwSh
05HwJBLzF4RddfVYy6wus6wBn1CBv3X7EWWynh57OQmXAXQcrYLZRVOq/VQZZOdb
XnvkFnMHvyZ0ztQAhrT68KCmOfv8keANnqxpx0HAuvIdDc8BfViOiQ9ZBQSkRw81
/YwfHcFPGIlvOFSYyIoJixYDoc031Y+OYMli0JqeYal4eRBS6/iZH/pIMbA9sLTK
gzr4dn6xly+rAm5Qp+ODSYgWlzJ3RG8g6X59UVJdqJtn4xBlSHbFKC49DYtzDLCb
uSufCGmHv1ecWomAtQVSrplT7nAJp+yiEN1TCHCFDgpjrJuEr9hP+yMLwokZKPff
lTLGF7HQ7o5NwU43thAx9Rx2e5J9hz5cPbojjJphP4xkfG4+6d6GVWqXwi+NoHDE
8hph9rWEc/zvMBlEsO507/g/2V8g5LvWQ+r5zUzXzcITobxpDCRgaASyR9F3YGve
yUaARPgLaDoaFw3r7P8Diyz2LgazsRijJfwnHHK/01DJRF1BLN40OzGwx0XUxP2D
e2E/2zrkv1yWBMbi5QTlKjoiaTExwmXVo3GarAfJEigElV6Bs2WNRTEkXJT8SHhp
VOGAb2D2bzR0Y9cPtK9+HoZCPg2ytcqhprSzI/26298MAoQNySNa0neQ5NmwAQSW
mKrvIG8wY09++i7e+LXrYW7gch2InIczuqqyx+98V5w9/Hj4eHeikVOup6q5xpQ+
G6mVD1P7v9hkUjlJ/tQp5QhTBhvNn7EDmO6iSvaoZoPup2TUbyfUf4LehSrjcvKw
P13/St0Tq35AEzcwwiwOjZBC3T+vtaIc8+KUPWlNceFgXpdRplWtxKmol32f3lkT
DZfr2/hE3vlFp+EvIB98zua+7Om0gmRCBh+/qB2NSY/5/SZrv3uTIl2hcAh2v8we
1pQCh/xkesqIiNaUZiK3oBFb92An8vIrIi7XzKPZ5tEJ0YBM6DnJnxaEtwQZqerF
dNfvqr52ReM7HtxOvdi5PZ1fbnEHnpNx8vSjIVmr4lMf+YAQByIPGGmw1TZu1b7h
6AUaZlNwKeq+UEfDPPPUycQ1AWn+5REhRaBy4TWWeVqP1S9JKYcSbdm0TeVikp1l
76lfs9ozgDe1p+vz6nhDondQOH1T/89w9uPr3tKdN4pRqFKjVZYnOf8IlzMyWs5i
fp+M87RbNzwj0dUqWyMJLiDSUXIIHRgNG+Ybsdf8Tl7RKRWgrALfTtF45QSaN8VH
wQuTi2hUnsbao/W3tKpLqqOJWtBu3QNSg8jNYlVqkCN/RbSSuyY4H/HM8gVn6hya
sfoH4jIsKO/bGld7ZLD5GjhQGhxoT+zk5+VqsW1TYMF5Mhmdse/nLGyRjgXbRid2
YZRd2qdqdvneKUQ+75xafSuYJxupnVpJle1R5Y9LMxcB49lA5CkuVA9B/W0HMQGG
6oRT1sJFAK4naFbyWGs5WOso5AxJahXLl6x00ZyzyyJT7DKXAh+jHfaCpAKlr8dZ
/pscsfgoZNBNN75SxunGwwjgL6tdzxwQhl2mZw8ADnoPbcdMbJJdDnFImI1rPXxC
CFzQcnUlqs/RxvQ+H/MjAe8Dbvm0C9u1GXaVrXx8GWl6zMTBy3xnRs/7K3PQrWev
Kmu8NgfrIye6DQVLUgEVUTAETs+CeeU4XBqyHCR1W0ia4D12MQxDyHrB9ZfNNF1b
O/ai4Lz7jPTVXGXui/E/Hvv+iMu2k5c6M5J35IF44PFWKpn7uOr3eUaAvs97cmgF
NopJ2eKcbzzmZpqVJMAvqYKUt43/mBqcP9Sx+XurpeqK1fus9Gi4D9Mt9KcXl4L1
PG/Eb+hc58TUBvglBhpAVEkyzqxr4w/CNdVZ05h5zn3ATlUlz9iaOkaZO7Onhflc
pL2JcPoWGFsb7F4MzOAceTPQfTEq5RWop8ltmJv/HRMOKwBOHz1vVEQ3EpGo692y
klUfpTdHZzC8CGr6tFP1PFvG6MrfWm/NdyJnYPakrCAzv8uW+WhXpmM8oxar8rlE
9T02/kokaTU+KFiBbd37a3zk6hU8R7ysLx2BWtpYDmWPCV3UBo6mjUyv2HZty9UB
UZBt1EOplMv/aYeYB496cc6mIKWGPxz5ypIzK9pLd0VQaMNFJHvzuwIuZu69r1Mq
apsi26ulRCz9TQvAeSxkKnMXW2AwnTHNAzwti8twHyrWGvPohCiMQxLXqNr1kdkk
iEeIuGjVqkW3YlENn/Ea+2zrdeYphRveS3s7jncU4mWs9QcPhsLsGtxFrSxQ6pgl
ANsNPITEpGv/uSTkgTbOrSRDy+yy+lpKG3z6ke1S5B4efZmml9mBqtud4cbqUlLT
nIjCZs0hPkoR7+aGazh9hc3R/tj1hA0Ph4gx0L5PCeDGihaQc8L+7C0PDVs3FM7p
oFrqyHpJ922aEWk6YjR9QUakJxAT89xGpxEOQtEUGAKRDoLIZF16GP1wQBpBYCK6
18l9oYfULk10vMHMhYRu7RI/z+RLexGvGGuFnay3KOZMUwChUynB/+2ehzE6peMQ
Wcj9KQ8do/65YieyWbEnt204MxbAzrCv7NzriBNbL5uX0y0tNecS7nrO+Sxa/Lt8
yT5w6sVlU3KKU4iROfda7Lj2lS2/UUmT+edDiHqMONI+Cu/cjjk73c/BftvMm7fY
akRtuLXU0GIWLxu1gX/9gC2u7gpLNy1rPzQkzmPpocF6faoOI9t/ypN9BdJPEV/1
eoJiP28gWbAqf/jxDQ7hqIJbBlQdX1i4mksJha1oFI7jKxHMq9G5Grh3ccju0xed
kHxinIXN+PjfJmv2zsjIV1rBJI0AjMp1QwrLm1b1cL3JIqEcJGA82K00tQ5RBglk
CLSo5ZtWbWht9Q7SpdSroUhurW9yJqneuHt7UXglip8Dvh8ZCoAiq/EgRDLyejCp
ANks1VH5xZ7BwhLyZ3jTiZyQHxnov0Z3NNEXblR1uVaOAGIUl0+RWltheIIDGPxo
vOVLBWo81xKK91k7O87mwTRzbWK/oUV9k3JPZdKLOl9pPX6Kqykj9PzA9kJIBBEo
Y6i8pWK+fjoz7x+/MKEX9dLk3WCLdNZz+ZayUSgFbWxocrGDVxCP2vG5n5xjT8GY
OpY+BdmPZw4EBW6EyJop2IUt7qGTAEFiY59LiGOiksk6WHtzQTWb41TecdNN20nh
qtBSkokrytQPjgWS6M377yg8vd18uvAXqaCTTSzPu0HUcaditjuUPm0BfEopcuGt
t9qKl+33FRYmFlU1KWo5QnAi/hfygWzSzy3/+ZINFWLtNrp1jI2sJurnHbgKL77X
JLql8wr5R4xtPGMFeA/dXJimbcY3zWnTx7hmCKxnfds/LZJtgQo/30cVihtMQd8v
+20/IQRggBllbMGY/I62ucIkPMR5rVQ/WzbU6wIekooo25uo5D4f5I1TC6+izdPe
ugoanYkdTkA1PUlBqABeM4a02BOLAkyec1Jr9ZQzd5dlh3aatFgvmmzebun/HgHR
6owSJ/XVKg9xHMBDFjoisvaYuJsKXyUezXSkRylX6gDG/gPWD6rSF7AnxqjHaTo5
tINprpLo5cqTtmczJdcLqtyCtq3Yw8S4k7aacxcol4W+0WStUWEgqbhbzWr8kt/3
o8Lf4eGhmrlsyVW6n9snG1wyPaE0XMrRX2t5pdukuNwoMIfp6cM79bxWkp0JYvUh
aG/xBgWN9A3Q+mZJmKK/vb+wajlYwUQeppOvsxVzDL1YOvx7xS/n0yOR77EtiyzO
fSOLeMQFJWP9uDXUG6l3MeqqDjagQTHGCbYzam5C6K8Sc+lEQ439WJE16vxVPMZ4
oVVmPkjh5vGvjXPDtGV4vrOOcpTbPDYiQ6b72NkcW55BDB2Tje1e65v6Asp00Beh
FofC/ODFMUVamqNDp6Qk1rJgC5z0tkl3DzHJVCoN976LG7BqU0oh8VXZZhWBKX0P
XGVnEicZes0oTctleUbNMTpDgEvIT35yLMoqL8MII7kv+k2hqtI6PEpsLWHs9EfY
0qQLWnB9uPBCButcy50Lr2Lq/aXVsf9k1qaSdW00IHU7ookmCt5U9F90sNaLpKiv
B/xr/oY5Y0YRb0xd2s6jtEDVE5sdQ7aBt8sVcoIaUxp53kACZGRviDeHCpbSZIi3
1GdP5esQO6PbDyyaRPsDVl6X30J3CEeTj47SPY4p8kEF0PphAqMc9wbl9rS9lhck
bd4enngc1Z5wOPlceD/2J6WnVS2SFIzmULYS6othk1yY6JSKIzlF9X/ZC2ur2+fn
C2Q/Ov7OzsquHJoXQ9Oj3qxuyD+PxjuqteMflw/+6uqEzh585OX7Yyg716n0FK3O
xSCQfhyrrAMou+f71XAaw+mB5yr8SgD1l5Kd6iKykQ+1bCLEG/eZCbR3dXxDLJlg
o15+O3M4BlANbmaD5fSaldN3coyslmT12tD+Memd+HMNkQBImKiO7ENzViLkXWX3
pSYc0Xw7SUb9in8xnSWbXwUqhE+HjeG60LJkCmgdhWPrRhFW3Lca0R39paGvFceg
fbxEamGUnx/apuOBr1OSTzliDwb5zpQvEJARVlc85tPQ7gPZoU/FMK0i3/2HaHP+
3RaJ1J8cqLC/JNsCXQltIFjXex3nTigEJpBt+n3IEcvGLemJufxAhnKq8fNmXHep
1Sholj0An0WahuKuewGZKeSLFI2KtY0cAFdg5P7gRwzyJcAcROLB9CtiR8gquXmU
fxMUCw3SRVquVnFudqHaUZGMy+R3qSnCoeW1lnqaLZcH3NvgGtnGVV2nxpyTj2wa
B5vnj+86B5LZ8db+F5HcbJBGXsT1fLBlxiv2XHN+8WNcWPD6KfVi/taIxG2QGtCm
OMfBA/iOCvzZFlXN1MIxoHbJcPE3aYhxYOLP/HlmpoRvlNZ/sAzIgOsOAmFIQWRr
+B3hXYXNR69oy2InYm3uXk2weNyw5qpwnc2OmbvTFIwMdXwOKDHOvus/WFJva8xw
SZRHO2gYdYirLZTbjSWkVuP7LYFKQjG1RwQwi3UktJS0xuJjHh5iOb3NS2d69eEo
2oinoNDnL+rYlHIBZ8YvRlSylD5SD+q4Ie8p2JhwJsTe6mugHZj0YNucyP8FSjwM
isN9GQ4apaZ0ZvjWV2AxPygr/WEhmh0tQ2MJ8aPc3pwf2Fi528q9sGQF5pyYorCo
sUhGuTTfOo1zsmgQgCfWze5oKeBpYptx6mhB5pkKwyUh1sCdP9y1d5jdP0LiIesq
b1TmlEx6vg4nVRVzmJ/383tZ2XIocbCnHPaXUnl6iGc2fYl+9qWmIm13ke4eCnUO
Y1lQooS11ZCBl7whUnfaCeNw0t7bwK0kep/dunMZHViNxcLAt37Eg0NV9C5/56TK
G+0FT56TDGPAqIu0ZhBstUybc5HjlbVlrtf3Mk60Xod1fg5IvxD/f69DI4RwnuZW
RQrQNBxjtRuP18Qtdib9o8XYzIU7KZYM2hsyxYtuYYivrnSLbzLAtKNiqBLIKMve
gWiWKyaGpFQ6hgegAXBhqHG21B9VtcJnuKjp6BCkofOjE+We4EWYycZbzLzN8ojI
JbkU4eKfwlyXmdvrEuyLjl214tfLijGYhIyqEmqHDIP0TkDxSf5EihrkRBFvZ7y5
tnhWyzRNP9OVGuij1L0dEGnPOsmA5ASOXKKFO2pRc8DN2GX/5sukbI+SEAEleP1u
JhEpaYImGp4ch3kIaXgBAYTWi01GsJrlGrU2JiJtOXIn1ppaNxF6PCbUNZaz70fI
FVYqsaYJ/dc4DfeEV43R5qbdJUr3digoFG2077RCzviIbW4Xih2dz2pLQ12l10Me
Mix2orRawhIS82xpZm7hHKqMGORd0BT5UMlCgwmMUa2runArbw6pJY3rCAdgwp4L
BGkKhyFQ3ySnHAzRxeFgeqvLjLnELr4XuAdQMflOaZ2sjm+eTPGHooOMPlk9MCV3
Voij+flpujWDDX06vyisqEzyYCuY87aeU2+w9gw9UF9oESOLxBQO5uAjy7eiREV4
1KPK7VRuhKtUwt6kLsDW/z8k68w04ZtIF78AXSNWA95/uOPs4/P31WcDCBWuXQCE
2sTF4Aj7SUlaji+L9dVopdsi+pjiwJrNn+wyzDikGc8bizEPRwrAGFlwOaJKfgvW
eul0N5D7ykoXzjzvrd+/aRl+UU9NIe0EsAymY112XK/YbCX4wcj7Jizg0/9WN9HP
UBuPQNvmPN1zNLBvb8xP0x5iuKwkf/9SyndbCYCk+1W+yaO4j5YCr2u31AhCj+WW
o+yKS/fgNg/hxJHBPcBtFHT3RlXLBxipDX6phmTPz+cqeYp/6KbNcaB7iKX0U/JV
A+DU1UXNeJSTc85WewaMW3KAqdRqaSTHjtEPoZULfMGl/tql97hmtZEJdGKzVIzH
q/+f8844r6dwk3gw4VHqy3QojhlXMtZZx4eauvx433IW6ZSYQ7LcQ9eswl52/M65
VbK2yTJ0oyzRThh89F8XUZ7QlHTLzGlKxVh8tpt46PBmIoP2WLzxOQLu3OIw4eAJ
iV1AnxkEM84aWDAxfSkUkULN5XbscZi7wWD/wDaHdjH//gF6QtvoWAEF3h1iEsT7
CKBoDw468DZvu1qZpN4X07lql2FxkYedLwqL/YOVCFB7CyEzwRzdtVKatz/wHJ+5
Vu/Ha7CE021RJJyGlU+Goyw8NHPB4XILcN2tPvSYBVGeQqDcpXyGCtNBmBbUY3rN
7rgyi/Aani/03P3EneUUNhgPaVOmAeZ5YmBgQErCT3Rnlrig/Bly95GRjR5fZgQP
0VW3dxDoJ5MZ1MiwfJxvCTGbvpplKPuDmHZqpme9H42V/AxL1FURiUeGvicvIUwS
OTB1Kf3KOPOPbJnAV5ir+kUat/Y+k+Aj+4IxqtajVh+rRItZotHTC2BM8hACqbZw
fK8qV8ZLdDWN53KOZjw4DNcaiIAHACFSFQ2jUCjFMbrF5jsIQX/3DcdJdII1JzcI
Je74Z1FlBqskmfiuBldfn52oBCml8zk9EOTdHmjM8QRRg3EmmepZH4nqD8WWxrkF
I4bGGcZK+MuutMu+ydo0J+bFotfEQEIGFGk31SSGdgUAU6+uF9bmOXJrKdVVPCl6
ZohgO7I5PyxyBq4kCiWJTVq6bOudBOckrtfxAA7On/OQeIAe0Rdh8wrB4h8AK41I
LmG1Cu2+HKMfhZqeRVDtJ//4PmsC3nv5ub+wI5AXa5NBw6TOq9UHItJW7Nd8T9Ue
4Z1StoRei+XFnpYj0M811zTRA3nvJfeL15OwsHK7XIaSqzRxy3jZ1XdOoUz7ZUaj
GvSxvc5ndbF4VwrmHSaikCzTxfY+hitECU7Lt6ix1jDjiGV6S8SyRaxWY1s3jydM
M2zc47fNYKymDw11ZYWfztR9jXKR808EQsBBYfCpMCFS8u0Pl7Hl4hZqx+dpAtDD
FgYz/ZdXrM4k0dgX+GFUa+JGhAwOzwyJ9XlpuA0AgevwR2BAmdC2e9Nx0YeuKV95
+L1UMXHkCvs0KSU9qbd9rXcn9QtfBEbu4dO3rTmKjbqhDtpwUJVSecxmbx6mQ+ur
dnVxnirlD7hsn/qyrfZlQ6+97ZpWIsxEmVnaWJfrsrcDxQdCxcpq3id03bPSGhch
rY44FHzvPCz+DsRgu3kbJJCmCuPHwaA3QifJGoe8QiFqh1xBk5pJtgvMUjM+gZIZ
wYYrmwPElMkfba5G3CbxsQVGvPtFEAeRegj6tMOFSh3ugE95r9OPKWgcf3x0qZel
rdUt082x9jLsUrjl0evc9/0bbbxQqwf2VxbaIiPPgV4lfEXqfkhbFSmUdc7o2ByR
l0D+MH3G3JsLKlQl0q8X5q6ufTGGOsxVP53Sm7fhctnFM60cO6lvNRp/YRlsCy7p
nFBj9pr21ZcvFyGbqnJOY/93UW/6oGVFyj+RsvttYJLN7Icppze8G9+lfv6OqZmO
Rne2u/fWChFedJmyKbWrgW+WNCzEQAWnQhWynbmmzMGMGSZujo0Oq5ji4L2KDetu
aWwlPPPfKdMKbaWtYfO6v783k3fXaoU8nC4LYA/wu285dyQa0nYmr/m47/6Ip3Mo
3GnYtSrIoHfrRpEpiaLv9CbaWUvdzWDb2rksapEm6n4VkttkYZLOgdcquTdS0MbH
D6ekKb+PSHVX/H4BYpWaNtunp+nPDlXDG4nylD2r2LUe0AmcHRuXDfiqD/3Kybit
W9qUg4YCzpHisUdXhvV9A4yCI5y9avwdk2Nhig791kOI0/PXORRHUkjVT17zT1H1
4p/1I3TpYekod1JkdTM7j5RQTSr/2n/o85w+1xdacfaFq5iAttBjdFXk+amguZQb
yXWzmNrfVbv5qceo/r5CzyY3dyJbluJ63TU/Ly+8THMPRgeYyIhOY75v6R4u+YRE
/ca/sUlXx4i8AnjiS7SeMSm5EmwJUhpbHSkMdpZxkrKJNDSq9DvzhfU54CFCt13A
+YdasWAPIuD/AcVwuNSUGOru9DYqb3jK2Y1SBWYcgSW3SwIOKZUwDkqA0w9bMpsa
6OZLjH3QsoaCukCNoXqLhp4T5nUAR74Uq/ugK1tGZlBVP5aOpecCfVyAQ7vhK7zF
FoWcNSWd4it1ZfSXUS1iz9LKNDMug++b2YWVthTLsEo5nQCyTwFpteO0xilVar6o
rNi7Mc8ZhKTV8yZ1oevnhEvCa1xIqe5soihVVsgU+RQTouN0U9xC9rUcA0oEueTD
FTtacdzgorvqCqi6m7sDLBFaFsP1JfTMEnZn+X2VAW3tjHhWuBAOnRyirdYGwVp9
0/kkc4qMNl3zu3EKujwv5PsBcsqZIlwfJpbDwaDIEVUJL4xd9vN+F+tkSmrAWyli
VjXu8PmK+bNKxqQRHkTBr8oKZgmXqRQCW/sje/qhz+6jj9TxML5h0WUwQMpu+I3N
8F4hEqGACYaKD//LLT41LjPSUzhtx9kLWrDIfbc1nrVwgHj2x05jCczBNvTnNwcy
Rw5Bi52CP6Md67QaUQCPXsxOimBYXjcnRpmJ1cS6pTj+dnp1Z/PsparOfiHTDdEW
wilJV81hjpHa9toZNbtK18eUEmkFmlGWUi9HlyY4YtqyDSiPKBoOrE0GNeOyRkEw
paMfVOUzK6unmV/sEMOYlV85mkorrQQv4gagtf+EEdBAo39LXCJZdHG7EVVwDJZ8
bHmnjj6kjEDx5SzZVrdyHR4X7dFjMs7aCw9vDe55a0cN/F/xkoWkCHJIeI++GXnS
5y8UW48Eu3g1iJ+OxELdoP/kGhC+4eFRUigE6hWBei4hnv+f/WYAFr2jx1LZTj9f
Ax1y4rlE9/ancWOF2s35bDhiYKnkYpdo5e/xKsz2yjEyncXm8r4MN5s1OrzrF5SK
5dtbl7lOQTBd/TCbKtoishiYpbZ7ZgAuTYD1avHd1oqYW7GW2XrlU8OTyRs4Dwjc
ytxSff6xRRoVhFBqtLS1fEjAvo0Aj+KYQLB7WTP8fuiIFUtbSCe47DZq+ue98VjW
eWNcVUs5sDYDEgzYFFfrSjOY1+UbYc3WJ7wwQm16nDel8w+MqSCapAEicYdrh4o9
3zSr2wpCismMrbXMLqAmi0hMc9xgReQ86UkvyWHIlNOsjnvi0vttaFvjIz6LjBk4
P5yiLkFqRav4Ke88MVW27WSzVHwPmKDk2vWp+xT1rkUFKHuUWVt2ad7+gutkuvE4
KW9LZ5WpGtLZ2PmY+Iiwh10OZ6TVtcZ3FlDGq36vETW7qt8Kh7sIo9VxBXF8lILe
XBjkETcWPy8YPPBr9oGt9ErjfZgBvyKUUlzECca1r8oIBVSsohO72khbwTbcmDGM
Hs410PMUDUSnyj/Fvw7/v6SYqJMSoOjcgc2CQBkdhleMx3gzz1CY+LmEf4sqvj6H
JNI/OCmnXWEVl9JCShtubBXU/lkzLCTWxwZVwXhfwf6jvJbxx/YSX5wPh4EPheKd
jpAyThze89NaLnkTOEk11RGsf6B550dnWtyDFADY5aAtrUrfWFQED9Ua9dkk8oUZ
Ef8sTFSIOXBrH6c6pqogkTHDtlt/rBJnsAu+d/hNPHWnHLSqoAIki9oAAlgNT5YH
sCHkegkAhJN+yif1f4S0A9XMw9Q66K5Bb5BLG0wvMUYSbpkBhD5KWjs5bizrsy6a
KTGhY6AYMVe+07TwtpQCS3dFV/+dfWgQKYfKsendL9nWmSv6POw4DsAl8t2J/pmk
3mj46P40jlSE/0IVGqEq9jyo4WkhdCtp+9AoXn/fWPa2tWGyIGbDJVBIvnKrCen4
GAsjA1hphu9kCKKBMAw97Nd67RCI/Pppzi9Rgg7KpggSpTioVekFYSSsHGjlH6NT
P4QdgDC3F/flEALMd8YcHiOPQfQqkUKRN0ZPtUxeC4KLOdXY/xMldSLyBFCmeBRF
ApgaLp6C/kZ4r8z0EwblfJiZIRkeTf4xlRFjJfyalF4rogRO1PnQoEksvI1Z3A/D
Mpda4iAUcz8nysZ/59vC8MkCzN5Dis9JvNGCTBxMLAG2BChWefQcoVtjWsqhvdDm
ff0QmBj0XJ9CCQFWKG3oA5GL2sxRaQaglvNeGsXG/7VZ1zXeZxRgPtXQTPW53sdH
9YxZFC+UVuT77f3n6f0UTnYGUXcRHREjw0vgAU+nhZw2x2ftHeJSDG64VGjf4HDS
fJdr9TfQMcyH+Lh9tNQehaTsl+l7nR28t4F9cj256TN9dopcbVn9zKZVFKrX1bxe
gr1A3rKQFMFRkZ9jhhB5RhXVGbBBTSO3MqBYcIWJpZ/NUP1+AC/7/lriRoSJCiyu
XWuPPdF7ppYlLzw/zGMzldGqywwxlOJiY7+sWLzYSYqySbTLl0duksZk+pNTraqz
ehviUHNYulccXsexYQmvjSsW5+rWznrMQR6xywbI4PAHge6v7WQmOtD90ZMMIzPe
BF4HnRedAlgkaE20oWi3RMxbUBPGhZ6yjyZSW3hfTYwmUQzcD3+tuDAo+ZtKsJZd
KcNrjM0LnB206YkCn69Enxl2kLDuu0JkTFN/ssGFb0u7iqhOvUS6y1nJydVdTZuS
dQvZxVaajP+Pyzw//tNv/n+x/36taV/GfemODOp9FNKfw+0qEeo6/nYUsqQNQSr3
kQmXS/m7rGdRwcDeRP0rFsV/K6DORpUIQOUWt0EWPYQUiRnp0fS4gqaKTL4+bctA
4tNwIYHtzpoKs2GX9QtL1augbaueGMhB7uG9BYZHQHfP1YuQtLaj6nis+DHVbwrz
uk7eAQ8vhoY6uSvdcdsn7AF0OsNHmBWvRP1QSD2otU/Zud26Z6jSubNuxZTICPCj
o25qQkByU7QJXE+G6Jh7YSRUCZSsvl6APIhSevsovIhSj2BT+jibxlGyLx19QxKy
tWGhbHvxbtJ1Kfu+PG+Er4KEchYYwikDhs/5y9jvqfxFvUxpZ2wA/5dWEzmbfCq5
FXFDZaqPmLcGv6dkeaZ+3waUKStW7M5iS0pcJKxmXBtgHxB4BjPm+x88XUaMwDFW
dEuPgmLca8RJMxnvgLOUgCDHLSUEmpGLfrkHJv6nx6IpBYqpZQKOoBixAzN+djBh
9LM/Y3mge6PG9CIXL43bw2t1FIepv2+quwozGsP2sLe3MFJWmN3x2r32bSfdleJu
IDa+oxQqAzlCw7d7JoudoXgRixWlHluJYn4lGPxTDFfhye3ZYpUFTR2TQNbbZxWw
dCBzI1o2y28iCzOtaPDq1JVvIq9Fkcg0DAK8DzbpCvaBEk3ZGFDO3DUt8g+BmEvm
JM/k+4vJRAffMxEShntQLHFc90JrTo1FplZugrzAiMJTlYvO8ZO3AGfM4n/D+cu/
xucDzcDH+BdRkGoxOreRF0KR18q1igWk5aVh6MvRAUN6GaXldhf6EbB+TezUPb3m
i2HVDfUFsyhPltDQmjcukIlbXclmSxr7HyrlrxotgTz/mq2BOpagYAnT/IVI/VYo
mWousi1T39A+b/CdT1NwTEF+dwT6nHMItwb4IOb1fyo+hdAo+sbGSt/p5cuxbdCH
x2Pf021/S2du1zv3VyarQ9ZPy9TdvvzxKUxs+sfnrDhCXuV+ovvArOzdApeJ8qgO
80C9sKL1D5JlTmqRvG7ysfGvnwsgjjwevX13LwyUttummbctqVqelkgLxi+Qq8Bh
12syQZMA1MNT0rhZyf2/2mH+gVomsED+u/HUFmYvIwCm2rv81PDnpKOgor35M2xO
3yize3uRpelKTnsJK4MY05vFj9pgfTySWuBIFIQYB0Ws2s2W+2q9WxGJmKgbFQ6w
8zu8WazV/VOmKA/dXYexJNR7U7QpeGtL0YnUv1NZ5vqzgsoKAaGsBkX4YJuHhdH2
t7TADUYxKa8AM4p6KtPIdU/4M3/VgWdS2azaySoacBJaBWFaJIBLMwVzuyDkrtrf
kT39shT73S1N/EvEEyUZyPJebzX2hz1+1idbng0/F/Alf4DBLy9dwCDmqBWwhQKm
WOoE0MfK9IavHh08m7ikvXHObm3goDcpfVkEuoKGM8FrXB6jC9TJ+igSUqgIrGX8
AuZwsfCMNkEffHaKutSgibMqvUEhyZ+/zXDbWz5hnhe0kgB2oI0KjdOSrAYYggk5
tUHmjSTC7TF78FIhhQz9WF/q6N8I11ip7W7nOUX0RYAnVD9h1ZsQgieyMhOd8Chi
RrKfxmqc5polsZ625Yx5+FfhqFCT1a/m4eMeh88e9pSS10klqSItrtCqFvJIxvTt
CeJMnDXFBQFBNxxg+33rVzZuoSzrjKGAyytVHLY9fH3Ke4NYnujK+tCB4Nt+6ivE
Llruie0ovRhO0/nDw5zz+B8V2XMA3ceAjgmqvrzlRqVNCu4fyBMt5WUusILT13cl
CQ0dID32h6u1l9Lo2c7+TglM8mcfZSf4akFcScp+to/1+DkoQTkKp/16ljKhaCSL
GlXaOUsu7YAqIZaLgPL4nqkrzMTMp/EuZKunhBLizG6QvKucxlP0jaeVrHBeJMay
C9t/EhOlllT0yT67V9tDW9ugGt9qECvjNmg/gcihKxNqMHv97+L+T8KmsNoUAD6O
8cKdnbCpUFWn1bomC3col0Wk1XlGOPbiYqYFYiqc8Lh7WCCZF6M4cBba9oJ3sMaS
Ilb2LNtvtVqiyrE0znT/ZZYyi/a93CTWj/yzbNchYE5mbiOXpaw8uP0a40+WM3vu
wBMS6LHJXkupjJkSREbjlw2/1GJmP7COY2BYTCRy/9uGyyEWs1UMGhZi2L8lCbcY
D3/5RZN1gE9tK23AkJVX0FRysZWyBZDWCnYRmpjW11pBRjlB8RIp7JZLGMqj9xuf
Scog8Vp3DYB1sE6VWQA7lHCdHFg9DXNH2La+iVYeRpnIGblF0R9GU3/+TYtCvrbt
HE7itQ8ws91O1hsS4kNTNvvsvOOSPiBuDihRilDm6IwELIewg4K1pIid2kQbwhug
NBsxhM36pHToMXoHWQ0RBkFeFtGanH7PyzqY1bxFebsSihaTddewW+htj2gIlm1j
3pilukBjTpzdF42qrUzZg1hG8qy800hDx7FWzp1bVrV3X0pBSNehOe3kW8/b/RuQ
TBqcXhlMzS73RBly7UiW0As83q1OP7aM2uVgu4ctaQBsHnVtPRTA/i5Lf45HTf0E
QTRCKAwnHlnuMt5sej9Wk1V7HcUekWWLzTIhonDO24tPTpEBiNM86M8VC2eQ5kAQ
upqf2CUanvYFaf34+rcGHiPjD1e6Xbi2db4DbvRNcDLQtP+u278K3LZ82phiYC20
YPw+I6CoCD77vXDvSz98QDvau5N2JBXde1tVuCWCkSGVMg07fV9LwS29QkuhmOUK
tstAmW1iBOwyAJ/RAoAGD0mnnEodBF/qOlXVuExC1BmBzWErPxZ4us1cXDeRXv3W
mXIeSsM+CpfuriQJRP5+FuhT8CClNLjyWrCMB5s0sjvaDwrdBxwOUQ+FhKnL1L30
/r89ZjMxH3Kmv1tRCwG9WSc9cKNLu6fasPJAsq2+x6I1IHvxGZJw2/UZXLnJJOGa
6hLRYE0JTWGDcRJq1fl3a5shSLE4QiCbZYDqjo4a1c9TETIJMwZrm8bwU1tc+jyq
hgYjf+CSTetLAwDUm9EpCftQmJbud4FzXrPKrv8kXNCDcjrDFbXAEbuzVLggvH17
fRpeQgb7Tl/afSTNMnndFIr0cvaxAH4PCmLRbHWTsKPEW2iq3Ghl/vzwmQ6KOpz4
ilYfzUTZOb7T2aryHLZ1bjPxq/NgoEWxktZ6DSNQtPXVjlLuD5CTb4+MZ3tEqNnE
piC1vNXzwV6QoXXrxmWgEMgF86uuJI+7bl56q1iKKquDvY9zYZk6OcSP9QtrQeHM
t3o5UFBOITH/cvVB5MdkpTL1RUDKNhATmWfog6DOylFuQEeIKOXyMTfOQxljbfxr
Hj9FNpBOTquKpYKrgqAoDFdiOcaOvciStE0lU5Vn3qGyH6de1zUnhLU1y+1/NASB
E8UbHCxyj3ltP6GGnpi8xi3bXSkBurV+Eqt0yvxbYKoGv3EAbsv/2hKDFrClhiqR
AOzR/kHNnZPHUJlT9uYHY02vpww5g7eceV0yEbMeG3QBQu6eozB1XKqtpT9QeAJy
lrT6W0RxWvpw35ToDVU4JrIFHQARHQ3Wgwob1l/mAWv6EaAWEQpIla7XXLC2tJaN
lhe3sQejQ4SE0gXoxeVIHIYJ5lOpZ1K9V/cYSGDAdkpUohLGlHXBBpzcXMJg2qB5
R8d5Bh0Qz18OuU/ZOtlbwnYWMjP3cxxji8aAUijnnuHSWhR7x0/6Tbt8VvW2z2ve
7IbmUM7kVkrcjKsmJfdhgi006Wc69AmxM7ZSfAdo0LsKJLT0jEtZfV2IwZCZq3yj
G+qutW5Q9wbS9OarQzFIJkLk6zso7dGX6UZ+uVRkher7h9GzQzsayfs388X1DfeK
ebs6a+AXp8XLqZrY75J3AC1d+GpURhMaj9QgIlF71bAEzpf9TwbyA4hztFZVgnOq
slLJT/WAFgQYfdVtnp5EHy9qUtovBlbda2gQLEsjIcwNr2IB0OFhlZ1sLRxVUVly
GrtVj1ywREIpe6Oekk8iiv0GB9rjldHEEhUmG+weI22OzHmcUe9sKUiOJGhG+X5I
N525Tksriw8KdIPwXiMQdGZ1OvESAoU8nRl2nDfMpf4PWtLJM7FnZbcgsLXX/vmz
BHt6ncDH/G2gOD+hUj1AQ9SKtqeZheWFz9suxZADn05sWW1mcFz/wUfEjeucvyvz
h5T7uOPro7c5m4fhYNd6fqe4RWFOuubDb51ttNyrWS8QqordOQ/N/6bLm678/Z1z
KBpjfiy/cUShDThlUzIUD76jdXJj9IBVTYmLzwoPeBWSznteqVhqrlZvqcdt+XfE
uQd32UA2ySmhKIndb9Ge/IVUw83XwZqVTaLoXMHpCaaxUyCnuZ7QsEsFxT1qr7GB
pESH3AMBDq4L0T8468kfVWBwRPjdgwNIWq0Z7RW2lDIO09lWXC7k7lTbBnzjzE1a
cFKQXnZx6DjNBZhkkVaUGFblSZ7zRaTeeb7oOJP/YZyIkO2CdKK+G5ZMTgewdnMH
Ij9d8teiDAEKgtV0GGTKll2nj85dCF88ro8D0O6wJNA1d3Ayl76DD97nqj8d8d65
RYX8bj3G4A4CKr8iWcdCEvl8spSW3GRgGvMyehXD2h7VNQ7ageh2ZF6Vy2frUzKB
x+rlp/FuE9fdKluHdgsF8oJXtjxzo/2hreSGlfqmk2mGUmIuMJkTucYcv7LOG6/Q
pGqZdH6Lvitw+a88F8UK9du4EAkyO5pS2gGIGbOyfz+GluZPqhHV50K20vZcx4zp
ZjmiC7kb8iG6c2oHbKfPHqeyaTyWz0Iob2D6FkmAx3MuUMVwJ5p54eYt5nrcx+zA
4VqV5CEV0JH2kJyukpjRr7/8Imt8ouZPB3OwDXeXAp6tBx/8tLeNQ8NK6/xxQCTq
b5P4S5P1s6FQoEB30nxcRfjfOeNu5Cyefr68iRV96GMcS3xYzs8jxWnx5NsnQCBD
zV6fmbXMi35/OppZwdludF4xjILc19kKGsr1p++v5o5OKjVoRsKxsFYvDNE9wq4V
Bwkl5knYqNhap4KuitRG+GvSisAPMakjTeLu++8cII8+iPzuKJWLc89FjMPBRUAA
ogMesac82GNoTTxpMCDvUwE7C+NTB+PNs0bVeWVcVHJZcw6EeKP9eX1G7V2APHJR
qkmFW6ibJvji4v1AYvDD9jm3jD0NHSD0SgyhRAbxMZiiBIi917h0BWVd/iQIC+iP
PUGZfgritlzRm/nnyR8+S9wDRMMq5MBEnehSK4Wccq9lb1O13Ma/eGMOsW8z4tVc
o57QQiS1VT7De+BXadMbRZjQumNDu3QWhQgCGo2Xz1o2osjs1FPdujvjIoyqAJ7B
D1UMLgPuSmLbi6SgaL3z1Fzua4G8SIgtehMKpuHQbhYHp8dkf2N/YJAd4i613iNR
Bq/ftOLN8ArP9oPSAR7CbU++XnWkHdXF9XTTyTWzF3LWQ4xw9d0g1N5bx41450no
FTf+/vjCoJn+DfySuq/ooCbfKB8QjInTHLIVVYx7xvsrjmHq4eyzLHYMfbnk1qCl
KXMoOu9tnv44naIe9vAucoCGSMu3bmcQOEcCd60nNGuLk3k0bz5GAmoXsGiTj+i5
xs9k6eWrVNEyrKHDEIqCZFfbjCJ6a5txNv08UkArPoMyLWy7SBE6kHt3l/Q9V/fz
irOdicOXRxIKaskmUF/95F6kae6engHmLeaqeCD41GiNK7O2sYl+FKK0Xln5GkUK
iTQGmXZ63pOqVzRPJtNWmhpypLEFfSeXfGr4ekYvsyLoWKdopjODzb4gF/FWatJ4
KIARrRfMo13sq802oP9GSkquW3ClbVsWj/XNGdVqh1uA2Uh7LBxe9N+2PJ5zy86h
SaNYsMx+B8GACBT/y0N2oJSF7NdYbhmAcl3NMU0Pljrh5DH2TChYBnac9AFqsSfe
AhzAvGXtAELQazu/6PgwAt/MYxiXwaQpJbqNKHBqQIpxcQhAZGm7/pbfKWqpqvIO
Em7pkCB1DTG+z6ym1nRNUemiPodKTGoiC9IW7d/8/fFZGRkC4wjC2u/5+31q+HNi
JrmR3Z2t6ABTHhKxQEz1Cpii7zcTVMwIIKLbbnpfK6EwTwezOkZiQmggMOY81EeI
05lw7BBns8Gx8Z5b4GuFQwq0ywWFLlDQPkYDq9zbcszEwPrnAvfY+CHRF1vOnK3O
ooyVU1zCNkYQ8oSHV/BH1tVNc2ZaEuaIPwtyeg0Q+QtXRcKBqgAAdNMGT7a1faRU
u05OC7H0su9wrNS5CFU7JYVtoXdwekEyveG7vY5Fa9iAYSxMn4JALiQ7BBZ9qgLk
WXRqYrgV83GEvlge4PHQKgeZ15P5V0xr2PLwvrFuds1OGv0trGiRfxhMNB6/Zvel
nmcd6gIgUE/KasoAqUnt0W0dB7O/DeAptlKDpFxQAeKkRHaOgbM6kK4nK3kW+rf9
TwUGee2aHws7UiF05yiddmbi/r1nCz6j83SKWkjOfTl/ODLIzVCxs8m89jHvb6hi
ESNNly1LKtlNCo4XH1Ys0OA26CjFpF5pfNmttcSGSpob8mTWnFbea2faw0GJ+mtf
12NHmTfvlKpcEn0Na0fjXJOzZt3DbIQ+B4KNTrUhAG7jhgm6V2bkXfptxXCvvK7W
3KvQooMAM/3VNCLZifqOWJMoMzVrqlkZUMU6AdOOxMZdYHjymRTSaP02Ww/f4slN
pVErBq336El0398uowdBsNEuNp6Pb1l6ywx90jAsYNyfAwAwNsPK4heG+AXQYlNi
XEJRdhqbV9gIWuEOxYq186ljKrwmViLU1dTobxL+5ws9qyuB1Azqofe0HAIheqqe
lY5ut6pUsPPHnMDBBldw3BZ1u1XRxnJrFwEalzrDiI9zU3JqAF1M7ZRlGDCD4G3f
3R5geZGPOVz3pPQTiEvtmyWIkIPj9LvtPpvBNL3Da0osmRKNlECHkxLTbZNx6b3F
6Ussyz2TK7HuELZDRGviV0i+iWCgJyHoZ6R2P9+aAJIpLXqYZBCrzCN9xmK5rIQS
XaZd/JjxPqSdlDkmHXPYmnFqZoSFV80do6yA7PNcLiSetlT3KNtJgCnA8kSPYoYg
pLqTrTrvFaYPn7FzMIQ/mt4HvT9xrSmIxYhocdBYXzQw0Um9R2LPGC75Bcb5ZyO+
SnbNa6sgzkl3vsJs4S7vNucbkIO5OZuBzvQYLfAp/RYG3V9IBv/y8VYbf5yT/8V1
Y+VnNEsBFRCAb5SZL7JAGtqQ5v2kVBAov2nC2jsU9Xeli8R4jYQYxwJpXSgb40FD
tmoq4xcYTV2EomVPvKAA4DD9RHA867VSvUBfRzY4ODKLiCJee8odfu5f4GwMVEiE
6aM7fzPF55+YaMt3QQCZTxWCThFqI/PZFBwRDDuU2P5oDNkC6al0MUK3KJ9PvQ5l
BxK222P/R50uTQpIiXeL/ChIY9sR9uKDVwWwo8kBmo+T/itDVE6kTfhR+7hM0AGW
3iju7YDQnDHTfVZ2fI626rZYrGE3nDCzUHu8t9T+DVo7V8dodwEPxoTNrvxbIoUp
keogAlXTQpQkXIHuGwHaJIn8FRUTJ3vSXoDAHiNE118yYQmO/Th5iPKMRfTs5PnM
CmPJxnNCWkOnSVfh7uDERrB/3EZMSwcNUwnHkLsj9U0vSjkTvBBq4iKkoCe5nb7v
fV8YtYndzwnMuFF9jwWRi2TRa0r0E9uERjzg54oPStksIxqCo5kJ19jU5J+idH31
D7S6Q/DPCtENTe3BlJTol+nXo73ejsjEQvpuhmes9E6XJ02bGPQaFnjQADkf120o
4yT4g09nWcVUHPqHEfwjvVXbS8slBNuXBNm8pl0mYKkfZmPyjem8mR7DoDYnzORG
deuT6gwH9WSu8pyNyVRPlHN1EhS5qxCSLZ7FYKeP2o6vaoOMeRPEYBM2fGBEnrYb
7l1qtyCx5ysZ+G0yxjqrJoQgM2d9J/JwZjuTdo8YzXjOumYmS9cwLcFGvsTGWPBd
3Xh5yycJlgiePU2d+JLvAZRmqs5O3SXF3WKlxhFNqOJnrqaMKX5SsJS7Xyg+GjJT
WSofRpTRCwbmD9RZhioi8yZIsaSD/Dk9bU45WUbxFuRHCuRS0wN3N+kNW7KqUZys
V4mUClCOpeNQwKgxJmBb83MMa2+PL4CYyP7/rlI6K8NT0DmBwCT5a4GS7oWOoRZa
e0QgmHwTUhVgI97JbByb2Mf0uJxpOVtbCIWmAsN5ggFKcI2wk4aBTTEf3Dl7E1w6
AQa4QZ0tg0Q1//HziCMk0EMF1ZaQHjSD7PSOfc2BF1/aj/T58C+KU/I9fL1N3tT0
SRV8SPXG4lhefhXSURmcNfHoV/DmwXjrtToqALTvsz9v2h1BqhkGiq0iJ/iLe/36
6Jh98nTbhtb70o6l165hkqoPXnpFL3BhTCSU7tfcG/6qkhOZEIRJWvAg4UFhx2Ir
pF7CkX2iBNztgVk/Ig8bQZGHFSG8+bqaJ+R0m/4npiS23hxqnuiWQOOhgDDTi0g4
eLjPoIpB0HN9kmQrAxJEHG06IvFspScVR9Hmwqv226Lz5JqgZpShG3SsNL9XYahT
Hb5j3F5resVW4MCoHiSLsGMeApzeFiwVfzS57WWB0blAACtpSItjiztA7RkCYVO4
Jh52XmDd0OLdDAD+KvCgpsX/EvajcuZlsf/lIcGLpw/hppV6tYR3+kfJ/rhexw6a
M1vv9H2DNVvA6wuIUSAa7bM4tbnOWzwW59hVB28IRngYpHIUTDElNDp8Nk/mF1KE
RJhfwqHget4a+Inkt96uB2qVyBJWb3XrlKIeNr/Se0gcrcbsfHaCh1jEF0tjxFg2
E2ImjDaSAGlUAfn2yzVNmNmndxd4lm9EokxRNG0sXw9dgQCbAGoElMDfkjA6yw5a
WblDMSmM47RiQ3abl9mdjUz8ktVZncH2dLAzMyY9yw5tA8oNHMq4ZfnnMTW3Vw6H
sDkVm2S/rWW7pxkRGZZIIxtmHu7uJKG15v/i9/lwoH+5+atrS7/mwm579qFYQarx
4nyWzOB2YVC71Rk2cYNSkRMtFKRJW5LCzuBl0MXN9ocKIvEz8vlotveUWmblO1UL
r9CqTXOgGhXYE6tyXCbbI4iMIZo9WB/aYkoVerDbmbbYt7vYFaV75DyaHkMiZ6+m
N+RYeHIGYI1R8s7Z/4R+vrw96qPdnVrDNIhzbAK/Ik9UFh+snGor3vRuued3T6zA
ZGp2L3kga6NaVNyp5tQ9p/mnx3Iu4h2MgznRaRY5Y1+D6sw5JrYiHDl+dBRc0coZ
Cay121XCQYFsPh6mCb/qun3MGvJssoYurUwmaujQgCRkavYuSdb4KNgO9JaNmKnN
YyacKYaNyAbm1MujUEylRv+/8D2+WJpWe72qSiHDfZCyxhqgMS0Y0fZkBpSlnMfq
BNdz34FhjI9cXWpn41lwESBQASR86ZhvsG78u0dDVnEVEnpid8f3C1hdYQyGXB+a
9JLVABCUshxzjuv96wi480J/3DuZko3MNqYx+3dZvYbYwG4jdaMY6JPgCUV3cI34
/V0XIpQKWNy9bFnNcvXmHnao7cw+5jLpQiJE4O6gnchVwUILXRbdyKgRXb3Tf19I
QeLllTAjlN2KSSNrEYyaigmhure5eoHhNu6tqQlXWUXlBzBHQLcGpiUltJy1xFrT
weUFrfTaKd8+IFjmScQmFmvxQur+JmRvF6NW3vq1xhwtR+njP1kB7SmEXhLNeKTF
uRCRXieFOb613HNznHfB5XRZwApexE7PNJl90wxvZ1aqOVl963rQPylMNKVjPcnt
HRyrFPKz6bubxj8IY/Tbi8iqOyYkGBZr4ayCwQcW6Z+vQh4M1ExUF6h6nfA2ueOu
Z3kbCaCeZz0u1cBVabZHArkbmT/mU+xM4UR5o3kiYf6cRdu4VpO3bRQg47MBYiUZ
hDhLUCHUmQlqp+yu8sfRa6wxgmVML6phV6HbtA9KueIhvVTHmz42LLthDCsIXY4F
/0sUFp9SbyHupFwOATxmytipFPYcBO3+L/0cnTjncgdXY1no2UJIu3ORKboZv33y
77r6V6J2b5Yr0UXChpDUUuL70M0SfiJKKlvyBbbVV6eJODqiaXFFlBdFI2IhYoab
InmrFU0o/J32QwcmnPbHdZSQxv7t6RubY5MW2cLdkLZ01Ru19a59qLJQjC+Liyj5
6x1rgCRtdA/raHrXj3wh2bLEbpY/q9Lf2/Q04qplkKsQLcHP+0g2N87KXKGklTTN
YuRiMNr7R+5BNucn3F/43IIIg+/SYczMNAXS37xXj9JKsTgldb/MDq2GTLA6p+xH
laNk2B3JgUxgj5cgk8uHkGoRDCEsZmxgMY54zwL7xP6EuiEByGRbocG7YaTbiJie
fYvEKyrlErzF7z1Dy50E8Oha3Gt+uVWHq5pBSQpXs68x2cdscfZj2g58rq0QBi8N
oIdqNZmwqBBQ2aiYUERgVb5MbbxSzylp9KAt6G4l6T2sjh3tPXOq5U/bFjhkqOzs
xekHVsOUm2Lf86KOuhEVsd1MbtBAICekLx8RHx0kNa0axR+yLRXB8nI5zGzdK2bF
haBVYr/d/vBD27gBVBlTWwe1OFAGe1Vjgr0XZWssN4ZEzhrHynmnuvhG5wIVbMj+
JwysF+O9G67fmxA7ncglQimQm1V5AkSj4fQmeIMThoJ61RqEsfmRe+q8bgZ/LnWO
SspFZbhp4cnh8CaEceO+43NS/UkLWtVxLRCsLmGvpbogp3UgOLFWhrJ+1pw3L0p2
7dD/jqEQbb9q1MjCn0pCyA1k9VO8JQnNnm9750BnEsVohn3uZnX2Kt0c075wYByQ
KXMjwBOIY9dyWmqz8F+STiyXCksuI0wKYC/8DOHGrhtx3uY6CMM0p6dSWnQDl0Ly
14XMEFYVbsoRjv4be4VaRSvMPYtz5dENmY85iVZPTkYt9pSZLc7i5waPCqwQK+c3
xZfwO6zBUFqwDuR/sMTvS3Pkl8PBzEGVyXon3+iYvFpXCyKxfV0dSH2NZ3jGfU2s
cuTGRt2nYlv3D3RzDPR3nJUiYwGhMIswDHBwrBeYX8Tic74ea049roIRTJCmduqN
Ve8hppPBE/+lQrQ4zJDYvV/4oTvQLuwKZ/8bxGCaCqrLa6XdRRf11k8I72+DnRQ5
ycc8fHCBLma9ULJW+1bJLsA24oDl+YrPwe2KvrvoROLZJ9fDkTY2oznhn7XkmT6U
gVJc+BOPg2LKTZoH450ANnTVfil9yrGS+g1zLGRUA/A4siPNYmNTz2joZt4WlidO
wECdRgGSj0D/s5OjrRKZ1Q7HeK4IeMQGVSEk2cdVgNP/17urzOMjsXPYqKGNvmxd
j/zEPPBDAlF4KVCGR7dgz19c1Iv4z2Y+giKWKIj2GFlIrnb8MApPMB7D2BwOv4yf
0BwnDNknYr2iTrEobCemosAipXZo5pbztQAXGkrBywS1u5mPBUyrTIKRJffS3qD9
Qx3OwzXsDHqZ9UU9hLGwuWQ7csT8jqCB1y2jjsYgvxG/0q9tMSHvCqijNftOyocT
9p4INtO4trnAM79yC+RAhySig//X1+qTsjz671aCFq6Ey+uitFkflmDlTrnIEUp1
17U3saDlsPX51ouVuM7OxOk9577SOHw+WOvuAPVpGVTE+/ChtNYmVeb6EzwHmrRl
e7p2O1mXioUOvqAUS1aVQg7FCXZSh7C9l9B6q32QPY4Y/q4vwxYxNtlMUMq3iMeT
Fexe9CZekGUM2Tv3isbW3k3ltnUsCUQOGG5adjp09nW8bB/Z+JHxLiyG7CGQvNmq
PDkF/WelL+KY80dEAMRbV6oQn8Y+1Ge86rsEqi4g2JJ9VujvsEcunfgt4fcDk9ZH
xZwqzVkdS72uLnbnCRAELr8we6Zocya/QOYxkA/C0MxCupv/1zDGs5PDnzTsu1jd
65PGBJaCJXgXejoFfHAAvqUejOynqDpNRnhhRXAad+h40Ykwd8I8qUko9oSED6tl
wyzIbWgID+r9ZRq4sO9mfkaOavnwJJethBTQDyGjmJEvtLNoy2hLai7dpZo5ehDK
o6CchxYn7aK4s0nIjfSSxeZVR/p1OjjbqwrYxubg5bb3DRrD1IfCtLdy6DyXDxTp
AUlcu7VdHdqLPc0nkRqUffciMTweCUQZojeAowPBjfwLkJRacDXxns0BVSQ+oMRM
+wrYt63VhNL+oWdXbRKqIBTJP1klvDemqTeFTapZJKLhnA8QGxQC9TQzWFHtqq9H
gt/ScTXrxWhL85+3Qszj8c6s3NnIRCTZhCFZtbBTmGAK8hc/JkAYUP/jxsfknNpW
BaPYdnr4ZkJL+HRt4YTDqhs1ejXfjuEqV4H2E+QISWk9OWwPLPvxR8LXV4eXrHuO
M5ma0HFIX13F1bEsQhgN+Kcsg1ZEspd45r9BiVSPFJA681gzRPlfaY0M0bmnemDt
ScxBsWrB3oA0KSWRwY3SX2evRySCoRxmZle3D/HSLC/5rFRyqEVn0+Iy3Hqn46mU
w3IQKmfN2OPGinwCB+fQ7xJ//8dH47XzjQCY3qBqpCdH2lNucWfa3UuFDjcR+QmE
k0q4EV0ohl51NpBoOUEi9KilqFftf5U0fWTOjchbDhyR3C4Pd/p8gWG2pOG/iOTT
UkG1gWhmobOQovjzP/Hxr5d4NYQ+/UaVnxUwIYEoYlkby8PBEvsdCfOZ6MKNZoqU
PA/Fku1ebE9iIzEqdTsTJjivkm89BHpUN3QUnPSnbdkL2S7K5QpPdfkOkQVv6016
wTM24Aymy2tT2/sNvG6aunDpCSdC+WsabxuC0Pb3etqdg2feN29tTYNyaQlLXZcZ
noDWNDWZ56oO8F4p1Rv38vt5HQEApi1v8lzHw6B13FbLnuiQQqBgHZJd76h19BdR
NcJu4CXd956xN1R9JT2y/0RLENomjIMHupfAr1EVAHibgES42qS089+sA03RAU+T
im/lEeE9I9O9KXDtBM7yLCzu061jAi3od4u2r2HeuhHXJulAjVVI8wReRaSIl98u
/Upwcm7iFwqu6RGoTq3UPOR59EQ0Arc39+FIo4t1kUHj7FXrGHvJGWx0979M4ZlK
z0RwkpDc1Bd2KxCNB6qf/e4RxC80Cj3WnvvYt5s2kO4iDbHPoA2v3vrGZjfwFqQw
tuAzYzsKeSp81CmLslvWYDViJXv3O1f3JiR6ja0ipRdZ1ovMYCP5UWRiDAa/SiPz
JxsDxYP4Kxxh9re8pDhMP6rZCkUKVJTB8lewHK1PPq/FkLPmL/ECwvbKhqxzVcGE
FBB262QLupJJCwNaJMSMh+hBD7AgEvoyS8Qk6+JSUBfotVb4Hfuw2iWTFVrvNglH
4+5qamkZN0X36ekLhm7bTfj96r1TlrP9x2CRMW/LMobo/rWlVUZPZJbW9Md+87xi
caHHpKEkw81hMBkaBWK4ZR39j+grUFEtLH3QbdwId6oO1soNwgEn5NejeQ9SDRg2
RxkldaPyg3REu9Np1iw+uMYsip/AzJlB7LEonc9j0E9MYjfXI3TM2xtrqfbttjce
uHsm52p3d3JObXK2b+g07K2bQJjFpTxJH1A8bj/4f13hf8Tkmyt2eXyhmOzFDufZ
JXowjNID08N0O+W4avuEoOvM/wIiWBtHZOVmht+qBYAv8Hg9fTkLG/Rhf7+6qCms
x8Fu8lhJVVg7y/dH06omXb6MCW8Df9VsO/zD8+eAH+u0bURHbuVNmh24D0t7f0vL
JnSQpKIGeBkZIO53O7Mp6a4KIN7yK0FSO8DJGSF1zTzMZ3Uk1MXdRPIoTmgIvDhe
EJY/SfLzW66FWpRGAihMNcIq2FCVLL1MaOHHy04kO+8WK09BD7j0dJo4vzQZrrlL
G+bWRhi9x4ryYHc4OYxSyON3A0GJoro7cwfOUJ9CTDCnnCOf3Ww9pmYE8A8Omqie
OtU1pRHwhlURoQQ0DQl3Bkc2tKHJoJ1c4xAYGgjwHrjqZxjVdQN+et3MpZXJwG5K
A1gUgnmhqDEfJdZUT194xMLVfbW57g5ir/ZFd9BFOf1yL9qvY/I8UwPNMequJyQd
1iEVoHOxHdoGp9gptDnWvb46k6xoq31Z89p8vka35BOAdE6qopd2OPGHoQs94ueX
cXCezRKBJtY5gUeN4gbxbSHam1R6hjzF/O9Twx+IZboAr+s5WyDU0T4S/Q+NBGqX
SgBLuqNtmarTFR5EBCHG2HgisLfbil6lx/DDtkDSDJtfpQfzQlCwa29H7Pq/ivbJ
Kdfu0BLTVcOH1SxEUPvsaycIEG9RolDsBm0YZsim0alG5pi1+vkaYlGMq/P5hKtm
ajIFVFtDUbX2n5uYUmO8R4xscPTjZCCeGG4obbANacz9c3nkwqAMGROP3EpRX3g4
8+nBzVa43wqpbk8tL6sVu7VxZujdxSJdJ8UOldiE5Ec+iINsLtnFNxENl6ncT82Z
l4OJLaisO8eSEBh2e07YbSLJl1JfQ+cVDLgKYDJ5BtjaLIHo6arqF8dTcbb1xAem
cj4OnAARpjlueh1ovGBVhiJeY8BAkT6DnCVsgVzpF4T/I/RZaDNYCS1vt7mkmfiS
CM/SDiGF5G9wuiqGcGd0/wE63POXU1QAtwJPAD0HdUOjUEGFpfK+NWbicGSkDJ39
K3q52ql8y0cccOl0YkZLc4R7kMSh+bsam/uahL2Ts66Idzb/XZe4blRjMrxw+Itx
HGZJEJc/WcwNJPm9Br3LxOK19Y3lASv50gowxZAFIJ8apbTTiGW1WOeeRcRdzMjL
1mZnRd2H2A6DkWxIFPf1O8mhmEIFn1zGU46D+4Ueu1XyYQMhI1cB57Jp7mip21Hw
UKoeC+WWWbzImGY2ahnUt9YIcESX13wxMgMWRkXD+4cf8JnMpoQW3dXoX+mUedm/
C30xs78xWryf+KSxH6gjej9f7DABnwA62LVzFgfGzrKy5gwwoU296e2P+Z3KuaB6
38N2Q02gg2DT3DD4XBjXXIFPcd5ZTj1KRgjEArwH2hEokMKrLemgXO7VwLdju1Mg
w4cBcnOlswqcI732ZISk7W9w1Hxf5FCylymut9XLYWRcpMuO3cjl0rB/n3OEq7VS
VvhZKdfjaf5QoRc4KaxfWTZIjHGqEKqItpbl7B8gp0uypj1ZjXvpc1nNurHiN7IE
HFXGBtu2IwvB6p52OpPsm8ByKRLwYIoJ+Ekj4Mts5MneEW1HAZDOE99aOCNASJO8
Y8zdb9ltwvc0qF+4Ook0zV/H+lOOS6SAhgmnX4+m2s7MaRdxT08RmQ9CuQvYdsug
e/yQUQFTLYupvntupeA8qKBL7Q0WJi0WBh34kpOrA24PUqUQOU3z022SiE4Q59H6
R8oz/mRkpzm6yMuNfp8MOwpYwdZXsJEqUZOez0Xbc1yyOSqog8z11S/8hUD35oW1
SAF+FFrD7N18enlFnWzF6Me7JXNNxWkTacdy1BPMPARVH34yRUJ1LT7vTJpVJUah
Mv/R+2jg6Yjs+LiEL9mzRXNneQR4GeSYWgL4zr4wOeRrsQSy8yP0LKVBw1BQbFdR
NS+xrL031sENpystHMl0UCPfzCabYHq3pvlYQQahFDmmhkXkLRJoG6ZXrDYKD79K
gOgoLtcR/GvfvHJGbilLa5WA+g2Sc2APqFwgvofNp856fH4TIzGksRYvebXsXlFP
u65Q+lZX4/nQEnDILGoGBoBollOp0Y8HdLtb7ekHmAKGFKfEIO6ZzYZgAWWRANJZ
yuRpN7ZIOfY9etFl65ClcsuFOfGv3JrSF1/mcQKKXRRmcJWtJa9nch/YH1pycmlX
ZUK0ZMIwDp5q8OeapErK2yMQhgucpvSNspBCEQTfvxnY2tigVotZl/QMMywk/UEk
5klL7hCichIJjAKqmYtR/aSbO3QKXJRvYyFuKhPbd/NW1Pd+QgWx+g5e4N2TZatM
e8wtRzNvQgSan8E9JC2nATdBOHm5kSmhMYNrZOr+glBWFA2L//Wb6WnrMHpEDPes
NTkfHnoungArC4LjQziAaeUPNiJ/a/irx0a7BSR0RjBWoOhm7S9tpR1Zp4oZXHYD
ISRnp3Co953X36JhwAKS5msr9zhdyRCkTnjKgDERyVKb5WKV1hM4T0cQSDiAtsot
B0EEQOcKQghxDKYuFuwrvNLCT7iY8sIkr9DSjhnOk7Z4dNTtXeYOKoEauRdA35F6
toSAh8lrBUV2ypno+c1BL6pLosDZWdbNB318Woj2nQr0Mm4VzmmIdlscKYtiXQpW
zdSG1TL66hyt5bNFVr70jOB0Vr3GQhy/glQ+lUaZU6g1+huGQH0EGOxrUiguK9tY
tFcBtXbXNx2caW0BUq58PZwxrbzyPsrXqBkFXyWqaIL5di+8lNvLvs5+HInX1BNn
E8dTHxH4hcicF2Ah6tMjsu9TQT1qUN2LCBhj4DyteLDdDTgaBUZuA/u4Y7m/73Lj
XTU3OvLDtGk8HLMIbrIltZuOyG3R235If3bpRCc0n9PzstgTWJMHP7VMiXSnENPi
IekqA6FtstgjoY5/lLNy3lI3nPI6L4Pnd8Uf4VU7qP6+f7zS9yJST5DcRJp7OpR1
6M3tYrMXAIPfHWm8O+G7rVZxtuS9QF6mXbKQ/Qv2xGvPvtJOOyyl3WJXLgDQweLM
BM75iAwKYL4KM0d4W1c0H4SNt1n+kcMTJxz45LvGhIhj31zT4bmzJDHDFMw1LnDO
E8mncM9cw9fhyHGEJ2YX41nNJoYjqs+ZuxTSHZQ7DVzV15AcJ0vBsIDQpxWl9XUp
rEU2NSN3KwD0DYGVTnJtm4IPNBgLCnVBSY39G1SXhBe2dHLsEmEJcmRN/3F8SHuh
eP9DflHIm9PoDd31SIYWeLjfcZQ4Uxo9IsnTqMfBxWKhJGkL8S/coBJp8EA4m9mu
BqrA0kLGMPPriveH/dyG90uoNVhUjVp6hA1z2yqBph20A+pGXV5E6HB1+KveKDWd
G8vNVp87fYo3HHiLksmc1UK+Y/IFnFmXTJpncqAgEzic48tVPRALB1HjscuzGo06
MtZXOGOX9U+8VoxcTUP18LHfcKPXw4Bq/k2yz7zCMs32Ye90GFJqraBE4RsuUYyD
vZR+OHNsMJAf5nKTrfPF9pqv7NLByA6GBHYoG2xQsr4rvfgPoBLShp34IHwsCvqa
d3+hl0iZqKHW4DOxexAsAymaYcZ0Oh+jwxZUfUGvzLN2vWuSxY1V+YN76jYxxqhG
SuGtBy3BwmYcNUZrbseFZAFnTTJ7D02PVbwM1jhj9CCoXZMLfFz2JoxS4+c7IzZ9
RKzm1SxEo1Y+MmtErphZ1t03cUaZsld5fUgjfcHxAq7V6P495kt/5cx0nNzC5B3I
Emwg/ed/beW3okGJJMGoj2ftAO8PBnSn4nJcJ4G3NqSyhDjk2GsAa+2ruqlYkN/W
hNXog9cxJNL6I9rCdaRWye0T6vGrr8kIkMavxzcd0X6VTVtsqlXI5Y4USFsCw7WC
RQ43orzhjEtmM6RTMDtAxifd2Fu7+VuzwQyQaBeKlEOnwb/oZP/AOKAg6wG1kwOF
phHK+979tn8Mi6s6P2al7vTWK4eKMHjQPct1yxccZWQX7ijrMFYP+QZLyLJld3ah
VWRZihDiCTjQQ9+V7dKNIK6TlG3o5MITt0Eg6kSZcihS9IbQmGNTkKUKUjVy83bm
iBzJ2sYlDQwy3Mo0CxBsZhVSS7NrKQbqLY4UNgoEVe3YQzGyrpo0NIC3W6M8g58/
Kja77Z+J25K7MC6Vs5Lvwfd0Q2TNaTg7+xG5fbMoTgPppqmNwivD9VZcSsxYcD2m
3BIMy3uyead/v4L4dCwPahin/JTOGDaicyBtBpywuzk6EeVBCXASmdFUblGa2e5u
uursZFXqWvLM4J/B3B7auV6w8EMVQNDzjHgKikt90zu7ZYvosoytrsPwYXMo5AHP
C1VHtXxr57sDgjajNfuTT/zEFDgv0lTYVxrNb8O/kozS1Z1eNTGSmup/NxI56Bxh
vDlS58nVtaPe3K7GHOdi0TRc0RSABmmvBbAv+ufdCgs8HC7fFHuc/vwpfioIjW0M
EFg9iB3ww83ZRi9Na1cAsXJf3fAEr38PevnDvkdJL8hAYNcRUG+dzreuM0WSxjr5
i7xLiwFJoM2ZwWjs3TAL1sL+FbN6Jtw3G8G20bICcFb5K1iwAHW29NIteW5qJsq0
Ec96wq+e6nUtNYNESXxG7DaQ0iKy27m4DY5+WJfdnXgpG5zvtQvG9jWuwDyp3+LH
S7J9vxKscnS20RaIm74nrqDixuO1M9j/SWLoqfNsfwqh5hSeFKJsph4G93kwAvxS
XVpAk1bMOvHkTMtQx8wmulU1K7uEKLHlJtWSds/NmGqtWzWzwxVrfWulvcFn1TIU
YGsDMHqOpGDrqCFX3e6N5kLxj/hig3VF1vWZzmZSwzcEtuL08LjwegjlziN5DkbV
JDM/u02k6y4RvZLmkb+lkLIRGO5pHQnYHCn3Zs3wl/gu+Z0eV7UVl+l6UtU/IcW5
ythK6N1BZYqChY1djOduCJslFd5NIDcdhTyH+sh4uEZmU/bt+GHBIcYiLxTIwShA
7OUEFRdnpdy8HE9kSu4OXTL1pfn7rfHRWp3Flzsha2dDT8EeAFv3TAywsHNspiaH
++T79r/OWIqN6wSMktXbLhnZL6+y0fh6NWb/nTrNvB/C5UA1CUf/uHudfHbnhmx0
HAACrbRknKv+31myfFrj2wQsWTosaEFiMHx/KnwwgHi71WEdBeVqZnOCBFf1j2PI
hXAV9hTYIns5lgrmTaFQRGr8m8fvH5kA8mYGTRLa3mO4DZCMVKebniX/6DPJgdAs
0uQwANKg7KjKUhIYLQ45z+rOVgnJfAvdmk11mjBmudMZh0P8wn4vhM3d4Cf1RrKn
JK/e9hL5CWMp6YTaAIPuiA9NG+SLpvLsqzxxNNL04q7uwjvJRW2+Ak1k28fbyf6m
jbVHcf4wfyGK0bCC4x3i19MhJ53+5Qst3lq+2SJcyW3M+ioeJa4aUl5e7nMJ54pz
OaoBMfApQ93oT4tF7qxjClHfKOA4w8W/NskjxzGs+cGEnOce7JnEJeu0s6PdzH98
NO9hz8IgbSeBLvA9yx4Ns1q63Aj/RFTUMgc7L1sPNtWOBPVpy+ybqmZlrFlbu44R
codrZ1zH1q5HEZptXIuZ3ZyMA89wb7lKs9fT3jpdVyHJc6kZEAMx4koXVeTKEEvJ
DaTXLhhyFG0uOMmJ1sye1+rDSeL8m8LJbO0AdcsGHjfTth8cc+8KpV1d7GeDgE07
iHqRnRjLAJ07lUVa0PIDMiFG2DTXJ6LWId6PxmzAdKhtIZhQLE2d1udKxs+tVKbD
TOmapxPTpHqsnp0wUN1i9pcOh8AvTohZyufUV3p/tI2SpHhEUvuvmgkqV22ESuCv
tkuRXYGCHFeoKheLduyNvyTvcU5WN+9ezJFsg1w2EqR27a+4tf6Pfc0Z8sUkXeqh
OL4/LsaJIMNJ/pwLdTyHfy/Sue10d5W+oje8hF5QZiSYukwirHF3RwSTPFa7acRx
cH+Q0isabTQkP3r8BjzxIvtgAPrEpiI7qvzeVZufBuoIhFK3JNold3w0/p4Hq7tw
78x6uffZ/BUduYAwQLJLBKtwAAkXAufx6ltnZPlm4R7Di9mT6uSXdCPkUvO8vXeV
+mkbIDY5XYwFfO9jylZhECTvsRLUVt2c5kXpx8fkMEGqJ4kLAAETa6IwVerThc7Q
PI0LkPwgfpAxjUqeRW0l9QZJ8dr7ZqMc6KGsFXAAmDekPp2J+z3hlAqzJNA51EWh
QqOBdKGhyKRu1tYhN12NT9JXm9OmBMe8QHmj6B6nax8qxZM/mJ6IhP11NqpHqR+l
T1TOlxIQzZdNjIFsOAELIjkH7lcxdd09q9DpqA39jRjK6DFXAqST1cIG61w/a0Qn
X6CIMj26l75Iw7esxPgH0awhfQINhGZ26hP4LS7senUgScRKl9yReLiI1Q2zRrmQ
4yXvb4v8ziVXYS3n3dWts1J7S6exBfnwXNPsU5HAnZIOByfAf4g0tFFE+mCwv8RN
3HT9RF/jecDOeiU29Qt8r/jS+yPl6xcWfB7qD3jRel+Gqh6xjEh3XE4l9aBXl7qj
OFdI/W7R4y8nNcIY0fXzq4z3c6Esyl7+7rQZLdG/8CVQX+ou8xjoqI9QaRsLFVjH
UDUhQU3Wlyp5RVOvLYUR9N9T6g/bblSZIUAKgidvRzSUw6dj1ayXCr/lA6ea/eAe
FGtXB/sVOsfCcBrlLq1k3+pUszvl5bCfDccG992IdZgQmvcWKJpSeAs0UJqLOL0d
KniK5Pn/vIaCja6WkuVKiXYyBNkQJvD9POBF71rCg9plHZSjacMg0RCC2e1RzU0F
aLAlk8g/qpX7YVfs2etGe9m6uZKCrQo/kX8+L6dPVvrhAUhcIWcog0QJQKYvl098
dx4NprLKedf6XWnSjn4xeB6ungo9c9lpkHWdpHimcRtOUQ1ZPqmDkuE7SItHtfLe
jr9yf5fczj3WTTYnrD4TtcAE0wN+MgBru0gv7JldcygMK7UMpGLarPXY/RWNqk0v
Qn+q003+PjIBM8q7dv4pQN59EM8IXq3wOrXMa1VRZkEeAe1RXPhjktgl8FrZ1k8O
mQDC0COSQ0IyQF8wirhBLvTS3mW9NIf94rAeg4d4R683GIT1SVq8vISt97bWzVPO
fs8mTxggZwtBcyx7BubYb3JLOb5t6WQ0PdsOXWiUitxBN5PZS322bzv1wfxr200Y
S7bd/YoVLmBvIcY1A7nNfX8qV0u/OJ2XYaMdpHGh481POdGiO7F5xitaDRVkIFS+
l4BODEarNEuFd1o3EWB7arhdbtPE66cC7EgLqNUybeScwob8/kJkl5EHieHBSMT1
XGiR00j70WNjPP0Gz+YyEovQ/R3rKvfDq/9Hykj/J2mzQxlr8psGPAY+p+v/LIFW
pb4ebwsfBqq/uQ2TavWopskOCtNGBJ6dtG4YeN1QaV0uDQGsn5Ei9EDf0oWOeiCE
KRl3fM0SxR76c8Zdriaz1GNdwHR9mzyfT8mLoA4aSZW0gwD4pH3mhyadl3ioABD6
nAeVKRAPeDw800/VOOvnKBO44en5WjgB1xYepLamuP+8/QIwFAAbZHuYpEDmR4ZM
kRDtA2g+eE8an78Bywn33h8QP2CLNQzjy4dzzbvImp6Bqgg6S3Xjp9bmcZGyjtxX
hvDmKpPGtVknOIZQTQxl4h+ISawth0u9gW4dSoFMNUXoVbbr1A4KuJX/eI/mZZq/
dXHvT+5w5zmx5yuA0XXtskS86MPooiyDQANanO0tKrrqTjtSAG6MFY5NdQUZY8NV
jU4Waq4QC/ZcudQ40/iU7/xyikWvI3JycjeLU3uui+gciVPcwv3zLcdwKjV7Hj0w
vg3HsXLgd92+evXKK4FQ/MXhNQqT+XUYn4qZ7f/nyxBUeuP5Pwd+zRC18hVA2jWN
VABUbeECESDL6toN5Gfa1Yrc1QqD3EUNVSGDgBzZWsdbFUHI4Rl0wxw6V5qFy0cS
Eu2+MzA27bWO4GVYzWHgXT5bkD/HknZF5WZNY37hzDu3utyirM9IAxA7KGvu1kvB
k9DSjePot3I5OnBfn2srESwUAmknLh06aC3PSjW4FYExxCAUtrbR6m+Qp81Pn/2T
Y1StbcnJT8HAuFpANFZBLpwI7VV855LA1hfRGdsct5WAXX1yf/PzjM9ScQxpnDsx
B+wjteG0yZoptRw2dgRAduvUZVVlIzFcHb6n087CoE4wPk8ntDNzabqrNdIuX4Wf
JeBctFUTmEqOIGt6m6PoWHYOS2syzRLW1ZNOahnxcUF2hW1bCtO52KGkdf7LgMdJ
gQhqeeg31EV5AS5TSxOu34oeX9oFhd+BfE/h/ecaLHrTIAmYcLx3szUH12x2RrBp
mXhrFzYpJEZLqPs6sTbaYV8IhGRA52pRrMqz9CPh3sVnqKotnFbiVIiZw7dyrN4z
18wIKbJnpHzCyJl9WE7SdiprqtTDCdNeAPTPBIySxkpR/dlEbBQh8+NsZktzI+tU
YmycBOse0AFNhWJQxIKBMYdSjqN/w6gpcPps0VyrCNkt9BagAAQKWyj9gvso/7uQ
Y/ukleL/2zN235ioQDf1e1NkiBMDnEPO3grLT57XueyG5DOsqrqGqu4BFAYTTbUK
KIlFljISv16JzJGTXqBFIKkAJkr5MVEVA1YNDP4i0YvYOyuz1RWesc3v7yFDe2Qm
Lt9gWcioYmixT/fjfJ54bVWwBqIyXk3ataEfkjkgbJOOYnFZGFmWQOIzGDw8s8Sh
D9+WMbtV2dpb0aisg9XpohTVNLcSq1I1sx/mjS9TvwIPsMFIBLjGo3ZBBVw0Zzvt
i3dHM3c2FlbiL3c7ihrhXjihQBaJSS/uvMOCMK60cvqsK+9+Dm1TZLbXRJ1QoM0I
9pd1Qf28oWdPi2BqvH0rrjGsxtMPxRIfszJUBoM6MtXDR/4J3qzLWYESzVKQ/FlT
wiCLYpEAeSZEq3HiLDD2F3+6RDq1oMs2RW5+S2oMQRpzd48T8vHZ4mIXxjtGeHcO
5leh8vcxAgoojIJ/IIgjhq5qG9yRRrTIJO/y2PlrxS6yVY7k6RPsu45jyyOcsxw5
r25PERF3iMuaWof2OxtrShWwHxGztlh1M3kbAwJMP84qCXZ5g3wxpA4likCL1aWq
tNwIfDeWf0JahSrL+7xpnoMRMvRirx+myHjcwoOceoPBL57QHvLp4iSAbKAi92GJ
Wm9DzlXJfQAcmZPtrhQ47iFUUHC5pwSCp4WfwBH7P2AQgiV2ZTSWF58mnrGXpzmf
rLqP/sz3lGKGvoZEHPf9Kpmx1Sl0L1bbt9heYL0vUV1p8JvOWe1WaBb3Hn/53XtR
7ilOKVHsYcVuxvpHx+z2ehrIGNTpK8r3DXiixPC6tVQW1W99yfBwmTIydRcs8jM4
sZe4/w5zdjRsnnBTpNPDv397qxW6KM4OuzcGVWGZF2GMvhM8h2eWrxn3l4owdYY3
oAH2LmwxlgkPWdw+Y8APUimtyFUcovqDqwZRXlSoBUX3r+agCkK/k6nHei93YD79
Z+WmovYK9OW2h74L5rjKGgGqT9aW6VfZac/yvBGtLRrRiAs8qvXx67/h8tS9A5Qi
wktaRtc9V7yb6/ADnMPNnAQz6A1sS7KyvVeLk2dpu2cJRDRVoNb+CVUVdswgfTYy
MJGFkpg2itlU92unZO8dQdzM9p15pNsUMx1No2XNinM=
`pragma protect end_protected
