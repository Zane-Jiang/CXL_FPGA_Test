// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
W/9QpsmP454z6pYU55BgH1CFzXiMAYhfS3Qy3hpWVJ6XQIXl21NNC5tVzi4s
A+xe9CdQNhJrCjQZxyWDBHJ91hIiYRc9GyJV8DRc6jmBY3FrJGppA3ylojo1
CjKOoEmU17QBS2mguorYODuYDm5vn6C32TWCzocRbFs6f6k7rCUG0+SvEMRq
1yX10NUnll/JMsYbQw5vqVC/XZh+pZlXKa50+gE+rUd+Vf4/+xPpIlY+3pDO
FpOE9WecrotbnkduUbOIZNEGd5putuNrXlSjXFE3ixZB1TnHKf75uWKDoNWY
Y1lxbJ9evy3l2/qpHJsQDQrBPLKhT0DsdwIUjIsiWg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GfC7v5CZZVjp/kBuPgEFHNjoGvPkjmaIdRgcZ32GeP5tm8pAl/TopWrYmpxH
1U4kJqmF4FK1O5OzQbp+4st1gwFFMSeabA/CwnuO33Mz+jjQJVddmPUfJtJe
XeXSdilMcMlUXz7GGtGqIplyVhCEZoAAp3d2GmXL5GKCjR+NZqYC0m6loI5v
wJRHCkJnNIdSbisbI1j2vMq6dA5dcGDuu7L9bdejmy1VMucLyFcksnk2ThAP
r1pbn6kwwJEXE79pHMA4H2Dd5BJYDNjnizcdbYaGeuQhQuCU3r+JK6syY5be
f7UfY3qlZVUgKMi5YtJm7XZTAeCZnhjG3HsLFKzGzQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c2C1VDGh1VE5n6wsagrNZrilU1bkA91x7oQOMJ/eT8PB1JYpQbOnFBzoYlrF
viMJG79IbyA5C5xCXHZtxP7Ui9gYuET0xb5VtUzmXAu1AEqse57nc3hELn08
cCIX2QDTG6WRftehFN5S69I8PUTq7xNmo0hPQrOkAWzoF1KiLt3XZjgIVhxv
nLD/ORZS43ka2vToXqML43V1ul8+XHvW9FEqjmjrpKftcxfxM6ZPW+f9VRRA
6JOJ18l8HLrQeFbFH5fQe/5UUaZ5iUtQltjkR5ReIHQPZpkwNzHeORcfZyoT
VhCurs1MnzP7q3rpn9u0pU1t6KQbY7qsSM+XATa1Cg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YEcDeaOV/hQt2lZmVFdLbYvQ+I2OGzlwqXYCyg9/hClyMeXZPyweWiHe2kOb
/I3BmJzfEEnvOa0B8C39nVWj9nJqzHcZacKtJTxePO40KUP8jHBuUEJXgzcF
pR4l89NCcETqVaS87/UBeNqghQv5XcJAk1znYzeM3iITkdWsqX8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SAxVe/1PBEInoaMKk0LitT7ZhaEsz005b7utpb08Ro5oQDyYg5hbgM849bsG
BC6szr/tmPy2vOyZTu5EcdIKDmaANmiN0MAlSqooawMWbdkti/mZWZ1d0wx2
7/x+OvwXWSOLDf9ebvM5mxEdYiUdXBM+JnR7p7IRv10Z/fIaD4M76Tp9i7ls
luDhwGs3pRZyxUKmzLOHZSSy33ovL3YN2tELaQg/i+7p84bHPPGYwQ0mEOjF
R9XhC6Imr/jeF4/cJkVXUmkSPXfYB4zsKE/uVXkFXUCjDa9abtN8MhhZJfja
O8Gq3Fz3sKQ7XfyJeULfMQyzkV8vldWQPq+m+euxwiq3sUdj+3HEc/BRG3y4
SsR1cdb2ltMGnl6sV5N9dqyhfv1Rp5eB5ocI6OdkvnLBXBZPN26qkUvADLfQ
9mrtecZdVzmVY0/7o7RmkOVWCv/ym+X6YG+1X9iR2kbAl2tEnTJT3QYawze0
tc/bOUkHGOZHPrLHa4iKgHG18nBH9aXf


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dQsk80xr9QB0P9wBTiyPR4dT4j5Sxgmxz+dl1nWdIOPjNplh4YooGEDvzA66
qEr4h/0qzR0GUiM5xUHR6GVpTJjI+czQNGSahKdMJmIZuC/59VHZefT93lG4
++cXcAD4k89Kuh7vrUdlXrjBRc54niwX6Nmg/Rdg9GAQ5b1/LM4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E6cE6RtXIaCZ1TwB31TnECG3jApX27ygEbHDd+G2bjk6pp4wQvC1G7ABwW2Y
/8rWVaCgWitAD92VAAxC1lMPWEASYaTpxpTJIdXZpmsjJGBcMJC3dedoyWHH
9G1TiJUMBsd/4uD3vOrAPh/kWOqAKwgxBkuo5qu9w6bTmx8KZ0c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7936)
`pragma protect data_block
l6xWQ7bbAxWpHaSogn2SGcLHEmzTSM0/Axk1dfW9GVc3RDvkSdxzl1+z3X57
agFqYfsraatAYPqI1zkuiIEiMUCZdpGa128IoNCPd8U6kGu2JXxKI+ZLgVFU
zYjJjXJgTRJtB5cC3oqH9zbZaBv9iMAtZJeOcg3GKMS6cMWpNCwuWu1DU91a
qyEbWvfgaZCQqlvrgm0x0R2sC7X6/+RrovxfMTqcQdM5UlxOSsjDZTEDKRIl
zwPb6EApTcVwGmDT3ZLwTr97MPeQQTadBi46trcw08NzqQUui7+w6Pi4+dzN
HOeY1tG6u2y7jzRLsz6V5mZZwdHwydQzZ1u/hmCF0bUa1KDoMTcU5wnTczqP
+X43wAFnju7sEsTBWIJr/xMOWTqRS7cW/fy2pI7AdssQa3H0grNzaTl3Z3z/
U7ll42DO0ROxYGU+MXikn9Cbz0h534wMXJT1mTrySmHbo+i6CXd7T9Cdrpnz
ikwLpnCiMRkAZ/ed8JZ9A5PrClN0Gq5+EQqZOaN6+Dp35ygRN57+ghfJX62s
cVhH0KXaggfHle/pxbjtq/z31gkiiCp2pS7Y1oFjbmYsVwrWow2aHUXviG9L
J7tMu6zY98pBAfMDQHkBQKni2a3KWSNXEC/qchFV35QFHPsJLcKq+0kW+r7I
7W5dGPcQw55NiOQaBRUyYcMy7m25YEWNA/s500c0abYdOugKNryArC8eZ3Px
N/tiI+yximoqIszmhF6BM/bNk5WBEBkRwA4UMMJys+1Mzuwhn+mRWm51z8CL
bGdqG1IhbGiqcEynVMT3Wlk9kgWixM2WfSsa3ymFon3QfvGcstuitEqZomdZ
GLPcqleY5f7wqIIVzXJU0iIQ9688tXPM3cGo9Jg2ujNJZTTDg9tEjF2GDjCs
yAmd8LC5SrbbPkQcOf0DOgs0T0/bdIOKC4MuUDcuUsmF5/7egGRxP1ayC120
f8iZOgt3zjmhTG8rvQl4tDKvz+dELv1kAYsfou89YZe93N1r4eQCBXKhB8e/
Rr4+g/+ALgrOkh6Mn6t2ZCXjf+ZdvEkj8/wYkSY3JMTqOdY+VWFl2OszuIgk
/WLI2+BGYwHwBFZz+ssllSE37/Oe/hKCkBh3Tw4wYECqgylGhLSEjffXoxUz
zVfmKJVT17jdf20+vRnTJGvDSEDwKfaxUdXpzFIVEuUZTwmfhtSxB5M/V3bb
pgbY+AlVB3yyg92nEnttwT1NuD7XjRwjz4wqvNmYg8FpKGgoKAhIGOgoXNGi
rMvjD+fWYtrMXYWGfyW88JVww8Mw8QgBlpY3HfV+ex2gHC9Rc8+p2QNvkWyF
kb9Osq2aH9vMKtJUJFaf1PI3JGniQ+n4DtggFPIcVHispBfnw9ZqIk7nPKIX
B4El+vRP/SJv8LlAQxAwQ7a067Ks6imtnapfRsvZK4I6yWB5HAF3tXMJOxaM
kRjcn9ns45RLUc6iQjsab+IN5TU3Qn4AuFGF2jrJR6XQBFRsPXo/M9zPWdhi
kg+k63shrZjmu9VLVwdK+tS5Fn7lIxNqKRVRpsrXD0tU93NgXH1LipyOpxCx
qCDhQ0UsQG3aq0l3CVUwcEV3R/UaL/ftVNO03LF/piyZoBQXkmGTf3BT91Oq
X8rZJwXrLmfbvXXTZ/MZgPbssuMi99rJN/dA9l4/YdVNIst4nTBs7dw4zybr
pnr84VTbIHkRif8qO7XzZwPlo920ILXYQMKB6Y6GbJfBx8t1jrWNQ5+kLhZ9
qRQtl5+1VEBtp6VsEDYlRCqwZ11ch0eW7OSeKiwvUGD+/x8Ceb9r78Pjd97Q
vgzkpNNq29+hksMcwK+7+zy5vSHBtp+64K1awQ4V6sJBGpB9IgNAb4nmcq2R
TWA1BGaySYqWLfFtRHcwJgzUNuP9jMxmQMeqDmOELy1FnDrB35gC1X+1fLH6
r4X+3pzbvl79of2+ZgYffzIpnYtW180kxmBlvNY++B+SwFWUxaVKNjnmGCbh
hIxu3/ybI/WynL3nSfGAPbrxn0duy++en88gHhh99BwksJYO0yo5SuXfgdA0
K3qNR9jYyYX8JrDJ4gFY4ZtvYSHQeQUX4A4Na7LfbrU0BcdRR0LEICrC4ljb
BfkGX5fnAdJLdPaDhDRo4PY3MVJH9SLy4Exy48gncQ5ljgy8xdQo+WleleLd
TlZ3kSs0HhLsogVpi0//4E2PSq8zsu/h1tdCgickBy/3eI9w0LR8gnMf0E4O
PKP65QQoROzmAUZazQhEJ3tV8Jz75i4auRdGqKNBPa7u5xaKZuQmDaSxKQCM
Qnl5gtTPa16OtLEf1Ldn2CEY+g5irAMrozCmcqbGmdatRGkGAV60ztpmcCBq
4LN9ctAtyYwdfpattKwUVx9KgI756AGJgvjmr2fVcSld3ctE3sg9UhPc+9KV
v0ImbpZZQLGTyWQZDhWLTODH2FPhq9FSPZwegRKg00YAIo3Qm0SgFMrho2uD
TzXq73aPTXuX9OsWSGUu5OEdJqX7cVM+xIbN0DNJKauVyqxr6Qt0HcltBxdz
BvLjnhFdhCQPP2Kw4nLXIXfSfXzj3QNK9pMd/RX6ojW2wagl+nZmY04KvtHy
rlixOFPvhcUF1M8F0fS/pQEuNImypnUy5kyX4yBRU+wDM12uPRgZMCh3debi
KTmR3cG2kyWm0mD5TVosaRBXaaSaJ7cVYXIsO5wnpDgEOSC2iyx9WpVq0sqa
xg2MT4heg/rDf8Y6siU6+7WUGY3CtRoHPRj5Q5Qy12LCvSeg5mdpvi1UhS8Y
oOi5uWwd94VgAE2RkO5komveJzlj0+ftx4wEIj01K/Tb5f3OWRtDEamWE7RX
iOb3AkLNSFGoK9hLVRrTumqXxn+O0LI938ES+Gv/ZvfKsrdjJZI6ejPYFk54
v6rPg20uYWl0ScjWVhY+3o+zUXjDkEJZRdn+7PXE79BvKUb+qdEp3t/PDUhm
cfBfBeLTC67DGEk5AbxWSl3L6TIYbUqGT3ESCkBvUUyw4cqGrzDIylQFaK3F
j6WdLH66JnhTdWe/dMUjUPgww9lAQQyNqvrYv5WMADLSInKnyw/17OQ/PqbO
2bZJle5Ydm7U3mAWRCzL7U9tB8f5OAbxHVIRheRsxLCgU5rFk2dPALeYQc5W
fGMKETO9ne/T5RYQUIVuPqnltiwEpdVU10xlWzJissGjnCat4HwXsCRJZFsr
8w4CcAPFG7dc18+aurNk8Bo0rjagRDsMTOlzsUy/UbfKD4zGxh/8kjMS5iVd
aueK1Q0Y59gYTGClF/6XOqGg3yFM1doIb3QwW8/JWlMQ2cU9ruBfgApYxEQ4
u8m6/QzaPDmpNQt8lu0rmUqMP3MpzkYo5T4yiuYKTqWV9RNxYHPZ1XkWpd6D
scYY6BG1yiGBaPdFZAOBHp8xSD78JnCOB2BzvQ1Nvm3GUBKAJ4KHck+Tpuhk
+T57kvSZqETMhsM3TjEkaYNxn861R4IogdJicylz6GapwKBVkyntR93cWfEo
EMM71oHRzoRDC1mAVdfCTTe2mrKg/QGVyzKryXRnWXgJR6AXmQpiytZCTAhp
hUNPimKKo0qY/ox3Y7fQt13E4uJww2kyXOfXhzANFqDYcq+XV1CnP9yInLdE
Y0BbA3yeNU4APvKZUz+6rCQUOWdkB9c2U70lX1RKNOGj2OT5ihej60PUcuhA
sEAFh/weBQ8RiFN73BJI+Pzb+qCY+cMk7tNQ39qOCCDJpNCVRvUFpmT5r5U6
Z3FFYwd/nif+qaD4SMubYqW45IxYp5kTot09hzgIk3on4DJWOujrwv6RtIJb
yfQ7N6PgIEnbL7xJncsQAeCdlN7cZP/SkGKPLuyTl6+sXzJ91G3wLBaCT7m5
cwufC3OJwh2Xm1TIgdNEXEfMZmw/CadhV5C1eaOOqbc9cLnXtaaBj5M9DV0e
3bGRuCvkQ6VtVFCeWAL6K9/5SgKDsJaqNLHPtrkVEHitSC6uLsrZPVihcOXV
9f+ruGaVNy41JvZMVX+Skb1svA/u92AKZLsguEvfhD2rw2H8X881Owz72rmW
O8aL+03p3PYjaglhJLtKOev515v0EfXTHTAt8uSiTVLMqrIqtbsm9hY2QI07
dYgwj67juaJow4uRKMQw21ZVKlRzl4FHNvgphe4M5we4Hq736NIvN2JAGBUq
dwIHIHowGC2HgRDf8vzBRLU88PnBuZv//FvJ6T/LZSSmm93tl6e+4I19SdmK
YhM23MuD8OlTm+sp5yWyIRg/bwRCMo5y1eRetqWRgWW1+L5CZtKEQ7XVSn+K
wPGCxL+/dUteUvK+XNr6/nm30wefYF/vCqF0vIXwMFwz0d6R8nYWcvhSi5LN
OA5AwBeAI10z7uBbP/sfXHxo0TBJHb0lWwx/u/YjnLwjPIHUhkLsPH5Fu99U
6v6nQi/eCFhALIXK1/6TDlPm/PQEQO9ndGCooAdBiOjgUaDezT6WRySvDSzF
ZTjJGY/aWI7gsDeiQzA7fBjHT2TaltBOR/xrpyHDqOIzVqaoGfWq9eoCZ4KP
s9XQvbkgblkC3i8UnqGEH4TuyVC+butPf/xSJdqsJ3ubuGa6yihYV6anDc6M
tRqbtjHSmEqlF3Rwy5O4/LvRH9sncwk3XeaKFy0NKoORQgst0pn0GASYSQmU
aYGFzRDVNzudJQjY13iHzlD0pofbEH0VhmyIWWI5X40ckVMDAclHMDyYWuvk
HpzKPnbSdGBdnWL0g0fLH/WUftwBOvXg/WMI5p0EYrT+oHP+amq+O4nf7LGW
r7mddxo6EKB8d8ihZXfqxryUOwsRA/YWue3JeSWzJubHIBW9MQL5NTkN5UFs
G7CxV87adsBObpiF+HsO1PTDi7hAyLSbPy1drhjqYigLqVajBJy/lJjj2AZb
/dTahZ2EDp3PDZDTqXb4Rrv5C3AHJaT4w3Hbao1AXtun/R43VDl4n0llv0Fm
SRkoO6TKDcGBAsf8zkNsZmKs/h8iGijnKYRZm7hdhQH/dEH0QOXqWPslKb+U
GmdhSBxYqxFHqDHQ2DMkqcbSRznfFsYabAHs5nZ+hDANtMZVcT07g7DffqYY
XNROkVvCfhCrb3KlewtZtJ+7CT9WX53sO5ADJ2FLXzahXJb95+FHlHzhkSdW
C08KQpSPENJdJWL/drwWN0VNzQK+MOSvpTist7THMkcnPY96jbXdh2/kXSYo
ZTX8WBpa+hHRwhJy9bkNl14li02P7EZFLxNESKtIbangf/DTv2P+BNJIWkNm
6TPaNo1ZZWe8S8xd5qZWLLOWhClPVdaLFO2CWZerFWgtYlxbvM6fiqcn+Zwp
FaRXa8KehaEqitFtWC7PLJuzvHM6ts7Db/Pp4CT3r8KENovEkdZhyCCYvm9P
FsmKzzg7KGfOmDfOVgFBESZTiGEbNE0FG1VlLonDuKZyAG9vg32AibcRmVtO
/sUlN7iviK8oCBKY4T8gMteuJxR8/dtNmHSccSR9EFKOFpGNUTi6A4VVYZSe
SgRDTJDVcLa+ANL1IPCw7ZQIKGpWLuQ3v0c8WKUhhbQLOdaE2xrIE7e1LIQS
3dCligX6QESSEPuMYMNO9WW52+1+duFCbvLpZiqTnCjG7eXN/kvl4fBBh6XX
GlJ4NJ+AOOAb7fG4/pZ/+/wq63U+Bgdp4dafVzJmLwB4vUrSTQptWDdphAxX
XcjV9m98KS38gs/yjS2ycEKf5pFQusKiZ1+TpOf95nwoSwBMHrZpox9NNnuL
0nPIkcWy6UDbNzpyEgG//21HOCcB2hL83JJcz54Qc2qMN8LPZM0u5VyeXIb/
6BrcwZzmA6K1kxoKse0tFmJCHzLBegVyHR1DrPomNgNPVz4LueeNkFwRUG9h
GVsf9ulaPvZYs2lugO3iVYEpx1MxQA7D5Ov0zc+eHvHTky5+YSTCuL1szeAG
ZwvWoH8PQWyng+Wz5ZDW4ZtgwlsN8nMA4NBN5GZqoX33kJsUjl78pO5fyGG5
zpZgqzrr4WCHbRAzVzWqBiGkY6oCE6mcsPxQL2KtDVKJrjbmM8yNXBSLI8NX
9pSBydW2AG2LwqlcpmXfHTwJf3fnwbWdvtumxDtQNfeQ1pUwVFwpGkHibRZB
T4i/tPe0/SkBVmxhTbjc2E3qjTZF9588dGIzp4EP7RGZiKY7Uqvi/aKN2fXj
bxXpibUa9ZZ8pNwHwtTvdv5mO/knjkfRH4jGR1AegIf3qtSzuDv3+6HVW/fv
EeBst5Be6xMFnTbkRC0W0oieKJrVmRAXKvloBFIGM/Uu/Rs5h18iWU85du0X
xsbTJWh5CAWELg3HyvxAkBmfLomdata2FPZQTgbpaF2M8LxEiwIjFeSlnEBh
zPticqt5U2FZ0fyUB4bkhvzXH1G8GWSxV0+YBVGH0BxoV6naSajy3N5zaz+w
6oiYLDF0KSlwxMJZrEDhXWpfngV2roAY0MvibzhMwJvSPrs0lcWFWc5j/rgx
dKCxAAEoCzPDZqyIJ0270rjJuJiKY+R/xGMJQArnLgtv77PeKpi8K1jfVrS4
Llmhlc8Nik1NGsc7OmL4bEtEfTdzI2p0X37TY97DHiwFzs5PKE5P0ic3Mo2W
ym7YrYpjf1Kqo7Pprjjy+sBtyuX+MxYpUF+8pomlS+EQraYrJD+J03dyOrS7
zkiovg2Em7p63I2uaYNURTiZAfxVmw8xVz4xU7nlX/DWI12/1GgyFoIHV6J5
IzUEQIzeMFYDptZMgI88iRlFVE8+5LVmdMZZgY4FpQnLJEr8aVKh0COmhFa3
7X9zK7fdLb9R5dSi15Gq2tNoRoEjpgSWCl+Kg5c1IuCz4kNGAB2zXe7kHX7H
OkNMMKK7mvuRUfLe98zlumNLuITqKyLu9yzK37bNn2tecW1eA+8ox8B5NuOc
Gh2vW3lT37dYh9yhrXtoM6rgRQTg8i12vtQ8h8wsuQD/FFEmnLfiyEqGtfLJ
gI6OFTAkaLazDSCRNHdViNIEXGysA57neZX9iWmbO+RshRTwiR5pGc4k3V/l
d6Doci9A8d8oCTao5zufER0NusjE2mWnEosOg6KQqP4GNtz0RtbE4nQzadM3
uHbeBZep8CZNPrVrkOgwynuw/uXLHxc6iMoL5sVtQdHZB2buJubqQamfU/OH
5lGeZfbxUaM70mVzroum3dPejzA3yAIpAbMlIaCLy2wT7beP4kr18MnnLhTm
lC639MvPPq6mMeei4H1uYrU+X6NPuZ7T61y4m/S4wPKadWTITz/tuaD0OwTo
cCGNZ7KlnCWeTl2lBX36S65/pvgamJFx8anAQLNHvg9QkSRZBLL+cLkH2ViV
en+kZVpBjX3d2Gh4USd3JOLxPPchvU5BIGAL5lB/0wHCsPsOZnf156/q1tZc
Iu6fFv8MX00tfFdlywpmVPXXBRCrsGBPY9523m8oAtvS/Go3S3+Nm/1esgWu
r3Jfxk2dqwA5NwulnOqUdVMiFpg3iwIdDO1j44pxcKcfRQ/Ec4fA/2k1fcC7
VWFfbvk8ZI4fI3LhfsAj/H3v7aXWolf6zbAqjQUWZiw+zwoOygSu2y+sKpJG
LkRHxmrUYtR5k3olnbSCzMMyUxX3wPIxSklje5cH1gObqvNF4gNNQ5sPKOuh
wMAO8QWX+r71+a0+TnTKO8ibFNJClPrZPM/PByTVooPDnNI1UxDIr3iEI9++
Gc1s4eqMasRaSfOVpKcuPhzUTfR9ut118XDHFWbN62P8dlkT/1VUpAITrzDs
yDjLOP7jzo7H05LL0ne8wiOGUaNDwRXCNsO1aHSJRpMrN5aEzRAPczRHiwRQ
Y96Dgc2DPhzwRwD8ZJ+AKV74g0PScjXLfLMv1raPFWb7BN2F8jrLU9LqN7Fz
PhW/8hskDApx/5+wz+gsCvCoyenSdvzFK0qXfw4/q5yczZh/WT00mlyEaudD
qel7URz6FEvkYR+/t6AqPr3odhGM3KSvPDb6tA+vGF67z0LmUwIFDW7Wgl5V
FUT/kwZYTygPeVMucD/SDpoXntFW3WuFPvWzri/82o7CLMnvOLC5Quc6Q9b2
1x6mfyBayn3Ns+DSPISBrhNbbow/fLM01WMnxI2RMMGmF4Ewx7ZjmVhcepZE
HuwQJZffAGBb5RiQSXjMn2N1UoRu4e5Ir8V4KNLUqkZ80Q36nnF+SU9s9wYk
4Lj5sONml+OQe3NsRRA6uS4gck81jCv6yEUMU7qiC0Beq6iVitssb9G5Qrfq
w+nzEqDcsnj9FS5LQYKq7XU77fnr2vmyw21TSUv5igImRw+NZurb85G8O19x
2XPU1Kad6trjk6p7b1+LRFdTiOpCaBilx/qqu7ry81lyeZbG+trJqzx53JMm
tVItNkEc6iw9Nw5noK+x7uXRAly+Ea+lyhCKTDwUD3q4i0rWSvveKKBURz1o
tQSP1t/KeIzQ5piJB4W4wS2qXZjAaxtk9M1fxoGr37VyhF5PmODBwkxmxogR
dcOofUIAeZRUdN8VR5dCdkrQSbVklqG3QDD+49fGk06qQrbZJpVrLZxDcCle
nVSaw2sQfZSSkKS0HeRfGItc4rzbzZxvbF7rX01QVPEoth3e6OWTmeaBSKpE
5nbCTGajtoXP4xGs9BkBhOBwmV5Eyv6hI1Upjypyo1Wi1J+kMPxupA57ZkC7
6fte7uf3RClIp5sudF8Pb9LLH2k6pigea4tJ3m7enG7nblHqAvizRpsbvE1D
ioeTJ4osC8Lr3s3zAAlCLVobmFN3ihZuB6Sve8QnnRiP0efBgWxbEeEa7AWH
+Ozdy7gG2h5nnjYTJQTnxoeqKH6LyIq0M3tyRtH7TRukuZ3Z88Q1k6elElFV
kmUpe1LmaKycNU693P8O6eKDK0t4HxhXaCk2aPk2D/MVHMWrkdn6iAdXpPrr
RVHcfAmmnNCSRTfDdANbQE1OylC4TPb4zv7h/Xyf0X+5IAccMHd3tHYVT1yB
SlQD1IUpRDJ0GgKztTkTIdSmIVsU1yxKIAK8pqBlg0gnnZgS6YjdqRZTnS4+
yLniNtgFsyNi+JAGoPNakui9g5KXI/nnSoeDIGWMV3VEsSKSATE/fTbqN9NX
WDpNKPkWQcEWwatZS02yy/67s1C10REqn5n24YZ2jC9RSNgEjpMw1ILoU1Vo
oLz2MJPI7uc08JgnC4IpTtYTTFB32ZWcSHC47JXK/CRwg9ficBIx57ahZErV
/ruCjNehW2BD8VdMVwvhnLa0m6asvt2+9M+6ondP/G+aUX0keDRaAl6h+RHA
cz+cJ9TjZB7D8iJyuoG5Hp8ZxBqQl8Fb8Kpm9Kl3hp9wERvoyM7dXRQzEWQ/
NpBgOqD2xY22vSdCYjX6qSCmf/8Rha2Ac8GhCbIEspJXiqdYYAKr5uLzs8li
Nl7zrQqUm15rWFgssSB9fWrOIrc0UA2sR5E64YUY8xR2dMP7vb3tETEj4u0v
deyOcTXA9KngFmdRo/1bxTaDcgbf//H4CEUdeNhZvGio5SiR708wCPxcUA0l
XVvnyVzLuZT9gnZ7YVJiSMOhuUxYQbd2DXTzxqYGJCkam+9eVS1AS1EziwFb
p+J7b1eIhDFyuT4Wl7j6HRygFGVXw/De/k+K17dtCBDJOSK4JJAZuvk1bsM8
hcnY6bKVqJLh2Gr8w9Wyghtn1uwI0H0LW5SBVWxdFBQRKYqcqiRMsy2Gsff5
x2Npc57/7wkmJ9GJ3+7CVfc2nfTkUNqAT37zWC31qgh5WoV0TAONh+VIdT0L
8n7MvB7uAX/3Bt3wisfjk55ou5Uebi28uwCy6l6ahSx5qkzaMWEDOFyzTTsq
NENiuaXsmwXlJR6M2l4RgPKuKa6IkDK9F0Pbi0pypfpQmNf/32dhTRYFBaHs
cfEdGcHZV3TNfGWtoxWUK2vAzNKFUqDtvSFYjQXIoOP5vzTBfj9tRgSL0A+k
ukvwkEW9wRkfbk2DCqCtaPIKGkbI3nnjPywnnbyVB8xtHqrWARrX6iQrLIJA
M3AyF5NqVAfjy7lks/cgDoIiTW5KTT5/+Yh5LO2LsseT1RnxKcohhCDqfMIS
PBkL/VZvRC9iJANcivKDEYE3XwKqUDIK+nrhaQ9UeIR3ieMmYW2f3Hz74vxq
EcAfiCbT+VhEMkeLNA60A7EqLV9MY17FhEjcc0ajwHcjyzEGpnI5msWthOnK
oEAVsrV6qy/71rmhDoiOQ0DGwLMu7eLdSUaH6t2K/QMWleY+SCuxNAoVHPQT
y/xs9aRU8VilCX5qkaixigyJPE8Z7TaK7LAbaGMOB/fpeEDJzKcHiAPgbVO+
48pg/QDxv7/bZihvou3+Fp4O26a+mQXYfPcK9bXMi9oWokOm8VwJLHaPGp7X
feAT2jA0NPfdgbHRe38xtQuYG7DhNF+/PYzDIx2pgOIzE15VKCGZq4r7ytVq
BFzS1wugRiTfw7vLeNN26ffacLKWYoh5E2aGy2Zb4n0+KlaNS7F5M+A7qMgs
33atkC42nw0gXuw6U24sF7Dyil8erdCXdOitb/919cFILzRmXtFLhiJN0y37
NgEtQ4hGsnR8LnEdSiWHm0XpJX4ztHOi7bTWp1Pqt3PNa3aN23MsPVTMuhIt
DFJp9+fZqyGGiisg+Z2Z6c7pqkPMyQ2O7Nm6WaVeKEI4kyJaH7QOihPaWdZU
78fTjV36kUNQ+7s33daN1A==

`pragma protect end_protected
