// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
T5zMuG79UXR67F3sfSEmbWIxBvNvsKzD7WPRp0FqVzou4wXb+9kq6xASnZ8PftcqM0cf7e8CV6Tu
U1ND3NF7WaZe+ucmjMqJ4ULu6GGBpRzuMuk1fjeBOD3PpeeXHdj+htuEQS76PqhVTqsO3BC+U5wI
PZSGLS0chuZS+6lTVbEvjHesq61qU8rqPg9z3UVUh7E++gn5ZZxA/rt+02v3F0lGGPed8R102mg8
/mgAQZXPRxYPEvJbVsU4sofUkhaWlO9WkRfYUqbZHv9A5fWjrovKCzgAuKFz7C5PC6Zw51R/3bng
B0e1QTRhTWyiZJ5PnhBTOIJjsvGiqnhu8nmXhg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 29360)
wgAtIGYFXzUtk2Ont6RTO20EwsRToOZCcdu/HJwPiM/uVD5UfiHXQz5VsbMnaMaHSfjwhtguavCw
hRFQ5iPYoZ2Mjm3gUulDe4odjtIx2wFA/iH39sFZI4wrp7bS8/j8XeNIykA4rvXkk63RokPwrQMT
Z/A+Ss4EFN3zOS84xWDkYVv/TtxviTB9JNkC6SUhWub4Dimh/UK5kpwg2fPF3xCfZLbq6mU5n9wy
zIdsq0Ka46Bj9iLd2gFqfAjWySIbh+q19OKRTbnJdOfxS6n77dn+6n/bXSGZTCYm6ejAaSZy16ut
4mqN0xxlqhwmDAFSWR5GfFgdYONUw0pKB+mExX8S+dPcRmfthxwjFUDR9o/vrSVTIyXEQC/VobUj
I+3QNLAk9SNT0U63ZibvQC0G260L4EjPFcxGrS08rOeEzoCjFfWnxijRHvI/Cb2+N8wdSnn3s9aC
FS+0g0gfSjp8d6dRWLu5xX5kkJ/PflycVicnJaL6ykDl67ufiTm/74y42YXk7loID+vh9i7YDjEV
G4zUGTzWl5Ytj2hf7tKTFQTMpiwZtMo3d/FHZM3pI+5Bp3YCcGvNs/1GOHQ2dGUC+DGgqayHtzlF
Ae+Xd40Az3JfHzqnjvzxDsslvhCm1VFo0aJaR1yVhngNFYSLh708ebKy+sGw/wkFK5na6JI34HlY
G3VstxmNcuaBl9JiO3iOZgzxvdJsYCmDbrsngYodgF7yr2uuSBCl85qWLWCtSjzm+e24Jh/hPH0k
FKyVW8xMuHUIUuVilHxrlzyju1nhK8Kc6RssNkO1kd3sXJ7EDBQcGJaupnTo4D6Gm9dRa2+/KP3T
KAyMAOfX5UkyT7byECqCOOQ7T2+31gN9uHb4Bekzqu1YBvLZ5ZR5nSwQIosEJAK7+HCZPqaXCtFR
9p9rsuRGXUDD+SaRsmP0vFa58drQ98ro5amLEDE8f3fFg8M3gDOM1ZgyU1dTDI3XRYvtVDFT3VqG
7gL4T35PxFCW0MZ9ipfKa+GrDtOXor1aS/DO7kSLj6JqiJQhrAq8GNFGSCDV5+LbXcc96/IPZza/
dfZE8N097LVCM6Og2DGhEyJLi4k8R/TvtIRDhetpWfOkX8kafWpHdag+tED/dHgo6enQp832SMoN
cSiZqdWIFOrjivCyHejGU6kWOcuAbh7S92rsyxR1LPvDnM1TOjXSVLJZ+hqQoF7QcjYtqa7e66ox
dzBDF5jq6PsHm1FUcEkn6TT+yTl1HKg7Vylr3Mzudxx2BYpLOv4PUaWT3UAsQjwXEQndH4QrWxHe
I0itxfJNljBoKALnbvMoa9BA2uK/ClygtZ4EEZdkMo42kFJhblbn3fKhG28ZeteiR11Fv8DcB2bn
BViz35cBX3Lfhte3N8PU2cHXoYA7LlgyVw6hWygccTkZ6znRns/O8RNuTOi8eKoow5SCxdnoqGJ+
FZUEyQqsM5vjIZf2y7lcTBZsIYEK3l+iav5HPaPdyX1PhCaiCaJSnhOIKLzwYN8C9edMUVV1M02u
6SPAt3naLs+IAWGSoU2ORb3r4TnHIxckCVMFFAhIF2ZaEWt+eTtjcy+RrpH1vDmMGToTQWeuiAGF
Xp7dtSNvUrMKCKgRu42gjUI2ERU9NL0Rz8kMJEQOl3P2e8MSpznQ0JbgdNyAxsZ8y3S6iqhcYFLK
7cCWmy/lKsfCgTivtdlEYsBEfl0oAZFB4WIyI6Cxxp3+QLR6bzVCGEp8nnnGHH7xMUd1gFhEySFF
d5BHTPmKB8jEFGOm59l/3DfXZyqMc5K7F9mXEJIlQ9q9sxyMpdiXhL2NdJL2ecA3SHOIlncZNB4e
/Lci9eICi4ZLFD6eI0no/H3ypmR7rmaA3efxomWOl2/Pv6xi9GEmce4T2smqPOhGHeKdESyY05DO
2j81F1KO4gqf9KKa3eMyDTHFngf8fbQx1RjnYcpmceoNjw5DYhBJo5DKEw2RdnbbSteOTia1RRSD
bhVXBRoW6GbW6dZENjiVIhahWt+T2SmEjG6nVBoYQ1PT1tDx2o8wKfjahI2gmzZM9XU6r3E03YNh
XLSPlb3BywNsK9Kk6qDGAaX/CCXclaa+nDdG3AUa+lMUUdDCGkyX23oUYS0VXpm5mRWz5etDuaf1
XdfM9VLwjlc/NJLizFvbbudf6v32kT4cymrFcV5q4k1r0kurIOOuqmrS8KSFzAhHkh2mmB5nFIG7
O1zIV65EHdjwydXmg3WwHvk+oS3QDZLeOqKUy8wMA5N6En6PP/Uars59VJr2YBqjeafZwKpLTiaw
Qwiw3/olL/1dxXrHcoFq2m4DuOEf1q0i0HG8XVxsSHLUSxmWSnQ/95ANMraGTAoYWKUhNyOVgeMA
r/xYyufIc1Gd7RSotReZUu+68ZMD0OYUL8++70Cf4Xdnmmsodej4KbEjmfS7jYqEt7IWGBgNHaiY
N+3fA3axH44T0DFmnvx+Anw7hJrB0k1dI7c+2yZT0vJn+PGV2a9dqGEP2a3deiL+R6n9b5nS1mce
LMUeX4oJ0NhRdVT4UWB7wiZR/48UpL+FI6vPX0HpvktzFYCfkP7ijT9H8XA1XuUf3Dst+UaEELrs
w21HQMRAc+DBZxr1dMbwohqxjEbTntWfIDRIWyrebu+ICBsIkH/nkrQVZhnaqs//K96E6m90WRkA
Viv/YHXcrX5eABe21HXPsDt5O+cziQz8GLBo3Dwb9eU6KJTu3KmDiyPrM1jqlbDSYnTxGbwFupJi
IFU83fY+MjdCVpQ9Gn8hRTd8/5F/cEA9+9awrKSmeV1pH3DO9fA2fIETI2zDh1MHrJTbldblUP/B
yt2sTYXbGuW5z5XLToMWd4HyBqH36rnDe2EMqD6VDaeeWXF3w7aMe3T0GU8YrcpoCqaJzXagoJAt
AWvONSaiHPLqxnpkScREbJqkAX1Ir4kLd/SdSsnUn4BYZ2Mq7tVOoRb6nfKUiILRSristz7N5yCd
zkwkirclScD+MnMgGrbZBNp22wqlUYnuzGsbLKudXxYra6CUVr9txCJe2cFb2Uf4N0fJ5iEIkOOZ
qQ7zoM4JKLF3c14j7qbmjQcOh8mHPcpS3NxgpTGUqSmFa8q/7heUHQK1bUYiGKQW3HQNdffZtUKB
OiEZVog9sapCsil7CyIL7b79DgWP1dlFyI0D1jm4dfSc2oKKgM8NVIfry9SUP6LRHOmQVOaIYavK
jI7v7JWa3jgBbqzfUazSkZ9T5fT5TkwyCEqLlDQNf/SL0RDXxIV1fcUKmC0advjNIlXh/uYTd4Xh
34szqumqWw+2L606M0Wumd2b0EQVmpdAC2LBOfLkJjOXpGAyFPLweRfy53RaUf+q/ZKFRqKT5qnm
LyVdfHeqvSbkuiILpN9srnKqhVnH8H6b1W6PBxs2GS7dB9Dd/uXRfbvrllnN9Q3JVMUh8If7BxSV
OkC16MyBuk9G64sHcFEMB3EDZs78Cp+170cDBcTisEsoRlupZVhQOeiwjo3PzOJ4pL54PBcr9t4P
n6AW98gpWJ4OBEF+iv3dsuyw+GJR6nNxkqRiNimZrUftmoL7UT/wyuDzPAkIrSqvV/d9JpiA7TtX
KSl3SUfdVyGTE85lG+1SglZdAod2U9mHDmnugRVxrEoPSr8PSUyBzCAw2RYr34V1PHh+7n5iycCV
cJZMUHwbIF3yuTbi5GVjqRZz+nUatUZrwGZeDY6STby598JTJdhjjgIeFusbbhJIh265rD06pjjD
UAU+aIU9m+Mg1GxfCfkP2mi1ekTxd0pOt4p0Fxi+p/bBkVd0TyldxGFWjueIi6Pj3I5s5dwocCxa
oYgY+ICIYbva6OuIxRZgzt+Eh/OQMY1ejfc0gvb0gbt+2XG5CiUCFMvrI6u3nzKYGPvhC1l51eQy
u4eveaJMJUovrecYlk3ZTRrptcPr3NZeCiyTuPkjlJSi9MI9YN1aycdQJ5Dp9zRxV6oRsLxZEmCn
nOoSlS61cd5Ba3jwelW5JLPIaVd5DGNWHq0FhZwgpTup2qIPq/gwbwmxthhdcvXDg+rvggseiVyQ
IFvU2QaLCYK9bTgXfjDa0LREOYmQehU1ABlHc7PrUdwCzF1bO3DgB9jevDWs0PUSWvNQFW9vMzRp
gntLYLEJJkvxQm6bpEvA+HmkOd+yx2hIKMinlrdmBF8YtsK5EGNONKmgQl6Ov1o/ctDxRJy9eyHL
vChf6cgdUZnmVDK1Pm0WxWT0CvsdTlGHq5Mc6A4oXfSBSW64r5s5oxEdP+A8jJ0FpErOugN6Q7HC
8Tm/mlP47gSWK+xeW7ExHEhegD/vk2T5haeJYiGGKZbk2o6ztYGnAMOnHI273qjhZoVkhK6UPbot
Dlp/KnCJQwpU+br/TTv31jtsfyS6YnbcitMy/2sf8Aswh3GYW46xFMCT1T4JtvAgAVzzkgbMcd6K
Hy5Z2L7PWU6SkPjY1wBU9hE8BUArgHl7p71cBqCta7bGZf+WzLi4GFTpXbHNASwYIQ3Ri+IHpEGF
XVbkBAbX3u6hRJz2fo+D3V9pBCKIhX2GNjj5PS/rkAW9fu4HqjrR02XoOdyo2qObBJ5EqRwrYVp+
wGtDp84AKiuNkBGCr+JQHl8vsRL6ufQDAckjaJvTVlUjUMajOtCoqYzncXJJzqpYWNaB6nfgWix6
91FB2Ayp6ubeHwoCvW4GSeU8kwqoOOt81r4V1K1XYA1W9TIODnFJel1tnOr0PsKDLW6PVvRIAqA3
KRzNGo5oasL4AzmUhnWvLiAbJRBZGzn0OK2zEG653v32KuQpqycsYMBAk/3ghXuXtAHls/v7n3dx
CeZfSdct7rT5JpHPFZZrPeUTXX5uxF6EkFaramy4pM5ShPgHZ9PuO+OWB6sztQuM4sRPdAI7l09I
HHNZqODdD3kKaQWjAGNcv/xI4g5QBu5Xm7yjC3z3ZqQ1t53NVkbWf+E8BmpTTead0V/lKQ9nJdYZ
Tlrw23zK4d+e2kEDtEKPp+RikYPIa7SWoq185ZUWKc83yjdHvMhW79ogadJ1EwCCtioLPWKHZWsi
yVt8rVIZfEKAVaBIT0mN0lAR2btvOq03O5znVlTa5F/EfkSSagbRRpYVDzCUUnlGsPwP4DN2REsy
UMClkTWEvlLF0PB5DGhyufS3nUJbDtcxlDZrSVaKhs4qrIrai3B2JP4/hZOfLb3EJGI1bs4SLZl9
LJ1CyuT/UZ89oWrODV0L6bsvbL0b5a/NRfuzvcUl3R79PIY1js7lqJpvvhNmMtDccIClwFzGeEq4
L1Al0j4tfONiCAEwx/dat2HMCTI/gJZRrg47DMYRhLIBiyw5RJz6p3IPtZNvJqg8tUUb5jCzpiY+
Uizbzf9PvMO79o+NXCNjvOhjdMnzmZHl+CRjHz7+0NwFWsiGl2dNXyXvaMt1EvLvxHaRaH86TetK
/nTAF3TVIdyaXlZVvmfwbXufZHQ5EReCPvv8bnlMfMbO+qD5eW0QdBvPb92RRNzNMxKb0Z78AEa2
NhYn4Vtn1DoeGJy0UNy7taXzkUi26cYUdK2/vswWa6lnXZ3X/tU0r0/z4fXnKJ/yNRzC5eKaZS5e
iobmoXDe0L/aHmIptx4UndG0m1V+SpSypHk9aUShTtHqijZYgSDEPSbaTOKTpnZy4RXyx7MqrZ/4
OF+vSr9O6lOUwGhejyDqdAPKCwpT3SBDBXu9c9KJ68PjOgfKB18Zq6dSckepa/0+UQ9JyQP7IgOh
hv2wnUnPRAc3tQ7yjRDjXFtec4XmcWe2ZNtiW6qColZMAaJAHc0y5ZZv/YWf1eO3cwuBrtMo7IbT
fRir2qwQOM0fcBOMIDedMdsptKWbF9dbNi7b1VwKEmlQnR5Xp4NCGsNVrX3Spt8Y0tup6tFXUrZb
OQCZNBQ1Vq4IJ4afJWJbj0Ym8XPucZJYX/bDZqqoT2+VpmQltpf1NadtahWwTAFa337x00JD3Tn0
kZ/WvDoIZv2v7hPRYRiW8+VRaAGQJOMBuWl4hkcUmij02Y7vNoPZ9pbSmKyzHDyaY0Ti9c1EKUQb
N8eTaW2wS3STuowWI747jMFOnY0Qjc9A/EcG00v/lYN9wYUv8fC/bfX/83EYOOK1W3vhxl/UVJDN
NOKmvkdelA0eJ40LHWlFDSnW43dE89K/XylRTUOAw/ItAzpnTjyqp2RZ0DrdPPH03R1Y0NdGmKEB
lioZqyp/DgcbAwQVvT6Er3oI+PSnnR3rxHXDUE0sTUyjv7mTPMyCVLiVadoLZkJFVnBkSNzvK/YE
UkDmoxAdXO/7/blFcM1LzN1KkSCfBd0uUTod7GI29ybYbOPQfkoJJfRiBHjfE2oiPUhN20hmO9FS
y28Vz+Y3vEUea5zkbliGzaU4X8JVuvO7+mMDMQKrb5e7XG3DMSjZJgefZEIQPEBPFZeqRZeJCXof
P8d6TO1XG1lTIaCP7pdn0imxXD+DmKrRBAUF9CAiLMfC9vl3baOU7rcn8SP7503bSCOPSMB4Eo9E
K8uI1hISfmKu1aKObau9I1Aw24NNOgjfaAsL19XdZQYy5LRkimjhXrVFW7F1NkItG7bUuVJb26Uj
Yj2aUmKyBcH7vhpxh03LZB3Bw3Ej3eGpBLISeHAnNhe0UQE0FrXlSx/je95lgUB9wusA10YR3juu
VVMr5SwpWZMcfc0EMbSdGD5mVX43rd0Jz5FjGxqhfvWQiMVkfJyzvxcmntuDYV4xZfAiTT+nAJB0
G9tG1G2wWDBLCWWemRZWgiSwjXqXJhnSqN2+L8RFdfspHZfpqynAQV8t2d3QqYs/cECn8En6ofgd
qqJLQblzjaVgfp8fOs5J1xzR+iUhsnQ01ZLFzgQIeAceyBYdIj+t4F7VIVi5PWqR2X03LjfAJ3ue
ILbTmCOiI12PP6O9FXT0TgbFW/0D/Mjyjm/dzoTTZb6KgTH6AYDcgfLODhbAoi0L+Gl+iMgewmDW
YceBbWVyxXLOKua5838gF1FaJTK7geI+BkXmtYt8OUjErrZV4cQu4R7QU8yM+L06sm7hi/L9qSvA
xRVDmXy18U/TzrVumyfrBOS7HBjokMFe5x6VN627QcgZlwgRyw05G7QFJckowxtbf/JP9kDNOk6q
pctjz0j+0CC42XrmZh0NdH7o5+nPuOPcGDOE9uTSqr4T5ntYAKvIUZgcOEjnhX+BMt+uKpkrjqUM
xO36tjP73AEAHoJB9ZTakyb7flnjZZbAjOnNpeBbIx3TpDLCDQHOdwHO0FlZFQ4U1tBalGBYJ7K2
RKjf+fF2INzf0K72HxtACyrNoDhCVGy8g9rCYhXewJ4TLx6LOu5HrLH3I5JLs2XjscHLwEYnc+s6
t5/wsEH4rl5UuUog+jPNBezHCMwk3GZMJzqzm2Tz6Avn+REu2TcOniSfmG5Vu3KHawVWRbLsvIzc
6tPu1oMmPmaDc5Mng/JWalxjOo/bv99xrijDiCvRQPaWFangbsHkPcgfiKxIO4AVFOaVxnjxXJqS
8at1fE/zeJPUgLv4gMKAOclISGehjHAJOjWl8fTS/Ift43QcAUIx1ibdh0CSMgs88PRkGwthx5Q6
TqAWhtxS8wyHJxgRj7akH+bU3NCJntwGiyreZM3ZW05pt3DyCzhC7bN4OwR5td3CpKgnT+bgy0ZI
rD2M2e00iEXuiAcJoXF9r+j/37HPYwY0j2sONdGGGCdud+L7nbZijNOXvrOhhw40pAN0G3G8X51Z
rYByMjvGLMTY7vDRBMVI7f0w6LQdRBlYyhHHt8TUxLlHN9DaJT0UgwdSi7mJdR5e6HG1CgFjmVlc
q7z7UvqO+xNMCfeRyijBlLAzVGWdIu/Sb84EH8DmDGSByM9Z4zz4GY/KxBW7gWjdxggTGgDxE7RP
cnDnR7UHYF1d8X6sdIUeN6a936O0ulDQpuuiYQyBippbfnthY+Wi7QF9yc1G8UGUTlut9uDOC6Gy
k0w8pTL01Rmo31ZOPKFc3HgqI9kvDsI3yeH72GBkeWiJK8N8dfbd+OGutoPFZkUPe9ykvDAeqwHQ
SssoPBtSCR8W8mgvOrVSHm4644OnpO6745g1olTbqIhU3sCVODRQipZWcPoDzjb+5Q9+iW2/yH/b
UrMk9lZTOfYUW3EAV68Sic3DrRuGy0ydfCGGkEzyFYoeRe4+F3b0/TjgVf21p2sX3neaEwQ7nNAp
ctFYMqk6xSt4JBvL0hPd4mWEXFztBETIl+Q8aCZspsnxvksVL4+IZq8aGXC+qNlDDDCgjLbgvrpg
soSBr39WFIsF/EKh0J/ue64NByeFOq2Hi4VYOYZk0pM05nUHjT67i7RvtcSqWAJrFLzh0TXvjtAf
p58i/4K0396QTFisv3A4yTv6HkDGSAhDfeBMJpPcZKq4nHXDkl4L6LGHgyAvUoNwpjOcWZ8ZmKcZ
SkwVGSOQbeKwpti8fPiTgQ8yfdA/kFloKX4Bix0A2eXQx4fIapnmvLOdxT0eU80bIEJNZmt4ZfbB
nXe4N6ERgQmVgbgqkT/dUPlxi9F0pai7XLJe2St39YzvzJVmX/Jn3pk0eU13WJ/3cfz+9c0BrGOM
FVORViUXCW3gKQLBoOUA7XxNodA7Zo9oxJvhvBnVMjeDxZqBb5FOO0Dggs04YXWJoexX9MrsU0vW
Zr55Ep/NzecnH0tu5/36RLZD9qE8cY3IoYwrcbBf8wS56+5ViWpeIWdvrB/q9Dax33Rp9TjluRqb
Ps52iDOUuLFqb82EbdH9yCXUGa8IjAaqAvbGmd7bWXZGgPiB7zuFZiEqvulkP6Bz6nUMjm9py9sc
yNgdfQNPJxkP8+zHjVEy62bTzDW47NBm+x+YBpYn5HtI/aaAtE+xQebyDQOeJSRlD5rfjglGwj/x
wLm1AkTt9vt2XMs7oBjk4IKDH9nIeRdbyxKiZBzYTawR8ifGJnXv5aUq42O0louPlnX5tzBD6MSW
/wFQtNI7OzBdASMqibuNq0+POMBiDQuwmY36S+tJTxGk1PuRdY9kw16zBEIVVxT7soECdCF/I3KB
mobqDz0j/Q3aAMS3e2QKmRdCgwSiDeWT7iY3XPa/zJyzxUhrrFIr1KSnCL01goxsc54RAuaJrZ94
TxC7PHlKwtld7pjEszanck4BNNL9oSbsp7qaDDPUVB/m6pTlXaXFb1oXpnZvoKlokU2jO6ChIkYT
AlwrPeKpUNBrKxlvSCOLcqQ8i8IhO4VXWwMnDC5w+zaWLoYOZudSa5wMc23W56jYQO9ysr8E2Reh
gF2gVBiREDRr2SSULp+vVdyVjVhG7nJPZmVdBeOXkB8+VYIfUcnaW9abe3NvFl7rfeVjS/dWBzhP
MHduHGB2r+x8ICNk/a5sEnTdl7eG4sp5S8vT13wnURV4ariUFR6XhLm/aKIBW01HaPrnhZuVX63Y
9W9GN/zo8ZdyPVvUuTh4Oc6y2OU9i8i4tYQKixE7WCsnvPSNteLCwTbopGpRx1g4vj1K4SjerZY8
dJJ4AZ31XOghtH7euSifJJZdkibiYMJMPcEFaVZ2Li1396vnmYpYByZp4rdGakld3NNqMfQEMqt2
bybiDhEbTlBuQkDqxHpxFgV60z4qIZyl3bpa9Ae1p08uBvDzFvlY9tdgcH6pgI5Fqejay+9FMQxU
d+MQsA/ea75sb7ukzwN+Ijr/f/b503TFJ903hC4hdIVASp7cls/bxZ8SEw7Zw94iVEpatrvCVmWz
Zxcz891xRvZMTGrntHi+STU5WHtmpJ/jp2vQraqMVjOxN3BTKPqQpsJMQyMzHVLUK6YktzrssWIG
BBcj4LTFibuGrttCryXuHEPdS7zEEuVJ5luiHCLCdPDf6ERlA3el8PC149j9/XAdQa7xQ4xJdwhF
1O7IhYRVxIi9OcqSKQynjEKKg+PmHvV4/HL+CwWFKFU/AoHlnntluyvNYIPokOaaKoiYmvlmE5GA
fYPZzBTjvrxLAikInH2OeuRgt/ExDRm3zZJVY2NuUC5ljfDZsXMBWxbRBst/bnxVlOq85Ivms7/u
CKXxD1vhXUjgzy2xmydGjn6Ym1tVlSZU4hzst7IzZPa0NG2Z/VvSlAq18idrzpX27RfR4WijrCvL
yht6+XnbjzNEYIMtGJUs3NqsRMQ/xukGiCkWfN1ytclB8KD6VQHoSQGBbuZ1zOLEJWhZJ/k+ZCPe
beVpdY0qpd1FtS6Hx99EGVZfAMTVPTFtYLPHZdQfUm0CRU+fTF5kmTOt5MHEETypAb/iYmmdBhjo
RtL61MhLlzrnAbe+0WRfd0mbukaAE3MX9isQ3BRK+5OzTwbTpE5NwPMP3xsip2Vajf0y2DGQLdQy
0CXwJrNcNR4fOgOp7yePER8veytttHx6Xio/3GDRIaBBwrjHCDQ2hBEcEk+rHir9tbaWmdPD00Zd
Fba6/OgkrEdyHvE6ksRJGvOVXsEKvbofo9NPBBS2/gqAj/rgHGqRt62y3b+tqoBp0yfw74kpQvMv
XmVjl7RRfO5rpQXVgL3TaH1qw8XIKSMBEzQWE/Wc/dm9iF9zkmKIO0RB/zhjVM1nZSORvq77JKWA
RQjUKTl9MgqjNxZ73CjjiNWxPtfrDOw1k6zPDPuoQ745jIbggfKrGVcDtGm+rW5uikN/Zb6lRppD
22bhLhwbrfiz8Ov+fSnMK8wIwnjbV6owgKeMRCwVYx9zFDa6MBjigH7v5OLhr9UpRX01RyAdb3rK
EA0b9bj1TWzXNwHacYPK19NXnnrcx6ErnHB7kF3EOMEt8iMTFDs5lB5gPb78chhwIHZqIQ7VvtrG
1oCADVy31Eni1DvK8etxQaEdpzLUxuVerBanbB3wtT0ezjNclrDgpuj0rCjLEfP5rCE0T5y7lQS6
wEKHywV6bl5k+KSrs6bs4SmIMuvZmDusFWd2k3ZqCLn+2wdgX9v0uo7i6m7DFPhBC4fM1FGkbcUc
iVojFvSePMI6S8mIabZhW/SLb5IF4IYbVYsf5DEWdiomfgTOkyQag4rMCyXaHo2aYGKE7aaao0uq
Tvvht0NLYIJKsDG9yNNV9MceGtQhHEtWUoAhYS+lFln7+7NB0RBv354kHvCGpsiezvntOj4fic3q
kQJXmsyp7d7rhUV56ZQMn1k80fqDqXeefZ3+Wkv6+KHZMBF+nPmLw6lLQbGVaEtoLq4hvXQEU75U
xov8YI8cvfVBXtxPNTD8DLDBKRE2GXB/Jm1GMtb9vvJjLSgXbbgkXNizcnKURc0q5jgr4e1KwcZ7
6tbez8Y5lxksZsYI0o9QzJXEQMSOkzhRQ/Isk+5zv8WriLsq2otxeay/KXPpTTlEX9u/zKtX4TXO
8rlhIex1DsfWIsQyabI8SBPB9/oU9J5zjd5jEQxal2gofYev4vqfr5oIEVMqeNxauDH5aVG1WQJS
+dudanvyoaDDQ0ybsYA9hJbdLXp7KP8k+olFYXjGJhPoussgb7wZcxTfo0D2PxdDO7RblcBKKQzw
Q9sax1gIz1IAjh5BD9WreQXSuPmQiuueCWoBA7665X8vBejhJu0MyeQXVlyomwBgRpZpIbI4KBKy
6W18AnAumOzUftwEVaR8I/H5wmZozUV929hmNaYwjSeXtchOy01BUxreBfu5uMfmHeKZdYVs3XTr
MSU442urJbcgngrg4JLH+RCmQ/yB8l8AsMKu8FsqtQAS4uFupMYQ7u2PuYZlHb/424/r6BSzcbY+
UcxhMF3Pajw6/FJTljuFQGE+s3M4kmtMGkJ5iLAQhmiDExQ/oNCYVVg9Sa9yN7HzLcM3z3GcZrBy
PY7GhBzJBCVwnGsBAQE6q6ZUrnQNmfhj3fe9uULZKLF3pexLceQW9vEpr38e5zZ9irSMTIU8NtVU
5wvrW0FK+dnYkDOviXVBkWucrX7APqoaWFtJ2Auvh5uQPfRQfAt8vZkJ3sXmjIDTVwKjkdMk2AVJ
3RcnF11SmUnUAUk0epBwWkBv/xorwgWLZyxSW+xBGbgLlU0q5tFmXj33U4n7aLy4d1lHTCmvNwu6
cYGHRGjwN1kbZGPk8ADRqDVlzXqzS6plXHUr58g8Lyzanr4rx8OdiFqducDyyYD15qk1teuGiXm4
7J9bR0fNiP71TMxqqjQtIn6usS9UrVQgVz/cMlFUK6AeR+UH1L7vK1nEI5PZO8FvdRHW88yS+D/+
6u2BxNS5VBxoK76oEd02enWbk4Qd2UA2KFFBIa5YnPVZF2OLwd30XCrlB0kY9UoOHAO2HnTr39Rm
xIakcmUwZLlgKyF0EFGxiPptZ/jbgjB2vMSZd8ZJO4KkN7oT1nEM1hlhg3K1XWO1IsjZ/fyJXDOF
GZ7Qd/Fix0mrmWPcqixkhtIGue4SjvXdThIFyuWAZ3uY+8j2X/nzMOPJxcPKeVTZpfxkmzBWJVFC
ZNL8rujBrSoWXJUG4ndDEycNd96YBNN7xGwRizdgZMF3uy4V8jPFLidZzOoXyIdxFn82pMFb/VZN
ZtN7BzWLhyfNlCGO3ByJLhmys7hyJeCaYxo1s0TGG+R1CF6BS/e4LBMZPss6I+VVkXg5QTMNnwpO
f9bXG9N0/l79c12nQrztzCx3psBd6VZKCTGwPDzooMKwmccPCanft72SYd7LGN4QmdVIo2pF1ypM
comSokewLQokcUQygoIHHOjPcg4A87rhAn15vhCLUKvfD10ey19e/4c5ryvdyEEorHSR3FX4ZXYb
cTZgmBxMzaTcsHdq3+v+WIaRCBIprUdHTvvglpmPhX4T9yMC0u8ZZ5AfHFsKahr9QPZrhqRs8wTj
uusc8ps2KU4fEs0SFh+65NJRBNut6mXj//JdF//yT6X20KVwy6MCG3QlTiN080FKLdGh1/HHWDMH
kD49qk6xlGgOBi3tkymxnnhmCkmqTJgPm2jtL1K/KNTAAg5GAZL+/559ZgoFBBfCNYNWIgIkA8Ed
qhRs4+FgxXB3e8qTn8vuqVr/4ihaRzXx/uEW4w5BMnwK5bNOKHefUaIH6KmzcRqX7IwleX13jPkT
bKV0LbWRC/Dvv98pAuvWBXQNDlzKdoEHpBudFC/gOUgavybvGgMc9XUigp3Y33JpdK7Bgr3WRRDW
dGnd5/j3U2UoqymS6wOr1bGgntSCecGLao3KPFwPHgDlTPXKpGIRQNdlUQrrJanFr5bKtGHZUoxu
q5q39WZWb9Fjdmtr8MY5sFTxxFCnthRyZQjq3F+wq0XAJP02a5sy6voImhBTZRmMLZwkSfYBm30+
lrqrJvftGuRX6cQc7Ro7b/e47FrisFC55TXtpZa3WaaoCHTLOYmxK5uIdorfRcnZtRcuEH14qUtj
qeh+VQSuXaFuCuIa01R1KjywFj9deZ8x/GykSqhLYndr/kqLKS0XiIG9iQ2fg6fweFNS2IlRrIGZ
aXHgnsAb9ZdtpM9zjROCwk06MfdyqeypWwwjXqhpu5tRFejTe+8pIQ8Jcv1IWyz+BiQDw7rIrTMa
BRZdrdSHq5QTrBMn9lD0MEYEE17LiDnvAcF+C1tsDe76HADB9fZOEmTjymLaA4UQS0noxvXlv0CV
G9l9QRCcq3DwEFbEPs3VRFHal1KyIZiz787z7LX0MSNA4phTyb2XqM1cmtAvkD7KZ9r4aMRTDN7m
AgQ37wz9VTcPNH52P0pqf4X5g9kJ6qoY/WqSyBxfoJoLu1loWTtyNjIleXbOPG2C1vDLI7fXEGmd
DeTd4r2fK1sURwt5oTbAzO+GHnoodUMUXJC4Fg1SbzGFh+98reQCXPMTKf6hk9uRCrcYrIIX3kgS
fkqLNbFlRv+3DB2gOnVeu0vSw0kqRfxA4XqDMDq3MHN9lynq4qaphitZCDPqkPjGx9z8V7V27NcS
zgn5cWTIPjRwixlxHYQFzJvEQB9RQrHezv6NtOId8V8KkQTALjKqfS/A5Y8uHdTs4TNMS7Zjoz3f
pFyUzYRiCTDbuRe3CIpxRnDX6EmaVaYErvhxFrVRKXEiAYxTC4Z2IXTBG/m/mlItd6QOXKTgoYoU
+/p0KDSeywsb3t6j4aagz1p0WoT1hx+R/KOWzW+mukJyA6SBwuXvxwU5VhN3GPEiGdK9uL+8T1OK
3DfVp1Nq2NVQdUFPTZXep7XWMXdT4tSRpP5isIppt9l6GgIflHl2UjKZvZGuH4jvRpwdLioTNOQi
4SKQUu30/Wt6XHETg8YvRxywykF9Z8QYWEQShrW9cCIdShpK9y5F5d4XObLMX+OycF/wRKfcl/6B
7vhAauvinJiPwY7MptXfJkJXeZK8eOsS4bKBCsWH470TEUHXGgnFQAUUPgi0EK8HFEfbTMKIZJ+9
qTEkfw4r0ZkINWEWHxrJWXj4FcW05H4BwqnK7T8bDTVhTgxwMYf8OBNVAJSs5e6jgPTni6xV9WoV
JqGlFrRv2wXl3gd7YA9ff1E20lPLTiYHHlCboACbmreSk6ABF1UaQmzQiNzt+e/eb4PtXP3QddYC
v47wFMNUILf07KCdROf7qym8xAd8CyGaudM/A+1VDRtj6OOETureR+6j8HbW49X3GkHBlBZTGrxD
XMEWa/h0h09+WpoVDAVpdEfEMBbIYUPMeKnT+2MBJE0XtIBhKe4hZmPbrXCNtArmtxkaOy+jNAsN
BR70P9D17NKkQdOup2QF/kOFYOhCoCZSEtvz0PuFaP555S2l3msah5n4+IOuxtCvjtfkDu3M4H7Y
0qh4rpiJvF7AvmzaNNuT4snz68y0uszVklHwQW/1MBJESUULQJw02gbU+eSsZPdribmOLgv/g/T/
ZE2MCsnGhmDU+x1p7URtnjIJWgx4mRIRnw0echwOByrFzVFw+eE6NJlEcWRSE6Phcxsbtkv0uMe0
kkqZxAeQCxV1ttO52qcYSCD+BXIxyXvkjzU0jxVlx7tX1lXhPokf2drvUwlvU94CrCvSY78QY2P3
liCbRndyNtiNbNNtfQFQnQ4JDijsUIkXzhudLs7o/No3RoEWYeuI6mAwBx0enpe0WXZK9smiF8bW
KsFPfqSVNsz3R2nzigxupyUVDhTJvHaHXu9bNxyBRAfO7sEI7pJ2+fW6NNyydSRCIgElkPD1vx0k
1c+HA8ROcknyc1PHtzqPLVfbr0cVuZBHtfEcG3hbrrUBUp2aaVTKIOiuzfBvPxxtiGV96ByWDaMC
XN29XVsbBvWy2YdAsY3GH66933zFykOtsiR5zLXEnxmFos5VIU7rxoxQFzvNiAkZFqbJPaRghdJv
XYHet8ZezgaQOAcrx1fTEJG40qQQKe3+6r0iRQq08wPt5IzLWx99yl2OZdgayeu/ecT4tTjHWPSw
th2VIsTn+uSYgn7ArE6LJcz4VJX3jHBjAfSZrNu+XACDZz5fw3bS81OKniZQgVzAeZYFAOxZ7Iyo
st5LgyZ4mMx9KMw4zLg9ME3fbsxcs39/wnrbYeVgmIjtjWbg5+aRKO3tylKSRAdTOLZXCP6shXsi
E/d4k2SrPTtFZQAsLDgpx9kokUCWEU3CsucawGbyASi87g5l25XKD4/viSrAnOApAgYka3gH+hZj
c8WA6va7CA3j09GRPdkzy/DME1EIp1w1kuwGkVwZHXaflGBybsaMDU3+Zj8U+S79CmPK9wtAO1Ll
stPG3RdpjpuYCTY9iialcvbobWpjQWACfl27F86zFIgmCsjUCCSh6CCDAnWJrgx30gg6Bv26x58+
1RJix0ReN1y0ozhKF4XgLXvkXbjN6FOrD/hRhOEVq47pAUHda2F5r0HGLw8AS2b8RDjX6qca3Skz
wjX0VbaCDF5NHRLK9y6E4wD5Nv26EOEhZjBu7hZTRQETz3jRRxK8dRCxpMT84+8ACiEkKmic5nc2
s6NL4f/NuxogtSo7qv1ezsCObJgq2828llk16RpPrEE3QmKja+VAEXLWdsEXzJ2MsVMr+5f8sgLt
eM8h6cnAAsc5illoU2xtqQhiHgQykQ8lAugvA0BsOkwTCR7+Fa49UbyoUfAC7tvWe/iBX6yRCn4q
JpbCjPZpd/nS00x3zWeADM8JwEO+30BKBkKxZrA6eSYGmWJQLb9up2gaRJuyqK9eFiaW7Gx2X2Bh
u/PGMr0qSIq2ViKqpmy34ieTxKo4JABG/YBKe8WMHV4xrBYimq54tXLYw1rZzdg3qczalog5kJmW
GZwEtUNQBec0+o0XtnkoMT7eHDH5adbrUDBUM3fH5c+tUrZ6TYcZUWTthVxkcGhAOGd5IpTndhzB
kc2XuSN/2PnIG5jRrcZaeqPn1gJjGtD+VWpk6bzTk/2kPpl323qYDRnb72LJKCGdbaeGR3+5lKye
PfhLdNTcqydVModCztdSlijkKRN3IUXBw7hwO64/lGoJQngqrUNanplmQERajqSUflrcY79ktOtv
uVF40OOR+RNcsMgNDCFgnD/fjvmNckCuA7QQ0E6MGh/fd9n9xeBFLVNdStMUWy3Mm6Oo8OVeqsz5
4wVGwQVkTiu7cYTKeEQhEGuQdDNZ9G8tM9ZubUeirxuODC33IoD7RCLyQBj0mIbs3p0T/OGkM7jS
HTtGyOfQoJYeVQgIfmI/+xufY6tpTYMKzTPikPcKr3zWVR8WrKR8SPZ3Ms852mUyliJBm4De24km
4aku7YZk+X4rx1iQDAiVM5KbJvqC05f+RxQERrwfj5PEbIieFgLMLZQ67XkvhefH4PumZCBqrAxV
H0MStQPOiIRk4CTxJgvnxZyMWzkirvM/os5AoTUlQMxxjLXbORUomua3GA3uQzTLknUHh43gcNvF
rNYXomM67K0xzYRRb/HMa9gAg3xohULjs57DvDBysIa4qrF/rEc3KmjydfIQ9PnYn5H2a0e0ZSZI
0Di005mPbuOy/xwAKn3Y1A8f5F5Ms9ExPvVbScxhiKBgKtH710VEhYK1vRbjl8oQnl1seKHeW02e
4n5/cZxILlgx+WkTnx126YTndFGQjF0O1guj0mg5hYOGWCq/hENKZwclgiRw9p4e3OI6VPzjR8up
8kqXnt6codMMHUAQpgruDGz9WOMGJwpwGnPybC0dzQ/njNe56FfvdBQi+Iapmlp2iVksnFOa/kxj
qmwKunTeZ+29HaCtR2soI7E7pfzx3zcRgHks/fOXZoYCEHy+aCdiXBENoPCBz60x46sUOQUDQ/JR
O0msz4aPGzSGXI0c4xS7Tj1WlYmJnmm548azWBGJLYnEfaeIpwUef1lsfEzbnJRmLcP5OTsrek4Q
e+HScvkrPCWZP5jHWJhEPB1yEtT68rm38Sdnngyj0Vq5hrnYEvQQlydwyFNKdNbqplSJ8qsYH7VN
ydgiaUP+jeCRvYbv++RAOv7zIkGr2Ms5de3+esgveNG+kkHd73WeHNjk3dcDb6BgFKxuYquwYnL0
x+0dXv38Pq/E8h6nwCQfcETl3vrS47nWWjc5cG6L7bAHvGzAaEHSpJM6YHYzeIgIc7cIl/xKBD4F
fSYP1RnjeBXWDzTyYi9jhJu7sajLKEFuRekV4ZdN8pChOOV95k5y1qKbJLagwfdbKps+Ax+O75vf
3ia4oXQXWxdp71wStqR4/1/hxRNfNIiNZzYp0hJE5HBxrfv/EIII5jscoysMHN9mV+l2CzE2I7WC
KJCv2Qy/TlA8PtzjWtomPeOMWMWUkhr0mxpIK5EmTZMHdu4qRtLHxln623c4qRlF4sKH4OzENq39
U7h8N1xDu6LnNzNEVMRo8/1jT6ZaZ5s/269l0b+LBRKrQ1rC60c4yV8fmgas+5b4qvKkO/90gASS
buOTYEboPqeY7eu5oKe+a6pIZxZzHKa8Vds21gj25fGoNglKCmkhPQ9BoycyzcPB+9nd5fvFLAp4
oNrRObWzUeltKG2ok4BLPX7FHUqUTZLYBEwm6H/ZyU3KyAPZxi8ovPsQjJAazIVdgcTxCv59zYOt
eSDOoSYdAGWXyEzOzJBxEmj4SWezMuXgHr2d90BQbUg1HnWWcvoKQbVHOvpW6xHMvhrr8rjnPlHn
tAyxHKBANDMQ1x1V2NfYRVG4+rlAV1POpW5/YKUlbjjgASzbiNiF8HPU44hRWkbH8YjX1wMpS98x
1G3O28kQrSSK9avgnHlxfLfDGRPp56U6eEtNd+nT49Z8pzDgtQW1aAcQeB1MIUxoKGS5KiGZTqy6
5n4/gY2Z+CqH8iv2A5xAbn68FkyYFz85W3CjBbA7Yc+9mVJ3srHXdcwu7h/Ibrub9dE8KLy+GjRc
l1g0eJj8JiN6kr7doa9P7EqMTRtZ8b9Mb6jBaY3l3hahyCAmVrtOcp5OOO/DgOeUzp+BEKYcv2jq
vyumf9oaFwfRwigaM1BvlguJhxI7JSHDmaVBBnw7SjQ6rLKudrnbxoemjKQ0URekzHlcQBeSGiMM
hMIOhmrNYw6aZwnO+E/RAsZg/UrHrPmz29Wtt22aHRldX3Z5e2YrVx6YNSiuIu+7bhRs0BooOBN4
aw3V2ncL+ALo1TeKrszdUm/1VhKUihzSfF4lKy2yZpHDPEAmg303opgdVijTT95Sor9VNJMm1Lgk
4S+k+KWgdyzBop2ULrpImdul+UnphQOFj2mgEneyp+TYOMKNyvhygHjHT8FjIJUjRZNc46zFgz5Q
cDDgJSsGdDRbwMVV8d37EYS0iEgZsMeQyfLMx8Y+CvtqREdQeLuBW89LxFx2/0Y8/PaLdKSwt4x7
NB0hg7FpXOMCgfdSHPgiT2VapuKAdGG8/nwFWYRHY+nbGTvPBBBB5KqB+Wi/srTszx5+4qhTv+Kx
BUAy1lOAf/tlYoO2ghMYLfncHlNx30EC5ugWvlC4JRqMbMelNcErkZlmTN2zTibdsjbUGPj4Xrng
Z4goNpCkAPNQNUVZUS+LF0tqiJwnMGpV4LRGn8xHE2XCMXET9hvVvZuj6OEToaFWQsU0BzRIceS5
QeM5tfuukFFl5Qy6BAnljokx5JuHXK1WZLvOOn1Lx7RmJx7AlDzkPCenORnD0BVidE3WVR7YGLKq
FYRfBQRhNz0cEB+RjbWKCnaDXKI7dNXREzqzh/siny7aI8H44XdOsxHvYgOhbQstDCAMuBLqfnaa
WUHV6TUCg/E94MelrkIWFQVci/maoV/rkO0DMwFxlv40UwpmXoIbzDSL+cyTnFb1PAwmFlvthTOf
Gndce8netaka3+IzTOpf4uwGP6KbQhdl2ANaBCucNnhjdc+eS7xpXgQk/0T+1RCElzGf7N8FSLd+
7Q4+X7NiphJKgKnQapuGaOtQVwrp5vyQDe+NBFlwvPjfKJWmoYy210A2ePhKpPK076dKc74RhsYq
FGua4cnM5hxYJwMqrdA+CZdK7RtIXKO8zYSyh7w1lmu9jrZdU2jBXUFedyg38MxAdv4aHSBqOOP9
nDM/bWjStRpvvWWx3Nil4gKCX5ZrmhHAOyCPmOR4Bso7EfBkhhTcsxVBwkDor4ozJFjcbuIOXI/l
lM9IeOX6GhcICc8FKXUS1RZzh4X5FaHl8wAJ/9bZYzru5GTMYOTEn8I30RQYD3S/G46t48mkqroV
AJzfxsF3Vi4DnrBN+rb2lAUAAw1ZNR6j1PO13tjFi/qNKrRQ5uY542Kjz2O06tCOt3N7s9qHK9OL
ZEVdPg9r6FgCVG84kyV1KdZCI64DIj7Vm0NY3LAEkJKDB0NmQAdb4bg2agCTNjtPfnDdru8h7FpR
K1PUERzJcug/8POntQdMKVy3RFjGACyp3nO7UMREDEJilJOcXYC1lYF6Hl2ws0MxFASgmnXLNi5x
0uXc0edA3ZYTcdeR0HEgxay6YG4AXArU3uKzvfHMjr+QGcImsPgQP0n0GKrd0meeMXPV9zSnNzbO
S1PhmO+7+EdEv7aT40if1QfW/S39u7bjLo63e4f/Qm1b2bHlfmB2tPufIBcITVINSRx5DnnIVB2A
6jtQd/EvTTC3rDSE08LapaaKCtQspoueh+nKOFzAh2LkZWtxTGxjxBFIf3ofFdPetWMVWKnHFqT0
RraZ2Wr/1Ry2QVyu+8RyGZmHpmyW0zGOGQ9jflZP0lQzDek7BX7WUxedJ3FCqyl5XekmDNFU4C22
RtWzo2KM0a+a4/h7X+Zy02k0Adzet5HRgqIpGNpUmeHGrMSF5jl7CYCz661vZ61SeyqX3Y6S5DVD
oXwOhwzEnMG9CNfacuXSR5uhCeI2kL7wpEARxuEwnmQSwWaCBgjWS/VpXfmj/4yq7kEvS9SuRV9d
iXHKtlicl2bnZTXB3LfLqQsdo6rnBg3AH3JIoifnVkEvTGceua1Qagxqmq7rZ1QnxKya88HACR1s
pywG+Rcjq7yql9pd1YJx7Im+7xux56ORFcSD5XrqxFaKZCev7Wjp8UnrgmkCpcghNIeCp/gO2+rn
Rfb1o0z0q/YHYzDVy7MuCJ7H9VMdghxxWH02LcAIhsYo9trFLWbPs3ChzYXp/R8CHbt4FMyoqMKv
21cUZ8R0vEfKlewNgAprEACjNmNPx7/pVVwWQ1E5vA8MGn+IffrXrcfZdsK1/zrFT9EfxLNLU0SB
voUImYvWWfiXK8JT76/HWY6eL83tSPaqfGv2Fg4ntobPmtJ+DpjzX2vbyLO3yuBzYyyF0z/Lsw1O
xfXent8LcWsKLhJnwQz5SGamT6LbuqjPQ5KIDNC5z5O8FMwMYgmIFOyA2UKcZ4WCFX3+h6eoMPtT
xo9dct+Wn34lSBqPELx8ZHN2+wmwtfjNh9OCQ14dlU/D+EB7t8qhgT7XOYGa3SDKS3rIVsXNtGDv
l4XWgrt2ZiLBxnWS2ePnC1an5xcTv2Yh/J5orK2P7ZZqVbGSQNA+uh6Nj1zyFfeyLeBGDn9xx2Vm
N0rYq73+/umtYDBB8tFOIvkstTzaPsIC552TTIOkHOnqGdPkrrS8TvIaftLFwvoTzSa7yYkNuPfy
jP78lr9DeMgg3ya5Gh0nCnaFDmqXmn3AgGezbbQqhcqOD4dwF3o3xiwAQQmUpWiIP7HfSEDWSK9h
idTdrZxFMSSfKnNrOGw5N9k+2VGscX8TDZgh5P/tdE7+AQfSuZGEpgxxGG8O8ryzJPGDDATkNQMC
4FLgRwWePG8oGqWhmbO8C9JIQXIybyijUUdc4Z478XJEJKC7K4+IHdEO0A1vMACEQi1vXEWtchYI
dk+lzkcotP22Td+ajHJ1Adb/9Auevhsg3Uer8n+Q9052DvvrYJLZ3v82Fyz7kJvwFYSYvpuziZIc
p+S7Qa0eGqkx08juAxajRsZfIMVtBwjgQ7cdjESEwJ0ykiVwQLD9kaB5LfiN7dp/NqLSDDihkxeh
3cSM88U7Y4Dr/LVizCNG2icdbSi30n2DHwN+x8ck8ZoTsxFt9NhLSShy6r0Q9hbaPXWKC7v1J+mV
xFngEuSq1RbuOurLGXSOIP5W7par1t5FO7oL/Op6/wnYteF2jPPByeJ4jjZTHxAVlSinqZmwV8Cw
c5frWL3dRQWyQZ3NG1OX1XmmAc4TsRQJtkJgJSZcHV9QqGIgbQCFxXpWDJWdPTuLgweeuEzzLzvv
mNNtWHdgC0wv4BNxk9yHr2tXV2FZmFmDhTEm9m4fAtDJSap9ZXa6HTnwOe2eInwJfyETwbhrjKZq
BKBM8zv2bQcku77WXHZw4YVQwY1GMjgnyPJ5xWayaOIst8xtuBsuRBOsqBm+qvZx9mtW1lRxRuig
vteJ9w6cPboe0F8CiGRkfePJWCHXTpnu0Xs3izSLD71EzcA2l0X313Z+FT7C9IPcTenxIkTbKsZQ
Y37eTvimyCJIHuGliNjen6WHwXz7JzEHPeTO6qkR4kJ/ZgoYOicdiqBoBXnI1fNOtuvOrjo29dB+
rTDUZCTKF347P5O1MPW9xQG9PsOqx75T7DfDZDVUnIhR4FSLSdj565CajR3qYQOcKsGI9DlrUoFZ
apQ+mr/tDFyJKb8oZiaT0PXdL/8p8IMq+zYsVRdOGvCo5aCagDvulgDzRnNA2aZw9vMgj7ZZcY/V
6E5kAfrRtP4YOyYgVb2oy5ZYWCswBmJJ0zbp2oAredCDVTnRcE7cW9dqDcr4HTBB15raiqmhY1KG
5E5lGJtkiOnkaarAYFHDCy/nUpx+x8TpsPXKtXHdWeQ+aULlIJLjIvxYd8XG/tRjqUJqQ0RrBSlO
HyrlZD+UBLjt1CbwyalQf/rBlJut0JLBx1OSGAbrkaAv/YXzNh7nAWaMrdjvQcVyanHl4gWfoYWZ
rxkWQjav/P+xqvuA1Y+HDNr8rlvfOIHiIoGPVGshLoBwWvJwdsVokrHb5SjDekKzs/IW0twnss8e
MWl3dcID6wVHCPMsOU3tYgzSJ/IhK0QNV8EnUrdZ5AWxDGq7koKq5ZKdMOln1WC6PFOfTsLuccIf
60dZz6Wl/ecBZWGd3Qvb66GyrDZ2l5XrITQo65jqIaF99KDu3DuL6iodXYRm0YGiTgiSwLg2ZVL0
tsBgLxL6ikKqY0ATPNdt/2NX0I5yKExAw21XYDwxc2nLTQFzXcQUZvBIejzl5m+qc8+4vGJsOgGR
FLdoL7KFPH1TcS88v6LssZ4StMC5a55MMNX6XLciooJhk9CvyxJIvIgHWVAUBre4Snyww115goWj
xfUvMpJPdXGOD49ml8Z30oQQOO6L21rwAD0i/urIpRZHy5dKx4pVJmCkxzTakxtD66SjboeveUXp
D1PA1pDenu2+NNdGUfp2zG04Ydsd2a72Wju6cnlCDNc+fGsIq6sSWUn4wy7wBaE6gvMMcWdxJ/kL
In4CQ4CX3/HGrMIQqvqQ4vGzBfeb0azMRkTXoR1w5Ni3KFwTa6N6vo07fcYAG2vToPqigI7WkL5d
XECt+a259vTj+dPeZiqDW8VglaoMU8JEFjWZ+S+/0NcTDpgruxvQ8fVKUzIK4ctw6MHDOcm2nwwb
KtpdVm4fv1YL17tmHMnH/24Z6slsifcoj9IG+rfbZLqjDsVnlNmwIsyOj6e7nmZVXMhVjEwTEyK6
w3gCLm2TMF9sqYKWHQY2tJAfxCgs77wqPYVZsSq5idY5o+G+P34ABH6jVCK5GRWl7HebQBarEGjM
rMwFlHiPtRRJ72sPKTkKp2j1FkXF366MEqO5YRfkz48uOFxCj55nfWAPPA2mzqWmZfIL0so9FEb7
e/I/3YuEZN6DBbFLLBJFAEz3JSDF2QL4cdgSruRn40Zny6RUxTdVK/GYapiFSV+0ms8nbNsgkQ5E
t/W2HCuGaChNPj4MEZOrzxmx575DftF/wFo6bgPYlS4z8ni8gEf6+zZSierULhYGdjWbevNhjgEZ
ZdgVxrM1lgnxRyXwKlDkpEPC2f/e9ZVA3GQdhbPpUl0YUEI7DyAke/ZnSMzU/8m2oEyYtJoW6xEA
UhVZ6LVcD3fL7WSFScg8CFZSQBOQ4nl2FALhNzH0cK0+6o/wIT3iLydMsGWZN8XKSqN0ArsOKCE0
l2kOoGj2d9EBVTD+Mu/+BvG9FH5IZcDNx3Niqilip4lNweuIo1qHfAzxVZ8rX39MIg+J2/1BgfSI
xg8y6ejvmA+k4NHP48CrgUJECA1UbzOSMor5RwaabaUyWltIFyjSaos4FIAehVnjU6/t0ASTkzeC
dSqjlJVH1/gAkr8gMqaF3tukKmZIRBuFA66AIJNDdDV9u8KrKr1N4SVLjcvVaGNjDr6jq6Q5b76/
XK9sIZpFgCkDy+0hZd7x3N7zsqYX7ZkzhI0knj+zjaPOUeCNe8SfJasWUA99yFgh+dP5vi/Eyhom
sJmtV3FETEEC6cCTiZBu+H6xtA+9SwroKdVeKYmWX/Z4TE0t2S20N9NE86yBCXCHtPLa2J/6Y50p
SG+ZRvFtYvCAkXgqb5j624zgH6e1TmTbiP4ljIiYoQaxLlSwV8Z4J/p4dQUJk1XQ7HF8cD/w8eJd
x7/lXNeyYy67IpcDLHFQ43yzNAKZSmZa/6BMi6MaHLHlryJ9XCT+J4p2DP7NvE4nBJxbObSJ9CnR
m378V8LNQPIWyGfYyUp2u89TZudON+JhjLFJW78fKSQKgvrpjOEyalz/pFWYia871sn7vKxxjV/d
h7S7vq/uy45kYq5RVSD4KVjx/GnWh9rOQ42K1TgR89EY7WgyDlMgJqgvmpd+7N8celhpkncM3ExW
0CtW48YD0TPOblB9Ah3jq82sCNFFHwrnB5NrAtQiE+KFFgkzXflzKaVQ6K/h9smqN72vzXzSCz6R
utoOlnHichVux992RopxJ6+OzEL/OZbxtAxyGHlNzk926KUd5ZKj8Rxv30+nK/HpPqhP4t6ouKv+
d/rqdK9rZoXdRlNL90z6XB6cjaa/8p3mwYXnDEb7uJxGoMIWJ6igVTyOAlHjnDHTo5Mn5d2S2Rtg
MZpazbsCG/S3MPx2EFIWD3iwViXJ4BNO+16keYcZJLkP6atzWeWILKTGHsC4uGpTpRWlMPz1OKZs
l0ohDERzos8C+btt+1Fw9O3j2ol+Db19s1xRRE0eoBfgsZdG9zk2afYStE+bRc1wwSOxW/sPnEsp
9ah0p5RFVdmd48zBh1sN9Grop3G5dP+0A3IT0nTtmT2KbgFSGmtUXFZ3Wtys32xNQ1oTg8mSe90m
VkyMoQjoOkbUJ28nvxSBhBx07GOZz9/kUhmdcDYjRVkCYquNNSGfkgICy2AEaHqEAJd7zSeBIVNi
cEqfJzfDa0K6D/+unVor0Db0EvjcUPxETfvxVQO2nE6kPMrMYLS4T39ZwVkGTd0ZAJjCVbW4GbPe
FEziFJj0YzU94BM2kwqhVldUXwZQm2RY7rG/TrDxP4kH6bMbkXYkiYbMyrWedU2dtYmqxJJRvyTi
IbmTiSioWKMpem0fE6MVCuEpEZAS+QrSRWRgPPagEua3bKenP0Z1Au06DY3L13YMmCZgoaO2h9mn
LDBUxIBgSClT38Jn8fdp5MWuvRFu2FarvYnw3UIDhE7j4tiAoAG9y7+5MX5IXzwc2wsrkogiKVC8
556GqotRaAX2Wo96CUxWf2ejM0G2hgox/4auzDX9S4sNJUodkjTSUtJ32kJsnLKZxt/irUd7eq5J
4VNCWcjz6EnhFSJAoar7B/eI+G8e5F8XTxBt3FrPfZAFPO6/3Tn9j9toC1FHTVNIW4EW8PIwUnkW
uTPtBTN7/dKfDHRR+lr7LCImtl30dtsllhxhCdxOrqDa/dFUKSMoaFQN6ji9I7M4VMm8eb/tLBFO
ymgex18Yy+267luZVbORyoxpZDCDC61ipwbNkuNNbiE7FlZNErO/C+nCLmlhCAybTAQ22cGQfCF5
i1JiBYOUkEdwhmfKVPg9yTNsJFvaRrBO1qlD/z68oWqZD3hzuLqPbwPd+k+Yuofnn1Y2sKvIOb/G
cyEzJ72DmXipR4h9Zvy9h2/0S9S7oCGD4Oc/f77/XQ33UTerCdqiDA68BToKfJqdkeYw+k0VODRY
wrS9iziN5nPlmNDgAEdiDAxW6DDQ+u0+sIeZLxJyinHDqR1gKlMfx3Z/TvZhCZF2LQWCWF4lmVE1
nL7BU9+mMKBNkhf07U1/GPDkTHn62eyNLSlmAJP8XM5vXa0YAdMAV5OU4KnXUx5d11gle8DTmfI0
owFFErgk6Avp3XCtipLJb2NfNkXpI+uKkK+go437V0silFIBPypYFREvBXFBFqlRuDFBQaHabcai
EL5KUPcg260FeEbThpeRwaYhmp80CYihm1kCfHumMwRMXNB/BzjvGThTpF6ZHQfdudMNI9eyaEVA
m4t66khx5I0eFFk6h0lHXAoP9CYnLwSMVjwN7dq9ldUF2+p7rYdrU7o6yRxDx+mCp4XRh0xmzs01
ZuEqy2qmMe617/gyza5vnXLg53JYb8aoAvWuAi0W8gP3D3sYVkNqyFnfHWE7NY+QURsGtGrR3Q96
h+XvWfMObm0Jd9DfgHkKJcOefDT2wX03t1CyHD4smDmxc/ujcExr6ELHF6OmrrjYCs6x3UrTInCV
/yVjVj7773i+GHbDQi10lGGmpBEA+wEoCodAZgc3ExBAy5GaA/QTNol9PdJ4qay1LOhmXfmFwc40
NVoZJPxLWrTZTOjDHpmWHgmv3dFqOvQgioC6mEZKVXL96yx7Wd/fw9UH3Wk5HP8v9e3A5aveS56S
QgfigJyxA0+3b705QmluC9ajJyhw6kTm7iC5prkZZOjnUbnEubMFlGHpM1CkqhDbpPuYF5Bnuaph
ZRD1vynkAeQaGZkRA+cMx8wNOe55biyb9aBgx5bGDewJIV+nahTysGAMiLzSYElTuAjY55I8s2oC
qksU/t+j2hW7/NPGDn4C1X+aE60oRaHbnubhKWEa6msid9Z0LtGrzT+d1aG0pXWygMbwW0P3io0B
T/oRS5x6j3xycLwNhxWSeucxjwBDo9u75BmypVrM+iEoLGgD+/K9QupTrz472jJbudC+WquFLcjF
WPp2flawNrkrkAKz5vcT09zvVUwsTUR+WiZt+63tHllw+RAXfCbidl++ZIDoxTOSRe7qs3JmGhvZ
HHp9f3lP6r9nnPIm+BrGQJy8kTGOqHznBU4ZMRoyD1gFLHmnOZN8E02PlmoX1ifhyEkX+lGD4+V1
1PCOHRjlKzKsq7NNHX7E5d0qiH9nGwY8mzOr/UQP7/4fxJKwMYgk8sUdsmHRjzV9dFMMOsdgSc1o
FXl7dH4AKTNZd5t2AI6tfgZ296eOGQmMIqXQa5Bv5BBF/tXC4YYmfqBh+p8/YUA8NivxDBYSuHhK
WAU75PFZz58ugMoV6aj9oEHJRqwI+83hK12TTUZdGvStKzyHhqXmGNbgQpQf7Q1VNxX2TMm0yJU0
TT3u6uKAd8rgf3ATEawT/r4f0HYAu0OsoV0krP30zUi8IBlKCyhjsZNT4YViQEDEVL4Y9rHJdHye
e6XA66rVvfVlB8fgvvYGzWlT8KCQpQYV0b/IRQPS2S/RtnupWdiUn6NlFsCT7f9NGfdWr0Pi/tsA
7edo9ALlLCx4yv9IEBVuIdszhnrinXXTtpiZEnapJELfmOwnIKQhuFz/fEXdo8BiSVIoCHsM3KwZ
AewzGrMUMeG8jX1r7Wh/uOJND2/wAbJrEfV7piLi63NTOuSvWGR7iZxHwuhy6eM6scft5fMMi72b
MXqcZUkpaKtJ1Or/VaXdGNkPhLi1ZbVOobD/AS4n4/JMjxS7u4gvwm+KiU0ebI3XuZ5ISVKxon6Y
clXmwYPZpzJFqfMzNl4x2UkcilSM9oPwx4u3UK1Mm6Fb+VOBtpyl3zYly155wZgg7FxRFQtV60v6
rEH2OQ5T9aIzdkEU1un1eXIgjoih5oUJveLtVfjePrKcIiKO0fwULNEEKkgzvayPfx6EP0l1D6CZ
SOd6wSDrMUrioRwAdMLqZIZfQ/yEbBrCRrByZCmSzVfZ3cV6+wZT51wJC3znbYzzrfJ/wuy2uq1Y
DjOlS+B87qdLJZk0Mbnpglnv4BbzudX4ar+0nLhjrKorWn6LM3n4ckMKHxoJaF99Vf+hrTufJ3MA
fHtlKf4jWFTye0jeWqM3YLv+LMekbpLzgMqjr33A1xeBZ7qwJy+lBtl6pEyD/5aEoq4lvlW1TWnx
rG6h2VYVVb81yG9WE+XO9uIonLIpDNG+jp9nAHWejQVSHw7TJkcvvaf6oh6gQXE1PFfiGOtPHtxT
KqpTKnGH4dcvJDig9bMl9CM/XkKNKHiM4IpYHJJL2rsEYNT11cdj54v6plxdW6S+0JZnJfpwnP/8
QK6WUHgKsI/kwFLvjH5WTahXtjt6nPVmitV/YuXeZgf8qpWcw4eXAwhx3AnBEd7Dszor6yvNmymY
GwEHTa/BifFVrgyVvqr0zRIaWPcS/23cLGKEx8UOmpeXfiy7rv9MeE4VpFDcrL6h2RWiXjwS6P4v
YlXJ4TslbAVm4ORjY1lCnLiOBMgjDaZhbbJZyGALQdSd1ydjYyRAMeYTno3sTkY9PR7RBPdnUYK1
B8ECHBS2n+W4VGyld+EnLxrVQWJ9ETkMuBjn7zgtG7RKaUEqOZgZdOJ5bynBhAuwpBuaxXPjwf9R
jmYgqznaJvoDAU3/NGvGQiO/eXNur4p35wesBA9lusjt6vwkS21lpatRj3ofFjbKrdz6W5EvCa0n
Njb6qeuHxly15YuuGyoL/jxNeYah6e1EvWnI/sKqSE9pzfldQXCNPlQbz94g/z0KjnYwNSGUZPbx
goJV+CmcqBqoFxAJcQReoONoOl+La2zMCMhp1nRc9cXVkF2An7TTDi4QkmVCgz0SY7AjfNuM53FZ
wqC9rAd12rfsgkrZJl0e0Mn1mLUDrJOr0f1PvLb6NtArQc7biy+RY1ac9jrHQmRxx3LLSWOxOI+Q
hIr+yVZ3MEEZsg61sGEht0HNlrIMRG5NeBxh/wbtSBUfex4i/Okof9hQUxoHFM+8DIy7gOYRLhPi
TjByJI8Psk6weV76K4SLpbWwp4m3ksI5ZrfXJvj9wsGlIJKiLpjb+LOpn8cgMz77HCadNUAevcCK
QTb0P0u670N2zJbpMWyPjEzKQZpXJWizzF0tQNxrwKB0V7UAHPWr6VEw/B9kT/UwEi4IJLicQ9LI
ypU3QLHRFBjiayB/ZyjbF8rcDDEGsyNjk6DlTtK/k+I3+cuM6j9fX5bgQMsV6LLwO5ld7x8pi3f/
PIKIaHytQO3os/7lyhKSVPSu48e+jEpbfNgpxiDHRfos08XjOw1Wu7D6hZNXaozIWr7xgCeM9mcU
331onMniUw0/8st1MgE9cuPbBiuiP+HwEBzcD2TKnwOq9cOJkuO27AJRGEEBczTi2fmZVplyaEja
N8Uc+ktRTRImW3VPDSiTTbC5pTn4cGIuZ1mNCTQXzS3CvH4eEiAhMPDMWKTfRpgvGR7qIbVd58MR
5Zkff+55DbPQKIIBiit9Yp2rmhZgUmzb6biUd8hBxVQrVRzvWTEtMt0UOFCUPqhjyQD1TV9DvGb8
EDtJAqiQNi2p7kZLYY3cb6mU4W8QMbDbLc+LiRMXff9rWXfGhHnF53vpYHmIoEc1//C5KJ0MOl+k
ri33eCpBck6HApsCVbJt7/Yi8/spbWIJZCZ4IJw2GuTGuhL4wYg/1l9vHBpDaQXNW2xffaEToJ/G
VCnyyEtev9GMxpWPDjXd7zke5ptCTIrPaw/XIRH1QM0f1RvrYSzziIXyZxuGbFmeP2Ok1ghQ96N8
HDFevpOJEw53OUr5mTVlcXy1IzC5GfPNE7ibzzYwYMPjbiesiLgEAGkCdlaU0AyuXdKcVmiCkrg9
lQArU/7dg8pyz+ESZrScH39lwvlI45Zb9bS6tORTS7F0UNKQ5PDSYKWDHGupOnkU1ap8I1RFL7Rx
O8P2tcsnN7JRd5s3RvpfvDJ0kD2GU+7tzhdZ4z2bCFuEB6v6IMn8aAcHRpk7YllRQf6OZgaCie8B
YOfnmpQx1dyuiMX4/vO+kGAlXxRp6K7nNSOUHvhczbbPAwoLLzcOX5RgWZP8ulIoCkUBfjbA+e6d
TFwX5GV+dbZZiZAeRPWCe2lcobHnsrSp1QWahwKxu1hehbo4HP8kEO1dF6bPAXDT2Iz7eRpHBNsE
uWr5FifVMYnUwWxB8uVOmYkwgzLQHoYCmopRM9go3S/4PTjp0/Slw32Cx7IggMyWD7GRgWUhmTNG
sbrX43dGDlfJpUDzlHIonxbLFYiOsDL9GpLlJjYx6P+OdCXa/p8bQ/JSp4sVAZDi1A1E3XVwo6kV
bmkWOHI3rWsG7h6YT1BsUF0J9woXqLm6a4Eny9OAMsGnazjBzK089vfw2DhWc+YEV7KEoMNJF/YI
EYBGVPm/8bnnkRCEn2Tf9WBSwXepAKt5KcekXrHi4O2tKUzF00VACfZiWiBgpmGFwnbxE/JTYeKo
8Kqxecq/yD3FXedgukGG9ccXdG0+I+M+GPTUNL9xtDVQbaUxqBYsO1T1oPHHrxF2OMIfgjzSt3aP
eEsgqFATlAixZMrT9mBta0xiYbsNoAPVCdnvIjp79tPAu+rAxTg5N8LLkOLGf7zn0n4bQAJKW1eZ
ggNtwOzS2JRXUMOTFtYv4Pkkpq/j2CkAv7ZE3iGfNIOOR/DImaHRyLhTDuJ/ZNsnAFKlkZBjBwEZ
CHxcjmGgqBUoVH9H5kfU71u86bv41GFAoqqdvMxBYwFL4g5PCpFrlM0Ix1CE5mkb+7bcqOOpe7m1
ZV5XybeB/N3Q42DR54otuMdCoAYR6YkN8w/n+Sr8kG1klHwJUnmhJYNn7bY6Gkae31tAcdVNgGWD
7mfrV7r8ce4XXSlcVSWU3ox/z0umtL9FJH+Z2gOFRayglNfNb9o8HYJVJ7Gf8sRKLHGkNu+KbowF
HkvaAZFnfKtrCW7Hdiab+UnktXAZasQVfYBu+oIY/x+senLhwm73tMcVT4TcnrXe9swATn5iqIsB
F4+HMRvyRSqceVsn5uCYd8OtQeNJ17nwaAcr4ZCpRBNMQ59TXqjsZvSAvSCdNqFSkGKHqR/Scw6i
nLn1qONTYOOV7/dABXhp8c197KzxcNOIXY3aQqDg7U4D8E7e7GTDdtcOdcznsU9q5EsFI4imegPs
zvNXJyQmadc/gk+oumwIclQys1UnLUUp8SjMkXXCKgQaPbPW0ueYAt/+DT/sGUKdyzAZ2JtB2/2b
tw47dfjEnF04fjxz/bDqnOPQq04KE+TDHcLPTdTKJxlIlF02MW9pMJKkjMR1r+hDiVqSPmeVr9gn
bHAGPHFBEpLEHjI4oEBW3w5xqOR525QNGw//ExG9r0m6FqBPw6MXTUCntcuikZU081L2MIBeG3of
c0y6YB+Wtn4EVkdSkNZloXY6j6690Rl2bGQFBuncSEttWRXdEv/QhPRhrOBs+x/ixxb39R/ogE/p
jH/c4XI1z/U/8q9RAgWUjHc4ENpSab7Yg26KjHBeJf2r7jdA0yQQCk1lbByNJrTYUSYbk1LtKUqP
aF4vt5opNp2q8TrjHXmnm9iJl8cBWGzSLlF6Fd9C/kSWqDdrXRZbJ2WAPHVmD1eGG+XyzH/wekMw
TvnaJnbsKPeG0aNvjFCzkldPPhwu3arw9nqTU7aNKxwBN/CfN3X0qmSNwJvHBWlU3wryfUhCMfgV
t7jLZLIFIioVG2B617zf0e8nPurrdauBD/bC9WfoVvc1Hv/kV0WKqoaRVffSVH26CeC280ln3KWx
COrFVnBqQRaxxw9oqzZ6BO+gQLFPyfRfaNR9GVpWiLSW9sJ/WeuktkqllPe6m+6TncBCwHVgdiwH
mMDLTr/W6rhvwMJ6Gsm0E4Xmrffus0DAPx3a/42nqQyGrFagRPPpAW11yxyJCrX8VecggGxV1uKi
gMQTKCtK+WjnXvQ1iMWTc56nEZm+S1lgIuZdYNxq4J2b9e7eKMjCpTnRNhCSUkxMVwtrGRwhwfDd
Y9ucCY2JxAeKsj2u0Md4LiYLMr/j1VhaYAAaJc5jg9qS15KdP4N7VUKRftKT5rFjHJc/ig4M4zK4
Ire9FYX5yf2s35U+btKbJkLUzM51L0FZAWPBwtcvG62WrkEZXHU59j2Kev+kPVolZ9tcZ06WORlg
hoLKMtkfLXZ0Fotw4lD0uSd8WNbjRDo3h2WmEvLatrM6+mmxALXk9KYYLc6KWnMhEi4j+AghZJ2c
KxBbVuDkk93QfauNIOB2AQlWW4rDVnTsLHGCt3vom7jh+qJAV997ud/Xnb8eYA137Vflog1+fePH
Di6Zj8Iwa+X8dXRaVrICI/31UDfm9WRqE6KeFYF0kUTds07hTykLyZz0sN8OByTw24G8aYTuSemL
SBxpnapt3cawB3oeo//6RESkYTXgO36aeoaPzHy/BHWMXj3mIHAkjJNjV+zHfvUHrJYTveNbV4YV
2pGZrf8swyzawGMI6u4H1414td4MiKYyjXlgx+Mkdhkuxdptbztli0QRzxkFYp3O3sdrRvIWxx3t
doPYcXVjcZpJaw0P4EhL4ILI1PIw+P0m+VTYEQWEm9lz9Arl5/szldKTc0dpNYaz9wmbFSF1sqYn
d6FfZGI3bLt2azHqiMm+PDJyQEfSkJfhMCPCu0skdt/XWq4fC6vMFqkaaNQ0HGzIQ2HbnGhT9KXv
097zdWo7gSjpiA2rCVxkEyTIj25EoVHJRGTrAg4Np48TQEa0kH//sO5bIHCo+VEKxvSLzchlUZAh
qT+C7NLVdCit98vdRuGNz9DErm7v2SQttgz22NmiQ0pSbqdi+8mAS2k2CYkepImMcSDDfMnlTm2z
Y7WkP9rdgOwjKPcGEiMRjLGh8Vj1piW6xGQiHXbRB4eorMNaL7tMwinLlHRAHpV8/zGjPMgoZJBn
wXAjoUT0LIXffhnWRiEDA5dOVy/2XB02nuVWBMOcWeYIOpNV8tRBxy9tCcTFDNBaKrFNgogIENAy
YXdz5bfriBYtaTdfGcETAhoeX3xrP8BG7eAbNfmi3qiylOtdfk6if51cuGxJKxL7lYo9a5vt7X2w
CTPXCq3nK/no23uxzT70cGEDUeq7MfJONi6YE2dIX/CwIhfjD8ezE1k8+Z1H515SalUIHyGtjNXi
aRa2s0rCEi19otEoVG6Fm/PUeQTFV9sJOasIQiRBxeqPUQGo8w2ZbIheZa3nHvKHieAYXZL36I9s
C6e1fxW5UUr/blfbpcLxGzfEiFEHIs3gB8jH9dkQB0DvCNwa36f4ARfy20J32jzmwHOk+EZtJ1eq
8rJnfVDVeaNkn9kST0zcBYlU9qvaVNbhwl5izAyUBfyQJd3KOcjBWvZR7Umu7MI0bN0hEHboc8bX
epibUkhfLxGsHcU7AHsN4lZ1ifpxvoThcQFCMQeXK30HpukRY5IT8idYqBjoHFN7iEtyMYJ2JwkI
xIOwWYaxQ25iHWCbH1zHLNoOheST6IUQwVbRWS9M1cF+i9DkghFhjNljKMVa7M0RP2TfxALw3GgC
J+ItzgUNoOjMrwtuCZY/uKjA34gD1OkAwdXLFUjp9pszn2w9C28BJrT5TvBH7+FGqppEpvf28ECu
4H/Kfnr2yzpzo7xTIRKokF2+PIo6TkNufrdV5CFJdx7A6yXW/viJn9Uc4qmipg+RaUQLc1983Tmb
/TiN7rwBIWvtilHZ6tLj9j8trfES2fjbc3fl1r5EGsWn72whMkLBZvQYcQxNyJtT8C6eGK3nOv7o
aR1MM9f3uiaaC6gASa9k8yscLbwHw5b2ip5X2VzJhHqWNmFjdNamONQttn/pkWHODA4G/Ff0mBuV
pst9dcqKxGBNaSI0rL9UJ2Gppozyfqnrn9YLHMw6odVQ7YTtkm9qoPBeuCkyz85p5/WPKKV8ie1/
rsHpZP1MdS1QgCUNXwK3vLg72M+LcaxDt3OW6bKsx1FHpncpdv8hraPdgPVjRGyzvQC7FBkC3kKK
fWrFS8IsZrCyyu/slC77WfG+MgdJRvfmHNMfnjqEFlrcvkBMSqFPenzDd0xz4F2nDjDwRs9bE85u
b3sihKgk1tUhfO5ZZQneCZdkS1WbWcpRxbY7giKolQ3rwYwDofnz/wO5vVCdAZegS1fojeTaiyF1
vOHo5cIqUXyo5ugjds0SrAOaU7VwHU1CCEApvyB5/evDl7v2XNboOVyh/rCEiojn+eoe0Bgkxqh5
9B8SVXn3Ty/yWjnGkYPWAKNUlzfpbWRqTf5Sw6cf/zbUYBeYAi8MLWAnDuhJm+NM/gjx/iuxMfMr
DP+qkGZ6YQujd+X3Q3/jlXNq6ZAGU30re/EYIOqD/1I9dlalFr2mDkF2oNKlz0QpVki28YhyLyLZ
u5Wfap9eJhg08t3SsQ0vv0JSUuALjdAk1MI5OwC8IsHKVSvPBL3zOlgg+9rkHIuXUMg16Wtv9CrF
WT140MG9soQyxJSs4DXrJ/4Mlhi9B0DdRK3h1DUFyEoMks7gZEkKEKcC0DJqvTx3BaI8mJ8GpBV4
4kh1tua+4cf/CuEhJ4lhgaDC4xTzTqxFhz1oyc/MfYOar2oxMWALNQSOgFmqDXQwUOkaYWTEY83a
Kh6TMKjwkYpv6HMgi4KdnV7albLfBdYruahCYSlAS2sj8P8L97uVlp7B8LF7JpBJaglZe1enW9VW
g8D0S0YXYUDNgcCA8BWb4DvFveoxqgZsAoabcH/1gLLsFXs5xYCaNAmp6oPAca2yhDu2ECR74esA
fo+6m+XEAnLtp8vnp5ZAufkEXsaFtTbrG3W4tZA9ZxMfR1Mp6DmI2RkFM6My+4ZKGhvZGyG7PGBE
UPuqOCXkncNmG23ZM/R/Be622P4I1SogSWezZcNOjvcZepEU5X7oybya7XGLg0oA9z3EiLcjb3ON
+atS7bEHMOURg3AfLaglBxx3ip8d30VhNX4VTrWbeI6+MyuCiy47QLsr+gFjTkR20Kr3bXx50XRO
j+IfQBdH2zgCiL5l7nF9Wm1vhJHAsKZGmcenXYNlXfb7sruj7dZ6lAGdUwj+zgryefN1Xg7eprGs
kAIFPXqJ48ST8A0nsB5U2Ehx4isIQzwYpt9wyvtYkPQiAs2mGq4ik1vYT1n/3CHs23WS3SeZYUtH
3erJ2CVM92jgzcq+1geqDK1cA8gxQ9jxnuMHjmVzYlEUod1oqbEB/ziMOQR7S01Rur1vU3g77K7j
6QmoKf3w+feCfGXT7TmkmqIVxCTwEAdYx4TprbLrMSeR5SmmWwQPt0kY4kLADQMS6RkizCDDsTfl
gA7wXdlyuHTKA2AZG948Q+Wh+S/GC1ZUYVh8ADQDJGJHpo0daf5tPVCq4Pc0d3bIOb7v6haBkmma
P7oC3QbymlsRXjFn6DOwyVZu6bXRG4YMyNfBkud87SYxj5uztUks9IU+VgcPFy2ZgBZHSGrXoC0/
8NMTm42rCw/Ch+qIeUJss8nhbrW53figQzQUh+6MwxOwoZ2PxFYgeffuFCz1j5Xpd4i9YljLay29
w5YnS232Y5lCVuLrpGTBo/EBzj6WMaY/mLKiVYT/QeUh7+dJSErD4zMssHNZrN6AcWgMo/anlJS+
hxkaaLrQkbgKIODRf6OygIjlOgf5HcSqkKtc/2zVTl9EJ1Bf3HdAOf/WloFG9mP0jgaGtpTrxEiV
3RWnU6vWfPniWgUgMJXMoUnexr1/ML5TmFL/UmihHrKHXld3jcKY6fJN5xSZ0N1BozXvGxwVmM/r
+f3s8Xl9/m5NaXnQ5mzRp7GrFjRnlnZbLC1EUefTbPIVi47y25HaL5V6mNyn5uGc/OoIKVO4nByZ
Fz2donEIvbamHCe7WwcMWcCP2OWuNrE5maD7XKf684y7tJwzj0fFrcVGiBYBK374a5ulliH4apb7
YvP0XiTO044BfkUqB5wAQ2ZHtZkrWdWs3Ytw8wGNhe0MHVDSGY594S8mREDyC8KwNmk2fyaoNsIX
1/OWgSP6gUQtjrxnokMm+zAQU/ao0ORsV0vWddCO51n4m9DTnz47TH9e0sCClR13nUdXYi9su4Uz
5uVEZZSNDJf2/Kpw/4FPEN2AcVpwIL0QqZK28kQaGxZ3kf4udUrCHaL6LFyNPMpj6CqCQ48TXY04
x5Q910heXdHFByzUQKCexUNB/HoHo3xYQxQKjfV32ta2R1b4GUYmUqvxOhZO0i9norenKFHbZMCG
h1tqmf+ny1EAubk/P8X6oYp2WO6kgOnVMZp7V3b326RXvH3tTYYeTF5ynCwv48SRmi24sqFYdmEW
3lOmSgoTQzAyRmWhRoQbApvkPmOAxVkMzKWwRVpf4f0A6Hf3uXOLmM+qyAipOA9b1IZmnlqcPuOo
VEdrdsxZVOTC3sAkP6GduLNrrtMuTlWjmNsaxx2u4lYTUvprAE+n9CTecVP0jMUvv7D4HRB6YeC0
7qn5EyM0Hci+WC12IwTC/zXsTnUtBKwXTCjc/uZEOopaQ1EU512UDnEekK/tvddopxIcIMAlHLlO
4PN4zB24cF6f8Xfn3z+Z3ZFGSzVQ8j7qhMc4UDyjtzEv4aXrUrPXdGkFlzENlSvooWNyW7Uw/es2
2wwHvtgOaLBr5SpppxVidwm/eOMwSbDQlsN95qPxhVpZoxNPOv+vnmQYi+tHJm0Jy7CGmUlNJSqm
Ypuee0jnSJ1vG1bc3ktsnqQHN1qp4ys2eCzwLCbzZ0XLFcYHu2Wn25+JZMNLk1pthwBjzoOmX5pk
sOfol7Jtc5gUEokqOHV+z+4h/7elOEGcqKHDCD3j/O+NuKPOZI29c8XtP6XAa/Z9q17n/QyllTQR
iQ9Z5wCR4fxOpISaCRkYovQluZdKm+8SBfZdTfvePBztz8uzpECa9x9LAP4k8w3w7h0ZiQdW8PFS
zW/xRLInKbejg2f3vbeydAiTGlTYbCDFmfx8LbxCx0EJG8eJCWPd9xfZS1HQlgr7vqpwoyXxF4S1
LZ53NkUn8nxK8BJ/f9oCbr3rrJHOAFKiLbNi3Ka0d4nLOXeQHxoFX7Hi1TkDd8+WZTvseeg6+l0O
plcGiokFMh0uR2zmBvntIDKmwkO7uCKh2YjQa9pQzvTqNF4dEIEx2bpsL/9PrjpzLu/sDEL3T5Or
VU7HLuk9NM/L/qlfjdSam5kAl2hSm1gZ1UGaRknBQ4Km6lcn9xweMMxP5zbcWAdbGOBvz6TbTgkB
7Yxr3ve0iAXDIkTDjzqzzPzfrumgln64Y745S9lNIo46tL3X6u8VXc1B3ED/ykHcXUn7a4cwGRSs
2UhxsETtC3SQFLQV2rbkILyWAjHTLxM2don9w69P8cLFY6uHwB/k+KhrYH+1jpOBSjVQaNAjd0jG
M4lrYEtDLvBZP3zhQ8eG6HaG2JtdveG6x644vuLCYph7x0SNbFIFsAkYYg8y0RzC/SnyAQKQ4B4j
M/bxv+raV/ZPyz/qWauNz8xN0WK4szeZgBMzx2iozxTbrDq0aV24Zzsi/OVB41EH2JEk1vKUzC/8
yQVNfD2ezj094WbRfIUtFt2sBX5S3UzfOpKMi0HSW5d+tmnpUo5TM6MpXsg397ERao+3FrstBn08
Z2NkBTzZot+9NQCuf+T+feYHVkJO/l5XmUJYq5lmlWe8Vcq7hd7x6umdZtyHel0RNvXeFYYSZ7kz
x/3n7eXnWQ3/ePSstwq0BrbvXafutCeWLDzv00WFeouxFB/pU9Z+UfjlkF1yFi0vb+6o00qrPmW2
mUS9F2smiArgolQxXgNjmTf7b2XFMRvR+VNJx9XYgqN+Gz/XC5ziOMQnVMoSfX0U7hWygn1oZMtH
86ywC7EBqdqpPMkXH1xrUEwYaBZz6DfUH8+Esw0OcurVll0cbanb15WlHzQICxD0pNZVQ4fTTZoE
jILeeDQFIyYdoRCGUlzUYFsFO4pdkkgiBAbZ78YJ89GS/yeyB+VpXb/9SMoDOyjc32PU6S24+Kws
Bp/O6EHWdUS+LVHMMBOKy6zfCG5rOQU4Eso8qJC/RTxQzylFYrX9nVUIOLRA0SySfzpLwjOHp21p
aVY/JnjKUB/k5Pm2j5YQk+eMwVGzNCyVezB850OQ1Yg+v9emMs0Kok5/obB8pmBAeDIBVGZ/1mr0
s/ITMNP+mj/1eRN+dwS6CZgYB4FQtaQFVU+R6OMjBisO5ztGqxoJyquJLCpAetUIcmdnPt9bvhxV
cj9mJQF+i+mKl5oLNbhcgTbqF0r+3hEDkSRbMjo4j5WSOWotKOg5IRXOJZXi7iMGVt0BYlBBbUlk
GGzWYhAdWecawAYWkOKHu3HUFn/GnR/zcFlFrq4V0W5KvWSoWxcHYjmVeTrK0RUatd/qz46ue8Mc
OrQzmUt4ddkL11I4f37DX429WhdNoCebG46vFEgrdoaGJIZ7Jx3uqbwRTPWmlRSgcz67h1FZbSK6
L/sgdoSe0V4PLAgIOJXRNsc8OXFWF3LPbbShmewFkMeOBqGXqhWQO5GPNh9ROh2HrIJrrlFg8hUs
ThqsINEU8qO9zKc+jsjPLXZY5xJ0Upkb4VdeWQ3umcQwWInlaeHxXdQpjK+wNAuAF4DYXCb0uBjm
qnTFP/2HSqk77E5YE++wj2vvqviRV5YCJ6zG8Xvnko+T6ne16siCTiRg9BgIy2Q5P2U9aBfmKQQG
q7ggWxHeXylBqW9iHwNrD6H/x6RHkBJEiApW6lATOQBrQsBhCDRVqsDjdFTEp59w+jAorOjbJ3/V
xXAnb+VKcSqMZauCB6Sw9eucp88+pNFsGmDSzy2dVm26aW45gVYgB1slXwqM8agjGuLW/EpFyqzq
+4946qx5+SvndH9PG2jCppxu8FyiXqfRhWphyhWU+I3/PtyKbUjDzFzXuZBVVWeb8tpcFWc1dU0+
b7Pe7UOz8s8uc5vTiKwf2e7qhVQscICA6Wh74dePNnXAjxFNnqmpC9HchGAswGWu/3kilqGzH3l7
OUKdjQ46BE0LXy8y7kdfV2J/BhNbDTKhO40YkF1+xg+mHF6iE124pcb8OrvA2w0Br0/265Oz9Lzv
PwpIkTCiyODp75qmeby3tSlS8ZALozdYuyC6PDBOJR5/rKACs9RmjKTVpX6XCf7ast8RFw/V7B5U
XennuV4GVLkjZYhoYdpzZzOI3AJvXNkyCaCcpXB6CbvZbhZv5zQ7B8FIMGvKKqJjjbvBUFwFEphM
8uWhBmk7Xg5XlrX9h/JOtjDa+4VjvZxiDnO0B1jFxT3ay6a22Lz8aww/M2d26Nl0dV9jNnS3DmUB
F7RXC5BFGGHY59PuR87AxdWOAo8GfnUb+cmHhPKiuScb96cxcCo26Mxgc3oTBa4HlLr48qiyEpTp
O+0XBIAoaK5ThwQVD3qa449OyD2uAFx1jMlpa3vwitjUmaGRinTZAmnGFIK677nmeUxJKgGx+Q4W
Rc4001A5LoXdPvHuNHT1VlNKFwJNybzB5VHy8yIztvImRaIOXu7/6sxxhAshNBCRjGeoaWhPf6K0
uC0wsYH3F8GoQrthlYMbc+vtG7jSKCcelMF+XBsPPyopmVl/Sf6gT9ZEuAeAertMc5Bga3waXIlt
4yerozcA6+iwLwqBmKJZZQwCK8ZVIxqnrkU7+RaXvVB3VgMNyNJtxNF6xRFZsSy+dKWh+nhkwaCz
KunKvzToqQz39KteSUKnvjJ7f3zecwTuWhrEXwhYNU5lyS6RvohuL2dt7oGLnprOEft49uNmKRsP
XgYtATN7c3vnZr8Sbs+q5j/wBCL/nREmQPj0exVTlk5btQPfKW4Fb+5m7lscFdx4aivhDFO1nf2H
Kr8BTCbLgjpgQUZV5Hx7bzYULCThrm+BNeTehMAvLNzqh9VIHRrfZNx09kqW6aWUMbpqsIObxYix
O+JokOTgYCvVSsGTfIDFxpN2lJifvVMkVViyDjMh09lLp6jePToH0KjgKNe1YI8HCJwqC5iSTaBO
EuvjU3jweFk6WZNflQLpo2GWYr3+4bAR8k9ZhUfQ/jcnrNPVkVBzUwYqcc6lYaT1QpURA45ZSmra
gKtU4o0=
`pragma protect end_protected
