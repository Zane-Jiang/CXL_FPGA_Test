// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
5W3m5aqza5XmjgiEUM2skRy9HrjRUL4mc6RjSYLiDAmtRUmI8jnn92pLS+XbD3AO
lAfqQrTScUxZ/qmP0cvLvoXo8hx17wePnjUwKbl05mwBkGQm8eqkzLEajNGI31Vx
0F14AOXwJ21ps5ESaG+hc3S/Va3B+Bl/h6in6EQkl6l9Jh6qSt+JHQ==
//pragma protect end_key_block
//pragma protect digest_block
2FXxPDY2gpkGOVKEMCaGsp7rcNs=
//pragma protect end_digest_block
//pragma protect data_block
TK880oyorIN0I8uWYXLsNKp4FlpYgxH4Z4YvIAaoHZAWqi6/99xyepWK+fRTU334
WDBA+tbAanoaE0um4/4MihM/4xHBgbVCdsQ6iGtP8HmVKkbC6K9pE3Hx2khX1VZt
Dai6N1bm6DUuTrva1owOeeGc5tMKsvTg1uf507/9a8UT4uNOwtnBgdblGmT2dSeI
635eyQeL/1EWmt+EzAQLMnyQ8JtJ4q9SmCm2EgXfSuk/D9mROZ3vNhN2BFCK9GWg
vD0gozUji1r0B+UUl9VnuKBSyHdQVTUnOd7hHkuYup/8oZrXhfnOmMMiED0+Yj2Z
cteF/WjdPKLLjP/EPsSAbfLMWyXTgBm811tpPuZJA8BuHWz11Yzxh3KDIE7W/65A
fOMw5Rveby1K+74wGpqvNmwA0mBbyP6nUeuoCTWbjP/srwKJeAbhrvkOzSvdIaaS
3gNyIMeSw73mSHRZPbXZIVj/irC+9VE6xcAUzjhI6Zy9Fv+dL1vd014dJbKRavSL
lOUzrjnzMYWZmG7h5SHBM4uiHYLXrTPNYiGdgUT2aMtdY3Xje9jhHYWOBWytVjYo
ShSFSHXpglVrvcKPJJQuDDcxTFzfrB3Be5eAVODpUatn0HnH6giOtrhrVBKARDfk
plT2n9VcJBy2Srlu0Hh3JT0fL95lzfjsrQPAiw4usXq1esxye3fTsvEYqdIsFRtj
3/31vdjqO4Ywc2tWmU7I/L6gvOmtPVklhXPYnYOF/LST2eS5jdvFejD4QidXRsXb
SGG57RY3h3v90b9MwinCz157k7gbvCb4/n4skRFg79CHrLExV1A+Ddp06EzZSDSH
ockUpcUPavF73ond9gwLy1WjrbFdT1RlXjU4wg9jed9yu/06Po3+ShRzm9dWJdj7
8R0v1WQvwcd+HZlqzl8zTamzO8857S4lZ5Lk04ZNaknfROlSdZCDoewLt2BzpfqW
1iGpkhxgd5mBlKrJkV+QbfznWAV/QIREGTOemjFJcEV4vfDxIWp1F41hviUyMRaD
XVeiqK9glXZn5ykhLJZ0O9GiSjZnDePms9yfmbAr0Owca/qOSOg+nGehL8MF9sU8
nkjsG52IZUL201+Fh5eHi1pRn5c9p7lTeZWU79GhpKve4BOy3Xl0oKGjRFrrggd+
/8oTBmdpzJ1G/H2NukS2dfsGJ43MU/rhp6iNaOzT/CnMialGGN25LePWEhB4HF1u
k6ncXkiDZaGRIjjzFdYSLAfWpnzWO3MxQ83kSXcwK5ioZlXggiI/91HN+isyfBlW
QKV9SCQvcgR1g9sSRpV3r/X/qDP3/mp/lPfa66jKFXBltohI2KIs8PWGH36BxA3W
L/rvKM5p3U5d87kxd9gn89sYRN6Kwxfv57qr0YghsAfxGHwdC8UVH0EANloKrpJB
xKM/RR8yw5gl8yPaL5/qyhQuQEFm49h3am/ml25K8Q1rsJq2aU5WFjUCdOBTzr/4
8eNo6NdaV6QILsO0BMIw3dTgrwyJK92r63x6HrFGD/Xg0VLQsCSixZ0f7A95Btsv
1lnPLJxg0TcCXN9LhZjSO4uh3GbtN6zNvw4I3xgskh8tBWPQbEuevRc4fTL3SKks
YXcsexC1KaXyHEwRjpXYIDbSQpU9BpN/VtrD5a5mS4fceeDx0ZflNQiR9HAJsspr
guFexPzRP4wy2k7KaM92tXq3kX3JyCHsDEAypeqVHQgZ3uguhR7GFZYN2toqhVY6
izZ961YAN4FdZHsA52+y55VyvwbFN1htdJGqaQa2km8TfIPgI0V2gFt77Ouj9KTL
djUnXLjtseNqlFUqimSbjhcF6uNoIDfj/GcL8enNbGs7BHYWYe0J/hB/jM5W99rQ
fE66D3wOsXKu6l4kvo2FqE/ZqCSvGtyuMOkR9z7+A43xImJxtjxrvI9KQyLgtJnp
DdrrLAgDAhoaYjcwIltqr4SpZgy840v8NLEXNis6Dp/7LuzF0Hbqdm2t7CYQlq4B
MD0Lw0d8ecuTLvDlhkS/T1z4OYDiTEiocZb9sDgN9Ob+5kHFyJVUbW3gWRknBLoV
SHZge768Pvxp8MINPHbIZ6MBjwXLNg5XyG7gvRw5RyJgfSLvCmswCwvKK6BTVg1F
yMhKPrwMJOkn67hZ+fXCySHhVNnTtIpKFnaRwOLh7zSrFfWvbTumYK17dIsL5ZNV
fW7qJpf/OR7cthfd2OD3ghB2fi8NdfS7g2SUPYNlBBzBJEAw6laFniZw0KQ9Pzgs
dcklt9xk5mx+8vjPqPcAtcw1SikHSWH/uRd8vBK/91/XlixsWGTqfTnW5nJNTVwC
SabH181xbtaxTCoLd+YgXwOn0q+VBXsSmkdKysSFt/p3m+A8+rf3wwNtAeDHNcYL
ACWinucspqbrrErSEcaZi07SS+X0z0jDcPVoM72XyBkAvmc/Odkasg/zbQyl3msJ
LzG2ggiv+SpV0fEPNZl3AimoLBGkD0QgE9aUZIz8X7vmkDG6K+mjPIc8BgSCphpI
MdaTN80+D0PepLcva2kkLIokJIC5bRZTeUrT08wNYxrRO0XcBUoFzy4Te0ThJ3nJ
O5bMTS7lTZ87KkTyHdzJciJxVwqs5kOJKik/U+4pdK1W07Az/fHHHyXOLPWCl9Bl
bWTTd+ZIHIQSsWjykAVANz6vJ7lhjSkj1l2D10Qa90ANXxtCLj3htWGuGDg3aGNj
ZurntP+Nglu/VqaXaoHbdBgTs4+Xk6uKuhYtf9qMel5EGu4Q8zt/RWQL7azO3HSF
C6e4F+G2u8dIiq0s+MlvDaHDO76lu2oZEFj9W8ALoog4qQp2ARGpgF0jo52PEsdd
xRvNt0T7nHWVuYvt3nBeNABXW5Jcskpv6KH96gb/21Gr0vxTh8QJ2QU8GK3/pUC7
QArA+R/VrjfE9KYiCxdRktxitP6DLtUSMh91bgCzTVp9I8+C2f4POrfmc74FLNfP
E/3tn9sUa6bLW/35fyrW7aoP0fjVqeNhzjma+m653ER6dYLAsup4sjXBgNu/KQRw
HwucrfHihkWWUzL3ZygKnwxHtkLIeYLEQ0FWVU0th1MLHLOrl1BeWQFBpTkrDg/n
2ra+s5cQwrjvT3bnYfpdMzyNxD6g55IOJpcczjEOXQULVLGGR+uOdrZuP/4JYdhL
wYnB6N96F+iXM8SxdHM8hByV0sy7XPKxbZ64sJ135bF5gQ+VlBETLsYs1+MajizK
pEEeIAHtK+OkkrryYyR3GACy2+1HrJIHeBH5ZIfLSItJ6kotRgNNZN3IwAuM2/ov
yB/2B3hK6E8DFl8XBwzWCZZ+f2vAfo2+1Z7x9shPPmYvGEzSuVELkn7HbxbgPD9U
m9a22R7a524D2hrr6LoTRZE1Vkml8OURc46JXyBnKiNPSMFHKKiZFPt2wXpys1ma
tt2bvnfxs9qTXL1esSdzADDEXAjdXZdBkCZ1W8PEa6fLbyPbo3OUIcSs//YLysZO
rCr80IxxVcs/9xP/xpPgGRCW/5aTrKWvRj4AyJOQqd7gjcg9LXIkM7lCXhqPmDcJ
sf8bH44a4tYNpgijbNcHYOZLS6nuYD3BkG0oHmLOB33Hf3EaNeNfDCl0I2FKTH2j
349Rw7BT2C/ICQ9YfOIh3G5jcgXwsat8Kbp4tNXoNHLj1Qlb1G3gcwV7JhkrGbCu
leav3xGWXw+F6RyJtIduytHe1xForh+fWd/ayLrQD1VhFnYHKcqMxNea7GRy2+XE
0O5QYqTCjlqmzR7HdpjuyVYznkjCrIvWN8N81f0yy/cZfqeq4vTiCkQyKKSBt/ZW
MQTLXtRC9Z0hes7REULAbtRPyWVvXJ1c/+P3zLBL3RaYz5L+8Rk29Px1L6Aj1OrF
pwCX937JbYu4Akeo9KyKLCxzL22vg/vRIQgWWFKgW6seOWyweegEOJi9yqQX5H04
z7FDJqwh/rdL4090cE4wrEpRSkmM9keSSsfHbtACOX2K1SgMQs6P6hjmZuXzrW96
JDzM54sMueqc6u2uasxWra5qIZ7LwoS6YeDWUHSphzit4gqfltLUfcQUTO97/B1p
Igl5bBbmDQaWm1frRCabKVdR18ztwEbQk6DZsYkem4m5dGV89xM51j0F1BSo5KSH
jUnJDlPAT9T54nlTU0gprH86m3znBOeQiNGrcGLD2DCoF5Fg/3uoTzRDW2CSDgqp
xP7/YTc7OLpzzgY7vtPBQIK/HdRRc5mRW0sQg83XfTy3Fpxti2CRLi9icGNPVMx2
/9vSCAyrWVHFOM/Nh530FYQ6T3GvJKaxvkaXoao6aW6+qDXld65lWYasnBv+diwX
Sly7QiNzgzSTQNCDl2PACgxM9BNDQGUaVpZubhsP7k4HRMSgYIcNkTskcrHgc0hV
gmTV+XjayL/HoHcWK/Xca/jVKsEevl/+E7Z508ssc0xPh9aAWsnvljr9uebAw4xf
hZUflP4NEQo1T1deqlSpkjbj1JxLlPr35UHPcv5FTDuMz2YynOy6e4MCI7Y6r7Tb
L5fy3O5Ux6HMnnMJCW/hV0Ox/4erq+Z3c4crgBiN1GuCIeFNrEl955VIOtYltVfF
aMpQ9AupWrOGvL0jHwG/Ie8kPuyDNAVnqTN6XuJBfW4z+Rgdv+8RdzVfvJf0I+ML
f7ukuKPFjxcR0JgDLUMMSD67/iChJMVjRzuzW6RLaUfeLZ5eNqH7AWyZk9I/pwGa
j3lYsxWQsQN3NkjwbthDBUT8XEZ6GMOmRBSgHe/ccm9kLIvcg803vkccQRbieq8i
rWnO0ytqN9Dai0sqJ+1w6vnNmQ9g3cD4YZ8v+xto62AW6CQRsxJ5o5lehKzzvKWR
6ErEr603dnPCLaZGpRH8++kGfwI7X/V7TgxEzAHSjDMGq6j6knGzvPqm9HuGrLxy
ZK3R7b437cnck/9Br+Vju4xroaUUqh0tJnBViMQ7Bm4Bx5pVBbu8WTXYQpe0UkWV
P8elvtxktG6dHu5mpoj9dBIOZZIT1oKZAT383nIJ0jiruKntQVcT/Mi2veuH9slh
WzNecZCD9H5sIrOPyfLx66P/VYQJECs2H7jvbAqEs8406EiiPrjhH7D2VybDTung
Zyvdgqk+0CmYjq8IPYYlzKyomjwmI6GMsmEEPx7X2vgY4Zg5tltr5V8WvVVBx+sU
OEl84eft2qdyfhT6mVQQi89HllWqAVxP3bjKegKLZbZK42/PwotKMGWq4XLN9R5y
UDA+PBNcPg4eMAJp1hTAuzaDmC4IgAm1TAofho7MJ/kigOg4DhgmyoYBmUMoy8PG
Ou+8JrAkGoUmp4j5LYJGdLEY1paLIaRZVgyj61kuTEuq9WtkXtTvFTTPqOMyu6ly
jIF+E68aym81Ib9059HaxnYups2he3sty7mEzgeralB6Q17WsTLb4bM4c/+CZ1Yu
LnFI5+SyZ4+Rzj00gM5Bcl24wOanhZXL3dSTz56YvF9SVyl5RCLXx3OvICBHnpPD
Mo/TAr2faQLpBcmoeEuL5GFfvRw8R+VGeabhwRXiiAS5WVIpZ1GEYUkoRFq2AXQN
QulKR+vENd8sjxU4OgJVr/nVfHuj5EJyskBD/ck5NvWUqp1dDsar11eD0/vAWA7g
fVl1AmPx0RO4ox93FOi9S40Jsf0HWrJFWTJ5jvKI73sBTPsOVwIOinHEx05/612h
GmGQoEQxSXpJ3z2UU4aEf4Lf3jhdOu/W7VHZMlubhiHUOYZh8my1O0uq+AcnjXla
9MURaM0Knw2nb4yU1/medcq4J39m76vUL7pbhDWAIqK5FAy2qFfsapnmDlY8ZCIA
9FgJaDMFrAtjaxyFK2pafMIBLR9OHFDWyGN0ksLAwJq5tsh7RDNG54Of4gEuWU8m
qXANdbTiWTxt42ysdZi0g9JFEZNUlgibf+q0qNLzE+SSG72rIDO0scpb1SUf3Ri6
ZLdAmz9cDTodTPsQ5kEvONCUAFl1nOTSUrlTd8HYCkR7HcRS/LvYepBMjnYNeviw
8z5tuoK2MbbpXxRGPTEwOy4UNWKI+nEE1X0P1Xzmj3tnSGolyrAPqKajx7brVWk4
ANeHG1Mk64Feur7+f9Gt060FLiLtzYco8HScQXPhxmVNA6mzd6fRuzA/PnTlZOMe
tK4fDCAUXFhcpR3+IRUc7VLQ+cNHRarJScSGgAi8nw2a/KNme7gKNDH1hLck1C0r
yiyQnTi59Z55SxGCfW9HRY0JjLz/EeNMFckdMCMufm8c1Gt9kc1N7RI+8rPXi6bU
GwKxuPEr6cnZ1XjkjO0TWyvaQDbyLd69mqO+nXc4JG0MojjfOE8xxDYYfuDdvsuz
TSW5Sj3vVWNDb5mdhRA3Dv8GKytVD38BEx1bJPvIc6V8DTns4lN2joJJ0G8Tux1f
FfRVzKADtpJF0MLN5Rn8ZcGNXY9xPTw4VgPzqT4oDiSS974mGgOFZjAzaH1xOAPN
85di234OgSpqKRXqMRSjuZj+U4vQTKsjBl0nbrYlEKbGGQ/wI7wLk9ajtRbTG7uK
oJSKYAhfIM8/ghwzT6Auu+9n+KTxtqEHctNlKBua2C7Gl4tYArdhdU0+h0Amzhb5
2G+D1Go35Uu0WT4PAGAgasNZjTXRAh7yfJlhz1dmVsZ9t644xZ0+S+ZphjhYvBBh
QVzAoHWetUjmuKpS+l13lxhsUelDG4VNFaYH/IewgVFC90cUNS0PSRb2T5mHgRNJ
Rmcdiu3JFD7ncupGNtTaSHzRC5RbjMutmJygvZ9tcvniEuHK8KK1//A+8949AyR/
fQdI3D5Y2waJAHOPwRZaGI0/oPfks2190Y7QYP2qHWAkGiATvt/w+BEZQRInSlIO
RzppnofwpPtxxviWmOoCdSIOv3mRIkn4SQwyv/JCWixo11P9l5IbCvcNaypwVpsH
xmuVXVSgWV3N2wiD+vpzKyL4u8gaZYHc0+D6rpToEGusCBz8wh0gGxyPymFfVBXc
T2UytUOOEvFZQ+U15+X+gjnyobZKh3fllG+HmFAkoNpBJkJSlDAJHwOKZe1XpxTu
DNZoRuuCwTVM5yul/hgUi6oxrknU2k1Rhd3otO15YzwOHCM36wetiT4lg2P1KmSw
bOvoQt1NdIzBhXc3pDCigPuyHTYyFdMMbXlWd8NEEWwe46J2yEgRdXi+B2ROrLX1
yRnragCwYKZcUAD9cCGgdACj/8HjFfZ4Zs18El7BzVigXagaCwwCJlXqSagYuzFN
rPdbjTvIKYrAaiAJMEaEULKoWgVQKuXI8dw3eAl/XyFMMNLAhFZqyq+lTVAEfIcm
yQYVBGn0Jnbcxm5224ivhHypejP9L1YgAo1T8iVHU9Q2OZ4xlrbyM3D+y0yoaPb8
EJjZbmMbnr9Ur54+JKoYqSuOGFJEf5peUB/74YAY6DOwmHqtu5r7xrqmCc8K6yB+
ZcMYnAWearZdUijBh0jDLIddK++y6IglmLSjG5ZLXJAcAd/sHjmFREa9bVXYxLYN
mA++j43rgE8/2rXVaxAPBHuefB8g7atLTOLHNchZ46VIY/r9p4ail9f+UtOkZYoD
K4u0AiL8Sgx5xl+cz1By5fAp/zFk7rtiTUE95CW0Pk/cvsbvfZBQOLxn0dSeAH51
2sVRejT86varhKaPjs/6dg6z1wpPlX9HdCOpFQ9DkZXrzlGGIzeNzlzjv1It8ruT
HFhNdhoghWsnllAJ/y9WUDbtYvWwSWxAiHB+bGwEABmZ5zTzoFnC9eNzd932zYp5
PbFFuCZiqFlBa4E6uOLep/e2L1AEtQPSonCcY/nqDIz/QEDVuhY/JOIQoTIY4N8n
bmJ9XI1MXZW368LKla8DhFucBHuTbmETn10v98g43peIixow35QoaGghu/o+qtkQ
JYc0RLiHfCG24e8y/BM/duhHaifviQ0X3hGaZ2mVr7WIwjgTOgzQC/2bjVTctKtM
UMttrq29rTVeV0lrez1KULULyyBjCQsjM8QZqFVgVa66YGRJhdngFaYGuQAgt/Ov
EnzrwglARnK8eHQ3rIhJ4rbMs7RkgFNKmDb69x+ylLvtyCuTZWDbnmmOVmH22PFL
xV7/cZPORW6eODRuIkdSJneo7zMYOv/1gKSpOKHDexYlWWAKDMjwBE3vxUqGhPUe
4ODrI66K3BQgDyBiWMo85K2q7I8ZMtEuKSItnaNBiBaySL1wiYnqVS/gG4m6n0gV
bcq5ijYynwPxY2u/xVguWNcdYcyNqURD5fxw7cC/HopIfhVVvbepxU1V7FklNcG0
RBixX/qNY6gebs/pLc56p+sW112mPVjbuihmxeMKbkcTlSZuGvRNYZh5E9NOy8qS
IKKtXPNYv1JqxXFWZGRFZaTHVifN/VwnC5jj6pCtC9TJQAHaXEgUNirtGoDe6Clq
CZ3rRKKMFEHEY+10TnMJcG+DibD1tJyr9p5Rlr0KQAjKinp5PP5w/FUGVmhoVuDZ
zdeILtipaioG7FRWg45tTKq+2luUQ7gEWhY06m6tb8Nrm65ktAmxpnndOMjv/nhH
0HMpxlH4hlphXtzEy6Wdv4BoP1D/8zbAvBGyqkiXWJsqzsR55Zsh4J2p1qe1lSk9
f7sufc9p/NP5xLqzICOv6A8+qmN9z4dgJs30Z6MWQFNDl+/l4k2tGwrJs7QS5URw
dPI8uKmhewkYeYhOEfMe01zbwhfs33DeVPR3sB7xNZS8vT7HHtzCA9+zwI80rFM7
JN5F6io5RBW1ByTdOK2FFmqf35K1uPgqYfPeR/ggT6+BHBo7nE4D1wYjZ34sdQvf
HzoY5fICjzsxEfpGj/SvJt6tmb+Pv9ieBnFb/pLxVKhR0Ns9SB7ON9jSBqK2d1bb
W5PFYBbAiJmPFSl2EcsRwhOHYaN/bY4VmH7Cpc9fgDpB48A+CIPjAKAud5y3BfXb
BY4zT+Z8BBwtnyNtIRQZGcvmirF4r5RL3d44hreqg67fpFFCqE0ArO7Lijevdvya
/1CCDQIoHhZPW4h+vJ1ar3nZHuy0jx3LRCzY4/Br5yoCcqKYKv1kRaf6ISmEB2dp
EaNTe7Z1pX4kiW9apcTimZbaynYiX3/6d1Mb0ItcabqNYORjy+kUf0CALalQwyZn
TNTYNnPmmLUoLOPiONbhIeGEgW5df9j+DBKylB3fXQS7vm3eT4gvsVXhogiZZf1b
Bv99a3oAMbYa24KJh2F4lvZbnyQUlKYtbBeHOzB5/tO9UDlMv2/L11l+if8AFBGK
epi+kso50YzligK6Z4387GDjO3Iv45bMPNIJ09e03Wkqj44oUlL5yZOKhV+6hN83
QaLIKQ4IbGdgF3N23UifCCYxUNfw31pF3HD8TN71G+0hpKicSDaNIRVtzpdzpogC
/C9e8ODHo4nNIGkrlN3xcvpJ7XnI/kQD6qItLn8x9VADH500+WjmtbIKH30XkLEg
mE6apbztCwlQoNpXIjAmphDur3Ppvb2NdcEmsyCIHWQsOyhASIe4rr3nXheWRBIH
7tIEnMSq2cKTCOA3N/VSxS77bZg9ZfNY3I0nUUZxhxAjNp1K8J0KQ9Aa1TDT75Oi
P4YjK90rFed6yMhbnwDoDR/ufbFOKpAf8g8asiKbeOpv8upLRKkifd6XxJYRTfV0
dANvspkAX2JFRofkYRMv5cH7HoEziG9KYMHpCPQFvc0/Qc51/SdhQwbSTEr7MoQJ
3+89ivizFYlGJRV3pt15iHuAlas+HtOQFull0/LMxnwzvPVZWlFHy6ta0grZq6w+
TXZcto9tSfnmZd+CNxyYWy5Ih2SvU2pCxOoOYl3f1qEgCG9E3lg61JfDLqnEakSJ
TYrigoUWvfuhZZc07ftJBnNFqmD0AROY/uN3mfoxRWyTlOy6MMqMbpGefyVv9CnC
whworjWDpKhf9s06n87O/Xv1HsemhPHmIoL+bkzZGWgH7nynYom+Vyt+TWEazdK2
p0PGzUrutY2o0zL+ZUchiIxeaLpbD9c5nR0LAJjGG9fufzj+bxebpc9iMQyCnxqJ
3Pc5zq6DTjuQK4cJCfiwWEkLRjQ5Wv3Z+kqjzxGVoSu5EnQyTVOKc3C1KJtCEsKt
FdpxqYnO1Ho8Ovm4FyKXeranLAbdo1NcW6m03UE2bSQ+XIXlFBCo2iJY2gE+bmUx
SSTWUEPNy6Ejl+qR/IdStg+5aXFoVaD0F+FTvihXVTQ1zznfaoX57ZfyOMKjCsRn
I+qB5qKE2LUNTvFpKIz2VB5Yh0BBeU4YyUgLWlor6V9U0hbeIDATNxXIfy4CDK7d
Q7f5tdOXDLJ+v4xrzDW3IMxilNCA8v/eVvYxjV28CoBNue7P/4SZu/8X5CfZbjWh
athe61xFXs7OcC/BuRZZW7EJzSf6DEjogG+1K2d5j1GlNpLc5J/t+B+VH7auQO04
RXrSIJzX77qPu3N/93e2P9NmF7PioeHMbG4QPmWrFUUWD25koeTtnE+9XbvaXCIH
cvJD8E1eHybMIRLxXsuPKaLoXg2Wz/3oLTpq/6dsuvk0QiHlMz6EZxoQz3BHkPKy
ATkKRcHR/lfF5jZfFA3fsS+8M4VEoCIl5D/xMFstcGURV612bW9mXpQXUrfhw0X6
fqJe+izEwOgp//FhZSgmfbllGFDPd+gF7rLm7oFjaBTYU/rYL3dI+4K7Bx7+hJfX
0Dq3hUQKKTaSdfUSnoQ1tTspTO2Mz40s9491Tp0jAFuLp59dV1gFhl+RU3U9Bwid
UWWm5DjusqlGsLFFTTZPmxCVFUnnjxNLZrd6OM0b8jUggOpjGkslV256tWg9Dl1z
ecYhwDgx74j4PmfdER6iZjZ/OP8Bt1/EN34dAVWpsxb0BRHFbXwkRQ9AlSp+ssOK
tEgXm8FNWXgdTvYBQcp5ZT6puU7+F0oZJzSoFYfcqHsDQ9L1+88pACAaKibsmc5Y
W4y8TGu7aLzpfR74sHVMKm0ynTCW1gpI0sZ1/WFk9LOH2yj0bwZYVpAdXvhekXNv
yKDA9ljMaLEU0aireMVSaAyNLNCeZwbYBAVnaN/5tIamBHOFjYBZ67k+dFHjd8IK
OjZ0me7eesjlz1mQIizAEYzydRVWWegqUx0/jnBqMjtmpG5kiubyVP/HjGMsofjG
DUq94jSv6ggPplf/jvw9hG4kqK3jLUzByeTf7WaA9+/lpZwJTcEWBsPlU89J1M+J
ALuASIa53Btz3inRSenxW5fjpBZH0zUcE5DnfgGhQz8b1lcSI0DDA6KRCFAn9az0
ToPyaTnicVHwn+9n45dOzqF8gfKcbEq7WN3Cl5Dv56s1gpFEeU4FWTbDYch5bGlv
dUMJ6bKH5k5c0W6/SlYaRCLDfXKNaajUQ20mSIl2T89YfaSdW8OWLjNUOZO3XPqC
dCC0lfF5vPx6qpNVxqCIY5/v0wD11K12eiVl9TmZp3n4J45djl6CqIQnsXvn2BRb
OhqfMhn8mVHy8fVJQXtc66e8bsmjuHH1+k6Vxw0UxYfY+roVOu3pCy9hPMFuJAxH
HHHdoYGUIGz5ZGdZ79cp7+CRAifCSAnhuM+JgEJFvmDuVfZyGt7S5FM6PlT+azKO
h18TaxGzif5Ikiuyptz6xT8TxC7200rz7kcjXoBtBEz/5VxM7Nh7FNOhjHWjVum2
3mtnisJGNzmTfGMG9kxcJryN+SUoeXWZuXz2RZzCZx/6UxjHMSY8Olaui/LdKiVG
f9np98UO8FTKwhUHqXjZBQR/dHz7b4q0btEE9pghuy9EQdBLWrn6jzLEWr9tfaEk
SwSRixub1hDcuqG2xxF+Nyf9BXtjFoB3szrTrOVPlL6b/u+SkiObGBnMh+JDJzQT
2kCUUO5cH6HlX+BCqYGbf+zBygspFM9UZUC/u9K0bhWpu+fHc2HjYNoPAsGubJM4
vK7MJ0RYbX6qELGdh+hJaoYCItLK+DtwXsaBN8sXLBzhBmKWRuZD06XGxh/l+URu
oesYrWUKX9wPyWFB8+j+jHVEg+SSmD6N+oepkBjBs8tB8WZnJhiKkydrCuwZ3I2b
IuzE2HGtYlYJDRwpye0+1h5kO8WI947Vf/136kvCArchm3WyYc+QgTE4OUgYt7sb
SaQe7gvhVjwZ34rbdSVlvYh5c2/2ItZtOv3uvQ0FKm99yZuLLlCo1QTX98Jb12Aa
g65UhO8iR0bF1f91gomFBj32hWw7oUD1uclmwtpYIJueNLHPMuq70TtCEvk8P7mn
gR0kvbIJqudJZyOpaLZedxXQRoNBbt3iihVOzYYm7Fg8ieHmd+LYVABYIH38IYoN
W9OJ+a33RoXJPgXFWuLvr6Yhg2Tsr3yMjjKI3GD9m2tWjkcK5UTXeK7VJmydGmfr
HkNAd3Jn7e0YIjYYgWGxmEsvTldzu8NcRD4A1/t56RUQYr4AY2/NVf66QK2WiiKP
+qE4My9WZggeJqXlPE2gRwprg9H+kzdlWcPzxWP9Gnkfd/qQbCG6uOPRFKm5vabl
ZhC6lLBe2FwxPX90drQIFS6lvU0VrXvTFmmUO8t58hV2PuzJxhEOOgdVu1p+xS8D
2zzVL8xcvEbCVRh9/57TqYZjsq6eOpn3Dfpyavw2wPIkSIQvDY+ZN7KBKEWQTUFn
oc+xemvg9Xhdx+RzLJBL03zeHsqptTh2xHxTEf3wKW/DU3ZimD6KAyxxDbNbvux1
3Lv87M+t500+dtcuUV+REalQnr0E9TfLf8oCtXYVEAX2e9lIYhdPRdr535HfhDVt
io7SolX9vBiwLDUOXV9VVvJyOWt7SDU5Izyb0GIoXTGhTyCrAvxw5peRi1Yp6p90
8EFkTtu5Z1IqvTJnlgB6PHzbbSoyXbDSXyd0mQeRDD9N57RGGePbd4wh6HaQgKvY
xOC2Q+Jhm2eTOC/E3/tX1SAt/nO80xM4yFCTgjDamQ2bVxzJXobJPcvIDMyPwlIh
6P1jIMXoMrul4+uXkkARNAA+GuOxIoRpb+lqlHjEh0tW8bzVtj9yVg941SDvCDhk
Z5fEZwhPdn9R8MTV7eihorgPXrzOJamk3C1wpK+6f1OOp5Hr0d2rLP2yEf7N5ak+
57pjyGiyxuvQkKh/zvANH01WIOO0ykMIaxi2S66OrNYIpUWeM1WoS8CFC4L9Ngj1
1HxHPSN9VMkAwlY160Fqqr8FZbYRodLa9345lENZRnVCxlKcyV1gsOdDo+JtVnRE
yS8SK3MKxIfWZ9DjsWenmD5oGYk7lV9YdZ5gJwX4xmogK9l9QhYvazJqDmfOfZ77
4O1ykRcGJFpBHLwjrv9fDLuvcIxJi9hdB/9KKrqICZ3mf1kh4vCrfzIh64XQtmNi
IFYcViTyYY6a1IbB54vV1xoNLcJynQhqIS/zENmnCuFmsuPwG6jSXY+KWlaf00Gk
deFG/OPFwIpdRtsWYoLfxlnYGdrHQLoUDMAMNhnon7ES6pu0fGzqDXR4BlAQ90uw
X9Rd6MoXToAns6xG7uL6Z7FqP9LjWjSqnZ6vFSfFutwMD1MXR6IAZaIFB5k0XA7c
UQhmwS1YvZ0/nApKwrNmvLM3qP2BhRymA8nCKaulBiE/A4Ry3mCy2nv/EZaWpJBP
g9phr5ckGNCveAB0/jB0/YPB78qbn8oecahh+kKL6CgZ2m9v40mGFpzMZE57D63M
2edVKebZX69KfnqU8y/MV2wgBNaM7rwhLKTEtIdv01o3hkSMI+WZWZ9xxXIhN2wy
/k/QzcO8dZBvY5HJHCKlZdLb+sEY+eWjkSdK2/sWMYuB8U7dgomIE6NThpL4NmJZ
ahR5iYgXqRwrXLkO22j6ELu2bvCB5aQRSO8vPa6RRWAQnhtehqYBUa00eoutBFtl
HUtO+aZw/+sbRM8IuWd4o6AVE4A5aNDVrDUnhgSOgZFOGOtE8g1MaVpBFK7UwjF6
MXynWrlC43QqOQWcXsWREB8VN9N77aKmYJSNV484/7aaQOHtBcBqK0z0INudPWB5
jrflYJQmfVlvFKmEBT5Ew63gT6HY3ERa68vSusSDWSYhlfe3zCaFl6Vl/0h3kGeD
uaU23TdLXuwYkXxV5VGHSCcoyEVcD12MyZXXJJYCP9aTX+Cc+oDokU67yfUtNmDc
LqSNo6IztyAuE91QQfgykMJAfNotCBjRfkH3X2r8rPVmtTQU7abcB2HsNCXTT6AG
QLX3bX46OQCoagArbEBL3SD+4ew+hecbt0K8Bs3CzmfPxy/KFNRkPSzCeugaNWeC
5OKPoil+fkARSssPrGEZ0tE+NsAIuzIYpeAHGoytv8sUEJRcxuOCL7zuae1xH4Su
nF/D3gPa+A5w3kYEARVAdGceSEIAPDYKRA48tYw/UNpCJrBRoTpZQE34Ry6avKlV
THcrM/R0wF+D1bJLMB4jHL3CMS5kR9mxCnAb1YA3eSzriGOWmyfL3bhPZwSoVcJB
HuEq9RTZDF+hj/SQ1AW7spV9eAk4/e6pvkQE7vtqpndk9j/cF4rCSKaMSvFiUWoS
F0BSV4z/H4/buMQvyZ5qOkcrzuLfY8bdn3rOhVO4e99/MhJ/ST/pyYbwes3Mrr6j
uyixtkvGO4QkdrMH4CTKx5FQj7qvg+6fk0J7WTyh5rERlkmADy/HcSDeNnlpSxt7
L6p8LgY8vP34cLOsj2BPuBXuJ2iM416EObwUVVBA51Qcg9vzeX5RxHsCVcSVCLPV
O3f7tBd3/jqVyQpqS7VSDk1oeGKBgT5Zz38+9A+uVjLu/2fw4kQXQvcNK0wo51nz
HtGMOVIsUVtUyD0ilOv2PPM22wx4gr/x34mvCckUYtaHm+FvXGAJNWNl4TOR3gfr
EkHsa2RY/ovsmXBuoaeXwyFZrhm6qpeCRX6bsWV0xaVuebtWDzHK5VC4my8vy7LJ
aRsgRLoqgbmdp173Vg/n4vKMX5fhXVlb2UNXXR1c4z8sHEImRYbyZumVQ+q7/iwT
S379cpFL4nJ/802PoNWD5HDgiYYS/eXvfBm5NIhzKLPJ0EPx1ZkKaXrWjtCf3Dgw
Y/J1H6eC+2PjXHRdO8x8UPm48s3upNc+b3P0CPHX3Dt8FFILwJnqnIYkIDfQ99pk
fG4F9o9WUgfts7O7mg6onh0KEVeHXsgk8WyGgqdyTemKoFTrDjEYk22dI1FjEOVu
lyNhZGXZFXxgGn+FaXgKqYUnSLhZc2nzxpUgG3T9Yj6NA1LE+zX0YlrusqFb0npq
eIvDDrq7t8BWLwTfMg8LlpNv6FXviYhheHuzo24LF+YRJgVlr3+BhjzxaCBeVeED
z23VxfwvcrfNX2cYxA2xFVa0uLWHcSeSPWcDJy0DN5/F1+3W3rLpN2FsXD3meBOh
Hlzv/BAcjkXqDWHDE7nzs5QN9NfevVyMZHT8rUS7zfENRL3P62nkUY23IktiC0HP
4neKoSjtV0AmLp1desq4jwZAdml3IRTBnI2lEZP5DrRARwyHgrj8nJl3GKnZ/ALy
10MykS+kiy84a1wpdEP2PUE5XyXyoJTyitbDNQmkRsDvKrS/XTZj2M+B62r4XunR
uGtwPnp0UJffStpvip6OEK1ePWK12GJhoYHqFluM0svqvluI5PTm7cxD4l7fKXNM
bDvvokxGnNyWKoNcSysfbFSPY+UPhr7/LloOQjjzwXfmS1mv2j0Xi3iH/tNRogTo
4Mk4eQ/47tsBGUXuPzaLPv75WzgJiFBdxEZ8SNy88ZRJQhwlHL0RWNMBvM8QJ0lD
oJkdb/qgvfORKaSvrRdlNSPwjSuYpJdMVyxUIHY/+oJ7rYsbwjrVA7kTRDJZpWjj
RgJ2g+qSLMRscYBFjhHqxRiVJLoODZ6A3XfShj3ReUfZqp6KrNXqHmGp/QwIY3YE
1PKLbbSmQA/udKe9aneyeR2PXCVJfJDNUcJjmL0avwiKZVoCEDe2xqSxy8kWtJWb
KhOzd+h9drY9nXJdzBM2mflcGRnTuyNcExq2fRRxz5oA+dnpcOmUA6LWgo/ARVFh
Jf5d4lPiVwVx6n0a1M6//uOa78h3jjRsLlhFI51pdjWmQMDdSdrTu5u3L/T31qU0
EIxT1e9qa5lUa7/TmGXmHfl6gJ2s0vs65xFHqAH/d4fJieyByZAaHLkQDJZ9myfc
nx7y6ZuH2jnXPQcOtUAZxWgGDdZ61LWcKD0AoillSFfxomc6r/EbOzUlihQEDInx
QLRpYBS882yKQynBXvSHDOzhwGtRBAEHg6OE4iUUSTnaIxz4P+QZalMjwi0OBFhg
wyCOFgxc90lMdzNn3dzB2SQ32PCV5fPGWnzJeRIyqh5UJFKyHnrAIauBN4btWwgc
wLTGO2zw322t22TD9qLq/syLC98FZj/UidL6DpLqn8rsPCn+QRu7HKeF2KefVSmy
YrsxOEN0WeDA3fkIO/izzkNJziRu0BWEf6HkydnOZuDED2EAPtpEgumBhmx8+8nH
g3J9OaFhWuybLdBJLbA3ebYm4LVfZ/9v8MZ5FeRJsWzQMLXG/WUnmjhUf7dq7gLj
Xuokje/R4sJNKqlcNUdfsIHLARASN/eRWZlTVHwc+28ooZ+FvjNOBmOT46aV5bH7
LSwilPNMkgd1Q6xZSJZOLSgWFpaxKKTRZtV77qbgq5nBrs75uz9fopEkQ9Xqr+tY
bXnqbUP/ZSFz1Afl8An3VzbtqYYVIS7Yimep2s8PP8ZsLPqqPSmSoFg6+6COmiBa
bavNZa147p+wyqwW9pWatQ1G3Wt8L+b+PKTs1NuhhqvXE6dOk7bRHRLL5ecXjOOt
gJ0isnS7AJMWozIAMNAyZY6K2lrssrVV+W/m50d4MFzgnwWStlRtVWQsfzbsk/hm
ig7fblTGvjYb/seYtxbRC3LBCyC//RoDgzdiK5+kI6do1qzgmM5Au4+FzZyeCFe5
6t3VpeeXWri792ho1aYGPnrGQu30MtQqhOGGz21gw74VgY2vfB8cNp7PBr9c0pMH
lgRL3jM5vNUgPUSkxPCONp58h3aU0heJ4mVyQIm5/WvDcsG5L+WK/EfJLdS0FN3H
GbZx4r3J3s2M90AGzbSneW7XOnuhVeB0SLZngdAxdc4fEW8EiifRffl7bQBHSIRs
RXVAFV40iYNulIUwfQ4VQkiDkTT2Uw2Us2mNO4HIewR/DB218w2qt+Ap1hi9dI1C
L4n2C9O9qc4UpRyGgE7SD72SkyEdxQrHAUtyY4+dDUFInYKJVtZwb+1YOJl28+s4
Kft2N/ndHwZrN+qKFbffXqMaks5N8kjk95tE/Zrce848mVpb/rFdnts99Lwnf/lc
tfsjSLCYVGzTC/bte4NNr/7pz+8ICB3J5oQEv2MfpPJ/9szDP/jCUnToPdE4GZlb
qa9fUkBwCT5NKOlkgg+xlBYZI8332pY6mTi/w4GLKGkizqUpLBO1jKY7UpyX4HWc
MxY5ZiDD8Efz6y0rRr9QGYdsRu442MLCwKGSs0TXf2LSzamQUHVTa2qWRXxG8PAZ
jEpgp7DKHJj1N1EUifjOYctWGT8KI+kAXBCU9cBsDQjak+kRXmjnbmpbVMUVbD0F
VOtM5otUH+HhvSGl5jKQ18DrxIJMHZ7gJGuBWVgGUFExWSvwVJY9UL4vj59zErtr
G+bER4Mucw5uWG82Zs9Inbzafvrm23kuTpKyQakFkkxkOzcFLV7Df0sm/jHK0/TS
8NFOUo+HCppWYcyV5XDeFUgSCAcHvmC+b8a5ZZGhu41mxqnhdHUo/cMK5RWa3uvU
XhQKn1P0pe3f6IW8IFlUTKNz54oSnW1a6rMVkdUepz0ieOkIvVvj4bC5q/bE7TAY
i4aEQ9gg9VJ1dC/+M9fOby99kSbd79NvapabL5YQYJIyHuR2MhdYkW+jytB1IU1I
qZhK1S7ad1DkcOnx452JiC1K7aPrtwRGBWrzNWlzVK0cizn3z/9wS3ZhpH9HjeA8
lA7z1zA0EgyGTdK7UwmYjIoj4bBFdsCJP14X+w6ncQKoF5hMTUGv85Qgh1XV6cvH
VEtO7qKXrMLDmf57LMahc5QYyRVjN2pDgBM2ex6FV69PYspFl9ffHkH2gvQSFkuR
nX2dSE/1mzrkMLMhF4e/dh4iXmcA1otrl05noCTx/TBA/Pw4NE0W2GOxCOnCcSS7
oKZcVl6ZLHfNI6Behp11QkGpC2R3s7tYdVPWvyelsyd8BsO8XcqxEig/2jK9njq5
//yT+CnYDyZ5YcR3R68Rq1yNqFp/Z5wmfM+VWsWCbbf25YpXkkucVP4FvL/B/zhI
azCwnjyNcfwrpqZoKVdU5RsF1s/vPahxpGTKVUyAMhkSHxQRSs1u2ICRXdhQQBeb
Q1VTgUaTfxcEBTfGtv9RWK3ageWJMm1ikozrDzrjCMHDT+S+OERDv43ezHUmqlQB
Mrc28WxMJZ+IQ44+CMb+VZpX8C9fDKJAHtVIu2ijWHWAIksl9guRskHVrLWBHAYN
4o4pEiZIl39fnXiDNYtU3cD5a+DLhBNLDbnZTYwjJrfryoYQpbTOBhi2MzE9VUHu
Hgz+PIbO2oR85v7JdsGyJvqDrZ1UMqLbOqCLHZvypl5Fq6LW13PDZoyn2CbgEb65
BP3ZxKi+R/0zzX+grmwkbuTsF7kSqm4AT2+BL6Qm7j30WcZr7Kcl3cbe6PL9Mbew
m3qmmRTddEkygjfuy3FuN22sVRKu+0FFfwMgz1oOm5l1Jzmn0xymi7Oj1+2ATujz
iibLl35u9qFNqNvG7JdR6WeVkHo1HP/8X7xgGLPgO9zVq0I4A/eg44KetIY6L53o
Lc44FUg3zFVxBGyULD0f4AKaJVMXR6Oa5dzhDxXWXlukBcrPQbcKA/PkCNwyeI69
EwZKvdlGvyusnKcjbRCDoq/3I8b9mafN04ibR8wWdDcsNoFLkRXrEZOUMtKfOu1f
eJ4Ma2KTM84i20Y3HtXFyPbjx3ifkIo9XzLj0VslX5l6QSlUbe/xf1vmf2XL65q/
coMpvAJweb4IM5hEuzyW55J6/i3HqFRApGXQA1fKGg4tT7yen8dNQZqgaZjrCnaD
FzaPVop0LyKi+ZCUHmCC7D7Iort9AhZj28/lOjv0RvjJNso0UOdQJkhb/Sqx/Mo7
uyaMBEAVN8+exY00fV/iGIm1Mpeik+0ECpLs48rsyEd1Tf2m9kmDl1JHBjfpbEfY
ek2HqHXVUmqEVZ/axvr1oSxv2QBqFBttV/ku0ZzXaGW7uxGR9BjrPQ2yvwXK/8TM
o+31RAH1ryx/U7GGfEZRtpnUG/bUQ5/mKT3xBofvn7mmeC8RDve31nl5rJbrjch2
iCUpPCcqbkDWjElOlQLyaYQhJxgTVgRgVg702kLtMefWSJXH+OgYBJVJ+y1yt5Ml
o87kD0LVA0ApXJGV1Fh3phNHDpcNsNOF6Puznru2/ZnGgNK5CyDFmKaxI4r2MhFu
A3dLAmHKsQGRL9ZyEqsdRFVC77QEquntYUOH6twj1U0EwNCnPknXs9Fr8WBBshns
j+xUvYTRBGj/JzxnqFeafxvSP8BWjxsxLWATgRuxn5ZXAezJ28Drj49xqxSM07OU
Jdh1xG8tmiYgIY0u2t8nA+QQgzomYMjleW1hn3AYWm/wOkPjQKEpjUbjAraWxwm5
ill3csCdfgyXsPu5lAXIj7SDeyU3eY04aqjSfoXb5ZM8pTeFXBd80T14HJILVb+I
tCO/2eXmu0NMG92tjht+nvQlyKbXBimQc6dQIp0xw0j0/hFtnQR1xuQJKp5iUvt0
yWzBnA6D0KRBU/jjdB2noWNEA9JY56bG18a1BKZh517peinjiUOuMVhGJcBDrCSk
YwIMitq9/5tS9TcoORkHiX2vmPIHR1FrJ7bmtoSbHCj4i9iixbruxV5QuDd2Qndo
G+RJxVW4ZIYsH8WpQFPgzIVg/0ChNXl/ITzM+j5PJkGixtJpsqkjrBt+TNacpmBH
3PyPIfo69WmIDPkIx0NQiHi1zUXLakPbCH4yArNo578WH/fx3Wz8RVNlPk4+vX2P
UcaLUqMwdzhSwEyJ6mYrZ8Za/8elucd9jpxJa7YS3UfbS12/vXdOoybvl9romTdx
h6/jSRFl+Q6tUspxAPbHDM6+ItIWsTRKsB9Twfl3iYx7cL/snLP6PTJNsdDcPmEk
ubn0+sXep8WUeDdrwAjOwbGSuehtT3GkCmPnjWk7IxwK4PIywmfvwiqAJ2UY/ZK5
xVsMiVVbKLlUOI7f2OivKIKY2UyBbaYke4DVaSiVfenx09RJBtNDoqJ880Oy/Kkp
d/9sB+loMiRDtUgEEmoPveGNavV6s8LQojXQXyDudSPJ4tr3TjWDVQdYKfhcnsLC
B4zypM5tVxFhul9JnXiapWT/fMRObUcJZpO0WH7DGkEI/m+Juh9xs2JLPBJOT3od
1r6QSVrx2Rc59+MSbHM2FU50e4j/a6M7noxPP/MukWt26EqiAT4sT1WRlV2nOTHh
bSm6jNh5ys6pp+k6EHlBuLApv1vEUJwg+1KL03LTSuiBfihQVaWiLqVMv/jlc6jb
W+HPoXUKUeMWR0L38kMVpYGqWVvZqGmOvfatOaqxoIncJItubkTSkWKzcOYiSewR
jACy6HELIiiN+gw2jbt78/ctiyRPuOOZYoR3V/u0Wg6qDJWntLWD74rky3Vnyy5I
aBjXyODGjCAKb3fxjEQiO97+V+y+zTfwNMDOPKw7gViR/nHEYlF3e2kePFA3LhmB
YLSqJRWq9aZXYmNzKOZX2GNc57PpzxI4bUCT/Hl53BiZB7lwnT1qGrmtpD/toFza
1SIMaBVaLarR/2B3cO71vdIwnxxD/HvnNOm1W8xqbaM3sNyeho6DuAyRFVQHPXBY
e3G1gFVoMcRdW6Lj6QD7G50QBhkICKUpk2wex4odp73Se2Bvnqo0p6HDTBFtMeJ0
AjsEea6OGSmU/Yw9p0fvPjIix2CcUKDd4GybHVa6n1wv+/j9MGZJpFdwuGsoxAR5
P9kcyJtvFyvfJrCsalNAgW8KgOPwfIJZ1yGaQIdSJoviO8c5K96HKs73uWLbGHZB
e+7IqQk6cY3rLLXidlmtmZkIvFAr8a66Ew9ZV6Mz1nZJNwKkygnwGEgqenOLnsq+
CU/W/05mSQvFNrIY6bIQYBZGyqXKjWXZ3XkTlJn2XH889YA0kAJodD+AbSu6ClMV
OP7OLbNlarR/CNrLy5eEVl7cDgiVQOAE8CXqZ5uBMqqvAjmU3x51BMY+6qHGppvS
XYNT5UozdwVxKhG1H2SaNqKAmuCvYISYf2ZgxzaAv/1HFQu3rrXnRUcz9IU3HYI+
FnJRqvoKMXAzr4xXBrSfuYuwaZ7+cQs+G9DLZEHe4WVSnB9voTskIp9qVLjV/oT8
+t4k44rLYNNqo3PK2CpkwAAJhF3Y1nh8deoZBLJq+9I/5TO5HmHp4sMhXrYfJDEB
pecJZy24HQG0QDPke2EaDLf6aorZRWFIKp4ZY4qSJ3kaLHd6fA/rDVZDh8ltgqob
/X29CX1oJL9WUbNR7AP3M2wbgcZlR6YHF/SNy+sMXIjp3LN0eIUXg59SVyrd2Ygz
blJqlavuxMwI7XxmWOB1T8xzNdS6lZPWPvfmrg2ith5Grn9X1swZ0AdKz+0Ll8Ve
PejzfQm7j7UG9bMpbgrIb00wvH8IjrWQAB1VwwlRSYVrGWam9uliBbqvVzMl0tLP
EhNE/RSI3zoU4eA/rXcrxg/JupvWGT9OefU57Q5Jb9Xqo5l9RUXVQAKlHut+vw80
eR0pCCJCVeWdjul14JR2fKZruFWlYFZwCOv8u5S4ooGZyXzGHpu7XQk3C2ieta+2
mLa8tF+l4wt2eje79tm5fi8tiQfymfgpEaZOZmw2H9oHSBUpq5jW0dhvokDYmbq9
v8UXyA35RT1SzDr9hbHUA2SYbFW8EUr+U1DuZa+YphBip2HTx3s2sG8UdlZJKvL1
06j9UZ9tyR1E/bqTSFwGOwhbEEBfCO2RH/8YuyXnRJ5++j2PbRss1qtTyLZVx4ip
wo3+NMoHqN6diUCN+ny8dkHtxeGe80t1psR5uPA+3UJggq5EcVTPMCiI2JWFSUEB
K3+eMT2cOxiNpB74CxZh7TEnage8/XUC947TKy9YhVCtUM5Jdoa+5xRIMpK+a+oC
G6IRbrLig5kuab9dM2zsRdvWL4NCZO5eidJDopyS0w8F8Ahhvp8l/5K5ifw5EEVy
e0LKlVDgYeHDfUuQ9UhOvPS0AdTSuWT2HP1WfX9sK0ZzuG6wf9DNiXgZQzHBRpVa
QXnCrskurpeigGRIZcCkM2FySzsTwzZSCSZWHfwzH/SmKDxxQcoaBo131C3MQtlj
pkBT3ydKQCLrHNG9hFbqWmLAzVvN5iZY2mWhicnUyarM90gLL1c969ST5pz+N6ce
yQzOBBPLVJu7p1OJv3MbO96FjXEx/0mOhj+Dc8wtp0UQGnk3kZ8h1TTi61q/A/xf
8hVQCOIFe6ORfS1ipMvZZQeuzL0vwKrffq4RibNcW2bOCzlqRqwd02Ka+IAaxnfx
xtJkLfqQ5irpYh0+V+SgN8RqHH3O8vl+My5/5+zgxIG+gYkCVhX3sAbljlV4bS7T
GjQFbkGyAYpu+8AS75wT4LPWKevojNynw8flxqYy6es3ysEatKhw5hIAUWJOZnoN
loFFR4JfSHIgcpSMf89b6rkhlwGuceCGlckNT5apUVGoIjax0Ac8VnzwnSWoJdZO
jYNz4stTU76ks77YacDAQrrr65xp4rXVLIWgsFgvv6u8SsthplWKLchLRY9jYgdr
4pUMH02TmbCqiSmaELniO0wejTn3/4Pm1OU3K10ihuHKRX0uIVTeNw+k/UEH6Kpm
oStQ05s93IMVKMa6nm4RG1RfeqS/uZA9sdc8NIBiQymj4lq9lgDSKXCQqEuiMpDl
/CkLTxyxkjNJQZTUfbeQlGpd4lTogKH9qBAlI2VERWtZObxYnqQNcTPFVzVRZTQD
XRzVnMoERqTghJO6yo2iY/PtDuwKMAgrLrTw7VEhZRCJ+7mYCQPUKQuty3ZvN7an
S4h3nw9dgD5HVH906QZT7rcugGivIjnNAnLh0ues1YEqVLbMPuDUgW+LUhK8805d
Ji+wMPXW2kNQr/PgPC+zvixpmAER1gslD3eTPO8h2XCfBVU2QR3wEZE73yEzuEfm
xwc5qDAZ/hpB7deVQi48xifMPf9BckYQ8Zpj++yxS9lI/izGuRxzN84Li/7i6mOZ
Jk6WYI66/VSerL3oeu7miMdwm2myyt0/OMCK3TMOhkahou80lHH4etL3BIniBJWV
+UL5Ot/MjOWjD8CzD1cBnhedpfdW1c3wOCrNojohZlaJFPT0HAaeKec26B5uU+Dj
+wTItE1T7XdZ5LHgfnmGypdgB9uIyqokaCZte11IIu2nDWQ9VsWDk9ykwSiCY2po
nDab/QLGvEq4dqLaWJ4ztL34CAyhXRD9E4YEvZmrnX2TWhfVvdBFVgjaSkGE4yew
kToly2g33W92zBKZeE9IUu5IvC7vprvyl/LkF9ybMZEOLK12S3h+Lsj15Wxwsrnj
3OKJICGb3yo4izGOx11KHr39zjT7XteRvQHVGrEnkYPrN74gQj0SS+thgz6IoTbE
4nxAAsm8MXlQBccJHJ2s3IzvOiOV3NRutU9ce9DMrmG9wth+gu7auvuzb7YOWVSs
96+R/2hlg/UlLzgbxidZBk8kCabZfLZ2/Q9EO2uCTe4zPM8d7hWnaFr3k/zEvcTT
mDhbUBZ3GmuKiecB+869mHhSjVXs2fU4YNAN3TXNoAprArNtdeoIHGbcaWP4nmcp
IqU/xoUiwS52PgfC1DnNJSrYInVITjayMR9vOHWwcvl2iblfyJ3glSUEi9dnHNNg
qKdfeAy7oxOsMmI+B1NYESX/cLP6c/3hLgveI5WbcvLDLkjb/X5NZK7SJer101Ql
VN4G2oOfFZx8l1hISlQtgZ/91Q+JCDRNaCCwDnRqib7sbiXCQarItCRfDjTwZdZZ
8wB0XQH9TzRsQwmyB0bo4X3WXjxUixxR1Gc1iGOAJSI7Vj0tBY2yftZW+WrNrrQc
oFMaprakloNs2i5kFe6CQZWna16l3NaZCdBj3RyHtLfcvhBq2jJUs7puxb59kdvg
d2LJBupZEVyB2spDRGxCDgthvn3Eu/3Eo9Db5NArcBwAmKsrmJ3UgSD/95obq39M
7tNrtkthKS2oHIbtBuPdDO6p5N6UCHc8W1Rj0rEVnQeU/RdBffVYjZl097/OXXKl
sJiPytS/iv3HXCr721LKtZZQLbe10RTSBIHmKasS73YU4w4MBMptmXvZHI87x5qn
0rj6z1ZFEpJlrJfq9svF7O/AzOcRTo0JMY/xr9O+F0FE9xtZAMJzNvynsrKM29GS
hW2DsMeZGZ4tol09N2tGYAdfr+adelzXNrArLgaVouXGPNnMczslFnqtmfOEWf/g
BKw/a5jquHxMOY/HeW4D10mHcUHbxteozm0ZxsheBMRItlQeS+7pg8TAufMSr5Za
8EdLNrLzgO5YKk7uXAq72m4PADMAvkgPVd33x7Dj9HRcsDA8uM5VV/bNe+ZaOmXd
HDuYHv3cqOFxJefh5VgqU8bp4NJqB+N6TVY+pZ0UURW+Ziumyw9X0nUpAcbhaD1W
MBcNIVPbJLriE2nNqdMwk185dDIgXKKdukDueBpHlMn39NROMPnPFxfmGXFp5CiJ
PLOfWyXK2Gqmq9JXYRY3Fu4q9SWvDEvqEY42qVI8wt7pQ3JZxvX3VdJK7hRV/4ij
DIFFFcyBDw32gJzx3vqZ5BDzkmhkxaFuHu7YN3HKM5GutGgu58Du25nLOeMFqpFT
/djT7qo5+ej5bOcRGfXuDeQrzKv2zsXp0T6jBuIY++ou9n1eD1n6AWCDlRTEYfCB
oFQOSRAlYii7qmDBsoIoiJ3xqsCcn6OLbsRykkLAV149IEbopzDhDdH3FElbgAC7
8shj41dX+lXlbarqnr877WbIC9IyVKo4CDX++e1YS+zlLWmXLkoppIWqZexPOb9Y
qmQTfYVFYiGcMxRMSYr+UpEPnzfsDBxP5kro1OnWczHpcE3JhCOjmf7LMsCKKi7I
lBgtaWT3EekatFUsbeTIQbMa8Glun2HZtyCgj4NJEagcOXXXbbqqpeCz1TEAeLwK
EzgtyFay2v2Vj7b2vZlLKGQusY6mPtGZ+bt1nUctCgT5aIeVUeqqTfY+bcVtJEW+
Fx58QHMn3v1OsAF6rXyb2m2JQTbYADu4cbmkA4+g/DBkZjgxHW9lClTLAfi1rxNS
3ZoiWlQy39U9C7hwiJqGZmpYnXsnpQXVd9+pa9MPGYxOsryB9TVHE/sJjVjTdEdB
FL08x2/ySLvkYccjIqURtJKGUvaZtOtwqDNbD1yodZm6iV0JnnlzX3yssBhficY6
Unk26QDKcH645nuzGZsRxoNRI3PLvOouDtuhC7losHCuSv8eUhd2pi5N5SzRpl6V
bjjP8UxXLwAWc2N1Q3FbnjWd/ymuTBZZpdmOCfkKzpGCrlZo5ZMiDYD/izDHjr/4
ilolivnTOt2DPLIBLjSSX35gLAj0bb+pX+Z8gIhVwmQqo0u9yVnWRgxpvEoJeydZ
s4HwxEJmS+7AototITKWgHDtJBKh14I02/H0GIT1rsSKRbJMNXRDOPXp8ea/NfUh
cg2XBRV0aavi/gUvr07PGzVzQ1hs9N+9er+UkyZ/yRy98+3bbJOEoxpTHD8r6iZS
lQTfBxHa62bhxDjgmmdtnI+//hq+Xt3n6YV5naoI8aV440rviENhWwVCk8eWTziL
6frC3cKdavKah77nuSS9LT1l7tSWjp0Uy+VgUutbHsISrSORYlxRuzKiqFl6gQiM
rVITXXQx86vDqmT3jog8x84ALiHXS1blPb3Z/QfqlRKfDnWvGvb/zbXCvHF6s8TO
rQfh1KjCKPjtKxwx3AQ149UVuEYa1Z7WYFp0gCkUpRHcKwC/zX39g7hjmT2gI52Z
OX+R+e/x4H3Vu7tx9wU5/hsKK4wHjD21GbmFCKmXEOs65kQxyGcB4TTQxIKASGQb
I4+sMSSDcrJY9y088ogVVgrWyRFYA8RbsGX0v5xeaH4ZkkZXw5AhSKB3jYMWXEyd
Taf8nTH6YucQuRs0sHjJLpj8kd8RE84LDwLDCnEQdHkajP1qg87pIfQvKE26H94+
6wQTdfWGvI7SL5rlwJeArTEOqCStlJRiYEAVHmH41y8g9SLyyKEN6toIYajpI076
MZEqIb9dfiPCl1IW87Y5jv3RtG+1opSgTGhPN/9Gzis6j4S21hZZcE2IgOD6nw2H
Eq/u50XxkMI4iTaZ2ORTCh/NpVa4m5Qii8PGBYLI9Mgnv+4IR5AnNPpGEKhETmEn
eOfUNhMSGBqb1d7BD+kOPg125NUTXx2MraE3UJe9h9s77Z2XmHtYIkQaKC1s/z2Y
Vxaaf83e3j6UahMe7sHbKS+FPPPK+5tkqKRtVT5TCiM1Q2eAl9eYgvlQjIgjvpMw
f4pBxBreWbpnJkYX/TROT6ja8ZVA5bljbr9MZqf/eA5oIBDDd0Gr2pF6HbwS5tyh
MXms5Q9c7YfgrIyqPEpfByaEboPloPuYANP/YkeCSwJxgk46QyBgVc/0o5vdspIC
kzgx5ixrFn3eXZqkHc4PZcLknJdLhprxKqNHd0cvgp7Q/HSUx97zNVNVrH6mLhzZ
UGEa6UP8b8o6FVIeDMLC36Gw0uay5ZWM1T7LXFPMj/qGns4q32UKXLTVTbkaqwA0
p2bvcqoF+fVT+yLcw9vQzNlYZZVJRcpu4cflecn1L+Jg7A0VflnAwcpSsUnynNSN
kG60hio0yDP1lHXUrBMRdQtwLrNpEYAsc6zk2FH6x4pVka3xIStmnpk5zOZla5W2
78gtcsQvALa3NpcM0S6W2AhdWjFhpy3rCYz/oYslqb2cSEDDl83v520nuSvug77a
+fSgtEobqqi1H/ndzsqvhJhntRZEkp+NLKQfQWn3TzSQ0Ps2sJKQLvVYGH6Ug5AH
ndbokJ5wRz9wLEgprMLxnGJkX/cPK+cFZDTkJLCyvdzwprHZzMQlmeyonN+ngkDB
m7Y+v/zx5/UVJO4X9l8RThCSDyVl51XSHm9f9MYWjZofedv5BBZodB2VWjctuLUF
H8rzHHUr92M1pGbQ43FgCP6wFTgCLSxO6HhApxPktrWhwo9+bvMGNq2OLiLYPZ8B
/Lh4tUdN1hu8YJl9x8om3SntdAgauJDGLt6lYvGBzlCRur4u5k5eAYgvnPzBQkSq
g2OJhFAo0qZ1szRZbYQ2ToVTj1/ZxIZN3tEhpnQ0FgpKvgXN44UoaW0jjmtH1p5J
LNIWEE9s8NnBez/yRCS4/0CSrBQ04CHRsIOinrnAwBKCRIbJgHOKGtxEpxEVXEto
12BBH8ZXc6Iairgn7oRisg62P+vJdM82r6D5xVsoy2jonAQPvJf5jTnm+wmacun9
3k8PhYozbFguWJxG7x4QqcggoWG5Er9DnJdSYbNfi2DZJtE/3cVT2md2eMdQ4PjF
RjDZRz5szmW6JDKMYQ3kfIeN8G8rHwHjGpnGOZDMYW23BCp1ZTwLzsm9LiMLHput
EIx2z8xN4div+JH5jAyB48ho3PtDXlUOtjRwik88YAkuT1OP3mt5YzKyESW/3aii
9JWto0PfUVFl8YH087NXM+mhxA5JY8Czf3cd1NCe3//yCVpBdPERIsIAOJ5eiOwZ
ipCymslsuO35M346X88mLKtwXQuntscNcxN1XBjwG1p9q8VAD/zX66+xjN9z411U
ar8uu2qbYTUIo2c+EWIcjLDkFaRw0UhMuKtu73U8YfMJG/oQLnXdLb6lyTOIAGuh
xL3R9duJWgCQeKVyw0SLjCrFc+soEcrIeo0KSfOofrTHShLand5yvrbnJO3VEKLC
HRkwrv/6YE3iKMmKv1cXMvQgq0m4P5RnjWBZEiggrop6bdjB/qGE3qUNd5xHVxKP
Hpqe5P58Bj0zra6+xKpG+t3DlhM1s6GzkH5sjvsbMZWWZuoCNn+H+W4lNcywbj6M
+dVfI817MNXjD4dCjXHi6NMTBo71x9LxiNMbtMasWtKUFEranLu1m8+cB84NjZ3V
SuWjxkL+qt87Dat2+BICRyuzwYbs+L9tKnh75ImYgy7kxl4paJ1g3YFBmqt+RV46
IetWYbJmlaykp5jp98x2tk3j94cqBGmbHNWexyTLeF15kdIFF0VhuJgPijAW6ha1
pabCifY3vkI+LJjUSdxMQJZfECfQ9+BVpWuUcRGlJf2xuc4D1JSfGp9RTtNX6o+d
nQUBXCaMXs6vwVcqm5ci6x2i3wTse2Vai+n5hKrHti4bvn/gP+5ATih5S70ustj6
T4KIbjuhlTjqE0KdDVr5Py4pUkraiuSgyb5zAUYwHEIYj06XAS2Bue5JgyB547vA
xEkTVa0KKQ9Z1jKljB1OGMic1DxJH8kWQv76cnaqBbZZ73j290lka8A3/NXjwB7X
fZtm9cPFHXWlxcejwJ8iEVH+D/wOH1ZwJQJXPJ//+7eGN6RG8+DkHowNuIyNdoYH
9WqQihfLnxDniWBtOk+ngqqYnyiVV0kXlWj/yegf0OPxvYm+mGH4Va12TbtJjLrk
UkCM4UAROT+O9/2QYJ10aaI0lxPuqEmGeufs+OznoJuyaM1FuBDBojnIhzW6XPZE
V9ShrY7Ees0pezCAwUx7ssaILJ7sAEHJVP+RbYosW2Db91lE2nR31KPfB3FS4Gf6
v7jYvxjARjYBcR7t/vaboZNzRCfIeBQdUOv6caUiZ+qoc2wHvumeVmLuv6ZFVJYC
nwOs0S4pyXmc0bdswwnOM6esNsQMd80szrKwsOtasXzynGXqhxQemT9KBF8+AXEt
ot5X4Ur8eOJoO0/LD9DyHmrRanIx1dlwOW4N1WIarzJoIOtZNA/Mt5aCly7e4Iip
6NDt/CmIlP9tWMa8MSy/5V5PqN/0aybhXO88F6oXFX0gp5bvPT4GKa7PcWTgpuEA
GKFjdWGbNb27Y6PNo/VJaXOXPzeYQ8TCGaGvxNshQkkrhNKkpSvc1YUIh2r2medW
B8pDZCoSDUyf5ii5mMtdK60Cuwr3nlU1uAhGqW79q0O9oTcEveW7IXR1otPH5lHE
jw8XG8Dm2QZRK4BUZb7rIl8sUkr6WlsW8Rd/zCDubz1+k0ja7m39B5kyG4LZph8G
tijJir9N9tHetZEiTY56AB81I9u9jACIIPhwG6xhET7fbTUZ9NbEsEw1dIUjqk/x
aumNlrbq/veNJxngH4hweYr4td0CVZqVkTvDEZQpSZm3xcPHBok2iDsrzzlybaBT
VeyDs3+9F3nwwZOky3snKiJKLau9zBl4eGdJCaY0CDZvydzVlrWRoHQftZ7JGYI2
mZTgj0NPbGthkyjOvtWvQxnJlmMN4igSj4zMe0IohWE9vqrXcqeKrUh4HRP7a0kT
xUqdAWL6g6pjF+o22je426MeBFwWuwQbhAfDNK7l8d4E71E7w8vSTjWELI0y643T
o88cxd1AyQqobf/tSFcIP3qwtQWjvydPtW9O20GJY1No/SIGW3L5BDBssNreZg9i
ICAIOvrTqJqhrOD2K4nfQpfay3K7joy87RFdxMUk6kO7TtxWgMBZROoTV3IyrYgW
Zmqh9u+Gjyq1ubZ7Wv03ow01NcNXD1roZbKG7sVAkQHI0svuf3wCGUEIDcZlW7ZB
YahTbUcbU4hmxDzQ5CXiC8mzB3bg48T6lwg/6WGN/HEIGoVPRAYoFjb+1rWrxzy4
mFi3IkliCyk1kha9DuAMwHbFRe+/WRx3wXEfmXtLTAou+2qbPAoLBar1zvdblFU2
RaK0QxQhyV5nsDx9T/GIt0jbP9OSt3zKFERcbWxwrwzr6ixrBt1sl4EfLb3LCZc4
QV4DXCr6yZxptr97b0wCVC/QxZilTpO9pJaHCFIgkm+pH1LC5JLReHKYACAeZQkv
PnIJy6jk9ZUEBtKplV+Wojqjy5OV+PnfuMbQkwBmdMgfW2qjPtEk1DRsJGZp2Q02
mpEV7M7TzA1vXc63GNOuVHm9XfBM/AuEyZm61kFzwKoM99Ek/juPhoimMxaNYuDj
L4Yj+E77aoFNcKXKMAVwm+MDdAtupOcdDBxLkLUxdumM0Pcozj+k5whexG9pN6mT
VXvjQwdDFMKHhZmP6bQe5XerCdj+Yo9N6/w01QgJHcJ7rBFybVJneXvVCFwxANgC
nvx+BaXuxg5Xj41UZhrGFWyHwx1mYaCNlg1vlBMtKDCMf6q9MImcIvO8jtEK5LG+
msw+uMw4t3P24UN/uvQIcs1mTA2ki3HoNZ8v1JDEIemxNv2uf5/VWFFb0bkoUjB9
SR0aqUajTKBcndCIxZVpfvYFjIY45ERa5qVdRsA817vO0x8+AaX/yWkY9uG8za67
tqXIt2XOLa2MU5gKHP2IkwA82BjwH0BTBvfuOmEgcFOvG9X4Z5Z8W6XEVWuOHEtM
anDtUA5LR1zukCvEyR5CL/MQ5KeG6FNpxY3IGoanmnQjmKeItTxZ6SnMbC2hqeot
ZMj8961hcLbqzzhDArXa4L23V97c1WXnqazPB72/LXA0xK/XFp3qNyJUPNBkRJ01
HQF2nSaql88NzpcSttfc7svQz+W6D/BXk85M8sfCFnaQC4yb0gc4zNOUQLSM1cnQ
tH7v/rKMbE7A5AtlHyD3YYh2o56G/Vnw1mlwgbQtekQmeYwbu1xUfi0oh8iPoW5/
5NG8bAlsIceI1fTiwlL6BrRx4gCHJ2IYk+ejN98SfEvIo81hpDFrpP3HMcqPm/SK
IcySSbHDh0aAh0L+89EIjL3/j0hXK6r3QthezEECwItqpDAinpP9VtaImZICLpC6
7Yh/JxbUta8J/occG0F2SN15sBYrKztJ4/QJ0aQLYE64T2JVZ4PqjHwJnukMB2pY
CfE7/Mn5AbLhtDSQJeJpErs3bAKGve92POpmuqOGJSyjlFukNhi1ziqR7ol6zwAd
DISo35hT4vcio8pFi5mSyNYUHXOyQKobm4W2DPGa143UJDU8JfCf4M6qVvSIBtDk
c0lx1LovXRRn0UUB+d46rT82l4OvwSCuE/ZQzEfa/Zy/qRNTkaeAeiXlOMNuFkPW
nEXqGUzDJFP9Xzp+zGuWUwezcgewW+XqY2Eg1wW11stN6God7E0r75z6R6CB1h0s
5wfqMWv8AJIb6gfOYTcsDKCYJkW1/b1VKGc7titun16kv26EXIv1/CNBVllCMUAX
3Mp6cEWha69GSqRItY+4qaFTMIv3Xgiu+BbVnB7akZSHCxSttJzICWEbrFoiorcd
ucti2JVxNp5/t90XqZU+/QPUd4kgAocha/QEiynA/LQYuzn4DMUVzE3aVmib95av
5wxK9kE17rZymNsXUDsBzm+J/wTBddxLPNPTZFtI/Rw4MGG9As8crc6GGdRwed+t
1swWt7Kdqgp5betcRt05Kbzr+EeHRYbca5O4fB9gkuYHWPiH3ObPrx7EXwahXd3A
lHLVX/2YHQoxEr7MmDgPi+ex9X7CN/8dYkREfFG5AQr5Hz4QZWWR8s7nEqNgou+h
pjg53fp05J+0B/X4uKRlBa3N9dODRsjMunQmoetY35uCpBxDBkaAm35OmLaMgfP7
YoUk/sRjlLAET2i7TW6YEk3YaRBqFVXfaoXhWtUPlhemY/Q2GR4wmnt6UB8TEEV6
CxHfZMR6/nXEeYLHdL7Ag+6ffnJH3IbbdxU9yU8CDfGAIY1OJpWrUxbeBrm9zN2T
8stmU5y6iMsVvoRrfJOu15w1inrMTKySK/Bby+Ryzq//tTe0vKVL2sQpceXQlkyO
Q7nEMhDX5iw1qA3w+O2eF4izjuL0BvTR7GoYBnNohcjoLV6FJAJ4axCrwF8E7YPd
lUn1pMdQWUsMG+hyj+Ozm8RFQJn0updW80tW6i72E9nMlP/xHDr850EBakbB+0ij
1leEb56ZlYPUPSWOD7+Knhc0JgRQpYOfqagpxp7bac0lE1eLSvAiq7Z2EIMUtZpH
kBnzAAD32Gwa4Bg/dgapDy5oyxNMAlXGxDaYiZkqgD7pfbMOQu+RSY89jOAyQEDz
ztL4vemLBgO2tTaxAPd6wUddrkEWTpgv8ZHP4kgobMFGvgq1mG8CibAxqeWJzbSR
rDImKzhrdwKL4gpFrgIFmuGJ/W4lU5cR2b6NpcvKmgfq7dnjwrEVwAJxhsvgGs39
bwXdiR0NOoDg+xyXkj9OBuAHxqbvBdQPeTFtDVz9V7NghGpyWP1hiNDE2GAhg+EP
PLLrJmIaB7caHLyw4RLOydzwxL0aGDwOJmsGcWB3/9/VofJ77UMq+IKnyM2J2G5F
12ft+NQ2HJeFcpZz9DWkzsK/5zcBJqTZhEz9sgxzgrYAXfvXNOfURw9ULWeCF7cx
pENBCuoZT6U26aVrzozI5KfsYGiBrlCL6QwBiWOIvdPfPB0S2CHgUp6k5njq9Qv4
fEqfDKdQbDU4gbv43MnTdh/jb43uPN4OjpKqFI4yPugR5tB3ljOXvzzQfmu5kGjw
q6ooMDj8G6aLiEAAuiehuevVajKS6I27w69tg4mYchLmX/zBNOsC+9LrbICkVepy
QJP6zGmZBRAcVecQB7cwA2DA8V8fHOMw7tEBFc4mrr4EEH6FvbllUHJ2qUGwK4LB
rmJJh9TzGthHTb3U08q5iaalIbpLDASwrITEJo4aekFZAL/ojlcYIbLlPaAa/wq5
vw8rmYxiVgU4Lzjl1UXVFkg+sJwHVQKdQ3vctxUvTDNtjnOZRswiE9ry1rDRADik
IWaE1xcta8Y7B+yuNJCgDG2TP/Geqe8LAIMy4UvIxeeNVZFuRcVxJyVPRyThxpSt
cnOX9p3eccG7fyWo1QxmhjMZAbK9AgXnikyPHDLZ1JglA1UoT3gJjQhTvQgCwlnv
mismJTq2KOE3ZIFhSpcR5LUMCjmfz+FtMAb356p5G5Q2eVvsy2hY5fh8poUsBLIw
+EuljQBtcd5ubu846xhO+Bn53BbpEgTTxc5wW1IdI6BvCn56u86nfP/9QEG/dehw
JD1i9PFnSvA2oYcVfpKQ79dZH9Aa3FMx1RBZAbiiRnXJGJ952ZhBoofm4cIS+uTr
A8VCt3BMVRV1R7rl3wruJOZlAzPMc8wqY5Z+hTGwxvOQTideCUrh0Z2XS3kKL+8A
Lhk96bJpM5y48E0PlqBV2rwol5lMno6mIKKVWTSpXQiIiZx9kJqJymbe4s/nkSqv
est9VO/O7SjfmXEGBtNmIo8F40Tdn+NuDFhF/YGzbXdgRN+hboWCPRZRNwbyCgi6
NSfvgc5sNpPqXmW86J1wP3kqHPiPWhEHZtlcARfOPRSBsvmiD4N5dHZLoLWIvbvm
ML0xQ6SVp0c174RZ2Y1e1xJZRpNLKJ0vAsPt4GgYQVSGb2Y9gOvHyOUqYePWj4OO
viLFG5jvcnLv4N/5slpC/GvzM+2S8/p7DEWuXfsMDaKXc+Icy0G1L+vBpTQYLwXi
9na1gZBO7XwpWTSAJsmIyRCrhVlfmAwPFBm3F1H4p5y6KV6uwRrB4iQWwKLhyWkk
usE7Dhdg7wbm2XooBuFLf/nK4byD2FbJSHvpFBKVVYR6Cr/UYA8drMfSsUhWQXMN
UMtxu7kCGU2McCb/4oI7jTVQwWvwv2Pv+ogc80C7GGwZC0HPT97+dMtb9dAam3G9
kbhNgZQBoGQ9Svrh7H0kmg5i7tqvE5faDhhyQ1o+o5p9yQpAAjYOJanNaP/TR09p
m50iPw7yymuoZuRQNB5hmvq9r/7Bonj3zaKKnYcVb9TcqxlskYyn26SZrI/hqxAW
4J4vxovHVypHW4V/yCxXhkJBWeNDsCRGFmn5238f6WTdNLhhSXo9ipJfWpMCZlkA
w2RpVx3yfCujUd2ze70T0M/ci3lGBrBcC8bo+dg4NxBTXlm6MnkPccVpKwKrgVvE
601m49iu9KNT4Uryuwh0KoIIfAGxYRNGbMsUTZycR13gXmZqXNkUPeJRamuOQ+RC
ZgO5gpzAjuOqdXXBjm7PGYPYRciJBsf+8Qp1VuehtrkQ5nvU2P3ezYrWGoFdDrWr
fBqwO7mKAFe8frIFuRmv/ZvpCNtR5h/Dy0m4T/mIRkFN/3gJujLIiLCAwXt9fAPe
HzbclLDHj6eR+t7Ap2I/ckonJ9pkIw1iC+qQzyOXQRX7zIScf7NEP60OorVmtj/D
NLYZs/OqeZMeq/yvddCRA7wtBBBvHuSC1IQi4bFJ02aD7mEHhGvFABzGkOg3Aehb
wo5jlPVo8zvMLt6eaYcN4TFwyn4nzjKzPa1EEllCO6+1t1OOPuUXXSY2OpdJARWd
ZfTSUO0v97ynUurCcrK2Z30lNFE2WcsDPwWvJitDRiv36BPoy2FGWAZ6JwFYBi+T
s9efR7md/Jeruhr6cI8CX6AqHxZmW2CyHAgJN4KUgu0Z0M+X4A5G1+K7upcqeP+H
Vcl0BUdPDy7a38NFzUbno6JOABGfdQuxuFXPVIjLOnP84xlrkfug1HxCjiNw/SU9
Fae0VgcF7FOYOvK2xMOxFjENasj9cxQPo/S/Z3OLJqh0Fucv7kaDgFWiGspxqd+T
S+VvNz3PchwsWbzwWnEwk2rfGKqmx7orPZKRbcMcEtQe8tWWwiCPyHQiyB8W0/ID
k/yJz6drltfWwCqb+gtCgHCady+KpSqQrnp4NPbY3DqSIvX+NTdnaYDyfK56tDL5
QP2gwCiqtUxulWgFUaxPO6L9Cc8e4b9uMc22CO1/DaZL1Qa3+NhQTWBGKM7aKRvQ
CJG9zRtkkAjeIaYrcmEm/IQAwA+GzqGAUsqOO0VpT6PmVyrC6J1dOFR/iGgtBYxd
AmK2G9wwDaO9NLVKTRWGCkyWh2IgxTkEZjb3K/hmkek+3515nQuzi/WZK2CE6pzm
lJnFaswejUJBNhRVivVcs/FDNg7vqZjQOlat1xx43WzLYDrBN5FTaP3MNgsdmI0x
EnOwszfcdDENUuzo1acsp+SrwavHRhE815a/Y2tn2d/5I04V4a2BQTPa+C8DsySy
0WJbJQ0Td4837RzeRaEode7LGV6W5jWTWP3Blk2b3r/j0vIuuH5lRzPvPSOCjBV5
RHxQ58BwfepIgwfIlJA09m8+4R1y/BW0ZxsnIgZFA9+e19Uy+w3RYFTyy3EAvJLe
Xo2X6zLn+DDhgWJNkYlJPJozNnOYI20QDBfAAuw9JnRrrwAgFH4mLC9+NPo8SjHF
bFFsINBTYQ4AUZzfKoWuWltEQf+WVh5yFWtfWv2DBvP4MIRJSC57KA2OiIIyzBy5
lKo4Jeur0LfUDIRQ/FGQ2oca+UdGwovcAqfUCUu9fUCpDdPMkDTFJ/vK8+8XAxIy
kTFWRy+ZL85AobcqeyPL+Shpg6EYGWFIb9ozfq//XkKqS14T3gJ2LcRf9OnybadJ
0gddtZycwzkfYdoKTL6gxd/bLdMyVnWTNRyPllPMVdyqC66kouIVdEspB2wkD7lK
yBo0zqmvy2k0xnii5sUYUFXdvah9pwZ51Ci5YqWtFw53D0nDnKlcTE8UC0K0Vpq9
aZnQxtQExk8TQLoLd4yKYc5JQAKNfuEusz2y8JuLDpGVtjbgxUF2yvZIS7BO59/6
1I+wl6Ql99LomHLNk1Ob6toZYFBgcFTTYLtJy1LIDHwrzrgnZEr+hB72bKz/8o1n
jkfDMlewhU8qjjmdOQwEQYqBWUlXn4rboEZDJG/GEkzoqjC6eX9m/t2nvA4SPq2c
54kXBrBa5VyGCj/E/eaU4rvUdLcsHzF4G1eFXZ/BOmX3K2ZJzczG96QmC+jJD/fH
BhtG7KaCfnVZXC2tblEqSV84qHr0coE9/mYw9qRgShfDaBeMPHbsEj6+6OW4gWhG
MK4NGNod+Y7QzOQfJtqy5EwVYxeM3TRzzHnWgg7w2HcAvr9UCDZssTwsHVVY2MzR
JtjV+S6VqT8SZ8WmaT3Oxa5FVGfcCEP3JyptOHrhjFi75pk+0g64PVG9WirHhGyT
w67NJsrdYwQoI39pd4Xqm9+ISc5qKnHG5bq3IOSZHrN08RFfyda8glLZDio9juUU
OCgT/a2t+2twZg3HSjt01nCdkSvskoxmeYF2Pdr9vJPu7//n5FKdy6NkYoaraZ/x
pDxxFCO8NhrkKH0CoIFn7XzEiV+tOJL1aue1MTkflH4em7o5g9661zfAoPRMz4JW
BuzNWmfFYoQdGYauLlVVQ8jh57gWafbfyk2zee4QD9A/cYnkbt8cbLEukcYNo8jj
vLmNQ/W0NoIlj4oizQ405149dVm2dO3kvoLI1yYJCnivJ1YYOnr/9WZ0Vyhv9TAU
q0EqNKw2Vx9yluuLlB/PkFqM60QrNfjykbZEM6bZWUmeM7VKzvXKDNdixLmANgBO
vmD+VjmPTvt/RoW/BxUIrsyz1FxFGBnO4T7lgxD25Xz48K4RfQ0vNjrSLr4PUvVJ
pGk278mP9PTf973h00M6MDGdYcSApIPHJ+SF9KHWHzl68dKdz4bU9zYsZ0h1U90o
vDbnYkii1pI+Fau1ZfnnHY/RxMCEtt9Z8avne/6WqFBilVjwTNQDi7eZVhCCCLpA
LcSZfFI0fVtspSgB86/RR2FLL9nmQXiZtHSGQxa8zb7+EvS/0f2LKO9uhn/9rMhR
3L2Nxpv+cg4r5RVL77y6JPCVINZYmbdWjGT/qstyvnHTwMTX8EcWeJIRcaE1mAMi
DEFzTnyuri/0MfaSf3xP1pw4liJ4olyumDhsQGfrdAIpGYm6esvswpbEKAqOaJw1
kZ5tI8hGJdtushwwxmIk8E6plj7mpaF4UGUysbIT87UcBXh+OWga6G+NudZQwQwz
Ob42sw2g4LeNrpZe881TGlb+b5RfUD9wHp869uYl+/nThTIoK5yt/wDQtyIskFqz
xdkr4pphk/ZhrotrvhLjBGDvIH7bkKO4kYDt+7XUrSRdV3wSUETd2PPOv90raYO1
F3UXQR6U3KqE7YIpycYZ1d6FxN+ihpil/O+mdt2A41Fv3oUye4yBU2G+ZLQTxVXC
bcWe+B7nPw8AG/0eV3AdE1S1UYcdOdk70WjX06NKPq4YY0n1EcrOxo3KqbKL5jDR
AkCcbTfz96xJz98nvF2PmZ6N6Ruc8qD2UGjQ5v2euAOl30GqvjsJzTyNxq2ZnJ6x
NQiSG6WVHUfBak4nLuaWwdz96l+ys2TEnmLJJkWG+9/J+TOuFc1d+IH1pZZPT6NA
ULbWZz8dYfHOMlukxU8Pyqn0juqUatR7d1yR5C+PTSbQXI45HrwrKKhxO5XrvmL9
luf0ZE8wqSiSnfuz5Wd2LPzCLst2N4ylJ7wHwzWsrfu/n/dTRjwz/fVXj5BsIPTz
pfNZCBlAoO9OTyYivNTcieMk3r1of5Sm2AlXyUNzbzQd7k7JVSpMCxBZo7u73NzJ
UwJfHJXXrUwSzHDLF6gZVBVwqZhNIikzmVJDks1ORDXkKlea0Zxtr0mYtGBsvl2w
kdEpVkpUT3+ANIciVZkizdzi2/+oNvLd7U1PtRezpwqF8C5cyJwtR6j5pJAzUih3
ZToCxVtiVIVjYIFYDg/NJ3wO90kfSZtX9Pxx9LxJeLMZt194fNBC14x1RKFsnM8t
zLjMtM+zI07NRmJPChMOLTydY+3jVhAsTQwmDgC/Nvy5W1A+J0bhTM7wTHb5Kon7
Jz674bTlNcwIyXZzWlsWE8qbADHRAP/jjf11S4ptmC5zRFeZ/gzEqE8yDanl1/aQ
4beIfxA3LEFNI2QyU94r7O2rkY3POKFCBhiwlEgb+Z6oJrIC1QBNzxV8lzfRRjNt
ySz1vwidxd6qm3whyPdwH6Gd4nTeEs4xe1Yo5I2mJApsfr7tpia+AQHqWs4vsGIv
+j8US30GPdNqk5QZ07S4iZ8c5yTbNmnlDx0P0gMsuaKMIX3vasgx7LWQJ5xgNxRd
nV3GtXRj6wHJt0iasMbUAgSOHeGxhtDjvPkSk+nxdYKgVjXNyJHSIee9Bg0Q6PQv
g2gzikCt2ZUVzFe31chn4Va7gpGSJfZdsUzkzDf2vReHeeras9hu/fcbvsfJ1Grw
qeNQK+WEFWievuNHMVAGA5ZN7R4nm103zhU3ZBBkxi5DHU3+K6yTURNTDh+pLWgC
JylF7Mj83oR1IewWHucQ1mCjzDqca8dah6GzWZ0ZjVR/Oo03/NMm9eVp3Uq5SMhi
sgH509DI6iLMQMbxVsjJfJ16TXVYXlvydfbbZyjmNLcjrqosxParPuvQNFl6yMV0
unWc5360SeaTj1crTZMRv7U8i5io4l74GVe+rZx/KlMLBGL5dmwGt0lR5v+GPUTC
g4Vt7OFqJsEwuZIiHDGp5SZw9th0P/cnujADViAFAVOfpBGcPjWAGGdoOzjbcr45
n15kxglH+4cIy+bP0Ks57yNSCZKc/iwpfilYeKsJw5ksCQ2SoE4Uj9n8JGhw3OjN
lqU+nn4B+Hg9pIVQ9TQcPVTIroooL6o/eiQaJGb7VO0utlOGPr08nRyU3Tl5ReQb
TgF08GnJny9MbDArHG9d61BbinlYS/VwfJ+M6p0td1pbpm6XXUFcM0W/lepAdAJO
Nswt1mSZB3O1wLNDu2QyD0ekI4M4cZCo+xHWpSHxLwdc+rc5FW/MYL+qjWwwbOzU
3WA/SAGaoBG2h2Z2t1LN8dU5X82mLjapNdo3rlFkVNQ1TmRj32wKb4YEj1fQbDug
SOnz6iBphAciK1mXOk7gHX8D784Vplq4YeLGS/f9l58k5GVlo8KAudbOG7Iyi94O
5+LFBK6pymz2GRiK6939svOIbbEadw75EbtxKidtrTmjC1JUZG+CBYTJb0hIFdWb
jSn+54gwlp1sT6duapFDNxGq/uvwF+LRtftjF4Rf7aSyL5Yvad2cZBYoSGHfnRBf
SG8hDUSMMIpWPEE2YGMsCIVut127vgr2H1l2EOj0DuMKTjPcWe5rhhzHOpFFI+CF
iSFqr3KakaTY15qaLpn6vzXcbXNplVoTm4siAPpk0lAeaFhjisjGNBF/YdlHVjb8
hFqLZpfcjOQ0P+AcENfHyMGkllUR/Xhw5U00yDCUjWI5oj+8zRQJngJJXoitdimS
507q5TpJXfdxHj8m+nH8Rz05d0FfAaee7+2brbqdlHbh504GwmN37GEe1gZQsj3L
fh/jJUE1DQNXPq4jDY1TdmFN8YEXAM4IYJaH/l35aTdYvPqJRR8aaHOzp4XI6xFZ
0xJOMJcC9g9lSsvYuHkmN3yGF5vfq3TeHR2+XQd+m3PvXCohYPE3EaHQzbRz/9/x
5cYZ3XR2FcQm0zCIsKZOAykntu4npKs7gt/Zo7C1tel8HD1seeTg+F+XO/kHF3jv
HNve7i8Cf7uy7Fd72tCkzxu3QuJnn2cfmMS/dnZEJMyJbn9BeBV1hm0phwXZxWRX
Jf9o1EvqP50vsNYbcbJEPt2+X4Dt7zTjPKr9PMbJs7bqlKg7AE86Bg6Ht6m9yZaW
A1N0hj5lReopRCEzA+LZAUs2XUspwMhCLndOK0nvoeCKBqw2zFDJz21YQc0KI/cV
SLk/4iuyKg/LEJoKVgrnbKrfXmubAI3Cg2xIpiaCGT2wDpD7DxiShTws5NdeZsP1
u/nsGhKFn6c/cckXfLsocy1IujuRajBuN/EBCZZT/H0gtF//d6cpdCbTtORFCH8r
dDxOsJHUE7wZ9um7McyB1Qi6i1dMZ5Aa0KfA6qqYFc6QLXNaCKf7wC5sTTeV4hf6
Jw+eG6MWS9TOp2CF/BbuidDdPW6WXVV5PeHx8E0DVsVT6vq2jsonQtVJnjNwv6b+
j79s6F1KfNZmymW8CQ7lLKnW85TxB3GeEYrdGs/WGKKEFdHX6/pxlh2QWavAsGdY
fjMZGF15bwBJnC4f5Id7TEtovpZNBsID+EqEDHmn7MDLF9eOpPgX8nioPzpFXNUV
e+/ZBlL6dpwid2ZaDIwxqn8b5VyaRdCWEkIMO96sKU1ltJe3POyiWAReYQoj1LhP
qBZUKeEYjWKywDEtlBuCi1mj05P8/ncLDE7Xw93JltkQnEVxNcQAcWWanQt/j6PV
iVBFazQVEI/YOai04ahqopX9XROC/4xS8roAc9vLewM6Z3XXz7EJBk8XI0J9Jbzh
KIlNyKE+sUdSRSCeajBNHglv5OELi3yMQJ00Lkudb5FEZlj5pF+0ShAbPN6sHorp
NAFT7U4DIfA5RCKlYu1QfiOyLd1sj4ShGjNvUzO2BqUfIUyyObFehwiBMkKFV8Al
M1XGGF7iQ67okOMPjWDG49SkSxmQOUPCcxG8I4+qMuKKp1WB8R0f0+qY5t6YCrDl
bbwfYC4Fi6EgiMcWy2KZgrPbFubM3rOwuDyAuii6028f8jLPW6PA7CDEKqNshN/O
5BvF+ZLhyL3AobrbH98Q7I/0p1jQnH213aPg4qvuArspSLr+9/wthdI52iJHHfVa
+He5FkauZKX2e9ShYlyqtBQxqtPSFknIu8xgoNLALprJMkP1JUdoQXTIGvu+4Dwc
ZAioo7ygTh4MENpx60iCzj4pdJA1s8zfu+XR5w0OGVrQ5UiftyLKGsZ4s4g9AZMf
jseTtS1zVuEOneJnazjfh2oUTapjC8ZyaxDc7TDbOd8ekWppSIz256FQx2HFmT/u
xksCEKBGSSQ1AFdBAtA5SXEerbCqGh76a9R4p452MsGe4Vc7zVKMFNyrZJ1HDi57
JK/iBxIs2RYmIHF3/jp6czIGPEUUifSTopKPPMfY+IifU1kIhqZ68HPtxmwGrdqF
n8am7CJ/PTOYW4BQCiZrYj+N6GyMgbsstmATfbD/g25wFwAQGUBMGMCpAJ6RzJ9A
2fBZ6jHyNHgKxYoIkzEmKhzY1Q2mzcFZ74SNlvib1Um7RSVulu/uPB5Ne/ca3o7P
uSE+Wq5GiEGkR1+BIzsZrnFQ001KSo7gn6mBJWqBmBQXXIdaWvto1i/8xQpA61Wb
5JIxRc86X7waBloKO8aYCf8cqT4i5linh+/DUDf1an5tpsCFi7AOqjnVsM/XmI4M
+MK4BNA05wQLNyRCyqyJ/y/XWMW3GKBfnC3wG04qJlT1Ca3oZzZjDPxDTP0URMAX
i4Y/sRQPQkEIujeRSWp/hl8RALFLrZmhvoQ4tW1FB7FqXEDEV/CD3kuGDSpIckuo
YtRQbC3pHBEf+HlzMLozx93hhu0/acs4kbNHUlzfPVdf9qFaE2fAa5VYg5Nw/Gdi
UEHmnMpTpZS07CkPOnZhulIkn3ZjBT37+fl7qknWa0W0Tc3nqnq5M5sxmSn3cemO
Hq09SO1HvRs1ti5/oeNYrXZVgfGxfMOXg0WO0N+u4oZ3b54AnXo+nIA4F6W0Skk8
2MYdDySKtwRJ8+fJWEbSOwxr1xiIJu4Inu90S7shxCPg9xbn1dxkcrEgIKxcwxyO
+9QvYjB1bNZW5aASsw3+8t5GNdn3YKZnkALpGXOOYDQyA2djwQiSal8R/gkZ4W99
ozo24JwJB6MDEoiHC2ULiDqLIIKRkncQw0N796BTnP9hl8uGFI2/aRlgyEvmXe1H
J7WONFrYtxGvjby0bZFbY74CzBMyShX5INPxIoRW0UUn0V/8reHFJlm9R/jlV/Y/
/lvLxbNEa2r38H5xs/uxhmQyPz9G5AObyAFdLP6I/pQgWWFbe8brlkx3wUVHxFx0
usoQTrHGrVPlmvz0Lojxl3tic0Qw2R5pCMXT7rCp2njCUifTjHZMmq62myFCOej5
BH2O6Vky66oBXcVp76mPjXQ50x0ED3vlCqEktWTx+J5RE8kHLvqCKL9PIx5sh7uR
qaOzuD23ZZaRCke19lMfUO+BjPFYs5ZSe75VFDLvOK8v80YCZmFFWDIOAr3dRGWv
NP6OOhpJoe6KZrmZkfepHF0nzCW8bxpCoOdZra7BusheojEaQRl7N+g3DJK8uM2v
PFtvC4Bd4dC+B84EMXgtquwDb8ToLlHRw7cao1Kd6wQIbAbpH5tNxGftNjENKmQ+
kzC+4plUCDIX9ayIipLGHkJE8rbuNYZpf2fEPd/QYtI/+qfH1PMGgTmjWMS1zT7j
sMCuE/5Qahf9D4JDmUYnbAIQsgisBB6QTwPmaJb9ZT4GIbcKciiq7EmiKcs8sEaJ
p9R7jk54gBODS+x2LG4PPGSgRCUJpVvXFgxa5OlDT+T1lpkPl9JyetKjHpiMaUU5
oKS7rixgBSiVdBT6E45RWDPdr/srL+CWX9qrEDnKcNwd1sRukx5BZ3Go+4SanymL
H2ylT1Dt+GxxYmyNQtXz2ADPmJA2y14ndXZ0PSmicRmAy8n9v5+yzlJhG1O2B6uY
lwmtGq7L1RaAr5B6d+PqYjKo4gcB4M/KQSCbOGfOai1QwRt0Cc/q4uWGgB/+vblN
nAHPpWKN5/gx4E5b+hvmAHMYHKqnuceRg0NEXCwaOZJVOx0DdIBtESDEM6F7Sq1U
LuoJ+otGIZKlAjVA8p0kUyscyS9i8cfBiiir7xlCNbDbVnY85d/noD8yf1WfC85Q
1xE8Dq3bRDJkPV5GYYhTYuu+UodYrAmCT5DGWotLQ6VhTg2Uap5dn5ETOhhMHwIf
OaiqMlowQ5dSkfAYdSfOEEnClZs+FWdvj1lOiG0hA7YPqAbWwwJ5vLABqdiBl3vc
zJU+IGcamMWGASDSBLsIVXLTs1FamdGWVoxcFXNQzIU8iehLZ2Qq7MbNRQjL70vL
qdHMVQMOnYRT9X4zmNHN01hqlMBHa/U6lEk0iDg23T9hNTMG/4/7eVIrdvhHgwJk
4VinaDqAH1MqEYEzb+N2+Myycn2wWrubo7WfVhB2n2OogogJ1CFzCxotbiU32ZbY
QnIfaZBKy59q1EOpC7WxdyqWHrTi5CqQfetxRgAFLKKMPHoyVzKBDOvCHT9Oly90
8m2bvEXQWvjdUSKOftIOl8Gx7Spe2maBHbwN/orjxUXPKe8V+QLcFo1OqXRikSED
GANUtbj5f/N+Fs9bRITksZwgdORf15EVS0uZaYFTFR7idTfFdtwGCkJtfRXkh7J/
JB1e6GZUP59dnFVfrrnuxCF//i1Xy8xh+JJNP+b2DSy3vu2p/posds9IqjGZO45b
pkXkii+tAW9RXsYtgUMWn2plFcAyTYi2dLEuvvbjOCcg3Hsah9HgUO8sCMBY18fA
UZQCU5p0HM0rQ1k828d33BqhS0Hx7FGDct8gWCE32Epk2kMHcAqtNhiNem22J9jb
xkXJ1hj3Uf0lfC6Ad4nWRPwSMKNEzVozVME6tbCJjOHQDwGLYq0lZS3b0N3vXPYt
bzkfAgrNkeSzNxwKJxq2aqqLCh8bZmOLnSQft8WFqdQAYYLUzI1Kviq/EYSyXkta
7h0aJfss/Yoe43lFoZU2uQbzDHhJzpsy9v0u1zhezgosFcMrFHRkO1gFKT3kx0XO
idIpbzztix3xNeiqX0DGauo35jUmMbpcPBqRXBYnpWRvVzcUXvrVpxUkiLTfISDR
T1lXG+TcNNKgIUFR3+o2avM3Bgm6AuJDw9SS3w4yPVILe+77HIJ27VKkWFWFgvti
R9PivxDLVGSNwDAxkaZ9PapXiuXr2wb+Ekcfa9MZh1PLO5QRVI4mwqxJx6fJQL1c
7iliOAxYRi+2tgiGgedYDfzyQAFbrI+nW9rNHxIseOPFaX+ygosyp+DWM7t5eKe1
5lQeOajhI4SZWFUKfxm5tBNW1fXjez0PfhlL9c0fVBgk2eTB9+KvswQmTPkRZCDy
SQbttMyEh4w6Q96vqaozWcwSzXfK5OoYSRLEfnUBZM9hh0Ff3ZaohmPkcO3z7EE3
hf0Cakhhrbp3fRFO7YwATTwNcnWLanVlH83RoX4W8g0RIUYl+3QstLhaNc/Fz5u5
PTozDKJTWiH5XjjloFrGGswounELN8aFuj7e//8fg9dHaP8uLX4PW1F8NcZKPWKW
MmCmVTo3HOyzmW75QHpiZmrp9wqBVv7LlZUGh6jCzYbHnx1qYhhkysSLVPU9ikYi
WhdAnElz6aTXej094qalnHeTjLD5VB5uf/M8C+Di0Flmr2WniH6+tvoaVIFWUZWT
XWjyjynhX/j0yioHp6KYV0fjvH/KXKq9a6D3gohzxm/7clZb9odimp0++i1YR7Fp
1ZSXrSX1oBZWq1aCj9Ctt5YQAkFIXRJAUQja7wEFKTi40epc8m3MTmt9BuFNHH6A
4qBeBZ2Rdx5IklBsGSWj603zGIWD4VCfubn27o/INZhTDUvO1K+aYmMdkce54ITf
VlU3RZSIr1IVAj+3rtXSRdB60jjxmZI9OVOKhiRiUp3X7pPDSTXTflYROpv8Uu2z
sktrcUq4j/ZcUcL5pstC76wBUOMgiUMHGtCv/BeD12/thz9/H2BUPcb1G3MmqsMZ
zjNzfjS5sH5pln9QBGXMbSbvseCstF+xxF+qkE9KOdnkFX3ISssm5u/1dkTORBVS
q3JKe7i/dQEPK6FHRHtku7ZtVrP18VhViXgQrHbUIh6+LTNcawZ4jeQfcnShCyYE
/NOyNBApU5CiIajGmuboCq9qWwy0LcoQG9PbvhFe+s7JCrS8mAVWSHlLDMWmeXpD
upD3kxNzMbhIZKwnYZ0CPAKWxzRdGsciRgYCMgJud4jCGxecefEQ+5U2Y2d2nZzX
n43Y4K2YDweV5oNHJt6lZt43S4EHF6I5tBS2wa8XHWXEAyNsZvqEwVzPgtFt9YT3
8kzrxdb+Zy5uXfguhF/V5+q0ma1HxYvkS82IpsunUa3PaASTu0DEUm9hSruFhiGO
EXB1tUTkULzNltBX/UQuClTWghBtPoP89iVl0z2liliRisZndQpz1vqxll8O2BEJ
4sfcYrK4Ldjpe0yhyMqWQIlq3m8PB/fVeFFLJZ6CQ4FAZd7BjgKIifqfH9GJhSrC
WYVYOgMwM7UIEf3gyup+uBtJxVGpMgeVCzt34FOVE/2lrACMZusdBYbyy7uIiHox
UxY4T/grxRvbVNg9XYtYSBvQLzYG54g4V2ynrgXpbqjEXELJxDz3ZS/DwRB7fTWS
meTTyA89EwG1BNomYi+R9vMSP80EDk8AEHl4cr78IF/8qhgqiTUXYBib9MPINGZf
q6jGQjLYNyzFXscJ37kAqXKSvPODOsrGZLOZJqRVuyU0lmXmb9n/IPyTxRPI2okU
1vPwkqCTn91Urzzlre2T3ix3l2+o8xXUj40VGZMiekl8TCs+FsjUjaLsBLY9VM18
A5Bfv0wMm1reVYMS9pGqeuu/HZ4bXk4FDWT53V5Y8G6W3opm1+pY9ZtVoNu28IC1
iS/1qzhc0Crh1nhVqmb87QMlXduVfZgfZN6tVHHNvUnwn1hBBISnNrLtOLcXqpHG
FDCiAi7TaRVzCOxKYhgks30kRrDRWPw3ioglztOxE0FENMnysCZ7yFB0Mp2GWnCX
e+9uM/guxVWN4AoWz74Ufz7aV9lBhI0bGfvMRZGwEgF41Z+iYjmC7x5rNK0nlgg4
lIWn8fF4EuWth6G4JaV1plvrVP3nHOF3zHvvd0g2JxscJE074D01C9Bm2w7y9iHt
2tpwz8KfYN8S5Y6pRFCEBNVmeNzcoE7TTIVH0zT6cHWwyfClfmBCwpcUXZypZWkw
6NhPR4fpi9dhJghbpO92OCOB+LleAd7XycDrCFzHK/gpKf7ZGCL5vX2kp717Za17
iPnw2eE+XrgiwHFbg+VsjMDSA0lo3oPCoLaZqpC0gGb016mIRK7MjRn/aS25KmfT
+xxpCRfCUUjSQTarbuWXZUIns/wY8h8loOeEbc4Ay8RgazK1rCNPdlZ5H9JkphnX
c0cVXM/ZtZ9Y3Sj19/rPTbNP82neZ5KfkEZkkpkU5/WdpId/SZQeiD69/wqqzdg3
i1OGXVSPMpCzEhMoYYbnbRzDGo1bMnQW+CHy6PjD9cf3r9YxIHlxLeG6ml/FJu79
AYXHtd4Ci+tGMiRJRrEvxmNUxq9rh0+zOpilppWI1vvQXpebFi5qMGIQriSOxFSP
//bLHmStykNqvhU6TtWJTn7z6QA3vuxDmQmyZLxTIU+nIwsJEQ/hJQFFhxzo0aEf
93GwLiup4VEIAEQzgJFWNAIee/KZqw8kqzSw6Wgl9Dc/oYRpjZx94Ytq5R+jfCTQ
YbBv64NLpFLwliFkp8wun5jhgcEV1RM9GGRfP44RHGHgHANE8KAWFQtc+i8dzXDr
/stFOF873pOjAW0ZSC193csia37SoJz/j/ZJJwCZWv3uuTEp07DTXdykmbMOCwY9
xbv/X8F0KR14xt0B4++6mI2Z56qYioTULdvTS12loR7iG6yT8Fp9s6dYfdItvUxL
Sfj2LvR4la/JJjd5e8fab05AZK1z+oEaLm+iAeqJrgg/R7osoY98t4NJhm2EvrBT
jlD9PJCuJNwYUE/bm3eKbb6ogJ8uGecsvHp6n2P6VTbrbgw/FS5QXTDATiwpvg1S
iBB+k4heRUB0I1Ks285j9I0/QDdORbqjVfQssH5b/Om8cxa/qiVrEqeIqZGN/6qK
AJ3rE2+0irsw8UvUTz6H+t4mzyCX71ABMet4PTSPRFfdXT5OYkncdYfOPIztdbtt
4aTl8GL6uMqbQGhoNGR7zSlyAxrh0ML1dAb558fljHlQocb4NuuGszhGhS5T66/a
Ay3E9DL+ad6SQNyeau7JGFjEP/k6PqeNLDXQ9mgWjtsJqAKZ95R81Efj/+MDaamO
BQLx0sp2XlxS/9+MacvukhSodABMojhoXqPYzXZt42KQFoip9+XiAqRV5kFAY4nZ
F2J4TsHRxK8B8uvYpFz+EiZ4T3ciKk3ZFAXbHAnFDGCTXqE1WVbGeTR4aWwsOpTQ
oP8YcpqRi69pMTawSJVlskL14ZD0vkuC8Sx/Wh3uiluDuSZb0KhSxXoI+OquwmCN
rKrfXhLj7MAeoyKlqpXHaOMn13aVXhmLc8YAq9qHyA+KvppdCOllqIKopbYF+dEt
K/p9IblFoY7fjTLanbOvOwSAntXZvPTuv0MypOieR+h8uiFopJ8Bq/eisU1Dp7+c
vOQXamYrjTNxvwwzbN28bNgGJkbL+fJrIMPcvSo4xpDa/BBGDbGal7B4HO5RjCRD
eRxRzjC7WNP6l/vJnITfKcjs8TcJBJOx3bdySX7ogdVJl4+4z5//F3D56Yo/DBD7
1D5IMJY0/o2+4ZuT4VM+BAL9pPT33WMwTP6gMSCgXpAIHDG8NzHQ5Je7PO+nBy03
QxbYw722Odv5Q1dFH3xVfhSiCeYST4png4tnb2QI7Q9wXPNFNBuH4aDe9n0POe8f
KHN4Rh/hTHuCXCb7UQg+1JH4OHpE2VQLgF31orNsmW+tlOOGL6jlY1S5GIX+NYrL
K0T+67FimildLLJOdE/fCcrdlSaoLSvq4yupr/ctFgnu/TDjTr8C5mwDd5CZDfW5
cSEr2YIZQ4vujM0SflIgv3ubqYdu0nBFls5ohEYwILt+pETwkc8ZIcVac13pzFp8
QZhRU1mii+SDKxqaLXYpTMcMjwAt4ISwUIu8a6EZgZHKyUZJXDDIhWyQ8f+sCzzm
piE/sAWzVzT8TqhKsZn/jedITqoBGzdhg+FJD+la+IFSGZJoV9hJ+gIG6Vwi/12/
8EgHn28Oy8dUDECqVkdFL1iTZVIy/VJ8n1SpGY/elzcGIqvYp718NlEjkgg2HUeh
UeJRnp5VNidayueuMVHowPSLOVGRZaTGb+A+aWTs5k9eWzeGfbx3z3iuhcAb6oEC
kueM2k5FHdFra0forZN8AGdKQvDbv+4RYf9sCi1EcqxCOds+7M90kje/Aci4Omtg
atWRHcHgj220kpqaM/xRwjnbhnIIKjBwnxOPj/+CpNPHt9vFj/529+PYBWbKsS4k
vFlzPNZfNHKNbGXaM8Aod7UuWXbs5sbUFT2zR6ZzxOsFsUaz30wQxinjL+g7ZLu+
ieuRaJi7e9wkXdT52cNzX1f3Y31w9pLjjnh40HbLYuKF55LiTU09CytM0IrkSVTR
pk9bR7FfNXLBcXia8Q/hoCIduvJp1ram2WqKRts53QfFikmhgV+1QFAuFFQPCZyr
kRIVA8LBbxfRwMe4BdStPNCI9ZKemauTiGQWGMC9oR+jthj61ZQy/WC6SE+JTXou
sXwc7KrUCokknyxM9QNXcerxzqOEgSsu8JDPTwQcLxfIb4bTsxC0C1Bf8h6VDWCH
3jcO0fYPPpz0FDFwl3HKYXtv/YFMoNwhm55wWuL8frVvuKC8dWMIJAyUC6I0waI4
BITBsZ7iqXl8SMN/g3kPLHhWtR+GJRt6srC0j5oXcKIdPJrGdZ/9oc3PKVnze0KA
fnEnShmJo3yoQp0SeOkP6MGT1hLRlPdeETRZPOeUw7h25Z2BMVF/9DBZ6pzYfFzS
3NYAEvg6XeWIU4fhtbK9cHosc0IpbOLDijshtPh35Qgmc8BTu7EJTr/muf/UbGIM
qTyGl+4XjFx9UQWaTY/fCBN1QguHmdzc8Wqaeg58XwOxAPLqdahpmq1iezWqi7sK
SmUd/YpoOVdks2jLPNf5XDAnqIztV3cidF0G+MAzW0wr/ibb5SLHYMRxFmPtraGU
9PBGcEuCjXfQDkB+0beLUDxvM/9mFKo2HY3usDy2Y8l+kP0JZTj1DzE7u68gYh9F
XXmyVPfXWMvzlB9Uli5bmsgoIfrLL5AjsE8Yo/ck0glUhnNIszCLGo+JswJaVkZW
BUzFMTJHUNvcf0FOXzVNibayXeHn1t/Rjg3nLP1riq61azXxmYxrWrCsKlkT6/3W
2+1r9jUmBjjSX6NtKE/Wa9h6H22xea66xgQDRIO60cdAtt+40hBS67qHJ5ZJinVN
hbMzhBt5pi8gLlrdpT66IX7tguMA3UGh9hxiCabDCDSLruIAaGhO18O0Bctpv5wT
I4OIyUGQKGZ5l9sQok4jHue+6ZVHXOlBcG66YZw9bbsMBYMrfSTSR0MQL0ovrkrV
S0jPjFTO8p00ikdOJTQZvFDGagXDNESTanwhnFd9aWM9TO74s4VPzHyjykQob8FL
fhm2vUYretfSSwTMKO0N4d4FLkcxTmxfeYkU4jw6+4NQoiIlCsLDabuh2p9sXHmB
hX9oB4sncel344yvQ3ilrEFiIF9vAov9B+QGm9rgTUYkBBW+IfdHo9N5jby/wnV2
AI2zsOUhZzXWV62ZrhxBpfd9DfjACTebSpvbPXH4GSbJuFgujjQBhMmK+NfZMTTg
xwzS/3hy9wuNIOdJ+gCXwJZwBPyvXNheSb4lAfM0x7R+y7uw/evGZuKikwqSanBe
8rJQn9WG8fyqHr31Gkcji82fw69/nEq/pUGKmEx2dOiatOZ5WXpl5nFzj51UE8EJ
0N1voMGXgH7HgNvUm9rrItGa7rFqOp6J7q+Yiua6q/5u/5yQsZFk/Leor0XPpZ23
6Xmyz0u+XN+zbflEDEgUvtDHY1ehYHIWp8J6Doi6Egl/chFP2Kst7MFJs16LRXOa
3pX4bGOmZ8BvCa39PPdS/+yQ91V1xVoobFMaS8UYBlxoMEijFDSBC+rv5J8IfdtI
8HoahsUJ4Yt3EnQU8K9FnKrLJvyIRfmcJ16lrIaL/B4bdU0iQpa+5eVGgx8Xpptd
Nx+9LK20QUajKMb6B8CA0AXYKNwvK2WgiEdv2vE9YDWrKoq8ICU37t1nRDrVCXnX
Vz3TMSE9zfrhfotw2HlpFmkdEOR7gW+7ZevWaQCVTdJf3ydDhlFc08n/NI/5vTXU
ia1oAEjPJ0lNU4VNaFdV4Uzks5xby1iMkQzQxJowOzgMuTHtFEwneRrJmavlZKjV
K1PS6HAVhaKFxgMZJBlFInaYot+JgOQEqqaGGEO8DVbzolNyg37sg83SzAur+un5
UXbYrszA0a8XdkVkKciZBzoF/HJtSUKh7PCQBmaRDagq//a99j8HGeNS/e7y9k+e
vUVP5H0cKGUBzRebfMtlg54aUUVZBHI+5WWITqHtUPYz9o/oJ6qLewCC8536sjzK
/bvmoeO+taxvig5No3C+CVkS/wUukjaTa7RJnNO5l3i825ulKszLeRecPkGueMO8
/VzTZV+MkphmYknKGMSkMP/RB8Q/OWymqHhU9xTRxpIeWlDfyQBACKrEJqT8fjxA
MNab8HkByadcZoFKMMFXDjVtkCdvAyB/tPu4f1J3bgiigNjooGY/hjVCDPlvsL8x
x9gvSHUH6um10P+2xoVsZ5H6rMDOofI1QWoyBxDfu7w38n6TlswqFHePG2V03RMk
HGivFmv0WH0L9UOlj//q21ADvBEbW+aCjZJgNd1X6ySh3H60CuY381/m52kV4cbb
9Dwp/+NQVwekOXjC+2c1DQr1i3veFmtP7VD9xU+A1wtofO3EKHv1Ccf1BMoPNMNz
4cEAxC7+Kn6e44dL1twMc7BHKfOV1tzShwwwNQkr37z3W5RommiLCd4zy6VPX7h9
Q9lQHKRO7goMtdC0Yfn2P8oppfeksvq1XXjQJ2fevfxpuRZjcERo8PU6Rjcs3MC4
VpZA65o5H2PtNWUCtFn6Xf2PYzfPhok0jmxHPirk3tiCMctwvLOvLtNMDZmzX1PF
LGNk1MUrigQmvLkisvYijwehOKyMlWJv2nAZtOozuLbd4KrO78kWK4fZInThsYZN
VE22c1i3CFgJWBx+CB5ZDULG4jAb2lenKDp/tcvZZGxGRSId286JhGptmVXpssM2
HvD/E9CTIRRMVBN414QQaCGplUsjOfYsHF354ec70U8FnNjXq9g+syWBfDA97AWC
d8WmSD1vc8daq9IrvQrPEnKkR208kShFGJqrMo0GDcMpM8/o9E28aGwUiUPVCMVh
sTE0kudK4VuaYuh1Eoqo4yXzMVdbJqUlPAp7CITyWcn5a5BjJFxBiZIWVcekjSLC
Wc2bw0oRPbIkyk1nXR55rmgM3HRmyyzKd3kFHkxS1o3ksvhlFHcGO6o/ThDFFNrr
vn9FC+w8xFBf9YVlXEzjleccuuY34fTi3aAkeS6RwXevTIkU3cvvqS4QLOZnbylr
e8H2McTOlqjl2+otyV9wwRFyxa8D8SWJA/D5U9dlkA8COCX/gxDlwM3IbvFdz3t8
d0iEiymZpf04Pc7kcsisGvIsukS/OZUd+2TpfIEBOracmmkhXT7M0uh1QXaJOOi6
8Iehy8bXysOiIclMXPTo37fnECsXH15vb9DbKlrPHDSb/WCEjzb3DGuwIFe4za/i
mK11V1jHdU4Ca0BRuZSq2N5dJjscYhYDhIyoOU8XjZVuy0k6ipYNjyIGKXVv9iQs
YvQVzL07LDscTJ5Z/REjJzFL2eM3hVDstQ1Zp0Q7oqgiXjtu7jFy97L6u+TtVAXD
B62v4vCdyLA8wkTLRwosyoejrcGOK5FWlUu7LLc5P0UqPizfFUCoSqqfEuNxvG4i
vloLCC9ebqyvdAIt7wFZyRLU/HNOVkBStX5QQKP8SxRFkVwrPzG7kzVNUhX/+o6s
Jq+xlBLLXCdWwPZDpmJn+8mT1MiS/UKrxvyUrFZOYselZw9gsOnCupSoQFUqVGeN
AFXZdeTxXxH73FA9os1NGTmm+xSEWOko9TQS+2s5LjK6j0aaEaGQWk1AGO5eCz/p
KR7laC/HBOO/v1oNsXF3Brki2uA6q6L7LhNFjYnw5oh8f8NqPVgUjj92LlvK7C9+
LD9/RRRrE8zF1bCkJckzdsp1mE+0ij5sZFiMlvqVSyWZQ05Pj3zN/anbNXCukDBR
TV2I8YN+/svSHTmH81TynS32F4ue4k0adSFoZ9L43xzAI/vNLwZ3wNFLw7QkhFHy
mhHaGHBR8X0nX8GigPl9X6RDfV/xUJQfUAJaleBUOtcoDpIJpOyYcGD3PBbHSA5L
4BLSd0Kd70rldNJlpTNQE71+z5x5JlWA7MmkFV+09w0WqM4SLqsHcLftiOtDIdwL
yZQOVpShBDZ9Zw5IMkDswgyBaWr75cqIX6nvrPPQiNN3LXA+cnwsILc1J7d8msBo
ZN3vX7Twfedin5SjtF8qOkHDc0TAzn7LdNxpo/pzXUt00rAdaIC25os2UXvnOXwA
VFje0AtniFRcARa1d3L0ORV3PhiicZFKtbNsjDDQYDimOGGIn6PbA4mChb2xl86S
+n3B6gwfirQQwGzdjUUEcrEmcHWpzKQ37wFZOwj1N+11RE8mSEBXzydXkuBYBwpP
EVZw+G61F1iz2TjPYfUmgG849Em+U8LU7f6sPKYXxHPkzcFPheA9yRxLMAYNQzRN
xEipN/5hiK/TRpIi5blj7KPHtTM0q1kC4P3E9tYM46pVhlAzYrp+b7zLljsXp1QX
YWmrOsDAVDqyAUNqENkYy3UmKcXxXRyIHXsqobNht9dsYDN7KHzZwTd02JLYeN1o
wwhYfZhjjokpKajTinwAdvC8V2+mg16ERdXf/pc50VavB6IkkwYd2PJLe4YlGcwZ
OmOgJY2MVV0t5DbSKNWRilF5MALraz6NdyaUacLRXWrNKbqsVjGP08O/A0SG0xnc
U6Y6YMCK3K8sAZgtW5Tbh35Yix3x0sl9dPCoJ9W9X4iJJlbrcwntOSZVLCGCD0Fl
IQ1JcEQqDTWDGw2Ee3b7HD85nPxq3CVj/+uhOoHJVFaUGYXfuOgRPKl+itxkzRB3
1e68MfgLU+4jSjwI1DzipdGzy6rO9I5Q2Pq1OEcScWOdXFp6UysB3PQxh+dZ4vv1
k2pVhRiQecvgc/krITqJ4vPiwy5mQeW+xjFru6EisVn0NOEwGKFWhUM5EJ2R+7lU
S7/+HfCfG7jV7vzAn6izj/TEmNR9kbozxvzJUaod+0RqY/TFA/jaNfsKQoiKZoQf
8j6DkSO7fBE4tXZiYyw+aHZrVCU8DjTI6KCvTlksYyxceOzxLeBoKzgIHqqmO/EI
xPKQlJRLvkW8l7Lxq2N4DMNt0FVYtanMI0qICsEZPqRQvSlOsgG47xQeH5CT/gNu
MjoJh6VbLgJmp+wKuu4mat8g8eZn6ajyP2WK+88liNXFW6LOsuVc8vdf+vbOyMfi
uIsaJP9/YMr98CLxXsKbJu2wvRorw+FvvLfaFtPm3Aoe78cjkoHteF/hojsKKQAT
Zq/aat7rzMJzzYmFJOW1o464ExG+tO0IjBqDpgs3pFPAcgScj9M6DeMsdKccXeMG
oQ7GYhD/PnB8xndyG5Vt+ubiwhb7/ufLp6s9LwB+FjXXZp0av53WLFPrBBJMgfe4
uZUoTi6+JCBhDB/gKV5wNUagXVfNM5mUB/oS8hm4qMTrs235L5coxUph5l3J8c5n
yX1jnPAJLpn6LrzwHt/LlPL/naV9WDeSXucyILHFQ4+R0noIztVAnFVerOQ2uUvO
hsJNiotnyMcwTk0UZnbjfPe1qvqQbF8wU6J44g6Q5S4PowQGx98Md0H89LKgnuhx
PMtscLqgYC7qkexSzLH7erfVGUqwVOJGv/hzkIOR3h6C/XzP0B294AugJfRr89FH
f1l1RMdiCA6AT66i1tJ/JL8uOd3iop9NU5rC6bg96U2MQHJdFI561l1KINN4tZ8E
ik7IesXzoFC9Or5YsXJYKx43a3lTDxETgJEWgG8ep3KGx6YGAhl0be2h5FYS0lYi
++uMXdbtK/2nxCqrSfFmUZhRPZcNX/YgdedXzT9UMurbZFtGpPhd85K/Nr4DG+Qe
/IC7/z5GFYBf9y0fgSUVaPLdSC158YqsLWibeUYuBX3LulQvu+1rpNTmcRI4MZzV
6h4ltb9dji8F5ZrfvPBRcJYwN83ENq7j7LoFjD1DIXTRAxzLzK9oLlavTGnPh1YF
j8NCngSVqao7AzsKlVKdw4fILpMmBErlqQF6gHuhwA6sAblUTvg6GeDOauCMz0Jk
cv4ena1l6wXDFfo8sOyM2Kigxq6JZR9lguIz4k2ohwkA2MHXiijONX3enN+Uc0mo
E6lap3I41J9Ka+gr2SC/X31/f8ksN/FGwivEPR0LKQg+tpmNt7YjXTDn6+cvOEZX
NX+Fs9it7DnTDnE54HBzR2mh1OPtT7wQx15NZNxintg9lwwOUP+0MTPC/RoNP1p9
KNDgp9blsdI2+nd6GYQZ2gRxRPxhPJ2hwN5TW5dQV67gOK7+ouh375CWS813nTyW
00dfrBCFHcTmwjRFA/2KyNm2EydyyeYYY6dO4lrOSq8hg1SeSYrTUW3zN4dCWxOB
YpX+ZNF848oOza2DxSrUVMLjyqFMq1C9uCgymxS9RXCsbVKOI4Vx10DcdDpzkV3K
lrLhWqgJA3v9CVyJ5TbPeAlijsfW6oC6Z8Fw0x+lkR9tb1OwhdnSZjGXjnTm0SMd
L63HyX+1LYOkUujb/PUqeCafFWiCy1lS+TctKyjAd1zoPSvitQPI1MCGT72womJ9
33KNVXcV9t41EUZgRKHMEWwlMMuGTQf2wSSmkSIdnxSvCCHXmXJiZ0H96Mf2kGIR
5xcy1vuMxzjU+lw7mAYfV0W5IIpIQlAZMGv0b38PPBrz3+9VLVg3lA2VKaJiWOwD
HPOsuwoUnbVr+1ufu5NDUT5Jp3DR6eTUFXms+ZQefD7bYHr0WAf9q79Mi1cYR25e
nTS1w1m4TY7UWzGGB//k0ePsVNKJpzul5yJC35nX1MnwDuom/7GoYNgT2o6sWRI6
g6mgTa0xknsa0IH+1qKA5Vwn1nO4yZIjEN7opCpMmRT0pZ26OvT2U9GHZhKdcUeN
q81XBb8uag47AoGohQZUd7ECCrS8901J3Qg591JKDxjwi48PwPwke9J7+coHYxRe
bk5iz8ix7d3imBymVRL86FAOTw8CO3+DQCu/gWHSwVNbS6bLc2MxjkGRZtW7p+6y
cJxl6JkZ3d2831A7u/Ay1Sc3uBUfmsh8CenvvU91UkIJfKj3HRKo5bov5JYwjCzK
uX+hxtlfWEKrXq2BpVXdJThJNordngAcU4Ko7EKGHQa39AeKaIBw43Ja2oEgQDBA
1m1fE2mxy6FpoyWI0YfFbmpWx8uFbs5UdLOw8syfY540Vd4wiGWXUxrELVUviKH6
gPvocItJFyV8fk//JRiS+vlw4Gvi+3nIfCgR6riUA3Me496zGEKLh+siZgo9ug7/
EutCasn3tPdUtHr6k4qSCnnSvhF4Obi9UmGvEsdx1kqdKSEU4rWo43R6DLQNwTSn
vYBq9E2n7b+u8insYTZukbwaU9eBGCgSyR38+bcbzyuMpRqPmBJLj9fGZ8IKgsMz
BIFHiR0aZwhGfnmH9/Kgmastorp5dOEVs9TooLk6oagRcLZ4mfmFBR7V0vo31F5E
DcrY89M+R7n0KDVGkm29OQc2nI9c6MvwL8CKd8ZlCqAdUMMlao1Gtksl2aEjPVS7
ayVgl1CuQYoeDtK0kiKJTUt35rkPn04SO/Q1tvxmwJBbixCaK0sVzOKQXORe+cHo
ggYZ5VCNvt1CK4A1r2hYLNHf0Dbsr9xyw6j9GA9Q7MNlf/L7KR9FLWcbcgO78fQn
QyeX04VjkfhqOeeZmdggXsIQ7OO/zFM10Rcy3Ded428iY8YlTjF8ukRpe9ZtSGY7
aCkwcb6XIi2Qa4ZhSb+U7u72R3G/nT8rX5G0cFBhTtvbgyoxw0gGr4LeMQ3xPgls
3uZpec2Wmw4TKxadCS3VV4GDxCJve/57pXeDHhorwv0gixPVh2Nj3b4MVr8PeB28
cznlKChIeBMhH4bOsaPwWjhMzQZcZppLbyiH2YNK4+xweuzynA6AgyAVv9VCP2lW
bkDBjF0hhLiPw9ALHx6vIRIA1qcebaiHKRkL7jykqQ6bZ5J+PlmI9bgzf07KiXLH
3D60ndLBZcgdUIt+HVaBWRF688Veq8Ap/+0l35c/PYZryI4U6+BODSUYu4XAuMWn
DZ1ZZnO26d1vTBG8rp1/N1b2Okp4+UoMcnqWAwkS888KR8X7McCg4HEDjoCGW9B/
Rr0Oi6nJePnuFZn/V/hZtco0yQQyKJ+Xt1zG6UkjDCvbBoPowkQBd6VovwGsZGWs
O0kL5vIeU0Jbbzw8UZDeI2VxLGhEAKjSA+QYuMJgZQWzoRS6S7U6PI/B0Rsf5WZr
tlFRFJ6PAoMUcq1R08lAYpWtsq6060Gz7OM9PjjUPJsd/hfPRp6t79BwSWsVRgbl
34Ko+DhoTVpRrGH4mKA3gvgDWUXkHbxi0AE6oo6sKbM/2x1prEXaJwO9GKl2nTeP
Ox91u4XvtryhJ1rjKeBZiE3Hk/dQ2ZLvVo/KtI+sj+jcx93elqgjsfBRtC8A+B5A
nbCB2vZh0yU1mGDwjDJu6S4M5Rkhy49CwObhyUxMoX7Za7loOZcFT5fkcVheIPCf
JoYbneT3cW+lB4VAvv5/5NESHIFY9c3LpcqaVNGtsio0+C4YvL96xlCw5uh4c2f9
ULHIcxGwSvT0OUurOa0wDdSy8THCWESDS5A/DafdEbBPRHs0zK9IttrS5GXCxIsd
yW0RY+1vtqHuAbu+pazZlDkLMRhd0YberHfaZReyyqkGZC7GX7uAOCWswUsbj3hm
Lwsd6PQha0RQwUERt8ycy9phZ55kZmQZeH2Qi9OYNnfg6me4s2GqumFymA8qdeB3
H+nBDMsMBalxULrO5gHhp7dl5ozoGitfcd6zEUbLnuQseQ+rrUtazphCAkbH+jHJ
aIujGrl7JtrbTHCoK5X39kHQ6NeZioqq/X1qj6QKLHQutFbFn+Z7y+WvAh/FE3Er
N6eguMc6MYCs4GuzPf/l5XviJfAmrNOUlSyZrxTnMZej5Lw5ffOffyH4X5aEEbUr
jPGtyp6lbiCDxjHoX5maNw4WJkDhKAvM7AsT3CzP6PiMUw3MPIYVXek9H8GKMyRU
psFUnrnEeWEtHyniiscr2HCULdTucY+k0VfoiLErDI/NtyfxJrNHv+bPQEj4ggwu
MwsS0YNWDezbsGPy0lMP7umiIQwAb5sdD6b/2YSSFnNPvUvSbxw5uVnCoN0G4ouZ
2Tu2zz4iR3MHUxhhZU9cPeCRFsC8q4wQ00MszPM5as982wtM7Q8SxaPkIHgutskE
zQGee6O6h0UIy8A+uj6eDCpdBVOzkpMJKzc6V9xJt8aRKxnyNlK1jZbjKm4HExo+
OJa4kknzQg+7wv3jjrtWShsV/tm9PJOeDzUd2Je/GQVJ5QaY9XnEOW5f7ECjrX29
tgNJn3ob3aYe2/5Um3Eo09MPQ3hk7uUrDyYYsYc27KAA4nILHiQmJ2EUzZ6zCo2g
BuWZM2gK9/MkhxIBmDrP6rs8+Am7DNPLojyxnimlpc2X+h6UsGmQuosXZt1eUV0C
m/2t85JXSx8ZPB4Oh7DKRlfl1BhUDblYcOarXs1G1AdJh23BReJPPF9vQicbiIGe
PfKBkgbVGRuVhurtHb6DiT2mAesPLf3JoUTu6TAtQasc8fExh8MZPSLNZPrfK5mN
fi7WyL3OeMx5Zzs7Ma/L8qbfvTcqOq9odMcdiJF4CgITnUbiPZS7OnIxjJXyB7Cp
Ywr0pXcwtrLPvyM5m1Lt2gS8OlcC6FmPL8gZOOPowWrAvfetzDSLlzCkkkQoe9ep
DuacUPrjBxU4LU3Jvx02u4A8D+WfQ7xfketYD9xz2FaHl5TupVJ87bVJpyIrBdvA
qkSNeUAN8IXCGnJ8t1ermiWqW8hEJUISJvVLRdipMpLsynl1ovBy1TKPkTLZ41M8
VFlqCj6XprimkOIIFCGsGFeJtpm1N2BUNv1WLnLt256X9CANIeVRsTPlEZykAs+P
cnjCepVPfpcT56Mfnfn/uHYYljRsYraR4Dj9x+ygenW/CriKjgfId+zaILoA4iPF
eOy1yCHYBz1vJPFugdfDzTnEqEoA3LK7Vg3dK59ayfmPH1uji/q67vsXLT1yOUrR
Zo7Al+bBYPLtWtgue4KJvMa9zoG6YGpNjSbBnoc6ay020URwuR96hfiEpALkd9Kt
p+YPfEI9SL11zkudaBkBGTKpf02and4FbRaNavPSAZBWhDbwYHoIA1OII5vBtROQ
um6DdhDX7MKgH11s4oCncL9bTd1F4JS78BNCj1XAuRpGhHZ4iY+lnfRI2A0rWVOe
sdO5Swq1m+GsZqeTPXBevOnqvA5YkKtbm3m9HMDQfxIEiczjK/m0h8LvyfJeurUz
ZkOslSvO6gpVKlDZoml5+a/ZgeM/+SlDCZwjhQcYNuCxKcH/6vbpPa9COdSplXWb
CLquJVNGn8tS69emiejyM0buxS9p2Lyo2SOWwzlJycSV4TwRfm5ksnmhtluYxsVq
rttmbkNULvHJUEsMAtkoe2ZJz6/G0nWyMc9wXq5R0QmgMQGE10z1bw8No2jA++g0
Ocqn5ivwhbYOd8qEaCiu9SVeJ5zZBHDe54PUoQ12AnpUl997rgWNQKd+hCbJ5rod
HbfOuUmAGg/d+rZg21F92PmvrVIzVvbDrteGegA4FsJF3jWLkawhi/NCbudipNin
a9beGUAYXgdJvGbCYevB92X6FWPJErWh/EoWXU+gINhWzP7tBU0tee+rw3qzaR4r
L7AABSd+20exqUULjCl8NdMrsUUsSqNyS4bBN/Crhg0p/9hNlFVtctP/Y+LvxXsY
z0Y+J7G8b9orTcFw/H8aO4yjnJIN/Suabychx5YVjAS587LIJtnOEUOVV9bGgyrF
9f1BUUxKOkbnb42K/ygOY8S9txQ/MDnYEt1RKFFIcOAiQDPROZpd5xy9/T1E/k1E
tVuQIcRGLHdVmjTUJrUrRJHdTyjVGDA6IzgCE9oA3pHiaiqBTh+Pgggz2duzuPK1
assCWDGgdUg3x+la4SDIfs6cXrsCUDc2ObwS/KICS/D6L7ONLGmLPMIZJD2ZFMd3
j5XHjMuNOoxtbs5/LBUWFykFEmHPCAWv/kdUTlOyk3A3+x24EXkqgLpQYvFtC9/X
OKc/8bIvFd6xf4Z6Y43+HhNVZHNQLxk6nVmGMdcp+3AH5tfcL0WunMCRJb0xts3b
6V4nSHpe5GVYEVrIyRLMG3fkTQXh9ZuKP4AT/3tN5BltTks2ibq+dYpndUR0GPdm
jNc24JicBmaQJtcvDwcjJ4QCwI4hQzTgsEbJDFAGd1afEI039inxadbcLHPdT9mE
9B6Y3dn9Cekn2yzCD5F2K3ZoOZbiPt4RMOJ478O5tW5F/GnkfQA6y22BZtHYMNRU
j67azp2XD5ENGdt2lrh8HFLZyNwNFW3iKn4s0T+bvZeSZIFX2bVcZqj5yszneAPK
3/3dXuRJVlCmx+lrOR16BxlJXH4n5Qvu+VQYyJ+1RlmXYcZKIaqV9g+8M8+hK/9v
ODfhyIsIENz+e/20d5uDE33ffzHYCeKrZmTJjtColKC6S3lUZJSHYZMJ/RVu9yC9
Z8LsCrQ6JNUHG2XdEhfaEOJ/6YDZUD1Py8f7J+DxIsst2WCGEpKO6hJJFN5Taf+H
tr1Pvn0XUZB7ZhC5nmRUaQdBqxO3zdpmC2aXg8ZEt0fl8GhkBF3qmSBKruzov6lX
Zy24Abx10aHUtGLGB2pZ9oWNAfJKGxUpaKfq7yPf0DN1Vzo0rexM3Ep8W30y5CJS
wqSsAiOs3RyXsNt8GZnxCdhcDDw5jV5eEYNdTlArta8ZBoFQD6nxy+Kg0qVLmx8j
cJmscAphIi75/3pwKzeKxWJMML3RYGNy5gGjShmtX0fWj42JnWn6Xaq4M+T4PkFr
yatyHT4k4t1pP/Fcoe9CEkINQCRApLdx2i/prC8QTPTITAMDIQP1aDiT1+wBL48V
8PNRwrdDo+dVJAKYJPuif2HWlVbbiZA2n/VUt8oaLj5r95kFT/rteEMr9CwqUVVT
+5pBoVXE4WcMwMOyCRVz0LPobDkyskTIMNbaV0mAUgPH7i/XVlt7IFzxGrKRCv0w
DQN5vS73Ojz8LRNpy67M2IVIskNKoloJCXFdsrSsS4aKl8vfBQGxnRA8PusM/w1A
87/hORS2GyTJXjntZLPmSJYVRky1PB3bC9bVOHyrzaqTl/CIDVNk0n4LJefxoqv/
eTkUvL0GSegqLWp/mS7mFn4FfcmLqLjC9ANSnnviYr1G64zjn94i6MBCBc9PBS+F
tFn6Lpyzs/PAVTPNJB++aYzch98iM37ZOjewVJQGjk/F1lkAyXG2XJDAcv0TcdMA
4zhlC6tc1nKV6ao0sdnmorvsMd8B24/O+4DwcjRFjyQ/5YJclT03YKo/S4ei6OBF
Z+15DorPfFA9k0pAXuL01fpJEVRJzMfVdbAti/z5MZwqChxy6LnFK06SgAA+/QWf
B1gOy/zqFoniSSJM1hkOt+ACBW+H1dii47PsGXMmBctpC49z6Y62SUXeDh5Im2xE
GyM3qTXhkqUUVr4Jl6lHtg0y+8miZE9zB+DQXlSZ+kT5wnYrpdCphw8rJXgvDTth
gYtSgrpgVOXuepSsCC45iXS5cGc8WF83jj4RvWzawqhq3IMyBleeTX3aaNmKICe4
r85rJd9IFHBy+RRF+BeH3enHCxC3t2cLqKx5KOB7BhXVnGtvZfXVD/7dfajUAPze
flxcrq9OPg8O5b1Jq92ahg97RPxPKAX8BVwUBXnnlnhLDiSDdeFrPGY1DK6iGnJd
meJQR3JVGDsXB2mf58CMNYUuMXhY/UETfwpEzFUqFpsk64AJGjS11IX17rfKA7Rj
7d/OnvtYnaIuL2qheYOUvicoM9wrhjjnI+qL2wWhb3U9b9qvmHQzhW8RE0HzDJ+U
8qzoLptDM/1a5JWR+5fhSrV1KHBqWRNYlhp8aXl1AiwEZxBKkq8CqJUd5Jat9qrv
Br9JmygJ7/+tSmunOwOdooHZFthXmtWMwIpo/eJGOM/lkQVvAomzz48kiBvtC6YY
DRJYH/ObaiGTirQKA2SNofecLipUcrnp7fj2I5nDXGToRAb3P71bN0Ns1xvcVSgY
MSgglGelxWnuPq+po074vpxU9quHvNB43bACK56Zv8bBPAm9PAe3e8jTMdFESUJc
9o1Gzr2FzeGpHMa6WSK1veCZvbVrzEFV9ao7Y+dXP6yHiXAqmtCbZhsxPlJqSyvA
0w9e2vsTs/FLLztXzft2bTotK5fRgqVlQwecd5dQfd50x53vVLXhOwUPgHnTjfT6
bEQcxcQZHMvrRzsQXDOYfaU0V23cUxNbRmSJa/NfGkAtqsZkRV0XiXwBv6Z9NQ3S
/AqbA8ixQ0+agjsTT8yEaUY3sxgMfqI2nm2wfxtXGlPhLS7wcYWYaiHSsrpx/xHa
5/tlPnAUwzGaIpDiSg1bNL7PreJk3PWP0+Z8VmrH0vzfCzfh33IprK/jxoxI+9Ga
2kQIsiG3Vw1m+ZiVMYfGTC2tILSYZhNBUejZZfK4fCFPGwKEw9XyhHqX5W0tjNA5
V/XrRve2H5sVcBoIGJqMexjIRej3IELTmYssniJ34YHUIBV5Zbr2TA5nm5Vskjtz
+Bn6+tZ29NPd+fI6Lax/g0d0wX9gGL2AQFD9bk4CmQeDnF2PsvmbRM/LdwnjomdP
G8HAIRW3c8Pz5Zq1WTp2IldsxuT/PpwqeA9UYYGeOJ8sl30FlvWvNkJgt2/rJ4i4
t5Al5w5iJAN1R80utEI3ejGuzzIb5ZWgoQbvfVODmPrd0kv/fdDqJhf3FzdF7AxC
RgE60t0MelfJa21HSmOqynGwR9uKa1FmzbP59LQa3U8rDPvAKqkgUyTeWbd7mDvh
AqqkCGuXdOLIti3JzAc+Gu/6Qsi8rkpH7ju7ynRdVjqH/Lm78hrFaOWatMj/xzVW
Cx40/7451mb9swI8d/qaDyraaP8UEImENYoFmO0covXnt4hmOTXlfzngcXSz8qtk
aY5c4ZN32124aYQq0R4zQrNTFroCEujTrIbpNJK3dxCLhIl40dn5umkHdq1QQP06
6MVyVTTpS1oafQ7SurodqQQLGZtHtEv8IuPPlbOUdVd7lpqdUO0qVrdNVsoMHoWH
Blm94dEckBFIsXaf6YHx6YTwgKJGBIHpUdrOLV6X9ViSv4Qfy/4iJCYWBFGkCtdc
6IXoZaMgCgMgcEWGmPPp/eSeM6Vi5clhVJK4FcaB5qAblEsxSKnvOGevQ6bdehfd
pEP8YEAZzUufalmmoavd8Ok8klaSnvJVEl0h/b4rzyoow2fQWXLsSQB2TqmN8uul
zO7gQQgZpM+4JgFzy/QHWfV1zkWDiWnKF0VhjL4SBVYoLHQCYE9ISaGU235eUhx7
takOpmIYfRhDR6viIvCY2mtTzZ8WtniL+cj7ufaVpoUvLTVH/E7Tpd0O+2676HUs
10LELb0WlmXIGCE9gtDcrKPcDwSpSsreiHeSoMI/5gyPucN/nj9ijL7g11GzI4IN
0oNZqeQxi2JuSClIHFi8u9FOTvfP4hB4Q3xfdit2uUTt1c8KVTUFY1ahWX+N+uPT
9viBgQAHUD3RTlyMObQEljKaHxHpqrYU9ALGjAlak6EAW30WTjdVe6W3lx3ljz00
U60zmhWxMhhgvPEatmIaQ+RaainEaSdfN+9rcUE73VN2C6aDgte2/eMQ4EZKOSHk
nqdjVJC20KFWT27Dwlh/lEiDmETu/HwztQLkNgWUu7FjMSIZs0tT2zRb/HTa9uFa
+J1pl8WCMJIALovVl5fYC3ssK86jMVgLoPFIDzbucnmK9wz4TmxdvW+iQpPiPVt0
rv4hT3SjKamEX6qIZ8iii/m7R/rocbg+P4ijZdE4KhfXHVDfVqzy2lsLDzcV/Hm9
TXRBJX4xk14rjT4dcsnClkzk4kBEwd8eBGAonmRaP/9KPzLa3A5MexNV6q0svrF9
ACIA63fwBKkRRvmF4RwkKwypxes+2T3hWkdq8XTxIN+f/G8VUEimeAC1bC8fNL1O
Chnju+t9bUb8eDwjkSuAefuvL04xsRLxVUviy7zNvUhAnaUZJGAFItt77DOpfoKJ
JXpCPeYrPAN4i8eVN3xoh/I7OTcw96oLkky870h0HnpjwF4/nFc+k605YGIkHyGO
pCkOQDvx6wQxlPluR2TMP4bKslcGXzEzSrb3+zHg7VzQDhEaluCHPs55FhlCKNcM
D3eLh2q4PUyeQOOUxvsRlocN4W/uD6fYZQTNuV9sxRcOppCk4wbYzlis8liwRt02
FtVnZZNbvr1BZapMFekFhiusZ+L8tKs6teJLvg8VhmnoOm8Jj2LeDA09UJNoJ3BZ
MOqoPMAD1vUWUsVJmAx1uI+NswYfZW4CS1RYPLNKUdwsTcGDMZ0lSe1YbjrgHQv3
WSAa5PB/qgMCti6pHkHOFwWA0l0iOxMPpByL2tjrvPalzaKaaqCFU5sSpNKibV+l
yxOmblDKg66wmPzcje6avif0kEd0aVeLj/fy3v8UbRGn8xPPO7ZoB+TSCmyOAqhf
UQ9EnAWe+PVivtThNvs4HAFtQfjxBm2IIutXbSd85x5+kRY7o/VJZrVCu4GNrnS+
UL3+HMT1QK8d9WyGWik8gklxcTZR9txnLGN9ZqbUIiMhO6LZTLaR4AMO3E6Ix5bv
CtIU79KdHVXYruyyu68SkTMdSkygjVKIFKJrPK42bKLo9zeCwVWjFr+aezSJKDEi
Wy0xx79XhaZtBzq8wekQfl/TkObteqDHVdRd5Pw5YgybxP44OeAu8EXVi+APfsH/
G3XEy1Mt4pcaevyDGRa726ThNiH/HWm7k0IB29tXYXsVIU3oAkm51z0WHc5gBtdh
ecONpigPb75FmFfSkwS+jxYy6zRKC6RjT+7mLK7UMw8yQJbpN0eeF9CJTXY7vrMo
OsW/C+/U1KKMCx0kwJfNiPJv3Uzkgp47l9tBFImRRMjOZrYBi1F40czcGWO5SYME
3H12l8TIellZJkXPTAqckcG2lGbjyGR+oxO5iv/JJqNvxwmY7SygkouFR2mb2Pfe
5sBzzGXH8vO3WBrdssKpBWEWvxQwkhwXfCq2wFLFmOb9eZCHEN711w2ug8Mn1DLd
m9L8qvCg7n+GkrxDZq+ST2CbpiGXUZmMqU5w4YAV+zs7tVXacmDSuF6tIauOgM+7
7/WdS4kxwoZTdIzAuFlXAvbLgo2zgO4eZanKnsAQ8EIJ9TDv4aM6PhDE7OtsLuo+
KY5DbDpprYYDOdSVBH/Xeh9xT78N4jPKjqJNo99u2OIPyC0VMoQscLvNFYY4hosU
AjjfEV045OwQj31axeOstMUFAHcIggGfWSe40b+ZWvT+THO+SdgikrwC+shEx/iN
9sXfnM2YLXW442WrOvoySqHJkJQKzDloBH1tDcojIBJlihUZKtDi0Xez0/8343rh
XJW6HJyFMpGusLMFYZHJ3kENEJhCxaWqfTRb6CzGUEO+tuISFV74C3lgylcgkDKZ
W3qm3dJ00rvzFYMLCWwUQoyv7/kX+xQJcjPb0rytap6NYobpoXGnI57dJE7d/5E2
MpAjM8cH82LfvvaYJqtVJKtQJr7MOrJcP9xBrQAmsMPDkozCpwzgUDzu0LCFueQC
PPPeGb9O8VmvBB5Q2X863+tUjtXrL6mNdT7nhiRSH0RUOTb0l5X9OEJp0Dh6HzKA
OjFXlftz7SvfWV6FTu3qKZwvKC+1KSdDeMf9FJLeIWoyjQdMXGBI+faA2a8E4+09
1EDAJxZ33LEGsQI1KQnGWUCv6qbBzqZgUPkAxrk3djJOwsps7sMEbMDvWHFWKxsm
Q+WkEMX4wIVmYrDb5UQ4A/2V0TcPowesuCvDu6R1J4ABd6hwg7dUveNO7D5ZJxJx
rQPYjn8kDNgtz9AWwhJnoa7gUNo3/s7PAFipIB5HA0hlzDLOfmZxnFT0w9bIB7Pi
FSoYdORNAc12RMc6kmVuAFPV89kQ7zT0KQsNjUPlQHH3KoKo9inDu1U788BYcniW
zISzM+bQv6LW++HdL+VjZ6su85ByOJbOA9gVxWp/R2D5T3EWP3D/93F/Z5z7J5X6
KGmZ+5SiFdx+6TBzLs8fBIU8R/S4uCP6Vl+QrS40xO32o8BW4Gc6sSonuErngOeJ
u2mUHRDZMBZ/iW8gxLI47YSJEhvg7W9cQ1px5hPLaJqn/dU6Inm8HuxwHhc6Do3r
RW8oXtYQ8/E0dC4dhPtVuD1VeavGE21/AXBxsH2tPkAuTVJ00ygKyu0EqAF7XnxQ
c6ps5RyCTauH0WJyBPM9DmGAGy4acb2ED+1VKQkxC7WkGVcT/jYDphKH7VspJ3T4
fZ9YvTXQAmro9wCQ+sOd+ANhWDXa+0+oc66T9oBFmzHhAD9Qn+UXUZzK7qil3MKq
dVwvXxgIX3M5eJj2H58FXz+sXY493uuJxL0hKPvXPczrCdBW2rOgEXCp29Bpv09h
qJyxgA8h364BVUZDRKobNSqKkYqqJGwtkOMwkPKB45C/fdKaohVCPSQbyB1MMKHw
b5a+Lz3986SuBMePUDDhov/p9jOP0npbYKw/Ptj7wr/dQyu2ujjIhUjGrJdMNlWW
85zNYUhnAnK0PgaO+zlOO18AvqX80yRGemTFUIegjt0PlAEc+2BNS2JF2W/cgBXS
ogEw0BaUw+ZkymLvvOj/qLdSPQoxALsuZZXSLZqmX01sn85SCZVfi85K4R4ykWxE
wXIu0griw6CZmoR27PcZsOi2NU+Mgjw5FqW/VjGvWAmAUpJG4rduVKMTYrPcFoFF
zDTtbhZM8iN5y6gyZuC6LZ9rGgMOUgVoqRu+N88FuxdZZkqJtT7qvTIYwwKt8pYm
cdv9tFYFHHyHony7SQVtdpjVcOM9pWArsa+DOLErqYUlmh4amQ2L9rt3gnqaeh2g
+9XvlOgKpCXfXBYCKl51ZVZLkpxXmH92uqcgwhz9LZRNmLWuPRmdS6jHdRo+7OP6
//MTI/5Ac7WFP1S4zkuiZNvC+HHzYZ/XTbfAY6ReaSLOC71EfClrAOVoQmHOs6XV
121Sgfr1B/Gt2u9TJGs0Djtskjl/L5OMRgH9Cj0P1muRH9hVkk83OUw3ThTaWroq
aHzVJe8V+ICVZcLwR61PVqufhUHyAjNyabbyCmA3aPi45ch015PxzG4OZw5t0o0z
ZpuqD6EqqqOhFzyoqmMF14NpwveyZT++4oqZlSx0Dm2F3FXeZ9UZZcphfXuHL48o
s8RjUittF+1ThUhV1eUwavSjHPch9/eujZP6JuJCfWKVsDaC6pqI/55EGboAyswQ
wv3FGql2Sp2/RTOuRe2KV3PHXYiU1iurXTx/L2lSogqrxoNqL3zZekKMznE+ttQx
h+wrbgPHxIywO7nFM9wv3lZ8Ln2tf22kyGK0RjT4olgPYmBv6iZbtwCRXoZXaF76
whHehcpKSr977pR/zlbvrgIXCQbgiHlkErXYP7PKqmXTRiCMDsBHtZK/lv99ytbx
9PqMQTVWP/4gc2OgTQytYOBcQYZBZl9lfL2VZ7asCJN9RMKtodWb1t90sTFOM1Co
C643pslTTdIKFBc+JISv8jFd/mvYB/twwuz1pBUSkWpwp7lbSUBi9Oqt2bCPCvVb
2aC2tr5HskH50EvKALu4C1uVrxFIDGVE9PupeNf9S6ZBBhbH2G25VYRt/7PIheiQ
HyL2NFBEpLm6x6iQOBJ4LSexNq9t9J1JnENlAsZ66hOtiFiVcb9CCFJWa1XRo02q
p6aTkxj25IsHpSxviikRVKHGtkqx7YHHU6r6Tx4tLlQ4dXNHfJZeBD13SnVmjGl0
Lc/PLQC/J7ygCJfn/ACg/sVY0MG1ecC5v3kLl9yBIEFldJoXTNwnV929v91KbRA6
Dz32N/5QLYze+kHEL+ismyR2sBQYhnW8pZmWMYB/zNX+6lp4pymY00/CNaDlPDYu
guJVtBpRHIcAwqODE5gRxpxS35EqHvzD8TY7HLILGEd3mfC83kyAGQbEHIswcjmt
8/8QSfO1QsBR5EmfYs9EzTLuajDQrIi3yZnJKnrEW8ti8vwGJqjlpWaWsK9jIB+M
IpyqImMox36zIx6GrPmCOlHKbb58iG+mirlTOsAmsQTqSfXq5EeTp+/DFjsyiUCp
9gXv5JrJomd+XWeDwq9+up0bLPoIm2cwYJ8CzFKtcz62lJ3SSynaoi1NSU9Egy8X
A5pH7pJkoJxrPt68JTxlpqEPqn1dgSdRQSOyIfNH1vr9h8AbnjLVuiEkfKV0YBcR
+EwoV1+4oPEaHJQJ5vPLWyFy15IAqfYt9ozj7s5aUKXy3YNaZxotTgB79CEMmHjf
+09xHl6S8bQga69m69pZwlp7x7eWhtgdOuOsDAK6a/f0KoiPkPcXK0eGMr8UKKwH
gKWtGHScVB71Yd6EiXqm9Ho6tkwCVmdruLD2MdqnSf2PgkBOntpKifJHlIwdiA43
6FVVACagUCfWyhecwKhbs1KCoguE+g7c3+zyN8V4ISQOkzaQTiJLrnW1TlzjVkDq
crQRIQqVivZxEBa9xdqZU1P6FhLrE/BVkLqxGXXDxs96Tho5t+0aNCpJ6ORkzjDG
qeBBcyIfrraQXINikWvUEfqsbbKnEP4+TADOG5tglr50EJp7afOWDsYj1FV+Jdmw
IGOwO6B7EEymQ3jm4ZeFxj7QFVDMGMZ+lKa9t8LisuFX52QOktr4YERPyxqyK7ZD
Z8CO6nRFvt0Xkz6QxM9gOiDeJFua8GGMH1nwwNmDhIe7JNIrAE7O0HMnwyegAXn2
j/LPlWFzU1zK83Kcdeoy8IxEXaXRUej/kzGs8WKIM+ZeHstDRBEcnCPwkb/pWW/r
nvCC1nR6T3Uz3IzEfuXfi2Taa4rkhydMz4bPpiGBfwfZZfYXyWLJOt7txHWRm98Y
w3+gwSLEfT07VtwrMAikuDazqv3XT843pImjqdRdB9qhAp72eqlSvUTvdcx6xSVL
nIWH7gU5ASClmzT1RExSh2TsesxlB37xMkzgrNa8p3QmxHx05zYYSh6GcigLHobJ
sqnLeFvx00EOCm7HCZCx6I8JMrfn9n5yQi9SwVOFfaoCIVO9lqZdDgSMMpFdRVUR
n+O7/oIYPJ5ADYxTFRhPtQtsCpRpd/peMsVdV0DHoYnxMosQpOjbk/74GSD0BzqQ
7yDmvTQ8Xup3Co+Tw37DT9j3QlP8sedwrnTbqPWLDGrOF+QT5aGgH9cq8A1tkKqH
0gKRlX6w4whQgofIwzLY6bWO3gKukTuweuPu6K0oIZ0/9uGLfBb1DZKimBwz7nPy
4milXbaSwnHLiLx7BPt/ZH/VrYSQaMvzInSMHY+D4Ny21NC8JyglEvzOeKntQw2P
p5iYB/t/P5X42aQVOUY+/MTfgS1NS04sST2m1R8Jquuno34n7yAQIO68lsDBDTR2
UU2CPTAa+F2iLrzGaUQPr3+lkn4Lgafdic4bKQar5avBSDVw/MnfO1pmcHp1NnPW
YD54NLzPqmBkq9EN0+1GsdVxuqb9patA+fYEJlwslLWaidRB5r7iVBJBeFe9inHj
cLPbModHs/p/jjhj60FT21c39tvUUZ3iy18d4l/Fn67FF6rjNDlfkepR3QpTsjya
06mibQ7MoGKQyXcqPipNHokh0qf4SmJF6LcbKKQZOsKeoOZgn64U0hCy70jvnAM9
GBm2wMGb7lSirVpbJZfOuA3Z12JE3iMThnnvXknbIcb1CQ/GuogR8DF/TYuL+qhH
gun8bd+U8pmiUSmgpsB1zZwi+KDLqn6aOj9gtaQgPxXz/yUAtB4sAStwF/Ur5hMc
YV4auIuiFRMw28HKSAWrAQ3jMM5fADwis5ruI9BMXalrFjxVCiVWXoizBPuPxL9l
Hhw42FGYfcr3mknq/etv/IaKzij1YqbsWc+OtBMTRM87vqD6wKJhOP8gjpHKtrIu
YyzkQ0tOTdTxrUSRA3RwVXBBKCzC31pYYRDrdtsvgBHx2lVVozFZdh1qscOoHisQ
F8nvMIHtzfQWsWjYt9dzg1vhuJHg4Da48lVYWWdDrJFI/C7AiAI0fhiu6d0RRt2A
5y3Z73Ly4aUefCFO6KJeXZ+fqa5ZhSmWhm6oYnilmIeaVh5tcFh9CMbrMF47qQu6
CMoBRZvn/aMLj1a6DqQsXgQqVXfS++TXei/HZwzed0aNiGgyzMSOqM9/k74hmOSO
KpHoseVMLEAsLOBu6Jlwy5Bi2w5RKJrxHjfERKDjJ839AervoibXdhv2Ggs+UWNo
6X4BkB7x+5nqV5evgGvad/H24mUs1x/J6kqeFc+mbQMw3NnZVj+q+e3eh3hSJuP9
ZcQXlMMlpeHcpGmRvTSlDjjQUBpxMz8sDcx9b644pdZVsby+9Vzt1XkAX+kSrY8e
DqH3/UQVSX/nSCClASLmSNbAd/hMCFM70wd/OWw7Mue/WlRGIVdQkq8DuLEAipv2
1MTjcSlvHT4wNCHfGGJv62UnT8Br/+aZy6tgxbvcWzqjN19JJUyurtlcEIWwCfTV
0vy2a0di/qMgD3Xd3OzTh+uXNh6Rkbjgc5HxOXg4zp6Kjkn9oBlnF0wAkmuxzkuH
5C0sqGmsxHpyRqa0JllNejVzJmuG0H5pVRWTj6r8gAlXeC1fp5t1rQEuXS1xRg8Z
wThUj0rjWnQ3SZyzplH8O7+kJh9cUdhNJEOSO7VK+iPO69ea+l1CwicVHIqZaOHx
qlb3/psPOjq+ydyTorQ3NtgfRVeG4tCC0oGi2nq+4yTykTAAhMd+7CQxGsjFJ6VN
cUf8gCk7pWgaG75K4GhmUcPc9novetB67isUtGyxxfuVwfdKt6lchaKtXyU8XaRv
w9G+9aMc/McIUiiazIRwXjmMnTC9Bpd6eNmW8AI6MP/wB9Qqyr0xwJNkotk0tt3H
d7NcK/NoV1/+tXLAGkjkHJFhZOcw2TizvWZUpyK7OE9pzccjLlZqC7dJNf0rGucz
osiPtcdt8fP/yI76UJyeAX+CF6YASHV3ZQIHujEPqQkZ7PEj/T7B6uxOl1UbfZsM
JqcRA/VMlE9fuMWrn2lHhkiIMc99m875YjSKM8gHt2OQhWGmGQsQKV2AWxrHn7ia
yFRs5rSSPslvKgZi/qKNzXNUsTRzR/4r5iPZOfUqGHR5rdZkLTptusm8BijdIoxi
QahPsDVEhpV2tWKhoOtZNbTOqqIYttS+sZDvOvc7ScOQ5jTZvIyqdqBkUqNlwbl0
t7XICyg3/+cfrfdPZA1huC74SfMGIb5sCswXPC6BNpUcjlsWjdI1jstHLshCOZX7
QYcL8+wPD0cK72BFUTNcYknJ4xBbnmrYXp321euE0sHDGljGqORZezAFDXE0Hy5L
C8q8bGii0evGZQ06Fotwoz/4Bqdc1jFNAREFo80wWbYkWBtCo+ch8bI40YnfyG0i
IV9MyIMzXmnTtrW4SXzPozTInBdd2aIm0mpjxRVkjA86K/WEnp7eJJGWuiAEO9yk
alxqlbnsIgGK2puOlA7MAYbq9DpMIZtEzeUGHuVEGfPNSLZHjjWCeGaizgflon1h
w5uJO+r02EubzBTE38oQsQd+cQiWaAV2ddVdm3z8ak+vdE8j+gkQbpolOCIb+dbL
MPOnHcZNusXKuJ8ALffcAH5j9LwTwCKPwQp8TJw2FtLGts9uu+aAswJwQi5YBcQa
QWokp3t1N6lfdDRqOVaMCYTUlI9IOv3AgzyUZIDr9i9iYuQXA+n3S1rGQmv1oxiw
Csw4pcf6dlvX8EjixmJmRuLZHo58z0wpUfA12iFnSQgY5aBh4t9WZIC6K7D470wY
UMAF21imGtiYine/eCqaa7KioJsYHwCZv1JlhyRGy0FC0WHEW0+0hIZIvG6tgtYu
F2vUv5+IJSr1CBratY9O/0ALZa8qeUjQn02KskQyj0Rhu+iAh+SP1juscU9zIMHB
u3bZdMRwzyYNJx0i69fFyF182FhJTAdo4eC3uJOluxSrSF9nnAxyecbFnOhhChdQ
VQFSo16yxomOxOymP7pU0JWsLKd5C2hMMUZdX/nYalwrtmi19yYz8Ns7+tBclIKK
Y7bLWW+BMkbR4CPcIai4Uv3hF1vuCG7D1ewDLsMN25QWGWOnIQuaDczED2JKYHWn
N0eerreB2I446Rz63BCxbTvU890uWTJX6Kqfwz8FzLMaMLLxZXvcE1T6Dzhb+GhR
h5ZcYbNd/WrCTwo9BNPnoZnweEQkA7m7k/jgRIrIv31KUt52iLYu8BSulUDaYCtH
VDHAWxrpwaos8e7a3EV4rAjpFyZUgEbL/lt6HaTH7kguJRg8ASsPuVNdeRyUXZlj
EkPaL94tFwKLpTsliY/DUFeQDhxA83ITeth7oR2loyiYUSoPO2z3Y53yq0XCQA15
+s38ImEV6c/7gQtFFg4hfE1yiTwkLwmieS4/xggD+KDzwpF5a/CkhjMmVKXQSD9o
ck+Rrp40+GnkBDKpXeMRMYzyCg+c2+Ltif0aN8QimtNPcpvuYNcwRvHlt/FdYV0g
CCOwrC24HKnadff8iiWExW9BkhHw084eusQTwdtJyhPmCs5ABAx5UOJyc/f2TZBB
qsD46W5zkCdRow1UUKJTPjzCKjKwOtA4fEmDwv1vhkFw6xR24u2wVvlGfZWRc5XR
j8wOR6lIsJnOAf/uHFTGy4La0JY0vmUcGarMJ72ZFjLL/C6pGH2epYRgeEncpzA5
EzjyIH0t9GVOfS65P29gaRrXCTCAJMqcqNM5j+rqURQUhOdDGiUfjWXeY3krYL7y
K/Nub09/zKc9zzoukUsYuIjvYVkREeOiD61PieUkiUstLZoQ2wy5fif4/cD8zzQu
OChxa5Z+nzpl6syvcOnuKI33GkCf8r/GWJ2UFK4esd5PY/4QbsCFMG/bNv+aMYbi
Dk9LyZQcCbqJBqHHygQtmkuO+5/JYohYnElTUbxNzmtbDQg8OikbmeZ0HLM9cPtc
iHpGkxcq1AK1Afoan0YP2VKfh1Bl/yHBulRBmaA2P+4Xj43CFCTVTq1ZgWCQeOyH
VhMqlzxRKMVzg1txy2MpuGW0mSVuqhjlAZME3PlYTIdfrErXvZO41vaGUuIU5i5H
SWdJe9qe1gE803YcET4URS/W2BubuSwebjmKItXJiNKyFkUg/VK70u0wVJYTrxLo
Unvvz9xcUV0/n+7y03b0tMJCAVHnhZsQlilp5zXwbJiIkCpBOQyM1DpZkkCztxk2
5tMdWmzKPaumJ/RjX+/njyer8B1ITrK7YZF6HYdw9I5Zb7PNDCTZ2X4iONhpp5Bt
iOLiRWftGj0jFHHUar93ku2dQ8e3c96easqpx+WPFu0zKG5JxTpe3x2tSXndrWup
H4N54YMQkvxg3H4adLFpSLPiCnz8dyK/cvFIRojBDG1B+6wAwLnx+txhYOKFEP7O
o/akbMUTCVq0BbBSE7SHAU+xkG85/kyiP429wDyc+ngE7PajFQmO1HX4xjAG3jSL
v5uyge42JvFlYAelM36IurVAoTW4Mb3r174kNcXqKV+8sw0WflSzs4iLW7PmDJzj
g3AojOi9CI+nSPb7Xu6GlWUvc1iOZJ2U/nyOOdV1mNQVx9CM8j2HFX8pCnF5wAt5
ETmJ6GFSQRumKxbuT7MLI/GDz9EKCC4KzVzKDTi4rVMSsRRfeLUinMNHxsH3Ci7S
h7isAuI0ldWAFmXp/LYjJEhEb0M/ygmxuBOI1+6iiEpxG7VHQH2WDUFZ5NzO4QNl
puh0duwPMqaf73K7Z2nrldi6ev4ABEHf2QH3fqvDOn34dO7WAhLLt5QfNKJARg3x
btkMLQaTkVKT978JJSVi7/36cCjam5KO2S9nXbF52KDx4YBgWE8XN4IlDUFLfr0m
DEQ6hn7j9q7RGAslMJqSpDTRknRO6iQVFU5UT5AMgDR7dDTVP98JTuLwOK5DYfhm
7PfJ5pO1xWjZJjnuHkkZJnGOseC54aIsN0i2PJhBidDa1cJ+aXbSy7NhIViZCUmj
XdjFKINO7gWAJlXFCeZcBNUKlSl+Tt3etruaXFr6JayhUCKr9GwFQ1DgRWixEASQ
5DIoRlJiAJaAdSXAiQuUscFiblYHx+BDt2OuvHxALYRhq+uD+QUG0jfX/oHhijMM
a7cdYlIuDN54nWmsUPCfkZrfrO0R8hWiWuVboSwpvHQXGmjL1eyQekB4LAhHNkpe
ZsQri8GXa4/S1DdEKHuOCR38InMQPyZxdg0GHPXmZPj+Lx87OzY5VXPVvxX0Qc7P
A1jIxavSGbqJPp2wfajd7XRCEGU5/CWAWK6Rvta+UEpIltqy8awUelSU3PFUM0fV
H6CeL9oly1e6MoYHcZ/sBDSDlCI40WDrQFklJV/bI6qSXYCcO/o5qgGHGjM2xsPj
QmXchI+LpG/ZMINHvdDScDhe2JWcKmJPejwJSzWKUC05TPWPY2jUIRGWaILz7Frj
jt4RMPffhS0TazeUSDi9B8QbLW+uDcBpOPqVqo1Xk+sK5F/pD+V93jb4wAKldT+U
NZtrgs6qSZw0H2M83CoaaTGd6WpBX1nHnHXCYEA/IKq3vLRkYOuNovroZtKPzmHh
SOIjFVFc6Z3Fza3SgOxQMCinOEOqTed+EK4qN3IE1/VPqyW2vTE7mw7T7EZVAMnU
Q7V2lVLpbO70xCe68ap3FwlPRZLbbyxZCGT6PbGlXGSz+ZYILH48MrvA7fvm0uku
lP9rG0hv8R8VygGcl00sTDdcdT1dY8LTCvBhuDsIbElA93ba3C7VnNN7/GnnownE
4s22azjd+xsN/hdLcr5ouuICulVxoo6MIK138Chod6v9ZQPqw3pXN2SaDjdyi0j/
Vv5+qpp9IbvsQxp04mhDHSUMGLWg8CADK7FpPDSbqdGw3T+2PmvJzs/M8hLckHvD
NBJ+g4lN5mfm98Jv+EgloJUlGN9oBbCOnq3brb//YMdItRXjqVp+VCvdSools0DC
cSZ97poV8oipm4CQ8q0o5E5LwiTCOy+wk2NISCwNm0/mEB6dMO9A3C2fyuQqZqhL
6u3Z5MOwOMo5eaZJcgBfDFYwpPZYomiL4DP1rCYkMJeJRzDpOI/1baLWSAcbOwgn
G6FuedFPIGHXzPPs9zHFIhk7pYc0bia9hoxf+HW+lrPBu77LpNYBWWk8C4p6pte/
xrCQDarCzl/KfqnK2/pfAGXwtglWTYu5X4WTt2sgJSfRFyRXcEM2N9/IRq5M4Sew
hBPwGKPiOoP3idBg9fEUiuK2XLmKWfcWr0XH3ReoaQKwnQYRO2TFErgaAp+CUtvM
DhZiHkHSXiKPrI3/g4v0h4bHDb6xt7D82F1wyL2orxpRDTlLiuwSZ2GAcay1X5eU
Hd5Rif3mmxHkb+5iH399scqKYUSXWIkrAbUxTt/UVi4FLjL6ZMycIut05bv5faLs
0ZyoFxaIUO1Kv21ft/9oOFU+uG5l4BuXwBXuQQjh8uB7J8y6KWdcWEbb5kk6Hb91
ku4QTZE/F/BbnQw3xWctnGMWpcH1uzuggJ/S3v2CnQv5TFpcgEyYQlDroMQ0W5dR
q1bnqUkVVkEReQnk2u7LUf6HcsyZxczJDV6NfmUzEUji2TGkcVKWoySgXkEc9hRG
FEe+dYn7ctfwJG0OtoAPrzKhIEcUYZHhJ/Rvoqs/SxM4r02eYmWOcJUnDAla92YS
KEDVUKXVRmstGFW06zRtCQhR8/RWRHRHsWLJFVcij8LB1khTUt9NBwz8oDg0uume
68VKX1C/zEiduAHgUgVAJbuur0eJDFrVU4h0p6l0fCKOZd7DZs3+GV+WJeAiDblr
jMS+gQckOJgAvF9wYzggT/xdt1m0GewwwtphjTLtLfHkJ5rALKoTxUGWLUYUwNi1
28Eb/Vf6tpAQWXOmh2rf699X59CF7jL8ssUsKAi41N6wImL50APZLLHJwC+AjmDK
xvcs13cupB/tlFegaaFxZs7rZ1f4VyOGfeSRwgm08y75yJ9Qp1jHBdyClLGLQcbi
iUeuzTKpnAr5YCIWDPfhciquNzMIXklK0mbbCLlhSWNYCSluqmZRqn2ZDxaNhiUJ
F9CaXa33y9ga0Ab/5emEuInvMfXacePnAGKN0NcCGziFZakf25ie/9XoSvUwlumw
wHCqBB+eD4VhpoI4SMolPydGWhM1STGQ6phAUiNkHRT2q/09HsM+MwPlzIdYwVTH
j+5ZHsC3TaKRpdCbjxGtn3yctsauaXTcD7EyWfVMVSH9Cq2Xifml3f+l7MDLhKlt
w6WlPqW3Z02rpsT1Qc354IdyAEPQpFrVEk8p0aRBMlIkvL2hjGMP4BfzPAVwY49A
eo5yEtto0W7nnQHp8g64ORF6mAYqmyJt9FvGOHQFgtN00Blt3kO3uV3+EKmjFjRG
5rXcU0ihEE4NhqcWMnKAgXufviaAqnvdIHLjmHDi9rA/bGWkY410TBSisiLO3epo
CEp9A7htwSPauYX8RB0O8Qn8JW+LmwrpnGV+7sZCHSBrUs6EUHSVOfcfG/HUNHQ7
2vXUXlHxA9H9b6P/vmXm9b9VPkRZfPkN0X0wgyUSdm4pACxzeMW7WSYqS1SwTbS7
We3O1pOb3FeDv0TMHaSsTrcaU2F6Mb9QDVxRuLC9hR3C3C+27HZaAgd4wdFAlq7z
lAQyF5+UlI+vmC9+Gm8Lvf0ppanItCGV89Y5lblD1FEuUpjODLEnibTala7QmEos
kO8VVTAzbvb/X68uBLCbpXTLUeNHw8ZBZa6mXHzRK+OVLgYy5l7gDkdnLj6Ab6Wh
40+BofoiGdqWheEzH67dG0YNMRyqz8pMAAx63pR/x/sHk/pwUj3rEMH3K7hA2FqF
6GtZsiLBJ23h3f3PZ7OrA41R7e3zcde8sm+cWu4i5WDHlz3/BoduuVhpsAMo14Pg
tHkfA4a3QBrLcgdz0dDjsbXT9Gfls33r2li5abL82Dy7evfC+5NBx6YZa2bpFJw9
TU3gUwjwKfryweUI/SGW7QBUDJeYRO+SZ5e3WLb8//QZxSiwZQ7Vlfi8NC+v7Tmv
Y4OQd2zxPsZnilJqCPqIZuhGm94y//oRsdV6ICy9xURb6sMzQyFx/eqFI+mefWq4
5Qns+w++wostv6zUAcWtEt/LpiLcvC6TGL/vwINJoxo8KHoNrBMPRVWpFCUnHUao
zyrp0VCMLJnWzFECrUZPThGqSM4a6bx37IVym8zQ1WyMxUgU1PZmHSLTfvHBwLAt
VcojpLqLCCbWwFUZ/zZRoyciE9UzMt3l3I88DgAEofz9l5aMUTZ2FwZGvPfAnqnT
kRmzG95s0OLiNn8faKNX+VOuyXY/ELZanz4qPCnLj4y4tcMEnP5lzmJTg098Crog
XVmpyfLDe3Ld6jvZq6HebU8klijV0LZiJ4KeipDG10HVTsXQWqwRrosQeLbuUaeb
iFzO/WlwODZrkDOpj4h6Nfu5okvH3tXQ3MbK9U06ptrMhnDNUIfPQOpBejuxkMhC
Ato9RZds84pX6UNXR003XIkbNP5rdM3P+JBeMu/c1gHLjN4iJQT1/0WsbmTEVmvy
ijGzqh9VVlM0xLU8mJ0DliQYSt66oeMtB2MVFRBmCnsy+KtspzNh+I0mNy0LAB2y
XbviqIYPmAkCq9wBRzddSPLo8Ee17FOmeut04a/7YgcbkuWE1/GmtUrE1irkRfhe
KJwPEjB6nRjjx6Z4S1S1ADjkOrVbMO8EUL9bS5Wa0k7ewJoX+uUV41CVfegHa45s
3J55Q9dQ2uF4uWAgUKO6PMXd/TfRHx/dmmZB3HphWjtBGYe1q+mZJiEDgGeWkaqB
i+9YIh1YoMRIvnWQ0ZdIvPmy9kRNGDqYPVpCPmO5ns11yN25zrlz0V2Ii+IU508o
d8/XIpse4/akobIY3LCn7vVKFN5Is4DUB6Tj487AuJcuAwDCIDxwXAbVcDELIN+m
RIzASZ0tncQMbi6UHVOKzq3SMberWx8F484OmqCVBvs5OKcnpAEMriABsbvtxAwa
Hj/Hyt+A2uZPNeVOZ4XIJkCvbTGX1cKRDZ3UpS1F6b6t2aDSr2gOA7n1GRj5FiIN
bZM+gM0GbuIwodxFhDZOrbP+48r7Ys354RVVO2guGC8bpNBNeE8+c8N84iITu5Rp
BaJCmhZnfGSkFO2VPDR6oOc8Pqdptt/DIr7dxnR2wjg8F0NCyA6IjefeF+UlWYFN
dvn567xwRL3zxjiRKkiZEFOlU6NWZ+qLmgHNFtjrzA911h+xLRvNo1ddJ2hPWUbp
BqEOZDALNwkiMJLo1Tkd3SVO/53rKB5op/YD4klf+Fgk2/siBmQWEPYFOwcv0eKc
W2kxMI85+zuXfODHyUqOAqUzHR7LVUjLte2B2Ze41y+9VhYvXHmkjfvBD4HIhA1l
34X9VN2R2BIkjttzBbmsK7yXB1QXdKkXHWdUv/XHra87cpXX6HjZylD2LC2Wp/lk
2xQ4t7Sw7wHPt4ZB3sEreG9YjB4HWLH798YfWXWbxbv3CtyaAMqBuOBexcpYuZ1F
cDQDiRayD949NO5DZMuaAVCx1kmpwvURQ9brwRU/xce5cKfzbQ+V4dPQkWNslbgx
GjQo2zXbwhApLtIDMI8i/360VqGMzCkpGuA4aw/DS8lXQ7UX1QxWny8J6BDrjaFe
/FnFv2eNzxqMxqXaZtg2sduLy02BxWnnbg63e01HD9HwGymvSjOppIUux8y4XHMx
CWjkvjke+dBTXKVcMU4v0LL5KpnHMfZrRzjBXCxun4KZnb02JBekZ3VtnWgIxHjD
3pNw/hGXpyCWelnxf/1Lxgt1mWIsdZ9zBeFZDRg/ReLFubVifdWTGWFneQadYKee
R3ffpKKzsY9Za9ZAf+ec7S2/Xa4PekprjPHHcoP69R/8AmGpYDGeOHjfDkHK55Pb
+E1zqAGFT95oS1conKtLwyLIotl37n3Kvjv340DRHsSMZp8l+aYmE11GsSYpoALO

//pragma protect end_data_block
//pragma protect digest_block
KfrxkqRG001Po/QIQF2JsI2JGOc=
//pragma protect end_digest_block
//pragma protect end_protected
