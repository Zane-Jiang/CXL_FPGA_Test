// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
pEwCDk9K4UVOJ1z29lH1pYR0TvRu6J5QDsqnHFvwJfgt9uuCM7w/NjIp6XUTBKMs
Z8vJh8lU6oIBzWFuMovPprtK7cM/3si2nVFaNkyqinIykwfDj2D0NZEoUpe1Kdek
JdjEH9tXtCZACVwmJ45k9YumVnQoNwEDZvSjpBCXt7I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10336 )
`pragma protect data_block
H3r+zFfX0lhNROIxsbXTwV3iCxrlYixmdF+8ZPBvdn1uf8roV8+hfi9ehuTaQ4OS
91HKxiCd97jxTa9x+eIp2bSLLA8WRr+o04JVAp08LggPm4S0e8uqKtIbA/UHaw7u
THdXMZZS76L43z0rUsqo3Alj3pTanpwdrQ+122RS4j+hp/Y2B8oyTbTDgDvh+/3m
G7klAJ5qIKqeKWRdf3OtroxkYvIVRR/qKZ8R4bXEBzoAroHwcwC0H8YKoXJauOfT
BCioYDdeo5p/LpiIsPDahFWNKB61UTNw2rq3NZnwjZ+yepsgsopcCkOF4yY/ER7y
XPLE0sM/fl4aKi6g/P2d0CNd76rj1uIQZAmvzWUx/BqK8NcKTspsKi9fm2Oh655m
C/IpAGd3txhYU8NuVA0zTmOvek6YvkccP+NdRjq0zUheJ3e0S/vh3OjjiV/QhOei
6xB10OuA/XCdeyE+3lXvmazTLHhkLYa+BYQpNXKHU7xCYPOO3GkWu+ZGhRkJfQ2z
CMtxb4cayiCnoiEdbhnGJU1Tstjb/5LxRXTDlJec2MSmM/Qde0O1/QRGqUW3CeYt
WykQiphSWIF6E13X1UN9ibvRbgHm/fYk8dKmNv8IBI5fx9/xad30uYeuSqiR7F9r
LqwEO5JiuYBCq0PlFi+GXM21jr5DBGsxG2h41k9k6vNhf68CzarFITAEp3p+HQgp
qTFYf2c9OS/W7Z7MVHpD82mU2afVTCSmwGNg2pLTixNUys8TZaj/YvZQqPzRb4zL
DQJKEaQhLNABV1O+Ogah/gaN8x/7pXeyfvs7e/Jgh6PXNsiLGbS1O98weRKYd1kB
HkRp0Pg5NIm5HFVoBCpouaMP18CaHosVnoY2bTQLKI7r9LRjv+FvMzvpLV7JKEHY
KrBS44eC7nlv6wP6Iv1IYRLurcHtfHJkvy4fOmvWO+A+MCSCJadIc9fP1vBt+AKp
Li208/urztUX0ZLYr/1Sr4GqVflvDciesJNUF2OekjdwWhngGONPitpsDBec3DSU
5e4p9mDMrbJFLKW+eVbdFNz52TR9UN1LrKQstw8576v6nU5RE2Gs4vUXO175ucGw
o7YhNvtUssQpN54Z6fguDHKGy1QTb1u7ZpqOS+wCxkbs5zQI15MT2pnMBjUHmSII
et+P/hgvFpSGwhsgTJp14HRw0UsQqy0qumovHgpI7ZYK8OwB64C8rjamv3zjM6+A
yhZVg0gmV/5ccTYxHWxm3ZIdBB0/yNhwBDc4dyjWZ+5ccOrJxRguVuHpjVSSFsLk
1LLhwp7HafPua0/A7UBDTtiQuBq0mOcDOXrbY6iH+mOA5xCSUvfDqleaL88U/OvA
e+i18EAuxJUOVbZ9r/w+yxBMBsI3DVPIDG8ZAPfKPSu46owVKkavY5b5lZief6jg
UgAh3Oe1ySIcxEDlneBbidToChgZx77fkYWcKH42gtgByesXB9VGzFsVP65wYWnL
TJxxQCyvMjmGZfgUTnvFP6pxSOZCv3p/4Px+n5wmg0bE6Tifwx9lKZHMUNNSr3X1
znuRPYrTqj3ZljafsVu/H2vXounKIr/2bSSVcyfyd4Dl/ggCnZy4CSVi1gaMvuB+
dP2ZfwaJihAl2mKCuJZCBwjod7pcvTF6Vsln0pyaVSQfQ4nSc2jy5bVR1+Cl1/SO
zatu8aH2+ts8zm1vGOddXxHGLg3P3RHix102ep9ubDk7A4qcPGhZX6XI3o6QY0zx
X3Pf7vS7DsLRJDtqYYFbQqrssS+HO8WniomKhmDnbjQtkWlelRc/0YrJpnLJZiy/
GVQPaza4M15Grj/n2in5VTDo+SraNlIsqPQv6mpDsTxZAv6dwg7RdCooCrVQu8bx
NqB52tP8ikaEh1k2MDrGc7mbL+4r3kBRnG8mDFzcOfv6yJxwa61Q0DSaAmQSIDwI
/XExfq69YMTni1zDlsQ9zLDp8JJV/w4lo2KTIekLmw08tTvX6XWcEdFnsvcffhPB
afDvBCfQXiREZsYJqx0A3Qqks+nz8mdsqm+eg58wJFd3V/FMsfLhGnaZl3P0MgYX
pCJcUYULwMecTox0Jq/FTDr/Ub55/laPZ6BvdYivqlpNxDHkF2jgrxajnO5BUsXb
KXl9jfSJag0aTRax1/0oDqPmxtWQ0X7OGHy5W37DUAVeMym7rnZX24maQUx5hWhC
VdaT4vAgx0icvVQUKhHu6UEMB9Vsj0aEMpcDTNQoqHh9SDvNR68hZpRkRczsbhy5
Lw7eKP7NeKv+i95P7CqQR1b1ycgxN/XpwBU2Up+SJAkCWO2MXzntPXMvz4EupyE1
dHhso6MtxyJbQTKus9pQNb488JTZKk9c9TFzVTT9z7NPewrmGQUqpMVpi4FC4PhV
1ZpLL4CyuCuhlhLX+KV7Nw2LwCBwuJYRcQ12r1c/S+lUyjqEUCb7iToVGI9Vnbwu
LBcS6VBLVy0lKd/6vaCJ2BZDpbgPEuINHL5/sgGnMPxojFNnAAV2g8jiKuyiJj/r
SegrhTkmDHKNbrR+6iZpIM5P0qb+Lf1UKn6DFn1EkmqEQWh8N2Vp5tPW+YjB9D93
Wya3uGUkYS1KZ7wowRHL8WA2eywP21O11EC4DXjF0CCkPFv795wsqI7C2L0RecBA
1CiDFzLWra70CNgWiGMkQhNUIjrbicx8iL9uT4fCmF/zwdJGq6iHbLxvD6Ek4jXR
41838xlMGgfL7g+Ns8YmSzbWSx/A/6WX7cNU7xVzHrRMHUvj4CmP/Ux3oYeFBssL
T9+sMPaK3DmNgNZTmr2zYSQp0uFobm9AgA1xNZKzKBAh56F/WaXRlj5OgK6OF6Xg
yMK2Kah6ev9e1FeK/t7r0t0+buR0LvlMZ87OWlUxRWnxcT5T/pvfVnvZkThu3roH
mJE7+qaL2H3w8TINIIcw2dFIjOspQjcH1JGntZixRPeecA8NUUxKM9H1cIFdz5Q0
44S2I5SV6JIf/2TP+BXCRzklNAZ/nnB257Py5UQPN8xXglLvglHtZdy4O038cW87
rq9J1zpGpdFmFkBdpwT/L/rMy7Bmg5nwBeNSsFXvpzixDN0Hf0STRmMRX9BVmAIT
2V5LLBtIvzJn0YXaU/tDA/6Bl8Cl+079VTEYRfOABBKU8/XzVnoiIPObXdu0MIVY
NB2FnV8RvR8XM9qBsC4IWHABXW9MR1g7+fF43yex+lUXpmyBfWoL9V2ao/OBVDIg
arJDC8iEUziKE++vjhvofov0iGzH5pYYppvje5v1oprdnw1AFfL2GRnssxs0ku+E
JDtxL2ptCRbodA9MbKz/RH2bw7IPvSQI7SfZ8UcxTORNFa6SlNOY3hoZC29vAtWD
TxYSt2ZEehB9VX/8hsiPZtH+IQE/B0alArgI83mu04pQZlUbdHwCurDS4hOUHGWw
hLJlaNYGv/8VMV8BY8lAj46SE4b13Mjd/qgZu/S8JO2QCyv6v6MUROBKEHYZPJ6H
5edJJmirLBgAZrQkVKHo28c9ix79vy9NTPMSOWMQTQVVjyn8r1Mkhfa8Aj51ksZy
btgtZHJNNGywroghTzj9D0JgkN8wXZ6SMXUOEzLYjH/CNEqf+RVccmo1425GRics
XfthjAfbVMmM6TGk8oTx59o4RuyRRDO6uNZAI5OlzMDlJKK1bAHhooiRpcAjVuh8
ej6pfCc/aIyDYV2/GH9efIuX4kyKKv1JU3+LNpjfa7Nb7TE0UWpIS0/Hl2FmeqWU
vYNwCsnqYV6ZBJMzyXd6qh2dzEVo9iEXKgZBonap84xpe3jrESVBsA5xEHutwYGw
SBIS8wyc7dNjOdx+r6EdCzeu64lXGXjnSWXWpAWj5mmOjsCJLPQjB08D0gtZgGwM
n7eWmDsR/rXY/vplFNZmI0C2kEA8XTPGRxEqTvBSH/bOX5ECQoIbsGAOx202o+L7
S6PaF+FjHHV4AA+ewl/VM9nH5X0MVqnMTaCJYWWKyYBYMNEngSB2J3aBcvFhJuYh
dpr24GhtdbfRuI1ubOoukK/86ZjIOI8o3HhErrDRojj5/XyRYO0TbkoLdXwg9JBT
f8gwdwP2eCgTrfaovyJ+uubgz1kM1qmN7MurDMZHtPi+0Q2USfwCGdgnuQhZMOg7
QbDjoDL1zIUJwLpChHfQOfXvbSgYLs4POvUDE15dUV8qFLGehThrXutW/xCBVBh+
vEBU/jVd1mOwe12CWYtqreS/n6lruKf1QLvUqbcymcDSe68NTVXzZJVmwJaxqZ66
FUDCrM5jPADIjeVy2o8kchDzNV7g0TJ8qoNMcDXN0XHCuYnGHt/TWmrv2xW7K9TO
z2JKDqgXfazKrgSyp2XS59S6F74WYrTJ+uAON77Ag0AE2jfkp/NSR18+H2vyxDEC
gnnYie0U7YLQhlCzZIPxhhxOPYjyQe+/SPShk+h163v4+83CoOEt0MghP9F6ygW6
QAA7sKTh4i6ut/vMu+ZO3Y2Zvx/D6NAy+LDeYgIWWkZMXSHXWKUa5BAGtnt3Tzuw
JSMnTAM91MfPAiyvNgFnQpzW4uR7ZbH7AVQ5ulX36+QTHeBqy37R7UDNS+QCwtt7
igXXNg6ukhT1cxT75+Yc0VFP3WBgrg2fzMJdGkgC1zNgJokW89AzcRrqGy2Hgle8
rkana1Zl5iu34lIbZSsIyFQPt7eMqveNTXZZUYsyNhmqKrPSrcxnWu+YDIAu+CGH
cUpETahGgJmZRrIeKaEFGjzejlWLBh5osYcuRJQHzioLNBcQljWwEeDUwn6Ggv9e
wvIqk4+3yfHwiLa1RY3xd/eBOymP/ef+y7ZBOGMPcy+qhok7RWZFfojsP1SrYZPu
USnYsyo+0ZyV6kVSFv24qmXLjDiIBXA6ev3uZq2w6Jqz0oLhyxevg4nYkeuEiSer
dI0ZcA8/Htl8qPy2nKMPgvLR4deFxaDD8iw+6UExp2dK0/Yxrc3WoXQWvfxR9K7g
hxuk5/L1CURnP1DTV4kfOtiv7UGzn7fNAmTKE/KuIFYqA3fNF9WG50qNYXrQHrK2
KwhAiM4myZkqfk7YE5nWEg7H+RRmSoBMmbVwDvfV4Pao35mVhxpQtHc+7b1JgXIL
tvWFlncS2yCkxHVaxp4mbzMFSBpnR0OlNwg8YVsh4xYZXXZPMkkH2Hz0IoBZpw30
TkmQOhTB7Z28aOubSh4WHWc5rNv37fHc2lAyDFyUM2kkC+OqHuAQKPdieJk1csDJ
Pp+wdYHSVVYQreULjs1UoJki46BUoHVRdBOmAcw5o+kKAiZyxHmOR4DXkMaA6O8K
QH2e1cBsI+o0mOZdiID4ScGPZBwqf312knvTPRhp1OYstPkBeomF8b92QMOtlQnA
quu6wiealApKQTQvI3j/z8hP9mOIm9YYfNo/y80+h7f+NQOHVKnTLpmW5aCpHM7a
NszFk9gPRDmmaipRid0xIvudnlTG7kVyb7EVg7Ff3SYwavpsUC7yULwWtKg8Yoll
ma+OzZQfstSNOjG1smN9r5I+Iu9BrtGXHuk3FMesBz8mUs6q5zRWzicXqDk2tZ8N
Eow2dB6ukfiUzcUeUknA74RvLRxnrVyEcb+/kB6cFu9GiTWMpdjBx/4qNhZ82UFR
8dSp1wwxft1vc+6qOyfe0iOnBS//O7G/9DDCHD4G6JwdGicCrBiEpxDKGYOR7hrY
GN4Hzo05rCAZsWkmLB2r8N+6XKs+wCXLjnC/AtLOoknUjyNKiWW8uZqLOQmH8L36
DDiMXsW+ecu1V1Q1Y82JTwppJizbj+x14HzBMkW5dsSvine1ZcAw07o3qDNTD9q7
+YleinNmZ2wyMYyEXyCsY75TRvZ22NJbJBOOHQtTZBPVVRX1fl90jNKozGbJEv/b
AtAs2bUQtvAn+562OpVcWO6GJNGGpytQYIqgUyqKQiohm0vOKz1WbHjcRTRDskIQ
D4+Cu1fmmFd2DydMTLO+vbE7v4PNsUaK3nWYNrooNlhBekrA9fuZD6UvfUpLZt1y
vE0sGLQPCj7wi0TSIf8CIiu+6JKYZMXShHxQaXYBqUsjCVYANuHJ7JtoScqqDaOg
kMJuEPSxILdFE6XEd16jZiUmU3Ua4emF6s4sTro9IurZWxvLz9Z5WP4l2OAT1Lu1
peThNYM5SzgpeQDP+bVt8TpcBJH3Zn4i1Lo04rqT7mcm4b1VD7z5i/oq8Dn22OTZ
LxkpV7cAW67DJ++FITBezbtmSH9K2SFi6/i2EJLLku8RzSMPQ8dCljJf06qYlgwg
jYclnf3Hn/WSCZ5YvQGiLe2gDGg1ITgtI1OGwWQy2TlcjW+f4z2cdSpol3WuNoeB
MUSe+p9XR+DVyz5pTrU/AHS1u5DuQyklaFXshSaMmeGy07qYXixoh6CqGgqXDMz8
VeuOWHrrh6ZO5VR432tT9Tjgea5+D4gNgoP5MR50ChkG1OPg/K6/3sw6C4tpIfvJ
K1oo5k/F++mOdA5KdrfmYc1Fra8W5EDY4lFPDvacjMwxuyOAgJiiAMApfPnfT+9T
mDvvi0tTOyH2lhiwCVolE6iAlqyF/9APs9fo/Rf2acXR5xx64eG4LVG+LCaD//9O
uIlfdpxyXpRmqsn4oy2H13I5oWKZe5DI/P2Dnnvs7K601rDQIXhCrSTDULxbAFas
wYqrU4ObcAHxCPZnayWNodzTfVgJxLvWnqyAScYpz2dvbbEeTdbjZCRx88o4OosX
oF9C4jNH+kpJJ7ekxw8SgkTQ7//jk+Awz1Kva/sm7DFSZbN81qo14qPZkkbihYCe
Y6iU1PLnsoPuCCrd/xFYwdeGkHb1imHdd7hHugDP0fEqdqljNrdlxpz9/BXPfeue
vXdNOpo1CQDRKinlry4Bg54CnuPy5JrnzwfzZA12ITpQdHvC9vM5tOi4l5IDavSo
vXvvzFVQs77IjCmtkKUGZDaSM1XK4Hvxx8lo93LV7njgOF4eAX6xj38L8UQyZ9Eg
s9LJ8FWtWkpWBCIL3UD2e5su+7q75SyXz9RF2FchqvfSBnyUFTKKU8snndzqidnT
l5VzYyAIXGNb5j++wSGkhaVZG8Frw0176ps6gWC2uPihGIzji30OLPcSFnkLMkA4
a3YnLi3E0nYOlxUwo+YEiT6VeNzK1QwnvZZahsmDGsk+3aP2U2djkNgtt437WY1s
p0osC9HPNuLmSE8gLcAWlc12Vzuow/RM9Xh+FWQGdo2HQsz6M2wbw7WXniz6l3hT
G+akWYIWtuSSdvMkAatuR/WnSOLthNqiUfHxzvdc2ZLFrbYmiHmCPrZR03j2IacM
hcbucwlh0VDTp/FzeQxqYNQLZC5nb2aTDUcG/H5xiOpJaP066lJFdD9eGdvjDnHD
gf4wJyNvDIrk4o8gxwhMEwLPfgtYIH4hy7Fub6rzk9fRoD6lteH/VzWitxE3/fYr
wAc1LbLMDp4Z7XTSdPN2+pkCNATB8tJJggAQ4WQWcapyIqRqNcvr6lz+t8X1FbUm
BHUvsFOm/QrcHUKlvStn0+xPQsT1FxSPvmk8T6vC2Fnc7xcTp2qvVsDW6h7VJ1GO
YWzTrkMc4Rxw4VffK7FRPRAi7fU5/xtlMjPOByhu9LTD/Ssaw3c2DXQLdcLp4UOb
6Wd/1vxashM389Rz3sXsVPk+rpx8WSIK0Ol03TPqFDhTPhAx1s5qLcEVugVclxxH
DvUjdhl/DemXgzInkX/eRUNdDMLeZSliDCUi6qIFknME6QIRxPq3nthLttlXN5FM
nvgkq96WDOymDwMdENm4Dhyow5QWJOenVnYoSATBA8ajXSS/h0N9pAtKqbYk+bLf
gDqng9zx4VRjSn07NdZ4qy7xpE2jvuwZNY4iuWZ2ScwA0kpYHi0rMFWEQr9ENk0N
AeXd+9+CIWO2D7bDn5oXTH4yeZDIEsYsGu/HCRo9DX5xFQJtXZMZoNVHwaeCYfYL
/CsppJahaYsBxqYZChRJSXokaxz09oG29gDhOZKpq6H0WboUkZfpZ+Vd9UM+N+ft
xG7aQPP2y0432FJrKU/8/ZCL3N0nGc0l9FI+BUS2WuxKNmJUA3gvjoDJINef1TaF
7r0uK9zcdKSoJOLkP1LcUyKENjjESP/fLRpz9aL1aLju5zoqlsJlrAXyu+jvqL2a
Ug4SfhSrKH3cX6K+TLTisfQNxu8R2by5Vp0NWH5+crImNzmo57XJZARjjdbnVv06
+sZbQ6eAnijwSCCGQjWEJGUaptMVMh/Oh6Wumqb6oRq8KwMADSEyLv0xkIJmYtvi
qXdsA6+A7ARdBIDy0wQmP/06oYDhPLGF0/b6Arss//8xFHmNRfO6CR69rYYd89bu
E5HAReCQhPpwfihTigOjfd2VQNtdXEllv3nlq8qRLYaMoQWwCrof4j+i8+lcvDqU
RvI/FQ4M2sdzTRYt0I3LFiBKJSuyRrCI5xteccmno+iZDzfqMNzrIz40z+R+RTle
DHl48tHeZ3/ubNzhKYtODLtOLDhbMgK7HqN96szSN8819J1aY+oxR3INBdxikLDI
waY5YRyMkdfdhAzQcQ9VeLzHgBBxwFOiq87IlD+Rt52mV74x/2UYdyQlejZzgMXJ
sscstbp2XXkSn4A0oJl49Oex39RzJ0AqOkCisa9PF21wRRczFMUuYGbFHMW57njZ
gZCckOW7vY1vEI7ggVgCtBHihz4Idn+h8jyH4jb9Ce6rO7JS5RIAK67At8aUfpWf
PwgO81FMKlVTWpgm+NXC7NAu45jYJ2b9hnfr3hde0NLQW0qrG8JoJ+F0MtLByHjy
oTwA3ETZJ/0zQGQmg5wC6vgU4d8nUQ9JLZV9JpanGxu9m9yqabsHdUtBWQeymqWl
JYysxQqOSCwZQL8MlmX70yVzGDYoGC2mCQIyNgRMHZbaSAqQ1FLZUvfLphsohU4/
fbIfTMpq3snWbw+s8vb7YXAyg/o5DrKspqi/lImH67+YsxPBJL1wSWuNODSSJaRA
cVgZ1Bo9Ig2dUOkrGPY59L44q8dou+60TnRqF3/mIdb/+qwfDpXQwcaqWNRgcpvV
AZdkmOyBUC+SWwppUF2cHiZwigUwto7/EzPX/g/UepB4esVVtHjF3EhPt+Qdn/ks
C9jfTn1BoysdJGDs8VpcGqijIYSc+AVf/RQDjhwQRzo7r9q7haQul/MEW9JjcDa5
e1DuW+MYGOLuNUVE4lErfDy4K4jvoHEwNvHwHk8LNcYKK59IHE0PodCrefvYOtQe
wUlKZjlyfSU0gyWaX1vqEJQQ29AqK/Wp8lW5B7HoqUxaiiuSZKLaOkTRkWw+dFdw
vzU2Z+gQ/UWMxkqvK1mYlk1RQW+K8jL+UKXL8X6pA8Ch5/TqEdHtCLJLtCTZ66g5
8+7N1QVvvjuG6rS8D9Doy2oEFzOW1PicAoDI8Gfjww4zrwUHhqmMeIg115URaqZF
j8azkIYrMWmTi0uuaQp4bKvx14Tisc/58ptFCickrnwzs5N53YW2grbi+/k2XhMm
yZ+whBGxDjiy0YBeHVy3fQW0ovI253iE21repQZmghgwklVy+qUMzAEX3oUkhwAu
Y958PrXvHBwzXq5VJtr3G+0+TFRDhc4VPGkC8ygYs8RBzPbvibmKxXXlvTLKvYAq
OOVOPiJnpnLTdwLmydZVkZmNBelH4uLjd0M8fLJFKEfzGVQcQrz/mWhdRfZtDdp6
kpzZJD2SIJ7GrVli/VWHL86HyVA3hnOuUv69euTVPXqjv4a84gOJvqbLjI09TZE9
ibBdqKBDOD/sAuohEb3+o5wzC4KLNbijv73GSuVhBS96/u8rZB26HUrjqKChUcYx
2jmi3qxlga5r3BLFBlkcqAZhjNV/8Hbc8hci2AT9nL0ISv9WTvkgKF3twA+ApxLY
CqH6fj1vyljUFcIrBBKvjeuKmpHgaS0/An0C/oYszc1FrVtH/XhHcwhsubfMv19q
3ZrWKk7CbIUYTUHOo3ZhekPh3in6tTQX/Irh1sq3WRkpQ2QtOpfeNbPSomR/uJ/7
6UYbSqPW4MnimkJRs10Ab6PknFvz5+xLvFvVttcJ/IOX30RkcK/2jpiQy9To1+y5
F/Zap1haYR0ArW4MB1MkSlHrpTIE89erXBVl7y/kxVtpDmY++hcC+RyMRqmZbn5J
VFOznnduERDlVw/ygQ122ME0ezRSm34Pidpwgx9MMLCqtW9In3vPfNkaF4FGuJ5T
aFiATBaI1KOGFQkO66WW59wvjGyXMGqm7WfyYe5YAOnLW+c3JXfNrkaNS6Ramt0R
ojDfEp7lrYXAIPGRWYTP9rBfdo5P3E4MCeGH1IUUhaO680MgDaMij9ox5U5QfsSL
T3w7Cy97OfDxAo/O83Bl3Xlr4kZPtxdX3lbjTHvQR8wwgrUCVmfyU4ahdGqDiL0j
50SVN6S/240/D9UXhaO/hqbdEHGCJTOmWK4X19mo2Moazhzo7+ComRfVE5RVrAsZ
bBHvZ9EoOaV4HwN4hAo4g6jNBn2yU5rMl1e618O9dlsvoTLEen+8F0SkGvurbn9a
ihGvHtHS9dOxsvOp4nWFJxwh2NxltCUxWLqIWGkDOpaDnEO0VucyiRu//Sn/7er0
g/IT8PsCkA+eVDPoeD+IN3meINZvdiezC4l6dPd8Wgmun4Kqmj6hA4rx3lFRYQ2v
p+t+PCNz6DVqhVLpiQRUPnmGYkQ/FT49uPeXu4Fyic2HrDO1a7SVP5iXtX0dfRUj
iym4nTRbr0gZ7n20MzlzbrJFtqBKz69eUc/bGObIIZphGGriVRdnTpO6idarcR1k
AvQJ1hISuhvO4x5Vmq2jJmguMKNgOkdq6csZWUzaIHipon6AkofNHgTtnBnKo0RU
aeByfrPaXg0zNZ1/yPiVsSQauwC6/QipyM+vbT3o+MTtrcf6l9mHcd4gwmbi/U3M
lYEfHH58O2PSXcPC1KVGhqDiIvRfv7t5908+ueUfiRMElCAEe4MpoCbgfHvYpQCa
tmJpPPMydPO1LE7MFauJ1FWaozSVVCwG+rmDwTK0nY6q5KaMdOGQXS9jpGKujbXj
QtPNamBMSMddr0yykMWS5k50Uij5EcpTXG8RjxjmGBbxbtF8ZifG+K4auIFtgJyy
yb8AgTlid1IZGx3+4s60FxvllgHnX08uN5n9ge5BxUKyqaKrGeiMF1nCIUIK4yT5
4D2VTpemNRCRTjy4EnALFVRHAtkwRYKCv1I/00mIlE4zMvP5tHMk3VI/NJi/JwMw
AmxPMQtvBpdJk9Dl6+bKXWKhVAYSBlU0liOIvFy2BJzZsjFS5W5sP2FqK6Uh6PRk
r73eYGJFP1HDkBsWDDsr/+X8u3Vq4X3WOSAtoSAQzAKazvQJY8LaPJTIi4WAEdVH
Mh9RwnPYTT91+NzfjnvOY9SGOjvHkdyFb3GsWbKO8TcWIPKpbZ59718Hf05KC2un
ELFrtnwovJ74Sx18ReEYZU2a0cVtrmzv83Rqrd7/N0bxzna402Psz34VxJzDJ4ro
H6OYLuo3Rouvg8LqIHK1f2IXsDh+F16fZPoQSbmT1YdZ/YiMFBmFAxzolg6vQM8L
NlPvliD3lechrzGmVCgFS8wyasEnkFcnq7ITEAJTX4/ablWIeV9NgSVyQTidoLTJ
ayovWghF0gf1ysag7xGVMTzNyabW63P3tA/udaXbB1u4Dp1OWUyEKsXfEC+1s7Ip
krWwN6reXcB89NRzZ20o7urJ4iONsXt/sHD/BEF5aw6VUKgyz7M8pks+PjJo1D3W
OSMQU7k00PLDsjeE/tq1Wo7ayZIexV1B4/2NCh05eovjyuqpiqrDyev9/yEVBvpU
g+vfCjJyYOtYUGevieuYRfEKj+knCdFXpxRXTaHNbQwmF158uwNrwY00nDBOlF1J
alBdCuLwo5SBIcgXtzYYKaojWC+swSw8eMWWuBiOZ7oNmKhmLg0wRAbP3iNxUDLp
3lsxpcpaDBryGiALZObWfMAqGGlWYz0yBNiC7XjB4rANhgOUlqJS3fqYUf9XmtJu
8itXvKqVlnxpdNuTKhBrZU2SGLoBbrc/w6PPh/1e8vLzH5JtjW7QGCVirb37bdos
xqeVTKDQBBFoY8ULMry23p8EG+x6mMoyAHy3XG1JaEcPHzhDjIP/ZqTk2+yN90TH
wcXBN5+KLk5aD0EQDdOGG0QFkCfy+s8MPEytPmC4ROlQYx4QudDSCorNpzo8Mj95
h8czQMlTBzYqcg4/f5bXctx0ZgmDCW/AQXBLnypK6N75jsRQjpzZb+luz3C4GSsg
0YocuZpeSR2XvLk2XIaZiR1P8JbeYmSrA6eXJlF6BIHSKT6qNVSoJvSAfLmvtuLf
n7xkH4cJtwEMS30ZFN8eTbtwQgRMI5loWd8y2CFBiTEB8tGKI4k6scv7zM1c5Yrj
vdSBlsxW5SSKM70xmAR5MNMzr85QvdOQChkkqsIrc+kh8LQi/vKKFo+njKsDQTmq
mMVn5TW3HR1DDZt8GjTGkXvSeQm9BFnts3aCNVRuKCnUAZCul61wW4pPV0wHbnWu
ZJ7ixuWURP/5Y5YvJVlnpWIa9uPSZcjum77nie2PcwkM16LZzchdh77QyNKwT4Rp
d0dEtlZkqmoi11Iy/ffBZ1JKT7FrI5NA5FcbysBcXm3ND6kfa6hFu0oLaZeAD+CR
vTMlDlxykHGF0GNII8BfyoqIu6z5ASMKmZz3CJnJrfdPFqMPIlsJnXrUX+0ym3UE
iXtNH/X9qN6QgJeBO6GfFU3RbWNVdBB6JbZdsNwqQXJPueAokZX8kcqU1oZXIjyR
Me+AggLV9JYMbKU0cKeDBVmi0QGbJC2cF+pCDAJw/iKuqhmXLHOMgHAnzi3eUEvV
DELRIGvBVU+qLctQ7vME2XsmwRld2LC7x5CqiOHenVuGzB+ho4yrw41uSALTEZiJ
9r44JGfI1tklHvo9ly7GQhq0YNG2e3P8IHhFSGp2O6JHOR7alZCsdToPL9cC3/dU
fhK4vsvcfvq2zUODnHRw7sb11pTpK1QMvrZI3zfJJMORB2RauxH3W3x0AEfs2wm0
2oYuu6nOnvBEv/5ZbAQXGq5TurZWWuBNWSsSZNpEmtmS0fdzV4nBpRyfKLjCJIxA
o4OPHRRLFTN6a0byOPwW66lCJy/TWDgy5APhVMnGJmeJtYq4rZZxvFp3rd7nG8C/
OdY1KegdJa3ybtnVKd7GBb26niOr/ObVhDWVk3wBBe7Vxr3k/zDjMn2NVvuyzMBp
ePhjMLH7Sq3CxdZmNcNovOwEJumIj0H8VVOKY6UaaOzDTgBaYiDfBjBUz8NeFZ4q
SdWv9BllRjUaSbND4OH8sRcDneb898Ij1u3fivUUdiRCuAFg2rPDC3mP3cgRCbo+
w4misu1/R0exOmOrQb3ZsjwOWo/tjOtbkgDt9wXNw6v8EVO8RxF2FcqtzORsWwYP
l9JXWmtg6R2co7/FvLRt+QYquYnDaqF6HcyRGlomCNITptvxfDpP8B3e5IHHef3H
U+baHqyORYHpLud52lGlG6EKoYELd+At0gcYezFybJYtHJgBwnx6UW6k3+UrTWlG
rUibxL71flecphOZ2v+TEJQAJrdRXyLRkHfHxTk0p6ab7UcnY3Cj5ewoMoUjnJTC
hHAGvxYhF228GtMJAteEzSAWHMPRJye2qFuwmIa0tsbARaCesPLcb9jYiZR3GZz6
iq4dzKlzcUW7yrJrDBBnAEDFeOpLw15jSW4IDK+phLWoKhYDGbcJE7WMKCHypXSL
jhYo5MNkKnuWs9zLHeMgimuiZaGwIcovhpQt0w+22RgOXfkQi3Mkcdrp5C8Tom8o
bs5KbDDPlEdFiu0vrsUILH4hEK7v0ItrEfFpEUv8ZEzxCtcjDtX3KpqtHz9GZKCP
PdK0uSgTBBYMONnK41hiMw==

`pragma protect end_protected
