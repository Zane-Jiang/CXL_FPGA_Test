`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
BRmzp1Ndjan+KnetM2NJ0CIB0zq5gtcKC6QBsB2jpWZgJ4K+o/MKtHLLpKaqxuA1
9oxceYg0YYxjRzjDv+gWZBYdJ5+Je4K5e8LiNAT+zeTF/7I4nJpdWJ/gqOdt5g8u
P6mFlt5HlhUI+3lfX5t/NNvJWc1Oov6vFxWgGgssc6o=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 99888), data_block
CjgzS3TSQky7E+wena0ZA0ie3q0NY1643z+WF9gjFDDqXPKdobAYmRWk3OUAl9jy
5bR//PjT3ABEH6iNnpO8Q42PHx7Z/MuN6qp9ofBUsVlym008DYNrd+mvd3cQPA2g
mMc1rH7Ye4FyYknnp8HHUTobkxb0TWq8E8ZbhX/JHz5yQSUOdMTdgjHhxp/0bdtu
PMEAhgOhA98VQlFNVs93abMN0Ynm8p+s5zXSQ8gbuyrvwbk8rZhdmTWSmg4HqAXg
1wGgPIpD/ZKZ3seKU8LkFgAYpC/emWhpIZ9ZG2LnwBb6fG/BD1l7hnu79CR4HAHh
KhKRWaZr4VjTKW5RfC+XpzGrG99taMZtO7CBErM+2ZM+3k8ahobPtxPsnRCZxT6M
wgNMF5OHvlD0mSAYL4DsU4RNFATkHPP0FZs6zuJ9m+bonBkeZhViyjrXx40I9SQu
W2sJLhSqdD21pjP433o9QeUO66ercpYX+ffdC4QEKL+p5AGn6hNYGQGld7upMrXh
tc3JCwPMoKQswoZR20lO1Pgsxuij6fjk/xMXlk6S2xyLuevEYE31pq3Bl0KruqXH
UfQpJQBZjYDIY5zUlfoCFe3ArJsfbztFNKWNtbrEtiJGcBLfVl5tTtihvZdoxH/y
ahJjQJtyqYF9CtuNiCM5Ngxy4XNsW5yGu3ntsGMGijcUTwDcy7/F7e71GgdF/Mr5
ey45tHdO5d4HzFADwxG2tlFcsabApMMWvdAxOmXWu+NGgmhGl/onN/xLmmnJLKcF
zY2Gplz2/M3bqEG4f8FEVS8EZ197v5jw6MjgTQlU95kXhZD4/Yurq/vuq6F3JkWy
U8SDcwz/+TDGbohcm7wFhJpCQwJMz+V7keumcLcuJ14gsTW9HVIezvz4QwLo7Q9O
mXM8iL1diwSYkYSudfuQA2DMTTTbDh6rA1UcQyRnvojkweWEIMJYzlA/w0pEdL71
ys2c001YCDILr9MFIS0c7qr8hp12imVWXZGFcpCiB2G2OZgCMH5B/mDUFDlZpRFG
xJ7gwCNtj2KFhf0LyfZ2q/jx3w6WgnzVOzQKM4mDOjMFAQdcvvGaQIlxMLc7YkPl
rbRCBANe7+iSVacd51ok3smBhUHUAwac8wfHcF39c57PCgmzxgfRepcZI6B14gfZ
5LHxl62aRYSmB3d4NuHFs9G7dms3YKSzBur6W5h7vtj7TmRRUKBog6BSQ0JmFQrf
cThTbVuvIvHE6fHEyujjZCA7IRyBT7sViH5FLDJ25KvtJhisk8BwcW9Bb++A81Qp
pBT1UJYcUCXx/rr/G7KLDWwgYlbHyzehQayHolTy/ibuAnd48i36uhFp4XA6LapK
1zYiORXrF23Zfol8jdVucE3huwiQK6o17BQG7tAlR/5taI4dT3d0gvuXO2zAgddb
lGLszqwpW4dCAQiY/dv0mM8ki76ozNb+SUPaKEQaEJxNnmmcD2tmANXQYSGIKnIb
FpqRTnoavAGQtFCwmOb3CwiIUoQ4hPHE3n440cXne+/8okWOEqf+Pd8yYslmPF3Z
AWiTKnpNQqOH3RsUyaqSrmod+wR0cL3c03/pZDdrM6enqQ9UcHxfGw9fsx9pdC6b
CYwES1dauWiyf9AvcvVrp6wtODAMqKgiPYp1QWSotmz/+tfAxMJJ6oTuKp/dFSE5
MsxRmfiBnRF3KypqBaqKcjMYybHOID3NZvI9Ql8VNXHg8HgG6kZmUStOObq0yWJJ
cQIYAm9UjU3Iyodarz/1zjBYe8h4fmo0jCXxWKXL5ilef8ThiN8p1x4xIxo/vocM
KJ7eSgv8dJREYp8QkjR0tv0h5DadzffZDrBz4XcnYI9Lz9sIx/qRCFGX4kwgwaRK
GD9dxLs5FsQ3mO4K69sL+ISc05cAAOMCoYyJ2tsuCvh/3xeczFUUKFRAijHOWc1l
xc/M9bsmCpyEdXQtamyrGRpa3Iia+uvWNImTBPH/gdKN9AmtAIukRleVZ0GMlxD3
eAEANA4VSyg5vKRlNdvVls7eDP/OcgBjN/yNlAOtNnGiXHvoAPsiRYyVf4QjowdF
YHtDUL/LPA3lrivmM1h9LU72qbJxSaHFiOy29a96G/1NaA3cJ13gkyiFJV76Evvg
mXu0R6P3vPQTN+LwHGyH+mklWg59lUuGzCobvtRW46iY7iOT77ruR/GICXGptCcq
I91FfhBUdFHiG0GQGkUlqkMd0TwPAQQ36B2Hs+0RbraGoSCa611nCV6cb6e9SGj7
3ljT3VTCWbfl3wVDjPwObb93JtkeL1215iwR3f664tna6p8TGpEVKedLuldsWV0b
uV0meH+FFOzQm0Jl7+Gz9eMJzsrIfWQ2seCA0lmXdx7XiT3Dgk+ygEm7uoGsZI5i
DjEC7IDFhT5d2xBBEBHAmcEXPOaZnsjElACJvluqaOmTkIHFf+SI9X2VPNaCptgI
X6XQ9vYnDiu5drH11N9Yxgw5uXPAl0Pmp5amrRwCnm7NsPxAEx36XavDZZ3haj1H
TEqDaer2aEzxKjhUQxkrVk78KFUzIZHNFpy80hd5YiyBpF46zHRFlp9wzRbMOsx/
C4XfQ+PQKe/CN+5oxCaWDAdl2SzNUCedtimLYpai9GzoLD4Lz88zbV04kxPO+eTc
UrbowvdVBwjKDaSyPYBuOBHyAOCyjxnELheZeOH+H0DcfRGcBmNBBlZ59PPpgLN5
4EPbAK8GS3u6jw2h522xZT0sYj5qpebfV4D+bpnlv5lAFrLe+u+yRCMZHUTmJfTM
u/JKdpc2spLipbigslYTO60Heml6GfzPs1BQm4zA4LP5Iq7H3TbZsZ7mDEszKRpS
tGnKDAM5sEMYZkPq+ooOAz81UgVK2ar076VfLW/ew1nz1VKpeF+nbdWSGCxM8usG
HCHW2gHlbCsIBSc++gh2sXKqNTCOg5dpnUzeb8P5dX87Dmsg5FqmGQ2OamoVBG0S
W0H1MwDy2d+y+tS9codZQluEkoHuWpjTX6P8fTqNa6gVWEbjYwyBbrXxMGglIlI/
QoVx5Pa977NyBUznouwDrJr+gjVAN7JHy6GzCHjmi4IkiMMkwmckK82+pPj8vfdc
VWkkKO/g19djOQlRqv831F8e5MhjztIly/n6g2vbKB7wLUPyliNOvkOxE84BeKnI
crLaP1n3bAuxcbj0JDZcJRvyVgUDf+yLHPktkk2yJlFpsOYOqylpjFEY9yLQo5+1
jOvXeGI5RpRHRwxn4ktVYvhxgzXnMVCOf8iWIfiW0rqRxlsUAaTScwDCN0ORv1lg
rnDuxa2np5/u7e3ACQz/WcDxYsEI83lM8iMTd3tFI+NHABH449E9dAHmHkfHV0Jm
owuqKVRSwi7YexUibsrks0Mv14ELThmpEjZ+P3lIjGgEBykfzDlpNP2nmHvH51mG
I/mW8/ROxmdjGL7SdmfB7D82IAbCHXCEpwaXLBPa2uH1uMnO/WZSMdjAU0xNSote
Xan1UK9N3yo1zsu6/MxY9j/r+fuRBj2Y4saumF/zmRjMuZUEcdDPxtW6ZqgSjYLL
Qkg4Z2i71XMW7BQMzLP8daaB8H4zY8jra6cQ8OJev83kJLaiRXDvMcTzZSWmu6h6
/ZrJIwOWppy03aQwE+93uDRVujfO2fL9nspbsnJMjsen4+8pw4gTiYRJ20IwBp2y
DXDeDGFbbEhJFNBEVei+CcLyFkScTEdfKznbxADUR431b9Nhfb3fxalQklpW/nuH
955g3hiYssDWdMAEtbdYodiVxoG4QOUz75cpUJOAGbDFSgNIFcETW7m3CBjT91id
+Kw38jGHt6I4YY1GlymbvLSmthVMLHQ1t8VJqN0+gje5HcUC305qH8h2E3FBtPlR
aeliP//uv9KxM2AQxLEuX9b7hZ0OW4iYDQu9GZBDiPJohJrzSgGtk5sIAMtXBxmz
QNf/SgNClrka8LXXqh8J2/slvHGRqJvPJLMaRSNWG9o34RTTx4mIkFq0+VS5hJy9
Uq2foSFk+NwWVGHr3Dh2Qq16Z3mc4D+RwFTVHtK0bRE4OSGsgtx50HSRxYD57gu9
Jx5WRTwwCqFf11BWTKkTj/2JC0sCENW1+gqH6N/hvBwTxavcBQ6UQeNEiPUvenAe
EHMuL831fesiOSq/cxR3Vjt1urU3RVVyokrL33V7j2asKtNbxzHr1qlTo5lAfZok
kT+z4ao+fuK3b4gjSGkd+M0obrYlGp3RFBmNYZnv6WgQRqzPoYpTCnnc4p/73Uup
toX25HImKvr6+DnViirgYcpYQA6ZjvLcSLWpRPuVyOa1JokaHGvtvyfBO35Fm2ES
56QTCeGrKRpdBiDa+Xpde1dPsaGCGfOwoRMBMsR9FbJmUX90iGq4xcf2S8eHu52O
ZpMEKSF5vifbsqWadpdYAI1z+nXsBH6ff5lAVNPV0wX615MSjZ+2kcyxoMbVUpOc
9AH3wI31TjQzqSj9tZ0z6bumhXJiJw9aMo562y0mj7fzzd1VbV+8j2PcVb7G3NTV
03sBo+G8Bh1lSLLw7PgIDQPgAVXWKEiHzZFAXTAl1Yr9oEDDvMNiHoVVuSx1VzmT
xSaTKtZehyOJVVGtp5OYupvogadp1iG4tkh95OORytCvWYGrycv3EGGQOUtQbqIH
gz1ubSnuCSSv1DdV38rtYHr9JB16NrEY+7ZpPDL3FmEBQ4styeZ/K0fuGA/ggXz9
f8hk7QQpLayG4h3M23FlAakHpM/0DDKIljXn8s+S6nZFpRrrIEX8B8Vb/unkHMkf
quFtgZYl0bEaDbtKu9fRNzRfOYk44DWjPzyuKO0600TAot+2X4urBW5WDSQx1V1u
/fU4JrEMX7oyqziyqE08Uixj+6BUoY8Kfb0acn8hcffqL/dS13yJUn0Ha4DvJ02i
pToKPGj4M2fVIWRsifMmV/wU0lt/dcbMdRmqIgPbhUv5cI12bAtPFtBLT9TgLrhC
I/UQQvPGC5N71OUdVvIxjeMe73PGGi2JgZVB4of/TSOwOEwQgAmQoIqI+hVp5x1b
tVFEPhpO4UOQMR605KvIrmlqdL9wr7b1cDHRRX4ykTtmGBFU97pOcAdLFxza1on8
a/KGFLuYv2yJTBzOHxVcdaiFjnsqIR9Bsb1pjSLcSDbak/KFrxe/XhFh6JOtQBE5
db/GKvSEGGV3xssXFHjgHPDiwC4tDaHM9gkSxWRmNkcwl5wdpxBDQY3W+awi39OX
+h21/pSNZ+bXJD/W+QRF4RXpWSs1HMPLn9vX1h05wEL8Q3+XFBflf78fAKZSVvPI
p71SJhx5JsAiJjfidaVQoIQhrvrypQ2XzfV4/Ls0Lg3lF78/kBjAZZx7ChgHiiI9
SQf99r2KxCS2DrmHZOYlvqY5OzP54JtSKGon0bL3/vOXIqqkMB5MJCfe//4qM+aM
stxRWuW+jwmpoT6W6ULHeeUm5KjjThxRDBELo9azX+s4eWVCXlvB1s+UNI/8/THX
d4XSpJdvCdeDHam8L0YkDhjq2EOvLDK8nlAkg/vPbc7SJ08vSytgtlLjI1eGuPGN
vT7jcUYH+fncGIKT5u7o4VTZEEPaIX7AUsQa7/1FdBJ7/2R+Ss7TBGdIWVELjA0T
DXbuxBIhTzg4M6sEEaq1TSUNG3a+iaXp5lolK2tCZ+vjrGRC+sA06ZkM6iHIfJt2
6+vrUZ7dyz2nGo//l7YvuarnF5Ty8iuBGesfeS26SGj8pUgL0o8lTOakrOo+b3x6
XhdTzGakiMYFCyNKZiS7mr8P2v6mMkrMKQBV52nqUWuwtvbVyy/TjOxuYsaJ5p0S
9fJ5iiAt9xkTLPw9IhTp8oYdlGPUe+pfAC7tJ8yv6irdyoI2ZUv8ay7gsHqRaS8v
d0nBmu2Ru1afO2/lnwYEKIHYqWi1Jj9ugQdiPBqXO0NDa0hJ83zKhi28ysiF6zK1
JRU33Q/qZzFSvh9iDd2SkWybCIZ1p+vjLcQXdE6aJbTMLaf/vtm1b09B1dMfskW3
k9FSz8sqi0sZ7rIp0poXiyOoX4octU7DOgDiG8/VygYme62jUUt/NOVAzM8M8y9d
k6ajZmGsqCXtLFw4SqYVbKWwNSy2gSFAkaWbhQX6mNUdSnLRKf17N8P+4tKkt0YQ
YxG+WeFTvpnrNcKgIceEZO+lJfgh7rI358edKtQx4iFYcNkVcI6+RCLSztg/On/j
nqUnLX9qhLefvN+nDpdWyocb4wVELGIWaY/PiAUTZqEQjjigjwnJ+xcK3Qt1E8T3
kZ9hxIRP7x0hE55ahHZHfgPBSBGRhIBw1mVf47UTZH51xfDU2oH+/mDKEYRlreoQ
9iaUzM0pJqjv4GIdT6XeXqypA+FaVqVKkUotAHtgC9Qb7ij8fNwB/cTJ47zlxW00
4WEdRLZqlfvnrlwr9Xce9uNocL68NVXVm13zNUjeSetCoxgbvA8GiWrjvzn0024h
+VDj1RrBAb/AH9o03Crxw8yNWl23Nq+vQOtArE3mNrwoOHm+jsQwQRj/4oGBx1W8
HRTIcphZY40iefWBQ32eHkwl3mQy/Mhh+Zrb87oWq169Yh+KV2qcC0RNguBhyfrV
71/EJGM+/R3qXU26wlstQqkzA+aJqYssA2Ko7GPxyUEnlZ2xfuECV9pEXCl6iWxQ
HDmHL4lKKhIkuQX3h3vjnGOZxCylZxrLdiaksYChlmrciXJeH/s4hIRMwpzj5if+
ZLlATKU3BzibyCGYiw6Yx0hTwS4E1lVYSPM3aa0Dakx1Pz+oP8Q719GQLIKO/79v
IELusvAHoeCPuoNpY6zszJlqp5PlwsWftEfdXu/Ma36OVooOPQ7vZq0ydURrvBcb
VozrApJTJjtel/12/t54X8Q53CLKdi2UktLjsO046k0YPjReVX6YXobWgtGIjoxc
2JMrZwmz+Qa+234Js9g8YMOAD46pjFG6jJvEFeQiCjUMnciwhJxSnlHYXLVclbkF
VBVKfnuuW1MeE/FflTXf4hiWkojAjbPT1SQRHqIr2ddAarCO9y+R9bACWUhIUcmp
hkg6UNUbBdiYpvzlvyUpvY3krJ+yVbANGiuh1aWDzfHvat/t7LHYNRtwl62hzmSp
cxUIk4EiUD37qOvhU+Q4qvGF0/fFlW38QpGah6nTcpFBH1pNdarA+sQ0xeD3LyK1
AbQVObOWCwfa36HFTCpiIAAG+tIoxNmKKRAGDbo39IvFv/HRXQuRMBHmoqG+HDvz
mzywc3g6C+/iuDFHQLrkDpf52+TVzuTPMFw3hH349+tDBzsiyGB+B2UorcDNUkJq
TCN+Ak0GPTeePMG/r49/DhhN+4RYumjKOOIGWKZa2nernNRKwDfRh/htitC1W8vt
K0vU9GMRq0RQQasoVwFLnFTleazCvUu/fkGXAtBjHj0+YQeYjXr8EbyFK+bsxd8U
zQ5fnEYC1Y9PEw4hxcSHUjy23LrKEEI12yPNlXEeIYAfH0wnzTsjPE5VxSXf1Nd7
We2+ocbwwlWbuGnPuDbgt+ckO/yn6A+yrf+WwS/sUryTdWW9ZNAUWlcLWOlno+tE
UIBqdharod5fBpOl7SfwB63KeEfBRIPOZayYR03uR7SvREJWVxbS3kteKHFOlf/m
TNwYGta0tIiN5KsTvOy3zcuege7ABHu6YcVMNvXi+vvPiJXBHrxj79TLmsqjh85g
nPZB2H1mdFwGzWFTTz9yQb17xnJujYwWy4nALMxHyjxsKKXjAkbS8iIQzHZtC/r2
Zd49iPWStnzIi4Hmz8GnbKqVcL4QtY1sVGV2b6p00puNIIKpOp5lmXOpdOGA12vZ
mhiUJCvv7QUr2MFBjPYxcd9cDgMial+t1I53M8HxnyEPT1is4fFzVItNvpWm5hYU
bfdq6y1qkCDSYKue6D7KmFpdvsm9zEbe+Fm7B+FDVNTC3C1ud76t2+ZXfDqHCHHW
fgrkyImg5o7h4lcv+6U3H35W6JDVRDweqv2zehKUSvEnt2afTY0LlGRbcKN/yEIz
WbXXM22/cZXFotY/4tXWRiwhdWcYAk8PR+FO65vG3H8hohYqJJAwe0WZjkDk03ZE
a6ura71yC7JFvF/ypJ8fdswr7PXJo+saxdN4Ea3VhDaNi/Bz7R9Bni6YEFYehZfH
91/j+1S89xXP0OOjcuvyTj5K9+/l2PNLswX1uVFK3KJp0uNE89CujfKxvcUe5RTo
3jxk8XJDzvVbSW+2u7QyAphJfFymKdNZzC/toEroxq4FPkauV9Wvk+91CdGgchsZ
NotxSsZSr5ZHoz+v08dXax+wJL/uNm0zuLkczIfm1e138Lvnf0mRkqYXZGgzW3yC
5GhIRDWmZCvQZ7ftBKDn95Xug0Xzk4+CusR5QZ2uLXnPwwPBotycuhe9NRnea6sj
egxhIkgk9GAenOJS49Pz0ivianT7Yckg2F1C7cXUCcTIFJClhbtU6OtuzDEQqEjB
S0hdrXJOAoi59KUkesMokDIR/ckzDbzcUW5R1m5LEQ+AZMXigFUSqDC+0P/8fhbq
M6yw+QNCv5JswxQ73uLEZugM/QbOFUegIUZ99D/LhnhWfvi/zCSzF9Iye5ARX6Rj
DPClE09hS5XrKnRU1gLdAMNL8Vt6FuM6Y9cGlVdVpPzVU5p4DUPuCa6Z00PfL+hv
1gWsYhqBQsqpPgyQ+E4/ZtE/s+Fkfj/ZydivxCBFfhgCwh49YdFXYgn0CKb2hF6u
hu03AXQ8PDyy1f4/Ay5YEIshH6JeTjYpYaUoq5eLZkNOtNZBeeX5QNvdDPRTTdto
H1SOf0gz0vuCN9pB64s8XLA0bqktGWSF5CyuWDXL4vvHP8e1yfc4aiKVMyapx+e0
pPVKKfLT9UOXppBSbyVa3C7VrbZbJnbhYtqqGaqAZ6K5KlSo2/1woIAQLH0FJJov
Y/hsn6DYw4MTCgPrLg6DpLnJi6gBNvr3oZQ/1TF8wa8KzGK3Qjc5QUIN2WvjonaF
EpgYgQhHG1UD4Ln/yHyK20PniF4yiDEXq98tTv27c8tAkr/bEFeHLsYj9C2PG0+6
xAJSuSyGer5WLBZc+cpHU0+2ovcSwvg40qjckR9KuSEPAFmtXEjf6ZnyYy6+o/aK
ytpfTEC6ViH0jLfaj/bh33N+GtMPgUz88T8rsxgomCtdszDadBmyKAiJrAkvyqV7
Nv7CjVAK+5PYz2WlbsVAVcmeu/UR6GpSOMSkGLMqy5TGOatXtWhffOjWlP2MxkSu
5GI3Vg/Ac71+f2sdTeavN6sjEobSQSonMann3ExmW6xpF6mE5aSCBtk58w5I+cSI
m8epx6s28lVYDkXXjLlWii7jW1DjQhOR7Hp0bKIXEn+/i9jqcNEs+rY8/zd+ywdH
5SHgW9hajrwS6ABcs2jo6hM5K7iepb2qfIMD7Ec4fvGmXG/ND9kfJXBy+C0WxZsu
BgwHox7g0e063tbVif4gmf43q9dgYQ4NAk9fNULErj8Snh4ZDoPObBp0xQJYgsiF
hiMBRNnT5PoVWWfTB0BW7x1kxISiTs9d4L+cMmd+sgSDSSAOgtYNJv8wbI73gUYl
gdIa52KhbQpIlt/S6lx+lZW+AydTkUKyzvk5K2AKkeuQhyQq6hRBi9Ls9/Xf0rpe
0k/47g4EG8bCqsaf2C+llwuSFrOnPK+XplWi7wmxy+AfXakbECbihc3sPR4psPzq
WBKfdexK8QXsg3YipcpDunJZSBHQhKi0lFE19eIBqHG01dr6ZA1fBVliERrPXvKy
zWoFYtQEjBTHehQChoyfj/Cml6fxp4fp9x+nfi3tjJ5Mvxbz5l67m3FImZ72SYhf
BUC/Ne6nDyKb1QMnsVBaGtAQUlRh6R0gYmESQ2G+Q1bHCuXIHLMFw8gxge69ZetC
/sfeULbTdAUFdaufDVJtQnX85/h7jCEj67b5bgyf6nTdUT1u6M+aFvGkWR+ZvaBl
lN18vQxoNlxvejygOTNvuDg7L77rift3IGuBiLdlyJJWTuWPGcjn7oQwyFcRWb2j
ma3eCK2gk4ikOGI6ast3FXAY4lAlW+osXHIUKyWy+Nk8Tf46o8wCNxD9lsz1pa1Z
RKEFaLn3IFZZA3PcFH8M0mIgWHWZd5Z6849ASb19294rBuktu9euWs4RKghWJ6ya
nfsD7Fv29wzor7rdKNaODEMrTph+a3IlTIax+RoaH3jQO+lME461aaRpWDGJNrsy
+8H7fsetM4f0QbhJRY8zCnw9wZd5TCsS2Id0PQ4qMdeEwjRQPrjM3sQiETfhlS7m
6NLZVtrc1d4lI9B1nQuZDDExrTLaIlMEs58PzARIltuw9LikvoiAij7eMbJoqayt
eZRE8kZ22NjGq9DvkbTVEb6lYcEewJ1RtFsUHQvGAIokGuDE8u4u8qBjjHmlW7bt
EISGqjYE0wKddj/jp3H6ZbtdZErPmXoGcQEROou6H8uM3uDU+U3rMfI4T9v8C1Vp
xACIE/AQNFgG7+b6Yhz+zwiDt0NtgWI98AW6DZNt08gJ+alPHsKlFFJ8aQXE0T03
iAr6VRM5WD4c2lhis1v/Bc6oxM1zgZKdgTl5XgDZIZUUYNx31cbAQNDQZ+BxVRf6
Gx/ULlf+Lh0pPhFMsOYEOMjuXAxJBovXNg0Hc2E7V8BpKBIQOzczr7wKtWRhLrY/
Vs+TViLF+po0adgRwS/+X4QDcDuFuJbu/U3nC5f0U+m/zkxyqPZJtpJoK7pWrZIW
DueTNQqzcWrxSBvamA90F44kvE6wamIMMo0marP4HizTZ5cVTrysXyry6usOXoY1
VXACDf833ta4PISxaNM3T+tXUduNIpW2li/oTy+btVYaVtTCnTn2nR2EHDvK2rOb
7SSWUBm87u1yycCnaMDS5x7wdm8IHmMjyuf1fW1eSCjN6bRXNQ59xpTkih/CICAH
V1G/78yYA4xvzGMcnR9zUGIu8uMk1AjYaXXQ/Btk72nEMTjWE9rx4UNynNJPeT6h
fBGD61Ok+pVZyz1xUd6FeKTfuGB0Yq+rmMaZxMaGdVDHlifANhFc6DhfZSR9uF2V
wIn71vPf5mewdfY0u6P7yWxvKsjsLh9Q2QdNCEd7IMp7TxSTzTolIT3WztCPwZi7
8f/osE0gFueMGjPsqSInphM4cgOYGf6BgBR0eJlXZx9pbr4O5cipFrqpgaftxqfX
dxWUugPGazzu+5cJudsRTiyaqdeT0+jKjAgtZXLiBgd8hJ3uqgBop+/72bsZ5lrH
us4TBSS93b6XmEqRxTRVlMFoJo3RLVT3JYCWFgBuHsaIDbM2wWEOUKUD64SO0FzN
1Mn/6POrPwe+iLiRlI8GUbSrXBkY73hMTPIO28uxg0+/OMuKN21uCLUNI6yAKTGV
rdpROWBJSIUCzUAuF2lrTYObnt2uwKL0pk6IvR91SJ2ccirB8/Ndjk3xRlGSmGbZ
BnlCazDaSgE0vJqppbkZc0GyweHDCpt4zoyrLdBR9DYiiCBDHzQctctMyt75uSCG
jDRVS0KyaEZLcGkzh63RT36U/LaCCBS3EjMvcf5jbc998fLbtYy5eTD7CGRQNzpH
PNmcO+rf6fQuzyamzhCPWoe4WA4kEQR7+WT4dmkjXmH3/Lg/jrlI4Dyi4vp7wBwy
nwprsqHUeecRi+Rw7yhpbAzOC+UAyZzcAEKAq/XpolUJA2f9cjcGOLGQHUeEaz2j
MBNpnxpJ97YzB9KTIlCQCi83aDOznG9cpQNrhEFYyKsKRnVBtpg6dfjiB8rkhDHw
go6cDcDasfo3p62pC80e5ooL3tN7XGlZI5rRsJdAbaLJ2bhi+8jgbuRlAg4boxqA
3UFJNwK46iZ/Udkw4zi0UCiDa5asq4UxwsJbNplfK8miD4yeg7Se3adcdYGVg6Mv
tGpIdDcY8xuUv4fIO2P5Me+U4k+JrOLah4efYR5ARZTFEJlA5Oy5fupud3PnNQ93
4wR7EofetDaF5Wkvqn3bDi7B3V+MzIfaigHGC/LIw4utUBo5tToJLD/HcUK+B1j/
rOcoHgWhTLyd0TWfUNVyIWZIk/ZW5GVvMCweqR3clvJ5C2Qs7exSox3MXmwQMvmh
e8WnzPueMEsCCo3p0gL7OagZyxXHL/0px+89+5W9PwXDntSKJRadjq2SBJJE0grS
tuGY6X384nn/dWRDXbaXCyUfKAS3gnjHvOwBrKaJPF0gwNyRoVaC0aoecocYlKF+
Hab2iH5LQ70hyAHNmnO6NJBrFJBiq7/sVOHK4A/NSL44a+xO1EXEdi53iMJ+DVmn
oIipgi+mrDfmqqaxQ2OfuGLmPpx/hf2tJJHnC4r7QA6oUTaZW0Cag5ozqnJ4cXaM
spazeFkKj7bR4hGjLN1t+LUnJELAKl6Y6DvHWc9z72JliPSJ60U4t1CgsmrhEh1y
YTAinYdcsbcNODJrJnHJhLlTlpw9imgTYJ1ks5+bqvM6BFDTLtsNUnIyikDa21Wc
ot5ChWAF8IxXT/k09KtNwtvIYhDKiA3aC+6iJY7Mn05Z4qx9oWlM0PJVsiRTy2ut
5wgyTUmoLojhg8fRtnjBIFNY5OgqH6su75iJNQmlagKoetmU6cq5VCk5wJqb3IGi
B2EM92GIsGFr3SyjqFyBmfpz9XyT5aTRCZrXGzpa8hor+pR9plkM9eN5M3ZQHDpI
DArh2Sv1Egr2cw93TLeux1prSo/3T/RU8SJksyke+7vMn1IpIYez2/4D8Fu+fsXn
ctNjpIPusDuE4SZ31fkm7atlLdqGVXJA/C4/BpOJnhpayPJvqeL3h7Y4FegO7kKn
WEnDUE6zK3pQ+vlUNBimZpAuHUC9DfhjIBObzQBBCDf9IEvwOTaNQMm1DxvwR2vE
ZyBSODQpMLUb6wbOcoOZZgVFTyAn5zDBObJ8a10y6raX8Y3SQKjCarutb429rSVe
w9qhamzDn8JgqMZCXlyfenClmrw65thLgITvmgitseW4bwHkQWv36tGXVWt8Rk+u
ecoaAL/Hbh9Y4IV5A7A0D0KKnowBIZa5d/89aNKIRdvFj7UmYnikFskV7RtucMzC
octTTq7TISqJi8NLYJdNZwNBhrUAb6aVvjR7jFqGQJqF9nmkR9sYnlFR3+DTeLTi
ZJ1yILwgnA31fWoeoJIo6QxZ4m9PfeGDxuhkrqNn1aozDB84MV0H/z0PzrJuoTTh
UZkvKx2rjCzavGV7iCCC4UIOThUHpqU4W/yK2ctznFLaqVtfxt30L6nqmyqzOU6l
eIkawbKmB8ov64HX/bwdRKdhdOokgBTUDudmj3BS3AONUmmAkuFVBClKEGM1Q93m
cnMeIx9j2Ii0RlV7UTy7kt3sSUDe7Oa2kSLo7qMKBT6cLqa0lmeWjML3ozVjrZ2e
kT5UjLjhZGqY6ErOZNTztQgQg35nwAZNvhSCRFhWQCBtywQfznUcZ2luco3VbW56
2t50tcU/3n+vLqBoyUjFFJE+gM5j0sCmbjn7NzHBiCg3hYgqR8EJmzszYz0lQ4+9
/nLHJZ/0sBd1+1s5WEbxQDZA//EtA8nlhdlXcez+TUd0BzSqY8SYowoI03BhbDJJ
THbLmVFlvnI2YeRgL34BXr9BEOyxFENKcBFXX+/Szy9XBm7Q/nbLOJ7RjXVcy4QA
IiQ93Yv1YH/WbrQXg3Ax+nz2inwBjZcDdvbuw7kdAYiVkOBd9C8UeNF+3IdxlEfI
UUOLMNHTDw9lMGt6ZnS5K4vEtBLcdfI55DgPxfcG162KKFk1GMo8x+bhL4hQ1kPG
zQ4MR67mhAIMPPyDOUa6EavZqj2Yi91/5zdwen5JO2mRRiGa9295TBDa9yj17hLe
7CCxIdSIdlp66f5jWdj1A41clcfuzigo2zXctorpSIqbyUTy53ZmIdifSDwbpUy4
plTDtAXQ7GgMx0ay0zdGAy+hfZ6oJqWq+PuwU4Z1LIIqXEYFE27aTwTY/62p1q/D
3VDjC5Yp7HkMIOsgKQ/1vk5RxG2e6QdKuzWep/fuED49obJBTkt5n41CtLPqGeh7
TuXg1j0mdfOa9nHoDxtQAvDN3NQAYbBAuH87GD0wNrQbXKLbUhweE+pFkChkuYel
oSt4ZqDeMMNaoQfE3nPhwhromkpACkJvPjSB2UUe8wTBu6jDYnTY6lcEotGQSimJ
Bf1SgEvY50BjXYjJxISjrzz50bgV7HbEV8OJG6uI4AvSywDbpDAHp2tiXsD/s83x
V3mOW3BzNyhM0ZOwdF41dvge+E3Ro3KUqXk7Ik7Eq67SGYgxUHukxIbMlpGI72+D
ZXc7NH71maMsCZ5+Bi858B2+yzJoQW+DP4weHzHR5244g3hlTqKJgSZeOBbniAMi
2/UCjaN0Obte7JeA2pPlbC2kUKNDdYjRSCxdscPMr+7aWPU3E5QRQLuZer3RWiwo
ORZjFMUq5QnmV6U0Sid7DtMQJIJdTZX2AemoO7BVgU7OiOyPbbEKnyg6oQ8W9Eto
KdhhWBBJpmlysGBf7wAwjr9X68VdXOXgVZ2OWFh3ikn6YKdLl4N/ydauJ6wFbUaT
TwTjtV433VuV1pYYhB9I8Jxx9eAUVm+XmehRTPcypttfRFMEuHeIBKm1Pvj2vIX2
69byCmBl4k8UPS6PHZBoHi4PG+JJDbLGdbwsqrFUr7h29ociixp09Ra+x65/MHUY
r1ltpnE3c5kaYboCNN+5IA2nwjzvh0JsO3reQcFGeGsst3ej30rNLP9/TY5bZ+h8
7IO9fo5G8fsemdEOux8P2ZP0s15UITdXuaMW3WY/hlynBQJUSdNvFRAeZ4PNd/Uh
MifB0iQsDX+kcsVqErRVX1xrWHPaKzmGKw+/tHZO0ZhOAUXHDSwmQqUkWi/1buB3
xp4J1vO6ShIiKSEj3C/XSwenfTSU9CaRZ9qYJoFr4uwFIhGvvzjeM9y0icayPk9m
f6BzcL9E0Sl7vvKIKgmmX90J7RwG8Rxg3mXtKDHJ47pGu9EiC1L4FjYUSqDE9UZB
erzQbMVLnIpKkCJVYO7OrLNKIjr9EYR8oiIb4uM6LiRI5vujIsvrkl7yjJq13I9D
aYSFMUJe3XLMJSZ3rgt6Z52/cvEuj/9kC5P4F/QXcHjU4dLA37EE1151bU6tI0DU
US73FzjSiLRDhgmRquDgqjtDu6SElKPZ2cKwzjq3oemdGjbqmIx7UEQZ+dMSUQaA
nQlRo58zp/h263XjU6JhAr4HHvRCFSMn89dS5gD3qmwewrhiGztdCUiHo5UYVjln
pZe7/eZOUPJuqgsQL2HHp9tXNbNjZ4z4BFv1XCdkRwy7AUAg0miGtgBvhGjP2lp3
4v/vLzRz3Ka8O5Cp47wG0WKHTdWKUr2DK3xsQyCPRBKX5mUgh2guWfqd/ULG385f
UXBF3pcVQ+f2iupr2NEYVFwDoZsw0XKySEMrbgdK0tZcbGMhTPYtQUTOpKz6YEm0
+G75QTXrHTYWxNxi8a4IwGC4ZB9f+7vmIofS3zC1B0m/C+yBiU+NXWX55IaY+UTo
Zn5N0MiZvGc4MjN1+tQIT6zUbBARq7JJ4+RybLemORUdq1HMSZVIuz2bK1Z6lP4N
RVR7xWty4Gq8F+Ia5QqpbvAXZ/w/3+jH/j/y6MflTYB37w187fYQ71fultlVCFO7
oi+PPFQhOUlSBnhnAGnkTwZC8f9xMtiKAVRLnOghb5rsJynLtk10GrnTCy5th3On
MhSd2wwLHVCIY0qhUqF/K5Pg+bk5Ak7bsEh3B/KAtP16d2GgmQlz6wRIh7C0lnVb
5CWkkycGhq7jp5Runw6nzySOBINnV1PLz7On50O+i7vypc6S41X8JJp5UpP6MHNw
jQGGLjd8/El74uSE0dGKbyQnKVCK8hYC/75E+ien0/6uplgYE+b0/wjIWCMv/Nlq
tW62kXhgLORnlisLY7Zznr/P6ZoKXYLUb36bjXpplZNKQdG2sWp6J+34HNkqhgso
pubNDDb8HVAMo2JYFcJmRudeJPPzChJYuzlQVZRB/HfMzyTGb5yub3zC9ZeISVat
Ri5ji0YsCWnnWgMDLIKKJQxJFaphE/pix+q8gBJIrl5SOoRcdRlMlZjYIdJduAH+
DURLgbfkLOkUFIK7BJA7eJBdpUU2cIOopK6nYne/neWIKHSRTOeXsebOEJpcO5xX
tA5g/7AoUr3LcU/9j4Jsajl+nu6qziPfj+WShVBwDLX9chLRQHOHfRaTdWBa1Xy3
Q+6VaK/90/sUIPiDu68q71hFxyhpyTAuPFByymFdn70HyEQek+p2MmIX3PewOnQT
Ogo3N1YhCC/a4aqyUsCB66BvGQcRNCViM51GCsjiCAKoJoyRkq02Sa03SpFVJ3f3
byw3/WGGtTVByHvNybzaed4ijvpnn5xiXUeRaurOMn+9fVAtN2HWzkSoaf6ef9XT
cLn03LPRADUsLeHjcnkWT6PPsh7Ho98Q6Y09JRqJ1wQVba+25UjGHJZkP5m7K7Tg
Bd2jqPxwj3XOQTzc2SC6RycmCtOAqGR/1aiLGis4MOhtrUjb9IyCydzNvTRra5Jt
Fjl7CsnsIdUq2D0kWnO7Rs+GnaBVna48luqtKobsFCev3So5crtyN9KMxqrdiNJ/
o5qGqq2LJog3L8ffq4Z1L+qbNz7r08J30skwk3BbyWUrgtJnbBdJ3wpInMV2eQ8F
livMNY84yIetN/S4e8JMZi4W3N+kN+9j4BNQMVvT9eIUVrQt/w0WbPiyF7Qz3GjH
wLQOvIFkvPdRXcnFmuCUwO8uWq+hd9DACv8jJm3nXxv+aRq67+xSirE4Il0/V5XC
MJnz+gbV7uDFDyYmq8QcVZD8seaavR4motbpAjaT8f4ZDmaBVylF33hKqPhOef3l
lXF3l95BHvPYFEczhUY+hz8rM8K0PG0F87548vFs3poPOBAke8hP9kGdd+u3YURZ
xgia2z4JfE+dA/URMIFGh2fa4wps/5rf6P1jtUFnCjZPzwz4b2TH5Db32YaVuio2
prnTReXetxOdck/KXtJbiX4A3AKnGgSvom6XrTplqxA5Lus5K2umJbXC8TKqLKhD
80xfSaWY9TAp0SSJ1d1dl76b7j+FOAZPSD3KbLXhIOyLWoIkBeZ2kOq7Af06OHVz
B0jwaNFq6AcgTj3tFFbZwnSPvo32l+PWqWZJaC/c5gB66hczeXyNAn6JTLVBVlt/
JhtysQtj7P+YEFXddKvSL+ClFDw/EUJ8hl3T5KaInzkM2Ieaa6pNVrBmY0hGqTzL
sU7nFgureTNrjLWp0XAHeKHJy+Q+d+oJ9L6QZA1NQExb5JAZrczzb7nzWWuZZ/QT
SoSaU7L1HGdjweuDh9lo65QC91Ftlg2WcksPd36fYEgkFDI5v0ottaol5Pa7s3s0
bWbk86WhWGa3gbO+PETO3C0GswPIcpfT9cpxTQDiyp9Nv+vCx0vjQ53gr25y8vaQ
JAKFHGT2UzlElMLiYAM3uG1YiZJKkys2MRpHWh9760foZZfy39MYeC74IShd+1gW
hBdy2QWJIUtfEI6xXCdxLmwGBpz/v8koniFoh94+4NXJ+lXoDhoDn2ISKBTVEaNP
PmCxc7O3gIWoXhSNNzwUD/vnl7IkfReBvY3o//OIXA6tUrtDEeOj3QJ4qGcIDnHJ
BSbqjrxPfKD1zgTbehnISsvveZYzUKvVDJ9uVFmtao1NVqfiYnuwfOtJBOttn989
sr7Wi/5r5q6sjkzpP/YkZAlZ5DOO5/35n/jlifUGsIh8/xWnENMNTnd1IS6eH6Sy
0jjicnidgtYx3m31bXXYF7+Yj+bH1Wz/FMj9R7eM67j6kHSuik96820nQ3/daboj
LoPWvOrsYxkoXq1s1pREEYg8Pmkv9pEjW96P0abkj4jSL4GXpidU8nqXZM8Bqyev
cgGLHLTutTF0k4Jorma0llNUen7y3R/NFSzBU+uqssKKOdQR2NWu4sgY4G26DQVR
pcirVfMiEv5vNPgM27ZwQPTCgYXnVfigubclQP0D2hgRW9HOdWNwrcsRIBbitty3
sqVDOnpFoqOExncqEA9WzCChwRkYlDkT66adwCULWHSDcM49qpbdHvHYa4uMaX8M
AzSl8Dzq4HYryyQu4jPCLlgiMiVlkaIENRIeGzww9iXLNuanGGMJsFh5Lb2qEHT7
J7Anqx3yJ7es7rxqFsYJae7Xx4wRiACZuOnzGthbToGc2BqHEro+QbARcGObTAoT
oMFIGl6CdOgGuHw/HPU13gQY9l+0WgBIFRZnsbBHzcskMGiExLi+nYO09IPPXK62
kFI0azifPDMGm30qw6gWRhE2esw0e4J5eUVDB7ThtdWV7EFmuBo3lYx2VrhA2Da/
X2kz5ObOcANuH/3P2g2VkgB3V2vNLWu8g33ekHhIr/YuqGTeyjk0IFFRkUvZ+9B0
hq/lEA9hoaI6Pj0jsRU3ZgyePaIplxQEP8/f0T4DtDfZA0Yupt697t3VebYVB2vX
dfXYxdcp0EDqDukIkzv79eA3pr0rZ47iQiDgBW0VwD/kt4idIPtYtI1bIOhRMS96
yaoEVID7c1dtVeOyjii6u/t8f2QDSPgiwUXahqjNWHD+c+3bi8yjGYWdygqpVRUZ
U6gdNTaCGL8Qpfn5BOnAOnhApzYmSbN/CvDT5I7Khade+EbjCNCIixC0c9xFaa+t
al1GHlloKoo8RPq5A8ZbzBihorUltzqr1v6vKiB5IypecJHQbzmCGDSM4WjQp1gf
o4dBaN/a0zfXuwkoUXJ296cBcXDPxDwZVvUYXmgnviD84oeoTVNC2x3EkiAIkaU/
xemaqQtBQExKmeqPUE/iGHaxUoUg/gA9l3yhxM8CS2bn+JX1sjkB1PoylKOSw5Q4
ZD1tCE19WBPSizzRQYGLb693IV5mGgZIA02u9wvuboj8iUcMfrE6J3NwK/WV7mKs
vu8GMS46z554HT9ddPcWgeqD1mXFpgScwTAAJn0GEIK7OjOZaM54aKSoy/BUT9ty
YWHxqnudry0yTM0bwZdfGXzW872weok01wjIeSwNPsMjzDHf4v4/DbQJ05pDet6F
b0hn39Zc+MOHrH8yoFYrWX5Fgp2vUs/FHycG3yLOEseKBaR68Q9KOkardycFF7uU
Tj87wqz+UFeviZt5E02SoIHLJa2L/V+CQiuHspCnm6QBXk/YMIq58WFKjo+Bp/i/
8Fw4ZL4kZTmOPouM7dN/+856xt5VHQis0won542n23q+pRhTC5Q3sgOIqwGbEhh6
Lc7KEgW7KyYJhecFrwyeQUBMr6Qns/tIlT98kyjCqJFPIzKoX41nC8q/o+FXLoYP
CQ777RLNp9KiZccko6VMIDKLyNJ3e1qP9WgUvdUZJGe2AsqUJscT+HYxNCrVt5yR
8td32iJFOKhOjHQ6VciEfU89O034Xsy1zs1BmVJ6/oXsQlxgVO43fWAs2WAUpiyE
4bXx/PTPGP5fgeCkj6cJAL2yvjfiMVCducdSUJY+wpJ/o8jhuQKFssM2lM3dsTTT
hIUJnOoxxQvukOU9gRrvGB9BwdCa05N/KAN99EabPNsnK+e2CzPfKzlk4PXdOpIF
iL1fAfHzmoSpYECNZatePUkchN+pjdsvFQJDvqBWY8M9LhnTRhoh7ourjidGFRpZ
DLIa7q538l9pcbVe63TK/52e6WR2l0gqGdHZuSZ99X/9Ph5iXiVYnnzy9ibKH89p
fipXarhderC9CaFmmBrtXZZiVpJVsci83kzug+DpH6EAineGr8tTUncd06RgjB6y
ulkjfpkkaa7sps3E0wQ+0ttByVvWCazoBU1bH6ZtTCALtNesH54csr6k0/vL6sR4
HMlyumX3UbaX0cBdgiYn/2HEFtMjYpU77RqHFkG3N9lZ5T33Cz1J5pjGVAmeFmG4
UA9VFHatCJbVbK+apFaMlsKM8pbV+Mjcj8KHjqxdnDPi4FvQ0j3Lo5XitJyUMYyZ
9LQqZfWh/eR8o5kN0FtAFzijCfGWV7OC4yo4yubPweJRI7DuaqSwMxtCcWB80DOc
mAvbYjAtTYwrBsUdQ+mMISgNdKvjAgbKZKem3EDK0dn0Zf17DkTOsFVvCfNj39Sc
GOUbLqyi7fChTeGTvolWMnnAaOEisVhG6Gp1tFHUtRceYby85T7ji0PhaMSXXXbL
fOdV8iLPyLb3p7xp16XQbnjAMySgJPbzAR6h5b9JT5BY5ln5p7Wt7JRYUXslSvne
5VUWMqruKRj9ZixtsixyQdppoRePOhxrx9kQCCy30K+NLIL4YDsOK5zT4ewjgC7D
tt/+/ZR1+hv6pg1SI/BNQQtPUlOy9WSA1fkbd4gVLoqIFsWOtCkL6xqhdGAaORcx
qKKqCp7S1EbNlO88UsXO9ZU2C4BE4t8TvKioswC+FjeObwRIfcAMH4nNWjHNN2Ox
yIUhNb5GXK9ToDVPR3IiWs1F4YoY5hEQKc+eaQN1LgwN653Lx3a8IYHUwWf2Tqfx
NRMCx4APwFEHwOtQHzbFx8V0PWdKBaCkR8JgVPTNRNJq4Win7x5EbhRStDEb3vio
oxwSKlyNszfjBJT+17Q9Z+g4xy7QsDI+66Z7k4ErYPJrnnJoqSM5at0sfCpTNwLf
8Fdv1aDOgaDu46kP8JQcmqFpm9FmrxsaFQZBo8t369tA4eplzQO+FTLtK8gp4p82
ovNlYZ2/ENkUo/M3F6jo+pSAYmHiU1Bjnj8ZjFsPmdbufx+NmPp5VdjqUGdxqgnU
3GXaZsAqZs7clnnS8GFwx3YvLqhZqi/BL9ytFjoPcaXzCBz1wukCnu+bZcJVRZfz
ISZQ8JdL93+7NqJtAMToTryMsrpCT/fUYVOUcfotnPbq0bhigI8KZgZEPt8iVq0u
l74rZB5bLxTdMnflT3siqgjsCRys9mZDEF67Pmfcd3z0Lb8I/Uw5wl1WJN7b8E08
zPfIXZCLAzGxKU25vM+5wx6fsxaMp2PmJ29ndTsTCH7JsvZ4jh3k4pwT5v2EacYO
M6N+F+QaWJa38iyVksGtkxiTE0mschHxC43Ly00TneccJQfEUW0PV/+HXp/C/gDV
hquNPabhibu2b+mKR6ZWW7PBSvD+Lq68pklLvKJUWMrzQgHckh8LTXzu9nPQyBKL
Gz0rQnNz3+TbH/eedK3THfRdQ4Ryhvc/c2KW4hW08L0gtOcn83e2R1ECaFp9qOU6
/rgu1dHLQ8dxrtdLPpzDX2kENI3gAbHRG8dpzy3B9YQ659YIhSwnq1BaVN2NLvBS
LgTg3VtPK3G3+nLoiFGgAbdbcH+dkbxFDr8cH9C6nrz8AXUtzVmsBDSvMomp1o3I
OlXYRepAUfevvL3sNoa3kCVVZepqFQvYFcfnI2NAHX/l3JRb3Y3RYNNtM9wFEN08
iFXa6lm/fXrPMnnMo777mEqrSM/2OnEs4PHDaG2uJ/j9OBYsSMyf5US9lcEiZz4p
0ngIhdNk9Rotmz9Zw5Ln90j10QNrUPNYfbJymyTJLim2ZyzTS0GUh2lZ/qiLHLzn
Pc3ezpE2p/Ts+r6rWsC1+fWo1UvYLIA4boCHf5lnNr4pmaMHa/XlZ9EU//3Qozjq
lLQ2ubPXemT/Pzna2gNFEI+0MokJCzbDI6P470YnkxW7aURttG72boY7B9rEppQz
gt3r3YF9e9dYSFCa9pj0KFdgElrrchg5Zlf3SfyfSvSwoH6I9Jb6y1DLA3kgJJX2
QFC8el+TcFNfOyHglN7SDRncaaedHMYmNjZNtPkcq74arsDOZO1erjh/KXJwZ+OA
8qpn1yaCVUWcORrdC0WrkZojMd+YV2JJEjwDSHOgnaG86ldLlz5wyJ8p8rbkXBX+
mLatiS1RIbVS1foIrVe5gfV7Zlc152Ojjai81aGYTtt1fC9xUXaju0e6576FQkjF
Ize6kZsG84ZLjt7FeVakbZU5fnoYC5TtArDcVc1DghNCf+SDfLiRKKQBRPmqhWpm
K9Ex5HPXrXo77cyy7QwthKOltgU8Q2rfh4nivTCddC0di5hfGr3PHZi3tas+2AAA
mNmEGiGqeC3LbqJPAEow290f6yRuf3VtPC5Q5FAqfJpt5GdMJjK5IN7Buzz9olk7
x36f3K3ZOuG3PThpxaS+hZR5qlrzO3Mps1HD7gaHabWfsAA6IsdyX1ypJaTkyMRC
xKkxeMTx/NQwHBg4fNwiXxabZtzkWdnl8y17rKHl2gFUIfyhbV1jjx/1sL40AfVu
jalYL0jTFW+0UoAx+S5pmexCYFCpAyjWi/uvga4XaHLnprjgh+41c0TC0+UpXCtn
YuMt9Pb0Bd5ENzH17n/59vozq1lJpp7Ft6nfcEXTqhGjkoV0GLtJ1i5u0tB49f4F
4k7q4QVATtmq040CzNkLaV9yGIlLlcSrhdFWI6aoaNUVyjOSELGGNIvxRuwUglw1
mr2uij3B+XIM7IEPPUw32rOljQQGzbwSlPl6ATWK9qjq6/3WHA+axtUD28hhiJAa
SzQ0D+jDapVHEK/RFIkBNvwmQu9Y2DQWaY40xFVsPE7SZ1GlHL/jXFU9BlzmKHGi
Fz/a4Gkhq6SAaSBKb0Dpq27n5rispwLhUezbSyDxtBp2XGtZ9fR3xZwzpTnS5gS5
EFzTFi45RU5tEOupXG9XcJL7nBBEKPQtBriAtUjhfEefV/1nhQ6FoiIrphuypTgB
T19yjefnZOkZdJgTVzXH+YSh2Bgu5Z4TlaQ5xRWEkrkijwp3IXQFQb10/fXl8SP4
gx5+1MliYgKDp7wbSuu+j8sRdLg7rILhMfBph9rgVxZ8wMDzsBVyxJKlDAVgg12Q
wR57K9Ago91vgt+pZBG9g49kW2UsJaDXN4iBOibRNCWI2Tw+74mfmxUAgzJyMKiJ
nSDiXF3ZCn34oFRCetNaOrTDIJJG6oTKIthqYHxAQwSge7Eq1DreVJiobhQJnUZw
37TFFiG+Id1QYhAFsQg/lTY7yuPMROgCMvU1t29Di8cg8T3dHag+OuylXnBL1vyR
QzMBqeT4rtNBhLhhTToVrx/Au44fV01q3T4JOzCLax30W5kNZm7eEOEAnnhjwRur
jDtQ67mF2nsqavNJeG7ZCcs8kfAO9uzG+mPdBju+x1SUiUkVJLRMPWQIVUXuB4RK
DnnL1dIg9vcrONLAEVNjy8iSMHDZASd+OxIEgUd8UX3RSOWHDxoSuHAlqk9CoeXa
LlzVtNXIUmbR/qEOy892U5V8YKfPfVmjvfDmmQ5cjXAjX+xxSQZ44FxiQlmEtN4d
HwgFh8/5Y4iJkZNu+AxzkxSiaEW9Icqnz6ecAyHqBEdmBQ8sU6OnPi9iOXAHwH6t
3WCxVF8xBeRrAQ3kiE8RAZIb9D8ueCoCnv+7jMHL7aDhR36qcfQGdanUHihs9t2y
Gu5G88qRCv1t0y/jhuaut5IGO8c0iIeKE2IPflwRm++dKBsDKHr9fzMvdTcDJajt
bAHHYChJs8nVi1xYqlNYiz6XZuuCdgs01arscyh2VNf3UOisKV31k8kgPwVaav4f
k16xJF/7DoZ7Rz4Eckhec56I+rTmZ5+qtUu4vBF7EG9mvxwD4YfYLK49h3IkIqT8
ol9vtUVHObDWpofJmJXV4wgzlsa+4PVOTEPVi91HeIYBq8yJD/lhXzzKZR4dwi50
jogx6fXvVWj1jEczWSdD4qmOH6uRY8sEX6VLqx7Uq6Tlm7R/VNGhhbjPW5Y0as5t
dgIsIZGQejY6tawIqdSWeTwJyC2YXh73C9h64wxGdawQVHX7R3YybProdrr3g/Fm
iNY5S2RSry3F/h9aS0uaim5zadkEcM1bW/rQFKOw+R2XfNUQEvVioo80ZUUgg8a8
FsMhd2P7Vo9lSlCPtVq2ZEICv2zRreZK/gPSB+drqX0D7XGPha5k96joCIn6nfv8
oxIf53yKYEEw3SQCkPz/1rOfKToOZ+vaOqeDrezcuBpohKT1uLMF8zaEhIOUYVm3
e6pNPPIFHncmByGyZSwmb/knob5EtH166lN88f1Mgw1NxWlM5AbEEwDBEw3eI+9A
ItCN6JCAWX1G/eGxT5gvISuzezlXnN7A6Ux+etcLdOnjk9cK1Ce/3ZoV6XhRSXwH
A98jmxDOhFUOsqqplrhfnnn8+MEdW4IuxLym6rbeGarYeui/m2QY8kEDtwe6852g
Qi2BL2SVPQZD6SWKXq1p20le1jjplmSjnr9tI1hjzHqmvRPxeQgvExkmmTXXaZCE
1rbeu/seQr34+ThbM62y4NNASTjrr3lWZrAaz2arVDsCrhpxjnYCMOnjBZ6HFiZi
S0KTXIBBtydy+Jj6flrZ4dPBAmoPMR4PMQddNeulqRmvyZb0Y8cGJ9IHQSHehcW9
9gPY4g2/eJG8YNONFGErHztxhd54llaQHJN8CPrsDWnDke3yZFMM+22sXUne+I5d
y3Qle2Td9OCxJM51hQq4XWo37SbdImapMonI0FDOOPV5bs/RW2cJulQqiXB7vOPF
GJ4WOUp7e2m1/fzMtvKev/dE5WeCpFLZo2xEY3yJu1xK7KeR8KSNgY/veV48My9/
Ge5yzdcTx5cZmupM03tcreYrekJNQh59K1B9vyczj20uWyH0w7E1zz0QuYSw+lsB
rp7YlYKCv6wOpLQsBD4OGUnL0B8wHwd0N+JWnE/cuvhdk2GKh5Acz+fQaXlmPpcs
/0diZ5FEANCZndalpZJu/uNAHat+wvsBVq0WyhSlJdRa9NzETPIHvKGRJ4eGGggV
exVu3r4tq5MT5fWtKcMEMxRG5WMDtiUFx+hM4V3E7Oet4bxdproPRSmgrArdBmlR
gu3+vOQ4IayDrpX5WRJDwGYOaWm3En+LPkFKP/4AcSLECS/fup1+UxqN9dEpVRag
grfvEvNo0Mf6xQjR6eKW4MaGjGCiNsY6mL+IAAFxOA/xFQw7p3jyodV6tl/ZGy6D
MihHJ7d+09Py8J/SnNtASGbEcc8F6lnPVPoiDK9QrajMm5APB3Z5zaStMD9DDUTB
KUg3EdlLzUQtvav4mYGHcN+OV6FoR8YaTjZMgkFS5OOhfEzt3t04tvAzflcu0MhN
9G3BTcwrtOXVtyqT4ew/JWZhg7Ll/mtChJxHfQoDqNLgnJYymHWe5bInhlResBUl
KtF/ajRf3CPx+wr3HyiJUiYkBpBg568uBU4YI1uhjarFX8HYUd15voXri07NBKso
M4XHva0wC/RH5ap0qpUuGZTw3O/BR5OwUbl4Px3WlvPSkHke3pzu5BqNPrryVgiK
K+L0d5Q2ZRWTi7ZrWvjmiRlPT3PE/Vn0YqKc4DBrYt2mwFCTr8Jkl5M6z0OqbYEX
aw/IvAV1Fi0aq7Dur7zElvEVgGVaf+CEBluyf2CJw99lTjKyG6VnskxrLbj8UKd1
I0RoGzihJ4kgMuai6KH4zXLsQ5mzNVAS6Y9aBz8K+Gy1O/MbludxOjfW73ipDLjT
xjcn4QwACSOLv/WDm7latQdTopb0mLWOpzdaEGa8KS/87Wd2u3l0z0c08/iv2jo0
/TpUNzkTuuNINAbuOHfJQDQyBRgyl6klpPnoAVaphALZdDx92eDWv19eHvdSgM6P
29kUX0M9G3+8BGwZlp2ZrgFgZKn6txqWu4TGRI5vbM16b28sgEktD0Rm7Gh9bDRA
JP1CpedLcMUwsWGwErEkMNhdvGHzHUdAQ2PrsKJE14i/KDg2/dnTdpKfWVSYKv5f
JWmouciurYBeC/NVFUWC4XhUWfj+c4pWndfRX64Dv8L6dzONrh0wVtvaipTmBqFz
YFblU83Z9SEZxHYqt50SLDltnbUQTJR/klvSIiEDE9CYU9d/tGf98RS/RN+V8iuj
a240AMUyAMWesTpXqivzv2CnkhLqVTeYINFfEQ5TqLpqQeTy7CB/3Hx3qlyLlNS2
lE+blRNb28D7aSEUdSk9qFgY7ZOz783p4rul8Ub54HPxkQ6AA2f6ygBrMdpuKs0/
UHe+aCH2RrpeKKoNxVT4ztYhB8DbNPDOHClEmVil5oTTyNOr/nHV0qsbueDU/baC
HeWeFqaCJ5SKrADHam+f8PyS1yC9VOgOM16KeKa7uim2pvjLZQ3aBIilq9rBaGqz
hK1XArSnyByrkCX+xB+vuO2HoHzeF1DbP8ujNAztSWNdF470wbyLr42seRp7/ZoI
+BGUIEqVO07nioObrGZ5wEgAzEeSq0Ien9Jr93ih3KGF3nOraakJCTGsjG2p8zlu
mgnxafyvhMp7M3J7rzrtg1i9RxqQRaSNsNxtt7BPlgFvwesM8mZKHxQnpokDvuxD
5pBsTCZrNC+pfBJTKAx5ZsZCb22hAisEunME765tYPj9GC+lJe834++C2U3tg8Oz
idrcKhhoMC5yzFs4dl0A9nwkMq+zyuSi9PheHUqmVUV4tDxDbHFqfpRoQ0ZsyBCi
iOBhVuy1ekBLz1bv3SaEba/juO4xx+kC+mxAGNuYa3kBHo7DB8MZHrgEtLx6bCYf
lVbXD4YJhqCxO8PnSLhXawqOoKTTz+8QMO6qqjw/ExjkR6Tox/5e+y7rVjc/qhpt
22vR57efGPTe7zL2nLZR4gPfVkqJKWcD8Eo0p1wpiGlYchJF7ZlIusYC5PpTgA+S
YOeTN9VjHgDG5ie9XZJsmEm1Dw+llrwLN1mkC5tcVArrsMBXMWzc8WUshBjQkSaK
VvOULD/KblV0tMSylfNDvcf7H8NuPUx+42nGd1OpZ6qnAVmSjA3TBsN0CcbJqNPj
Zut9vZsjTRAdOqe6dO8keZ379bcJ69DWDVV5zVvuKXbNRCbSAjx94i8/xIyUWFGf
8lFLUfCsxlgXN3gA1hP8SgygLYdnAbXmhysZLZZtBWuo8aZcNIxLHQmyjskRN4ao
O+Rs6b7oW8/EBFiwoG+D5M0YFMURjSSr8ZX0HjBIx8dWxmYeXG28vDFOdcCmr3+K
ULP8F2Ifw81c5/RwJbpVcS8uPLo1UDm1ldiRzYYUz33YSvlhD+7RF6dMrCiGQqcy
oFD5gvVwUbpdIyFNhiK7qXOVyrSYaErjC9S4Ntf57FXuzh9nWCbgWUaCBMkgp9OD
uAv9SpNpmiEYJYpGuezvqJt4YzlpS2reCdLFGDfAJsQEMHXC7bOcE6a85+lbkYCE
9kmQIZGfQXrbHyzXcDgyipP4qf5sXCQ2ubuJh0GG7NriBGjICIZhCUZTPwWW7B93
GBH+FHo3aS4kruOlQ9XKJNHgdNl/qaBXRXd7UWBN3Ofo0+bHJuGoTMrnOudTQmZI
YBSN+E6qevytV6sv0ciQx17FAKwTMm82O3ZTtqWnOQCBcdgWMs2GSAzzUx4AkGle
m4IuAa6kcoiayzOH/z3JovBD9laOSZNdXE+42WSEaTKzZGRaBEzHT27+c5pSAmbB
Dz7D/ntGnFjO6LD6Ob0a6wvNO62naJnzherT8Pxw75d9424bAe0brj1oHodJFiIc
95vZwUw53F3SkE7yODNF3LHVO2bOtMj6lJN97GS2+sA/bdcH8VmNWvEwhuZ7AOPb
IEOC8w7wIQf7K8dZp93RBcQo1DzaBmr1XOxdkEKIU3z+q7z1WNaIaghqDYidB6wa
MscCX8I9+6uVqEcA0hqYamU7RmyehqxfdSZOEzzsC1Od70gk/FNd8Qp+/zahfrGz
Xs9quLfEOaL1wEAqNk5Cz2TRCJhKWPptOTTezFO7tpbC03YzQR12KcXPIWLZ1DAL
SJognIX9b4PITekYa7kKNJEW+6i3gpx17N22qAp7RW5Xs9qHGUO/MmqhDxtehPuz
wFXwXIeZfI1w7f4o4VHBO/P3qBdyuSWasu+3HecYTYBhqSePJx7Thy4r0RVsAfeH
6Zxm6CfBkZpWlbBo8SMvGfHpVQTtFWrDkCHDo27/kodWlZ42b9k218+TQ6HYmcxh
rUIbIqmVE3m/O4vvzlRt0ztY0jlGpPZnuYq4Qik/l3MqgtdPHTRnHL5tLZpQAEIR
Uacx7ATWfhWMjgR0MtfyYFouC74VQxh/grr9CPwrBsdAHrqOr60Ikd1d2zcEKa10
Mn1ogZBVGok8kzIPnB/rNXTihVrpm6DWvPiV6ezpe8um5A3GBgafHomsL5KVMBif
XaJv5EWwzYbmedizf1JgxO7RMhswD1uHIugg0vGpbWfoxzHsRJweoG0w4EO3oPzs
c+gWf8w2+JPtzz+xK+omJ9Kb/e6kovDocxVPNFqBXnTTk9OZ92vl3ecFiaDszMN0
z6QAzsv4V0u++GHQTjaeMn+FC+jaLzLLviugLWgOlFrq/XdMo2ck7xE3eogzSQ0a
dbTvKW5jJ3UsU9auBOxg5TFNosWSdQTIEM7/teILStGSL4uOFnIffsYKM2J0tP1A
47OXgzakZEOiJ/DLtfRcqrZYVQvET6H1GFqbh6deg+Je4JnZAYqQUtuXG8OfEIMw
qH5wVw/T4n5HJcF+df7CxsKsn94VRbNhEm3G5K8klFUCa5KoqrJ+QVSmNkIOQ/L0
mW4ziKo0PbRc1TQlHiCK4sC8tOHKrGoZ+CsKSmgI6SvPgzp+zEnWgDNFRLIWxaiq
hrJ0N0CB2It8w01X32N0WqzyuOH3UxlIwe1O1Lifo54mJV9rb1aHjba3quGSBEDs
zVhenwLcYeZsdue8rOJmXNsQdXoYOtKgnR8G235BC7qFumcZ0lOyLVxDOq0Nx8MD
ywkr+wcsfUyDbaA3++TsIoqQoIqpBX4k5BiQbeIgZu5XZ2zvpiVweDQdM8XneQ/n
xhCgCHdogDya4hXMtsBM92AcNOYnuzFoPfU0B3fgWSrF27DItyjccNOn+e8fzfgw
FqDp4RHvC1PIUaBF/vqBODbNYZpo0S8/mspdIVtwRHhGBXnStrHK0/nNT5MV+/eO
w9Gb96Qumf69UXaUbXglhJ4AqAcMb78XWmRXttXRFF9Bx0EY8Jatbx/TvzeM9HZB
pTRn4x1C8Hf1exoA4SUTPQ0svCAtrQ8I47ENzHuWoWhCm1Gr8V11WQtjRT4QmFI9
qD5TToeigCMPbFs22C+s0U1OLv3F/RKwZP3FRYZHEXVhDeKA8HUDAxx/syQsOTll
G8gWWc65DOlV8O5stYAZq1cKEVZzRfHZdw++PHv0BaC2Qr0S5XBD4dNpFbeiAv7P
Metx3++rwi9av2dbuKOILSjeDPyfa+ZiGsFHVR85xFj4X5FNg2YqeWMkcf59qKxH
TJ0X1FsO8ZvrCziGkrqEsDVTWlldP1uAj0eDUIzpVggUHgFhoswZkKWM59oR7vM0
J3O7apWYR7s70IgS7L5FywQKFf/alwIpnaKBWBlFzxkjOrElCEexg3/zrNN866LA
IsCiKBFMKEycailINqyrP4VrHdtM3v+Elf5SV2wvBJfk2U59LbeDO288/bWukpnA
CF+bGZki+lFpid15Q8DSOSB2Ix0UtEKGAz5IOcog/YnX9ol3bOEvDFA+zqDv1Xw/
gzWzaLL4nGO1KK/AWjd4qr0UPNmEGIz7IyTeDQCC7uxfBu6QU+WiGlKXZct1qob1
oP5X8OZd4JZMVRfXAAG9hnUE5SxaUh6hRQWRFjRr/jU4k41aE9h+SzS3WplVLL2Z
4M9h9vIkB5woOgNdGIVjmyXtZ3ZaIHtl7DD1LDRRLYbnadHp/B8Xeel6U+4a0OzO
3FLXi3zQZYftdUuad2ZjGjG7nBPVWB+S6/5dXw/N6HL9t3LFq7n701GUELC/hzma
a/fRgHI6j/3BUi7vqQETsaZxzBaXLE3PWlSmPBQwEy5HgiBNd3sb3UvNJeuw7HSd
UekkbGEnbBHpV+CfvDmoSsCrSycgYymMWYYgwkkkcMtVsmPcOOitGZ6jiqOP1p3k
TmFydf7ykOiHllyPqUmVa4M+gLfcCjTRJBYA3yitWcHwpm3Z7DM/AGDxLkTR6w2X
HMoCofg0izwP9n1gbP6bSY8Jo7sId0KMi9g9IPSPG3NPku2IpzkhWzMiU/3bhBzj
7ksk8CYb7kw0U3OIN/H6eFGSMx6mDyoP4y26cpvvDX6ZV6uLgSBMT6mjowC/HH/6
4dOF+Ee6OJ7S/UXrW78q7OrvhL7UZ6YAm3eHnbA3hpGqjQ4+viBF7DHSaVCivfJp
N57GLcofTt2SMCejzSTE1FVWj7diHIY3W5UAoDrQZ1V+INvmtN6YhbTS9dGsUKKU
ne2pMQinS6nFXlNKn6NfW7VrplHbO6SV+2fDDmVUxGuaUjvdJUjRGq1Xm749bdMT
Ms2ZxlXGDtWhX4R2IpkTAgYI3dKNB2qXSgDHMgmjUPo1k0GrYc0WZleVWTFbyc07
KzFl8n/uHNv+nGzvUzmost2gNCNdAEwXSRi2C6I56RyMHpnkwBOztYsI0UPTyUvV
Zi3r+cjBnjqwBK+dXV+ksFWt1UTdR6H7168IIxZxJ4gkO205JVdwyxPeitzvJMOc
9xJrWiFPEHy9z4bk7fxxqw7tLtHALO8yg/g7rf/PjpmozD0PEjbHTNwK90YUoPM3
vgZyqOMDkLnbDUrLlkdhPU5gXtHEq5xjnu8luTnEDz6Bp0IjMslj+JahcuwCYNIY
/nj+TEAeonDJUFo2tJRtnhOUY6UdaJ/19MuCN5VmCOBGJ/QNv2Fm0LLC1rtENGiu
6eAXtxIbOk4cbybQgn0ITgtuhHO3NLGHb97F/Yy1x1Mn3hzO6EtDdapLcH8LW6uK
mV7b9FBq6uASFYi8mTmu2+HhqyZEX3ZstRKCh7yEht9uvALMjHuvOqLKtxjNDoXQ
Gbm76A+gWOMDbYVijIRq8QxNHLTqG+Ahc1rVPIRIdeIXEob+eInjDRxsyp5ZToW/
FkKeOAq+YZmRLO/HnPoewpBiVRT23KSEpkbAmHHKEAJ+VtIX2ssV50ssUFGmh18j
VIL5xVwA+1F4JuI+DzuUjPf8psWz0UOk7Ns6v+Oc/k9yY5Zqiumsmy4h3FnIOElJ
6h5akFeswJf0QXH/uylfQnCNAwi3bsQ/11ea3peWvWPHwMX9j5feyIZeABXp18JY
p+1t4ZR1D5Ct/FUZEGVf81PSPySlQ0MiGKbdECbGsMbTDrGYQ/X1CiUUFgid3Lri
VUD4fs6n1cNm0KzTtCWzDI/bmK2JxlhsQR2GXUNP6eIgtvxth1AqHAYFZoCKC9xt
X8sUOtC7o69KWVokMar6qta6eT0KKfHbVkodmD1HWzOWSxkfMjzlsAJM3HDeSt6v
oeuz3xDPhe+LRRqheX5bRbQOYaB/LllA5I2qi2MCth0OfmCslIpT5gwaibOVuCmb
dnLRcHMfPAq02rvRPsl0qTFjV0x9p4oUMdrdJibvPvH0epKbrLkZGv7OGiBg37gp
t0oa3vdDgkfVhCAz79Az1hKgjTyrNjyk+13WT73gz061jILXhvDOb+uhlZMZXQbr
k3CiL60ZratN/r7B346QVqLJcXTGTiT4zfYIIZZiKxNHXz/lbElVSbkiyJ88exd8
AoRc2PnLAk42vBIgJVHSwC/PCZWN6Dx0bu+llxmwMXaxIyVs4AlklFZG7TB9gxNx
1mcVfSNwJ+C2bKF2DSKUleCtFVGaklUnsGz0RzaYlLqiuQUbCr/hIaLw95roYsna
Hc6c8JRO+0oF2AfEexmF7ilVTcfnXtFQCtBn7OoPWrTYiBpOZ+Hnwg9eVJlQTGYA
bG0sySHYZYC0/OdXeJg/U/TbIHrnJWnwCX/V6zEhE+Nrd1WbErqqulAJg8XtErCj
RVa+SRqOKtpNzYPk8GOO2/dYnk17QlX3qKbmvTD/wUJecZvzMtXlg7NNbfpzwdyZ
iuRIhDnIYceDTtsx/xL9txnz6dVwB1JE11s4EP/8Jz9HVEEM+20GlO+iDJUAY4ye
5ydej7yJBfF7+VgE8pGbbDecLrtW7xeLQ3bJgcp+PF/3MWnUHW+hp2OYUtHnX2iQ
Wb9RpT2m4B1baYZGgjWmvz3979NtKB/0jfH5nxrQ88GXtkYwax/JqxbXypVf5dIx
JiRRWfLJrY1Ea4nZ59mtbmUegUrJiqQwthlGHujNGyURX1zJEINxDJxkJbDnbqX2
5FEYOTmVnzpmoUe3kk2ouY2Wt7EURpYlVHIx8rosvNikh76j804xTT5Esxoh/WXf
HjnuOWkWXAh2d/huquVHkF8XjAsevBixIjkCoKO3DMIwRJdIoxn9Duue28rWmELL
DmM+ekI5qIY2oFAE6ZPWaIGAkpe78Mz4KIG7xFzgm3z6CLR6t8OohPWfRRc3sDoW
B9Q/1+gVnBptuocZi57KeCSnAcW+0qIxsNa4d7v/0GM9PN8R6k+rBUi68a6eOYNM
qTlquJfJRdZ1zHDqESjl5mEdgx92aA6sw8mVltyByUWK1JyWOwJUwwM/9GqGwpJm
xdvFNQ321qi1tkYLwuL5ukiIhdj3B5IXpxLAXzk4e5+n5IXOVKQMmEhSpEgatTCy
3XSDusvjiTUlpz0BwAhJ/8OP4rKSMyxmhsVK+NBhmGJW1tO/Wdr7R5PPDTgrXWgt
GH+qrQw1QdWE8Z4VGSLEPr7PKIrzXHjxY7PiKtU/Qmo6PK8BHSw4Dm4LjEiG7pzj
ii+c0EKJZOSMm2naPcjhJxH20dJSBHJaAY+KLkxslz5hYNZ2WHCnYBD/sUOprVv+
3mzOSIPQ2KqYkVfA/6AVR2EaRo9YkgQkb3q2Yy4ngpDtHzMsnwpKhrfh7r3u519t
UfZt/LUKMkOeBjdyyPlsYI//bs02ER5gde7B/6h1TkguTGzNFJEUM+5LJgusnslS
m6RWeBE1HIGWfY5DhMArmiBeWXxb25JILSX2nK/nV2amXCGgeE+TddQpzR3LoytI
umjSHSAl9ganDerFFE4t3MlsVGGBj/Nfkl0BlBw484f3/PJvvGmhxZNbFeUkOQpm
MgJzdQ7w6IT5GsI9HRUjeIVYULsJz4q0Y8FcgxRQ++/YgKwtSFxlmyO/c8AocQzZ
YRh3dqiTKa2vAxDzwVlaDCaFu7oLaLottptzndvA5lKD2CkDF/WG25hNX7rKWLJP
O7a80Ntzd5tqn5W5WZHs0CXvKsyGkw5kgGZubTavtKpDzEnz4b50hTyLMbdpLJpb
riYoNnj2HjbataEEEfnXF95gSxyFbooumN0+D7lwusbpP243yPzcFBuLX4POVwwW
9mH82D545Ia0GAnkfqCSv8YcOEYcjnK5l4vNFecO27EltwyoV2g9otsD5F2PP9Ny
xIan9XLCDawCCEsUFUEK7JaAOnf9q5mx9qK/V6I3/8IRGiyLrMuspob+upkt5Umo
gQiPilYX1+NBTNmqvAlMR+lvYN7fB+75TiAEsiWwnu8scT8pQ22hJisUiXcIaTqO
42JMoSJUseUoCCMiTzKQutG+vbOeRfplTRLpzwJeOWHoUrdCoAlZJUqZrNnVNULk
lNBIpyVq+59+H1yZtC21qS3YUJgnZQ9GY/BMqigBCvIN++y3U6w6y2EGK6fHb3kM
+jYdPDIbflUNPHrZsUaJ/HUEtDEhawwmqfL1KFbptJuV3hK7TbaNzYQiCsOMdd10
SBkzhuGn5/JlmFaUA70u9hqFPuygUBIwhoohD9NpFP3dvUQbmcHsJLHAD+MQuNlY
GJMZfzi78dtYvo2Na9rtwHQ0pFZ6xWPu0wIFtKgJz0MUZFjBnGj4Z0optr7txMZI
IKNlEKfpdzwU3QBNNS8bcaJ3FV9J1GRKxXFsN+3A1hVmpOpoX3jRqQad344AsSkq
Wc5Ypl0dCeVDOY/0j21LT0296+k0jSDJkvNrZCICk7Tkk348qgJJoDqvgbRNSxBK
hJ8NEX5unrzB0eB+8n+s+9jB4L48pVnsU5CDMZRI9KDmRmeBMjIN9Iwf5/lZ0MND
bJmmnOnfGGDP3X6SbQQzN0omqR5Ld+U8zFkL12NKD1iMSi3ZgfDc8IZHG3Cub9V4
Jb7DdDwMU8e17u6q2EqoOpSyj0N2PlRARhF/j0k1/mstQ6z+eEaoF6eA10NoL7T1
bbe5PU93WY1eK5YHr95/kMh4OpN+VE+CprnS6ZM7M/BsADptk35pww7HfsfGgJa9
DOI2v1QvJ3BYMBfLo4FdfnmaGEf5nhOvjP9HGDR/MjAZKycryi/jo/os773GL/KJ
c2nXZQyumkXLgaeeosLqQNZ3j+AKHiYw3uoen/i0VrAIBqgY8yJ3XHIMWR68lmd4
zzwKG/XP2nI/d4PeC+2iFe/pEYS54KFaN87jg2tIYQWnniQFSmfvo/qnQZf40unC
c9ccsnas7yTyw/pZ8Snw+Y2uwrHle6+POA2laQu/WnuK/x0JpJR/7zh7gFWTikNN
yTKQZ4RdKSyUJh42kNgc9EsaeA3/0pVWB5SqLZ7R1hYqfLNjie6EeOP+akp8kpsM
3lyvuHgsYc1MK8WP7sTEwvHNS6fn6HcKo8aFLSqv+C0VihSX4dzAvDa5txVw0SPd
QKS+D04crkPNI96BTNsbbghA4oi0dpX1pZViCiUWEd/2daSmeZjShdTfPUv/fbvH
nPZqfWg/GSFeKcjDnDlY0vMJ+Q1IPgx/EfiFhisviXtoB06HWFnQE/DI26krJCZw
pOR1t+ePZFf5GmHtODxsFAXP4QUf8YA+gxNPrZOw3xVDxsYWNGlzZT3tP4rJyLwX
NH9Mgf4af9eO5mpyYrbieOtSk085G9MrXExx79zYqLhVtq8AL3+4MNjk8PzckXP9
ChZvcKIhqV2sL4RmWE5a+wigEgma/wjLezGGRBrHrvG/rZVwMRzUqFWEN2pjieo6
ifsmJJWjwdXXx5p+b7s+Tmok713wgSzfZWIUh6mECLPKmg+rdhkDHRZ/+LEOBBpw
55zQfsrDSZo+S86K40VEqpgJ4sozInP7aB3ssIpibCPFlHqk04EkA3E7EsisLft9
lBcNNguT24/Dqwr1vSVdsoIQEqRFz0PRFbnuOpYScHJWdxPuvMFafUHWjbzBNOGP
ttmq52VN+a0kEofjKpUXYlQoSoUF7qrB269D71L1lLj/IqIE4yy/ml2SKJKDmq7C
8BOeMTuue5Zm94ELkZPKveNqHQnjxN8NQ9S35/SK0gmpIUl7KL/iNj+4fS0f51wE
f1v/aXgkVSyOo0WFEoyCFuKgF9xutXM5U69kLtWuFMUv7mFXZ/NLhmVKBJeNuj4x
I73i7GYGSjkYebnTjVRLkPxcFNPX+pXntwk6HOikKxaVAP/ppPEWFtXMaA+7Sg5g
8Z4g6Hnd0Od/4zYoyIggtqC7nHeFW9jMSHdIM8jAkHVrk0XKE0SSvENSMLplLnOS
Trq3v3pFq6o6fDWDKwABzMLzYV2YP+LPIyjJZPLxL9DfMpedRnQRMQh8XvjlKasG
Ndcc7fpshBIs7ADUXkn0bvI3QnfuQFh3IfP93/gI/vLU2+g5fWhnv41p36Hltb4T
+i8G3PKk3oljDJM41iUamINgftvKFt+YHOZ0xfadluasH2tFtjApOpIz8/shY3Bh
92ze8FtZk/JqOf5Oyex1O8SMbctBPH1UjjG8ryPdlmKy0RJ+9U90SELFJkfWOa2F
86eI0Yjtuzs/qAYalhfVECN6u8PA3wMu8ANeM5N1DcbRpfmH4JN8bLQyNrEiSRDK
cgURxfHENDzf7hkge70Ld41PCG+blmsisC9zAAE48R31HBK6+y8fRl2NT5OLRbq/
odOk9nvXjHCIKZ8OKJEnkrChqggE3HDQ7V0KIrAaXYzDbuPeHDfk8VFKWlHbG5w0
dmKc/6N1vYdq244H7ThJNSXQiN8n0kjGqxIurS9zIYf3jDrPhiN1IAqfSDfeCqVD
cNzwx79oiaCWr0b2HKJWoewDRfeQ45oE9vBLRPtQKcNXCWcX+ajDOcL/n1k/V1Oy
mTRGI1jiEIjfa+VooEkM6spX0rBqAoegQ4Tuj9wYDu1sEgl0U6FsfTi2FcdwuLOc
Ui+l+pf01CIrhLZGiZ5EnoLPC5/2xgxU4Btw0eHc7RHt461D6XASaWq/g4KXs/7O
t23dbggyuehYy6NIz/wSAIijPYNfRruHVEBSBz/YONcA1wVWqW27DGUb9uv2Pc32
Oo8ROXMYM/mAQgAM40NNS2mbxGabfApz0tQDMK2DJHQLQy1gSLs0d0uhkZpZ7VY9
s0nSibL0gKR3nxHVInoa0fmY2efub2kDHr2CEN5NBye/Sh+nCkEvym0g7kYp9ss5
z7mR8mDA0T7AHFp802l11fpZah7LP205r0Fo807ZyHCa4+knNSOTIv3UVvHvcIC0
9xijlW/F9ONLAtT72tel8rypzaVFhpjIYkDx9GuBZ2iVerh8A3c1UObO6/g++vLo
DETKyPsStUYXztN4+1iG0woYKPymVdtZn1lFFKypEBUiL0hDXjdVg/dIbJv0cefS
MTt8NYOMJqemWppqBiETKk/iy+wpexPhhnz7hmHRIAEneWQD3lcmHamOgllKZZ/w
d0sH9/P0plYntR9Q7WcEhPIlMZTmp19XaTFPJj5kXdyPvkYTEi1N0HZaZuLUx2lF
diBNlMZxHFzNVI1UV+y4Nme/l3fJObCGpcaewNSt9t3LYAMET1+eNB9QndFiVuij
74tR7f/cXTsZd1RdnGXP6inmpT/lm/EWpkd3vlZOklUsP4+dwhbkHwlJqcPjU135
jM9FL27CRMGglH9sgpqmdwGCDp6Z+fSs+BxEWWCdb2vXTlg8Z8kU977O9iLSGJQq
OrK2OkPOWHBppbaS4kcv5MEWeNLOuGTlhcT/U9NSQ0XHOq9mvyRb2KIfjDs9sQEZ
JziNuV4+lIJQ+qWsiwIiogelnkI3LhoDwmjTiqW1Jld+eCmjD7pbcG6qSg9UMP7S
uKWG9G1NqwXlwbKtQaovI1qcFXZO/bOYy51Uatx2uYRP9DCoPGiZiX8Eh4Y6avZt
Ms6uDFsdCZjE4D+fYFeOOlQKtisTGXCzxmFNwcZKuhLGfFibkQstg6cReP8tPYm3
+QMivLVyH2E67FTF7LP/o7OqlUjzXPYEHz0Xv/LFUz8ybIqRCpcPAyeWOdW0eJbt
+Jv9AJzZaiHdB03NYLx89rg6zzvkKUPAgiHTukaRlsrEIaz7r9VvBSCHyDjifKQ+
xwt9M5oUFBYGzMZpo7z62kKA5Nb4SzAcz5AeWWlubli+iF6sXDlp8mXhE4Bu9agk
oen8bBtkSm6LU7mvelNLluCfQ9T1JYJU9RCBGkJVWgHRWgex8e2Vx7WaNs9klWJr
eLKgjwzHRXno5Rvus5yHgqX2X2PYWDY3wpvdTQrtcjO4Doyr/lyO/wGuLhC/Gowa
FRh7htV6NB8L5kTzRzzZ/8n94kiuHAILmXL/SMdHyti9bbNe7CziQKG4+qcq0Dpx
pwJr0xLTRrpt10xFZ0XqkATMayJK7EKsVL/UmRt88AihBWDB66ZDHy2JfPQzO8+P
vMbd1MSRR7QRFC4QgTGF9G/1NcV8Ol11H7nFfxtqohWJcwmnWMCxuUNdPP0DLlQ+
UGDng+8bezPvyAoboYCNzsSayvS2u1IE8HdaBRImADQfwoDi15Ond1ob80v7syNx
wrtX6wgcmEHXZprqfrgiaS6cVy+/jr7jklBI3MfROjZjZZP+kkqE1A/4IzNbnCEp
homezNm+vqOogjExTekKYIP8v+YJefTfOAjBrk3su0qG3ji1lFjGsUhXniQArREt
nWd9anSvlEjlfej0lWN3iDH5GlHbuemKVoqKK7amk0v69wZ+SGCnSP1UxJBY6af2
YSCbqE/t6RHQMDdqkhMPUBJx7WJv6KoZzIu1CU0Fx5vxhf9oZav/M9RJOiigPKUt
vMLLm/sdVIXoizEi9KnSbmxKIaMEqJCnYVW1tg7RKaIFwz1kEBV4o31njuRjUP2g
xfnEIG7KiHX94ifnA3nUnkOf45iozLAkqMw+GGQHG4KYadqRuvHznkYELrHeDcfo
SCpZe+vNF+pSSNx7a9x9PsmAFs3wQQIDMhJmMlZikGj43NIIIBg+l1KP06uTYwcV
Cw+oVpA2H87Xor6LsUw1Eg4TXVD0M7lm+Q/Vzed4/lsHDekgjQKXQAN9bThJNhU+
HCNtS8G1kayCFRaGyx1O6ZtuiOkO2SAeq9mbg7floX8dV3fTE9eczTAzBTwnl1DN
QT0+h9GWtzWmyI2mzk4r3eWaY05ETeMWh3vzCc5sPVYu6CYsCjJvy1WBUMBKsnJL
qoh6pz2fV2wnYhrFvGNaE61UX92vwaV7uliNawtwt2aSNtIX7ssv5eDtlJG1hZWm
svis+blNioBZU3exNOEcMiQOC6pO3WGtJwB+hFpecYZrPYKVTb2b/mdSs8OaA0PC
SkexE/gFw/Fi9GUz7+T1cXd+aW09+ZyMZFMZhHcoo8/1DKZAfGBvYT0B2VDvRHw6
452PQfXcwCIoZjSXe7N62CWcHCTalRw4L40ClXKzpbcPVac5uAZq5q5zv+T9MC5Q
KerW3yKg7wVWe05OTQCEesXaG7bsg8FaqE+BA4lnX3jWmUNclwZwJqy/b2eTMBYR
JKDMf2c+0RezoDvhKxkn+sp3eQ3aYoNYnsD8wvjjYBdoLKB2F40rj299+4pCYQqN
pOs2kIRsMWzym+3m/RT3pD3Exkq9WS4TNVkQsevPJ+fFvNbuSr2GR5/UGOVfDzuS
bQgqLQ/1BtfcU4DfnIeXUu0csCKMZrBNTVmKfzp3Ym8fdUw43Vr475CsjysNGogi
kn1nXbk4IaMh7Hv7mRtM4JR/TCldHnmkQ0pxqkOqF6OYwuEJKnT73OwCaeF0+S2e
Se65UIh5htIRUcQ8M8NhNxpb6ReHSnNmFyL6HD5mUydnaOna2lKdfYoihrUDzzWY
4/p2ugDuBggl+D1wE5EzBqhTMvZ6qkgDuXpN6iPI8/ix2QYL/Np36Xq3Vhn58g5S
eLdIPML7rpIpVs/2N1h/BxmirUDw9S++CwcrstiR/iIBN6GBFIww8HfwXEI1CsIb
Cexb3ZBWgCEukaWAzl0XSycF27lfL/dBlcr1yNBDzdSvsZCDhRC/irve3BQiwfVF
4tOoeNSv5KzGmxhUiF6ITXnbXeGPQibI2+oY9/tsTGtF5L9FATdlOoNTOqjT/m4h
MY42gSCI9g3GOiSLnzHz27dNUjI/WGPin31LKP/wapHSDyIzTQ9DzyNcLQA5D+/s
YlBzo8jK3LSv3K8eDrp5AeehJWk6z5Nf1QXsTDn2I8rBqbYn6plOSR25pSvGzHuy
xhQPvVlEcQc8B19cuk33opXmCmY4tVeUx/2lYG9LtEuzJpHipVtJ/2oNC/GLkGkQ
eh6+CxopJkKJQgDBYcb5pX4rcTIX/pdXWI2vM50j9Zaskq3+93UsHCEpeiCxgdRm
8hFlm2bdeXsgXKSgV116c1nm+Z3njH7kwent4eVkG0XkTuTc8qxu7Rd2zFcKjkEg
JIP7kwcTQxNXRPJXdE4Ehet3vOVHNK8RRWKIJjaM99eVyiCc/O9DCjXdnfrNflfC
cu0u8L12b2NTxg+JHtzzmubKBxB74s3o5FajJ4ZylKaqx3ADm3xUixppchWIeO+M
KPPv/2IicEKb+yCH0nqFd6/4UJwMup/D7zbe15SSg6Zf4pQnKHSXqkbMKFkqpshq
2c0nweMq2f1xpJf8/+UMtVHN9d/DQtYuua6AVzM7GyLHWwXRhR74V0sCmHjIC0pK
zawBKBBbNgHPaaLnnbHET1hhsZLnJ6OLI/H/TKYw+IRu0K6xsgPQ4G2FknSsioAJ
qJRPa+L+V345tN4tvgRz+zlVhluBuH/EH0GhOa+bhteAKs2QVm4gQs4Y+xBIr8e6
28HARngeR14S/UqO7HENiTqh4/Nk/V465/dVoOEgYDVfOjsKLKg8i75C0plomcD4
2DvkanRvoITBrMYOw9RUtE7YrXezPzX99FNMiPehWde7k5+8dWRtVfn7oFQ8LWva
/LrrIAB7hHa2yUfnRBx3jUb2jvyO1/Q2af45digGuPkSbIVBHK1A9KnuW/3OYD6f
lCP+9GCqoE6j+qKmX7mu62i5j1jLn2BRAhU+XUxH2tFVLPoz0Ocxwi8izPDuuN2m
Wocx2cPtLy7E+LR0T0DdhwQAMc3rhAx3nlLfjCfIMAdg3ezD5kjEuOz4DeG91t3Y
2ftJ+2zJjzB+IcTaOffdZPfuZ70DxgkyHgHSK0VAor2ENWQrUw8ZxlQ8g79vrzmj
DdQILanjCsHD+UriLySlyg3Ze8Q/g0mgePQyzg4yxF1scejIPzlQGZphFJO1x2pD
KSapxzLBFY1tDZKxJCmD+5+w/iJ7Xd7IRmmpOn+F8GC6uh/iM3QHOZw6oUcnNmry
q+tjtA6Begk0AzPU/OxSnC5L6HPEwcG19JoAHd1yj+ohX50lYS7x0jL/hE5e/kA+
Vo1OIjlZpDLksof5CNb8zZBDSMQdE911WtdL0J7TQVPr9DMU0zZ/+4hYJtu6rMQR
AVhKo+IDsBqagVSos4Gmbqf/kMVunsLVTl06hqw9Q1aRm1r1n4qsgi1wnkkAOywa
qhxWG5njcuDh0C+7pKfrGZSyOZCI0CSqAWyn/FTxfDxBEQ3aC3Bd1bygxtQxwX6L
3Ggmfi2L5mQ148nQwB3Zy7MHllEOD2UxJJ+3GmP9hxAOVmX/D9AHAHrLILqiTtXK
dzTOSDB1RWUutGjg/q3Z1hyi2isdcAqFWVSwoT2wDwTV4J1gZ2AxMcdqwl7CPg0v
GP0Ib2sHu4jhye5AEFuPR8cpXX0G8rcaUG5N7RV9ZYWsQ3zwHZpdGAr8BPfsMI5g
4L3Fucm73u80B2YGHN1Q0xQwVWVwlPJTUgIbkhkK/qr3y+JQZG0G5b+XU8iYLcY4
W17Ig9WWYwx6//ErMLN2Xc09nd5TrN4AEg4gQQW1biPRFFGNPNMtsKXkrprASol4
qcwI0iO37CjfNYTr4gwL1iLSgJo3XR+gMQS1YNMpd8XwRTj6ume+3y45j6mesp1U
/mulanUBXoDRC9zCghcyP+jOx4n3Ga85/YUXPZImf3cKaVYTeBEUs/1P2MJAAJx5
y+wCog73L1F732lggLix40J6bVAESFgUCWpYDtGaJzS/wpmKGIwKzIMxDrsncBDE
HSvD2CEVoyAsU/8SVaHs79jRgnKIKnoIOn5Cy/sIiSZNDpTnN7darTacF9Xtxvqy
jqLaMBR4tgrGk3KKadHn6jEZ4taUyHwM5uNZ8aWKGf36Dmxkg3MsgMLCiW+GPxH1
Ahr5PYB5b4KNPrXggtTDu5FiRwIhOiw2xV8zauUZI5V3AvLUCS/bkluqBtTSjsWb
/Swn5IvP6U1WdTw4S9EKH/7vfJ3wb4pkBToOpaMigLIJXGaLs4XD079G6wJg34+Q
WpdvuI7yAVIB9Oga9stmC3p/cN49yW/z99HRip4ngcVxqQdQ73K7WiR7nmDf8NMb
699b5K8Qb1DVRCvkyWqASFdZOGjRur3alHJLTeMp8x1LzJi/9vXlM4T5eKdY3rHZ
/sX1KK/H6XSXLmjREPFYtZBnYUTEwaBGmnCtaL63Y90WVYWYdaA/Cnudv9PHqaYq
S0ckwasnwtPF+jSmDOyvZvnEw2kLWUkCmxtFGjwxi+JYhCRkbCnZuO/LuGIZa0zL
J0xM2MquXYq4i/+Ycl7xDxowPNMAAD29Rf7dyqNlzGg9YnPVSWqBgBCMNbjh08xr
8CyTNTG2yz3uNF8fztNzo5CydNepKTTvxpTyLpWPuHdpGllm+2qc13os+PuZXUdi
fnxoXeApaoxXiXKP8pCpTdNkoYcOr6Ry1VyTHLHDmNT32iWCmLtD93Pojsd7AeMR
xyhyR4NXQ/1fLOo24OENYq7RXb79JqCQkTaE+2wjtGog87sHuG3yiFeiHfOaka6t
h/jnWe+aJkrNKtW7ucmrmnMkQhdYvc4DEr43yVgH4o9J0bdRnksx7vjfBJmNTaw4
9H5CN/nQGU8BNxVRCIU/is6xd2Kkm5ZZK4LMX+YMJBxnn86TnfEMtM//1KMjoxUw
GzuD+XcB+moeYghGIuSvUtw1Q7DjeIF/uHJZM0c4jXMAxDZphCQ0ztgg6IUNHHAE
/5L5P03lttdU3eBeatIVvc5r8zidpgehVbnSbbr9lQHzO5KP11diq+IM7XkYWEtM
FRX2C2vf53/ACoSdYGFpaFiJ8IS34nVsCB7i6AIGT9Pxpdyx8BRakIvpX5XZKoXF
KRzfF771VRzkgv9kfyYUcIt5dyGRJe6KBXHIrFfgHgHMhEzawymwngIfjyX/es7J
IM6s+0WV2kEg5rjCqPeB9LYXD9UlCay00GEvt8FExHS+39Y5QBYkV/o3XE+S9wSi
yldiw46TrbkvKvUhEkTkouE0++TppOnh3UaJzqK/4Mrho34nVFxKPz1WkjBu/Loj
tjn6IGB1VsZ+CUH7RbA54Xccu7cpvVRDXTVCnrobyYFIU1s3aXDEma/WeSkvRbr1
cT9uT5ITA8ocs/Q4GhMWMPeCv9W6sIzpoynCEigli69vw0GjWOluWu7iqRYOJEWT
+0c673yKTT52qa0+3LG6edb+ceN0aitv8RZpWgBPk4KQl29opN6FDJNCj+zxkoam
LTo7O5bzOUiX4ymCgjSQPf5ywYZ2H+xY+eXxxzjHpu2dCXkyf2LxYHe20wUVFtgq
I17X/fLNPWiDgI05j7k2si7Phz5NAZtxfAw41fel6XN3mkrAxRhZNC06am8CD6Bb
XChbZZKHD/U11ET7W8LrBy4OxUTR90+O/+drK6E8B1fVpsfAivgc23Q8sWzrVOk8
8CNtUZ/IsnV1hSdg5E6icqkFhMHRnR5a5y2ATXnJ9+Lbyl47yhBCsBflmpkwV92B
xN5LeapxJ/YrjVafAaPjhYCiP40HmcJdsfd4qUHZdWdJNaIHQ0ozEY3Qc9s8fALX
ZLX2bp4lsaOe/+ggI/IgZV4EyFgzGGCXkIxE220IV1Iq/ni78jU21uEVQBd6p+O2
mYLBNJ7fo26rzHad1zlsPs1hTCGCaXtOMvzvDQdB7rfIQEeZCJsemTIktFZlwqUE
u447h0/gkt6A0KopLnGGtEWJ4kMDNP4bN+tvwVaYPayuq0bBaNGtXOzL1QEvzhl4
A/GBE2RSvkwymQMpVvXWxYwue5eNLwFZUHlqY8VaJj4wB90jhOzb46fqLkV6+r4t
6GnnpQd0/NIhQvO6etS5fZDJ+squ3JYACd0ibeDKvSu++kFsV5V6INZcy1RpSe5O
YLcVTUvR8QCb/+DSBPux8o05FsdMTr9TZKp68Ln2BzFBjL3Hy6Rhgpl+WsyMJrMH
bYeIRiy98vz8Hk2jUI9VLZa/0SU3V+D4n4xCCM/WOijCdKKJVfKD4jLNjbq4esVs
FPrsK4OUMVaGdxAi92+eubTdUAdG/rD9/+WuCcpoM70zcRrbWmZrHhCE0+0eFTpI
SVfc376+rbBpTFyBMxFEukwzXf+ScWx0r2REs29RISN44U2k7CK7O4X5TttxZmLn
3iMvaoj8KmP49+mPaBJHOyO3cpewCtMPWxBxltQit5Ubv9ObWu9HgtkvV7GbG1jP
3RASNUMqdjTXoiPulE1AntSc4KS+Vi6GxWE48fgUaSgAwIRBQ90IuEG9c4/xn8Pk
KUt3vHiWLRgvict/XM83ic82LfIMeH7aQYg73h1qcRmGXuBofXc4p0+iIT9zE+wf
B+3ByroQ48W5fmr/YTn8TIdOR2IgcP9XVdI4MIV1gtEBFFDSWKlGLfxSonZ76fLp
xBQ9uV8jR3pooJE0pqlrcTAaRSBw9KB8ip7+PCAQFlpQKDOf9NlZIMBp1G9jGv2B
xJqG3rzD3qhMG7KhbZ1wdBZRX+cnQCFTgY6kUDCI3jkcIWeL+JZ/7JxhH1Lqf8bh
REJiM8TnX07WSeaw2VLNU+rxWiR35wgT3V0hCl+LFClHJEh3JQbAwlj3o+UzW6GU
RnGOezcONzBWE7gQbEuQTPNW9yrTypBJl29Aa7iMpPlTKXw3oR7zW5xvJYdaLcnT
dy8GXDwuBycfxMpYsCvYJkwRQTbFd33KssFxioVsOSNoS8pZ6XHXmMkg2VfQ70m/
SntIOaPs7U3Hnn5PgK1856/BL/k/gGcOojJzQF7E/WXPos8Lh4gDUiojwIcmFdjh
vuS59f4P0iPokj0NQgg5cXi5Z4hIln9O1aXA5t9BAFlMLh8YuxRjHclvP4E3ZGgk
5cNxsNnawYLcVWPR2EnHHIECfqvus6dB0sgLVOul9KjWxRdf1DfBwSXic1jHD3g0
9Omn0Z10EndYIR+09sX6rQTcCMHQbCjJudwYSk42f0Yiere8gAGpcVt+OtQN0m2r
XpyxZQhWVtTl6F3kEBszn7+CjvfplON6zVj9AGcMR05/5/EgYruo40D9snfvweBM
ulj/NqzDLjJK4au6dflwG7hb6NWG0JDvyO6tylld/UHldmtDQAsJo2UhgLdljSzm
CZGI/bcLd5/eONeYFyDJgSOPC8pzWVw2BoBwj8mDX9QiN3TsawMD80xJS3gXJq7x
L1JYl/u0RlBOEi72VV9C8Sh/gJxwOSpLnKXBPDkUZ9/ztzpVejCWqbw0Ge+gouN+
vVKUBVqN52gftyCu75WmX/ejviM6aFTgNnUVv2C760HYElpZVp8EENAY5VLEYCeL
SASNbpS2SU8E5LHwriVKYAO/BWZPSE2zf3HIyvIwIBegpdjBWpImmH03lUvq2f/y
Xtw8kubeIcXesrAQCArEGUOcyAF/2s/c9SlOsaUSsjp4ti71Q7WI9smk+ld875yx
FWzSLNh10pj7i6ZdcV/kqaLbn9uxLYVehbyaixE3VnQaRJTa/i3+92a3oxdu6gH1
KxQ6XhbXPu5ggEqr3K4HELfW1gxJvow1+/wzUCgmYv064TAPYupjS4/4wDpNSWW5
tb8QJMke+0E5mAksl8Nx5xvja91i+tTOMlWiqA3BWcJcRy5rPN18uvrCDiYpTZdX
TtmJfYqzedPgnOa/9LWVQnzWq5CyhbJfhuqtUqiYLgjO5MhKk6kBPtO1oEvYKYzY
P2k/9xXFI7HTatVCwLH5KKw4UrN90XTjQ4itC6XEegH4iTJAs/hf2+8fidZHa+xu
4KeU9I0UgO484XuEeKkgCgtbbluS9mtnx3g/FyILiBmMZMrHHmCrNB29HgYbshZm
Ti/WxKzMlirql1RJMvSKOzSkmnuRA+vvMGRNR2v/jNYaOkj44shHXZ7hdpqDc6Ic
t0TQAVEgq+n/fuhufP3DjQJcQp3fIz8p6DEWYcJg957MlMaHukmgoCQMgNtcaHGB
3+20MZCoxF1WLuIqDHPhv/GR+gwGktUOGUo/sDyeL3xbSQv3sr6Kor7BEkOYddhM
qHIoTQb0cAuAdMbxcJaFFOrvGIXrNthFSksTeAV/7GRtvoAurM3Uhx5astN1+9Lf
UsWZk8IkEU9LugnQiP8QAG3HLrL4C4SsdFNwYZs0H2/By+2idFw/hYtqf1ujXP85
eGBd+Q969BSNbxFTKAFg+gRVdGB9UtyElQP+UYFVE6bA2EMuEkfMaAF8I8U5lZDk
4mjbuOerJkAPZWMKye1XvSmj9cQIvY/ma15lmw9gDw2GTyDOG1XIkwE3j74RaZzo
ZfRnzCT0aYLmTsc+EPmoaOHWXJi7mo5GyHbRr34pDDeDaJ4Bt/UA9FIU/RJm/mF3
zCB+E905lYFr1KO0PMspiljDeZPlO6dRvlbAqsyajZI4IH34uP2yU0qUmUd0dTmB
pRWjBH3AJO4puzvfT4ev9yyU3NDoTZo6B2jlRc3hb2TP23V3hiFnf0qv+pXyQOwt
10uz/VvLKRmEirLI+Jysf3UaTgqP49qj00XBUrKSrBl67tU+RHunTo9/VFcbVGms
8ZusAoOzTKcKxkrr7giI+a50UzecmXdW1TirggpcKt9aotC3973bsTpnscmCQatS
W1jvr8GzEbRnOme9gQAYcWSNq/jzv+YtALouKfu0lDHQcUGpVyH1d+rHj+0fIYOk
fApjfplkZZVTP61XttbLguKYsa8owJu1HWfrjvDnwvqSNnPNhZXrCHnKtaWWPOhS
f7Z+j/KQWKw/vthUhGfpCLELd6VqDtdxWE407+bYgo5fu6vVrJUlID4BX0/a01Qs
33EaToOdoT8wFDCsEvkoYIeGdHadZjdXZGGOlqszIUEVxeUCdcInaEfJ8Efu38y1
UifzMIV9cyZ/VZPmHD2/6YQa/4sjQh0aBnaLtSsQ5tR03VBap87PxuVG9H/PCS5i
oXJCBSsmeigqTgVsOZc4vHDX4BXnJW5r0WKfxNrulXjfAFxvQ3+ctx2jTdSlYLIq
Q6dWWovErfPerlZFho08xg0jI66/McHmleCOZB2XbeTIUlzKqhFBSS/xUizRy2s9
xzTF9zjrda2OC2XX2MEW7QZGORceLsOuxpzDu53RhWdgbDmAjLslQq2MfmJJdUvT
/bX/C0dXPXpfzin7oPP1TC27b8nMS6d5jJIS6tTXOjz7drh35Hf12HI/ryURlZtT
VDzeIS7Ft4zDAQsC6dGb9cOVQDxOrdZrlrC+aLoEbEzJxcODLZJEs3p1hdj/O0Fk
KPuQoGx4NrbgxHVfWu3px3EDKmUmZkeCMNpBL4r1HJTsPQ4ZVB/yJPMiem3QRQlZ
aFXq0GViG/3dIcPE2QegGtGFk1svpMGPmm7L7aX2du9bYUVZiMqL3OJL4dOr1Iht
p405Gl5P/LjJ255wxD9obHJnISezXUmugnw837KwJG+jelwfxB5iKW1vtf75RhPC
833Shs6Ix24GTsXoJOnPa11KlpMTihnDBZeM4assRd4hw98mCHYjFDnj2gaJFRyw
7/kyD6TkzUO2Lc9SVKqcJB5hIXo/zEhixGbuyxAuRIlVzKey12UCFF4V/PCh+AvY
zqJGQzp5QUNkb5zNU+mgDSsTR7lOd2TJOqyMImswe+JHwKsDr09qADyCTUu/i4Rc
vI64oJes+NWl1av+0midu0Y43TRn8dqHzJvvENptu2hx7dc6O9ycsGowecYdamy8
k43EQ2arpgM9Rcz0n99vygp5qg9y/SAZyYtmsTAFbNKdgU4oxgDSpygUP9o5k6dH
Vw7MBQhzXZn247uX0X/XteiTHBjhqNeK7OLQDgJjZ35vPpNjYM+/GnFlwSAd4Mi+
/GCQAopr2lfEc9Cz1xbV/Ga9nLETA8CPJsq6oLBFXGCAyvjFCS33py8wsFHYVlVF
/I05/8/r/AyZk4ruROWelW7KiwOuTOl66MBzhfEuNlXTaIy8kJNJB7Dmr2aOCOFC
vQuHCERj3Qi2ACqpBpgA+J0F63p+CogoTLOCZUEv7TSCJOIbczEwSQB+FNDqr3V7
SICa44lNj/USejQVO/EACH0m0X84lx8LeXe7A9Hfo8Pn5akIamrGqmSkBxYClqib
0aGPIG/tOdVn/BPDvLPuxpuFRVp7+PqLVSc112CHyO7XQOIAviuqG8iQ7V94+5s4
5rSw/gpnoLCcWZoukLwcPVRXfrZTCGJx9FXl3lvbVJX5e4HKBjNus5WfzmG8Xtuq
Cn8YHF5CKZ/MXJY0HM1tdVA1XWEKBTWyHrCoeixEntfR8kKWWnqxhD9KAO1ibpaw
BOIYaf+OjpLS2Db1ojy/wNnxwINfH/qmeyt3znrZ7sC+udleC+NJES0pLtX0Rb7o
T21jYIzcGQt2EHXwTeSH8rRc1WLOTgE/uWcns7sXEOPCCuYld68g4c+xM9+RYr0n
Q1hxb6499g9LzEV2XVubWYCFlG/WHi9/6iyT7a3iI8Ja0EZnDuVOo/Iy2OYDr+wf
LV2hGBJcFfnMhYEBwmo/Gu/4LJU5mNoMnu1MNAcyUr9pxD2SdYZtMjZZr9IitShh
huZp6ASBSIln7DfzMIA2DEJ7GbP4NzjCSuVjsLge82RrNHtl/41/2de+ju902IoT
iaQm8VxoG0JF4XMP0tmAx++FXCAkaLWQHkv2tETfbsqylNRXU+fnOW4+rnp+HrkK
ewartCCOBXu1xxiNdtN0wdm8hBq9rB8mEvDYqFjQlo5e/awfyMH1KVvYAaY0+z0p
W08JcGDbOdQexGvm9eeRw/ctrHcD66SxdAPO69WIZvnBhl2odJ+lUFVej9sTroUC
OXekoieF/kQ9Y1t61l6kj9+4ZQqRw9eV7XRFpCbXn4OkZo4H5zamuuCi6sM+8s3e
KTsDvY2FW6knrxeqSd2tHxiHyO+ueCXHhScGnFGgaJFeX/z6AaSGRB4kudZ4Qni8
IrpOxurD8fw4ong3MUaM+pbIgox6IUVcfXkaWc0xx7XgUB+KCbRf0cx20Q5M2t4Z
SWnzGBi9F32Ml6joirw2w2PnWBRJScItWqgRzF7Ky3/FpCb84mXXnZ+IY6SHoibB
icnG27r62xlIO9Y/+rv4EzuJnGECxBF26QAfxKDdUtwEiH0/9EYFZ9NcfSfxr4UC
I0v/ctlAjEGMaZSmoTtiUmv+paHm04nkW8lfHMOFF0KaDd0/n1FjA9qHJYbAl9pR
ANUV10ki5uGbnFGpPDJeXBNZOMT3oJlJiwDb8JzjuQTNjpuVPNADtgIaK+MMLCHm
z2k8xC6+dMA+6r84rvEZnjCPpjd3ORiJ7Vqsa0qUvcUaYDXXvUm/6SCv32zciJxZ
37ygWCOWCn+p9aBIUbH9f7ePR0Hh8UwpsgsfxL9WC7cSlLnzqr43Di10yX4foNlo
svhRZJWIosoe2qRziM3mkYKsphehpOrvSZg2OfgbLqDN7mZAyAdi5in16EQvsTvo
4G6yORaTk1CYYBYBpW/pCXWXkx5Lwpu0evzC/vxGSDWhkVV+eIvjhOi7kdZODXuz
grJcmxHRnPJUU7qwKdWktb+2GQSXqDjmjzwjsvQX8NVLzaaksuDIEwtmDXSyRUD8
ms4De2pK8e95y6JpH3a3Zs81fhR2i2Rmgk5Ir0AccKbeu42WpaLXmWVG2fpH/GJY
GmTIA8J6pMOvTC1jCxFnUevQ3oYb6/ceMnxdbNEO0dB70MIngLE1YcHLqEcUIE2Q
y4g4aXici3ttAr5t1APYF3AjyGmJoIXaGjpBXXrztD49SPxIjYxfcU1MdwXHF0+Q
iJFDQar2WvJfMvMQG2XMy4s3zjN/cSDvdDohp5WtoF72DO2dCtZmR5h2w1CCym68
5kobVsEQk/q6IqaPsivbKcqwDfmFi3J2n+x904khyUgoKxMra7OHCqy7HF+0pZ8B
i7otdK0EH/MDQL6jpmwz/tvYfcJCMtGMbNV1Kvo8s3AP7cdAELlfS+NmybVdloed
vZkrgH1fDBeYaB5H/rkMNLF1doKJGXtzVgm7/8OGe7sqbvzFdnL2Dmdk36wDrV9U
swz71/8ILzWpAI6moIAk3t62+9cucs4EZbR+Sd0dP6yCjrjn0O+64I0g+ytVlD71
pVhc8Q6k91jN0KkSay1VqpNaYsM1qZeW5Zhr8nWtiMdb0bvRHL2mYpZHYOijNOK7
GiWAXpz5fJx9vwu5GcHsWMjoqnBcthVNx4GhAq5S6v+4KuxhFmWKP/8blW/ekhS+
MIC14lohCjITbJEACbTp5YpJW7+DaNgqhIdmw6HIFsySLU/2dYkecfrP5Qm/bzKP
hWLvq73zSPHx91QK5m1+QRoRWmAumSjpw3b5d/2//Kf3UaaTGG72fM5sCPawj232
0f1VxqHqOfGlJpycfMFrl8VQOa+XxSoguHeiKrrnzlnV0VpgBwJjW7HkvhMDZWU+
lhiu/guiJCPAIJ6Qh+833HOx48Lc/bPZjlesjW7l/Vr5J0TPfCB5KcRjPe0qd60Z
mdp447gulgggqbfInyFjRngN3BnappAV7zWywkLEQftMP04uCn+r6TiIoE9kWOIW
qQ3Ha5lnwqhGqLx9Zy97SsdphVHHZ/6EuwAnTHUcjqJHjYFdJdZgRvfXBnikmEl2
M8o+vJ3jgC01uaVkbXqEbaP3eiaYj44quoPljOp8+ddHAwwglxB41CK7quR7uI/L
NiZyFm2yh3IoVIQJRCgx8E1eQPXJHG6DHQoi9vxxBd5UYeoN0WoxLb90aiWhx+PP
VNfTexFtV/mT1qs/Xs/ft5NJaElBQM3siXd1SwhERtMiqbvrxJ3o07fxncZLQ4Zv
ce7C9qdmBCiV9AezyTdOJdTwTKJo381V12UQ1YYLkJVWzT0tBsGqqzIVdP/eBohT
pbSUZyndgvFpTvuzBu8PJnArOqiAtQPhW2MftH0wkAlRT6cLhOtnmqszrzk2wCZQ
legah9/zDoo6eeumvX2o16Ed2Vu6TLbXxguqur3sndT4WlqTJUhJ4l7fpSD3rH3k
/ErltAr4mfKwlQPOJgi+hgWUKfiKU6+5rbTWCHAvKQbxxp5YdnnF6urejD5V4loh
9+AvNEZo91G3KQD0skuCDYa4bmSRNnEYXN+Lhm6wBIAvPWAlaVZMCJDJzFHEmCxk
bp1Je1vwYZy+pZofaUiHdW18VLzhulsWIIu8wWTq1zd4fsT1Ka1szvFSnA2wRu6J
k0ecRm2rYgViwMB7yDw2Em7iVGAh4hDLEKTPyQdP3L35aJ/7li+6zjVBRiEj3UZr
Ujhp7YGOmGVU9LAaYoTpIOZHpbcgBEoy+a+emZIsIUTf6ayxS64nrhrx5ovySiBH
ToBu+6ZFfaAkd9o2qkZzUA6RPqjNi3Ewe6L+Ugw4hqW0Ox+LqMcy6QM8Y1pl+ouT
FayOzXE09O4nDF7fsYsXxADsWOR9g2o1KZKvaZrvqzS488wNz43TJlGLgfDGMEYv
I+c/hk67V4rLOfs9ENB1YRhrc8L/xFzUdflzjZxa5xvO+n9tVYlY+Cbsjj38Msqz
id0yFTJrW+MZALZpVtbN4LfmqIsc7CMSjiAIYGQx0q0mqiHxMmb9+oUNGk4h+7Yw
0FlY6KzFnMtpu5AmcWnf/Grbx4OVeuliVa04CL/DxJ+Z3ghhB7W0vtGgqWWbs+QV
SwkqtAn1Fsu0jqfIAoowSVanpoJWyySYZzyfrdHVgT65n/4R7LGqrPUJJVcj6jC/
O9ClvtnNHz3eWrLZA7YLQR4GGq8MsEj4LECkRjq4gxNtHWcDz+PtNd+XvtDhCRrP
cY2qY/u3ZCokIBV0dcs/rSE66BsSRjEi14HS6PCPezcvrTmqG2epAgK6zxbthbac
+2kKHjvxAQc3kpWUITp8k0skqT1N71jxN68bn3mxuiuUnYu4jpFMEEiOUgFt+01P
wlA5HVXDZXlr+OYfr5cL/0rNsg9WtUfy1a4ef8lBBGtm3WzjWyfy+ANki66tJYNk
v3Gt7oqLnOJGKlMGyW60QwxsqzRoaes+w/BoB8Ej3k9hCKOHh1N1y94J6+ru+5A5
9biOmQSa2VYdUdmx56rxNDAvxiLM01gTp1gLyc5r3A+laKStP3r0YBdN3224Z9UW
BWTWItRkcfgscR+lFbLfoRQCrsEvhurIk2dK8DwicakX6GB3OHrgRfyN/UUxy6us
CXOtNkD6NLQXrEa7lLE0N7ZGIt5obX8R0CUhH7vhD0G845RMJd8HD9irFpIGju1+
MysHQC4dJbfajfwyD/+5+wP8l3v48AJczWnqu6j+sFLF0+BTSSmmqhCls7fjpY5G
Ros9ztxfGxh1lVHz+fbIxmFMItMDPEs8EsQaQWDy57jBT3/1pOCT2P1oEqiZeyfD
WE9lkdoWdTCmA39C7DxKt80d1jcEwmizsWLwNYQ2nvh7P+bSUja7WuV0o+tq9AAA
MgdJ/M1g0YJz4aJf8rrMZssV3PPun0dRXI3eA9bj1RJNNQhVBZdkwIFHfXrIjZ+m
vJa91jcJ/u8rT9EG99SEEgYyD+Pgek9x9sSCmi+46oSWpnvGlfEmuFY7591P3h5j
kLc1AmMQLD0D3BtM4cjDYMFcLJUW1Z1skBay8PwJSFAlsC2e3vluo/gZL7ZseFZE
kaVpqMTViMM1rkvF4xexxXFUX6IaUXZTBxV+UlyoiAXtC6Z9j8W8U2SKmAqCeauf
PKAgtwk6zYo0g+BaFnXC27rB5jHGxNJ6X6Mm7dd8HRyNpKe7DSOnuxhDLu/ickP4
BSrr7s5O8QtSTpLuto6FZG1VhC5BN7XJn8mH2zV7q6m2qqFoGXm7KPuVieA4BTND
SDtzFzXir44gOT9LtAeecuETb8TRvBcnzl2SXiT9skvJ4sjR02C6cqaTg9c0X5eg
hBre/erKoXedLT3jYLB0kv9kCPI2Zigd89ujdHnmX9hGJlIB6r/o1N2PxXzt/Fnp
2k416eUt8XIUM5/1zsLIEo2Rejy8P7wPVGm6gyCVli0zeYVUkKFu6r4ZBb55I3vq
pLD7OSrDJbFmxPSLDmtvLzPiObbWHkoIBdMculQxllCpboRRjD1BqgQ13NwzEfQy
NcBWbpHATjbkYCnH6YTnFJRDPWiPkLM6NldO0pg3qQt1rP2bwaREt1Nt2snlCzp9
/0dUSEII6VYQXuQlEEdwpwSYvDDiw7h9WGdqGz9o/l2u4l255w7jSdVJOwuDW113
k2wLDAOcPtplMpC34FMRnqBKZwbbOFIXAZWs3SBNDB94E/bW0JoGU/4EdlFTLg3z
asJLQfamYpG2jdT6o+sRgkkmKkWJVBYwGLE1RMNAFerohlElsterIUd6UQov/47Z
ec5n3mycK0nd2SObxe8Vej7tX8hihNLWM0zFyr206OTbl4H8fLYwao7g4734AXCY
U0cbbmw7n8Ik0BGe66+8xtBEMTRfI6VPrOGjLEZvqPEMkxh+cg1aPkoczFaP+9xD
Hg9DmFjlKXJDPF2umb/60QaSMJ9wkVveVllkY7Xijoj65E+QNMiwbIayMhzCgZ9p
uuc/loHx5vT8k5JGAIlEjdD4YB7itdzg6hM98ADxHjREWMn4EvZ/ZHk1yP5m+8dY
6g9obF/tB46kKCW/rnYCo3ZlNsJV1naGa+D+Gl+bmJIiIe+2ZNd9WxlgvCp2Siym
fBgsJQM+JP2pgjKFLOM8yR+HNjc4AEE0OltZ7Ag2GJnNKp5kVFNkCU+P9F/y2eOV
+qJux2RTvG8W9JkhJrtu5C6ddU8cWGCXT3MBD7agKaied4nco2+wk7Y6D/vVmNX1
wFECd/Tm5VyS5EklkwcC8MGBDKKd2pHfeOoriiNXJ2VREtxIA8jgdnbV3TF4IGnW
lIwjxq6phGzq931BHzDmO7pUnQG2v2DEUh5dPcrdBI8tnjSSypVfwN63t/VIMixR
kKlbTDwAjcnmfpfwIqGLLVXKGu2Cp2c8USpZJO6ECImspdWpandBWO5nZY4TOd3Z
uvU05bvDibgm7hLrUebWUurZSzmBZINvV2hQvo7QFE5V6kNpajxhaoMBWWCYOTyH
2Kk1KxetqAIrft7itC/W/9zBX4ONdti2matJ9gMUI0s7mmx5/uzGM5XGL37/GYX5
hqbglXfGpTfcqB1WeINK/PHozIe0+DZW0OPURPk7oDtgS6tJV0ZP41zfoZoPWLAL
mXiM45PBdlHONMF0JKLx9efJeODtJBOvOzA3F9Yn1AYM17NcBAJl2L7OZv6pLPlM
i9e3+lYSJo6jbuFJxQdYv5c3t5ekfgy5/CWGYhMxspEb6EDlH9/yNgDwkO1GY2ma
LFClg97ZaZCIFsMzVWYkMhcwhmQ4Da6BqoINZUQSVQZdIlUo865RNZmphNlwgJZ7
jjkdA5n6kWrtTRYRyKcmIjS07hWxxziV9wrBCCA1RetL5PQeQMhjIKoyUMTotM2i
3236+ekKBHFTUkLuaRM5OBnrhFysnBxIuDQGAFYjRciqyGhUEayu2x446MCGn82f
hdzvF7sTIa4lNGQmykz8G6VOYZqM2KbR8IWxjmP7lkQ/cMsjVveZSMxwgbqIJu44
wPPTGr8p564aHALaXVi4cSrgkxyBP2wrQX5cykvPQexIQ16uFGR2xHEKlgmX8kgO
3+aXi3Tyh7nxjOswRKLLllygEaciznOVOUZs46w3WDfS2d/YgG4slemybkFh8aRn
NGYqOj/1L05F8K6cNOEG5ujvgOisgUjOEA1RYG1yhnw2gXCVdeF8zOTTrtPPG7/S
mgSxg2tNntGm7GgeKCNLhkgfL/1QE7ciwrp0qhj8HsUUVtDQPSNaSP04gko+bXEu
yWqNmmvz7Me94bPlvtHl9HeoqtGJVZP+ZW9NgnT4uWvogm48ioGMPa7quwiWlRrX
N35hT2XgVNcEaub1NQZjgp1Pmj80QtlgkoS801Fa+IEBDAebcgXqwpUj1/F4Uvg9
RtC/Na4NuPj4D/9TMKhS35Zagr6MYgC6V9YJllUel9Jr92ivAgJqGHBJdWjOuSNa
LDOBbsirinVUpkvOw0w8ynzM4eA/P0WYclGLsJw4/MSlhdKK+IuyaCWzWDJGrWSR
Tv3jNjVWmEZlCxxhniS9ezZd/09MSIdLWg2SOtdknXoQA27BJOmsoG4wqKa/Rmc5
NmYnAjJWjKImfgUSEap61uK0rMu4h+UqnX9zhSD387tzn/2t1GIMDdE3HSuk1Sfz
S2wOeBZgesyX0xgyitCR93I3bWTYtFTye7qaIhVYX902ejEJ9cpuWFAUmb6rxKD7
GGaAdV2fkkwKTBGa4HaNIkAdDRHbpthzOULis4uKGR9MQRoV5f1EIDyFmF5JRfq4
dkPzf9cJsoVheBnt2fujLGV8fLQbWwxXpdvi+MGLvrkFzaDbYmY0v2PbqnANPcYN
Eh1x3OstgVQM7Dl8xQllwYiW0nMCKZ3Fk9vclnJUx+qNmfBeN/vDbvSll+mEarVa
8/lGUtLgh7xn+CSTvK4ZgQyfLSTUs2/B11tcZXJWBAl4Ada5fDEpAR7VPvGyyod4
/Z+DEsB4MKqO4/EwnF1tjAfm/gUKr8iw5IE3iUGhi/mCUNnarBLA8FHYb40sKwtb
EbNi5+KhdJf1T4KFaSNY4m8iKolHmfI8ufFFJ8v2S4iP4JeCpfsf5lt9IUuab8Ca
sqBNboVgjbabn5rRr5Cj+MUjB+FSChkoOETOtdG14GJVvntA0ZoNNCsA2yWgKWbh
995HLnOsQDlzL+pJPBFkb7voJwL/SYqTirBh3ujPXYXK4hA5hz+Z0uJDP8/yh3+6
YZJHq/qWpvzFZHJmAtMs4k5hsgLh17flD9lNJuTOL5cAyQhHmLthuHAL6B8x1elV
oD0yFqnB2J9aylGK+beXsAEz81LRypo8YX8r2K4Jikr2f6xftt6ejy+UxnBYFz0b
AvctQZH9yiiWYoMRouqW9EMi4W3YEiAR7+XqGHHdi2ilUuX3v1UpqObm2PmeZP1O
2GaCkCDqbJ//YSIDSZtBZ3BGujmEh8E1McPU9Xbxp4LDs5u3hdxi9yn16rXnxF83
CylOjjJ8qdqRj6jmEZkcLPS7P3T6LnI+AWeXyFdy1Np18PicYYFadK08aXyxsJfS
Ag3NZbJmUuV6H06NoVYEL48VK3GV5kFkczpwxxRXVizHLggWPBah+7KW4bSaNq6R
CuyZ5nNgiIejNvd5dT+lDjkbSDamKm4YeV6C9BqE5gL2H4sXwbsZ48LZUG3jmeWA
0SVIWwI7IYNvLPwQpjyDtxnZ1FA3AzPTFse+YKuv6JEB0mVB6TT9Q9f+RXFXn015
/cS9KJGvf87+2/khqV29dIrvm/2GOrtojqsFTYWUDmZMUnNCoHqMa8jRgN6F7C01
d2xIIXhmagrJN8lC/hlka1HwUjEQPTo8YZfZVltjkZ6gWiFshJ5NhPiyHs6Sx4Gm
3o5gvE9JGMe1kG29LEd2do0DenwPp6XjuE/8xgPPQR128y36cNWJAQpa501twZNr
XGlImmbko1dAnTt8y5PoiJgDLppQB6wYvHEoqJFA4n+k6pdKny6Ut/ZnxA5emugo
mYxU+5HlNHpueyQYt3Dj4tAEoZDY35oJk2cfEWMqZ6ETY/dsH6dJQO0+Z1V3uRli
4lZydl+BH7CtL+t40e6ut9EhyKlkeb5oMAZviRTcCVMozsY+abV4PkbPpJ9ClD4S
jtoseTYVRvovSbt1aWFb54639OUQCvERyDl8ddNgIRuLNQf3AEkKakL/r7h53024
Zaoaml3bYP/zxVb5HqN+i9RJDb+byH63yzY7dgurQ67U564h1YkxcZL1fLfFRR8j
Q8Q0kfTxxD7PObdKr/HYNDdtoGwwkY+Ik5D3cOh4DP9MHXlgRpxkzo5AGMj+5lql
zwzjhwGIZREIVD63E0yHDbdwjHrycsc6P2zK7nOYvidiw+S/PoC+VnajSLcZiZ05
0QQ8R6yhSjYo9WTuWHSt7gm+6aMRACFZP3JI8G0wGrmPu1u8osoaDTF4Ct2KilGd
p79W+KIu2zzlxtNz5LHPPx9Y2YTdKvQnXktLB0hg5m0EMFLrSlymbvSOBcYXKuir
o+LNoVf8860+YH/mz3BPWS2pdvwqYoU3Y/F+gPKKSHriIG6tUAn/9K94m0lqdsbk
xy5UfhQ5aHN742tgMuckg4+0wcuZ9QQbU8wuYg9iT3nOgn0H1CxpvhI0eVfNDFgU
7EJUsxp4K7/xJI7x6uc+NqWY3GvMlsOdi6Bg8E9QQx+bp9Vz6kJz0UiCnhlKof/g
c7lbJLGaVk4dWV1b9UhgWuX5ElUOH9bsQ/MdR5mXM6/H8j7LbVzCGs2GZQ6hos4l
pOzE9AfmEe1GHc4OWPn4ZvEpqnt7iGbJKyGCfhAvfHCuOIlr8OSBLIj3XsVt+81W
q7xdWXsM6yluWm79/j418j22OCA+aZSOMshaVrrdVXOWqQbp/OUz5tF+ZPkyg8d0
dK+UjHECz0GgMWWZJqPyUGEqxaBUWcFH1ftEDHW2puu9EjaAn8wgtlaWmQzDO/RY
oyho7FXB54ydFqUXwrKSEAOMUHj5TgRuG43V79IOT99FoK+kKRh+6uUF+67KLYB3
EOiSYPLiKZyxS7qdv/2JfY4rMAPaMTWrgKkvBMB9I8Ch8+mbUiK2UoIHvMhGNsjD
+Z5fdPf8D0vEsxl8u/J8gJGl0Pt4LyGSnvGH4ViCMC64vR08I6e7N/x6NlQLYLK9
LHl9G9ADq4pYlsr/zBXGZ2JM16jWTn80ht1KrngQdwvRiNnxBHT9dsrxk1vwH/fc
465k2CnLeXQgXCON+WnZWGAD7KTsPe7SK7wwCrkm8Lpo4Sr7tJvQBX+LnnfAR3Rh
vwM1lhqIv/qA04zCy29lyPOyS7xjmLzfXZiKjkT2hmVX2H+/uk0AbGJQpZTzrmUS
1kKVIbfHGdCnKQgtsfN+L9KEL2Zqlt+nflqVtbbBMFCBDLOnb97hBRP01ITdEAii
gIktWU6ea00HsgngeCiuLXpi6zyUDlxDIBVjKj7sYADSzRS2vwMV31CgXD+SyB9T
G6QsrVPKU2zEI5v4T4w/5N1wTvBT3I6OZ4+BAqrZMHWj/PYgu9ODxIojZ8xWWrxq
55OL6KyZG8OT66H3JkYD7JqsuTKBWPrf8h+0Isi/aEvbSdW1BXyD+wbyUEkhqxuS
Y/KhnwrWhbKLBBHgfWh+5Ndxk6xLamKppO4FU2fZu1AiVmvhH7rCruS8WzCso1pw
OD749cf41wePyOQiypaRv4BrrZOoT3IcjTWKu8lf7/NfRjhqyOYmXpiVpAYizHPs
OVy4HutadSxyTnp47aA2Pji128DYzn3isa+t+j08ke0J0Kti6D10l+Rw2HtPVEO3
8cmc5g7MaBcd3ESC38SVeWdFWD5ltuyLKZ0+g8uv47Kb0V26TTgL2ABUn0COhcRz
7biwKnJIME9aSREbTxG5Dy3PvDNJUmA0wT6fzYIFGqmJ8pyhxidvKai+JVyTTNLZ
kJwU3TGQoU4cZaH19EGXmlQ+j7AI7mz9r2nreSH+nIx0km1+hVDH83+ws9Lw4zld
AP3gyay9y+bQ8XDUPeEDnJza1lJdeX4KXnRoimKoG8lXMFBFF2dOtY12JpQ37H3H
X2wARfO7mQNNQ0iT6aIj7bA7qj0CqSt6srzMFJpzjujeepH1B+Y2zr3BXFLhltXc
8+/rXQZMjDFlzVXhBFOk+a9HEy3BsGfwvYJbHatzIfQ+2VTPkk+H8srB4gfcJV1K
Fzxsf0mFUcu8IUR4KqchyPkQ04BAM3Fm3EAHoiXRzNaXzQ3Z7O2ItfbfDbfSTNkK
3E/TCYXkb00F606w58OpruE86A+773yKSMPdR+qV5a+S6xmTeB3Epu3I6OXSB/Vy
Q6N5EZFY8k035ejItzeBufL3P9fBciNx3feSLTwi9irHYaJo6UIRoXMHGA6Dqv3h
k/d+rZgFXMb4HyokMVSUl+nLl/OJGt0HvlfUBcE9kxQ0Fd5fWgzNB+0bKHcXgGZr
v/QE1itbLWGU3RJSmZjLBrTrsjbwicCHa6wsJGPOR1b1jAkQb7kjwK2eEpeVNcaK
wa2W8tGo8UoilQZerao3G2k/W8JXic0nH1hRi4G6/k3vXQQG+OXGthZH+YZk6iNv
flmuOiQxSK1JLpg5lBfwCU7YEy1ma/UwwMYsvhbvqg64GVKQMKyphP6hUlp+lPiN
5ntf9iUBrTijZId4e+0JjDDtnjCkGFQ6XLrzQQInfHguCIcFD7l16MifPHkvOwV9
XOYQt6UVRDtcY7LO1nV5GmzLj/FUUprPaMHKO/Gq3xJfdCLWZVyUNeikhrTm1mDv
r/8pGJpZMXS3hx6bwaJifWdljqa1ha1pETX0n9EVu0rzZ7npd4TdsXbKxRyL5rwC
8xSff+ssb/tkm84divaGr+7+fScSCALYl8O7tyf8DIkcmsanlcCqDsrTQ7NtiVas
eR5KYIWeToeN0eZ+ZjTJf+y8eNxblL90ifhEKdnpHlXVD+I3BqaVCr9U+rCOx4Vy
nrXyvEtgEmdmkOsIIJLo8h0VeI0bTdfYhYkbEc/pftjKc84hwrc9BtCyQGmB1l3V
3knuHs0UxZBAslRpR1INwI6LapQxbP9PmeOdTaRnaqzMMFVTcmA2IWf0x+DqJvWu
9u40G8IQeTDq7kJAP3ArO/Y8uYD6g4WwLYkuHhUkpw3g6DSeY7HXbSV+BWf9gNR2
01wtpCMyEievrXfIyuydrMG9bpwXTtbKQe7oQP6o5wjAp85db3JPR7oq/M85JE6l
n1kHYFnKiwhct90GsMa67GVgUoFiyRvaWygjByZJyb5tfb2rHPB/TX84+8fo7SmP
+5WAsdVsr+69gqPPTpkvB3+8h76l+KJKHJ1l6CUsa6FGzbish+7RMiQd5q7kCTNR
p8uOKOQ7FQ9hPnZ/eRkRzJ+p8Ra7r5VxJx7EZpAOfoQb19sp/ubm/CLgUGoBbY91
oWxRzLx9CJcYmfvHf9aYkCQbjGgrI/HNhZvHvEa4f6fd2WAGjhPN/0Oo+NjTjp0K
C5KtW45nXPy1NMIagKcpMXLYclEq9LzAgMMGhfAS9MRRpuVNLYDrJRVrwdireOLB
8/yxhJepKTRGGLdh3HqWBMvLtutl13/NJrEz4OzI1NNsIVU7fGfIa1lJKZCvOsx8
kUk+TvSxVMaD+BmweyfqSPCUh8ZK5gtkjzEzcAgKXQPxo7C3Dh/R5+Gze28lV/vJ
PPrIK3eb29noKARjG8coAJgrZqo8VApBngDsW4eK5CV7oTSwYIF8NNw3KBfJtAZ9
nDvI65II8RG5N4h13wlQ5xg8uQrMfOV+1lESE+97CcDQ0fH9KcKZEu0aaDc3cvPt
Ec1O6x+21UknESySRxMJiMJYEgNxJCwl5ktSyirYeouHDRjD98TYy3SoJUoNv5p0
Aw++oyUsE2/nDSN1anXMYN6KV9U/SL8zsAqMYZqSs3Qko13c4Wm6TTQJjBN//w+r
7pYbPJU7VphBpiXip7Kb6cj0CSTIoF23MFjlljpqAgTBinAZeJo6PoH1VLzd4lw5
NW18zO6Ewx09L4KI3+LjLTu3n9dxWypMfMdPdshbGwE5zxIvJOyVlOrbD3j8kzNX
mZGQ8CPu1cVCKEWrR/hZrQkRXSGT1ZsNvFGTJEBPogEZ44Ta1siKgR5kaUjPtEfE
Y0qF8I28HC85LHrrG2vLxZSbShMQqhykACqZIPW2QEhgwccLbEILW7GVeigrH5nm
jwPPE7IAbsvPINUP/7KjwO0b2oc/xUiyCLuT/9AMOm/whMbEZQYqtmMYUPCeRA51
cuxzGhIiL3fQildxRATbwlsKnsnp56hZNbaVB4fx4M5xfMexzFpqbvYiInuAuf08
YyRmObslnjiRpO3fo36yAhYyxnABQ7RAcLGdqPe826EEq+w1zyFNf4UIE3kEOg3V
IWSr8BSOVw1JCbTOtVLD3sdgatwf1paPuxjBWUqve91wZ/T4dkpTHPtd1yYOAOod
mevuJdfLkTULdu4kvYOuHK8o+e9zGREyRSMXr0VgkRQBnZE3Ton6VH5Jrr9RGUGB
+nKJsqPe+OlHooK/BiPjxZ0JKnYQGI5+vFzUeT3sPr9tgDw6/c6ug0+YH2ep88Jc
1+N7LFPg4HSXOu6DR8F8bdh/fzVPmlOrOB7DOUIXeLEa1F36bIhuG/AMwz/yNdoE
d8WYzOkdAjwRAXZkPAI6ALPJGlnSnBbtNGQTW1mRCaxIqNVljloSnAHI88e4gkpW
RQtN0iUxdoSwtALeRbwNzDGmKI8fTJsAkqoJKdtGJL4zvdyKI/CAc8jU/NWxTQV2
SaSoXHFkJ7a4owpS/Ed8Bfu6JgB+0WtrsadZpXpUhT4PseGsbFQZbXs+jhfAgpGi
2108rntXLxcXyorXVj5SIqpFZIwJgEciv9TJpwXp7r8SZQtp8q1N1ia5CBKmNNw8
3qcsFJyZrX3WNJ1cL8iz5qQHfnZOn6w3//nLM3JGjp0gj1Ao5DToaPvNqB7JowEf
bhBJkCo42qTS3LZzzsbf+2FIpoL07D8+qE+sekSjquOijhMYnOU4vuR8VnqHFqIg
cm43+FEfrF+Pj/7u33dC2ry1k+jQNYzdBS/GbrBjw53UkZf/cBeBwlmFkb8xa7Yf
61ZXNCFqvbQ/s1i46R+TZPCBpceQLCYQE4mAp/UT1DRTi3166zj3b8mJnM+rUsBB
eDSltyMEYG2AY1Y6uT3D2upXap2Vl2xH3OQ8FRVAt+bsPez4eLMjoI+TUdJTaboN
dhlhC0akSkSFneRiWk09O2kylsYHx6SyvgsUSTyG3qlDe6B3sM6H8kDrgsS1yRDn
W6hwujx4kk6kplT+Ct6ncy8H02lSXJ2LEW0jCYHS4oaYvi0vNs29m9gGhbPKE0eT
G8/x55FTyDPmEm+tXHNM3gyqd0lm1PsDrvtyPGz/Arp7sbSC6n04dfcLoS+53Vvz
iidIdh/lnVZM0EAaQCxmEEpagSGoGSEN7c1J2mpc3iwm3O1X96HFzgsS5Do/mpgy
zglOARa7WpB7V8f0JH6UC0Eum9s8Jd93WFXf3yaTsHO0LEy6ttjmZmtKfS9AchdQ
W4iXHHAMLGzv8L8+u/3QI0gmHbWhvx11M8w1aH5VKA8g1MmsqthOZDwdwXJKSX0O
4kzqKCLAiX758kDFa4Rz0Asrw0QHrD2YI7MBi3xjGME44BMJ4gOXcnfYE+gV3G36
lGnDUp2uzTM+H5k12UxzFvxWvlGtd123W5h+HH5pOOOwSTKGmSSIfPB5kG212xig
K+zJylXHa5ornp/KCzuN6ei3S7zM8Bzi8cU2ACp+LoX3qyg/hhVgtrv2re1zZgKB
g/P3SbpIe0dz965rt9agVvc7GDGNUJs5gleQCoIB3IgMU1PjxAW63MweOxN3gmY/
cClolVa4dpvrJBHH1GVW8j+jAA3OMd2r+bdGjrmS0DhamyRdYLQr7DBmg/4TOu91
saqRp5+1gIpFZ2Qdms7kUNbASiXeY/SA5+kO4nEVaa2Ntjolzq59eB1bZiU3toRa
w07lBog+d/wbcKpliIP5M8gXNqCazzcX0BGZHlhL6n7tfQwzEbIWzKsaAAU4+4Xu
tDu966OnzpGOz6fU7AnwI5giEF3nQvBy8d6MU+PU8su0b2E5DjBPU5nQPUK0nnNg
cu7uF7ecTPFpjEDzJup2/8f0Sa+kNVn1otHKlmIh1l8YT2XRZLyTMvJARbF06sNW
W6ilvZv1np6DYTKLXfSFBWTVxvZS0m5F4D87JnBHpr9mRQ3GyGo12IudpFdo5dSi
dfVfGZVDEnTd6tUK7UAy7rze6oSWfGtGLbq4hs03nkAtnzOhgPCPMF7B4E4BuXzN
cir7MrcTuCLtwFelqMGg28/Cw1c8NGBT/6+HH8zYm9XE4/OZh3eReaQezuNd3+VA
wm2zDYfAs71UxaX89DKh8yRpsnYP9xTcSOmV4ZOpEVgrWb4GkN0RPUBiP5TRfcth
8fpHdWhLPmurvOhaxcFc7r73OFuerlJVTxrLMNnATV1eiQ41QQj351nNlREdGKIr
TyXIY47D3SNKUbX+9tGgcDzFS6iILnBH2OA/PwQOeFehuCwWK3Q2izuhtpc2WUKn
3zihGO8LukwGS0P07fQERWM2OwrsUF5bmxHgXhXxQg1Lr4Nwfh0GxD/bLL3ejzGy
pLAjohc2KGG+iHpyaIjfJDt3+7zdYV/WEiCoFyDvsnjKOMRVC9+zjTRwNKJH6O/K
ru5ZHbjlIF+9Sj934FsIm+GGFV3sPEmih2T/dGpurBQh7gfXV4Vx4/eUp+ay4YCb
oHImVlJfW0gQ8wMCzJ6BomHsn/YiYFknkK5+7RYdtt18/ufCtByYjVXzHWgWyxBK
vUPkcZyBHmw4/y9LBOIMNSLWPyWOUiDBjjkLJQiC5Je26AYLm0hlGwZTujhAtxce
sqFg5BgmxO8nYq2eb1w+LjrtC7FXN5yElGZ2MMtaw/0g/yKb0x/baEJzQWKgTrju
DNOMdjEWnlKhhPhLqdVGPPK1WB55xuVKKfcYZwOzlZEifvciWWEqLoAYU7uN3dwf
Fw+V7vhAhVEZ/leU2VE6Dd+4KuxLFCrCMjfj04f1BADgKz61475U35xGuEib/WBU
I9+uVAaTpMAqmUlYdkuCYnPmQMAAVxQ+OxEOTjt9SQzi5UVg9CAYEx4mN1YqgKZR
U+O0xTs0ABoeS/4cFNqhin0EK5AwILu8d7p+JR3GpKUQrOnI0oCrg5smHzluo7RI
0ZTgUEmkOt76RURP+T4AOjO68yQNFUofje0WHxfRwJtEOVa2DUSFkgGlNAMDlRv2
jnUNyEM+OhUcwreJqaLeBWGczrOT1ytDYKxqs1GE0ex1G51jYfmkrBmYM2+y6z6O
fz17IMXQCpDO/UiKStM0Y+HVfZ70dd14iVIFa/R6hTocDUHniOs5/q3bTWfrtNrn
K9NMAaXdFWSy6feIdQ728pav6S433A0/LW/JTH2HNDfFz+IeGbSQ5Kus8U/17vPz
XE5rGrHwip5BTj42lotb9tKSpO9bl3IwccEfyn1PNqJLb1LnzUOGUqLKerGPuQtF
LTTBIYPk9TH30g6X/QP7MRJBScVEsdP4+Jb2qZ9Z16lE5oBXshpZnO42uJe+25fo
QNhq8ZMw1kp6kQ5Uk6erEQnItkd+9LuPQPSGY9R54wZ+yoHUp/HekkUs2IpXUS+I
XQLlEhblIjc7JZOi3zcEdO5OW4oMJD6477cncwJx2TF+fyklijEi1LTvq4JM/dcy
jId5P4yzQ7KjINADAJ/o5iaEBKLqUGB384eZ8+VdwP8xREz9VDL3sahxIVDwSn5S
ibeAC5rfj+jmjDoUxaBkHOtzO/ZLjYrB4rCBwe2W52m49MEPOSLsBfhwplAB6Xfr
evM7ehpKfFkON9r36N1c9NR3bhetKGK/43Xo/kE4hrpR3yhSkfZPbJAJTwueevv0
+5DBbOro6peldlLHG4ZGsuOnm3hh4mbbxKV8LswMTG5Z8bRwhw4b1+3pFMhlgcqL
AAV2SL8Fpk2Wnd878K7OE/cPuf8q12tc0Mf9m185Iu1K9hWhXi1BUOZqNVocM6xw
v4r3l2CbyosDX32ooPbr4IrykYOddprArq12+tgAjLErLstw3ng/zzq6sIlgoqbj
Vpkz3o9BfffkhawsQS0wzxzstvzvJTIU9Q1M/v51rT6aRDvChv8Voavk97A1ESRP
Kme4SVRakd8yHvCe9HPUU7/L2dld2lJv0VKMGp/Ho0kjUuGOmMmYzvteKWyvLCLy
QNaGdsE2nUIoIhijKO40Fheh3SfHA+lPcZacHAkBCbhN5XVfDQICmIs8NPK/nimW
BUapP9Wz9IfksQCyIvxrtTanPz5Q6Etw0WljI9GzgPOA8zEXMdk1vkaR3qhD1XaJ
w6rd7s+MCf5v8EGYiNNgay2hwRa5s8f8b+6C0nV6Zx0wMs8EA+wAV1qtMacpFQd1
pEnqi2qKSs5y93ZxDMQ/ybrBlUH2fxtu/KzK/q7xFJQ/sX+sl16PGunjGiem5RdR
FZ3HcmYUpwLa6sy9iqSyx59Cj5rwWMC/Cg6P9oh61jAIyidIegDQvmQKbS1L+cD0
kXfRTZfp9MJenPmSHT3Q9+ArC8QT2MaR/r4k6ZwPUSHCZoOkVIs35bpP6w7C0pCR
/afb9pmyLz/v0YzpeYVkclzwsSIdBr7RuMAnjOZQhje0m72GnxRJq+kT9k4u/ZvL
KHXWXy90na+bSeTF5eOtiWOqgKR7Ltu8FpQBpnInVyvZw1gvAYriUWrr9o8E8MxW
O4fWMZgt4fVsnjXSqxK/mw9dEVXw3kRQFKpjPkY7voKBVr2eWdbUXgKhHrwAzOkn
sWo10M86avE0Zt9ULmx7gk/Dztwj7NRNrhMq9SiN74Ys7/Eo9gY1rzeS+tOzk7cf
PytN3IW3w2+xvYtDR5bRUlFUvmnQnRKU2X3lpvPYOS127yOzT6+3Tsre+07yuMY5
RkyG+tUYSArmj9QDPsTxnnDpCf1ux9hkmdvYLMiYuqJP8pkFsxwHcUcIo6zEa1Ls
3ghYOVOPNqUKsX5qSBKbQKwlXj9Y0Rg7C8rI7HX7B3TE9AZJIaU57xQBdGV2M+2R
q5Uq0lw/HKZ7aXp1TjuogaPNocBDLkATCptZ1ThIaa1Sqq+2N89eN5dSVvk8PO7F
Q3ku5u7FKrVn5Ie5iV0mOSIFKA/V08nkoTdgtOEqlbbQaJ9LfaFbP+1La7FEg+Sa
dpfFFOk27ZJWAxsk4YVQax/101I/1LhYozIO+YhkaZYbrhu6FF7BysaYjjscQ5XH
OdAnbz8xNWvfVwMkH9l34krqcAiBu9R0MklAECh7Kpu/wILXI8O6Qxuh3cUVbP4J
8T5BIcf3gObHprShocs4XFnVmoguzvqxtK7YxEC6AZuKuvVsgeGxFXe2j3KPFCzi
MLn7F32TH0V1EM+JajucNcBm+Swcuo5hHAbvGtVdyStD0iPy9BLVhaDbQ7WBpC2A
VJzBjnx5fO/bbzM+8JdXBwlOeoRgUftqUp7SW68G5wFBYjVlQpDHsjgPtD69fyqk
OcDH2JVIsqruvwVhg2DrtpufakIar79cdpyXhI9G2mzuUQX5dl+DcVxL3K9oZauX
7VUg3rYHCf9cuQkOqe1kJkamh/L+OD1q48Ro8tWkMcUnPwmNxtf3rUIxe3MD3QvU
RSPA9+IkVt5OrHV7cFUTurGVO7YBhxU/lNX/GKxvhhX35CM2SzbXIwN86VnZfZkT
7TRwWhur9vOF3EX4nREDMh2yqQOJj/BzfhS/Q1ppU5+NMC2ZLI2ZXBOgdNvACIOP
Ut8dISgsL11/peIlfx4xkIy4xH4tYDstExeqp95F6K0Nj0HxaEkiAgGsGFAycNWH
OoPryw+4B05Z43E4CfmITCdbNOMARrAlD8KXwKVZEo1Qz210ImtSOXDHExEaHfIf
YGLZowCEcmjfOD38vM4mvAWIdZsFyZ/gart6ceCRtBtKQFb+9jYbaYjrtoGl3zMd
PAuiCSw6Xe36nQE2J2ozwtYmmwnR66ynwxLvnOaTYYEZvhuTSfDbG17nzZbqDqKH
QLrgT2b75XIeT6Dij0Ddiga/y2lkjaAsEDfu4Ifl1X6AVxY3Af7zjtEpEbxjd5Q2
CbjxAJlLf0OgO1l+oCtERVM7cjhb7ubwE1OhyhyrxFbkpziKEYhxlE9iIW/VRKSw
NPQxcEw6ebG6aHWJYFsAYtazYtWS6cbwZa/fimPGCDsWLaIpFWVP9Zs85GTHUD+v
7bZ3ZRzxLeI5u/XDkU15k2ZpVsnSYUEud9zdA3VkcGyLSt0+upTUg21OJSM2722K
vBghxab9VsVdTWaflYpQttU3EYqgQmDytJEdHd832OhO6s/EYn9bYJKxL6xF5mnT
ONBcJ1k2sZ3qoCMpNDxeV9ka2Hu0rQ9bdF+FJpqC5H6DhtxzUZ6GlYn07Jg65xgz
7xhVcWT43foJkI+ZcSJxIQ801rVCddrj3Y3QAo0zHXgfZrn+BYMdXSlj/Rg1Mb8L
MrleRloe6zKvb+TSaDzb8zk5PV+Yv4mgu+M7TelR6+IjeXeH0dZ1wcqQ4az0aBCZ
vZMNmMifmgjhgUa/jYYpQs92nVeDAzxIiCoFA1puH9hGSDSo5oV/99ndfuqPNzCM
D1jxvRmMPZqqj679rkniIyiU5qe7bb+17jZP0+aYOb2l4xWKc4UUhWfGF4fgfSCF
j+g3kjAm93jzGl0xMyXi1tgGJfj9+cCR09mMiJUejt7abUTSgBPoltsGWExvl31c
UN+lzLDOkH1Z4eu9DtJLi/6ar9Bph/UyZBfdXOLDT5MZku6/+f5fogouw3MQOPnI
thNXqJe4JgPiMqnfhu5MVIbWLL7YDPw9YOzdfNFR1pIN/M1YITQjNfCQaqLsVvuq
ddmEBtjHAOtyCpkiDRD2Ti2Esp0d25L6n+YmzEHW2Axm6DyKQmTnnEK6qVh3clC7
AHKo/Hn/lmWsyrzmRf2ykQltsvwT34BvPs7DDLpEXJzJiaxcLn2so8LSfl7Kzgwm
xeUNWyao/pkSxo30VNZCZumBY7JJ3o/lrQx6X0103DTrwJ5PbI3juee6vkMa91ob
TWnjDMLcaoB4ky0llQiIZKrd5gL5d7X4pzwTm5+zZPtVyAe2tlFyS2rM9EIQKFSu
FMlGjCD1ZGZn63pR3oS4aat+0/E8ifH44yu06wDRis9t9kWMSlLDxRiD1wYegqtT
jfh5l9d22QSuYTUaux+1Pxj1qIsnlh9YtRgmuEpGLacsHyoUvB3wOMnzmF2JiOzq
UZlVpjUm41Lbwoy3IPCfwMTnuOzASyxEi59+RUUf29sgfZxkRhzdcvQTdYhYtxAe
w9M17wBQufd6r2G8d0O6jI1S9tkZsljPIJHQ+e0+g36KnTP1c4++HTjByO7EjvD4
2ftPpFGPn193hnzgOgyLU6tfDjtfWEPcSWRtY8Kpu7J/gg/Ac2RGXACvr/8p6rwE
YtG+viecuhFNbOjqbP/G0BX5wa3TrVGEpuJj11kWocET9EdumcnBOA9HsTgAeTqJ
KEfBolTrlfYxBkMS+z2KD8tzSdz2i0EKfbvy2t8GqAcILOjQTHVJgdsGQ1nCZLCk
hvaWn+s/vsuAcQvPy5qyXswRgLCuVohB5F9YDM0BboAHUtRLmFD+3Yr71yX5Lshn
MAZAUwwr1N20Z9n8VtYGOQSLADcGXroSGdxLT0vlFiCN/5VYBbClTDPQvG1gjjx5
4A1kPtCWTkGtVu39l+MKsbKG7k/ySnBNuLvjXcCC0ZqnmQjuEKOLMh3ya9gptcWL
5NiUPM+UPm1wQAxJVEuvNx9kUNdEwXAguM85UGOGkgl9pgErbahHcBi+NN0YxDXy
//2Dcn3UmwHET293EBABhSTOKWlxvs8UYop/0FdxDm5zrOyefw3tL6NSPJVgoDHu
r1e/Djeh9XZobBTBM0XOhUQ/5Rr6QPLSLqngYu/xwljc7ZFZKZyaxJmlbwA+HCbQ
SY9wloxekDE7a36OuQ9PrHzbYOAYzJNywsOHowLsxPB2da8nP9JInLwvKGhGQSSF
WnfUY6vxuwkbYuQiiDwDU0aPBEdT7IRPTMIdu7sPCCq3g+Ff7BtnrAF7oiVUjNC/
xh2iQOd1A8pGGi6LTykbh5l+8y79c9ilc9qHPrY+LwTItY2mf7Xelwc7GGwyxLAF
MonIpFMiTZjnP9nu4vZyHtD4kv1YuBiz4TthY8jQnmlIJvYRuqbu1VdHdA52W1h4
9vktY6HX9k4C+oH0nEP70xgsyiCuSpCPN7oFrnLwPeapIs7/sDhmOIz+DTtIYI7p
VKQsE2svsD+0vrO7cDvVKbBffXh8dF39FIemOYH0ILMAbA4rg0mbQHmeG33WyFE5
uuNYsLgnm8bV//gVEMoo7TPUqFz2LmRVUxf9Txq89Lg6myQqGO4xCdNHIGK0k1Yn
+WiLhbn8h39Db1LZl9jaCwdn5lOt4qbF1O32/pw0jDYUJcVzRRSxL4I6hB+Ng0gM
C7eel3A5YP3HOfxyIQ1+t/N3lg+zsRazePun14HZ+sib+QBuoMhGrXSUPpNhmgkz
VjoTC9xYwPqe7QjgFNI0u9bYEKSKr1rScv5rd9rQ3r5r8+9GpZx+YUxd7Xqqu0rx
iAjrAyks/ebR7zn92NfGw8UbSLzlpexYLbCTTrdiePq8OHgTNRHyQRG8oh0/rS0Q
josnms6EpQ72JjltfX2uxexblDV6t4ABxW2w6JYEv64WwXnzuZxpAptHv5SX4w24
ZGv/iI150vQORRpWI6xYsF56ZkVc0ApjSDZD2ETBrqrlRDq/td4GUgwKp4+C8eYl
Da4m9LvKLYUkgADG6U4/OIms6slJ80NrbZ8Yd7PsYdQC0C1i1XE9YnDi8MiH8i1f
wqvyCLa//Qw53P++Yz4uJmIDWJF4MwO6jYrwA7YxHAaq5BYOBbdK6YlkJvhm2s4I
K6evbXDfykdQrIjskNBFSoCW7AcLbYCyUp7iwQlWKLMxvpMKpcIUSoO38f+bBM92
1ajwy6xk1vXPp1Qzb7CrDCrCX8X5GNTQfjvHcZo96zQcXzImzqQDoewBS0+oSvVw
pctP7e/JAfkFqCh8bphpDBRMy/YdB5uArN6xmbeNRo19oLNAuA6xvfOHNeULypo7
fh2G6NaMmDOUw27P4e8FIvsiDY2qZMtomiGTmTQJClYCZzDoJKSEJ/Auj0rEYYYX
F6KZ4bAWLlQ+YSIPCKrQMV6BpYMoiaOz82JGjcREWlwi2/xTRMvBc4/UdmBHKs8W
vwH9UluBE25AzMciQTZpdZdf7oHEof4aQBItO1K0zgF0aXiAe4T7ul2WDfPafBqf
S2KrECOQs3qZO0K9bPS9KVbcqcOSxoNDxTwgsTgdaHo2OlkV2Sv6xXN4kAKlrw5D
WHSB38B8KdwmImxNoY25eXQiL2S4I5YVjfkBul5ocVBneW/iP90V0L/Kx9AcckQ8
EVvbv5GTARqRj2ABhWRj89RNiOECyp7w8oz0+9rENAppyBgH/yph8JgdrFPfQv44
rIcI3LiLogZkx5KM3C32Q/EFp3tsMfSgj0PRLnVddg4j69K9nIX+74JRs1hV8O0w
tKgEWGU8eGJubEMhsZ0yUKouX+tEksmQJM+kmW2jh+/II+0SwffMotQ3qvdUUNTQ
09J5SYJEcDKAszBSwnC2rwgKB68ikO2UNhtjRStvjMs2wGFgxGX3JNhCkMU6v6bc
NCKPYGU38P8smk0jHFgbsMLip7dqnK/482tRYAsM7YWXvK5ArSS3v9oefUhEZKiJ
8tG7QWMAqgzJUPIeAvtJI22SgU/xX6qf7GnuD0ixPOpfWpo9DkLA9v0xp3wdKcB3
mKs/nnc8Dozn0TxdaBTlxB0RYQVW0TyFYufuFt0EGYFAabhZOfoXBgoNCZX5UGE4
6LWQKbK0rAZemTccxTBhyThAl/q3FCydtQNAUrypp0bHtKLH/WnRMItOuO8KZKhx
0b+lKmAczts9Ra8yfQaWrMLTj0cPZ05Lx3LRBeSOxgVGoBsRUac22po6KKzx+VAa
Vp+qB1bhPrp4SWNh0Tlw3QrLrdLBrU7eIaZvgwNYi703V66XfIlIgJKvujj0jDqM
ua0lq2l1vl66kK+wLbUoJVTGSY3zJA8WNaHGPJ7Kv0xSOoDwAH6gNkNdaNRfKU5s
ta7em/m/BY0b2xtvcawrZ4Kf2FlMtfoDk9/AuyAf3skk0p7snwYo3i+Q8EkNYvL6
UaONbpZsBn8YuLIVrBY+YBL5LC8CGRyoSh2R5FNO158bY2lfWr5jHaxqR0qJ8qSp
GhKTWHjZ9nNvIeymDs2DO5ERhh03rBsD8mZ4yw5Jx0+6WBYR5PJZA2+CzDqlyunR
FINkOy6qIFrpvGyjqQY6kq+Pnv09SVFXC9ZXaTNNmMTP/2Ucjn8UmZpB2MbDmxxj
xbkBTDKt7jC1InC0speMrfHHFCp3lps6jHuKJtNM+ffu409CkeciUASvcOcuk8MD
40lpkDJr8LZpx3sQC9+8zixvXKkvt72Gs47roLKNWBWHNReA17RYr4dXsQNGWgsC
SbW0caJJNYXr/2URGFwvbAPJb/AmuJHs0Zwa2MXyFkUMd8EZ7RNnTWU1IVovgPW6
GZ7JOtCAsK5ZKntn4+7RfWbjFB1S9d7FqJnpmPjCViDcyvbeqPidSb8mJN767tSq
CnonQa7o6ESBxWi/19X/gxev3GjvH2kdnc3lrtBRmbpMEJd4BJCPpfAXHwRDnwf2
g7QOvcPMjcBtsDlsKXM0AMvdyBPPYY+Y4y452XVarNqznYl0NDvNCEnZGqkDKmMO
eF1Tfb3azzxozURu+OJIhvL7CkWrtSXgEuwlSD7mqN3kDdXh6NgoJxZ8lThHxfKc
Uji0ehQYSRnGhALMxvbyKgecZoBDIkmOB8v53Aiu1kfErwDG8DgtC75fl0mELC62
lAqYE3V+qOkwvxXtebBvbcB9DgWx6OOgBdS7QO2SYGaVHfF/PZeZ23KMfZdDNC18
aNhly84MV9G5Td8AarVk8ZskD+VC7nsiTFalu47dli/vzgYoid/P2RcxW5cUftB5
6le36Wr7GmZYO5GNMFWeJX4SWTK1chXu5ykMWXkT8EoKY5Kwapqe+Os7GV4jDTtI
aPWUkmTbEla+q8ohMAx/dEyFykeuZD4VlkKfDnTq8B6IiN+GZT+cDSlRVyjgw9BN
Wm0uGKuvlKiylwfCsemc+CV79MvpcJ1LLtXFNv0oqE9kJYvfsQeJQjZhSoXRmvmo
kJ/We4qm3RM4MAb9zf0S/GCrFySEc4+Zm78ygYHU4FGpMbC0wMiAdObuIrEaWbuE
xPB1uUHoOkoEVUGOUM4np0IHpOCKtLMPMSE9ZLrBFkVpBb+LJ7ntLQ3ZsewiO1Uw
yEXP6HLM91bRpzjlgwbDi+zVKAu45xydoN+Az9cShJlEii0HxrOMU/6H5497COrf
h3OzU7vXU1FxCfGPXk/iTrN/RgI/q8W7laTtpGnoXd3qZMcF86Y7I3+dMlvpac3Q
oDBUq8Co8xVbANRLCyXe6NLYEKVGvMJv/saIJ28Xrj3+kiXB/Vo2NGaj/1DkSYcb
HaaXeDUcAYt7UBeDFiD32gzKp0ntQSlGu7gcIWSJanLKBFSV9pfFxpzcpNUDjMFu
U65n9wsONC8Nk3pZ87GIsbrubtU8+1hvbrC9bb/n1gyLMffbMaM5MT9JO/q1oEoN
KDI+tE5sqpQ7vsJNgasxzf8SgPHlJbBUEJ6j9+AM6NHcAx134oP0T9ihBYUdR17y
XtA3SAxPC6pqy4vAoCQTcDYM69/V6wugkel3NNMVvZ6H1uC+O3tCl6NV13Min0YR
9cU9P6hbxNTsRnyCaaLDr+dUTobQTR9M6yFkTuhhEt/YWQ3FP3Q88sehwOh+9lFJ
6eylCoMBpnil9CTjvBdYgePQ1uEjJ70zen+j4lCwIcmWrCKwtY0s9JaKJuQSSfLW
kZxt3AC8T2aSl1w2nuc3BCaVFBeUteJBbED7ClU7EPStTMH7lFD48QH6yBr7KPfJ
ooisRac8gkY4kmpzWh80FZVXNXb2zVcBjW3tfV4OW/JOkSnhSAqlkigI8kRxb/3s
+mD6bKkVMrofjnh6yrdGV83cDPxvZxFg3rP2WBPq34BqyjRzZDjAD4RFp4Y1VXeE
LLdClwVtdQ8xselKJkjTQAzDt/kg7gis0Dj0vPv+C+bbMwd5Rxsp4+bWMT3m4M4X
pmaeqAo8oYuChjd1vDahshXxD4QaWSclA1twpAu6eTHMes4AHVzZFzJHdvHSs4gn
XtyMPRltfLPpuQRlhR9bWtnwpe1NhGh5Z3UA5wfUArbn+N0gWnEBfgujHaIL4NL+
DQ/YWQW3DauO3rNhGRdG+i9fF23IvrKJQZDNGuHbJuAkhoHWFDRWtFdugiV9kzbY
IKPerbAV3HO0j/Wh1aHhJLhT7KCmFznPZ7ufPSrIAJGAfFMeO+piH1fHRbIT6giB
1u5iIP9eW9TJv4ycYinKMp/BPBSODIWAD2W8jpur1ytUl6JTregyp2HuvzmLbQ13
tprkk2zD4089cUAG7bW9uAXViPuDFkgWlOhbJwM23sDdQnhetijEgLJnLX1UhwqV
YlRSKX4QXmk+T/agvyIo2mKayRE3oUlGUzCYY9rXG79+3NV2IVbwRSjsDVwla3GG
aN2tGhD1q04go+l0ry7OtPw+WL2A9YTz/Y9hw3snI50epjgs6SCc8p1WCOO2qivn
ai2ZeA15Zv9An4DbZPTKJq24EHQBl1+guK9hqV0vFT66uRzQ2Li2Zu8/Tev/2l9z
+duXATDVsue7buUKjzefT+J8bCWbpDCiaYbnOZZCdqzxP37tkFuCJZCCFCec0OHg
sohDzIaVGqiVRZrpV9o6CVctJ99Tt9hSjJfwv/lqeZZMADUDWS5QGYY4YB3JTO60
OBOgKMOu3O62UEbuHdOf05BS0J9tAhIuCdsjdECMXgXRpzE+T+DRZpK6zPTG1Xv3
VGN8QQSORLwRxnLprK+VZLz58HKJ63NO/xatGTe/KYZdxnaSPWwgSbw5F31LsU5d
U87iJBeRVgu51ABKNOwC+IktADewvzd218HztmwO/T6RAmPCuO3JRsdP0CNPKwBE
HCYf99PxxzPMeVQ6AA5l8alubv6IbRVDpHPdmeV3sFAOxp6ke5GzAmqkEwMTvc7g
rAPcYizdGh1aL9HMQgBInrhED2YV7Wvw1GAsezvOEq2p1YcZTdMClBFGz4BCc5Zl
GhrGmpXy06nY6DQlaQVOoq9rHl43SU8rwr0BZGL+dQmIqMlNTADLD5UjHr/0Riqj
2iyCtWv90RbgQ8PIeDWz/uT/c/xhXoS6gw5YYUYAFuYr71vXOzVny0cKWQO0TK4i
rcHwP6HLuxTuIobNYElL1W6QCH7rX3SHPoRI2xE5ITOeefdbQffQWpHkpfBxSZ4t
D2XvzAiE8Q6SPCJC5fSyUUj+nd2E0zlJJAGu5410uqWJDQsOtwXuiNCv+EAFeEH7
/vTHII6qc83+MW851LTCCrdi3lvd++ZtmZKKK7hp9IzQzOZxpSpN/pSclDvhwzSV
t5jJAt88+8+hiU4cxWMBFlItJEC0rulQB3TZcUQrc3uyN20JZyFDX1Wr+cowF0r8
gPxa2M8IHhn3DdEEJZ2wFjecGD6opo6yjNO+M0yO0eCJEAhdrslyJKkS6QOW1quy
yLHw2avotwDbiQ4TDRZIWoZNyZxtj9pr6ra1cKR8U6jk6oZdtj0jbp2LQnjYEGgj
RUcLRnwehVQ11Ng6S/8R5fbU71k0xaI9Uq1KB39xVgx0JpKmZEVw/2NcoRRi0ief
ZPWPBMjvXwSUXDzmVB6MknD7Ohx3YzvdQbs2x+YEJmFb9mVR/FHf/aabAwJkpjEO
Pilvyr5DGqUonigSUL3Kb6weKSub7xETCPg4jPhN2d57k6zGlNuoFnVUhTWmxJJc
Lnza40ELmFdt6iOT1KccD6/rf10NzB69iP8SiNDhDB7ZzUdwdkS5CaUANlFYQr8s
PH/bMDFVX36SHPXdC76Gcjf8KdVcv7JGK9ZSJUURJeMCbsFyAWq4mt6CAXtPnrKe
2YpZeaqXsSvnO6P20sC/NUDpxX21bMCVwaFsCl2DHAoN1svS66xXasK6HFHXUPX1
uL58PAkOJ7Bujzr5AOKFktUgIl/cH7OaMh0JPN9ra2/+jlQwBTtcpFnXZvRibbWd
pVcLe0VSGnCaSajr7+OvQDh4kR+nsU5bGnbzyThtfIVCmeymueZ9htAbNRVKWaPH
YAbdTwZYKXBr734SAY7dFQ/vythluC9mNPamDyYPQuMyOV/H/prbnpqTKPSuxo9o
1cBjMN2Xurew5K2JTsKQ+aTq0fiCgnNP2sSYui9hKReLpzBGx69UMs/pwCS0nUNg
WZ4X9VvzwiMC2bfkNrwNLcSQCIEoMOoCbOlWzxAp39pyMfGx+sSikBg1/MFcl6fN
1gFthpeg6XTE+nhU+0zsCyoObWwjl/D+8UvfDEiGIXouNR7rdoAgheag0K5DrS12
6C6zhbKVd91Z1kdywX6HVaIcaXUpYyzB73Ct3qNoTJGG0SrUStDMBTn0k6S+DUHq
csU35HQ1xHR2avdoEx2E5iOINFWMQm0LIrnoa7o7xQyWmnNs69HVcMf7t4XaMBJa
93TxMPVvjzExdYrU0apNyIObr9a0P8c8ErdUsoF33E7HsWlqpnByAmkzn8+hVvmi
FY/W3YzwuukTrRduvKypoUC1+Ay/C0a+zaACWKVwib1ndKJSmTYeCKPIBJ8FJWqH
Sd7+iWDGWzmuuedE+YLD6pqB8sZN97wRQe7W6KMcICeK0NjsFYNDq7X4Rl5QmTa6
Ylpvf/g8fnIzDbJTdhCdx2h55UdVFUTyVhWYzgHmaM+3zkpnDcPywLxeADhwnAff
2bIFLvVe/Eoog19Aj62GBdkYIX8BrmuN4/TTTqIQLhxlm/sMDqpXEAKkDzks5y/w
UmWsw1DSTQYmPoEERgioIjnWE23FCr2An8kdtEuaXwR727LcPHnSlkKaJB5PkQgE
anLmXy+JwbeuaxHP/XpUBxPR3NsmwxE1D3cw6x0Y7YnFTtH1z/DoFTeI8hpKIRdy
edjZT1I+gmUhRnWakjJ+Pnf202Q+r11AahLthrHFUEFzYZ4Cg/MKaFf6iZGMeQY9
BJXhrQ21FiFJ+ZPvhJkOyYSUyJntqP8Qh2eIrHMWcRTItReMPe2gVZ/98hiN2oVZ
5iazxieIgEYlsighvzdTU0qg2+YxNhA5dZ/W2g5XYbyEvDN0cf8F7PREw/er/Svb
IvYIrabejJ3SIRMvPXX//3XvLw0aXL7XsopLnypUKQXSUkpURKcv3jj/pcQJLnaN
gVLG1tCWZo9oBeRSEqq0zmMMh+w9BzW9kPngdfE85ZmIhfK2whMY64k8U37JIOzJ
a9422/qiBGdvja33tDhiIPWGkdFRpwTXOgx9Kym468oLx5ftl1rL+KXb+nYj43lo
Fse2s/Icywsn9gYGe6J9SC4D2Uck7COL4AvvS58T12TL//pN4nQuVR6046nJh7bI
sVuFBGQCnBClKubVB29OLTO0EwPdgc55G4JDzrDZB7zvhh6PJO35gqyDYlzYpOqR
V10IvL1P5D/rxpNSfQ14d8z45PDHrk1TFjJZrdceW2JjAxWu0XNwaDC4gfNki6u+
FtkCx2NKVrmBGwbOoYDuClfK8hlqNIC0dsl6GiwB0DKoYHPEfMtiKK6rrD7608YD
UoN8SawttlRVCbgGNs8JkEhtSKAITWns9zx56GLN48Yu/mdlBcGZyQMXUikkvyvn
p3u8Rbk66mcpZeJeqbvXgnX7aWGOGQwuojd05SW2Fma3BG6zQhL/mpxcGckeUt/R
PuoMkTYq8kxNwAJVlrtRHzX704IJIIdpnOD2EFyVU+shzLla1NhRUkHZfJA2urg8
wH56VA8oUqF6C2KUBYVd4j/iTLovf+dGMLDkNb/JBFIvbz4Pvrvbp59836VpavSU
UVKXUefFdNlF4nzY1k1GqaDCvJ6fQs0wlz+v4bLBChxLzOXBusk9AwUm+FBBCZPf
6rg+cCzSK6wAyWw8Cp8kmioo2SkD513RK42x+ai4FPu59+WLtTSX3NyLshVqZtne
NiU0CmvOJKFJ3M7jtIcRGbjLFe+IhjMWqrr+IHktTc2GjvZZ2PMmJP564PmuMJ2u
uu74Fprj23wrQx4sg2Oup/r6D77hCRblCKZeI2ENuAWlEpzUvEbu9p6/srVhK1Rq
TwiCxygzTDRm9mY67//BKL9+ltZZyHZoq3wTSKaj/zGV5XQl2DIBN/J+lxkRAolu
u+DRq/NrE7GCcocS719GQ76PEtimXm9DJUHtb8I80Wy5s9oKaTyi2p/PQpJCi1qz
LNadNLip1tdS/3u0lPqhEsNpiRSZ2pR3qZulMM1TdVBUseeJqdBJYI+ymEynryj/
zfpoeWvqy1Vxo6np5ZyqqhdbdehW/bSJooECutZ9y8mBSn0sts5kTVZN7faC3pdo
AF0hC4akBJt0ZWIjt7d74133MhRDUetQWrcgnZyaViQ1rKSN4+NL63sM35B6SpMo
EYAPPdq0TtpExYHh2Zkmh0/XF8ml24Bi0+ftHAN2CZWMhlZ/ImUZcPyCgzdKWv8U
TkZuNmHmjH8MQagoZQJC9x+YmNthqccr2qc6bLVqJj45gvSRumI7SHmcsq4bYxfW
itxqLZUdZwyX6Bq0zimG4Hhk5TQV3/8okSqmh3uiE45RmURYlU7FWo29j1YIZ9pC
StUCp6Q9T3JR8JJWFN9wVs1yrCtlOCzqwV3N1Z0WSbYpH5DP8nXycL5cRYZk/1fJ
iF5Yx1OgWVOBdPO7hNS0bIwYmeqfFifDefGsNTwPToub0UluDvsPL68Eoam8VZ6k
NGQjNXmeH3jxaIpBf3/POiQNsBn7Rvd07hL6h6PpBejZvCjaQJec2OQEV8XtCQ0W
teWZTdsu0sQkmh8AQr6hyAPfmL29IQyBWhVlah0DVcazB7eHvm6U5mo0hn2oJ3mA
MDtH14bD8r78uR6o4MJKEfASAp94noM5USz4Z6yjLNnVEbbl7JkhfaH0QYsvGY5b
9rlWfY9I5xEM+xwgPTnnbyQDGQ5lpCmGJjYceEgXKKjm+kUYglu41rHFAB0ZStxH
sVUiYXRxLNMFGdqqyj60bq9NPXRc3BGQO0jUoNWlU/i5r8xQtJsXwclasb2zRmbQ
VqOxTajobMIG6I65Z2o/H53ugPNiujVuuqp8vQkKAH8ziY2NsIkDElK5rXlwtpFi
jjauOSF/v3SbTgLaYgNXFj0Qc/z7yCefRUrchJdFoVru1URa/KMQm0xOCJ2AbTZh
RX25fMoYtPj2PI6ZlYzLQJxEmCWSxM4GefPvufaK+c0sLl4SrwD/hj5pQH6TF/ls
6fNEDd5QryGulg32d3aqpIxF4h6cLnFFxn0vzK9dD0hdHe1/4iuE69gnC8DY1TNF
aDopgoMJHb2GAtIso90ozN6S0fk/ISnHQNT/N73yRweoBW4iNRKUAk16ewIyTpcg
kQWFBNLIPdx+SpsSnN5IkXsgTvXUSSZRASvY90FoNdZNBKw9m0CGLWw/KMegQiCu
tPzRfZ0kyT06VX2mzek5P2P+hE80qIIqmj+VW21+Nf4H54PNzr88ObC+bzclc7lH
oU8Onq8sbr8qc6RNQIeTS+3X+pkn1QYueZ0NJPWOLLuRmPkmwJBlC1gsZh0qJefm
arQWUFWfIeMjH8ZomWMIOdgUexs/jIwePUfUO5uEOOlkDrdXyA4Ywf1hYHpdi2p/
Ctw4mDvYydhpEtrZt/dRZI3M59LH6SYYINjUVOmvep4W+Xl4S6KdwS8EeDnyaIZ2
jSqjK52gKkGi42s5K660ew7hkbtra3lLmO+TITMaUWpZL8w9MixwkqEMtEtlC0xf
r9luYFWBSZQw+iU5CCjCkNcif8kJ6a/b6SzvRwuyWOzEgJCf5ye6MGTzkcVh2BGO
ZnYetvpsIzFU1leTJFRIXDVYjxvvUg4z5SHzTqKSx9PMg2Z1Ow+299z0DSYSWfC6
uJ3syJp4QipQrMusy3QUcctoR4KoIaXQpTSTb8HDLB6VAc/5HkhZ/+cq2PowG9Ng
Mz+z/dbUM6dNR9K2ESmVHEShXvXKNiF1GEWi1rbCo04q3xqSgOi/JAVfh6embbnj
XxFc4D1L1OMo8lecIFk5R6iikS0Q8o/PtP+BZ6ZaNJ2LPf00TTqoYlQc5Wma2ldd
ADxSs+VkDHrAurY1bRFTPKB6euIq/2l5msUljtyaujlR5GgBNoAPWRJ7ISwpu3Cc
g0ujBWR0mN/ed+ndJD4+I0urB5NnZek7dFlRx1BIUPeA65GS8Inz1FeroACtN4mT
APf6jf9dj4jSGmWPx1iMXe90+3YY/IxRmI2IZM1aQ33ca/6c74M3tK7UDJM6ejm5
cw8KxsY8wRDwCnNLeb7sgRlsPELIH2pGE9nq834jdTrXzON97qYQI8WzuXyMaVB8
loS2duYZu5Yc6yzwe0O2a8D+Jj0ewCNiDeWg+zlxIWSKwf/SmyBfaEwKa+iAPkSE
ol5yvg3t90j0YNbuP0kXWYQI36oGpWn8fKcnLbU4oHeQW+MpxI5EF+mbyJzOihix
hcbo+kO2XtGeZbKyiZ5ORZDnd+GjnLgG3SYJA4lvFJe/EaNelG92N10bJfmfmM2Z
wcAVuIXcG/zMrxVzRdDS8WBWM5shGt77G7R1mgK3o+xWQeSF6ia/kTHONN63acWa
6lzdiOZPb3jCGncHZy+nEImjmfC8Ssg+SNkVZ9E5ApVg1tff/lQpl8atHxlE5SRh
UstQgfCTRuYKGv7h56z58hlGC/6WaL6+OxSlW/JdzZd+Kczx3bP6P4KW9cJcOG01
O7cFP4N31xqpS3XlEhtnNmKAoTv+biokm3L1zaoHRC31ZjrM1MolOG8NE7xcMH8e
OwsebQPy3Y3ol5yfCkRFbMJTnwtm6t8UOFvNeJnSEtB+beTy2ezUymrReeqvaz0K
rFzP0MAT6kuSeQM+kxKGs3eAsDZ3Xt3t15+NTNBSQpHsbWVJYmDc7V0F5oNVn3y9
58HiW7GIiuFVvsTC1AQnMIAQATcHcp81TDdxPsf71/etxbLZBKa11RKxxmCo9tjm
LS+JaTEOOI/6MfQRFw/mlB9AKGHJpBlvcHXAVQBSr649gwPN/5bTLz8Zbe9Omk7I
GhPvTKhxau5BJyDTC/MeB9DGdAM6M8WMsytLFlQYiEsH5CO+4SIxFxbYN27/jQEg
jQwM2grd1cFcq9iy5mUV03Jk8jGBN/IgU/apnTmdX/vXkrn9DC/wpooOOEu5n8Af
5j9GtRo8Y90Jz8E7qEHiZ0KBFUxaIwtbx56IBMUpMJm1xTZoegWSlIaXV/YQpC+f
vssFURje8mZfmRP47ai0kcD28dV4dateHHNG5sAtQwbf3Ly2rD4EEIkO5NdMMpxz
Qk9+pMN1Gd9pQ4PdGsY0GppPaCoWOFwWT18JVpWckWqh8XyIW5KYnLzdPmE038XB
QPBdxWMrc0H9axCOjCP06c/HEDe25/0fdRlCSxd+na++ymeqc+UI1ugVQbmDh7kH
5eKXiqtYCH7/gD+paTxCyancRedF8WW1VZJErRK34Dr3Kssiab7fcVzWS6dqsRcT
6CSqeVv5tdw0pE5DhKJlYgkOqea5M36Komiq3kzYtVBt9BY5kk8cfyiA/ZX2w6jb
s0wIl3yNmHRI3aV1gcT8ENytM1gpwOH/hgyQ+y621zB5rBi5l/b8InznW4DW2Z+6
GAx4ZTXq5OyUYF5YUWskkf3EQI+dRFMWG4o7uBNwjzCvsViGmEk7UQaDqOlgqpMr
X2l6tza9q0d88LIKhaFeDVZ5KQvZ7dIgOSUMxhkXTVJ2Ues8qhiNzqr1kwLES5T1
EedhgU07YoL3DaWLCQHmWg9a/KQQW/SV5xB3w+JHZmLn7tEc4NJhS9FKAXCK1nsc
WKo1aIW5hqUSp9DSrRFLekUwCCgQK9dN33JBN6rwVAJswwO+zT4qppaXP1Z8XVd2
Q7Q5fP471PqXcBuhl7/6l8MCG25cXqakyjzNCIyYRTLKzguNM0AMv1g/YeDxzpX2
XVt9wr/Cktx1Cg3UziDy9AhkblwjVn9tOkhThEzUcQACgxaiUmJpb1ceCMLUa24b
zZT++wDP7tgA5q8jmSSnU2pOBSTkLm6ywAm/aWpsI8eCfYHu+SYBh173b+s8UuBp
cBH+2x3DCErKpKRpS9gRTfU0AyK38xCJZfxExILE7/gLSPhHP6EoItIWB8Hpxzic
m92DI0AjDMaPOwTpmsJSvArfavZrN6Ci21W9wjjaxDN9PAQtLKxp1WXF6cAiWX6r
axX32Vk7KeD3As+hu4/J9PhL5D07y+vqTyu+stb+VAU3XyA2upK0LeJOToX4enSc
1g8htH6nqcMhZ9MIp0xIp+bcngwAYOhi4BjtWNNkGxqUuvzNJVlmTqpK4PoHyOQR
imTxf1bbELvoOlaIuPQpqM+1t+2agGWwWqQXsP1ugs7WTqGwyH4JXjVmZlXZ9sAy
sNaK86ufK559ehUcXZGLbcZ21ZPSmRR1xwFi1h9A0uGynnHRGgmQ0abmOJnkT+xk
XyNYRdDZHmtVj3RbPjeyMpx6YykDFWG0a+HUpZJmpiVKTtiggKTz6B++GcXUhlPw
tprp3vwt+KXzl+NzTl9liLjY8ovxcTSPdD1Klqj2+qRDii/Gu88vcsjdt7Zk76vp
JwCrnD+HVcr0SFQv4xy9uHs+O9Lfjqtps1CwYJ4oqamXzFdxs17J7WR7VeYLpcbW
BN5WRPk6UWZ/PHkQam9RrF6JUPgFU8w9vfa+55GGeAAZRKTCNwEZPuwnW+yQ4RSw
GXuP2o4hmAFo+i67zQFdiGmD7FlBUbJqirZSQyts1xj1QwU4znNFLIu0OtUN8NqV
CwtzsuVYSuTXEk5i0cQuw5r6/WgMGbTyiG+AFxKPvGuOtkkXbHxHNapP2FcvQMPj
/Z0Hb6/ysPIhTJhYl+5oI/GQi80pzQgmL+WWZP70Z8dfV/+RyEBkV6IRNUctkpz0
F7s9vKqzTuQjomMMxjIDbrCo8MaLAYqdNwS5pruAV9D1bgMPRr7ou+0I7E/gi1l+
T4OdhL1zqiskWtXaUVQ2LjoJzmhAU5QOnjUmGdx/ZpYS/uRSB9pMdQWOWsp6ZD5H
KtQZP3DL20WqGdZAKdKWFOs5LOwcSOf8QKaGUTCEXC4Ymh0zyZ7oZUAtwrnqdN0X
yRJTLhH9l2yIPdq7FWd5zZjk3G3M8e1TEL8Yd7SxN7LGFlGeW4ovsys+eDWsyIbs
eFW0QJRY00kZ1NwfQTOsAPOfSvS0Tsa1vd49KWM33cYqadSoWnka4xpqtbpUHg/l
xNxocGPFv/XoMFFOTIxr3R7Fxb1LMmRA690H3WsEXKaWixQzbim0tJQxf19YnDI7
hCv+FGduatXm0zjDiRVoZkpxiEKPjacykqD5UuoLd1I2Y8KvmDBoW0fduVq5DMZH
9KCCyNFhQ3HasoIeH+KhwUyemqX985vcFjG/Gu2EtZMu/4DNbupeo+UGgr93Yhbl
6em+UoZGfFqXNlPQdcprfjvpYmhcczaf2NvXu1+d35BegXOhyY12iw01pE+25Iym
yxMFq383+2JCE2deQ8XB+BOh2tfYAF/IVtfb31GaFuG1j0CucAQiKcx3QRXw27ci
xoGQPaaJtdScy4lOSfpS81Te1g3NaOb5CFOvLh8kA+aWBrIqG/N9TScRt22AqRo3
IiW43Jl01Y1e8T/Uhy6K1SNa+SJqSJCEYw2xcMaCnw6BELaIJ+jHiynUDsOtpSLC
MJtpfG8qtVTo5gO+TYNWScfyJk85EO9XGycDwjlml/TuCM7ZJpREWQ7v/tOMS6N3
NRhRjuDzoLky+9RxE8G95s9PKWJf7+9G4aWY/cmQrj7ycLcR50+mdmCU9ibXAxPD
uPMlUcWJup4hvYjr+OZDfXay/tlFeG1axv2PpmNfaHi+pD3YGNh2O5jnIJj1IcGr
YQfFtcV/8rqKxDANK45rPSFL8943OzVQjhZG1bBRBvgfpw0Chb3/UhhIIlu9SQNZ
w7GZtI9WHRdFgpc9SRHorxIn8LEc94usF0qR5nIYzndY1z/StepbJR+jqC3rAzil
eWTbFmj2Z4UPSlo6hJUvegNwNf2Xyfds458XMEz3Z/nrdpYw1Ru656z4fchmZj+C
K1F8q39q+rvbAiwPynPJTfH1BtoefaduxC5NXL4nDecXCGNHMwsmn0p3TmHpfh0I
4aevjsFj9fIJ9e/p9YB9X1J6HBlkUh0RdXDR4mweOt2EXUy4+kHpTGKyBUSne1vE
vxyjoQ7ImG48+Wr5rR5LIjvNLj/3n4KYN/mY4wtI9t1QAA5Yilgx2+rTOC9C9lYq
msdBPJE0vJkgI4ZO2ruXSxpvlulbd65AcetYKOmd1ElwT4Q384TV2bUqJFV4JS/7
ExB0vipRne/UcYBXY2zTnT6ZjEvITEH7/Lb7aRh0kSFXhXFPK8N3HDAOpc850Jlm
UteahtaQ6Dp0N+69+t8YRa48nODdANheIpNoV5GPUPVhbe8L3N+mK8HAH8OZAHhj
faW8jhD7rILzUSVpLwp5dHdpkxQn9H94EVZsmsvuDtj6pkkN+0yFBpZmRxakCpyD
arak9xcj8+4Bb+2qdauLhqtC5XWi40cHGxkF5ebjMtxmtlbehKxsXm2jSoufHWv0
ss937otcTIL5rxLO6zKtuwN9/FfXajGl7gAfEZsxaGKVHF85ZHkGyZTSXI1jHO54
PF9EkiZErK31kX8zJC1kYtFv60KIMJnOV2pb94oOkKXbfejQ/VDYgctam5MFA3Dw
TLLez0dO9ShseU0umCzj0QsUz/GWH8ruy9PWb3MvUTJaLvHkVPB4FQhRpItQOuaW
yCdBR3k22vdiFIagJTkKEuEmu1a32mmXEk6CycInyjs5x2o3vZNwrY2oG6H14UqF
xaahLVqoiHlV921yX9RaGhtOYwD4Ds2Ju5BLNlucyDE9GAHaBHrS+X2EURgUx49Z
vTKZF1V5fUvUfMWbkTveUkLgIXC88/oz60MYX8XSnMGV+cqMyjMj8S+o5pA4Bk6o
EXNu79iNHYtd5nqrNe7K8o2JFwUFRSWVNs6nrrGxHWUYgtVIxZ2LwTQ10RMH5G35
GK8HR4kJnUKMs+6emgLGacybFyafCMSxUAFEWLlee8+k62rVODmsB4TaWI2lkbTg
hK8CXx7duPoaOQ0RV2mqNQTJhHyxdwPlMe/VHIMcCrebclPB2b0y7Ys6lsxPaXhm
1xR81MmXxOpV9MYh2CqxES1s4JHLTSnWfsce49mqk47Y8w87j8IXUcm1ya/M7IXI
fvverkvpJakhStLhvAEPQWNvwwx8R4BqWJLPoWZdMocsev8DuoSWrFh7DFUM77XI
j+0VzduCzeUuFtG390NHrqSsTeuatYDEldHGiUuTOQzUMxKvv/7ndU8y0JkN4RBz
oQZ0vBxTRPdf6HOpCKvAvDWTuP4sBA1eCjbHvuaTJFfuGCLlhQ30O/tdWIpbCnwb
zzru+Q28LcNYF+xYDj0EUJg2cxD2pKlIESrt4qFu5GDnKy1rlfPw7SYwV22hq1LL
zddKq0tXWRXJo1ElLLDdni+0nHYnU9NkiNjHL6yEiwxItlBZonyCxXslinNO8+Ag
UW6zA9IiRhKwmT4PHv3HYaOlIadWNtbE/5XdTmLDzp54q+vtRnxl92n4mG3+Zf0y
ALcQLhUazWVL8hmt9FmXj2bmtjY0wQ+TKSQ8E8wQCGD6r2tBvpeW5iTEXVujoVVL
MPl12Gn7BR8hO1qKn7wtbJsdGMIJBhJ/geYIGmqjtFBeDbZR48OOmBeECE/QeOOA
Nd/lX7gQ05oEYB+Vs3wzPw/lCXZFWeV+NZq2Wk+QnXKwYaFO7jhyCjvPjB9Dz4RI
uBdESWeJa41acvd8NmUBTiFtW0ZnCXajHe46XLx0VNlyOeaGAa81xqQpm4Qjq7xU
77KlKG1NrZc0NCxp+irDLI+tAFN+ywqd6JVVKfGz03Bs/cEWsK0kfWgXdZBBKq+f
N/5A4+e4Ts2pljxi4bdjDlxnAFnfu+demYEbrf8TXNukgGxHaEmQYL1RsuRp0iHj
DQaQKMby9+Sc9AYVgOyRhM057jeFnWQMK9pwwr8GoOxNd+V17gKzy7IyW/CNdtjn
SBIHRnwYzD6sK0IeXv2C/GTiCAMe5zrkjOlECMMp1OZCz1uD0mUcBnWap/W44RAP
aQZsD0juxN5cj2vePSwJMG89cBe3A3StMlWbvJtdRRomrKgltovUUO0h7knwOomj
5efqhOE2+ejVL7lmjzVmN0v6yVD0rFulycF2TYksdEfl1UytlRN8KhF3Y03nRufv
W2tj5Yyg0BQ4u6q55Ksds3+m/D9zHvGgxms52su08ntwOtaS3wceM/x8yYvyPFp+
+0fqhZISi6NA0mJXAQ0xaHGCQcgcefPY8jhpjCFofDqpLMwJ2XSgJPs9b0ZRU6Zv
vlRFaLF8+cnOoIQ3PHfnYmyZaZieHwNKrZtSPVnHG/zm7bMequAJl2roDmXIzt7o
c4wgqS2CxFlo20YZoHYqLB1HTQKzCQ1orjfQPjo0qSHwEGOh0lm/zSOVamEBFg4k
a8Rehv4p36jYxRjKGxx/dxt0jaWLXe4q2WUpiot7tpwUpl5wpp/6BfcR4IfRUPhN
0dD6gFrpHtMMtzdzK5HQWO/jIHX0fvMyt6vBsw8ZfxqLe0wFY09tnf+vCfkIW4Q+
NDoT6xoGVq/sE3WdFpjw58peCXpeeqZn6lQIPtwdmgOeiV6sIU/3T2mcPZ0Un2bC
s3H3Z+r482//i+UpWo6eErjFoP8rjD31j8pxjzrKn9S81IjlzZQ6rIlc/lSFKQTR
NjMxGCv1fIp/DKnoLVjVHQXCA87A1iABzn79cXs+QEzN0WqAF4UZV7Wpgm4NgO5E
vYH/otWM295GN3lOIwre+Q8k44swdZ5WPib6KBAOLy1mpA3/rtJRnrBiW6MWWasg
nJOOC1HmCW3dxSaSJUZFFwSgpyWB+0ZV7V7pxbp9G6X4QPWdowqIBOl9tG6wyQmE
yw/SqvFdqYcCCxiLKfJ6ggzJjqe42HZifey+QrB+Y0HJ4cuhfOBCTcxgBgdHnG/2
fSrMeMTSSuV1r9wv/L98iH4N4bwSBYWNq79x8iqRcouN2ZeE36gEUCNVpHpRIpwa
12pChJwQ1kldoKVTkHa9b6NEKFO3LFuFORJIInTq3va7M7VlN+w2z8EaBcoHwFtL
vOavHDzJjrCSY8OQW4NYON/Xb5mbtkd3c2UzGv02A2KQn0dQUW+X7V995nA1S8sJ
t+WcxQ+wvofmDtZXeEqctF1QOCEUTBPaHvphfxJGHT8V/ZEPsXlo8PQalYj5aoap
Y9ZEiLnA4vWJdkSwzY+p2y+Nvky5INGSbr4nmJu4VmJHNA5ViJ/Kr0lwSDPwzd+p
vwsxVkHopbFQ5sGb8fRK6X0S7VUesCpqf+yiLGrXSVS/aUbHn4Wlt6E7tIzJ5Vxr
ZF8xLKxDqhKP2i4tETVz1zhHW3TMCs+2NQgyiaOrijLBVHQvU/K/kSZV75ZTyCjN
0CACvYFCij4xb7Vxx+ttHIhdhX+1sR4jGsoTSFRIurFTQiJkwmsNNARrZfkYg7mp
ZkZEahTsydlR9LymicoPBsdpG+NE8Pqn5CVBz/d2eHjvhuCQDpOBHLuyD7CzvoC5
j42Opn7ihUtlABInh4iU18P5gmZFoDobCcQmB2AldbfEoSATvwsMMqFBx6sIs+k0
qZpFfDyDFvYwYZS+l8HSot8+u7T3z8ifK3izo8AF//tCdGNxiLcS0sFpKGyjnoRE
E3lNGoOkqRAb4m4EGkWOT5Gk6MRBr7nDDxAowQqxGgedFAd/ycs9m5f6PavCHZwK
e+ylIYxYtBZOyJtr63Cu8VvjyO+kR7wzrJVC6wfb7rC5FZa3ZjeWCVoVNcOAQXQy
UmkPAPZ4bcBJJcTAEN0QJLSGZPG0FcZeFn06nd+Fj3B81L4nv22dr2+x+a3mtnC+
nW5V93ZjWFSH2ItED563G5VrBZT+qLSPqQxE85m9UHx7fTvEm6gbzt0sd3ghYOWb
8v2aSxt1P17wEENqas9QJGQIW0s46HNDvvNyayry8yXYb0xlhpqRywyEe95f60Oh
ZyT5GtBP5rbcDlGitCBeJJgmGbdESyCCFwEW/IJq3dQx8Ovl+3mwt9vefqYkUQn1
8w4CYebAwV5tLfgffclUiUE2AySBSJKyKGWN+iqgNJBDS8W0L+oKTQO/B8t4gGvw
MwQrpoXBy/zOmtOuRPWry+ttUMh8DQ12uh5UtnmDo7m6i7YXSL/d6NVZb15c+NL0
eQnlcsKwoC8TMqaHC0NdHXzcPR4mSFEK72qAmRnsJY8+ZQ9PfpDU8wKyyecNY2qg
sqH8gNe2xFuJK95tEhWHnG6hd62QvGJjk2kyh0yw9wdOXMvimUy1ftN3soxBAHnP
Q75aaEuxT4FhEMH1B4Qc3WribHhW5Zo+diu4b1+7bo3KX+7R9p3D4ARQTiGtQNj3
FTS3D9JEzPNw3uR2v2VzakTWb1YdbBKkuV32wLnTvPdmER39mQn6Sqstbw4sgwh0
WwUxlvOJnQmrB2c8lceRTcC7+bQql+ToK96XN16A0rcgFfTdroCY2FW0ReNuWyO/
Z1N5cMwmIFVlbXR8+PAq7SIgb9K3fKMEq05uUEyPeR7dA23CJ98Pi12iGHV/aRm0
F9qZgF55ljHAUYxzAbLr/O5VygZ4UbX7aUKqBfe3BrGjHdwjyZFYjFLcptfulcNJ
Qk7BjyxrjU23mMwIUiaDVAAxIHfYUhdtdJH2cEswRId637BwZFoM/frZHb+7h0VZ
SWHbiSRrr4267AdQ1Fxpj/b3ZFPjAPsGXJMKJq3lQe9ZAM+degocngSjHUT9T08N
avmDdXwITjH1kkW+XhR3RqiBvbkn+lwtsWf23xEsHxUj0ibJpofYKAMgsEfsjQqu
9mdpcUns8pu54zNXQJBDK0XAfRsBoLb8hLs45964YSYQ34SOXtPMl3GNDKgq6Cpy
pBwogFRYUIXk8NFGFAcobhu1MJAqrGJq5TeC7PQYwS5YwAb0RW9QeZ97Qmxwa++O
cqL3ZXzuY0s2Ltko6wU5EbsvYxgLbx/3/Ce+XeI0bszsI0bNJ3BvF4k/6GY3D8Sb
uW4EY0k0BXUqvDTcuToocapotUroytjR+4ay+QsEolpuNmXwjKXasUQyfJmf271p
WV0tr17b6/VcpdFJCpDSDy+NRoSmabQCkfyDnIrVCGQ01QNbcEkwLbtkwhkJoOTf
7HzkWdAwXhyL9Se55PLWyEaNH+gujInwUzIq0osvmdI8HEm6xOwRIE+hDfUngxAz
IhO5Ujo5BSWFakyMiGJ9QBOhoSbRb3UQ5ihgwTWCV6WSZq2bqZnI2/kFYj/15SQx
Jd6orA/mpS2YEJZGj4zoMQHqWkXotFf4JeTOo10kfrkrM8A+Z/y6gVWy1nYvXGgV
ew9TfpgLmvvcRApBCr9OEndhjCnETUeSoox8qlXVZSl9TlVmMKEMZQavrnKUOcwD
ixMLwSinPyA8dtZPr3vlumzKG3Sim/3AZvC1ogFv66R75jzhMMqCis51Ss8iKiol
2Usq1thwcXqANk8d/HInFIJJUAI2dlqw1DwAO1Z4ogV5Hfd3Q6xrpxE4s3rIiGFn
c1pAm4dgGHzy+4OlB/U8Zt18G4tBnysaMoKoCUjBml61UNpLPbYVq8gGtpHSHKOh
i9jH+GMzuWpQIqBa5imz8xte7vYG3on2XWboAD07PD1+GP2SCUu337pDRac22p5P
LRym2OHJEix4a9hcPUPK0CALlS1Db7AKgMqTD3nr9hD0G5Y1AALZA8EroryEcwj/
oXVgzYofCsx3OC+oNKYsK89RRa0IBlakEgRqdcM3vgMlB6oDmWEA5Pc91GcQW656
Rj4vAjOsrgDVrFKj8oswXC3qAXbd3vMoMVfh1nHFZAmXPIedY3XmG4nxNyWD1OA8
6HdkHxTG5DXnrEX9EujT+A+0Qu/jLEkart9AsNlOdfVWXiwEZpRn6GyYujXHEZDS
3+rV5Uqi2cERG1vCUIh9b06/m50jiXtbPFKs6jnnHTOYFPv9A6NCKKpQXWIQlN8d
qAe6SzdH+YzyT86taNfylZAW/601sYeXAO+WqJSesb4dhGq8kD2XD/LN0aFMQP78
2f9AxmFGnocFRTe+B4K5gLNrs/keFETXXekkPHO3PEO/WqYewv24Luoibnr2JwKn
zo7n+FRsXmmpKWuUOUkeOWc12I+2SKh/yC1cxXkQqENF+TObbV0t7N0E+l+KkFAB
MFvrJR25Cgbtl/3zv9VbsDtMQpnJIYnFHf3R5Ye/BKTzYbR5fyBaxpARxE8x2hGo
mqpv9jxieKtrEW+uXwuvvEy77hqnZ0SDO8yzm7gCY3b78W0/iNT36xnz7vu70zWM
WknYQleez4B6+rZwetj6lXdjQ7mb/Z/+U0/q1H0GbQ/GLwzwYS5i3Klc/Xl43nRA
WSvMhgDKojoM6aUS3lJNlIll2BhRVw9njMVxB95YYhqy+7AsHRI/d5sTvnXlYIw1
Cri3yzwtrW7o+xxoMVlJCUQBknxXRlp1Y1NoeY/WhVx33PqhltDls65jiv6ayfEU
GKmrtpqBGRiWAX81tZLv2i/GYJN1iIZIu4ccG8n0jepxib9KAbfrBQb5+wL3hnTm
n/64h55JCdkV6xFtA+hH4NVpWZPARQRUgS6yOFU6178P/zqXktJzPqZaAl5eUxQ6
bDD92DYiy74L85fb4vYyGLUM47rX2nfCQ+V2y6WdAccdxWs+maXoJ9uhd4QbNUTg
YjX9lRvSz4MHpIt/SxxO+h2tbkBRTtBDgeGn6HLvh7D3B1Oc7VZIY0bxELDCqFIg
8rKm7xy64S8t3YgV8JSGevIz2bwUQgD3HiqvoahqHuzLZb+O2DCGun5Gu2Y7pnfE
SxUjFuQW1ZquW6mw8fNW/F7Jiu7Si0ZnKcpDKyX8ezzjceu5v02UtZWZ7bOa6+ua
9+0vew3mNaV+Fe7+KnvnXr8Vuu7D25y53twhVkfuvNad0obZDO5rKzmQvtXzq8E6
N5ok6r6Q2Ydvq4X+bwjHqyl3OF2N7XnhqaW+s3L6u1z5i4uH4UMR63Bu0184jY3p
QzPULGKNIG796J0QcZM+hlY8MbgL4fit6PqbZZwWy/XOfv0r1zcSxXmsa/lB2xkw
dqkNr3mpygw5mC6LQv3gVsSK2HEo3vge6ufJlJ6GnVSrKrSaxk2QyFdB1HmNlW1h
riOJJ/EQEBc7aKdLPwsXo+FTvLy9qoCa5ETxfCDp1hqrXTU8Ng2GkwINyHvc3jOQ
YXFcoh2AN+jCiGC9w2fpii8/Yvj68NkpSVLP6/ByB2Fw9agtdU35w2VeOilmAc/5
V1LiPCpN6kqxroWmFTT2IzLnVPNwIjU3mhNMvuphnJ/Y9vMDa25BZsAsSi7KXc+U
hjxKPk1YgAGCqvF6OO18QFtP9U6np8UczwZMgABSKxgLtOn9M34inPHUED8ewvWu
u1eyr5uoA52aTOmFEBXRUBxzCgft6NjPBcfyf/iksypcYDNIJNLWbKflGOrP2s6a
bN/vi7lXkZ3ZPTWzhvZ2eS2uLNRWTKBD3X77C/DKf7Mb+TzA3Ilvvnulkg7krS/Y
/rZoem5Z9Ut0abBb1Yda6sYsm/J8XgcuKfXSSbbgh7HsdZeXhM471kqAi6GO0K3h
uK8wIHS7IJ1lSXNbvXjeJfv9cLW5n4bpYJGsU2VT773BoTvxDnev41537NOsqvvP
8hIzP9vOE+jxBQ5h2PdejnE+aG6eCeO7k5VQStYka34QtU6IFjLnPydY/LHKS/dQ
YTycjPIbbloxycZohW5Z8agVuNJKaHFbpupsnEkZj/F1Fj/YAXY22RkYSdeaYTiJ
N6xIESW8BT1r08PuX90pT1KZ1SlxaCQc9dq/mUA58t0pC3jLPGnTLvdbnCaLAHE9
dbumeAU5TqH2V9I/ZhtfMGqbzyGVcg4xQLJoHW0jxApq5anhE4KDMhEN50q0Vbo2
NW/OewlNCoZtKlcZQ49t5UFNULiIyEdbkVVHxWGkbtFrdE4H7GyXkKE3iw/bZ+nB
EZE1jras28YVqzdf5Bn+TOnLo5sYG0SPXFksW3tb0XPuoJcB6CnR3/T5nZeSLp3J
XCm8djRBoyX0i371VmbEjpUVZMvQl47gyClRDsf4JG4zj7nj7wUcUdQ8TvbyZo0H
M2MEV6B9V7Y4gIp++stYrrTNOr1KKSDHe8+zQLNk+vjaMw5DcFOqKeRQ1UKOy1Ub
M6nqD8cuZfXMqIyWt//TA0t9HJ+9A+MvHbTTgEgh1oHr3JBw5snMy4eK3KVNHuIn
1hHGOnc5iWZyLFRzewB6gQ0if3F46xQr4L+d53/aMggapIEHFg6majO+p6VBjXs4
hhWd/VG2jT7YSCs0hyQQu8WJ78s6DZ8NYl7AbdbeNF/ALT61ky4jLBtq5Y5kDzNo
d3ZiuZtkVYQUbQ3A+IpD6bdVcIKPL/oIft9s2ynfoG7PfcnAoh2isjSgDLAKV8NK
EZ34RV6SrLzvmtevJSbaDCAeRtQ5wLszTGuSFPMAF5Rp0zoZ10vN2FalbLE2xgfp
EJglObYHo0hxVhBUk0UmXhvG80sbSUUkPlrAq1MC8wZehSXRcewmrfanJjxvM9IX
2Mv4UWw9ZJi9Ow0tBc2CueHAagEBXDSPP+rfQtjeausRdvIgk1cgZqFyugUvRN21
cpbqs3uTansLhKnpY1y6m9HO7qeDzLFxTKEDALAftUZzsfysYB9nxV1Yqvv4A1u+
appVyD8YyQUyoMTNepYY9HTh3t9pVripJiZpaYGetvaOVt1UL/CIp7NAxuSvql7o
++CGqromXHe4QtKFEMfHnq6j71YAuRvWV6Rxz2/yusu+q9rrAgetOFV1YMYbqu8m
mjvr7VYbhLrd6tYitnzX71ymCHt1+DyvIpIG0fE/YYRaDW1RFAnUlk1JhQxQNK6c
KHRaYs7w9Sd45LbQs2BbctlmK3kb3+9ZV4eDK3c/GWxZrDdIig8jJ0pj5K7rinf4
dee+zbaBfWQo3uMxssMh6lkRYDm4hlZn5x5rilof592RKh0UOptNVJQuHvWh1Gk7
hploeadPGQGH2GJJjDnGwikpMa1w0Ni7hQe82eu28YDI278Cu4aHmGNnoSKKc+i2
aFrJX3dmGlQo6ImfrlBQrAjg07+znIZJ2/yq4mrj5gCrpD5tiRiCmNeE3et/KD5y
fm39qX7QXCJec2ykh5+bDzT/PrlycjyAjk9QLQlNK+9iMuh1CiUerIX8Edq3vbPd
h8s89/F8hpe2rMHGeLdB6fL3onY4xwNNsSm8mSFUf62AzZXOslKt6YXpZQn9P7Yw
aAShDvpk3h3F6aDxNKImEMhine8JLPzwSre2Ih/viLUYMvqGC3Ow+FDR9O/CwxPj
r/p3cl9xyfenF/vCZLNYSvVBvV7TqhVJrYfaH+0IHh4V8jx58IznxCXFuWpk2v98
rErZJEUGhQm91NpdzyP38SztDmhDYW1Li/1dCGI8DI6CC2dwGY8eSIx9bKZb7MKI
PxDwJKrKul9aZM6r+6FEieD0WOSoe/La/6va7MbQfvQ4ujPnqipGzfB4JO3QWgaL
ZZkL0TmRb0v5XrJPMd+Yznn/7VnPCgCznmHTkzTD2c4Y48qeZhB/T3TCuyluDfe/
V/0RnVuk+R5nAoAxyj7FpWgE0iE04FfWpwk09esrD1rIhZzw4PSDn0jhNu4Do/Pj
3ARtf4cV0RrrHSuUMYJizGA6JZsiivkGNcWj2yccRodQjDa/v/b6TSVHllpwupa4
DGhID2u75tVBzPbUFslJkY52L2ZME0gnsEpjnl93nvnpw6xQ/hYC8IMBlfs29w9p
80/41ktoorvHH2J2vXuVlzp0ADahHNQ5rdYwEcyewfvvewceDyE5HzJlLehljUr6
miyTaaufvytZw8UWbXzwpbNMdz9HJoDTh0MD+uxBCRfO37yFM+TxfynfrhNC+ubD
+Qv1cvTVKstAc36e7opIxcKGuyysxN1gNyUWJhxd0ToLAt15jM8QJi+vkI5Hv7BR
UIRZj0qpcMpu1xYqQ1han4wb70QksAJNVJnMAwlu95m4p63M+GkV2V4DjrSEIiau
jetuyQEeojEiczaueXlcBLHCs7d+FnRAOenIcKzRyTH0qu/7RWYVdbN6Az6kAY4d
aqzrtdvl0vhJUBmo/5M61F4bAfPa6qtiA5NSkv/8C4PPUvtuhSPhlhFzFNYW4V2I
NsqdHUp07Vpw+YOAVCFO/p94VYOfKRqax+e/nHN+nNH+wFcI4PpET8E9Isdjt9DP
gKmLqeEBMrE1jkCooUek6KDLybqPFP5/bPz9OO9kx6yKhpFeqAnBlZVUxpEDNk5x
yiC6wEZejCYTy69WDD0hO0Yqdv/+LVsCXOXWh8ydx6Acb3RL0Sjsf7IOKCH06FPh
KJgmi5RFc2uiSI4X2Z59szhk6PZ4Aed7yBm3nghrS4/fhTovDilpFPKK/REQCpRZ
er5z/r3fKhaoFDwJwQQvu9jbrIi5yoFpxyW8AxND4To6uS+unI5UchzqNHIXqjKc
6+DpCzeGkfan85thAwI2vMwWEF7GqEZMJi40ByJl2DG13Wwl/DK8FpeqhKb7byZh
tDRMfXPYxPpx6PxcNYOuu9Hiw2/ow98kBrI5HRnoxrU2eWtWeMWrJlGps74rkpW5
6FPW/psqxPx+bAX1X0XqA8U1QUY4Vgr9+n4OJT37p+zldQ8nzNoQFznPqeNB1ngg
oa2JO2j+QtLBhTSGph4HjA40rE2N2lO25aj2vnVodGqM4kaKwetIio3xSde1JbgR
68TojLuu6qn4AAq9zkTe3PhyePdEXesfqK9Sbg5YcibHxqQNsO3DD2NWrKllMFDm
I44WynTquQxKtCPNFyBOprBwqzxyluZc6h5sIBfW3VCcfQfqoyFe19USXxMY99ZJ
L5+13brZqn5I+agLhhbyJ4HJ3eXuFDY37oiN/6smO/98Efb1SuBODCo+R47FnaMF
K4iwVj0ZorYl4YITZrk33RmK7QUzPM4aaUtonISVtlYa+FJTSiSB6OtJ6c50gQnz
cFxiAWfFi/jwEjgrwLrVR0AvqjEiXGi3bu+gnzH+kep9m1lThV1WGL4RCixuKJzh
pwXcMd1c9Hi0c3OyzC+QITp6twz42hbejA7saYH7I364BupoYyK5mySIIHwbdyMY
mV4qgiR403LR9MBZjlanev0OyQ1QqgPSoy4BpB8Lnpvas+Nbq4Gwe6l/i1RiJTA+
R4kpKPCkbUqaE3aamSZ1FBdjPch+w2Cm3Fwt+Y/j7hL31jJnEGtrD+5XvZ2lr7QV
wgGkCTBWgSynjvQSBGgajLCGvpwaobZxCR8JYLWKn+VINgH1D/xr+sSP8OBUOjGa
ha/52D8CrDO+hRnVp4SeYJTDZ7TtLSIkHeYtURySsW/pGjfV8w+6S1EOJISKhU86
Qy8Jx0nTylf8b4brY34N7A/4YmOg9WUqFxtGRUD/stB0aEWbRXzPrb787yG7kJNE
eqIOgcYaKzndtd5liP2LWol/aiUnKvUFZBuZ6/0Yvj5IBGiCDltsihVW0aD9mXWP
aexGPVPcMH+Bb5OkG4kOixtV976ghX6fo0KVNt+Qd41LBFHh0wbhtczN0loYuZOH
X1dnueCpdMroZdBRWZT5hLvYFBAHCOqiF3LbdNJew3qxUpi4XdtQmmTGSG7CHi9y
kN66gyey2gFtsWNj4oS03yi7voybvXaYPhVZMlK0WCQl5b4cUEzniVna/OI8T1Mp
FhEAEFUaeicXgcsc5QpZqqqNrT236JHEz5i7QFWJDo/hNaVt8waScvoui2JsC6Z6
8AMSypPgAC8Cble85f4eX9qQGDLsGS7ZkvJFMNgDGQNv8YbRzWxD56TlBLHB+sLs
pNJjK3ZqXiiEFu3p/xiEmfPT8huXjmcnKnwcCief7XaLFalLWjLwKpw5EPNH6Fae
h6V2jAp6m7o44u7wPMh4CKoSQVfZ3Dd1OUf3yF8rxwldwvluzndSrwaymnTeTzv9
fadmx0B/P9S+6hnCFuAkfHZpgBlbXc1UGdwzNqC1uMsog7tWNRRxqK/85cR8wXy7
NIHW501uRVqnnJIUmfKPaBsZL5GfEaYWBSHc7d88RE3vHessoBjR2ZlLHRhzlICi
vh6kMQTUrU5l3ImaUPMRZU7LwNN/a8+PosizBrdlwcSo8OIqb9Rqk6WpmmHvsXB1
kxk6zAd8EtgdRBe7Fo5mvAPyXa7cD5DT18uZJ2cz2e7GIOJTl+f9nSH9Elx7Lepn
3COuG3wIItAy7PQ58/6ai0qyGubGR0r4zdqNUA8oi2KoYBMH7lB35V95IvEbEBF0
03Tov7Pa0EmVvYfw6DQMau3/zScJQnQgFQn3G0basRDgm6L4riiYII0qThPQbXB+
EcE87hz8P77U+GTEJLtyb42qvm68EWi37uRcDQPcCTR8+QBFHdMZ0gBNgWWhl/NW
ujdL9OoRw/c7IoeJgF2TIKBfcPWiCYuV7Y3BtICCk7XebVFNT0CG+vbT9R0sI4EN
sLHPm3X6hMhPNnzHLox9mgyOYSRz69hVkD1me4NXBtZvDJhIy0ufNWfdQ5oDMthR
KOnHV4TA6fnajliN9R3i5TaJf3roG7dIshhwz0BWwC/RmV8difrNz7JbNwdn0tNy
zSHkXTy9xn5nfB3NPGYWz4a07oUIvpMMpqkuAplQzqVKFfMhX+zBOJIyOalU4cTq
KvLnVW7PR9+mt+DAZrzCmdxI6lPqP5DJ8MsnTS3LkoZ5Tdxkl0nrCd1e05a9ke3H
76Xz+Y5rAVdodox8R/HIoOIoxLWH1sbDacx1rPMeUV8ml0UUSe5nUKnH6EFkvSSM
wAfeEZp1k2Vj8DzN11ErRMuCZirXV6134F61y0nrqo4U8ZUh6nr2EzNW8NVx/yFa
bF0oAJYij8m9R+5UyKsUGAYZktnji84spV6Svxk89aRnw6xXyN0kgs2NYKGw0TSB
/dkOvEtzSU27DyO4ra6CsnYNE4kVlIglnoCoU/ZKoh/TsV5bcJTPcqqpXPnpOHgr
b3jP+S+tt6bWN5yELAGCfHd2CQAMGvixZJPLxxPrv8SFrMjX4AfHry4qWLSehvzB
PWtMsSJiMgNNndoikEfF7pv7UO3z74sixpKn5AV7N1WGBwPRRzhv3H0rW9mx5SVi
XefO1jZQJyDTBNsYnY+6Ujc29iapOiFwC3DhImdpBAqxMxuazjiF4lGFCjt+vNVD
teX6juClQs7RrHetSsjpXCNsY11BSU59j4pGTbEhWanEdhWMbwXIRB1Lpw4coyS4
+A8KeirUqwgbmv4ZY4ZX05At3ILJ3yiwgfgcpZcaD647aq+C2o0f0SPEfyvciGVn
dkw3FXqPh98dGGkcIyHY2FIb+y367iZL+uTvOJFHOYwDqIH7FjQWL8GQdm4DNatP
zTFAzv2RPc9D6fiEjDclNyjnhhjP2O+actHpL1b5NHU7qh0/oaWdDOm8hIUrmJK8
R594I9GGa3tocxqZDzMcJ6c8yPHwGSXXh7gGyqFCcIyPcG67ososXsw2I3xhf5++
2BG9sQl8In0rkzJ7SgAR5OMpagG013Ng8lmaQGaDXvkKv+xih/pk/JUbEP5CqQ+V
9JFEUvUEVn5GGAh5sVvBnN1ISHb68Uz0caZS+qtMRZF9ztAbcHrWTkOKRgx+ABVU
r1/PLBiIjGL68WMqA3uuU9JJPNsIYguYIfJSXtYNBEmbgpaFQdau52JTvG4T7JDn
e2IywXfzRsHzTGTo1hlR80HimLndvEc3GK0GaC356jR+Y0yO53qEE/7hChVMhhZA
dbzGnChBEc7HdFVXlMeK49Y8BYeqTbYb1vQ47D0gigiO691G+2MKqR2oGN7egaYo
9TwFqW+aDewcYGhftMgspMBhQyyr1MxDI7yq2C+HfPl3lbJRgSAuOBqAnVWrmG59
hIYdWG6nE0/rXMutdh13TEEIElvkKc2s2cdxyo0rb0CPCfOqy74SLxjetRLYy+h2
Qu4wbh91uHsk0jvILvrw6XXB4wNy7TOJSHqID36GAO5Ymk0OEhXVFuM1mcHRuvQQ
3jerS7rSTe/mmL+glyDAIgThBOD7uyRGXvNLbQRva+wtu8apgE2P9W1R1ezvqiRU
0M9GBuKCzRftXVrZcRXXIXlVMKT7MKAS9qFwCjADfZyFRuWHI4gXpfJ7pTVA3S7G
+z/Wg7RyoYGySNMlDr9Zbq0V7q9tpfTVRB0JW4exHhFn16j/Z2eEfj2mB/VOmBv+
JIG0NSSdeGZdyEG3KaVOphXl6qk9FcOnp8r+vmpbZFy4MD7XP+6XKgpqflY5CtWJ
EklsBFuaDxlgibc0PiseFQQgDqFOE3BC4neuelxCNuTjCyldcylrmuwECGUQ673A
wz2v5MQLMTq8Zmb7p9TLplTpm8oaatvzEJ+G64Spy138jpRuU9bwOCGHhgEhkX5F
Qwj3x175KYhF0QxnUsRj/EsZgW4O3wfTBU8JGR/P6UUD+n/kCO1MpCuUdA51CKgq
7mfLKggAZiqNRMUD8NF+kg2IQdg8KVqq8uLsaZW3RxP5OZYKw5lw7pPfHP2Lqk/2
AVC+5nKDKs1Cf0BRKXkbABxCLzgH/rzCBPyusaF+s3gI7aJIcbg6f11sCcQhogwf
G3eTNOrGXHzVTy295FNrTFb/J6MAagGZZNKd/5hBVrWUgfa76uMmhj4jQRg0HdIk
5xJr4PN5qxQo/8FhVgM1F1oa9NNWQlWt9vz1OcEXpw4lMNU3jYlC4l2Yaw2gmGcX
NtJrHW9nP1Q44U9DYOMlRG910XfNFKzVs45N+lc+9YWRD0Tzq35g1Kj9l/Ki/zvV
EHvA3TRfjHCZ8aoL+MJcEldwLn9Xx7Cte0+i4mXmU6hKOgQaHSvyB0wAxjXh9p/3
ixv6jTy8c0xSLspDAJsgw5jn54gB9dWglDc+zjRlUtikmQyLKFCKNQa5YDM8AvAF
21fdPtr68WQETl9zxRMyjAAKZVZBeCMeGVvHicSyc0c6l28puT9iwxno1+Wqf3AO
yb44DFMCfd7Rz1hp9fjVUdvNRUhnR9eHKlf9vOxh5F5lsq4MfkS3yQB39UnQxACL
V3haRq3Bg9FfunErpz8KKYPUeiFDa5H1GosCG42AeMKOX0kvTUPexFYFuY2uoEwK
NMrzuZU4vI2ROFuZjdmL5qxqTU38eYtGjAde5sLEDREKhf6ve+aOt9GpgvptHTXA
li406IkVwY+cSgW8ocKfOPLnlBKsDZ40IsjypWoe5AUhDwWU3pVqBIQwt0dcMFib
0zZsUavxxXkYkTMrdPqjAxJ7AuEM/VUW819W83gC9dZRAEG54LkFci6bmimsp903
tKKyj6qmYbNyeczlqgwtmdrVX74y8Bwz6CQrvg3zlBoV9gtpAQzavo8YY18AuxP5
8EyZnZYhpepOcPVjeurJV5GVu9gjQgDo/3+WVT9rrhWUeFSWkMuZcE2gAq3jdafD
j4VD3S/OX/Gdpk9CLKUXR146cfMCxR1XOsZkQxR0PoJqmorPFAJYHElJvfZ7UQFp
XsX11hwziizZngcE82Wdh0gAGYAtaZxxJgdcMz8WbJOp/vV94SYyH8vlv653/rdm
e6aQN7shr0mNpYK8UcW97mTMaBWSfZ+DI/h1GTUj6p83w6MF4yjtYtDL34BD2tWO
Qus77CIfHKN4Z4kS+4qhJisijxsJLEzlztGrR7gcruEfm/lun1d8A2wjBDTJ8f7/
cvO0w/CpGwbncFhJsqc7F/dq36ey/r/+lm724oGC4cNavgUBBwIGQ7gMXheeJ1wn
8RSnVzpNevZvYEIyxCdKzrJhaaU2U6SZGTgaoonjL0nHD1Y2NIdPmGHcB5ynKmB4
z1DKOjeo/dRsflAPjfF9UZKjBJOfpX2XUt6MaTjpVM30wBXXslT72iK3FkLfGzSQ
ZtFr7wseny+XerPiw07SZzJA1KolnBA8O9CJGj+A834pKqsneiXg2BGM7nVCrlBz
vi6XkbJjyHrlFlh5ZNalv2soLbuBw91W5KLyQjhWcHo82trKGxcc1jxq3CgcvWZj
G4rKm4GuRxfDJfO8atSqeMDqroDvnuwwJiUu9dV8cZbaS0NWKnQqPnr+xk9HJIAb
3fiCKS3VAzoAxYjYYYzosr0eIjl4WeWR5QTvWrlxzFJjYRSuzxA5zjIY3rhhcGf/
ZWkEisKiypz5EgOB40XDJPaTORq9LlefhbW5V7Qg90qyljlhKn3i0i+mk0R3K6ZC
C49UHMvKZkMLRDjRvXaXYxFof37PNyAmY8l9ojWCoP1+E6QBZDLatQRb/PsLGO/W
KXLfDb9S1MJahupcUsgBsGKZ5p0p7bcSrMFQmc/lE39Q9O5TcYVTV1nx7lui+gY9
AAxI6FHFruJi/8bM3+FhcJvM6GLZWgrn4lok6mvgUfF7wDBm9rM2YDmjUSiMEwDF
mFICPVwwLNROfJMa0lvfUehUC5GYsRvuf8E5AGNrLg6ft1HlwPuw3x5U7uV6cTEm
NJWxXD8CG/7d06tDJwxdZa5KEJbl0exfOOMGJxD+5xUYKHnSP1buL4/++XupGXT4
qnJLQW3MgpTyJ27r0hP6RCsBjl38vcGstGpreoIXlnZLXz9bflrmdLa0xrDlGKkn
JAHcuVDKQbcg/8DfEyQvwNaStI87oLD8Bx+X9t7rxseQ8DSPKn+Oze7Tz6D/D1PS
9BQ0l1G6/ErHmnjElfYFCWM4hNIBu1wyY9rjNhhJ2LmytqjZEQ5lKmks+mi8mGs2
aIQe+Yg2DK8B2IEPnX2pOaAfVrA/y4R8F9TnmqYE0z0tCslXQ//SgCykqBjr+8YQ
km0NteLMOmZQxKyb9HAMF/phmxrbWAftOmNYYcY5Z4AWFgEXWvY+qYRZi7B/2263
7j0PRIs86jGhe6x+LpPfC0bHKfBbA4CgooKjHFSqh0nMgl/OPazrqC/S1pUl0gfF
WkLrh/M3UeS43I49Qi5bTvUwhcg1vmIYeU4hN8W9V7QUowJL856p4l1hzilveW6C
4wAhnfheK/TJUVPg1HD7qafY3FYan29gJAVpKugS7dgHrjLjJ0NxCfRR0MP77NER
QOUSp6rorIxfoad9ruEx1h3a4u3nOL+orwTZ7PReCKm09XKIMMBWWsResTIEPXn/
VjqZLe456I6McSn3BAnm1jgfpvzuyfcZQi5WaGzu0kNzQLzpxUu6/H3kR647xvit
6EElzlfzFDQoRe8AB2NuO6M51A751+KGPaUfbDfJzNNUpW8Dem8lw31qHRbiIwq0
UFFNG9DgM8x34mi4UExmXjdL+A7hEa2YqhpiV6pevgfT6IyHsGOGfw6+88KHlM/E
K10FETz0NKyvZwDz7sOjTQdxAzyfI2KAZ8aGWCiRka9SzoFEvqB4BAn6qBJphRty
0T0tpe21rHlt4R8UpaV0tOcbczXULa3IoznqZSh0YCQVZMCAUGHiM+IZFsLENsr1
sfSFFblEPNVg6YK1qNpOVon/1F0+fBWPzUy5xleOiJ/f2YjPG4mKxb7641Et1yID
GrAMR5/ZR6ageqJ/Y1uy//st7o0CxlwNt8GT0SYZic52vNpD5uFjSOq3vwXcTEUL
UdY8zDtvCodC0mawp2DsteQs6oo1M1LgZxSanssKlNloaersVe7PP5Ks9mYQVZCn
7HBg8Ama9QJx3iXAA+uFVbOiskJYdYPUxvTq4OAHBYvPqu5TLS726Ztc7DJ9YwCy
sB7OLCVoiEU7tQZLqYQH9SQL+7b6SMnj47CaRgjJlVWfLiNU2mPpdwKyreDgx0Ot
83WpaE1rp26W7tOUe4NRUHwH1Ao1bS3XmP6rJumlEF0hCd61od6qNAoOQOX8Tu6m
CwLZPfzljTSSlFUaiKj2kGEkub/5kM68r+VsH2g3YYp2DFsvZbIMjqaV/6Crm2Xi
oqX0T/38puTNh1gCCR0DyCUFNYp+El4xKBEOaxEktCbnh64exC0XgS3tleKInNOq
5X+SCS+9G3+n5BSqDUJYg4gm5ybArSIGJb4PLgLgwKU/y1yJhImsIta53zODZXDu
xQvAo19pGt9VsnhYgO/AmVU9MLntRvbvCBLmGoGoFZ3xzK4EeANbPJf03sbY9C49
mZOVvl0ImEOph/XVEVOCiMbSE1i394iykWOrH3PvvOJZYfnaVKtp0UuTmtg29b4f
f8v+RlBK7igfoPoaGnCJDGwWZdyLEcFX5wpuYdCaKM30upcmWkmkR9sw/0bkrOvx
o5vm3Z7w7sqjz657OhxoSqeqxlNctlR9+kRMX6vhPODx7/t4yWdm+fdrEiuMfYNO
G6W8AgA7sAHbARfRItcxJQSpV0RASv12XmrfkG7JxM05OsZcRGfV9zWzyZGslNVX
6jVGNAWeC9aXsEtuVkkd9myaZyLHl5RN3jlcNnkhxkcfpnjspkvTm/cP+9q0CpPz
ZP1PPs2oqK5tdqoTzN5aApoVzLClSanS+v0zCadwBoleOOz7s5GvLgCBqvSC8CGh
6rMtwPHiuUmLrZa93FVMUxnp1Vza3wUiAxijGYy8Rfz1ogdRq2lV3as4zM2hOeTf
4C/6OGalusyA21O2Cqh0+Fq83rSqTNk1OPj/c/QCHRck+V5ivx/NrCoNkyctG7jR
I41g2xejbqmswc/C5vtBEFDxcBtCuj1f2m6GgQp4B89OUCmK2O1CrmMmyXGd1+ey
Nu8G4n8e3oaKrphhkPmp++tE3xbDyu3bK4cp1JhgUNHpN690BDVboF/1y6Ye7LnO
EQJqgbkT9gVENN7CEzYnlVQnKeDrIJGnev3VLHUs0ifqc3eT1lIuuLRGzZhNnNG/
+oZjuDBpDwlla12MqyM47aNEFjC0TmrWsAO0P5fAZHDef0/MPSMYOmBi2tUo+E8M
zXbG1Z/rxRLCxAo60XvwOhnAGEMq8nw8iyDq3zGBg4TdWt5aDXzFTwEx2QyEeOIS
DUTOMYxwYTFOzughRbMN9uhVh3cK08w7ufVVRbv9zJ6AuBb1TvwUyttDI2dK+G6g
oaLlyrJqgHQlfx6S9xpOI4MK5MxrBnWq5tu9CgGuDDteCbX8dqt1EIJWy+9qcyFZ
p7V7h+hzKZr0j9JDFIyMVJBMWPz3Zfqkfv9o/MWS4+T7dEJjcDjfb+9yvx1O5+kL
ocqmQOsEYs7Krq1EhvxAIw87N8a+2sM3Zh1vmdjqTDw8MQkoCjpG7ltrgPdvUHPb
GH4dXC+h0AwPJpt2pP8RUFwcOKt8IIeGr+zCmEJPTi/Fw/9BuxAyM4EgCKXoq97f
egRHaDZuyK5nXlH49Udx922ZOhL6q7GIiCmAPB1Y6HoT+5epoWH40AlAsy6VVDTa
fzsKxJOmH3yAL53oVMxsNTiQKV5pltbezW8LCuEt/pnc56XDe9SDAxwRNJNiG3xS
AcOp4K8yaE8aUm4HsCyDkbMoTWu5O1Lra+ePsz9AiLQZ5t+izT3ws/wc5KExdoO2
7gyRLBXRdSvdRZwR+Njm9093c978LnfDUTn6j6+TlUZfizASLkfiGoYDtVoUbm7Q
EXeCydHBKFuCELUC6BH9w4EVPNmwfyORl94bIYsUBB0+2NtZM7FhrV3osVn7L2Gx
n48qjZ1ya9ZW/uhizCfsPmZYbRD6sMVkTuwOc/UtH5L3ickexDxwLkmeoi8yNe8I
e+pUwmBgMkbfqUd7buuHg0ZB0NhD3CObklkg89OMsa8QmmO0IpPysOwTfyw7OMuU
zdHubV9B0aEvtx1LoVqNUd2LRpABYawU13eRRW0OqvmnhYkunwpmRbQj/t3urAOv
VcBPDbiYfIXfYGYxuqIxa7LpUQhjT2kOjB/06Y7m2FgtV7KPjLJ559AkhkCF4zbQ
vH4Mgo2gqBKpdpr5dewEzqlxBveF4Mm1eb31MGj9O/E+Nnekhx8ICXiZKekFZKL0
sgqJ+wqUej25sy5LsVJ1OCsUBDZxI9TgtmhWlzu2+HRIVC97FsIJBsyZd3GpZMsQ
5ec1ob6zoaOn1oKXVnIq/dvhXCSjx4V2SSWfLVvpDYhAIX6MjQBluwWYD9U6ZnMy
i+2t86iOKxZ3xOtGAnuxMViP5KuKS47k/PWAmR+f3bRN/gz6CGofHxCtTxykMASG
+nNyAIRnWJ648/ZxusRhX5Zw3oARODvxzdEpvwkE3HWoycwWxBgR9ljgK35elBdS
lH8HMrbOfR1rU6Dve1eE47uYZKXs4RQLPHq6t6xRjQGA1NVFFcwQc52L0XMmJSyz
HLRX2HGNoHlt1XTldNIcUgIw3/1sEFDgJo5ubmk7G6J1ENTOq76nblIq6HA5Wcqe
sy6gnOGkGQKGipBP3E1JCKuu4pQkKUbzRtbtOMYvdZhERPTtHY86/7rM5/lQ6nCk
dVwz2N58gxJN/FfKVT+BuP+l2J5kRgUuZfU8Ra/x+b06R/sNTBiR3BpRf/JWiXul
fdS9/TTqKUyOSRnvWmX1mwI6YquPID9L6OJMG9HqAOZcRTUD498HrNLkpcjNQ4jy
W316e7Z2xgVIOHNc3FpC+b6+4OeL4CX1TphMDv8od7so3147tRdQc3giVmwGTVPm
kX6ZYRzARMvwZemPZotU3ecX+zqUD+BWosHFvAK+s4hy7qUliSB38iN3N4EDxpnI
7GW5MNdhOLOtVbkDXjNiohbuEzDx8dzTep+lcEZU42BsKalXL0Oje7SwTbXpV0jc
pnwXMPaFC1TUozs61uuBZlAzjtIA47+83HH9dCmbl8fVns1JpNkBWDs45L5N0LJ9
BnLd4K08ElZRiV4Ds8KRVrwhBaXOZfupy6cxeN1VDD1/5B9QCGrrmkByxJn+wuST
Ap+/7LgW10FlDOu2AnBKRkCmAYzv0dWlXOPGo+fDUfpkDLua1IdC2nCzzb4aH2DF
Ggm5huv9usjBDcCF+aG6t+kEVC5Xn4ocf1ZGsqM1BoYapPsNcm4wVMHbsQa9KBLi
l3x5ja16Qn4tYkEk7lsrig7ajL5savtu7jsvEm52uOfWqHQ6YFdM7ezigUaNNG6U
VJrrqoJbVFVaEwbt6a7MD/D6BX75Pv6XrJSvaRMKrKdVrnba7OnKaDDeDODdRQIe
PaQIFr+0VKqGkhtqdVpc825eGZ8GdxRv4hsOAulYpCjYtVwtJhNaKNX+ZQSZPBFe
5awbqulu0d6Ite1vBo+wwMVIRnp5tdAbwXl8JJ8ZAfrne75lbq8QcaiBuK0LuynC
ChyJ4x0MHOi8OrnBVLA9u33Dbe5DgkTuHBDk5jHvneR+6gDV+L7Ee3VbpIXpwi6A
VznDXbOJzl+Z4vHPW3uxZnX0WrViatoVoQz1GZ4uSbsETbI4AB8exzFhzJqr4m/q
DXmpYsPfGfg6DT51I5uFIBI3A8phF61H9gRw9jc0Lvd5QO9cvgsTRlw72esoJO1j
W9G55Tx8rudmaLops6mBBWtXF1HwlkQ+xsZV+6UVt7AME9FQ9Qn+e9lkGReBnXhf
TdK0M9gBVovLxZr2bEcHLaheazndJtCXf7i+yIG4b9DEjBkuDmkf+vialK86ixvZ
tqww8AQAbieydz44pkiD4XyfB0vjbGXefbU6/CxlaUDQf7p+qAXwmUXkhI8V/34d
zb0rEHAxwhvf9yXcb6Ylhd/t4m7pkyFd2q2JnPJ5psqac/J+IVzrHgkwAejNwEqe
esFPc6Q4UjkHmqPyEkYsSFfcccHsmG99jBNk1SP/7/bLuIl4UmoIpFH8lbRioRV+
NLd6EuHlojYp8Bds7VKqz1HfAHC0xaWxkTl2U/MOKIhiEiKFd8bGd8O8ykKLFIVO
+Zov2N4lvx4YhqaWO1ONjvV9gCYRU9dwC7K09Bn6PsVMVRJQV/Qy4I9HdJxzPuV2
HHv26FmOW5bkjJLo/cBq9a0Vcj8DS7mrbblVItW19XxJumFl+uQ83b0zIiXSpsrX
k2Yodg2GcvSm/lQsKqrJubyxCQUs16h0lRs8r0DObLL00tVgzdCFEXlqSMvSZcun
KK6CTPbdMB1DbjoZ7PkfvHfFq9Peyx3yNHjHMPX+Usc4v2pwkLF71RI2de1Ifnjh
HqHQvaVXXOYAHlYCENs48ZkHm7bENQCQ93ALli+1Ko6bD444ZTMVkmo1ng9ZJPc3
IZqqb1cr4Uf658l66pDQkOa5RyG6Gl5MHG7naCG7GuNIfoToeiCSC5J5g8eAhdRD
ib9Fz2JmTI/vO5QvRKFdwSd1uXqtmaFfhLcNLVjPJahFfkzUVLS5T7hU+SHKArNF
/6vw00fyu1KfhZzvnG8PzoN9mlrMEIiAiDpDg2Deo+gGLuqXDFTfimOJYlgpuXPf
fzifWpyOL/t2hLoJC+I+ODYMqZeanOu/PjA5gtyLgouuK8iaM4HzvNTtsoCK6Y8K
A348M1mKLiin0hKZE6nV0aO055IZwSz2F0y+4cZQh3VVf0Ki08i4kK7ZNC5wSjIC
9qQcpvNLjKWFf5wYvA8sr/7BjFshvh8u7LwFdEGT9ndnXt7DdTFX+X/E8VE2Q7rN
WEsGwA6b4UUYW6VhLpRJ5XWb7VPggN9x5kepOpmTMM0P7swStzIxWAVtGiIjoib8
hwt6Cb09zy670xkxPEHwGxjEtSjO2wRGrhlgV1a3wXKRajKCSSLNuXVXQC3YMgMO
mUwJjmRJoVyAx3mmMTBBIP8tPtBVxAc/M59ehGCxU3XOBJwHkW3n4vfXKMA9lJOt
Y0WIqvVdqR76IcIpmrYU/KiHNDVU99QJQfwGX7UiZ84TM08xZz2NOrAdf/G33hIY
jXJXlWBnB0JQZLNlObj7d8617+HoL7/Yoh3XtuAZ9lMqSuvZ6BSw3v6FcUwVZjGf
wmXgSGvuvSsIctnlEDU241DByOa9Ef2vYZhDJQ1ZgtTq0XOO0GErPOE7SgdRRoj/
AHqT5B8Wvcx53rlzn6Az2wFJkg2WVlEOJV3PDOw3Jtgo+l1pLcK7PYzcU2ujr/pX
JrNAojRlqMw2qIe2HSYi6kKFLNwvVK/n/O3HDZ7jXVO04TenwmaM8FCFaktkkTtp
pmgr6zM+2nAqbFAXNPHf8COZ+addFmjC4tXCZxIDtV/fc9tMxG6MX1JTwMwaW8VS
nxRpjwFhfgLwAdRx6mOYhAN98JWzuHlYWVBqsolFFRy6X/HoBDM0PD8bxHe3ik/N
4jGz6ig3DZ6l8nC5fF5x5ZvV9todbzcdDo71AHdCNDVSd9RWPinFUiu1wO/M2joK
gmrh95LseleF0g22l4gjWI0irazOh/NUEzeiVD0h7WYGdx7Xpa9r7ZR09hAnRQju
2flK6pl9aLWv4J7q7YRK3/wGmyktXphnYDjYQbrZduSi+zDEygc3PhJ1631BzaO9
IqDHfGF/+N4DRxA6/PRTjQGeiHp7Z0n53xHmxeqfPbBQkReD+xWGL1+mcto7lauN
lsJVaWfYBCxI4xUzwV7hq4SRCxxJD8/z22ZTbdmvcJlWyhCDJB4trvS1zQmBthVj
cYrv1ZiYT1q63i8oE3SUrwHkPzy+Wg0Qj7Ka1BmopUhxziSbRHaTPoDJL/A/w0eQ
s/N1S13ErxMzjdMyFVjBmqpUs3+keoxziwt+SWea5lcacQrWX7UpTEEA3wi5fUFx
Sfa1j0Qn1NeTI+JFYH31QHd/cTrQpwnIn9uIf2nOpmuIGSejO+9g7Yc9YY0S/6oP
kdRxJjVEISSrzHnGe4j1xeKDK9W+gq4On4innhlutJBjt4M4rOdTCxRIMpNPcNYP
3tnQ+OirYpzLbmFZX117+FqlBGOScuZWd+jbvz+qYOSqf4+dI2mdrUi7pnNZPjwH
1u1Xo07QQx+AtF4sDjm1F6qEJbUFFdomOp7FnqPgBnnTI6sDRmkaaoyiF6rrayG6
2aRfLaL9AJjrPsSbxAY/ShV7FyEB3x8aaUUmceBtAKNV7dJXqEF5ZK6sdQ4qBGXv
rQx3GVy0bm26N2gGJoMwypqzDku6I3SRmT52HX2OJIjmdqdJoBfSe2oXFa2Dh+mR
XIpHdXDlUMq3Ql2EcDBUqP0kt48tM41fjC9mvibMQeqxJRd/Shk29gs49He4MFjn
fGmXp4yf3HqsoD3gQVROZvrHmniRJcwdhwTCzujCsag9QvZo1UkqNfZju4Z9jQJb
EFFKRjZEJew2kOs1gA67mFZehB5hFEM4sFflIdjHRZascr/vjhExTiU1sNze8Nfm
1eTSV3M2uPvAI4Tc1tzaKl1vdEiY6aWBvFCoolTJPETydzVPgKAqRk8v73xm6GTd
/kCSkJ4GX/r5LS7A/l904iYzFhkgg2u3Ntwhbei9x540KuavV10wnjMmR63zxlOd
WfOjIFjGTYPn+tH64WBzdc9+owQsaqnuYfcgDxhpx4Z4HagBMrhkTe0I82b2fdbs
CYJY/D+21z+JkYgXM3KTiqSNLnUxyUR7SPNOyN5Kv1b0FBBqWloNlbVDeEHDUjyv
S4I6SRdsN+PNpaFdviRwA3hCw1iu/p3w927LyKfUN219+TvKUj9TG0ggWjGd6iSu
mHaODuVFlSvRW8uWtXAD+szd7W2bmiylAP5vHrjlBv/IC5Ftg0UEkovaZwhS0DUx
C+VnimuroYzBloN1xF0VR5c/+8iSxMEtLZs/1GcypsCagLrRFGTRaJTStu5X0fVc
zTWmPZVnsouBxcGm9o1i5VHxhiHLM/g4HscSfHcsgHGvasIHRjNjPxt2lav0K/OT
yBgC+QyYqt7NoTXs5HdBMM0eK+bLOSQhERTG0CJd78KEPpbimlewblRCjO9smGyn
7XLZ45wX8PpjzQJex60CT/3HM4K2+8xAI/h7nMhJePXlfjIc0b6vcMwHf1bG9FD+
U5hAYh4M1i9CPYIaRPaQKf4Z9yTcoi0++q9zQaiIStkNaWyHjku3Fu6FXP5Rc84Y
c94qF6eERgz4kFeP4oVaZDXcDAMEIrofPBaRo8Qe/fJgRv7emJUX4P4lEuq37p19
ZKg8fgZ1I53sQny1cREZPg1DlyGHaguJySEJ3t8DfEXGmA0ztpKT+WI6kYSp0YtA
FhpsxOfdeGm18CNEPMa9XkJCPYQq8EwPJh+YUzXPxKfwFSs8PN6s92BTgQaPj7VV
J+soG5I+v+j6lk4UMX0WZ0ZGqc9hi6EbfOv53tbVAr8B/JM/CdbHoGdsOGisk+CK
tL+lt9YtrwMmR9IOw77eLeaXdt4YeJGZvYGM5zzOhBDlAcEB4e0WRssMJ6FJbp5R
z81RuizbcL2pAnbm9v8rOD5BE9+UOYVgFb08g7+OaHO5xjOYLEv51j1VW2IDQNqE
U2kceSJgVQlcjXk/cab3qX07S8aoVxjr5q9WIi4KRVVvBQa1Ecd8f1zHl5ZG+HI5
WNAacpHZjlMnjG+ERhOAwq2pobgOYo2lTbnmeuHT7CdS4DHea9dI6gtgR8cE5spK
36IVeKWrQSeGmVHv7LMOb5k9z1FofmRD/sK1Z4ZA3HtX9kqUdNw82RwU5Ayz7I0d
QMpIdyHtXApL8fI4kAkDDEU1g1la4wLygrupGHKLLjvJSzHN/ci0+PWPVjTwYg63
LjFPAd8hhkH6XvE4adfF41MrC/foFrhdpibFPGBBYgwg6dq/tYH07fUErtAe9TW1
2mY6WHxvjr+1gnxJBp4xQ2Iyf/cGts51oShd8Ze5XxppAIpKrqckbJ9ZeoRo6Y7D
L8MWLl4vEWweMPT47zGu6+arWTO36Dr5SC/hWi3A/HsDwSBu8ezv8MD8C03R+ml4
Ew3CWHUDgvaZJHrRFuLGknFPB+7XH/4Hsk09FSjirxfBAs5uEu0WSFs4wI8qdhPq
PybJgSjh/w9fL6jQtPASnPGwhIMkol8lutUduZqvO9JMI7Xuapos0wt4WZC8w/DF
pzQOF/7M9uAECLkbkv7XmTIwMFH6tdScNIxbuDLan0T6IG7QKczjH5g2TAL2xyt+
1WyEj/QsqG2dn6jNrxyscziZ5pDvpJQsTV0LWDbOA4aJ3HwjSM85GyMEtAVh+Y2M
DiH6LoQcVy+eFcokv5EMz8vWuoVP7gf353//yXTyswfx0tAWZegNYo2lZKxL7V9T
qxXy1J9GVvZbxQFuI8aAPCbTWeP9y0pkVkv+HdNuFAnQoJrazhVdAmnrcNHRTrAW
qnajiy5/FaznHrmSfxw2A3qxbmUUEBAPKGfrw67vCY0SD778Nvyt0Zj/lciapYqI
nO8QcCb4KdWCIoNX9Jr9Ppq1lCBrTJ7Iynjg2+Kf07Yb0eRcplpP33Mgc3Aga7ei
txXcEUK2saTKCqKkT/gvibHYcR8eKRwgzvDYwHGvc8lKA0Gv/Sx0DZ21LERVaLIl
0woPA2M/G37eT6nen6QgpGJZsnFngGM18FB1+n3ZPecTyP/stK3kR6KQ+lpdkTbC
nweTxgxWxKvzbobmTX2c7NKP0QIIoPR41FrDcW6UUMoGnPLJV91HzUSM3g4AM9sx
/yOE7Sci6XKPDyX5sjGkiznFRbvsDsbVFKLrcz6IqxMeKAPVC8Cd9oBzn+bv7cGU
DmdHYmjrECoJtf1DIiTR2VQdTurjDuEjSPFVX2pdRiYAXZW9ULbiL3/NPBwO1Epj
VNBUOxSt3x/1Gf6ZpPw5/+k1YfoSUNLn007rb0efFtEKiJmHRk5oCfZEVZVfI2l0
1a69yTz09DAr54j0vBWZ3VUuiudHsZQnIcQjd0OqvgvkBrB1bEY84yyO7jIIIJ4U
zipjlvZRC3tKiZo8Q8/nNuiretn+J6qs956QFiG1Ifg5EDVVVjsc7B32hYJxyFbB
E3J/qqDmNbiUFDT7sVOQ+icv73kZ0R92gvI75wtbvUqu/dNisc8p1qx+KQGiv5bs
UeU2qWAnpncDAC4R8JrS+m6LPxTS/u2xgGDzcFrMEuZG62KfEYWQRCjstPNFVpvU
oD+JKICa7Wx8IOCrzFW+KQVw6jxOLiNrd06vWj2Y9CnudL1b9hxUu+hnManga/SY
BfK1XDJIz1PzpUfDtXIj+hW9LxOp74NaWQQnsqdH7lzSCxnAXEFx6BbQBUZiMUjp
l9ZT56wtY0chcgmDJhvqgy+vlVLyveJw/K2HtiadVZ2wKFUs6nuYz8NMKvt5+mOa
1swvd3E1Kfe3Gq9ER+kpS8B195tTWsyCDyql8LjQU6IsgQcgHkTFiaUFB0/MV/J6
Y9OxLcXcZpUz3jkBc49N6ZGofZy1huG6SWrBvQ/dp+c3E3FKBMs+goDIUolsWtvA
aycMbwhrYJwmTTnZLIaNAGUSCNmaEKD2hxXWVwDONdZt05172R2CEKUno0UpdSrr
hsJj3vpk+P7D0zYiFQGldD7Sss0GS3vYcMtMvYod3zX5oCqynYxAKDFpOasHPtnV
FPbWWcgwMbXMuQhryeyikIYBuzrD6KrL1wJduf+MWgTxUfp3XRSibHW+VzJJ7RmB
WuiYhDTcyQagikdjB1BISXmi5FnNJHTQc9BHkbhjCSgrYCeo1ZSkuQurzkj8uc4b
wXjPu48gyEN3ov2ezHIZJE14VnAEIOpqFX5ncy9VYFJGhJJ69CJFD4mT6goxw/S0
mWdKFD719MTFI8w3Mivrg0n+jgiMY7WA91f9g7GrRypOaJbBo11JsdbEhIAcZDBR
vfWSBBMxPtFSyMyExqrV/QpJ5g1Hss2Kov+PwyyAVTNltCeLuXJGBd7/tRwIQamT
qgGTl2SsEhrXAwYjy/U57Gi6HbYEPh0p68nfme9OuoAsr6tPyGKIGpapVXK2VITD
yq91LNStsxbrEWEJ60muYl7KMfIWLgNFJb8TSrHMQVoBU0nfkGRA4UFO+/ReXlWa
l1Gnhk9voqCW4+Kt+s70uUdkqSe3NRCdxSEvD1MN9CWo3MWatuvc3cqz5mtXzXvz
Gj6mBHmkoztFKD0d7Rpz+3jUpt7TceD6jsM47+BtiFKYg1uynCPsVmtrcIu0KI4U
krTUKMl37ShEaJTOoimtJxbHwryMBCVN/ljmkLNSC2aTOuUXqy3Krt4rt3K/veD1
5BsxW2F43eKcYg5OOdTHgWrH71/AZRiPLCR222ru4fSNoUvjb8XQY3jNDxa31vKI
yEJLot3OIGUxdqoWLQMP3yuV5d5O1+LacSO2mudRifbv28+idn0EFCf9Ze9Z9y4I
nfMPRPigITndX7NKM5s15/pwWEcRURLsq9nipMNukSm9qmE7V4XGmMgx6T6GXPfL
x2eHEZyAMS75zg1Z+4Xjc/c3InKeEuiIoHKJDdzQnFQFh/wbVF1Kd8iZa+D+LyBb
K2IxDxznbfB2OCBRGyq87W2jAVjnYyRNfbntaK1P69Ri/f3ldh4U9LNCJMdtLjiQ
XU0iNNPQezaY6h+gdBVBj5XwAvW1Gd0tccfu0UnehfkU16rQUlHf1qGJeA4WV1uP
1N6asKIhTd606LLGHLxfsdKitePx8ZhgAz15eCykMpDOr4x/tZj0LfLMzbahcFGh
RoZU3gLE6XF0N5dp5UfVao/GWwcmX31MtRrc/vAfWi3MNQUrnwFE1Iijp8kKwlUA
wv5ca22aOFU6MaZLHDwvBouN/M7m9y+se0bjtMcRnMM5rFXlyQ3TAur3dYriegWq
yRL++uGDjq46IMA4n0uR7tOk+UT4Pq+v+kj/DVUGfd2K93qV7aHoMNkC/o8eUvt0
HQWGOdZMVD4avrM6Y/rYLhDz1XHbKF6wRJeVQpY6C0FPpUHX1ue0IF/ocPUYX+ZC
NyLQOpZkQ8reDSckvaWE0nDLkr9rMQhaM+kYFV0HfZNrOIWU5nAMhIccQE7SV2WE
aenSdzcHj3pbf5Qx7HL+2G0zxqxK05W64nTb0nVjB0V8h9Rhw6Y1EqO3v0qWJQbO
vAKV6U+wjyltdkH/eRKvTnswjE+kL4SX81QwREmnnnnPK/3/0fgYNEVX6dTbkae+
weRMI9w7X2YA53fNimr3dtooGvuTT2FgKLuAPQPulh6fKbhuEwVkI95YatMkq8Dk
hnF+N3g+7erGOnGLCqDLYhme9M1JgVjc7mBZPztMY3vIFmP8ZM0EP9dnKCbFCKWa
Th0qsFKbUMv+KSG+vSW1UF/8nwAsyyxuStBPFRYzAVP/owPDtX36eODk4IJFGKDc
z82YVON1LUHd+ZQEPis4qI9vUrcnh0JKqA0l4tRLP7spQq7OshYr2n2y6xBHrFsS
FxXnhuwHz903syJWmmNWCEQcqbjJ1yD7HaCOIihv6Ayeuq4ryohBd2GblBcOCePi
Q1CnIgEnyhejdMI821x7V3wCNQYEBU5/VwutqUYfdCka7EHffkjS7gCrgPUAAzps
/Mh7ugz4yTLAyPqA8veu9TZSuf4aA0tmpm7f2h5xJLglb8fmInM4wDFEAw55sJHZ
LE/t9DJ9SQXm/IKD89Pbmmpbi2fTW/sQfpbW/LBGyahOITfyvKQe1qiElpe9ezwP
+Nwmefdbr39xBFG0VAQQho3qrFqA83yJmh+HCXe4EZk2yjXwbdL9f1rtqXjkGxui
fn3qHygQYL3yF0CopkrJj6oXqHFj9v2bCI0sQWQ8Ad+boC3NJ7BEqTPB9Bn5h6UZ
euLh0sMAcGIiN/taJZ7dzEA6h7R4rrElvy2V4Vt+N0sOB4c3EnlzFSGk+uXhzrof
4MqPoCJkyzCXeq2fo7lxHEPscua7v0F57zMEZPpS3JXjVDcvQdDOJY7f8uRreAtI
XzUgi7SrMfRKqs62PAKndcXXP41ZFU/BGsaQduE89UGueNzdLl+YiGq/Hx+r288z
uAoz8GPjyasu+7CoxoXhlyDdlUv3mq+GMa3PNMcDL2/IySscA+QspVPUszM3uopW
HXf8T5LYfj9+bnOhM7E7POGoanvs7lMo49i7d/dlnKrM+k9GK3hak4NlGUC7j8RZ
1RvdKo9sv/M7BUD0RbRhQgZw/A3sK7Mu9tsX5jlXmgjziajFFZUGoIV6b5FodVPy
ftFlO6fW567NP6xPWWtKUCUSwUCgc6Q79Hq/HBBfGLYYNbiOosalBCDi92PAfx9z
VBylebIF1CyVqInTU/6l8Axw5+xjrh9d6U8/qk/R0bahiWs6xllaZT+W8AY3or4S
nSUZjuILXgCQp+/zoQPazmZ7JX/BeWXE1WKvw8Gqv9xX2z0qdSdE0tdcy3yyXlCp
AvrhlnyNGgeFEaFc3fWX3Mood2q+Eld3i+n7QFz5wDN0RqFMk8eQrTiU1HTsIbVC
doz1f+Xnp5/UkcrhYDcwuLpwXi4W8L8jxC657m9kSLFrMt1X6+s8qlGS2MUgETKI
+g8e+zjsNuQOmoHtqM+xRjfv4bNwBOmhOAzN7yRIjDhUUPXFWjXlOrSxAO927UeM
qg5EZ3FcWZ3FP4IOZ4Bxiv8JhMgxzuh73Ef+WxhHdTooXb29qjE3UnEW03hD1kbs
e0ctUIvSo3FHQUaETguq7rjXkWzYv/hElFUwoetMxPyqwURQX6Nx/p4tDKT7m9La
H5AtfwzvUnplahd/TqOEvHUQv2Eu0Tjd+9F1730c48U8GWaT+agfDAcEkNGsCk8n
N9NcmmqxDlHgSXoYkyLGtyuIsU7lXmLmW9BV0NGekiBMcC5/elYwasz5E2V0XlTh
LKzAEk1d3+59wwhdAhZIA5/zbiRgC8X17LbvZ3SmY7vPiypwhifrv44gBmTX5YHx
bj7fLudJvp/6lOSPbz9xqv0JMGcBAYaFNfrmRl1+7uD2Qnsa21NK4c+uBZdrkh57
umfycEE1GDKChmLtIDQaJlM+Ho06MU1CS7caWvNkUkmnZE9ubBGXkhAyPI+t2YZc
eOe1Ivhx3rXOOB1ru1svmNQBUpuSwxV2J8DO5FeavA7cZ3v3Tn5RraeCXOnTs3Nq
22xH4Ib83im1o9tgDVQVOSaLFc6frax5Fnt4A2BbvRWM7fUu7l7L1r8fvbWlLfT3
Q9Q9AsO9MM/OfW7YIUgmbjBMBkW2UrYBt60Zx9uSK1PCGsSrix/74C/Pczn0qG/9
tfX+zynJrScMS5c+mR3sQx8L9L0JEXwUFRlNqNEioXRnk/Byeww8duM61ZizGaCc
ZwcLzIAjaOu18if2RsTiEF3E0dOBz5AOjzq12CGWHcnZy5xqKrIF52CSEinD3sy5
jR9dU+B/83YSitWmUlgF6Cn4xkPCuhMtQVx63bOQu/rsxPUxDa2LTVy2ZdMs1vUT
weQyl1AylUhaI1MBCJ+bstOzDtYtnXLA5m2b5yafuBAYePxQgf1k27FLp93WDkZF
epxYgacO/YR4B712bLL3mP2S/Gzq/baxLqicdWW269ta90JsyZbJC+6KxJVtHxFF
R0OeUbDHu2Ve3zs0Dg1jMNSMapYfqRhDzRtnhjc75gdJqSz1iPVfPfO+QLXFCLNn
Ny3+PEsuBIPnFEIZj/bwl2JCGGGDL5opFcVRY8FFYMSLAAbVzypWBqeaavI6/3f2
PZf+aa71GPZNEL4CcdgjSSNHVZIWf6UpBk3FGdB3nxlGQZIKOp8uEbWSzvQQXxEo
BSm8mRStAiXaZkri/akbhkSXzsuvGKqwkA7d3Pu4yItLdPhH0HMff/lvR45P0Gz5
zHAuh4FdLsUpGfMwY836p0vIBrZ236+lvCZw2SQwgnp4OV9063Z+fvZMK4Hgdqlv
4sdLJq8TiS8QpG0Ni4bPqygtwfCfi2AJniF+EzNZlFEfa/tZSyNWKdvJH4TfY/kK
GyPIUfGUz01kRA5VfeQIJYlybb89rfw1xb6Tc5ljQeKx95vyhh3YarGHz/sTjeSh
yD5L85EqAIfQ1KolSZjgh6QpOjtEo07r3Y21eBbOkUsLvU5hmZ9Yp579VAsiYnSr
Wvh+UVJjS2zT2i6xkNeIMyEuqp4C4xDAr7aC7ARcVxNyh2KNSoiYWb3O+XBNLIMZ
HAWJqnYaKLamHFUpvm6P1ZKKSNv7sur7CkhDBX0KaThVM2qHAfXgSBncCC/E0eas
cKlcUGKF7zRyhUKbiUJdfg/5UHtEk5J3tqJ4JlGilTm68egbhdTlyyhWeOG1N4ak
L7KuloU+Gee+4FNDk760gs63WJYKj6wEBRQUEHP6ZVUiXbXTBil6YM6T1DiZvvGn
erxUE2J5M8YfAUWcx4e04V1xAMp08Fz33hhmzOGIbRqNfOqgEkQpEGo3qQcNE2H5
5uWNGamXPqkO1v0g7nzCJFIytp7vQE8JSu7nb+zlIFOuXRJEnn76e1akvBPUWxQg
diTDbAmtvvumR1NzSVmXiXNGXie/M6PwLEYtGbuCIyxJ3tOGOFRrA/gVqa2Wrn7p
uQeC+WKTlOuOQteTju5YUjuYQbk5h3vszN3QDliwspjg+N1R6pBIhEFV/wtrKFlt
2jWioczKpq2mk8q0ZGSNyQU4b/6VUIhsbHIevduFHUPJ5YkKWD1G6cBOYiFM7GL6
5yOLNWhSzcQwVMVl49xHdIB8bZnzlQziOXpIdpskjnLngDhFgIgQR0RNgU9svdak
/Is0fHn4hkH24p5h6ziGnFbcw4ovGCPjEB24TVxYXbPQ02N5SbxXZQslmULCVFkC
xgOlF1vAbPes52kb35IgIWmrPgVN+kTMrvfS1e2abmBoJJQj3Z+Ok7cMYWSzVru4
kZbEysEbWOcZ/Z2OBjw+GHxEuZCSObzWfcOm9cyWHG+4UoGKRt6ShExvvv+lt3Mz
94GwXAl/yITqz2fvVRGRtOu3aS3v7auWqn8RYX76eXI2gafDfA208JqklAHHO5Go
IfgfFcjYdfa09E0wjpz53KuVf6dr0XHtnFiyx85dLtXyTpGsVhYIzJBR8K4X5Jbq
CosplMgfhBqK31sbFvk6W8VTWoNLLx27L2aMpWbXC1yx5IqaEPwr2LS0uO/6i07Q
2g8R0Blui8SohecBsEIo0/JiCIMWNgzYePjyh0DTBgdmBciw56gvjFbry/rL3UcU
/xrvRKIw2gNg9suDA+zys0YbLsaMQp7gXJ7QDI/fP7o998ZBBHTtBu8WBXRf3RgK
82FbaXsO71x7Pny2V4VMbBjR84YxhwQgXwLY0kggAPY5mpiJgIGigMbsD2qaCZFC
3pwMnTxnzM1ie8AdA+Qb8qWpL+Cl0T0bfrF1Vsa12HFgZw5inJvccUSYgaV6hcff
V5N0jct6VUTIJG3odvBfxL1MzEVNutosv1Bar5bcv9W4Qq/B5mjymHS+P/xynlKs
mWRN6BA/Y4jFMv9x0n1ViodATdWR5zD+GIDKDz+UwzemaHG7OEWFKotpps7WeZL3
a7nwTOj5v/6qGG60HYh6F/984tC5wBGwIo2DTaCQ5b4v8I9Hi2gQre/gwl0DGzlf
s9IVbqmSoRWE86Kx52YzFLJ4+xTZAg4xl7PfQVvFeQWefP4saH8hA5qx1YGXUZRv
gi4/3Bg1TFpdKhYoHblIlaFq38ppzaA3ap/kgyYIJ/oWvirgrESGeNf857RMKom1
g3bsw1g8aBZzhMdyarwsUdWjUHjkNHSMHcvEysrMnvl3LpyHhLG0XdJxvAzoSGvC
IutPrGuuBWZ87P91MVSME6S4F1i7/YgstGw+Hy/JQEw0QMxkN+Blfct586rpT0gL
Rsyn+6mKsWPHWGPNDC6v6EXUcE9UeNd8ryrUwvqDL+zQJsqNXxFAm/ZSqWSwStwh
pRymaWh/RCM/yh8kforpRkfSnabN432VpfdgMGY2MQKomFh78gSdaqGi3163wXXB
lNpGiovN2dE9PJ4wdRi4VukxAYe6PoxYqreeWZ/Y8N+O6x5LLb79Cly0VhnZOjz7
fLxVTgcY6pIC/7EjmQDBRjp+RtjI3xSHk1+B/LmpdnErKcfwyBzukeXzd+03VHJO
LCxaIgt97MJYljBXwa+cgtIE0HiBUP+XxSwTgl2eRQuXnnzMsRdKVg9r9TwMAwJL
Q9ikbYKv/Z1gUcZi2BNNJwndnbwoIG98//LuWLIfrDyG3KxGfc3/iU/zIB0Fglcb
janIcS/yI0ahUUjHS/eXnHiTcgvPjMNEr4pBF4LArxdPtfnBfP8ONOWfnZTw+TF9
RAJ4nFX+0m3Lng21xfDd+6Opz6lzsuON7zU0PkKW8fDVnHVkOPkwFTrabEnAkhI+
Dy4kgUHklsQz8vTKQs+CeD2mtvbqefEOEWhr7NJakUT9hRv29d1zhUeFtZ3Z8zzj
TH16Js5kJ+D2sp3KwYV7lKtQKQw5MmoyrSbgqKnvOKA8kI1pGEiFv/+l4YQxIOx5
3ctkH2Gw5bLczVdGQD6zXbQfxoefQQ1hqHErUaMmD75gKl3M0KPmyxDak7OvqkPP
lVEMd1yEU6hlx/Gtq4Ld+x6EjMmu0K4OlWS/jA3M9dey0R625edizmoG7l/ha1yP
1xFrv2b4UjqrRFI2Bx5oxR8E18TiN4Jt/EDIpP+fGszDIAyWtT1nZ+Jdo8KyplGh
Al7rHYdcCPk4/PTBjAgPRb1A1JGl/3I7SKqBVUAW6Jvq2HvAUqToZr6c2bt4Doaf
TX7/pmCmbYaSKW3wnaRL26WIF5D4FvyePiTVPBQcWu/WeTCUCesjwmMwwTTaEUe/
gW6LfMQLhn/50nzzZ6CMgQZTwFBOsPl4CzgmhuUIL5KR//1AvZEe78v/q2Qu5K24
BCnimpPUi2/rg6ao1ojao1YIipgyLQKpVOXrRh4XZkAAS3Q5qC6ywecpWmG+4vcX
1uJyRgTBe+FnVx9ukb2uv5qaVzuo7PzChNucavPseASYiuQVyfJxDPPhfL6wDEfY
zCLwM7uSbfZKmyf2mnW0MC88nEOZJN6K0wK8ihr/iKGHu009HwOQfM0WhRQQ0TsS
/ZriMbHORTT4AL7XcWcmg4KrQ7dXXhE8w88NAhLlHieYRPFGIIXwus71x5OyBew5
t+dT/XIDdxZmYOlv6q+nYZLoo8SKqrHJYUheY0093p8vkLwHgE1yKpm0C8j0GiFr
QfW8PFcJCfBiiPIC25f+fhV9wv76nDEFeISj98T6PHicvHwOrjgo1T5OpG3cBqyd
UKpmKwnnxmxwk1JGZEgF6ZR4K/OFfNHd0TCNR/zgqusgHB+46J44XgUpRxqsLzZk
Tos82e8pn1O9OeQmbCRKTU3OoKmIeoDpOGR4yIy2h/Kt3ylh1PlseyFGW1NzDcdl
XSDIwG3F1bQFE9j1gMKrZG60QB7xiUIZmHYloCJU8FqAStQ0E1cYO3U1Td15yKg/
cQqLKHdf3IS591gtCZyegfrSmgmD1WzVls8s8gcPXO+debdZI23Aylqs4v9fQKkR
ljzLCvgI2akk88c5JcoJwy5mNt6k209V4mW/ow31bVwNbbP11N8XgzQlsFnpCnGT
qhyMpPWHZfMEXtiGsxiCysvVv1hkv3dminERFDiNEXcW8WcvHb3Vw76BoQN0OkRi
XNnZn/7q1Vre6nbYKX3D/WbK++/3uGDeWvHWEK+GjPPHBfkRg1arPgS06qzWX6gK
x97AyJhT7w5q0Ntq0rmSM5N5tf62a/rQblT/qwZxBeqr5J2lIfWIfaI4s0MMsFeN
eXEjIzRmXvDcdVWtk4VXPJ/CywDc8SmhLJkH6GNPE59rHie/jXiol6aTQLqf9xgL
x3T9Ommhg4H5ROXET4bQuf7I87o8/OcwhL01zj0x2I0HRen8pKcsVDsBdeVC4ToR
H+KXSCfoL2ijBIpVVDlOr3Lv3AkxeboIq8+3MmsFpHtS6UFLpTFkTkkOQWAVCJg+
iMDtFN/61EnOhSPWC26aLf9HceeUdEYpwri1FliLS6s6f5zHYE4IIqT/KXT8xPt1
FWyleGo2+NcaP7tCdD/UXtvJoRvN+/zmaVFqLeVErqsmWhW+1EBWQBwAetE6HJng
DMPtOCL6NiITmLbFUsV3CxEkv97W368Zg1RA/UEVeR/URoMiAKa8kt7swl+L2qpg
4i6eahBO4iFSWWby9F+pt93yW1DXxJV2GHYfqGdTvlNht433q4QFgDrgP3dpStck
6g6oH+OrQSvln8cCNFuo5xQidsOqhE0UuLmY8wbstKiHyueQ/po3hykrU9pzjjvH
BgInfXQSApiPfkr7T34vOioeKks5ovc+alyFZzQFjoE2Jd9JI8BZKfWfiL/jNvJe
r9se9jxvSK003HMPTSGpodbryAr5MVtocvGRjdTgsVB/8OsKgj7WSoLdaYeO3LXn
bWacQDISuLzubPq2ArMWoP1wOECKwIYgfWzUXSEmlUHCrgyqqAh8Fg/FSXnb3n4D
baauCGsFy3rfnzQlJMhkIIFOayyWOxvZQEUkP5aL3sX3QNAUm3QwaS2E3t17XWig
it6NwpmuoDcrA3FnHrJD83pVqvHoTWcKxzEdttT+jsNeRgMnJOjuMRlC2jXqFOjl
w9EHHV6m4bDnE3BHa487ek9e7muNIqJyf9p6sYUT4vpRn4e40Dmqn4JzReE0uhaH
ewab2vuqXRVGi1a1kn8uiH9TMup7n2o6VURWYm2t5CJWbUzrcHgqaHCfs3Fcczia
MYiTwqHTQiv/OM5IDlT1LHElBby7oubsKo1Gtk6Qbqt4UuK1JiJQFBX5zLH453bs
bE6cvjEjPAqJmW64Y3HFgFrWORiBfk8TG0QSx9AmAIAYMd5sPQ/ixs1b5p/WUwuf
RCXyDJRuf0ifMhQDqGPCUM3qbVQMTrhXHXT5LKZkvPKh6gBdfJmytHOeYtDjPoZl
SdPMft166NAzK8RwuBT4Rbkl/CahpApdv0uAdffn9pgSg61DaEE1NA194TG0k9kD
8ooPuHxmNO1nsP4snP/+DZZ8pQSpW+DezlsADgpneT5yuICpfSZGF+9i0DB0iQ87
J93R20G5BEFE093MC5QFtrJADpKG5SMp10h0ktBi9RATHQdMMd4p3Q3M1jCkfnlN
JgvxsJsfVxCs9b+fC8fMdhQ73bq7DJgqtVqk6x8aoEyNIttgLWfaOKHMtYsq/LnQ
o+KgwoCiI15Y61cm0JOQS6EW9/kZCgw0nPsHCLp8wOeZlHSIGVtgOeZTSwlIlChV
+gxIVES2TLNGdcJVQ25QO1dsrGvU045UXIxpNyKLocYqfZ1CrOSdHUNvK4WH+WYH
yW9PTrMv7CHZB25INCFIpbjBPob5e0SyYoImhiPCmm0gsjwUtsqXLg6Yc8vcZPg2
sUICIbcRrLXH590D4XHXafvnCsKGGRo/z9Xaui7nIFI8Z9FUP4SlY68y140jQPqv
bEDZoytnCPPg1pmHTbZUS+A8Ry7QP4zxU7Di66x0xpbM+sJiUh/NMtoMZaGAsg+Y
Qarudwhl5Olb4NxxZal95VSmUSThQw2jlFI1D/A1f4ohKsnsLzgJbLtSRuvBzssd
AF0iJQ9QRMH2g1cdQfWAu3Nkn3uP4qvmNVxiSpK5huRXTa6ppywtkwP/Ql4q5Eo1
HW7PZafHTBBsAH156dKF99FHm2jBJappiTLtpnWwTl2eVuYaeyZuW8Dp09+0ziA7
rbmBrWUdB5SeJBgui1kZwITyCw8pMgrBLs/SHO4aXPrO9DDD6M+Ecuxee5eVpTqg
t9xD+18e31AcK40PGDlyWpHJ5Q4ncd7NM2+aFztaNgNhIksehO120gCo2MluNHbC
p+wT9HjRnO0cs9uwTekcEOCfsVE69QROe0XSTdnwxkN/iFS2Cb5AlUX1VIaWfmcC
WlK40SXtf8b3bQGxlrDx80JFvMssb2mM1huQqmk6FTyGQ6Skg99gFvS1ITfhEaJW
HOCH1BvZdVAM3dIRgDdWtXByMmfJNkwBpOZdnRe5446/1n3p9JsKg7C51lGALU+K
4QcGVR8tTsbq5gxFoA7EOOoK3VU2Bn+s4qJmTHmOuuBva37jqB8vaSNOlgzIoKz7
QEdLpztIT1EF1eZXlircp7F4DOWh9MtL9CpGfYTbnxKKqYwVolu6T1A/DZGIegTa
eHNhBvja5PF5+mqvKwtrcW0CFQEAue9zhrLNLAM9WrHUpmv1sU98gLCcsVKkQyKv
rezYu30QLGz5pXEPcs9urW20VClXbNNradcZ9jW1PcVCMCIpn/p7fE5rXBRzMWzw
cYahYEA2JMhgJvKV8/nL3sJ3Y9BCygVVD9XS5CG3J5Z7LoTCotAGoopf0ueuvwjA
/mo+IUDM5oP2KgcJ3470JuSkXpMH7OKiX3TA6VepLe5AZMVr251WhEJGmYS3ZaMm
EFmRgWu1zBh5aoRczY32i1mLDhE9LBRRJb8/NzO5N1oButEuuSFv/5k0RCM5kkUE
BleD9URUOmL9sGCbTo/iQkSrGcBG1f4Ss+4bOdPPm5I3iXvyTvTHTvvu4CTeCcoF
zoXN6KV0LiOwJBhJQjjWYpEtcgPMLNjXIvL00c886WoEafQZdbgLsFhd4QcMA+E3
g46yCiTq6kS2KAt5RncRInxNSeavXiDQoRtmfSKztnh+77WRFECLsZVw3OV4fEHv
dJnxCNUZqnpBPDrCmLcOuCkssHDVstLmDjnLpnhd5tibsu9qEnZFXA15jjobcT8y
3/Y1WYN7LaRhEwLY3emNCAJ5cKfANWTNlBd5+0N8uIh5y3o32NPJ7qqbT6xBYe8q
tgpBOBPFOwo4AtiVz8xlKvaedCQlSfCz0hF15uHsUUJLbdYyN0sZfKieJBDOASJ4
U6uZxXybbJOqNXAo8pWWHMQR2CM9Tn0pe2F52ONpIhOQuLQBy7a6ZQg+bhtAs72V
uILGZ4O4BTlW/hEZco99Klia5wZIgxGKztdw9sJVgvmdMl8y1WLWXmyqIhj3k8iu
Vu/JHaZpmWv5PWoZ1RYjV/NqsFZsI9fjzVNK62eARDW6KskWmE8Q7RID1g4xgNuU
ZZ1fDiJaprFX81jKVsca0Rzl2xeGQlr0bLA6am1p5VyfMQvZwd9fGyCAeniZd770
+/niyx92yJ/lTCac4dCeOg07JnfP8YjN+ZxMUbTqd6pvffb1DX8N+Hnkz1CXjXYR
I1EwsJOnuZhIedBk6hhzf2/kF4oLOnIuMDO2SstbWNXmI/kvW2Y+odCWlUnPso5y
80Cg0rsHo30QIySZWDRJHGk2Nj5RzWWwpD03tqwiQ78cx+pVk2paikvAbpnKMDnU
OnjNz6u67gjo9b43sEzRrwGe5Myq30HR4Jh6uTj1+J2W/p8Rm2DZDygktITXrhWZ
h8k/e4nivuXyS+3LAAps4F+CP2vjHCLvfZok3f3Ej64gdY86OnG19NeTjLXZtzSq
cG57H4HGRjlA7HOhqKsPPySEMzjFMva1XHR4xwqLZ1lB0XmKT88vCLJuPAEh2k1e
NFOKfqG/E9SR3u00nDOxQev7U9qQ0VJgEunlqYwKFJYxQrwtokViCriAklz1HMmb
AQUU/BMi44dwGI2ioQa66fPaRubG4XDOceSKdaw1jlFacs8Z37QziV4kJyrV6+tU
IddIoAfRasBmRjQtY0P17Inze3zUaF57eDeK0nTjc5X8rUSxN/kbEu2lrHy8c/9Z
4r9lhPzyaA1F5k4C5iRWKjjgYYZBAmR/RqVb6IEn354tFS/o6zuc2cizHgCWq8kA
yLZEJoO5qpDKhy+PZn7A1LHW4Ot/kIiTeEy151OHD3DA+5FxbPyAMXB0pDdaG1gy
JQMhyfWUoMbpDTPH5QQcTVJEOqyIhhqU/0QZ57ORpA7hVNrJBOTKT4qT9z4M+wIt
hhvhAyjmQKDgx4j89+3XqIJoNHs2wCettdvNfsDMffaWAHWMA/81tE43OKD54tmK
s6IZDKEGSr5p+22LxmIqoqY8NSUmUngteoNUBtiyMcd3HfKr9UFYgGTIJ2eT1tL2
henezzNTmrP/8qVk6Jw2hqfqu7ujS4ffONiMyQJ99IR3sOb6fxGwl/AzOtkeIz0F
9FMYOIxlcsYAgnraMfOe6Ik0wvpgeknHkpRxT0XC1RL/VAYLYDyuWpKyPXep+sZC
PvXOyqQclgkddQ9JvGVDeWxFKmGyehbQMzZSDZJyF0bAJW5S7B/tX7HxhLdBKqMs
Dg+A/uvb3NBDSNPbmAH0VsV/bjLxDhY5urQv14Ea8YNOVXJLWEHMifsRPJtCIqel
oDGw29V46mO5Li7BC/jc1CU0W1Ap/TVJCtIJjtp0M6apPcG/txbnD5d4cRIkP5L1
WRXNz3QWyLsB/46rDY9vL3dvNfZsA4yZkNPiUn4tULRHyMBZqe/SrE5zorMY2DmD
JMGZfpqiYWkk7CB6OJNhH8pxsIqimKs2RajL9VB3J1i1qZ4MB9vT1/5fcfSzqjiZ
ZzgX3blIHTZNHoDKDowJqijGPV3+x5qHcmNo1OK9QZGOK5phznt2VcS1pJ2whvz3
YUakpQKAfrXdo8sKM3krjwvmiDKzqFGK5HVs4VridkZ0SwpLynk+YXlZAuxJmQIy
SXgwE1V4bCvMMe4qBX1h6GcqBCCtbKnSs/IIRV+klalbiqUkh37jtSGCXCFejW/o
Xks+MTq2d1GcSXn6YT+Qr59jPJRyClw6Su6DG3fgKhu4XC64nz8venKjGntuGs9Y
z+yNiSrS+OzVFTJiQ7zbUcr2kUHTYqec97SJ7ltLOtduiVVUqKhHThl+/FRtM482
ZeRnXs7tFJE/VnbDwBsEfiEREqi5Ck73Jj9YhuZJd6SsvPfE48jj251FxulXEQzj
FtwfINQXVgwBlvyMekb2O/mdCGym11Ka1g4sBNRc325JxMaPozmnVpQYWVSlZ0M1
yd8aSImWUiR9L+M29AsSm3U8ac6vFSDxoB2l9b+LmbgS//0czJW/wTh6LHskVehb
NqvGrRgrScxbD7RbdcgzZiWUqlxe0KLKoGrUIn0ifE/NOOmbYV+iRQHA9fwmT9oE
DLbwdSaM34RxZ2+eUYjVSVthrKdZ4gZJMpDI2JMas7je4EWeweSNCeNWukrWt66c
iSL6h2Onl0qGyIEIgwDAhYYYdKMYtbqnimGFYV974XxGK6KnsCFpgUh60Xfq5mvK
4cJNI1+WIqvikorNR3W6yYxe1pcNXXzHM0k1gFp91fEDg/xSfQkKlXjHtCSrVdJp
6BzbwGsS6dFXAOMg3/lJp6IRQSuv1OZKpMPhk3ZyQCXkBRwruUOd9gV8gbI3O2kL
3QRlVYZfUeuFxVW0MoAcUlsEHdydCCHSOT9ULgALPn2HzrcIMfYZBsrqP+BRmcCr
NhYzCsxIF8SwTB6paLxjDlRtn+/C2oMLYcSDj6UETNy5lYg+8l2Lfq7iEls7KfUI
4c0mPbGBebTmzHBZvgnKwg5hqXoJ3UJ6G1vPTVTodUxhTj3/4lgKfAuBQ0s+P8WO
27JS/MLfDXN/g2dSOzqRucBfzK9U/3gOniP28SjWA7WnAaLphuQ7mCB4kgG4HceX
6Ae1d8g7G/O6rcrRL1Kx0g1PuQVVHXD8To4PbO/3elGoiAtHQc9XouxezxMoZIp7
gHH6ip1YS7TiZsre9IVMlr789wC43egEbXce2qJTztEm7nUnekThm0f4c1Rim4nL
tvZBb9Xd04H4/tUladZshKe9heiofK8zHDGFVr81VF6Np0k8j+qteOO2myjvIdef
r0I5Otiksnw5O/m3Mb7MaP85/LFTB9gDJRrQNN/cQSHvVxtgrmlpCKgQQ1GHTK+y
KzKWQ1gR9WO7IrTNn57kvn5wK9U822ixxh5S9zxuE6quPQMtyN6VTwrYyGX4liGe
wg8StT3zOg/U6orn+4OpVlHS23e1bwwjZmnXl/pbOUnO7UzCK2D8HmCN35rZ9wvX
3ZFlHUXU2dLr7t1J8008shENnNpgbt9w8XiZIfLxTrnAzSSb/WR/lRTI45vvtTMd
6cBS3VyT6Y7l/VleJyG23Xr5/yHZDXFi4M6YrkBr9FP7+jH+saaoL7SWpjgEq/Pj
rtYp3FxIeFQ4II1GhecUKPdaZfxbHEqeWvkM8UmW29FvgbNk0MGn8/vAk18FyiTq
DKkJ8ZzSx7GQvYjj9Pxybx+ssEG3vLwbE8YAKAW7zL61uKP1wJPtQJs4YzjTUQVe
TSxc4ooFKS/F2DWbnYzVvQVIprUTscf36x4AIyeoRTkAJHPu6S/tU2ptSpvXQco6
C/+gQzJMRIHIsWhdBv1b2pfeCckM1MBgPwxcZhPvAgeIFAkmxvTCgcC14ZiNjD4T
n5iWB2Ee4tUWCpWZ22a04U9j6a9DR4UrQyAkq2lvco/nE65RMaHaAQaGN8etjAo1
OfgpqiiyoVMFoanT9y5+xXtjCVMtYis68As7sDNW9mXxagH7//EiUVP5fU0T09zo
goJxSq2ZpX+1iYWD+NixcDFiFioegptdjHtLmGlioEJ19Wj2v4vFwAXAKwmqqmUC
o8GPFHOBu9c4Uttplabs0Bp00CzcwDzTL//NhWOnbJuw48QhwghaqxYDsy+Mfddy
5w3PVu+hcqva/Mqsz/gBWeNTMgp6sEZKKLhkXELazH/n/5GiM+pnHyOA/b26XUWI
89FOStguYINBLE6o85FfhCoXDjU04lW0LroxktBEn02tp6DKUk8b+zM/ZGY+EFxM
8WubpN7XkKklEEmpOkTcNfzZjW3AN/Ufw439QvAaSlqhMUUeqfP7Umx4OtqOkx0G
CkNzUcW/Jo58HHd5ucQ/9uNwUtRXr85auwiMVfjpDLSY4jWSF84SMac/2PtA6NR2
io7nfXdrt7pBHp40K+Zpzg5pv+Um0nRvgbqerPa73EGeC7BJUnVCKME/UViZgST+
mKIXJ80u71zpZ554hum2DH6ZSJKyYZcBIIohjMG3aEQpcfleyd63YYZXaZtHH7Gm
W6ydgmg16sTRLRPoRoQJ7Wxrp7s6BPo74tFUUwb6F9wkJ/KzJ+HbW9Pke/sX2f8u
M4wAnQgx0RiJSRgghpz1HDEOiTbAKm7uoQNkq//i39sAxgs33eLv79sL3qApNXhE
/ogoF5RdtIXc8gUZ2Lfu5H1VGu22WREoeyhbWpHqSigOhSvoVghlKgeLREfo+iBV
xYeIjVr8tWB2j1gIxUR7lUQWcsCrgJr2DZUNBWViLWZYjhq4+y7qksqIsG5H58fn
jwEfdqdkmX/vRSci2lI359TDgCSMbm4dfVjs62+pPnlcmncELajOVwNoEYPEytKC
KXLRvfq39nQJeBOQfVNdnf+Ep7XIVUiWKS6pBMDfG1y14SYHJkFtz6eaSpXHDlOl
cuYZo66qKU/pcetKR+llLBGpvRAnttQpe29wDqPlEEa4yamtoQZ88i3TXQQxt+9l
LX4SDfE2jycmefaBN/tXQhg09SjIte3sdgXOzfkfBYeEp5GM6j9xCLFWA4ivvx/V
nw0Lhj0zwfyDcAoy7fbMkREmLSBxHZIrVNSLSVYpPrB+OSuDPkRkuu65Xw11tkeZ
0X6Xaxmtt8bbxNP/uJ8Ix7FlStDdnGc+BjCW0AvpB6ykwfVKtRFis9t8ANfPcACk
j7CNpSBiGVdhQ43m609KlcVIyGF3bNFLyhWvsCBC7gNIVGKr4+HzKVeIrX5IAK67
2upVMSOSoQoD4TYlA3R86ZAP9DiBkBmWY81VbAbIgA7A/Io+xB0xnazcFfAUG88z
9kvZ6M7wMSNhUB0yaYaClH2coVjD0r45EyQb30+nh1dF0yLA+77P4xCbutla5JCh
Ei9oDL3NiS91KDGNb62qY7rjNRiHQBgnx0LOrJTibIgnyaPVuM7ZwhJ+TIq7F4MO
ZIZdtHjc4v8U7GGnuLYwNt02rAAaJ+ZcCjqWlBmyjsWG/kBUU+n3EGWCl5AZ9Tuu
LpKDktdEa6b8DJuifcTPhJEssTDlxztxwLRYpMbtWFDKXhPryKKQnDo4jE5ZVQNf
2sqjFpqF+Q5GZgYY8nRNXkoE8oWa+KqIuJMH75PpbU5YPH8Z928IBTsiDWOPBR7X
hECxhbdXJGaxOsO/+94VCm/Zvu+LVVDFAkxMhZs2MQ1tR8t/d+f/ADAQ23CbNfpq
pZseaEwyL73N7rodsy0sedu5sdNX4bWi9Dgph3WCMKUjg10NRZY5J7zY6w1dq0rY
RKx2EHluFzlP5zNtXVcdXxGoSjKZ7e/AsDKAUUYHD1jSKSLTVeOlhki4gp5HD4hF
NX5UmtwqXvXNyNfZwklww7TDct7VGdwQdv761adCKDq8Q3tcU8h7/FocICw5f+dI
xNNBuu0XSuz9oSFoarh/fN8fJeAe+zNx9ZkV2b9KBNSBR+Uff9kRovTuChDRB/Xk
qBtOfNrgNn0QJ/vUMcWbbleEBmZR/p6vVbTdGnF9uJpjw8o745FoLVVw1+xNh2zG
SskHnr+VVI4/i9SYRN5pezgtwuwn/IQGDVQN8U9ZlatZY9EQT8PEqvWUSuX5Md/8
L4GsiMPtba+lyMKs0BwywnRi12LRwoT/mPqCPdQw0JaAnU6uXyqqOdaEzAJZET28
xn2+trE3b8HXnXb+hoqJjYcUD53wVZDxTGQzDE/ZaZEJyYQmkrhx3ZK0e4+wlk8V
vOByvPAjbU8bAj8a98jFXfkh2MV/PpdJBtaOGEI9nSPPg+pq8tBK1VT08urf6eIw
1XCv06PvsD453pSIE8ANSeAwLAXn+IhY9q1qa/czBF8t8n9FWz7owG6+7BG+dXdy
7hpS457pUKElHD47+jiBCnpwAzRBvaNdd9en4bPLdcrQkt9UfRRMmyvuTlPGg0dL
3kRLhCeI9XfPyFwtn9781n/ACZpTQCdRL0Xb+yaQ8geR/bOBtKgyTt8XUVxoWACW
o0M/R6mnThP71PTPpDWoZqnNLp2sqzlJ87SjiUQ+JG05PbRC/quj5kxJT6dxYy+o
poi+y0irK12pyLP2RiHfFbxc7nvUa+AhnqWlb34P6TUn5RFWlINbwihfnleAqbPF
q6q4dCRDx9RABWuJ18+1wIOXS4spPesQ1v/2I/lcmkSCaODCB6YC3li0P7mPJqwz
BF5wE3m6G/TbLE9p/Vuxpil0TO3ozCWWuRGo2MVyQWPyUGJU3H70rhC968vW5ufT
DfuvI5pMq7UpQTyg/dNe6Gv2e58xW86ThCcCWYlq9GSJGOZOtYDRigzqkEH4/kE8
vgUlFoXTPV52rRH/C4V/VN8Fvc4spqLD62XjrRTeWfQFVh2kY65h3qAIlOTIR5Y9
jenOaGmCtboK3XWcsBa1RpMtA0p2k2Ga0tCsQOjb90wLZ4JfnVrAL3YQ2+TabkSK
ohG3XmYMK9oraTSEo0bq7NJHUqyolpXFueBFjt15aO5go4EWO7Oy0G/rj5XGkKxC
qa4CpvAtVheCgEcmdCqu56jRv9MqHBcPc2KbHLGuu4gvBarTX2zL0v99VnLhdJL6
a2hSg88WvXnqLAhrFJlkJ9DSL/PTJM7cLaHYpHnBQh+ue7115DwpsGzan+tr2Quo
lKDsh6ykaM8lt1F0dV+5LvAwd45hhfDTVnxZJhRX7fxxnlpsDyi4u1iBQ4I7/c0x
/dJVvbhRRmzmBMpmJTsXxLQ4xQynqd0Nwq5KpBDWd8np6sQquPmBuD2gdvgxtFlY
+4F6n0/MiAs9meke0ZT5QAyyDkeAO0IRLoiL8Lf3MSBUPmdQj4TfOOwLRerz3kS6
7EYB5rlCdUl5G229xJxgvMfidF9VvY4By8ofyLUrR8AAvC6GutpZcmn53x9Zv0uf
kYNlan375lRIbmBBT7rjcIkwOq34KLdhZ11ZljzpRqWpy/xSzhrIZNDnA6u9eECl
pbu3u2LrO7zlF8NClhEZtt5kqnZ+tQSGFQt4/bE5H32yEn24bqXGM+HcxCE3nXrw
x0NbVylMuSQqY5Jq6Th7WEKrefa2IntaUIV1owX8U0t2ZsG9priOMWc0RR5Sx8JA
dXkfiWwCbitFMPg27ejBcP83jh4xF8TkM9YXso4uoMDAfqf2xIJJuxFNObmT2kq0
4If7hGLegAiouAz9kWNocMmQpr+zfdfsYjjoSDlBjPklazRpL1lEcDNUBx7rYCp3
V8wZs1w4cuag7PgRw+yUHZ/mO5uGnLJQcvJQkkyBSVWzLYPAo6JiRLj6Mq0JNi4k
2l6m7OKog7yd9cfpRx7sXQkUn9pmxgVDoCISuCToH02Yo8C6umtppWd5bUu2LZCP
ezDTd1voVX4kCcPFp8YaAXc1Qa49BiXuBhZsOs1lQdT2x9X+P/0p3dUnNZ+VpPyX
bSdVgtSP+orpUAf2/MEPuFfKh6c2+HG13ta0XF5saRs55INNaeu+75PU/bxVH00q
6Lf5oDsXT76Bx/hYwZHwrWHJBfQFt9E03VQazHiHtf1OZnZrxV5+IREWzz6Moht8
4qF72JnCqZ+uffEg+fDuVV0QE1VfMZzG+f7bzZq2Q+rKOY8nAZI7DU7qNcKjb+fC
swGzDLV+cwoeX8InNOuVUUK8rdRYfjlXd6CfAuJMj850mJyZP+mvO4LFM/6EBKZY
qvDlzpLcyWWVaVPQHVXb36gJdB6jLr7FouQSFIndlwLnw7e8d7AuS0lyu7JSzL3K
G89Hnqf+F7oi+beaOqNHZ+NXftJk9I/bsmfbEazUz2TO0KQn73tY2bxjOeDomtj2
IOFEE5e43/2BxA0IEZHYtk1Qe5oTOTkmGa67UglZoejzc3gAutMBTwY6jIMiQK3H
XjkV24KtwTup8yYc1927UsDCGRVXCL49JSuZCkPz9EaLHJMN2jtv74dgZYXkFHm4
t0o21rfRyDwAe/J6zxtg6ZC6YxFkBp2ulOOxLzKkggsQ0xuSmwYOEF3uSF5fw2kO
9EkQhoQoU/IB+VPBKz9J8QFk/rPAaESf1Bboh2Q1f1dXVzdeYMVQrD94USzKGkjx
TUGDWGPJP58y/ay7OK720xXXlI+zVot4pS/aMlVv7iOE51NqjeNsxKqrUNX78wRd
RBKvaPpH51lKykEZcc0wzsD1MGH0abVihfuJ/p4uaKqCvKEyedN8MYyP3BPIHPHn
JgPR/GwB1j8yKRcgK5VX/mjeKLmrB0AJ6Q9uA8C+htgsh8pmFFxMulUBROWZeBJK
NcfUvCfdjEXmhlfF3F8qIZBlayxhnaiQs5kH1ktKFMBQ1D8CwTiEzPwI6GhPRHm+
gcHCpxbOAkmUlDaWKweeR3VEHGbsjBKJ1Mua3oyzpUOFdme2WbYldCivJqoPN5hd
qx0I2Ax3PkAZIP52Nwqscae+C47c7g6/UUqqjp/Ev88LrNWqx2zLeXsf0+kChmQv
aKuKOSS0iEN8BkHVW1qu5mXr60SCuOVhvGnGU7GOtIOtAFfN67ZErsOn/Y3PGvCk
KL7ksLYPIpZ7gdO3mxTSmNjl7CFPgWCRvyPm8/TvL1F9hStSV5bME5rg9M2BLZep
bb32Q8rTAYyR9mw0Am8lpe83Xk379/pTBUAokNvTLR6uYMOgS6RyVq6qVtYMc9aA
p6BBKD51u06IkLzI6ZW6MTuNgfrxobRe2Bby5FALBqLOUSgCtA7xKRJqR9qBlDlj
W15LilKUQCkV50AI9if4KWUWnSBQ6+lFfhU/ocne2HOqRCdnwy+geaI+mASAvpQj
CdRQoZzU9Q7iq005PoyK/EqtXjFksYIglrIKowiXylJMXlfwIsJNLoiVynooVcWU
0IPkWUSp5R1ALEqhQ+ampI8+c0PJnPmCee3Usk50K2KvOxnNQ+noe9N9TapPboYx
SE26VZvPIetM0sFAV17H7zqU1CQjhPGVr0lyH9Z9CbHMvdY3QGWNxPkp6Wiod8gJ
d04Br0C+YGDEKvDvdKiAqpML0Ycnb0l1FgmVDTs8bSkkSw4u3yJOpaZiyWr7rFss
GoqJ41dnog3eh1f2I9DqdUR1r2sr6yN4xFuYVXrYc8AlNH/DNVBXW8Cp/Paa6z3b
mcWQUsHSit0zileSyLMGGbATs3L9Is6XeHn9/Yb4tpjfUVGl/RgZF75botPBpAyG
rmDY6Ksca13nwUxHT/6zEat2JJTPJEBAtC8v5xhezkA3W0F2gED32YFxVQbrRL3f
9oZ4KtaKB3udcj9CsiPNMWHNzgznX+O0Q7z73n637WITDZej/zhXzBYeaWN7WyHP
Mw9Ugg6ygF6iG4F6Tzhf3dpfN1/x91YnDkGzdRQGORYxVcWDrJMW4TwDQdl+KuBv
d8sDSZ/I3FaQ5fl874EJ0R5kFXH+zCmUoDV/jzVoAbJqwxQlAnxD5bshV9ls0FBG
5l5Yf0rpynaJCIuxJJLR9Mq+l1gu3I8/yGEM0Eeh54txi+NRI8f78q8sKHWsv8Cq
LPitXRUCHEUhmdTTwRJ6WNws3qsCr1A391ortVlQNoAsrBiS+sD8kcWv1yIhoYuZ
7xfGkEWez9VCvvEzl5gpTys8cViw9Wi/ntyduoZOXz4YOfVlmexfxYi5JEIt0/6A
mKDBmogq7PDbCWG/eeDkgrmaFY0uO0VJj4DzdM9cXQgJOueAQGd4fnoVRuqUwQce
8EaOGk4tdtRhvEKJS4MQOH6STn+71vo+u5QSwROu5h+GXrhX7C7OK3UdO7HxxLC3
asXMlq77nAjZ55sf8RAHChK+e+90sgz6CbgZZWpCJO/VFiKOG64V3YSgUd9QNlDW
zfrKgOhy1jXp1tWYrFL1t7ZjvVtAOs9FCvTKXJ+2FlzkcHBzP3aJFrI5mvEHF5Mm
IpAJdNtDWnm/vnFq8j0OC/BbhvXVc7MPehl7ls457AHo0xN5a1VKvV/3YIDcp+vS
KElgI9SDmsbI3MZeg69GVyv6J2Y2RU8ieM3JVsugtRTUTESMjxMEGPEoHParqoHZ
F7RCewjklmHaPg3UobzXCwY2m/ldsawOIYYdhQ5uK+xh39ybCSK7ukSmxw4u7K0P
IBwGQXoYwrtzwkZ+5ZI4Xc/xsHdQyravIMkuoW92tdmFYHrad6ViwVInE5p46+tw
dyNfbTFEBKUWDbgzk210zXDPTZbhYAFSUVW8xrwm3tZxn1TiZOKp8983jcsLRlA6
cqtJW+DdbQipO9a9Gvy1M6Y1kAEJ/gffZMH5VyNUN6sSurvc/yFhoHyokuoV8Xos
Y1xQGJ/+wjslFdj1dMITwx/OUCv+CIsuwf4R2FUgoQuMCTGWVAPYG++CjLM+PCuE
lUN7H+4CLBylDZ6H/VfNgz4S7F0AAoDg2Maunyey4hBtBadYE/rDnkj5+H/0qb2v
v/No58Rmbar7GQ9aPrLhNgpDm+mHyhlSDmnJXBRVy2uZgv4AloQkiRQjMa3DGHTP
yB/Dh1NxcvClVYqnoCTdJIAMZAiLqOVFvVudYJQqwqCEinpArEywiUY2YVjzqTom
cvj54ngfck3xoHltrFkDdAC2hyRAykwHEQ37akuGErt4i3o6y1YHYZmNvC8ahkHG
epUX3ORUcMgeEqS1NB1hMnZSOApbeX8nYE/ySdjQYqYHXdlifX2Ufo87REd+K8UZ
mviRO4a0UJdIS2WBKo8b8/VfqhhU1I9nB7A6GNhiltPFyF222lNp3HG3L47qqoUz
mWufdHel+2JLkLXTUKSNVs5rLwmv4sJhSBmqRdGeZtWHdIfADOR5aqZ4HBqbKuYq
CxGdx3zzQDSX5/LkwpKM4ExjezCyP/0OWcBpPYDVxxJzuo+16VN1d6fmCWnG3IQW
E045Ipx5gudJONc2BsKhxVdrZuQyk6/hCPQVRIOfnQcwh3oHDHt6Qj/4w5eQNyIx
/uuxAif55UK7Bk9N61jX3/7hXfF5cnsIXErG06J11iucLo2EfmkqP/ABRKTz0EpJ
HIJj7P3rUb/8k74jpOOoQWLwMVOlDZC5dceTYdhsIue3vI9iJiFMsgpVEOwSGIob
bAe0hLswxp4kSjkEuRqNy24RvMGIQYW/h3S0WV1BgIcYtcqupe/CS0PxUGiRhA23
Uoyc6xXjDGzIYTFl82TEpFYdLX6gFVLRxXnKZOyqYkPzWlKkSyN6dwuOOHf4Cdmw
cUoyprMVDrtwzc/p6CX/d3N1eguCeQy6v6zJNYNXpFhpfw6NoAskGOnwgqqhh8wE
l1hem/WrslU3H0Zh+W8pYyPEvVpgfJOC4xzaDDX4D/mNMRMYJviE90z9d5vg/kBs
YfyuQC7zR2LNG8QA07yGw6SfuPRB+pO/B+tvQ2EVvWG8H7KVyFIdpMfRieZjDe7H
Yy/6D9nCudzjplN75/CeBsmAm6LFfBWGoYYqV0GQEby1w7ucMjl/vLjPzVEfnEMH
k746yhLREzPzTD+P2X8ijfxPoKNj5Jh4oQ1tjghJbRPYsgzpaSploTMD4aBLV0Gp
OCs/LzhLIMeJ7xGLlBLXugkvXQDmQMClTd5TaxNBwuN1WJGSmGCpihB+H2bWM5rx
NwwyaPZ6OFpJ+73VQ7c/cnbcMA5n/4XuC+oUKPakP1eiIWuEk2abYvi+tgAbu/nB
EDQIvD7DVKNv/9LgrfeY+FKoxRSKp48JUSk3r5wW+gXFMyQjfgpXnyWpD6Oudhm/
EkshHXq5lDJikJkGUnZlp0zslZ1gF95xhJcYZi1g1lIf0DBPJhD7RvlJZz94gdL4
RsmHP3yyqYo72K5U0OrqdC4DwwkROYMC2chVN6QCpikXduPRPpWpdZSLnX7S90XB
r5Prw76GAlQ/1RKW7b3nPvZkQsR7tFaApyhswclPnvcuGaUxSWiPUFPasb4pPt5v
PYA1rBl16hADtBKbWgxb2T+aHccFOGihnl9p9v585Wpud5xN/CuywbzGRKJ0OmnO
uaM8bdjrfH0ErQCoZAuE91AsmsusCzix0QLdREU+veUegu3oT3LY4qe/f1pQ8fNp
QEhXoeVbypHipf6rTPfP3e2j4eMSm/yJrPuJqSJ20vjCQpK5veMeZ199xGIJuupu
8yy4jxb6005Saypt0cwXvdDa3X7XuHLVnpnM2VBj2E/XOOHDxa0/n1+EjyWZ82MC
JiANV4LHk5aFM6lmqvuV3063oRXuhGfimPmN6OI3oYmgbX/fNH8+2RMpqOuaUY++
6+l/csW0cxDtPcATBACLBB+YrhwDCILTHpORqqmC0f1PrNciJnI21SpVhGPQEuXD
FywGlrt87H8PFouwEIPwC6WYWx/of7dyhlbUhl6B+L1AlVYS/R+sfI6079n8wtHy
cWxXViMSpxf/4wxvIJkLky2xEO3c2iKPnHlpMCTGbpj5CTMmYz+UPDorw2L1MRUn
3BCIjf3QNDw6TJYJuyXWzaRvMD9AqWmUf/VM1mq7ScQAEQmdjRciCFR8/unUfLy3
QVaBtyNWX6xsOYRTPrelIFgG5NMQuWwna4PGAcQW42HxzM2yW4JVH+20yN2CTqrR
n7+hG8Nes+fbBjWWddwF2E0NSxJ/89UrZS9M5sII1zryBAf8vZ2M7u8mlUgO83N8
KoBs36heEbNRuAX7xUmYKmK2PPWiCiBYmpUKKnkEF95YuJo2p8SiY/eAutNbd4su
/cfElIpYVCNiICi1q33Ryvu3mxOvP2EUDdrCFaIp+KavXrsznkacX2T+DGr5gdrL
nQlWCnQFjwibZflDRB56zc4ICbmi9rusdzE7ok+aG4G7/UPbD42MXSiE3xsW0y+x
eRJHl8TEU/itMFhUvOD3w38RSrLiDg+c9aGY+sKzqyzI06EQ1hk9Nf5VjdR/l3+l
xFc5k6BdM2bljZAUw44+ESaRBZd/Wo+dfsGoaZie19eRww/Q6OKBXS6tKYhEH3HE
fDXQmiZbQmCM6e/+5h98Kz0dmskZ6EAhtHl2Y+72PkAT1GBDidGxxNtVO0cJGrV0
IAofU35Q7XKpyBAf5N7xA/BatBvi7G2OMewUkWV4nw03/AggE2DRZiRiCMNjRu85
Mo5R/wQ8l2YqS0jd+E5s/aKqhdzWMMqNqBfRvnsKEu4peiqQzGch+D1tPt4A5kMH
LgoVKpDmzChpXcvQvFnic3EUMaw4AJVTi9j7uP7mJo+8yoempR+78aWUVB3eJ2DN
TMyUdlKGIBdShrCcn0iVr7uEsS+kjBgDzbHQNT1aWpJwhCf/gFpnKYtTJcBRKbUV
g4O8U6ywe8qz+anG7BD+HZ3AXysxzn6ciP8ZgpjYxJfKAKkgjoBWu72+jm23xUjm
X6/A3FCEcp21p4f5GylwY9+0unsjOn6zxqTb8DAfrsYWPQg8aVzw8/GyJ2omxzGa
G/0RdWynEt1byLq8x0Pf5I4HCvE4CUOHYdj+NRxcH2xss92KtnHEL0Vlt2p24Iaz
DlIZNJ0hl2p+AyAo/8x+5JLN0wW4N7OBess6NQlTL+RRG4v1u2zuDkSjBow+NNgI
`pragma protect end_protected
