// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lBv3GVliY1qjDztpHOrrZiOo75kFOW0UFvoGJvvH+tCNhoFwriPiKDf564M8
iuks3cniWG8keDRcvNokSl8UX8YDI7NnvNsBC09bT88GlSs8cLHvG+LNFVqL
Tj0feMKstognhES6TEZmBurlElEtSpEgcE3sd3V4i+1bLfpcnhRju916Kdyv
IVA2te9Q5YNMyI+tY2IPcP/0cPtrxgSPqESCoZpyUmW5f/3pMDnRag1OCwTn
RPoze9Jzv8otRvrRRXijCrA3x2PPBa1OBaz2xbTmWaiokc2QFBmV2OIKfSM1
kyhaYYUZrB10YViyLTX4yXFMgIT+CLllREPVWA2Lfw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ojd0HVxCjwNnHPUlYz6mDrRJYDr+YksW4s6LcDMFmw+WrDqr+9AnrbmjTgIE
pI/261ZQGB6DlUHYmvYSaIbbSS3xsua3dLo66N/sAtb7ZWrNXyIWsLEWrhen
UMB8c92pfaVL7F1ahm3zmfLr41x4bi+4v08kVmuL+GXgIfnHTRqBdY/ZcBck
4sPiklIhuUaPrfpLrjxzJJbCG5nWhOT1W97FIJRwBUHwlondjbQvRIZvLSFt
lMKu+VDYxDGjUFiaEZ+bvo6AqOuIhofsYOd2iS7AoQGxVLpAaG9lCinZIjVU
ZPZH9HuFpyF+8O/cBx9icmcLodmanFdOzlwBnC60GQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DcOuMxkC3dCHOcWQk4QLcFx4jkqQBIrx+3DsdFScaTVr5yI/aNorctytPjRc
n9Vrp07QSslgror4dUaieyk+HN4mCht+FD3jalxAGvDWUvhYWmHtkHqsxmZ4
Bk5Rh1qKJOY4oIDLYLI2IO2hs+Skv9+ah4CQip8r0LJnv53RASJAmfsVeWOa
3KgSWDz90KTvFDK9CjbNj2xTYUYN9WFkJd0uOhQ4bnfvHHjkWRAPZADCMSld
YBKnza5p3HCFnOueGtNm8SSS+GeGX++xMtEKj11K6wg/GIdFi4KswqFBI6fw
NtpASj5tBS9WpBLqd1dwbTmiuIorouPjw2ZNycCX5Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GhNrlMtrxHizWNMDsD9b7Q12WJlRBRB5hoEwqpwoiFtndgwhDPtaOFjQuom7
VElwL5hwEA2ltpdK0O/wWBXVa4bDXBMW7cif9LFZuu2jxSh6y5q1ZoA4SnNT
q7n6nfiAFWaxoQSTK80FMTHo98nGE6WnB+/1eNeqI9f7iVNaFZY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cB71pJF/KTMk10psmGH811rb1+8O3iShPnOMGjnxXysTTRHxCZxEpiH4bzr9
k+qBkWgTs+rXPMAi+qEqs3j75kjBmSt+RF1MJhKbw9wcZS/MwbtqD42Il9Mr
sN5h99oBptI5RMFXOua7naP/gcwc7LXnr23nVJWmwdLr6YasNTtmxIXOhWIW
WDkHz84DH0S1smQnvWVTEicWxXH2z/CiZb01KOPRsNrTVuYj1NfUC22K+bK0
J5+ADTRaPvMwlnlBwd3jbMXe1m/wmqk8kilBDjMZwLHoc9Juq6OLR1hZfjSU
EBbguj5yGDC+9EFwG5ozNEGL84T9VRftk2fVWOvQDymKgybH0zJNgJ6Bwe/A
oXoyqUkA29k/b8xpH2oqYwWzGAfJZ4ndVzte7vL991VddW0xfB6Jx27g0osO
h4v2oZK+O9r8RQ4zoLcxLyhTtQ1Aj1gKuSg/SnIBwS010XyhQFnaPAk1hDSC
BWU4+fnFBMBgOM82S/BqFqPlMPfrB5MX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Lph1T6n+UlGSq4c+NfE7EbIbX0S/jnweYVqJmE6sq9gIYiXdJX+stebC7NOX
1fP6II0CgZIHP2n6YyYNVIy4l93UY8dDeOTBwTZlpPZtcrk6VmmpYApgIbrZ
ApfTGN3Z5cTZSURbQqstXnfDXaZvZglwSX527ut9ZFxK+8zJIf0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QQbCpzqNZQqhc2YbSzVnMYUWyDr0fSOdpd1zTulTHFOb1hlVUdcxvxZ6XBrU
TJAmbtmURsXcsAT7WkB3l/gTmuR+pWnUU/qchkaQn3VHnAJZDq3CDSxBHL/O
YKlIZTGkTxxpMgM9CsABkMIn3dXkG2sf72PWKbSGEn+1I7fP+Po=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 30032)
`pragma protect data_block
Z32aTPQ7wjBfbs+NzgRVa2NXAXlHOCV6YXMc1tYv2H3SNyxatoP6t29jqziR
yZCFfwpc0Til7QROwjxxql2JCA6oATuBbgKZqo5Hi2pIbssgBPnCm3+ncVCF
Ww9SY2GqRQX5sy6+OZ/vWXzUdx21tjqrX04okxsDVKOfPgffiRu9hjd+eaDj
SnIV3m6nv9eCk+dXoRTdtDakNJkOnOwjjp5ohdIIsfia+MGqKZjJ35460yGJ
OrNWUvPVTt1X3trg11j5MwtcjoJZgWE88lIpV75OrTXSeS2gdEQuA6m69/5I
BGtq3Upcdj7btXOGiQTNivca7sHb67IWraYnVeCzaADTAeydXU7WU0Ca2gbf
S33Yd9e0MWVOBYASPkVsW+A/oGiY3d4FSqkKE0cnG8UwR9tJ4BhgoskLVnb0
MHj2h6M5Qokvuw2Clu9rhRQHmxglAyIx1IfVTQbSoasf5MvQVKq0yWInW99n
4721eL64ALXIrmg60OJb+dsO1JBl2osdvuBci5NueTjaxUG9WZCLDTI92Ql9
3vVtIFs6fpVex00cMFgtvNYRb8RmujDOZD+cXoLVQr8BEz6yxSrUIfr8r2EX
24EHiGlBCMEFxPukOxt0HqIPdQTCJ6JgGEYPKNTHrWZrvQj+QuiryVwIHhzO
jypET9dy7hXSpLkBRRJbZdqYzrIeNbz3K5/rAbUFom3G9+6IopNLScJNPX8P
a+DJyaGA6xvSGsC7m7UVD7mbsB0X7vBr6pGw65ilyk7tFmJ2j7FTtgIfrdw1
grm8AK+P4mugY8fmbkQiZRRM5iuqBOrwAAZyOHn4x0cOnm8IHBsSzDPJUqpk
eGFzn9Umvar/Bir6CG8zE+vTnCFMPnUkPGtGi8vEJl1O6g4n42EoGN+Hv9m+
fp+l1f4FhOjY6HUpSxchTHhY8R7PkVAvxkWmIK0c3OnEfh2qr42KNpCUXRoV
GunjHBYwSqv02Ntoj67KcZeu2r5ne1PcKzcxBVI2DYB0y+blrvzzSGuFk8bG
+GgZ4gva7Zxba3Qnq3dGEEcpTHwX+tyeSC0SZRngEYuHLmEb1nI9YZqyzzGO
W4CElgtp9x6zQtbPDAxyS11lqtXQ+8jv1JDOhY4cSummyrCpq4O9oynaUNfN
YwKwUuvu2ZWiycl32cI/RTPA3+Jxx49ZMtzRjw9W/IW+i5J1yYfmWuM7KYLQ
zQIy8Q2+x6/OC4CYpi/dhnpkP2eUcXujcK1wSk/OBAOuNsMjsB+bkeay47gh
aZtRhSfROHwLRdZa6brjLOajwtMhDrRkK9IOK8dmZC6W/kdjDpv6c23/yIyT
DvA0vRjONBAYC2zoEsR04JEdBCDEmgjpqdOzuhP6/6h040bCruIRi0C1WqKN
cWE4tpXxZvfU34G5i77G2TQuTmwZ2ZiOXdoJ31phK7+olC0o6lZj8TooNgYz
8pKHtsE81Un0HJTBNbdeAI1uhKOXFd0zAaQPDtmyjHBrfYx0BY0rRhfFsAhI
Yeigid7guZe47Vfq41iT+7s5ozilo8AMlgpMNK3CUUtExN4FO/+egrzxd8M5
bUlozoK8JxLIV+B9RM/MkPOEuyPF0K3Hlaz5uVFtOrXqBcTOxOAuuLLOy7Km
xEyvQly/kZFyw4wcalnPoRfUXD/EaBdEA3Bix8ZUSzKCnSEmm3XsviXpsX66
njzMwaD9QEkcsrrNM3v5gb5Fq8BpLdR0eGtN1VJfFPj0gVx7i+pSwz3BAOM0
LOO+UNkfsOj1D4IZyJvlB6D5r1aLQ7lc4wqrae80cEKeCFQgbLbELrXolVVx
ENEQZmIf5Ry5JLEe/vMgGfqKFRUc6z2L40737TJEcGa25tCh5v734X3pO8w5
wAG9kR/vao2/OM4D/I25BXBlQJxYsrQHTYSUHNK5H0WOf19d/6C20COlytDt
ATgpwxlfF/qHmvdLdUhCDE3UVd9Bgj1O32u6T9DPOLzA74I1bxkK1pK6v72F
7+qjwkrkNL8/kMXngE2EWvj+mAFaVUp1dHWUqLXJgl/pyE55PVD+5hGFzXTA
FaJ0bw7opgU4LKdwRsnc1f5Yoio1/ERIJ2Ns0iWafYNaNHqRN4JKL6q5FwoZ
ACcYkjCk8/w46EKT0U0cvb2h3thTRS44yj3mqZxIGuSHop4Q5njIvQhYVY4r
Y3u2ltdb/aCHwocSj0n3pOfgMFe2olXEsOEWdmMP+N+EjIVS9VfPeIjXUcaJ
yUv/MWdHBqrjZjWZk+KEGK419iKnV5gY8HrB36K2SxmmyYcIDJmPId2PGm2Z
LnU9G9QKzeTnhQTg1YziRVblcoIaBeTRPC4AW9U/yBTduf837synHFcc3jZ0
XkGYtqSWeAvISdeJD0CYFEh0pCzGulbr7Hsvd31jJU6wAmcrI7wS0SWqvf87
LnKQ5wstb+sVbur8PQuymGeBRbtbUDDMgY+uIS8dQXK8ILLGMZHRrfTbxKQM
7XPOM8ArC3n4MQ8UDBFy46J111Wub9Q823zI16/QKn8OqBcqb4tF/LsRKCy9
3FcLJZ39zGZAF7sPySMH+aXbCIWmFsdd6L+LUwjyJszEgEmArRCHzFHk8Bcj
lJ4ODf9M65yj4S/+oMcWSRy4Z5XXIlN1zDIUPkzgDceS+eZX/LDxXuu+OvlK
z9E1NeMPJDEdX/p681I8fUwfk5T9pedUHrKisbq7MGyJ/oCMDNlPm6sGcql2
PR1CKMS5AttDyHgFuk87Aco59lOXq8mJIFhU6rv/hvczRuMhgcsSjetG0HQg
FeJRRpuXWURGsgYYsGGOOD1eU81oTNxCgkWZhurhNzETo4yPzuO6D+fRlwqk
iSBhypN9lHDa+XP3Z7fZ+4quynfbtoApYb45xWjQ45O5ZHWP3CbemUwFOTYX
cH8uLwofsfclDqpJ3Ue1Eyk6psmPUH1YK+TtryHwY4hKWe6UT2CiDm2xh/gg
N2cDYkLvmwN66qkut75gWPVnwTLgQ0Cres7KEyuPied/vj8+lhLJzDljYZ8G
vhHBCUHwzByv4E6WIS/xPaNp6DLJl/ACMJcPCym41ZCx0R+tcDNhuPNHxzk5
MNNzQ1t3ozdUC/DjwxBwygguE/uqLs0AZXaXUN1avAtMOgxlrs5IPAVDzPCb
x/RZvnvlP/Ook14UcKAXsmWTjWafq8dM+y0daWmbtbIoV6xPglTizkbfq5Wu
NS5moPShbU+vCdqjWIWg7L9FVEEDHMMnxAOnHkvmWqRC61WQrk0TayGD2aYx
1IHRlZ3oUZ89xOz/twxv3MNvi5DKrY3pSEPIUVYI9OA3OvcAh56l28IeLAW6
AmrPBHkB/ghSC6dWJLasFWkkbJrVbQ6tHWct/OpbispnNpbeV7M71d2GKHL6
BMli/S716w/inSoO9OodxaIJKvxxLL15UK38LNQ/LQVnDc+PFN39xud0kEpG
ge33WRneY1KrXuXGSIQZ1qxRqtCbzZ5YOT+Mz6Ai0mSopvB+8hJjV0C04JAY
yN9R5GpDNsfpqGcI28GOJUiwDk+t0KRzcrOY5+sF5c0nBvxWhSjNd3olbG4U
P+eLUi7+NQezZVt1L93yn8MPhX6tTbqtpgtQBQI0SgcLg8rDfbZM/wGbb1zv
QInaqzh/guPSW7FiAHdIFtNI6FBYWjfNbeCSWgDAiJldYaml/UZTxh7sX5KO
Hf7QPw4omPZu+hB0UVr/3P7O1d3nHsPIm2NFJVwffHwVD36y0KV277/QD+qS
QnY1EDAriXX2EhlVsX+lsG2fiVPsZ5Cu7f3r1XtJCp5Xl5lN8sLam4HCaDuu
SO/FjPJF5kjabSgeN6c19qnOhqUebSUT+mG4tA5TfV7R8e3tqAvfq41W4ldW
t6Han/pxXJ4OL8NGFvBqMltiai7sdsLr7g6r96dIJ5iJ4TMcmsCjbet0tvB0
pWWDN9vnfQqmNUteG8I1ufOMHupiX99RIYcv4It3lcAPit/vY56lTUehpnCy
iZEa9zZVQxZm4a8Cd4+JkGCHeBKOAjGeNU7RgFw3J3t6IpBdVvLFScqknOmF
Q5muAbV8fNI+u5K0+rQnnU2+fkN84QlQzAM3aebv36NTzmrqihquzsouDf8F
S9lfsSHkRLD6XRIFooHTVNwbfrX2rv8MIn3JPRDzUOh0D9itka4DDJ9xaPYr
hQi4QoSqDOKNt2LoVU/YLJuwpEdgUq/CaMElbF9dHtFsNh4n3ssn+LSy/5in
OaDtsTP/1fWeG+BjMQt/nXjqhMKh1o2r81xFdEcey1udP3Od38eHtXqSwsO3
+9jhbxn6+8+UqIrJSJjoIatnSfSYQp2MS06pQRsuek3JCNwlyJUBTe1xeGC6
zYRwO+UhdboEhWAbM0Y17MttSa9U7IWx8yku6Ayx4WSuS+kEcJijkt+DJ2cx
qocEK6ONchp3skhkCIeCACn8qlnbj7A6bRv/W4QpEgD7LF7a2vK8u2crVgmj
LYm4h+lT5AL9lIHi16hID3kALSPmUrW2pp84PYMs6udEgejFGKmeJvXevNlb
5umVjdguzWdR63GoFG2BNzWAk/j8ZiP98J4WuJSw/S0iFvD42elx7IRGIFsE
mdrz1KRBPV0/vL2r54ek0sE+Mfy24HvCoUSIeMaU7dquIdegaiMy0OKjgktm
8uUnNbGSEzLDB4nKNRbg67cnAPciGAPKzj1UC300beCsb4sCjmWDCOWOqnaG
o1Qg0mVpPr6U9K3Ie8HfLqQDvswU+9Dlm8O7l0Bvs0CguebAvSX3kyn+2At8
NIkjG2fMbaDE6rGo9zfLw47ZFkxquvHfK5jg6eBUXPiIhUhWWqPle38Z9K/0
xTNIaEFMTb6lKgfhjaF9M8I1jFwjGNRSskBa3mV9vJsxPDPvRaib1KQC4ByE
MG7V5VWXBcvFdOED1Mj60iNj2snv3rgYsGcUAdtWXVrdtr5KydQ2PDt0t2dh
HyPr0m7tKfRsZwsFgjGu0O7o1DjZgvXI0K28UzVHQr88p3O+wBoNX+T5m2Iu
/kzxrjRG4BzGa6iI64+0SHKXcREqWAEbWcntckagIptZC+jd4QDUcfq/kVZr
O6QTwOZ95qo3eH2akByEVcZS0ctpb1P2NOIQC+csleffn5t1lTpqNPSZcz7z
BIiq3LPSRrh5l9migJ6g32ld2Y2bQrtbnLNdqs0DP+6P68ena9KiWTxZDKPX
u+zlP/dbzBER5V7lx7nQDJ9Ma20g4bHaLk3bu9ARmU1VIRvNvEyFEszLSAHK
VWrugr5QojEYXpvcXeHnyAdbdPhy4dPMEQ2wpkRPikrSpcCY0XvlaczrXX8N
3hUgFaLD+Btg9UuaKq8VuTw7GCgev9ILrNRiBp6e3KH4iozGkHGg2i1l9BDE
MIYwhvgurl8+A1B/0hU434vD7CMcPoMnIdvOA0idHjEv6TGU2lxuK/W/iWZz
3hkSLNyeT+a4HyyhdQAlrW41JEJW1v8MEllbCJlZMoNgyX0uwdLShVRSetk6
RhtxCEYFeSuV06j0CIbRYfOAiwKqoQaKv7r4VfcRLx19Njq/anM9nWl085vK
aN59EQSDzwp7TaN5qOo7RMFtsKSRwBsOD1qGyGMfASJGoqUKJIP2PLsipWVc
zCfYLSktjlHxZ/8E0H1oH8keU0mDlOOFNl6lp02AxC9kKAko008hkazog2Lf
nijoVgXS4MOoCJ0NooiH7yIItHTb4Gq3GkTqnMuyFT60EVZcguiRBHJvQWep
bN+zCchxUwa/Cri5p4otmqSQ6uk8VGZwzPRkRyQ92dKROjfAiaxeLTCLC9o7
V+5xmqIP6aAltXDgPOYAhIK+1mT9eC50QYyZ6lh9l9bej2N7HA/OsYqv7VPy
9aPavDmcsSlKf/YVtSgKnPDzruBhf+x6mn8AU77sOnjlf9JKpblPa/M0I85I
ZMiPHtOnrsz682IYnHuCR5jIcG/7STraZVWY9Dt2/tTwHPJ8kGqQNg2Pb1Zj
vCgyBW+1nfnauOox8bxg8nXkKv9cuYndnqGwA14dOPblPKRHuT0FdHd+vwZK
+66G8pLuUgPRvEg5rg3AmB7+98RqU+qm/KSs5Pbtswrmi1lrOIPlUzsZ9KPw
Jw8mi4B4ucb4IdVZ8RFGw68UWvZPCF/rLtUvHMevU6pon1XoEHWC6qmBlg1Y
UOhn4djnzw4JlL6VJUo/7KDxwOLcj421N2Yoxhd4gLEtEysQ7Pmthef5wxhH
LMsGmdU+0LqPYAHESW898mqxNElq26TlV4C9ujXdH/19lShm4VHx70VWzSNr
ZKSd3PcWH7JGmY/0mA1iPRHp4X1U5KKWq6kqbBZ94kzllGaG/W2uV3+uExGA
DNvfk2luRJuZCnM9V49doP8k34owDoy+1X1KvTVootitr30OLMyBjRDoLktq
umcyd9ci6U03SszlCyJ1wNaNgi3VV4CKXuCctVqDZPD9DWbPR0LH57Lw52AH
wCSD0EocP5ugo72pveePwfT5sdYiNYjWB/kkVcxzzov07YU7y0DK14P8NZ53
th5coi2LQAPWDJLiUqP6Hr3z+Buz0Bwbn2sHDI58vwNN1WLJtWiRu6nmdFv9
ddZ3ZYby5X1w5NyUstaeruAIedUIy93gP1LNy8sposvguki40+lmrW9iwOll
FjOLiImbE2qtjv/me8Sbitc0T7hrmw2mDfuPXbbptG0+L+19qNGM5q4+hokf
juCHZ6M27fTZXmqXs8YDWZKTCtJC5gQo8CfcO8aa5RQRkusI/JrkkU1MLzHG
PIZH3zjH5FkWiptVBp9Ws9o0+u89/Nf8+evxJYCcu3wduq77e/+5wcXRwMGD
uL04UEy/UzqpVRe/N+c66VerM2kQwui3WfSvQ8UbL7ZZWJd+wISvsqMqZPcF
rLSgySnpHKAv9OmDbSVcXCBgrLcW5Y6eSRVGKoaLc+FpvN5DRqe1lHZFvBfV
3TqFdR20+K4WtebodPOMOT9qD408ZXO5VyiDG+uGIr81Lqw1ZqZumk8k8qID
/ltQMNn6PF4bZghMZhcOT9Jw6vAnO0xbZqdHrb/xLQbK/J8j/aeG1dui17Hw
HKWkxOpmfKYwrLZw3kU99GZBU2dm2IuwK8/1zHENolaUaq4Z2c1sOELoiuOj
ZaEM0kKMJ47/gDFvLVukXgfT9dJ4YV+K2jjGhVWVOOEN2DW2NVlZ9rB2kc0h
0lfnClxPLaULvXzns3c1Vlxc7UiI1qK7yLjgW6GGgzicWnIpJuQXKtEyifYW
l6Xc5DivKNdqZtn75LUvePCxmefclPWspm0odIkCHPvfWNCuADq1/oEg6F1m
qum4meZBDSa8vjDcwt94DPLiE5atUkGnGCq77YoDKFE9DfncHlgo/bRVm9sE
zIeaLEA2ovlhUMZ360ZsF8yZUAf9im8hSV94hF8M/wWiGjZhuNuyWHuMFhBm
eHnxBxDCkUHMJSA4pnN5DLRC1WmJTEaOjgDKM1ka/u0g+wH3DtsMtvL30oqM
KzvKOtaf6i3ivX62X6txSuzdX4l+xkciiaB0zFl8cP/Xhz9eLmbmLeh+mHUb
Ydq8m/TPlDz6YvpVNA8D991N8n8daDQeW0dR0lgb5LPTqJggNIde3dkoWNUL
4JB7Cqj3KgajjKPg1z1WtIlNlpRWPgYXBwWmJjkUAHzUglhWpA3Iz20f4WyD
YSDZUJ76qCdqYSNltFHEl5VllRYu12hi6AV14SIqJObTzcqihnSq3WUm8CU5
cVwgmN69/5c1WJDBGnn7oYFzMzLUO45kxCS08LFY3wuaXjLya8kcGKXCabIt
gp6v5XIObQgZfvvzsheP6ClR7brQo6b5IDnYBitInoa1qaD8mZfDOn/08xbO
EbpUInMRQ35AMNuTwf+/yWlwMQqrGCGfylxKwHLtsamSUvT3XkEyTHDsMHNq
7JxScw6cOYQsuWj76pLD9c9AgC/OZfUd3b4amypC8qBS9v6E1hn/omf24fYT
VnZ93hCbZOpEViuMfhRUSADKPauJeDzlctiWGnr3MpxvHJAR45Qcpltq8uYj
0RDM6LF0qrUGzs/YHqqurnUKIDloaZUOlUgpRLBmtKjeanNvi1xNGHCyTegb
job6L45lcv/v/98U/qoohKNQKK8MLxhj6XqYowjA3hf8KaE8ccdesnTVVIx+
EQl3sfkYy03nGLqqON4L/ciPFQW1WHlpXi7E5WyPQmxXm8rppyJ0JAqmJ7ti
myYOIDKn7vIvllgqjxefulDYsmO7q6Z+kexxBZfVJnKdRUZ2BK3SR8QacdyE
aEFWA6jou82h+GT/s9AUka4DOdOneoi3avD29+QAZOYZEaKJjm+2Re10aD3c
RDfDEftOmbR0P/gTRNtQvIN+wa1sxnes0/E7n7MEZiyftGaHXb2BE9s2mobQ
Btkg1rIR04QeWOmxblR5jwzPk7ft758enVrpPFUwyOEouF6rOM2t4TKqbOCN
pEjzMVQ89VswkwpamfB/T0lp5QG+Cg3TGllX4e60aH1maTZ3fvo0ny2gfMa3
6aUKLTCC5rTeNdE/IVLsVa1vyZHzVbS6i+AMlvyfTC61OPzWDiRvlItZT4f3
EJ7zlySbwllI3IP6r+6pj/2St+q6Xp5FiPq+AEgD1M75X4NqQdKrHOoAQ06Q
4GjyaIG31v30p4vOD1FKlEiO5Wf+I8HyCMBYfaxdioRcQUY+2pRQdmxmQl48
thcaHoQZfu6h7FJ4Y4Z9wlCFp2NXnxVxgWhiReZ50dOCCab92V6AjimR9Mrn
ES6gxrRM/CwKbD8+kttXvkB1caND5MzE5M7SyB96bi8J3rVqOMiYaj6IZwn5
lc23bAv6vP4ouGk2UMQdaBzpmzQ3iq6EtDXXiPLoE8ZZEbMlbn1b7dgjjo1R
2FxMra5UX0jQE6GbqRhk6Yui3aJKNJMvIpxqo1uH1z+6ep907/LgpGuPOKbL
WKWCapVSjZKuT0uDZdz35EHcOjlgapMdrqt6QGQcY+0AyMP7seRtWktgrcgL
AmnMtTcrEotcET1gsAez/Qkk7p2F9w/w1+4ApM/BZGrfnMYfnufAtdI6f4D0
3UwxsE6TXVds6AES/zshX6HQWDrTQVw938l7gNpEH+3vPtct2wvMA988UpSv
nEB6NKJMFoSsNqelRm1DEHvQYvpjJ6/UlbJjBgTwsbT2Ty9kmQwGT5zP/fQr
7JD3veN+IdeAKVcNUN9gjQM2Da7RDYPmjVKyLyQRC3vf9KNvMfCX1U2aceWX
cul0j/UzpMosuCZsTAiugzSMYQbRshbq0Mn999RdjtbPXxWwgn38r8p1e6HW
ODwx918U1FUxxzOxPkgDtvSLDuxN0M1Jk4mxj0NhzCqFMvkPHtRhH0GtbpCu
gyBm+l6D3qPWI9peBmQUU8hK5qv6R2LK+gBpa/AqgDFtUO3OhDhmk8nMSyLB
sdKzcSACuXro7xcBHEQUsJbXk0YKUUmNAh4RaAeBFpQhNnNna1oGeBAYlR65
iyyveRiTya/4AEp6oCzPIyiwLO9lfi1QUpYwAwgvBhcqKwYanCSuT4LX9HVv
50IplGV1nGNWjeLiWFOQU+udH/j65+VVAaCwwz0bNA3JGH+cYNc6F+KYVGvK
VhX0FgK05FxwXskir1XNhl4cvsKKTBPyL31pWR6MZ3SDhygfsrSSA9QMsp6H
c/d6RB8N7qEPzAPSxVzzDFtkNRC9D3NP5gsFdiLaSMNh3pal1DS2GrjH8RXt
S2Sjh0dH00hbBOHisZi5c7lpFqqcJkLXQCZloJuwob/ksswKoBV/xGvxGlu2
JG03PlHKok4mcEQR/relFpjysSBLoZleKcG6Vug93KxIvVZXgLGJMQe/fiqU
yYyabvfuuk+mGjWjdFpIKA7NtWENcghdE0kwJO4Y89de95KIdd99xYGFG4Hf
LEYvgA1q8SDnDp1pWw3igQWkD9qBL0AuuVDePp1+IqIJw+U4qKo5/VC31p7y
sqUWlJT4OkoJeXOST0YtaIDRO+GVdAslYA8nzIFC3yJbPVyfC0E/EqKkHGu0
CCo5QAFbqz+/Uee8hcjatDa1JNYGlGgBch4FshYXxLGTa8P0BRooOY7ElA/X
6Ab+t9YYczNfLd17QjSiRQkurCzN4qn3+oI+J2OdY4fMO1KbkFpaoWXhts38
tcY0lIIbPm7NSITYTgeVh+T3m+DHqskXrDOMaroXuH3uN2otdyzbfo84nzaM
m1g+BQKjpDNY/iyzA+7nUesVoLHyrvm0HhJw64qq2o19NCT/6BWgnr0v4lzd
L1e3gWUkp2DqGQtE0Da8qlcOTN3yUItrr6X+Ac+Wjc8vFkB+kZaeJ0I7+ITO
NRgLD+HuzYawhYKEGaKpjYEBzNt7zPkxvCLolQUmfbm26UI5aukxK9ayuoF3
XOjRyUYzSg6A+SjDgX4Cxkv47cpKpU7L9FzXcSyuoJmbvn0PHMhDZ1RPX/8e
75VAwg/B27Np5hpXBbgkugKD8ZoeFcaKguZWwSNHsKAaVwkulBE14VvV94PV
x2DGqKDDG9LNdOOo2AYJf9axewS3Gcklcy3G+sT79BKmtcBDn/Jru5dt5vmB
lX13i7NOH2LapVw9E3I+UEp/HJacWLOe0ClQrbgk6TdW8/DnvTZvTx/oxSIk
Sjd/dM5WtMHKq+PUGkA6M7poHgXiJ8RjZXJ19wwVBwPXi+mtnHr5PZScC5fm
6rPUmMtPwn/RdRyJaEEX3CBXiptaalvaWDYO3sPy/06VmekYi8HWcSLxGcyd
Cc85WvChoGDXT3txPp7Hxz3TfZv37koShkCig8pR07k7/3xuUcUCAf/W6dyj
9pIzj+qO+cphBzGFTMjogocyq5e0+XkltH/tlLn92tXSoERUfPsa1rMyKZuy
5WUCtIs5xmOlNRk8tQuk1DLZQUgSEPGzhBbQHh512rtdbu1bhDRsehBLmbcQ
rqD3VklOHzNMX53yFUfS9ez+m908kx/x91tdqKXPc7iU6gymld3kD6X2fcur
brq73WchqMgaPtskGhnVIBDMg5q35c3gU2/NBUmj4oSQpapOoVqBzTf3s3MF
YXuPXf+QXRgQ+BpMvGvm3gCTwjc6YECbuzEmRRpqtb78GpDMnenwxiDLooCC
ai4VWeNjHFd9bTszx/3vzMvErnkdt22lL1nMZw+A5TOZLoC8ku0LCoSy7mvm
IDXu1cSzRyDfxZ9b9ZZpa9PoZn/HZ9wi5LN/0pJQshcVFsjVFQogIsfxiR/1
iEHVUfr5AxMBRgd/jiDXYMYXbt5iOmXva0eAFtLyWCCn+xEkMldGVMjCgcTN
uijBplAY9+RV3hOfymdTjsOU3E0Bv9v4rOmndakyFqSFnNNx5ZTNCs6QdubU
4vPfjS4PCuS7daMKENMK0ha0Id92FmUWOI4YQ9gdCfgExKlBx9U9ecsd6bsR
Lf9VhDD5GFRLUpP4f2eDp253nJhZiuq2wCerM/Ik21G4ycUisT2/i/okY25+
+QJNobVLCjtXvLoc9kPufgOXJxgeApHoDZOnm6s/1M847X/RYcLak2SLrep8
Si74KJ3Jza0JChbmk56TYPGrL6z94Pt2hIPNuudgNjZkVH4LDzRyY/v7vxqW
9iLU2S2BhUYntlGDrwAiMxAUPJ7En/hwIqsQb8zOVtOWP6cDgO5IFvipGtRw
yfQtnNtnA2a5c3RRzR+vrdjvv5ebZQomv2ap3HNCpT+39Y8mTu2OJ/I4MWZ9
PqNpd0le9ZGBOYEc0iEB58IovbF0OHxPIXZNXV4QhrMpBvfkDOXL3NBQzcOb
6bvHQdBtz7CdTr/fwPJnN/hVaHvaabaWPISOggJR/i0fq9QV6boSz/L7gOiY
LQLX6+k726rxAtUaxOmO0GMVk3ZQaZoGBzZl8hztMPcKdAfX1OGaxyyHimSA
5pGRoeh7MrRMy5TLrXDEAmKi7STwDoM5a0YhPGJGhccSDWZi1EaAXc7tYwxZ
uW1639kOaOLZQcphBt7z9Cvye+9exWrAYx6z7zdeJXJnfrtmRQ1aDuSx4n4E
RJ59YObhaRaoCCP8NmIPJzdJyW4XH2fKIzWenUsH0e1SUxqN3wtAiTr4S55U
sjfBUopSzSBrL/CxaxXaKt/s3Zv5AESIejc14UGjyUGm61DcpJdg2wFpP5OI
Yc5tO3NozyP2fyS09btWohdfCtLt2r8Ync+PiNhk713GkoaiuCPetS79bZqu
UZrnZEB18okX87z3gVYYqAZIbv4hqNqWUp11ST2lbk4aG6+VC9Eq0ho0l8Ma
2KzlEz51Vrpe0S8UsdzHQ2nON2G+FuvKTNPsj3v1FNUCIyExGMjA4vgbYueW
G2z+TBlhuoN01OMO5f99xaP+Ex2CIQiS4Bv4/s3ZMqWSnfPdsulBL604G99s
w9/PgcfO2u5SgP1j76w4bBXJPHgCm1mYlrGEfI24arQ/io/l0APJFKquonEL
Cx0/at75W+yugOrkDNcWAA7JcG8na4pnMLqvOlhL/EoN50FejQ1NJO/wuH2i
U8zmbEPxBCQCBrli9nnaa/WyqTMth9PIZ4wWjRZNxP//FuI1yOtB/3sV6/tq
rY7ILNL0Y0Gi/DK/o2Aj+j3KM3oDkJ4SO+ksPeELX/5w96rbinOoEUIvlkVA
W6HLk0S96jsvE/QD7RzRf7XLz1I+HuLZhgzctBwYyupZY+nwX2++riWFFAk+
g2EjA6jHhIUURO9GAzeMwhrPvB49S3CF6TpYBjTdBr1cMkyUbapIB1qFoX8L
rJ7L7Qrd4yqZH4TO/nUDPvNNf6qmA20N1rxFd2IyZqylOc7IHBuWYxwmACqC
GuSLeyAD8gfjOwJwjIEOPuM+8cLh3MkSrhazzo+lHo0a76UhvTwo1iPBIQz7
7VAMo3sfvmw6bPxR1tDcRijFgJD4pzat9MkpwwO/HoF10GSZc61ZdCp2ROXL
MB9t8JtABSMCE7qjMUM2xfhzzqBrZeeZJGJVKXyxWS2BnxNWhkElyWgSOSRT
KMdis3t5T7kjApLIhqlGznpwQlJRcptIry8/UNEP9lrBz3dVbWK1EEJfOixn
M8RFQUJq6rn1bdS5Jhpu92J2iT0bhhaElJKySUoaEhEmSaj8gJ/joYBxq9W7
5FoNrxVzyDJH96Q+nczkSnGA3HN97NbXQ/QdBWKKm2OAjSLhLVTmB4b/G5IR
h1YViOA1mniI7pimEWhhZT2c1Gc7OsH4TV02wlK8qNvxoZaZh3GMBtqWIrsE
AO2z4kbIqik8ymzG9/CvWUDNP/ubqDkHRMj/SQydNDIq99tmCrmFtoMZ37IL
ojWjEy92KdTmK+BgNwt4nYKYqJQ90c1k9jU53WNjU5jb4Y7inDOKICE5DYfa
iyTF/bFw2eHgtHajncedRKkqGGvDp7OPRYBlqt6zHG7GL59ae6YG3TTNdcbA
Mne40pqb60tINQKp5TIJf9nbTs+7Mk/EE05Unsug6HrusmCpD16LgK8mTTRC
HLZaJgYu+0z6NvlhYKroaolvGAv0OIhuFi8xYjoefkeFTTTOvUctlPrxmcKQ
TUguKyI2p282JC0Z5vZFykx1XH6YhSKu9BIKsRziE1tXbR0qtFCSml4PFmdM
2KwzMyZA9lFuBHsKJa3F+Xt8jTwOYrhC4ebsLJ/i6g4AjR1cuVyOrczgn/qc
XbroQ6RVJ+66peLQp/n/cDMSPgoI5on0qiq0Gy9VNJbyV6V2TQX8SQKM9zWP
dKLlVzxdo//aFXlWOayeQyGEf2Gxd2wNsBo7GAAWsx23/Br0S0rFvTdwdr4b
2rUPSBXDNTDOpw+TO4QVQErYYF8sKPDcCQEgM1/CpqTFLcxXw4iE9uCSFrR1
RvFz/sziOUXnOEuFlAHGU6bgLshy6YwnC1MtcUlASUVLv2M21W0KlyiMmuA+
BMKgjYn1bIOmysKtKndXu8yfbUlZFE5DsugtK2NDpi/VgSZ8CzrBEjZU7nF5
FmQ7BqmNhRWE/pwKop284HOE/+bnBKMwIS7lQTD5fF6X6WjHA55LbG4G8lwB
4+cytX034lHQTwZCQ3MAV5X2GTxXzr/ZFQi/laQqa5kTmPTweetfx9JSYG5v
NoMM8kiCgwQAVPaIF2VfvynM6H8zYJQiig9jn8W+Re3x+2pNOSc3S5RRS7YH
KJ2wIMULKbyuR1RIrShD8wHIdID42LUwGH/6N1XmfjVTnOkXWlnQ1Gh+kTs5
lp3unfx6pBTEf44ljvOPuz1bjYvi5dCTN3dAGbP1xVEIDCLfIuKxib+6mbZX
tiKVFOEIIemjAv8TNfUZ2GQ6PSy5KqVLNMK+lPIF5zIXRwB+B1AH+HkiGthL
eux0r1H+XjWUMBxmcMN9kwKK0gIAcArspuhvdy1RcrtDd6bgO2yG3uyc4b7H
ado1DduNtzujztD24gRiUDxQvTiqd78/Xu40jvm/B9BBJYThhuyhdq4hL1Hw
6X15AN8fUEHZu3JTysnpvrqekKEFJsZABgGgeOwuXd9CQKAdaphx75WDlZsP
x1xQBt9MGzOypCosX6sM1SE0JagzdPPi+AOuOjIGCRO9mv2Wd2LwRPz7NEvt
Y+8hosSuIkBT9halw+R3ZaAySedjizpTNYmAAe8+c8fwDYaaNhRdk3ZDsnma
Mf7G0tCpyloeVH0+afmKhp/eRkn/kLVwSh1cZ5SuIAgzvxqOadXExN+XbZom
4vxS8czaCAS/xceCiVHGDYouWFJ8jcecaKiTemMH2GMdZ4c+9FTpRIi/qqw+
X2eSbvhblpUzUtBGJ/wV91PdXX4A0pKh8E8t6r7Dx+HqzC6l6fAmxZiyM9r/
bnXiIpoMv8tzgdiskXHd4bFT4QJ9ZwOIpAIVCrHRvCaChlCrUq9jIx+twrCw
pbZVyz/sNiM/wDvR2or26gk5gpXDZoMdSbfRWVVRGmBOKSbGI36EpVE4Qvs2
tpSHISUTv1kkcS/LTPbcxpFZt6WOynczFuE0k35RFos6OEU9CKlel5RNh/sA
buINAX4e33asBjZdU8zytFMr/WT0Gtx8kIP0hpHwqzru54eq3g5XKX/cI0T7
jiwd3yyjUCKTwgOdLcjvBw3Jw0QdOct7AGSKtkJ0TO5/HOXAKco4s/cMU0Ws
kEri3r7Ovh/XkkxHlkM274x+ivrydizcVs2LQCpdKMkK2P2ozWLvDVmozy6a
bPMJqoZ7LDVAOdLak5UKGD9LtRkBjADQOsdiffcBLDRYsqGYR0Szat/vetaf
PyjN5upSunXqxynXWGwsi+6IwzLIoJM1I/WFzhRgyMUjXKhfVKHEIn+4+cdc
iibZSFarvECq+OFz/SN3/62wq7cq9fXXI9F2Jjw5RGLynIHsPdfuiih+ydoA
U3LuVsmDHKjB6kWEsXBGwLdN0R1NC9G8Pgf3RtP2RTowE5Sy1OkketLXTKWx
xe8PyuL4NfA+XNY4mAQLbkk5zpFDo/PBn6Sare75nkF9H0jolrWgC46Y/WCS
12nyEIwQceazcZ0k2Euwra+G4pn/ccb0TJ5tadgGFDU54Z2UOYVyboV2e2Ra
DQZ4UcEiBSn7nSDnPkH9LtrmGa4d+vfkWiuHEPYL37WWEyKSdzJyO5QGFYmn
qXZnazuGtvqnSXLoXJrUer6eoGL3crFENn2xLFidd8L/YydsdBgkE/jGOa9j
D/FsDLBL6irLEN3aE/nYfGg4UxrvGrtBYnzS2BLvD1Y9V/rlhbzHLkFWMbiB
PyVtdLO3OIWDT3c3se9McKzPNwGSr89MJwbKsuw28UJWdtZJdEDBo5Hrn+Di
sV00unKN+sNBKPCG/2GIPnCfDHEsQ6ZShJ073AR6qEQpUDaqE6u03POUjwMy
pC3G6e6FaPX6bugsWII7eEToC/M3J0I6j7csVVIxBK3LTgnvDs+4AJnkWmgO
L6On6rlAxVIjyRdapHKbM3MO08dJTEyWGAnVvvnJwZvlRQTXYqlYIC/pBo3N
xaowbHktosO4pNb3R3wgB3m+DpxEyoQ83OckTZ0rCsMPAY7VFKC583zIZPvh
z19z5gI4B1J/4/Z1SEuqfL863s1kd2KpdnkTEQUdjIBEFntOTZVkYe6yunrN
8dzFb8z2ISeawQ4rr5+pNTfpXSyT2V+0u0epQqueCVjIArvt4xdhpT9GaND1
IWjCUGuHoAP33zosA+4z29oR8ztOizVxhdzOuojE1chVJ17bGlaBAv5ym87B
UTLw4KbbMc6lHUNBP1o1JdYM0lFiEK2pKsk+Co/OKzdm0ex2X8PsAP0wh+oI
v1kMr7r43f9PcYnqkDzN9hp6AFGiq3NOoSPSp0YH/jraJ01E1s3JGXp+iRjT
JqxaeeL5ijM1LWZ4HgvF7WhKqJxTksY75BvmjnLlGmewPu7aQIvYZfXMs0Kp
LKHajLdA1qemhF6kPl+EgVk/RS++t/4FMJCNhTUoGxs9ycpg04L8Hh0vTayX
kmlUMEwgW7/+XS0xT4rlQOaWkGviQ3BFnRuAp3TBuCuj0VcNXTB+Qn12wxAa
Tvwu0tv8pF7hSFexWw83a+Shl20vSrVbiNE4bx0EBUdACvi3kOLTHWHTXXtT
ER4dcSmUR8XfYZoAMzgmfD4qFmojAfXQrqTXEAArW3OQkxEIuVBOh9EbyU12
04NAAscUnY+t89dFYJQdXS5KbrW6nF2V8MQOppRGUnf03I3KOC2RUtOIfA0X
zvaKkp8uNIOqgo2MjDEADEctnYc2Mvkt1uAF/x4oVFwOkab/bk3XpNL4+n5l
qQ3HeVMsLNd+Ah4YC4gT8u+AN/bj7CJR0V9G3JoRGEec1BtLf5QLU0RBW0ns
FuFvMAbu+Ynrlo9n3DE8NJGEweVNBAlzafnDRIXDH56qoOuFwXlJqGxRAx++
hqCfJ1c+cxr/GUrdJiXDfXof1yb5EbkYLMyhFgUCdTnFRSvNV/DSooWVEvOT
st6pN3tygwakgFWtQmvp0r2B9gDFnZ8hsz8QW4+SnKuvhA5HyF6ZyG71MFhV
SHfnBA8BKpYf6yzcdtKM6mfxnhE38rGn4Nzng2/z2VpANoPImXgAZk+Anb8q
nkyjzdsVPdIWxl6DqblGXb/3Bm5TTOC7Wneva9C/Tsa3OCkzHa7ZTRUjcUjH
6mYm7J3KeExem0+IETZkRwx8T+DNYbewQaiQE/GTSqP+oH2DMzXk2deS5uDO
YTGtkbiTxpx3Vj50fj0gXxdhn5vA250K8HleFqX+06PNiWSp40olRky3ut1n
k1OiKvSHIhiiTtOCNU5Qt+0jPVLIxCscDCvTweaqvSk6TAJy4VPU2ng+SwaU
uhhyjg+iHvdRmRub2m08HQ81MvSrbeGvY1T9hZr1L8+Rh0byhmnDRa+SY1N+
wAKGtoDPwzOTrc37Iq10nxKEAbeVwAfWyuIwVtbMC7KqE4CSQk1hSAcfn+1/
vINFOkd4xi1c0kMvCzPkdaxBbyn4nKg86cjHfoO6q1pMjhTLOUGU8mPkLoqs
ftATj9yeMrZokDGr7LPJhB0+/752q4WppCQs5eosXzm132xR2UswgzWc/DNB
1k3yntQpDexoHdzGnnLf8DKmMRLZIKrj43+LFLcIkxRfsPyWXLtCHAOKsaXq
pRDpWU/8PjMHukLdG3IBXXsRT7yEEbeuzZdgMpjhEZVwzgHDX4RZJmNFcPZC
RxCyPvfVbq6F8ftLuXcmXC/D5HTOxz9glmZfBKU3y449/5Wnc+nWvI9h/zOw
VQsQYcNUAT1SSNP/L6Khbfo77detB7wBbBNseVWKw+dtas1mqfCLbz2TPSfk
czlrVsUJv3BVzYyWP3kC7W/+JMEpdkoTk0kt6LJEN0yYmZj9hhGlmSU/KAt8
9BJmSbH6gfgjfpnsxQmJxnkrz6BvXl8RWWv1lBQ+6ZY8DRu5ZVu2KeVkK9r3
2tA/TEg6XwUQNdxWIq8alqE+t84Guu5gamY46Szrh1s2lm828fi5dx+LSSw7
v9iN5ik1ohGmhg31jQGO/97A7hugCGwAOZSfGcLXmmrfrL7miRCoGmiaO9f5
usDvUrZQf8CeZ9jBdAsGaSFR/BQlVxhN/I0FU041Sye9KeOs5FReETq9o18h
6jqvlNcoHBIYwb/n8Hx2fm5rcQ1CkWmmHEwPHnaHPj0SNGLu4wvnTsH+ce14
daMAn36AHfthHPJS7Ys6nbOOmFR9DCregWhPj0TyPub0lCbcqdVhaN6DlKMg
XNUt6sItf0rk0JUGgEXNlySSJrgxsgYvdIAX1NRhhin0DxClT+dPlZ9f3Upk
6MQzlB1ZlESHv7Zibndgdzl+/TGw1K5KGZEwYZZs9o/jSxQj+kIA2vHJW06U
iPTmWLTQJwsWRlXUI9R40IhsZiOwnB9Es7G36H3OHVis85wF54QcSWLdIXEW
TqtKCM/LxPevIBhdycjYuJ14yk16D7aL5+nkrgp0OsSSwVj+VXR8+MbZZEhe
F1e9d5LR2tv6I/lNjqvByghsoEhS1yVCd5/B0dyaHxi+KmdJ2fng2gzVMZVM
nMY33kyKBrWoXrCmzbeuJxY1zlo9rH+dlqs2SEVbMbS4l61j37U1wx9zL6T8
OiCKoEg3PvQgq7dy6r/qcAUEhQHfY01UE/vl6IFeMKZCe90+JHecbaF739dB
HcdduIT6XPWZrO6aovFtRGocML3uHrGlxIMUSgVw7KdCtHgy3V5N7clr0c6m
I0EAk6Q9k2fwk77EMU0GAqynAJUqi7d8LShCUgXYOb7UZSHOsPnNMdmlxe/H
C02GNxkd663WxZfAyej65YfAswMBcfHojLgjXmnMUSIHqQQ6cIOXPXeEmA0r
Jye4xV5cBVjlw6lTwErNp2kKsGRRoS5E079VQd0+hWSJkgQ3aTCQk2052xca
/MF9VX0YbGKPidR86KO6IPIDTIDR8Pt1z8zWGTQ1tU8L70oE0T8vEUNDqPEn
hQwxSBBtf7vP4W/sWX1jWh+wdmWqX3W7AVeLYz6yUZeOlndeWAoIGPwUrT5a
YczCNuXquG2KGrKhdpCG1edPHjvRtwZ1yl3pHrpczUQ2MJW6SKkXCiWsr5Qb
Of/myDymDmmafhycs/DtMc/1TwoHfkULQqeAPCWkQGme9RF47QRzOD0nieTB
9PIYy5ktzLwtpinX6huz7p0uzHBcDAbyb14QJZTBoMEDZiVpky1EcOnUj3pS
bRETwgMNwE4gjPOte54I2pcWpIz5yYIEWYu35CAYHzlu18fZJk7owLuTXKzD
IzxI8H8Drl/lThc6LvutM/Cdx8zAIrD4s4aeKbJtxl9ci8EPmTamwFU2P5uo
4wUVy8II6B6FIXNhsCaKOqicwHbFL8WaKjec2BEc7aCE0rUyL3nYd/B/sJik
Wqrsnal4QCLBeaH3BvlWZbDC4MDu5VTYuzmdQcJT5JgTUjg2j3s+XHHQCSYB
h0H51iFvO3N19QJHg+nX2tnUoVT9eT8WITLgCGELnolWb8FIr9ld+bGxAwT3
dbMnxMwfc2GTskP6jL/sD8MgkZzr+PP28AudESrc8BtWtU2mtzB0BHtSUiJp
eEr6qg7HkhRMpityLXLc2jnIevpDtTt0eCntED2icckpRk3vMxvPSmHUJ+Jt
ZlUh5hLnuWM8Du67C/SAWCf4rSKONetGJM0rSVE5POQW5UqOj7ttJwonDQqh
w0MXBAg87qChCcL/Ye2vSIV6NEIv/GYmZK6fSDbkpl8h6d2TMCSku/o7RtdM
TbS1u9aRogzfNyEHwJiqrDeL6l0F0OjMPVUQEDXuxxCgGdbN57G5kDw2HxKb
e/G1T9EoBW4zaIFbQ8fX1oyFtcSuG9GRer9hs6QldXz0RGX5feyK8KeOA1JU
buRki+eO1OwChkPxhHY2qzH+DYWEcwbCctrqDQ+k7IvJArVSx5TNwrWjpqDm
jWhicIr21F8lKcStjooYGl7poel2IWrfy9BMknF+x2VU1NjtU3IkyrhSQZIm
Eh42VnzhW52iBcCFHpxD8OTYdUkLDpidQf3Pgc1Kg0YYeHqpxbDox+3XdMNs
/jwCXdZmKKs6BDEu1OQWgVvZO5D72lMsP2gM3aDFO8zuKkutacDGSaaAsV4c
wJB9zxOrjCOCQiHkZ1VIJYGdWHIf4WAG8eyGX0s6ESrDOiTV6jJLkf6xPAad
OREbAzIcDIYjZkvUXPrvfiusweuKLko31Df4C/z0APBF85OyKRBNI4EpuhiX
pUUXVw7fQWk9X1O/HvApsxnLYaWILOOZfAO4k2gANS0XS1ZfB7eYfUSvEvJm
CJk6NkgBpFmw7jXtp3vDwvD8DyiDgyCzq8raD0ghlNN7q1hbXYFZ84ZaUZsx
RbJ5dpS1rGjgUoK3BmP7LzIM0ad/k7kHmo/XDaElIhIwIKbQ9QUalojA0gIP
MFAzkWqMn6aqBTZsYu55x6BWrvVuGk/N6pPgLEIiqVviv90vvBfSka6bzM1D
lEwuGAxjhghoElM3LDb8KFkvb2jGROKqu98DHb70QJotoG7XniRjr97K4Po2
Umzq9Ud3YG8KxWZ1CZcqsFANigkk4BmEUy/3D1CFj86OvSMZYwmaxQxSc3mV
PJbcn1nZDS1YC6EwGZ8U+BJ77xfAHNZ59ELCWLFgV2vlUDy9YrGJqUSW71vx
/wDrQgG7W8b/hElCa84IKKgQDgiQoVyeOyNFrjg2C/JBkbf+RoXvB+gJZNk7
yARA9SB3m3ezk8P4RR9l11IXVxcrisGmBTRnnAJwHfhW4mI6JgQn2lgm+irq
5iXPchPEreMokBeno6CsRhkVFpXsnPIs6J/H2Fquk25cLLnQ3Z0EdiseUF87
VtcUpKXoGYy/uPBKfbirOsg668DrtQVPcAkxHHQKMdEhdUFtemxD0m5/VWFh
Uv7WZtOBeJ7bjpxLL+oNW8hR4M9lw0zGX4W9nTfuH7cZNQ7irjCvs+5WX0w8
cjesqk4AdHPiQc4StMPbb4Xsafe4Z8Z4wNnFfGYbURcyV2BwSFpLqNSFRjYG
nr5homS+yZzllj4e8j70pjbIqILx/Q19gKABTg5nXaKW28VSG5qzTS/UTirP
56DWUW5UbYDZM9xS+h8f/W/sC4UCwGkiisvu/NdrS2dzNJO63YhdnZCQjjfh
mh3ZRlnKtnSBNhYfbf1HILsdci1VTFyjxsFTBrZTnDFaKBGAQtb/iL5/c2am
7x1kbEhUYC5ZMXvDPZQe16TOcPIjtn3KOy3ytIUCjqv4gUeHHvKc/YhxBgaj
HrPSCacjvihbpshGYYoKgntfYtOPF55Yct0dyoU0CCzBA8X2eosoIfbITNFF
CprfRrYgn896lQxE8JfUywLbvz+L7rDW07rmroS9FJoBgVqEAiYFA32H15bU
y8HcHoCVnX/xH00Qz1dusm2RpJ4O9XZGIHByJzjBV49mQlXFoQ7dZYiUF7i6
WVIxU6HROLxKSRZ6ON4cw1Bmp3axuSBsKERIGmQq/gKlskpxsBd5WRk+e9XX
9c0Inhq4Ht5YXyCL5H17Mee0WFGU6ccJfkJtONDzRa42iRt0wc+yrpx8zygp
QLb1C0G8kcDJYqmZgkVlTD9UWK3wQbp8bauukeTs+m2z6T8Zr6PWc5Qb9sHm
OQyhPe7K6/fTowqHQMhnYhrYeUotGQYRVgn7aN+eUoJWVvlMEdT9SQ1hxdw+
0lHkHYFg5I3eqsi/iCP8K9Q9wY67UCWZ2XmqrX0RKjmdvPmXTFNt1Y/FUYQJ
VwgWt2n/XgdgFZgO4JBGOTxSrn6sPz4/BYzq2bNhFENQXBXBB6cJ9POu8Npv
najAX1FtRyzWdQXpsxJAjsPZjMKT2S0IgwIjMeZG3K+rWnXZAqKHWz0D9INg
wAkqOqYuAC0E1KNhkvmyoD6nNsYB+k2sWqp/7hRvZ/fYuvRyaaD/xhs1TWv8
REE3+61k0E7bgE0va51qIwPM6V2G3YVFfYLj3yt5Wq7Hptny2dfVUsy1SbLb
CHFPZbp+a1In1qof6zXRVfKteEVddl216ECBNQyYBZOSTfHvdN8gKSVgQrmJ
Zfq8E5WRA+7SInisqYB3pDQuomzm6VgdVPSiTSFAB1a2MavqcDUxTJo6dFgW
2fr24r+bQgZNqCej2x1Coinkomm5OXrxQlQ3XV/xcxdol0TGKiNNJddMmKDs
bUHRxku9Zxpro3QbUKhKmfDLRMrBVrRuhVIay1QTfHSZsGpiJ5WMPerjbfdf
L3F+k5eBVe7366TxwRGccEFtVBUYk162dPELUqDsnNlWhY1yGnnIM5XkB11S
SQ+mGrRypjc5yx+HaJEtr5xJarZK8lkGe74/oTYRGL89FLl68p1gAsm6JMKh
mK6z9RCo5Fpoiob46G115FT2rhevaUMDTH0Z3GDb7M4PSoiP3dyUiG7NuSFA
HpJo8kVCIp+gM7amNMVZn3wo2z96ZtaU9LpJ/7OttczI+Gwy0hDNk6E+4zu1
BTgkdt5seJtlwtmOhkJolTb1EevIGcbsWBclKJDCC083aG3muuFdOUBIDbWM
FQFj0zUJ1xzbzzKGAT+mS/nZEiwxx72goQCy1xApSbJM9N6XAJT7nS+tOqv6
CemWjQ6XbTW8wSZ/+bK5vxcg7cyOk4Ewduj83n+g6mKK9KfTmNpOqJVmbV7l
gqRql9rHz4exIat5LMwEMKEt0VnkbB5NPlvE2HaBzA+lOjdyDAxsHRfbP/QJ
90VPudBJ06iIpoFsgq1kl/7prU2ye3UkQFzBbgFDGxuXkYPtHbTRtBgOQbLZ
1kYaJbIufvAm+sRu9SbEQk3kqeoAuaR8Ovc8Jk03Hv4Z9Ctk2AiIYZ1VNx5B
zYGusQMVNsDYvBy2jjIRroiFQfd74Ugqu0V+dShJM6nry5TfNiue8nhahocV
T1xaxeA6X7ddz41m2nLPO+L0umGraUiBpizuitrPiQ+F56rJvf2rQdGZsgJ5
D0OXnehf1qJrIt3hxOBu9g8x5u4uuE1iCJ4i50t88OkTBf23whOWM5HS9Rom
AYcAMott0USOZqlrYiSTpCEOVBQdnx0qPbMfgLyRjEqogfwmQUqIF9e7Lkf+
RFHL9Jy6stsLtsm7B4KUo3OpGh5rIwz9MkdH5IGbOAuRjaLWSHm6mx66j0To
I8JOJfhTXjciBPPIlFptyOl2jl1FaU5z2M2/gpPUkjAOyo7Tnwm5vQ3R6qX8
y8PrvkpCZacG9UzdjfUa5meISjlvSaCSJ2ay9aQ1twEhdHtvaF/5KS1tv0ET
t4dh2icjyKYun93IQCQvjsPvFCV5FWjI7NMIefUMxgSgpugfnc0+WNZ8oW3S
cqLH9NhOjY0ZdRvUe47mkr8sb8ZxhFYhHKZMgngSprgElyI+lPGDz0QC+1MY
hDLUubma8djHYELICklKNi1zDpgVBiNflTOR1bRlWuaxZMDIQnVsr9Z4AVE8
aFd6ejzoBk7oS4pLfxTdLkn2F3g+86zL4k/OPz53wyYtRd/ob0hIMo7j8/+f
1tl1aU8oL4CUARxXWw7zV6shyOx+x7mmqspdR1cdRYB0A9pi6J3PBM+FRndY
SqGFVOzbDJ/XTzZ2I4BdmNPeRF84mLvevo7johm8j2aWpYUzHzwrjbKi3NR3
EZkTfnEWX0IIR4N+wcbIDHJXZYiXYBUyGrpgvFhpRf00LOvq473JAn/RYKPv
aRGJhxkzvZx3ENS59WFNCtV3ZTu1vgsqjnoVpVWU78QwH8dOs9LUyBdlRD5I
JrUKGNHpLKv0HWVHDc4P0vyejiaRuMUJ0m20p1BtMWUbO8COID16DxAyFQw9
0Ky7dB0qWRm+Y9/Djni7TeFMkbiZ2PtjRHEv0lRHPf3cGY5I6U7sTsiGrj/z
qU98+6KooitmQ86RSwi+OeTz/Ed86M8WGSyxQbvUsjVMr/lMMn49W/SDNLt4
1Dua+KHjEkMa2RfRpOBn0NJiM7swqGxtVA9ZhiZtqdsfU0x7jwR+/RfmZbsw
2ocBRV6eGK88h+r+xbI4sa72hCP6tzMs1UWMOEQm+Xm8faR3HxA2Qx6SkX1A
k9nBBjreP7Bj3sOvHAR2QJH50khKTMoXrOq284/dQ7AFDhy+hyxb8F5rvVVD
gr2MixsNrGHTLPQ2wjlEWQNNRMvO2Gog81GFSLtChqKXfZ3GJ7ahVlH5xlFS
Mx885+B/v366XtMEIPzuQpvfssYfFhY0ormXXd+xvmijiejsm8uMFxqLfPZr
e5tLrQu4uCbAXXgULcfQAFlSDlcN4YUP6ocy2V2b/2mQHVGp6CxG5C5t/mqr
DmtRXThKnDFlJY/Mz6uHsObH6MnQn6b0fZCY+KLJUBFVi7/TWDlUmB1iCsoh
cpHAFNK8Aak1Pn2+/G5NVCfuOSrynKDX0UObQfeq4hmSAw4w09CBTl3mz2pz
Nb4NR0qzFQjEJY5OGFGhiWpth5+7fN/0Qtq4C2HTu4+QR41AEkolgMy/pQyE
fdQHuNkJyPx6QdtRtiMuUbaincSnzcSG3JyVkV4Fiob2Ed5eRntXUnoQYfPN
OW8SwIoBulhj5pBaWe5l9xgd6zahEfvrrb0aMYO6ese9OVzFZegHwGtA+lcu
/etr53eqpEe31XU0i6AO0EEO/tdz9hyQVMNHJaiXJVxofSsaNM1qPwAlVRK1
hmzyYyS2q6XeagbAanvacxHSm7gxQ5NSYy9bxzjGvPwvz62xSpRCcxAA93t1
GEzL7tG6EwyDDbvS9vgnoP9E+6XbI7+/DV/GjvCqGWsCd/c8hPU9mvWi7gcc
zBp3WMLrIVxC/oqXI++DKdXfUP9pxBvWWokGYZfIlGS5D8YY222FzgwSXKUs
lTBk8V1YteQtT7s2m4RpiwVIw8FlYSHe+6EW0NAYjZT9E6Zro8oitvqSFSEP
IB52jdNCgjoBCVJvi6UKV9J1rbIiIKejo/49t0Mpz0pDZN+LRI/ugQ/A85YD
ns2nQ2dQJU3W7BGRF1EmdHcZbRl8FwIv7RwHhET9h4T9y0vF9jIX7xCryheP
2iHdCS4IDTh/7BWOSMCKr5dWqwlmQf6sxE6HlYaLk4f3OQUWjTa82j/5c01q
4CyqS+9p8keXTLGAutZAVqrQphku+GQ4wYYUVTKmfs0mUUyvoQvJXNHRtYzZ
QyEIenuXCt+wlCOvjMq+wObOznFXtLqfJALN9q3+PxSghHCzwFyihV307iiG
Rig7i8SYnu3kUM49m/Pw4wx8Hu48BlAVqdHOtCOCPpgAhYsmMZEkfnOfNP84
H5YPzRv4+f4vTFhzJO6TlsBXG+pzWHScmDdo57oaHX/q+3XkN9Kvac06PEO+
ajrde84TP6A09bGigu1F8ilzL62m2TREuN2+q5QUv0Pm1Qc3fE29eLf3Xb3T
a2Tw12Vu202zqzYCsqhaYagHVm4Rg5eDySk+/rH4CFZBPFx3djTyFF7gbyct
u4qyWHq3i1YiILRiUfVr4uMfpmAT540L7CXsFysAj7ZG3AL2S2Sr9FFkPdeq
HKFLP17GvZ5ExkpI0sedpyiAtoxV2R4DawJ3hQ3sKGvmxU6ExKnT32xYrcoG
Lu4jeHyNDz9kIlWRoi0YdQ8NzB5mAbGF6nz/ZK7X1nx/xYj1/Sz+l/xNwE97
Up6nujBwfXOHDmiGSedurcQr0Lqv1bb1KBzvH0SzNvfhU2t+AD6n59Z+FcnT
QEsQ9+Vtb4XPD6cdAKKFf0gdgvzSNcScJP7PTMNci5rUtAIUZ7ExN9NvN53r
T5yXzJbRpjW4VsD70rWZEWKhvP05guo1fINZOF9l42yWjEjlbWV9hs6ZqmBD
kKWexTiZ73srEYtG0IyZ6DVMbi7dYf1KPv2DwBPzJ9SxwG9wIewiwnVdXBEV
TCvzmy07BkzO8jUOdTsjCZmIa0eNznX0XdOStdIe+ivPYhmeW+3EYYJ/bwF5
0sLLy2tNgL7e4ikxsOQHqbNWVcbUeE7TdW87ZQcYAndLmN7GofoXATVpofYd
P2kIwThzqXND/aw36Gd5sZ1fQo2rc+/t7AgVlDm58YVmO0Wxngx52aVehcyq
0IB7BpnpjCd9IQFB17z1bRYA73crSeOIg6Fz/9r4zfeyRXFD2X5KAhoG6Q3o
ORKdXYNc4xw3K6LewDb5vLEtYo+wWXYqksTO1DROnVNubDstx6J5E6irARqq
QSliaF2YjTU7+ACU9FGrY7W2J3FyRaJjjtcm2fA8av3xXzruiwlwSQsY5uqp
BYKY4SG5cz7MtQFhzG9rQSDc0+0Pk6pERRIw/nbsRcIHyRzl8bCPMWiLZVpE
LsANK78pJkzmstgFub8jBD0o2q91Ef2rGlMCM4N/XPvNvpdl+UIKaZ54KyC4
ZPuD+Poujd18yLGYoAVrh1wknU/GqGuoiKsCrYT53pVadPjettesB+HegQMH
XtEa/WJ4n2K0x3TrpzIMJ0bDWWVwg6Bf+kQnnn1UxvLyLMakWdqXKctDvUWp
OwtNbFcReFF8r9RJd3OizsCYHkM3Mkv0XnAD1NDy1YxxtA15hiwC8RydEY1Z
Tf2yuEPL5uiTHaIWTGsjc5QupbJqPAjywqjPYOu9wPj6HBwsnMO/JeEnw/t+
lXPsrDOVBMxNkOQVZwj4SrSSLiSXA8zJNVtPIuiZIHJG9Vk8g8MvoY9kYc2R
JAA5euRcf4lKQeb0gbBGWdq4xPK6e6DynoQ01LH4DgWdZwrEkmVjar4RguUP
5vlEsFbbGAD9ZDTcugbQCro5s8g7eOLDVwgj5BLZDQaSQFjkDLazwrY9q07A
UK4Li4N7swLgC6BnBP/RcKg36vKi37X/pAPLwVjq9XYJQyTe/UTed6UBWReA
F5i82FSKmsZJDDViQV/3AFpcORjfgxyNVeLqCaRB+BXYj/Okpe9oP+eCI4fa
blJji7Yc2mlQL+hCFZZn+48aaKoJGCZ3PwpsGyULnM0g7GKv04pTyqvcDUkk
K4gKtKFPFsB03sMlKt/TCZiven1Dt19KazNBsVeIKncjFWdp5BrEihPWHeQz
kab0Uj058CImQGGXvbg8619h7njaHux1l46sfNiUP/SxI5zlPm5uTyDgp6an
v8nG3K9V3wSqUdzQrXkzQD+c1ZT9HGP5merK5KeZzMXRdpHzSXxQzc22n2C0
8aKNQsqq7z34Fjggo38YqO3xC2K7Zp1ms7nt9/3YiCf1twutO+coWRSO7XQA
euz+o6dDfxqXXGyZO+2doKx7zT+FkGH+g07Q/r0Mjwl5oRcITj1nDoixwcjW
Rl5i249CatYAMVJRUNav2+AgA+Lu6/vmwOlizguD9OEZjK+W3FNuzi3IQxJ9
mpZtG6sKLcshsaHDDjP6Fli4FQo7qJBePWn/dZWcog+pVUcMXfTceE+DsySA
8GJU35S880k8zuQFSGhh4jNJrbiaTyJ4ASGPiVMnz/qw560yCCuJZDlqwz+P
kqUIDECqPij0lbs+fXwfU1DPt823tprGHtxUvZZ2dk2suFWF4+qg0y4BVZZq
jlDoHr/QWi4hnpY0R/YirlKVoTcnFWbeOPMHoFEaQT41rcawnls3FnB6Ol2+
60tg/JqekWwV1pUaEiXW94TUT7nPChTzElitGL/FUWjODqqpuBAG6UA0wMZp
9X9seJ09J17PNe/6zVsxTSoTwkUQwJyadfkTgsRyvItOTj+MC809asoCEYEb
rieLcq/I6u5RM8QO53e72b1dij6cMbLUKJPnw02YVc1Z32glptcvCXD96dQ8
MF4wCC+GMWPbCroszZ9iRFwVFrT6ccHFJiSpc076cZvN7P91HeEfqpfVRw/w
xySsh06AC3ZEItH0E5Y9U0yf5K7/QDEzmfznNQzErGFo1O53Bi50k78th1+g
MgvdfExlF+QweRJmud7dLzzB23qWA/wmZOeTL85kGWH/VRyJUdQ3R1/5xnku
NhLnjd6tlE03M5u/VipMT2hSpIPCoCnRV4TqL9HZSpv1NSE6D2ESyih3PP/5
U5SGIuV7zDsfpky0MJsskKt/6nlWi8EHS93eZC1W7oT8+bHFuw0hs9t2+9Vm
RokNhnCjw3Cdrp0FSHhYzCgoEnFhrmK94HZPKebU1bxfudP4FGhwAzyuopdP
BivqoNR0pVkk95c3j07wbzdp7aEMu2m4/THccmDTO2p+jrKOeaRmyR6pk68J
NXG3brg0u3JDT5i9RU1pErjYc9HMlEyNBnYtxSIyjbtwY9BTn761hBQDV+/6
opkQNOCBeICohDFN11BuPwXAs7BaclkO6i/Hg3AakF7ROyFYybv7ZQWKOqvH
1neUSuFLrvJppSHzKDe5E01+X2/r00YHICe556tT3Bq5PQmEkq7j0coiGNv3
LqULVxNa4+CO0ro1DGxQHEB3+1JlWxVYP3VLQMjMcDg0/rtezaIy2lXO82gR
xqqVlnyav0JxqtEFLNn7/PCB/JjoQ8YZ+Roj0LipwH5HdG1re/tqFRvC1Fmw
uM12chgYlvPtkIkc5Euj3nQo5wuaQ0eyQ4u9dr+6MqIjtg6epjlANhw0deEg
4dYzJr5qu1stRuoJ/UjjW3e0bhbG0WJ7i8ig+JSrIU7KbbcwgiWWZOFJF1lU
m4/g5XSwGuaCFzS1qk1iJjLk3oDzK3WGBgQo4H4bykij+0fF9+g6RBJLVVUh
LTG4zxI5EUpvqTjAHG8/KlQ3iYHG0IT9EN4zRI1bGOwr8rRodaagwIUv2xID
DGgjkjVQ+vtHXlxf261U00lXY3AlH/h8g3YMWWTqXwrjjkeHsTo74P71C5vR
PjNikHUf0PALKm0Nv2sOZqMMKdT97cxtffcVBk6TKh9vZYZMmGy94UC7UnVd
ZHrx/rQ92QBPfhLyDiKIZgrID9R3mhNjI1kcLtJ7V8waSQtHN1+1ocan4d5P
JpvS7fN91f6cq9D/0VMjQsoNUfAf70KvOH7fK9RRVGNIjYNeAjK6CGwj5R0R
nuqKIgZbQePtL3382OhBY9G+4On1kREbFWeJocF0TDnqejXXjW/rVqt5PS7f
JRaKxAcT9tYumkUQb5PvcTV2dmVtn2r6pCfw8hQ6ldmFymA8l/dyNNNm5o5M
k+L7Z5uk8Ub8GvJqsHYhnHJYua5ppYCubktrendwZ6KVF0A8ZHMxtYooBzVi
/Gyh5OscIVxUIdS+CnymbyzTq2eVZec85OllNqCBTC3c+ejgMJtOcLKl3Ol3
mzyjLm76kDSLiHRlL89EXPT2lgV98F5YkOI11cVMYGHbuvLgNZ7Anub1wOOo
PX+ipKUXKskzd2iXN985VbUIX2acX0L/u/8DFPRJbBOpQZx2DHKKOR5Oy77A
i4ZJrAIt8oILf6fzqSbBbLFEdQMdHMICyvgDI1j51DVYFUTcPT8ZaOS+Egnm
SH43bPdm6QVqedadkvGd1/HkcPro7ovUySoGLjgvCrg3HGdPh3MF+ijH5frc
8b/n0JexG5kPN2FURKOhJowZda4AM7uqg5ONRYmQ2HAr0vxcG1qdLVEZFOWR
HZcKqRzzpZnVEAaKf0tZvZFr1cpWY8ymKyWBoJDIz03/pkG7zuA/sY0rnKzE
Fyn4Vf2yyiqG3Yodp7EQXVWXax/UZLEoRMJya/seHtwShf/4G2GNc3GYD3HW
AFrJ2qgpA8j1fSQmCjbdiFtQWp9XLQAkXrOoQbd6lZLDEJK7YOSuOb0c2zJO
dZB+s9TrdkY8agu9chwexyZcRYHnod8NM+U/U4SJzOBQcBzRcKVfGWUynJzj
P6/WO/HxtcSOnA0RBX5ZbF91rsEUwWL1t3j79TcPNI593460rD9EBc4X83vu
7yfb4oXb0DnbrStu90YCJghyPKR+SLU5sOs+3zZJxweiNR7xwa9G4VMVAmEU
YUr0fh1vGjipbRw0QYKtF3tDcJSt4tClfEc7YNalxAGUB64+gZ6XpfMXmVYw
ZnGpgWCGH/vY9wdDXlN0rQkAPuoiYfk/wzu4ko/4OOm0Vs9En7smDWiQuEKc
qqVoJwnEBFLvnifhkeR9TylxTXii7wSYmEkHZnIq4Ar6X58bHCkX95I5OL66
/Xe1JsC7SodWI3d+Six+GHL1ouiVLho3G7gBTrrS9Bycosde4YeGw+Ov4YUi
2VBiZQSaGXw7eB8akc9WCmbwKKBdEvjWLRUEEpcrkCZNZ918Sfo9QuDoitgX
g6NW6ttwfHh08QhOSmS+Wn/OElgBAiM5qdiWTx0xUsuOrbMbsHI+1QiQv4em
nXx1ztsirXtxuGwx8pD6syu/jKIupZNmHPOsL+vJ/rd8hs7cLWhjr8SA1pYS
S8J2g7/PPl3uImouVRCYr6B6TKv8Spzyy5EVcTOqhm9+yEypxqbP6TW5Uh+Z
d7fHLspZdE0YszkxfROx1838FkTwe0Hpu12eNQ1mrtMiPon/QRPSA/cqQ9wY
+OMVVrScKdkDx2Z5QwXxrNPXGTBgcDfj1EAmSEUArpy9e9JHr+7ymNzziH3e
nLah0hc/YKOnXVB4n4VpVkH/SGIT7KH1YvJSr9ILIp0ABtTFvEBZiOIWF5aI
KzDAHkmxM+YdykjVoiLatfalq/5QrmGN8IGxHd1e33YWZTzFxVXiekudddZe
3MH8qFnGw8BatSHrNIXp2oi17KB+NWzh8eya/hDtJaMTcJ/VH+9gxsoUCvZc
v3RibmmmUNOp113WEPYU7xVeqEqyWlxJC7OU1S8xC2RyqQGSYxW1vWsF6dAk
GrWt77ixjS7tlDqJB9/ntDcdb+EvoP9DUWArwlpElvAjdfPaj1BkGy0Zvm1J
2C+2ed4amgMN/0fLVRVG3XJzodj7iY1Z8x8GmfCGq0/96haQCiVaaO8nbVfH
MrfJZOofhTmo3MvM4D739b4a4XnQuRqz48j4B8d7jnkDwz4zzavWUAybLaEH
cYoChyQu5HkzbVydjTsg78mHrnFn4HR+2Eh87Keys/OvoQOk1yg6xk1OHofl
ZTL9w0LBBnAIvlsShnZGY6psWH8WF0fpG3PMIowuWC7LKTPGBbkcRkaamMzc
gL2kYqbgT7rGC+FHixdj+WgZc+tbRYaqxR9Nbv0qiESsO/q7so/wydnWL1lk
Q7oKZ+Qdt80rp2YJFmkNKNHvl6ShH5bXgEvGHCxBwlPTjnATTo67a+42OQAW
rk2xV0Dj47ExDZiA0GwOlx9fi9hhqq10rfIf7oA2yAkzzDLPfK76mWFxchkY
3HRwQEsl1f+DoZaJ42OA1eVRpn7Jmz0V31DsJYOyUWk4JgEQfaGtb8vwnPv9
LjIyKLVcsmEh2Egtc24PZCKO919BREsCsPYdY0gyBPMANf9D+j55BNIaNhnA
nGyR5ZZbSSr4INt4Utz89NDfFJznFNG5DpOzEdq0LeiTUKGhx6elsWEKuBJP
7523oKrL7rYBrwK1iiVSuE38cWrBIzspzbjWNpv0nCc8cD5cMPkIzARC+6+T
y0AWBtiQqow8bLrx7+qT9cOh4LI6WyhhwvBSptq4N8GdweC+5NoUmEIKbMTv
8e1s8FcE2kPKb01NUc3G5MKbupuCOSlVuhTGLlZTI2ffbkndFNkX+e6EJ5kP
U3PnFujoiU2yt5QtCiJcI6RkzBkQ7eDpp5e9LAT6MIIojpNvFLye0K01JZMw
ln5ntFwor9WoIh3Ukv3Aik2a23mHcpneO3GEgnU9/33bhzqlVcbup3gGsXy5
LFamAug3K1Aic/iPzRUZIURLcjPzqK0Ocup4faz12iBsRivia+VeC6BPFEiu
0q0KHRuk4B28ajNmOzgMQKclT2IJVwlT6l15jo+v7o8YHr1fVem9zKk96RdD
DZT+6lFjT1YGkbBDVqPcOrza/OM4faU5vQLRlRf7kSfwdmbVifEvXgUvwKPk
JAiGyVBIrLrnzAradFcaNRj7hmn8UZSVUKIN/FzyD1ydH+hmQzRpsO7Tl2TZ
+Cqs+dPfAvDOTXNw//5NR9LuXJGeZ2vvEUmB5CpSzTiywZRlncS8ec7zc3TI
amL8JCq9iS3X6r9I21Cc0fwBwkJu6O4WdlU5askj9zBmJRqFyx/Uz57UhylF
wfhK4L5kEkfwxwond+Qy9/kezB3QbWSOFN5fOQwBvujCNNnfk7Uh2gzE8B12
5KpNl0k+daGXwM9C1o+z2iCKEmOHYqraRNzgYIzUGdjw577YMD12UHvWYPx9
Fnj2CuxugBuzHQ6tSQ9wncDlQBZ1uxiwJdWOnUtFWVWydgubyExfemRjg8iU
YNhdEd7Qf2Oec6VkmzPdYEe08vjL9GPefcVMGIIBiPZlig1LKfjseE4G3KS0
Tx19h95PxeEHWzWrj87EZW86lnPScvSlEgpz53gtQTrrvVtTA15pUuGRBDRi
Mu3iriYjShqJUXE7TFHMhMXrO28/hQ++/ZKtyvI5c1Qtoao17f1rz/bGhwW3
PutfCUTZKLjPtVNEU1PhBpC8RTIAITyoEW3Yj1AvHBbwfSaUouaKNrx/yeF/
Et43IfmLK+B9zEEx40/pSl9GpSIVqR8Tmlsq3oElG9xlgQHidLZcYb9db+GF
fCNecY11C/8tZey323g+igl00YEAnETEY5uh06IkTnb8tyY/f8kcQ7JbTL+9
NDBtX/bhGd35z6glwFfc4wJSzOLMWGzQ+bdFmpas6Psu0zlMN4noEHsd/rkv
9AwZ7n88bZ6boo6VDcWAzyPu1ocwxGsy6lgNoj6pZP4UQms5+SOAJI3GexQY
GatkZoH03tIlIoLC2KAgGNwBIIdOGBjJGLDnE+0uVyFGyvKWgochmcbpBpJd
vy+Zbz03crRGrVfO9tX3ihcwYAMR7e0hv8sox2u1nHkGOa1U0askHkcmBk2E
pwIy/+msvG3mPEUF+hYEJnN5kKdm39yV5tO8wlfeDPDjFWhT3onf+cjHQLJs
QO99X7Fib2u0b+WAnDJF2gvJbb9tbsk1FCnN+YwltmP9mxuc0KlArYc+kTpo
t0D0gOIl70c0pmN1I9J+vXMZb9GukqctAz4ifaxV6nmajmqpn2vQD3OsHw79
10hsWm3RqXlWK5qdtnH591omgG428o+xzvZMhLGnmymEt2kwqXF/iNlMIHot
XxvTexOBunFl4wwK79OorLDnkY8hw/P73p8423hexZKM71KH0CwGkgvPX0QV
9AeDYIAq/+VMIdKNDqH9ZuyLEm2B8pePBaJ89z751MmnH+lBZ72IVzzmPlkV
XgThRuBnTIo7PlfWq5TWn1WQAlvmpORXD+maf/yrMVjsyEAVP/qV4YWiuo5B
aYbl7SVzRbbncakCE5JLthRAGkWtH12dltJF73t4+q8Nm94NLlL4bLrs/Giv
PKy4J5xyO76GWd91BzFnHJxDsi/CizMph24nAZJLqvMkvAcvWp/Ae6/qA8B8
ZxDvv1SZ0nR7lUN1sMvQfQ4lcJm985y1VUFfnoqJj0SQFTG0S7QbwhY6xsPR
sJk/TaHGjzoC5ozub4yxJNCti+WO+vc0fLJcg7mCotXAlXLanPKifGpTANDN
39xfjj2mSsKQyJL/R+Z4O6VRun1sSXRbnsmvb70lUKnHw879RHlwIUtBDHV0
of2kk5K7ElwgsyQKWNdA8j0TfuyTUHAR3XXYq3qA/yqsdRDkomR3gz0+FA5G
krxrMOWd+WFEIUGpu1VpMIP9yEMFXQHEs+RMJ+4pbAgdIU3mNuMSNhzHbLY3
t2D8WS8Yj9KxBE/nFI7F20+DjCs3kj8GfcFe7jPgrQn/i1TNZCjbO9O3hfjv
8ZO0+B4bBAbvyvjJERE/zeLlR/JqdBmURXy4yjVpFZOkL1TKl03XFxp6Zboj
B9/OgiTsZv83UUoKn8N+GJ1Tp1Fk+qdkCbaB1ikvWks64QeC5iTFr82b540Y
08jqnsl5S6rSElumZCrgXCYxepBjY3E1B3qzKVIChCSwDrwjS2d9ysf22KuS
gRETZYzngjPN4kqvmSMNuv68TZv8TRONBRg9kqww55l8Z6bzjYyWbKaRb3mB
gpt5oc+bUHdmDk+7d1cdAqmWJKXdmdC8xlG0ZuK897+jh/Q/ghd19Iu6Q9Y9
5qbrmM8g1pc09ubCTaZP1Lk40kiRLuqRwNQuaQ2FSMfdiHw5uMfo3GCeEmyr
qoWoihbNmTgAgDasLKxBoueJsESWK/myDReJFoHpEBzQydykrqB5M0AZBSSO
Yf92BAdtbdIzb7M/IZE7dx16mlMPUWoNkgvOMwIdUEynlLU6bqscAyUCD7mE
jS/hLEUHxO2lTBRD+n0yUgQQs64wwgyG0Gu3/6rRuRfiVsMpbnC+by7IyvVL
Mk5VZ1+6jeD3u5vJMAooW+BZwm9DOoqBsOH+aakPShatEbZsS7F7vmSnAOnm
VFPuAVWnXcmCd3wAnriBwkxr84x+H1R+wPu4thaNPoh3fkD35cKSmExOmML/
zr/GJcxYKCEhCoestyNzjkz9MmC8X1//rPpJzVE2onWLpkvB7cBArDvl8Ge9
SB57QgXuD3jZzoLakZdK9hvqvH1Km/TahafaHvoLr5FQZY7rDjKYlXiT81DE
U961ARVGe//nDwFGf2tGheB8UJWyToz59PxipArLfrlDyl/I3TdNtrY3LjTS
FbTggkHifjNiG5Lv3Gdlg7Hl5WIMLcnBJSXcB+Tpkd3q6mlm9Gl/oTLEkE6l
TdXSieUYhxuCuqBirrUsI9KbEwCoRw39p+dem7Z/mLiU1tfvGfhluxvhIuiC
0/hJGAvUZ3GRPeFgW3xa6PvcbPLGuvHxTNszsy9hqJi0TgRg4CUe4UWIEhdk
bzfjVpsCPV7mB2B9tpRZu1TvrmkrztKUArbBEF43oWM8sFNcdI16c2fOhYtW
SeKclUJ6sDbGs4Fpv4Vc5Y1skYr71D/2IqyHowNMineNe7Chfcj9rUYwspJP
ui2uTAewdR0HOjXu12xEYBJ+ZL4YolKQliEONMW3I8f2xpET6kzXKXF1lwZB
UYFD01ec9cWLuP7TcjxMndKotJcAfT3q+ePuzE7dOksDPm6x3w4R8LCk0U0/
ufVhgZpfJRci0UWMQE/mTYD3YqCtoTLVmSV7ZcQF5GkD1UmumUc+K9ekZZ1Q
sSi+ejoxryhZPk6JVRWIzyFQ+TcW7FL9WuZbTNCV6Eqg5LBKAkLm6dJ0KoEq
1I4BccJzMDc2NF6l9z59qH2m4Y2rCRK6l6It9cmaNaqsKt5dCO81ZjTKpcet
xZI6cnfYDR3rju7NMtT0I8Zzm+kORGxU8RHMKxxotvyyhARWdeMQzNI8KB3R
z6ezp0vT8JMDzIT/5p/fzpTfsMYWVe3fMkG+Gx/t8uB5aKIQ/KsOYBFOYixT
/9fDekm7LLuA2YjqkQIYdNjobOa0abS8N8y/U84cgB1xoEHF2AupcpZMxQH1
+iOKmiJdxYXg8FRrT9IAaGZ1VPwptjfq3JNrIQ5CYLesTFCu65MP0BqpziLc
7BOx3E2ZmOJIMRPVF4HTGtEhLAG9R26UH6sAUn9vsq+fKWZQH7iJGOiC/PYw
9VjVIRK5tM2nXuIC6YDWodSFpmIuL/XbstRFlDukn045gFOfYD9LobtXLSV+
LOZNMG66G5cK7Su0JRNrKQ+2vErX7hoyYiI0dB/DEIIBSxhdOEvdfFyG9b/j
YGtFGAKyVw9OzRpN44D2l4O1t4L6okArJ/YrqD2uetIvDOQyaafMbA5Y1Veq
PGvLPQeQwxxQ4deOgq73BwgDjTvFappc4VZ0r8TB6hu9UzTSBANXMBCIEmHH
GAEbMnWv+LY8djj5nwfiy6uDlM3Rc95KM60qP5VS1HA2/YnA2CAaCcITsn5j
pfYTeDfumCswlWnWTRPWV6bXH21JX2R5FhKsWiqcCHuikzAD/aNvNtyRpVdG
0ilVL4ODVd3JHm9DZrNM5jJ0v0oYDslS9/pAGm4c4OFnXhG0pT/4K3nvajIh
UDZuCv4JidRuqvyO7/9Cd77J0uSKuuNnTunDJ+4Enj98fZIQoTE5VxFbdKea
fOSf5FOqHDJQnVfDQwyY0tCsafK5S/+7qISogc5AFstDD6yg2dp++8pveNCR
TyEJsF3RHAC8uisQcJXUcWb0DAXyeuKomnfm2N/0meLskEyKCYDw2RV1JmtN
APIq0YpC6gm8lb1UFjrZ2xtromsMuFM4JIsMEeOlPtrx6uaijFQ6yH/Xf9jm
p1TNSO2MGqDGjcKOw0G0TQxHuquWCSMESPHR/PAkhi/G4L9uk68ZW4DInK/8
WKhAnIDPgtnqrztfoczpKHlJjn9WVBZPlJd3wuvHnI1epPEBkOgNLVtA+rSG
pVhkYYsqSwigKFk35Y8B7Ho2YL6N7Z6S7B5bSGo0dSanUcmMHRgm+FHsw4FX
ydnjsJ6QLsWcc7XlTrUtg862VGpFbZsvzlzvGCjxRrrWFZQVeK7fQdfJlRMg
G+F6a4FAHjgwJ1YPH0dBaF+PAbsqfIVkag8a4O2uGf0NttaH2V8WvB0l6OyN
9kOlITvt4waxLHobxg1Gvsekd5mZLHYrZ7hMJW4r4MAI2n+upxC9uguZrin+
Gi4IPbDsNXxlfwNZLvivLtqhL1wCLhlgSNsni0R9XhQ3ET2LRHKOhDfXAEdw
V4aQXF6nFEArp+/7EqdJD69RK+qI3PCo+ThZVHkUXdDr/2ixOuli0qgxtZzy
mPPoxoI+vwrQBnqcC7JJwP72lxwp0ge3N1J7TTPzOkGCk5sHnnw/ABuis+me
57M8Qfb0DtEfXZ9v32jRWOB6n2GFfBE2ICv/OJc28TWa6FJlvqQVk632H24a
DW9hlVzrc1IL4PY8GE9CuTpbxElEZQUUrl33kYmqzSiCk19kqwqrZ4cJIDD6
aCcQ+JTpq5z/Mnxz50ghp0ivm9/TnMcA6IzffyeaUYwAZfTUo9gvxglUNrrI
KcdTWWW4kgF7TUAey2/D4qVUIPgiOxMY82Xnij4WLFE7D54YTZrwttcTDZpF
b2cHYIEfu0WzXGGKhBQK20LEQYfneWWIqHwXX63v/K6Ln/lEsApta1AxmWg9
RazJq2jFj35i4EH8H9XWiTjRYVMgqG4YoBbC+vIwGBynznlyYHW60aNU1nyN
2uVzF5r7ah5wdB8J0b2SVakM96dCMxAynkd8VvuKbno/WW0dvNeEwzR78bXT
Y2LcrXMKjBfIEIXtS8uzHopsk3Qm36cG6FhiDIkrtvNd55P+yjza1nUUfmrX
ABPili3pO12odwe1oVxlUdiaL3002L316d3w/3YuE4pWQ1saRYXlveY6L2LC
vnLWzQEOG1XEkzWaJBQSOMWdxWOLTkT6VkRxj5Lswo5+mgjap0M1V1aB1PmQ
vvetploEpf7EtE21S1ZTfd/CqNUd2agudlK7Obi+9TagNezjYBBp7SKDlTq5
beX4DG9buwdraz5Cy5HGwO69BzG31ETgvn4yR8Dx4Aqcce7mEa7JLVfioKYr
on3nV5zb8c1iwu0q4fFcSVlp2zESWezY0CDz7XJhFOgRczKgmGSRHAi7P+V0
gKMLUzOgEYyjt5i/69lG1nyX6zWYMHdBqKxORpP6zwmOtB1oexDQgI+HRkPr
YPfHTfabObzUiizcDH+MyvJCOJXkwIhCbBKyulATvV0FQ/prIectVcIO1EMK
dww4jMMrkv6FBQm6tf1rnaiZiTJAlzKTQXMhKgClAnSLCFey+AFX3D5UsLG0
BGJz8XK6VDMJQxVsZrzLO4Jc99Wilk5xCqlgnzVQIqsR7fTUZ4en3j2HAbTA
1iw4+AEfkK4106nTSP7HRBiF9uo2RGC1NRCWb2/jY/g/EYSpK8FRVRJ99tEq
TlZbzzfsWeIPA4l/z0CuEG/GOmRzxu7fbb5eBQiqZXMRJPOl4ZYpovAk1gco
NJL2Hn44dPbLnL6acC3oabSDT3FjY9uQ1FOa3rRLuA9uEto2P4s8ntxIMjf7
hQFcOWvCgvH96R3XkxrMM3u8jV8iF8v2tRGTCMEksPMIqsdtX133+EBufC58
L3Km8uWNs2SL917H020Gk+Pc1K8Oms7kf9ZwU/AiB/Wu1DFtLwoYnAt5e2Uj
01142oslg8xe81CAtg2mcUj4iaYMh4MQ66UTuyj3G+93U7ni6+INU7SOLsa0
TeV7Xt1gdiPxmrJ7XgbVuA6c2QemLucps+Fa+YMKbnWLFHr1CSLNK08bGeF8
tF4XmCKg/ntjw+PkjCUKNRMfWEFM/3i6q7jMSGDw7DqMJTCBywFrcv9bBb/2
CuNi4lGSXpmRieE+lWXvEro/RyjlJW8THJl14hY+vvex1txTHe0vl0dolfoP
7mD5lBY0rRtTSrMtbOd/ThrwGG3zv9T6GzFngvrporNWfJs/E9YHbfOaYAsT
+V7iqerC1O5OI+tErRvqJW9beAP0APK9190mbRsKSARHro7biS4KKJzUqxFv
dEqY/mtjcHMqUQWl5VCqzuKSCcL9gkKyOr4N7qLipgjRyDHT05Kf+SRVxSbL
OIXd3GwqLzJfbhdoVcUSfyt960UAM6C9AJBoYkj7iS7Q4UFsAmY6KhoG7R1I
OOCCae0AUZG8B3tQ863HLnKXodjuDSPI9cNMQ615JuAMbL39B0kecaMevTxC
Fpne7M1nuEmfGcVRYzDLxlRoUIMz6atPRhPeJl7PmPw1hUSerDTPlI86Gf59
g57L3EG15+5LmiWyyJ5OVA4ffoSQ+FNltIVjWsoeon3b9bUSFN5BVunUdPr4
pDPdhhe8tIEuUWoKTy2i2ohMpj9U+ZslvnCzELnYT9ft0Z+s4igZGbSZ8Cnb
StmlYQToZgOlbNeZPHvT0JBoNlsKGW78J2Kw9JvrQqjS4uhT68IrUHMaynt+
BcaozxemlRIAAmKf5C6ZAe7ABPV9yxfV+YWnMcXylmE6KJRN/HdgCq+0PB5+
q9oY1YMBlrPbJM3q8SXQSqNtoKWyJyQgRLtdEn4NsdeoXRTP8vgtmKSyZTiF
Ffpm2jxkskAzJSHPuJnoERZR8O9OLYmu6Y1ga2M0S0Wg1A360DRPGoLTbh77
hEhJP9jcmfhTuOzt2ZWuUfPrewmHaBwCvPYVbyL/PzL3XjLod2BUKkXGyUB2
hj1xXp0YCwKs2YO2kxHyJJabKCaOPYHu92FsFsI55svhlGMh6cCRnQqpkTkO
vylLOQfH3fyX99mUwWi1QTzvD7No3DatFBGzJCtLOg/HW9SJnkBKzoN20FqD
ZdZRVESi7jsbcuHrq/HoWTEaECclLMDgu9LdVg8jyFoJWMYJMNMKvc5Gr0y1
l0i71YipfxsmL5uoMRaSiU1buqsawaaUnxjqWdF9Yly01z2v9ZitZfB4DnTh
I85jsxu0u3NIKv3Wfzelj/0FxHYk1IxDiqJBviYtgF69nJ22f2pZB/M1RiH0
MVdr/y0y+5WfDES7JwDBubrZ96w5Ub7/HGc4bmew3gNNk3p0nM6L4/GjkRYf
nNvBCeAeqpUHo+LP8swNQBF/sFbdbQmd4JmKxfOS8GSoC8+ImkH9eTpExBYW
uKmUQgoBsoSOmrfKfzPPUc7zY9SvDo1nqCQLGMuezFaOqqwKCdDsjkTpI8/q
vAJyaU4DLyIyFDR5sB/NzIBKnusVij/GVYti/Yn6eXa73RJREzc2Yhn9mKNz
2VfyZUxY+I5msv2DLdeM0sHfeVFuq54NhiI0uz4UC+u2lhXDraBsH3yvSLiA
4IMc9Xc1njpmUsvsgR7o+h8c7lrdR9JlhbjyWX+Tvx4LuORMvenMhtiyIFco
hUJGrDEYAYc4fx9H2CbIjBuTlU5Yb32NKtalkn1qBD38nAkPbUQQ1OGj1TsQ
zK9nw9m+kNmD1hxs+WNsfV6TLanL3wLsMOj1iJCu5y9zJyIZC+8MCBhTwRE8
oTE1YFD2KLgAx67frNbdCGe80FLmPKv22qqmRXFirDfTDpE5qFGxTZCWe3Nv
wRWdc2VX2NcLxi64waC1cplt4XzW6/leHrgiRGLhY+Nz8eodNQLNB8n3scJr
dOAZYdl4BEbcUf8aQ22xLSFyBiOhzaHmmkGa3nYKyRbrfa8OUStvJFwkbBqL
1dUHYVUSx7Cze30XcjBIC09gJ6w6iun/6D+di6mopG6jNXWqXxliZNY8IW21
URE/owN+nG02Iz9lTkB8tRJwE8I3Sc4t82zEMrdcxDM7XuaWPQl+bIfOq2of
2H9kkKZo8PaGP7FyVPWMqraFSWkEsnMclQQzZu5DjDP8ahwmx+g2zan+Hg4w
OsUnloeWnO3x2X6iGSeQnI08PxFRQHXHNEnqDlZWtd0owampV0+GhFZSLKKU
DauCnwoLA90Pg2UgT4d5KK+yfEfKHVCyGcqRNiOWs4WYiLYUx30XflHjOjmK
l839AMQ1AJ32po3dzsJ56wifue5nRgUfqyQAOXFmyPPAGYtbpaJ2mZlC2Kg7
NGr5J2Iy2UVCmZu2wnD9N7s=

`pragma protect end_protected
