// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1n6sijSvcTUnqXpfXCGiR+JkmWRJ+fkz4cQm4qhfwMMMKKIWF+DITP1++T4k
kYRBF5XXI+hIu1O5TWgb1xernxOMbU3L2JOTr6K+bUX5oq7k+U/MJiT7lRoA
Dg7E7Bv+yASCh792D0uiOUj5/+HWSJsYzDaX2/V4sdMcsHrx10bi3dQPke+S
pG1QUnclkbxi8anXQE4Y3gsU6ilnBhsttYcPOXtph3ymQlwBwp9AMZQIF+gu
aPuPsWuz39ntLcmFfIafgsCHpzrdEUvPbcHlwj8DxpVAtZRHtiyF4TAX420Q
FS2JJsUtgfRYcTPDVBnE6I1hp8Arzrx4XdN/+sQPMA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RNUOH0P+spqZO1nAp6Vo60qmP3L+9JxVQlXz/6mf+zZ+i0o1RXJvIqbGn/3N
/Y06VZjpUmw9rsuJNc9EoKTavGhquNOpg07wDEi+L8UxTU7IXDRkDfzUI0De
DyfyeHV9VcJ3Xc3VabWfbVRriJJjt9cJxIjo4lvplBkWghKIDLUhXUOlByyO
y73/TXUu0H1+p2SEqx4T2xOsTf2bH6w67ae8D4kT7vB65n8sNwulgt995ElV
c/qE3FiJ39zZ4SO9PgkPq/A6I9kJRtstjPcBJoyZ76hCM8dnB+q3GVShcFPg
zIQZL+b2+GzwKpuD18e7bigmYY0Spgqi7gIYu9zqNg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IJSmRvozuaNn7YtUOYfOH07e8f4+bZTr557b7QTn8vgeSRC37UxMBWZzHFlL
h+8T3KX7XL3CzlqQYhfX8Yd6idHur/q/nfwrYZjE1VpFwISXDhHgq/30SPgG
p2OdhclOAokFZau+8d/Do67ohYAUgbhVvInBYwQbfqlBvXX1du9dc8c9B8Gg
GFYmS8qi5vq22+JopxxZBegyE67Wcv97vL5Tsv2Amw39GXj5WtmhKvJ2L7pv
9eqMukkZT2BtVJK33+fKGrxjuNu0JbP2RaZbrfhLMI50/84MlHjMKHIacOHK
ZlZ4EBTXG1SNCzNXnPDxMBr0OAVlQMds5Og7eK9Hgw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tGTbOo5SgAb2zMBfuLkOnFBUGiiRDBQFiTKfxFlTr1Sh+ciOFsraRCM0f34y
33rkfw3rSrQQeH6EEc9zal9JCdEp2xBDCnYeqHPdVVo8rfwb1IpsQO5MphTU
zNzlt48t6FO/NvVOwc+lwCWFUQjjFKQ3uwvnPhiG1cFcDJhVcwk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
xzy5TXGYtW4FzrNZAklAGWMWk8zfjtQe76vEGq2j2i6RdGoKyLG6EQ6iFAOM
quoI7nW0TzOQjv7yzrx2TCnN98qcJ2StCaBjcvzw7lHp68DZfzN2p+t2dm7I
NWXkD8xm5LA5+5Sk/b8F20FJnvWzOZO4oz3AWgqKm8ITlDKc6N12WxR0AMQ9
+VXe6yJpmvBp1kUYPFBvpjFua28BXqJvaaVn59gAov7Rk0NCdIebPqaZGkkq
KL/gcn9tu6q7ar89pa6YIhTDoV1gygAt49y2aAnIFfzWOuDNAcWBbnKqZ186
SmCbDKVfVQCOECpYY822Xq1/eIY95RmYiNZKXmXiH3U55HGivFPACcVPJlCi
7evbyRUII4rWbl+YF6KfHL53PQWs2evWvLvipLAMNBryW2UnrLtTIoke7DIf
PLlf/6IrSz14EIHKbD+XC6iTZQ4TaUJhaxujIP9Phgqv6145u8ZAOq0iLXUk
CpEHJWBQjYZFevqscANFCZaQob26TDoz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aKJ7zvDkjH19xlmBCLvVsl0Z4z4sM8QlVCrpBkIM2Q7QOpLVyW51+0ZtCZYE
hiTwocZcQDZIbSFC5v5aXTL0Vp6IfM9VY+P/u3Igms/HP11+Jl4zDIKCd6FA
OCj2lcRNtsbj2mkIUQ4l1AWAKffZCdVd4HrMZttzWbY9sEgCTC4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SsNl8SPfJ3nw7VpvJi3PKnR0x2XqD2rVLGd2wxxKV0vvtHeBGA/6TvXudT9n
qnbsteNvr2roaZItJ3rBqjkKITLKJ8IIs0SXnui3Yz2b6bbrGIbyj600BqiE
vsT2Z7G9mNB9sZ6H06+64sfSsOXXf14wVhuyp6qtEDv6QW6Lkko=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 976)
`pragma protect data_block
JaZ1JrhaxgNw2jpLFDdFErsYkNRlMNCuEvTSb2R7TlyW9H0ZWTBJznADGyij
OqOTFAioQ5lIo3lliVCXI7cfhalFwFe+rmEhnRwMfhCRjRdn1Lirm0/qSeSx
wBBrQL4H5tZvaasFOjUKl9HBp/IbWowRaHwXuaQ4mqHBwDPjYQHdcVB5wqcC
qJ6YDJI0HZzISUnCAC9+93g3RXIk+qbn0xbMiWon4jqxhX17FK2E5dl3lSRj
xqaeHgewFsKM1MOcBtvIB3gs6wDpzmPEGuHjSOpVi7nUpX62PxBGYICkLyhJ
pMru78VkrwOQQKm3rIatj4UBP0a++zGI6V6GCZMkhP5Amoaouy9KG5o+ltpz
CA81ZzaZ44JoWwTovUbQZJusfmhoTagTl7Vi/FhvpE2EjiyekuzJrS3ofYyk
+x4ORvwgrnGXbkQ4U3G6Iga+mX3EeBvj4AiVD6EAQpD9znh8Z1cai45pLpCc
IGfpKz9OTAQmOuikHT60m809RvPZTaDLI/ECxZIgnjeOwUW4jqkUNMhs/MM1
k+TwFPd8I0S0mB+6ZFcZuZQmxV/QMoS4VNp0Txo9v1dTX1ZbGfPjyyYeTHcq
RoS0DUD1gVHvY9rmrYWvqFgF6VGL7PTgNZIH953Wy8wk6KUvZ3pPp1rE7Ig+
T+IxV1Wn6d62eWXBXjngMhnM/DWSIDvuco35o93/Zn6h+p2vXiarmw+2lxjo
Kw1WAoBvt4idTB1WfM5xyvslVXIbJcfUL3LiWArR8xTP4LvmeTq/bzUayAgC
xag6pUzup4IgZBf9anyBxoBo29PcIlasRjefKU9I6w04kuUI4+ytp0Q32xpq
vUONlB3U+CviXg+5SHTwDmLBEpYBU1zTbZmiZZpPT0SnNPc8Tp45/EtOTi/5
433mvv7QPtbbUsXZ1MLgtxw+s+fQuO2sJ3L9em/FZh8ggOnW4Fp0YPBS1yjx
DAf3GjmMxQxSyj75h3LuFOgGb1elUtASqNbU4akoBngVZ9k4oexYCpTleD4g
/6Lmw4rZJyo0eER7FO6ke/8szgcJz83GB/BhpY/xQecfZo7+IBNtHdiakZPI
7vw7gISoNTGGSPw2qYmqLzC4VkNRwcmJs+jfQP/72nqvASdvU2wY55CV60QL
GpFhGgNpd4lqhgBGiE10LQ7u0uOsdk72oHGjsErO5ugt0U2J65+G81IjXY0e
T9YOa0Bp4M2XVWIbMbju02Jlc/9sgm6hT4hPUurFnxm9lrOdBuGV17jxToA+
bYMAaOcmcBz6tSIL9UgnTMO0GqTXn8mTcEdicysnCg==

`pragma protect end_protected
