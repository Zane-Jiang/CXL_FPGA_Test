// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
R8pqDqIh3NfJJUBmOhxZobPKfI0+XPf2stQWdPg7LHnT6W1/DYavZSGYZ/Qn7TYB
P84gF6VddayzOBtIeO6xaMfFU9wndq6CRkWN1WY5fQZFRupO3JmwhHxG7wZ8rO17
g9io20wavRVTyrs1Z+07eW0/oijPOl8zy8b8KNt4CwuPEBvO2QZV/g==
//pragma protect end_key_block
//pragma protect digest_block
2GrAC5VNmHPqo9tMYnXpWBEyzp4=
//pragma protect end_digest_block
//pragma protect data_block
OQ1LChLRTRtkuunwDlulReCsQTER0wFguBdvw7RViz/mL5Z8vomrXJhYXC17v9Gy
PULs75ykaRmKGrUVKONN55rDaz3RbogOzhdg2LjFSMwFLRjumedS4uTbyMxkwfyP
Fl8de+i19mwsKtU3PCwEm47peomBD6ZfnkYzYSvi31gnWjJgLUd3pzRiv7xFS9M+
Xm1Bfi7Td45A/X1r6l6onvoXbFpZIjC7xcXx5RvhqGnZvAGi4hiGu73kmjUBxns0
Pwa/xH12zic0ohZ2z+ebBgC7heIiapgOCExdBTGNPC9AIQJFzQcfgvhl/S8neRs4
iZB8GfHDxMt5jivmNj9mvaZq9vx4qj642n/rHNsgcc8/AOThftGyltR6DGiAlTY1
CJsS/DGqY2aOIoPakfthJ2IDdrV2H1q7x3PDrfmpwf3WXaM0qxkBwraet8czNRCm
nM6cQvSx2bU72rXVOK19MudAsQ7Y2c725XIpkYhrgVy3VMybtnqhYpFtuUuqKk3Q
JD6Msypx61lMlN5DB49fviAQ9cnKxhRxUDrO9qFLFrc+dLlFFtjBu8QuXDQcW9eH
YskIEmxmY9ERBT7rIkJDsuelEJJqmFMN8fMVce9l+X/gr396h+GveOe3qvsa6qpH
98UeY7S31vz4MlHCwoZLzoaSNGkDdOhwJYhXZ1yJB0ggDH0+CFapU85nwrmw/GaA
TUoVhuWAs1TNRgbnBmtGYFRtyFzjJP7t85Pqm9TtjvvOqSAMyRnRG9p2wsyBxu0d
euiCevDnxMsuHZ3EVTc4/RShV6ugSNVDYu4OUp6nVDUFIPeCChchBP4GsoecV+5v
Rj8YVP+/KuUVf4+F6lsHO6WeaOcRwOGBcdSzOkUYffNI2ukzWttI1TEs8PiED8aG
C2SlRhTLFRpr7Ll4uG4IN3/+qW/buyPb6A9GJFHfhQF0mgrhPWLtMjLnmF7EGQEB
zDrsKc11z4aqHqlTWew3y6nlsMEeoA911/hsXvVrRsFDvm6ozoQFnlq6Hehs1GXy
mMg+NMoojUC+20+bqxwBrvICaLURdw2CVUvufqxZEct3ulEVPp6b82RF4+oLqqaM
D3vZDta7pE5O6PU1SygniPTgsgPfFy6pYyskAWJ5sEbpU5kMTxiG+U0g+NlRuaOb
oow32UBirmm0t4VPeu7pZJjL5mxgvOs8C2KlSAiL70u9pdV8jfPGoIdtmuhMqhMV
M8N9GIkZSwWfiNPvq0/K9NJPWCtbjUesIbMHBVm34oKevM5l33cXbZ1pLhxhzEle
ShEX7qpd3Vry1GGcBzgqCZ2jXzuXXaSmg1eDcJLZM2TkZTThYQVyZ4W8CMa4M4ID
SBIGCe7JCtWP7JdA7ZK42yhJv6906i29JAZ0mS8PO69OmhFOgI/oIdtAC7K6NS7U
olhLnROLn59zQtLp79UzlBu/K5j95KMtEW53gTanBjwhusoCrwp0u8nHUZhHvxze
xaS/t6tFSzM1jKJZQDTw7fp1Kmk9iIt3KAOWbjQYfPYP1HmTRuiIVm0evlAwG8fw
WnpUhKNgF0b8EAJSpiE+Dab6WViFA4xTo9rUZK4Cp43pZC5Ky4okvVM6dTYHuyHI
C4VuHaGsG4HzAhk5cEIF2ktEWj07trXT/4UphsOt7aYW0yOE2NaXPn7vzL1Tf7H5
FFPlBlVfT58kOwjVgPmK3WNQY8SEU0GbvTDcnPJOr6tVW/IJFV2nnfIi07sSZgAn
AcKzTK0YTNB7uLS+klN5cM4LHHRgy63z51AVrbYKX30bz2A7kpKRtX3j9e7FDm+X
MnJC8cLYryemcEPMcKVPbAcQCo81F88LGxZPa71afCAdtHBiLLFOiwej/mElmcWO
Zsp8DBlJ+YwxcDFUixDT0vizu+S9a+uwmWnLqq5yRPL1MJX6EVlgMOfdS6D9M/v6
tVwfeoZj8Yl+lcGuS2PhihwAHrbUqTOHLvXuFgdBO7Y1Y6GKSTD4znTZhTVGpICs
ienC2/nc9g5q4XKc1wAh7VY8gZUzfjoWTrD3qJLK+t688LGw1cJRhcLpdrXbWFMX
zq+pkYvjCYAcYNv9iVeNv5kAGnRMtkz1aE6QbwuuBcC1iYX0M6qzx40DZcBCS56p
5RN1GghkgauuttxnGx/p5n575lmcejuMcEdZHBnfbYoPqUNZmaVYQ/VJJDGcYE2l
pCaeKPfqcmenhSEVGydA0v61K1MSrLhrHzfEHBdQtVrWWJqofxHM2Y+4v2OBO/xN
4bPaKtgUonICtVEADeC36sTMb5Is59mtEmRhaqeBdhAQYsPV5Klnpn0kyz7Ljm12
531hb74/NoawD8pOmYbcziIDG2eFw/T5uCXid4KRqqm+ho42p24ciqYt2BPcnGXB
sY++UEpOMnsTiFuAf8ho5SuNcfFhbfAKB3NnHG6DTR5fY6O/JyEAy52e3fjtRNn7
bEVQgF3sc1oQjXa4YpK/UyPR+esyWbx9r+bPBHvBITCbKuE2Mwx6gK9WqOVpy4AW
H237U1+Tz/Hg6ZNfNCUCnafRSH8DS7pCmMpWaaPmK3LuX5wObLqXL1Hjp37kPH9e
Bn3j+AovTmEYZNPl1Fm+WJd3ZHcZZz4Ff18PfGU7yfo/4Zj1W65vl4TGAO3kVW3z
uMRUYOC3LzztK1BmPhIOX1OkoTlqt6WztTS6SYYetu4Eyo+gB7OUD7XstH2DiPot
Qga9WxKrjf/C2sPSP7dt8JBNBET3V2D4jh7J14OYsp6FREAEoTggoK8CJbdG1c1Q
0RB24t0MuYxlCaPkjN97sLAg4JKOuO9kXFtXZjpR0Fj7AJrlmqnbfFLFes52ljrt
kGnMiHrdx263aT9N0OrgTTAqi7o9H2kTweMP+R3NQvHjv67CCvdqwjpmRyRQd9tf
vaOrhTwignsapt1c1QyZaUyauM1zjCTOlw3GBN62+jaOjbkcHXks3blO5+DfvNf0
fSkI4HRnnWCMQlB3nEqzrl7I/MKV6amJMQA7nzupU42xIVYEyRX+9vjiE+WdJ4o6
xljafY4jUVIGcPddVtDkWYlLo6UhS1wv9paQkx1bjEOVY+dS+B4oKZ9yaC8DdNYk
dS39mNd0or3wfQdNI3wvyuF1y/mr881yPBCkBZospFpmv/zLuAEkbU0czwTs8x0A
xXJEPtXMguDSAgAr6aAfMCOIRJbPM8NWGEXsBqqdLkuKsfJgztLg7QmNSdiD+ajf
0LAnU6Dznf3Qrw7MWqYKZH1ViFMBljO6FkY4XlAjBisrLzZw54iONn0jXaUecG8b
EW4wYCYIRHepEeoM5/+Z/Sg0YwRQ4EmORBSxJnAr2voVtNlZCFbS7jAvt+ZEkho/
K0tWp9XuBJZS+Y3swfvFw0rKBPwAPoX99p9/Hirg1jIrHmj1mk6I6e2+kxjq8Ptp
91s2T21eyXcgKWm1kpjyOblYJYdZnoACSxgc/gQuJVSpX5DEnVyTNHbTvQtgI2fE
oZpCtFiMEyl1rApO4nxnoK0vH9mypAj62vrvhabAMJUNMnX9URH7muVfhmNyiLaW
6/1OmxtRAFfXMqIV2nBlR6aG2DZMAJLgWJkAV2KdL2Ah2/I/GkudwLf7SDP0hhHd
wzPrgbacG+Y9zdobWoULU29zhwRFx+cGO2STTHH1QwA+f2BFPPiheCSsB+XuJ1AI
yx7fvjKAno6Rxw0FaxxWZgeNHdyyS5QnMg9MrNSpcc7WKM+FRH8AJWVqTeiiGiQw
bNFmh/Pqdxs6GpqTHGfCYAtPL7m3HJ+XLNSz/dmNXfPR0bsOE3iDSDnkJf81O0Ii
aGaCQysy0u9v68sHfpcNCDjH6JM0il62RgmjhY2BFrz246kV0vskMM/vC4HcnbjH
Y/JQiV/qfrsDLNTWRS2AqSvnZi5JI+9ZHBXkWiKDZYKW847humcNNrIAlu8hr5VV
USaBQ6g06XV505rfz1qhAfrJtvXKrr6jIt8OcO5scU1K5avRxTUJEtZJrs1Y7pOZ
XlpcE5T4vYBZhvlA+VyNv14x1UPdOktiVj3bcJhrgUXSR/N4VPlZyx6k+l96eGv/
lLq0zNBsYxuyFLkEigVuJfio00DJXZirTXcO2VFftDwHJ7xfjDjxJQU523l7WS8f
0bT9tQKbFJZfEtEYS/74jv9GgMeJuU8ATHLqkYhG4rGpAaXS3Lt2yQ80zOU1iqfq
n+iuBXv8TYGayNzySQFLtA2pW9tGRjL/MUGcZRsAbdDc3jy4FBRaQNgIWsHJV5H4
NkT+oS7ywLaOVrktsdh57kO2iYzkxR+CIEFLCTVQKm1YcjC4dx93IJWb5uoP2Udy
gPQcjI6ZyBiGoHXxzfPwVLA0+yATLenZG2cAPSSfN6Aw6HXWTIQlIC82KAdBdGIC
qj4d3hFNQvfeEnzt659pUL75TFD1hyIWFi+Azp+ITeZcBQnajaPHrjQuJKlOKRkT
1ItKFC84MYsMOIaKRHzHzG8yPerCJfkYA70zOIHL10bSa4iMZmN75fRAO9AjkiH3
l3w/Mtp4nQTP9XHUfTMOu0fP89sZY8B7yJHJZjOcFM1csKImR+J2rKCI5jpS1wiz
YjXrO8sF7tay/HelI4wq3WiANXgFDxTifIf5ql5l9w00OKe/fOLZRK5F8H3krCGd
p/fEmMDsA2QgFopVMqQ4HmXwbGCIjlWTf8YMB4BI7bsCd8gL50SKt/KUXNxhF5DP
QHxSDrnts8xWPNkHqs1Ideki7kQJ8Trk8q/967T1neu2FdKKYSAACuj2IQOZ2jxy
clK7uWnK6WNK/V1b8ll8F0eNBG1uRlPN2G75DObCl2QXhYKmVsyDTK+fP81V3eXX
0ggHBzOlzKOiWGyH8bZjGTSMh72D5U3UN6lk35DoDoOIxErJMjDdNRGMohTpYSAd
J4upaqvPLgKEgQwD8L0xIGnWu8U5JZ95DjcD/vopEE+9OhfkLE5Q0GtenS/jDhFB
gvH13c2EAxiJzvrFY36WtFjGfZl9lPcJ9zFJqTNO1/4N7HnZK9gO+OmQcVj+Pwz7
lzLwMaPjIhZBaQlBYNuh6jx05MQLtGKQjPdEVCKXSXFuzBf3xYO6mEiax3x3J4xT
wQTBD0JWZw6ClleX5b9ccE9ugevfgwgzgAbstfXQo1e3OE0W712Tg9vMtsOkxKwp
kXX9XTxUT3n7/l3HP4rrj0OOpOo1FO258JLs6UNurKzzachQDSg2VlNGQ37VzL3i
eaDsz2H+79RbrrWKuzdWNtSwaua2SYGAJEk67rqrCgQ7voCRSVmUVGamcYJs2GMi
lDMf432/d75ue5rsQdKAiUdWEZIDpW7XJfEgiJz4vimIR5iiKezCXIIInAKreLB/
490jW1SFi3AaXwpRHjq/GrErEs3FKYLSxyDx56cW4MRH52i04XQQSg1WX0f7Pupe
D6mB8GbleTDsA4BRa+DJS3wDq8heZ/FB6Vy6GcpejMGnXUXdv9lAnPpDiY/TLPn3
PvlsVad1OqaVsdVrnNEo+8uN529S1kJp29X5b5Lj2UUVh2VF5i4M1MkkQF+kR77S
NyPrk5mVpBCtDx6jn+eR1BCElD0WgithzJcaiUqAcn8UVX4k7b14dw+n1MqgdAkv
k88RomKT+DLQ2QEPnBqRw/k2BHVyLgchf8loS/TI6xp2SElfuyRXi4pII5ecuAoO
H4nK0bemLlq9vCFIUnPAp2lqYY4a+8OWsld3VAB7qQElsOA5yt6Bx5c5oFW9yPOX
AxKQN9eJ0WmFu3rWwxqNh+gkxc7vGgI5Gzhgr3X4SnDQSc1LtZJUisoUTy9A6z3W
kZg37k084vL0C+HYoDFh9veQLSZJHgSfrJV9P7653oQDJNyOQsySdlqtJVZ8ynlh
anLcoqvwNedqjmOxpqqqHgr7irXt7e+VtESyy60rOWwZvMzrp1x+ZA0if+WyyRlR
yH8JlyGLGTQ6dv2GXDdTmYcGhXALd+ZWOE9dfLGjzvs/sD+G2zck5ftOb8Qg0jAm
KMmMetMbpAxjGBehwerRt8BuGq5xWr6Ap8N47BLfS1Bmy92X7k+Vo1TqR/RhQzeI
WUgAj/a2B9abh4bJyeVe/kjrpr1GNpvcCaqrbZqzQbeYFpqile7rKcRCW6IhGJYs
bs3PnRRVpTuTL3qtDZZeXuBYfSrQjSyB+f8LplwtGpkovyXHo/7gqOzrzS4RReeX
9y5ESJGG+madUryjGrU3SJmFyZ0fCZBepb0yWwuAcPWnZGxO24bkoAfdSa7GZzRL
u5mdMynK0dkMcaIDV1Bmfy9cKVRBM+/JzX7YSRtJeCxRiPspzrI84Ir6yuLlvXHW
o12+sX6ofc6eB652zw3Mar+IlTnwMeAHdjA/5Swj2YJHpfV4rijOC1cJTC/oKqk/
GoqFj2j5YKGamIMjbJlbYoFZVi6ub+QDgwLoHMtnuCDdJGJBb6DY7+LZsC683s9c
ckktSdjEa57pIo3uwwk5ZhbD/s9apOf2bWCZXgRE3miq+Fgdxhdj4f7flhTYhA3D
QeedIf3W0cHxA8obxGvu9inTBf/yyg8ieuitP/6ti+OR64DsiIwYb1q3wqkLl7gt
Bluvy15pBd3Op/zA+D0AB7q+6nVijaQ2sQ6bzypHEdSquXUIas9gocUH+vygFp0f
Tzufh+doUP/b8CV0m8bRehFxLb/c86VK8p3kfiymiing1Vfh+F5uTTWtmJ5Hh8vZ
Oaa1GVJBaxnXGKJP3oGpudNQenhM5zJd1B+LF1cc2y1LsCXsvoXvDHf1s0an2kbB
Nv80oq4sMswysgJFT0y2Wojrp62QdIeqWFS3amBAuGrkqPnQb1okWYQkQNoR6Wrb
VkpTTcuaP6a8Twb3Oz1fbVsoFlI3t7rrglK0fvfI+yYpb4WXMJJvh457eRpA/sEN
/FPH8M6H6kXgjLZdgUfsZuzne8eP2frYJU6h2CiD4B9rpY2Ngt2WQADXtv234zvZ
QhkhfYvr6Ast/+9FtMkX+FT4l6y+t9OrpxZAOFn1DqrqQite3wrYyxTza3z0dZkX
UE0impHGvZ1/RzSM65fxErqpuUyvfoqPyKJFHD6PUj2frnIPv69MAWa5Pl6Adf9u
+MbugnsAhuk5/LTB/cd907fDM9uFPEsSMDIk6sDP+VGRfIaFF7VVd9EJcSFEE0+w
5W8SJxQ51GuqXZ5SVmmR+oGdA6NhFIKM9nqTU2Ssli/z+Aut3fcpYAV/k+iPiQAG
Qme/NugzUXacxhdA/HXwG/U8/eKRqTFHkzIHkyRDhfd9m94UAXRHduSl8m3cXhyp
Ez7zERcHHMvEBcV+8gj3NeInYuRHxxWitFI02qEdNvJSoNNvfKkZLlcTW5UAxpLQ
xeZAsIOaO1sz0O5xOLmiJSEBCC0hiZN8omMMCEPsXpFWvbH5oivd8LQhNMmvwoA5
weiq9lJy1FCYBNaeTebQBAQEBq2es0l0iEcxrbhZYGI7O7C+Zu71laBLrxFtu3lB
F2tWwgJB+CpI32zNbEXXDFfImmO14OVtlxaoiruT4Jd2+N3Ah1V2o2id9fCHkI/7
Q9RVbqU9+LfPe8mz1iecyg7Mu9Dx77u6gvcQo4XtAsVxND+A4ADvFpW1NEfLfz8P
DFEMKFG/S/k60dZX33k36bctW6BI1Ps2uEko7QECitK3LSHeXmBLIlY8I9T8NLwt
g3MKGT4MOJiVnej2grilDWW9rLlIcgx+srk4Kpf5AEF4Pr+5kc7XTsvbUulKkJb9
EUcUqfnPglySpUd3aYpYgA/b+xgCQ6HI2FCUKQay4Xfa0Qs9VcJyMVl7ibv2mB38
8okCSQfiDTln1RJQQUQr+4i2y7Qh570SGaITx2Sfglkg/A9LtOwh4yNb6bpB6yLo
jhSe7svn3NYwhDXwDdyBp8B6tDpS+czWJxYtkFe4TylnGP09UxSmyhi0PI7/I+4B
aJD7smWxayWnSmP6pqEHagTjN0X+QNxpETxckPTnba4iThO/ATRr9DuBz186ZsWC
3soaqLLI07267b+YIGhrp1h02UqNPjTRRr7tnkK+QE4MpizxwVMq34AM+3zUZj9T
85Jd8Azjmcd84qB9KjRbG1ZjyY4xqUGMBybCp5fF9DPDKOLUV21qSvcN+uDdgHlM
i9ktN6cQUCxb/GAxcck22bsRZOuLfIZ99wRFAIqWGcMDdg78BRqcvOHkoKgnsWRG
NAYLSh3lUXhnSv1sMqYWuvE5OraSYSpqkD1a/IUBn6o9gNyGQnCyRzedAhIns7JB
yGelVztVzXjSecn/jJda5VlTjN4mZsr40RZ8PFUoYmiKarkjcaYYCqmB2SFzKkzq
w5//KaHUURYzQ4iQoc8ZohnRf2V9js0MHvQTA2I4jfz2aEXug8GXlB4b4zObgT8N
D63Kkdj/pvO+/S85hLDI/CekQt9avdkHE4Is5Wy0do7KJqxLfK40zSdBlKZf6no2
pK17OAt70NHpNIHLEsd/maWw6bQcr8WK9PeQ0rD9FKvrZ/tM0b03AnAXwDU94f6d
61DqzQeW9C1OZR88cruXtkvxmk88816yEnJWkQw2qhrLekCwFfGr369nXNKKQGN+
A3xsmPuYIN6py13qI6ONsDlPLLm/lX2XtYG/7QK510brUM6VciCsnTDUfqJUDq6y
Iz7QlZTExPHtUupL4tITmxWuOSFLpcNCI8TIZpKsZsqKU/n4fRg5ojQKhkJ8px9M
ON2a9jf7MWBFyn+cyvI4+w8ZSkIq2lPzJ3+HBr9KBUsy9PuRuCZRuRr1XmKRkHkv
qd61wawVL96zrduU01PNSzA1uw25eksJjj5WV8unxahilfDKvP5b53FFy3bNblLn
JEwuJ2/9RS9EkY7kbE7tidJnf4F1EgHpJA1hY0wgtdhfU0NpFUpRyK3lEm8y+r83
LYjASMPgjKv4yxYm2uNOczOjKbWltJp4yP5dodT81fMpPDQ68KNbSy1IdI7d2G9W
IP/xT2H7/+py3S+H8sBS0ZngxWkZD9lGcEgYMN2l/dgHHOGWhq1vMSWr1em/X6Tm
fiUVBlYUMjBg2AheraUa5SK2v81QOVXf/AqZ2O/mdjLupBz3+nRS4Ow6pmEgFHTX
HZYSO0Uu7LGOKS6/F07/fgf2NMTsXTdhY9NCOaGF7atTaoPbLf1PdNxCKonOTdiP
GXWRiQsvN+c3di3yHpIJZ1oqiqIwKlT+iWiY3BVihTAVwCmIdd4KeOkCZfugRcOV
JcWzfrT+NhBzgI2CJlgqioYZ+ZcBT5Cm9OHQ1SNWEFlVyFEcfvgTxb0AoLz7jfUa
lP0LXE6iYQ3ax+FV6u0U49v4otVq/dCM4BWZwZkyGor01Zn4CXGlrCM6REzoV7+I
C3JUhAkxe8PU18ssQ4Ihw9j/D6++EL5EhlPK8hTR7s5LOMGVCKli6hywYMQs9D7v
7YEzXVu2ThgyDUCuDDeuph747H+7RPrGsn8+SHVuLlH/7voCuf4sNUbjlrj3840g
5S5ZWbGsrSP867HPTLxUmQCtRFOpYOeVn3XE66ZD52t2fq3lXKAUVTEv+OQHT4fv
c64D0DM0K256oMRp3Nqfgh3izhXp/X8MNv9Goa3C3BXLxOtFKIz9RtMEbm5H6DHR
wZG4iZSCd/u6/LEeEfk+B8d+iR2MUkuDB3RWSKVX60u6m5O/ospRIvom6shNg2Pd
4JN0m4IQSuhCw8x0FKYIJPRrDczFsdRt4UbKtHtcxA6W/gUf7wuFRr9FwLHFX5eH
rBzWkaJulwVCDY/x75FplhvZDR6zFpLGooYIjMfZnrjaLb5bo4JjHVc2YHlByYlz
AgD0CdfcqTyTLnK7gw5zkLjtRZdmC1iB/P0Ga73o1yZw3YbIQnmxV4e1tcjObSos
C3QnngBML3pLDu0KpkIRfTbfCp8aHAg0+ce95Fgag8wv659+gVxCWWPMeoB8BKVe
y36oLgvxHLiYzCu/9LRJBQQ+Rtuf8F1Owu5cec4lcOBdMhRe0Bm1eHnsDY+Avxyk
iSwRDIBVDP1t2HzrKdgadRexz7NhcjGllBC4+XuBdZin+ZJfg2EcPKcLOh3QvZC1
IFBAQFeW0bokS7b8jvcqk40Xh5Z/DFSIc9QEelvU+pKxqikWOp2LShCRiks2bk0f
hQvN4Wbjd23+NKgkxtqUbXtIl68GiQLSoDU5BJBicWN/ctPw/g5bQ33KXSOflj2F
Lbb07nVJB724gtVy02MnYOAQbowbF4vPAJ/xNMbqo2E=
//pragma protect end_data_block
//pragma protect digest_block
ldqB93mJGpNzGOfmbU1D+Q2OHPU=
//pragma protect end_digest_block
//pragma protect end_protected
