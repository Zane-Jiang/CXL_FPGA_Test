// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wqZUxqh4eRMJbp8hkzCA0pPCmGiZwiL2ipA6PCh/UzVgROJT0nzfPgI1jG3+aCJW
2m/0k9aOftw/PAMZQTz3AOFf/MlQbTS7DtvWGt8QBGnOHtheUaT+9ZiBXO21Fham
XWGNYwoawlEFbmqOm3y+eitiNCggbQCaupw4lCWG5uwBvT1SXhUayQ==
//pragma protect end_key_block
//pragma protect digest_block
JjIBRlA3PyBEhM6Tg8JUOJs54FE=
//pragma protect end_digest_block
//pragma protect data_block
7JBftB5NnCgOVhaorOheZqu/kw+nvSuWKIGSDyQ+O3OG9X4H+eqBwUtDchDH7lTx
a54FTWQOSK3O+jmYvd0dN+Xqfo2/Et2q0CP32lz91cahVJj1l8pzTXDi08O0SZys
ccGnaUTFNg5zdUKe0ccWJHM5paXWKvx1WN1yxAonQJbqbfquToQvehFTJxGYeX+w
q+6ZVl9agskTaMN/uCCVO+EMEXZE3RxiTYUQVrtqgAcZ3q8+Po6xZknTII7+wOsu
HQr24Te/k8EdWcQmcPibBKiFMfcfuCubusQ6B0PlMhP+CVN1mnYfph7VAMOIeLin
j04boaQdhXuFyR96sbZANvidS2jTIijZL4GbxechteNVWfs10d1B6ACe3lH2nK1D
ZB6HORJpTCT09dln9wctG9gmnzknKIy9barAtTuGLponkEedaRciq1/5zeu0TFKB
lgEymUmCl1blYSmbLKy2z0GUjW00nx9rtMLJWfJYguTr6/4SRXpuWWeFbvIgEF8t
7nSYrfpOF0SNHQGQt+x8dKTf5RZSEkQjSnn8cbs2Xh1LwyBNX1qZXuWYekP5b4d/
N3dExMDITrYf7uU+S+8P3DVcc8eL2SX78PMQTog3keCd+S2hNCxSUM0W2JlY/iOl
Md5YnIsOvZVpNfX5+XWqYxCoswc3MXxPT272vqTLKY3YUPK9EFpY6sJlFeF7Sxqh
vYfJqi8I0bsswPvzLUaux0VgMJkh1BCWU6m/TOWpYS/4L6AxcxzYLjCBRsAA6JJT
zTmgUSYv37uDNrNs1vbhUmicnzsmrm114Iljwnbx3V8W4cyt+Caejm57ZWK8GHvA
KnM8A0bRv8CoFWz1QDg+VDNw8VKyid/vHG/4Ep60iTXeXNTHrlSUL1JzvQrOQJCp
t25vOghHs0iz/EPYgVj5FblIYQOlbUcSDJYmsy6Mf74J3MFqAcn9hmEeyZzynzcu
GgrqCjGNEpoXa9flh1/M1BJ3FTq+m1qkndwXdz/ABDdTcPZjUZrhIlGm1pmDQJsF
C/XWXvh9HFNxg3Q54GXSOGDztTVwB9yGOwrSflDE8WnGicw7G7d6T4QRmow+id9r
OJySc2Ih5V4EZq07ZsdsieeHGHaSafb7njhAhmliHtcQ4osCO8NU73VHkrn6qp9R
BGWJ3OnWpnwyQSkkU0flX/y4ziNSDvIhrCxh55AyLE8xgUh8JvOguDAqxy/+gkz4
YpH5UxLtTzDGRqc3K5pj0KRAFZCDkZDNj8LsHUqA6JvYiqiv287M9DfCr8y7v5oM
9tgGvaVRQRdwoB8wjNzfVshhRI23XSSmfghJ/bxUXLxsqijS7naYqt8mLwB7fnTF
NZ7oHPGqygf9Sb8hLT40SGFNeFMI7w6qwmxC+WAQeMevbccd7zMjq4GSJKGF6QD4
z9f70FuQ8bPXB9tIvVqFOT+EqVT8QgdDUtQ6sCInh4bt69ByC2zxA/jTa+lktyPl
mqPnUvhB96gS/paYRjr3k+wUifqZJM2sFSUeNo2vikupaSzYJYBYxq/AhceQNxGs
zV+ZxLleR3IR28L6iecFX0FFAAR3TYnejKB3UmCFWGpvuHxWuUmXyY1pM3VLJVo9
9N0hsWdE0VpOe4oDqwhk8vBKD4R8xPWmRCqsuh/Uy/edab4ufSVeiuXcTVAsd6TM
G+XfHaISfgeDqJ8xTLwTDHSoZ5zbch/Zp9GIO0oZ9d4t2CyXjZG2dLj6RTw0wdeu
7pk6rgecTJqz7mW7iKXbnuxNbqoxMYeFmZrEKW+XcN3VEgBTnFN2hZow9ff0EF60
kep+oE2rYAayW6EqL+JD13/dumX5YmOwyR9rm6Ewqs+vWJnspVdvzvk0S13n5E48
m39CWouZUGmdrxEk9ym6kZoK1oOXFIPvH8SVAVPy3/eGaPCukeIm7npoaVX8paRg
5Fu8GrOBrCNLl3N3MMmXL2aDvZeILRa1Jwg0QIFLgHmcLZsVKZftty3mlUNqIsnR
JA6mg37Uq7cGJnNrB37xaM0nkdjDRhReLzDPsXhTZOTUEvaZu5PO2w3V+28XZMtn
vtqwLe9q+6D7lvzLV6zj4cwFBjlp4PBHbfcg3tbXrBDcPVMNacOXy7Qi6BkJ1Oy8
qY8j25prZeFvbs0pjdK96687IWlQ/m3+V5qcyRis7jFdgfK2J0IRnu+XUtQrJtSQ
x9YNNcHNpllSPPoI03hdQpst4nkUP2P1lTOhtmJgvKd2xJfOi3CuftNSguTKJTyN
Tda9PGqdOr6BRev4Hv9Wj0ZZBjzpcvCFAXGagrPddDtA6zfJAZ/ifM7USF0ZGWgc
49dwmMmvhc+9eA2SfHIYTAbloRwgklGDbbJEbFB6lTCHDCRd/TghpR1E7x99HOVe
kpAFVnDYaQiTcY4jyQATbdy7la3If9Kq2VIoIyGq7VOE2MEq+c1g2+M58rPVS9Gk
cMiu4QsC1EAzqoncuIOPbeS1IUzCPatsOstZ58eQtSbu+HwUWQ+37L3vZsx0PMlA
Ci+xi2LQDZgsA67mXm5RskUoTQ/p5jzGN/BkAYDTu6NOrILa2fsAYHHW2+PzGnj7
DDGwWyNN1dDCZMgHeDGgBnw4t80erm956Wo8kAWlzjoX8xKxgkevOBoZfXJg+JHP
ZckI5NNwQPdCg4nvQmntjj02fa3GhaA+7U8FE1H6kwVUmAY7dBjEcgY/FMgmnF8O
NGTzDwTjIMZMu1gJdR3fkYV14WmAKZJ6yuRDa7lfPZM6S1e0B84v0t4YrctkZlNu
nRqiniGJtfaR0xBbX3rXll9WgGZcj8hejP/8PWsSi5hgpq95kOsgJdl0A9NSUJeF
PwQUDjPZhOH7ywFnlmLhPQYwUpxzBY8WvDRXvlO4hyLzhqLoMBn5r5GIeH98QCem
r5xH0eVUzLmn5WhNHiLxEEyzFcuS/DkY/LwLIkyvtleGZj8LSKUbVsS500GjYPGY
pSWu9E1j9AI9NgaIvZZMwY40af1jO3LYQvfpw+eRBUOxD1hlmdOuPgdJ3eYmW0d+
2zIaQG31GmtcZRujQ7vEtkC46xcK433FRMgT9y+DL+PLl5jZ6LidRRbWYS4SFMU7
CNyn/Y05FM4tgmPuiFE2gPKQ/ikmitlxgohV5u4Th0yQfkxucWaMuItS65tZIpyC
vfVW6pup29FTZMpI0frt+5zWlS7eiJ84kpy5eJtOlsEjVjrEmsNcH9OhEm7Fp9qX
jKfAsGM3Toh9ZPTFOo144zPMc1cuWAwbYgkbLtW2782ifxFUszROSE4Z7i6Xe8C1
XDyEIPIeP3kjsC+ULLAhbw/HtICQHuT3yEf1uDiPMvShTiqFtfe467RTIMdMp9yX
vsCf7VdYdVdiyMYDKudwNzsYYbM7uRYPosAAXue8f23+IbIRMqEyrR+vNFq5n8P5
7EQVgMMmxDwNiZxLZvHiJ1maVNxgj7QlC2xGvFqGuPEHBxhy22qWI6RzCI53oC0h
WE5Q6u2ThEmSeGVd1tDcUKnZjiypL9yxpCADMBKOD7Ph6kHMIcfjXOyY4c4QOorh
Ba73Ek2P60N9ZJ2c43dcu9/LWzXdhkDNBRLy5RT6q5qcz2X3934ehrvdGWtEpLvK
L/NDJPE76hfIWCzvsgd9C0nvkJSJ8AYxXww4Rutx2VldQ89J3trBU6atPahV0aNn
xwLMLH+FcZZukoMMI5pEYDllGX5ZCh19bt4RYE9SDVPdq24DhVK2jqTYKbcRGmPq
esW5BwczVLsrAHwkUGMzr0KIcK2QeDEjMObXJZIS9ggi+vDQLN9TfyaQIgAubtnH
gM/DCq4irtUbQ3MstsaktF5rTgu1Fz97JeDAutK0aDJ2FF6quA0M7Dyy19zikXq/
cD4+/pxngd+4/RFSgupO0+SbOFmqT8YGB7uPvZ3OAs9ki8l7R5A/VJNVKp7X4Sl1
kmY2e7aR9MwhDfcVJrL8FKvSkP0KoRw5cK49ICKGai4FRQdNy0ljj/paYGpiHETp
2mYnqgpUG3men7docr2YhtCXHo2RYuli8ygMxApUZ8I9gbfj3qtcKHLIZojDTLjR
6ERSJyubZP7wr79PUuxLubNfD0c6kRqBDdlE3ujJujfm1+UAmxzmAFlCACQ3ViG3
p/IG+x9tDwCd0Py/jmgFtdqThNKviLgJn6ybS5u6RDzFDgTmEHjD8wMv0JR8c6MT
P3xs64eDBgp/D2Z98VRNdDOUPZMJiVGT5ReDzcq6LIWJWMkcULhVWHRtH6rgjY+V
DQ3SjOkVcSduuA5/sw/ONBgci24haqLTlQ1tTwaggJ9xJkgprnvNrBptjEZQW7cn
9eb+fgQtVt0U+DwtkCNgr4Y0fnWgaLG+jzSLiP1v1CxRFfCi3zYxzORDj+zmlDpV
3qXYBU04dBnrgufBdNr5MTItMux9avql/KlEbzZiFZTYfXLaSzgCi7dEpPjGvaHh
uyqe7hgplHkp5pv8Kg1oPw4a0uf1rdTRpES9XAvHOrFQh/6aCDjXlBSOzXANerNc
I1AM7bgjFhvTnVA9umBlsN/AwmWM+mXWYWB8fjm6EZXE3hZ0JgzRuRM1xjCbBTMT
Bsg6u2LR/FkrKvrIaeOWdB/0OM23VzLGQWLufwgpTKmCB4suc94uWcJzbfEripLN
ohw1qQQxutoJVwY8wxFx8Shx94XP9CquiyZoIO2Qpvhe0+s4UdKOA1gY5sM/argX
033ni4QhtqFJ0eJL1E1kPh/GAy54/o6iODHWqKH9wiqmcULDU+ryqtBQz73S79jJ
8ZJ8pngcnOkZ3Pk36XMjQed8VwQJdO5ShvcGOsbPeCKPBfc7qr85uFHL2l1yvy73
vgMJuV8HkFvX5ck1YlUeDo/NDvkaje7/q+/wZPlWwMyGddpnIvVLq3KNuOgTwsVL
GU6GHq/Uh/YLwczw5Z8IKs7SJH0BZfyHS2H0ax86adqjhHr1sqmRxRm18pHv1tUU
dqY/xew/EbFYcD4sRzGnaKYg5mvY2jtyqPBLva8y7SHq8Kcbkh2BlEI30dPpOrwj
gqnUIFmfsLSFiApAWWZHZDrNnzcgXnOcv0qQ3ErpHdeAxdh8kJdRdle1oE+1z0+m
pHpD2jrJ+1B1aTAnh89Esmkqr/rUGi9ctPcRJi8z3h7ktPDWMlC+yXkKe1n1B3Gs
jepm8ftt2F8Gsy5FxFrI8HDD6evROgwpDIGEnEzd/qsgg6UWoKaPDfLY1CaDRdac
tXCS471AtjKYBebOfCZczXbq1bGAzXj3kNf1A5ONk7MfwrsNJOIV5gPAKMBQTqtp
J6u2Z881xXRUOrYMzK6uzDM+pLQvzkYXGTMAiuUXKs/pCqfC8+/iSKOR/sJ6QcbG
3VUxEFGRlJmg9gOfuEE7r1cXfI21askaUYIqdJ3l1jAwArfIvP/KAtBHfab7svLA
C1M2HfSvOe7LHbHQKYJQ1MWii/v45fK/0IqiE3XL2lRBAjrhKKgGgqkZkFE43cOb
87tTwBx8jAC845Xryln1Vnp8i7nJwCFsjeiMexfZGEueZudMWqoGqGLOVMH4806K
l4wYmXWWXvc/chbaICdV2tvRUZc3Xs1jN5hBc5epjL/8aND4prgXU2yJu2sTMXMU
80z+5P8IOFnwORrdhUHzkkPyY4YPr0jR5kRTWE6ctT+cgBdywDJnbW9a/gboNl+E
vORF0Ba7SGtROizUHboA6g==
//pragma protect end_data_block
//pragma protect digest_block
g2uTGfDFq+lXh2G2hrMzNzTpheo=
//pragma protect end_digest_block
//pragma protect end_protected
