`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
M9iQ9RmWN/ocwoShxqdmsmiRyYz1togyrizJY/zroFZPmxZmlFhNAWXt7YDR9p7i
SEAJzFlHjkKP11NAw8KPLOcbQl9uf1VfNI0cxFLt5aNIfZ6G8zoZ2DcBZ59Sr3V+
cJtCONltMJYEcEm8HrIOZep51SQWm/Agen4L4fqvjvc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 9696), data_block
xfF2xeKOYYIRPrBGHP2EKOR/f/KYT6vxiXiqLi+a7tDtleyetClKaLb/BYf3ShGG
j7NXuzO3aqmg5M47WNw9WfmwV4JTuI6RCio+3OZUT07K0GC2cbpQ8pkMOFk6qulp
GyqIvAccuuehzxjVlKBu1kf+QeTs2MR4GQ/hMDX0kQiOFyN5hYfznjl3hwQPIbuT
L/netaqswsLopeMHnmejh5/79VeJpM8J+zPYMIXynNQDyhknjJZBhdg+KyEvWi4B
v3sr9pAs6x867Zw6o3fFHarKyiUmzpBusU4lwSwi0Ov5inD7CII7ctAP3oB14IBX
+lwND1RaygHuWyLyG8yJxaD9P/3IyOqF1ZMP/dAaiu19YJjFvvVvao8YJkPziNwg
Kx5vT4TTYPxvdLLSHRyZ14QE1/y1aJzcqBN+/6gGXmj/jTmqW36os9qpoNPGi2ge
kfnkT2G1mx4VpbGXDZxMvzDW5a4XiuJ5gxH3ElmdXmTSGUJ8qXYiUbSqHfOj0qhw
1XVts9yT/HCoZRjrux+8jb5ndtQeauNCdUq1eFLme2AS1iBdOg1h9H1DomHDD6WW
K9764OOVkgWwaxxfaJi7DVguWnt4SiExqufyimPq+z1kp66IXU9EkF9hNmG8KK/G
H/5ByphTE5scVLZglmsqE6l0gJaAYBBsHSpgMT7CO5VbivNKA9qhmpJCamvLX1S/
yvp0USvC9AqCI66X0X4amwlEctPdizRM3NyBPMTjNPoR4/YzWFDQ7aWWKIpDFT9G
eDfbKvTRGiwzYpS71DQ6dIzeh5re/pl9YLUn1j4V5AkzZQSQYtJi/STljtexH1RA
Fk4V7x0QU0tWbI2AJxvMT4C6K5vDvFUh7mlVirqfJ6UrMkeAlvtBFMQAJI1vnOFg
fr1I1/zeD3HvKNRgo1JyDSJkz6rupu5oLslBU76yNWRjIDi7K6gko+/xAcwl4z+f
osz7nRY5q5CirSoChHH4/E8QdqoHdgxAyFH/80cazEGpWX8dJQfr9TX9C5i5ti+4
setlctuWcEKtdd/DpHFyagfn6kd9b2y+Oig31vVtu8tGAMTMzW59y5qQYe1EbTjV
OB78rBr4870/XgtfIhHbAoMycLyJYYOhw41ihI5VXTVo4E8hIvB4HSXAv91gsH7p
TGmVZyxOhm9LitYL/svToSx8Pk/5UbGjWB9NEd8XbFVN6Sa94bKHBTY3DxF9iSUw
QF/nJUrsedxoLljTU3ltyRqaJZexlCqG3s7x+jzC9ny1zaWbcmwI2SbduA19v0w5
st0Vp/zYPMVu5z7jofD4PjuX8DIiHsTFk9WZF5xlF7HgxHqEbus8c/Gd30Y+QUE7
p1+4MFol/QLxL4xrrOExcxdODo59S4xjc4QiABWLFarLNApuJmYpv86l5CmV4Z66
23Z2Sg9viAUNDYZBt8cin0x5Pavbw3nTFMBqNgknVmgdK2eTsqzE3vLEy+RoxAgF
vv5cyVPZI0Vu0h0M2QIzMIiJTv60l8jmBy8gVQscX7r9M5jd6ZC8enwlP71xQkaa
OFeNyfUoohIX+no8w5CkTtvM3W4EhR9qvfVVImCMGvm8wpxAub+b6T19Ha1gDZc2
1vEc1s6Mz6l1UDVMj2eR0NH+oRCNeyoWXlATLtGeYtgae0Q9nJS1XTsLW7gY5Rr9
KzBsqQ/1JR4wYtvzH+5rTU3NQxEE6vC1XC4BEiaOuEDComGa4johjm4XImVKADCE
i4GsMyaaVrn+z1expm//CYkPTtX6u+TtOAZy2f7yscf98C9pDz7uS2xkqkJUOdIl
ZVThDQo+0GlOEF9Eh+pKTxB9K9/4Tab96clINoDpYV0N01Z7obkRqkd5FiGEYqiz
Gly1sNeJhbQGfLtA8uDvHbgOSvxZ1vG7/TRL0KXb3+EwMT0XZfYaRQZFyKoSqk64
K1K6a0NJVM7R7H8YWbS+HUVaSiuUewibRgTGqroSEyJ6uS6YrsZU11k388XV9inB
5/oGTKe2VTyo+hYfHHxqCzZg9t82T2nyhaV45MAoAMuzVwd0u49WL3ESrCh/vcGS
SmcvNIIm7IJga/zbaDRqpqroq3ryZ2VpL91nCzITBB5BSa2TkrwIaDTRfUKevUC8
oryoCRMlVB2C288dRrY824qM9RcLRe6JmDKIaP4k/1CY9Cs6DmZiqWIbVRnld3Ch
EKnldPGFQtSRPkBUOJeJPhbA2/o1cP7Fo8dc4778N0Jxi/i2Ke/+DS6v4zbEKwNc
cdT5ADLvvcKD2i33qd0jHQrmjAuGvYrrdSSVDCFV/oKS0O4BRqaT3M/3dgM9u7Ia
gq0XImOdY2NDkbUyilsF4aWyBzTtZXxE+4BLsoUhjQoJg3mvGq5IECQdGZ+mMh34
GL6LgucUOA46DBJPjyekKrENAdZC1FFult/4BuLJKL2fGineOFMQLde7fqiWa1o6
ypEhfy253c4zNL7+oRy5OWmmDBryEL1QPw55rSGrpesJgGjIOYvsEq+4U0Fr0rcY
qRsyxyocUwyVFV7vxchnL5OHt8OT+JF1mZte6cuV8tIJ5RNoR2TyZc9Kv66FO4m7
olm+zQdetjR3AtJk236PwEHPDBeFJOX3DEmR5dHnSfl3rbXwAyi/vOZo5H9IXrw9
p2ElyPUr2xdADkpCihX01nER/siObW9rWuG6DL3eYM8rYgOKZ2TXo8vWctUQOL1Z
2vybfKxFGe91kqBAStWBczzswYHQMzE4q3RTG1kdpeRSMbLwGQG8wflEdv8msxkB
0urpzdZmfPyvoof4ijZaisX0gwRDoAIl8F22OQ6ZembwMN9whscSl5QIZ2p+j1ci
EvrKEfVqrDQBUzW5Ft2RWIdpknhkcSgssBUmyOtTqwKaUT7lPYliWforDAqFnVuz
xUJoxqlJ++zwMsp9U2CvHEv8TX9T/Kd5Mj74wR9nyzvCba/Zm+Mt88luFQkNCV3M
SuLp3B8eF8SAyOljW0Ww2rEAR/+kS/AVpcuf9YMnRZh1o693VTThstten7WVfJ9W
ElTPCyd36I4eClePdzdoBi7QFy5G4IkADsCxp0LREGuYXfo9Oh8AXkSIbTcrYRZp
Ui1DtBYV3NNQLmlI4lnPK+AQZRrJ2d9fCQxc0PF/anCB1WnYkf1BDk57YEjvONlt
TlHxquHMSAbyIjHtTP2vJMtcAyHOVRI8s46FuKdQuvE4Q8WWl7YKNuNpOU1GGUVR
yfjR3Z5fTKgnYShpK/HdTvN6kRdK7v/yF6nuWjYGazipS6ZHJWwPWWcTkB3nXk6m
DRvMLBY410veuy+wTrKD4f955/r+UEbsVNBD+B60FwF+e38TXNcePxu0Ah0PazDg
kUmv6tcErAYhufff2gDsS4ag1s6x7KkQUz4xn5tNKbKLvEw82Sz8sUgHZ6xWnT3T
88KR0u1jxksYnl/7ZvTwX3DYJKgm39g3wsG280XaRG/iBtn6zRnYfs2ubBaB2W9e
a2CrQ8Qjq/2IelaByux/VO1EVFDBjurNzouj1eCbUn6+t14wPjeBAsDwVVTsuAVK
C8AbaB6KGaOy1rgPmXw/8Cb7/gj9UGqbrBUm5jGKT5V1izxoH6DgBLnx4GSoRkhd
JzrYdZS8G0agV0oHibweqoJyNdr9aDXx45bMT2nCnNwvijYSUpjHhIQauf4+CEO8
ZWdkdjTSiBEzDPahXoHTWbTM9qUepBLySurJrA+CEWKDO8Lbfn2KB7gD1W0Tofg6
PSJyrS/FrM24AIm/4Ao4IzoO6nTg/hqjZdAE4oDa7aNap4wuyTDx4z8ljJHr5QJQ
rxCdEHCv6KTLEtbrjf4edbNe7KXdVgB8xavA6W1f3cJsHsFCMJhNYejR1SHHQKIt
G0zU+WgHQAhw44Ych9q2JF9LZA62V2UhvgBi90XoCvYMuKfs7oNPP9Iu8hrPS8bV
Semt0bi/STGfGWfwCNZ1PL8JhrCMTdfNhh7V18E9GDdbw4Ju8jDKDxStLCvZQ7Vq
VMA8oUUz8qDTzsK5ZckYGZTl4BOPpKIZr80KV6p4idk6pXPz9HtQOHCQVaqaJCS5
AHoVfXiueokAxP8B/6oYKN8KZueYn0zJRGUtpM9Wofwtk0BQhEZuVCCQMyIMfnIR
Rvp0Agd5yOXWSdtV7O1FCFLitxV5EK4KDRGKy3UYt5p6/VYb/r3Iq17RwEsGOurB
UUOFC5jSHOjGLenc2Q3iBajbt8cXbaRlw3yhwTi2rmr4I3v/VvodPSEizrZfPmpb
QKmC/mPDI/usznkCRVdzwievJ4rVzoIgJmbagWWpM/ARPJyEowqnrInYM2KT5maJ
nbTteHxDso3Cs2N7Xo+kBP0NQt12oikxeGp0r05tZy3VuWXCBhX7ZISYiqTm8MpH
sorazQHEHrvKwn13EaKxbqRmmp7tAcIXQXx/MBVSeJUA7iYEV9y2KrWBsAS6SaMS
QnaOMt4FZTJ1eey1uHD5pvmC/QqRuvVlD4EIHTP1pXRt2BUXR+ne94vPzhtIeAnf
DeSMrRqbuEbwI/gHKCqqtyvIyRDPP/6/49aew8gP1kROAPPmO9aLHu+jr5IZbWi0
JigXh5myx1OSjDm8MsQx3MxOY7QOIntbD2uIBl4SeUHPxeNnR4s0Vkeg7dakp5Qx
AeRvWjnevv6sakf/3MhHdMv6chlHf3QvAgUChh05jUXmrHEZn8tswc6MuOfwNG9u
H13optIBFGb/pRDY18hfLC3gSJPWbnIASpesaV9NVppDDwJ/ArEpLSfoVIUhnetk
ittBfjcaxCWCjKBbrjBt8rHKKG7taFcUR0s9hdV9pbK2ozI3Si71M6x6cYcT/WFH
AhzZvDT4EcQ3qe66ru3Omcg7FufPlieRuHN12HeAXwpWXaDSrVNf8fpdRgZKqQ4W
6+DyXRvB1l1Sz39IqraWEaVXwLl1UkgZn3UShvVHVMvWk4L9qn7oxmTbYjp+QkSj
t2LkGTVe6UnI0ZorWySoFV+JeVq653aRE+JRrxMDCbsuJIBrk7cwevrKFI4nWl5p
wXCccNqFhtdRWi/V7izIiPez/xpTGMnhOFeL1UBjlFoy+YWtWO3HBPw6peBPQA8I
lX1K1WN5pU8wWx1gpiyXKhbDS5N3/xwdFSALbP2HX0sPaQkN3GFYk38fzbMapzJO
YhDqFoVzMvNoa2OVjMOYzeZyBRxfdlPKV/QubOvphXknhkfuFfRkY7Wi7yOm+4cx
v+boWSbTMd4Ux3silQEbI0ATTJdSNVpnaBiRdOQvTTLcF47ok6wdIxwwIIYKC5zj
zexZC+E0KC+YOAe7wj+YE+rtfyNHo0YmANKxhxgto/88fqOCSS8N1DZin+wa0tOO
DYUB0ap5+BIcUoDjVaRFGrv9n2BUl6/AW6GzWwE6d3go8ZddplIjDK2MuAFSRtXz
kYJYca+S2RR9Fyc9smDdosqF9zcUk6/tbsOzc1Seo89xWM+NnlKIIuDIcufUEWE+
z5NbMFQZSawYMiO5SJ+W72dLo0RMJnnqY81Xxot9Z0h1PNd3+lRuIcyJPOVi4KYc
/ljLc7M/aAfTNg9Uy20WlfD8/GijBmeK5tyfvOgdAJW4kdIznYyp6FYMk400Z2CD
gAOUd9OTxzWQW5YqwEX7JsoHYBDSv4YAYfAe1cEaPMNEH66xDSETKwXqrjlSp0ue
Z088if8w3+HiRRgHW1dZBxnsYMKzyCxn6oQJtakBUI7Yo4eJIecIn/a/vExE4B3a
rVO8SM/FUg5P02dusKVaXy6jnOXOXRv7vZq4BMRAo2yvA1+bRgC8wXVQmW7uxCZY
LJkPP34I0w+Dy5IpSKs0Nhqa9R48JXgZ/UHWzmKmkJQyAiR/AFMseSHB7IyZpUdB
pXd2HTaPV8SAJAftFcfDSfnFBx1oAhpNh/KroqkeVtyuMUr3IyFZLjrNIi04Ab/2
5uKbr7BsfLz50ub7WW+lzSSQcjND0o0fnQDMiNdwWQ/FfhwyQ73WiuLgbifLJySd
8zzIxEyg/lVL90vnVTBgUUPHMaQzQTM/uPPfDc9yQzQbB++oQl4z+Vqk8b8kGRfC
zZQ+jKiSCQrUfX7ytUbwbgSaj1Yq/4GM0mTZJe6MZHaKhYAmRZ9S+HpXJhRNPj5w
YhUZ3/2wZcywwa6BoCnUiPyPhhUQJN9HmQitKa7Aa3vkGRuELUMHP3ZsK2Nm7zm/
KY+KGmPDK5lCV1WYHohCWaTROs59/eyVyy86WM+UA1Va38aJnb4xQoR7BZZeDRoq
FxuQOnZBrp3VvUX5V3Qj2kr9DAjNtW0dLGASrR2blpsydyG0+x50kzhAfmWFuo8A
34LNMvgxzbBvvI5B05OFyZXcIAlxglI6ID5ZXUnnr9opUN/Z/tkzbhyin8VBQxrK
muGbdeqQJ/IgE4SfOojuKTouUNyZKJaz4dtX+To5S5+uFxIUrI52kJLPZP96El7S
bKeFoKSqUv+INC3O39DMzX3FU3nW04R+DoFQxTiprc/yUFh1i5PW0ZuICrst8eii
NdjpEwNBnpN0j1KG+UFsZUDz5j2JX1Cg8WY4BIY4QTJOB2t9KaADwPl/wFTKLMaq
wH2hNlpwMj67ffxPDBnU0OkIPCYrjTLW8ZDFAALy9dfoIsJSxC990S/YWvmpdgsR
OLoST/1dgeQTjFrsNkA3dezA4bahnW0wlUcZscF+QOuVdUChfCc0qjH88IpH3wWi
1Q2ESQa+2vZ2IX2JuLmLqQea1hFRJSPYXjfur+mjKhYx/cC1DgnSGT0jkvLTtfm4
xBwOgx0L8BmyBBbBkR0ZccPes37w5sOIUq/9rkI4Mo5Zp5xrpYxnTb98BEpX2FE0
bUQn8Rf8SL69PNLg4Rijz8tr4he2dARaJH17YciL3VNExlu2SvazhbZChcLvzDpb
igAnAbGFNcl65pwwlthqg7Ry1+UxDzovJ2UbtvE9sXcAXeVHcpsHlnECSsP/uCyW
7maS5tR+ZRAMmBDSrJJP1kQukxIAMXYhw2yyglkiSwbiyIlwfv201F0bJLUZ8g+3
xRzN8np1QbsuOu6BDtDmX04SwBhP0Z9HaWzjUoj5y4Nlo2NCRYtXV4DOpm317uqr
QDdDKxsBFJ/OGXbXuRLaJvzx+ZkXk72hQNoUd1rAUk0H2y9vyfk1dUv2AjTDFt1d
YS7/owOQZdMVDMEwFp0wIQ3nxkQsTbtLREY/viJmjNY/3zaDQq9MVGzB5Pk4Rp3t
Zja+xlyXKMCilvDn47jqAYQ5xhn80XfjB0YKIwrnKmruXxBIAekZZFOAeLZ5MqeH
fUMescb4/Fk3GM1BpGFnzkaptaeRgol1yV9EFbKEd1k04EerU6ZLIHhIMe6xCk2o
UObBA4LYQQazaKB3EwiPU8XFOYFzOBWDZ1+1xOr3azLMkB80eDWAdMq4Wrz8gUEB
E/O1f1/bEMz05UmwGhpyen93r+SFNrkDSb1vvItJM/Q2Utb/7o8QE/ER9+vg1UbP
Ufi+D6Mjb0yO2MsGAToKtxQVLSzDk9mXtpFC5iSnVlab+seIDZcsSj5sGX8BG9rV
yZC41uTEyHp3rfCPxhzjSZGcu7Sl4NMZja6UyKG6ANvQa4Pi1/DWAGtsHbasS9qS
plxeD9p/uAW5aXl0jXTV6KX/kB6EBZzG4dSP3qUfEfKuyDKNt5PEGgSnDh5HmM8J
fZVWiX8SJvkAEyc9nd3lRmMm8W9AxcXzVo+SNcS8/cSDvJ16yGcmv8sB9QxYhrC0
NWVN+eWz9yZHcuOETs/HJ3/+MatAxHWhjbxgp0yeb1dfCOzMyiPm+i0JgnP61R22
r9Cyt3pHS9F0ytAKT/5016eEZ7ssM1+cP6SNxgQjc891/32Lv3NpJOy2eYbjXcFX
SpCUufEpM9axCg2j175G/WcXSE4MBrcoLTQNqjgdVAhb65JrGrDKz1pq8asDYSrx
z9KiXQ1PJg1Gz18fpolFets6WfATMKonsgPI3sxokd0iSb+Q4uwyuEsb/ijNtQRZ
xlkSNR74ZIbdcPejeYtoXWB5+Wo5ZkbBv1BowatAmDWX0ZLjJgWppOgr7Fi/6m5w
k90et4zRy5vQsT3DR5eIYyeMiWex4qoelpG5muRSPThZPX4/qfoxPJRt+8IyQhQ1
kAoJ/LRbctYb9P7DcOLX3yKEnIzo+F3LlktN9UndkF8VxJX9ibY/wc3NSb7JoO4g
EHJzgb2lKyayXrwUKinvKWl3g1ebFz/ZknUWWu71arq896T0rtZ7Qz7unAi6gdU/
7HgT7ph+VtjXMO5OnqnYn1wO3/ScIW0hm3mCG6ngGwTp0BPgozYqGHlT4e8diCzg
MTMuZSHdoeUUyjJcg1cPYxxAyTrKTLacMaBcpg7zy7wafMdRdzMBojsazCuYxSPz
KYhMYhOrQGn9mh/ZBmuvanGs0VfaK1W5Q4g1s72lzSwAu9l9ZLmN/Nnf9C5kNrXZ
ggZU9tbvH/+GViQL04YnshgfbhzMUyjT5wjJ6IvQVL/+AJFHlPZMtUwlgz+jxU0c
STO8JpdRJKcH7SWHyaPzotTROTJ9dYjq4M8pgnySHw8byIWFw/NH/EnvDiDCYwRq
mNwxpnZkxknm/CFIY0rYxAZ7he+LKcDbvT/yLqV7sfaNyB9rEDv6HCBxUN8w0E4L
TniWk2q1/FNnBfwAa0ySSDDSJ+ndOVkvndjDMSb81vMKYSTmONruebG5YK9gyc3/
0BpBBpWLQGP4iNl6j8krTqp8LCOeLwv3Ws3cIXKiQebiGapL5yfn49cdomAXsf4R
Km8SWHi4xR/PosPMqYKaSX6KvOb42uaP09Z4/xKaBF6sKFZzlAdJxy795wyMXHZr
iJPuJg7V97+dfKntzeZYkhkCtxqwxCTtNFsIlxDkWMniKNdll/sbzSb4pBEHlps5
A1MCif/rhz3ZFfQL+J30wa5NWSBJU2N3k5O90PHPyDDCNBhbxKQe5kiDzmZ/VVba
M618WAxKEI3ssH2sQUCP/hixeLb8S1BerNYzs4LuxMdNHeM1ScW6qdX2Vrr0yKqe
TUSstK6v+/Xjs7+k9FpFD7sAchlGWNr5AbGWgY0TPuCyKvemBnnm4CuhHCDccOBP
dX7P9XHKo6kspAeDapv0/srbt+EMq3GQeFqJRTjnsbYJAtOhlkP8LO5BW0rq6Oyw
dxZKP+j25XcoX6f0nMpQwKz3bQRXfj6xwuswLflTJvDMsVS4ohcmBya3O9yDBvFs
8JHxdsZfT03XedREWnLiZmV9onNqPA/WwiTrHtNVhPJFGd2uvqJi9byIwWPhXrT0
fkkutKs8lIDRjj3DmNaOw32HsdOL8RBMyTq3tFP9fZ+zf8tRxmNJ4cqjpeDrligw
8pZrOTv5EMvjfWDmxmDfWcuO09TQZKPjvf+g4bBPA6hnlZW9yhkQ7yrAyDx7ORYo
DRVKDtAGcoJ9yU5H7jBYahYz8JUWjOEDQECWWEybe1CicMnt0xbMmwKHL31NZT69
mxGeC1o5FEBGDtwIwYYW1hbmN/jVvuZTliyr+BzCOLRxflK8YqSXkIGQSSScpFl5
FQbcHWnQ5PgoxtOY6a9T5KY3RHpC5A/ELaA9e1WgdsNv1skmm+Oq9LCEg1GT00I9
SE89Wx6H9Z/StT3JfA0KJvFtJgvolwyBkOCKU3E7RG5HBH9MdvqKX8DJIm4xodxW
KtZO53NAfXjpVIaqcXUA5PX6bo8/VzUFN9PMMFrfPfYof1h/XR1EUP7tsPyRRWWC
vUY4uBo9Y+QtRnlgbUyG6AHhZ16Z5iBioWTbYi5KTP2DUUTEOlrCvSYb6qwYAN9x
aH6bqB4/mxUEDj643gCECVPyK7IOfar5ddXtX1MrFXCY6QtzuVPg4BAcMMAaaR49
MzfteAXx85a36Gs74oTM68d8xhOPe2M6fH2xqi7tRbgptus3w2QtHz3gQhfW2MjC
4wo9Eq6bHNmlGsBEep51l4QUgb9KnFpK0CdBYX8FAY7bmJ5JvEUYUtzh7JQ3cV/s
YSFR4dOaox/76YG0uoniY4Jkh9zq8RIxAxCHRoJ3OL/1krAI7/28V2wEmzPUHb1d
Qdm4/zHjtCyauIcPPvq0GUhHNSggBbJIbI30dKKdbZRZnrZq1SisS4UEmlKSM7P6
1QnagTwuzwljuLI/3rhbL9Z8vVSnjKuJcWbpo28bmKVeVWgqLWhZd4h43fIKepe/
bE8k54gYF3vQ6j/XGw2+Pa+r9XipXFDkpvv6NXMdf7GKgHLLe8FQMqnWYH3tRXDR
HMeykRELFuM3KE8olmtUXyhqd8mj+vnr9PHHDiIP7vOl5RXBJpO9dltbUYIrRr+J
fMpMXtT7LbRkvQHPmAQFGdBQUuU5UajusUynK7Cx2soWxuc6lgONq58ESJCWJHWW
mh5s1HmMqvLxVodQm+8sSIHJwRrN0VdBB5qlK9qIfnsf/5m2BmHtjUli6xV+1b68
XLZygzvHZYrf05yspXE7RNdWzifZ1cfURZWVWCkNL61dbGIanmf1bugIDF0aBfcJ
CUlxgFf5GaKOygm3CvHVnhyEHBGuZQgm4PyCLCicXU+b94XJcomZ92UBmSRFEtUb
NhgEDg+mAztmwxCH2oufD5FOlKUNpE2NNMVEMwqhrFKsIBsdiCBKr3Mik48yJU/7
sgGj/njo4GoWiVHTU1zvHXRe50O1zsUlX9BPBo9yvGpkMRp3+EvooBB5WnPk80bq
vht/TB4mbfcLm+uao0ZGU90FSVk98dTjslfeaqGQmoRdEOMvRp209VTKkHZaBo3m
AOcwa4W2g7cn2QKg4/WgxiPJp14ifWNhkDjRY/aqk4hyYe0cs7g5K1rc9c63fQva
ZL73Pp0pX3OUemv+ji7BkRlvkAs0KDYncLXGihapfWPOiq8k1nPTI0hCmASa1tu0
nv9xVD7KENZT0+Z2lYzwKeC7W7/zKgoqYH4jqi/eI6vBAKJLhBqXFASOe3YY8+YT
wSygb+pm8lcwzzQkP9WtOpVtUb2IiYBW3hUtVT4HbBPoKak7VH02hq8d938diNhM
05BdoezlZP+MazI1FIJQ7siwwerCgm98cAJ3FeYl8FlZrJB2n8jwbO711TaypSZr
qbm1TwRO6XE165L6xwn01CsGSl8JCksa5XIVCeG7HFvRKfRifKYJTVDkJTf/ZYdP
2bosYUYFmX8A2yd8RkmF7XSRsTnTsEW1/5wDJ8MlvULhVtuOuv4ZYqcw5L/FlGhu
JwmrRIwRzZ8ow6I9Sn42MIjCuudGtOoyPIB6f74/W7F7M+NknnwNc8U1ZB3OG/yP
tX5Z5kn1SUiL8OuMyYA+AqVuWvbe1UDDatUXUGhnNaZx8waE+w0Ek4HW3qS1V2Pa
zyAYJMQHrWmezZwjYkJ0+dNWw8VqH5u1OClQ69YKjOgmVWwXXjxCz2bjaY2SXPo/
7pnvCONRTN9hZRMr5aCmnme72+Qastc6SGdJLa/iMWD9Rsl7q/wfhHQd5wZ2qLp2
wpP17h+j87le2g7ITpDi8T16XEEngUmWSP/Aje1gDqJ6M8UrqSQLbcMWQMMcyOmP
OSVcwOpubULPedpyMNV4s3x5V7morR/b4CfppeltV3mWoh4PR3/BH1jIkzt5hERr
ZXuj69RIYbi8+kl1lQLAsCv79IYrs41Lf/Dg/RWAbzKgnIvvIYmriwvywK8CtSxY
kBhAjxvuoTls/1Z294BXUHadUOC10IBniCLVumC6nWVFmDvTvfOX/G2H/bwZY6mD
vwqSc3vcBk4SzXerSHy2VXSoWJwuB4iuCDGyo52mfeGWJeQRmU0aDkFCn1qlZQRf
bkd0AK1Wn6uAVTMJs2E5Km3Urnn0B3hXqNM6amF+MzQ7EaPQwkzzBnJhl9OZO6zU
Nz1vT831BoKii1dO2zhH+ivwQux/CM3NjUrk00//QWSAhwlXctS3f3d8mItdR4X6
nARtdkwDFecquBJvFjfkuA2JjYlqoQ771H6vcO+ATagNXOcvzJDoDyIO15d1/Nz8
+JWwlX/lt+LIU6eVtk1xnxyBdoTH1maIJwHUvoxyXC1mc+S21pkZIQfEVCc5Q6dM
NupdK5n3epabNJ7T1jMnOspuettUKaVWM2IHJU0o000x6XYWckNJhxVmgV5jZsvN
M3u5AurI93T1I7bcgDrlMhSp3nlH8r4N+mxKeqrqyk4rMNSC5oq43cx36XM2k2Lw
5ims/0TVyhovohiK7E6lRMHa0o8nnvx+n7+bNmZnzCdqppdtGuxJzhJqWF7MNH3G
YYDnPC7vZoG7ra82cKdFSSCYrWg4erd3S/3fFC0KzPI08yuYPCV/xrI0/94r5cPU
ZcOwzUTO3OyMc44i1c9rKl6oB3GS8bmm5XOeIw0wIHMXZPCaGfnnsUmeWOtfzPYr
Ji7JrCFXKGOiyOpwmbY/b/j3SOkDiBTF6j6tF8nDVqkBV9ehz/NXaQ/Ah0qibIOH
Q64cgchPQ/oAdzlPKNrxavtA+SgX4vCMyyPhutFaTDQXBSgwuBJjAhO3f6m9Z1vn
6vQdEhNlM0L5jNNy7zbBkfcS3xR7ceUrAd9UxvwSRI1C/WRydOAF5iMqFyQhVKqD
kKt89mw9kKfhYBsqENb19k4U/YrTB5QpYKESr/JTphNc/nyskih8AjyvsF45PE2Z
0Xxm8Tel9xdsAWJDVUm9B+Y+whcwkI69CsrqvgI4z5+4mmlJM1Z/NnUSrtg/VWe2
SkKzIdr+vz+TQy+AwUVSqM6r0c0VmUAwFV5nRkIMLFaIHw/OQEH166e4IKiu1KGI
Ok5XsrRD2+ErB2QCEhzlCkkeIyo8GftCbwhT+R4H8ZSF7OO9NpV7HYh57YuGe0Gn
rNXVn6VBDyeswtm4ZkXGGlK1UqZhS6wbTS67JYyoU9DE7B32S/O3BU8kQYXH7BWU
CCmoISNGCNzb0T3R2KHW5v2b0lceJ3eiUTwLkC82k8v6Pna6RrCepRk7fEbYhhMK
ij8snpBk29EMN3Q3MjzvG3YGvkr5xwzavedooud2RD6YHSu/MsWcG4AGaQI8UtED
`pragma protect end_protected
