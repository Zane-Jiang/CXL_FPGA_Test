// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UuflD+ofMLHlYOMTcUxCeOcpuOv20WP0Iwnx4mMmQFCWfWK+O9u/UKsmm5LY
Otvl9CVHaTPclIEj6yXOHmSDYZqyx6Nykj+OBEpA6fzH0/iOSOgOGwHzYjQn
wp4lcZfH8bINFTGIy8u7BbpsubC6R/fHjkultJ0xrhbj0O4IsfLuk4HEEi4y
Qa4yXBPUORsIkTb+zAE14iFjGcoPd8+QxkI1R3KdCaDy4wSCy66o8IyuFrsW
bBw7MIEh6LrqBNOHisb4XIho8u6giyk8SzfJKg2UQnmCcKAzGWsNCJiqsAL/
kJMnVtbnLax3l1R1sqghQt5s3Hf8Sem9BVChoNUToA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O/whr9QkQBEz5Y3wgnauL3Sf4TrOOnnSl7FmLkINCS77Oz4idQx58u4jI7sZ
TxpDXEp1yZ6JoBBJ3nzCNvsiUQU1kbvjQxSlaN6grR2gcDT4sdd5wTGm0SPM
sPW5+P3oTEpdOnWwHlhHYreUnEiUQCXrMrLpi9yISuS/vOTpcvNn3wurPJdg
xmwiDRKDD8i4zYPCBA1TRatVnOdMB+8glziepg0bAWlNoy1WItmhWNzimsF3
zY2ukUp733klKv0kxSclhCdF6DcastJkoGIXLbJ6bNsDpAyfle3a8WmXFNUR
xmmt2V1j4FkMlfUqTi42ExRDi58w7V+sygfYWNj19g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KyMXS6NxEUDv/y3ziytpnEmY/mRj1zRfnCbl89lfV2+rWFlKELukiuovP2kk
lGSYtbruGKBEDSusuyJSfsWJ5kKUNIoraE7grl8mPi6OhL+tYCyFSqQqxuG1
s0VnxCCtFrYE19ZYgn1TWveYl+ip17WiVm+Rp7e5qDq7IiFOjEk7mfuSh4V9
YolKSgG4/drSx/YToSeCMd2Eh6HNtBlHGHqAxt/xQ/fG2FtvIQk9E+FYzGBb
I17Zny0CSq1raBENtNckpkmhjJco13BbkIT00DFOBqq5Noz8amwOSDJHRz4i
TF96O8CbEJ3GYETvNHxu66L/jBKnn/8FosK1fHxpCw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
U/wADd3I/YWlZNZub0gCRflnk/JPqi1UPkK90hCzp7SSu7ldfYPWSe0MKfKf
UA1OQCD/bznDxPI+Dbdlg/TRwoYSE/hcCucKXCA0Wz4ju42tzszLo4Ux+uR4
52kKN0GXLy1eu3kxPX+h9kvBEBwUKNqo1CFOSP7NuEKOs4sgpv0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jD744X98m8gCakMmwJ4XUTC0AGxfnNV4EyTWp/gY8VnwHhQRYNFk1qG9A1po
OksO5Y7hmaHGV8jjdc6P5Kfx9VeAfvE7jhpGds6V3Xnbx5Ng//kO3IlF31+/
RXerup8LMKnW3Dd4Va+sd0LCV/cFfTDN2MMKXFgaDq59naSXq8SJ49qULfdG
nt0Qw9iIPOoDs4CBHw/oNlGe1IV8d56Q3b/3dnJ948ATGy0ur+x+O6mM20cp
ahtZrntvuy+6fUcU4niYYLGk0/cho5Lmzu5VhkyHaNAmR+bMgFDp8I4kxZbY
2IMZOg0NrxL5DsWWoLUJnAIQfaQ7x+YipeQK8dTBjOOOf7dFgVBPVkY1tux1
DuqVtdZ81kQKn+jrsCCCJ6ofaYuSw6zBbbSuGR2Y2wSUtpq3lbEOP1u/Gb6c
YS0yeq6spcF5KjsySGKdJpo2Tn1Pj+ssnjcCjBeYZWPPBHEuba6jq1akb088
LGC4Hto0hXe23yxiiaPZC6d4dpqh9DN0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
l9cZJvS2fWGhQOAsWyLU+LdtqX0vLHoE1pK/8nqtsK7f6T5Z4/YMW4H+hbTD
EoKy6MkZwL6itkBhC3ODipyaj6uQCmDSGr3a84hxzG5iWy/TcraeLJTT+DIH
VdFp1PPcCpxRriEVm6CCIsNEIc3zKIOwEV+EFdJPHO/mzNN1ZnE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Veghzfkju4v+u7f2LHc3Ee4lujENRp/EUhh2X3pB7hpQ6CxcZRcPdSJHzz0B
IM4WCYVw25koFk57NWAUR8PkO2d+VAjNYobBRROO8wajVbQrHpCjh/7iLABi
gjly6hr0Nslnf5YD3TroyHsAMbuowG9mbphPY8/NkKJUi4R/SDw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 90720)
`pragma protect data_block
7zGn02sph5+6+dtSUxs0eD3yWswZA0436dclADU52K9oAknmOCODlNYSqdcX
v9/xQp6rMK6uHkZMfduSRou5hGDwx0JbCHrb74XKbKGu0heduzcJhCcraWgd
O9ukWScLiGb7ewxH8V3/pR+cOzShiSXpSCnxKfs3mA2oreUyMVrptE3y3HIL
evL9eWi/xUXwFHXAJVzcnjpveNgrFntd7wOC6UK5S6zdY9KAyqudoQmuPbgb
Dw1HNOPCwowfZVM/7KW31VToyeSumu+n7mQf12PNk2B5NZxrGrIy5xcDvF2N
UyyciF5iBAb8RJVjpjtRKUilouLu0F9DkWf2WRPTrQ8pGATJFW4vyoOoJscg
09hFCLE6Vo8HkrdTkMfmIyYWjOPcAvRSqS+ZRsNpX3DAvKkDvG9+b5/nuClG
BFPbeOc7qygPP7wX+wxgH8XRr9q9e3HTCC7SVUAFyJ0DRAEadiizITd/A7Et
989WVB/b5g7oAZco60Rsdh+oJfmArmWobMthxyH0fON2DVLp0Y2ejJyoR9Dz
4P3vydyKKYmvcQ6miGtMz188DNJWZjeuNn5ACRTg+H+mOGIFgnG+0b3RtYit
dDXua2POdZdd9NRjd6kDUv6ll0oYqIAOMQw2rPbtcCVItCXIAc5WUKqfJIh2
LjDJXGC2Uw37QyzcqlnEVSC3YqP8TOIdmSs/0XCTtIoU6lbE4CRE6/5NBzbU
H1eAT5GHVdHOCg6NFMnm4pCyVOOpo7leaGsweNN3Voq8sXQWZPzT9Ir+Yx9n
BLZyNUh7gHBgA/K6zGhgAPtq7dx67hAKd5MXdaVGZFmyTGyN18+57Vytd/h4
YG/td/GdanHr4ea4yFZIAnivoXoDtlXS6FMyikY9PsVkeKaIm2np0QVLGb0h
Y/590pei/Ie5thYWMLVZ4CWld4Kb/32gTIBQnTkW+YvJNt+Ai/LKkPgsIc9z
FgpeuJR7t541yrpQjfvgcTkmix/UP8yQl2ZqNwHz7HrfaJhh8nI4b4Ev5j92
evHtmySNzDaqBN2DVBaEp+lqWJoay/lLlkwgf4jafyN7t1a0AvzHUw8pQvJS
o9BloW5rGW35fGlN8T45AzRp+7i7faAEpFfwkn7WwkAy+jpwtPT1cuE/F97z
WIoH1v5vJLphfStA8ABGzHhMtv730A0Spcc1MyHqShBaNNgaJQAibj7LRDT7
BUiHc4o0BoFMY6WjRBXyYs2AU0D4R2WHkMml1GyMFcS5bgUeIzC5ow+CNKpp
xkZCsCbMWF78i+39NAJuxpG7o/GSTpJ4jhTZpAsM0zjGeBenudZpkR2TxvdE
s+MQMAhYjl0oelmUt+wmNUhEUJ/ybMTUifYWb9vm55LciC8n8sGD/WgGeugC
5e9W4d+NlLNI9Bf0yvGf9aFJ8mpCRiOuole0OiRzgKE0othbF9E/0zh/SAQC
7QM0zF0E7BEOl6/zAF+YlFXmDliB8LF9ZrWp9C+973L0MwhZNSWy4k9Ogb8B
ROtm0bJaiXmabZcR3p449GWfoVFeoyPsVwr4J2x4kGhYXiO2j/xPZCeN/wyH
g2by569JGs+zeOtdj1WyattvQFkQmRd7CBOU39sIlNJM1S0WhKFRyDBNafic
062nSuQB7RiC/NvXQU3DO9LSQ8bOH4Qqmn3Rff/yL2E/YNX9XY2Hvg/Gtvzo
rHeFdOr91rcb1y+mo/5xHbpC6DxYNevB3kSFoJfjqbpImElue+fjDzXAbzjD
U6/FwGKw100S3zSW3G4JWTj8yJfc2Q/wX9fT7JetGZfwFQy0rKYU1RzpEBS9
bxmmTkL6nqO49Cb1eD7keEmt0YtX8yYSK7lt2XkEqV6WvKgf1Rd4747uiYk0
ke5ew2J8OqlSGTTz++uU+KJzmlF8pIczttAlh3yt9Ff3vE4D9QpGwv9dld0H
IqOVrFeaKZimSu2voqzrOl1LNUueaOiPe/jEOG4UPEc+o0G4FNPUgVe4ongP
O8qnbK5yyC8u1yiW6rK32xgIYBAciTM8RWuD89+qvxMEf3EGHjdVV4R1ZZTK
cBYOHSVnVdVKcyIxC4ftWvtYnmWT+RFw7V8zDX/QEUeTk8t5PdF4uibo6ES7
9bPUeJ9E83vu100pBqqZQQNsXvmLXi1ikEKpW0ZpF0I6SFA+i8if1wpIyezF
IIRf20PtIOHRoDJRIRz0WxYBeKvG6QAHW0H51NPcL/Pu69FsDlhnPVIviwPF
TzgJmqohXKFiOQrGWVILM0HuVIU7p6sj4ufzx6bIHgaRMaCXZdUV9nu/m7D5
Xi4yw4xKkfGqtHd8wCqHcvsE2nyRrZ4JHNkKM7El+j0df4Ix7yG8/e2qTrwv
CyxZ4hIxDTApQfBj7Jaz6KHzZzbAm0fFhX/6IZZ/ZFjtJjQ1W34P3I+qGF89
jEcL0/Gh+kI6NqcM7MdDsZdSWdY5p4+h7hCp7C2YBJ+dciUGGgoq2CY+G/oQ
YfTuZiXhlnDWspvJ0qdntlZ0NE06p1QBxh6D5/S32kWPJFIMMYCqqVjRzLOL
oghktVBHAVegwcgvkhGXnVwwDWRIuJeO6fYSPFGhVuGyl2Vt7hEy/O4o5hsO
wPv8fU2XFDpEIrqCB73Y81v1x3YV2UqEBkmR7ohRTWOMlfTIjXfGL5SA/khs
MEulnK8oU0xoCAh9kkjzBkZccMHm+yVzHZB/USV4orlE60pHJXfQU9Qn673F
TBpaqIPawPn11cZ3QPLA8ZnEWKj23hvyumK6JPVsP9B1OeZ1G1/4LT+s5lim
xmlXYIFAD0/qiyTPsXfZxM7xxd6miUQ3lC3K82/F3QthPNGrBa1UBHTJQHwd
ZGYf/wTchkOA859VyLCYA9COTRBxUCezvgtspmdKfMo8pIeWIwmsv7vbQS9F
c25BwEZ+nXq8mBGVKkO2xDl0UG57I03NhWAS5qp6lsrVNrdUokZ8g8KuMw8Y
F4T312ScYOUKwalYqfy/j7+qox10xu18P+A4f71Umqf9i5IpxspYYV0UqpLW
wNuUepUVVmoVBJZPZLA+j7oYtUfXARAwJnQMZbdGsXBskdIiTv1XCn0XID0p
Ar00GZ/CvjdNjH3lQSgonL6+8pLuI9g56LQBTJYAPqYrRw+NBjWxkeap7cw6
l0sh7CC07UHLm7eP/E25/p6rp7+EMz42j3xC+ViAtN6GdyhTF9jiYzrVp+12
FbcCVu8KRut4W013aq/9tyz4cr6Q/hv2XS2fOcyJu8FwSBcnz5yqrVwzd6BW
MGvJhyrUdeDPlQoyquoLxN+vTx7LsaORuSiUV3/rqTpib7aAVLVGbc2o4qI/
mEQTRL3THJACsx6Wji+TCBvORJD6aK6gbb3F7MVu/oBvL0/vNOzeFXb3alj2
0Wvv2LaU/jlqgTFgTdGTY+ufpqBPfKa6KLuhG9biXt1HfX7JCiwWxWO+iIPY
iGCxqRz5Jmq+4HkMmfLQmp/ZfzdxKKAdHyUADIqk1hawK48vlI9udCiHphr0
v76ztedpiEN6/+jmlg3EBSw3n8znED2xk7nwoyu+pOKnMMuMhNCEX6wEalHx
phwGY57TYcuHqMgqm4mIw5erRVCHL/YEjhl9wjZpf1AHxL42yz4c8dHhEECL
66frVI7wWjKrlRBxuMgPt4ZPO5xAGAhBAxjobP11otQwaTbgqc3L6w4wSfQ7
gw6wCGqD6CBmqoPexsgGQdKZXxgJlxGtLnfRtSnWtGI64GYiPcUlsfOtKuVB
NWsVFEbqlwRfq9lfanKITKRGDhzbY35yTadZaT+wEPd1WEuIMlZf0F4hhzMY
ysAZ2fC2CYxlHfQTtUSXZ8MFDPuDC4obJ1iPSFL7ng8IePMoXTi8xKzz7MjU
8pn8FAZnKOBXnG4iccB5W67nu5pH+1SkWOVlLv5j4LFjd9PuuaRC4TP1Dp8z
Y4Ap6mTjzzy+oC2C9yq+jns2TeFm0mn9+5iU8gmD8+MATrEGTXEllveA3A+s
C6K8XOw7lLXUr1+HQup/btpIP1wGN7LXwVChSG3ZwEAbyi6wviGNTCqBiygV
za+4hcyvr5d1lg+TX3FVgumCm6bS/XkB5SGNBvSaY47TTw7+Bof6L3jtPgyx
qaM/q+Xrfl0gcAgPG7Xn9tK8nS0BwuK+akVHuEGZDtHB0MnvHZEfljD3EZKS
+HuPwwFPONVJeYd5ShGREmZ4IpWcO2DC4aS78o5d+jvtDIoTwXX3XUEOkSyl
zEl3vlHucE3RcpxQ/nQH+3VxvCUDVsca5R/Cdnh4se/LBHWp2BZ0zFjgSehN
GekhLwNF9yZ2UuzycMHtm7X172t+q4Nd0jKmfz7XEAnuxxpRWO3SJ92F91qy
671e4m7vrZjFeGLPgdxMeLDkQQid0yOmdZpENzcJml8L87xN7yHZRMl/ovFh
+IpKeh84p0iHVxlZ9FbEa3d3v+752WAnjXAgIBaQJVbSZKLlDq2wbgqdRkdi
hlnAlk/AG4ffwzcNnE4jJkeQT8dkMSPi8+JaopxQJ7g3p49b57m6JzJVtR/F
LIKboKJ029d9SSDgcdB7kQO+odNaBy4VrCKW9DV89/c1ay14sPIBkt9zPAJN
V/EiIYJiGdj61BRe81Sh7Wuc5rRV4KKHvGhoFYOAuncSp9rL8Gk16L4LNacf
baXOn48j4G3gU3Ihxf8TCM6jqareHY0Bf2YbjuqFUujEwwotTGUB/Dg3R1Fa
j1QUny5KPeU5tjadNfWFA93Ao1B/i5ZqOt5o3g0dY7GdwM6ZTwTc3bdSbOoP
HIpxihIEnlQRJ+EQsC8ruXeM6Olnx/GoV+wIqT3LIzkybhj7MnSoD5FNRVAT
eLi4OTd3qt59QTj0ooYhcRfQgSRa8W3Byw75f7xZf90dV+Y1+AFioINv0Rdl
U9g61oPSMNWzVfyRsQgerFOEjQNvJV8FsNaxRoKyXhn5VUkrjPaSr0MRTqpJ
kr79KGY5aH8Pzh67IuKinQ6AeAmII/10BLD6YA9b22XSpLXjtbqu6R8Jp/T7
g0ZXKMx5R02vLztDQn/tYTEwS35n+tHivcqV+2QC25WFXTwz+QVg5xNfrypn
oTZs2ELwQAumdl8wbhR1xWeB5X9e+alwWc1qFzLvbENIZ5TzyG4EOyNvZso4
heFwXGC+E1t8bxls0pZJ2QnjeyO04lkv6g2boTk8Tlrm0rKT8uValgWW3qoH
iSlaJoK7Q7+YK9NrcNO1Lf7uj1KSIxBh67vUnij8O+bkh35pPS72SkXy9O3s
VGCieI7i7sDiseFmimJgZVK1sJ1m6RXZnutGo3gm5+Az60RS2lYoLuGPBVzK
NuvhHH6SdqZ9RQN1qJ5z30YV9qikkYkoH0qqBWUCo0EI4UVrJOMPX8cXRccv
rpTAjBX9Ah/gHOCOR/+AY0vUo+V0nSSz7i1hn+s0fKIrTMI24dyOz6UadnIx
RbZwC5R+7B0WDvDvVU7boUVrvCODYm/2XF0l8cCuXqB4GkINWjCJbGquC8Ed
d2/0U4smczn82jcsIC9XmN0V5DnoBHJE/rHGsSXeRX2sPFCrccJqNNLirMDh
7GqdksegVCT40+KyySUJRCb6OhdNKnPVTl25+37zDA9Y+iUgiyyXbufol9tK
ks6UyDGupPi8xMnlwLd3kRE3ZRp4kZHKxJ3mYIJ2ohL5pbpLmBod19YlzGTz
fxTDBYyiHXxgVnC3ojWng2DI0JL/+koU3mbACZsyKYNb1UMIB/DZCqSHyep0
HZUGBatFzb1kR+NDIOaqUiJgNwsWoBI+hCiX3aJ5nCs1xnGgFGKIqwm1hzwb
lgl3BvnLpARXmL2JRutnifPXjFieD+49S61hfau2I1ZfEQEwnySY2YvZJjSc
zvGb7c+8HxenGiVQnnlK1ELDdrUt9lTHnlM7N7Zp2/sBQmJ2lzFDwAam6cVz
DdAoTcKIzXhr34jqaLO+H/1ltTZdeULfVKigcFS8wfQV7yJoPX9rgdIul27s
siINGzNHsInGFqo3DHA+6GYewMiLNiyIEu/vFWvL+0nNapaOZKyGfR92/Xwg
jjbg2lomAlD/aTuzcKmOe8Z6k79D5dzEh/sUuxsL7c5RsEcwXJc7yN5KWAN6
/VST99ZK8vmBVg2FQgq9OLPytHpDN7zmBx2FjMWPYluIyVNWxDE+PLI9azOp
c8b9T7fzs+Mk+RI2k8Xi0f1oR5L/3eTph+IBd61RE3yCk+BnFBTunPUNsaez
cUptx9tjb6FZY6NP82fTWk8j6aICCkWWSN/4GogF+eUkG2HuPYxKMd6ENL38
6E9582TxAMeawjqM1YME+u1KRnuREpPqggW17yOBUNpeuk0tXDUUAv27VzKP
naUqkkKRkH4gnenDUgScy2BvTwJAgmXMJ3SiAlB5RwgSlBCORQA5gKdUVA/q
7B0OASEJyKxcoRpMUuJjW33aUTY8buUvuq7oDxJA8lzClMO/hSrSY1oyIj+4
V9Pl/AO567DFZDN1CVAdlsxWwS8eQNWXIZz6fIJUEZqC+84OIMHjlPe2I+Pd
e/iOaR1FQvuC/G9E+jDUmiTjq446Mb6iPNYLSZPwUKYFhbefAh+jFmaMleZG
8DeUP1woPA8/WIICbDM0OsjTLn8w9125Vn+yshVLuDZPosUluTQxH+nVEvOD
p1M1BH9rwx4ZipBGV22jJWgSCJO+wkIUhk1iE7Ep+ciX7dfJpey7iUR4BT0Z
NEzSq54xpyhrKAVEAzlgqQa4bLqRvljiuRQJYOegaAgMcgpUmso82jYwYwTO
iZlk8FZyeV2P7MFWB98W1/ForenXB3m/Rv2WDRfOP678gWy7LSc8QxUz08rF
mJstAjRwik44/CmHMXmcKd6Jz8fBpW2KGxivvVe1ComNI42Baxz86abkXZKd
HvvPHR+WrVn9+UWmz9/6X2Lb1PUHODM89VbKupyFTmVSdl6Fb93iCFSX6pRE
XWMZtQJpgQhWL1qwK1w8Ju2vU+XnDcfq4vfcxFeVsaaob3vOVZtjjpTq/oNv
gT/MaNXUSpp+TYOCOHncNMwzS5kP7o/N5d74r+aBJp1aR5K2kcGDnQfMxf+q
KiEQVB60pQ3eHKhpOPPvaDd85xrg17PIcP5nvjZq9R9i+/n27RXTstGEylmr
R9rcZnkg5O78GfEAckPTFJJrUikUBZ4XJNDQyCn7yIkyw+km5Jxn6IjEluHQ
qPEyuVJrLTWYdHPDG2DAZ5KHnNI78KMBdd5pT4+A7PCpBCHUsH4RmtL++dfz
rG5c5hVjy9L0tqgycZZRnUU1X3s9RW+7678Po8zzKUl2FLE9EMKUydN60bIV
/zinDzVP3fMh2No8cqRLfp8xM3aQlspzpfTPw1LAdOSIYDbA2UFWwr0NKtoZ
knUI6HoKQ6Sai//MjWOFrxItFU4zQPxwDYWjm0hI1iTsXy3/h742pJe9nDK1
7KkUyzBGmsbp1H/m4N5hissPf4xwAo0Dd4u25F3NdJEBw6AGAQHwJ9q8slAA
Wd0lbNqZnA4x69S33DN1e5GcaGQAtYZmIfd58zmaWE3uBNNeTN0iBbLPFksW
OUqAFF3C4EZhIFq/p7tEhMjwixcisizLxmZ4EpB2/a8CNu1lqTMKbGhLSCac
ZqTZzKzL6jJEhztWDblRpwxQNyembCaU1JFROrP2LxGTyGeQFHAyb8O0beW+
IowChQA0oswHA8GopEm1dHm1o41iQdntKQGdvFb3af4zT5Vgd67QDRucxC9k
ARWYclMY8lr+UFL0oH0ooTwJN6VbEJlntHel6vXTdu6aRm7gIyqOSdonhN2o
mm1lcDx83lA/SjYLdembGrJ7/POlf4/t5p9hZQs3bdg6d/erEs1xLYpmXkPw
zwGhek8lbI3Q8ZTfKNpHHOo3LOFwrLLg20j95nyuqKtwH8KOxfD2pNK+PC2Z
ZcMRxSuX/ndQgMbR8pPxhXlLe98v29cyv7uTu++vntRod2uTtVOXoT1oDpsA
Q0RQ4kFa2pMbMAZXeQv9B7m3NH9vtzLyva8bHYs4CpCz5E5woKZCzjim1jz2
sW4eWhrQJTFba7clD6Df1cYBAGTH0JORxq4TDlB1bvTgkKXylkLFWZ2ppNsB
8XQ2CiiI7/pWwKUwry/3fg/7SuXy4s14fNbUqeZ92xK1PYSMUG7UzyCkRfej
aE8mpD3IC4tQ7tfthzNOpfNp7PGb1HZxTPyv/pBmX5Rjo2a6CQyc3f14gIY7
Fzt2NS3ehiFIl4XbTc3S9ueRq7CvFbh51vOhw9Nf1h6nTqiIiZwO50RHjcZA
d0KnkQWwyxLWOLICgot/M/+J22nwYJ0AoqnU0N011Hb8/pbG7iIL+sQ03gjb
6IuwFaQQzSBlKGAtb0WGVuN3dTXNyeJDklo+NGQA0p/tPaQq8ooEbcUKGDVi
ZFwqyN3w/cJ+aC10ubHeVqeE5tuc0R1B4yFfdkysM0tmlpPufivY3GaC07Ci
CHnz68dvCped54cJzm3N3GY2VT4Pa4/tik9JtnodHNMR5HcyMC+puxV5yydJ
j5NfroYn78oT0+QYiOsbrwpJlmhV5WeShAhYuXPN/k9juGoRRfK6MPcEFi/i
EzlcPzh2LjFzxyGyTmYkyKPmyAUvIrVCtIpkW7ae1xjOEsA6E5M93nAwf39F
g6CSjG5wkUiiYNCiVQNyep919qjBxfGjysbDrvMrP+56nYj0tARFhT4nSwmy
Ohtury/0zoCn5bOtJNP7udFy996LuOnv15IKqsoHhBVD6npVMgzTTactPVQg
RNCYusUGSdHhSvHBnP9LxHhm+f+BCH5pMxeBVZKNCBP3VKiBYhthCzY5FVxF
8J005Vc1m3apqBUhVZpxP/rYQiogcIyOVcpar88VduHjb2DnOQSmLGHqhf2/
deEAfunRYg1jG0RHKukVNbtwkr/SCz1QwKXa8BfaQxROiWhEebd+7t+2OY0B
bnafvFI0XEuGxi4Hd227qIMwW3dxN59z51lI4QW0n0BeJYf99bamTmmsYx3r
AB6qOB5YEDEUdNr722snVg0go3XcshXNOnsByCt2W3piRC/LWJWNZaQI3PWj
YrBDPvutUTRwajyExdiAZNdpPXcIkEAwLA752zJe1ab/vpuhJB22W0eCOaPe
YGPAYIJZVzOXIiiM3CUCvqHJMC55/iOGWsU/0Z6Jk6Cm++Bb3KcSXtyUmEwt
z9848ImfiiQcuHJJpnaga8kx7LPLg8GgBy63qsUhNB9uDtv4hiG6hDNlj7IS
MHjIP1Z/H70/zRb9tppxpIEYYmXmlH2hY/0pqrU6ZD3noeyOM20cnEPK1o7o
Qt8OovaTCYs4VhaQ1XUawX9bmg+oyamVB/E5OuKRotdKlAGQ6X9T7xdQdgiz
9KQInWC5aFc95YFr0MSLgHh0HayWJtKwUaKbuPoUFhU4eoSv+OUpzh1nu3/X
1JWIAhWi+AHQfpy/WQMeYObclKDzTVSszAQfPJgSW4Z3dxSBC34dZqy2V0ND
okKThaBY6j5eIScE8EJXaA1pxritxVQHLpCIGEUwEvyTnIU6sQw6LjxMUHKS
UibP97LcqoaqaLTQ9sAYFN7t1IKo57VrigMXscTOlLouOvu7CFbhaSPgfY/Y
fpzfwBhP9b33/so96OMuN/pr7XU/i/9IZPyqS63lXUKuoYLo+YcMFJMtLAsP
R321Ppo9H2K2WZumyitvFHHfDDCjYIRlYOP04MxMVi6G4xL1KT8bIGqJTzdN
RUf9cDD6QieT9hkYK9WgpCjLcQlqRy0lSTaxG/C8bxOVEHBtgnb7ssbSIY6s
X8WTgXQpJGE7944vjEVUGxc14xhNYN7r+K8h9rXlwFrelsSmrRIBWAh7bhXk
lsaL+w5hdeXR76bTJUcZ8zbp7FLnTX37LyznJ08sL074gFbNfwEo4mAwCMIW
2FfBiFIpzcrF7yMcgTCPFcJszOLYCpa8v4x2nEcSFZ8tzW0DuRp8iCm8xNsO
z6kucGmEHS7B8e0foA90+yhLrkzXlJB8OSzBUKv4zB0fWbXUChST2hsznLMc
1IKqrT/gpAsTF3YB3tnjFY2xLX6MgJotTTib06ZiL12ie5gjAlfdE/oLlYTn
jQ/jGMX9ehFFAvj3p5mENppSqOfuMZsqaGB0u9RdAiDtRALHWJEe5xXz7T8H
ZDyfffgo7CnJ1oXP85I92V5z4HdX9vuBTvnHHDe4j/A+/Uapp/BobXn0D3XK
VT1VZG3pIzvSNkJUpfVF4BzUbu9ZazoKDnui81LW2o6vWDy9dpoJNwi+1Qs1
OSNhs/BBgy5WpOtMh2IGcyi5lTjUoW+hStrPp8VKGqTgXYfXIboUrTigItoQ
0443GJmjrwgxfjvjihTkUa0+OajPYZKsPgWqW47X1y+3eGBkK38U6YEF+Tqb
IyHddVlo7odQZNMbTGQ4jXAUvmE9mVRaJVuSSUZluQmPHbn6cMypC2dPCb52
jnmpAU96N+PazisvfSlznYbv8c2+vkQYzbMS6N1UQbvSXPEysIHNjPmGeFna
JMy4oA+Ln0e+lMi318a6vgKGGtRtdjuqheI5OYgqd5WvfBqhXowY6KEQgt9v
rjKNHNCDYu7IDstt84EjuQds01+AeOLvB+kuLNlw30AIuOBfJD3qwBLriYWC
GYlYtRgHQ9kMvK8ZmLNb4OiKsK61sNSw2aTayiIGKvWyv8h7IRJbHcDENNoZ
eEtxY2md4ZpnMolfDqFANSm57ic7lhLLirK8/RKjTbD9xL0IFBJYUygIKC+h
5OXnSGwcVbLNiPYT02s/JAt7ny1pF4ne3xIc3sRSMVW8GXu8DnOvNiLSc974
5vHeZLO626LLnjw/9VoN7mzSv5dUUAEsJovTd734cVUxxOrPsCsXyPwcnO0j
8eFKkPhwCgpKBmTdcgHU7irAsgS797qE8rQcspk3Mx5RcxqtpkDr59z3v8pv
bLvPJX/JH1K25RguI3mEGHk95H8YBEYApUMTBCX8xWmU+R+ubaDD4YHtKX22
YEvCVZt9pMlIo3VXXLf1i5BW7JQBzwkAU8GccZK6TgVekqQXAzbrjJQTwFRq
zEFYNG+HWpvBUUdhAdG+HCnLTZwzVdZFP7OkZUc5d3b7Fus1turE1j9JkCn4
WM4+NJMVmEHW8FM6UfU5lRZSAp94d4xdSVXR1SU68HkO0e/dSGsm9FOZ7G8y
6M3yjSKcSaQMovQ2/rC/1obeuTm7bvSfrX2RiNnJgyOnXJu5hhLa9ozsJnLh
0zalXJMzxhwmT50dTx4+4OIlrJ6eHXinOX0Qp6IGwuWgHKCuhANwxymY4tJN
CAzqt8fxaqo4Y+jrR+etVtwOxY615IxjDw0lG7Ew2rkhAXuqz9V5+d238G5w
2NYMoh4Dty3NREUkjwRV0nNvx82ATaPSx2AHIuKWhNRh9JFfk5W7A/CPflsG
kccNSnegZR0tcj/BodYZdZnHZqD/CNN8FfrNRjU5E3gpjpIJsad8Qmnzepe5
noD5Wy4IIv7rmOG+SRJQJXvsL4TMBS/iCd95424beCXPoWzDU1cSqhEGi6CT
h83d5gLwvT0b4I/WoLiKz5OSXA2AjglkbodUxdVGezwsoGfMLG3H0OetS+Bw
Y3Fp9SmeFxPgVvGuOIi6CeWWTEvgFbF//tPac7FZGjtmWuZSsilRIs9gJ95x
jDTC10LnzSFUavmM9IMdvJXbiRjAeWThEKkvOsi7aQCVn+ETXqBhvyTeJKGU
6w3BcnRbAZohqR8owPx52x0CQ4atgRR8S/y8w3fgZMBQGmiRDxPoHzzG0mPb
7uI9+cfL90w4Y6M0IdvqRYd6R5KV22/2DpCsvrhJcJZ9cx0fhN7Iz6RnjEYs
Arq3OYmS/BSx7X9s8YP+OvpLl05ZSd16NgTUeHhIdHoP2rz+N7+dB7MOrujZ
eBiCNWUJP2DMJmezVsB3Yro5Cbqt8ex1zmDkJfqyumUweRzysYg3KxNUui/l
Fb5rRrcQ3i9f3HvWrlVK7ZJwJ+CTlGRMtada3EtzXV3zgGLqXzZPZwbz4vW3
FtNqDXkIm8E3mCcvZLdcWG8oSvTO+wgNtyXkKkGUOlDSgMaLPTWBBunfYb33
ZxSKjq2BygnPS3vkfYDE/lt0u4GzNsL6/hGEG1952FYxOSvIX6d5vhWWbyVw
78do6sb1UevTZJDkmZiHpIOZtqHb/3tNSQyaP7CVpKmtDLc/tD6Yzo6gr4UG
vnI1zGQ7OvnIClWOnViXOqXEdOPhLrvLBiOBsZWURZEhh6TkTcWPWJu+HqHp
sTQzLOvD1rdipDMj9tQngg6y6oa8IgviP+Ni97KlLTQLMKVDKT27rBvQxn+p
/92UWeR5VZTbURy/ATaVZcCWQkJhYnEVniCnkINtj3U0H04oQfQ29m0pJ3cv
oM3vtO3as7GYGI5dXpMdAIMauhDAHFwMk71HJwC44i40LW7FK5X8lZLb03Q+
B/Mg8aT+9wCZ/stbPbtHfM9zurPrtimZcmjXbBWO6yODpFfG3Y9Cs2Zmjfz1
FND/QHnFc0Cm5kFz2g4FgcGtl3dgQIlZaymuFvjYIIfbodzGxeOIOuY1pDB8
xYSjz7oaULcyR9g5oF1VReLMFnPOor25/x/Y534gXjkJjz3ZJEmlaUexrmRB
UyL9iT6VoamVR2fJMqpsNVN7be0hzJCco2jNERHfEJlI4oYe1xEXVtDWbcru
B2ePaq5x/Miia8VF3XkUKRA9U+lE6fSPDBJwRYUsliBSWaiQb9Dh/7M2z2Sn
NRsiNFY2sL6TX0wq6UEDc9NrFNVaA/gB+ZEi2alaZeMDnwDYRRpalyB03RCK
F45AHM+F38q/6jH9t6k6AHfEg1Ua72x5DGNU2OR0PzipXjMtrqtxgnvp2h2s
t6bQA0XJvIbfkQHaB9KxfKOUyUVDGPtn7c7pwRRYF1dXYlqlogvPThYrU05F
FX+wGDRLnBp15BYCOi0CwEsSwjk/3bKBFqP9jfIIbUCuHyhccrM7il2rWTva
7b1Rn8kkQjPV7EbeESGcVDr9R8lPAW6pqg7v2opYjAjLujp2xi7cGKi/6umz
gZ5U7ffHlTzdde6CLy3qKnWZWrWSGlRYb7eQ2X5PLnbe1VawQZt74OvsuW5l
sTvWSnCPmlAATSgtw8qRY3jO4KUC7or5SHZPh5JamW3GUyRb/W9CgTMjUoxJ
2QGIYJYUuCz4LvwcmfzqjkR60JZQMWTS92XYIGaXrbUPRIxLeTyCMP8WcfKV
+SdbHIUsIIhwalpfGEFYRt9ONMZ8hn1Pg28YA3G2cxeqQ1AgWv2wT3soK9wR
nAtcHwr49AsbtgJhL/vFnToX/rZ6Q2t8lRCh8JxA8963Fa4454osg/LbPkWV
g0c38RfasXmxpDBChP5AfvPa/NDMQS/ZWedv0f0GjUSMXMI2byu+TGBHiZ+d
WWLSSqa97eQbHbVkXxOVOP+2GhocBAmyRDg8du4SiCrveySdbLcrLZSS0Rh7
ofXgdZQCn3fdEjTYg0Gs00Q6HmeoHAs2120gU3HEk6ZKkQA9UBSsQ+Qm/CRX
S6OIRdXEIm5NIF9cEHElGlXVRKiWGf4t3HG1tL4AW+8fMaWeTD/NGDL8Swf8
aHZ6WOkC2rXp+aQ2l8DvKoxMhFLXJfiZYvbPF1z2BXJV8rcYKv3qfPHZ0VDG
nIeYlyxjUoh1mnvy2om3QQgyF6yRcB2Ko1PwOpv+azih+K1TdXpM50oRW6HR
UuYmYUbLYd7kQ5+E/p+AaE01K/PqZ3ihYo9x8xYN8EqFyGHV9LsiCmohY9T6
cupwyDkPjelZCI0Q/OhZ8mTRPv2JQl0MTORbw03dQ+JGtmVC3gaWuHBJeBft
WCluniI/SDsjpq3PvLmYxz36/eg2/MpO57fJlnBYWwzcb7Xdhc6J9UExJPWf
ALZ87GRMIiM1t5VnJMZUAg/xNDefEpQd4rr7ypc0C3cVjOKiUPHIPy081Ylz
dfi18PU7J3RLfyBCVkMIjGDsPO/2dxTRHQXlnHIGtmJyM8mxk4aBvSPAsxrW
SfNAhOrrNSiI5fJBjjIuqF6tDFD+S0nOHNM1zPqEC81tdH4TB5Ps9mWMLE4f
6MIUJpfKvIFtgBbeVPce2a7fG3GkmJv/FjT9VzB4qZ/n168e0VPgNTfym8Fx
7fzEbdmveVgwBPIQLAUWhlP/VlONjwGQXl+G3JsuLKm9Z17dfAQzS7saDMYq
m6Yovu6qHMW1SCwppJgNxwv8NHTq9nB9nJfN/JLPtYreYkBoOoVSGYlKVYwi
K6ZefP8/c+jvaD15rdWSg3kReMsIdFfg397ce70DnlgImDn8u3gx3x8spXKs
62qLb7vZd1hcskS0IqcHztoJqq6WzHsYXt9tmmvbcW4Y0VhxjDKXqhjLFspP
3Ptyx/gxD0P37qQb0png1N8ufP/qbuIUUQllGmbohC9S+9RiyMLvox2bZrBa
z/80RYdfn+jyLhxVYwDhsUW4hrRzbethyIwLi1ABUYlPGIS8F81e5FsG7sC4
B0A0gNGdfhNNfGQIzpurQFOnitdgdTWVLYLLO7IOCDpgCvv8Es1mcCN9T7hc
0ivwHl1BpciKnmRK2ds60EhXtnwAa7cZIptvXAQ5YlFwMWMjHWrfjpe6Z6aE
ELX9JxBRtF/BdYRW91Y0hygwpyu4qi5TymcEntej9MmMCdKSVkPWySKxi7ww
0OOHh8Oy5JvnMfhSa1HgCY7xOmkpCEEX6zcq2NehH3GrCWwFK0jJQdUm/1iw
9eEDEHNlF4rSTxpI7N3SGZsVHCYEGL0HlK5hMZnOK1IrUL6MFDU8aOmPzGjy
9CayHY6cO7MMWGgGBbT2tFFqPsF5nc5/UxDijae+Axx9XTMqc7aJvM7UdGn1
4GCeUlnZbs/FxjQYUbbK+kM4C6mtVHeFIQjPV3btNT78NBoiM40Y+MeJtRhn
9LBDza4dRrClMGO9TK84yiSoxtsG1D286h5Zd8+bLUF3DkyRdOqtxdTh0AUa
Ix4/qQSIxLlaawkNVh37dHZBvQEhL6Hc7oi1QFOj3MykKQO5KyOSQqNHYQT6
WBaqOJH6txFPMwh9mal7t2COHUaRi+gFoNiWBei74075k/xVnOZz/dfUn/ii
ZcXLzNYBButl3HW+OYLM+dZxuTJ7lGtuJmSigHmxndhtM4YHz60S3BXpIgsd
Z6jN/3Q7cP3xnALykNOM2FpLoxcx5/XPd6jZnyD2HtOuqvlSqTZ7G0YeeJ7U
zz0IQbOEVQwjv9sMfztbZ66VfDz6mIqnKo+4xYv23MF8jW9Nqvc8d1hgrmRs
YHzAWONOlpTXnTiHYfhZ/wyM83mO2W/bsDbdIbKJkAODlDSZniY/wUEB8N67
K4R1HIPd3KTju2g+bSPWufgx87bjovNhlTU1TXUBwg3WmJ/JDNZH8Vxds+IO
T2myL2yJnxbUJG8WV9GX8E5byuV0fobfIOWvUYCu9g9eNyZ1RQHVsBFHJ39/
S8pQewR//hkyOMW2MoDfedWSOO3sqHQ6wWU6D79YeDlXW7+Z2luKloapQOQl
AWVT1U66xTT9MruissEscO99bYbvwqXB7vigvPQ+H+1G+urgKa1ksvjPStNk
vuqvK/iKtA2phfF6QON6CL4MZqC7mPdhyb/pp/QGLnvj+fwfBU+X3+LYc7Tz
ux+SuwA8yarLv0gWwCRJXgmyB1eaeNMcR4Z037p8+lvrq4YL/HxFu3fcdC16
ORatwOzVBzwYuWoUpjZUdpV5tLi7dsDXnDWoLJc77WQ3JQJ3RzOWrUBTvdn/
3jt5xAhVF5JQKuX+YcbuhVzxrOnn56EsOl2+VbrG7OzpJaJLBQ9VH5G1FsB5
sQaLo4JktFYxWVRW2xHNB/M1ZgA8bhYzwi72QgLXeNPblcdohVEgRoPwNTHa
YLtu3CK+r4hDTRVXeLxxQRAT0swbb6pTAVMQT0Lq71oJFKrZ3oszXFBMVKss
zf7Bdl9sJ9ejxyqGdYWZRq5Plmxh78Ik31SARcms7VfAgX9a0TaLPw+1696W
wPzukAum+UFX02IVO5PAPLUUYMQC8Ks4FPiWQoFYPHBflzkb9cbszMgWuujU
Chv7mu5xGmGn7S5Rn00PYyfsozIHvXoOr3q3qStPwe06JyFEdIDipLWosW4h
/rTiHPr5UYLrjkdwKySx/NnclkHEjrRJ7SF9DzJc/sKk69N91dY6okk5jY64
ft8ebQkKVX5XWQcdVjy1MH7UjR6XbStFmp6AgT+HqqHiOozd6/vBTWd1bLgh
1a1w0ozPJGxtHUiKkUrgrkxoKe9K8lOFekM9B695JPTLQcWj7a/kWkm1gceR
2Z+LbEvuEjWa+bbcu99EskuOOTJa9S5uIY2T90exlPUB1qM+r7meTx2Nkmt+
Hm1/4S4fHNFPtKji09Ji/s0YpcGeNEXh0r2SNIswRqUAktSsogGfpXz+aAs1
acfZXTe2b5EL/CqZ6x0OXNm19Qvd7LBRtR78Vx0atiWrXiES3PgaIoxxRpSX
91bEshLV/7NjqApkL67I7JtrdOZ963qQNWZLYWC3d+O1O66/X34DCEOYLOQ4
K8eC1djr6kUx5ixDlMsg1sIhWGqcyAf5PmfU3EN8eOFnfPBcgWulgU7sOR5Y
TOizgHeLxhnQD8qa/uTNy7/kI/CSq9GKMMbhoEyfV/22ETMZLdAcK2nvyYXy
Ypn+LyYrDg+FR9ReARziWX5pnCh/ikMlp0jget0zXFZn9s2R+CpVko13J3J7
HJgsvcS5zjc/3CJuSfse84AtSAYgaOPiSKxTCQGuXeklCFnuoVuLb/cVpkmC
iFAIr+EhMqBptVHovrE/AKD6/mNIVEF8rOMfCJYTWAH8hRVG1DAh6FsuawY/
hVrc3Hc/M9C0DXObIV9lkl+ZDtYXFoHyITtI9LBIJhso3dRXaj0rq4C484I5
GaLJgEcx5kNvRX0O/NSH7fVY+4j5hpXaNsATFywFduXxHFihawpc22jyIv92
lspylfPWMiquf9TYD2p8qNJeMPE6owNgILj110HO7CpcxG5HC5zHJw3RbZoG
wAQhaD2t4Vl8lB/fC+RfAEdAsMfmbHVfJoqgCoA8hojYjELGpV1n3//bFvpW
zNO09Be8rXOhLJ5lgl3O90jifoeK/0U7BmKfLOIgPIRHkzwaj685VcWHMw6s
qXE4ZdldBBUI3Dydf/et3tLRdiak8RzmiIrj7I6Ho1OtQ81/aLkwwCeLYBfe
WXthb1WM8CoHFtIl2oFVlVXgkZRyrXwFq+aPAxS8dEucJy1w4whA/CcnNA2V
RB1OUGrKTEspf6DoPRyBl6/jl408A/9LrxfYOMb/OI2gj9VGCJqs5DfhH+xX
drreCFVHR6RbVaNvNAt9gGLmu+hTMxIL4nLLJbGySAKqY4BHV6VnB+OpZKTr
YHAC6lPwaFMEWxw82VRUgzniPVROiED69V/EXar8fglLG1//6qIl6ZyKwbtX
hli2ZcsgyaU8RBNv+RRIGdur32/bJ2JsxvIuz9NaJFMiYFKvVJNiQ6s0jC58
Voff09TURXPDMabr08VVe8sMikNtbXcnpHUTAWilQcdoYzld6gjlsi+aP2Hw
twhkVcL/9L9aQHawgK5vjI3Lli/tcTeVcTpijBW9mSY2XaXypx7CeVsbUO08
cCSdU4cvdlYipkpwM0wBSX7oe8MUn00OgonPVWQVWaZIy4sCeeKBDGl8N1JT
fZDGZg2KfYFfrGOsObUmWPyJviyp7EUJ7gsTEzVsrOpNnJD9vj7ztyNog8q/
+98Q8bjZo19j7R4DuCakjEJ41TB76ZaI8WzXTyl+VRCQWIPDvadkgXbOuT1O
+mQrXuZr7YCJ+jF4qah+1H4DZkPLgGHzLRld+CbXlSC/KxvMuZZgQ4pCphqc
pYoiqkZLsazi8fDEvHd8EST7jPClocZYFLaDcylBlngXgHHHiSfOihIYVvFz
xro5IrFXmlfPiipVEL9G2X4Ctxo2O2pEK5ASQO1UVpu2WfTmGZSL8Y7LjfNm
uu+SMkCg2/GOZuI0kzLeINX//fZ0MEURMAfOTdKt4P3z+SAXiWG2V81dRSwV
rF/NStzej3J2PnnBrp3vwmA8y8i24HyC9VUM2kRRhgpr7iyXFZA1LAj4VjdJ
rjkCSiyFOBtkSGLzdocEH9de2SJaNpQgIg982q8h3K+bi4o3NN3i7Ix77Tvs
NPK4caw5AvZ3gmgVfmbwZZPun56xwNNoVWr7hTc/HM+QYOWCy3YrHOWf0yu/
LsMIAtj7pPlYJRcT90q3x7uvx831EUZzpZettXLlxGz4nWFWsey1Wdl+udcE
EGtsDNj4UCN0OcBwtL0Kd4vq3fdG4Eug5fN4VMQYXtRHU7SPADqH7w1CzawF
UsbwlZgEfldbCIy6VsEwXnVlUjXET9YK64Uipgy/PSvcYkg1BsKWd1RXvUh3
Jh4/iXIqgE4xtEwZPTGgsuTnEKOEobCnNKBKX7Zf9NWw64iUncuMt7YezABN
WkkSHQpnMKVMo60/ckJe+XU+XVQkI2OriYNM/Khcl+FYwdaVyNgvQc4HJOli
97pW6rpMQiEcWCeYh+A3rBw36d7QH2LXIzhgRc4MIIpe/yxlGkGB3Cd4NluJ
/xQzaxVpYUYRWRtJMz4ixBQkyK2vHc8ZcpYCLiomwFS7HomfjIWSAI1uKTdQ
kBk4e7IQY9dHsQhbcxJrQQHAF/oQFlnZ+h12bZWO63MxNN4RoVrU8v++D+bk
Y2VjXqUZFXk1n3JqBVbjb+/3ZPMh0uIuxMtFqzMWPQ8i3EsBI2QiYROCW576
oBcpncklwgTPegIyDGhJwZLKfDuXj02v5Yx4wl7GTN7qksHuRaUbFNxQBibm
49U3cZbEnIlJGTprpBLmPadUJWs7+U7SIq3mw2ZvibfkxMzYQeapwg3Ul7qs
fy1XBd4xyKxki87Y2xL097WidAxpX/Yqyy/Q2HKx6KjyQ16pn4j8zo9DeAyr
7lehtfpwCD99WXqcNsGoXsyNcdFYVfKBXAJCoxtxnDniIe9ArHuzU8QBv48e
90BPPkMr5s8Yolj3rwuOoAb/+QEQNHZJ9S7lhGwwWPGkkSQGJRuwwrwDJsal
1PxMELNV/ctJ4hczyTjnag5Q4583NH/5QsuE1m8f1OY0FEQSSRWY5cxeFpvc
WFygR0C81kTlpEgqqhgVGRT0FkRK66K2caDlIxUxI35ABsdMJGsr81jEYxDI
X89UG5QxaIyJsnVGQp596bz3OpGStrY9Cx8DXd31AO/kq1+WLXo+S895mylH
UXuAwFZld7MZtlFk+2udFBDTTFU7Y5heRenN1U2+Tk4L206Pc9yw3Ib6v9rk
rOOf9qb3hA0cxA1Blm8YJpValxUVmA++ihm4MY1QMaIYXCMToM3/9OtbcpxP
Ds6Klr0TZB8kg7Ftt9X2qzMdEx+E6w08/fRdtVEh1mZGCf4d+IRnf6Mm/lus
r3fdT9UjYtFM5nkMv9h7YJXWlTtK677Ea7i1Ss9kxBSwVLxhJaQU1PPiCnnn
TjNYUvA/uOjEGCpgfbkKZLSj/maPFePWYoSYJftXrfCXLYM09JlHcu3BX9vD
75oJNiu5p1CQsuvXHooa4AtArFAv486oVdDKWZnCsXqQmkCyNgRl3RwDCAuq
U1glB4kAAzEJi9MZNi8+PUctKZaJCU5lMRz7q236NTwN3sinB0IEg16uyDSS
41lzczTVuWzB28V5fEd2b2J4fOOeTFI20nnwzotlbvWScERLacl+Lki4MmbD
U0mK+ge3CdhGnD2NuVnqQIlBsUP+BazPCk7L1RgVveov1lc3RsVEjmj8jCkZ
hMKIwxiZysKx+OipGxSHB7mCIr0E05FlKDlnj2XbLLgPpQOCa0kY5UaM03m3
T+vdspUfwZbJV+pdo6pOp/5DBR87hEkVBCHRsiv5rHfDsiK915+9Nq2ULcdF
PzQeyfxBGjEamVJzS2SNIkyDgtoSghdkJg75Rhi0LqedXmPIwGfnayVpW8HO
0k709w1oG2wUuAhjVXff2OwqE56KNqc4w99TSwy4hFwvJjBvqqWumJzy505b
MClpm4JYH3XQejjFnrEh3wDVfIGsid4iGCmYPPueBswsfPH/T5Fs6F0ZDdY6
olxpq6hOawSuUCiuAea2t+HR56jya2qUUSpneZKgYB/TLfPq7iv14k424Tuz
BlS7lebwt7IAm3q8dCWXcadaJVXYYtSK9fByg3d4LHmHXYVAVfnjqz0Zrhxj
PTAIYERmY0M6/5WZ+Y/dcEfdm0ZREVpx4i5virb/LcGcK4QuRxOCdOYlu3kj
VZWYc8NI2xGimmtoWX3UgwepK7Jt9SgA3NeV3l0SzJyIzuHMAmxtjkle/Cee
78yvHD7trHBdeGgT7pSm9N3T+ZDFJcIvf3ULbTAxUtirtp7YbfmcBxKzYw5I
Du4VOPiyvZYtiprSpSTsTfUTyst1+uSBMwjJtIm5DCnUy39KvUgSOmw3sOyT
SQ/7UICovzNl4brY3AMPnkpmjzMIPM6daL/U21B8RB/nj7hlWYynLvAZn8gR
PIRqZT2goQiXZJ8HInO9SsSDIzTDUl7lH1tZoSkLDpxrAzc/2QUie/SCXH4T
Dc6b4I6xDTvphHioRZeHbVH3hyb/8af5ZUBhkGj4Z64MCDgv+w9p3VTau9Ma
ELnCUz0z5xxgN3O4p6tGWclslrkYqMvpF+UOjNmrObJ6m0EIXqZMB/P4cKlc
rZeGyQppIj2fsdqgUqN2fTKQhY13kxIa/xyKzL2fMsN67sch2b+3ftzrBjtR
FNyfje7tk4ur+frGEi89dmO300Qc9BOOfnZX7EGu0rdMAB3TFmSFuvVFtCzR
VT8nVBReo6/q1J007EpRFnjiZg50+xZfo/Hfnn6DIRmsQWbuF88nuB27mR3z
FziYKo1d2TXaKjSTEheYpXK/TJaQVxZsYDfuSj6F0/q+DLrw4s5Vado8mqkl
dkAmtJA1hTNRETFEUU3b3BAOD9MIiTn4TAzlK+EuIRfgF5QILaWRKEXDCT8L
6tEVj2yYL64fnadSHl4H2F2LMjho6FyRkbuc+MHwR8v5+uGhNqqCCpu36erW
wrPbFlud6gU5bEkBIyUMQ5GzZsXyyUJO5pokNu9pYmWnbfaUwYPNyB5vfKQI
nugFbdT9+d9dkfNDqSnc6rDsdsyopVkRQix6SZL71Ml+RZLDppf5+ASgFn7T
lu/bxd7TolNQVJr+v7UlPpZVGnbW1wujUdp54ozxT0uzmSngOWHuAoj72rYl
x5j1SspESy8mYGsDC9liX+LSxf1+OE/HRciX0kG31YSBTKpySeP4KCFDklc2
TzhCdQFSguBAUNHVF7h2kWrioVguDFvbr7xZcLfVtowq0W94UjePal4blyjS
XghEwgKDeZddgcXK08G8V0c8seyW2ZVh8TvJE3OOV0boJI6sTBwl6WZSWGvn
UC3aLqBXwvOoVTrUHmO8GqEucz+gYuON3BB9NiCQT+pU7Zim4mhD9FXVFjLN
/ozM4LSvkBRzppaBlfDIciFNp8NE9FGFv9oSwZE0wZTTe7hbhUvz3G7LRj92
9L9uGlbVKSo22uybQ7FRmWaMOt6nRj7KcTOenyppI+lgY76oWeV9G3VBvoPr
tHcBfpWjAhycwfKNiNB90OA7P001WeK3vryPHDnjRucIMG1Cj2KOSRxyDEH/
CCqCddcmNHVRLERJh1T+BoqQLGPrz2LjIO2Q/fCzEfSr1xbluJG9tRXhIbyi
3iVQSFFG/pgozw726adEIxoL/6lJhgVn4rzaY58M51R1+w6obx2KF5IZXTfd
SzMjK3HnTB6ZiOOASWRGlL3coEl1vXITqoKQDaV5Ktk52gRn46SqNUk9wXnA
ro/d8P+hZdk/otAOLW/Ob44syOCkzBKSVxnKoo8rl7uwcv2EIF1Ccp5DjHI+
tnIVeYNx2PTtgLjST4aoEiB4kF59tKyKSCOSrrxPScY3Kk8s+mjpV7j+b4EH
ZB94ns8DC5LSuRDF+YSHo5Ng9VLYy8E8Fo8GONOB5P0PZW4evgOpVaCbbqE9
Z1o4702Gjit51nlu6NJdQAmhGzdEei3U/HBoAOS2LMg48iihdSirg683oxA/
qERsxqYvMpmu8tdzziT4BrdHbrFN/agOE+as4u9KEsNWp3UKuzTW4rqO08pq
j9mmVhJA6JunrFBRzsT8kfb3CGdvTb41QhIzioab2DdOAhk9qr7TW9nkWLKO
zXKuIF0B1d1FhTYO8SEJp8uaBpCga66FFgCmnu897oDJ0m0gYqg9rjvAJq59
99yNyRR6426Kw9Jl8l8bwBYK3MnwWZ6zYFC4i+/Y/BSENBTj2fEfoB1Fn3aP
VxTaVq9+gUwhvOcS+AkTbXJmmymn6JlDbgFlBDwMtg++Zp1EUTqrruBumqUR
CPeTVejcPEiwA3itTTvlbn1d5dY2VMvokJ27NygcMKv9GYZGa10gSwZp6H+m
sCQOpU/bSf7O19Psc7SJjea6laFS92DGRc1QunRo/Mp+SRTprRG552B4QJx2
+zZgUu+PN4qm/gls6ArJRMRwCMtYF8RECHnYqnfsHXQhVpX1rEPiyP5BUyjx
+ZDuHKfOK9dZ21EJ9eC6XTaeZD2QeqVB1jOUiULuZUHoWgbMtllmmEiucBDL
FDTgkImGZoPqZLQmjPappFszEZuINRhlAreQaALDwWAOWiFZ/9NuVJVIm4vm
no3ozeIPp07L33dXLLl3IK/GQ0pgTT4vJkxogZyniPzKAz5oF7YUXaWiZu8q
M/5WHRy7UuahnbRkUPNz1WxXj0a9qY50SQrmrjdlS5qH7oZlqhXzkaNOWXTQ
YXX4WIUDOrtWJ3pNR6Yh3nq/PZ0a4soAekaDDlzh9P9nM7HyY6i9UZV0ezt2
mzUV6jWDje9Zus6pcQLmO/VYwYcztglPwzNaV/emnE86Ae4SNSuRg59+895N
EPdbBgelX3nQ7CMFqURm2/L4fqQhp0ykUBqfm5dhWm+La5OS7fDLWHXF9aiH
Opqf3EGfl/1PGST/CCfYR5X+I1OOhmcjNSJlaUYPPT9tg2cGRfQNsL4pXBdx
x0HCiwTTWRWvbt0LrT920dnXgq/LYFlrjd4JzwR0n0b9WTi/S1mAdh+N05Gg
XntpmDwQKPwbVMf4gGbgHbcVr1/a0GngpITc6C8TmbHwjcUVZqVAiertUwjd
s3U8Ni25OoLL6uymxDOFioy09S+M9clGU8r2Q/aAYT3drfYOdZH5GiFriynf
5cI+i2c4BvG7VheKalh8q5vlpv3mnNeMnXkB9e5jE6tfq8sKmORJL4lvMvQ5
5vx+GWTi6rDsnEZdRwjsVbZJyCIGmHI23Yymn7o12SLcBDR6+yGcPKo2uvAJ
Oy7OJfdarUouSdyMKVAnQtRvKwz7915S2VYMvxgbuIfFMZTRSlh6XtIKQ/of
b7vBbXr87MENebPh9gG9ungztadTidDVtnBNznejfKRo667HoWHM4zsnERqS
SzIaeTKvLzT1821ucjh9G/grcjiEh8df80okS0xZYQnaV6CTpjpItj20Ehko
UdYoGH4rNnDuIrKXQfZFtnxNJedYS9Dnc21x78STAD2KKV2fwaRMNbchUnre
2aXf+7scJsf7mACk2UZpwI0FuPfVqfh9y+zYEzTgkvsNjPnxZ1W+MGVLE7E2
m979w7qF728hvsRrJ7/qVNANZtiBm9wrB/fxcfgSgJ4KtzM6ZXtWvrFV8ZCr
bJH0RNHYWXDCcJzb+RFQWmn3dfYRx6AW68FASXwPxSGd810oW9tq/3LpGvv1
8/49HFhy0+FJ3S3tu4XfMpUDXBne4pDOvW+RNN9phmnC3U1u2bkwHU9unw5T
zlHjKPxzOXfchjGLhNfn37ER/BEjuaH3jcgHO/ADjEsQEbzjOvo4svZ7UQUn
++cOF/bh1Di1OEdPh1cw77aiInBbqLViHOpZ0l1b4b+IvWATCYIqHtsAb4A8
k+p+PHqDtzmKdC9nn5qD0BtoFZCqTVL4tzZTQTCM4cuTOmTygELKkIrTw20Y
mBh7Vb9JAb+ImXEGr2JHuDyHmsJ++WhXJ0+1JaamXOutUhjkZBiVT9k1Jcj2
x8TfZ3qRKUBd1UMmQVBfeqEOBElHAsxaI4TVtaaJEw0ut0q9Tq/bR0iA/C3V
1yAHc1tKZ88DP4cFp2YpWrGv8vhtvbK9ShqAklY1NpJp7SKJj8IsFVjE9QZY
CGrUqgC0HHysbiJNpXVri4sVTWApSSxMajHO8ez8iE+5jjLUH1CMDKkBkUuT
y7X4tTxlkDLcUbK2KlpTsyoc+IZ3Wb4RAvIZclVORttldFuojIo6FDANre5G
g85akXmD8y9eihEkiy9CU07oqkV5j7H6EkWqlRkpWySCGNbV1NCK8KD2oldS
AkSKwZlX4U9FrcamFSzhcTEJMgzU8hxpJJq2snFbdWiEvZpubWbboxEFMU47
W8ve8Si5BFEpi01FnO44e/oATTOIbA9My+4oCRSsJzIOqAP2JKO1F4KYja9m
ru9lZZvtbrYW5RjkpUNUPQDVZYQewk6wHxYLLhf+5Az8gG/2OT7nK6spu5do
mZLccSn3ciChQmJv19qKmY/qTvSVlhZ0OpQ3Jbk4KsP5i4PYVzxN7XPm6VPw
wme9D8URWxgqvTVO29prk8r/RnlAg9gY+CVU/MmHGp9dQ7uZe4Pj5WHd+trI
DNVUxgQQgE5NeXhKoxXRAIXROME2ViqDjAarW8DaO3MWc11aPBfEzTUcdrIW
P0kHtNRonb4/d3c6TrOtdoiDmgn5fh2SXCl0V7il+sc9Hu8AZgfIkOMuVZKb
RgjOWuYokdyPNB1PE2dUGwzZ+rkXV2HPoDhWX2UBCj7C4pe0eVX6BqNyygCv
sbtZzRhTt2Oi/ndZwLNLc7Imkj4Ab6X/ZfXaxsiTMr6g6Ih7WJ0kKUOA8eGt
gh3Mo8imgQJ8Y9hCzSUvyIsav45GMGZldCWvq1F+4Z2uxCQaA/Ro+vpgFWAw
2CTzZsfYkgZmwVi0h2WhSUJGgw66A3VUE+Ko1WdEB+BxfebOhNlZzshpJ71J
/ehU/50HlvNQiTgwQJ8FdhgxVVQN4Wlv5jvQ6HSY9RXXfjVXO1cu3b1J2Hx+
GgZBUfhx7TVOa3ef48F7S0oWV3fjpURIRxXMawqV5xk269jatDci3Ujvjucq
oVmDkbTV9/x7ATt31GpeS6pPb3xMrKXhmYQmRU2zUgHsyShAuLsRS+rYTSKW
r9K9T9epaQJuDtGSY4cvDpmiLxPeNiIvpVf2zZoIfbHkT8Np5ADVh4ivNd6c
YtTtc3IlQd0fcgfAgtIbhzzn+XlJGm+NCbjZ8PIiWVZ07iZVPQAfCD144FE6
frmeBUQrcP/a8z+BJgU27Drl3xSHfEOqm2kBgMAZHA/uqCXf3tQDYX9zFP/A
Bs+3yeox8zF3DSo+0OEBLSUe6ZGsQoCA6KHcs26ASZin33aChLEaxasNNwwZ
v/tX/lO7OgxBoTuoA84EpmxDGPvCE5czrufgXHUwoTWZTl6nY4n0qCJPjjHu
CA86TVQogqVjmcYz+J0apUbbrEJah+j7T4mdv4QShd3Blb8Nm34S2T8KT+pr
YKJZqDFVcbTBWA1Jzrt52Etvisvds2877Z04dKXKHO06xx6F8PzhJJs3i3ry
cpQ4gGkXFFjqrJCKz2ugn2xilmM5cvreE042eURT+l5OyUvOykFVVDskbcoh
kPpPuVd4fC4/MDsf2HwW6AEQ6rc+tFMaTOBrOJYN/eiD1uVmKZZpBonnTA7y
rKThRx4f1p2eLk1vMP9cUb3tsIGdG/V3vZr4xrmJSR5UTV2gpp8FSoBTEc4p
mq1rjrUijlNr42A5kNthfZR3iOmFkIkTqKqtQ6gx+bBnu2mShAgBqMiQ4/Ge
bakPX5RtNXNO7Zb30kT1n7QBKhw4F4VVKLvGA3Epy0GZP5O9L0F1EECAcSgC
nNVhr9DAKMpvsSGVkfX4Zhddpl4Bjv6L6skXEPz3D42a0q7u9Nh/k0bD1u6Q
Rt4kgebI8s42CfqxYNpNPhgdEGjHD4ify5YXnjdgeSzga13GjZ8iGcOxsXlc
somncgW9NugaWplWQlnKCpRUUD1gek/m2DNLLPjC8Wq2jShXlM9nNA8HGnNx
UgVA2nOuEItrgrZ5PWoYsWSyohcf43MY5xhJhaMF0M0myIAweRJcer+hJUKg
SEQ3Wmplz3PO+J5+LWwmPF1pwRgD22hegTvYl73TK67xdHGj0sBEJrtji3uN
BAdmCucQ0PxV313ZNkya3mJ/4h1/Hh/Ql7cJMsFkTGbJMwFpqNtGTdGmyHeo
vUgy1utC49HoERymKSOXobCnhtl+2zQkko1kdgS4u2ukiP/J8zqFeCjDMv1X
Vx+PCVHZisBtCHZ95ZiB7depdy5zp5B1Rkpsb4wTsp0828Noq90fBE/U3VaF
dMydENMDh97KpsvBqccfiXWp/aDPnzYrNvOVhpL7HjN8TkAf0tIK2iKzG11J
Q37wAvQSiTSNs6ZjuitWPm1VyIMkqLemo89krWWCPmVqVMYmPSqopVbSzFd9
g9XfMP6ySNuTjz+odAJ+moBjQsdO7ND+3AD1wjXkDoL94VEcQXLrUtccq9lc
1PphXRoEn9SBOc2c8mFtfOUe00qqUAy0U42cCdUWuXjl0IueK3T9j1hHO3pB
OkZ3y7/hjfXWv4Xq5x4P9BKXYOcOeiUWTT4SsC2Fk390NjKZK3b9RZMRoCuE
i1vlt8aIpcxj1bfRiAyZWQmgc9AkuBaDAn15hCLkS45XLDzXKoF54KoyzxBx
ZVcxhdkST1+cEhXNlGZ8CFuppujTzdZBFPMxD/PESiUceEp3LIWWQS05NlWM
ESaBoS7IWPwehOReiRdHBcPg/UlHrq5Ur+VXyxZFYUjDExx4IbbR+ph+JuCo
MKbviz1+jTVRtNfaxxI8Bc+Nr+0v0WCupO9278THgJaB6Q3mP6U/I+QLwvZ9
tOsf8HcngvmrLYEh+t9ZbY3rKnWd4vHH/DYCBsuVZKpMnyXQj8UC2nJGJHFI
9PJgtzXvWwRH+5pIWO0tl6bEX1LR9GXRoxbpwYLrJI9AtAauOSzuAGZTu8TH
94c3PKNsRCCjqXokn+5QAm9PBYicFq/ANxkjwn/PMQejAn7NYG3+vk5bL9P2
1pkg3+gAu/PXaOV5ntF49hB/jky+qGQfiLDOzEaWJC4/EDvzp9EDcBkhk7c2
AHEYUJAm/035w5mZ5Wno+KjJA076P+dUJBTM3NH8EQvxLrkW2K2oiZ4I6k/Y
uc9h7qHqDcNv33mFkXEfcb3tZz/FfYoW0m4G8RoBnTjX0C36HZ07EDyoVupU
xkBiwhT7vEfWxIRG3yW+1//h8GXei0T03cE/zsXCwsZMxt8YY73zlFF4A1ic
NiMWSWE/4pCNtUFiJ+6HQHo8RgZtxGwflSaQ4fYHIfjpX9+UGl1DRAXb9gEm
8P3r7ynzusYtSNcN+VzB2ZxumEd/Xjm02mNDX8gidA8gKbSyANmHX/x/iG6A
YNJz99ZxJeA6gtJtTFslMFieFxXQTM9iAXyN23pQ6/tTun3PxU5UdrBf0ArL
z+40ZXM6kBTVuTGJdoqfErK7RnrB/yc/iSrLv0LdOwRpWI6vmwen5I8VvlZV
aL94Pqqnv/5imkvtcTKhgyPxm+RJdAEVXkvRbGFoPKAu4aplZsWk4nHEkHfE
r/Z2jTFfgWROrt7FQhkwYYAukJ/raZdQedGIfZ4j2yQKMjsTBf4cqVITdxr3
SHS9OfGPwcrWNm/spX98Hl/qyFAd7rz+eXAizimReFLoeMhCNmwYoGjbfOmF
Sfojl+iw74E6xrQBLmo6+69nC5RtDitfJMnoEO9PnWN37zjfB6AhMilFBytF
+yuBs8rjm2oMk9iXuAiahNqbs/76toIu2SQ/ukj3AThIR5ETlk0zQRD5Tzv/
oWS6kWMkd3Dho8rgERMI0IwtxEbnc6mXgc9qY+1c1ACZGs6u+2zTcclhM6MN
TQRLeWLBxMrsnbhalYefz7NbXIt5jP01MpoIW/IADla9L1WfrSUUi119TT1V
ZyxYyORenkfgjiYBfvIB+rJPy2woEXgYJ7AIHISdJlyV9Q5rPGqlM+GWw7s4
IxlnL+47ZhV4/bK/j3p45GevHv+GPo1J6ARvFFKmPXWNSxY4Kz195geNPOL/
wL5gpTp5pn36TcMqRd9sOFeqF0e3Q4dj0YaKgWwdUKNZqlcLiXT0hDLu+xDY
CC4ifoCZkrLZLCh/8ZXAXORfVnwrvpNCBf7jkOV4yG1rMIW0Wiy7SqYLZMT4
ZheJeV82SLv/LYDf1k6VF0eidt16R8fyvIT+fClVYrkk7+28XCSezqin5ApH
T/R5Tr6rmVbAh1cirSFvMnkWbuGZ2eFsefSwkq+XViOkd+UUNpojfY5oOSTs
mBMbJh/dvfFiQ8ORfUHcwqNgbEPg+/3tQE6SaPduYk8m6KlKTzW8yNcvR2QE
MSdkilSIZhQqWGPyOJGWorHZ9VjXinyaBtdoGveiINDV93tJKNpPk2+PicRo
NXhYzOIwj0Ehs89c2woXovEYCLnqa8//7Cf5/8mdUG0hJvmkCEebms4he3Ro
YcjsSqIU/073c7yQKHRhYrFMU+Q6wKPv92L/dZGp/zPeNaIMpMuvUM0iIYaG
WzfV1VTagf/nnVhwANewGo3lnA5rQjH44JahNNKieP4SebrMx4Q4RyyPtW0n
QBX/hRj+m3JmUOiL52Q6Hx8bEpdIYkGRa+xT2Iyfag9PLCmHPZKtP9vphz39
om00HNxZ7PSqXKMy0FG97Mem7eiYn1OvUVbZHKa2Uis4CucUfazsnjKxPrF5
SbTapvg7EeATqGPGSJ0gum5KkxjiixV95Ng1+zB0542yTfF22+QfN04Vxjzq
SXKQ7NU33VUZCmRA4V4/yO3TXQOCMhGHlfs0ab5I354kxO+al/nWWfiP0bpL
+9XKU3HbQIWabbXi/C1IQzy+kJzOdhtysAKZ3p41L9fNkETwFbYY5eqcRtEa
6m/D/V7DwR01caqhX2h/P9FoPRv8hQOlYHhRFZdXTfDOzZyVtCS0jBoRAFbA
BGnDGUNhl3RCCI3vwIB3G4n0fotfyvcc86jWLXXLNLp0TlqNaPm7bztQwSR8
vWV59QKGEC6uZv9988UxHDhF2eWKP63tMJrlwq41lKWF88a2fa3ttO2VCoiu
/aCX/kMrxQLf2mZ1gB0MB/eMSqT3fu58hcvV75XGqJM/tbNqhvqxT5cCM480
3xHeuLqIjbMb/AMgAbFsj8zn7Zfz2Cz9j03e5/1tDjxkJQOo6VeVWnitb/aX
xMue5lPbPljnwmlTor6nKV79Xkh8D20LRtGXZDbFuRtEZHFzSty89BRIRP9N
Ty0xTcts77fkPOOT0Kknt3SID9kwMYy8BC8yoJes4eau2UKfqmChjBMVc46+
SrOO4gKM+7ZHodm9tdcuXy0zmATlusAJZVzyTSxN0/gCNaezdzlxRiaRPB4h
5KWM0bZQzyGZHH1GrIoWnHJM4LKoBlPk+pUxnMcSGoEJ+pC542SlTsaQWxN9
6QwhBNBP8qoswdLw22hFVh4KtjvZMcedIqri2A3ZhKAXCh3HY/A4qDlFLOlk
FEYXwEUO1bKFtjsTKZsI26NGj5eOC6I236G4QEJiSh1RRx7ENxLH/DZ4HcPU
XgbMWtivc5A83AxSZu2QtjfwEc1sV66MbM7ZgUTa7zObM9uixCwUNg9MXBM4
nqP4D43UAsvOvYhlfF2HwzNg/J7oBLlosvPLRPyE0UXLbbVxSl3J612w7dra
ZBRc5H3FqST57RYwiHTml+2TOWxQ9PhWohAwamsjuWUUQPEh1p19j5F27IIc
keZuixZN2SiK8G906az+6bYBsA0yerOZasoWRfwVzdGKbiHZ5KP90/qUSwKW
TC9U/t9JMdwLyY3mv9DV8rMcJgaXthdgQ1yWsSCdpNuu7u3IjBFLSgwWFQRa
vAf5u6cZ9Au3o+ZAqwgec8nxKOpydV7TyGJJrvfrfv5OXX6a1HOS1LOTpCWi
iUfzL6yMaUzasTc1poHA6VqpEB3wKWEGNDHJ8l14PY5i8RU/AlGwBUrvOb/o
tQXTic2rtbIvFbPcxF5UZmGQP0OzIB0AlF6BkMniHtVFbfM7MLWznJnsty1S
hEPTaFi7oami7aDLwaDac25hzo8tgkbNyWCMW/waRaOZMR+Lj1L8gS81CY77
M/9xq+cedrKDp3I0q5csBnQBkNCMjdvxEDzDBmy3HoxBr8/jxw6V0pIog1F1
BLCa9NUfS4YOtHNfKkNlLjTQ+Dh+bq5LcXbuCZJknMU3sQHXxUSFLYfebn7Z
u5tl5X/oXXZGYsIVUBaowaecVyUQpB/USPJvBjuVMqDmgVOB3T1278A4rneN
RWgeMjdXU/Fzmd/GsZ1sXuhp3Gq0iHEbAo7kvfboCY4rNGP/QWmQtUeompTn
05ciAaJE+dd+GW5acRuPahI4tDkxbUoUZ8HesxsQbB0U4A+2FzBlwMrfft2b
QJu67vP9TS5DoHlKTEu828J90Ns+H4Gzq8Zi/vNhVqj9lZBixoFJ/YshDxLt
RFS+N7ZA+cm5z2Ozwb2y5HSnd+UKgG7DUQv0KUyqNYGeBtx+ehtwWXhOStNi
VaP8N2a83tSr0AOLxgEy0ZNFH4tw8vWfsxqb+gNok4Y+cvBqvc3hZwqAowR8
tqhu60PPBENaKhWYKJ1HjVbGYYF5a34OLWQLCbxiI5xb3oKlcm5G5fLdsxkH
mmCg7zzJOUeJeFQma1w/F+hR15rpO2keL091hDWSmBE96ZpVqGm794mr/TMm
hcuFrxY50reumVqOESJEdLCzkauYX//w+cqJut3xcgY6Vqs0TU5ZwFsRR2gW
pduLVpOFaTDSMcb+03QgSZwwLO44VlEwyP/ytE9BnBMUJan1teEJR8Ljq9WG
geFSp0Ru836KNIoICsEF0R+SjgEpD343e199SuOKduuxPsZwwScwDfUTpcuL
roiGrDdtXzcqfdCDJP0RozbNUUXnj6bR/DB3zIDUsySBVSENebEw8iwhgSMq
kPfSGDmd0ikqRshJktZdqiejG6eNyas0YAQYcNjmHlFHVOSELjWUmmzBSkzT
9vuG33ltn2lA9kJIyRIgCRT55Pwm3XhSu4jFnsgxe8tvELjMVe1fw58MdGLE
nw15L79iOaO9PysX/eqr7HJqpNAufYOG/Dufdlsv3VAuuaqNz4B8ousKi3ZS
0irJK99QEYRUOjd439VUj8dTyPXhq4I12ia94OdaqIT6zT4Li5cE8bjVzEZu
+5ciqjI2FRNYrNHLyuMg6YtFhU1fC49hRyUhgmXl6rCC4ISWMWQfFIqJ8Vav
oyPLY/mVzIDlKWUetjwpULn6k9ZcMNQE4cBQSfXSh5Jdb6sqdWCMkLIfEKWz
/Ck4q/CQYnLCJbxnOMN536cJz3kWD9VFkyrY1HkOO5q6P1NzH5Dx4zTbw13M
hItMEmUe8mJvHAhdTGsZ5BJlpk4pveUSGwfQ/H6xf5UQ1WkKKr8xo6DoqqK1
7WiURbKEEO86jiHkhQQgej/mmYxWFkwO9rsMae0IooR+Iye/WFZWInaV08t8
LAXdD1MGZ6GPSzPA4lISvzzk8All0604g+xnKd8T/6Hev1W9v3P9KDv7TMR3
iNffhP0UtEMJjeR42PO82+te0CL4zYokhZg9QuMjw2DzQpMdGifvz5ngMUbY
SruwtTozIH7dL5q476w1qrlyQ1ETlMZG5i2DxIWL8eedpMXGkrVvl8mYcCK6
pRefZG3EvvPeNLkwdbjEL2M0emxdBN+Gl5WMSyq0FRou51jtdf/tZxjXV3Yy
oMQeAxleMMC8Ynr2+uEq2Nk7txF/u4oBiKe4cywNgTr7iIb9ZlNwq0u5UuMg
pfM8pNaU1nCzww+7yWqCPGJ3WAxGTJdNwE/R9/c7NpQu22+Bg6Hh0bm4Szmt
9BEt/FezqKm6UqID0Xm4U84CxlVUEJNyjFXJO0jp1/bMIE79X22XDzrRs0iO
EzicNYHXahHl3aSlMRS2BQ+1V/btOQGIdyLVE+pNWy9p1QyhwaAFww1hfM9/
ZMHGdkrUusxSeRbgpe0h2WRU+CXWjLFPgmkgPfh8K8yFWjs/l7El17SZ/eZd
RCnwB2vPp2elw1ej4GC5HgI8flR5GikxW/K3P5e+TLqrOD83cfHCr8YKV9WM
oAp2y7h7j7UJBRgc6UFkBsHMJcJfAOMI4HoVY9mjXy/NlPWt+XjA3kqrZFiP
pIyYD+AgrKB4dD04tXVFlHNhS9bq3N4LbkKonbn2ldbBIjt1hpVHb1GRljqp
K5HLlVG29VT02xP0xPcIEi7rX4gKT0TSBUFPJBXinNRGCpm4JIDJBuCEL7Mq
F3wtLyPbTxLpYbUmiHGFjyO9/3Os+3lNRGpBKFXQ3SDYLklMsSIH9XY5p4pU
9DzQXS6A+h2i4Wvgawlfd8VCHarcYsDX/nwQRMU7FmmCqpKa5KURX6rdHd7Y
WObj9EC1nOdhcXo78281030pLOmvLSme0HOAOK5eyQjork7D/0Mw9umJvHhu
xMnQXhe/NakKy/F/x8qB+arvB6h4um4zjoeHEXLvgHMJyvp4MDpYnQUaa5WS
vnw6B+/XJeLQyGihOcfktSlXXaMiEsN4hkzJIIRa1euFqZKtNffTm0aw3f2P
EIYkZ1rUwrD8I7l70aKXs2/LHVQh87NGDFDnlkMT3gyY8CQO+BtL527HJEcN
t+AZ0/SImAycpghsR1yi/2keHbo0gVugv5giB2Dse0dQ+6HH4PV4bmJX1HPF
sfWx4r5ZQl87eFJetXPJb6geQ2LZKZKl3VPeM3x3j8GabyR/UwU/rRIKutBj
CuZrUkGqHicsJ3vsI8ncwHPKk22tS94FeAbOPYDd1J+XEwKHmLq4Ff44DKOE
5CtAkGTVCXUW2v6rKAvmb8VluyZZeBfJEF7p00ntyLEV/vV8rg7IxKmvvmwA
PbxE46SfBgwg1S3PW1pgkip1hEn76aO9pjqPBwzcL4scRTvJNgR0NKT/QBLY
oPtb0HR2qELtb8xid31M5KuDDlfJWLk05isc1Jg36xWzs1K6xss9s064jyld
BLH8aYFro0C6k4Vr7WxzlMfxN2RU04YOK3iXGEG0O1BhxxPaY4VvTDcxjLhd
wNN3W4ZFYII+WfOTs/fzQcprKXS4LuH71qA62JTrc6SxcyCcHnmuGpU1VbfD
p0znlLEiVuG1QOhgxKqm8rHVLYIimczvc3GxsRfEq2VD9UpMCYZ44bkVZXpa
SoPD8bzPXn4jpsbcdKkygGP2cT9aSAfijmGpoIaA5tAEeYVRGSAO/oTOZb8w
Y8McrMoeJo7tvaDHwWWBJ4eLeq8Gd/SfucxzuZkpYa52q2k6L6wMPg/6r8Iz
3ukXye39JyzwD1pAEKwVIcXlc4n9XwclhT9NW+raQVkIlhi1MH5fh9aUNRUc
uMTLX0PxeoWAmODIvMuz9D5Yp43nEcdbDvjTSDnubDphZliLYWmlO8+98wCX
KaB2lXJ7akxOBK5+usA0td0gVFPNcABPsBZ4A5DOxfL6YqQL9MbklA7zfU7I
kL2JLEdQpAuvRmf53UeG2NaECQ7xHTkJdRpFLnOCdejvsfO456kZGcSukX1C
qpJzAUJ4qAk6AlFNwTQEn9jf14bvAjFB9CoTaH3jTEnxOIkLwUmcrHHQ3aci
EQAOBwO6Es5W0qJ0QhFIcAbHAzcaD57O2uwxuRR8IdrRboLK0s1HnLbCALqC
3Pjs0lrog7wUEktiZQiexqY676vZxz10pVQswST72PNua5gHzWvRMtJCCBjj
HiANOC3t9XlDmJZVB8ITEqJ4ywjA5wB2Cu3KdN/qRvLaMkOTGkDTAH/XLxd6
apHpn+FOVXg8JWITH5B2Vbok/DP+9XrovkVjT21Je2Hc+IHHlxNfohsSUX13
C36NvbVVRgyQWHg43XvRUeuNcHvWO5SFlBAVHxpfHjrkI4YS0AYQa1dF3C83
jC/MPYpQZ4mrr+/QabO0C3AK5EP6URK9m2zu2+sV52DkCP7QA5eFdjNwhElP
yaQFxmKiNd9N6UOgyPMu49T+7cHT053CkLZgfM6CT93Lmt9Nkr5wBE2YNEN+
09FB32F5rRqZt0OI7yphdFzNmZMpw5GgiY7/KQw6qGr1iy0FXOoxwG8XFxYP
FhnLEAJ4lqTD4xfZFn2rj74sXjQGM9SsdhnF++KzVrXKwPu82Ak5+FDyMW41
53+R6b4MkUdrYErKR1/NYMvy2SNiM8rN7haN3AoO/gvyFhBPRsQDTdo+WHN7
AXdDIsLAnWrk0g4W9Mm2LIGEarBHmggiX7yIYGDnzFkSdqKfPup8qlrkNu7u
P48WKyXFt/GyHwRttc/1AnQrKSR5NDpccEaDJysgBsFfxU3q6+k9VqS3a1o3
DSkLqhnUzYdkc15ABs6Fjb43zjIbdmyMtkXCqnVyGWNjGQMafKbXudpRyTD4
PaGt+8DqjKXfQnEMf2lCQJSEENpHmMQF0kelmHlWfiejteWjC1Xkc2803rDs
aUV2F0k3quQO78Z/uyqBh0pzUJGk6Sjvz7h/TexEtxHf/C5YhNt22deElPJX
dgKEpXEBJW7OL0D2xrB899Gf1El1ZGI1p+PcPYCZLHKc5+lwayNbSrHqG8TC
gmHEsnVcjN1i8niN/I7DucksmnBKxsCLmtmDfn94hcAfZ5sMOpbVXKgAjB56
VUSbjEQ2mAKYttWU6Jq6k7YdEbP9kkiA5ojifFRsnCS1kxZQhQ334tuLl+pp
WgF08uTw9eQYMuoOspA35K85340FhynH2l0i1hc08M9g2MP/sJTcbohvcQ4B
kMcFd091izJV+1cA19qbJ3ew3tGd/6bSF8sOVulV2QZgDtyXNTnvEiFnIou7
vt5OpGC3h6yh4a89Dbl2Lmt/3KJcxYumUdQQYnbmqnqAC00jg5xxF0SyF5nO
P0Sou3rVnOAoPh6Y8jUW3L5IA/3EKxmXIKFiWeU7oXLbLkI06w0fTtDI2COP
vZn48y/ZRUu0jxI/wyuCvcqpcY0pELRoT97EG+3UWaJ+6I6Wsia/OXENEk9p
WJxQ+Iu/5mbO3BppAHDtp4ZHtOBFAPpVPKkL6sya7yhL8907gQ8UuR0ML76T
ffFXTEaKG35CkaSiX4b+mq8a9QQHdtaneX81PsvZ51rIN/dHV0OgsmKGE1cL
rtu3ecvnNoD5zvy/hxAs8qGMS04fRp2mVKXhI4u5UV6uwUYvutLZMrFXdIbZ
Vbs7er6Mw8GPc4f1x/uMoRVH2UJ3iXUFNIZeLvy89jrfIYUJtgT/0vB72T5E
a0vQKhGU1sz/uzVdJk2SIp4QmoVBWUg2WbmYA4LhknoUwm4LqTxmso39qqFn
BpBfrBNUO2LjRXhcDqfKobeQAoCtMyfbrjIdXDnjViKZJz2GA4YPWYBuwwFX
4ultTK82Yq5OvFc9LmLms7ynkHHBuaT8rzVFQXuNkPjGK4scAGNClVHRN0h+
n9MPUPyfSeeeSMv5mzVVA7ZyOActlLVVwoFWFSax7SMVC08eTBhTgnsUEV8J
ZrbslpEUKZocvcD6iEfTGLGL7kw1nIEn+O2yOMTRyZkYaLPaPaFEjrwy5Z5s
EjBnO9znB/Q1sGZhJWdRWq3u1yYqqcaQRweoddrK3kp+pL/n6ooNI5r9LUT+
vRnmvbvW8eG1yGRkGVw0jbq487Ipf87eI4CIgrURbut9vo7/+yFUZr96FWpE
04KLTVSuOgn/qXGxpAu/mSpve/TOznB8zHeNagpx3gKaDivfCxwzuDQbsfCP
NGY6To4QNgSSlGcczX9hP6TYca78FRMiek6V20a5aGdOKwZbfYUw204oqADg
fak3aCUUOh6BlmDkhqEYENy7BWCbj39eokgvccKgkmLuJFhN3qsTqqTZ8YJ7
A9ivwtNV7PYIyTxkD+/uJJkOzphbvUXpjpCzLe6GRliN2obuP2mFwEqwr0N6
K+RR1aXnt56ZGzM9mUuoGhopH3pnz1Z4GoZ/kTXsd12bbQnEBEZMLNiVMh6n
Wjmnqbe7IYOobtWbczHV9Nk88cExodCs4uWo91X4bT3GhplX2+DzUZvFFkAh
Khvjaip1HWcLzMbuQyvjTATdJbvIHnjnF4x6YPgfXAxRjYVelfKeoQ0U8KYC
MoAaOYdEi5mEV1OanBgWCIjNYqM+u74lnowKfiRbZL9DjFic4Nkl4x3sQfPu
Of0O8YNNF4N/fQwhkaLK0UznZr3sSxdMqSDMXZREkVlOuK6dh6d+/wTUia3I
j5o6ZrG1kKZSXwyUer0ojyn4xtIa/IwpGafIOIhGRhUnoxSQMoTxOThtua+9
gEKp1TbiUPM1GOhBPTLbp01wuUpVjKHmk9ADGZhPe0Oj6pPPOhV35sMGVHiu
MrFpMhAiifFMbJa2MriyBF7n45aWSKSq3d2HAikrIcw0sGkJD3tppBM2z55a
pavko+YJ9n5COszO58fYHm8ScAjqUYX9r4iFVaN+n7BQNZ/vuUnQU5JGWTpH
sQORwsn58bmzues7d9P5XZ5OvvkkyypjuhgxSqeThT0RDZ/t5g1cu+klHMtb
IzdVTssdgGUDEvszdtb9k44DWpGCNeO8etsHu70DZhnO9gh2wOiXy/Cl4EgE
mIuewEOle1wCJeqHCqxDo16qayEaUH0p8BbDnljkVc05CGZXF9MveVUrygBd
7vueVO3CVys9x3dB7fT1SBdqfWcUX/r4N9y+pxe8B/iAG0SNAkGDblaA8J4u
ybMcoV1zE5Rd3CkhfauekYR1TrzGqddCMsYy+mq3p/9bQtmp0F4CwYfLFHfP
a4Khk3P4CfeIhQI7ZGYj+E7+vLq8zK0GwB8odj0etoc+Q8CBJRIua4zI11h5
P9Fi40BEUFqIfqScd6Lh8cEnoHJrByf9yWRumW6BRRBHeOs7Tc655NAPEePW
EQj/M1O5CkdGHVbGAfZHNkS6ygXiGD1rbZ1vku4r5UZMIcxb8R8WFol+a82+
4T4zBa23fcPLTdoZ+n244xEP6zq3Rwh6qGmgJvhGiIjDXF/UDTQ2bs33WgWd
r0L4ug9Lroz3AmHhlsxiiS4r4TOXLrRnx6IYr3rpJdwgQExyn5k2PtNYAfNq
Uwuw0jdsDF1vpMn4FQYqouxfKwdN9hsMmpnl8h0j002aYWTKfFXpeDIdSD46
9L5VmpROFAgKpMTePHrQEMc9wnAv8EltxAdqcfDX8rc1dnMzjlMFJmBuJ/zA
tDTPX6NUNzROviFkgPzOHEl/rFSFC6JQKwyTvEMyIeYoTu/5Y0ZWzGxdUWtf
FedlrlS+lU1qEXxV4D9T7ZYp8tlh7bCfH+kAvszmXYx650P1wKCt5rUnTx43
xvQJ4O/E9uk74xd8Dc5sBtCCzacLStx0VLXHKXpY0PIyyRj9cO12FwUoHg58
6wH3wCmMpuxwPC6tdP17vT9DW+78AfiOyw9HXEWGpylEMEBvXv7LZY8A5t/Y
3fmAcZF+8GZ21jE3MVU4zlKbuO4kw2LrPEQFkCnnqpBZ0w4gYdH5++jy2/5o
zH5YoPl8eOmRJomPPfJzCMpjvpVxa17HwnfMOybAsWZWepWXo9mLV8UXpX25
3vDZAw9K+UAL3JPzJCC17kvlbWxZVIEDRuQf2ZThjArcQ53eNhmQIDOfOrve
ojUDxW+lAF6Oh5+uP8Qa+5IdxswfLt+LrLg8Jb3+/a4+rQoTY78h1Z21Gkmo
2pK1HWQTJzShTUuHhfzUBJ8O1cqdxS7ab4SOGUy7k706yfIDZuTnh2WdEgHy
Cqul0bHuTE05uDUnbCkxyowqPODc8xaYo7lojnSHPvo6yiAnDQ+Ykmlrs12s
30DGC7T3W2F0Kh1+YEolYzzCxds9lqukrWDWwzmo48VMLEc1TIz0qEGtQlqr
ZSYzNPWNCXOpcVmsSQByCyOzBdL8ilyAijYgu2KIpEhOn98LxvnYRN8Q4YBF
i8IUQIgBa4Fv9QgbB1KLvMu0521nnM4ZeAORFgwLD8d9DJbi3Dfp5EfZEkvo
R7dFIqAXVmU1y1nYUfyjN97e+55oza/Neg+KwKxbEjLbuF0dQCXIOTz5gHlx
NIyNrdjoObrTYDGjRM9bwbhhVpo5S3cn1ZiFIHQ68Ny+kMGzgQI3dSiZ0HDg
q1eQyk/g15CxaVha1bMXsWNSBKVirxxCsetcgsEuGHF0cwWG6HkupwOGpq9M
O22omY3qS4LAZ4xtMCMw/7y5Q4NMCyz53oFfnnDnbEoYIp3M0iozAER0k5Mb
PF72HnxxugsE+FO5KS92V0Ncjx4IFcoWpaVZgBzkCZMVNB1SIU69H184JgJd
88QDjVdiaZ58DD1rKMIWrE21LWtc4EkfJ9u7Xb/laGgz4sb5XfGFClk1ZTxJ
66U1S/bcyac9IEs8K3zkIiS//nrHsmn+LC8V+lq+cCmuO3ypuuKvBNwhd2Lk
zsk9sDDZ59XpuXDeWBXIeoNX9K3mJTQoOWIGbK5I5PF0kP9bUypOPkuN8MxA
lx8MErQBXpyUP8OFsPHaQRxSj/m7Eel83xAW/xcyTp173HQokxT3HwOOvkOr
hKlUkXBau+DOP6p4NUkEyYfZlWXzx6Le3FShoBaEWU+gbPK0QMAhw2qiLYC2
8qRYS066zXeGM4lJcBodF0IMRbjosZGq4wmTNtxb5FRYYJxXLlueXl2d4Sp8
zTEkEc7NSOxAXZJIlsZcAWTGOP1YxkasQiVBhpsS1Si0luIzjQLQm2Et/lqN
53S2RnOJ0Ke/7kiMONgd1KqPynDOzfxiYh55BkrBTkfsgEQsLgHklZxHrMTV
MMO59e1Kyaaajdb3RDguNQLx5oSNmm49dHCU+KSOwEBIRxGa+FW0GChJiNzq
fvfGazEtEt3SqM2cbRS2f3lQ6pkn3U1dieNwLgKbcZqSMqm38IEu4dtHENgL
WQKBYMWcf1v/um0iBsG0r+nS/vo/wlysvyoVCTfK/ct0VMHV3tuWI7Y2LNrJ
L8x3gEgGuvRn5UNavGdO4+0kvCLuVnGdrUAfetLzLRyZV0DA+pOSV4x/9z+Y
8XE25eVTOpigZe2g7YeTXpPbJ1s9lK1RaglLNN4ECC+EVPD3DEdQn/K/4lpA
bYW53vlwIh7E+YfjBOh9AdBDl2AwSV0YX9rudrbHlqvCYET+Bntx9Z7eF6bf
rVWoaYEtLcRQRMDSjQsKU99khdOnuRVpn7rUEUHklcPBzX2v2Mjjmi//uiEY
8jotNOJEdCCGXEmu5o0PVw8nzlUgFBYsLS+k5WksumUGx1w3d6dHZMW82L6L
RH4VCt2Yu8ihgvCHCUNbRcHJogftUINVsYPGnAXMtnKA6dPACo8he/v273GP
vF7o9zs9I9Gu7uIYns5HSJejFcPBXlbVxpIf7qOxbAWaBUf3n8VzGu2abyjB
OPYj7jqJOFdip9euePhTuKweii0qaDDrfafLe4hJLnHeUB/ydRh8Ss5+HWZu
qvgBw0DNsl6atX0v/GRI+eF0qmPGnq118Mt+CHaFJhrNo2UIwr/1XDl85F/j
YSl3oobqhtvQ/uVCPA0i/j3WKrNJ3C2GghvplLSRY7X9stJJcwOy+ACckz+V
JM/ePFvcWK4x8+UXEC18g83zJS9p/svF9mY7HmiUnOp2t4v/sgZFJbLIgMrr
P2TGFYQaNFjjJMWcJ7s6hx2VUx7NEvZGXosRuqs1EdjGHbMtR415nXJwbm2K
uNNQJAvhNcsMm+qxtUTY07kUG80daa6d35qzmFIK3UaZ3xTS0kFu87nEkT2m
HSpeHuEsWe5ObZEek3ISmMvVOZZcd4D0HlYEgNy6RZV0J9DDrVPoHrgKJB9t
oWkmEn1iVtkwY6LDKsEQw+LBUJvSNvKMOsc65xfe32/9vyZyMgZUeFiJQSbt
XusBcHR+gWmLRl3zXwfnIZyPGPuL374QfdBEvPt2zd5Baf0nvrvjrHRJEqF+
rXiseXDwddju6D6SuOaaKtPA/z7QXRoFVirCEYPA484PAjY2bpDuEchDWRWW
UfvuYKJ9/ODc8SLfo1DsxcDYi7HnEa//29Av8RX/nKzX7Y7P7tN71NGDlMMG
T3qRWjjOLN2hQntIl3NwWOAQFgBOf4UxtPH6lMQ0zLQuh2iQTrQ3UcrzyO2o
RU5r/taWvXeKkHTJNNt0KvLwouGG+bFIFJSN3Vqn9Lt5SuUiWR173anZrKu9
kE7RoaE4eQ5io3KeBNqPGbK43EuZV2VZjSFRhk3QrjOmuQkwQb23zUCwG0K9
NWIY4OjEFiRY0bfxeFKYz1zrCabwVW8CLSwbRfpu/i8K1tDnKXa3LYjgjine
nfOknappVoGoeZwf7vf/cBljbqX+UH3LdVM2Ss+szTXsjxMqKj/+lEsx/5Wv
7eLGajRVGBVV6Rug0tLCHfwD7tsJoJa6Tn8P86rgN212eQM7VTX5J3cw6ZRc
C9L91QR6kwr4vG7EYk5rw4rzQr0iwoEcG7vej3HeE96Lc1hIVu3zg+jJ9B2d
z36SDsnrzj1vVrNnMVPLBjAPcVU2rd77P+CHeS7HqAaOaIe1LQ4j/ezS8t+t
Fj8Fu94tcZpX6sztbZG1DOuCUiJd7R/wWLBdTSMm1DJQrWWWMonTRNnnTJMV
x9aav7q2BJ+C5r30L7WthYesU6pNoanwTUQU/wnkmxOmP0dE0Z12H5iACTAX
zURGdX1JAAlTNp5yNKyPuYXWPCfNjleKjJe3bmdzu2Ymg9G/SokM/kWacRTd
+SRLZuTToTNpoCOWf0jU62NPqXz99Om9qST9HN6zOT+334k8fgP6/I1oyyzH
azjjo3md3zMHjqCrmtCBdgaGf/gyHxjIK7MLZ1k1BzNx6H3w8xmN1Hx4onrn
PnYB2V4D4kA/u+7JjYF/MwuKitBJIeznJYiKxxtXNACKr1pEDe4SCJRUnhEF
OfYk+fbbYOAU+2Q7wREFOuM7vPYAP0mD6U4DBDSnxdFszIraGDs869LQOX1d
+DHa9XiU+PKHSetR2XcOGj87RL40POkdBfYHvx05tjICK7vPYmNm77ogZpZQ
Jlo4Paq+IYi1YR3E5GjtdMNEAOsbO5YOZWJQpPx48dep+zQon8nTEZZkc6K2
q1qC8CZp1h1vMJ/kUB94d+2SQ2Bbjlkv59bFu25aKJlHq4LNfNfLYKxh/9t7
R0duXO4jj6B6r7FdP3uJd/X57MPAQ46jluGdNqmng5Lu2iyLIWOTX1ozqHfV
psMSiY9VGkaN4SOfZscnFo1XYAl/M25Bs2EnNBMfwqK57swtydjaoXgiOgjk
7B9IzHTPOlPYJM4owdtcaP8IBnUECrX1PAwi44hNkDtgOMTEeZZho/tZQy5a
ZNneTSnxlp8KMrWeSJwNiHPTSE47cCPO+clxPlmDlb9iRkyeaDJHNTxu3TQe
qW0Qf4hu3vYYDGMEa5iPSvPx6k1u9nUyYs8+H07mZ93eTKOp+t8l560iyufM
sZp+p1Y9tK8L6p/RFEObnBrhAc6q/UXJLTU/Mh4wqUTvQw5mB9YSTDX7kJNQ
Hf48dlfwiK6d8uradsNqmDJ8xdpuIzPzWFXQae6RSqkQraFng9dOS5i3uy0E
uwG3Xq4tS9Q2sRIIOKhzbpsb9jxkPoH0n2z+qZPxstDhxZ+vu4zn4/0/Ow3W
Gggv6VojPft1jnVBklYaJthreRVesdeY6BMs340khjE18pJ3R65TDQDQEATd
h81NSZPjB8Pxy/iyb1r5MdusZF6BfnH4PhcFT+RmC0rNkp36M44peB/uKr7y
p5j50a8hd+dezRdeDHR/a6mbfcBuVVP3kWPawSGC9nrpJPhY0eE2MLuyoiwG
JV2QJZTbA5KvhSEeuefWYL/Lz33KVHUOoUX7g9AzKzrsod3T8k64kmSJXIQh
eU7FrFmIG8rN1frsnZh8d4p+0Ig5WIkG4ZZNgUFF8LTXNFgyKZsBIVDTxjEg
udj+Wn59xWO+/05j8F5LsY91D1c/c09cxBSQM/2/Qso4TmymOEnPx5U5edxf
Y883/YvzXWEoPs1zkZGXPmAl0KA74Lj9+V2GXKGL0SZuIa9CLokP22p4AVUA
8Rk6kVsWwVWXF5e8sByHGuOclSuP6P5Hbl5UpmF+iCPx+HGp9/6LxVKimAhv
G5xv6lGDfWpBKMY7qnE67MpqS8hOR6/3ZPzT2doHtSY8LWFHGcqvB5k6woFy
oQ434mTK/zA4BuIYhS4PkE8fwubLQptbID2VXYlbWQgZ8aS1lQta4gJgmcZc
HhE7yX6cMwMMK0Ct7USsA/IXAo5k69uJiQG5ZTd1ZK0rM94DrbfiV5tfMN7u
B/7Jsc6VJfRyZkKAfHGrQIr6b7bijIZ2ZgNCBGHqBKBasw+MHI9LRjdges/a
AgcL8E9csscgIJ5xXaJkM5Tn8NoMbaWLsyUO19i6pKGUSVlc7CTx1DOS8ltP
chaODhZu6ydt8p75HDLSj5zYN9Y8n2xOluglHZwbSv0H/a0wcuhvSyqKVRe5
FB9tsvpHNuHwTktdHChgznP726ZIWROMzFfWlbgzzayth4vCAHJ2VMHOP2ni
/eJQ2sUhc8J9GuGxoLVS6Nbp7ia1jdJswFMdfCTjvSIZz66XW3bfMvWatUUr
LvrHmobpqeTzwk6yDio8ECDBkCInOO1o1Ays2Ukb5IQ4kKg6HNMrN2JR/NLJ
lyPj/Nzk79ti9XHt9vbU/gj6D101cLm2rFI/hIZpnIbB421dqnh7jjeT7N7h
IjoxdnJtHPMi4ZfKbNcsiyuF6KEJCIW5lhBkrGqPh+x34yWs6AUy/CiZ1oMj
eEUu8OSHOSuub7+dNhcOttZC4L6SQDQqJ70aopX2B82q27U/qDBOuFrLD0kK
BKknO40sMP0JFtXKF1uYKP7wGOviv4+HxL4+o2hqBsnqodES7ara7BLCbXsh
RQMfeUgcvjRPiN20d15VGB2dsHntGcISR9dR4cxIQdKE2ZvKXr/UgW+l8zQT
TbIM47PVLS3jVOJUPULgSjqzuSMk+AXpk7ftpuO07vitZP2QgnLTbr2WOwFd
kTO0qQll86Uo/KWQWialF16uB3RAfb6Gm6aHRkL6QcDtEwYND93uqtV1XsOX
ucMwuv+tdp85RCBENHrdxB1RvUZUl82C90wI2ISByJ+MkWByUXFG9txdIYu5
9CrJmaWIVXLtR6LorFFwD/HlHOqXUvXjmCg58WjP+2dCFIzDYVj1m8b1F0vX
GG+535PLTjc94/gAfcJh7ppkTb9SVEnIQpgPDJDc2KE7gA5LcVa2V398Zr/H
dVYj7+8MR933j+9mGOPZDIjGeDm31QiKJY2EhVOw1sYHpveoOatnhf38veHX
cio0OWUfQp8dXZxd7wpt2sIXpz7k7XIkavY2oL/pG3IJEVhGABRBX1Kl4p9I
GoOdbu8atFlu4DosKQRytxLjqu86ESCMFfyqEEEF2iEJlUA2zop/vxJAV0cX
VwWf9DxENzoUcucBb5Yp9scby0GAF+M+FzkLJTqwmXdkdECpdisFa35bUARr
HcAnmLSN6fcJlf19oYtPumcIm/w8td+9PAOW9atP/et55ZUByi+BZ/00RbVs
Mq5xIfi/yNkPwc4nGVPiHdpImx5En6ILuENDN48KXCtlrdYLqX8Nv+Sh9t3X
8tFjzISqkV2DZ7rnZjR1NSDUSmbeRW5K2OyI0Q9h5naPBIL35jl+Yno7aSNf
BNB2Wpln0JZVrSt1guVY+e9+LbYVBH586q8tiCCr+i8GMojVmIU8e6RwOv2i
P4aJ+iUyVpnTF/LrpnmJ4k0Hx8bQnI835hgYStkl3Q/x/l4OJK8/gn2GHiXa
T/5RYtdtZKQIrZ8zbYlR++8+LpLqtqKauaX0Dgtgl5Hkc/JMYW1EMjx6oG4h
60RwxxGZ7wGEzykdrqql67HiVMhJnTI0YLLf3iSyuLGKVHbXluEwXhTLqT6j
p4QWmHpCuYMnkWM2rvZL/paCGO/wazMgcnWU9ONpdd4hbVf7k7s8u7qK+9Zg
w2BHchx7GAUhkOOU9jtbziny3Xi+surO87CkTeZYSgGUef8D7ReRxdGtFWUK
17jO+anRofTwKAtpurwbWxpTr4sTVtk9TFC1iODi0abaMs/kJwvBqh03+DUn
+aOHsEMC+bYL8d8RE/qr3FfnfD77vLguQFbfJ0t4kmNjOdN1Rrzy1RsaDk08
IRbJbjKI7xsJOBuvIqntxG1N+BXopBmh8POjaNbYI8Z5BLz/jpfv17kpiPuo
q0+tS6lJZ0gdK5NrJZXpTuiR2S2KpDcj8/0XByxdNmeRsA0CQkbNdmijWLyS
PUMqyNXD5DmNl6Dhnto+/Qgt0seb4CC4o3FSr+TsUioavfIKtx0g3pttYfpl
MvPZjCMUdbSt51KORyAKIDe5YX4Khb/nQBILMRJPAW5zADDDp3fLTM4sU9Sk
tLgCK73afGMD0W73tRWLPzS6APNBAxjkTjxiBc3gWABUPhrxrtgyqiOxd8Q7
KuvdfV6Vi0FZg+1MSdsm4gzMGoQ5sgQnAaGi+5ZqOn1r37fGImGUhR6MMyS+
pBMCrh07vZXsgbUHtRNXcvDX2fmUoA9qX6ymrdRlr/2gTJ5CzTitQpGEW9av
3fTG8klVN7BKdrYTbZEBV9Qqf7v40b7kUzaWJV2GG7j7w6buWo07fOyO738Y
25ndfAu7eGhebWqbyWKRmSL6uWpC7Ih2d7ldSChljjPBo74QEJBAB85uOTqU
s+eDjf9k0nD6tOOr0oma0h1B8TcLqCcGF1ChmAIYiuYFgW649F1LHBo1BFzb
ktydsWp7crQOkqTfACGzgvFFGJPk+xome4dDxBOKpkuRjGkosN5U/A6rjEgf
EPUJDjq4+p0BpRocpw1jl5MkHZgqAt+y8Y0mj4LFiCIN6x60Lfn1C5Eq1NFC
VCYCi15ylIVTLSHv6FuTk9Q/8iAS+cIWb1GCJPmi6hB0pBgHFt5NdPrN/zfO
urzrGA8JZFWko+6EUOcc8DMd1ZmrW3b1Nvlr4Kx8Y9bcB//BGjxQyBrDghPQ
gTtZcqfIbLu0ERvOzjsKaMhnOMJDdXU1/ie5IivBvmYzhceRFlRNA23gbdwx
4WoLVqX+ECDlER2mcdbBHjC7wMtz0BFD/cZYhNiZLirOoQeqVJvuVh4xhRmK
mQpQIoUS7ahUhskDF6HonW5CFeCftnql59QFTcsJd2ARegyq2MLFUgXaxn0d
onLFIBIy/o3Ly9QJtEH2sWY13UD8sklB7JFAKghYVl4cjhn6xvF9mmt7dw7U
IOCU8Q12Zhu9wpW0GKEaSSyNJMWgp+vu2kY9AM2Oto8eElqutViJmE3y1dQh
PGnfVc4pSpicjI0hPtOImY6KFxWzUiORHxpcei5smJdvzEhfLOyXbguHFuGn
peyCBad///gCmTipp/pw46+ETOUIAxOe7kbZBEKvFlFtxYmSF6hhMd8ZjKUk
mesCgERVru0k3hRocmY57UtExjQIPvPgd8Jy8cqJJ3A4xtQVmzJEGoGPP3uz
eYfXMPt4C00Osr8R3UDDzzhvOvvrboEKJzyGXT+UpOVzsSOQoL4kvOV72SaU
0lPB3seu+4b7dc1kjnRaTM6yVa5qlGho8qsEpqyNR4OH2FOOzaBoMWGl4SJV
IL0/4bU+M9Xyy8ajsX04fX3jJBwnO/QS1LGGEfPPmU5/bFJeR5ZK7GhYqaGH
U1kpELOfcdB4ByN/OcYaAuRxLxiHQVf4XiPKD7p8DXp7ZTdwD0g+BvFEoml6
UVtXByRh9GYl3zLjMjQ5ZweeEtmrTiJFIFyMGd58Qgj6Ze4llRaawFANOICI
rpWBReFyAbWZkcTFQLxnc4+Ds3R9bBU/fJCQjpr5vSbIvtVLuh2fFAf4a1FU
MXqmdt6Re1evfLFSHOSsEdJK/w/Q//Y4tGqSnbuWPUBcnfUby6t6HZ8YV6qL
ziMKdRL+31cDwOuYUWzRpQEjNuIR9KfOM+sjLMN3HAAfnKuHCSXLu0tFQV8c
uuHabx0zg5bOoWEIVSvfgicAa1lTi1ZYI/UCjTSVKnzfZm7YixTB64i1E2Q5
JbkUyysJzZIe2IVNpL7hbTl69tfxBWJ25JDZNPsYtUc/Mo188Wiz8daJJWwj
s2+aQvWFCH9PhJEMwO1GEvrKH3Uln8ZQawdrtTumKBPA5rVaCKWmtqwHFbME
gVlspmk6bdB+eIIVxLJF7XErIkm8TWFuyVTP1uRiOB80S8L2rLlfw7lMeTA/
Br+Corb4WPsSIcPqGVXzOOvozhVB48P07B1ZR0L8+D+u95FsVEm4cH6o4DKu
TQ9vDO3iiO/jUcmd8X9NjVs3t4nbPrrCmxSXZpzywq2Y9C8bHzd/7Julfvbk
uwg3vGgVVogkXLgGwPDcMr9AKEOS7qHvdGOvoa8VzEd5Klo7L7XZ3wUDOB1K
9ReYlLm8oyVG36DNPQpm9EvZ7sg8faUDu4xjE4fRVXO7YM0LXsSjCcV5ZduH
oRMrFO6xYzgrhT1qtZMlLd3hEEPGlbeQbPOQojxisk6311J0pNpd+kHCp//1
DPNZ5dg28Ue7az+IdAw7CL847ibEacCSr6UAHUtTy4nq23Wc/4RsyielHX7W
4BRTkHZr30bTYbXrNba75gQkGIsqKmrTUIA0UGlGyK5FpgkjdXANHKPW5nQp
P0Y/1VuOgjIpoboGEL4yTBdbuAxrHPteGbYSUXtOsZtGAtXfBuU/jsQEW/8g
uKazPEoArBHyqG4IOoLgh9kVNm2MrMtWZya5NgZ1d50TdAkxDFYRggIx+kTJ
8qzLSpOrBJR9NGp7IdU93YPti6BR4fGLKDLXqEgwjoEFY7etvPo3tl2fNVbs
31vEsDJzzQsQRR9Y17mBvqjCPZcAYKg8ln9bODZU3qnm/zOovpoleKwYcNLY
1mwq7VjvLjMrqxfDUMozYsAd1rNE3JEYQHSll5Tt8jhi1xSQ/WaDo0CSxLzZ
yZg7D3TdoaS9fCjJnBQcVW6t4vPp2EPCf82w81fyFUHlQkxqTldgqkQeUtNh
5+fPjGYx1N2aaHAvNxe0zZI1zXIsoOuegTX2NBheEC7tRH14I/zQfuN/L5RC
c8RVCtk6EayQbQWL5B7JpMsnjE2vScJ4Kbgm3z5nKrjdUaoYH++M6A2kITa0
QjLeSHor7DZn4oEMvGLQ1FlhgnScC3wa1qv4/o9Lsg5HqCRr2lfvUHr3BD93
WA3cBsNtx0s4m5HjROcZElwT8y9HnLzAuLEI5XECfQ2PHgOi2rvApManXZV7
FjCLkOFNjT4tGN8upVxClVOdKStFmHoOgLKXN7S+VRaz50zdxR6eYu8KrxN2
zsiJXA2XWa8qaMRkWlmZcqcyx7YYglzHskHX1j8hn8DBHcZEvolSm8+uo0nT
3L7e3ghxeSPK/GHBh9ngE5ZWEfXMxMmfkGe8G1cSKH3M9E0XA2dcW3mR9FbA
3d4YONtfHR7lgbr2UfYcAZ/blCDZOiJ7WmtoOFP0NQsUvpBfcnEYWD9xSkN8
uYo3D4RjuBKwvVWe5SKnM8ZFKNBb/emXt4QEnID/p3rJKNWtf1AFlgtKj76E
IZYqlBgfH//yFjBsjZYNBl2m7VFDRPxv0oPK6S+V+h46/5ZsgVnzJ3QXwnEh
Grl3NnTVfQ3I0A4B5gLW6esQJNnz3jEuwtOeB0bNtXPrcd35uJDI3oiwuZje
xRs1ENdrbQGYE6DtO36t3g7bmf2mqYbPmXjUoI75oM9SuP9KMc8kRawFCg/Q
CHaDACjN+XAHfesXeUKQk/uzMKnkIZOoubGw6gROn8vPjRYurFFVtRPA1V8H
3Mo4AhnQ9UASWMgVEplzp75aF8Ag4vamrpJUJoCk4+WpgR6i9+yehLxsAzFC
o3L1mIcwMInA5HfqlfaLawoNYfRU3magz81RMy830Dk8wp5uQsWZGX7wBUet
8jNUC1Hlj8R3sRGlns2Tzy7IAFJlUWshNyQIiiIUpyKUkmr+Wd7aJQOkU4OV
54vRTJEI0xEXqAMGLrvL0AeDI/qHk+y9TG9Unuzi2uoYQUd0g9qYmXDSsAvG
wqFNjTmFQmLztkK53B0bYHA4qsHmzdM8FN+xtYy3lGTZu64jcVsqzIn64g8z
zY5wKrXx8tQuQSi0XT2j0F/H/egqiIs8qVyk1XlQuXp46+tPyR6nZ8/ik/cO
heLxMn7XQzsRz+Qa0Q3Euqjx0qu4KWbL3/ITqX5yfmici5bzVYAeRpjM+QZf
l9Q2IJS152Dfqx6bLQnZFTZQTUf4JxT9c6lYMjnQ8JpKWdCR/mf0OOwm/ho9
CfMHjgmLlOobIVWRTMi4MY8zqB2AZYMmwHKwCVHc+k1rg5gSMBpKQ1AtaA2p
IDTKFHQ+DSgbTWA/MaDcTpduZHnmeLVGkkWZj/wzXK2NIzYveKD5I3Gn06Pu
j1mGLN+H8/dbDD99Kou5Q71UpjUMI/GSapw7bJZGGAdEdVaCmdC319zLtxd1
JexYi2djnqFEC2ucXV+YaLCHo1q5HH6R47wyg1kH/pgZBN3rT3cxqigeR4yF
Q19278MRcJIAajUJSN5iljfHN8QpMuITLGI1QYU/+jWTw6qgs91gYEjg6aFn
TUvnX/Jm+RCxQO9+H04Cc6rU5wK0WG5vSD2RDWU/6cs/exx+kr/KU4N3TdYa
f2dOzr4dSA1xTtF7NvHe9JT2BvYUmSEoMBt9Qj0KM7Mgr5Q3kPBK9EQxc48D
CVH62F2zA9oGC9Yyi6CcJWS2cZ7YbMc4kFS9sdh/fGN6tJR/fIBbsvAEHOAW
ScX4F9g81hHAW7XRHHclQgk78l77F0kBWC7ZF6IXCMjzFGi9tXJcHsfEeq0/
xH0CmyMCUy9ZYNs9On69T+M5rZ3GIB+V8MVFXtyps9MNf+TKeHvdWkUBC2wW
JPV9Fq4fL/atmLL81SxEG3KkXNiUGl0wnqjmcWVcyOoGbpDAsVPziQORHKON
quwavWRyiJWZ3/Txu1mDT9sKHkZzCsEEFtLCtis2TuKh44ytr1LH97H6c3D2
qpmNVrOm8vHVQy6pRcwJvHwgJmSS6i0jN7yvkx5cvZEAyz/Gbee1dBrs7v4v
SEtzQBxAp/p9DRR5qtWvfw3JAKmPEt28TU5rsjITVAGIkbefs4jvLLYP10jc
7CCvIOjqTSCKFblaAwt7Z9POUhDRV39pehBpsEBdpymo20a4iN2oymGbhemH
i1Xv8qbKBeJbKmIdHz2QYtRJIqI49u34pUxKsy1wwm6ttw43RsXu6Lu6VeFv
GnN0i9nRGzJzB5CIGux7g8eMOgYUZcZq6F45dKFs4lxzKsKeBC5rdQLYipgJ
jz/qKZDa+uX4C5UJqeeQPIBsSvjLSH6XUag0YGptid3z6WNXpKbqzLcBgOXf
w8bFk1gskXmQznv1UworvmF3RiLK8s2kzwZeN1LklaWbyX74whbCkyS1Aeih
dzZgFlyvks4drSIuDiDldT18WdAvI2EbutlxUc70o/GMSLnP5Q3Y8j6OrACa
ZzbkuSPGjOFjHNZsU6nG6FD/aojmyRQqfK54UHmCXQzg3gHPtBZ3qUQ6q3eM
NcAlciNE2mJ/RreOCw5ihSEYf7wSFov6ChjtmBLhfN9v2tqquOLlJLyGphdG
6V+i12mkJqnvJq7U3K1su1Xvab9c9oppk80i7gAsaKdh86ieCEajThe0WSo1
niJTo9kj3K4HHBZI39HH/d887DflLR/8PTUK3S8E1ZDo5SrVWzFT7m3vAd2Y
rsz4Xd9Nm9CpreHnpv8u6LIT3qs/kQqTIhxZp0nGRpxKfH20n4DtHp58TB1X
RnzaNK4kyjD4sbJ4CFMp8OVEzWyn5q4jxlxpA2u5Z8F2M8qAG4pwCTGgT+b5
IdSSDdcNIthAuB2Bn9BtAyXGAphFyWJ8+qDkj6ESMIwS0HBZcZzK/4AMEP+4
14HZW9UMRQBMBovJhestVeBqEWCLMca5/DaokGW5X1QFB24+ur4l9M5NEyg3
cImLVJ/BQhz7iVb9JJ4hHtZgj3jTeNHazf0SckxChQuarK7pCFC8OtJ67Atm
apIV+p7xTo+fq4eIbroi4adtlJP6eyZMVo7phIFscW5KR/v+68Tfel2uowia
MVidZheinb+kxwYB1i5CNeLLtvpUFh1b/tnSH2js9tyPt6XVNoeGOzVH8rxB
STZQl/CbtAUIhtZ3tndhGJJI+xBYljGJnrKyMWCuDSXOu2DQ4+JmZ+2aJLz3
B0CCQR+1dfIw/delU0zqksIXdfjA5CtiGKdSv8z+2Qfn5+wjc+nBohqEIzL2
pmY+rG6+PQ+IciRLGo5N1rqWd+kiaFC3oQRhaTOdiQZPXhzGDxQMgKKqHpHL
Fq7WNFb3BRJo2PqUgpA3anqWkHt0P2GVsNfao8g1taM6dOjhwzAW+haXiyPD
nSCcp5naozfoks+gth8k9M3kMTf9SZttfyeMWB8OOzaiHcTjEbZMtvbBBmGY
x2s31ZhcPJd+CIEP+sCPhWkFb/WU86onFPo3CDT00o2g28sBinLd+gWp0IUv
D7M6xJO/vZzJg9KE4UgLhIB4NGDm75LBcQQNdQjsDUICla41URs6jRQhfTt6
HBUPhcJ8L7YIwbfMC49Evw5cFJ2wH6hcppnMYrzqCUSBmLHeMHBt1OqNPTal
8PNtSiHvZVn5gIMLr/MZVGoZftQtXGmGoBrV74A16bjX3L/senIhtzMHNxzw
eOrUSJ2L6+keW5Qzet3X3dhkeawZCgPio9Eg1RXbsKQ9/o7RUNVTmbYiRe5n
MfzEubLgNIylz4Tzddmufu3FoUIYqclLPHoMvMWE3zXJxrrDqy08avrv87Um
ixi7wrCgU+ijw7CPSjc8R8YJsaY48RFa22956bHyXk3M888hUKxlxPjdEXQC
v3jUQd+zptQzakaBaERuD8ufWzfD51igqstyXkoacXOTHe/07n/HWlTgyGIE
uiND0ZXeNiKkFewb0TbLqvcs89enzsbKvpryRcLDAS5YrpJ2BoMZBbwAKB66
2H5tuibPZSJfCrjrhFp3hAs4vv52TVDh+zM+nMpEEYEBJeWvgHazMuw5tAcZ
Jvy09b9cXLnBcgdxa1s9YiLvAaHz5uokGJA2kYtInhmjs6nrULMGJaLkOThD
TOZeqoPLZJBfFgU+bJWdJ7BUa1WgMSmT02E5c6ft0dZOgaSi7Vr7+6sI0UoR
nNK/ogLEMDvzW1YRAkgMtpuLRpeQAv+O8g5wW4eWrM6Sc9buRXlDt5VUtgwe
SaLS0Ju1Hn9Q102RmpobOGO0RPeXlHTzO1CE+Eb7IHrsbtwn4xogIWXjclOn
GtT+d3/+g7BcCKzjsiJm4Jm0JxdcDQD+VjhgFxunH1IC2lw1522GHTM2YClk
UqCm9URpbGk66f96UO3unNwMS+VsmkMW4qFeDoGZ+EwGD8kbH4TKVx09bplV
xecSn8vK/QprEbd9vDKmZ1r2HaEUwB2lB+HGbCLE21OsYuxloXGvfgaTsLDt
I6OZk2aZCc4yiy0rLPBOvnuInIXvcHBTKSEJRgpbb9RQVle/1Ud1VB8IEGCL
BIk+EPA9rPEVzKv8BbGwi2NlesNhnYk1TsixyDxjLzU9ruBVZAIK40ptRPYg
qJHvsPkfEoeE0asV22GrpzE4I+UwN5wbr6ZcY8uELZouslpShrpyfaH0E3Nd
2a9wrsaA0jr7VYXfNeUG8SeMrVWjHZfAuXkT2pcAJW6J/9Xr1dyk9xgqs4QW
wLw5REJdm0ZTYzFeDrrI0e7u6N8nqOVI0x4L27YqrUGwHaANfBbnE7lYtWp0
5Ix9iwJ6DVdYLNMmZzeK3TkpZw6a7Q7pkwquK0myJCViNuAebElZFBZMZQV+
n6D2QEo8ofh0dBFmOKe+HXdqjZeXML568+RvzsbCHuRolIPge3yYfuyVFBUM
7V7BLxo+Ox0Qtb1CQVtxoovpTFdf466/0HQN2nHR3w3x7J2SYBJzSmWI8J3l
PfDKj7Bx7znEvVdH5VOLMIYGoFhzwmbdJj0jiaDwkJ/Bt+h0kCNjPc4Kf20X
LAmKgL3qlzVBU8QXjzHNL2Xluz4ZqvT5lGJR5K/YsdoZfWkAi6xRxvtZ0Hko
4TUHlcZL7VzodZi/H/NjfEr6u2AbGUhoB1HwTkoEJY0AkI7AEsY1upHZDziB
BHSS1WlzO095QzMyV7l2Iswtc6NYAhEIls8fxVn/z5crimaJTIjkyWvlJ23Z
pb09ITWAnbtTkzodyBFY+U1RLMcQLopPLvWAfLUReh490/9u1RL5j6Laaw1x
9VyuwWe0UBni5KGmxtZy/k7gfE8ARkdzQYUJeYg0MAzbOXi0tcMhOLTVirGG
zmsEXBZ9KywwyiQoZ8sFca73kCbf58b5cirCalZE/MFbljesxDO5bbLfIjO9
maGT72txU2BIfGUzY99Z6PzTkJXNe8Xg7hBKCqKINfhhjZZjI0fmfwqyp0sn
u5jap7xwRdtdamp1a8fiMRPbXUsALQgPIfZjVBFoLzl8tZXyCQ2GUNcPeM2Y
/nisVLHFGz4vASHpbG4Wuq04MaEdw4Wru8qS1F3m9kI5z4GTYGC732yxANmW
LUD7nNVhbDnb25eag8tRpOpC2Xe15EpAuYKCcEr9vTKmyq29/M2VI2U6Roay
q2JOGvLa1s6J8veC6Rd63OUWaozy6xkJh+ZFl7NKoI5uTeU+qNNwrkxHeLsN
k8CNcR7xibl75G/OTGT5wHkgVIvLcl77XSLt4oFhMPYXDQCqEfZeeE49qYoS
cC6J8Ltomu94Z3Q51JtQIhwt3spZzZ16v5VLZS8JKEfhwlg7vezK0I+zgw2+
osayUHaKoGrfDRLytzO6IRp9RKxyotcBWCDVges1hHU0Y0e1HbMAqHfkVL5M
9ramIxvSBQBo9Z2YU3aPMA6hsGHNLOAuUtgE9o2xnA4fgIZWkkr72/V25ttK
EniqTIafapJq9e6iUuRO21l4vZlFXL6T0WS8WeYHKjiR+ZDkZ0E7lQxqaIin
sHDgk8lNrVTUIFiHeWUO7Fwfa55rIaKCHdotGVdMKH+jQvT9DQAo+bC7OUkA
GboGcFtH5ttvbU68sx+DVtIrkrMfuuvYY2vvaSWQSIkVczat7KvLc56KMuHa
jz3oY7m2L4XXr3+UvHT/RkK02jrw+MggF3sYjCcjw/TuG4LXeXQJ0NLFZsui
47fZk6rzhOpjXYZ9qx2OZQq6EN/b0VY5F57Q+leHrAqCGHTRvHJ+q1+wvSkj
fctyMsFDNUfElY25HBxYMpc4rDvXRkL4HRRqnO57h0Z7svaNN0mHHZBJPhe0
jReLBraGqjHeYmQoocoKbWtFXXBaLwoxbxaEPiFDqMHRwn5mQDLTH9iy1wyG
u0KYf+8m2IAnfJwyZw5w4khIlnSFo398MWFWPPZa2uFfijbITfMU+612Ck9M
BhredfYzm/HBOkAOgMWzpvWQS1PBqioaQKoPtba7uHjmvqmEHIxg2NNV3L2O
jSAWmykKMqXa5gfTyfUHcW1UDoyPcmaq9ita7kqIwLiAeFgcEW3t9E78xeom
hF8dqUuvSbgLWsovPDhkMbXfnaEoOpk3EkV3tinH4YrrSDsrjzDDOjoFvQWS
Zej6bfxctZPMJqssAd8YapDv/owiUzgtwj+bBz1C0+XmukmWjOMz25w+SEQn
i1KHpn5LZo6KYMGU956WijFwuMokCbFEFf7ZNO/qz11BxuZEPuEJVRKr3bin
Crzq0gKn1zDd31bRGmeqgryIcV84Kkyzznj1veVEYTEek/fiSBSggC5hSmho
AxaT5w1PIFk4SABJ+2hRdOi+0Xi7cyht40d+GxYsLT4WPM7aaLx3SgUdsTO9
rC77Hso0645jn5pVgUc3R0ms/K6T8kZsA4bamk6QVq7ILOGQTdi1elmATvYf
cG5KbqleRyYs+YI/UNnI34C4I9+ian9Mz6W25wvgmV16sbtulpLsJ9cSwMM7
wAgn07tYPURh8k90zW2XGdmRZ1U+MXG/KeILYMSqEPIvKzrGAj2tDbGOk2Y/
xf2OGtStj99rLyRC1gi0MxMrjQ610m0dqTQw/gwRMbYUcvqg3cAzr5KuOOWS
bwXfbtxM/r7ANhBL3YNdueLXyRbLUGJ8hWDZ6uz+hO45dqTZQZLvndEM4PkN
s1b6dbf7uuBqcsrt2se+whoft+p+WOGkeUPPig+crJIZi4sFdQnKEoOvoOA+
/c2SBOP2CtcmbS300+MFgcHfTZQzxqdbnkCJDBgW4lpJ+5yLu4mXmkrUXrLJ
ejinWnL3ix14FFQlFqX0EAwGqPEOkXLExwDTk8OhaJW2kJT2ZKwHbuN+V5Az
5CZOIz5FBru5h9GdWFsFVDoIXEX3zBcDIDlawvdVJ9QmQeQDDrFwAR3/+yff
8ro7wXZkinKUyEctMwhVjJ75IHJfmYkxF5B3BDRAKaPni02rFKJF9K/DOZDN
68/KDwJJEI2w3bSK5rIswWjiMPpOHPdcXFOlRmK6ECUk1ajwBlY9UBwClEXJ
VV1OV/prz70JuVmN5EpASAqrUffWcouiUwkIao+43BPZzHyQvc9Ji/2Xr6KK
bUyr+JHatliELfAHUoQOGucZnj8B1qn5+mhEK8dTAxo5Iqjnl5Q4K2pf4Ntz
itBMua1yLOz7ez9Rsf3CPtLwLGGOTGHRjpLlv+IXIWmXv5okPGz8HjV+mJE0
M4E0ToYAFg2L0+1P39YZ7wvHV/TyLrvdCIW1onC/K39ns2TGcOmnlpjLb0aW
OMnGbwItKHl6wbfjZ1GzTx2nN1GcMoRZkwyINsV9C4td9mr4VBeBRGlg3qFf
NqXplHIIiKd31ShiV6LrWOhRZo320nucF6hGpOauK5TByTozu0M3sjjXF6xg
jJpclFwcG6gGUhK2STQNQMjfNwNHwofNbihE/9I7MkHGuXXPFtZ0mFCaxM3u
b18OTsFmenQju3t5yp1aNRVqp65KW8vAhiofvmFKlTTVWLGfHVfg3wG3F5zk
txMpjMPjowcC+9YuA3ZGtNnf7vNlp1twLslI6e2wiBed/EWT/aSLdhhfrs7T
u5boZgRKjrv57zkhSUPyS97trveyfX+HsPmP4mvnJId+SlFUp3maIA3EMOCO
rXn1snwQmo6qJo/1jkTsHGy45JPWCQ3Czf+dnACi2Zb53rQZz1wva7JM+iuM
o6koR32FYqddgOZ+4/pvUwZTePhyL6rKfNM+jrifApLyfwoefneI7hk8N1eO
kN9aNTr1flGUqwJZW4TzaIK04ZIui9GhTuxpdMZp2kHEWyQdiFKsC0GFt9P0
lUIBrqGa4HmXBUeKaZufF/5kIkcG7ubzlhhBEbfCC251vj0vhLflsZ6LaqGZ
geoGuuruKbVIl/FiaOXnwFU/e3rjLhXxbhMcJIU5o2QfIVmxfzQwQNhUWpZ1
UB7jHeTpiRlrVmMZYVTbXDB3jaFxdETOgr72NNKrbznoSElxkhYp91cZklD0
iUZPzNXN2HzgQlfavKxdea0VZJFhkfC2mDEzXk3lUrPnzM8YK1bZ5WqPp/Mf
Go5fbCHYxQzIqWOj+kEODWtrq/Eg4wB1YlSWTOuFBASD8WIi7lOa9hUz43ZQ
4EJPLhITb5uWwzbsUTQsHOldbwwcvAcd8EbzflfrbRpAMYX9j1kHfKz/gl86
VLOY/Gzc51zzZIffJwgDAi0zg/Z4l98cYB2LZlIBkBAMG4pUX2dYX274/E7c
WYVFIu7oSzSQXcV2o1W2JijltPP62YbM6ZtTsRD6cK2ZOlR/E73/HfqBdYti
/3kl8j9ZFkz/V8h8CQShpP9fpQH9apXvJIUTMgtDt7DGPtu+Nw0bNg0xZu+4
Y/M0WxjLn6fnpXdmT2joHwxGOuKXiLU6k/PTlF5gQcT26E5eUKFX7I2Wo0KC
gwuAn7AG7KkCacFQ1ZUCjV4HiEAPIXhJrAMrOgTTN/0nV/LVZI18V8vBB0ub
G+u/6gox50QepjMv2TteswndiiBZYQ+bB5Olt9u/gLeHZ+wKHtzk+CxdQMjF
LhNXuaE8r0OHuCIeqDTT381BuuDCiBw9mU8wCBWVXVPs60xzGfnNbJEiPIVL
ouFso9S8B0cq89YfPwYOV30IijeMmQw+4bD0NtcIkCc4AxdbM5VtE/zfeUJb
79/A0ImdjrOxLDrDbFQg7adMvudSLVqIofX5Hk66fKF4qEegFMVjQCeHGYHx
7kj9GbRXtiZlvdXkC8gu08xReMNoN8O4+FOpnCzNsFYJ9hYESY/BcgiIT/kS
8LQqC2JdCgdzXTnUEzOufLkbLsyTwQOKhVJZZwyqH1WvsmfNSdtfAXXRfx5S
mJt3QYXmR2lviLkGlvsU/JWOo3B6dV0LaizYnsPY4glSlWkVfDqIj+UUCemY
fTGBlSj/cQbFfFHZ8jZhRaWgS68PfWlmW5pR/NVMLXGF37K07viz4xk8ZTCM
1ssVq66gZo/QXmbJIzwNz2lscF/bQvxeB7Ot1dKau/EOHljwFnPIx1Y1yF0p
eNqaByqbeDdn1l/05UgJ34nvolh2sYnnHB9jJJteiP1dzgwCgRbrI6+lUDTZ
GVjJvoKhA2RtuJmpukrANJ/IMMg8H/C8jxEwBi1j8GTtYK93QEjzhGz2dN3u
BVQLC/FrY+AqokuHC0HQ2RCUm+mbRhs4ILrWI6IB0egq02SfYNe4vZ840LWG
Oxw6VPMNkbLZAM4L3AMXLqBn0C45+/aelH8hdGX5tJHi6skNNKTX4zzGGl/9
FEsIHh3VVWzHMO7sjrf6rAo+8StGlJSDA29LlyDr4ksEBEsAE1aGSovtEq4P
CUlYsKie+wq/UrqGMdpuocB8HjeX09VPBSanC6KHrYnffsVqbhyeVu+LdwHU
DhXjf3ClWbtQKFPctApqkm8q/HQIMMN4vGaY2244CxGFQE6bi66+n/pd8tpQ
lx2umHR/BcGk8jvtrC9ecIcOwNXwX8mnwzSI+SaMg7zihhZpduW8i9qWobAA
J+0lKD6o3rs9Z9P5xekj0y9umrttbjml6uWdmBedTKkDYmeWjKgoH/bwVrn/
zK/AW9Cp6D089Pzhsifn0XbzqGfnPhLtdAbqpAmysjer1v1np6XJNGEB1oRm
+1LbavP01u9KHplajAdI2vr9/wtoPDZxxls6f2cdJOdxjsYenJtX7Mg/1wSC
RW4pCm2feRN09m82vdmNjEtOQJN596TBVHltDWddCBSIISnvnqOnb9Dwq5em
vmXwAr64c4TBRVfAG0fk9ObE69lmaeY3v/18xqcYRZhiUPBqbYyNXDdNp4Lc
iauyhpSdiBGeGJIYl3b4DfpwiXC1ISpUYzO311enaGdfp2xay9CSzhLGNPip
gPJ/1cZ7Q9HvGkcjs/tJp5WeiGWC0j0bqGicYAbboepWFqh73UHg4hlZFLwX
EyS0WVr/bm0diynlCnDAPrWIP8HkoOZfAX7QeH6LYxOJUHN1TQshbBqN7w/R
myQxGEl8QEv7auc6qS7L5Aqlp9GnoQSUJpna3qjR/qwtEYfylVLqsR2AL30i
z21gCwf8GNODe2UU0ZoxMB6TY5tWEpfXV/1HPHnKT/3gDuDNuikVWkwv8upz
pmPoDsj0dKFuhpOWZVYO4pJ0n8owJt1T04KY04+CQj2Xa8XyzZbcXybNnDs8
RgyB96MoKd+kr5DzDeDKlT9i+e+wigK5dWAAZP/V78Zb2aDteLBpH2Z6TixN
3h0stdhYlNeaH3zYl393+13AhoTsGUd8NZkGVVnYVnsTCvx9GAzoXZVWJLU3
hRY2h1UNsxzDoby7i1zsrNBF5Hq/ynFoiKs7Jpo6WTZ4LWmfG6csJ94Fs+f+
5JqMdofjIrC2jSKAc5HoqxhS54LJ9h9707H3vThIZOuo+gMJXorfgASCoi23
GTtYX+l6WiqQkFA8F1v2lle/gk0FRpM/in7moKahynOZQHUhH9+Oiept+HLR
RTuKEfDk0hNfMj8Rif1U74ogudPYaV0MiYIzNbMJzLAaUjUDnBzPzquQrtkY
V7FgAoP3An6msdC5TDO5vpzuYJZRURcvundQtlicCmjDXZCe/QGkGk5btm9H
YEcggZSBPr4xjRum5UudfVhURvVM2TQuv9EFN6ZTIMvUAP6UOGJwGAChv1yN
FpFAAXAwl4NVaoYzOTmDVjWqE5GgYlkE/qriRmu0vO6CSOA3lle0O0spmreS
wn2dmInqjhKdsO94t4wPEqldkWsL8DV2NLuqLgfPiJEETjOYVpW2rjbdMEP7
ZHmHrao63lVvVzOoKlcmashCFgN9UxtA5l9CS2tZ/Nt7V1ClWL10UhkfZ11h
ajWImbB/4G/VAhWWj7xBEYs8I0C8iMSW/QHsW59EfxcRR+ncr8eN9OF86/76
cTTybEwBMVINTsxspwNIhRzEAh1guc0CzC7wVNIH2z2Fe5RVyfyQGmrJLY9S
ffQl3fLvaPSGsoLsKyF/Z/QPWeeD8uNo8uxSnHPtBka5YHy417KrA5Z0Yso1
KZkYbiqlSKR6q8jKccnZEo7HIlY8hSdA9IdvhnanutqbJG5bLRp1D8gGSGQ4
LxNx1H/L6EGCwS5atPEqxhT9FxMd3LLuJNmA5oEGBOzgHtVSGIgw3dea2vmU
sI/Kts/hlKIzpvLPik+b1n4USMiSFeaZKakOSdvGPlc3B16onNQj3Jrr3a8Q
tViWaFCxj8E0L9LxQYR+93kQYXM1HikQNu/kZWMZE6xnnZSXrhlXhUBiJrlo
0ZFvjZwUBgpjR0VgmJWH4ZHjCbnUY7z7tSCNNGVzGabRViKmwFyV3GK78P3J
owG1pfbXXSbQ1fi2PWNEj53ARewhQC8CfWf3Qh7CzVTnoGI6LrOkfsn4vJEM
4mMUVvLWktJ76tcHENpetj3zknshw26wsuFlrGeWDzvmnFmewlcl0YHHTWEt
SdrVr4V/tZr7czMT5mE/cpROWAGuIQ/6WjW87Ybdd7CQ1tTj8uO86hrWDvZb
e+KIwNlqV9kEDxdhjR/dmeyU/4vk5JrFn8QCbKIWm13YKdKoLccufmlz4i3x
3PyUjMLTqs+jZVefQHh6TU/5KKQ6lhMxdzIEv92VvDQlSU6qctMiNEMBtPSz
Sg+6PONFDob4sxcvJVYzAh37oJWAfrNEPyqCQNFHATRjw3LYV6YCrnZyfq8l
97Mk0GNIp4pOdyDQPy7ox623bhAe5K8zJJcmfSVqZtN2EOKFSRA5ZZ/NIHos
wpCEfqgfLlLGUtEH7IBQ697EZmgzwMO+PpgA5TVkVc9mKD8guns5HofJtVB0
qL0PQcUmAwUQ7PazW0ucCwLzUvyMK8xsfSOFAGlngUXIZNgDPVoFpUqgtU4Q
H7dcBO1Jj95yiJ5pfN9UsGDzH4Fpmz+M7nSwI7Us3UpssAERAbdlfLo6bQnC
Om1VQijosL2tnLpskp5sHXikbl7R487zTZo6rgbymasokSdpJ6ImeF9KpA2f
BfZPMWhOs+NZvHHO6glhUwkTq9WFXyDnylta6LgPOjAdAvEFLbxdteM/TvcS
zlOut8KvFNIcSKKXqTMa2U20gYSUYcM+YtxIqYd2woTlbd+HbgVrVdVV+ntl
9BvPK0lcBVUwoCwLYqKc2dpBkaQjwLg2Hmm4BpTuF5E9977q0O2ITlvBWZ6+
utPzVZHIG+C26QEeqjq7hLEFnJHiuseMJRZAZmnX+yo4totxU7wMN794/V5e
ZmvhvPJX9FqIWrsjIe5f+vVrq4Wq2xLejTHpT2GGc1IO7pB3l4mTrZI1uNW+
a/ggxD20KPQ6uIWZ95GXmGxsKNJjx9FwmipQfSzdQ6v/W6Dzkrg0QeBcVqFz
2B+HMndIxAq+ADvIF06eL2PpIz3iomp29wMPmIPaiDeiIMVxqWncoP2m3ar9
JGhtcG8DI8aY7svFBo9+G6Z8wSH8OgBcYig/9rryr+XqQB7KeE1b6U3Liy1F
MYQEW+B5/n8U1MJraq7tJD+sZ8HKJvgskngFWz78NGDfuDasWSfYw6C2IMcg
mJMAjB1U6bQtTSV4HzUzfg5xR6UhscpEAQEhGS10DEA/sUknKZuw+nQrJjmF
86KktPEuJSFmZKjOMwUXK1UIzNXQDY9QbZLlkY8j0uRrVl23/VS2RX3iQJJL
9AU3jnHkADZowJu4GPKU0ZYZNyEqc6dp1BbUGDAwT3JjJ4m4bkDKxrKm2JXm
/jHCoH0UEcIbIRWSPqVkyiB55GrYm8ZT5217nGDJX/qFThHHXobBTbMS6ZZ9
VBl1/tEOBF9Phw4tAoGc4xl0oWglEEVDBQvQf4vMFFwT6dLQcn/TMfafAhvb
9uF4yyqZJ7es25Ywu/WjyPcyn6kBvrNnG0iTUdgJ9iXchOGewjS53wfh6vAl
4TBvOogi4WQ/ptXrYSjUDWO1bhQ86y4bE4KWK+sUnrsVKgbyCZGuyiI/Qw8V
XUCW9PDsdp791Ff/vruT5UYayabADVmfcZt1O2eOgD3uy4M+vjOerhP9QATh
3OtQTbvuXfXbWNS6ehAwAVXLV340n7u5jc+ZUJrMXYoBAWMJL6Oui9elWIPg
Ih7c52S6FN5lR3fNMsxzS6IMygJhbLJcQ9yQR/hWJio9ZqbCknA5Y2uo0UHM
1we9u6KBso2R3X2cuvtdQzIQa2HvGvdap/eXqeN7WXJ1fAU1FJrx0ezKnK6t
29Fxe3LNQFAHmPX9hWG7Kb/peE3ZAyY0tKtT8PDhW2iT81711XHpfaKcrRFW
A1kNGdUSs3B8GoxWRlN6m18dTSjpxXjZvT2E8T/OQ2xvPvy6dIOcLFkMDgPz
JaKiuuMzinBWQeRsfJy4sCp7QLV00fsJSrEcnPLCPCq8JR6i1WC+XZpNRv1r
l5tThjLY79HKihMyNwe0XEgCMMYL3HIeZzlRPou8IOqIhY7QY9Z6kEoEE1HP
9bZaa/VtZa6GGagamq3hs441O0cnKtzDEPy+T8HLh6f9PAlQ7+YqZWdKrTWR
YRj3+rUx7PyMN6EUpeQkn9mDBAC1nnhscm238QGO1YufO8SADa3RY2kz/Ewp
rqV3sq27bSnE2jnbjeZXaJrRD9Ga9CSFTxrNWPWbgY53ou/oSxBuiMFdGM8q
cbqBt0zmhp73x/bcF2jjyyqO/lhauGOfoJzkPi/ywHIiM4FTFHWEH4Mkfmoh
QsFxlDh+FqGLkKezf1YCYRBjp4qKFmeFN1GRsnkT3wDwZc4WCHvXUHkFN390
hLjeHLzyTGKuo0PuBfXh4WkoSElBYq1Z5XOlAJe8qRCfM/YBcl3G7ZjUb8lE
6FkODOS+SywwOEB94qo2qFAUYvyMRYKbYgy5m7evkoRNVKVa6B4pu9zO1ic6
C1mhdjO+G7YCY4qKLY8dB5zIsyZJl1ylPeZjFZ7EOPsMk7jZUE2a3+qWmk5G
UI4XiL75Xs+ZrITuati24z2rKGtEpk6XRkdN+CAHUuPQJq43i3/CDhDn8zHn
5Qy78iXMwSPVhpJjlOinNONmO8+y4UsPN8VK586PbJx0SasOI4mTSvgaUwoa
3zpuZsnehbza3XBPFas7uHwjcXxrvwSzymxifq64A7Ax1fyrnTJsZmRgeV65
UDo6uuoNP2D0GDa6scsyaXmRbsxAcntfEcbBbXimLJ7Qy6LGNmzLTdzJqBaD
SdSI1WOmn1uUdliyel8uJLOcQh8WrlO2c7TyBjqEeJ4vmb+SAAioa1Vkrsq2
yXYWStGmGgVo9av5F9vDhijAPxBJ28pDMmmXo907SmmDsH6l124KZh0DfREE
OG/6V0orQ8Q+zDco9eTGnBsFWKNL0CQQGBiUDot+HfQ0iALWS1Me9eKKQBKo
034CdcbO624raYU9FO8CFiOpc6FGSPc2tuMG1fXQbVgtop7D9yk9zBme8pYJ
s0qme+dR2T0V44VvYTFCV6lzBTwD1z3TOKMcknwPfNCSgDwV+W6d9TlPRVtZ
TFrBriKi5dTuPbK5gr6dEYoFigVqCYeVrLPXABrGSlB6gOLhI94LSV9LNUgl
u5GTby5Hl+X2J6cz3sGzxXOiDTbIWiQJghamCXEBT0fvO26ke9BIAuAzLNgf
yZmmYtvLfYaZQE7sFyAnlGe9+2+maS4LvKEQ9P0Lbn5AE9tjaM/uHRZrwKXW
lI0CeXRyOIFh3lYjIcgVqnJTNxCGPwNHI4YZuEB91fEH4DcuXky1E5JZTgUn
cdwMVBzI3gyuZcIfRRQs6h7IgGiW2nmDJgeJyJQjvhfyqztnIPtzgHM7+ihT
LqWebHec/nPmss633Ew+Amz9CLkbRRDlVSNSIeY6rXUe5KOlwfrDJEYxvLlb
1iw8jSN2I2XgcW/8YbXHVNeJrWM/wfkj8MWou8GcG4h4PPyiGa0ya14TeyzB
64ksyDkA/YJLOaDntdVSjvPSLm9coKEGy+yig/NRf3+Qfur8VgQ5TtkWJT+C
ljouj1ULFL/zdlEsLGL0UbWU/iLity5Kg+esDPNXIjIfKNJBPMtLQ5Ikaawn
1y0rknOTUTXfGrBX7PSutABTTAwLOs/nSjtsIgHipTfq4ndvn6IZOCI+Q5Hu
C8mmbO2jXAz13DrU0NMjjw4bOohRA3DSm8zQZ2JSz3gX0tAVnbwdIxngGiPP
p7BJTi9z3i96gaHey6z7aF81CiQ2Aj6WeuAksAf3xuvkQGnEdofAdyOb8Gmk
BZ/MOMUg3OwDfHWbEJcMnUcM/RCMQDqwdfnvJMMejm5kSGhyqyAzs0SJxwao
4H4cFj5iLwSxgezFRkM/zkbhWknTnEUkeLqvmVZkP955KJePupbldgeCINeY
rjv9Fyb4HpQoH1tw0I2MYHoKyKJI9wcSG6ntVsn4dgbIBNQE1inTf7lZ70kT
x3v/H2OEKpSJ2uYqjhu/1fZxtdwbNgPV+Td2DZcR4dSYHXFAJx/0jJQwoYXS
64EkoiAqChZ/hFtVq+04ysRYalGOLWmRZLRst3oNoYv2MXVdFNipFSfI5rZZ
5tmsedDwnuSYK0eBD+LLhhMxtaVWMPPrcneU5N7hEVQVJMGBGD+fI4YmFFN3
nHk9suKbk25JRESLRtADE0fycof1U4HoEjTUwx5Q6nZlNrENwMnyX3YSPZ7n
WigF3k345LkituEfKezfRuOCelMA/oQeMAzOCAQU77pQhapm1EDqbZ91h9ga
W87VPDeY3gvxO+hK3F1ffzx/YBFJueYr13LItmrtQgWCGGD/5H9ndldpoyIY
Do+YxU99DSk2H1H401S6JrzcOTxEClA3P5O0ey0/Cc3XpLYUMIqlBrQ9zwf5
xH06cWadWvsmckYltlGCm6OR1DswXcRR6TpcQOpsPSVWjRY1QhcnGorCqFIs
8laRrL3A7gIzDNynorlxswqk6FOto7I8zNChcV/SNfx7392dliXOoVTVAR2u
9FU3T4wVOj5xJ+JsnLoHDi+bPEohYEWLgsT2g/PLPLNv1adMaqasQ6Mmys11
jWDZVpeyu1Cmw9DitDn5xCVggugQOaYIIhVMQesXp8DIQHmXHEzSPHrBi1cE
pqWSSkqtk3lBVo/AH4zOk0mNQyv6l35dGmG3cK9eWMWXbykGxGdFztZt8Z0B
UXaPDVxH4VKhs2/mAQsdc1IQEBhCJHmDnqstE0smIaAEZSTBhEYoB7uPklV3
exbhiKBn9aIoHAQxzBUi6X6hT+EQHs2sDSX+54/5DHdlr9gDD/M0WlrHSQfy
7RNA5O9038atdFs9WYufa3b8bAiao7flT7l91/Z3wdoAXZg5BeSwWJH186wI
/01zoDJNhtszV3CzphBWue0k4ccyUF00V22+/VAdUouWZWaRByQZm4sOaiwE
2B0pTEAoPEFQc3LVvp0qyekzTkwxYSnvpGdBHGeyNQ940DDig0CYYNM3MBJ8
sun7gbvDHDFasOMhCeeN442zQUTQWabkpFUO+GD/wwhYtfdn9R87IpM2THKK
F8R9zBOTFJJ/p0l/MVAJ+cjwjzSp5717xXGO2dic04uxYpzbZMHGlJ8zK9Fc
12CiMqy2vqemo2YoEKpyCcvb28YR37diEi82XtCIfzy+2OiGcNHSxEWhViM6
bUcXX1hpfDru2UofKoK22I2jV9BzVlaW6KRw7XwHx+nsprBHtsVnMQQF3CCV
Jx9WZzWFxZyMfNzV8JfLSCub9Lpp1sx9tLMvPqxXeSnnSMYXo7UVCB/WaviR
Qpbl0EKYyC4DK8VtbR7vocV9RARr52BHEjEph0QTr/QpB625S//HKK9tduJ5
oIpa7Bfxqw6QgAP5EJKBbWT5dmv6KhbXx3T9EbTBHK/6lUkhVIbAK5JR+5Ny
+GNJkS7dzE/3jOKU5ywllpTTzb+EUesPO1R9qB/fl8PcSU6EHEuphdfLthpR
YuanRv/iIQ8SqbzYJXW44EGGjFgB2tAeMmkfwkK+s32kKAepNmtGcNDVHZom
nxf6S9+JkgwBzsEIlIcYp8H+FYeiLButXg4Z5eKxmCdF494zSQUrvsN+hPYJ
Y8iXxLGf6RQHJqw3ckjgZxjClQHDNPNfcgS+jHde7mWb6j9wpY9kVvPzOhqe
D+p+4f5lwCM47TA9Wv1coBba5qI4tMLfKYhrGhkH61QFMx2a20I/9XKb8qAi
eSr+bIPhvqZsv+AJW6gQNSNc/vvgiruTqE4LDh98qneQnezVq6dCpQ5zqgEO
f5kI2rwqyDS6mpFnegYUnA/RTmp9IEysNUMzi1G0dqyGTWBUwAEv4mHhJOiM
/mTT8k3gQLjfsRPkn6d1MPz9bjzy74NhvscszDMx4gIcFFXH0ediEJ1WsLQ5
NBneQ1UCrFQHCS9PdcrbWrWwz2NXf7Dip0q2bwuyot6PaIbMKh7ugiZ379jo
5n2mTwVpJX8vD+qkc8f37Z+apHDk2pCQLKJKzwB8SuW5YoWwBAzoZec29Ce/
6AAc4La64ibh0ADUgJQWTLyudyz8PQ/lmztmBGh29USrS7LjeS3oSbRQxjQS
5s3DbtWBW52aRfMixp5DAqMrwOo/cCJRpkcswsanXUlcnGM+aAx+X3Lwwxn4
oyQejOSyWKD9e9oL4MJiOvzu3QAYj30nHqD9x+ZWneHoflvb7IEd9GxWzfKG
H5JZVLGzJRNAGHZ68xdSF7Sy9UTRb2DhxR/zUc9E5HQh/PqFcUYZpq3apwVc
h5UzNVg2pshCy8KOi4VtfY091bllqkEBol4+Tr3PxXv4ZWoelPSAOeiiuBP7
FNvS6Ohd3S33MDbN1BfVq053CiNHVc1OhSPlZLw9tawLEgbNNHCswvZ3cSPB
StWVKd2Q9cNhL6UFTFKswxMLEvR2/1HEqQnvGRPRsHn5z03rXSw0clPMRsEP
GJ5GO2MlqB71uAsa5sQn4FrhnR2pSksiCvuJ5QPWwfy0IaPsuCc7e9nYLhhL
W8m0+zUQrtYmxZxN2E7OT+tZAlRXhd1o3OjNPFd9ITCrFQfd9FQ+KeNtAvV4
gx6OiXIpOyBMNlFGDt3JCPch+5q9+wYWM5Vlt9Y5TZrY1vIkaI2667WLRxxg
pCinL0584KlfzrmMtFxuschxiBxcD0VDd9G9n21rnSlSDFV/YDerisznx3Qq
vE1U0wF9yD/rgCdcEcE2gzp3wioWmFfoDeUL9OAw9f+JmcdJ9T0BXKW6Y/Ck
lGMaL8lbzcdQc98pWiApL2nc7Ff0h2N5nHNOPaEd5AaZSU9oJTim5nOwapHE
v26NeIT4F2aAwUH361MQYIqli4swd9DZk7ka5mWfHV8bYUbaMr3twzyr25Z8
uvh+5ziOGu9d4LY9D3s5GRU3ZZ0D3CC3qcYvQx8MDhZH/FqEJdfbU6CeiLN/
tUapze02Z/m8LnOkBh/wPoDgdl1ESGbGbeJNtOj1CknbhLGoL+JcNjl9TfLq
f0TYwr1X42sntsUORrv1R7EK2x9o5qBAghiy73fKPsaTQcHdgNDb9xLBooXd
heMxfbVjW076Tidv79s32tbufDG+jGbPeeKXVt9CxWj/wPMWobYLUlSvatRq
/jbfM9bbUxFWHSjiH4Z+f1P61j214SmHfTnDgXXS4gr/Hes3mYUAQ3oNCLj/
97GVtv+G1lgDBxDGUeQW4v+v39tOiYumlmfkOp3RcpL+vubtAVpCtkXmtmyM
tbJRYslak+sgM+QHclFzN3R88dI/FwnOpxj+qViedYWkf3nKosjcWbd+eLti
G1VzUrwgiTUUjHiIKEWq4POf9kczC2/qAcnc908Gn033Rj/aP1P5YtCRFJfx
FeH/ITza9OzaBB+KRbI6iUdmCTKMSQMspweMAR2C46g9ziq2cPiIQBskowVB
6WnhrJkRGWpIM59YuXLclXshvCpq46w0d+NbJlzH/0KtmjIuC6pfLtUGKcam
/s6ZB/LeNhJGhDWUWzTH1j3gGoi59fPsRKWM634zpmwjrpJMH+xYyUUH1Rd5
oKk5eLBSI1YHM4gnXgMlPPBQe3ZZpBU5BRYD+dFABwxd/MoEvY9fZNScvLHo
oVfPzlkdBrEn+221HUJ9CAlsQvH0EoGtSH3nZaN+ZyEQMnrfEpKK0j9GxOo7
4Or3yVPgi0EL+7TJhkF8zW3YTT4L4XzQKVprstCOCgL+plObI6y4Dr1FS4Y9
Ij73Is9TOVLQpqarb9PkiuMtIBR4jifSqiZn7QDp6oJS8a79ISCNBHWoCkfR
fM8yTESDMAIjUfpsg6zchLDI6FoIjvBe1yjElmwWS3t0zSZu9WfqNGIIYdEM
k19CkaxtyKV5WvWMU/NGoMZBVtJFRMc6unFqQDA3zXb9AA5oCJ7E8nOC0xly
RewDfy7jvrCFO4KYBtEKcOo3ykUvc4YEt728TC9tPkWPoS/s5r2YHhSm6yJK
KA7hYHXGgVBlZawPvFjwLPJoge/JHEgO1EsRYG4cd9X1IVsnNhSlZM1Clk9x
NBtmnkPGeidUGZJIAgQ5Gp1sgmHwHrFdavt5ghRRwdaBO/3ENZzlGZ59oetN
WRMfpy0okSaBi78I4Pj8LDZrrKP7qnsWYZTN04vz/sYFpg2jf43wzbXwJXqN
dajPOed+oRb1inURddSECrU9Od3S8jU58cvARV83/MbNUidaxOVXPFfc7D9f
XEwx9gl1BJN1y7Ga5IAAsJ9LECg152DDV1yySRfKLaR+ytAEdohnL29UJa26
KfHmE0xgnxAO0wA8yT5xQ56yrGrMfAdrAv2dfZjRhr59e6ERlFGowgOzrohA
IHnhkviqdklP7MyzH4UveaA34W6mWPM96Pf566x0J0tJh71jLj2fySGRaTx0
pCHckkbg9w31AK8tB8l0CjBuFSFWDAIHDxx7fkFev2uSkFjGv2cLn/Iy0YvU
DWbP44I5IEttdeCZ1q0dsBvd7XrjO3VIYfwliKvDRUx39zHJU8ZdGMkHVaan
odIyGoBnqfNgqj0oTPBrb/C74G3tsRQsFSTQARqdHXAMM9EhFpPnE2JyeIjd
9NjlUBSJ25+pznkgkVlX2sE0I1MfupjGGIDhsviP01Q86ilN2R8osa50+n6W
ZZuUCDuT4NiLduMDDkrkvnA19fP+hfHDudGBQqFrUY4YgPETNj+PCI81i+1t
OWbDFeqFnEoEU7aVjbAd1e0VjUgH2A6Odq3YbXW7Q/tJWn5ukyEUXGFtYuCS
CH8L8r2Lh+PuJG7X+5gI8uVQBzqLdnPbiCpFk2x7CKWZpl0jev1v+ljPqpAG
CE3yP8GSos6hQMeSdAk5e0RkMSAm0vfyD3/oVfGXPOLcWcReq8Tr2fFcdrNj
7JcX06QHMmGG8NKZ5nvGJpHLr6kctsamxnRdxRBy2VcfREZeBSJmOISlekGB
3E2A7DADp6creP8xEOz+ae4fKSEgfsaSARFVY32MqLv/7xSXpsIyEM3gycRz
UTxvS338nMP9gNFN0bbzX+WQhAhhUCwk9A3u0DchuYeM4vahAiQUkZD4iiSY
en4sqaVJe2yxVEq0YnBvCT2aoVGE7GPKosL7I2GVhmYBO2ac04JNJHvDKjcU
L1jpYIpi6qhTm/a54gJIqh1W7RAOFvk1cpJlhctGFO8FEkVNPMGZTWED8jiQ
vqngBczTh/5ouraZi1OTKvD20+TN+8W8bEU9EXRaX3q6Wz5YnocyypVCmAG1
kdnFAIw96GwjBOk4q4W4eZaMbCdvXAtkoWGNMOvhgKGlerPK6O5yTAjAKV5v
8zqg8jJE0PkR+NsUo+87nrF+fL4iIppGJsNUS/nU4dKJCCCiKBYq0lb9Qajh
TrG45Co3BektdRtSfllZoCGySNJjYDogdqnY+4R/X7BhIf29KnK/kN27IlQc
zmS21OaRiPwWl+qybwMOoVZ6cZ45OPmzyGHdzvgqVsx56kvPaFfOHSkuwiiq
fo4nma4TzIV7vT1gM47kNqEKPW0cYKfoMFgzL7O8pS4dIgcP4XZVPskcX00j
NTtDW9lDCJPXI/ByazmpVVDMM6eIoUFRxdYGB+DV1pAHaW0+9Hh1xtL86Knv
RUlWq5FKbA9vrIDauxAojjGSkvFXHybvUfpArtjAWk5iEPwc1FYfEiQpC6C7
t99zm6H6SARcfzNTBJ5wQkkVp+Oc57jxz0GzA8jVkQUGa5jQmPPv8mdVxuw/
hyhQz5Wjq4TWWxBLIDjdN2myVVmuSO88mz1G0KvQoUSUu7jAMReORMqLMxZ1
UTkFq1jsPWv0JOmX3EFDscpyRiS1Ixqox4mOW5OoK6oTnEj+KnY8MaPvdIgj
bsjJNUwzBM9WykrV62j8lF4ZNmiyTYID8FSYQEgFwcFw9TnS7pF+ID7J72dz
8tWER8RFOELunPIsGGhy92DY+3uj2GCf5vCs/JP2LpL/vwyx3g7MtuTLb/h4
FZyMIzhcZCfYR5nVtx1WsWWPbCPESZfFi1ABarcq9MoyIg1RafMLqPXKZHw6
7TIj4+EXCci95p6Y579WY9Mo6wgKdj2Dmtqd5Clu8Xnh1XRC8cprIC/8hw+m
7YK2NDA80K/C3lyg+M5mlBIDc4eW4ia1uIf8z20oNbdlpMqFDFl/YpmDeaI3
48eyFpf61exRLq3nyaTQ6ZPC50FI6k8yHUy0sls4Fz7fsTIMETwbg4zUmY0O
DPcmvAEptlZgcCCztzbIrom3zyGESHqq4p4xjRpeH384MH8mG4+qOFg7cLP0
0ppmMcwAD5grpS8L4Go4MctF7qZ619JIeWJtfSkmpDYNI/QAmLx5gklWKuKb
VYeluJwhWO1ehHhPL/8aGV6qgHiUL6trtC+6A+LfuohYPQ83+w1jw2rmbWky
f60CczyG8Uu2B2wNjF0X+Ov3xXP/VACO4rO5gnIGvILGVO9mNoSErdNQKai4
CTSPPhF2gZhLY28U4cBP94IUASe+yexroMiRhGkp4CFX+zNV8mHAL2zeGsWs
ZCPIgKDlv3vCBqvDk1PbZZncxXzRdJRjQ//Ijg+Pc52UmzqyfGV3okxrweyw
cDiI11dldaCs8qiwo+MbL3yLvzXOMSVQedvIlZzZdNEdkgeLvm3+u3httQZm
BDmo7dgVbbyYFxoOSOIl9gy+Qqfqtf1cj8+hCtyFLUa/BX+UHJ3MCWoWJoon
BsXK4W68AoDTuGbqAFSjFXtXYDXF8CRFNvPYepM5u5/yjqb0+emAZjSwD6QI
O5qPBxHGqVwSloxUXyJ7rAg1syf/FC4mFvW7WvO9nWAQaciqBg4cBO3wyKVZ
78AnaQmenSq9B4IbR1aTlVeKfGJpNy1ZXQW5PPGapNBlJIrnNNzutikCoXfb
csCiWVCn8xqwbbv1Prhf6Yp+7IIMTEWFbKYrj2uDsFvE2wjFLki3WPhoVrJR
msR3QYyc4xmRueuAo3njksBznrvE2kCE64eRnZRgv94tmy4QRYt1T0gcInkJ
4kirp0PyvGdXFlZP/pJuy435ih/Iy2EqgEiNJRTWRxIbF3OcNPvU++150Our
7WRoxvJ032uQj1e65dd7jI8BppLSK8Knsd9WUyzics2jFgGAo1qXOtgNo7r7
rvMm1mvZMRcpJi5Y6RLd13owriTU8uaUFLk03/EhV4QQE54dIJuSS7g04Q37
CqrvPd5mHZm4brZlFwdghF+fg1uY2Vwfr3R6WKpSyZKzt2oeydRAnjubwmLx
gNS/1W3pKwP2yeBPBKkaT6Bf7uXdKiv+7Qal/2h5gAmJ32CdC3o8IcMQ16AB
ZtqL+26Fj6NifhWGR5wzQWNVZjTjGVCA4iqcHvuEsyBKeReYyODsRN7V0dUx
olsQ1rgycoFetEjLbHVH9J/hrsHv/CaFe3/ObEDQMBHfCX2fr4galrL/3+pm
5k8sdOMpHuroyxTrXNneYsxI5MWJtpQTxepJcL8ZufvzSRiuxl8iCkFNkyHR
dE/opyQTtZqxACjKoBr4Avo7oNyYbcZWuY498aEIVyCGl+1zP9G6ETlRiL0w
OG1rA+7+evxytqLegUzkTIoxPQ/2nBnLBKNH5py0pUOPVsj0QFcL87SHIPMl
nRF/WEfT87B4nR1FN0eR/G5uC1MsZPTRyOW7WZChBKEdLT/4iKiua48zbqz3
7sgLDXCKUKLaPmad5ubC5aiPTNh9kaEgCX/NJeA2CkQhRS9D7f1xRffvbZzM
P1tcfTDkmy53ax/f8MVF2bRlZOaDY99cAD7T1JFhIGPaSPacFOD36h2KB8aQ
zfT2excXqIp42lslGXmMcrkKyzIYIw+ANLuaz+RqUOr1B98vw521R9ilCKjK
I1rcGjAf6rv+hjP/oVJHmikSm0x5x9LVJvGNhnDk43emcFLWoy9BqYnG+O0Q
TwestDNfEzfnrplXExZQMSRQ0pCzg3HpIW3B4uhK14j0JzVS4oql+N6qonpT
J/jMXAB3emLbjx886WetQvQ2iZoHopKJSs4FeMbr1+ZPZHe/y4fTPzkMh47x
QMQjc6c1def8Pr1RY0juQMMh58psgnJzvNSvhvxsxP0rpnAFGhk23djvAuwz
GMrTN135Snb+UPYAL13mspJgujf3w8kUSvalMQKwC8y+zzRsbhMn7hTfyW3Z
plmPgQ5LFfKknjCMFYDaeIi9hbo6rBdvAsUr2X69/ltlu/9hRW66g2KmpBoq
IF6/lEy+oAIHyvddDdUlRjhAevUMIcyeuhApxBPSArOwCBZ1YlrBqGm1img9
mJPXCIauC3uWNcZ1cixqGcUcU4sv4Ep84VRErzCUROnkp8PZ53iBHXOFNXrX
iBaVCN1FI5mRhtZMVqcUBD85ic8S5fZ7B3ZekbJS7kY9AfMVG+wNKMkVJ3By
xX+hnAdYSJjlr8i7OuJ/3QiyAp+ijMDMCfCeimQuwXg1lfVIrJsGv/3P7Ngi
2CV4rMwDBHl06tt3FiTo3oI16nHTqzPgKFoWECd3ygMWGDxFUge0Ul7pPcmH
6J1wJJDZfAj7rL9/VS44NRE20NFseC60flEXquFyEXCPiia0JLgFNZly7BCX
AIAtgvDsc5x9AODvsSPAPYy+k5JncXD+a+takUhev+Uh7CW1gHEHC1vyrFmp
klfLF8pqeS9TE3mHh7vtrXZR0wICHaRsfeeD+935wdSfLqb9XeOFT0+sVES5
gwbuhp99kelZBScqGuK6yTRaadqt+mfjJVUQMHw/z+1QmPKUiy9TNDo+wQda
VrQmu3eTPTod5vXFz1aDepfevwUPoefOMs3LGYKw0arP5A4oa5SMdsszFAKD
4HTlCCuLbaXMTpAA5XTVv7r35VMpZSCUuNaytQfEBNBhXGv7zp6hzVr1US28
UjkmlSJAsvoHq7epeES2mFxeZesYGHRL5Xq2AZgPzVkFxuPY9u9JcnahOF+D
40Wiwb/2boghXdFyHJvBNbRKf6RFb2uXjPaz+uEvwMwHCiiw5jPWLrWE1Uzi
C3IShZzYFQvXcoXQghMuSu3ag4vkHGbYyvoriwy6Q4z9ljmcvDyNoMdaacO/
MdqlwCYbcAtqs+WILQbB+6rSTFLqkbb1kHP5ym93qC3kr6LB5IWU3VeZMeyF
CcuDdDaUYPQIozpySNUA3ASIK1gwEayURvSdaYirY5FuzlBYQtO74BbHb/hC
JnyU3d8k2egd3NY7Q69gdsTGO0yd3BGQ4i6jW01kAQYOZY012GSDDTgB2AOj
q3YxmYIZ/kP61+prHJfCekEth7vSWJPBBAomcf8cIRccOYO5QwkucJxCQgYy
NH/69K9M/6Qq/O09ED9UCiIvYLqzbrSu/Rm5TbBFa21GKHWvY2AI6F/vIhhP
6kJCYaZiR9YWYlRZgilOhwmVWz/jS5uQ/XOXW3bZtA4FHnMwIPXvSjokvvXO
/lgP61PBTl3M7+gs1wQjyosN2QOq6d+j2A0BrzpNfYfvRrJG7qpTDZLdKWFu
6wTlSUhEhNBnSFdgXxlYxTXDyLVSzlQ7pNTRQIy8HvSDkBhMh5oCJmJJSbay
Od6lDlyKssgM0xOHFNL14cxk1nbLBstXoam3yU6y6nZu52CCd5LyCkxQrHJT
4cQPMcBK9GKIlqrrAdGhGr2ZAnhFdjKzrezncmHDbSThVaw1MG8YZR14Sf0i
IsweIa81WlH8KYt0rEsx74QVtu12eaJKEMD0rVa92XUWRm7Wo03xlgMUziRz
lEpxPmE1Qkmo4J1V/SptJUoppP+EyfLlsaQvPvKZYzY4AcaBRaM3bnL3zu++
Yt2w9yw6Ex75RaS0DO/E3NtA0hl6nJssjdUPKVJncuwxQSbSzXdpVvxZiqzM
TNsBOEwDfXlvPSMjrXwkcNYh42H2h76LZiHl38v23uULxKmWkX+bv609YCF9
C2Dijc7idz8z26ai9FSQlNf60QCOHXLh41/DTZ3597hOOQjwuaQAYYYfoMhe
wp0pgZqyxKDTxT17ecOHqgQIfX9hsUEgxJFibYNjJU6DPqoTNrRBAXntnd6O
vDGDXPThBdnUVIG2+CXuqJHz+hHkwyT5X0q24wEXSN7DRe1I6LgIA4K3wL3/
y9y7VtD7HifT5M7Dj23v2TInw8pK3Cd6TkPBOaPRWuEfeeOiFZP8fan2NfVf
9BqtCjztg7jBg15AspgkvOz8BKho4WYkz0DxtnRNkfVDw/8w3paIaeuyhc4z
R6UB4MYSHxZyYcuxIO6keRAnfi4wWSr6RD713oRqlJISXTNtIhwhz9UjeUL1
9r0BzZxkhQ8W+LcI7RZQrDW2jvJ69oBHnY3O1t600wTVQdhVXdzpAZtN/N3d
gkXLZKBLCKvW+tLa1Ey6EOamIkBtAgoHsC2XcYEZf4G/MEpAtX/XJCXkYFnT
RnhlzCRqNRTRYj9IhRwA4E1uEvPAqjj87tTbOWNvlWjOf/qojT8ERPqdECI1
sWWB1EILGgHnRCZ8IA14DIoc8CXfgiy8Q+6dR9MSVEBQHXkrcELfRUsYefz/
2zZhWTXlukEc8GBIQgu7vzqpq3t4vcVDTmOPlNJc2pbRKrK95wup8+KgcOif
gfiliIY64OAJYc4l1JRa3u+sxQWH/sHpQJK6VhBMUQywyA1AJY/Y3K8hKsUZ
21Bcc3oJ9eOVicWOI+urGRe3CxvXmLlstcFxwjrpMlZxx1lq709rb8mdtZXK
oT4W+GWY701sswk3VQvITeIPuYHMMP6ADZo3n7Ux2UonpGEDLvqxY+HKMLrM
IJUZPh7M8agfDjdV/u9ZQSdjeDEk3e/+EFJuT1EhclyUL6xvK6uGRMkML438
EI2/x6u7eWP8vupeIvkz00d12jQSJ+U6koO3Kms/jCc8n5fqQRjtJBaNC7CS
fF2L96urt1aTNTU2ZxE0vR6B59fC1SWdAon41kSlxFpWTJbc/cNusUiqKExt
1kh4LW91XTyws5aMclzsX/GhO8ODJN/5oofvQyy7/Tk5EkTr7N87VBTtSImd
YxGx/quWUP4LCSwdnKLK8QwZ5cefvsW1F3xgD09oCE/TzAx4Vr123eAHFLTu
ZeEKw+lPAGwV2ajMUL07NCUBtxHWzOGz2n0PsBsy9SeUEUOTUiVp1+n7O/SJ
ulbHt0zlhAG+rrZzQf+NAQLg+JPXPoSA/F3VUSWVh+doZHA63kQxoY/Ud/rb
9unV3exdDAnOMm84gK7+qfVPlJocTgsenjxdB3TwK7WyrIxWjkanuhjzkN2X
tCqceGtvz++xi2d0ENtI7cYA9Df9hXt49pQARCPjtugxzMfeFxq6eZRcf12T
aXgsIoQcroz+/XZb+QkALIe/4F2KclOQsqlWwz9YKDxIRa2syIo3aEpabJS+
IvB17U4wRkXewfJdg1+DpMQ04CyMgSqfmuI8H0sI8VQhM0wWOWhIw3fRW7Z6
jvymeWik4Caon2CwtzTZDQ6UTg+cP31Nz0k2L6d0EScfUuuJkgHDE6XUQQiz
N2bUHHD1fBf52ZOxy3llv5dgNHke5oPpQ5dg43RVYyqVhjBRvnraUPeImljT
lGnSyxCoTg+CWvK6yg1nukHr+ce651mgRpS3fXSTcXyWBCBvE5I5H3mhsi8p
RoysTwP24bvaMUAmkLMkl4J523WTBT9lgFMhMGlWMLBqnUSZIs/JvwBoxs/8
J0jtbCFt7FiX5eR5gpNlJR7SPv5tZbby9fq39l7RXw4NZ9FzyIet4y1XqxNC
wHCFKB0hIb5E73YJdRCc6/xZ7zIdRlLcm8cIl9JhpclaACU9OLxm+WraQFwB
OvfE5AOfXd8aCLGqAJqdntpRLl1iX65tB0bKSxElnA/OT26JTZ/gPGt6klmp
y9mzxe/ytoO2T9gzy5uCZz/PSVumTnmZ7ZtOizl4hRIkdPaPI0sJyREsSBCB
nK1zk914ZCJdEBLbYPHFd6+v1xX3e4AnKJWvhqmjaOBTZv1coOmUWj9aDS42
s1UJJmXublRqWFXFQsMdQHXyhhISfVzKh3TjLh4A9WrKNEZJUMU888jGJSlJ
hMgm1SLGP9ocpv3pynWnYb5Kaafhaz5MpJLwuQxKFc8P33/slQtEa6F55tRI
cNx3VTR4Dxmt8TupJ2KEw6BcUTxBWIkxsAMwy/TRzE8ypQF7YNvbdDv5nOVk
SeSIenseIU4Aby9w167VdYBeLF+Vse0jl0YU/3XE8PhZJYIm3KZLWsW3rd+Z
EOaD8Tfy6h71mCft2tMCwIdXnEwB8qK7GBAvIBjANUuD0+WPrPb5q+0N7cDq
tiiymLNOb9zTJkAEF+Ai74VW9vEE6DWSn5iiohuhtXsavJpAELQY4A8X6pua
buT9eu/kEuB64NXrbiHm9EhYHAjNcvlJDpFMBRLmeKBhWNA/N4ToObXZZ5gs
Vx2Ki5nX/X+KY9ZXAxpjh/J3fhNu1GA4TB3CKOXZmklgYQGdudhNCa6RNzUP
mdRG9FviX8mZY+457CJOfUo9c7/Mxs4FeGSh1XaweGWI7LCBvvfWf0dxYBOm
WleLqeGov6vhBYWGrw+jB/mAw5sv5uY4aNrwTof+eU4q5mqDQBiW8Bl8JdmI
mVAQ9DpKaGJ0llEqut9APcOTi0QRPQT4A/TZNEZhIbt4LvqjdmgEZS/6ubdH
Uk1oe2h1bBCvk0fMO9RX2PaYaQa8+L4BokAmItdGhkKy/aVpPRafjxTc0vx2
d5ZHNrJ/++lIqmsnLHXggMfpGjqJ3l1VW3faP3JEBoKNXmFItusKAjLaZGEm
6rsvDiokze8hfchSr7XLQX94EGFy00lkexVrfPA42PXzn5oevCUS5Tkku5Yr
ktv1yb/MVY8ZKGypE4hILYV3JVPRz8p14efGRrJCuiQQhOPwIZqSKWZutEiH
wOouE3OIj5taBa6aaUWO34+WdxkNRN+FY3JtgkgjmV5C1RKy85nfRUNOBeT/
iromkn1lh/vdZSSP5+XjrfZlCkC7fCVM5qnl3MTXw95FFyqs4PMZYMVJWApF
HyHm+hUJKsZZ+KlG8/sPwpVJTNhzAuysbaazTFHL6mqQR9czV9eMjbWZV1/+
wcpz/piiiideUfcTe8C1t0SaifO6qaac5Xl7vFREyYCRHzux7nuAvw+1x/ya
DbSI5Ob97YAe93efvpeAxgDYKd0LC5GrtNMdmyAAtVY52vatFM9n+1KfY9Ud
a0fp0sShFVCJtYf4YVHc7TnWQcth76AYYAxJ2zmusMMIW362xsjrPHVqo5Dg
O9oWEoCAXGxQy/mvVUkwC59jpS0Qecfssehd5MEXeV6X6nQxasyC9bO1fjad
5qYT3Rw3sPpqkIUUYaq/7npTgB8Jb/zQVq55xm7NRvpCtZHrWSRLUkj7Io9S
pXSjsnpMLno60r0x7nLQZmneTX4BX/oGUQ30FLF3SZvaCZESwcj8lvpuhwQI
D7jiFE0kdstK+cY1KGA2IT1WQomHBeBifaKGmP+wC8DKXiRp6NV3YM8iGBmt
EKfHDcEgbanw9g72n2AnMupty8vix+C/OKcbAwzpXNNVo4Dj1Lk1/6y8Xi3s
PrDcxAAGjhyI7tELFeltZZ5IubggZzOPI+RFXKya0ykrBQt0vK3cJQICWUzE
LbPEja6g87WUzZtT0zObcxNvXVLSqx0Eb288Mt0s+Tj0vw9+4DPr7ShWKPHM
NAOuy8EGnb+KaW2QkWdVQgwDw8uOoJTwk5QnnzjJI5oEjiM+xb+PyZ65rD3b
FSvh0HT1/KABBeldShM+IYmis54Y5SshE0OVFuA51oPeEF4cNIuJanaMuerB
UQrY6IzlSJw8ZS//3pORlia3XwA/r7oSZvD724tCbkoO+udj06SaqnfeZl+H
peQaiyJvLQAr5+BBiR7wVMuw1dqYx7y+VCSV/dpLmmbgJEqIYsI3dRPKVZla
YOdenHHtOnQBa9nXqocZ3GFTt8GIwBkyealPBrPUhrPSN/4aK7E9QtME2N/y
qEllbyxaKZ5nHcv1AonCO3B+Dea4mJBfuqMlkrZlfcZNKM7KLtWr3ohnmzuL
gUIm+fnZqXNE8aqHvgQAaKSsQ4ExVG7kBmRgQdgkTrIRWa9s4NyFZuDqSk3Y
+SMtiKy9XlPyoLi83wft/dgengmEWwwlM3L/pFNF2D2IoEf9MqhDMYFGJbhg
xPekgwd6h1IBWBANpPHflaP3hPwgVxL+mxETWRddifw70HXHUXCBSvktLWFw
x1JwJ7WshhzuyYnTurfyfQVHEw5PqXhhlv1cO4etDFSrzD958rSYKIARFzI7
eJD1aybIf47Qpd5xDtE7KN4gmAkiz2PP40iI/cdGT74EzY61dRLJuKmfZLlp
ylie7x3Bj+KLac4ZOnnm6DqT+wQkHzBONah5w8Mt+zFokgH3bPd1HpvpBWaM
l4vUFoqQ5c0sweGDh2qoBgPEBIoBbqCjSOYTJromLmxlRsmSEz30mDH5opyM
sWULAuxVrEp9Eol7S+Vr5tL6q+hmRpB+v9NbnOjwAUHRzbhk09X+7OFHsMox
p5KwIsLkRCUUGH8QrLBU1zHeGw4Z46pflK0+94g2op+5197x3qXc1vHCTnu9
r101vYcYWq2TAeGDyRglvxJXpJ7tDctALQYcWH8W9vWKc2VONB+npJH3rKGo
JRB4Jk8V+VLvMHVxSiNxh6BBIu+h74e9f+gZDFRr2yeOSXwegSRbAfo5oWk4
cM7UYMxMmSBeo3QuNhOhnneVNZCn/yC8/OOO04kfOdpvkBiYAHTvO1YMIoQP
59IkX/cOwWB2STEn5oBJW+h9i+ui9SrenDji/LnLY+ApoFY0VKNse4doQzKk
LChNuHLEjLYrXw2sk6LHBaDUjJZLP+VLkP6h7KmoeiNpJxBuVlosEZMoQYcS
8h6MLzQHjMsXY3k+044lf1nSoX88Pmw1V/qGvACh4F00jb55O4ODe3LTN5oH
b127WwdHao6I3PqI5sMDBc6IHSjkUKhfQwj6+9uPowTnjrMeBVHTbes3BR8S
VcplOraATRtxMnjOksjABDWlIf+tdzbP6nqtuLn2X25JZolaZRDqzGdXakKa
4LRML2VyyK/BxChExt3oEE7aLWximllPACLd85yq6oZb1GjGAsv3WSi3lqXC
7uBJqBlJU16zNZG0qok3zSBO/GBpmNtZotMR2T20muPHBthgHdrMZEjcEOeC
XDbPGd+sMARFfk1HX+HUD7wxFBoAzWOe5FON4mwA8ZNMxe8bGFwTKaizIK5l
7/ogxIRwF/opkcx1Japxsb+BmEwHcSG8ZPaJtIsAVMvPuOaBq3DO17eIiC3Z
kwwMiYNnD2l+AwoKHDduuotNTlqQxOstd5qrMVnhXNN+LI6yMkrWUf3VDw+s
pJQdq4FFhYI9+cEwSwxUgG+UkxarMK2qUbP+qdSEim+tI2z2FDXdiqDoWtqG
2KgpJ8zpDlI3wd+bCjybbstAA+eqGuBoOQeJx1Rik9oC8KLK5nS2AnXZmBSK
/VA9hi954yz/4y9HRt2aV9nX87WHge5OO4ghtWTuiI+USCrVPS7w8utxoJJc
VGWz26gV1/YFofzbjyhVCkfw5dDpjSHoDZb73vowhqts5BadPPFDyWn2VmV4
NvphbVS3OppLZupvzq2WDGooCw5w+qW0Y/M2mPMoTE9pWTyQ/XoVSJVgp3KM
/5NFzfmfdQUUHdym8h1tFLocsfeO7I0GJABORT+/GwSXpvoWjVbF59CTM+xH
sBAYj0cqvCUx4b6vcv21SMDtojaZzoPO08a1gxOpH5PH6tGVSggb2Q8iRux5
UF96MpV7NRXYNKaYOb7nmVwCmS5eHmjhL1EPB/AWVufXpbOuduLHBPCEXoSM
ziOU6p3ibKyAYkJhWQ5jx6/7yVzBGIHM9keW32CgKc0qRnBMmsxsEgjJbiYc
RdppTkt99ARPdHmXBygqyjsdzjPR4sSWhCn0AfswaqdVH/oanM6BBcnjcOlN
+fhQ60NZZ+r4rvNke67IX2AvV5iyrVWfcmvX1+Iwljx+Y20ToSCJK8t3/bV0
ec8mgUbdYjZ6xUBc2xmULtDZKQxc9LfrE9AheCez/5QP6F28A2uLy0fsOYt4
7rjwLj13dCzjPmIsqQIsLTbQzUXQICn60CEU0n3/sKvP3/QKiIiHZ+9dufnk
LZ8eOvjiWS4P1e0JLAh/kInLm6qajOJjJUFs7YuqczNWsgDAJbyqbaIeXwNd
Ds1yi4bwAC27w1jbXqEbYyQqxqhhYjtVOFgO5G7wRUeEQnhN0h0gGJrJfH8s
KanApU1ee5bhdeR99AIYcHnZTnfETG358/pUM/13d/B31TSKmFWoF/dkq8Nx
fgSD8cTCY/GR9lb4uk+gZxoyGXc4Q5OHGmfZraTDob1NAFrncWUwtsDBxi2R
v4fqLQJZ3yhWhJgMYEO5UIn1d1Rl8+FrKJzKmVBhLqLz7tRYUEulNkf3xxPD
rbv0N4F8G7gOPbL/JHU3NtvLyBI+TbC9KBJvqHNVTF0AjzJN6LpSdoUjQO6L
7ZlHHUBZWSQVo4+T1Kdn9L0JC944VKpY2V00eruLWAtgxHP/5bBbrAs6nRTV
Qjs2A6jvFlNO4oujEeAhVMPI0MOw2IV7oR+lN8GFFSx7d/fVWl5FVnzPLm3O
vFTqTR95XSFBptAmDf0EU0TjdpdpWyv0n43syH31TqIN2nHLTD0n7rsobZ/1
wcr6eDfb6/umW96ll2V1vfhGtPvmH5wCv9nSoi8bNgNLfvOYAQaMAWH2D/3d
lVMKXCxIXtB4lX2f1ySPiwYcc1lnLgLLWNNps+3VpAoe+sNAcV9e7AwuRRQq
VAtKU3CtyhQiPcv2RX2TQmwSJl9YZgRDHqiNND7eQKhyoQijsUmsbjWEfb6d
37rjfnAZoH5/mxIPKab5QABg3Uyq9HZiqQ9suuhQJGXavkScZuE0r6XXaAxO
Wdx+rtSv5CttfPWKMtfazHwecxHVi6AVINO2qiTBNOs2mEkUgz2pRo82bn6t
R7QfW1CsRmyzjAqKcgFAmVhTjge+PIjxta4XsDJWl3vM5b9Hn4i17xDy+1Bu
zrQ78oroHo0eNKeE8OKhhwFSELWkJcu3S/YdjBxPAdFAkzRH08LsL7UPHAtX
OzKwdak5GzMEjD0ohua+zy+NdgziJR0eT7BqGV9kR/50Don1VLw/ppP2vEOL
lk4jbILLgnLdXGZV+i8R2p9RFtFzBJIQI/xb4dW9cGFprDUMbX/mEueTnlIk
PKH4cTSK3s3mlHqOrXqdlX7d9Ekf6bdhr1je8ptCqn9jMBSCfi93mAlZSfKc
v5NXKudMR3ZdiF/bMuRe5sXVMEmpEzFEmBd94NxB8xGMGXFc+Wl1uaek7DHx
Yl4k7p+ghvK9/GUeGEuCpFGbgj2RgaG+SrQnrnIhMHuGQyzuqLeAyMyR1LtV
PhacroqHWfK/CMmTBYnlE5Id5cxRZvO/vXA6PRoaeyD8q2GsAMK23UUqxZ8J
ddmPkqVa/rv5uI0AlKGImqE0JF6dJR317rZ5a5heNGwzo9z1u7MObsR2LV2b
TAIuDV6q64TBOLf4sD1oxRvOusrujavC92o6CCODndU/NElUbRf+HBYKDfgT
KfWslmef3+4cDb+MLGaZNhyuRd1FPoidA0LHiqG1HFaUoUqHEVRl2Joc3sUd
8Rpubcivdv6ENLRYX9eUo0QI/AzlCNy2USj8uw2nT5YjM6QqmFgpN1vbmw6z
Qg053f2S85hDo7u4z8/eGn3oG5T/sO0de1KQBVSdpcqg+dU7VFZqscSDuD96
XairHKQyZXoc2yKge7XPeI5dIDlRRPZpO3E3I2xbcV2VaIguGRSc606nLjpE
kw6UivGSnlU9m9Zlg0oCGl+iBs0nFYh36EpZYDiUyV0LS6fU3d0ygF7JAC9b
Cx1iRAdfB21yfEyZ8stBNntup0XlCd2igh93S/ncKWLKhwEhx/AMwJLCLqq7
UVcubaNv8IDdYX8fR0FrzX8EoiEvl+xb9t6rKQ4KCBNmZavxqhyfVG81Q6cP
DXqq07dhPLIyOCOGdyARf9G6ngHvu8qlPdSFbOn46GQYEbWYneirtSmoiHJl
iaT8esp7kZtikCrJ9Ar70rCzMVOx0oYHqwaLDpjd0dUWYNgLg3Sex3X2SEam
3Dkrz96JDBAQihnkxwdDEZJhsVycVsD6xv4uwDrrJ/O8AhsZUqQ+UMkpyfuP
dN9SD37BCv0nEpMYBTQapyTAVLcFOmete4psPjcX36glzScqDNNEqlzBqAt1
cH0HF8jZYa8RCh4zB27OjtzwSGkz5OycybVHSoQAJkJbqMJZRfZ4LLuHMkex
rq85m+VXDz/6gBEC9TDIlGeD9LpUTaFA4yXgLUl/HkC1ag5yRqMNHa1GOdGe
bHVEBtFkCTdNQfG6chML48JUSMnMNJpngsFe9lnavnVm9/MOTUapCX8OZ6tt
Q5pFwZPNQnBXmm0JLd+colP9EguPB9S9jsdJ5MprvDh5eR33KaHMth/4G9I0
jRx5lI83KQEOlZxg47uY7EQmOfQ5VZFDqScplAy15k1dpUVZi3X7fvJbnuIE
cRV1WEqOfgpW6o3XrCm8QST5vRmVGPY0m8D3UGx9aBT4zYbHrvdtO18ewluN
LS/LgoGawLisUP4JAnEtZkXcL4gjYuaw/cvoeKRdhp/upI8EbzHeE+iQwaAF
5FfR0szq/kkR3rjtOS1WcFR0krAZBBGCn60UmccgUBDxZ2U5pYo8jOb1dI3p
aHIBD8gJVwpP67aQsDQXdWILlqVz8LfMpuMNUNTuiQxV0GV31FVOVNtaq7kG
Uqfh484OagMkjCH915QpccTvCVbFOWs0lL/UelmMXa5RyVPueU4bcMRG3elM
o7W6ZUlVSUNICn4m0nIiMTp0DWOhF/jQ4o1zOElvu/4GMVutjZFS8yi9avIT
ZlcbarXUNJowdntOwUOfizZsItl1+h+jZYmKBwvG2bruMHP/zfLhWqlA3ncr
ZZgqdxrdM8f9PBOyjNG/B/Mhb8ZONS//M3fdTExefKSpwWC3HIMbyUWXxE3g
HQNuyt9+iJjnNc9MctMzH1gfscrKtcldGsmozUpeXrNbETxEroihiQICCwLI
5n9qrQc1YEbJOm9lMq/UzbDVOFHv6bB8H5ur9Vwyzhn+iLpy3DCTZ763oDDN
R8Fk4MNLDAtthlWStxPSAfzgBSpS4dvoQsX7h7ylOXHtxAasY+7mBL3K1pji
Qo4P1aDo1LviTEjWXegw5XFSV+C0WnRuPi3Y+0jcm+MLOB5VfRAKx2vd82m1
qp6BKzscgWgDAsIIuFBL/1jioD2N/T+S+hlJII0f59u712nRAa5UKX44i/Fv
3UdHW5FAxjuds63gv3RO9+bJK3nHZeA+EN0wOkZRVQTNpKOOyPxNkKyDLi/Y
BjfS33VToK2EQSRkY5+16oQDdDg5nr8gQjmGRljdTVxM5/OWnPctUm+Zp0/P
s8BywbhS4p5DvZm9bsLhPpTsuyifA5HdpaIdAqkrsUKhotiK+BQECnJOpxxB
tw17Ng3enkpZmum3BU1o6U02QofPXjKo+yYgnujsGMgkWqJ+MfX+bOiKqDzM
/mVGcVHg/9FY0CsX/3n3Eilnr0POcYJE6AmFyqla1dWeI1LUHgEXgkhMQ8H3
pC8fPz7mry1+ayCbFdt85HMooseT+AmxaIs47WUKb9AtuLavVH4i+S5jGLLz
3v3u3hA1uZzJ1lKtbxgeU4fw3sb+lHQ4C6AJnwCAeCEgdU1W0FIDne/7HOzn
aTuGEm593UrnBFRU392/6zy2FPQMWofmF4m7ChCgTT+6/1j5LD1LixKn5RYw
j9xwCmnjeP0Tomw/sQKbtZEj/9LqzoB/GRJzt9BGMrkpQ+nlChO7s51EAFRK
wIy0BNBwEDNcpOzQLt5DJ1m/KBDt72nRJT8/89SH+1JTnZeux+50GOYckydJ
9XwEAVd+XilRtqZXUJhS8XXGzIxfLzcDb9no51sll6ZrpbC+l5NzE7+PDjHm
bH79VhmoDZeQ+xXSXjeyHe8Ivq4NJuyGGg+5OkzHP6uyzAN5DjlNnfSBqVRq
kWtt4L6gwRDDwr6g5bLSKdwyiAkrdkcZK5aKVmHlf/+ZHALG0bTABDWNTSk5
9nxmjrTP7UEA2eddLRtjxJ5ZkIqzkca2KaZi3409CeNCrH0AjmvWmEqXPJNI
5nA6hv13HTF7Yz5R0b8tC20y4FpTBO7w7jY+etoExf6Bb1JvKmX+c8Rhubyk
Uw2H+cEdNOQ+NobrjCDl8tagxd9uYQbxY7MdiM3WESxTFZFoWFLQO0XPDa7m
tDnGC5wlCSQFWiaIhXJBMQJU/wxpuIThR0LUJxeRCtlhNcu0v+gU2voYzU/U
FeNWzuKGguAaPnfIuWwSTdzB84p/B54KysZw7W1V0w1HyO3TV7ZeyItdBUWU
jz8pZfaiuAjuMZ+tHbVEiJHeCsdpoqLmWlrnWq5KlOknaczazpd5c8gHON0q
zonSjZu8mkRlHXvx8LU4W0EFU7aKH2pJ9/Dpg3QeJJxwixZ9ypRbby9XsER7
SyzW159CnBfkd8ca8LsKQ0yumU17H3mZ4wwjwYOOZQV8Aj4tr7kXY2OExiUx
9hozYgUpNNDCcXmEqicPT4qb3dbkPHOPq83UtElbn+284+aGofUic8vhh2aI
CV2VdUNVSTHXEDNXc0yOsd5Mw/Y7jLL+8HyEmYca1IYVYdB8DhwmLjE0OmVr
vvE7dmEK3Dif+v97trejIGRkmJSNu8M2rBXpcMl+nr5RQQvx/ZXSGxFQ+3UF
5v8iFFePdOnjRWRcGSoEJ7Y0EA9Qk6xf1517xoTdzN4gk3cWUGOhnqbngjJl
Pad5qUxLrJAjOaisrtfX8a4dntbPeWS9lQIwFUpZLeWGAvlDF2vWzqTLpd9p
lpUuUHIAr3OzcHQJ3Q2hmjkB8AZ7SY6FkIoxCxAaGWduxK22qpUxSMNfAaAN
3Z6U/ImtXGHgVO/Ri8gb3JKKxQwaWuSjKmRT4NrtVLTRqgvzK5XD/8JG7sMS
+Y8USrcu7tWdgbsYIUm3BGqYgEFcxGKuvEN0ATwoKUQcMVsg9NgKBYtVCmSr
EJyzjh7OHx36VgSOlWy2yBE5iTVogC39P7h3QTKjwnymcEhXHjVOLE+fbWpA
XocPlCEWo0v4UEzyVw0cGyeNjtyt+wp2R6sGBJP84Za7HoBEOCM/KQDSdNGN
obxW47iRWx266LbDf6x9tpU+LFmAQh6wie5ryJBvRSZe/sB0JkRl/HiF3MPI
gyK/DdTmFDyd6xpQoR1Jj+NqqKfboN6LuUeMmzeL374ElctRDNLljilySjZD
hLhmAKQvGvcK16qFC7bjen5XRZy514tMgY00VSmFrz4k4xUPhzDafAZmwau4
jHWUgKDwm1jaxgPJrpjGCP6MPFOoZxg7FHslVFQT59dUpg4+vU8jLkNLPUYS
oWZ4qc+wMKbQJq2KuZL6pucSrTfkQTL58TLnuDuvFHWLVMAI8evoLvJl3IbL
sNchwpaR2F214OolN/Zk9Pbds9mnog6GDnwi6BPOWvo9hRdis9ZnYVk0JSC1
/2QUTS4kYGVBUR+gxO7kpOcJJY9GE9qDtHA28IRoajAg44jGt2oFifMAyxpW
MSsOVviUGWdqiRWzArpTThnpKwc4U2aaCQdos7qDHynJ+nJObd1EQh9oYvAg
O11cXobmspOA7UL7ucAHOianijJSfEWSn1J9UM0zwcd1c129lwuKFw2gH5M0
gJXZ+Wwsl+M5r7vN2GCcSgTWCHx+FFYb6UOLmNNMBGIkzfhqbk4dnQhiOAqR
2TzOy138/rKy9pMkfjS1TsmkBZqsrKO0+ny2iUc78+4zcOVZD6ygrJtcmUUn
ajRA8I6HpwWMbQ3ZBc7MulVlgquuLr4+pkRtKoDNBrcoUK0OBdEbk9SfZVQR
QK6fTvMp/cKd0ba8Ii6WFlhllk7iU1/ocLoOZBDzqlabIIfeikcmmTKstW1n
y9vTjhVUyoxHHm4IGnTxo9n2R+dzZzRklwzRZKj7HTRBAGSASOIRl9m7elBL
ErPCUYbBfsAHa6TY+ZyJikW1AhCJNgdX/EoVTXaEwwHVyPWkNF140Ob+A6kM
Mm3/67JQzMkUN0XXuoLxdGTrR2rT8ehouJ65k7yjBxZtQApZKIkPXKIC4dr5
42qVOepRbddkYbDfOTPaiRjSRECOZ9TFfEi2qc6m3wxS3qXZl1+RoEyHtANR
fjs/rVFH+l1Xn73Tkh+bESPqnYgmdHqrr7fkeesYqvni52krOqiwKjU0NDtF
c/DFkbu4WwYZUXpZUF0GyamdjFLmcaIUcqBQF4pvpYwzi8hrCuF2qX81DCHH
Pk65NteWoRQYN7gs/ClSQ7/uy4Nz1TXo56kVzuFky6HQjchlg6r2LrxOyXSF
epujaVGL/ESPCtyCwKIH4mK6V1FHcNQ2TUuvHIP8W7VOfrmgYb42yGd+4q7n
Yu0pW++b5PEX/rGxK9wSzAEGREuPTlHPXNRMPNK6IPQ0UriUZfqvF9QWI0dW
4v3sH9Y5MEiWH4/ujQ2GntfjqZrvU9Sjn8sZWf2wAaZpWUtTVHsANyyb8/ck
GoFteA77U16i3ux3HYRB+d+UB25/r/qV5p4SUpQOVwzmsorMFHxVBj6i47uw
b3eSPk9avviefkIXPdB4pc5XH9X8T4SV1Va7Al8kfMBSxR+9CIIy16YDHTMS
uaeTvEEvApkASpuutQTHu3hhGO2QI1kZKQ83qHICMt0yjh5SD8Ys7zIH5DUs
jUaWlJ/+nD9DVXzqrA92djudIfROpXv96ZOSPEIXWJM2MKX0O4nHDoi4++W8
gZxECXBjD4PRu1D09X6I53zNoMiPwPh27y/htYm1byUk5WEYAkO/n2q4BXZV
/1vgs6v1N2lHXZ6LaPO87+n3k6f+7JJX/4ikxBjchYpXXn87d4wYPe8f9xgB
oWimNtJla/Y54ZiWaA4DekskvzOj0+2S2aZP3Vy9Hr62mGubZuZqF1wpb1lu
0o1fM9GHiwXnQDUdi4z2W4MFN9jHrv8NymVesKvlzsL4rKNoxxCHxaOtwZ/N
lwq853g8N3745nd/y2rV11d8wecbhkzolrskBX4WI8/ec94ZETtAu9F055MS
60mQtN0DC2wUvx4ULqm4eRyqvUQCRpggriUliHQdY/Mjag++bXnqCYDWo5I+
DCzOV9CrYOUqrQbmB7Y8Ro7pD/86lt2/Kf9p/8juhLHHnN56jv3XnlbtHx4Z
g5eaPsXICtlWz5qwdvK1cPGT7OOB3AlwdefPiOlqj6mCLJW7k6iWNB2mF2r7
2Pbk0xahIruKnB2QusvEvD6xz7OkgHLZjJAKvHS6z2xPP07yYuKq4C+G+h2E
88Ibx+/CIeaATC35ESDxSDIZOxz5/HkrBblTgmzRYkradB4IxR7MsAksA/0E
nKEKurqKYFGoFM1nqbutSPNKovDLxHIVH0++sjJWCywGF3KrToDyV+3JkdLY
Uk6dDs1GeLEgSfGb5HOGctYBXeiSo/o1YcouFxmKKgQe2xTlxSnqq60k1m3Z
60LACCuE72OJsNWf/l7u79xm23UPiUjEFQ3/2lsUeRGsxukshjrFKgH6FjLS
2V6T77TGIvFqeWO1uBD4hO8FSx9BzM/Ja10bhdTBMCPFIaJjw5adcxznM9OM
Oq9TtvKiPK0pt8nKJRP4vcYVHEwTukpXKvZ+ft5M6w+1SEmnKxENA92BjeR9
+uphcrQo/QaIauVAWorBgmzCFZ1jFSoBvHz84Z0LAl3GrTzatTTimgNiRSwK
qe2vGu4fLxhXxTt/81X+gHHZPRa+7XU7ufZ1okWTEkGuS9Xhxm36XNRcCVbc
nK9jes1RS/xfijUTCL/2dV+OeKBQYe4Zpt67yEBiYZ1WaEfnhQyEvj+9bYqV
UQ0kPOYjDx5TNvW9HTPNgyxZCatJztvpBofKHxbhzzSJXcBJlh4QdwTeoA7L
1zya2j/h9jpHMN6Si1lNJLVcg7NevuYGOB3hkvHtFkf2yG7jwwFod7McOG0w
nK+zugN0HqJ6T8xDgPZmcpEN4s7UkLwexvmhXlc+trBa4hCYtHzdqELTkp2L
R7LOEDwYI+86OdQ0T0orPESoJdwNjf49dejg5XntytcZZ+jowQWL43H3T4Kc
foaMKU6+W//GlKAbKQMJleSAPoC7TTFac1LNozAou+SVA01s6u2pMS68tuyt
t1UJ8Wx403lIdfGlmREQoj1/YBOhUstaAy6gZqKX/7KcUKyamScmJN9+gbKg
iqTgXZca5j2WkIvzeOPIvbe3ZCim6nyJ6Y1vwYXRo/o7mWpHQju+FWOY++Ob
Nn/KQMqY0MVw0zrL/f/1ny7QVhC+aqpMDYYv6h6lh2ElqUZMMmnIvsApAFkv
of3PZkQ+N3Mr4ocfRnVh9cS/OqH0+lHFXuusu2O7zD+tN26VN0+GWdowBmAM
Bee3zQ1EyRV/YwHSjuWXaVI5jTNk4AQ3au/toL7UmjlKBxpsM+yVb0bO9PEt
K/i4LvyhZfMkd5NxwkY40C0OvlbbSXAgFfXxN6RuxQAQI/3/nPVTqqsaGsTu
i457uD2H2MSbRU1M+d99NAzmpOpc6KXQtO01W4ibAGYwDxjE9Ch4f8Y+eDVH
HCBM3V7PT8nPqGtyeUpPQt7ClgrX4WuNv+s0qo4H1lR75jvqy/Bw2DAgEL5E
fpDbOEZjTafhOo5j+PTDEKJLlKzIA9ILjkJnT8VlJma7g+AvICciwUnzR+Ev
q9P3QeFntaFIAaCqJwrWqZMQNKhCRZtoQF8me4OSGdyeqvyFxatGLuocVBEP
vRKKK0Ks1KDLGCWlc5Cdy2lpJkISakyf/6U5ll5yYz2YiCO+qrKHEzb7Tyeu
zqOEpJZ//OAlzU4fwQ99BnwpAkCus+FuRyx13rhDVPhMANUPHha7DKo/sgHZ
aaZMHHIFssEKrJurzPOP8Pqld1oJ06jUn/PSOIPTGjZ5pJM3Dvgj91b6rYto
Uxd/i3YwJqSaqnTzH53EcY/9ghvfZBi+evjboGx35hQnw/xPshF46DXles3N
viK2OdEgl+dQja0CKA4Lv5RE/joL2SoBFZIfE+vy8MPV6hsyssPDSvjQ5lWn
W8izX4EcDy5nOWqBei+NFvnF2Aut8YAjw/L0pE8/k5u9A+0ZeUgSzvC6wsTw
T4cYZ3rd1lLN1S+pZ3AJuZ1wui/88jhi8OOOlAl9UqF05NdA6iJzfRX5yHTP
yuqe4Wo8b2R1IMGxV3eyloz+Fa3Lac5LVZS6XfYe657WiU1AYss6hu4cKbyQ
pzA1O1seZIqZj9O1vQ9GmnW/RlgnNRy+rhlNW1DWXzXgoQpiqnI7F+r1gZ4K
R0sL2uVJjKIn4G1VUyuZwGX2xrgLM1ID6RdUuHpUHhF1ePvnUrpZ3lijYxRn
NvUEdeoIb7wBSn35jQgrDbhTkuEJg6dKYLQm+lNWDCSvF/f9kkg2gfhrFhTR
nuQ46nY1P5WXGxmy8SQids/cvT/bwp7QlwDlNH0WGLcy59JTnSCeL3wWicWg
NlgFaUfKN0i9xbVfEqB5tC+97TzIG4Mph6bUbWXEMfvT9UuWtN8MU6sdhHCi
nFjQQ5Jo2m5Wt2O1zN4HxdMGvGiN5vGNOYOzGe4d89UYv3C6S2tESoIHBtQC
S+ffgblzyRIkELD71BoUKycgMP92/12qjbNkm3fzfl5bP5E2EtKQHdyTP3nE
+CsKLp8AtCTnL4yWsBpqmZq+8scO2irmA/aBuyWnAcxisxq1qgJhGUouOhNE
k00cuAPXRdFtGxcvaGrl6cnliWGh0iv0G26cK0fozIwyL9ADJJJftjevmDLM
rpaGkafo0dEatW2AC7T3mSoks/PIW6Cd50qe+he5VYul/hoNbQk5/CP3YayB
sXL+WJR2sGpKGksNmtupvpK4LjCwd6Uvvm6j59yUHV8Q8Ih65paLsrH0VVkf
HR+ChE72NGrRWaqfTE1LxwcWZWKxbiQG49zyJYt79za6qAyFbezgJns4wv/8
bjE8PnVvaw3Xl3Z9cQ+xOYleJrnCvJDztLHKLjnFb1lBbGTRWTsI5LI4sSrv
po9Z/ZblBreXIhsMiE4ZAfCDGV9Mbmse4Vil1C+s0ZzUj1lBrk4cbGU+okoQ
LzKBIKsBzGKzDCK8oCJ5VuIO1vUE9pYPaCSWsu1HGl4TCkAuaV/5/5USX24B
tw50Zw40n3GZFFS+0RrTai9jnCr+3gWV9g9ENonl1FiZbV8uJqS6urOiNnCr
65XVDOE/8sFuvBzGVruJWWDNWaX3JiOqpFIoIsARP287mQXsji1dxcmkqqgA
PcZBKljBgnlMmynH5Be43dFpkTXzXLcann6gHuvpD70O9U+Sma6uGi/N7Ghf
c7FZ+pH+MKIynm1XBw/SO8JSy8xcNw+pFDNyFfQz+oGDH8B78ISckBCz6CTN
CXIfzc0hgR6o3gkiBqkudnWUd6KBEzgyhcj4es84d6524t0SYjTUiq/Y+kz9
VUQp6nAaJ61U+mRc4R2+dSvFlPOGCn/2olEZiqqSsY7Ez4gKkpPk5JApfn7Z
cpIYpZ5Ba9L/yjKG0Z8wKtRWUkAqzFedcLQM6TJVF3PNAD1iZpJRt2CqRZkS
pP8EhqoA+9oCZ2oNSkru6tlvjZ6WKKbX3+1rHl0IBzaW+aod8eaZOyMij/jQ
yYhwaNY7KjEMddZ2Hij9ESdf12mTNY+C4O9pxUx3hiA9W5jV521QenRb6cXm
HdxtyC1IV3541D4kY4jKTWmoG+sFxin+kRsXJOnU4gJvL3GJbY/nlQRLjHFH
IrQ2mESLW0NFEG5lcBE4n5PkAi6SQ7D8YWk7FVVvSduKD5mTW7++P91KIuCz
7MM6FjPIDp5h4I8CixRTJL8yocE9EMzkPM+Te/3HY3rpYlTZn29GZ4BjnsNI
BhKkL77mjbqHRvjzyF4Z/RoxtHWgsYRyOMsvQ1WOZyNyGnxkfJF7pY91G8eV
aATKYFnEym71aPBVpSKXDdsyTGwuHelv/MdWblR1voWB+JU8DkBTWJ4Bxs3f
e3iaMXDC+bpV6tcBmnOpLouQkAkl6jkaAXNHoNDzUzNa7XRdlJB3teUp/UG1
vnHD4LD1adCZ1OlFmW54tM6DknLJrCOYxd//8uHlxqh4J9TYvFYHm82VJQSr
w4NbDqj6JraPZwIWnnLI75iaYtHj8qw2gGi5kFhiGzGu0QVcSeeM7ZQh9kMp
S0aU5GXU2kfCBvpQeImMchiOPJWuN83V7CJoYZLto0KL5Xf1Rj1x805qEBO8
WS2PlcvW0NwPW1tkNeOChXp9fiv6hFs6SRnMwikXv5or28XlzbGIVYLwSihz
QMYAgUfRWAZ34xq5gWDq5Fy/JHfa4azoSYulEIGrFeBE+gfrEkW0oSAUcyDV
XQVM61sj1sjYB7s2ldgPrnPGKBSh81T1Yh6aUolKiob2raIWlCRO3t4jmW10
RuaUwkLVVz5xKB/MgKzUYEkRGzV9s2xWTq22+4ZTRdjGKOv8Kw/1oOiy3mL6
UUbKzewwcssjF/OKZLuD3Z2/y38HDnsPtxztpZmTdacKAFqsC6ABbyBm/1Lc
Xot9RbsR9IGGCQyOmkSB7+xVENfDz12FwTod03HPXKajQHhW/WhWFzBIq4Q4
M6zoJLTAAg2J7eDuG5TBmRgtE96uUEwd0OQwbH1QTvu+wGNVVqiwmzWoo6PK
7DhWXXBsWbra5rOhfRl+aP0+7oWurGZooH9JeWWgusmWpmsOYrOpm1naT3WE
3xYQ96OMf5HCpRcnFbwXknk5CxcVFDe+aRB5K6dl79BGZ+2hFwmZZMLTuht4
5zolEvbiYFYxvIc9E3a3u6g/S3lxTBWGojAL909NdCYLRn2n2iiJIrovAKgg
r9FCJSE8i3sqNl3xg6OAASUSz7TYjQDlJ61d4uCAipPSbeUCPu/J2l1phlEX
OMk2DSesjJFFjbyAg71SDemRYjhWI6HOXehnZl9lS/sLDjctGRs023HjCEmT
Ug+PYqg9YuKLb4dWKkgXrJPa+6qkzrfYaizBpgM7rQN98SeQu6RLgNIynoFl
y0L6hi/xjXXteERMQdzyeC0FjWpqUp6113ZYTfv/MQgZFV//ey2vUKyAIHAs
cIyp9Z8uXARLudcfreh0UV77hMeU/SI7p/VN9nc67p14Q49FlD4tK+7DrXcW
ETU+3UHg5vp7CatyWnOUQCunWBpYL5ZJe95zR5eZo7/k1ZmnZyHi7IUlLPGq
O+2BkWU1iSnGbrUAJtXkyut/WftRhqd84t5qbzQkb1A1vtMUTOmb4kpGGB8C
ubK7YO4ecle6MFnUG4C33lpDqqyQev9H7RNh5uQ//QbacmWcl9NUioBdgg1C
1jsVklmGe6QrR4OkAHzhIhISBTZy/WCkzcibOVxtpiN6XANoyOGISSYFGokT
dfUOxVCx54vzm4HViLl/EagI4udW3myvEg9k+pESTiKbSReSf81EjWckA28E
URhlMQx+fhkn1m9pmgPj0CKb2Qm8FW3p8oJVqG7h6CGHp4GOZHtBTxm4heYt
rON0nKoWZR3sj/K6pVAdvnrMh+m8qMqpLGGc4H9EUWpFQi/Y/rxsMg3V4G7L
vJc9l5hM1MUay5Uyw33NWTUZmQbxOgubEmQAPJ0M60A+lQz9FZ1hekGssa3G
ZmIX/HvHvWrzX9Gkgx/j0NZS2PGBQxSamxxF2WBEU36uZzXL8AzFmh2TjZIZ
Hdd7+X7GmWm3qFy16SQEIyAmeTim9ZicS4bwvpzpgRfyruBpo/5/LOCupoTo
mAEgzaJWIBqMggFT75zZCVaYbIfu9Usab21Ydv3yyiW0RLmakpBGq10X452R
eHKqvNU/Br3nNGXiVVWf5Iz48ql4HPvFZGUWxyxGPDpUipdfCn/D8S8HFuA6
eu2HSGUOnh2DRvz8EjlVKUzqxQW1/j/gNMs1SdbzJ6CJU3mN0VRHZfvy7V9W
/1VullGbryC7Em13qHzHN9eB4Nc1xaCmL99+ngubesrJv0vtnVYhGRAWW45D
YWodTOd+Lq5kBa23NV7BthB3zIQGCWdBZD/6SY2kKuryTwvfR8o7o/nwrb26
WX8DArfrD0B7Qg878dL3pLlDkivZIgQAlsEMTYpdTpt/lQ6dGNUdrN5jiklW
20ECoMzeGOZDeeEEr69NWu3hWjNvxCy0qVNFwyKDrFP1B+iNk/x70EiP+Ua4
abZjziJAyHO9TIuzzvSJRqueZeovGT578Yk0nTav3M69OJRRZ0+7Z2YOcl7k
a8ah/ghKrGFFil70R+StpnWttam9YaGg183KCSFdjMHH+fiTIvoBHrtFpgDT
Nn59rFsm98d4s1oLdW2hTuMJc2rCzvSF2URbwoYUBkKkE/hIAl4+6fywCtkU
oyDRNPgABQcUGsqDm6yb7qpBVJsMk8YsGhCs6Gs/h1C6LgZH+QO+GP/bxcr8
wBCFs10jx08qlW24erWSD52EOeexYNNzeqbGQy47UeRM74P2woY2yl9ypLpY
QBfLdcZaBloSxOqc9wMjhBf7LH8YjMOKiLwQ2xEG0AS/Da0IqeRu/c2tHcA1
YvcUFIiQUk3G6/OX17OxZ6EvgG2Frf7tMZr3CrdOpHUy3iM8R/EHSP4UtycF
6Y0doat5q5laNe0uiJoJ8xnYkS/CiegKYDOrMM2xxBOsiN83p8vi7/Z1ciZ2
8gYO4WQ0yStrzQSUfFJspEkJpkgmKmT+p58eL64k+ZZH6ucdHHaw/dHq4/nS
OYiLF04B1au+gqrZrlaFcxxtzxE2U+tehsKmIytpvEqIT+lxwlMqoiI1H6pX
yDaootorqiAZMusi6c14yn/e/SB6p/Twp5BLSuVTqecHTYG6kIS66Hd367ck
uy/9/wj1XxEF2oJB2IioDD/xf4n86d8xuVrq1Jq26vSB8n5iGvEH08YDPxpV
oIcVSPkDDfab+NFIYIyCooVFyVydgXBU028wxK1moJIrgNlzD0fl059dzJln
lBg7PQd7GBCdsK3fymiVRsRYKNk3LF6eWKvY+8xi7MpL1e0XkwFGrW+Er6IA
uy6ffIUX8cyJJMn7JI4lyvE8H7xiAk/f/SjjUyDwxJ487DJXRb/dAIGKlFk5
OgXeoFchTXsXIrU3edlX7NnTy4wf+3GyTnYTNTfmTwEyOu6v+sR0ejKs+guN
tvsZK5u0PZALSmJKf9kAyp4Ix0LEz64iKQF04eYkKLabi36H3rwmnE+UJ9fY
sGd8o9WW8Q0ct428US2TpNYed4c0CCu02mkzCSr8BleLgk90wjE/zy9NAzAs
Uiv0dAfiyn2TyAqTjc3eFNQCa/V5ALaUuMJ6MUMUnx7TKmehT+fiZmhVNYGD
ix5fR6b+zEH8qDQp8yAK9v4fdKmODmfaZ7k/JuG6ocqejpOKTz2MIaclAxor
vi++ofsu2BFfXWqOIE7hXzHRr4qRwSYUFGr1sopoHXJajfXoScxOYasmDXwL
ADglsd6D5KtHCWhgTOKV7wiXmaXeVlsVrQ4TG1V4g783RGPz7A5nnsadIOwi
ClvyLelk4287SnE6hOZfliKrpw3J+bCrG/IetAWINOSTkTgLFMNg8r1ZNzZL
1njFBXjLvqF47DmnyjO3ftu6mDw/9ta8Fq62Ce23AS+ulfXdReHg0BfwHnW8
ezMlTRQNn0AOQ3S0rfWV9DxNss/tTn4EV9LiuejNu9SFc6SnGXGx9u16Qmu5
tlB4zsJEZUe9/S7+nTgj2KALf7dZbDqHKmE5k8LUE8Mtgeu/2LGh44ldTZ4f
wa1RmOCNcR3X0iVleQ6pg/w+ENtDHKzVd7C+YzPCf10EuDp0ag/2fKG+7L9a
oIDDp4h2gyBl4Ftg6EcQu5/nwS3uVQU6v4ebUxLRiNpCOl8l8ifmYM8+N0d3
o/vLdKpPqKWzip5qcDIFM/4Uwto5Gd5tjdewz4Zql7xaRWdZxWen1fzdH162
Yhos/uxJXAUp9Bo8jIf90XmRMOkwJPTXxdoPYRlkhkuQTiw1jwnwWJu8u9NO
d3EcfshbaWC5abRITvJd0ljiJgSDVO8iEsRa49aLcYPbVQjVeb1odr0IyJ95
UtPuf7ScSX9AIh4XAhzjU29xlrYE2a9g7tbyTvC+pG0d/duUe2FpzC06Rfg0
psub5Lf54/W7WHnn3tr7KFw5Q8CjsTR1wInGujXXRpdpNdOxVsQwCGxndZM+
wXmD1UoKpnTrP6K0G1RS5lCxRkJf2SLpOFr0jh89Q5AnheuW4Gc/cE1NaIgX
rznRRfLEf6OG4MrAxLH9obL3j7UtU48z1e/uXb01e+zi/6yer78RB0g73gU6
TJlXL8ZXWYkgHq0jVPzdDGh4JKGqjMawICGcTc2tXGq585Dcz7vktkr8qdxJ
fMZbBiZqAHHALl/rNwR+K5zB0QBYhlfqd/IEx7P+pjvgZxSSf63z1naoysOk
/4U7iwwhchNcknZTHjZRDiWGkswSIoh6vTFaegtbu7pI5GXEEzGQjFwnQV/P
qkbw00fnJrLqigchYTZLMqmMv0Q1zUPEIChsy+tOW7BhcX5XrcThpCG2yqWa
5nNzcFF2YgBzN4bWWzca23PX/yZUxF5ZoTZdxy3yLIsKLF6+bGkOCQ3xdcJB
/Q0oODDw441hdCnzplEI2V+/XK8jveetYcKdI6kjS1uU3ebRtfyCBpTOYnua
zXmxbHwo+tq+vmIpNc3/69Ng8DcaBFScaN9+WHEyBs9+QLqIGS/mgQXzJVFC
K5mKrCq9+P0ygmoBQltc4eCF38XVPuIH4RoP+kRzmOO6k+aoXpuCUciFwLqc
3YAM7Ga2sGcd1OQjQWmCER2lqiPFDqzDqMlPVkZGh6KYaZFg/g0KFGm6aQ+q
zIwgkGpY4I3xeclYV6U06e3Logh3xj8qsB19+AOpQjQznTVj3o/ILlPQ7d6B
l8Vf71fE5HU7ljEV9yIZ1i5SlDpBrnSbu3Dwg/I6gTqYmxsAchXSIAPvEJNX
zeO9pd9BF3j/qv4u+sKVwY3oEgCEcZRiN2aas9piFKrl8t55rIAWSXMgLDfI
GdOz9hmWlSN+AuzwSkOWc7auaNMUayH78JLkraAoRrkSrsH3NBOknUxh0Slg
dV9FYmmzN52oZAd/aSsQjw/2ijx7iWRaYwHeWEfsWa180x+a5ZvD75dX/RUl
L6Y1fWTyY5NfiS7rLdVVRh9xMSJnY8N9TcUJH75wx6tspkyw12XKwEVEjKYR
ytckFRrBgYevm2u7XDoShJYW8yqAjhajYOGkecULEGQw7TW3JYF+piN538/S
n0Er232fPTczFrmBdIs5OtWJxoePNZG+X2nvFgx8W+AoAMaoBzO9z83uxGhR
BRrA33i36XmtArkjEgiJ37N6/olwNN6+2LQgn3txcanU6ire43COMne48SC6
AIi+Ee7iRn5VWhlbjNhNk2qerdjpxuPjBmNIilVSAfBRDDQ1J8J25k2FEaLL
drgaxlitUTxjFmKGZY4K0Za6+3DJOUN/A8hnmZDSENINiqlAAFIW2k1uEQ8W
yMyYFlRjRSiURwfYS4sFYI0R67q9Xqywos4XzqiGIgDLl7QEEYuOIF0RVXrX
q2aFR6q3Ghv/1qW6bpKMaZSuBVgc0Xrg/COFjb0QU5kHSHlbgbOgLBzGjE6Q
bTqSNSEwwvc2AmVgxu5TcCP4JyqXVs8SWRTqUlTlTgOusOOZbBKl9wx/AIc7
e/8lLTsrmIrVy8NJMaJOW7NW/0gDOrlafiMU7NQQmNbVkTUTesOpLILbrEgH
D63EpJ20xNin4WUtqcd1/BrMNO55oP+gMG3PvSOfW6d8S92O5EhJlaOJnlDi
GyTFgS+Vr8FDg2PBH13GnMBiLm6uEnm9ZbQdYe34Nk9tX5zmVIiOkdg7BnaM
cqggkEF4lMS51WGEwNlM5zt6uMklPgIMD3CiOaowSiUOX2+57lpmn5qoSZTU
AE1xL2k3Hw1RHyEznOAiBT300Jp7r5wYiYh+3tSCH5147lH/GiPcGwBlTn64
ksd7Tlv2lCU2lpNJ8j/Gld47QsXHmIvNbOe8O+O2Lg9+SlDDb7BIrV36Z1Uq
NnSiI+tLzq24lc69ZK6wW8k8jJMjonOK3xP5lNZxvH2SW/TXc76LKFUeaQ0u
DwyP5Y8ATTJOml62JQNJpaqzLPh/92QFw14K3qRzTm9ykMmxN0Avs5jy5ZZn
yupRo+3nqg0BQOfcloM6Lp0Uc78lGKy4UtAsrbk21sRHdjXgEVLdvmk2gGui
ftbhU2Epr/yuQ+nprm2fW43cdS+YoauzTY7jSdZOKXg7uuxQ6LJbHVVxPocy
5UftlWYtGRFoVK5cfMrd3glNeZY5QhCyjusSQ2GIwTgBOPCmD+RIzm9w2kTx
rKFMMwPa4mqTVZJmJfdtgNx9Fb9snnOMSzdyEHzFnYC0Vv+s2mYaNN+E67LP
5HbRIvY3vukypCYP1XWThicikxFqsWAf/EkcrmcOme9VCSPMJ1akDzrBqSSv
uNmtsfg9BZ8dijNYsC72gZQKqAFZER/+1sNmSwZuGjgy/5lIgn1FhPXhoQcw
fia7/ExwHA2P/QA88CLYM9D9AQfmBVOfjCDQbJxW683WKt9nP3/l0WhBy1oz
TJRvjff5GsFKmC0/a+QMm0pVCjgLr27thv8cmOAQ57vcbvcD21sJqbskCycO
s8DBLeKIv5wlgI44jS+uVXVzUdNVLgBG+mPzVuGPP3Ih5sqIKbqt2uT9PuOC
EQvEwcuvD0eF6QhnL0p1jTPxkcV8gx8f7/uFyrFwtMNEdDQuG2nt8cxUlpOW
9EjvczyNsUABmBs4DsmugwoIL+ppt0kiy2/XTuO5jatJw/84kQ2l5Nf/wnhN
kVVhvOl0blVJFNGqFZrdCuZFtIh5RXr3Auv2+liM9ixtgyaR8lSVdTjVuW7n
6Asp0tzIQTskl9IoPHKJW7p5nzmwIJBGiNdlTx8NXf75cfpZ0/ffQzHIaSKQ
QHDdqAT9j8U3Zc31ZpiMW0OvRu2xFohzMGwHbF647hIckwtSRggmrWQ6YzX6
z4BFlGiNY+7PxhTF7vqkO21N1hL8nAmTqZTzM1lnIgOuc2M6hbONKO0/73YS
7IZfbl3pEqzzt79WgU9rUPZdsdlAIKKQ73tNv2s1mRZeIrA725Vu6jrNUl+R
uJ0+73gQfJoVT/q6VP64TRm5YY+Rc6Pj/MEZ5SzE5D5ZtoSj8rOXoweEpWyo
GnChaJ6tDX4QQ6jeHV1jREpoOpE4QM9xDaXEp2T0gs/G4ckvDhrf/DfoqAMn
4HWYy2+THSM2Po4SUA/ZhQaX2avSvjqXYSDYObyXOPU/hLjlJv4wWVlFzABi
bKfBtc9XdQtPIGqp3+xwBr0dgkku0+HnxO82CTPhFNVkmcLJLboCheikp6zy
xTzj3/9gkGuWUwXQ3gQwI+i9T7W5EsQriPGXKetxbVogZkvrm8fqzNzWH1g/
CkiTcdNvEswmCrlW+SZHP9ZewsQdISwU0t1xFciyzuiyYkEJx7XniViw1205
uL96e8ol5iUtnVH9Q9cm7h1VJupsy9H9bGsr9sDDm1IeLcDOh8hkgGj8zpPt
ffUAQ5oFqGoIo4MQBvNjD4ta7yzYy/wdRUgwFx5V9P8VBl0wAExP8XSDGBNw
jtcATU1imltC8ky4a8dytmypNeWmPNYxTSjr1CBirIt+ZvEJkpbvX2kG+InP
gP6mgqvv/Q3wgcBrs53SK/AidHQ3MkmMNv8e8Lo+Jl3Z04KHySdfVia2Y87M
KeP0JDbbX6l8vpAfathxjQMM4yQFR87XHSoiTWOhuD1pWKIe/udsNrNoUzin
DXg2VRHjkSYZHXsbmsLCik0RIHFsMFaHbLgrJMzAe5o7MpUUEZqWL4EUo0bl
DX09QSvZYGtt5rJEURlK3DaoKj4S03cKpCGkCXcLoI0f9VZM5Gh14y9xUrlQ
Aix7BOQ+Y/mdBjRFPYll1p9ZCq2pD6gmJMWAeUO3gmY3Eu49DrD8XaoRS4mg
n02TZN6r1XKY8knoPbsf68RCxqT00rGy1X9O9M0AnLqZDPyrym1GRWC7IJkK
8ltUxDIcozAf5VpaNfDI0ipkNF1Bn3WgFF9uk7BR+eJbo/qg9yZuJQpCsFlR
1oCRs7klqjHm1BP9PV6JeRFTLia2mvotv8HUC3IObUwwE0bpZ8giqxcgI4Q/
KG4zZYywvrxBqbifkYXhkni7p9iUqP5wvfT3luIHowv+cEYmRHga8pzKv9d8
Tf2TmmGORUn/9+neYeLShQViGv3lNgem7epQoXq2MrGWvZIaRlA1aNqNBaBr
NQIOnUGlTZK2tb86bSe+no9dIsGKdMoUTjBSJKxVD4oTfsCUewpy4Mh03bZo
dOjp5WQFjAhl83MPDU6n0QPZirX/eV7U5/mH4nxboktTenNGl5BnZOh+ORVD
0n1DBih+y2l2o0xfAoCNdzhEgXozxJMmoKbfMkjOjXSVIq84+lo8CF7JC8n3
inThGfIYY89XNv08rK/cf2T9YDutoVDcV/1OhkvpVNPDwshStR23+6ct+h/+
y2PfIVKbm+D9rIew28Mddz+TSWP1QOELwTCB3hc7Ex1+Ebz61IxWgi0ScHTs
XxfcvEgkq8p+ZvSpKutFRMWXf6BigNRKE63EQyE4kM+hjSSYgbMuSsVe2MKj
5Is4r8xAGBx0yiiDZVQWLQ6CuvLtOpEVPxefYCF1s0bzUNXuJJ4tMi75ZWJC
4vx6+tA0qbBCgrdX3EWTS4Kp+HtGMa/4Bcoh0ZbJr05oOMcJsqsxmdvSk1zx
oBIRv1ART7GakgSxCpW4t0aZqMVqPAhnz6oiMqLiGLco3UHZUjQqoUWB4eoR
lFmoUFarNOmB+gM3HCGz+YRYm0S+y/Kvz+BoUE0TKWnNramzzzBjsyq/Nxj3
xnQF/oVvfM+t52y3Uflojvws7s6gdfOF2cLQlDa/XDaity4ycUrl99mJ48Pw
pViCpJjv9SgRLK68/GkqzfKAifYVCH/2YQszQrZv+XFmALRT4nnVH8TEVijj
rm8DVr/aP6GlyuAsdgeKa74otrVuD1h/KRX+ruTFoVo+uGV1ekjj8oI9Fvx1
2q7Qe3WoO/TQD9Mdiirx2h911e9UfbZS4UEzneZ8Y3PRbVsDxXW6ihIpUFJ/
yLmtfCfM/8Q7YBRe9tONC7r7YiK1tsKGLmyroZfJihDhyhJYpbnwuiKQH02j
lWHFkWZ9PTom1lL8Iut00H3nHw0uywkKfPsLZTyUhM8ZTiA1VJ0uURf08ZkK
XbXYx3kL5KmO8944E4I2d5x5dZBeNipeHltqwCOgwpH0i1F58KgZyHEcqbLa
FEBkTCGw1OnPbJUU8Mt7gweWNlf0PqNMI8JGEyR1URXz4hDwQHqRdelXn7hZ
OsNUvVmtGEgHujuRAVf/k3aTdQtT2oWo0Sgz6YGYbCaUKZ6Qz0DR3sgoPvUJ
anw2IPgBdAM8sKqbHzJW9pQtXcuN0/10QExDmx/Ts5HWnwin3ax5YuCLI3t5
gkagSwNIUh0GsiJna1GIn8xWAflU+/idjzzTUf2yN28mfiVk1RNPpeBaM8kt
YLVk3SshLOreeoiQl/pQAvRSkoPZqtawa6YBUAaRbijcVAUAtTNCb+/c6cLU
FExS0Sixe+rGFH+6KvCXGkKoG/kazAz6p+yBZGUd+m4JYRLHlesX5EUnlUZY
cslyfL0QL2H7DtVDAflcsDjMM6fbzuGm3lQc9KXutVkpOq+lH/f+09dRvq+i
2FdtecnMllI3Dj3YYWcAyILH8/dwYCK9JS9xLCVK1KkXP75xtieSlBq0KTKf
FZi4AgacfovATh8FCMbk+BkgO99C1JmC2v4LoohOzL8bKuOxFPRJwOKm3Ohl
PGzjHIGpOc2UmvTXL86qUrcopgTM85Ez8PuOM2jcB7h4gEBPa/XFq36Q/ctA
nW5C0U1uRwgf0krdk9qQor6vNx4wC53853Bmi3GJx6mckpzf/bxvyyZ1+ciZ
v+kNvBoG05ThqfSG8ZGcYB0auQyBfDHUGIWK5p55R4hHEeIGc5CDaJmhdS2X
WkcoQJfY+36xJYKsFPYcBKq4gmolh+/pD8FVSksKBIiund3wYQ/KZHhw9bKA
rSJOiqyW80dK6bvAiFixUlEa3zIpHByUM2xi51KayrPLdO2zMiYSyuT/eZrl
mt6fjYyT3dSIBuYtVUXjwKsYQm8mcFRYaJuS83oEWwXCOUbB7hkrAGJt+2cl
2EWyr8QWEvN1CL+kFxcBBnQqy6mrkkbgtvQ4IgW1NBL9m/Qu+W298qNcxzce
ET/+NEJg70EUD/I134Eg7lbrcS9sx+SVzIrHWDPC8dPFllzG8RUDD875KZ5e
o8k0UiklklPrkMUisiKvgc3RAg39pPDGJ87DnPJzG2+TDklAh3Qlj70m9XYq
L0HJNcgq3DkJQ5Du7URpD1IJ6o6LbarCD2Rnmd9GslSwKP5JMwm6BYaZzWnK
8OrlGSz3Wk7UY56FYGYeWRQNve2FjBP456Kzl96Bvd4wFPEs7d8HS8meMsxI
oTqUmblxwXlHC24SCk16J2Q5iJA/uIVRBoWWxIUyvGFMzKAW390yYQtzMpu0
x1yH++toylwP3bTYi5iTKRgPDp868oY7ovI/GonlzdG9J503aFHcNO2Dhmfb
/yqT/yf7Hs8aKElhI3U9jIvjV8dCCf6fktoKZMK0dBgBz1iPHGWv+7rmnNS2
J+TRU4zpL06/0mk41h3Vvgowp4TJlrQepWn+v7WozWcRuPWnbglvhTqjo5yb
A/yQPPboyziHcgxrFRd3f4477oVzckDxbxmFzOTqEX+Br7ORy6YNCcLvHVz/
dGFdGe4Ow5/Fb9Nk7NY69xX32dZrrJs0CxRyNkaCnB75f0dziUk7PZJztb+v
p62B/UdXvcXPqNfDIUWsfD0B/SGJXV/xHmyFvw9GZCEu5yGWIYK6CvwZI2yf
4xrSl1vRSzAgcDuWz3SSpOwcYr+tNkjgWY51o/To2S2p6KxgpruQU0iL+KrH
f7JWiKjoBsIPBhDoZXrCaTwauJlB4YKb5mKppGHVKWlhH/gOQF5+zLEwcVYV
GNRWaryzShy792WiY+Dn6jEoyYl+nsBjjVQ+ddv+JCX8v1Rt5AU8phj74MEv
FCzcu/KHgb4DnpYkbWkysU02FfLAF36UGh/EfaqBgZT10ajvihrjCRhFQ8vO
u3qj0/coQzIN1/SiLMKju7zmdx8eOYbfNRIRBhudfsVMr++94tscO94mzAP3
krrIl9QoPLPzeg+5gJq2GA0mF19xouVhfuO0Mh30y0WGzFpWHfksd6Mj0/jk
bKa6THT3O8yz2PLezVR6QBHQlzLWbFqSDe7r/5g5Jw2zsbSN1MhmRWlpC9ql
rnLSK755WXmN24TfSnLWVP9FSciEb4IDHUkWKm/ZyY5aCr1A4tbnah0dWxsB
It9VlAP90EyHbgOkDngA+paQBTecBHYyIdVvdG52y+BJ3Gyes4+JxTNyYS5R
W2keqEU+I77/nDpRp7vPrx1iadZWHKlodTOAT2Oi5LLZ3SFcAw6NfKg9E1WY
8vulPEWH7ajt+Y4KqbZWRebumdc5+DQ0HUy2jNXqst+OUKzfM4KQwiTRgwfF
9wPoYt5c+1jMTVALx3UgYKb/brUzQR84jo5mU9GpBiQlc4bDHGE8toLGVLFv
AeZy5987A9vll4Hmh5dtfbKIj2BP4J9d+QS9l5W/TRock+Sa/cEbNlkfbeBx
x0rK79MSVWkloTKmljCJZgZsa9WYsbZhP2LfDgWYg56LKqbWIRg7965EQRiO
E1xqhPzdP3VF6BorwTY1Cvl/sPGVSyOuSrbb7iLbZgyofmaklT7jilidAc+u
6jz2o5KtfHiB2lVG10hNYogYwe6HLSabOo5012U+OsJbCLIy6ZyVSm0Ha7cE
0s/6acNbv9oKbyAbklf6VNPwXll7s0ZKHejcR2g2F2TLsQKvrbr0gJQUmEXn
aTOXC4KIjhTodVssPGDrJC4SojrXOJnjFCzyKDU5MYan0H1lEaKT/h5djLT1
ylIR1Y6px1Fk58Qzq6rrfkn4t/BLeMiI7T0KGetWDHoPbb4q7ow8QDvPf2sJ
huHmHIz1P5ZNQcWdahgOawvOVn3VnInuBexMKcIq74UMBhnYcaEskcskX8KE
PG7xLbyxj21wfP6NDonEBl27DgMmUYDJCdR/jvxkKY53ErxCKSYQL9tuNtsF
Bpffis/kOLq5kpruZcaU2KwVuSdjJ6qQAWKS1UPOk0a1bAWOrt0hBAun+8Gv
IbBB8g8DRl9eQP5ggi/8Q0itUzyGZj19CzolgS2/NtJJZ/r9tl7An9zRb3wN
FEXvNiu08uFRkiafSR+a/3M0SoR72Pj5VN2B38L5ulS0ybbSqUOTkC6GtCBm
RGnt8+1oidZGkewPgiKGe8jy5UlbLqKNe8g4AzrjvpC3aNTWjMzxCm7BI6sF
beLyH+BXELPZ7FvrogZkQsjYGkvtuP4aqEIaWIr6GedMpe9QgXE+hkNmB1Ui
7oR8GF/86qagXvyzLgwdRcaCA333yPmxeJkQV8gIQpECI5J/Q2KBnaQM7Vls
4XMLxTuP5Z8gZCVbX26nOGHIDIe0A9r2moGiM9doT53iA5HQaZEKCitNrndk
SHMAHRUxWQb4A/Bo5P0/aP5u0xBUumIt4zQ5kIcdeBiRR2Ae4nqQz5AYz+fL
JEARDJxtr1kOrmRx3Y1MZfsUfSuqvrC6WpVc4MdajDLFgUYjOWdRONlcChvw
nM0zE+KZSIYAjzdyW5Df7HOT1g+iSnVmVWvkCO0eppCidfmFhH2CwqTa/plF
Bhsaeamn8qF5ZqkGIX4kjR8DheXlKcZ3yFQZucOn3AYEmmcotm9ItUNfU9D/
bl5UAZiXbUqZP4XVvmQCk4keW7gvZqoCK3RklNHlZbI+46YTLKuvVdC/bEO3
YoJRHuZi4pQl2tYQuscAzh47zMfEP1kSC+56V8DwmAxlVRq1uxfrA61b/g16
KtfTbtpZTEjHwIJLj2q52j1UaecNL7Rs+MvE7gD0gpKYOZtlWKmOThcCp7nx
YjuB5lQVkfTwvJ2EvDgjjfztQVt1mmDd7T9VmXW5ggsC9Slf09dgx8cK5j5d
fZWglA3QZBhUpJ4z0vLBu7xVi/04/x/ycuNjUL8zkBq1om/2L/7iyn0LnDlk
pYixv4EjlbF5QIAw/wcGXJbMP3G4qiPSoT2KPNWjVkUwRkWfRyUZTeV1zVl0
yTyZxw7bhCpkNg0bzFjyrkim2mAepnecNpg1Tl+PiVyhmBO/hMN688s1/Ltw
6CF2hq+D3sGNMip9GC155osLHJFrhqQbagBT4927r75wKskv/U/oHGfl8dkO
zbKH1EgGkpLheShB6/2vqJhMds1kG8UKdmc1JrdFaFKzKWe/YxW4A1sQ720k
BAwVNugmafOAsQPivS3GL+oky5/kprr/8fSlPkQwcDuvyC09+dHhisK3Z8XC
2DAok9g7WfPqKo1mGD4ZYP8X+megtGD4XMsEBBg1u6rOr61uWH4a71jRGPtO
p0/Ny+p6CcJ9iW9ckeEx40x/o6556F7A2LJU/nZObtL7Z80dhMIO4WxgQqB4
t9hZuOptYyRqKxwr74R3v6gGWcbgyxrXY+wUksAauSCcF9pT06R/O2yrhzJ1
XnTviTR0PIy0AdX6P62gqXUhpP/9xX9ofmpulS0Vjkl1UozDUS1ixb4cwPm1
wYWapv/GOzXQLY8KxwgC72r6ZW0T7LsLPV7fEtlqENwkQ4GFArF8NkhEjnhL
mab4SFZetTKIjaeOZgIgi4qqTs/2148/igZUGBvTa5qxJwSAHhSFCior1s7K
QdL2Jm0yWZRtKPHcNx1S8/q/PGax4J44Bc94IJoI3drbJBi9MSdno3T+Y5Zk
Di4vb1uJ0sC69imre0sTzuCz1QRvg0JD6h0J4SFqWzYFoGTBSswVNTw27xWa
t+5ktYMhEeZtobzZMaNFUCLukIVgNYi4wAb2kjj5omOhgnTRESUphyYkjoiP
sBFLmnc12AnA3T2kxDdlaupyOXPyFXmw9YIrki+gME1QgMAYV8t+AmvAB5VW
Cf0iquVmZ+m32/mIIWHcAL0XPxdXYfb3OIj+zjgsnd/OcuBVpIMCNPaFds80
9MR70OAcQMYaNctSrZjnS89KsAUpikrV/J7yXvUtfDRLXxzRovRKQDMEc3zy
Ytbj0lNe0YfFWDHh4pUW6Rc0WTvY4vgWOoNg9doISSRqwQd4CYCxSJtA+XaP
6mbezH5QkxS9PZw2cbnf/uNVB/pnV/j/U4g7cvzSuBUcLrp5bILXE+xlHMtd
7v2lEvslZPTHogaDEiYFjx3IDmRA8Rll/2dRIfLyeYRfmJVGocB+s0DNE63n
s5T9uFd0+IN9EIUhPzRPcYZ3lKiRVR1vJMVuUSi3LWHqblAK1XN+de/ic8lK
4+rzMCW91Sk4PZGVSgkFdJOhgQthVuGteZl0legaGdSd3EsoNBEXTUmyPtYB
FI6a+AdBY3iiXUby2CIRyIw2ehhDFSJtTLXwgUcQjhCN9BtjhHWxUwPYU+/0
p4hlBy2hwa17REyD/RUBY+3R92xCafz95IyiQCa82N2hPCHAaxqJ1yHu7HKo
U9QJQHA24oOpW6YJ89NNwPIJHdasb14XAcmvAGMgs+nC5OpeDYCqG2rROrkO
XnOBmKA8aqKu6MK/EMtx/Y0DGDa5sQTgJm4+2nmHRsqjBmjoSQ8ZsqeXDnqy
2raAj9ggClMh2O49JyTwJy6ZKxTn//Gud3BQPBWavOdkn5DYu5rRxkI4GIaN
hOqtD79qAwD0Vwh6g3eNysUMZm20FSp14aYMjuoXs0tK2pIAbojMYGR8jDyZ
8Qz9xqUgZsQmPWCMgOR4KC1RXXwTtbIL5gxEUg3w5IZX3Fl51bXtLTK9k4cG
V21F3ofIebKkAElIc4O3QmnTqb3aNQ9WIW7RAipNImD2ezjkmA2SPzMu8DKF
7bT9lcSmPx+oHck6jQ2TW+a63vLTSJIqtR+v+HkWoQgiaB2A4UYP4Ku9Vewd
hrs4umDmjGhjA8AScnh5p1nmdyp1nUTR3O7i/e2fwND0BZzi9R71S8E6Fqcg
8bRTre9lFkMAz/hxeioJDvhV7RzlHAx2LXdyBVfJg0oT04JX/t8qItVkmqrG
mjeqeorX1o68BQT4x8dfJjKU9ku6/kOipjCRdoHe0IyQyDAF4p7+Sa5/di97
CeugjBXi10LJwrkWcTnOR3hoembVFf7u++So04jFPIOzFrjPHLh/GoBKNb79
zEPL/PqbPdI14X7qoYgeuT587TJIFX855KXir2bP4rggvAPxC2l7bvNjT9+2
5Md6sI/7pwQnGIjV6v9eKC7nP5Z8FMowsepUGdd7WdbEWjOiYTrcoD6Ja6Hx
2HrFgWVT0RHvqgFSDEPI/jO4ZWJGVIwhg0V+4kbUwqtsUt+zLhElB+0HOdEK
aC0sGl0rAHypkAZlIq+tQGOKt663hM8GjXpenJ79D3RcNlmSVRqtCgFXGPPw
F/GDAlXZD7yEDSpRj/ggzt/2s2fYborTXWpoz7lmLc6JLWFAzg1amYlCT7gE
6ijDtA55Q9gbeC1ISoW50Vs1qRUtOwPMONrCOLSFp+rrCjEk8Nme+s25JTKE
3houU2BqONz50+l1FezI4+Q67TQWxGbUejqBeptfI+Ya03zf8pug0w0ItyeJ
swOUFVxlwgtEJznqcHZe7ea08x6hBJ7kzCCi+O2pkXZSfmBzADrd08nepAGW
6g3eQdRTsv/ZQHwvfYPXNH8479hfhmNqegr5Hu1e3LgVj5KwIhTfgV8zP0h9
RGDjOvygRdnQLq8exa/yNM5Gxe9iZt5bpZfwUt/okKwmLFnLroBuQauelrmt
+wyP9crtNwAc+nbD91dVpVG7ji1iYq2igTtEBeKJN684Nx1MhPhjKZ5KhTwi
EardOZWV1odo8OEG7dSQn2e/wCp4UVQPCCQxvK0jAo9zpww1kKp3xFYjZMyd
6OdGk1OkhQ77HS60kTYqb3EradcA3fqt67yK1Rx1PFf+f10QdYrhMa6ivcXe
8S9nr5MP/pXaSD4gZg74IJLH0KPr8/+FOqnI3pYBvz5+QiCmTnRAZaHHq51z
t0WdL/TRYS8hOBbn4/CClY4pq4JUGOY3CmVS6M+C2oBXBFf2hkzBCVeFAtVl
E7scHpRx9If7kcIqKJDR6mOgF4O02qBHed80cpSYOMydC2UfnQHNUL5AyWlK
WDujKqOfEHElK4zyBW0z7ue6v8fWhPBl8xyGy/xzmxPL3RwbnYF6P9jjnKW7
oRIyc0T1XNdbd+FZoNpnltmUR1lgHUQmGACdWDb1ODOuUUNvo/ffzGOGdHEG
7MibF90LrZgv7VQgdED4UlDoZKmH/u/8Qb3pfdE2s/vSdQM8Cy2qXfj06Tp7
wRPAC7cPpSu4Y25bDlZbe7ntutGpk8WNZIP/cF3N9DjtRFISIkljO1KjW4LD
R50DDjT800sDTLmwdCZtdnst6oj1BHLhO2cIHIoRd5/WQ6F1/nVKP+/qcKCE
rx14sBCTqkK77K/NNDflZS2j7bMLgPGOZp1RYUHM2p2yxFIUX30RuauhprC5
KaWS+sDjteg+5gPGObewYHUDRDACbHsDnIGldoAAS4LXXr25AfEPZyYzFZe0
lhl4Q4KBEHhmU4gqwZZl+9izLzPpKm5KGfWaei/gyPq4IQj/6wyS0C7fMGKj
0+gafZ99F3fM6PyCTCh7oU3AtYvXW2VaP8GtEYfXpRC8WZt6L9A7wwfYnANZ
B9QYTSTDh8YidLhl2qFOEZbNuH83sRUF4BQJzCQgdqshe0L1RkbfRIbwyKFt
UpFzmgjsUX1ijE7vqGqZTOnpHxsIvY0Eoxv/vioERLfZxvZonBvq2c4+d8mA
zUPQyn2ye/BQYzsjA3aV7M8aSfrjMbxgakr5xzJw9KCnerV809b/tUf7JCc0
BsczCEahOLexukb0qEflftG7sQxQvo5W0zGnsvbGO1o3lIS1dvrK4GKqok8m
zeQrbUMQRi4XtpGdL2KSszcOZLlykn7kmqJMX0e1oHDFaSJxBae8I5Nxzt/d
0WRnLJ7/Gl8XacLda/TrBcgL+Xp2jkll5Ov1MZctO4fsWSKyiDd+nru+p8jL
kJiFfhFK73KitlV3zoTotwkne0bl4sJ5t7pLdXpSIzcCS4WV/uHf0kCYxG4g
3q3qnBn7hPN/iqAcwQ96bbv/HTKdrA7nPSZJiqtwm54AmAz0JUokGHtVhWnr
IR5HtfC6zd6m1BacxWM9q2OI6uhaY9cKL8NfvnCSmKGS65YBEKjRzDTMF7xb
uAEWtPjoD6aug1TewN3NcTwPhEpjoxHEBRr0bUffA8ne1vvwtE36ITK+7gri
G8/2ambeUU2zKFJP2F9I0P5SqkvT+WF37c/J28Q2xmLphN6HBMKuAQ6p5Aj5
qKerNrdZXEFGuYI/FMSujdpLvrXOG1Dzd9msSdYsfekZoBTPisBSSynxerr3
22Co2wXvFgIyHy9P50T1LptgrarOBMNt5zR1IT0IkWev8a6IFkE3y2YH62Sv
N6H88kL/yPSWceCDzcsO2ZKfau7GcPmUQQy6a2VTW9oUxrzGconO05Hb55Ff
8Ats/4jd3qY8ptzbC8FjpEu9oxwLR3PZsmrHUH68UED//iV38RT1gXizPTLW
2me/f8DlFkgLvy1spZkTiQz2fJC6sDptqAw/3ujsRqgxm+VIdxs8z9kKfQEn
tN0Ffac+atRoi7cVXffVVYQr0IVMkj0aruozTqbXVjXA0kBXatshufhPHLTB
/Xa6q6JybTcEyfXL/oGCsO9uQOEcC28HbxzKy1jYeYHuN2CYU1AT+veSth3o
m+aQXV9eKTkxIfsYjjMmvd5aGe/h68MmNxH4eF6cS4DG9Q0GdgM6okvMoK5A
dC8RDIEerllYwL9bUBNGjLtEpnofjGzdGCHjy/mITGwuS/4rxZpzQwVpGFBW
mrlcqj2BOAMpn7C8j4t+/6eW4NAqnFX91mJNhO85EuCBVBMAWnFjRDs94Or8
etlK9flhB4IuMUDE5Ji09xK5fTUjzaEB5W4x5r4LDBJG/s3IOms4QOvufz4u
lsHsdO5RCzTylXw8ctRqUb2fH31KstsCl1OqN7Os0z0TgMH8qF4e7zQ+wLVs
jS81rnpQaYgOqnPv7Iq2EZxbabp7xhJRPrIX7oesSBJgDC33dVkNyaBNxVOn
6bfbb3H5mbhH+Fpymf/MQrH/E5tgPMxWnfCt8DYzYCeC1QcmWd+4X4Yq0aHF
LH1Akp02D0IRPqQIiXNj4LRZtP60yLLbNqN5yI3h9INOPLwWmaY17K0JYEbs
HEpedhMEsQWVGrowWnMGD4vvTNQye1MhDBak+g8u46WbD7c6WWnrrd4Hx1bV
DhFp6v4a64nmOq/ZBQeTOuEfjRbVpW0MtbFiUHMdYtGSYpWt+vTvp79LPsF+
XMq1kez6FcF8Sv2cAav902iUW5HRQPsGqJS3m/Kso1yUUt5eH4pdswvtjl7j
u4YjMcp3sGGN4Nc9A+jD7zYtkstbsRwRgStFCdsJJjXqbHLOBagKzls4cvJF
VC296hV4SgwWgeRvzXWdbldCt3QwOF4BFVrsFcHj8uiRqfUkhoGHwaL8+r5Q
wP1LDZP3RpgNj5Imt8gql3mIIpWr9gh8gGSfH3sxeAMeGgVgn3kRlqEHMiI1
bSBbkuOlVskaxagl5eTTMTkQ/Q+d3iVSamCplIE5JdV6sE82M+j0WJpKkhaC
hMzrO9kleyLvG9UKYcw0O38CJ265m5PGFarKeydOIeXlZTyn/GUizqMujAp2
BAQPfxmjamtzu/KHMEULNgdrHbmaOkOxYn6qGInJQARI+/AwXf4xPiU5z83R
CI/BZ5Qrw+tuypmak9enxPdd9IvY6IS9ejq2Pifj4ONhymasG5Io8V1Bmaxt
YxssUo/Bve9zPP4to4b+gn4s1FXdu4OvQXyAAm2txV8KCQW123pCuATPjY/J
34xqdOghSYBm9QaN5heJ7FbU1jQWJrLCB1jCskz2pgVmKWildb6d7beWeQIC
WRM7Q6AjpHcPUYHbJhaaCbvbwZV1Jlx3EJf4anQoqMXHNgdr7G1b7kHedDVb
Tx5ds/vWZoRHZKO5lAQYtsQERL1pT51whcn1TeHZUfM6bKF48jIfuxzKPRPQ
2BARtVjScLAavTDVc5gOI7N7Ws7iw/SiSyXNGvOYZrevFXNYRSlIluenuEE9
xPOrjRgFWlVHxBfiUsccQXadjdc8HC2sfnEbsyZEtNkD+04EJYH8r2MlG04M
Kj8CGXjjei3PoE2y8d0MWUHfKn/PKg7eNG+9tK3MIm0crp+nco9pHhPQQ34Q
Z5/m5RQ1twSZy5w6BsZV0ELHhRov/PbfRmlx/Olv2b0nwQ4HhUL53RjU8GE6
Gu84NuFzIhnAdt6XeSN69MlaejDzFu7iLpnpPdReyZU/OnP7o/OiKu/fl+fH
jjZZO2CF1QEFECDRE9MaWSWMENJ8i+SYe1AfDodXuH2+VgP5fAPw8+uLxFln
msK9yHGFsImSzoX5PVEBCHWcjx01Cg1S4/YYgyzx/mUZ0MhbVuh2vV1G30Rf
WqSFttvnJ841FlsVKPzPj0wT45obpk5q7uIiJBHPw7cM6mtaOlv++nAHJpOO
TvPSsBRaRegy8Y4ceQYyqpoEC+6+AGc0zivuyAA24Y5t8bwJjGebPfZTNzK8
V1nkIrek7Y12bJ5YLN+nr697jdldi3UD4NuwwPCqZ4qy4nHGWZ1NjZjN38nz
Kg9u0KXd3CU645fqjRKarvKXNyHylWTgdPWM8Qa5+xIoUbfga2MT45JbNSzn
shUgEIYqQPtjzgaUcMeovhuXidRyic5IP0ShLPy+7iLuuOVNynJqYXat1Tbf
SziOM/ipgWuPsXYO0Be9l053/TuJ/P2p4qvZbj9OrWTYiKbsB4kGG1syfWhx
Rsnv85xgAgnJ5FZ2lRByBtFFs87NbzOPNclMDRYC4ndY8YsPkpuRUDdnxYZc
5k1TbhhEb5AiuNrimi8D3reau44ZHr91uv5MsrzMzxhSrQAXRqC+HyDeWhYN
n8DWMoR1pyNHhMHYyPGtag+NHaOvQdRqd3eId7xHWHwk4xKLxTpC4OdTOQse
7jfqDFsugNZg8b7phWcgpRKhsHHj+YZyM4OkIM0GbJiaSobMbTrAm38WP+zQ
PVSDsDKr0A4dKPslLgid4YwVNNojn6ku2lRTQ0b2+Akaf3ZYei0Byw3v0iQD
5k87N96ZYGswgtzURZyX/lxw33KmFDxD/wpDgFk9bhedBgRW4EifcC6f+Ro7
xZzPOAat9/RbMMkY4LwBLL8383saWsN7ZTRktW6hmV/am8+eLahKanQs8TNX
olly1J/TIY7Q74BvafsDeQIieUI91dxTflFUD8Do2dn3pJrKDadrYm1Y6MhR
iTbLlyAVsTO29g5Dz0Aj5n4HKMFhc48GYq91Yk1Pde8NaNCk47iX3V3AyBa5
XSM6tS9OT5D/A5nWJ6dMCyMcdSe1rj4/YsQxmnvwR0ByoaqJ5NBKap+mXOSa
6xQAW+hltWSpQAjH0amldogEXoP0tXXBjJepaDjzA/TBsxK9cjxrxSMO347c
Qo+3ncwUDqQZPxd2dy98j//wl6Oo51q0VbIOaunWixqABxF8IWwgZAdC9fNV
ArqStqYEOp4M1XNsyTIr771FPu+3hJOYdDiZuPRCtuvegSREVhYRsLX8H7SV
t/FVW+YoriRAKQ8VrHOq7xfBgtm1eaULajyX8ROry8M24vyzwP688BaF1tLe
JPS9IAix3NGIs9D1nUI5Wd5fMLybOT601CzQ7nOgPYiweUVgHKi39CtD/wvu
eiJrY7pqJTsY7YwgqDnMHO2i48Gx4O53DTrbmdEkn1DLHKeSvBawaHOY6OFM
glY5GLapiMyHf8RljfYnNHdG5oGbDAuJMvrlU3vHclVkSoPUL2FFDQuyCEnd
N7cumSdLD5Cp6uUWDzjgbNQi0WJXdiHLVyUbDc5kbilyxNQ5AMNlwcNr9cR+
VF5ayVGQJFPr1uOP8/zAuvYJAu7kVJgI0ZI49O8r6g3FSRjpNJIgbuxhwr8/
jkw689utJlgoxgvniifyLBCLbZ3nfEHhLms0/GX9D0mxUKq0atcxfhYFL8VL
dni1t76Z/OhnbquoKb0RWZVEiTPDN3og7hkNeFZ7wpoBqGVr15MLtU0zJhUo
2U8YQ7t9mm52n3c1vIB5dtkqPyhZEaeie3be9Rz4VLol/FCFxzywHmiJamPK
FT9FJP5ZLLVS6NzEOpvaqmkHCXXWlcRqL8fuoTrmbhnS/uOk2E46vQvCrYRo
Jo+Sxbtz3bokTKYzJe994PsPXz8n6qj1CPw1AdTgFhhfX9Psy5nII5szQzKA
/bCbGb/aB7DAfZ4BNs1SES39uLKq7iAZPPRqb0cLRwqCIg5G8So4KDCexjvw
pam3NQTRRmHpflH8aL3+R6AG9k4S52NOts+1hGkk0OBP9RGY6hbi5aFX5Ps2
eP5othcDsmyvfa6nbOEux6I5y9wMyU+iHrD9Du4O5PCvaDwMPUHvsTJOGvDj
TklM0rRiD28yO5J4uuJogI6VQOJVununj9OKxFJk+/HaY4hj3ubHLanlNUfv
N160lijbMO5tiptPKWkiDI2JVqODGtSXxowAEmX45uTCCPuU+J9RyzvztHIL
ShgI6wmHzOJXbD2V8SpKMCYzxkmltlCyAOyAzHSPpBcZdvod4Urnamvfkb4n
Mr0oSnQ/H85uUQAYD9VnRHULQjRCK0f9DmsV3cgVrscvjTd5wypWWhcz/EHC
qa0O0chfcDtWNO50BePb+BtYDkM+GbDawgGwbJ+2b664pl2VHbCHrQdC3QC2
2y4StfVv9wkJGI9nynqEM3AHJSyArnkuw2E7j4+c+UbIF8wsrpKo0dtmIJ+Y
lFu+iYOqauKGzPR3sO9M5hEGlXGiRMhku/g1QYAOAyvqsFDk6JZuQuddZEAc
9mC3kEPI4xNSlyqQmg6XI39RYmKLNVwYb4YObPLRIcT6mabbzHIhgSYVMKYN
agJM13rBd3VYlfWYu9Cz8+dIWv60Adl8bo72W+BNSrwAoZJqOybPXXLodlag
hACPuZTQL4rjtsHISNtsTDNcPawLy6XGrReP/JXW0phKI6xHzr5wFqMI5xJM
nOKi98iIjObN1CAZJIZN9gO521OSwrdV4YbG8mUI+CS7/54fp9yJQnFqQSZi
py+ZjBiXluU66OwbTc1ZZAHV+uYLiRNIHLIQHuSymaGqqP7gsXyj4aFDS83C
7bXIEGR3WEHOcQEYKiY4itiYD8pZKlj6jlbXdZjO910RG00gHhCeeA2MuLf0
MosgHBB03Exrc/+hvUHr8m2/4ZDc134ZKFpfZLLLe6/prsdW8r3dUdykD56f
G4XBUJHCm7uinvNTVsBqEjSqMZo2LP5kbIqn9Ng7quk67w1IjoxJM1NkKvWl
Y0QjPsYe61e3Y3By4Z2egekglSx7zxsA6Av5S1lYjl3jvKCDG/XRMo6tOI+9
gslMgfAuAwbBelOgewRudXk2munUXz5pNUUn1YWcFipYc5rpn++AeZCPM1x2
pI2wn28ulCh38gh+Jaa21HZAGBl9SQny6UcmTUJHw4cfEdMuG8Ac983JqoRl
KEx9Umfzb4kcsTQMHQAOXYYR5F8F/z4LUrOylNYFxRMwlEHIMuWeBOa9F9kN
9pwdzsgsRC4kOtWqRy5thmNAGj1qF0m1LxXcIg5cQ/Yb0RLL0zD9dttQq1db
gMfyHd5Gck/F+6FdI+4eC1482DiulOwup920OyPl2ZMlM/NETfd/qmO/Khts
rBW88meT9u8p/gO3l2mZ/uUQkkxM6aZSWAflvHX78UFocNRuIS7UqBpnjecj
MouvP88nwLj/VJyqMwpZ/W5cWo+6dLIKh5FmkQ9VSRpWZSilNz1hd1GlLXYf
/mYTzQeLRA3FQcrlsHjaLUMLaWeBzT/i3EStIfQiwCdt0R4N5ygyU/a1NMqr
gQ4hFyjQeP86wWy5RSU2iMd6CaAnjfuAT8FhADjVX02b6usj7uUSd/wEdfhN
PVSAc1ddAt3cJ8S1XJ32U+qtb0bsl2n/JAGPXdYT40h4xa6f6b5UawOyw1re
GfeuXj7xXRthR3+SSV0lcuZW2xBoR3bUz1p/dy/D3hdA9SJD3baVH9an2rPt
1AUnwHoDz6n8XX4bLDEGkJC+II8d4YjOusQe+kcFyqwand1dBHUmylBLxzpJ
KwU6WbLh7DSyI6YQPgbiX14VTZ+PD3ahfI9BAtPC1lz3aox3+Jnmt4oOHPqD
jLwH4/6Q9SKKBwcOSWcxP/EevwjH9uDBecpZYqQxcKohDBlfdCpOKtl6xYkP
fcrzjLESycdluwN2otaSYJZ1jT7J3rYpXPAJjUHoYMZe4mPfA5stNt/SHFgB
W7hTviOTmlAnZJNDQy9U4VJDDauksyOIrfaqRVlrLAg504HZrXCwEe69UKzj
5rLMl7Jvc3yT7KKoERP1tasgvrOmaMqdDz8laRdAZbpDp19Z2fBLl9ppW1PT
SajH7AbVVgJKxjI8RAggeDEdR1pIXKDri/d1m5282cIhqFx4nSYN28xlQzk+
eBeDWIXgRvvYbGwd+dVhRu03Wk0RfFKINqUoMna18MXUxJqOusREVQ0/dcFP
uvTx0VQ/rK09BgvCDC5xF/Mh0eGttDNker/5hVWwdx022ZOMOgNifxYGtefd
PN1fSQalTWigE54IUwVAdp3fqMzVr97IkIIuOfwJAcaTpqKXZImXE3eOLgxA
fpgqPYrc6SgXcGzbQKPRp0nV6snK2Hiz1IjeljNK1QpBZE/6vsJxnU006FC+
HoGz6IgSeHvPLYzFHcdCXlPQ6/ZbPiuWqddKsnxF43aRdQkdAD4d3fCMZut0
ex1jhqUqfMeSx7hksOu29uA1wdLCigNinNTSe92MAXQ2VDMIuJ3VkFE/qC2P
rpYl/OMv3uhFIkDtjtr9AZ2Gl+39AegFIsIg+tHNrwCXVIj+2qBF+BpPr0YM
5hzSCiuYyMqKxAYj048Mar9yAcjamqVOy8FHDcCd15N+vYkfGJUC8tNDBplG
WqoFAP/qZAnV8Vvm0J/lyQIvKK0PaybpaGVtksZA4EACRsrQ1Oy4qluLJRPj
/iDhNSkowX3gau6c6zVoCzoQMSD8Th3+VxB17Gwi4YGGIViFFp80i6Mi/s7c
Humldl/nslAzBgqbBOg3QexiSUQe6tef+e8504oNy2ek+SlafZhUUEnTMSjK
vEEnCWJreysZTeMZeKRorv5uSIrTnOfzkl6TixyHFQbSIVIW4qnhIOHX19qA
PdfxX+CjR7BdefYVpe+LT4uIyb+2VrT7icuxTpzvXk26XSatXsmVpN0nQi5G
hdg7f5YqzHRtjuIGeU+DaN0vT+lCWutAfhBptpMGAuN41X3kXwtZwLzClgML
PtXZiOVjCSRNPOMjnh8chwPnKlYT4NJ0rCZmqALFBaetEJXsq4YrPHYPx/My
+MmFaZRctfWfv38kmb0x9NqqhmhX+rtmxlkQ4DTL/hnBz9TbmrkDcDWbh1wJ
dnPku4sfKAhFEDsVeoiekdVrjvF66JbC1fWXfzDVj+vHr0/iI7K6v6o3XdGE
/EGh0uU+BP7naB196fK44vmzWZOQEGm9dsNrMJwtOpNO1vbaKBj9p18CqbMa
97FoF1gEVOdcB7oh6IknpKj2FDCSU2pyNvnAJjx7cI+J7WmHNnGIOOR8+hiq
WXKsKdf0nEB7wVZAOycMndDg3Wyx0vCn5RciOz2KYIQZP+KRj7uCO6a8NrVt
sARL5wIQFPiPD0G8OtI7zzE28VpJ2OxBa+cjyg6DV8kKT7B7/pRG9rhA0rOC
2oqa1R33PicUgbqsnIsl0CJnKUVjDVulkSGXh2vRSOBqUdk0ykrkDXnO0/2k
7a4WPX+wy8ZiEP+sOGI1EFw3J+9osX4PZYZ57ZlfkLS5QY+uJztlZarVWfsc
xwjvgfgBfCm8KvAF5hIbtbHJ4qsbLDJwG1V7CJJVI8Do/MOlrdXwBCtSot00
z6vZ8dojm0bEpn7iPR/Obb+7GZXaGcu4HYhXeeeso+jjdSa+JavcSPlvAbx2
FoTQ6xHs+Vpv14ZQBNjfFYjyEasWqe1gCabOVbljSOjc8m6U/ifF7LMN3eqR
gHaDEyk775HaJNFW9fHATVs1OGZZPr8VfSpOQhpEeS1oJ6tHvDu2V0gWpihI
A9hf7KoqO1DhCXCTDYU3SDnzE4XD1wNwz1Z+J2qAZ6DnUEFDBm1LnE3KopTK
m2A3N5BCa+f4z3mR+Bsee06x1DhW8UI+exKTnLJdohagDb1TYTN6BqnYcTza
J1HOC1xmcrSgjGmN/iI4yH8fGKjDM2YE3pE1dqLwjR5b/y89CTnyQNhZKiLn
c+p+aID6zIWHprxgjlUhfkx/mCT9aHJwgTePfVjkYoX+lcwnq7IMAXzjiX7g
T/yKdo7spQYYU9NNGmz7/hRiyG8qCmq3zNkJvVsAx24khWzwty+eXNgdwIvC
mDfDzl6bCyV8eKH4fILuFYvUYR3SuAUY0QgWeWt2GDmx3b0PeLlnV3FY97nY
IRSGDNs+p8sIirfefmczRJdw5X0JKVAtl5ekuqqqH5XhBDr1GtNcW0ORvPtP
mnrWZFvaSgcO3vsLm7syUFO8vW9I6rDBo4I5LWwBMQA7+xImCq4Qgl3BHNtC
ZXyPVxaVonBqvUEp0qjWkIbm7HuFeaTJqv5dcbH3A3jNjne+e78RvNlVBcqQ
lk9fR/v3s9KxeaRJSV8ckYbZbvYvOCxt+kRcmcgLv/Kv5x4iOhkNATnndXWv
lYQrpYvXmBIfXfWmTsohRpQpWxFi1M0lVrife/2hg00bquL+C08YgEbNT78J
LwCN6Q0aWcPipUQu3lXNM6iLfcjiuGKK+dOR9E4JVjDDI8LXcO96knWg9hoi
G/ix7AH35UfRDSDCg/guXCTP28/kRqhQ8QyjVcdFae5tEv1401usrP0nF/WR
/WPVX6WerrMTIOhskUGfncS+pDQuAKZCFYDCSzoDnDUSsRgGayK9dh7OIfNR
hvjj2GIwtG0Do+cMFF45aRQGInKfyPrjXWFhqsWwXkt/Cf+g/JvVOGuZqrE8
yQVbMN45X0ZpFXuQjY/7FdxlnbcauJrfVMDPfGP1nDMDo5EhIBxcf3IcHxM9
GuTWwLC/x80P9FDJ5TDMmsaW3eifHJKYFM+Ha2/hm3jNaG6epL6UATj3/lpv
zyqsxRofaFz/jXl6VyiCasFJJ/duMaeMABING0cxWnQnEgNb7e+KBE9CBaTa
U/DXVQF9yKNvWVtu6ZIVQiwqDehWnB7MFz/lwWMfsUy8L+pa9xuw8aOFKY9L
sxghfTdRa5K1mx4LT85qQBm7fwPkCoORnJAkLOOmiv2L9wSW5J+PK7Z5+e9g
o1QbsdRnzGGxhqdpDICf4fmXOQdM0t2cJmoM0ohvPzYZ+y/Rrqu8vpAz2f4s
KT7acmLoj0qcgas9XT4Blh7gqeZ8nbz2BYkxpE/4Vv7yRJBmOGCHShpQD8N2
+LRSZGNJK9i22qHe9ZUoT/IwrkP1DrlYDVQ//3u+S6g47g9OKx0qXInVwX7P
FL0elZ8pGge53ZAp5nT+BYTcidEi19aI3I6HfxndDsdP/vnLx17emQEFW7FG
jbR2YbWm9vW7gH9Ds4IXCkrKbRm7u9Ncw7/4cVgYtCHOv1y2UZN28uF7sv7H
jZmZzNKY2XyfmVfBtLDDKHTVo5D3yYM34CRQDvbZeLQzxmELNo30vao/0oDT
SoyuBuyCeKgFwetR2Jks1IxHCIAPwgRNcMxdRreK/WE+7ok8RQE0kr+oWq3V
FSfk25ZeFYWd4R0q/d/ZJFqEc3f8/+zXdQ92JT02mC9YKkhC++cSgZFZoDwc
JYeho30Ql673l3yYRxGRJQmfZdTr4imN8olgzrTS4U1Ok34EUebO7qe+qweY
yp+x+T+vnuBZgtrbSD2XGYDwo9jpMSh849nbNX10S43Ae7rv1MaWuvfG+RRh
a7pkye41qYFspA4yrSSF66WsNiwljQ1hF7yzHos+GYMsgAlIEwstYnHHajda
98+NP9ItyC0Xzhiw7NSkLUiILz/MPNYj8CByTi4td9NZ/Y3pJgJKPBg/n0C7
Ebuqb4NEuNUMKROsnwYOcMAwlhOqmkWAsjuWdMmewQ2bW1hgBAajHOf1lVCc
F03a49aEfHIJhWM5nsUq8m3vzawkSKFuaurHajiMCTra/2TBRfjg409yol6/
U79v8Vvd+7EGRn/DUE8g34DPfVpKd9GLvmoXsJkvKby+LY9tVs3tQtPK4FEF
r6MEXlwrGw8XfII4uj+ki6Jr1fz4kYXYBaq8mCkNfDDze7L1GspBsaJKfwhb
mqd/eaBodmt8fSvwfudrAxb6ps/QjtU4LdV8unnRMOR8yCXPxltWShP6t7P4
/cDFLRGdsGJcPZJGebqdQTdRBxaccG6jC3M820vFjOqLFP22SZk1qMrPhiom
88Y4oVuCXp5YI3EzHoxfq1TuCd5b1Eg50q9+VWtOqH+xVPwje6fQ2yJoZeUL
uPpbFW/TwTQzXXuysbYQjNDoM1QqfV+XKiC528QJjRRMNFxTSCoSW4LiRO3S
f+TpMq0AkbfJwd+k3ZLSjtya+h/xxbFhhEC+uz8YvRNzDTBGPL9UKf6SAfHh
naRAmppm0lHg7Klv6g9qkKeJtUNeBgxV44Om/MxcGQcAXm86WpSs0jZdCKc/
fEFfBWKWtCMvWXRFzU67K+K9imAt102UqCTW1y7JHb9bP7VZghGd20SCwIKB
bLeM4iDYeuxWDN2xeMNaLl5Sc/NE34bq2iD+QSzvPZS9fxSTPs5O0vkjsLTs
EeFrX4VJR3G+LMM5re7ovT8leDFW+kuuG76hnDHAHo8gjPYwadVrA1ywC1qR
MovbY4/LKXPMP1GKV3W9tgjGsxh5wxBr0d+uc7YHRNTBUBFP6se7MmBbhQr6
mO/CvK/TkcBu7c8hd8nFoYyWZl2NsrQTVpPDXyiFoid32hiDCLyBwv288ZGy
tP3AVEvMskeY+qWXuBExqfvDkoAyYuuHCj5MQe7Foiw1kcYnKuUTHiuNWq0f
dtvS2e0z8xbWqhJ+WS5KU/95AsPqdx+SeLw7Vzb6pfaMOWwNDX3FNdOLuDbe
NQli4pr8M/6b4tYRYzyApIv+esq2/f1Iz8EGPlc93q/wnjBO+9jt3b4xiono
r4ksGjDY83psFLIcA8EHBgJHdWJWNIJJFuf7VUNnpb11b+V93SUPfyJNIyK2
FSBLmK05EomsKvucKCxtpJ8Az8LZ9RcHLGzUuJgTsVGOfUdcK64oPV0nsZu3
UFERsGN7+9bj0WDlhKp3i74RLoXBsuqOwmDDyZlknPeYSsUDKPd72/mZPlYu
Y+4ZaPGZPtspwxb6CSfr7BRsoH+SxRs1eFIdmsUtX8fAMDRDXgUsvjSXePjO
GTSGCTorTY4sBm4DQFHc1/kbD8IcMp7ECiLisLpQBRVBewU2L4TZqzFf47oZ
OH6ceyfybszF2yyN3OQSWJL1/fJ1gRD6pOFvMyFV/evqOKAGRMsUDPaF2B9f
vthfGlw/mfWa6a6e/jPU8ou0ylEkHDMe9YKVL3v2EBo0DFpAmMe2i/9gI/jt
NzouUi4YTSYlXnYSxLGhCTYQxGbyBDoo4CeJsZQb3ZPvLI9yggDSB9WjrMgb
X+iYizgjU05Sgg5K2J3nk6A/MM378P8JeebcXLNxKj5TDyybOXu2Kqittj8a
yEEm5tBInBg1AxfdHzwtU4EkCB9mcI+pZhWYYh+g2CA9fCp68icD7lhUR+W9
idMuGTP02z8d0Lj2UQdSaMvnhXMEE2mC/nfUfW3dsp/ZuOsGegQ5wqXciWdP
eqHJv5k44rEt/8cak9f72tOfEMzteknulcWQLoZbHUbmyki1HAiwpqMXtDfb
QtIMVH29XTnHgdLQyJLF5j9wfa9oX8o49vWxt4dRBsuQxOW3eQaBQxf9cS0N
Z0RWPLs8cOTLuqqRscvmOncSi1UlaEJvPMmX9ODDMX25VT3oDbDUSi9OYVIl
RmkLnQxFFs8YthW/cLpZM5RZ0xC82FN1tOe0uG8q2hZZgm5qYyNloIr0BXgr
78faAimyCnTDQL+Ds5KWXq4ttdAt2Kn/d4txt8kagbwY6lm/OMV4m/SlvzFB
dCuwjCXJ9StbIXQ4sXIIW3h4c2bHKCF/2AXnj374u2inHmLXUjgXNtwqgPCZ
qQA074JMERvyGNZfXtBjJKrEK5k+aeMkddTI2S7VKAmd8XFv8un8w09vV3m1
jvNKAxkGJt9kFImKMHQ2wAfE86Uvk5K07v/xV3yLKW+zSJcPGOlDBMRNy7az
NNGdtWlQs455Et0IIuklFB1okyWI/XNvtone/nyMVRu+GXknY6Hxdt/IObLx
79dReY/Fvi38tnSu3IHkdE6CdSAo8ZIXhhj8HJSshmcuNCha00rBbJANOVye
XemZn97wWBrB60dVpuLoULhJSsnNk/OT7tmuTGKgkZyvoKWI4WqGyEz/D4qD
9+U1uqST9IFnRjCGjr6qy4VQjlOjkTh3xY76rvkb5XOwYKFF5xmTZPhhcNLB
cYsKudfxbAHDff/NMqsCryr6t39sZUbWAN1RH4HOcDEqld9TS9zT609/GZ3m
Lvwe6OHn8AFhMGbBHGI52a+G2rMmB7xEVQEjbmKqD4EDJGASaKdw7FkOYjWd
bXpYRgyTJinR+Je3go9xG9Ur9b1YNReBwQkwxjt/nyrFNNsmi9lyZsQaI1Tj
bJmzwG7jCDIo/7euFH42//Z4PMjq+HcbthJ8kaMNhr+TAHpZ+LMR9Pqb6dzb
U+tNLNG73jrHQGqY9YalkCrdaPjm+rS0QbACpDGce2MsCFVcXYxaOam++oV/
kOk3PkdNO7d630xYNBK2sVJs1ppAwxaaDTodNcR19CmcSwss7H/Gt31oO0YN
3/hry9wgXmBl5hkyJ80jS9wd6wvuXiIQ36BLH9Tg4wUu7+A5QhTKUKwA1Crg
KARsMdbNpb6fTJxB91ukMgUJnB6GNUaRsMl+N2uwo52kniwEmq+HLkrVMTtK
WI4jEdOIoifkJDvKkNUTuEQVMawe7m5Apuq1UE8AatpgumxzBtU7KnFHCqLV
P1dxWgxBvK2KL7oeF12BLciHhpReezmZyCJnlhEVBuF4K2iAY1/mjm5qfBC+
bJUFe3ADi5V7QxXMnROvdDTMc4lvQMm0bnNEOBO5jhuOG+9vJIGgFQPqW/3T
NubnzTgICDS0Gycaqu9ERS6Bm440lH7dFdv9XSqNZlLTiS/9k1fzuMC0RNJ5
TUf3QjoPlLyr6EvHMqORVlFfuRyTUSHu5dG7ugCSYxZkwnwBc6d87l37yAmt
CEBPwu2r1D+qEjl+N/A1GxRq2/YtMMK8LyDZhDQcGRkIN75tzCMCZSY0FpN9
ses765Nsc8D38F6bfOChiFWmRLscUquBwXmlaeVsfMz6JmmhKcr7ezxGY8j2
t+BOfONsk7Ehm2dLguWHvIYbeVQt0VdlNugRjFZjOpz9CneluPDiOCZ4+b6Y
stG/25l8rKRYkFqYuik7Mt9bfC0UPn6u6t2n+LQhTKfZEEpN6pVwOisnAB4u
KvjcDfbCjeww7u2686pfn/ILAVfzNnHLHL26ZXLSfK1V7vJSS9ipDrQxju9M
SjS+mRCAJoXc2Mdid8OCGHyfi6Qg3OZpgruno/lGkZ/r2k1lRX6qX+xFby6i
tscUcKLZhruZY1JKSSyjZGsTY6EgjuJMfMcxTzj843SOwPSKMRK7lZUstDER
YrniUv9OXytOfnTiUrBoiILtw88OkIEyQdphZ+dW4X+x3zQTa+PK2Zngk9Gp
E0YY6ZHaxjfdJIws3U2f+XrvpDSTI15Hrq/dD6ZlGAN78WuR2rzmMYGawRld
JpwHQ5HrmHUMLoLUbK/sgY1byp6nChrUREHkLIA1hAkfluuE3p9IassvzzbD
JgzOpjUTZ/nYEFrFOxeA98SguqTztxwqsaPy8KrQdeagw2QZX8tBoXigmPh4
n3dUIq4Mys1xcPeBmOyTQUvIjfa1oNO0X9uPZ152+d4fgek31cHKdbuQIyvU
/qqriGD88oQ+imiumgV5EggtcLEVhKspnenFowY/lYTbEDV576j/GPdQAX/p
cWPccBoEpC61VGEk5AJXpF0IgYl9msGRjSxzaHPbRxaM2zLMIyfppelgpyas
qTCPN1FfkLxjDI0NxJVbZNwPcVJfwYxHGkcu/a4ZtFq87P2GOZ8K8j6BR8Ym
gbZYXE4T3XtmgTxma6J2H1IB7jL2VMl8WJ7q3YzGWeM21TGIskOioEQC79YG
ZIrweyIlzzdQ9U4GUrjYqfkUKSkxzvuNHcuQFlCbJOF6/plKj8WBZUKdmjRj
LbA9MR+hM2QhS7ngg4+buiax3S+TEihOZfvJCtweTqlLKHL7tyMQSaq2FFdd
FpT0OM65+ke9C9/GkLIST0x6DtGlrU3lzqfdvaZpU50U81BIDRM0Mf7FtbSV
Vchj1pnrp28FWQdAPi0D4GOnE5OY3+Wyjmaq0oAelKQiYO8cMbr3Td8mp+by
Dak9hr6KtVzihh+26CNnPFKMaUgRYJQKY+deRcFbV9jMcrbAYoUastLzss4e

`pragma protect end_protected
