`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
hgid1VBwEDZkd4Ianf3Blf6bzI42Eryw03AYPul+9v5If4hJXQ3mle+huIxq24wP
4wGWVnBkMom4uIWgRUW752jw5V8jRNw6M3lFYbVRRN7VteT0DXgZgeR4TXY9QrZq
TJMYPnbcPKmkaRdjB8bjsphLYSa8/l+4JLbXZMwldSY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 13088), data_block
peenGVuYWOKB0UI0f43hwnJEmkLnRWO+viCFqVkIAU8IxxnT9AM+KdJJVt3JfkM1
l2vE4nWISalVPnE3HQvfP4u9e/YEvO3NmqVvJzQc+iS4wzutQN6JUKsfifbcJkLf
qmAqPhVkQO4gMmCJgfxuCr6BhOfxMcE7LkPpIEPV2p32pGNgw6BhOcLWHuC7ycaK
TOUjWaYcE5iG7RRM9BLec29vQ9fplRTLwybIOwdQcjGtBNlaLqQmBz7tmyv845NL
JixHhSdmH8VVCw6eodCOIsffgjyDbgIo+XISXIn3KuKi+vnTv4L92cYX37/clr++
a55Ip1QtRQBA2ciPm/LiiKyJkKHXu/utuTulMqVlXAvWYywRG6OHfoAjSvDlQN9Q
UBg1onDmwy/VsLzmmvIfaxMIm2KklAGOG8prNLa3nWyBErqd9OM9WklHQTUecHeL
vK+wYFAnp9j4Pcg0mequHtFwsoiFSFv/fCrD+qzgt/wRmeUvED2xOa31u8I/w8iO
YR9HbwDt8/o6XTXISi3bZzr+IRL7kVQbdpupvnP9K0bBVYk7LXkG8tirJC1C4o28
7Ef+BwmZD2GMKJ4NaRUjaFcjsMP4pow2Hh0zUEOynfZxrsCkMdtp+DCyG0YahQaQ
xdb+haqCETzWnybPSfJ8/5dYOewsel1corOpIbnECj03N2He2AdvqozztwRRJ2wN
lPUlFzo/Iz5qRhQTlVHy33q8rcJ63RQ5T6ay3/S0buJdx5cjikakVlLMfocOqwLM
wa1CKpCJ2hRa6nIqNWlGBcW7B0BsFYkZQ4/R/aDNuTu+5iHsLybQ1tYAJD/0f8sk
rXP3Fgg9B7VBfIUtMLcSU6E2pU85QMGmW/HGXD44LpLZ/285FKHr4SzPExxulMsk
bvxFazKh9CcGI0lVNpLBWaCvjVTRCoif0s4dQfdRC6YC2PAOZRShmFDcK+JjQqa/
4+JOlJV184zgx2McQi6Uk7XJkTtOyiK7adk/HBDzxo6V/884YlZpX1VMQDZoxagb
s+Ptxf21/zpg6xb5rBekQd6LhE8/u5VSjk91gwlwXD23arYfes2mwi4nSMW9Lymd
wlWtrUF7uaovB3Hl77KbA9/kwwcQ/X2YGymPNITupMEFCvXZFSloNVycEW4Ip2n8
H5kpgrUXyWBrXvBWDpLuUaqghAqGeD0VU0vWCllrDVRn5oRb1iNJTO5iGLo+W67+
uqfYpHEjdA2Z/2cznSy+XQuJDAOO8eyDkkYYTbV9Ec7GotAG6V+IPPsm/Tn9wSw3
3qLsL1vXGB+n+vLt9WwnckPZFMmj0ePXVZHs6F5Ld8EIQevUsBZM+fNE6ZTMiaHI
nt5N8KxqKkFh0QAAyidWMSknFWMKQEpwIZVCbrBFqJrI8mtbA6ca6//ozgaSx7fs
bTvodtUumuSvQvgTzqoMZcY2BjLKiJWrIgGI5WovAjyziSuIG1ttijEciS3oJaFC
XAHfeS6cqOBjd3GaeG9I3Q1SBRTk+qIQcAiqNMsn7PMg0eq3xA5i+QPkIcn2PbYp
oUPBVd7A98SJstQ2IHDsWQNEhsW0DgydZ8FPAIzNNkXJi9+PrztTGCsvSfr7imnd
xskyPoHi+Hy7Si57vTXTbJnSj1mTUWSZn84KcvAQfO6Yj2ewU65fSVD57lDimGwe
WRJ58yJGQz75/GDsIf/EdfRFVZqELfb/3yK0dhAHY97vLHXFOfRsg4ck9UoJ3Tgk
Od4uJ7vcpEqT6mJRXfO9LD0oP6+Y8igZ+tb7KcOVU8lguJMzMqbfwrpZijNwLoUK
Nn4HGgOk5P9pulAQbN2l8eqKaGjFtEOWfwtjow/bIeBmYNhLqODnG/7eUIJDoAIp
50F1ZyuvLdtL85Jv6BWXktBKPOJ9ov3JdflWEKc/7TSc6BP8eH8LVWLvtFCXFX6t
44DjvbElrEVeVk77wxY6ImueQyUFY4H6NNQGKdME5Q6S6cs1w6dtjcaOTbI2K1pW
CwuKy8bVmNBuMtS3k21Apupc3TFH9chsqcxMjHNzdJ5LrU75hsH/UG0m5mM/2uUd
xZCJl3t/roEYdfa+2jEZq05LoXsngAM7oRfEpZSNYei/KIBeSaYqfiR7Dzi+fZ7H
kBaZmlJacEKLhpx9Tk4olo9KuOeR+grssrd6JXCeQ2BVUzqm7IqODNL8XEAf+fmF
ysJTb2+IUm8J5kCU8ZK4D+lyuaoLIB/47on+TadHoreau3rniEh6b1PmKj2fPQCi
RrUspt0B8IqVj67nuPZf8aCjIBUeSKbLHdXbhVXCScQe5y7hmvV/bLb/VN8hT911
b/R+UPvyHlOgp8PYMzTUNL/FN8EgCtQwsMoJUSClzXsUkQzHVviJ8kmtL3eYZtRY
bmpjDXL3LfFuZxKUXJGCcH6vfXn/3dr4XKnCWFV6voXzDuNDD2WaaxrL7Wy75S1/
G20woXAYmDfW7x7ZOcU+pjOvoxLQ3wJQ4USBI+1XTDZG+SK1fy6GSKtCmEGTXR0H
N7KzITOxBqLclqZPGTZm4HKrrpxxECSzp9QodZOi7Pt5Blo5XTl/RTT61dgR4zRY
9H+zCnVPvMm9czjWyKyl5e7XcLckN7Cn+1AWIT8aAcP85u21uqdpSIfvq7UTukV3
G9Q1y73R1qJhRXXSnKyu9KKV3dJQnQ8PoaygjZZ/oQV12ReG7w2LvVD84SWEj6SQ
rZeVGXi5Da2vnaorWIO/j0n2fi/M3V4QF1tPdb9gqJohkJIfhCK12EshqrQUspE4
pDDvBpQsqYan8y3QVtdxLMW9FwOgKRpV6Ewcsh9IeYuNH/4Na5KGWlOqWphYibVQ
hxUitrHQz9gNPp4wNvSgz5ZwvLkWxm5+AwiKLTymu+tPXI+Pzv2tXB7iLft1PBKh
LjVRP4CLCWLS5iz8avzGvLTF1GSPesciBa1kh/p6J2fWr6PoLFI3wC7U9ZiJS+pJ
jvJ3rOa3R8Q4obtv/QX+nIp4aVOJmRUVH5ajFZilbCzDWuGsmq041YpEdg+z65lQ
gAetS1MTaEQZdmn/T4HTB1OHibBh8q/Z2Kg2t97yrOewTgqoZ9NSRlg0lJxHb3cX
v4qb+woBZEJZhsADU9/p8YAZrirgrwMxMyiWGYCtzH7qPI10PYevRkhD21C1ro9S
Iy3jK0/8bUVEbDJdkrAIaTZLrZxB4SSWg4v89GZFAkarfLQFoxfcuBhB38V2kKE/
N1Xaor2OpR+C0DgAhzoNEsBw2ZYuRIHNGDt/Tv4qOZSTFqsGPip5ROFGgaJljqVs
KeqaFm8ClUW/x+WjlfhOeaCBn4OCw3QyzWPG9IWeKQeV4gNuWnz2/VU9tC+FcVyO
Dhbkrw3WxbQKO05JuMAW/cq2SjboF5WpnHqZqvcFSiDvmTIyMtX3qGNLEnflThuX
I4hlPTNZ+VN57ij0dKxsv9qhDf3eMASz7gUORwMsX0Wu9uyT95DN4NW/7Om5Bevu
pXn33qVUtqObQJSqTV5vUQxuIuTUvB+Ctg6VLYCpUmuxvmuwF8tISQup0oQN/5Pl
byrlXce0w+kqL1BFOzwbfGzM8ROHM8LvDL8VA0CE0dzTDmwpxiqk4Ugznoviz91r
INlGjxKNUzwc8H1mPkZnR6FKgAd2wvuPdfqVp24C2D68Lf+bPnaVaotHIAA4aKwP
lCmkWk6oXbPk1/OD0Pk3kOA0CIlFenjqzX5VOuB9tQ2rxFYx8b+bB8WycIP9SfM6
p3RXFZ7t44Cpw/rd9PsbVsrzFKbRuYF9l6nHvry8xsLHAs5Z8lIeBtmnhAfCHvsF
bWsWULL6eDIz2Y0ph2+2vRnXII4rOSLsG5dM+Q41wqMog87usniaOi2APb/0bZK0
zLjkSFBKROJ1C1znfQIjgAaLyHCO60GYNk9L8r2WJPLiU23Xg68J2iikU4Y/0qmC
OFq6bAwnmG7TQFUl6n9GejaJG7Le1M+RYhhAtqEE8SkU6ZVrPDpffLUHnaFbGZkv
BJ6Pb8wbAWAYZcAsfAuWpbVg9g9ssqg2NUdLoiIrEKHxMypIcuPMY5v86u/WPsz3
APYs4HcKH/LdQNw16ckvJrZ9niIkiuAMhsRja/nFvMsMv7rfCpLRh/YaGHU/znd4
xVoremoOAaCbbX0U7jerb4ojrkOaJCWBzv+ISEunjSN8v3i+azpZUETWK1d6mpP3
dlxsTBicDeaJOKA+4aDysrmYGLMzXgDdfjMsebwJ4OSXUjwQwKLhSxmTMdzDPspO
vbIVmRyo1+CIa//UHuZUSXQX2M1NcHkaMjz9txOfOAA0Y8urVBSOPD53SbGwPHKY
DWXQWrAaWHwOfnRecoAldVKDbmJIck/FidVQtgnyM9oIKnqYMjhzuyaiCuf68OGg
k2vTLxC/E0KgkC7xCv/hlylZZmKydgFmd1z6eAGraHwMTxt7XKNdZEd5eNik8AZg
7Ycj5Og1UjWbUV9Hb7YCNvU+Q+qPFKHZIvBALAAzFo/xj4gBCwpLVUHdr9OeuhG8
MZwxD1BiIi7tOwohfpJg0L6PpUv9zLBbgSZbUir9hfZoQyEmZY9EzxszNu5C0IT2
cN/Wv1MJikHjTRrJOwKwCHOgBcm9XSJCw5O5GLA3hKq4GDQdGivpBvRYRFHI6Vy0
LoKmt4SlnrYRkHtdcD0Q6ASvvktRMEgkTWTWPKtf9yNhefP0YVlfg+eG6PGyN0qY
Gd/HyKGOXNBX6jB2esn9q0fC9QCRY+kc6KbwGQibSWetFecnYoUP6Zaf8r3g1jQu
6LrQjEM9CL/XgFgfM7uySWLZo+P8Mc3MU/mg1eYa8BxET3mBLprQPzWZuDtWPiyQ
IAofyUzEGXmcRtizuPY2W8ElGk0rrGcqBXvTBEXFXrtVwJZOQLlvS5a4V75i5ztv
n+qFZDCDoOjBwOrPofoZtrBcp50vsFAJYDOTfER8vN580AM7uB0xZ8nUk8XFV96E
KbuCgrg6CvYGBxIJKKNOElWFjcYxouVnABPcN9xsw/fNAMKx5dEFW9styuaCcxcg
uvWCvem5MigWvouYcl2aPxSFeQlN81h9VFDThW5RPxTuUk26iAXNxq09JKC992qQ
Fgo0r+BAQoZPvWuoDBl+Pf2M67ZK9yDyxsm8La4Nk73S4cBy/jEib1iagEJQP9R1
5f68TcpX/eHeSBMTmJhClqsCGnKAJYAzvaDQKCprqllTmRxGpKZcDqsDlFV/HBAY
BJJpbPTllW7iTzIp5U0FvWaAoKLKHmRNWNUuLuFpf1lqAv2QMHi+bKW9wXivJteR
KbanVOZ2fTr9illXN3uLh6x+D1sd6Cfe/R0hUks24Csst14i0oHaHop/pOMiKqWO
jl3L6IL6j8PJQmzUdO/hC+CNxGExQPhB2fu4myYAo1qYVJgNEypM0u+ZIHIJy7kx
f2smBvCVgfqgddhlC0W3rEseYgbS69f3T3zWoKc43RY/iBeN0q8LkEGOo0gwdmrU
UY7fZQbFC3VUw213hTzTKq4MpUGr1qQlKtvVUFgtwUMEhitWd8kSRPSQ5cWnD6hc
Vu2RON8AO1CCtoNBAlQ0DXk02OnB/g87/LGLrYd8cy3cpjf/IXoCwKpLGIv1I9lO
AEtI1k3FEypJ/0Korjjs1DctCmJK4CQ/8Tz6MvNoif2X8OhNCLNfTwxvWoDEo1J9
MLg4FenORQP+LDoqCFgQI5TkPwIOktuL0nc4MrJnJ189r1XrY1D5ApZVqRSCSDDM
6k0vcoocYpu2gc7ZmeDoDjqnQgx5jDSz1U8iC5EUM02s9A77FQxWlhUNdF0Y64nK
J+kGCF0MyD5Pq2UcZJVvZA5V+T1TivagN3k8mPVih1ZpYqJ3L09CWczzV43vBnJx
P9cOj9AzIzutlL1AvWreOquciUrTq7GvnfhF73+/vYia1ztiB1jzO1tO648oH1zw
+3SVPq6FtqeG5MUivH/JuwNGteuyQ+od+Fe/0HjyFL1IOSXbHTmLQQhGbEbNOF6b
Mys3lzqmFmFT8RFbKAptfav1iHMsOekYkQcdzI0/tgl8cRZ9klrqyMinnszNeiZP
5y7g5Nv8huNRnF23A/hI8GsCvItbOkWQdvHXpceox9604Db2fAnP1Htf6obzjNgJ
fXTR5Z6bTO4N002Xp+HJohbMwIgWgXgM/44NVGoHWbucecJ0jZM3VkkzQXPeVpbJ
hl+ndOr7dZTEqrx2keRzVmvUwzjc4iHKIiDyeeJUOPjcM5BadzahNcKI5ZAVrRT/
5WlV5xLVT2+i3Psz38DV6RjKOmA1MKA1q+0zB4KUQexwM6dPt5rkhsJ2F8HgV//E
JhRqeRLh2UrggY/Gtl+D0MlL9rLdhmm0PH/Al2/+RSq3CekAtTgQfuTBTrO/Zl2r
etXoFsZL72eE9fdMMoNwWmrrAw02WpngD2BMFgVJod3nnEorjNAKEEvRT8kU3CEQ
XIdWG7BPTx62TbaRE7MrVH7CMKH7/EOLkrr0kUXXLNYf3XOcfs94XclHDRi+Ca15
i4D/aDBHcq64dtYbtYqci4cd3T0Gpe9HzFRLswOpkaDH555BN5A7m75/jSrigELa
d62vraebk6yhJnniuM5qJSo/jiIjq6TDy/hOFGNL2qFAiXjPd2vPzabca2rjS4wS
PjE5R3/xPz5G1kFVeQVnD2svpPo74zPg0Rwf3/CRRsVOYC6tOme1OPFesN3Er+qr
44BD4LH55REBcq0omLgr1bkrDRrmp/SqQsEoM8Bw3SGJLJ1qQndd3BxDoQ3HTe3y
2FMPi6hUM8tv+MNGMQzR9/GDPTErlOfHShMFJPwahjULUXmRn/Eh/+J4dqKcug2t
bnUwqivax0eCRTBL11rqfftCJlRt7etbA589NmM1BEr6/30mI43l2UdS7HbaWo0e
rozENFh0C2LNHfVgG0A1QNKTTIzqjAkDGc16EVShFX550+rUaa/GOHnf9RjJOrB5
QXxv6+YfasNals2hE0PTewLvv7QViGyp6rPkeFq6MwPyxegAD/fbNAsKCAFtwYeE
wU+a/Apd0nzQ8dP/s5T4ObBI2N4uF/oukxBVyI+L6FA31QavHDfkgwmg7QVwQIlv
aVrF9pzQnPJpEqhEdYWhCsDh6HohQG8bm7Fpz+/qQDxmMcebYFWKNUFA4tKkPJgH
wMejBSmGPPgTyVu3ky4oPFBxb/VqXToIL4xgqnwuQf5kpZpbwUPaRPatZmyGjO1Z
fyU/cJZ9/1J7T0IyCQ/Hz8Hufu55a1RpbFjR0e2eE3gcVbhkCLKa9v0/jhxonsKR
jA9gcjP4qJef5wGzN+3WBrUxO+S5GpKuXxQ44835lmuBxOWwvsk7LzzWXRRkAyWE
OMFBHjI7OQsSRmRUisHxICcHPXB1FzyuYHXGPwyEoSbUSISsvpwoiX8QxFGGFKhI
ORh2scAh/ocyqCqqUCwhFsvuODRbM7OthhoEUNxzeKytUsV4eBwehc1c4t8ObmZl
0+0IyFN3LyREWcCoEfvHh5F3gNh35Pue57CmIMOmDbCz86f7FzF6BedLxAaFx6mH
BSCdDMF/dxkJM8o0bs1P2PhXXopD016342iizcqsXZ9mHFO3We6aePKHWIr/bnj8
dFmvR8X9Tu9I0UGf77sfi3qh+/2C8frDbQj4Ddi4w2JW+y1Cg2vYWZoaSUbyHSmt
req9PFH/ZHZslMEy2RPKx7BXJFh3WkDjsmEnrzJBufcA9ab494z6NRX7tNbNpg+y
peLX+NPIFun90XbGH3iMk8/CSHtF8wKLdsIlM79kYLLUSNNxvuQ+CbkuG+XGkpJb
buCm/Kh2mqzXcIU+dl5vLdm3cANPAhM3zOEomcNP6vlkKdvVA3sPSLhTBBTaUx12
jkOSgh9iAYETxC8rvVmDvEdaMnB7q/yixbZh6vt8Y7sYDwizdmgujJglOTqmUQt7
uNANQkFXO8w3SL/IOh5ygLfJ+TbErTs69oZFv97x1rl5LJwQ7Ir05ht7Per0l/Ly
Ke2QsEyQZJhJi7u9f8EVnbL6hqyZlSdm0pZnxog+ep5td3FbjOZEL7/9WGNDlfYU
8AT8Iks5IhfP4VpeZ21tBSyHNym7mmSaN6+kbGA4S0B3Kw2uAfcDRK3ZB6HXYAqr
Zgu3+151lEIHOloNF9vciXJSUSpjFbRgWJI8t56Z/HiNotUxVg9HfKQQenbRHO8l
/ATLQA2Y3ma4Lcxb81pMMiv90wAtALg3ghMDAfdcVDZtJkFrLRYdEegO7O5riMYr
uwwFGKrIv9xBjTcjzuvvO+2WGKXQgIOmpPn6GDb8BQzd+ZGetTPIcRgOuiTdgDZF
tiAlToCQfe+IyPxlYWH0eWFP3m3fR7z78llExenOZBJ3Geeyx+ifxMQd0SOdvhG8
uKn374F5/OgNRZu6zU5RPWpCCEMxTvTGlJOSUhxqiYnKoupXi+J27GJVrkEQ8koc
wzup4Cmd9OjRl2VwouMlxb6+OjRbd5VTYzdLaItmUmjyFhNdQEILFl51AZvQRo2v
abpO6Yw5lbcUBqFPbZN8S1Z9Y3t6ZdApOIjp926x0T/KBgb+EFjE0i0KtS1TLbes
J+SnhMkZLl30quRbBYbrQB7/l8docSkr9r6BUKA6fgwHvkbGccjUEHghYqbTr5+Q
cJizLuCv/PSKvymXxXSGrlr1wu4zgMPAO5Oqll5o9VRqU7OJkLlLUuF8bVLQGPQm
/91g60VdVVGlMDJHVlWSuWJdIsOc03mGtr3DEGHEyQNZvHNIpBpY08LUTqyR/5F8
EeD+tKi0NI40N0bA6N8hvBZ5g1zV6C4tWnLSOUUwNXiZi3Y0PI79g4GeKEmos4bk
wRoqOB7xOb8sh9fQ+8I6LD1IcdNWsOYuyh7pHuOKdf0V9MB/FUZ4s611zdAItPFZ
0XSYk8OycPfl46WxiOGTusSRDjMgO1AkFZXhXZX+6OCeJy5XyxacKriOqjX10l5d
RuJs4UuPeUooKDc85U/iq5US2UV0GGzHT/LvRnoOyaDAmEYZZuCR9UkPAB/8U/Ei
Q1QhviPG3M0GlLENYsPskLmeoD7krmb5IiBRU0Y+Snz32pSyzmSsWzNziuWh+YqX
qohTOhS3D62AZFDE6LFrAM2T0GUVwPoXCSA/sPu47hvVOj1YpmsJLCy21ueF/0R5
3o+X0/ZvvcNlcvyEDxbmPvGtvZVGnKVMTs3zKRxY4zb5cPk4E/tUPqSyRpBmDo7x
j8KsFUO4FzeBPBt0JeJ4SR+ob6v/l9yJ3Noq8kPPYYl0+OXkS98ou2hpjIPije43
3CGcFYUX1fgwsbcu2QGlgkD7F8ffoDb0pi81B94vq2lza4zig7xQf8m1aHPNh62K
e/31hf58vyk/EYHDvuMF7fRAdd5fUdQv/hXsnA5MBDy87/keI9q+QFT4O0oPus3Z
1YlFplFr9o4YRdIYy2tjvCwdMw/5YU+aPVjCYOAadP81yT4P9zNnTOsUtlKXl7dk
mh+jMgfJHEzLkLYbPfDv5PKp3aaNtTDMNeoNWqfG+Z7XWJEeqWh3ABKV4pzHc6tM
7n6OKFE0lvXASufJqK4Bl8966Tn8tEPDMGFS/x51YErk42zAjIHgegkKLF4KjE8h
H9kBnwQR3B9dZvs3bYkaLayZYNa63Q6tSlirtPetuYYNL+Q5+1HghpPAaKCQ6uhC
1pQlkmss6f4U9PDgaKTtrySyve6dnoxQgdG+H6h+QlKL6XSTZRPnWYkncW8d6VL6
z/a8h37OBhD1gD/c50/ngh3CrFM0Bp/4H45YJkaxtmiMhb0AKgJMo1eg//rhqnW/
LbCkbs7xcH+ERlp/X/dp1ODQA1H/ewruc8Y+mAhLlxSvIg1R7tj6EdOIDMHuf5mE
08pCa2hs9sR0fxTELyKLcKyEDhttK1X+cGAtCkVeiCfLQwG9V6TGr7AUWy3Pex0A
ZdGS/kYjC8TD8MwlVXHPi0RuFU8s2Yix2XeYePyhCFQNlQ8A8sTsYZBmF7Xrc2YP
HwR6qNwNQ2cs9vSdH1fCXzZIYX/8E1hJ5z51MFnEy13KWgDON7DeFtwGlPfY2JI/
2I1hel46nlgPOut5CjE+qP++QELj1cZSurtyBRpzHsLp3dOy/1H+jXM/lSoKbs9q
oSih4xKiEDC3Kc6MK95CA9kasdxxP3+uY2cY0sqWyrkoaV3oeJXkSHR5E+RGc6Vz
r6AOEWHA0M/wvlyOh1NHG/RVj4Mm0gEfvMK5cbtT2nDq45kvax2FGJXa5G+q6o0T
g4tbSsHQhPNVbpidl251vBg5wK75C8jVW/72ao8ne4Iuame89vFy/tiT76Rm721x
aoPIj8C8adRYr4qISwcKAIqSS+2qp32QmmQ56nIPid6MPPZL9C3t/Le1yU+L2kYa
sT6i9+nP5QPD+u2Dg8JLGv5tQmegSFJIyVryqbXwVsA80BuPczVcMMEstRVs9SVT
gph5Cx4/RA9ARpLdkepf5CD1zMq0cFHtafZYYZG8Djj0fZ/qrbCF/PMfSJcqXGez
QPYA1LE3FPaaC0LYthYNTkjVhU4AvOTP0GmuuoPQ9NYcSWxkmK3pBUm8rNOLD70O
SCq01vA8MXa5qI3VXF1OJYZzFoDWbh3NClVSYWN+L83y9X0zeSox0H5wo187DUxU
/hHmCKbVyG3GNIVsoMwujPhBYro7IDD2DqR8i65POERE1bdzGm99Szc0d91Rdqym
kyV5E9l71OwoaqRTWN3fTScGVrnSwGDSUBYSID9bRd3PQtZhY0fkF12bMenevWiA
duIjwlLj18uHsPSeI+gmL7/7dV8Uhw1gMShLo6I6kRIEN61oPdJGl5PsM8E5hPnT
NHmypxlaxbp70EX4b8JkmS068D3VmO2nm5KfOdLpkDMwcCnt3RGtwjouDNTtnG/O
WRBWnHbrUWZPbnpFNIerq6zpLRHKRVQ0LZR+ULENY/LW49JmLnzVQHSdwf5JmRIs
yglRBD4LN616aGx90Tqdoc3Q6qHC+G6MfLIKJrZdzpmAlHIY7ctGtujjNm4zXzVQ
/EvaS9a/jFZMWKdobGeVk+YarevRrj51dZFNRA52sGOjE6CmZWjDcQhMiXLjSn5g
Q5YPhh2d4K1jWs0jAPt0hl3ljzDXRAlvdH4yWyRPf6+GywPmvWqub/wWr7uCLVCu
dV6YsCySjP+tYpinICdU6Lpxzm8jkALg3cBOHl/uwxigC6DyIhFd1duYrqvnbNbE
l2z201rmNDun5KdsGgV123uLlonEZcz3Jw01jY/20c3e92hzRTCfDfR4nCGC7QTF
Yl6UBf0fd3Fz3S6FWExc9vRgI5GUc6BsMWpjICHP5DKQpQlrjLJBWy7TNg/k+61g
keQzBrJcGHAY5qfPBLDdDXmnl6xIWHbVp8iJVzZGwn6k7lWcQajiR8WE73FGXJXf
tUM7mR+eIDtJ3w3NT9lWMPE8mybgPomC9xWg9QJ6wXx2rMpoTcVGhmHdsbRmIqZ4
oSV7j9JLQxMYkdpMYcZYHfFW8TN3R/X9pcmUAoA50Qysp14N2r2xirGuwROW/UFD
R0EzculZMe6nN5VvNPUZzyuvPsEYhSafZVKeGDZ13VBpHjHgPjVexaGS/JbkNRut
1ctvqoq2q3VnM5KZchE6QHhcJk0GtqkgCeo4EjlH+cT++GWXdMpdGEj2lweexAlL
7rHabW/clisZJty99EPd0gaVZ1uASPO3eHPwEcyjF+hR8YgZlIvPWTHte2PhdxPn
oJCLBmhGKqyZ16MHureDPmziZel9+JJ7SVVeVKxk1J3s+Wb5UWROMxM9u4AcfE7r
JUbvM+xT8dbAYTGt2EF22eRKwV74HmD3WdeJkEV6MdzgYMeMJEaP1YnPuQfzigqj
Wi4QKkzw7NBmdofdVt7LRJsCRe7VNhq/nRBSd7mOHigB9JQAwYAkjWvmlpafyPQq
dEzkD49lt1fl9We0m0vxeU/+5FxJmaSzzgfuEsd0JDLEyIDp4aEhp5st0V54NTWb
7S5X48NNF8CFqx5yXjnLImFcYzaFB9IH3WPS+49BLSNhkyulO/wn8lY8J3Z3PU47
E7L2ol3q5JX6SAiCMKdbOiiQI3Ke2K0YHWaAm/aDH57BVuSs5TPUufzkvjCG5muC
Frs5VgaTsV4Ytkx9VkpMtygvv48SS00hihf5Ez2JvZrMAF228RzxDO2M3b+lWBY8
v6ce1+sVZzBNaDxcwxQCw+FFXfkq7e9TKY2jwHupppGmI1JufPPtn9vUUPN9YHlv
lwP3n0dAUe5y+l2WkZKQyUDiqViArjGyz3UL6pbv3kfWEOd9+JK2fKWRD9U+yFoK
tYHAdSS43T/dJDM9fcIOiaz1P837kCjQ4huIooSiGCE1N2h3HQyv/jZEzED6S//g
on/O+GXc9VhA/niAcOnUugbq0/rTKi6PNFBlZG0DzdKOlNX4FOiCJKxQHGHNNvVR
RxrJ++p5q6vKXNkE/XLftVSHei7rKdpaxwvY50NSw/w+hQCK3ekuOwETakknUD3i
777ulSpuvGkGFPJTzm3s3q277QmRx624dKXNeu0ZuJb0v5QQt2AWDCE6yVRjo/Fm
o/tno+AD9KLad4/9A/waGV7b9XiN03jG7qNFtEOn34bXjrrX8B98Zj93RxyovLFD
7CdiQcqpbqB8Zlq7YM5+v+8P7M2JADlKAsJ/FLMmGIGxoD0J9CFV0q8B0XuLbDmS
gGUL8E98pnIGeGZv1FcXvsuzhOtCqgVcGi7xRC1ut3FBdsWL+wjrz1+gHV42MSqV
+rJE4E7//vQFkn1zQXBvAiQ5tt67SEQ0Y7tfbedzzpd/qngf2XmCZIv2PvrbdGXk
IxjPieIq5v9QBhwNEtM2Q4DsWsuKYd2I9FuRXCaQtbM3VOGkrSylR79IPUQJWew8
KUxObcrT87btGP1AfkRlJ3xwd66eTLOk99dCEBNt4DFlejfZ6nXsuo27mHoLIjOC
Ler2nE0MiYA63ZHMdhRKyHvihmSC53fCL+8N+6Exg5vVqgV/7L5+w+JFhec/NKqO
8wPlDYZBSSH900p8gjM8bAdt1p5ii1scFBU9tBBmU5rGxmbkfc6WoACUbZO9i5Kh
CjzFif/ipLoj3EN1/tfwJbto1Jq3gwMiLJMh/6iNEs0P90bDLHbdzX1uA0l3UQm9
bjx7LW5aS3wV/Xn/g+g/ZhAHe29xgnDVJLKn1pyVQ1WG3nT/tBcTyOgbNz8nbfjj
iq9YI8rLvAiS6WLwCRVVdvkCf7WoJOh5dUMALv3pkmJGPavtbuDv5TeBCWSJhN3b
4YksGDyb9WBpw51GzpjochhTMub87jZ1cSb1FiCLH8pvAiKCUuJ8yD5fCLzqLU9X
TXl8czNLPk1CGmImgqEP+X9O6nMK6LxEGspeS6pYACjZAlRXveT2SxV0P0RTej5P
JEoWXDWtE6aaj/UYDTzAW8/JOJ2KDqJkPa2XAuK7XZwXxIFsZmZKkFAWe6V2ZpaY
r2YDXDiCx2LgYSr0goxltJHyKXFvcu8oLcI5C1EDw+XSZqb9Lx25IdTLwm5yhADx
66eR6ABzet/PspePZK11d9OZSfTsiVIZAZLnqERS6N5F1GzcMTrr22CE3LtZ/4KC
XlcXigZ6oA4EpjET0Jyc4B6Re7JJT8378HPfcdAuyaqK5uTVsOsue/F8V36yhhdc
rRpneQuQ/TkQJU59DUqN8209jNJixcCQ0guPoF2wWTMG3goVzyQGRdY5mZaAqcBg
hx+yqAu+vtNNfXAIFB5kyidqI/MVNk39vCn64pctLv3UTAqbbuUWkIVFMyEn+2cF
q5HgIZpbiexFRxdxFtsXQ6k9MmF2rzjhGYVPralF8AHdJozgvpaE5gUhd9x+2dK1
kdOTydD7BRsFnlsKDByKcs1V93M1y+a4NmIj0EUjDXnOtf3bw+mt5GwMmZTisAMn
1WNlz3akdPHEAyx8HioUGHU8koiE+C3PSeIHofIvl7yIl79Ajv6c41+/L5udeDGU
stXocnq3So+sxFGVLRpxodDymVruD1vb1dMAE8f0J+FTSaLAUcTUHTVQtA/xhd+G
zA/ceK8dZA9QuzEo96tl3KUnk5okJk4gD6zqiSo5wmdshE/Q6snoY5YaLpD+B7SE
YUyFaeKPdI7p1RnWHQo/0hHQWUpnsOmrXMYSkdvnDR/7oPBWHOnBWe/qpsL0pRbv
DjZxwePQdO30FihwdCUqxyJUki7eHK6zN80XW4Wtt3O7Wj8PZ46ZzDgFqs+SP9VS
Wmq1a2QesMwEYVw/k+gOqXlVPes1ODrypJXhwlt2y0RNqoStYN8LBmCJrU4aTrw9
51XE9c0v1BecEwqijgQbafTza2qvSOnck4ViNy7FiYEerLwllNfKR7Jo7oKtkSnl
kG86wj5ccd3SQZhRc/gY1yYNZSM+FChikjeSSdqLpUQ3gxfHkIP/DYQU+OktXeS7
XXyzzHgvs6LV+9niZ1EiXSuUJWLS9jZf0BCRRKBINgfq16fQO5VFgHx8r4ee3BYn
MP9xGL5qMPduch/VTuaff/Zte7nVGublCHiY1T14hdKM0aABJKRIpvYKKT9JieFy
dFl147nxP8YygY6od1yfLmBpCZer0ZdZN4oq1LPtDl1SKVGhvWJXo+bRZ2rQ7nb4
Pj5lCTiAeBPF7UjplmBkl+W/ukDohLEb6Ryw1+4zpSlu+3yInAozwygKiltj9D0o
VGEF7R/Q3qNGdx+u1xHCrGlqPiJyWAhvsUmiDbMX+Nc16syKT8KdEfupHTDaMlHb
5SbzKNMoQoKy8Vp3DQ5RxR0leX8V/Q77wZ82StG/DXf8wBErKxekcdLQ0/tk/GZd
p96lYQahVu8qZ6EKHxIIwtPlF9WFbYNOUtaKoNg2DYEjrSWmBVkW/5W1MhNfCDym
2nuzCtllC3Ypa5/yH5p2cVvBkLVtF2nT5+MpRTTg4UESuTgEZP/LYNWgg8AkIHE4
LQIQG3vqVfVmCb6B7S9kub/Beu6NasXvhedig9BV9DBhMIGp0KG+tZ8Zzyx3ALbi
CKXGQvuAwpWLAYvYEquaE15ZVvzEJI2GjHhmbeSb0leruSNCNw6UIDG+keS3qCzT
ejcjbQtcsbcb/ThHU6+yFHlAEYNTUzVT5xSoobVcCEzuIxOgjtA7KxUatVLmlmRP
irHDDmxLGgF4FtI6euvCG9rzBp0jL6OPLZe7xPMA5oRBOfoO476UP66+bLRQCmwi
yAW6e8txmkDYJmhM1EBkzqjgT6o+w9FjiVNIyZaw5ylrXydubjcTgUg4bVBJgxPr
zdpi4iKuiy+LAR5NQlfmYcOgHRFFcNBF389KdsKXaB61H4pvvUXs8GDUlv3qinHt
EJHDHc0xKMOkg5A0alX8o4fBb/ACxxWnZVNZtHVaikyO7lQQ7qM+zcyyzMJz1RJ0
JI+IMQYTN7/TH7tauVkvahPfeNAcEJkMgUTuioZGoax/BX3lPXAz/1BYfVCfe7CP
p95eV2SitKhSyNWa9gyCUjmUaYn2jByP2CwhzAg/DQT/yc0kvZpB2cdyYkFe72ZA
nBgX9Z/WCCdhi59idPfWkUcU4oJIHxR1oX+vdAZCI8DOp3xaDnaFyAeVJWvhBR47
dJyFLOQrS24vbLd7IR95GGKRFebEWbbkQGCMZVXFsxlran5vSbHfxUHSwh5cGXB5
3OEvq53TBMLn3FGnjbr3Al0iL1pwH7u1Ywj3qQBEH6gAqDeZ4yzL15bfjlUS+O+k
YFAh8WekhitjLBUj0IyDrqM6n9tlVoR4iIKwWjn+iJEpk1wtmqfJiHfINWEBWTSR
p66pXO58wypfMx+5zyBu4sRwNubRgmbldexhP7vY16pV/KOP+yMIbSv1PNtOb6cz
DHSJtucZgTGMZAakU8RJukIQH/IGrrauKpDU9GRy+aaVU4n0W7Uv/wYGaG3NdkiI
Z4YqN1O8IZqvBTBAPhV67rqky5pvk95zLHduXclz3CXm02X5Eo2pCPtF9x37NiMd
qdjCeX+30ukF2avS9gGOX/tBEupWlCDGiD0Hx49qV95Ef5xIWOms5ivx27VAx9Zn
w+Y3/WPJ6zfJ111EicUoGYHdjKghvzFb0FsoGCO9Xn9U6nglFykVymChsALLFGkh
iLa/cLWjmHt0fMqx9IJFDHuLk6QFx3VxNYV0u85FuIechy2lVb2zbsQpeYgZ51RT
R02GL0gzRs5RAa580cO1envxm+ILW12SzR8CBQgt34Ik1P/2DyJEtCwbancvK1K8
b0LWLZCcdvEhutRmgV1mgYgbqBeJVlY2y6IpnK2yDDlSrcVy8ICJFWPMMVRhgl0p
9A4+REPyMjZEie3oy5nG7tAIQ0SKb5q662L4mvIarwpJw8U0OKzZCg+nDmauvjps
Khk4dQY5ksAwj4ByKCte9EZ6Cuvhj7etwsnEhmjFwJfV8Kx7eg8APBGvS7kmC2Sn
bDxiqthpyggKSIZqheXcav7LADrWVbK4g//zAinDDXW4Dkskle8pGQBLogBzHtth
5AiIK/+IEpIzpdzLVLvGZXnGFfI2Ligu2TWNcwTavWM/GbpuCSXaVjBRLglDDYzK
3xaKmvy56Y6I540f/AKAizq/AYIMqKb50wlNEp2WiapRdVsNAP+DFLTYWFAgfwx2
gM7TDZh5wGCZuKdaSOXbdiLbMsV2SpxkE6gCmhzTXuzvcBMwFbZR+GIEllm8m7GS
Bbxw97XpFMi5nHgNQAzCxe9jtfb1X7/WJ8ep7J/usHsM09KZcVTgC1au+jUvWEca
2O7+qbMIb2nZGglzIbiF6nit3CMyHhVNvA4Qnwjy7kHBIsilSBv3qnmOsQnTCyvt
ABVOMh6nf0Fo+xzHRh01y7UFksroyP3drmzppcVRX9wEL9GlLWC5bsDEnoH4/QNl
fcOsi+xjjwMCWC+8keGFd+0LDxtnESMq5lgvLyvDLbefEkBYHFrSEOemav6aBuYA
U2Fh86HyUCWEfJZD4zBfOOeSgVGOJdwRZpQ44Al85JAN/+RXMoKvnlXDKx/RmMh4
QGpOrR4drrU1D67uukj0NH2SSS2q4VF5F3Je1pEgVUnFph5q1r/N+Ehmc+8LR1hx
T20bLneHPH/OweZXJ0HwGBMTfabZbZ97sF6w2K7lrT5x/H6reO9DsXam3oMAh0k2
KA5PkRcLp+oeUMJNLbKZyNnvI0aaewYtuvwPH0Uppt7xg245joj+ESehivawEFd2
ZkFT+0Q/zSC9CFmJao0frkFQTO68fZQ66E9uTCDc6TCWg55lA3DwQRMgtjHi62dv
igVhcwjMzvoIbq6gkF9N6vo2u5o5F51Dwrp+JQgD8cPWkajy57X/K5bW/UMye7kc
xQvtYK0aliKezgyO6v08uBEdp4DQtH4RLKa5klWzcnT3tQigkcRnXfToz6FxEHlp
Lnw3f4KHApo/fND7YquGu4rQbQmdts07z/A+YJBpUtBzq69hfEikpncrxviwe7V8
NEi1NxqZIPhRBz5Spnkqjs8QvP62EKDzPbP0of1ugmnWDAQQjhaaWtopDD5ggzBv
1atqcteJuub3kQnTg159swt6vsLkbhJzha0LqWobIWM=
`pragma protect end_protected
