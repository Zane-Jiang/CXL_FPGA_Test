// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NV2UPxcP8Y3CN9/q6JB4waVv7DEtJ2ucKS9KxfQZAfT6ov/1lJfz7bxG/q92
VxxdiuUthfkVA85A/XYQyJF+ZivPHYgVtgtkSPNKz99icghHS2qspzXnvwGR
eNlL4PmqXJ0d8PfMx7t1JOAuDAf44VmWP0siQWX8fITXLJfLbqnOMqF8k6Ax
m75uww/UmqV0U9GxTw3m0pURQnvqWc49rjtvxGH68oq5bHcv0I3h89d+1BaK
purr1B14Akqh+yVpPIRKgwCu0V1WRPBBXc5Q/DHNjblLDiU39M+fiIUMYGGw
q2gPSfDeaU5FuUO5Ip5MauGZxQoTBFaQsN02/mav5g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NJhx5YmA0yatfdJXRQP9nqqbdumexcQk5SXFD+qa54tEhoc1kIPzn+/9kbxt
Lm0y0FfXZPSDhDu93GrYaq4eZyILGiNKZqH8ZqIb2sAD13am3EnZcGKG3eBw
zCJ5Arl2jgTQqItwXjZ8qg/T/ukLNOVEYyzHZ0bTMnYqNDqrSZ4SPsKfv7X2
prUaV6FhRObfg3vHsMMqQa+kjfSJ0CWIv1DsOYCVJ00bN+7SSIPuAbTPJw9E
alD6uKJ2TLJcruA5StpszI8YjRRt+pmM06iaukLugevbsM2yvoOqIY9URX/h
mXZ8LNLZlWDpN6tEf15s/DHpnXuR25RfY1PO36sSog==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dtf5lO32a2Y0A1mc/UIoujKUOFUnLfvRXUhZXWq/c6wAkRwPgjMcgxm8TNdo
G4l4SHSK5vXcgMD1Z5NATWBIrK2faBOgpjWPSL/Wa1WejQzSpl8GK5Hi7Byu
UgNBw3xQpgmLWAHO/TXSSh/XmvL7wGC4C57TyOKbaf+LNi9h8SeUyXNRSBhx
FqP9a5Wp7VvW0OGbRc0+zHTVa47gRTPllhJDFbnS3DkjL6rZXHArJoYTLE4H
0b72VC10UgI6F+gh/ETq/38rAopVYG6MQJOwb1j4Vv4LMVcHQl0e5BdM6Shu
EqMqgup70KsMsw9RBnpvSRqzPYfEZytWrQ/MNFiedQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lDaNurvXrwpv2uWDg0fl83l9ApkQdcCnU7eJYUMR4z2YSMlKrTNGPOm5ls0z
CTR6q0lUrWcJX/8FPnX/w56N6YpvsaVQQLt4a699zWIxMDfrRZTOZhfn/eHd
0oqjSV+VeYla2+UGyQtLJJQBP6/m8V+EQFP9LhpbqOkqcsASQLA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
n7YJV7FHypWp/2WqUiodytAaHXANsdL5PIHsasZgQgUBe40BA5bByzp1y342
yg/nzs0qr1zfuKskALuWJsVfZyUeK6mckNYi8OvwaRuvFuzlnJFDV9Pm5kwg
ILzn8e6QG4c9JELKzQujIy8hMChxZhRXpHw06n2KvQjt4NWGtu51v/PNZnWW
gAsuYk3Pu1o3KP0iwMa0DqM6AbDn/iQmQ2L7D9Dq0IfxSa0eko0XysFFta+C
g6fQ1P8sf5+8RfoTUGRRHYsvhfq+tjynyvdVV7r4zKdW0ZZQ96eMyYsObzYc
oQ7jQudtnovfuQB7wikVvrJSdE3crpPTOa5UAp6q5mGYbA1hgt2t1fFIkMGf
8DSR8SaJho0499C3VBbKKerEO3UpqWvoJfyZ1U5b8S8UWnCM8GCpxp+nlQa1
9JIkUmz+xj7Mnrblseb7bUvE1pUu6h9Gyh1vm5bVYdF7oA2HLIDZbQCeygeW
I9QMBr+kOT/uwbl0/aiCYnJwpq9VnOgo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oHTc2z1Erj7p3br+vFhxmM9CMOH6GmIq+dXU8B8I4o4/uFTRHweLYrfFstnr
UAW1gPmKYXcyrJS4lcyeVIWP2geAefNyD7fq0F3W8qPleM+WbA/E4lJEuRI2
mXytL5Tv0z3ZkD8mXITJlRKgiFS4EljNa0/yJnuXR9RHA53udAE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jeEZkG50jwoP3MHikEQkfeKFtOcq4MF+m26tkLta6/ykv3Ymro2sXc7mmuLG
2WKosk1wMiwDx37nKpjnlLIUoZZqjxSEnAAz8f41twplgRlbHdyej2ewLpYm
tIdf/Shwq2hEPUkeN4eCcW5kq/p1VkL5zSM6nyI6hm8XsTDmTKs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11488)
`pragma protect data_block
S2kJeSZhUiqF12MAbGngPraDENnM2TfimuVrY0gSgiFfpCuFUtg0GGPRvQwP
3UEQzpqSYHtr4l+mL02BBkycx+ZjDTloizxhsONmFZNN1hex8MPGoHt+uoCT
Ziyj8mRr03T+/XOAtlcNFsNxvGc2LpLRBeNGpOvIE3uzVdPSAyzicbiCoXYg
G1949hS270lIzJM6GHgZIZxi6FwBduh6t5dLXrwzKj7nSlbi/kOmugaZQmU9
IPicCDQSFP93Y5FkIp/L2EzTuKnJRUvNvdKaePhUwbEad6UXXT3SzpmgEjts
46DBOnlKm1a0kQg8GWduQf/8aOkjAVBr+8odDT6GKguZLJyLP3UdsV6WYoko
+IygdWO44/Dq4HW58drzj9uegZGCO3LGtoL2phAE/wH+pXpI4jypShtfLiPM
KFK6gbmWLkZ5ypxr1Fy3qjVy30mJUWz/+4nl7iY13B3sLTSLUkfMiuKKYySX
EElN2b0j951raY79ch4npGGIvqYcu/p7y7ZCLrXrYHFtggkzPyfdiIyAp9FB
6O6YmPLDHWwejJ3Gfo6jZBNYxkl3vsKsrROAIKK1UIPfgE/vCVrSzUQfovM6
FSQD8d7gO5AKGUXZAMnnFOdOkYPrkgepX8+MTeQlbKKUzYdQNRiEIgf6Gofn
ocSWe39cSeM0a6VQKuNg1xXxWIXUa3pvvru6/7PuD+a90wHei/soojj0S02r
SAc+/q9EEtEhFMkLYJlzNbR8DGb6ZK8UPFH+Vbl/XKhkZ/n6neuGy7cfuAVr
JHMPEMgOLMqfejCtfkJALPi5As8ocSbVnJMKruqWOWAJIMgBiCngRzNs2wO/
QhSHZd8xqoh027920xqS2EKjFZi3G8kuMyIU68kDGxHAixxy+GtbaHODclKE
yRXktW0agWejFlQuA4LeC3HT7GqkNtDxzeqHtlOSxYaBr+uFOj+oPkbxQv0j
axZZ+MdT/AF82zgVWRPVO9ZMhL8wvq/gdZY42/Cp0ZlGAzX6QQ1aG0ftu61R
fXlhDtmAFk9y8tW/ZQFgYd0xuAQVqpFrDtUQhs67aUHGfiGGnXSgFBQtD5Qx
DkG33bcepWP1ur5pRgPuy38EzDd1EobG+vvQT2YYCCMTD58Qlqi2t+J8PsZ1
NjhO2/WQv84TG87VVcq8mtSVyxA+AYhj5zK3Bv1q8T2/hJEwGAtFXnWHYQ1d
YE8HSoVtNs7Why3W1KbSAL4WGt/aClgYDv3K6+1K2du1r4SloU4HSEMax7Al
YnriZI0O93c7obBOPwiaPFomxRUPoXGc1eT46/d8UmAzy5h+c5UCeoKyjCzM
d3iBseWCvHNjG1iw2vNUNXnQtKxp6YUDir+YkiDS2bxhu/ZQiyyYxeXR+kgO
BlHmLX+yPu4Wme2iIdhS2JS2MeE4khz3hHrwXdYrINTLQNSc273i9WbBG5KT
NswdC13Qn3VqbGMsrRdlQHuqYI8C4iY+rL8tdPqSEDTJPoa6+trcPLc8AxDt
n0VId/oxCpTVt7RDFD6ohJQrBKWJrrpujTfyXJREGHUHv1dUg95fW++IOVrn
iIYvNryqJpnuD7oJgI0W1rF+711VYiFA9PyxpPEl5XB3YkTssQwJSRPB6IDg
25m/6Pa4Cv9pWA3MYF5qSjqvwBHj8sP8PklPNT+bUAmUF4XToOqH6iVZ+cUU
wY6G9eOhSe+KaclTI1MBrZI6yEWHLJ6BJ4Ehlw4q1+UyMl2d4QYoEWuiiTfj
W7iTBGCcTod7xUigdeYsO1XOB7KWz/akaHAa63o0Rd+rVLiXxP9pzpXbZK65
asSPXsfThtAuvepfmz82uZMkjsF3t4cAE8w6wLCjKyfyswEE+ZA6syAnzVYC
21pxpqB1HOrXp4gEg7OGDZ4sctufgqwNL1BlWevFA7rxl9HHunenRFficU2+
XvaVjifg4rjtC5A04JG67oZGN4ypD2cOorgEptElSUZtJcm5IRi6gJ8igqf7
aKwzz7xLizXhCYO7ds84MQzxvd9zFVnW98HHhUGiUBztFdDbLYksIOEn7Qnt
JjMmUGNYjL6zZn9c91XH502Uk/mxnThQcmIxNJ2Gvcqm6KAweSRoBRTxIdnO
XEA1W52+pK9dbnl0aIJYlvtUFNDPqoGyfukhJKg91IdIqKPS2myznwT26D91
6i1mo41wSe0SquH7E93IJU6xwsNk2LTj1eUOOAnnl7udRmhPT94QUambcG6a
YOtr3+hnaQmNmUC8hNhh70wRuTVWpups1iaJnK96UjhlPp3Dfb9b/dORbtOg
Fm3GYd9Gt7ziDnIaH1uaCTWGtU8sCMUgkaPXdV03PnraSsrrr2hppJ0beLGa
LP7T/qEb8PEEFwPw9fjYJr2OoKZtOvL4J5BDfjKBgqIB74dMjh3pZ0tUT67N
Pfeo5ZxFfv4J8Mh/SXvXVjbUPLaAkbkdf1HVrqKbxvRbizsdSn809j0x9+E1
1qwBbYvpMed73tc792hwOaTo3zRdGlv8N/rlxTGYi6gkReefFNZbianutJ73
M4uLmupE5rFhJqseELsn/Jqppm1NJCQ153nGQyOuBMEmTt3sxH/wvMm2/t2T
LLnD+auauJPvZA50YZUjQO9EaES//cGS8G2JWA9bD5SrdSL3Q4AH+OSmeKIh
O9QeiGgW3ePjTS852qB4C/EDyZIM2TPXeoZg9HL3CJgI1yI8cKUYC9NbQ43a
e0UbtrcytpqsaHFLQvs7mk1njVUXAnbJRo4MmvfwErbQMbKPpRi6nIzfGLUR
JexiJLBHXAI/mWeIk4Ia4QE1LQmQGLcVt8JuL71lQ9MoXetoP50WIG40+yUq
NyEZimyIbZX4FtRti0/0oX8deM6vXDU+M5fAqlojVaMm8nbqXCQkShEMlH52
l9R0duAHNMDybU7mugzeN+y3pegXlblqIs0ZtYo25HiDosSIROTHOHJORU8d
MWGp7cJ6X8ZJTlLWkufO1syBwrHxSvtxfyMMn8JfTdImfksQ7INF8RPgmu3e
ShDzLeVhqqT5AfuYvjeKrrPGn74SllAuJXTtSY0XRR4kGaFFcNrMGiPPG82E
OzDW5SUFvb3oisZwkmSeulqWAg7t/tX7VwZqcYTvDt+8uurctM/iPumN10QX
+17cuwlnMZuK/7yxHKsSVOq6lcOm+Qn8c1K1fLu6stntZskxCCVNJKT1Hyrx
n8K0hjApQVQNoujqiOko+BBOqgEwS/yblqAKUjwG6C3gFr1edfazTglAAQB/
6xmXnB22NhVji2UN0sxGvpYSiXq0FZ8JGpS+H8foZBlspFrpJYwTITIohKGz
G64YK3PYR2LzwfpInS7U18aSXV/5+7tpDijlQgD1y1yNn4R9BGYYcL4IacXq
YEC1U3gKOLtc1KLMM+xhMkELPv/fhoO1vpD2v7pk4rLDEr4MdnF9ZJH3jG4b
F2FJwOlgoJhuuJjB5SrIgkbYmcFs/hgZuZcBo3y4CoHFvs7iDV5tLXQeC0o4
BTKoaRmdhiJilAClDGUzvm64cptbJCiKuSwdv0oj7m5QV0ZVMAqZIi1FV0+9
Mx8/y0bAqEvE8Jn/s/Z6oIhNC8WLhQmKSJ6kVe10gc/FMUn52hvIzKH6JQA/
qwUwnutaKgmNJqPr8ijNQ55FEZIXShsNwkDW3031ehqglhekOJe1kdDu0q6j
z2FFIcWUWmeYAgIoGAt5N/bDpXzKCWoeiFnMkpe+6BxNAv/S9u1BPnjzcFkm
d1NDNsJTzybQgGKE7l8dIxlxCrIBZ69GBU8Hz9Ff7A0tVP+1/chbmkwyB082
Eh/L7skbxFn07h8z8WAITchHWFYefntNmHjWWh3YlIiCmA2ieC3B3IIBsinR
dm34tyrALFJQYo3TzeunjZid9YpbEE03uTs8wmuxeCpq5ZlVZAN8CJnyLJzX
7f+QTsk3Ufy2U7jbIJwGMTzDSTOm1+NcCkg+Kix5oa6zMbyclqz5DV7HVtEO
9domCRu6vg5+BXAUKPqAWeZT6jpZfZ5UI1RcM+2ZaYhypCAz09AzEWrXuBXD
J3f8P7hYE0It/EdPxDv+2V7zuo+It4XFOtnXP+0XzQJkYDdg/1jMeeUAfv/5
FSqxTBU29fz0yVpxRZZoC0ro7d8UpFrdzIOylkd+sFo4eH7xMC/V+FdqO9hz
be1ZQ0UlIEdR2cyd5gm31x89DHJV+DK+khWcypLomOxslnoLNORHTpChEjNL
dLGz2zs2bDzYowpWu69l9SLdBqHtHu9OZ9F7GJdDTdcVNn5P+lc07+rM4MQq
386TA3voeudL3gnUQWDiJcMoXF6AQStTJOd4/xuOgWq6Ee7sYhQV1Ss8aOU2
JNfPWF671ogAxsTh9Jw4JLoytQ3SfsnNTwB5LeAhiYHQAHWhr55+Za1Sevo5
WuQA/YSt9Wgqls3GgR9GSTwGVWunp56TvU1IX6n9u6qsZhC6uR1MSxuZt8wi
H5e7TZEdOh7eDV+qJ36XH8RXLXn7tmxnQiYaL3gdIcWtGNib/OTjfKwJ+VsW
Mkk1Z/ftGyBrgor3KcP2pacRpBkt6Y7uWD2/Bm3l/rAfoFVNsUiW0j79jiHM
HGcAikx9zl5LqvcQZU1IeiBJeWWRSotC1sSkPi31lvG6HQG5UmUzWHcnZkKj
MB+w8uwrtJPfwtwajH8P9m0KlC863oxCednW0B26odqDs/rF8b2Xl6Z56aIO
IxNeI5cPYFutE1Bv20kBzHXx+AbkmKdQn76GjzHk9rEopoX+YB3xWnHWojCX
vbeAnsKevO+5+F1ehqRq9E8WlXtRo9lLyg1qDbGdEjmWWWBDC4y6wYiUsr5v
CGyFCw5QtnI9R+nGd5DNT6TMFdupOgi3PqLgMQ3egqskQD6FZkVKyWOU3aMp
6exzbjXyaKRiln8mDc0eipZvr65NnlQsB4j8EzKy8cmIwlXmS+kv6oQjwmMu
dbBPjDa5tI89lVENk9h17LUR+6a3UqXrBe534x6Z9+eouNwfUjZD8Ar50npo
PjjjQOX7AUuxs5aiMfTfXlIXOg+c7wRaHLpvWLsHJNP8etTYWQIsLa3AYEp+
PldAtS6aaGkqZOuAzt0Y7dIZcgrPciWorgxPhb2jdJcYYTLwMOXbqUuBmbed
UM8bbE2RUxTyEJJinAvdIIx8X7ZbuovocriqUavxD5oc5AQL7jOFoVNdgzpg
fpYPehbabADtQ8M6iHzPfNeEfn7jdIlX7vxXjRWRoXaIjEC9yUb1SwxovGcJ
Pee+awA76Z1iCIZ5oK9Ebq8eeymnzFgMEA6haHw/Q6OPP5UKdkGvMj0SzQi7
7Q4+fTb2i9G98/2mHcW4bN2khC/Tp5L2AdOd8JmJQuRRf6+dCiXrgorOsEND
SXtIuiGlrK84pWU+E64j7ltiJ2R4ZDyZ42x1GTxZZyPBrHFsXyQbRb3WFRVx
07sCMCxTqbHRiAMgnZstrPCss18xGP9N6lIcYnLfC55PutGjTwb8BP531xoH
Gr1+OfrfmYafFj6YHyMvGzWvI81EIS12KxWsdJQl7djGE7s62ms+XYCn58Ea
6BfS2067pmakZfwqRvXv1zOkPR5C0PsDTj0xxI1X/0IERXM1zMgeqs7UFxq/
iJyJ4dIZZxrPNcpwIxsm83j5gq5xCl9aN4v6TmDo4nw4CxAXnjyCQYCGCUVy
UsUfXqjh6YxgcNCcBLHzBhv/VsP5pJdC0Otb+HIT4mIRktESZdTuD5z7/aHV
PegE/s4wINw2q/4ytWF0BLf0RgKGR9bNTs/KcG9wwuutwHCDFTxlv2gSJZgx
HgV9oObJcuwEIze9V/a7OIXprytS2PxLDThU4wAJU7rmG8PjhQKkG4d6ehmu
zSyqTcnVUZnTeHyapc5SXd30059SdOdh8HHxkw5Y5Tnof5RXcRCnPnUbfDkB
XJ+V1kyaPSjtYUkfX4gAHY2+qfiFOb9ZIGjQA78fZ0+fvcgQfo6ZY5vZhcIw
c1rHap/QbKwmDjK5tj3kX79wxHF8Bk0csF4B5uo0A1Yk5Q2kHHge7B0yc6hF
olUoxNT+91WdOyp4e4gvPWXGlwvPXHHGv3YddlZcq21V7YUi2YalU643AOFC
SvdtqHvU+4uTIZut67jbQEnvOPo4K3UrdL9MkExoiLr1/Nco1BDC89UmNMI0
bntYasvLM57ruck6S/HJ1Y7zs366vDV16dM9TDWWPLz5DKVX4WAhHqLdvwyD
x4LKf1SvPGzspIdsmOvwgj5dAoFtEcEwFyVPbbOobmIqxBun49s9UEAZ1z5E
sEi7VPRdtPhIJo8tBstWCULvuWT6TgOw62rdo+jkYm3yN6wqkckXxSOs1CVw
OmAiN4WD8vX9mSuh6F5+bCeExJ97JomQgXYX9FhMaIQO9M8+gJrKVFfgSboU
ImqComauyppgw4hv1IQBNZcWUo8qvFAj8GW2Ugv0PVn1MtUjlV8JCgOXT+XJ
Rvcga0+51R7rTAdpBYnY8YpKqBc+d1d0q/DBARU/9rXoXkSeKzhB1+Aoc6Vw
+jLUQOWrdNvaQgd3jJV4biIlf3gcBXQdj7iYjtCEhH0eBJAv2tgdpcgd9wFx
+omnLAJGuQeNMKxKNWifdWRyFsET7ts0PTA//xXTo+/qg5GneiBGVK+CJDOu
SnwIMPotfLO45mQafE2mmeICaowegjTK5wRadn8tWkt0zJNwyGwIVbC1DKtp
jAhy0voyrGQkf2CJYFErt37r3n+5ndlDvUZZPGseWxDUPOJmp/YKYF87wmO1
uAWKTiUvY/zL0tWGK+qB97xar/Dxz31/j+jkoxOviXqN+l7YK95Iya7UrmAC
4nj7D3IxdKl54OrYpMT/rui3B7zl8pvVnMHPEwPp7FOqdOrlXTSnteEVNWXJ
wH6ryJRWFdane3D0hN4pHztu2gAggmf0p6veZkWKAVtEIxUW5VkC3HCOeznC
t+qg7pbx09iKQyJycEi8s+1vlv6xbJtcVbxptlC0879GdCsrIqgiXczrggOx
jQFApqhuZfT/zZg3ggwP1dFEmPRMgKwolFqMdTDiwu+tbQ8fvRCjWP+g0P8l
biaktyizTeRnH/d+vfgSjp3nLxmDAjLOtfT1kTx3n3b8h0d3bOl+TBB3y2Xg
Ba466xFLDhzKZvjIw1WL/aSXIOLRpAS8zmvWxCyXSE4eJicR8iH/zwO2V5T4
pqNGghxAp4MiFz8BhhYROclyWLzRFn9KJh5yHaHITpUCUhTpiQeV+E84bAFa
bRBIdw20hT2/yo/n9hfioiDdpsRxMRGzYY1WVsjgA2VdPmTHyx5ibQqBYaXg
c0ZcQI6Ygz/dHdm8Hiz+iESl/dhareP26bn3W9Y2zOn6dP5ucexY9EzsBWxm
rY2RqueEDMNYvPeMtGCASXovUBzfxkc80ooGUYVOs3IlAjDgFgGCQZgrFZf6
ibUZkh8eNSlOxDEhLasnrlOi/Te2xvtNjCBWBtO/71knE1c0NKPSMQ/rpIIH
jHhHwurYZBj0STBkt53JEJ+ypzsum32ME7Io7+N6N1N+ZeVKQihe2eLeCXJL
6mD4HcsFirno96UFpDU8nbeFL4TNgQEhCVyywp8X2ySjSkHXt48kD+fTgURW
szXcf8KOb6Z8ezerJGWMK+CwtWUzB320jBIICETauKxvIKtySV32hwQbdyjD
IQAk4NOPznOZhTJ+K56jYwDL1fwfFkE4zZwt+9zcJoIRdm39jGcdlCUJmwqt
NhH3uOfQeRUaIfjA1PI9r43AvtgvwKOY+Jjf4KW0VIoRo4/6ZWjfot4NXnen
kaF7j9VPp7/B7u5QEFtd5hQYjcSQSbXNl/Kl828lGaP6+BIWotqrDDNUdZVY
b03tEA8+aqSa7/autNDzBCbiqWEXRB3u+7T8zPsod+rcuUeTfGgOtkGwQoma
F9aIHbiYMhiyB8QtstblvgDoM0A3hX7SLMVYcXmpsQ6h51w8+kT1qgy/v5CZ
WNMEGLL/hu4tQeCwZYAnBBN/JZFpH3wfxJVv9ZZ4q5h0fVCs8SXRHACh5FI+
3SHGDy5MUV7QeOtrh2bLRO1F3qslUCEwdnp8t+UC+2nQK1JGuz7kY5f2Ca4X
LFtjcsYy2GjYhmCgMFQpN1AL9NWdablsLVj6e3o4u+UMLae6mdrutitroH3N
eaMb0gwKWafKArs28H0cLvy6Qo31RebJeVVlD/VKnGrrS3flnszmWtmz9Kwv
b7HHsIGRwwq6BPwHSB+pEIwVf6LPel742VBqspj07tQztb3UVv7qvY9hP2xn
IF0WbQF1M07ZMjVpRwgk74Nx5Yj3PiEnGzdyeeW7ooxc7IsfW/e4JXuQwipr
AgtsW8s/Ku81Pacv4GGo93c4P/zYiGoaYlE2XYuFyAfx/X5Dp8tyP4PfUTzn
a30QLPKqO4SAH+VmI1h8oFbyM1KCb30DUD53rycSSlNS2LC1fV981vvlBpVo
zaOXBR4MSB7+BCy4dKYjuqAHHkIIBPZQWFrTLyocgha3S8XKW/2H50InMmGo
8Y2hbnMFaAgPZ9iiprONylTyGHnDGzIFGIQOuS+fScVFgPiLpI+m554zzdqb
Hzx4LvTYMDjME10ayXqTZf50x7wcPz3RLWf/zbd7cWx7C9JL0aHeZajjA5Kq
fOTMBaXaNlO3fDg7mL+F88wHdMwtdJlVOq/IQUwwOFftLvvPvZ7KO/8oP6L2
9jzKEmgS8hLhfFO8bfXDy8sF/mwBCvh00TqwLcPb8BRtcU8ZPDoGk5qsycVX
hZDROk3rnwjH7KfIy4kDVfIkuZS2pd79VkMCrrsrpbnSGiZEwUY3rQ+kTs06
X+mdUgrDhhmH6ZgMF0Tivhqw7wPdKZrQW6YapIwjjxZoKLEL1dP/3X/vcrlW
x+twdpy06DfuHX53ID3dJXPaFy/VOMAlj2+Rmyd3sTLvw6TZA95vAufEfZ04
pMhbywoR3hyjgvMgXIryseSIXa3FXVCiiIsjbmeS2/MO3bhFq/2+vq7KYtGQ
B9JYrINEm1RMDwg44X8RAKSBWfNLPHnsXqkMiUNgvFp2XAkCVFyXGQ1KML+V
m0Ci3PWaYUxF3cz300kiDnK7b+HDWrVno26eeEzOJeiMJwLMuMC+ca3kWT1f
DcyYhZkSTPYLcNvUZ5gxR1sSz/Lkh4LIwa+GqEez4N7+lqMvoKYnsPgE6EsH
YvbM7IlQ5ZPEARAFb/t8DNUdmY+B3Wj2NPd8Zevd37ODdFDOs/RgmETTuEkH
Us9M0NPZLDh+TZUvSOFVP6/IF3EcmQ7LnaDKhOEOK5uVY32JzENCV6A9XXgD
KwwR+k+1Qq9jrV59l5SFT3HmUvtuVG47gnd9p+Jg1nHwLYfNPEJXI05vAdB0
WHOV1S91js+5Missn/EEYWs0+4FKvKOWkF7YalsFUwyfqsM9MvQkaxxeO2aa
icnDm4dJiRYYLIuy2a+INXfQk/KijdN4eQXq0MbRUi99NUqBbGc2Tg4ikPwd
TaOpAiY/TQIa2yUkMIFRc9KXgT1n5nQRgxkWd8pV+oJRfAju3GjEvq1uNkhM
k0O2rxb1FMddin7yPf+YfhS2+L8XtqV1Uuu5UaeHKQ0HSoTXgWUkV5Igb/fW
7pNVs6ldCCP8XMfRkSsO/joBt/B82gpgZvRZMy0eZLWi4B6M7Ca+JX6qC+/v
s9hmmGE1P9dBZTfzvGEvmGGnUzi0UT+8MeLRbtWchuPCD81/M73ExtKjlpBM
QC9IwbeOSQcJkdp5ku8cJf7hZ12FVE4CsCRQTJPeqqTtXINX5ZL1du+3kW22
jkRdQUm9LdUp+Pj46wXiiCuuSRgvvyzOlzbJ7pkFeex3QTzZeOpc9Tecz2h2
/6uJSdI2HCiruj1EW/QYx94benUzxqb7Q7cFvXY71Al6iwcLWxp9PJ/oz81r
h4CojTikACntWb2AWxWXeyOrjL5VA+/8JLGEBsKVJB83uiAoKAbYLvHZZVAy
ACeSOzn7szFbh26ff3oJbc+QCRgFlATQlV9mfxTNaWopQn6pxlVdyOpdyQC7
/Dsz0NfqSMlMfHWozSZFxQMQlZ8soRgijtO7LC/Mi1Qv+2pKt0PuOfrIhzjv
xz5gEXn6gDIboQ1J8XfLkr8fy3muGwOlzutKKw3T71AroERI6EsSjX36Q/H7
OGc7kbHDLUQos6Se0OOvI/CTm62BYgGOvB6BfuEvAb/Z30TtQUU6eoMADBAm
HWwGiHi4MQb3W8gaP5wLFn0zCXryUr7H3ZZ1QUFhis0JpqctZsbcEmPWESeo
7OPi58ZkND+96ylZOjwuy07+nMHj+wzOg4QXMuE0DaYRSduh5dHQbUOQ07gB
KXYyZ4QH1dFziDXdhz2z6U7lYgRGuo40kVxfJuMDp4MJqm6ICarqX7Wf4O7p
fKPtylul/wsdDVHiitSWk0D7tpcw+rS+6auje6iheTnEzB16rJHuBZHUBqB2
y+XDRLPIEIcmJTqikdD2vYqSGMgw70LK6UOTuQuanpjxXWAvoVXBPEHV/Qvm
aXnyM005HnJcCdzdG6S/V77lBjGiidVUwS/UKMs1A0O2S9ux1tbdkG6p117Q
qgiVkgmMb00Ercsnib+sSZk/8EumoyYod/OYQUSSprPwhMTPY/CqVDzifNmk
evFt2KRFThChpRh51CC2o8XVdj4d0F1L89qt5QFNSOmAoRLmgg3opxSuB+lA
hkXDOIDZrgxvVjSl0tZSg5Y9tIiSoPL4GBjSBsGvhg89wavkj3mCJYINb6vc
+UbLeH8Gh3eTkuNY0AfiTs6i7rfRG7nwQqIq8AaPr5CWDu3oQoesTrtRh7a4
EBGzkecOUfTGvWezI8fFo29D4QluM9nh/E/LXOgp8QYj5QgDv0SWs4UV2of7
RT6oJsyZsywtoKFavrPgOezZI9gJsiVqGd9FIGhHWuKJ0yh/S+CccFzzD4Yc
W8eXvDbSTRtwTroIe16inBXTvHQC0tpANqaUhZrHlMhCmi2Fuk1/67c0dWQj
RZb9pRcHVci7ynlv6iLOqW7Q9HEemSWy6D8h1gTQPW3uwTH9rTeyT7pauXI9
tbHiIOLGveodia709tAlluAu76RDSSu9ht7d9IUbaJRsM1nlEMcZgpSg6kKp
EXvO9MgkSKeMjXEJJgj4aJBwP9R08B+Rd0iLMmKdIhqCSsjUbLWMYpUOH8hF
HBgN2qfohDE0U01rUHRQjxGOHbNXjoWyJExvTs9Lf+bdI0ogE5rivI7Uwm7T
Haf797KuThc1dpPfjCZFqik1S3/obhk51XBIB4P1oX6qyocfSPLgXqduRQB6
i4KPVLc/SOLoxqz9NDUpL4UYAlzid100ZH64AqE/TPVKqidcmuZ1kbj3sMXb
q3rKFYf2ar4tDsp5tje136RxMOxMEpvF99tjXbyQm6zgA3Fhc0l/V8pSE2fk
OI8eR5k+24h2B12aIbpbySezMm95cG6oru4VX5VtVSpWR4+pErwMmipkNzLv
aOztesbLAgY/HeLqdYiTjJ73/+oGqBH2/wCNYca+7apzWoJ1zv9V1UHfImm/
7BOqQkwrLiTT+3Db+1CGx5L4fAve52oeX1M+bTFnSC6wXfPaIeAfRh+355Rd
3Xuk+Elct4RJxMSwgBlNuTeZ4sbjvTKVrfAe0HYr2/xdIfi9GEXWPn9r0ZIO
SXjc3S5bTxuuTXBct0EKcIrGVedT4qeDjMsTd9m3D2edt5AYk2ajOxyGS2rn
VILf5EJJzfxK+KZuGCTIQkriKdvy2E4obXU91IYUG+jw6jj7GhYsjVkNiFnl
HBNBnnqrvXHiKTRVCr731jZKenvMJ7AkZl0NyKxs3fmOgKk+usjTi9t11x8p
gvckbjOGdBORxISvHgMt6zYczpkYACTsTB90M6+fKxLPvtlDTYOvEHhdAP26
x5ajWJWTcCXpohY8jpBnKhBIoqhFGxbx+0mhSlMXyB/MGIzFy8KF6gCjmZN4
Tdq2duNLa+t5ILrl0lbdTZ/KyoNT/c7l3zdlgEyEz4OIaS31MMP+wR1MGpeg
wFlMf5hCNahOiROek8u2gx4+gkWC9LNQNGo85i2nuJJFNfRnLmMDELq7FQ4e
FTwkL8UT6AohmHlg464lL7pTJf5/pxVAJswbAvf8Azd1gdYL6twSyDbBPwmu
dtg/3jp6gg5EzLq1evmQm3u6Sd32BAyuVnVsCkD+YNUiPYsP4XwvXEdSqfh1
qlVBJ98e4VikjdMuUpTOnMLI9dG0bvhDRyIqtj2Y2k5FMQftaFDa5lcrz43U
pL/B9JZWs6OlaIiz5tNuuknSJpv3C9Lee7yatcfKmWWiurVU5yJEJ9d0XTsv
1DMTWLCRklxBIXd2HLWDDMQ7RRFBD4q+LQr6zeZxeoNXlREQwZ0zDtGVsuil
TlOGY3cuHI33GW8d9sH7ehViA+bCj/rDKhxMKWashpcxb++vOp3UekFtiyRY
7MG3Y1uhfhsiXD/eKxHpjPf9ZQBJgtNgfXGzb1Yfwy6FhaVs579LQqWfqidx
2va/3p6MZrtRe8N0PYnMRwx6la62T8qLFfEKBuebXrQI/yw72BOfQxw60OWE
bJAcqlKZto6+51EDXS3lpaJj1gCVpyXHxIMCdIjyVP0D+n0/Inrg9crqFfgk
1YQWIejbbDq6Z7r7+mXgQzXD1QIkbNcsuBDQSq2z5ZBrYAV1XpBEojStdc/9
S91JCTSlPklrXbQJwqI0pFXrlllrdsZpXh8Djsuu1UlDV6HwTu59bAauvsCY
ZkwTRPGnIh2ioYfoJeo/9Bq1S9hhu8TcZHzUPhRcD0J79DMuSFk4acYKj2u5
7PjpEz9iY/1cPyr984Au9KOt8Eddy4JDJNWESXSDlA+JWB9pNxiLDp7bWr2F
KEgL9K+qdFaUYbOP2HaP24SGU1QAb04Pj5t/a1mr40ZlShaMADfgXoSHYhVg
pq1auZ5Mgb043OnhSQV5CSXHB6elBlxrQmcjF5VzMr0PvrJUNWXsi8LQDh+b
Ay6EhXlj+TFSDZoY/y01w+ksuaabMasY37drGS8hOyxlFd/bD0ux2yKArMe3
yLV9pLweo2ibu8OzmdpCLJ2mFps6+Qux/5U2JGOGsSSFe4UiOGUBd3tk7Xte
nl2IKLTQtGNbp4By+wMwj55llu3gJ/kOCwpD8iPkoUYmMU0i0pzNzeMbW+tq
1kU6iWwm5yDHLgot+6oA7cwTJKWWYfYPsJ1Xnz9T9kchEk4VLSYKrE3QlcLN
5Hek+D2ukT6/aS3GZc2Jzw7t7Lbwk7CnN9guVXHzw3KSm1OuZe2GNpAALV3B
A7VdzTEcoeE5k675vcVF3n3nLYBK8HNwDmRxq9yAbuFEKDu4H6C+zE/lLUay
dNEc6YXl8PJ4IzaiYdQoDfc0MxNLwkZVSqH3rbfh6paY14FaCsbrfVBPP2d4
eCnUyTnuhD4eeLdMrgQxzZF8vEHvXVVO1frSTkIXS3Bh9MK0G4reo/huarcY
HB9NcwzZ7FntlKVL4uE/XFKqBj32eLxFEeR1pniiYqEgegt95GBRzfAfc7aS
Gsl3IVJjqW+/XcDVhdSqPtoyMsXuvXZrrX0JThERG32300P+gAgew1kpslXK
bNlkMtOURwiQl6kcNq1BEGpHm1n3RGzxoe6ZxM81xujFsTIYvVfZqpErlqG9
OT7KWO5cYDr4WUx0PybkCWSZlUQMBQbpzn35QK0YM2g4L7FurtO5dFPtFYSN
BJtGMIINI6cAMsBuzIgO8uDwQeL3EynARMWtBSXl5o2de1iISDe2XWzB4VUE
6BDnsycjbCpRvCTp50fsZdj3eGGK87e9wQUWovH2GqZYjCewQAZBAIu77EZV
fNgsGX9fTCy+OvC6pCJ/7M/+H8/oPHLFqXsw4kGU+TpMsCeLJBr/IxfOlgYs
j933EK7fBBcihqjaR9GCpdynMN8ge6xMdoNlJXhnAONSmRqDN1tkeh6p+uKA
oi3RafUy5PFHorLVi40jgSZBHckNGFc0WNiPsl2V6MgRL/a4szRHFhQXdJhy
0Kl7LxV/42Wi38GnKGRWF3t+910VoqFqZoSEc1Z+EerQod0b5Ys2VFFB5Vw/
ZnJL4s9Xa8Nd76IuQxpxY+rfkbPuOAS9AkvdmipzCRUg3485z1utfWu68gT/
tJhRz0xYsqNDS/ZyuJqWYR7Mk5dTGArmzlBvdkw3Yvs7rh+KU6Ab6MAaQShQ
NYDcCHrlTGYNI9w+efVZcm9qnP7SIFNcuxCLqnu+NRBgHTmcY1r9s9CDLNom
9ZVcReKtN/x+Zr2dm9zamDCigTXGspv1t9EPCC8YkXo/2tiFdA+qh+xqIs0U
Y5ueFdmh9hMVswl1xvbEiWcs+h2CbjUqUnH92CTYFsrseC7a68O4eLtvnXjN
YkN1yTEBEeoG96xwKaRc6MMycsQKuQvyVW3sBE2jOQBHJB3EPlPo+IbTDp9T
JKfT4syep6sQgzOI94teItraUd250YQ/MIHbugMT4HYVWejvhHG1d53pBUX4
MfhyCxBEmZLxJU3fgxCrcyBV2/NGpLnvfXQi+lV37LYh2PDVuEnNgp9EqPPn
fWM8A7KSUaHWmOC+5CYKMAbP/2Lhl198VJc8hz8hAokHHxxOgJ0r6q4TWC1U
WfhYl5SpdAAfvlziX5OUDxi3aAuCorbBSJuxtRKHSeAZgng7tMvGqza8oGw1
RKDuXKl+hGKpU8JXqwMHup81dRQp0YBXw+0WsyELpZFHAZ6bxn0hbozzpwS6
JqZgIWrjZMs4mDMDQUrG6xqe05TKTIea7POHpRcw/oARHpy3TB/395Hg+8Yr
+tZGkRRydS1gi7zh2DakLLVOp8IYD+8bfR7AbIlLub9FfJG6MmiSJ3iEdzAP
RCw0kY5qHxSx3b9qHLQokCGhswMcmeNrKsC3GPTb7rcnKYVwT1RX4mLUcmEc
ETILNQEgmDsYFwcLidYvnvKMVxRgs3WaLpnAaR1eQSY7pNO59Bxu6abjBVQP
jIBbbYBn/QElp3+pVlRqjJgB7P519jjDBVpFA0L69QmqpfhWIe+GVRr8RrHc
NH5qstkJ+zIqFQgnMSaMhRkHVQU/pRkpxSj7try/vv6zmR1e0x6IrlD2tVX4
41RejOVjf8wz32R8Byiw4d0oPqI1ALUN7k/j8RSVSV4+nV7SLS6XcfXX0lI6
WSgJPCO+W92qi53qtiKu9IMU2yhrGCrLy/eDxTEweCYUT4/STxPtxS9DiEp4
Hy1/b1WEqpdrGHemsQaCyqLjP1pF9/KplhYSNbjUMmqRWMl5lE5Mp7905Jna
Zoum66ODi9DLEGunOxU3Mj5UPEtprTQ7TbNU/macY76iSqdDFE/U8g09EOkf
3hCCmvrBYk0KNLwOLV8pJwZ3n1jpA25KXGb4cv/wP0BperM0tjkbytmVnN2f
ZyoJE6aPXgkt0VTJVQ==

`pragma protect end_protected
