// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HnTcbYQzYDF/vC+/IyY81h20OmLGh6YwImKoOdIll0R/8xdBuVwz2bTbu4Kt
Q9LzyoPmkQh3jiCN0O9eIfz4YMSTO/+zA3bIgJS87WuxaV+yAXHYa/BKDzZU
xyo91SDDrKhZB/5Pom5nHhC1s3jBXpy4oPwIjdOO0C6b03HuqZ/PtohEhUIe
Ax+0IPfdAz3q+XjRlOphJrdK9aLS08qwQ7gdX3bRJJPkqI5bTSinYEepk/Oo
/CD2ISFyn1E+t7hZJrwbc8Jz9qIKgmDvIg2Pt25aiR2TRxHqC5nrm5SdVrIU
Q8rUuPmm9oxoD6H8lEEnDI0LqlW6fsVsHdbcROL3wQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jmSXQwYaXtW0RrU5TMcGfNpHX4Nrt5GL9BeDiSmuphByHIvetAE6wYkJ9tGR
Lk1EHcQTWoFUUGCbTbXkOvv8lUhstBt7FbDoIAJHWBcpwuG0Iu9/mm7ldXm2
vUXc2SCTBbdtuTfHV4SFEs7NhbjnCJlq8QGhsznaUTiF0WIXgFIIpmpH1eKw
8rghL/ZP8nLLx0F3y12Km5zBuuHCfb74ixV8OWQ5P/Qms5+6DtbQROneitNC
G7g7Rc5azUyyr2PGx4RM8ZlqvGsPMOxELqWy3Q8qx/vnZjuaoSZCUrER4gAN
npmeJme1iw7Jo2calKVDQiHWmgZJBKfu2WaKU7ugCA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ehs8d2R4y2IlBGW8uwDnvP+0RPwj8ZPaUFY8COhtucEV45nqMolU6UxuL1XI
9QsY+zSAuzQWsFDpJrLgWN05XbQDUBOtRI4fVO0wZTO1nZkknACRLS8qv84w
oSL4IGAF2V5livYeQE363KUwWuoR6+LpSMaTgN8c17LI7RFDh81rpwUOiRYh
Lc7kOc5+Q2nn5JCZTGPa+jxOiNXw3+Gz3TzSqFjb909UZsjCBl1+PePVo6b3
nhuxU9KodU7q5NyQ7G30xbBV9t1REm5oR7KG9jAqwrK6+cJiqnNuqiJtI0lM
UerR6azA+5riYuYKw2UCSmHAjure/Ly1On4gRXnduw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qffDmewN0So7xkkkUOqM6TFsYOzqpGoRDGGC5346KXOnoVcdBp4S6ohUJCI/
qtSA/MwuiZnXIgU1k/WPTy5wec0I183da4pAdWrXB9Ac85px/9f1jMJxDvG2
sM6tLE+WJX/x40oJCCBxs2RM8d7a0iw3ycLv2eRd1nLdTzpYzlI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uMeH5gI50bC1JqxMPODXFhoNhXzUYze3r4T20dIL6FnhHE79ekIv474HJ2QE
PtYNGOMeB0n9QHIV/VxpynW+OL1bcT7wVXQKhhQE3dgdghuH0F0nVXcFl7gW
ljcsToWDpNbQepnyJCbR2v0zqNUJsHrkaGwmwD8q8VuKZxVFm8de2tNZnlno
w4I82ew1u8KYOSEXrcNVcSsWGpCuB7JL4uYKV8tm56s0UetUTegUoQDWRoWs
rHNf7vRR4JknIJjrcCgT6g+xc6CK1mdMI24QLXAjMQjfgZu2NtRJSJcL6DnW
1AN/RKHbJ6sgcFXSMn4NBeqUp7KC9gQWBwQ8g2+m0Qe1+U3j1Zm5b2sdiqkW
u5DBOeWp0NvHOFN1nDXMViFmhVkxoOft0LqMadJv+CKCUntsoW1MLWEyK2GA
XWZ3Y3vcvAzB87bf6Ok4bRt3Tw6dNTc2UtYOnksHN1Iy4ncHm3+p9KdkP2QA
bjxhdDqfxWFgHWzXefizkStQIX0EKtpc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
A5SeCTfzJKxOGCUNWtIrsvLQTz3k5a6rcQrWYVuXjpfcHEkZCnQDzQA+tHSt
c23ro/tek1p0+BP165jBom+Jry2QaeIRezG2xuHhWGQbCdSyoTGlRx+hEB9O
jLKoI0HT3D1Ny5B63+oPOwcJEX5IS4cYqfIJ1eNgpFBEi+zt/V0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IBEtew+2J9Xtt9f62wpBWvZK7OkZlwNzVGOgy0qMkl8JXNj6ZkOCKBvmH2AJ
9+ppe1MlHLYqrLBXEpcoWt72vYBX0YkyDRnJsflmpE53v69x5JqU9SGYihG7
T3bXhUMJs9ZsGUMmV3Si+3mEW1Okt62l45mQZiM3l61hVnMCL2c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
E7mQk5cZsZOMp+s95f5wNpbvZ2+hGBwFtoOy93IK3jxwPfB4w6d63mMqnA4q
/3n0vHA/lRcy6MGib7F4kaitkYdRRqBZn1Bpkn05Vb1tXZYIEKx37ENVdppD
CAWq0NCtges28PdHGblGOzZjfat3zpi2rE/vX964h5zUZ7201kY6maro7JgB
FsLYKRWnOlCJM6LiQcU1p2Nvld46O4sg3ttTYaPiv5vpbrOWDDMk8h0TS2tx
g8OCKdTLLdm00iYlBQq1Y2qWUc1YmMXlbGa6oY08IsX0qV8AgoypM84D/iTn
eOjih9Eh+e/sLheBAx7k/UzXXov6BfmXo0uRujdPhYyGUQL2fKuRB2NlWkbQ
phCBZ9VE18e8KSL9+AuOlYEwXcFsdjsodbCf+dO/PtcMRjgYXTHUo5OWzgTZ
FerMO00cu2al9yxyPHwXmWB3Fmv8QgelGQDuarURRNXMbtR3KonjPHi4U5z0
19mrCQr9r/TJUuWB7Cxo7JcQ4psMQWhS1FFlYvQ3QAE/QwcfGuNnapFoqgU9
nhVaCmzrANX7OZZIs924bsMKlpdt3H12tXNf0F4fJZm6RJKe9Uuy7n8UvrHQ
QKoIIekH3PR18PydNxbxtpEdCII1zeKUWvHqVbBREsDnpYdNCt1X2Bx/PbM5
Z85uewRhzC7qAkcTdbWEanO3O+jjXg5whhI+kCJs7Eo1T7pgl4z9hfC5SQj7
eMW72CC4ReWGDxwB/+XRPCH9ogQ2uAGJCx0dE1WCYZYyCgFswELMHjRd0KFK
E0Frd3/AjnvG7iT+iB/IccvcO8xzvW4vZGEwTL7mrVuxEZ/AiYwgGFpeSGQS
wr3w/gb8oFtnpA157Gl+9hu7p8lHayEHxQqTA/XSIYLx2i6reddo4b/10d3Z
Z5TG657WMVy5WNcExibdP3Kfjo53NxqZl48OjEMa6qttaHV6Tp/MuKDav/n7
0Tqnkmi8ZKXXJaduCzP4KK8/i4Byi9HwE4JTxiMobQbwciLCyHcjCOCXL2N8
d6kI5rwhN2TNW8kK28rJHxw62rAP5otuu+6fp6DnZrVyD1zv2IVpJOuXQyiE
Y12jmtc7+DuLnoqDUR5PdgY2HHZIIOXGy6ZimzwlZsu6/lu1YFhqPhpCNIyF
d6NvPwDHEQcU30SS6yGEPldMNhWaPP1brQqlacLeblQqaGzthuQfzbbnFNef
sqZM/V7ozNF2OSBvGuto5UF47BDYeifV8b7Oz2+ObhtWqd3g6/1Ql4Ph88kS
ofZheV+3BQ4GeWB/hN0IQze1NoqOzRBQnzRLAdF/adlmIywBVY1rEZkU18Yd
+EAavp+BSnCZ+BAewjBRpEikw8/enAFsh3ufzZ4n8innl6RdHtrD4+ZO4nDb
KZgQr1fMVNtEhUQaxSVwkZ7OlGKoTtrJedd8JMYUgt/W5Dqwn6LlhV1+QLZN
gKV1A436bgJuYcVcL4zuIV/ZlzhEkDtheQvbDdAwQRGD/qGLNHKF/exvW9rh
i/AsTin2M//zE9pyzi7llPZZ2b7dR8zfMMkahveAhkI+5jSBUO4gddd8I3bv
G0Oviv+aGAEnPWVkynnCt9PnFvqhgNVZjluNW/ALrOBzMp678e1rSM8l0SpP
ZUpczbdjiuB2YIIYhcnrWe31SmyDkOJhLht4Nm3CP6A+TrYcdhm1TGM8FXtH
Oucjok/phKZ5juFuRXFdE+FhhVPXUPMRRWhtwV8MWrd+6m9oSwEn/YILQfJ6
cnSQ66znJA==

`pragma protect end_protected
