// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
NgZv+SWu530e0LhXv3voqhoh/Ln2IaW7A+KZsTod+sXuhtUecilvrgna3jv7bNo4
j5CmgcnYtdm9NtRntIZvg7lS+lo7NnC4aaIhn28HOGoQQ2xcyAfPRkPbRL/LcTr1
iAk538mU0JrwUtFv6703IakhZM5taYxbB/SzgOayDO8omo8mU7SaBg==
//pragma protect end_key_block
//pragma protect digest_block
mrsMKT6m2+eNDQe3vsMc5cR537E=
//pragma protect end_digest_block
//pragma protect data_block
BgwxSzQd59zKB8PQ338I90/3pc45uHUKhueCI7FMmjhISemBiGLRn2ySodweF0Vp
z/Upi2SHNpfF/bUI2crYDNNQ7UxqUIjKn+fcIZNRSJpwEh686MthVPqWhTkBSe8i
z7nKvMJLZsD+H7jOHh3sGtpTP8aVVtHZ+0JmOpCCt99jCZGdHa80ytUGtQjOitHH
twNgRHDFEjdpZ1DVYtAuE81mDrOS2D5HHM4cgpdMSx4bt0KnEmlQ7c6DU/xo05Au
+UeCFGVIeNX1Z9TU0MyvYXU2bsJqQZpjw/Da5vgibhMPWPw+welxs6pHKwrP8w2K
z1WvT7NhGC6CfzFcxN5fWBa84ysgDaHgUAkiYgQNjU9zrnFTM5XygpKN44ShfThL
uLduZ7uOiamiteHUpVFjcZVh7+U2UKfhbY/EsPsS28qXLUBip/J9oD7KTPa4Bwwb
nT1kc1kg8DUHWGfT8OWHhvzhhfB5AJYDV2esPjVytKvhZEm5UwIycg/lnJPjpA8l
bxha2DzSU/SSMFxdFhTGrO4HBm5LrzoGrZD9NwFYai0eX+6gVHQb/4EQ7UiA6YgM
eCdB5GtU2F37IBB6CqLqvvVxhZgIik89iBDcl2ujByjJuEA/1iEBYI+DOPJ68kDO
ntKQXwGkYdBQSdp8hMMjd7Dw1m/qzd9o3m3L2/ArVRAOzyRa+phadpt4rkTz3TUE
wbHxXbIV38fd3dgUirypTzVpcChNKTwKo2G8SV3WUtrwwuHN2xHJm45sXq0UOnBa
irF426WnKzNPhDCulMXUqgtViL+aTkCVCn5t46B4kAk5r4xNKYS0312G7uMIJbLG
nwMqaIGxi7kFp+0HfWzpc2AcoZisfOBOgWYl/vQpxUFaKb4tnbdHUCL8TAUwi4ld
8YhTO5rR2tSAaVcJWdZFeEvfa9n+ZLOAFFWG7Q0kM/fiY2/exwC/sLRXQQvymSEk
noh9kbYEg9HcZ06sWBLCFJC3Se7/3z9I1Td9Bf/y7JDNGzAWTji9dl6NVk6UfCOk
++BEpn34DuTgA4fe0mxRRQX+UdPbOGPmFJh3vDFciXIsNIrV38NhqUInuhTDoATf
VfKbuxrOk809ZmSABsB/rkgwTqQ4zyTHrMA/2xV98yTAsahNyGV1rkMpWD+ox1J6
7l5mUz0oNiXOdGtZ5A4grkmJgm4vUZTwiNGbnPnTa/j3LU3ek3aVYg5HfDAtUMbi
c5OD+X5ESBt8s74FQpT5LykeDv9p5oS5MjYmOBxBZUoC1aoIW4MUhAL+oXy4k33n
gnMXqOJlHvYFVGLx0DY7tDVDQRN4Tz7s1J+r1kADwI5dVJu6EyPc5CU+QpVEqK5R
8yYGClmW2/t0n8eSFfdCqUBLF3BTVuux9l9eZma+2P+DORhttkK+wSTszVJsnuI7
Oo2LdN/FMn+QAiBpjB5Ac9DFuj+JVF8sgkUtERCtv0UhNrDcUG7Y510Y8FY/8aYb
ANwJ3fa5/RrvDOo4hkD9F3Snp1S51nqmEqQlvF2DwjsOciBsAGNKbQLoWXx2ds88
8Gfk/KWITm8HL/0tyW+h3CCG9C/zCd/O7O9vt6jteRmklBfQyjXYRP0yAhHcod1l
JHuqtJhx6jZLsLIyBBdfOf8GRZgRkiI2R0IV1m4bcw9NX9n0cqjV8oQd1v/kuKcR
MKkLOgLT0rVfp+xddWeTveDM7EA4aoaNdR8QydHMsC+Go1z33An1mj/RBKC0VfCi
obbbbJeFVlg2fkmql/PjSdp1iEdeaGUXKqzMy/SVNkrD+U0lUqleF3zh7jwfuvge
8XwPEY1N7Aw8Mpx+zUoq4Foryh+bdBo/l9tzsQAp9BkhJXhJwdq9rT+5fAhseGY+
QQbYnEbyWZrR4pAjVV4FrrnpTGfmIUMfptennehugcENAs9KfoAA3n3yEpzBm7uC
p5zPmaDq6n0ixspCvxS2JAU/IYn3amAYgkwk59MfPkDvEiFXQDISHMQTxVzlC8s4
QI12FV0lr3IazQvpmY6AxkQHAv0Ux7sPP9XLvpclxoosMulDRnjLlirkBq4O6KbY
/WWbo6NoLTE5huL80ohYulJH33rPr+K9SkjC07vd9MJhkcZmSB09o8oE+J3AivWy
Eyfud8VPtd3h1GHjfKUBc3w4K+mVGuKmW21WFlbemqCuT/1xFGX3II8MHjglICwp
sb/a/sEdCZqPYMnuJCc1ovwy2FwLdmNVWPhKyW4Zpe/u0QDK5jYJsBJn4qssridt
2LDmv5KOTri44za7DlXIfHNvtitMudTnWV0jgG0HG1oYb6man1d/nB+i5BQwLXso
J5kSaYgb5Yl219LdOO1NkbBH+u/rz+1LzrZMGJJdjGzrXmOWLTtovTeWvSTt1+Pb
YK7WnZluzRr8jl8HYGba9u35IHnaHdzSz+4t0uh+lGuRuvLXtqCARgkpR4+yWFg7
PvN7/59ge3UviKBGe5YHLqO/AlLWUbwVW9ivOAJ8etzRKGmXj0zyr7sZpOJdV3dC
fTpe5TU6XensBAE2DHRfwHe+LOilbSxyqaT6UagxJPHspUEdU8tFHLIiwJpcIvye
XIXeIgcYnbfysTEaA8+YRjb9yl6sHqccf/V+TNgIrPkiXoMEZ97yYGPlStIsCyTy
8jG/jNxc7xWTULsv94NdL/nL27yVSLT49Ka1oLicDp4E5xkEMr1kCcC7LApi5Hy6
3v3POwVhlXRcaGzQpkFFpS0Sjhb+n3kSCQm+xxKLPLp53OmbjPo5HFtdZffH7o/j
WtykmdJidwLdWqOUpsxnUH1IsGawN4vtgnG4Yy1Lzuk3HbQ8ZLXEt1JHZr9HhNsM
Z7bxiuTUvzR5eHra7QGzBTpbOzZfHY4dHc8vk5Uap1ZsMRZzvjPhdd9M2rPzSxDX
INxXawZNLlQP/zGHdiBs6dmiJpmvn2b7QR3ct3UnrZlsqVfAUH0YTmDwDcUWUENj
mUIkXCkXyX9qbrGUB2y3ynbVI+77ApOuZM2CodPXRCJ//gCQg7c9bmsi8OOx3tbK
3g+uom7f+Mkums4X4vaCyrTMIWLZrL9mfhWAkgekz/GhekuDb7ZGi4hXd/C34W7d
ZGGO1oDw6Ig/khTd9Nc8guR2ZaXTvaeXNtSo316FWTckMoo80IKGza3s8oUQSuMc
7iEcuLq8UY++5bpxRqdA5/0pDsrOtFG1N6hOpD/b+BI=
//pragma protect end_data_block
//pragma protect digest_block
tO+rvVGhehdt/GPD2S52uC3GS6s=
//pragma protect end_digest_block
//pragma protect end_protected
