// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HlKtxsg2mI9R/luKASIsaLVKP/952v0Sqte09HdPZ/B8gL6SPpRYUGjYkKDC
9aYXYnKIbfhzn64Z4dv1Lic5/hON6WU9/bpCUHGbxiD3dbPpTKZJviNlWble
WnRj3ezk2+s8fjpqQ4Ij3ZVKU0tulr2wSl5exK7IGptL980wryD38UzZsPcv
aUZzyfPe9BuJMdvzeCAbZPbArYTW9QGOi4Qcf/Qw9QP9www7zt+K9TqVo27b
1pLsdw9i0tkmvoGW/T0h24Ruh/OGL/gDLimUlIDAoKM7XXDA+0OdDRCc/MnE
53sB/boo21ZeEfNQpywFI7jjM+ISXoJbXVlOJNh1xg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BJkgBdQz+404iFa9BNTXyKcgmNTnBR3A+BtrCwin335oo+gP80AaLZvCE3wJ
QhA+Ol0RWZ0om7GLEokYaHlahgXVNXWEcZ/+VJAzyp32cEbESNePpjk24kh6
JbvGChoo0XFcwswsOyJ/TgyRDYCB2BL03cVwuz79XqNJ9mowARDy3WOmbYVj
nRd6B6mSZfYymr91G5ZIorNa6DYZAM4ZycWfTaGVdZ1IQqtleqB2GAiDlXnQ
IFhGFpMMLqQaRG3H/Q+Bsv3qDTg3UCZfw1mZ2NZsuoEmzk8E51J1aEqahDNt
WMKdyjwiLZYqzDIm+pwa/m6UvPVECH1hO9Xu7E9t9w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bJar80ZzrGXBjEzQO+dUoeIo2h5egHiFESNDMGXyvChSQPwHzvr2UYClhtFB
AKDb79rsifJguPc4ezTa7s3/erJV/hbLsFOXxhV+MjQV7nySyQpnyIIgJpx0
RCNSg4F89onk7si5Wmq5QgknhBJq4OI0V3iJ6UjfZFJmWNUyaoZ6LvY1tuxr
4HKNjS8RCp8mYPAnJ8NkxHDhDC/mLWI21uel/rZzdG3BJS+xwD7wRDavjoTm
Zdl/39rSM3NRFPGxuQV+aQiRhkIeMITApoYyxG5iD9d+8iyBd1NhgFCzoD/M
hY4vLu7Is6WUl5W/Lp3QmZOz27lJ9WLWDvJ/7dIemA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hEi/L/s57+MQcXdy7sD+MihcduHZlGw1K0AZ/rvWdSLud5vgD+MCcpSaCJC5
nOtu8Fl1SHM/YI/hPIc4hHDgKRxUEF/i8xqHnuECx8F0Hn6IG7pQFfvsF+S/
0jMbjlgcwirsYwB8pTgaoJu93RWN1ch3BgRfxQteOOoMyd8ZCi8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
P1SAbkB3t/X660mfb4AKNETfDqMUS7aoALT1gjdaFoIdi4erHqdncfwXPmDl
ms9BzToy0Fa3b0+zmNTrIlR0NhXmCl1uU9eLSFf99E0IE6AG2j66F/stY7sC
OPaq8amPDqGJvf4UvRJk8GpMuxbno9IR85XvfiEvueDFI+Kbh1LHarZTIl3q
E05LmeC3IMGgG94G8H9KoJ5L2XCSO+e42RLOrXaTygmhjX7ftSid4L1GOtzk
II2uyzY6vHoGA64wy+Tz5aJech07U/hzVA2v6ak8RqpF5sJ4W7QrHzL0Cwk6
DP8fLFgVxkrmdmCmARX9w1peg3aDIG7+6L+wkmPuAWCji5QAuLuf1HLYrDw5
haZIivLT+mg33DawFkGzRXUEMeE0M0HVw3van2HjwmgAZOIfKZZxEPp6L/YY
LNSqBgHYrrJmAsdBQds2LoJU1y8al+fjHfk4R7u7ASWvwsQVlZgKfv19nNui
Bk+ml1Xtjyw8kpa94i8nWLhYuWWolhBz


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NLhh/JozS8ENIWJvlb2cCHhfbB6QgAzmxzAfSvy1rZAMnVMQrmxuvkQA8J6k
v028rS9d3bv8TBekStLndRGeZMGkdAh2XZxr21g2rPCuzGL4W77HpP2/+Mav
Bbs+GGyOdxDqMbvVE0mTHV2+maZxJ4yjfedAq9FCA7HPqmCII8U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FRKq3o/o8tPasNP+ZUDOxwvC6bXBpBUOhWuktjR2CM8HFqy8FamdP1C0JKvx
nPnZCTutBUko/beKV2HE8IrsVQYLOFEEwdoX54ljHiNywX2v2R4o9+A/15eC
uwcTG3yOT9WCVyenLep/xX7SpaqX08BkZxFks4ld8RWLuQ5npH0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1248)
`pragma protect data_block
Fp3eu0Wk00j6x3+vrkErnu5NO/Z7ABI7PiOtyjfua5T21EyObqrvCZlUzKMy
27v7G+OC39l0r52OJ7Cmfewlg5e7/Ue+U8OS/rzbrJAEIv/IGYY8B46foAWD
7+627yDjx46D8ul9Vf8u2X3hwY3bDpX1MhOlic8cpOqefikv4dM+UolVCvyd
s+rcO0qZfPTPfB2eQrPoZmbufOKFcffjIsNaK4Hhxpu4Hi2QOAOio99dd3Ll
1wpZodqXmjiSXSbI7igZS80GLF6QOuWEYNlYJCf1mPdQ1ICwYuUA3Z3l+ldE
rzau2JLQmnwOuLib5ooiC6LupD3m2AA6+ETKV1Tdy5DlNG1yJNLg+AmAJSQb
6n9QzMc2Pm+jTeogn4HB1mJ6mlSOMYtB+cSKOsHTowSQ0Mr7g0u+M+jfMXck
tLCk1AGak+A6iojgC7eKPuVC9XQasw++tIanCP6BKiKzKwxKbMIIyYgLWe4C
J5u/1vmUQxUh6vOd/BssA4mh3aPQbqHh4ZUapdFuLJe8nkaAN2u9cRoS56J5
23z9bG78LgFL4S9YBln8+qlrVf3qUzj4troSjyEL3dp0Qypi3W2+ypo0iKW5
ukbKf1CgGciDpCbqhI8Pl+NEBxNm/VmVMN2ImIBlEBQNKUq9qfFCuDgioraT
FpRtvA5uRMwh5ZV0ozrl+xysxoKo9dRYlysoua5VDHkZ7kSJq7VkIMzc0jze
hu0XrfafvMSWkbgDy8CHYbs8c/j6cRI+H/fsJ1LMtxz1E8txcS69hrJrJPm/
bfljfL6/KALhHF2gTEqSKOvPQh/YPrq2suZE7q5GaWKFSYZF+E8yzHSiM02l
FVYFDZHNl8dIrX/yUbA8BfpcN9q9rbTgPSIqAi2F9agJcZSY6iaQA9Cj4Uyz
L+hJJ9Slev8Np23aQ7VMHr6roWWSs3X8na1vGo3mmyQBOyv4HlxZecwXJt4g
11mIkgOYx4yFnuv250Bfw9pnaZdA4nCD1B8FLMYTYAV457cE+/npIMpz6SLC
36ks8NGQWSXAq4hT4n3LraOUJt1dCGT85xAqCbE+34RBwvxvlpIcy0LyNu1D
x4sc2BLp2NTCDWR8ZXdK5MIKxhIl7RkPNlN2KHmBaofNBy+K7NtpXCDdouoB
ePskqu9Nmpsu2ieT7udnBg6ISZ660RIk95flaYKPJGLwD7boIW11AdT4UCvy
N+FoSEI3Oa5IjqqwQsvQ8vAGgq+e19KF4nmoCpSm9QgxiUQUyKOT2MRhGVf1
uLIDNCe5x2XXhQKn6eIdoIHGQwLOblAgBtoMvKEW5HaxhbdzkWmQsD7IHGI3
xFjZyUJzlub1YrTAEIfwusnkdMh6hD/s3TVg8JsukrwR/ANioMUuzlxI5rRl
AxSw+0b6UU4g3AvE89L1Vx6KEgH+blauwZ49EPoTeK+7Z+Ku3EQ3xbfr43Xv
tukL9TSZUtEDmgg0JQlqJj/cQI3mSi8+EPbKV1bogWAWX/87BdUG+/kcK/yg
4qzhCEXHgUEeLmTGGi1oE29tmwgqlH4OPHODKQIegrTLz+ljL4TkTvaOYe+S
04rEys3me6Bxce/AyU2ISIA6BUg+f1p4xCE9bLXIpsoqK2qMyjhhEhYd2ab2
RpZOV/EtcZRMszZZzk4iIbrq5Thkr7Jd6Vw2sWNBZGrB

`pragma protect end_protected
