// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QtBaAKGGS9hi6FC7vlWaQnFDR4VD49tVOzvLDVob20ZNwTObujnmo8NSip/v
ylMRqtF/7+zPRxkClHB7WzQny8wQvgIELLsSOQ2JRWvke5TEasBivuTISILw
AIqJSpkzbHw0rMER2agA9ldjp8PkKpW0KOv65hX5DHGRodvXgn8Y9ErAmw5Q
i18fCWYQARp5bNIBp+lyXDXM39c9AzyaKQEJwXNd0dJAeui7YF2xQc00uABu
UUIkL+SGYsT90CNaHAVV31ZwCYsUeiEIwiKcY6bVIHFRD6ouO65niuyE5J50
yQqCLEDyW+QcmekfuSQuuvcnPoAKWlpqK+cGVOwZEg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c99GiVofYTxTbn3vo8sIbEAeuTBAVi5bG9etVdmHBoQTYXzrrgZVI3oWqeDD
DhgJglYd8TN7r+pBKR4ARFVOd8iwBiL2q+1cy2z6T7XYl5+xMcpL6Fb6ONZX
1p/c29K7neaVnd1ZkW6oKNYvaF4aAoeUfLCFHbHxof87KoyUXH4Opi2dAQHi
x7P4JLarjMBEUNA9roDYfUxol+AUB/LzMOhFpBlQivKqbJXzeRjaCyZqgPB3
6HyqNolE8z/SEy7Szgt9LbRju8UsMMTNTUYs5dZfBagJjLj6XeJB55OFnez3
UrsH3XoSpm3Rr8XfNvQ8zL52lX9bLiUpO1hA5ZNqEg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n4FABYrSe1fV0yQV0i3nJSyLqdSUTB88zTSkYpI1rcA0MN2PMUb28WEdvPLv
wsLTeBcMC3qWrENHjPHn4mPRpBkpshNQSv+02hQ4C7dhFTRnVLFWacfkp9e5
RRYVAbIbcPe6+jz68soM2SgVVUJO5vQ386Kr0OqKGHpwB9lEls9HJtPyqLRU
536jNWw/kOEtFxzj5GsY8boAGl6FZrgcU3Iu84Ld4OduoNo5fy0HoB8e0/j2
vsdkXpUTnxjMfG0kLucKdJEkopRW3VrSFxWhIuDnP58lyuguj2JcKdqFXUiQ
0Dm9klU6FZI8TOx/4EOHYBQHW+DDAgC4764bTkGgxw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tJuXWh6xRVa1uSdHpIyr2FUKsNgVe+6vcHSdO4FcCgJLVz8cTnenkx9ZLpR7
92YZK8+K4omHr0DviNbzbFIlDdCYW4i70kBI+pZCg7p8KmNByvJpKq4V7Y/c
uH9C2z7LmmYyqwzhj+zWbukV6yUo50veFi1gUFhEurPSloj/9BY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WMC187fEs4d0joF0J2LwS6fvfLwpZl0dQYXAzMdfy+T4HtZjQFM+Deu/9HqF
+xgj6iAewmBnbfGuEWP96dxOg5NyBRG2YcYaQx8wuJHRl2EmxmPcs3U+RL8P
rReqhnkDTC9L9TtodOmPUoCSOL3E5mbqfmI4JVyXbrLuG2b2mo+XybA6csLl
mk/os37VQ8s/LDFzlj1yxrheNVRLWy1lcZikZFveA3KmgsxPyURx/IlIPrB2
sxmiBbCBuYARwqfPt/czXHtBmSDbStL6mf6oYD2tJcZLnQNoccfwO3cob9wt
coeryXxxLRAW0bXodftUstrBIZct8NrHdxaN2NJX888bm4hPs2y5kuBrCY7q
l0lckUjaGz/g4FEnp+rxdtRofA4D9ZiAmO92/iQrVWpr/VMQhYvkQZ7DCOkp
+9mfhQ4TkYladsMtu11e3VhzenKaJi85LX9Qu8G1YcL0mc7+o77D9syF5kOH
tI3Usv8q8GUaBppfGqbp2lsD80FB1pxy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uz2R9d6GDbWGzBe4x0Qs+Wjn75vS7n9Zq9wuVpbrKEnqr31xQ+DJa2v7zbMG
+5vqEigx03t7YP27EL1QPHP904b9+d7Da8fce3x3uHY+Cgmy283pqRQZUwHz
TCpMXN7br9UOWRG1HDTMEPell/QzqfhtZnvCIDILfsJaBKzC5+M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TlOW+TN+nfT4TAq8tpJt1uzuE6bZ34sNQwrAobGQFsIK6LdTMsRvjhvl9oZO
JBcT8jY7z8QQMd4TI0tcgz57l57waSuG7Pwv1S06Pf/L3fdYwiH0Pqjzhs5u
RFg4pGaVi68PN4BOR90RqY5Jw/0PMER/st0ciETlb1PUdiY/Zo4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 35184)
`pragma protect data_block
4mYwTtHXlF20nHNPfnSx66QQuypYFUMOs7iPW3hAVh9zhnL270JOuMS+SInv
YgU/9d0VgWoM79DTi9y/C9TdUBUWe68OL0TA5gDwE2xdNzzg7U9cSt/cIiuX
ExAAzjvCxQh+p+8+9cKXS33l4uYQfdIp5X4LTrtmTZdM6UG114JqNQWe8LsQ
ghYcJjkv7iVSVjOEuCwizMdjtiiytvIdcK34VHTUiWsx9tdvBfM00mIDKTY+
DT1rhurOdXOihx4kkF8BG4Tk3uBbWeRix13ne3foajYOn8aDZZw1opbywN/M
Pxw6155JcA7IVFIcAVGOVqCeMpuvkGaNR4JBkFs9JupdyN+DZDK9gaoTEpFX
SraAB6rcyLU7IxcUNsORAJPJwKnhnzKyTWjel3bhVfMe5iMhJ3f4OkAq9IJx
F94oLzGLa0IrLXwiY7lSQ0o55+56gB5MRimx7At6pFKqDF3YI0hHAtsW5XfO
wycCQJ+maTXaGXzEzcKBhmuWI72pvF2oZs3Pv0PqpSwrT29RoWkYeCM6Ibo4
Wo9NITy+y+6mz8ujpwc6iP3/rtf/WOjsIBKlr+jbFkXhVRLxf75CUDaDUPNQ
QrVClwBIQRT0h98lAbrSm9IUkdOxXm0ZIGbTiUjSx+M9gIkI7xh9ubWwZySt
3qAK4zT8DcRM1XL1sCEKAlCg7pdwSRzYg/iHBN/k5rBGErXMnTdhLZ2Qt/F8
MGYG0iAxhkrA9T/LlVmgBVv8/H7iRyF9l3TlMhgTYcgJJcJZ8WlOPCUywNLO
hk1tnTZi9K+mjUfORsLzPOXUtYO38b900QeFMkxQAgxBfVcV4LtnH4tOfkWW
DNRvbwNXqwO1Gp5mXJnQj1+r8r8MJxQthnBmwywtu9fEVtGrm4YtOMa3HpyH
+pD8IOzw41vSCKuBUmTk+XPW8xz8wVr1TLfNReZ1/vn8PRStLfiJbIBSmX4A
2aK5kBSbOWVIkre7Xs09FuszxHsFVy9AOPH6sOMVoJsjkAm/O0MLRlJ0rTVY
K1pHmWrfWFZE328qS0y7EEFQyJyay7Sqh488ZcOPdTbh8BHEvP/MZIYp8k2E
n9/cMXevNGMQC4a2thprleJQy0pLMycaRItejJmVVoP6zIcT/k7XRtBF7YFv
g0GM4QvCCRtAmRCyKvDRQjdzX4FYKUQ618vvZ+HURwdKhDBS1cbz5XwPOtOI
MyXr16WMNJXxQpCEIzbyQ8cawh0RRXc03dZCjp57UrlVHLkkwjWuRr5KFTBV
OSaxDDF5cwOgGeajFiiAN/NCjQyEf5Rqt6pUq57Fnh90eMo3ZwcBN8afbY8U
tfXLJc9OiHj6kvnjIOQrh2PRY7HfsnLMqoOXuErDAqyfn+TJBqOJ5JobqDM9
Vcvsd23gwZU5fNxU8QpJxJlYD5q9ECh87jxrXJduh7ab33P5tcLXVjohHvUm
zSUbDuTrgpF17WbP0DnbFgwBTwJ0z5ubkX5V0JbZ/MFUH35cdOSxjhRQUAI4
jFId/QViyZ+TwlcoMTQqiBXtxds+/21C96OcVJ/ntcKhjnvFJCHpaPXE+ZLa
+5TBj7pn2GLN0cWeko6LD27HiTRl9wCJd36R9ZLi812TaS2MscMbcSFPUle9
gcIqqoAzQGipHuNINlMnu7mxxfxP7nTl9pliJAkQd9dGGPUv5xgV+xu7aqHs
5KfQw+m8NhyxNAiHGkaL5n3tH3j7w1y//uZ4EEEgkaFBe4axBgqDodmuj9zU
FK3589qxecZY6hXNnLJVba67NYMFsRPnaaOhFRX4VMdX7Dgk+Joz4l7KLT8R
g71FtPz5lPsd/Z9MXDI+PP/zarXT8FtGbDfr4D/+dDFXCJ6Ae2hmlXkIC/WM
0MvzvHxFWkGFr9kI77CSMz9a5aDEUJPar71jCIoWfMoLeqiuCRtwxAhkf/G3
Z9cuQYcOq5n2Bl/Kxmcj0L3Agd6lbIoRei7/2/TiWY0l82SUq85aoxv5IkPZ
jwe3mLgS18LFtcRC6w+06T7AVCq7HRpSf+YBv5D9TCgbCg9QAZKlyoe10All
1yQxty9FJ5eMn7ssJ2xZObYK6B1KYoFjzVz6HkfW9H7WauHKnIYlf0jgTeAf
n9gmqXj4CGtTyvqyAXuBGl44m4wDQcNdogQ5Ej3qA2Z77+KjxvFgFsDX0ZGm
yUmCM0zZKPGMux+q5PWA4JIRjBC5K1f1fHzrbanyReMOC+djAvbOWtggKfo2
dKFZCicjHU5Sj+LeW8/truYX3UiJjoYzi3dauYCkL7mjSn8bUBfRBZvgv0d7
aRzJ1pyhpPv78D8Bs2T9x+cFaYRfq0t0vhJeKRI2Zaj0j70gSt6CYjuu7xWy
ilIXKoG411DtTioUW03Co1Hch3CVaRthkCn9QSIMJpmU4MZ/hY4BincBFNkh
9Jqf3ZcSuKVrkKNRimIzz62ST0adszxs1sqUWOqGUU5WkDJt5jCNTh9v+g7l
KfLzkGFfdBtnR/CCcvtNoZQAP9ShvA+Hi687xUD5VQsrsb6WYS69vzpL+aCB
nKKl5obN/QbQL4BKnlayms9k6oQvTRBKkKjTsx2ZRO5UWTctReULA2qVNkct
WsPjJwxJ670G7R/wFPyzjbZPNox9Gt3ZDL28dBFJT+3UnOhjSGTFBiuJvSJV
0HGORQQCgaiv4UkXBWZCzwAc9z5pHDuQkNOdDhA5ZfpjuG1ljmx1u8uVWtws
R0wfuUmYhpmIAak46NHAED60GsYKZL4ETCTyyWYNZblmCWfqfZjBoqiyMoWk
3EUzYK0G9OB/GQQ+555IUBasx8Tzydna7dXLmfd4QbCaoAZn6y9a7PiiXG6a
MpU4smPEqZN2b8kK4o/mRb2FSuCTUE3qvguJ5NM6Zh3bYfmtVMJPP0apLJn1
VqE4Tpw9nLQt79DNRYTIFB0Ec6sMsIiqHrokB3jqSueXREo451WXz7BLnk7w
LVZI3KkTexx8ZzgjnGmfO/wCgZhQoIHDU65aq1VgW19K1GFcOj7Jr1J2N3lQ
fNQtxhs7qmUNUPcz4qM9rFmndASM01y8t5jJXE1MXIIQ5B8rhGG05NfQ8smL
w5sK0mnlz6hylzYxTRCJoOteF40CwbYx4VmN1ikPv8CX66Ve2QxKS54SeHRl
h6S2PBrUwWpgkbPWABt0nra3bLhAOWOylafdjSGKS33fgzt3RGTSssgGcToK
ZbgwM+WpYGzc3zwZ79PaiecogjzEEJytu6YeVFArjO6ATH9oq1FItAcEeZUu
wKdkuwAUn50Az9UUAAEIcSRvLT33QC0KYsGhN+et2vUGGZOx/vkHOOQ6/b0m
yU/hyH8gNWqhPzS3lHE1+KeaGemIDQAei0hxNFo6GfaQg3DaZg1dJpVzZHo8
Ykplt5bYMDbaJHdxwOxJ8SKhSSC5ff5JzQc9bgPVDq49yMsZ9Lm7VRnXmVKg
U4Xb4vYovx2qa6jNtvmYSPf5kO4uBxq6SDuBR9rc86RoUR4JFv1WfqP5pKvM
83hWglsz7HSG8vnzrx4jbZYAR6u3khZiIXhOo69xCOE22bwiEfgSnZ5/vr96
BXu0Db6vW4MrHMsf/qhb1Wq0Ze876a+MYghCXduUy0gJv3zvh1VoViBF5OZs
ToG4KraY8u9JryYETVFQbnFE8aobyfqg+ouvuPayCltP0mLE5GzIAYXx6hph
IJBuRPB++3G5373s8FP8Y/Q1nNN2IezjOTL88kr/6ook5Xzqi6Q4SEEjHzbx
0WjieZHHDi/oxSuCxA49zMRf3zivSmp8emoq7EkSSh57ezo6QnDDV/Lz2DQx
ThKnK+TsZNU0WhMnjPAIDgMbpwmOO+L+UlHQAJxWs/2hke30/bepyxbaTJHc
8ZUmvZVn8E1PV/SscTrOACVA9V4S+buGX5c5p9XN4SlwN8qxphC1TtZy+yci
fB4bhwW7ofcNmIn4IJLjQIF12aqDOj6eoK5HxHpDJDev35sZY0mL7NcT3oVj
MIdYTL4If9RJsHfRAwLRRRLQPzRo/Pmf9CCCn465BwtZkNsa9XjVcN9ChL3g
gKZsFdvStfRRN9AYbxiNKIUZBg/dL1bje259F7JnCNRR242uPW1y1qPQLIYz
ek6evUjP7gMWXDukMzY4GpFN3MJ0SH2sj0XSoL5pKf3yEss/muOmAL2iXwIQ
MjEJBbRiVWImafJE5ZuewDMOdnx94AD+eb01pKxEnoQZcagylf2qH+tgbCc+
z/XRI7pznM6b3wDjOdubB89/WTJgquOaj5OFRZRwbujhDrGCiRxDemPWDfc/
N0KSu4hV6ID9zeYMLKn+gKOe/8H1xIpw/SadkI3CzwBZT65zozZLTNttkNkS
njPIbc/IeCfrjIa7vT/YEFq/zQ6oWVNZjZv2xjAjw9YivFN4MKbtLChpJ3JO
bhNH6WlGsgByOHmgXs9VVLalk0hW6U757e+F6pI4hBQ5iQAdxgwR35JMumFT
WMvnrFH24n5XiItHnm+jkNW7cuuxkjlH5/Ep+9ZwnZto9uA5crREaLHV73ze
M7Avdt6q/RUdTW1eXcDYkZzQKotCIdU0AiLnBarYuveHOKOAP/fGTSV/5Ks/
XUzJjzDvwtzmfqQk87paNC/hK1jnmaF5P/Y/tFATwESnyjtnoOKrALT8ixwN
Ip26GaBwQWEb3u//78pYxJQhWSmqOnX8TzL9DAv9i/i9E5OGu5bNZR2twq7V
JxBsBXrjqXwB6CK5bB56fNEuMpMsUfkrztTS1c8IVyVNJ52wnQr90IJUPKOm
pJFWd/E741J97Bzqd4ASPj4+bYnHuE+v27WfpaRO9OL6Jegjf5r+WK0N05oD
vxX9vb985TlGSx7gMji7UPR3u3jyr+Fiqzg6rCMlfmLIHxbVYQDb7N5/w6eY
gokdWi/fpuDxaZCrqXo6d5K4v0jkUGjwcB4HDgwuz87wq+LmhEJquteZWVPN
IV0TuQepVzicSOKDrvKHLlPiLldp47dX4oRalfg5b82wlwr1mhxwirPHL7AF
zywtHtNcDGF2KTNaagDOCwN0XeNTWB6GENH69gWUd+L3MJStGZr11E1umsoE
E/AXvfpXbgE9gpwiHKt2CEFwecjCXPqhD5WX7SNul7yyVNYdrPeGWAVO5CyM
i/tLz7m8cXbC6rgT06xKEm47vyAWX1xtaPmcQ21T2CVwgZMECg1lwBl9yXTn
cXt4CRFcZfybW+b3J1gqFrydRmZrmCdX2yJGTG8UO+ukUDbB4XD7SNiMiqlr
QLQmOzG9MzZq6jta7uK4LihIsCpD6b+MNiroWBfESDhXBl4Y+QdKq14/1Hzu
vTbexWplpbQEiWIltw7gUe+yM1Ur//8mqHMF3ko9vHHesqi/1TYPQt9xL5BC
V9eZCOOKPcPs5rF+CqZ3GaBb+ChhC1CQTqzyi5swBHIu55mIj9q+SN2WbQs9
YrfCW3Fhs5BYp8JFW5/Lrx0KDd+QwQA4ryWFsFovp6WhWRnKXCO0IBW9G6I3
7YJc1IIimg8F5774PNq2skqWgUJdZfPjXFxCdVez0k1mX3jloCJOGRp1TObH
4ccXcmpTrw6LYF98QSsPRs+WKfEEa2uZRoppxnGMTWHTOwFdWMkNQQrYntl/
AGlHiBmU5YgkNYo8zjzuf7QPXNTaSNcDX3T7yNNTY8BbzK72tZ7tKPQEM22D
eYJqPS4NNuZR8Znqh8IanRUiHQqHmjfzqROTyldbiOUUc4uSp0UKKrN/BTtA
uD6SgLRgitdiTUtkHUvFE+4eA6wbJz//Pr4sNqP44B2eTfVoy8ptv/xwdCC8
tWondxi2FZKnEn4qJwoVX+TFer2c57RGSeSSr4CB4GQwajSgEdZJOPPxwMt0
7H5JO7Sqep9ib9p09+Gz0Ggf3zJ1r66b4Nvj7sF1S/A77QvenZJubuyhgAJM
8z8pex67NCQW0ht8se1b2mwgIcjHrcA2o3LYTC1Q+m3lyn0cC9GX9ouoCnlS
mRIQiScRRvPCK3clKVTfeaDz3t90DliqSk8rsqnyT2wFLlOV2mCxLzppPBZI
C9U2czT65ogD7YuVoV1uAKKqW4HSQlu5y2e5Uj6j7j35NcF3cRmHUP7i2gAh
gB2DYLbu+UsEkBWqet/Y8JH3nfYR0H22/rZ+xNTUYaX0ILbzhgP6RTIyer1H
0Wd7uqJeooSEa3/r2RUbjPNtLiBEv0Dg5+dzcDRMxm0Ohoa6GPhwurlxYyyX
35l+8QV3Yey4rFDx3s9MNQpel6eUHA/0n76jQs3yCxRmy34uUYXFw7P+shC0
OF2F7oTFVfoZ03/k520pR08P7/FvXUkkETyCS9CO38jJALqR726ZD/niEFtX
UyiQrq9PkcAUDhhv0j9bIJDv58xFUioF8QstSAn+ypL8D9soWdgNyf6U4oKb
rVDaMXtPoBqSJ6nG8/5Es73CcgKsVGVQM4suzDOs4nGSJ8GAqTEr92Jik4y5
pzhwjuqA5WjvllDIQUkB6BI01KW/Ss2aTOCE4yMsua38DhU1bH8jmD+NdG2C
jExOelF7W4D+P6ftGMv0q1C2Hpx8zd7bJQdbBSySaVOT+U3ddykq2D2nYw2I
Fxt5VOOOYA/Wd8o02nWTiTRVPKsw4HPVHJO2y/tHp/zwOMOpZ6lYj9zSSlHj
zbwE8D79T7bw3o7Du5AD4UvC0k5M1NYtiTXHRmQJ/oEjA5iikJZocpqf9Evk
p9+Lpbq3GG64x2wv4lH20ENL4ZzAnjloKygOkJu4ozMjd/CpX60Y9kxBv3S+
TGgLdK9m77iykotXZI2Ed3u7wHw6/iRUnzOrj3Ep6MHEW5oiCwju6Xdv2726
1fh8RZEFkdCzW/hQ5NIe2OplOBbEL3zaRx+kJXsIS234raspa2iD0tXaoT+y
/KkJtuPWXuNKePWtRlnhPpD/ylJDpYdc/yW1aFruQA5GwN5l5QcviQHhjQ8X
Gh66+5aTULrO0EC9TnTaAig4t/uG1D2g005+EJeJ0QI0UOkk6u1RaIeHPy9v
zVKL1N6HzhJ2GQQvJ5SOoBqyoBYw/cfN3qGfjcyTBNvX5FDj7q2OlpSrG5yp
OdWBP8XEh+uy4zKuKnuN7VRgGd/m7cBFWhAUcJHTFIId2RzEnxDnvKUtDDx3
+JGy5krls4B8ChG0/twY/jFD/lkJklfzbi5Ddp97u5kjg6gDQ3q4vFFdApEv
276+qEnmTSyyT4gDQ7NokkzQ4/JsWenZJ28Eo1R7oeRTCjhKe5TTcBw3DLey
kOSG9nQ5O9su+O3gDKYLnHc6cCLkDuX0WHfYewwRinw1ILWquTWbElRARhLj
HhdGfAu/ue8YKuKFbSwf7TpAOSEejStCHX7gfoAdRhpLjbQuthBKlO7l2zz7
B1xJNkdMNE4Pf8rFAQyhriAw5uSeQRtuqfGwDkcXcsID8pk+SMcPiP0ljonr
U2s5CwsFOlAey092uN1ElF4otix81k981jyahgLK+3w4ZgK1erTOf7d5LaML
lSK2dNQ2VblpV605Hmra1o9UK0YwWWGb75NMDoq27eGlyEgVUboSB6lhoTd6
1ILW7w7qYUWMeQ36E9gCClbFyZw0psoWF2ss2NYKSgMdsY2ACfgVacNG4gUH
CMtErfAu8dnJZZJogdeF8rWXYzQ15lYfeuuJHDn9+9YhXOwZiWD2eCTN0DQ+
5kLweXtIUd1lJ2SiZTtrxvRHxwppZyA1/y2Mdq2cf+0Qt8mLzyKXqXvesjpG
AtFFdxAxcEByLkUbLGMpvG1SrXjZ/XPmW8tuxKnkVviLqHsNV+S5RrIlDFyd
WOeY2e4WXRDRTiadH0n4BLbRcaDnUL8RAk76sXNobXLWeH0RheH7hvYOfiHh
TUbUiuPnT14M1EmddYIV7XA5xVR+Tfs/g6QJox2LArD832kH+kardJde6SUz
K5Cl51MkYkUfI2GKN2XTA8e1GZdj5ryh/hBX5xcasKZ6Sz3d+CCKQLjwdad7
5muy756TMNdXrUcd8Q9DbJH1kzA76QX4y8Iq+02O6OfcH7eD8QGCbtcc8Ten
gAA2ViohdE9+3KMn4lEA2D5vrGgUCJos5Jhsuhn3sUFtPYukljjSrVnFuKR+
P1/fKny2XxwFBcYCAq+43TQFYijjHqjpJJHC8s0IU4TsZ33GMKNVgefNZFKR
cxFoS9ulBu22vXyk8d9q1TixTllSZ0qLb7xniiF8jm4V+QVSQyxmUSVrVyTh
pIXuWjl25Yj/3IgTz4tE3CFX992IOM4Ng3rdvHAOvGdDM/nmFsBiGLVpv9/C
56KxcDRATFTMM2PJ1yISaT5jXd5XVRCDBwiEe4pl2aY87iGULkgC0EW7GX+b
hsCMofF7kpCt9dhRoL2vCUvY5L89wpnAC7129pQd+leC6QdDUqBNZnRkqA+7
lbpQaxagEXTmYKD4CxM1kx5yf75IxV5qn4oHusmga2pEdj7N6zqJp8nTxmCk
ubH0V2C05Ky/EpzG/HVlzuHiMChsKMUVFsW7heYqaVWLTjYlPFpxe8w2R9Ub
JoorrHCpvedAx23Pb4aTYfpKN7MBePTFE0pVflixPKqsgQ+c0hxURn3VSW94
lDmNJ7S5YWs02eZK9iMphRwKcVnrubKSWkk03MiZROPUdG2kn6g8+n1iKLlv
P5FzQQSHRhFAPWR2i0uLmHVvzOSs1xRJCbig7hTBl1Ko9SulckpgbegZr6ub
DpV4HALGrauMXiMliqLSN3Pe9JWgNOEHZWRR1QMyc1iz8UZuRpExEBeKDNYd
boDcueIJs7GzHgk9nx4BxQKbB+Ljt+bQDChTWJ8uFsQVgPX7T/sf/kyTjZMP
fIU5HWmMsy6aCFOp+cklJSd4MUgUf5j3tT4XZ7L8gshXhLUEK4HS6AnCRvQM
cS0obZMTKE2XTRuTcqNTgv6rEHAj+58KkfnRq2vycpsN6qAgVchU1ncNJ/hg
7hZ1hogx9TxocUk22ZkyaU+63KYgi3pavsIs7Hib3RhWJ0f8/5rrad0ZZFG1
yy+RTKyWKDgH9HKIIkX1rMeUuJXfuzfTO0lejfdagftosIEr2US5a18vPYFU
7FioLFWKjWZk9QBUJ3/3ZR/uQJq5JzQy7/K2h7hTalWpB0aLG7bfw/pd2qnZ
qg5356ZiFbqFL53Mty3F7OghzjCU11Rr7BML4TNoFle8rrrLddRc6pQNfFw7
BbzqeVlpwqclR7CK9W93K0x9dUQ5tmf0Zx+B8sS6zIcyfcy8wnW+3HXcpxNk
xYKn0grhSxQIzChpuVD3yIOcGR8yGap70/Rrvt/VoZt5kefJ1L/n+CS5aoBy
wxoSEFHfVg0Q3+xAPiGwKO6PsLzdl9HdB5Pn9z8BHRjiBrGqVu/KnV7Ei418
W/qdd4ZSh24MhAG0JLv79EhnDOP+gmMmJ8QOwjLzHYKGs21JRmfqyPH3toPA
bVicxvHKr4BV8ireyd+GvAnHgfasIbB2smjdlsweKK6Ptcoou/m8MbSY80sw
wQqFl9wYye2iokAfE2NAFSWHsDujju9KLvByf/aSvEbbnItCXE1Mj45Ixl2A
tLCx21vz6EcCvx5SzFghEHa/ghsetyDeTA+kHxSTrOaq7g3PmOF6EE9L20xp
9pnNx3DNUGHY+eNO/982d7HCLpT8aBn+Ev2NNW9p0WlHQKGtv21IH8uw1uEM
2tZLiq3Z4xZxVyV3xya+UDWSWjEq03vwBkTfMhPGWGXoAiI+as1nIqiqFIRI
pBedazs0xBPjD6Zrc5oXo9DXxGXtjWt8rRgrgYrjMxu6qrqSSSJqWMcow9S+
t6h5xiNlJNZQgT7D628mlKQn8795EC20Ytp5J6qKc0WtIR1vTUtauAhiR5Ot
dgtdgzQBCElcx/z0Oa0wcHeBzrS9QJQ6ECQsq5AJgit3lVWvlImfodars637
0xVTpD4BYk6JV6i9sC7lwpT33TgXqvCH6D3BV5yCZrKuFZ1rAlF9n2Lue6oV
+J76H3BZjmxc2VQVreX3vGu1xLRTfJ30UygoAn+tP/pOZtmcBzGrVrem1C3O
XR+lZ4uH3kudGYv9Oni7u79Rrh+HowKnZ553Iv6dfheg4DKSnEceIU1Vgm6r
15UjhhAaKEKx3oT1ZhFGZsb/9ejrmYjIz3pZH9bGGt1PQr001lppNlP7lhyQ
M/ME5Go2wJ03PsYZqBKTYBlpMLJkdQUO6JP88TS0S2M+NGGpw/krO9478Zoj
lmLY8iY8SdHV9mqV27mLpy/AorJDbG5sOFVvuzpKYCXK8oqPIETqEBYa05ep
ZsNpjzg5qZd9O/J5PqlogeVTVii7v7TJVK40NYOK57jfInxoOQ+1qlmJkW0F
w3maJ8SigpTrzcAbP/+BexCmkBYjHVs9K/1zV0xjCpZXT4cpxGJRFi5v0Dkd
XySqLJjBi5tP7PdTQQQ+Pl1TG2QKAa7d+SzcH7trOViwGjvkbiiXZC77nZAX
6E3JQCCnHB/tH98hFmb40X9jgmzzYHp8tFLWXrYXYCs1XhL6/AE5bfGJXkml
6ZCVngNOiqSMGl3mgvLaEIh6gL+mw+iEwHsxB26gAHUUEZfdhW+5oZbe6pI6
JO5TMUKRvuS3Xy/okAd2sBQc5ZyRmnFFLi4wWiLvAdapuTxgibLHv+jTDuWx
PfvASHRHR8X8NH+AVkdqlN7Qw4B1kUElZ2V0lv8KS4JoDWGGyqffUJljMLN1
QT7qHvuP0d0VMoxy6kCVWo4n325EbxjM+Qi5fVac5vJhj0Cww8OrRQVdFonC
0kwowwSMa9IZ+seVbNClKtM8VlkPp/ESCkJxZ2mnt8hNb+a41SJaHTVJpuEx
fqTT93I1ALyQe//Sor48pnPSWw7k81e6fE+Orsfzt4h5EWpoq4oP4/xyQ8Es
4fGVldzlCCJZt9Fx366LeZiX61fZSn3UQF6yiB08V9EuGdzKbuRt31w1pKju
RWJUJZJmSn5F8aCiLaoDWKSNjV6vNzxY36ifrZaPagFPszAF6ZetSOQ+e9HD
ueIXSiJLBFyLul8/sOcM/qS79OwTbuWyNg7ULIJfQNyAMCGdBh854uhZXgZV
OkWbc1JF1zm2PTLPJTX4wn8HZSEsbEAm9DHGhV6c8pvuIp2FbtwrhND4qDTH
N40sbkVWqQfATn42VuAKoMg2EPueFc1a6ermmlo/b/3Ea6E72Guo5lKP9MoP
UYPQb/qMOBjROOFFCR5WUzsxO+oha938Ef9lUW9wYqlWqZH/gi9tmq/QaWpO
xzPwd96fXhVOYyhPp5UKqcWDAKtI+wCZzqhZzEJo7dnbfUuo5ZC012bunN0k
13Z0ealopDcI6xoO05KqInwlv1qIbn6aGDFYI9dSiI9akTNFBJ0rtoUEwuSb
L20hOKcTCNhrav0I76TEbAPCowPhjD7gNBfj8dBTzASFX3laYi18Fr9RoNSg
ADPt6nkTIgtM9CfBfAN+vgBaaxQn8SRqqFjO58MSYFQESDv2RDMInuG5uVWS
VnxadQk+8/66ueZrqDHVSmsa9P4ev8dzYnCmnOafcWfBAVbBJdKqJOi5Xkhw
/arPMEzn3Tqml1myJIXAKuXFfcWu5ptj0VCMv6vHYE+6HymfzMEuMYpWXeJJ
N99ZFRyukjKDOyxlL7Q2tWJyuIFpnkbt1516A3hkWzUZAr30+5bMkJQCoNOO
RH/GV6KoV0qbopvF6yIPCjBEEL4aXCORz8UQLJXYJqFB4LGuswUp8NV1T5yt
Teok7VMI6ICLNOSZudHam8BQrxlPsQE9ddT6eRdzc0OyvLgqKbTCbjRzgPlW
UtK+LWdkYuOJYijSfDvTXbrvfefZAwYJe46wm3roH2qh6D/adHDetqM1UZ4q
6w1HZIGBaeqNlw3EdNjJ+una8imwxxaQ9mTnpQ+/pJBaStOGgmhqQwCs7Ts0
ZtDRi+QpAMCspnxrZeCdIqVfyuCwyFzq0Zp2xndwPCJvf0HADTpIR4fZFxK9
5mUQalkJYGRpzMnyRhGFiEAjAmU8cwuZf2XWukS2eWiRTHI0qwVLIZjmZUeT
MO2gc7SHLVLd2WZzgT1qViVZcHbmgkV8NqqkBPIZbuLstMSK5mVPdSydCeri
N8kZsuyaGxmvZRk9xhcQxjS7iYT9hpPnAP6M56JU0glGC6tL2hmpJ9nYud3E
JkPRCKrgFFcNiQVNIeqru7JAd19D3fR0ix6n7GB7ms8w7PehfpZpjIERmqt+
VjWoR3cpfhmuJTnhIXWkyRYf+u6mjc7aoleY3f9ZFR0c5x92iqIQazXNDlin
OVXGu2FQv/C0lMtbk4COEpaT/B0hWnQjfYLhSjJM3Mi7Q/ld43TyTiKyzMqz
WsQAWsueJDEQVhtplqFrZwTiu9u1qJIRcrKnG1TfGRqyGe8qZRmRrubvJai6
FQlk8NlhXTW3UI5domf/VHKMzlZksuYNqAqIcYV0bfeCydO3WoeWDKCSUnxB
xG/nAHpyOYtZeuTcbcODoxMQtO+GzkQ37VSou6lPLy2IaHBYoh0cH59bTtOI
ohyVWXVXloc9m/gBv+IicPdG9qopggkn4Uut+Z0zihRlL3KVK09IDvsK2+r/
hGQW+ceYnkeE+zcZeoEx7/uaAuA1QjwoxMrbu0z/8Gg2WGPFLB68Er4bgS95
bmC8b5cwYZHhcPWgdALkN33MWe9I+kAjHiO+E9BRVb2AZ5zWYm7+HV1qe9VB
gEdztDGlGEro0pvRDEjpiwkNCbKPs+prlPjrftfqqIQGL25fjvXAEXkpwzTI
ylw7xisOd7suTYgQT9NrgJ9P/992VU7BcRDM1Mgk6PZ5K75/vZbHyFzy0buE
7M3rEice7QNGYgmlOyW70LpL6pGObSszRMu00hARGqCAruJg8swMchjxVYvS
4KGCm239sb9Vetooe82ZhDGq42J6tYELGVEWDXr1fLFdzdwmHpm3ynhtjW2x
7O1KAov44lsdrNRTyiMhqwN/tnADFehTOLUMSEP1Ux0li+lKCDkVuF0YBtX9
9sOSVtFJsnsCJ47SUybN/APiViGJ22FNU6FJ5Uv91Ch/2FJBdYDCobSD6IAW
eCZBqwfy5TyBzOKp0l0E2QZqRgaS3DtFBNhKc8tim5ZDNu91R+k4pOKLPxFi
FnMiRriSZWmEVKnX5Z2VeG4sRx0FjXvOzWIiJhlwZBPmTaip6BnHhSPLxaP4
Vh3T4tvh7LI/XmyJKK89c9eF+wXwl+ZHW0d+6B8yNyrDADPz7ycRvdbKmzal
Q3PB2yNWJy+pdUxGs3lXJ6TE2UYrobEXaSKNzjtlA/VD+y/RVMLuDAB7+Ebh
DNpl5N0y346TvPO4CZm/au/5QzOIloomHMT9Jv7uo0Q+fOO0KPGgdYINo8Gj
6gqfeuU8+HVSCV0KbBgs1C3L67Gi9MMp7igT3nkmPtHx8IXUYHKuAIYpgjDh
8/0I/QqKWTpZ/HetYxHdUTVLs0AyIvoL0oyNOvllBsZsKzkgRpvkyfN9W0LA
5QNTiemSES53oci22QYkdcZhG7r/zUJcN3PD926a6W4/w+zoO60F1wliRsSv
F7wQ9dn++81FwMgaOxiMvRF6XNRpopKW6oYzkPnIWEGGnID/NV9Ux+2cAktb
RHcu8TKRlUl3H6VzWwOoIL/6usHpzFCFzi/YjvLwDYEJEo9Fa5imcrq1smBX
6d5AZfQRulw+rCJuOGMcTAca70j6gCagdEX7ipR0fYmcvJxlWvJZ/zu1xeGW
2eawJpC+i6Oz87PRSLeKUilxrbxpyp+0fORTznxo+e6ROwAe3wiMgEEws6Mt
QMhTP5YkAfdVjpOyvZmUcw0pQrPBGTaYGJT65ivrr3tlm3bVuVlADrz7Xhx8
fsNlEJg3I1QOb21D+9YulXtCim0Nt1F4aKlo8KxwDK5k4sQAY9NAIu0nzMvc
0edV+jX/2j38AsPsOaHpkKjl6R8XAdtyesPXofJKf2gGd51l+cxd/W0uymW4
6fBEZGO7g7mu1SKrCPCgAbExmWE9XJgskn77px8Y/Ujpe8HJj3iEUpYAwFFe
MV9BZ9hFzqrR53euQGelh8G2QnXJ3GZoWPrJWwNwF1K8Geh/94wynwyOZVgj
pAZyv2vPpYFZNb+ksmOc/fwOILoWPnqjt6H6qXUHTrP9ZD4PsEn60lr1dtrj
1bBAE8Is1X87fg1bFrdhXQuG3vES2hUW9X4IwtY1b8ZGuf9wjeTF7X904cAr
hrziqrsUK38AsORVkO+zBKh0y8UgNliOIujJVvHTxP//ZligACcp56nDcg95
/ASgJJqg17eJ+s1/LIGxVsObwkEYPUyS0eEuVn9z8pqvFl5EqpDtAddf6N8e
GI25/6FwlHkSuwt+f01f4wmmnyPdpjk3VGqEVUuV1h11QIjXezX0g04ZRGSE
WqCRwNJWnCYCM0Tj7K350C4qq/b8g8nalAEFEO12kJWsRJtqESyXdvpRiBRR
e6zTgMtxQkEx+0PyOOaqWRlU6LreDHHpuZnzMrCSrKI6rn3WzM4AqZySFgNQ
PC9u1+WyIn40wlKHb1Oc7CnlS0MHIWS4L8UgElWNcU8l2Ex6cKbakdHwzsKa
sPgd3OGtWLxB3vm4EvJaCFHgeTprRUuEzhWO/eu25LbKa9rce7cEZRhldjaZ
AK/6WXUacMAO2sSxFgFZ1I7RJ/DpXXbmPilq8H8sPg9zOZ+Twij2dG/T+gp1
XP80uffDo/KIX437OBf/Q7NwkMCPKJXi2S0CoUL/u7miB6b3DrDFI0WNmYtu
APfMw3rOYY/dGtStIVokrnqDOpME9supc3ZSb2nI5dMXonu6JJIOW9hTtKRY
OELKFUpzGW1kA8EzwdouOXiVQP0z0BVDhiX8d/5EjCZMNduLzT2uR4AaJyqW
q0e+1QE2aEFVR0x0FfHsnaKEUamUu1AYFJETxx4LBnEJNnyRjiITVRG5MHJ+
8UPz6Lfk6n+JCUZjNIo13xpVqpj7csrRIhIVggKsOWa7vR47Ufikh/vcMPg+
36oQApgXBedIfgTan3tM2n3HbJAmiZn5hyC98QX0PTzvMvkii8QOZdR6Z3NM
LLzCLQWJDTZUbU76U2DOqVYj9NfB7Ps2HVA4yzN6CrF8qoHR38/sb1fZ6lUp
o2hpmAgSfMvQt3yAafTXSFlhnDVhF8pgLPNVaEOGRWOceXWw3WusvYlrG5HE
PaUTtVTcY7Ur5lwYxuIL6rGIYQZzvHCN3Pk7TGI5+D5mjUoQjuYGZozgnv3E
XLCdqYSRA6woeuqfxhPyKVQdeXibQox+Um5hEaSfENcBWJOUhNrt98UXiWPM
jOZL6qLaJPR0/uL3zkpY9gm145ulIVmAkKYxAbLpl3fbs495LOLflPJVusnd
VUATosO9UZW6ghJ0H/6qvtmsFIE3vJamFron6Bf9rtIyycMWbYjkbIN9MBUN
6rW0YlkKrcSqQ3Zr9JLZ7hSOCl6nQNw4DB8+NazIIXobpUjcpkFVcv+g5+qB
WBJX/wg8FFHUzXoH3T+dKWEYzpb8N7v6zA/QVOeilmOlA7GhImifN1kSFPr4
8zOdzjN574FoLV4Jsknr9fp0G0KJxke6GP82Nrj8UX2+zt0BtgQ0wap13TMH
Zy62dRQJ3pjp11Y6QTmnomRzZTpa46Jb9krD+mGlQ3j/isSRXoROgBMSKKl3
zXsVSzEUFbwrRdBmjGFswE3I7C3WQGQ+/tOLU5x7R9w0CjkFysdeQyEzsApT
qJaJpmqSY27JD4PzyNyr0eHArbKY9/jm+rnKVoV/45z1FFPYzIshPyRfq6GI
0i9OF2gCRRRp/f8s9U3oVHX85z8jY1WKFm26mwoepb9H1uxCYW7aH2DbwFy2
vUZi9vjnCVLSS/9tuPh6RyCVtWCARNBcFAuqcGPxBpRohTA8e/JidKyqTvo9
Iap0B7he1+yx/BY90g75WO+HpnHtmgLMTwi5kCqtLNIQKnTLm8r5Nh6pqQ28
RlVf2wqncRUTQdmzbmqTsNYhdaKBGhHoMf5dlhEnebaeVOb8zCCfYegKedqW
JCA5XUj+XxgachahUZ03xRlVvyCX2n5Vxjwu+aMF9XV0XAXP9JOqevhNedP4
h9jGiOkoI//4K2jI4VH0DVHAu9BDBStPqtvc8QqVRU6FCDqqB7vAfnGBU5RT
HHeHp7TfmHDAcgccDhjQmwFL/uVQle3C5WmDfK4hSs2KNXEvDnRiR8+hVZNO
7KrSJwxx0CwD0FzUs+g9rd4OzuLOrIunh0+jrcq4uuypQuCwszk3nelRU68c
EOlqkZouhezN7kS1wbjymxwEAiR97M537RoXW7VCBGOQ0kOtu9wUWQXHRNqI
2mJrA28+JYR4qWyFZq+/NzWx/6gzadWC810z+v9fYnngijF5gFsfCSYoCuqs
+VgoIUaob91yy3tpsexFSt2jzsMVDyAJF1FgDMRK83othG8vdFLYuVnLTW9u
qfVXzqjjw1ZoNs9rqjg77/gKEewXDo66GOpzDcb7ldQ1TuDsrEP5cqb1i72X
W8OXBgxkRhfG93v7s9L9JcNV0vphDGfMNCpW+2PAVwyQ4iVF7tW6u8WmRGBn
6rMSea2uqxNiOQfv2WlcIN/O5f+10Hy3eIurrapRNGxS1p7GcKxclekQ5j7B
6/r0l87phryWiKdVRNsosyuwdDjZPhHEYRVk0rO1V4ZQFHwwdPly0nFVR6/S
kezZNsDprODJGz6IDGxuzPKRhEYJ+bo4J4n9h0x9MhGaTd+2eTpxWxy7Shex
X4Zw1t+OpM8TjLpQKHYAiHRLQ9/rd2z+wQ8ncyxr+r4SV6h80DuncuZ6wOan
oOL51fWo1VkMIRjZ2/D8pGT23osKTWjXAvPjvH32aR802J6vJsIKSlJVycOC
x9ad2EvBqTkhioGsGbVFaQRwGFCDcX0SiG+uzHUPU6EX3IkrN26Fj/d50f7C
qkRl/ydp1Vw33O/C3y3+JQk+fixxjT3L459YBz+XifXLhfLFx+x6VeEw63Ry
1MlyYY3QTlKS0YWa9ie0LoeFIOpw76vvdfCDNmXSo25Se3o7FspMJfz1QTba
GezlJeVRIazYNzHSreCNfaRHn8LQrIclR/K9acjOTrL58dXUr+RkrlMIAt4e
d3Bl/dsTMACNyaGZrGUUS8KvAls9aFVv02h8ozpTTdwYeHwZmSHkSFXJRggU
1qznwkwIxA3IEAv/Rv8b51COdvCfmsDD4zngPCgN0+0rjPSqYIxPZIZ/hvlC
K4EH6wL7rZ2hSrszklTq+LSb/66pk+Z11NI6Tl0f2dpXyCNeyicWwbdtmFZl
gIIDM9z9gArDOX5b99k1s1VHN483mLPOAKg1aiJJDe7aAn340qtYF7W04tT8
EzcA2dO4LNzf66LET7WqHTzobkqZ2nI8J2znxfx33J10wKyXoO5yG8Cabx1r
xPb8BxSntjGKPcyfbL7CcTsVP25AW6mQ3AJECSoT03WYeKahbUXoGB0ZgFNn
1GEMtKkYMGsMi/ipjZCb7Rcb6tJBhCoBF8F4uzweLHWwdOY+U4w4g4xVoFAS
ldqeA8GtZ5LLYtSZp0a1/0ArfwyfUug4jvSE27Td2+cAFoAZomWRA5AahmfC
+KohgU8iiyirNj9PUErJPO5nBjE5YfUXJYEW/fH3lUylVdtylmtVi2tNvaOi
gc4RQkxsCxJ6BCR23vfLhDE0n/aElwCIRpde+tEzyPK3eO6osUENbz3C15LQ
2MJIc/Ert/WxVS3jUbKb0NGR6wMJQvKfb2VChxAJJ8afiklSn6+dUIjcwWLF
0j/adOB9dAy30O3aVEK2cQdZWj+SHohBCk42ahp9QDiZ6/Ht/gg+EKH2z0/a
tkvW1WU3VHW3kU7LcsAK7FLKixuI69CamyIiuNQtFnBDP1TE98OchHiPAxqo
uWoZVJn4v8oOAfYbBNiSTQTehGjrhzD/NhT3mkPArYGQZkwh7LyWkqNtyLaa
9Wc+5j6u6MyfhTR7GwDACQVur45BpUh54xOHxbe6bJnl4GGYnbxGhRV2Kylg
++29fbk/OoF8Phe1pXdm0QTViqerfW7niSbdJuu51om+KJMcWPKHMXWrDb6B
InVTQMcBKUmEBPqf8BRP9MQj15L3WJZ+Rmee0IvG3nwOeto0t9rm90BtXrLa
299UP7NcEttTXqv+OV+5T/BX+1KySIzMroOoSVhcIMP+G/N3FyWk+zMzi7Ol
woxMrpcxgwa59cVEhqoa8ulQ0tCOIjD41CKgiLavs7BKB7CfveQcZRkPDLDk
9/O/Vkxex15lbna1cUxX0azO3x+i+EWTCSAjpU+kw+Q89u79QO+PdrbV9uqu
AnMWGrOjdLZONRRbTReQvzHkjkdTEh60fm/Dxeamq3Jub1VllN/fso2Wjrrz
jD7qNgrmqbV8hVmwKpOJilh2T3J6A6CTw7229ZkoAwAn564X1QXqTTk9bh4p
+aP2ofHZuiBJYkbYAgdClG9YrkglgN6p8Iuex9NnJWUJKgAKE5uZoIPGtm8X
pna/9sBbwTIpocgixrBaWf2F+SVj37oQnWZOm+/NifbCEFh46maGIQf5yz6X
xrF0RJGC0HyZ8UFEaqzq1dXkpZeJPjLNtBH7BFUvT4p6Gc7NtWCIboXRcOwi
3KePUPjrLw9JjxfXh49ZJ2TE34kXVkLpBUR2Y4VoeyGUlfrQUTh2GVjeBEuH
6rbyD7KqzDbMJ620Qh7IbRnBeYdb+pAXlE461X3GiSMfMe/fh9wsVM2+ZuZA
tpLJC7yDTMYP739kZDzuX2/EW/o5ALnkXtoLZuY22oHKQeY856+sbmQ11x8I
PmbbTx8ukO7Ar5vGEDEpP5hSYPsjeqzg4cWOVuwkgjR3Ap+AkSF1/wQtYrHx
XOA7UtLSdkcL32+yBiF8bh6bKBbnhaw7AOT0P+JI987s866fa2OGUhDVz8PN
d5uaAt8Lpn6giXgAHyCg+WdThED94xkt77svAPSDzdWMauSQuGx2z/FIWvqG
q0Dma9++cl8/c0XllI6Pk6+spb0idTRuv4LajOYdmqRMRvCEQOz2zABA+x7K
R8JNU9L5o01cZyXqkk5dlDSBRuN8+n5kdnTkRLIyTqa7PdNUqcbnEUwSEOz9
TaRZgLCbCWjDkVOJ/EyQxnW8FXnhkZdUpoZmgDRcLkWrtNIbiTUSYSdCa/ld
bRTTagoTpK+F7QNo9esRdOryLxkzyDYSO+UJ8tuBd9Q37hwm1LPZp10Aoq1R
vUy+yWi2DTKx8+1VQErBSYFixNQWHPzmrjjxd0UqeRhvQTuDXsJAwd+OEqlI
kOgVw2NdGm/EuDPVD/hBr4OlOYQVUWYGmyalCpjFVzyvg86wXBK2N4ycTgj1
gPDc8q9Au9pnpbv73CUAj1p3E6baSEj+lOJGVMu0VWnV379F0ApKDJbWhn+c
5PnIZfcT4XvXIEKMIwpZCnUYnl9Nps12FLxz8z7IqO+Wz7Dw9gAJJe20s35e
at0HSq+Dc3FjmVL9CP2+WpAb3PbSnTCePz6vRL6+CqDaBeZVK51vINZc5EFa
S/0e9wH/pLY7Z1b2BBuqqTbbCCkirndeMwFSQtx2FEZeIbtbPEZ6oyqnZdcf
g20IQDHA4sfEIB4uO7qV7drn0wh9lPOwMZK9SRNsw+ZTcCkXbVAvUInCmTRJ
IgNJAdWCdzSBpUrCqx0K2n3jd0zYgFmuvLtcInbiimexukImDh9/jmXPhIxP
BLqPh+5hARWr0JQb85S8RYuDDrnxGalGrDKEXE0j3vWfg4GNuQLFMFpQ+DuC
TTgQ4bkRFKNcDjWDikzLJtOkYDqiuzlW243OHuF83giZLzWzk1W58W92n4nl
pIleNLsYZst4sgMtVMClchaZxsYmwCLV83BV/eAVQkVkyIpx4y15EsXq1VYi
T9xdmxPFIId/s9LEGTWkgD5Zvs1TyW7Z0SQ4PoNAG1p7T8n3BBgmkUpTMUGu
RUe/XA7kXMpVv9sF9Jqfyt68DCDkviJre5w+WvrkX9GjqWuX9FwU7kIAXjWs
M7j1wrPVEFXuT5rZcqqrpG/cxb+DZpv9KdnYbPYGv9bfuTZa+3eBacXcM3kT
X8p/2tRLvaPIttULsA8rzsUg4TeftdvDSwtJCwTAAvy9EmcXSI+UsY5Y3UvL
QY3jQ2OvuZ64oYJoOar0a7XDvuADLAwZsuGmxVHAL7uFXlZQOIG1HLtjANXJ
QxxdvLvjzkZvwB/o2s1EEcqls/x+CscSApBR7SrANPli92ekCmw+bO3sLA7F
eWkobDaJ4ZnOmbOW/QyvSZ28/7J361u3Daio0HsyKg+OVgK/j9E5RjD4hbAk
eS5FVm5BhF1aOp8A+i8CXIN9+qj6WuW35IhuTHky2erL59glBhqobQvsB6Vr
ZVLjRg2HCGc3lhns3rTBSE2IeamaLh+/Y4qeh1+R8pFN3Kgdc6xVGjRx5AvM
FYl9p1Q3HVIJHgbM60g/W1bIxhmxZdu6TSvkBffwL8XV6cdquCbcEScfVKIv
9dF1BatohTTjlw8jBtUEdF2bRUkodf9ALi7tNUOUlo98ghuJc8fkwVx2omUO
GbrCXj4kDRvjt5mIZpISiKtVolqJjfgYa3Yi0KzSxn+UPmxG4vE0v0LzHiF/
pQYCcHUFu+c94m9+H+sHaNGaLybPWVcRnocLOk2XiXfv7NPsmIxznF77DvSc
NoTung3qrgYdPaMbxNxPavXbx/sb8kFjz3cK/5cxKlXbqV1BXtuYmJ/n+Gwm
wPjQ1/mX4rcMLURcP0gYLrdfPVsivMVhdP9/zH3WehNJar2aWJ1qesgHvVpO
M6EzSH1ZIElOY/9XIrV7POSIBgxP6aflT0Wr2FpafZ0/uIIJC4q0QU704kc+
1PRvul0ZLh1iFKOs/U+gUtyBbydHclZmadOtris/RdbH7E+jDXFgp5mJQTbi
PxevF6Kjfw9tb8MQBzNTqzhQYZT1zeFywmR/05Ya7+yfkqrQB419FlhvSv4D
OS6FiVByD+stD9x0g5PikQz89hghir7jSgV3HHa5GvEoTh07quc6pT3GHtBz
6ayj/iyZ2ffZPpNiuSumMWEDuAnnxfbGO9OzPi1unONokaBtYctucnz7hbc9
KnjN6pkZdtgp7RLPn4Zr8kVtF/dBVVavBapvmeuey5L6a2HdGFv5z+fxX6nt
wCZRJ7aXCdMcEViwHWuVFIB0WJgys/yH9zlttHvKxB02CAU1WZ0ElxVmXy+z
GwbSi1fytLvLsFL7M2iGBriCYDPFPcCJ0k/T24UDJR87AbK65+heDz1ohjkF
5nAT7xDavQOeIapTUGUXHeFd6CGekJoPHRaHsGdMq8itzXIWM8BShUuTceGx
fW1qcYhpymDXYrCwvBA3AYDZKV0sxZdk6CxWWQjiywW+cRx3tOhbuU21nnMT
jVbj4ODojPvplOanbRugX+7Sr/pHSG6yhQOGQw+5s9RhafPBbnIbtE5rXvZK
+Ny099J1IrN/yAIRiKOoIMbH9p2N7hcUFLas11CPeXiMcnGFc8gFddlAfMC1
u6YjqfS1Ys+P5rLdIgW8IuQienn+Lo/0OksKYUM4R6QGi66XzCQpqjBkFhRQ
dGOf9q1qfnKXpri2qVNYMxqMgcNgajTGZxVONjqoNlFyDmfjHKoZKPEuvF62
77u1lbxJ1pGRmIh8UUsh3K89IIgvuJyMQC/klPAVT8p4L7xigY2VYS4HgY0i
wgIRIHUZvBIbqq/JNhHKzV/VQY8XlTDoSZ0inzeJnfmu0B8/S5dRQXJ34ywj
FuTZWVeryl2da7vlY4Py79vydD1jdWmO0pEsJIDxg4lrF1fBVQezSIT+ywPx
KVRZFkLd0f/eHC3H+0irskV2IZEHDM6raoyZO89XoppcycvLYFWmYbYZAum0
Nd2/gLoox4WhLwKKIFAD1l3gKls09nj+ij4SSzQ4IlbRoH6eFnw34p4uOBFd
kpQgo9UJlUiMBMn+2vypIaX8GEGlxbj2hR9o+89JaosZb2txrchdFkbbEbGk
jy5Z2+/Gwo0/S61SlF0F/ZUGhhvpf+YPFyvKcokVERNeaqrC+pVhHVxJdGts
IwzAbiHRCTcWpPr09tnrFkek75PBdE4nm0+buFtZBfBcSbvFS1BDIqUWSrV+
XiOAPYhN56sA/Z3h4p+BKO7LVh3NTFbWvsS14RsUWyULxhxRAR/wmBJArxLT
fVZDE52tTySoDzuqwHMPHTS1rUDqgddsenbkzUKTs8VQjDyhzjpA+ZZ9cZmq
aHVtlY7r2ja0Rfo/XRaA6HUnTWw/PGu46LZNJwndahUNHskU1Hf7a9SOkCRi
NO3yBz8lVq+p09+4gPgAUuIkPQ1hiRrBSqji/TdLTpJZPBC5mMH2mhwmpxla
fHJ7iJeCnSykWNBaJ5FP+awqwzQCcx1IYq1EdmTHU1yaRpahv/631uPppEU5
hWDNjyRbDmO5DDqSyBHf5hSO3bL5fbjecF+qYAoI7r514J4EYaRmoUJwAuqp
AkI3gz6LQeYE3puCdngdMmmXRY+7yHEAlZxBQrcYd5Y9Sdk/7msTRrH2Wt9y
zw73COHOqvvo+i8zPjiX/nap+TBDEVklQgaZ+2z2ePHD1up3GAVI7lKzoLzi
ntotS2SgdYW/w8ZwWjHmXm3pTxR9YdUgQI92uoeDnX4i3NXjXCi/UciQLaKV
AICUbnjl+8UoBxMuRU4tTwhR+x7VJ44MD9V+jBSLdSBzYQ5wX4xaUhMkP4Aj
1RGzV8oa4Yh3O/ovaM9nx/3Wm68VIUPlR9ldDMUVnIFpHanFPBOYlqk9hFIF
aRADaKo1ZvoIk4k2l6SO4ElUvfWCm26if5uWiBdOFy1aN8e2HzPG8srNfBSv
YMVI3JM8tah5vtkDZ6yQzxlNgOGxfrFvSsPjoFQS056QlsRvthEOkTuBEjlp
iabuUpbUEZvjRzq5CivfVw88BYJK0tRsWFoLtj5LhViVV8fkvk3H2pzT/Btc
OiLeDQZnl1jKlZ09m2oGiSmHxdm5vWfM1cRzSFpBchr5kgjo3PcOCezIxdVR
z25YjynkvhJGuDWW5O9elfudA2itNSpu9ALwZ7HUushbT8M8FMxxWSDMBeaW
cnlYEOhoKSRdKJQwxgiVhg7LVGcPKiQFVznxiTfGPS3uMGKCkSlcnAbkDk1J
qPJTHdJbDBLp7IP//H6HqoLsgZZlzOI0DePseo1uYet4NQnUZjppAHaJmYDz
C3+KgVXS+etxQzVcPXEilIcZ7Ek0TEU/JGEOcCB+D7x+dCm+fKjeznwE14Gm
bKn67J/XOIWl8eiz15Zhv6EbCR/i/zPHLcKhzhZO2BoNOcklHwSG5tcD5Qhm
dGoV+gpQEI+JU/ilk0MLeXCuHHS69f+Ufmt+1o588d01vKV2fRT28XRkm6db
lEjCJlLV6CS0+57/1CZrLOmvLtOKX49TVk9vFsGvSke89uLvuEsVTOnXOitM
R1uCv83XaKgMZF+DkLkukE/b1h2mHAb/v9KKdjb+gi77cKAsaxmuvj7epQox
mKlBd8yERT+Gvb47YLULs9iMoaQszBrWfBolrU5QyBn99L8MRwouyXRAWUUy
m2i23yqUpWbEPBXZBLwg323uvy69WKkNHycLYLVFPovP4G7FeNTV3DF1pO94
tDcv0bz/1o0jDvH26j3DgckVY2iEGuveTHA1TN+lYxL7ecl0cZZcR848nF5V
N1fpRwZfXxJ6hTxujNP/3XW8qgr5jR0KFh2fryi/L9guBn2vpXr24B/MIreK
WZIKgoUFrewItrt7Urd45c7RyMwH0Ll/Pi+zRlPbukBEFTuhIwAppw8ZwGKt
s3XIEEMWUvwZJJgZz4qK5xh8KzOOsjZYGZfqaAbJz8MRazCQHEtRK45WC6UU
xDhqrr5zb7xSpqIKajFitSgO12PCroOICfK+FgncrLHT2H1ux+t1Rj0AKiui
w2UY5x3Id0Vn/W02PYvPOD2kuryCFtyriyUgRhzdafTu8ieHQfEEBu8ICvLp
iHn7vwLEUc4YK1UwwCJnpy5eCepvddPYvqwMHS3wnI99QF6VQBxEH9LSzvk2
WIMA1nUvvauLjWd5KOB5tAToEgcanV3rE6b0eAOaEcM6aV4N76cJUIfI7J+W
93HDsFOQG9glKZqQs6I28IXIiYA2fBBKp6S1w/XhACY7Lyc207+Dbf1PfWC9
uFldnZop3vKVHpr5IpR/F3R5Lrm0/hsoolxANibEluonibq+EiFYiClK8m1d
P+g0O5iqOzskzaabL4b2RoMp/kDDaOZL+geAZW6X9zhx6tRAWguDBZFBmalR
4d2tTxLLVDL9UzEV8ZoC3XTToEjN/yH+VpL9dXYtY7pTB7Z3arsUhJ8+s9FJ
vPzcLmHxYl80LmY5qDLLOVekrmOLnEB5yK0ORI65yyiHCiMWFtgfhmBLiDdq
1iQnnyF51gvfphJhhF0CBneplY7nABB1k/CyVCN3uLApdPz/9pz4NF9n0r9I
hhxpMIL734nG5AMXowrjCo+MNQWSdPQ/EyccOSZNQvCydNR2dNOe445eKfRd
dpsT6xxMGaIyeO3hOegkdnqKeWNX30ZbJ3RI4FNE6SEKxlXYkWDPzXowUegB
8eQmrNtbtJIS+P+5QC9S3EXp1NKquqEFtSd3TShm6pORvHxxBd6ga4FFJvJQ
v6BuRVqk3XaprhbEhllIpvQlP6I2hWi4HeRM6yOUxd8ZrUL17J+nDGtB9kuy
et1Oc5ZLNWenOVnUvb2JJPgubIT0wHv1oJryzY2Br4eCFNGt+Li0fcCnRnrf
c0IQ/jsCvsWHR1zTdbIk7Kl8IwW9DSc+Fx2Zzjyw0qP8BbezYUJzthsWF/DN
uSVFmNCBH2y4bpoJHXB+FuVaDXZhuQUUbobBLmfmO3dKJicehshSyWqmVgcI
MLTc7w0C5gsLgnM60Q8fEuynF/6WZJD6iI1oGsJguqlcbsJlMZInCaicCgFg
2EOMslUmFJa8jLp52BGymQ8a7Lr+FsVlEL1eImDajybfhC6MB5ziAcc9zof9
72srSDRSrpGRjMWYHQD3w35DUdUaN3EnnFQKCQ9A7pjM+B9IB/+LxTiPIWb5
VmiMXskFI0cNZRIU3O/5tQmaMKLKHwbhI/xeQtFZ8K75Vh4/HmmTpWUJkG4F
f+Z51lmcVSrrVzRXI6NuTn7fXLwlN8xjQXNHpK56xkT8K2DXZFNrHSGNiV+S
uMGvTm5FlweX09z2PMiGbUcoESVUpzti6+k1wwVZ8TB2rZ1MGVCGuOEhS05W
Yp7FW8NLgyYCi5ZXU7FwFxQsNSaBRJQGHxLVLG5Yjdsh3K0zI0vnSLOFoTZS
6QVJ0PPqMJrRWAa3/a2YdcPTwGd17glD5vdIXjPg3YkezToWWzybLas1qFJo
xOBSjYiuSdI/Bw/k/mlCe1O1xEriBQgvwYI5rNLAVgzCXhrkEOJhyVNIwVLJ
GpuyLpfjST6oVmQnB1tGR2I/fxTOqlxZT95qtg8OGNwQXS92npQM2ipBQSgN
trjZz5MdyNVZhCCjNLQkTUwtYH1W72009VTD684wNg7D5WrABqKMKg92ENAR
nwwGh+bhI4AXRGV29iYSBGj0fuOhhcWxonXG6l0+CEQU0mQpUPriu2LdCKxm
hX2mhwuk3Z9WgXsAHl3zL5p/PcWS9NZ9KeF5P5MrsyoPwTjSM1sU8GpXjcL5
4xDVwmf3M3rG6l3VN4t/eL79MGxcgSm5Y/xW1rchV2y8RDBP4mC9jbLJws3n
6F7top91TGNbjQP+4X4G6NnxdE8V48QGH4ouYPsWAAx6HIVsqLQjV9fhCZ2L
cpDYbLz1dmQ7r8OTeuOzzJISAkzD5I09/5SRx/u+QlrVgv0SwvaN1VsxnRq+
MABDzh0scmozFfiVtalTU9zWaJ9iARdhSBxGg/CEi9US8c1mA4rCaCSCMbAG
qQY1b+f9fdtcXq6L5U3F59kuOwPjQsEEuktuozRndYwQGYbFjxMx50r+737f
uPePI7ChmTOFt4LfkfEUvgRGdAIhVncs8IZA+HdWZuCXECi3+P5xLb4imdKV
n3tal3b6jbQgaaTMbvSTMFaO0U/hhqcQWnp4TsGFnq7hGmVZmO1frehX3CoK
jaTnGccSEQDL/AKqHAieoMCJAC3E6prQjnAWPUFgQUqQqzOI6vrPTxg7eK+C
TkpkUnntGDRq+YIVo/CLM/N95I3AMVhbSFVcFpYYFvS67J8s3m1eAYjqsFIK
yoZUHZOehFZSvlhzOTeXd6FPQZCxk5KXI+9LCKdV9d7HBqDdxpitke9mUGPE
umKLYXTLl+SEmFniSiINpiYqSx82e7xFzL36HnDjZPPiHC7SQkYi6P8pOdfE
YSQa93Hb5RIhUFvJTI3SuyXj3p2lQv7sd4mdBSJsH7tO4KwcW8reoRfY+FoS
b612XO2X5cj6oVzI7mCuTMfaVeOwgrgFsdsB/sgx81tqYUN+TJrGp7sKwmMD
xx7TytUuFqP6Vc0lKK74jiD5bjDVNwiyLFF/PTUf3KnCHyYMKr5lUegMFWiq
ehomGzLtOst7OMhT0rbG3wZAtTsexvTjzhrVsp5PKLwfiwewPBFIZAbjx2t9
ZGUnAjFVqICbxIVti7CP2en3R8l14WNqMP4zkyOys18xxIdGs7iXdIyyLfkr
pdyDy6DLEFWyFu1kH2LMc8xT7W+qqdSRVsnYCXlXFOLIs8Uyez2BZL6fcZ0t
YrrJIPk84FP7ng1UVSwncMii7cFZwjiq90YnnKA8TDx6xLeDLcfBLDT3Zldu
b4pIvbEX1esoIVCJdxTNKxyz/bHmX2hVQYDUWqSnNnArA9tk3bOvHM0JI+Se
Q9s5FIxPvFpj32FdiiCDS8FMKUWGU6nBIdf07Ge7gAT3hp5mUwTvdAtIJ08R
SouZq87Ocls9k4RUZkVKHoOPAruCiwDYxRv8NKBy2YcJLeRQK5K258Yrobk6
gRwFS0bvvYuBgJxM9u0Wk0QNhusB1ktFW5a/1EmF+385PA8vIpZfb2Vh+KCw
0VkAuVpBDj+i1GjdLjjUTrwhWvrvr0o3s0BeqYIGo/KJ/ccTWUb33w3DxHJB
Be+SX5MDvUGtym+3lEdzEEy7UsH0q0rkS3CJRZLECtBX3yygsyudE6w4m3jk
YkOElKmJoE2WwCGuH/7R9N8V8KBc0ZcDQk5h2Cd5Oh6/1VlFQbW/6oLJVAc1
9yZNYrqdbWdmYw+6CabgSo+ZRxpIH+e7Uck4wJuEh9WIWzBQTvCeQ3eVaZ3I
SsCKZ3VB5rlgHJM7MqH69TcaM5K23JEqWmvAmCa5IoMJy6OhGl/HqE5Oc5r4
Bf+JBKobtGa95Yc/BeJbijV8TBF5kC+9H4R0HWRqY4l4HJNA7r2A0zrFeWIu
8TlQWldx/SFxpJPOtvNl6GP9pR+JvMHSHr8astBqUKkva7/kftOUch7tgo8B
H5SGuwvyUCv7Wx6WvZ5NyjRq9mJeTvYvg+FkzHG1Ces8SiSYPnCqqBoIn1ho
wr3vvcXN88eZZCH3hfUD6x3eFO5PoFM/QuLnYZcXBcE4ZX4g6cICkSsC0L1O
iPHXB2vDBqWyCy7grJHHtnawepxj/uonOtYJhnkowGat13ACTOiwdtkpLZug
lh8C8PUkqASQ1xvirHXafYQqSQZ+0h35cYO4rtoOnmOMr4tgtX3TqxlraLTl
4QAtHC7bxV6mCvSxik7xrKxEi8fERHNqLnpPuw69bVWow+bbjRr/vMuCz6D0
TmBtcF/Kn9KWn2NB+/Nb9S51BlYtM8wTKwszuMriRjhbrFkS/LBNWyykznYJ
HB2P25jVDpeHjwWxV57s2b3oA/wCcsCiu13UMMe4IQn8aHl/WsBfqJUcvs7A
MIXMwGZACbL0kDM3SaeGmpJXLD388hOnztuUJUq0s7MLtYm2VtxqKE0W75sg
eVJJAYOPo8mPwygzXTQnipBSk5vkpNgMWN4ZSrIKtPV1oE8WCSLUI+yqHfbb
wNdQVwMgcapLdiSCwVwfxf5z1fczqlVZG5G56t0EpttltbRWtw9wW+VUea9O
OphSc0Ca5P3KRi4f9fqihVjElTOE+3pV9rgU5kcWB1yYz+ZjtsXSiizc95Bg
VMagkjHxjKVUHf5nT6D+mO0NS6/c4NQmrtkUU4UFHdD3tp9E2xn/OQNCTwUn
ZjZ9to8/uwLqLCVW9t+gVNpbM0wUYLZSE/lTqiYHy5o5iQByAntAn6neiGeN
ZxeYI7uLAVGusnIIaJsTSKlP610R8OmgfeLOcv5hwDYD7bFcxk49QYxZ6v8X
9sC7gAs57hzoWpGOF8sxgsid66MDlGBLSakXNF1oBBvh1moikk2ZaqtZvmPk
xZdZSXX8fqv5Ff6amp9bdESnb1ywDOJAk1s62f7vkqlTQODvyA0QbYOLVkSA
QTk0AWF9IhM89u7kyqDvueJExcEq/UHvoJk2gLWJxGNLtwqDEe4WDJt3lOJw
P7r0vXd01RDORe7pVOxIYwUywWJx658UyQVfauqQGmu16eszoNdC8YTKHe01
WPlsxKh5K22haY1Rei5TnmfPSqK9lE61CCTTRQHXd1TPxwhEup0jFeTi3z/V
/mF50dSCP/AyI/fhIXFcy9Es/iAW6EH1CJ9z/wHtWF0HBW7Nd5Opsqrihwy0
MPzIHbz3zxiYP5WmroSrJhQIQ5mzDVoaX3J1zrXdLEC4EVLW/ixt+fFUQNIk
Ea7o5esqp3anKwp7qTJ+RcNdZQyFsiZ4SeZvS1y2BLR3hcoOZYn2Folpyi2q
YrCwsyIr5WFgqbyXJtqcoPvK5R2Y18avs2jo7fL+RmJQbtAcOMtyCFql3Yg3
yLCr30iunE6EokHDNPy7aDogvyY9mOczPhkMaBtyqCr0YTnNtGb9GMhwxCs1
SO5MYWAykN3moaB2ikE0BiSoucV/Ovx57842X/2Jan/pFzQRglqJZHhOjIJo
Y+uCsE+YpdE89MMAD5FWc4DQetTmNRx/JLJa8KhvVoa1gk1BEaxM9FYZ+Q4w
ntu1/zfnDmg4M0m7aG1g2+Gf4ZG8oI0Fe22aXfomV3/iga/72KoiybxWZXme
dfNooEq/Dgb3ERfnwxHm7ucNIoHfyn+fvFfdlYwY5uysD8mEiNbt326ThkRf
58TRFljLbBonCTUKbhYl3y/7z+3Ol7NuaA5WlVlfSRQnnk2HltcB50ASOvIs
YHXVu8V56I+O8Kxq46jlPOYcE8xaFwZIwO5bNqUOLSc2/pB0kCj8urzqcLsS
21YcOSuannfdQkMSBhNNRP9lHvZYFmzfZf1BaM/PjaRjpiBERtR/GNtehwNi
fBSQOYQNybN9N76cE2Iuos9L3MVjFJR31M6n3xRkJKBdgfa+kWwz2DOY+WaM
SUNWDqFz6EXTfBVVCJ3XJG58fGWtsm5ktd/Tyn07W07AXU4o7WouNFW4nZGt
4Xb+WXBZk1LY6V+0dh33FkDMvCSVfVtFz3n2T778S3uIZdFlS/jzy2cV1+uE
JazgCc64+MhZLHOQKDk1JaBu50ngT3HhtD71LBVLUb/JREOYcf9VqO3QgjE+
U7/BihJATCKcaIZBeGH/QwcDZYFn/GVW60xkhvtAtYhCpOZ+YfeAblnBbjsn
oS+sBUhlSam5xy1II8Q3Hhglz+2z3IpTZP86f7ZatTTx3s7DFE/LzRZNStuQ
QV/1J5cSmnyi4UPka2+KU5gGaaVBtMZXLomnKSup+QGGGZ0sMF6iL6xFsq1f
rUPcpqJHmKNA1Yue+aEC9HGRboqy235EBmbCzXi9VZ8UH1oIYaoEzS/v6FtG
MKbANrNdK3UPBCMVc2xtNTT6zpJm5gQ9ZmBSru83GLN5HPlE/sh+obkCqoM2
KtYrv63SOquPWIBdw2HtO2J3YTah6haATiZf2DZiMuiDL6ZKSza8xY2Rh6bL
CY+YFPqvL0A50L7pZxxZ3M5yKqrrn/R6zRaRZejMRN9Vgq5mKV90M2jA0ZVU
B/djE+Dtx+rcEFofaPA4afcXMtCcQb8EaU8KNvbDibuhjyx20ybZQDuMUb3l
UKqp/TDiE1qWS6IA9uZlSBwnwx768KKYTPpehiI82RrehzKN9vf/MikjXJje
lB8AdcPcWdhXrZwIE12bmEXelA2G2UzDOb2uGaDrfxPPIO6Wha9mesZt8jhe
PgNgTrL5QXRiuP3erTFaLffor1laaHFuvKZ0F9lln7nnPAmuzMrTniukmgMg
xS2dTQP+lKs+g/lx6Vs3MKrtsh9KZe+4ak9EnBGrgLt/+ffWSh/Hd4Icc9W9
Hhd3xL5C7YdA/GuP+P/zhwuw8l+F7kBmY9ljLQJT/KKCmYUPB7WPubUgfiUb
OL4j/XRhPH8fnuLsWoLo5IG+EwUuHgsuS9M5LzazkDu/LVvx57os7XaphqQU
WFLFGyPPOXbQ0cMf5Z3LPH70p5EpmXqGo6n2PM1yyrD4S5b0dxKWS4t9bZhb
caNu2TecJdV9n0WwJbo1GaYw3NXMWpJHM4xH18JgJ5Lu4XLsUg0/DIiVgASu
NBuMahNhrhxZTE57Aa6BqjFdomgPxwBvH2Ul2vpStXWsAzgGxwZwnZmqZbEc
7M225gyVfLrcszhqefnvd1vzSp9Mo7cxPtcdr0m4vqzoOQHd55JL5dDKkg2q
mS6oGNmqrZEZRTDTJrOcOAFwGP1ItpIJkeq+m6AXPZqg8pqFt1+a95poFJsa
XjuNLNi9oRpP/FAi0rDIanGFmGrX30mNy/rKoJc0H1i2z8kXfdzkC008NShr
OPK5KPVsJJ3cjj2MRsbIzX4PLkgQNoxCcgSUjmH2g8FvcT483+sPDVSxJI/q
fwm7ZpzcJOeh8jOgtUHxOTQhYJuf2u6UyYKbYh7arzZ6mPZ9NR7NTFpE5tE1
0+Xw7da/u5gX/f5nxP10I5SP3pxbBZWXEe8l0cO5/cw8o5RM+QIClfo7gyvv
OZDNJueRA+/inZHIZsLFWXwKMpFnXcTPCRAOyZwbIun90XN0ufzDummNM9FJ
j5TRZ5fJJRAUmtmvBQ1P2qVVVZy7JNpIYT4ln2ZzSCZE/Xqyu8PAz/WzEE+G
OHcCp+hisPJjVqnwSLKPPvaw/eCPnugOQZuzlutkYfHFrBtmdmRJHvQjiqgV
ukoAv2bo8GPJjTJDZwDAyr0ZMjooU+/o862wEw3bVFefus0uOULlpaR6AuVm
Nuz0CQfTeX9u3em0ZbPDPxsOcntJWKnAjuPwU2YRUd4X7iXQlUsDrcwSvR5C
v0BoFrAW/aosbhjQNACKz63Z7ZxlJ37jbE7UIJxqOaiEuF1+CaoKrvDdMDxL
5Pmy1tR847bWdI8IcmZPuR1eiOLW2Kx9/sh9Z53gr43vWqbmzp5hdMVE6v4T
9vEePM31ZEk5r3m25aJ5dJQkTaMhyqqFc5/16PjtOJiq8me/v0iLu+Fg2ytO
gS802ujtFLgW18JY/FiOJLbwerg1+wgBY+WbfI6wBehhmsM/yKHsdyNDNd/Q
ecx+DB6LzwKFKiaeIuEgr1U9WlZWsjwj78JRqzvqENw9axHpS/FqW8s2IPxM
ead5znHgNQEKwCsXaKhqavHUpKJdiJb52b7fmdrmmz8QRXrLtGKSmuygCpRy
brrhhw4teaMCKAlKzw0cohnbUmEjLDgBvo0rYlcaNLCUMuDNfkHOA/ox46zx
Gt6SOSkTUy0vH56ZAY1C38N27T0SLU/6fPFBWXmqnHYggD7TiOChLdbMWWKg
BHuEms46tGQejGMimsjC9Ou2NWYkX4uh8VGAKb4UJmOwVehYlZ+pWM8Rh/CW
so0K2rZ1fl9DkUOyEmMNGc8IPZXR4AASs2aZnu3gqx4iSvnAhfQHDU6eQgRJ
TMan1STVgrRGpK3uf/78BCRLUKknGokFc3zMiXyi7zzrzL+KruDHwQMGZfIR
lz1ZYAR/fSEkFwGLWDO7ENIRl1KXNZTKli+rVZwu43O92nwEVkirBIJDzvwY
Javm9vsmVbYLCaiWQKaVOiQlxQZYA6dhdttpU39JWIKmy+OavZU0gjvJE01d
cpQMjSgMzjHWqe+R+ejcS6Y1oYbI9wIbaTrEjT1wjRI27E6TzpSEhXQVlfxz
GPghlmwGfaVIsSZjCTukdpBTPvFSqS4g410sCez0RaWsUPe7b2u+FxP9Gq+U
sAsqHm1wdIG2niySUgnUjHqpGkq9siWhFJpsae3N6ocz2PJrokgcimBk0JW+
XHOQt42e93VTtJlKvhLGVHXs3lba0vfWrjFc2vbllqGNUMFGrcLTuwuJovBs
QTX4y4ljFjhrDCGednfNC+o7VYgM08uR0XGnV4qFahVbf24sV2iNqbbDAg/P
E3alC/Qv+pPUkRxFYkZoiMHKd4m4tIm0SOHueyyhAV+bVZSWUE8cozzW0HMA
rnY34cXy2A7cqxD8YOH0Dp2wF0gkQZ9GXrTyn7E1w+uCbICxMKXyTx510i0V
XZWkMRTiyQ4/miKvuHlaXC9gjozBRBrsuz0ycmJl5Pc5sD05EjnFnREjanIG
KdMBg0SIWF5MUAnDwQ4S2VuASIR0dycMokdPV5L5EpLw8K12eX8jiuL2VbtS
WqM/VjT7rlFRLCLZXYUg+RsPLpDH3j88syBpI1VJIMpUNdOnt+cGAFPOYK++
tKVPkn/XdMw27hNAu9fM4ogC+OAOdBz6ckljzfzxlgzJPD6WMtwhT2ZHGxYc
kP+4YMZJiOsIKDEV0+ITQKjUJL/WS9Bk/akFjSFXa44Xf7jjWdFc1YeELYuS
GyW/1dWEj8IpwI42vJmOiAhpJwb4EKnWy/30VM5dplkxIDAkAFIvddh3pOAM
JVU+uy1J/k3FYSp04xbOdEYoHUJI1xXpbSwzJQaW9Qq8ktog692+dBY+pk9y
GsmMXBWTH9Fr24Vm9jC3DyT4Kx7RQuBDhXlGkiJegRnU1G85fBx4UBLjw+tg
nzSETtbixEoho2EC962+l6zODEkcDecv2dNWCfUgENWoV48n/E1UIaUaGAsV
DNlqIwviDp+FeP19EOosqMMG1Lxybk9pSR9ciIqLkD5SohCyN6sI0bveP6ql
U+6tiAKacOyxoVTx254O4ySECgT9A3Xe7FUdFo8B56YF34kkN5aWbkSIEZ0N
bFZtvYXPCOmuzOhgoBRo7N0UaPovYUSObMSFoEEc6l1ij1f6C7bea9MYWISW
k8fQH+xHZXhoJzqkI0nv7iXGkW+oFwBpbF32k2f4OILt+hP14rqGXhNavnPK
qsxu3CBvX7jacgd6OTmuVLUX+e7mI1wUoesh7dQs2/al0BVB4K0EYEoEYJa5
ig7lzPVImWbjs32BVLQA4TsSXEVIPPajp8XGanDZMILluOdyJ6v/+SG6B/FF
YFRpVcp3WDtKk7cOeA6i0xHkP+2uef2EFJPZAug28VFPrXC3jvPiUWzbpX1M
XbbAGRV5YPVUERzu6TmZdTQylRThGPRwia7pmHgeOSOJ4AeS0hwPkW717A3u
qRa7ZeL+JRkuAl2vpTLoiuuBlGgZTP9wt9a8egARbJecibeSRHMcv4KzIj2S
i6Kpf5Ta1NMcMBqb8EvG6C4nfTa16Taybd8t/eHo3PoN1ifB7J6x1/be1rny
yPwC/nx70Z7wBQwjQ3bnfbp/oK3tBEbn9rjwD9SmX+3xlEkIyESS799j/XcF
I/gmQnr/4vIrrSougdbGbKRsuicN92Nqk0JKZPww6Vis0U/Slw9jBIdhR9w3
iPi4DMC6PlsSi1sJGAbHtBpWlJP114Fv/CjwC3tn/ZI75qmZs7FWhNc7NGZJ
5otEXaXNLSNO+fo/C1Qt+SKbEHXl1qp2dN+L5+xgXOuvfw7dDNIUrB1p8QFq
LoDODfRR/drBwCpx90FpABH8JI8FxGNcBKZNayyFG0e9bMlD6r45TFhjIFT8
KLfq/Y2KVxZ+xf6mImhtJ7sGhVL0xjogV+K9q7C2VIxHCDb8+4i1iIx4c28f
kbwHDuT8jODLRbcfzGu6JVom6LcoPBkfSibwRGLAEn1qyxSYPJ0frWqcPNQv
H101+9JJVgiNI9ioK1YX2cWJ4kPeNiczduftxfyWyXk3t1bayBQq3vUBCK+Q
sg+5vn6bnpZmtEcgR/otUAlfRvyaY3gYfNeiPWNgqonKo9J/EaDW0NX+21d+
aMGsDBBy7L2QMXBv8u2VX5UnXgU8UyIjTAH6eIHAWoINOlXiobCyjNO23NhP
rFzitEPlPWbSf2AWlEt2QVMD3i2WPGWrmXZ2RSYmAP4RkT62JDYE9l/NinJF
PbsolPrCJe2gyG8LctBlh6ngduPIZkZi2LPNfTW4cDiHQG6NJkMXZ/6D6KFw
1OBEmwz/EyxJy41wlHzBAA0YSIFZTEK9ui7BXLGmGJrUf5Cn+4S6vi7Z+gmy
BtHEnugMIav1dOuHLf/dnko/xL3OxJp4C8p+8IiXTLqlScwhoVJjzNfG1D1Q
4hKW3jTqnOcaPs0DzYLX6U2a+mgMciWWwYc7bJ1ZvQqgnm6MYH6bfAe7WjCu
7hSJqAkQqgmHepYyYTiBkba7KOKPVL4p5duB+3MN14mY8+Puf0emG+yAI+Vu
DEp0jDOL6+sxeRQPoAUqePlpCinESXbs1KMobb/d8DVUxdF40EWnEnCZQeYc
dxdXYD4N4twHJiSbDciNP+4NE5P293EPR4wNQc8RVqWqty2t22D8GDxs8jLX
PLblLbw6ToqOMsM/cR8maXOixv6HBiuaEZcZN4JDsV3gGxmn+/qoG2H+P8eJ
XttYqpQ2mkoZrUR2XA+MHAx6miEcbmXdf6CnJlrazZtzsyF2Tj5W/SDa4k+I
1fl+eOas3xIE04WVw/alxy+W3b2B1saXzq0QY3uSRMOqYDUdCoRfZj6bqjhv
moR0zGEGLQge/x3+PVBOiU3Y2S18D+9cL6VefE4/vF+vTDdSFB2g0EmdAlba
Gfq2agtBv6ca+U6+QOHkGE6YEXFEEy3zFM3vlRMWhuncDk8WnLM0Nihj+l00
pP4//BMkTRN25cppPu/1+gQpgg++QKagOadnzgFnw7yubK4VGLt4sAbIxQOL
C+7/cLKJPwXhY6h7yAn1nOiZWKUb+wmx+52PnnKD3V/oseDUFDE0e2VHM47N
1oH22iaxwkn3/0eXq40388CS6hmYYq+hOzGLLTvZaK+Df8I6ncQ/GbuLWfwo
7K9thGE63+/+7ioOYYlN9a5oAhvANee2+9NOp2OMjDpA/NkfTLTHdcXjJQdK
njgkJXthT7EcyAwiaRPHK6StxU93fi2UPi8BIQVFigVk8+7brn84w+wEl5ji
LSgAcZ5BzWfafGj4/jXoxGeYiQRSxOO2+3nnN+ycFH5Aojg8nB7d03PLDko7
FL7ThgiJE5s5lZnqeOv4zVvw7/qYoNeuT7rgZiAwGwoz4XgJbkrQ127DXzfN
Rht393r53EaCXfVJwUFBIo90IrHHGzh5FjohnI+IqOfUQ3M9wabMRkwsQZWd
ycRfFA26OeJ4xj2ivs1zGj/Vf9PdQPXJVoMovlDCKyb4L6HC7aGUAvrgI0Ha
Eaww7PSxTHG5bAgvt0nm3FRMn9bVqn1JJLyFBTCwg+Z6bnZu97E579OuDa/e
fAQOxV0ftUXdgIeT6VeP2k5oUw/5h0X3Q+/+g1DEPk6zyPxma2bpR4OvOqal
VIlwehW95Rity6S+/8vRMWon1ITSCTd41LeP6P0cPApMqJYVplA8Ounw4LvI
qk1x5IX9Niq4CVxVtZmG3jdzhrzCwFwe93ZxJ82ff/+VRoklRlQ5g6FmrPIX
FNyqclaLIzbISESy6LqTq4EYvEAOC0dpIZ7w1i1/dOuY2saTa6PEixSJZchV
iFJvWpf0ZC+Mr8gccjxKiy1C8AGwjwcRVC4yD8nMQMvl/0BkT6xWXyiMpsHV
VE8RuYna2vbG+rh28KdKbEwPNVGKV29nYt0KVF/N4V3N5sRUGmDQy/WrIh6U
EoqLd/b4itWUt4jLJVImqnukmg+X241oScydtmdSDhzX0H3DHVHFfb7XweF7
S/NbMnSB27PaOuHIq8SSVV0iF81jGabUWynr6xBeMBpe9l6sidn4yxX4Zp0+
LGwrBmfKymFm4/04Og8M948KOFiSw+2NlHdqr90KhBy6INxXHJhKW7bcfB+M
YCC5opdn+PairphnT6IeK0yKSLXG83H3+dCxM4lbs6qDd4pU1CbItlHcm+KE
QhRCS3BKBYWI0pHqyLxKlLA7GBcrFJ+f+u96rDfQ/faK/1apUqZmJehg+ZWW
QquVRRzVGTuGMEoz7psCD85CoZg4tYMJZaCRuOBUiXmh2vnSdxaWsvyLZAJO
oDaIXDXAnGw+5LfrHLlrkYEP++wyZ8iONWVUscoevVQUnGJ9tPGIK5jQiaPi
Qe5oQTTlkRBrIPbwistCimyG1+yRVH4HEh+0215cd3JtHbkjYGOHGo8UpxXw
CcnDnxZyyXXgOJsUuPoaH1IYgJXhyNLVuGbeWJ8xuitgUVRDCRNC+W/pQPIb
vdt7bdRc/j5ycYMoiKurclGASqpjysq/IBy4MbneLO8URT5w2HMMPT29VxIq
AFmmeO6G0GccX8vNxQkpp7JDZ+3tVXnjOIIIrAScKfmhTcklQLL6UpHb6YPT
RHhfXIX9n0pukceOqpyLftE32DadpIsMR/nqBkeKDrxj/ypSrrqlH1M9/Y/A
Q2hTagbwiZyepN72pG7vbkHUIGfZkQQdLZd+9kcTWvyZBN60NbGmYFBKf8MP
sS9AZDVbLn3zzO8xuq5IGdY9irXLNX4U9ukF385mhI5GgbyMCfQwehfJ4Ip5
SOWKUhi1D0qfW2aXxyWFuAGVZA67I/mdeH3ISmpoY6vVPEgzSTmE2MbAGabk
SubhEk/cj9hB6q/yGeyqDV02+rRV0wx+tBr0Py1wntsKLSp/ZuSwp1BHP1+C
T9IzfLHhxJc1pLHILKxZSVGY5z5Post+kKjVchCPfx8ajTWkbet8dxvjwT1q
KdCXJHjzbk7bb168XME4XpHe4sOS0GGL2FqLjRqfdrfAAs9zfsuzOlD2Db+2
sGwLCZAjybXTYpedG7A0LohTuItBVSvdpnavbPS410UN9gLM6RnYmdWn/0Nb
7Y/cTA8moh7Hcq0cAjXyX12vulk2S5jhaPCwuXPFbhSkP5S20STQ6GnwhnR5
JqhR0SUvYJIejUJlbL8vrxz01ATCJMxb4GP1GsFVi2bcQdql9ir5NJXYDURU
wnAeuJ3ZSSweR0OZ1qTJ7woEPEKD0bxHaBu0ORE8fCOii3sOYrFQ2Fwdn8nT
RilkHiZjZv+3lFMytyqMh2Hi4LIojlF0h+IUF9tiQyG8BHq+gZFmSxGCdzFa
+ttc4fYO3URj6vZEjoN8tOizv/Ku+BAieUdDzt1MlUc2oaBJe0OZsD98Eyys
ygqKYQzt4u5/vLxSupyEpp5E9DpEHzmuVK2BRGnfhAGmG9G8HgW2YsazYxxd
4LX+v9z2EM8lbvG7s2DnqrWfhUbzlMmqZFwhfzTpk21WYgBeWTMUV/3AuoJB
6ksh81g9UBOhH96iYbc2pT9RwrQZkte4f2OLjNb5NpwHBVaut8MkIngp4e7W
ISb59xmWO6tHrfWNTQxEQjwSK087uW43VyPU8FWZpE/bnK+nKLllE6j3tMD/
ISEqafYG5YRsDMYmxZnoY3WeOLGDETGVfLpZ/aCHKj8e6WlspCSFQ+zqbfrI
9+8uLPZSZGq3z6WgzJeExMdydqYm61NTe4jok2neAqZnnRhfLEtnSFZEwnYM
+JzVzmsvWjOfYXNSc6mx4NL2v8RQGr+YQD7oCor9Y4lrlNy73aQ0iLSY/HcJ
zGQxLKYqP8GMzzOzQ4bY+bctgN4ERnMLtsCiUEjAhd5sOgN4Azby7VMbNbfg
CtA3aUKbr/MJ9+jMVB3wBM7j+tBTEDgmccs3DIda88T8QfVE7dgNJPvLU9jA
ZvSN8DiB7fB2vvzaJa7F75WFZHkzDsRvu6qeCNp74TA4KZ6QvaS9u4Aiboed
Kk2FV4gDeoSAcGA144BLesBjSMUnYeZ2MShyz5iI4Y08pyNh5MdP2oQzYf5k
StC2cckNgsmIm7i/aixnns/r4kI/jLxpCl77VzS+6NevkjgTRWuxDSiRDICM
MMirkF0w/Ws9xGLBE++cpVAQ1d6hwNmKiAs2MYv+gouVsvIbDfJyfsQsCpHV
AxeciUgLPdVQivr0gd5kfZAuxfS9Dwl0W7ZGj0P+d0eMybQYZFxesSNCbUSj
Eg3I+yKQDHNuF97yZGEO+w1n7MnKHzxMtEGlj9R4rLTn6xgK35cmv9iis7m5
6vHNiY3fSPBCJhOA3l4GAzuQDCuCtdleX8HRxDuZ4yIz5vbQcrjsQgnE6R29
/gXzfhWO1StNI6HqhBQluFozgftAixmRt6tieg75hcl4A+XiH/AHLNkdUOUw
Fh5IdUumMI0jBUojFqpBufaiopPtoJa8nkE5WJKgybUAL/SyhwAeegW7YBDP
pK6ZmS9yc9H6Mo4dzBXrzkdPwRytzBCNzrQcu66p6IKo1XdidO4B7NCg4m2J
biF1vwJ0l8VFtPBU6C7r9mfnr1lLQ7dCRXW12klFADnv6ZKW6VG5eiZe1zoN
kzrxxz3paGSpqZShlt+zWDDMvP6mCu+fC2lJbjZiOy7hAAJN9rbUBiWILZzH
Czvbd8fmce9FoObIiPnyXfEHnlmnABCVjnb0YNTIb3jeU2u8xeWy70fNbkIR
WFV+050v6QGQB1IvTyHILQskLH3yAYrJhy2l4LiWkM47gO9JkA4GnfiIZAVh
s2sBu8i3ipl0/5cesPsq0NMHES7gaLBwWfi4Yd801d0E5kJX5NUUkOKSHIYb
SZ7JMF9ioxLsJE/C6wM0f5/kkEnMrmC6VYc6jiRunyxssqPpTSTPhQppG9sI
fK7FRhNl0Ba2de6/xlEJkydlHAmm5O8Ma3kdhe7uDOApSzCkAuSv1i7ZEi4p
lpHaAnVZwqIX1Dm+yIUZdpb3e3JNmGuOMNZWLYa2Lj6y3c2wgOyH2rtgtAch
Wj/+gkCMMcXoNLKbvj92w+wfX0DtSjNY5jRJQ65MVO/cCwr+cmrkxgB2lCcQ
ygCZv70Fqwr+LawpwSyYOdULkZVlCEb1RDxut/oRQiWjb6e+N+4Gli9jPN3v
EAwk8D6ohfpQRwx/MNBtCQMYCxZ/d0PcvxyKIs6tlKlQmHD2yG9IWWejr0Eo
ns4HYsvx0WYAMVMqfYHjgF+FrM0NEpPbR6QW88lGZSLyNqfaJZXuoUbh0XuC
YuAxV8t8NQ/WrIy8H9kgzPRMWPClVM+1vG+Qlk5Gf/pSrMfgL+t6QxgzJij1
H+2eXUblan/9xXJ4Ompim0DZhWrg6JxyylOYE41Di37D7/80KCIauTWhPBrg
ueVsJPD1KpVwdVVyKJW8QGNAUQRZ3mbpsIZkKmsTgy9LbgA+ebarBaycle3+
7CYRSBuaMJGtVjN3HE5RR/UKwocaZf6Oh8icGkeiKjZ/eL86/jzWmf26jzYy
j0/hEbX0oKmT1Gw2tCoYK6lZuLzjOBXvXqEHVk0yvALko00HUOeLbDf82nN0
GpRQTwk693lJmRBt0qGyh6+PFTogS+D4TPhjYfQ6QD7jZ+RLv9dEL1UjmGJp
RpUwJxRz+gN4L/q3efKj06kCQTS0h4V8z5GlGUu3TQ/Pomrge2fsHo9bjUM+
EaCuIc0lq/m3SoKMjmF/FIlS+fYwmyWDMDfv6ncs2U5A72cYvMeeEfl38HyB
VXA1z7pS+jOW3fUOPHw3JOOP7x4M6fQ+vtINY/1dhtqgRfX0/b8vYcClI/Mb
8BB26cJeXBjWXyhBrWDCPrisferbYZWYkoyjWj0zrEVIV0HdCw8X2Br0m4Fj
w2rXUYFXNXmU6z37POj63tlrvqF9DzxHADWBlOgALia4fXNfn+1yenLc0ECf
TaZoBuaZxRNDk9WAhzHeCDczsTWodxH6XT27T9aTFWq6qVdr5NBe8zNy7IYF
ysSaRtdGyl3mpj+23EnXlRRNbfz4iOnsc99wXCxKYp/F7GzfAp6xGMmYOAAJ
5JNUWgHT6DWiavVezU+6CN0H5pxgN1DqEb8bCLb89zG0iPd/GNZjflfETU3H
yA1+aTX5cXD+Fut0TzsarOYHTqvXqZu1QxbDtuTZ0rVABhucomkXmykY4/ws
D8OyrnQ7DhrtfHKk2BUdfFrorKGG01TY5/nRz9nXhCHFt8JC4Kqy61X1bUT4
nqM2qlxwMwYF1J7pqDP/L9eDIGhGwGRa9IbpArMPfdzPZpq+ls+NpQjXK7L2
X/iQQYyhWdQ9tj12p3NKtnK2ETtH7OXO79Aby0oYlonBjYDIRrUEU3e3IAdW
NF6cqwmFC6RIAmmT5r+W3BEnp0WVj1Y5Ebzq27wdHG0QfR2vIP1sUIEg4Whz
HjeolV8swIWaFPW78VvfaAXKM+gEiuvbr02i75YmAQO2ROBfy9ib12JOUg9K
g52f5aP07oOskRNhB7bIHQkWz7vat8yWxN+OwkxVz9qAk9eMN1hOCEuF1OWp
hdaHmfI2PM4K6pdeBEy0aygmEq/AwdbwVm2DpYniN5jOxkUw0oIPE4eKB6xW
Dfg3NSZ5hXm5tViR1BeMiobU7NTHzEV2YUuB0Hug9nEB/Vtsy6/vMqsK2wIX
4v9BVXdMZPjmzl/ATC8qFJ18mGZjqO0ljSRzil0/FsMMwSm1hA8ivyduNdnG
qTxP1PZBgPyYjPA7kR6ihX3ZyA742G+dj+o2Lro450Wl4g5gqDOXn1QUE3ts
WCVGpyQmaStLbKVDDrTP4isHT71scVINYmudik/jTuovwrdMtCAsU4lljVPG
9N5cVQUiFOZLMJUMRQNKeyd0ue4kMVUjXevIph/F2a8+PmOUG7yMmx2TqoKr
HPI9uDbVsdxu6BPfu92sX42ChOKvGMOe4BcceWlvnPF8pFxbNWhUVFof46uI
4lTD7oQVqX7tZtHCZ+AjXUrfk0i8prQPi522oPjhUrDrObamYU1ktGf1fEvf
2mmiu2myKcE98ZQbHZQGO97PLwL7OYOELu8b+jD0qWkLfRnGHAEfRNdBSv1M
Jx/D0TrwXgZqY2tswImXu+rkd4DElz76zTUlcBlLcMz7fAR+U4cso3kdCgvG
7hR//idNwT+DXI1phU16UWtNXkXGqRsF0zTLpqlt+jcsZUtPSWG453n3wilB
L5LWd53FIy+AsgZUPVEtiXPLHRYjGsM88GWfEmXkMCIkaOeok6QF4KU/Fvro
XyFW1ZFtxX5NEA27X4/zTm95hYkJzfM+L64HCSh09EDvLBvEj9kV8IYP/aZ2
odrtqjIUqjYOPoIqZqYpRm7XFUMYc4MQ+m8wnH+ssWRJImG6PLmC8XsW8T16
6UphD6IBXfQHA8IKpdGARLQIO3X5MURqjEYkw7o48DnQBDiHRO427kdpEs3U
HKXXRMUrwysDK2Oln0R1bM6ZgNjgyH7nSIkRKEiZG6ZFT92+2AjKIRb4o0IO
usnoOVBqopZRLuYF1inF/CIxgB8kYsXIfx30jKw/lG3jI2YHPTHoHcCLeod0
T4dAX3wuQEiYBnbMxY/LWGMD6PV0uXFcYuaqLJDHwHUn4TTYFwBMopLviSSd
p2VxVnWExxsIYde+cqlyGTYW0SXNfN1M//TayDJ6W8q1ReNQiXXKPE8ndyS9
429pwhZrldix4pYTO02rq57UEeiINTO3z2fuUbBvVHERt1M9olkpYNVf/0Lb
J0mbmFI0ChWwWbA6cQsZgPI/RTC9nmrgZxpH4B05xtvZblMlnRw6CAq85U3A
dHmpMR7kGs1Ou3e+eohrjEIbDzDJ9e4Xo6xuEg61zCQO9lr1IwDN2pX5yuu+
XJmr2MNVeDaxv6NeCncL208TXgKJfj7uYstqteFnPGwANuwU5AUknFfkVpJo
K2TjgZVrjU0SYOdyxvk7kKIP0miok5jPn7j70LbZXHR12Te+7qGp35TosQMd
0hyul978dTNWec7heyC5HucNZ4n8WtMGtQ9V4ECiNo0wFQYVFcnuErIICNtr
2NqQYWpCZcPy3YGS5AinvcrOWyo0QyAH3Hde9Cx30p7TmC4MOqZ1rwhyOIuA
AH/ngUcCbN0T7NLeS3mq9VPp3XmG8vHy872MyuCwQp7a5WhcV+Eqr5NwDSCZ
yzlDtL5Z9tyGc4jcye/8jk86GgESfzMfm1U5cOjWEQ16SLjthTKTD/kcW7Ti
AkC1lJmNrG8WtHw3a0k02ImV8pqnl4XMtXB7biqsETFmCJWm7tpUv2qQfMY/
4SE6NdMeKYOvO/cqDsFM5tVYwzlLAGXXRNiVEO/HDZdosNwXkPD2pORGks+E
vMCEc8dzoBvPGRqbcv6GAY8C8kGLUWBwPdrexdAm4hsuEvVYad64YiaMXnGW
G3qJfclkk5rQ7MAFSjhzi+2idK45gDXPGvOmW+FRrEgHldKCkdCBlbUMQH1U
r/1IQeR5LbJyHVZnltMA5P/YBXTIYEldDqzBf2YM1BH7vOGg87Jv5x4vR5Kf
6t0LnqmWk87USbDUZNwAFaFRSwrm7Wk+AlCr2bXebhv87OUlWBeKsSGV4Uwc
KX+hToQAlynwirXX3HH7+Dk0H2Er1apbxsfetAHp5swbCsICD2UBona58IV4
IPfv/Kt3z0d6/dJ4zu1eb4pqKgQYo7DYuIJWYvMOr05dJG9OgCnHJ83y71h2
uxMpIwpJAf6bY9iQPNK6PoOOzpZEyRFdwQHs6cnJ7N6KwIc3v+KbRxLslh5J
p+ZvbdN3aBboAwhK647yKGUZn3nXIwU03N3JAGlWur9aoIKOHc9Gs9wjd/uT
VbqgZrZWJgPSwgym22ITzcXNs4+ZdBmympSxO46Wu+ZteXp+d6aoqnuc4hJ/
foyv6hd7k8YcNwXVLdYBurM5mhjZWFKoeHg9Fy9u3csAaiUkES2tuH9YJxz5
u7TSXK5ny2s5fNwWxGWDN4o5DX/0eC95VhlrZi4sKqm7qEYINSBh6kwloI8x
7YEK0r89Io+Gm2YkPFoIW0VB2JWK/OY6SfGt+zkVq9oEDomPULbKssqsamC9
ln/P1zMaXgRHIyFrDOHp6ySvG+4FKRl/xYtpCStAJxlaYSVps0pWIDHr38CU
BHbOU5tIauCy2934N9hqxgtdTAluVqHhbMW4tzwWEWMp6yHqu7FqbKyyOS50
Byge2l/C+LSuOhq0ZBYIwo4yR7hVRAKNO963MJs8REkssZueE2aBR/s3r+lM
CkMgGfYNrt4iVPJURjuh3r3nwsq4oV0v0kro4VFziJ1DI92MpSLPrKVldtrf
XIxJyzuso4Lmp2ukxYBnhAqCma5lZs1aF+ul8u4xW3WuS5j65kvbV6kSFmVZ
gEZQKdYGec7ZSzkBojggGDWwqJNuUXVSCdX6tBhikXqj2QHAkth0mxUfzUhw
/zk6VAvWHxPWqhqB+NfT7tuLRtHC+2VoH2KtWPAkPdnbgVWkTVVwhFjraRoh
YrBPEumfshPTlLPWgOHmzfdbVHL4w5zpjChY57XeH/pu8zqAot4nhE66o3Hj
NtubX/RxGtlMdidNt3qu8S7xuTcpHaZ6s/d+Xbz654JDBbIwhEtprmr40kiP
W/ZZfflrwoOEqSxL7Tg3ACXSPcsAZx8vAmyenelun+b98tVjVukcg/bdzE6k
s8YnIDNDzice7RMIlS2UXXH37GveMg7VwfeQPGo5Z9Hb2k4LtkynI4fFK6R6
caqFBjbW+piIFs0aSjKsUaf8141P3C3P5eSX+f7Aavjs4Aik1zTGd1Lot8Ao
x6+d4cY6tBKPdwKdTNmTOA16+onNfsR3sDtHB2cO0BZjcEhu45plR/pAjcn6
mdlf9HTh4fbyeqYk/rWbc8GeGKUHgTuS5azVBUSw0jLSmwkEYbgxKgSW1gop
cjNCa8oSqBj91Q0TVTKyMooDSp5JBoWYXdyIXRJTMY3Wcc8/21p4BdShWWYw
QpOgaJlPYQYOCwyfO88s9YA72yhtMXIQAjV5VUljNZkj8ZyLwDlJ71AuuLs0
V5MsqyARQjkd99v2f71qcmWiRr4fW7pyxg3jqxnXMDfFdqRVzst8CmDbeB5q
s6hIsaftNraAehh2IujDzzKRaP3n20WLQdPXyXbhLbKKd+vCLEjwfviTi4lU
0Fq4hUpknFSmidxJgTyz/fv52cTPRlRQw9HXuMhGMhTcN7wDurEHneP17CDS
JdP0xta0uwaumuTAmgqBjOl/IbJkERYrhugQhiM6aLdx13/rCU+XzSsMLdS1
3x/IRvwYbWpjJnoxElMxEoPprovf6VFU0X4gX9hJybSuzEDKAXYKndz2M6cS
Zl3Xivbksb6F0ACO/l6MjVX6gpnUESDG0BIL+bfGfhuPwOenPaDg/jDNX6P7
eByjpH9jlOhayt+wpDmjxiVje/iwH0vImRRtLTlpXz1++dxUKXoV+uqGKl8g
1Xi3loKgTEVjTk1Rl8a5hW2cLR36p/TiQIK+CchtxfXF5INHFUS0SfdLfzW7
bms3TLg0/ys36P7eUX1ce2UXYWyyC2oJH4dpETXAlF6oeYgKtFEGhMAvMeij
otJmOJDE5sSiWk6O1+z9gvnRCxCMpgtsCr71pGExgOOcgOJ7Cy9ESJRFHISs
dd2ejy6B6d2qQrTnD+7crXC41xJOL7v1+v/sIYcWc+kD9JPXMkVh3zIRlugo
ziMDaFJp7sxw95asWr1wzW/lxYBEApvS2H+g40HsvgsD8kWzWkJxUDh3LA4d
CGz9F1F2/Vpkah2DYpClLW5dMEcnOhd7o2zed9gK9lwZoUaSl3jArRIm7JJ3
KWy9dk6SjXOA47U98oKaDAY2dSqgi9jM5CJF3jTFjBG8RA7ksyQy/+W6mz2N
QQ6eA0E2cJ0ZXqiH3BRqlcpNT8qBAJ2z84/SC8gKw73Oc1bpWO0LCAZ0D8gX
Spgrk6tYzS9OPTrxoQ3Xtu+I1henkzz1ZpjZqt3p1/64qk3/rxZefqEl6JNb
DEyC0W7Zp6SdpAjKswUKuAPZejd9jux+ZnA4x/5lWrrhHz/Q8qXqa5NR3I2z
JBPWKV9gwm0MdtwCkB+Wy3CQJZGwr5AiFSc6jIX2hgZIOI7Qq3cA3jrbVLNT
CQu/3KkxEAV2k/KWO1HnHnYI60OPAWvzQIJ2MB/1dW0tk8EvDMDbbMVC2oCf
8xa2jOZEtpzFGJX04A0dNAhwajkMyEgAo0Pt6z8hxzEakRkamvw1NgoK5UWC
XEjJH8m9zyrdS7tyyi64FHxtwqjCyYNN8usuf3kzaoAOYSO58F9r4pwoI3Kz
jzR7cKOg0/dfP+p1aQ1/XJpVvCrfrVw67zU8+gF0KWilJOfaACC7yKHTvK0q
ppC89ihMthmbWfOn3pbykWYUhattp6h0QqT4+mjFM2Ek+aVYWBeUIQcwu/IO
C+KBcku/zQk27hUNMBql/fnbT64g9do327u1/s9bllFYExHlb8G4UofcZ5fH
W9UUnnMyYZtcisL4/9IluEY5/NJax8qGWjBXDFxJ6SzjuUWy9CYrO9mPVMun
F2hoj0ZNTidTxm/xqsDk5Stef4f0/nX0cG0Y06YHyrrY8/waYgNfGe96zeUG
qoXNGD+7PZYset2IkZMu8pmUANDFZRpYSv73eHzb6y43Md2TWy4ZM9Dhcx4N
MsH4m2sZWJQdFDBgQfQu+REzHsiHcVrb8adCmEHxgc1vfibiVuiCxJTsnq+f
onG7QILRD2X3E9WgEf2vWh/8tRrpfZInZWM2D2jRwuyQmGU5Ka0w2izt6sry
VQqa0LD8YsW2tPrKhYVOOAPDWEPz6dQLMVUCRYyvIaF9aUGvO/1wYsTfkhoE
EBkAVsnMr+yWfFsja8WD7tqFhoTHCdBn9G9v7WaRBvpZZqIN+/buhC62gp5/
aYCKa7unkOC7s5660xU/IdiOTvWUCRyxgMF+dZx7N4vzLn0MVPeNhw1JwsB5
DjACFl9sNUKThoK788vUUQeRhZbuLaJOm+yxj9WMgQADZAngYEo98HUjg32f
6CLZyBIGYFEAoZIbJxw8IJDzEKyzmBxV7tg69WQKnxMR+pnbUxPctAlM9X/O
F89wXTT4j7zGwVvKEnBaQ0YUnfb7sUrj04OPYZCfszrXG9tz6qxWsotZ0PgO
uQcJRISGiFMGDmI9P0BY2JzWmH4+v5GkVgWjWCbtyJtAxbWcBmBHFk7ywLit
3O1LGj3N2gpqAC5fvlePRY3oujZiPTL/1D3trAuH4YKgn+tUZX0eIoHow/7k
SZxDXz+ivmUIBPSeyLJlZRTljOuzk2qqJ1QOe5dQ9pfxJppJ0CQzlwCacY5h
h89YW8j2IvAir/eC4TDD8Mb3mFhoE+2KUbpzrGgtEm39E7RBnQqnowQWsCAS
lK3NmmCe9jfvl/qR+2kGEZq6CuO/t+vn8XPAnEnK0vkl3hZwNk+oEkcHia4c
HEdwS0ximfJEY0vpFmv1PflwPuyR3I3ulD4Uqrbh37pp68WJz3l8cqroIiQB
pSHsN3luMPE2qXK5o3xUgr+WMkvRtyE83gtOmnOZPBNEv+FP24FD++dNemqD
qy0273Np9m0+V7siFkG2Pc2T/8xmGYJ/TYBY//pcODiwbkx98bCD+zh8rM8B
EIQbWWifcXGMU4VPawX4eD4JlFaJjQbWqmXMes8IbQ93tza+ylVpQbvXqzbF
UiV4ymVoxf4I2nZD0tG+AjPuGfGFJ0OEDsRse5p1mvf2QUIlP2e9y+2UWqtH
8JlYpwnXZ1IlrREaI27jXrwNGAog4xiYLzX2IXMjEA65u6hyg13F60KuxZVs
LazOIyQ6FzUUy9FNwU1l49HAVe23dOVXQ3zflkPW+DRugUYF64zC6Av1IqOQ
VQmLUofWt7bzluJwRnIb+p4DFLz4JqdJrzx0OxjWT5OsnK7z2mDzAsoLhqms
7/MxqG8iBlhgl21hWfpat+t9/D5DDRUs+j+25lCxh7yhAwxvRIQlj6W9C7gk
cSgczMezQp5F6BPPhnSkumSeSfenLOMTXptsUdrJHklz1zEFITq/ymSZQVca
6HMoKT3f6ztTivWLhLrzQm7toydWE39eeu2qQ9K3j6/9FE1ZLpBXxfhYsdaj
ObzfGb35tvlGYIyv/mJIDQ8ChYyxHPkOqtVAJNJxrHg/xj8jtvJ5o8uvPa6a
fd3oLAE7LoFRk/++7wt+Xo38YXWsTOuMzWcLl8HgIuvEWlbc6vk/

`pragma protect end_protected
