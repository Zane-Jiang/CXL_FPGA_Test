// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CiPpC1N6ILxQHp4Iq2wHUoEpKcBSuX2WCno/uYe6tyiKkeIzpUGpgybcGFWotNGlXwbjgyCedT/3
Z7jTltQzLqq4Meot2GW6IIpEb87srkgfWapfIyCVSteqGGK/Hei6qaLMgrHYOOEsAdGIKtvMx4BZ
eutBP+pL7+1AhV7x6Fae4gMlkdvVEmLmrDKpggRPG8yTeBCV5aBWeL6mb6/t8H7VaFwJ5W7Pp/b4
g4KHc5lvwp+q+gZeQqg+AaH+wyTKOm5yzlrkDFKnejtYDo4dquUi9L5N3r5TPYWcSibUnFTQ5ctN
7j8FjmJCJHysUS8Uc/QwEx/e4gpdAZrHY5EMAQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4064)
OtP6YaO67a08DTlsnevv2gJLMJl32oOIEvR7EJ76Fs34cqUHb87bw6oa+pVr4RNvLNaVNZyVRF4A
0rL1R4gku+0M/oQm/QhyHIcDURrlmE/PWBxJ+/OOFlzp/c+LjFAf4dDg9YXgwJ1yJ0oc9273aeuU
QSe/gubn4ieO7LifUfYcFaqFVPhUhIs+xpp6KQGPw+grjTuXjdX+gWggFNZ/mWtjWigL7UabrEhJ
pqEb8Sw1zIc91dzdEiDcZBeSm0IzKIN3AcMCbPOSogQkEqUG3T7NpPTeufd7kJa+PFkAWsd8Ls4k
0dJnxzSpsDadTyQGkF3nCWPLYffc1ge/MPhtvsW+H28eUn2ER1ykYic3SZ+kdSKgV3iR3H4yERT4
qtxw9KSMXTJ/+JUKlvJ6WMpQTDmlA3k8clTT20zva9X6Gom3b8zrBEkIKSQtfhSHqm68xLILBiBu
Xsw1t4lviuOC4lfq/fLfg2RGjU/hMQC73W0TPZBduBX+MvO66LV+GD3bS2qJc2CqgofNPR2Afnpt
AOhRAA4o+mb++qHz8cXNlomJz1Z4kJw9DUZayfUyihHI0AWYHuDgytJ390BkuCimpHGoTGGphU9i
OVQXtXykqKiFr/iJBeqIAEmhXZDkYUzb0W3P0x2b4uu+iaP1chJUUtsrGGvrvwPLm8QD4+D/ln6i
gAiGdy5HWcfk49rKPOU8J6GFgsFKOEibIMylzSU6Ajzxg/xAt/o9H0gjP+J58Kp+HE+HXvNmw6cL
tIWOr05/25FwukOB2t8NXtbqGr4o1Sq+tbE6uPDEgUuZBBfZoOIPjw1AdLT9RVIPKUZsbCLoIpwQ
5pS/OKy+ebhbaUpZwlkZEltcmebFecGH5kSBAj+xLGSBvrGFUsa0VQX3CGiLOYvbTn6ySc9yh/MA
6fRVTZIQF9bDg1kPV0sH0CX/f4zUmEv2lkmQSOkzSqOIALsQeMsXdDxS4sWccDtD1faub/B9cfJQ
wpAj2/gs3dUXoq3aOaozzsH11nVlxQDYxfbHCDAH9jRisVZSI9faW0s/uNIEnxAtVS5KeVAsI3Ej
IN7hQfcVOLbjn6RCyqYWAflEFyS+1flInZaWNOb3QQ1JbxaorKBnKsa7zvEOe0TiPbJogLR3Qs15
y/60ZE6ctBunJBB/aguodkBzhXYJEiY4NFXKwXyiPuMBkINiRkaNcr/GT0fRaynxL6s/r8Lvf3jX
fH3bbHNY3C5b2W9pGXEvSejEyBCu1G23c7rBGCC6DxWwH8ePvFZSNSlSILoaS5R+ll6l/cMd+l9V
V3ZBYxJGHVBbeD+ZjpXE8Sqkg475LUiW+3lCwlIEf5LtDFSArZ5yYx9G7cWqsSRNaFMwhZqMu1qG
2kICxC8iODMMqdOBNH0NrMjUk+33Oo29nbR3uvDfvz5aXC7tp3TUSb+w3Tz3HDrCyXfAeIVaKa3d
mRioec6QjghimecHzKIhgYQ5ssIbXTbKgJUyIkYyXfjFXTD5qzfPD3ZtNG2bTqmgyjkpGG4vAprf
t3iPOQEfETB+87rNDVKFFi4ar6OkhRQsK6K0LcdXqQomOhIbSnUZFLj8sPLKQQaXU8xZ4jsPZ8JI
aQ3joHd9iiGHsgQjkX83khp181rvq7O0pFigaTRIzceCmp7bYKRZA2l3biET6djdjX8KeAmvqv0H
b7pn9t774OgYLy3Lz+nDx0WXXbEJ+UaFZvelcIzWSInoNTekhFht8+QLz6lr0uZX2+3aA5sxPFsq
csb7dUtnmlioy1sVckejatzr1gc4cnWcckHvs5+TEhIlGyUru213LB7w1JilTN14RFc7kbQXAHw/
3bfEpPucCiAcCMkcF7ipAeKV1CtEQcaPv930lQSnhzp4RT3QtDM6kVo3V1wps2c9pT4CMuMxrMIX
bfO/ugNcYG1TbtWptlwZ95jUypb6qTLNYxnFz3tSMu5tp8S50BXV8Odz70DLdpsOyxKXHenKmj4a
u7pt6Wx828ipNejmQcNm/SP7TgXpj1Vgc/JqK3UX91ktVaG3yVnOeC9gBdvKdRsougpDcSyVJZ3N
rs2/3pmpX1AUGGoGfWhSK3RqSG9Lds+Qe3+Ac24nl6OSsfVPKLJTR8EhzfZMoIcgZr+01/hsPiZw
ERlbbKuBftY85g7QxD11aMrIJJ5lC8n/htKrswB8QLo2kDUbwtjYu1Eg5mkCoi42KkevnmaiqMZg
/0H8Z3SU/LX79wQqR6CZuZDBY4axV7QxEHokcvyUwqUoKhptg5OsoUrfXEyVQ63SR4ZMR8l0lzki
LTbmn21ivGGtmmass9cAGAD3YX1lub1it+ozPxQpAkQd0thoE8/6CQE7QHpy6iaRsYxyIYn2RidX
ji98VU6BbJC9/DwkfHEfO6y6LFKx3XVKCZ6zXP0RwLqYJJlI8iHYACJG953JopqFNpntgCsr35Ki
HAiQDQxLrhyV7ZkuuVW/dgu0Lwq/OH4myWbuetme7nq1BMU2zVScmClAaHtRK48K1VAfkTbQDBP0
iOxtO9cWak+tSLHSFYCnMi/2sdZPJBl7A2OyGFLtfQHRIH1UOIhV4BgMW949e62UzyNk6XeKYMkF
QWL2/aQCvTiw17VV7Zmm7g/H9MXVPwj3GbY2VCK3SBVU02HcOPFNBxhSMKy8yK3VvWOltwWBAudO
JAJRCR2FAEPfB+8x7XUuOUgSs8hzoXtog5MFce5ERRnq3LOe0DdhMXFZIWPr9LtEAnbhpnUkzFUX
w1xJrkjrdcSCEnIqm5wxkOVS+E8bIQZR9p7FoKkMaxQ7BWVmNSjz9oJF3Z5OiPGU0Rz04rfO6CTX
0iPzBbZLWXbAwRwkqBhX3Dkksdf4hvvEpoeqaXy/MsoqmWMVx5H831NtI9k/bYJNq/XzQTDX+uSm
H6hQycxN/pnQxazhH9pvptDzK6M9kwxGDeOPx5yvwk7Y9ieZXL1e71vWxg5HaEdXvlX1IxZeGjDs
eQlMrTojRv7iKZ4glv2LUiXO+BKx6Wj5Ual1AT9Oek4ggNKLsW/CyELKBycQ/TdZGOSktiTdOgFF
QrCs2a82ogLBzaJNMawRrAwbtCfS4jXDb8SGf16/l+/xpHqk9SyZRfgxeZVkF1d89mpI1s6X3KLU
eWIHt0XLdluvxDHPeEmVHXdyIXjrZd8AMmCsa4srFAveYdF6tMZdy4CLbGGfbjmYamRhKpACPi9w
Ncl1rPIm5JHf3rKADynj4VXty3g7Wz7kEnWg66f5KS2LA+O72WeuADzaDWJiDeyjEWAloWe68axf
Ip5rH8BWAyzAP00pRka/a4OCSMzBhzMM1XpwXN2LleVR9VbV8yuNkG8Em9F4ody7hzpRPohWZw4X
9G6e+vte4hr8UG/7D5Qz60WVGzRYrgK0RYfkpAM0Ls7HHg8AYQj5sYQJFCE/IoeGMvyvGJeOAMiQ
WOriR2JihXe4j8rMiyJQg2+Ka1YzfFHgrOBagbZMBYvKEfIOymYxmTQu/44JTmTT6LJ2xWnETqBK
SCVx+NYOH7pFmHgjphBDF+r+HDxfllqkSLhWj2WQO5xQHqtuwo2OtmjYl2fOCZIlVgGzmeH1LDeJ
K6lW8OavnQzQaYKhM6tBO2HqjwmicPFo5reEpxebruDXxEgWq5DwNy3/3v+eG5Rte/20FrVzsDKg
hrlFC0XZd2yjdckzLnxetKN0LzPX+ctq5v4TuIxQFR1fjij0n4Ir+ejT/B55KiQ3YwgN3mZ3fsoW
RSV4S8wQsllntHpavyrqQRaQekq+aRd5Ua7B461uS4yqcT9G6+qFpTOXrvcBqozdB+5e+QF0I3En
k99R3VDqorrUfewWnT/p/6D9RiebfKhJDF88YJwFc23FxhlYBvAQv+MCA3FfGnHO3S4EEULBUZHy
+Q+8fXvslvQ6295Wd+a6xmrE3WjcgEv5I0gMWSGre9t2UBOtZVDD4Li0pZNgF+p3IER7ZNj8HuiT
igzvtvUkXUqWRh5EPAWw0wp8YEhBZyHaf4UXvmYv/Bz3PcVQ718ZmdnoxDVQ/AG8yDlqB0Apjsxt
FkgTFDVdsYgdJap6PiXfZzQ8AN19Fxu4cGTc1sr7fNrLcAxbTTQIx6039CxdT88KgH+eDs9FRzX7
Zbz5sHq+A/Dpt6Puqf/cSL3StLI91441aDeaqdQ8CxcFzkIc4+N+EQpK2q4Oy8xP7hlmx4NWMsag
XZQpvU3LCwNUftrp72XqcRWXj1zhT7pKFB+njH3YEGEwvGUEArquSKcYdMziK+arQkZt5l7l7irK
6jL7A3j3eoDAK2GA/O6MHLigSPrVu+Q9xTLsmkrAgwJYCy+nlTv9pR/NvrwjyOV6c3Qu1u9iR8R/
wleiJSRnE8yu5SbL8XNo8bNagz9kn7dEArVz5litZGHP0HuyFuTlHWpCa/xgwjqWAjrk66ueBT5E
xaasAnZhbA/TAXLtl/9IDFFlTov88eH46LsYcgPcWPLPe4xLAHDWAcJRYTRTzVkmaDSwSUxUMvRX
H4i5F7SQ/tK1hreXEJyAZsIWQTR5+RXOLrdukUVPE+n2Zs3wnqwpyKu2igvFeuySI3jfIcmdH6pk
ruJb42JI4eiuABc7Lnd7NboceGi/eF3yWJsESgBulA79JbDwFCVZa2Zg64qIExe0l7J/QRfgUU6T
33efzx5C6/mTICFB0IF7jCZBMyR955EXuad+SlH8stSlsRxmKud3CMU4s62Xvbe/EKKVHm7LwS7z
4hB2N+wPqbdBMyCJTkuvlPqiaIqCloLo3jnLVrJkkCXCI5MuKWw05NnyaRMjBcB9XW8cdnRBJKgD
+Uq9zCqY9GrGYIEEnM2O1wOQZSgiF2HmwX+1/HJKbR+OReBbkbo8gEkf5IBCA2NOaqyeSgkIAGmh
j5yVoFoewvbZdKx4qSSUu3/ofRpfTa5QnBrpIn0AaC2Cpb5j4Vp2RK0LZEV7/XuQnfLdtfPMg8kc
mO0w+4Ouz9LbWMdL10J9lZvIyUch4eDvylnCzQsYq2AuSkqFdbxBRkPx38jprWJ2R9JNlTEy77My
GRkrGb65e+mksLqzrR02WHUmKuNGxPVpJk4qnbqGbZuWUsPZxMZNZwNJ1EYst2jKwuY23ZQ9v8gl
HqCpNGpwMTbwYxZNU1S4PUkmj/Hyk4fOMG2iX/vxtjngmDmFpow89raBY7scEg0mhK8f1wlJEptQ
QqOYsu/bPdESf8v4Nc4KqZBSLHK77zPMVKY7ZwU8cARsHT0gYX0Tvke6ZXY0rWjEeRyRxb1/I4ec
Z8LmTORmAp0SbZMt9qPSbrl+uy1PMLMRTK45GKLI1joi6MTcbfDcwcOK5DmPp6fGRi1LJsWkJ4wa
ypc3CMRcTxWTHEeIrgoZS65t9BLcVsYs/IkCt0lZPcrIz+CMUxTcl6C4GoYXFVyuaMJZiCEA3Uzl
EaokyiDTVrtv28HUbMExZiI=
`pragma protect end_protected
