`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
hadvZgedV8HchRTiWDfNaTzFVAx4pGxeux3sibLWghOccGzlCjWnEnwoYbvqWguO
8K+32rJ4p15+fLlDydoBZ8SV4kt+g6XBTcJskop3vey7ltvoBn+jRXEHe0Iyl2qb
qfkYw6t2JX+rMP+cL6O0u8LdC/+RpvVSBhs1phWWHes=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10928), data_block
g+qhaNFnbaCW8qj4TbPsFDQUTtEXNMjPGMLTa56UtinP0IYrjrIulBp451TX0+FH
usHg8u2N/qcvbubyCz3O52eBR00/rjsk+xCi5QR+WmvJ3k+lXK5RGf0UMPmwxEcn
Bi7MCtss5kAxdOIHvB/nAwYrHJPG4gLfhUfA6lS4uEz56zBrIogROJnBckijtY8q
M0G/wAQ2D+hqRSa0EKrboIl2knMQOZoUmxgZc9aAtynpCyTJ4mAc397zLfbaKiAY
/yGDHQkI8HN9+/0zDTByeTFDavlOdYn7xE0dfS2XkLVJQV+LCrnfGKrhovs+TSrX
sXzkwPGCyTrUd7WFrPCajBYyAo0SWPKoYVKnodVfaT/GpUhxNcqrdl4de+UhHJuH
ctLee/2y1NSTbxaYm6jnbinFJhHPv4O5F+rXJWOSArIJbiGJ3JuImz+NPZBSvcIB
X54MvsLiFQQLpueO2hlPOz2OFK5c2/GZXqO/g2iOGO5iBm2JSANawWx/O1GfgoAG
ud8EB8RGVsQcHwSqSNnn8oQMe8vVlXpnmobvFzuwgumH15jVm82Kf4AWe5jUaqbv
952HAKc7zmyTYbSTfr4fX9J9dtJQy81lLceAgDK6lzbZ/AmlLu7Ijllrv+lJX9sT
f9Sl6AApb+ZVh7RoineSOpNKxFquCCNZ/7Q8XFa9A62lD3I3sIMvJMOeyv3FcKC9
NFjrLwlvK7q7Qjo5QCNhFvfAPVHxTbWsOP6w0GX8Anc7ftikjUJePJLooRLcXtc2
w54aIaVqLsKWXTcJmLsDI0nqqVBQTxDK0uHs3KqivKSqwt/kjutfzqv+qqeVvjzE
euCnzvFRt5YcOKNmH7m19e3tFdyZSN6mV5rdV0VMCi3hrGR3OfYd8dP8wGIfdlZR
LI77SlpAR2L7LArAvCWrj9aXP8zJlUSDSHXbbt371HzjuVqzV8di9N2LrK66asq+
Rc83qNoRqiKkhWCbLQax90b4GwNpEsAhL37rJZaClkXId+cS0yAXRRDq6i7Ee8Ch
gxmcMnQZK+aRx1tfl2nEKP3ykPUmt1e3Hx2oTPJtC99iSXcnZSGjxly1XAzMqHyP
XxjlZJ7HHOWHOnhnF53d2kDyATTCRtPVXz+b9fxSFoZm+QCOFtFR925a969TT0RJ
lUqFjohhtUBpsyJqJgeSzjk39z3//4eCiTawEnKxdVDO5jzoJIiGg9TjPUbLScSM
S7x8k/QoJLX1hbitgYSBp1dvgcVodh7m+gWQW1Ow0/sxdi0pNLelBhRkyj0LAr1q
zhB8fxqV+IPpO8mtdi9UPM7x2TdoH9ra1Yl4jjmp6VnVCplTSpi8/U70Gcn0rfs1
TArdhVsSEMov0EA1LTmZHlHzjemEQiIFpD7BF1wEF5b+xCM3LqMgptzhizLDe8Bm
60Sjgq+stphoQ8AWZbSbEOOePKmc17Z8zepaOVaYaHpLywb+5YyyWeZbjgmo98to
FSbo4hGX2+jI0LZ9+LWAPW1/c+56uYXf70AxIW+0K9iWnWHrayHN6/8ItACzX/q7
KPrg7AP9gP44kE4DmACCHgikwdZ75hD6JsswxVA5bbq54ZB+GaMk5CdLLv7Vi454
G6AIoW3zzAZeMigBBWKadU+bdRmqbKYXzglBT9cn6dpP0o7XQ9GwiP70dq4WdyAp
bE7JhNhDh/LtOahEOkyyXemyCZa4EQ8/2M9aVxCxRKGP31Nk0ErP2t4ewRsIojVm
53O/NhV5/4cl1R3UplsazYcDlyBWaNCIYEEMErKwflULGgxW3aB0GUY2GMq7fqQd
Lm+cVvY42crBMQvG6thNGHwlopnAsVq16LqRYTqUO0X1UimgPMzNTxma3dN3i6ge
iOQwIfqEc0GPPfumySAVT4sG47yuBmppjkzGtglTamHSOVEM8+LJW0KxdZOe4O9N
uCCaertTvM/o9QtcpeZIwM5fYMT/kdWcRwzKiUZAp2snqm3wq/0MFgY5XbAR9u1c
v8pJgdmL4XJOsoEbfLpSrU8+ApAOUeA/CVl3UAwMUg5O35QE8Tpu4ut0/JaqOEEV
S8T5MfvKZyXe0iMWmhdJbEkp4S9vIxGAApyjvD076tCB2ih9C0dnmvr9dDuZAX0+
CEwSxiOl4GhpFna0vzGP9o9PaKDzYdikHZvObka87EwIg+qAQhHH5Sc43Md3Y7Fk
5L5I0D7jsu2lQtnC3k5c/pLR0P53zTvI2aOtHa4WmMfkqRhuBD4BuQYxWF+sPo09
miWspIUJmzrSdqZeUvqrcv7sWOgo0R6ItLDmL92n/o+T9cO7wTDSVB/07aSFuAfx
dxB3SeBmPhP2OC8e4RqaxUNjtzlfOtuf1LWnBZJH5+p6N9AKESNDMCgfTRcX8Hrv
QtQQfcmuZaMyXhw91apMRM1ZeXq/D3Stihrt5/R23lQawAfTck5QTyvaOEXJPGmT
Knzz6whh8NYiuJkd6R9oz7kwvKp/ZLH3tXhiKu6PzQM1TU6QXNc+/ypkMvB6Cvqi
ls0x6ERRWs4b+OE5VBoan9JTv4JrX/qVXSCWXpQWbcT9l6WiES8U6JfT3fuCXoum
RCJRKqDj4EUp6Z0EPcd5QwqIhOyeW1Cc8n4FRIzW2vaPAVxogoRgPupR1+LV75Kw
LG0B0Nq18S3R8ZaBIy7tEvXnG/RLDwhgujQt5ybvBxFwZcG9bYQcnQzciRnlVsVp
hYpus3cHIIG96kxv+zMz7mgcPB2dLSXIOKPPok3bKiFAqDTVsZ8BdqyeWtDUnH22
SkOTbD7eT8ZAnfg3lyY4LVeZN7cM67gdOVmdWhiKQ1K6yo+H5d5meR2bkTP9RV7W
cgv8ENp6MubhBLRCOLwoT85FHQH57NInBSkE5VN0P2VCmIqujBDPewMWfq1NR238
NQZAdWbc5u+rTLEQOG1lynilsQlmoIkBnLc55wLTt8jwYJJg+tqIB6TBv8Cuyrnj
kpitBV+ySzmMnrLnMLohGdaWvWyQFC3UIwU0bpp4+/M75LaIinlbZarKCHEdSWNF
pFN+/iUI/A0LBzmJ4oo+YLd/XpVJ0+W7sncMNAfVZCg5RwT7j96VrRYIHn29jgQT
ukTeIIili609V3D/eH1zHjYM72wgmV7It7H6LAkIKLqzyKqmKEapaCPHyl1kFmxn
JqHlx+nrMmd/ESVVAmgzDhksp7TcEaMJd4xUIH+R5FCEnHzyMq02tebcsJGcfBMx
TCQrMGH+SUjjawTffh5Ba7NENdaLQdAq+ZcPJaHI/RzF+X6hE4ff73xc8ccqaaqa
JW+7JQA1wh4Ui8jDX5iRWWOiXeBSw1SVO3mlqDhroiCEEorIssMUx8DAeiRicqxN
FZV/Y4mnXVys4Uk0iV9Go0IM5/Ia2oDNJInXqA8o99CLGuOpJ/kN94T2rknXrJwh
JsqoRmbB9AZ72cI7hDBIOT2v3aqmEheMgCYj+dTF9TqBjCVB8rfypznh7wGyXoI1
CJgIZ4KJ3PWzk7Ntz6q5pLZjvEYszVq9Qpn8TjpmbJKARJo/x5EYqJOwAcMrYz/8
SW19ZGCaBg+H5Xkv7gQC+KizBvyFCTJCCwpQt7wdwakzPy6iQ/knSy18LutSFOM3
wEFfZytCD+0mCs2uwwYbzO8EhRzSjkECQcf1/yqHWL/3fQ991XxYOvUU8/VLZJTG
9GzhayPdGOjCZiMuFkqOFIj8vMhDgZvNwpXCF5ByUMaVVFbFcT/b06/b7ltUvOUc
0ySDthg4+os3RGP7MoHutdFI0INbhGki5XYVqKEz59wAJwajAOtDt8kZ8fVciHHe
ZnCV+TwxJ/3/UY4Za5hdGnOkmCAB0kffpCKGb9RXMndkSBA+GDLgRdy85Ydon/+r
LIrathARR7pRBBuxjgfelaueyIg1S06v6SpR1/ipJla5XmluwJSatmwSV1oZklI2
Yod/Z6GGhKY5xqYnUDXJLwGz1aBv1r/UbwE+f4wuBTk0+wHhF9TgsXbfMDLBhLYx
oafAV8fKXUMjf907ole4VTIdFMbMwWeFWT96xqvYd9B0OStTiVu+XxYBD1a3v5wx
anVXVDqVLdrIRKDlHR0JUzNgyZML+NUYZg5nSk+/1d2R4EYi7yaAZkAQ0TBWzGMy
BlMMHo+7JyATQKF/AQawB0/J1vZYIa++fY2h3y0orz2v8bEINjgznVZVTgg+JWBM
bkDz6G8qnKYKBYPkALXWaNVyhmnuXcZZrouHwNCgHdnN4D1oLRhYLNcJ3+yLFbX9
5FxL3qZRIaMAh9claJOkyfmp7NzD/ZPD22xadNFmMTvfLCUjqjActSyou22lRAHR
aoUP04vdaQcx8J7TrZtj1X8sDBxfv26fm+YyJ5PN/JPmZkspnVmOWlu9R/jqGTMQ
jT5Tbfh//Mb7m2GoDwZ+jtw49fMVHijNO0gAA/0Z92Wv08TXwaaFSOukc0ZeFQER
691TbXZOHlI15hDTEKy9pN5DGvUhOVchA1NtGjq7RNWxJ7UhFFwcuzv6JY4JwyhM
SzrndJyujNLHtHatKcYNm+9XANYLSltepRLlECiohmLB8BX/r/2xK7qUi8rQQvgE
RxtjVn3nvWt2MuCkz3AZ+qqtirLwtm5WbzdcGw+BXo4lEtfwl3ubal5s6fHwYvYu
hhsyi46h93vCFPcnwaGBpJce7sQjdE4OV1YmuvkA8+d8gvcf40a6lVOrrwC949xM
lBkpH5OLkSCLzKV3D12T9eubE1ge/bvoUZ9NHh2Di0/P1+loVtfEmmhq0hsJ4Ptk
s8LFIfJPv37kK+iQAhG1ObR1PnXcRVefBjEVFdZHa/qeL2u7Q3Z6JUEBl/hO3dR2
8/0yXGNL+gDmkwxLRySb/7wF0VjN8T0+7uQ6pkTa5wYVaZaSD0FggmcxLwGRRhmE
tOiPgVpdMdfSTfqgE4qo3xhis/FjewngVvCxPhFk5wyKoRO4kYGvr65F9NSZBm1G
FDkfDCZ1+28JmO0kpaeNrYQ2LwcWpN/Nc74Xiey2W+KVcTVmer9vsVrdX+cIFZ/O
fUVycqvnwv1I8sUsLnXAi+uxgi8ogDkyTPxL6yjiVRAzKdywfGWXtDW2gNCgoAV4
FLGs0o1gBbpZIZCoY0ml5BFPlsWirtuXJd022rUpJUYScmBd5VtKjp+nhEcnzvmW
edOgfM0CzRh//qWMym7eckCygT6jiB1sRVAB1o3kNPxNiw+z3XOhEnlmsv4Q7p83
MTTtj1bR0z/e/BaeIfARIbwdQfY5tFyui4aPlnemng52o4rI5FbELDZvR3UFgDt2
frBPzhxGZ4sLvrM2/mFbel7HIpz5X9i9tq49ZRT9CQ5oduo45jgjiLuhlPkvjnH3
UpBTolZLoQgN9rydfH5TCJrEYBMPkedl05adNX6AtnkmLHCVMcRWQ+Ld4jv54mxb
pwoLbMWYYTynKLgioBWOLab+MNGjhIQVzsTXWR/gG21UnZGu8Ygnqn5eQhobp22T
L3Tk5jbpK0oyrLuJXMbZ3n3EJJu6GRcEHJIB+aufIKoAeja15Y5ZUHiwOIT0mEb9
ScfPn+XrdWdFyKimzj4bmyBJMfq1zOSxTSrSmvj7OcN6ltDE3Mvl43KEy/+MzUoP
wGTfWvKp9vb0CzzPxy3vN1oDM82w99uvS03+kxjmP40+FKHgO64JTpJQnp9mbBKl
GKJpsv63S5n2ITy1bDLYY8CpDy6YpDZgcGAyOe17txfj7stCGOmZ4700g4bgW8GA
JUgCsfv4K/TuilPQ7mCUGUMA9pcpsk2jOiNv2zIRyU4niBz+uP9NVU/HLj+UkLay
7medWDyqWWPMA/zDIKLtM0AX9nIONXZ8Xt01rrXGW5Hn89a0FnKOHseIWPuQLjdM
E6ZkQYlZsPwlICVVJZBsTXlV+b8OQie6tlg2LPxCmqNGI5Ua6IV4yK9Jdr845W7U
A78ZMFX9qLFeW3sxlx2u8oV+wgrRgrufdwSMhO7SLS3JaXsHeee0i9Zo6okaNAQ4
LmzUtTnDjGDZvgL0o0QYq4cjfDhyILrHYTuQ/jQlCUWUBpG+oKsVa6O6bHuoCB7K
bZqt5/pbnCsrlEH3WGeiVr/91gNjgQG42mGFyO3ZBqjoncDTF7ABxZEoBUz4pifI
4QxQKrJetUxFn1ZAe5BR5AzQrR+46ioJyqBeeNAh17O9uVMcMDWWFOCAmmOImkJy
hQlZm8UY+YUUft9ju99wDu5MjaUp54DPgGIgAc+tAt2/DAkMB4hlxniwtuXah1uK
TmXsFMBkXC5MPzDYlwedVMxsXuGtqLMjWeQBHrVxZlG/lnbxVszzM+GipV+vh3q0
rGXE6lnW96/CZQrpDsccQTWWx/hrJUOfMenuvnfuxpNtc/7o1PaZg2/dGk1hgCs1
HNIkkfoOq8Ei0ibEa3lx8df32OlWS7m86fmsWMf/8rTEtKFChcEHMXAcaTaTg1qq
P/6FOCRGuw2R3de7C2LWQd1CeRb8m+zYbO7T4m6w6XrndL/qolyFoj6zdQIh+NmG
ID4/4rApNZWnFe2B2RXzYqqDv2V1B42mEYKFRO4owBRve9GvG9KoI4Ip5VAXm9rf
d6TX3pw/NqJ3IWVpQNHtp8xG/fpJCfwV33NWCcYtg25CaCms3vBlLQpYBbTAeUAR
yt2CUogbhYo6tuyQ16DgOGzH8Wo54HAN60On+yqvAfiKuDO7Lot78oup2SuCDlEr
R/wBT7sz14+OBOMA+G79KnHik2zUAI8ZvyEuph/tfbX5XJ8PGHLRjnHmJbjQNwc5
lxc2IglsXAgmAuWk44ISfIcqAK/snRfL2XhugnA8cD2YUa5eTg/gKGOEzyML5YN8
pALUdbb7iAdXcxUvxRAhipCY3JNY7W+ZLghMMu5V1uQeTlNciwCX2UnEQW5EKT3N
YSMLmlHWGo6EornBOVkY2Csd+4quoiHb6Z62fB6NXubDgfzTMDnyUCKHIXB8MyAR
kndfCit29Qpo6nsixDawiGHihphJGKHz8B2buK3U+wZwCPHKOPIahoZQDUX3F/N9
3vcwSgCKmzJW2Fs5rwR7SzhDe0rzxKhI1fLWxGFLN3oIeVIRh59NHuiktdZJ4s67
uEZKSRu5FakrUA1uiPJDq0Xh3V/sqryNdR7MVAfSNpe7FrHJUgpdNvM4DNpv8kqo
+kZaS6Rfklw0lBHgSgyYua9qRIJrPEoh0i8FnQY3F5B2TOh3EHBopE5TU0IOnTmp
8wXSaps+LqOdjiol8zySVpsKMtLPdKWYsNGT1jIogEqdV8ybdYRjIYMX8Lksy4c8
fZOiS0sSBNu1zgJdis+PnVHvlSLmghGzvoAK89uQ6h1a+U9TgAdFHGNjwb5zFvJH
TG21VaSuZHLTQ66Q8Lw/QKgAj3UnqgqkcQQ8ug/hDyQTFO//CnBAdIC3b+yBrYHZ
LDpXQbAfJ9CiounTFucea3jWPygJnYLodgsVBM4FmzlxBXlYy9gK/2bPjyEX20xz
OJzDlsyh39C3or0BVBbzE1wzrKgw1cjmMYBDr5d/5SAsR/ZgY4iUie+fWtiWbw/b
rMWcHrynLAxxniQQXVPksL5E08JcnyXB0bKMqh4zw01gToarAkftf4TyOMnccKwy
xpKcOHDYwRRC0JFXrkIcb94a1ramwspJE9AzPAlGf63HuWoMSNAqrBGk36vt/qk6
NEsEla4eQzvzqF9NMPakpznfAkj4UdRPUeGWMYD7VO13whKGa2ZECyCBu+8hybeK
eYoDZdz2foFS5FcxLbMpOCKsnByStuimgnKW0pta3LOVeG+RjzxqDGdNhZwg8Czj
OGGykZqQeIyqNX/2kyjj1v8otMmg+BVvjg8pBYgGuT8KkF3CzMGS4dOa97n+nDE2
NMAV+J4fNlxqMYWkxar43mq9OnjkONUla+EaBAi0Wx/aY5aj1kwkeWx0Wr1ZT5fw
GlCEdMA/aQxJiHR4Xue95NzI0cuTObK0R+MoK5cVSfchtzu/amX5RuyPssA1mW7N
0eV8jHPYsjndwT4v6LIgi2tOABZ3coxBYK+o/qlNQS7QSyGDIjMER+/6OwvWHOvh
DN/pldrJtS+lZEa4+LPMZ6pN7gaHpsMsXU/FW6Csd3aIhtBOI1KLwfwVaNp+/vex
F3mzHfUMXfugZjcjxXYoiteEvYENM9hd03L1z63kNZ4/7f22rmqaQ7uutzSZ/ZV2
2zNfLDz/08gX17cXW39MElzCzwK25wYzrlS3wceBWmJOhNQrHBXoiEXS4n1Csool
qHKZGNtB0bLtlixmtxP4YXWjTJe8Tfb9EzbMpvHoOuzezHR8FeMeTebkFWb6wkKY
BE6UyVlgRCFEmsU2E1RqLOrH9qTHpvUVoh5YPbDfHRQlnmleNR5dV0orpPe7ty4/
9qPhfdwLnmGpzKGCwFcIwAq6D+JNIr0CkKep/CeI/Pp1eQtP0KIdl+q5NYQpIm79
V5QgTH6Ys9AXnp+QHeQD8bTpW+MJJxVkHxhWiKV0cz+se81/ZgSfsNVxNQjHj7lT
xta4l3BkatsRFYo6IC/8tG9gsjF0vk3eJkzuyu91zibnYI7JlZHFCxUQ4ySDTnbx
4eKrrEPF/Bf7tlSPI/p2zQWvl5fR5sHj1X0hrA19UYCflxKxwUH1cVVN2asC79aP
znpsN+FBdkgYMK1NvJs8UNUdALM4p52S2S483xD/2kw1V30V75/9OwXsEhC3AoCt
6A3YYbJv6wqFkweHSdyUXgljoiLzq0060gVO3wLdUaaGmGqsncf2kkWUZM1jDvlk
UYFMmBbTZ1V6biRsge17pa/r4B/wHgYDFiEmZ9JmKSFWSmdoQWbj1ewIogmPSG12
npytOVS3OWeCJTEGEOc48OkBu95WQ8//zuZKfUX5BajiSIt6gNVo4A21duwjxNLs
rcDg9lbr+Ogp5/MYRb4jLKXZs5UxkVZRL/E2X/91+2kVZQbg3tOJ6fC0ZY2HFZZo
+DYJmnL1FAbOuhTO1NCwnhbp88QOIiCCUi1Q4FCa1pLpWGQnRfHbBojYdk0j9wj0
t+2j/x9XNm+YoUNP9HTBcWnVpXAzT8ohuN9YyzYqUBdRLaOSNJCZhXhYVqLT99Ol
Egt0z6JQSby+lWvXUeVr+4cXwqp2O+LeFGZyyk4RkxgsDlh4XveEQmLf/UCR1xeE
xs2FJY87ULPbgpoZ9r1183Y+VH8qaAOV7Q24xPpEu05v58EDjz3by03cfPJKKvM3
As5ArSvZTvvhv/V0F6A+sZpACgXzbA+563od48Vij9s77z2sCNwIGUwXFo9TIBT8
B1S52GvIHwS3SZ+fb0klYrUY+U5J7OXE3riAWZuhfEg9S0BkPzEzH5JGbAgNwKkA
wBQMWsv5gU3BID9dlE8LvEEHxu0TPCltc7RSOq0CdK8HpmdVRFyHKeTZnlUmXDqV
pqNKa7BSeF1Ha79POmQHkG+S6cclXQMZ6/WvhbnTxdtd6RWI6ukj9dHAIQT3oCiw
vqzw2I3cTS1KK7QJHBBs9JeaHRqw4Hz7N0Jpyq4NtJjPyPcB+W7ekNyzDJMyZC5Z
3vrqA7peub1b4rkYYyoK+2Pd0psv6yVAe4BcrH6u8IhBg0U0iMqJleqAocxBvuFr
13Uh05DzgFCroSkh3GVXOk/1i7xMADbR7/e/yUspu4uVk5ZjbaqqbjFN2DRgDEaC
/1kD5pk4OZ1y3VMHqfaW3ZPqdwlTPiOc2uz8tKwblFGAhtQDXUiCUzY6JRmjJEqP
rmi1HRNBRABmuJRlvBO7ZoSYzjq48fGUkMZ0aLlo1mylvkQLPwGVkmB7o9HQzVvL
UpACIyg5mtGO0TkHnN901IG9eK3guvZgEopQdod/DTPzKAghq/we9RLIl0kTGXia
9Er3qUZm2js6FLqmfBB7jpZnmhATLVoRK8NmkkmzetNmSCFHW/Nwi+/gzvuHZgnJ
xM1kkSItSX3FU5CNm86iMpb6XHFpCpULDEl2eApHgzuxQt2uNnhP8GU/vZmVFVlK
lorCMrBkV4c0A/9rtbl5J6QUNdLmOOZ8g+B2c6sXGzcCQw7FURdDsd9zEnSMvJtG
BYRSXg/qcdssFFFPZ9LyvMZxtILy7r7LJSbFjyny+5N3bYirBCAJLfYK5Pdvo0aR
M++79UXA3+4TosypakhLuaByug4EayRELdzJ9/GI2U10cMIwTV7hozZ+kYXnuvHr
OgXOqIe1v2g0poUnPUQcspgpSbLXyS4f2vxvbvjH+PcroCkp2aS2eT4bsC3GHMN4
7qa5sG73c/zgAUbbDA4ub4iOlsyVsglslTjQa724eYuBAa0yPNBPNgg/GAE1VFzC
JkmEB96jvgriasYFSczB3x9dDxby6hFoJsvQC61XJ/NLCUn+y6itgbxiTXs8dOps
dd8QwsYADOXT6VQ8Vywzebzs1EUBu5bIsmuCJG17dsUyTCacAW49DQ2RZpN+3622
TGI9HCl0qStvhnXifxTXB7+U7ljcwlzKCbw2a9J0xdst9MX2fuGoz7UrnrS+/l76
ZN2OtsWsFiCZfEE4EBP8FcM/n+fSrmEzJucSWmGFVYXwnnVG1JBZzLczxPVbmutm
dsiiU5oU2nKrmeBOhBYZQYb/N9y88McHAqkiIZpHkGSiWF3OIM2uffHQQGbS+ALU
AiCVuzx1PNdT/PtExG0+RPFc5E6decGhbfl4zy4DTFQ6690y4pfFsZc/EL5Jvi/f
8uGXXZ6SZo4zl1E3uYHoiGHA7iDh8tTKahWul+TYZpbykg4so9TfgX+wyRCBX0kD
tt2xMB39BT1wSXTx8EYM2cCGHp3HsYY2hbJOkUnvjFT324CQdbVksi0OW6+1EYTC
27ej0TrUsH6gfgTWeRrHXJCMbXLgmva5uXA5FtO2acm5hb+b0YBpEWRzw16zPYVb
8UPZShHc8FHWM8RJ5005elU7o3bh+pNMfsUZ1BBw+e9fq7KH5Bq/zgRoHR6QtUdG
rVgDLzbx2vj60BLujeyhfTvdaYDS6CoLmNobrnizlJCj5b3CIqdFuHAn1G+MBkuC
au+4qmVDQkqNcIZPEWr5nebe7QRwXa+lJ+5jzgDttpuyPFnSBIIJypL8bSbXuqLm
/burivs1m+/bY1/XhS4KjsAyajuN0UudE7c7JAt15Amy5Oi0gs+8rpoLTk4GLuCS
xUwROaTUVk/PDcphH0A+ujmQ2nGBuWzxHAW3Vw0vqQ/v+I//+Okl/yr27HgDS9pr
67pER5s2do5pu5EAZUhOiPTvQdrfc+740dw0nbAPVtcXMdtuJRIjpt5Bmi9QJ6wy
KGa4d22ftUmd3vkWEgBXNdlmbLJwcygSDaerpU/u9RrnKe0jvGXmVrcKQD9PYiEw
VsYFgrUYnvfRQfGd/3rJGxWvEtsEbUONdGqVyXJZ02pbwPrRUEFJk2MTwJl3+/F3
SzePgFxN070ydfSPMrS0WO8mzWddIUeOIF5YHRG8PIamJpD9M6EYtZxbxeTm9Z3k
OIV6yFy5l1qwLuce7hqSYOm4ksU8we+ZDitW8gcn3tzEyXVkyYCD2F1hEdPW30ex
G8UsyWPSSpUPT6uPoXNXDdeCOdc3JzGgPQHZv6Pz2vZp+Ius3Z0T1uGZjw93y56o
wnOJ5GpP/xrKpCDAuLdK0gIgYmxtP6B58G9n0QR6Ag03Y2RFhTaWILwAqI56LuQM
qFctup04bcS2TJypCxowBFbbK5RwiLPLjzBo4H9YbHkJIC1agtBDf7HnD4t9gv0R
4wVPq135tE/B3WIoy8kAgAQpaPZkxiCEsjPHF5wc5txcZ30pn0arFwr+VXABlBrA
IK31Im2UBdm62EwGtqHIXCJV3XLRgGapOUMa+7MGNOJxnlFgB7Dlk11LcigDoSzx
umNHkGdnbeqXfcZfODqrBAt4boxP1n32B1yaOOGubkQm2cYIJG5egNq/bRo4SWmT
RDThbQt/QbRXwSQWv0sau5wD+M7a5gg9Mh++dljewguh1wfRqqeRnHB16Bs9i8Vv
uSZTdRbT85VJEeeP2U+mZiXwCNaoFKZPkdwbAGMyOvUTPGpRpK4waLHal89UT13e
a8nvpSSUCZKJCeqMr29Z9yolIHnWBHoBUpGiEmUVBl/oCRMF3llFVRT7yqCkmv/G
cccP08odgilDRjzbHjaTqQOKPBr48t82vvyzzHk/U5D/pGIhr6iOtDu3gV+sgyaN
k/Z6r8jvWFZ7W8MIWh1aIGykJAED7rtL4af6pBHWuZiePvY000cbsOm2ItOOabEN
b4zCTTemr0/REEyYPgb20X9tDMG77eKDexKb1n7fkW5n6LIknoaA53YwsEBunaBv
dyphbmf39kMR0Ec4/BHe4giFK4TGtpYScHzMjyw6+Yg8B7Pv4g4HmAw/VJD+FCsV
sO3gaZnyRrCQxi+TYZO3F+Lcs8/ZlBTOZS1KeVMPNCBJkpbfHvDH5v39lvXsA+qp
N8+vi32ZFVOfTD2NRUtlbPbgM7A+71mvfdOnF2MIAPIPaczNy4ISo4aDcEBZtcSv
PfcNE3XBk/fYVeNQhrU/+L6OuePaf5NRGfIuc6vx/qrY/oKb+NiTyviQVr0Oszbk
UaAC8pFZ9Uql+uTqQTFmZ8L8luAqM2vLk1GYuVjVezWQmdhsaTSGVJ0sGaivC0r3
grcA5XkEMlS6V8o8WRs0IQLuBndmIGFBFfd8jvRqt99SzxMZAPExKqDAZNNHVUYZ
IUVJqOz37XjU5aiCtHWIlTi27bO73omnEQbB1vlJPF3WkBQ5ieUs+xlyoSndbtpR
yLJB+zt7WCcV9vv8alSv/sGyx+zOdUit2zAriVUcPircPmmlFqPVaaEPBvFXrMiz
SUI1ZxC4zw/14FzU43Td2b041MY5HpIEHQlDaos3Yu/OMnwIakQs/Je6M7dRGW8E
bznA4Owp29W1hXFBdTQZuHK3b5AAjO2/mjzf3A+RX7fKdekD0qifVIh/0HGKIv0E
bSEY4q1cFoXRYNgaNas5dYcqaAsCRDZsQCb0FhK/Z8PK08lKUeSjfAChPXeQ3bSl
emq/41CyFsW8n50A97ehyYzBPILmRiANKWc39ZahV4eenCTdrO28SO8b2DNQM4/6
XTnNkCY7W+XnSvCbft1+xjwy6ak0yXslhPHLYtlGSIhRxd9Ik8fhBY+dJVOoosbK
aI2sLqFgboVpzCwCrB2fl1WgWfer41EBVA5gPCSTv9NaaxwUa5meibC0jCHKWBzt
AcO5zlsqp2uDGZV23/5o70m6sYPvrqDIHvqWFtPGS/QnGuO1tW3+XaOc71tKVK6E
w08hOgwCvRmBtzEs3EUA2B55NMZn4Wo9q60fY/mpOuZJgONGTBOtw6qoEqnE0WAQ
B9P/6znI7Yh2ePaxJQNGzPYzyfkOmLv6y/NPJ0elFu2RgcdSpGf4tQW5tL1Uz26H
fc7sto6NfnjxZ004mvzyC3oOiK1d9fUXQqpeGTvqzZrXhAtzBeBn/kDWR3iz6LOW
9VDVxQEUKQnevfRYv0Y9S17kUo37Ew2Qz3cgnAp+2yuBvLjBUN6I19AakN3ApvFJ
rTX8LRazjrgg2iAc8quLhnYUdHgr567CtqCsuhlbeZXNKiQ0T6BYE+kMNnnUZUU/
2AvnxeVGObcn7TojMLMUTiDZU4sKUu6lnlw+rbW6eRL+f1NrvYiioyKdDg6DBKgR
9FeU//ZUwhRdAd4WrXN5vDtQUxItqo18fkkX3C4GUz3Hjjo9X1uv8XZEqz1iMdTN
4qGYEh00NB/OYq7wnRCotTs395rzWmyYUGv7WGOcewsqvR9TxBfKWD14U6Ff5f3A
L5twtFFL65ZCwLT+KZTT1aLpdjswV4YJMYVf3sMHS48Lw7aA/2ZpjIEGs0Qrnxou
acA5/A2x7cotK02pL5RQZsTuJXGx0fYLM6GPylJUE8seZT4mD0U9nXQhFhPko1KA
kTlz5n3KUBKE1FQnorkic3/MDxMAs82on+16h9duja1UO3vtGUzh/hSDBnMnuFV5
jsxwcVSbRGpRZy4Dp2ZIYhPHQjVNNovihG5KzUCznykX1VCxN1PtZvyEnL0NfL0n
PBRgU6IlpGJZ2jCGtv+PKllw8fGOa/S2Gck+qHNxynEurpEj94rBos0c0Izi1Frp
eTTovMHXPlvhnoqRxL62VVOXY7BpZ8jBZomIY2oxl0+0QH+A+Ellf80G7zj4p3k9
F/uJwwM/aPtx/otWZ3FTH3bnw2d+fMX9Gci18iGuQtkv7n3wlSow6PQjuJRHyf9a
AJzx00MCYC0SES7MZcq6AHM9GmsLNSyV577anLfdFpcsY7H3Ou41Oq0eQy3vyVWO
k/StIQfjDIrezv2Di7wnChsWhJfduY3BkX3CNJ8b4NF72nZfUqwwqSIss94p1D+4
b4V/V2HqabxFH9p0JGM54/oEzcJoUqrR/YNJ6W96brJG2xkYpaDlEbePE3D/Cc2w
DyXBmmHLS0UvUccNvaHg+BZI9VzwOp9rhy96DPrsABPOpuH9VLS3IN3WvSPRKx3D
rNUjYowRSANPnZDWUobFrdNPM5a4TuW1D//swMmJT2QRRY1WemkaejfWwCgiKsUV
5BYEzgYkgjemw0CBd0x7Zc2442uScmMZjEUaorhftFHxsHx5NbFiLaXpW8JcHHcx
WGbyga8Pu4AX2jEBX2rOfPZR90uWIiK05c7Y3TvFb9w=
`pragma protect end_protected
