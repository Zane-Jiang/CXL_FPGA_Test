`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
OiEcW83D0fXDhoh9jEHIlIjKi1pJvYQbruVRcGIhPOhrn3w6Y7zzDDiahA8Sr7tc
SfpYYbk4pJ1dRn3j12kohnlGqtkFceOjtdGpuy+k74dkOQB7n9vrv/i4PxGAtRlj
y7eqG6z2BX8CLRx47Ui6hmKg1uE0lm+yOtNCVBsTfME=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
OPMFPXzyi9HI/LnlV/kxbnKuxmNIq/Mx/Pej15h4HpiPbayU0FsekBGEtJAVwZ02
PKfI3xHMJ3urX4GTmKyLA2CQ7bZzp+Jid2WxuUy2EFQ0euPlwCkf8Jytp4obp1gq
jd9NfXpDrSdH3xQVPE9ct4ZmVD8pTq4zO2cTY/1hK1DirqcmP5VSnRi/4o162rAK
DnvrS2061Egsa4d8XR8fBe8vH0GutP9Yv1A/eD8w3XGud9/aTQ21Oioc0DZRAg07
mD1Fht4nHhUr1Tdt2nTvkSYyboInmCXDrSpb5ybO/FbyjHDb7O2XrouRAYimMWwa
I2wv2bS7ZuzHecdMEH7mc36Bk19gU66ndPHche3Aip8+PfXYqITp/BEUN3mNtszp
9ILeb1UFwrS7qhLe6awuY1RoBUSN/yBKWzsHVss+q2Ii2AFb4cnfuXpRXfTT0LgB
E4L37nVIqtQ0pfO6o/js8qjCuNDZuUsTNgshuC/31KG2MTHU9RKKHYummqwNpWkK
zJmQJN4+DxT5Hx9Q9g7il0SlWvv3iOHG69/BOXWgBAFVifEVhVCCi4B9+H+K/QyK
fG/Cg5KSxn9/67kzHMk38qSRlNvFlASq6qY4Su7nFRkhxscUhBcnRue/xR5Z8OOC
6ziCQ8AH2VIlZj32E2qNJDirTmMx8WPzZDSCwwJBfdd0E0mDdJCDlHUqN0Lcuh5Y
yENTKnJlec/ph6pKdZtaHaJlGcbzUlyzwJg1zxwSlbgkvIfSKfJcytXnZqwtJgGy
05F63us9yEdSjWhlc9XGC8w0/0nDaDCpOF846PQOj1a0ZaBMnVQoZIrN6W98K+hq
xSG/EB2h5abyucimZos3NEQn6qxMaEWWEIv2+ry7yMmjEBerX+pru0qmaX/f1XDT
drQ9Rz0HN8tO+zOmXNOg9QtNH7y2Fx8IU1yFTbS6mH2tXDtrsYWViVWyszHMR/1Q
gRc02AnO68VGQR9/5IjCYgX1wpSaJOn8v6pcFYLKVRlSiY4gm4bZs5e2P9soI1EU
WS2osKu+Xu1uSfV2vwKnllLMuI/elu1XYM+GQzt558e8zTBEf7H4WyROC8m7ostM
atVh2V61i7OzJsGsAym3rL8lj0ZgUKSgA7cL+SrmDPEg6rEtXMF4B/QeK5aqrXei
0i66oAKYsiE0uiEyZU9Hr6Uk9PS/+NEkE7f9lzD5nbmSnOa3Pu251ex3QDl9CbZ8
isZt5cCwja9JbtT+pFelnQJ2/3dL70CCwa0dtf2wR/8V1AwFsSwlhnXmaFb7RvpX
wsNiGjVXjm9RvzOs6IhsCd2FEBDJ5hnPIDDbNmA5imM/8/64962Ex4UuOKJ/S8Iz
5DfaVnwvGekASJh9smqgtO34IkwOXnAw3NdSj3OiBnzgCbMK1V5nQM4F2MkxV1v4
XZyEqECw7FaYQXdXzuKRHZyhaqU9wgTCTrjk3bruvYeDqmGGLBj+RStzBbXap577
DRR5UjGiAnYUg9hZJP7/6AXMuuvd/gaL2VVAwjxC7y3kcSdGinJUTA3dtUZUpuJK
3Ky5Bko3LiSDUkq7Yt8P6qOLsPV4v1UIli9N9Loj45CBV6L3mj4PPcNFxjqTJivY
cFXsGvf2XJZV7UIsaKLS4mEidi2iM7qSIOui0l29BztdAxrDhB85xaf/kJ4siih+
FjSgl8m9KSSnwQtlkP9z+I7tpDRY+2norJLI7vU3jqFQqdcz+SxRJOKFgTDyCkF6
cmiklybD9ZCc14Tt9TuoRLT1CUdVn9udOouS+Vq+qp82YVLS7+JVRHvOoXTnRN69
DZ/GMTVDBfC50Cj9Q93bpJmIMgtbfmi8zmkHr1Ex/wgiJ80SR4dPNX3/lW1fitph
KTJJG1j/wfFloQuyMJsjNwpwnZQ8CKL54lCd2xhyf/1Y3ALr/subuUm06A2kVI69
NaIRwJz1yUTcDxd/tiTyn7BRnu8oL1kemsviiJADi8Dlsdu3oGOIA/DKTAji3Iqj
x6tkeDh0icjrY0n6F20GtmGBCCo4Y+59Asy2s5v++G5NjJ7K36FDqAXTcdvRLxnA
iUX+xk3JBbXCxf3WNpMJCB+hQNiKxkSYu3lMi7VJA23nGDOgWXKsCMq48nkCaQIF
feIJpRgWPph8zOtZRK5YbPGSd541AqfenBi0HGlm4z22jzbbKykNblwsh6MIXMIS
9kP7VOH2yAFcckd/h+uvsQF4xPLUmNQUdXxOVU80PI1GKaBqtlMwpM7SSzj8a5Ca
QuO7Qg1TnSn3aFa1VRc9HCwnlT6fX7R7OnyupAbWUu+umxZKX2pQo38GW3buA3Wi
tt2GoSob7KSDQOcljCNHXFhCLUo6WSkfhOmhxjrquR1KgBXDtM9E5C6CsgBv1yea
sPpeFTAjCuNKZHM2j+HCbqT2Z1WjJtd1zn+l+7Y+pTCszpGB132ZGkm/HHz9YsYb
K6gYYQ3CkbE05Bb2K5xdA24rB9eUpkRsfXJugdBQ2F4sUzIqCXaYaannY21Grk1a
njU4tewX+o/9Lrg2J/+PY5cojpudxdigi4QVEL6uO0bOLi9OjtoWU6Y+ablvmyUt
1B6Mtb2xfY7ALzM+nlUaNhhR7g0Vwds/OXHqh5ukIWqKf4NDxpuXbTBDmkK4n8fW
VRUwEM2ObNlDzGcJYGXXZAKzpH3eQ3vEhU5R5/+OF118C0u+lj9m1+VNV8VEhy8x
rYDqn+SaGEsEVjJUBs5mYMdE+LE0GGNgLMFc4Eee/Dv8rv/ql74uk0sZleI8yzTg
UCYppoqFlF0ld1QNDqcVBqHnCAArz/MHnLnKNKfAuSy0YSf6c1XSauIb+NXkp4Rz
BT07ItUGW4S4x0/eXw+CYufoI1TxmrgnEvTYRyDqQNw2sgKwzbK6YHdl+BG3MNR7
Y1vs00WlhyoK8RoSLxW5xRZTVyczftj6V1iuuzu6zlxyxTHrwpMIrVpzTMMWuKoY
dc9dQgUqhOfUMbL/4x6XmF+og5No2/V/WQtBVi5/yn9Wx1p5W6VjrHTJeV/94qvL
fq2NLdz385M2XvOTX6yyDiHxE+k00PeESYHnMEL5XnUXrZxjQXeneizwlTTNYF3x
s6owmZ5zh/mn7J26qgPseJ+fD7iml3lMn8eyDxqxvTRYDt9b/HSQAsTEIW/jsVBj
p27bW5Akfjz5ISCfnLQ1CJCaZ+J/BJlqQ2cRx++0B1yYupHrVo71i4oszJVsiN9p
hMdpOLUgugdbWMo0qQfKroRCVQWMW083oiwFAZo50Py7YU98qegfr93SN4Yg2ggp
eaByh9ExN6ecqGU0OOa5wuEm0XHqfcssyn3MIPI1BKT3WW9v0dIIrg6Qlahq+Gbt
0QOeW2LmBeaM18by3V385kgPieN6SJK/0tBoGKjteq86i0bBXi/GGRRoZJFAeQud
Gscrc6Bw6R8zNrpYwcAW8S95MHgNQoBy+h1LkzItNkPoJlJrO9acZt4HbzvpQPTQ
rjgRpEIlFPA66CT7qMpNgivbv1/zmaaWN7YfBIuA6Gj72Y/BO90ICLQkujcT3+wb
XpM1LHpMwii4q6oV/vqwyiY+OBY2oWboBFSC3cNpR9voHDce2WmPrXVTJuD1Wblf
owMlt7WJMCj2Yd/px6scyl0qcaqccJ2h5neBLOL978Yxy1sx5qmEwidxOEGZdXNw
PZJXnJrF1EyLbWlpB1CoJ8lXtwOkvvSL9ItMDH84qe+gEmkx/Mac8M0J+6Yx3F3X
SUNsuqy3BgrpexQJzVl79O7dVrTVMwWt70dm0YNpFNyPEKI7/SazYdDmaS/mYibA
/nnEpobak3XraVzYEJo/vuWkRSVkNBhCptRq7vShc6Et+sNlC9xrtJpfu3/6/bpx
UiCj4Gjubj+5TD0Q+6VaezOWReVgzZzwDb0E0t0hkiP66EMKlOo2Ipr8c3Nu+en/
aaizNrSd6CyvKpr4ius0012Bkoj9e2Y5Geeao6YNgBHwgHe7gPWBYNVE82ck/YsO
xuWEZ6ceCh8Nkyk4zp7Y+FIaRnIm+CSJ2mPaaTpenOZ20bTxav/kSzLGeUtQBlTV
M7+ecL8CVARlNi/MskhxaoKc8TSHcITOAxhpP7RpDIGlqVtqR0KSTwq0uV9SAiNZ
Kpiq/7Gm8z08/0qmLfiZXZvVTGZh/mLHXi0185XEfA85T0S0MVlNxEjNA8QAr18R
D30VoaBsN1d6UlcaQJfAnbLb8fb0393psWrbcj8MdEFOiO4ETyvKr8aPw46UaIUw
eLE15SXNL9AV7bg+UhSSeFiyVcxyMpvCtq91tR5Za9zYE5RXvGRLrVtjuyiTOFeO
DtodgJqqvg5xRX4BcGKFZQdDNIAF/UsMbFskF4KSKAmTE61cwUjVkKtpO+kUyA06
tD/YXzHUB2N0MVOiPX4fLuynUTQw2oS2+qOyl8WIJJgx8KQ7HeIrZ9VTxXdYEjgz
EJ91mGeBdtrKv5u/rC7zIyDc/kOUjVMr1Oex2Ba5X/RW6UdY4HIYGmJMJuhWiE/K
pWrog4ea0GtRNK3QiQ7vGEzXq0+ZKZYNPfgttJ0fcgFh2DozlsNf9LFx2e8WaKEZ
cvw6F8ud+QCgkxQwRS+R9/KqYFiSISdpKJZ2ulOC/nYp8aIGNLGKendxtahkHGan
J0Ch195L/M8XiwQ+XblmSHSEUXnt/lcDBNZyUJuP3/hGzPhPyplpJevUjGhFi+WJ
0WAsuuaiaTzm6mfbkmVkuSfRvW8Ybsw71YG++miJHkQum0aM7Fzbtf+1LtaVTLFD
COchP1u6xVGq7sjaxl/Yn7IC8/xvTmKjGgeiUaDj5z4N4UWVpMQkLZ8iwAStS3ml
zmJg1ZutT05gRMNoIvYxewg6S65vaKLVNZJuOokyduCr5Ncc7VkfiTLZQJfgPOqj
ILRTk0tL98/hmSUsZCDIhCtLVBaqnU7hs0ASQVc+gktXtX+9/F8sJkDfgpKJEy+k
58YZDpUWJEYXsky8D6KxUBbiKXUhUa12DbqYFMVySbtfgDBJq2pDnfoAAha7yaGv
biydQyNOvs+vpUktrN+vpQ9+h0n0AgY4kIhr9tLR8m9xu+vJ+xkzMFW/tbfJiPwO
b3j8YPXvqVQKedtuo45wbZN8pIamaOSZX9zAWvGn25GAj2XxWYzcSdeBRS5rbCyL
zB+Xkkm1lUatdcDC+/v0wLVhM3w94WmGU3TlbeCzJ6/B3My/8DmelptaxK25zunN
qjWhgu1QtLBve++Ba4dzXnYTm35+FwOO0CpxC1kAAOqpfY6blf92W54LijXKtIeQ
Ue3V5irFb/KEi+XNoZA8OpQXcpB7GkJl6S7aTLKvIHV7u9ldK1LZVyQobbTXt45A
Pmk11HpD8YeOpSoQLfwYcwVz91CK/NbDuvrAe40jrNx4tEiJw42ObEBNHQhje3HH
9lnOCbfGE1YC01pKpJAI/gbm3N2C42FvBuxmL129pHyCtbNRYmQnFUveQVHB9/Hs
zpCKg04/zDfaLyiCFjYN8/Ee0+NQyUkKrH1XULEHa7Z41zZlN29kRa1BvJ3dbA7f
icGftmIL5pWmmoCpE0RcHC/ZlYwLJwhgN7RZmOBPjisRmhex9HknRAVLeeTSYJVR
Pc3ryERIrwrH1kKOM+P0NSW4cXU/E8v0bSDspHsO3XrePHllzVcnWQ1VzY+2fh72
QLNp/8DecSwj3wEQOT1LDAnzdye+hynA2zxeTKzY9gYSdAHlm/yh+it8kdFos3Nl
jTuGTkOwkOVDfgpx1VHg4a9cNOS24AirNkKl4m4txSrXTFr8xk4RsN0zAYgrfhsd
I+5DQsU9rOnGEFNZhbns7jCTw4687JgFB5lB15kpDl81YPuoC1XF+gAV7SdLzlmi
Dv+FVnoh+Ec8O5oNSJetjzqaDgyY8fqa3Zw30d2g8jk7lktHMbDc66FOAU7Ay/k0
sldzbejqOxjkt0lVQwSZFCtAaOUqs8wKak2xHyuZgc2MvIRZQR9TeJ6jmdwrd+UF
0uwXk0wlW5sIbQPFo51P0K7AtZN4O/NS3XdktauelkizL70EJBVvqbFauYdUMj+M
spare8ciHa4DXpWRr9Ajq1/QXbEsAi684XF/NF7w6m+MNGMqg91H4IzJXSwQn8SE
qq6iVr0/O6m0T0g7hjEP9pztoDz/thO0qRBFToRcSVqY7g5wqcFZN8Vx/ZmPLXGE
Ce4aI5sefBeRGy3XXp5fEM0XVhietIKBY60zrF4/OmG78Uy3ZGane9PRDRa6qgnn
2CuUHDX2wQScOOcZqUYB6WER9UxBixyIKNTBfu7OnA2cTzDAAT7dapL8H9+o0m3t
CaXquCxSeFg33aFCaQpn0Wm4EFfdrDTvPJc1xFWRV/nGoBy2ESaRbAQweqNzYcMr
fbp5VQ7mf23Mz0bjl8twa47T2D1sLOpi364XrPv+sVpZGd3HrdhE5QXs71ULVy0T
mF+HgSx4lpmjMjFVlPjOtEtKCVamnIxsN1+Iwgs9R6xaFa45BTiYEa5zlEOvjpSO
4KTgcT45RTyY4uV6ap1JZ8gEs9GX5OPadiOsAKp3edeLJ78BrlVFFONnHaIiQDEl
oXbhGkyW5IRK5+D4hlqe/E/rzqDPKVhQrjCEaUiN5if1waeDZQBV8bkeYJnzl+PA
9bndYpJm3ha53XprI9lYLvv9BA/Jrl3MRVtWDAf2bmuKuckxzNi2TdHekpWbaCU9
LDl7QlkM/gfEFKmeeh+Na11BRLiXIHz9xN9uryiQ9GuWdqYhKyZQEmHwlR43VJXh
IvcKTg3Ws8Zr3eU8ujr3VQ6cTet1huEpUIzut8M6MBaFtaprmhhpYjExtvdtN9yP
sijB89uJ4BH18tg6Wl2dh1bJZ+ujZ8YRWUOSsdijZVUimWJhgBUUiUyypoqpG7WF
JGG6czlWDQ51n4x9wQihYns+ka4ffYZwZtZ3HJp1kjeePq8pT7HW/AB5LHYkC5Md
kiyZZ1Lw+WLEHepOHPmjdsHz9Rs62Hgz+a8ovQijMZf52oWf2M+8U1MMCaOA7lCp
cky+ZvOUwIs37hC56XqbgdvlNFVRTeU0saRPXn2nUgVtlPmQZBJFDkpxAfRrTrJi
9uQdWsTEh3JWR53crbngeDvCFPeZbyIEu9TxnS50CdP9Vodfzw289YeXewKPwYm0
lXMitFLkg3F9dMG+NVgtV2xFiSQ58eHBr+lAhdJJqApFTDWwM+rTU64KjMa/q49s
tcpqul6jknJHCqCHiX6YlQiDMP8AW5W8hdE+7z4+P7JlOVVlOYvHN6NP2Sj/e5LF
Q1Ix46SV4ncrm597Y10QgWWDDYvFfVkvSRTYoK/8ddz6je+ToOR0Q56ncPYjh0uF
qmMq//8wFv2NwDiRDmLkJAQNGFrzi0btBGt4Dnmk8eHByJniEM1gK0s+1ueqp7ai
M2y7FvRHtzPrIvFr8l31ZlDgkuNSAU8zQKbHUTUKDQdEo2YZaqAzSntq679KTtZc
+5cKNh9L4tklUH4xshVwIj1PCsB0jKzz1vbXaHZeIrbDbNlzqQIenNZhQUlA1TVy
tumjfFLw7DQhbxhLimKiOAwncyq08vZmSj5ux6pDXepHWmI1vvh2yPZPIT0GQo1X
fsnH1LFX0gYroKJizC0/3k7U4rEsN+7uMCCtvwNsV/e02mPhSMsWZa9aYYr4mG89
TtNwqEEBm8Wsos59PN91jFMEESIgOxcy6F4v8tHI8Dv7OR45Y2KzdiLF9281N427
tyd+4RdxgGANYlGAABxrs62+y7RyA+WnQ6Vl/WVeyq8f+CfoqjXEmuE4ewNi+OpO
cYWNvPSLJIvRJPVDSCDRfpegtcQyv4nEn1O04372rK3Nar+kVim9c8lFitkiABc/
H+rANiwJzSuUdkWpYaAClxv2qZYTAasDXvU0x+/laOdq2xSZJtwvc7UD+sa71LFb
0DMbZPgQjjynHWwXyW9qLQ4OW4OMvIo414BMjf3sRv2bS1FPehgsp6Pe8u5FQf6N
X/HSCdyquLn3eU8IBvkdhonlh5EE3Zz9lFX2Yu6b6ErNh/oscBoM4gaYsUyUrGJy
DaKDGUjGdubr1uuSLV5Bd12I0mfOd+lsKANvYxYwm8v/b6RGp3p0cSZnuKsOhLjA
S46UnOjX7IX89V8VEq5a2sf7bdgDzKjkPqwumC1hXgkwsE54e2MvRZRsRCYYVCM/
HBCnGh9sOOTK4vEgIMD5irHxHThyj4GJdDQYdyyoNMbkrL4x8VP2EVkwPtsKgVvE
hM4zZ8bRFdJiLlYcRcifKC6DARpbZaoTHez/xKeUa72z6KZjE0MfUqNtxc6xMbBt
AjxeVmcDO26YCHUUGYpWweHwszelTrrZ1cqnOgbmrMRDFnuWTxSWXEHNrKU7qwXy
HfB5Fk7ckMfZwKKmmz7BPeXBGtt9gLjMvTtv7/R2nN1dargoBFSG4tcbCDJV9vFq
XD1HjNMEbIsJDlfzRcjsFX0YA5W1Ts/h7L2iqask23lj16ZcYwzEn6RbWq5mjGeX
JScWDxqyM+NQsRq40945U0q1fuCyRV5KpXMEWK51Im8SsmEHTvAUf9Hcomfez4V3
ozaKopugOnecZMsLEGvLjJpRabXFnTE5Ex5OORVh9Oxx4jeStQJp8/M1wnsJthyH
EirwY5Tcu9LuLUO7a+RAT+MSDQdvL079tIC8D4DRxq5gNFIrji1/4jUAFjO7RGru
YcL1ECXvn2ux7GGkfY7OdC2fb7EgAhXRxIhwYmzpSmYzPvBZkRVAdBRTyme6b0iA
E2S5UyR5o9yWSCiG4NnQgMUJLA7tB56gsyr/FrY3xXA/oAOCeoy1irRHSzdRvftP
FuJMl+LMDHf2sMFRywB7RsCbMKB1Af5t+vkfWkAPlc+Yok2ofLFv1JSmT+Fhymzg
Gb+7R+DgFX49YgNfnGrj6ikNcSbfkjLUdTSz4fKNv8gUsefWHj24B7e7FaCDmCpu
0U1Nub6dipKmNCwBqBmgkmOgfoGznG3qSqHpQmdbY/bSXm4wn4+HFys2QaIp660h
1qlBGgW78Jat+vluNvRdGlZY/vZ8kIxTFdhAAGq8t78HPsg2EP1tsjE0PE9Lit/l
wURSDn/KQaWmQzEOAO1Vhe2uDiiAR2UgYYjNecDIbVi8pP5kAFnxPC2jPxvJK2Dl
6DTWM/Hgkz0bth15cmCUYpVzMu+9sMnwvqFjBZBItF+XeZnzfN0Vmuu9T6VEVEuN
ncmaYg+8bQkNPZfWsm5pYUFuorcJcg5LVXAWJfs33JEzyAjwpDexyGxj9e+iN7Hv
QbdOoTov73kbSZKxC+MzOPqUh+tTdrPqVJz4YETZa39+Qb8x4DlHgZ9686VvRb2E
CBU95kn7Jrm9X+3rzQXzIpl+l1sjuPqkzMRd52ZziltWcmfVHK5Lt3iAcGENJOMI
eW5KkHVMMzZGUDPPJKn95xhUvUlqyLKiwEM33M8ZlB1nbAR5rYQXFhx4P/pLs84l
MMrXC7tfmD0in5BBgwgPOc5wuSCYrKqQHfZZ/yAwMUA+lj3iOsfiSfpYUnjd+0BA
q+pK6ITHR8GB61cCgbk0m8qIqgL4RN4K76y6dxr8NHIXRCOZb7Xt7E+mMvKvAH4T
oIXaw5cE2frxnbSsyPHAlBMdVmVBdiZ20JroFyAaDxgb9XIChehmgGfMFTpEyQ/z
fHa4NdcetOmU0Lqzk6oIXhk9OlN2tm+fRSHmyaV1IIh3p9hu/Ga3ieq8vJ+rH+qg
Rlx6ht/Upot/A4XQYBXPhbguXFLi2NBJefbzzG1c1FLO/Vg/CkZNWZSLqb0iwfm6
zEG2djaGX3kDUuaFvgC9sMbCbwvNNgbCJWbbZuOnyzkyURx/iNIS9UBGsONE8ny7
tmNgmAjbo4GSGPuyQ3ZNykeLcnMc/hSx2sMCNSpUzHxGgP/BuLGNGq7VMc7XLQ/x
U/k+QfDzSwvcJHd+q7hDX2dA4B/CWLHhtEpa2SBl0WoExZdI0Fp1Ow+wc2+UsqOK
8FZnJiz3SJ4TNggzm2yStaq+eRZv+uwDNOPIDDr8GWbLwRKk2T6m0PesCPVEFq+J
lWN1LLxrnBXqc6Se8NHypcP6MYf4cok+iuiERVA3uzjzrxOXMygUtp7WYyTx6jMY
9B3m30L7PQsWyYMx6PSaz6eRACnr28J0MVJ2kwfZnsutij35hWQf3/exRUb9ExKP
QlnPDhtO0lJFJtRZYe/k48VpSUhnyO3VQuRp5WNBWU5oAIitY5Yev590Ab4yd8cl
6xXG33aLjnkT+YfePB21jpzY1JTnMz2pLbhprhHTLMLXjRv3T2yUI3f3HdGOB2Fo
2fIsORJ8xbFzCE0ide6SjDeyfDVcnW7DhA9Gt+Zm+O3EVbuRhHv0Uv492HXv7Hro
HBKpZh+pmGRXz/psRGgZ4VgOh/YC1nnGb0sogVoRqw/tL37+3BqSJBSM7xNXbwaJ
PjlvyP5FYtNZzBMzvdRIfk+prOtbCAbA3hOP2IMO+/+3daNGE6QlaRiVHrRHWuXm
CsnzvDQS1g0fvwAF0phrcJ5mHSXVSKgODHZf2m86RqYuCh8L3V/ReXmOR0/uwrt/
mkkx56HcBvuXP+9ld078LQrr5RyHHszypV/z4AZB770fhOCA7WZ5ztzkkv6ZMzc6
PbY/IRdt2XeNU8mOvyZ7zjQ1CKgRkUvdcMzDQ6IbK2Vuti2hIqY7V7qIvIUXhWKb
Jdye632ZZHVkmzLboedI70yJ/ngs9/NwvMT8u/gsm25UF3+bW9nIfQbfYDjPm2VM
Hh1biQyM8g3b/+nYtnl4kP/ObgOhnWAmDXPqxBPIBogHZmTTXXNizdKICjeWbOHk
gAIplgRjQpSBJMtNvmqzMI9eQrGgiYHSadO5hCq6341bHZNjwzvp29iRQryIInae
U2JGd/B1Tlkga80xNrQOgWIiZ9AfM6S+M2ocuTnptgST9GQ9QgOucuFRevib6OsX
LOl6AIUYpQVcZKzg14BWi51wQ3c2uoiLxPAfkCrmqXkXyKI5pUg8+JuzUd58kPgp
T/eB2+CVPOa1YhMOsfY5ZIBviv3IwFH8Hu4EALVJx1cE94sjxFCB1+JIIxRBsqRk
F370WziRK5kQD14oDv7vxqHTnV4v173wZtEOSLvinB10MNgSit3NiWsmQT7AbcP7
KTE/tiTtWpzMqR+0Dsz14nt7jjh7gJCAB3mPzSKhSAtQGyQ8YEoKyJRVCZVx1gDr
AF5Ddf6P+p+Zu2AcxPc5LQP4doh1tsI5aekAnxrm2PG3dGTz05pCqTRfpKZAN9Ff
ZQJq+BrVs++iIrTkOn3zpEcDqKQWMK2jvhA7Pl3GyrSo8PBCqc373g1bLkZWvCHd
27eAU1sHaEW/2Iil6nzghgvsUPSibkENzKHfAB6lTevmDGw2PER7HbOe000xML6o
ObXW619mDwARkqYeZS/8u/hVRA4S7EnlPFHkZPqwJSGipnOwo06WvdVLFcKNPyZ1
bZwyUAHdWtifXy6e5ucRUCgaaduS4DecGn0BJoP7ems=
`pragma protect end_protected
