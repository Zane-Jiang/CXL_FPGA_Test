// altecc_enc_latency0.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module altecc_enc_latency0 (
		input  wire [63:0] data, // data.data
		output wire [71:0] q     //    q.q
	);

	altecc_enc_latency0_altecc_1910_azqkyey altecc_0 (
		.data (data), //   input,  width = 64, data.data
		.q    (q)     //  output,  width = 72,    q.q
	);

endmodule
