// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H8LvBOa4cQM1Cs6eDU9KAA6uDc79fKRu5g9L1IsECsrf/IpashnEcjFLS6u5
lcx1DktPtVRpluAsc5nwqnDfWuU8OHKqNiQiZC1mB3TXISypp4qgbTQsjJAu
ATETJBGTTUZvrfqNkI/RVDLIf64OMXoygGlEHkQPOMfW9/3Qw0FxXgNl8cZv
+fQW4JpdUYCAqfp04A+7GfupbPe2vMFiGpfDzqgADJgPYKjEF6e16r0U+sMH
/RYhQe//s5BJvNQxLvY0/xMcrrdSSwBuq7tSxRe0mQizQyKnk2oC2csbV4oZ
IpUL7qQwKkq4bekUliPRT0lH3K+IxKtjzdWs/aLFOw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pCLxH9suC7qRFtik7UHYVhLGrw26m+R8va63z2mh7EnSZo78q9iAhwF4Ysvz
dv2W95xFk9pNdbayhIR67ww+2sJnSsENYechIgH2iAJXg20miSI2rXoWVs4t
WBbZDwOcBAO8rqgPoiqBo0qekZuo74JEa92QlwoFgvsrTzuaVYf2tQGRSmS6
aTr1VnlT13WXmAA3nVaWABgDbKhiQuR9BEUgvPAcBIdzhwU9j1VcCogiBtok
NWxqZql6S2O98sSFLkG381PI9C5h60E16FgmAauac9P2FjMQuq3yTKFT9LFy
FZroqGBjTke3YnKbexVIJWBPZ0VhMqj7wMUT+5B6xQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U5kOK5kOMzT4XehwrsdTmV1JRippq4kkuhHixtqO+LdLOzkQaiqD5UDBL84R
TiN6mdopgRwASDKn+9SJ6AL8lmHJZbG1iZvSjhHhZ8z52aEuilPBNljIioL1
fphhe3WvoztScPHNOC7vb4K8xgrT3YrdjRGhUWl2p4jXFP1AaL3srXybLIGp
mVg14Hk1q7Yg0TrDbnt++yGw+XDg70FJn4eQ7DEMFaEZ6B+GiqfZocuBhv0E
RF8DSKnspYNDqE1tKe21/zUubPfnLxfUb85PIurevZXdp/u4JBJWdmfTv/yA
oTo1Ci8YYFUkvFYMtau7Qcfv7xniKwlpV0HJsTZoHg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IMkOK3JB7nO1hagZbIcOKnaghu8c/LPIO87/OTFlwvKhq1ymR22/FPvd6JXj
Y/g+ElZNZRgUzR4qSDD23pbj2npqwfYZc79I+zm4qq0cLgwu8r/KNGhuQRBb
AaWE29ZREvA9pIQ/idYbmSG388jWOzxvTPp+KafOHmUGILe9Z2M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
socnWyvv9rfBRNgAZKDhZKUiei0IuYR110q/gya9QcDr5v+jRgVPKAeeJ9hx
5MeqBWdwxFq1kv822/0GPoiUuQevReg7iGzpwHQV8wKuxxKJ8/Bvf369OygH
21RNMV253FnhWbc4Y0dEqWRe86ARFTztjXf/PMDwOm/5DAEUB7HuS6OENP4Q
W7LTZqlG9KN+MxzFbC2g99HRuu+Qj/xO1w3e/x+vhkrldG99SASW6JcCmWyI
a6lCOTnSyGm6cvA5W7pHQ0EMPzeYKR7z216f0gYLsq4Yg5RQyP0vq5+doo2C
Ug3BzVxVKl3PnFcb2YATfm1lva7XqZtaJerPUbwVTEP1jNq/Ozt9qAzUxAW2
rOT8m+B620LgoKSiddnxjovcgZoABXsQa+u1zc/sZzOMWg153WmPKl7lp67l
dBcgGcQtfsmjNk4JIVKtTsLW9uqOukz9Sg0FTa1mtIO8rmjEF+Q+Bd7hqEC7
Pu+IUkjmL0ug+o/vHKHrToEKK8n16zEZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PQfv9ixLzGuQ2gW0enR5597Vykw5MVyX2ybRG2lr6pWpSF5NFcGzwl1e6eFX
KnlBtLRyGY3iYzlmiF6BP1Nvh1gR79WIxRlsPJ0DYgDm8tmIwkVY+xrczjr7
ZqHIzvIDkDOhKYmTG5cc4s+CQEXEgOu0+J3g0JCnl+W1/YF4de0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K6zAH2mKFu2iUvHyd6GxlAayCK54zkOuyunJbrJ1o7d5PA26yM8jEPgehNmJ
HEl17XHt+etOHpgomQmWz3Dct2yIYxyKlOKkN7Ad3kmYjajKC9SDRgEsVZ2d
GJS876OHwn5CD/cFs7tRbvWyHZjiOhtQJIGLGzRvcT2S5l2LeeU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1392)
`pragma protect data_block
ZyoS+dsxp+WzJnr2RGpDC7f9BTsW5kJulfEcQLztEoOhaBixQsCwcdckpDqS
HA9uSrVpwyK+91ogzbje7DsLFUOSf+jTZ+gelnN5xkFI6vND4803Ki1admqz
vETgfDYid8hz1Qi44QHDB/z8374+VABmQqWvamd5dj0fmAcKgsnUErcL4SuZ
4dusac+q8L/jR235xdDvgTIieKaGjbZHts1T5RS3GS1amruGISU2BMLr8bW9
pioAG+Z0bIbyGifafGHBDyVTm94vKKUCZycSn6h6ypsNXdTEtN6XfOFBZGMW
iIlUr2QNkc5+DkgU7jzVhzRVFGRQv6CHsn9G4/P/ElKj840Gx1HeSwZ/ROP+
IQW2Dmi6iIyogy2W1/HjqOLX5SiT7P+HJwngkBTD8UKul9ppcN0rTNyfpbMe
aVZULGhDydYRHOcQuVurK/eSFHeDGIR/aBa//2L1vwoavw9h11H5csDzGUR5
wOFMZyAYl77Sy+eYIrUvZw9xFs4P0nUXgJluxZT8/C6Yuzjuwv/AnZsW1c5H
bN+qSeFlc7M3Fj8RweJFe5tx2jM6SSs2zqRrHjbSZtoK2SHrZf52CbP1Gxuc
w38ftlc8X5ZDFbzvgBNWC9gpjWEn+IBWe7znwmKuQ0Od+ZVEifQYKAdouJKB
7bdyWEom7TiuG+Jq1L6xdvg//6p31PAZBLlvsenNk1B9Ouw88o9sqD0EhP5X
R62iUmCn2tcj4IQ0FW0SX154i52ta4L/3dtTS07RXZwCpa7UkMAhUg7U2mfZ
0ErjMyZ4iqwWThfRWfuZagok9zO2uVR3olfyiBVwRD/V4hwmjSBGC8sx6ubq
gB4jiAi4Zg1fyW3iwumFjkiGLhNiMbjeKRV6R9LKtP6WUVOaljQMhQmAYviJ
h8nj9ZTq3SwpM25P7IVXUcJOIDdeGiNCa9buiosdolYFQN0GSlRFxjoN/UC8
pw3ZvaQVMpPyNc9ZUUkzfVEeyr2nKkvvBkkSIVIqChR10MDhyqbP2VQQKSEF
m/t+a0Ny1bO9Z2fv43dUkKRBw2BmzWS195swNhmjedWvziW8unZKEicxXkfq
CaGRLy5W7XRcGf9SXRmCDKTkNHjem1HFS9aGHX5lSwL4JQPYbOQ+eccEf935
s0CH8B2iHNdn6yH7r5LCfRKzVI5VaRjAlUZhWu0mZ+DxuVYeiD3gfnSFzRQx
wvY5//ebteXVPqVLg+iQYmNwaQMJTDcTq7FedI2dgDb6/Fwype/DE2VOGBL7
hF9uCxLhXgMUlCRm11g7Dm/RGwK28tktgawYoDFUa9/+WUUA8nzpJh+iSuos
ejBpV+YdzBI/xoYoznhcO6WaImyiCvQGx+F50ZiRq+sxarl1rTKtiN2EQu/k
Q8d3uJ1vK2TEufu8GGLGLBDf+YeFkAt1shSDZdi5gdFCSQGUiOYyIe3nTFyi
X9aeaJrDTr0Z7riWkCHnuYos5sJFqv+Tw20lUYQTpaPt+y1I30CyOyaN5SVT
7g5iJmTbyLVc4COROOhgmboGbtZ4Ne53wMIrmG3Esgqb/aXZlcoiBPfYpnx0
evYGQIfWuNWz3gIxc2PzlovNYvB36j3DNEoX+ZXip422v/YNLYobXDwadCMg
LNJECC3zLR1G049a63Fbbr8+zXHUGVzkJdXnFhdT3VfNtccoCnH5563dZ8Gw
jLw9qww5QtOLEP4CDN1Q7cEozybKHh69BEqiA2ck2x9PP/OUmmbFZ2vjwPLk
QqdbQMCcwu8GPWme1VbC5beBFrvWP/7qVl04q8Jw/Jv7qLRAsMsyHbAdHPym
X8N5oCzkAivQdzSg2cA3eTgMaX0CTPXQmdMDVuYc+djx/etjGzr5DErz

`pragma protect end_protected
