// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
HlNh7NoJwTI/f1UJ9wJIeJdqvlNpGbC1ecYdshW09XXnIzBz0W9LOb/+IdW7W34l
ZAbGOHCowCtAFPwzO7y2Ko5tVHirUasjy6ZuKKSSEWm8QoAgWe2roAdot+Xz+vCk
GS0KTjPXc2yJ3M/02QTOP/IxKq7A/WTS+OvX5re3EMpEtptfk61ceg==
//pragma protect end_key_block
//pragma protect digest_block
v/yauMnHnvsw+XczmNoK4AgYraA=
//pragma protect end_digest_block
//pragma protect data_block
cjgQHSxYdRoHWUBqV8W5CdHhnIagmZ1e/AGs0V6zFVYYAKIFvCmiIbNw+8HYW4J6
XsLPZ1dT9gj+HTwRJljMa3lWvWC7ckAWCCPWXOoDzw1CoLBz5qcvBQC/jfnm8JIG
tGHWJLKckkRd0O2jSm/nP0fRGEGN/sZVcrOoZ42vWoleWrVIL4iMo5F59dlLxKnS
4ysUannSl8sFuFE/OUWSfXB7NjzLPrYq7u30kl9wD8SLj1KAtWYL8Gn2jVaMxhm0
z/hTkbnA/kbv0gV5L+/RsL6FqHL8Rjv/LPqwlgXPfSFjpaLu8QRibQodK4IB+ktr
pvOflTwEgn/2cPj09IJajczuyxaZRQrVH53sZBFnh8S3pAnpkGjAaMrGd80HJBEo
a0R+ERztGW6BJdRhkfJW52qwuyh8Vgo9hlWu4/Sgj/n/j95uelCAeDpsaiQWJe9X
s9PBwGn/4LaLiX6m2Axgpc+wyDJDXgtXGYTaEYKPOA/31DNb1nwEIrexGtfTdE8W
+vNFiTNT4raDvUPFvD12+IHQUgv1GEOvoWUDYaHSRHNXd1HBefFkCymrmBjlHZPg
jqYlbe2RUM7iE90f9L+ZWrKJljeqidQiZ0UtCzy5m+k/DrhLwbmtMui4qUmJgOrw
cqluTA+5d6DKb/o+TQMHPhc1bzdfowQItgtZ0m9u8oWDLs6vTzR4RL8s29spuNNG
mqtYVW0kk9GvlTX6CqL0w0JROHe7b8VyShHDK563tpVzyrbedg0Sm2xSxQuC4VpD
B2VBuNoD094SAzgU6iMV4ZUlkW2qy44fspCQPdsX92wFs1KgGEIEpaAIOCdvRLLq
EWdlDCU/EhinUxkKkmjiOdYNRdg7ZmSvZVbP/iJrjBj8dgTkaQ8jiGTXWAGcWRNr
qAdGJdZ0O1vjVuuGwtYLbt/8T4YB7sAdSD69dVHCiGKAKsIjkAPAtbSzMUqYwsUM
eAaJVm3GcpqALh37qqCtjDNbikuqjW9D5id2j5O9nqsTmuwiD3skHW7g50OhqBe/
O6hF+4n6aA3RmJGC8GZiNbIZyb4xELwkCi95kdtaPdWuFtDi6wba6ZK6nWYzP9tm
q4jK42rnkTZ98pr+qmi3CMK789Ekahe3uqwStBQn2DVb//d6O5O0CuT8m8RrMGsM
ZvF241LoezFStIL+BNS7eybY/ktCVGqKq5tyPgrR9AWqBQzRX5BN+Y/fL6kVwO9Q
rnLwhpklMVOX8gUMsVJ8APIoH8ms88p4vdkvv2VIwmF7KGmY99Ux2/L0IIX5VWIP
UuXcDwPwp2aru7s+vNP/mkQe7od8howDwgUc2/aIIit/z6Rpdzezt4u7yYQckley
Haxph7AVTAH/K5XG4OogkDNB6sgaH7wWAAMyZDJze1qAcu5J+KTQoGIZm7jRQKBk
nDNK9nf5gVWyHC23jwhaZkar5uRwYtC8mwbiSWQpM4w++q3rZ9a3QsmBz5E7ZC/V
J8eiat5FuEN5ajKbr7g/VExX0a3p2ADZJ6ZoFcjMrfnhqghTKO06H/n3pby8SRVY
UdFbKoPdrnXCCJHAEyBN/AquCaXG5M9DseVtoPePZi3eS0YIuhWr9kAmXIqK5GJG
OqQyKao9YVUut6E7I1yrJToRvfC+mwM1Oz/8tRpjsopoKjbEGq9G8bmPeS7Su2ij
xbxmlxJwM1vO26CGkeNtXo1UIH2txqgedNEVK5GbEORXPyhdXJZgy0u6nKRYtP6/
w3ECZLevKUnMaRRS6sTnqphxLkpAGxDfy+gNthvx/McbER92hR99apCEpcQaMgr/
uC/PNkC+kGSgo5zdTl1Hcudh5RZIbsYURMbtI+ztl/Nr4EXJuh+ZkBpn0cW2vZfZ
FYecs5qEis/dF86+4rwjFGhFaSA0g0aTiet72fQSUo0GxiRe3xQstGGFMxCqqs3R
LB3Se1JFw05gqNXUNlqPIoX8f1K4mrIifk08gsrW1hsXyGqdNkMjjxf1LhiB+lQ3
VrK+VRoAIhx48fkPYO8cLWKAXVzB6/QuSc/DfC5ggtv5sDaaZIa5d3PB7ACK3wgN
cahKTfJJcx3Oo5Du7OkWsLpMOVkXzE0eRZGXl56O2hJArcFp29DkDEbxJaHS4SPj
tLukqtkQuNWOqMJ7q9TxmPACGQLWsbEzJIgTXEsoE4aYeeCRlaCLZDgJofHsWgFw
YeAPSOizAGLSmDE4oBV1wrhPW7MtPUeuSOqHIYm7PIinbhL9mQu0qKI63AnEyy83
pv5+44ksBFSqYTXNsXAM6TBTmhRALbWv9GFHBD13BCvYzPUH6l/0NRbRnQOLIpc3
2+wj3FAc+V7RhtONB/o2W49XvEMY5jkS1ZDdjcUpjy3h8hhk00kLq8FxaQlVS0mK
nbukkP7igu7If3T3RrBfdZALHsYM83cXjx9tjqEknNuafGolehz0igV3UWCf7NP/
HqNVcncbuVepVyjKomBUMBLYTHQ/Ipr2CDG+x5mMptfmy4aCsii8H8c1tH4ClRuY
41C/NUdAdDDEz0c5BHoVg2QfbtwqeAzmuCZSUcDXO+JBU27kfzfuxzCWqfH7b9G8
q7/XZAXqDH/NBzgHLGTE5E9po1/qTGezjaDiEOCs5SXJ3QVtk7RMemmJfKUHiFQW
erWnEnnJByv1Qr60XuxvtCFN81yzeK/iwqsxKfZlFF6dNknrqyYLMDpf07I5m1rE
80aCom9exy5pEMz5aFBIlCachmqO8eOe6UyGATuxsrg2N8K20VpOgRWN8atMZMrU
E/tF8EBCeY8CPrfURfDwGV1+mtHuKLkhkL6wMdE5io7ff0u5Hs8WaaZPkJDBYZUW
l6V8lnR9+CH3LsJMjeC+4ycGrLa1529urscKsKl0O/BlYHv8oOtQdJur9qktrDFW
SwgiRI5QsQmfeAfjgKGRQTSSx2L1DDau+nziANE2zJJ5weM4bIj6Thi/tj19zFPv
hHqx0jcwudvE0HCBvgE6n594k1cHqyCaWawd+FkjNxJkaMMshDvfFuJUOPmDwAAI
hQApMCBDbIUvxyOiR5l3BHCyyHiidKZcC38STa9h1DZsFXzfkNC220xPWFNyYZ3K
tdEtoHmM2LZNobaoIBYQ/fY+6/owPhBbZewlWwY9nKIDRpIcerBAVJ4DG7kCu1A+
NerPRFB9ZbH6/ChrLb1Bgyg4LefoOGrPprZa0v7W/gz9wbFjsmlGvi2R60unjleH
JnoIHts3ZTGvoD3aJXPWbFDRTq9FNaL3/le59t45nPWh0Be6sH6z2vJGfhiwnMSn
JJSruATZ4RzSS5OtDoaZW9I348/eQsXlkV3Bx5WCcomLBFNsKc683f0mkFv6/7du
XWH6vXq+IEQ77Hm5OcgYsj94bMPVs/L8jhl/9SNaViy6dNQZy37by1aH+fkoqEw2
KFqgRXzPaF8EnjqMBlFIApCYRIX+Z8ljmtXIx/jvKYabXsQbQpLVHGWJgZA3hKzH
suU+GQH/ynm4z/YgUpXSN8FA1ipoavF4Ua/rkDCbKOwaWEsyW9nFkyiomlaUz+ex
LVy8RQS/spuquVuSjGlW/fdheGNlUWz/mjaZ7F6NdvdeQw6i4lcy15m+Rt028cC1
bcQHLOvFvufQZym/PjcIRR3YqCO5WiuZZEA4u9Zn9FbcHWWRcMl7Yo3zrHz8NR4e
oXiAYSuTSYHxS3C6jH4/bhqArY0Co0fBNMAaQKTz4D2ahmNX1HjmdUY8eTBbVfIO
8/LSo4PVmGdlb/4oU+aWTr70a4N+F7Mlp00yrNQkL15gziSvom6ypf9lSvmfduM+
fg/iZOFd5acLLbMlirnyVMY8BIj8D7O70JDo3PgVssIe2Iubk4yrTROQvLbL2XQH
UR/NrfAdtp9XdhpwJMNsGYc10M/6DtmLTUCqGOCzRVCOAll/4us48Jk4ncfIQLVA
D9kA1FIGddQH+MyAm5IYoEhKyXyAfmQExsviiCKIo9Kca1LtZTTylltM2agmZrRO
9uIy+zCn9BXatnv/yEJPWOqplROVl2lu6Lba5kqWBijIu5j7Ln6ELXbQhmuhYCJH
+M+JhgoE4iTdRbbFHl3EUwBEMQBjBm2kpSlaKmee/HWgsFkmAVGmMnBZ+XT1HFl2
OG+xqzw0uWykui/dBmaM8mnM5an5Kg6Kfb+c1zlCQffrExSb9Inz1NELGDBq2FV6
p65tGciqzLjbLcI/mCmbIi6KlBTOnj+vewVVEsm2cNGKW6+NCsYSiBlUlXSyO5lp
me7CbWaJXlCndpEevE3k6VVj0Q3igHVocQ+XJrgplIBOSToXOhg5QxhNh5iDuUHh
lJvMr/fdJ70PIoWeK5YpUNgjt3+7ZynCGnNdbNFPMiMGQRYErhdP8M2nhHwII+PK
nTMspn+ev6TNibNX3Qobxt5vFs4Uc/6I/qqAWnkx05FALWthBKt7oM9qKox9h1A6
m1gEn/OprrG3ifvSA9Yt7Nv5rc2XPIxjVs3EHq2d4W427bsf5i3i9RlqO70gViPf
LMcH/x14WhWV0jAAZ0jWnplQ5lzQ2japAYTaTAdo4sfeDVqb/iJA5iqotY7Pg6Qm
7AZ/2k23RDjSRDx4anADdgvp2/aTdqDI9aT5jI1DiimR8tkxX1RSS9clHwokDE8f
mTFoKVRWjmWkPqV1uhN2r2S2DPU3w69tVQedXNvcwFCRNMLBsfnXVz0T+nTpP22v
mxFRohjDpUvuEKWSs93Bm5x76IZpY6tBWiIU607UG73OoOItQs47kPk+4GXtA1Pz
Nv5ZLK2cDkFeBgrj2Uhc8NM6L/MDpLovM6mTek6Xr6HMIuPOGWYErdfgafgCIf1F
rCGVUXurv3BcHO3q08Yj8l2S4dJuc++AUwPdR2tLMCVCAauiGAk5IaEtDdAqSSfI
QcDX6m6KJWoom4pqtJydD23bmu2EvGyee4+8c4gHMv3mcUY0V3UWhQakKyGY4T4w
FHbMXn4pa93Yc3Xzdvv5f9g498TBFw4S2gbZZwSWuNrvWUJYPxz7j9/P5QP04AYG
DkwIvq5tul/6py76EhN3EL4TXmyy8yuk4SiNB4SFRk9bEHxbYrw/c95Wh8hv/uaE
cVrhyhXvLS4Y7vXt6fSgVdZ6BXvAp06tC+iF/suElMDudypHcjybKOrUJQXbKa+w
zSmTI+Xp5nMKKrl8yrqNw4ZQIul05BzsJktsp7nS6a9iZQlBydwFAQDiej90wZ6n
hPiOEmLkftkZDcAYBGjkknJCUyWvmxrkEleXvjqFrBYZ83wWcdj+hmtbMLp/H7BN
w+dhIl/w1D50jW5gmmz7OuY5ylVpQe8yvKpoMFZY4FKGJsgmi7KGVgMAS0hXm79F
29u1Jig/d/inBA7OXUjIF0H8eK9ZSDFHOwIgHk+w/wuBQ/ZOcdgxWuC4Y0YcbYvN
+VHg08fS+FWOZD+AsdN2/JU6TCqjRSvULCfKRp4ymmPBCymBTjNoAtKNubuLolo2
T/d1r/TjZk73nV4SduhpDxaEq3C1LxGQF7EDR2SRaWU7arOUCCP1LJ1TZQFbQyky
KU/hCqbsYj4Ki5zIKoj271YaUfl8mdiY7ynmwPObs5POrcex3xzaivPWQA3AzX3g
5mTS0UxvklN+9glugkoEsigf+YFuf1COIH1hRKWri6dyKZIDl1BDMMVYPONCwRRF
JQzo/7JH44CezpnjxpuyN//lPzGXA90b8/QB10LZ3Bd0ESKhIYjBgrNqDf8nFVwz
e7Uhs0VKrg7fZwnra3YKAkPfVqZ5XrsItLbL/smSy10aqamYGLJzly9mj2bJtUhl
36EAYNX37YYuzPi4KoT8d9QFbb+A4dp0Ia97YIQNMaVzbebAxZBCfRauU/Yu2DR8
UGucrfErtsXB3XJjtWgga1r8eg6ftx+gRl55OehXGPtLs1Vf4XnL6S3c04nygfVA
62ZB87tRLCzXu0pKMTOFJRF1RfhvB/xihySzJB3IU08zHJlry7dqspKn+zjoTNyl
fRG+KFPSgk0/VkTn0oR14DHCawYZV5o2JG6OD5cxjGf0sghCuobV8Shikw0WDIYU
aspSCoA/rqCg+eItPc/IjJNICzbws6PQUuWBHI8ezEnAbglip5bu3O5PrdjZEOGw
86nVXfso4KH9Dw6/f4QLDqhWsdY72uwRGddJ0TuxHXUN0vsDw8aWfHNhmAPNve0j
SJtQKmjwMDOvVit7xxtT68T7YNbVQqMFqlxiLJkkpRBLsnG1r2uUrY8isuuj2cbz
QaNGLY7Gy0vOtREjxY8bR82qhCSD6AbEQk+WogHsJEUc/yntY7RV3b91KLiSIkLR
VmCCMVwo7nlc05y5+CDYbtL/GKzcDPu7jl2TXGT4Qtsi2xycy9ZzjajpomeuXVW0
NRLtdm2yJ97LBq+IKcQt9sLEbJN4+G4R48F8bdtC2nmR/aFaDsfSDsVlAe07EmQL
Og7ld/GAx2N+WQLXuL1OSI27/NuDkuCtg1Lhawa0KnYYDWqo9gh9ktcOfyEFbUgO
0VlpQ5IEBJcLFQncrWBILmTQ5PVcq2g1IOHD5MNOB2SWVXcW+ghN0G1ujIlQA8C2
6gqKzkfQBt/vCOQTewiMynubDwSldbmb+gBodejQerexHVhNv4HuvdmQjgtunfkD
tg3kFLbWOtLcv5HWtgFntZfMmAPdKG90abBuDvqlDDlOS/weisK4en0HeXkX5/If
AVqJyxInWbxmdqd8e/LP1Avqc/G14WraxetGHEIAeB96nm4GSlEynFpf7AKsfump
DcfU76Xm4f2UmUk/q+3kx7hENLKJa86vgpLHPLHTYftRe+E4eoya6vFfuOBYuQer
MH9wEHhYniQ4WsoRm9XUZH0GgEpgZz2+2Um37apc6839PeBsJyN0cFPCm1g21Nrc
ZOpFcg+6J4YR/+R9rD6ekFIN83MCC5TXU18IX3fmhKLgE4WBo1VbMd2bz1kAKLEv
/s1SARpSXtNVpgNBXDcA8ede+0zAcjFOvULiQITnyWcQZRd/AgYN/jka64ffxW9C
lI5GLE+Gft3rMN9pPctn2A7AnzL+nyYfYTTYP/L9lFeELaANwmI8tcsnGGbOHsA2
EfETI7sU9lWyLIqQDRJa5vFIotcjeMvzjmeHuVZV06lwt5zu7RMT6jUZ82WL7kaC
evvqi1eanNbstu8SOnQInVQXKNoyONZN8xC2ErW33LAfq77nr6jMSsuj5b8ySFWW
O30uxEPiCgYAHxyMaaW8rL/CQBeBU00o/SOGM9MUxABCsE2sH8fL6sNDeBA08LRi
LRl9f30Djvsp2bUDyXk4adWIjVPmHFKIMLWwBV85PePBarXeWvD7eVefiWbfE64E
iNw67tV1rhDFgtmQSnhu3A3fSi9IDXZ5eDVhqRDAKGq/hqQO70zHJHmCm7T/WQt8
mA/LyPBd88hnebnRE8gpsAntmHa8AzyHpdmiVd7FvCOFX2Pur8uiNuFvlptiltVB
OWB4xDmyl4JegiElS/YH01YkVxDym6wt7dMLfiF9DKMHGl6pOhRg/7Zd9RYPl+aX
7g6W1pRdP1hG/te11kq8xH5sJIgwoSEwSLTv9Reys31697L2rdncWAHs6ojVony5
/Lxi+TTZjNJ0UpzzVzwb2c534zJKxRRGFcVwKWkRgVfKvFv+8gBfdFn9t4r4ShQa
uvBMl3X97P1spowuTrNtiCWzYhIhcMZfWriYb3x44T5HWgvm1pDg4I2yfmb1xy1A
oQHfZwTE8xdtC0NTWeDWSKpIVJtB7A56GGeK95ItORVE15n3pE8dqVGGW9wfPmIh
FEIhQB5bs9qwy5a+/3n49wJ8y/nOynNXK8/Oc9apMAgiAQS57Cm+50mniL+fWTpy
EcVKSnOszKSMUKmUlanmHIz8yI/njMvclzDbzvoKsAVLQbcUTux9T5jiy+F21mya
BcUaL3gImGHOLi8zWB/bLfpqC+HDpQvrusZta0+le831b3Pgi3eKYrf5EJQPmObW
HLjS7ZB4R/jrCmE/2DsL9Icpdf50ZyFdOBSVlKlkYwSYjCDt3NXdfOLlfALbDSmB
YN91DSWRqiDRA4qKo4axqBxyWaSUGEyBkZmeD0x+R1RZG4c6yHVkXkaEc+ns4Uv5
xrgWO1VYDuDI5bXa4nN7OzvQDokUWquFOi2OEOjNSuMp8gvngC7y092czikAMEzm
1eS7y8ua+Dd/MKNehAxdpAC9uW76DvT/DuSMgld4v1P80G+ILAc3P90m/oPgZdeD
0GEY9oEylTkDm/+JjeWAqHCZIgO0/7StP/FUsqlyhB2+mwzsgg9ImZ5TV4RVc7s/
Dxlv+X/kQJIHfn0w05GCKOBl19vfvdPvTPfcSFFOLx4heV9rhLgg4HSkVnuh8Gcr
xwi5UfoecY3vegQOcmImdaR+/HOtKBPh68Wjpx2OIyrHLbqqjxjy5m70zWP4W384
TEOOvB68zrt0wjSXRMSXTRby5MlSwBWbdxaYNRf/XJ1kh9mJD6ScQG9Te2K+5kWs
LLAFS/tKMBz/PWygVgv0y9psQFOnXw1M54CYvqw8DuoBP3ejPnPc7acRT57CwLgX
GmNqNDNCANaFkwl1HUoEiyPm6Li37+co6nADY8BSsi7BMgUs9kVe1iOMVX8RE44Y
o7tOY18HmIjuzFdjTq6hTtqP/7WPa0y+yEmN56dzyG5W1H+A8w51NoCPwBeh8aZ3
qps7mO4g4erOXxbn7v0QGtvnKTNLzVasp5RA+VC7Ejw16T+47TDZLhlHo1ev7fPc
zQ+3z/BIXg4AGYO/kqyJCjQt71TSycOL6j+Su8uf/P/0G1jaAwWsSXtP9DLwk/4u
M+QLdxlv67Ams8M/A6dPCiBj0nY2v9XXRscFz9cjYyvZCj4DSzNMzG9unkgiMUJd
MQWYADckQsmzSmjfJMFNk1bB5x0bmTVAvPJoThBiHXw5WcBiLjP79cOF+6wfxlMQ
X5CmQBpW3I+34BA4d2MV1yLFSRXTuw7yJuvCef0QN69za1i0mW6TcWX2tMhnyDoa
t4UNlulLcm5uQ8Z5BQuQA6Ouf33ylwhoEvjzs+8FZB9N22NqGkwCZh8dz1IfBh13
nEJStaUoT5hE8SbYnMKZgVZNJlSgpAoCPzZueTwv7s5x99PuVcfFBsttqQm6ifKt
lK44iyBI4miS5XFtUYFB6ZggxCzp/mlugwYPNLni/YfU80NAzXkk6uSf+jraHFa8
zToN06kaMbSWOQvoqmaVGkGgFBlbjtllEIB4ch0mtGHvKVi7D0druGf9gdMszu+V
l8nPnUcw5FZlMPpoBSKiO0P2pXVLfk3SSxIK5mFBt0fwe8Yyr7+FrLL6sQDoyElw
pog3ko0auSGv1zLyyb95DNvqWLtNLgvpbvybVnuDbKfXctDoP7sBb5i2owt7EPAe
4EF3aCNsZZHicOQM53p5cff2sGexfyG7jI1omf+pgMScKYJkVE6yAsJ66R7bOboN
7uMqChI3rgeTh5Egbw4Tm5Q7AlhWVEM68TypHQZmMol1+JN4g5EgvwTPpK/QAba0
PlhGow+CAxykKLUZdxpQ43rafjm6pm8TrNQ4xDrf7eevyvgexZdcEimarCJDhjln
5zg5EQnOGk67CmuWf4ILHQHdlhWZmrrCcgHZ5V+IRhjyhIwBHfX5jkBlNSKVioWW
KBPJsNMiJkMw87ZruWPqiA6qp7pvrvY4T2HkqT/rVWi5x9SgQE6sJ1ZZ72yUFKDK
L7OTmvw2HZK7an+Dczy6PCTCn1Rqnu7AxMpU6dZuAAdWbRBAmh2zK11umC8nXuL/
ES16DNChF5pjxboygH1JY7Sti/SePsZztxpCp5Fy1o3f0OlhcaXpfvbMLK2F/qSv
ycv1zbiOZ39W3qG3sVKiJKLitjYwdaGcG9Besx6bJg88QbMHeTi/clOtiCf6nh3W
E50IFu187tpT5PZmbQULPgxrRC6i7YTvSc0nHFyIfzzzpFTpKbjWHMd/9fcNHa3w
DGsBemrHvqecqyGxF8Bo/HLZNL/4haCLqrQjxjn9emnPMVd0c+dmNU6TqWAn8np1
/+XldmCPeiyHBeUuqG6XLXtTAzylyuddurEN6pEIXD/8JC6BXc/EXlpXdhwnau/d
9luxKDJIau6uhrx/IJCUGxSPsCIKTzaafPhLnI6wKnN1hY/+kCtcqglAC9lNQQBj
2g8/16ngRcrrxh/5WQtoe4dsda9L6hV5lDvg6sPZq9YvnCoxHQwSY5MbEl5+ij/z
tkvEwFAb5dmvRpW6fHJ/NvQNZhTtSzcpP8lW5HPshamZrhIShXR+Wda5wnHT9/Nx
haLWIsll2IR9XkZavyn6XfI59vXqdhzKkD8A8l2CJu2Cogcw1fn/YDbILOPbiFyV
uWLQdq6mmTh+Vpn+w/Vd3JbIbCBDOiv4ls5vDIbaJdl4aoaPtugEViTe6JwV8TcU
Hpbo5/Sf7NasMENHMgFsPeCVerI4cS5SCb0FFlsiCAPqScQMioSi/HIg2hWxKaPx
JbgxWgqqLZ0/s4jskAoRmMffoT2ITEb7/M/ttd43dRE3gbR4fSXfjew0AgBcrd4C
Ptk7ZakaxwW8SjjCYeG/4fkSaCeM4+v/Kjp7rkJfm7HDvmIyGfxl/CS0YACFPbMq
gELPuLRKYuBmXHK81ZuFoabJLFmhM7xTIkNlR4fsBsam7jCQ52gG1Rl+p6IQqb19
jGUtbwWdsljY7yJbJkujTUt+PXvCuzK81Ad2DCNha6Cu6odqMf6dY9capsoTkBCj
wVCRZU5AvA6hULhhhqs5cYNA3L4R1Opv9Si5BD3d07MW7ufIf3RbzlYXWEf7lXWL
eNq9r/Edzgcppt2odFQRNTRDM/8IzqhxdlzWPwK3L4ipCom3hRUlLe8TsCLiPMIQ
IUmLuX0dj5EMckkrD1FZC2It5Dd1pAvL+8XmahA3VSzk6p0PrAqaBrixnyM/mP17
e9dzWhLeg0QM7vurcNU1W0Y61LRWPexDdvOLUp+wnZu04xcMt35+mpq7ZMDvwBgJ
RVHwVwQUhwf8GK9yU7KwIvupH3QU4vicScXEIfFiVLp8I81kNAqJ+i38msxuJFYQ
ESHsfAayr+FqxpkXCWuq/CKQtCvsp49GIalw5WTsaj2l7RZf/wuy2MVV/2P2soI6
Mql34DA/oInbEImfMwdNYVEmnsw3qtvXJRI12nD2aw/78c0pcgRQVff1GlV4jPaN
PR5n3tZYMNy/QogO+haTZFlKGxWkfauOHiwZqBjG4pt4dZeaEZ+TX1LyAeM2cLA3
ZzEJ5Xwnc2xyEkNDl5rmMx8muTy/IA6zrgTda+snlkH8DiUEY/IK7384gCU5we1q
sKxnmVSP1jFZsUT9/SlraBHJCvFiJU/8UCDtfcpZyeFsb8uo5hBD8+fKmqTC9AW3
/NQiw37TSfiMHVqfAnreqZbnsUVHfyXXIMuLTjBhPtdC7iohUMorG9oCqTitaZF9
Dy52X8EROMvA7/EHA2MtTZa2W13q0lKQUq3FrWgeTJ+GXuzUvjh3VXjSZfSfAzHY
bh4DyYq+bjCRCRKaY/YhT2pq7l1USv4HIbarPYlVp3aPELje4xqGOl5WM/rx3p6l
eIr6n6M5v02ZiTMIGrnOEjmmn8+I5Dowb7ctm+8odEEG218l1+1UvayCDj3lVZDD
sNvq+SNTtiWwGo0UiwrO+KgkKBiiD+Uv0Vt3Gi9GhKGpM18TvQzCkGK30PYojP/3

//pragma protect end_data_block
//pragma protect digest_block
vF5AmcypASaJB/4tshn+HmHJpb0=
//pragma protect end_digest_block
//pragma protect end_protected
