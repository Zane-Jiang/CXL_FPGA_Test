// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Oy0JV/UNY35GsuwqzH0E51dzqxHVzT0i/FAdgtFPVp42Vs4+2vGXzVSGLB7SeXCx6Q+mhAJUURMT
1WlFi/XWZ+aY6RVtU+h8Vglmd/CpRoVuQOrWrd/6LbBB2WF8X6kRnj0nfgydtmbTG5rYx5CLmdF7
LgwfWw64YFdoXHIFMHyHb4HfQa/PO9Il7Mu3131T++q4uWRxs0wKKUHmWue0+KNt5/vGgJqg0TSN
9MEWjb2bVqF8tseMfyF765Zl9OR6CA1q2cNCjs5Gd13joK7Oe6lhfSFtSzCxJifFbF4t6YoWz86X
hYeGUteHZN83b6ArAXFtX30K+9kmla1jyJjqRw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
c3uP0U6Vt81NSfsQP2zsnYNVsJv+mjFmcS0Zk5YSki2/2AcoX20n2L7urlcpNER1l7G0bTQyhpAe
GEtQVgdFg7ijmNr+s327gCaXsj0loKCb0uFr6J2s29EJRBVXrmBILongHsHF9nYU74/Xi0ATEeZ5
WYyx8fPq29OP3K0gkdkopJPC3mqPq223ir7+jtTD5R6eealvIDGV1gmCDlrSDG446a0rLInOyw1l
FNM8Yvgv79LXP0bLCHaL2jnrjQQEJzsHESIH6z756HY1TeFkEXlvWu10MOneRbsWVEkq5ud1siEt
vhoZEYhRosziBwkICbmNnShCoBosA8IwVrWvv+7m5iLq7AvcCQJE+CjIx2INPcb7bGiATyEx+1Qm
FrZ1z5pOPUoI4iGKqNY3GQEx1POirv1FDjy0bgJEHROE5Rbfi2b5VqG/QvS5e4ZcruyCQbVj3Zo9
jw4yK9CpUO477fCROgU0xQ/UmYpiXYDG2JlJb0/iTIXe0lxWNoq8sv5QBsHrel7HBytO4zCWjoUn
qBqcnVNUPop8+Y5E6IJz3tm9RIIM1hvkrzuSqYAucvat06l/wiPN/dMk4tFBIBoiCACqb12n9bou
fVLLDCpLF8idjDcxNXcSwX3O/DWTeYm9SNFpdHHM0Gg02b36b/Js2f/iuXsVwrymbdEUgL/zj4DH
1SHsBywcg+hlg0GpqrO5OZ2e+1TxT7spYT70qg/0X51z8citDBbeQ6MREri8YdxMKctV+s1e3F2C
LfSu+ueCARQVB3q5E6pRdD2jHMhRdVW7KlhNKvIKRnHllmESTeJXgc2eG8WsG60mlMT4jaJ+kvXm
y7LHG/YNa+B7MEi+34/i5rzSTFlru2ModORoqOu0c2Xl0KJedPVTzOIOdjaJVndHEsgENTpWN8IU
dhpgd7K3fa1dCps4uVe28vLChPt4BUqTjWkbBrwWdACbvaavKHX8nHMxJrgk19Jdu740Hf78uQD+
4cfpFMpMAyKCs3FY9GxHacgOsOSSW5GLUbC/nrV1C8ay1s9nXAn5Z/gj/F/hTs1Hs1W0okOaAo4D
nR8TYKNWCom0WIZ98QaOrsueCIwcX6lqKwzsMktwNh43u/ODcfK6NjMe5fSusSdTD2J35pYRmhe8
2bd5a4W199STY2bqUud1AITBWT8j8yrXiCC98fe7D0UehyegEqsEo2fgQ0rkvC0amEWhxlPSBhRy
zjz6t2k2PMH+DYjvySMnvlzqQN2gsl7RET9GFhPA7zD3djP98jipCaADuljAOX3pgry++R4fgBMc
bTQOhJXJ6oa8oMatxK7I8iViPJDCrZcXB9Q1J+vCynwHY+Hs0481KAWl0znFMYvO461q8JVENUQ9
aKGIhrdZK1FhXcN0sQchQzkIuzO+f03JB8u7aFRLAtqprXzEaNrhPx6wUv3ckvr0XSHa0oTkfzP3
+bF/CX12g7iYwMpieI851yRTCaV9ml2g6D7qnSnOUoBwdolTcjVZ57s5Qdf/uLoWeM8JVy4jxFet
Wnnh7n5g1V9qk3CfoHp1d+YelrYfsSy67pyVbYWTbyZwdWfEh1witAmPvovGZbjIHwCB/9mknUEz
5l30Ed5mvLYT8YDsv890SNGELxRyBnjDjqamdi1cfZyqXTyZrIM/3NnA1h7jeDsZaCyzK7QDm1oR
7quEnYGlr5JuNOVboPGqFATlzD1QtPGZsbpBVFdCWZ2VzGCnbZBMMMfTRloj6bikZ6QkR54CGqko
9j9yEoVYaix4UebBRRLiPLWSBdBsN7mUz1Glf6c/d07tTeg79Tn5bl7EpkruY1KNRbVhS3xfYHEo
Mm5IwbAe5+lo3MdreIsQ0S/no0tX5WiQxwk1Pf0sTuzrAX61gnDZaQwV9XCgVJIrRAQmU+F7nLqa
edvS8FnC71PpIKwdngkIelxCuE1A+iLIhDOCAIsXV91Eh9Ksb7tYMgXBQJNZd3lRmlXWCC90XSfR
guQYope/M2iArjJqg44qPoiTTFx3jO8LsRTgECTMQ6xieRdlJGmxhnr74XyERlCORmgCFni/sZ0v
nkv5NHJ8IJ6D2aKCJNxxe1FWTnhrgS/f8XEccPpccyIV0FnrglGPYfIYwAsdFsXtFGPJebmbAxCR
HjFKiSgLtsoWxivZBq6JVRXBRfHxCFYWTXSMG3BZNCBadF7d1QIFWHK6TWOXbP/d9YcK7ROwwdqx
6EvckeDrCczGaKc/tmkK441O8BHtXxc7c6b8TtmaI0sjF4tnG9BkcUR0mmwP0OX2D9evUxKtNBg8
qWI7m1L5JAWNhLO82HmEL8BR1jK0rSvZFgwOjwQjG/V596MRegnFG1YpYXPPcvMfrPqISmSoFhjq
3Kjckud0SXkya72+C/T02moXJyY/ZmafBKi34FZLN+AFCxnvSUykJyySSU/3zC4IBqMGM7koCU4r
1F2jjs8X5VCR13v1qkLzujrNNswktJDYmL/YB9JaEbaVN5kCTqo9ZCEEopsC9qFoHYX529L8QroD
qCiTHdpXNiwQ65adOaKKEdlqKKnD3RF7evP7WH+f2o/AA5dT1jw+rYCAUk+jPPoFY8wnydeh7Uev
ojTSryJdHxdIpMcobno2D1rpfDMUIiVZWvknaAnLAGOWSwFnvFbmt2yAdPPkdAk5gNKEbVOxrBB1
sQGSPV0J/cWflTvr5mHpJQRly01GPYsIObl8rGeKS17mb4IgLY+wJ1h+5VYNVy38DKD39YKJMlLa
dDvhIRGc4QZnFyO9wHFeCDaeJFg6IgF0fdsdLofgscecQvOSWq6DFLtVAm9Il9uNXagIyTFkeOaq
fAZo+tlqrE35D9JkH4W3nVqaAL6+evxsSHoXk42f1AvUtBoXWIXT4mwBhEC59/WkZzwdxJWQFT7u
H9MVQAKAf5HzbvaBR7WlniP7Nf9xf1GvmhDqskW+T1DiacqbHiGXxbI7ORgsR8h/53O5XyWeCd/w
6JnrEZf/0YKs8swNi74JJ33JjKdWyV+7NhAzDJFlWK+IrT+fXFPYc1BiHIFLAt1cDaBOVPwPiy08
UBgF7e/r17421i3ZH829zm63la1PhV2mXATyyPykCWVjD1TOu4HwXH7ngMuvlFF0X5mYbEPsNM7N
FrjVvF2OT57roQjciN097CIOv0BoenpP5W9xZ0dNzYscrqvRNLcEVfebamDuKkdfZ087omfXoKSJ
KD6wg9QKMeCRVuBteQzhBYioaz1TCk7UpEJNk2h/PKEW6uq/FXmN8c8t7MzixJ/8nzFXvKzQ3nJq
cOjHshoLdwPoYOJF68z3j4cHiFM03B9WBbwcM9alKhC50+oZhX4vsOhmu3CDGRSX6+U0KxKwJDpb
wN2i7n+LHI6gKCB3qURKgSt5FtNiNdFOmBaKBtyd+J08jxKj+fnXtqC+dFyAaXhbw8ZnvBCXTMwg
wKWW+3wRclbBrikIA3oc82wC2PvEW+qbrsyuYx1JpHjc0Uqk1K1D9KpTYfMBb7UH0F5WasaI/QE5
q6VVbvA6kOhq1ixaMLdeF+lLPZ891rWQCSXD7ClvWuudxUaisH4KNOoIs0uObo2SZ8FBStqkIZ8X
DhokJxTXFs4gIuIeM5ui7bIInEUNyAYh55ZCPt+Qwkb2LtJJ7F7ODUdICNdAJSr0h//EKWMkyCBw
6Rf/eX0xlAYlNkIyR9CA97kimw3EsT5zBv1J3HcpRT+9sRzRCxWlr5rDENS7sNbz/nW85Ah/uSwX
xrEFyuTmTGaT7OWTP84ctyzmPZdp5oHptyJKMMe4BlI6SK5QOcusHl029wN6OivcYHREKyalbvxb
pz8iTmW1ZVPXV5m1Vx5apdKH3x+KqWMo5lcBJNahbIEJVBliCydC8M2tUS59rQxZ/X+X83oz7lz+
oz2/8TrpMjzrZNq4kQOFwknhNNVAc9biwgnbD0judgeLYeeHcVGEUtCJSpKa5YQW2dqF0ADcbBr+
Xioy9osRiKI6rMRI/edALRTHwNA3cYw7mGOh58S/0JnbZOqZh+hpkWdZqVl+Tixy8eFhsQw8F2+g
sE/moMI+ZU/E2/UoSf+3BV2zCRL9NrCzLL1vPlVR3jPZUNPb0eVMk0twWVhKWsYn5e3Fr+mHp2PG
Y+OOsuO0gb/C1Jpu2maiNwoAgATTrW2yRYv6fomtd6jDQNOaXFLqjGc95Y6alh7u6j7hHi6nQ6Zt
NlKzp91OGPgAx5J1mugHG7cb0IxH30K/6DHUyIbcLhB21+kGaWgnpp95ACYGON9gnRWO8qx0Zmcv
9FzhrGCdY2I2at21F/0haHIsplDjnvL2642wQf8s9yJ6SDANVr9MyxwNwnRYSdLOP2my/+aG6x9S
PN7d0TjcF6dDuy+/jgPpmzIdAKk1cF2nI6Hi/zLl16HgbWcbyJxA3uySGQUic4dMdCU3dgXM6FGP
JpvEt0VyjwPUBoU5JPY2zx5FB603t98+jgHkTCs1lZSfXmvAQH3EHhtypBeeaLLIcV3BW/rF5tFl
Ecb/uMTWmaFPetoOBEm2zMxu318tdlCOX/EGs+rxbELmhnN/JVhSZmuO5+cGDGIRwsfzfzyJZL+h
DREpFwMY9ST2CJSGIGuwiTL87gT+7GuIf11/Be4xE8dEJ8nJS3jOy+FlaA9AyWLMABXBGe727+zS
s5XKKRnqPg6reX87AF5lR78qEDv5gwLxbty5FBOfVsKICs5D7bbAsIdyXawYqFTccLwzKKi95MCD
7td8YN/tlyf2i/3AiNxTIVDhYNf4og76Sse27pBPN0/M0ohDpVqZhdWw0hOhe+174DmEYpRBr+ji
YtktRRuRFU7Ugkc/KGCH3BPzC6okwbP5ECuFT0MhkFb8d6paFZdElYDEf2EQFh4Z922Eyz5o0vht
47ycBiLf5r15udLKzEg/RffjSU3756mBtdXXpzE6zZxM4+p0VmU8GwDp/tggj0iblVrFxYgBzx54
chR0pZv0dY+nfdewq3kaImUIYVy6z7KWtA85rwc5Ogta3zvEa3f/O/ayv1w/tSOuUku/H5XqRHQq
HsG6aposkVLyToNqtIEsNSMlCYojcmSsqm0bpfECyVeygrOZtsSLP3LlHFKJUOed1sn9kDOyFjst
nHVA2t0TfthBuq+Onmi6gultCbcDoJDFTWM5WsfKpX6C9OgaISwB9VBkHGSpG7izkk8HyxyEfWdr
KdDOU5f0YNocbRxKE+ZyGwN9g7K7x+uThPhZMxjL9dnIg7uy4OPfoOYJY/O2z6Nt2ZZRxuiN5iUa
nmMoBAhmh14iZpi2UxZoCYzDOqw0Njj/cC3LUZi3t28I/DCnwh8NwkAK1F5fi4BESposo1SL3rA4
Cs1DrW+WFo8oUnQW0dqKtFuqDso5vaGheM7VOgfIYgq7BDDljW7f64BEXsFBKdiVq+xo0INY3Ccg
aQea/M/A4Fw6Tnb+Nps2Atc71N67kMVVThj2Rj7SHKAt7Lu3ONGFImPEAP/iGQjjAvFjw4U7iWWr
cwaCVxhamk19WzCNVj7pekb06YPGkggPWx98Xc119bhElEcd0TVwYGBFDnwWCT3xm4a7IfYICN6A
dDXp/HNS9wgf5VP3Ee+DytRs0d52DwBzmaedmQ7YKKEO+bs15LnpJFennzLbt9VnwRKRP332Iw28
R5fSsOW2pSzRVQaIfUQossa8WDdgFC0XWTLegdKbE+/4KmsMtbWHTcmTVElNygOqZj8Zi4aCjSIp
ZvRCnwkVH4zbNIrAgnMksAIxjfOusyeC4jUM1xIP5U2Qv7z1GsF8Uuv89AIuu+ly/XqEJimKIgTZ
MQR67T9y8Q+G0cF+ff0iJSDs/omsEwMpFumaayuw5yR1XH/uOzKvNJohijFXUPXdAmX1XKOkdSnv
/4cecBpMco7kLBhYHTiLE9x2mNlFGwk4AnOjIx6VYpY+r01j/OIePnIH0f6zCJmZbh91QjPOvEe7
aR5A8xl8NAsnKMARfyQ3fdHo/Hi7mOAKxAtsnLiPJbDntvh2+jA3c1eO8B86Hifoe2MAAHpt7fpR
mEc6BkSFIut5hg53EE6gL8997wZHCvYcQLlmzxuHdbW3EuWB8p/VTLanvtNF0VCvc6U+P7JkwjFY
9gRALSlo54DURUEthWzEzNO5vaAldd5ei00eljlr8h4/+5deCKozRb7hKPmocgraO7tid474rFVV
vZ6J7aptoYiidPFF1O0ptsJLxFceaAnVG3kLGxiDliog4D5JaS+9bqfskVSCcTMp0lemLqDM0tYg
ps1eZJXjBdfJnGekm6JPsCdKUEt1Im3xcqrWz9irw02kL1X0H0BI98Sso5satY9DMT3JDluzVFyj
9qM5yqB9kcvHsfSyo9TbQEEGh6hbZFfBYBj5WND0qpQsHr6mhWmfi5hbui6rfJnbjM6dUkOKQvmz
ujHDMb9x/FKTaRIkElNgI95CCYW8guTY3tlh00NU71mbPccwTwDMdr6Vc7EYncFo62G+KI6uxWPC
0WJDRox1e7UvUyrvjpxCwJDEn63dJVivGrxtAnA91vPpi6dzMG2PNgyxPMC611vq+4jxDoBdOXo4
BnxfuZfqcPUW3FnRXIFbTYOvty7Jsy7ssHB15sWuxVf6L9FwnQvHLzJ0WcH9cO1FLxbFhQhBGARD
wzqq4q2Y52NWnh6tDOC5loyYNcJlmQWk9nFCGCMLgStVq6cTxHah0BjVBy0TPwKquy8g3+2Oh3H/
OpTY/+A24tqFGB9u/IV5Zm33QiWl0rfNSsUtCd+SsSJRNOqevU32RQ+HwJ/Z1kYn40etYthW68Fv
fW7OwYZ1Eb5ftXJhRVEqZDoz9i/ZH1soZzAM2kpN9p8FVT+nonwVK5E8jm0IuUQMLpKgbn4CJfln
wqpYVyDZ+qPvY+Xeu3ckKQm4USUPmVtfWu/iOZMccL48mSB+ZWw3JWKe2xFOsl+BuoqHm66R5ggH
TziaGAz4j7keZrFL3Kj08YLIOXIJk10h7L393wng+/4WOnRupKr7pKUUAD3He0IJeAYYsaKvFxw0
Lv4wmVM6zIkLhCMIsWt8RCzQp3bx3oZ47R3KwDJcULV/cBLsgg2BYX9MLx5EPWShGy2O3uQRXy3X
Mlcm7+th9DVw9n0f2OcVuikeOJnyjNvHl/CE3BAqU7cXjdnqROTOkYdgH0WgYRfdUKcKoe3qyoL5
J5vUQUdFHn+CBFDItxadIQHVsX6he/Pl0995E3gqaoVxr/ZkIsHaP0hdTCupOhTdwYPsrfEo8nhJ
t1BNWRIoOmCMbclffXi8BzKsIWVs8FqB5Lq2MiiAtiS/PJgq2nmWzi5ipI9N9VmwpESgMTosf3MD
GEYwqjfPaW014J1OI6cfML+NDlVdOhgloTYu1U/oEn5M+Fl2ux0NTSVbFv0if9CEoYDFKRAFfzzu
iz5IxK544xuPibBbKJPlf1fQdL+cdwRdHE/Sv2u91ZSKiCXhdC3HNsX+9MK6AftGWtOb4KawT+Kf
ViANWeCSevRCk43T2JbMhwPIaVHiOWN+7k50iFVE2QQWTYm2sCXecxDEJKoOB/Uyuy/ogBsbEOlb
o0+Yk2U2wC4AJiHtRg6pN4ydmLA6keQUz2votOGiz1APiDiw0Fk5X9Hb/9PN750zxRuSkJhl+WTf
vWrq63LPVTDWsD6VnUE3cilmVAMTqPc/xjyDobPB8J7hwiJWcN+Ry+B5d9r3A86JtwMEMQzxWCVo
aYlVhcq28WzjLzSK3gz5O+73tplg1GZGcIOSNhuYBVzcO9M+AfVl2toD3aVKshFYnnb63JlRNvkf
BzvclOjkRbbvfztp7E3OH1lnO93Rhz9YWJxGm4tDD2o+plai5lES0miabUYw4Kl8wYjkPdT73ySi
a1zQLzIvZgr4FqslvoLNZfvaiGVr+8G+26DwMwrRfGA3TFR9QwQIBvNO8ejk89wrfdho3jg5dkAv
HZisPonQHhBosDWLBW3m6xFMKViOLdYSctxhzCHNYeQ1zEK/C8RQbBYyqiAxVw1gsg83I73TbuIo
hQ27KyYw3u4qZfXpCoLB+PG/Qiz9Yt6Tm1X9dnMduCyUilSIPB6BIiJBn1bGCFD68AbdEU9QORGv
vMBIP1oTc1ImiJIebNhJdwKj8HSOe280Ln7kj+WFp0vUP8zKGlSzslw+CYhPrQCdw9utwoGauKd6
Lmk7m9PcZg1jGZlP4zCLlLsImDr3+ceurmyO5BpvPTwIBjfDFe9qBrFcyI9i4ouj8wl1+B4ctxHz
i3gdi56wXtHQZsPWJMkbffBPSqHoAgeHbVD2Zo81pJL6rqMuS5cm049FYQ4/MLEzgPFTAu9kMqg6
xIMvWSyjWE8yXjHquH3jYLeTnWG9taXPm0blDPAMsOx9Dl8cdVnOo0lobiSqnn9bxLYGLyDOPyvb
KhDEKq4u5B5dsj/tBabf4BX97CkaUUMBytfYisjDwLNpD+8vY0Vc7ylhSA0G16k/WH16rZGa/XK8
NhgceJ68bagbQ66fgDx+rEnJBckoF9PxPMy5RztBimatBxI4+8b3W4uTVptziF9h3msnDfqm4f5t
jbGs7NRgnsb/n8E5+B/njdw+F54lpPuF0hPYKHgQPTyXvZyx14wtC+6qd929SnpEEMYoglUEKKxb
GKMA+UYcDWsr6ySSSpKg7xAlsEeoD2Fhr0TdNtsycNR+lQ1vHpnAMjXIu/2FQ2NFOP1avm0aeY10
zvD7rF3VNWWR5fULq6OoXHZX45umfZpaXrJwHvTTR6YC+LRqjQ5M5+aGoKQb8823QW4K2WYPO+jY
YHUZU9AR+8FLJ17s7o0Gr250okevPYQk13Wrdrxt4s8FnUYoqgm/M8F7+R6963IwueyUd2laoLP5
Zc0JXukY8wPsYPfISnshL4m6fOX73o02BIS7MOrQDZgzMtWweZdqbWnBKakDdxjgi3jgBX+9SgqX
04u68L57u81sKEug3E3Orh21DxytC+KOxmPGxHHszwowRIzVhsqnCezdQFYyxrAuwhXqPzh04N5y
XV/6uxakaKe2sI40p9eAtRqffpZmG7IWurwE/8xPHME/4b2PCVOwuxsLd3yPDhN1cEni8TUrxxMN
tjL3ADIK6UPDlBhIGJ3n1qFqRIJdfqd63itGpPtgL7PPivYawvv/AAM7G/2uoDWs3Fhfcn/Ylb0M
lbEafoKGN0JeQK5hlAtFkCzO94oUU2bTn2JMgHZJsZBv79Af79nzUzTJtGD+/krgBc3hDREPO4Ut
EV/ZQT1iy7ZmMw/51YuCGOdrAbJAEvTGIPIuLDqheGCeYxUmVmAfVFzpf2fxUyxZKbU1I2H/YxML
a2Z03+fUQGDtHDwObzfmuzfcL87S0o07f48cNmhwXNPkh3bwnVDaM0bifju0oilNa7o76IrwDHsZ
XvBH7Oyl7Row+rjXHpkH6s/BmzKmSuXXwyDbaEJkT4dRxQ//zU54/gL+TlxY7kDLLK0YFjrm9nsu
1hBilAqM9o6l9wPpwyJrH/iPKV2DdRl53GbhuSYCLeHEmP7JdKWPhj2PIdcUsGKHoBj+2XyI29l+
YbYhWavKlR25eU7DwH2XUBki2l4wJUWkQHYPGieoqJm6j5K65dqZ2fQCW2xUJZQxFf4i1fk7gnZ2
33F2+LgKKQBrZNfmhA+Uf0Rg3rFtZ6OqKuMDiHQMWIF+pWJBFwXpdsN+N0swYLOgZzKUhkZQxsjc
FZkRL7eGw4nZOiFwEBbiMOZ907TS5QGU3Q7u0K//hPdOnv7RI7xqoXyHubz/gELhJPEw1Pc+enhF
Vl9xkSt+5VkC/Vg+mLe5avFpQ9pkje26/OsXFh5IuuGM/IbE+TQ3on2wJSlGXB5sQa8LKrzqvjtw
jxE1W+5gSDTNdYdIORQWGFARUxRLcm5oz6V6+b9uB3XhElrrrJcgPLUu0ZJs3PF+yK7egkLQzv33
RThk06hX3RJsgDqfteb/KZwH4nMJKIdDn9heFWgyWURw6AdvQ/z07lD0zUvAtMPMavIBsNWyzQrG
LYI3yqPOSs8AikDPI+7FIbblkNe+WrXTsjRbkopSInxM/gqQFsBFi0+xe9a/kNUT2GQctsl2SmgG
ZVtg/j60g19dzTJr7N8QXqsBvOmRG+Aab7S2CppOOjPP8/PmkvcQas+TmqwSADAF3WzyYUuX6qOh
7XzLxQ1cnpfNN5if8Ln6Gwy1gGHdU3zvFX1AZy+34XTAaQPmzopnDLMETv9scpNLm3ra0zW5/fkC
8l1lVD9xOWDrpmU9zUQMdXyfJkDgtcJ8q79xZV0a1Qh0OT5Dehecnm3MrThYdmnsFbAN5+W37QHJ
o6GhJ41joYNsozmCzXGm8375S25S+c58YwXXZpNCPu4UbJiSoeW86Qr2BYLGS3fFjLxz7TQ6CVny
ilDhbFc+P40qE3LNMqyjNKW08G9bT9w0Yd4vIJBv+FaCqSwnNjHTKq0BbiVC5u/MS5C1jIRZKemX
wrEozc7QnQBTl4kVGQIvabOOW7PR4x2gqWlCXcmKZ49wy3GPH3Kgk/gP8o7pclV43dZVFWlse4ke
x3w6pcfe2v6SVvVbX6Y0AZOQAB3ps7iKlNRvMr+B35ZsHTzHd0f2CRAcDFiatn/uIIM1a7KpkzU/
ooWXBdHpmIxp5yUdfaOveNH+4fOdNF4UFPDTcz0P1205Z6jjKVgo2alG1A2uq5EecECkfnYwh5p6
82ebpghzChHRREGVGwaWlJtWGqQBmNj8jCh1L0Kxh8mRpoBhQ4+VjaDkJZIpEI2lKVIU5Mptqla+
oAlZsiLchgme0mqp5S9zaRTic8EduAP4bRoc5P4w+0ZICOThmgoZLLqRxtFaVlhPIHLpf90j4BYm
Rv8yrpcuSQ9KA925TFlhNKZ7EV3deJB7nxwx0w2WeRSlCCcOitqKXKodRZ2+9cUY1xAoKl/W/nzp
NxUonKH1gTKyXC/JqAuS97LEBqutx22RuFFIjn43pg57pdkeMQnDd6Aq038c3kP3eggJ1Z8M0Dp6
1BdzAeCvzZwl7oKt7OqlwpdTBQq+vvyzZYUJMIX19v+OsLakTS4YdccxlY7vt+9XMCSmNn9V9twz
5f4AaSEKgkwTgkWDpkUqoX2RIhAQrnNW0SX2ceErPE4HQg9DBQ38oMF1QjQbWjwjIiPFhuuQdk/X
Z6I2+EG7ZfJvQkGXUL0Vve7YJoXdlqMbIRZuhVLJJFUU1fore542HY1lVxeVG+wRKcrejRpqKhj1
VXeeccWQHtWrNPkKPhFSszINhw0rhMlWD09APyt4s5c3D1YFGHcgGFQodn1ZJOO9hq8Mux3UVV3e
lW12heE7vrDe/ddz3mvS+RJhm2fLYJAHj7T3ttlr6gpSZj8Ufptl3uSMOrCAl9DlMRtqhgiPHIY2
P0hp
`pragma protect end_protected
