// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c0E13Meacfmy40xV/1P9Hxka9gVIE6Vk4CrvDhV13DeB7FjZsWICQk1gIfpv
oZEf6qD6f9dUbRmVGqcjF26wOLoDDg0s2cRTVYigc0FLKipLz+pYwdGikXEu
f6cXDV3lEFlrTMptOAvHPawEZnHfuiIrvD8KV6MHDzYQ2juGw5FN2NkTIjCZ
qdoE9hhihd/h0lEeQrOJLc9IEdZNj+x3LpRK2+mKTr2Cuy+9iI0HJ3VG1UH9
+D5Y62ounkvppEJSs5gLY6a7tbfoXeFJqCYmxcj96SdkHRBhRpi1uOPUCVud
X9xr8oZcLTvSDwAYCDX7JMvyTXw2pSeUFDB9pA6p4Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cxfmRv3ZZ0TMYoqbwAOygaBGUOJsbFf6VSM0zQaOK8jGPC7tO3ewt0ax4tmG
SV4PSeJLjBRGa1xmH32nyJG4oqxihrX9sSJucaeNuU467BXt1vQjIJPi90wa
hOxCYN6gdrkQgZbOQUco5bxN951XjJTCa3W+G6CbVYDAA9yi18wSXDNbkjeX
l3YKefGqmTFGdWh+ULs44ukuUp/s1GYRlJEe8wVkIDW/v1Jh/xf+w+J1Z9fH
NVH0MAxa040fMw2KK4z0jffJ4nFCKeEoDvS+1Sd7Z7p8BH+13Js3+yuFOL4N
jZGIgk0PRerXBpDHXy4voV30HsM9M3fy3SYOwSuegQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I8dxlj4okouh6goCOVmZQs/G2SRy9EoBdyWd10oLIpsnO7yOo7XU4lgYBFcH
JZ0kQX51ajblzmOjkg23rpz7LkafYQ7yvNWsmAX5n93dSVrHRxJ3c7he4kVP
PQDSXxFSPAy+t3XpZ2IdiZ3rcWDjWymELjEqCrVYU0jpR1fvVXRzlmCumezo
Yr5GPkWFSTcSzB0ZMgB9A1z2AWRgikU/b3MQUr3mkv4ETmmhbwdi5o2ftcs3
/c6o5i/JOK4WdapH/eJJ6YoRR+o3OWpr50NQazkecX2kJq4QqtsH6u6zxU0H
E/lVlSjQ+R/Zh15wJJcWXyFX5p1N2VQ98hwdL3u71w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QaYy8HRwKaGBQ2BW0CRU7LdMiy79wBWT59unH3537rOeiVXUu7vn7q3HaFfJ
QpqIqJSfw//elqxX51rIDHvssyXJJbv7XAI9UTeflZJ7RKJYQsf+Yi0VPYPB
LVipVRhhqpyETUH30kKEO5bE2vtqyHSg9tvKD280AlAM9Of7sMo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
BzugwkFBzF7DVCr/w+K6fWDpMjK56puyy+Xj0F0Ar3C3CfN/8SrsKldquZ/4
z4ZaNnRYkLkigLuJlLk6kES8+DBebNftJ8RiOxDGgtQ/NvnSp5c987ueoMXG
QjYnbEB3XhYA/fM1o5OeleWFhScMfF5Otx/fCiB9VgEgYTMcs/EoA5eF9Eht
U52GBy6JRAOnDkBRwPBo6Src+ecdhNX9ZDzcGqqyeh2997+XpGsp52hvj/To
R/lJbOvcFCon1Q0gciAeJTMVUPUzVS3RsxZUt3f3lkKC6hJd29w0gD1D1K0t
DaqXABJzMAtlS+DMwoyWgb5m1WXl+Vig5uHkEihG7ztC01mNCiis2uSIMCEU
nY5v8fQCQJl+nKiyBP1kUOS3ajsT1NpEXh8oLdkG8lkEK1IHKq4WZb3yRCDG
nP62ks62sikf4dNT6rTtKI4mUhLUVswW41lA9lTFiIe2fhjKbnpKO85AQsmX
JKi1OTwPH4YQehKG1gTYCYzSozYccIBH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B8eMX0fO5RAWzv4d3EcA9OatQ4jkKZw+IzwB2UG5XT6vUFF5YyQj9E1hxaA2
hpR/djx5DeM51EwWRCKhYMLol+uFTqY2HZcFrMmytbxdN5H4Wk8jJuFLCr/9
Qbp7ZS/5kes/yEYKDAq7W5jyHmVs3ipnlXD6JD/g4h+gpG3O4xY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r9jP1QWYP54hPVj8+DImjDWMqWufhZW/Tqv9+23sTX1E5KWgMBsEndtm/psO
vvAwrT/u4Ia8dnexi6XQin+tiZ9sUoWNaKmGZSosJb2c/ksfn9T1AHr7YS+R
XM5aPaiW+V6U1EYJcDS04e8bpX0e0AQeFSFIBfvDdEnRe26Gzbo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1312)
`pragma protect data_block
BJAt1MEWZLl5Qq1AnNuac4G2tUJ7WSGUzIIa+F7ZU2bRbbXjbrs4fbbtAacV
7ExMAvPnDOS9QeUZZOgZYpnsIGZ2IIYLv9KqN2BQqp1W35CAXSAvrDn/C/Zd
5+94jGlCDxu63XC3hfL8Q82z2q+BE64F9ZrTOOyCC+gsaCtxhfw049g7RJfx
+rYboeXilfYhE7GWVZb7p4ak/pid8kV/cPA4+vDn/bj3PMPvMoun3AYUd0UJ
JgjmrdWMBhLenqqgDXIOzEYO+YKmNApiqyfx9km62X0l5DO3L1DVVsQkwuy7
HLh5FgCyj3H4YPEH3K7eGGQLSRQdc25RrjyJR29iOUpv961rOBssnO9gA7f/
nWIcqDzKfj/9VumjFZRZxbhZg0ONHKofUAAfQ2HidnF7v0SPukyZIJRx5xQa
JXAapZMwF7TgiViVCfR6EUk7Ib2f1FarX/wWyaTFYD1LhEt3ZsDnMFU7yYJj
tT7U4WZGhw4liDZPzhpkHn/xegV5lTlBI3mtdgIak7yM+odALhZW1xUJ9ldK
KbUdKzw0pDOEYv3UtIIunQVWiLC+qZt/MoKFAa8XJvUh8c6Y2sgrbC+5iQpS
2N33wdF8Tz/iT/QsZDxIDp8Ag0t5jZLtx52P+m0ce0KqjsQvzZFX4GKUigIN
v8y1Zqi3GONyJGpkXdeOR9lPegS/onO3BwCttwnblcSNkkXy9uhhvOp/71nt
Fo0jV+R6v7vVNXGBVw0ODT8hTTAQz+I9Y7BIEMawz0osVgYuQ/cefVz9pLkR
itsD65XHaEXTXrUjrm/GkpXH7al+VAp8f8vAL7FLQU7XzrlpDEztiNG2xL4M
IMiixMoD5XysBsJtZzlcmF3kdMm43cyjuwHIpRtx2q5t6s8L4+Unjr+prMny
tZd0gjx8bScKiZj/wfdde17gZ8LYGR/tY5ghT2dW/81Sj+slyyMzc3k0sXAI
P7G12MfAEVMy+fTzJq+JHSoHzVwIvO/kjQqVxleJM8xmxW1/9qk1sbsmS2oh
uY6P56jqScF/0IJqiORhofPnfuEsG+WrO8zxjrMz6ksk8aczvSQMxpcPPQJO
91DyFRtbiE1k5nniyKP/j/A3guzY8QHFOfchE4Vhlfk6CkooBkAkbqZ8cYaL
Z3I95cIcLJhYy+rOrSLguX578JymiAumm5RWWR4e7NB0nTT6meLE2/mne6Zd
KpGhztvTQyBfuAMjHQK+NFtg56OY+bPnY2//sUgROoUOSiMSQt6ClEK9k2E7
8camdQprWk3chQDceynPIyU/TKSHdzNvTnZgWbBzIgWSqBK88Pr23YiKbbkc
2l69BNQOnCh7oPK8CWz9NHBReCKoir1fNR9/GscAJynsJsWt4Py1X5GJWe+P
us3D4OlL1EQYmCjIrWM5Z+8gzplB8zJq513ASYUzLtciZiHiFA/mCZ7DDiSP
kYQx2QD1l1ckHiHpAWKMKrAdf7cfeLvxRB4m5LrJmptQ54N9RE3zltGnOgj3
/giCwf1aZIIWTo+wLvPN6uL4c1BH0L1xpJdKEO8NutbjXYUwmLH3yDED5OnM
zxUdtX5r5YTCoZdfIQy6qzivtN+xy3Z9+AGpQxSvN53Fwgbmr7UzRJ2B546N
Q6+gmsj8HxHsNyhscqrxD8WsRB36MHEwWNaiKgyKvOFNig2JEB+xmva+VAwa
EOV0zoo+CN3uVjgUx9QkBtiFlTkUCALMej2c13zUGDCkIWiBJFOeB6sOP4NB
ZLzYblV3Kw==

`pragma protect end_protected
