// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
yZtel5P57NKfZy1d9TE8PQv6ArJUyOxg2XvIjmKFk0nOpRSrhLbRfxk2Ywbw
Ibz4tKSViGQipnTqBLT+b31gy79zlB/WcNIM3ePaObMOA5WFokHHBKg4r84q
sDMMZio3pGxx5/1Wp9jooOE3jUcVFz8igKN37zXMVDtFrheS5/Kg2Yvd3t9k
FPv6vGTttWt6D/Qt8lmxEgMPB18goYTz+iU6tpEQZYYJ5yTOhj2M2E98ald5
4tlVY+7/1Ds2O7vYdFZQRJDax1tjY4GrBEdPecnntTeiJOxYTBMp6nQtF5k9
bYaoJl4NAPv4t8gKb5xNEjkKQ4PpyCt0ES/Be6Cuyg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RSiwfVlH0xm9Fr7X4+hnAMRNb3TIG09vTatzABBn4sqdYCI061ABWuy3a0b1
VOMviA06N2IDumVYCC/EyED0xbvqR4200QO6/J2KHmZ7zdBJvrCM5UPPxsR/
n57Qa1rxEgCEKF2BtsImdFd8M6SBP9taF7pBP2rJjdxRfdFygNMtFm2l+fnz
c62xZOvbd0Fd8apUaVJKR1TvfMkrvtu++IAHPBUA4rv0mrht4EGWv8SIx+7K
ho/cXZu1IsK+2hTopJllz+Esy/Y9ux6kL5pB+h4+sh/+qAS6B737owCDHIUq
fiGJr4E14AJGIM+9hnhYU+p75Z3JoEFCV6IgyYqZCw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bywl4OyJDNw63mUSUaymWnTy78HntIWYEhhPcIU7G+HQatmhR9/A80JdhX27
LEozxDN2dRv6DDfiUhDPejFF3thy5qDXcbYl8gzYyBgXRYe0OdQ8960ADvuz
ZfVMUOROk0EvdWMAjNBf62iBwP5bOpMMjEpn/Ctz16k1Ne0JyLiQOqplfm95
VMe8qZoQHOGAk5BzKTXuLVUyTDX0Px87nAMJdRlZdu+iXbzIESbpEKkAXLYJ
73fpOuas5VB96gQkyhhPaGRe3gFBvaNtCIucf7xkZCGUSpYDjNp6nKbVslT6
2ayue8SQAyxssMVzq3tCLgnC5kZRDRiHXEUypC3zJA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q/C3Z5ny+5VU6e5R5rCjE6G1uZGvPjzeFPBGC6rICg+a7iYmB9xOzLAx7LEk
gqGk2RmQfarF/HtQs8fl+jjmGrJUetJdLDYzl4mI/W72HDdXQJhlG1G9UVKV
Vrmv1t17D0wblLeSrqJnoRd1QbqCcL8Ci5OtJnY9p2s7I9qJnhw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tgKEcwCcjPnldbQC+gfrSpwkX3sYDIsdFfR48SnZBZ22VCW1vkYPA7OvweTX
2lOLUxekeP0SMz9GSvsn4eeXWEablQvLg52SvkfmMfBWcsu/ovi7WzSAJCgI
1XIrKn3PYwNG+J/brHtX9WjbbFaSTZShWJGW/TIDTbPDUgl+A774/DXFXXny
Vjzw4+zxwD1tIVyuN6d2R7BD3DZUtwCbXf3j6R1/n19/VY1K1UHQkq2B9Z3Q
1Q9HwGoIJphJZpBHG4PbqpPLYfYNgC0P7mhW+UYUpqsC8UyJu24GwkBU8hWC
n9vcKbZWWlzTBWS6TX1XFImNJNVn5jCRKwDMPfUdhH8XoeQ1v8URjn+v4Mv2
UXZYfnTVOBifOd7sjX4Bw3WM15BEqWbsATZm3by0/BwEmKxLUYURgSKdBXkp
rGY0I+udgT42lBEPFtdNRqywz9Ecjz6AgleTAy+OHbsUeSK0uFmSl9wk/yVt
D9VLz62r6ycltoWvIAoJ1LnDOKWYhuqy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GbJLUqHQuQ9f/be6eCNjeNyk3oH9FjKaHIZd9A7XWf7ZeI3++mRXBb+cuf/z
bnPxTU4d7BcvtpYVsqD3Jdhhk9TJIVYReVt0QbZHwIT++W9v0ue1Ese4Tk8X
kuXCggfKm6BuaNyXWbI57mTS03i23TxPL0ex6MpXVhlkPwRxJP0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Khdl+dqS7P/guixlGY0agmLhRi199jCz2lIx2CsQZdTYI2SjoVbLtd1uDBUT
PdzyStF2IUSSg67JOs6Tci/2Ueg8ULFA1HRAi0D7FRrm53N2R+99hyD1ggvw
dkq+j06o7joGaOTSoWI5L7GQQ73XZ4ZfQmrMM2uzmM5/1ig9T0c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46944)
`pragma protect data_block
OivTdGat4CN+Nw3ovpydWHhVL6hu3RizXw4hPMAGV59vGSz9Iljp3EsFerey
/BMkbEVKZ4Q9zT0ivYrY0kKNCJs77Neq2V2CdMiGi4GZKnG6G9iaD/OHj2K7
pxfSNBDDWJQy7yDmfxsp6kUYGGBymHuozRNEvTGu3xXKSdhE5WwzPosIT6Tz
Nixb3EKZsKpIsekTzBTN1PX01JqR93X5pwyvPJy0wtIB+SLscDJfu1zA7BJ7
ADO6H1ktdiXYLFQFwD3ZfAAYS4ucW9wW3dYcwnYcFumBb3xrmRwm3VedVOMe
sgtZWoumll3tSYjiRSmdmR1/jW9bVI+spqoELGCqWwMcfLpEvD5Mjn7T++Bv
PDBWRMh4j7ciHkoUkF9uH7wKthu0wP8ZAiRilXdZymN+aaLTPxUz6Wrg7DPU
6K/FXjzoSKGcCW0u2c9r8AYkooAI19/WJ+1aVSA5Bio0JXMzhgYaJ5/1pgWF
tBXBSzKXJ7IwbXzr/be6oRQaRX9ykGoYXvqZ/LMrTwneJTMnUYHbK+Z+qCe2
y6bqXDUXbpQg4RZx8pvXQ0dlIgxQ+rpq4RZFpFl7xYU/gfJLT4jr1iR11au3
0oCRgfADE2b/npoK5PIo63tgfNm9FVssh6GcOvmmWWzI8720PoFIwsIxfGYm
W4DKV+68JJAwUhFbsDCdf/aI7V69sLfzr9dLdNUxu36YGWvJavdlGKXljYoH
w9FubTIrvAiyKcMgsBqLLFvJ79r4r7P4F1yxiQwsPtFV7vlmQx9igUjvOSAG
G8CFecUc90gRCTi5brRp2667Hqww+LP5Zi7bGwac1urDfvzcvvM029u6fSLQ
A59EU/Yi433flLBe42h1tMY+V0EqE/cA309GHdjcGJtRkqq3VP9fxh9x7mtt
AKZeoODHa6r8DEq0U8k9lGTiiu3XGdc/ZB0utWx+d4p3p69NHnFm5BZVuBS+
9W/OB7jKllMUJWihuw9giM2lx05d6Ym+BCc5M+EkUUjxRw+S+MlJlsgRgrwX
9V7tkyb8sMGHxf8tUEz9KxLZAZ9UmC0FlDRkXtj0X2+3kfDw0ymdnnKGW68E
1BDPkkK0zcE1Yi+OBF7g24eez7s1MBiTK6KqvdYijpxIWicrFTsXLHqYLXgn
yRJh6XPCCH9QCcOmXgJoMVAc+rssPOJWLraIS8XdUcJGM07mnoeobtw7F0ND
vq0XMEw9HuYpBlkjaNmW4bxByV5j7gpkfVP40iVk05YXCb94oKmqv/q+s09s
XA3BEvwugmL0E25tfXnWNOTTsMAkOoqI0dd4GeOb7RkzV1bWUBrsdThr9fJn
kPX4dXkx/F3zScIFaaF7rsJSPsCpijiErg9dFXdKjT6hrT8P+MkvaIW78OAM
a8UcMcwiFHowk7/eOG79l2v3TIvyNBVp3+Q+gWWLf66AnyWWp0Qpks2B23Fi
3MQGE1qeJ5DdJPSduXbl6co+VMRJuZOPo9Z3R27b5/dPfyM8NvCV1TUmYC/K
+nYJXVcq8bTJH+mhFeD3FHXT1xfi/F3bI39b3gfOb46MaxVy+I1WTvSIPXxX
pIVxFGL9oVvx/wvsv4+hW3FCBVsKBjeX11U7A8oQ3nF7ctsroXFBvmTbFQhD
y8ggWsUHxc0ZiH0ugNU0NGVeX/scTAryWEcBizsmwniwXQOwxaUHU0YnoF+Y
m4E0DuLfvtWmHsiCUf52re9bZMnMniTgxDjz4hSe5kLGZQGw6nCtSxy6Ol61
6Qj05xT3g0d7MTOviJmmo9uD4RIw+4Ndd1pT2QhhsZTEks036ZIUbTeqwCCO
iZNHMwArVuh8fluYhOuNBboWQB8lluBN3DEo50ctIMl+PnAJdTxCdJbUJTJR
ZjJrv3H+F7ciV6zkQk3tLr/pdQEKth2HdrwC41VS77ghhsTsakHp/yfUlZ+V
0uKKZ1bxruEBfh4NcQmbaWBjAgVC1EX+UCh/giHD4yyUbNd4c/T6rYbZyPD6
pR0EOUubVWJgve72PSauf+vlHblnCmetW2vv72tAev7ETTg5Cc1ChIxrXqvU
uq4IBzNIZQDgpIghPn/17KaxAWy9R8OpftXjHaGdG/OrOIZxZdH2Au+hS7Xr
il/CrSNwW7K/ch0/YjDjJdCS//fBSTcXX4ubqdupJ+3IgASzr6G3GRDZw4Tn
z3sFbSZjMh777LFivxkRyMxLs9nQ0/vq046LSPze+yFYszAjsT3SSy2nJziW
dFQLNFaoLnQLdsFwx/8k1xCOb2Xdr9i+jO/Ul7YvEAttcXqvHFJHP3q5UiHo
0G9DkH0/+nUMzM6fsxXOoPWxKUrvTziinTVhBbPN7v5afINFYZUl85QK0Pr8
7/uoo+JYILi4waMsAHJowFFc/D0zMpkDrwl/gpZKsCKOVlru+zF4qwJZqq8Q
rVsTQAl9ZBKOown/bKr8mrlwXVI5nuWvNUm+SeRAcksar+0ao966VyJAc+4i
sJWoehqtG2jGEgoAvxEld2oa/YEHaTfBKPKNIY9+uHfHCMmKmFOjOST651L8
Zek274txnmaE7rbzkqnDoYosEGiP6FMUB221CbNNWb07RSY5ET2aWwUdnms+
gy8OwLCa7XKvHxkRkaqXZCmw5i7I87LYjNGcWO/8OwKz3PvBhKbepEhwxGiY
a/wG05XTtMZytur1XE+pI7pdvfMPcZC4iYeO9RbfRnZcWTqqfULVhzF90Mx4
Dwk0ZXVSDTA/SIRnzocrguP3X4lR6rMCAYZ0JL+xgR5FbGQBkmiX2d2AFWiz
wM43BMGPKqAEHNd2t8TCDMrqNj3nT2ReFEmirwNX9AMuRVBYi0DWyLQJUdf0
rRbT2h4+A/hhKqo9oHqwKZKY8iAXNRpRcPhVV9rK/oimyRu+KuKs0K7CvKDm
q+Y2HO8kMXvlpd8ys/hJCPAkOd5xRn87pae+2ijz1NRIVFyN2iNe8Eyxz29d
810DLWMkhSkrWaOpZslDDHuPhhwUJRx04ef/4+70ipR1CAXq+dW485bqonlf
JVVFSpDSxxplmpqwKsFzLsF+KA/O71TaaUHl+WmXlx/KG4lNvIruou+kX1vh
rbF+AsajtZYCG2t5sXePfHNVN1Lj3gvePaZVX+eCQX3xbMrl4uH05qiBdbHb
01TdnF6Tbhumnvd3CTFMKf9/R4dder6KZmUkkpx9+ExqLw+DOdipaKdbUBrq
DnjdFVc/6BWew+bGAazdiXGWkRlrAWKu5d7dycZR8lB49CjoyeZl0LwTB4Qp
O6ES63H3qHjOrEA5TJaOuKvd+qfC82f67Q1gW0W2L6xWunnFk++uBHKEQYPY
Jcf0M0MvTTWjIW1XqQ68iC7Gkb0i0RU1iDiUWemx8sLcgN8zd/mi9BBGDq4E
pyJw0Y6nrXiS5qW5xuo4HbLeTf37Jq8k5PS0LI7oAdU9nZ3GYvTbCn2YJX1+
sfSfGwhj5o+bBJO4x77EbnPJXxiqwvu2wZo0gc0M9lvW3l2UtKS9TQ4r8wBN
DMv440uF5YvRpG66Az2mTHujC8j7VotDYHk/9opXXrs2VKj9c9JA0bHcy7AF
25kJWIFGeiSwUjpsb5r47xmoMAi4quMHVEdKF2iv5mvzhlBJIb6ySZsSx1uj
naNZnhBmGK72o/yi3jv1AMQ/spZB9Sgkng3ahmz3tezWwKLw0A/YMJtbH8m8
kBLyAKQkUQjN1TP7UtzA9w+m/OAErm1mLCuVxsHTU139W6UuuLUVe+JqocG+
C9sZjN+LC44xCxqpYlqcuMTjRAcv3dQyDfhO9VzSD9nnVq4voRGGFT8vi0d8
QQE/RtxGTFlqk9bs+WU8nNMvoEgRPmxIwDCwrV/XJt8Y1XfHjEW64aIFz0sk
lRb77GwRJgbAOwbQ/56XoZVaEnn3SdQsX27KMwXWUrcL6q0fxLJP+2iWmiqk
N3AxcOUFX2vSsvSTPxvtRKakwnAMcOCSwvpTsODJoJoc7yxCVHIfI1pbatea
aoGHsXvOi8Rs9cF1EoRFbjoX7Dad4f/Q4ENdud0iOa9gB/+5N3MKBOlKZGF3
PgmjtsAI6B5FfNjBlr2EAUP9/xpXzt+BKhL61Q0cdXY8CGx55AkRf/VtcCaZ
rUES6jyRx+DpC3hhgfR4xUEG78JUzZ6XnYQdwV0/6J+StQt6r1rrwGTLuCGR
KqHNIcZ/bnNoGPUcgIT2X2Y/qrgSviK0N7CK1MsG7UQfvILReQx1rBw0vOC/
1i1TkIg80tdrqrK57Apw/YS/mQvXkOlt3ulrKc8yhZyXOEgoGMoz/X/4844p
kk983DxyRiAiN2Txde4o1T0g7QamByTwibrzLzE34qAASb7DZ9UUFI3bu523
bZj8yZGia9jFPWTJBTj4tn0fyxWgZk0yy9dMlqFLQZxo4wKZr15MECK+Xfyn
UefDvrE/BsB20o/L+UQw+eyhDEGtITm5z/MM/PPiSVwQuI9+o2GjGx5V9Fg4
UNCcirO0GCkWib/UXVWEiFV045R2wGi7256RDeDNuKkeBBZ+T9lYE7cSjdk8
2oyjAoj1PbcZ3yjrh2pBJxq751NBvZqoAXfhc6IACcxufVfv61phpTTA9rni
BXcUsAlQKAoPU1h/I/aQF/o/zuHfk6/plF25IcDd6vIqYcaSU8xAKjK0Whpx
7Mn07gQGrta5Da1nJR8GW4b1CjZfR7VFNnNEy7mzp7SgwsQ4/MeUgvjMbm67
hy5hdLFKuZqooORfzKhXYd+2IbdegHx9coCorPkO7re7UUZ6+SYzKDlSBo+7
eW8Et31RUsuCYc1OJHxMlRL4EznldV4GwpafKgpjJrWdbAs5tT3MV44K+SWV
rXh5J5Le1OOfmuWUjh9xsLAH/0bulbCkK0XtUdxDPjtXhCX5KNLcli005ued
Ab44zXRJCoP5Bxj8ImOxvalLMPYZdhNo/aStCfrcGsljc9g6VMg0ywYSv0aU
/x2Fg4A+zoKSY7zP83uAnYceK6Bc6NYK6eLx8iVj4esLYt6oBCS0G0ckDL2X
AszTKNleaxfh40FAd04EEDRdJ08V9olkLUHkY/X3f1L1hHxRgxzkYrCn7cLJ
QH9R7m/W5p2E9qYxu1kPDI347Uk16ri4D40bdlP5omQNmW+1T3FDdG0+Tw0D
28i0NJQ/u2ML8EUvIoU062IFj/MOUVkQpbPl90Cdfzma8oxKhAC5PkYl80Gk
xK1a/hQKCCOMvjXS0qU/i/W8TH5QvUHqKTkoRTRwVAG7Oxy3sH7WUkRUO1Uy
WjQucGlRxllk3yRQ1IQbaSxdZnoa8u2WYRtr7g1fG39imI7/nX0VEKqtqak8
NFelYwPtQaW0PHSfvLNTi65SXRx5QBZylBPXKY85sTX+W2nPQmrjoeogi2JU
Wo1foFJ28oYmDtzXIKgjjwUVnM0YwfDcw4SuVXmnqyyQaGFfCKwayeiksQuG
8X4omE1jTTsqeYhX/xE+nE+yyuSQUXQ+OeDPXffs5V7eHMN34XtdTQT7GPE2
UsAySSBkBthYjhzj0QugnvgjfNedxuI1iZ7OA2MsxPImIL54ERh0y3O5FHKv
Hi4imVIfWQtHnfdoFU7nqMIJOPwS7fJCR5driFt1ct/+uLHPkQcLXCy1jF55
FsN+fa8tC5sub50iSFZ0V8ooBOTyQHJPig4tAgIBjxiUaaajjBKq3H5bkRNj
ZC/Z/3X1yH3Vy008ctptLZ0Bz0z4uFh3apiaedIWZAkCmynW8svtbswB4vOW
1rUSHv23P8qWaUk3jRIr4FkHQ7VVDjBG+HKgKpoBbjcJheD8Xpxk+IYzHFkC
uFNSWLwX8UrkGur0FoJX9JccTISS3Cg/RqVOPkvmLEG2Y4Fj7XhBwftLeRb+
SaR/1IIVBYgGuGOdtPcy1UFS2phA5rbUdiyMEkOY+mAYiIaBlF3WHmhHLrDx
gJryy0lLtA3AF1EmnVXX55zSbL8/P/NmSWrvvTjgh3rUqA93sLAnuYKqWiVw
oFjFW3arGnVk6Yt2e6cyCcTp8MUY65T7tpiTjlUz5XfaKHzD8s5uOBaXjSGt
1EY0ricjc8Dwg8FzXkdNUlBNCdP96rPYftmXj/lMhnOg+hr7q2zx4p1b1ERp
eddI7Nc3BNLx05wm8cP5rztbDinlR6T8RkEkXM9219ijHWG0747SbRSkiTih
u+ujsKefMwlaTm5z7fPLTtGd+Lj5gIf0Qxir4Tq3r++RVtGm9X667mC1R3jC
M6KDPlbmFLWdk0wxKeazoxpevx3zIULHJJ4MzMZhLW4Fbnb5VABS1rNLbKEC
4rkwrIB7mAX1XcZ6MUoOq1vJgtGAFOqpJxceCSjLltRzG8p5xx99Twyo4yct
ZR7WzJZOskOYfGxi1hUGFVO6JYWX7E/48ZhJvF0CMqTPQB0HV9qzGHSXSl/j
9yDdo9dDsvglRuVMOnQJF8YCQjr7He2z7UNtJwn8uPCOcw09ETLVqaIR+ECc
nFgcKffoH5DWvW/lVnxLoN6966qj3EzU9L38bXr8052lF+o4KQxkiOr+Q78A
lsHDXcJXk8+9mvI8jEi8vki+r2JIa85UYYlnUEfGSB3oG7dNWRYvykOL83KR
2Tvv/1J75/0c1Zuf+qyLWu/1t9TVSRIxsPE7wslB20yNCh4RXb5mdpbJ7Ug9
btc5pv+0JeU2jx0kKdoVouDbFYnMQFo1TrNBBW57ICUZaI3Rhz+ekJAjRTRW
pMa+Gpb0KaFa/bKGg0ekmyvkSUyO8u/Hl8UHxifKgs8L5Tr1Dc5i5iPrHfbO
8nEJwpzkca8LD9FqLX621KnO0bX7SEu6FqTAeC1vyoKDa53h2f6BXNat8tFb
tp9WSg5R2wHXklNTTHiKcTEudSmPJh1/IyeW8x5hHpQENZCkAyliEzpZOLT/
P9W9YnmXU1deHT2AqNPTJcTZ7jcVQy/kC/2E2uU8981ECnjVCe1Xhl5fqyaK
/tY0fEtkXXaY5u5ebfV8cAB730Pg7EEmKWQhbBfndF7/PRq3YuQvj61m7VF5
WvHqxU1Jy3aXnFIuqP6wHptKVuIEngB2oQqwRIoHXfyxRT7rRRmErvEgpMX/
4PksLqcF4ayPbNU8mu705IMmP2Ue7E8u6OI8lGD2H5dJNuFCmxbqfylgfyuG
YuKeKUlGf9BK0bJVjyCzUOvNBfKN46xD4SPublElAvVQUHphgrt8xSZsQvr8
Xhek+YMaVzwtQRZghmIiAuYnLE3G5SJ5FI67TMvd/gSy/2a1h5cHpQ3X4cYe
CAgLlsk78RubF00/BUz6TfaBKQWO3+A+yWezchJlastJZtxaPvsfh9NB/JHD
qP4JXCfc5ySEepIurA46br4MF5zWPMgA/TjmatZbK2VkRVjWFLo1Xg3pVKpD
QPRZuD4Li2IYHZf/wH4pXPhaOQ7fyB1Dif/Ka9PHB5aHBGO25R87wO67rCrf
Vd7z/Mvevbi58T8xtmAEU6F2+gciG4v6H+FDZG7ovcxk67//IUTN2HUZvtM5
4SCp3HSL3pYM9lyRLbfpyW4aE1u4Y8NEUL4/BqxSapze4x+KI3kw1BWAxcqx
oHNo2uM4R97R7cgKQiAohftD9OgkdPkuRtn/1zTURiKeNH2fMLrxLSRCoG31
7cAqXqWgvZYnJQK6P/cCSmuIl7xQ9gpu5xQlkDv/j83rP2K4G6wKPLWzF4KG
Lvfw1H4YOQM3zqzhNcfX9cxKfbkU0UdtUL6g1moD0jh34MzYnDCcKQswtRD3
0YP6eHE2F2LUP14mprTbPaXXWGPRzXQnZPUltnWqY0vBbMbvmLfjYYmjVNGV
v4rTYSBpM2k0DRxTmI2iMByxnpadT8Rb3buNI6hCuZEOirP/A3T00eaA7ojn
rvcrBXCpONcnhKKGG11cZ7uQyJzVMVdzFgbfmeshzGTDQaNX3Fyw403xfCUe
x7NUtOUK3MyT7XX8yCSFSUcm+K1zCthzxq8vlA0KVomsxwv1rfOQxpL8x11a
A+mwcgODT6/TlNFilpRp0S59+fTPUZTHwvuTZSnvwbTFDAID7UaFzw2IHOwU
AvYzp/26K3P2qF7j6I+h1SeLH57yNhV4SGVW1IMMckxsQHYpCytGn8lGvZWT
Lfy7CKw5MgSMw1vr0atiBTdOlPO0wknYvetl5aiuQrgZ+YGpmQt6srCGG/bL
Mu5s65LeXmmPjY9vOE7JqIdIMrsYIR+ol5x8TxVD25lpVAkPBIDG1f0leebI
GvAe+5uValCD6Gl0Bplca9ZUJZ3kogaskxSpFm+0LDh20Z56wyNUpT7HJkxi
wf6KZPnT7R7xnyjyzutkYR0oOfJzeF8vNIzjLQL5fo+zmRhhx7vk2z81PGuN
66LnV5i/y61ONuA0kB4fNDqYUfYwfc0TDACT42YekFResNgtuyXPnFpmVLHh
l1bda+bjxuAjuW2bh21J0vqqdFHSUTSaOp/2kqJ2HpbXbr6dLMs7eO+yTcTw
JX2XcoAsQ2aMvz1qqRL/AWlm31wdrjFDzgQ5BiBNQ7QtJl5LVzYAEejVC/7t
k5zzK6izdzZhrL4xGApRoVKxftQpeuV1qwyt4eoVrfOQgldMQAPhMJw+4hGa
rX2eSHMnrSopB+LXk2fu5CvxARA2KO07UDqX+jZrPjuvTAQS+tBB3tYAGBd4
zNPc4cjuX6/gAfgovOrlomw4lebYKBIntdap5RV/7WsdMBElRvUK4qpxl+t2
w/Q+AH0dh6F7IfAIyyUBF+YnucUMchbzZeNkXRjiwPT6TM31OVb1Lactgv9C
oeWziOyTFnX9zcV4qTwg6aLPAhbt2uO0uVWxc29afxAUzG2NefXwm5u/IiNo
m2DTzRXPC1HTVH9/IBqNzBiktur2uf2kLMcir1LAiZG+W6yb0JTpdue0HOAl
OBDXWpFhx/0+fq8wS88/kgPpoRCvRrcGKDAFu/xfSXMzHbpkH/Y0ocMQAAjP
qtt89nbkOKTVHqR9tPgwAFO4DFJFtoBCYXrFb6lXtGamUVWP30il7sCdshJt
sZ/h47mO+7xiLsAj5jDwG8FzaJQqKGGfVEKWgAYwMlIPkO+WdVO/B1hqPxJj
ldlxxVHJYAJjHVIagVmGbZ95fVueLdEabAs9Q4Xc845BQNjzJw4+ItiWi19C
VatNFMUAAf0mzFUljYRqcPzkdLdEi6xOYrdhFessJAipr9K2SEq7NUq9lonv
qfubUedAuo0DSJiiKreH/pUB/pIvb1iON+Ir2+uNnngguAplc78TOTbRIYGd
IZFX6JXWNCTxBwp7x48KZKgJug7yVOlOilHrxEQqEykIZb/ofHVyLSmrGPmG
G9w+O3EWXo76SZSFsEovE0I0lw6VGsQFoU/Iutfu5z2ZH/0WjEuJFTFBQtLo
YX2oUP1QF+MQbvRGJNkhNF+o17UIaotxl2lIhZTgTC1r4hAQ94BQZcWNHHrf
Og5FTWSCUL9iHGuW8yXr0U8dHckS9eXa0Wju/Gp3/jgy6dT7d4SQ7ccEIr3P
edrrF+dwiwwIi3PbY/uiDeMcVxQjPgmYgrPoaiEjbj6+5dLE2/8rFxq6ByFD
sUSibpAzcbk3bA/K2s6HBWay/c3AuJgkVjlvynCGLAdqkYutOdmVPRQJIZFI
PdPIi9/dBkowIJ4x0xoCetGo9SJDGXBFo0xuUOknBPsaYIRfd4+CJ3FeReG5
ZjHfA8xR2+P70L5lN1kjfhU0CjIkZJLcmo82AKgfz26iP4Fzo7Vzt0WGgV+L
K5TKNq+Ng24JXWUkwAgCXfd6Msl3RNorKO56dt5i886ygWqdEnVDyaDkntWb
V0EoTi9u/NSh5P9qiaQbZIsnEwv+Ih1b8l+9jKqRTr19AowlwpOkLg4iazIU
Ik1aoauixB7hPNqpU/EHV0q/sJ1+TS7cTjhtPdokgEjj1tY+wCkiwAPDRbXN
ikq05ShQQ3auS+UiMrpIB3cM9pZRyfrR7sXJCXSd2y6p3msvGOVs/GXMhZ53
Y9HmuOcsnywfa73Y4AZt3u8yt/j3rJvhETNgVJEnp8g/8sFIe3WGbDf/LU+s
FPe3t2bUB3ROs0Z2Pvp++PpcPHP3rVy2CSjzTUzEa01n+GWT2dCTXFPdJ3lP
NejxRuTUmBp9qYuiXAnhVXHBWt1WEFE4e5ZFFMluAgqofQBu0PBpdNKJjjyx
vd2+P23dyZJ5tgxDRuuex6SHr+kruZpH7fIkuG5b1vAdhp3ZPatJuFmx1Dn/
xe+mcp1lssUIiFmT52jMMCoEjsN5BMCTixdswwqnmiJxIJF8IyT8mj1CBbry
Cwd9d+K8GH3SgUjKcfiR0nuNfQhKNJkVbM8C/wB43pnMj+JA9ctouDM3jhuj
MpFi06pn6U8E7f0881klNOtfN9/0WL8WfUJFaREU3bJdxv/u0qUIWxQbV8UC
pjlB0agVGHy+DC8opFwYtxGwXSfVdtd3GpsjhfiMobewY8JkFiXvnDZQ26wK
KH6VgZmnVgjKmSj9ofj0JcmVf4i2j49aVuu0vFXdZ28c4p51dhsqEKHBLEzt
t3430UNrYd6HfuoYxU+NZbkeeo8XhgZOAFIrILq7szb3m4qrO8DhJtgeQtIw
8Pl32SSlnMK7Uir4I3y1kyWHLLrV7I9Sfsc8q/pU9er5JYfjO/+H8WZqJ0/Z
H5bQJSVM8/2hKb38CkIpiTesqKKBGij4OFy5bhNnP8PWu1m56urGbC2wh07G
JxsQC2yoNuQowmHPPaPTYF3IOeRE3fyyFN9k6k4E32vWfwBBBKbZIrlPPBjW
KatxOJ0oFucbA+2T4nUN9/D23hCz1pVVPPoCKjRIGHGaqEX34Q80/ozJ2FWM
pohAb2giomiaacHa4dBMjPnipBKUU7vitM2mLC220ObIomJVzBJMC3H2QyEY
0CO5Dwq2FZBRKysamj43/MgDrM9tOhQ8ZZGrPCjtklbBy0Arbj6kdirL62Cz
HCUMKHPcPTJHm7SukoQNphrvazuxbjOPprKFi/JB1igcJlKrgCY2rroL3JMQ
+/sDqA42NsV0jCwCavR9kUH8jROUwCyn5rTJbEtahcpRoG13Q4e//IM1TBqu
AhvxGwyO8AerbeZye10nbxCBcmH4vR+MCcrIaIUAyjiNjYbAbGe5E1WO/FYC
kD/vjED3LV4wsnjCa77ENofPXyNC1+Au9XfW6U8CC8x/kWOi4U2uE6/I6NYx
qvq4vmvYI0T9eUukVYPqUWSUSe1lYB1XhJZNbkavw3fF05vs1rZQu9hIw4zn
TVXFzut/KG//+8pUiUq4xw0ATYSbS6IgFBk00+d0wYZ16skyJ6Zic99AOX0z
4EeZNhsWdPl6E89IKOEUWjQfLGyZ1TvrWv7VQjtOlGAr1FBE5AgLZOOgXugi
Q8h9BOYGqLsTaLEM78D68IOCal0mauRGD9TvvJ1RZ346N1akYjsT6E5jF1Xq
NqV3DWKti+dOmHVJxmPjP2ZUL7qD8VFZBAZ16SX+9pvAX51rYMPzxBEjT0CJ
3Y9uNfMuVkSqcUbyZkQVRNMNm7JVYp8G6FbtdbGPP6vdAm7EA0oZ9Zusk+tU
mfj0mflBEprDUkSe23Z+T+AlWLabZMerwvDlz1NE45/w9ghhhznwsWglD481
CkYU4PTDHN/M1PfDE8Yil+4CYNefbFhYfmyuTIMDPBlbKgfVe9W0S6QWDhfj
3qy1csnBNMlE9VPXI++M3w16j5s9i5X6h8F/X198BVn9Pg4gdxtmH6MYlxzP
iLpN7tZWm/x7PE9vLA4EdshuHULoxCyJ7eju9QM7oxdvEz4FcWCy5DDieG1k
qrYFG/VNqjS6DQGQgHWFvEVaWwrGJA01795tuAdpSuAm6nAYCNFpTm/tvkHT
3SgzKLldygiibRZMEMdebwJj/XuIQFz+SetTCOFBXCWW7bSbmlJfGwBTT7Vv
pcfyZ4zYDTQGpq47vIgs3gJ/dz798hiSol72hEWGanaKeMTVUFno7R6CM0ZJ
5w0VP8JajgV/1GriTO0vIHd5aW8rvUA4EXmImSabwK4hdpBbQ8R73JGeQdJ6
wKPui/1sQFAqmbRE16Lmk6EmAjOwLNV6+4i3YbznJSn9D8L+mJABqJ0RE6a8
leGB9T+hrGDcm+oIY9YmIT2htDWjQQ8fcEXaLFVMv9E1zM0/XktH9ChpQIxh
yc0ATjIU28DJKXDV5D5osPRWAV2bs33TXB6XaOGvcHhUmgVL+QaTSuWoEkA5
eacQ5WoHyy7awf8TlF0UxKpUpreUxBjE1bgkpJVURtT02FC6mPAN8uSLjnXL
8hXf/azkfN2OSKgpMxqLlcXzg88uB5kxNHobOPYeb762BY9+lQQw1R37aR0k
xuSb03EuSZQ9BfhajqiT5lAz1/VviMOZnZHK0R8lWE7Wq9jbJC0dwVMDwNvw
sueL5KcipxxSqUQREgGiLUuZGep4cDNdQ4T4u3ZxXrOrhDb7mIqHAeFutYAf
tLdTnlwDZmMqC2foI9/VDZO3HqHrZkfx27Qkh9zIEjXueUMk4/TnZ08KeYmm
rf4U0d/bM//yOkjtvdsiSNTsLKc+3nFIOaF6UXu+HhgBA1I8P8M1nht8hiRg
bos1kfqD2+/YJcrWSvpwi1tW8tkF3kyR/aEQHuAmrUc3YPgFb3OP/sf8Lbu8
MzzYgaZW3vsfHcl+s5+VtYsuhpwqRHp740rRNZOInvZwm+N3bubowAN2dMU9
EF6diXX03QsnRz/K0uHmMj5hpiej+d2pHOn07WSR4g1o7JEHcBFC+/VL8TQV
2J0D2KI0oQIFXNswCXJNDib9z7mueXvfaFClIAyiJabcWOlDD14Awm/ZZbSF
6JiBdIRuIHUe2lnBeJWf4vUPli32GKrCeTC/ZrgYOFbqGgHKlujIZ3AGjBbJ
xykJFEasA8CzIc0Rx5+D4AH+59XaaMnfGV3t+sjNAzVjKXB7JDlaXnWYKlVj
SuQKFCCzmfpiEm+QNjfirIh9xu9dW5mxF4/h7aeNn7tx3PZnr75AhLBC+PIM
Ae8rIkV04rX6AFUccikfxnaKx3LGTRoJtkGJJV2t9F1V9LODpyU1ypOsDM/7
hVjVoSt4uT6DUhZDl6n5RV57bEyayRXohVMcPtRwgFr7YuEQHII6iMb57Gnr
JO5a6yJrkl86D/S4cQ4B6nyCuJKXXCYEmBd+/7sIizZqswr+JlhcU87Jl67s
xle5gxm8ks3tjnYiCMdbrwdXbdmh4l427S+9B8jmDK6phHOgiPQa7O7XqqK5
UTczHh3o32KeTjSx5ln0UXTSP0nml2axLlOS6g6V3M4qWEkdTkkR+JtLvb2B
ZckjNtxSGQI46n+eXiI6PHMmx6sZcrpJ3sPoJlUBhPu3e+LyAeLyNB40gsKd
ttNG4bsB3riNXnQkQHA5vhxGPmAl8YpEETpfM/Pf7iSRM4qaG/yRX6C2yp4f
JFvxTux0Wyr9rRMpFX7o0rsEitV0EKsH16ZNo5L0KQosbRUXN/YWZOV3yEme
3A0tR24CJ7oOnOyd5NSIqSloR50bqh8KzldXAxYCQREowIdnehh6jt/mUTuL
q6pkd1yVEBXyCp+Bd5rUJPCNDP3yI+u2qONNebyMgKM+BYj8pi3SDokO1JvP
YQei4fELLvKUN7jPK1XkXErF9sKOnVo6+Hd13gRXv9U6OqVfx7vvoItHhkgj
oTHUUNUi/hw+Jfpjek3csXPeV726dkOUNhd+sNrvyw/HHi8L/QMiX8DfLrZv
G7NrQavXZLfmtRifpli3iX140pynMSmche534pdMC+shu/bHGJOJpAF7VQlV
Hc/8OjD7BcTil1Z8ig9w8DgdidXJzx1szQGQn/0FSLiBeSVr8wvnRlFLX0aP
G831hiriLnmWtB9MOutCwUJrZV9knvnEB+Qv4csTuIZWkw0kqEfyGi/4rYE8
KdmLpKw7oj6Xs4lBGa5JdpJJEqGfx9iZx1+tIbESB1FbM7suiSSo2xP4C9sT
xiJfHjNHqXEjnWciNkr8PYTKNVP9dQ87TmGE25maCeuTIcXIgi6SfBLgF1AI
tGqKVDpzEG6FrGUmOywvFbI1MnThZeV6coWSivU9S1iKYenXEd/MtUlY4uqn
I0/H1yIw6luvU1L7bakqTjc6+qfdLDTs6B9Zh5EiAN1F657tLU0qJWnqvEWD
/FPOmIc40pUnnXuWZkJNroAcenMBaWO35GTZ0K81WXyercJRAvSWmN3+BPE2
EzFQg2wgaHBA4XrTV+usIIh/lNMtB0wy1hnW476nbHUaL3K4akYQ1b2/VJYx
qG8SNIUi9YyR41dSkvC1B2DVqkgTZfMFZgwCVFfEGu5AFENM2IqN3xqrOVtU
oCAFzQ4V/jxz7sCW6nitI5q+wV0t7Y8ozvqoNsM7mwO3eKWIWGBOLrw1x5fj
NygVi38ZsbYSwDhL+EPU+hjxDAPxF3r9zjc8hbVXTOyAmOr+JXBhdr8MwH6w
yyejJtcHxgRqVKErsQadGW7DbAynpX1iUMAv38k4t/2QH1+CMt+7Nbe8SkOr
ZsfXZAcvR5piUrnfMt60/kZRQa0ZpNqBBNVNQwivcGhnjMg0SQBNRapHhaeM
qdRaj6yJrasPdZD61KPYjMDcInN+ibtBo4y8w0lNq+PvOBRpL4U2RSuvqesB
1cfjc8oPJ3HC0AcurYvsl12Ix1ObYKqU4CgxkucBlsC8M3X6N03cdQ3Bz5Zo
wdK7T6Gu1fRURGII1kpfys1SiOvMMVsvXIWyHuuXxkLoGh9n474pinwRytO6
iv9cn4rBdDdtEfAW6h9wqjohefvuvtJ67SpXHbYSJjMtAfJtMz2ZwgDkP5dU
QivPDOdEYQ7KR2Rzy9X9hsttm+7aJ+Rm4V/v/CYAt9+o/dwJYM9HnhkGJ2iG
HQWqNLJxYJrDrQMlTuAQISGZfkBRZe8U8DYGLCcq9LUs4FFENvhHjeBleXLe
wAjjxuKr2CHVH3BgWlE8xMSiMUMYP6qwqLPXVQe4BuPMEZFld0vyeii0hybD
HjtholOAZa7i4Hil1Tieq3AYfrneBkuXUiVi8kMqbpPT2GRYm/U+4Xu0ATa3
bZofyNyFC96diJru6DYQj3cEj3otx9fBx96L5kNxvRxi4yECKgFs4Xw8Y7A/
+34Ihi+uqAXZ8Jdlfd7asRU2jGz2tXiZRoKYJqI4NCKhjtfLLru8P/eExYRw
iH9B2i1F1YS9buDQBYm+DBAhXJg36Y43z+UZH11Ng8iGTf9xWVjyJE/ShRhV
/mUpsG9LCKb0qa3bOSF2haPcy+G2t7mNOLuSltDh9oZsz649OYFFrHOlhzjC
0W+9ahUr0jJ3Saf1PLIoyKrQHtv0BLyVjvvHoK0PiH+f5iSu9hv3LG6zpn/w
5RKela+zYXhi0MsAp6ykyT9u6GMvBt4Qs3Eb5+4nq01UkzoYKBaLqY8KLf5Q
B1cG+kOQcCgRy4CEoob+HWW3ZGYInrIhwH7VUXQfZKnq43+PyJaryOcYc0jk
DaE6ta04jgDhkLQ9ySRVgHhhk92AjKuAv3VpgoWDSTYn0mK3HsfDUWYEkkwT
a8EFnbdmrY6gFR5A5rDFDiELaf7uIdSAjoGxSGRBTkXEE6my78Ku/rcehUcT
itPzh+0lnpXBZ1xhjy0TkxFB9jPsHRMxeRp4SQMW6ftkz1baP3VM7KYm9b7T
JkwHDIv/PuEwVcnW22TCabI+tKAfB6cl+oH4v/CFKI0rRwlyqbK5BQlIiwxf
5Lg64d3WWJWEcUTvzrTmbhA3bP/w4gEqOBcSKIWeNcJzUYTca0Pc32zcMowY
jLo+e5guzacX7y/nf84QacSOrq6idSITvpRkrVzSqVzlBMnqDezGglU8Ik3/
9L65l+LQelags9U5zyFshmJL/9lJMARvcu2M3tSMepME6wRLA2xJLbWFmPi/
MQJ4oupQNNHEUbEb3eMR+cffZRDvMDNns32XSad2sLhnzJHTMSGtIYWrgnjq
8ppmsDYUYPnY0jz77Orr5H0ys7CBAHQInzvERQ2Ncl+iP7ELTtV/sb3znKqB
Tqf+7qrHGazEXCqOSlGR8gQxNee66KPt8Z5hJyQiGI/1IcvprknQ2o/YytQE
OvuGGSxXfrzAOnZ4ykOmfoIPpCjj/k/fXoqTvLCMIfATVUsgRiNyxaNgE/S3
kHTuuhNJJi7S01CmGmpzjIVOC75eM4K17pFF44n6qYqzdz+r3yp3EpGeVuQK
hUpRbVuafkJ9k0jDWxXT6HrU5CKcWf2VYXxSKKc4aYE2Jx+pKmRnG3u7EtjN
IeFj3mziT66JlhoOQUsK4vAomFs58Swkstb+0fevbigSfq0h8HufNeU+rgSA
VgLWkamRd1/qj1lxWtM2xd3wSZjg3bAStnlWXR5Ojck6v8Ch8KiHAP4HDnBS
B4PAFmwbC6MyjASn4UnaTwUaobEhRd1X6b/QhA6elJ9ppTKQG+ZIDU8JQ1PK
Ghs/3HzWi4kqXpLo84Wt8+G9M/gFyMcJqc4W/Xt9pUm5t5A329S1b7frbc/U
HSVIZu2GViPHDDds1Fkr0TDEukjO7nuxbRszMtRamLTS6h4inFM/+2X0+Hpc
s9wKebDGamWUm6dtajdw87hGDX01jU+aNzDVgIVRRJ/RXoEY7mUrABG+zpWS
gTLypPg4587TNf3rir3NOvfrXrsBPTny7a/D4/A3KxHMV2qHumAdXT2G76wv
1c+ElMjYCQmvokdIfTtbna4gFCrNifQbMNqTWaCFwGwYe4sRka9dnOW9Lzab
2gDQLLOfnSPpiD98I+en8pCA3OKzr5m1xsOW5X2QXmirxD+nj1+LGhn1WwQZ
X6JZLjDnuxJrodFAQ+KfSOEqmiI6T4JIvS9wGgA8aQsSip67CUrUrF2YG8HS
SKrVVGHxwNpn/9HO3F1JVTyWlvtk5dOWq+ygJ6zap7oYayqzCNgGguAE3Ua7
RhmBGjl3q/6gtQT3RF7MOjaNDDYas+gfiK1NIPUVgPZaAWpHVt+NM0qKQBuX
i0qqxz2qdE+Q8oMnnK+msqiCCo/gl5kw04HnCelVkPI+Lbrds0l2PSqHHsfg
5RnFizArms6p0ly2ppiKzZBO53wbhsPRC7PxvWE0GmsKu7/Mzleoe8MRM7Bf
DPMEkt/TLZb11io+EosEjtSR4AWw89Y0n5GZ4HlAjOIanKhsLN8xP89jGeRA
KsL1XNsh59/1Xblu8lgdsW7Sd+uuFuISBiN7kXeknsVXDIBjL7bwjiBGLXFX
nsh+gNTN4a2Jk57F6tNW2svwv6Lmma3hhWRLBXhGUGzVgTCz58jJR78q/esk
dXqSudMtuLFEFP6bmsreZRP+LMvG0a3GkAe27QOrPaKIeyEFGSNsYt3e6rst
WdWuzb/LtelKOOiY2PkSLLPWNdE6SO/eN6xmqd4R8uI9oIWXgdrQ890dtPGz
8fkoJ5L5WM5wO92rjBcAxw7ecif6AZIu7cW02qRvG+IsZkaN4/J7awuweAv3
hGkByAyuM4mhpu5PCkr2RBv2idszYOhN4U1f5AcwH/1s5Ynq03BjWvWAXfvL
TIJj+7XKBiFsjx3XnYO63kcZqVtAtpDniqy2sbigHcHb3MHYCXSFmo5QVDli
/dXeZXdw4Edfr47izFgmlzHV8QJiAaW7XvNgJQ7ePg55XZeejdd6SRtw+wLH
6QjzxmcUxT2zfTY7Et/T5kANB1mzk6JRLa/fCFl+QTs+twJNAbDbsh5feDcF
jn7sDxCyfsluOTRiJQhFQEn65HDLZetw79V/A9K7g8IFBVt3G2+3roQqRHm9
9XUkqo4bLfVA5KZ8o9wQVo7ZPNAEwDAJVeD3tnjgvR96DftI3BH/qT128cPS
mINxjr0ykydCeckzTs15dhXoJQP31p7QwMS6N3VXA7RwkQ/GgaopxD4th2cw
3jGMnSKbhjzaEPDPhmseskZbGR95WCNt2+EmO3m0OQcb1y7o08X7NAs0l5e0
RkYvN6bPd8Ov4XC1NoMCdaGQ+CU3Akg/FNnJvrHlNZrrp/ZJZeQ9P32DhxT8
xBUaVD0j+kGYZgRAJZezmSYCkvkVfTJa8z0VJNHERZy1TCOivllCm8/cLXBg
kAaWGPZpCN+yMT97S4YsBobWEc/gNNM+WAu84L+i1xkVCjwys03iHN3bEdgk
jyVp6pxAmNMeStN3s0PZhcGmfitV3SZvh1Np2IdgCuBsNZPMLJMjxgFth/W7
WR8UqBhQ40QwujHN3Q0FxjBxjiTayXcttx1fUo+G+8IYQKhH3ElAKFxDIJoN
FMgoYbpvyHAqS4b7lcXtWFbFTlYegBWbsFM6lacXsjHy4KhKMfQjfYKrKldM
GZDh7aokNO7hi7zy8+UQiWE/1YiLt8rhf2RF0mHuII13PbPT06Sdm2VglC+s
+75IkGp3RB2xhaKvKC2J62pPbEQlQl0MTL6PUaBn99HhbIczof8cGVCVhciq
rnAXRj1rv6ByoUk4S8FNB8xS9dxeOz3OpkxUtlzbWAhYNjTPaHyQhtMheoq4
YhwIKYL0jiFcOfOf+ul9RBFbh41GnoD6vMAca44EaTf32ZFwz/FB5nc9qUFh
kNh+hKKPbXB+AK9vqjeXGXcNptECjUcldxnZblAFS9t4D7u221ygp7hfkwcL
kvW5ngwegL4MW3E9B+PS+U4zUD2d60AzbL9NPSRfNBI0aGbj7Uc1IC1suisY
2x2/63dzto/DLUIOVv4R3lbRY81qlJDQuDPM9cAjyx4epaVwFCoU5wA1iqb5
AaaNpEbVrRdx8QXdcKBSfsve2FtI4ivq4rT4RxCvtHov3vUs0N0U5gBTHIU0
7fMFNr0vxg+HDnk0OiOPqZvJNovgzycZFVLc098gCXnlhGFdyyHW3HFrd05g
9M5fDQ3WJcAtDDBhqfKyjDWDy+fm89gn962Kw/xbkD3Y0WZiqXKKogwu9uSG
X6swRqG5q3Jqk2XehRCi7brhz8Ro5WitZiKA5SSZ/vXCsKHsqt8hB5PpikVB
qAOZkK6R18FigWr7td/G7nUC96MU4kLHNC6pFeMC+j5e6cCJsxfkbNCM4ic9
lvAh7TZcc94emm0IclVWXPaMm3xJPVGdM18HuR76a+sQT63EJNwwgsaEfVU6
yv+UaEqlW0TonNbkPGxgsNpDBNwXZeFGdCxEfZKo8vOiRPgfiB/9oy3xvfZK
Z/YY4JhHeRMaPLWUe+ZjsktlKjH6hs09PczSbls8XxLDmj4wM1Z75yTxCeyR
V4CXlJfSHKIVVa+2DoqKs1d32eFzNkWYmWbrNzKpSaDcq1e9Vj8n6/bdSV4n
lmjtXst6LcGxhPgZGS0H6zihexGi/3LlzvW8QDMAHH4TMtiDNjhSAXBWdb5F
0PGezhoG1IJHo22AkkGCFJ90cxtntS0Cd2IJkBrLmgFyRGj75oQn4p9KGavv
Fxa5FnKGr+D141YlpskKcIbYQZ1YQLWIIkwAqo4/RIw6HFfhDc1heljrD2gH
QNmJpNSODKxIBb6Q61PnMb9IIzDKNZp4ABXY249L6W/v8Ibr7+a3JBHnbFDT
2mbOloMmPScGpv9f8j+iKOlun5nBXnQn2QNnjxBkp7zxGTAkfwHqiADxqcNk
HkOu+/gz2TZZjd5xhuStIUnAWrtKYCAOzfaZLL6WFI73748NfyTThyK5GRtJ
nHkmHy1MW+dpy/K00Qk588KDuNlkP87bnZA7g3qlWuYLdY3AXVUv0YI3DsDZ
HFlRiCqZnXYWLq/zFBs7UEsACNQRPAQxP7Vum6ioReUVVZK2k7B/fJ9rg1pG
iqMV0Y2ME7qH3CgaHmXCBsDtfPwHqPbN+dW2kRaXTFks7A8LvcgYDx6olSf4
Y/SlwyFXadKxFmIxO29w4PBf94eSMOugySV/A6MPlRJKbHZ++cKHT7boHQKR
FHAOUmyeoKOVM90YbCqvDYnxHiviFijneIqHEWh/UMUdQfDFlpGZCi23d9VR
i6R+d9MvDD8/pMXyQYAS/O66ANAiJZKfwW5Kh+hJ+jIPZ/Fq3WPyBx/SwFb8
SQRd4rh6LmNl/6s5KyrqbBcfrxo5eLi9xjMaRG6SNmb+9LwoLKfdwOTQiZ1t
ZGhWovydv3l6kuTLbnJN/we7jWQNU6rgr06UpYo+UwL/qc5w6/O0rCsfKzh+
A8a8SF3b4DkMRr8rrBCnGPPIAGl9vHeN+r/YOZ4LrQj+uO8oG/ezuR1okhtm
OLJTgEnP3HUst5sKmghFw2YBA2buYQSbVxm2fVQRJgYQXwozTGYJNbUChvtC
R3Zj4thzxAReVIsR1xGD9tuiIJN7QQ8laapxrdesYGnhkf6vPpWNpsLexCwF
TvwNI/wDN2lw2DoURrUqGQ0a/En16iHsD2+dEQn597gX5TjRgTYbi+8noXx1
3+6W6HsnJWEj/BVL3k2ZeDim2peVYygZJioBOtKgfN7hMYhZdGMPx95D9hKt
zfwC1qK+l7TLdITbbjknmps/uxNhB/2GSpsflZODl+1Fa3WFYbsAS+ozX2zR
J+o7vnL4rbaZ9vnie5GHFnxrVhDv6eWuWZJY6SY94300LoC7KA1k9dMgot/j
Vag6bMuIu8/ue+FW9LdYNmmBpJZlwjUD+VG2nnAKSSuagQBT5K/36AOFVBNH
mkAhINlyoYCOZQLM7u0QI4XUogcp/jr+y8Gd9dwJUDiJvLmru/xzc0KQxqAl
nzB29RSdDnVvIL2+d0+6symAUOMv2mmByJvWCopjC/JY3UB4reDX4NTjsfsa
fKnxG32v9oQ4vSaZsaXcnwPlXVzfNJ+OHJw0Tg/ch/5P7aJvueNMg1dfnPB/
goNwp1BnfrdxLE3FP2HpbBZutG1xz8liocmy0kIOAxNwglYbHXqYvFlri4ld
uvNis5hMf5u+JgNEDR6qurYyCTsxDegFRHZPzPy8jelA9JEIJV0/XNm4YQwj
EIvKwM+SUCWICtRLisjFWXlMB0E/2XgtVwCuLVoA0cQRs//ZdZtSJS5iZIQm
FeuC+ZWQNHK7byXfnbZxC06HJDxC2YxS+P7ZsuDJpoX1weP7PQyPduKw5oLs
lv1v8xLy2p0k3YVG3oAKQ0nieZuwjGSNprzsiU6HSb9RN2AWYaJYhMaHetsv
qh8Ma0bIRZB5NqjZU3cIU/fL37z03HoVKbBSIZ6TnJhSww41vlg5/MhbIeJ2
0bxmGDvPvn6LLmRVL7xput+dFibsuv7xeHbIDtFzbXvKfc2z07TKj2tzSB5n
UVbysCWDSZooj6+gnchkHmj6qCKgzC4sa+MLzAcWWZKE3bqW+8NT6U9awt8p
1jP3FsoddIPUf/joSXcV43Dx6PP9+7Et/FNvUFNBo2/OmGtkvrdPjybUN2g5
mD7tRpMIBPeOoGcpHKgCM/aAc/af4hMgriulNNnxugdYfFb3iCrx1VSZrD1R
dQVHd6py+o1sITIrkD2rewlauZGO9nSS9d3Ij/xekgKpN6IRcjfUynprRvuv
5CBPvhy838Z1LiWt1yfS59r30IUTjrRtnDsqMi9rDVEgRw3iif2Q/5qbHrRu
3clCTDrfk3/CjUHMWuDhmiKMPiERPZrFvS5mG3kRt76IO3GsogVGN5/B4lUy
4v3ru9JSdmuz0L859d9VLIn14GjOBTjGGyUwxbS9ktjnC98cClmmlKwLDhYf
oUAu4UHivqcstzZeTAKxvQjHi5yl5AkqF2lo5GVKtVatlbR3z1u6kvaNWin9
fFfdRT654hWnW/gwlto7ci1SWK6v6PAaO2A2TUj0xHhH3JLAHWBNDxkeuQYe
QLU/xM1K68K92nlFZBoc4ZBg4Xzc0Lb6i7jLpvxn2hm+gu1o5MZgrY1GfGFJ
ypHS8g3x8s2LVlbTQ4msp5GQKnOrEamm9e6smZK8AsNF0s9Etd2nQCJTfOSp
xQs/Yhgf8cTKPjJcyeBmFzZzkNxqnjHHFMeFwB9u+P4iTeAm7QAf+DXBNEXT
Bo0PzsG6G7n7Ab4vsdLD4SGotKa0qES9pjaDHHCeMTA7dH/5+ckcl9we0sa2
DhhrBdge52bqsKG6lFBADPdMlIVQ/x2co7HR6n3jRM5wlTlCm+h64tlUGXGX
PBNafUSMK4nGVe8pb489h/EKe3xPqe5gkHUZP9rGwUiHeLJvlqFAcvH3gxCG
8bREwN3nEBIHaYWT+8LJpv+KXHkBeisf7ZdzL2Xfd395Z1OnD3HV1uEtvmgy
ZvjTAxIbuSWmT/JeuirlfsSJJU8+Nycf1anLp0tKDICL5OKurdhn8Nb7RCQz
Sakc6aQAa4ZO9Hz7CPJTUh/iTMTDlz8U5aDG0pd6K6ab76y8sB0G2aw2r2L2
637IBPLwqDvTg/z0aZSr79iINjz1XXr4WhQMvO+d2Ac+54jfiwMBb89iGMNA
TyPlsVVTrN3ThmmnAB70TDaZw2SuShB4Obx3GbTtj5z5+Hg61vmFY3al08j7
Fe9VBqXZZL0Ov2iHnOCouBCfgKUOrOG+hUFAGr5OvbRKv42FSmepAYxlzw0F
ZEQ7rmY0uAxVxx0BDnxvt0QDxpiQMDXtIyNi63DScoyTCKvH4jp00rsmUdH4
jNrd6kPcAGphAbAyIPpxUvXiDSSb6FzjoPk/5ZaINkZcLNjNfyaxMRcXVdTT
aIfqRcAZLh8BEosCPbNxR0Sj7ukF+9pr+RdeNT7fKAyOQPAyGa/zUzrxc694
2lZ0IY38B2VUJSAouj14bKeaS7SaVWE1q3BerzCOmmQHl84IHoZiiXQ/j9D/
AHsu58u1+8kfe3/JKjGDyfTj3T2SNMHMRVE6DH8xCNzLjVxo5tJ4S3j6fIWd
ZDqXEZqnzbgvo8/S4+/lmWDDVfSFkNR78Nvxh9u1s0CD/a5QOLoX0SkQgu4r
tWds1pTGUSZLkAh7SRDTahxTy4dtgcVF6/fi3zDx7yB3mnLgJzRfem7Zuc8Z
fAViV4Iysbk21xnVqbSUVyjQZeNwvt8Z0LpRz3heE8iI198iyTemUtQ2C2DT
Cp8Qquz4LtUJjOXuBy86SqBDFXfrU6v+JG3D/deNBr73hRAbVZezDAOzErEE
AD4Xg9Tk5yJ8EHG6Cax/T4R0GYKe277IwPGEdO14gZ9j4lRNAnsl44ACb0kn
jgiQndCL2O1HTI1miAEfY22xl9/M0teS3TdM5qehJOKuPpAVuM+RpB2HWlfG
uKo+63rXKxnoKY9wU7bDhcI/Fud8o8ZuN3NcplnCy/+5qa7wKjqMmcfK+xKs
emr4kZ7313Rt41kijLnBKm33OTGRfmf7hAOLECC32x/hlvHcJuSd8TkVXXi/
E+NFNp4KvDnIkUm4/6+GkpHF3KJ/fD0/nu3nmI3gysDdBMV631BiTcywDCIX
wlp0ZuBtAnKN+OKUjNYje8pQ1k8Z7Ku4pSYjA4JUup6DOulRDq/2HtDQFLG1
GYXOcDALr3xBiyQ3X52P7s6h0DieK7qvsb4PT4lzK7Uz+/rztoWrd25c+ia/
ECQNqviwqfx0YgKasyGtGIif9UX0uLhCJRq0IhtQ0yTOOozQQO1igClVWBjD
YnmJ0gxGkY+EyeSq4fW3vCoHpPH23pO5h6hv2ey33dbaTbyavgcXK6+MMwZr
0hZW1e0eAb3IxbsNW5IFxoeZX198bfniJO5xA+IeJ7r1IlvjhgUj7VV8BFkC
oRERsCyztWN1j9E8P/HkWX7HkNljarVhy8KRM7FZHOAZ4zyrfAOKm/OgD15Y
GYLX7XpNPZzTvibRDvVgU8bBZrg6T0n3jpDL/FKE+dTNuzpd6Le/37fJQ/3g
d5WfgsFv0Ir9RcK9oQLNIYLnQMoKD2r5qYvdE1NFsBxF+2xFKIbgWIuGYxjD
dqxUWSy46Ar04iF8g3lAJN0oOCNpntCxJeyv82C95n0eVkxdQyT5ezuBX7dZ
L3j3fDdxEc8DjQ5R2OFkKmq7AT4y7nzDrJVvksmLS+zRsHcnOahutQ5Q3e+T
FYs6oE5VGvYItj52b4FJfQH35hsyP48WHM9Zg+Dz/7+I93fw/8hTlKoERtgq
dtuZhiNIldEjs8zWpY2ABAOT+mc2aAQRkmS1uHXmbxBDIvhWm6a8t16SW2Fi
h3hWaGSZKHXKsfSYdQssoHt3l9jDAhHF6oPg4xS0BXUwEBGwqJD+5oZgOekG
/85AFBbetzXZIiO3kmU2CP1uhyn6maBjG1z6AzePYaTg2g+l/ZehjruQ1I4j
t8VjZ4UntAYUwf7c4S5dJ2djVSYpwne9bdYRe4C6hlD3Fqg8ykERuTu9GQPy
SMYAl90EilSfDGQJm3N8bRQcBtvjnjDqCWljfXq4hlUGHo+aUJit623y6DQd
PBu0qaDloRCR0PHq0JFeDstPwtANQmkESphomaNosfVrjbCYFUEM75M82OyF
3MQxhvxuymSCMYM6QTi/SePaymnC8qxT5s+HlQx9eWh7SXTQH0ZwaDKyO/Bb
Is3vfgTbkJcjPFKAnij1HSesAH0ItXQQAEVd2hv5HMy58/0IeAkgGOkIUGci
7Q/H2FiQuEPlmHE1YlAQZ+FzPzK6nT5cIWyQOI8Ido1GpbVWvUOP4D1KvFE/
/n87ZIBjXC9pPu/aBq0Dvd5q0FvvaTby5SQ2639lr0ucGEjiBobSGTC3Qhly
Vqbj3rbtuQbt1pM6RLMAnXwKKvOFMz5hBHSYDsXW4+6UWlWW2GHKPFSZjwC5
6kHO5XYLQ/HwTjT8S47CqZqSq5nfDSNKG1IclnD2qOdES1s2GzB0ZOFlS6XP
hImKyJHsMdB1VHlQ/EEcjPD4+ISRf2AUefech8A2Wkvupm9PTUkJZrr4dWDd
LE+Mahh3qcfWINbHpkBH29pGiVXCGgHjmV6mxtQCBhAQIJ2zfS4x13FSQXWh
YenEtcfRi7gDEtFgcfiNZnjP9tBy+H8y6/U5KgU7nAOCeg8r6sgqD6xWwtHu
gSZuieNEMs7ByJh1f1eUaTM5hWvxE3TzJBnL3eGB1OxKkebneSz0oDY7GwcD
KaDA+4MSSGed2wG+VoYjRIlkWne3yw3wMVLZpM6VU0CK7sLS4mTjLSgzp8W/
DAO8QbNhfABQ10gyz7RobgpSvDJtNbgHu6icxBRYI6avD6PA8IWNiJZAfpfi
bD2Ec6gWe4d7YSdA/TSxn8pVtahiKONB8Tjr0dOsBMf4bGiW/6kEqZDxFIbC
O9DaJ6PMMBTCsWCNnj06ENtG9WEHc6xXE0zkWWu6GRaRIFams5LfRBTaacAJ
WuSuZVj72Jai+bNpAP+E64G3rw9ftSQaSewV9OTUjey1RmiYQGRltGg3hiLk
+E81UyDeohAVgnoBddw2dCISHrUQ880PFTRdw1O4SbsgqkVpNy8Pyg6r8K2T
wg1iTaBE8Lrg6W8v5GOLySYAt9FEdyYqC1QUrBQLwz5sb1dgQaG/1o8mCvU+
MTx9pi9S5zEQo6EhJMLUW19Wjc+86unOdf150qp3mjnas7dBrMN9p8QmHnaX
OOLETw5VppUp9y0FKym6f5AalyxhG7ae5/X1uERujD8G0TIApON38kinau7p
c15Na276a5/VxNIcXJ/7H/i0iCae3mxltrhJkqiWvWklhbup5T9qf844AgGe
7uPrZD8JCzaPLcyVf5bylXZV8U66lt5uVa80gLcGkQWdJT61udGJ0kdhbsUp
kzNNbYTUmim5MAL3onYGWOpdq6f/Se1meJa+RyIqtQjg1p3Vb7dmn22DSg+U
ZqTXsjnTZZJH2k2pRRaA0KLfwj/siH4XJqRzDhvJBRStL4amdItVDR2DsQ+E
xbZ5z06nTayW44QvBxGiZmEdu3P6OWWSgAGOmJCpArQWPcPYcaxmoptrTL4b
HpvjZG/VhdZktRuKy840pfW4Le866HqGBMobftx/meinlat18Ha1mXyatYgn
KsQdiYXlJAS7CEuIjmxs6ViO+0gVjv3PRS8eN46uO6s+N4P/H9QnnUGwlegc
amL5DWj99ZxuJlVo2feA1SompTSI+MO6KpzXijv2+0OeCuQO4dVnwnWY+TBg
8PjBJFhtfmgdY91pB9Oii/lyxdsxDqjdvMbFZfZTtJ/qj1huhubN0at+ID2H
pGewzAhHqkst0F4py/Ato901i2tosLg3eeZMX4sjI2RjZUOHT8c7mP3V89Sl
rxYZWdIPPgVJ15nXVcXARd07H7i4BK4Y8a7fad1cIdLVYTgYM349OxCUuSxG
vxGbXI2seEUF5nIUZ56epJFCt2rNv5DXyRI7yggTZp3CDU0oVTnF9Zqd1VMl
NNygwS0sam/G5XlGIJkfOCqWdDyoX+FxPKayxwktKN58v8sPkNtHHfBaFZWt
8g2F9+I+Ig9/oGeq4TsFT38coCX5QOyB6fcO9u2phdRJIxGnqwcMvTQ0ZLpn
HDC8l5YCT1nB6zQeQZYMrCnTGl4xKdR780GwH4qIJj9hKsqONppCih3b9Nye
eTh+svHHxx0esda5mB677ezKq/IEnPNG3f0kZc9Gwmto2K1ZpgQECC7JNCjd
9E8l+IhEcaD62cuon+eCAyUTLpejgzN1lMvwllCeUxM7bMFQj29fw6SYUqj9
eozal4ZOoQ1AqsWWcZSgJHpjLWUDtLDMm1jADHdBMtPzUz+SwjfW+HHO9/Ls
NL8RzApd487x1t3E/LUIZCxnnm4uFm9LDh4CDlwVNFyN0dGj9fjKouRoriDS
JU49ZRCWx+u/2LfJ9r0MIPUxZ6SM7/pKUuYYJNtwFFcmJVV0bfL1I7WTGe0A
Jf8RZbQ5xga14RuOMBPskl85dykvPes/98iVvjfeqkkUguuBPmRj0M2yIkFz
pRU4PnQxmh+Cp0yVl/AVVehiOX1xtzvucGe1YXQ6y1Qk/atZsQRhw51vSPKD
b6qvOibSAVm0W/wknYhE/Y2IqXyWmMrFCCD0zlhYWsNOb6di3NUo0p4wXg8Y
LXuhD5OS3IcdCDl+t315VE7F9i+5NqljMN3Qi9QbI9YzZyGM/nxnRisKsW9Z
yj9JeUO/8hNe3QjJANpHBCd93hKYRc5g3MWT7KYPHRx7wM0Du++gqfYDiT2W
i6rBStOU+tnsdxDowGGIE4ReSZ4f7vRNrgQa0JGdTA1Ft3pBlRp2nOxvu0SK
FRO03i6dXa/k0/5+hrFs5hRfGzCfX2fxN726E1viSDiSpUexWhI9whLi07RU
AGG3nHdhfGBdNT3DLZw/L9g2Xj431VE1+ECMKQsEKeT7aAAueOWt939G0Hod
0276/7p2nhYS9hEu8owS5OiNDMoKj34X/CEfOsZfpxC4OL6LUndj8utSawOY
iOdydwyBbiuagsXDaJZZP48OxLPdEDam0r8y8ND0G2DCJfvzcutjRyAshmVR
RjnQCX8jrIKyI9H9ma5T29SxD9fFnMC3OCe83S9Hlq83+CUX+lZ/apLXYE+O
zHVoaRg+C0Dvigjx03oi7nIDvIrw/uJ13p44kHgAPz6VTKgHxd7o4ZX9Qi/q
oKhUKZTsPl1dHbA2mDv0vjApQ4Hbf+fH97hJ9fMs4Tbl8jK5pDSvZ3k6yEqf
Bla5lmzCGbzHIcCdXAEzEIIXsLnZVVaxvlPmgrClzela0GmofFBQNcLmznrH
Q90VHPTfmuwx/O33QZZk4oQgw69BJ2A12JxbeV22A9FbpsuZyjoulhRXSPSK
ZSCz0B0ZQK6JkZEThfJFZ5OLfsLRAoCPAWkWf1Q+/6U8y4j9gOSEp6in2/kP
cAbC2ZZNfW1OaiKXA+OjQlqpZlRXjHNGLitY1VTV8SnLsJwbNIxmJklJ2seF
1KIAzIsxJe0UIxHin3TlPBvF1ZxGorQmTegLyWL6jgbyt1Pxcc/jVeCwSgjM
XRhBBfiJsAA2gW98M4hwDq3rdo+Vl7nHWa6uhdUFFoTVT1sz2GA8jdl/8VZB
0FkciNh1F5oHLjaYvO4h07IlX2gMvuPN47WC0It4/+b5F4a1W2HQS7sLuNwM
hHhfxXMP00y5UrzSGVtOe0ZaJxzN3Fvs90HnzzsoR4skfryHjCe8S/2jnRrS
faSIiZXFe4le9PjU+WDZc4C/S1gtyKR6K8KcSdV5szbOeqUsE9nlYY1biXGq
d+5D9mxMrQbjc/fKOf9mTZy5ePzEm1gqziBSySo15Ihii5G04o3t3hg13Nj6
AO7PSiFpHWqA2+ZEDCU5zTPcZojAt3nU+7psYdiJPQAwUaferZic1+HOulx/
ueC0HSFE9qLHiiyTsEgsr1YvAFQbUUk3J6gKostve3gwVRzNUdr4xKy3pv5F
oWkhDENF7wx0UwNQbuSkGuGvAZIDzbYJMz06wPb6ZxynHcuT5sQMogg5BaHf
QG35QgFGn3pdRHlHOP3ges/MmDiNyJiDXiRD5S5PqtQWac1kB109f8XBsGu/
PdTy8vIdJG0xF7oOp/rcu8Ajdj83mwmwPegmstLoPGtdf6KHAMNMowKzMCs0
q5qmg9y3goKtihuC2fnR4LPl6ZvHKa1Y+FY1b3usf9G2I8Iv2zTaaEQJ8kSQ
QT3o9tJZhK41Xp7nKKC6nOp14N5pmAvOPkyfRZrhEZFiCYeK8wZZb0e8GM69
eB+kfW+67EDxCExK14BJHfKG0piMMb0Qu9agEs8FgApA3fkqDdyQh0YrUTm8
cKvFoY0U/8MVRO0QZnnt/q3dKhU4RmfFb2sChE4gE/FxygEbiI6yRoVqrwZ3
yszQdbcyIWB9EZlHcjhq1e04wOBEwt5d//vSNXO5In7xl+8LUkKfUTsmY97r
3q77tRMCgo36v2k1EhLCZCPfjS10EnDsfPMJrg1UBORTEre2hjiP3EFW+XbL
VgS4rWamUPQ2YbHVsveah5Pcj+YkVrRiZjdKV2v0XVRXUZYbYEQ/F/YdnHTX
Kj9HEDoVE35O/w1mcRGCHWiizO5vDur2LJGhlSKl/WBSsX6I6bb6LV4B3GWa
+bF/bq5riDh0Sj6l06RWgbNtMAOBQI733jOENL6NmxlzCy8wZP0uRigeQcMn
q/y7Zbl7i3XStUwx/YD7h4JmgxnJKnnfrzHEf/TFXGwGP5+2Bo74XYA7aJbs
u0XB7bZ8Z3MOTWRhf/BZEn8RZDUgZ1ZjaOivYXWxxPbGrjSmOg4G/TQ3bbnQ
niE/0DukIVtsLmsOs4J8yBrCRCvwwuMRaAdytp3jvphHEGpwDY6mqfFcAc3v
jDvuWoAPjXY3ziTSEiTToEeSfaHd6zdVNPnFbL8EuFByhXrO7wpsAl3BTB58
5LSHrzhMJB/KwYXdL5wnICHgY+CO+BzKjEJ7+/DlQyJOqTqTq+vYa2wvFvIN
yz4cHlLnNolV1myL6W084cf6gFpVjYE8nWP0ZsibuZ8UXyEplsb1esaZQlI0
bTBRoj8tQYs4llmtY+iBzfXldqwgy115KO0jOfAMom9l0vYso3CL8HQHo/pO
pRGwPXsj8fTGLrbNibqZfv+STrIaFqKX652/V/jgCAky7wSMTHintQ46fibO
bqzKhkWFy21feapOL57iyIPGcnbMAeEqNOAZUhqNgNFMnN6mqH2KaLL9w4u5
4n66rlCitp9wzSBTXktDZ9BDPatw89GskqJSn7CZ+M2UtSEySDQ50g/11g40
QLY56nmD6wHY6u+827QJ8NdJ1LS/2GBXAGP0Vzve7YPlkAMZXodx0ouFUdGN
dzvp9aAr3Whpg66AR+xfCF5SgtM5BbRQh+8sMbfyYs3RLUHgPbsLCOvIClMj
ltAQLjDvxe6nO2oR3VPVvc0/i12j7YiYuiEv5fp/0DsgRvtJCFNhPDHrccjh
TuxPjC8sbL0DVSTdVFiveeL6TuE9yorkCoMY83reQfrERBpvbB4hgQHXXez3
/Ava8hzY1fEvAeDqPnMPIbg74d4qN7zf57Orul5VYl/oAVMyNcarKsUU3slz
8gm/cZBOSCAOMNfkNH2DufZtNlUxuWEhEQ/bT0fQ7zn/SfevTvjaToKjfXAA
Kb2gRmd9JfvIAxN+0J3ZUTolwD6eDzv5Ek5tPXkztpwV6K/LcOt4AaMBGKae
ZSvnzHlbulVaMzmsVTfTvYkxbTv06Acym6SUQkNohA/xZye707SjXFWoisdb
golu+x21CQKl1YQYtJU0lhLMgNlC14FVOeLQUk9qJnUQ3LBusBINsMy4vM6U
mgtE2YTgvSh0hVUGsGmZScaGmHAGzBmHdUeAPQkjwxXqW8xDzCSUBrgUfbMm
6Jmz2yOBy+5hju52ZAb4RbBDz8YXOS+EKsP+vaQr9wiS+M8SJhQvMgVrX6hb
pj+nRdGcvriBCxBFnLqw/VREiU6fCovq+Up7tKSUPNYz7B+C2LU54HrYHsg6
uKErNeHsF9oKtv6E6rFILHgDwJCsrghn+Q0jZ+9ZNJmf61qDFI4xo95y5TuH
/3KnVyOdC7Tt69aYfiAvenom9lJlF4hpVRHtxAim6kcvMoleZRTJiuW4mRdv
csHeEkeWy/c4ojvO6J7AmRdGHIKenRPRP4O5d5UVjOBEqoZ1jMJACOpjfj8u
E937lvAA/nLN1rbnyNKOUrtq6/gB6X/0uVfbRShggAsVNUSQsQFd53GJURZs
am9hNTL7PQ281tk+h7VT2V4dPNeX/jeJdHwNQnxzjbAoz+kADwFqvdLqo60F
u5TKgHjZeAGAqVwlW1iJF6LxtWBh9DDZyaZbcNqJ9VsVe3e+K9VaNuJgno6n
re7/9ifS/FGcabw7eKsmwl3YlMkSMI/yLi7Zt6L3QhV3pz1SVT+gH6P9G+n5
8aYfNUtzkYQ0qHus0rpU/1rBefhP6v2PQJP84rgFU47Ecetv3PNaG7sXO1A5
czIoUmWyWmICQNrel5u7NIB+qZsgWt4qgKM+uONHWEuDvRdUcRxeEAD6vT1m
QS0BPc6WAtUO3yrQOqbU19iVBvDdfNynWh6v34GO7P+Bjw0wv7D9UTHIoiZJ
li1CWaISWg8f5XFkByKyJT36pbrTiatMDi3f7Woh5s2wU9Pn/2JgUO4eP5fB
D2nDHjL0XDFqDACOFAKvqFgKUVEjmnC+DWGAO12/Sq0Z3/WBC4sETW3uoOuQ
zH/ue7IDGEmwgqStZluk802derLfbDCYf4cIjKljkpK7Cjt4uBqA9xDGy63Z
uVAE5sPC71IQWzlqkt/0f2PosPXXHjwhyfJ23PdV+sIisIzkqbafwJs9Wbt4
KWI2Si7gQm3+0SjQx/DJU6B0U3D0fIrv5sF8xKXlCxANpSb94fOR3G06tqQj
IoXbpbWxsanMsyGn2e+P31N7oTAnlPfm8QRaXls9crhjgIVs+4kV5SNHex0b
6yvYJh2aXnyeygRyy8hcc5Uovo/lCy7k/Oz57DWVljT82qqbWbHzufCtSYAd
HoriWlaJuZtXx856Cev3R2Mr57A9KStHjX7FXlb0T37cY2Dz0LqxCGr9Mqb6
Qe5bZ2tCnphYeBodaAScsemQ2GTQhQNBTc3dygjgpOCKTK0URHIM3UXYjAqI
swgeis7S3k/u7mX+FZzkAmBXhQSMh2pAc4pIhU9ifct3YpedkYYmpYJkW0RY
Zsq2No541IwxHOwPUFot6aNulEDoELvkSf8KPcfpClSQUed7tpct+5mNdPsn
KbOwhNxOJBPb+WVgIK7YcXZag3/sClhq+gU1BbxD+2fcPIIMf/1JemT9DCeZ
Jc/+P40/R/5rgVP+FOmQLg2LEThDYLP5Ds8jVUhef1hs9stVyOOWkunzZt9/
HOXiRJ8BgGms5CgWY1+BdDbpxMBZOLKZeeGSjf/4DSzS7caDC3wpfa8bciKj
W6hJlPEXxpQVsNrlpbF6198ChYGyy2VnssTWEzaW9OpHcXXvk/wfys6HdrqH
KdyDK7rogQsyeCAUGtzaCmJCelR9XlDGu+OtchPb4s764j4Xj70aAeBlkH01
YQ2S9bWnvDEut6zeuOcmj11Krji/nGK+eHOVcfv4meIlFLj0WX0QhO7MRen6
rz/nayuwtpoXLwMDsxCVMZLT0GoAkUwoCCysqcn22LxOUesSlv+zjOwyT4xB
XsVIllczSqFMTS7idYsRyanyzkGN1kOIufZEQ1T1kDpauG2awI8jSmXAI/YU
By6AKWGlYjaVS1ifm1Prd07EMgGkaTCiqwL3okYEHaL5g3GTpuuZPH8HU1ba
HdjdlQ3uww7NrQWOfmP5RpuM9Qw7YoDRzBhkgTyBB/+zwTCHyqeCuYtKDimg
Ox/66BF30gSsno58TQaq/Ft1w4iCn6Kfx9rcmbUf61TpA5WnARUESNhSAJYp
OyqcVrScq2AevJhEW9GuV3zlck9l1IXfQRktd6x7RV1XM9zxeZUXHeO4mujQ
PtId75q1uE/KLWV2GHxrF0ek/ty7C10tHsVKdp5sTBZ+m9WIS7kGfOWp6Alq
fqRXQGcIOvMpE+qDyPAMojVkOrS7/WyhIkYdv0s53VDMMVaTMNBetyX4aKNB
rWEtP4HYyYGVpP6wsyrIddd6uVCH0aPjonpBYgpfhm3xwzk+aHjoweAT+ay8
DZOavBfpVoJOys7XR5Wgquw9N91k4Rry6DOAsfYSPhugpFp0EZvlB7yQ/faE
rGwUiA0/Qvgh+BtvdvS2BWK/EjJT8Q9tlb/FvRvdnag3Jhh39wDGOSIvD6sy
Vn7nXYbX8n3lbdPi4/YlNMn7UgCAF1efmjb4U9S07xnDOpdqGE+z2/P3Kh1F
BcnB9yCfZbW2jsffIdFu2XRsNvsHOOpdLFTUc+g1pBzPxWfsl01DXYEQYCWb
xeplqUhGjSeZcD/Ve7mEDAAw3KEc/f9FrobsBmmDYkRWg5KR1zzmcHSSnOB0
mcQqTMCsIwzaw1PEUxfZPPBkP0sh8hWAvLki69sWWwd5jBHfM8HE0x2OHhWJ
L6VsDgJe/xX+3He1TCoHjddd+AP1cmyfqaKcFcJVOhJQF02o6Ny8zCFpbLe0
VSu1n+WcJ6fF29yCTXfrCMvV2w8b21Jg3eBEGjwPi02ZAT6YR6Ms74Bi5HAk
+it0twRCBuoWPAJlNIE2Rd6FR2mV8G4kfddJ2b7i8KhTs8kmBSYIPay7dKwe
Hu+v/jx5rSNKBkjUvATmCYD86mfnTFHPKXwwz367HFg8aEmSnGE543o6GBY9
cg1MID2C1myyxN15mT4xgE+u9WqiDfUkeO30ndbEDETarsPEBw0VwfuEPZVy
UtTOrxBx9Xy3D2xdXvm1ujPW0KMNugpuzQ0MuVx1GLuhWVfVOMFYz0fBAwmN
w86AMs4FiBIRv3VwPCzmGSmqXwA8IyMo5c0wo2nG4OoxKH3Bojx51iGNkU8/
1fAyW1IMwg27cAWtWGG/mziyy58l2uOXtlRzSMFT05zilubW3v4Qd7g2GBPP
h5jasnfUkviOjwV7S6b/naov7+twcUZnMjaWHg6RFWSHvYKOC/q3Uxj6t8//
vNoNLy2y1tVdLccZ2iTE7KTG34riGqluSCdSfM4d6QFOIEVO7+gk95PH4NKt
pO22SdaRtMDRdmDcUxbnlS+Y/ekWWc5/5HGm1aIt2s/8mXziYX6ZVY/tqYtA
/NrLPLnKrsy9Gb+Y+mSC4wWyX48v1CuSFq/pAOn902kTrcYudXcRTEJ1IzAf
Ex5nhwAJZ8DjfzvVKeiUVgNFlwhOs686Fii5otdyDHIWZ88BSbcvwtsuPvgK
OIkpyXShzbQlArh5lHwOSU4So9WSmkRjZrfHCb7l8JENWvuDymgXoM2uASuM
CgJGIl0sJtwbix8/ehkmrHEtBTTrV+likI+JEhA17NyZDlJXnul+bHiOreNC
QTpjUJfmJgNAA+ZZ14n6b2iyDaDINmr/dDES/bloH1MSinhwIKiOBnvRC93o
H/X3+5FOs+5LejjCgAs9Fs8Z1a3RkiGXcyMPXGSYGDD+EQrUrMi5x6ad2bHE
hEnsCXG2CEOTWYgAFbMPY+IJKQiniA67S4TzVkoI4DVVb65ITMlDsWYOnllm
wvehk6lRGtw2ChQTLN3mxHDRF9ojd22UGp9F4GMA2N0I9XReXTJuPvapCSx7
JNVNmCkzlPw+0ms2KCvoq2nU8+4P4wUYMrHoFMUvLCI6REiZfJpS59TcjOsS
0HRaukNg/YLayMYYYwk5UYg88IuENsR2tJevLMhmyK1/cwcc+C+KChH+NAB4
2FSO9Yx9LR4gD3+tY5S06nFlUaT8NDMDTSyeHLPh0TK/0UYVKpIJc3AipVac
vNDxnNocMx2LOygKH91Z9zKoOueGiQ4Oo3qYE6FXA2ijFvpWjPYHZyi4XOor
hkhPrwgQQUHW0cy+BP7OIHqY8cP5iC88NOCMp43AQdtSiEoeFQyqhaQP1V08
yz+Lw/UnGNZqLCeo2jnrbae+Xo1mW3Nl5nBp4+CC6OKPURYEBtG7/HHFedbs
E2t+JP3ddabTVZjeYH+Dxc5+wwL61anXbx8XEMpJad/R4CzhdRRrEqxCj1Ja
q4qBX8OSbO4pAs73oTlVfCC6cW7Ok4SecqkS/eHFRqSIQmCc3guWTZq/6yxl
JUBrLcHqq3dQCqnoJp9qsPW0LKZqevAoKsBZJR3K4sxfhbrohA4u7McsCFcm
9R+vdY7+qa/0elIrv4I8cTDCzIxQ1PzO5AhxYdWQMrV39dE6tHn25MxBVleO
Zu5qfJGbjg/Goazuj6DptcBpLVdTwEOPA26a5smpwp9VaSTzF09IkSrkP1vY
Sa5U2hOvVWcPoJwc4VO/EL2E1liZbXlB8QWE6DOEjD05vEMs0MzxKx6pva69
41X+c7wUMRa8w1rVXA1A4NPVyrzkAHvNmpAdSopRSmXE5XuNKypjrMszmIOi
HzQKMth1vv/6O8gvJND9mCPC9EAp12nVBehmhZjfUgftvqw2NJ8lK/9Ksyup
m8e7LJjWUgIejqrJjMFSF25wGLDckNBnOrR8LKOf1Pe1sdGaSp7ZtplajFiU
wvnHba4aE3ZHs47V0eyyPA+O6h5b636haBBOISIWvggQvo/O56snaTsblcbM
pFo7XEh0GVSkFLRmnnoJVRcA9/D0Ou4/hRPN4ny+ilr85lVQBPxM5H8gDBjT
YfA7p1sPrsg80rphDj7frV/IhH8ZwNVUJNl2BKgH63iymcAswa3p/tV5pAwR
Wby+uWdv09GzLI2KgF3zCv/vxX5Xy+BPNARlC1nucLAl6mJCbuo3/83Mg6zM
EUZHqcf1hO6F0xGRTBo2aP9kHLzeYYJ2jHzSXCtshCPsJrOSKX2l5ZK6bbyC
w3FvqyeYMs2bVpBEAwVpq2zV5vFEWsfbhiyIkeVGwMB17EPVzBxz4DTNopYr
zBRayi+o+OHKjg/K+F3NSWH/RAezIFqXjPqcVIMfncQktC3QlNzGw8m2/9e9
+Xx9qFdq3WTni8ZlSQwKc5Cd00GHMtSce/Dy81mcmGloba2JghwwWnwztUq4
uans0UBkdoL2fa3a136NyyE358Ebrq7k2/oV+vj7c2x32PI3yzKcYC2Mj8wF
YyV//+95sHloEgTPXMUbsXc5LLlkmh7fGy7MvkZGxliEhS+b4+1R7rdnRtfC
maYfR/VE9Fo52irY4sg1r99yn1dOEuJhbPxsv6mTmwJeyEj2WNDroloW4qxh
uFHcjmapus2q13BxgFzEgE3ff4G30lZPkpmEOkqy0vJp0WCB1J6CXU+Q2Hx4
ZqjRByBnpnGNh8zMdj1E6szhb+PJ5mJzDMplt3fbkKl/M2aP95P5wB1lnds3
4TPZO4z4Rh/8kSwu6+wZkZ2bEUWtmH1AMWXZt/xKMU9wXwKQ2uUv1A8UjGaW
JnTeAtjGaV/HfEg1ov7Ox+p251cg6ZiVxHiDhV3XvILFDFLfsGXJScEZzfZM
RMDe/KGDmJuDFw7L5pOC6kRsgkskC4tc2lFA0Z9KS4kzJd4nstsLZWtJ2SQ5
ZwEt6EXGq7N/oC/7hqI88LiRsJlQoeZGxUXFU+oFO50/KP7JrNvNSj8q7uy1
9/IP/1ZbfX4AIF8i2uCY956SRjQjgr1KJQuFjmlYPfj22QXF4oJlOFK5Ejxi
2mSBCs2O7TbuBX4EL5/+H36E10ZUiT/QEKkRrLkFaujXYBuZicLARif0WUp+
CUFng3qpFV9gg/48BJ/n8q0umtgZmpzSK3q1+HPECUmpTA9T7qM0W5RtuRGe
+QOtvagcpHYyNi9grTlei4/5qMqfSeGmjSyI39ZPds7CbPaeUA8IMLtQdie6
PNyqvrD/Q+ZghabiehfuzXjtDbedXT2BX9XNcf0SMRuz5gb3sDAgVoU6n3ST
/tLKNBRRAmpnSov7t4qexxdH/FAmZYTqHM58CuT94NkKMLcbxkpdXrx72rit
xFnVU3zOGVXMyA2YxGnYqeBEELZbAtSlDPuGnvYBC3/RWHpwWpV2JOQEnXaU
5vV1lCz695gAT7yOHzikW4gwc6ATocXk9b66qxiJ2sOZnwhwjqiOnEXNVKle
j8QhopqQUnrxc+l9vmUpaKtnx3IdkCdxLg+V2U62CK6YDYRATpEGfWA2weZK
4++hhwPnsExREunrHPkKkio0r6nGEh/DEZO30g0qYsTxHxcTe24fLNGWmonz
T6XddgK6gkoA0GyWnX1MGKsA2/inL8o7yp7oUcntuSKjEePJZ1kt4uWaIZnh
ChV22skfJuKzaI3RW4vqIzq1EInRqxvzdFPAXLJkzX6m1rMV2gKrniDY2s9I
qXxjrPL3Z3U38MCX20y8mj+1RuFNdAAzjAUif5KkjybJ6ofbTof1HRwKmqLq
G7a+5bFANXJwpF5kXTr1MYSjJa2nXJxO55TfJiV2TiLexS03K39RjWaTb7l9
qqxRfrcwDgEzG5ApQZLfZAZDnmtzkdeCanEl0e0j48NrndbirR6U2hTBr9LA
TAVHhWSyn/Uchki9TlkrDYM7sffzHdByFU8QDQQo6KJphwzkDwVcnpkf53h6
P4nwHsY7dXKRETXXGg2L6bgow1OlBBal4EPjjbcSNxN8HkGMlkkSeWMtoxvP
9AmwgK3h0CAf1DJPNt2k/Zt28Juw1YSnUWCUuDM5dpKjlCEpIIr9fSJfR7k4
My89bSU5PvDBQZhh/sZK/R5hizBGs+UFqGU5IUZD6xFxzdJOYq7lG+9Cqccw
s9BPcW6tLVSHMQevifecRJyB2hSdTTT5EQfrFADv0N2ARBlKrGds6T8puC/8
ikLNpPv0tzgwNASLs0bPma/81Ma/sgEnVNHtu8Kmj6ZJkwuaMHyGGaipC9Uh
72TzPYLbKOR3CI92CJBO07J3dgN0v1FdPk9m5AtcuGcOaFgefjGpJrtWTYoE
aB+TQeA+JCc7mXcdiGOoJ/LgI4cdM89Li529duhgHNgqEvaFkFRivnon/vE8
NpWa4CFV6dZZ3XECCwlbnObMrbqT/BMAiPgb03sT8+Nvs6lkovNeqo0TWQnw
r430OTnAJ7Inex3vM+zHmh0yTPirOE9LiD53wUFsyHQLTJ9dL2LLHTwOp3G1
JQ2goP1P4yFKi8eyLxCloivZ2aizwXOYLZrlV2TMr1tfugkTPIJ8Ztavokd1
d55vq2f1/X4VncKq1lNpyYYMAyGJ9WPucb6Vo5TGYohJzOYqPNiw8OTn571m
JjjfF8nB1ZYFrXXDSQQ2ZDuiHqpca9koPp3fXr5EDKgtoI/hAdk7PPyVxMvm
EC41Llxo2BVyxP2egZC4e6MNg3Q5Z+ZtqsE52gdhWOo9OVVmxiWyoCy29PIE
OapX98429zltLKyH6CbHc6w0/opG+DPc4C/50Mhpm/0/ckPvHHeeVxahkp3B
XvzaheoSrJ5nB4a/ZwsBelDsZU45mUFDz8ISPfoE18VPq3hf8Srg+N/5Y7W2
XrSWyMjvzBTFJgMIhDmM0XUHRO3dLXqxFri+tn/IMJHBtJy1qB9v3E6f0BlE
6fdmV/2Px+6C5vCPut0nC16fFvogs5tJTGlqAhGfVO3frISsydyIOqfCaqpA
2L1BRwP3mxmCQDcFSV/xcKn6wgub/aqhDDwJXFu4fiAXUTsQbi+/KekIV9g/
mB2O99d5048zwCakBlfyqMCtaDZs9v+H++I0QvxHUN8glmfmkwqdWKpJbGnV
ap6/4/qRVxyyKqP02Jg7xDwbYTwR5LRL5U/VKaOWYE0BqS0azy9DCR8C+1N+
0p+rLDTeyVYcdoWg/U7sx/AhPPZNNyTJ0GiyaIc+5Y0NnHANrXPdfYkyVo5O
UGPzi6Usn1YX1f15Pl1y0ecEZpsyzHU7tzMYHLZqGUthZ68oN/Vj3lr6lkbS
XhITQSAFon/x9r5kAl9ckiZAYcux0C2Tu4cFoFHliO983uxyGLlQJhSyPrTV
yuahjS8vYL+3fLJlhOKroaSTnVCQYA3v2WjpPC5MBcqukn2lOP2hXRYW0483
s3T65Ltjd2U00lnD7YK2abtllxSrTpslP7o0yyo/fP5LmwQe0wG7SA6eiUwk
IZErq/buUO+t91Lu1BrCJY/TImIzIrD7TwMdj5Ck+yNTtTniNkFgg7dRVjuu
TlZ12nCCSejqOew/+OjRueMAARS0A3FJAoDzE4SiXvPik4Jb6w0/l0AwFt5J
JxntOppUS12I8HnAyrUEJUS4QenPFaAuSgKrIwjq9k6wFjN6QBFDBq88x+Ao
LhKBC7+vHvzf9BrctDoOsWOQM+7yQESIncj4NNAqu4vmUWuj6s1wNty9J8EK
ccFx2anL1KLDULjpXB/zA3x7SUg/c2kB7PeJjLy4ps9ekpxVa99/NkThZ/NJ
1tmO7tz94kzuk6Ox7zQbpY0G6pt9vIjcewl1xi85Npaot89Y4GllATS+czj4
uikV6VIuUca6HScW/HUGoOwvzmXnaBH4cU0bxANxmiSRw6PHP6TgUNW7/hMr
86Qc/JdIStGzNpHVfF/PQLg14u/d/zdBEA/bxG7yhE0QIiSgc3iE6SOgMhZq
SLaFRJDJbc+S/IcNPpDcHAKTMLdJQIBkjVEyMF1whzrBqu8zmSq+tvOhxuJp
AQHHuuna2piUYnPKV6FIN52l3jr85XTVT2dSE9Ts4+Ias4qStyxvDtoGKZlb
/XeDq8qdlSfkZmufYsAlOyj70b+jnpQx+7lPmAU1RmyGrdVzWIy+UrDxP8QQ
LMFjSiKl9OMiKoAEo692EDeY8jRa7TbudbX18nEZmjQV7GIhI4cvmWKQkSqv
09n460hBvyXGk8zQkyWHF0czH5ew1jgyp+QzMVZQ1fxfmr1f5jAadaN4CX3/
6VXWAeHJkESej1nkfx40jqUO5a1epxCy29t26/jCmYgCUvzSUIdlcLsaWEHW
ZApbzFwWa3y5F2Dbq6SCzlcKek70ackoXz/UVMurUIiJ3ADSxmqGy+XWfxZ0
eQk5nyz2b5ncUIwipAQUS9dKTFpcgl5rnDT2nIniqxMCBii54dnUnLK/7vCn
Av5GpULBAvIsqbnYStjy6sR1Aqh8n5kpOc/74qWah3l2rnXgt8Gw2sL9QtiW
sS79QZNC6fy5mc0CnyH0L7TX4sSbSCVeo7AZQMzYSerLJFN/6OXeYAsRu9V3
6eew3DNn/+yeApYhuYjTJe8k8wLD5WwLeNoj1Mw1MBwWQsm44/Uho1IWQEdU
bKnqE6Hj3KHdl1ky2kpXCNMRTokI1s6FvCaR3U6a86ZUKN///0qgKJaE57Lq
VFWJ2z6HdpDhhGHYJgL+zyf0GahnfeED9OmmT41to84hZT+kF+d37CiSyw2m
PibD8iDzzdGZXKSy2v1oPkSEorePOXxYBOUpIDqIyWEVuPDttmVcCtMrv/YK
NDbDOpfERURTwJKep9hCYZG3zoHxg3JtHpXcaC0j+LaKA6OSK6Qf+4DWCa0S
UCRrk4UOGTdAwI+25UqjCP7IT1dZFo/yU3lyQ1oHG99hK17wBDL+NlaZGe1D
6Cbw7EkIUPqZYsI6PfiODXwMKg434dT5UMlhIwkJ6mkSdEkoF40r5P1BhClS
UzJCJxQQbgXJmH5kuN7xJhcCnpydcr8xSleNkCye5i3NFJa7Mgwz9+x2U8kt
Wjn+DPOSELYGoHaWhplXrLXjRqzGOagHUtUC8kcbvT6U5de1AbyN21PoFj4h
Uexn7CuohQVOfxjC7feHyV1NQ572EiHzVj/s7ug8836EIreOTMya4FFXog6K
g0pkKTkJI5WhNsSRDGCBPNoib1xICpnbeIt7QlaibPaI3Q0nf/CIFnznaNoT
/sbSirZGJKUWrOL6JLEmVn7vOH2OeJb0D+SikZdiHncC7Z7IyhkYT91t8iN2
hCQY+CE3sLEnBujAiWAv0jsKMslbVPWM0/u7zXgyFUblrXsHY3X8KQIsALu7
TUPu1fHFRdOCmyaS9hPtDm1sHlVvTP9QJOObvmKbbvvr0tVirHiXYgESuXqt
/bSuiD/36ZivE2l3ss8sshWW6MhtgkkVJMCHYEduaj7Ym0PScoNgc0RcH0Wu
ersfqEd7vfhxseRkiu4FKbAxfQ6EfZzQrpwkXnDAjgqXuuwimncKlgoaZATM
u9J26VUDWIYzOwnaQWNChJLBJ2wnG0pJf9cBmDJcZs0QmliPB8XBvE0CODPU
5WHP+amsysbWxKO1f6+OtGTBqZq9xzzMwyqqW20qIEZ0TVMmtuEp9kp1ws3V
FuI1eFm04eL6cz+R4B14UqlHCXJeoViZTgYJjH6HpnSKyQuYCSYb2TxPoA7V
nB/tShoajvhJwJigONVQOFeQfMaVdisxpH2Z+Hzg7ZLXBrDiA1winmBrg2Dh
xcu8JX2QY3badiiBl49ihXJE9Dx0VG0a3DKwubf/0sFn2m7jERw0DHIHGBDk
Qf1KflPtlGXyP9iRxF1waYcdmdG9PsK7fM09+ZlPcfFLUCBMuItmmfPbTZCp
K8XgtJFiJGl02MIkQ8lb6bm0A/zqXqnBgXO9+IR0srukfdjTsGvrt4sFFLSv
RTB7pUNBSTb1cm8gTC++/j7fkThuoYv8QRdWRfwc7xxBIWeyizE692iVZVdk
Tl04YhTdBf85J39tU3np7v3GdGP1JMa6U9kppmP+E86XB8mjSDuzxX8QfMIf
t6wXVzPSu5C/CUJm0KdwYqG8Q6I/q5GmkC/mzdHy6bYmqhDM02bqzlMcedAu
RWZgCnXfJ/0hHdrmHY+dVeOfyZoE2MvdZf0Ke+Hr59Iht/XT770U561Lntkt
lV4e5ZVNnTaglefo0vOqHWSovT2zgwmPN6tvDwz/sC4SK+Y4RwHeihQAt1gp
jKfryQd8cqmAOrgRMqXVBi31thX+FCBi78VkUkV8+mag8r+tteTSVrwRj4o+
Du4bCMyDmFVG8fVwE02Ctzve3Msv5Gej+ysyMAmiTTmVLkfnFBW1onGsso6Y
LkHuarvkXMQx+sghhKKujyXWaNCVRtsWRacJDBdj8QVNNiUjAPD1KCttf5dJ
rp3Hsu7b30mgbgr5L2EbTVsd6XP0Xl9eGccrABDwT8APdmkMlzIn2fowhf0A
fi+r95SXIr+nEOsh6p1u7SKNoKKCPpdMBQuHywd/pSIlqHBU+4T9Nay/Nydg
yfwmp+lA2V6gn5pXREWFrQTlwafWqU9N/zasPPq6iD+MAtDM6a48TQVzoWmV
2Qm6gq8YtxpwToCBXDTOSp41UCpNqKLRdeXMXd9pbOl7eUTefKFNWKdkdco6
X1qYhFrOVIAmJoO1pmtqbd5Kt6JW2hDmbhxEz31cnbP6MTlfKjBn0H3SgE39
TItbHF253QHTReZqszi83pD3D5dD7yDMOCTd+FH9In3aER+6DcbbQ4LRrjVD
mQL/IQGn09TX8LBG+/Xe7gpxKL0S3akiJ9Pftq3ElwzaJSYuaHZ1DgIjaSb2
oQLunAnDWXNsr2xbb7HGGUpe1Kab1EZje3SV29zNtpn64q2LWxdrX+tjbTcq
RNAmArkYzN5To93BK4A9HcD6YnAVuek6rTj+thssPNllHL2XA/Q1RddGfgsB
YzyKyy4PPeTuyj3sIT8C1uB2BAA3Z9OLfDvE9JmkQ7MZbYTBBDD9qW/NTHNI
cVbm96i8T+azaVzKhUcOm/ueQUOFWS6czpP9+OJCnOMbP+qbvpEBdG0QSIFq
YQuBSYsM14ai4Pmw3ZFCuSIN7oz7eUBq4vfakUhr/9agIhBkK5MLUzmh5mje
I/XOcDl0yuiY8YPGJnFFFEtYW4zfsYLbVpgUVlVd7AMz7UmYqyH4cifKirCS
AuxbcA12SVLUuwB42b7uVUD6UZnHhh8AMuGMk6y+NmTMI3oee8WFkiPwqNZJ
kbJmO5ALtLrwOnWkpVEsuXl5Hx1EQAERkecn7JsqCH7j1I81N1yKNMh7KVti
qmXUgE+3ECoTRV1krHWQ7RiKvqL4ax4oEATj3NvlxKwZfEFMptre70DHsMwo
P0T7/c0ewFXNTzXnTRf0sz/2ZEiCH82SBZ7pbSMFlWsNPuixC8EJB6Kt/tHZ
+PCAHAWI1rQ+1zZYkvSf8EhHqU0O2I9lYTO58enj//801LBsmcN9dUsWFCl3
k8uk0gQ+0sTw0H0ZZICJ2je15QnN3ccOlnAgB74aDPJLp/1rdFrMAKeBQV28
CFpj4Eemw8nf03P0/UtQ95F6lbKOC/rLWVOSrGWplhiAPnLV0IR+hTy7wUbk
tOscuZDX3HSPAHS0aPBIcPTfprC8X5XGnxHoDN9d5SWOlqCdQ1H1+VofRuns
KnB2IDwBvqCEU9oAdQmN/mdNdSccq1tgw1EnzxtqyzJXxJvQDSW4K/Xe6fhW
Tr3SFKbiQzbJKc6THohVNs3SN8PQmVYZPKsAn6xFO9d13O8mmeM+KolXIYkE
VAIZI8Vtz18EYddINsWFJ5APemvZkcyW7kuG2d7Mf7RttmyZIc+a/9i1jDwA
XMoHEd70Hq+xD488NHJ2hZd3sH3uTaFQGbpci3piKe2Y0WgtoPg3Z2kR9w3w
RS1gONetfa8zrQzGYYx1FGmYkU4YJX3bbnVcTwPznYPPA6Uij9BtZz7MlyIN
MuBTr8oLpxjlT/OwdJdMMBpviNH2dzxPWGxtx+61uQuXJp7LHasv/EaAQ1Dj
dI0pq/lvlTgjbWbHmlqdPzyfeo/YPmuHJoq16LhLBOyN75yV6BagP1BdWWZp
/BIqA+Nhq/Ju49DaHtbE/nM5/U6EP5yxLcogWlYIaDh13Cas28y3k18Y4hAF
GOpKE8IMkJ0IF8uKugNh1EpFPy+ouczHrFkECcG0bTnPe6wtxVvjBUCFInJz
6szIYPxkllRTfw5sUCpURaTOg7Q8KMhqSvRwAwmFvtq6lD19hC62Q2I8wa1I
hFYYkRK1muLnrJR4ZMS2IH+ojbBYnUw/npXDzWLT+vElZJsSwHVbVbUAbkI5
uspVERYviiLZrInRh49bO5xIFNZ9EuqPJDLirNVPhcZlPPd0By6HXF8whH7W
H4UBy1OT2RTKO9mIbNpJubRhByCwLC+sccof+MbHfj7TAXwPNMBONDsXZjgL
hNyPPj2lCcUPZ4q3x7SGQp/w06RxXEjvT1nqQ+2kkBYTrYwPKNU1imkFpWec
Ccyakjjv+Z4uFdbCKcQnY0UW87UU87KlTryfETu3FbO0Lcn7x26tQZRdNIeA
N6TqlyynQ3pLzjQzyc9YUeM6xHLsFX1xCIXVyJe6xeLK3DcnHXzGCIPS3V2l
1klmbpB93QDPeQTIVbm/tTmMPVkB+/M/P3j42mzxrStOpMIHKSk0unvsEtok
rj1WUIY4M5Cx08zwKmk42j0Uwwk/MNVz2Npg/w1vxPA5tfKIyFCaTR27V9LE
6LQmKYpr5JyLN6HK9nqiQqTG/N6lxOhjVEhApigCMzERbGtrrt/6PhLkQf4W
i9HN5z28PIqegJVZ8kM0rXe0ZDsboxd8o7dFOieRJz7BoQfSOz7we13HKEhh
kUdmtoMjn7P3ckM+8PCG8lA4LUN394BWdjwvLCykzK0CTzs9iFBvOxExDgzv
O4/sm8hzclE7tDqVfhjAL6xjL2OlONv8xUkcsj+foV0cYJeHz6tgRKFJJu+w
6G6EFGtvFHBuLJ7w7cDEb/kZDnnOqKZNNXADWTGENLxldnJ/cweBtoZRpm3X
X2Xl8NKTKMwB7ojJoIVX+lE28Rm1sK8Msdr4JNZdpZLDZqmEDM+PUYGbyKhy
fR/zgooray+3IMSarQ8eQIAgmVylFIHmtMbeOO1xzHCXU49hwYBuC6xoz6Up
MjSPEijCoP/h69NNQjTzJkEpjPudzJV/ztFPJSV0cK6/87d8XLZgAg+yoCAl
ILg4uH8SdYsUpzXB9tNP4gLbrk1bzYtvuaC2Na0AV5TLE2r9CpG2oZejjPvs
BH1SfOAMdnwNvU5yxqHOQdRQZiG78ZtGRw1EZoCHw/0q2ZKXkEknQNv3Zh3L
DBKf80QXW/lZKM5bYlhRZFaQ4nsHEr4exc5n5MXMh+3WIVupL1Mcaw50aLzV
OskHUBM1AfiSZBxZO8h7mZsRszAjfE/JE8pWZHrv/ftDtw6NURoElmBzq6V2
9MqBsCNi7tz/guu42DxkIPNcIRnG3akFX4TIIIZByDT+4IE2dhVkc8V4rP5L
oc6DvrLSKfelnIwYDtMkFoMGfKvZCDtfdji5DQXzaL2nSLk5O3PTbO9x5O1X
KwwR3CX2KZ+qEZOTIHUgs/vynnVAU2lNu7uwb59q1ovJ4rH4FBDjsyPmIfgY
sxNYg17qRzd5FjcshUbhbhCHHcDb45p0eQ4o9TI0njJ97PhF5RZ++5RMuYVA
nMvKYB0PDQ+jKPkAPzkUDA9nNGHacC1MFvjoogU9znJQH6lNdlKvTqRxKIwT
wPHicdOdOskd7ZTiR+fUnxjtMzcWT4o8u8cHdjEuoApX7lSXa/9TLVJKuzpg
454Q85o76aokyFx672H9NJIc2UAlc6jtoKpG76S/AOt8NvBy49IFLd8NnAo2
UCcRLBpC+X1kjvQtWsOq8ykXBkKXBQttvdZVE8wZ8Bc+UGtEbdXbRURXRDf2
nbw+aMtrF6EXsVouT/PkYsRaiTPrrLvBTyzNZgTvYC0vDWfjFQr7NEPWxDRZ
PkvxHNbgSOB1MZYwePhwmJXUBYfcnfobdXPuwtfpkWNUaqcK5JOWdptyell+
/uBXSYuv48J63k2X5ZqktSmKwbGNXeYWPHbeMH+f+csCZrlDOfkuMjZDrVD9
y+7UKf4tobX0BxT/kpnaQffZjJNGIi8QpijkdMSCsZdYyd9czhg9TT7wD5lm
kYX6EjWFvhpUXWRQbRjT+2jp3d+ogb9DAAv/7KyRBvHDnx0DRBeUi72yZohE
aKE2iPipW+oapJIjZ2vhfsg7BlbVi+RnzCL4Euu/arAXe4p6LBsD1ll4yrdZ
ftt9ghKYM6K5UIkVlFM6AS5gHF2fmBa+MQVXMZRTzA0+xpF7DfXkRhzzCn1Z
aYZXgwbbgbm/zCKV9lj5ryNEgoEd8omLE56/6cQiFsqaCQvBssYvqLlMd4DV
2RHtAkjXeEFIOrBbwoWTGyzaX/X/e3SHfJdTwmwrbZwxdWwnHgcsCfi4LnL+
HHbtrgunjoV2qhXdgzPAOaSMUd9669iKQhGD87dfKqpsDqtjIu+3nY8uIu40
r7sVJM3OG/OxXRy9K/D5YXASGrl7OvWM/pDcaOW5HYT4Hwwm7cE+uqCbHL7m
HhI22BhmR4E8YlG3h3aDNz/zdY6uv2gjBhXkikGBvR+lu/YPEvAYDXI+O/Z2
qeSJH1WkQEUdKZp+eaMbDmvZTuEuMAPNiCpl1DFTyl1m9W/EfKGHfTYkD4ht
zFqV4RF4XJSrbi6EYn/w5VchzFOcamnLRoWosx4k9ErWW+KcQHViPuzKEKDH
7AscXARGcJ45y//I4ddtc9nufO828fCE8w+CqoPA+rfxznZEO3S7ZBk4PfMl
mGlHLqCzXvst5hIlMSGG6cLWayH+5jaCjnMH7GU2kxNkW0EiCHSe67rx+BTe
qIiiU9uwzmlM9BTEjvB1yV2q/FNpOyv67y8lP8FbjY33E4AR3J3hQXBad2+W
x2sKW2jQwd/xSdqJSs5GQRbkeV639RCa9D7G+pV4L8B/GmrrF8GoicgoMoff
rqcws8HnsDmf6XGaAMdplq+4wIi89W1R3KpnKkhR3yuzhklSAB3bbHJ7h0FK
DnGerjEsf+fNyJEDOBJ3VCuFQ3+bM+l+GTjnyv8a1nlGCUjDb6ceQcxEHCtk
6aXcZzxV7apoSGE5dvYmziXKmafU0HgY3NryqnaVima39HxRO1xjEqeqBHXF
TD+82S6WTRwCoQKwJAxS3Dd+IjzdjcEUYz6Q4sTkl5ZgKfa8vAg8ueccUKYg
Z+ls1zdCuiDDXVqNxT4LSSJQlw4++x4ltTDhkL8A05NiPUYcHh/rGgFguY5D
Pt3W6SsAhkXkXq5MpaKObbJnqjofKMaXHEUfBcAEstdv/+1O4AnNgOuA3xns
DZcu/+FDA6CXxNP3LEMX/JA6NTJFt9qJZuCO/yFwJLw17FK8yhC+ixsbzrne
ChZ9LU7qy9IotAijyrN4sr5o419t/MHHD8PjzEBBnk8rBrj3h6jlaVWy69+i
F8NqVPupnqFZzvcSoONoAZy2CNM8PLwtQPXUCfkw/AqkAqICHu+e5vh8bTsf
0HMQ8lqlAbrQ3cvAPoNCcy3QM7+LbPfEltr20jaHQWiXYGPFKVouhdehRZRQ
4mas6eDVI0MQeDH5/ROaRvPxE8mrgRgV7pjcv2chuZyFVUQvVYLPoi6p/scJ
FTeb0vCWtZwuVz0QquKa8DxNaGX279j78IZ741U/m5XsPm3qddkUOVZUn70j
LuXCIuLDPh3scRjwhmHQIWD+LnIMydqK0xeDrmrH81KBm6OKmGN8wgIc4HkP
8U29RT66Og9YSO4eeZvQbhIuOpnv2dyDGft4iib6QjttwAPW8e5tMaGUExuv
3lNeBnzBt7S9hlNbdq3VR/fWyk87DpGeyPIAvvI0mu4lx6vvIPyopZap5gPB
rN1yUlaGluFhAB3PFQW8gE6s4lzUsP3XfDZvyCxthmRLaxRUNwlTNOPmN6VN
qvtosrprlSM0NzWC+XCKHrRa+1pPiHR8Znx6mx2beMwFCKE71pj6TIa1bthe
IInuE28pb2xqFheOVsw7ywAmqa4MgDSmERtE/StEf70pitO4ZqXPM5n79B58
1EpUh7TWpmI7fFKnjrcX3ps6Q62Ny/EMFcJ/yP0BuRfUnoWxELWVHdVbhxn1
FofXUW0HGpfbJjeYPLpgqW6hARFz4nYUTza+6eiwG9NOxpD+LGLg/kOD6Ass
OJ8+dgBqJk56KrOJe6HOv/xWcOROGCuoHIHy3QD1+bySnIcOuoOQAKWI53DO
q2BJViTizymHTSCrX3TBzLjTUSfb+eDcTdajYIVyaNNL32tUe6B8nX/Qf2Zq
ehIEYjBBvkp0OgoGhODBsOjZCr974lFzS4gcfNZy0BFHGYlCAYVEEp15/433
d1xchkk7u1Hq19wH0k/2n6ByCqIVz9/Gc/CSzd0UnhgUO4fX/IWy81qBfXqe
c15QUidPZcRDoerQLqc1u8svucPQ9In0HI0TkupSLE00POS7doKrGDfLMGQq
uGxLLWEAjmgb6JRLiHdXdfUTUhtV/JesaJ/S0TqrZsTHStG3jyMbnSfnYobf
cj5TwT8dgH/G8xLwrxut9DAdL7EdcqAhuXAyUSABiROSpsqKX0l/bcR8Yake
rUm+1TxvFRNscS65eZ9ifLpevUiopsFTh9/e+d97sKTFivcsblilGO+5aOAI
snLI/jqDUsyzB23FWNExGypxqqO98S7dB/0gkRmVP3gkOYZnze2128IamO93
2ZoVWLlQQRWoijYHd5X5eELh4U1Jc7JfvafOHvw3y6WkacWAhFQAVoPceJAt
E+hF1tSMuP4gqDj4Sd1OrmE+l8PoFb2qHsj2esMHDrCFap/V1gtyIxqsFxl/
GElJmIvHCr8ws9BpmASuav66BCyyhGmkX9ze5O/2Oe/2SDAVBLQMtYpo3JmA
53xj2GZKMEZoDS5SaLbSNvSlOf/FjTahsbEItMEcrnXFNIFMCBhcSrL0ij5X
HYyahT3YrTEbLassP8CIw1uIc5uFG92f67pXSeCKMw8WDmPCtLfwdyfxUYEP
zloSSakry4vRO+5fw96LhExv8t/wTb1km5j/H3zfvcYrENu6k8oLcpZ9f55L
tayKAfwbxWgxBJKCp8df8RadArcqgCUSmy6lfgEcYwmF4E+B5Jf8w4h1cyGh
uy0AUBVc0ge6zn8ZVLyJ7U00eoIi/ixdnnLEZag0Tf9e6D4cOdZn+UvUf3NQ
wEjLgVh1wm7Y4rTtXWIIX1/Nw75AtKLsehIoqPGbHtmCwbdIGFQdEF+Vq6p7
YTSlkvbdPHYeAu6WZsNE67XMFgyGKRPCokmkTEtJo0kiIHjlReWhdP0C4jIG
7RnvDC29PUFOB9uckbc05nm0CfAg3kwfoNV84QGrnU0kFyixEcskH6oh9Ksq
5e7qBLG2dC6yh7xURSZZXKbRtKL1HYlwGQgrhqVS0Aneu+Hcf38e+RH1HCtY
Z8HR4fwVMdzHv9EgfXSZ/IIGInXLu/YeEVc85ifdglXjy+ah4D3/FfcUxtqn
VbbfNXgmMui1PnR79ldqaDsjaNhzZ2lGXAM3C0V5ZABLyysVgN8xWRsqvusu
sjS45wuMDMiiSrwnhz0GFwk1LeVBl/Z+g69BUnbFVi+glwHlLAddzbeJCDhK
F9x8N0/qlR3BaI4eoqC6MJ5yu7tsZIFxdM++qCsrQyOuYSaBy0iPKqIDgx1T
kYO5zyLcrsd59P2Qghe7aLGdMptgMtYX4tBKfArARxrgUVdQtS4/Z41+G+RX
+nswEm1xQy8oKkJvJspA/IUpCrvHrmS2UKZiH121LN9HfoDIyUoPdXexhPh0
7xDPOUC8EthK750vA+mLHyAGKLnDIhW/FCdEw3UsSAryH7k5xVaJn9BIU/qZ
R7X+if06UTBrnI7k1/j1up6PIw8pqvgX7HwlGEZxlyNM0DsUxqFzGC7xcbFn
MZKnXADBN8BQEll7NxPnNdeiBXXSylz0yCknXMRG215uIsjMCbL0JR3ZMAX4
U2Mgk+7UkncOCk+JHKcQQ0aOdurVksYCJf38gGNRg17iNuKTafiHpFUM3g3/
HI21MyzvfnVPPU0ThhA5NPaq8NUAuhxbHAySkjipnUaoElEOhx49w++Sdsox
1ZtETBZo2/63ox6nsYPDwHJwvVg5AaYfoHAZauX8gb79PrMTkyJuto3qxbIu
aQUTan9TMG/aHWt6EFhgdWho/2S7iLMV4UxI2OU4hwQCzdI6QuEe9NGigqWK
A5EmyXtkHGaBDKrqI3tKVDYnhC+aMorH61BAWLpnke4PL/56199HkaQhbIoS
hZTc1i2JaWWdr9/qtziuqjenPaT0lpXFnse2F1tsFyK+nRr1tBjCA3B6LQ8S
thrNdy4QznErDvwuXH34lwbjztqwhI5Tx0QlWuj3zqSp2BaMy7wg/WpDsWHC
jDo0iMOV4H6/20p3+X1xONZsmxkb2AnI9UpzMUn14eB1Z6vJiMx/c+YKPuTw
D04+RZ+91UmwtyQiB/M4k2A4gNRD/18OE23KR8ZfgB1F/eJ5/I6h1TeAHDS6
7bR1V84i4rzH7pZ/6yPjnnYctEZbggCJHg2ux6oqSMv1FlCRbLHbkZVqQ8Ro
S8dsSL1UZrAo7JUZEy31Ag/MpjMQ883JPMKfs2PrKPFDrIsIZ6BezvFXP2PU
PECRa3MdIedEAbZKqyi2NkX41R0octO4ECiUJQkF8zk+c1y1R9QYPd3WG+8a
CwyLp3yFthm8SEeLmPVosg8xKgvofFBWgCjhke6mzRQLMxbCMwirZWC3Cea0
aEVuMSrTSx625EIFnroNgApygafNfi1Tx7+lOF+x9+Q6BU8/0XH7xuHe7yt+
Hd7qMMNWVXNG3ad0LMs0KzedBj8nelwL9ah6Ou6ppJm28S680VVtBxBJmB4q
4jrVGAgTDsfDbL11jTxVkbsPsvnNogG7NWa4kM2HHmbeDyxbuBoFhRs38ZWJ
du8zqYbzL2e9s6F+FyqtAMvmGMcmS++ecd1amYW8qYvDIE8KQ17Cs6tdPL/w
EiNBM4VETHCDvZ2PZYsO3moea1xAgq67mlDJ2GKMF3kqaxqlcQy/o2lmKlyI
/1wL376wCbVEduo/QH7sLsWI+8y9qXmDbMPBI3otE0Oa93lxi1SRcTaaRZPi
w8HVB5uoES5z5BJ7EddcelrSYWyfnCr6jFshiBzsfs8H0RascFYyl+ogZAU7
45t9Z2GSX/UIV4HZvdVSF0xpZQPyZj13SMACMjHNqNarGUBeI+NspVNcEYWB
z5Kqh3gR4kFE3f9TYpx+F9GcYErFc5TqIujypz57Wc8GzaafblUHOsNAy9TJ
YKkhNC7ePUU3KXreHsS+pZ3BFKuyWpJRCeq8a6T82rGfOmceBS6/bOyqj576
N22357Kf6l38UsXQFodEoBk3zi/sdkuW/v1d9KuRYTTlnRhqMPEfctGCswFS
gS2e+uKQyzVzWUvs8YX1CN5lZwMWuTDPElzhp7o1/VM1kcr8C9IztDmCN6Ka
iuTjSI+ft5yl5a67/qwl5oULVkVGtZ7rOVbJrS/LnACi/duPl8BBOGwci6qh
CbYOo9oMqaYfyOT1oVNfquZP5XshvI1TlszQLfBugESACJxQvdQLBHBh8pHf
DjfFajojoQovUtFF7B8MdeWbxMMPwDQJ+39E7lCtdLHp8ZToLE4ip+yTecHW
/nWa06OKmaxOXK1nqyBSgoeCaM2pTCLFJ7+ad+3CvrdjKz+/gKRAc4TLRcBL
b4oyolCWqKhcTzAaL9fHcDcwqjcU2sRpEn00aXlSDh2ZulSqm44TaCZMpJo/
30D+IrQSom0OiMrMe+b8uxLGzGEkZAF2d0Imb9w51GOpo4Ozk2PBhuNJpZmx
EAo0MN0cqK+KvhsjfFkctCp+RLbKU94I5okLbBniKIjfKVtm1Xp0rKpnE8+U
Dmne0siY6CcmkGf1pfurnByJB88P8aGF+1i0pMjgHa+xmzNwmkPY01OA3bh8
DjQ3NmAEUiNS679ZAxFePq4r7QiQiDik4N/s4lth8tEvocYzibtfyrB8gSms
UF3BnOHrYljchmYORRgcncn4KphNYMyk+50xUfZruBoMyZ4WF0LSjX4YvEXd
5IXAHtlaQ3BfAV12LOLkXeiH7STRQQGVFzqVw9nXeGGsL0Zm4xYGagJT6pz2
PjVf84PuydXw4xIJtErxty7SDeO1nz8iDrXcB/ye4khShn9cwWHPWPRQDQS/
a1IORlaJWvoCpdIwE7mjU2ND6jEvl6IO06xcbXyZPHbEsepZ1BqcGWQOG3Wr
gk67IXJnPjoW4DHgXZh6uyp7B9yj6/UGCSaqteiUndO0HyIYP9FZAwtcaRzV
PXAR6DBhCiOo6NFOUUNUw456xatFOGv6aj4YqhIscfnMdlwh/ppcor+ixW7C
nfChewCkaUMuuYmoQgv7cO0uh+i5me095p9dknMN1I9d1Xmp2cGyNpkM12AN
Lec28ABLTxjiosskWoHiTsftXRTpffjqsHqIZI6QLGPqk3DNiaxWzcDIzWrD
UN7VhE5ESnli9ipMuzFbszQ/fq8a7GmY7CGsLRYywtOuvHFWMm79RGqB2IT0
wUBKgFC1Cu6RCK6jwSvBZYX3zZtyQE3acTAOVYnDlPuj+YsgxRMC073Hfd2n
GliaMcgC4m9kZgzeWrnTySRAG4zuYeX4AEG2nWc7kPiiOrNTfUtbIvv3K/Ds
tPzmrvCAXh83KfkfVj3PYvaMUh0gwAo+sT2ikqCY38n23pBy+vL/o3ng8pQj
SxYrkfzyaWKDSKdlrnHbwv3dSs/lKfgDZArfy/qxe6q/h9dGsZ2fC1ADBMi3
72jfEokRhBULRxU4tQqcagWVbnt1ZXWxAmr+pXWT4iHmRWaQHp16WCxpeF0q
QA5ydgmklwNBMAmxT6spN7xi/khVDtu3ppKmF6Xzav7BKPNUVST+QcFXQgod
3NxmFEfjlTrurY/C0883+x16YbNw8IIUEeZUOPtcIY5T7KdP9R1Uoe1LTMrJ
z8WZKTzYIsapKLodrh4GWbyCfvf/K17UGQUKcoPhsYJNP4WBdA55tGqJ463r
O4Yp0LURO59OzlrNL/BHoYCw8iX+CWxJ8z9CCI7JSwf04r0FkUfhnwOryc7p
iCYwdiNz0vKdroKmzKE3Aumu4HoHWMrwm09PtvbaG/0BIiyISz3TYXvDA08N
NfsK8Z+LqZlLe0g8VXVdbOQYIylI1GmyLWQRlbcmn1awGQu3NhdS5e697NiM
6IstKEnC6W7mZSfQU9KNb467f1U5I+Wa4uVceSMsWL6NgbOtQ69viZ9tWmM+
dVDbL5N+XMExb7YWPZ3hDYn7FR9cgQO78xHebG5cgn0cO5M/6Zzb80EkmO9W
/cmpm1FI5DzIEs5GhuR/CbeERrfztOvFOdH0kx5YubSsHc6NI4ssj/KXaCrf
RmBvp9j4+lI5aFDEfGV3IphDkDU8poIO3WQjXKFk1Klm1IS7Ajksj4NRzk1k
y47MMn7ubNOi10Kzxr9swCRufgaC3J99eY9rz0LvnNtt0WhO6y7DxYMlHno4
BwCsjeea5UZHqEajQnK8mubpSOxO+/ki4Gx/448v7L6PWWUX/r2TgWqqMYdx
f5JlJBqgdIFEHbAJPDCCuX87OSXjMyPTOEYCuuJxM1WbR9I9GSd7r2HHUk74
Qclv+pj/Bg9+KgHMgbfH5dsVd+4DfWSEMcUwrXsEl6CzyQFvYpFn8J/ze9MD
e7rtNOExu/IGVjJNIQ88lKvEq+Jxw7qHRx8MhYlDfhmsTlb89WgP7B4BMLAN
T0UNp1NelUiC6TlxkWgRTbNvVtwKrBzaa/5HZrqV4KBt4oYT6auJ5qgyBumk
OFcD+rjchRMrHLfX1itINk8us+n3fm7xRo65OjSL2KvOISfwJ2LKbK8Y5oc0
HujS6Oh/9uN/XeTriyaDHJcfYM3j72VTYrw3qzVKFLOyV2oC/zswwSyZ52FZ
dGXcAaEUkJkSz2fnhmnOLHFA/C4jC9F0A41OTe21n/jkmrn4WVsA1kJvlCjL
n7/+JSfiwgsi/px7AAPNJmVejlFc1ua27zOnZIM9F3cEy6xfW2NTwEwcQp7Q
z26cfGD5tbir/UoW1yQfqOc23QmIOM40dg6Kc/mxY5TeLVq5p0dzVqo6Au/a
Nlg5RDsKTxqtvA1c9ellrWA+CdJRX84szcF5scuyv6MUO1yRVkpt/jsLBci8
nU/fkULR2tN8/xkECx4XNhJiN1gM8EH9ucYYcpqHTaTOF8WqAUALeldK2sY7
cs01O4PeN+1aEhGm6RueltNdtjW7WHLcpv2I2lCSut0noC+wJcKlUPHwea6k
B7L341fV+5kBJUbfymE8wPf0qjQ5kOXURtih6MD5MqfRNUZ2h7rQhs6Ctzp5
f42HatIAX8BiBmziWJziv90P+3gzOyIZGL1LsePGJKE9QyFUMHpdoOv3xRLc
uJ2EUqxX8Qaec9lDBRAY95QNXYTdRuwclMYhzxEzrBPCpCHeRxTjStqpqFJb
XVIElgw7lcULZrVkqU0vkxvAKIlsn33Sbxuw58aDEH8MtveDZRJwAxvQoHNb
Eicv5Lg6kjk267hknLW81B1s7RAMkTm2IUI+X73bQpyzkl87Y8vfEqMIJC0W
ERYCp97sSg4YnzH2S/qxUVg0F4fzG+9HSj4vJeoIqf6RhMtnj8tLZfMMIhJ9
UD9PXcJaQXw5uHLZdpvgTqa4AS2Z0GPSK8LTgV4dk9d9s8MN8m8oezTf/gnF
mJexZij4zVFefqPVSoeTtZD67K10ZL1AMRBdfhXUBP5obaLzNs3bu4DqbuSZ
Z4hirwrsrlCMfkxdSp5xJJZ0KGJsqkeML7oWJqnXlrzVeaAC119DFeNJ1bWE
sT997wYGBLfrkKWXiKjbBQDNWRHri7sjFY82mwxhrbHytSaDRzxhatn7cMbq
6P5gpaOk577t3r3xhHJ40X1RIH/fGpBuFVUdDWLyGlY9A9l2kKojkYx2Gyrt
OxJrDNwG294Q9/iitJ7bgd49XUWfS7clYL/sWgNWXxrErUQrvjX8WEJsvFAa
9Jwz6wwvax3dPyfx2IWDq4FpQkBRr9gUp2BbFpu861JQGTZgq7H6VoVVkV40
mjWSb4DkiK0N7D8ZC10/R/RMr0LbBWInd1A1+RWvpTaenHiUSIuCUAP4PjI5
V6JOGL96Hsvm2Jd2OrxIEgc7/3vDkUkZ3ba2YxfhPrDKzzYsZvL4HXyxCP4L
r4w1xyUtLAM6sCb5KNhCfJvBj3m5wy1CzpZn2wn8oxzJP/BlRrrzbncuBiQP
12D009A9gBrGRc6bUqlMtb7HHVxK+uoZV+tj9eai6V5ZPOlV0yrXV65AUYRn
veLt6uSKqupTtE3rjIoyA4dFz6NiKn2yAACGQYZ6mo2oZj6HKKXkoFb9fo14
Uk3k0ncMCY/385/Ad1z4WdixLVc986ZWosCMNoSPwdFnWP3dgbhadBTObc6K
Q6qSpMm1CfgtsTybODqmHAwqO1m3vll8a/3oe6tW1eKAYsnQzmwZNEjPrm5W
9Bjdl1jVD6BBWwDhFsEQLRkDNNPqN2vzMu5CjRSG4rxGLFRtGhwTQ4TRIcbT
p/ZrgrOeWsVeX/0bnCmduLdcawIiSNwhhKR8EAFHZSD0/TB2XThDMAi3pglz
DNkUWg0Z3TWui7ZwwLDHfYzKA5SflDVEw/kSzQo+XcQEnZqPvDaAcbiNzptL
kjPl2iuS1N/XitQBP+bNDSntsgVQjEzgojMdzZkkGnwNFrhgOQOfwukDUY8x
7TZkPqFCy9Qdz+k8RNEwYA42iIWoo663tHf5sSe95ssLpfG1xHH22Fb+OTXE
8kSpqU9AtTMK/sEAa+o4CeFEH/S7S1/0sGwg/HPp7ZTk3fn3qkVFay7rgRtd
rlBzFrX2zib41upl/rUNR18rR56U9yqSmP6sg6RrcKVyuMvWR7dbTHcgwaYC
YmJlXpp9rNX/DuKNhHCpPCYM55tFk3oaswI026hMYFrKQOr9JMY5cPpqRSFD
X5YO8on+H00yZxuRaiEVYvucZxqCL6d8/IqWssPGiTJ1UX1BLegI0RNYHm7V
JsQbo80eGC3EvwJoa7bakd345XWMj2990C3DkeAz1wfK/EC0N7aUbOMBizZm
ibiIjqNvE6MKn9RxsEOo8X9sArjgvG6RH7/kMf9ugYXKXwv20AO7eGJfy3ZH
t+yPP+PuViLj/jpqW2z853qr8/eJ/XPSha6EVCj24+TiC2qBLGixzINY2g6Y
9cLCB0A2tvodIy34POZx9wX/0nAbEnoZGPdBCG5pA7Tm3o7A+5wavUnd/tTu
fnJOEatjLVEWnFpfpdpFqMh1fTCNZzeBkz/TFnEgtBMN8Im2tmV8QvV23yWi
zy4VtTM6m2iPporimFkBLA6gvLkPN0EaOC0I1jbrP8+BMhh5r8d1VLXhdkgI
7tNq/GXkSMaRz3yPpqcXCgDE/QK+NXYcL1r3gBz3pjVGDBKpQGJl96THd1eF
/F96PGPQsU76z4Yolb2VbYtP2KjZxdpXpmbVdTSOtAhlHj20qxfKRjiZft3/
mPYtVEl2BnZoHoWTxhURWBf6gXdzXZqP0lg+a2/cIvFivFeBnhhNzEFILNgK
h/P+gQy+FUzt8Sv4pl8qxTl6UXvQereru5Ag0TDir/79SPWOL4/CfIVFR9gc
gXIlN10dmNv9lvgYnm4zxQ9m7fjydOGD6Gqlcr89kSJf5tjChmcDWYdV2+KA
Io54gTFQJ+lF1UFy/wozecEl2VPFwP28pz0mpb0mRgQ5uWw3wFeYhIAxqlLR
tVA6NOzT8yuw+EfW6N8/QPb0n2N5UuDSFAaQHu3pxmlGkFAHJxIquu7FpWFZ
5SSxdhNcgIguXTF/tYimrk0YUpg+7+Ktl5tO14R2nxeCDIbdbk+NjZb/zwiu
WIEOEq2XRrunr+CsVND4QpwhIJKdDuXZqEgtdS9kRLBwgmPprTnKPHJTgp9F
XSEPU0QFQx8n2R6oAw+ot6ZfkRVIV0+S8PrFjAIs7O69yTTjAQ0wua7/5wjk
mShohfYuNYd3UOCZDs1KYM8kE76AAtq5Lio0F/Gl36xh16js/9gqd5jBf0RI
exE1HkcdW3GL9Kx36XkOKvwRDYczPMcGvoLl8jvISFISQC8y2udH9nu/cekb
pmjMex85dxn6FFCxoCqfShFy3e+LPDUC2h+t8x+Kp3UMCfJCc6+g2LaIVvSu
NeQYso0AQhHhXg+6XBndKkB0fXeH9LF7VQx0+W6IYlIu1FrPuy0koBn3Aq8m
nUD8GzuhAkYFFgu25xUbFBJl5HbpjbZvTPJWnH8bQJzOkxMWotk/639eU5f4
LMpWjVExbLhqc3EI+QFWod4pgfAwC0pn1T0LzuF51oPWG+jeNihmqYfWc/6L
1QKJNa8QDLwMdbrAGt+9ERDvP8UVlM1ESODMEE3FLZ92Fd1BZ9BcwpgH8qSM
bQkLA65qPsm/3B6usnT6g4FYtg4wNQ0t3f562iAV6aU0Y1IL2qgp5v6j/vuB
kMpXWKlD3KXrEk1snxmwPyosWAOaoZ7UPhJpkdASfacquzSeNN1gwbzJpwMo
ipmPZmBb5RserIL6hwdsyD9NtMYQXGAPuovJr8rELz0TVbninTP2SP7EEpy0
XSUu1bDzit3fHQpcxqYVpMLdTGSwKuL9lt787Oo1vfyl3QaMXumgHttSxFyK
pn2/KeNzICRle5f2Jbd0xb35FP1sTLPHX2/OfnoT8vNG3qzkw8tLCtA680M/
CAJ4ubVSBkDRWmMmmABR6ift4okTLvc+F1jep3+LpxxL6DkY0uWUBLp0Zmuy
NKoAm0Pqc89LcfzW0zZRbl6PXDQ0ImevYhwbLPaLBT1KkqOBgQ4s0mZNwb0y
1aSLWCfoDcCcA/VEomapgqex+rbv05CJ1B9R0nLozVHrezlJAz92/blGfo6R
VrmRetl1/H3m60ZHuHR9RdLOgjutBNfVOh1Gh/YpGtnXjMLjT1zL3eypcpUX
BOTb5I2x4U13upCTtCRSIEchymgS9I0JoKL1wN/4IRapnjU+rlOX4+xeiP8d
bRVB420srF+dbihCY5SDQAPEFJtl86lbHsaBQk8fV6vQgVrwRmk4GJmdIReE
xpExmzfe5tCTdTWoVJjCv7xpIZRmJCidreY0z4GJmYidA6JBHQT65fJ1PfdT
lK8K0kT6I1w0wosYstk4A9qxaAxuV0xczGqVCNWeirckmUcnN+6DxYaGiB8p
LUYBBq89/KH/ugyEFqXwbTYAijbTXVznRTPeT5/EZMQ0MqbEcGYC4B5tTqn0
Z/+HPFMNE/nghOyvJBHGcM0sHHM9X/EAM8UQZlRopoAFE31kdjCTllaXYy8P
Idqf8PTE6OwyFGPCSzAq3aKYQ66URsHChxRoE5uPEFRQedfE6uMIHIfeVSpb
mrkO9ue1Va2mE7Ql6aRGkny82J7jFYA0RM96NPO2F3yzpakZhPYw6SvMXmsC
FkucK5RAW9uJIgktK0UoMy+Scb3XMWY72eJ3Nw78NKac6GmXy0MPR3UihrAJ
wC7TznI+cnKWO6lShN7TYDdcp/aTjPPz3YQUysdErx9BA0VljqgrEJpx0XhE
xJfikybl0RmIM3b7b0tTKa6iMvbwXC7kZ8JWWWppLJzCUWe3JJZJmV8/Ja0S
9OFNiYR3LpXYWhWBTFagMJw3+KBN7QrOJm5sDy8Wm0hVSCJJJsbuhDaL2vmg
gmty4HxY6OcbkZDm3lZEZVmSWY84TqmoOnFLBevC6XD+m8F0TdMqi1dfuhTs
mVQBJq8MsbjeTnVReqwq0Mi9IO5KLgEEo7DdgnjCGudENO0dCn/uEHxxQdDU
WE46Ph/wpyTh6PU52tzqdx0NpDYNhUrGEspN3onOCbrDB80mZ3A/s2y5eQaI
no6MNpI+G/qPxwIii7cBLCVk7ZjC438iTuxB+IjJwPXTGHBkdYWAeveViANV
IeorwaUdoSzGgf7c0mMkHBJTU/NbEv7Ks/pTZPbOt9jdZIicHxyShEUgk7K3
Dp30x2tMu1v4pZSelg1oXXiAO/hPJT37McZLxqtExZ8HDU0jgSkSEXz5xPNi
uxWQieyAeGSzlY5OV51/bm71175B9RaaN0vrNdMPEO1mfjgLEyzEDft3bVGm
c/9U/2mAfn4/SK7D0/wjM75OYwk9IOM1MgarvlkJLMgYLGPJI8CsFRY7Yqo7
LxTl4zVrN6lj5hg9xy92mi1JDsPOjOYeo1R2cjW0xeRX5yo9QgbQKgIEgf8/
XXjcS82slzkrylreM5ALagB40IwBilo47izEz63fne78xoEp5uv3D1YgNE8U
66/8Qs69cMVQGemc7ZPILGrwV1WMz5oDmtbzut4PY+q32dQHuSaLWmbABq7J
8ObpfKxPc3UeZRyU1GuWHD6Mx3Alj6B0BWDQ9zR1XjQyQoG21MaTraQUgJOE
8kQi8Umd9w3XbnyPwBSvHP+ht8w7kSKUZLVgPKDDQvWGaR9TdDRk6MbPji6J
DHA31ICrqW7hD3nQGkwPEUZ6wDhQigpAxtvQVpDShKOWHbQ+ioKulRuIJTe3
csb/XICSoqgEKJD6BGJlBQ47YYnXH9fSYndVl2uNHxNbQmffuO5U/KcPCzlk
Azkix19VPVkxeCYOsuM6xgHOqrFYAJUO8Jdt+oQtipcDeBw2dD0O4coyubva
kXHCg6U6rWH35+eNohtek+FoUgGVnRa8tSHuPIKfX24/ZRbyrv+4TvljvJ4P
t0QE9JdniVaykwf82f3/l6S4PbUxD38j7OE/PTfAJNDFAOk92O7VQS1biPXW
xx3LCeFSRVoJgwJlGwjZWbCYv483KjGy5yThMl5EHYHoyVa+0d/602fzoHAm
KmMu2jx4imDDWXxu6h7zYFHS/Ois0Z1ALnMdjgjYdWhlZBXFpG0Rx7Yd3ZJF
711RaSzMKO8JwyW8lF2xB2Mrr38SFMOiEqVLXyDQOxPFc7Mu5g61sgJlb70n
SVJf805MfR4uvlzXlnRfBQYylfeQUTI/6Bzh8Ct0bZ5TGq7h+4zzBlc93cl5
oD9NBR4WemIdhiZ1ybGc1iQup1wC0I5GBuZu1nTQKwYTvwoqFYPN3fTr/NGn
L9wSQ+sUlU0iK41TzuQCvufM2UBAsD5+CNcbK2cAD+nng3jM/ejqmaWUqO1U
czRBBIDANVe/Xvnu+uILg5H9by0DO3P+tAee6WULgfDJXPRdu8cdbJV93UyV
mmSBF5bzwtuBKl5G9BmUvwf4bPYuGrvADWkjuae7OGTOWiQG7xPKLxjn2l9S
sp7JUVbuIaZz9HPIePnRx+ijYM05Z2CX3wxi6l1usUfvnnxgWIaKkVr1UiAL
6rD9dt+oHzIQQ80+hJI0T2NkZf8nKiLJFVumeL4HnAIcXqsiV0pE58ga08dx
O+/7+dcoZmh5gL0TgCFq4BFow8nQVv5m/zWTSfSl7h4EUP/+QIFGhnTxQmIS
0Nvr1iZa4rW/3zmp0m+T5gq8Jpc5YQbg5W4oNqOTTgyUtSG9PWdKgMzT531z
+sSWE/0ih7j9+MXGi5R7TQHPL0w3uhy3tlK10xWD4uF8FiYojNngzEbYLJZ4
qteVkkh+xEW6mdSSCJEPGl9yTdTfqIfoNBkBGu1zDBxthJmnoRMRhafeG2Au
vi8neUTypMRVM5bmp/VaVaQGKFakyDKu8yo9PBmLkj2byV5a9nk41bh2SahC
gfroY+L+gXbZCw4t0IAkDEBmQfgZPEgJau6278MoRDHo8fBr0jjxFab0iEN1
dcSbIHwcx+aF3dC4Malk0y8Ne6Nr2JfbOvo0671VcgmegbBsAE7pXzDXwtw5
r4Dhgx44A0dM2S5EQMI/kby++zswxF4Mcf1pau67L5m8yHyEeB7H2tTmpi69
GV4/hppwVHOH8sioPuuTogr1a9LxY8uFyMKle3KOOoR/TwVnDDWlWpzpK+Bk
p1BE1LcoKpaf9IMSd5LrpkGdyPXZwcObMrFKo5Qq2a8Z7aIwHgtBuOEbr3mk
vKg/SsRHK0oqwL+psoC8EQ55nfjTuZK9DXiZBUXXOGX0Xse15XLmtKK1HaJf
H1s82/Soj93yot/j4i5vCYbo/8uF5HvJ5rdJUSaN2E9zGudBr+3hTsIuYm7B
pc3cRO16JjpQwOuq3HGeU4p6gxX/b55Fd16P5MIP5x+IFIhRk4fk4Ttua4iZ
8DkIsSs11I3qpFqCEu2ol1OIoQYHRLDYygED2wSK+H1tfLelc7bu2U9dzgiF
wHXhGYxegzSVCltcH4pCprjU9vhP2DzrNUlWCS2m3f16Ysde2VXQL4AdN2oq
5IXNnASn36kSvs/6+M1+Iu/Qe7kOfg60/lly2r3Xi3gNT1rW3v5h06HvJ78f
Zm40omRnwTNnJksmOqkkEEpGxi4n8dDXQDK7eJWjhyGh2Po0MaOmO+KGO1RU
XtwxNr89eBJFZm9qwZk8QlHwyM9ZPRWi+XMt5S7mEfpa+GhyBZkYd7ukkjdz
XofxPGRUfQxhJuaRARN2PuAZEYdjdwEzmnebhspH9W2K8J0HQQAOCrYrLcTg
LXSm/wnhh0zpzWxQM41Yogqy4ivKGcZtMP3SNpL3VlADwRtzOG20UvI7pyUk
EzIT8jNnF/JODAO3mvLMIsKBtQQnSZm99GmSyxyL5T9ju/H8slHCIrTmrCWB
3lbS5AYpxqu5UZA7TgD10+bpL0NZfnM5+2CLBxvAbZqeRS4LkvPY8S2l2LWP
DS5CQpKckzLRVClS5TXpttMombgz+kReltwzik5m1J9+RAlCaKfQomoHWMzS
6Zwbkf8kGd+76vnm+md6qy/H2WU7dPUpyLcnfcUcK0JOJ1OH6jizvjxLKI2A
N1K20ocjsuDEaSkGHoC0Z8BcWZk04SO52FZJvm/1rsnpSFdwmEpsrX/ZmpYM
nPK7qE/mmurMVJRjw0OBVYeyjtjFNrq4R+Vbpc/NCqxtH3N5F7WfvqNkfBWL
2OxBEk3p5YeOidpa9dBva/Z7YCXamh27CWfYvlcYrtB9QHCCHYbWYpmQAo6Y
ys5RE6KVrivEXvUyxejMJMalV46631B8kZrnhZP1THPhzQMShJtE30Sx6n9X
ubEy4r7lOBHzUAXX0mkhXJlbIJhMiSuF1fiRUOhUK8hd+UUEHzb+dkaT2OsR
BJP0CWS4kN1EFbPduq7mFfw+eW5tCYYyPXQqr3uwoMCdWD1aEWBkk0MvX5Mm
RyWd9dPmSZfHTzyTGqD/R12SFk2Nniaomz8kbgTJXqiL12EsDrtHCYmstUw1
jm9s2jTY9CpzXN0vTPHCaQn9MYHPELdJrMQkPVc16YKOjETgR6w1FGAJY1vb
F+gX4Yfy1zxVipLiaAbi1/28ObF5i9OWxSoxR4DghA8diU7yc9yU/grahQ8e
BpV8MuO7WpoFGw9qd815p/KvLkOblcyQ/CUMpgFSu54bYfGRkqACFwb6SnWh
WxwGh1KGDwBauGmCqbPu56S9mAVOJl9CoKVUt1tSpu+2kVTPFxu2v3Lyq68K
dORdect7wmj4a5HN3LHABvgd1niPFiQ8llfQK+wAWBwLwzJv5/Okm0Sqecpk
RLXJ6DVxfuXmDPflUvU+DhCyYFXvFi30QH/SKTM2U2lP8m3bzSppx2zDXd/C
BT5Niu4+sOxJj6eQRGDqTh/x1+P71mzd3rftbMQWpiM/+9nYZZ1eAbWqSveJ
kq8stxHhLIuZ01wVw24XBeRXXySh+/qJsT1A0Kk6+fWE3uUpB+8Lxmkid4aw
yf9LZgZmX/SoF9avW21iXGrCnDAXUXab0xrK0sqGbROiRNHtAsXYF8Tly91V
uMiHFotwxDRHzrncyB8XT6qZnr2yur6Co/lhbQCo1n5FmI/96mIik5sdCN/g
PjhIUg0RAIl5o9qbLDIoFHl5IfiL5dxbWPUsGKLVMmW2h44dZynhL4F8TTdb
GMh1x3csGDzp73vCliHFDQGSFG3U52MCkO31WgDJDMRTVBDRrtIsNUtMC5Ky
AMYOdwgaU/BCo5JKwwjeGBMw4Vb3Zoz+4rak6tl/pI2EfgGtkQWhjUkj+OUU
hbUxX5laAZgl2U039RFp9xg5vU7SkM8aNaAs9mFeJPoWzge4gsWtCWYYwApU
LF39gUkU7qgn/0Wk0rJ4F3vNLK60VCvfb7fFRNBnDb0neKSdEJiljsOiPByu
QdtynRYPQrqyZWLPkOKzs1bAZBTTHMG3xWGQClEDh3joZUA4UM1ypjgfiVXp
uKAZyWcKORoe83yeNhVRiuD3y0MiCSpRSXYp+/2Y8n5xVNsn+HjquSahCkOC
S+DsISfNHSLh9Adgsje23dp53xCkJK55LnwjWuSjtZMwGwiHKiVc26rSGCT0
lbr04VuiuIxWm5rhaWTDR4Hq6/ER2+NCvKhG4q9215KSYwYPE6mwNkZUyADL
+EnvzIN/haxdq0+Eri5ACSmCCFvi7TcwmDyC6nauEZmGiLhRux/iTOF+ybTy
HEb+qOkFjg+YKxrrkMQmU/14dR1sn72GSOY5eWg0IBhjT2lqfLMkmIMjOo3A
JcrxuPhpNU3yKjsOw8w9kNFCeUR/eJtzpB+M6DfH6T5ZceNLF5jDktgU1Y1K
vkv+dNuE6OKT1PwBQOywdshRkVpIr3bPq/Ro78Ecd6LYNBJChvVsO91mJVHB
RGc/fUQ7UodwPAiOE6oAmjCOkLo9tSVpTN/HpzwQ4v6O7B/b7EjoN2p/QDgt
2QWf6EROQrpksy3LBpmOn3Jzhr6vfdTkpkZ7nX8xGmWvK+7JAgSCoyz0W/AO
gwyW0zlgG28pwemS5e61DZc6Ipqrirkbl3BxRAvxS1xEx3ECqgxBK+L3P1zi
Kj4N8p6yTs9IVhB+9nqoMoaNCi2440QTU7eH0mxO38gHrJ3FhqxIXDey1X07
u+Y0OyOUTxL0p81DAy49ztJCmGC/7ai5dydgSfXRE7rGNzC7aQO9hee8MA3C
MdGCpjqDIW0C

`pragma protect end_protected
