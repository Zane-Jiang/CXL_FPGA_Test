// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
GaLXsiY1syZR/a9bBFTdqm9abgFZgHXmq73AA0lMhdpeW55NRraf+PHYWrR/xDyd
RznG6h5vCuGu1cyb9v7RtOPtp7siCJVzu2ITnlRD7ah206DmSDM7fY6VRGyb9UnD
iO9OI5S7nyy0ITKSyHvdTKcSmOxMLZrLdsSbl2pU/ko=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8640 )
`pragma protect data_block
t6lu8/AZdHzmRQWTEpevgfCgXcj81rxjfxwm7ZTur6+8DNfdqCPGbrk+g8VOfvkz
SwC2toHBnbq85QK/tDJTGBfYH28JI/s80xV28pd+cmxV0/vywOssg920BS1yzgn2
XMQZylQRsPLNBRGBZRFtKTr8ULbbjPE8nFB1dHM7c4jdoey9OcIHjXmiWqTVHgUP
f11sNWHy5BVN6dnGyd/o89zlxCQBP7RxUVUPpL7sfFRfgke9FVe9kM382baRMXRY
Vd8dX+qP11MhOHYR5XcyX61YRSb5NZWr3Wz7gB8jEHF56CD5FBAE7J22YM+QxAvh
YEdSQE3Cwkdk95R5+cAGcabKYLWtLSfJUJj3GoZvjc5STKA5xZ7pdOd+Qf4CjNDg
tGHSzVZ99mTbfaaL78oAwNZHP8c1S/+PG/rLrcjYBehYgncNG2L/8EWlnTLR3XvC
eLa7rTsLgzEWVJhvrH43XtBYcEDDK521jUkJ85ETA9BTs8zOWfU3hGni/H0sAo97
nmrcuDgp1Pkhf30HmzMhJuWkqKXPUp356Kr0kW0avc0ntw0yFXbrlpUolnArYd7Z
wewz6j05+4mqmkPs+ZiDC4B5wZBQYKrCfHY2TUpWjgD3Z9HIuxtR/fWOqbC2uz1z
g4YjUBqJTFIPWmI9akpYJy6e6u/k4OXuhCU+BRZJoCMmTWY3cdNgRE7p0m7KqBlY
IiZDvIb0f1DOKQFWKykxzl6X5Iv9HLi3up1CiMKm0sgwQYnC38/u+/nnzpMfgHG1
0+BB9/XBXfFbOS/D/39R9tiIDOty0v9e2eOk7nGeebnytx5x1PTuueg6leQmfVkQ
JG19PHipge8BwjQy3HV0+XnHADm8JXGelXgjp+xwdRUWGMKgixr/HSv0hy6nxRx3
7C9E9t7L4V1n6cbJqSWexhkG6zr38sCQ2crnlRNk3g0tWAv2OM2pEJvjofQyOhpd
ymBCPRoNNR7Wa09acMR5d8pUWdkybvAvuennEdUZ7qRgL22qF80fZV01She/5KKp
/3xjv3kWEV2cEskQoldw8urtjEA2SWJ49qX4uoDEH2fUmPCsutWDJlmIhyDSfJbr
RwbeIB9G3tPsgZb7xC+9cBXjNu0oQtMERUjNg9SHAGQ3yQ3utQoLY6PnWrNNIdYh
B0gHOJxITjeNHmGLt1PxIb1jZ0/jPJ7cL8ZBC/l0xiEeujmmyMRWQJpGJEe9LQ5f
ZEAwlUGKQx8CKtgNSAO0z9rnHOuoQ/q4NKH+eIrjo+3snC0L7dTcWTpPglRYNqig
QuQZMPpeYvZ9vS61RLsYvzD16HiC/4sJ6SC3mK1CtvUU7PShHw5rlrCLv2CXodOD
V1Py5OL69zxtbKt/6zMfF7+GMlNA5M00iRqGpJKAwWsCFPemdltVofcifJzWcZu4
CWcc0SvyFW3VesSRTHBlweo7vatGNKZ5OlRHEExNLEeqs+oMhQyuBfrKtslpmqG+
VRFyQTcsFritclUUCiK608VM/mJ2C182NKaVbaqzF9u+vcizF9cQW8lPm/jZu3Ao
cm6wdUdOKszhAmlfNykjm4iiwg0N6E1e/2Aszct21ufVIzHd/Q06IIdj26+Q8Zgi
1QVZvwTrOiq2zT6lWUCgj/61Yrt9J2Fn6VNXrwwalmxIoyYpwHbQgsgLXphmA/ij
98S82A8Q7o4Is9zd7zazuGfd/F41cJcHC/s19LatOUySenmTZJLlBNM50U0lhOOc
cSjKZziZAXE1zNv4z4VqcA1vUhlL8CrYwCYVtHOyaaLikRxr7pwnpbvwRIUbpWVQ
aUEYOnMSJFW4eCds5pvle2DYCjj7slYFH7aQQ0NDHSd0VIxnkKXKOlb059Not011
+APyPC0Z9rgzVIi54aGZr8XKIiPWOYkzWxQ8/Ajam44BkUnjCilRoiA0bwqyq7ue
DZtngZA9ZG/Q9QW4wYeN74sFgVqGCtYUwh3lbuIuyxY7KtqGlao0CQQBkmdrYBOb
lZZT/wDNMi0r76NTUO1wJEMKccwmOJtkDykp1ntvhga2OBGVwbz+NIxEJdQs6xxX
ZH3GjLBdsbv+73LXd57G7zsD/CocZNVmuSRxTj07ww4SKg5T8dvgIJBwOkUabaVj
H5Q3JkvepbeL0kWy63EBHobbNB4wYAI5rLEUecl/M3YWeHOXucfR9LF2cgzYYtqX
wiFlREjgKxv7wLE5KYfm17QL0iZGnJmKjcWI+2W0F+QWClQvNVGwbqQJLum7nucA
+fuvndLNbVDuZDlP+KFdXMnsoVN1OOlPWjnekmWsuGKzYdNRvpPF9tDUpUDEGI5e
W7s9JpfjGR2Nhl/a1fW5DHHeyo7gJJVJAYUHUL8MGlGom5cxk75Jv2acDXtZkRUi
6afUiZ2TEwPlpyg4qL35Uut8YnJ1mc6xlo5ZyKsAZiVvPWUV/CsxhuIDbbjW00Z1
c01axCN44M3FlK3NJnIs+ZRKj4DsBcl9yfv7tnWSfx7k+VVGxVQ81p1O1W4kUX93
6n2I5Ll+cE+DYQQP2RhUuGbYSY4h0tQm48le1tCGtdjDJacl+e4KPLTQzmjmFwnI
x3e4TuBMd/UG8+s6cQm030Ctv8zOadttjiGopkwwaBl69yQVhuKQiqGUhyTI5cdm
55C96iVwDErjrR1FyXz0Jr1h8/9jvMvij4kr758MmgneCPsU81oicQUKwimjDdm6
PjQy+NZXHrRxFelVeDb1YbBYMAzjipCH5f44wIo1Nfv71aXHOlMlvcsPcAmoHpoI
+GlErJKE9hNcjXCftMPDx0xQH5bJ3JiZJ/QUkaCg/dy0X2eA17gthd8srlQzgsrV
F5H7Un6KXVN/kOQN9QM2cZaBqnojT/G/DMD8VTwbGn9pNkWYcZEtoa01AeaFsQOh
lCPrPYtJl8jUrJH+cpcw0omb9HIPbaiqyU2sBdGBmF5l0sIfY9wW+D64iFr2W6RQ
06YCmtDNq3GyvXiw8QH1np/6CWs8ILl2ia7caHF01FgJAXEHxsDHm9gZBP/tl73J
ByS8Kyu1F5VESYXdYJCUr8LQOPmiOtjtOGJI7njjf7bBLnUT6kh2SE2Gk609JvZQ
PMg/I6WeCW7ywerAirv2pzYeL+yc11XRnEe0qMaWhh+6WFmIvbu0+nXkf9lDp6z9
A8azEdiuK1CCcKvhqgP46C+wtOeg9+qEdhkla+BgXEoqaUAxSvwbSG6ROx9PfW90
ldid4WXo6NbanlRCIMovhBZUhoviO+02YV9iu6tkgtl9qdcekVkMT/wPzxM6xhQj
Cv9mk7sE5LwhdMGxhKup4V+xrKkpOTmV7bB+MyaUWX9gTxZGjY77N983LGf0YOT5
0Acl/rwAXSwdbDx5kQUgPSP+Aw5lIt7DTP+TB35+NGG5tocw/6rH8sLZ3NCx3puR
avoXd2eOrYqdZoZFaYT9saeHHYp57k4UXdLvji+68VwsEcj47nJjY5aiUyMZZKqz
x7JUIVJSJ5VibZmqeYNod04Mr0rGKW2GOi0FpHTa5BHn8waF1GdTYSi8Uo8yqxGM
bZaz+WR6aEgKZrd47IUGWaF8uzSHG1ewlUSAN7KaenTprUj9tePrmSWL//gSeCDh
VzT7fASwGTg5H3Un4qoY8Id54xWIpKfJmfBaroPPa/F5iEHSpailZi9gPsboLzgH
Tfsq90QcVKkCobqbcYj/ktAVxQK0mm4SaKznqIaSbWlOFzyF3TkH1hkA8ETtaX3C
4K4MSFzqyIWbUezT0Dd3aavX+cUALH2ilvBP456JSjoY55qg5C6EVrvPRXB7lyJR
FgqOz/LbLMjbCsLTjcaXCNmhykM0pRjGYtAkfHOzyaOZVgyEi5oKMdRbK3CjRwzq
ZxURoxDK3dWtn1bVskZevmtSIbaoU8QJrB7mfktXzm9HECMhvlSAQPdTKXHq05I8
0Tr1EKyZh6NIYH6GdscyBEBm9AOuKPE/Y4pAQFkYGbX1YQ/BUO8tlM0y2XVo4JqE
lDK3Ck2kYebeqk2JSPbucS96leUgXAJdQJXgR/QvMpe+Nil925X0cZGCvN3NZBht
mAF98FXXina9wMRMU+2EmqBrXQ0eg20AmRJVDoDpbTbYbQieHK0yXp95i6W/6GUv
KHKunGWQ3hMYFFAxxAk9upcMp1EzoBNx9aMd7LxTQVSPXvcVl2za00NFHMIoB34q
TCJByPjuPm7qfEwnjtweRx8hRt/HVw1yc6Uyh8UeHQScuyTJW6CIkySL0KBpcdHM
uuatv23spBg0g9I4QGVqcV9sZqk2/Y8kdZSRXU9fbpB9n9MfJ8gCeuHXqKv3rxjK
DmzLFiy/TV6u1QDJ5Llo0aXMNwlTLCvCk0nfDnftF/JrdQv5AuGW/wqV9zzyRd1o
T6MGRZA16UCUvaDB8eWFNo5o3p/P1B6XL7Dvddtf2tgNt8dcy0Ghsz/j5fwQmMN6
qMIU7NSaxW4Nwba2rVmBu2AbudWTqC462ZS3UeRSV9l2aegLr4Ec3enzkrL5Hb2A
92nJvwRcUI3Or+xLQDR2xsmH0qjSx2n9dvHNWs2n1GcdpSt7NX9trlrCXYKvrcDF
RQ6+M2G9rfJ/Bm7/1g6iJ+bipo5rP/WzCHYD7b2pzWNrfluu9mTL7O6NtSG25epd
KK1Hf3DT/AhhG8E3onzO3tQu+tnk9E94wTy2cbevk3TNNFux4CXILCSieRz/KQgs
whxO+L9T6jHjU1k7PPXhZ2rFWEcdRM1EbLvt6VcrgtzWitXs9f8QVn/L8DHWbyWR
rBRnfNi7s7g+eFVWUOC3PuldDGYPgwIr7ZeS4UEORW/2A35lnLUvE60amEuCJD/3
gJ5IQ3Dd3QsG9d+033xQV2HXlH+BdHKESgsYyFYZqYTRk/nBgAVIhKR1LXf91Pwl
cL/T7bF5oTmNM6ioMbfkdEiagZ9c9/SEiw6z8CRE466zUmGWbDahS4cvaQc7L92N
R9s0E/wsQKrOHNYRufjPhtRr038gOwK0uZ48G3lW6YWU74BKP80mza2VjNq2XhlF
Ubs9iJoLBt69NylIvA91lxVL1yPXAoaXGOoLZYOYagbg4IUeEOpiOlEQT23X1I6Q
gbUGR/ipa6VQOA6TDpHu2Y5XKpvkofsv5bmHozCbv+GjhohF9e3hj9oVrAk8Ah+K
Oy7yOP2gsbKoM9vks3d37jxr983tHKeDmfR8rHxtD2wzHG6TBQG/9NFOVbu9VQIM
YRQ3B6WlQN8DG0FEuQu1rSGfB5b4qp7eSvjHv86s70WQpuTxvex1v8ochBdKN9er
76e4jy3pkHlPFLaPpWtVf2NAZccaytHclxtocEPpL+P4Zsrqh+OwzEF1HEMkVjdN
FLxo2rkHNOgfUY3ayAw3ft7drR2oXqRBQR2dEULvbWAiJBlcgOKNqX5UisVRysAe
1rHy7WCXBftkqGbJ3gRPOj3nkN/tfrCMuBvsAAQNp5W7wFySxaEHhE9f4oj8VCYU
LjV2li0kORqd2MLQ6pfv/z1fxzDtik+o3RRzP2KPTaZVIefFS4DCAlH61Tv52Xd+
FZRx5ikukCZkx6K9svxOsygurtFMO5Tc/MF1IT0m+AoC/bh5lXJ3YsteB6if+KOK
XJFPfmzwnXfxW+5ZOASE4CKE1kfHIXVDTtbB+u3fcY8P1HLb4pd4XLVwUNmXScIb
WyVJ+hQbP3SW1eJvpxXwSFktvzy25KIMseeOonSMmuPzSxfABDLSDFR4U9f322nU
oAgUdVeNJTx3pUHgY9jrraPIPKW6SnrGbi/fqAep3RDMToObR+3Rt470GNExXwYK
mnZMRTg0rDgu36IGsxHy8XEBqm0ygfJIL+/Pnqw9SJbd5+CJ9MeeJTA4gUJxJsjt
jr+Jn7wJoMfJH+nl6Gu/YOLMR0Y55ORxy03KeGFgL8/1uafhBmYSXkg1+m9s5LB6
i4fbtTOuGvT3Z8+oHI9RWw5W6hBfEPvpuHjh3daHa4VV7pCThNphthkhmQ9XpxRE
zMS6sum89InMsnnmWt2/WN8ygHmZ2BfMhX8XOAfHpZmM5v1Q8/IWcXDh+GSEceDY
soMaGvOeCbGegfRxjghtOPQZ7o82nFXHnnAS0Z/8OFmqID5TgcK08eI6vL1DmE+W
dRLkMPGSrKZxPRomBhLydrLuGJ5IKUgPneAs4iVvjYPfp7rkhyrez7hObDDHprAY
HYIJbCYLLL7YIgIhJkkhvdFudoSVBkF8V/Ad8tbrsvWLi01VaYiZTVssOCkrkL/Q
IWk0hue6fe0BoeL9I02lV+7yWRVZyLqgx90kMYvt1LmI505kMoGzzKHvV7wUX4U5
F9R+YNosDv+rZ8YsExmoVXsCAkKT+kdVIUferDp+4jjRdI8RJVzF35peiPfNrH2s
jbCeUXxUIlglxHN5/rhnoTN4VzKGtZcp9c1hT88yJUgkY7YvpEvzv+dgxpu0saGo
pc524SexmgfCl+ClK3Gb4RaanrFnfC9IgsGN+JCHUrhRKQcYd/ImNlZwbvmDZOFV
AdTZnvQOsMuM7xWj2ve5v+ZQxCUlZQDVDA2C2CGM5Gfwh/DBnGmV+d784GwO3Nj0
fKONj0Q9/HHYoeGifiGhJ+/5TiRW/o+CD8okngGKBSMjen4IHdv9dqcusORnqhHG
twCjsjyYvJ9xS0kKWXY8Zp12mXZHi34h6IhLpn55FZDz+ffrzFfsAlzpHjR+5zVY
YtEVIqVsVqxBluwiW8VpMEkNGlS0ZADd/vx5KgSS+BMdb33mhXW7V78JpJrjthDL
ev120INpmxnzJThUytcZ+4+DmcFQwFIG/KZaCtIZp1pOhmeM1i4J4rSmlYKFclYR
dYW4JT3eBQM2quPB8OwkDhlv738lv2dLhBvUb2fZY8DRpuQO7mYYCHzXyR3q0Xq1
4qnW0Wzu2uU5zP8KGNVR0esMzjE9Pf3fgk6cBysFpgh8zDEVGjHPjEe6TzH28R7Q
OfdQMt6HkbgNytNgWBupSU/wdARfaNbvePK/ieKVngMojW6UpITxtfiLdg6q4D5x
KD4QnNTLtUVobUagt/wPtoX78W0ycIp/t0H8nV5yF7wxpec9S8vpnUHOslaZDLoH
mbREDV5WraIOC3fjwXOYT9JfBEwRNy/bv1NipZt9KeUCJNmnycGZR3TLwIXJ2AYw
B8tPZk3APoQFtbKKAuMNDa/m7zDIL9K96YPibazKgROveuk0f+0U7UEj+jtTfyMr
IFwjGEQGOZHjgmo1JhsmLRp9U6fP1Jg2k1XGunh68HkGHcJxetIrXDuvL+ns7Cnp
YSllux29S2Rz9gmTIEepoB10cDTyAGVpTOjEb+igmVWb9qSe88uC65xG8Z5KcmLh
tL2rHjDGuBwz0lH4tIiVKjlNTieNampZMc6Fp6bFpjAZHvptL1OOlmX0ShGF9gBR
62JSG968HH3I8w46U18Do5LVRdzlGYrBv4nS1h8t0uLt41VOlZJxVljmZ7KPjVY2
xCmn7yJ4GzUTVtDnvqTiZApQSJ45/QBZ+GCsEbYnerloR7vseq5qiJBc/5qnisxu
OnQYZZw9a5DRFDqJwDl1Kd5un54bMD+XYqnR5SYz1bxLFiQiHUnSI2Ps3kDJItzB
jKWnThZe+YeP3KcK4H8zQSWdyVzmTkUzsePLP/nkwj2z+8ihAMkpLZi9bq4FcjlW
R6WSrFG3QR/g8CyyG5VPyBgrtvFUdqel160jZgySUpJAme+/2Vvh64E6iHLpAR2t
4NNhle+SQ8GCjgto9H7PNwx+/gk1rDrx/74DWEnMVTm11gYlWQJs2+pOSIVJcocX
t3vbJeU61TPjBnWvuv0sHcIBm0D32W54tx8uC+bm5LvKJxwLvHpnaYCIKFVnk3lF
WEL7JOrgo/Kk+X36pCKbEa1NyrW/vJgDd26jOqcW2nKnKnNX1PYUvxuZzTSDZ8Do
AHvdS84p7R2PVl8QG5tw5s6HQzz04iPreEUrDr0WZLh8IxNc213g2wCAKGrmNAUY
JfcsQFKbQn7qim8DN/OWiC4uqgCWGIcUEdii3VmCaTRPEaGtO082QKsGEaRX+8qC
r2SUYXBxgEvAPJnkzD5ab4h9kmi3jFwI0DmuU56seB+6gxv7jLxg4xWLBaFfrJAb
fgxS0N3jox34f2tQqC7xCItjKaC9dZyxsCZo0S6ArJFKyQkm0sv/tlnCUrA8eLKK
keIEl4GF5C36c3czktyRT2SceV6rvKwTOxkeqxVwfWW3pnxLfAl5cUJXAl8NvHhV
pQPm6olU5ZFBKifdXwGJzHMp8uNFzsHnU8HvBcKuBrGa+8giz6t7kkwPpWVKffmj
iB5NVwXekYGGlwo9xe+njsUVuNvdLeEtHrlJjCcAIyK8Koh94RjKOnezmwPEmW05
tR7TX5xATQREp6O2PORJXUcaszBJd6x6feh0cGcQcCtTJ2QLi1e1MBFygJAjVr24
yJBNvnyxw8bNmxB3YMHnTP27CXuKpo6hk16RZQT8/ZnOVBmBsABkR3arNPvhz4+Y
Z9v0Vx3YQuI+heQ0W1Y9Z62DQBWC/2IdoNq+nDFzfPrBAMOMN5lWQjoh0qLitrq4
yA9GLzUiHfm4kTqK5NpI6eyIMQlZ03Al96iCEQCIuAHk/Y3KCQh4J+icV4aHy3jc
xwAU2PLWGCce/T/TW9YGIw1DpKdyMl/FjWSusQZ//2VPJu7/jiVuwesdy9/sRoiH
EcdwW1nGtExG0L7j/KQWEnoSn1aoJvTpTH0rqXLjiLhLzyIRqFJqYwgXaF1AdRcy
SR1vBBCliQ94kg+Q5z/0OHFqztOXdsHvm9vL579fl/jc1klGLZdpYUIR7V2KpSxw
TXLNRd6tGFYcTSx3NBz7zSxLkXEFJv2JSeHFSouxrsMY/0cEmAoyoPbTA1OISGAi
mJ5C81KBA9DbhemvM+zw6c5Q/5jkyGBBS8ck3znF0WireNI9xpm1mlM1egApYIU8
RS3V5SEkeGb4b1TFNnh4vRfrspiQSb/C/5Y9+Eu9yf7A8N9pT1I2dV61aIUlUeS4
MBsI2CpkUHTSxelXWsbTy5Mfx2L+5xemzIIUpTCfbAU/jNkM7ARW7Pt/LmTRAZWZ
MFknsf9g7LRlcA/cYth1Isk3LTD/pEOspE+D4aG3YAFGv5I74JcCScTJc40ujKvn
zhRmvh43CwuNQ8EFPYjclAJKXAA7dGkTZ5HDFrtY1bDH+JsfFR/dascEY/QwSoRT
cBN+HT0FB3L0QfYPUXi42PC7btk1AQaTcyr94I+O+BGnJfW+UA+Jt7L2y6RGKRab
AXpqwsYkXLbliDB1TR8JoyfVgvHgbWXBMjLzt9+3/k6vOWl6TCE3V7/7DLiecWBz
QX36brV8j1WCJr86+3jukMv2cmC43sN5BFe+LLu0OYH6j/I8i1KTDXzx8qIGTcds
x/gyYT/hZQg/hkuBGYKqFe8XG0FwUw1iiiEBMQlR0e88E6G7u5whd0iq3nhfh5cb
WahM6SIuUl2di4QR2Ws55kIY3wsB6+kEHHHYD3+2oE/yfYnmxNXCni1schBlyMMY
OLswpFY33jCJBorCyKuqbQM3pBy4ZeEVdc0eC23kP3fJ0TTtE8UDmCHI9qxigvMt
nR0U58lQ3Vh4E/Ex5H4wgZf3fPujY8PAOJOzRJQS8GissLz4K98/eAASVpwxfkP3
wdyS9DySIzmQTJ3PNLW2dJ739WM0ZV5N57jQaY7bVdLSbtxQNTisiuGuuq3P9doi
QSR97WRnExmL0VgW8gb7CsmoAiEg/MNyWFiIRyvPTMDULsjOZUBWE/jjYAztgkoz
qR7Xosh1hM6ORk6TDXIPn2Fxaydohw2aJqiT6A7RzIxynALHtavUMuEsWSO6gWQ9
rPz2uu7xAA/jCaS9sofLMEMKm7v3BE+vgon+5s6jbh24MotM0MLYgQlJbolL3r8t
LzrIyjZsDjtOEkdkIzkJI6dHcM74/8eJEYeqdMyKseyndu7StOTRvjTzCVlAYxiT
vJUaam7Je5uJgiWrwMIIPmcwBet/Ff4s6mdqvjT1BP8Pq6qmEPcbACzINxZ9uXkN
2O9mjjraJOcL+akxHPJlF88WRI8Erwt22XDaAlFJvsFtHPmhOD9H9tk3yUqV340V
UhxKpHEOsyJrHEyD4AcltRKTQ8yof7eWrVS41aw+bhEDyAjNTUxS4mhTk1OTuq3W
7+QwUK3l99zOP7plBRJvRU7RKVb8zxdc0oTtS4FqM2Nvn6ZkORUNrk82xQjJrtWj
1USx4kLUUQvVFIFnLYbRWULHfkcyqaDeA284Te/4wCx2GsH5X/QBCT7c5CUZoP4Y
+M83JLFr2kVcN7PX/L6acrAJbJ53c3zEV1dHUOqyUQ5X5LcZVlxWWptOvJ6GA3AR
HUh9hIV1yolzRSksaYzJPauKTWFtYSQ4p7fKMAJni4bRdXVq83BgWE8saa0jA+7/
3ObgEgNmb/9HLQn/892az3r8Opu0p6S8RCTvYSygiEAHcyediW+FhOS8d7L7XSnG
DCwiX7C3s/vI3kvxe4Bkp0PAh8GjthiSwfYQfA3e9xR/eN2TczNp1f9Yrs1gqrsR
1gLv9kWMAkr+fvFHwDpdTFHxEPx0TgrvytScC+YU+FFuWr4QmdAt6Fo1HPMtJC1E
M8RH3zr2/y8OrAro+YJTBfrJWJa2NJWEF+2HZfdVpgAvR5KtzsOKGz2K1poI1b7x
91Wzx0VXmnrBpbyOpo2KjGYSRUIzZdPVPJjN2UEtm1+ZcYo7TjBOpVKiKVd9aG/O
6eN+p/CKdjdyJZiRKUeOiUB8oAyGm3Z0m1/hupvcd23l8o1GjF9ps+RKWdsHyJIM
Db12QKgkgJijYfimC9/Amc7HvnFcwCmkaoWCTncQuoTmWQDIx/V1tVnJ1cuDtkIM
40JsViGtEdourzQ1y0XH0/zFCXvz/iehRYeLVQbXJrhLiJEENn3oki3pkuxQvSpN
yXHj/3wSuPJbbO0YAiUPei+2Ge8YGADshtxMsyN1QIKFlIK4T7sDYmnrBRteXHiU
ougtkwCzpKyeKJG+B1ThiJQs8mv12XelvtvLksII7zgs7ig4kSI7dALhDN0ykL1H
yR0Z6PYhpTEbPNGeNKPtbwmh9pw+bBZU+Re8VMfc5gV4kv9tgKdUaX9eN636Sqgy
551irpTo8BOkkL8Og2caBcMDugxNO3J40OCBreg75mjpkVVFBaY3zfL4Ano1iZbU
XDtxDEYz9G76D1q3FrR1qgVFgjgmvpxAcnipWbACKBSoA9UDk7sh826WFJENpTVU
tmy0a49b/zLjJXsp9Y3nMnYA1EdgEtTAVSTvspjboWMFNeJ76aFg8x4c9sADg7nX
FNPgimeq/cg8PqGiS+xt9mCCQBTB9wZ6ebDRAXYyegMXIucWKmQqUXeRHoapaHFh
cQJzqzwqXssc5YYZfYR65NbKV59LJg3P8CeelA5owd3GtZYtwFvcf5qPROx42sda
RHaiBJQG6Ba8JazYVOTD1UV4i8Wps6z4hbVvFFT5xdeEMDyvcvLKprwbdDzvyQZS
vnnKJyo7A6kSGOPPDWg70huKM3BSCl1LPTZlBqoKLZgRYRD2UbQBfY8UEaF4ub9H

`pragma protect end_protected
