// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
EpwgX35RyWkUeUo300wY5tcrDqEkfMZYt6bcTMDStlIHU4MTvWB/lTGkNQ/kBVtZ
LOMrJVHKgkdkGpHLnM8L7DtkMSFavZgJM2OOvrF6jNMBjKkrEwMKgrSIt95De0/s
M+9gyO8076ISMHsE2zW9VIAvTe2ef4Ygk6RqnazPK+s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10656 )
`pragma protect data_block
sgSXo0L7I0bxv4tjKgDFDJng0DgRBFXpZCXRt3nSxz6jiY9TGhOYH0mJL1UCUepg
5x4DEuSYIR63FbVquwj4mzIP/4DxRfP5PeRZgj7UxGWSlIJWfD2CZp67b1AYOZ+g
+cjT/B9XuHB0qOys/014MHWCGoLK388Xe8b7iXyjRqR0Be8+xzdsw/pZKeIHJrhg
olnOoe2DpI5cTotBLHDxjbgzZt4SycDFqQIV1jO9rzaxrBESMB1o/zKlGe5YmWOo
MnzfQ39z2UTkeHR7YRwkf5IcfYXBIksP2msAn/gH1b0afk2Ga4YM2byC6wYS1cTt
LUow2HffJKFthvSePShS4NISe+nMmoDNFKuCt1lGNHSIMRa2flTjhhDoiCYEhOV9
zoalJZ68GG/NGNhlMCIkbGt4MlL3RE8OlYxK3jgbnvfj+PhEfm+pLplADoEA45fr
UwhUfK/a8azc9S/wfBWJ1Qc1VVVYbfoV3jFGiL3njupMPge0zSnIa5sq1IIV/ngw
ggw7P9KkvroVd/vYXeUN1+jku4ZNXpPGt1It81grcD59DjrJygkO/eAea318O1te
toTo1pwa/BVHRtW+uVGQaojLkZJgPu3VRHgB2cz5ajM01DI5vrbvkyB5Y6KEDSvk
b6X6qqKRVVBWW4zIfa7vXyXCi6yWT1kF0kt77uHqDzxOfdJc9Rw3eZQvHoxC0Vxl
Bj2Ny12yUqAnJnFLXTqD1Q3ngHvwtmtPuLwuMKZGP9qza92HVI0YXndq8RmqvPIx
DzLC5Wq3f2d04M+5HUmtyH5ZkwcDr4t58Rqzuwjw8fuuYBHoBRAGuS+VgzQgbAJe
RGAYal6E7Ila9tAjQVWWCf6Avf69mPF3f+anD7X/n/VB7rIPLDj00cQ/raM2WKLV
bLBx4n4HWGidhj+LmjoS2eBkuqfcq1ec+/qdLfD1nysndRAPiS7HUtYdsp5zBDvI
HKovVVXLPrWeKaq5nBQeLAvlxo96YBPbEedicn8AhY1C4SOlQ/e7QkXDyXt0ZkI1
k8E3pf+Nr/pG6HBKCDCnH+wM+RDuOQTt9TYv9wM3V4rH5htnbxtfacP/tUNGT+Cr
0Iq8YD9pOxrvL2QaMirE+IW7PcUjqLQYjymwWya+IeYUUd0Z1Y5ujy1qdMVVDpjY
JcoS3Zxk7UEnGKwrryR66DxJOD2szj02a8EvTz+mVvfJZI8R7SLSaKu5/fe6H/t/
8WPQ3VsN8aAr0m7buAe/gA7LbhPD/37A7fUdg+stVYZEm2OPVpkQ8bed1AA+aVgC
8ebgGULiYPNJYJ64h+aYX9TpXOQwa5cmZujEMCY11SedmWdUV+TUkRUNXYphJA06
aNxbRk7g/MzAiR+BUY/5+bvimAEZV+8/7buMIf6zPjSrEpr9OGfekfjxfbPv/uOj
u0p7bpbSvQlMxXrBAOWyMXbAnFVI8vKbtOY3I3OIrEQURyROlUNzIxmPL675/rbz
FqjN+9K+aTSkm1x6fN7+YDG/BeMPoPCSSlchg4iMhUbNqfUjtNWUp+xLSyWBNnQC
YrE3NzaakUQNOAGWeW+8h7eKi3LeL9KBUvrzkQPAC+rMZ38+NCOJ+QFqlXIyOYMr
AH1qZh0rgf2me0wlTwGw2eEBJyNP/zCxflUZgyt/7/HTisWtkWlXa/bV0KF79AB4
JsFW3AfNlj4FF8MINb+mEDT3+8L9uIRs3j2rYF8L5yT3wyCK2ptMxi2llp6cHANY
D11fsQTj76h8bGvju6ypBvMiEiGOWXa4Iajvlyn427ArcMLGDPojbpKzIIi8l16Z
NH5GSt71rOGTfqlbWzxvzk7J8QFKh3xDuNY6tMFUUDficNPSRz3eZwa2oR4R/SEI
nNObo0UqsBPRfLsp+2+H5DBgTS9VOH/r0uZSmedc4xQJ4IoflyzQjK6yBNpuVw13
o/HLkoN3a7JCtJ7qur1+R0ueGXjol1B2eAr2dsdxJYq6VyiOSnnHyZTox2lbQTLY
YBSml8i1TJP8ONtqcUGMmKUAQP7I6Nt4VG52g1sMPLY1zKy4gH2boyTzBzYpMldW
ztISNE46knMVa5Te1/UML+9lTlByqra7vyMjY2q7Oq1lhWOt7m6EPo0cBih0Rruf
sFGCT1/UvPZGfhVoWVlxZYy4kSjsjHjSrFn0jMe+O/QBtIgI75Bbx2mB+wqePAb2
ejOq9XD+u+p7nCZS3wqs2XX8lWI7Dv4Oh6h7lr/63o0KVpJQjx9+I1+9R6NSxW12
mmDpiBHRhWawad3ayqitiOJ64qa4QkCWbUvBgii262dNBZKsq/h14tIMQgU8ivbt
pzol/Hqfgpazs8St1TJLk1ZpI1JWczQYZanBfGdUO8+b3pxVKpt0PbXbNdyyIOZD
9V8bKRnw4AzCLGl5DAhZB68tWZOHAGvEgIZCHqMHk+N6rvrLxoK5pm9UzOQ7Czg7
wn1qseuKdZD92VyPKf60EI5Y4hlECm51aHUvAvrl2D/P+pQkRv+K6N70uIuxuAnh
m3qMIVw09Y8U1dz5cWxZRGOJxRyiFYEMuOereA1lLxKstwfDTf5jWvVZoTzuNKPt
PKt6d/JgYyvDsI2LoFx9vjVvoVRsy315+g8LL4kPDPAm9CaCAkIa5pKXZOGlK2oB
bjzhzeud1xsVZM+xArzFsRYKn539fmcuZuhtvekRXBc/qaA5x2wV8t+VsrE7dq4z
t5Aw2iwFIyoTvqaqv4NNsmcEEaypG0TUH4TI6SCvB6YGagH+LhByAuxKRHaidauo
X4RK4Dhi4RWlZxaHuHhhnFOubdPp8sxtCqMYMhrwk86fOIOgqofCUghUANIvhY+V
2EW3Hf/MJEd7oQNLJPcwT3OTnkiWtBTBpdnLw6pUMbMIZHPV3ZHH8Zc62BjAI+a1
fcYVwVQCWH0cNcMaz+4wRWrgqyeTRymwk+MLBMjgEYOrnLgu4V+osbCsXq/P5P8w
37uXAPD/KGNG+bJUyXHWxiwJkF8WD6lXphKTubpBXqdtVkILoKK7t4K9BjcxsDDZ
zn/kKXHeIyauaFRRFglu23WbksU24a11aAN0C0SB91R8wNyjKD/YChuACvReomWM
RvXZEPnh9sPpHD2fxSMcpIWuJ/QfaOCT45ZJ3TlxF3SWtmyDfjM+k8o5SDAZHdf9
7GGM+SOJLsDmji+c01ChiX9ZyJPrss0F7k5UAVZS44kjBHf/8GkXNUEjFIIp6axC
HFydFIrrS7t8VggXkLvWdn9r7Jb3dJG2MJ6ocmaZhFyhUdU6SMM7/5/MKHp78flN
wFuDNSu9znVYc9Y0nYIQTZDMD+Den8qLYDK84wP2lGlkzNrO9jFn/0jVsWtkyFKi
4iUDMS5951f8yQ+ZCrZSy0DV3MKH8/nMoCgpjA/9ia9g4PpPd7xsKBB5+mqsXMya
7yBLGJDYOWCMx110NWHvFxG5MvfUFbTqkXPfBuyW0qIAp8lafWvyj7S2cYtD7a7k
zhDDKG4DhcTzmBde0lay2x4iziVtzC/6BcT2pGFGSPt2w3jMEsY/CHT2ExXIkDjd
YD63bYOc1bmCrbjffY7C3S/xXz+DmsonguNlrUaLv5Mw5KsFmq1AvZRIfHO1TC/r
KthmErO7TWcD7oeRtz/g80L3Kyb8vLuU6x7m39MehYgzIeTN0lZpUOkftihhnHRn
UKEoHRpIm1Ghe7tJFhIplUmRM+Mz+nM+AF0VPQ/7O/lRFCg612wNhr/Bwfps8UX5
+A9zdn9sM5QT9w0GX8YWPqfhl3wxzsZnS2JSdVEMRnbwVrv0fxDZeCWghbiWl7LV
itLulh3NbE94TH/x1QO8Uj/0+ZaKhLQXgDPsxcm/u/ore3O9XRwqUpmgVzGAm2bK
Z8M+u6fwBnm60Itlm3UV+x2NynrrWkXs2wHiWFQvqyUTLsviZVSAOXBkjPgwNgpx
uJRW7hX0chxI2cgMSPCr+EvybYGJvKVAMYXcHvCJszqoiMTabJ31VFnm4jKe2Wtn
EVwAp1aK+jH5w4sJEW/H2vSwWOy9pXvLwPTwv+RRuX4oAAKN4p/kgm6ve7HYZ7OM
ulUTOWPZSzj7FpeZ6I+MGwf3x4yvgiLfcIr3/tZI7xl2vxHaVL4RVu413Hy3GjWE
oA2m2GBSN+cTziWTutBij/Wh1jjOR6I4z3frE4tCIjDGMKplIugcZZplgBl2YhT7
jO+3Ar+fMOlVhByEbfQMA97TcBpg7ZM5ESzN7kkGHQ53GfKWmAcAtMYrUrUuzz92
NTSAVBB8l7T1n7UyQBWowU5a++PMe0gnMTU7I3ggRfGVY6NxDat2uNoQ28BREML1
qwkSDaOAMIVgdIqENr9RL4kNyQKmbCABC3U9msUGUjg3CIiSQYXZY8TDldLFfros
Ddb7PkumAhR24ron7TTuc8OMzJZBCMQBhyg0NwJehtTpf5grI7YDAiMWGV9NQLTC
q0RpvJtX+XXhH+sDnrTn0WL0+SASACQzJM8tdeDfRx4Dl8iSX9diLlJSXLl9Jsfu
1E7ZK4D2PFddG5xjCL+zpesWI0NyrspbETKVkYQ7XL/c3wbLmZoPsLh3LLX+v1dJ
ypiqbjiJAYWUGe8O5v83vt+c0zwUOKoB6GTTTm2yB/MW1IQalV29fagmO3CoFjPe
fvsFnlfJ7ul0MbQsuNehhJuK9bG15+62L73l7oxFZFMhWovb1LxmM4I+QO9wF3vS
ZNdyWEGSsQNa5aR+3YsYCESRwYN51Of1KD2xYlpIhc18Fxj/DSuWFvrGHg0fD7G2
t4tbeHnK3IQ0tSZG0MKrYViyGN+Yaad/wP07l4J64JRExic8oMBqaesuKh07pLen
B/fAfuuLKzn82tfgddHwPYbSnVMF1o+l0vM0kGo/phcyAyaoJ07SBeMjWLW4bhG5
vX48aYeDXTF+cxHIGCqBc412hdz1u2NPAhYYqwZlnDf8wQemnAyGTwUrkhMPY9dD
1wjQZT7xJ8JUBNcQAUUObM8Mdf69ucDvL0gYzvvok6tEE6mwKwFZbQDe4IdfUdY+
e8lOChmnHakv3sc4VmfLgJeCY2da2gvqi5mfVjiJX512yrmDPEsLwBn1VMzXx4Bn
5zVeuoKkOoMxHtksVMhCg7v1TL0Ka5BTR1ja8U2o8Iu1PjwG8sWYufVorXMbz3ol
QP/UQjObYzhUZ0FIOZ4X+nLGn1bxy3lNeI+JbUAK01LWUgIVoFH0Fo+sZ1CIdNhO
VdPguD4q7XNEaVyndD+laf00P48D4qX3qTOkKuVnBkP2FCBYSWCdC32Y+uiWbUGg
OIUTFyhxP1XH0dIYoklN/l5qK7nqea4XSAFlho5OBAugRVvfuhV23r2xFQZxmYBg
iZm+QgNjuhdlcnZMx4iSMNcZIh98uPRjQPk/5mi1rX2tD/2rZ4hbfFaTtT7IN/5q
mqvG5HAqVkEg/xG4NxaRJTEUet92YIg2HGACqsLko1vZ3PboP+CLVaf6btvhs5av
SdAAQOZHZRSrH8iTgGJY4oUNj1axlEf5SlLeJqUikcvPE16PzUXrsNLfy/djARF+
iTu3delj5LbH7PAjrOYzgciPj9475GVmqzfL5WIa0J9jjAH7TTL3PCxFf/dPVEzx
nzYYIH3oimF4NZAgxHcbDm6+R60JRiXKpHTtlOh/iU/oglBNQpZ/6M8KcxPLMr3q
IDxTMcRAtAtDyJ6z5364x0Ji/bQkBO1j+DmKioERr+kmyhlK1aV1S8MVkUN+uLzU
YdHyLqT8fuEsHF5VkF4hlllUhuy8wWulJhRU1hb3WyWhqvIF2cmJwLsKj4FG+24t
AnBVWTEGAZqIwL24KiYHNZvpLKtOh6SMjFlevCHzuswLkElYnzVvwt48eaWWhywi
hWSQ0u9XXKTyBfd3v1dFYVCYr4+zeROcdvJhHuNVyWc6KpsapzuyFFv+phERigVW
TzQfdXDT6xYGx789X5yMQK7TnEcdESGTlHCxw34yUMzPpV2vKO8KBew0QbmwlvSK
UHWsIEdMHzVdDey+k2RhsS8/dmGtP8NCEoPNsKoq+6yrrMOkVpBnoJgrNnBvcRq6
4/NMbF73V77zOGXKhXkgz6xRqD8Dn8D9kkZJMDpXQzzVn71PqEa9cll6Iy7wqLB/
EDge+IcolM7pnbtetLU4woUD5Xp1+ztRTfz4fZtfYGjWPyGis2jF1893ghveQ6dz
PI1fZBSu/Ss328ml9ALVFUpgVzx9KP2SxLwmEZybf1Z6DpG/HeyasHHl3XcwkBVY
/33qJd9hvJ2RT3XbATBm3hl+MvCvqDUJun6weo5Spi+dpZKDkz+wVu0mN/coT2q0
dg4o3nwSnRMfO3dG9/VPd0RtrpUyS9oNjFSk+BqySwvIdvrNiBp7AUX8BJ96PTH9
s4nwooFnVD3mNy7Hz97Vq+BW4ovM5ax44FqkbzfsMdDT2uWlCZBIBvXEUdRmXMbW
z9QdPvjd0Eg9tjhXmqbaaXJ9WPJbH+ntpXkk6XQr0lyYOdgh1PDq4KUCaavsT6mv
BZtvKYQIdFniHxiwVyGw3TIHAB5XDPSkLrrsr+ZemZl17kSECsvrtsR6hUep5TiW
BgnBvOkoHh+O1EurVcisxmth+snr5diYA534XuYZzi8yjsf8ykhxiDNMNEzW28gH
r53ueqed4se2Vo3NqhsVko0CJtgI1hQ50PzJhSx/ocMqzOOHChb7IDcDUdB2Tz5w
5UBiRRufMXDss5TccsMmnb1hntrFuDuDfTS4wltZTD1EnJxbt66VMFDBtObFHSVi
HaY+CSDnyekg31y/nCZTdPJV8iawegOyxASWi+wfFQzCh3boGe0KWvYI9A3DjbTY
9NIkBKYTT+2i0Ln+GWeD6ZqQocZs4G/uxM9ZlTx+LmU4B+ElZAJIEcEScDRdtnbg
0OZuDezp7KORFqrTqx/z0+VUrU7XfgcA4DD1HMxiUP8pfDn4+2UQ88QB15tztJbW
RS3mADcKPM6iOD/6iAQ/Vw2s8ZyuXWW9ZQbZQpeLBzsdllJn6yv9aSITfuIk/Zaz
rSUPvQyzbdEcz0fBZ3qUdPFxmeo6fdh9ACOEhZDQ8pCA6VzuNUQPbliy/2OQy1Bt
C8+G8xGMkqkm+eCyOc3RI8kNcvFp8LUUWMuycY3G0oLaQGdO8kpvf+UcPclGDTI9
w8Hu83vTEV+BV0FULZxUG0aWqbNkCkf9hMmtx5MPdGLOda6YsopnVUQe4/fe0gTM
PZlgU2+pX5ThG9Y8D344fSvF+FzuaRpfhPXT3mqvksyop6POrk/3ynRa3Ka4B/v+
UBRAHAj+yGKPuDpTcHU9gH9I6U6bZ74iEKjVQ/fqNcbLLi5OqGlzVGhf2ReCbwCY
M19lnDTsRl7pLKykPO+fGM5nz25sdqQ6A5du9UZZQEv7UlOkH3ZT2kVvSoHg/RSu
/Dp+TiJg5CR7WmpzI9X50QEkXfG+aAF7H0TYajt1ZsI9iDqWiHOjJ1XMb3zB74Pd
kwjOn7UsikvHwqzZ9YIDrTG+uihUi6MR9pmfS7JJpyX6OdeXKS/fMLrWB8eCrPEg
/Szy2Nv9XFl0bAsikJiW1Xqrkbp4h949ySOmuawV3Kd5ll9K62H0pG20Z8UbfKw5
y5vniPE+9MvpHWfMPuiJh9zfSO3DjcxsvRe3CeKPJ1ZBHomESayAnz0AUR7HaWEv
drUfGZ92Q4oFQAYI+b1UJTZIjIu2UT4zEa4bZhRLP6NrXB0PTaH2c2+vFEmejaaU
ZWFnbaX8gRnzUKpx1SNbFFnV5fsijUCei/eyv/tG+fqlD5Gc2Q7sr2Yhta5uoohM
hO2Xih6H+43u0XmzAHczMWyiTiX3ccf2+5E3TYFExE/dbnvqrYuoaEMEnipv/1MF
7JeioKuxELHpgK8GMI3FTLC5Tqnss3ofGYZ84dUw/iYgnExxCArT6WvBpYOJhwIV
fgYfLesztXa/3ROoZUQc9jQD4SiG8b6pvVK+mDE+iSf8OHVSGurMwSNyuVLT/Y6J
4jpX/SMXwMrfavRwXDvlVSTqK2JepFnhaqDjMkgS0SRt/We2MCg1htWv/9lI4N72
boT6txW25SlzFEJoOuFr2sX0q1A19UXSfuBms5OT1kmhbuys7SvnpdYVxCmizUo/
IkB2PsWi3APDhRXE3xCEipBjtuuz+Fa9RbkVFHZxeS/5LQKv1ZMA682/grgltPCr
fjnMrAzTPKv8yZzyrPpVQrqxUPunuI+s0Ys2uOVDou0tW7KJVXXYS5vC0C8bUf1x
LqCV1bGXkTklLdIlkTA8GP2VE6HWnw+AXZrLmpv8s8+vCRxSNKpPTkWnYPsA1ue1
qrO8mbszyhOwJ1KxaO11uFz6ylm7Ut79ZI2CaVUPJhxsa2PCIjTTwpl8lAK191b/
qaD2Ze5TNlpoTyuA4Iu2ztmdh0I/u7CC+jqu+Gmtms0d2WaXhp4+sjQ/rOoo1wjx
Rumsg4f8B1PhWTu/toK/+6a1IX7yOkbxzTIjK2YAsqcWuSfzifOANqUIIXZmMcn4
xJYMgwPO3bOWCKX2URKws/5htFJZD37v2MiVLfbk+M9t3ESUxQtpUiRShKLlATiA
Ho7imAo0GvTlJ7IYW/vuuSXJMItclc1mDOWzUPjg560XUX1J+BPR1deMrhUCfDe7
7NT3IQVp+lUEMQWhdZyu7Kf7nWYHziF7aymJELRRl/4Ubk5+i1mZO4HR3y7kSGZd
ImxfKZUVdQWWMRcHzDOvrAXWmHcJZB2l9Bm8eF3r+bTrrVAzn4x1GeE1H6juC9Ax
6UUdEPPae0R6swDbzYhAbUAUhnXhWA+qVGkC1g6KUH4NQzN04E1m/14Iq3dUrvV8
mSz2sOYIoZNCHCwKq36iol48L7RCr6HtQiTCHg0OzFLFlH3BEABDQxfyUFoW3MKD
2mhL0J5tfBF1D8D7FcVymjnwQRmlfgWcdC5DRNM2p82TbIDJzdAXQ+kGIdtOizqO
+lm9SuMaj3ZQOKy09U5j67TUxo0fPXsL7APgrDpKb/pju/jI2amOjUHJTDxiqY4e
7EG3ekuP5Wo9sICoMO0e9lgohIeOodCAyQuK4o8X5N2F9rKsuYosSSRWUlZJqA2A
IlQKCBAG1wCAddorhH7gYJ8HzzL494xNIrriYLftY5owww8b1YFMcPdZ2XRX/dbK
J9PdeSCqka8YCc2UG80Cwl0QZwGbbyKNU+KekYjpYQJVRjhjSRkN2JJDnqr70X6+
ivinO/hwQnMPJ5qb5RwdXH09nSgJm/wogag6Y3OFdJQdvzb9dVMGC7tbVVGoDguo
T5nwoarjQRsVHzgAyUda5pegF/PjauZjlokcnDveDmdYtwxadyLH+hGimASFw0cr
svU58h9Jf1OvlpixNANzyuJLrGxiztVL7yGYZ/n5DrH8eDMFupahC8sw3KQcu4Fe
p7IPrpZvppQG0li/fkNNQyFQ0cu3iqw5AJdhtxUueuY9N3Or+dhtuqU/LUaoajks
0LfEnNfbdLD5I0vP8pZFU1e3dwb+/4JVSIELzHt6z0IInQMT1UZ6yzX7AOkPYdJO
p2SOOzTs3NPx/FXeEV/Qo3C549BHVmmKeVK3Ot/x4eSyWO0WpJzx8jnQHM+6apE7
43uM1r6RgLYLsGWnSbq3nIIKmVBF4hZe4evcoYPaT6pukKLEr07Qt6VRra23Q6yD
yJbool7Ftw3+gQ0T3IofYYM3hDy7SeVhyF8T3OJBblIqw0s2Qtyzlw9qRkjuctio
1C+DeSK8YnmcmLQJOh4hPmJiRsjQ1mtWcS4MjS2VesroBcV5HhephKAkBECgTxdO
RjUAoOKxTzPCcB1jdWkjaIeHJvCSi/FPwP3EMl9ke8DGF8Zga8GLhe7m9xM14pUa
ImpQ8ilxBQqKZ012AnIR7OekVonsELiHdO/yfY7R+vJpTTwYEUe8EAx1/1nU0tSY
FEW0XwGZ1uxF9AHCp6nEdwA3h8AEYQMCxAS07nz/KANo2TrrowjHB1DlgV6pwa4f
7JxnqSY2ZsQx2Gb8B4+E8L1jDbfiaAeMcpXM2qbJvt0AeHf/BhTKEiwffl0fDD5t
pRBl2Y9zoydLP22xSM+3Oa/B0LqULKZj72MUkCBRVq//BAtggK7rBkucfONGqAbZ
Xgq+bbQrX96N/Nes0pOtKG5HNR2ISvyu0IB73bgHQVWCdFoGCa0r5XDVW8NJxUe2
W9gZkn3tLsyw1E3thSmf7yO5JBMZL5IKRveMb94bYIlA503H7mu012yhghKHYwNC
N39CupzXoDmtQV6p/HYntxLdSWNP8BKCd3CjOcG82gK9TD4YdMSVUsO/R8FzC0cA
GXAOLq8+r5AwxGSoHOTnXJMV24DcjB9YHvGiaLgDwtvcxx13YIMrbgRnEH7Ti7im
/ZLpa7v2ZNlDfDLfp1i1CEGb/+8S1HN+4TsfqfygOgzzcEpELtl0ChKMbbHKXr6y
beLd4JgUszbMfq1Cc9XhERDyQybrV/Inl0FglwDGET/2nHVSFRdwmY8Yw2jbdQTO
ujYtEAiOUZ4e5twZisStYHEDsn04idfxcnzXSsJyyd2sGI9nd5R12lc+o7mFfNVJ
D0PWnsEUEUDGlInbSyQ1Ox3BnkmUQyhnIuPJ7s1U528zSxikjqItDpLMkmelyobA
UW/kb+jNu4zrDdil6ljidC5G4EdHaY53R/Vm+X03ZpxpHTzSKGYgpWygSgBG33NS
tqyXU0qVJbUNXNHdk6LtZSEWz1vOP1Lp8UpD/jA8xh1IYV0CIHEMqT/Wq59yakAS
lQoncEa3Os9NIRK/gQ72fXPTmxxqZOX1Eub0Z5X2AVXB/xPcGvv6Xfn7p/aKOnll
/ISsCQKozvs8FPjQZDekIJSp23sGlKhjuChEQ8VFe7oAO4y6pIr4m9T6b7Flp5jS
8lGVGF7zekhUv/Tr0l2uBBIm5Gxtntnzdntl/JepwwdZBV2X1+4FkijtCrD8bb23
b8nZF3kbNr7ypmkfb3vyV2P205OMTu02ETQiw9vVGHhUTeLY3CUcGoyshdo6WTD5
WbTiOUetzBLrgnGm0Ey578KP9r4bBaoDV3y0x6NYn25GwRUI9cRep2rl4uvy3huA
U1QJcnaKP6NI/uXKsMgwzmWXLEh4XzkZgWQS8n8Qjeo75XC8RnjCyEPgpL8P5MSV
2Wvrw8UXrIlMNZENBJ91nbmr9aXppMOQgvj5K/S7wWUtTrYE7ZfDJScoJ+EESLhb
/cnXoNPW3eh4Gj42ak1CW6BtVHjGliVhEflTZSzjGF7oOpfaWDb4WdHxNUwM9Pr8
xflkB9REHJoGmtUsXV5eb08RhUYX+vY4tQU/A1zf4ni3Jq530Uyceos6guh0EcEV
pL6eCTz03zIotOgWdQluqSu45tJ+mvWlDC2N1UpTOAtefm3H0VFvNK8cyvTCJqkJ
eIzhLBnOi+JJqiklR6JGOuyGYFiLJxtx1tNq1Fa9lTPCARz+/0SR/Lj0HXN1mZ/i
gw34E+SoGRAFfBZDqELMGCtpoigpyCD7PbI/yYqYbiU53bFAMDseBjmHgLn9/f4U
OFO8kJ+xhJWM3Co4cFe80UYC0pTqPTUlvIQEXn1zubwqcw2haIenYL2JPPLly6QE
zM4VYXeZGp8d0XEmrqwR1qV1bZJtSjTTfAEA8f+RvmVV6B+Pw14YoD9c/PtYZ4f3
0SkBJs4FgFdYpYW7gIlFE7SdoBXGfHa+FPu5kGJxBBn5yg02Y8bZ7mEoQuWpLYB0
B7XfcA5K0+pnKHh7tJ3SoSwn+HWv/g5ZV11b4vPhuEFpbu3pWWj4CS4TV/WFpHi8
2ieya6GdlbctskA/b4gxqmWgcKzkq1+e1bEWK8uLpMszmZOe14AGuVBWz4gf4ORv
TZ6jpkGPVfjP0EnvjnaHpsV83rquXHqEBPURzRc5CL1FP0AkqBeahSZUF0BeSeX9
cz3ulZlSs1T2pAXbgFFs25y22MjacFwup7PuelhCQzxnthwcpPfauX2L7W8CRJas
+/xoGqvpt0fIsdpZ75bPUU1CWPmweysNGWhDyysrVd/9PRgOfaa7BX1xkAPHs/OU
+JA6IDUmDZrO5uzl/CBQ1r8bJq5/qvAieWyPXrFmuOPVce81KKIE2dlDxd8y+gAc
mXCZ59d5VsRNsP8WAMZ1vRQxyOy6Q4mQI3D+55Lz+Wqh/lgWB7I+45QrdVBC3t2j
YLTZeK0/oltqp6jtagFrcsw1iSAYJkIr92JOEmkkuVrsvN2VNEvWKBp87bCbbrZz
dWF67fcNzWlE+jPwWPNEYG+RxILs4T36VY+EIxGXLFg6cXvIZOscT5VrUu6XBpwZ
f/uVhFb7t89+Ko7q/U15aZBnT5wZQv3ZjeNUNhhNcu14woxsdeD3Wcld2NnEYNcf
k5RzDeAUEfNNutFl4675ibYGbu3yn44Q/ogQ+zH+qAhHqIIbnlvHNurLRPGFw7Ro
sOkYDLlSYvV/aS2RX17Xw+b5CuUAxuvVJdUJ0qXvVWhfW9FKYWEb27hj5pHuojbO
BzGhIYdGIHTejlbO7k2kk5iqDWDl3LHHuun2osXUzDC9e2X21xZvQ9xKW3S3r7jn
FnfHwKilNxkDLqJK0xJBrr9LPtaAz7e+cj4Up8yg5SagZPvOu3E6fXTBZ2lyaZSQ
1qc1qkZoNoky+py57CWhV1vyJZ4PQOZ3GZj3E0d+iN0ErMUD/pnponptVVrQL/Go
vAC7/vobAmT4rZ85esaJKg7LMca6u79CRxZsSRVqLcmRneFlfl/itRZ891S8MOnt
0A5gHOb64ZGwGB66Zb5zyI4w5luLom0UzkW8PA1w2Fnzst4V5dwMlQUJkldQ4JbW
RmEn2QsaBToVHtq2xoIqkHXwh9i2w4/25k5dK5/Q1DW50zoEnJ1wyWDHLNN5a1Vm
eygfpHQy6znLkrqKAIlZxnObW+pOeNfocSSAOtX15mnbSv0WxAhzl7agWMj0aZNn
ZM5wCKSlj5v19y03qXbX5t6kEJfMy12yCda6U/mtprUo0yQ7F6lQl3IbNuHqiZ8a
+uzSUoG/dxVKjUIslkYT1+n3uOKZxndXvjFsFiTXqSUqAb684nokNL+sLG6xXbvU
unIvRFUfr3HugRQlVY6bSEzmpfHVLKWnokn98rVV3vVREMViwk0YO5adkfGLlJgC
gCsPr4WJfUNnd5ox3siKgGgRxffu2EtDzjKSSJOoHByzXuMYv/tdIxlmjoQIHZ0d
G2y4NXEG0JgJL1sz35T4P6b7MBq7s+woOg/VWygjhoZaI96ZKS9h0d+Eh5vNGQvO
gdkrzB5TdYok1cV75RMVfl56426Np6YyPst4kxjwHGBHPiAhaSn/AysHrDnE/o3d
uC66T3HqqJgZPzDLzNmU73+IbUb4UUkI1anOq1BLMAAGstEe6F8XllJgm7VQvbtb
4qUhEuOLk3HqVWFurJLRu/Iz30md3WmhAWA2ayVTp6Byq4MBP2IxPSJfnoR+viJR
BuyieGcIMqPFs15B50jwOPQFhS+u8S6lBkZTfcfAOrkX9JJmOVujYjGUo85bHueb
xgT1K6CgOyNkdhLmMeZ7W4NPFVNhLj8n9U+EKDpjw/D5vFjQSSJaRDfA78HijbrB
p1xurUN4UO3HY4Qr+3k6aLAH3rYewczEYdlfUQiVgopvG2+p5PS0BNjJUbOm3Cqe
/gEwzU4Si2C4hz9Bruj4MSXnCws8AAWlCZJlZhb6Q7BOSJyaScldO4jwXaTtNPd/
3NCDLcDYfYfAExrXduvgysYvbh0BdgP6++QwglO2VeCmfCJ8ScKaSnVWmjYPcWJp
zqhGpwJfRpzMVSBQ6sgc/PaL/IhetQnOrv3V02NIH7fJzNvzPOo8ELQc2ZSUNg+j
j1cVobX5M6bhMN9pulwCp/O7t06oMWVmeMfHBJVoceabmdjxU+NLNKdgvF30Do4c
gzJBTimQ5uSLZ9H+TxRYZnPFEsLZMXpOt0LRAeg8anNKgxFBH5QHN0GloCgXvyjl
JMwa/bw7oAaCnbbikhM7mwkZTaJrQr+qK9/sBfoiD19MwrRQ5ENAK/dc+q2pCRm4
LzFtjCq78760jx1XfJfFsNErYHEG+d0/uIRAHbCQnel4PgAOhuZggRsMGtJsQIKl
o/Yf7YrUp8ixJLA45/jcer9+VH+GG99p8higeX2Okya+S5ExKbTPlgf5BZT3UQZr
htdY13aeizShmBVwS5zRNtbnlmTqV5njyDbFT9oclfJzk2a65lCylJVZ3E5AKKFh
HJQwOn/IPNBdSGKHKhRNb7WwKvtEYbgAKCm/sv0SVLTR9pL1kv6jmzMjYxiCZRWu

`pragma protect end_protected
