// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V86oDhTm8qkd2ZbAv/m7nStgTEKtfoAxnUIvLeH5PPCSkcN+C4RT2GYJriSg
HQ7ksbppfOUguZiWCUQurXylo0iQqDJ4/mdPDLPSS01jfFfdYrmnp+MZPcet
3mY56gQiHYei6Znd58R+KMYF727sugTGowvdaLmzSOnKrMDNwGkKywMyGgLc
8mc1IcRczZPqnuRphLcjAR/qj+H5vnHiYujPNC2aLAftQsETif7K2AxUPUoB
tb9BEyVNdnvUzB6VLGCYbDIX8psdBdPLg9R1cqUbdqavB2HHeFeuh5ju8LYL
l0wS0q1Rrc1UR2A4OIZBXJ8El1JECOfXDUTMqPTJLQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GrN67wQV4pMruFLK9yJogi35F6eFDeX6FsXcd8Sg89hi3lZhVdQuTRSZFtp/
D8WjTHZ/bIfQ7pYnIB1FUEWiO4CGLCkAFmhoyFsIKzPqbWPcqFwZ5IH0YxV5
V16vF0GgahuaZZS/jemVt4ARaYsBDTj3XPvFD0DTpdC51Ish9sSi6LTGUCq9
TkZXcJrgSvvgWaN13E50nYljKV3sp/fVguQJN8p+EW8QbBvwLxm4i3bLXK8n
dcN1kAwlUMSrBpRdP8A1l0y9ykEwkFGO32JXJFVG3GnWGSOm5tYDRKYFie+x
6LBGeE3NG0WRqv+Bsv6/rC7QDKan0rhDAznuDqI5IA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m7ZMPVfG4SrE9S5HdLeSpiO2bb3o9odc95ZiX4Xcr06kabJg/oUUpL53/yUk
o4PKORgycRdp4rMgQglZzLbam3GKLBxl82gUukjImbFvVPCU1yk9f97RB9DP
7p2sEDTYOH1HR0WGQrOWsabUnEA5n+ggr/AK9fVosmm1/JdjnOgm/iH4JPaf
27ZMKNmD6ADubkXgWwLdne2N2xeiuAA+o4WiODCmos+owOAXyrRskPlOawfw
fw/1lpSEecZSYgSLp474n7WkCit4H6qBHfb4tdFh38vy0/BhwR+NKPQt/Bqz
BmrlNCn23I0WTzWSbj1ZMKEeAfwlJ2bUlFxKRx0G1A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CNNG8qURIB7l/cz/igovAEzEgBZ3N/PFjOTMBrtaqSBWij3YkmcYbVN0VuAJ
jXLqz+zVoCxEZDh0NpUL48ldLnCMFC/UVfF+MrBZtwvBbLqc25eOLb9KtAQk
lKStYRtPauHeUBMdldixjHEspLdFE0aYQDhJVoaOO6kZ1r1Pv5g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZTeJno3U/Nc9zyeIvhJf/tE6xfe4kMSk56JrdCUxNzekN7V2kM7nhv1xxAiy
MHdWt9reMlK/ul5u3WaYSGJAOJKC06l94MOD1twz7oT36ZrgJ7dHKfa0fxlN
h1mPPJqxcbk28Ss+Gj2+YNJMEhsya49YOb8pUPLEve4ik2oqp7Mo4YeLy3n+
g9y01+2NhoM392OOiHxPA5oQOCGkEadMQuCb8SCzwiI8Qbi9l3WoXovvGvGu
+0cEX3nemuwhlUEFD8oZlUe3sn02ed40ff4M1k2qj48c5got9hHCx/QOajcr
RAOQzupXdGHN1rG0IvwsJaHbzYH+9jyr4nezFvy5CV2VHtcYn4p6/tGLsZ4q
Re3oZ15MbbpBRMNkfL3eJQO0HLRDCCu8tkh++vPo31jIXqA6K/206YO8dYZG
in93emMkHmEv1mJ50RObQtxaGL2+IGlx/dSNe/cwe4uLvPHC9k7p9+i0PeqG
7dKaVja0ECkg3Q1ePIPKyXGP4E2+xnJL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZQoWZdEQ105w5j0wKRO0hc0TdDYCVHg1NPSezTk0AQgkb6qjGHM2oKUIeJ60
ezbSE3esTQCtX5eX5ElBItRcM/MC0LfG1BRNblnWkyWOd/lQ7HO9EtjAZFAd
52lvUb6wcNeGcJ82zcbaKQoLai+LQAExMftcp09DtA9w5+jruTo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d6oze9uz2w1xeT4IFHvct4EDOAF7X9gG3H/rMVR9HjutZ7pg545V26dzV1Pc
CtUfegKkPCkt1bocUZSYDmKNoSM87orsoh69/K5O/1KhdrO9FcFPpkZBng4o
DqBPs3Q8GAhGhnNRAd+KjFBENV7ALFYS2VlqqNrlfAA/0OTstww=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 66800)
`pragma protect data_block
sKRIi4yafpBkScuf5EsZM44ADZlUavCSJNM6tbclkEhK87BWp9FmiE8X0+vJ
9X7DnKhMr7OLS1rXqmxXCZOa1N36apyNWiv9eG3z400L+B3rZIkrWRYigHl6
cefKU8HEZcYI/Rvsjh7shpUaLdMUYj8sRv6hzrc++0ABUYEuHpZV/T33vVUo
BvrP+dFAjXQHF6QdAw1ppJFqqxDZWr1zLte/wQSZIJdkjyGdldcDra2nnVdf
yb9ElW3Ukx6yjn8MYJRwuItKs6NcQt2IBNEkhUc534lkY09PlXV53Wd/kEI8
cXQ1PUiEW78exXaa44n/e863hvo3oe4kd2PM5tPgK+o/KoZw63qb9yjaj2qY
Oy9MHk+iHpQDEqa+t43/F3vNi21Vukb8FzKS/FCLV9U+lkqv9ZqhIru+TbCj
eM3YywB9W1Xbs6WncKJUeHFtSWXAvUs7yv/ZQsBG/iZfjtJwbEfnvYdMzm3t
fOO1uYvF/l3YBJv86nnyZZ3CBWUvayDYw5iEg5rPF9SZaONNCkDN85eLxWsX
d5PqOTpUjfrTg7o7GSXaxTK2l77FlOrIFctzyLbtOT8zF2GU5Oq++ZyjVpEQ
ekzu+QdDExgEiEcLlkNjkFUOtML+MxV1kdQ3moo9mrkgxkikU7YQBGUVa7pb
E8UIjVaoayKK0L/m+ECaFjO6XUna5CWfZux1oM9K7TbW05tlMoXNKpdLsRE/
tc9rI2noRGlMh/Djbimq6a66ZRWYqYSwYlfTkjCJEIRDryXhmZLhl0CMbUIQ
uhkSUmsFY8xkDhTg+PJaYpk5SnZU6JUQRixvhkUAPg1Kesme5Hvuww1dZZmv
+BFs6QP6QSL427x1IAAG0hB6swDnLQeyKm/Qzv+GPmTD3LuwloColbNWONMc
zvF1Zikm4OmSUrWrnc+94UaVzsRXOCOvw4Ux8aRNSWcx5LLbQbIRre+IrFHF
bGmVNUdlDG3wYqB81+gNsQ9mc1LS8quv7n/m1R4YFlup+05Gb7kMCF4xOwJs
NF/9vgx+in1zf2MK8sDX+j1eG0c2TLXqaECdvBeBzpswqcQ6sQ538aeFR+TK
OBv4wap06SJHnt6EskdQs3WqUSN0IgJZwXMQbfLF50Uam/OVLaGhyqSCHy48
3AASsVctKRtZQUfLgknE7eaRrxYqpbfQ5CnNXuYxMkqjZ5rHPTCeE/r/JAtv
R1Sorn8xwjvvAc1uKApYvJ9J79PA9JAaSyKG7/l6VfdJcJLxokV2t8TeHra+
aKA/edjNFRmT2bFv1xlYBDiqInXQROLRbTBFjYOTScZOEVElOeClAZm3P9SZ
XLDg30MDVa4AlVc+MUxfFlutVdHvobMmhvBrNs059IvjX+Kd5fSXvRL7qSgW
oWzkC1LRqqdxZTsJKmjQhqas0GP0j3NRcMfsLI7eghxhypVyUXqAxZMUPVFO
MRNG60w62lOF5Je1GVXCnnwAl+dtBA86hfCRGYk9PydHZdrF64SdIr10/IT4
5I2ia0ScIACNQ/PBqkkOWRkzL/3rAQmlzmjCxYbSIzN0Fpz7/h8jgpIu0yGL
md91LJabNgcoYUNt0As7LqMnJggWt/t4cP2O8qnhnvjL4uE2SLRFjse13wB9
e+ulPZ9FnLC46kd3wkjDraP7JDBmUHeXNiqQakd1+QvC+JrGoRUYkreSgOM5
pcF+Fa7uxiqscvk+xYfbgbH16X4ILhjhbuWmsfol4pUvQjP+pgKFvieon40y
Sjnz2xCZIRrQ7fGO2M7KuUFS6WzZPygWjhM+BVjXltcj6Pud1glCPeLjH1ZZ
7o/jCMIORqKhbaJFxZCIFlCUyvvhBHmz4mZQcPt+p7qnkycvBrKzhrwL++Gv
1vTlvsnxRQEgr9acfO7doMgahGNlurJZ37aC8rqdubQySIPWW46nXWlhvVAg
yDybdKX78jUpbDM8pKiPcdB2UTwLoRYaSd4tYfAciN2lBIK/jdc615hbyoQq
AnkVMhfhFZRmxi6VjNu4NGc5RYtdnBXIVoO2IQ7BFjG2roapF52FHL1dD8DK
HEXRwcVAH0JQrO2eiJqFpwE+MoE/uBqJmvmv77cvWMi1Zeq8nGAu+wTMdhd6
TKqqXsJxVXqtu90RAZO29ew/ygnsVImqHlx3vYk6uurqRpmMKjyvbtlIt44G
/Jgn/LHVzl5QqBcasLqQiw0Ji4Bftj5sR6TxIR8icF2gFZjBZEutOXQUyYkX
XkoBbTfywKwWnPJieSFqXfpGngZpI8p/oFPdr8prBiYRFeA0gglws2WhD+pt
NapaCf5zXXqlPO6cOnVmO3k+w2MOkS3IVD2Fw4HiNp1C4/hWRBunHZ2CIBnW
QiX7VxcuEo1QUjXsYp6q+XwbgpU0IpjzjkqYOaMcURYDHDPQvrrmASJ9TPh7
W0zXlWrdSZtBfEVV1fNjvVqgtVP/+uY78MF4L3Pq5zPNCwDDDdFMDA2VJHK6
+eYW3AOZPFk79EMsqBoUlnjvp2m/VLmPJ79PJE91DBPMi6cwgQO0+gzpb534
H9AayihwGp0RZ6/GdPSohSO2sRZm88ggiN55u/yGZjqw//G9W0Mj5DefEQZk
7Q9e7NoYrXvpw4/JYFgQWttCS2oobCvvx3k5goWjxD1EjYfkz1JhqdkDo6qz
0QjTSwPMteAQ/YRAkUaU0JGpWyl0gRhZ7y3RDXon7JPD09WZhYnQfOf3+iy/
xAbmqtmygJ6i/QRgEiM1AEZhORguTbxMDjU80BvGOqlTIaCSo1s12bhyuU01
TNu0FVR7lUA/1qpS4R0FiWN/Rn2IOrPVwBGoQ7HzuQafcI6SxQmXkDBlsFrq
H8YFRtfAIIVTbXQyDdnScZUGoguYX6lXyakAAh62/z1rhvz3XBjGLMweVubJ
AMvBDYCXPTrjD1sZcft9Q+0Vi+ZMfHqtdgdXAzrC9Rx6vAaapvCP1Gh7GQSi
hLmRKnCnjw8TonpiZKoKTyUhbSpoATyBba1updHkpnUbYmnQoqI0tFXEU+qR
XjPNqFJso2r9Qn6CQQEtAZg7GDCw1sIgcBrry9QHCzMQvC1ebSJ/dc15qXg1
z7Fc+9xn7od5MQKXUvflRVpPJb369XzD7l0FcdDCdNh6FWeQEzRNphK5SJMh
SYB3Xxxm7nIo7XsBS7DeEMiYs+yIap+WqGw8YLsWX6BdaL4HpJjCD1ff4af3
Vrgrq11DxdQTzZtYQsuDyNSyykIF+yJkrphsjcx8CLrWOcW2CWoWgIqDCVwy
cPL62vlM9l5C3n/QxNaXvurHnhFy5Jy1p5ARY8LEUsWYCVx3P1QJRVEqXpmC
M3EEhAyQGNbg9vUxbKwCMXKkfGYDb4P9hEGOcro8D2Qm8RMSM/rMymz/+fEz
nSEEeArufsnjGD9hmXnlzyEgQXdz4RWjGaljciviIvOBal7YlJsevb5dfZ9E
huXxi+rOMzb1w/4gl4h/lsLys9btlkmgEkGW1B7Bn74TDqYm13bMBtUJ3ZLu
x2g9IDXy7rAnOfD5uMKn6Jlv9m09DZx1m7sJdrEr8LAnSWd+15Q2fopj9Gzd
LgU1+L7f/ls7ADRnEfbmybMVEu/6J8z3HszrSFA0GUbPq1QpYpBc0jznIadO
ChxMGd20pIbfmMg+KZa4NZbsnF210/HGQcRW152E1xJijguHPl7+67ptM4+r
+g22hLyK2YijSm21rQB40imS5NdIhnIOrVGeasSyQeN3+/ZoZ8TD3AXspNN4
NgIEm/vPD0KHYkMWeueXDYfvsmiXpUs9GzhH/22CuWtRGsRTDc23wu37osx6
AdK/NC2CfSHskFWmVeC32fd3zRxjuxDgTkuXF051Sv1N/nu1sLxZ+/IUDrnL
gCPbqNpVcZ9VWTnE0akPmDKhbZWmZLnpnWRMzyPUPFiCLo+uAaMVlX87GPgt
jkD/l8DeGwj8kaJv9Lfq2JqjlHLUyuf2jcIchvUFXWZapvO5iAR9Z8WEVuOc
XbkZByJX+HYl8Dp9T5Sj7hW0mmPzKyvq7jL+ANmhahbgWcVtW2O4qdgk4FA7
Tt/21P7g6aeymsyR2XKSWJramolKi/xpVfteR4s7mslQngHc1+T7Z2jY7/dN
wxxisONiM8BNXvo7lADidX7AyO0saWyvnc9uLPjTGu99ya+UBF86MpIicgdj
yKDMw/KnxRbWTDWJG+3a8LT1Lo/c5R6zFdqrasLRMORKUag1aCIUsQlA0zjq
hOli8J6lpWNhy2Gtwb0Qv68UgBZSPmSlvIeafQgqEEEjXVksu0rqhLinloCR
2bnnBobxatmRghEV7BQB4dcd1ZasM7RjukchaIkHRhCOSEA2VSeLE9V6W4dJ
Bj3TjfrM3Ioa/AZd5tUynYYOdeZDgkPvJCjbinj2LNRzfBPKyYCVgpTwiIes
yo3w+DdTX65TJLgrlrPsQX1ekrZzYbCGrKXs6t9okQ66h5sgMIubwnV4Qc0l
y2r77ab2J2tMQmeQLsAnsHJgnDitXUF36krt8F8QgbTkSJXkgvVBUDS21Ad9
jMeOjk90MtOrKdceY3WKKMMf3ZVKcuE9HNVr+nsJBao3UXR3ltEKtYUn8wN7
y3qUgNA4s8f6Z+Z5lU8XZhEL0Nr5xT1GK7M4U3IyviGcaSga6sm8xf9XHxTt
mS8b/MtPaSRkZnY4b8R9bexL3525BlrkDmjQy7VK3YuKi5sJ3lhaHbnOmxPG
GG/67EYANhHt4n1LukOFEuMPrR7Bqs4S9q7pL7BC5UR1o279Hiem2NWjgZef
5tTvb0lt/PZg9wR5Gm8oe84ywCr893465817+I7T7CMeZ8cxWyBogUrYjPXc
ZP0xPiC4hDgT3iikS80EDZB9uEJJBO8n/TRwxZ6Xui++Wf94y/4GFrFfS/89
vbRA1BviQYh/xbPn0+2ZN5wfPEjrg6boxK1cxL2OTuBjeo3e65Uioy5LBbJX
BRq2RZc6tW/dPUtUaGuMvsHwbCwY1pLNGEf2CBpJ/fBtW5sG2W8BjhTZhBp5
/P+UL8rTqB4myhyWBHEXE53+BAe58OYuv1d1UvHg1jZf1Oq9R2ufwmSGjyft
BICoIL0G5kVairsQ11riNBFB4xK0yTxmNW41o9zyVvThwPkfmw5GLrVVxAKN
yKf1dPHnqsdwjFPlD6VWWe2mwl/evsQ/LHaQr5RE2FSdaJzZ5mL/4HqWMUPp
boePTnJD9/mKrpmdClUbqfpE7M9ZV77Q1Yj6x3HuPGQux3O2k+DsDF1evgku
K6ksXRiKw+V25iInAdhZC4j7nKBOxit68MZB7S0bbP4r+f9yj85QM/epFm5L
SIu4rjYyBzEvgpV64ShPpPtwTzCzlxAkJkfM/Pdp6J2RjGVjcDHBxARB+e1p
mgZyFVIyi7nHnn+iTT+kMtJsiU+VLfVaYusKcjubD0R+sG3WaNn6NPpNeIlG
oAIwfIkCfixGAu6HO13qm7HEsvouOEGNWs5ZUxJysOuqAxp52lNJX7mmbrhT
OryPthyDmg3X2B6Tk0NaPEL38u2FQKJRHQ++ra/N8ZTBSpT5GRsuJBfBoMDy
RSYs0KUDyBtu5zDAES2GkMuD2q/HbY398BvK/Ygjmdk549E3RAJews9W0qnE
H+0rIEUm6P1OFhiXUhLE3X53FP43nP5aG5ijcevgHGQJZNAoOHk6mKQ4H3Wj
SduMVNQEjDJqLXpHBxscY8ceti7+kY8cFXdoMbZZnIy4skefizn0JkDgl3yY
sEUuTPJcTYGoNVKf7DOlUHH+o+CNN5fEBmtuo8l6ADy36TcZ14dtTgADw04m
4NwzPneQVMiPjhEUub49NS0kgbabS8o3VSKG0PaU3jKSR8TtEiOzJsGLc6v5
zNxuiEeHR6pucVu0UoXt2uOxQIBkHJosb2fDpsc4HdpSMlkymH2sOyl1AZOP
BXU/oaI4a0/h8+436OoOaYvL1teLLOWkuSdTe5qh0i52caaAtdq70BiU1AIm
oJBAITC59soADU5C6M9IcijbDvHYK/nj4yP17E0C3mXUyDhd71eyYnOumyiV
xH1CkntuEXkNp1dN4X3CxGlDpxUqnak/lxZ3IXkCyhNDgoExcPdeNIOlxbmX
YXYmIG65WRN2JCf5w1DsX4AX2UvU99SpPIvVW72fILtfMAqG1phhDAmLaZqM
024CMawZXjulGhYreUJKWLnq3nQCuzr0rT5oA7DWMr2lLTubkyZl5t8zY6FF
GBQ3KpxC5IJS0B1LaCgBd+3tIDcFPThUepQFEJRmnFFdJZOY5c1VqblGZuVh
ObFpWeQeWbGk+TMs/ASIYFT5Zuy7vV877XyWIJF6rNdVauMcvM9gbG6Eilve
0rAe5N3Kff4XLmItB4n/9Rd1+DdA0sYXRQCbYG3Hs20UqzvEbVyVQzWOuIKA
PVwwFFv/OsSOBFY8e1I99J8rqaSQX3/w6LeL7GW9r3WU8GGTykU/eLix0BXC
MGFmB+iHPrvw/5AP/mhLBc12Z+n/MdUcrYsoeqn300M5Kd+20w6fNNWJ7I9G
R3viQFrNC+ek+OA5e/KF65PTQ5qX+dkI//8tVLVToGTP+5exgCWs1KO39GdW
/lHNqI0gy7Cfzf88iqNJShj4yd1s1v02D9eJtUefZkGVO+2deDQ2huImXUnc
9Z7a7xXpivAb8SP4EQeBPN8ASXa43B+tFLWHa6Beg1owKfFgE4Ukd3ciJX67
xYg4KR8RsG0ccss4nIsK1QhbeZJme+t2wGgb+WdtO1Sr4mfepTaIt74Hhym2
P8vVDj8jSzyfD0tKeOe8xrQ7bV8IwlxiyQxqHmzxIlFIpK1BETL490Ft7q60
OLD4E5ykZosvWfjgVyPX8dlGwzGrJ/vA4u5sRrlrUXH5nqnxJ8f1RtKCjlQu
2YA0+oxQdEE+loqGPAs7FAfDC10QHgRpesFlVGS2r6lOBDpNfAbv6xNKMq4I
N9PfrNCpTrq/p0uPBztCCtEesZVec47DrSYfBbm9J8rPxgdX9jWCjyonkAaV
5LXEmbDvgMGPKhUXPQeWSR0qMDvQpJaAt8oYRMBVt81iEOp0YrPihM8pGfXe
u74xSjG3eh92LES5Zl7YQkkaHiyJW7cXuEaI2qF7yzxOjQNbjqv4d1PP54q5
J30s++VXkRby0QQyD42Qy8rg1xID9h2PTUEuJoxAp0yDZIn2HYb5xJfpdNXo
AwXNwENMv14ktLwUoRra6tWKucjqmKa+N0cmWQ8VnjQzOcbth9U6JRb1uzVm
UPBqLaQ8HEvXVc6hPiWWhs0eIvjbyhNxUAtjUoFE5CVNdr+773AufaPci7c0
ycQf68qTZcs5omsf3618/eKBYylBpC9KA9NFyGkhog2BGBmDamDPzRKuBBk3
jzSPdHvzU3KsIy0iKCDXN2OIq0FvvtubRCgApAKZLHYjX9mLE+Y36yZAvg4v
xcSTGgytQOa4Br1kw98/PSGtricv35TadwkIZYuX0AG8fX1/+iYEKjWnbClT
05rW+sQCpcdcU3ZeuP92d6v9tUHqXPZ5Tkz8PHm55C3gIOgPpf4ndA5o7d56
phNSGtShhzIubuz1CM6PIfGgLHt8JeokGiMlAjZYWqsrSR1YwHDHXuCEcZri
8mGpACvGTPXG40nM9StT0FBNsmpP/2++A0ms2ZBu5fHxxFBD1GWl3MAR5bzC
bQb5zaThmCzEw2rnJv9LuzTNT00sJXozP9KbFZcd53KgJbNZIqX6YDny8XGw
M/IMdMYAkn/exmkPgeSkmuqh4l0sGsYBp4bPuSTGOLRqwb7sugO1dmfNF3Vh
GmWkyn1GnmmU0pW8BNfEMgyYV9w4+3Kd65lplEOAqw/7lopz6gyIOoDhMDcr
ofBVxDXDFTQ3dP3LlR1Uo1X5QFsVzBKDiw2A6W2l6fqmtO1o38/2Wyl7oMgq
Ra8mHqBgJ0RvlT5E5l8J3sgSu85kMB7a7Y1ZK0wgATpVh3GOHxtAkD/7p8ci
rSqt10ms1JynyT5u0zm6nEckRJit6XqJS7v2jaSyMnxj5Sq5chwWl3v4Ka5+
vFYKw7kO+M3PXOGJY3hJTgnkisYfJbJAWp13QshsYgPN08F6/xKDX6u3ZO63
bnkb5Qj2kB62qmIIs+C8hPRWMp0KjsjKvhlBYVQ09JwXztIKrAeeChv+a97i
Iz9OXz5LEiA8EM6dTIVGKTI5fAqQwG1IqSavOFVkSUMyjzknTE44sG84dHYX
pOoJlWWGqxrd/jjGYm2/yMeMh3yZQO0A3DoL3osyAOy2TofWtbEDk1oBC4up
NPhB7+/Z4tWXegi+co64J6mTpqKkGxYFY4ph1wu0XK1rhejUQNWfgbt+ovIi
uOYIOKPDJHQwZce7squk1loC29D9wMvaGlETfJxzuDlexGuglw1SCE+KKH+o
hSnRzUYtAkinVoD+g3KhLU1kZfhK8riyiTdT7w6ssnm2vdoC75G2twnOXj6R
TMIs6WgyhX09NRPe+92Q/bTLP5nkT3CV1791958VKYC9qXfc8LwQhnBuFSLQ
08uJeTxpJw4RW/ZX+ZxMpPy6cJxjmCCoYYAmqmd51MkNasa5kkMQeMKH4ioi
VIoVu9BeNIO/ozOsom/ogu3Wp8eYGcIozpUIbLMkfzGypS5EMnRGsy8kWx6r
9+dZHK4CcXD5UMb4edFz9ckdmiQKy2Mi7pBZEqoxdAGi2etVysMYMuPRZost
JKnFCrNXJd/bRavt67S/XjQAX9k0DnAwlXj/8DG6mikxCJw7757HVTImtWN1
2vTj1IcXR0ZhwoMvTR54P6eRqQPL4UfEmsQ4kHpyVJ19skv5KyUF5WvRA4Bx
E4EsB3degL2p5RtJvNuhV8EF4+Q14DchORpiv1V3QOtOgJN7EZUpd0NCvruq
Z8DWCngMjo7O7oXZhTMTCvNX+PwyDXNcUOXArGahi+OKn+jlMQ7NwsgZvxdl
JTYGZxLmQFF95QVGZidDJWWq8Olmo0qeuoc6gv7QWuILdmAauE96D6tMPrN0
MumQr/t5jd6f+CaAMjIIKVICkIG8aI3oxYa+DLRLVMujs800cDVkONbUB4BF
y8joQix0HGCjEjKC1bkuy2ybXrI5BwRtPMEwr1rmzotfZOD0zqC2oiS8xD+T
etWYsqLK4KsttTp3ostmBEUJVUsQsBu5A0lYsl3spIphe/+re1vr0D1fCYxC
OZkxla6OPbnpdXcpzhIuoKwd0e0ZWIybACLjL2SEg/aB8tcn3FEiaef3CdTH
gT3/PAvU1Onm2sLNvRfKZK5A3oR888nwmkAVsu6iVAJhiYQmJ8x0xf9GbO+B
ck3pY/CECV4qtIa1Dr6FYEJOpA9d2bK2TN83HT3tI2XLZdSErgdgxZvOEo2F
DTSAzYh73Av8wVqjl9VDyJoV26D7qGCENxnXQzz/5HCyFstO/mSTT/NI5XCq
8hgKr+6vkEgZfj6jveUorp0kqbvF7x4pnF+57vwwN2ZwEzh6NN25w4e8ImbO
PvkbnvuUWSbukw70Woc7QSPKuuNVC0SEJlL5ma9V8KV+m43K20f7qW/v9/F7
MhYlngLX5kwfiCAJzlxYCLy4TEbzguYUVo/FEwk8i/edY8hOLyuPT/IaSsjy
hTqO3003MJJW1sVPBiMbza9niMT3WGLDCVBbJWOZ3AOkT/nyp2VYFtci4/BE
WrQ/+ct3ioZtR0mAlNH9rFwwb7Cf9M4kfIrpMoZIM84ZybeP2VKEkFM347Hy
YCJ6IV9H7oYsWYr3XJ7I4EJgVy3ftTuNWQ0n6Yxh2ANPQJ3Q8qRiAlwhaqIw
18tyUm/6+uGeXp52PPS99hl0o1sofpjNNaryOGVuQ6xkbEGOKgqs17jscLtr
b2FLBa8ceeIBpwVv1Lsy2uCxAPhA5SO5NG4PSehVmq+IcZAleY6GdeivE6ZB
uiOLogkcTv3auWfETKrz58+fJXg8o8naa5aQzavNm6Blc/Y3pCwhKIj3rW+Z
frYJ+yARorPa/wzxeHlHoa0bf6rQ7X/9aKYMHKk24/Qc0c1LjIxisNKK4ZdS
7u5qkD/P/wKQogLHLtAsMb3RafhlsEjHVC5sXzFnm38DJhqM2+emR1pykdcy
ZvUBXC9VEpiKo0kcJoGR1iRWkoBfSipFtjkyWg6r31F09REBnLyoaLtz1SG7
fkEqCBvyQLZmx+UzIfwM/4CwisCN0AyXWhwiQstriJGMSt0/PEsif5hE6e7e
8PUkXv9SjGQwZZcTONmsu1LdvTQs3aSOlnnOoNSOqJ/1D4QnjaTSDXyNGo99
EprY7839Un9LgEY18MAAQiiOutFs91sXkLw+ZdtgvKDcGy2M5/VuyGdFNc9G
/D6awXUN64GAR81hiEynGu2Ooli5i6I6Z4LikhcxZC+SwsRqSpR4zdNDpOVM
pq7Wb6xGr3agGbwP39IKoEalb1JHO/zBbVz1hM20cPrq25879ommUkEbrkxj
1hFSy+WHJ8YRyqB8MVtPU2bVGGkbNy3u+Bgn2V54Rr2bH+DB7g7+JIH9u0xN
Rwl7DiUR7EIvoZxUhGs7nNqsmmnGzjBUdcD9UV/tXo3ONc0Buj5V7+1qhrJs
HLtX1hhdS/CiJuYwjOgU3vdb5uxYLXXNK2ntpW+znYc47Lni1VTbAVh++P8N
0FPO8jebv1qqm/421ifgmwVgkWlfFqLrHnmaKGGqSgtHj7zIniUYZQ58I0Sj
8vWn8Fk5gzFjO893YB5q6x7PX8MsnCQTwT42HAdFCDQ+Dva5G3/uBmEQdAFy
ofY61UKaJDMzmPQMAx9F6VkXh6P8EcGNL1NW7qiEsugbdhLnPC94ARhNYEnk
FMAApfRhyDYEe0LOEp7cbyIc9dLbMwhqUvL1W9imOuJt0mFvTJo3upCIhBXd
Mplz9jv6DVinNYTM34/0SUcos+bIurSq7ZJkxqSFzUBzlfe6VaMCLW27z0lp
wld+xTxZRC+hq1FwCz7hhUGdFu1jDKwIiPXnnIgKIl/+4Erhyz5RJvfyt4aw
+Mn2Na+UV8q24C8bqVA2h03tHYEfm9Lu7OYM51NGe8/xLG/BKXMqaDcYetFU
VGfE5H1H/IpkRtTuBdEP+sP8YTaDKPPTeM1/8QLr2AtcsxCW6TYlOeKnI9r6
2y3JQil1x3Y3MeMztc/J3Q0BYk6fn9RFu5b98opFRe9g20+9NOBWBksiGQcN
MO+K5dwHJ1oByugljCZsi0emOZaIsjTyqnsoK1rT1ebMIAq478S0C4hAe87o
EitjfTvA30MiKA/SHc9yH7z17baqxKV96SQEU9+t9MA922Ne2sRMQ44xddox
OX32guHLthQ8nILoVd3H0YMq7D+6XdnPrNQ/Ibn51lCmODg6lFt0BoHmmweF
z27OPFDPhHjlnVDuDfuGHrowjfQxefJkp1mhil5n5YFFhy5+LonZ7N0i5zQL
TByHLIj0VyDRSqLt28MPX1mxIEnb3wJHsxXD2Q04/bwoHwbYt9GW/kwUA40z
Y8PoX9VsvZ2XCYcP5QTUFrKxy9HqkdR+0CJqKAfJ8mprXYuj+QNlmdyX1wXT
U2HHdH786vUs1N/WsWTgx3pEGzky4uHfrSybYRVEUkRbAnMPAcAr/16aIK7u
hK39Er3Rmy6XY3/AM9kOIYTMQ95U8ic6LEervpd1vTrt0OgGq0bq2eh1QCUF
3bPMnegy8g0cpL+pn6hFNBmMISYek5W0dUh3X/vBjCB9tTCdsflDfsCmCBX8
FfvAdtb30SiGV0wABD5fEkRgJIYufOda3tr+E1FlPMOaI7J7T0A50QKc5Pcs
FuzKAax2q7M+i8LvD8ExJmXL6p9EG5VCSo21YtRHIU3L5/WsasrbYKC05EyW
OTYL01noP1w1as551AVLetMNsdJ1uK8eRXlJG8fkZNpmkjQYdxNiCHcenK9A
d4VGDBgngGGw1bB9YxMISILZnFxVaQT4WXVSheyZzeiZ1SOXP/GUEviNZHTI
g7wv8BWRsUfl2nerejfB0aURVXD/39dE/Hz0EZkDSYy7we7s2o6qOIAr3Ceg
wkCkCW/pqONkT3mTrXRgmEnC2Mtnsr+dqjMdcNp8u6Mx6dN3U9rcRyUDxfNL
NlRsVF8KNFkG6hI5qy/Wgqv6tIdl5nA4KLIdrMje29Q1sblsGVmRVF+Bs4td
rmtBXGpGFSwA+k9+0t4OsJTB3oAzXJ6rwLqjJixyCo7e+N/a+qsrB36ay2ke
PnjOU6gyXsoGbMXQA6SU9JUfOUy+VShaYK6J86EOl45PONx98zCkpQv66TnR
rXoUfjZ1aKFLHYIWJxCWUKFj2bK/GUtQmDrLhm1D/P7SRnW5/P4CrDEmhMjZ
D382/RUOz88ukLp8aHV8lCSrJpWRsc333NbgmC7d/odKvxG/T5fZ3eau0bm2
ejHCmYEYyKOvEnypdwIGQ1tt2JUIc5p7x4lcWY69mnSC0WiaAPfWD/z7uOgF
Yj2h4U0ganphap/Nv263k/sO1T+SqgHF7U8zvsHHUGhTmHiaAVoLP96kf9cb
vP7z8emRAjaNyPLbIvUPg/Etw89QW9GP7uDTq3Hw5fRRhmB50bge+u5HyElg
sOpFme2R574IznDGiCU1laaZ18TzCIGMYccSriBNEZu/c9jQXTMHD2rji97H
ReBbStftiH36Hnk1XpupndCNZDZVUSySW6Kgzb1nF1v+fAnfJJLYVVlXG4fc
h3b5CdMq0L60zaL9XIiVRBt1uSWuiDPnNOXg/BGP/EygNFCs0gbwjokEU8gx
pt2irTX+h5zJK326cRoHU5sy2Zp4BuwD/dGdrxoqLp7bhXqk7UsreygZuIn/
xnWCZ+b/TDnOta5+rKbv35/TfnDeaM+JSbAWBqwQz5LADiCjb76pYKcYxfO2
Cz0SUPLhko6S426eydBaqaqSVVB3H3zoBxw/CdWo+E8HibIUGfpt0/vt241Q
AmE76VukF07Kj6Ie78OJCdv2w/4ySiPYN9WFbNecKOsZ/GoJuvAF31OiA0To
t3LqKcRuEVMPRmcE8Cur1f4ldQvhNDgEu5aR4jm234RXJAdremi3mJa/Rxj1
+xvIt+t0ju4DNl3dVMk6hgfNUcWbVNJB6rO8dYbrER/JQEQwG6xRCCi52Z9Q
Xq6qA6WsV+ffhxdi52Spiwb10qAGs+QdICgECVOfJtSDWQ4olypvCJuOovqL
c6uima6s8rShwbFdGEWDzMbfl87w+Yg3P8c/dmHJ7+iH9/hLnRC9UJzJD/0n
RNQAn0CFnhvOT5R74OddqtHunDXnRhLAk8R7kHnLa/HV+Rhm52eTeHIlGs5+
AkwF5Poix+CzjcJsEsmz1OpR9/KgjmOlN7sq0qmQcUANCR9vLcD7hDnTcpGY
8UK2pc7escfAqUrYvyp3HNCxwDr722EAgu6IGEFSC+2B9lGHJW1axaEbEyjp
2FLGnEMfw8P/XoaCMZMB9lU1xgmbwg+rRjpXdfDaBjsbEPF0DipQy0/YQeJB
1ng9CMbHDIMEWFnCI6ueLbAldpYBqp4Allh6ppCONSJX8iHx7K8jVKehr5Fr
Ipk/5qMwQip5g2+Dsxpii+AjVNKhPd0b2VYzcQJg6kTHqXnxN5Rlq0+SzfdE
e6AnQwcziL3v1RpqAwy4FW8a0BEaHES9KdZPFoQYCkGMSSu29ARFIN9Dgt4v
kr8itJYsWWWi5DdEju/azF21jsjzgivTh6Qw06RYQLp0NFpcEVUSG4giOmhl
uqAOSUHuOXHF5l1u8BDSxxEMHCC3M1nC4/NH08eWIOiiFe4bojP5OZHoNbxU
U1gxZV7IHQYFhzXClUjcfnjVj2pnz1vO25Wk/P27g+ndPSKMVokAhLePWNxG
uX41OTFjyIKPY1NBCqQJgjDlYdwsJnYVwTShW85zq+gdxsHOjZ7vRbgYXyGc
h/eLgJjIXe8Q1c2dLV5P9kfSjnYZdHEGRJ7D5jhfESykgQtPTaBwA5zh52Hp
vnx+CP2ll+U/oMur/7HB5iSOkz23uLJpSpWRKpYfpiImSHnrOFrqnPlajzu3
Yd+tGIQdAYQXMo0wWXi7MeBDRYYXPE8SH+PuYL4QHU1PkMBpHr5P+t5sGXV0
CBNQGPPdHlTeuHtu9y/lZF51e8UMvO9VE6iYlYi4udkJMDDCW4H+si0BsTJr
SqmrLiT5q2gBO+urasxmw8M+Jc6eG2KFdEcmEayUX6z0M9p6RK3+rPir0fKi
HUMv7MfqBLbEA0WgGHYiL+d6x00vIPVOe7ECzYEwWzCsYNDE+vepoctZiU3S
hCxUany5dkCHCRxHo9BDyQgKdw/VdGdOQcthHXVC3rOwp/pbLAqxSKscaFke
dQlF+JsJyFcqZqLtVOsnKwDzA6REwFbusHd8H/O8ex6phRI4Rf0MPGZRrycN
MEkNVmEs8Ve7J1lxCNCEv/2viWIq7kNxLDFMUfmXTGiygt1wn9UpmYgoXTpE
ZLqiaWgtnkxYSoOm/kBY9VWh6Zr7ZpUlBoR8SLuJsmuJPBRwjxbMm6+Sq7SM
J1Jtz+PLWmi04WDv7U/uaOTHuilfsYEON/yg5nKm5IFagCXNvF81suNpXbZW
PECNQTIF1ZNYQhBGzzrmhFVULARNjDXDo26eS33tllEW/bDMsql0zayve2Xy
NY0idtC1WgddLc+fVG5DtOkS4HyW1xI9+DRwkF6b1s+Yizwud93ZhZxz+Z/2
V/HZ2+Aid0mlKpaLtDVFX6lEUWiJR11pXVcu8T0YhVM95M12nGmo6UdeLUn4
o6mQq3Ux9ZbMNeKR8ZcKGDOAH2jx2NCau60nfHP9Di4oK9jdVuYtukYor0IR
N/R6jbCvr6NMVm3WKWvkRnR7nCj/goYDUcN2gQRCuVqNHw+nS94e/+wCksLf
TuZOPOsEVAypA3x3q2xcp3z2he/pEWR8bC19A66HBy7bgieE6xysJwt59gsz
URvWb2MMgEjT+XJH7nkvWynFogexqCFkca6Xh39zor84E1qYMsikyMtsIcWk
hd6rMhMXtOfeCu9fPvMbDcFK2110rf5kLHJKpi16vGDyT8PDHKB9uSh8eVZ4
lecuF5S1amdvZVcx5nwx1n1+femxKvcj1N+qAjHyvO13agc/l2EfIBTugbuf
UBCJ6p0a7TjsSc9gUMAHr8mYJKNew8p2LaYxRNWTu9wKAfqFoYbQKis7feRe
nihEafukSNnDprOu6PuZNndhrWeK1bETGT7lCPTHS1BCLB1kt13slDv0LTCN
RiEHheuzM+zNCdkpLAKPxguO1WJ6tfsDoLSj9zglSq+RuYr8cENp/+X3LL49
BJ3yeUxZm7HQZZflF8WegCmHv4g/y9OEumA0T5bQPUFyTHX/gh9Jd/jaIiPi
tKh2dctclVAN9V6xX1yx+elWwetjzS6WrZHBL8McbczMcdc3gV/PNJp8JSax
mp6u7Z54DalzAqnC312PZz1NAyj36iRktQhgeU1O3a136Ra5vYtWGwwyVd/f
/WDdjmbRqFwxKe7qTPunzbZulDmpnfl9aLABgdGSKhUZEEYoRAJnAFCHpifI
JsHwnl/xloSq9EN+3GoJHhmhhgQOvOCSJDiDzMxS8T2jZPQyFxsJ1F+bVP2m
DXMV0VZ9dh/9tHHMmlNOvhLscwl/2jDbsz2vNCF8JnVaY/MsNecTDHQ84eX+
0BXpy1Am6xRCrNPcG7khwTlT7jKj0c7mPzBHMtjPBYEAnT6lkWFSgxH7k4Fl
ylDpHY7xMVPjDXNUX3KUcysgZaki9xO73qovKFM3EqZtTCYf6ub4TBVcbwu+
Nyxkmi3PDyNpJEK1Irt22wrk3Unsxokmj48XMXmkqSXVZ6prcyZlQ+1UjhEo
UMyEb3gFcjjopgek5tAxZ/Lj27iKYyHBBE3uj7BPze+6oxs7aTVDNR0sBJo+
xxlmS41gScQ/J6S0mkt7OdQORw7zyXnND3/rjpEaJtGNTN5Vxk7y5Hv96Zod
JoAGN46Sg7mn3kBnk4jmQZaHXbak6zwJxghaHLIKOEZ9oOziKu0eD1orSPh5
g9zddE4dvXd9vWEI4mMx0s8MSJb5ghSTf9w4gMKXk2Cb2QlC9sVLjWy1/jpw
v7ibtBiuw2g8gPglDysO1zQ/3cCRkCHO2c8gWZOZUlSQ8GWxxJiuGEU8wP3a
zoqAgFm5MALX0ueomBHIfPZOMgwtJJx7qvhC0YVwhE3Zi7sMunuTondE2ITC
hUtBFgLR8KENuar9AF0uLqoQ0JpnSS2Qitkd5Vh5URCslbQgGeGmlyBmiV8S
Xnu/G6pH8nb863Hxs8/Y23H93iN+v1+PBdo2quc/2GlUNYR6OqzakKI8Tu4b
c6EBbdayR3hiZ3DE0ZInF1XsPT9GauCaNLHL280zJL5kSsmzQz5jFqtsp82q
VpyypdwfyMX9UlJW5mo3zr866qHbrtso0zKXzCzw7qNUc167bvJ8+LN1gXUT
E30ej7/SIYBrzun79hWdDZuhmtUWEOMPup9tqZ9dzs3LMeKSj3PWLoQipPOy
GGgbZxrLQUIX7+IIbNu3paFWOMyB5VOjSWuNOI9KMynVPm0btQLWU/tYCMV9
1uSyARK/IP4O3K/qY8rWdjZLvZ3vHquD8NIrwJ78VJrL+sHkkQWQZCFhK842
+MA54tNqBZM0gF71Rdjp0m0z5bAzXFiV/+8VVUt74kx5Q/QVeyflgmd3fhnB
izxMIwug1SG4fXEBQlLTakooqv812vnkCJtP4xBgWRnIeLJl1RKi5w/kF0pe
qVdCP0GA10dSznflv54PJdQsgOkI2rCpkYrZ5sVUG/DLVMw3jdR6d0Dk59kl
i4RmZVQPqdEFOmZo3NVZvIvgmNdQ+A2vI7dcLmDB7mR5XwQTsssFR9KCj6j/
MmSzi+esKVJSnjYOw/wuzZTcbZJJBP5pNMIrtC6k45+JpzXxc2JoKYtuo7n4
JTbxqAa0iKYGdVEifpYxvbwC3tCx2JQHiAnC+dDs63PwX4mUreSD322TWhq0
C4tzPNQ6GFbLphHO9CgX6YxRJUJeNUfW2QZwhKIx+T/grqdZvqNlZ/YFqMfx
n9CrPMFYYAZ7na4lcO59SG85mrla1dEvwziiftaGsdjqCDAyxFJovgoCeAil
5QBkFJ6xmYmB0NWCDvCkqvyqiQr37bga/rdqjR8xaA+kY9RtMEqX97O3azyV
iaUGoIbJT9Ts1eKOe7HT7qm66nPE2eOI2q+3zkJUWx9tZuRdn6jyled9D5z2
0Z/X/7JU0XB1nZ52yjqz10ZGnjpQEZfjTXdDsRy9zII2b05zdz1yq/dqKh6L
hl9VFPH8l5lXfkJtY9f3xyyGcfeCo4KZlzbqhSYfs1ipnv97Zv+ed+LR9Lik
ed7/L92IlBMbDOJ+oKys2v2aoYk3283FSnvOiuwEkkhkcYHZhHYe1h2fo3gb
ua6j5v+SzF/lfK6eiEbjRg7f1zazr/5aywoa3gcYSc6je680+4G7+7zvqHfa
SvRiVlZ11gtKubncsE9/2B2+T+KV8gzXpmq+iYjdZLERnEebr+1E/ENrTAhk
aswm6VyjCipixzdvDPYnLIlkrGhkRng5ZKm8avCbOfhvTWHaDeceN8lqjvqJ
pUb1lBOMWifE8n5jXxa9+y4+AzxZ7uatb2rNmiFD/Wbk6SNYadAN16FKnZ0T
DP/zuiCDE7ilACgigDL89X7vZ319/zLj3jcEQV0kIvs0lZ1KSxluDHWqQdAA
2m1BGD8Ph7qVGlonZY6beMmcqKrechBLEaKV8GXIyVdkblnEHBifmjEQ34or
Ou5tkLqyN/zwU02cDHGaSrys3xCaYg95AjccmNmNpz4pXS3AjLy4k4vfR3JM
f99MR7nCVMcGWiq7ugzpCuyCLQVdg0h4JbYTlm9V/ShQDS7tiPNyA/GuqYH1
mNLNIoqM2y0epfKo54M+GFOAy6m2uIaEyBm+UERSKlMgOLRSrRrXkGS9U2gH
EV5dvsjG3rWJKTu5rbs3IRMtZbFbYk0EOiHP0JiY2SxyPosIOKAM2XvwbnwV
9cA4mUJ2gHjFuaTwOuYBlSL0BIZsYscIq2z8ce2eqUaMPPSiZBleNB/7gJgL
TQJej3RlsnZTNyUicEHIYuJ9EuFDAywWUc7aYDwCmZgDKTHmh+6ls3IpN3ol
YxSTwlrDQE8MPepEGOVhpV0UKV6eRarFJqQ/HQClLqlKbHOcnki850KoGMNv
WzV7A9bczl8Fi+KxizVK1Hqq5wLsFNWFsRTt6DtZc2c8uHXu+x26s/KQOU9Q
hH5Lyk4CnXR+umldzwfgeYDt9IfvzZo5+8Tgx2Z1YfulNVD7qsqDeHWYW5WA
HI86vTnY57VbgVtAPMGK3r5wS0xmjRVAG7WNBcwSw4QSlRm6y92dgJpBVIcc
cDyXN5a/aOvFIqFebpQBWHDRpX8EcYtAIfp2uehN2q4YS+k8jH8zOu0diMCo
IAa1LmBLro0NrF2YO83RD9LMqgqx9BiBHizpozffKr02e+GXUWQyZIwTQDiC
v5lBKnlel/p7occVhLvHhst6Hxc0eoVJMlH45veASj6MY8sVOoZ/aLY10r5C
VAjs5+SxvFLfobzVRb97fBBiLjvqDwJGjpl06GKGt4OgdnP/jBCeb1fj7kZs
EOI+aj3VAdokorOwjmYjRcSQGtoemkkcBVw3G1i5ZZyZVUtlcurqQNXg5Xcv
KGSmRLcBZTHGMZHdtp0XjwIxPJHsDspzRUo6VLvscLjapYblKNeVn/jvOeEn
4oimLvU+UhTuDBwtKAdmFCV6xiXPiBok2+C1QJBTzeK1LLLVAgEUN7RhiBSy
VJ1cRE2CEa4GSXrGslzbOdG1cCNX7mMpef2vD5QkAKjgo/DFAmlGLuZYWEo3
ZCe+5sM5JoU5VAeZc+0ZImqG9Z7plZXbnCSNYCas2ms2am7a3AVWIgqwWYF2
c2flSbuQVzTY22wlJtKb9dndudq1teaLuahO2Yfi8BkDZawYFSsh5k0r/QuW
dmdE6XyJ4fkS0ninhcVIYFlKv0t9hMeABGbpUysyg71a88hALry/0P1yGY7N
C5ZtblMUcGjDlUqLVgvuOP06Y7FK1cdi0bl3t+/OvepJSTOwVMpgK+/LF3gb
exxw15GcUUiIzMf6BWRkRwOQTIKHW2oUrHKYkv/gD94JkEl2pKyA2NibEeAz
vEpaIJRCeY8WxpdKoLd0+WHLWPCHUCFmZovJbIdUs1OSLfoh+SNxv9ognTca
wOBNbIMdbtijcpgCZ+c3HxxiDXcz8EzGTJXdf76p2RA4Lj0HIk/G2x5pur95
hDoEgoUJMLUMWcIH57j0u8o4zc+aZj+KFmJ7Y3iDPLhOqXo6Ton7QBW+zIli
D1vhh+ZJU1qrH34MDnsFrVN8EA56mGeE/0d2TlR+OyLuxwwqXjDYIRALe0MX
LZrMaoS1zYV1dLbMwBwtEsa8dESZN7y8mSOFhVqqpGjwS8mRYtxx8hCc7n2p
c7s4NoGxXU+Qsk/d74Ml18vnnqshcPaHei8TNiNJhGHDxDJ+ZfAFsfWKxizK
306Ix0f593f2kJag0hMI0IIFJMN98kB/iZGkkehuWx879QtGgUN5tIOln/LM
z9xXTzumiISCdsG49Mb4Hk9u86JZWfA5i/VpW0ZEjXzlHmj+Z65qHG+6GmgH
QTOYBv7UgEHVtUHRgfe/Md6M2isX3kMYqnyBfupTxego4I0bYELcyYWARCYd
qtXnEASjeB8MKkfPPtozcsV+eUYTooRTOrA1nyrkaVuy2KQ3LboXJVF0EbHv
4JSeglNIHSDLfnznYDxBmgqWlXfvUBZZGCWXPOqYWn9sZ6/Jsl4eKRlFUVc4
THMurnQ498DV1nQ+91AXosPmbxr/f405LQrqCnKtjVUnrvPS1KL+Wd67XzaR
85PwWbroA73xcYN1qj5QiOivuhfbMjuReW3jSt6LSnD0YRWs3Z+E+NjgJ7Y9
0yIsTtU6T2pkw5WncyWEdO3lmt7Ua9RxcOLtiGriK0rvPvDfvq3Kv4G4nY9S
GtphOw16DWZCyyYnEgizTqKax60zN1NPuH8o0RzrQEVcH7TwtmeeTrz0224+
QHMTEBF3PZGvQO8gbdDuHeqPl0AIMvJBqLhuEmRTqQHHvq/FJWLjywfFXTtx
+CTvfYywJrkBgBz5wRR/SKQOeUb4HluTMm6pQnZf9XCPMDLFrGdKenDsv1J3
0bEwyDfod/5yIf6h4Rc/lgp0O7WHlziRk2vtF401+1jwhaCWSA4skCMgPTlR
b80fzELKoirtNcUUCnpRTpyp91QeicpEFUR9TAph+Wsx/3UMBE9KOloZWROz
1Q6WNt286TE77+5CCvgl+dKBKCRsY8nWHrv8tP7MBMM6CoyuSg4AEHeQuxgy
j1MMkfmv8CFSvSl9myq0izQPmzCp6ECYvIZvZ6tgrwg8Nxfu/+FFxaRkhFxM
0vp440HYYK5I4dpgWYXLdKcuUzh40w4yfa8VoJNudVNn4wBC8RMaTBTF+9Uq
cBWvGclzV9oxjhyIvX8G0s16ez8dHROSIakHvwbfMtIyvFy3CkC/kVYkVvPc
n4Obgslf4R9TTKqrLrumhvDEP+ij6WCRqIXbrcpUNoNU/RLWtQaSkH03FFGa
pTrEZGTAvKHCo1UTE/iIowIgdfZs/LnwU+itYDc8UantvfXL25eScK2f+iJU
LbohC3NWpANiEHg/Bo95cWlGkFhegs6h+Dv2hlJB9palNm7wMKpTGNn8O2lT
8Ui2BsCqYrxKMcbq65Qcf16HqHVVXQ1SL1uI/LMItpNTlVplla+dVSktYN5V
QQlL13oF/hY/I1JRCzJhXE0AYd0/8DIkwVDFaHH2K4WGwI+ryXVQVRe13zNb
E7H8ACl+fWbLc7ZX0s/i6nY+TUWZbGT07VfUZrvCtyFBtcWHEb32ZHXOrO9X
DY+/K1qP61OMnFOMxI+vKJ4nNS4Z70jxq0NweC51JN13VdauvRCg+wqEp/We
gOJgYZrwwBUYbVCY0YmjHvtm/cd4kmXRpgce69EpaWhmLyD8oAumWId3glaG
dC80ElzyFs1aL+y3r6XWZyF2HCbPezEvveprAqWnph8gPESxH1MWVzQxvERO
ZrlvFDSmZS40ymxxMX9V8suT9tbhJFK0/USqWouhbG//A2CwsntTDi43G0yt
W/qti/sQMpNHUmI7ECvV24Ryoz9WuFYaQKpaEYos7/lM4pErkimQ1vZ5D6BG
od1ij/AHs38mgg3ep1Y3pKS2//EVxMfI3Q88HR7dxoDzOcgjuG1W7uesUzYr
+kC6enZndsyCeuy0l//vrJTRbjccnE9hKW7nEpTywDv+AkuUwsghMUV7IuMo
LVjUPux2WZ+4V7mPhr3y2C1ZmVz7abQkDmg4+zFTz3Gsaf64fyE4VVlXUJ0a
Oh/6MKhrylQCNW3rdEl0BZXskYXW+r9+g8jEuF12wuTLsunYVMEkLHG5xVkp
Oodfl1bksYUf8RDtDGfdU1cS/bBHeVmOD59UU4DKa5iV9N2bGINtE4+/0I8h
sFj7ftNze31d0SWFze2zYxAhtyem57HC7eG6eXddsYleQrRn5P/I/ZZWdjeA
lj9dWQzvoTLMXbJGWQCQCRzyym19VsbZZ0j59eibiG0B4tWLJcUAYKPoeGK2
ulD/hdhWmUyycB4oGWoATNZDqVjMasE+1uXqwTrfWdEdS+XIGJfkrr6EbK5Z
dWLQkWES7uV0pQMKvTB3UrT++b3XItAOLZOtGy35zUuYSNXn+99U41L6pvJA
BTxFU04Ck6XiXOS8pWRiinIVNIsk/Ok2r5sBsbO+SlNIckYv3xseKfEmzhJz
wS5NqLQaeDqLUa8xbFZtr1i03flaKn0TqkeZWN6j8k+/CU8lD7IugWK6XfDJ
hRXCqIitRUTaZao1qKlBYrUn9+XH3//9KW10+WtMogvLoAXkqJpHjzNvYzk+
FyKMkR2OHcemhLI0AON02jpJmOtsui7Han4UIKbH+GNJ+UyX6xx2RTU7aPcN
w8OcGlDFFONRe8Ji3ahT3k4BasCHF4GUKnUg0XOkLCbZDAPfdOTqgYIQiiTr
WWQn1B6T59uVCIZQ907jHmBdLHElF/xphkmw9WNajLRZMQPR/Pw/byDkigMd
oH4MShJNhQbXNRyRRDw6EgTWHyKAEKRBiCPXCzWrXpH/20aIxWJXz570Y3Tg
JOlz8jB4VjIiWh5OA3QlZ6UvEvQS68AQF40yCzZbJlBYjQAbtWZQDUoeTudf
BhU2G2c+H9xDTkVt7YVIa/uH5IkGQQ126DAIvFByh/idK45HHR0AWCgGFgvi
3jvxj+gGxIlbL8cQo3uO88ZPV3RSW7kPDAERROLYVxKmhKNByFayUQAsbVCc
upYBRF/orR+9zFRLDqKqLSh8uUrh0uoIHEijLacEVBuPyJFZhXjxQ8JVfmhd
IZAw7D35K682XBnPrKbqZfudi0pLN+vj8JGgDED02xW8swfxwAifO3kxxPy4
lCQLIClXWwNIlG0GVtBB7ViHiyqkMySOmvO4GbjkueSd5VkWfcQMaOw0xmfm
4So+LYV/FTfTT1dcHkOoosJED+ks6F5ymSOVwTh2mhXBQcIWDqjHuEgSJSs6
hNIVj6lLYU9vzk8sMMmNcDX1gaOhlH5m8JdOrp9c1BXFkcfDn4zhDxeXRU89
nDk4Idoh1AV3ffiKxulqUPKPuhPONgOnkKr6ze1xZbXCy1GxbUlTnIw5G7t8
8iltpQhGK1QzU7V25TT1ZRP8UDRGYR4RI7Zw3Y5u5D8lV5SUVb5sK2FrHAd9
iIlN0Pv6mRBsDBAxsGEc0+xksEtDtKgHYzxsjELPu8vdvPaZvIB11vBd6V4n
1VqAil7xxkd+iTHHjZeqw5JVCfwbz0BPT/+d0XdzmBMLwj7ByYQ6zGiEd+N0
W0QSAnCdqSHqy7NiCsvawf72d/rguZ4QsidQSXjJwRgN5MTG7FA+Ll/zsmpd
sbTclbm4ww14KmtTPZMhrGcA3fgVLfRid6aLQc9Rxe06T3+LEEaK29vIYRuN
fRNPEc0eTgrk/QFvj/1xoE72j/P6wiSDTe0qV4HuYkA/VPYWF/C5YodK108r
TmakD4ATWjQ5B/T6YlU1uVwhSZE1S04nGE1zRGT5o6bKzdX1keOozrpthVTX
30OO6uR2+NYPzP9HYkvKDf9ZT4Cms7QkSxAPFOKYuBpw66MBE6LkRdX71BYv
/0ffLrNE8hhnVFzVAEwy/1cYEUNIRacW0gMtah6cGKMIeJilNzAc9rIHoFad
jr0VRLOxbLkKYgkSxmSB3k8/vclX++ZV4cmMh87IIf+n/ktZXmELUo7iHTgl
4Vfm99GWZ6xWJwpbpBM7/3vuQOaGnuk8zhoR/F4lhSRXFaUsCdbDngyZoRBE
czteCuas791WbygHhFOeJso+lcqi6680AqVY36FpyVIPWenWnF2AYhMsB3bF
zeNBilm95iCWzn5EMJlSTP934d0mU+bKrrckyzh9igmFu/EMsdyp6fR7TTCt
agBv0P+uIIv/RHhZSH8ccIY+61+AdKy565Y9LTmZRACl6I8xNVyxxlm4xOgq
aMy7Lsbctv29XlHIRV8Ey3e+OguHZaT/89OgHDDZypzZLm9BFRUXZpXtt5Ie
udlmmztFoFzHWznaFI8hEYITftrLRhHwA2r7ZX03u4DSNe9+PZBHJt0w9gGB
6FaTUkHj+wQ381UpDHdmR9vG/bZN2XASBqUOIYnRrjjdh1Nwlncjk1Q2s8Q4
HQAvAMNTAKpPDF4f44WehDS2cjfS6dqQWX8RRDCqzQ40wbrzOuCJL/pfux0H
p8/QOCg61AxDxVc3EgIutpuQuSUPyddhAuKrJinsHgcNUKUz8FrmHOgL4gZB
V9Kc/6VsAxH70FagxgOhmNVvacnVifkK1TisqPNANw3/N3V8po9cUL7d2cva
gdCWFUb/4q361SVzMvYNzFBZM0V5Q1Vt8gwu8AxAGHn9DvqGRG5GjjeqeJET
nBpLx9jVWE3YXt1bOM11z2UqkBnGg16zuruzZjbCP4o2W2+TqS+GzVPETXLk
ixIfWJ1cLPfMpJFUNcOripIYWDrU8b8Jv7f2JPnsYOwiKlNYjvn0oSxc5hVo
vT4MHnzxAK0UBkCfxZcC/yJnbN9gX5+dygzsTJfZVghgYb6laFUvBxar1CuK
SwoHuDv+rI5xwTtKZI9H3fSgG2SDE1xuFQ0MhXmr6YsfEJPjocqG6/+HAFfz
LcSv1K0u1n+2L5ymomebmtLq+frsS/b52qvIkjHcKStIFRUJf7lU/alf+6xH
P45XZZBEhSzJWT4Ol9oAbrmLbAmPh02Y0WqArqJ6JzWyi1Mawnx6KBi4VC2u
dO+DRm/jX3nGXe9Ha6RdCphvbgYxZ2RZ7RhAPDUtwtMRyx91ibTLp8KGZszn
89GlPtum6nDxckMzp4G1DFTodSpVdnfIvumB+vDyf/R/55nllvH+BgM9AhrA
qy/4Y7g0+WEzuAngexVmWeMFf45QHgXx+bCHiClB2ke/CtBRQ/Dbfk3fVslu
/btowR8Ef/JT34lJ7bxjUbxegb5WdX1ctBSIwM9Q3vzxgnquOO9cTib4wWSQ
e0vPHAOqmIC61p7euT1V12me1vkCwSxB9lOGN95HezrM232/0g3pk22VJUiO
OJXmTWmMkWGePuxm89C7JM7F1ZYHsSLqK9RDOOV/hxF24PDCpAS2vDO+QuK+
CNO9gP+MDcIBLiVGy0rLcVhhoBAZzV+g7XHax/u/ckkbbIApxSh+MsWqXeKQ
1C0BVYF5cVurRtwk6RSmhlvOJBfFxHc4Ir49E9HLezToSlsHCaOayjxTgMTf
Awdp+SVoSC0ZFRP2AA4zMwGUKwCG62Du0C3uDA0YWJPN+fS0SDSNOMs8IJKZ
oODvSKP1pxQPs0v5Bzz3YsjzIhKf4V3QIzWx/l7MseQ/+k+IuGKxW7kcASiu
J83nA3Xc5jSQXCn+nVbFrmMFWPWDmjzYXmR8Ikz3SnMedUwQAVuxqq/3ksvx
mBbJkG641I8lOYCbZC/xtFiGsc9qSGVh9JhQCbOghKc/wrVXgQ73O6972s05
PBb7ldS/29wYfAw7V8H5f+4DqSowtb5zBxiQsARAlmzi/Y522Cz2w/1Lakwl
wiIhkL3wYeAwIFp0/yj1fdZetJ8j9752wnccQMwJLm/JZuDJIuJWU/bNJepM
yOUqrEhllySI/jPQ6lcNhWcpxr6F7c8kznMmfWZvqCHOuBVaNTTkmnXPtb2e
qCtpIB6IQYvf8BUPNI39fVyIXqfg7J83KDhVWgeIbQXGO17aOBZhQnla8stx
M8UlgaGc7Bym4dAf1HLzIjG6rhXM7VUGfTepBA962KPe4Wxx8/hX3PVa2j4k
5cFAW4WYILvPCprrTjm5mVRuKCImms8PZDXkdS3kCZ9tbHFXDbKpFaIWTKsD
fGPSrKTyAYgz3RyyDCSZxZ1ythsiVYkuLuUtw8FdwfAKJS18G5J4cI/a/6t9
+Aaa3zzqnXNOuSE+VuSJYeYhrXoHDvGbS+JMHQ4XXJl6ZFOsLmJJzLRzMjef
OoKDkqwGr01qhXhal0mk8KCxL2GHaOvJ+r1GCNSMc929+JV8HLj1Cl+isyTp
+2Z1syluZYkr3wsLJ/f8tB3aHpc+83tv7I/f+q5l2LXiiyFJ7ifbT85jKZAu
4dKrWQfCFsUMhqoHbezf1s/PfdhQJLA173qJvdlLpnf21mlwNwoK2jwKLPVY
SJBmM2pQeNzuha7zwPyIB/xf5ZXYju0A61YWc67dG//iL0qBfIifYFVmfeo+
eGOA95xW94WKyYEUY7uQ+L89+09wn/WjeymbAZzjh5I70IflpFKC0w9DWJ1R
hIoikGDnnDRADLjkzsjAnhlPeHkwygcoyQpDmx5ii0vkcSqYW7WgTy1/gSZm
A2kVFhoNcdVueNU7NFUYR3X/OZn2MXPlKzAMitzmJVvf8RCBSjHWobc79y+L
tx5c0iyyzZIhZ3sTJ7ST0mpuy6FXzM7pBZE9XmHi0TfzERxTP+3lufVzk8IC
IxLqERB1q9r+jiOhBC3ap8xkcQiEiHcYQDkQJj3e+Lc63zgQzi71x6f0u2kC
4q9Vi/zGs8+2HSEZU/uxfXxSMDnyRn5DiHdpj767embhcUj1KFim0UZZkd5U
XEP5dw9sdy6wOmqasA98DYGVdf7X18OczukTM3id3R2jYjE3EXPqBVDTFfre
84JIUsuFHqzTP6ARu30FxRoxOp2dFIWldHpPH+ncAcBTVPNbpWY5LoEBQheq
AaPNvjMYiuVPNECj9xlilO414tBJWPTL4J/ENOVW+IkzeQ6atZAw3u3TryDC
FStZMygNsap5s4V/lfsnqs5zn6pC47DKD40eH4/p4x9hAy093WlL2nx+Okfr
nEsxyGb8l6Oz110S+GbIRmfPzEN+tc0CtgWmwEUZUEeQ9E9AR76PwaAB3Pew
LAnhr+482nRZ+dxG3ZQer0fN7mL3f0UDE92v3pYb6rWBdb9La1v+eqkn75Jw
VS+WC+CPsF5TfdS5cDNrh/AiTDU0nkHVBVjIGlIPZQxD0ZoxmSY/M8ElhGNc
r57Sz4l2jzUACXvTUoLr7DeeCX02TLvKlhVB10TbMlobNK/IvMqN7lKCC/0q
eBISD7tC6APBcTPFLCz/vCS2TOZHci+Olcc4tlihN2zMmabxG3PAftNKf/6Q
zmaQh7UBB8Kbay+08hnSDbk1ifDvjxX35FEwf46OSFYvQBdiWUci4T/Th9HX
ICzhShnxodq443rrFTrBE7p5CrHl8gySdjy2kxPp1Zvvcm1ETYWkDm09Qto/
43ZZ2ZrucU9drJIb3pvMiM5q05RjWePqgpGJhLHtNkfxhiap5nm0lUX91HzC
fH3pllXpRW5LevhbXEFaiFUPTH5vSZ/TU0Hivbuw5oWlw/L4QkEvvq6uCYHu
u3j6wQplYQqGDowJbQN7M5zA3vG/GXxlkH3uNaxE75qnr0aWULZZxMEkgw36
Xs362BpjGAuNAkDrAOzKEGwaXWPuYg3fBWstNEsW9wkPBmAufgKfCMWwX408
y8mLNB8z7NdmJxeZa3eTVyqZQ36fbDq/mRcMDz446VIFnoLDvnwOB68kV+Jv
aFcQv+GeES6ZxMMgyjVeVXAaZO0bqAnfTA9bWCETQsqeTiOUrCwKFBC98Jl+
P48bBOUavIcprxj28sWyDo7Dk6vdHpnzw+Fe3MRRfCUEDJyGnu3BG9ZhG+AS
GVosciUDxxbXaOgYXgTFeftj+JN5E2kgi7GRyzHRGX2Gpclh2hXXpbW3sFLb
QYRFyseuw6noJl0zwtVoMSX/m0sZK/wN2fCWd8OIhyls34EWBOjfhDnXGbYA
cKeEd+Obd+N8aiAEWU7bSihqyf+3Tdidg6mf//+26bonodT2NvWn0v21HXYT
a+hsdqgIr9luqT8fM0Q94DZIwECPRMHKQ3bVbycsxfzfn1qo2GYDWNlKAvkx
To30mg4TSa2AU0toLkfP2ahxCWMSVA/fzlYKYDuNJ9om/WunPmyK2hUxctx1
XZ3X4xFgbZ6yzjGAyK21nYaeosYOKZUQyV7s4/EycZ3+5YViOkep4FNBsMoN
F0j2wE4eQ9Qsykdv80uAXVk1Une96z36Bl97HUmXms7Rz33yvVyBoIlxNTy/
QWcQRcQgVz9cwquIbh+vqItDCu+YlceNjsPJjoFVVdlkvqg4c8zSttCCS17U
61qc9+IuJ231YyBXH14SRn//Mk6hSYbfgzc0ADl90pFNKuDAUU/SwQ9x1DMx
9pj6maN3AWnuVYh101yKQzDB1yx1IY+SaZ67ui7p+ra5pTCLYfHZCWnWYBzW
LpQbpsJrDiy+orPFW7i/LU5bTyJbehmGaygGirVx0J78S+ZZtSg8b0JqV7aB
ttyckagxo0ehHQZVPAJ4jQX03ByzmxjovnmOse//Q2W1jFrA4QKoT80OGm10
607IupfAyZt1tVU5I/HOMwWIKE65UKMnrF1KZ1wm4TxzReOhJwC0vqGO793k
aOS1hP+uQ6hlvluzsDC/BqsThAfu21q93opMKRg77hia9nu/s1SlW4hrViOq
c/IXr5iDXwQY0Jca3pM7k30Yn7TZJ5ThYweQlvnVlH1OociGfP/mqs31Recs
dw7xANAbezR41h1MTUgOT9g7TR2B9q50YD+Un61Dd/kX7YsmapwHtptAmx6e
l2pyZEMIgnAo81ddgnptZir2dKmMUGrxGu00nQvT3H7EXGEJF4qHoEdAyaXK
CQ04nb7On8SU/yVPtOS1gCvNDdtgHPgE+PaQTXyex+fWyrjJJFeZKafJhpA7
ZseHM2R0R/an95PRku1Q1bavjECiCn5TS4U9Lapm9qVyhGG8gDCGHZ9Ajcbp
2mcDgVw9HlRCjKxM1NhSdoM3wwAoOmjtD1Pu3rM2jhNbRyizXBHXSog8dxi9
zbsinJEVDFhZVST1Ub+L3jUEV/M7R+y00zKm+W9mrWIDPSrQJUsMLLqoIBUV
TcV+MUeMl7IncL6Ptn+Tto8+yN6uJ8ubNbDkE4dHBKT+WmU6OBj28anOg9r9
fgcjhFamlJb9lPApSOQMo2fVhmsL62RUK8O0HBlSqW+HK5oaP16cokfm0AO5
h9M7RrwQ8dxBdviRXk/LXGZ5qt1sn7LLodfo8SvluYGmaNXruxXTUPMhVvFf
w7ASLp3FfJeUy73/Q8i/aySY6LO84kBXr/ZAdFZ7tvJzf1P2fP/8Qmlsb03b
yUTPYBsuMM82UGSMBCn+uwbHmKIJ55yHPq6fxeDixKivKtfPKq9C/EY/sQS5
of60szN516kpGlAuEBDW8JvHRRb5YP2La+bVTzcAuYFbYRT7V5ZrG0XRZZ8c
pEdG0Ts1PhKWdGXQWKYMNOkH/B2l90QFY+WAQwdYHaGBUTWwQZxKCBFQO9CD
lLdYbFqMv0oNyBki7INDxt5LG/X34m20yd4l+6waVpbHROUnGVCjHPNcAPVb
CKwQk0AJE6Ehxd5IQejHZtKEXpOUPplZQEq64A71DRorzSileeV2/hu42Xs0
4tQT14Xiska1znCxxLahNWuRUXd9sk0DWRH+e2UKRFarsfx8szdiqFka90Zu
9dzqVam0Q/IsUfxdk2M7GXFDjQ2ipeXaO6Sp8ezQLJktMEPzwcquCsfAtAg/
FN69nkkYEVnjN4fbP/s3sMHjCkIOF/b54Zf7JiNj8PhswHeJz49gNhQytix6
06gq+3MBQJScXNC02pkR29221kP/9dMZVjiuVTs/C/wR59TTcA9tYyLVsIvZ
4hwvR/rSf8DHgDqERgtXIMxN2LUvP7hqCJE03KGm8mb21DQvaVbHOl8b1TAL
Z9m370AeWzNxOG3xhLpFkQIFrRA15HAHIhwYZm0YWMq+FqfST2zleCS0qBxm
kI6/lzeY7KufncuEQIk3mpOfI34tJlct30XcE6je4AjOCJ4Wn+Ypfh8Qo/5v
XdGKhXosihRJQKpX+Jc9JDZQldTqmzpTTE3Bv6bgcgr8nGKnEk0OxQq/7Wx7
HIlYuxCql4FQTr0+a/hmokTyRe9R+V/p7cX+rNUW3+1o4UCIS9m+HdrAXaMZ
6yo9DMUOE1fxb+YHJlD5EPwWixAYSXhvji6bwgZRqhIdE5zWrgh+y3SlpTE/
M7D5Ku03ojzHwaml63lJZl/VsIT4jidHxFKGDk6N/W8VYO77E29AbQcHQtML
ewTPE6m5oopyRqOh00p47svrI7K7XD1dcpUKuyPgmyLaKz8py8d0FG6LhNiH
2fLn5Y49LcLTF/Yjkz2bp0+D4qNN4TFOG+TypSxRYCtvUNuxE2EW3qX8D9hl
YO+/xULc4sZD9fkqvDQpTeXlVU9PNZUGumGEqUpTkADDZ8cqAv4avhXUaIWP
RT+zYaAJbOirdIu+FfYOnUR/fovJIVL+XZOlEPpFlSd3vHm4QxM4VVNdM6NU
9c3CkEbbjvmkTSDhAwx0Jvz7EaYb+Y89ThJv8KqmN0aJI4+KD0/abRDiVh3W
UFFJYKHWkelOpGW3WvoaGD/s/I/G1BinvPnVfnfCGM2bSLya3h7LabdHH3kG
BO0e0iRFrefMPkL98bwXzqOGDFL/Xx0YKMvjcRFSFbTA/2k3S+yZMVFzPDmU
Z6CVYh5WjD32PDJK6xmNHpTY5dYHEq6jhtVFd9D3db/PcpbiiONJ/AvYPEG6
u08em4JGBroKBzRu+86dezjBpbJQ1E20tk/i21HMB7Q5aAPqpj9CRuy8nuA5
Hx9F1OM5Ky3ieUVKwnKKCxGPuNQ80BdYObXY0FlkKRTWLgKdABR2c1jMfZbp
WL7M3IGvh2GYAhBnvF2dFeGEHiRwCVflIw/c0ibdFRgBUhMWDiiVImMV87GX
E2hiiPt+ZBTLyYxsNX+JpBbj5LnlQ63Dg4IObXpKeDNAc+/L/XwA+yxNa9f2
J3ZbTKcHDeezbDx54EOzl8ZTM9aCBF7XoeEWCTEkVvrjnkZrVvsutERa/rrm
RW/WG4fNT9K4fZ8CfAfMaDlBcEWpyyVSQx6NtcvHNFQtXSqUtiimNFJsBaEW
WoByCtDL597vB6t9hhCL9mI5mN9y42Qz1qwXGRkFvQq/gjiXcnBCEvCiKPkq
ERbs9hZ3QfyYneRcufFDI+tnLs9gK9aPbdAgSVtjPa1fwINg23zUtJkVcw31
DpBdxgrs96Qujh3YdciZwT/BGIgsoFItFqayCP5/oCw7OyqKuIZ1QskhmaIg
kPSp1xKMbxnHhMp3JZEqnvXh/6kfe1J1rlPITYzJJsjLaWQK52l4W90hzdcO
IdPMfOnapmH6reVCe8vdmmPCVaFFnHTW1Qsuxrn5fADA2iCStibR3baTTmUk
EKCqVNBg3ShFENJktEZiwao5n67OvewGB0MWYFlTcVlp1iokXILaU4sWt7p/
wGnU9KJqyb4dmLjOzsNrNKK20U42wQPg9OGDYVgb4zXQCsGEzPjnnS/9dOdJ
nMoPoyX7vEmb88P7GoZR1tAYEKqCZsqrESrkIaYs36qsFkZc4xXwRl98uizY
BMK8X/9Lh/QO/wa/rkvvJlFonAmyVPg5bPVKywlGS1SqgN50R8j+J1vq2Cfm
Vxz52Lt2uK0+xIa2l4vpqfPSnmV49vuY1pzNN79tJUdWKL3bkZGJCqkZN03U
KKGhSZLMIRnJYiZZSzbUqteimHjcBhYX/EULU+EafEs6N6eBOM8mzmFIoWh6
O0FCcyRrOn8ozcXn7teRMsH+PxUCbqsQhuEdzicMRIFvuOw6prad0+SreUH3
O1d7IZG5KR1GyU9Nfj8N9SdOZJtpbDBmQGr/NcGPgCJ2ma0WRRhdi6IKCgFy
Kx388ugyn5MjpB+JVS8TZouZ5SUYvY2TC/9VO71iQjwYc4e5aP20RmPUZT1I
fJrO0MiaJ9VlaJWiY+kwt7whmowODJCXbKU1AkNAcpb2Oc4WoLX/i5ZjsnvH
y3CgF1VnA4cXxXa7MNb1E27eSS8DYY3EkcsqeBSmyPTlkW7GXAYbGOZoYToD
9HBXLnurJ/8k5LAl5dawHhkUL9e/7rOW4More7agf+tUdO6EG7F/oXC2wYw6
puHjQoDqXfAbXRyVAouzrqzXCpFoFt7a+ELyUU+j8R8VU/4sMp9Bj3pQwYbl
dKRQ3nNkdfsIDdyrvK3BVHJzpv3z0Tf1MIcXDGqWp6JPzrZh2HQhS1wlSs9x
POb2hsjVc0eN/s8ywfAH7+exxdl9DMJUBKrn7jtABgtFnVbfISFAxUqJLCyg
Ekm/X0uXuPdZY7bGoLhlfbG1LriHDrv5el/oMHXSpeQa4XSUzdlyLoi/rbBe
2hyNuHdMeBAD4QCZm4tk6VRStBlRldoWM08ck0aiI3yDYIcbkmQeGbc/s+wR
6mPFrocVV8RVHfWLmLqjr5QFcjmi0K/FgTyv5nLznrIaX84jzdUNPDh5Cnld
rb0ySvQjr55KG5AxMnZUAvDq/KV4LOuV4yo+mj1e+x80XQwCrZlCgyIiN3XF
lO9rU5bQ8jsaKwiURffS5tMqYRZaXHPrAE3DCcumAFVi3JwxDlBo6BntgMYP
5Gxi7whFuCjNnaNFOUCU7PBQY+/kp2MQq95JmqGwYgZ01TNoSjJN8amW7odP
Amqyj9nIaNv7gCF0QvJUUc0hSUwuFR3BmTQY0H0O/QxCOqkAyRB+o1lpdCo0
+t762S1Rb7DJ45BX0j2WZHbMzYKP+X/RnVexptbKGrQ6Syc83X+j4LKpxklz
rjixzb5TXckk4uHqAQX53iudPe++nIkbcQj5zLCbrH6Vyf308uwxXZMLX5wI
pa5WNqvDQeZoxPcxRf+BNIDOOQBj4Kj+Nq/RI+N52smLR918j1iavHgErYEf
4QPY5dRkYx+iSfF/U9y00svy7Ilf2uBr7iB7Jce5ludtIFk/74MtW5Gc7urQ
9CpII12ppzV65Q2H5q2l2FNnrlesuDpBEqIEuMSei9BOVycwsZJA4sC1hr6i
vz74MKPwQeyuZEq4SQ94Ki67Yb/pJtZYXh61kc3doEzysVbviVG7xo7UEkgf
rnaUcskPPCwTSdI0r1j9ciRsBbvXmTQetkZhjrpR4TCL1iOOKez22yTpe8gp
HaIkenI3LbxxEIrckR4VHLHp8nI0w4+393nqfvK+oExCSigffvHcJkJiWmS2
N404DEpMch2Rb9J5y0WaDCylhHqT8y2PQz+MEcO3gMttXMb8lViQ6yT0sXcB
qxbJYnZH8tFwy8zPkeN4m90Qkk71OrRWwIkM6+/DAxwwvree8Qn5GRrFsK9W
Gi12csDsqJp0B3suczwnCLS5i0aGDCgCARAAPF3SFdr/bZlOkt8kL4plE5T3
n5TAIjIALWAnu1yZW5Nr+p9kfm1d40KkX7niGu3JQ64F1dIfOtIbnmgcPaHQ
35RmbtffOv0ahJUxAklzt8MMR5cuBvqRGgk2QToHYQFlKWz9dHHaLkKni85E
l1pb+L65IN8pd5phX8NQmQriARO7deB3TmbU1tsirx7N13jOzDTGHfB/k5pq
XD5loESwT2y4y3Rek+T3MW1TKnHADORxuViRfQ/7GBEnldP3NZ4Akch4zYRo
wFHSctqcgTNwDdjRTlzeNuVRgSd12HJ4CI0NjTfO+xvQYnsytzdeYPTK4s0w
8yd1wxFki2xvB8yxKgsSnAX+0JupV0xkLP2CnETN3eFNm1eyCaN299AOJyFj
TD/1RwKCueYZnfxCUOyQZkdOhs75sEb+ABxRJvSCipgihGPZT0Te3RHiBd+A
9JL/woPFroixc2HJuzuf1pQEemikt8rTuNI/ctgsQ3Gexhqw+dYavHTP14dm
FcXH5HswU43pORe8lLOztHvRO8CbZo+ne08ln8gUGC4ljIOgjytVc8GxmWBS
xUaIRqsN+3toQJxafuVLoW58kDcZCRvWaxpPGKSjNSCgCzV9g75SYocVB72N
0oJ/YGNjyB5jqtKjfAkax5Ipz83mMrUkN0EG0uUOsTxUkOO1TIh0rrzI/cdf
0tQSguPVJn+ZnXwtII+aPdpY4NKJlmQOzW208obML4qEDd1NCFflOdomsYZY
moadfVhW5mf1bwYnP3Pc+ogL6oJ3GXLkwinzx6YNKmyR/5aVZ3/3I91ELN0f
Kp8WW20sF0KMXFBMbu1UKnFxtva/niWNX4h2g4Hk/CUg2DSl4zkJLt7ywg4/
fRmfPgwjSy3U2eL/pw00NzD+dVzFUoceJTmgzOHWuJ4oV2auPleajl45jPUI
cJEcq+x8xP24Izlq6YvGzcdTDrF3+ga0zRO3NLIEbUdwdit+NRZhVcJJT3DJ
y8xHN6zfE63et8KbzxA4P7n4iWw1R5NpveqbnQ1dXHwaMmUDG0AVFaKURRwc
9kuXu8sYXxnI6CyI0DXxwuyliQD4aKQseUaNvsRp2ijLmm4MTUnhXv4kbgnn
m+7rZhwdoVbgyMPXyjJC08G3I7nj3+MyXHlXwFzoRM1SmELd7c/PnIGXkIeO
6NOj5I5D2i5T0iGhJUK9VxX/rBKct9dg72Yxsy+t4P89xdbE5Y9wExBvcfJN
14VqocpZjIMI3mECTtOpdb8QTfGqW2mRHTrzPHClt9dgfFj9xAcLSxYzHICo
6Iv8xWiMEKmDGIrL/lRvFqKB4+kJHPDqo4kaIPbCwP5rIrRK3KU2KRLSG7S0
vD/a6IGKVvOsidlPRJBNNkXIuQhfPmmDJoifqPS4NYFo1DcrxaYkx7E2nP1/
K3N2yKq61SHfey/3QBMhUU5WsMV3DDGadlmECO2cVD2mfPTFYlyHQJhUhOlv
QEpyvxK1x5/HQjqX7xMRjdb0jOz4XfdwGvi5fclr8WzMfV6siHnOLIqgdRwc
pUnAs7reBkRAWBZPQ/1ZXhg8WlFcYQfc1cC4QlXjPWmjiS3o57OFcUGzkGKR
ValpKAc6K5W+pwv1wfaXdhqRloDBmjPr44sIvPjz4BhkyUEXwTXv3BaifHBI
7Br3MzwUMdqWRq7ZD40EXhFsJywos94uCLtyz59mq6ky5/+IY/EbDshRtMvn
F3qoDodTRzFrJtuU1ROt8ttiJy8ZUCPLvCsFvmWDDxyDfG0Wsb0a9xcTawoO
Mc8JbVKc1hbxXwM6cd7r5CpvB/wELjK2bWGmUAq1BYq3Up229+3XJsW5+76C
yznf1EpD7txIPDsvRJqCWEn59gAsl0duN2wEBQjnM0IEkqptb8LoCHSvyPhJ
7B6f6pvUvzmf8fjE/qEIE8wqnbgOx9Cdh6MEJC7HG33MBIbrqdpKZ3S+jNo3
/6Ww7f+MkGDuaCggVcX7Pwcxq1K2kozSopduDqrN+a0pQKXh1L/SReU/0ZJ2
K0HEgHWy2CGu1srilUj6S/HSfHOQwj1HRHSnUiLTFE2at8BoxYl5ddAijY4D
JAnDTH1Mt670awW+G5fabHWErI6kSYKPLTbMD+PAp7Nte+i3ikdrWHLSuVEE
xJ1Yv7nT1GahxWcHxjXtFoal/eu6fPjy0AlnjaU3sRgMfE2mzvEJPwUO4art
5v045Jtp+QD5NJtLyM5us6Sa5KjABf/eTEAsMxLuPmB/romqP7Zb/5QdU3Q3
TMbF2hKyBGWNI/ci6xrpCRIfwMdErOTaeqf4YTZRtEyb5Y6eiNbQnRspcDn9
tzvmvg/RkLDEr4Qly+5aIzxI4QkS83HEBSg1YSTYwzuhQg09r+FacUgZxjCV
LEfT+PeEBnQHinYzYYeaKrTLFtGV3u4/5uum4lJqwZrL4CvPbR7n3+CzfZi5
qmTR3PHjpIglEQ4js3Nk/9Qf4UFySoBfO9Y8Y92kqK65IzS9D5oVus4h1a54
LFOofvb3+QNfBPbs1MktKYFPHrqrboogqJYIRHvUh7jDYWICVK6PYwag/5by
XRv5kZm2H3zeDBhFEjbGIh2Z/PFD41lhvgM2/oJ++AZQ/7XeardYzph3PRnQ
Zy4046P8haQLD609vs6a2y+XVOCCWwWVaN6A27vJoLZ75ZLHYm7SUdrrn4jG
2xIxpbYj45n0Z5/NLVVneZbWlXqxrf8suQKjadgN6aFiJUQ+S77fLqSh60CZ
QtAsIUTuWTKGyI5kjF4kudaNkXviZ5Z810ra1yaoMpJQSyml7xiqeNMwLJzg
8ejJHXObCZpfyzEJkg5klQJu2NhlpBzAaOphlR8NjK//yuMAS8CaXYQ7D30c
syq0ZCu7ywFiwh2UkcKRaXWTI1VkyWT5veRzqKi13N7uDS1SNTAMfJxiAL5r
toL0hjDINhCRerim8hZFOj+1NOmpyZ43c4UO/qFB10FNnANXrZfGMFiZF5ef
btq5b9mllHA3lh6E5jxsP+teAbHJpWKyiaPk+sqa0pbDU8arEpqBt+rwWYLl
j5yTjV2Ik5Uqk+vWfNk6sXONjnHl3OTYcESEojxTopsoYo7itCUdMohWJ73P
92mwlsZlwSxO+Bu49ssoecL2HJOhCBdGiC+3uYdmp73VyxIOFlLWMiQlJnuQ
Q0lkEfH03MudDxHooew9JFUXJokh3PCMvbT5N6BfuaSUxfRG8837gUPazpVf
+rGi1op4K0IZUWJ9idWMIFJEsdY9je+s0Cq37ZGgTWJHu340XunqMiXdXFyU
J4h413Eca+DuIH3X4+vXFEMV7hsp9HyTDKx7SBuVVkax8yepEqI6mSFby0gF
aXuvXLIVvyBPmYDBG93T3Rb+0s8NAJU/o9qDlefrs5b8hcGrRcD1yBCjuUPq
BISV485/H2vqv5edouBP5ANg35SsMZT3WrgTc8HKPq9EP8Ih6c/laBPaYoy3
/BKEb4YUwGTjB+CP5Eu3uZBwKjIPkW19oRcLRtudwiTltx1WX8cOWywYgn+/
/d3qpNvI3CDSDGiAFpXvuKsCI+LWCbGHFOEWS9SR8bAvF1BNXu5io30wsn8Z
AOCm3dnFo/E5fd+NaRXdQcMnPb+kX8lfv6+atzc2A72AzTIbJX5UMYIrNly2
FCQwtrs3Yi5PI13W0DvW67YCjfvylqu6Tcr3B0jWQMIcl5wXUSugYig2UcaK
STiuwwcDFLXH7TzwHkTNU3r5yGxiqXboPWfJNs+0m323U2PoiKzD76M0UJO7
i/fDRjTVyvbZRZoK87hKu0eRrTXPxPRhdzYfnx0ah2y768G0xk0u2K2rgRB5
PZCyym/lbljeCux0qjd4JS1CDz31u5wona2/noskw8OHqBQLJoCAFjCFVzRK
IulvF48ju83PTHDUz84CkLGeaBcjtwiUirvx0bzY/g76g20T1DWRXcSU3zAB
5V0lM1fVsrSm2ugelXSDoQtmAWI0n1eLDdITAxzqGt3U5gJH0Dyp7EjC6IrN
28PdkO+2X+EnSd8KxrEDNKgnTYTvSKLezXV0f9R5Tg/rn3GYC5uoTl5anUVy
bv//mHr2PHxw4YhIETtxpq1L3p0RQ+fPywlgYSasXxeBMhEeWbC6twQYf+2i
5njqyq2iR95CDuhQYXrWdStC+MFTWp9+h5iXi+Pj8OI4S0AGVFkzDgk5Es0H
5qlLYu2n4E5BkTq8d9sKEnrs+htKvhyFFzs7dLbzByXbr73MJ92YHruuayrT
OQt/KxHuW8dFSXUWNd75H7UNyVvyLPesBJOEu6ZKvDUMncs5ujsVjEPOaN+Y
9C1J7lEElaiQUyil/Xu9wbkRLlScTlLQNS6chCEW/0swZw/w/KZnoQZ2ukqE
IzFTJa50k2+QxSrJ9ajGoPEaR3trjNxrQKZ81RB5aD+lsWHuPy2TyVxc5AR7
9A09WiYQt+lb53LRE0GuamEBir2bXu/HZ7iCIF0DX7Z0ZxTbB7tQKq+2xRRS
qGf3BgN5e8Qk/UZjqvY60dmpMfe5sr5/YGCL1yZ+sRTcifIiLPc5WlLYSudn
hwfR0oJ/7KIfF6CKW5mhiQuXHEniAzkf5uL6OjJ+UvK/OYjNcdjn0GLtn+EP
yC2rQXYhRvDd/K8o6S+TRbDoIkwk8kgxRnkVle7hEH1hqmqFvwJct0G8IpT4
M/23iK7xcFqbg4TiiQ33FOLxuE3dKmXwJp+c7p7TsHhywoGRCcnX+ZiBy030
s3Vn7SfMKZSLMAxpXxThydkdwJ0ps1wQln3z6NpqIPb43k28Hnt2hcrWb0l0
Y5vsQLrktZHpRbnDvfFBftQIhxBVk3uJrgM8H+X6Olni+OJBv3LPbA2F8PtJ
GnhR1zaospVFP9Mc2Kqk6HClfzuuwvJXOcBX1o5yD23V7R1j/glMagrRitBb
ZA5uk5LEEjWrRCcsQNgfPJkDRMSBSC/gEKWlsTWec3m6CiooYdIAJcyXWsDT
U35D19XmzxGV83SL+hnan2Qmmw7pmkqN2rFiw3MT4zOFnDLJuoD3CAalj3z8
Y/1kpgVI5NYXC5eIYyAy47TyC1lsTzkfEky/ZQxuqhP2fY+HY2zHu/V5Nik/
fx13Sg3n7AeJc06NL43sYF6wCqK6R9BBttc/8IHv8GVMWcedvWDlhbfll3RC
MN4EshoxamEmlfrYrRf1T8yT/kGu1ZKdZHd8J9YW/81xLkFV2FDLj/xTSiod
SfetGMp/MVq3v7yglb5WyiI9m8D6nR2t1g3ZhJVvlExfmaQWDljeRpprW422
9x2M+g5T/dEWJPlda0xOD5+DvRC5FBHUnpmPLDXpt3uy6CHJuiGHp+DX3OIq
G5brfIQIJ2X8fuNBrXwu+FfZsfG/sXCbf34BLAMflMiKc/sGd0zuSPP2E+Wl
lhqrxX5JNgCOXq6//O7xD6hwWCjKEetTisPxxbNOTk9RaPdHydH8EJA9a1XV
p0V1rVN5x+/dXNap06J5fC0WPnwAkc2S213anhJqBSVC05XMFmDW1KWaFIfv
cK7vQoeDs6jiKqdVjzy26ZN2ohmoFofMoI/sUYlyk3nguYjydQWufotfdS8K
T5VpuNPMbfjgnzcVyZMyjAaOVj5aBrpHdAl2S42D9k7lYqoj/vI+9ZHSqm0/
cWHIoUAsteKVRi2XiTbzI1ROrU96i/Hv8Dmjg5dgyxrla6LBblRKL3EC5lNd
qfNoMF2JoEbsTTbyfELkIf3bbUenA9bCn1oZ6T/gIptaYgrxtd3UOgcjRWUY
EuW1yKbVV1eE1rqe4uwLrTpYLfmGPBBwY/6LAOpMlUGtSCMf7AiF4VdRp9KN
j/1r8Q2b5Xge9BN/pGWkAYONsCfx+xTImc4fthSCDKNt3z3Dgk1M1B5weEfU
VUHpfVV8kwS9Bc3F7O63oyXII52Vzcxk06jFSUyeC3urcwhvmuRzRrgHptgh
Jl8G6p+j/RnCOkddmznPfQFCsFQRJEU1TXuQ/kb5nsBIJzp290o65yiwN/iN
KkBNArCEaGsJ4Gl2ucnn8u/YDMduKitYPizxILEEqI4skLPl1jXiWzeNheRm
7kvuDmmWJHiWg9ADqYv/TDmzMlk8HQh4QJ4Q/qQwSPo2qSLlIl/igj6K+Ni5
NYsYy8ZIPqd+OGvdwyM1FgLsuDGJOPRUDNAkogxRn6wH2Iv9fw4oCQKW2cLA
H3X8qmCd4JZvBI2DS96DJ3JKrXvh/bGfkC7thTKy5bXDUWmtlR3xqssk51YV
RFteqAcVSnzxveZH+kzzq0z/YPbV2UeFAYA7K770bsiIp3gF4lAWGhoHIlLx
yUmp+j9Tbst2mBnjgsiOKKv9KrbP5V7JKsQn8Od8I003rWQ2WGHjIjnsEE95
DDicNpQRaKIYDZo7aqpcYq7YmyNIHn6I7wYK2HnDClHqkR93R5ZFujvwrb4S
tC8Tc1N3Wvmf2Alrhjgwtj7SETXUpBTdLoxPCPKdDwkAjhIPWLFqpZ310AZ1
vdcTe98m4uE+nr4g8CTzY2rRThIjCw1EFG2h6mLjKbdgidRvEzJolAOvpU53
8l5YT4NLvJDWpe7+Y2ZgF91Xdh6eaneQSc/+rP7unOdhPnoypKG9tXIZwbNF
ppnSVJTH7e0wQxtqIlc87Qdyx2mkTT0zaryCzgenAUASuUM3HlNmOtGCd7s8
ZrsycPaP/M7Wrfb8yTkS+Ee6J0O23FqBsy6BA56KTGnP5KgdqVA3jqTklP48
QDle8dbfINCQJWC9LiqH06cMLlNNi3hGnxrU160CB5LzevfnBkTnALPfX9p4
Ih8Ly4wBmT/lTjhgFMFRGsLRQzXCa7Jg326TKqQ1balSicxD6ZrzAk3/GchO
qvOI9M0YcBe5wnH2sY09I7iL05IYtV6Gp9qwxMryOB/ZWQ+rnpOEhCZKk1OO
Vxzb+L96FqQmRMR0SPFKf4mvOI/WcRD7IZRCNODwyOGSk/488oDq5OhEXyGt
R+pNwNdEWOjOOkhgnJFpW64Dg10iCY7/0E0dkTNpXhZZ8o6wNP0WPaAGm/G3
cr4NDSgkBKExjUyJpcMjpohI1j82/zuGANt6zm0FWpmqsh7bhD6JX/NNGNaZ
Q5Ov6mWj47YhTvb5Rdc//+1cx8/mVaUeQU2pCS3dbfkBtvlDg4ukfRH8Y4WV
XIBN9Ne6KA4ucGMTZztmbmDUQqI1n8vSSkllrHftLkjaOP4GO+53Rl1rYH+Y
+GW4E+7H4bovy1UV10+kuGKs+nHdgGxxerdF3zY+zLEw68rId9qvF2gCIxc6
m2voML39fZ1xYoJcy3/KWTZPwj5UUOjFK7aIF21hVcfbbEiUClgjKssC+nha
4B1vP5BC8FOCqU3tsU7Duwwtfegm6/KXw6mTBl8GbHH1WSOn6xKjWRYb3np7
lbfjX/5HBGPWwt/BkF9+K4sEMAO592VYzczC6SEOkdhfrTW5B2SDq4yyu59H
eRjqlT+M7HJSw5vVNWPr4dRmyQKVH7eKiqGJiDdhR21yowXTb5MAro+p3ClX
vnIRRKE/d11GZIiDzVsZZ9+r7hI3w3jhSX7MPuuAyFVLP4lqBiW0eIsiMOqo
mAgVqKWLiwPUEUlaEcnuTyTmBPZUDYw44q0MUWLHi6WoUHEebLIecKQJ35si
GWqXH6wJWZlV5P4yU8603SpDgwHJikY0B1dZvk5wtzC32clvB0/muE5zI+PK
4pgvQmgxOQ+WtMb1/1n2MT/8khK2JlQa8QAs2cCeCzX2MJ7qgUDIdaoDD3EW
gGlJZdvfzCZyulAdnX4v7/Cyt68ZXctPbHcwTPBdc+X+0e/S6Qbcon9BktiT
uhudhO5igmw83cTtFWkNsKaYQPb7gTz8mWkus93xW9+PJ4wdEPWWgwGYZ092
wb2PSrPp9cnBjmrpqAZuxs0UAcMHDvyZDcwH+zK5wAh/DLQtumtxim6+FVdy
icenbDHI/PJPUPfaoKu5zw5kCAeJRTCOfFM5YzA6Qxcg5/FX1QmfXS8wBoyR
cWXGpj816qDA99flEN1nuwIy4bsX6K/JhufOPUj7kuYS3vPYivJJ2WX1SShQ
ppnU2achg1nVuDVTB5js4vSeiPU5x/w9mAY4mPfjI7uf2H2yvGgNSbziupF2
ECdF6F9/Y2UtL9nzxud2pgu5OeDEbrYcmMLkrmOmMcJOem1vkND5WU3LWNGY
DAJZpCD0skk0YIg7Jje3jHtv4tg7HdW3cfDAyEfGEXPRFu7XMSl/0IBZWvWi
7dn0b0UriAOU5hxDVxxlTLYWGewpvDmKHaFOaCcNghw2v6+rbtkMAmvDd8XH
WAfWY1n03IuY7J+AFI3l5o4pVAu04owER4iKPrslEdOGxfY8zPuivCHJytDH
httTXVOJ/BHaRH/LNgulQCIeld8LHfzDDj2OrMH6YiC0HSlKYS74PDJVP47u
DYalNk+daKkfffaGGaR16v4z6kBbBIG6F6LxzC5zqx0SsMmjPmy2lwLAvvhJ
7cVAgyisbsH4eUsiDnJ83BP3M7xiybmb8di/ywvyyFHbpsK5gAsKcYEhXh6K
IYyI7CHerBmdQjNtQgZn+8OygIfILVbP9OL+cU0JVfxEdVLl4+I6O4SLuDaG
GAdSSrYB/X2wj+DZEtsb+Au6zjhWHPP7P6g3m/n7CTufkw0+mB5DZXH1Txld
Ms95uWtFNb0d4rqoQy7PPszh3qjCNwHHN6QiCh+QWc1Qv6m+5S2DMgz40A2t
H9y2BXezzaEheoIDVY904IHVqG6d9kA73zyx/Fdbazs75ylOuyJWUBeTYALG
rb5pSYYMis+1GuudmGWSzTYidRR5DugCh2wofCbov2BfpkwGoFbUhwJeDTsX
th6ID4Q7a6xvkmMaeWrUOCa0Ny0EBXPyC6qckldMZ399qLM2TMCkzrTKabtb
yF0pduKityr6HrAOLTRPWvEwEXoUtQj+jt6WfvQsw11RXJ0JO283ss5CiHrd
8TjQMt1DObqwMOO1Clw9E2AlXyTc4hOk5HMAK4JSRTV1MYQfgwxzAZreLFg5
UNGSjAn2mdIyljwVKBBl77vqutcKje8Y55X/dgh5EmwxqQugMCwbO6kKvupv
b0hvT3TIUFRVpV76/CfdZTla3XCkqF97o1C6oTigHvdeRbJ44ScRs0YLqISL
vooeAC2M9k2vo78Soxv0L8dRd6Ce54/9U8Cgmpk82XrBMKgPMxI7IYC5BpeB
FE/8xtbmPH9izIEUG+9e9msg/H3nDGtIOXh7f7g3eWDGuaY8DUpRrex+yK2d
rHA/yUS2Mbrnhs/vPmjweV0F+M0E69rHMV77qbCphjahtKLU5di168r3Rl2E
o0KelroZYGv16/m1cSDRa0FmzDLpUkGQ6diFV/wsbRQzLH4s8mQPNMdh06PI
nkLNN+u1foKpA6WY/OELPQ4QB/SwACq3J1INwl7PY4NBBfZvCDu+fUFt1F2M
2qc3X5MNhbuv66f0e1NiJSPE1JzCH5+l9bing0T9AlRq+YVariOC7FsykjdJ
KaR8wLsBPDrdMyIx3nOQaz4p0qZqLfYVwUXWqJ7gSduU/z5AABEPN/JuAbIW
xTHU+w0FJvI8BNcFfd/0rHsuGe8UKMY/fhVWjwrbBiOJFBpdv2xnlorWytzC
547FN8/Skjl/szQCH/ixV+Us9OUWg23E/Ov8cb7V/3H6v8AWA/kTfJPidx5i
KADE5G7e33HBfHnA2AxCmHSwF4FkVcW24tCHJnlOLSZTKudGn4mPN3qUSfic
LyuLLEzgucG5+dkGkShPRbHeGFpX9lYzP3WdMiTddaZuOypzX0CBCYIYy57V
vHONEELyBVYnqyMdnAHaVd0+U7OF3Am96jBMQRZYXqfa3uI7YRH1e7ek1p7M
2vpdI2+DiAB10ir5MWpvT9jdGE4StB6YuWVvjZRgbRlu9jQRWltL9sXgdqYf
KK+qKilrBcwycCMgkFz8dtai8PMBCkpie3bsRNEC3EpvFZBGVm2T1bss2Jpg
4RcDTFDKiZuLw03TV1MT3uNrrYnuRkytcZRROPRywUrCOMqF/5Xt7KDr49bz
qUt4GAGWXr94JRuycU2sySA6lMetVbOk6B9EvD/CGIfmyxW+N4aDcbtPOEot
bmVb7kYgDNpAjcEPyoaQwWfn7HKHKZpk2UkwQmGsCNiP/bphnY/Id50FQAEE
LZdbleaX2/w37qvUQUIsc7A6YNX/a2Iq+4Kk4WUOGHR8Zru73zjcI7pR1xgJ
JxiMKG6wkjhtkp24bHIyviehQGqmx6X/53D4I2n/91r+/R0XAdPqHIYI+2Si
oAbz5xH6PmCqWc+kftk4cfyPD+wVp23I5sJY5YiQ5PrTJi41pj0Yd0dhq/LH
UsC7BDnd2AkEleiZwgU7x77kAtu7STtLS83BYu6/EdX9SXLNo/3hLoOgq0ud
wgEVDndVh6rfCp1IzyOe+9lCZoNke4r9C2snivGAv3EfA8C/c28Azb47eGXK
mS04t71OUsJoqtmumN/rglcmBBJTmPJdNTi4ms34cp5aRk3bM2vqplclvr0s
391tr2KrsJSoKJ9946SMZxc0H8DKF0LXw6W36NV0j0Rlg1Lzu2kutnFGV8hl
lLY84pkoVFI3yuDD+I3EtApjQD9gT/d4+EorQ1kJmRVpRkYy260ZQYLhGOmS
zZsv+bvLLHaQgN7qLpOTT5/C4LCuotAKNnnpQe2LyUipuBH3q1mYdsDAk4aB
Uk5syJ+sd5QaHpJUb3QzoSo55blnyKvT+jAuAm0y4VhSA6XSz7fWb7Yr00YP
SufmbTszefyWeDNPhW2hZ+Pi87f8ZSaCK+nfx55LxckOLK3lJ//ZCeCUpHJa
9rcPd7KyQHCbDalTGsdaYVPP2RIAgFDy8/Zw6mLvOMWtYf/mrm4XDUmYazYm
FTezcqUyhKyElVElAxf1sgxQltiUng3ZN+1WhX3zDMwLTpb1bByFKQrpUxJq
F2oT6gSotUT1YulamFXcM0MQ0M5oIIpwoVn/tx9QYe/qqbSfp1zDHOrSi0tk
0StWEQsnRvEmywHWefWZ0+ps6ze8Q7mgUWVgEEIMUfYkD6UbE6U9Hmgp1wWm
NWYXas7gqjzGDkfjpGFpyNMoS5RXT7Pz1GDWFfcZJsUi4Rp2oGZuaATaygKP
kluxnAGJ6fjlB/EN1Viu5uv9VCsx+YzKpPc3+rNNWxYRlNjYtIkhRb3hFbsh
AnIaT6QYXsdx3lShQ+SgU6Dr04MUg0D5RChZNxHJtpAiKOcaJyxcfRxYnaFz
VyI9/ysjatRUPJo+wlxjn8l91I6R/CpLV3TnhiHinlRKD27tRLFEWMCer5zi
MJriQXpkOC/epHtoNjPRY828PZbu/eqiFdywGG51iDk4Ktc7O9GZIN2Zd3eN
tyNtcmGF13egBWbTohGF3l3Hqh59yTGSWNHWox+krL31DuwerzupGm4m53fD
MtLqPrAjOx7Y808E3uDH0VTTSSSQ/9F8X15MNDq+DzN90KH9zcNByz8aB7tx
FZnZp1ok7chanKlvzH2RYhOP+VP3ERLBJ/4J5LxJGhA3CqFe0kr60QLE1FFy
nnV/NTwj8V3pkoXREd2PkDCk+nCEMoQrhV77h2HuRyXUyjhxdJ+/kuTbBlth
IfhB4mAS+MDy5oev7frUnlNHCgAoy4eHzETcXe0Vas9PazLBHrx0yHX5eOMk
5z75ME9xdiiihiLEuKZcJAjFscUbvp2vxr/wnbcjiQCTVCsN//H1oFfEiuYn
UhrIiZr75wpfKlduX0Es1fHYHFomBX4wdGj7Npc6+FG0WPeLfBJvE0fEBSJs
lPixwOu0pNEZSPY2PJLWW1VA5D2zcmhGzSV4GqJ0Eg2TxIa5RR8HRuxe+vyS
HV3uyGdLDVRaOOdaL35nEu4HhHtVZgoenvcidU2wdUXduVcwUVofJyDX2gxo
BLlNODKSH9RWx8OlUg+N6gQip5sjXxb+ejNlCNfJwdqESt6t6qzzlAX7R0Lo
3xJ9fwQVv/EtqUG4NKijrc9Yibfe+lkTqG6iDnCYoQ0C6DfXtvWiGsl35a1G
+dHYye/xqqhp5BXTbnIii5OceGs47FAFl809aC18ooFyqoHAIaxaPTERUKDl
20KfNUbAZQRIoc/Gy06cv9d7dXB+1LDFBXT/jOv6Naez7i8gzfLlSLkXytbC
pbUehEeS1keE9hRWq9B2fQ0yT45Uubqpf9o3stwMqrO1dMsRzw+9X4rv1cYf
klE8cOLYxncc4pn9uCDxXp7GUnpFs6CvYMMC0fdv4tJDe/rRV1iKzeG30nk+
ckOmPHZoXSOTCci/QnL0pg6owTHUXAg011fHqjHHQ5Ew+515fGT/teRA0guQ
lrjRoS3T4kxrX3ABOAr628BkvZE24TXizNZsNx4iNilTLiQysZtnOj8fo1h6
7nccXL/Ke5Pj+MRomvpDrSJrYyo/PiaYuml+XNmgyOG/uJWwAhkyuamk88z5
y/eIF3Hrd+Z6Fs20Qcsofh5SHGtkE3LEtcg/aPK8yggy+3lUrK9w9bUFoxlA
SDs0EfSamV3lOmaI4ZwV0pX2+ct20bfEkjTYv1j7aa8IVF10GOPFSWLbZTqP
OCNfNWJHdg8VuI0f/B+Rksj6NOYC+UQzX9IBrKqCfzSSUhyDG0nCaJGKUH8F
O/HUG9QRXs8KtL3XK+tn/uDMnW8+tD/x4zIwCbR47c0uKur31s5i6tzDWDq/
Cc0MmX10ga2ZZKx0mXuRXs6eYHJumuCtTbauZPLO643YHavTZfnsP5vtYZDv
IJycfSixFyIzgg6I/Ia0+cJpbtvqDffS5fsR6IqlBV0hQoT+J/zJzY8ZNNYw
7bHTB8kv3wrl5grUmT/OlAgm64JAAmRbZ6OwnNTx073jShYZ+zy6yGOs57GQ
3JHnww/+hbfDAn6oJfqc2Z46aEFFrUj3vvappstupnMuxN07/6BiiPoORNi1
qI8o5Nk/Xku6db3CnEtF/Yuce3SRPIogsZP2Ewp1hr3uEdTBrnH0q6j5Sy6h
hcHuN/bvVWsQCUFPufmpw33MEnG4mE2NW4zVlLKB3g9EqqpWb638nQN//oFd
b1sLuSEUsrrwpiPAvMxhSuYOVHkC7jOxkvj7+l2TRUTJrnYF+BQi4MhxlTfH
V3M2ulyGGWKmBXdKk0KC1mtcHK2yfQmhESok5K8+j1hEhcInyAC47Jv0hnMv
2m1KOGvFAaxFD5m9fiK7lJmKh0uzoTGWayCVz0x20wB/cai/6aL4c+4lz5H+
s0ysI1QOGdWBY6nHgJq5ECFoto+nEO0OispZvnUeXLHmstZUSgnjL7qbilrQ
pGnKTlwjA9Ygy0tnY9WR+r8deXdLaaxO+/lqaZ4eU0OCmQ/loehGomWAHGvx
lRgrvAqwlFY51PEFzjlZmB3RlAWp0AMfTs3ViBz0rw1grYY9bNGNBsuxEhOS
INS4+lc6ueHTGzUCzVlNRv/Nn+Wi9pGNKEPuV4jUtpLj0G0HnQ6Uv9k+eD/H
5swuhl5ZjqC8rFdSncPYGWmNJWfmbd0hn7Sl3if2i0TCf57X9GJlnI0eYNsm
9gM9delq6NqIuTRM/7xA9aTzfJ5UbTBUU2SOh9Q+Ssv6HDBbCZ1ruwJax1qT
ykoJ7m/9tTXV+VIJ3Cd1r1FBrGiraLJEtOjHZKKT7DCpXEjKKv7x+D2IGmTU
yupuca9JR7C+hNwynKjfk/P7gMllgCY3O/Ds0SsTBt/5LqLDBOirZHWkySlY
e50RNtK5LAmYYAPk4kce4zSmMNwD745DmuOPT/j9uMMWMkC53ppReDQo4J2r
obzjqI7MwDiL1/izRquF/OFi1xFmWL+naeMC9H2sOEXHDOkWiyIJX4lDcEiI
zElQgBEQ2kPO7LtM3oTe5eOpHpBUqi0q1AZ5pU8VkjvhzixHHlzJsoiyRdVb
NnScA9Xwcfa4j1rw0BjFh0wgecF0X3dqMNpsNxQX1+MwMHKbpvwPp5GV4VE1
R2iHGanRWtBWZSh428IyEjDfFmcAzg0BkYiwfx2oRFX98Mz1y77xDgICHaXc
MLGusRR3W8Pv2cUKdPR7pKcIa5WuU9LtTXGIXK2kWcIYIsBpfzSqfTg4rOa7
5Frj3ZryVD2r90GlScL+2IV19w3JJGBgDwWTJgO6d+h62hfM8GIIG0KmAvPg
+hlrZXinItlP8CB488caIxRiCSuULIgIH6MfnisJYqGdnUfUmG4YoLrzfguA
xWSpuArkNvcUZoqMP0JAHPgM+Ah4Jao51KQgyh9K7pBrAFPLJ2WCmwesHH7p
1gnw3xnXBsWAetK0cMxEn+LncMkuqmcFAzfTAOKGKVtEH1CAci61OmseRXwE
r+mrlmRAkn4C0HDgJmzEEz+zgdU1iD941HjBdGuezGMpQG7Ssp1YMvj6wnVW
0C4LL0nutXihLFCujszO/fhdNYNgIA6y9MWiswMX2YQQuDOIzugn+iI+Nx4p
gM51N0Oza/W4NPCQnpSmVAnV7uMryjxJbk7LReCPqlEApAP2cdEHf6x5nC8/
hRIabmpcY0Ztq64LjeHMKZQAQdl5NRrZJOrbuV1S7PxDgRRsnqIQceu9Y52m
AnHOGH6istm7U4rgDvVpm9YdVKxTvXa3UJbOPfVu44XpTokazJ24RkVYB8xV
eehGCOlrY2vi2/m4svJLOvApzkhqjc4cDWMhGzB91mKxIyN4XPy4frE8imuu
TmkMf0mfZhMSoh9t0NncNTkvkwEUp5j1nPPjxPAYDOy5gtCUd4qogTBF5DWg
+y+FAtqLCxKkPg1Hl3TAXorXClqGb1lJ40++0zqbFrOfQANEWcVr4xNRLkbi
BXLWmYzwiCYqnRB3D8KxNQOD1MyVgkYZ7Ri0ntT0wy0hKTo/1UtV8RSBFwpE
V8dS0LbFMI2pT5UUSZfgW0Wq1NCpxDpD+AbSAhCh2b7KsnGft/PmjFDdKgAS
N8ClWwSOp+SoBt+LINZ+tHvq9B5BZuk8MpuzkYeyya4C6KU3xuJJxfqvTmVj
cPSbAH6puwaxd7sk+OFjMpGChpDbrzmztyCnJSWbRc8rorWey22x4mqPKqUo
FMYfPRwQcgWRs66hWshZSeizioGVnssJOLySOtGdPhWfa6/spvFKCi0YDBfQ
tnb7Mn+UxokaExOiaoEgpRnbCdvtKnBy/MoVp2uDs9UHLFD45/PcJkjjI7Yd
KI6y4+yFbuuXfQxGSNaDPJ/RUe6DvOayllWhZpNcg/6/VXnTUzyWSyYgwu4k
rX63Vpc9qgjLDtJYp3HiLiKuMVrC/EJSEuNEndRyJ+iA3DjE1BAmcdCv79q5
bGJZxlbl6TMdmIWg6ghkt8jyk0AJ4cf8lXdNSO3GNa8t69e9SOFf1s1STMT8
nFq84M4tn0KARrjMNGlP00vfaAdxvWPxJ7WQYK67u+iQaxYFfMU58CUnsYPI
JTS5ZaXbZqcIm8d42Ux48sQn1Yscw/EGCJhr4tFOMHudbhjc9STTkCABoFKe
1gEI+q9ZgbP0mLVuM5nh9rGa6t7MSLJer3K2Jq7fPve9MRPeuzV8Upi9Ko7I
fDsoDIASIBx2oXYM8ifpan+mtFJmz13tu5vC4JEHd8qlL21DXETuJhbb93aI
QiMiNOOTKb8dHJAj4kATmwiSSwPZLjOu1Xs2ocwbOnbqlxVgJViy9Xs19h9P
mD6Os16CJElyz4R0kjWnz5VmHBwEih5zw4Y28Judf/9Yyd5BTpX0BB7EKHtc
SEvblChpqbpfyv16UdsJX7FG3wLbwMPRDMZfj+FoQgK5Mo/Pq6YHMOOsCAmo
gMFpBkjd745VzAJ5kBXVaVmYF/gt8Ba/5cTCmq3Zcnp73F3vWingzvICK7sT
03RxY8qQN84U0Qg9WAKHZNhLb6UiTJxF2GSG175cXk8itswqP8C3KqSmtEri
uoQxwfb4M0V2mT73aC14z+Mp64XY9X9BRRnUAz/a1hWQxQ6S2cl7RWU8fDyP
jE888aUg2/8wbRzp/5GR/G9ktQRN4l/f4sJzJvo/OLZ0FKNtk/+hkO0ztvVQ
bIQ91J5GeiigWDbUDSlbNlY1kLtYn7DknLMRU0F03tdxsaemjm/qwr1+uGKL
GcO5ZAJi1yBbjSN36xYAtiuco2htj42y6DrHEDFkEy3xbP/Iy9pgjHEqE2TD
qTq/pAcEbi9xe5Y6S2FftwMFZLtjwBUsCAnLbXAyY950qR62FCnlK7HV0l7o
XX8zXn4jXVOM8ifozc9mtwnkDWf6JMVvXPFMVHRDhOKGf3mrSKZJnaVKjXqG
DUsgX92xEe5Hg/iQjF+lqxrze/+UuAMiFiY3WXiOOWgbUafHtZ62WFKxrubk
EK10Um8oo7dvKfDcGUU7nT6wMQQydNsSVYkuxU5X9rqEO/9yZl8aXAMfg7wG
c/iMrqi7h0UkPm0ui3mgWGAkI8IAmIWdS16x2s6sYdzHj0zBYQEmhnrkdm9D
AmWOaGI5xQ8xT0UF+SVBzuXsryrXyus5gnMHNOCOfmSmmpQ8Ju2gUi9voaLi
gX+MhyDBMAiLdyd77aaP04iQD/JwkVDTQg6BswyCsg0uIq8TvXtkw98X3BdV
ub+w+Pc2425UXhPSEbfOWVNhhZodzAYrzkSogNSQmSc19vpEqcVU+PdiK9fl
wmdm5eEio7lBqhCPOygTT0YJJ3U2LnAjmD/O8PjNkAodckL0DViofNXbL9YF
Vua60y/HuE5CXlaidXoEkLb86X3Nh0v/rS3E8cBWZXEquyMwTj8Hc9nViYCx
Dutl7tJk2IInn44l7IR5VbQV6sw/2OYffXmjYzr+eGMNcod/WLRc/IrY3tBC
336LXqW9DqRsgQYdw24DxYV6z1xyN3P46wtVexq9oCmLZ7kKePfIHKXmKM3g
fnHc6vXrzhyMWt7hOtFYd4TCbW94fGvbxIAHiz41hlIsTJGpMx1BAMF3cjbC
5VehVVCEPzyw/3VJrMz8fCDGZWjOR+5tAHItZ8+qnr1hqf0o8jWBOITm485X
n4nrkCR+XmFuEe6GIZyC1swgS3nM1H7yI7ZEsvTaW7G842P6KX9M+XkKLc9H
T0Wopf4M2U+rTCYQfnjEkkDxyQs+XhUDpfCcjw8ViCF0BveqKrpsre9mh2bZ
Bid6GJYRXtUd53A2l4VgZcNISTIYetv+S7+wA3A6EFH6JxZN3nTRm19K39Fa
j23obRmzmJH4qMVdOIWJHurOD2mv32f6sQ4ZBSJtnIdG7T0LJNDpYKfyrehP
Bw7y1J2lUBbi7wJPYuWdiZAO5xQzsGiBfq2pYcdm0dMxwe/Y2bCAqcz7YDR4
hpCkI1Zd73gfJrnVZ1526DnqenCcdD2qFL0y8CRXpj2C3T2S6zLFKoEyVq6u
6GK7nujM9cERzbAk6+Xw4LsI89zDjMUES6UGXEiBIxVLG/UzDxwz6ygWsgSF
nxs16CHfdujbbfUgAxHLDyczRkm9VE7ERCwa/QzhLfcjzQ9gbm7Kfi0/w5gd
GCM4Op9Q6jvNUfH4SB53nt4jUb64red0j77RKsbvFhWvveNhyTY5PHpn5w9H
WsSBJIwJ8QbWWxwM+3ep4bZo/DXwIDyRvK6iBKE2dfskHE8T6tVXSzz6fvhH
2S8+m6UhcFlONl9oxsn6sNRnsyYkbc/steFLqYobU29OPJYZYP49N9yuYB2j
KnpehgVjapQguLuF1p5hZShQ+B2/SGoIh1Zh4jFIytMgluakYZ4p1ILE+lt6
TpCDyYnw5rnzEdgDA6tEVwRVALaFGtYU5Q9p4pS6E5ePxXoH3AGzEU8f0Bpk
cjiITxIujZQs+j+S5GG/y4WRf3Vv7PSKd+bkYdVSGG77qnb/6VC0wpnjVbiR
if/GaClgzWDRMYVZ0AyxYtkgsRkES+Rgv72bEYFPG4Te68XZCVwMoOec5FK3
J3wiyWi9eIdtSwYW2QuR5YZ84w0ZdKYe2CJjjCEKhgkSs5VUKxv//BwFFMiP
G+f3qiUaKa+VM3sopMn04cYD88+3uYoga3MaHD/S+PCBoCQIn1Mc9o9h2ymN
qVCvtyWdvyggpODjOFfecFS3PJxp8abZ20C1Vqb1FzLaW0O9HNbpX7yqIEC+
gzk7JGWlD2XIjv6oKa2ZhiS062f7AcBCTVtGsTLfOJSb84MEi82kHDyb1Fdb
jE/9aWLbV44qziz2NqTpnpdkZoDBLQ2olg7mQtFlbS1IEc8EhmZrtVitUqr4
uz57w48Kb4v51vEbAxjWxlLjUZSnTZyboIOG401wwRP7gKYn1MFOhQkjBBMQ
1Zvzz4GaQMwyj1Vyme6pcBk8GmfOEaya4v6jUHk25N0HI57sqNlsBK4dRBdV
9jivelAAzkcz7HMQHlpYbGxBPUC2c3Jexwf6ShB+qmVTbVWy1a4suR6lkLrX
mLkgZP2cbSDc7J4IbWHMM9l9SgkRzJDpv3+BM5MIlnz+vX9jAeyr88v1QQ5k
2AsiEYuK3tgDZufzG/FpKVby74kggB9p/JgXN8Goe133suhuJ/3M9ICyVEYn
YWF5umfFPCitTnfXDoyIcWv+qKKAwO0Dv0G897lDhb/l3C+10Dza2xFQko76
ZA9aOjXR9vm6/LIVn/YjK/tG50mlmcVL0fr08Hu7X7OXvnKiEwGRjz1AF4K8
bnU9rq+FJAS/TWlg0vmT5BldRtu4h54VW7c4xrJNw9Pv1q1t1XHSIiTb2lLn
Ox8QoWeJt0ROxX8wNd224mr8q32V2+3qV8+Da1Sxu9axT3inp2W5yjqHsh9d
9cL3xoV9/UNfDtrLpwXOJxJCVvNAM2d8pwFn2y0Ual/8k32kx2Bl46kmT4qZ
Jz3ZdhwpWtJGZZcIwE/lAEFXdw207/Wy+r57l9kc8Cu8ht8KPwW9qSvjXvFV
3H9TZb28BIgJ+iLLPYGmZ01oN1SziIW34fyfespTlmXzupNH8XerIHV4Lh0q
Rll5MLUnStTNKbnbUVCpm+B8D7PoW/bbwjDW7sLrBQYkJUJVgZMRBoa9oH5M
tXHxyqOq2wRWxnIzhte3j9adw7VbzdaCI+nLhIkIsIC+zKDZSFGzCuTgOeXv
8ZkN6kGM7Tf1RErRMtR7hESOMPjMEgVTQU1lHqptcq8JquoplgXJbI8aohxK
/XZuNf9nMWa+49b4AE5Z2Fo2xVBJ+DAju/kKm21mdJMV5se6oS9mYImvlPox
j4TGiaeFmB/n/m3kPV0pBOw3nTdXNkRtHJ7QChn+QC9JzeHHI++gFUrSSiBw
XHJfSwoKwFM9NlCnP4oYRg+DT6yCvyK6SNzOP7IlU6io7ZRmR/aDVMGrXQkK
mBTAoNLmaLL/P1nDv21VuZsNQmKNz89Gbwaw7aSItB2plU+ehmV3e0oS1eqL
sEHU9Xg7pTbc2PHzwwVcvmllUa9UXhiLuZpDMis76APxIA81ujyAAEXXnN7n
tuwY8Q/CtTYzcepkAgMOW7C8VRo6Te0lWkOWPmuirb5/xQvR9rDEa5hS9q1n
YsKKonDry1B5YPgAT9wjkjy3E51lfXY906nuRJftL9QXoMnfBwi0Tvq30sYg
2872enA+tpk+rOd8wGv9hjjGjTtFSzPRC6lHySXrdn0FQSFbY6NrDXyv9bsn
PkIocsNrpsH3GNirOnShpM2px+MxnPJBTNA18u+JJzU5sTYBtAACdSXYRwLi
rvXr4iV1LXS4twGnW1DiiFI6dmdzZCyq3VO5MrF5yiTewFbRA2q8gXkLTfQb
3TeoW+GuIYmU9evL28JlqcNpB6NLmB89SlEEDX5SpXUimUN+s1NjW+xb7Ags
JvaRgC0ExJIqe0h0M63b+wLkpAc9SNKxLZL/40tYwLGRSLgyNKbN6xEMkqxA
d59OTiff8+8zHiE3Z2F6TrUUWpWXtXoNIykmBjMlJYHQZveeF1hRkB4YLGpt
smZBigifcLEl42R3soMOzxvO6K9oaqnGszlM6tuae5lODu/TX8AoweQ+m7cF
o+YmseZTa4qWbe7heG7Ugq+Q8zg4tlhF4yusdsgM8yuPrmhJ7HFeVj2udHt5
OqMIB2sk5YVXVxAsLaUl6zOpNscPg83agMcGftsmbNvIMrDiKwyzgAYq7903
lQv084uvXEK8XriFqVrAsfJ1Nv7NHxJogUJ6czJKqqkvdhH3Glt0MOru0M8M
OyLrGuzmfCMsaUf+2gCQmgD0XBdFwrB0pt/ES7KXYiZrKHf72hykyBk5GJ0b
qMPWmsJ3q4uFrGBlL6sK/NYWYfesJZK/DySAPpuDQAVBCPipEj54fDzIZTV0
ISiJPqO6OJVPTR7ehsykUvAovM0DHgNZAnMHQwNOHmxzKnHUZ9ac9T8YV8fL
0IkIyRE2WFKB3LcMFmQsqHALTvJQ+DeSJll3jQ89GW55jNaTOELTWWKLvaTD
WKbEV2cpW/jBnfdaI7dHLRBXqWhLkLvpxymvh6XoLyurn/VFdnCZCHsa4z5G
EeHrxhPvpA+7bxQqDryGBk8oL7uSLDbWQhuq+Sr0fd9SOf/1fp+Tec4H6OU0
E7gEV5IlV0ncRzLA6XoilkH8om/i43GzEvKFHY0zFmXyuxq72jEuPjwaX97j
Yof14O27F/xRS2J5OAJcpvfRRfS0OLWbiZ0mHDgAuAs51DY72QlnEsQGTktW
lO7AyVZ6eeuqEPvVwdu9GpPKOVNoRdQUlxF486W2QHc1MnebA25Nfj3ss+Pf
S3j6cAnZUyG209KyH5y0bcXVs/cfgD1nSKcX3gY/VhVefnyMBULBCJd1MF1H
0cn1weuSaYTIhulncMEhYK6dRl/Wf9ln03I+EqM8wsc5dq4BgELmTdjYYAtp
Avy7lm+9pphLJjAOXLjmqX33MG0DiBnxIyEpZHX5a4e2xIpcZOFcXIFBWU3a
13n5uWsGg6OhiCPrnxPNhKhsZVi+ar6K3rZrCECcGp3j/PWubkXeEw31tIdU
HVRr3qnitJYRI4eQOqylQTcuAJFDzosPfbpygEyfjCIV0xgPPoSntvM5Ad4z
G888h5M06NE4QKCwcsmFVCmSE1vrwBapnLqjaRnxHq5tAMHEuml+Pm6b6uZK
Tm2ZiqKkXHxqxb4nZ2UIG13OL0xwhQZ+LM02K3zcPf5A+beK1gklbLLtrpXt
PDOEfGYsvEhxUYyM6ifYnDTPmskVuSvLfRnAztkAH+eaGowvzxCuYheAreGt
CTYluMZpxiREm2ZdgPSGHkkW/n9CFgp3ScTGoPBSIiYKiYJL1itrCvNrT350
ZKfmLMC0uPtNyakOsBta/oiEzG3us2SwJU+DG3MZ6JpUCoATd0jIWJpjII8N
B3YsnYahmMRvWcPHt8aVq3D6zzR9asjYM2m7XIXjkZpeUgvbOSwc0G3APcqw
uIjpMtBQRxPxN/LBl9tJg5Q76oXY6LcbUUBwnZ9yLcY5GN3rv22R1EObAlg5
CF/mtqfmPsGPr4Pkc8ffh44vy1iTdjrcq3bqhWU7zNhS0ri3BOWu4IMGgckx
WqtaCOIs8HtmxVY0cx7CC882//CBeRKOaIF3BXYh2w080K/qfdw9BtTzTEME
bEqct4+ruxjhSGPFabdZtLCJ+3wMl4J0Ejygo6raN5sHdByqHd0IngCAMhh5
oCGDJZcPMxavasGbK12yAJc3bulBhCTATd0+NBPAI9yz96M2CXrU5zvcTChF
X6YA+7J6Em5kDQc51L5VDbNpBpGofJZ68e91mcDAMtgL6ILDAnM74B5Ri3BW
3JxYX3XrsuZHy9BDGPklfEmuWT+hUXRLJmnp2Tgxhd5uR3dqjhsV3pViZ68Y
jY1c7uxt2Dvf32WXen5nUZh0EI8KrMwnpKH9YZ8O5gNiNXI92ZgMLnbdVo+Q
KEcKH4duzAK/MjmvNY1EMxWt/08zQJpUNS4RGimGn/BZV+AsctyMjNpI7RS0
0uHOYWtuaFkXO98nH2exapafit7lbyT/y3sAcmXKD8wuLMy0zjwAOpjtxjtl
yIQoDMk97Xoxggrby7Ub1U9NSfSpAu4HBG1fqXHNBo2jLXdtOeb2s6Y2+Qqw
TCNfgYV92BzEOxIQtE5u55I9AE8X1I+HQHEx08ZSBda7NJ/r9O35ntQbyWcH
ZSmcWTKt5zmc3rAFgnClkaOhIDWazsqaxpSclQIVSUkCaD2BCStlD4QY3+OW
sOEhyVnfGMLQ2cbgIAHhNtCxqExj3+46VR/D1NcUiNBYySdQjPyx7S3twlja
c0YQ0fVJP337p6VPb/jolz3MppqTtsbqxI+0btJS7KiOnWqIamYwn0+bnku6
xsotLBNwb8WsSk3I/N1FUDWAtXRZYN9z4belJIUgLcLYxh9rhuZ1bYBmZd+z
AZzwJIX8dayca3CBLPBBp4jn5/2fYzQBuFEhHBdfqveuBMFyzvWRjaGQVAOc
Fm1dt/sTG3+OAgYsBRsNB7GpTDKVgvcLYHJDAAiCnbSTjji963lfbtFOuSEr
+ivvbnj5knqbgU7dS/tKrgGmNn9RTLJJodPtNhN+DWye0trrjeqoHkWkp8cZ
B7G9g5qXmyrJ58MWf0cuVwZ1wlXbry8qRLxeyLaZjOC53I/J6T66ipfH9s/0
uwV8PrLyiQQw8sd5FRSVtfJDIUbFSwg7wKLOPeu5vZAGzD0rMu6fFihCVehM
BbuISxAey+zvLwV52ZffftVhzBJFwGDFUJApYFrPmLQonqzXBQ9N4zBt0uer
PPVbB5SAgTiLtXsV7xApfZqBoAEPoXLpT4dphnsRf0qNvt4ztAlG6VVdydHu
+66mKBBt/lFhaolsI1I+R9VnOR1g+XCMWkfByuARVIVHm35nbWD0ZhN4ldeK
csV6pEQ5pzb7jL68NLpQ4XRmRUfAiQCK1Kwbw+UT+Mtf/3Ln3feK1ZRS56RO
pHnQWzznsJ4oN4wmSRDMokd0Y5D9PqQVZEqCbVqdH4SJtR6AJEo7eOfHcEWw
gOo+xMDCoRCiyeA+BZtL2qliKXEhV3O+rcKFhklowS1oyEvW58AJkj8EWl18
Q+aK34P+YKdvDRlczSrGBi0+WGF6NLQohx/Xr8a3y0Q60GqRSXmMe5UJdnAy
FHLiI90VfeiSimhvgQlSbiKkT6lxSqAMwF62o57kvsoA+zUMITlmDntfNExY
c3Gg2uDK/QBgEuamtgLItWv/r7ESlLIfh0WInUb/A1s2vNDp4NhHHgUhTtOh
DXJ08KgqoO1x4tEJ45UoAa4mIHs9iTtCGaEWc3yb4UCmilrDiwPsZuhP1XIW
Ylf6sX+Sla3mM4nOOY9ThM0usQlw2ZVMOBMETkg4uIt1NE3LxRM5A5ypGkpI
HTZmA/lHzSl3HaN/xVlALB/JX7n4RxHpijTY1fQLVKSa5VCtpU/jF6ZmXrPr
5LKDgW3XcgWE8iCWboJIpwgKQWnUxlCNUkCa/hCy9yoowfnseGtoNIi6K1cs
AWVHRU7zAOGA5FoUfMPPcawgKmzWjiyh5TyNL04MFdo+DJoE2DSd7f6T8LYA
YyqBoMhciHt+aNwsOikvgKUWsnTZNAaCYnGFyo6BjLd45J/hl9w3vN7mmH8h
FYD2+gyfCOpCRg94fAkm+iylXLxkMyfUTuHAfOFwo7+PGYMdo+6rGQhGhmyc
drDij/lgY7qlQBBOsdKJNbnhqsdb60pY1lBFxGav1oINbCeiJU6Cu19g/mLv
79XK5jsvPobQHY7a0M8NVmBn4Qzy4QubANX6DW2G+Ec/FaBYdkREQMQq/M3E
4VqE7DVpWvv68ZRzkIMJxe8m7PDRWXrWfZYemSeRMh5piUxNdFgwO/J1MHnC
mpKxHFqOPMwpZ2iMu/V8pyuwjvJcU4ARa5oGljIJ7PjpWRvO+43V0u2jqED8
ZLG/wqgXmXNjKsI46rdIIov0LxxBuHdMg2reXQ22/bVSDWx0cIVHnzNAd0+C
H0VGb27HAXAFNbP1gcs3LuVIxjz6p4yVc7llC1BrcYYQrwoBpWIZn+Kjmzxq
iYbZ2zG3HjFUedVcG+Yec07Z5IhEv3u0mSxNopLCt+1VKK+LF9gAMnvln1U4
QJCU5Vbe2vY0ChAcK7icBk+SU8lYiFmK7CBDfi7ydT8LnlcTnNcBq/RMkczM
Cdjtc1fzC+5ZkKGW4/SvDZ4HuFq2Wxro0SoVUVlbE3AYJIa6QaLtZBz1uYjW
Zi4cLEAevHhG3I4qE9/IF4aUW74MA4S3T5JiTt5Au14ogFttr2Z97bpQJivT
x9hJ/qJfez4srxAVul9ShmZxdBAiSIL2qdyFVWtoSrlxin8/3ZBeo3EVOqdM
7gf9OwEntloSERPRmIecNa9MUTzDUi8KD+Oea+e1uwevj/WWuQcQuXx1AM05
fT6NMRZpz8U9l/Tng6r+4Ywk+pMS2XRHV1T6QI6mOMkURCXyNobBschniF+L
S0VW5Wlzvg1lNVUg/bhTd0V9nVAcA8t2N/AMAiJrRZhj7WtnauaU/b03BBgl
mTwRVi1ofA9mPyTs6rVa5210LxuO8hO+/TFMzn7I1SRJ9hUN0j6dzt1Hs3/m
/NhCo7aob+rRSz0WXL1gR8UNHaSuLTWlb4ePqbOXktSgIiPWDSltHNVhyVl4
ktauVwVmA8Po7qeIDlPV7leZs91Mrt4JKLefpq5TaYHxRnButDVd20AiHcMD
uXWIYAiso97b1W+5H9dN231mAtlVfphS6NZ7bDLnim3sKkEpNas+ox0n4uYk
mLNOvnQHa/IfKOfRJHr1+Vx5QhmWbMDIaYAnl9sLofVbk7SKxteLFOdF096z
LamLLPQKw2ss1FvTez6qYKsiF9VxrLJRZG0hf/U9eDQFFGgoK2uI6Sy9coW1
+44wXVQmz5N3eJRhk2mBLWlpXjuhgNIxx8Oyzfti+2Z6csncW2Ehe0Qh7ydt
HPC2ihd0MSocmEcGKZacukw6WtkCwwTpaEb1TY45Gwy+ehoyW9STNySWWHlq
5Mp8x7MQZqKeyZbd55rFDHZmIQKm8VajbNRO4BOIfYBEZyy56eryEgiXby2/
lCZU5nbBqNzVtDuLZaDwvt75WaCsE2MvW1dNkbtaB11UvQG4ebxv0BC+7AFl
Y96OWsmzR3cLvgtni98P3JPmlZdrtCwKHjP5g1V2OYEyCZof7B+T7k2gZa9W
IutA9x81HCU4CDI/SNy016PuWHXWv9ucNidgkXxZ7B4k0A2iwIjKcIV2YoEE
J09xL9lTt23MuS/BC7yReOIWhknH5XtzDg/LNqy7PuTZcyR2i96v54tXbFqA
x4q08qwWWqGaXUn5M7LJwCQpgR5gBRKMMvqOOycyQeLH4qRBiHD42H6im+Yh
d6E+T0kcAfO5LezQLw956n2XpGo0xG6ae+GBP5cbr7e6LGw0XBpSImvMK0dB
Gz1qsA2hpl/MZODWhmG3IIXfNNrg99LgH5yVS651kztNtlu0xPHGX5zKTEia
m7AOyBZu7mVZdT/zoFkCixLrCX75gWdJ0EepqjISUimE+32IjkFgWEIXPprl
JYPpH29sjyxoeeqz3pgp3UjWKlyV4z0dol4nQcfaYmb8l2dZBQAQmY5HPI2s
ZD8UqdSC3T8bWPzexqLGY/McTIDwaMvby4KXkQemUoiqMFZrsRXCioPeMmxG
CKj6HLpFA/2flT7kDCE6Y2lZ8+zgEU3rOpNI8xJoZWkhdOcBSXB+yPmGxztY
hcWN/v+tchbTAkWjpPXLBF3J7IEPI99Pcv/pwl1imtTuC+TYw+HgboEtG6Fv
/VRuMDVoOeuwRJh7Rd8Qz0q0sIVmo65mCn1LLVbnOP+Yi3yRB+5FBr1hyn5E
Z5HcCqak/qm0WcCU/OMy4pVqC2iI2Y5PhNwQzJ+CmNbaDm8WJxJgnFsE420n
iGzkN7XTa7PHQ3pUj82Kp5KSfrbw8eRvRr9DdTN2jUR6yeJaCVuRFjoiKTOf
I0kEXH1oE0ebUOnXNVkbv7OEN8i3xcm+xZ1u0xi1TaBG9Qe/Cfl88AcgJdbA
Z8weFBLFpqr01e0FmlP9B8f4KTK4ZAT2f/hWJSKEXIEMASD4iMO7VxWyT6km
H+MzKAcm+drRv7OJszGmI3H3ZGBmaVUiqAfLDCZ4hE8WLWKk60zV8UULVx6L
Cn1XAiI0YkdslWHdb3LfNH7bvsQhHZLZ02ZzXl2qz3V7yLZjVAfqx5EC2sCI
ATbZw8+De2z+2aT8C5LAgtc5N5xM0oeEtHKemMbnSsZKW3RYQvmlCjPv8sPW
eHgQJGlyM4Owmcv6jpEEGAEV/1rNyl6EPp/IeCYiCh7gYobtjer6Xk3mZExp
Z1vsIIJVsRFk5UqVzAdCD8y5z0s0/o1MZHGnguliwSWP+1IBmdXT9U+CfHPW
7qR9+gDyJEoHsWr++I8xAmQk8pcXgCWc6N1zpN3hTAqzbFlCmHf/zK0pq1fB
b25mdQceL2F6eiLCS7hEx80vAtwtfZR0fvKHfq7hBNYD6ALEfv1TwFdkOgEO
HjQcNabtlbxDlghLybCrZ4rnLjiGNEmYWPHSHLs/ZiFbrsamnNVn2yQnG6xh
B0PUW0WGKZS931uAq57DMcLqzJ0+Yf/UqWPgUrW8lfvmHIwvDgjTh32cZYd/
JQhTpKmHudbu/9RvhMKBsPGY4/k32oQszGSPIoFkaxoHQiO4AX4UZsCxNMx8
drCA7HCcUuCC1gtEDAYs3B0HWxvvx7Onu5FYDRRqqSGO4pW2dBUCU4TkNffV
im8LsZvom1LNlH7qUR93X1DoSV2X2FptA24AduyBVxBztlTiy4KvKoMU4i7J
yuOsF50nKolbaiL9HkUinVJWgJo0PVitue2ztNj8LqxseP8FnGy7MaD1QDRo
juppbzjT1knkFULzaWmUSemuCRikW4pCKRhH0tHJoOa1VcHWN/44ozsaXjdO
j3dqm8877pHII7HcTKUo7s5hCLwQGt95MZ1Av06tQGspVZBpv4u0B7sK0hb8
pFKC31TGEkrSicxrnT7OAm3O/UG6JdawX/GdvInja5HYF79F4dGtiu136e0c
uLCK+iOZaietw3SwF1FrDrq8oBBcUFObwwDzav076R1iS3c6rVEi7HG1aVu8
R2M/QGv4kdxxZlZiY1I1vjmDJTJtuveUAL46Un3g3prluX16nw6ETEffLY6Q
lFuerrFSD1pH2ASVf1BA6HWRRJUmN3+AbdJ2XrXxz6PUS0ZPyVqXJVtZsO49
YJfaZL7Y5kP6+9f90mURL94AVer5J+rlkcZWOf5a6S6NB21fUeE4jX2Q14I4
X57BUzBDwMlTmCyBH2Gu1PSjgqqwaNlcqRhXlpS5uwM49aa5zk8Nmm4oKc1x
udQfxDZMgN1S9F5XdqWwE3/Ck7mDQQVsdJBBqkb1IboYP0bQUG3XcOqBmdIo
fL3nAP/hnhOvEwTlV3vV5cHhw/5+Wsu0h9KjUCuRsaImorlNhrX5QkXZUz2B
50eHrKLRk4S6+BsXcRb+bG//PFeHcxcZO4DSPWKJZdGpYuw/ajji4Qdpt0Tc
e7onWrSbzKM2Y2P7hlkaZpMC7PMVSNDWbGd06e3qbBKuQwKy3OzsApQ0hx4m
fKfyp8xMXtPF5H7jr6JpKhjKzyaKLLtPsEbxY9WUG8asMr9hx535RYLcQEBK
1XnHQXufpjOEs/zjJ2zZGMeZ8kViyoWdzFVlcaH1MUBLQfqOXCtd0AvWmjgB
1di+RzUAGDzg38Ky4E7SkZ8AkP1ReV9M7k2hP6amxYyDMmllYQPSGmCTdsBx
YOFutW23Oyi56GWqpp7/9KI4LmiKwbNYg0J/JDBrGbaJSEInoYy92gl3j4jZ
0BvhGYlU53JxUCCyGv/zv9F3Vcl2E0eg8lJkl4JnNdnn44aQAhnt6Br8REoF
mBfeBZI3chFJCmlEkf3aA8od+/vO85/5YWrdkv4BOPh+974jHXuizw5jyx+l
QJyrGOApGPVe19iN8yyAbx2J+AugFCglSeJKHc5t343hTg2Tuzemnq7YCcXV
EpSEzO/BeSPdZ6sgO+9YWHjyPO2Kc/Um7A3D/CTwaRFONZbCTJduFt/4gjKq
tNka5fWzPR47IFEqja4VD15sC3IUKQJTxjD49PYAdbOD3rBzGZStAPEW3QTU
BGugpuAWG5Ip2uCHWQ96GPGkNqH2l5vttELH0g6pdxApBSGt+OTg8UsdcmJ9
jiMjFVmaayejaqtJE/8VM+Dixv3fVIMIn4sBZZXNhQzFmf7/xap1kNSCr9jz
7GjOH2EhzPJyEwcjjC6tkwW/bUqCctEEXdlr9raOlxd9n4NUytFHvpQ6hKeM
orLFla8a0kPxMzx48r8tgSIacoMP+6r8KxklkGT8+DlAwH1OfKJptO2edlPP
uh6PWOh95VQpwSH6XvKXireiBJmphbrXOon1ygAFq8M1Mtuz2h1A8+LDrPCp
WtHNSFvjXmLYL7/EHw40qulaeGztu9x2t4OqIFpvHKH3CrddipchR9ETDLcX
29iUBXz/Wk7bHePnbhzg2ZI93MarYl4UP3cflQE5m4Um5KP9WGVVCAW6aUAD
8TeZ9ucsmJykOohYIdMkB86QInypk213JCgFvzlFoJ3Lb9Io16o4zy6ABZIu
xUaP0oVqCbenMPpS5gYUtJXHt/obCb/A3lXBJPSRRu4Pq+O+PY4FKfiegHN3
6l4lDWwWglhr0XHZ92FUJsMnzk8XBDMJ7HpOuj3HMgrJmn21n3lujRownh5+
KQoANMnY5Z1xvtI3ZES8X3ryGfEuTa5Gs/jYC5KARaToDAZBvPHRhvesuM4K
BvY3lV2Fu9po+u2/uusD9OmID33053LJNdOxOGSXO2l5gIrtN6POD/gmT/nZ
4s2RjVgo6RQ7Hd0xJguLUnoDA24DapuyS/zpiq6sbBYbtQTKl71hZY/kceXx
RyhF0wwRo+Qq4Ba+nF+IaiXdxSrlfUkrMiwQnKmHon9zXTwXWndLWJ4WcOKB
I3IYigf2Qn3ckU4vlPqqKPh3ZSiIZqbvbsSvMuT7gzL0uYgn70tsfboD8c6U
BirI+sk7q5u1YofhsLDab/nTD+0NDdNj/u8r8Pu8t4DUiHx6qSr8PsfQzG1s
/fN1Q3zSwUHa7gBA2raMIgvFbHjgoLxCo5K6A559vdGCuF+rGzXd+0XhORzc
birVYLPTPFhBQmN6m3cFWKLXay5oMUasql3Sw2x3KHd3rF1lH1SRAhhh9tbe
NwLJpQADvtgXh6OoGNJ2Lm6KlzMoTxF2tFTFkF6Pe69np0vV/7wTrd6QbuiL
ReQiZflKAjH25BPFSO3v+2o7zBqjQUXzUSEzY+qmCC8FPD65Ugm91PLclYqa
hMrlhw0Kf6wr4XTscJZRN+I8aQ40rio/Tldu4h0t7gb3ufBSL4efnikar4Ek
NlDsD7f8iiIgt35DF5itZhfmi3+IIwe0XEwfhxDKlrpWZDKp2abh1YTIEEYV
tdtgnnIzHpf9iHX8BNN5TNJEfV00ONXBEJftZhxmuKFL005JhfmUPX6VHBvP
NxdXRRMra94i6quZo8DAF19T+n0DdmMd6w7mYQiMoMZTA0unHgkpKAD0x5zE
6Z7jQ2GcGWYrNw/pCwGgMsIpK4/doY1mAhyGM+o+DcXgYnJN4caMl4+c1UBS
Ylbphw8ygrnlEqCTqzLbCevUJr693dTvv5js6rUpMoBkZmHM8o2nHpViBWSr
0+5r3gpbBjC1SolSN0GTuoLvC487e6XnXaUb+RWz5/n1DW4pr5fCZ7paj+r7
Lw77g5xM0bg5PAgCC3GQrNoVFFcLHZ0wDyYDHxWA2Mja3jOo6Lkopzx2ipZp
IOSdR2aTmx8A8p4LiftLRtHBFSDtK4kyx3932S5VGZWd5hiBrj/AE+8Z2Xy1
oU7itjm5zHx9cCXMvU/VOhTWA61/U9Tg2fnNtqqoUIGJVFOXLuW6XvfO9qr0
0jpBXT3jLSEdCUCB+uFBv0PeSKpTLhZaP6/MHPdK9SiwAhD5ejzHiO+yW+fg
OA/9I2SU7B18RoRAabFFvNY+saLPMWJVQod+o7Kc9lLahO6Aqs5PpWyh9RPc
kLV3xGICRoPFj/Yaqf9CX5whwZsLMrBVCOtaZnvsz0kba6m1nGMxZ74gi/+M
VGKVDaQyVQIvEjwwfxycrkMBikGexFzsKrvxBBBao2PDudN9O+tQoIS5mXgG
KKsOJK378nF2oacQCarl+Nq1QmyTcvMnkTva3fcxj4Tu7/cX68AAdqNBSbaR
OYaKUzeLfXnUXukWlU4Z2dI7f2QEzOvUr2DrWih/mC23LXcWcDj4Qe+Zo5yT
kGBeNMm3pscUX5Vx39N8MhCI8SF9eOach3D1SDvrN9GmgcfpnMJ9KVvtOIbU
Es2Ty7kdmhMBFMveDU4l2r3jGBlRzfKX4P9w3kIGmsQ5O4GhzlDAuFax+51c
dJ5rCb/DeFK5qd/mJUctpFNIy0LsAKpJ175g5pb7rjYNAwLekwYCT9wbRyxk
oL9k64NlDUXBdq1omyVNGpr8miok2hkBA9uYGqQWyiKOV0Cta8uryG4MtRGW
/W/ohR5KNQ3FSPjQlwLyatwUx6MldqUIMWnkb+0YOD9sm8FAe9+Bkbhkp2aX
CC16pdEGb+EQywh8h79crPCyp9ghaz0Y3v8vYDsVpXBU4W63GNpxTwS8Uaam
c8X6ItAkbHi82bFBkQ7bA5ECChrecKFW6MHgKS8O6MdYFj5v4zmZEftxAyL8
OYOMvv7yi7l0al+2d14pT8uUrhVIcVF6I0HyRCB+CeXytkQrMlqysG/pvWL9
7DdbubxGvqZsP9F25Z5vBgPbTGyFBsbNFdvT8v5+WK+Qnn9LOyRz1ZDYlU4g
Oy5KJC6hPZ1NnXJRIKnsWH4GizCxATWldx42sSXtBRO6pMVwQbIeppR+Y1kv
Ky0Cj1ljhJaG2YOXQ4eosQqeO8riDV6qgmVKHlIpK9PfgLCM08Cn3TLZti4B
nQH/y6ehm/EBuONY3fmX78q0ENCZfRkeCfWGZfqGV2NA+9aZNfpUvYkMi1Is
ZXiWs0+l1Mv3yJEKIvX1CnP2c/K0G0iv4ADGDBLQ3yCTyWCDpZJPBMuAdOWc
Au+qwwYjvthN+WYfBjwpxoR7SjwySYZNtJnMmi/+ndhfp9HSShOH33VszcOT
aLuN+4vV5TJNf2x7OQDzBi+VWp8TlZEnuPwb1ztmRzKm0HcVZqiSYSJPqwWY
0sa9GgKALM0jGeTdjSrlh9uzrQ7w1cfK7G5bP53JMF3EfLn5b0oyA/U1H6V5
IHXMUZgN9XNcg7VCcn9xpg0RG4M4OIVQzGdLt5Y6wU567p1CzDUwiZPGp98F
LQipxQds/6CboYGnO6WKg3HzRnuF7qjSHHa24iQWFt4Be/FktCfe7OYoibWe
GZ6rU776J2nAkhly19mfd7pyfHMHBSjGKfHdaZCJfurDrWxssNPh2XmwVTT2
5iHhkDWmkLJNC5uG53u5vleqnH5DZF1PkKQ+O+KjqiI5A76MDAjGLpk/RE6s
D2RghEWPYNjn3+U5m31eRUvvkNUKvcS7auy4mCMxadrJwvjE6QUqJTCT44Tg
FEK4pZcJ572FBNToCJuzThD0EmoPQWCXka0pAugilPm6lug8DERXzg9e09OO
uYBcWIGon7v66EAWkzGJDv/SOobZmdgk300PA9Zh6jmHZbeAQyO7Px7CEGWe
bWgdV6ksyWY+zdRh+ae8jSDRSjX6RbU1YnGGb+GNYU5exWrYY3G7pfj2YXBC
qSE3JJbfxoUiHRqLaw50GaX2WXv/wrHv5M16Z5+oL7sIokGkU/AcuqEbbuPX
1CzvozwB7/2mOtx5SAgsdqeYkgJ/YFGgIVT1RUfPibYwYZFiNx3OfS3S4q2H
wEYme3hFp+LSzn1MVL+SiGaMf6hXhFtvwahCsRyC5pO1o0ecRqjoRhh+MOr7
YbcXW/3Yolg621qHZE8u5FACreiB/+L91DtQa+K9DjG6UZsGYnYLK2fzhyWK
7owWWuf4C0tGpyafiWj1fYOCcBVZ7LZseq3F+VniQ87jBmj8xXpUpMGMUdBP
iyvRfx75gzGpwAMJaAD5eZmPrmE9S3rKHpNriJEz/7S7EgDCt9VZqoF4bbPS
EHCsHWfzJ7v5u1Lap6AtQn6bKBKP68azf1qmL1A70isc1aecDs+ynr3NphHa
5pTTpiedbjzXvSaTRxmvgkJJdIbQwyedG+BWwjfl0Qe8XQQEnBTdQcaI2QtG
/1AvauffDJc+Cj1Y2CGWo4LENaG+lZzYXs5dYXL6kR2J2b/1Nz0v+14tsKvL
bYCGNxUrMY2PRXBilsQ88Be6lmc+g6x0k3E4u8ZgrXc/zTkhlEpa+tCH6q+z
Z92Ghmi45oZaAuqz88Zq7OFuUcOA4hERSfaZ4zpzzvaNmkPAB51Nk2Fm2bwc
4ffNxpHURpC4U/fR8u1dSpXsmCtq3hSQnQmHCFIMePy0qDymLV4rmgkQvsjZ
IVNVVBGwAZzLvhkh1VH/R5K6jB66yg5YLQdHOy2dDoekUgSb3ggFUPDDcWax
B+hCLJydTQgRoV85imyZN8PObgc2fFpZh8eewL7Zh4r9pbsizIx8Ubr80BYE
BhHF4jOD+BzogACSqw7nigb6VdbvKKbunzCxx3xKgPTZOCu52PT1uTUM8Rej
fsXCm/2/hc9l0UyodmgT0VCBgD4lFocklKRTFU7fuH3oxGHMdm7IXeH3P30Z
dR/5qivTPlyzORRX1HuDiUdmv9i63suWVXtY6zzVtPnLIRyO7tfSNgV9zTA7
hgPpqPwz9n2dqgDuKj5W+FQJFjMj2XfiVO+9/ooqIc3OLLCRuMuZq7t2PeK9
2rUB/X0GPgExzgxmcRIUByTB2U7OsnEn+/5/H+cQScK3VuYZ5XsBx7/qvzfO
AZyEvvBhDrD8F0iH2polALXxsWxqnd79jgN17+OBuE3LxM94afg7hAjVzeDL
vpH44S0sLUlq1hNXXOfTlIcw9XDCWkGBtcJNImGUOtiP+qCGXgHYYD+7OnGQ
XA4TQPC3J4X1HuJovWWABwiBCrRTJTIQUSRpNw/jTYtT3gBM/z9YaJw/uOJj
bCLmiJNMpEuKNwL4t/GJTr3rueIpu95OPJcNp4IEBD56yWspZVT1ar55im7l
SL7/HwoJ4plCQED6ilqrc8VABt1M4CHYzaevUH0sTyeqUypWadoBnI7qXzuH
oGc5YQJX6BOvZ9jpTziyvB9gdiHEkXVk001qlAQ2V7aBR0q1lsJbwIjcEhfj
ObWTnAloTQBtK6TGokQbFoH5ftZ6ar315EVPjN3FwOY0eS3KaBsOYF5BfCyX
RJFcVnmkFqWWdt7ZkDSXXf5mfnZsGzoQWtFURjuUc8hsjnYV3ii9VJ3/fD0g
ZA4HkyrE/cYL+JA5q3+ybqdRbO1dbQ1Uws443WdBa0OBOPW3o4yJ+rkHRQ4w
yO5Fz2svjgtbMXajEoSWI4S6N3X8/kJZpnXfwJlHH61dXNHL0KUcbqQrCXkJ
Umg8KLoWfWhncDxN01hk7IZh4rp197Fm3tz6aZ1AhnAkEAEdfVsOE1gNAsC5
AJNdXl6lR7mmYe4BsuGQtIuR1vjk/1g8kJbeF0RsdCJW2jC0oqQ1xvTYpOb2
3WhBuxnZXE7dlBtQJCwk9kZGsOPSNK60PGKmA021sBf5Z+SpNngLUh+5UUJh
mwcPcdHUPVz53k52CieSxpHJffx7hhLdiDOIKI5OmEJwG61/SlMWD07OKgJU
VPbOCWYyDFkbNt02g7ZXGW995i3/2hQHwGA1FMkBp6P9+yXw23raSA2DkWFO
SFmnZQ4VTRVjGUSbUjSuomd0SBKab9qGxTEQsdLbhnN4emOp9DRDgHCwqI3o
3YQI58U5o0jDN157kbMvRYt7gWX4EvmELy+Qc/4WB1cYammAC8lG4xzjdHAK
xiJTtD8aIqLwiYDeJDVzuiguWrkq1kLgu++VR5D1JKbdICYws4x1/mirinhJ
KAecEPQb/06+qBNTrxWCxuRrCh+gEnB9N08DVSIaNqcdReYidbpp/n5zoIYX
RRZh8emS1fQzDmEDKzblZwGKvSHLUOLKw7h8LZdfzFcvU6Np0cYbKMaJcqh8
y4bZ5U6p1/CCAF3N4oJ0TBPDXbsZB4JbPv4BM5fS14uw+CLIhzO51Iix4bEW
4ExjSb6nvBZf9xmFv8JO3lFANXrBx+YfTqUjerb3zOZKuU8D9Hp4NnEkFj7U
ZLgKmmQKzzyFrkLPa7kB5lO14zFe4BfY9Yc+2dtlQb4RhxkbQe/+ogXmlKRV
icfx0gWbOMD7Gn94qDxOJRX6DhLW8I2Phy4331JlVXRVAgKhVS9gso7W3Dv4
e/w4A3CzC+Oma5T8+vtmzZgWNGbkXYFc6OoQQgrNCaa9ZcPTPhe9+HFXzRCz
c6L5r+e8srzhR4jUW/1GCW51pEZs8bCKlcVEL2EgvVadVR6jyvImNBiVytsd
zEMiGOlax+VmXEEQwXp1ExZBvNUphpHpNRUSSCfGqUdkXKy8ZXu6k701jvac
01GXKsCGFT2R/xlLcSfRSdiM/t+H4Y62YUX/9fPSXvyVrnFwA8wYWF4yKhHW
D3Bv8U9WmtNxdjB2J/6WNXea1b+q7flEepj0M7BNTFnQX0haoe9ncQrfNLrf
Xtza+cZ6Y92/j7lEICXmHillJsAGuQxoTWN4uFJjcTRCEndP8mULnikmsUyp
4dtJ5srd28yMxaU7umkuyktmn4hQpXLdOKtR7BGXkAf+6Uaf8K2ghEO/IaPc
VcG1fRm7az9o6U/T1HXcr+9qBKI3FnSnVudxmml4d6pKp/vmiMbmHF6voidD
oL5OYPF2axq2xNPx1D43bBq98+1gVNIevqbgIHOQYi/mmjbsOQNYDdRfC40Z
qdGJX9haekOAZ7WsN+Mw4nLDWQqeM2q8ihy9PPT4jFAKigP9uVW33EulQOfT
I+OHxdpSTwt5/PPLCVS077lGWIkmg/Hmppk32lRC96b/J9Mf2+bs0Ma/2vUn
ep83RC1vGTqJRdlF2iS+9o0OHHf76cO2D3SUOa5toTiExqTiJziZLgvwHHq0
cNAKJLM20SH5aKRRBQfATDIbHgfpstB5YQW7NgTBO/Csa/0C5Yl/dG7u7l0k
F4DFljy/GlYwJdFNON4nO8Ws6ade8pVOlowhiAJTDI7sKPRtqJI5gg3Ah309
P6IfWi8V0c/RG48bQdymjvv0S8tLS8+0d4qD999x3cUVq/MyFEx43p6Q1Myu
mvHn0bpF6ajhPOB1j1+yM2nYq+MydYM/pKxVQUcKylwwcYBzWIBa4Pj252F4
nM90KZAe8SKlBfCDSWi8+LpwckNOk00jPOMboeAyov1bEbfTna1MeF8n+Gr0
vYGLJWDaxJK4VewLxUDkLwGNd50daxqMdK0zl1x9RkPRr6z52A6aFgkIrM0O
+51klXLh3jMde9SkC+Ann4xQPHMmOdL+wzcwHoNSqIibehMMT5HwosjGoCrZ
aplOfiUiOPitdAn8/KS+7idSUWYy21eJHBuALTlFv00U+FBYjJqqIUJr6B1j
zqZwKBgFUkrHgJQxKlv3zYCJMdIWrIRCxt8tdTc+IK3gR8c4UJD9mbV15z/e
KPuYWpdKUjov+P2JmgaL7pSa1AOlbit13N23eeeWFRbofqYb9knEXeqq/0fl
g33OUWkPHPHDp+nt601zjqwQXJ8hBndLOM5Vmu55zv3Oq+xswcjeSxR4bNfU
IhAQCaDhyq5/LQslJ0Z0x0CAW3rNjZHW+VzqiZeDLifL/m4IwT/eZlENSwpG
KgcjrrGIt7O5OwMWtli7yuwCK5KhIQpdGcmindfKqffaAJGD76AxNwttZ0jp
k3ltYAJwVeZBMIV3u3U3E04pKsaZ5rK1p8+jZoAYeu3fDAtwIALfyO1ittcZ
w8tuFVCl5XDX8O1D6C1alRbZG3oFZIL0pD6IeLDU06C8jhuA6oczr9Cspv6S
nJ3Mi0qNZaS3Z+TXqun+YpHWoIJgSM0r2t0HMuu0Ct1zxQNKWwfwYqpxVNys
4+9kPHYZkeH6AovEi7KoxN/9UXHsx0rdx4CtFAdQeFOnq3dF+IP0SiO3nrJJ
adPdYtgE7o0LpotdHF72G03aIWGpVvxY0rhLAZ6t8C/hCRsdVpm+6Ka+FLJP
VbmAsqCQyTd7f81uZRpgbBzoA6vzO/Ej3/YK1LEzsDJhK14s4xr1VlhEdaXk
QG3iLJw77LFuFwp9SHNDZ3F/t83+mTFubew1azZCuGryXirgBKQJoOCeVCfZ
1tI1SHMqQVayHO4AGcOxvT1XO38YPNC+nC48QaJBKzRoa2PuA/fzmOR11UmT
z3IJue77LO4EcIeyxqkbIf82WJP/IXZXC+SDNp84uSJU/Cdv9LP5xLj62/Nb
83YY51cbD4/+1nHsEJEaZI7RkQUmxqqVzltz1o9N2LbSkR4W8PGqD6pvpNRN
uyjWZlH1dfXjgHZkwqCYdzSPeRFvMtOkZrDgkvQ+uTtRB7BqDTxVrqCvAaun
nSIjkphaHNMhFJpP2a12aO61DRbwFLIaZImLPVIoCjmqdqKA0cz7Q8Ikvw6k
PSEVm5kijJZBUykJj08Z+yThqLu2weuRw0TgDrp8esW1NLDQy3Gz78UJDpWG
+/iGOwDOrECuzvfoiqoWWPEy6zMu1eDdS+SEcmXklx6ELGTGlfre/vITzErn
h1rnpZfGGvxWeIgdtLZ4Bxol3vmbC+aQdETG84dW0SiYLuAg3hw1XbFBUr4a
Khi4NmHHASI3bi1iGmrxTqCnf+byFYP9/htpA7NONGav/SsDIE71sOpvvWRI
n6qXpBdOcLkAY5/JZCdYW/Z49p9Z/L3YaYYu94kFFi+luMMUZ6jFrSUBwkX4
BbzvsLNOyFKrvKHNv7+wBtNWEdaP2xMJanZxIea4nUYZGtUGlwdzGY2hyU75
rt6tqSJ32smnhL/NQfQUig9O57PLD17CkuefUnPC/T/QkyLRmZa8vA1gWG5q
vruZelcsh25Bm4M2s1npbN+Ow9lurV1X8FQJHrBiJDMpmzK3OpQrF6HtlDpF
8w/ZoxrInS7kBu8kLIsvPe3wahaiVr+jrhb76/Hb6PJ1ct22x+y6pOc3hWNu
TfC8O3EDNkvj+nUuKB0U8NZh+XTP5VE8C7VpFG91QBCTTdq52m8K3NlvBsCI
H4s3EA/Iy1GOlxobRfyAaCPlVCUhYvNzSncQ1kYrz7eEa4Sjy9sa5e5ePdp9
sX8j7iPEJgYWGqBpiZNNjE2tEb2b+YbmsnQ3eLufD++6A1ESqWpn7r4ydbXU
r7iamXwR2gol6/Poi8X+b26LsPjEibqow5FhXg9I460xiFMMa04O/iVgdQnR
DSEbsdQ/wjFJkhHQWaKKWu17rUtC+cnWljpTUorx8iKGnRQvf6uJj6njBX5z
QhYdXdBF5ynha4OQVA+8r3c6goR4rJ5dJCm5bV97Xe+3+QbNLhLpZqvL5umM
m2Nx38qZjhkuQq+3eN3NJH6W8oB4C9rwgA9iwEQTMAtQOK9bwfGqsEKNmau5
3pNVZHdxB5deD9Cax1cNVYgsvuP98FYwY0FjTaL2yzrUdW/bCSIwvMSFVio0
rSf8Bm+wWXpBTs8xxq/Q5RzOIxUJ91rgKEoaiJqqQn15oGEwZFAY0XFNAQsh
B/Iwh8cCFRLm5mMibE0YbOGGRHOg102aGFJ2DEHU9P2/PRmLiAD4bord4pQz
WNMvjTpithHHKCPONAdLHbyyDeIfpzm0YYXPoF/opKQesKTgCe5WnfFuy47L
3GhrjnW3h8yBPrf3eqYX3xgIVPwW0SQF5daOlCHq1kadQF+imPgf3v/hHNBk
72bZKWyrkQNjb9jp6Bmb/QXyczN3tZQNhImJWm5t14flMh3O4Vw/k6CGbK4+
8zwbUzJie9Ez+S26XnDQqG5iZEJ78ddIpJr2tFLogMAppmcd98pq0ZmiY3CR
Z9WIetOjRU2lF4LDI6+Ccoglg188h5Lzcmo6vvDaT/dYR61CSmx57oG814e7
jIRB/t8DZElemItlWsRtPbrAkLugXLG+Upc2DfyCVrdKLzkbAoO5/w5MgR++
HQpGR5i5IBI3DmYc1eh5yMrm5BSedrLmB7v+hJ1BOSD2TlFhYgjjK3BXGUgh
n2JoWNRCBLaPC8TLQDzNYe3a1AUzGb5h4gpb6RB742MmmFqoSX/cD6OhSQsa
Fe5sXK6dQEB8ykop3BQHqo9fpx1PFwHlIdY6YIv/ez+r4lYI4BkrmujBFUNA
KJIYOTFGOBBsgS5JiMlEHLo0NlqSidAp6norzNA0Q8iPivvu36A1oX10TLSu
IcvgIno/GDPncgPn57wB4KT5HlKKv+k0VB+9iZhCS4zccOcC1/TpA6u1zcrc
1nkA8E2TN5rtZUB2nVaEE9QYUHw5do9+KlxL6qPusT+Sg3/3KIq7WWjEIdzm
r8BRycS7zGqjV1pQkyLnGDqdWphW9+RzMsQhcmFBFSLaUpBtKLcseTwfRx8v
1LKaQE4nzKptDoM2Sh8f/zR5+gLUCpMyTQczpskFlLWWgPcTczTquDCU2beb
SGuFjKct4DfdFkKcQtyjHmCzibzClGIlQGDh2oP0mAVFhT/pHPozNUDJqqhr
tUR4vTBmy9qYGNo6ZUY1NCkR88IjiJ6EAV5Sj3nS2l7zdEhWbP2TtObHbLgl
c/aIJETmWM6M1WeWlSXcJwNJAHkeLoouxVt2v+OiMsqzRNUQ3tdb+Khqf0TU
tMXXOzIdu4FUrOF301gJ9L0K012PxB9znrQdAbTi60MGholCPOrjuG5ja1Wt
6+s6xq7ShEm0e3Q8LgDL3Z7EpaIsev32NLqfdgweyrBlIk1MdkO8Y2V8UFYv
Xcrbmpgzx7hZyGYUuaM0HgknsQTz8BOtmxxggXWT+9q5Ol1AhQxMh7Oahj07
aH6Jd+0xK3JEZIvkvz+nD1ekyII3ELavwUOsd01R7d/95HQydIQTKroSwQjY
8C+JNyfKVQcHNOBxQqjoWiF0i4mHlENQHEJgxwXgzPshdltaF/yZMaAmOYNM
o2WokJ2YLKMU80zxJs76nAzwcx9Bj0zxQpZ6FLVz8/kPolw/uKbIhxvhG/EH
dKZAjFZJUmUKtGWQ/ez3FSsyjqH72rWrYxPXpR6n8X1AFeU9TNaF0ez387kJ
/E928vtZkIyKCGlhKxYVNq8XCtigFZkXLL/1pEDqnEDaAMuvWy0r3evjR9cG
5HmYI6NBK2Fo8L76XEN7MGKTGObKDieuXQROc+vt7yXqyXVjK+R7Hctd676g
DtgH/ZuMCLYH1fTTcpv5Y6P2oydg3MqtSdQSy198C8z7Z2/JrCBc0d9ttKs9
FuB4/s8TFKRrYyR/WsIdL6/rv8gNu8tfAgWecXtO/fee6iFnVRuRnY0VEiuE
bmxhhTXnT9qLFGfYpUyuyAE3tc7qH/Uhn3Rus/VMHaprmKKrejpwHyYx/aRg
ewiLruEcKtwvzTe0BhJk4ojlNLJ1h9gQdkMiaY8HEHO/WnuCfITDdSskC/bp
5+JE/lmZplbRSqw0soh9WF/Fxxwt4SkPvgoyIpmw+9Z+YzShod1s5EZxa/7v
2FZIB0OyALIF4/5/ONXYH9GvE4SM9MR6k68j4FQXrq1KLM6aA7+Lk6ogqcK7
1aIVePEpZ+epoVC9TzLXH1lqHsfhW1FXePSaZxcoGuV6W8MMXn7Uoi6C0Sad
TnuAEoxU8fRlXsU9lIlgw91DTx7j6X4LPyqD6GmYhaDLEnEXrATgD3Q6bnLz
IlG2u6Ozz4aompU1/lcMNVa/z6n19OlRGDuDgs6IM/KMaOvBPHo4007AwIAh
hyc0SQh0pMoKJuLCr9J0AZS0iaT+iRAALXgRz/XPL9Ec16kQLX2BvDp90Xzu
OwFw6ekHP+bt4YgGxkYVYU8oWAjhrVDwAmtnoMnph9UQuuyxl8U1anpqbOnb
IsRvwb/Pmjo8Pv35AEOe6s685Z0e1JjzD2jXgw1a+qpj1MfH0kZScWtkPUu0
pgXhauD+EG+IPUF5bwJFwfaOXxKADKQeirlzcYoNl95KJ9hh8YgntVrneS2r
bxiwWpcMTnjRGWiIKL7lONXHdPXkZTe85nTz6aYx+fokgrIWhLUxX4smrbbY
herjqaTl+aMrK3IA9w6HmINMcjjra6PUbzYFaCIiV/RT6sW4YsZF2iPbMJ/6
2iHE304xo8srNyGovlKs6knnHu0IYSsX4DEDhGtJyE9WkslYtEDLJmiSXBxM
KKmBZhiaqrzee3IyKkzmZGnn/BGt9wV6P+1SUUeC5cCr970lqiKDr9EBY1dQ
TwPanpl+GhH8h/wbe/ymO12l46/nTdyzdJjCvvCGh2JgjEfXY6mqVLdeJzcy
/r8CTTxIUrf4qvSjPBZdcu5stRNhirh/i3q5bw1asOFv/ApLRcA78+WLPkkT
U4elNqZXlNZvLgqZTHeSrzWvw8abaKynRR/DS7aYUk3fZHfUgGsarJ+J5qN1
oOJk4d6Y57a0g2+hljT5ViQctOSAMGnRDe/eMTXWM+2eCotRCUHOW+DDqFu1
tvByMq4obAtX/Xen7vZ4U7M9CJADONeUrmAkleiJ9PvIdSK//qWcKwo05j1P
OrSLL7B99sGjJMJbr3OwcL2RWbd72BSfnke2Gg2suXK65ahuHkNTIrgNgVmG
57Thrb8QhJGJSVq1B7XBUHPYO3uGjBJnrAx4nd8+LnrFrGix0WOyi5v3i9ZT
5QcPZE1XmDuOwPzhWCorBF1keYdA4bI8aXymKUpLbj8IEzrUSV2x5hBq8wnY
wwlJ0cC7qTXykt3YE1uI7wg7RKT2PSY0m3Vk7/A8nHRhKQOoDEhJkEIBb2vp
6OkQR2pyX/6MjH3D6lQ0nKIkjP0dLosWpz7ZtK+VgRKVEnpjivTu62xXFuJL
iJOoyFYG9WtuB9rUmcmUXBEKI1q8lzGetlxoKpSN+YdVe8PfWB14t23oRURP
two17fIZf1qlw7p1Enko3X/bw2fZ25e/7oySMsPWe71wu3w/dauTH5UcmTsX
f7W42WmTXkhaSz/AR+71SSdMgTmJNeDH+JS1qIcNk6UuVDsKWFHvxE89Z3gL
7JqW4Z9R16vaQp/3J7kwqd7pVukotmk0azz86QkbpFZQwFD0ni/ETS/YmO1L
n8UHYkB4aqtD3fLnrkkyP+CFAatdGhgwi8YIgS5NZoNfb+2njLo0rIYQ8Lr/
+NOOPBoQPvka+1EiAvl32hp2F9PV8RH2S64Tr3z0qSFJxvfwmvnferTctqN4
8y3G1S3bJ6ZOY/Du/QAQVkRAG+mnowAUyL6tg7f/rpCm9EXMAX2o6BjoSjAx
FxGOQhQz3cggyUxyZ8ufrexg+xSfkJk6GIo38y8YiPjSdVwsUI4JkfqlXGYy
NRlbUWYs75tD9ZJ6bTbb5YFf0IDbIT90MN1ynD9IvtiMvVn9pre4v3v2FJNA
GlcZXMks7nPwdQ4apO36aZZo9xCcYtxXBHwWW0NEiUVJn5A/SBfsZZx8l34q
AVXxMMmHhn/OI5m7r3+bM3dFlMY+XtyhYdzGoqB+r/7DS0uHmzDTUdh+87Pf
ySVMZ/9BoI3/ZvczvbqnEqCZHuVD4YEj0k4bt+NqHvx2/uIEDsKcsAlwbTTM
Qog+yeBZE5IafdX7mSVyofmAKUh03T0LSCe9VBXMGC7xr0oorkVsz7cZ9EmV
5Rb+B0taNjebPd0JAQ6rKSGGqXD3iyseTAdr2EJvZ4676skwGrgUgV1INHX2
fn5TF+ct1XAqXohrkQ1Rfc8ILfzR4u5W24Zy2PIJdivnfp5Ve/FalR2b/Kix
CXYW7D6ucIMJRpIvfs7/EGBHnRl7s1agZoiloBJvlp7AdeRpSP6daioVop8y
5PffON3r32cVNoQGTaRdYjPhaIIRsvRUnOxe7/CEFAm0FYa0gF/yQCEMG6gL
iL52Ms1HnZmcKj2r/9sw/5uam23/m48AMSZNBrA8w1uiy+x2A4p+F7Xed8iR
rKuBRceaBtSOrfbxBbgaOoiLDT9aOSsEAdywDGMSnKUzucSOfWAhkM69uhWi
8Y2hAiWRFOvYfLIyIAiOzn7Rn0x7JoQnVn4C5SreqCxmPv1oiybS2DDafWtJ
I9PVSrQsioDcHvKQT0yFativqhJX6fMOsEoThmuqrcddeEu2NKFUWtwec5Fm
qORQLegBBjF5nst6gz3akE9k/EqnrhH9KQHcAfWhdHAacxJ+cTBlCYI/tfsy
MPfHZ1BVruSLl2EnmV+5g9NWDnyX8xuvZ0kiSkDeZwtG0X8LafGlUh32Odpo
u2ZkJo5ReKl0RXYVaUqq28lOwFWh6ZUV0Bn7+e9wva8jzuQ6evw7iUoNJiPb
R6+WX0I17irwnL5S2t/dUVUW0gX2QiEN29PBXoIORN8Af8Q6GaC2TTsP7HGj
aOfa/Igd9OdyY5F+W1dmQH7yLtdv8fPg6peu2i+CY9WPfxSImAMlKG4t5T/u
i2NUnVq25PWQ8+CfHyAPXEAF+8PCt+pevvy8nD2zy63CAuAzsJb4PhQ05yVv
WOllD51Ud8sT5zD5kjXEFTMTt5ja9pvZo7AGRCNtAjVi5jlwLjiAinvmJzNe
gNx23N4pC9ZR3nPblQ10k9Fje5DfY9e47b9KinwDpQR5rbslNQ7Nq2rC7lcW
RdeCLN/m0MYAl7j2qiGZiGLw9z6eyhVuW0DjvWoimOsXIXjqS7HzR+ksdYso
3Zm7fNEcqoPwe3lRleA8lY3QZ9MNWpGDpyNFMKVY0sDqGU19qhPJjl5O2IzJ
YBGjxpwYB/weKYI7C0QtbzTU60bdHqEJuMyTUwAwccZK9AdYyPEGpH/+X+L5
vSfv3VSLXeX7Z52LqBVsKrrjdydPVtqSpsOoW5RGsIJR33mZifwhvcoNrKo3
7/c5sjT495KdXek3lh34Opm01GTzjfvKpBSxfYOdtjrrSBsnATNHxblZmVNg
YZa68efGVomQZd/863b1/aybL4uog8I5LcNn2ONu6Az9Zr8HtqdWOH9w3/CO
1m+JKMOcRQY01vhUU6ORwgdg3t0YjcB1Ets5IijKPi+5QErKvR8XW33UqtPv
J5yU2ZG4eAor0jpOayoF9xqnyw3miV3OHC7SQ8Z0NAcKlxtU75Uv9BNC+Rey
uJABnft/KsezNj6DF47+XKBXsqDN9o9oaRc/EhLFgLH9jjVPLM5XkOGuLslF
FwfXGLP7gyXVH1bMPyzwevns3Rl7ZrdMTbR0eEqLpG1Z/xFVK1I+Wr70rouf
f4M1S/TMLzJYuZfNH5Sj+jnT1Ycm/AVllVHtKPdJXIpzuOq9qDOMAtHBsBuD
Bz+tqT6cPLaGJ9MyYYTB01bbjPH2shsSxyWs9FKoBRqVQm5I9WJwvzWLCyga
y/V54J6yGDW/n3srfbt5mxLLaSQV2LWGBoecOYJCdwkDaKA/XYoJoAvmHAI0
f0N986Lwia41ynqBKf830B/UUNcaQ/WomIXrZDvQm+qa00Gg9KzFSU46YeCz
SoeP+Gxz7fZEeDeKYmaZFh3GIbMz0E7RZi0aYwyJZWPWLse4EYR96QOUikHi
szAYTwKwE4H7ev6GPtcie+J5clct0GhjaXji4pZsR9g95Wu2ow6ZpnAQgh78
9hyBQ/cjTQmiQ8U/As1iZRkqy065oI3365wgQ5p/MNX9fq8IJnrJG0HYS3ff
J0lgS3YfllotboWXswdJ2bwK9xO+mG1ncZuK1lMtyhvawHMq0KR/bC0oXX2y
8gzRFWOGrirDHYBAx9Sxv3EywyfHt4/fzXiJAe5RfhXKfPB51YD55V7VA1wU
CpSFkcH1Lv7O2l70tHNpeEnrFg/m8jGPEmctbTFR2hrYK8H0PwmbLZItvHS3
n440OCBASqaHVNfVLqJ1tQHIScoRF/xhaiA5MPDQt/eC6S5Cd4Q6YN72NPp5
haOs9kJfYA96G40xFDcxme+bxqLK8GVVuJUYsE+85cZZV6Djo4ykBFCqKwc5
XFBKhew9aexNRx+jwE4LvAK2l49uN9G2op6PLowg4RrJPsctGYEZG9aAeZWi
Gd9Lu3/aVwzcxYkfSQ5u8x3Eo4oRt48w63XlZkObti1aP7QyiErgt9UWP8CI
ERwa+kuJzQWeP8c4CQww9hcOaPe+mfhcFb8D6cQ82blXZGKV6lab+LC1i07l
i51CxhuFRIwwx+n8wR3i7zU9QeO9I/wYZrwOoxoaNSGZMhwoi7Spk/TpIi1r
130T89+gi8jpvaTZGnLOFg6ef6PEQQB6FiKKPii33usaFWuCSv6BP0CrWOUk
5VuA4bR2N4Xj365y5/kiS+bCBuE758zwHEpFG5vFUIorj5Fpm7wdvV4KfIyC
tbEzBmup+lM7n2JHk1pkYhO8GeKbOw7agSjqXbiWqbp4camwwyKFnzJuVlfk
4mc7G3Y7LOAA9QN77yFLgQB7YKfgSkxPibUJRmvYYwGrTFPondvvbgI8fWEw
aFyB8jmNL8Tr6+rrK208ppwqkZGaYCHIBd6TQG0+VPn9AZw89l1AO63YQCcd
YX18raXelsWoUpnv/z5au7oET+w1twOATTpoj+L6cyUV3r8TLzXIL7qtCiaH
nilsKw1+1C/5/rZhMntFzrmpFRy4dI3dsM4sV5EQ0aGzTCAVXDTAyFjurrK0
CWaUozUdDJg5t2mlKSGYr8e9KyBpd9Q2EL2TIbuTBVCmI93VHq+VSQCG+zgN
PWLUrgkVwt5brru8KDwD3/4yTLOO0vDeK/YLvTMSs0AtVzup9wzCTZ46AmGQ
OsNrsIxUI5R6qRJfPcyA6vMsYS6b2NVOVG4J/KVBcVtvZ5cu20hUBpbbYuNw
rEYl1xz2cU9KHAVmsc3P4nqyuILkPdxBeazmJlu3DJgMakUdXis57HvYkR8G
bjYsDX1Lnq3D7IkNuvffuqXVsMp8SUbX/FNWRwjT+bVGr3nl7EBFfzVsvr7s
k9+kAfHZYu558gtpwquqaO68ZUb5dtbrmGOkZrOhgNaE3as52uMsgkTuRcFO
0miowKQIvUh18vEmfV8oZBzQ+8Pw9tCZ220URlwimK4wQwyinFOVCrV+AYSx
7uJOVUqqXXzqVF+mr9kiDtrpqzSqKfmHCLzIXu0plkjVT6c8U2Be5ejdx/Xf
ICw3gwayYO8WSriHZObj7v+/1rwjyf2uvYYrg4exEEP3Smjk2TKrpTpDPpAk
jX2AuwO3wydIr4mt6B5Gy1InRCarQqKAGrApOnhuvvoiXLYS4sqzdsGlDYQz
2zwQVQL/XI1jsM6IOujRznhk3dkMhlJuU0r7tfwWJ+oB3m5hPF9yXFElhMQd
/MDtnGJmXiWfYRXnM7igKfzr6OZ1hc1pOhU2WDUxkUErU1blq6+fMekSh/v0
bBOpfQqoWrC7WcGjbyJPOe8ziO08F/aYXUGh1RX0Ahq5/+V0X7KH0F9ZZebP
NdrFJUd5XevWM2oaILGJ87Fjfej1yWimZ34BfuuNwlGklv89NDLF+R0M7Ivn
pYDSNN+gEsfrcw8Vx5wDoJxdFFdS4ZyWubMZk7uK1GHDb3VvkYxrcIScv5qd
axWdb5U6jjj9VzuznFzl04coHPxxwZ5Rw7ScBh0XKOgUnufiAC6JqeGZTTAm
VvywWbjholhVwXsLVss4wm3H4QjHG+iAbvqkEuUF/f+O+Z93PD7/0vZUMBAs
LqhMBBXM93HW5W3Mvwah3NvfADvmu0io1y+kILfXzp6urSHNsM9VarqC2Hpv
qsk8gPxhZcvWlmIn6qFn52WC8tigFcWUWgGnYMEfgYsGrhX6Ic55VVXPK+gJ
E5xjBdsQ9eEBzcIRrF9hfON9lVEH4SbMHoSBpx9CxQFJOqQfQM5LHnDbpLLY
mnrabh1TQ6VgY7HAxW59vmq7YK+dOh/XSLIR7fHwoACPybmm9zwnNpZ3IWKr
CDagGT30UczIMDWwp1jMD6K/slDFZ3jslNMk9NDJDiirY1p3wubpv3mODRF2
IirhTOA0f+b01uiCv+xGBO4bEmkJpnQ1sDCjk2q6V670oMGnluLqs79Z65jf
7KNRXctnQLlTrBpOZ3mENkXilLdIym8JJ/6Gpg0U3ylhkmhQfofKUEjeJ5CA
cxQvSIOY1hTu/+D8qLyXwg/UmvYmcN1Uy4eAWF7TrmacIeB8VaVChJtYTu5K
5HnNnS6WdwcA5B6NORqcRddzKLhSRAOYYO9ObLGylQHywJwQocpM/ADq5+gF
54c7U26A0x6rso1+YrKS+Wv/G4P8J6sPfD2DsvODImzRfRj2guh/iJsXVk8U
KFcOCMeutNLE5jtqe+XD/Ccx1yxPYlj5/dDkWdWJ6FUuWb7iIX5Npiak3Y3L
qxsbYdalSSsK0rnziCC3UE+2uCN1ks/41+Kbp7d/L4wVibzjkL1nClz4nOBw
oQWS55hdgrnGIUaF1tqOSuGoyAsLMRiEHNpw/B5GQbjtfLEpx9FWjnJ0UO3U
jOUyOMlECt61/tBrwTbflbtGUNTG9DEJulbN5CdYoECQ9yJAM2CVSLa6t9vW
A1uRiHbFILmoia3R/WGrgMxCRgP2dfQv4PPPAeaZdr62PTxZbjoxlrtzNm4M
PxOH8Yytixi7PglVI89c/Ciu0H7HH9R8ohQ5V4xBF9UIUovHYCn73GfK4xkZ
VLSUXul2gK7YoVkKjIYqvjAXC1fNJa+QZf1RNtmnVqD0fNMZTl89S0LJ2GTv
kC6qVPApoz+V6IFs8Q76iZXSlA5CxMpbCWPuxgyKQHkjNuGLTK9hGcwBtl2o
ePU0zj9TVSNGq/6010UcVuCDD6CCsQZ/ad4xtcvGMSqHzrdn4lRE/L6/u8Lt
AoTCTniYq/G8PHtWzgu281ggh5nnwbrzpAnj+lu1o9K52mU25E04FrcSHNWt
fBMqYB/yxLFMAMyoEJHlth+GuqMML2wCBIwr9zDgvXGJZ/ch4o+fUogXVhl9
/IhSyWeMkA+YGNWQenqpOBzI6ZfB10Y1C/1Hok1uKrBniMv7mKf/DTdKN067
elWdGTm9Krqbezh0EuW1rJDHmrXDmLN9Am7UySqAuwvB5U8sbsADns5JZ914
QESTJ8aGkh6Fkkl2/U9+kAaY20ZOU2aWSwuyBXdVrzelcm68lBfAXxyK3Dgh
o6EH51SGhz/pcrkzYuMSH3XJAw33RokJBuq3gQhHZHU3tqgcUa70Fi4YFO4G
NWyviX7izFfz+tX1rb9Ig7aVQ0hTulCZe2Q3lP0QyYDpp6cfYCSF8du/nOsH
ZZ0hGh+BLRSD4VfllHIv6GyIcIh5StQow3FNXJVtW0U40UfaUHWdZpPAKHhF
jLKrIpq2zOAk8pxip5X8XupwyYd023c88+JW0EF9vfv524Lv1c2J3UV9HzrF
5kKPYKL9jF6q6QI5nwpJ0sWpVimj0hC0/vaxiIYo0mFLkDM1qf9Ng7+6OVi1
ymbXi6cyy8eLOLGYbRIDUkXLE1f5ESXlnarRfxihDBUNli3Y2S8J/bTt13nU
cCXZJWhPYl2Tm4OzrkcpM6AzFn7wMmK/kRk+fN54JLW1MAFLiqhzXT3nq53p
HQelFkXvmnfBJND7WT/7TV6Oy0lacF3+aV8kWMbuDSt7K2ENo69CKtPz7xkm
0auElfYHxEQUBXL+79kl2WM7BiizTeMQB6qWw/73aZ15HQl4RNe/73hiwvgc
gPDOqTuJMjYHvemTTeqNY1rcTcQbTNQRKBRTR5NZaRddteqolsOxndpmnPSY
lmXG0365TuqVrQjO4rZd+48wemy5ico38gFFp+JNL0qdckbMdk07IIUu632l
XX9PFZTNbLbO7V0n6ah5zdTaZdqFndOOoOCkcG/RTXrGwaUv2/pwDIRtnCs4
9AWp7uD5PekWwWxv8PKH2ezdoQAqQHMGeDwYm8cDhWn/e1SoFIh0ESGgrLyU
FutCt99psJXwt+wT6AmBsnX5/A/k8YtxLayM4aEg6IUr6SiBx5HprQBPgBL1
aKOUTCHdcrenLApXc4vOYcexgNHOutjF7fkuUA9hc75fgGeqHfOR9MZwz9Ky
PABSeWrQKzCZrn1obxTKBF/FPQJdWGEJ93AQL6uGjukEXhsj2ZajpyAJ1vHI
NuCKWa/xeDVYQMj8u/pd3e5s07OkARBPObZLhCA9r0Brhi5wVz0hrepIF+tj
mA54bYFUfS0HPUD9wpmmharKF5M8O3eqfNcmeXyq2SXBPfzg5OQTG8e8+h2V
2L8m1L1Kj2rNioYp8EOx66fMcz+JKD+ln65+2AmeBws4E71fD93p6dMS2iiN
47/b6qO9RCv3T0LZkv8Rx1BRCmzsXund+NpjAOphAoCyKEAlUMeEIaBuEcW9
PRpfcngz6rI5IBfBwKnoBt26myWDdj4N70aDRyrI23FaMekOhPVVpG8E35u2
SRSCO2Vo+NB7Bf58r1wYHZ72wmqbEGeFXUqGKiXPr9E+xPpng9aJlkarTZit
wOJtRka6408oMWjVE651KPtX6YUK4H6OmFBUXjoPPPDPVmuYsgUTOsmz+wmw
DujgUoWCUxAxcQO4nbPDRWNXNzZ+Q/PgmLoB+6DzIG0PZXE/fl9sFt29xZHu
+E9sPghCNiN4zJpBgIO0ApD2cB3vrWMB4PqsJs27kB0wxZkrYxTigrzliIwm
LQwjZVNTr3VLeWzoOxrZokbRlgAHjeO3akydxV1GglxThJD8zNM2i0J+Bp7b
bux6UT9weAEAL6fzr9F28aK3KrX1d7VQMAjpFHBIHjMmjE1muegwpnlvvtkO
jhxBUxeT03zkJ30itd6p9/UwwHY0s5V2d6ORyIo9oEarCo/6DYIbiwBlf8g9
y9/yIvSp8W3lrubddaCXL6smXKJLa7sAweHomTP8RlHf7yf9Zc4dwNrZWK/I
nmi37kia1VkLfNGVZhdem06daTt6TbojYSU/VxV5MOdcVxe/a4ZWRmUT6VY6
krfLb58CkX9nQoAkFQuSaxqE4JoEgdlQ3nJlLiz3l5qfin00ZuOrD2XUbkgf
ZoPTbYFswvBO/JMrsY13Wwci+cPyWvjBSWSA2HDofMQcqbyjAslrrElJuA/C
GLbo+Jdi59vX3l/C9NZrW18YhG7Lh/UZgq222LvYHnYyNjRhe4PPsmVYcyKy
7uzyoANSve9SVRZ21pYdchIeyklnsJDESz2Q/A0IdVnfpYPBNSkHHFlolHEb
mOxZWjQ+CtgEdy1AUR5ZEL9sAdanSeV0YtDUwd3uy/4Lvcb+3AWjaAoeNaAU
H5bMiCh93g/p/FDq9WaGcoRtI8h3qr+a2LfxA8gkJ/8vElPXzh5M3yVOxWrU
zRhJIRIHH7gLiqfJaslYKenPAZ99Ry0cEiLky8wh+owNDKQLlDhgoP+/+thr
qpu0sXXOYjbNq/fEp2JVdkfKzLDG/c7fLubIv5MRnb4kQVPK//yqY4tEVKFA
df2MJzh4+fM2ujBFkn2QhROzEWqcgNq2KeqZt0i8x+MhD+Mkkpr39iQyStoU
6k02Okgnp/1Mw9TQcwL0W6iCgPzAU2f0rNJ9YNU//gDVNyjWDCYQjmX0WQ0h
/WtS2D2VGS1CWYNRgrKWgu1Y+H8+ahpnN+f2PMoDLitIDiS5yCf0v3uZ4UPw
FS7oAlCIwWLTbhgR5y9taOz2asjdrfW5Ay50FDXR06YI9XziPP3W6Jn8fomF
grvvY/mAJN+iCkhUUQaSnO31LV0IYNmLmDPOJ0tnspqyxajzPkmLCFN+olPZ
4xgco8QnLz+nOgHqSpo1HOU2ohlrth9vR6CAbVsgy+6CDA4wZWL2qRqYY/c8
JoPKyTYCTdddfI6uV3qNRWmRRGz+IuL+zpOIwNNKasADbxPoTiCPcMF/Rp3E
fXVwfwCp8JwpIeSL073R+cdN1HT2I/CcZ4vfaLsoM2dj3BsdegxWjmync8/i
L0ftHQBWrBDhbqUaZeEzDl1MkAzkVUN94OR2wm7R5bnGrBPTkyCF7MGUbUlP
neNX7kyvmrw7RrZfcBBrBRsKIrc0X9izASnc5BRAOa+isNSFLoMrjlxTc9aW
v9u2pTQ2G2F59nrO97GSx+L1xf2JOrBb4n1O6F0qNe08iJPiD1xyopW0Ixon
IpsNRn/sgYHOnyemKYYvFihE3gj783xMyNCUG2hBNa3KkdJagH04rcomLZnK
ovpBIsfnVZHZrn549o9xudolOWewDAK7tyzVQfBDa4mmVK3JjvkXQXvyfeC4
k/A44klzlgdPO2rxBhGiyU79TaYRQus3iZdsSSURhpmrDpR9x6YxyDfJHsje
ufbkgD3mcV6o5UhB8V8HA0R19HqBE5ER9QFibdvQ7hwJKfKkJGmSgdjeNKSU
bjMErmq6EqGNR1Hz3vRkUnX70UToUFgk8HnFdWKFCnmJw9lHwpej4vA3RbH+
328GclCJvqVNDaqVkYkC3ndhncs+qwgR8gadfgrI4GjLw4/sHBsw94tpa1AM
/5LRaRnbd3pJr901pinuq+YxdsPsrn00AZJyVq64U1x3zyal2fkTEfJ7lUnA
XUH079ZsoYJBuJ87w6CXKYRzNSyovYfXxIoVqazAm23k1TPdK2+1fl49p0nY
k/th9XFYOXbgxkkSNCL1Gpk4mBOn6Nx1HkKhLq19eYStbDJl/YGtLU92WTAf
bC/TsIVaKG6URsNcz4i5Sn2lfgYxwa6y198avlwoBiUC6lj8BP0hzbZkXpjf
u1AowYFTlW3VMMnE8J8ND0vFp+l23mLiH5xeZzhH18hWcZSQsBu+26wVVBXS
/QCE4au/SpxsKTXUwGszTr+w4uryBW/9ZnTtcfo2jf8i9IrGx4NJWKMJdXuw
l0zglbfIRmSk50QIZUBCzO0B5G3IxV6urwEXoTmCuDqfm7Plrj3MEhmftMtS
QYMfG9/vi2VNiVevFEr32ELvj12Rm5pKqaCOvW1rs51bHTM5VMDNd/ioSm4O
9v2fERuam9/YjlEnewh/MKXxLO861sG9+f5Ev4PVp2+ZVejsMFG9G2/vCAL3
2ngv2ljmx2K8JdaL8HBL4TZh4zzwXcnV3M/ConGsmUrsBYqy8Sjwi+Z/6ctx
K1+vDylA0gy6IN+lsMyFS80U80brC/SoB/pZXpaLqQGxTiN2QFmP0a/sptYP
dJVz3kaMXznl8kgb6VnRjMJO87wNux2qb8jX3fjUWQ2L09ACs8BohJKDQCwO
R9EyUKZJqauRId0PQBJIFDEccwGXx4/j13Viccsju+s9FkmvWgBpg8QxtDj/
p/NGarLNBkRkOFleRE32xxqRv0HLbjBjyBKX8Dzitw231Jt+YL/caz14NWPi
zwlZf/ddkPBjbEN+O1+pvTQz1Nvr7aaznjZCEc7xFNry1jTlfx2cFhQssfQa
C3JrNJWjT0uLN0JrQjr3nan/ORxSRe++dgKmDVrwEM9qBgzO+d6Ru+xkLjGY
YdBeVlvL2b1F0Pel2ik2tr7SGJzxhqFOwfH7lOb5gZOd11J4K3OirNuSuXwL
5cqayWYLPVBYDlEVGPyfCsDN6movtY8LYRx56uBZmSyLv9S1MREzOFvttb8G
jSUFbFsokV7LT1okqB6nWRxAfbhxg508RcX5w5tTrfXXcnEmsygwj2B4uAHH
5QOch9gVx6/1UrDaAJAhCH6btOsDoVR0zcwi5YW0hbvFIBp5DRKMycMDPDk6
Kt38otiI3FdVjCQQ8/FX8vmQy9C1F9ZKyx5D4XK7+6iWYNLsuQcBPhqeAY3h
sGFy3jtSfDoVVmC9sGmkRoFYcnl7rQGq5vYUbDP50Ui5D1LiFjxnyfTso6cq
7233/8exZsIMIcEdyaSyx+LT9aamVRIIjM3siPmVZNKDgjh5kZ0P2Uzjqzpe
g/rgpOW7x1i9VPuf+ZDnmbwNFWc5qwS/9Qkj0bu5Go9GSXcVDsDjbigHWVoq
Ek38uKjs5Lg1mLq8gqSbonPPKfgwp8MfUveyTEOvqRB8rk4ec6yK67aVsW8a
sa+EFs//iyoVIsaOarejJWBJ0zs6u5mfVEHh+MYiRrGo+/6bYU6g4U73NZrk
dONlTtPgCZptxKCWEGtxj9QmcqPZPD812aY18f8mFIUfEXkUS3jUP55CTFRi
TWWLd2Dhcqz6nzerDNBGjR00RHQCfQaewvAKC4dBd7G+A/Vk1oxf8uKo66Nd
MspOQa/bDEC3jZpaRBgDyHB+Envu2Ec/E8Z8kSG78DEYZhwo33LpGw5Acia5
uxIC9DdPZixhOx1UUQXkgpwLH91bOQrF0FFWrgB1vk11P5SpADJHgU/HxgNq
XIiRPm72pPFkbYRLz+fQk7Bp+tc64roFRbcARqHrqzUwonR8+IRx+a0uF+n5
hqDXBQHsHRQa1va8bg+Cs3QhREx4DM8SRYipVPLLARwVytVgoI/VwVHCBGmW
wAVrT8DbFZEYtDEryrvta5yHBFYJ8LOq+clv+PnZ8PZfHJr5HBuWJMvQOVQh
wt/xLrjN/eUrOe6CE797kdWVMskh/fWK153yBCxELzkBhJZ+cxnAkz29VX6G
3uzTzhdkV/+/JmCM32JsR5kAtkkeZXR5776tKPmNK6901dz2MhKWsA1VBnnW
IHevLJBXU4mOq88MiJhc4kiZCZqatfK4YJAzMR8wEaKBOuejz22QhDjPPJ7t
3IERxZEDdL73wiCR7sT9K3y83DZWN8X6VxNKuWwVZfThRE2JLXZnB6JNiKNS
8c6hY8iy6WyCy7/ztgo2xdUGPpxQqDGpFcMh6HljiuIz9C8CODtHcS/1j0aB
wakIaAK5/5ThGrKEc9zZYcijAhhnNd+jPXBFEfHrB85Q7koinLu3Wz23s4Qn
ZRTv39ZF3D9pWmzXHluWaeH8HZZAvooA9xvGaaal2quHlPTR51muAksmbONi
AmCdgB8QOvES0hbmbDkTMBmBoQevgO5AVheF+a0gpTGyHV+JWWwi31pDcOfX
4dyIE0VRd+kin73bk600MT79w3/FD8f+OklCAD0wErLaBrznCVE1B0LOnTZB
tBs6Pcadbgixn0IvdQv5/J06IW7SvIWOftlu7kH/dqCKddnHtP5xF9amQdsp
31zjRVzaYINvmGtgz/x2GZ/IIyNYQb3P+FX2FnqtSXfdMAhNWhAVHMjLqvTU
+CTKGcSFOXRCpomGQnEXSnYhtprKi2EicVH+tGFmRSBJOGsTqlWSiP87zAIf
bANPX0aBBlILNIgYGhqkXTRqFdTgZmp7cmx43MYehcuJh9kU7hjRRzJPTIMi
ai8BGc+QGI0lbq3GmB672V0DB7wggMpbf7duH4ND1FP8UNKtdQdcxEGJJAxG
5OiR51OMfiLtqkRFZT0og/TRSyQ/0w7q72iRLd1KIyef4xvdD/ZMto0Vp99P
6ijPzwUsz4FDO9l5TjhC0ogKecnJp258NemaBkEIdM3fSKaO0WznvEOgBlDG
EqoBGmq7KVVU8Dmqvt4E4Tm16EfLye3aIFGPhFdnFai31lDS1ECjNcVbY7zg
rTxn9qOtlgsIhd4fE+/P1evUlrZE0PiR4KNBhPeB2FKQkJebXpGZEqb23EK9
JqOizcUyOEXarECrN/n0S8VoNJ25ZbbVRTnSEqCj2WkmmQz3g8ABnsEOBpuK
k1tXG2xs/5e/a+pu8gYqS7Mv7CBBxc6mp1BVpWJZkgqVQW4GRB7bILx39jvx
ZrkUwDb+OBf2Na8lbbuE8m7fkaLiREZoGBFtL85coLs3ZLK57iEUsTwh2xHP
Uan0FIqd+1lBsb6N7Bm6s/YVHAb6yoyn2XxwdXfwq7jbSZFXaij117U4bMZg
bLH+z2k+NYvPKqgdhqtuHp2bttGSZbuZLA+RM2alNjlshfb1bz6cxe+Ua99C
ujdebCXPWc5p1fvGx9LpnD5De0xGJ2TA5FkSsQgG5I3tMsgWHFRIbTnXTiqI
1tbCfBPYSJr/c3nLwJF4Yi6qpVlWwLzLi2BiEgkfA/aR1WLZYwRzdbr75zRi
EFxZbKzI/0ceJEld0MWyfczISEf5s4Fxy9SRyUub0EtuNStAYxiErBM7Go18
S4gptC7KHr/2tFjDAPTsEVSYfcbaWK9odNqP3A9SN2ddPGn5PW5U5pCvTBUS
UaxVMEI/hB1BU5y4mPJ8ijdyHUT3VEcN6g6Q/ABqX8NigecYh41wXKip/PCh
yDPHdR3pcHMu98m5cp4Yx4HTiqO4SioiMxj3HLUimqdn4A+6rchOjKZ1i46i
00ad/rf7OvNKMmDyE3pQAeQjlo+FUOTUSONoRFWBUu8KXnU5MsMhYXFj7G49
4qh0SW60o14TgaM75aVmIqV2jCUHOzw4+keGlZYcXj7dcuCJNYxPT+ajjsHV
01btsROjJ/GMHm4gmCI3ynawvhwS26nChnXu+0SpKmYrhmhnt3lB9PJpPHzg
nqg+FA95Pd6xLC3b5dt9cgSCpwVprDZ5pxB0YBVo8EV/CZosFdeYbHO/DpJs
oIrGTsjuljKaQNmfgu0+8QsnKc9Ef+LXdqvZnTkRfWR9mao1qbrcnD89wLUk
DCqb2p3vpgQI7e6zPAIESFCv/+tVnke8Q8qy3s/gBSwHJKOR9n1oE0qoNn+8
ydD9KuBo4a+Tk/vP8F04ds9l/eEml/NYpYUkri2RHBleUOjFxi2hsH0VehrZ
j96XbGzqvII3XYyWq/a8h/m6YW0IRWsjsHSbUTEL4GUqvLiZEcyfAsfeYBF/
axtcRp3s4jHMPN/1lgNqRQwOZujQJCBHF8zX+r7KgrHthANlto7jpPj1Swk3
z1+tri+a/f1xmnKosuKoHK8Gk6C6jiH4HVZu37JINQEfWWkugcPljqbeXY1c
uK1VcECCMBqufMh892OV1Uswu+2MVoIjZRnqh9BbUXvWIEX4CAB4yR1FNEfN
6kwU75poN4wZ8OaRyBSD09nPF1/vrw+gudJeM4tAxt7wyoL6X8rZExMI6HkH
HSS1nRveTh+4VRd9ptuaFyz5ua1bcgcfJWD4YMhjZTCDxKV9tbAvXHOMIhsQ
KIF9VW2I8AuIWrLUM8txy6LKHvRX3KSF6LZPYBAM9SX6UtMh2IvTJchPsjvf
w+I1RiJPqYEbkAQU4XjZ897PqKS5BUiap3AhvKDsNgyfyLoFqY0E06884Rsi
+omONQ6GTJ6ZHXpE/8h6hhL4+FexpJHlXBI7sJCid1MiBCfY+Qo9PkQoftrC
XH11rTEUX+rpHy/GYhiagIueVcG8mPx5y/dSbgIkW9yNtNoIap3r7zqv9heX
lySSMrOmf6mi/v5iwpcftsjgm1CQ0SJ7K+TJ7fM/E+lcvBKSeWW4+cBwcBOr
CQGpk4/tywbi5h+2mPM54UPJ9bd3BTxOOfvqaMqarLFPbWgNMb6NRqcAfpqi
eGU8Jr7nkWu92587p18zHKkj8F91QSUb45Lmq7fPPN64YUxwqNoPWw7eG5Qn
pJ71n1P98pGC4S34CnCZ1BdRX9Qjkmds2sxxJxHgzugO3SGqPuB30XKgv8Y9
ppS8D3ounsEsivbeR6B/EhJ6dOSvH6dMmdlb1ZfR7/k5ovRzO6ibvG0M7aji
+NJJq3lmyG7f3kcr65MOPMdwz0TaSXydKGy/mY8U4/x6pxeSqvrQIQt2DpmS
KaLfYzd2EpRoBKYpnUeEXyM3D9oUytjeAHZG1pQWb5ObbKgvWcgOh1DJh1i1
c5zFbll23Uyaa95HZdndc0SsjwNm5qco/MxKxd+M1wvZ0iLL6ZaIb8aOEomM
WXMSjasyEpZ9keGudghwcNOimPe33bQdl3P+sc7WtTAdS8wHhzd9GZuh6fwx
sPs8oLR9n0LpB0k69JUHn8Vw1yJU9ViIZZcpbmDixNIpmjwPQqknwTiDk9XL
dCRexOXWMph/fTqTMBbuCIac2fRhnXsJroDfUOYUiy3dRqmpY/0tEpsxhOIp
tFAmDdYW49L71HGTtvdybB0aHlDhDDvFF30PGaYr/KTXAaEaO3Lf5c53SluM
7u2j4mojsVtIpzaDwWIe/PMcirShgqbrzBlbhxu/Yw3DYISm1r+taqAugIho
hWQIq+cXW9Chq3THzgBLZGCtSay1+EWckHYgN7CFYS9h/exUTDFxAfWtbclo
YXaS/XuRHLMvw8J+vJSpdcR+hbR4ABDXjYmRqXvgqOvOflTtrwiaF7xvWNUN
wWZ4IpXqHSrWzzMiLoM2nMAUCGA5NRp7IzdS/vH1ma/JvX3RWQxK0E/HNBTC
v+Rx7Aa234buqVnBx8qnVl3oxhK9rXDf4MVDgJYITUNv66q9ntzyAY5qmX13
Yqc8YnaQ26a4RGjxyFlaOHR49cs3S6XD4OZ5gze5chO/d/1Cs1Bcp5zrkeoJ
rgmm58TUcq/4umX1FypnMdHq5RcGxSxrQKSoXfU2z4XfPpZXEWkGUennolYW
BirA0KQpaAO2KmKiPPX0IBWSW3rDCMCC9S9794bkEF1rcC5KXRtZaffSxw8b
Dzhz0zbhpp4Sw++K8OK/p2ALsK6GrpSc7jXM78g4FFjTPh9DlJBQALC5oj8s
Eqn3nZ+iN6PWETs2LbTobGSManJv4a4FmDeNEh+c//hn+DzfLMC9O6WPGwnw
xPt6zHLQ3VTVU857d3zrfKpQ6O9cBWAFhkhoZP/BawkqdW1vGDDA3jJ/LJto
1+TEjSdwqHQXX8mRbTb3tjr6NXGQ/pLQT4AgOaJBU0pje0Vf1lQOCKmXO5Cx
0sLJDbLQhp0bfx6lpbaMeMROLVUwMMJ6N1beEC/uMGdKdacz5Wm0v7DWKLSO
RC7+97gZKQ+dPezC0iIB6bZuqRGvOBqxWn2GAUBDFyfLQ7OV/sERKDMG+nEV
MgMmaG775dt87Rn5M64bPEYwHcnzzNGcExj1iLUXnh6Z/NuA1zHtp7KpuS/9
i+RDd5JnZv/IVtcn4aNt2ubL3VI=

`pragma protect end_protected
