// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
BFoeyHFl9VYW2XMQ+HKBu9bmVYh0leq71940apZQK5mf8pEN4uMmNctTixlmt8ym
EM996WURDgMqkC1wwO2pK5UvVtOg3OJWxaZK6n6T0p0EuHUUM9+ORqp0Ypxg7dwn
Ff1i2Wx6QqGVbXrLhlwefXZMDUxWC1cy6Vq0knEFZ7I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7408 )
`pragma protect data_block
lBP14ruW4K9cLiGE0FPTQVbkX3JDXx3cbZqOqjv26nxAKLs8qkTNPJe5WP3cLoIJ
huODSW2uwOpC9i309BsWGV6nJwV/ChQvrvwO0DxvXq7hqMOLBoeUU9DCEFSf2qBr
4A2zOktTFPuSK0V2hr28IbzRFWh+X3KxbGgdfAvyD3tCFEZJVgt5WpB7smqmUToX
au7ai9vnajIkqg2yzFtsvekQz6X1Bw1KVADMVSA06VJZOSTJ4GxIRFJCjFACndI3
zq2w2Zwq0V95bL1+uaw3VAQTYzqxSk8EngF6h6bFy5VeclXMOL8g4BLyL0A3ea9P
YGxJl+XwpZHbVH7wWlgujyUsBytD7kNWf52pbNaHwr8ILGoXuHQ9zV5b3VGhrQAJ
NuyMfiWkkUw+bPzHKIPe/ur+8aSR3jHdcj1p+nYz6rh+Y/bR5xUChV6vy5v4DvkY
8SR3dJIi7TBX4BIwFfiqUO1Q+29xni2ZOhXlalcDEi8p1dz2ZICV/SoZ14TG3m/h
kdWEZSUKhFNoZuutlvcgXHxYEZrODqbebW7ZSkRIQxxTQz7DIom7dwcTjQGPRFbA
am3WkoSIpb98XCAtxG6XZ3QdIMazx2vI6qFx/U28lQUpNcLrMTHVlM6Xy3nVE45w
7Nl6/5F4QP7Ey2TUCM0tw1rCcWGhyOITG65ipDX6XFe40jyyyA4Sw/Fk/mWGdDCh
6gt2ybfcim9Gm3B/9EHVbWQ2V8IHm8AAfXf64+0ihY3URuRlXVrhhGx0IByVGC9z
vMiY9AK/Jv+MaTNn+1n7Bq31XMA8RHfdi4Rq22jLeFTeAjMpCBZZsujtWf3ADw5j
ZwRqrT9TC/4sojmYLbhsF4Gal0xXp5MjB0g9flNicSABT+Uv76LWpsyMs9H2Nhtl
F8T055JIDCpJiLiooeMrzQ9Q81U00sdox6btKqif8caGwUyhBiIabIC8jis8CWe5
slLt1DLv/SgxzsHpjmrkM9yylxAYw1i3iF/ugEYR9rCtNhPRf6xnS6OB3JsmRAKY
3hNGZVGG8UmmCe/n7rCe95TIV/dTITZnBtreNUKIuCnjKTetJdfZ6nDnfT/bjb7x
VmC+a9UabUHAXEwFJ2hMSU0mBv9xSTTG0tr+/3VLVRokl/fgQpcEDvtnoqy49t0F
5rJjRVmpyJLWSS4D0CGL6gXtjGpv9IpfqMBfkm9ECDRE1GaqD6YTU4AwghvQVHNy
5DcaOcfNZFw/AY208rqBxjSCjy01b1StL6Mi/a03VfJDcM7X+mSJNXFRTVDgyChH
/JRSWYAbQNMRtuI8hgKC0/zkZTOxMus2zkjUaSVL2shPIJ9ZHbTu++s6lNprCXt4
cNHQZdJ8F8azSSN7xhdfeMJyn/Yspq6KHlwRbp0lLcv8J/ERGSKBRrTp3hMJhKoo
hDfGoOAc2fC7ZX5+xIcwWi7TTE8KcyVE7xTEwByjcbo7+n4CWtrO/z9XWQBUeJM5
x1PNvprBcl9Fg+3l9nqcKHJLY1POCTFiyGIhI7+KDuL8ycZeXqiOyh08A8sv4CFk
CFGfMtmu71cpiIn+SsgYK3bbY6YOQTTIHI2HP96VAqjowORASj4ccCsrKVu/e/6o
AwDbtkcE112Od2TZlKlPeZ98as46R4eXQEgsaCnEiOC4JdE8xe9TkDjyXcXh0t6V
6wQ0lBuRzlZhSSXOGQ+hI9Kwr70mNHToF73mU8LjVXAcYqD+zpq7ecHIFlU3Ug+j
RDodbDLrdIQfWcLijlD3I30bO877jod4QIXvybUWSXWwxUopvgbpxRy2rKN4ae1L
tyWDyWifJ5H4CyD8zuyK6JgLRcttTrUyx7rY56UqL4dWnzdVYweNs7u9cAuyLQaZ
PTsyow10kfqYZ/5sIhu1UEzNCbFd689GT4QbdSajkKWlA2qZDjzKXK3g//IawlTM
xjFWYlbfKv5n9TFdInz1we+ilgMpH3oO4W6izOptChjosHU5vKDg0S/RLpo8dX79
tcWNZVPMG+B24K0/Njhbw9+Vieq2Z+lHwKDrp0DdMrZTq678V0HQPgu9eyORw5Jf
7AQPvCJ06QtBkNfEK4W9rS5OCPyh5MZ3b4kdusEFEu6JNiOxe8kiG8Axp9sWKeRa
vaSsfbZXJjWctGsD85qzwxvbTBs0f2Ln+18e/zsZelZiE+AmKaUASIMgLC+vs170
dxjUzJUtNXF5V8U9ygBx03+Jg6ihKanfT6tVPCN9x4dcLS5lXwOK4I76i7Lqa2c9
g0OZfqsx5McIBvlm+BQqyQRiVdjKSFmYEXC3rOjGLwGF2RTlGhhrLEUtjYIwE2RN
UbDnZgb3stdE686GFY9leweeLSENVdpMpgLT7ngcNsprrifjCvodECNP6mo2rFTq
7G0OUpTlm3BgGwwF9/zgfMCC8Bi+398Aoxim5LOJBGLFRfycAhlyqjntJQs13CYh
st9QxHDhv/HLEswGZb13da27x/CtB7XzbjvbdG1EKmQOUKqjBQkb00unzFM8oduM
KDKjC9qq2c7dbYYIbNoJ74QUYi4NJMGCTe5NMD2uMEOdGfak89WYJGS9rHw0aRJd
BKge0zNWaucBKjJnfvIsGysuTQcwEIaR8YFeEaWmOQ7SWRv4mZGKkyVJqnsue7Gn
U3nQf9T4lxL8F8rR8EUcu/48B+zg8qdDE62HVwSfEe7q7/FQ6NW6U/daROgJToqn
kFMF/OqSz6DdHgD/ATNPFk3HbyM+AVPtkzNv4sxhdtZlebDsnevuLzODmw6QOlTn
QBQqoE3wDGt+6+apMOOm90nkw3R8Lpaf1K0HSFfSimbtruBqFMZ16Qx5LpcqeM3s
iDhxC9wAhUqerrgwgH1LzZYZNWyUPm37ByY0vW0nWTtpOnGgxxBHiIk5b9Ev2eEI
BTx+6jNTfo9RkL5hHLTMjTtKyk8bNxmD1/meK3C0vX02+APLthPW8rmKZOPX9MIy
9mz2oSmfmm8SizAiHbvExvXG6wTsMmPmsrKVKJBC6QRZoIusTuzS1VpgHNpGOdUF
xQgRnMTGg/5Tlw2JyzalIVxMGC+DAFGtcLKosSdbylNWDJn2CsVvdXNBy9k5ku3Q
kD/tMu9cRIaO7mehIF3OgiTe6t1e/5a0/AIVnePOBnvs/PjAY3886xhXRjs/8gGO
F9oRG9mhDKscQou9cS6aqnU3HrAL2CfAXzRerZAl1vPWUT367axIq3jmmK2uyQMA
ASt7/rcFlzqHxT9ZQLgbZNkge+iCGxqUjR8GjjOAn+eRurjjmx6XdnSt0jU0Go83
y9uoFyb9dmI/vCLIQ7uEEt66yqTRIQO0fBAChlaqpGQcsZOcEguSeUsuYfq3t4aS
HCgzSIxXnaXgrJGMDmoUP1mMtn5V/b0oAAmLYiyVnlctvyTv68DrOl4PnzAU/Pt9
Adax1yJzleXRudMChtvsXsDHcXb40BfD2DZHacs3rI4iHF/UEDckm3bdyZJfZ1Di
C0IRm/RWjB29G+yTgDZOM1XpZml8VCr3ROZdJ5gOKSTpFBSbVhMOnrhmFJ6vChFB
aksuonzCAg8lj9LEHdTxnaKVzhcqojXUvIjH5ED6l8m91FLuQ2g9VacgzUj3u3ad
mLL89TWcLRz+qDWoXzC2Fox3wzjYLpBzVUywZ40HX02tQf3elhR0N5iE5nKNj4Y7
ymjAjRQjgMbXteoQj5mUS+sl1OypyWRpoyR1n0LACyTP086olrVtCviD5nMcMwJ8
4awIAJ6Wti6STxGr2bxN6JVtjsHC6lBjKRyi189G5oY8Owe4qFYEh/UxP4A/I1Nx
hv6sx52T7eYHk9LL8gqDIjxUS9LnMq4zE6t3p9dgbfPryITNYGE0eb6nESvCARUa
1JJRHqKr1zZVVaVzr6bunYAN1Wzz7h7iTW7C4ir4EQPIjhmZOu0oSxq3oENmi2qa
so+9dO3sryTL+zvr8IWZMgIX6kNLVFNJzXKnW82cQVPDkWUlBZVaqYv/NjnAnk9y
SUX7jdcot9hiO0gJ1+ZmuTi9nh1O6wuNoJ/21D/EIim4aoRF3V7cB5V/GdKLJePx
50/eudjPWhHy3Bdjcy9Qe9TwIKQUpORGLVANTv765cS8Qc9fKZWHnsDPNrUFqgem
qi7iVWhp0VTc1oneMzq5ro1FTVi70mixtXss88McoVw/hiCRofbHjlaShJ3/Pi3/
pQX84uIhL4BLtpdrDIlwyhcBi1XO3V6hvnVdKrrzgFkb+Zt+N/odE0IozwM0+pwY
rxdY2tgI+CNkED1lo5KOhLaA5hjZbsNGVuCxQ332HnMR8CB9+s+a1dmwlZmPJkie
1RiO+5EXF7DN1SXYIuED44f3sARtvoe8R/kqjKaG4IBuf3NgYEbwZ4TmybtViF3u
K5XSk3A8yRfMANIOcOShDbNm5fRbl2vM7rtSBomsfmA0bABaV57OVclRdbdfhK2H
JbgplcWHwgLbU7zAmFOQ+p7/SYoo+eGeXtu78pI3UXCQVxs+UFbQlSs9EnF5aqg/
I/oo3oXwjnhvBxjpUoOixL7VOxTSp/HoJeliWFyg+7uj3TIUdtcSutcL8uZ9d2sU
/lNPL9rQkdX0Ol5PJ3GJ/CSMp+8GIR9y8yOZ2A4+8ZqF8qSjPTkhgP5APjv033W4
bqJs1RDqmTcVlir46BXvsG4gOcAUvW0xtDjSDRUUA5O1dOjxax3QsCEFEIMKGFrM
IP7DxbOj0sYOc5cQH0ZGjg0iJLamNOeZMtNRF+oXmfTUoIDOXk1lgTY/kjvLzq3C
SetmoAOxa1PkvKV8W3pGqeDGvjk3LdBzptC6+wssbzWvmPlyoAcyIMcXtdjmRweE
xw6DADnI5bbpNSgz5YY7JnIXuKFzwe/osOKI9Q/HdQ52mSxu93SxsdU+eH0o9PCA
PbLkJOjoP/seklvBoR/fJ+onFQJer5o4w7KlCQ/Cl/LJN79DdintUBYFG8vXUvCD
+EWzqvjVDU0mPari3GHlbl9hdrr38+Hih8+fGPJYBbQ3Gv5VGMw2cjK3KU1NZZH1
inrDbev5gjgnOYP7TtIcGCtUXowqd2Qh+Et4RA4tSjibT9DIfs8GfDMC2cSCqubV
7ucnGNcwQn3lC5XQkfhnRCMBHhJnjCm5KxMF/iTVyVmMjRQuHHY1sWQH6RvzFDTZ
9aREBoKbnCgdOl5WiSN+tVvVZ4baA6dtRXjalNXUIatXmYC5Swad5xYY5JBC+TUA
FzJTQ4nmRCh+dHjcmKdJxXHpptlnMeL8UxCDs4LGvpTPcgDAMgfURPedVih+QH3f
EFKecTkSHq6Gkl7pMiSsY1UhdFYw7uaxHHuX3zb86ujJi8dA124irKLZcSQ0b5sI
/lhzNc5TOQVPKy7BCw+J+QDbOnx6UBL1V7m6gWPiLIMhh4ExKpmXfnhML5erkkS8
dpLgd2/T659CUdZJUz+Bvr5U0wlLSUlq84XZ4IAEXiAf5imxwVa40r8bF54iPjqI
Nmekuof/keE045K8UxeBQ73V1iGHq/jDBmlnO/BpUecTJeJ4kW02qSeSF06AfVqC
UC2xHfxgPQGjSd+CmQZv99zoHiwdhuKAnhOZDSPQKqlibubKjv8zQTDvEZEf5rGX
4cdCdUvQgvayGJ9++Kbtso+hZwKuXE2jMe47bK5d4JbAW5PbgAuuvlbJZlNVGEiX
dmINSeEHIhLbc+uJ/Y8aXWF2NIfNozHpb+2m6hXIIHFzqokwwOTisBwwq7j/h150
+eHGWoajz/gUQZUFm3cLclAnEFdjCdgBpCG6iq799p+3DfOeAGr66aVAFrqyUuz3
ry4mdNORQNzw/F2mpG308C4OBFV/+54B01a3Zh849d5FTm2EpZrFe3bEO6Cx1xx2
0PCqwpn3UAGpqSSehQizn6EyAnxs2euyAiIxpva4pmGVQIlyiinXlFaquQ7rPpoE
SJpQf6mHjnpl+g1g+WrgkoNTYPTGYYKOP79kVrTyOlu82eKC1UrKa7Lj5g+yI6wS
zZpAjxokD+JsQucRJZqDsDe3QW3Q3Znj6Iou55SbROrrHIewoR4/Y9H7BEz4EPKt
KQdHLkP9e8pBxuoGAijahSViDZ1PJP7S0sWW9eq0Z8vRwNl76znCZiSHEtE1iC0w
yUJTcwoXrPh2iULVBteFKjCP5i62YdE0gkkNns6nB5H2U4e68PhR4Uz12VLka/BP
cLDPLT82c801k0PjAhusMsNeqFcVgKM2xcs1FFS6f5/+aTeJ6yGTE5UfpYSgxb6x
SW+D5ns0fgJ4Wk6sBFYz13eqDeP0fK14aHEjmBwcJn7kUV4tJRudCHMOWJcfYGBx
vRrd7HTDI6fWFzZk760BVlru7jkw0y0NRb0fFTT1tdUcUxH+BJoZqDii4ArZvCAk
jcqfdybxc8I0+9BzVLMQ/Yol1NYW5qdS1oXJ7cEsBKbNhgB8M5jOkgqJf/QDeJJw
RpTATaHi33A5B/048G1As51QErAVuQ41/WP6VDKILgUJ3I5CSSLcr6FzcE3b56eo
DLJM/hGIHJteLGW0zmafFuNgfh7JK0dX+jSj/NC6IAbjLNE1S/4lVGgS2YH2gsy3
/3MF3bQGF91KkNU1n09LEi+h25Hwe8I3ovlAvUPQtKhuAoAUbZHINNTi9yDPzrUB
SNVdb4GrzmIIoPPrHrK+S0GEVyMthbiOUgLTtcf0fYjHsuf4fQCxtQz8U0ixQ84d
x3vSochExQvey+vOKaUpipeGn0DJcbx2OLYgwEefseDYCrmyOCpD+dlk20LeSSlA
1/Db+0y14UoP+nTgheVw0Wqt5BvTFMhIee2SCl3L42kvgnyMA45OqxMk0VrEEQdW
SkO3+as3v4NZO/ure1g0NNoak9O7v1+OpIdmpXSZNF1wn6s1q1U3j34nB6yGz8BD
YxbWJkIsTcPdNHq6JvMEVnOGJcimwB+Zq2//6cl8gcLtBLM1JLk7xKqcDppiZ3IQ
2NVAbZ1TlFwM67QZVfu1DCo1evs8k+xqY6aQrY6WoLQPHQ5Ucz3WniomezXObztl
srtfke2pAikKPmVtEAunOTR8WtH8LFJf5NK2/a2POmuUKhtXzax28V8jTspiluYa
CtOYYWFCFgZ3bfQwEaJ0mJUNGGGdwrg7T//gd5ejCU1xTKkc9vKbYi6/7yaZxImi
3wprIrjt18xpXTr/Y4OMDUskTsrJXl4tHS3FMnxM/L+tU5+ygQ8tsOswUZjv1Ewc
Vuy0VSzoNGx7gHuIsr6jNsyXYD+seUDH3sQfs6eXrL1z8Kox31MMs+EDsRQv8VWM
Gl4q4jAMXJEo39ve2hRJMP2mUIjBUIbli3biZhioQP2p+TC6EyXiHPMzyNUFQFG9
8UUMf+ZEN5xn0g5DIB+83ruXZ2bIdlKnZ0eswGTWcLOPqqgaBbAoLdNh8tMNtaYm
DlznsavlgElSMvhCNpbtckDPIJsB+9hWLIWxy2hkEFJmIxnOpdeKuiU9E0833Frg
U4FpB6ERh+h4MEgsfpuTnTnzlf/0H1Qnt4B7p0pb1cTzkEhmJngO2wJmydSTfHIT
2w+X88T1wwyHbGH/rrF+BlxTG1rYWuTwP03aSf/W9e6l5K5t7+QwtkMR3tlHLUcC
qwKrTok5xRqadFxJ9iOqx/2bUMshhbsASbeDk1/3wVisO7yi69/eYlRxliZMi9ex
jBSRrLLN6O9e2MjqWu3XPjvQ8RYSM21JAS+jsrcxCBSACEw/VNeUdAjqmGpXo3QC
Cajrx7JAoTKjePtMRGgY9huB4al1C/BzG90+DemICEpSfkG1GYuYZZ5RvXcWFA5u
/dSOLXVXE0kcYFjHmRnqEc5MsuciD6B3QZQhz7o2nAJvDFahPQvmtF2MdVxNK1tU
w7RqPl632+q/goTrM6vMoVnD2rFPc36P46D/3G3NxhIpHj4TLj90C/i5k9eeCAwS
i1OIk5jPHSjxtVp0e8sx0k0zVUqSYlx+CmZBwWEUQzZ6ioLoT8lWTv1jofUkBK0w
vWII+21PHS030eq3+EGDBIlASA3H/ESon57my8s9r2qUk/mrcDBUOFBNHIIjBUd1
5lwHrZI7nkHGiB2+qTt9Z1qvdrT4zkeknAsLoRaZmOugyb2zfnX8x/DjGqdjpVTs
vxmKmTQvm00xSDuQ7isS0XAk4Jsjr0VKLpZUWM+uAC4XBw3QuoXe0bJdeZTuBxCm
2JOR49xZynadEsKCXjzruP2P69aWjp2PGtPuZiK9E2DfJtOHdvvNZkrTmwk5RdHV
7vZCoCw2/U1ItQrDH9W1PyaH7YY/yZvJV48cNxfI34owjXtBLqptBAsyV2MvCUlG
pZWBVNJmSVvy6/HgqaEnS3sa2c6SUlJuHM/nNmwKe2PS1pGrbfXEYPPanO++BUTA
yUAlT4Tt/8BMnTrqkphJEksMsUr326aIQboeheZCdrBEIZjizPhcKdj2fkH2YZs9
DOiD2PmlQ9XchrPOh71wkdFjBdaVBU/JQvzVWccg8PQEKCYAfoKqeumsrVacfPZf
SCGYtNBZAo6yuBKD6ErF4ouLH9kOYMqVSSaO3ZqmbcM4IYX39c4wYKj1wNqpJvQT
++pnKMEnpjk2AvguvPKjEl2lpb2vvIk4LMusavtxJsd1O9ACJ/L7XACL3tKK0NZR
QMXfgSvjldKpMlNGNJR9Vq+VOk8cwDnGVSlBHVbQs6eqprxElFIE9X/mVfTP8wyV
9xDyzAVP+Td6vDuAjzeQ4Mp7lAG0tqawdYfnK7AcLWjekzdnYTY5s63sZnHDlOIt
U7ZXTg3k7mW2RTdiZ+7fkyQJXk6jWlLuZ7ioCCw+TaFDXb8sthSEECJsxu8glfYu
c87/Z9HXiKL0Hi4wyh1o/AMdVwBbOaKYrwgti6qEwLqqIHngW3uEYFLbwjbhKWqh
4ncvcikR7UT5SnyhpLxD3Y7YiDx8BZRXWnhV44I/zAAYhwyN06XZfqXdQ9On1K/h
2v9BHmlLCNNmJANcgnYj+zaNpfu5II18QSurkYoulH5yeYTjOSAFv08vo36ZNgYS
sWIs89mEOWQ2ZSA8d1mh9fi0vlKy+XXB2aScDKqMYbl4yNb7x7RiQ+nEPSnyG7pV
x31AIkfNoxrcDajmiXSBgFNGU3cMSxaYMd8072qicjvMTJap/fM0Rlibm3CdlSi/
x5LY6uvBACNtCOk059na+2uMDySBeNFsRsOO7gWgLgubyJP5UehlnZOhpVxNOyaa
xCjx30AH0lJ1jTWLu0OmE9OiLcnGVwnCEugmHcIT19+InoLbRLEyfrp6x7tNyMZV
iNjhS5RxqXUXUI8X4kvYfvQS+/GRgILHI/DVDpvANbNENdtpjzPkWkqPAW49tS+k
eY6l9tz9gFJJICtnbTDHenwFF/uBQXAqHp6OZqaMyAgv4M+xPHf0DGYhPxf4Z+C5
rRYq46VlE+7YB26G1oiHhB+kvu8GOG4EonWUU3hgxnu+x3NDSVBJx7FoV3A4snbL
2AIxhxU9ThIGYU+cKoHf++eDPM6JH21vISgcAqpQEAs21YhbrpKQjVpYb36pzYa5
Jby9TZHpGx+mhotgY3EfwnbDz7uFgaqciFEHLJyMygGSBsfR5YPWWAvvXJx/vqtG
xt9E8K6hKiiKUxQBvg6LeQumksJEkNc4MyOjhbi7Pm4juAowZk1Z6FmRipIs9J+h
dSqcx7qnabFScBOyAI/l+0dJJI05WQ+iyw/Laxk6m8SWncrh7415RT5lT6yUY2cz
rhyL6XJGLarx5fahQoIbJM4LMYBfIG7EK+h7DcKX9MQmKpPMmIPMVc0LJ7WN59IF
sv1R2NKYJ0niHlOx3rNzBMyyCChA86UKAPkAJb/fi996YcHGsoOUY2806IlELPR7
MCdd54iaj+6rNg49wVFFIo18k78o9UxVUgg3BZCBHrvoGNJwC4S127DMbwgMyhIB
FNYb41+TBypjnHyc9Tizyw==

`pragma protect end_protected
