// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
2OsTS7f89ahIcYd3W4YRA+BBK3NVppgF80PpKp+OIDKrK43+2KwxjxQ/jlCQliUA
FhZSmgiozYJJ/bcN+gPxMd32PvSdR5H2BvQSgLgDHAPl2As5wliLbnMKnf5bOL2S
67aeL8/3Q3KWQB8UsOer9DNtyLdgqHDXjHBgBJShIHbvqWVi6PXoOQ==
//pragma protect end_key_block
//pragma protect digest_block
GlyZbdRvAgaGph7Zh2teb3i2F5A=
//pragma protect end_digest_block
//pragma protect data_block
8W+ohBEWr+ohFC5Ou0igvLr4DzcmNCpF1jrQS6JlF6LEaZHYGjQAGD+h+TDK1XAn
dIh/9lUu0nnMQO3T2lxv5tNpt7Il+oOROu/Zzkh5vhaJV2oZMiM8aOalkypIRBsB
U9/OlKaMlUkE+9WpY3Ib9j7camRVH8SwPbNq9hrNFqWpODxzgFZQxpyggi8VoUAO
rdU6LXviPrC2AuzFFPqFNXj7x354IbcXGl0sTHYT7+JHpGCp6TRKxNlI1yedIbe+
xpTXgWRlC8pGA4n/R7r3hOXFePRU8jbEYnb1djtT8IaF8igDvadYiSQKdIFWQ1G4
0da5XE8LT+dK6qkDg+t7c13LRlw4Js+G87JE9sD/CWVLOMg99HX/7wO8hNWq/A65
zVOx2NzcQ5CQdXrGzUwazTlygngE8/toDAh1O3KXNvZRN32O2wK/bMSzP1vUyt/1
UHT0m4yqJXdOt9i7Yojkrpp15BH1y/8KiPUFelPPoJ8vOJlMxOxIAC4OevTY+bHZ
xZ1fBybShSG/lk3TKDHvj9m3+Y6RDm2wnnS4u65WeY+tkid09ak94lvpFfejGpn8
0RaHnFb9Q/L80T69AA/vw7LpZmLZSm2W10Q9eYDbTtQNpWY5yluqE0f7/ntrJaoP
fZcibaZt+JKU+bH09cY6EnF4fIbFugTPetVggrAQ8D+aGaoRKMyNshMM+c727+I5
OqW5x7KTBolukqXLD4hL94SUYCTgM5z5u7ydQBXamOj2tcOIdhwTQ7/VpjLwUIzv
Ulcd1RhrLwCgYcVXSJi5rrhIfqK3aq+9lMtUeN8wY3I/CZwHeEa3hPPYgvJoYOC5
QFrwlGyxHmebaiGAiGJHo3ZLIJoBPt7woWEJCeq66gd9VZfqKdbwEFI2jn6dOihZ
QlqMjoKc+MSiIkWuSQYGAHzftlRqvvlj089lD8LIfmbgjyVic0YxzDqa1gvbJjEO
9drL2enuJ5EJdu+q1cgDUdgohbFxCWgzlBtcYHBujqIQexMLna8aKUT7K8lFp2iP
SZOlQjyleQdEc+iwVsMB8rM/RLfPYDavuIQKUbz1pe9d1f4w/7elr55OFhyns5C6
WkoGfhqms7GuKnYy0oukwcIKCzlG+RBt/AWH2S1AlRZ+YUp0V+sK9R3T3fImiWGp
c5xrpxDmqZJA1jNl22DfDna+vJhOzV83LzRyZ5ThleHpqd3LnRGpp27XAdcRwfZ4
a2c5MiGtBmCQaGqKr8iXO7rxJ5mMZhA2KZRQ1jzg5Hv8NalKT4uKOZjX22XfD9bX
Pf/AacuuqxdwyqtxS+5vaGDb1uKPvNznF4FE0IDlM7e5AZAV+Jbw6UQenjv1HjcU
bAxZwxAZ8RfUeKGJcCqjyBeYqdjD2rWUjb6mjkLbrjM4vNgZNx8uVVERwiUu2Jjj
GBXmDJ2t3E8Me9b4ZuKvGRuLR+c5iQom7XGVa598vu/8VbtRABTHTpYRlUaJwNQT
WJVmwRv2JGLMfU995daZxaKOU7S3xQ/v8klnMxtqFHsVb7II82C6euepvtxkv7iH
uATgkZtpjdC1vvFeHmFLllc1DRggXyJosFWoIxhVOdAIuJPsPKmzGV2NIRVdWXNF
PXgZa30Pj5U2j3CZaobmGH96sIKPpCo79+0yonslF7XGN8PN7S4tTKayp7s0Yiry
cw1RvGUcH0R04+swddVlfaUBLjitdvrnYMn0ITUEZC/NKdwoxHIkObq0WFz3cnd2
Yri0P56XCgdBYC/DNikNK3LD8/h3AdyDb4kQFS2o9Op4mnCXlfxic5QllvXB/N5p
Vk1V6YDl64AoAbVnFxjHY+2pTf0ZEIQq043KHl5p7IsMCacy2fy1VLazHZF4zDcQ
2fau4vK+KavhRQiQ8XvtwYx7yueTQBaH1j22Mk8JAjwbRxkU4wMFJmFDrLlU1fIN
fU+heXJDbHSRZnDciCSwIYIEC33lZdXk7V0yohuAozcAHdbKWP/OExUWYg1cekxk
yE3BzJuiOy9N77GV1z7EThVqeMmGJYPSlzZuqgXhfAmIwFXIcD/kPmXUvovvOxjs
VoKu6wABJI+krM/clwojoa5kdkJvnr04MnQ72+CqyGtgYmXPC7SpiOI60CfseZGd
DN8TiSLtjxtMOSkJGBZdUhV9RmT62rF+lkNlDHRwy4UR/VEYezxH62jb7rZrAifY
k40zb1B3LcDbp7NZjP9vUAtuTYixMAVOkeYMCnPtTu03S+fj+tVGmioHLxRbhVWv
JjpnpH5n1GWhkKxd5H/yRbY3lWmFsQaunguENpptaiYV8jmkb8cx0CwnMf1Ez+o0
2/H7IG6zsm/exA+jNKufpcDWuQb0awm860BrtBj2pD0r1TX5g33nUUPxqkfdA07J
qVno1BTlOse05FRF3TGtLq3Z7hNQTfv51DCbqFAgNtrBxVl+16/JbzgohvoBSHpn
caoEcpuo72zW0uHUfSG3SGs4mH41iDnhXBGRF0hUksd7KuxAwSQtFezT+Z/jdNZd
P6mIIk2MPF4+Scbkyd3jX+xSVGlCDaCSZ5Cstxy9Ro7LMM1xvuPGfOuNfmusxX7Z
pb+RxAc0GINMAtXKcvqtX84OXMMkxjIkVIerCs31268EMVXOh17sejwIWj/FeuWU
vYhDYu3yu2wK9LftqCovHN+r5nH1skDfzy5WGCT4ZioDFT5jZbAQzi03cT0XPjuS
Bj86IXgJiipr8GWB+qzfR2ro0vWPbMeb6rM9ZVsROc8EeC70ftq1fSCDvHbgp4ZD
RjntBBlT1l67K0ovXvSFSvzPDN/0OCzwT4ZmZJWhS6+fe3gIdAJCKlz15Gv/6WAU
CP+k6K+MQ5I4pPi9lLNRZyUrCKcXS9roOZaMnXgsRTsWOtfZpG7T6r3gy1RWrN7f
NoKC0V4uznt4Gws0t1jzdmXH/tsCHE4XvPfuQ/1kRkW3Pw88yqHOkXr4AmATd6Om
1SHFe7QmgGQdFQdac+OSMgN3SrbB6mmwHFZH6OjRW9Yx7F7wuhEtZTIIUWk6oFf6
P1c2OB5dTzlI5d5DFXtNbOpwMHF4xth7JlE1FHqEo++nSN0a5yeWzwuIVuz41ryC
3BQOpcwPzLg9JmVmBzNT/iaFf54y83PlSNxfMi9RQZ2lnSzubGTAqR0IqE4KNmhh
Sv71ubUUZopWb0ZJJeH46wvuFniNs+XmiAiNPNAa2o1Z4VPjUpIEyIcuUTP9JGQy
nPPr9ox7zxUlMgKmo/PfWJ6HC4ntlfvxDAZEGENcxUuBpJ9tc/ms7VMdg+BDUDp6
uk+YcZZQNyqMLksfz+v9S//fDOsNZUNqYhH2tkWJRSvqxdyhV1lRFjRD4iRR7XWJ
H5kIK0sPI0uqjNt/8jMXfpAFnU4j5Uvh5jQsrVKfoC8a2InQ8LJDbJVWYAYty3K+
5dg55ZUnxNjrs55KnX0UELxwnllRjQCwy3LdWtY25spyzKYV5L2TLlq6357rzVyw
TFswyzSnVTfdps8x8pJ+HqpnAbQqWBJ2hQ9ketYwVTtlCJ1NJ77NbPO8hVYip+qk
pMXyhSEDn8n1bLDugsvu0LablAhH6ZoTkYPXn0WtcGEGoLwyWTx0593k0foYdB62
9MV8FhYE3OKqDeDlAdmuFM9IePpDpn8POFSaisq0T2S/RG4FSTe1csughFAiBXUK
36X7zdbG8YQS3GJCkHLOp5AkoUtH0J0TyIDMtVlGnqfVkADzFikBNMxWcEOmr9Z2
QbDABTORPYmftTtdBicsMt4uAIrrxgqvonXW8KZPRf4ga0T5XK7WzjgybQfTkzq5
24N/aPKB7u4gzDxeKQ6rP+g/2mAmEGSKfK76BTL32aAVSLwJNnvb0/XsA+pyERZ3
dOSOC47UDk+NZJ3MyzfD355sPCiVxWKJClqoUcQ2B+Hz5gMCKB3DaoSzxoGwJyfe
stC+pUiZyE3+rkjt2AUxHGa2v/q5yjFSKXwCTgk8vr8/MjBG++4JwBMQrMUKe9ZU
w63Et9pIjxC8uWzEp7oBCpcQ6HNDNzQcrdks1AmZ5r8v8ViujUnEmtlMc6XYD7aB
90o+TQWTOVx/EFXgbrarN6qP9m0pnDxdCOEcWdDPu3nAEPJQVtywxNRhdskknkuY
lAaMuRHwM67G2CJqA9pxxh9rF5yGHmlRAYoMYkP6bZHox0NwjLMasC2idV/Sgpey
ZVyBA7FJkqVJMcxP3v5DRFuOTEbFeOttKSyK5om5ICstpOvEPfGRLi7aM2EndNGX
/z93bdgWLwT3Gja2s4+I+AmLCQkiNJIwCEkGzTa5enJbNjdwbpUIp8zsAxEr+rSw
Wn0GDr7ort1nnJh0AifEsXZe6eRbqTeoVja5qjGji3DmbtLSdndm1IMY3a3jNrdP
0M2vknZ/mKMi0YdT5VakhG8w/u3AJeidM4AjPpXNA5qh476cNib9L9Yvbv1ZqPv0
MtpOUjBg1zlpFDemNLlMm3o59/sfaqvdg8xkZYPz0XMiYqxZBx5LZzSwQqWDw3ZQ
rXmKmK69DCO60el3gnYjJ7VaTuNWRAi/LH7O6HAQ4CT8Y9IdKwSVVB6JEHA4X06r
qXeLW0pqEQKVuDpWtzZtyB4wRD9B0yV51w5JrSx/t58E8yfOMURCVdbpsF6/vZgS
7iByZssoi90u77jWI0V/gwTtzKWZfbkDQRVrB11cutzmZYcnV3U1WTyRgb2eTjQF
mBToQVxzCXlcBMJAs06unP28zSwOHZRI7CkEGG45HTAVlYaTtmkp/wPTOGI9Qz2G
FtDJfjgYLyxlVs1BYi8pTr8ATd/gZU5n8Buv0dwwlLCKH1c7XqxpAaUNGs+cfeHJ
OUITjZthJAUD+2J3U3E26ecoEFw5edtA90RfBALgK8fFiKLU5BxQdpGx6kRDQweY
8oYYIrqXM5au8repngBxMslClH63t3urgD5NiynZEl/Zm12H1xwk6R4rIm9z+BzJ
fBvzKYkmxvOkl8r+d59pTkTxTQBDN2wuWhPfeRJs1oXCwoWhKNSfhI7++r3BgI1A
rFHgK2aXJ8LGi9GcseqxFbnptsn3UuBTt3Z3N8qKUVYtEvh10aK1dR+LtYIF4pzI
h9lyRv/Wm1Zo8IIJjgQYHBBcgP7X9pfGwJrJPlBWxMIBR0w8SXH+ZD+zuDRZaoqK
TOdfQqBzv8uCmr+1YkP6l+mBkck3n29OQuB2iZpVo94O2iWyyJp8y+AI0HQYUwRx
dAuYwFIOFted0f0NeNXN2WoXfsD3Y6HTPYBpfe5qMvm7Ts8/OBV5R77atGOuNEZy
FK+j2v4hYfzKgY8gG9pTghgj1YQRV11Dbo4V29O4mVF2JLoCnXM6X1oxe8XG+vjI
bz45J7DtkeyKr3H3jQ9jO7bPGK2ZekR+T61A9LmVtWyc8u4OEjawVYYH02vbof0O
cBdUBrw9ZbxgxS0NZL8WwETe8iwE4PcI+SKHT/DpaupO5G05o3Rr3GkcXRN93JJA
Dzxef5YmwlHDsQXGn9sOM/UCI2VCDWB7BmS0BRjcRHh0rw8PbvNKIU34g4sm5dsG
OLnaNyenV3jHVa501l6mPT0oAJ9zeyAjHn0sX1c7yp35V9423tayRkGUD8hBxrKs
UJGSscOk3tuW7OyPGt8uCi3RSDRbh+t8nZ3IHPTK1RxlFZ/riSnvd/rhCtqu8JfZ
3WTnLw8WDNhxgeLwesTzIweaYrDz3h8o67hF/foXX5Lo0XBmH3cXjkmIYyNNrtgM
hdm3k9EyZe/fpYXsx9t6llQDCwG8wBCVvXBtTs+9gtzDBgcKY4mOj6+zqMvTUNr+
908D5axEEBDW56A4/bW9q5WsVvMlHaadTD0tJkl0oXMx9izJqod8S6lU6gmvlo/h
ajkbELZvVKcHwXZ0YE20nw5MWChPrOmmV+W8g9xbKoGk/gWvXjwlMb2VvsAyUHPB
plJADRmnv7XIiku3CpnJgIdsh+HkyeufEfmqBtxXsAPu8dtKc2wdV1Sd1fjz5ACu
2ODmJK/24L1v80c6lb1zL4euEpi6xqoeTN9x+RWjtc6zoQ9P7++CjpSzDXU6hFvW
biUM3haZTb0c0dtEu8mrwbad17b8SfoaEiCm3S9njGwI8QWzJ5buslJfDCuwpaAE
BMRLODv+KJ/E7kBdOn3BewA5i+zBpXdXBOnTs3o18S6U2DPFi36rKtFMlB/k5mPl
ZCKmi3RUFBZHKuGe9KzpYBWFx7C/Ysu/dfkedvvwPbV3QM+cha3TWrFFbne8tpvD
SXSZtB3jpFMcbPBs9BUyUxlaIGxceYspxhmwYJ+CdynRlvAhHyQTn7aFyZX8Y6sd
qxk8wpwtxX9Q/eFq7Et8tjBGWkIAnH6MM6UhLWZAuhSs+qRUw+5jzRRCr2RqB1iR
Ynw9UzyuP1Cm4DcQ4HdcptvTh6j3GAiIU+2W1dTldIFBC/HhUifZl6xaF85m9R0R
9huuY+7eIo92VEtri2F1rQYUZCTNVmNzFf4jik74lbEIOHYiisFVfJdZTMSaSBih
xcrVhLcXnJutvpdjhhHgVVDnZ4EI0h72J+HSuWAQ65xS4N1VBgjKrvQGWtF+qNIe
LiawtISFc3yFT16aq4XsaHZU1HLjkJW/zHFNlA5ch+pR3FGfyurcvalrLBbhvuIb
+zg2zgq9aEPdajJFEdgdSdJs3IvPkxeN7V+Lf2OpjR0897b/2drJCKX3f6V5JgB1
XRreQ3f8oay6syt78Dy2n+aTlZVx8CojphyAMTG1wLJiNZzi2XWI6n1ojbDvdNTX
yeEVPn5Fdl2hFXAVL8t0ej6ChMoFxHh38FxY5aKXOvBxd3FB/p5o4V41laqaPX7J
Bu2n/v+YdG/Kscic1aFeepGJ4X+wgY9PjPmt8rE/o1TNFFkkK7KwHAeEPTEhlLYh
XDFBlb6apGvZ2SlV/2IpbpHSASCnyBPGRtQwpwog3UkbHZmYd2mrkA8E7NmZYuYB
Q4mP11UBLpNU2wPl/V3u3l+wHU7AKRVZvoWgrFFJd717ORQm+oF4s2mzp/EU8pBP
p2P5a+sZFfouNWw0qiS1R+L70ay0wXNx2FIfRzJ/WVPnUKvTjEHGTVBf7uMIxljJ
O3T31isi2IALCdyLWbLsYE0893KRktzGVsKfMtNBzWjvRgZZZ2l/b5HQtGCCeYp6
m7EkAr26GLL8ICsuUr21guaWExigbzvNfiavSG7fHtrfFcj3iMo8YG9v7D6v91o8
hz6583tZ7YRjgp6r+mTcQJbCdc3I60Kky/QygaWBDvxFBjAZQm+LN9pmnjyhI41M
huF+HqmEVVwYw35vQRx1ivyxjNELJ2xgHlQaUeQvxYslGrP9falho0hQWI+jAf3W
J6LWFwSVQron8CVzdC9GKEYzn1ReGqbHHzr7UgMRRecBtV8eKHcS0J6j87v0D3wf
Na732hR8OFCb5m4zK26T8zsvFHMY2qU9nn/SBI0PUWMGAiv8sTdDlB66zuFTEGpw
3i18k9ETLNq4z10ksC/VD2I8Tjl1dpO1uZtlkDAiECaxt/Hsmqe9UZLfEBCh0WlF
EKDd3MCz+6EsVp/Mgh8zLyCg1bm4lwCzKOHb/inRxo7lZsJa72Z0jSbCFXQojcnV
eYwJYIEegd5BIxZVeLWDOG3NQciwt2/XmpUhu1e9xoVLBjVu+vsfOXJ/Gli1fDN+
pcc7zs3G9VBaGwrCfGEwXNROi6qGjHSYOZLkvc8erQF4qGlxn/H4a1gPkMrqASu/
ifwPCCUq/tdbPWH77AONkAnMvRQ2sQw34K3grSPAK0NNmm34lDYB/+Vwg4E+DdtC
XIDnkEIX5iGrYMrIVQtINrImYutAKIj+JscTJphKVlnT7xPlo60rYC7vYyPDUL57
sXLEHdseWlDG45y9Not3OZop8zT5+Xrp+kgWi7M7VwWyjrjVw5eoz1ZTbpVn1t8a
dMpB4Mz0UTQ+15zv9/D1RSYjbTsB4Wg8jnz1Gz8Q/OZyxw6IhXQ0PU9M8LLJX7PH
N66POjlF1aOeGE9uugEh9PV23tOhkiBqFogymTn591ZRKcYzNVcSPINrYWrNONR6
IJY8v93q+3YsIcDT94041cRg4x6dpZFuSvDD+yNyR7yBPfXNCxCZyES2sssAujbT
p531yF6v5CX4PjoU/T7WW5iJcSYpnVsF6slUjP0DFEDZ4nAjE+tD7BPOU6wFCJwV
qo8qBagFyM1VYBZWsAUeOzQk7jQ7UclL0bcY69R1L+pzYzMJ67wGNrxouLifW/kg
WWG/DgPpxrrRAvz5BNFGTxBTGobFwqTE6IbEU3J37lC12opFiKxTrq4uLAxHDAPJ
R+rVprbPucN5J4NKuy5poONxuohRq2OkYZSvsNGRwk4+5AoIuaX/t6UyZTQH24eT
If4WNE1Jq/0gsHNPIyKESUd7oZGVpiHE6Rso9M2/aEcWyEb1ll8L5FjyAY/N3YKs
QpZ+zK1e2/USdDX0meolnPfKfMM0uf+Qj9mm5aa0MCDlL8tsCjodNnNN8C7yN3JO
Z3e4z1nVD/WLe50UkrQfltD5AVpOynKNHvAN6LlC8prsBNRaIZ1D3U4uG0CSr/Az
myeg5/ZmrF46hKI9mVzF4wbdWHGqfvImSX+qLnzIqU2/d11AvfP5XuYB5ETeJsEc
2l98cgX6Lg50rs3RkSNT1J9Uzrm2wYBS5wttPjvlBKDBNjioGwspuEEFhzkukCPA
zRQzH0AINrj3KfxAHuO3pE45v7RV4je/I8ffyKj6lklPOhf5MYepmx6Q22lrQPOk
pOqa6Rm0ZAM8hm8ORDfc0thxIjvAmfU5HaqG998IXaFBKYaU1NEXqoPZ5tpotS61
B9bNc3D1op2cXR1t10xskssh95vTXjTdJWAN7o6Q4goMNmmPzlIVTzMpEXGPy6eZ
W3ReT7hYxHzLnF4L4RQ3PJ9Btd7DazHThBNNUivztFUsibYjlGfn0AT91h3Q7LAB
Jc2SVBDrpXrzPYYTnA++X6NLDG8T8EPs+zb2fpYiZeeHogkBQJrhvrBmgQJMvkna
Lbd6ulpvDy+tNQkErDRgbhLd7FDvbpwgc6Vrx+u4eDlkC3hDupmtcy1CHfrKuUVH
/IMEdMUQFuxlOzkcYE6lvW5E2UkvVPGu5ZF4CS+t7CgK/QNK6fjppLaMIrKX4sRT
rxFUyfHY8Ru/CKXToxnrRfUryIu08joEWn6cq+lw8E1IMx6f6LkLPIFKlVoM+zAt
WbN8MxMe7kz7vWW+kdFljZdTLqb6spefkWkd1lea5hdZ/U3xsdwUQ0IL6uiA6pro
wSbBaNOzpJsh1wonP3vh1wxgK+PirnGsd/t/lxUw5apv3bbVzEzxnQ8Pq0lnwKaU
+wlwvwRsfuD6pCqxNTTXJzJ9WFXl7fPkwysoQD2xg9bQ8VuqNC8hoLgBiMu5OTdd
NfMcQUafHeC/HaWGLDaKIHKZhg+a2ucRixa+xBQkb4UoyEwAciM1B360FHXLn47h
GXevV9c4hg3p++0Jc6GijSSVLSEl8eDjVhF+s/OIxIQ3cyoxbYJuvI9c4Zqu9g3J
x9sqUd0UaEBq+Rjw45dHw1A4oOHuQH6aVj1p4j+/7ZGNAOARkiIajoguzk+RtC/h
c40cqA2WBIdtUZze2n83nOmM/BNuX8Mlx9JeIXhenPBdfLB2qmeFl9qkhunFTGNI
AM/k3lqeHSH5sKy0X6JYg9z6iBu3lgrq4BrYVwRC+Pe1PptYs7dZb/jCd+WMYIKO
oGZ39Ix/INuvySKbUKQel1oeOLkW4pjm1r5jyE8QuUodkT0t/q4barYbcUGPqBiU
bXQmuPeuXDXvmiqnIwfCKAGCm+VWaPwUKLmvyTGo4Mv5X9d3xoWFiwwKebw8wTe5
o9iU/3CLmIpNOSwVZmOA0L12xH7Iv1X249rClyUfhF1ZMY4ys09KEgZ4+pEMEENi
k2ZG0k2xczF0he22B5ShaeDOVj7S/TsxIAKRg+iv/l2ZKs9Jbl/CqAMqna7fKJgc
Uplx2bmhG6FwKbApVMiVkYUN1lMsTFlA09FGfuLzLvK/+iAa3MqjzieXgTTIJgAZ
Wcj0tJdnUjs6BUJHtzX9CLiMozRGdZucBacKC4+S+rl9HmGxySz/gWPWlzsNTTW9
Sc4roaIAy+kKnwwBSZdk+wr97QOEisdahhkkHrGJtnMVmlwvuuKkVf3zjzB36kub
NZkQjJEbtqCDYKEUiKT1mfpwCphJTSb2k4xzEX2lNIjnR1M2GGA5D0azXbxsKD7s
+iPZ2PWoiCq380rTjEyCvErlt66X0BZH3wyJ3vhM1Y4Obg/4jEeAub42ikiEDgvo
r7CxKTJBdOPxH0DkMEddXorOgM5i2r9XtL1RIhdJKryynHYrdGJFqJh2wEzJUu1Z
ZWeBSti2uU3TlHuBz+oCt+02Tlv8mUzWiVLfTfpNCbK/j983fGSDbDLLvZfkX3C1
8qw6aeWuMD8x5qQAv9mq9zfrixmi6SLuGqc5DeLZ85tknhv60CGIJvGT6739oJoY
wTgvuARj/mdsgL0vqyRQrpZXoNnIvQ/Xa+vIxKxWyVgMSAF+T+ub0MRJhkpKvub5
zouQ82ymyvVPnZdhZbL+mNWmiDL8LBiZooqdXYzUNj8sMN1YwGGRLLNHvhmvmoOE
CsP7lfO5JIfhWLcUfi1JCPQ3celR/DFi6b8J8cszmDp+XyqmY0HRL+qTZww6o0bn
I9n74rtFUS8DOK9Be6BgE1sNgrpp7sPmgOwJd+2ClcxTYZlgvG1Yf3ZAEuINhslj
xcO0UD73vR5ZVje6yd20YrMfszuQCPzy7Fm70SPFVrMCY97qCYD5FlDJyWLzRHJ1
aL5SrNb93qQMOyg41gCpuYEYYRV8J/uPgTx8rTCQCG4dtb8M7wzO1AO8qY85n6gy
Hv2eNaeJbjuLrj+VIdULvw+c6xKmtZMCi6gb7iJdVSi3C1ZXUTdJ36dhNCK74nCw
nvLVkmad2tPuFPhWMy4/O45LvSbcPtWJHcM3LOBHHVEkl9KLOAPK0GqBNFdh+JZa
9aJyO44bQeoGXGgfD0SVja9scy/PdInaS4IKHV/xtBpPoFu2kAaNoormyP1jafcY
So99wlc3RPtdru1BD0y6BY4fCgmM0JHixYNLJqMjSe+bQUODvh6AxUzVu3PUHB7T
ps/IH3xVs6/7dkuUkgVcDQPd1eq09IRdzMzOWf5zOKrtj8TGlgrrn6gdkwzB72lO
9kqO3hYA+n3unljKGfuSp6oneysqFpJIhGfGLzs8qDDnl4utPhq6IZAKe6okZkCx
MaQJWNON7vFstMjtPyMeAhMzSbNhZO6UZyDOIEWLnRE9ZSlgV30Kmi7/mT625A4s
U22eJ47JPJxUtZ3c5r+mkjnafSARY4S8gxytVRxprAnKgfWfD0DIPxABV4QhbvOW
3LJ/7agQY5ygK5xo7EuZ0zpk0Vf+/FDw084Oio3dKhp5GN+eJN1G13bVh7Tn5qx9
M4sM5ZDZ8KYrNyed7MK2caDApg5bBfrgzdLxOBNvPemULgV61Zzpe3GQ8CEKJcxw
+IS7CFSFgi0ZXXJJEwyW3SOVaAK5DEa1J5YQQt4AuylCojW5qv1oUt6gka5gLKXE
CF2e7Vd4gg4xrv+GiXyvm8COdSd8C/uGOBifQLN6yfya16PbXuIkFg04PAr3DU9l
+bRTaTH4m2Nahc4Z6EqDX5uaYSACAexhaUUTFxHfxHfAEoREJm+0j56R0HA3xwTE
kngYQ9EHeXfVhQpgF/wbLuWS5qgrGCM7Q9Ebowb8UtWyvHLyPoiaBq3hi2mZRMLH
h4jun/IVd51Sd+10iM4li23Q8p9cr0HsK4hq9zOX4uGEPdb4nqeUhruDIRTFzRrO
P3QLAhpbf0FKHBdakFfOghQg8FdugyRd29VIIr8s4TlF97TBDEcNEq4ubqFZNoUB
8FunitZdfhAO1bVIq3totVQ6TeJrmUZv9HBjSS/J+sPugFBSMAAkHXWJk+5SYOru
hw3vexmNVK6EmiDoP/lE7M4W3ZLO4iaFtGqPcapjfI6RYHt3XLzauzT4iERzVH3N
AOskO57ib4I0FXc18Xbs3uMQGuXVNvoH3NjnA5b1J9j+ZswKKdmexLOKXNUP2KBR
SpW6zUlr9mooSWQB/An1RRNMfTs444G8kexA9TiBTUbychKwRC4ZcKNUNUMP2mg2
k8md3RhNuL2u0vfsMkFeu7eYWsWi6KO0lVCKgGPlN3jb34uAnuSj9oj3OgVMb5J6
UYjROrQLLTLQ1gbgljwxttIO+A5Jqf7wtE9j8SLld3/P2X4rYix1xhzzd9ZH8rUp
XpL+tCtNBnMn8K3ah8hWpx5ZOhf0DqiarstuyKipmk1kpLGdNQFIRk/yykuK0Kzw
TsddGThfnZAw6um4ISAd8U87Pqp5KxZYAl1bQFXO4XzRX07M+2gzW8xA98jhoTY/
/qaBZhwvFAKUE/cSv+2gOGZaywP2SXPeWHpVmyUZRZB61JiaH8qWl90l31SsXNsa
79hx77tNwGWCR3Edu/58fuEmLqbm5TFFk1Qisg2mOoJALMR1wVM8qWTHnB85RixR
lrWWsjbNKLAdnIi9q807ZgS1OBM3BQ5hERv2CNA8JD9saVxEOWYSIcHSuLKek0yk
6AiWaeys+LHU98adB88ADG3QWVM7LWdwxRsfHb2HWb74fX4mPyBRZuQvMUL6+rSe
seXnUQFtrri5cvix1PE0LVwIyIrVWV5Uh2fsofXjU1uPeq2Tv7Mc3TnIieAhWk5M
+79OJ7pLFKWF6anyd5oYMybVBbu9kYtukoVZI8UZU5giqaIBgXIvekI/jFKfdFMa
IqnxWgSzsYlyGFSC9vsnQSBG7KdiHjr6ix8IhEfzTfwZTlM7CaQaJDnDCGxFqG8T
Ny9Rf+B1jFpo0cDAtwnWd8EeSuy7tD1SxZ7Iyo/oi2sJpzcmMvGhq5MF6qYJXFD2
gBy893CWwruf1wNPPxIMd6tbu+qQ16SZHqljmHMBMStp/EFfoJr6oV4ppMu4B0/n
0lSeKVbeVOXkx0efNQeK8ootP00BmvYxcB3eT1CeoYP56oGURD0vrpswfaxWBnFM
7rE1zpBNy6wScv7ZRCAyGEh6MJSMpP3Ha7OoZH2O/DGs7f3nkMd+mjvegedF8GDI
nI1k2FgQMdvXq4RKD8/x03B1nlwDsxeMU7TGZBKv+IBTLt2Ol2AwkCM+MIP+XM+r
VgLSniWqxp44d/lFq16VahNiu9hnhn2upSSo0Aol+mkgIcBp9vIywyn6i3Lj1uxo
XrMA1pYCqJ6tBl5xvYN9oQp9GfNor31OygD5Vq0LHOetHiqsinzAZRI9rUum2EoV
dcmLub4B/unXgyforC6tEesNZUR5Dgray8VsUBJTLfRTxdAQwwOhmn+Q7h8i6PDC
ied/w3GbZ+/1XIfSOTzgp26UXkGlQYyBhjvJLMinEnIJKTbtjEsclXYgWrPxMl0B
BF2ay4mrFGMIIL6ku15aMDUBWqzp9xp8Ok+JmTLtbcbrDaQtFK6D5JdwosBQM4Gj
mE1OdkfpvOQlzwDc81B4XGLw0zljAW8QCgnOkXnK5CxJ3xZQZzBwjo1xcr6ajis8
mMN1TbrBwIAkodN4YrUNRpReleK1RgQFCIsilpHyIm/CkMIgFu15Ssh1W6Wt/Mm+
LNTX5LBzKo+L2SA393nRBe0IprbN8u5sjSotJ2RRzLUR4kMlagvT1JyRZdCWem4V
Wcjw64emaRZLWpdYrUbD+xcrojgMcM4fLdzSLXz/z1L51EAlnhvsD8EOn8Us6scT
x6up7zid2U1aR/xa/ep/z/Rx7k7LmJM72k69S590t8UBOgGPRBXMzyUdBgIDap8C
e2ckoTom8vtAzbPBufydUj/kTti/1TdCZSaU7dJsgb8NYTF9gQVnr7qHk8N2VI+V
ir0OoyNlRzHjticTfuykRvZGBSELX+T7/hDOhyff7VkTe+QqeReDROGwdwoShu9F
lNaIlz8/osVO0JK9IO58APfivhQLIz5BqsIZbOx6ztMboCbst8kdQ7mUuWx2Ofzq
8EjfYZV9dWVsqBVGZlrWD5IRqLryluuecxdXCI5yb/ogdMYuPCznxASlU8C9fybB
TPNE84oVF+XOBMsLK6ZkfVSfYpkj+RJoiS6ct5H4N4m/A+xBlKgT3z/T582HJZkD
HWEuj9/J6Hv9su0NSTd7doptxdPGgsR5jPaWXJv40RcruOliXOiGrMxGPEozrEda
SEMrjEHUrakFvaeSEfh+IUOjIy41tgN2RLl2xU/V0jBQYpcT6bsYQ6JCbmsAZbhw
vBEwm+95JgMXHioTcwPH+VsYoJJbgQC7lJmcZHiqaxdb2DusfHnJWhU7uejT/lXN
7wNQod9UyFnYn8P3FtzdRIqku9wrhlzAH5oSWcXnk8xRkqoLep9IAfdWSfMmTEfT
6gMZq7YIbXcbVFNaoUAYQIs0s6HgT9pdq5YC4r064nWAYBYysecPDSy1Q+TyMEIV
FnXKNh7yJpxIdE5l9wvd9gNCIB3iscDvmRwRk+M8aWnEW51Xxopg6rT/jxoJ1LTa
Y4fMwAh6cybaJcKndcMC+pdrSDMUVh/s6C8atNzdTnv7BuZBGQe712Vnq3ICVJxz
6dUydgRacdP6/rQShr3Se2lTWAZBKK3NGKov0ep407w0QcYj18HOKZ+ZxcopvcvG
qX3jA/ERpUbzLNQe0tTrtw0o5LDM8R7asGiUT619aRtkJYx3UhZ5nFcghRLDsRCX
zFnWF0JpkpSHNzapY73iGfXLigwwyJ61zMA5OMzu5x8gWSaa+Fm1ZYRpdijXflK7
pT88thuoKAOQhlTKPvhAGyHTU02HWMgG1Ej3wR7erUA65PXliZc36LTvKzhEH0IN
y9+jqE16kr72jMBcLve6DUcJMnq+H+E5ou29opFNyzNjvoECQWX2Fn4vQc0qmtVM
BHKF/qYlKX2OvC6OF+pdQmlgV0uvAt9rAcHJ/PpAllw3JPS5t4MSrgPDNwkLogTh
8fmdovzCVxmsCPndqWQ5bRdqZBTIjGJGZqrByGJ8n+cAyngucdCebTI2cDrIlCA6
e13Ay7IrqhMrzXqyZglvRY7QAyxkv3Xm7mFv5iRbQAdd39WeM80AOn+r7IemD6jE
s0NuH+5+aa/+YWm53u5DOGh7fYvaJG9wYe44Gxv1cMJFlr++fHpV8AN7plpzi3uN
b69lzlZFDuY+tfxCLH+85s2xiE75rJytiJPmbm4AGjOJ8MkYZNrmHsZJLOodlU2e
jF/VICIN8TJeb85KG13hyV4UfWK9mphKhXK/4ha72x+LijYChH6AQXKicK++r+Wn
pcBcMnrZl/x5wvooCoq/xYdHOqTrse2ozB39+T4cu5KX3pd2Mz+WzkN+T/ieVolF
cJ0fLwHPD5bQLfvavEiazI57Gvre4mi9DXl3yp4HKvKamzdbxgbibD/i2pEe7w4G
lgs7MOBgCcxOk6CvFGbMI4lybZ3xAQ0b+ti+5JElsQxJzi+6eHSTOyd7ebJVznhG
LAOKBEM48uYx2kdXJs5qrkNh2PGw4qcSLsSAB70oqD52dYR3PytpVWbUNAFEdktJ
Vk3DNLfs5OeOQsr9MUKHUnb94G9Omyv4SeNth1wwzWx9rouj23peFczAin969IO/
M8zw/IY+cRJEeS9R4Vbwk9eEPvDZmpTSwVddu+36qDamXirNgW7QbCxc+1VLEpB6
3SuhoIFtHCO1sk5C6zthEucBCKi8aY0HrybRkD9oJfHenOOrDywItbJcmWVR2YmK
EoSj1nh/GyZ+o/vZ/I9Ynh6FE7I2ed+Zl79z6nZBgRFDeRnGZAY6ueZuxo4vKDZ4
DyJlYREfFy1S+3Gx3XSD5l6Md3r6rn7ENiEoOA1bLMQwy6a1SwVp/IeszwIeVTg5
BuC87mHkTxlJfjkkH2O0mCyYPWQZD+zRTc6mWo75jfPysalUYdyUEiNpJqKAFnhR
qqbrzM9x7hW/AM+KfZApKiOVUGAsuq6AWwmamrppvAZr5OYE34rqllgkzuoabicV
AVZIp5C3fEOpPrlU334435sLb29NesSbtK/VeX2+sxPBamQ1D0QxPtJwyBmD2Vzx
Yp5vBRI9sTmdr920NNgZc4d4EFnXwBBRkmnjR9CiSA0wdfMsZ9QToC7zLwoZVOfA
pYt8YAY33nBK1LXZ85W8IBWOXcxprYvT5PM+uo5KEuY1P8BOCLTq2ogvmLV2VkjQ
n3kjW3cGYhrT51i5ATMD/96qDt74IYxKyHbnh5Ia6ZnFDXdjTuBsZNYHRC/DLRpi
ufyRkcj1sXBKCOHtkOwv/1UNg4GjxR7UcxRU/arUQV380FMN7yfgJZmTnhbqAfAU
Q1o3wf/VoWoICFoY9alWd6NA3v8Hk2uLFiJlsQ6lSnapJwGWDDF4h0dIDbh+fBdi
vQKeqUdNLde0eyHuxB1FFN2hQyScOLBzvdllBw6Hlu5/aTaUiMBW1Te1X4ImYsvW
SRNVPGR6+EEI857pivJ0bGHwR72mxtQg6Ww4+XvqhktPGTH1V1w+MmTnGUIYFGXy
V21GJYx1UPn1NpFREVlwH2FiTaZOK/C4rn4aSYAseuOc4E6Lzgi06O9uvNqkPFSP
0rs9M+/naojcl3E1NeIQhmp5URFZPhk0YQqDr/zjxDAlfFP0Q7E5VSg5V3vdwhnW
GwMTaxlzUf8T4nT0Miv6rlT0I4nGr9e3yISasvEonsWc0FERGyA9fqv1o/lA11Vp
yc88IMgCvKpJvOamBcSAUOH96/w5e0TCwyPJ7+52lSrBngYdw4Vab8ecsXo+SdIm
0j5ls3syQtfghUPCPEvXUf1NPFbkRVOrOClVOeOeuGzVpEHy3GDN/JHB/bX6NRq3
lBqsx6JzI29HLmyKSyIX/gKcsx9FYeOodsNSracSzldZ2NlZ9Eu6vEh5NQzWw5UZ
rqUtvLJhoy1Wl323cfN2bPFYS6Ie2WG+zBUMedyX8jzlURsiIP/8bp6a3Xjm+7r5
3Wz2j+243j1wfG3x/0jmQiQJu40VuTeHTzAybgen1hRiSarIilvi5Vy4860YBikG
ZtwAn9nn4xSp1y1gKNH7eRh2ojGk8ExQ4E3EinE/HDqSfIi/JqiAKxqvI+Me9hmq
KFXtIb6at66AkfS+JyReab9a0zYi22RDD4qCzaTtP46Pd8u4DsdDic6SEbgrA9aC
sKEO+VVmiOYi3eTKxJjgyp8xpX5IYD2iqHKhCSDtluDmKTf6fx6hjdmKR7KSZtXu
UgPIlCU9mENrsjoAzD99kLVHdFNPC7uXF/fZ14S3qZziQkqJvKGxg92BWl3I3fXU
VREvgWWyA/KUEGZ6R0cs+IDJfPTHX+7cFFoPF6clHGgLekBa3eHZgoXlr1IFw2LF
I2G6Ioawo2/46/zHzA2hH2kLy1VVgqQd0C2FI++4DQjh+I7O91oNXFQNpv2zuQdm
T7ai2lC8cif3B5NxTEnZ6dU3+CYoH6kVRi4lP3xMf5OfslIN3Lk4agTrS4/vWqJZ
i4OhWkdRK7x3FrEh0a6nipala9rojLBokqRIwep97fGWUHFyJraxCB7vShDIWKEG
GWBinzouF0SF7x+qtUWaHg0rN9B3KSoKtwjLCi1B+MbrBRtbf1cXWshj6B/QixJJ
nongzyCiwrFJOozED4mXc58YjuErcXSMrpREdTgZb5bi5fCz9yUVuwuEzgZSize3
YbIZsa/cRDk3o74zfzw9RiQIJ3CwF+4RumclPwl+j3lwGMVpe0i9dxgnRn/VAn+X
l4IZENn0mbLR79TJoJ4lEn9t4g5gzZAiV1X/oMSw9n7PAdOrgNs7v3ZsnTq3NZow
/b2tE+VDUwyRuxIiDjlfhb8WiPd9LjE+GuKnvVlgWIGLwu7fwScSULP23oH0Menu
DGNp6PCoC8PzrnqVgyoyG05iqY3BwfTWW+hlGP1/AGtiLB26rKD1uS+EfNG0vY9A
D4PPajZCryrfIimHDBbtjzpRrwx4fSiLOPBABm77QvVxJNLGftIeq0T7VHHcCkvy
G9JA2+3ApLtrVKpNgo4tNRawVy2VuXFzyPCkwmC+SENBvTVWxqF/FOCaJtJK3GA6
i3KFbA32omrwaAaRx0CH3is/0D4K0T8wdAeL59M+eEHMBXfJmn37R5GFk/2VgoNF
OKjhnOHcdvYHZYBLk4F2L/ByTzFhJt/p130a1RhbCOhq7ZH1NXhQIo+JugmT2u8n
HZS3OudZ3+CUluCHTISFv9AfVAYZ6dljlaTZ3UU3svMt2X2MCHMQwz/pbWNBnn4C
KUpw15I+x4OpvCsyjSlJFjmLxumVDFhdwwZcRS9NCkhzs8E0wENS98t0W7/Gj+93
EV70rI0l8RU4g0xpzWNw37fRl15iK35VR1Omob/BOSrmHbpbSRU3OPHS5PHFP3Gs
gyV88ZgKckFU26Qj9moOwqnhYFKVy8VXwVe4FbsJwr8gN83Y5xaRc8X4Xq4O/e4w
9tYwwH6GQ5pn/WW1tEbzzxfoCbxvjnDk6LhGCu715R2gGkasHn1XZ0ON/gfyiMMU
Iud88w/ABFTULS2sDeJQ8DpvrtZSiR/7s5Rf7Ror3UW5xMqHzQW/yC4N362pHoOk
tHUQ1PYulcNzDadn0jCQILHrXxGhxbmJDmL08sJuDq8pqYLHSBB1Ep4R7CTBl6AJ
oeHiZmo3Fe6RPW9iN5gVjdWpDB00JhnP2D+TCci9tLBUGggP2FKsVFMZjUx2dXuv
MxMkKD1kt/aKpCGM35Sfly/sng7yaOe2kswK1/ZyBjP8rEjTF3ArG6wKckN3il6v
WjxrMSbdnq5ojgKwf+RVid1Ue03c3/Vc1fr68aGRyUOP3UNwYLSJ/T1PQQbaqbiv
Xi64bBM/aW3RDPP8tW/uzxBlY6/g+BuKkejfmXODJHnWm+aruRPCLdzidHnVO3Kc
Wf9rh6oNjnL0JPPvwwIhYBlfPcQvEPUbM/JwJW1AeEUHGUcpFXIaL/8oKNAe1bsv
lBKO2z2kwKsph03qJeTCK/esc9dsbywrTfnnLZ1fIgtYO4h4szBwC5vgKJgwN00D
+1QPYt1DiWnTUy5+z0/1JBL/hXTQv7kiig9lpdhzKfhsY/TgK999Y8Jl75V7Zeiu
3OZdKjojZVxLPaWWcwVAH5BEl3+wcLBF0Pk5MG5OaViUil47IxOq2Lg0NPxdL/Y6
teHJqcZFo1w69I+vHRQqkC8DAydrq9cCw2gieJvLBctEf/watq5H0M31KZSVU9qV
tMOthj/99o+uLvCrB10QKylMLedN1Gz5IK5uOKqsGz3s7uOmHSdth41xcWJZUN4d
aszBkB8cIodEMOPBOUtlqs1wwUiFdMJl8xn7fbKSKtbXBaxTj/GMLGgGo21Fk/Z2
CDei0gNKQpm9tKarrcDFwBGVcLc4d0I7i3lDu4QDmZafR8rFTR85ZHxJ38N/8vCG
v+MST1z+xiMzU9u2G6Tz/oWRBmsB62tsgPKSVx+DM/vm+DIz0LksFaZgwLJpKCYp
flsswYB1ZY5zqWQD3oGJQ7vatOTSQXgObQXL/IMsWPP/IUb4V7W0tfJWp7YP8lE2
hacdStwb3cTVyrCFLLYQ+Gqnn4j1kDASEtT1Mp9x6oWZxGPtorpTNUeNI8BFEW5A
H0T1TiqEpISfAZuatgXRRVttHbFS7a4fIvDBrAVgCuSLv/z/mejPwSIOcLGkBzPc
bAtPHrSUYRJCQNE9TRoGuyC6VTobryiqgql31i9OiYRS9B3nDVamhsxwANmyU6PY
hhMpLyvSlZcAo5YCSJdsuzLaxSw7mZ/46NnysJU+U81LqFUONiWVtMhEwWIUo6Td
FJj2Uak3KCn12+zMnCIcrMPQPJAAYBWhyV1IiSsrd85xc49Z/+JJivk81fHtuOzT
q46QkNfWlqGv0cuH27f2IODqUG1NWVQvNiWiQxHHoNGvnGx6myLbWhMM7PcmTt0d
wbjnxwyK/v9MNAlVJlR2+/EbBLufpcm/hguH6jKHvaKTHsw/c2MpayxlMGJwzBNL
fUTEwdJq6OCQF+ChI74PCY+i/63l02lTMiL7VU/UafM3YDwHFeBpHPl/IdPOdDgZ
0fa30Mpik5ZCrXOr9Jid2pJ17vNTw/O5sA33zwZ8ijorNIW0PWfCA12p3UnAAuk5
Z0ut3m/kTX+2KI+xsCy0WzkMhKcKSFTizB/5Uhqusztmpn9H88SfGUfc6g1FJTAq
nM2Kf/rD8ohqDbkH1goFa6kby2Bwhbz6BdK2s43i7OEPVYdrZ6js/eLLkUz8KvG4
JkYj6D9/wq0zH03Cbz5XAzyXytLxyz/CiTH6nWQT2rLNQgtzKfZCVF8oHeCK593m
rxewS0ijKnFoEtQPF70LIuD2JBYo4j4vaNNbzxBBb+XVXSg1GcdBMsGgS+Ayx0ZT
fPT8SSLFSWLHgr0w09bzq5YSz9OaFBgc5g2vIP391OuujSkgD8AVqH/4BqBa3c7r
ncGBggKpsferIGwpZNBGw9aa4csWogK1ZKqcmZFPT5tCDtGU/rwD/xc/pc/HiYG+
pS6sTH5JSjfkWgWURrgdOKd/X8IX8Ap3Ee5ktXT2gLvaXL3CkZoeLn/cvPCHuCOk
yxZmtmuhzBtOTEtbsJNvSPRCVthopcIa7byrel0WXMCrro94+UVE2wT/+NJMNGcO
bgJCLI2uov644BJxGyG6+Gsf8MsIr7oUXwX3EczKZZ0yUD4MUk1hNOfKKsz4oLSC
PJKI7zYbfchpBrIpyRK5GS0INiZDzDHQ5wXtybxlxBk/KweDC8fkp/VXc7zjHOe1
y9yv4DOZ3uWP0EgNOhWHIFP9wJqgqj+JR3RBkyEjU0bu6yRz429SgBAzWAv0/fB1
u9umBh6NBnTSO9TfWRj8XY8yJBN8xlITBQGZ/hpVUTaiMHPvjfASfAMBe6y5RdXq
bHj7cvLjdTS0a5TKrTI7yxTqdpV+CKp3M3a9X2RGe4O4OZNPTjunHbrcldENNJeZ
tiZPq9Zws5KEvsYPX30Rn8hnTitBZt2b3Vl4kfBE8HiLAZKBFpEUBQ4Abv2q8ZU9
/rICqniIfLZ0XhORs6TA3/BEeHkdHoGhNx01bLsLEecmVjNOTBB1f2KNC/q5B4/t
EEXN3cTRZtGoSZ62vNwR2gm8SYL746t0khXtnETtXLB75QEeo3KLhkwAKirQy+mt
zZh7hCAOMq4MxA5qVeH2XkpVvmv8RThXM9891URB8mSxeYuf6akzohJlSJmCV4JS
aMDmoYuX6N5oDE54cqrKtfrSUpjivyQvgluih94Jy6rIf73q61FAhI5neibiQfTu
JBt0kwqw29TBB1pNRTfrvVCmlSV1pWKcA8nV+J0tQMz06zlTaTpcY0vS5vnqGfgT
2UTikIEG6fdZFdLwr0OHkBSzDVUoF3llQ67JODuLhHLS4ep6WXIRfY91ORjLElzP
723FDn+NCWpzOKjTdzUdsUNEwCey4EHOU0WW2VAEiC230MPkA4q2bzWQiqfbbpAf
ihc7cIt4JMwwh6SwRXmdsdmUppUjhKng6Z/OTCmZM0KkZwIDJU36z2LWkfp7sXOK
49xpTfcIcDCoUBJTamLtC4hAmsnkJZ/BtmilC8Wm0QVTUiPXylki0PIdWa6rk0A/
3OHFpT9dv7JC293GzH4PlEBhJ/kBh1gJU7PGRc3sSijuoxOe2gX7rPu3yUTebtgR
rED2oVEDBxt9yMZjYRpV1WkNjb8nJjHVRni+5q7NpqlQaskqrkKRw1MKzDCwtTyw
hyrYJ4pla6mDGRCUVGUGqeoIJI8qYcIN6atbI2oiYbwM1av6TmtJO+fu3QajG1tU
+Tvb+jm4Aia25+W7OpUHe2OQZ6XK4G5KjumMIeIP8FvCYyD8lrSZ/x6T1OxLSaqR
6zVAm5dlmcfUjN5oTONDt3n2aqLT7ijrFxB/x2gauSYrJw6uexRTmxQydui15+m0
94ciNO6z4q5Yns195JpErnzT+oEvl5Wg7mo8BfOLyfjaCljktcOrP6sKWNCy8FIP
giJpKTtgGa3X7kJygIZXejDl8lGMeGLASUjALuUwo2o5hTzfe/2bd46TsjENVQQJ
cagd6AsJS4VWrXhcfQjFtyWxaNzamugwgy6XdKIsPcgbwxhm6IPUtox7TNSSDVwb
9/NtDV5105OoG6D33/Z9//g6IF78hawr+J5wFnBX8pdM1HqmcEkY1yYtiNY8IwNd
LWTtMr1y7oS8BvKREnKH5y15PzioUbH5pP4dZvb7v3kYX3KXCAJQDKrA29O0RIPy
M5LHysQ5aCmfGoNlINH8zBfFacP7YGBAmpiEoZmKTk1Yvc4XgSCdmSctMtpTDZsd
uyS6oxyknIJVHPyBcKn/wrHI/mKnNvs2oP8SXaKCD60VofgmFEKm1kdZzAYruICG
L8CnwvQ70HBzGJtXIOX03O04D93JnIKw5eae8FQygbBXCFT0N/jBLZLf7RmmtoVV
catRu1qjXbJ2y5CVFb+TB7jP6Vn2SRDBXylOnl655RSDAx9XZp+39r99FtT4wbcB
yVXixWC+7S0NIYjLcU4JmUOrmhQazTjusWW4U/Beqb8nHis6ogIICpzXe3F62WA9
4K+od35Bd8Hos91Pqm0tcxsizS49H3QYXatesTGxNNA5L06H8Xa22Kjuc9H+LW92
SLZxUF2lFfEOGSTnoCvddtKbopcJ2LTLSSJU1CPI6o7Fn2zK2hXU0Sh0tbiUhKCz
zauABJxfUYo4UppxM/RnU9jzeBaVj7fEpp2wG+NpnY6YQqbPuNwHhyg2Chmn5Sr4
eztQFxrGfy+AJLD1Is5uigzVO7sw6j/5KPGeTNc1sntJIWBeDmlGwtX/jjh5u+rI
FVzbkJ+pix3NoHInHrGBjIAMBPCKI6r6vsjBJx1+/Ez5RTc0KLA2bDpRJb+61vsh
4IUO93oD6QhSTLSmNNrHoc80ObPlhH3bT8NYBcuMYRLh/ivh2bV1yRc8bG9Wx0Ck
s+pt1H8tBgTbmNedxVDZynHrzndjlaWPMRRC7eTYY3d/CSBRiwECRZrEjytgvEsj
ZWg2xPm2o25sYGF7ICADkLsylXM0rFWS/62iUBHna3GnoBj9ZHbhl5TzmKaXaDSE
L8smt+PeuunIhBw/WxItMN7EEBI9jNPyVwIhBLMniyPOM0wm7R07t/vACgz2y3vb
gQodVACGP/4beIdw3Eg85vvzMR9jXQo9cNsGuNtAKH0lEjfk2CJcHF9oPKL1LE1g
QwjudcPfzT3rT618SQaVV17YM+O9QMpUJb/MB1274KZHCwAKigm9XSDzIYiHjr7k
AT8/enE8knDWEej5Csou5B0vIANNvyTzUY9Zlrf+trW5JrbYyFYyXDRlk2FoJuQx
KghReTIuQb3giEzvN/ljvUsoW+Z0Otg+W0R7bUvpLS19JQotxK14XQBBCGS4dCco
caFd07Lp1pB0ffyN/1zy781NIeReqFupE00/pKcGgVqx9jd3dd5m6MHlDh2GywtZ
S96h35FjjBFhSf2VLYP6f71ir5tvjYQ5yqGKNJuZabIfW9T9PbwoWtAjDBxQj19k
1/sT+V5tW5ThSATFdsa2fLj+QSvrMNqFcX2EdWMl3ACkqSTj1MJE2r7z5fk+H6mU
lTn0wipnxRhUn0x/vVCGKLVxb59/Px6reU0ASwXBU7PCo71joX4Wlszipj2L2caq
CYMYl04NIAWtmiabdd8qkH9xlBHVJWqBJ/WLqNH/cqP20uu0EKOoFrdRlRdjO2Jf
O4Ewsc4YwPIa4B5N2zHR8hqsprnnG2MDcrsFtmpVXYViuY/jU6RWJKwtQOWo5mK5
3478ttwM+dgUrwBIgRG41c8efgO7zRoVZ8GIOlGqk+lCcGpE6o4oZMqZrwxEqTZ6
qWHzPifgc9IyDDmgTrazidwKU40Z0OdtJ2sq4Bu5gdt0eVv4wIOVEnzs/6bYcu+q
fVqlEqWbzHQNi8O1PGXmOTGx0aNJtoiem4RQ+udVdeNDSbymhD6K71+Bm85TMTVA
Wj1WxiqPef4DLlBQfXOmOq5YR/ujE3Cx4dJrP9fYBJFPuLX/1DU9rD/awYpdHV//
6/l3fygU90gdGfOZwHrKlFkQMkuL46ccLMU1bq094p/frtIwh11NHlyfh35MwhGl
jyUonAl1SmhNDyN2dUd15Br3RWkKySnuCpllRQYI2jZjKDlkYXrHpqYz79Iao2pb
qmjnU1O+atczBA2Q0+dviT6MsttWcxwuMb7nHc1ozYr12O/rOeWUzA7RlBYsWh9f
SBNGwqmXyjG6ZiStmDEjHYbZXehsxfLZnwTxjtzPuO9cS0yFK+4Dpp5SVmsHJ+78
6gpvpfSmcmlASHJrmX73Z8mgRDwgZMXDkjJjAKzM/gaGrrYoO3CGjmbQegAYk1D8
Wthwt5MqKvIIJysWn0DxL2jd2UagiFW2sjYD8MEeoUiYbE3V0djTIBAfQiNDJ6VM
jsk7/sZmqMxql0bdW3z3LCeFlzq69+675MqW0EKWGDg7RK3NW7x54FFO/30GKsSj
q1mNHQu8e0j+xUApQgU7K66iWPd1MPE5FsNAnmnWY1KCG8c1sgnJ+x3GeCwhQT/X
dmQhoZqn9ScQDacd7oWf8yXaW9MJ1k4E24g9xzh/DCsDe3QGTb86aema5WU+ez9Z
K4POL0fiOWbr8H7sDSy/gOPjg6ocYHDDzoOE21B6XqdYn0v3szgXUbHykBDNggko
BMkYMF3pj19BqGS8xxNap0i0gRheo/0Lto9f0CIZCLAvfi9FtFhZTPy23EphEk9a
GjePbZexU3PCB96+aBBi6LDMLEiQHqonb0/lUGliVxDWTTMRfuZQz3U51OjT8emi
aTOW7matzqyXOQjsdeFvECh/lMVMlUGiYYY3BvfV9rr9GQgJjwIUr6NgjdS2TbqP
eiQZDRdXEXSur+Z2WDjPpF4mv+6g9OvHLYwuwXJacd6t/u5c5zyQe/cFT14wCaL0
Ke42U7k6tRW1fYlverOKYLQ3c46poDiKXSOmfDM/LZvfCD5oy/Ra2Donk1Ef7sYZ
1W+uLJmymrRHEdAWTEf8Qlpr4d5Ie1VSqAAW0nh9o0N6mKh2rMrYSiONoIBs+sHd
jNeo4GU79Zsgiq7jgoLTfOk4fEKhvGIa1Q1Edqie3NrkC8HdBxFgYY8EELuzK/WT
oU4gdbqBSPP5SuSEVAwDwkqHAHVnycoixYVX0R9a6kp5r3h9H/tWPo80KFmWePHh
yEX6pjmOGxyGL77bRVb2C5swJ8L8WQZo6fULO62KkiMqhNV4mXN6tRiORm3E/5Ok
WGL5oCpzy0iPZSGWrpwau7REBu7oGC7sci8XV/dmvuQuzubJ/UadhcA/27hLxbId
cAXGYLzpar2U22heybPGXG3hoeIOVRdsiFcRiHtv+mFZQttQfL5F+J7Bo0RY/Hkm
7Y9UTQjZ+XVJ0gkyY+OVw0gHaUuCUi6s1yf6OXSjnIANIdaBIeMC4WnN1YkQStnH
0ZYkr3rk+Sw7z/5qGrKxM90T630G9gQcd4szwelQG53WcaNuNH8kNZynJxGXq5Ro
x7qAZPVwMQCAx3sNpmAY/SqC3DJPq8kpB5axcee8kd1Z20SUGVzPZQIDOb89kQjz
CZdCrajJTpTQHmN206X6HutEH7+S8kh+ZkUeZQcFrdcgDphHLYZPzluF+zJJAMT6
MwwbW8U4W4NCOsSnqnKZH2t79k3Zwiso6tPGYnO8c660LkO006cFxwKs1fpp01Cq
yEa41JBwoobUoa5g3WCkmTUviqAeZikzyGxr+dqfy/JkuKSyuAGmSEA8kNagT+6c
KUcHp+UjPtd9PHRTZtMeWhyLz6xmVVNJaqqkbNFrxP860CTn4GOhrcHwgMfx2Np+
qZHT5FfkzS/mkqDMT2YoD29fLtmrZCaM94auQnn3rpNrbU85TZVhKabadrNoaNzb
vfCNU18+/Z6yZy40RcBzRSMtkB+/mfVQZg5aqWvp+XIczgoz0OPEmxRx3tdBYo8F
Z1dB0vbfg81+3TKH7zY0lLY3slAgpxsBd/dQWz3mFs08h2FKCVcluZldm5EDWFbg
5FwIJI4gjxE/DWKvE0gud6DuBs5ZIAD+3niyzzOXShqzd+JcrHV2YSXwEkJCMOz5
P7ZJk0t2TEuCiTh4a+ei2KpX6JipQxKrR6GirsjeDJwwEbAu9Wyyl0xPoaVKycoN
Cydtg45RZb2jTKi5oWDCPes8QjWcKasiYaznThwRQl353qacjPfPaEqUoSGM6aeU
qXoqTNxq2BTdsvADy5fDQxpFz4bdF7iS/lb4jl3sry2oEp0OZsP39I8/WaQUUy/5
Rw29HqwzBMOdYxqTNU+KGIGb4D9GfjTq7n5JuUmwddVD+Q6stQ6Sxd/h2FY1l0H7
AJgWQ+vlJw3GCVxOfb5xdykzNSvYoGAwlgNOOdYWNkYiB6xiwSFM5QHK+4QNaHlm
ddMIt/0VU3bMNACaMD8PyBHs3tIAdViHTAxj8wA7ik1zvdn8BZ1d3DJkChXQo/b5
GkysKEHFVnvlF6bjnRk/bfFLYyqzCy55pYVmp91BXTKzE8KCVY6ku2RQriSqJloO
NgGFPoWYZssiGyVyDfvcV7IugW2HuS8hTmqcHM3ZUWk0QrDTmWZWI680x60s5LYx
WcNum0Nw8lxYNRQcvZIqcWFouoNycnsU6IZF92WFLubk5i5BXiqZt9gKOxIcOUwi
+5SdFjiC0MaONv57H7sfrLVOJsLT8nC5sbQSTgl8libloTDOtC+WBw7Ch7e7YEY1
Ho0oS+RSp/WB2B0f7zbpgKToL2YUQ60uWNQNdHXoy/VnEFOvp6MccEQWQhNayk+i
WLEbZDWBbJbz/sChMitvNDvMUp1bXvMH5qnR2VHClVq5Yx03Dyl0yBc8bmPlnlGY
TH4fYVDkQSW0egrE8/56PR4rMZbfELFY62g3Cw7VnPspZNvQmYISdzfGhJ9EZsMA
7MVLz9kjVaks3fe5uLUHAFhszgEmPgOeAsyXlPJTw5IlZwkf0XwoFDijVTnYmbfC
Jn0aqPlw6cvf2q0qpzuf1O5guK9OMzLi2USMK0InJ4wGM4BgDdNN0SFQD0Tmsp1h
SluTJUL5OrzdEu3a0pIIv2WvTQov3+7DXQzJ6Cw4134RJ50gSMTDQRnK5lLdVh62
PUoQZZ2dPyzzzQKyd6qg0sntq3vz6CwT3Ase5MklYYuNO9GbuZBx/4FYG6fpo1ua
3/od1goIBwKadqe1FXhr32zSI8dcPJGJxfugIzhlZIBLy2Ah7OUGhIDwHcLSetoy
WJwOd8hwz7Kb2XGK1RkoVsRZDpbc3VA1C41ZhUmb5xUWeJ/hEmEGHMa3TcuEFw7q
lMPYxPFy1IyQZRnbDaHkRsTDeIbXJIJ2urKivs6iYqTJArNvL2aEMHCOtx08Wou0
asEcA9nc+h4ZkUPP1fk/Z5e160/dzOV204qIb8fx6kLdMH9Ixhh7f/J6bNPO5lXt
h9GJwnc4xAxnMOh7+rAe/GL3k/ptn7dhVcUPIv0qCTNnQkggoLEN2pzExSGhv7Hb
6B/bOAtdF5IRqqQwbWiGjPPbIeEtgWkB0br5f4o4oP4B2qYoLD7TkOWh2Mp0lUVS
1KfqiC/5T9Bxi2Uwmx5RcU7dR5XV7P+tJkZ5/ghdb7n0DhSSMF29EFrAfaAQKOo9
TZOvDdq34MwVVD+r0AGadVyWhrfCbs6WXSAHN74OGXs/hnIPQtrX/QyWamJ/ULO9
KgQeNx46oC+wO9Wn6KHY6qpZSEm5y6mEuSGG6wl1pkWUt54A0x/cM3/yGnJlGpVF
Vvc3rxpX1V7nnoroIDqbL8IJmr3olU0s0+s3bzVBbwv4+hCv8OOEh6k+UUEOIp7t
LJHHFdTHfUx1kBk+TkrUZQ+C8xueBdPjdG7TuozcwWKIsDbROv99y5TSL4c5TkX+
f/8Lwg3xSqbHntAZ6srPzSWJWLfHMyJ4LNy9n62CRqmeM5myelnc1w8hFYcxYIbW
ohLtCnXz1P+IK0xhndyxkCuokpt05o1NQdggRKuKObmmaqwMdwe4iDCyjKRp59Qd
PZWTl+b7dHRVcF1K/bVDJDyAbT0l9I/Ba0o8yfdGmq157akkzDoqR37IOqilP/du
Kl0NzQK7jX36ZogNIy9TVKbE0Xmi/DCc5QLTKEfFf9JlBUS1DAxlb8oRaepr0oxT
g6NAxKtZG3eRoV+/ectVibSW/TkhIrxfURuatwQ3/jABfGIAtN4qLS2GHZNRaJdu
TMNnjPQ2PhNJSDVbCWCM7hVjU2IqUuPXw0FQesIsshIXT1NqoXlsonjoNYHd6hpz
HMLwDg9BdqJJC4+csOU8Gf13KJ4LgNcoGWVd1z4acIyxEoWhHeVYbtc+ofeggVzs
eaJ+tB+LN6t27GdoYHMiBRAWM6Gy9oCy6dXZgFloZNuLu757w8pWffXvwtm5edg4
rWESmz5WADT4fccOyKcex67Re1u+tktwfXhfuQAuxffMMD0AH7lxFf7vCiujPGGD
aqqFir/1JLUjbIkh2ZR6WIKjLamQOtfDkEtmZsbI1/oqxxYdTFOoUzJhuUjcD5RT
KIHPBhIPpdlR32eKIQhh9IyQIK/Rs7H5o9jd6H4sferOyFJsEFz5vCY/MAeGPVCF
dMdemNvcdVKR/Zs+ZSr2NRoQFLNyMIjgRnWhHxZDElUJrT+YcoC+CVmpznGhIgCJ
eL4kPirrrBicgv+ycx2WV1h1embFjjOvwxn2bErgxDN79nhKJlZ8ep52E/HbTKEi
MT2Y1k5NuB8JRxO0BrqOUn6Lietfq2e8VGAiIUUkiIcsG67cIu5NkT9L1OE7yqx6
0t/VA1NrM3Vl9sgg+48ydCxhp73VXJzfjNRxpgXTM7xo9xebJoTuePqMHnqy1yEO
a8iwxueFN2i7lQsqtJL4+TPOHCpi6B7qYmM05XdS00usMjFgSCR/ArA6ZTbK5TLI
imzRU8b/xv9+znP7zX4JCGGBNt7rLLLnkzlACy57cZclDPhALMc3+TWTU4FiGz22
jLSRdYlH7Cjwb4tByST4OnAZnPTCkhouiBRAy/Z/kAO1W2jE0UOOAXwK008qKqli
8aq6J5oNNa1Hm+mTURTmur7249wswqpFqVatuz4KzSY6sbnlBa0EXw7MoGU7SV+6
ISr3Smk5ZXnsK2icjgXpGZBe08F3p5ArEevWQ62tl4YZVRoK97YmgryZGauXospK
bUq/yBg9fxmYRR3SIihD6nfXn3fWw4PMm+FOpMXV1wBejHWWRsbllTJSKm5+e9RO
9iAGWG7FRKptN42XHmWban8eRazrZJzvfkxJ+BeRyjeqR/1ZZ/FE284pMrOdUtZ7
YXw0eORLck0jfK+vB7PSCMEMhzxxPVyJEBbfEGcme+C+3MMse2vRCVbk+W5NnlSh
3IsXjgVm6a49HNMsSlWg7Ev+XMiRWgXvi9wrAw6Dq2tVARRLYuvOXP21DWq2JtEt
XpJ9y5oK24cAUR97ldNI30Wy22bbwZ5dbAbc7vH14TLt+qxhgC+lZFcZxgn38JeA
enmIBqw9bkGRhsvo3fDrMLdAMGwtKHgzjadUSh/fn9Fes34YUzZWTvpTkNCJWbSc
Kt0KHKc0Y8rd080urrhEXMCi6HbZMTtD1aHEyV7TbwMQg5zr7dBHu5Pzy1oppnNp
d/j2kuz4ShehBAjqp31B6P+i10oP0M2ajX3D0r/bM9hK81bsnr9/XmKBmZrLOcaU
u067eo8JooQTBDR4FczgGF/TZjgzJv9BDtGOEbu5GHX/Cm6bo1L1sRZYVtZeqf42
+JrBmTJVTcmtIbNgieXiJ4lZRW4l86FJ3S84S20YG62xW4MM9Mm8FwJzkOJrBqpc
b0FVHCrAD+ncp2ThiOknq4c+DNbSvExeUSbHVwAIciWfcxOEDIvoujOSW962nmBC
QSM0hGFIlp9SrbgR0G1kkkPjrJa9Exl5YeQE2pNAF16AO/UcNvHAnGfvuL4ufP3i
VdnbfsrfQTqvX2qktsgUhZrNTiDshfXqXdMRe0j2zoIDrLy6ALWwLKGuv8rU407o
n+XtG0vTHJLFXSFAUypeWGzEPlaNn/OM+IVPd5lsyQyNfl+LrD6BV3h54ENsrVTd
bIQ+NJWjxJd29YWncf4vzSZLH3Mp9hmS0JxVRhYayXj2tA3qI7LlejgFYDy2fqFr
ZWrX8afs1C6QQAH2zs9FWxaDyPS/xCjCbrZ/KK4yyOiNSlpVvEKJ59esJg9K/MMv
QiQPdxa2mTxuQEX5FsyGkUKmLZMwpngZNEjuwvduBSHjCKdt9qIeZ7u3sO4ab83J
X3niLUhrj0xQqdCXOqzqcaRWEVVjXbVFgSwYGAr4y5aa0sonNf+y0TgYmU9DLXyp
JTIdldmsCe75gEuWoNujU41qSWzNjOqOEy9skSkVIL18f/6lVLUMiWwIyHCv2ziI
ic5Krx8VHVyELttxUZUon5z+B+mc5ieRSO6udHFI5Bq927XNTTI5aYRkYCy/AGbK
CI4YM6m3gdbzzfx7VMOxJd7xSp/w0FlU1GwupP411kzMzqoDdDm68yV1uuiUmgHS
GZcQa7Lk4S6DbwDOMlLnFoJ1Qfl+L9NyR4eK4jjno/kp5Xhov5Rh/mQLbGfFMcqQ
zWgx0l3cbjSxb9NiVbrKiAur4ArYjRSQ10iflGcYUnASuLfWOD2xiCLYtU/gUG1j
iVVxiAFWTydSDYz2wuWMynRm2lkfgn9vhhrrPJNfTV195Beb5S7hrJw53IoIXiNc
buOI5fdIbouxgJCp26uc9eDWkZVxub4RyrDtOp+xWcznI4LEdH5gh+PPAE8tST4L
3FDqCWgTdbRa6CBGNrxxFYU5mCsMg2vAWUoxMtwqHpwdgZw0ns506uHxG2bMOIyw
w04ZJgLLZXQ1d5OkSe38NK7q5TqHzT5xnVX1ZhxrJ1mZpJ8mlA0R4zKBtncoKcll
Ybuhjtz7phDdaoM7Ilv+gin7DvUTCZ6EuGCM4xbjwZ1DZnHOvbe9qk/4fSIh6XQW
bN5IFU5U7ueBHNoOAgn9kDgumqi7aCk3A6/YS4WYv++494KIbg41nl3B1a7Rvp5H
2qM4hXCDVAy+whNSp0pGv96fLxHWiwFS55IRGo/bKwfBQnxlgVa8h9zpEdByRgjq
rnVLl5VroaDDUJam3va9W8vpotw46Tp8HR5Pt6OFNnULb6geu26/UxJ1T4n2ZCoR
LYhFhpiAbO2gcRgwtM9kQznvymPaI9tLdDQ2FHtA+iJdiwcldHGWgzB/5lfJPupI
0ivhMXxGq+5P8J7iagrIJz5ZfQi5xCb6y3P937HltxmgckGYqT8aUq9ocbh/XDJu
vk3B+4GCYk4M4YqX6MTrlBywE+YZAkSdOwEufzts2mNhQMLfKg/1F4gLwNpy/kxL
6cXGl6HC5246lHzfCndK7VjoMuEaXCvuPNdGd11Qz9X4/DOTymJBdIplSbkYOQJW
aBX/0xHbwqcCxUJ0/TiGuOSzjOs0RwsRcYzoTQvVFOXz+oSDQRrmmqAXADydiOxa
d3tPJk98j7aHzNYoGk+6dW05bboKN31l0uyiO/Ti8AIjPTr5I8xAhpyuzqdImhgu
TfRfhnW13B3+iMowvtzFR1Qx1nFQCjZtC7WBP6iwvv88ID8EfX6VHmxLFMqWxBEQ
RIQg3P5uNx2og9NKV8U0uFY2go7moodea7Zci8+QSp4C3cYUrXg0XyfGkJZazv+F
2qaFBJUk6/opQ8avm039ArC0b9yHVEXYiL1hvDGne9oJM4A8BmGG8Rui1zIb7rOv
EPRK3BX7ZMsA/MzURidyYIX74BUd863j3cUJrnaw+oi/IdszDYReTNXGViGnHLcd
Bg7g7heWsWu5YNucCDr4n+CDupl7Cj0MZojBuzRBNq83YFyhUZUhrd0jiLXkvqyn
UE0BcuSt7KthufSfO5+dfOipv+Hwz5E7cmAD74bh0Et4Jco01SkxQcK6qeuwOuRd
40zzsb8StSwOLQ6SErvb7vqSeNNCXtUQ2L5Xe9MmoOiA49b79Hznf/FoldFIB1YD
i5hZbGhsASWPK+kbHBPc2LFJ3Kk89gcdpws7p6AclGdFXakuk6pxOqsTEEPVhs8m
8PzknF52wIL+QYnVEFE/1mc7o7NbtnCZz4L2fv6BGctH5XWVLmvPTTMan7eZIFYR
29/wf1MKVdmo9NGcEnCyU+7Cm2kBSKLWy0Nly24C1PdUzzLNhK6FoIJPRv5Umt16
pJ748plwMWsZWHva1q0ZbBPT4L+Q49sHjdpDL+s2WiskRIwiY3dnEU437NqF803h
Vxj7yRSpJY+m+mm04pM43bBjuKqMsMcZ5fJbFGQs2qy9xQaYed/zeFJQ0+Lte/+g
LyGAdJmODfVkoNbsB45hf0NbZq9V8Naz+Rhc7IAKEGpcJJjRZ4uhzeeMYlp5aWLy
vOEgP00JmpoEq7z9pfW+ON6qyfzVWuzQ2yX3UbVXLo18nAAiGl3Ra3D+O6/LouJU
/+dnJAuv7zTDbhZVtqwlSM7ThnTCUT36qiF1AptAYiSXIFIzcBwsDP/17hIkDlfa
d+0QA2/F5tz72H97WEx9/WEnXwh//ZfWRD1sQXmPId4eRBnQLc5wAqEwqqpwztl3
RvfMnyATtNNKJJi+w9sYbZxyOo/Q6xRLYOY5pFw4f0k1oHQMLOzoumdCGphBLDCi
IiQ/W0PEKF+O+mar98c4L5VGHYzNQfdqXy4aNqbEPGCdx4nAXf4keAEhKYtED1gs
sEkw3/wDelhQcjd0Xy1cOr3k6vKoRcndazr1NiQ5FntTHRR/JNFZRqeZDvE7jFsy
RRg55U53puzHnsJG85yea8coed9qcchHnBN63nfq3UrR1qRuS5LCi/U+cUXYi4Tv
4PLluVoBlfTZllrqKFYryX+gL7UuFynSlqXuY9YTljp2aOTU+/3PzgaT/5R/oCAf
GDksD52Q5zU8Zx+QyEdZVok7mzoLM0ya9hRw6sAKS10BySa/5rHO8R+z36UDkfYY
0AYKl+QkyODrNxquaKDR5V8Q5ryRtkqo/Bzup50SxhDxFGwkqV1VJCyGfS3afDRH
RoHyxcFvsZgGdleGtQSiGWGyfgog894iHtSCkVd31kJq2ILktgyg2LgopVfhueY4
kyJzeuLNa4SqE1HF3DnjsnirBVuHez+UhlY4I5OPvYhGvIHoUYHYcLANVEainGS6
zyPSKWHkavNHVTa8wxcQWWpsoB5+S+hZszpNPAN/vSuUtNYEWL3DG0stiLaFGntG
33iZdmJYzCEIoJdyCk4L1gIk7Sz2mwOuGegIVfRdAQMNXpErE2+4oRMTSKqGCjA1
H/8NeioYln50JXEwkV7H3nFiIgt3/Aq+XeMR/EwF1WVIiwwK7BfpU173gDFJOyok
VYuFw0wUC7rNu6Imc2I5OX0n2sGqRqdT30UMIbfO1Q+gK4kngb9A9qmqXEVt6z2f
8yD3isM59HzBVjYeaTTHYmNT/imCMpfMLSXh92b/dtjugACVHspSxV/TEk1euRzf
20uo2aUkuDz8/R5EyLiRykW0J7LV6LNzasb9g+mgMCLMgrqfqUhqPJSIa2gMKpcu
nlFV8Jo7qhPy8zThC+GY3cdQQq+3OvCgxgAzKoZxFwi7EEK11ZXhbpolBW6O2bpV
N+TM4sOlTsRfIZSj1c+8eqYGH+UmuMHDBBL5hRsCBvMX+M6DNrm3EGgx9MYJcBxU
ZMMsU1CcVvSSO4dLPmlsjmf3ArI9IEQR7m2R/bejySx3JyYyOGu6OGOSOWBepDBK
FASnDDC6b5HkW3Sf5DJDj036vRX8g/YFhw215ShNHfBzsYtml3Eo0+rfSJuzZPwg
mWQaLSa5qHq21WwqV0Jb7c9pAda56dWPMYw5V4XLc4G7AczzI5o7m95czuKSQCeK
nBEyQGIkJSzWLWbUs7f3LvpYgXcuKZXSW/cv70d4NT+mwblM2j7fKuFXAM8A9Wjv
jOKXhS/2DoA3i02pguLGhnjRQAhsrm732ytIWcoD9F2KWQz9WagFol1TfMGFb+Md
kK+RsEY2LugBb7ZyeZxBvtjqiS84muw4z//Zh0W4Wx1Tqn6QMx2yad8Mc4sjdVr8
3dPgd3eWRQ3OhkqxeedF2SK8RL4ki3Ux/l4ns6qCzFkD+KB0VKzADPmbgH7/xSsv
8ox1CHCJT0QPm5PqnUnrqCgE+cmRIB2A9ABwJyI4hVMi8WsPJhTfTvjjp+iUHgQ6
vDiidqyA8lqESGiyws2YKloRinpq1CoJq0oSUNHx/E7o1KR0Ui/siwuLwN1+9GEE
ENv+P3NZrMHKAykqMMwJoy9a4TgRNJmTP4BuAPaJwAngiUndMygU6dAsqSkWPMPt
yEj0iQTMc3wmasu/leltxjnVlj1Ks36S8DfqP8BHhQndbWdeZ1Hxjzjg9YDR223i
nc0tYcPbezGmIVdhn1rmTIufN9sVULX1dg4V44jBP+7wzJ2HzTDiMihuO5BN+4+b
34NAn8R325h7bYKngCCXOjE5iGkNx5AhhiK4cAKlX29UngVMcVxJK4LceDInHos6
OsQ5NAqIpujQEw7IYBk1s656CZGfydv2MUb7wW8k7h5+14GlWWfTGzkNUac6bh/S
FXc9BGc9cfsHrzNXe9Ol0uetYZc5qXbwE458+9eqb8zfbWPrRGvAq3sO+GDIJGXl
h7XNQXuQVPi7hjRG2JCZowwDvTzThO86/eKVzZlDwZpsb1/ZlDh+f4Bi1gEE75Cv
AqwH6pA/48b6xmax7zofNIIHDp66yMv9luExqFuICrF/Tn286ks+Qw+k2iyDZdZR
pmzfpMoY6gQJhsrmIpXvLYIgrqxo8Ru8Db+b2dwh2w1oHs6PMeuPdROjmzFwA2zr
sdzy8leHdUPTQNXtacUg2/bakjkkhMZ+S8IlMrxUa6Vxi0ZTrlqX70CD4P6M7pMa
KjsajK7j+RZ3CWjphifVP3wPiRByRmtTJxTh209zsSm7lJ75YgEqu0e9QqGSvbJy
nTlhcSKdcxMpUlnay5de1CkPdZBU2onKHk+z80uXThD7h+gniAP0mSzNQfKCUX+c
OlFKDFbszxRnU5365TleGeQlYbbQnoBh3eMgM9S465qTEw/9ZZyUIa31fOiEeZpR
Csbn79B/mjZQChmNRXwHOHqKTy9z7/jbQnF694vYgNCS1/kLMSXVcutkqrXWaAXu
U5v+BlCsO84Gl7I5gkJ6irTZB0jvNyLfAHbZZo6Qba/bz3rXRBeHUHR8voOLuN6K
44l98MeLCTBnjObIbeMgX0+8AS6ur06ZEirsmFpAQTMa5SOzID3zvbjfza5yukK2
d673yLJUt78bMmBRdLBNdBPgqpyBfNrSkAMmn4km7eYKZuJTJ5BM4apzes8mRnzh
NZHKT8GucFfoz9F5VPnJtFhjv5IuAaLtL4JwjbRaHFo7AuFEoNUKMMsWM3UKLwvJ
5uoNV8L2T6hTGAZNukZdcG8sq+/LOiL9x+qHZTt4f6LiFjJBqPWDUD7oeQFANxMI
SrOxLwVrK63S6YIRYjpFz7lUNQW7YPS5NKQTfmoyA2SwvL9dCCFP7ItUd5mikvrx
jroS69GuK+zuMw9Rr67oVeIOAPhF2eEG79ij1X91ggimYJm3RWsY5gXYbY1MOb7z
nwXyCkWvBGlA+i8p1ybpdOdP0lKRlWhlWT80/xBJ122+T8LjdoOS6q3inrlmCmCR
FJlTlCEfLGJZVPDTb1LEA20Qr6KrtfzUyAFM+6tIRYBO+cL60Mgutl4wRr1M8cM0
uLRYLTNTlNzMJNBlTUSRtYAxzQBPpZEL9ydt55JWImqKOSM70mDUv2LCwwkCpjrt
8+xa4sKfdO4M37RTKJRobjBW8e79Tv3q02QTXGFcyO41yUXpMj+c2hfWld6j0uns
C3V3+CLXaRrTE3wF5rmdWVYZMtj2n9y3Le2Lh6KKxuMhPgn/YLSpFNOh9NDJRbQs
QRzAsoQxX2E5KuaJsDLqs3s3ZE3JOrGww+ghFMDKewA8YkpkTId+LmXlhSxwTsYR
H+ICw5ZX0xxZ0VpMr638GDRtJ1JOc2HFJdjJAhF+KwyvRlZ6stvNRiVShng/JjJC
W6Kb5WlTAaF2l4/6hIhUWUPFYRqkmuMmOb0P17e/KYUtYNW0ld2CqBSMvR3jnH95
dA2Pf3kRy/1nUakrba4vS+4qSpOdY4gK1Gx8SLvsjk/ngY2bb1/veGi8gEHSnnBn
Cu0SwZkLJgYihQkqiEVeS19WehwFDUqBm9HHSGMnkROyOJq/EH19L2oZ/1JAR8ib
8YleEytQ5G8DPn8nYQhD5JCXQHCeAZL9hRLgbBO6EKj3Pr/y5VbC+Cvzi69YZj0Q
kRvgNK1yUJMeL85EKpRpLi4oKC4h3qhoIS2HU+jalDhj3X8W4r2OMjFNtvB3CaeJ
j/J+BsaLlPVrF/NXD889RUf89M9J6Li50daqaY1+axtUTRCBh/z+44kXcKlP/8vT
Dqp7kYuCPMNumtkq4raSncxx8a8gJGCSFGebCQMGPiEk+4kI3Uc6RQGjPW6zS1PK
0lEQW92yibIaYfuq9XlG7VdYzl30iXMeG5bupMb978OlhYwls3eoah4xfemN6VP0
5TRKEcVtrir1+X0/Lvzv6s+cfkXBy3n/Cn9NAPDQirxiT5gODNL6A1hjTGbJ9mFD
X7RzWCTdjUTMODcpqhJX5JiLFuyG6MI4rwKTlF1Kj7fSLQVgE48TOWm65FWnFG2O
we+ykZNsBFRnce+w3kORdyAube7Yxz6kwxfb56ehCk1FGY0utpeRfgwZmrHfcYCr
crp0YLESR6IH6rwN4yXXa9kIMjKceXOLc4su2Ly67lPW2AgygLJAqYNcMXxFWLAO
Srh2fx3amyK0QeYvd6TMJn3QAS/e5lQasuy/C8E12YyVeC5p5VXP2KrbSTNDop3j
w6ZDgNHLhxaRpakX+7XIPKEs3vwLdI2LAWEuI983Csevmi9zJmY6pSshlOlN2ExY
7tGFCfI6R/WCtaEBYWugd3jNUJ/oj3V8L4S3GZfS9juXFgZPprMxJMv+a5lz9PQW
G5dkd0ByWcZLH+EBRHlpoI/bkNEbyy88J2j1klYfVXlIOkOcN1a2c5EKvVv/HHpy
u7JyhXPKCjUf8RP2Yu87ck7xlSy8+vt4eboGUA+BEfsWNWug31jEUD2wBYHhl1hL
OcgGuqtk6w70Zqngip3aFOp2aGUIFKfJjUXselwDcQZXyC93TU/ESS6K7buEhbts
XuG22hOU+2X0A7B9j2YVROnH3djfNTS+uMY5vamOR0GGiFQ435R4mw9yT3WVHoCQ
gZemyi8wOQEHcegmSgU+rosrJ15CeWMgGNmJNFMXgWmpcKErSBwfzAJEacfWUH55
79AydLl9VqJLX36prUx3ahhf96YvtGMlvSamhEFPYt1OEdcPjyw+oR7m3KQE4LHM
xJpgZ65fv0+wX6kP5N1n2X+yMVLbXYGS//eEOh440yp7kxRrudUX4Y47aoNb4m0j
SwZFU1eimro/1LCNpsGZQV1fwHNddIB5+iGv63XBBx/wOXrhljAEt221ZZVsIH6V
hmPmhICS7vMmGAU3B4vvpW9kYwf3TzLpknMadTpEWVxWkKN1r+PhiW85FSz/d6z4
aV8EB8aAwU5KgO5RfgtRw5kgIX0olIr/KiLd8u//s8pXSGy7bEugk4mS4y7xMgSp
qD9+UKEufIZLUhsdN3x0lTPqS1pW5r6sGkfrSMfqGyOAidelBADeEqXxfy4ZXqPm
JJTbDkbuDwHnSq8C6Bv8Zg8RDp1QNENrHpFYfx8E5cm3UfHJCCPHNt+t+LpzMTVt
o1xS8KU822Gdk/NqPj7AoIMke4+FeYGkTP0JWTHL/xnVrI89dPXaFUSkRzJsfv0f
NEmJCas7rZQ2iBYQXeJUQE/17uuuCi8Frer8XAA54aVWht9CnQ7alaRRV33wk9o+
nseQFc/WLhPwUfddEmauxW6FyjSzVZ1MEBRlJlf2t7pP26SxAN28fDsSg72H8BaI
M7iIQU7tF/4APEbwWm978daWYryqnlBj06iV3PT8eD7NXrmwn5IqClstQE1IkqC7
OUfnO0Ry1ZOMAMgFnWmtzUR/6P4vaHbPiTcsEX400e9a3BgCNBfrlPACrSqxE8pl
4cluGx2de6U+v7lWjSLPGfgcRaB9lu23QlABsdymgOxzgdFw4tZqePZ0UDBU5Gfd
efYCcJxjNRbtSBvcJ2Vq2OPW8mQIVuq0O5Zs8IwkqyF8C8N/nVlp6T6ujAYMbDQ9
dvcnMtowHrR0zd/uvuLWKAMZTdXBLmI3JESHh1aeQTekUsN/YFZ5lU4CdqcXs61Q
RaamojXyy2Twn33sg4BgSrs9DUzTHlU2S6xUftmooGiYRUHir1P7BxfHjoE7T/bY
ENv/dgPylt5+/yw+0p8BRaJr1NHuFlZNYkoVdkHjz49PpRozDo+jtFLDqv4hG1wO
H1KLlwT5DdzVghTYhKT6agulg8irFQK7pbcoHfmiQ+jJL1t3d56BdUJOFWtV9/R+
EPsffwNIeUxVdlL9ZPuuKrpCn2Od6y7ecxOyrKm3OG1mR4qgu+jsyiyyS2tMrVY3
c8Z1TTsHIFjMZEeL82Gxo/32IhgFkJc3WsfemlTPO/KKlWA4qccLqmVdZtYeMY+T
QqiJ7DdHgMB49k4Aklob3UVzL9xL0mr/V7lJ0mtnze9YiUtk9pZe1P2mDXo8p1D7
WhHinYX5FGXIzBiEQNasORQtXxIP17MYzdnwK4LmdmdB+XBZYLtydncRIKM1hEYq
Sf5B3cKUUb5CeyZvQ7pn7HQ77PwcGeHHmuaLFDrl3qKpAPWGHJ+5p+R+IebX/v6s
qs4r3i/ni9mIWqYzhOkfLIN4WNPLr9Xk+DIOBQLHGnEtIyxSyguQZXcptaW6am2M
FqksAFO68BqQ55Ov5HxTXvS/aEZaOLcgxJIBhdFB0b5DjJDVdh3HxDOyVBYrZhjz
qXUUt/bn3Suw/5Um2z7SLD8O+ZETNvN5n851Fya3VfKEIcLpeVKVgz4BlE0YxyIN
ODnXxsmczt8inmUHJ6itooi1DDh6K/xdYWoNiPtzu/ZUtgVe6z/bJTAeAVdSCXGN
ZFjkhYiSLNP8Hylrx7v2zv7DaLeGyXhOKsdQxP1oVGrQwq1WQswom+f3TSXdzy0o
iOs8VdKeIROro5hOhLuWR3Tbsg40RGPsUr+VF6M9TllWql+NoCebblkmrglYCfb6
e8Xs2e7ICLo8QDXCKHNAhDFARZN3Dv0zyQLi9fJkNqUYrDAPEkOL3Rm1ozelOCuH
2EPjqmhloJK94PSj9QPjRwCu/PDuGsOzVeRZuMeigmc240e+NZe4yqbFhqW4YWqJ
x7AWjluqIwYicgX6NnWxHknc8L0qkau/V2I1sk2nQIIMHFxdObSgEL4yhVf1rw9z
Sq0+ZVfnbVjFtlLc0l6nj26VbIZ3saCseIQ7/Nzyu1U4cr/W0o+Dzr97lsjF3kx8
1+iL5jF489GYvSLwLFiv96rdtifbw6pmca6S0C9Rlh34ynAStXrzsKeq7ThxuQTm
LDN5u8R3at57vefASvmTpeo7RkL9usXX3OUi/rfJjCMdcprTobwju66N52ebosip
yjaMJ2kR0Sn+yczfLekOz4uB+J1dBqKBpr/UZf2Ev0UrqLfvoCr7XjD/vQOlp0Vr
J2nOvHF9T7N/twUOKAh/eJc3XKr99xGDm/4v+2UMaGDN6eFPgHY8pol43tfAOL9R
RC3pgyFEhO+vGrI7EXXFZQOfBEp5aZEd00jF2qR8s59YovJe1DJphtPmv3D1jbr2
tDtaFwQl7+MJsvwOf2Q45M+sBi4/ZkjoEWejsT3iOMskoxKuKA3R902OglGV9LUs
DUbfh47ViPJIhhoAkzrNmf0OndVgy6e4imdABcxqkT9Iw8HZBGbGZj0fqAKPYAeB
PL/DqhLeTBT6cCol7342KIBKnv3UGwvaTyNt49pH5uTDIwTPVRpHFaXnAWohAyVG
WQQZXJq16s7LfJgxzIt5c08GBuM2TYKXbxm/NbjQA6uySfvnnNOuHENskTczTfQz
2/IYo8pILME/nEGNbBOwLadIXTRSiBpoiYZMk58/Hf1eHtooaWswNshjfodnFGih
M9rpynA3LXjGD1ZR9/Ri+Vta/CLd9OxP6k/bWTqRwsRDaxEZrdigL7uKV6JIqLVg
/0MH/tELiJmJbi4vZ6o9oScFi8dEhD0/RyVbLQIcfc4TKvEvdF0YKKzNytU4V3T+
G7mBTEG6JyL4IpZCta+NRlQfW9u0hLbtBQ2lg5cyahNe3+TDSyFoLD9TgQu89Nwu
ZhcAFUMREz/086PL5/uy5jn17cT7cazsqNM0mTFNwUZI3ad5gPdejL/aqkPP30Wd
MUk+azaqf/4HpD6yccBpSQYT80Nd+V5PjplCQ/ok5L6KQHavLyHjhwLuBgYM6Po1
Ktm8bxSwIbbe5XHfz1so5C7YrEM65lhKzQYVBGGc2ShVBv7wFIw0qeR8xOz7EGca
ghLeyrvssaIGWBdloPGmZzpbtx+vzervixkGPX8t3Mx3seV9u9Ot7kahD9Q0eWjC
KPyPkFVY1gXpKrO9qcbxM0A3Tn11PjgS0RJTZFHMh6o9DZuvx1IS2AxDoFtI/2TH
rrhgSN2DF1EN42K7eFmX3n9XL6iR0WzHB0VWGo7Js152MhiCWqtikTZ71rq7JPwL
772lXw+oQrENnMEgx7kzBMLqPruAJc7PjVRYulchPbkyMPGqAkOvX4WYNE5mfjxK
czjIn1T1IZTVB8uhEcsf32Rpy7m55V9wAIKgQ0VHK+aBNBBZsrE7hxjkpt1ORYmx
E481gnzQqt166ZVVYU/klCuRIOFiuTncMv++RGV6HpJZsvrruM04pVSo0MrYB+0w
/CDACbA5knx3eVpflNW3/63FKWs31gL7l6uPpwchMN3wBkHC2ITbWgtzm4FhqJaz
UkOSdHWRJtUiPs69jYPUoja9ztvJ42CyZkUU8IwxH3C2tlOiz/2l178sj6iPDFUg
SMzoRTyFKKLs5eopjjIuMdVadZ9WYDppo+7qVnoP/mRlPwzc2bE/ZsAnrN08ghq4
aCa5RJ+YreDUZ9p4JJDWlNaIkty7q2YVhMsqaeuQV4eBlL025UsmHVFIGY2TgleZ
pa0tCvUunzCXng72imQxCeO/Qp1vHp7buqV5cif0OQZfT5K8IaNDuZTLFMK75tFG
78IKg5AR5ovWPBNhlxz2tUp0JM4ndrVBprJzBeoNfPMyW4zArV2wb6+I9J/jGCkx
NjLtf50JDcNKs/nfzpjuwXsVMPOdzGF1mGnQoeEhy1oPg3T6dyV2TYD54fBe7gQP
ehmfvghYdmCWUwxydnUzlvGYPDzzT6fnYVkuu0OeRlx0WPcrTNXp1h2VyN6ZOZDu
gRb0FElOZXw+9RJ64SohUDJoM46qDMsE8kRa249mJZXW6evR08FAYWk9lxCmK4Qk
CCtjuu1pxSBiSDPoFQAX8Q7pgBW1Y30SDg9PQo3UXdoTYq0eDnDvmpLTu98UPgG0
huwaSEsnA6wKvsu0OzjUmSHozBRNpqRUnugtpepaSPm3AQVfQyPzE6EF9uyaPARS
86TyPB0PdzYISRTQvHcBl7jE4hRN0uET3KmJmiOI0xGcPI6OvX2h4lNJ4b/FcVy/
G5wJTE9wT4yY6zyXmf7LUcNKY7muZZm0I3D/NWxckM4hDuPesTqvULUMBuq16Gf7
+s4AGLQMLNK0kBtelU4B3q2K3Ne1s8l4siWg0u7H+2wCYIe9nA+PTUAIcL2fPCwH
sc7YLy/wKxnJcjcVgM1nNhkZBpVLWlSYtQ7Qpmz9FwhTQy6qxlmpd3OZzR0hhv6Z
4YSYYYwr4xBUJrIfeGuuBvLokpcdno0NcSIAUZ/v1yLULyO9zB+MypmCTjSQEWz0
JK1RA3EVcEZjDxoQgy4cb7EFz/H6X1gPpLuiG3dpqpUc3vnL7whwqwW/A+ni4pTp
eOh8rf8n7jRvIr5E09urVoFYphZ+dgJIiiNVxu6Kb3/PXwmkdBVfWLE27RFSpB2A
NO52m/eJ4/b/Qx8NzUy++eRzkheHuC+mhBSQ2L2o+z25BzUJ3BjQOoOVtr7CCJT9
6hgR3sn+/MptE8z0GHHV0uzOM/HoZpJIdgH0q7hYt3Kib2c+DbnsMmw9wSKW9gzM
kUejKlHQutGCf7fZ40zADqN2YCvt1xMsuGrj2R4xD9UNEtcosCeD0nFrXCI7EIpl
4jXVx7Zv0kpYSfE0iwBUMuSowQUfUbKLyVT2BLAcP7lGGtGPEMOg6dYMNp7v08Jj
a9+TEcy9zDePyusZRo3/hkAR6+rnZmg0gTurBDOC1Ivxlb4lZEgryN0fP37AJgiP
2edyoJo5fWeVAxWAZ5xE3hC5L0AnAAtBu5bfKBP4qmrlQh/PM+WpaLgaodwxE1C0
vmW8D7qox6AhluEcfB4R8FReCvcpeq4f+25az2/QGwCWUS8rx9lWaePauFm0L5ME
coDgxF2wr02ogGCuyOOkQFTNS2YAm66ZIN7vAacepAxF+5UBRO5qx5/4gS+3HgSO
Mmlw9np2aW7RcxiUy5/7GUEY4/eYJ5iI6/bW8oHkIloVHz3eRtkBOv4/i7iepeeo
2AGGA5Dp0r7Wwg35tOz4GLcR1u329ct8EjlQrdC1nZMXqJNcJ9crFkZcNB3jspmF
lskxC31h9iLymWSkA+VUwmne61G8kpYSec3C0lr5G+R/JrJC9PogtzIRNHHQSVuA
wuubalgnGqsF+xjnOSHvooCrEf2u4J+RwdG1Rh580hXQsjqiTZSUUm/qr6aW5s0q
ScIO/M00HbzMbbLhmtmC9kfByGTTxR+n9+nG4IUJhGD3+MLLUbsY1UDTb/x42lXI
1hVAwXAdxH49qOeu1uuZqAtLwNuD2K5+DftFDG9gY9hKMe3EkaVh5ihwczjlrOBV
ummyfd5qGxthl3LeDvR31ybxOO6PCAQIfYVD+r+au3i+FbFIDCNlmfxjYuWsPvyv
8pK9X05d6+cQ3LCRuZfjgP1Z6n0SPPZN0F5riwWoQ/nMTfAKs740/SxutHpyoA8e
jg3N7/7Y+PpO7dX8AKunumCGQt/N2ibocR3yxKfHh+rX02TJJuyXn2BWP6MXy85l
7LqWoPwT2yB/Q7al99thylG+5AAZdmUad0KWcGZa3h5uNPS4ElaW9y13/ZjTMZ6N
glTceRP/kqS8Ea4+Ed14jmnHEcZUNNGytotCOWmsj2HCGAgGDNTyBKF4FCajZ+AL
GQrRgPFP/VSYa1SFjF7IzydK5e9Js4kUHl56VQOGY1hAw4jHg+QDCcUBL+dIU9Gx
dhXy5YX9VpLWmXHfD0VYyFvh/hlk6KZdCPKomJmRFnIvHOxjfLBcLpGye3yL8g9v
VlvMq9BAvidtG9yLMH9UHRwLxeQgTb7aSZgqm8RCaEyJZyWOwzRsYY0lx007/jQ6
A3SdNffDZlMbZktrRsLlcPekFJYJRmM2MUa5gacogIWPXUHWXEbTk6kBEyDIRS4J
/OhSJqWiS8xrnjDlWByBDA==
//pragma protect end_data_block
//pragma protect digest_block
RHB6KSnNPLdmVLmuPiMwQIXLeUU=
//pragma protect end_digest_block
//pragma protect end_protected
