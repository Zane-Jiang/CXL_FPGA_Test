// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0yAwgdUO2dCgQAtCki1eqv1BpBXNq5hKoGqxdYs4eMnY4kSXW2Wdq37WLckB
zHXn2zSToKifaRXQbZP0owbWLPwGFuw5R6r7u/UXCH907ujoKrHOqDsgNEOS
OqoMq7SwfVlZ3qHbHGe5bnCYBXcL4wHFh1Jhr5aQ4KEnmkFGvNLuzaZK4oWm
REYiiNX1+4/3bQgnZrRqCxRHursU3m6fGh0M8oy3t3S5FkyT+jGWgUCXaslz
TiAjvgtAiND++RVSTA9Hb4j9ok/hjBD4Kxt3F/SsOiEYsu+mdxwZ1zjN8Rnt
6gNneX2SC/6hR5E0C92ArQWNMYvemtaP/t8610BkZg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LOzXWmFlP/4LcVfgPvbCblZQokfmofhxR/VfPw1onFhzjZg0UaDg2c7P0QY4
hE2SpE4i1UHsPk2ezZE9n9+fhJOqrUm473y6QopYsTFaJc61+3yAzugS0JMX
53AsBKDSsB/QYJYMwJyMat57S3jg0CMoamD8v/ET9uRBiX1IsCA5LR5aVf62
IuDmn+Cv/tC++d4XRkz8KgnA79wEWFSdQmQ8TCagRRe+ziTWqzgZGByDZqpS
t5/KYIEP6COCwH9zt/+YZfsDc+/yNoMXDuoFT1SsHYnc9F8PCMGWg+iciaRj
WDHrWEoGxmLORMTYXHGCdkGn2R5fU38Rc3Df753TJA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LGjKg3YdrNADNnSSVr07PeNbX3CwG27t/YG2xPpmFziYtiAlyU+tGOpNKq4R
0bzDgW/vnB0zh6t44phYVCKcZRI9o+YBFc0NaSg4CpPLr86CCXYXNx1eMKZg
DSEUE7Us3HZ8PbfZWzb0wZOgdSEfJPIg6GKl5C+JwKXjQvAw1CG7He0qY1fe
2GhbwKzpUWQUXshtP6HRK42C7NlxCzZg4ZfdN+2uRuJkS7jhOExJd3/sP1Hj
SEVJfUFETpjZIPUVvyj3N4Y5m7kDz6eg+qcfZKR4gNdGYoFdL+zQ/NGR8cl0
Yiep02jWbzlcwkudFHMILOk9vvdKbBwSrSRcp4hYAg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RE1fc4S+sxZK3XivQ4jffbBpbUrmhp+eeOrkN6FUuDrKfHXgm6DSoRS/buEt
OosLhBm3lvPtlaJXcq7zNkqHgW5mgTPwsCMPq3tCrNsyh/HXx+fW2kFKLjMW
2L7YEVZCeFhq8VnY8wUg7xZzmHA94aJtFtwZmhOcakMqVw8ltfo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
tfxYc2JFXlKb2PzweU8tMsH0wae/UEyMLdV3G0mU3RrD9vkeoCbZD8/zn+yA
cSEjA/VitUUT8ju2/RrRgLu5sMZlE+meDmxm5iw1der3UoruwMbiaKf1x2Do
NjGKlMFdtSBTWiq9oAM2Q6tMJJ1diK14j3u25U8ediYaSJwg7+3GuL8FAmc6
Dc5DWMbHokAzS7rH/97VVvvc46qCBxIkzjGDoaJpvTbr5F9+noKTvVWfXB5b
sTJ6/nBpeeypdIZ4ev62aZRutQc7ZAm8zm50GVFJ6UCJRPOF/l9srVT4qs5G
Mx7poIAmUY7cnOG12v4u32g4xi49T/PxRDcOpfE2LZX60Ec47rha6BV6c6Aw
khFzcdgvE/j31hb0NML022Fs9nYYo/+/fk76TBbhvzoxjUdz70ya8k/ceLh5
64oHJMx8QkWQn7Vbfu5ede3aeujk7RGsOWw61j0KyXiJ5sKap1+5xmbrawH3
KoiaJmLEWuJM0ejR6qkqP7cwtbwRu8AN


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
upBr5kqPSmyMVIEYETeZYrR7x0qRrcYJsIwew/5QG2e5AqviwJh1ixCfjRL5
nOo2//OhRT9u2A3UUZVbMwG8Dc8ZOvTzO1aiqnJ3cEv5IJDBIb93sTMHBU20
Pu79wqoXC2JpHTjKG4Q+3siUi7EyeNLZoGbTBd21Qr7CiMMndZ0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yk754kXsayvdssvQvWNtyycJrGhY7/bITFBiuR89WjoKZdYx0eDSXTc/hVrO
bDoFIMR3cTYI+0MyxftY8yTGzghRaPWk+nyfED+XOyDT1ypW1moMi/uX8vwf
h0O+w0RiGK/d0j3RkPwQiUP+xMcOCIEYCDRddwzoEukfxC9aBf0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 150944)
`pragma protect data_block
piVkxn+5DgMzJ+F9OBAeiIjBp9GhXKacft15QPPd4+sFRPM7Zt3zWDMF8wGJ
Ze40HltscG7kaLCYnlFVAL4ruPIslrL59lCWT2vcYttjR53OmZ998IdtNTfz
T0IU/MjwTJClEURdzJAoWuWy+6HuX1xlsAQNE18PS1ZaZL40lsx6BddUfwGk
dI0oE/WyKvq+uWJkbSdD95UN0DpZA0VSUOGaYOKoNZObAsioN9fzry1vw+gW
swj8tK0Fk6Jz01nIwAqerI0zsgXUX4rWqY9UOhQMQOpIruc/OYOy0jEkdS4L
fjJMdVzbRmF7w6sLC4BiZYAgvZTI9MkvSSpbJwlp0RpJedDdV4qA3x/3OCCH
Pe1hpBON/wnwztTAKH9ljFqF1TmzzfQq7kpGg1/FGHmhq5RFOM/Z43EMDUjv
o3dpGjZXcWNKNrmxNXVu7MHC1rC+/QCcEdxaj1pZpWi1e2BpnrV06Wh2PLhD
+dqFrTocLgvYns2QI0mOI8u2c4zGYpeg9S6pXwvrfr/Vhfcm1j1aojptsKV2
wNi429pNiI9L3kshkJzn1m4Rnz+27VaPLvgfqH7FuV7RnXT2+t+jlX9vMV1s
9/JElB4LS43y/MH+Bu14x8lwCi8GsmDi+/vZ8M19kugcWl/UpGb6EBcb0TaE
2uflRrLgfVxYESM11k3FvV6/ENuC5mwAQfDhtqVTK8SMQlx3hYnXA7K/SE0r
4yFKBzhGcuOYQi+WmtDZtM0WncnVzvbIlHeYZL+iQnT5cwQjNdtD0nWyVefH
2i3k3zic78fMjlplJj1RKGkv+qgD2r32GUTbSQBAEk6L9gCdisfnbbvrR32S
qVFzX/YUqTAfgF3rOtYU/t2IuNAJhmBZ24w8oRPyaSd8Z2FXvNdabVM86CW5
axT1Kuj2URbBoq4eW9vMShn0F+ZIOvSaUhi5POvNZhg2OiOKqODBT7pnpJTV
sM66XGp/zDw27by25ydG+d7iVXr6TTKixNSBh5cgsXP/7aRyrMPgiGHb9ezR
Prg21rJ2xy2wPokhELJbpMbm4no4GpPPJRbqiSLDG0WbEbw5wsaf/JZDu8Bi
JN1ZqaKMMcsRxWRucIpnXFV+aFaAT9bojcSbMgiFCqqLiqvBYq7L+OXDrH5D
1zUITprH4Gr0yH+PmL8McYI0jwY4IhDltBPzpYsrbn9XoMug79d6eJZRNKKY
HuOi31LRHMeQ+QsNyUWItEDQv5rYOWRZI/5GlKE3m0RyJIR5j/d4BgfsqrTw
vEswb0nrdQ6rQ9dYll6fQBzutEZgLmVuR2f0KiXd5RFRrKR0QinqiGqirXW6
+O8rDGb3rAna+kpUwVzwNsVjL5dHyLl9QgVOLSfnkJEei2sv+KJjdWZ7WmsA
gso6qeTZazs4dLyZHmvgShJbAGT1m2xPE5r3VPzpnzOZwWFsqxZDZAnM8rx0
dqPl+7HRxDpA2XD6kXDZdvsR3Bs0ppgxZCbpqPEo1IRJMJBaIhxcD4WViT1+
c2R3Nwo4CsL8InpDSIwAqEFhnSvBmCHFXOUo0Ftis2gsAkU5tE7rHwmE8d/f
EZzEN8wBuZ+cMPWc0w5lT/CGReD41jODtTA05LhxMnjDskM161SqgfUr6ETB
1jK5er2ChBy4AMrFc5UDiyJD0Bw8Z2HNFeRjBZYGFEMxX9EY/A4yKQj36W24
1kqYrR9uPhw9HZ710sYIKwLvNoL9mBZlyGLcE0st+kQ4yVtYgVVmQ+rjLwHp
LHAq+lPk9zWRW6sHRLZ+TZeg8ak/jR4BEraqI7ty+WI1FVaLRmVE6EKDxfp3
TdwhBfh3wVvAB0gOmflSACLVqfzhmwLQhYJrsy6ZUbU4V9wJmZ+HvD8+chiJ
kOPWeTqIIofH1QeiIJrzqy+XPUDuTiFM5h4kHa4APUVzeKGpCrgNGjYnuIVk
XgPYneU1SOrK0lldTUjL60bQgZazVCvlXDp4m+7smFGQRDWLVWTH/gVyrTRx
BGX3gPBNLcMDQZBXr+pGQGu458llgo+dkDAXN5XmQbO5XYe4+qRknL2jv2k7
C+9ZEp1I2N/5SUGOOK02FzxD38nRImK2phTabDg8mVC1TyOTmuCE+EHWnq1M
qSZ+4jRlM5955esBDAaQq0UNYHkOIJLTxjlIv6/0hKUcRoGyTrNXXeNKYg/1
/Srd3MLDXzMX9OV3QW5nLc4519OdZmWBd7MWnjrV0hufsicLwlH8XGePDer/
4XOx5bMu/pCJ3gjPXmu75uXDQBS2lw/BCdfgqwNdZV4zl6o5YbUON0ELqGe/
UJQJP8c1GHXGLJlih48jDlQbLEV8yE0qkxwjAoLhHIZSUlDO352CQbjySN6e
6DXCKVpfVLVe6Q9epfae0sTnkGv3pKpoAuPt43SfBvictBfoWPiOIlUBa+36
R+Ui6zHHmRRr6C0vlkuO/g7Kzd8gUS6q5I7AlJqCa5gBoZ2jJdK8PTisma+j
Qt2n/BWRD92E097iJOySO7UIDQYIiRWcikiCHdepA5IciuOMxKrnAnUXqR1N
Ca7/VDsSu0WLbrTifraFZBaemXAqQBSW1L/FjyKiciG//caxsfj8Z7tWxRo2
MCg8ACyig0U0OjNrepuHMIjz7zg2EXV+laSUMZwndA/85qLappqQJeEaFnVl
91oLpRBZ+GZpGxU+IaiB8JB9qONm6FiRFbrljO3ZO/oiuwh7CdVsIZChfTr3
StxgIUE76+O3S3cJNbEi1MAi/qUuNmfoTnsDKCHZ/6ObmIqZeWuWOhucZ38t
qL5IRygzyee6eXUQgge1gqDe5lH0Yt7qT7IbPM0GvzD0stou1+cqkKPUfTQM
995RX/utf9VDSWd7FBVI/Ewvsf6xjIAYP6qqv/FOpzrVr0oDJbMvxT3Zush1
QIYU/nVRFbP5ATmAxA3atNWq/ZTrHHRnlMRpL6HOdVHmDsnSS5e3DDA+4v8A
Z2+8shxCiIxTSwWXj/CZnlr5U7fBJOYew9bp4dmcBGsXLh7GG3TOWjNXhs0r
lwIL29rJi9nJab5O/JA4RoEFNpfy9kRTOsmljQXFO3VbpAf/o9d+iyjpNUu2
F3g/Qnpr674OKheG6vLihMJhc5Za93K1RCknxpKm21leTnxnreprWTrWVUCT
gZ75jlDu7Jw9QG+92DY59TQhyonxzqEi0Eqfsu9bgq7mqnmWOPKJuhVbs2Vd
hNOjLszqOTKDhK64n/ibzwI5bACO0aR/WAUY0Bzm42/I7u5NNRAgyLtN7Swo
TR/ecEiwyEvEeFm7ZCwBQrrfLW2FHXq4/ZSh1cK/leftMNYIe5YNEzNeamjs
BVcb+hiuRMM8LNVF8YCtedU8HGF5vo4NrqwuE8IU7UA+2bMiY99CrFAzgVZS
w4EB63BIl1TbaKzg8aEpW22SEO4EICpcMmgFcxWlX4go+I/DxpiU7tbvAvMw
a/GYx186Fdi6mSM+3zkb0LSZ6Spy8d0fAeHClN8D/t1mGxJfkMpeku+iuupO
yA1v2OypGFnHdWJyyhZwW6BtZ2Jioa29DBp+XdvxXN6PTB9i7nkGzVU07eOz
l8+whiSZBsZ22Q9Ok5glL0RZCY/Mga+84esBVLx4XZ1FfqWEfkLoovTDE6Ez
yoiod+Ud2G47oi4ZcKJHfsTNNzbnDA+7NOpulTDlKKVSQ+XuLmCayXr9tSVa
082d+zfIA7GDG+r7APkNDrJ53zPOAqmFJPs7guVGJGrHavbk/HUcdPYhCdnx
2aGSx1UqZplnHE08c0aXkLXZeSCqpIRcYjUOr9MudW1LKjNUv+EesXUPaS+W
N2VqafNREzu9TBJfIIQyLuFmIrECaW3J4q+LgilguI2wZFQR1QKU+DvdRpVP
/eRWOHkbDENm7ySE4GNgRwQwWEIY2wQ0XPDxSr756n4os6cHUHMDgv/qFAWJ
aPCK+GmZ/mJf5QCXAQvH1MGH7OK/PGTkMSZFCyh7aNPDO5pHsG0elQ0jbUk4
MAicJvwlYvY+ARTd/mULR8RwyL5+o/Xfgll0/RU0Rkul8uPGVJUpTSu3S/ru
9z1pZnUbD8tSNCJp8m5Zum7ICsv2zkZrNoFc2+gdOC7e+qxUZjV04MfWGLOt
qPhlzNnNFHn6pbnc9ONmTjAr/JtDecjrj6OwXG14zzu56O1sSRP5yH620ADX
Qp8sFGof91U2/NJPdDNgiwt332bmaYJsicMeJyQaOXA4YzhPRlnawYApyptF
2M+pe5LlR2VJimhmrgIdDZLG96OPe0RSYgvUHrSqREQffbikuzPH68oJ9AF8
sP/ct+YIQyF306QfD2f1nad9Q3pqEsQ7kMLqB9a0oHEWAzpK/YaI0R/gSVbI
Sd4INXKfkm5/wez6i/5XI5gqy+ZQegxzq/XF13pQI6BYSej7pJSSodi4Q+ho
pLenpsvYWZWLnPgc+pPyfrDVQpUNg/3/epTrsBICddRAZ4ksqEi3D2WMHqYq
5y8URmoQGvJQZwJv3uPt9dnGPb43pRheaOp9diWdzEkepXCWW7EtBMxIgyas
S0R+90ejppUopGIzMTyp90R4WIvO7av6JFwUIBgdQKzQKc8mUzfoAwMRFonz
xQtbRFuUMNKAMXJFU89wRIlaVQq8aFxg2RIPCUxOp5/TSPN1L3b0iQDDY3i1
1AbmF5xAM+3P15yXvp+wNjpKTP8r2USQJLYQzKwTGMrShLPK76OW0TWa/4wB
wBCPBGnYpBkGMlR08E86KrFlDFmdeTxU+AdBuZ8Myw0c3ZVgHQBmlqd7a/gh
XNUPN3blNWbVivEfXu9dFCCYF88FNmt1IrNXs3jnf5zSwM7qNpMKTSRiEPey
F2dLmRnmKIsylahUfB4tsq9Da+dBl1qknWMzqeoK5+7B1R9y0MMguFWMYiwj
Pdz7ZQjKxcN63luJlbEaFheJ0L1PsPVwg8crxRyT6llmpFHnmKrrSxjXmv2K
oJk/1gWQFy2GElHmkbeqZ5Z/BjuQSjnsCX/25/JRpjps1b23xRXUuvKj1lPM
KGr86WH+SW5i26XuNkDLlFb9Y1rVB67QrPTzFHNW9IBgE00XjCXrtrurhweV
Xt7aYE3JxOM8t6HxmyYok+Ng26eSy0iRK9QUPEFb/2dMI5hkOZtpYSM7+NnC
MGh4HVDtakGfbZTuiltV7QS0AbQNoOHDNO6nmGaD5YeK6kfaa/EcorrQd1oJ
1/EngL6n3J6MfoZOa5MkLagiHYYiV93X0JvycpmhJzyjByEY3JPlYmrBJhUN
cM5hx5yqJ5wwBDadyd9WS+VsfJ/yLC7+3mvaB3PtICD3pQY75JkSJisMZ4q5
yBYbn70azU4z38feFIDpsogYPzEu/Mj/IGRbFnZxsTgnxD46LQD/10VtVtPz
IP2jARUsJg49XoO2fwDKqdIylAjx/kiAmAwqP7/jEbSf3Hl3b0oIS+ElSWVG
JIukalhSJga+tS/GtwzQSX3Fnlgcc1iTWCVj9FeyIMuMoegxiBBoKStkhpqg
rX8np242+OCaqPN9zBVXb/tK8zBevpL3/MFVZPsOqx2Nd8AnNIOTmKHgCM5X
OXKRRkarL3c+o4aWONeVhs/h1AsY60pVsWJ/zEo0OFH7nwrjSoBmQzsux4uF
WXM9/YmtlzbBZQ/l3Lz4gsu2FWP67UUcQfR8kVNpPFknU717G6gKiYULl2/y
bZph0UQUEfBWJv0qyomEJh8UnLA35VzoAn0BJCYx5JAAlu/aTNqxtPXSCHki
u+ymeOSilV5slWl3HEdj7jp2DCz2cFI/P5FWmt65CvM7HrPHdJ4J8qFhBRIF
yC+uJ4tWVKYF0ryvjLtem+negw436K/LGOJwSULZ010kFyyCN8hfMNGRY7A4
DddcEv1CPuk1Et+e5aEgufzWUWQVhlURWJhJOaLljAZ5R18h7s0R8vynKfvt
93m2QOwGgX5rwrERFlYvSpIT0jhqdsMIdMCxLiDVluWCSt6+MrH32duri11K
PhD83LA7R0sBZo8Jwasw3A6yDuMw21MIexwm4BVNZDHTBnZGYuh5L48X+PJB
M8aCnTtF8qAu5yHkPQzU4H2vUUZ/RcMBlMGt4LYcJqo09cAK5yY1wIGV4MSB
d2urX654scbdGPt3yuytbuhI0i71jA/wgTsIRczPQ2kzoR6j02N0tcqTNi1X
EQT8zH3yHrYXslHl9oV5MlwbyMJtL9cu6UhKW0xeBvGQsEZGmcqRY917/V0v
uCiPl1oOG0e5GyljWrKsjZ+Ljm0aMOZgSFMmXx4ssiIiH/aa/bM7MH64ZH3j
jndMnyqURRB3MiYms0j2i9Wov31JaBcdUl1/8nbNGGPlU+XxqyiB2awiBsqc
n18nL1v6gFZQxHowPm+XtCqrQsG7nDosydAeACAV24ez3Piva1vV21GkbIxl
lCsEsAL4KgVqsrE4Q3VcCPIpIDYLsPa/7AcrchNJPZNZDFGJf28M9Pv5DqvG
KtxvtnwK/G1ocoyIzKfls3OgKXaa0vErly4n8tPIKxJtczjYQ0ALD/cM7huH
3a+FU97L2AaWmFTZFr8Cxxth6DaLKY2NaeBGKzdMXtMtUr6OKZfi109I/8uh
J9oGtNhazx15kueiXuSBoFZLY9++a/7C9WGYeObE56I3ymnMVadxV0CToCKi
YUd6Sz9TlQBF5yVcmg42AH4NDnBkeBv8LU2WGQhTBWqE4JnRgFbeVY4mr9wu
Vqv/44FbkyDiYLlbJ9uNw34q0UqPSFHDVmVn8Zu8j0v8MWt3oxkMKLU4UzLp
x7qjrJYmBY0qcBjori2zwlLYzH8DSJPdwjoXFXKDwe95PB64Eg4oQGcWJ6Lq
kmweJKwM0e8tD6NqL4RbjWE8bTxRGU6g9phycQIg7xqbIsTzRcyvuM2eOQqt
z6X8Q/K22w15fwiL3ei43VNLef4QVD2IGdGqu9BG540nTSkHM0YOObiOc1JG
My53VQFYyW6KI0nrqAG23a3Qrh30ZFMtdQDrtdLuB2UxD3OUI0yX0YLIGUk2
o9Mj27H5U1Bt6LnI4t9b7QC38ivXQjwdN5cTmbI3+XQ/FRCxDGlv3/WO35q1
Pyxhbw7ugIB7JFkVofoJP6pZZsYr070FZUbnjp7augvaIkgE3my7KQvCaexW
43BBTfuLzI1qE9khLAMY07YLJkzeyv423i+62S3WIXZm7eYfL2QlpL+uxxUf
7hOg9xElA4xsOEixo/KxAB0VciBHVBas4J3bC0tu+X8saDhS3c8LaMSil50Z
s0umqt94wQgyflV82XrDQ0GFQt7+xZLW95faPtK0ONDi74MIEAT6i75TAf3a
E3G3+ryV4a8GimbP8cSOM7SNySz6tWHw9zm9NY8yaLlToISgwaA6vNuCmGw3
9yiRL4TtvzHwgELFS0qre9rQx67XYAnJ1YntLYB13YMx0KdiuDXYkyP01EAw
qnH4CZLUleB737+9n2KPHFjxSWvPBzAgizVdZ1hwLlXWesNNFz887gETFc5Z
x8GvC3gXDFqNcqB1qeA8NX+efRNoqZ0VyS57ji8SUPtPKWoYX8hP+Avibe2E
Nn9INvJG8lLUXek/h9qT/doD3n+5OxUmU0GtV1VPqzco/8uuV4XAVajpGau9
EuD8Dj/2dhpqEfQnl6T31bc6+pW2QG/LrNt1iXe9j16L01efNzzahFH5riEv
/IWJcQihXFtx6/l2bNbYrELUHlMJ2Yr1GtkWZ1UoYkIgrHPT9JztgRCDsR0+
+MMF+JPUKV2Ie5eDu1SjiI39CZIgloA5E3+ypCcy/4t6r6E0iaEqjIUAdKPr
TyzJd8PtJ56rHmHH369H20N8vW3WTQkDjjXAEuBi6yec84PKQFz+WxzLHHc0
dXGZjRGCbXn1C5+lf0xY+gp6Ws8pkaygGjKBxK7xarynb3g35TsDXuxHGgyW
ySWath+wdoByb/wJikTNz0vPZBaoWxagZu5uvnfSFfmIhxFGOpUZTccTkFjR
blsXu4MnoCGMxWCNefNtLlS6ja5xvXn8joAohjvH+thyIBlieX9Idbqyn0+r
ULGB+t6VG75E2QooToxMS1VTRN1qpaRkj0QkEEQ3UAtzYfOP50fnpJQkBf0s
vAa6tySkMjIMGuEoUpBWtzGij7O2kShE2B3FFC+ySjHUujiXGbtV6AZaqCKy
rEAWTtY8XP9m3X0St6b7be2SJ/pnsG/RYuV4CfeurGiJa2qc6SUAzyjjkvm7
f3Gob3ocOoeSKKzAhyq6My2NHKRVLIOMQr2nlFSyoduDIaMtLTboy8XUH4uw
//1dmTGipiDLoKr2UhUQ1qsxyY+xindziz1OQqkm62adF56q5ePOTDYIX6NM
2iagXuMuoOtD62B1KF6EEIat8zpzIQ3hBUlq0g2bY+7SF1ddVrAWXQa1QLRK
ZRJbKTW5Ah4BJ+2MtlySoLi/Aww1RDHmLs8Ii63EPMfVzwHROqVbFMRGbrvn
25KcVvZgNkEvyrbbLV8+/px0tWGArBGFtzb2YNl9NPyLSy46II/EoQFKn0YO
X5uoMojj5jT58WNE0PMgoWuxyqpsIUUSblsCYRr8FDMmk2gkULltWrZOLbm3
6SZ+W57QcQo59OPqKqmCMQMnfm4f1QVl/sI6Q/rVV1iumY2RzJemO+EgIGVg
iJBURV+j2jT/PhtsPcqTxU7iXyhLIkaLqHbe8BeOrxUbcP9OPJum1beAi2Pg
qZUcRTZ7UF90QzFh4waS8yF/sTzqCnuQGULvukElMt6KNJRFWuLj8RprmFAe
KHp40WGyE0objkYWYZnfIV7++cjRIU/Epbp8hHaonHoRrCyc9QW59iEloqJW
I5W1CNZF9KPuSv9HmeSkaajhr9xOkt55k2iDE72JB6zmxqWXodQH5qY3cDfo
rYG6KMde5XouCijp4c1xXtbyE0ZeJA9qSA5+qeIEWj9DkfL4UKr4rsHt0Cnc
JgLO7hKYyLwyBlbOixZ2BnYzkjSF6LVZyubu5or4/7yG3DgTGYwcW7ieLg2F
vu68M/ne+vv+JRfja4TOYdy3UoWgphtbCYRM1hDZh1tn3o0eIjOFD7yxculO
szUETsCWOZtVckqPC9v5BjsfnNcd8Q+Ih/Ryg8QKaNBmfJyGeYWs8OHKA7c4
mzD93/8+v+rcqn6SE7obgFD+d9e3TWSqVtZYOLYAcQURB/hzFFcOkQMatOnK
xQsJOBI7xi3Ppx/rGIQzHiBzMg/tjPODWa88sj3+Rs2Qn0CfjK2QXQDEJeFC
2ZdYnODRft6ql9fnvsvHU9YYFpMzaN8kZpAzOYwhYb2Hqgv7AfqtozCReMS6
7ucLRz93yjmAv/JL/J0XQoJIi7VGj5FVnxJVbhLTtM37n+4UXxy5WCJ9YS0j
ki9LjaaHnUmzN+t6vQSAk8AQ+mn4iccwEkSr89qTaZsOaT6Oe1/IEqGHzfpO
FZBQ2FGjGplXeDc2zMoC3NXAyk8vH/tSuQDvFcVT0v5CXO/aWU72gmFuVGa5
VYR5uI3D/tXjN0OLpSjwfD66l8f788gs5N0dzIAnpUIBi+3kKrHkumjM9ZFl
PCQ3GfFIx6RtMuYZQDzd7wannp1iYip/fUHK3WWet9XDpWjyZw4xV6Cp1O76
5spqYoofCKSMCe26gfo3wVxPzO9tuXSmg+di47F0n3hIuiekCBigzR8fBzh9
jklewfhriELUIseTGmLifd7BVm+t+Cu0p6WkhF6q3TrX+aUmHZ0s7iI4FVki
PrkDVUjZTOA5fjXsUsPT4PBNQJ8jpBFR5Kg2V/rGk+vUWzU0nsc/kJ6P27xV
Wa8B7iE9bKjVo36vgmKehzmA8YuZthghHQkJTv+6ZHm7fJqQd0/2VFNk28s0
NigNEEpN0C+CB61fA+63xiGPwTLrcX6An8j2vuKjv456D0SXfywvV28XkD1V
HobnwonDIr/y8gasKMJruedvGMF4RVDjWZ6iuPtUBkoUtE62fKwbvBoOQuZ7
L2Q3CS6+nipvwiZVLX0pydrcin/UY/xmIGVx9YdflVjEmW5FLqE3eJiY6msu
5Jgj05931D4zFqM9XuksZ7FrZp3wI1XA8G1gkZs6EIu7ijFtV7gINICQJbik
qTzLYlVDGlXR9wsy6LbRD09U8KDDEwfb0lRZRWkec5a+JIZb0oex/wY9GWxN
s6mvK3SzRNZbxUofc8sQVezWQ8b5m/J/UuVwiCPlcBHJo/JrIc9SGYLKfLUS
qYqtoGX5FubLYiB1k/TB6H7Ip7P8wevU8xMjr2cjd/j0m0RyI+L5hXs6sT1N
epuVk8Hz4FtLasZSzx9WTpzWLsadbBUw69qCUEHo3rKRe4gXNZEyR8RSuk/H
OfAAgp3xFm+AQi5XoGE6etdYAHqV1PqD9c3DpyaCTHTyLHs73G+HDyk6FQti
4GQBA9RhytQD8iF5RTLtVNoP3rJLSE5LhRxA7B6iFCmPhioZlZmDwbNrancD
th0/7TUlVS/x1m5MmGkGLT8kCjSEs90r/qzNkfKSsPhaMMGhY3S4JF26hghJ
E7zPe90WgyXXguTJVXNFny3AQ3sYozq4+/LsoRnATvKCa7iVGNd3y59WrOlu
LdzOEYj+0ZuYptTz0Kxm8NYilCBxHkveOL6IeyObm/KPeBNAGvQs4X2dBdxy
zF5KTZPSRpO2G+0t4omtViDMypvBpfwnjKLKh9PCio9i+BDdNFC1AI/e7qrE
SeDZIvk2k0VAYRPSbpusPyCptGvwAsHb8kT80KX3gQBBvD9Ur0GWXG7MuzHN
HT8PvdzP2Y1HTBB8xVG/KuwKJ/5DrE6+fHsPruOVRfVMGOeI1+hVEK/+Fcsx
itk68AAHZqPvXiAoaUhrrMBxuAkArk5EsAe6AMkH8pIHadCW20LYld3Bd7Sf
LQt4s4veyHDzOqOL1Lm6n1MXQLbc+GVxv62ThJ6pgFGsBpidCFy2+8GQ12CZ
sZyHqaLa7ADppOAjBdw/dA0ESSBMkFBNlR8VSD7OvyZdaPVPzQWsKeGZdBrY
AdmuoMPoPnrAk79oeUZd2tqr5xptTloOyMmu6YsK7+fCWWt4aJOHp4QLlMhy
IUlRJcD6pwcD1ra9Drk0F+zvZLD2S9GMPsIzKu8UDR5u2L++x5nvih8Za+tO
nDJ4cESRgLXAYiuvLDsHvMwpo71Rw1ItfnwV2zQubo/X1qeXxqdZdXn9UJq3
0ZJMm4q11ldfXVP1qxjPQ7g6jssiXSjahCj5VWnd3MX6GHAs0k+QH4b+VmGH
LeXVsycBOhppwk45EFLTgP0pwO1Ed+9mJffPATt44SO4vSqEUcTbpWH9rOwt
Rld5wgkRXdoAwYFNGEEmcksyDG20kfCl9oWFUIUZmPCfhgnm3rzbA1voa4Do
qOlVFE+dWAdiV/bep8bN3Ru8L05CPcXiQdg6x9DL2lhGB9mkSFEvl3JocIB5
IeTkGcm4slqQcGjAb3MtOmctfhVx2mzDmQVuM5JUGggYSjq2e2sIrOjGpFCz
rjhPs310zsHrfTO60aDVwYVczGpQOUzxpONof6APqiUPYUqrQZD8Ty6kosDE
DrXM96wdNMojx5TmoI5+IEAQEJvUrLE42R3p4rjT4uQlVH45j1I3GScVCeOm
cUi1KJUmdPNiAtDWNbXvnVEP8ksjrpj1Txdzd6PSkT5bAvttO7fE9gmM3s/a
BaZ/gGiRS+IyAp1QLWNZspC9VFOaGKmhtr7+OIB1ELzB+GfNy2OVO5BlYBbL
UNo0pJ6ZU0Ln6ELren5B4l9n/yQ2NF++X8DnajEClN5mrHFV9+PIJyr04A1N
zPmzFWthnCbm6rsvtKEdF6ycUmKAEsdkgr1YgbjRToX6qlwTCztliBkbYLI7
8OPegABf5q6ExjO+BSBG9XmMlmRKN8eIMo35A2jPr2utDTeAYkdp/RwYzoBU
vonSxtA7wiDtWFZWQwx7A3JzqEB5NjIu+LGwV8vAZDMhglLwU+VtZR2BMRXJ
5iBIA/w9Y+XSC+kU250PwmfqKLo0pKewhBvCD+tC8vWlONNgeJ/dEmv4xE8q
1Wmfkgpoxeap9XERUl6tKRAEljCiLKJ8NdYCFeW4P4GqDUMYpiyNIuRUIHt9
qLUZ4RErJuhgTXYYcXYZSWeDXYMZASDIBXCJptTeYPabsTsVwWHZjiY9AmMM
l+VVU03AzrObGrlZ1UV3eXeIKKwVDxoksQ4zVmRgvm/8v8/xtyOTSKLUpw9h
oLUlfYeQr2EWCAcsk8GsMrz1t6wNDCAimQ11qQNDVzM07ytBFtYniYp6wbiB
uFxRcWf3sFIeR+3/y2TSebsqkR8qPy3qjvi3had344yE4FEvi0cGg0pylM8u
26VKwDmJhuv2VWw/wLsmqVxvMtrXYOrV+LndSd3LrjPd6gteeCO0YQ8k/VSN
Vz7pC19p+7yeM0vrXtUsbppqwQdDQRKAhICqADvQ+cerqXnU5jw2hgMSIhq3
MBfrf+jwGj5/iMcoUeRXL21IIKtXGXxebFWlxEefZ0amLpC6VZ+vEDHHwd3z
W1TLOZcdK/aFNgTy3peygS+nfc4mqil6L9wZJzIllJw4+WtpPii5hs8kLX19
4YxCrtN1hmrBBa9hMCJNYl/tetBzo3VdXBx4fJYCYN7AIeRIdkTunNaigBS/
WfwjzJT/oR12fbnEtI8XpoXuGwjCZD6s0wHeZqAhKZmzXrKL0I+4OgR97VMa
+D1ylBHvrg/X1V5R/NkJnZtG8BJtHzZtwpryTsR+HSZ7ZgbsETw07ZnI4TkJ
N2oyMSuHT7aiCmtJfjSnpXhxA7vTTrfqFPEYlN9zFgEt93sXn9YAIp/9kKCe
Ut1dhy8XKrcNU5VMUjBoIZWDR/I6POP9o0lt/JQnjuiaPVuTYISaM+uspPUM
xDSQa8VQF0s+7mJ6LtTffE6mhCsxPnz9ol4orxqPUiZxW7b8x9ziK8Uvkj9+
RoimKHlmPUOW/p+0FcrdsVpgurBWQhvh61XxexmmwAvpY/vg8pGv8Ko3NO4q
aLLttYwBDiUyqB13AavqJXAWq2BQEgzdpPT4D3Ybffh25W0ncQckbVvTDqeV
lonC6JT779yqoawr3mexeYulygEDt3WjOrWLFvNmk449z2gBJebQrpo0+uQI
6TkxWre6M+kzISDEV0fyGENnUGIuLUW/K4rJiPfVoDZXe9Ox0cai8PXCWAh2
I3r3EayGpE+sOMxp1gprFLF4gtFfdl7686nUqquAjikLCsOVxltW8HVWBJSH
7iryR07Vkd04mm5Xoz32Lqv0750KZ1J1Wneel9DhOIVJ0QSFB5bfyX7BM4NR
3213Cch/lQ9HObB2I8mBDp+Oauc8AVDkpplTjykHYSv2nNAzaYsmOrHIVtfw
CKgcLrxg+zL0jgUZ5CcreVv3PAUZXedcX0ms0pULD+f9WGVl3Zjo02Q7VaDZ
ecbL9tY3z+EySymUGLyWX7fEsIRKYvlgbBks5fw6YcjsxDYHvJWEb2DnL7Vk
FZGEJQnNoTDCVuGkVvf7xq+XgFtIXB0KYo2z9/g63O/xmKYUtH9tG+ZlCrjR
S4QFrW2GqAVLw05JWltVJIdr5IB7dWI00Th2HnAk69aYjYeB2qGfJhahLEI3
69Kyz81wjHl9F75uNnfoYKfqpbo/WH1FhOXp8sJAJCeWD0jlynGaKc1FoaxL
mIEIiMe29rrNXLdu17KKpJUWbGgaKtJxUYxFHPTi9fyvN7gcKaDwHTirBBmp
ybUFilj6bZgZS7+7PvsXru/drtDNvp/tNOcDewByfa551cex+eoyeiYlFLWS
acEUpH3cAFnmFTkPBSYtob4ev7GF9eLxtSSqRJF+40EepErGUBCrWpLXmyql
Y2hku2DVYHAJ6FI07D5AISpksMZ8MA+B/8X4OPSE/ll8gQNe9MNCnCHbt1b9
mxlUSpSdJA1lTpnxtTehqgc824nDrxQf4erW9E9JxLlnivKomTjqTKJGzfVB
tHt+9GWCu0FAYTdH34+/AxuzI7bdBor+XYgD3H4fnv+2xU2+7gJnFgf9bpof
UB2grY3z1CqMH9MQ6DVtQOoDyU0lfMBZIZeNW7RFaTooTP+2tz2UhUjLms/R
Ao7d4vhsdvz9wWzLg7Xgxz0dMPctSKwpnN3DAbt55SdJz1uNYMdoQiz+OHh2
ma72ncBNDI01BBT1HIKlW28aoi0q2IuC4rhTQyI/VlFqjPFaqbTgr2H9+nOa
yQaf5RY7pWaGPTxpuFYKlMJ2UROqF5aB5VZLQRjxEgyVQqv+ShJr9rb0JbPk
lPMyotKq5BvrH318/mzgtIxEJUjREmO/6uBvEWmNlYpqF6wBJ9GiXRWoYga1
DdZhy3ulovt+yWVwAl6A6g9AgFSMaqI+QkGoeZUvg4w9l0g/HjklBfHq8J84
zefiOt5/S8nQA9+Gw7TBFMH9dTv2fQKtv9NfhPNktkKNNa3HfTY8PRLhef2e
I1uK0ab619OD5T4klyW1DY9zU4agTxttU0vSvRidRE8Zcu8rJpp3YwGqN+dy
M2j1l6Q9rVeMO6/J1dMkz3UVBJZS4a1YW1J0HN0mUrSpISLzqzubEZClWsWC
jcBfdzyyLCEvswCCg4hWTQyXIuCHgHgHk1JYnLPDKexqgyQJtSBY8sWyaKmN
JbDZQnPHEB9ytJGb9cMiINdzuhASaKgbUrNXScSG/bXdOAb4N0v3T4h02qy0
tj40e6BfzX/7+7tXQ2uBnz9vlhRcSgtGmzLBcSQZp2/l23tE/f9/jp4hqtBp
hU1/9KXAW/aRfpe1EPkBKUT3EeUUbUC1aRlAj3S0YTdiUdmkWV8AelNdxRAE
/LVftijcHn2igu3ePXGkUk70bdCAN80X96IrjmE8p/MwZvTUnMB7x1ax83FM
DkRV3k8Qtxh92AJd20siu3BbmzzlF4uNgmfDJq4frT4J3uZFBf2OESW/dASq
GshuQQUKOMU4mQvRbnVGfidTSuMGvJOB8deT9FuLpHl7pDhZ7wRXPZDaL+Uw
fAAmxUOxiwSYDCgO19VEY3n60hALoNGO07k2V0sfxUIj0ILWOcB5ki6+x13O
AxB1EaaHZVqoYWFBsrUGRo93Yqc/4xtQIgcHZ/eaBsUA3yxaFSWND4rSeFzt
B+q3DGF+02MtcLLX7NynRTKz071E0zGtJhpXsCNECX+vW/fRgSHPkGmlZPez
oFmrW/G2xuw48LWFVao9tc7ODe1zEweno3mw7j+TwVtT2XFEDriyXP3c3E/T
4JFt3/E4BMgpBDzMP+iGt0JUZmeQgJ272FSBGsGlHXVCWIiG7BeqVd/6+Egu
eA7VbHmkfn8KqBWI6zbXYs0HIxpSEXOAk3T+6zUntACyYrfd9/ZQtcsVPFHE
iJkuE1US53hHH9EkBufgwUrw+9tLjzH1ahkRE3m9BU2oXDyTtgDlEToow8+X
+ZhuaTxFm5McVBM42B1F1mqM8oDJPZ7dWoizkoRYTzAbE0lsKBD1wJG8D8pb
YBi6skvL9jgogWKXQ3uR6yqRx4cBe2iB8hAOcUF1GPmRxyuRBwJSD4ZhmA1j
gaR7qOcmbbtjaxctHyx7gePDOGEt3eZ/fiJB4gp23jrec36GqKNrz6dlkSA1
6QI4ym2tOGxkQ76401bUTYxwXGSBetCftI0y6l7jzwfyk6pKwMZoJI5JCOhn
lLvSqlhGohlHgXkoc4WdmBg1unmU+KFfIiYgGp06Tlosa3v2s3/fQrcMPJy8
5r+KOLpdGSNxVId6ODQNAwxaEs23QGeoqNCUSaWiFvOlYpQ8vwq9J4T5d114
mg/1Azxg5E6BuaHaEYQErmODwmZF2Pi2/c93Ta2UucLKb7Dh8SOD28G78Qm8
k4AmlhZ+DZNTAlL4L62XcvO7D0ERQf4hnl6E5CYLGPjdH3DiXdh7WXCGko36
gwVrD8NS9WBQPXDQlIQNZoWL6CC5ddPk4WSFfTlVOCNzdBNzscNXT/tfoZYp
fpPPhSO+U6aWvbzxTN4Bd2/XJHdooWXfHmVOSsq3I6mR7KqVsZKoktgcp83n
5CKB1+7JBGXVBthNxrkgxY84qIMqTDYZxcPRlQjaHihNDrS8/a8RD2qcth3R
71PN+XMTJANZYDuzqAwLSKyY2ATghPTq4pdQ5NT/7UvHjGqcag8xkiTcoGn9
6Vlcb5UAXCEvVd0F8ljD1EtKJg9q2NIMABsrvyKThdHwlLU/W5cH9EoXZF2e
OmX2EAkqxpmG2iwhyCBb3IWKSQ8eekRel4SpI11mhomZCCMT/7V8iRIMyC0X
OnH8qQSmlA5SNift51lqD4/g2sFFUHlkZsmDuuwLUTnSXYXJVsfmR3jbcZM7
krxSZPWIWloMIYA8DT+wJYnpQfpwmZx3zym9CNflIWb18KgXk2eMXbp476ZZ
8APDwXLWkiaIBCxea6Za1xMHtRcXrGQP59LtDU+f4L+LQbFjUiHl69PihVZC
HTOsSKpVWEuIwzhSst3D3tfr/5jOUm6lgTMp9sPL2Be1AYQClj4qssvhRm8T
04ObeLh+M+przVh/vnk2UuEjH+ZpG9Ih0grrPDE8Hw4U4BsX5mPnBdMuNn4F
4WL3Z/sa3BS6PyBQIs3ETtwpxFwxeLsDj31sX3M8ntQmXTZiu3aP5A2VDB3Z
98YZLI5L8qG31A9V0PWtYQhFWIDzFK2fSLP2Ubl+r3KksqW2aRsJe2V/N8eA
NYFrIvC/AUnQxJLujl6c6PKJAzSqRgRCr3jHnkAcWq7TkEac74WDxnniPn13
aQyHDORwjdpDur4Fk1tRhOleN/0E1H9Q49NhcmkN0rpfIYA7afuvrYkkie4j
b05zhQQdR51Ley9loJtWqxEfS74FP+ZFHEcJRPZtLBH+COGXCHg1Y+V1gu7b
Fa2jEAUawvcOAheL8/a4YcHphXEsGZvFXWQe7w4uW/uiFQxCTv8ZCqZkspN/
UxSOKimYi91HbPY4jeqNnBbJtNZv6UQTnl9+2JyMenHDUUqAef+p1I4GDeqi
GeZ1KkBdLgIm74SyG9fXnN/4dxFzLl3lw2xwND6yhMKY1CBL6McYBYaKq8id
1vT/US93rWK+nqq8kD8J0PsD9YxVIbDGjQS1uuNZb2Gxl/etlNi4vA0qn/X3
Js2ge1YMHCNYRqDhqRV85SpxnFmpamsbZhAqTfz0jZEjYaNAYcEWVCNHNgt+
DQpNqu0OUlrsCJrzBJQYboKa0ArSg6OFpK1DgD2DvPUvDwR+cWeJsileIXgm
ON08wG8lfszPp+u17OfY0dc9Y1pCaSR2mg0UiYsKUdJNTE5fAV6uD76uGP4N
fg1qPngTFRXnpcTEtQ7LXATcpNfwPRpUy0sxHwGvD/JZDOmXhGFpJmyqzIPt
ctB5WgnTOG3ydASSB1vO2FQPeRZfjuvxLM4XpoN4qRznmUZmfl84z8p3pzbH
U6kkv2sNAbT8R+LOM4e5we4zxfUNJslwUslM/ExD3lEkDn0yRXa4L48ihGxD
fmGEhyRsv7VUR7AtozgNVXtwGwciYm6J4cnsVrVd5NYHEV310I8i7oEsOWb9
RyagHZzncLwDd1MspYyKdYwWrKfMYl4ruOMC1l4QjUA38eSxtPWkxvMqojLu
ZMzz/rCW+WiUMeZRWDyAXF/qGN1kzx0M4+Wo9T5dFNsAGhuBBwWxcCiZq+82
GFgzzvMYhXL9A6drAUS1UVuicqY2HK9iTS2pJWVWOW3Urogt/UjjuveBjKti
5Prj0o9D7pUYw9430pusZr5TR8w5v9DhNbEiwL5c+74DLxkTl0ROMi4coGsB
LEfn9HDPHAlzJ+OU2VAas5JxXpAdreD+UGCMALx7KsGULnWR2Rsr2Lk8J0tX
xh2sURoTApgMsTs9+vjyF5i+fvyTXPL4DN2kq1e5YI1Yokf/fuuZYFESEOYC
dGKLT4bi8nJCs9FI8NFweMabaAQypExUvuah+ThL1MNyYMWmaSEzdSHNqRIv
kJXUia9ZcmzTuuKtGZ0kVSek6nCYvc+zbltuYVF0UOjI0TVR0t/ScV1fPioA
vQ++rPd5Xyyymuvfr0GZkO6WkTkj0qbEV09N/R/ZQZStOkpuNtNgxFhbWi95
amGYpauQcnEBzO/0GC6HJclfqHZUm1WoRfPw0icB++U48CfSuHZEnim81m1L
Ii9Y14keoN0HqZck3Z6vvOiXCbLXaYQENF0xR3P59dqMur5yqOxqaQyagrmP
zbg8x9BkVzD34J5eeymgbRq9gzWWL2oiPV0Ner16FXKZkwdEola9ZSWRucRW
G8dAtYJqutMPiJHtkGQ0iVQZljhoJQ664PkbnW/7REUkCSG+z5g7fObAAtYY
e1+w9qdahtPWhmeaHgnwgBwZg3cOLWlqaEnnb1eppG2BLw5GXmjcQxE/SagN
tfeDznSl7bIW3EATgWdvRwGT1w31+NBnDFWkCk+Bw7QVCZSC0ZkK04R+swuI
kZ+6aln8aQ7zQEMUaPbZ1l37qnRo8MkYZFNeDbmIKpR+THwZ3K0acj1Krfj0
rzml/p05EgXSej+M8LnOCzSVaBh/NsHLbnqR+HogVlfrCCYBPSktAAoRixyJ
nlTB3vuawQnFJctUEzh/WlEpYOSfMVM8RTgCuq75T8bn0DyJJvizw/c2H6ZZ
4AT4IUknkGxc4hQIU2l9Z3UtugngUCXrtgCB0dPfmEYiS338t4mZDeg/p0Xe
fVv0dUIzpLLLmfwoGehirtdATkOYAyqg4evv0IlWRXeqWYopOLrOuiLpq6Ey
YDQJk5sWmwu2S9Iae8vg9vFflk+MP2b0GqPLCxDNE5d8zsLrd2w8rlmPDbEs
+3q9HfmzclbM5zXYB6iuYg7xYh7IsA1vCVn4zj7FMDYg85ubHP4kruFsq9n7
6xGnG51zl4ME42pudiektZDBxzs05BLckH6FzKPjWj07wrebmdy82C2arGyY
6cXhJjVgQLyyrm08o53ZWskx9tiQ8oYthMOMwo9QJJghEQN0H/Fo0ev1szoe
iopXYbVkEZiEsMDSOvyeCXUCh60q08wJDRfA0I/4T94+dppnJzq+4kvN/NcO
+uk0nnn9BKhtbymt93QnFezrjbNRlw8CrjdRk/JLP1ji6tEingbApVkjPl/H
LxgO2aQxP2P1TUyilcSSbbKVVO+jT7I6yBmOW4ub9+HAU1AJYz0Qr1K+wD1r
EAxzQ3FNYf3tfQrZ5CG70hM6F6PV0z8kPril2mEAadQc2NluivaVdLhHFjRT
0AWFozw8hAdt3cX740g1qSiLPU3M/bqoDOF17wF+tB3CWtlhbfuSCYlWuvQm
/V6Ju3aO4XgknhbtrNXRscxapWCMbXEzECgOPR70gubSSajoNp8NRf0Ec7L2
alpk7hqNNyL8bKSvZKI+ulr21hc3fQDrQUMUhvJxSr+y2ZD0a0ETslw8FT4t
jCuDFovbNPSxFDFlLmAggv+zwJj6hfxI82QV6uc/GCFKKqjdNlayxt8HOYn3
qSZuItgYIdtxzZ8kZrZc/yaaXUb40K7j6x/Wa5X10RUn4Pdru2+39hII5HqA
F3kx+Z4Xo9txZfUVXCoiz0aYuUxmOlUPoXen7mhzoosYvzy/8W5bC+Tm3Yxn
Ja8IWdKOiBbYe9ZzPTjyd5FSTCQvewklHA6iJQdh9+AwuyGxTulfI6qx3XBx
CD+L1BGFBFdvruRZjwigk6R4kyGTPHbCmQ3Q9dPTzhabSEJpr0cvUXxNMrha
rtKce4chIq9WzXUvMDRKjLhJPL6mGw0H9mvFJZjGjl5CC0Gb8ldoxC4WNS5b
ZY5V0e17JQtk3PtziX+E0oSeQDBb9yIwr51IGZnh9wWhxyr3HvQfvNiDIlUr
+B6sFGfJjqMn4IypydIi/6UXVh6LDsQhFl4twnnMuw1PW7RqZJJXfCsqe542
eG71Zc6+MdHqkD9zVPL7RL4+2ZGFvqrO7Ma25irw/vgha1ZzZyn4Vu0TvP//
/OEz7xU+9r9ip4VlFQ8r4iAbl8Xxn6xIpZqvswNRI4SrxA8Q/6kATLWwCgq3
PhwesnyanPvtkVbq0Nd2mwsR5nHz87gKoLXngw0wdxmU9oj/HL7ST46Cwm0g
dbMHmzZaKjOriQ7vGg1B91K9UPyfrpXE9Fj3YbqbblZxzC/wTEu6Nxj0yDf8
wuaPganMzM3DdG/pI6azI0iF98GN2vnU8nMXfOjhVeMPNhE/Vte/pCHe3hxD
MgSw5ChYm3mdR1fARrNMfnkLcV7ZVi1u5tDr4M87kTDp3PXNAsXTmfb3mzA8
MRezY6xvTxCa6Bt9keVdbzeB9s9fl94/iNPaB1Uljv96NZQeQiRE6MG16tMq
PuBGznYwHJy2p3+SWcBgVy+qqnzJzzm5A8ixQszZjm1JV+Qx0DVPt+kJGLSL
i2tyX4ju+YPB9Sif7iNbp8AefJQ/Iut4E3AQPQgX7WFzYVs8SLc3wZAnNlIP
zGNbUaT1YKewX4sapz5LsCYmWfJEa1/gpl2C1FzrXxAi3DxNla3RYa0BtB7n
aubjcMUHQX1g8WdeJNCJHOIJ+RzDm7b45Q3wI/u7XBiOQL8Oehoaf6zceDkx
ZGC33vd5uXrOfJdYd85f53VtLNFzY9RjbcbaG2O2LVFLdvHFAdS6aFWolmex
7Sgl6QgiXgcj+62tjNJNZQXBA+6e7zAMOfvMqw+i191csOfpRiKHJ5Bk3gKq
V+9Rw1HashW9meXzFHC22dTiYevBIDm4c2p3gnC3xRMIEsRQjfYybgRfFrL9
bIPlQ7zscVahDdgqtlSgNDwIycf1cT32rwXd7VvhkeqTW2jJqiL9I7nKlmFN
smwsREShRTokqswgXXwrlrC396QkWl3YhqhToSpYkg5K2bmjEhuCpsMtvCdS
WuEurzqCS7TkOdkQ4JymzIj+ZlGuQz59a52pO/YvOBdfZ2qpB25nLNH64z9B
G0E9ArxRFbDaTrQ0rjdG+gXx7XZZvy96v41fNM1AMbVlDyd/vjQX1zo6yDNs
vW8tPVibBXC9fP2L2APwbyl5T/5ZOIx8s39GFHUCg4EWFE9Tc1StJRs9VZYq
F8fkkyj3KOFmqqSivre6WPO5Vq39Pewa8EooIuKVCXmJVoxJN/kCu3AErz7i
a6c/qpqlJTsQ9OHLI4DvmtQF8umO7Glvv2xU0WhTSFgSo2/G1iDzzWxOuoPi
Ac8V8E7GCauP7xwMdxycI7GB9DIeanTcJrVP+Az7dj0tqjUxEdCSjF/xWSUn
P2mFDK9bsEw4AX4AjpDR53v1NMc29oQVLSyZMaqGSn7Ci9SZzqSbXE9+ZR5z
feO1KSJbsgpp8PpvCM+PimYsHDgIFIuAbW0AdZWfB9qDkQbv+NJ1FkMnD2jG
qESXgpL5FHGH0pt9ObFeVN91jUP0ORgVmJxIWQW17BiuDhB/3jurzGVQ9Pjc
OYoqe8bcRTQPRsfSQ+Y+4qmfuBEbRDGOqZaRtuiuaLjZVmAz97JolNMuBMyy
roV6BpNxwRli1JMsahjEFK+EiD1YQnZ64e6jGXZK1noj+PP2bUkISTxy//L+
JSO2VlNu4Gjkl1wqZx8k9eikLRAuBTKQ91LlKiY4iZK23Oza8iRFxvPb5K7w
CHuR+u5djVLsxrhah5zSOr7fIskcGnv2IwfIVYzZ9D+ib+MsBLy6wRG5lsJH
rj5+0gH6TncrvFtibV3Sccq0rImtgiyq6UYE88OJcVQRhS3wzE38wzFGGZCC
AvORVTpTpPAoDeN0PsJz50Rw5o1B5t9YAJpQK4U0EtnzH9hj3IlAM3mWsakW
2oX8PGPSjh3QmE4CMizChI2p6wXw6exe1dyUHCynIljQuS3qs1UAzSPqHY+b
QwbPfrvj8NmrECg0PEaNW/0I4p8RPF/2QuqFMv+n08jpgXvJ3WBhhdVjC3Px
K1qDacCy6zT4wFwMi80DKfFSPVjxqB6HxKPeX+AP5/lDgLgBk8O2Yx0QvPbU
by5RfAuHKttnj+/EGNbrJPTNidArhGvWgDDJ4DrSdBc5fjt4HChho/kkzkUi
jpsRoeYAUZ3QyXm5zOQc5tmWsHA71UVy1G1ytDMcFlOY+o9tQ0mKmA3A0UJS
h+CwRWsT6mqWYACLTH2uSHsxljBRliXIIc2zmpyON9M8teyXD+Ypc+xb1suF
wvdNpmKeuukAamtSh4m2XQzw2+WT0xoRthKi/keUdv1k6wuQd8oc1q3cZqp5
EU7YwcmRgApiXpN0cdTftp4N5JchIXL5PkjVSj/fzTgD1I5e2F3euAk+UN4y
jf6do+6VawCy/cUP/z2FKRs3ECUMvTvztpvORH3Xo+5y350Ff/n0jp/qaFlF
RxWyCN4Ncgn0/PheJGwsMXhZAluJFRBTO2x4bThFSSdSsoh1kEh4yPuKX3zw
ncUwcidAOtOsOlA2XIaSB3lXjIuradNoTZsXiPZB+Bu82bAdaY4pEDhwh/fN
LsjxnPHaY5iljvtY6sa3lA/zZqCCYDG2DB9l4DaThvgplayF+USwYEnV4A59
uA6c1ODvAwHLb+LmdBpbadGtxAccLmR1JIbf7epIwbpDg2Ul4KKct93GI8MR
2Kte/ZnOweb2Vs/okftNLtSAfU9FnLSQJp3m7bwqKheuzuk8lAK1sA1R382G
fLsKduvts5NpnI4tPhosIVwqrYVDlJStlyqFBc/XwrdwCesUWprWYnYPQMM/
xgNmt48MNur5cxEEyaFBHeYGXn3NXkhY2NiAARtyF9HzhWJ32A9v3Por8sJv
PjjiylWgT7E4ur48Gf9gpKhAQHQxgxmEFmPNABnT18t0zES4yBz6mimp0wAJ
qI0ytpPuNewUF+a0kMCR36Rtfu/9fRuFuxpBRFwO6ya1D3jQPrTOLUq9FjCf
r+RNkwm8Fu3F5F1zDO19zpxDNlzTnXFoS6qugBu7trOQfTmSqzm/ZrcqQlNN
Y0/PW4caSLKA07NqUjNHD0esngXRL+m05M38B4U4DEpwsp0DRbhOb+qfjqSc
ik53banczg3St5x5chXUgFe++RBj3xQ5nyPDPYS7YuymtPLJ/5WUkejYruAD
UUecrWVTyDAmehW7NvEe3ZEMUosb3jEjG4JiYJjTIgGg43nUUDJ5C6c1mB+i
gsxKan+RBr3JVkELylTCMDCBo5fVouCHGEfeKsxlikVT4NPsHSm41Uzt7Ibz
HH6BY3Fck9WvJfF+1Fi5LQD4eb7g+z/xlU471yKmOQIAetj5qJY39c8NN5dX
Sz7qnhZUiJ015GbnVVu5KmjtWbeAQ7lJ7wR8IvMhodVlv+To5Xm+zh6IWpv7
EszVXKI6PdnnVh+1ksdqMI7lpGcMlZJ+4SQNVScX8aoHtDEfEp6MKsArj7kM
D8udn4ia4arnKrvUvfEvYCMzzGwzkxed2CC6sYQ5WypHdZOn0NsbdE+dL937
JoWvZZXfd0JlrYhwGpvgQM+4J1NBifjEV9yHWdRcctE3qXdGA1XZDDLOJRHz
+hc7vIMShH1Huy1TwgyvKpdeNoES+g3c4PfhFYTBDraoKHN6CoBqcmnrBf0u
o+Lvt6y7SCjQtUjequEIhRfBuPJhW68Lw1o262p0uiBiuPdFfSndho9c6lu3
e+LPNSbkAcc6u665U5UT/0jV0y+b9r6SKrYWIfs4XWUgNf6nU5t81w8bhqqz
cxDrAWv6d3n1ebVaWh/Ogd6Ar3HMqSNHWWQ5IvNraSP3+MGVovLjHF2PyKJN
EgGdIL33GC+8RY83rLz2mjCL9gIn9eX/3L5adDFSc9y0A/JWaoMbWTjMQl7E
aeV/H6OE3YI2IxYLeb8ORhPKJ1oiyKc49pw2V15SjicIeTn/5dYtyXkJlOc/
cUgXWNR+MrtBP0H6Q/U1eD4L45OEFgLkUD8KNx/s/1H5Wn2223ip/9UwVGuN
N6wlK05a61xvrLcj7jmWQwYJt+bivUSlEo/fYIWu4Q1QybzkAloHWSH0Z2NE
kv8YjjXdbnNjCkOiQh6Qo+uU0XVa80TMnFPmc7S9B90fXg14gzO1HGisNbsp
fYx0IdpefVn2i77vqjZRc0s8eYi19E28YFWLi9aVxazRaJK0B7UxCVQG4ztv
HKwu7KHEq38CY12N5pca/t4rsQCn6QYsvoGYqwSWb6a3PlxQRfRGGza+kBET
sWxlRuStGxDdsDhn+oXE6dwsAJZD+CyFNWho84tdLj2CiwcNnGi0uuvpLyfp
ND5gQkXzCg3W3aK6bz0zBOjRkahBswOplQ4U6rzcNAOaoOVCa04tBKzKfnVl
xvM3a4lQj0ef+eeDBgzPl/YqQjMeX0NVDFfmKkmqjjUf68hJM04Rd+whClu/
y8BSU+mOEH+Ag9z5SRikFOveH8Pmi9ZMuuyG4r/T/JolSQvRCWdsyiq8YxjY
/LvZGsuusTD3djzVo10s5ldh1aCSViW+HMz2xhz1Lim4fkMqHEDCZyPXY2hE
mjE5jzLrE6H71KJoPSsVcpApCSFRlFCsP/kKdik+xTd9LtXsihVe3pSsAO+L
Rwbjw2Vxx4wuvWPnue5a4mXiW1k4B7CfeTbmCPMLXBEDvPekHL3FCnVEM63B
MDFnWdXShGNO/wPuX6VrswBffERsneuQ30cdu1+88N6DftHl4kKmpbZNimsL
3uBlaSBlTwmf5WjoTHwBI4KJUMx+1jS05OKWlymHclh35Rx0vPM5UqkO7wGa
+TBYTdlFyu2KxqIaXIi1Bju7mZ95lkU8gZewfy6UhCAjiOM/FdNchGu+uwW0
wP9SG2BqMgE4gj/aGddQEEb/yUuS1roW3KpgnrQ4mQRQrKVHnFws1+rgYBtx
ZoyUpRg76Ne9BIb0/EIAHhlfp8kI/cWHYuKmoGKblu60xvtf/vzCcBZ/uqF+
AuG/OSV4y6mLkMhZ4wsKv4OShrJNHBrtyF3MK3GaXxLwhzYqzIiVJgWcCOP5
HgtOgSVSfepsY/fchC+TzXtm7R5vOv8Lpuh/1gZUC6BnnV5kZih60SvYDD4a
fS0XEkAmWGUm6VHO/WrtJlHkVdxDbgwfh3amfoFkAmjokZWVK0sfDPee1rfz
IdAZDIDfu94KgQ9ZgspB3pZR38WmsB5RDipXWqzT4rkYx8huCVUHBikiSkEx
Yf32LZ4Xro+CbiAStumBssjn50ucQoCUY6BlM04vtRCHkKA4Xh0UXjzmCDVw
dn7okbNyEDyXQt1leQ+I/yOlvh1hgAZhlgyIOo+UiWX/Rz0307CddxnaAiZS
OI2eoGNOajrfIAkT7Up3a+bBdowxwffUBIRT27zEICuyuRdSUb/vFnj2Dfn2
Ssmop6cl5RHR7naFeRNi4XY6Cwre6aqwLyVNVFHZ90kp96IsZFVhJeZ9aDpu
4sZzGTRdsxboRfKj/I+Jt15fsH7r67+WybThuE/Rm4NB+hbrnnw9fMGKwCs9
I7HiO9tEG9P60QnNTiX/N7qOImLB8k5mTGTmi6RnB4ex7ZRMsSOLtC2737UP
/qbwTjnQL9Y9DxsaqdM2ZfZlYxVHzI6wj5r/BKJaSm1ELL/PGS0etYu8M7D/
K7vhPOG1xG+ezWStSRBzhGbUZQJwN4qHLWujpHV0lthUP7DCajr5yi6xaY0C
Evxuqlyz32k2XmCW5VEJ3eE9YXVPzSOczSWYXeOWANFOTovSJ6jwNmbuSZRc
l6Vw5QMPrP2X5ej6V2it8tUZ6BLTPGbBIyuiOWeFOZ5YBWDD2yGpPubmswpD
E1vAfl4au0x7MhmZLHeAqp1CMuOYsBfJTq12cN89qZ0kqe6tEukuGzUz4ui+
+4UaR1KOc4kjHub9SKP2sU65Jep09Kn6EPCpEvcsHqGbLP8DQQpnRVt6g/tl
gP2CFdXi3NV247nq6Ygx8CIMA4JMcM5YWOOtw3fmYFDLxEK+g2VWx5KcnxiJ
O4Fv+gI9vI90jywoHHwfJ3ImqB2rr+kjtpO5YpB9mi8ES0kOA+AnlQWqhpY+
VX15WVBDp8G3EOQZpxA0habXlUA/FM1VKQAy4+wQUcVkHfu/bsuOuXdS7Ntf
aGR2hG04vLEycPaDujlFCQ5oGmSpx8dAANp3ZeV6ez4SNLRuh4B+mgzse2hy
sfKV8XzDfT5H8WMgeWlQonnmk3Jw27nVE11Mh29UzIbX8O3sWui1cX98ypE7
6SpQpLJ670EBclOhiDo3kP3Z4cQYXjm6qvE4m+lYhBt0827I4VOCrQ4ru262
jUGWZrm/qbxUFBSlfPi1WobxIVSovDijECMInuKlsVhe/GjSNHAFnOClTqY5
EB9KxoeXfZHY1H7TSbaoSTOAvT/MuGt5RmTlcyVSvHH75KjPm/NAJKQqf7T8
PpzwfXs+ZWqGZT0wNBmXRKOiLynBxjINsohZPinCmb+aFlKIJjiyM5IyBdzy
XV+qifYfW1sUPYDIvOba4kH1STw+fGc4RqoXL9mi3T+lpYe3izpRBVILp76Q
7V9VcVmwylMIwpRuNViqGrAZvdXpMBVHPMbeRWOZnS/G3wf5mv20NG1mQPP2
Nam02bJ5W3rT8fTUYyOy/NZRfxZvUGCuAyTVmspFiNgfR38tjAsHc7xVJCtS
CC1xbxiUXs5aIpxrf5o6WHVSKF7PbWfUk8ltnFxEtpxUo1KC/Vmkf5XL2xnk
wN9qCoR4385JPUZdK/O9cA7+IqqO8PJCzcbR730NONIUB1f+TyMR5PG/D7gn
RyTPsgTCMjdXzWKWKpMBId1lhVdkeYqDMb/LEWpBsTZcaShM9T444suqB1Fi
FIpg+sTT2bRvVmr0/9WQaY2utaxAOUUocnigi8A2q9nEQK0CEJM4q3w5d7Ey
+s34/GZOkDaH1iYJ0tBizVwe9AfAbrU0SsZx7ta8c7VjK3LMCtMCu/174OXO
oEubDJ/xf5/7sElqmsaa3gO/UJn2fKsr9soHtmO9iH8P6Qei05W8LlVb/3NX
crYExvb8img+XegwhMvqzfxSVYglPlb5E/pOZlYs9Y4xV6W8WFeGTSqjVSjV
o3uNczlr/tofUZrrbT4ej3yEKoNmWhqVzBxNFpVG2yi/w6Ap/xS3tTl9f2N3
Rpnc4MNlsAIdpPkI1kzWy3hrC400XTmLKM6BPPJrdThproA0Upg8THioCgAU
p7ockGK8t6X3tGIH1GDgDPei2/RTcla6K2siHYxZGMbw+KF/rPMrgGcvZlnS
Ovb7/DrzJU1TfGgraXeigbsVzYEK7FsG0xEmXqXlHfrnBUo5dbHQq4hGdyjL
Qk0lI8DU9XRK3YzsP3H9zaYQSRQfEnkv2Ohxul8TuIN+IbmcHxqb7h7hux3D
rtb6KMGjv2L7xpO+n0YNz2DY4jw1CrrKt5gQ3ED8bdqGDB3ACEfAkuNpLSu3
JBXXqWL9sD8i8OPl9ssa0ylvrFjicpREFqNnlsselvB8cRJUnkHmunWVr1jy
re5A5EEyUY2SPY1ln5Q5Ca7ivGq7u/o8BDEO+bkYGqSdKys4z4M8eygn8/+G
58vQaBd+U+pCfiT5QlpxrWoUmlTf+gSQS08FHHidLSMDjC+2mckGWnRcZMaP
Iiyjld9oBc6od4sJN2JpmwM1vXGUogOXus2gQJL1caWCY8pqpmIBZHlEkOXt
BVn8SJw8lQNa5bL6srsJnJ4fa3NUmUm2IEcSjQIY/sKaaDy91dk3lZXEKRjT
303cHLLmyUMLR4mfV4BivJziWbxEm5PG7HuL2I4orQcnj2mWgVa+9nfeE1nn
Yh5iiMLV3cuHqkgZFe9ROAfyQvdBE+aZ8VM6iRmEw8LtbMGOk1ykroG+EoDg
u5lGvlMGf2Tm9oD6XCS3d5fcITXOpCWYO6S6P0nYIhLxCg7ZSOp8gVdSqcLy
PiB6VRDZ7y2P/NG+TDP356NkUgMjCrQ76Ua4gitFoHAMJcbFnLCrw8IYNg1c
VWUrNpQn3uPNSmTbuSqtnuTfApYgNjJAslFJIXaMlQv8HfvpD3VTgxBApTns
Ng6HL0OeeihBHJXUDwG1m4uXpky6s+O0gGY0f83KilLNziTxVxwBGkNM8+0r
2otKlQKivLImsfZFiaReeBxqz0QeDlgpi8g3ePR+nCGpTD2+AH6/AlOqLysL
J1uWI5zMMbCPCdowH+dtu7U/Tn/oxrM+erAHIa2uy1C4f3Aqr1dLC1JWF+gH
uD0cXM/3ZXWESooyRfGZTKQOq3kuUua1s6fJvQdBWd8ktBulSpX6WRYmyZLH
UY23MyQtNf6DgUvsROBmWzNflDr7fy/Bd45Qo84N+H1GqDc60SkyAClJx5Ml
XhR+YMu2Q2B4rRO5yLWxEaLpMG4FpCcJdhhD7VBL2iMjbVrhB6pAIWtdj2Kz
nKL0KcW0Bx8ExqLbzOVXxiq6vmHxiGDpOl6qXirsyyicZ8A6r5hih+VfIw2P
U8uEDeExyqzcpHOz16RwIsjrXOd9gwCX6CxEO3vrb+h4QopdFuqYVDD+N2/K
9jvTncpiph3haTSYCOEgFRVAuE9iHdbeFODMcTufDxf0q6wuSpVKEWrzGbOV
8AaD8+gExvqqjx7UFoIxSu1idyhWdURZjqfVgUzCmOrh1284lZmI7zYvS1IH
4oja256dTGgGbkkGLBbXEKFdh/WeJ45+4oq4F/72ev4CYF5LOGab8BMPAq2w
nkTGhwqXqxHw6ZuVQA3epFmT1QOZ2DoLcXskQqep+uebdzu6MXbFKF3nhXas
Ebu2VRs184B95IGi9tk3aoCDfRZzQNupP3Go6SWxZaZztD1BfGzOuRzywkt0
nAiycA/9/UF+5h5XwOXWXWyTbSpejdju5xOe0bH8MAupv5wBNLEkNiNNin19
hrzzqvoXl8Y+eAhougIZW/2riDdmS7TfRhUiX/8Ogv+OcYTCXC5hz3+ylJxi
4IkJwUHZ3FQut7SgzLkw7Q6Bw6iCdYzPTAHHRIDLhWepJvJNO5BOJn86u3GH
/E9wS8xdymArvqUANULPDB4BtNltb8A/ROqqNO/JnGG7nx7r+m2CBKJjJlxR
XrFPB8x5qyPikmce3hsEhsrWzDsvbNj1henmTIQv0bXkt1kVwRwIw3j76zUM
0gMuPtS31L8IU7J7WpRXkgd2OxMRcApj3TSICxnd1dVFqmi776qXn537KMSX
vOU1ijuQwZsMtkzj4YwNtLgzZ6v6CiZMZNH7JEwwbVH0uasNEYnSZByYSRmi
tq7JnFo6S+kNJ16XGj0r/19icQ11ZeXAiOH997uG/vIqUSEySQlpl6h3Kcm3
K4xaUmhqQYzLSVrykuR8gHu7NvwWLrp9dhcgs6cgaBXGF5SSV2SVGQqOw/jZ
sOKtWMiCWF0ixOqadhQm7OEejF2CWNxU6acCVSsTvjJzTTXv3xbUrg5s6dhZ
yDw70S4sL69TXuZ7OSHD1YL6CCFmonfv55o0w5iUaKRZGtluKE2dmfJy7IFi
D916lABRn0j1W9/MPoumxiLBRyHjVa8hWKU8tQYeDmTVE3dVkXP6+ZOXYx7f
HA5nzLj1TuvLnV7voIF8syR+0Z7Ea1wLgyZr+Uodl91YahiM04VYS1nQuQa+
+MwqTJborHR6OTYsUZCgiemUxE+7S1st9S6pZHm70+UvMecYLz/T3fsgRRLO
ZCVHS7JY9OtxYIJwx4vnE/mXteOLWCZylzA7Rico7UozlbmRKRimUBETSMgZ
FN8JtR0ub2Cbm77jf1xLgKGypEo1TbPbDjj7VL86NnMJqVNlMkvYeeLpplD4
N2fSYP7SAQAM+B8EsIFQBuMnj+414T7MAtgUp0uniMPTQSb+8MWFgARUS3fV
+OQq3GsndcKwI9iwSfPPbwRGx97rAvsiI+XISyiSpmtx1uUtqh5Panxgsz/r
fVAXgD7jV9M3xC0K6dARx/xyY9fDUB7l9nM41JNibgaVMY0oYjpbpT5rvMgJ
tkb+xqq4HGVOOOdMcuPVLcRa3O2lt73U2T9K5ybJ1eFPay9HEpkVliMSUcDH
h0Cnkq9HlJGhtUpQ/ZusFAH9NaZ18NrNrqZqL4Eehr8bQihJAVAG3DRzi3Aa
KAsFXXJXzB+vnb5cjGvzdLWFnt1S5rj7I86bHbf+2Jtc3rWMTM7FfExDMTrV
lnxMZjXJNP3zkarN7HINZ497qPrZy00b32svi88BF/0TEvUcVmLwjF9EtgYE
GKtv9fkGwdPs82aBc6x1O+UveaHZexx8LRasEE0ENO6WDh/odZVsVrT6viCO
byBTFzlXkFE8KAdOFR0sGL/9DMvUiYIHHxOMFiFYTpPPetvY/FsEo659mYcm
ThFQXRkefl9DHOYgATpWa80FQhk3eLiCl9a6I++YNPNR5Zm6fl5MACJwtzYU
IaKRrjOyigiRj6nREP0o4YHEFGSdS/EgAlUwIy6iSQ2dRMLG+FLUXCgew633
lBCeKzIoyOFDGV+7A5OG+2A/q0mCLSrZeRkKURM+ylwxxR1dd4612L1rKO1g
7uM0m5jV531G9G8QN8/6zsAzZHox1S+MtcL/md5dnDftgD+8JMVQTCH+S0/6
7+jmnOcud8WlBIozprzwG8kvrh3GuxUlV+fBF6hG+yIeOKtX4qlggqeZif24
IUf4zQYOANcU+MBFdqcS9FhSn+quW+29jsu8rm8fLVTEMZEB1ZNw8wf038D8
mi8W/X06AVf52v6p7OzKTE+LxRTR2h5AnRVC8x/sktkbZyDwDIGUyyJER0Z5
l7Y0z/JaqTG97EnyzQYdUlJgVMnQWLK0l90dFl1GaUaRHIFYYU7mVdWXnY+v
Yj+sZ65+H63BBEcVqTzSAjVgyHSAjOre77TUHfFnK+/N1M5DVolu8PH/vWKf
MQXzNz8SN9BEoHH8JM2l8o0amqJFUKDrwBQwNpWLeDsrSN4n5E6bdW6XWlvj
G1elCQtWzzkv5Fj707bmi7t8blTwv9MonSVddNDXMSgDHtWT+OIeE9vVoQZo
rYTwyICAwzcXJIdfSd+8ZZTJpCsXHZsXRYeUnDBbVkIa/VrYftnkuZKHiCnS
xLoiNVBINzp4dAN9JB/jPt3WKYoelOBDe8qTZ0E2QguABv0O5lLw9wNs4IPG
NdVgKlCS0LQQadYUXf1ZB4OTfvJnfO+438kKeMNZJIrrgehpYI433Xa0Ymhx
T7lAp1ErSJrM+2eQUcg/ang5zVcDPKvFiw4hWrZa7kHxVoWhu6rEoy3Cys4x
iI58d3WpRZyESl7aC8sd55hhsg4suKYws7R/MqloPiIhbgja8YxBAWJY15BG
S3++KaqzFgs4uYCprq4XK1SUyMDyA9OqP4nmX0BX1sgtCEOZ+X+hTmuDWrzm
fnYbVdQusyr93pqGFVcJOxS2W4nl7IknklXNb3STwcS4SP+aMW5BHK6K02Jw
rWcbJ2oImyPkSK3LxNou86/mQG7pxZI+E7GqxKO72qa4ScVqMFmDH5hcTIRs
XSFT02iNagTlu6HXWmCJoPXJ1zUZKzCwlxFkmHB01q6ecNzXrEEN9u9H99vy
FPfp80Kq3WMf4ycHVTYRvRTXDuhllwWTl4NVr4JCZF0aBCtkpNQlJgkeMrrf
1lGsOmVfdzhBh8wmTzhEiaBPGu3c/IiUXrEQUCQA9SguZghe3Mh6TUbDB9F4
0mSEV9jhItOr2qcuS/knmnpclfKTEBKhx5Hq1ltwiMCw9UeOpJ2pjyWO5ZO8
XqE7TsyH0vp2nTNJv/+YgLMJrB0vwycn2g9FI8bH9Prta8b03FZ5iBuQAleo
SqqbVB3ZZcWd3M/yYdAvVtH427NbEnj6rt4QxP3PMWd7uN35IbGuMdJkn8Iu
ifvJa96tAaiLd77EkE+huUK7xjafX4CVRifNVr838MMmvIB/0UTu9SZ0OiKE
TZaosM4H2R0IeFbAfVbxpaB6GUh1zX1iQHMaX1/9fHF7xbeLDB7SqEJ/X/hR
U55/cu0GZMQ6aBLdgKrtUwURE9MPfVcxpdasxccmDiFTBPr3JlEQ5vazXtOS
JELxxzA8zktA/MFO77M6Hcc5i5J/cCRSde65wLxc3xLJ+D9F/iDgyOX/xJvy
v4HL9v2l5OV2DsUET2WWc6d7tEQFYG+bEFIEEpHIyxLwq1nbc/utIikuTamh
Mj3G3ikO2nuVHTjhXKBg+z5cBWtmW4l7qZMPVBIW1M9nLyCx+nxShGk8CkqL
PGiEiTeCbdAQZ5VXYg7WN156Lq+LcELTtpc12M5GyHsweB0SsSObxRC5Q2Rm
3wRSG1n3mennWsnqQSUtLeoEoSK2dFfow9T0dLpVgfjHpwCdh51BccZKb6sq
td2vhFrQFEHIbB1mrzxtEOYRv+HqFdo5dksq9spZo96hk7UCD48N8K5CObMK
/xmp+Hp+HU5GSUDonx3b1xQIpvQ76LUnDdmxiJ/X0HlZF7pCQUOfpkakYP7s
46d9mE83iGoS7l77gccZaH1zMrXzGRZQO+tMVn2Qzv7DN+OYkUEFJ5su6lSV
ufbpmt0y6X1kj4NeSmYcUW2faG3ttymJMJ/EJjzlR5hvk92NxuWlYZXOUbC1
4oOkzQjQ1+POZxs0p2EL2APQM1VnK/c2dBp6MRvIIHVhHWwyKJQaQZp6axng
CwA3hE6ZCIU4vzfVIYed/s7o+wTJGn9wl6MQ1MjJj6knSK846ZU2U/kJUmUI
qQGRqoTsHAtUB6+rGyHCtTgL4pScVuPHEbSKefe9P2WoExAwSmGmA5BCLxh2
3yyYlixHzD1VfgUPzFvWMvq7zGEc4T78HSVLCu4/M1nWzttTEMAgHRiT/AA9
mt1xkdmCJFvSZ94aZMiS/ccqAVdFqfSe07pF5imAOwL3zMA03Oc9x8BQUYhe
Mo8L0fd3QgkyIGvpi8GM9LJG13dkEhqk8I76S5M8uYgZQTHwTD3T53sz/Grz
dX4doStsm1SDWgiBXWdCP1xXukJHZZ3K6JDTguppgwJ8AMdegXHFY5cVurKH
p2HQdOxeTM6FEDXGn4VbS/I8hBFh7O4YBi8Y7kxIBbPkInUjl9TUYSzN9INu
LDfmma6x68PHeyfOISnAkEdr4X63IXkSYY8zlsmyAqCU8zB2tqVUixiYFFWv
/AQWZ1lqpOkoApx2X2jsCzxaVRDLC4u/8LyMWOXmWQ4L59NPbd7MJnXytH5O
S8wDdZX11wTzshtt5E7U8TNi0euYh2QEEN3wTZDNh9RH1SWvBacJMwsQLvdL
Y8jYrOdegrH97G6rRpurKFltwfcVFrWnr4uGGkQxNLq4l6AV+SGM6Stxe2sx
FXMhOJXl0QcXGescE1F0jpecpYtb/MjNhwCAXjKX3C4Mt6sfXd5y8RIJK9NR
hATIc20ZJlaD7LXr9kEyAZdaJNCUcpsMGqlh67vFy6H/eDhdLVaNE37w2OFS
dEifOuG10aejq1sYBLFvmXBJ2CHv3mKj8CTDbfd4DUIlCbQLxRuAUWRK5Fp8
Q4+GudHkZUvSKJpzZ3gFB8Zt69P50nS8uRJJNeKUBm42OOSc2G5whCIiTX+A
F7XJwjcXl4X9BMLbHqstpZC4Z3DUyPrSu+eFev0eOUm2wYD9RBWoFiXS9elq
nfwCeLWZTEDkfCKtoLcjkxd2qrzPTxISOhf5p3OOmyv1gRI41bCQvBlxJ9i2
TB4dgmI6/ShBD7trEtvCW8GpfaIcvn09tKE7Cj6yJrd/AsNWana8NkV5TJCn
h+zNXiaW0K3gzfjlaR0PUkJromvB9NuTv8YVkYN/uRjq6eCwvbvEToum4QC7
WSuj6zq9E6+KZEm/TauXuYiWSU8rwmR4cCNKoKFSsmfnriD0ff7Hz9N003RH
951SUB19ShbFQKvkX6WZl9OmMKdHg8FOqZVH4qVNwqnbxJ4q4WEa79K1U+F9
bDgd2CMIxENReWlYyWB5Lg/anL7Ypff+5egvFiK32uNgufbREVsiISoemO6+
tw4gklbHE8YOJH6N8vvwYhnofPuuGeUQnLk5TWO+UbmoSwMq/jQLSR+8PVM1
O/LcraLxGPPgAVaSJKeglxYlTS28AMd/JF1oWN5IvyAZLuJvv0d4IAWCc04J
4phZurlPuOAMrvvbP49GycWGqRXemubKNQWFsb5I5DGTpSW1rb1whVKUEr5j
tjmd1LfWMB+vothz2uFaYNNn4x1xMIg4HpgdY0WfC+kpFJpEzJbDAR4FPGYh
YsoKYhmKhY+NcGTJtTYqzcC28sR1icSb7iqW4W2BCWmHlibhlS5lWG7J5se5
yOI28t34W/+YpsDEf2aDk66+NEar3buK1TnLMQlsg8ZkCB+NUU4pUpEA7JjY
xJL1xdLSwyBtY3PuBGlGknbswrDE4gLSSJDusJIXXGVIy93UDHaVRPMMV7BV
ZS0rGm0tUq02dqbFJHBtMcoKJhAHt1QZnn9M9rd4ibVNUx3vkec5zkrpo9lo
joA8Ynb0SXrKmWe8CCKFKRFYL0YAnbNAe/l9QwOtgsgtVUvYIWr5F+p7LA3G
L0A5curkFMU13Bc0aCnKaUYzUW+MtE9gAB7MNz6keW/M56/0tlB7ZzIbb635
UdUq8/N019Q0p5gr0It2FxxgQ6Jai2kU87982v5FjIU1qC3/cFyjVUDpPp8C
ZCHN8BzvqRnrDHnY6MDDfDHoQWAerHZpTWn0EkR6M1BJe0ZUGfZFnhzAh2Z0
Ngpf54YmN/utjPnIdaoHCemiO9aFAG4LiHZ7tyeOSd2uFhC6ivo1VsIIFfdK
lmmmKUymrZ1OyCqE3kMwHawuc5IEd+il7A6PGPt+kTPiYOUqYJGL61Dd6Bog
bLojZWp8q4Qo1ZGxlAHk0DoU7Ofk/m8eftOU2c02By+Vzy/2OTVoYoxnDeHW
Z8UAbsP3SiJNuuLdzKGdJtcszMpUGfUwEn52GLkt08QghVHn3yQ6EL/aPZkD
whUwajm+hE6GWopXhljMf+ZiQeKMVmDskD1K6IZNdXA9VKZ3Nl6OSfR/3nGU
e+06fFJwffMMPMSx8ZEgD37v9gJicqK3YuXKjuP/dnfwqDhfFAB7wsIAhXFm
VdFoGuZSmXItoK06vANY4KwTTHSacuMpMlNRZq5QxxkrAjziDFi1o0jhtnz2
t0MfVBQiOx6O2V8Fz6XI8eIdFlJpObj5R9iaMoXCmYTuTzTADwFuRiEQhNyJ
QN6ZI8vSyRXHt5N0XOaCxUduXPe6nq7poOairdIPqeh+Nn/XwhKfzGH2QrYc
jH9OOb48feQi5jy1NAahTRlS/IaQAKOeYbI8AsQJjDQPPP1PDd+Urk6GuiLN
8lLdyEydQ/HwWuZxIbNd+rwXW4zsHNOo0X8WIjL0FcVd8XSguZNAYN/w8kON
aT8otg/BoxtptdLT3HFlyssdUCxOX1gY0oZwEgmwX4jHfl6ttTSa7VTDAVH9
gMnvkPLaOxh4xMK31X3KaujEqvQ9XRuUBvj28Z99xD3RPLJeeIWbSzoW458k
AVjpEpwsVim/pfyGIgTSkddn6/DOnxQAJeW9MabtRqX8u2/5h+igTlTnNDyc
9jWYVbf1KOKfJ4f9lEd9N6XAbN0V+TOtoF3gmFZ3br06ahOESrbzrIHamxsL
+GQBf9K7pEocJjEOtLcrrLl3kOcSirVPJ3KNht5t+4DWnEe99m+/rSk8cgcY
HNmOBw8+cJ9r1zLNF1xOnCG/h93jd8ef8jS9PE3ojBPdNM2uRI08NMiPq4E5
NnqucqnnQQiOcTjX1mRmRCyMf2fcf228E3/C79j2zAkWRRDreXroW0tivQN8
CWlNv8DAGVSiN4+/vv1JMoW3QlnX7CFE0fmGh2jVF+C7T1avXUGk+7IL8U8s
WHxMIhhZDkBwn5WdWxzTZ0WKGQwop9KT/i6jb20ywrCvb139Qm2cbS1Mygsn
MO8X1ckJoZWWFflHEBc3Uu2d1QSldxDV6VhH3ZHSg6TIUlJWcu2LYN1KbbR/
Bl/f6JszQhfvio7K2pYwiq7JjoggUAvBbW1SmCQcr3CPjt0lhUMcTAu3VkLH
HxolkWfh92514q+9xQxXGO82ZVYARLJbn3Y9k6krCSLZ2AtOvyfSWyOsCl4Y
fwznyl4lMZBxRKuMettQG/eqVYfYZr+cfT64vkA1CZhuOyg/9gkbJAzVRd5q
zvBeeqiYazZqe0sBH84P0uE1ivC2dMxCeXtO7UM6Hd1sEcMv6hpg8zBh7ghU
jrzmB7UPRAFHHkePFNfZ4feKCo/dXwC35rCKU3qBIcN3ijgfF6gDGjCr3h92
pf2orYrh5kRYOOOvw/I6lv4MLhg4UqG5Kzu0bK7/DHSsLPxH2BINKC24kU1W
dJTTyXYIqX9Kf3E4n6Bx+8Y6iT+s4Bs7y76wEppCAEwKn285Hivzzk0Cdz0Y
QyoDed0zfc7c0J9g8m5w9Ew0uezNWX87aJE81ip8S2kdZX2fWgb95VUyuVCS
cbh/ChcA7Ilyh0O69r5LfPgTWAusyGEjr70Q14ssNAIzTtE74+HoaLhd0tEZ
tXihnaXRLpvB7I4RmQOhCYEFM/iF0stf5u8FLmd3UCXnkLpHGHvWjxe9FrgL
CZTlxRVHGTD4K9+1MQRnyVNsxvnGKLk8pehD+Dcn6oaoVBCwTAUQdQ3ZELj+
hEd7rxWUoHZ3v5ZKnbpW9WWdiIzxOvUdlgrIfYXftKPvAbCYGYFo44ABuPHW
F7PA/rLiA3gYwNn4Uh7FCIx8/IptUfB0r2E2rbIEpshAHmdPyfAEX12BEyrV
/D2AftexRzcndUcYW5qkzsxJnMMlgDe2WvsBPsXITCJ+HJB2v7+06oRM21El
5T8svxlIF8z8huZip0mVJ0iOrjcuCAR40U8oiRoEFYJ2gBKS7KV1yCOUdRrU
pYnjqn8Epkv2M/zsFhJhOXNYGA6apclcHfatipfUiXjIUji5vvMB0C6XssVy
UxoadVnpHmiZwTnWKyvH3iKNjXYuSRjYgLHRaEYLJbwitPb5+207AImWWb6p
qKsr9xIAVgkEwPFj5yVyZVUYAs11LgipfhiYcIjIRTW8cEhzTULeks2NCRxA
3GxeucR85T3+MwHDejEYuasqACD0XfC1z9b4Kmq/Tlz5Q4f5tiJFz4EdhkW1
d14jwGe1aI+98+BOOnH2KonvpNVrcgoHIUDH/lmAJk6Gc72cD6dhskrpxhHi
lrSRdoftEW6kBHbwqUhyHzZZSmqKOTMzdroTcqAJcMaZB452Xmz9rup3KBxm
b3DLSishFKOcdavbtrM6MwehJwcM588cJTEAmSAFeBGPZ/imuI9taevrQhXR
oxXAWBYo792AXW0eeiUzwDLEjhVzSCQ+NXcUWmz4wvkMdMtCfTLzes2jZuiL
ck1sm8Dz3VmLqcqOTqiZ6ZFJs0SaiOK2Ji/xQUNC7OB/r2WXuV/S6QEEEFth
CEm2VaySGpI7lPbyPVAxUtfw7xrbZnf3vX7OEIFef+6TnrxJoER1t/5Z7fFn
/qNchWAD/PWGvfnNgD9WJ9SkZw05eFH/B4loI5L5fms/6KOHR5ZpmwzmNBxC
wGQ/lC3y2KXkLhC8pmVOajnM4e7beYFvRMW3+KgQHy5eL4B5CVuW0zLcZf3x
R3O9T/y6vrOL6fEnYTPaWY1ndlZnjSNHPiZVaSHs6Sy8S2K4AFQdtnW+Ysf2
bXgpPslGUhMLlboG5MTiVNBn2NPIlCA0ysT1ZMn5HFNMR4z4WBCIcgxfKkyn
+tuOPofFG4QztyLsDOI1eDvwh263JxnDgo5Az3njEbRyGLcN1gdPKtJUq0zQ
aURnmjswGlUubJD24R4HXRB6s3ac3qW5LLV/QsbBnv+WrvXVXsXTsCv3d9w1
i5BusqpDxggi5Isw9hawuT/RVCqjI4IWWXf9v6HO5EDmE1/QkVojFUBiLrkN
KRYQKuj/x1qkd7OhNLdV0tHUxJbTOIULa992hHVRphFCuga9YHFNadt7l32e
jWcKdFnRDvnmxe8grbFEi/Q1784C0ew4GKCS0B02/HDR8YUN3OWSqd99/Ft/
JqKzArDmsvyz4Y9QTzIRa4dg6bUDJEBe/5vO9ENUs8dQ0de6gDkcMeo8S02p
Tc3JyNV8QMd4i6LnIkOTd5MmjSJfKCPr6izRFfqMtqzRoL036OjvuoNY9/9z
PfgqXC6nRlvjP+NU6wG1pq4n0eFc4ZiQSyQyyx+aTF5aQdlrRDdlOvl2mJp9
6PLAVmML7Qyo8mmMWQMvRAyCr1nmGxCq9VgwPJ+LQyblbCnxOG0llOAg69iH
6Fd9P9/enHdJSMmdAzYBIPJsHVxj4A4NHSxfJAIpGzp8eSaSmFEModzc+5Ni
MZpa19XJ8SoPlsx8c/JtIgexP1iTZ2dSBLR5KEPTgJJrOgrShxuYbtduNyl2
eHTZvUYJrgpIjEyH40Ll0itjx5nLsx6zZqyVDyheQUbrPw9JezrIRinMKB/6
abSfzPd+2Y9jZEiSj2E1dElqxG/3Z/2JFOwR+rGDVcXwvMxVP804EPYzanSa
BiohAdcRFI1u1eHJMYqtuoYuJX+c9UtLvJ5roxULyilAT6xr9trPmJ7GyrK7
gVNL6dbTrM8xmrbdbSBPbrO5jxVv7W2jfkUtAM950W4vXFRHVXlA4bm/RpQ6
mW5IrKPMDxxgEJ+wxsWCNZiMgHc4OfPonKVXUn0v25mYoHvmtceFLr3ZSZ/f
HN9rkXIO04BhnaX8NKqDXOttPLzSMbcLE+g4S82Lbl+XMMrNiGyIfmbFoMOs
nQmiJFuMwbujOgTfSGr/CCKXIDEHijeMoeOfPMRfxntB0MfGiH/Kobauu7cG
2sa6e9LVOqhYVEPmM1bydeEGSKopqhSeS0QCbVOIi2wjHsG+r1PEMd0CapA1
EisejCqRdE+ux+aRTRlFqJ8wg/WwJeBNKX8AYnH09szTXrY8JPBxg5Nx7M3K
l/lyNwzMaGUHfstKVzdtntf5K7k+1g4jsp8qABSHnzugQIDL9QJwIMpGxsZb
L0qJzfAMjYxkUvpghqs3iXqDGaSLgttKVGUWcb60tCjaS2CIo8jPbnXSLTrO
U94R+Pk6g5YP25y92z8UK7JsYkJUphdHBepyN67Vq74qlNfTWr4Q+OURKM+6
meatnHJ2lL+x1JrqksQWVLjwPwrIYRC+NgPIntqnNfqniY+VlO4fiSqyjABn
0Y5C5lNwYGzAH1eVdxeIJBNHlJBYjMBri3dr1+vMOs1hv/xEYrl0f8ibE+uw
r6ZZJ85QNRpbbS5rxuXdPCb/LFWYWRPY4mlzq13PfV6XkmzEMV3QOpQsv95C
Bc/loauYG9kdofSRfJx/u/obR4I4Rl41atOK8vrSVgEyHZbXeSc8pKu0q/No
SdmIt01D3/JYWhLX36tiZ1KB1WVj857zgoHYPI8Q5RY+f5ZBBINEKkm+sU5D
DG2BtysoKY2HMUbMl8aQ45LSXzrWElh0SitXOqEmmvgoC+sI5GNkOX6XoJ/B
UvPn9TW3C+S130c2JqlPVVR5Xqw+bbOcyJKS+BceLX3/yos7tJyYkSMoYN8p
I2O64RzLsJyWBF0vfH8N9m56Ay+HYywPKHC0yvLOXIRmJz/Zx6fN5gJG8hyr
guJ33wQevLYtXX8nMyaj59XlrOnvtDDeQZBG7X8gJc+rSvHlNoRDqzGqFiPI
DJcH811qQL3daFvdf0eoKrEjzHjVYDm2ZlEPwiBrq6opznbS5GEstiWvcyBN
B/8ZYBZQIZOUlLN0lLUnz0QuxsRDTL0f1/5fgql+V33Y2i0UfAuKffU+6gPM
yN+ljqQ7g9WYTm78Jla/C/+CBCORRWVNLsGgSDeITm3aPe4PNT/87ff3nVVg
NOrqoQNcN++y2bNoyPLafT/iTzaOa4UZUNA6YBlOja3KBf7p67frAwnlXddX
Zf9mzU/qS204aeJM+wEsMFiME3t1mhsOrsXX9J7dREqCNV053YrV/Mnfdrbo
rHbizYjjEvVsnM2rJfOpGEyn6R0gtoNEVUaBWiUTgnu9Ce0av7wJ4ng75NVH
FYxNCln9bk4DW7xLIn+rXxHD8EtdGIZGSIWFoxxLJ5WiMqDIq/5q6LfU/Tta
RVYSFOtQZVmsFlql7tr4J1mR7/HnDR35iBGihaKofAO7ib68pYqa+3u3xe5+
vgcsSvQFp6iE+yU/rhLxMse1QE8Tn7Beqzu43nrMY0A8JX8/ENaAcJuGPZfo
5MHYo0lHNa9rVowcJ9uOTDSp8q/+8vvdma8Y+auqelOLuGCB2qAkB1C5e4bq
HzemMpWQsUUmI0xE5IdwzxGv1tUsi6/2LT7RR9YmsLm7eMLWgTDxEvVzy/3d
c3rg4ZZS0NoEsNukO4YmvQWu4tjrRne9weui/mDQDtyIGy30mDpVpy6XyuFS
YYh5I1ZKwVLLXssgZAP51YXgMHT3/b4Oz4+jQXcenOGDB/51KSGmIn9EAxvr
CNWC7eWtKbGJvJwmHHvfH8ps7ntUDHXdxCMcTOMVWU4plD7RcJG7MkAhVd9B
w5frvb7cV1nUiQqAW9+RqbvqOyH8M9E9dCM00zSHR0YfTcUkyF9LJcxiG25w
hW9x0xZ+Qai+aTFbUMpWQkMsTv3EIA9Xd8qgqpxBVyIg2FjHc/Gdz1d8vzEN
Hwxr+YmRQfstkW4dBLP6b7grncHfzxTMi3q+ZakGwXjDQ28hhM1vCtuNuuiT
9NjvAEZnLEXRscLIpcy/jGxX/h/t7lP/vKeBLOh9U9BcY62IYMuxIU+jYZlf
E7aZwXyNMdThgsiCrdV6MOJIZiBYq2ERUGV4CcQoxASumfrFQJ0QDQLpeXzq
E1lIkNZd9LlD22BiFqON8T2YoQ+fZ+5D2HJK7ff2ypwNbr5E5UH/tR1fVGg8
ssyVAv/vrSazvgR7kagYuL72DuxTupYg7Fuqb7wOIxLSFZL+nOT0peFiYGwh
rL7DTHTiJqQnXg+n1Gmwn/QJ9qjkgs18NkuqUG0zQqB630a4bK/Yn0iW7sHj
lrEQxOkVTdiicPnVPnzTT61Yl5R7zBAXkJMQizMhu6Tw+6puz2amYDAAnPXm
yVwrB3yZs9VNhRv9ZlFvZRWMOzL0dyHpW1OHOcmZlFyWTOV/06TT68QuVblJ
VZpZVUHZFMSe8k1hzBC2xrcjkCngP5kJwhXewpWq7yOj1gUU/RAa7AFratN5
0YPRgeXeaF+CmQ3WtBqdNP0OILwB9UMaGDmvKTcKxwCitG46KI7LAPAZG7tx
c6nceFYUR26Nz9vsd59j3UUOM2uPDu+8vSyykoUWcqZbL54+rCsNg+mce2uU
xF91iS+hGPaEUzdvb4jwtBvHRUbCo6wX9dT3wfwkx7hm1YlR1yfgjbfHJ6f5
hNeZvs6sHLPWrDphYVsD4wNMnQyAi5TsnnN4Bqkiw7QwMplHDDEzgcm2Xa8Q
m7UMHQA5RxQh62omB6OnpiBtXXyZW201a8QsET7MZ2DZHl93zNFK6814pnE+
nryZEAreTnGrUMDfdHrYsiS8YYO/pOZbWXmejZZJBv0eBmq9ugWCtLdrW6JC
JcRyMu9Nn0bAoP5uE5TI9Q4IKOvHAKmASM3LbKfkY5jfXEihTpFt3DwP3U1c
6c+3DE1pqSfrlQOo0oOHkrnFuEG1FPdd5M2WOQ3K/WnlpMldNt5GpNfZv0HQ
5CuoxmOY9vZ7Nf0+CEuFL21n6G6C3QPMgYq8hI8botzWfuHnF4SZ+OK4s8YM
50eedhKYLMcU8NuFG19Wp16tOuSE85Om/CjyKj0IP1Y3Y4ogNARqYhKjNAvs
E+SaZDk0s9JTwM3rwYb+ii0uvyW6NHDlNYo9dryZTlYt6iqF9Dg10fd7D9xT
o/M0jRd5+3AwKRTL/2vALqWZ2J+O0lfeD68hVRLNcPQ6h7ePH8Ocd9La90rt
x6jCr+moIYDNnDfRGZ50cFpJw7U2yIh3b7MMjOjpNk33P00Zu7LAN+MVQ18S
PLtTd8nZ6Bh9bf0lZf6PZtE2bVXz46sUe7+01WcxeRFSV/aYZDqgpwm9WVaF
alFG3mu+u2u9fo/oDzFWuOLjJqlbfrcAbLpkjhFFsz7B0ZViUyPPNYuphLCP
1c4t9D/tdyfD2I0PTL+HUqmPo/TPDdhM+mZ29iLiNoVLlmyJATsfqbzedfBp
EeqKSxo4YG/Xhfo4Y/mhBeXeGph4CBHJUipQnEzsFbreXYagvl9KKKXbbYAq
wfF0C//p3Qc6GOUCSUYVP+4tFtMRDx70VOM7VpmchkuWdfthknP+YCBISSjK
W/QfV1zsURNCX7mGj9hVIj29dQQGFUfOz0gK0+6y9TjlsZxjsqmFJMVnToYM
V5VN9nbmRE0qzuaRGh9klDZ91IWi3rvlyVF3ikGoHIZNM1TcfQZgyPcku1u6
z3z4qShhehGOfaVlp0Ezz8I2CJGL3BhsWOwF6aKSnb2Mq4nafHERY3lWUTMc
tv3ncedJ/CMM0STzCB+z0lzUOnXLcuflGAJD/nhvjerJ+tXx9MwuUcQUrlHV
huxcTYo4XpRE3YzHE6ok1ndXP45mS+ON4xHOlWg05O6mCzDJAA0Xd2ZIhzFq
rJub+tNm/olItapB5OxeJwDi2XNtd2zLdc+bzEzDRtz8LHLU0fX5KalYcJr4
Vnj9SgyGdOuf/PwMUrJWeh0Yekci8uZaQ+YwF4riCmzA/jA97DvCZWGf/XKf
0r9N5D0IYF2DMgk777dzgwy1D1sINJq3ERr8gJF9skNNB7Agoz3VY3yKU4k3
A4I+orfoz15j9tvkoo0W91y5Qi/h2PV/4DHtumGx25vQgIZF5VK9Yg/sE8/4
m39L4tpqkH5lYqBYJ0RN/cxmAGhYsLdBjdZEGYNSBuEP5VN7uLHpjv5BQSR1
FPcGP0qLA14lcnkOmCNrVdDp9KkAwCwLbxuCaUiQR7ZrQJRkq69WP+26oDPx
YUvN2lHCb+jsbIxOXUGpoNONUYJO0ScBVAxBAGQl6deHb1VoZ5sy9BpILzLF
foLUpxQBVDIogvVebfi5s7S/4Mjw8ZX4PEqzy0+miAcKv1Z3aQzLqyWWdiea
lIiMBf0qDhIjloqX0jFkb1XNyEMm7Si8D08D+CzWcIaepZT8L7TFRbo/PRwR
tJjhxlaOISdR1IQbOPRl1k038WmEoWaGE5J9zlMZYkPOqxfi4sz9jFnnvgKO
grLy/4Sj7X0msZzL5I3tcuRT5WhmfB/7aw+30luIiYpQfd4ErtsgmQHPOYOz
akhE9H4jxUf0pZ5R1SjTaiZTYYsZ/Xv4zHe9QEOuzgsYNpSY7k8ySxC9b6BA
qg3+wNJcJ/5VcWgN57V6yNTkMRzUWSRDzNf3s3PxnGSwtOqPVwQ2uCVqahxu
2KR07Vd1AqE1V77w/NLUa9L4QE8ESvy3DTp+bIrwU0XHhP60BL9S5bjPHicI
cUCa4roQ+yytUwuoCEWmtf2N0Kzq2F5kVWZCKoJd7IQ824qWSPdkDOk0b/Qu
1uVR9j7Iz/+h2+aAE7hNDE7bq86oKwhXvUNqWqzDkRJ6WLNSi6Ce/kaAFY/W
2ZK1WqDREkiTL/Z3gK+pM1tSNL3AuU1XnhSy6OAifpc8wth2IrqBq/eicS+k
kVjGPyGvdZfYlLnlRGNRt7xvp1G2sitf+Fr5ZecScpwg81tpAwNwMTFWB5c4
14gA325OC9806iB9wlshQPhZuNO2omnWEn+q8JlfkbB6Uhss+O75y+ru7Uz7
icGYYywCZ1OvH6Dz0uXugICXUcXt1A3kN7YDwf3Qt5Kxau1TnOJicJ3cXNQB
HTpSR2KGo0QjT+tfin2a1fX0NvdNJkG8FC5QciBERMj3M3+m81PK69H36Nel
Do23nFed0H4oYbVpGhZ/bH8a9hTZV/ZHyOYpsvp3/HHGDsLd5qqAgU1VKvll
AxoPkSek2jG9rv3S45WG/pGkKdP/UjCM7YUSVttuNEoILOApjWGHrJLychoZ
soVChhrL7eKLBjiAAFpDz//CKzUcrhP3XIXgiZzw/dnnPt6ZjfhtnpUXFGN1
5zXKCGvuCejVa4GnZYRd+ErU+CM9WmR5MjPz740bBj+uQ3nqup9l/5YmDpo5
KZ58lMK/KOd4udfuanGiBlM6+pbONH0JKkHEZJC3/YquKSPZKN/xfv0Lhcva
fRIZKzUWTmjbJN/a4HVR4mtCl57YVOV5HF3MIysM+SqT4RnmQW0N9ooFlf7j
uJijnbWPwe7lzbGop01ypj7hxv23GH4YcChyCL84IryvaNFldSfxBjJ0yJm6
DxnHAjyKuBEjqh9Mb1VmlwMyMu3eOfDphLqgh7Y2rtBJAkICBeKsA/HMncAl
ReLoa+IHZhSfHr3lRgEBQJGjgd6vVFRs4DzQCa+HYPHH79T5gYEhh5/CII0g
M37amU5e7VIqPxTyAo+E1oGOtYI6TRssT8HITNkWIvU2tmI4NnVIyggrDSvp
7ev3fcDeELNZBb3fWI5l+vrAJk6qj9sENeQvpPpikfb+uuOtWcV2Kfi6FOP6
wHIFHOaAxLV602vukS+xGYFhHuwdEqjf1gJfIPbuTeM3mCq6X5K9skh4cZh5
xsE9mXejp7eRTNPbI+ltydcGMVZJHa8sZhsKqduqyOR+Om2yQaXUAp5etbot
8l//73pR98MSYUZc2WJ/4r4HcHwyL5OD8xyML1DN4TgZYt3+H1md0vWjqYDq
ga/mIskYbHFM9xyh4+xoyizGvI84o+TXYIAt7HyGc0ajdIzsP2E48GHTCdoz
zWONXxSzRrYQJAp61G8oxbg4y6fh2xxDl8ulNByl6KvF3vLUfIF1dF1B4S9e
nEP6pjTACD9O/BL4YAAFp97oL1qQYN4IWNt4Y5zlfBIEIYz4hUbXwKnfSwd1
j/pegJxR0FDVQVwHzM9GwNdpUWwG1wpRqYfS2X7V2iwB+zhMlkF4mhfWIbVB
pynMn+2zpgP8vCm1pnAldqrW4GuUiBW5Up1tiLGlC/GjtC8d/fYdVrMW/u2K
RfPCVPAk197JbfVmifvR+hbRgXyoDuf6BXAsepytHbIerQISavvZb0X4NSLT
vSTNMc3o1pbdfRVFqn8evvb310VZ+eFoEP5214e0z6AvNwjJLLzzEaF+/mIS
SSEnkCvgbhnQJie4cf/paxhIqQH2QSMpRpXNnEs6rZ1G8h6LJNKSHj6iv/XW
s12N+75E/kXcjpGIHLFfxAlVvy1vF8FQuLQ3VimJY6nSlz2u+FrgfEco0I/6
E9Q4a9zZmSbcz6MngqyzsNnOoH5MDs6wz23Rd7hKBReQelPsEYaLwBOrmMY1
i4DT+OI9kqsfGoQWdQqyFuAXn9ASP7MNs9eFxe+dfyUgFfyi3PrA/9euKwI9
hSs2qSEhp0yegsakBDwiaHdBMlWYrTQXzsAe7in++cvSJE6JJE0RwowlPM7k
SYtFLhi8SUfkx15VjMrQ4q2UyugMSKL68/SYEiOsgaDL9cQ7byvTbMXkLb+v
iZ/VLAj7JRvygS8uFEPWpMr+cLFHsck0gET9qJRHgqsPwe1zSBvsF4T8LNmU
/Rb1g8nr7TMcFLKi2tXsaQ2ZCtLtGW0zwKqwefbyBfioQeeZdCd8Q5RD+NRw
Az9kkwYSPhz3qWptH5hnDIuyIXwzkX8KOiojPjmo5y60/4emWoUbOica/ftp
jWF0pjV3fi6SF3GY+u5v3kjESvos6X/KC+47jeCbRy8vcz72V5N+DAj8w4ey
vOtYwHZZOtRWD30wbvrc9bGuPusdn9PqTd081K/VZcYQ9M0ed666niLr8upj
RYQX3aEGDwqZwyfzoRcO3RAnTpOc8EWG5K90NnNXCwWLNjxOW3h3Rd2QRaMJ
F4gIc8jMyyAkNOqUWturf3x5/t6q4rLQiUWyg+Su9zdI4dmVW6vKCBq220rJ
KEf0du2IXaXJm31mTh0NhclGwqvgwJnmZ2D/ciFJt5ziNumKacSQ8yIJdiAv
8xQ88GkzX1WiG5Zg85bW1h2WC/L80RLJnBfQUjP25XT7Os9+lmjRJtxuKqoA
ZvXJFnXueEKUM0u7MUb/s4+HgFt7oddiHxuG4qA5wehfMibIlz8XgLVyQKNJ
BjGQT7X61nBoMePshU6sqwbT/OhDu8RzqFzuyI6+dWYmwfM9ouluQ8RNZSHv
t/3PpfzOI19IzGGeqcB8DGlrGQEFR1dNuaEsyYbmD5jKXvIJ85fxj8rw5o7F
zVDLUs0IFimmsb6CRBK9bRXMrDVa8tdD90LYbDEjjGpj+u5nEZUMTmxQW3tx
c9N3rAxT4qGMH/I02N3WaOhS2GldnNCdgipwmwXB6IIyOCSr/Djk39bLGmHr
S1A2EttNyNX/OcGwYVY0nhB0mHOMp1DcsJvapnTbRzFVM0RRgDDuAVOLdsgW
HBjK5TclMAQv5c9aK7cbmnXElujGt0Joo8JYiBHgvpgVzdbqNv2/wcR36ONk
ikdZqhEk9AifYq9K/Wzm2d88prfILQ26WFuxcjTyaWX5IwaL4k2gCcNi05G1
hO0iPGuwDJ8ULsK8gZB+c1pDR6X0gG3JsgZ7kM/ijGNWWXf5PH55S9CVbDzq
Z3LcVNdVj9jftP1yZuzA7S6S4/zQ1jhbW5C3Sd3YhBzdSXvDrnRGD0IX+bg+
/uqwH4cZ+5j0ao47Zzq0KH4M4kADs3AYrEhaGtXbdQHi0Eo7JevFD5wN4v5l
miNbo2mekjctyCljZanAl32U3Ty1WHDeUm7DT083gxyJTPSDBVxB3csHmx1H
ITozyyRkHqJ8Ov0xDUrqKH4Yufoedlv9jNvS2S4exO8sc5NNXraxKr5sMIW7
1a7HGvgYRFvN5hAQFiaypcOGUWuLnGk3esp33pJ9schEu7ziqX+BKNDr85XR
xAmi3rz5CNaVIuaKb7jAu6wlHw4A9RYvwRAcsWSmOezhcdrHPaDZdu1hUKCy
tyF5HXQ/g7Qy4RX+8YG9J3otByJNPXP7wNUh6rDwo5SDJ8cidj/6rj2zhmzS
OCTp9T385M/HITNEnlu+l38f8j750NP+TYibZpPXvCz9eridlJ7tAE55K8J2
hqEw+UQZ4AKxKsF+81tYI9SQ+q0Vk0fcjBi+8UJ1lQ7gUiwY1cnq9ynOY0qT
tFYsWumZYIQU+1TKSp+MrUcFCO8spFjc/2YJC7ba4vfSdt1zEAWjonh/H8HX
B+qOjFnerDkRuHU79zN0fqBQgtwH0rLvf75c0RvliX89kdsQ0P1tHmN9mo9k
gx3cX/AdzMZh44700ANvEHbsiMHMx1XR1hws4S0Uqy+Kh9N9IZ7brQxzxmzN
xyHFGB3tcx21goJRlTDEmvRXK62Fuk9IRkhh78MiENTV+iS5Zxs7OcjmXVL1
k4Fo29b/CVkVkth1IrCk5gD/pcfZLoaIQkvCVL+P6kPf9OTjxuC3D6P71M3q
tpn9u9TeviRrG16gUyDP/DQgK8/tKfbkl9pDZhm25NMlp5LzzuQqxp4jy4Ki
xLnJG8z8zjfSw0yW0Yz0j5QcBjCPrneSqBQNJkRIQq8AA5qahOS/+P82U7Vy
dmvrD3Wm5yjcsGhFYnHYQfjm2rGNr/yt7Qc7ckMd++TzjZ0DL48E+x8RgXQ0
Bk5DtA1Qez53TcRK6FMC3fdE5A154v0qYckDhLg5mQSxHeb12zuC3RJMIUbk
MQyzLR8BeSg+zqPCc2RRUgUYTWO+H4jEhmkdSy7CUuV1/XIgSk/Hk5XafkQQ
QXkzSCiQ61uiuqTLPCuLESRaX9Js0iyxBxAeIQfnkMTma9DRmeF85DhSmdck
9Hdntg2eF4XLezzVxfCi4bEbI43Tr7+xriGJ9IvC1GrNQCg4Uf43lCnzdX5i
7NizgyiLKx3T/T7QITaTZPPHXexg0IpEX/XNuTyvO298SenY0H5LqFISJHP0
wOuaOJ9yKJcsW5dCUNGEsli9HkpgBwUIFDBs0edZojvyfTbS+0sNPGjKQyE1
C8Tu/M92Y6X7KrBpLNkvrUeM2clqYwyIsAMU6uV0JZUq8CdAsWj2MNje03zs
8gy32ZLeVIwQpJavwsrycOhL9zDqu9cBA0Hy6L0voFX+jyjIloEqn1XD2WpW
+dM3CqoE37iD/ovoqBuDQjFsu8iBFBA73IoZzlS167cyvb6w/olXFKW/9oy+
txPAg+zXsUry5QnaeH0/y5hRSBBWKAHGpnLSyb+s4uhmm5XN/6CcfQ8irUGZ
N58UIiyrzY3Fl0n8hvgBHqwCy/wa6p81eBFAlbU2Kb3tg1guM44ZrVhCxXem
1wQ1Z6UaHrLWxVavsMHBj2n3FXi1JJsTse1d5qW0hwBFZef0iwuusy22vUZg
ex1O2/S5v+TlpVMpNp93GFdMMBqcyEU7BP1poPgudQQ4NsNbrvnihYh/9U6p
klLJeyvf/Lg0MWX0rS96f4nIiWXEWFlE/oywyYSA6cL4v+VsesFmVNbZiDDU
UUXu5/K/MsrYbjXOmytajEFwY4LY/gCE8O4SPrNYcQb0lQpia4zODjyXCQOA
rus+mI896+VF//8XGUf6yG6qg7vx+BfQSA5FQTvTA6QOJHgC1lWy//m/Qwv7
Se42ve5DcQbBMIyrmflVZhEPa+cygAqlDMaXl3uD3kEIvIxjML2dzBh0/fFy
BL+flqSZHJ+uIbsMXqSsJRoqew5KN95ytnpjtGfzP/ddM/UvikwwEORM/81K
xI3iY1ScW0MtWC0uIj7Y0srLneB+q+ZANFyGSOj05wlD6sNGaz9/Cpcx9vZS
6hZJrdsia0mWwk5LRD0JFhSk7CtjclMOTBVhAm3GlHexbFy0I44BP/vI/x7r
KDVvaUdB3u7If6b3gaMiWx+ZniXUsQpB3Kpe5shO7+3F1EwtoTLz7HjlNK9x
jnJdzgMrQ9KZIok/8xLFDaqXd031ZduUt8iRJeBLkwFbLXOFGumUy+RjJ4e8
ozbg8LWet+X5eU5zdtKgQyiU84GVXyOX8GrORXqC39Y+Ubklaw/iUefJvN2x
YgglmZ38/SU+IJdisYaozpv9kOEWeWJxnXuo926Bj83STRRelY0kYWzutKOp
69Sm7G8LHPLuxJCieJyXr4UtQwf8PjY1F5nAGWIgrwjy7w4EsQ6VbMyPRbPN
rjAcYNXpEv+lnmNIinuFAOH9iEKYa64R33gOyMiCIog6w2OsGdtgYnStwAgs
u24zxMbaNfe6KOy9n4ZMrgGo7QWvtl4KRHDgiKpcC5BGm0ZqPFpXHybFRxQz
gBBmHhJHyPAJwB/Sdt2Ex8dZX6V2AScfgcs9j/SYf2abuXlA+1QF4tFEpOXx
/Y7nT0OaiJSAWYU71n5yaz5kERZHdEze7EpdUrB41Z9SLjsr5jYFFLdJxexJ
3eb+zR/+P0cJA2yJv861HSZatp8iLrbzMGlYsbyI5zukdiw9SeIR2gBIRGB5
rcH/EJ4fEV68cFBe088CkaUuFXsGMlbF3ciKlTJya7Ffp3P4qAoP94aeFl5t
Sgt6wXXu3eTlFdXAOj4quJ3nRK/PEQiB//vv58O42MGZBDvleEXaFQuhr4kq
nBb6PkP4vszOmzchRSzRu1TwJ9y/E2+8auVpaBqwApcJW31LraFhJGAA3Sde
Qucmbj2Y/iuJvVv2MmnxaandQvMLqgc8RJk0vIaBOErfJAuPbUQuKq5FBqqX
T5+/cN1CFf6+E9Uvt/UR7cEqRthv9HUkL3YkRk3/zvlMBBzaKgqwdIgH023u
CYhoCR0M9yu0ulAsOOIxeE2erDFIfxTmqfMbUTRZabGLg3ICuJs5vS0TQgsb
XW2hwu5OSmvmmBULtmxsGpog1fHX7YwchMtyCXbwvNgNOv8s6hhPOGZyvEsc
AwQ3tDTTPiqZroK9flg2LPgiMH5wAyRS+sg86sVUj8KRqq5i+I4nZEep2Cdk
p3zjZNQSPuRI72iLsOsDzgtAPWtK4tkCjgnnfI8yAaT0eNg4ufjhe0cUTRs4
9TR+vYDbHWUyQDxkqWDH2DA6grPjGcdkg+wDP42mV3FGYAKTRgN46l8kJFXd
uKH7XmNSNxcYqStg/7M9uar2WstM7GUFYxleZBY9R9b1WYSyhkW1WtWvG0JT
DDWP9TC1KKIOj3nChdJ6bXNdz3wQV0xjl+qIP9FK2m8k++OaAoGc3TfSuUCn
/lLvJu18Phyen0vjqxq+rhitl6QCMGra0z49C9EKbb3AlXii4H5Y2nKjWq4i
MhcHJUumZmo7qJWLN7e4P2ajjTW+wuDyVU/HqX2I7wliE6rj3t2MoCtLnWoX
VGzVxp1ClQMONfB/clQo9J5EbDt7CTSN4ILNty8LG1ihnMf4yGI3PIheUQBc
HvlC3w8VC9EH8miIEuYZMaPjCCTbavQN1fLcnzKmkR0MBHl9+czUwoCUZtDP
FtsCP8GwLr2g/qFovMNq+t7dAdY7UnT22fJwGo7vgx/0NU/7Co64JGQNZVOU
vLEha1PYYeFkqBip3FGf8pAIEew2xr67ggvvo3njGQUEPoXED3WHtHacZou+
YLX/XXmc7hdGtcw6dnKbl2Kpezsw7KfovAZ9hEGYUUX0XCkHm7gVYGuU90EN
uOg2mX640RcsT4xTakmNaDXQTeEKw9hm6M4iSPRGEBc19v8ZdxgYqesZoQwY
zsCXZw5P/Prbd+YhdgNTTAKNV5AjvqvXN0PHwjtLH4KcN3dx4wknB5IMlKEQ
bv0sXcPqQfrihP2HJco+kk0c2eJFA5aQbeSPScSXfJhofg+e2w9RvAA1wojB
XtIy4NV5ANlvtwSxyvMb61KP24vykpZnLvhiATTBIaw9QPZhxKxQ/i/svcCn
tASaokU374LrN2qeYkgMh0FBbYhgfSo+P0qUqL2juJNektRMhdrdLYFpnzjR
uUNiDGjgNAZ96WPPH0SswflnAEQBA+/4juEAjUPclW0wMCg1MkZTkQOzm1Ka
OxDJxj0rJe8Q+JMW40i1GjizwHklv2jzp1O8b+1sAMRW/oBbwfVImwmiVq56
Pcwql53zPfXdjWD1je3AHnPYltOtkrkeIyJH6fLCsRIKXFlrjCY9YqCinq9h
oEVTqOrKWA+RoBz4Hfp6KKwFRHPcYpJ28fDPjS2KHuR5YPE0SzmL4FR4auEH
KySZsAgHnpRaLI/Q83ivE9UUFAFdKh+FvBZj4u129ZvNolScOwkPbAfIZsEa
nXEhzHryByTF43KeRKbFTFuZVXa4pqHrFInwNvwKK+rVwDhTeIP7AA3ZsB0V
3gyw/jHDdidFPU61l4KOqR/NA5lzL0J8xpw2CYK5oQkSTYhN4+g7HlzQyoX1
CidrxOpL1hg16pH2JPH3fQTQDk+7vJpPJzWVuJPyGBnDlitG1WVaVJyIZDBO
rVcC0RG2lnQRahA1SdXFo4LIR1dTJIFiEJI/SA5+5T4s9NWNJYoicwq2Tjcg
cPpy9qSdwzgsJ+fu+jKr8GK43W887Pk6RjlBASm0BRcWqNrwPo8hhSGbG/Bq
LrwctKk4QMcWiCHxtitWa4954GKddBMa2rGDBuZ1o8A1+bJGnLz1mSnVVufh
PVFCKZr6XXe4kJD/cS6tMoVTrh6az8bG+xryIDp5kV4lfY5k09a5sIO63ukS
kGU33UkNYwXXx0VwSrxS10PRpmx9z8N8sAEn/ADqifp0mc0A+W1uxR9Z4wLz
8kRTEKiawy3/J4lNz1jfCQHQdSiK3ULu/5DgbKX6uOdx525UDbAGLinbXWda
mixaXcg/iS81+oaO5ecJ0rXnm4tlsjN+xfdmXn8hsHHNLBh9bJo96uvI0m7v
AcwmjQxmj39RRdwSmYaOTVNXZOCa4xOTD32aGQOURQ/tgWjJykSmWWb018Yv
m5bTE4fO42P3GBO3pDFcKKZKrfPy8832KGqMK8Tj9vQw1dsl4xqzfHiybClm
L0CJpIi04LeouRtDUghgMtQIiY6iaPtiC2IurM8ii/XV4gipE6jm8eIhcAdc
0r2Yvocx5DyPgFKsiCT7jC95JOGhSjSPcDYU1yrr8HZGsK6N58O5wAo57qdl
SsdeRwPvOkosCSBrpPbkhk12toR7MmuihOIukp5JpnJat33BpUWpSIi1sULK
aWa6tefeu8jnmWFuNnRRNkcV3QgoCZP66Mm+1+uZ3DPruvxRaU3ydYAX8JJO
lo+Axk6JQgsREHTPTCC44AJFsihCEUt50H/m3pun5qmfrbhnNZarrC7cLowz
2pt71RaHZpIeAaPxITQv3sEJJq3iwdPYXmirRHDc/EjXXThSsZ95H0GP3fon
k4hLU7OaABGqgtc5Oj5m3HteZ5pXPxp2FpfY9heU5jCRFySvIEIoD7ioRyGm
GOtjDeXZlZ19uigZSL6hcNqkCt6X2MqC3C2iSJb9bpxQFu7HGuYRnr27ImLk
Y8x8xzZ6BwUSxwOnQHzdRamVtLWSKPUged+bOyxePmU7ABrlHfjN0jUe7a5G
3jVXUcslG9cNx9D4/oI7yiSPYdsXF3VDYErGlEX8/uGhHdh+kjwzGcZFF1bs
29ihPiRJg41ZxBzDBdU38gtpDHjP7Fkie5Z/9WKhHK5dSIBjxuSikVSNsShJ
tP66hgdiK/jQGi1bTW63w6dMdqmgQu9fofMUTs3fdG3UiprswY0wrLy8uKGb
VDSWiRhRRLPLcRuTPIHVkRQxtjjGUr7YR3jOMIuoM3NE6kiSRdKT5c369jFQ
QFTS4fM12TaRYzYYOG4KCNnsxcva0AnLUTdr4AF+dISFJ6rDNh6niQE8xfcl
YeLLo+6FEcPypLClpnaDXxkkWmECpKt2WarDdKu/tvwyxc+UozcQM3B9vequ
cnS6n1J3waNNCFrmEpEwY3V9LtwGWOIGjgU4ScT3Cdupp+GP8oY297Uad7gy
dDoINbBxXBeGlfNNlXiNz1dZiGEpXw9393ck36nr+R3xcRCch3GiULvJkynp
K4oBQbUuPayON1GGg+auh6HyqSevl6Ykuss2/yIDACbCyfZxaosOgrSyEl9Z
JVEmCZUMiZyc1k/8IkPCpRRw4euhoFt3GKGuTjYBx5qTpjWBoCsnVVwZ7HkC
Uhp26VknbvrmzdwPlgkZ7rxv/c88CAOpGXbm3pHYquIGgAxvuk/8PFnTNIv/
EW27LTlucbEhjFn9YU88pt6eTCnM2OYQ8bTfEZYuk9V9DoXWCHC2kKA37Lg9
z/zxHZeySWhoV6hmcimy9TVlHcnnXS5jTNe+0aWaF+FOdNI23OJpBRLGtyIx
snxTsaZcaZpBTcxxLCQTsprzYzXl+WBriDaoXtJOzjjO/mZIxHeBskxVdhVx
tzZKJGiBg7Ixn3iQetj24RsdIsczlM2p5RJqkfc/+yFGolB/S+7VyksUYSrZ
u/PSpqmlirlEXb4jH9H8d3FbEUMXuoPq+3qf7seRs8PcQoJJofpKGHLMEmJM
EqCXGN4/qGgAFPAvsTzoQHxSTL5u6zHAEV5l+VTt4f6MjdyhuQmgd1dmKq3j
NrKMrCqtwlXUrvGcDL18oM9XZAz+ecqUOSlzyT2RIxc6InEqo2HjAYPu4jd4
5DWn2Al/Tw7ElSImT2Okpuwv4YlU7jAkCB8ipb3OFHwY34jATpuGUuwgbVjm
UpcfrOVsQ7C0VYPlnrlmLBeRBjjk1HhKxlm3RXgiOWNCMF+hq09K+Ddj7JJa
jZp7YRoaTMyatVq1vhI4FBKJ+dRIwojvVmEc/jGAn1EeDXEVlXdHhu0m+M0T
w8YI0buUzoE7NT8yO8JAlPb2Gx9v1opt4Gb4A5Tm3gxVj2jfnEYZEFRPq8yO
pbGHNEyLGGJAlbu20NjLe70qneSNXg3GG6FyrxprAen/Qce8ggs8H6/amjpP
iDafz9M5YHKwr6q6c9iu6MYfELNCwQV+kDi5dLJmRpmaMH4kkA2G1O2g2EIX
prQwE/bZr6ueYYaPXFfae6ZRh15ejMmZOAQCbsvojFOPx3nGzh61ki+I3qfA
un5IZM68vfmmSOFkw4Nb+nSlcCygYjLIwYU4RdkFO/p3PWO6yN5H1DENk7aM
6uPPFPbkHiDs5AEh/o5PtgUUsgx+Qeap0VKLWCXCqPi2pWQYeX43L1zlKm0f
jNcdlfS74ZsQ9jTSJD2sXGc3vBiq8hNSIB/f+cAFHuZaLxNVSKwhPflLZO+Y
XRZwIIi4IjNh4hyF+ik6J83+DTaDcUK5PAXtumxx2KRoL/G9vljIye2es4Ey
dtqlN5YR8olF9YEgyPtHIXwusNBTTQ/oUSd6VUUh6WoXEC0PVzy6YbblDZL0
8ReY7zSTcMbf3Gk2P9xCJepjBpWGKlC/tSb2Z9ZGnpghqSZCASgnCsA8H6aL
P0uROhEKIq13Yy2ZDQOUNA4Y2Avf/MVZsXLtk7fidOA01wWL5k0pWSxtI7Rj
zmgfvXlJGZXDRca/ZolNSZYDdrhPhmYViEupm40i4+d6s/wOHyLh8KoT9L8h
9nlHfu5dACH3xZT3cjzO0j92PZHfxAyfc+2N4lWzdt5x69pkud1drKzR5cTk
4BiXzARrKERuZLDfUxXlt3zXMQRgpK/badeG+7CJs5vkr21En7wC+9nNoiIg
KcBZ1F47LbJvVE4hEYM2SJZ04NG8CY7zuJJG28RqEUX9PVRKmJFyBKa1ltLj
mifHmk+FYZVm4Nf6zZ/UYMxEyK5h+wIK9HXnX0WPFftI1IGS9lOgbzJ3+abV
mL6JgvFYBREBWCRluVEUUGb4FtLaLvOgz3xSeif4OsRIrsROcGQb+0JS6yfr
ZsbkdbZQOO/vEaWDCiJMez15Rtji/UN/t55Q0MZXRBt5wJ7d+8P9BXhJ6yjZ
kgRkYayNA/FoHOPIggCKxmZTfN82rGlGNg1KrQQcd2im8uWqKGCNmRN7usDC
SqOsU7FILSZSXZvk79k+bcHD8bxKAnEUm8Xu0SwQsF5Ehc2geQqOmTbuPWqG
NJglNKfVKIyB93m7N5nrr41l6UY24ikXWlMh2LCeS9SLdYd/TXszoFVHxVvG
sWoeZ0Pk5WNiiusOYvXI8juNNAjiApuYqNA4PnTLA4izQRTlvmTQZ7gpDfGc
fbTqh+BnHKq1ClQKYnb2fYgZcbDB2lETmQKoorU67Vsff2CeusV32RlDyAWQ
8dMInngWW9tVhpy6rXBWp1vcGE6msyUuvM6sj+GzU0ZroUp7Ro/r4iJWObB4
92p9hVjmGwAIYbU7RZi4Wvnusv73aD0UtTy2tS1ijv+bp4tMKI0VtcbEY8uo
x9Q3KQzbGgh2qVSQwA+O6P+mgsMFcSiM/y2mUeG0xAdzQazuzaOw+SsvcMYr
Hi7v1JyOam/pawzXm9V/7D+KeiCEGyM7dWmAO6ZeA6kH4Gho53mpIrv+Px/C
JyrxIueNkIy8J91Fy48B5BR3k9r60byD0dsgOqY4FXVB8HQc3XW8Y52WUCn1
lfHHrfsKu11cLzU+5N2pxrr90MKi5+PBh7NwDsfDC8L2bK7rspBmOh3EtlTd
+S0t/peTYvrk340CGFEBOKdIFDCkFFtjIjgyJX5oCg94OwcOeqy5OVgKLkUk
BRB/JVMK+HuOIkMM9FimaPtciCrBL/hB8oeRRng9SnSLgxpa58oLqtW8MhRr
69HVmewnsB2b8A+6nSLK4fNux/7lnolGKi7DCMKu4ui/PRjlKeGej//bxc66
ieufIxkrbOaMudSqdG35l3+xbKikc4rycxsWrKZExPJ8R6Lru/9V+BZEP1rF
aVyFhglEelbt3jOVGuc5faDEbJ4QtZTO99Mup/V9yOT8cQ42TzftnorB57OX
cthAm6yckdvWIRQ7lZLDbywZrubGEX6XJLi4G9kzEYl1j7xMZ5713TYTIzb0
BXc4FB0NNWawoBwjrT+YqvEMXq0ybbon5Jup/PrS5HHvSoVaWS8ZIzvEOLY9
QTSuSYSQ6GkdBJgHLPXU4eELZO6l0b1nDCdB3T9dtEMP/ZRwBz4czOCMueCV
FSVZczJIITgN+TS4y7Uczcq883/nzPhUMvrkNz5+wDm12VWBoV+4lYKZSrZD
sZBa7ImigfnG8f3C4Vmeu5HOlDx1yTLGEoPz3M/AbDPEUToTzMYwSepquazb
C7ZKX9ZjDizddPpy3awIah1nWNDRMxdyRjDbsomAquuVKOFPRRFWRWdKPFM6
sMJs2xNJs3Ntfu2IKV9FPOPa8pQqKTu9m8FH3EMKBouxthDNaUAbq7WYDSgi
oXj2XYBAuxD/J9QvptGf8cn6pCA4SaxeEuKDqU2sJnN1wwm2Zw2wIA74sVZI
+9t5yy5rebVo+QO73mW3PFhjgdw4nPGbxAb0LHLPVX7NdE+y1GhUGc69rbBc
Cz1ZQKh2hj1a1TctTI6EeGdylZ9TbeszW3FSmcJQNz8o4GvKbG5p4JaExDsg
sOQCJBVe+fy3YkwgqW9cYV1QnfqIYUuHR9Ble5rIXPg3+pBAJgxWqMuedSGW
NKU4vzWur8+n/JWi0cPTCIaIHYiyH/kZer2hHXL1MlN5rPSw+dZKisk0lB7d
cSM7zP4usZvO0M4IEaIQtrvEU4P3R3kBWwKFGjiZIktxlQ+k5U4uO/TfZJms
AAuSB9MsB1Z80Qxh6N/eMYpqhr1ZBPfoo2/mm3dDX+u5WW8I3YpjcgoiIaHa
wFME3uoWXqCqhq2OQB/qjLqBf3Ux7Awvwu/vDHO6Uyia692Oo3G+vrlqXJJe
viX7E1MNCvwkCb3t9wx3ilNoQbPmUbSZYnEupeGmMUj23McHWW0BjdOE8Tr6
son/3oBFT2U9kNBhxPixBWQrpTlNJ9ZmKgyNkIzDLQew2BXdqV8vLhVwFOH8
mSuTi2j/2HN6hzwvjCPm4FGL91qSVThkKS5rl1p5pbhDVtXVEXxAA1IT2Abl
kkL2/afK1prjd5u/0PhGvj/4Q4nU9ucr2QFSTa2QkFqErVEYUv0+eI1jZybz
3jpp+pE34Hw53YNApjxMHNJdk+1CtPBQ01PtIkfISpxPq1TRz4FOLR9Npqkt
4DCWXrauSoNJHOrZGtnl7zGyP41AihijAszNPtMkziRkXos4/MWYz2YZQkdm
0xCGCP1RakIhTocC9BKSt7BP722UIikl7Bm2qOeIpNIlxJYDERmzkLDPVHEd
r7b+fEPREcv10d2E6vYR6rGBtB5oCYRq24Lr/5g+GT0HZ4sCi3mpHQ+VSIa+
X/Mt0UP29mTNSMTe23ZjHxO//ME9MghQgsyQdHrwijDm6htRfZHo2GO2szXy
96lhs5ytO5iRzpnQCJxU0gvNnwL0wogC8bhzssjIcGqyA28Sn7Y30dRFWHFX
LNDuQdQcsKjJDAIFntU11958xPkWN9N5O8T6+78pEwidUvFIqKBthbcVBgOQ
cdFXiVwKK4VmeqiW1LVdCJz6fFnBVN8ND2fteDmkHPbYkVUQvvk+pjdkPRlz
nggP8B45evV1hK+ymVi8OyVDEtSbD558Q+Flf3tMJO6sDbJW7t4tO2TQ3kjB
e9C8HbKuR6Y4TJhO3TqmtMpKNeeL9ZdRS0bUYd72Prqd0gxSHjK2sPqf4Bxm
hZPqJ+VVYeYzjRKSdLLzAdijna5VaLtr7NcMIOTn2sDrdutMadX+mWfoLWvE
fvXLKvc44U0Exmqrm9r/Kni/pnPYMTgmytJeXsHfWU5uslab94hDx+yqhGuY
EHES7Jsbt6L+bPmgyF4mLDyzgOugS60vH0nnFiPcFuYPunLKJ2c/bvbJU6x2
RJCUx4sU7uVQCTwGM66Xz0I5QeNgIWSOLsQvBaX0lgCaCYVnI5XTGu5CrekU
e6PHcSCt/gKdSsox2RKRAhJNA5+Ujtwu7qJ9igsY25JSQeYYUSxkXogRlpsB
qgT2M9cTelxyr0Xbk5PAYvU41dzu7q1Id80CtifBZWG5vKslm/lJnASetYQC
pREziTtZMwuyaGhkKPQhKXyukU09ta1eEKAcO/5gO0539HyDMI8W4albMPA3
qAuwnyDWAVPr5+3HTjpsjpkevQ9GOG5grWFaRK6rvSdLl0Hn0v/HSIijpMIN
VnlNDc99Z/WO2O8sOQQ71tcsF82gZrOV4y93ytZaHZ+JhD2eH78sV01nNE44
t6Gl2Hc/HDfE9lhAq1+ryBnOtDd6pgfi7UOYwMpuha3LFW4jPtBozIZV+/8x
LRBdFemKeGa9p34UYpekg7MMInIB9e+GupOP1d7jPIRs+41N5BcJ4ZrduZyv
14f9YPVTdO2TO7AO2UJEGt/3xCPDI7kCbSaYoNPzMZ9+M27nLbtw6HfLffTR
hBr+RVsKEFk6rvXw8uf3V/7HkGHFcjzpuA+pTn7xQd12U3wEZ3qFpOz/uHxv
/xSfyZLOrkKNy9t2IdriTpFr+8IYklaxzG0h3sNnvNtojeQP08LJLJPJsamk
JBPVk5yIu9NUw/A+7ajwkjMEoP+d1+D5Z98eVn+iR6rTKcUtOcM+j/ae3/SS
2pIMKvql+cAGDmERsgWfQ1PYFZLCyermUma5pGR7loUF5fxlLDZeexlvcwpz
mcw79mQwYmwqsmxVa1LqnNgB+2yN0KnI/JFx0SFEJG7znkgc7lIzuA26C7Oe
9EiYFwfrITZVGDkO9qSanr8UetY32G3OwEAFLstXLAGGpCl5DMncdXl5i2fO
T+IWiMZF5wWDaqEsDmzGsLzoOSOOoyBhS+DjW2zOGIbFC8ugQjaAtA/hIKba
v5mQc2XvH5UQWIUSQTa+d3TX+RNUyWme3XV/0YDB9jOeu6pPVQCJc1uiuU6A
yRFm7mFphXIDTawq4re/bhIj0TrX83EyUkiGev4zN+i2EP+C3EWuA11zcWcO
2CPHTHqh+2deW6T8BGZvaYHz3Sj2A1cYeBbV7P595FYunZn10U5MOuheb3FP
4R3rtkB/nC0QpDasCESTzos4KotFaOx8Uh7bMzO0fikuJuf6GNZGTezKDiR+
58eHs21ngckk5PZf+fDAVSpt6/v60Fd2y5NdhaT8jg/aiwBP7EcU0VnWhiuX
6hMbcXNuq/9dyNmioLcGALOpNCTffawjR40b/1L+PsRZ81k6eGs/RIbJXDAE
92euD+YClGbiXVbzMSqTJkMvdhtYcB6vR0HbP9B1b9EEF4F95SwRnY9oJ20S
bQqHN6DRgrLGvJlQJLGWerVIafCQN0DCQkg6LiEPhxcS/ca7ziFQ4csyBahV
NDG5lYxEbY0LdGu+d4hyoMdRcmn8g8r6oucqCsl1pHF8yz/hbHbNTOCbxa3R
Ib4Xfn76cuiKp5KeVBgkEikSHSZ/6pqp1b41Cx69p9gjsq2hLMK/gg5x/Qp+
CJmnFJgI2AxV8FX4QJ2fc/xVIBaYMvrV1cj6saJRkah8safnRWpm/R+bJe3y
K0kVBGRKisbffEmnB63HNfS/j3SA7x9Bwzf5EWD2cV7Y238Yy+xlXKJ8V7lP
T9W93KvsAHo+ynbcTLkT8H85Rnbatrx3Qpok0t9RPxo1AWFFZlyvmnwO179V
8G+HWAV0egP4/V6Fo78bk2XokM8bN7j8hyXdJOoN3b60UMThmJoCHhNYIm+H
LtrboX3KmdewyM9kApMTpdNewGw/M31fXiGg+x0A+qM3INLPCbdGJ8d2jHJx
Co8zlrjY6MEqXhFR1UHxxNLm64Ne0XV03jAv0LuHNdakwYxtXmUGcrixPZEA
Zl+ORRITi3tV4hKnxNWmspCcNjxPZiLTnGxFeeWRVwoWHILMXv0zdWLOk5zr
WbMQgadV2Q5X+XY3Scx1+LhwMy+jW+RkRzZNa1EIOuN9OTk680C9yqrLtHuW
iPbi4kwTW8uVa5wJJA6u1Xxbn1RpIv+vY18YfJ+hoqXjb+4UofYXKjF9iucx
k4GEmYo6wXXsStfYrEetC+M4cGw/dftI1q0ooIIxP+Ebu+uCsqDuHTVZpNwr
FakxeARdnMmp+628x9T9H8+QFojwSsHhU9iSLnIVV+iWut0+IBs0L7AZK6g2
7pTd2ggSrKoKUVs46WZdWBNfuGrJ82Bmw7JXwDkjJqwk2jr9vIKa8koFXhJI
vKSA5BpJrqN7SJ8Gzl9KS2ujpoFV/zVbk+2aXJ9/7VmZQ1vKvspERKuBm9BR
/7HshGAXFVYVIMZH6R9iSDQVQkuidspbbWYdkB7NYigydnW8BLN3rXwD2XW1
AdgV6Bs1iADgGiTsi6312ZBoLwbB6baPQfcVoUsBgQbg4F57FpFToT2kpQmk
DgqrewkqTrxgSbnb9nrFabGggStCdEABN7B0Ep57OAVTcjb3dJuQKa2U1COT
K2tU0ICMXtDVmYTS9tRFlTg9zjDrdokR9+/XqawMKIlrOjeAZ1ZfhTDib8Y1
Tm8hMS0ZISaNqs1ldLavQqy5JV+vTP5atU0DXKrqy4jqyLWpWmAiodEC4fSZ
6zadXK+qse7UvUTjIPT/ZdCJlJwGSkVbdLPRWPvww/87KaPqh/ho7bz0NDrK
SLDmRFck/MgFFD5c+xiNnxyKTJlKlTN3SifHSegTRowo0FcI4HkZcZr4gqrj
06SIlBeOlxJg6BnUJnPjeXFUaXhUJBcjflMLL4VRXuOjkxc+UEpKrYBqlQOf
VkqgQY3ke9Q/mjns0qWe4YmBDxEmGrVQYiWe+zJwxf9obase0ALutmzxUZ7r
/K0XnZlANYScYPk3vGyHkAieIFNankXYsAxkrC/DdMiqj/67JjRViZ3Y/r1u
uqROOeKPjPxnrK2UjuUJh4vHVEfJh4NL5fgb7aUb2Xzt+qHcajGm5YqGyzI+
s7OqsuxbFH2riFg3T1+iqTs7g1WhyjMwOBXgrpHs5IzurZixdsVqH5fHDliG
P6v3WJ5A4k2hBgFyQfNX3dALEmCdiwOj/tUHSAoRIa5zwg7GiN4y/FlgY3li
cZuG2gl7pYLBm4GRbOW0fmRX7wUhwNrqQpq0scnYXe0j9paDMnFcZzJzTEiO
RcjdJB0sXm8twAuk2FLg1Yeh+UqHjyPcmdxwy+bA9L/95/k/TqIodlBz0HtC
/Al9UffdLJROlI5/+G2aUSI+IylqZA1MhuTD2SH43wFXuBuBknXmD0Pqi7m9
irDiLAUs5s057Pg/En4RqbBSPXimZwOI4WPKWMRjzUD2mCG9kld9n9MaKARi
YOoXVhyBVM1nGNRFhvjWx1HV050DqeMWkI9yyDkxI2azNPy9GY017XPnSC8G
yDs8uHDzxujY5JnTjySgtQND8L3MYVSgEzwx1Ldkp/QRKaFBo0P9MCZwRy+i
m53PCxSIiBXQJYYIJMELUqfcblSWlpdEpNXEhthEOnceOTmltXXFENFPmkyz
tICGzfXRkZZMNpLGxhimUXYl4v6/CMO+MV/yt8JNF1nQxLtdmhSPANr/06DU
9HwXCDm7l8wAHiItBTrsgl6l0JXap4MBVglKrsNxZSQOB8wBSrEy41SXY9jx
acCrg2URQbuGByxPAvBjX9tYACubyWDFwLO86GtUOvaniUCo5hIo6BqFqW4Y
+pgxESoy36HdBfsVHjTcn05P/VSsKCymLWsbS6QfdkqbxsasByDrlRyyr1zx
v3DqknMSIq5a53huq9XAhr1+L48zlBeK7epFBSIM8ArW4Y78SnZEhnC3cW5C
FJmQexv2/ivN4vih9ERHshOQzuz/OR5CoGWcpk/yv8VuheGdGUMdUJ0sOyEY
hAdamUCyjZCrvFMFW4FLS4q5vavBrRU16PRE9o3tltMNakf0t5wHkoMLHZSp
3pjFlIOwkD9mVlQbORRvAZJUnZ6YBW52xqqQL1WpC87HkRoY9u5yE5v/MRYs
6SejBYNGpef+xJq8+NHjmR/Ur0CelbHyvBGwxkjoUOLSqpCFG+iUTm4C8jEM
oC2AglVTakEEE82jYpceN1hUxg6rK5Ahv/ocoyi53NSMJewuzjnvog8XrI95
ueRxMBwgqcqB9gnjkI070G94qWCMmmiCbAgvR1OgSwj21an9pMk0UT8Ds85f
/PxxNd72DCi0haw+DO2SO2quIoEpM70RV+QCuqXbTkGQKZRoI1b+hFO7Ayel
+W083+Lxd7/QKCLEPz7UTqYKNPND7XvN4CC33lcWBLScGvirySCZPPzF25y9
c2rHK+HuCBdkbNEu7h5EhPnfFbXCmPB+4fVRnxGX5h2Q7Z+m731Bh2aAY60/
NnN68MvCOPUmQS9pPOIpJ6Y2VcGraTDXjw0DVPu8cMGIEXxwNZZHUnwTXi5f
qnHHuSYM+kvQDlALml0MoEOBevRrbK0oOXdGJgMmHaQNGTpfGStWLOYRX984
rn+gPxU79i5leyJMkkaR+IrLfJAmZkcniA8f9QM2ku+Das/GnzECNimVgnZY
k5GS/BJOn8b1LUC3jMwT4ikKk/gMyeOrven5G3rin+KA8moltW+GONgGLDOx
lZ3cZZk/O3BHortL4vkg/omiDCirvlLi44RoKI+mxWJMptYKJDuy1gOTG9jr
9pt3tRxv120Km+9J0uu1z3re2KuOF38KP64AftAsolqivfiTOcyZrUBBSK3/
niE+Up0oS4VgVF5xJJfTwLJS6m6vtaIYlE9rgS2x2wH9P3DXSxXKmFEIOHdB
VYkmbktStYna0Dy25JJONsVrdakZc4Amdz9N45lDirW70ZM9uvcbKeisEYsX
yFLWVjVQW/+DGvz8nzulb2tQc1LGQ29Lf9Q1XLsKR7mWZo1obz5OQ1ya4HDL
YFBG4uun+kg0O8wvY4aq2KleYlIPjPXV9MT1WcRVqfDQXcu/OQile1Z761C6
gMIXXYYn+3UaUIsYUgvkQWY94Ux729P5LaHpM7RNLFibXuSAyIPwjpbsmOpR
EeotDhseGEMKygzeY0xbt+QcJPAFUQ5ggSAHO/JnYSGaj+My8Iwbf0ubOuC9
keihTnO1Fst+xrRP62oIQtntkXVLe88LJrP9OZ8EsuNEdBA0pMCxdFjO9IrU
C4ZZ02rgo6Lsaq3C9827Yx57h5LJ/qNqdK/zXg4OrdqC76Az50unxDWDJtpb
KnNTS5U2cfAIUUyFSt+qC2hoCAtz53djqa8Crn+/+bHf3qBC04MOnfm9XPz9
WMxGsAScgndBxWrAJ09lvVnEowiFxYGumIx1MbxCoxi2V7YJty7twuZNst96
4aIm9lwh69RnIRiDEbMbnxKeeh7f9Q+wIaUNwcmNa1+v5KDNXieLFdjeu3bJ
rmYBJpMykQCuLNATehYZUxrW1gEKCsqc0aCF64KeTMZ8agr9RcAQGNCrbWZ1
ewpSUSpYhJsX79M8q9b5AdDTG9XAoglD9VLEk+o7vNMnZOeIcDHe96P+g+29
DdZU5aYGrXzjzM03Yrkj2JSuSwiT9/2AlnUMNRAmS9qWRIyhyE9Bx4jxLDaf
WXbq4Ru6L19RY2XzV6r7XtNMQPEMqLj80geVv2084li6dzWm9F7xyF6TfAfX
QwyX4Td9d99EEZ1zxJqYbsySRdHOz1UQu86PV9+jLlRqS5dvUD/jY7/xxaXZ
cUB2fkt1a2SFgybuhpWd9uYL6j82qAWDF89xjsxlgKxMg0KGE/W5JsE+Ep+L
clv8H+W1Fmpwjqeif9R9/JvxLYHwTDzkmoeEkLt8HTY9EpMf8FV1wDH0TJB7
RMxF4gVO3pwcTCem3rEnKg8dz3jBP6x8jZTUZAZeDnpI0kp9dyCKqrLe8CsA
k1A7i00vjYxiN/3jAq2U4BWnEftN8foAKN3icv55dQI6Gq8koq6rOFXDzkdP
4hIUh/B/EzFowwPtNDyzDL3eUVWBQsjBeSjhvKopxkcM0HPOraLU9ehV2fOj
lWzUAnAmucL8ejxv+8gQKr9EynMQQ1+/cZfXT8Bz5UJJvC+vh5rkaeraHFe/
AtXJ7Edva2Xn+7tLvQzCo5qiqe6A04XCnBcYdA3h54nU0QIOtkaihF4b64aR
klAmF8rGFOENpJevtPpIkH0k+SX81k2pcN3wRNRcILhV4NloSL6Rk7vSoLjr
5XeRUuscb7xjq9UaPjuQ6d1qrsCtyYZci6xGTOskgf56bsHy1QIKs5wS1YVn
c2n6iSRVQvD4RNoBYa/n34k511sX64dW9wPEMfI9af2CoP2qybM9PG02SqAL
cDFVVcgrh5Zp/uZyFte6C8ZyKcCm4UgW5Jas8dipupcs166xzt+r7dAaSqiz
4kNPhNEDQ6wTSIey1oUGPTGscBCA1NG7db+vlHajAd1rm1ij0tf0N6It7Ei2
2CdFcYVZ0TxUgIYfmzaR0BfJ6UUXvwBjDWUJjJ9cr3dNljKlJb9j01DY66TV
jUJgOp7vkAutt7HMv2ukhEK44G09/QjsAfPBQNO88SPEa0I8sULFDatAgJEK
ycJI2z9ZTXVhKnewtSOML6T5jCTRfdbB19qlpqQu8U0mIO37dh/Kwt2WBZ7k
CTwtPWXiNuGr5GsrvqEEpa0p2NA+ReCXvjn5fEGrvAVFMZnc9OZnrnwvldGc
tr4NT1BtmU22xzv9bh+pmtePP2NxGyYBqwrPFOLWOVndQq9woD1S+oSpGzF+
WFQQjuY7D/8qFKzmXXgPFvBDb4SNRy5YeWYyfSMWj7jsZgNGEx+toP2yeTND
4QD0W5q+zvdg4+XaTLlwFAEb5+FTYM8Q0M06A2J/wLqBgNJBi5Qfh4Ckgpf6
MVOJGxUW84oe+MJP6X4YjcjtlTJZkVn2kz+E5wzrfiux6kqdWf8Q/L9O8WMp
odaZArM5jfp2eMH7MHIjglyW4Qg3mFEhT5BQe8e3P4XpKTnu4WljwAZ2xBWK
w/lebCGvDcu6d5VxglP/ySQIYIkBde+OROzUt6Ylhj/i9EYJzethi4KUww1m
RWn2ufDblYLXfLz6IgSL4vGcbph42iD6qx+M+4z/sNsrOiVVE7PiLgcnPvXA
T7iaXd1ELcc4CtOX8IP5Vj4vhG8OrGudTEK1uij4Zb5pfE+yerVBohe7NNMC
l6RFkOeICygdWKlo5c2A2Qo0n/y5riqhfd/fEUaw4iEEdBIyZx/MNFm9fWKr
rq1+FaKId8fa7K7SQAXg4jJ1qRHw9FEXl2cHEnMCsWT+c1v5hy5M/HeZx/0+
X+YjVWftSxeflRYX0dCrL617tbDus4URc2x2VcMvS8w34Q432B11K4UaJl4b
LUoOPpK14caZODpYX+pzqN4R9e4HR3flJlbuXL7/3QWReoueVEjJwKRa84aT
Jigfh8BfApTMmJJL3N9KJxZTCeqF3rNLLvGMxfVEN5H7o53lOobq+/XqIxpx
EemDgjEdI0w3MASyWAnpJprgrtdTrDaIpp3LzhhhzPWqTuzobARGVr4k7tEr
6vhS8hN9sCdjjUUiXjHNSoWwqsYn/GX9oCGExDY2kJQ4S3dVWo7IEEykj3sl
k/MLHH/xyCKsL6BdpUYH3akxKAGzF+ez5PTwH6lIz/yjnxglN9r9Rgcw3D44
UslApj92LTdeuuQZigQPRy9M6Ndio8UxjvqmUC9SVvFk0xik4z5D2vSmv+OJ
S+A5VU6ohGB8dpS6MuRNh6W2S77jSC1IYRgs9pZzFmr3dAz22Vn6H4Tib7b1
h1PfVjPciqQuvzcvTd/uVtDOxHI/OIKYRQoJV2XORM/4W8uXBk9WO/RHSzjO
aNQaS475iXFtyMI0BH+/9a7vx/NMz5GCqzrvSjfI2wyDRGFJmJAjih2avl7Q
wnWLriCvRJdMbtYsZM6buaKcSx8ENykTRpe6H5U+5FJ1jqKLcujrXNzEIifp
bBeunZLabhNQJtTCYpvQ33yEw3HbPyAgWye6gzdO7GUwN6IIAsucyNuKC5/p
A1197bM1lyqD316wj9q2qK+j4d8Og4gK5UKxzy42FT+5ahtR1K/FpGAW0tKG
MDUL2Un85fYSE9xHGeDKvKXamrVxHJMcI5Y0qzEqzBjLn/tsBCgJ3Z9Aronk
farJuSTixQwGkGv+f2uHUXuDov+Yd6DTEDLGlrd42Qc3ggL2MsULW98Yqy65
ttx2xuhB5xxKHzsSJYTaRGlq+KV0YoEsAMXYY2b2g/DgoxSM+iV1mG4hddZF
XzCAC8TO0rRpicPfOPyR67DalowqLFk6LyMXFXTjU/oS5RzpZgukXINQVSai
DIVSSjSOZUMzr38wajtgZ1Hph3vRaVCoN9bli4e3kSiO64K/9b51NBInok0u
h5i6hbrvlI8o0OpN58D/uIHhtJFjsFp0aU+nxoQ6XeT3B8kugeQ8QzoGzBuC
bqrTDMwXtsU3WuVFpkBd03yymWXM5bgZVhGJUJznt1FGKx88unu+Vj3kafsl
O/b+2y4Ygl80CkyMUeg9+3j1WIauqDjXOtpRD7uAMGNqFCWHy5c4TSA6GyBC
f53I8LkIJaWlk7P8ML83nSXWs9kvfwzsPvXwlg/XuuU3zwGnpKSocWwcag/m
10PhsVUNUnsBfyrQ3parCZl5AiMdfaZkHPTI5sRZ0xRGJm+YnorSQtjPXOVA
jVzH/PgN5Fg5oFoOB+2ztnxtXUPckbqIwP+AokQ3cvxg9dQKEjj+G9/Ybo2I
453J3TJhU/Mbq2AEw0IwhGYnlF1HjmciKN0WK08oGcCjcDYIZl+sWyVmmLx1
tP5hgdCkSTlQSTYiXd67lrwa2eHAISOfSig98zqOPQZyZcwCqoI2rVNA1NZ7
sOZ5cAvOTAUmXaKSh2Wb/9XUZ/j4grthOv0+sHB1NNUVAZdQJa9YhprD5UfD
cnIOd+jqWOg91oKiQmBsPgCsOYTzBiIX/LCrF2traXowEwgyjATDoWtaIdGb
/jsF2cPt7q4Ut9MpYO6w4BxM5K/lqgAC+taL2AuVsM9O+vvPR29gRb4KKq14
8SpyyraXqsFo8634+l3J7XN5kCyPs4XIbW+bIkxxnAd6mDwCRZ4uBgKDeVn0
okntcrxiLbmwpPIPFtWXplI8SFsgREvsiuCauZET4uE3FdJKEQOVWxK8sRsK
nitmtEIXwmhCSajcEXKkCpLQVpQS/lXcGzt5GqIHc81N1nA1Ps7nkzripjgO
dOi7Jm9qPc6kSgPgtZMA7xweDdpJP1J0tXyTPvxgZmxj1sdhmZrQj6NwSEuM
d77SpQQ9QmVkhf78VB5rNXnhXZQsWpwbEzSIAXSjN7klQlXHFLl4KhNgEstg
tOAc/78hujnKlLUN+KKMtBjfHsKiixA3cB4F4eDxLv/maiBFyzCXA/sSGIfb
13SGtQeis7qlu2n1H+SjN11sIc28fxEISgTpyqF22R1DJCU/vn7ic+0RXlNB
HDzx9AnkGQxk7KTJq/JTs6F3ao7FvPp8yksjvNkNTEosKFuIEgvIY/liU68D
7gGXlGNAYold9aMR/0Vy7b56EHdbqr4R/7YhVAj5JVNxQPx8dS9Te2HjKTta
Q3n4PmfoU6/CnGn5dTP03LH99lryM9dg2Q4UgejkdE4lETe6GUe3NaehzdBM
PHhdDd408zUC/HRWzr0+J1paADaxpF2zKv8/sYHQOOC9pVek2ERWbGAsn23Z
2OgOlVrB7sCLTwZJlejm9n+B45jUg7JmS1TxwrDqAjeuGyYmUFMfzgvp2aAX
qhnAKSHz21FkWI0u9lHq0eR3IVDnCTbxDgZOKXxF0XCjbu0aNCa3cq2koldA
2mmGg5Lq9LGN9rSMapJQXjIceH80gFDCAtQKDAbgrC5XqWdHpJ891oKgzoqk
YfJsz0wEK3YKFPfxjSxzSO1WsL8uc+wxo2+Yiekl7up8tGiSfa2w4RfJNNjA
jFqAai3yAMELKT3293Ut5XS+u8Ax6jsjz4jLVJDGpS4UTImoCNIluz00lqJr
zXtTD+ujK0/gGXjRa78tODJBhJpf5W1n5hVrqj3YEba2wtN7uTS0RzSC/g+w
k0Msz+RwVmeQwsLNZDnQyp3e2lg3YI8AHX37lDgmJibnonPvgwAXV37Smw0D
a3uBMA4dGN6zLxj+kRIksbgLg85S8BbD94+4jEBRSsmWlPVvXkbsvSp9T5EL
gHhZIxd/xX9OahSNNGPDJ4GC/0LmOiqClXVs1sgzvAj45U3TyB7DrOO4Cqfi
npXOKP9u0+28JZr7bEnsYLzjPg5ahpP+Uk+iMs33Zr3JR+zH3i4M3Vl5OSao
BK/RMmraUQrjJl71uYhi3AwVROplZfN2CAXuboklwu/5xC70quaqspZdV0lw
0nXaZuO4LvVJrFYDWi2ZWAI/zkbFmY+y9zDP6zp2gv7EVcvN6NLyveI8xGJ5
dvKRJkxFBnNM4aXXUDRqLMgrPEHn8o7AlfZ8OPjqXf75tyFhycSU9x83UpfP
0IpXJU2CajoJ3g6C4D9+BmcYEQHIj0vHyEPetZUBx73mWGllh21EDpplayN/
tvUbHSa9gNsS9VrQ7Wg2t4w6A53AP15en4f35y8FS2SYm3q6DWnCKK10MQi6
FDcjISXqpowN7n9pgwJV82zAuUKMgDO9rKi2C3G3YTS7oCDbZWO9WDYarKHB
ttxR+qQord2PXeVK+tJmbYhpNefXSGwV6geyWYopwu4haF1B8DE0l5hrlXCh
2r3p3gAXwBv5BTQtVh9EkySI/bWO0eE3bvf7h5j27U/AY504JVayUtlYezZK
PaKsKZ9pTEIcwSIURTU9xPb0d8oukF8X6NMGxBntEYnSdUiTixEqZ8dtDhbj
7OEjreHCnKedJ2bN2u8c7yoFb0GWRR5IBFYCeSToRYnQQye+pIa38fc9dQ6G
YSe0EV8JtnbU9HTdqSM1k36k9VC8trr1rgj4Dm0eXbnAcDt/JLTsci6nHhVB
GeO9y9q1jFc7tcO3Dbrqrwt6FkGh4Q4G9RQrUMfELLNCinzjYOOlLZfyR8da
g+yhHLrMkMvCqYqruDs+JMxQkAV8oUeptT6iX9oql3eJAi+6xqLFFcoqbAT2
MPLkk0GGV0nxS+T6izklIfvllmpiDu6Np3eXoM4UrpwluKwHJ0LHWly3qeRx
6cxhIWzhZCwdhmcetAOl3KbY8Xd+3LAd1iD0RB8LKsJLD3b27w9b9xyrC3Zu
TErhDzUh6Ohf5EBgMpO0/hdIQyRi6dv0OitlbuvxIb0F1w86116np9f/rNJa
+gYJa59iii4+QNJUfGforHzTNyamaEDP2wFeexbDa0SsFC9TCOn+u3124yZ7
+Ydi5M7kvJZG+TfdlZ5uOVZUKymehBGqml0V+Z5nHEHLEag90rUUyNNGbBOU
Qq2DyAzYnZhSLbv7877MekQuSGj/2LcdwzRSugd7cWOAMAy39o6DjFnhUd7C
7RFlhrIKfLaVeCNqdLP7WRRCd3GGaTf3kyIN7Clhb8RcVpDSCseyMqIJsk4Q
l8JINL7aSr9rmqR8TmIu1V1VuDoLJQIMNskW1GXry9tyACk3qyAj5VH6d6Yc
233tTrAMqDVqMon/gF5DjMOd/4eGSsgYVMVHOeHyLO8FuwgLSCwpTQ9KqSBi
1FMCGu2iqE4Bq0FcZW1sREc0KqE87SGfkfB58TRoP9PwFSLsnJ1EVjSOw+k7
oMnbVoXzD/fKlvY11Rqu4Mglit39tCj1h2AsHYWptj9y7bLqxDx8dAmwnBpY
mNbZb2wCANLLQhgoSdAcsttjbkwx81s7TFQFGEDSpNJbJ4SJauOtBctp6RmK
0ihZpaA0XX2M3RBtQ/qgp2TWJUdyijP3OLouC2LXizYEIvUv0fwVE3djvjTI
IalpmVOUvQi3qQ6SMwoyvFT5IfI6Tj9/kN+eUymj1ep6OLqUbERoV2ycfC9l
BldAAZi1AewouLQieZZHDOJZ80FMFZksRMsOMRrR5cYGybvGUcTn4M0E05x7
TsvWcwW+RFbNT+I2HmVCmqKIAv1hBedHl2wpQd9t57iajqjW9VUjqWXjhBRD
N442BdzekkxlWthglT8DVB35CxSnMeD6Q4M1IOwjiOUQIQKrc7DROs6a8E8W
dkgcRmOEEaC+ElSOvNvlvglPlNLSFzwl1ATlQpxFOZV2cV+lCTQa87IUgp/F
OcWvyGfJ7VtGtKxDDV7HDNZ5jywktMFEZcb77SXJwLKjL8TMOLzqWcMt5uN4
VrWlRH4YVFuLa2wPkRvl77gsMVLgNamtIOmKXcUmaWPaIL/PpEX4hf7fYZfd
jJsCnej5W3ukiL/6ZDU35XOmN0OIrLI8wxFBlRYlIyM87B7wbDrKzpqQvk1g
DCtJthRF1WgT6fNxDMgUtCAfwTAMn3RO3Mmh4RqiQ2eIqr6jjwsxBYKVIIBt
xYNtSjw28QkiH6o2aMDtxKk+VkeJEI89+LQuknZJ8x7pVCuGy8mXJ7AUE2+4
fVdiCkrYLxJfiSBNCUxEEJRs51LJJsSWtk5hpesBY2bRJ6oIIwScIa3qPLW0
QfaTGTSlb4kkOfixpt1/VX3I1+vP7vPXGTq38u1mn8tgq+9Qbx7NvwuuySKQ
1ktDs7tarorILY5eCS1LzTjx/9QYon/hMzscFuaM7249DA4x3OIpnI2jxtgE
6tPLSeH/QUkKjhs9vvacngF/SNWF4syVUanx5+z0H2qfuy23hycZswxgDwXf
NFKJ0fhAc3pItaXWBN9jeplBaQcCdhvKNvhxCpOW6LLIk/HjcZS5edpBBfiL
P7+ojHRig+u/yto4mBf1YC9rLinuzUXCv8XgYMqm8u6JXCXQ30Jj/Hj0fD1p
UJnPQ1nIMJcuLJwl3fOAfMKHzCgykbl+UAyc2q76BUTKg+KBkGuQ4OC0a+ww
SlePHFji6hguqwPsihcs6p0qaIpcV/rlicDoDmscRHX/Es8v7v94AYbdc10U
bxHxOoVHDD8ftMnavQyRMglL6FHzFYRVhTvddVMH0vN7TQr7l0UsQ+GOEJ1X
5JmId4a9vZ0Cj0vwNYOXGlAAaQs7DMsdhmmA1wg83zZvxWG5pRzbe3CV4C0C
5nOGjZA6c/Jo+f7Hck5d0u8R8RvQOV8bn/uePQQiL7x8dCVYG73NQ4GByCm1
QGNlrwk2XzSoEEhYxij2vV2r6Jp9++auxh0aTBaoPW7gDQu4PeAB7xlsYAT3
/V1CHL9Qgf3pNY58l1E1bOcGlYOocc+Jy4jGV98ZN37nZ5Eto1YrZgVaTwzw
gowKkgKA9cTVdUYKGWY3hIwKu+PXjMK9AuZgjCJZpy/8ulor21fgl0UulYKp
XpsKxfDxVCNUd/DjaTOcDlnYtShPK19cgpYFBCAutU4cZDBBXc0ZADaUJHsb
bMekP+57qGJwe4XADUxo32FpnTnTAgWb6VSmzHn7OV63vCuw2+ZBBjwImjnS
3hjpUOAxn5Uxd7ZFJeMM1D2MYTMsQ1dujFpe8uWCLNKPseHu96O01w1Gf53N
IjGMb7wlmcy3RwiwpODX/KiImSRsXa0cXgRdrnkovYo3+5jALBot06pCHfc7
Q0idWC8tsZCczRqzX9HSjop+KdJsQBlnMkBqcuTt2WnRU7pIwDj9TTJJZSuo
FERc2SfJxaVBJGtYPpT2G/hzFZuhmVxVqRP28+WmT4o8ZgPyxVWr39pZsPyO
06Ru3apnhFsOMvRHUNdhivJDvqjLhFLaRHfLzfqR87kRbD8WssvOGBh122it
KQ9uXAfKuyp7x/LPhwZfZ5zVj7f21a+JgbwLQ4PV6U5/HLZCn3PooxPbweMt
4TJbuoECOj1krIU/ym1+rZDDIx3OiNU4C6szrDeELy+xoB7cgCmYtb1Io0um
xKIzhA3Xc6bHR5mJDyZyeKXTAAVN5eJnKP44XSPDJANkeOPToEWIXAJvu6Nc
ZaTCmic1haYeVl5sDIBtcIlrFnyjndRA2yzoXRpgu9smxofAFez9RqvHr74/
/3ez+phmjV0AIG242nUzSEJ/pZ4NVFWmAMKX9G67fZqkKFmd4Fo/0HB5G4Mr
3Qxjp6kcwZZIGTcimatsWhXGasPg6DepndV0FRM1XmVPTxrMuAGOY+R9lMEV
auT/B9EIpr/eBUonGV+i5+yP54WwWBer0TEslmQu1K3wK6Qep22dO0z1Qq33
tafIYFMBSy8ZCX9OdXRNgTHuk+BqcG9/fUnmuPp8vef2z49O8HXjDsIMyOIT
JAq9afIk2UlYeuyDMdGWM1Buc1HEcld60WtDnCfq3RdkjZ//7tLkDci8XaG7
zCH9wGLtYy3sW0JvdnMSbN1pgGsLYfVsqVRpsFG+PheHyXUPz93wnXvfg7AO
COCuIMMGwqcUFaDnJE5jzy4de0MY8ws/Fd5TxVJfZnNXeTvotMOr4zLxvur6
OwnLL9BtGuosGSqKK1oK3ObLhhoHqIVnv4asjs4Pg4yoFudwdcnAB+i3KBqo
Mzy9wswCm9fmV14eOmvm3sVOVGsYYpx1KD9BoNmdmuwm5ureR/rQsJDaw0bE
PaLM9PWfjv2ccKqfw+2gw/Gx5MvUR5vYTvlhr1gjwHxMUbixNATmcgrGT9Fj
EqQksw6SpaA73gFkdr2j8PGfsVCtXI6B6p4q8UQIdO3m5Aj1q54MeNiVsY+K
1F5Hdc1rTFWF91lGN0XGdwVunbQxiGBgBHQqFZJ7DX1rC7sY+pBbMWwdqGlq
fpl/Hb1fLZuO823Hey5qIHjPon8skJYxoIydnojxof5beAA0UVpWWF5dUhus
FMV8EYxGZ7b6ql4pjogfjaRXeInumbiQtA1Jcc0xT6gbxe8cllVLDotBmWli
WKY0WTHf03FMbnd1yDC1+aPTO3c7Oxsvdh0p5fHtMUAkBcwJf+QTSvcHYU/E
s1Y2s5r+fMMrsr7+Q5ZAuKgtoh/X1r0BG9DUmRxiIQo76rLZBs7XDIGWmp0H
GDkJAE7p+MZIAf/zz19FnuRVtwsnyg16AAWAKx1+cUudPPjOPtpPU0M1v6vR
CW3r2lahC7hKufZzxsrJwtCi/+SoNaCxrH9I+9f8uTbFxPoiM2f33ImpEpg0
uRZmVk/0p5tn9cebRq0JQ6xcwaKXDBnAyd4Cew0sf5tqtdB4zd7DlDw+zLaD
O6P20unIQCk1A/W701ErqiKwBXMK6EX5E+GBz6Stp/YmBW+HbwL1qIZEvlwH
NVD8IQiV62jCdeZC89ZRZDNp4z7Tor1FVbu7LU4RYtiBsOsnvmBEI8JpEGXt
4kqh1F55DnMaraEyY2zV1v87xBetKMcEA+/HTPQLqJCFvLMFUfoE0+hAuDe7
1n7xTPYK0GtFszU0eb04Q1K9qstYW8lmtZiKFm+5tOdpRIA4Y2blx4TSMSuO
aYd+t/ChA05VffK1H8JmHU2spuHvxZ+KbDmIVJL+3iVI+KDyBRBgfovcyr1P
MNSqsSBbXkdExpbkPDpIhBYRAMAH9OogiLuzRPdvmrpGdOnMl5cEZeeTOYaO
D3JzKkTuIF2njW6skY0i9HsLMVv5mbzSDo+bWUrpk+qEq2waNdHueqhqARNg
h6RiaLW48W6fnFdF2K+64JAKXrbbdG6+zrbc7b+IqjAlVwZiyHv+P3vKbGFs
0/Gzd2g9e70EqyfsXc9shfKgwauWz7HCt+QFKjluVF57jVythVqtd5MkqfaZ
t554fp8vvs35E1sAKXGCCq8FF2/0uE6jH83mdehKmocXwkb1I5PZZYOVAm03
qscjTGpAAj2gMg3sODAWDSRn3ant+ej2rUFpv3j3ih0ZPRdTNE9YZo/6p3H9
/fBm9irXpvtoNAukNuFjqpFRk3Yv8gemA16MY89LsKbyZBZKEal9gdKdcFal
H83BtSrsYZrvj/v8yrEM3xj6E/6OFjuPY/LTqnfI4Vad5NyQeITpJBC5YnK2
0FW+09EilivnXKifAmiaptFwtblRG6Owq36f90QjYYY54JRf2CXYVQcfQohq
UPD7ELcULIb13ZJ0fcphe/nYa6vQTzJXqIAFS4emJI3ALId5p8+iu80DpUv7
p6+v3ubhf68pRwW8Zp9FaNp778l0TG8Tqz96hjMGPWlZUvdyzB5sBxoBYKxg
Gfr7PcEd2ubD4d2YY64hRs8Nh2OAAYHhkaiuLgefCytcQ0MrVeXrTxo5Fb/9
jN5t+1/gjUnVSe1xrFdQVSlzX6Hr8zlhKaYZFjdleUe0F5IhU809gsalE2Z5
kWQ9bz2BFrJ6WhLcCsA308fJ7KWLX2SuairxT9ySbliBZOdcmO66Z8LROqpy
67tSPv3I8RdbuuoKJL+vKN8hSQ5sg/tVBXwnp7cJ13MtAySWm/xb8KveZJiX
0PqFOtVDXBqFZ6R1FZVyRF8k8ER9XT1K04A0f/dqxnOfeBsIg6/OuH2IRRGS
bynEXctWUQit1FRN88tBnZ2us41+N/8krUQEtXeK7xqzAr8g9dY0+dLGj1/X
/765CDC+AUc8R4vTsIZ1ImX+lxQdMkDBm7iJFX+oMbCecGkO2TwjgtkOwIRc
N+oq8kf1DuyCiAcOCjziL/RWqKap1hRYAoKW3As0O6BMaVHIsK9snhABZFXD
i22oTp+9ZsxWiMLTwu6xRoSm72RhdCGpOV7/CStcjy4zi0bXbP7MSBPJ3uT4
7ESTTZ/42tOU4mbUXIP31ywAhxulIbg7Z3KWvk/UlJcigN1Pt485VRUeFU/i
22Ym40ox5rNO5HqxCn6gz5JKkWMsx8YmZE5eJElBPR2Y4Mrg0KDgQGyvBF80
aJLVKalGecaMPeypuIr8Xqmx7KQHmAWaTeUR2//soVXjNfqz61w9s950h6HJ
k5O/yUax1UtiSMnqjmroeWWYh+ITQPtPrbfg2+yfU/1JDBUwMz4KzJYEIzwI
6t7V4OYynnV3rF9oeOfsAPNjO3sh5bDUgsx4G2oSy0qPi30re3CiGsELAClW
t5cAy1Op8O3uH0h+pESZu8T91Kxpuq5JNfHBB7n4kv7n5k5ZPBwJ6SwfBIzw
8IFPK2po/AdCwpN7fNQbjUqLJ0RCNm5KxFp/YV65kI24lvUNwNG0h2nYu5Zp
YEmblE40e24rJPZjAL/QfxWEGh5W7qJVHrGFdNOb4UAlHnEWeoavvNEGEmQZ
91DEObMu+5Wi5Tprz70Sj2BPJB1McGiPJ+FDfGqNMcGX0yM4ICxevIpfN1St
mBRkhoFnfZS0jL5GpzUNDwjCCTn7u6f1QHqRYGCr+hVBvszl5b7p0lhwagR1
XAst2BdwfGNtU0sOHO1rUAuuBKF1h1WU5HSoClAvWh6YOJBoY3GuJ8nHgNUW
nootyXINr2P41z7QKa6y6Nqb/fg3qlFN/3Lbmx+DFUO72yV92oO18fbyN9vp
tWmnNLUn3G9Hih9XG5syQaIcwnEEmdJeo/QuCaIeMbQCT/V5mRTUFCqgj3y3
rv1hQI3WdF5sT+/nqFcgMSgMUEAhVbwS+FIClEj9mGrxRr/64tWNdKR1t57U
w9MEUdfCwxdhRo6WP/XaFMCT0NZBhFGezuXxe7/9U5/H26mj15Op6Ev21YuI
/kbhQm2YVOqtEjL2eoBCzMUmwOrEKLhnkYX4u1n83FuRDnYDfHAhlUD5ORUr
l00vkL9ppVR0XBIEMbQbarXzyg66JO9RJDbq7TV1Fswt3pdBu2XNB6A5CngG
yr9OY5/FfSxJoN9+/dMczQ1XfuUQRGinxM6+umk/c4NFpD39iN7kfEkkptmM
bZ7V22nfeWisH4R+zKZ6ZqEuYg0cUHfM+S/SWS+bVqasN41g355faR0z932o
F58oYh1aTAsUifHJFyunTOm7CxV+Znf3M6VFu4ta09zffEPfX9+6He1S0OPe
erTlRPLOEQHq97J3JLyz5nQbefrdVITsYk311D/pE4fGkiUp948FDLdALiRO
St/PddtCvX92W2HBW5FZr2QcAN5IOB9AiIBxBxJY87C4kZCui8LjeYAW7w7d
jXm3ycEpIXQKtaAXwTRXdtu1QHtG+knqRYmbnpWIVGSH+Ez6n7bfeYv7ryyB
tDipv1PFpbDkA8LMZ/WQy1gQzzceeWGIgW2DWIoC0t/pgggATGyqdMx21F5b
SQOF+o+Ven6hTaLpYemBiLQnZ+ad2BSKU3tiBSCOGSg4WzWLsaNi6TNxZ3me
oYCdUcw04sgLTA8F/L+eU+A1HFXgqJXGZkd9GbdD0XTUZ2hC+cdi/7PXP06n
3ty45x3xcXTnSklAW6bh5RPnTUMiD4ElTbiOwdSLFMndp9H2qaUYHTcrT84y
EJWKbiRuWt1RdgYNbS4AoryjpzxnumKzsjUbSK4iW4XLUcZp2O7fu7WfMqj5
skNc1K6rWrPbsQ67+bQcinOx/+EfjKJUVzrHPz/92GWajPJ+abTVRhqF0lsY
Xh0SNsHISCioANnMCdKzX1TrBPbRVe1kKxJ8TPKtFdyHMHf7siKjUAEsNJKW
Z5PvCgHRQp1JVmUIT485aheJ259vzHlUGxmYcMk5xxTOetj90FgPnaGqsW/n
8iZ0Bo7qT4oPzzf+CERRQO6KgjtC4LPMWFzklXZeRZTjx73xdnI/TYlOw7k8
0RxCA3eWa4CULiTPQf70BmcgD7u/rt+ygCwYziD5sJ1bI24CEZvCUXqAt6ly
HjQoeJEWJBoEDxYJA0tjz0uVSzpNWULPkHAmoSRz+BZ9jKyHVHHhWeApe1mL
+PM6rtaLVjgCVKDGMTuGxY1QFGXp+j6vqvZVGjPkmGfDhfVMcUXFMcA24XCf
X2hLfbSZlHaP5FVRCCS3Y0wwRMUKGeZZXhn6QnkP8rB/OLIQKxE4VBdX152c
58YU5Fq0rdDG4UJrd7HhT/jK/ZE/yW4r0YnmnAvSDW1+YQ5xA/Szo0lr8dff
FaR9M+Vev47bORsJjVhDOPLSKSIHaX3tbfbH1lyE7apQqb+f5FiKC4T9oSh2
G3QFfE6IVhu3CqzZiqtCvfBcLiJR1q5ZIctzsGXfrYW6sEAyCdQLpmAS32j7
qbOhzlxiRp85DCVpqqpfGaGjjji9kjMIF3u+Ho+lHVEs8gCl0Ckl0oAe+DSZ
5QwnMYJO7waCQ61idvBNodA7kJKjk7rtjuhntFkIpvpZ0uAXZ+D0HsqbM4uQ
JrsCD7/mWj7puvSYhBCBv/nixXYuudMJ89SQjvTeSjGiG9AwUocgYW9Sp22E
sucBFVLAE45RR5CyiOBQLwpeasLfVzgGzLDxvzHhaGDKPm56OZr8GfIRu8S5
f7cE7bxf5DGj3B01e0wP+mT7JoMRbh7tqn1SaBD0tHiNUiNglaeTWdKjC6Lh
ri1e3emnH+gYSn8BVbyRr1n937mBb+AxbSpLsXK312jA8izu9H3M/y3LM/PI
rywkRQn9u6T5O1lHiTfT08euw9L9h5/HSAaDRZ8Eu3tS6p2Tqg6OVLu6kf0w
Y4wmKurUzf2PLJuwvnAix51vUCuWEXd7itW/GOXsFUiutEPEgyC6xeE2Ji7E
7PFzoMwMQxPBCtwH3NIg4AkYoiqkhD3J/LhZYE0mWM7E/k5nfmMv6cMxlOQH
4mSGSVJqhnUd/p2X5/oSYIhocyI01I1qdVXuKKOWQFe9auxus+R8jrRb9ihN
Ke331gWPwe061P89dld/OLbPlsXCtvaLwkAyQPAjK/UDRBxyxgtInJqVtBy0
w7UW5axui3EtfvOXoH3i4mVj7xZ4VnvoGuijosZjOEK+XgFN8nm3XLGcTdKo
36b3LPhozUmjuRnweCstMWxh/yh/Iu+V3RXNbGPkY1BOYxL8pKmZT/WdqK/r
ME9H7skMSs4KkBnFR+RDwi51IhXaIUUAjqXUFhRR1u6gUewe+Sr8IOOECfdJ
kdHZzl9z7nKdW3RIz8JLncenvVtXUSmR8W+4l4aSGOhf9KSklkvBpOhSGDzg
E8uZXl6Br8aRIHGjl2kn/Zy2+UrmlpSEZf+M7hqFHHyXI3qh8WTf5aBCmDXL
9ea8nBl/5Q0KdTIbem7Tz2fknnkrOPkhQ6G5+pBV2w60/GD9lrx7OObX4JS2
EqyA1kpyhaOmo5+dCqN4DvpCLVxiCqk2ncFHg3ScGu9Y7f27Fyp9ELpSy70B
M5vkgXcAU3kEojZbBdcYaYBSUkPYOD+fcCpvwhH+SLhfWDB4sIfe9uX1P886
0OY9Fz2Klj1snkgJUKla4dTNr2NElvCqc6IG0sCnrK/134Y36Qj/dZ6ez8Kg
Y4JoKpjdLbrzRANgYiYuh+taUzmsRv8pHY1SY0aGZKAfU1mlXuf/u73NLANF
WlE9/QDbdyDe+9qKHZ8I1VlhNPrdgajoX4YtPv0COJl2EM3M9HdNL+KLvITL
6goMbSVf3cpHxHvtOfXVzDPvPLA6KyyghMCyfBxOViwrPY2q7dR73aNUrRWH
eVdMqHfNBSs/9m5wK2jQp3pg8JgXklBoiXZ+i6f266LNF1X3jKlLynyh91/s
mxm+sodU9uZdG1FlsvNNxaxKa+PwxjOZ7MtjVYCoPUZiclVL32ObHra7XOoH
CoL0gSVbaUmRfls13/dwf1J34v3NnI4eqAf+judcnUDfdt9ViizlwLnoaIiN
Y/DQmAwZXWUapjLI82t2vLCGUgNAbIoHa2EOV5tOy4jOimBtFlLcH5VICrPl
21MZ9WrgmUMKHd/k0Hh2An82wU5MABhp9CwQp/+mP1A3Aq3C7fExNYDNcEsR
0AhBRqY+qFTXD1Hu3L25FN7eJS5vAOXVgUhjcyVA7zjFAqeZlp4tHUVoPR9Q
cYPlQSCpLTRBeyaglgSpABsfIje2HCsowxa0tkv6DRFmBiKj0Bxainfrrd9l
MsLoOw0DCQ4521ejZJyx1zxE/jIdTFjiWqcV4QNPZmzzmFEUhk4FiJwYKfof
8Q1Ft30v1pdAGpZ5z05mhK3YelGiPKQlniwTGqEYkGyxQ62uOQtiDTkgq7Xx
TMynHp8oEGXb0RPcouSUOQdUYPriNJap+zmLbRzAxg7wVnTzff9xr5ZX2VTc
T1hTMrS+U78XrTV+pdiTE4+M2pVmx2KhFW5mDOlOUuoGvXBn4xnjV2IovX5F
CAn5dn0YD8yQB82jeyfFUgnn7QGoifc1U8mWY60s4w/PiPbiH2GKEQFMbKq6
nTn7Tu3dO46vG5ae26RFUswIGvZGt9xasaImM1Rg3U7IPasBDDb4tbyJpCfL
qcMg9nB3eK0qJY5J/45SOcnH0E/xez75mFtOWQ4g0oqtuuURo2A6rVGaHBrK
2ALQVL6I4IqtFuop8LOzLzQ/HmQJcLZ/y4O/QSZkc6kENd/mxw7+i3fnOoYK
Zwr6/B6orbOTGCDc5PwchTZeTWkNIXE4pl4Ox7q+FlOI+xHFIXX7YhApHH5Z
R9U8ptxSV1ry98MlbDi4KHanNy1Tku68xYMzT6KlAJoE23hiGqcb0M0La9ZK
l5JXRcbl7F1fVVASFGprW+JEZgVRZEIzL9S0hQaTiCSNfhOlNIZq0SdBlTBp
mENcWGJzgWCekZSqPQE8YL3OOl9jC3WF1jaXRHvtuIG6999OV8v/yhzxjdUj
dg2nlZGdfqV8+ykdoTiZ4lvNq3MOZunZSdf+V17yWLDd5KjkqZcx9Wkq6VQc
XUfhm7kpvjF0dDxGC95EY66yE6c7apc90szr7UyBZRVkFF6oE93JrukosMEl
7TAldP20kbTfpxIfz0wEmjf4atFSI2RGzAl5OUtDRO665jEJnpg2eECDY1sv
QcpHWtsF+/KIRkiHYZi4Xb65568MSO0bkT5w4Pd5VMvalzoaU91t3ABznAno
W/DVjXw2X5zk5ey+TrVWTRu4prwzQ3ZGjOkLN47aYcB4TqxIXPOl11jyNbKE
PB8BY9jsczXUqec0ijQEAfZfcQwF2NYrQenHQ1Ps6eeXtWrg1amWp95fq0GS
pfXvwHd6KekPZxWtdCN6pNQczCUog9fGnfbWqiqv35P4DSigrNFBVsvJGgDS
MHv2YSDok0Db7bRGeMYbbkp1WI7PLlKf6zD8BsoVkBmRJ0UwTQiDkDYlvACW
I3nm79pydTTj9vWzRGDUIeIrMAKvk68CYM+YCbjpFYzWiYiHAudS+fooaYTs
6JHHRgcPBycpw4hRMyh+V7kOPajZcvwx2OPE9rs++erycUXCyowIGAqZOwSO
FxzLYzKjRSvD5PR/VaDkQTMK+o/ioNKwRQnfGv8rYEfIcNe8avdBcpuywy3K
ci7Mo6EW7q9q872S/CPxX6zsC2eB5UR8jXWIUk05iMnrjXEeP3YxxN0p2u3K
WP0bVyX6TyNscQt3tRs0K8+2+YGcV+7vD4aYx75MbeNi/V2TvjjkzQpdO5e0
u9e09+4Mg984oRB9gSMjG3uxMMFf959AefDNHWAokAnuoQBIvTF2os7hruLE
YRqnQz3xk58sTRjiVFWuvrwdliSJS4V4ScdNXF9xq8s14OwXZAvQwdEZOZ90
WrwU+Z7KhzUV1V5z5RjBSkPEVs6aZMcv6aBSwl5LU/Lr3rwskwUjmOXTFn5a
d2LExhke1UPFWxzp40BAtSw1g1ZA5KFeVVJUJZRRaDv2iSizbP0jjgLa80YC
PsmnOHDIrJt4hjZgT2TuJ6MtfPTQz5D46oAGiA+Lf5mRWcPekS+tPdwi/SUY
3aNsz2Zloa/4M9FttcZnD9MtacWVRBBUO/4Q3kVAqQa7nnJd71JsOWNuunAm
coFcsOa8t6+7IH3Zrd23UTmPltlCpcxDZuCFkq/eJfwwv4LvDzUSVMBVo+4D
oYU+9vLyT4P9IB+hLbYWfqMJT74aXD8zOVCWuDgmakGkgK9vj81eay+IzeVY
/flxdWV8ERRJkiwnJVGUuSU68O7Folae9/DpVxN346dZK8rSEGqXeLYZOAVS
apmVeryj3EcehEtVpw0KSyqkPZNo09CUuEhwBvukm6+CZPSOmNiORusR2/TG
RNpb/ybOeyv4/8PjX6XJSFrg9Pw3rZMuN8qRiGp4CDQKyEZSzZJewRr2moFo
ibhGkc5vz1rcFPPxfm1qeV44FQn9U8gx6j/41emWvqg/Ccxclp57woKOHAHm
psbmCFSlGingBqiNYEmxwf09OrLXCgTcjwSct8GSI1zGRSVYlZ1vjLOFYyHv
0YIyPYMw4BAua5QvYhcgeJlMN8l0Zdu5i6KodXfjGn5HRx0FYWAVE/WotUY3
2SGbqifVfUyliEWOwqc1uaIBlP5wgX0atmiX9tR7IMGy+MvGiCXmpxWNqBMl
5Yg7iKKP9Ff4WmxB4udhvqeHdEXa74iDtX/28Fejiu7asgTHoc5eP9rTEjJo
C2lOYQ+LGeTU2dlLQD/3+kxdWQIOP6tKJn9MZa8a0ZYKGNISHpqbNINZjBCp
vKaFOCN+jfMBtUBppngB4BTwsDujZbcjaeQwI9w30LAtu8vAeRhzgh3nHPpE
selOcPQWmh9LMKFAyhuptem+IaIaMI6M+54HJRmVKVsiSdU1Ivjf7AtrcyQx
dagMWI/Rpk+nnkDBhSw0q2Q1c+YKiuOPR/B3Gh7d4/l/y7qcgiAl8jJ37X8i
GyAJk5Pw94tfrSouiAeQM+yQOz5a7Tipt2iNyObbvKhB4ycwRDSATU+MoHaq
ow1cr3ViQ7vJbOPsKT5Q9puHhJ3Tbq3gHnvUKhoemUvXTsAlxPlnqkFkVg49
Nd9G3L4erQoIPnpUJkilD1f3F5LTUFN9eoeMv/3kT46IsMX+AChJCEefof9j
rsKnb1QGhj9Flk1irpD9TQI9Yhnrc4LjlLu4EaVN0j+UcssO5oQ0Uh33o61B
NxQKMkkOIXhTywQIDF/jCCXhF2qZJolXMP2XttLv3ov3n4a3mlcI4Ktfheah
1q6hU1NG3z/aYrUW5VZ8gLA2sCZPJzdQxIWu61hQeyVYbCv+YtMVzLiZlLZe
NMWqFQsFORtfMlhEU3RmMz5lDp5CsORMD5katE+Rda0N16s5b0Fn43F9ciVt
OU4HjFUmxWwDuALUn0odyj2j84YN95sMVKZys04WG9qMNM3P0u3nDTLH3955
vyVrxkYaBJjJFTh3XXXdF9ON+cp4n+dzOL6f5GsR/qg1oE075tUBAqlUJ5Ca
i2jyVa7x4onzqWeV5WLN+o3QnCskUmVA5cv5y6I/mL9zPHAbGSOpY7nzkJnZ
5xGHtc2FV9LAiK8bJu12Z9ODgUiJaUFmAwwZqeCbt8lOVLkniNFo7sx65lLN
RdR0uaEaG59OkL7CaiTsgkVeAlTYpb4j0AF3yTA2tbkTT6Ogf93WooMGjhB1
qZPp8WlENyANcMxXB91laSpcOJeyWG1qC+npELyc9ZPRlszO4ynvMYUEFL1l
AJn+IEgvKbYqnuHXrgMZHOZDMUwgLkFBG/ykqYoAo4I7FMCr3tRGT6+QdncF
17ltflHigPqfEteYnTML5td05uexIh9sGv88Lgp0fHwx4ttnbzPm+C/QVLWA
pUq9uiosl70ODNhwPM+gyaNFMNFxOeZAAmwlHgqblDOWT4AWPibIA6OOVWsv
/wsgFI/QYkg5jMzitR42MtQI45R315I7ZB55ik8Npvaol+xLmQnXDJHONI0g
6KH8iB7n9n8e2r6DHsQHoF6MoqA+O2AZfcZeJdt0exdZrD75RR9kFCsgFiM+
zSQFkguf3KrvoUMnD9pdYUg/MvTaaRyxlsSbpioAcgucqDhg+sqAOGcWKGKI
Y9+Rkcg5OIGO3nf+I/GT41n1Hcd2MuMule3tiklQHxRr4hspKKJKv6T3cZLE
oEd/EErOLS7qIo7Vz/MbM6wPLlrpJogQF999r7pGKeBFlJj9y38WifE8sxD2
9h95/6gaNDBNOlnqECE+v9dGooe3M1JGf/OqciVrZ4+4QGjC7pbt4K3WPPGI
r3nQpgJyfToMXJIX/QfEsvdAWvOQ/ATTkrKvMJM7TM8mibfBqfbKTtE1AEte
i9AjoID+WbDgde1vEIDub9SQZfEh/a1aiSXfuzZi4jmSoafgub/fUFDsd9J3
iQprP9OSjojeghj+TJ6H86yATQVq1esjnLlgccNvmXdfjp7sXHHSEmfRZE9O
yn1zcPqi+ulkIZMLCCU3P6DbxFGTUD8MJYO5tjIWBGI5cCg/YJs9099/KToD
K4XBWmg5Bj1k/NWqTQ2Y2hIC6tGeLZ5cyTvzkmFMCMNmswS6mWzIKHfOksoH
5FvgS6grfm1ydc2a0QMOM7aN6/9r5C2E6dY8z5GUm2isQftZ5Nq8eKD53RbZ
JWRSoYohgsDNIh8mZSe87xY0kSCJg33q3vIfT6/A8QynmG7m3wmBzKccksRK
jK1/LgqXwgaBZ7OVr0JNlD+Htst11iFF4mUKyDYB9HZmBiUx3d0h0MQe2Fwt
tIeWj5YoB5lZuz8WJSV8PAqfFTB7xkAkZawQxxZjpETWW17lggU+TF/kid2a
nNlZV6ISs7xIf6vb0rcbfVCGP5PBZPNWa/Fi6dsNfabXVj9AIBaKlwhiAruj
RMcvUlnlFAmWlsizYqiGrAV2MhfywreuPXSdYHg4esQ0dVjkVXkMqavkrcqP
vUrh9P+WlfdzIBZEJNKYhhQ58oYx/DoMKUTaoJtwNOnJAhDYvoqFbGCDPyXs
Rt5iibW/U+/QNu1H9i4EpgHjrKLK1NjGhCa17+i+P0nzUBOXhF3W2hecttym
bv/qSZ+6W0vbRUzEY/Hjh3SfAazh/2Yp0ju1uGrAplQ/hH+HWoyifd4229nQ
+oqetUyGwt9vVHb7LmeelBiddrhgGcdopTUcqZz0x1Bqpqz676kzaMTYJgyI
uVxPf1UzUFNk07DDrEFQGDnsJhutKcIIHJ3TciXcRkcs7nlewgxPP/beEC00
nLqZesxSRKMyEBqx3OI0NNKjZPPPsw+HEBrjBIrs7xS97tL4r5hfdqPI4deT
M+yMy/b7tzDdZIrZa+tLcesQ5Mfi8S/O7s2f9lwBbBuK0uZQ7+LMz1ovF8BN
xwm4uAEySxFLG2m5iRtEBRsAkIaJ2Yv/y2BV1Xkp8+cMwmMe6ABjd9gBcbf8
lSDhSY7SmaDsEhyk3mvOhbpvNZvPxKVT3jUDC1GOqppPE6qfiLn2a6VHuXqi
7X33Cf9MUVkPQOFxG744NgLbVvlWunrHyrFBcLrqsS2N6+o3/4uVLLojPuOs
DY9fQwcGCWVLL0QSDx2CN9QFJFWilQoadFU9rQr0vsb9Rjw1LIXInvnUggEd
ehbfrGhQcwSRuYpzDCeBzA4j/sNvDuWO0UajDIAJvUAlUy4qVJTKJvLGYRO6
xqVnb5pN4UMGbXlhY1nDTDN1CE9K2NhcLH+Ingy3rZ1WSfIFE11fJ9yjtImZ
XqepnN4Zggx4XwUWMWJ8oIs4QQ5s6cxIbocwLOTHIbkEP8XcLY8DaeuYNCZG
mSbgDCNl1WiDWl7sg+qn6NqJB69l6JS2k1lE6aKY2wXqH1sqvERA06MJickO
9Tw5TiRkbDLytwbOaG7xtPYbeIeJhRSHtthglP5MWBQ8IsTwaevF3OGmDs5R
ToA6q8Yd3FOzCCoS/47ydnbFN0rbKeNgghAQCG8NhOreqnImkKbqG6zZ/9Le
loQ8WNKVELBGoEV9T/J+h9RsHElHTBTgHhETx4urKKRk116bXiAA/bVgPOYY
93XCu+2Bx5BKqjAfqjz5amm2YoUqOl5HEjChKY/yQJblVJtRmFpDXoetETvX
NCUqR6r/C36UJLw55aZgMf/Hjg6mct9I7DTIDJe7oPSRPEgHzWPewnoXWLmF
m6dYIko+Wi9wScPOqOvs/6Teaq/Ny2Vx6DOTiveVUPr5vxGxM1NU+yPfmlKs
aEjvFKD/F2YQBYp3BvWrvqRpH4DIAA/G++zh4Q/ThhGHE/umDwkWf23jlWFX
Bc94sq7bu0JirUVEYCou6M98mLNrMRlIGHdougymVfVUTq59Xj9KMQWBCA60
0gx2z/+/9kxWVFsys6lThf5Q4Yzj85O7acHIwDUBut1fkvQQl4I7lJ7M90AZ
efYTpgt/NG9c7FDcqA0yxl+2zmcUM9aB6eTJWOELExlcRO0BHaM6EVhvdzpD
IEer+A456QDXwhP/36LFNuCROPHo2Mds1WGueoneKrkuhBvna8Ce1hmIhYjw
i+a/paNpTdY7r+8tK1Nbz7l2Z4N2h4zr/j7pLax+LbDCqcuD9Gwh5Z7AYHxf
TmNB3f+jbdEq9DKhmGHS1RwPWiOsLy/jNCowCA4kH0h7MLOeSLn+wi9bZnDQ
9vhESvWHBNFRIA1hZzbXyKj3/v0WWP/Cc7hvtAuipRexe9SNQ+LHEVTih9Yd
/RefK4Suy5w997z/kJrDZNPnKtekMkiih2O1nNJULykwXEoSd5MLhXz1C+Uu
4drAjWE1DRORQygMTcYZ+hkbN5MlrpAtf0eRW6OJNWN0cO91mv00mGbtMkCU
QPAiP6gFOmUam6JGr/liMbZOLamnH5DWqzVALyNs5S/28C5fCPosy3qV9GgJ
eMAJ5d/MY/Cpbnx6wQAELtR1M1a+2y64WmZZLmoXWUAyZeVy/rHvxnyh7gs4
yJgpASCvdll6jzIavQ3aHBhLQ7aJBnOczuaDfxAZ6ry2xcQ0WYVxOx9Srk7p
KhVtsiMifqMke/fNxgBVvQ+2vri/JRCa2PhojXGad/QMHgesqooooNtWZTmR
SFIc2QsabDI+CYETwOYWfL78PATXzPU+h70naF0RXvIe9kebm0EyNt1BuY46
Ekp16HOn9QC9s6PH2kj8pPJara1d+ANoxHk35/xSyVWwMOTB/nK7sAEvnOFK
vbVONzfDqHaWId/EDuEB6C/wNhy1vfJg8P5dmGFzqpxbWIS9PyMM8q4zl29x
3b1d0B4zvUOCqoJMw8J7K2PvETr9RnJe5Nj6e3/Z0cjRCpw3AoIPL7n5U2UQ
34nWBMrHYVbQmaaoxrhu+InnQFTFS11ArAcam2eTM2dZEJyjMDkIGRXwBjIu
4K2V0YznZ/IYj6VSiX+Y60cpZJKFrIMl8OF8BgcgsQXhBpjZTajf6jQ2oj7n
/U0Vy7+z0jVRaXJYrHcTfhAM/2xFvi/wpWvG+h7fVDhMNK4UjszD3ME6OY3B
ZukhCJFQAY+31dp4dBxgHdiu+yuKtMmyuOV4kxMa5KYIYgmtaTAAlFPugDDd
Hf22k2qp6A9jN17oPCf9v63N1TRgpUQ+2QgRIdHIOAo3yK2Ua2zaYsn5XHwK
v8J1aK/rwtzt9XiEx97efThkEkX93Mpj/ODPour02tNgsDQrYVhAYDqNJQ/9
EyNiEyb+KL1vEvizTCLkDgVLOVW173zW/YzJNEZBrVQkW0ZohbnEt+RF2rn3
7sCwq5037rgENhAMAyF8KnVku/xYQbRNK7vvHSLnMCuXEn16iVLv13LOSJq4
Ss8FB9IyyPQPDvzUH8e+unPc0fNL2bEmWW8q+xArB94nqfw01rFzR6Ck6DIW
DnMV/vlcry81GnI716A+9AxkzoD/F3rHoNqWnanliUECAOD9qwbunPbRvRjp
MWzY5qlT8L/JHrU3vwdEorXj15cC2MxFx/8DzXoyyxOa3BEYPBamdaVuNChA
WHzITFUuAL9ZQ14+P9NIzi8HPGEdc6pUXwiYoFaFZdJBqzXmOkuhX5UzsRjQ
MNk/S0UxOwbNb0PlkSa18iISaEaS6buYQROOOlBwzFNpjY0QAiCyWFbCRZ/e
+BoJxn8o/08+xsYQgrAL9hfz1EeP8FWHIrXHSCAEM8mPqHQj3XMCLhcYH8v5
/6Em7+ZgSE+3RZpwsR24oQ0VpatbfoXj6kUGrU3IZvRrcDS6ZbqTwRDHBpdL
UPf3xmcyZKtgHJm1xAfcswP3ntayguUsaexD2v1rQtuG8IlPQnCIgIWfBLjI
mxSHWoJXG5vwgHYofxAMBK8Z8PQx1+HCfu45IbQLEdy4oxZrmFLerOZxD+fm
cGoLI9NFKaUGiF/YCIdpkunNLpsySlVCKhYiN98j0pYN29XIAKPAZp0uNnd1
CbmMp25pfQYJB6scbyaSpypvhadADp6yQCiVq68XSOtDAp4kO59OqVoMqNE7
F/maUmdEsh+QwHrOV9VdscYo8uNCTc6xj7dmB1WB3YQvyBM7vv1QN0/JGd9W
wPriP7kFVYRviE7n/cmzBTUpK6ygiENvADpaWI+tbFG2czhqahZt9AOR+gAS
cItKayc74oxQ5IMSbkntNY8YDCmJ7mgaGjkGbvGktTkyRt4DjUqGC4k2Yl3a
lq6wH1GDEc5qm8UJN4+KNQIQA+0o0rxcMf2XeQxiFwQLwErOLkFAY2pboXSn
QioHTrKkcM7xlLxr850bA1rmNiIt9nEUVksuCjzSSoacDRdCYPiOCnR+LLrc
qyLfqoQnQ5oEHQcha6TCxccBTnxoHbslqkINWkezQ7G9SYcjG5Vpk1JoO+UD
RCB64M3b6sP1uEyq0L4ZhqaVdHvGW8eGql7/21O0GlK6vObPSd1Cr8oAg7gi
dNNhPfJ5Pl8PVYUAnxrK66BuznP/7f/cs5QWxKNRGqVmf/rjOdase1gBtcHb
Jie0wtCoLa/ZfnQxLnQCoKkVFkRa6RkHpvdatdBrrtQlvksd5RWESpTrvSe5
UsJ6OIAi/pB25qDJWTMEmD5xQoSk2AGUm/6yW0URAxSFhF2OTS+5G1M6/M4D
79DmAcdAz0jm8zl22feNEVs5TyZGRVjsjS2M4CB/Vo07IN7AkZev7pRe9P36
RBbGgakXonTeKg0Wkc8uVdcUidS30TDat2X519Jap5w0MgjNBnpo1kA/sb7s
X5e8A+Js4Q3uyFN5YRijH8BVIsFlga9IIaajFlDgVSkTq7xNj2C6qM3TJ/1f
O3Fdmhz3phPumc6IS4ZFSdFBC2kKJiyDmuKSdDx7OdrX8BjgLPUaBguzAbYm
o3BYNrqN/m/SgIcDsb8QZ/xEXQxqFKOL1+FTGUBcA2OxaEwCbdXNRCUhZ8fd
YGA3+VOLb4zjX6EZ0ftyqVR4WFxnEwD4KcNN5snbGzscKgs67GTwW6deW798
ASK1tieTsTzKkJzPrV1Kxv+Am3khoT5ZSG1OPX6uQ5wmZaje0tXzAPFbImW4
xVWOEiRWOfxQ2mun3g5HJEsuqMLRW5v3RecYNGaiT9CmERoz4aFyEJ0rfvQV
AosElpCDn5SQ2PpZ2yev8nGdYgilIFRmXGrikP7Ye7a5s6npnUMdXu/7t+lY
jk4UQ41IdTxrRXBvTCwZmc0o1oJGcuOt8Al8rhMxf+5jkjXBoyrqrKm4O4Ay
FAjlbVGirHcBf8oLkjW9Akex9HVIwUxTziF98XO1oL8gIfpIXmFdpAQSkrIG
q92iURHGCS8uTubpBEgmzTC5crELraFpoP38g37DcN7z/xveqosvuwwqwLGj
KgAwL2Q5M6ZfSKRREZU4yrL38vM34SsDuWa4fDhIpcy7M7Zvg1Qr4ExXfQIr
THwpDUy3DTowhS8gj9lG77Hm1jiHN+qj0MuE7USEUD/Rj5T5JPeOErWuVsue
u2dUvwk9eZdI8ao09T/yHiXbJIXEtzyjumKa6mVTCe+9rat+3/X7kMTq2k4Q
1fzPdsU5bq8qJbsVd7DIRPX57i96UGgSRToFfODAdlHw+ozEgt7hv8MoyDuj
ogvwDemidTsDDTRG5OL4efW1BgIYICFnSO+8T7K1BQBmhSi5xTgWhbIbD1Se
p3bPv0QILiEbHmtIg/OKiJB5uibMgtfjRDNpo21g6WorUWcfg3BnAXf71xYI
vOf51b0S/l/JCUqoD99HPFWG/AfAbS+edsXutn86xbJKErxGDV/w2OZNL6bd
voUKmvfJ/PWvBZ4edaD4tDqMmkSerXp9KqC9HdzaIrTo9lfyYJgEozxCm+Sp
IaPIrgtTzbq9RZTSCUYmbmqrexZtfNNn/nCbu117LqwZCCIvFug2FPwR3APl
vrAxZa97CIGY+4qDtZmgD4mg6M2whTMn3FdY9sxpP1b+tzbP/DEe1d0XPvIc
tF0UufxXHwmpOz7lQXWcBZMiJfdqkAXYYGxKX/S333gObtOVwaFsjLEwPkEd
O5wrBbS0lHtlpHuRBAFZv/Lu51vGCRGfy5vnXVXkNwmMWMJV2Uo+GznDbbbD
+6nl33jTGT3Wvur1Cvn0v1b9yjRkEwyALglAn+8dh4Kg3/9V1WggfVYKMBEQ
g8l4sFit7DmouvvmOHv6dC2Rp8AxOMYZ2FFHBigauMt6W7jKiTobwayPopyr
fZPxQijOwyT7mIOQwDbqCNb0C/H+qS7qXkWTs41ynNIhLC2zQYViwraldXPY
KUNckRHii47NWlLWHMi6aVBTY4EpMtv/mo+88B5ERRPBjXR2sa1lVzm1C62P
j4M019POCS65tAU5nHaawVcI+rantkD8Hw9QxHAJ2fm1G7UimoiAb0V8Gl+R
6wOU1H3JSBS5bq7D85pCemXElTScThN2z611Oy5MJnkeTkk/0FWxyJiS7Lyx
XDrYrHNpxAx243cyhX0LPFIy3hLgOVUjnT2AkljZaRMcrkzlBJBxz39QGa5r
BslYwr1ihsxGSzHTRxvwPJRV1WIuBKVraxG8RdodhI2DdPAQj9Vb3satc530
Pk8Z3T0a33ueKFoWCVTWCPhsZk74Ur9Xv49PFAXrXpC7ahdo9m5bug23JaWc
lYSUHQSd/p4unJ5KhSxBRT2N0gvSTIk2heF798RXWwOWTDgagOeYy7gQ6Z0+
kqsMB4Y3EimdgTcmpoq0ny0GoIppLUmeRNdSxpUbYZhbIclHHe1jW695UpiU
UTa6s/NCIfNTu30PuOAJvmTsvxPWeC6Z+82hU87nIFzBgi/nzBB4bRQlIShC
FnUwlfAXwHCt312IKAu/2n40RvP3m8/JYLLgZ//jVn+Av36t6d2SLk4LNcg5
EI+6Jz4quoml1UcnCjDYBlDs0dKJJWMfAYE34QEGWt5juBWMiIhYaz7/XQ4b
d7SuVsXT7/Pp8z22SKLys65bvl7F5w3v1TMrfFbIUlh7NIHjzcv1d0fHX705
pXwy/+Bebk4klD8iAWUqMjSAgtK9c/TvpaqXHn+qVac4BpNlJYL87UMpkSAe
QVX//DEAc/WwVZwH+5ycEUYpDpNtkjFfB36Ca9hiD75xZ2oisn39vqHZc86/
s/hhNG57oslMI177bZmM5zZEAdWqWo7dxZq/4X2oZQBeer71pEY6XfBEoDtH
WycjM56aV7sRNjifZ+AYoV0lBXHw4lZm2q2UXWk21AuR0aPhYDCZERcXEPJq
NoNcdzS+evTUecG7y7tyepGc/3g9Nq7eWpZdM33tHai9hO0jURs++b1QISkL
PzXhvxG+Wdf18x6DlAGh2DqSwxDFhf4WiWcqy/QM9HrierWhCNxvXVR7KJwh
eVuebkFRLIdckgF+DMRDOhSHqKSHuDq5uV5oBlVFI6qmLllLxX1aGJ66Vua1
T6gFLlYxv4Xe1mzwD5Wx54EfXuZL5C55eY0QHWMQJ09xmHzv4pbBJD4ZbpJN
azHR7Ndral61kJPnEn+5NLeDAvKtKqTquAKIaCaJ8lESnR3jskIlGKUe4prR
Z2aiogXX/c3lQslnOZ3jImkfbG0zcMlbz9jMiDkmPNiGv7EO0BF9/gvpfTfR
lEAiTY1qnwbQpqtbuQ7Y8JGIzo+B8svHmD2ATGKK/RzowI5ocqTSbvm1vHqQ
EU7foz8wY7jKZf+QZS2rh7Jvl6+oQw4LgDtQm6Yl/Qs+TIJzopaj+RvkD4Ox
U+lTjQBZjOMJGweIokWDkhlzMjAb9xHmlUFZUEbLhsnecYYMQ8JCtnqA6Aum
5LCYRB4P4ENK/iMdYc0OSghh3zEWM78ae7sLQQorfRZUpuMEM2URJrvh88uA
x5k/fBYhU2oSt7W/Lj484SFccyny/PDZkIKqrmm9TuFYdeXHUDzyveN7dJBW
rQrdLMG4cbIZEzwZPT+ZMloaE6M2J+OAsNRV8wmNzJWwWBIQAUbbenzlrXUM
3flcBYn3ys9t4hWY2Nx+QXE8AEQtdIg3zQVsLfsHgIqrDKKLNk83ip2kx3R5
DWj28H1m2fe6ND48qjsHWA7hqBn7ccnO/T8nBiou9+0jLcWW3l/Wy+3LSXZC
h165I2yDi+cK7nFgKiolf2D3pIzLKfpylAHZYxxIR659hvtAGz7Z+hc1fZOi
rtHcoGutYOrP6Pnz6L+puoAOZHcNHthRiYaHWHm/+3IyAH0dgppFzVZwOCRR
tDE7ZgHBv1SpGUqNTiWbN9cKXJzSundCiz6b1u4UCw65ogTZ4fUkHgWBVz92
O/yMqIHwHRSqN6VH/YXzy8FpAt8CIR1BVPFHJFVLPFc8xN0yPluDyzb1aHR3
904n+xmJQjAHwtUFx7mW4l6wZNnqxwlYDvIq4c0IBXMmNGQUy8IE5MNGvh4i
wmQ6QnXQ1G4WKJx3SZV2vYNGlDfaUvE5kOSfi4GINjdrRZ7IF/WOm4ZQGFt+
WD6+0td7NuzYjneWICCtdQnUDHnSoPiG7ShL7V+PTOKCedDdFaQIMt7PlCGO
HEAn0kXNnyhXG4shVuCjFjjpis5eqbmMmr8hqMjS06qzc29ovrBlqk9u+xlY
DL0UaV7ps2hNDwLQ1OY59EHdAg1xKInla6Qh19S3I+wE+yU2Ld+nB6BjSTKG
2IIiZmWwwVRQ0sqFlvYQ5sqBS//mljchkgjtUaxkfwtIg0way6RBWTtfUdMf
C7LVc51T2KN4rssFMNH3aWNGeQcnUzIHy5ytYb7UKovoO/xBBJqItS5WCdhZ
8bRgPK24ojLJZHKGHywZsnrVFLnR3VQYyw58HPoWtUpaMEl+tLVWNhq/ZnKT
NcRxhluyYdhlKpTUK1KfX0TrKlLnqmOKa3fZcjO5AIv4p5WNeii9oqmrGt33
BMQgX+LgK4/bonn2wGivpRnpXSkIee0LIZPRw4brBrgF8puuzOWDc5ZmuKT2
d/pmSL8fCrOOD8ubSLoYQiFpp4Rx+4dq1CGX0ikFOx6WVwNh6lvB6yznT40X
xFjDOSwjTZMKeACJk7fErgFfThW3sYWtuUoYOO3es0ZzzRmJDKy6q5K4RWf2
FUanJEqldr4wS7vBHaNbQ85nmfAjh6ziFxPpYPLH+c9OesrDl3KVVy2Y6NW2
PNeo94BSp9Cls5nqSg1zSvqzBJNoKAai+7T8QGjTTI5XQLRhB8fO/ZHBi5hz
JtO5E/1n22AVnITBxCl2Wzd4FI1sCrSG0JmJgVOQntU+T1cQwdCEJH+bS1wP
FXI7ZjdRR0ACwJBxSWLfFeTbYDTDt4nVeFvmiucf95eZj26NjuH+ZYxJ1JLO
weOa+KVYiMLeJlOJX9kwB9hO22NeWQXd/DmdUgncWPRLZ1uFM+u2gqtQokgD
hDM/Q5+kKzU11N1WOv0J3P1vnf4QhecOkeayZmn/9ZpeLKKGx4xXfwA6/zcI
Ep68T6btkjw7CR0rZbxKav/BLDW5dejOkGLg3HNac9OkjHkDH9XKisBT2UsE
Th+i9EOChIW9C+vsGOs49yqyzX+J/AOAFhgWs+I6cK+mrhyzsgzNpYBqQBvc
f+LSO/5HZbxdC5hgNP8rvEKZqYvis51bK2cXYBp2zpR60uCPn3gUwT1oNFPP
RUnwQU4kKQ8hZYZMqjWljpVqrw545cp30lUTtyLwDBH9DI/aY2EbtZBJpIpC
WApOK291joNZLV8Y/YU6bHGjyImYxHVSwp27QYvvwWOiNSaW/DNxCRu69ZXq
NqV5bREVpPMP0/sFm/4AzETn17MTLluO5cI3gHxQAhcLr1rpPl+iY+wvGygw
eleu253BBRnYrfKCGj0VxsaxfhmCO7WTKapVHq4GPhtxnXJvw97pp61tfvtd
kqg12qjJ7moSjXIhC+fiL1c1D4F7YS7yGf0CxcJXdv8LoQphF9I/UlZNmv/H
7r+EoL2GQoZZkQSlNh6ArNT3/tfYygh+p9Rso6/W2iw7OJx07z/qfpGkPJ3E
kDtywrqhTR5QIwLMrI6FEIqyZHvuq95XP6kwZg3gys760eLLCRmr9o8a6mQj
eTEqMuMOssggMMh/8XweTbqOA+V/AWVAHOREzTsfOZkD215M0H2o/H1XI1Lz
wLiRuSM4jnytgDXtWzpHJAq+G1hcJrH7DzOsq3dAL7ciInRoQeyhKkQChc2E
5GTq3ZKcn/sB60HH/6yIciGb9giC7Opnmp23ZHHURE9bnRr5EykskjfBmDTm
xs4zZgDscmDjnFCNHMSpdQc22bwT/P/bDc5pEBI61C2T3WPYyvXIAcnaK10U
+rY+Hf1DdWnDWcS9LSz8CmXyfbghBP2Fz1jUhHPoP3zvijSddbd2c7aht982
anTYrVId9/bjBiKxEd0RJ7BboqCoBDOqsZi+UWwGPSEV3+h4M931FII46ENR
ZPVuUT9jHWKkKBE7gXo6tDcrQktErqt5L32DwQ9VZgbBnuk5anz1/TrMQjdj
YyxK1/zLuaDVaXPVuP94WNm6ZaRztuxLUF5NMLYxm9hJpHMaT3qXO7wUmNdQ
gKf2pcJ2wRqJM18rJ1lsO2E/w3cBSR7FJc3+FZcuZMOAflQauVtxt+hhEyXJ
vPTR96scq4y/FN3bNz/Bb8OKc3GFY11etMeBb+7IALnaaQwPCka3aMftX8fe
M9sGd3iu8HKv0wYibBlY2glgGI6PebjJulBOMquCMoalmDsYnDB4o9tkMpSt
h3j4Gv9+Vpzpu/GSbQ5ru+3ibrblJlawH0CdmpRlS9gj+87WbAbO7Q0df18d
d1WtdUYjk3Sqp1B+tLIyVFAAwTxap0a1HdPK6J+KgwDOiqjWyR0NOiqNNio0
gt4+7aEymZNoTptWjEnMR2oOz94gi33tVGB131A4raOiUpGchL7tIpfjK2h1
sjJqYQnyXNiR09RhVlJCfBqRUiVw6n4Yb7/r2+UZNjEqhGb4VwaCKAYT8mEZ
5ec1KMqkN+EyQ0kcaT6wTNx2s7SpbPgmWP1YHqEIDNrSXdQFEyszzHpa8V2R
lAKR6+xVsiTLiA9UiciQVT990+aGTsGofBxx6O/vrblERWl7jBOQEDbIDq8u
wvslyI520TvcO7RysRFCRdEtqsEGMJZwOQ16QcdMfSatjL4Cj4aL77agRYx3
j42ocIibqGzYmKZmCp7WUJz7qgf/0JTY0x/MG92CkAOrw+XsJ23GwDt1zyuB
Yo7BlmJ4wLpePagx7DfHp0HJumcLHfb7TYd9DtFmF0opougMRIFJ9qzOA8ud
lAkiDiQaRE5weWbIiqImbcqQkXn5nO836vHURgYF/gxFOycx4uvX4yql7Y5P
Jz9MMsXM4REw/cr2dYwM2EtxRZD/fNt+TJMPw6JTQH1xkJnQUsRcNtvcqYSH
7FcWpTiN0J97OU/OfkoPDr2JICIPie7mZgf9H1Fa4fnIoTWh+uoAi0eewJzh
zs/AqHtCafMLTJd6liTi4B/WA5vuInIlNE8M7SW/yR0LBFcPZSdX3i4ip9B7
6kpyOKHiI3A9F2rmZUyEXdxbdz1GMY0W6IMR/aHCJaofDzn+MKTmH9zZADl6
UxNJTtc9Bx6nK828Q0SefQ85EeqWsCZwrkvaF1LJKShUzUMqo5y0rPFWN4j/
Drk5o36CVkMi0HicKjGhFYjpY2ByfADpTv9qA9AzFgtB5htc2BtTJOca95ie
E4afQyZ9AKgwd+ndAB3D4WZ9gHif/sAnBIZJZBN+/4zkBzl/OdN9d9VhIrKU
rktJQ6BMJe+dyn0hVSPqqT/M+i4OKDo17HpWXQeeTJtikybp3ieLREmYkhYC
YtjOO6ZXvw5cQ+1UUKFPo8DENKYG997MzBFQDrt8VQNx6GkpE/gZjwgdfeIT
JWrqUNfQpCErq/D2PoCA+r7hTZTPLfUcNOwa37i7AtOk8+VW/uNq7IuTkrAU
ObqkRRjnGwZehCRM+y5Be0sZtftLYPOV9QSi+oPYVy2ojiQgDSFgQNunGprN
skLk/znA/PAgfaLMyRPtT26TAiQdQh3vfRQZE7M3G6BoUXu7HxdW+MjZ0VBL
GezxTh6Rq1ntTi0GCAh1JTG/qD4sCGGhULjNZKkWyZllcCYMFJZY3ReT0STC
vzEwtb1ZQPp16CNzGhRqpP/7EeMLqJTPnh41cEo5pmKNUAXxL1A8rkaSYAqF
vvgQitATbJcBqTu1a2XjPGITIPVD17Zkm2hU43S8rDWILqGb9onFVVkKW5bq
64/ULT5pfAGyamOsqB1HVFQ/0ggcd92zGr+vanIP4DXsj7hg4N14iDsczISM
pL0d90F6ASbHJ7ZO/GqBKvRW4Hi+1zm7irnZP0PBGqn0OhHy39ax4re3YP85
t+nW7YhyWe3W9fPiaKdXHd4iAajRBEXVaB0rmsHyicrxSag2UsC9nWVbLUKc
tKZqsesLX0cqngGrEjfWB0FORUXYu4BKjmpEL4Rw1ircyIS8LLD4T4wkpK5T
7Wwf6IUn2nZtL9ZMhQkLLrBYuMtCas31H3uIoBQsImADRgKlDxSUNFQ8vCNW
/ns5mKEER774PPyVJjfAA6HVKYNvahaLIeDnQ06gvXDY0MgXllCIoLa5AYCU
rdXhSbd/CraEQ31AB69DrB0+Sf9JO3b6tuODu6jhBotQxEzomqKy9jSTGMrO
2JX8DbpgfW9W7qawvX+vWOGGWu7jM5cATnLvtz024JBcAFRqkQAM696HSOH/
iSkbBlKoxvjmWLgroV6zVgRdZx1R99oMYxSoixX3WVW1FR5MN/OMcGgbbBKj
nL5cXWd5cJD22MnVqe63J1jjWFAqxskk+GmeQdjBcywP+rTdHPzoOavjdUvj
o/w7Q99w7d4aZ8qwgI5XCZ27CxJt6JneJ7ixzyWGWpZ6CvTGPpMJXII6QID5
H2vfJvYLMnSwBKrDgsuUrYQYyqWfPXBDw+RNSAu8kZBwSMCkMTULjp5jKe+P
LtgBwxP6lkbiPcu/KPOJxx932CeL5wbfQHmyjnZ7VtigeRLSPObBlolyLVvk
e/1FAYdvwv+CWWj2oI40Gx5L9dWWeTkCP/zBZgETqNedWlDNjIWIoki+d/Eb
UbVungoEIGoMcV7wOZ8Q3DjqJQgcdp7DmBwYQ3tMo/okRqBXsmNEjQ8ZPllZ
W9DV7Xf6ipdV2Gj1dz/ht4YVCRBXrhaaxArk04Q8fsIhqUTg0aos1dOR7FLN
dIv+QiD48Wme7YwadICHiOI8/aF/JAlMgRXc6V9qlD8DdsGo6sh5fsxN/kuG
0auqn7/nfm9OBGzf/hWt6Tg8sJhsf8snLske5S51nWOA7JNmALCg0YhjJ+vL
XQWqivkc0eGliN6ThARhLR8efO6WNDaPQYE8m4izY9jbuFzGUkjywDFp5Jo4
TEB5jMLJHsMvwF0MMEhJJFBqR+Cc2ERaWKSsD58y75HAyjBCoOPqdhs5PQmu
/FUowC3NnhNQkR1WLnIKQ9FLP37TiN9xUWh+QII6MWdZiY3hbENdLvcCxKx9
9JEZpGbyA9acvVzCA8WzNF+uYUzNXu1qrlnLmLzv3N+xzAHYYbgIs3/l3pQN
LhgoDfWFcLcPB/AypTafUeEMUWKkdmXqSTUdEZL8rqhVxcfvegTQ0gLymIHu
AD4WLhw8Hb7I77JQ/5Y6szETKkmQkchgYRKY6Ebu7WV95VzgQar6q5PLmq+A
2QLNJ8RN6K41BXGntIwtnd5Dk0rrheBLO97Bcl8Ytkq28ZYUNGhz7JViMu3g
T0R8oM5UjIWOr/wliouPhhFMtNRxlBkkE7nlMiMgsaFSAnqGiS4/kNA3W3cK
vQj5pQYmeRxJQR0kK91/evbzu4nqQfS15Mn/1toyeS/FW0VHsIjRxdYuZJ7c
jKh18cfeJ3Ku/sGHFgPf91FzrpOtFfDKHeyZnCqREdjkgxLlzbZJECqHTrKr
NMrNS4ZPR11vUD5sJIOZIvJ14qLgaUYa3l3yX4nURp2orXaSzAZ/pxzG2r6/
v0Ztm9v8uXC2gd+EGonXvTHc7A7DjR1uhZ2y1hPdG67gmte3p+aK1ftsCrco
NRGRdFe7npU/p4f/XLmRImcMzHuFnyWuqcSXYNvmmP7qXkclKu69dECEMe2u
CrYZCJK8RcvMSRTVDki7uAzIsbd6Sdg3z54YQKNPQR7YCfSGfa0uuwyq89ro
3J1iJIldWTBLBLRdza46GyFab+PwLIjZgNOrpos+E9mzxgn2SpuBpmaEstaH
pMNcEhq38EVAFYScU/Cn7EybH+ReMBRIUc1r8PKipE7s0WglDYOQ8F7wkTEj
yNQez/dT6FweusUeG9ssVsnsVe3JoNnk/0Vo0+9++AG04jdi+cjLysYEGw7f
L71rIMdPRjvIW139upQHW3AlAw0FHqrWUmaGfY0B8XkFUQ3BTDDDaMnZcjeE
m+AiJjrWhan8wYXgFySE4UXOGfg9xTG4xYatF8mbCiTmx/cDoGQb5nMAXLeR
PzdIIMbTsLaA1MJU551CCNv7ijdTorjGmmtdAbX97+rhafGb2xBnDdsh89h3
tTn5psG8/hXtetJL8jX9xm70hiuW9pAvE/t/VmlTMeCBDowwIDQbFs7s9j+s
lXn3QSgnkL64bTvzxppRLmV62BRZr6PxyiTWS/pnPCq4JnSCgeW2dIWLmxRu
C0jBZT23Oss8LqfevLDA+P3+0ZmG7VfuHztHp6k7u1QphoNAzQkVJToXD6Oc
8M1+GQQEriypLtes+SW61otR8M7njmsXXo6jXvP19okLsJCrSObm2N7dgR5Z
6BDVGK01jYSbdVek5TLpKDlNSF773VmtOyWnLX5FlSEyvrqaB39DEtkwd2mn
toWsr8DrqI4pwfcngdgf/ZEzrO7/ZGV9M1pAqPJkIvEVknY4yOWfQe1gwXb4
ON5KsLCQ1ysm11804FiilKm9ZtZnkW4tIiEOu2ASkqinj2fvefWWW/P1dEYv
e71yv6RwixIAjv6tajhoPLLAjYYHMcXXiH7rYZM8Dwnyl1SryHss8fJP6eC3
7KFnrTGqoKE0gvGpPJPm4ZJmoAgsWFwTVwQrj1ZgDQLmyN3bMxd/jJxqMdr3
o8vAGsNh7DZNOdbMmNv66rbd9062bdjX2SeZRrPo5m6Oi1XKv3uPzcsMRPgo
v8dc7mmC4JswsABXun3Cro+aa0LQTepHyK12yccZDLp6TqQWOE8bQoz0wOXT
s5RslICEhJZEQAlVOpqZwb4Vq8cAa2dKHG5pJggOQcsR08IRDKkRu/b3Xill
yWjNyU//3MzYxRPU7j1hCciTvcLOZb60WoK1Z4quY3FafHM+08bzetOMaq9B
JokjcvAqp7YhcVmaI20rzwZjKFCzJuoV+fJgu6v8cXm0pw647dYpLr5RRQoM
8pIM7CZKWsXTfwZSjd+2HPO5NVyipXbIhuEnu/sLi5TJhPTgsoeh6JgevGyf
lY6xSYKdiZiflmoZcj5U+qtBDzUX0aGh3eIqWDzxf2DXR6G0tJc4vnaBthAK
VkcltbBVOHxSzdluJPs2C4mIcMfaEIkVQmcgRTgq4xrrl563YoVclDiGLL3O
nETAPNMpI3tUTev0SMD+ZOkq5cep/P7CJGh76XoNbTfB8DRaG33oyA4SiuLP
a34PcEGIQ5Am/VAG/5t7jmaM52ftLafNHzbZTaf+1M21BeJSl+yN2LpvaA7J
cAk9IhmwqcE9pIImhErLlpJ2tQ1mEhGM5rqkv6c46In1xkA0ObA+ANOmVXLL
4Hms+58nID/YD1JwXIpHpZL52qF/K5TVyKUCNh8oVQnoiRMi5MpSylnIFD0N
kfyb8zG/agPzuk8eBNlPWFtOanQX+FzxTMkpQGAyUCD26cu8lU9HrNNVx3aR
pG73nyknt3jks4FnWod5X9/jCRqTSAWdWBLnAnHK6GQEiKmUXMiOQ2RCpGtY
atjteirvDTF0ynH6osisR4fO21Ligjb25F5kEWQbbT/ZqKFQ4QpsgXcLqyBK
aOECK7mL/Q5CnP336Rc3jyBQJGaKUeMvzUlDio2MJdXDKh7tmBm1XgjSpRBW
+cmF+AG3pciFIQZ/up78xBz3VR78D2LroLzpJb1LaL4yZKKW791coRSzTTcz
QXOBB92TkE5pxO386mRTYkyU3CsTdsvNvojlRDNWtpKGjHzOeiUedtcDLWgT
e2QjJmTYw5DeSjTno7SepkeC6fcoyVKsxYBhxsjZE4jcNv7CCAacoCHrhX+f
FAjNOvDPUGVoFv9arhL7i3ZCAwd+oxXcWlab8iJa4Hcqjy6j36hm0hCRdfVl
LcMBLoMNV2bVKkpPIVw6ENW41oTgNB59xOpEmzLQkZIXQhuq9V3zhhbkDR90
Jf/5tt4Ynh2BhqF7yyYKktPeuWfyYsk+NoN1E+g9XIQ7ulSmx48VScfjpocl
K9lj/dJH58ibv19OFAyyrqNAof1+KxDvhz0zbj8kWkX53P7ZKu0TCRUrxm8o
oJpAfR+/Rfnx7ZvhNiLmG6rbbFzjG6/Or8pcpUshc1jG4RILGc5/0IVkDRAZ
+gXQZzeM3SZkC8SH/6sdOu3VDgdXdoBfFVdh9F1XZG7wv7gRT+CdxZD5JxFz
PJG6HDf/kyHJCfvqDBMj24TrvBz/vkWi1X7V4XBGCVSQ3iz2N70YNc6lz9CO
Lm0somsFQi7FHEoRfC+nmFlL3b+ILKjirO+Pyd3PCXvpoG3pgPxyQC6tdzfh
QYZVKp/hjKzOp74A93tgirjSmMYOqt3AMB/5Mn5DgTXCq+Z7VYhqS728W6tH
ck0cGP3R63tYj/LZLVquAbjsxdnFuhlADFwEmlm8ggtNmd6vFXZWndYUFE4K
4AgXCxXMPd4pyTHNSJmWWctGY3i3duM3bKL291u9kO6Fvc0Po+/9p71WVOjq
BLlumgpkk7eg+1n7ZRyhNj1AVdtkLJPyfnDN8iDYEqT5KAmcq5y/ibZygtPA
bYMDToflSGGJdMBf94TGm9kITnNdCmCBeFe/Q4xGAf8IExakjE0PjY0Oqm6X
LzOeZdVehYsx6+DEHH1rDHSyUblCodkTpr+HbwNeDvVFZCAxa0jrmTlhHzne
tHrMXwYkwHGbstlj8iJxApXZWBcAfxb8FLafOzOFPeZC5OPjfiigsua9tKuw
r3YEbIfsJladVHv4LSBs61kP/FqxaiEBZfN7z2RnN6l2nKvRlCzcX5rp2Zch
NVzibzzW6JYc5uxQQR9w48nswyBQ22HF9HjU8Tdc4D1LkiifKQ56dVJwaF54
NmEaCOtzOSk3/b6vukCr6wt5itvTwUPHxLbNQMRsE62xUha7ply9KU3FzPeC
tH18RVt6QJ/1oGI46TeTlf6zFhBzAMQy1/4ZT2HrxR8rewvrwfs0zwG5vCgQ
bcuA+tx4wCtn1uV+4Lh1s1xkc4zGDNbROLFW3oKRJLW+9PhPvCPmmqL9+eK3
5/kLHi2MQgMT/vpcDsF0hu3ShBmd1BXwj4LeKwLDhO65NclI6c2xpd+Z8LIE
u6IUI/K9XQZ2Draiv+SYSdtHjerZhznUJj52/tt78Dshmjhzn2BL16nF95cZ
YY0QNnZyChFFpc5t/T4FK8NiPHKU8lhmf7xiU+QojnUD7J2nt55Lne2TznFo
AbLLfYrT6ngfnQf6D8mN6NxXb1g2K8oEdNPTHJouhsxCDhPdXiXml5z9vHe+
Q/sQ/8TUFqPvr5yQSs/vBlyiR1ZK9Ghq+nF7o4R5BV0Yd2k31iNRsP0ia+XU
OXJ+uJ4fqklVB46Src6syvDRcxXql2n/E58Rn/BK7USG/Ys2nFuzopxndsfY
vNBhbqkiCrg3h/6V+rNMZMACzeet3whPEqgIvp7C2UdI5jXgutw+WIfKykzN
aLG+qlVbRXFW4vSIGsy5q5FUInSOKfmMabSxF+tRBy87uh9UtEckgT8qPpuf
JkhV5w+Sj26wkyvjvnBQabmQe5aZz0HbA5SlLBRYt5fXKA1xHbhNxJosucKc
ixlPBc6XmNWXwcqlXIfPRlnY+EvaswrSoduAu2stOQhQe892WU3u1bYUt1z9
0Jijt/OAZg4UE8X4WjtfCsOoZqNn1/FbfHdzDABWqXzMF6pdB7oj3xT9GKb5
6vic4uKtkSUDSdYPJ16/QIlD1fGDDKgeJwhrtu3EIrJ5kTcZF73fUQMRAVUQ
wTkgmAPlp42uTsQyez7clS20wm7WlskbaGISdHjHQQPCnawsiZ5WloMXy9zQ
Y4Le6OchwnMBShIdl3MLg+KwPUf64HazCeNwnUC+s7d5Y8Ag/YlIOVZjq0tJ
JzDcyqbZZSoLO38/Sy/JDAcy303C1yndIAcG9C4dqjvBDiYHVCUPRlsvkzfv
foqxRGdKRqAl4KvNsBjRhorNwVop4w1YL1g+qfto6f7gb2l6MllR9SEeNrO5
r7/1r0Ox0jEB2VUp51/DUuKfiSOIdmXH/uGf2sRaLjMHzGwodVf0NzGB2uB/
iThzvfytM/38+PithnU3ja9LTQvz0BP54LybxBbBHEXsllefkHNy/2AsFE/F
zqOA4PeI19kssMI3pZn7IUY+jYHPse6BkomcgmvvAl74gCmE+NsZijzBgUjB
PKk1F8mpJAemE2UbnjzdqOdDEDagHurVLa70hrpBbBQh5lgMuRno/kiRKgaG
+doqfocqgkIHwT03XHnfG0qMhQzvGfAS5EpeL09ar8ILfnDbRpJRTwHByd28
Wj8Hd4GfjqQ4cQ4NXOHIh1ye2921WxkFZB21t3B6BHUe3dwKxRHBDiIA+Kb6
IcvocuiD79CP+CvByax2eek4nGxEO6YKRLDwxIZrYwIrXQG8O2YZsZM2NTN/
1QIh3LRfutiip93pA5athsljoVROB+6mCvh/kH40sL8m1i6SppIckshhx0Jb
SGzCNYtusunA4gMZlqIfteMjTQzgvGMXqej/jSq3e8wj53UmzQohwalPvpNL
wqYLSwT59va7sCzSYW3DAv/tVYJrCOTSi9fBk8v885kiw75TAQrFE1IFzdz9
TFtgh+qeO4cfZq7jB0+5lgGD4HIKVdDprbgFPt7kjX8MXJG/vQ+RfLTm+Z1n
X9tCjZR4axAaWWHUS5nw2fyyYVpeQh1SKe1RV2DKP0BO4MtfQU0rySPEEx8y
lORttrCy3NELBLwXeZxmpDAw8xRP96/p7eAbA3IYyn3Y0YowsaDNy2ac0ZQl
SA7r0EwlZl62u6yF2dFiWvOLEo8b7XhHWskhrl2Qx60UR+1keFVRFbRaVXkG
KqyxdFGrM16MDV/oEM58xNh6qa3wAxawWqeit9wkh+Lew2Pe6VBmexCz/zzr
8WPgb6OXJkQz+0bgGm4dm9NerGC3NMjT4wlvCxrZfluGdfUUawLEtNBDQB72
HJUB3U/UOVUt6M0aDJXYaXWe570V4BkYbt1VeF4sTdjTHCy9doG7bQgpIxPV
j7hnHHj6XxgGnYTjIQcVvh1fPdh9dFfnMEZHGCJXGr2l2XGWM3Y2EmMj8A7d
a2nxcpRiZVwhoJRH5N5ZoyXvYuMkZnXNefNtTuIWd/eR4pJSzrKABGs0n49Y
zQoalVSE928/GGPpRxNfDPsxWW/GPekUpQCw3WhtNlrwxTtGOHoO+PwDULKE
08c3jcboXxoAgiJ3cxHMZU6sLSbxZvEI6btZcZNrPYYUSOmiRmcgJxWTYsZ3
4CA9uQgAN22HwDWlf5uFX+04AJXRsskrFaEB9+sWNDdzVpsxG+6M33TnrJmz
e1h6Du1nr0vu/3tLSHc2BQRlIDhYQx0H4XPTvPlCjNgsexi2vJ1u5kL/V51K
qp/ByQjkPjkY2103apK2NvpWUkzjMyJ8RKeXqzmJS1e/cArEpDitssSanMDy
jmdUl71DBDMuGLoNxKvWMe9vhYAokihb25izQ8qxFRZ5cpgLVxGAlI4bAoy8
2tmimLu61lRS8Xrv5MOMxORxB9QQxkCfrrWcFABVE/MxMYFos752LEKtJWt7
fEN6lkHSySFfz5pU13cs6kp0VIVpkh1hikeSwr0bkO0fRoZtT28BBYHsIchO
uHXs4V20xJM8b7A1eeOrhIaOsALee2HLakSCFzf4kImpjtwVBTb18xhbI4Jc
gSev+62oGpAVZX3QiS7BAOy2KUWBDyddwgDUESSuNFm3mx/TpOgrdDkvJT6W
NbKHL6wSzVqDyMJnECm4dLRJMm01qufkPLhPeRATxBlY9WZUm/D8q7j41Diq
cRNupYXYmf/t1i3rS1m040i5F0Klwlf8+dcXHJZO39AJrNA6Z8z5+Zlhucu+
GMHhSTz3S57QHD4V7eyJw/RBZ2UrkcCwsMJJYqm0bERQ1rhlgaptXDQFuRJO
WilAAe8f//j7cSZCg16q5N+UkndLSWg5VPZSqusrLji9T0RhaqtHgEDzGYfi
kCMaZiiVyBpwAgFOjiXbiOUQPSJq81SO1XbnFiafJRFL3onvthFxH1lVfnl6
w5aR9gLg5LutIljO6TPROhtGJB7puubiFiHkO9lILpHwItg3dp2EnSEq0KdR
aPQnySp1/uNzERs+7FrZEMKg/oEDEk+7EFCsrvMgz6iCODJssULFNUUjJalj
hqm5xvvyttVYyj4oROUt8Ul7rkJQWiIgmAbH1fULt0xcpzNjQpYbYPJVBX/9
s8g/EgQDE8mWYm4Fy3Jq4BghUA1sdQZok7QDdQAfZWy/v+VyceLwMlP2rhud
D28MZbaBLtlDGOoIw+vttDuF4NViJ9yHCYAXKD6oTj7FXOMaTtzUdRm5vRkR
QPlSfpzkzEI6ws7PNYXDXNrspa2fNlQgjG4ThhGzxzhE4Ow2jjHVh2Kh8GlV
feCHyNwauYnAu/txvpTdDMdS2lexpnPwkYw6pAsRduRImMn+DlMJSHpJCeGc
k+IPyKEVwjj+LQM/qMzIE3+ryj0CU36zwgQ6mq2ralfEcHi6MXEykzLEqYq9
KI911qfzQdGdTSR+mBW8aU+GXTca1l3QDJiCtNR4lXrPaCNGfYtb8YavP62P
OnX2dBoESw6TLZqM2uf4bl+yyQZT3pvxBVfvnM8jhbFcIGfRUAhq4uO5XJg9
CjDpkRkYE+v4kHSMtpNxNudApPCLD2vLX83sTtT+mCA1JDxvq9umcUr/BqOj
Z3bAE0bmigHbUCEUslfglvQ7q5MrCRE5IjsL54+teb5dNZVEI3jYGgNg32kM
mTUjO/ah96TDzxj8PviDDvcjUZco4CG2O4w9pvBDYDEiWXAQasJb78aoBKQW
7fdcWHO7wJi9S10MbkTwiDW6R0bg3Bvy1SiebpH/6Ack59zz2XBqaa0htHni
QZIMrFoSXgL+IBX8yJL8OKb2haGkZa/FZVQ/amC9rfF62yzQiR8Pyo6SdBJO
qS2f9DzZitBmC2ZwupY6i+wwbwh/m/JwtEeCUNbm/P3+6VDwTCVyrmedKd4H
GLLlwg00wwHYY5wh+vH1qRK1WztZx428ANjm5Gkj9ceZ41reDlwWpgw6m7e9
0hKG9jtlcdht2w9aCUvItA78j34gdY2dUpTEluSeSBJUTa4jemltjTUxemkO
GaX7iNjP246suTpQoICBR7gCgc2pnrhQKY8PCg3rfbMsQQGROSlkl/ErnUoY
a6P/VpaDGRFfiQCFAzPE3w36DNevIGEQXdSLNAn/YXAMdtkvnevedZ989h2A
wmtZNhyUsqLswxOTVrH6Cv8A7j0UfHrsr7RVs+7XyHsYSELRGRluvKM8CPmo
qRRcGM5wqe+WOTHvyCkyCrcUGaHA66CET1T6jvkg4L4W3M+OUAy2nkiysTru
McMc3i7HVKECRIvX7vvIkNVNo1kNzJKu8hw72PZmexpZ2gnQhS38Bgr5OP3D
m7SBRELd8TZiuQkkDS4bmDbFSikUAORs8ui17iqy388bixmoJwHmvX1tbJVL
KJATJo0/HS7vqWtfeQWFYU2ToTAxF2kpBvDEC0LxXqFFaD+RstvK8QvTdvjx
wU+gH83J5nSYa5kLOL1dCFNt4ci5OE8Q95et8H4x0UGJXXuB0jpKx0Optq58
vtow77r8fvh1mtnGWk+QzKUSy4dHglndOmj6hr7Tl5GyMheMf1rFWA0nNi2k
OLRXxx41AUCJfRTGZsoMvmeqjvVNIuRu4v2I7iOmtq7M+nPuyIzLtsrkf8yM
PsgWT5mhQbMjAUFCKZbSEGzvahRlULwMYmjqNutpc54H6Ph6nyMBchG0bISQ
khPPtQ36TIJcCNrvZ9zpeVM+lnmDsMV9GHnfF2CkPa/jHHZ34s92AqItXQx/
YdbZZ6Tg5lyTQLR+q2QAhZmM0cx0mYaVbwZE/0EpmsGnHalSkd9PRQcriPH7
Y70Aur1kKHIPdBXQCqOs16UK3MAg+cO0SoBTfEGN+F+nrVKpSZzTyLLGi7uR
NjE01d+b425uHJuz0gOuP3SdyQ9h1mEtgi8bjHXv7gIyGnyywdf8lChTKDBb
mWX6vJE3i8RN9uyHZ+ZoozBjQCkCnAvWaoJhCEXGz/mwD148KDWsp2R88l/T
nD33OFiwt5ApmSwnAnNEc/CfFlg1j7grJyr+yIhup/QwVny3jJjsemxzONmO
BnrTCUUi0pbUHgBvQPmmbPSkbrSn346gG1KSYVlGHfLIlQuUkK5S2YC9X0v7
+M2nABtsu9RSTvAqfx+cESJnyDsNSvNZIWsen6kWqbwDOMZxHsgu+/8Ycl4G
49WfK/4ofcAr7d8DHkZejd4cXFjb1T50mEWECvhMU78jltqMmcmQVMihf0j4
jv5lIUVMak/5p0YD9jqFlGITIVwireJGMt59FwaUMn0BjXCrEz9ch2Mh+xhp
hetuiqLThQO+NMCa83a5Vn6nDCXGW9lt3BnwQV2CqQhasSDG6Ssb6M/2bsfL
RW+6cx9GCBgTOHAeAq02Z8Kv/Ke2UMMpa/rO9SBeqnyb2rQjCxDM/dA1eLlS
VXi2nVlrXjQ3oCzTBGRa8gthAnXal4QgMozABPEjyUDWQuO04ywl6WfivMvr
H6g5gRxm2PX6OwjhdcBEBOnhS6MFPNaF9d9XqGneceXG5Dn06lG+Z9TiVrbW
tgTDXtQ53Q4MjXCvdl1aySMiMzD8RBY9jEjefD2mW0RzKJm1KL4dW6NXZttq
n9iNvfGSs8q9bbQxxTvolmd/m5d9Nqo15z87PaWpy6Jlp8nGqgvsUVEOIrSh
MqCuE8jdOyJRHGSMszH3f8A2QCW/hO64UAwBFQGMqO1VcJqyGqzhAUf0t6Kp
AoGDzvqo19A2UpDXf4sZ7IznASNpymD6cZgcMhINICeiIKFzpLsqRQcVaNI9
V9JUrV1ynQD/7dfHKxe5igE6Sv5wPWJbj0eSh2lR9M3gGJYzm4AFGAHYa8WV
0M8iaPNdWyMoj2rpYzywgxaK1Tfu6zRlANhqiTwPezHJ8HJ6qlGW2T5X0imc
wG6C7Yp2/iJQXU/aQeB3zP0GAmMuPfTn/mGxJgF2ZddXG69fesuK82zMtuKg
Kz4istIFeLQiQanI3bSJjBOKA6Em9wVx7+Sx9/qtVW9gQXoTCfJ3Gwup0A4S
IK76c7bu1VJ2rLcZhZp9i8P4OZlLS/4ppMjiD+Mz5jlVqpro4yMng/R6o5/c
lWt7ZP+yigXT9NIg2K7OGzSL5sgOTXHugnefV/qfyHnHLkW5t9Caetiwf4r+
3lgLdN5bClWkWve2/N3VHBsbBV0nwkuxglTO9VOpx2ra9GZDwF9hlSIM14Cz
+6L8HdSevqoR0ijUipliEejaICCL9LpGvbcOKn+Qd1Owwu8Xm6WsCoLvK9L2
D9mj2O8s5cQlI4FuULpjbSvL95JmK/6THNXNFcQ0Jr6yxcss125db81saQ7b
tFmgeCpk5jLftBI1dYFJVhEvwhXwnd9QBlM7ylsqQUG0jLHWAp3Aom7BkD0A
YO3/C008l78djqtfhXq2JnSFD5gG6qiroRgQB7SlaHzISlY61p7H20lwofWC
hcCwHtVtxnpORMcUjqawbdY1MMcq5M3oU+6FGjUdWXrGT57yKDjzDM26RLw/
hDQ1RI+z94hNFJ9DOjIM7u+ryEgCzFqN4SK1DrUgU7h9hpuBtMD0+ZceFfcr
kDIGYwthDsK1FBNYXqTEIlNZqtbPhO49uakw+bvGRod8tyCkCZ37WNyR4+GP
k1Tx9WY5EJ/CPhte/0eGeEK+YmVGXHtls/caEG/Ao5rpp7C9ae5rWNS0RUNP
sbtdai38KT1D1Y/lJkNCGq85wjrUWCW2B+qJSXdzDw2ppAOm/9YO4JruKt+1
5yd/giLkzCLKgb0qptaPI+qSWu9zWXqCV9OZwrb8P4RXkjmOIdw4cXf95vBv
FoKf4DIE8DOD92UCS+mNNMOwKLqvPIYMaqDg2PYcfCSg1XCaOg0PJq/EWNhM
Tu1G8nc/HQ1egcD6D8EEj5MAdOME7gH3EF9GAyh3KGIc99z1z8skAFzEqkMO
OnKIDl2Oey/Ux/pmUJdPkMplV4ooq+16Sva3thsRMZpdvXxBQiCKIl3Eja13
pxmtGgoxXpEP3JUEuUFzaS6CUTi2SrinZ/1vLEq+vtqNVGRz7l9H7e5ocXHG
DmJPT3Xp/y68YbssIyRaSizaEK739nwH7ak/xiIGaNgZG1O2sy4xJfSFUd/N
XrpGLmfovTOT6YBOp0eY2nl3LQ+f05QhNctxb6pGwEhcyZQguR2xqj7lZRnR
nZgXpo6LoGHeX80oWNCJvGVpbwtkWFU0a89J5092NNyRsmiJYeITONEflS4R
V9ko1cpluJGmLLWxIpETs/Cv9NinDjp73Gp7GjKETotGJf3AgQYoQak284Fi
DBxIY/HWDkU+Y/DdQ+EfNoW6HaGpHukpwW0EvUToJhPNnJLMikikkRiczPy7
aZCRQz0ORB/uF5ISQhLnKCfmwR6Qu+A6PqDgHxBLY1Mcmon9PAph0K/myWSQ
EiDwtS+Rj/gvt77KvlMwc2j98T7oMzUqPRY9kzsO4ppa65npO/L5wOfEo62D
f70SJL+KxRfqv7Sdq/f6IKrlEiu1fz1BcvJSdvs0I8qYDffckbZyDDKRPY/3
9XwK9gp8XOV8IuICNbNUuSkTX715HrjJmqBGLaUGDscqR84Y34SxFrUigyGP
+8QM68aBzg/tcMFNGjZw9AidpJd7Gtx0atL9pc2471SNyhGkz7sw2uUirP/w
+bygtDnOt0RaAebzx5iLkaXZz1uaYJs8mJPVrxVI2vflBTsNjadJ6dNH7Bop
vNzHW1ekPnk+s2ct5oUc2eaH6Oe+WY2LwhAvXFcBb0hWs+ojz6uj6aP7AOUx
hXHURWnBf9BOcFhI2/o5WxdFvt+n8weQOV++97wnF9WTZIVUawatyLuo80oM
aRGVkMgQ4EYvdz8YdbYR4YORSdFKLh7Vaq6pFuejaHewhWb68kturZpJV4wP
UtqRVEKg7HHhsivhpxC+XDoU3e9QpO/fuTyVLxN9T+Bqe2+/iGZG557Deack
HN/z1nk6NLDcdPFjl8o4hf/7MqIaSVLF5lumTIZXnfFTxm0S6tcmhZYo5ejx
UnwKosxPKN4sgl5kINmbT65DVQBVfuczivUh+p6rYb8vXS4u3HWyXTxu2iHy
GX882V1SweK0XGeCqtGy6MQdVGyb8hnEt8PyJ5los1NkXm7YSuIduJ6L59AC
Dyd0b+OLzi1uDUSu01kaG3gT3iapyxseSZEwDOgSeM+GftdfZ2f3g3h3Iw7G
BYDw2OAkoowh2E8urh/Rob1SMpngtdH+Pg5+1/DRbPLvowKzxJi7TwF3aAve
sCpmJMNQVJkgi8d8EyYv8TDJTqh100rAkTpDvRSgRbhEQiY1kG7kHhw/9DIc
UnkSPxazcmEsrpGHzPVTj4F/VAW3BEphmPNnT0s19bXHnMNp/QIMwr59bVil
cDJW+llDMIhC8mfUJLZzBFvQS5CxIxiyXNZP987JluG4aXlzoFeMzNX9sGGv
KhrCXBlyU0mWGpInE6VvJ+thT4yg4BOhx8AbBs6PzLXzgGFUDXEiJ6SwZVZN
pOUGMQ32jQ26U43J7Y0c1IA8+7L2LXdEyMmnltw/Vp5/iDtWj2Ls1LPvNfLl
i9K30ZHTQ4TTpH4XQxWQGnrhOQcvuzDzeZACuBmYw+o5N6OEeYwBFZY1SHxZ
xY5GJjUPI81M4sezoySgzmVZJ3o/8wsO0P7vrJQofGsU7hOmKvAOfNtGKdPq
ZNfr6E6ZDhzz+uk6AVgSpNDwWdebCOcwAU7EyZjJT7K4OOJODrRNy1FkFZFW
x/01TbnvLb4govBx4HSYNEh0sVIX4Hysr4rw9NVc+s2Ua3MPEgxktTdLNjcr
TFI/d2FL/KdcvahzadcQgDLChZY6kq3QoUnVTdjo7i37kG3wqV9KHh2qVKAB
pSMyVJSDZDrOpB+M56qYHAeed7/F2UC5oV/2qz9seXFFHh8bwhaiZXl+psBe
/pz3gBu5mrtQkQD29km9C0CzhUAMLcSVcg0n9A4EIy5aFr+yko3sKsnSPGyn
Ie6XCKL9w0+RnJWM7iRWF5yHwHpUIwDh/6/htbFNxcrWFIQ2xLuWNce3pHuX
M8ZKpRD5WW4Le8uN+J8f0htPGxazj35saPEZvldOsbi9164Y7d8sXNKAv8wK
hUFP3XKgVAjxzaDRXOFWyCGvvKcYogHnBqQFGwYQnUaCOu/NzEeYKvo00pxv
euxGcMA29Xp9ljkDcRw+JTpg86dtXk0c8xbjoZ5EnKRDGzNYAd66fm3XqB6z
Ugf77ltunrDUvVEeZW2tlUs/6agqyOmRN471X5Ax3efcop97zf8CnyjJ4F38
Snqc8FWl8y1rWE5lpCmxkWidfj2lBl2oCmYqQr92W34qjUVus2Y8umQwyOgo
zOvYgzP6eJIMSTebUM5bJYig6avD7MOfCQfsSqPbjPJbHaiFsKaC6ORGgIbR
eTEaN8F9dz3xeTq+xsBFHWjHFOumDGd/7cty6Dvf/OpRhKlN3L+MwaZO+Uv3
TIFrYOGScsZ95cmnNNOiAzHG8hHt5xKO5bJKT+6uOxUCNvkp7ySKyiITuuOP
5ufG8xdlm7rw5gB5dy7g9KFWRYR13KhpR7RNs5DDU4XaKs7F7CnhkqoJW4Rm
VBEoIW8/uUPWQI5cgpSsG99YGSwKIHsDl6zVbVmfXsKtxc2RfAJ1lFrsakSk
LQ70rqd56fyckn2ji4HCB1YjYTLPe8II4bVJcmrq8agmwjS23ceGFRlrCt0v
D2Ww5OLrMpBa5dpoTv9Wxko+XzTcKAVLSVBN5p7CE1iMGWVZaj8Kg0LRScL3
X/Ng1GnG//jI/92LMXLDtb/d1cP5zFqj9IbpD7AxSCpWkEpX4K5/dlX2UXvP
3zkPyxu2cQAaqxN8S4EASDBZWenhgjuqoJj4h2CT06uddW8wPD0/6S1C4UFL
YV7IEerVXW1UEkPCcTNlCpXuQ1xNNNviFCYwxugTCfuSPzRXYQg3O+XkztEk
hisVK0TPnGaxY45gt++RQoy21Y7vl6dK4bQRGUhCK+ul+vomfEBp8uRIwAuH
5pqOPdm/Rys9mEdqZ+4IT0tH4iTEvrN9+6f9b9RYYWiQm7M4LR69BtzJQ36m
8oqMWBC/Lua7u6AAvceoADMYxzczcHBofyP9ILPG9vWWnqdPW2OnoTZmtPD4
tUZ21Lypbin4Z/FWi2KusupqYNW+Xx0CRpOkXTDfVMw/3iSDR5CatLCZEIAT
xEFn1LzSbxj9G9FsyDtLcijzdqA4dXhAz6kpPDHcnF/bf1t5iWZMrTTUCSl+
MCE8WaCjkJ70z9DfiLFM058e1XJTdGImctWehF/ga4A4DcK/s60q8wy9c1wG
jpqN8EY7N9W7a8aPl3Y5r2pXgIcEghKJ8+ceix3A/cQTt5JT2ne1dEIdhVt6
X+9v2gadHXpVZzU8GTGlKO0VN9wMS3U8MdR/JPze9Aq5dytILIMXpfIftRGx
IoQPqfZroLnTxcDg2f+nbGmbcnpEx04euel0SkeKu82adm3ptOCqeKSz6sVF
qRBWGjEJrXf+E/ZNk5+CAh5rYb6C+TK+bjBpwfqAXhyl7iBM1jrS9aua2GI+
X0edVrrE+iM85C2MNOwhUI53xjo8x6rE51btQgsOBupGNuOHTjX8wyLfphHs
f1KqeymqgJxBclErTj2IHzBNJjDNRKZNg79geTDmTsXixskzNYBpMMG3trxI
WN8KBePEOBcoFOhQMR3chy/aGnxk9fXLUGvGnllmdceRZ5ZbovmeQtF4hzaz
e30nn0nWPDgYW3Ajez8o4NZlyOOKarDRJbowyCG5A1d6H4E62k89u0WgwfE+
5Sn4HVPQYj+rngUOFmt06Ep6J/Tz6szKsQcjHOGtcvQSqfGdWQy/qFeWuiwi
5Gb3rUvFRfO5TbBLsqmNOYDzsMn6oAaaDsOqZLdaIA426g626j7831l1S/e1
XiIBHN4rMsty37LlpRFZx0EyQlOm07/3WKbdP3ad+hw/UnDt9OReDCgmduGn
90SowQ2rAeTfrUzq6kG4t+FJhX0XqB8U/IO8yeGz2dBMvSyBlJuqP2/xJNXG
/Gczj7ylv2/CBBnd2e6xYGDhGfREv/WYwZvg6O+smAA+I1VbDlo+YE/yz35f
OpvuMCH1wuBkTcyxjvmxxfBwWiAekiMkgACEH1d8dEruc7wjxNopbIJrwspv
3Q1Xf+i+/Q8x1MCAKlaTBEK40LiMdh7+hcXhhZepmr1gm5kOz6WZMKUQtyOW
b6M/+62m17qDgN1NtqZk5pL2nMD/VpaTBF9SgVDRLvRdcFy1KTphAjRiB74g
kQ7iTFDCu0LhUrlQHMSzgXo8+EpT+sRvzWW7bXZxQ3XuUdL/JPz+SYvhI28d
KPj3I2/ArJsRGEqDZ8mh+vh1R5/fv/4K4h0bKtflcB4NZzuUZFqhp+7IPVjE
c6ZLQPq7A+6HzysAmyPhYwjklr4FFpxTto9QkAVAIJ7/r/HqDZ878OF9hEeT
bPJq8T/iIPGtxgzwpi1WAj21IXSOaF6G8JGuLwbyxXAMeF/2lCY2hIsVfdgz
LqywT3mtgOzKcWKeXts4dB+Lj6xqWanjALpXbYu1ZRAEQg8EzakNuamM4RRa
D8GMkalthwTeaKUk4S2I3+uI10xTOgW75j20Zissf9coVVHEuFgH3R99xnbD
50MJBxo2FGAaHo78X/whHvlEp17uK9dicNa1QbkfBRZ5POCvdoeiMiSF6vt3
Z78WVEoRWNCr1WdzkDe2Nm+xdp47lQcPx+TljCU3mHqhqSz0ldbeOZdWzUV3
+G9dFCNThLj4KOsiTVV5r2mjVP6/SWCKFa75K3fkWLNjuwGbpHZIiJAs9toR
gq8+qSlgIL25EdQ2a8PLlLfoUo/lWvXz7SwMARxvEN8gsP0EGKs0A53wnbwe
oeXXb0l8onNko3vPVWSzRSl6ARtBbrhwMq6m9WVV+q8uy/F9M2bI7X6IvkuQ
lTLyEi/KmJA56++wfzLMNDRLBAGEwdd+4+Br0Dar8cE8z8Av510TdWXf4Hqs
Wjx8rWr1uAW9anoFu1VAxn86UsQFH8r/SJsSVdfWo56yr3vjhy9Yk+GakDRO
H6539Ip/PSxa7rWh384/CJI81LHdJcPeI8P69cF3R74+LRTDbLUhKqgOf/e/
yQIrGcGyDt/04uYhrzk6SvZO5/+NqwtA3n0uKjjYFcBCNwWbMVWdV6YhqXrK
PjQgJadGPLIMDj4ecmSCcn+U19pvq37QiEFWieWmu3I7juwF44OAIZTBktLA
/mxndmQ8ZdOmxqOy+GY48rwShCa7ciFLtXwruCull0L5hxygBY+EvVzeyhbX
OACJmM2sGiVPJ6zuBdA2Zk/Q6TYiaUPHqvOXF4Xe3r1XiMN7MKrIwAWYzL3S
nVDKKKRleox6fcg3zlTZzhEopzJ1q9oJp4AsLZ3OtpWWakvy3Xwm8vri8Uz4
lPXwoVwbCIilGBuCTlt7VOTggdhahjk61x036WJ6zUBqEywL6EYIpXW2VNGw
3p0t7HLbjkX2g3jFhbS22KXuQys/v4w9e7l+WTLrtwVYaNKAJKIGBRxEA+xi
hmdeELkYqqwMpBU3KdGOF+QNlHAMh1rtHlMutP+53Th8mDpcyqL7VJHK0apD
D3o8zGojalvyrzYbqXUV42uQw5LkQswPdRFHAogd25cpoektEl555h0Aouxp
RsysjvGjRgq4Z8At4ugCqeLQxDTyt1toTBi+zjCc/aZQvFEi/h0AOdYUg+Q/
aU1DK5mMINkPy48ULJZUwadmwUhAggZtNKdZJlSYnZce6kwiSuFew2FvU3WM
7s3I5/Wm8lOWMofdFxU057rJ2qYsX0l9DPuvlDk9cmy9a61K0UyHyhb94ULo
NzVVLsXQLxbbXBcRYms+V4+CZxKncNVITx+yRwBRAa6dcC11WVxB+vMiRHdf
NivvuXSGP113gvVPTDKEj5eMS8Og/G31MW7TfEjNYwOWjQgkqbUmFLw0DmeH
+CgQE3ASLw0TG+Df5Z1iNYtDyF1/SLIk2eRvmneRQKWLfTCLPWnQJfAdMnas
KUttU11RVN+Yxu9RySUGHgmlDV0goEeYSF+qOSJEzGkKte2EtQCKcA6OlBJw
9Aj/rpH/wsFqOEIX74I3ymziVNId8+X454uHYXtv481Z6COJaxyoCcA9lbD7
v2taWRVrUaVgh6DWd90Rofizu1HkPjxpJfYHLKf7BtuWjMLTSI31v9GXUcn9
qH9ojw7ZF4XOFTFWqNueq2GztCOejqnOtWQqkijmGK4nZBPXm447NxOrHlB9
4kqHSsUsl+xMHoYNbTrxzf8BSQJWKt6gLmx8DUZhXAR/1KLFJInrKvI2qUm6
h9F1t2+TLWcG9iW6Yq1dh8Lyc1lE5ZDLnyJCsqbYAsNlxaeAfPkpBiFo2Dm5
eubWA6lHebL/Yi0mR+R3ddf78J1XBUvnqzEvGQQVnezUeH4XgUgaBLJzZoSq
R78WLOm3xzOjWdgl5ynWaId8bcLEZcOHq2GBUkfBFOc9wBHIdfbXNSEbCGyg
tLgxtx4xbcvsnjArOXneY6UpQSiAB8oqGjhexGVcQAu/RL8UyCRVSwBbzeQc
z0HHSghZyorLhTlHz1rL99j7Ts20jQwxWWMBxg8mT2QtwFKm0xPMBrU3Z6L2
9W5i8yWLFdPiunhRYlqVJafDmi+6Rwdn/eoc8f7C2bVegXS//XBHu9X0Nrr7
D+D2s0JLVdjrQjmG2+u+izuUPJabYrBsKTb+i3bUwgF2BXwCFEudAfFHTZl/
U9HvPd/vF6K1j5h9/pqSbbt7ZiXMvB6diQC1cfTVPsGaKTn6Fa17W2Xry17k
Om2j8dgw4oIk/HyvR4QxEl2HDb4wmOJm8K9eBH4G53lJ9gqXMXDexWKogv7k
6R0V1vt4x4KhZ2K6KnnfsqJUQLE9YsGurxBZ99CCBx/hI9+vSE6Epz6VVpMw
M57QXl887PQpSfiGCcfBvMqPMDKj+g+C/c+GNK31XaR/IM/AMonb1eDQp4zc
/CObHCbXHNZ0AaWEBq8Yu0W6/VK8Bl5Ic6A+CDLeiZWQcVVasSE1ixaPQL1t
U29Ts8ZaOxnvuo7eJ692KBicXmTRgydhTPTQ8Frn/u6QVEq+X5Baz8TUDoot
XelN2jebFaH1haw0iHlQ6PP1ThVAh54oGkLXWcLTzB8XtK+VU70v9gjp7nDH
RYcoH8frQhVZmTwnN5/qKMWi/VeIhz5OTl9S6lfN/2ssK0O6MW45jnsiqDhb
vYjvMEWGGBrhlziKDA6rr6acYSLfEW7h/xaTHp4P/YurYSESWeIarK+5nVzt
DjbyQP09zSV5EsM9l1jsnOOcEFNN5L5o001PrcEl06G2cE3z46gZx0wz+R4k
knYNAHZnom6ypGwuyOeSMp+T/VqHUhMzTsO7pXtuR/RJsa//88yEfStDUGBE
4qi9VbMFjaOE3ISgZRBqNBbBBsi9AtlAvi9LtosVHYddKRRJ8lhxhNCfNz8M
qCszT+ArweOrUvEHzbfgQHUKvSGW2zLinAXLJ0FK9Ks9sxMEoS+Fmfc4Qp7K
5GKh2ADMit/Xlr2IpKeS5R8yfg7NNOPREuZZbNr1VfNasiz1yEWKfDhPTw5n
CxSr9Qps+Soms8aWoXwwNWLcYnieCZ/lip9/qYtUR9J0366E623bRiXNU5h2
Ao5A25rrqByg9RMTxwhU28ujpEQ1yfntIzJUKSNysSXev86RiYymfGdTP08D
uXV41XHb+lL3tvnSdwzFiscdcQQNAMyz71EKq/uFbDMh/bFE7VouQKq2POqI
BtakGFPATHzDeEfZqIAh8D5pAWIcwrsl49xf/opEoDZuB96v4IGmtACqclk6
D8ZvBx0HmODRF6yDhztJXWECxxFhk82FTBZA2fhcKu+LbEw2W+rjF3WZWXKf
LrhyRzcVJUMuLNuGxXRU4+cdiGay4ZEZO4UiUVqJTFwLtXXwQilop1derPA1
NurrAd+qC3iU9OZZcoYx7CqVxDkuF1hbvpkIVMKPZIbA+EiODXhmx1aaJlkP
zDIttOnfFikOYL1lzGU1HazXUBMyery5DxHMJi4j5p1x++0VaxZQkWPlZytD
eOSDfYdMX0LbVGsEEBO5c7wA6dxdZPvIzH4HWjY12w/UD5MnLq0Exa8D5rbf
fC08UPcfxE6ilZA9142Qjmr8VqJQEkVi5z4+6n9XXqDY+iVsQWU2lqtNAhr4
fByUK7dxTbaELslUNs02j3l796baUYkVXu48SzqMbmJ/tWtNmPfrubttGpQS
6rf4w7A/LNrtfRYxvoiz/A65lXmytHEnmo7FpHy9lmVbdJ+AlXpK4zjCpF9v
DbwA73gqyyvA3v81IbiRhLMAY56wKzgIZ+XX84AQYhvyAdpFTk1cuQYln1+r
TueI51/Wb4CrWODigNZWH0V/yrAGoDYXhUlhJMRRTjgysOYwrhaRBPQXBoCF
9SbBVf0giEG2yIDodfNo7ZjSNgqDc77MJSyv89Zpe6kAQZlT4SkoUz91OE4O
p7l9H0RP+If6cXD62yL481RoAIp2/6McYFUDPT5r5RImNThxQIZcBwVGVMar
eQt/p/UEEBddyQwkI1X+Q4m5YZ8SN73wPpTr54U1zep9aMavw3lPAb+Ug7et
YSDDf9IzDNzG1HdrKNgIq3fw/u4CCRC92f10gKxif9X+05gX9ZOv+Dv6xha+
6WKqfPfkHbhH12eCNj2f5USClrSMQi4SmK0GWl1CtEmZYuA4Lo3MGgduHUqF
SZGpFjNnhs5lEvYFrIY+rQ7p7eUB1s6oWe+I43aBfWW5uyxtwrImTx+rCwI4
i/SPJqxP4M8+9CInrJPX1OQGX+P9J9Gq9Vc898ZSZ1vRTJXsarQVoJ28r6yf
i6XKvdSP5DYxv1ZSs6Rd39rz6ck1KV+RjYclXkd6/TyzyhmgRRBTlMeyB1BE
IrFNTgir30BVnangLk6JnFfL91DTvHxbNY/hu1lSvxUiZMw35qEST51ks6qr
8CLLkA8nkvK76vBPi16GIeL/2ImDFdjSKaGQfHUh2owJcD1mAdMk1ZlMHqo3
3LQo1S8bzKgOJgOjFG5Xk9m6ug7jSVE++HDBj/mkyzsoOkwL40hkEcnjYcxe
l4OtHwkbyx1hvQxl7RVZqXM9EumtrKrKPyRAV89EcjM2PEHo2hmmNb+ustky
YsNXtiU1pfiMNmrs7V8rx/LpvhdLinM6MChTIKbsTLoDIwq+2ShP0mS6g/4F
1UHoY7aBUysIBuhDbYAgSRfIEJTsSPry5n0QdlEoCKImR1sodiPaXFLxQlOr
vD1ExE1Q/RF/Aw+sveoP4QB4ea9y6M0GgiGR/wzNFlDa8xrWo4kva6LrQzll
tNZbTLjgubZHP11cG5KTr5fsovkOtNLUTo1uG4RRMdhQ8acivyHYLWgwhsI9
xanECrzns6vSpJEk7WUReusSB3QJ1JSOtMCf6br5iFEt8MHtT8G1Y0xsP/jg
zcuasBBtb/y7TM9NsKNmhK+o9VT7QibyhqpPje32LHpe+nLefm3KYU5lbCOD
0Lp1FzHKtIotuoA5pJcmFI538FUw1HxGB0uyb9JLKhC63Tc1I1NhITFvQzed
3XLkp/UoQQ+Kn6WmqwS7ImIfJr6lcEheGSl8kK8JMHLLTwxd0tiOg1qtuxJE
OsGnDJrswbUytJSjwJhZ+w2ofHF9pVijt8Tltuf8y+adkHsuuMiQKffPp9ZL
688zc0yArOn9LfkbgrilBZm4IHwgEqlCuWTfPzQwYAlR+V2IgrcGUu8odQge
AHHnFM4/3HPr7Elav85C0asOAYUi/KVG8+zRO6RUd6gZT7hbuzx1Tw+eYAtN
Fg0sfcByUikNtnTg0YHGF/k4Rvpg+T4C0xuzmMedr1mLB3iAPlSl/+quaNbl
CqnfTipTHFgI2pcge8iHRLAsdDk6Lkfd+DfBdYsA8ZLqbLwJQ09LUoRJa4Ok
eAUvUSPD/bizfwhfkIzrWG9roaglcM3uPO/4B4E+TXouz9siNIE2bW+1ec8Z
KN9sEBN6200wiYnh881vZw93U5QMU385t4xgtt1gtN1MiRsozEIEQ5zamgFx
HoeBxfsdnuhyt6mHY3MQ/XT9LWdoO6rj8zEFbcFYIda2t6Lfy6w38FjSN51v
hRqWTrFQ8QtIj6AxbDbmyUlkUfacMeP0nNoonEh0YTXWGph06BbklUd7G2YT
Gdwk+3zOlgNC0EqQH+LeUkvqgUd6IhqG7sTqhD5V5PlCRjdDqjRJRqE/deN/
8WoFYQbJ8/x80jiXu9t5FbrxQFGdq2E8zJzKGjV1RrViPremszhS6ZD3iZwh
KhRHBl5+dZkQqpMPrX+jhL9dFrFdEL3IIkWR2LWXO9lnCCozGDxO3owu/Ha8
AIpGuYhjCflKOpUlGsZh/OJiB2vzr6zxjmKWRJsyYWkjNm/ic2t5/U/MDtOl
L3P3/2FnNa29kgeWJD2pi8elp5MA8TKVam9O1aZIbPBNvOMxl0PY1Zrnrp4w
qowEgND+FH3DocMdb/yPKDLMKQdaCNmd1PlCdY6kxXMs/3TBILO3lHMj9VyR
yqZQgr/ltKHMjY2LoJC4EydQjSPBa3nPBGaaDem6HZXwZiRd1nbXNul3CYDd
CankC7RUry8HrojM83LCcndCLJIN6sm6NrdAPLjfZ3EqtnAghJeG9MazDyv7
xz/StsNmsaQvR+v4ZsMTC/pCH3maMMH62HTHFgtbQrsiZtfB4LeHfGKKZvMY
pfb3pBXnSIBSYSRqphre7K2GAXnZiQMuLe32Bhaqwedk7lIxk+pa+x4jGvVp
/IPaWSIQE5+NOIHMR47Dq36TA5/BMWPIFk/AHqnLJjEfO+zqpC2QdH+m77EU
OfsvlvryodEGfhVDEswJ9086Rse48W/4vHCLtPs4pi4t9vjaI9A2DnFKjOEx
fbpkqkrKfJ8YEKUvE+ZGKxt3itg3rNNYokCLSJcIM1y4elnp/hbaz3tIMljU
/tJ6f9thZl79vbdnCJELmIH1fiFlVj+sbCX/77VpAVPmSu7h53M/uGqO7YXJ
fhs0PQyEtKLF5nAYeK2mtpMYLNJcwKsFF5577hbi5m+rL/a+EQrRtwE7IrJf
Cwz9l4aIdWt3hZ0fVW/BaJCKPhyhZbXPw13Mgb4d9/Nv+TO9oT6ixIZuu5b6
+fRhv6r6WkjNsjHkrjF1Hr472IKJF7ahXgyH1aVgL4P8eLAbHdN9GQr6Sf1w
fFg1E2V0zqxoWxzOXPWZQn+y6n0YcchljV7kFEs31SKdj37LpTGJEfh4fO2J
kkrc3+0LcDPcrnDkvQ04IbCbohjcok611AmX95AgoMRwoWfb4VSO07ZeFVG8
ydRjftir32nAi8C35E8BxXqnsC2fzGgXQ3XVRXhVIvhe6nY27fiU5BSY+ymJ
7dQSl+m0kM7EfKBtG4eqWI5ciiEXgCv2eumxC+VqNd0XxE2YCvjnp4Y04zRp
ERJQE/OBR/pTCb3WqdJhZ0eZKj5UhsciSvPc4Yf/90974oRc4hynlYhGUxWl
qnHQq+iKv0TqTQ2DKQcVjyjPR0jCvXMA0Gckl4njn15fcYe5ov92/1znXEGa
efuQXoBLX1UII12PzzbV/8kHqeQRxcbM4YyZE4G+leAdxgIHgxUjziq4bDw4
0VgrWA4Olyf4w6RKiNoJXkUWfqul2MxUpugii/XJS9AJ47M0SKUfKmq10tqm
WVJJ+1DWUMmxkIjFIdB0SxQ24NALO/+vi0IVY6LiMth72NmGwtAvKCAM5OTA
okPj0FKTe/BLcCbYaKj8/HOBK2LwEvP9/FM3WjEWmiDMimYQ2iHWImwRQzAB
JQNYq057Cp4ITgwKvMtDofSREf0SuIgmnpITnr/w6KRFyZaTIwSkNbJXkUQe
BxpkNxrA4RG0yHPPHtqjsa8fJCWOM+u7sHKr8Ao/YBa6COaAzu2fLV/96BbV
/un6hotuzn04mJLeCO6Ua+A+N9oVY3j4qqjacD8OMnRUhOx7umWjtVXxCv5m
tojHm+76q94TEiA31Q/FxwlnzD3evnHlYKOsI91Q7xP4rd9F7m3hTQH2q6Uw
CARvXJpiNGic/QT9RIRTYoy2tBh5i8N4KCaU6K8StVnd5ASdJ4aCTeg9FHY8
LTOfPkeMY3ZxrT3OvlG6w+DfY7d1l3a/BatcK0Wbjlq7VDm9eBtdkTc8/+6b
tJhQx8nx/IIPZIMgzzRqy0m49N/XsTKIebO9uJEfvPtCTIiw36cASXikzndr
q8WA9HjDrvxmv9SdNxmwXgYEGfmZ4mvSAfpvtEHQwYrfOrwjVkJysV7cmms4
yB2r3pVlMx5P27SU7SLjewmcXpOfpbXoEAXfx5D35iAkb6eW70TqIu/kDXUK
O383kzR6opSIRSDyeogFRqvNTlITRuDRBPxJaZw2Ny0QgD9HdPRhwE7tdt7B
5euHBReVzXhErkIsIQvRt6LkgFJwggZG3BKVzYBA5ergO/jSZ97ORz4WMSE9
7YAkuTrpj2pJ6WlGwb+sDRWzRLIicw/X18Dk4jZxi+y0GiOzYke6EuLYelUk
RiD0nVPQbu/xCpR2m018xjePr36k3iWPtviO4L63h5psPpfnpkPmLRGrrpcF
+sAFqoDyEIIxDMpx0fRtZCBK3hM7R1MR/EQQBY8zQgkab/cQy64kCRtjDx9h
/YUsc2XBPufzdXHmoDgp7bOr3UF6qKxFHKcKIkN01A3ddM0SuJH6rybBDWT+
TLvpHB9z1XewM/9+fEnqlnG7RP9VNBKZ1Rn3rPzxBHBqCgZQ6HmBtuS2VJsA
ItbDhKzfDSQaGg9dxzcD/VfKVXUNEZQdWMndakR0hjzUTuW9cckAJLcswY3K
6+GXHJ3VrqLPjEG27h+QaUSoXdM7iyKOJoocaJsuZQ4bL0eqesAEkWnxb3tg
w+ijhTw/Ir9bGemOD5wSnCty0RJSndV5+NjvxgNB6YfhyvSxxWkYTWN+s06i
qsQdGR5GyHM2JZ7/WZBnSr2lJqirebHhm/jTdoG62soydjcHQZn+vSC9+idP
391DoPpwJpBAehokhqp5q2n9SXtigp5QwfIuih81fqi9n9dzuEC341rs6+0m
AlmJKAx3tvLNXHn0F+BMdu2IuzwN91PKvEgrF//TVvEY59IqOs1VUJj88LQY
863nnF0Zrm6WdJ3W+RFzi0lsHaDpEgFJRd/qHiAd+e4sZQkGam+3SQUkGej0
cAb0EqdELIRHRbGPoToCJv07meq4v1+CVTZJkmlxMyJjfXIxmLsImacONZ60
hw3IoHtb7gy8ek6NKTVVnsAqPt+MupdIUvJasYsZ0DyU14fYnfQZDtDoKPKm
LnqiV4Z50fdJ45nDHr6X2rS6iPwtvVqp8sPH9n1IqrYVdFWLyEZiTAS+zhyG
g58O8FInqwFopDjav0ngezNeOQMCr6ud9FG+gO/qNsmRXGvmyvJtdjYI9YHf
zlWEiFhOo4wTemc0XNqNf8Y9Sb/v0l+BIfEkDvvjIF18GnufNmhKtUWr8PYs
ioy880bcM0dcem+2W+mG2e58gcLz8ah4iQ9AIIfBI8wHZgkB6SEBJlwjEwQV
KzscF3GZkUMErp3gqvoal270wvHgT7d9X0dSCgNPfkX3o+pTFH6e1z4Rn70e
dZ3uegufX7Y3HXELXzUSYz2DLReEXfBBA9c+GW16fpFXhX9zYevRNg43QWs+
Nd7OzsXKKlhvaV+xM8KNU5Ru1qbfwjTf2xgStGLX6+rNU9QqTUC5L5Y1Niay
qxYnZngIiEenUST58OuPA/xqVoPLqAwyvZDpwGAOdJaqVOsn/LB+8k7dXduC
6E15goPPdjDfrWHl4r0ClxUDf747ghwIF0ukc6IKlOKCn49J/iGbI8T14VnL
y+O2JU4C4/n2XsshOuSnxu8L+RD1SzGzNG5LyHkUqBgRxBTZ1euGGxaPLgAN
LEU7MYf5Wj4MfLt3mcc4qHzN10T0DhdcPXzT1EYahexC9inw75DL0D/p+8DP
2tm6qAOBJtFvy0s6qTVpggdOvKmxSmA1O+82mUWES8AnHd9jnqqtmkmWEsmQ
2FhMwKaomICuYX5YhPEBNEEeP/cnotG7gI6hLSXvWDyZIpd/+V13USiDj8g3
9ZugAfYkyyz5eCV0w9H+uaT6gqLTwMbIAdfCcxRlVufchcUnWACU2qzLI9CP
0aSFCLBji9XKo+re//XhmKDc2bqP3XmDSBv+jes9BE3ru5GPhcBlsTUXjbXz
2sOIjG6vk7VhSXk9U04RgWB+ZlZRp9HR6iXDxZNKJccyBejtJ1nbHbPFX10z
05ShhvS5+zwtk28kLQNLzgwRMnbBsm7VXHWnr1OraVFiIazoS9EnjPC9HoqD
iZ2QS/bdTAnZxVQFcg7s+8RpphkMBomqynsYyen2qeoc1xIRE8B4YC1oFXZU
uj5PbTq7pK1YZnMpAMtpWGglql6Z07EHwb22IcajGleOGFKruWSXuohnB38S
+pzHgMieNCTU9p0Fu6UfClnCRE/0rKhG9jJFneKPNdcD+P0bdOb+sXttEoBq
Ouvc7p8+B91YBfq/kPMmxLK2b6aymnD7+6PybMbCNC+uyErFf5dkqM+8rEht
AbpuQ2OJgnRMJ/y6GC/JluWnl1XA+ddvQyjToAWn7I0e13yuH01eqQPI7NXL
8AlpQRGmi0Foni1jP/ijNwmqbwYjcEbeYdMIw2pPcDFjo7I1/nm4NFkgVjwp
5tRvATFjlOgyQaFQm87mVMOQQKl8BJCbbkQW4yjari3H+XmNaB5iXQhziI18
LyuKF5T8lfZ/2bKhvRd3XEVv/C3iJe/ALpbriRpEN+X6kF3LI8Ulfhhwi/ro
HvVGBFOWyYI3jG+o2VimeXrJpxYNdyQz1tUbHlG4KLVUmhGskqgYzH2FUpGt
zEHDYsJxSNZaZUDsmiPDSClplBIInrvigkm9pavhLeQWJnx6iG1xtBublQdg
rWBzL6s+AO0mGvLz/5MxsYSjaddm3F1wOts5kkoNR+i6C/q4EzQiRMQh6YJO
kfQrfPLpchjU3hGRTp+XrDUT5wfk2omqrx9W0j8zST90e9WrJ6wsiBPEre05
W4PAIXglNzUFHbUqB2g86LFr9s578Y3pAw6wImaWp5bU3HTIaC/n7S339FKh
lHTQGrpR6LcsvoUSHqkjuC+PXkP93xi90Lxrrzv56FzQwlDyEuN0dC4EMTsz
OuEoO3oji8TCpmlFlGJiJ5DOUm9bGK80iIPGj/uaOxV0zinYeN/bIHKNwYFm
+PZXVp6HDdT/VD3zncgjnTbs9kJbdQWIb9TF3aVnxkYob9R0R9hjQSisu7IE
HvWsYZpq3x4c7qv7IapLv7BxCloddtxmEj6G7TvpmOYy5nW7PPutCePrj26B
mdo5S+dzCT8cvBg184WaJWKwrYIoQ7Wmq26TrVlXdyzGwJi679EMF3Jmcwrv
jURA+iUiz+7QVFuW4jv8fC7M0D2OqEmQTwkMkfCk+ruqbYOE+VVzx7wa3upM
idEJtb9VvXYl1JLGLUmOlXqakBsK8lTANA9836M11sVpxM2YZ6rLjSzp3Dve
BcQPlOb5rBaiXVjt4TBz+XgyI33Hz93R3EEcuMgdiMNm7Oggw3odYb7820Na
YTPZyPf//fi/9TqNPMUvKYsbbSbJ1V3LFkK6TsrxN7yF2z3LlldGvzFIFet5
RbjKaOVRLKe5SDt5ADoMotUKMRe9JgXAhO8zIGxYnGhHgQoBFLyhNrKdqse8
T61XtrJLadtiFxbivUQxvcfJl/XK955EPELQ8t0vkFMOQBXlRQnaDodZ2f8O
DVGw0ZvIcRXKrRN473ozLeWhgbBX3cxiamEct0H2Kt2g8I/FV7d+L9kmzZTK
fVIO1KDvnkN3/UqsbSpfeaxPjezlI6COGsVAux/CqGIU+5oWWpSlXHzQ4IBD
l3JzW1KMUakoZfSXItk2ubTdca36WuwQx6DG3ntEPNoC8UfvAGWUKi63eVDs
cheqIZIfC0pfXELjHzc7+MusNkIKgw8PHnLOj0hM5z29t1c+DOHx3IUYS80F
yXlK6RjQJeOGuZVjYwjFlhkAKaKTk8JJ4zlzLlIxk8Nk3IWIj5jHT6qnLW7r
cadLjTNrBtG7GhkfyuNFwB3xuFE48wH6yX1OEHQZwkoqAHXtnzaVHe3EoZVy
7Z5FuAfjtvwmFnqxmrCnwNiWRQM/7mfYKtUTnuVehqc60Ht2fW/Rn1Ah1dD1
CvHEh/eNJqGhTv1Xx02GpOeJ2+15FlJHG38h3iCSswHfTJGd0dieDaDAITBZ
wCIpwPj8G2AlxUGRJwwLS3UzORJBKl7lcuqYmMS0Jh0jpXiuz9QOc7NOa289
mZKpXTknbm61pLUDGXQRJspoHKZU977vQ43RSniibJdXo+zatGc4WkLjwIVY
QQc0V6c9YRR88xbTaw5Sp6ZA32jDQTKZh1IeUV8w/gMR3/twwtcLD99MGHAX
uB4OfYmqyFj6A5frTl5BLoSL5aUNjqJPNd0nD7/9zwWG0kvkv864bLGDMppp
tx4/pXHIz/E+ipIZ9emUftHBHniHdv0D4xBcz397BFnV5IJpl0n3N6lu2U6N
2XsMl9N2Wvgeec2siRz6JvuhIlJIxRfqlOcUP0kw0p7fW76HEy7M24SRKu5a
EcxdrZBaoV30iNPmMCdewrt9T5/WoDWM1MwlmW+64z/oAeYVllark7zQehwL
r+vTziSbPiilZPmfSn/El8ut8beNGcSM/vxEuwgSbEnLmGonPnemEiFisPbZ
u091eYCqK2lDmNeOLiP8cdibsZjhjD2mR6jIZq5JIsSifAKZpK22jtIan3Jx
0ExKQD5w+Rm+JE9wZFG1eym63MKnLc/AJhHubgvwD8yLjPhdq8OvhfYdhHM5
yuiE0QnK+zmf2dQopVHwc18cdz9K7RaYLMFz2TAdAwNdvsY2jTeQh7iskaR3
UCN+ittwOGUR0nz5BnMABmsH4jXsRzAzUjqSDBa2OKWKl1UN6l6ICc6wu4z+
51rwIa4SnUPf91CtV4h8A0TuM7ZHEXjeQoJQITvML7Gv/+8vTLbsd4aHT1ya
hl+ru5lljBtRs9FcowMLaXxfXRDBiUDz55vW2FKY8pgtle5cRL/nZnZzroAV
J8yfZ6DLdGTxNYW4s4VaADA/Z/8Tlnk4sj8U9ZcQfstHKdlahMx3cbbmqgVZ
ePgLuoxgDWqW+NcRZjZ1BMzJBR/xwAoQMsbE3ckYHHG1MMAZv9AV8wpy4Uod
LAhdOB8y6ZtQ0IqsQnklf/3r20ObyAFlwMLg3W9nCzpVzxCHo/RXr/F8iQPZ
dvo+qmYm+yDPCA0GcNe+Um6AtSbLzlC67XWTRRmOsTcv9N/sxuxRZ/euzpYk
7jTDKKpK9ltIOiYxdEtZIwcvCdP3vLiAnT3TUS0lZ7DlmKNyySx/m9Z/Ioek
8M0goCUPGBjW6Op9RvU6qYfkfvyONl7bDoxLZ4YrMYgAuVKdTA4vD41vUvzm
X6jIFtaAzdG9kIhaiZEnFt3hJp97eMW/te5gcFgmDX+ckaUGnSRVgDHk3FvD
28itq+KN7k5P6PYJGnjdO+FbySMGCPrq6IX9vFzE8xbmdmkyB75eU1lNCltA
k84DpkX4mXpWfoiw0ULGPkF9OJK4Cdt8C3SS2mtxO2IGe4VOlnUEHhlqWz7s
Zn6lEinAYHLETttWFHZg6UmFzP8+UZ1d89wWJXi3zHn/OjcLlTDYPFlIbyxi
G6mEyyoOx197BArMeb+gjq82s5ytUbSfc2X7ugVmHQixrMCKOg3eWGnGPS6h
SqQg52U+fXGexHuX6IQJDGXhLT9d1+IJZ0UJuJnw2WnmZQ9WnNuHsHRxdlii
t83Cz3+eb1HT/OtbiNqDMZOo/KSSLePD+/0UcOAGZJjGLxc689Qf8/DHSsfV
flKWGYgdmxs5bhr9xdfrBVZQel3YAj2ExS68NKa7HddTqumlMmgLRHXtOdW/
JysIaw6bVwHgnHOAsqoAuKsRQ+eowk1Fk0PKwLGt5rgk/arIGTb6G7eHVtIg
pVWTMBhNy2KtrIPDkDL5c5BS3BlPn2Nfb4J8CcN20PP1O747De18gY48uDHg
8K/7NGE0Kiawvwtz3pxnn+WeEyZ7im7ZRjl4fu2MypoGgtsahETkB4pIJxoe
qrDnK+2EdTiAB7R44ArqTdYilEw8wGPwsB4HX+CEBaaIBvCs3tptHiA86YmL
061NMSCB++6MGe815t/YfspvZD+f1JkazaPbcBmPlujma5SyzGC99cvbt/tT
MhcydsPGhT0f9pewdTiCt5Ze+eQllf+nULQWm47hPEefegG6rT9gBb5QM69u
jemZYBsnN8rnixFxWoqZozMaY78n+UssXA4tODEQfbNXPiN1VddlPtCapMmG
WT3sAKIWMN57+KpAKbXt6VxNz3g24vMt6hLSeMoFu2DVaUqv9iZ9zeLGJWSW
Pih9YZoYjwn7B4ThC7Qsh7KBB9fGEWjFGxPegJeS2DJQ3rg53hm80XcdSPdj
Olesc/wAgvzBbA0rRFYKCPftTTi4gW9i46j0bZONIikxpF+5eQT+M7PRiccM
QgIzqssZ0HQjmd5BXZlq7qhzs48qotGSs0f1gGT2RfuJrMTWnuo2UNaL9CMH
Ph/aeIb75IqtBqjEh76vhMZXZhOO5FsaXJ+86o6VgJq4WDt6+9nPAwckbEj0
vEwbd6OFQibK6zXzf7Oa8C1g75VEpuzJJVcl8+rSXBBomuJjZ+c6PQzb1/Mb
6MckwEHzcKGH8s9iaCIXgR1O2SUenmYD9lwNDOjlFz2X6hc85zDbfoCzGYL6
LfMVz5xFesy9wBS6h7aS6UH3vCv3wniwMlfmKYMz/SIftVw6HYQ1XEcyrHpj
Bn72hD9HSr1xPQU0+o1T2zEqec3RhpXFC4j4yZk9xeMMmFcDqiGFTu2hjrhs
sd/ftflFaH22kk76Dz5CNHlk9KHM02fPv1tl+cVuhk6/4ZYqwWEK+RA0/uny
+9t5EVpGuMDopqGdz3UfByPi2/++v2md9PJH3ASYEBG+YEdENYfk4SOFD1qy
h//TJawoVzwEcxKNz2DoJT1Aws3jWUof34ne4r7WWBpA0tqAtpqZpX996hOi
PRun9/MigMQoeKjdseQyRKRIjUnYn/UCJSBTwCTa53VpfMxafFOLDQsa7gDe
u/g+jmvY/FaDyuv0XHabmUNbKR5Nvk5SFlqVVQjngX09vvH6oJl668aBip+P
0zubMN+64KqvVNKFm69epif/UVFu2z1HHYQ3pMyaYaCS+MAMhcTMdSH8nD9h
UzYgAHFjMEK358VTA25OV7Kcfda1/jRiOoMpvwECFHHfKR1IjqPnan0QK2Sg
lf9KIecf1qkylSbaeCXJy24EG0wNShZOvf5iGjGt62Hen0ugvl+CRt2O+DDY
/HASF10YKs8d4BwA8A7yJQeYx9v2AVhD45vwOPDNh2ma8SISS6v9BKZhmjWs
3RIZGoiqDsqIXPgB8T++LDjDlOInFydfgDBqKZDXqHn7+nu1EnaLyB/qGmoW
Li6BsdKt/wekpgV/cvo1dHC1YjYevA5l6ClTW/n2SwouLMXoKP8cwLQETKg6
7c3pMXFzjuysfzUmXYlSZkoujbOLOYQhCRvuGC0XKeelWxiSlCXJwVnsZXED
gFjrMVRKFp2uy4jDr9JcifSN6or96q7dxbh5a6UoalGpQuPwew+BaF2BZ7n9
POy4Je+8SF2t3fCYqu6KInp67ZC74FVJhOjd/FFtfjSj47Wpp4A+OQIYHG/D
GVeCfVKPDPzkUoMaYxYQel589s9z58fm5Re6vSbmS7SIqkaOBvzelwj2ALyT
BxEKg2rT6RfQ/Ys5l90KQOJScNgRZmi06+UgdSISJ2kncCw7kxdqz19et24U
PKORAFXlOtx9pM3kEgB6mlTCtqECYSGPatSQp46KI3XdyP9J/eX5CVfBV8CE
u1oAYZB4CbaPhsdXj6GkYrsfLCUGpnDq1qzALVB8CrcHTLSn7qJ8pqUj7/h9
fGcBfelUt0J+TUWkskgYFZxhrnp40AafYw/fGWAQ8RWyx0J6vHO/Gc/cYHfe
EM2gUIQkNdaVl5PT9GlyWKkxyqO9ld9xQbDak8IaM7naUioDncO+jrJtRbUZ
nyjv6F1xZGwHz9yMjlPR1jnbUfqfJlWSopncArx70BHwrQtYvegvYdvMrf1u
YE4Yw1pj/T1wq6+MLqWXPi+eQABK1Ce8eBcSnNVT2m3HQF/IrHYNFHATaHcr
WyfjFv3TcpgjUcGpzeQCmsrJLTB18X+Yr1pZTSzNKtDeToVQFrGdnUtNXLo1
hXhazCzAzHVBtut3DBD3Ege99GY7fJsH8pDD6lroW2Kh8eIC9ulaBSL+OWl/
Ixv5EbHk5aIIB3Sa48XXe6TeBBJk/9VilN1DxkhzNkYMgBGdCCEPJapdN2Th
mc1xfU5d/iZg/YONupDq/S2YL2xOnOTSEzSnNQ8HTCQxfYqgTcpLQZRfa8yz
zm5Be57oI6OZuTSKM9hNuI3ZUTts71KTNUZ6CH+IHIMob0cBDiLeQEi7RJQ0
5u8vyo3+yWrA5EYmselxMEzaFNU4O9MY1WOYH1gBQkLjt10X7Q1U5CeIXj6S
vFn/6wDdFjalMMHE0cscAc5+xCCtt/wOdzZJ85e0nkfULHEMTWTGcem6x1XC
u/XAZADzcEHWLGwcuiAqyvrnwVmBAIkiZxeFnz98gOMm9ZowJekUi9lmpiqV
Z4ppVUS/C2cpdi3zQuep3WpGF34GU20MW5XBeWq2m2vSmnjSLOmSV0wuCw9r
SBr5im5W009gx9Rty4ZWX3E87PtITPU/L0EXP9Z53ZCsvBGJ9292sNxeh4GF
q/H7DqMSO9H10DbAeo2prCIm6/ufvBqBX7vUGyUzdpeMP3XGZl19Pm9/qY1e
X9WPk9ix670hvNKOw0dAkSSdCd6shHro0NDLc8iH8LwPfDQB45ftczSgZ8Bb
DxLbixwuUz4nycHaDMefRDeShncg2z60eOF/EG5jAVUYapSwYhFvrNBUbsjv
O3y8miuq6l0hFv566O2X2coqjKOKhPUXhxEEe5U8uWMd44VM6/3mSrmbg7nP
wbDuuiFaSLxhauNSCSbHm2DkTYg48U7DTCLY1wKoy74/aQTvUOCm27m1y6Zv
ByBdqfkb4ctDB+B8vUvZGoflv0XmXwOImLW3b1DTVhHxTh0/fBLxABx3V4Pp
gWHWTy+VSv+mmt1ePeYcczj6/77rD7smhrupmDcDwjFnzfEyVfoukXqIjT/J
a1yNzsFCnhTev/3G3+5lOwWhg46RzyFZinDcohRf+gBDLM7rRiXblKCKOTyG
VXWAbX3G7E1t2US8xAKwOF/8cIMW4zNfTkhqDuj9qJtPi+a4lZTenDG37Nx/
kfi3J5zX96mzZH8teokv5MWErqDz/xIyTVfmRitv2rXxGDflUMrtiQyIak+F
WQ79F0cVgSbJrYVl1oVryzKfa6uICDgWtwGCy+EyVok0IQjrovgnSXDOF87Z
X8kUZ+0T95M5mDfqRR1hagW530yH6Zy9Qr+bGTJ2Ig0H2QKaikDGbl8yp6+G
Ov1OviZy8j9BakN7UKxKwBobIAyASZt8+6wJ18z29BmJvpjSih3gURO7Hv3K
DoFRQZXR+UGqyTR5o977VUDW5pJ12O/86+BIkDJsF2aNfHSa2rPO0N1j9cld
tKbkTAyJVHVFhmgcQozyJ7Vcec20NWVL/5MDCiGoMzUZp5GMjYYnyGgYLoee
37MY2W4PVhf1HGvg3sy5+30s5UtE7nUYu9ydLhAAYgor3suM3txAv4mJDTmA
62Qlp9/ii4ieGmFgoZksriuJ1cgT9M8oNZ1L+PAP9sL7Z2eGy8L8wmdgE3iJ
2swmIbkjKdj4zIPskuwEX42IQhS7GVn1v7bxEcMQTQ+T1vBUHaO4khGGSQKC
QzmAbKZQarj0oXca+DI076x9q1ufOSiyuNcNL8TAa9safQGIkqHFJIrSHxnZ
F8dpqaId52pGB+Isr4WsQaBmSUiIexei8pq8+6hHHA3AaDJv9OWw508oQcqI
RpOzNuuv4QtD6mKn6gLLs719q8cJUrHyQnUvd/alVJ/BjPvo0er4uBQaDU4p
8wGXQLW07L09czN+jxCyIl1fmmUdf0LgrorEo4nlAgOYUXGAzD+OML2UAauU
TyxM64hXlXBsw5BgBJKBmT52UvqY0npSTSFdHeBNGxiNklOSPfdM7CaZmtI/
+66slbgt+l0AMgZ5TpCf5KPIwRgJdo092F7JoHZJRdJR7LP3AydjWpE4woK3
gdrA7gMoaaBdPdAt8JU40xxsFmzBzKSCvVzRDWb9eg5Z881Xoj2dRs/ZdG3d
ALzP5J4NDdpmgj9Sk5zYZfJtdK0spOaJmJmUTifRJ4Gt11GPbsRBFTeygwx2
/aBGG2fSXJuXQZk43EBe0PSurNEDC50MpaFsBmYOTuby2O0aCq+RhrI4ddv6
G9b0Xc09y0oqlEUWsc/iFg2si/hstOu36F/GJp+vm6KH30pHkcQrpw+KK1Rr
DyxIwALPxTzOpRWbH4xob4y/nygITnD8gcBgpuhH7O4SK7BU/ZPmB7Zf4vf6
OsV+NTbT2L38zr3Vf488QhkmvZOiZlXpct2c4GAptQaVZ6vZjzC1rMhpRCKM
LPP3242pui0Dgnna9n2xzLPM+GrJpfC4ZkFBya1tgU6O4PopM3cGovLoHKNk
EcDbilnksIn/qt0ODBo8XJIk6m9WiPHTMLWH92N6lr8ztdmHs46cJDJlSn6R
MR/kMimMF/jppDCtHAkDIA4c5lgB38S5RnX14vg8MrREHhUrsfNd9gbdwtLY
VA2tqKm8xs6ZKrG4sGbr0brQrHztnI0/bBvdNf2CvSDtHqcakl5pmj/H1dOh
DMI77lc7YZ0tlP7dQXn7KnFCKGKH6qajSgP7m4PqbUHG3g539SxXZ8QiBLKl
yRO9NTPEpoLl0ERg9PEkRe+gJLrzztSr0CUjmtE2eEqyDawU2BrdCKBpZJ9r
uwu5xHjOz89ZS/cVWBkYpRL8JFUnTg1bCq9fI8V74QCQbX0OLlUAsooyw4I8
VP9o8T1K+pu5d7RBkw020+N8/1rwrVwO4rZtUHEBLHUMwdd9X0VEjb2qzb+5
d4OQgcBAfPR2zESstyG9eMTI/XCMlBV21oBxUtfw0wKFj38gyv2Oi0/2Bp7Z
lMf866bqCNz2tKXCdZX+6cVJNE6oQIkmDOQvdxlJrXSr0Q+yE70eDsrvrmgA
mMW1aiQoI/3Po+5WhmmeMFB/Zzvb+eeD1LS6zP2v0uCSSbpoaKtEc0sr2CV6
zplBqhGXnQKoiGgyiZjwnrWzQf8NOANwnp2mbW6ZXJhENQgrMcCV4+k9fa5g
dYOpwRQpHsKRETCpHhl2E0X07lUt94B7wg3OF00DcgfxNK096L7Ci5i1Hb5c
nSwLbyUjEDuwwmeDGtuz4v/vbjdGlS9HPk349tGQhwsZMbPumxMcuIPGvsJN
1a0zEsRiQykLWdC2/iNLrpxBB9dzj0fmCPJHmyrsRgQCk98KxmbIh/KTitAT
vL4eck38H7RTr/oEF3E+NZeB2fwexgu4o4W7wTVKhnUYeGDcANSwvyoLkjz1
ReMeKLTwiiAnfIgM/BC3z9dzBcFN9ZfkrGeTObOaQzAfjkgcLqBT/0Qr99rL
5zt7+e5IwPo0EoEzKKQTX+RkXVYH8eL/3y7V40gPLWxv/7D7pSjaTekIkhk1
lfMV0+lxMIeuvbgawgXg+SAWX0PEJwjIlBgMK4elDbKTc+DqD5S4qt19IMeO
qT/TUzqsTzFPWs+JHswewm/igWTrC2vSewGrLeb9mBLCFBI1/WWh9eCEWaPY
odXuCpEISCnIqmZjsq5KPkHTDKR1aeOf9yjFgiQq7d4smdLFya2kUcox7Jrj
7H4LcWoXZfhIZ619r+a0oFo/6FXk51tetqyerTQ5uSdFIRZP4QIeGbdHMQPK
8zw3CDOeMvcH65+6tluWSa3FS2BrBe1nAutocOJV/wul2hgUWSnca9S3W0iG
B5I94u5TPgzbR0kSPnruFhFOCPG0AZFwtRxPVyFFpCHB7w3z1P7HFE99iVw1
ahxaALbwzNomxcQ0eX4g1iN3N0cdg7rZZB3eicPAAf4Sj2G/CbmMe4x+nz6L
5JLwAn243kiWcqo9zOVxaU16YH86nN5ULRCPYzq3JFvGcDNFRi79o2NBJ/Qj
XrhPp00IuzpzQpS8fKFxWIeBfAhXTHGF+UIHyYlHx8dwUjvku0xkxn7fSGIh
dcQChomHDzEFbgYfg/zUz6gK8yXmUgJ5CJeArbjEM3GMBwVVHGWle+Nn+Wwc
l3f5l3ZhtVMkV/P/00XyzD9T7u8jlwoh6gfYXP9O229mlbzLXFk8g7CdHGWX
IuJn48FVi+V7QebCniOedlMr23rVFum12JlzSci0R0vmIAL0LyB6VYEqsW1f
ZceW4zsOP8Ov9XO5RLJuKa2yvsAwxfvKLAiiVKkiRgtBj21TrHJvYW54TUXM
Jtnyd0QbylReARUiJ56nki3tCXf+1Xejbx0XatoGSFYCpqQEHQzmxeKduN61
x30echDErS5k+AVJbruO2RI2WYzl2lYJUQNjDTQfgeW1ckPDDZuhJOuh1xPr
S8ZGOEJg3XoKB99iGQeV+ybpabUyYXTBBv5Wd7M7M8MlJcAstZiUGHyvTz9m
cZHguJzfTGneQmzm5F10CM1KV7pIHqqJW818a029QkNeqHkLnUJXzm0pIFt7
enyyVfYYtfC5wXts+E83x9wxmYzhQgSQY2jTjgSbL8cCnsbbcKA+QhBneQMH
kZBj5sQLB65CCEsv5hNT0syzKzCDZhfxD0yVVdo0GSLl+ve9YiAZu4fxlOo9
1DZWTCd/5CO1ApB8mSB7iCmcEp8Mr8/1qS32X7P6d7sXJ8gTmvaUy5sGEVUH
hH/IaQdBuSZSh1p6rwgfxEUCmz8JaV19JTkJSjBCztZm5rSgA8u/5y6BnCrK
MwmxzHfh1RAqUmYSCzrVdsb2HJvIid+ggJ2c+edayB5ZXeaJlqYMJomPwkPx
Ej+Ngdgd/gKCPxgtfAP4Lf48ZjPt/+X8snSbPB/+9YAcvt1DUYpDjRuy3EMb
noJs6G1aYnDeFePgNcj+4cTjPU3Gac36LUOxn47/BODTI9dMd6ErTe7Qkg3O
FL5Yg/xPvxvZHaSq2g+oAHtsVg8SR5BvPU/AXedrDDPLo23sk8G4TBwL2L97
1AyrDaR3UgGNuqXZZcvaVve0d8iY1KCiYwz1qXM5RpPf2UQQOjMTJuCHsVry
EOjcEq7DbhLrEPbLoUoojSqoi73izh3eXXcwtDExTxoEyb0yS3mds7p576EJ
bk78MA9AC3QMCGnDM5/coAyolWfUvFXIUT2vIj2QvpLSI6MqbvfFe9gRP5C5
ls4JeI3nnX/wQDQ/xP4qktiGHEyTah1fOaVx01Vud7F783jBMXOcOsxVfaYA
U9pYknPT/TWf9/1EyaeR2BQOPQRZW8No+L2OqrR11c6dX/1sfhnjEvcX/5y1
2HiBG4i5uoKDPVMHnbUN6zP0PtLWLAXOEKZw4M3wojJ8iGhlG5t2V4YLIlaq
Q6I6iVTdVCdCSkl2tKSRUyB0jxbBTOenowKVr3BFm3w8pj9Lf0X0eLA+m6WH
FOC2TdKtpStffR5O3tJtvouhCgrhWHAJbkdvH/3jGABLgnFz8iyvKNox2WIA
/qbSXj/CK4cWapQRf2zC0zwhUBMRyabLD2bp2hwxS7drY8SnEB5V12qlBX5E
CGt0uNTbNWTVJmZZAzuspPSyZ7wo/YGdAqPXV4R2NCo0cqXYzynCtUT2NyiX
5nk07K2B/00OItlZsk6zXgmcUnRdi6fXH14B1AXy2icKM1Zwy72ATOvSwQXL
DM3Fojul526SKPS6JSagIpt2xHupN/tAPfrnFbP+npmeBjYlUM45R+/7Z7nC
T/6mDMABQBUzG4+vAcXRZ2gRl7nr77j49w1Hy921i+prgTsBftHAvD4ZZ8A5
JpnOMCWLdK5xpXIwTPKVRMHQgHuebrNj8CxtACV0XBsKCdIxJkTPTEtzBYh8
kAqmDhcKQmOANfxHZpEjRaXibbm9yfh8S4LUFtQxk7trU/ko0phWtz54e4NL
GasKl84Bp9K5xLuL0RN6rvAOkgyZoXgsgpauYF7aeLcA6HOog4WI+Y+jXvaq
JsRS8zub/j57uNGEts40oR1H7bkOjN7LSSyM46Lkaa60BV+GHyCLBLm8q9rw
jsIhOAk/GocXltZqOXvfLqE9PkL+9T6cgdcMQ6r/2pqv9H37b4wT1rbn60z7
BymK5sx11ONVfZGsEIIcRbYouCpP5scjPxXgSvrBw7WMPQ5G0IPoFatB613G
8lnL4BwgbG5GYv2rljVoZngW2bAuuCcgxBYGHVyn+GgicG7bgAF7v2c5z+wW
luSa/kIkYwoXpL3707LAIrJA3vO5pK/SdB3xRukLyomeCS9PqHbdu5SLjMkp
/NKdS4nHwRo0SIGk4bGv6jzfawA7o94L8whQIwhllkH4hGyR0h3p5x7aHePM
7izenbYZwY6fQFEZoDHO8dApEyYk+ukkox4aunJScteGnLr1jo9d3zemkvOu
JqLt9tBZiMz5TxTJKf7NAfTQz4jrq3V/kVYzUfBabnZQwoICOykQ4/31nPM8
TXr5Efm/q/xeq9SLMbue1D08m/AVl44IoFp+5V8bBlGFBsH4LqaKIDv99CkM
YtKCyAoTtF2WhOaDBm9vrYSksHfFiW3Rm+Yz8HU5wn5F52QQm8/exqh4K+gV
wnCp+2qgmgwbhLcXSqPpDQIf8AdJPMLfuJBjlxsz98qMpTq6Z43ZIu6TkP8T
7i3xEA9iwKx77wWyLdRJMKTBtMGuyF/3lj4DvRE1lMQqhfvG2uzF/9PRt1oy
LQewZepy88VXFpBMonVW0a0LqYe7M5PPIDfaEllfAhG4HhORiVBc0sSVK8L0
iXMCSSmkufvOlki0HR55KHzDme30iCIF+UK8OwIZzsrjmizeUOo6wFnJLxS4
gbhfcY2yDcKnzyyLCJzf9qBXyV6Q2NkHkNxfx2ZZa5HzG/9REtcJ0JesCpjs
G2YWaqjofYo7MFCnzIi/7uuK+exAlfJ0xLw7diVL2oAekPl3kssCLnpEg41B
BYL7u37pLLWP6sGMrD8sRpWdHhrZzJP+PkoxxOPylZZMlvxC0oX9ZoFJnKn6
OzSCMM+u5hoZBYaxHC0YgoChBNfQlP0R8n209C62HqIWtqyOfJFLXUuOEaJO
2n0YRp3JpCGWLNq0702CMwuUB+Erv5MyoPL2NEd7HCyuGCvWw90YddpfUBWH
22hTJXateRegUsZ9PfHrnjvL3XfuL0UB9heMjyZxsk5MnQKFmBTxSS+FU4Cr
ZTBVLSxN8Dacw7O54ZdpUUGJTw5/jLa3MHv66o8EqAq3Rzzz4w/GzIkSkBW5
RQCBdVBAshhpSk+7KPgz0GmAknJ06Ng0Cd7cv6A0B82Um5ed4EZ7ZNse4ocD
8N0wpsV2wAJxLfYM0zsB05QblywfDKlRE6Xf9sve8zq9S8b0JbGYsOQ+Hlo+
9f0XKhWEf7zPVdJlgkNiasSog0vIijGxytrHNTdYeAV8G4/MPsFmdJdN5sEg
n9zrGO0bjeSyi2cfPL4OgOmUX2rLB68kc53mYUxZFTTlI1J45KeZjiG+LRtr
p+q97Qh7zjwsCLoes0wkh8MM1rFIXm6lbvUR+uA6W5LT9nFfgHtYbpltL4wm
acPKqDoHaIx6owVTgktrOz3jv+fn3MK1fVYfIYV2NsGEYwp0VymPzGB3JXXp
5bkdlKQN4YgHA9lMVbtaMB1MvwruuOqeTSf2hNeEFTuMt0mdvWBsWzBO4T+0
nLuPMqs6PRyDvuuszUBCVlkmBksxCPzGhj75Q/h3AR5McgSst5ndEwv1go2t
Yrz+uTAy1ZiOD6tEbqMsrZmwPq1qyNLtCzg20j/TDlyW5WcEfKcfGHfmDOny
x7T+BWghKHhIGcSXg9YY2PrtB2UBZ/ToV8+w9retoZ6tQM1TzB3a+ksOG+Rm
qTo83AJtOLct+eG3AYFHvnFRaMwShuCE44ydqcMTQC48O2mIWG5D7s6aPFyt
UTeh8sUTvegaTzJQvGpBNilYgqiZYlWu2xlgKEtqbwJQx0/rVoLSSDFhAVkA
KEPfR5Nq8vH0yFMTm2aXNe1l5VpklgLEmyEjK0PMS1HwbiH/oobikV3Zd/Bx
tnMpdSswwyUSquBjWniqESTwGjGjukhsaL5WRuSqfmXNR1krEI3Q2LV4ZRZZ
Zo+pQowDgvyL9ZFMEZ/kY5DFlDkv0DbbIhHaPkVTAOd9XkLfDC2zcozvIzNt
8L6gWLEy1yFwaFB+jvDwVp3BQk6vLrmo10bCQ12ctq7andkMR+0K4JL4T9Pu
ANX1ZcWDU0EHQOeZqWnYoYCrDGEgsNSYMpPhq9k1fFI1lQ1BFzt4bAXgm2CX
i5/+BWSzMYsYhomwK32H0JZ7h76IyB/LXhn1Htfv1LSs4e8cXP6RbjTqOFa0
zyVWB2L3oql3y+cRXQPFQjQpDy6CmRF9iPr4Wkd8Pd4vZN3RhYYGyyEMJG68
ekDkPkde9+usl2lLOpCqasLrea5/ll7yMtM7uAlVZzBb8Zmnh2dCk6Pcw1LM
56WFD3qN7y9q4yknfUzR6SX1kp0fYMIByBQnF8GdLZs2I+mRoaBvwALoRuwj
cuvYSiWfCSEkZrf/XJgNSem4VQVPfb6VfQrSgs2yWu/AsYW6BSO1kXQi9k+J
CwKrIB0HYjUBo1ItIKYjUbkbB/cmmLnI0oOS6vbz2fjC8sgKUhpfYPVqqRls
Ad+Ci9SmS5ay8pdQGvXCKxSZ7MjCTmYYlD2JKe6mPJq23M5e2udgxe/qFOji
A/oRYExvRLJxYTgmzXUGgGAp/VGzTj7WzAybYnftjzvUrXyA0wti3/JAM2yc
LZ7y7m8EI2qYmkfsfjQt1ti+CC/nJFH1BgB2aWeUzu8t74Px6qmNFD5NjCoO
8TYTvxrEtTbMyKqqpCZuu3rnmgAyyhJCtJFvaNYlxJqm9Ok9d4GNpGBCCiWe
Igq0Uyp7G5xt+CGpOQ6JPj97Du5xIH0ymefUfc7Go7ovuDxx23Cm/oXD3H2b
gliKUNHOW0gk/0yHnealMcANhFpKRiM4KyxVdtmEl93wBhqkpTZeSBBwoWlV
m6ruIcnMiCwASGnLbRuzzGbk6zjlPd2Mzq8ZBq83axOO+Jdt6lM6Ml2DLeC6
45TocOLo/0TgzV3K952+v5DWu4nFB5OqssAQDM581DN1jrpE0VVnlHvWZsOF
3ocSfACjcfikrAbIG+XLDtZ4tW8PPpnU+jJ+FjDMxrTbeie8TSzh3WtegkPM
aiCSQNTbhEaiVvdtyed52GYoCYEtwPAbIgEbZAH5wlZaaBOEVSri9cDimdMr
BarWZNWC/EO+4jvJ4TtuKdqVE6u/ijn26om2AS81hkOc99/zt9JbSDVIfbkL
vZi7mqstHupijM4EGqNz8FeGbtdqcFsqT0wYwNOEbGBIETikWXp82A5ONLiS
8B4at3gnQ4saE93CHdqSgjnRjbTb0b3gWZk3K5EwE0plAzrQg3+W4dz1sy0X
O+IlzrgKt+7CJEwdByhR4mHli8CtyZKx/HDLz8qaYjlmunEO8Sk/j/+qqTUL
9y9BgmMrmp9ke5rlTZAQOrNHhfHS1TJIfhXrgBEPOg1flncqy79jUpC25Bv0
pm1KuEjMZLTTBo8M48gXdQfHlC5natSHjK+oXKKXa6HO+OR3gnPM/MOUKwmY
0/EG+zlPHDS24WLST0NKgdexGZ15hBgm4mo48kpJFHc5aebhlCubz3D7YprJ
b/+41VNhUVcC5sdNvWoPZ/GHPp4tQpPvjTYu263O7cg5hsclA8ghYkrRBFqO
idCWg8yvWkJDOTZF0RnIHhTB2XkO1i1W3jcGjAx+RSFuAe7Nby0iDKrLZqq7
EBi8+tHsQfO3x+WA29rwIHuN6QBVWE84yhJ4wSuRFkw9oLCcHD+ywWyIScfq
gviLzvDOSwDRj3eQhP/1/528uucb82UWb0UYO/ixfrZrPRNdCizUgyJyEUNI
gO+3VYUZsR0XL1ra5WM1Y8ABP8W96rauvEUMKv8N+I6kDKHdqg80Xd48l4JL
1juJ14QcImR0McZ4zPX4AUU6AzogoJ/M0k4eFkEy/YrJGZV0iGEYnd3JdhrE
zvP3r8Z+1I8tHEXMkwlDME3neejXlALMjq9o4RJNCFPRRCYxXzWNl5X9Ay/3
TOC0q5OL4JifZ9igFxQQm6AmWPrrijtAfd/LirUl1xGrYM/1ic9CzP0wGvdD
EDVSwVgXi9szKdDN05zka9fK6ITXRylkUjIpDzgUjKH9O7wovuUP6CkVCOON
J50hB9wVf5BndJnqXm3JgYWwCVnQLa6tPwzXEWd3wq5sORnljtwGX2/o7wzX
V2LMpNuxWgPQ5pqMHeQ+2ETGWfBfPmNp4BXWCeWfo89DSIdCJuZojIPpcmQS
eQkvvvzgQpvTJ4Ow2nsBFCtd/M1ALXQcUMOOP6DVrtB7RhbMVPNIAb5tfKWC
Vgw0LBiStW4FKYQd1zTyu73mpkFBdukrRvK9OWEGL0krj8jHvIbrCt19XABI
rT5JL8W8sSBuArruamDZumcEAA0olVDXuzzznuLRh8UlxJdxWDBxp6sitmQ6
he50K7yQriLDte7Spxw0L16JhgAWcz/3UucSHlo40mAaUexswd71mjOGcrgV
0cYvg1diMeBPcDPULPLTNja+3JDS3c10dWdX85qA7CRKo9CLdQ87bD1ovyIx
2ppw7hGWc811FpWFctW8r6u2mc/ktnxh4FcmEmbOavFUjq6gWIIzcQOkiOHt
NSnGn1zt1GDhiFdBHEY6xiP1HnljH0X5rS/hOxXyOWtMDqOUquSMDtiEfj79
qKBkVONGccsr8HBa1i4Vp34VN40xCnWqnLo5a6nRXMFxBXrfKSO/of6FrXzi
rBzrOxcWQC4o4cZkNyLjOQhig9NeFgz07SXT4WcIT4zvrFha7hmDOmPsgVj0
vMoYyMkZtJD7mCHq0uwxiTEmPdEFutY5AweZzqOFq0KKyDRtV9EmsIxfrk40
s0zt26Rk3t8hut9LPh/H3wq2UD5M/47ul55j34/8UR5ctRdyKMItp9ty/zyb
kzaetzo2ZkgkBzOX+qY62CxNon9YlgnTGGXP/bIKy7UX2FoZTALKQANhIT5f
4ydRmcZ6HTe0d8LKWCxOoJZHr7QH4QdoZ/hCTSUo0FWI9xUOMsJiPj8/VOpg
bsuwschgoX8iDQWsarp0FYutZRp37qLpzMUeU9DeNz4q44hx/opujEHjOIjP
PCuNfRa9bc8yG+44bcNnya4vf4PmPqNHcRez7VnWhnMpvrPawH1qeYaTEYTj
m0ztcsXU64X3c6+3IdJOyLStiIb3ua6nUfXbCrhSgwPbSyojtstAcrVNkOYS
4WlEw9GYExsxGS1J1iZ2xNFZegxqnxegrMsCZJGhBTZI/B0l05oWsdlYq5xQ
xA2nTMxPp2ezsDlK50g01Eb2n6nNeO2n1pZwwSyxaI+LdpUfFxMtbhQBm9T4
cMa3WGqpSm1sHwZyMHm7OOvI9D44CFGFWzASAU/BPP8Svyr84Zo3obPGz0eE
R+Q/4tCiTacH/WAAGl0Wewx6eLw0nrYGHfPDGVtOlA69yHQMRjuvn6OMig4j
+HLowygBjaiQqsefDiFfyh4/Ci+4ZJutpK6HwuWgAb+tcxaiJZd4UxucaD6y
BEflbXRBws+Ay2y8xOcebeHlZe+h9wHYHzqzYtvvwVCubmypBpTypAnQTaKU
jWcxF9HlkrTJnC1T1Z1ufa9c155VYCYcp6GGSt/yYMRpKZ4rsL732f1EMKtJ
Y/SDNK8+I1HrJxN+bOsPFAKamqGFi5UXn/7AxSreNJxabfpmbNKSnms6UIlM
samLCCwekZFnVe14ny1g+YAkLMkazX3zD6BSMMqOqcGLvKO7Mdyz/7LTfIl4
uaMbooQ9c4aRTfEuRwnIC11aMsOaEVnaTJd+MCTGv9yqKg17ZwnsP6s18fQN
INkM4ZhA5AxHhlTdUIdw/ZDWyn4FVAPL6S1fhK8j4u2nGH8wsr4Se0OFBWVw
0Y/Kspls0i2TvEh01K3nzu3tmUKJmUhXT5s4uccbu+FMz8PhZJSP5Kzd6Zbk
/NA9ASlOAkXDGQ9fTuRf5RVT5jr26u2VhwHmpppqug9eKyc58xqXgRI4uGqy
v1rACW4KE7zWOQm0ZkwLxp8l38D8mJruaYImU/GHoCXJgEoUifZO4TsQQSYs
JlsTjts6DKWFhUhgFlMJ4YlvKFciuRIoV6gfnEnYUAAFOFXLsa74bdObnM5K
ebEhTHr4BuOIDutdGMaXm3pVkRo/BSkzypCLgUkTkswK9f//Cv/UtdVH82fi
KB/hDbrzyzMUaDSnnx4frUQA2CpqYwo5+6Vge6j6cq17R+R6BCqRi6Sz27tx
ro4rRjlu0BlM3ndjBpjKnvR22E2B103HnwXsVyWUzEV4RFyxzF2OTwMHRemG
7Ulp7f8FmRTvBSTDYMklxA+vLD8983l1wHTj9K2HHRZlqRHpuxOzD4mMYfdP
YT663GLMaqntNIbFxEnlPhhT6jnWehMbeLMuZIbHfiPnfF4SKrr0N67ujvn7
g4PwU8zGDMwwGW5B2MJw0TP+XRS6uJ7WtYvy4nFsROtpY7JNRhIUgliTMvgo
fHcMPneT7p+ZOxMEqVS6tqCjT4F+YKi1zV4o8JDjVEWP7IgTiCukFTjaQo2O
wHZgbEoBV/CxUSnye/OSU3Y3EsWeLFAQaLLc4kRS8G1UJ6yQI2jOyN7nIPCU
ffMrkbXJC+gSKfFDMUMRQsHo/eIofzqRQ5g2bxUh4FKVQpNaWHjLsR8ZydDH
nKjY1qPGpp9KCBPDBtN29X/4oop7B0mtH5ta+vlqKZJkLqcWd/RmnIIh9n1h
W+7BviwqDo4K+QKNUztufx4ff7T245uIzhL+5TQYyywdZGIt3Its2OYCivYK
Ztup3n/NiwzXJ9daxl/KsIB0FrbA0xO33/Qz1VgEl39Ku8OmofB68uHhum29
EiA+AaQppWYb/kus3pb1AQdIrtvX6MXnBwz9vOBGV4splXmYaEbOtuwZ8Jtb
YiHMxAOnfqoHIWxHUDPh+YIviMhkuGlK2F6xR0f1div6eLIMfIRzPVias6Qg
gkjujMsUzsxNmH/hN94VjPII18Wq7I2nL57K0xlSqMzCuUAMVLAE2OiPGmzz
oOm9sXpyflxAuQAjQqBRGvMtLpNy9WcaJt/yt+32uKmGrQyIsqzev5LiEfbw
V6WFtaA8pFnXluO1PkqChjg61Ay+Oz7oEKS4XP9IheLVgE8mryiQzFaNCa6g
U/wIJ44cQx/jcmz3n5cfQNTrLjmLUWQSPdKjcZocyaJvA2zMTLD99Uj8liAZ
Cg43Wwyix4RsVWmFYJvSzoG8OPO1LrwrQ5A3Fdm5xwNr8N0DYQtpPo02GiVp
RHl1xYkpmD7FVYSPso6w+S1DJQrlT/tB6bk9s+xXJLnXh0PaBOA+mEWeTazq
Va6TjHdLSsduUdr3y6DD5Ylp6DwXu7YngZdWPDcHJnIEAxcyWDLJh7jGJOWU
Z8+LNsaPRm86XFA/WWhCoovxu8oc8GvZTSm/5YTTUc17f4fdZO1I+Z5Qeu1X
T9J4JHCd+jZYvObKG2e6IhB693AcDXuNxgzfYvgJRi9Qu7INNbR52yZYfvrV
buh0dyLkWIJX++xXRcXBB/kiIzzywn5fUhRHoqCQQiyqGPkKWqGplsXj/t65
khU4cdBB7O+KFY7YwzgFWXRNZKK9XwGkIQ2oAWiSQ0lYrtdTCK/n7qu7gOyz
z286c/+eQ3sZLbfo/NRNwvChKgpmIUIVMtxcfdkdPNYVmei7oL3KClZAYzjy
/wh5CJ1T2KEvjnFyzcqhvVXb3RzSMLJu4B2G6ScJtR5QgheevvajZ/venuqh
cMC9HahY70jPPU+aFq1nop4SLW8CDjwdQnB2cQ2nYIWkKq7D7HBUV88AvRol
0PgHx5esAp0Vyzy2oTzCU4BFfPwqfWKZ5UVJen0z+RZVZt2gPAhe2KwgnJWA
eDPt41SEi7zPO33mOptNsttZcAH55jNbLOH7gooNEIGYuWw0klM+1PwwMnIK
u3yW1VZ9QuQlqQ26/RYnBWs4Q/mXJnkm7nhSA/ed2RNmcdO6xGVVIY0NvjCQ
YCRiQm75Va3nN89wp7TW/x2d0kWk4kUMDDHbDiRI9O/ysgre/Wglc+aBN7SV
xgHlYJKeplUERNgsLjcrD0TIjsl1cUCwnM5ZjMJLGmi6ZkBW8KpS9ixuEnR0
0hd1mbA+VOD9jOc/f3t0xu0WO7r0Q4w+783cBXofkoieI3e6RYcpHU9Dse8X
SRKRGg0/ydpU07e1zrxncblrQuEl9jlAkqshFakyl3M0b1nXYM0tl/YKqQyq
KPYT7+A8Iii+uIDuAAoSNN0DcjsSh7A7y4ifplkXtOSTMw461ZOizfBomT/y
v3VE8ASAWeRyONpPKZPAa7h0+JXQLJp7h7jHMFtqB/xIKq6sOcdVasjldDBW
35euyA8jFQHbo3XvwxsKNTSpcKCfXsr9AKjwUQt0Ux7ThX9gXClPQEbIECG/
ajzYjuzAPPoB8yfQLla4KHBDKaYU5EsEho4ExihTWCk7RzTnxvzgouLGqaaY
X61gIj8Skibp7W6Dq+OYMjJ+Ex1g/7IHWMLiUnISCcvDbtVcohrRbamnzuQg
D0e74iXdMqfwm5qZwCxbxOaE5u/qHRI+CHiEqlSS240FhK3dRQX0d31UCayG
7J0c343+YsDftfuogOScKnfPh4riG+tLVU6D3uteUIpfiWqopjDNtVbrF2L9
VNPpcmYGVo6lj0jr3KT/m+FVKpRD/Tdh6JfJy1Go/upvhjkd7Sex7EhbpBvP
yj5JwDeVo9UCmcvVMPko6Cno+iKysAepUKeT3abLCN6+9+4SA1tB1ra0bIZA
Mcb9DXFZJVnx+x2OoCNKv6V0G+oLWUHQzGMANfgQR6m4r413xXDoRQVCDJLk
GeWv+Ux6luQYpnO5WjozgO5TJtfrSh0ECfKkV4rGXrXJUuMIdlK6G9OejGgv
4j6slXSMrxRAw0mbvZZqlH8SEg2W2PbS3raaL6FEXZeoRqKSGMNrir5Q1VDy
ORuehMi6tqbuo5tfE0Uk8n4jUqMer7rI9JsDFeyd7EbytPeuODr87bRy17hE
EDZVOMMRAILqE/zmBUR8i6pUXFC6uZpacYlFbU77KjhY5WRy2fRdiI/Gmy2h
QPCoplEgZN+7b3m2IGIWf57yh+065oerhYSrnl9BKqvgs8qlloMnY4M0dLoM
pxdCFvQfYuLSSCnwycaFzCR5/vSv3xha+nDsvpn/0/wTMgddXu8f0neD8fiD
IRDkBJ+TIiui3BpOcWrT8xFT57sw/pBhAhz/jTqKL5QZdTW5XvHGOkuU16wB
wHT0mN2olqKkseQzMhAmwczKlLDXw5dBQAp4LfeUhpkFjf+KUUM2UBV6mwTQ
io3DHKvpagPv92cIKHhAUj/K3KSJwpiaR6LjVlPifGeWBlskJjoR5MPrWu2p
jrNrE9VY3QC80os8dXSjO8nLDLFbYs1o+3yo5+2UQqcMDu84v+hiWlQlYrEA
ckF3E3C/zswM8IFeGkX/ngiByjwZML3P4avMsxNU6JF58ermNOpCYWU0lhLx
MpJoTrMXJtM288PZeYxqMcMZltFNYs5itgf9TXMZVI/bt1Zn+D2FiuNIYrJO
UwD82ocBiH9S1QCRq9IeiqPwg1QP/bRCN2fIx1W5NDh8z1xOb3KnE+wRMwax
iZwZo+gq+YtbMiONL9eI4UytK/BfR8rUhElC4/31uy0lwDM2G9lJ4QtKiUuq
wl8ytX5few+cpenUeeXczTRo8UfXV2BwU+K3C3qHkpoU3bSEY9gIv2ewgf2h
EXS5n56HBeWa/TizR8hK/3/f+cMfYuEc9r+MA7CdY6uAXYKTRf2+fNj3cyi6
CnbJqQL/CFB1gykEXZvvSRKNyoVGE5Rs6piizQ+NfPMtuSVeDCYyqnp8eMD8
cbTqgOTkOssJHASRfdemWj4zxOZqt1A+jGp1/ioMrSpKaYaIAO20gay5NCAu
fWzA41KNhhjRmrJVk5I3j/T27/wac6IZ3iWUzw/Plr6Ityf/70C0o9L87o6G
/XM5Iq00+AlX9xrP8ARgFgkTpe9iwbbZ0eWcrbiht06n2apP6CSq86exF3FF
dEmrWVuHpIiRrhl9LE3gtCwg/QqcwPrrIj4u4qNR7AjWJZh8/Mx+571+z9HE
SbEpEaCzJWU+k/l3BYU71CGd2xjnE6Hq/HSzvpbC6Bc15dzNX4e9qCX+23CS
QJmEQDJupQs61zPXRcFfBRL3En5ZPOlw5gFVuqOFHjRHvE8qSQjGU4tThKxM
uswJVNC3oydkyaBSoR+r8ewyh4BZYrQBqfsKcNMXKtGVPxeKxdfAnIhjJBsA
jECf+jc/HJzpXx9FnLhDZYNgiC9su+Ym4qUi4x0tBTTNnr1UOxhW19/gDlU5
04BgSTsZqFzLxrZtRAmj9XtKy+t3DBBbfjYZoLaJ+O4ahOIeNgl27UaorrKr
O8GZzNbbeWbwD/1mzYwIeLwPkzjFtqIiYcASLuKnRthqtZQir/dqIYQBU87v
xcJ//TXNFyiIsIJsFRquXoHJUE5BwfJ2ivncs2jEC0iiTsSq0+Ydci1bZah6
DMcdaX+KtjOllAKByUaFf+uZD+BF9HTOsPpFQTqqIKCbvcjgVEXYp10dOqp/
zOZop1Ja2696xbcWG7FrqnAPm8itnWKHHYsfzx0IS7ZDGbH9zkBDfAp4gmyg
L4I4wkVckDemvIIadyenREL0KaQt1E4MGKoRAB6hKS905F8y38oOSMP3AG3Z
CcJ7Z7LTvj8NDwtB8iTZKv36L1o1+gHYTYXDvt9v0OAV3QY5iHo008RpOfgI
5HhbdoDnCS0VYNgHWZ+FImmcZVYNajpU3cdt19gO8mf8Si1GILIRW9J0BaQ2
Q69DJ2Frl2gQ4V2YG9dV+hV8/bOMzt0KZ5L9IDMkpM7R3PrtqqqyRfKyDJPh
cSQMYILhdCGYmIb+lADdLqsHSonL8wom42MSEFBaRG0QPJcDLoeArDhYg60W
NMoi1ii+RaNm15L80BDzplF+tV52Utsr+ntd64gqXop3PqyUpoyvNLScpiOh
jqBFseu1DDRQiZoxfgvo67SuPa4t5KB0C7A6Wm0p0npNAknQZ5grgWnxy0MZ
42Jox9Q7yiyRTfUpwSC/sqKo/Agy/vQIzoYZI+26ZsZTlFswpuW8F1BkWf/D
JnRjKjn/keKAWwbTvHwqLU72TJv57M4oh5k0Axz9dGbkxkPt6+H6KDYnE42r
ffdRRIRzYVgKikNOO/3uiAX4gLRzv15Hqz9B7B46+FfxhnaYPiRXEG8PydmS
e5qSb0G9p81dgwj0sLG6W42X11Gd+xl7ipMM106jYfqg1cBpf0ay/KcJTmx2
al/cHKX/IrjaLYIqigyHyLBjEBTss9zN7e+HepS1BeCGiQO/4caK+migvIqE
NlOicGy2FDlVTxfZsXXysPRFM9T7dlmQXbhRdwUUUoUF+v79fKZEYDO1Wtth
03uNBiKI+4jl8axXw2/4XJulWDif0uAqNL16aJFk3O51X+R05vG23T4YCAcY
QBco6XMAuagyAvEZA38CK3knG6l1jUX5WTPc7oyDFk4se3KhKSzTsROq40VE
jRfmr6cErqwgBXcL5dzzo+a6M4xOT+YP9oM3y/Mf5SPhgNpk0iFCclsutLrk
9ozA1UJiY1dGIozYStsiJmwqW0tVzp/mp3SC5NrErG4pPo8V23HNfPM7/ERT
SOrStbFp4ToeAe1EhjkAMXZ70p7wP3rizZ29A2s68X/Nb1MOjv2kFvi150nJ
0WcT8M9FyAlfVO//sBeynYZcxgS/x71uLo9lsPAGP6WZRsrqqTlrMMUmdU4u
T/WE2j4iFEw1EM8AxrCQPP5M/pXOUNluclnJO8tkugmEoySuS018m6dAGHuv
SufmL5lFLJO969DxxWDIWwLbJlB/eHIhdfF0lrRXDomav85VSCkZtNqqQKii
Eaj4ymh1tkvD5Bxh+RY29cdFYCEDHs/t5QKwT9lMEaigkOzs/UufvEJix+9y
0h1MtbMPx/rbmM3prgRTX15jegtDOwixISxnF49LDYA7RkxNRNClIxG6mVWq
52kYwgMQl9GcS5+s8XHI5W58C/30ZKgOZJ5Bp09o+MFYHgQj3LvtMSnrWP2L
NGTqvprT7/fCzh4enZMbPcaW7OzY0M4D1HBQF+9Lfr9R0zvMRdbEGp8gztGr
NrMzhEj80rRVP6aegkQi3C1CMeSVB9fS5AcVuystv0Jc2Cdbhbfc+wOOW6ih
pBs1uLM1+pc//UmH6OPjbLMj81csrCRFQB2vA7Lflaag1v7irCHxESmUB2hJ
nZtjB+/LKAyLCJ1WDfHjGOCLbYI1mMZ6dMLFt4rTxOEBoq7j9D/QWT4bKvqW
V9APMX2aDh5BxmFHhwezEd6zMGb26PNQ/KfKKC3bDWxx41rvX+fNEb9+l0SR
+yVRdwmvU66sVTzeto5899CeqE5qtTjF+i9gCMhKADJByJCkp39F2e4ULq3n
acD6oh0AQkIPp/lqvZOZKPV5Ybqd8oPkgBsfL3ZcpQEbv+LhcccmgMPAdoOV
uROYZ5NXXJQwMEgheebNcFNvJVDQATIi8NJNjYEuM0mcxbfjAodypkkKvpDR
A4h7oH4ztyoqlTVCqQeN9POXL8EAoqTu3jl58/sVfEeltnSiLN+9Tww9lrGk
kOPJSHVk6DgFdzmrIVE1aITgxE78yITX8UGbqyE8FrmUl17h9IE1Ab0R/Pk2
5DiMF+5fl6128hRC7c/d8JWMwDL/nJ2/2iUaGYTiBGNMkIow0D76AicRhd4n
rdoZfWFmXnvjaojFQYPDkcIbu7ikvnbinqTWbHt5dS15z/d9E+08pnxko1UA
3g3VaU4gwl/3CyhXmO8dCa5LD7gBbqk38AVPneKnu5/GLiSJ/OewQ3iC2AT1
JIO8a6qU5egN9j3IsxGRlwbRheOWeOQ6bHUAQBB7GXaYdtoUrsVgHrQdPF1U
Z5Nz26+TVvjlVaCvwIBUwhO+lsUN7q9y4SnZPwsA3clArc4wyrQKyEQhVs3x
M5x6aT7M4uhF972U5OsTtcxWDNL5GzC6QCLNHo4w6pP3rPlxl7OvwAUkuroz
lQMvqc0Mk1E4NY3H/JFbnvTXlxuUv1a84zmACrucmxkArW/n3nxOyINQNGdv
iVfoSm8FyBWOVBFzMiT6YoIZnau0WDQfQr3yr1PXaG9iTETQdN1D6Lhcrpb+
0rYkFUb/AEcUXKE0CikqZzkUd5ixlcu+9CaZwDatTZglvBNqu6iO/blS88dr
6aZCw66FHzCyG+KJnSjoEo/BvKRX1PLEc/lD87V0fMLR17xZcBtCVH/76diw
fdRxw3HKD4ss6B1lWffxkSmMW8xf4vftQtDDW6cv+123nAO/4XhziYQ5jRCY
CrdJb/PqRqw5NrQ5vEc0wpOfN7j1kuCHVdpmGNQhYCT6jA7kQadGBeyu4qK3
PTFAVddn1Xtm6jwdH5uNO1qHYWC49uaREU4tw9+aJMwzUMgKY4Vq3WZx3Qjh
Pm0++ABDf8YZz8RA/h45z5SMGzFvTEXxUpSrjFbCp3IvrBq/L78wI36PdZZb
CKglnRCZiyLiaTmQ9BCg9VtcQHUSTnzA3S59JwPKKn+lJm3xlK3VCUjrGZd8
z4Cio02t044gQQ5UwHlyuS/IO1Iz4nkP02wZtXzSfZM3/pFerEIITjkR45PH
wpRIbTa/VKZoTEVvuwAKIJER6Z0oAJOnU0ib0W1SkWPR83swSvgnKV4hjEeT
yNXC7qAPtShmXx/t5D10US7ZD/WGJJ/mT0crOMhx/PK9UNjipOYwFzyHQmZi
BpbBkyxXRv+m/ALt+qWhAJHH/BBlxqPiwrXZPHf3F3y/SegU4En3qiER9oP5
a80kkAA6+MvSUcl8fdV7ALcVVp6YiKRqvB3QvlKYMDE6eYs1UNr7cMl7QqzN
A7eQrqAQIUapLITCFfhf/MOMUgXkc/Gb/L2iAj7RQALCF6bogxP7ZOJI/k7I
dbdxArS/nmRQuHHj31O+dB5v7cuJT6AIiDeqmzHugv5knfkcAp2/6U59Ozwl
el0uine0Lo8oRJf7d2aYag/+02Hu4IdpaZdBlozZpo+EkmCMN11OG557vltY
aQ2QZYCke89UP/7ZV60JnZJzaVLRZ5N8DwOq4UG7k1leD5yKnKe97RlvYTDq
85mjw4Xxwmth8OxCk0Fj0RjA+3EGHFgmy2CLL1SHqpmn21lx1T8Vz0aY8XLs
vDJYAK7qU7qS8h7wpjTmfQuqu3uxTNSju0DEyiIHU5azDEEaMHJ/zRIuvEaE
+FRCJpepU5bgWJuXZcMVVLU0nvkl3R3qf0Vb4vP3/O4ZHCM2ltI8ReXBe5sg
/5k6I4ecZtM0LV6UdDqrbYpxjhHH3oCO3o0E/9ualyaLX1iccO1xtjdfcEpk
Z8lfPmzEqPohae6aKt9qs7p9BmG2jSj+V1K0KEtXIlCB2r2JVfYyD0jR+fH7
/WVQiJchOhPzB6QChQtC6N7jyIpXFkLTDwq4DmXMEsBU81HTRUi0kInr4yYq
PD00t1M8cQdGSSKNWKEh2lI+Y3YQwjPaPN1RpUL6eSNt/tx+TW5MSmpMuJMP
Ux5zizrGJAkZYDYayqx6MiSfb7lY3BGoKChLKERXGNy25cgdxwP0bwKk7cda
56V6PRccw9GEzuru9du0I8ABkMgt2rXrDEwuZhuOzIa1Jo4wykD5tNz0dBCQ
vaAcwFjfhwreddecIdDiJ/ZHc2brgpgMQQ8pAmlssPusVKFomFwkn1eFDt0U
9HALypI+sozTEj2KGwqFbTA3RE7cuaV9gUUym4VOKpdb9wdyqDr2scvqcxZm
EWzYZ6GgP1a+jrVbquEt+is4fsZYOZt7EKetwcRtZk5VdmvadPXIt/p8Fuid
wNYq1iIL5FvW67/bdxE//Y2LUwJryJhF62g2DzLVftdqBNQFSIzEj8SMzrju
5WtM81aWD6/lqroPv63d3m20as036W2arIpNISJTGiYHvh97oqIHHvW8I3Wg
AglhbzINaf3poSgu4WDYZ6IMRPv9WEe+88uCZCKtDShm03japGTwGIwIsV0I
qLtuo5Dykpt7q5tbbuA8BA1U8edtT/u6cg5oLTvRmnWbjgwtlUJXCyi/1RV3
zUKkeQma7ZcZ+/yMPK83Jv82cP3eZm9wBb1CIN3BM+vRRvnUsyY/3A8eah63
USqVma+Oz5TH5d4fERW3uKHRORVME5CyMi8JybrE22T4+yPbUl1yT6USrxb8
mL/vL6uJk935n5rnd7nHnQxgoUoeCUol6YVswflg0dCXAvTpBCOywnw5WvCm
hJaA0wFBVTZ9T0PAlIiwUij/n9ymRf04GdRMrZyyLpTiUT0U+WutK4iSI1x9
MExD+uqqu57bLZZAEUrwdkiZhkZMJ02GVj+GAjzFdXWf9LnHwnR0Lgg9IhUu
QMyxPScrduOP7v90EBlWD3uw+viT9vQvv2uMFIz0OJ/wUnuXfHC5SZPwC2hl
i9g4+o2q0EtcELHSwGNUxYpYA6nf/XUdKrQX1naKeFJmRRZgAn9x2uoTdUtv
wpA/BrqqcfyD3ry7MTw653t09VzzXlGYKL4lqPwork7q/94N7Li88xaT61YV
f8kfbgreRIPxInQ9mH+65muGV2aMpynOvSvqqlH4PxhmbIYA5Ky54dpykHms
KXsb49UC2nfbEJzV1q5SnZWSgs9ODDkhb6bfGZq6HcX4TWK2N90QIXv0MiWe
/rjHnph2StlRViIqEUd8lkI95fhSuGGAXW7ZEB6gS6pwzvRYnRAqzJ/QHE//
3OS8pk3c0lpPMaSz5LKtZpRZOQCYGcefkv8wb1DLNB8GyVT/YSz6x2yDb2Cl
koX4tXm4NBgebt7sOgz2KeAyaYqSbSEHgXvYQrcfKs08ICYqgHbyj+8hMzTR
goJQK+pFO7tLnhRQDy5iO/2/b9nOw48dGi419aFvmauLS4fsD/JceZ3JaF+8
SMuIxPAz8VvvmLLC8MIdRdirTVEX5sCzEwEW6Dfos+uE5y0ERx9HxaC7OIHT
+hc8ZSkaCTPJVjzzDVxxSvlwwxhDCt+NnSb64MXhfr8Z3QHD9yYul1DuK3d+
SK/PaXTot2bMkkiSQEh9J1eU6KCDb1GLOzTSYUo6E8Nu6ienIXbmXpEr1iv1
VIJSQ8K7Be5M0I0Lnn3tywgiqdY6qtoJa3DSPYsX+1YadF3AQlee+4PbGTob
3XfHpWFEQihP3qIj98aiVXz4sCL7FRYLgEmkJfop8I9C4XqDfwTuJ+mqEIOX
20L+tdOROVLfHNinzMwjePLwjilganvCTKuU3mAdADNFjxQ4qdc++aIGsCC3
FfkC5GP0RBgybpW8jDasTNfCOZiE7YmkbgKe6nsBB1PnnXveK1PhhQj5qmqI
OGOnbfJiuhoVlYZtfyIM7ur5SVX9M0HIa9HFDLJcN4f386fH7+40hahiyYfF
bJz9V9fvjs2/nsWTTTFMVDUUlUmo/XpEsHyksaIGFsvRUeTC4MtwyWwFhncz
cTzuUu+PsDsHojyjPfbYo2eoSMTPf4efdBPkV7yAMtLm0kb3mxYSA8u0yPBh
wpeg9Pexq1wQUPQM5uLAKZsP/97qO6tHDLEsE/fdwOtcAnIec2YhMYcRi71d
fplWfb59Ngm02M0KlGkY8P/22E9qDAir64quM1U20zjHIojOZiBqVjITuiYr
mLeSPOYKqrOapzslmjrfJk7K7mB8HORqwjxnh4v2sesMx6yZhRE8f8r/wdwD
jdQSqSk5ob26vAU8/tKi2Cc2hG93Ceq+5uAs8J0Nav+ypjdoBN5vfKsgI8LE
NeAqYcW/X7JBUQXvJeN2Gop6jZfMtWnFvytn43uumAvyjw2sArxdOB+qG13/
8yCralVNVTKWQyDG2N/LQ2QL5V0cgwQAtlAVvdMS+qfNKQqVePj+7ro7Da6E
t1ACDMySZdo6UvChLDcbNfyayWYAp7n4pnml4wQEw+pCZciuiL3STP9swzFs
qLlUm75KSgVB78g/+Q53JVYPuvDmJUSE0GjwFY/k7bT1XlF6oWSeTPgLua9s
F7jc8RxUlBiCYns22cnYeUvU8Lugz7Rkmf+UJZ1uG/IDDZ8rocw8yFYY5g4x
v62RrieHMHjy7/BsfPSmI/eQV+ppHMScM9KzlmLYjcs2ymWZpcVxqmUQLW9Z
HzzCfFG12xNc7UNHscTRV0hbkfWAdSEfVLl8d+vuaAY7luAvPBUhNx1flgI/
efuIYOPD5qqoF0fLJUk6G1qmhmGLT4KEVIxAY/2xWuYA/lVaC/WwmOiG6F26
NLlRMfZEw6u5mlWYramA1prQ9r9gAamo9RtrtnS5X6Vha15I1W92PkFsv2nj
BNAc7+C8aHrZcI7qNV6uf8knJJAWKMDe03J5hlxyUHWDFJKuyBpMuChMi1DQ
c13F6uJ65wcIG3Sle8HMszeMh3e+BrrdsTnfX2BpFigIHnJsOg4R+kXUfA7A
drYl7FLhXb3wqYHOU923Q8SFKIWYlCj8ZQZY4oBdQVFjKbDqNFahnGM9Ct6L
1VGhtJgDO+mKA23JnZpq8uFsBfs0t1xpGcE/elMepoabSEyz2uY9n85IDzwe
0bm+1ycgUKYv/Z7fNoKX5Z+KDFXGeZxjkvHMWw+eKkB7DgguwJkulJ1JbJ4/
QqXmRHwm+xPDsnsGodnRXwrVhUreIIQ9K4/CGE0BsKwntdiZMoHUcvnJ4/TJ
2mJFRAZ2yvjJnGPgeumYeCgr9eqgVokGAOGVlJB72aDJsVfY1Rgk+Nbx+ajz
ZiSqyNw/qbiSmMI0qoUAF4Cd95G9UUQ7mswB/r/fnj9gRloTjH/jnQ8gJgmA
sjorPxM1ikgIxt/CSHzZEUhvgNyak5xgUblXHQ9ILvOFp4krpC2fX+qgQKWW
t92ZSXuZ1tpvZgVKQ+L/Xf2g4wiNnMP+MIPd4ovKWD3FHcjSZGBSlGS8Ngfl
GFDRMQW52llsdjeiTAg6BQb6J6r6mYGAltyfl6U6pm+hxW+xmoT9sm68Kh7A
lRLk1fn46W4w6W0vt0LK2OpmebzeuUEqggZZDZL5OdoVk/mH3eBqsbR6oCb/
cH6V4Q4lRmqq2lP1rlZxGoz9SAeoeSCGu1pKJwhshVgMH5hAyWjohrkzXG52
+hGG14lT9u8UD8h7sJH1TBzB93a/0QdlspY0QRdwwQECBEkPjqzKlCY/ie84
+hHmOgl90InRbbzPBVJbNNarfaulSSnfvkzWTT6X6A8TRS6F2J33fFL7DrnX
Glz73PwIpyAp4VdQwjKKN6Ppvkk0tLX2+bjewEASU/nuIDWr5Us53vZgqbGS
/WGnMqcfIwSYPYbLoWvxDehXlYFTaUy3XPGP/T5323CDDExnHHYWBjOTgtAa
yxzM6//JPC2UBmGrbApkS6x6OXtBoLpGaGmHLi/hA8dqyvF2WA23wVKqXk9x
xBbwOvf5rm71oHVXwpCnh/tpYzn9n1qjyjzNjqIlBINlHnzFH9eX7y/ZSu5t
OEhUe1/ZZDZMxrKc0H/bFuCMgXVkgydbmx/bQQngsRNNaQgBJV0sht6PB1BR
XLJp+2ykdxusSgFrPgaXsgkXUXD4oxFrSET+EDg9BzsaOGLif2u7JFfRFBLC
nb457QC/Y3O6WrEmMmzNcxtxLe8lFT6NWPKRCIN9sYemUP1VkVbHC+gaq7r7
Uha6q+L3Uj20Nz9oj7+sC7ROv0TT4stjrc9V6hsuLn70H73/DHWrgkF/WCmt
nHvbkLjoMSccZSSaWfpJzucAhH9jXzatytbq0tCrYEUgm7Qf010v4OMegrIE
m6Qa0FfN2uW4VL2wiaWNBDF+/V/IOXF/DwaZigbd0S7QbuIyv1gq6zEONf26
Xmi4C9vusN7+okBoIwFVpSLplZ0pVmIuMiIQooW1yMjBxV5dU2BV2PrPgIUP
7ysFHrOHShh/4u6VeJAXFGcUKZPLnk6u03Mc1xFlLYP+lZLhiyehiZWkzSXq
B7abNI5noDMRIPlAxTqJybt9/6jX2li/7IQ2eMs339UTJ8ylqgouyMLU14z3
Rv+VREqy5wVmPi0D4fNNur8Z5WPkJm+/1gVfSJvaAo69sIz62swDOI++Vd6K
e7G62OQjYrm506mZlD3RYi+67VHnsVEKu4fot5uDVk/HxfziA7Ofsy65S7my
3HOUq3Xp9RN7b57SQnLE8f2rlR4WT9D97KK252Mn7RkO93oJVWHMVf/wUGF7
cJUc1enjW02k7VbSePmi5BMKyVhVahfxhhoqRj5+k6uogQMHYV4VrwZsebw2
9P7sSanRJTq6p9l+x3Vehv/3Zdgz3OwzQZHc3NnrmPagzArDz6gd8OWQ3zsw
S/WIEmBJMgvA0ZqTsoSh6URuquWzYivNWjKjJ65ERHRqbyzPO0hI4CfD2qP5
0mY0BazpTkbUYEB7ka79Nmx28WCuZe2akG0MwdwzIhK8qnyDRhY2fX6eWH1l
GbMxI45aS2MMufMaHXITOSvaIDSd6yQG2qKDKybrrWAHbJGK1KO/5kwy8Zoz
fbnGWM9vVZvYf9ffpr3yFSCTHTzxV107clvEPxCgbbSU4eJEN6C/SWjm9ze1
Q5ofS9QBhs/xsTwDeol06qf8uGxRobrJEgz/RmpnCYgCH0mFgTB4oIz9367Q
wQf/Ow4EjPT1BiIxpbKj+o+9ujH40CetEJsWNEcYgfrswy1JnjxnC0Q98YkJ
grUYnmr+kvBzFx6wAtv3TPrzDCRx0PRrQLWvcRe5CEfK/4rejXWMol1bnjU7
32+7dz7HmiBzI5fFjO0dG0c050sg42JARCLoE4WIgeYEBgE7E/yZI2SzeQu5
t9pEHdaWpQtzw42ya3ON4m3JqDKYvpibkT5JgDNJBX5FR73uP7+d7C2KHs6G
ZWR1FZ6f38H2grQeKACmKN0fhaA24RbMZoRxdMIQObkhbIQO0MVG+PXZmjfe
sodLzy5p0JgXGY3Bz1+Relen//6VJpDaXkbytStGsCzws3eh2wu1Jc9niYTm
wq1jH67bi4Zmon4OuuMd3Jk1maCeEFa50zd7W70TXF9s9NKbi6uH3Ac9EqVx
R0QmQVZVdUOX2yNGUD1KYF0T/VSRRXd5QizC+a5zUyON53L7DzTjZs9blK5T
juiFdCkA9JtlpkyCBjOygFifoOYnNG0Q0M08vkig+IOnr4sEKIOcTuyp8S53
hkruVXPFp6wpG2lMyvzMDNsG1l9NRtyeJjxZpiv1Q3MBA4jlqgCxXoDwZKfm
Vp0zah8mhNw64mNcZM4LVY6kVpVhHZclsqUUcNs4h2nNO1G/at3t8J+C5b3C
mBUCjtLll2KxrhUaPIZ++cDuHWoa7APxxdeZq2m8qP5V+MgkBSgcyeS7P+wc
5fTOAaZNh4/7e341Bq/WllDUtWJDbRF2ZQ8L5zYu43Ek9skUmTn8H8EPJvIs
sPBhSAD2sQc1T1GJYNsLeSiuIssBr28jYf2ay9xFGQl3SPGFtRB/iv8nRDHG
VQHaddp1cfaGUkLkmbXleNdIrQWtGbMm66ZiNuIdh6UClOLJ+GGLgtIeTaRv
nZtbq2mmWbKNAGPZmcnPfeLtqwWg46FwZ5DZ2/0Gm/5DtovE2pNa+kfESxnk
Z6tO/eKm9ixOtN6o0i+UCbNhNmqdQshIcpIQ6iLD1UMcorzNv9iEKAvsUbK3
FS2MnP9fsgfU6cXE3U46gKYkF1X+Fpj8yV+MnH/XM9mA4hllYjAl5AxAfQGI
d37jY/4pBX0TQuPjuno0i7A2NNyunShv4GWzWldJ2RiAcSRVq0sYSiyWQ0/J
FkaXSNU3jHOCogFhFjPd56V+V8pdNQMB1uQyvdc9Z4DZneJaykI1D+UzUtZD
tHBZPt3uDKLw8g3nP8ZoNFcZRtzXsFLtGG5Ss5RzsEJe8zew0802ueBNbez9
Zo29E2+kw6m0+KHfDA/YbVTu1Ze+RTjphea3g6z3OVusCYSG0DXX/63tt+FQ
B0A1KlMMXKIGAUzVE8mls05Zxq6mCd8vEI5421XHEP9sfUvO6IN0EHuqXpyP
n6n7cNoZDEgK+9pHUKcDN5YF12GEsCKGuwI8C0yn2/H/lV9UY1WMFEO/lPz9
lH2WNfq/AaduSQ7shxvQHN5ACRBr5GPyLSdgFXh3fqi9h3NJD6F2OoswBenZ
8/lQcix+RMEgKaPtwassTZgJa3OPzxyK6CEtPjd/zguFrRdU7DCSaywklHUd
KtGRBqo8FdJZKVrz94Z7DVeRJNx9eqDBnXSUqP78DjZFB0ZD7uf+dGDHHMeh
OKpwPGbFmN5Rh2sD8HlbwTYoEHgM0g6COznEp5xVec7WLLzGYEf2ylok+78I
9VlwXgSxAtrZVVmyYZgFyeDFfM5VxhMnIMfDQ+WnbGdPZoVKwaQhclVIqhxD
VaVEyXvPRTKN8BV064zE8O71xxH7lJa/C6slYh+nkjqz6tLax7+WnoUpQASs
IU6hfwWiRcjhuLMqrfY/XkRHOxqPmkuOu5T9GW+QQJawLdv0JNJm4SlSsehy
MTn81QyhBTOt4ou70qrFAuGj/5lj+XzmyTg2yAguQw4/0Ec3Q2CkRFGYu9uC
ofV5MD5fqLMS8SHPOjvC+T2xjKSxBILMoTens8Wb8SPSjXOGngMgvWxAyl5K
bsUuFETDzhdU2xjRQQvWFxzmhr++/JCn3Lkf1rwmO0NnMiseck4+/m8SXA5T
aTo0yWZrM2G1fyNRsC78fz7xgd9kdpLTiX1Q2IJ3ecfDTptAoQK56h6bs9P3
xYN7prXwgHJrHLRGwmalS24oO7Hs6AgR6Z/LTgbXH+FSAdOHzfjUFW9dNgeq
B7jsfam58zt3gPKBLmIzSloWytaoTkMQ+8SflUhaxsmXjrNxWnhZE5LRDI7N
HKEgJnu16UKifwPrkHg0+Dd9DXZ9V1TzC+1ZQg5+Y1sqBAiK+kLRpjZDQO+P
iy9vNYvxuD/5+Jm+E1JtSnKc8+sxrNcpePWyrJS19SjsLEC2rkh+8szyxxHG
7ussYkiOHbA/daXaF1oSq9+6Es99TcB/XEByqX79a5WBVjdm44KRRAkXzZ9k
vuyBwqfJQRHWsgT2RrH1engWSjuWO1gx636SkdyUuBYmMWsgT6FrglLaeBaz
NdPzd7dX00xBzO/iDBZAq+GB4MiokSI687K1LltlOH9kv6TD4fdwxd/fnzXg
FwyArYapiRYz8ND1jRwHWxZ6gPK6+38GbtNTacT0LvllqCYHvG2LiMjSE1wz
zGcduhp2MllrCyUOTSEiF1ie4D+Okl+xDmx3Thf6dolmXOzvjVjgHgVSVwOA
LnD0yypMDH9rVLYD8W7Qm0f6Wby8ebx3gXvS7ByDQl4Vk3Yhwb4T9SlzzUOk
XXibzy/6+58iMFjZ1CvL1o+wVXquFw6IxqvS2zIDCchi/NZp6rBXrF/QAC3A
JPvr/gFMoPbo8TMDcUGnXMNza3TCDVflY4DzcFhpFmWMZ/yvg2g2d6PxvDe0
BEDTUEFAOsK9IN5wNbf7H0OdlA+npTZruDrq9A/XxNlfOD4+H++chXgsYN74
NwPUYoBxUVQ21CbmWTCa38oLmKnAl6gwUcl7kl2IZjkqI/dmFmyfnV7JZfwe
K0ZzI7dpvVTG1BQZtGm7/Eyt6vh6wbtAMW95iIq9O6nCHclLIG4UhkspL0OE
wDtj3icAbgeIYKEDLyVm5h6nF2kCejByt25Q6lzTOUbno6zkQdwqB11ETNz3
hmGBdZKdKVS2cKDGO3JQuiQEpLHt+22PHsGvnn1vepS1EAL9xFfSjmBbNNV7
IAduT70BgUqcu8U5iMKGtxhUl0UVpzyurNolQcF5zC0jWTFOx0cPrSE8iTwI
H2OtXHlkKmmZwfNbc/gfoZ7IeJAM0kNBse9ziza70u6cMpf7y7c1gk1LrGHm
RdHXC/IXX7vPMHA5ezU454V/c0T7u4KX1/jv2RPy+S76Di/afVHIp9pUuAkG
zMKhk66sfMNBVfbAd0p8ClwCbkzJQAlg+dCtxY4QkTXMaxEULfleZEsDCYnl
ooyQU3x0kXOXjGT4WfifeUr73jREIrPioijAxjDlyo+vWv7R0hFjeSYTkzkh
rcjSv6dAbpsvuFPRt4a3lQea+9bWL73ylgatF8pVrcBkw6lfLSkuqw9cpBx/
PjJorQAJ8ChYnejgh/MlN8GejkoIdD9A9cmXBbF47MKtYacl1TJDTcnEuJ3O
/o4f6w1YcTMmhzPTpMXXtonhVwdTK6siMhjzq8GjK0WVvhrSwh2pjBi3N1fH
ZsZMUjoj66z3x7BAFduQ7MLZ0Ae5GV814V3mYZF7XQI+M7kfsZSHsnCUbXWD
tvTRWnCSnyKa/SlJUfGl/MmjzjyeMf7brtV9o+UurPKLXdSR3Rh6zTu/k909
ZXDMwRqUrowQSsH0UL10mOxIHdwoMqRTDyxB/XUUyHhKFAk6qvW9ijYLmEFG
N6LDGy55VtGrOvuL2DGSiUyEpHsXnkpn0DDy3R1PMiq8Y1WrDd51Dn63a3cV
eVP30zKI3W/hOctk5x3O+fRGQs8mSG6johUxWx8r13jZriutfaoDxLuvoQSG
4MrQfj+mH7fVBRgq0EE7PCFsAKpu8VpD/7lGdx08QZFGyONFYM3k8JiVRhWC
es4Jr36aHVd5iBQ61p6rkShlfITcKxaB5+26rlZFhgO9grVIOdf7Cqde/aGS
6cnebYpHQix1QkKGTZcfPCXl6A7mxb6tdW74gIjc4vpTPNGQurYRRxz+UE39
CbPr7xjd/Dz4y+6Aopy+D5PQpfu/yulVJpnl5bFtxEpdED//GvXSBRHoV3Ps
jghNmYNLM0KTHUva5Lwk8cXmLvNQbS2wlSSqs4VEQdS4tSSOZ9rKzHsOXCpa
Hd8Vm398PAAXH62WL4E2vAptyhyQVq2XVeWNJTpmepOY9di0W8tdXAr3xdhH
yBb1ujyRcBYxJIpxtNyZHu3Q+Eg4hm/l1yVm0673YyM9pnIZ+1wQ/Zmo7iGj
QJaktHaTRdSD1Ye9chzkuNAALWD03r2a+RbaBvE+Cg4Eiit+eYioNwJgOrTv
vG2w9SDCDVJFMC3UMwvPqSqwbQ4CgY3U2ea+CO4CyuL4whZ4Qh5HdEp2CqOI
k++r2MdmkA3g0abQuvHHwQPv3Mf0aBbnYjFlhuj4UUqJ1x54Z03CduqwkL01
mUPm4Oi7Rg+mkrxPC0VZpoFFG3zjuXGNYxhpaKOk6urYaw5A25Qhzf/lENAj
pkA0k8IjDT6PKu+Hs3JXVkYjPZLB6QuPPKpxhUL0D/bGGYtPAM2P08IYNi80
YX3kUSKBmCIPacCvwKVejkmlw4pH8/Sln/ZWRthh4YrF1lliIlHe2kP78wJR
TCnSHI1vw0aZSVOU0WqzJvfcURdudhYXyAAHmWRIOGuOOXgiQanJ558TTYx2
1f5NKhpcLMBiVOL/txUc9Ya2W0uRjlKmooKPu/tHr7njjzoppXG9jnMstzD9
/MOX+mFegC0T3lJE6AoAkbXjUlN5JMVYGXOk6XgdAbgEMklWscwXQ7a8MAUG
ogCP8ErRKQmj22pKgKmRHYjWpS+ytpFEE6ULXLOuXL9x0MGgmcbg6bvULnyH
bs4VAcGta8Daj4XZKdjMYZ/5DH0IzEqlJ023DPqGsSBoUcXo8Esb/Am33KPB
lwKhgaVekrEKYrXpLJ1rqUi/IXhamrPujjgfGHJQykSweV+xsrDl+DkNuewq
/sfuVBqsfxfPDotyzmPp6Z9hmYybuRO7zK/QimWzvIctKoO7Fkp0YuTuBDHl
EpNMHUBmCUIDFLXVpt3TISE+3ozZdMGYvk2DmWnCVKNhVaj8obIbzrDhMT7r
DMrFoiSZdZeYtHlK7JYtEAK69NjxIzjOxABOH+WpFqR6QiEm6jvu6bYbkG9b
kvDJ7sFu0VC7Yb0DhfYNKzg+FH1vyL4oagaFIhYfX2wmfvp8o2PuHdrN3jIt
8aI5HujgHizCy7nXl4FxB/jMMPefMTKs1c5c4SsHsELfIve7gKgPlt3ow7/a
+fz0wBS10F4x3YJmriXnLgZZ4GiOJD3wXGNk/0Vzn13NnVArsbZrsnCyQYld
xwIYznIXQAE3UN9QUDsOkMwyJkJLSzF5KMwf8m+buiK4oiXcUb5mpPcB1EcP
GXcCA0AElacy3DPlqtNdlEUV6NBfnswkuy8NXrp/Y5yWcuaTuYoECnLNHJuM
FHSDo+S06Cv7ANS5bjACxMDf2dcLhWwW+yMS9hdxcoqXvcB2J7HOrJNHokbq
Aco57eeoGwONewIACP4ilAdbaLkllLfNmA015hHB2rr9y3OD3ctkluxU5ZgP
gNPhnRIfW9W9uV2ox0/tymd/8s9gnzgWEpfYzRJKfbiT3Y3zxxjlXdAQvtmj
q0FVguPlaok4LkAo8Mho30B+ajNqzncEWkJqMU0w/ybCPwn+/a6B+oaZsdF9
704B74pNKSsCBxx+Cy+Pil4U6oiGd6S8p+5xPjk6mUmL9XObgYpxQHAp5PEE
47AthHvkVtZLpSNd03bdygNF++iQPhb52139pn/H340MEtFG1vx4RzwQnAjH
yT5RpfSPq79rWtWD0MGtr+wjDp5lC5fTTIN77xQYqRq/4ZiZB925u04sa5a0
m6byNQlac7ix21W2EyH0AfmqQVFBbIaE8TE+0BYcQeGAOsAQoY40qtq7xzil
AxiXMma5Td0CtCThvETEZiD6NAc7Mu5cDsnAohDxGmHW1zPuZnL3pcx2XJPD
k9Y1v43QIh+G4VKNUuC7kr5d+OcFU0SNvjOB9huDArr8QppslIKnHLxWnXYQ
eXNnhiw+9s7aZqulPMDXkim3neHq0uwcg5/2zhGqEz1uCRCSnRmlu9ClLOXF
xEAy72oRsXDqI7mlsH9HKBqzFRGRdaUX/r4ypoqBit2aTFz0ZNfM6o38qiOa
ize7gLtnnfVS1qP42NDbA+Ez49LW0cRJhUGVGYSpbNBus3uyxfPl+fE+65a+
cMbSVDnJ3P/gh1koJpw8PwJxPXSujxdeSso0M+KYDg2pBrtfgs2elNLct7AS
Dyx54mpS5RgVYgaFEksPBQYU1g4IVsm/K6enMPajjTB7XsPePtMUSsJTm2qA
d1rIltMgiY4y1k1bQqXYgR+2MBT/ou9C8ENFX5/JmU40kdAZBhIl+CKBnwEU
R0kcj6yJGnDruro0cL/E5wAGdNFD7mtQhvamU7gyvSy7SieE6DZVMhEUy7gB
nvpz0HLDrLwPGnJmv2D/cSZ9IIwGbQke5UdeIS9Wux/HFr2kvimwyt+fayGx
YEh3JM8zegSrvDsSVyRf+NeC8dCOxVjcau3uZQDUboY4/3K+usbhIGA4yiFc
txH+2M/Zi4Lys6dEGjuf+mVpI4EvgjXyTGgF1WxVPPjBIzr8EfzOxO588Lza
mDSVuNKzA4d4sZRSkmL/ti9vm6lE5oZE0hXvgm3+46fm4YB9J2QsVc48LD9p
8nEzK5irGtNfbP4u054A+HFJ1xjKoB9DUzQBhK2gqti+oaCB1ce1fiAYElq+
rK/sDrxa0yEY6zLgqL2iGvTcP+1+Pk7FCBIQ+YQC6B19DS3hKSC+CIGxJj1R
6V+gAntNLneDz+on3F5i4Xq3KPQUNgPQ0W8FzGB/n/FglF/b2M9ZNV6qvp4m
CxMezv6hX1a5T/6XglpA/1WtFXtHc42JlYzefRlD9r7/qs/6aHLinOjnE7Go
wbvr2wT/FzHDQmS/JxgrD47+iLHsyxbSqV+pDnP9xRQtHeSkonGYw9RPP7fg
Hb2/F7MHCeP1K/GexRJe9moybgU8LRoauFtAE1g8gyjd3EkgbVxlSrJSIyDI
MWQG4wyySk/UBxvu1kcERIMsIoZCzBb+cynV6/A5R0cxzE8MiEWze5Esk0dJ
iYxtIOAnsm3lyGT0nkBlSwWtoaUosP8a9BnOYE0zELvRI5XUhyOXzLf5StoZ
plwJ8izgyATP0jpNo69f8BgE3b9s2YbdYjzdN49nqGPkvIYUgo5SLHFN0+fq
HVSQyOQUiveCC6JjshypYLEuyfndniS3p2WJyhEbdOhJg2jiujVYGAN4Zxug
D0lL09VTasti436EBG6MYA4i/+Q5ELvqHYarzlVfHTs7rMBu/2BDpHomrufa
QjeJujE8iHFJP5TLE1rBFH+dzRzgUNyno9EtU7ufnDRptm5RARqpX67dlm7o
nLjP/4sYwLqzmWktHl9EGI4GRN9qCbsFzNfe3w8Ho4YdDGX4YrCer5PZ6l5s
OWNR2/SOyLDUykXXH4/aRzX84/nPY+nM3w3+4qnsno2iq1AjL74npRmq1kVV
ic7bjziZ9apydKqLIKCEeklCRtCgbyMMh+JcFgzGt3tkpVXM3qUbk2Q9RX6v
RRgkXOgOcyYISrtW5ZQ8OEVeMNZlpq6emX0uJzNdeJFg2/9osLy3lxYP0NC4
lliMYiufQsVz/xrAGoO4duakX/G3kcDBkLDJrjBIgx5mPFnzk6lvH2ZIaweQ
QLE407sPDvnv1+HfblEy19D3O1WNmoUDJxozwlbBpO56boBZG98C4bo562vk
qHmE8NXf+Cm+QUF3DvDT34teOM0GNTOA55emNUrSxpInkX1LebohaRVvM0OB
LGkJOYmXtXnh5i4fVVW+gGDjcJJQDnR+93pupUEWT8YKjjQ5R5LmHK6gb9q9
Uayo6xPBZjx/NWiQuEZ4MTPO4GbqoFZOB3aoMEJzOciPeRYmuKGCMcwxctdl
ESQWonys6mTG9nl9+Jgf9eXxbnsVYkiWXRwzuyMMbB8euRBO/EVt91GJKAxd
8AgtdO8WAg28Md2732Bh8lOgzPrKBOYnMTddwz9hYdi2BrqmiZg41d3DfdpC
kziREOJMFSazNRqrCB1XXxn3VplHqi9X8flqM2Bvw7E5lEJkGqW+Jf/qOfvI
4wEZseZgWsx1JLGYOrID4/F2CCUx62caM/ixxWjy2VrStwZX+3ZjyAqvWWyJ
YA/6uJclkqHqe1eIVtusiXcCiWvt45uNvTmkxaPPJ76sCqXv+YEuOL0ERnN2
ePMFL3p3k7H0HBw95h/Oo8kofYZ5bwA30B0WlgJnhDoXa5Ys8FwLBw96j/Ia
nWgk2ZxaUL5zd2UB2QjioELixmUVHgL0q4LmyorvL5cB3wQ/AzujIS99BjwP
we8fgvDqsJZub0mBv1Mw83Vt+4v6YutpJI74pjU9cwEQ9XnnzbMeoMJ0py7r
EnYlIFJgS6jt3afmyYo1LXAUHdqoFepRdkT1hp6k+V105604ZDGS86lCNySd
77Qsq6TwOE+V9RSlPZ5m1M62cTIzoL8DduCOPku0J8HUmBs3wWSbkgib9P2o
irgF3LJBvWk+Zv5bY4w/VP2LirFuSDUplnBuywnQCw4BbgM869ajLrFdqaPr
SLaRU/RfZ5gl5KG6ktD8ACL5Z2ZsntOYFKx6xHZrQlp+Q0+op6lpfbvLII4s
8z7gXurAMCeyBPYKixNzH43A7jqa6Qsfu8YmnRT7s52caw+Mbfgh9J5EEuV6
fXSOBxb/Fmd1tGc5zcQ+r3clsmLfaSdde1l6X/3qz0ZJb8Z/9jk/CfBaVSzw
ABTA93QFDdttpBFslEqk7Ia+AWM13hG9UBSu5h0mzAt9VFDJzPgUmmbs4zZq
fgQfE7GFDyM41ttpXWqO7PgYovUMpTxj/rAV5u9fC+WsAnuxKEQT/pUmNCvh
+AvM7GK0NWQy4koBPzzuHOLbVXTCaxdDeEAxT3RNACOGk6tk0W0+VhUuy6pY
TY+WfK8ryWXLo99AdjzoqbdQkOmiXehRj/lduyeHbQ0kpMBiv+71maXFzxSC
pbj4P7mxyL6Qp8K47XvpwJZYJPG+8bRY7pKHtCtuJpdQwyVneTvQChbTF47a
IT5yvTUFlkEnxQo+JUYH1kA04TXwhW3ni1ZgV6y0ogEc8r9RpA3HcM0fFw0v
sVS/xQxUcw4EQWksrGdJVuyFwyRGc9kRAYWnj8xgXt4y4MwToeH2AiOIXYWY
KPLZHpzunmBQFxUocl6Jk6Tuf7NtsW7Xgv3N1FFrmrPs2g5cpHT3mi1nhqmp
4tPM/B2y1jdsxzB5atbCb1QjZPx7mKSwqN7hHY2SvauWZL29xfT+i3CN1w0r
eweYEkNzJNE0azIZkyl+Op8bv2HX+sZ2w+1kpe8ENY0Ca32Orv2EOf2xV0HR
aaiZ13Z2S3aachKX285nfKldd4yWvNtCicWiX2KQ6EAfvzbwKzutofN+fLi9
xLs/gX0CuAZVrl/e4CfDf6F72Cb+DpM+28uz8+P69dBQyN/sxhgRTnKchgIr
08+2Gz+xT0Qjc7Bb0QG868y9zEncmjh+infP4kRJ79Tv8+mwR9FR7FwMI42j
Dr7fwullZqN8T+VfspW+yKQWsbdUZbFdMvqs8c3csc3bMT/HA7kawADfwaox
dBEXdndnrpJcjdMObHW3LE/WjD/2yzhhEnxhEPc2L8UaL7QAJwoxwEW2l2Fj
tGuMTHNCvJUp2IZBRrvBbhfsJiyK7sWW0mjNYHUhDIHVtv7RTJBpP1cruyKL
dcRr2N1gq6ilvat/Rm9Rb++yTq7Mx+z4ra9iJLDQvucpldxfLQyNtptY0cxF
b6YlhoDf2kMbNqV1c5GASVL2BZPuItmYiResjsPVtC7GRJF00EyHcRf0UJMs
ksgTFnGr4QBhOueNrlAxA8tcCZpcL2JVmMzfthBVWhjNkHS+sndsHXlU0gGu
g+wXyf/pE6ItREewZ/n57PUTD8JJKAUF0lD1L7x1nL6/vJ2abRE0hEKoRjSC
iW7r8+EUNdwuFFI5+0TFjstJSHDdoggSyq9iuwsRaDMot2upRjzmTxdqEhMt
0QHnrLBtJriz3fe0UkVXgUwdjrdXBjFPn6AcJlrJypgtqF8FCWq4hSjJBX2o
+u2AqLmiw2c655GzGLcTO9xf3wop2MTtgi68FTZecC7w+cOBuk8xswX7ActO
B6hmzuRbuJ+zEYb0gPwjJ4D9vTcxBOq6e5amLON/+8Mtm6oukfoXPxxPMdl5
blemwCumt8f08CFwB3S6ZvZBI9PxadWb9VJHRiHs6wQAR4zkwcPdIdVl48/+
ZkXi+v0Z1zbWYmbAmKLQOACBLw1eisujMV5UyqrAZnb+Vql3v6bnJau1mTO/
9gstwdUl+uhxh4xe8eigFWHNqvKEhPMRec6jgOdBixLhvXE25aPQEZqmme9P
UZKbkrdYflCcN8hAMB+LctgcY98YVIDPbl5I5y6JVscJpcwz+7oGNv0faGmT
uwOevMrdtIhTocjI2Z03y/NYobEZZPSymx2wlO2B8oM6rfPtGynAsm/dhtAj
mHoVfqGFnpv4OeJ+wfpP1cDiOWJOb+ur8cOnh2dXpKLaOkpWjZ+KFLg8a9/j
Klk9hNy+jKSAaQTH4d39UyoPM82xWdHtpam3xfY/jzaWg9Fy4BUBTAMOu6al
3Di6bHiEgsaBHSKAzzGa3+WtUtvPkqaUZPLdUNbj5rZkE6VoyeSd3+Jt+XHo
7KHOrRaxv0q3pat+BywyWIh8rsYVMdgA/6zMGwzaLXZoKNowXozTylirauA5
PDLeF9YJXHYwemAWDub4FY++1HlKU7ezptwym6lefd5Hb7yf3zDzNpnGyXWS
Bekn0F2ARrbyIJmYC4/uLuTAZ3UkwHrsFmL0S2/tb/Ws3VbESHuMmEQyT+0F
OeHQ6WJ0L1++MpGcmzgrb6Ff/40DRGqI2NajJLYLMp72AFYgVoBRERr0YoGl
zg1EABknMseSIvn/zCiYnSHzbu/kqAI6yfhhc6t+NODkJ9cectxuQN6bGLET
XpO2qxPCdv96QcHATIpVybPBTtl1AWvZ2Q/fxLkQft0tTIIwIK3zLgvDMxC5
1bMk4SzDa0/F9BILBirVpX/l1rqtC33LRJjwdSY6Yr7/8Ndm83MAJ/szeSNV
k0PDf93HzZOTMo3iXLFaqredUId/cJvF6ybFvxAfwVzIsJY7SElrF9DXer6o
CXStPHVaQyzd17+LC385oi4a7M74CACnT+atZFa/aJ9+THvCGZqaf0sKX4gR
fRvC+j3OOeWfWvDOtXIPS8UvHSOCX1XyuLN7i492Pn0f3txw+MrphhpBZlvL
xTUUgAyrsfF8hckFiebyYuOHS02wUTPIRFo8rsfcyH0z0ElvzPkEzorhtEI7
f5/GAUH1upfHCycUmnPOKEXnYLfE/NjyVGuAl1f+vC/DJFfNQezhE++fy6zo
76hwqzHWO+Modcmb2FhZMniMP/57MuTB/X5BSouI+vrJbMiIVS6gs/fPv0qy
uz5l0Ci7idt9VsZXmHuPA8aC9nCMGgcPyTjidzuSq1nrXOeZ2Ey62RgSqzfo
N9LTNdz6/Umn7m1rADcA/uz/R6Yg4BVhu7h6Z1QtM0NWYiySa9JjbGAFXPmy
6Tf40IjVw0ZHHlCLJPFxlGRmz+Y0ooHRw9LotC4Sw0camrUI1ObuLt/uvMQx
i3Qgf9yqaEVfsm/585zHb3PwFpS3RLcY7uv4RQZZT7IJY/ttSleOyzu+Nf7Z
DLs+HlEEAVU43oA+aMOcZP/PtcT6Ya5H3YIRHja3ZYX3dWUIqkoh+y93Cw9Q
qfV30uhQcd2Wr3uFxagQ5XVbpVMmqqdp4SLg6yEG/bChTzvQtDMnmIST6QLq
gU2p0E8uYk0lxDQftcsd0L6YGUS2W58fhirw5RE+FAyfbtlNdXx539phPqo5
ecUAgwQ1OkBPZMc2IajxSKAwnO0aW4WPdJHTH+eIGv4t3Il+7gviY6IOl3AT
NX2VxiGTcAw4oqnxC9sn6Tbm5Ik3813bwFGne42BQnjvUBWHQruoT3oTB7A9
eniEHBVeuS3Spte6U+JFr98sr08wYj9nxkmauAgH+gIACTlWg9UzyubM4+xP
qHDdEVfdWNo2aFUjV7ew24oJ8ppfhYHmlUsJzGSrFgtDe42he2LyytrFksiZ
YVo+lSHOyILHtObdX7v8WkHNL4O61FgoREGXo/Yiuj8lFp7koIbhp5lPp2jj
GcJ91EH/DNyPqXmjbMyRvI0dK7bFAzyKJArOYpIE9dkboOP1HfBfzISTK5I4
IP6cCC8jHGKswfoxSH5xsPZ8cj9ECyopjWWex5zt/6BdpdAqWg6CUPbinnPb
pycnlW7y4/SrS2x1DN2lnSxRGtEERpXxRhCqVjrPz13DQ1HEXo8ywLeG/+Iu
9lU4NHmmH3B1v7YjqteDpmufApQ2X+cVkpVeh2VC2SHaEPv/SRifaEO+Rcrk
1ucXmf+kY26cDuF1H7ghU5pFwRe1tRZ1Rk9o/ydl2hH0ga+HL48WHkPjDaS6
ngNRGvo5CDQrwXx00pWAG8V3eSI85pjrB2+CRFcq1br2T1FqBI/f1v2uId2V
+d56JiLz6bFUJ6h2IXcWiX7zG0GppkgYXSLSZARNZt6NHtH5JW6ro1nCJA10
WIKEUTetCLmXFJc0bKBjVUcK4+n1BXVxVz8T3wono8eMahXszb6DX+LtU4n7
BlyCqHNJlspyisjmH5QB4YJHFuZ8laj8TiwQb5VrTTf/2x7o5QbeK5ekrMlk
OdNrWEmwKQo7D28ihryMKQD+H4d6F4eQYEcvZs/ck08MyuU4KRtXZt+AvhE6
rJiwXuxYR5UzkCg4D1IhLv8U+lyCagaTT6JwecTRszT/qrd8GfSV+gCx7gbe
YZUqm53g7j0/oglggvDLf+O2d+CaN0hGIJHncImG53/HeWvJo6JLwMrhh98a
NV2VcYUwGkHgTK/ks7FEAx4noj+73o/ornjgfO+5+MCASmBMeKGBdvVSUPQG
wjVuZBi5Jq+fDtrL5D3J2xLQfWO3EB+s4SXx+u0FJfAQwrj/2fbOa0CCX2cX
euobrXhmjzXhNPKrCkrOrzcY2XzbTSGAFFIG74AldjLgqM7g17/0cMZcfUEx
klwUOefz7jF+iF5yni4bUp80s0gWbMyN4FZU4ub32VB0Vco6NNTTDJaOQhbo
bBzMLVJK2A07FXaYJgTyFlIjRSKx+AIZdm6C1pxQgLACvnoMq14ZsGGB97Vn
hNNVwDFrAFpIuAGhNvU3a+0cWnkbLpmdOjzOz5nv8KSHYz03jTA/Dy2R/2fs
Tq6Li9Ff2WwgKrYfQZqs+sMFa7/hqxUGYp/yrHohPVhPQBsSdW4yjG7G816N
8EjYy4AOLcwfbVGGHOVonUSCS/eIH4kxSAMMdYgr22z3/Bg1Bb210IAci2sF
22PJeVSmNYGlG4VlSNsN00hfmfRMCthdsD+gfFdsKL7f04PNcib22UmlW+B9
i4etz+lTCJM+aG2yUTLBAZ+PwniVSHHEp+hFLirC+H0Zp4iMsoCD4u/9S/UO
0VqRIWw0NJw2H7hA8uLJpDfXzt51XRbQkHhTgYLnePR5/6CH8t3Epj9sTwWy
zYuF1T+PQEhY3EdpVjikyI7vqaItGW37Lx1c2ypuuQ14uqyKqxovYyUCF4iq
VHgl7Xbidd6zo/JY98QHyH/5pIn7PmeC8b+XoI0caPNS99YfAtbzQvb6KV3Y
ph164Telll3lEJcmJDWeoyNyXsEV161jwyhDpzWFXJemYDN+DV/CSCiydyBK
ZDiX8HgS6jpxFe509AS6f7WeWtUGToLoA8kS5+v2TsjaJZEcvOcc7J2r4d7o
u9WlmMXIcN4H9gPyTz8YcJnnpXSr8c9B3tRJoNMfNeB8Zh3H39sfoMgMz4CP
swOdcI8O66Ck2nKcjdYzCT25MIHOpfKRzbvzQPu8lUi8i+GfDqxzpldC6vA2
3ld7+UhGtyChAoh5VSLnmZdHmGlTs94NhN9d23IA1LAHJ6dHG/k9crNoV3Pf
V1uzN4SvIS0WDqMMWQnB0LerQCzQBGOalRWvrusTlIvJYNB7NhZbovmfBFi9
zwnzeTq6x/SjLHcgyqT7D7eLL6Lhd/uxF3MWtmEhdRRRMQng/67BzROV5rVT
HJxYj8RUxUPd1nGbLDwbt/aFbL5BnfxwgOtfn4dljpZX6ZPdm4tWChVtvvkC
txd4TLPhNAd0hyq7sj8acTFxX3my2RPXADlCZFU1XmG/TUxBmz2pfF84eAtM
m8B4yT1XsUzxlMpoYUNidCSg0Nl5Pl519G7jbQJolTk07qEqlvilItZ7ZvBq
83sO+3T9PY1ZZHVZvDoATYtCFAFPTR5LTdh/5F8LBjAKu6Db2JoNrz9XNI10
O4LZrCAL4RCh5YpEnJN60abNRexRiFVaKTVw/6rv63975Oxb4KHJc921/rak
scYImWdRdLwtwUj943wcVkQ1t8VsJOvzM6+dia/6LuWfEqWAwzEKp+BzTvh7
TeN5eXR0wd6gtCL4yjWsLPUEugLXReOfZjDxtQrP7GA8AjjTdeuHPZuD57lJ
DUoNv12ObLtDG6jYbFNV2U7wpz53Wg6b6QROfrOFEhgOIJOMG1XBv0bA2j+V
S/K6J2Yire6OjBHZZIS+QOb6RgyZNXaxaeoJ7Yyebgy10mAZT5CYkRZEyRI5
kPGmD6EpKo+QL5FbAh8Rl1yV24mb/25ksom+pgy4tio5LHJnp4iePHU5cqb3
RJg6uxZewKGCcz/yTlCBCfAre1RNgNygFHRIfZX/9xACvqhO95RZpo4kD8zW
lHY9luxca7PICzSfwpn1fCemhm2FJEjZRnI+l4gX7+w6MZoQcun1/a8izbs5
0cgAhPVcxqXOcda4VCONoAFxcX4VkV7Iz1DKb3TlON+kv+Gd6FCrvbC8+7iJ
NAAOAmuNNX11ZrfymV8ocUb7RL5Z58qUMamA2K1BkcHA6657OmMoR1SM9qrw
PtHISB53Vwvz7ZHCgOHjPsp1kQJ7w6vrO/oMe7fqyh3CjOs6B4AiXmh05Vgt
OmKOVxI590Xqw49Yac64us5i+LMJcH4NRplAH39lBBy09KqAlC7Q5dwGUf0S
1i/NnWz0l4dyMWmLsBxUV27AGRR8lRRYMumHB5X2oZxaFMy7T4B72G8nm82+
xUiSEAyYrBX2CYzoQA35fMZ3NBCJo0MgUzY525QckmxiMtONCOpO/J8qESZH
zILaE4WsONVmTZEsGbFOa+Vm12hXEdX6AYieBqDa9knmuhOtrzUcfzVzTfkg
CgfJ1D/cSE4xjIy5XZbtV1hD0r8C1M20jY4yhmTQgBEJeumqSUmuJWpIQNxL
/9Lh3g/O/4HSj6qZ0woHjYiCHM5aJtPgmttide0qxS2QpYdtIjlfJgfZ+Qg/
PraCMNtaQHsUzK0AvBVWDS2c24jDJb8IuXpBSWjDn8rv5R+gu9123m27TVFA
LLg44G+jrX4qHlW39zkWskVoyfc8d6CbK2oGwpEOrmzO+sA+0PAOjYWqfips
PrWhoSZlAxvtcTU2DUoyuZ+7yQ/0M4z8586iwG5AP/LHSJ1e4rytL8GQDecP
qwpQI+pAtpOjD/eqlGyKOlIn3Kd5zDsPjLhaId0lTuZBriHsEmoZ5LErF3SR
YfyQMUBBk5MtzIo8IA6fg7AmFLG25kmezXzBPEKrIBGvWiEJwI+NycWN9Q3L
kmK8uzzyKsViyCKxye45FS0DKdulnnX+Yier6/U1QRA/Z/Rg85undQSuIQ5G
tFKg6Dk1iB5J/5SjDLIedf8wqGHtgYUYeD0sOSgGRBfVcVgYh8jc4szJqqAo
cOZ5R6JvsUg0g+c1H1qlv0RdoUIsKrHSmkhGv+mN5SO91P807TVLY+Tzt3ok
zIgxUq/lOM++Hy9XPi7pIXLlxG76EN2haE+8P2J6F2MY5xtcAQQlUI1jnfaa
NRygC6Zdt5T/Ha6TMZmmK44dUzPGOEoYqiMUyg53pZTMF3Iwx3gbio0t+haU
V/T78+7vW/H0+P4SKYQ3VdD+BMYC2BilFeMg2gv7uKNso0C2Q2wtIT7GL/mP
VB9lhy4aIS2UUr+A5zvqQH0wIs7EpcuZm2+9fLHcu7tuBgxn0kD0fo6AUAN6
iKpqsr59fdkGIJPqPxr92YfZn0LGKptl+BWL/CqDUuOnIK6f6YcgktYIu8s5
OwfrzQqNzI4VgYgcSe7pJFbRGUJZotJXgUeeSvfpegxcqg7hGN9aREa/UIrW
cQ9YAjA1nyXGU8dRR9zMUE8mXkOsDKIuk/RqT4HNQBm9anBfB1gq9tKX+czJ
eWUlb8dqfLyk5klsivsyj+rwwlZ/ohTB79n0K7NQADoYWjg/gFGWUYhbKYcl
jfNKKJLsUJDa97lJrB/lHmYkEVvHrzszuTEaDdVQYKO2L12AcAd8rGYXK7dY
ZCxtUvCwRvb8cTwWr49ncjun/XjgOldjW7Ldy9Wx6t51gcRhy8YB74bP8SFZ
sw04EKdWdUD/sIYNIpKnBQOJ38SHV9iOYWc+uBv0nbulUr/Srl3Aroa7hrnk
VblxfRnmopdcbcFXJCru0kDiQGcGZOuGdVkhGU0qEx8iJIb5OVpgnj8PNsx3
ipBkBmAHPH2yN1vprDWjuoW44wEqyI12V9WvB2woZfyii0REBTbb2VW6D4jH
qqdRLOQL63jKhKKpbwLLcD20TCZx1NH+BznhecUq/TyO6CkC1lM14sUSIPdS
+VN4IDNivCS1xd/naC20l6Y0+8d0hFW2E0+YFfo2VibhAO6AvHexupF+ZKpw
RMvEVGnIBb/us1VgXTRZclyP2+mlWm32vR7V/D9YxGI3tKIpRFYK8AEo+yqj
YSAth/6ODaX6H2a9U4HmG3Hk2Wkk0feY/leVE5K0dMnhUtDZlJvup/GV/vvZ
ZilMcS5RjNp4RSXChFKcT2UfjLLNRUUKzy73oLlFQwiRDSd8Z72a2853jJxI
ZLrjY41cxIqTTwAlrVoCZSOISwW6sTgKIL1uH3tUrAqu3jLXN5BGnTy9+eRY
oLufwvGExwhcT4NGSTNaGonw2MOqM7EZl4XbqBG+ogcKklB/iRK19YJrgJmS
/+2wdx9mDY9ZQ7rs/aXhLaIzgOZvtX0FTmWdOU8qXUAp8ggU8ltqbwW1ZM9E
+SNnVekG1ZibQYH9N/+zzqm8w93C8/Vp2EaqozXPNIgDnBVNln8rFq8FGkmy
QAlcYAwbKNA+amqi3LrpP25qwT/NkO8OlOu5LywxytsRVwjo1uqnV7n3kiEM
6GcO52ExTxn/c3mKOhsF2Jj1cSC9sWQXS0F691HtOPmyYig6M12B80frqrqo
cHJp+mKf6QdASv3S/FOEfQ9kKWHzx8WsbuQdG9iSkAz9tuJh9kkP1jdP0Upo
84vv1vaxNoSd+At3jal70PeEiJjSSEk05zLealwczVA3JNTpYLKQzGyCclCv
K2IMLTcZyTciuUa2+F5j6Qr0JIXhF1g+uyWi/7glDb3chVVOs936TNX153s5
RGTqVYg3/UcOlop5GrgHnplh3ekEbhIa9OZjukJsTUcv9nzHZoamqRW2Va9z
HwZG34pRmmTwVHiie1jJSAFqEFmi58VGdvAd1JGmS6MUJcUbMI5BwtRZjm8N
vRqy9QiT4eh5E6UxmOyH03rDdLo+MkKafFxLvaVaoCkR4nCHAssBLy2tMQNb
iEVK2x/nQ44tnKzaws4CucdQQqt5dkj2XDL3F5BBl00brkq1vTtvuFES9ndt
Ljshmi0RZQaW4YTAzB7o4D8CIbA2cen1TpEs2oC90J3P04IQKLFtL6lAeJSC
LHgUhG/fuVgvlLVne3oypuPQ11tBH/K9T1VfU+Dl1SnGnQrm2KUHp/wg5oqT
i/Ux6vwemTzZ/maAAakWA/5pk8uLAJsbA58cuMVGwokBU/8mIo0zwllQowtc
WgPfOGulKGIUPgs6uwkiNgUMEyj93k0227t9Eg31xuaard/BTQDXHv6Yoqf4
1ma2UN2ubR1TyYzhKRdKCYYZWhzql7c77M9NSu5BdNWqwEA8k0SE9kvBtX8r
zZW+4pomSSpF83Qb2N1fckwCF7IJmtsaN60jqCxFIn6DMjezG7has7KrsmMN
KKbMIH3QXmwwSy2alPcuJ06FjjTqMmwkcqfOaWEv88W20uFy9gFOUtWWv8te
OO5R+Z23x0brsQqnkqzD8eOs69kn7pfxAz7lUH0TsICKrf8OzG1OGqN9yM/E
sUtupml7K1HXP5LLjrruTg4xWnhPJ4C9ILN2sY+dM08xImj/glmu45+0YEXg
21Q1PL8yVtyS74Bkl7rMe8yu0ZjiNzbvt1jE8P4RkzHAxThUfPxwQq2tINRD
QT4nE9f6B2fgRah0kC4JhbXQ/9k0FeC7r6eGcwn0M+Tkr1aVngmeWfU6aumF
nysBklpxtyfLhGBL+q/oS/dRXY1pHdL9832W5HnnsWn4ycK06f79bIQ9C075
r8cw3BORF5lvwpRt9/I8kOzIRzCaUmkdVgfEW+fI0bmLRyo+Ec6mhJde7x6x
OEN8HKmabdHXIwTep4pzVJwv3BDZ6DDIWST65W10sNbp1ZLA4GgHKPMv/VWG
JEJEQXo5GVGxZibeUMXzltN7AXII2OWlQl8qSR5zawYPx9pb1IfVu0IqP+nK
Ab5scrRrCfsyIJwYqHc/wIOjfNkyA/LoCbEqXcN2EI0O1bkVEXx5URQ4AXDJ
P6hBUGU8nWCeTDxEdSy0/sHZtpdnuKkJPmo/TKHZBn2QgIKYfvHuSrPk8r0O
Ja4RTe9cz+Y36I4d/ll3u4zbRQqa50CzVKZoAOblIQBtuLLUU9kBIxfSPfWk
/8JI+ksdc5nMt0AgH0M5DIgP+8VN8iuJ48znpTjdiGmYjuK0DCULhx2vynnv
QYvMw4OISi+UwhhE1sbLRJf5vIlUsrjfKzE3i/zEYUKawF/wS+wiqVmt3VmU
PDrlzWXbH6hgkEtoGJ9wuPtBCs18/i7WNe8hhHitwiZhNO7OZo/VGrzzEv68
nuanMGdlYyQ7lg8gsABtsSXfbUN8Ir6VdFyd2to5AOw3+QF7WCFBiIDhDFJ1
HtxHa6+php0G0IIlUSLHDfF1FFyo4uYkuE1IHwmGaJaxCKyTgcQnj/VDtA3i
Z6xw1Y4J6FGCnAfCggoQ/hSjwkRnAAE2DAIenYbtKKvl2ksMSsLM2OsH36am
gpRyz1Nk8hNh735ESwW07SIx960ZU5kJR2g4/M4/P4EPBDmETSl+BZnXByHv
pAKhiw6Zl6/CXUF8zB0HP7abwkTC/eM4uE0JndPOAOZtx0RkZH5EWm8leqnL
9Rz04UeUn+++VfFjAXplDkd5RjCEq3bvrIxjH9h0Rkc5MuKCN6yiud0XU14K
tBXZpZPhMNYqbm/hx/C8uMwZ+GmgSCzwA/ofGwOXVb2B11IVdDMb55eq6VGe
OmaRKlBDvVph8lw/1I0amCO0b2XJmi8C1lBJ7K80dLz6y4h1/Jzatp3iodD4
Z6w5n7mdLKwiKyGFdJgcWFa8/ONUQ2bCL0Mvu+40UwFMNvwgN5lbtMJFbcOv
eO3bApqvUPP/pawRyhysRCpjviFLLy18cyf4GAuw5vqilTe211VelSpv9eT1
cj9OXFuBIto8+LUxsgw4WJ0NDpQLn3P3T/RK6Dq6YjQt2lMapumfQDfLseGa
N1CQBoNICMgE1yGHgwHJrlD3gBgQKSKGIykaM2AxEbGOrYDBUCWVTTrZIQm0
Obyxe9gcq/0+kdk7KLddfoBAlJD7o08bYpcV+NOQDSoSVfnT5JJ3iO1ZvBC4
f+lk2vXn6cmbZXdCyqVAJTNIC7SZq330R7pCwyVTXc9IvAl/BfjiJV7n3FXp
LLMaN+Ajqo6hPvKf+9ra3z+8PVM6G0hLwlGCTUMbTag5YT6Exny/jVVxUhRY
yhylmFGZnF+V/a7UImPCdDLk/TFs2oBYeZJHDIaIGpeMoVNlTz+V38A6irr6
Wpo5CwHGG65LSk6EubpMLr8s3UXC/Ib8uJMzoOCeSkHE9nHWQ7q6PV8+tofX
gHOexBF1tutijyl1GKoKWZgHbdE0/Oiv23yGibQUv8b20uho+mwzUdKsaHI/
wT9OFblL97VXIzkd2/UtwAwK7eiETc1nKTFCGv1FO3Srh0OhCgD/+Ok0Ahok
0pEFPVb/zazYwzMynxtcNof7eFMNF7WTmpOaNhBGImB0v4yrLm2dG0KG6Hin
SQyRFpg2z/n9EYw9JyfzrJ9Fdq5sa96Xl9BbOaAHWBIZnBbaAInLjs+my9i0
mfnw096Cyy8MQ1e2cWcC9p2RJ2z6twOJ9Tzw6GmHvmonL/a7ZzRMdU3SJ/hi
inKjk2WUFJ1y8q+7XX9arDceK4J7toQ/pCwUdsn1K2a91kDULBghlJYLNoWI
oAaQwQCEHNqVz2/nVMqKLjam4Hvru8lBgdhpjM3DpT5ja0SUp9V9wHvwjDHj
KxuzE/sg9rwnrRYxU0sQNT6+LhyI3SGypjQmOzeZF4IVpRuznN7oHhs2zimw
hVHHQRGUWZrkBllGGvDuInGlN4kStw4qk8EVSp/htcxluWiH4jCqGSe3rGAt
fhbWbRlqY8XdLMMXhveWy5owb9ST4kaKSumhFC8/pZZmRkK+Ip2AmvbiMxEx
g0NRaKsqQGb84FC8YIRqlc5qbnoPtKcRWd2HJ0haC/I7HpHrzV1WpSK1vbD1
ECFARYi6a6BjEvWuAXtM+zxNyAeEuh7ayxSBHgwKNlgH5lXttangj+/HxjQu
Mp90yMsdhmsrLmA/862wKdALKfwyxePYTjygOAIAbbN6egj8pvm8jK1AzeFZ
uNNIQNY2Zi5CNckvmH71n0+RI+n1ON8yP0OLHngn5DUcWJHEsRwD/Uho1Hip
jtHI5cRxqpU7/TGNsykAkNPKqicW3n8v1+ucoZ9jGbKjw9hfp8zcJ5sKX4QI
kl4PhQV3kFaFJbaptq/a/NWYMy3q/rSLWRveofhMP9bN2f68J7jWUpErSu8i
tV2exNZHmoj/Wcp2oIoCVMNIvRUFbQZT59wDJ28z3j6u1tjeh6NOJeJlWhx0
GUyI7SPHUPIAw5zUVqGbaOSOpOkjTnNQT8RZ3tnlyaMZGUeO1bQGmMBHNYnd
yOKOz978upsZIvTUOfl0MfEL1WmYWYJzjTuI42jORd4TBeWwqSLwQpyHVsKU
tPB03CiP4H4Q1GhKQfkZZkmaI464pvHCsP8olmWNeqaiZphQ0xS7I8iqluCI
D6ps6lh4zLCPl7RARXOzeiIrBVPUonZkeDGYPidZQJEWBKNCOLM7ZtubYNl6
xaQC/O9WkdZkU5ts5KjE4wDfeqkWES8lN4JfYCfphNTiu3WEFSOjdrM5+FfF
wa23O94/R0Ot0GiH9usup2UxF4NGfr+zCwqJMYQ8+A4zJg2CAJ/8T673sRGw
C1tqcflfFLAY6ogSuhE5nZ+nOQciJfJmDuSVbP46V0B97Xjxt2YcqISdkkeN
6DgihjV3Ccx7o6yxClMdbKkvc+0qrUM4FuZYbekuOrRXbc2gsmkL47BY6D5V
c8yTUtVLXfXRF9wt2bymht8ViTJUcju8opWvu0poGDPdfyRSgidNq4yZsCpZ
BuSd7FxhWmUAbLfDPEP0Mrn4Mvq2HPtjWQf9nDPvU7qfcjJWFMwyfPlHfc7k
/BU7qhWApUyFOUH2eqvthkpZs9vHLZt+NlnVoRh3ocolcMp59K2529mWEdPI
rva0Aj+qjyMeCXcmw/hLun+1PxPy1jxxQTnq+3q5KYfm6iZDCPclydqLxv0x
XfelDljM37sDqbzJp9Q1bnaELbYwk3GWVQOoCR6+Xnf+nmxinwmAm0ghHMdJ
9cAhDDE4UGMugivRreZCSRlVCaYI7CbmHZ7/cmlSG0QcMuBJTjDdufe2Cx//
rTVJ89opqX6I7Y/jHKEVJ2iZMVONR2kjwqeLtADkpQzMbt65O1nnB1ti2Oby
uxE61q9SjKNm646mbgJelM2SX9/Wsa68KmSQ6TAqMnOx7Xt/UnzLqgHCdWoj
p5ZFjJcR6pP1Tbw3Ch0OzVRbCHnu8Hvk5ihS/g/5w1Iyzsq2VBqjKn3UaNBe
VVOYa8K65q9L0US7bsP0fJlPpx2Sng5gYEdtmWfy5TOKFfQyyGFF47EIMeRx
RRvrUPPB+0UFjrCRwiJRBIF7Hz5izxELKngNK4hZIwLAqfZB0hy5YdcH/yDG
X5+5vZz1Vb/pKnVTqeDLp/IAyq9YzKi54AFzE8nypQZ5TFmx2VpTYZ+qJzCV
3LE8tsPKMjfZejVdL670wvrrNf52+CaCmRBTeG+PRsGrfAT6ejEF5aYCFrvr
4RjItNF77wdOG5FPepZFl5opVAMa1Zu5dAIhay5jGDRkMngBtt/Eu0tAkuLg
sCVHuAq4wpXQJBhLPZrAdGYdK58sKyhvsdZbzLiM+q5dWY0WDSLVjYxl5kaY
ssI+G+Mwbb7GRdpRTwgkmy/N5Pifk/qgL/j5fS0kAT0j4QQNtl12J8d1sQ8L
twDdh3fsnSod96WC/ktJ7TVPwZqUGoztkJusBpJ+wab5H6OxaDFRpPmmJGen
6N3ylOWYTyNdAT4nhzbpmt/7PoR0trauFzSODcb8UtXCMp1ZrJ1Tz4ZNjje3
czDC1h80dxKTS4FQ8PnsntXUiYjUmjJb+uuFtnk3yNY80L3Wqyxqy2/uwqYv
2Y11QRkFUkPW4oY5is2d2ZkN5U+xLkgEUDxPX3x7qIJ5ngPY5E52SyEFTpEq
z8F7In8ZEaJgaNjd0455tQboFnkNnT2xvQRf9678PRPKcc+oGCKebnNVNgP1
ex0ZLHCylQtp3N8uh3MVgnJmrJcN72oMzPm4be8ZAH2Hyb99BiXGBhbMbxhY
YvK+UzOT6O49pD+EUwmv16EHVFowB98UPJnGHLCO2tjjOa4/PEPbFZCKKJbu
740JpfGeaROWetkFeFOf830O7AoqIYUdPniVFxqg9YruUWBpFg9orziegyY3
8+6uYuHmcrlzJzD6rz3ENe+rJVnoBkTDYqyoc7DYCVe4luYJXVRBOvxea2hm
xhg5BI6GLBom01Jx2KINSrgCeAisUkfiZ0AVplkmpiNumH/p5TBldCRACsrX
6Z0ZbKpW3IGJhUCG0ti6I5AQyq2lbqFfr9NikalSfP2rwVIg/rYXm0HFsnCl
TgTYjxWFGtkw1nk3joa79tnzZ1ET4VZzRCh6lV/Jti3oRKB2uJOiBWaEMPsi
2M+6KRtmEUxA6xGU3rPA2ByX38OV3trlGHjBKfgQfO79ki9Z3bFje23Mkzq6
N1JXoN/e6A2kxs/TPdbl8pCuFY4honaA6edJMqFSXXJkMiv+HIrYjkg1t/wP
aXdzCMhI836igAhBw3E9CLZsXQDh+DZn4I1z4hR3jaqzDwPiBRgycjVZ3pOR
ptw3oK10j9Z7ynxrf84E0M+hppHYUjDfr9/PnMAU087tgHGzpRTqEHHbNcMF
gM2u32fEpOidBPy4MDzk3iTFOUwh0lt7GwUuKnSDivZ456SFaiKVExh5xvly
AlOeOOssKKMejQYq2S0zXzUqEtxsA6Da8punUAqXvWPfXgb+4NLdglb6TIY7
63KHit7ajhsmuPZhZ10461NEKeMUGyDopIsWOD4oDbS21IJ7teppI2m/sTur
ZsFurlMwdwgtvFfg0j0PET2tsAWN2tNcZxnh9E8JwJdhouknQbDhb5SgzizU
nABrQVBFF+kVjIyS67UFqJ8cC/u3GAKaPaLb5yOp/OOL6zh7UerOssHisPO7
Y8wZXF/FYh5CN3HISyBzzwM56pnjsNY8uGU+a+MVAdBJdxkeAMcd/4dcgKT1
npIM746lU0swvaILUZQ7GOM0bdUShknaMhJSrbb32ctXiWVxYRyOM9J+LIAi
DWXrl8lQiLV95ovd7ju9sjdPKW5nKhtrRCAnHLJuCQLJiKIEC/r5r2gVUWUt
rzcmi0h3dtbEqQPVIYfyBoBQ5IYG1Hk7BCoer/ty9vqlop5dAEeORXb7ulry
Cvz4qmV/Qq+08M3pweibmXnrlmsKgJkAqoGhWic3ONCvTUWegx98JyRuDr7g
xsxQV8Dl9f/vjjW/U5sT+zvtDSCpChar5uzYtXSivrTomdMj3ta4ihB4Guwu
zzmJn9jZ9cXn2+5piVfOmurreW8nCoQCikC+y3PItnMO/pRZUQy1+r12qIK5
zBeiaA38KTcaGGYzYNuRe45/fJA/NuNXVCMSd6Kq62xWT9ueQflvG6kuMRn0
folRdb7x2m04Sg419kbB0MAPy1hmkzbblHVudi1Gm8RPqLGiML9OSlriTkbn
ISWQHx7c5mg7e2y3X+GFib6663UJvgtbd/ApDXK/599RLzHuv7v5zyAO1KMf
pQhthSAPB4C42/A6j8QgeDb7ItTyoa+vIX/KrQs+u53w2un724NplGhAKyeo
cFzi8HBljCHty4jBFyOOItP4lOLWDVzWcxChsKPbcL6G1tef/P8fzIbyNu93
TEogXjLZ5fSPwD43taX52niViSpcF4x3PmtZ/VDPjC0bZuMIrb1Oa8LC8rny
JJEB4Z37/99mio4md++jZcqjfVHi046+xOdirBdn7wGRzBF0Rialmj/8hvRt
+oCy6pHHp2ukRaFLM47XBltciO58kii7Bt3Crg+bP8OJDFFvlfhnipRrYdmF
HtGsLRTERTa+8FJ7qdD7caQPuNWkTlgAfrGpYGdceH6+uVvdr6IB9LHKxLL3
105Y/6GmGitM2DyOyUUQ280MJuneZ4GdQmh18sv4nqeHNQl+b8pgUWSn4snd
C9hC59rRMIiFHAZz22gka8BIPWE26aNDI13Pw1C4dirZ+hbWsIGl/3q2/RTq
tDU8pymyV6XQxwP30bivVsCxjnDS8J1oydNXgU6HndJZUi7rAOw+PBqh/OAN
Zz/RF5tcSwGGzIJP4tE9lMT2XMcMrAtOKZURlANpa6ocF6cOXag7A4acB6EV
N5lLqQ+jCU+GlBNazVH4mHojzCrO4nIBOYymsHq9FQvJujwusANy1qlvViG0
qQFWjBhuzCy51LoQXDKzhUqG9lD7LDVMV34Edw9sIeefcwdSj1kQlbbvTY5z
Fi10CBo0dK8fIM4/hrIiEdPLwFrHuGy6kxQZaz36BfI//uj+RUjYIOUCnb9M
bqQYJlnAm+bdUmJOULUZTiTYwpoESRv4W4t8Uq7/5DxaDUU2DLglk+FTu14j
MnTIF8LoGlObrm6FHop66JTLm7HHKo6DfrS6oA94GihVmXgQ6EkmE4yzX5PY
9eU2c6fMHpahkX3vWqqBZ6tl90JZrVwAvnSPf9wdMFaBWEfoWFRg8+ZscaBx
3UzAKZQWulUUOGd1ZA/LhfauUUio/FBfV2xgWLCnEArhC1z//j8T+eO5GcTL
J0ufpCiYChh6dPl0BIjhHth6SSWR4XGunFqMOBvTqjhavmzQIVOCet6ubvy/
vGyaaWTeEt4F452nmW83XdOTGiPefb3rjQUlQKVKUJW9TknkO2iH+Kxes+4M
pK62hO1RO9lkT4TChrthEbbh7v7Fc9VLJ0Wq1J0IKgeRMCa5iYFrKDqvKWUN
PpH9OsgwRn+hdzgfPhs0LlmVmDv8VP71W6sCP5R4Y5ElBtWkUbP+pjUrkzGu
LHg1uWzl7nr2N7F3x4lD2sYuKx8UVklyI+xKTXUwhYeF1JkL8TQkJ+kXVXFQ
UVTWa3IqXP93oLCDtifRpZ1JLJJSEFiFBi1KIV+pvpdqzYjF0s7pPm9OQK+v
uFuASC/GBR4yCOYPQAxYqtk2qFGhDPGUvpYhpZ9+Uub6SheckQbzlU3pz9sn
JTcL0v44GVrUa5E7xUEzhcWdCbaNP1Z0W3VJBeZUKeZgFTKDmaK4j+vQRKbI
JOJiEeM5zgBKjCcI0cQ1pQrEOYbhIqMvSOUQxldmnIJj3XM/UhZ80yMrrLmb
hy5LwpTTciv8+vkazw0cExukFHfHmd4hUu4onzE8Mdq/NlrkKKe3zWd/VOx1
I8mcBHLnDsw+drxA13mP23UD3ezIcLQxxoN2EzpZxCsL8Ur/OEo6ikMZm3O7
fUS2kKiK0RVjVYdiu/d1X6ra8bTHHAlCtnUF3pJ8U6W33sCnsFSpNXD6aUXM
+EGBQOg0hA7xsj4flOYPdA711K5dsvOtUE5xA7OfJOfs/M4nEDf+4ofaKLMy
wsQwbcGrot7Aik3O4K8cOjXtiOh/LQSbJHCS3VhEmnt0zvNNH24XUgwIycOP
+f+OyL6kRYGok8yaZ8WnYXD1j0Ms/iiT9jlJA5YwB00dJpRgaLQsFNiypHqh
APpGuv+SOHiTunjox4BjuisoVsndNHSkl9k7oRYUGsO/sSmCM+CxWySUElQW
d2OnepBSkM+O/FBIPbQ/uo+F2OEwqs6ZTWZEueGrh5qHLO3qn2ervSV0ifX4
Tp9dGrv6BaOTJsDdxKnYMs1Rkv7XesywpYtMNB5TJ6lURU2TVGEWWHyVdzg/
f+u8BpRBN2iTBUbFp7mwRSkM26LP+tZhV08j/kH9yoUNQDF/IMZx/csFsOqF
aqFTAxuWCW/TOMWXX/67X7FAEfWNX/h4SqInLWnbb/mNRHJpiNsV6/iKRzQD
3A+donEhwT6MLe+4U0WKoxGUqy/0aaXEauqWj7MRzAJAjPA0TR/yHsVg42/R
kktf5vUHDo2c3FRc6fGLN/GaaSNqisG/vCvXfzTF7oqQZA2NXJXaIL9HvIM+
ywbF2tBNwzSECjbWpqBq8Wxo98PX+xdkuVs67p8cLZlyhp/fHxvbo5FUOCO2
EWnQvYhVcMvzdO1FBUgzmdOi2Wr+Smpv0Pc2m3Td97GXnudPHJjNpGH6ehZ2
ydQRiQ/i9S3Fyx16QPTTA8jnhbXf1UBmrbAeZ4j5dy0a8p3eY4udDqVoJR8w
P5liptkUzyZ+BEa4icLTV+ANGjHgxUD+9rEBUAGR7XSiD7eXH8XmHsLGHw+c
6ASy8J5cyFhmR+KPsG5zrweFvqdQFXkcM8MStns3rvjm47G4Il2Q3DEX8+EC
2RTcKJLo9kPw2JKDGyrbqvabkqPEuZAaDuiRJxBEkbCk1S+A67O1MKeQDYcK
tGsmvHv9YQDv5csb5/F9NVYu7OXvfgb6YBzY802LkGPXWflCcdLlHllSJ0IL
z7t0wZAdPuuk/B7qNuJnRmMgBQTE75k5Jj6GDmVC6c/TT8soD1c7jI2jHR/R
oNb1K950C+4ysQloJ9A1oDo1jDM3OiHA5f7EY5foWfXHyGDNDGYqXoUOlw9G
tdSSDBb8ssd/bsmbmnyhNNn8RkfyIq3AgCzYuXGCzaBdpqzU1MV9sLJB6Tg4
lw4qWr0DyxO/NANf2IsxrlnDxWvgvvNXTm3x4xCJL18msuLS2OJ60CGdqnc/
8nC/TSjxX2QJ+58tpERXiZUFNwlvBAuLYCvdL0TtkgVwFZa73CEhhWSa5CDl
OSv/VjvhT3i18Y2YB2IlzlczwHp4Q1Hkz7zGJ+HBH/UzzPcNl6ldFUbACSHz
uAK7W4fS+J15cMTaRsjJBK3FUQyFO6bGIPhaBfSHETnKY8yzRGy3EeM7398x
ucqDawhJMa8uXo7YBNQh1IslFScYjMD4exal76Hg0qbFgyZ4QHFbmME5aRIZ
eKt7jO+/MVZIf0DFsy0VAJl5IppJjmFtfPRfwqF5jpfh5wNgLM74EaPuOsEY
SHR0vWRHkWPCBSIwM4I17zh+JQZ5z2G5EMIwx9VgO+2bVlIUuju/MqsfK+aa
9qI84VoTI88KeZI63Uuu7H4BmNvIwsvZ/3sdCsPPbMP+dyl1Mb+U9A5aGqOb
ptt4qGbB/a4AxSro5FlbODZHmTFrzjHCwPO1IdGgMDWtLYAsFgWAI2EAgnBc
5d5y9hTVJYaYbzep0m2R4spMTHap9/RwhNm+LY7A2OwAwwGDhEvOEgOzqpds
zJSdh3llkcZLNdtRLQg2eF//qEinxPvYPGo3p7hAogB7tdkoEY/i6v0czcQR
7PtPyvPNkQVUmpQk3GwnrbtgOEJ2ZI6YIFzGWNtCjtLjJmysRtZdExEfSAk+
IwghRUUC1FYL5LfqHeviPlojZbqy1voEg5ENKiX3JtgLW/E3MRWkihzcX4pI
RoTcxfN5NRtVDkpKpSGk8DpV9Y8kLPSZIX5khT1dX2SXkYBqU2jJrPsPIHJy
h+ZPqeXm2uhWQiFP2hMirvfKgqa+S8IU8boItIDNuLlvVtyFsxHWUQshUL4p
5k3ujwpnrVhB/8Q6jOZwr16gshkeKHMUk9scGeo8eXSnug53b/llgU+GmSi0
uS1pH9lYbQtkVaFkQ2nbnTqOOVCyFMzPPE8eCSDdvIEbFlIUV9AeXgymTjz7
CdfkLjyPJr2T6WWTL4XebI21hmMAgT8fyMSVEHsKXhjNSnV549QzBm3iSwMI
k6rsaarEzrLPoTYm3G+Gs84eihOIfknmIMM6w6cW/9ou2cbCJEg7AWdKOdVx
0lDyOM+yFWgRb8Tq/4c19NGO1tyEQg0d0WsasS9KxLaGhtuuAUTdmV/zbv7t
Za8aQcrGldyXc/I7d4ssemPedGxtHpN9DFK6URXKnu6UIZQRhk2to2mWi7Ft
qJzRyjUR30amaLGyiimMOxWLqezL+Y0oyU4XECm0KDSN2B8PpoiRxJxRbOOl
QlYIARvf9duCqU8GF7qsHHUiO+0m7Xjd0smPvbG+3bVMKkzZQX6Zkpl2/Kw8
1SB6/1yXp1c4+/PdtqaBm9QyYONQuUZBAH2agQ36cbIi68ErXA0zd8WZoupO
wUPDHqFhV76duyYLKJVsTfISf1If3rpwXpN8wmbg5j+w9SzLYuEtkV/OEI21
ElGDR4NWqXfTOunW31so298arVl98SvJHaouubt/1kiQ6e5RWQpAhz+nLsQx
gqPLIwrMTxK2ogSMFOsErmIDNSD1Z9EsZ29Hn9LkIZyfXlVM4BL65eGakMtI
GN9JnoRMZCCSC9MSCqvQtrQXJA+lcJ6sJCmYxpnMFBzz+qqAd36UFMLVthxg
LOZe5NLynKHN+KaYV0JltL3VRHtf4aKRU1dnK6hoD2dP8qsVh1b2JjL6axWD
TLx1UWa7pGYdpeWFyBsVZcGKumeaKWo38WY08/WEK6yLRCbf//qBjHa41SwD
jMa9qgAH5wu5Rx26ErnFSkMdLlWqFVcA3XkbJWzwFT1ytq7aN9OUplCc5bGB
oHDsJjWtHcpgDtF9AG713Bn8ZPgr7bDmgnWwh9+kOvx1dTW+Qt9F6C5CSpzX
WdIm7Kv6I3qakp9NJgVrGFL2Wy+qbY6qcsdUA82mcjxl3s2nh05oOpkx/kPj
e0p1b9P3KmTuLFpT7b7xv9ghaPdYnJ1s6d6llj/t8xUGlxENzsOKWuWeuAPB
z/rOBlhkFdrpdkLNiGXaY6Xf2nIIyz3DfIS05/H8AsUFZiuh7jmMA6xHNCwq
gwQgdGuwaDfJ1JyujsA940zXiMCUsNKGyyh6iD5Nm2+KENKHb9TejM9xttli
dOBf0U5l8weg454I14IaQ0DA5pDPoVDFNZoh06DyHilcihCxvozoLFxrFp2o
Y6Tlr8W6HKEQMV6NRWYUWA8qtCUz6rf/u9xGrFZWA4K700MegjNieKkyOOgj
CbsIkyebC781JF1qfSVi/J+OepSKo/VvlGL7rEswxXKvkvKSPq6QwLd2srU7
4KhwgR1cLbVZn0B7xwAEoNjq1uhepqXhguKVkeixbj05bn3UdLm93uY2ZgkJ
7mRG2VPhoChjhbEYx5ljbalDJfht2MRm7UAYZXU5618hwxfLdb+qX87ftlHc
WxmaxFRe9/gRUztM6REpuTFZdUfT3PxrZnYVPWE65ItVsU7FpCh3vmWL+6wC
uQIXy5GsgFhjbDjkVSilwhjQPEdaCRyrjGuSUIoBablPCIG+BhW9EVyTfnjq
0Hl++uS6qC3/J/2/bCH01p1wGAmYpL7bSI6//6cRJAfqjIufFBZfsrnO8Zp/
AmUxdFzDuAakTqAFXmHw5n9Ccg0G1kaFMeZ/d0Ew0x/zCgfncFpNcS6bJOa7
bJ48WJ0n+fv945bVOO+Sdam+7fol622pg1L3392RDjrPARcxeAeFABAO2V96
gGlgxRlcQ3GC71f/1pr8Coe5N1l3Fyp0MLRZa0WvWiE7iORs8eCVBUVfdhDJ
gAHGLiG+jnkOsw7BH/2XE4vlYEIqORI/HJfFnBosD+s4MpGy02lbVws12mYx
tf4Lwv1OTutsTbKZvKbpg05PJCYOxVLJ54kCW34VthF92lzmETn96y1h7fJT
0Uhhh4eUwoIihwWz+zlV7G/FZ1CTgHuv8e/HeSkzxbQOC5W3xgsILYiswKDg
PerZFlgRD50etn2OFy+ynAHqS7PTITat5cNPnofcAC+J7IN3A8BRYd4mr5T9
NVMRq7JhzIX/CbHBfTuqqMf9pB687w5yqf7wQUwsVmd3cTuPj+xjZEwkb6FY
ycrXu0L1Qm38XyYHay0hhhAYl1ky9/igUEVCdO+GnOx4qTzm64eyHOqLEySU
+579uIduHw+xrDYzu3HFwO27TE82ZO9v1yH7LXyho/zOLERyxOq3+bigbA9+
nVo1kB3SNjPEijG2Y2JiGN8WlOwQ0eLPJ18Nb12wthx9svZkurogqTeV43SU
90/k/+5l0lRt3NjhK1HviAZnX5hLl4zjO1cr4EsRbH7X3IukAYOD9ucZ/uut
tAzjszCEgqVJ5ZleUbPm3onJ7gnMw8N8kUOui16/Cd/gqalQ5hItUyUjq9Vi
0NlM1poaGd5dWgGZpG2PQVc1AqsTvRotK6wZUW/Pv+ct2iDXwi6gQkqXN0mz
rxEF7pp53XdOqJDCMJFikBfs9oaYq8ElnzVEn385iUVwX7mje4llE69bgk7w
6lnW6BhrdaacvRR5IrCUMiR5WLcQ5a+AFC/FeR6NHJozKyx8ML54FTNSaO3y
oN9YX4fVvoOmuDlh0j1IRwadfN9It87OdnkEgl06SEvn+49p4erZD/HjaKsy
Txg7DNdxxv4Uy3gzWBEFxjB5V+M4429xM+KIt08+AdE/OdVzUJ7stnj2ZKUg
ZUZLymCRpgkkQOJl/gHz/tkZtgHiukzpJc0xo45lK4HwMTiNPihImAdxEota
p7vdMWNF91b9W0HJORVwYndvh5vmBzdpNwUIOOqIBhjfjaekjqyZQHR7Fndw
DKXF8rMsbTLsa0xiUSOjON4Q/aVxMOgzC/dlrwDLdT/aebgcCvyzFk22KNdg
OFiZRZQpRMxKZ2qCmro6k7uW/q1n8gHTKW9d81hl+Kch4KpCybdXrZ/WcNiV
PAxHsp+Gq/QN3GkmQvxMD5tXcd64rZ3+Wk0CDQKrk/f7Lm/LgW4c1F2TFesp
DnHBuhDZulHDcLO2cUaBKm2h8o6D173GOJyHghZW3m4c8NJCEP96xf4zMEzs
HMNxbWdzDwdsf8vtiHxmTZ/YPKa4WpmmB61T5TZCsHgWCbnpw3p0MaOBKH4r
4V8LuuKysAdSHaUf8d7QaQKCRhgDa+RusnFsw9RstK0IhvwRgOo8fwv8Xvke
H74pLsYajlbplW82iFkXKLnWnIIlW14/K+wWIUkLP5SLFFs/Dr36CTFNuESs
KxfuOR/QiRrzpyOokUa27kfxg8+Cn05gh9LZSGIB123NyM8gLq06pcb7TYQz
F1a7qhhwZtJ3KfKBvys7mWc7pA4htffGaWuNwySSZ5RQGeXnBYjftsiWvbYV
cmW9nTpNIfhBPrzVnP70ooeBRQ63LtqfVtbrYxqXVcA3A/sCpjNJjQ8lGrl3
7lDFJeNWKYc4W5nJABqtd21GMSEwlaykxLBoGwI1dp5J1bwx/pYGmZBAooy5
j4WioBaJ9siPQjIgQmYdey+BRVWRAXUQyLjRjz6IuyZUuJqRp5Raw02Mma3X
TsPYY3Bq2IoIo6nSlE2veSFpfCXlN18OowTuBX38uuPSSiWHegAqhb7L535d
ls7z07Hwq6mUTxTGoD/9M49Yu1uB/uzZSPucxeKBky8jnhXXvV8mvdZceJzm
IijAhKR0Ppy/GgGpDT4tqi7AdtU9QvRli56bwbr4XbgwOUcaDQabZjNNbANS
Qg4g4ZryWNTod9qr/wpmxJ2nt3aNaFAhsKMwpzB2qG8eP9nW0zkQvKeBArIn
efdmaie4Tfkc25/Zwh+rfiCsRITTINKFT8cGvJTDW1KGoQgbLnVop4ahQr48
NQ6KqadKegplqgSFSGrJ2AMoRZGnqq4J8hr9qY5YDqGmX45Ope49IicFkMgb
EQyzoRYdpQFAxLLDWUcuyJa4YrcAuCEie0bm56LcORpO51j+9tVzi0rn9DX8
Ohn8MMEZlLnEz69f4DGsEdXGzW60PKHhfslf1cvQmoWsG7vkS9i3nJ/vjcDG
VJy9DBMXGgmvolKFKaf12VtahWt0W9gqpITY7DxpjzYk7oy/j4yo4S+h2Wpg
sxWGwGTO2oypJaLYiGfMqDGmeniiZZR6nKrzw596Myk7ofKd8EDnIMIjYGJi
XTYGUpB0QaWPYIKRSMMhui99ZAfZCQ20npmAEaR6Ryi5yLMndzKWfiGkWqPo
EjuvlRuJmepNR7bW5Qfdi6tKdOOQtSDO8UpGk2UVjiNOvA0bV8mVMA0w2VXH
IBgZp8ttP6kl2yd8q7f4ptMbKK//S1+OiPGuWolCy6HfLpU6HJLwt5HrYwpL
JQUVL41MdW83oL8UQnV+nLf6q7Q3JrnQNSbyZws1+VA1aOIFFxZ8N22sPIqk
jTRx+jh8JWzsVOCC2ubIeK4rJS4IEVMhR4SiP0OszS3hawFQjS9SW8Lntjv3
wJLSIqhfiyJ7msqgLL3RhclpXoAItqhepAbDjP4IBQ3z9Tg5DRBwyGdnVv/o
mg4GDsl8Qd9s3P5piQFKwrucPka4Bdlw4XJ0H32jRGfo9gC/09BcdA3xCry8
GFnIGo1IhM+pCVtiVU4/fW3CxZ6HsW9y6fEC7ZEf7OSxvAHpPBtfbEVypFGa
6a1MH06E/J7KHW132k8gcPzpCZQ6BEq8o8pSd2vCt7WnNYkAa2R3Gff1A8pi
6Y6USopWvZLO3A5YR/Uo+E0lbWTWUl9I0EOsnZ3Hiyc2QKXaD35Wddtx5aT7
CQsXXpV/jSf8XvYQpnYHWvkx5QIs9K+McgCXHon7CFZKwhVBu+IC9qRVmQaX
su8VvFP5dJgK60l3g5qhwD7TagY48cfSq1vaZf2zNKiTDemNJhYfXnLPCcur
MiuPdKY7JTpln0fV7UuSHi3Y1x+ZJDWvOonyqFR6XKjTsAzyPw3OrqdpJwsC
iVJs0mSfCbbtz5Lp4NO9R7XuRYN/fJ/7g7Xke1yehX8uTWZVabS15BOqfp7D
HjZDwVGBw0glpkH9eeh1zWCJv3JaPJvRLZkIs2X8BT8yjf+dwtHVEtr+OZUD
iPuBX2jqGuf+69Q2jsiBNnlipKGhtgc9lye+DZ6wAXUMdfDgy1UWAbrbphsk
MSkrqm3J5ZiKuF01qD/mWfk0lIowlVsgkQho1xMj8KlDjEJz4bndYRbjXvco
BGI+wIeIKNaP0KxuOTA5svqaPTa1BUKmpaS6WsVani8m0D/TBLnJgIwYZIyR
ZrT7lHPU8dolWAZAmuGgeNM/2WfFBDadZswxIuR54Yi/F0TQMxjdX/YzGeva
GKf2roFcBKrru5sHuuSRNbmr6E8qkHPsgo0OoYmW+fbPpcqcpQ+SWEc2zZa7
lSscR/quhFhU7IZZa9JEcxFo4ggq1dnDWSrkI3IP2oIweDfROOsrus9sNQ6t
Hep7emXUyPiG3MCopjKICbLExBbQAfjq6Xjc9peGBUQg5bWHdbgpJhLxYTSS
mirRFIF5hjVs/ZbA8W62YUzx0HxH+W/l0L8656RtbgD7Zgh93c5TcF+DVGYe
0u2AmqTlIMtXmB2iD4RTuYJAZPAul1qZFXdEsLm2sJnu0yjnKPgvadqfgx8w
VtwTDnLK93KUBPLmKLkTdEIKZGqBFu4+3Odyi0WfdP9EwbYUY5Mri4Zwn5vh
FVftIMoQaqX1DiDrKeWex1ODuEydIEqug7EUp5rVDTOUstJye57fEVBcE5c2
pwdElLyrG/cIxBrR5jFLZOOoYuDtO78uKQlO9v23EF3vUWtNRm3j3DwSTzyR
qThTQJgjldWBLO/05rwteQnW6sIAiksc55LNIbmJEgUQKRxzDuHPbdHLhL9z
WJMRwrv/80+rcpQCojrj5G5Ihp1FTeJglsMfQkVZXOkl1bTbNXIfewJX0Cw8
CEY5p86Ad0JgTXKtc9cpYHZewRqGWv8kPgMCBCbQ9y1hjkUSpqfclitQneXj
iXV7AdQ04Ufy9rtywcg2Ua+Pyl4x87Xfs5AtUaZZH5ZQHOsz1gqmk3AQMU7E
CQ8T/iXPaj3FekJyzGOph5Ld8MgiEPSGCd2pNaMghljY0LPO1nnjar3LHCDv
qfaZknHeVthKGzrz2ejPbpSDsgzatrLO5nRFOHG+/wY3/5KoR0BYIja7dckV
x5C2fJ/nsKdAn+Xzqf1C3eYNZE7NfHUKAWx9FFOQ3/uYGokvY5/99AWA9ODM
KyirTGAn9fiYVOeLAUsq04rgOo5HBbXQmEdfOanQnRhAdIi5uD36ldKqczeZ
K7SFHhWP/UO5YlVDbjhp6+WGJsVVXCQELOEGBDhToYJHVHnjldnwrCPRYsmM
X3815i46egZGfw9gRHklcmTXUJn5Yv8rPKmqB1Zxdt+Vlc6fzp9XSAPuZXh0
9FJSykV3/81SU/3o3NyxHFrpwD6/KxsAHIYh8npqv13aPHfKHyl01SRBzAti
g/2nGyEwj4pkNHlY5oe+cS9RDOG7JT7jlcrQaSNPMcpJgOvnqzcca4Hi+KPl
eiG9qRhop6I4t/3/ySS5PwSB3MqLpVcHCXlSYaNAXEDINQn7xXkctZ+hRKxn
8yAxsLcTkjFoYwH21pG19ZJ9GvpSb+at/caAMzh605T7p+cAAP27IZjz/hZB
qmlo7yMg2UqMCBXh5mL2QNCDed1czqD4hSjGd4qwzDkUMD+4di1c1Kz7t/VD
j/x4Jj1XyUE5AH3a/ubEiugFhIR0mmQzAJKPDgE5oHgSVofjs24s0rh0RM/W
yaCqqFPoEyx7RMHwlTuS3zLEe8v2Eg/rt2esrzc/1U1oERNH0SYVZB5HsUxS
7/R2rqn/HOOFYPd5SKAp4At3DfqGZq/r3alaSmo/lqA1jXnUKZoZ1ITN6MxM
xu7kv6hleQJ3EWs1jVct1uwz00eVfcnpxLZnA1y15u/ouIZYmAiMClThvdEd
HSbRvokq5nf4H9agvK28WdbyFUNEZzuXf//0zdmBPx2zIcbX5uh5WnbnGwJD
jOHnvsj56aDJT7oRU/RLVSG291eleJBbK2hfTHhV0+9wUUe0lQDD2oWQkhYA
SWFtoUi+egnKbdwPyO8e0SKnrw2Ih8YBo5tR/+mxjv0enlONMZNzlH5yONxx
ukLYbWjTs5AmP4otnNoMLjveyZzl+LicR1fbGsFry9O0pjjQH0q2d1jiP3HY
e2i49o1isQdBjIabhqD8VsIzaWgBy530xLDTDeCzNM0oEwNjfHZabBSWghp9
Q9pKnwWyIu1seRruq2NRqVhFw3M4FK57DDu1xUAUJO0zQE7rhGZfYSaiDrYE
yC/XTxyAn7YWgyChQagCFS9vKoMX1ih85BJem8WimyOOMbFhkuEi98LgtMJF
tSOO/0hYDP5aBJ8mOh51cBN1TcqvyiMfnnf6ef7F388Tpvfs6BI/8nf9gGkv
NbnwPUf3m0zYIdu2y3p6ZtbeaWUHL+yzk5S5CzeHDYf662cgoZwvbKzevlhc
GHPpyWoC8yLvqGVtpq0O5WpAzci26BZpxjRXw0y1vpc4hTqiqxEceSneoBrk
3JSuEPLycF7ZLyZk83D6FvnBxf85v1D4M359zFmBFk7i7q/Nxq9fJLLVJR9L
2SGjSVh4nWXE1zqtxFtsO+d3Y76Bq89KtJ4AY4YhxOMJ/QUe2JlfHekenJ2h
3mwx28+cz0QuoNv70zoDIpYQIG0lgGPYa+nSvFVes99zcYTB/uIETr218GM8
mWaY4Zw97ZLGvdnYegkNBZNT8ZaTJoRCUYc/pugETADFwFCU+VCsFFhBd2NI
YPf1H/t6mE5yzaymSt+BNqZ5x5GRlxhJiIvOocZfR5FxpWIBdssJJhb6ihkD
CUAAxY4Q9CmmJEcrJqOIlbozkfK6kQ2zEpKaRKwHNcDKcz7eASDlylfJIIOe
BTBTzZo+/AxEOiangCPco1PqQP+VWJ1y4gQ04VeJziywkrSJB8tXrlvVDDQL
tKqcgDaInZCeFCntXMkRts6/o4w/hidvnQZlWnBsmUbkdkcldkbs+f/nYsCZ
+bi0vSgYzXx6Ewf4faLq2vM7yedvYWUKkHAv0aIiq4LwTX8w3C7JsFT/SUhl
Z8KenAuyKxferg+ENOv7vLX50Ron5bTdjeDnjPS5arj4ibSRSZxgknMg7pmo
YnF2oL0lFiveQv4YqcwScn7HMIn/wJElKg5du4x/vb6J8d0OgvG/ghmMu2M6
tjJ05/URbrFTOfZ8P/5zwiiQsH9ADFkUK+Oiz7+OSlqVAHE10O+i6+0UeCtL
GPIb0dGSVDBoz7glS5OCOasWWm1JyIzvB3edmf3EmbQdBriHLIEdxD21dzWJ
Bx3WtaOFV7j9csGB6u/po5apN2uDiZHlV4pUFSktdoao1X6srX2J3C77GEfo
qPXN5UBa+LhnS6LLyF+qh0ZxmQeEL67fHCmJlSDQflpJ/S1EQrqSAC5OqQdc
GFauF2p6dslvffAq8Q9HXv8fCCTsH3Pckm4x/vhBW8sdCwpPaDA/suWUUUub
XS2PiFHJTWZl4NiQUYB3ILfibwNrzGguUqTeg/4ftuFIet0PXmMzQbeDsbCH
/zBeS0mbNB/eim/K2TZPjWxvaxYfwtMKDDRA7wGEe2FIDi4SrR0hJfjq1quq
TImLiUyUtwLy1YrXm6KdJdV+1yq6E/JeEYus9nohatiCc6KkXCiTmh9buQrx
JLZiWwx/DmAxJhYPrgVS77SEYrD/k7euDrhSZvwSJeJYg0yzggSo9TAKafjA
SGxrEya1zWzDJcYRsYKazu5gYbnF4x2Sz+WkTXpQvS6ioeDPeyjfmyM8b+ie
H2dyk2OMWJ4Lzpz3zK+ZXMByuEWLhfVdk54EaJ3OCythNRA+mROa+N6x+rLZ
TIvvzAJgm7pt7FeL6uVEOrPbYrdCIMRZBOwA0n8HFRj3AGW2wn4g5mvbOgCw
m74OX6ZBIqKqfg2EdFpzPDEIwoQkZMuacGlb5hWvgXVm7qoeNIwe5PDiToCl
OoS1eOTMCZ8OTfE6G9LRbrTOwrGxXXdgOiObax4K3XYXmsxHViaCmKLb41Dc
HD2I5eAOwUJers5WPGlga+Z9AdfxjA2aE+V++DXHg13gtaaitLuib0OGASoo
gUWuaDLPqvr5Jl/IzZufMGT2H5aJdAVdzKRSXIll1pHl47jFyiNS+je5UXbl
mBeqcIBDKjUDclaEiVjTveKnxJ1y8gHXthcmq1PQuxfSk+S3m7yxXsDquGTZ
UIiM+gDE+y//RGx/Ln9OzJxB0Aj6nWlxPmQjHpgK8kjq5cGs6VWAsG29nkX/
B9DFF+IPvyq2M7YTnptjzh3ghI0i9He7YHzq6DmpanUvZwcXeBwko0k1yYSA
IPTHYQbP/eVW9HO5KWe8oEPH+kxcNtv9OMOGY2dRK0ERu41oVD5o0H7QVROM
BZsvmfNdCurdoHuAZCnCegicANCMJOeBuTYSWxWANVz1JDyiQPCcgGog+hf5
wieSIZruspi2ojXopJV5P6j7Hr+FCAXy9uyJVs2ESyC9Qg/ZRhpzJNI88WtE
7H6xHjbZixzsXYXe6/BvbdM/8kWERXIejSmdcQMvdL8+qjUfyMuQPLfMaxM8
xhTklOFw5qzS/jXJT1kXULVoFDsKgWGntvU2z5/+Q/4QasN9Y1xAOVQn5h7T
cWlzvG+ZQ/e/ZIT6rfudEqXIRU4adgNJL6tqBAJTtqdtHdvRC6+SxdWDx94w
bUvebMKiwT0Zl4jn7gDMorfIx5qGJeoRB6ObmZqtEDY40eYWiX8YKLw7Bo/W
KKQzo5wwnh8vjaq7D7N3q0u0OA7GmdAt318dZwWyH/jXB4rp4+5pBLFZpXZT
6J3FpiJrK8A307u4EFQOr3SfCH3cz/8dprjsU6zuAb9iiS6r3o5II/fKlKyS
fO+rnHF7uELSrILZKZHlCRjv/rwhYXysL3XCZxjNooU6pa3iCq9MbDCou2RY
q3vVDsv+z/DynMnRi0xJJbTqZHLCGGC2V0dKOzqMFIxevCjILZ64Un/z3Jp5
NyIybn2+gNmnf+onWGUO93Ds/OcGb8h4S6A4KFyCz4MUb4kLZQuVKzCNl23F
Sy2YL77ZAxzKAE+J19jDMvxQXysbWjKvk8woNEAOOZQuTJ8UIq3Bh8Nltgus
TyuAEYMzaMrxYVBBfwOagip1a0Fj1v4wD57S6WBsMLOxZLm9+m+Sq2fyUT4h
ZEe33oe2sjH6FAj1G7yy6woe71Hhs5eJJKGCTdz3PhCBWsyqenK2N05/Mc7l
Vz9Z863rikrwqm9i97XHNiWjyT3/QA5qAclv5URKYWzH7ad90KmmFEFEw2aR
Kj6MSPMIC3wVXGGWF8SbzL0mjb7Z9U26YbZ3jwH3tT6RGHH65kvwVkoE900v
rozx71NI0rOcU9M0jcNr2EvvapUNUpP06WVhVi3LNePHKNEA46T4nfqsFcmE
h+hdK37A6sW4dGQf+ovNkKsScfqh4wzhVOjvhl+vDTErEPvIg+Ke7piOXJix
2qwUWsKMvP6v7buJ3wE64mCiP3P7VVr9Svpc2IjSjcSbrdmqjBHZuMM6Q4De
RASJRjUCrVkDYuCSTadROekvuKw0HdFZjFuCwzVYGa0XwgPvr/biYBxsEVOi
urfLRGw9seJS4lrMO2NeNcWbHfMIszkS+ASEui0zX5kraihA9Nb0NxBqIk58
X49fUJYUzUOwGg8nMCdzSWWi57cv5gVAR+KmCfihOZU9J99SKyOwOpy8CYOF
BUtEZ2k1oZsxiYym4bIcf1JQf6GzBcLv7rrHOHItI2qwj0k3MWhIVM3zOY9p
s1OA0z0oF8gScoLaRSGLaY5FI9rWEhXRmB9sClaZHhZG2RziTzRWGSDth8yH
kCJMfl0BP16BjS+teXZBsh2qWGYfVvB/kJYFAcij0yYvx6rMpGfnv5C9qxxJ
PLVAWk98DPKCQb/VzfQ6lpgL2jyrRX0Awldc/i6n0mQnrA9NKp/SvwS5gprJ
CRSJXW3z7tLwAl5rGKAwpxWUFVWNmmCQR/s0DrDnoXe5+SDCLxLfmzQmXvz0
L5wEU+ggUXMHBu2vo8jgqPMU3VZ5fUnULQ8hkhjIdxCBXA2oDbJpOXSkm3qH
LWDM5tOyjZY+ep/cNZUet7BpuUfAhtIAc2FlUI0Fr5z54vV2MQwkPvgOxyVI
hhBJJchy25/yrrWSBx25YHZrvbmwnQgIm9FGx4WXCYQCXDOr1PHmdDIUNkp1
D0Q5mhYCM3x+z7sn4vKIdSxqBIjeFVO0eUIIyW5Gc4vGU+4bo2AZhzLkj0o2
HlxZxRG8Y1o8UXrCNskQEUFVDnNNuUlKU4smxWZtyc8tbUFzGSpgwgZw6ZLG
+dkMAmrl/pRS+0qnIzJf732CWhO231AWPjogndZue0xP5h1TObG7cc9CScZD
w0lgSPd7dItyr32RgZ2ZuiiYo35+wx1jFZri3qcqNIEjPXRvbhYPNDsOn0jb
tDZgMjWHmGlbeZx3/kcGbatTS27U6t6pnHHnDUCC4kGt3s5Dc25BTDKXSjqL
0JitMbyrMfFpI8dD8iScEJwsobdc8t9KF3+FiQ+iMTY34TNMgII21Zq4wwM2
xw4gvF3acOLfu/0DM1u34uEYXfGxEvJQidVGlEgVCN+kpChGcwxvL+YEEbN6
jZNaF5UzkzFEoDJ9BLhV9R7LJfvti2pt8haeSstYxkEasIZTZj9PMMmy0Fw9
fKrlJ0FgDjnkgkckDpvgkSYraW0JUDwJ2iAQ4MXVZCXFGjOKSQ4SeBPVfBns
0Je8DUakfzD0nRFBjOd05lkHscr/7kCFG/SK1TSM0T3F69lLAzvCLjYBt3i/
4WXW+iWSRsCzS2TBdU2GEJvFWQHdzOx0CMFpVmiwLqdH1VHBrhy5D6dhNk5V
G1wLJPwM768pnmmoJeas0fktK0rIOd5w295vl8zsDLmgA1SvQX7NpVLtfvpl
67I4K3ZPxfhhxwDbkWoxP7hAHC/hsXh7ROnwjsHz4v9YRzWHFJ1Ph826cp8d
vKeXOm2sK7dY71BZ7zubiq1LKTc9J07Mmg/KoQNCjIMvOn/88FViFX1lCEO1
MolNzxTjxXJl0odMXLGISDp646xv9kgfypCkvhBRZhvUidMhuCxZjxRcpC7w
AtEROq4rRkVQ/Hw3OxRpfEvOiumKPl169iuoSzxD44y4lTA47JxIgfzyUO6d
5OkSmdIqEM6cXOteLtR+dExA7bNp+uLcFedsPdGCDWYh7MwPDL31epxcOABa
riA3JenvYEO+c6+d5fD0gKZREK1ofKSpiAa69iP9pXRbviLcNuqb0mC875pQ
p/PgTEANkEvyno/5No2Y45qnfaAoVpUEGTXCJvoh/Q0MDccEMIVt4uOJBpXQ
EgYd92Q4CTqzD9a22DlgtjMbtmdwnIGOdj25P2h1AQX0fu0YGRF5pWu/KYEE
EGM7Vddjij1m02gKuwdv4ORwOril0GLb2+Gu3kW9qrDEo9Hn66M9l5GQO4Zn
CxFDfxJ70oNiftRg1E2Gu1B/EyjvGyl1QJh6/q9d90SqJ6wGr+EcYmaH9+qf
546173YeMZlX/LRqvf4Whn9aqoceMe3iauM5jV8JEW+Mabv98G1ZqmnpLGBm
TgrkHnpaokGt2faERzN5MfN/xnSX6gHxU59I4fnLtOHZqC+EeDX74JCGjGlG
/GCQgZWpYH9oim0d6+UZQ1pKWJlKbMBgSd+nBBs3GNSKyd8c48G2h3tcg3Uq
qRSNbylqx9cGCOP3t99gLFVZ4lEiSDw6AkjyfDWl4hKuMFeiNrjTFeLgWhsW
Ckyzvlpm1S2LAnJKjecoqmO7Kj7wM6nbOalShjHgsN/hTMS2ZnT3gwntA81Z
fVMpS0hrhzgIa8Yxj6MChC5TgoxatBTO6sQnGlUyQ626Dn14WxlCLKegjYqZ
CVLLzGxcqUkLa5IvCkrcMxD1RheWCv7F5s7wkDq3FAcdK+49SLxJJxjeIv0q
rfHTfXOtdhYs+mOdUpew3jn009A9EaMyIP6Gt23Ohb8cBY8jMAInkH1gZTIu
cNtO0suTGKCXJzaCPpH+Fj/QwkOQgdfkMjZ1ulKBmGaG6EBjJZqAKX46PEBl
DkSHQYMTMR87IafSPnRovPIHYtUsCBdxS66pFC24jZ2mW/i2A75CyWVKFCTg
8yxpoyXBcS+dlb73ncEFplLNfsfobgqSnL/WronkX3sK3TGLnBd+QwoUATJP
mDWWfyTEyWziOYJjOm/dZ2TA1sxQ5J5bGX+6h1392MnT8/9OCDywRnDhmdr9
u6nCiwDTPkTbqshOuRtmWUmW9tzFMI4eDmBT83sDGTxDfDaG8XYkuLQRlo9A
jRV/G7OI/iNXhAQf2DfwVjYe0Jo1SVsbExkpMnKhhxe+ZPrsF4ge82a4AOyf
tGfjE3s9oO9qYEoXAZeg2CWU9PFJ1V7r1xfYD6Qar/Xo5eGbYTfW0xjKGYxo
Wz9prse9yQXJD3tNePx3W0vErUOqMnBQpSJ5Cf6kz/9orUWh0mvi1DeiVszK
NvvadSoq9XUYMVsbHL1JD74HaL8FhBfYDDvRqMSha9nnQKy/n1rciWJu3Cpq
8sP2kHWYRrQokIYXEgE5ihYKC4boEAtBfe6Pv2nekWVvipZWBcNB8ZeZqqjQ
W7Buzn/JTD/IelIHNhyq8MAmb5594D7wiBKC2nAyD1fVq3aOhauTnwLg4OiH
jUSDZ3cfRGWS8CowWaqz1TqPk3RyfXEH0T44D6evPDBdJ+W5XE4BiHeELk5f
j9lJBzJTZCJGBFtyvysoBmd5+sNAWmwQFMfdkJ6LinlklwT5y+NTvYr60SCH
/2mLZWqnPcCmqn04T/X3EI5zYY9HbCKOJLkwEZUPLdqvmKHi3flLWZI3Ch4q
Y2p6QbRA3/XeFT9fYc6mN0LVYVQlAptSD7AX08VWyNak17YdBdFO2w7MZAfl
w/GKnTDmhZW5EMDZU67DQ9Gr7523CmDp5d1rN+1cFQYuP50GTB8PR8Ds1ZJS
/CSKP8LvOBYYRFRuUu6YG6GBmmfwvTe8CVgCkYQtOkrmlWOnMqRkaIY7YsZo
ZWXpCkaZve/b/5O3Gn6bfi655NnyaqYNlFnc+s5aJSSQ4JHUT+KSnIG5ODvT
mMMImaXyAElfrAOuZ1zpelw7Mts9FHiad/hjh7dwIDaHtIFtXSA+LXAwFPXG
paVU+YbOr/pEhMYsXqni2m15/ubH3BKKtHCBZnoJP0i7vo2CxvYUWwVSwoMu
bGZbznMkOBpP1IEfAp3+FpvDeY2CXaEEA62/73qwe8imdkhlh8nQ7qFEvk7I
cu+rxtPDyCQCEUKtxo9YvBtS/rdqg34nbclbOw2GYDcXK4yli1wTL1slvw6H
la36fz0PDjJ3HadtcnsIS05fssmWoGNdcUokVzMQWVUvY0WwBGwUJZtrUFrS
6KfdfLtbOpRWoqiTPeZnNOIOBzki8LFouSemIOVfUQIT/jKODuK1bq4TwS85
cqftl2mASO4o+gk08FHFC9s/p81//qUpMP/E7c92OMLK/9F7p0vSpZISdDm5
pS5Th25IYDLHH1IeKXK3ncmnLvOTyplI+JlsnjlvSITaAcK1fxtF1wA21PCX
cb4jTVQh9slJ59sIGxZizcOGF5c7W7c96h3fqrIaELzAILoWeIGBBZOka3RE
TT5MPgQc9C4283dhaL7j+Bx7Y3648rwfPKLAln2cRFfoPyuXj+8ble8HDrA/
390cjVwQRERs8+7ScJjEX13JxJdv3pkGa5EkuEqUe7qgK2r6cKh5KOTC65wm
DD1rPzrEWONMqUQLojjl4zJVLl5Q5C3wyyAE6P76Iz3kmRUOcDyrskufJl96
IAbc5k7yJCAadecj6RoJN2ehdQDcJ/yqFZIefgMsm+BpcDpAVYh9htguBf8C
bpoHBeuoDkNJmcTnyyQYt3/JvZm0D+UypTLEJGQXzjXdIeMLvrl+CTujAS5d
JEgQfC0NXE2ub22cviiG4MZIo7tLl/az+DHdp0EH24j7vIFypAip19Nv7cTE
xhGNxmhN+/+BnYTqOqUu+/vhgmM264WQs0TSMZIGSieI50Mrz6NC7W2XOIS7
aQ4XUveGxAhkG0Jp2/0oCyCefvJmt0ViNYa+Ms+xsEH7VOpdVwxHybB1Bnhl
waRl7e8if4yRLBQpApk9FUb5MGb82XZMrxezDj+cf7i9hbUTNWEGAmMk4bDt
pwoaX8iruJqLgVQj7HqL3pyDZFtAPjkYBOe0ztkczzsdBX4MTk5Vw6wU7/aG
qzUmabCWEO7LpucqK9hOyquHv9z43EJF4w+R8PakioaYBpFPNz5yAtYfcvFA
tHN19nNUE4Rwo3JMR7cuFbBmgL3lJM8dINN+U7/l+/bgYzzUHfeOhjKquCVE
X0xT4L8Gy/neBrNm66Ek3tVtSQs7H+3jxnzjtNeiDMe5Y7UNxnnT3vttOkdc
kSY+L4UHWw1yW0dvBPpn6xsHgQmRjzuqaatNyTSmSHTuRnqMcDB6JH8jFT5U
38swazlvaLygAoYt+1+fALYNYL5YFyC/IrLjtetbM8W1KjBpSB4zx75JCd0P
1bA6UM8kox7RjW0KCGTGAMrsmMJ0Vqkqxi52lYLBDq4NE2SVqLDFwqevoW3n
/z6bCV+LNYtmaxSKze+3ODuZRCig30Oa3+EetNQWuVhXh5H/aRA1X7j+WM7A
PtUXx/TW72vhyY77iDNrVg3Po1gxWmXXpaggZx5wYCx7nkK7ZUD6YBWqrFi2
/V5/PpHft/ZkybyBLGx6+tl1bXEnxke8Jc3+1rkReJb8TSaVdxZ8hksMWcsJ
Pj0yjZt9/wqP7PDJYXdHE2y1zv+fcOQe/VBjUJliit24htkIAnVITsIrU49g
SNIXvcSSrCpMGT2rki0Q3Kz3yxT0QuIJmk1CveK1dcgIA0+ldkw4TKiLwUtQ
WdiEwanOsiG1HxVnd+VQjNUqjwqDokpS4MpTPoIzkfXpwMe6U8qlUma9zNRj
EU2JXhjZVOOo4ZNsvyZjpcWFtZpRyJixHl2RqAeEHqmSloXaFsvnhGzgBfx7
m9wj/ad6/OLZ/7VuPWOIXKx7RziTs9hMQPp4wriV1YFWc2JAqiOJEazY7nf+
t7Bno2dv9g7LQLq1zcXQn5ksObjD5Kf3q6aI/gDCsmenvt6FZT7KnCTIudnX
eAzxNNaT6X1Ck36TUy7XfEhwr3ZTtuR6+2++Ssdh4zy51tDaOlTaxp6H72yX
xGrSbDFnxrbcYsIdr/CQV/0ZHmEXngT1TG6CEZdU/jpVMlusgZjPdodN1R+u
RGT9LYxcRHDOk62NpEvagb4fP4TLTuvCEh5L7Qq2Fit9utOvv4vHpdFb8WLZ
mGmFmca8BNn5q+LfU6VL301m595KNPRXndyM5qqUu3t49/6AApP+fZLInzxu
iKaZm7y65TcWG80a4xLo6vQ53ZIx62KsEhnRzYac+wAWfkOchrKBaR+8zaVS
lPU0raokzHPQwo3vMd6/bWbc0d364zXQ1F1XnpzTwUXJ1WH8l+qHiNY8OIit
z+otIYD9izXJKjxVEJ6Ii8QVqdd79fQjrJhyrywpLGBZf/H6n4YEu1i0ekHw
KY8gpIDETI9rcaN8OjLCu9gOhUHDe7mDDQ87pU2Zo0HL4wy/AhWtSDWVesnh
/kOln6QKpSBfk24pNKL6Nuat2V6JRbdfFosf35R7B4tyX0PJYyGrr0+K51wY
FZ9YNT5w8zd28jI2Adqcad8o896XoGBXq96wyO6l+lvhgaUF6SXv4u+YodoL
O9Nc/vGv8pzW3pkv2/gEXjaDwd+J8k7PZ+9VPOkRO3Sr2fzcEB3F6eqrY5sA
N6STa+TxYAixBiMZLqjGphxg2B/hrabBXOCrGRDRg/NBxAK5YPwWOFSOsKjd
p88FP018Wj6yZN9OBo3TceW75wUoOwSSfQEBBq7qHmgxeUuhYGshz4oBSnVh
dDZLHlp8W6lo+YFqFpRGoRY/rd0Ld4NR1OBotAhNrXK92YPZsY1KstsbFiBT
dyZ/7oAfpQlmziefpxGceqicU3mFWBI+HY3HItWMbBR127ViO6jzmlVljhdV
X5T4iJ5VAexicpWyKK2pa9gWVTzov/zlx9qyefJ7zY/AxQtH94/zfFdbO8Bd
OfFvMSWSLUxMwRs0vDLD/qQc3DflYsbYePCFj+fF6EgYcDEb1WWK1B0VH448
P0ZdE9/qRzfXZR02Xg3FZ7Vi5omTz+1iizQCJ6tN0fttdtaDvWwnOucotjIO
WG85LVkQRbdIqGQs5gwRI8NBBJVG9QFNBetj9jNFAc4fCpi14guvIDOJ0tQA
2tmkrWb5L1jID786qCIK/3tG7aZB8G0TFZGflANQByNw5YQtUk65wg6R1otG
7EOmZufK3Z7F2rri0WqcrMYIf/GLOOyPzbcyo78VNxAzdOsp3XI0JzLyGgCY
roQc83JnBMkQiutaFcw7WTkbR3tJzuzQ/f5vPbZ7/cbeR4Wylm3eiohJ6Pkw
etZn6C9AqAUkZ6zpP9eWVLsuk12WIde/EoicYEGkPXt3FCDuZOBl31WKUgvM
dGZTs96ayJRQ/4sIyi/J6f+NsgjTLOhSmxKBd+oGe3EOVs0GnuCJkq0PQwIH
XVRBjMo63z2w7nAr30Lrn7aSlR1dcpETufhVikMrqG+a8hyaCE2MyonNlPF9
jz7if0IEqpeGwr+afDOBwV2+9GYzsMeTz5xv63RPFn21QLskTTuwoHrFa4+E
uX9h59CypURE38m7a3Uh8AFzCWyGsQ58BjJTpn/5HHe+d01Rpdq5ndxM+1GQ
QNDlfxwKPpdKgQbm9xvGeS0TnoXJo2WyfR5OiYlc6M/PHlsNBSy0mRfrzCFj
TSzDtGzcYG7z5VWI0JLrVp+XoMi0QNc2huHi7Jl+qrxbx6ss4Vk3uZYluija
lmRZKD4HmzbPs7dqRKLeWpE858ij8OPs1fMx9bocwZkN84J4SqkKuk8fg3qC
Po2/mwUXL2lVaxfaAYqU/JizoXxIvs2WYkXfSZ9Te7146TGpIdtuom67eq+k
sSWKpAwHoZsy9myPC/PbD9UfOGrta9lKNqpCGTabXZ3TjKdmVT3QB86hJ1RU
s4AYl7BsYWu7O7ZGTDP6O9+D/D0A4ReepmfG8OJLQTjkp/XyfSLvv5v4ErLA
P5zhwzAva2aTfMmQHq0vRTTCwKtABslh2iMvlBNSZ+eFU2F7RDk+w1MVAQ5A
Kw2MY/awDr6uTvHOmRIgiK/Rih21IwFsQ6Y2zdIAmikITK8JsiFwaQtdwenu
Wa8Rb7XNXyAF9xOKtP29rCtxvYRkIYV4yqh3MhoTsZL0DSW5mCSh6FXT/cEh
xvdAQOOl2oX7aa9whTsQCyVt8mKwmRPKEsmqHKhdcKTFJpKZic2QKaSYauzV
97GZmZkl7HnWLfM1foX5hER3T6caQ6qseIscb1A+yntEzm1v++Itmpzkn9Rd
l0esKLeCpzr7zI6DvMcjQ7R3EsCHoR8zsZQw07IPM/3OXQBNnJPa//TsEErh
SxTvnaiqmctdXkIlHpaBbLetA/pEDfyWMmnUmMdSMQXe94fbli+9/hirRrbY
zThguIhE7oXmzioLbZw91bBdZLWz0l38gTGNjRCF3En1LB1Q3eTrqYbIIN/K
3FYbsJsYTvRUBGP8K7nxlnwFzIFPThSwALBm5QEy1hThsNCYWcjTCIMI/usa
rPEEbhU6/9l3Dpd+Xu+jixBex4RoNF3HyvCgA/qmxcx+Lzx/xTNd1ItnMlSq
OWxNP2A9mnXpxU2U/6vZb4A8aVXdlm/1s1lG+mUs3T4KQ2t5VSx+G7qyh6dR
1W32MepJUtAM+yCPMnQH5FwxqZVX05HQiWmYual+hD1tNNtidPvOpLO4rPeC
cTCkErBdnL8iiAICZCV+AMpPbVIOrb1fI1LOzVyI7TNzPTPvNCQ/463RSSgO
wd1gdYdpdUaWnNAmCP8NT3ZgvasXXCYjtYVe61W2NuBBu7mltStVkr032rYp
G2Vq/WtAKDrxvrXen6lEQfSclPZn0Yj9bVTMyeaU7cAa31rDS0F9fBQRGeN+
tLTsgwRPUxpIIPINaBEPzNXMosjQmt9V/nEB6DZKTzwmvqqMAC+p1qZvorkk
tiJqhpfynKi9Q4GB6vQwTvb29MDu1KSkSycmBdKM3FpzT4gm0EkhE9RMGsrc
x2edqm2YVoLaiKev+OgPsn+yyEXNZSrqYCaT/tVksQL1C1jSMn5viAsrtfJP
DaTj0f1cVbMm/BMVd6fRi4FISvBZmynNZ+xZ0s9PJU0JbP5CrvVHEHwRmMEI
LcGkOzZhkjtnkW2SlfHmZA1JDFU2IWAezPpIrhBoEx5T1a1/bZSq1GXhRAbj
Gppio0OM8ilGvp7kTD2TO73BsN+VvU2WFYS02rVHYpIy7RlWNg+uBWEEP1Mn
w0Q/Getfi+wvX41n2pSQUlH7OfA4G/2/KA5lzwHJRz2NdzZWA31mj7sJuAvw
a/6IrKUOPPLKhpmcLgFnc9LIv8NA0BhvV2EV8X5vdl72olWabZw5jM8J3w/S
hbecBgT/+R4ghjzYzIbQ1h1auMR8cYK9sXvOxXjzqtw6gaac2UIO0zwbYUVu
ROvFmRiL/y4+IPgEt1jANPGh6j7KO9Pk7QRnK1NdUFGSTgk9Qr7dl68M2hM0
yob6XePFRegDZZxzXyEdHOGCSARlTyEc/5GtUVRZZ+CW3gGcwRoG57iDJNl2
Lrg7qIzHvJk1T8GKpojA5HmtuTdyDw8NKByq61jCkaGVv7SbFeNI4YglhRey
JRKM17xDJYesZf9sWF+jf/HBEdiOKQUOJaDCu1san8IUBn05cse9WgrMS6uc
1b9jnoxkfouYNKeoPYSqg83C8vnc58SoByDEQVM+2LIV2g6M3c0njOozhdE3
AkscxRE4kX32cw50AYqm+urJERxVmy0F2ercMFy1tN8S2zizEXbAyI5iqNWG
8jEFVGtEatCj0qIkJwNOYwK0BYR9FFt0qUGsGVHrAe7yrSU7k8Y+KXEOShXJ
qPOb6sPAAvtyU/oDHhTAJwJsbY8bJHlnlUWU6Dj9zRSrMI0makzjCv1A1cFz
xtMUClCDwksqhQNOT8gVwKo9IPScDc8ZaHJkA5szH/IZ1HA65mvBMAww3kzD
qhMNYf4U6zsRWlknC123A0iNY5bzEEaig5JM1sY7lTi1iNXxywDert+jXOb2
QRl4n/PLDDIfnBDlO+kMpHk99zys1qdzaKlgG5Mu21MMU90sbbe0z1AGMPjx
JDIfboOOdYtv+1d+nL99GkPKu83JXyn3LPd3nDsaEoMarYRtdiswYKKXE3sV
M1Di1Oa6AStjxpPTXKW75UvtGfbAQ4Lx9AXCsKN5hA7X/gTHyYbAilqboBdf
mQUkzkHVSHkSz2zJhe+bjv89h504upubbT5YLMceCeJO64NPWyySYkrWjsZ+
hONm8LZRrH69rGJlkOMd4MgfarhNmYHd46VHNt7kObI8xOKRIVxZHjTYOUOR
UPEk77Bgd3bUInccqjRohu5JnNys16jKLB48p/A4bYYNZ3dICMXnbn6HSl9d
j6oFkU895WCSf4ZmqlcmBPPdH3Y9y8GUmYcCeGt5EvoahJqAcTzbILzB6xQ6
lKvii17AO6A5/MkLAgCd//Bx/Vgx5S13G3wz2kKfK/C8HoSphbOQBrlJ00m0
GTigAi4iaYyLEQaQ/JxDKLElEvjmPzsYCjxvcwQFplQ/KCPapjuTN5iMGJKS
lYU8wPtj5ItSC0YWui5H7xbWj50OF5KjnxkXgiArl9RqixUDnysIH2Ius4tk
UtJ1j09fI8FY9O39Z40MG62qU2GmQi/tTowIZ2QNOE+1yceATJ7z8vh73dHM
QRLKspJvdyC/9/fkPzrgJCx9uQaG83hzLJ4RniLmibvcFRA9pRnJJTFYO0nY
FsD9DgO4bP1d+mWlDAEpqjE1AdtzZZgN42kBNQWRBM1hgIPYbm9zWWnVh3Xw
5YgUi9ZZPP6qIFm1/nw=

`pragma protect end_protected
