// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
biNqVsUgyltMHW9kETO6M1rv557yYe1q+HS/3Cf8PVcXUCYF0D7POXG1AsTq
GOvYQMub1EfV4LyGDNfz9Wd5ULuMMMjgZKefv/TGaU5GAlwQxBDXq4iFp/hT
8HrCVHUlWZPC6VzH8DBPKRsQ4hK8VvBUiCqjlgO1ot18shfK4klbT7qXZNE9
QBb0ASFhZ93VIfK4Igy/gmsa7RX2drlvbhZs68WNEKyMkJQSF6TsArfcMQ+W
qwC8CeP/JxxEen0NfPxgQuvgI8Fv8Qvuf6kDQ7s/C8ieQzDEjl+Tm3dTDYKL
zhtMpz3b+JFUN2a5+gilQVSW7o60lwkdu0tuKQ3gIQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
F95c1wIIb2bbwzk5lC5LD7/IjYmcj+5sGPEb1fsR5l0ARZAojTwNnZ44ZH4/
1Lhbb2aG81uib121FjicANxUNz6MtZkhVI0haiBQn/nEeANaxZ8Dn8pH2S6Y
Q1vicIoOhQB7hQCxEnkIoFO8cmqr0ypf07ntNOncyar1X1fY33vScO++mWzD
/g1cGZhBYPHP+CcN6F3WAPdgnVw9qc5ZISkOSDvE7bJ6jTKq9YFAbRllwrAK
m781ZsQJbaqbCNMMs4s88DY7bLsYfY+Y54ztLFSVv4SLBNRIchRJ+9VxrTfO
EoItTDqDKJIsROh+XI4uAwfZdvyNnYLRxzDMasD8VQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dqNiq3KFnmDDT2UoaLQKfRkP1aVl+nF9KSJHGfDG465G1v+JvXEFhONRPbpn
kGEVIqh8yNaIp8BwMJU2jjD6kFrpeOu4sYiZqGX0Yb72WpQEB+XYHz1PjNPv
eyR1ZBz34Iy3ylSFTbbpYbcMoW/mPOxM2ZtYhwTPuUJeUrooVjMBoO9psSV2
7nGSj2A4Y3z2hgB8Cer2+p4e7qOFgQzEamy7gMFX/YK7r8Z3q5f7jwoYRiJC
GRKofB6ABPHfLWgJqeGCYfoQDbi1FOulS9xxYCFzDK3yd8n/TusIFYTvQm2z
3x4RI502TnsESgtHHgsDA3T47BItqt4qtnMSa/hS8w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UgJ3ZB722ymYQl4fzC6V3ckZbQUqfg4qpvq2xv8QBgEEoAygPci/kO4dyFP/
/SA3brXaLXGFbl0ch8/mMAqOOcQ4ckIoNr404uitqBkO7xPFJ2GDVzB+KtTl
CitsiKgL2QJTr72tci0Cv7g15SRI2L28K6nugXpMKtVqLFFZKNM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Is3DVpPAxCSKLRAu29F19Gkox0VAUyn3S62CN29by5P+hR9Zir9m4Yoew3Tr
RhubqCAdyoDPT1AwF6p8BBMnQ4cztmW2jsXo+3Y7MlvUtX63cQ4fu7tDbqZl
YSXgmB3ZRdysWgM9zuVZ4TXF9stkQ2UA78q8UjvQB/UTC3ZOjMc4PzuFErVY
IfpewyrnhJlu21WWb4o5zOrKxBhtSODU9K0SWjmXNJJX7EyvX/jdCjvWzFD9
epNEQw/ybtm09A8vnY5Oifea34dCgq7cbHr2nRCN0BGOHzfM0w2gzTsjauQu
d+dF+/3zkO1t7pxVsYhRSI7RlbKkR9qOY1wSIoYfKbOM4+OtG6jMSrGSLygd
7t3g60ZJggz5a3gmaZcTjpGn7ji4chJ0fd+t3AVyIwOWL60GV/yfNpdNi/6P
eIHA5sXPGOOyiU+dziY7lDWQixmy36Lj/NUn0dV3vuraKZfC7O31HA2ZTsfv
I/bqO2NRTyDOZAoUJNQ3gCJMX17icVKC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e7pYUm5GA7cq5nrscz9lKyFj4MqRFMZVlT1RghAClWHZpdYstCYCJw6nKglN
DCL9hN7A/xXSbQU3I8eLT1xJdlDSq/gUMYprvaPyrUmF4n0Mpgz9D11QzwgC
FuckVyP38dXVCTFztdIJYZp4Tkt/3hVh9GeHWcx+mPeMI2RPwn0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
t/1kcDCm5GJ31mYOLI+pvSWQkuWd37qp+rut2GDnl41zMjiblu7i7C6JG9DI
3FyESw/JAuOV3lU0kRmwEetKoRsQrYX4uEs4Bpd4KpSyYBfEs2D/OYlL6tUx
dpOBPZwn9TioPhZspn6fX3oxSD3+vVftooQJ6vTUeNJlS4KdI68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14752)
`pragma protect data_block
5s3azNSOuVt6ol0+Fh4wTTtsSteDvP0LXdDVBXDq0CtO574kZcBCjoe7F3qT
Z3okZiqseAQ3cfP3OkBOKNar3QGIZAzJwTLJLtP2DkDxsUBwEuovf/fb3JAK
txjOeOlwQorOaoIls0IhAq7+8x4hdPlQRU+02r2uLS9VfOMM8ZxYYhz/1NDI
8e2EMg5Wn/S0dd0Ek4dDSRSDyNnD05/98q3ITt+UywmalR63aIDRW0tqxg91
6rDM1LRptDvCGZMMWSPbfJGm8TWTGwvNjIrBvtVdChpJjWrSFBhRUkbEtgbF
qS73+iDk6tjVX9R6PRwx++09k4JfakWUBxnTzWRRHAjTeAOcErogwZIO48Vz
rIZgZXGrnCbinmDqeREa3MMH2piOGWcxgD7geQz1/1FfndZ7CnwQQ0AhaZGQ
NRV3PBmsN/sxXJJV3YCGRL/YZ+7ver7y1jj2bri3bIKi9OL0gwmWJeiCGI/f
W4E1uiQxo+BojgnoWh+KDzSzKPkP3I/eww8zklcLYk+I989HCfpTE4UjbgVh
JLzZoxUe828brkepC1tMlX5HBCN516grGuTrSrRZKblnTToYZxJs0He0UJnz
26wYr+mnvSJ/h9776mz1c0ls1tVK2/Ozu6HoV30GQDrsfPDvRZ+jAd+9h2Zf
tIyKRpusvlJ6zCaVqvzp3Wy29b7ZTejF+ql0thlQOu9Q+oSfpGZ/F9cMhSvp
d3/sJIcV5KOiU6bejrkk9QLvYU5j2dA6lBm4sxHOjgm4ehN/uYZzWxjpNX3g
wy/XBpknZ3lO5ZSmk+J7OE8Now06vM/f8kxDM46ax3aB8klgEgiKBFaN8N4K
EUwuVOfJ6QYXI8YcX60T0AbDVs13GLN5OoxKIpobt/sQeXqWomGMzZzpn0jc
Cdxuyuzl6ZD5DvnH9f1yVmMd+REOZ5uCAcRZy88p/T9z2/NzXZuJlGFQcabL
SxF6BwTW9zJG0joyBm2ZejwN3JmbL5vgzh5YDqaBDyWUiAHCE2ATmjsM/rec
fD+Y1Z6p+MLwE84ZS0Ce1hACgkaEqjLpAgLclhGn6JsZ2fDYxiDo2KjbVISU
7tuDKC6W43Q6ghfLubF0rKX28djRcTWxp3IpVrKTFE9va5Cv+KtLe2c8a6nb
MLr4xEmthBWc4CXk7MNNo7nN+0ToZHcCr0yZznh9thktQQt6/5s6wCR/vfdJ
ksYQvU1n8Kw96hsq45IdQuqhz/xG5N1zvDK2sHQIGmDkzvKZn6xY3HE43Cw3
hsuYVD4G83MR5GFKeQvH+JIWNeJFboCbamCE2Ag1Q26mXqqZGVegkRC48Av2
nRYm5l7v/8EmmN2BWOjvTrGJ5jOxXH6dspJYd+38qXBcReIci9R36u4b58hl
KSg5nfyOcX+MgIjcRJH2TMkflBEYj7GP+DqXC10E7RZGwFofXvP1yw6OR/Kp
iaLM2ZwRbLOuZa0Xx6SdKsAs/ireVhaU/P1PvShBxewbplkOYcBgT7CWC5fr
Y+JrCZDqoAUnqhBweqCVGUwSYyW2SOjzxFML22kIFsIE80b/symPGemxIhLt
0qb8Z9Ia9bMdO0Jw8ToR6AYrfg/QETjp3dgiVLv2EJhH7gSQQhBeoWzP/nVK
I0jhACXbcygKyYNLOiqcehOXSTmrRHDXFwKhyRRPB67K3dXCME3CzDxI0och
wXNEXo+RIRPxHtXFwjMTpaTEr12xd2hsyv3YHEkPj2Im+rI0YRGg1MSakZ2U
8Ovlu43kvUoAAOsgpb9gxMILTNON05nHsaT42Cb85D5uj2ZidJTxLR3PiAh7
BMwyGuaGcjfZAFNOk/FdaP6AxUTVModtso3pq8rnK8RosdVN3/CTebE04OQ0
rfMtEbTwInfs2Eza9BjfP6uZMyTvuH6fZFVjt/0a1ay55L7xavKIpqyVEfVk
wfVibmG35u9K2qIACIzn6f5bYZn2TPF9fNQezwydRkT9Yinhvx/mNG7dkQ8Z
NWiTL4cYu08PJEfeWa1ZSa5MDPxhKf8sgi+UR4Qos/ahVktv5ADTrcXJHQGT
t+/0bkMB7JRKd7OqbJU7gFAUy7FhtqH5F6ftj2UUp7b0ZY3F4q91p8qKofRL
dVlgObhLzQpOkNPeYr8UP3WBro5KVFCrUL/mAN/gTiCsiOrBz7ofzF0oqHoa
E8W/2EUj+iaJgWC6lneEYF0vERFRXr/E8puqdUuseF6w9VuSYHcRCynbCXAY
hW5S2LLwGDeuHV1bECAVy1mnYAPbwL1YNys37OG+Pa8mEtTtuPQFS4DaFUdy
mPiYThPsF+27n81OD/40jBKToPqqlE4Vf+WWG2M76tQ13g6p9KRLTnnAkLhX
GAcKbyCm+Yy6p647a4HKIYZFK7ZElAcTr3GtMZcJyzzQwfYIdril3T3ezvEM
aPCIcuLbXQMoA0e3jXBNDyJIc0mGrHtPOyWa7C5J8cSAP4m/A127xDAe64p1
EbDuvOszQAPBdCm5aHMWxybSAxcwzkxhUkeUw5LuPtRtJy5rZTxSPvA1x7uY
JFUwKs7YgculfZ8jn/oOOYPEFMWU6El2dwUDKazhc85KzTei4rdHa/Fk6g+O
G/wWZVEKG8TCRqDGYRwPhYq3cXsrxuDDuml0lHi9X7fgew59f5U6G0BODcbm
MpMdaVFyc3EzimfzJN2klhuDs6YkOklqMmFvph3EVFl4+XUUgovh6OGbxsSE
kThmhzh8gdPyXCoQTukFqkV1i/PHBE9zm1Uo4pacz62uiSrUtQjIejMPTiXR
Im83x1TW5/bvsQfyiSxjyriIaEq21AvY+0lPIeRdUrZMr8A4o/u9VciRi6ya
26xQV2wG8G528BzGZKtnHRiO21b3b8sV4wCVISYO1Qfhdb4B4AZ3dnX53YhN
slNlYG3w2WZo25DE72H6w+DKQ5WxIWb04rwzG0y2LMydKChEBC6E7hhUxPE/
IxFywYbzdKX1galz7suzTdJT2N1QNsZfrLnPNjdVuVz6B9WmL5Y9vwxW5K8S
+MBFwo55bu41pOTDzRYkPC9/6gLFtWQ0vkqiFn677tUQLw26b08hTTzUEstO
RPEHkahYMgRbO28AVkHcx5B66JcOZau9E4ZS7vcRwMKZfhafB9lOYynk5kxb
BtKKsvf1/ZT2bEOvBj6Y8XBOP19JqxiGCfxpN5iu/0+T2foaASIwfoJkyAFu
ygjhlEvEUHI9Fwc/7L7msgsHAZStZJYs8E74pqEW6odEclvruoikPjMLS9ya
mhasyWFgVLfe6RJem63+XQM8cVXXcGXPVZbrBcGhvEgxth8ebBEX3o70WjVQ
uS/xiU4ohhAjMrGsOBNcbtdoJdz+xdBAr5ym05rUT+uzFpfcCLBv5qlYADhG
EpAROKa9GF7/S9ErvO1b9EW6/U2C0Mhn603eqjs7SczXMkYjALNOkEfvLW1E
g2n8qHqvmhwKDvbAjUex0FI7gBeAzgGmkpjePvEST6oSr+84ULepwTWc9vhC
okHnXl+yoDuzHY390fOfAWI9tEgIjLnHtjxT3+0mkMrEJh859t3R14rhf2Vu
7tmY5OUA8h8LtARNcQKs3snsVyAwVIXfP+vLINGFHYpSeZjyOKoEtf60aZK7
u4mR0niOSMJJrAi4wx+abBB91KMHDXDxC/7Th5ajh9+0SUr56yUi0y9cqTF8
Llmpc8WC5Gt+qQdKNEqKWj0EjGAWsuY46D5yvpGL4goxpsuHVtPqmrjaa+7h
cRsP06jyFZ8A62jpmG5uXo2ErS1xWxbPZQuEJ7EOedeB7xM8LGngZqFlyDRp
MhCVU7Bs7RTghGyXJfmtxYck3NOVNB8OED1DMsa/2HFquj1991mt0fXL7vY3
azTnWa2jGrgAGW98G+6ncpyT8Wldhr03h2trf30RhXsvnN0EVq6jnJNbOkHZ
0/NaDvcSuPVUBVgm6ayCyvKltUr+RcN7CU/X5rLe1zOAwAWy0+r5vN0cLEgm
y4GBW5cqvdgbcJ78wI1GjSSMoueC1Fb+XkQj6P/SHSQBQEvQ7IXHSfANjd4A
2LKW2bycAXh6ctRJzgWcq4Ormm89u9utrnePOFUCTTth/aCPPGMjmDtTFapK
gHTarsI5clKuJmPK2SS5q2WYLRxdUTAs3I3NYe3VpJHPEyyOzMCHF0QZsUML
oEGwvTDd2zGekyYBvQyaIvbViO6ylRKI5v60ia7HTBv2CzJ8TlJV7Tp9puVL
o6Armo6INMSt055WhI41fKXj+ttbqh2xU57CtrKOfc/Sn+xNXfxCdsf5Z6Tg
eJj1OcsoWYzm7IncQH8pYYTM9dcdBwGA9xk6Aw6zg2PCq3A0YIa7/0XAXxzi
qgKIt8bi6kkjlapTytQ6s4VAK5fbdeqU28CVEpJB+eQN2zVnaFhutUpnB+kB
FmI8AKDS7A4mELGLSU0uwbeEHj+1Nfanx3etzYuTb08M0ESNyYQosWNYF+5h
wal1RawhL4z2kxsEE9M+Ch0x3yNKrdHzhhIv9RZh/HxD63x5kjotFTdQXipp
+dCeopBdsKtqlG+O1JeGRt6a0p2NQDtLmMgta5kXL6Ko+ohSNc1UveOkejpj
uDxrFOGDF0LTdmjqkW10XZmWVahqnGmvqiEWwwx1oJI1fscgHMLxSKvmkP44
Z5Vl0cLDohiVA+PIgDuL6xsYUW++l7XFeaNtPSlTnzoTKxnumLhe85w/6YVZ
M0KbuLb7I8xhWhy2ojbFjOA3T41ZdBLQ7XSLRDHqhTtaXfXtIiPP6/09BFd3
zX6xSFIwi/VmII7HvLb9925xjl9P/Cgg8X8zr68J5hRkqJm5AHGSN490nRMG
D2+6QyUGd2GiL0oAQlppr953Dbaf1qc9hBJDVtRvpuB8cD4ZurHJCxcAFUaL
63GEtp8+3J4Hz0HE5T5skuY02bUYwyrqXybVbF9oZxRAorEBhAnzxJPDZaI8
zREDQbtLc+CwFVFmQP1UD7+ZjjUddQ5BsttcK5OG2OG+NQqjMc2ulhm7gYE0
+LSzmACaTTRIGcPbcuxhoV24bKuL0dqUorBXVfXqE/pScuCGiNKmpeDCUWQa
ZnZpMWPAIQZF+72hFnw/KSgngwJP3Oapb14L6ud8rKsV4Xe05pGs0mTRWCrc
ukgCc5QtQRuj8YI4pHwah1dfZSHxYXV/kABYrQTwrSaJdkj/gAsX8z6C/PEd
hTAQ7LaJqziQc+6kBBIOTAEampWBan4uvOFEUS4x3SsC/YYATCL1Yfg6/fr1
TwFmgIs5526WO82qerGaPeorCrt4r5Ky8yNSi2Mk8BhBenZs+EoSgImbPE9d
S2zJADW3uuXC5oYIv2a68F8jYb71+5+NVig2eWAZANKvBQAzbikf5BVEfSa/
9dJQ5WfnljodvGgSnbAah5w3Ya9rLs0q0gEHO2zRsPfbb72Uz4ZI5K0Q+Bsg
zLrDenaGN4ceqHHMkGmyDYq0jgS9cM8fVa9si4IVx3UJdCT0TUqc7MtQSFzA
u7BkuxxZ+BLXu2THLT5EiTHp23899SogBebF0oqhEDQrV5o1EUhHtAmo2HJn
bXaqbNPIsbCRhYT0rGUNUu0RzJh9YViT8FH2wDPThzl9gvYYiR22P2zIADXi
Pd9GhY3RMCYpsV7Aa1FQWg48v/JmbP3KISlFnSJcXU6O8TKmR5y2vVj5CW5I
lBejAwRvCtUDQR85Dj2kC5PpKoz9qHXPb8DY56m5Qc8B68Vk/zKgqCFogW2/
cm3RsiF13XBUyU2RvGS5yXGhwR8KOSqG1tzolV9T0t6tCR74cbOX3bKJPAjS
5/62tMeqixk2HiRpSpYL5dkuvhT0HhNUPOTftnsg35rh5UOX2oQ80fUmINI6
tlo5SnBUCMWhSoyiMesf3P78rFSYThtba5E8tsgHYZQMijFJjWObD8Wk6tMS
nUrY3pAEr/1tXORPLHHj83HWjgvYqNATp4RWuPz2H2Uxx1t/d5q4uYo1RtV5
2WU3wUVEYXXdXQ6naQRXxeXRFki3Tu9fLKaVt06RFFanMJL9HGbGyvdDP4w2
NG1ZxnKEmtv5m/jeknXErstcxiPcncRXG8CaZjYUvz+vDp8+5J/WxchMC8Hs
U2K91rnnGmX+RGqhuQo5SVe9qasviQIb+BcQbGYrLpKUZE2xgQzWzT+4Jw9I
mlR0sr6O5N8lWwqKwN+ngvWKdVut35tluCOnLU50JW14g3znNnTpdYpuHqnE
qOY3bzULMUI2qgb2zWQru7skxSbbP0i/yF65JQ0aMCjzJmxOuS+S2+gPJK45
9/FYW8ApuqIJi6T+vV76iAEdBTHjvExYDXBtBnOjcfpimcipFqAWyKLZVfRs
MQI8FbKx+RuKSX9pWN1C3kEgr1zzEGWWP3dNj7M1tydQ1XEHF+FDTxgWLnPg
CPF1fuG3gEYkIZ8SVrZW8oo2ZNjo0eeetmxTqNut1nmrtyKz8vDZcQv0VbMe
A0M/h8NVyNUmbBHc18HN6YTHFrcDhSe8QR0lunC7wEpkPnH/ABA+ytjIIPzn
e3OjVOt60tJGm9b1PcN08WonmeX21BiQdF0SZaAIZ2xQBMTHn1dy0BUct7Sy
MbBmzKpWRXYwvYZpGKKT8iCpRi8aplLx1oBMURySWhzrB1o13Di5uZey4HHc
CDVDx61PDnmyBKTTx9cCzTx++RaFtgHUlF1xJulSI+molX7Ybp+2aWNGOu9p
FRmCkPRSMWGzneGnTk5j1fFTgvvwoNeELAYu9n/5n2P2a+y1u8d+Mskd+ZbB
uZfM8hHR9mCY//xmEUT3n9Mkk6kH9BLPkKrry9ZpWCprkw211C0aQX/mxGKW
ZvU6WdQIY5a53TKh++bv4woUICIQ8yI/P0e1g1IdTNKurhzwDsfZQH1tp/FZ
dA8jpHjFer+XAPDqe6t66JmEeWgwzLNA3b9GSvQp8ucEDqctprbq9Bfsllv6
rlp523hXA+sAzTQg6H9sUjuejjap7NPWMH9mVLXK2ya1CLFUiHktrsHmBtSw
D3UECoyZ3z3vj/2LU8BM7/BUfZCqCecpoNa7P8LXqJlEmqgcne416roOgqqS
JbaOVJ+w89+oHUi6/6nKeoJZYp8FK0dAOV+Z3kbQo40jiJa2UwYRWUFH2F9Q
c5kyG6smxeWmV25tDKfE5NtUKdul6RIyI+nPrbH24gMWTDnP3BIfi4VFu2/H
2+aN1IAZgFQ6lQYmqRfeMaJwBKgtAjizTEwWyb9PfUbjvgKCi5ac/9yWhx/c
477g6+UA5VB/e6tuvqHqb8RqUo4FAARPWgYnYQUHwxanuzZHcpdCqNVoZfo8
OQSEpz4Jogiro+nCyZ9iO+X8c9aX41RT5UFMRfdl1IgKU7cPS0xMRyXEa/e/
+Py1lDL1213f9ya1B344ExxPx3WuVI5xG42+kNnsUh2T3/yfq5dd9aealIcY
SPQjlQbRe47hxt2MeU+ka1T0mf5r4Z5Gi3XHoBWXfqTE89GPGgn2+xg8Tp3I
AxkakUICv0QCt7xUP7f0tC8+31Uk30FQjAwOE6lwg/aIs6wuzRbBXWOACOhf
2Ktso28Da8eyFXRVJTZ0287O7ww4iGBbWwSn0ARJHrgOvqyZbSgZUkj3/DK9
ex3dX/pVCEMOPhi2/5xoJXqj9EWsntVR4B1Vfn3Z/FWYD9HeENfZu+eGd5HD
acyw7xnC0GXV9Ww6Zd1JJacmj9Sco7dsa5WCyN4CrXUdYBy/ZDOEE/XY0H9e
U36HqSlqEiMWjdBFmcNpDE5vMh4B2PQ3kEILCwgGtPAkGxHNdQrVMtXXY1hY
7MBhmvJgtMybzwJjvm4B2NMMg69vg3tMQr9PzaSLRoMSSoYUQw3gxPIJlPoD
0zWO5ZrOcysaLPVD2IJuQph6qGYtsrsrGRwO00XToyKhY3QudDPHL8t2Q/iK
V++jzAb2OhlGyBKGORidlVXolakkKD08oxIqaXT5JZ2dHsQjof/icbAwejHx
2CSWo5egTec9sWwr2ZpnHXNuMz/WkfFR/h551Y9cc2bplkLr6j2TnVyw2r0A
acq1WiBtQM4Rikh2dUWt1AMAzvMqRig/tqDTWIWSEXtOR84Bph0V6WeedFeA
gxDhJcd7YeHyZKWCuj91x3wp7AIKQxc7V3xP2j2vfEs9ThQc/f6CfH/ouxx/
LdP2ads7nByAhoyDQ4P5H5MSXhG1ZXPayeezzqQCd88PheBk6Q3e6y2P4fQ4
Vb0xVm4p1czD0NzeC73UqrVVNAIRuHS7XhfEiIyAW591Czrdb5DhEYrCEyCs
AZ9scygcx03zqTUaIhEbgEjJOKiiSSls6cER8Abko7WrxClxgyA/YY5TjWbS
vKCWxJdeO5HAUO7oJgYZ3Z8rnadGp0uOwv9aQ00GV4/66L4fCkfbxY5SiqnE
hW8OuuQfdTpcyFUHlBi/HfTbpl2jRkAKfaSgzLDQ8xQz5mZcTJ4ioo/WCeHG
M8Cp+DckI9v2EhmkMYPdoUvZoos9PWATbE8bqCeToNwyhqX9UFL6deRbWLGV
0IpZQPxaIDF+zBR6wGpfSbJV7Y6Lr5cCSSLaOx3t/ae2EfadPBjyL7nnCdwe
GZFFC3NdYQVF47ZsBSTnvbX4FyfEw4MnuS+py7q0VH6S/EkApIZzrXu1aiRt
WafGbHRQ855qWl3JZ9v7ZQkhBuq2995K/VlBNJUiHXowocIPuUvRy3Ce5sMl
IZDNfmxeN3DuwwaBtEBKtBy3sG2RyUSF0WLi6tpXddnSL+K8FKgvI2NCw4s7
HP1xZxGVtYrekGWwynreRbU/qca6/pGC+X9TwuEmck1TOeiTkVTDmJNtjyVK
76A01U7O3BGpFrvxhpLgih+CsdPyvynVObXjIpxGJl++baZ0Jx9dhiDo/mOM
TD67w74kw8Mgk0eiSMPuTmntFxxi1UybOCyAOoeZhg6yQcN1sYeyLrjrPdhg
ww2kEC+SES/1XNpvSDrG4GXLzG4YR6GyQqiCpitcRRBuEWM86Bd6QqWKKcFm
Qo9cq+agT1C3vIPl2B+XaV0COO0qGzyMvtnklAq/DY2z04zeAUu/SvIqyqC6
rTE+GrXUV6qvlhYHVLNuBHNYVV9cU/U4c5EvzSrwkvCCZdKzPZ3Mjcv6PAP2
DPIhzwq9COfuTsbPRiRPgTqyB4KIn2WI01yNiQeXgCfcqkhJHwRDr/5DzGz1
gkZYZlyFnZ6E6k3hnwgEe8ezoHOSdSPaRmvkSgk5ChLO22nzfglQNak3BnHS
gaUGfYI7bCaWvI4ahc5LJMdDCFRNXgkLkrNgMAurd93kmW+8zLpybXgKwkAg
zaN0/4iBBuafK2F+SbeoYAdbXGYUccafYgRyY2yqi558b+ChPIuDSIfKDnI8
uKDbFSOEue4YgxxTJFS9CkRoJ8KBKSstVfCWxIha859Mz5YwL2UlggeA/E30
GellJeVwqI1e5V2xcq7M6YQQHPJkNIlQKMXi2EPdAgoOS0eRKfF75K0Z0Ub/
zFd5pREkQpKYHmOzZBy9LXHP0S1eV6QydqR6ijnhNMaOsqUm0B7i+kEvnfwv
1yzJLTStFhgWDe+DYPvu4QWPkxkwEqPjQvId6wI7oWlEc83GEOtwV4P/sISU
zUH4JqvVU0nOdlRUjT+XWb0/D8RsMcfFM2Y53Jo8Uz3DuHEzczmBMMEoypBg
lEqxeai0enoBEYnQGVPixPaTSbHEnijrPkKis+nj4vaymHF9RS3zhwXdlwIF
Jxb1/SdyL9Jg4Ic+IRB3kGdSQ7sJpH/iIH9Sqt18XrjUFzKzNEoap8HqH9xS
/rD2XiKKBljr2ODiQSUTWgCxKxdGwKOhx+ALoymnQZ5kgJPuCkCLeNnVi5SU
c178bMqL0uZMXj07xL2Sd29aRFiLj/FUXRJk0tgKjk2H9X7zC4cbsuDXn/am
SQvVSkhmGD6Abye2v1w37mbY7np2fL5IVhiYoMRLlBKv+8Z/JaafSRu2aZQy
fSDNnB21jFu31Pa4RcabcPxqJGQ9XCwdGKMRfG2RMWwfnuaOsZkCicEJZi21
3kuq5KN81urIPkUdlYPSdRW0d4oQ6fjYvbsRBfQ2EMolCbWda+WD1rYBurF4
TcOG2GlnlBXV9ah9ootHv+ITVuxLdviD9QcVfHPTS66VYaKeFBNxKbre/Ban
hniGVgavlTjqjeiH+QAMry3xWt68x7ciCb9R9fJ0F+2oykmt0rNgxk0q0xdO
fytMqAs2e9oEecto1urtx7Eusre78cw6YibCt9t8rIr/hIO1XEz74ROgJ2tM
6KozAoGlnMnxQxUzLM/nqYVGDEUbmQF1Rfr+Va82JVjAfxJn3f7eJSzQGonv
SRzZD58wrvtfkjvFbjYzAuFOSUctkdRmL6jb8yIZohR/YRYkv3x4rijuLvNj
iKtwYTOWmHWpOQdrB8jT4gIkXgdi9oi1dD8NmXDHrod/XdUsk6VYZGBYBNbn
5XHRjui8PIAdZaMm7ZSNi8Wfj5/wO44kQnfeLYgBRaZmncIYaYtW8UTuWI2c
0eKl3Km2oX4T+IoGH7qGTwSOr9wooNw4jW6JQoBfCnvlCExRoBPUA5g8UX9j
fwyDbilKZmd3wRN22cW47AlI2g/kPvGGLhNy9jAo4kGPZBw7b+y9WO+cVlve
i2JqOc80FwYi9zyH0yFLVmFam+DT930iQokodZ8I7b8bYk6y51jyp69SMWSz
sXJvZIC+q0YNxQPt8BXsNFxxCMlfECT1W8w0sLdioMIaFhl2ilaFDzVmIVjk
mHeblBQA6+na0gf4Eqv17LmLJuIp3R8Oh+FUEKOGOH238FWeuk834rYb8RPr
MyacH7F/F47LKyS2Ct2q3r4HlJ7AKpdFkpfxKY7rZHaIR+6iPFjtJKKYa5Zq
lAeXIiW9K7RqerfOFuhxNwLArs+TaYL/aQet7tSGbacP5zJJuPiUEcTFmXWG
yTgrOgMKjGjVK/jd5jGxivB+iuhcEPNT0aJUN28go2H5rgYrThhqmrsyEtmM
QL3Vqra7ekrVR/cgxbRbKl1tsI+vkGRX3NxxhWxRcQ1XIh8vI0sympbUi8xB
rfz0MCPo9330ztKZV217vpKaL1Pgog7td+qDN5lln4SY8y0Ec/zOv6K5z3IS
yZYZywFmBUehPINkKedd3PARpgnb8W2TMn8IQpaly/S5HIKoaoi1DeY9zswX
X5w2urk4c3AU9G5XJN/jMzb1iK/zxnVFUgAOmAAsM6U4H7yj84+I0dsUh/t+
LOhauDFi5dWn3K8qo68UouFr26ud1LnHNJywkLkY+DK6Jl+T/nEAcptwIN/w
pqK7Py5QHi73bAS9uPoAQfy0yaaO6nfhtiZTbr+fUdMpmkV5FUbWA4cccURC
CLIDonc6vcqvuXLy1j624dr2TpNt4iVMhXAhu+8ErKIF4IZYUeaddzI5Pm1B
zZBwWwa7ToqZlJvg7rgKGZ2rJUhbChXoBc1xLdQY3MqrSvBBzdSwzdwHFKGX
p7OnyIUbPIeyQ/d3QgYcxCoJH4TuaMoCbPadtQVkmhfga4RKQySrSkHngEVZ
WmXPD5hLf+JBXkPA9bv258iaIwCu0q6cflXVP8Ca0a1NCaY8nMC01M3oZhKs
Gau8J5jrvizC68z4igPNBAQwEdquSMCVK6MXi3jkrD6Egir1awbp8xs1phMC
ktXDbtGFo4sxa2RCXYpggSjhCPicnRI1By0bWXe10EI61OOwSdCqVKAwDtlb
cir+6lbTzc6nzq7jOTwrEcfk9JTMLVH4HsWDODyTpmlldKhm7T6YdWmgBUlB
HustNf44eG+IWuSPocrS45rzp5lPNQ7j/CS4WOv/VxvJ0vJC3HXyITtEoQ8n
8CdaANdeE+Nern6uGdEkWdE6d140wI+OrRK0Pkf6vfLQXp1wSpkKK3LqJetH
9D71+SV9mAtg0hYvCr7bOlVyLI2zQcVA1PjqsSZYevcvxVeUW1154O5KhTkZ
1NFFmsm+fmNdZPm4OxqajnHcAZB4saQsJscxH+ehqtXr4+0t/VsaL6vx8dFl
cyTYuNrIh6E8ORArk3ExZBducFnlOMAFQP+41qoS4BtR4WNT0hiRe04c9R1B
bt+oNGS5xlzKY0XawqRNBVYUx7RsNRhj9hmdGr0DawVs1danfXplxgkdaKXx
crjsBTUxjYbDt2MEpnxDFe+jGQA+AnXO7wBdJrRo3ur9Ak36TPGZnIzMcpkq
vJYGjZX2tHJx9lO9jPNW04NNkTmRLkzyAOop7R1zCtpxR/oOzV3hkiMHhn8f
VrnBcGqDloTOML/RPVSthcpCcEG13UzsntepzyzeFkurh9w73Efl57EaAeD/
6KwaogKmJFvhrjBgHabMc8+kc1VxElVUg02HB7tLsLaH3N7HIR0gy3myfw9C
ES2o4AP4eZFETw5YXfaheNP5rzhoJ60r5S7U2fxncmg8JwpfdDzcWZ0ZV/IM
v/02gGeT5HAXCm85r/MmX+6T4JPa3tO12xQ3VF6kcUCNucAnHG04uX/DUxXG
Fy/jZcLE/nZBWjuJNaIZbhuQ5FSypyv4i4668XLJSdOPgfP7uixbmQDISetn
d/f6KFNgpHtkXbqkZf4AkiAgTffNUkSZOI05st+3rG+K33gzeRosBkkcLBxT
wJEsqOTjT8gXw4q2hJrWjlv4JC3u3FZL3VGRjqgz0EUJfj3/O3rUn6Qzum54
US+CqZqpWRI3uoEqfVJ8P7xQwEJJ4gRHGpl8IRB4SwTOINWV6C9D9aqRTTFh
JCiZU9YYF+5V8OtTy35HsBJEsvv55RqMgY2Qs55/MVAGrHu9uxzzmAx4q4bZ
W0hD/h3X8yy/9Fcfwr0hdTo1fUKMxBY9A3Q5IkTkewpzZrKu1QoBBfwHimGq
0tPFtBD8b7savQSEKg7hZkv5ohkpnUAmcCjlgXwTRfMHvgJEavIJpNvRI8FG
VcNn8rUyNG8U10svT0npUtH+SfPevnJgRkviOxmFF62tPEIF7cmHgtaLmCqk
OV4PUVyP3NnaaVqEbVJyIRNuc28aJPv3HIzfSinkOGi55pSzmXqUL/Iyrt2F
bOdYuUy/ugtgFvUdLzLVxQWGHZdpH0s+o37GNcSIwgvMwGPfdVlwXfmnsY4t
92MF6f7hX+xnD7qiPtamkMEHwdpLqTQI3hnGfBh/nMpgk2LaeUZX+UgL1RIF
nQ1v8yJuBO5bUzXDb3jQK0hifTVz8KPqUuVFV1aXzrd40ZaDHDn9FIP8ZESR
0pAsaU5CzG8cueyFZX8VjmBI1HcsvPH+QNxsVSVQrfjGDEjuwNquolEsa3v+
JdjpSfY/8iyo8VGVef99GH1AmmkCDBvzZYhjcBzgQYPX+2VHQli3cFHp2gNZ
kfFrcHlBfOBrh8hXKeDRQ5i5va1jed4p25WNhtq8RP/OOXp6Je847FPqWuc3
TJPDrVEqZYrIlWVvLzFdlBl7S33W/dkgOb7vxRRJ4RHTnAvhTVLAvjPpx05v
5izYUw1IA+uDa3b0qoa775rXdt+ILRBpag1c8D0weice3CjNPTCB5RrdfCnM
84DURDHr12ivqRnjh7aymYfCXEGFVwe54YYc8YVzVqchOossZ43RvJX9DmIa
fq5GcrrWkE/j/oh96Np1JuW6br56DNM68TXZGtBCz481jJj06GUW1zkyCjwu
tEvAriUmaC5T9CDytH7WhcktW39wUMJ3U6icZRz3gtBsNbsTn9XRpsxXLWXu
XhGzTilkK1B4JqTxQ1o/g6K7XlgMpqcpNmDBNOYoAnX3UwM3vlSAcEEd9R51
+3mi1jJxaHyX3a3n/D7YV1weRY37vDr2+4CpV5U0fxxhAGa9bZ8iYd9XFUC2
1ecW1uZt0yIisdndIxbY0SCWLZpeNL0dBOqAlaaWOfLLa2YSm/5u2W+mZ3bB
xiUOZvaopOW13Xz/9iEzXTMrgLJU9PxIMt34Hb//O44wJSjaIo19s+0Y/xDG
vVbZfv6+Liq2HQSyXsfOvv5ZA0hYfsii2q6bvTpFUrITDhVmikyuQNBFhfQO
PpEDLupE3ha7FpFIVt8qA+oP0MTOG0hUlcI6cakXen7ZXE7Fer8tkeQUvo2v
Z5K1L/IPnorqaOQS5hdXjXZqrjgXp1J8e7c5UlBo2m0yxgaqdQBnLNecm3N1
UJMl6mPYgBycBRN/zu+RrNctme9cw4RLPH29oxavzXlLKhVKUmAxdH3EKdws
J7I56qYnUPAEYwDtG561zV9whhPwJV351qf04hKGsZSoeZpW4a5TSZHoG2T2
yNkypD1cIGhdsZRcsmnfgZUL1jaUgz8y0Jg5zF3t66ihefNBDsSvat3in4ut
/0TCimmSrmwSZcHp4UsYcd5wnM/uKJ0ESThHB3Iilo4wKMD+sT394lm/sbz+
slsdv1TtFNSD9kVr0qYANfPgip/70GIIBLeGFc1cjafBDlW4zHftn7D84Lln
hwzJb6ZIXXaUnS/gHpKIB3XQ9NftW1wcXXW+ODdaPXJiLhzJM70sF3bcb7o7
DXexynnWlW92oA8QnSObe4+3xykg1Pwjd7zTvGVKuT8SAplMRc0VXkP28Rpr
0Rbzblw78n1c6sDUy3729UOCl0ZelUr2/eEZ5QN6MdgpGwSZFDzQe/V7eOd+
Mw+sqMCIpvyqHEPt6mzLS1j8upqdcSdhIntZ1spL/J4oKmKvDf3MFe94C/Xz
vNGvRrSqqFOSa2HiMWbIHsOIuasvjBqNKP6Uj04HS1FtklMRHoY5mUeIjXxf
oIaBgycjA4Sib8CxQO9GkgNtilDxrjwON3HFeIH2ObzE5S4iKknDnzvkMTyy
xxkE+TROrRe3plwpDxMp/Cak3iOwB+aa+kN0VDZejWMh4iGDn9AZncPeQ+C4
sbkKIcTJHerZhe1FO0PtPncmt15pgxZCX7jda2FW/GGBIxXJoOh6NIkiWAs+
/yWJq2yKDaPYb3/6UgWJlI6Qi6AlUk5Elc4wnSBtBdZ5r91WxZ7t5kO5Bz/5
hcELn0h+83QUzxwcuER80DMAMpMZX+pa/wgMx+0ePzwkXxUh7ViiWXJvOYz/
iVxHLo7qfyCRXjQ88ZhTf1ZuIxm6fMRJ2zr+RK/33a9AClGZZy64sJ1o/JEE
JFKdRVNfj1oFz4R7hkjzLVJr1qLZ4AfEQXHbBDDmLPbadKhSnp6blDcpl8rh
9u4YecKwzDiJr1oTS3TtRfLZYSBTlZ2Ud/WHflW6PdxX8+BlDU23wHofh+hr
L5a7UllpsvRbkzkGXPYk/i37iyc8Sb9VVamwHpZQa+Hgcr6QG9Kw/nERBBTC
Luy+9M86+G5wDcbpv6cUTkEQuSwZrSy6e43j08rHDAXT4fG1aTg1Gh6jjQMP
hovCFxcB5PQyOFYrXr4ntmlcuSJT/wecBKQQ+wKopfQ+3HGEGFay7FsauTx9
NPUoHvxJUd25mwKLNbInmRjxcp5tyjGCMFKOf/nJ3mJnCmh6DM8mu4lXV7UZ
t3I20UJWsIol8Na5S8jPgnWaN2uHVzOXIZZNZPMOvJ6kcyiAt+3txC+MmpcH
QpkqnmaI8ooSscZ/7X8+82GUqRYAVcMfjTVv2KMktMYcXA5i3ZvmnjRRsChq
KKpZwfOuFeZ6jKwtcFHQsuudNwFVUtw02pKDGrzdvn6lUKxTE3ozeU4cIzRG
D9c7E+kawi7VLKM9HAaqt50zOg8JcaTaWyYRRcYC79/0ei9IFyIRLfomR3MI
rIi3+zsCaTVsRiEIBzzxYfkU2ko74t4SD5aNaHOM+Rvyp1vJb8yfQQ4WrmFW
y0NZBQAYic9OblKDwc5kCdD/GwwSztFTiJUENumYolZiNL6f/F/8eQgmaZSj
OO9XU/G+fdd0SwKwejZap8+vSbjqNKgW8laPD8EEXHPp/Rc30hBGnXtW0gue
su7/SbZ519N7gkb8BaBtNot/uz54xspKymR7+dy20xN7KAsLkXgmu/yhee4+
hOcnKguyeNRvdFgClyKWTfcBUqLyho5/h5wK23JMJOm8cr0qg93DTAP7WL6u
4NADPHbFKx4/RMZtFmG7hDXIuAQSFscOIEQNJm0LL8g+tGn3JFweYU8s+Vdu
2MHqiK5E5osDqf03UOZmBDvv+wQzSnd3sS8Tz8CjGrOui4XAQVoVwbwSDb+e
sINU8pcrbGrXRvBBlJKhuFV+aJY28LxPynGZkxCT3m3Q1MGqJ7xjLoR6R7Wa
QCXhD+STgOeE9rvTzA+AhNq83jIdgQz3jcXCIMcbaXur44HWcdH2ZZ4JlQfR
RukajMgCS+8s4z73z2zhQ2MmZrUMWIfp1SFUg5pv4HgUfzm+DYV/k9yooAC4
bQ3vxG5RJ97vWsRADBY4EVNo/9GWzvIp1zefZwnpRblS2w60puEeo/sIvKAC
v0IkYOqMPlmHbD6puI5imBiK8YWZnJQdU3El0i+/4wrCJSV43VFvgR5/KKr0
2/M6lltbbAoTRTPvw4YL/qlV8Gu/BVVqMYdwCWzdyiO1UU8gJZBjAMVDQ3jd
l6dRV3l8pofHramb4VjJcrxZlz72aCkq9iudYe8OuMR3+Gc/xOLtVmDLe4hD
wmAfx2wsluJgBc9eHvgWhO35W5OuZTVKqYRFkLmVA0UGjTg+IWWY6n02BF1V
hwP8lreqiyKycwmKgDB4tB1e44i9LtJ46/ZHI/gnApd9BK96SOvYhlCS6itF
SZS+Cd85/cAPyRuFfHw2Mhm3BXyvsIUtBWRVwtaRBr3NKczJIvC8MuqJ9+4n
6XuUtHMGM1ijCkGRtYQrrbx9chkJqtDZ6UNUTBfe8WACH/DFOvOnM77gbX0V
en48iOEd4qK8vggiyiel1SQSHFEH1/SBLMpffpOJDCdmKI7uo9MuTA1pD+NQ
JSKfth5Z+Ym+VJBg+b5Om2szNmTOr1xUSmr6GT62qm8cCXh105VED/T/gZg8
WXM9IuO/p6BCcmQQQD1uEsn1Krx71q5jnOl1ssl97k4gwIaM8KsgYDvNS8xH
FQy1uBBtLx1rRwasnBlXMgFD1/3bRjG/8MERuEvnXcq2RYdiOGDovCBPgi+O
d/cGIPJTEInXm/yp+ZuWmwbPAosHgVTmleZ29Ct3CmuKlCz/xifZCJsRZBEt
e8YqR5eTPkWPRtRA1bzj5Y6nTHk6uypdMjJW+ImS8J0eVpR4dpbJZvUTWJL+
ju514q9cRs2xmTWwUrchphf1zrzGLtIJRAM3h7cqb8mAvbePoqSrjHTBN4lV
bj4PqrLbdPkj+e/8MSqnvgXphOVhkoZgGGLFHhRcyVc/ilXSZVJtKnqPRN6O
fXqUqJ9UnOFmPoXqofcBWSw7FLgar4Dhh6LlYibRSvBTlnDJdyzBYZygQbo+
vVrbPxgD8zkgTfmndYLTfq9p3j02X6bQjWyJftNhJvmIwFBZeYkSXVzPN8vB
NtNp6G3mLNM/rsd9haS4X4TSVHloJ+3wFKGFHZ58Rsk+jehurKpZjOZSC8za
rmAqvJtdKsyANys/uV+kvsjWp3Z4YOjqZbeNVlwWnxT/hbzM8yEQfgR7fnfC
njPtpqvlqh2pde7WzKdl8HaIo5646PpkRmWnL0eLvkrje2KNkG0rCssJxe+L
QibTGnSHpB2Lb11w7XsXw6Q+HknZ5cFZLCfzvvEErrZW7YhA1I6lS57wxXgs
PYDTD7QLhMJ2szo932QUG5eBxw1qwB/O76nZUOnr8HiNf+DtLjlAVDvoY45M
Wby23KjysNvmW7x4ccz7dyRFD9LX0ZU5jRmnq1NZlJLyxkl4TCBPlHPOO2u+
oiYO0A/RyWKcePMT30vBsz8mbgUY7xn/qa2Ccsbdp63MDZ69vceZvlrUWab4
v5Pf878XtaXp9C/ZyMd4+km4AikVM8R503LC05JPiAWqll7wQ5gEwNnf96w/
8HVYEp3n/9fv1t3K/W/BWY0Yzzmaqil2Te1OfS0tHAV9oMM+iNhRliik31mC
MDB9Ih8EMR1rVXlUclneKIuJZN2BKLdnGsaj9wes6YDgBbjpHipR9RTUcjuN
lCuegLaSQy+yDuWKH8LcuclYF4fcpSkydEJdFPWV6yeVUNY5LEm6q5VT+STv
YkfQbT5EoQaLKhz5ZgoHxz9W8RsD8u+gYomtmgPAyflODVeddpkB0ltqWjvx
uQLV2M3UkDjw/zV40hrxFMXQd5L/tIbS28kz8AUxek18mTY0rjHT8Q7Iuipf
5Z0AT64V7Kph555VFYk+yntRT3SeFA8CjW7ylYK8E5Sf2ypO2cNAeRqbyJ8U
trJfuqV9fLtwvcg6okt9A7D5OBLLftgfVJ8oUoya5vI9MZjOLZkIO1cY66cp
8UTLwR5Qggd2JgFab0Wnq65sBNfW6KWBn6SLVBb7h5f6SN//DqHQRKXhQqrR
+4zUovkMvHNBn4Az5CjtXYq3raPFK7KKvj1E++cctuFp61Vh0TzfD6RkfV9d
JnLDNMmk/EauCWhtV3FbnZvnySDl1NR8+LuubMS7cnVwt+drye5uu6pBD+V/
Ca6t3zPns4orvKyDJdPXrZXDoBIqtLI7BcE2ID1nyOjhdphKp8PjZvUHKTKj
F/qBb96m04SbQLataptnvCQqYuMcoxckhxgsq9nEZGSj5LhL/zdoxPvADv5F
IgX7W6BexwfkFvB+Yktn7XXZKRPGVNawjaPoj314fLCJkDhfj98b8zuyA8zm
PVk/TqgKb26o7Sb4l/dNi9+1IGSYWQSR9GMdwNnzGsWheQiQNkGvNZNT3HZw
eiMb5NshXKh8jFPq8iArd/StjkrPxLMbo8kCa8E2VcjPqLwz5w0E3lQfUF5k
miXTMxSEbDhJER0hxS7NTun614IAIbv8V7V6ZXEq+CCJyaLG3g7TW++rNkRt
Y5phzQINQ4Cn8IG5h5kjgxAmNN+bj4efpWsrv7D3Q9imxzSj3KsQD/QWrAkF
9/5cyjftdIU0XfsTUR/J5nbZrkRCKFUuH2j3eUp1Iun5wCHbPigoZkktOBTT
8R/pmERKSuKvsJ3cB0uIu4XTZlbl3lvhwoyoRGzey5G4frqhvZDu22LZOQIH
cizinNMkhZU819txIx5uZSDDWP4f7EyMc8yBDfuu9j1ybzV7qc7AnU8c/UZM
Ob9jAvE0NJeVeSFyhoDiYgS1w4XsR+tDxVpEnXTLWLVDHWZtVAQPAJuyKAdm
U4Rjdlix//W0/tjFxg91rrGhxGNeRGm9x4tqKmVk8aHCoKfllpfWN+/up67B
XB5UMgpfYT1Y+ppv83NvmIxJfi8TTpAXeaS2+Tdc6T47q7+H2SBap4vbTtTs
u4gk4iBXIzu3BL5VQeHaHOe8EuQH3im+Pn/NmE66vgo88rJV6DGhwMdQHtlA
WVz9CLuBuTY2UE/D7guSfD6KB1TU/lnioFVUtg8RdSs5VEc9kA+ktCer+kLT
/MhISRfpbo8LHhCkprJ9MKYP4U7w0MwNHI+Syg6FRr2Nr8pehS2xvsDP9SOS
gpm3aA4wMQ2bdpFsyKHvd6Not8CiYjgy15q3h6NKlMCAwGB62MMFPlVzE9gq
nJRzAD/h8vdIb5Bn7MMJitIUX0N1qZToTpiSLAUbTgXYmGp1s9csjMapl1Uj
WOk19GbjtKdlvOxBrsisSoEjuLG28O/U5Nb7BuH+2mEnyOGFgA6gqJTJyMDl
obZHrSQsQGinhKvVmBbMMNRH4+XTNi+/NtwLWNdsKR/ks7rGUhOPJWrSUaAv
u75oEBFKXdfjK4YUJ34heC6tX5bU8/R2Od6MZYmJ14x/C5iWATh5I7dDVNeU
vXXPVC4v54JXlTwKF1e5IzsYwBXAlI6ciMiLTzZE7qEGz5jfiQ==

`pragma protect end_protected
