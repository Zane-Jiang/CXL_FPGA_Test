// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4dpVi+ayYc0uEtVnJcjwgZgN2T1VPDhJZTmXPtSEbM3taNypr6Xv5h5XBFRlfzcb
i9zcs/60RujCM1uy1W6o3Xbqtp2qcbWKjelqh5+a4HOR1ywmXGtyNqudZRZrr0bg
GOqM+uS5SR1bnCbjtpZ5gCSOnP9MoYaPlJ/4mlVRtc0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7376 )
`pragma protect data_block
7ECXrHqj7xuDl+hBxqU6hEbKbxrvU1z4CZ8HyRWtBvK++Fo7HOycclZ7BTIFG9RK
31Mk1p8wH4+mLjvhCVj+k+hyO+wLfFsetsDDk1p7Jc2oGlEGvrQZ3PN8NL2EJ0tt
LHshu+bzlhtISr059qArEWHXXf9AtGHssUuM7B3PnrI7sgTWpGvppYdA3bh4a4gt
wAgfy9o5qqqzwqjHcuKDc3jK2B1WGfwTNZe1otcibrTEXqhmtQymz1zqxeY4U/e5
mtCHVH04ljAmqqcvQHA994xZV1F++4zucUj/y5WC3KRehSS+K2BlTPeZlYoHMYsf
Iynn1ySLxN6ym+THtPNAyp0tkAc1gUOmFrL3tZ4jZGZfo4xo/DWYCTz0bpJ0tHn/
57H9nxEdAO+n6bOTKmi6k/3JTwiaYSMThbWqQ6w6bRYXcC1t62JUEDYkF+ESjhHk
E0fdjNWqE+AilrIWzPve2WDHeWyKL2+JuNreKSDIlchbiuPEM5EL8bfuPUWk+jUG
piIzdwsH7UR/0EdtbP+oZLuNHWmiLFB+OydOHe/tD+gdbcYXOFSN/CHB0XgnS6gJ
TAXvvKp4M25p7Gv58qTzyrluxlTY+rb2c4DwIXaZIpu0dyNUPWsJbE8uQ6slgYYT
4I5X6ju+houkiEMOCQHnJKLwV5AMJB46xL4aFgG4OX8Gqzl4bxtGM/N/sqYXmAlb
3zwoNck4a0ebsDNDICb1XgyEPbpPoZWwOnK5SmrJYgB0BmGeVIOcPnGHT7Oj7wb2
Txa0iz/r0tBGcLm+Wgzpp0uE8wFli2CswTrU2sutIpmYF+8UFqT/R7mOrNFQF5Qc
FTSNpi3LbJLGJ9K5GDVoXOKvc/JJyF+EiYq/Z+KjaV4mMN13dHj8K6Y6DSNwM8vw
nWoH9NRgGCwScPdEPYCLZM8A3bfUZyhQAtdhDWJWalPnxOmxvoSdICizxj6vu27f
t3++D/mUaqUb9CvVTyha7LkgejMYoSIvI48RNeMgPD9YtrAnr6YpwdbGs+4yNWgo
0x3WhNU2pxwI3JyWNAi+q0+WxKfDuj34VajwcoBebAtPEHvvU2kwIq/TmGSz2KXP
GQqBZZqoDpzvlN8Gj/Po80ZOTAHD6PjXC2khYp/uegnEH30U6QZSaWju73pzKTt6
G75Zrv5voM+XFsiwPGTk8Y9koXH7XsN5FEY1hV9k6mQHEwyn2X6v/LzmU325MWhL
vIgaZAalqdro7hcxWhzmD2YsrdQJJggX+FYkDnriw+Aw042hBwytp1DeXY8cJvXU
MNnKfHvX3x0ikau1AKq2SnXnCpzinFyquYXx3fwUaS+tpksVQC0N3MjSXEs2C+Fj
Kmo130U+t8ECh+zYFrkaxYPMsQdvsxKmbZv/feFghAXIwGXkLB755nCmO6AyA99e
uAtPMbpoe/kcBs29UMYvJDcU+fm8FdPccr3WdFHzr38zVsVZgOyMcFGo9uaPFua6
F32clfUaO3mggiQWe4URoawH/q8fgJNqR1J3PJEnkLJxy+OtE0y0GX9MyWbM0Z3N
RdmTY0ioPllkTsc/nqtMohK4svG6/cWxYRlPC6X75fXutTZzDdCsD7tQWUIiw6EN
tG5X0Fq2PooymQVU4SMcmC9/z3rtnmfw5kdMAbaYegDqEUSlrqGLE2rbQ/Bcnk+q
5CI7dxM9G8/d1Hp7G7DMVLDDkZBp6urQEjcxJpVxBmDOX/XHzzJPbWWhrlkAHHOZ
6Bo7Ib2F9OwYbrFpdWjULd1sxr42tJ5/4h1zfKD7Vovu5cTq/dr6Vr/mm8X5EQ7J
SeNeO5RkUwsvqSnImj5Gj7thNH/Sp+Jxzsvbx0HwRetZ2YV8gJr8t39+kevgXTXt
DSOy3hENBsocmIkCUWjtTvGm47gzJ/LkCefcn8w+Qd0a1C1Mru6PKxBEIFTfh8yR
xfIjLdWXN91UC5nFgjC8XySYb6zpSH6m9khjxn0yH8mPd+lYv62lQ0/KS7tyQ352
/dFhXabB8yzfnDqA2f5HPg60g2OY9KM+V26qmdds9rzhHgzGN6K+cSEE2H+XjUtY
Z2LYBbY4Y5toeTynmiU2n1SJ7Xakf9WsRQ4vDZvc3DH4gs7e9eMSzSxPCDr60bqL
NNMcmAlPRdT9HAFBgmy4DTQRC2Qhx6utOSmnIJzJWUqNqHGetTyZ/rvnK/CJtKbb
5wPBPY3fxy1SGk5w0ljZUd0zc/SoECJfmyC/W6Br8OllXwODJzjkoyZ+CLQRnbS/
5BmYZ/Lap/NjFtkG2/Qm9pZ1qhrQzTLd3NmaOhaNeKTluwfSHNrNn5MM0BqmDoVD
U0A0eES8sg4F/kpWbLb+MPGgcGlIkv8TdcgpelzsfnKAfE1gbhSjEFRuVXU+7sMK
6rHhwqbwHS0yTU9Al3aTEXqK1ADHqgigoC8b10zJkLtD/hpoapKR3ZtTOHh7V/rL
uKfpQxICwzM8eAeZhsG3IAXiEYb9pDQNXbHySN5ZI1VTwB4S+HyGh+ibJ5WZ5U8u
zK3gn3Vke8zFgVbbJKHRrtmU+mmtw4VRjC0fCg/2E2/9WTnP1YAeV4qNjOBa5yWU
1MDvgss6QTnbE72EcamhlsLlhUWXEKN4umls+/F8AQQIv40K/TI+HtrnRxKcqXos
G3tiq7OodNqkpjvrYIYVcOJF6o8y2cMGdBtggbD6f2sGniZfGTGP9oNzyLiApKtw
U7COvF8/CyqWaQdgDTiBL1mWEpjrLZFW7l4mcOh99VSbj7u9glCp+NnpQJO2/zzr
6pSmh+nfJgIq1+JjNnA5gWwpEnwksSo+QGpA8RMc+qsLl8LmUddDNw3KngnjW6At
43pXbWnSRbDKoK7TZ1GyAxQ5P8ualOQkAEK0GaX2ibKdRAtw5MiXnJO79HBojbW2
e3/xEBFLpRqWYIhnxHj1hUZvECyxkZJUD3WuFyiHjiAl+VEqTOw0ceJJs7tLhNj/
mDVkjghvWAEYKStLaZ/wRhhBCRzDtJcSctlb1GTaKl51myflwoMNIsWbWNU/R0EJ
7ORPAt5bQJ5bM/b1NZu4gZ1mBzgzioQJ4r0f/892BEtM39P6H8Z6V8IAuPyzg0k4
L8kOmTk6tz7zsLg7CiSW8bce7r8EcZkbIUorRJ3BLXC9gDjzwmZOZJMQc5/K0b2X
7vDrVAtoKph1p+Qf7D86AuG+by5Umc+lgZ7ycUu73VcqmB3FMbODuVg+8RulwFC8
aIdBxvRAr6ZcvfTdLrC+BbcDe1yiq1kRu74eNWuMxLRDTo0mYANvENK8IruKkuI9
Udf0Qf72lZ7KxM3H3/VBHWk3uOG7ygtaX+bd1QVM+ZnncgI61ppxzVU6Xjx4BZbS
GY66siNG31j0BDGthXQXJmape9l0or+E5EdSNHwI83IQ9pibmiwSADzh0rTLhjcl
TFq0A4oFXeNeHenpE3evioXICCE+ABn4sGOX1CuKu4Janx7MaK3fA+x8AAq9dONL
kdVc9NdtBIeU3WXMXTjzSfg1D2pD2rV7KVny9Hvvnm3vqad3AdNg7uPP+ylFEBuk
c6m9x9L+ka7LYLto3BAZ22pqYe0+WiRLAW5GqtSS58zs3he7iZ9HH4f4EbmxE2Ja
4eXNa11oG94oamPDniVFRb/nNW7b1tC11CL+xqn21SwHf+rjPhLHD89uIgsxYqxU
H/E4xFbR5Z0QBsyB0eYhI4PRA4lx8a7YgP4hP1JPc7gbkJZEBcvTfsQ1vT74zqN4
bSpDgqf964V5kdq2i2GIgrAMoGcdwLhh1zxgp06ekQSa3ApAAeK5azUDS934TWh4
PKjWQiBsQhQ3E7Kb9IN/7ExAgo/IMGSeyYt7bl8G4ZlVIsBJoD4cw6s32XfjJw/B
Ron+QoMUFO/+9HSOMKKPQHIG2v6HVpOJfRY1+8X1d0+D2Wr4N3+PoPxSfkHDFDBE
5m7tNtpGIDZl5lgMZS6KlZHmzhh4a7ro9GucRC010eI2BzSNyQ5rm0ntzI/A/urK
3X37dfKvaZQgKItDmwfA+X0d3CP9Q0OwNrbBgC7kSbd7nJERzQMdmzTg/OqPBpKI
0mwE+SBEi6SlTK99+2pEEvHqfRnhk/5rKTdYU6WLojvpVLdUN+YoOZjbxxuFe/10
036rozwFgn5qVUaEwzUxPj7LZO1IAOgwrqPkRAvetjUYA8lcB9yqMldsIwMbRdI8
1zQOuD0i1L+/s/aPoc2JBNIlbL60cNhq6LeDnwDEODfQhAHeON4ntwPoGVpU2Mrt
AuedKPXdlvsaiBGEZV+GJNsbkxACpPRHS6Stl3XFddQB8snV05S3/4n2htHtBiys
T+A7lr1GFyiR/72WFIuvLVmkJJVduxJgivqBkpfjPSEUz2QaHbpXKrbRlykS70Zu
V3kPt7hKk10fJSYO4TA8Xhq88YiqGbJMCgSXumNAc/Vfhqunl3vLERROrlUkP1Dq
d1rXQIf0dOZ5zLpyuAEhOiatF9q7XccvB0QZurjuzxH5rqiIRLKslZ0+cC9m+Gln
QZDYU6Q8JaGD6ESBVGOmDFlipg6ON4rhoAXYs3MBfWIdQ7lJtTJCGvQnY0CSvR7C
KgmWONOzNSXWmr9YuhXsPT1OuMBzlwdPEIqVIvCPpL5RjI2suOoIYFYMaGhTNrYB
XBJjFHDj4rEsnSB1S/jAylJ8cTyxev8eKrgL2rLL6wVjEgyq6eFQbKqCyMVS8NHA
OuyD6ounIFYYra36ho1wY4OVjNWiOYmWLS1YQTKwGhmDrADob1dA24Yeq5pQchzK
gHPEPssLSkmENGAxgdV7z5ZwIJjlrCvGiATkyXErQ+ZNbRpWmo4izwmmm4qqbtPX
xu0MqP/Gx3voFAMIqRK1pdT5zfYYqA0zhgv2aEbTVUBJA8zFZ9+gE1pjiV6hzKvO
JBpw3cAvhb6Zo5flwMQm+W5F8JQqrW1T14dFCMcMAo8D/guPjfpC6tTNGKjtHX/Y
Fcd1Sni10UVf4IQM4Jqc/0q9Uv3+DLuBRl/mwLN0P1Gz/bRgqrfnsgXQzT18qOoG
CkgboggXUwOtMlZq/avPT83ZWlQGZugSOuHj+yDq37soLz12AeNU4MjL389gKWBP
hzAl+4R2hj36iVHDeRa6H8XHiHZOg9YFC70hnp1UJp+1ONrhO0C58G2+fZ2DcYXz
2cEHGyp05BpEfqLpAq8dhVl4Z6WLOScQCuQy+sEH4cPliHqi/vZxfFpQqgWhgSKD
5mpQEfG+bCZ2znyg5dLvU665TMT+tE0TacK391fwbnLLx825E++083STsVnS0XAD
VZXeC5OCpN9i2zzbq0B7A4lLYb3HWxVC/TmLxtkEkXH6Zhs6oPKtuLy4b2apWFPR
sA3NbvCoNE1CATmSiRPur8I96udL553o+1xXiBjp9zBA9vLNoe6OJUUtp9teCDOx
QgIB1vcIb4vR1k4ejHBBy6qmBK1TSj+K5QTiUjqRYiM8E0ix/IIWhJuUAyMY6sxl
zwFLkGYDpWi8tAYb9zBuVSeCgZVhEYQXfNetBdYehlgLdSPDPbcT9RCkroZZDTZV
MRWWALzvqmEy6ECXWROnDCjorgrdXiHRWWtFkoTDP5MTwOk5ku7sZMlrhhSHkWXQ
8jSY9ZoqmETy1uuFbpVrZxkG2tpibVaFJr4Quv54G4BLIyyTUPo1i7SeZmdpgDQc
/0YSkkK9R9YTbGc7vMFWG7bQy8TLk3sM6tf30Q06M51MEJ5mikucbaBk4PgvR7pL
Df7BUyeLrzCx84BUEoItelQcDJnTXwMvIC6xd2/sWscsrcnRGrNzCZXojk6g7l2x
81NRzSWFCYrLGrNcrgFY+9f8hyM8u2tgplOlZbVCUB1l/6XE2m/f/2J/zE6rGxoj
03wVpMCv9MsAGJzbIymyRzcFOTKa/al6QUEmyXbcbkVbrw2Ic/rHPPPtQtq9Jfny
27V99DyH19GELPfeZ3Gkhciwj4FcGjIHgzvUYW+DKFbubOrD9IJb+iWovj7LJMnn
0vcK+yNz1kraAsQLpgXuhLdzus97stSGs4d6ufR4PiY5st0K5kCixFmx253KLvY4
hLCOAZielHzdzd1JZSEXwk1oR7PRKF0Ee/tW7ThlKTyzJ5S1YU9YTE2se0wao4SF
Ui635isgUaNwFpdxk7nt6ZJ8nP2j/Ipal0m0aOCuzokiHq/YF7JnRReZflZ/Spqk
TwPCUglpPG8vkXiFRYTaL+5gUqQuvLCMkceEQhAHWuHqJw1Lxpt0osmXbegi+gTM
wkEHbGi9OnbNKa1RBE8nHGLGwqta5MwrSYQppxa0uHdsReOZmSKs701xqREEnwsf
vcv7T2aSFu75T1WK9iqZnkdouXRrYG8N0c5aR6UjLwFQu78O+CfsKg4TmGTUVrCQ
JrSwiRNwUUFUTHwKpN80GW9fr/z/HhLL5ZiFsvtlm6Z0vK/WqgSiuF4sgkXgd2Q/
tLJylmDU/6iZ1eXMqu/waAKVH+NMec1YByvTuHuDanxhoR7/RcObJq+y/ZhsY+VL
7qfSOkanebqMbI/zs9dseO187VOUbw+pMFlOrL7YYqQ3VmytEoAlEOFVOZRtn0c/
fh/GN7X06cyit5V/q4x7AdNbngod2yAoKBl9r+qaIepzOG2mcoTkOP6stFdcWPKJ
pyePMwHUyZX4kGS0ZsvAseouvQX/bx6cB751ZACp7cM+DcFZpL5xLfQW4KVB4Qby
bVLUa5xr9rIGTW7mVZjU3EANDqcq+mgDyri/LGyIgZ9FToTZ92o0jqL7jdwqHluj
Dg1iGM7diuCUF+bOddhthnIKiYFV5XOYvdTOEYSjv9j5c/S3NjH6xeceUUNlaWs4
p/wOMluE1XkA7pPd+l+bPNrq2b6FvqKfH0kUDFOQnityH+SloBNzcE1/OkzHE7Wj
ClFWbn11KLFGJJnCOXlvuO+YWmxaEqylr3ZqfpOmRvh2mFJLt+UBfXXFEOxmmJL9
0ZzlrI5K3u+WCW0wNsz7ck5WJ0b+YgnHgME1Yu+FrWE8Jtdt7MM9NmIiy6W8Fi4z
YpHFkdXTIHuOWyxYjOdcTtKlIxIbTZz2zg9XRtU1n4WOs0+DjE0z3DydkusNlkXc
0WI6f2kJJrMAXtF9O07fbnfZR2vpKav4HWpNgcHCyCF0GTYyWaZM9uwnAFkqjr4i
WerAvLhpRNMwutO4BxKmCNRoEsrWMK/uJo1wik9/9no1/iPD8rAaZcEnMxyev0Uv
s5cj3Swv2VJdKbcAWo1KZoo87d4rbsyb6BwqcL2j/7gEuBz3pvgaVw1wMLi1nLO8
o2AMYZOeHY05jn1/6I5E9oa466jv1VstZDAfC3oWBimb5UizIf8JA1WRHrzVtis7
pRL7XzKKFinD40THKXjRLO8+n/Jd9gILMpsHpkOhSX6FhLBHNsPKscTQWM9FYexQ
GZXv3KqGQXFk2lzBSTOcIHU7B9zZ0B2ErsYYRlJlo5//PRs2E7k7bhS3MiHaG5lI
wqyG/zJECFnqJLqd7h/49bXJP436fCYlFfRn2dwCouD6raptrNDpnAb04iz3qTzu
xbT7eELG+l37qljrlzPYOf9BkzdQK422UZV9FOjCo/NhgGhYxzK3Omif4Z3mI/ua
IRhvjbYQm+L8GoVQfXUbwAo+sWEKeybZcnh8TvUk2pjvIDTQRijDZuSsJn6cjA03
y+lUaxaZ7ENHGl1qvejWkbg5dOBLCXCfj0jzAM6OHgxurJkku3FLINXjRSMk5Lkp
nzNdVHclvEc+dPxN4WYv/9/AATFdiJsZ46tlkJiKeqcI46tS5cxhSkd4763Xghj3
1gSSikZkj2MAlfUuBE/a21wN27UtsIsjw2wNgE2da/1FLVdq6dCCzOA4JQivyn/c
+0ik9IddTvNqUptu6C1LrsIwebqUomGzVTKIDaJ5QIUrfN/EEJsUP2CJO15CW74q
KdO7Tus5LZH/ffEsgD6GlNc6EHgghlUrEdZJ3ywu6d9yRZO057DA8a8q+CDVwOcC
rXnNZlynDbnUNPemPcucu4Cx7Cu8JBWXSvpbEEzjNPZFwq8wQpn5Lx/PGg6ManVi
go3t0CNvgs0V0soHgezeZGmpUWbLteeFbrJiaaAe5yafJOwUBeuA3iGgLsTeSPSD
KKxO3dqFaZodE1n05Rzn+VcZZN8pz4oM6JKquoMFY8Gryi9AM5bYPR/iBCjMSmnC
pjgkpPzxUB/soLuAVmPqK4cmul30PQwkIc0WYvEOEOUKhCiXEHeK1RYbVOeMbtAk
oJR6LzpX+mbH75ND61CdQjlx9MxZvR7VYO97X/HPMs5K3LvzZx4j8+3AmTsD5tjI
ddR/EGI7UMXJivUV9rYlFFdK3kMjpIAC/6Jy8oOuyRsXFKbPl6Yfq+YzcmcyOiig
+JW2nJ2Ck5xtfS959BswyOUHjt84Rbvrmvu+jAj8gx7uqpBDnk0e+cLBCBzK62wE
8OhaTWK5+moJjT4atZsCYDbzzLzPTWP1tlHDE9J1bazWeMI/VQvQ4qjob5Tvz4+l
laZ3BXaQTJOV+qQYg6dSD3xYHuBtsmIugIf4AKbGEatekXfJ/NG/SkFGZUYbpCCX
AuJoBhvXOK0l6h6F0Fo4HdP0DSpHf4m5aP+GoYWfRy9EAwtdCARo1dp7ErfD78hR
RDB7hBk7lZBX4IvvaFn6fAfzcgJu9nzTfQq/oVfKbBY3db0w+d2ydadwkxA8c79R
nbDxsYAd2yaATm2utQeUIr3/RbgNHzeM8FDgUe2RfdZDTWIFg7xcfVGfTnbQEGn/
1iUUIzqdLrlhzQlfhxDmmpKxPMBZ0M0Ay0CuGVJi/5wRr9F4zk/AIxA0jR/R/ehY
19wXgCLlMFbMbiVjGUfrj+KpAgwdU73ZlXxHROcJMZdEp3TApXV7XeI7l9Q7MWtC
f71uJXOhN10zAM5S66zLWSRlS/A4FtZ7gOiIQuxcz+/UU3aTeau1vuGIlDxjIoMY
ztj+TZGP9iXyk6ic+P/9yMLpC+YiC8vdGSVEC8642qTKwOSg37WbG3rjLlX3s13z
xt7VjQhOZ3IkwseN+ogT8AIVfZlZrVQpioSaF/xB50YBFV+DuRAvIcVc67Kgnz2C
PuGNbIT60bdaMOlHQIjTuYN/0qM7bJbikpISWDiAuGVTh3E6EnJ2zdXmoQx/vo26
dZQsyNZ9OXROK9KD4xYMMpcEUfI3vkiaMUFXnK4Fg+S78OJEnfrv13tjoCMDhNSb
iszDi0ba0kPaeVvsV/7EXNq2u7Ixp3+kh/8OOLrVrPuCOrMaUqFZ1dzV2nxG7b1N
LIpmJtCawy7/hsaoux1BN7TVaOa0KOZSvYn9uhu8E+VlaEW9YQU/BVuRhbBdouu5
+QvJl/g1gXeO0j5cIXUoC5v5FyKK3ErCkWf6iUg7YqXdzx16exz7dl0hVUmhA4Vx
K/sL/Aoo1e2gyR527KT0c4AKMwMM1mCsQMqH9JgIrqVhNBbooMb3uvOnE+DE1i00
yf2FhLw63v2VoIv6O0+G8Eo+OP3xWGBpxZDkDem0tM4C3piJhfu9Ldt8EMBUtJdH
ayuliiS8DX4MdRr07ipYsDtxsiYTdwg6uvqfPNpy1snWv50tjksKwoi70tqjwf33
/hcbNYJRKKxWjCSs5xOCo/R1+uchkcZfjRYv7UARuYu1WBfzE+PePLzrN1IRuGjO
0s4isgXxg3qJmGFfjmh+53+OQo8z87a3nALAUSoR003hMoYGLFcrisLEBusR5WnA
qLw/HYPUKncxiDyNBlJaNxDVWe66DPzNmKsA1X3IuVGUtTgMS482z8Gyd3yvfebi
ZCMQtWSaYEFhsF9a0LASSb4vd+jacbNAPgns4+h6fJIajl9sQVt63tASb4uvWBwo
NVKkJI1A21fAMlUQ9NmA1+4mTI7flHZ7whsaevH8kXk=

`pragma protect end_protected
