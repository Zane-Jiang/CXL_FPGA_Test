// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
OykgVWqg5o+sqA2CwhAG7NxNtqEOFby+cd6SidzjBiB6s2MtuL2ARQenvUatBbMb
GwqoMM6xPSF1/9e323Wj1txV+5AwDGSV2EkHV1U06ALry4SQwxmQJEQzUk0JujoN
twu9psNhvpesqscx6cemYuXpQCWqf/yVrj1+ReL03wY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5472 )
`pragma protect data_block
Fde2M25mB2Gg1vonc/J+lvuC79bVfvPVFBjdK1BJCXN/b7erzeRv02I177xKbRbi
R1AplOmGyYaEsLTxssv3dzpD5o0Qg+ynXCsklmXDOFMivq8h621n6YZsHt3zYoMd
1acpevpVdD2Z6ycw4cdqI1Rrb8M99K1iVzhi2rNfw3/ZPrcjPGnX3EuqapFynmpc
CVxPkxGTJSdTwpN6C9ZQGvDE6akrLOvE8BtZFmEKqDKL1qnhKJ55QgYfov9brlOc
TOQVwULxbT4EFZcZjhxDKXAuJA8xqJ6hkDqEztVV+QPxXqPC0yhDFaae1bLUjTJj
G6kc70NPlR0R99BRiJt7cQqOHFF9FsKzN2A/KDFgpgllOuY/6siSfBjaWXd8TWTh
RzXUQ5tkb1wU27e/7taSNrnRRhs0TvMwQ8J25qfSXKF2hly+YfgHHzoVQd9eXOe6
/qJnBoWfl2zYIhbp0Ja6ZZ1gJ17pqH5wucpUBsqkhuMpXcP3PixUZBTt9kbGMFCV
+oZHE0jasn1vq53ty5RAD5cXyBHe5dkVZB4AxYd8GJrLWz37/eAU4d1Z8Mkf2rLZ
L1s4LuyXfVDusgBN/nrRmTKGTWTy0FSP5XKgk4fZ+UZ0XxFnrTIOQHfKuDOeMQyR
ALAsZC3C8FU+941m9IEOafsz7mxgE3PTlfnpgeFhvgQq/TFuCST+sNm/IGOLxY7b
eX5bzfF9udsRWr+zaD4fqDdgyV482o70skdJrWWPB8YAyYFmK4AD78Jf7ieD89UN
XIqM5rho2JqJ0F+fm8CGPl1N2x8tdLcWCQxJ2W6vkx7FzHRgKknNKr8RGObEg4BQ
nANQDo+Pr9mp9/A7A8eSFL+5Wpx/hgnfrq69VA22MJotwPu0Xv4eqRljB3mJvud6
kLRmgwvdWvWpNIkxA9X8uW9kLxiIUtw1Jgqug8op5I/eq/Zk1USVqb4Qp70pFxX5
Ou9Safkxx+ylPqr9qopby6KXR6YDcF/AKKCJCADvw4UUwwWi626AUbSOL2q9bhsy
O/KvrLPQ3J7mYn6zA89ymcFpuHdyLk9v2bg03oc/huYphQw37Sj9rhh3UmPPIu+O
2WKwneYUAljzgVhUkeSWJcHoSe10drcAPcEJEU+oHn+FgA7B+6UV+hhSLux5bd7T
icZFwVl2c+c/R4LRhF7GK4abQoCC9V35ZHe1/2zQJtc7+X8Sl1KeyDoElHciSjRn
ETEaupbUpl+JD6OqtnGLvu3tuP+PUxbCH+U71E0JBTwVJpTwX0hKWGE53fxbo70G
e15roo216tctmpGJICBNpVgYFtDy4aasrlMFBGzLandAJd1IM1XaQJvYoXy+RYB4
mx89KRfh8Ob9dTV5JmSdP23Y5RZZ2tRk072YWvYLHZaXJSZsIQJzsyVVa8ijKSUf
X7ZWgBbvaYPzukW6zgNdJ+S4aimqCi0ztE1RdSrtb/tDqLLcd3IV6VC+QLXwWIok
FjFcDUjdR/n7kyhrb+jMmV01fNym2+y6c+3+Tv33rtUBKP9zunEYUbgGqhdjYz5H
OQmbkxPhUV8WFpUQEs0v/VvwBPnc5JAIlkFo9o5c6FjpxxfPD0dUMHSluvhw9Xl3
dH4BGoG8c1zihmGvrWGqvmxKIQhf6Kx/zYoATmcbXfTrislFpo/F6XxkYGgZVTc0
2Dl5pP2El0W7SIvN5XsmDNF5qj/VcREnqmZLdjV44c8Y9HlSKF5NGn3Q5XIUx2XD
zo1HDcj2WvEPRP6u0u0tlq7UUyhlGLrgvQT3PfTuLvXqYWHyTS41qDB5+1t9Yx+i
ELotv/lYrDuW+ejgb//OwBCxBQOqg1rGNCc+ZsWOe4at9e6g1Y/lysQ6d+grj0Mk
Mveu+9Zkg4UQYxP3nEEm2l3r6Lw1K2cSEQ0JnMBQfAdvyIMRsLfVK+ICu9TO4/Gf
WlHZvr1RPXsKN14c56i4jC78JAUlky3G7leTmL0webevZQRJoI9OHMKzwN8D9Bvt
LtdtXW0R3ookdiGxUF7krkCRD9dQPmIXQTgmFpK1IXs+zmlXgJhkkg/FhCYU5Dmg
CEYMnOhDAFKebqZAPnNIeUVSO2sGsomtkEEo88ctCwHFVluvKctI6lP/PlLkCUML
krb09OJnwWQG0akfn883KUue8gYcJuYgwfY0FT61h7q+ZHS4UmHSF1RiQCgTt0Pm
GyGkHjPrj/eH5ld/pC2CByo8hSC5j2Hb1HaOclAHz5U6KNRmblVTv+kVG+7I2GUs
b4K+ooD9CMwDLJxTIX3YvQgHr3jx9gRi8ni3dwSX9Dmifysamv0jQTUZsxB7YBDx
TLc2ujddf3FyLZiM/kqg+a9LaoKCtXUgELNH2VJKj+1eSbN5bk9ABTsRrj0oJF69
sbXVkUlwdayWVia0m2LFnUpvGt6ppoaE/3VqRRORIDjqXyGTALANG3pjksd2AECR
BAU94duDRu95X3t77Ggs683UbSPgc268023vVBd4p0y7JVddE3DRbSDi0535EZA4
WlFaOBF20c/bknpb9a+HCevAK5S8bcrpt1SvQ/g4RIfTssSXf9ZFer7dZP5bYbnX
kipUKHsL1AN/hIVIwGxQoOodbMIpCF2FDdw+01vyuQWSvzHphv4XrHA09zd3FsJB
69Ee9CwdHErbMentVNFBNY0p0wuygGVV7F5VdA2Of6RhTQEa2abxVwcWwHjvgjOF
uofCqoQUB4v6alKrIii7zt14DHgZJylX2TfgnhDzLEpELsCdzdaHD0zuk4g2Ok9a
Fiy3VpdCiiJRbAPmwYL7owSx3sgo5BhDEVTDLHiH6fd0alF5JvxnVkCSqGJOOGjG
E0sfRFRZMb+oHQM6uOx1Um/B4kNRaEYITcJ+YDCJD4mTQIF27jiLi9ax64Bmii4Z
J3u+3F/umKEYI5Zh40egzVbQbNkyKCDbexp6F5o2fOQhZKlPCLII6pHizeVk8gW2
S63qVopyP5uvrbH31CrvEeWOMyciJSEkq4Bi020zFhf3+3gKooh+4wKGuDBD+trx
MLx/Z7CuyxGY0knblWgLVZlf09FayHcQ6FlcHNc6V1HIaCKqFCJhKS9PuoFPPLYp
ykh9NLpw1+1tTAZna5Hq7y+9p24ApgBkzlNU4vYwHVm0SD34gmg1ufGfYRIPTXN1
ZVk3pOpiwGd29XlBlAl1ufPKE08Z80He7x/1MnZIAMYC5T8gF9aaw+D5YdfCprBP
suclDGx6527uW2NsKxodqQYS7jxNMSpIiyaWqVT0a/8b8QM5E2QiTSZX4Y9jG+Ki
vEQIaHpF+PeHqSzshcW9Pp75HdEuah4RnKOf9wqIM1uCkZTzshtDjhwB4zQ66iQa
BbxNPzUr1pt4tUi+OJWJvJetWN2uC3oJ3IvmVQCVciu+uigdxv10g/S4aKtgBXGv
0n+y5TsyWOKQRorYfBmnUGCF5BqYTPFXSfS6BIzaU8/r3LEWxqoqKCJM5ULv+ejD
uqqIg42Izlqd3jpX+4YVN3EfocyOzBReV5Od9Rbk5M+FxFQNjgAHm8GIW3XGvwIx
xW1YrQGI70RPvy5lvjRol1gOqNSwCmdBJsPrmbdO6agcw/i7rUOddatJp/yP0rmk
xqExoKJppZos4dW8rozaiTvRVPSupmcJs7TDvBk/6WZQmtU3k8vB2ZmaQ8SK00MC
DTr2W7hQ1/epwNYrZLm7Y+2wHH/KNOdA3C47rNMtSS3soIAxR12AvHsI+3BJwdKf
ZH0kl6Q4eX7rqScc9xcmUndYgziGr7rVJtDjkm2eX5vsAFqR8suvNFW0bJd1HS1k
2yGYVu3Y41MKxS3hvsap9K8qrmxLBEdK2pJXij0zbAPtcweIShXt3BrzszkR6CvA
ei/rxQmQCQjXnh3ktZSfjcQaBPTKGnZcMtLwwyaZTyJHCSKHffqhWcazoO7PPp5g
kdppd11IXeFvcxWQPEmn6wvVAS75caP1iKMB1evv0Vz1+wcntqixY6vip0bvNmwY
neoTLfDZb1i/fILlhk5MG6Iq6mkYPN4KXwghWTcrV9LoxiU3Taz/4U10WBVq+Qfn
2D3hO10YPUA6/sewX59sJv8BSgRbWd8P3dVwIn27pSYeeL/86iBTL+mtTWCli3TL
VSWQzXK1QGRVbxnSkLupixa3rn67HPNtYsB6oGBpP2i+EqY2xVaTSAA3JgRe9XHF
iQZtve6kBXk3nQ3KXi667LBB3N9jRtWoFPFmX0bz8oPZcjUBtmka2bWVRMgV87An
nUUTdt2qo8+IIyJgAnszMer4B/Nf3MqPOCdYfIpMHcm0OJwE9wwwRBkK3nVXskIn
fRbb3PJ5pLpObHjKkswzAz0PbZVasEVIaJ25w1l4kdPppRCbjPAzU4PdlAGWCJ9L
gVFFIYKijYYRH28JHw7F5XBfPGmdjArhCm+fYN/8ffNwTdyXteFd+K9GYNT01wsa
dA2X9JcYOL2rEvjLpVnsTEoyZ+SSy2SLFiJcLzs/IIz/nqPWPKKA92dwYHzDG1mK
goFfJ8bK9ABd51P7qfxO2zyPDooDameaVG6DRgmZCcip7OX7+vpJ250LpmIHKOP+
MfzAiHKt8muJkmM14gol/tH9YJfzH739U1mm/DXBKT4BtZWqzZV7nsRqlr9FQNlz
CfrImnWsC972aUrerqpB7lyHyArqvSG4AlJgcpgut7seaNbDmmpqKV1nqtSnti2L
mlNW3RN2rmOi9aQdDm8YtBQUglyIVGOT3ygpiJGRcE/u2rImJlv7NYHUstr90vXF
ogBP7/dDZXiyQkwXU83ElxdYfEcnzvIWqV2gtJ6ScgZMlp/ZXTmm0Rza3AVyyWox
u7EQO/rydSfm7wmlcHTgXadhX3uPSYFusM1T4OiX5ODsjyrhJt8xWzHgkQ8/hZs5
KOq/jjPQMGrORj2WPKR04rXu4ZsTUV8+b6CoX5IdYXvHSfWcrewHeWygs4+uTOTU
JWT8C61ySC1fL+5jk5w8EgO6E1y7F+5ACLF0C83sZcrUMKjamzj0NVqh6ZG5EmiP
YqRlbCYyzhNtLa06njSP9mhiEmxFF/h7rd8K5WEexwlTFxgrtuUD4M+QPYkI/l77
boziy9mvSvSiiA6koSsJNi4yOKMOn+OGGHigpHPt7DCkYt5uFpNXnDzbIE1nXPQT
PzmwHg3ApSsAWm65ph1RH94ylnaQGsa/vjG9JrfNUTly+MIe0DCBHovWuJJ8ymWT
PSPcUTnNNYa54IMew6VP1M8SUH/sZL7rEflSMPXsthLWkb0BDHfg4bb05QCl8r47
3TcRWhADlJGFe0ziJA/llkKap6qOmwowQNexMN1jSftQMrorjfqnqjR+qoDMEdgs
JKxUFm/Y75A/q9GUNTKg0O7zXi6W3FC2YxVF8+IRU+S5hs+jIiU8eN3rlZpCKQZw
+BFzJnSGW9rxc5846jkU31oio997uruk4jGNWxKtAKa8DS7jqVyvpJd5ktFvTQX9
L8q2G5bOhEkyvv+UXhmXfxbWBNsYWo/AJCTcWfe4dWCqI87Hoj/Elzv5DzwotgP4
mhZ7UGy8tjIlfgb7z9ivP6RR5iupH3sr11xn5h//q58B7n2ZD1psm5BuL241T9Qn
ASQV2TFqW+qHJZdbcXU9Z672Z1CfkKxB/ybRsyfZ4b4iTiAF6GaQeXPTZpRPwV5M
/FxujrpDFyZ+7jJnKfXymRRUp2oBwrodLC04O6VnWtp3+paJwVnoXyd5gaIReTOM
vGDGZbPX7s1fDWVQruCndV8ehq9nzrUVmQodpM0ItcnBQqH/giIxJdHnyQFh8qpr
mTRpUZfiThplg0k14E6MkSLw2Ato77no6QUGQVlGbV9PUn4DHEnY81wM5aNVQW7f
EMGOAcsHXEwyvgKfiM3D3GfIHTVA87UqFp6JlIxmj9BswzlpPnpMjYnwYML9G7vt
bHse/XN9YCELvO6rpsLAHW2cTl1wvW1RRX+WNlaPppO4+pM+LL3wk3bH0eWGSHoP
RGih8iC30wrDzAXJHSCMy9LdBJo78heVsReyrnCiUnH6ularL2LGSl7kxkh9FyGJ
39AsQqqXJASD5kztdvy/GK2IkK1N/vRXC8kr1VKyaFmPx1FXNaZN6w2lLJaRJQZ/
++FKNmvqhL2b7NiR0MXLYW1PkgzZHaa0k+K/C1jtqWH+kGkaLpdSqNWKf7CWcHFa
QTLN1iplHpXkTQnhHEYIBqEBvtFRY6qj78CnVNz/Ht/1ucoqXZFLrt/2wqL4pjJk
KoEndNpsxAri8Yv/VX/My/hi0xxTRUOftkC+bb6TVBsJTzxMEbItyZVQVMZIJ6ZH
y2HgMEoEaIeEgoaRjKMx10PttSxjrzeop2pKswisE2itjPedI+CjDUqD69JeIVt7
/ATNs8B+YDXkkY7CBNpzo4xQ1ivhpBP7797sLFTiwqxrGX3DHFDrogUZwlI1vVeo
B/kdKfoCvkm9UBDQwi9HlczhlHwvutSlS9AN07+UT+4EkL9og1Xskq8c4+rFu1kC
3TnlUmzewrs72zrYnAktKOVqNLG8GdxuBghno2xJTuKDNO60WlUeEEDBCPS9pTHZ
sstgyPYFqYovOna+FHlslwLsVPGed5QPWV3LpUF2TzJeY/YlzJbh8ZADkuzR/e+J
TbtTeHQ72+w5t7I8DZdJKUmjTQldR9J0NregVQwGX4Mu8xNE5Q8Ax57GLD+YgoXn
OHucl/8wt7GkW1X7Yfc5+bibsOLgg7vSsSHQcrV3xQ1JYIvWfCGFG4dwFRTC2VzJ
SiNyf7D6hga1V8LVpfhlN/6dT5cGfScxUrmCUthjzaqmJGxmFv6ZXcvv6EL/5ISU
58aPAcBssutRuwqfqMDlppygUc1cODZRVK3E1wtFEZ4fpvdSMiI9Ipgp51guuX5r
hAZTK7vXlbNxSjMKcRz+POUMA7+TuXh70IBzOemjLrfnG+Ci4Hm4SllA8VaRH4yJ
TbBM0SLlrchcMRIb1Hh5qlfrzEA1OJUMzZuJSHUTqROtnrFNeJSJWVOrRVcRqc6A
d5ioGTODv4lPVBxsnuq/Y/Wy5g3YpjgxggNxeQGanCMGYw3yQBTytLggU0V/0c21
NzzjIfAJNMydNuXaP0seaqkGhak4gE/vn9I3VSUceYZz3H+p27KGSDkQKFiHQoZ6
LX3mMciAeg2oD+UUBp/d8Oyk3A8f2NVE/pBQkJhwW0NGNbfu93MdfXQSi9dfKWCl
3dUpIU7DqQBcvi+UDn66lud/KEPyTcoVPjPc7+P3F30PAbbIJReIwaIst0G+oa5R
CSh8sEijtQOrim2ERscePlCeznvTgu7DqW0c8Xsl+uzzAv5XjnwGjrV7awz1qhAc

`pragma protect end_protected
