// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
OkxFMoSYNpvVwFtgzQ+yPxiELLi7TmPPp63rG/3YTT+NbnwP0QHGuPo4X5Emo+EV
rrsCWuQ7rmOZql9/u5oowWeupCQE6s6TNkfkEamwdikPEkaDs4ZGiz/m50l/CYSw
5BmVo/B2xrbBATTf/SqbmuIDMK1mefs79WcJejsI+pMoMLf7RTiL+w==
//pragma protect end_key_block
//pragma protect digest_block
Vd6XP9onnZiLenQBP50/WHx7Z2Q=
//pragma protect end_digest_block
//pragma protect data_block
SP+LfJ99chAGWeB4F7dQAtmhWcc4YGhTr1uExxFS4iZ0+cs/jncmntvG03ZAXa0O
JAEffDRtWxaOIoB+0B0zNyw0BsRWsPIat8Ut8DNmhckFZZhcEj5UMAv8u+Qa6gAO
yh4QKtq97nySUgxR0A7EAqPPg+eqoamDca7Tpedg0zJzWMHIj43t9AoGiAWsHG8b
jKcLf0kSjiVXGjWyEQHv8rku5FopCi1u0+p1Rp2yRMAYosI74EQeO50KURB1792Y
vyrwy3+9bR75VBpC+toWcsRrQzlTrw5oSy2ccNf7pyLLL3i+IOtzGzBfRHbT75rH
oRIw1U9WOs4/41fo/hsSyaK2DkMX5UnUnfvqdOcwyRE+3sqL9bizgKY9zeUhLul6
TgemvuWnZ+U6T56ybsJa91LSVRk+vJz77UOx+mMfxDCPOUBW59f+AJv7K5rKUpj8
os40QXqq1LMp+1uNUEeqs2/J5L9Cxbodc3Bs63+3DXt6lhQJetf25xITtqSsntmy
aqhepZEwIxmiu4Q2L8L3xTablqL41At0aBCFQYrtZakp4t9PnbOYDW2DpTk4F0O0
PZta12YUILME9i5/ivuKbWTttyM2GCP59FMbu+PBxHaNhEh3QWA1KH+u22tQndPb
k6VOQQEHMJjQ635qAPWr61wZYIjaryje3CqqZvM6OeJt6Suc3MzQp7IMnEbXlNip
jSO1XwvZEUbC2n3im6/ACozs3MwkqUKSl0OR7+GLOVAx3RSVRo64Fzc9iK8dl4Qp
2DSWYbsawcpqyBzCBDvOIeQWyO1k2J1gzl3osBhG9FIm8Me2uaikKJIaxiMGWuEV
yT38nGE1ryYvxJYHKu1d5XCEM4ke7uoDrYNWzN98TA/kbOmLhhEjgv0wq2+Rnntn
1K+/FBsMDNXo0cMv9oh20OeN4At60d30gZWNFaBsu8/lOoOyKKSI95kgY0Dvlfw+
Q9IhKJDtgxpj8xm+ggWEcGsiWwkyoy5CuPC73PwI85uo+hQWK8KAL75sq22hgJNu
oX0qjCwEidMX6u/3GmPOi6dLaKbOCpwQxWQ94PWDBGFw8PRt+dFR1qYG15o6xN0M
m7/1hlqy1q0KpcFoKASlY6IXiROwq+Ly9wKe5uG6N8ZO+dWmCEtwX8NAXEQqJWzR
yc3Ygt6jjQ8b7rm7YwWklN4dU3ZOZEZX315++oLBmpMydQA4bHuBW4r8NP5TlQGT
kvbcji978srv2FPzaN5XusOmiBA9btP+O7K9SyYOH5ZxkbwILohokUkXIC4UFB96
N0iMG5ZJZCcy8Uvjuy+77lE7p9jZMxiskJIodstHuA077FprX0XJNBOMidumAq8J
huD/s4IbSNPBctHQHfooBkXcCsK0Y7dUjmyDpxo7tAAGfrx11pNId/hcaBShHjPI
ApAFsuNZjB5L2f8i2VxYCEKfXKiIbyRFczPYkRJnl0u4ZUFlcWN4Gx3SywB7WrQv
8VAchvbCGkb87gHkCVVLdauy+HZHO2OiT0zLpp9AMETytgmIe9TZHzQNMWO0s+JG
dTCJscQUGKKxfz93YJIG2y///ZFoYjNCgnfKb7dwgJC56WaeAsXsT4wFOZf/b4Q8
tG6E2REmP3EYOS8kQyn29sNxw20m3tFrrwfRyqvc/22Y2U97a7aN8F5wEjkacsRo
tdxoJmAFLGuY+NTI7c0Ty8faC0ocyEZjgYRqK1+yVRGz78rZFC7qCcWHUzx6Hqp9
u9sTIRGNQkASTc7LtqyG515ZAqi0W4wf81Azy5HiEb0joBkQkXNFlBzVE5vgSNCD
PLyNOCy8ikeSfpPeAV/g9jSMSlo2lZzyl4y2jm55MujHs+U6fWUVsIqVUvgSYtb1
QffkdUaQc1ACKLxUXkVzLEi3U7Wgzpy/b6UD0buOzt2ZU5f/b4oZKHECbTrm7A/6
+mtrd2IfFebjudmCuc4k5yS9cDv1M1spFS5PUy8D/2e4sgZCUxL39uwgUzvrTfmp
6xt4KWkn1WqYwEE80ph9QBsvwRqASGutbc7kSL+tCn+SqEl2aN+De/RbY1J1EEpx
GJlQjw2n1774tnVZrF4wlF/MF0XtP4HVghGkBfCoApKLuK/bIsy5nbiRIsvWtpz3
jfii8byVoIsuYADlOW/tk/gt5I8PDyPdMG+d9fhGdEG9H6Of6EkOjRFdkaGAMTMu
vClbHTpxNPqqhlw+tpE7UKZ7eGiCYcCwanyARdPWLfzBpr9IAEQ3PTyBmT2Jt59k
eoCjZW5n4oRqxujP2byLy4An2Q3tJvVqfNkXa1lw6IGRVzbj1lNjRhhjpPl2qfeJ
JG/J0gvoqxn5Tt8ERiuiZrPJWtlpWl71s17QI7IsV3L6spZrKIOPdMU7JMy769tg
TOGwZw3jBvklDFMqv+OMSFeDOZazzmSGw48Be2ZBWqZiv8Ah6m8ZOh0z6OMYPyP7
y9hT4XsK2S9mox0f1YHwdrV7j0KUTe9ApfYUa6xjgkI6R4KhjaYHTGfkb1pQ0iFd
hllJWc61MhtVeGVIL69rZj5tZIIxfiYYRVJswMGCAOt6K+IgiEUs15ehHVy5r1fB
294K0fea+2nBeS/5TIJtEbdIgEVmBBdv+rrU1QXUe51iyNS4qHZS3w3hdKSM7uHC
xz2sQsx7bX+pO7Si3bkGxvVkQ4bp9W1B57qvCZaLLlAvfXraWUVh/CyyMfHU8grC
mWtFqg133cV6ocx//IqVdMrcf9n5eaJi6IFcoEG/ytvSqu/J8g6M2BqC88ndk6Fs
O/z5WATxhVq5mc+SYKDOx/vcipfGWO4ciW2R/PrQfUchkv3Slgx2MLOURZcFsK6s
B7z4bnMwgwoGvsi0BmSe4m4hlh9TsyGmH1zOcU9IZYZ+nDyOqNXZMRkqwjoemr2E
WJKZL6LDrypgQvfwj8UaWzRSZbaGlo2/IztC+foFBuEHBORVu5KaR2V6irOWMeBk
e2XVuM8Kz1h1fdQyWwz1VsYst86QVYwwrLyW8Txcun7g4e60a4zdy4JRcvZt0r0R
roEPbEfWVO8RPhBHvlWcGrDlMI0dymlFk0O6wla4hQP9UEkGh7Pmx0wT4Fh7//jd
XRBPvQ4zBYKhqe3eEwXYj52cT2SVO4/QHmd+IwqOQKWhUqw9jUjsof7+/BMdj93i
WDSKpjcRIE9wDywH9YMlIPf6Kryn0G+85XGYTaFVFp9aR9q9ui74Q6jXOCX+vOvv
9/cdQlPwD2tyY2lnWh8JdaaJJgis2/n82eD2E2517Dkht/VWCZnJn3dVkvleyf9J
mbYluzw+hBnIUGvg/q2cFzRgDaZSqHtsmSnSI8tW2kZWXwmIAU/iXB+Xg9/tJ+hk
Ewp6TzpM7Jrqlif5j5f+qV0xN5N7K39J2W2XZ3pga3ZEK2N1c2jKaqGPrfUO/HPz
Gk6gcdF+hfGGDWtRDT0lZ0VbYj86L/DV0l/mtuoEnoaTUEEAuU5cip6pSsJDE8JQ
p9pwmgMz7v0TKuvFTRIzAFlqGL2MyBmnjCptgippJXXlX4QJ5pW31uw8xHhEdjuj
1XG0FFVADFWqTlnnYwI/Mkj4J2PqxQ1C3Z8vn9sO1897bKrJoV4AzxHdpdfC/WrA
S2WSYfXE+6kLtxQs4c/uxKfQ2pcsA7ptOXkZ69KmXBWnPUaN0h/bAVV7cZsY0Baq
S0ZzJRTeTxp9iswY1o3jwTzt+1cu+QLOuibH+I2m/Kwzhw6Bm2gzFVjNbdXt4EcF
W+n6IkGl4ORSqZJju96DB9F2eC2yekZps83ZQ3kpauxIevYaiF33CcSSpFZ9cgJE
vjvY7ZoXxyTIR4if3P7a0jh/KwD0vCj73vfe5bAblATUIrp+0h46xNjvf37THg7Z
YyDXmPS4rVscdVI8GkSMyva8VdtUq5uMx431KjAAMTkUgxkKSirK4waz0Mfl0Oth
T7FY0tLkXahy1xNvHur5bJ7QrIVib5WtniHIqWANv8/IKFGV8g1KujIMOM7v8pX3
e21frNTUI810L8Zuo9CMwJgZWUsoFtutkFM2cM1jYfW6633dUOjMrPHL+tfrf8y0
uzI5JCwYgOjHoxItBuWPPsLdCiRKW+DS5pXclqnf8DPDMVDLyrzIpwub/5I4LmjM
wfhS+Vh0MVoU2UKcmD0Z9FqFL3WsOVWnlKVxWm+bRSPO01xnkwkO/JJ65L/SwXNq
x8TVK8Wx0p0vCFHldQOaVzpcnXMm5rqzO2Kx1oiBSpcgFH5Dzm4OY/RNnJNe/NBW
W0U7ulPC22QQ+1BCJxNGcYlLqoScSEQ21gK0GmbDPV6S5KMXkxVk41iF5nobWDgt
2IEus1mxjlIj4J4ggt5FX2A1SGIAub+V8pcDitm84WQ+PXxmrw49b0bzuHXBAJp/
iPy73ZQYLr4uEy6R0u0B75Cmls/mMfhzWM/gm8euBlvVncUxTqWzN6PjC4skwsEY
W0RtTZuUTY/aeGRG+/YJwGfPDmZ1FZpNbhvCv3YDfHviKhiTtplREVZif2RmoiSf
lA65OuCf+Yvh5rZaIujRNB9scPEoYqMM8ngdjxKu1Gqltm3McrgkJbxJQVen1TT5
rjXkqTsEk1BaOogA3RWDk5AXzAFJBrBviwF6HvOpRQaYFBtlncX4FE2CHjpTOB9v
Q8UVVoLO3wXrU5umFeJnQFdpDLtgU9YN4orCCiur1yPbDIdgYlN1r7J9G0XqK5pn
kZVS8PVk6X0RFay3uDXmiu468V1nhA1qtv9+YRFFUPjOev7RDJFPdDY6npItEVcC
zWFipn3eDMjuM5ORDjH7e0K4qpJMiMotenP9NyJtdtzDJd9o4jA9PgFdH5WVryeH
4ergoFPYP4q87j+Ps+ONoJ/NhlXN2k88mSewCqbnQftl7zsXU1M2buOrWEKQHVXZ
uqRsGk0PsfL/Kggw62X/fO/q9mYElef78BrIwBQmQEQ2BHU4/s2rYRyDipxkM1Z/
bt+b9v1y9AAYJ3oCP/EdqQIh4nRCmfEpRTo2/qjQdZZ5vshgrYB7TRQl0ezKG+eJ
qHJbhCJU/5xkpfUGMF8SOaAbglcCfzuUmqP8CJls24EjzE4X+V+4vZaaAEB2RwUa
7q44moQP2aQx8D4juTFs8Km3ebFF6WX6mT8Ge/ivdN7pcGas/DRIy9ArCrDf2Zeg
QuNKWTROEkV8a0w1asuyxmYoxIYPvOdYzZJUy6GjOgX74wvIqO0BQeZAdLsQX1bI
Z37cI8k0oAUa4vHWWjhkLsWruDSztKXQ4YMgDngKqtqXAeTK6J2DY0KCao7J1UrP
cHFAlsmENZt1ro8QYZd7wtmdC+q66ubNpAB8ckAJlvCz27AVwD/O+Szux/AGe426
1IRw+89mw+q9IKzOAQ3mFNMxqS32qr+tvMkmeAqaw/m7djRlGpvfgUrj6NqJ9hm3
JURKEhWd2rtOsa8uk7RTQm4lSgD/XvO+954bcX2wYjc3vsxRXLFj+X1H/EdMvBgU
2L39CQiHFPXEZ2Kyk/VdBMJbzaOivMqp6M5jhRcwSHM4VBySqchVqvLWJMrT6+ce
sTDej5VsWPlAgW3cROYDKhoWA7gE9wiu6DpPJVo5dMqvpGybSMw6xRb1apD6Ys3J
l2XtWR16IFyOr8jBrMthbxpnfY1s9EpMC5bdgG/g2E/5Fq+V0DJ2Fdc2eD1VMS1g
FUhml+g6DgRj+9gxJ/Akn5002hRe5oR9CK2LduPTYYE8ecj/2Hkchicte6LzrN6G
AdTjB+X5vMI8HaIh1/EcqQQGE7I0+JpJ7MweAXjvfVAJFI2j6w+L6B5LC28k79QR
57M2TzTf2XinJGCbxlOyyeZKFhJtw3jg1szOOWUqfeTyquE9WTnF49qeGZEkqV0v
WOdBYFMU5StX5+d7EA5EsjRbpJ4piQ3j8lesXNZGeewBn6iL1Un/q3ge7kQcmyNe
3kPaTMdKiI6h/XGXM1UEE95PAC7papWUKgJExbJjiDFCXB/5cvW6O6+2lH7jCppy
LBrUf/1bQhVDqAd4ZVDvg5yUFKyHdIHYco7NlFB+/cTAa5/kAYxT0GUYmS8GE+m9
A+h+/4nHumA4TndiKqhVFTPOaccejyodFMiMJkFeo8jJ0YdJr+0wC3ijyfpk7vQR
sZtVsvAc7MqDOyU5Yf1FpX7cNR7h8X+EeJsa0BRZ4gEXUSHR2WbeKb9bepT+LtzK
T0xzL97gvcDbrEFqoZpPSEHjaLRFLQuDPxjw/wvKkrEcP40hb5UUs6frMMtLB5KR
VFp2pyTamDigMFiB35WZ6cSAGMahzNpFU12Po4b9tEkqVDE3CLhJnhVb9vxd8sNr
+K98xs0zEhat2Z3yoCVPRNQXTpHWcebUaUEZ9usAIN6lRWt1PRVP7Q/fDAYTZPzj
p8/ZKtz6TcGdNTJnaKZ8rSdvTbUFb52w1EVaB9BUpqHBN4ex1SRf2OdJRIREYD/p
WqNUuKSH6rJ8Vf6CUJJf8CybfrXw86dzxk4Ck/HubFnfYjJyejIOThW0Dh9qe0Im
Qn28ZIo7gBM9UPhoVeQLR51HpIp3wbVKuLkNPRo1r2l5EiAovRCARROH+ZCp04hH
0B14k4g2qBu1mVFnU4VHh+IEjz5IdXbaNLofvhHUJVhqAAYtOxy0EZ4Dj7qv/dl9
RWyZrwS+zyTDf94AHoEdeA==
//pragma protect end_data_block
//pragma protect digest_block
4+J3jcl0ghpMyyArU1D/koBRtUk=
//pragma protect end_digest_block
//pragma protect end_protected
