// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VbJVCS9oiFcP2q8+i2LCzpgSo8h3EzA2D+nkjrvD9ca+0KyTKnegxMJ6fXBh
3p9BVpyARQh80fJlwDVYfkmtXdOjonCtqLnmgilGMUBK4GD6sFVHBuHLnBiq
DF54lRKeUdIwOJZnwCyfvi7mBul8tDWHa48IPQ3XBE74Z5rhdPW2WW9TGk/D
F+rAzEbCcmg9sxggF6GFhELVe3GNKqW6Jc76gdU2xuBp4fxUq96iPj4A+U8y
pmxsbF/Wnf8Eaq0+x8rN8QqslMBTHOAOTW2suv3tKQWPfBP3dOamBRgMemv7
RViE1KaANFM0kQPPF3hJZNbDwBrMPnoQ7yJyV9KKmw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Na7VsMhIS1gOD2VSLEmSNZwdnCRzyVmraGR+SamaUqdu468BGlm3qixVV7Vx
iP23sK+O1CrUaegVpFph2+PEfaUP1tPlgnmkgkLGRufPgXQC1sivV1WiJrO/
nTygahewu45ukZZp2lQE0Ji+A6MAMKTzgY4E1bbjfJfIieF70fsPUoEwVR87
sCnx/Gm/M54O3WCNvZaywQtWmHdANW1P0yKUVlNdl6vFOGE59P/gpnXlc+RQ
8bZmduv3YEgT2fWT2moAgFpOnJtaZt8HXCeACl3W1VlgCQWpcLfJjvzuRma/
ynhBvW/pELCkBzelxI2E4b/JpiRNeVSw3h/qgQRoSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D69ziMxyNTqlRrxNki8I3DksRgVu+sDlAIP3HNCGKlHX7S2iwBgetURJDpv0
i6gqSDkZdC1gOGEPkFH7JlM0FgubSAN92tSsYfLMg0TUrFJYI94FhKABJImo
9zaBvrTz2kLAnPM7ndYzB+D+uMUYESXcZLl31TQqji0J+9YPbuu2jYKjUmyT
BradVVVwkGNoxNYsHarGP42blDX7MeXUdcOEZNpato/dhtmwxIrXNmkDoWf5
E/7fikQmRTF6Qz7W819xVgKTDrK0/wtL5VHf8+nBYiyh1H+Yoy2mLRHyJA6N
pz37NTrPApsCtOU45+JxjuWwhn6FihPXV0rkVo+Qug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
f+KvSrw92DzgjRLb0uIaFAnEA2YrNMdQaO7AbEhCgJglv9pM7xBp6qh7SUMX
z7L/vXHg8HcgXNXquErEORlk5NjIzxBxL5nhgVg/E7mMSs24gz+bI8tZkzXX
nu+uSfDRFC5IDSoM4xE3ng5pHq+eDSkG95ACMnazhpazowxhDfc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HxfFeCOaOYrezDnbVw/85xKn3p3e+77u2ubYnc1MzDQXajb/Hqcas2dNIXts
d+mZfF1XtH+lmKHvjZQZi+HwEJWelcilzX9Xn2evRxRFd3PX+/H0KeScdWEY
Q3IZDaLMIY7MeJfsIiLXLwC6fuJF0nfU4r3boV0CuwONL0mM/xsnBDLzaG7+
93RbTujSSOEGXCLcL4wyu1lrlh58KVESzZYgtVOsyz5CBKFQAGv8Ke54Dk9I
Da0AN6Xx9EvyKF+KnSI3MR0MG20/aHmfnQTBwmYAU9gXnokB1Y/WW9yYu2Ul
tuCx6afM2KAF5C0vicOKxMiQrtMPQHddfgzdlNlxUY5qyD5uRMsROLyV8Ffh
sRsqGMAoRicJxOZbpVIohMHCAHqUM5IY4O2/PmppIVynrN/UBHYgtgdrdGta
4bRFyPzSQAxTQb7Hi+eR1rvycupqqwSehPbKZvNYojEgn6c/Z2d738s437jt
fHkjuS5fW2tsxn/wUlBrM2UVhKABcloX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SMWomeRyzAlA2g8fFmPnF9fGiXxbfEHoy1aGbJ1FdrSpSCdhyeC30t8LYUPe
OKS/NvlEpUkDwujuvDVaIqSHBHR6ndo7l9XEm9Df4bA7hj1/FBwZIJQ/sWTX
R3l8Xv+9KoXyu+1/Pf8KuK0PgiEopppFqCNBxxNOXyADv40ajFk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eoj3aEPKPbbRGKiwndHr6TI7JQgwwIdgCcBOgoPA25HNoBT4KKLdCYiJHiNx
VH3pqepX92/pxZc/Ea939Uq2x7fmRsFeKT47wb0goiZDjyfEZiBtOQS3yUO8
xEqYn302iDKLvUd62luEUNrwsDV06PT8iZIkVtJuDp91YDyJmDY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 77584)
`pragma protect data_block
Yuo8JYtoa39QmMwMo7yclsLalrr9PgPfYOo8vv1Gzo28aanRblgM+EvaaVV3
vdF4qLH7B79muJeltMg4TVeDKAukHMrJCiTFG/2OsvLlGkqV19iI++zVYOP0
BEIVd0KfsI/oCLOeo25u60w1MJ3X9Tm2TMSmRGXGTfNatPkvBgJ/H/EAmBEb
zzsDXVM6XU8Hpy6E8jEBocfFFnxJI3BvWr0ZxNcfey/1a2RRjPUdspesGbji
gelGNdPPD58w7HKCy6M+g4lLPNOe2TGaMsa3DqAxgk8SyWUBa5j7CpU/uPqR
9xcNesn1uSQ//b8fntt9+HMMU4sl16tpPUhuwKvxvsggw1lVXjG732NNShGz
Syv9ZZuo/JkXu6PeWANV1as0bBJzR4XwPR7C2cSF3citQhyhBHD2UIwolHqb
xVb8Sa+3wtDMmoktbfKv0LOx6grFwL4GJxLPz4xmBeNnl4NFuEb59DvV/sIS
mWNBsrUNddhxZzIkUIbtu7kwSVowMD64RX9qIGYCxBV7qjL6nY/kGQmLaaRz
rFyUtHhRktJYMnoJ04bo7o/Z79c5GEkXZ3M8us60PsOYXHGvaPXcE7KzvzMw
6Y9/3R2wxFCIxL/lOLYbL8MlDYtC0oV9BkOwpXsOPZMS7OQT100w86OxS9vO
xPZIo8hPzdJC74qIEpVqfdFRDUVf7gXeisRz+uDgc26BMHRY1LXd5Z8wtLtf
+ORG6eHIU+KuMRKd01/d6zTbYMIeK56Q3cuXOj0jDKR41CnsYxxQTCqXq+jL
yTuRnp9CurcEnwbM4wDknP1ObD0+7v1Mk9vHg8/dBuUkGg94uPnaLNaKv/HH
LkARVdEia941VoArtGfy9iWVjDnrCmHnZOZHYYgxICBVbWYf5U/03289Hax8
5br8bqZy7ojyfae4+FAdIKVIpoi40Re9mjz1pXnVdPcmqlFfnf4d5/2lDIwE
Vqa0WsiVLyYSCgmn6qi36W3qt7vaStAoBMJesT/HAmROatUeUKsAh3BuWZqi
eDkbo3pY844b6S6FVqEGbNvHChrh1HKj0mmfVokf7yHjmnUjLFmyBu0H8aaE
lDuDAuIc8MWZhHdam/4cGZtZHQ/36qtRbcERNz7QtgmTmCG3RcNZdfCTI7IL
rv+nuYZho8drq3daHryoA8M/T8f4perbPCcTmWTOX7zW8gb03SxGg5EAp4xs
T8pqjo+Jb7nQfrd/P3/5zTtuUYQytnQhSMJ/Z3aKxLJsxGrYokCULjIKWb5S
bOfXciCZJvnPDpTIHSEdd/z8OGtryA7QYfgsazLwFlhdn0QWVEirNmeVxoKD
89L5B8seQ5/FbRrDz3pJ1hiVLNn6XYNGmOvO8PEQ5SdkVF1bDv901H5+yQ0A
/oI+VCqvGzEV1sQz16hJ5YRRgY0bUN60gUeMDYqDkavT4wZtac3B+X3vX8Uy
IjeWFwOQNyYV3dfEV3JPgDbyRhlQDI1Ayc7ITMKWz6UC8RxlGEtz6wC1Xka/
oZ/ktCHAKcH/8OuQjIdf0Kbeyhw1N2agnclKn5FF6gTmthsWjzjKTmAfx6vr
CKUTEryxBpx+6kmMAtN2CYKNA5522IZp6ea46UZaWwD6yVwa2K1KmkZSaPje
UNHEJSSVWdej+K4q5y/cabG9zuXa4BOHUhqTJ/Y6AV26H98VgVP3AIIKoSDp
uYTlRx9LLt9tfYeW2lmPnIH92CHOeWwwnXKZWwaNu2A6gHxcrkJ7W8V5g+Cr
ENcyidimuWDfdg2SPgkfffbSmxz7d1lMAv9V1nO6W98+sfhjrU9XMhNHtdAI
Z+nA8yF5cdQWEOPkB08aGjoUxiYdmRsnQU8aKyHTKwmtIooF0akC68/re5mU
lWjfWX2W7TGCcP6H4fSXuU1oT5BsL/NuHGQJnAGtQsItaDQyTZWSN5l/OeFE
3bPq4aCqrE9pvy3opMyQt/KVlw9EVnMaZVjmLa08UaxPYjwNnMVVji6Q9gKL
T+uqVsnFaXqd/gCbtlZXURL8NbUpMlvUYqnyMNO0LnV5ed2yYKT/atwMLWrw
E4MkSvtgTaLbHj5SupOH3WL4tMAYsabvg240x7Ffr6xXPDcDQtTTAhZ710Zz
XC9O43lZdlEj6arIGnw9jB2INhBeW31mXfXuAmqVs0guMZYCP3tZ310hjQsn
Uz+TF8MOUo1J4IWuWeb1MuMRQPVx+PtNI1RQhWZSgvZ033g5+EXvDOKEO7Va
9A33EE9jcRgPtzHyPczcrJres2g+eDCe72Icds5s7x2efsVZ2gpHBPWprKyn
9j/2p77UXOVgYwf3HUeejpSn0iiO0ZZZCqkm9L+LxB7NyxmBbiTa3HtMEXiv
2YPw/8ou7s/epxml8/Op68Ng0Rms1rxzJGniBkOUmotypD99tXBIrKLEideG
h0BjETV9ZxBqNdVEc+xCJ9ToHm0wwuNj+1RZa6AKZx9pzjIduqANJ8BboT6N
pWLp+HJuBDm1k1qRQjItjNYlJCQliRorc1rgR5zcVdLLqcgwnLpTW/jJ39iA
JoXlg0qbgdiQ3rtIErsq4pk3vUMCl1QL6a9oEJp8MV/AzYAgL7ZSO4cwB1wf
c2BXptzCMvnUyhjpSgxUPL9i7hF3gLDsT7UdDG8zWXZTTSpNQF5I9JB+h/bs
TZTPKQIGDXsXxe/cV2b4tnkkZ0hNbAf5SkqJ9Qcwyfa68QugdnPTqocS4Hq6
l+vkLvdmeKG3LXWPZ1ysQS4cBoT6LHSCiyElRrjF2dvhFGhYGQS5kYt1drek
BpKl5Jqqkz5FeomaHPn5+ypuRpe5NnZtWhiRAZKmYYQ09/FIQwDnNhASRiWj
Jb4HWTAhIzGMYwAHuiG0P6MuUJhnbD4G6sZvIq9UnHS6FHH1at9+xxi7X4/x
sX8AOAxhWkzaYNQXStb96XGt61+Cqk7tc12w/GrNgzbz5kvz+RAJlCqu0Cql
euP8HuZsAvkdcix2snqWK0xSmA+EDx5m1+wsyWYtYXv4zsjRqVoz1p97E+iI
Rae6JjWyJjfcrfm3lP2U8T/+NpbovVEutUdn7A+2jgNiTjY72vnMdH19GgvQ
6p2dNGp68GflufHPO5W4XdpWpbd374VPYRsJT5cAQiZparuOr22bs6JNAjt0
0y69PUr6od1Fs1kT25PsP2hKhy5U/OFBZTf7DC2Dxv2JXggNMjf35eOzCngb
oyKPErbEbpPeixQIx+A73TEkGreHKS1KOxHYWOf+qSQ5G2zxdtMF0HSkRy7k
JKO2EDwj481isKQkmEIwEBN7MgWc7hNs1e9N8rZnwmEjwuOlIQajBlPw9Ws8
aI7AS71GMVsVtMnfh+l670ynSodEG4aiijpfGZJFNgUQFvAyZigmrWqwED/k
amPP7/6ks/P/51NyfGNBd49YPPmLZZ58kND10EdgXEtIv7C2JL+RE8mVNPIa
lLERfKoDqa05t3bfDXNMLTBfX7JzaYq7RSBwYff5S8AeEAmh+R74oIgQCdBN
TBnAidE8mHsWtFsrPafLL5Gdt/V7XliyYfPbAm0V03ZPRtLk4Itr5K3U3Ivp
j9ETEB2swHQstAprN6vvFYermKSt3HXYSLsRrycVCMaUEXEyMj+morTfRzJC
4jhZumk694LZiLwrdh7jk1c3vHQm7Gk/Vl45SXBh/US9RXf1ClayOa6sDv/v
oU7tFynDr2MQqadz0tHPEhpfLWZ8yJQcsr9svQux2LoOYflGp1QBInCYFvMI
0AVSCNElRYjsFdSsjboaa+On8Lnl1zaQi+HyVlcVB5LTejm1tJBPCp51yO8q
V1rQISPobRh4q4V8TLRT7YJigbo8OE055d3itMEx3qoZGIQ5+u7OMSUdS8jp
8oanohQXe2gzm+yaAiK+t6KXKFVQZ/JmJsucQb0EOx7W1Ex1iSxp7eziIivt
wEwb36exHUF8NxR72BYGZsfg6Yh+5xUS8KDKps5zGEO9geewJmOcc4juCWEc
VpWD3t6lbqII/QXs1TEt3lIgt+kGs75lXs06ee9uZ37FwbjWI4iEbisn45jh
F+wnGtwJT2Asb8LH8XU5o7n8C40mb4XVL7Fubf6dBUt0YEd2v7gqVZ6HFuJc
47twdXNVQ6GKlM5zgK5gsp4T9Ir4zpdpxxvdgfZxm055P9EIwBAw/FUVVsT+
7kloBnI2MDAUrXnhXeQik98fXNRNRKFCPjkV+w+iHjAdc6FN9BxwOuENAB7T
UpZXEqs2xPdc0e3RSgwjnf88Ak9ZN/QFDH7XvZmU+c5l/OuTgP7CwaPEKWic
L0RLC7DEr753OpRQYngtGgYilwzTmaf06ubV9GT3izQPMPfYvkayzqWX8N0q
Dp4s5AOwo+FjIhWYjikShrQUQVE5pKHlVm96+jw5ddTwi0oi1apeRTPD6UcU
rjlVOKMMMVYyj+sUrHGvUC7EhJM5nqXT3sBM8EYL1dWPhyCMp3EKXFbKvVQm
X3dy78xCkyGmnexXHBjHHOvRVAlBnHw/BmXbm7EbymmJf83Nrbn5Cie0cGhS
8KCpRlcTFRYvwhA6wvbyfNXfWu98SNoAUzJrOKbnT0ZVzD2ci5GROnw5ZJ0T
f5nNCBTE5gcW0lUADDLBzxa6H+f5WOXuGRkK0ctXmDcKlOOorkNvlHd30rlZ
XaT7BCQqS81tp7iFAWmwmWHl23nzZrGFzwPhRz3F0ubwG0SBuBSBUl5UZ+qO
c0GuY7T+V0zMRsp8NLAdt60S+wJ1V3FD6b0e2jHaGI7wHpxCYciqNKfbyYYf
/N+EqhvalIzprEqshZ9qm6dvEY+xZ2jUAZUr5+2zTeMjNiXeUYRmC/5+PTrf
r5pH0yoLra+dqWjR18S0B3DcK3gJWzKiI7y/YAOnwWHXfEEQu7O6dL2J8mtr
Cc0oaRKzm496No7KHmLoS5qd3f5ZUyqbATMWf3kAKVjEQEGqqZd4MdRGNOAJ
1YjGPAyIQoEJJ/NQE6SL594WIdNTK6WL4GejJmRaJaDsaQfqjeLQ/pTKNZPs
/jU/ByiIWiVQG6xr5Ex4WzulduCwqgk6yyeAEAhqFPe5z/JBTcL//qwiD5X4
sCnGhy8leSbhE2KvMD27CRp3Mh08SG8n5FvuUioMXxOgCMVxO28P+wYNeM0H
Z6DMNNr8pAPPT1orXMpA7k1HPzsvdSiqJS6pbIKGToaKNz9WJ7J3Gm7uEQuT
SIkpZszaJEFiqVgiWpkSJ/fw2gWDWyFKxcl8RgCVHUQbfReSj997PUgNvT1y
IJnDR9It8pACmvYT3eZni/UUHkbCyKiHy0nbPTSalAhSeEjAeWHOLxqyEOg8
g+mkKteCvYZKV3clYnb0b5oOYXS/pCcit8g/BsFH0eUGZmxQKos/ZGtEARM8
i6AEaSYNffR4j+uVgL/1XeRzr4iRBFsSLk3bk2jpdB7paKMuHHSbQofaIHLT
Ya8XeoL5ayXNdP0nlBhEaY3oL7sLKT2xf3CAZF+UAnUIibZz4tJhi6IBYVvH
62JLokK2qVHZRG4c9ubkxbhfT7kPW1q5lq1SLdCfnTaOt1M+K5yI6prrT58s
K91M9Dr/E69bRx35nkxQGGEU2z1LCLVnSqF1mvRrLIjgNLa4ENMq0DBmAJkW
bX54gGOvFH+kILZ72i5++kCC1+4irS895i55ZPDIT75Xz8/0gbnmyt2GhCl8
tsRS89bTZkVdLra7gb3jqFC/pb4OlQbDwx5PR4dQy0EdH5hgvWgXyaJ9zEJs
YObyFJzUQk5sz+cRaUFCdjOuQ8GJZNn+5jLEFEvTlongKMq7C8+UE49yvGn6
AMF8CMP/Ka1BmxcIFjVdso8ynwqWj1cz2jnb+5fBNSXX9k8vuoifEbF7KRpy
DPomLatqQ+nm5+8Dqul6fWKZHD/FqeZDJN8kUyu2pLW/nzn17+MyxG/Qj+7W
p+zEa5J4JDJ/NSmhq+qMP7uOsr3Vrs+mY1ajd+kbzoH0GX0aN9u6ccoK6OZy
Sb6BgYXbyq6MxFdUiBUkPC5xV68xrgc1kabKj6B7GENs/OHAzwxlFNzh5Caw
xPzrKSRMygYM2HzEkKzj/B49AT4ftQY2szs23fx6xjzAE3ae1g8LyFbuWF3o
F4A1ygTN8gO8RPBsS3P/SF42swSa5er+Ys46FZxDmwzy9HRLKFeW1fD/UMmj
2O0mf4LR4/Boe5nUWoqYS3e+EeephAP8JvjFg/lLUsBzu+Hgsh0QIgpSAb8u
Ztq1zFHXFFtIJpzzm7581r5iQogUMMvZkEvFLuWlFCQ+yRzvZ6dwZRDSqB5Z
R2OAI88wR7Jgnwi5tsjAqV1DHYp9dd7KmISB3NQ8rd8JN0hjT7wniIGXokks
FzxKKgayQ/VYZvGpLKzMj7gRY0vQPd+HxDHirzrJpusgTcf1t40wNQVFhX92
cIgm5XW4zij0sZ1WC/3WFwsC3JACcBBN3DTJ6LBn3lmHFM+Euz2E0+71A51A
fiQtObk+uTWqqZDKLzB7HspbqWUU53R/glZFrHUhSWgw0xGpVzt4IFQ1j48n
SmIgJ8cCNxJiWhKdN9ui7o0H1FD4C8BxY8vslAXbhmNDBNRBXTYp+rUAk2jj
oWCNxuSbRTIaIX6nrZXopxix/k9nhemCSP7gy/JyVjqDWM9sTy3HnmO00lR9
ekuiii1Y9FDXMUkhQLU/PyGecwkxJLZnDhGfItE55Aa7VUFvwq2zQJZad9IF
Mtp8IpqTa1u1mR+9Ern/lHvNf96Ovtjkd1uPro2l2tUaBWS1NPAzUE8XED8x
8UQX1KpBDehUO4IfBrT24iZoTblsV0YLkaLBb/o/tnVaE1XcbFHeM1+SBrvu
e3DsqRhS95xzRrh719/fxivYZ0OQxRGJQkVie7et63uyCFBgKkbJDTE658GR
RXGlz/V8L++wtnpRulUjCaBKoIJAQCWoNKKw6x88Lg9nvJYW3H0Umo9u527M
IYiupDR5fru0sRUdUJZP1IGhPx4LPTb8f48sN5lnh0KQzIxYu1cr+C1joCQH
Y4wbH6rENjpvAAGt3N276dE4nxGlAYr9RFYVOlds5mmS2JDREoyN2mPNAIcP
H5XZNYeSggD+wrzUCb6owk2DkhIWs6ghZz5r/TKS6LVuFLs50/6CP1wOX41Z
QmC0wOkudIY/HRAvcMqEjFM0D7p7KuzN7MTEo4rATDqbRDGKfr99T5OAACV0
zPsHFsJ1xAGaCNTJOnEFEgyzp7M71pTQFuroWsrR9gGOfMTW6hVAe4IGEAwk
RpD6Iz5sfdyg9vcx1eCq8n5UGmqxGsyipg1Ce3EFUaAzaDcUqMy8DfLg1Umf
JYNMIEqNPuLfYT1YNAurcos2kAGU6PM++j6X7R5DQJnGfzhO3T6dB+pZP47m
1qBf3fmA6EjOKPgoScLO6yQ5iqg0+2RJbl6/pB5JuERLPI1TE/KTSwi07MTn
0m+KYuRfBQqOIDfpM5zGl74YGYJGd9bcAY1BBKRWeE4tRPW/LswP1woni1Rt
cJySHlqq9jLuHKXyq6iitSu7hKkjgPCmBU7m6lwM10PYPLrh/HUUCuAMMLuX
33umPOmWpd7vU4X16PbfeIgate27rMAVRToS+D7kGUqW4c8yJdb6AY665KyS
XcKcVDWD6JqO5EZV08aqCjoJl4mnUcOI459nb2a6POsS0pNILn3bV17+8RTM
Xd9tYm3PimW4slmCIBX35WWQ5/p2xujLgP8gxyzF07CxLG2WXs0yeeRJOxui
3vyB9FKwiOZLPB40vK6uhipsqwEZCUV4nkimjO3vr67wG6HfFtpLm9RhJFTV
rnPzazmZU0n0QIA53s23IsJ8wPfcVp2uX3eJjHdaPlOT3EzFwwaOuTpYu1y2
LkVOPF3D3d8YqHFbgpwBmEPlF1AuF0ZuCv04ZJhcXAADRpOKnLUp1h03tCH4
7QAsvesuhQXxN4YjUCvSkq6gYtS+piDyrNFHkQQEoKED+mQQT01XamIBFedY
b05QAqYS0h2VUOmd0XaOIyGSQy1ZHUfZPJ44CxsrGQ0GMmUquLTwaCawaXyr
W1lve967R8cMWYm1U/THu7E/glMFJzIt/m/176BDPlaaYuzZrsk9eu8Magat
rg1ixu2tbET0+ozGIHEFd+bODn45StZacnm3Rw+UdA0KW8wt7AlCJ1UT8/eu
Fkl2IBmmPE8fAgBf2EXsYHx1gmjiueEaBDkq9ldg41+qy1byOZiw/kLmi+NA
DfHqqFKtYXmJlR/GYpi8omhwr0jMbzBIBjMZ4yG7XXfxRh86XQBowJTKM6iU
pQVqtjzY4Au6OnvcZw+9O4sFPQ+EA0W8hIZvNpIl6sr8xM8zbWEi5ocyr9x0
3kh+NjhAmzIm9ufdHjKk9EvmeCWd19eOZL29USDffx0HoZTe6FS1YAhISwGH
nerLXevwKOQAR54cl4NdPK6vu1CTQEmlkY/na4ZMtoveN85lifEB2ggNOGlG
3peCoOBaQg6XdoP/Xrg23sj4Pq0WAQJSC2b80CRMCkmxeT5kLgOfV1+HzOsj
ZEui/ffY8GQAsw6BFKL+40NN/6GclIuNcfHNJ29YfeErI18j35SwD/zd43fo
E6ZR7BsKhn1S4ewgEYoQuPABKMqnQi1PiATOfb96e5bEtgWHwjkI7PM8JNFx
G6r+1g0IOtBl/jK6hY9D2ItahJubU5Tk6RJeq0AUyD85zP345XVZvn6fvHVW
ZKe1aRe9JCTZEpB/sfCwWvFYDPpgrp1Auoxsk3Xv6s5FrUJjB5+JiPiouqqC
TnnBM+9pSH30diKX6hKTtDxIw7Kf2Gby+wCFXItt9iEj2qPSjFxNNXT5FpQ1
MENcUrIjmNB22bEGm1r3PHY07hgZS6scThRsCBhd4VNjyQ4aMuAx/T9X/IiT
GvCX1bjUYF0Qjrs25OHUa6mHSfrMLzWy4x1pApoCnpzdUKXsjp7Et1ILcPJC
cibxSq1oo1RJ7sO98mrPmk5Ldzda7/m2+ywDZcwToRF3BCrkce2oKXqcRzDo
JLWG5UQONBpy9IDu48p7fKIaiFYfraMqfH8EfLjaJxOjvNv+3FOR99ScrzhQ
9ZbMZUT8fTc2HCh8o38EW2HrOR9/lqs5r4gx9yfctB5tFHq8e/TCbWOwo0mV
H/v3aCufvVpwSzS3Haae1qP8oSh4ZOo/Q8RwVhoW8jcSIJ6DIPsf+XVarfHX
cPCqptQOONdn3HGyPOmKl09sFKPhA0c0zBMeh/LThz0V4wLdfwOspwYbwMPq
s78HfAyzDOJOl6v8UPNe/QCEQ96fGmE4OrWxO70GPj/TN0AYtphX2l/fx+ce
i/GovEGvAE8pqWNl1JKrxwajgzHJ/5pfnj/oZSZtsfQfg733oxw5Q3+oxWOM
o858IHwRrBdZeI5yVJY4Nt+Q4/dTKhjvNiKXYHXk/xPX0LK53sOlSDBZHlK1
Q3fa2ByKDCLrM5016ltxn9pkrCXn7zwXJGZPLm/Yt8JTQkZPfZNdTH1Gin1i
fdCI1OjYjPeEWmbUjPt33Q3ciGrPb0s+UlX/eu57F/EwaEjttVE1fVs6qflO
+2beqJgd0tRRAK5SNTHky8yzBKn191yCNwDp9k6RXOhh/fJY7jQAfj/PibMp
b7S97/geJ4Gh9zeqe/LsuhYypyhnE90siruQH5Pqf+E1JSDXSIxQMJtLVqrT
FQUYl4+/rbzgWsjk2EldrafSUVBDOA/8gflJUGTJUIZa5trjVk5YGhPWUQnj
15yRwFMQLB2rtw73ZQdMD+WS0SqRWuAiht1XcYmx4lOJyArruVtMgVbihCfi
IBIxmNAtNowII1tLMvCX0IGbpyPUY7lJcrowicQmLDdY9NF5zBKfc9YwpOL7
MXS5jL6BAndcWq9AGbMyy4UJ4T0TlTmGC/T5O46MjucjQMiKOMEpY3awHTvC
1n24C4Am9BzuohuVBPswreqyey2ImW7NrSQ9lN1aUaFSr7PxPN8SiA/tjbgF
vAdHB+jU3a1EZuit901FiAJT/B0/NzaNYkKVF06sH96kgcjDLOpN9HiKvQLO
o4ho/vDVQ3l/fK5yjuPJgHxCRJb1hy5AzzLoCbU00hHNQT/0bkdReGfpGiGt
HgUOZq62crrH2Mj79Y4hbYeSJtgZ49ECmurK5Tubu2zgqKEkiMcr4nd8IC2R
boaZLA8rGPCO1G68iBAQWF61ixusxrUroSziP5RzqxSsAMweohSka/IXbCiB
aidyUJTDM18dxsyI883ga20qnFXbYnWF8N5e1d9pk/aFFVYwSukIcV+soluf
vv+IY9PVI2FdAR+JlauOuLZ5Qth6x/J/NKIzKxtXgwxHdZuLI/VQY32jN+rC
nron7jOc8VlaNR1qy6hDCGz7W+CKyYeKHG8FSNgTykGJTLUt/iReMyrr+oyx
5XUPbsEz7QK89jSwV4aLGOeei0W7y9pUyhS2EYXOWZxeiHWfxkvJHosWXsXY
jqXrA/bZdsMPDp3vRi4OgfOxV/kgU6yMexfcllVa/oRuYNAom/7tpJLncQ99
65vYlBfRBaPeuueTexKY8oW43hq/mT0PKZWIcWIzaNYYWDk1tqDDfzuClXsF
xPTVa/B4PmgReU3QdouJ9UCwbA5yY7VTSA+zRxKXY8s1QH3jjzOVkh4DMTvg
YbebUrg4Ycd1MRiWIn1WjwR+HFeikUWs7jKkw+ZZ03uCRKvZw7kkNACcvivZ
1WJ42lFZXFwn/OYiKOkdCQVQV+oXSIybZJehyhyVq3GAJp1UlZNBNLgkexQp
EhwVVsO+/8ejiCDTpRS3ljor4g0gjGYEq4L1B2IcCikhgJWHTOYz2tS/WRHi
cUIEoZaFX9FTRplKO+Gy/jWNuf42NyMn+32v7BRHoZJyq3uxtHa7c/LAemJC
8wr+e/WKyUgT4drMOcOf/zbChwEmvVfXSRPJCG6WRoqBu0Tw3ydhMb5WruMO
w/boYm0EGAyvv+iK6Ch65jpqrLwVYLNC/0sh6YNkHB8I1jPkr0P4CSf6p1WA
dI/YwFGKtBJFKWwTzIMnlATyR26tH2jBG8aFgrMPcYhTyZL8Hg2t5xKYcF0k
3oOK80PLHJ9tg2GwwkyPqgFUREibx88De4UwB/rFgolFZxO/i4/ess/AjDxa
CtfAhjjc3jQJi6bwT8EVQLGzYfX6MvlWoRRPJNUcQBZOZHnzx/tC7n/BiZfT
jZ6PLiVycJLmSdj4BqN3QQK7m/otdjEoxL6a53/zDmxP9c6We81KKMBPwyjs
yHXW3k9ksBWoaayJ6gC6sh9kKhV1Fv8q42prmyTeif4k3dZa0//DBYscHrSL
EH5Xq24WX8U077leqIHKZfaILcarGUjKy7aNFVzzc7RLSfuOTSYao/vEzItE
i+N8sBiTu1z00NhYwGHHtXBq8hmdxchm0xmoJ8WEQX2kV3/WumkyyspPcy0t
fvA8rsv66G9S7nhojNsE2bFZTe6VgLdFkhtGdqgf7MV48cn5gY6pOYJahtfP
vWOZH+grxpEfo2Y5YLsg5giuNvI0Ed4F0dpYLaALfVUMwkok6hVeHz4xelHd
PDGTJK2j5oZnBy9yZ7NNkJ2njFp7F0s1EW5TS8bVnNrBW6al3lz2BuahEqK9
LzNOU5lQGsY76M1QV+UCmVuDHRYr5BCXYPmvsjblpjK1dcLSns+jMLGrEZvw
kxMMe/WGoKXCZjJBu0Bo+JpbIOiGQ4v3Cb74JWhF3C+7HuseYJ0AyQxSRqTt
wrdjSZ5rrLX4bpG+2hHx6sU0ONQk5WsQTqISsYIB8UbJo8TPXStLspZwd8E7
b8UkGRw1RufHI0hnaw+TQDszLH24nzrpiI+PKXAE18Cv634uVtbHz2IDDzBx
meiMzWTcOnvqNnrbxnm/fA7wPqJWHjzCDB0FUkU6XEjN1WXPZMwdTV2rzfnm
MlVXFjXYvIEJHvdjeI+eWJ/PjqlDtjuaDr6cPC5HpI+Y/TuNrU/Pmqi86z0F
qS7rRd24tbrC2TRIzmTTtZaSlXcWBb4QKJdRD7bF/Sy3NU/MQAW8iZcm5M6C
FTh0MrGqJL2Yb50PBT5OdQEgPioAITF+rYqecUpBWKIEkQtAAc9A56wU/9L0
9ztLrloEWgl0C3c/IE+64yyN1atsrWta+qEO4uXCyhzV61RbE8rrrYIVrLs/
X9+rL/TBNRC5L6iSGrm6KKYSmMDyiP+O5cgf8KsfroMDEhPhA/w7AKBgPHqc
nTqQrlIoXlW/OQfEjtxuyhTR+wn0E4sBSzsJoS7QJANHxBwgtkb4R5GSC9Po
kwKNucFWs1yIjqcFVfm7BGjdmfDxwFiWfxYzcp3Fzggjltmdjc1BThPEnPq8
3f4Lb6CtTfSZ1O9QRqARrj3JSMO6ExztUhBS4jGinvLggEOXIFtJp1o1egZY
TSF5AlnSIJVWiqXHNfnRSb2zSzs0o15Qq6yRdoS0x13bQiPgYrbaVKvsaeBY
5iLHI07NKAD/BpxV3p4G9S+t5FWdRqRxMRmDQM9UyIw1/T8rW8LjUDqUpukd
nMBx1hHlfmBwppAp7gLxpz5jg+5VGJj83PQ4u0E+aN0NOL14w56BZ7lh53yL
c6iZ8WPSXK+ozdCxxsWGPoAyYEZpIfwWpgTA4bkR/aEtDZWm6waT2a4j6hrr
egk9LKyq51Pom340RgRDLvNUi87ahRHDMb+XRZE23EU78yTRv6no5sogpk10
90Nof1VvhOD+QVgJLkW9iwlwc7WNF9hONLPounwbeuxoGyIcflJNbwPcpfPZ
f7tTcaQrt60EkPPF0Hd2OZTk4shDcBhQuUjeS6tZXUzGhlo+qLLzdJ0nNuXQ
+QfmBtT6nPu4kA1u62UNzPWHotsqbXXd5jfHrd2U2mQtmgyDiEw6vdho10h+
a6cTly/zlTV9Q4NL+t2ICkT9uDJkwXdxwL5PsKRdvvxezu3Ub4QLSsyzPZWs
XRsVVzeDkqDt9u1lhfUqR5gOjS7Qsdj/D3fH/XD0aZhaYEMqnMv6Gz+EbzJ+
taSeel7pBrEEdVDwLRw+KBaVBUoqs9fgkZt+aZqp4xmrhQbfiYO1C9mLevko
nnm3JsavcvFpeHHMB6Ug0e6dY6mKCTh+kPUY5IzrAZLpuDs+r4uvLN3sUkl6
eAINAbM9uRV9DIXelDo57lpTL5+IQIirRA11DCfANk+H+003HynuelfyOEq1
ZCGZlVuszFc2JwfhwcU1LOhoBDO4NBNftpBZU2VqoU1fIw3q4PHyNv+gdN+v
IoySuIY/k41I+yfNM9/JoW90bQMm0Cn6OTqurK4xcyjtkJbl3Mq40b4ABfvs
V6l2vX4cKcm5mHRLGJHpe2Xc/o+8vEBEXSuNIeEUn3J8zBpnRap1tUzzZrA7
XvBHVmMWoRnaTcDbEzKrrH8aoiKYK4zzkokKObemIJaM1Ryg8wk3UyJzNyNz
tR05099QOqG+/YE6zELs7IimtoAn8Fem1bAQl+2NKcnvZzntVVlQgLb24Zg6
yFLx8vnFUe4yTonrTZXHYthCyy5kcVQqDoSq7lj0WBfcoHw2kLYr6W6H6mkP
wFzrmB5n/mmGjf4rk+EIlGVzO92AL+EYRyvd1QyCctdTBwCYWEvmU9qImD2N
MJWsh9n1x1KOgn0349fiCqFUxSuxtHAfhV8aOdvZnJBEQjkSzl7y9t0qGhiC
bKdWKVEhyRcEC1TgKSV85OPdwwPaebywX5wkqFZ20eWNNE0V1or5Y5LQlKzF
/DQ5TWj09y/b7h3xwvxIWtSmiy4KijcK5ArgsTW14x6SvLKdUtEKRnTwea04
ncOhmxUi3aXvUaJ4iQz3OSMrg7F5gnnKbLrLcbc0mDbTLDxg7bwQJQlT12H5
8wxwfY63VgG5FptxHDmd4XyiUP1Bb28dH4ltINapWxuJPQgjgMROe3JV1/ho
OZGHpcG2ACCO9cYyfuH5pxAFr2d9dvZKt9rsxApPL+0eRvzIhzSqM5t7wkjx
LVlPun8rJbww6tPbyc8BvHFKddHPOsspiOqsO2/GiYOkP63kzMw3tbsLTMpJ
wxwL8ZzXIN7STB/TYuDsjWHv6bLEBCVnFe8LaS6rJKwQGVJwNYxCQAdQKc3S
ETtGWkLxGFiUHOxs0hUr4PXhP27CIz4wvyncws/1daNopGzZ4u3Wo14638oA
UB7Obok4UjciV8YuZe+EypIgyd4eueyi9OIPuM29mhfNhjwLFRZhuboGEh3V
cIuQ7iamzat2BPq+7FjtNIh2uzKKr/XiBnqVFk9BXhGWCLjuetqbeL/EZuII
l1di8iDB9qnrcIPloGWezk6AmW3nu9EKhLTOfC4ftCSfEbX6zaPFnEgqL5jw
CVSOYlfxoLitEp9cuLqc5pz/0t0SQnJ8lqPN/IKulsz+MwMqMLMvBEwLMXp4
JmwLuJBFH+jV06FKfmFzlSFUA15e0eFCUb6gPIp98BemzSGJAhCrA7aFWtj+
1HAm4EarcvYvJOjh4VZKxth4l073U3+qT5hI0RVoC8O+LG8eF1j7uFuaikbG
T1vQanE0bLqYPgr3lYZEEjw5IZuU/wErtVWlM2j1aCPJUY0wP6U9xHsBMH02
tu34kdkjzTzEf30BMhHCEz21fJMpjQ1kCv2xHWqqiqm70c+GsTEe02JKsI2a
i5OVg7SbDdpLmX72HMkaNQiQo+417FAkg/QU1YTK8jxOozQUX+LAExYTaknK
QxtoaemMhGm7RkYr/lCBZ77YskPtOzBkxUiqdKiSC2rneS36mqx1/oaJTiGU
m9lkIG31W85NH+z7T5oAAyqScw3C7cgEAYMwwjXo4mOx2qwxN5ZymBpHQz3U
8fLK6fup0N91cjBsUGw2DGDEN/iKnpJtmNv42TO/VsMK1hqtfaCu7nlg5bYP
XLaCg+S97fsIFuxrC1ArY4FmjNE4yVsgbYohyF3B7X8rgXALSwfwG5ZJXio+
wa7WKR6pgK2wo43XXGQSH4OPiSiuZRcoDqLUQiMg2s9HwdoSZKA4EYU8RSbn
mjZw5W93j+9UtyApeHIxrLjhGol8ZieB39mv+JUvMLdqOQq4kTUCbCnX9as+
Mezka9AyOXCo3xwRGlY5oBsSj2tbVm/t3swc1F4YNLz4IHmkxv6kmyGsBQ5G
M01qdmTLLCYU2FnL+A0F8DP0hd+3LoVmFbwUiBG8nW/bloIeGIY9biEW1g9Q
11RdwhcsWoOj0ReFV0xp2v6Uju3vcBXDBrRq4AHhpHKDq0lYMZLBji67Jcg/
Z223dVZ+x110/LGd7wdJddfs7gB67jephRsTWCeZjEMunOoVcHWj883npYL7
QCLUUPFwRczA/yiM8GQl/7greet+EeeJEWjvFDm+FANWKhDNhmWpnoob5IQx
mmD4Tjp5uXD4yen3fX7p/ICUTf/TbTwjvz61kEN13v1ePGd/Mi6rMqsr8TVG
S9lUduKe3p7vq1IICkbRnhEnOCMk1ALTxNTSV+jb0paLHOUud1g6OdBTwDTW
0KTKjXyn8oD26CjLgpSvrdGiXDd3v86y/BO9wl/fa2hGdCKDv3QrP1WHxDT2
dIfrD2RYSDx6D1/tJiIN+4PGz+ECnPig0mUndhjJVVKvaZ7lynzJ+c86m3Or
rUZ0cUUX3SMzO20n1IXmQ8SLz2ClaXyoh/zk0swxwxwy0WtimQjjNh2AdzJG
L0CB/8w+QdIg8OmdATr+91GunlIdr0M2fJu0ErAxbn69kRxtWBCcUeJuRBj0
zYFzj+oWtkjQb7J3+YrPvOTu81b+XphQDLli8P4Y/aWpbQk6wOkFcLbEs5Y3
htE3926Jlx6IqBehMUqKr2uExQYAUfqyUion39RGc7j1VfSHoxGw0ObuMRj1
fvQAeJn2bCQ0ttQGiabeam6meZ9XGfnL/OwHFjgb7yTaTJ2pe9GbUsu4Iz/r
ZveidJToOanCJfo+ajING0q+QuiwXWVXa3N60ihS2qznbV9aJ5myACnmYQRf
giUIj58H9Lph+9BUT+lgNgA/4aO6a538f/Ky3xv1UpD/qUs3t00Rl9fY6K7S
6M0QKHNpAY/ja5QJknfXGDJ6j3cwKiK7YKo3ypOwo0mHFW25W4inV29cdOWZ
LXtLTaDp/saAtlcLP4BKR5r4dy0jUsxTAbYe+Y/98AqPzkc7XvzCeFVYNo3h
/D0WCPzYSrCm6eWforqQYmmjhRmu2W2ij5sxDr3ZyQIqAn2wQ915uhxWckc/
2YS9kZXEUsogQwrKdBNYVIUOVDgstrH6+zY8oGNJDlckEKBiS87kzVPvM/ei
T9eDXPZXEGg0yoA0bF0J9sn958He1VzoQ9FgWspJM4E6vfnFKbus/PlblcGi
d3R7tFG6Jke7sfJPsWYifYhCf61FXcyH/+wldC6fmx1qkIqui3SNBkqdKKfu
U6rC2SCifsS2e/r7Fi3qmX+evE/a8E+xGzC9VgIj8AbdawwWFKBuBsr0kdi+
sOPmv+QDbHDF5DQF4+IB9aICPhfyRqLb7oTh6tiE3LoambPjv3uBANFs0KxR
PywEPDyIMAI+2n9RS4Ms0AOV4+bKKeMnx+Yy/80EmLfytsyiwASaSZhyvsu6
3dwqM2dgeiNOhZ+K4slr+rYI60iI6zhKLlvGLq1hvOfCAuhGawK58k0avdm5
IdIju+370kM1hllWf1j3636jBvOegmu5I3mtQ52FjkaOr4KMxrrd0DhfDCy1
A7W5jNUnMvVjeamf5dBgIwWUWMoXhesonAbL79wwMzMyg7tMqailOHFjGm9D
pxG/3zkh0aqWhR0+oW77q8fNiyHvm89mHP2sIsv7xJJhPuQaeh+2p7f43Ayd
SC/iBJyuZqMvAojLgfqv1IivrtPbcnAaV86Y7Lw61earWcsLnIX6zZgP8flb
bw4jLJ2obQSD2X42YmY+psnpQNsUmek+nV8F/fm2rih5yD2kLOdNKvpQytuA
kJ10s2Urr+v9z7UjESBHgo073LMGWqTNaG4J6YB9nsuluZqHbGb7UW31/Ae/
Es04a3nvwY11RmTdFsil9nLVhklTVlYr47mL7GrfHJcgZ48+gmx4EdZnqCGa
sgb93EjX8O5xuSxaJlSIQLSIOiL9wNYaw1Hl3W0Q1855dMgkGXJI8JhhA+Tk
7qkwRGdigF2cm8OwQDcSG34i8chvAOaHJe69ZqQGXsapWP+dQcqLZRVro0do
UQ+7YTlCEf/PNosls3/moReACNyFR5cCMPI+8KgQIVTUys873+AtPGyspXt8
9wwR2DW3IUeW/Z3vMyBbHDtzrz0yZrYqy+wcaeZF2U5edr7ohEplfZrlkDmu
Fa8Cq+fMDUwYvuYSAaCWmjkzfwoGGpqPemjmqX806sinxFu0+Au4sBLuxMx7
YwLuEKAx23dfcodsQ2VVNsCRVJfRi29vzsD/h2hImfFCYH/VmxNDITgdiyJY
EJ/1qGp0/7J7QhgABuHSU2taa4CdJkpZuV3faxMayaufyfVGghTs4mfz9NvX
2CnXl7yW4cE8GqCFs+qcxDPZ6kur9IACpotu4bvjjAMpaZp9TE6vF8ImFKhi
IWlMbXBviRJX3fEE0ud/dr/QTw5Cz9GtSieyE1A4p+fIBOSgsguafk1w3+/E
GQNvMN0MT1wnuUuwG3WldHVanMNl6JHcZGYjtkMo+QoD4ZNtfrEjnvEp+fsF
afiE9Q0JVfbCfBqJSlfcIZQo6RjVVU/nF6ADdJhzd0u7CaHCB6rH5+Fpjk0e
FvuE4ouLyOnT1/Gv0RxEj6ZQtbqfmJiadeT2zcFJwVrojLbbXe4auY3nNQa1
wDtOggmXA87VN+NpRgRuVcSmfAGEMXvkqQT+rapsDWO7VmAWL21GMBohy8eu
lV+ltP9WuFXC05MHGY7OOufqi6f+Ari+pvM0tjxQ45pNMKBNdcKrwrxCHM9R
X/HG6Q1xZ17RbvGFZX3Ws2l0T1q22sHcYJTzjz3CMAaig7+tnPZSgoHXlYcI
PfLr1rD2kMwGIrNxsA78x2sCyJIGI8qMJKqBUR25tpqA0OyEZfLNzF6rChQW
gQVqmYrmr8i8gn4Pd9KgNpZi+JKWQjS1b99plfNpzCw/NQyBolXYjmu48oeU
x5asbfrNWNdQnTzL623Pnaij6NeUnlZBfPRhawT4ndBSe+NTy95yw8P0aD3J
vGcLNvtwNP9+e0A4N7+eXCuuxgAeLt4NNoJAV//RTT6XQTJq9pVH56SY/zIK
HfTNpyx/Wajti5qy2S7cnQVKFtvPnVLoc76u+LCkWLzOB0VhsSW5pUZiQ2kc
GYVzD6gBWixsuX9rlARW/3hquVCJCVWxC1h+ZFJGjTFJclQZh5ds89ytEfZl
rTQR6sa6J8UQTusnyCA0GzKkXzszVeO7skeqjZggFqeUg4XGVEJ8Zmn1aKa+
y9F1TQwAALaxsNGkmQrqdfUNF8rUdmxf5tpV1mj7xn4M1SGHX80cEG8CTzZX
8oZszA3+sUtZ2DkqhAc9Kvg/RhMZ0Tc977mOeXsCeMHmZ8Gtra9HbpRJmLBq
u0ztLclqJpPVtWGI43mXl1V7X/HmtPu6km9mFCCvc4J4h5XT9gT07W0xOaVl
izGVs1kQt1kwik0hTH9V7pit4s2OdbB1wo66PM+M3UryQFKs6H6dVQVV83CQ
Zi88cWbdcgEprLqLhtGfwM0hx4a6AP/DTDblfIyBIn2uKWyIJ2ps1OpHDq25
vALWOR4znvR6XZ96m8RSj0lOd0JB3YXqCPZXpoPll+RGfoL08Meu5ogL4pKX
57YWVvOtK8ssNaXV0XFz3tv4ykl1JrU+hg4jCy1I61kjTwrubcM+gQXtS63u
JNAKS+EEvLKqaTL5c4tfHCrvUxeybwAcWVE3ptW2d/G9UVW5W60T84cayVrO
j8huYSttnhRuXchuwCSfYFPsR3IrZTOm6GWNyO4KlCEseDTOYpB4nlGRWcox
fELwm1A0kD2bJBBO80pXUVrEPxE1d7YJCw0L4yoVJnKufGp75tr+QO+HsI7X
75LDSXOqG4N49dAFoedYIuDBujeRnA2zdJj/g9PCcq236TEthwKagEq+fp4u
4Fb9OFgjsEzgInLCi6j44UNwaPNXkX76CE2kZ3+XzaAZtaGiFUQWSNgqgwrl
9V3x+BOi0x7cXfYzwuBCHjDQSejAjxLtrUOQnSnarAT7CmcQo9Le4a/lmxwM
gUV03gJpfZkyajsd3nvy65HGCuZgIyUPyCTbDeKPrRj6gvjAvpwS7t+8fONP
x2QLdQ0wFguVokWom7YE7DFeoLe9PZgYD27XTRh/ZhqHvpSLd79Z5mbJdC4P
zyVbXxGhpLOyp8XCK1TQYsLPDpk8ZdZiL29CfFrZu98ch8Fhe+eGYSXgjuok
7PSSTty7LCRkZGK4Q9Wzz5d9Om2JsTqNzekWu5wustUexeI93yO8XHV+KzhS
F8E0pvTJdEgdkWE5U1i6dtzXqW3hZ+XEYygrgJmD+bpVX4UwVDJQw4VcGMaI
ZuowR1q0SM4CqAIETis6DGvdn2gQilfXGU4uu1EValbtN03UWPIKhID3llnL
tsBH5flA3K14ZCFPrbsHZKrObdZo6FqO2v2SKF2zONC1dYj9ARPppZJullBl
1Nz1IicWRNPUZ6jGbXBEfeGa7lTuzjryNGHxGV3d1DE3PGwMOhomgo5fo+mA
i8rbNlYu8tcdmz7RgRwV5tSs9XN2igVNYtyQqE9cnWudLtoQZbLnUB6iA0WY
ktVl+qay2gFUMubtuiFD+8Ymt6smFdHryCJnNfTeRNuIhDbLE2JsceqsiZBo
diV2yLKYGDC5UORzq90z6t/XcRngrImtKrIqeHxlemPMZU2fnbIMen4cSUfa
xWA2QUVJw6vbSFp0BvyQjTWm+OVZcg2BwHvOcEMjMFsbNPEtdgC8MXRW02I4
KJneYtAVQLpOxmAPhTI2FbJ0tg5T9FwU15dE2cxYyhT/r1trliingqFXcjDI
+Q6A9FpQSXs95ZKbEgm1f21tmdJfPjLZnbGYRNvKSlM0yW7A6gpHPN35kPMs
VWfwFoA76wk+9i5F1tg2hT8jqdZvPYmspomiw/s8n0mgL1dOT21vt7aaWxwo
rKl/YupsjoEQ9iN5vQDVclYeqvyZf+i0OBljhSyiHh9V4vjYRp2GWOgBAxTD
8A0cZmA2rCxtU5tlvRg+ApZZ85J0FRCjakHdw+2EXbn2stj5ILJW32F5UZAy
9fuD+DkevqmqI/AbdvRU7YLzoz3me4HvelUmqJKUylAtrLSRWStMd4SI6eno
A/oHWQD8/0aBzCija+wncGWL95aa8DvUalhSoTshISaEQyEolB7l8XJNQaNc
SaXIKwwR0zgaUzkeLUVbvaayVsjuGIkHrYiWw/OSecu/JnFYdntof5q7AzWD
jcaRvVoe4t2SLVrqb/rTSoIF4Wpi3g8bVf8cd32pg5LjBMYXlO2Wlc6sk3Rj
LENRnq0CeJOxPcuub1OAwQ4hecrMuEnepY+yuGyvYRdW+QFExKWCPIxbEih8
EBS1Pbjv7sxNoepMGl6HaAvPYpfZ6T84RhZ8ZuKdDlkf4gsOj+zXL0xoc6ZC
RQToUl6Jc7Q7STpBoFkzi9vyx6kupwYji3AynoNHyacneRy/Zn9yuEf4CzJ1
PmwhaJFOti985wVGb4g3Lylfvhu4Gkzkocs2tZ9/LuRIljdSUMYbjm3qS1N4
OGGO/pJgr4d9k+UkLUYtxD1EabwRuF8xkzhO/ZI/q8RRVLym+WkzIGXsg57o
VisHO7G7advWcDeyCCcICnnOP+Lc5cyk88q6jcs/hHjU2e9Dw4WpBTLT/CVh
jrce99I7bV0U8HBAMsh/jJmHZiQBkEDJtT0M0NI0DpJWwY8Sy6yu1N1+D7FG
5uXJy9mM699n0E8ftGDPMoul+wECizDJETDrYQLzkOkrZ1qxRVANVsBDToW6
4FsH6+r8olGLa1p2HH/3vdndt2r9ZJz41OvR6M2qNJJxD6Z96r4BiWVbbOOX
DCW/Ot249fWZHJ3wR+OCKndQq68Qn+gUiCbOhiMlTQxezac5VSe0wcRzsaMR
rL3cq8/EQoR3kkIyue+SMFJSIz1pBDvdM+Js9X+1bzc0iZWNik21GbSymTGe
L7WmCdGFVW8Ode+BJ/j/BMK5XxsubE0TxxAi5avONu+PaFzTMTqoxQoEavaz
JjkD4Dd/ImruWDr1y79kG0qL+l7XN8llCR5s0J0lVuukZMYmKfOfbQJKGSTY
+5yK6plLDg33OjH79QiVVhFzMxPz+PL9TfTPZAkeA8hGDEaUDyR8Mi8+EYiX
uuZVKWs9SJW0b0cOta7V6PlgC/3OJvkDl0si4VVk3mydHW1LXgs/1uxEUBWP
RTnK9SVbdT7pfryUp1SjUtrEAOt8VvFOT9Bpofppklf2AJViiMwOd1LSv01m
QPyI1KtvHrIVuHSmtQY+GJSMSR6M7yYieVtZBItHjtIEio+TyO2rtXrjtxDO
KGNW4otY9VWT/Bp2ZF4OgFIawyjN8W6LvxmYOOJpCsGOx8rYmPk41a3xt7L0
92ry23tvosb1iUpSNUbdWvWt4cBj7zrO9srdXjdvDqAyodL5intd+RuufPCN
Gbp/J/yK5ZBR5vsA4aO5uO2fHLIjApycDYsdulmixbVseFwFvUWcg5dn84jZ
7Q8STTDTnqrCG9g1CbBqlKDKofeeymTf5NtRNoNGLrYQ5uQBGEGA9h4oM15I
coRu8m//D3RhsgnVZr5S7u1Z2km+lRg/Jck3OZNfeP0xlr/w1A7WZglwR3Yd
OabkXIVlDaKXKMPdgh4dTfR9Vikka5Nq7jbW2rgEL5w2vspZ+QNLm84sQj93
zQodYtrCk2opY5avx+Fgxr/2Cwou1DVqCPGcTDm3bcmzGwFAUiW6BCh/xG3u
TWEolF+mQiKkzo3sBg7Yg8E3GsweD+dPnpRa9016WOEClpHEhpH2yqXfaa3+
8pUYcNsqEidj6o8XWu6FyuRQYfrmpWQLUIvsyk3KwIBCX4lwBV/U0/tTaEGg
P4vvl2cL0W9sD0lll7e7pEhXtxH6OFmhgbPB36L0vyxD1mbFD//mHaWO3/PD
WVxFudsooJdsZdwI5nGbFGX4otfkXfFHk1Ow1hPLJaIEQuRVW0KpvO2DQNWl
fczR6O6e+BoCCCXn0DGixDVuDXHhmxjFTQ8aTsmXmHL4K2YAVdoYGswGHWxT
soJSKkADUwQeWj18PMJXfS2k6hVy8VFFQ2qfsNF1z7JqDljVZglTsa169GU3
DpUd1J2PABuM/r72JS6NMjWvpsZnGdseCx7r2lK2P/rgrFHmEOHRh5LAZScl
u+uAal+nUIqxk6UsHpArt1w7TWwxyRM2Zej21Ya030Q3uPMSqUwLR3R2l+2s
VXdRjw+GlCZDN8LdBAjIeykeBVPjUC1H1w5EF6rDwLv0bf0TpAyIO9URuenG
XxV8V+oZTI4HHIbChMVNGMT7m7RmDSitQHJ1IskvCwvHMO2nIj3UVIyZBq6k
PS7l/gCJJiNYUF2uYyxeVJ7bph5QHjHqbtwb6JaDtrN5q/K8rWHxlC642VxG
ThXnZA5ep25K/tTMjUO2sxSBZ0ZE1ygGFPoA37Y1eHXRU73s7796npPZ6Dos
L6BFSikrAZaAzcfcI6q9WBk+anme3ZFOK78TzOGQ4EwdiumT72Y3a67pfXEW
dBC2s5f3ioRovzYNpEcfCZuq9MOmXkND6WLvKxtluNR7UEO1E2ypXm95qqoH
OpXiSPz1Ef1oXISTvKfHLxeJ4yKpoLkhG1bEYpfiERRQtMnP7icWMeeJLDqe
arc57lfUd/88ceBeqDA8rRK/RfiIw+SQESBs5fZlOJUxYGrQZQOnPB/5Ujt/
e840Uwmt6xM+1WaiqorzbCdjdtO3ExBWxE5HFOOsga2mDJcVU9t/PC1u4BgB
nn6tBSZ3ZQvL/OcI0oB8/tDnYFqh6PMuwvvtxE1XKmwQO6wpCffVc8Z2Zp+6
cekgFyuouwzDxlccj3f5cfRzf1xBCMgJwHSBQ78RgQQp3dxYQGyclEY3r3o+
ta00XmtHybBwlneH5W2+SplALvPGkyRU0ljegWerkkeS7vw3ViPFgMA8HjHA
IqLK6rBccGGOSrwiEdb3e+byC9VTllBaA/p+43mlrZxd/MhbzT4hG0cnYubG
L0FpWtDulUtc0Rnrtt7+B5XgYJstf57+O6cWG428hRhmt5XCfEAQoYim+qre
RZkLLGZenc7Y3JGtlwBGWe2e5jn8vzX+A150qdNvtrCIiiD6OiTyckc2yLuk
WAdgj5oa89mzLae3FEEwwHLE2C5Ffhp5mQ2sg0qpn/EsY46I31vF113J4jm9
vBR17PPu+uVA9vV0GTvdRjTNleQLiXVIh2xLkkR3h2zrrCt3Bb/W3K6jnSLO
dJhaXVm365PZ8CYUKtylERY/DpzPPawo/dl654O7odmk5yOo8dZj+9sjwypU
o63cbFieXDgCT7QZW/ceMf8uD4WnDyMv6myoSEKI6A3SdgfGCK784qSIgYJC
z4LtMh0Ux+d/lFvqBqsRk+VEFcSNnHZ4tvdQ9uexaeDr/KesVx5Wp2DPYzHi
Bf240bxeXUgbPL5zUMuq63Pa8YlNWr0klF7hoKxKAz/OKv4rBbnKig2EBd6g
8TC7j0inF0V+2aALa3RVzM9ahhSHNGIO6wVfYbQ5B1y3W5t3XYMfr0KI+FAe
itPHxY7vis8RA5/+rcI3ssYMVmPMuWeuENMigd4vR4B23fET1I/XiDRPfgXt
+wD18e5OrJg11xit1+yUUvkZJ/i6rS4sttj/1Q5lwsxQrbKN4FI/OjaKmmkn
zydJQTBSil84+FAh+8wV/Hu9SBe94nahqWhvA4P/4fj25442wY1McWvJJaBn
ThwnQ9bYV40ogjt6gNMAMY7IBylQNVAoa7q9PpUHQSLOAdinkoZ6hjCqVeWi
TeS+ULFuJAJ/JbHSQqDKbg8GGNPHaIzVbgV06jDNned2gF70KARkiynMy6I8
aA1HoB4lohNBeSG4pYbDkUdYxy5prOVEc6GLvEqKTR2Fty0pydMwZPqlgP2J
z8R2hFnJUgfFp/1agfadgS+uyeuHT6dqNUZIstreq8Zg0auSxYzqXTnghnsl
VgZXvuXKS30/dZbYb/s2pw/JEo/4UpSdv1hQjSBiXSUXmyCmEIvHc2wbxgk0
DQAFTWENZiG6qkozt+kkgWOpEheX5rVcGWwZsr4LxCMqTSRU55Ux7OoHcywf
ZW+9sq6aeuUGxpTxCzt3gSwFiD2rYsSiesRjsk6KtD9LCi5ThPKZxGeSP98G
G3HfxCaf+MGcZCdQwqi4DmHLnWfjsS55JEhHYk2ft2VWHBiJCJ/ZLk3eu+kP
CqtAdxVY6OA5pmIECZm7179JjHasnZ6sRrt+ZaRR79hfyTa25HldEAPQhkpD
xeNWT+HrUaGOr3bQLJ2SQIheFdh5vendx/kQ4S9T1HpZKAaGBRkxozwGOXZr
oJ3rgHxjS7NHcmVY62y7U+TxF6cyhoi+43NcAKKBE8nyPpcbYG3lAw6yGrT1
OAXri7qUDpgBN/FGfxnsPciuGLHv7F4pA0SIuguK5NwLSRydRlWtujbkeIjQ
4nLyGKaRNfdnfKo20jwto68RYYt/eaOFDfFyjnW1ppbGQirCGy08sKtsiAC+
wDPl4A+FoVivIrDNBbFdFDikdXcNeytDtfRrfHDCVHHPxFd3wt8ZyLBxiA+y
U0Npn62g2t6TC9NjYgJnLcb9Yr+wj/WGO6YIOkgdQO9xlq8SW0rxDvJshPK4
ztlPQkdxn+vqqo1Y9+ysN9rWZqQetz7Z+2ZOgaLltRimxcEEDhpyjkIsYnPj
9WvITii4BMHLBCSbmTDKLEZoysL9r6Sy9nQYl06QaDeoWXLlrnCShwSEB6nT
FHhjjaSL7OAWxjcjsI1HEacmPL9Q8AI4FC4+B0DA9cICVe9e6Rt+H8TuBCe7
NX9oGTOrcKymBj6ArrfkxJsCZ7Lpe/BZhlUT7MdcLOUdvjtZqOYF4CS+wuf4
wtAhr0slCRS7He89BKgHSuKv92sguUTZt1pV5HzDiAAEt0BHIJMpePaLHm7W
oUqSb1zgpmUBUTolus3ruJcRXs/i5IXl1FJ6FSCPDLRDPN8RvAvq2Se5BHOp
f6SwPF6t004W2ihRsAxKaJgp6yMzNhYEaLlLsIyaivGGg5duWm27l8mCPuOh
vGzIuGrG0kF5Kr1on3YsmPLRw9ELkugc1ffNGq0G9mCrnxp/5rwBb0JE5hGb
93z5hRTe+a/1v8T9dOSbgA6+N7hHBtu4f/8h/Lh26s9Sgn/0yglPHub+fXld
1PE672Hteq63GfbpjgBtUMt4Xj4ct3xet33uvJAdIyfaM+bZhRJwWozNwPzZ
FLKz4xjGe4a9nSYBo96SsRwUNxBqbfZ6w0UPR5SS5JD2VDWiTxXnAhxg5w7u
/9JL4wxYQXwr/4U8m0UL7GZw5yddd8onAfCIfzInrM4h03wkr8PJaSEwJ8Wh
eqD/HnV1PK/rafiasGxxwk/A8JEU8Dz+o8LwHgCFIxbdB1DUI+hkJm8A03Gp
0uN7WajaIyi8X9ih9ceKu8/cLOl/iXysPyq/sMv5Z6SMVBvP1iC5tVMmpixL
wrXC4MT/h4pqQ0WMIQdmULCpi9UIBlsekiYQmtyK6Oe2H5OvsXs1fu2tQXkE
7eucSnp5JaudocHx1+qg8OcqfPUiAaCHUm29uiFFqNgMWC+ZJaaGl68DuTVJ
vX6vrfA1SSTswGV+n83emzMAtSDvDFCxdO2iQiIC84ec52Vl+PqDUaQx6AYx
MEoz4jbuyt2tFP8/VKurAOMZ+CuGswMforbTHfuPknir54ISGz44uT/0ivkU
Gi0nosW3dDNTqjGiu8I1O9QeGDWdf/dQGE7RencE+i1COAhZRubrKuifL967
cTjUs+87RoIUBPLy9wBQtiQl420c4e/w8OVIagCjS0XXNjjOIGMa2SxEMckP
OiyrJtROK2DQnPpsP/oFWbZckaSRqWsmoyQd8S+MtVAyEF6YP4ulcByc16Pe
gFkglFlDF5gLWlSnr4RIwrwZ6jOJXgLKPh4mDYDYiq6nSekG2NV9VfUP6pfb
FNtekFA96OMLAMtfh/rJvYtQYxJ4AIITsqf3BZ/S6JrOKi6yjL6zmzrY2ug/
yMRKrGyhlaUPbS4UGr8GdHJhuu/8C6OXGUVGP1x5btHlPQDpQgIWrErx1SwN
BN6TMxiBhEl1efLpIX8e75z6+NVLyY6K7tq+1vARG2xDPpetZL86Kibgdffw
5ZmjsSfRAtK0b8F0yxku2huryU8uY0eIKiKnrh4cTTU0UEVVy4EhdmbFT8Nm
N2pZjPic/MBlRV3MXI88fJwWN9jXtAHbI4l7+3BTYXznGr5nWNzU3oHEIaEP
HY8MCuFIsiLyfq/L5T3SHhlP1bsSkba1E+06ev02aijjzbKUP1buGqtxrorj
ljDmQne+fVXZWBtHprSqXPLUKl5Vl9iDi2wtB68kA6uWyaLIpJf+5flPyyle
pRi8FJMjpU8gq8lnAH24oIAZIWMaLojqR5w8QwsNhSPwrwNbuvXyCxV1FhBF
lrRwEkJqOEQva1FYcNxekjkqyxhyNAgvPcQzJ2jAAszZmojhJ5dcBDxPOPj7
qnVxIG0UwkjHx0zDn2u27+53tU9QZrP7SxQzbD5C5mxy5spkY5bnNnzydl1l
IIc0iDtJAeyypM2I5E0UVpjZ/3U7hXkcz833NAbxssRpqVDXE5WMrgiPZBrr
FYS3ff0czknDJfXangLcYEIwwQTC5BkUFLuUpCJ7JOXCSTGHW0+y7epTLH+3
15/TXj2phVaVdzuL4gZxl18zBfzrdHAHVjQTWHrPPONDJJYKAT3KlCtXS/Bz
darhfun5Vq5KDrGbQAsY+1djZBWXMqrPL5h9oWqPGIFGefat++GjGeON68Js
aPDhNHJay+o5z3uJf7/uwge7nnsjDjbEt5CA/qv8LvgLbMsG3e1Qlqd94Ckl
pRe3CkoR/8Lz0ere7w1NXfMV/qz6POBplgUMSs/0kHyIyIlijqRhuZagvC31
M1r3iRMHCupYJBlzlZ+ucrpt8w79c9hes/GIXsKlVDuAHKSMxw74jmnV+cvv
jAW28eO3pCKkw4ep3vJhglCR4P+O6JFN5QbU4VPSHJNGhRa9iEtQAIWiO771
2mEvAPhlAq4mCkHBlokjqwglOImhk+2sF2U5Na9/e/8YfWlzmVqET5LmWcrn
5FBixMqoLEtCN7qmaZabZc6tFga1s/b1INZjxlaBG9Mqp1Jxeave0LY2blzW
efnbbgGS90wvY6FpDSD46fk0NlAfKMI1YshL6Th+55t9oLeOUkTJhYa/I4x4
8O6zciYzN5r4fEQ21A2sMsfJQbXzG9+HOL/ArBiFUozS/qKUWiLqNuiV7qVa
0DJSxCdQurQHxgQ/NsZZardA5XM8h2bkCiCnquYyROSwmLeoENOaAHeglALq
oB8hrzobLptYpd4zRp0xyuCjt4Beh1KAfdesz+//7sMPpbOotOCVSr9M6xs2
tmzp8unTza6DhGv+9uqlld8L6PendW+63zisgo4SzSLmJkxSLW7A7k9IlWHT
ikxvMIg4ThnIFQHL5Zj33dS8x5P0KZK4r4uGN2pDmNgRU+QjrcP+XIeX0xQ5
AR3k3YagW7maDVRWZ73R/2GtlJXeCZYHuxTIAhYc0tPc9O3IybPhDZfsgKi6
GtKIn5W+mAuNMGrTH21haQEjwBAJB8k0jlDMeoKQoF14WSEe1rzVODdEEmIe
JLGgtHhJ+wTNMhkDrUnQKBwR7iPtvNYnRO0WgOOirxwkYeigotCywiCp2cJ4
H2QlUCol1YOlizmfoZxAe5yGcfW8eNedn5Bel0T0YWt3yc8JLod9VVgaVuy8
C+hzP0ZsNxSSFZlLVEGkBo0C7e9Wxza0SHCUknHKjRkQNJFC17HIApKr8zyf
eMNv3zFjGQzRrdjm17lX75FWCD9ol9+wb7+DMJ/jHY9zNpFtVutADuAgQ9Ru
Zahah+H3DAs7bXNovyMf4X4icEEeOKeQb4nXg5/h+cSQPNMka5fLow9auD5d
8fjaVOwj0WrqMa0gQkp2Qto01t19XJmB2PpKsN2Ur7tWENU0YmD0g+B+v3k+
g1qxONeUAg4hQaHBkQhvGYK89FWQWcgqfd8XIbRfwNywlwmk30Sv3cGaDYbO
TB6uKew2xZN5OZJy4ifHsrHSazoOlE778QNH7hl37BCMBtK7y50tC7j8g2f1
hX+r3aKZcnwMHpg4CJInNNoA78y5OS4Ywz1ZrXfbDf53bCcUWcbQl5++ScKa
z4qTifq/26twPqMrCAqDZpNKXvlH9khK/CKrm+Pg2V28lbjGtAmbB5zymDQ8
bApT3okK1RBYOwfGb67P3/Nh363YKfibyA4YdnCnF5GZbMzNmdulUCjVAo/a
iGrZ9KRxfanV8a1PZIrF2L9f9ZCH7KVl99uvDaHxh/dwN1WNVYPt2a//NKJU
sk4MLcwlizJYytnnof6Ylswt2LZ4NXsxP3tQ8eIZmjOWS7Bi5h1vYyxyqGpG
SR22vGmki1tag48AzqJ1p30uloXxVoZ9XrdKd5xn9s5bvb4vfcUDT93mMa3a
h1P94dvxcD16YXcqnAZ+8+ebVJESd6gVc6RUxLoAft75ghYqLOiOW+MNZYDz
rxbp5QL/mXXwkj5OcJS6KqLq5pYJWhxCDvocpOE+s+LiDKtIBKvNfvAshWtN
bG4wdY91HoCDe9Tk/e/sVOfdqityWtJ8zFnuhk0X5US3KUMclIfGrP1Oval7
11csIgMwvHbufKnFgfudbqGPI7B1uQgiUu2o2k5Fj8IHsV42T1AV9vY1lpye
yLiQV1g3bACoMiKfgLTjAxlPfmOdYzleMgfkJdoRIyujTjoWMGuSDLVljZrz
j1XsyRxnNonv3Mvf4ZiUXqJAX8kvu5V1F54A9QJ187JOepIl3B+sU9elx9q0
sTG1KCI+8u1kR/igYChL21uPwMfhuXDMw2t3RNSOp+Vu8CN2g/CV75w7EoQg
VLWRAvgWTWENB/imYbfpAFUT6Fp96r9wzsJ98PX9D8QX3SI1++63U59CZ1XX
6RczCycvM7lXeSf4liCTthGSWB/kYITDwygvXLB94mUS1TjZKEvZOunwJ0eh
12tYf0AXdUcTQ7pJlX1YiXdkVvWTKu6WBW1ZCjNNjqjopudPx1ttBY7p28Bk
+NxHvw3Owt+/bB1u1PIWTGNZRyBzTRmX1sGFTUqxJwahOKT0wsr+N65MHSZi
xTNH7ZwgiufXjIb2s5eYYS34gqtewQNkdajsBQGmmLzcExMGwULaIQIjysam
CAqzsMgGpwL8xg9/sqyV4RljN8H9BtDW4J1wGS3uRmtoOR10pMx9ZPnZ88h1
QeM8SFgyhsrsfE+7h0WwnyfQ6ZoiVzDKsiV0VgHNP8RwadfQbSNjSRdOhgh7
vNUV03/D1PY+2r7C3Hrm6bJ9cwRKZdTXb8EQdEgksZvVI6btyfg6hcIRNpyk
dmh07nyfBuIlDfuMlW/0t5Vb0B6cTnOsRHDOZg640B0wJR75PniGXnMNeNRZ
AWkzT2wCdWw6bzju0BBy6Quh9ewxXvUESlMVLN6uM+fCtD5+dkks0EOi4flP
hF98Uv8xyWb/u0l9QMV/SX/YZQJyrkc+6lOQWytQn4t7s1SjRhnvzU071bQK
BYyaYeMCS6NNQJng/RmXkGXUouK/p+qfge09WrIsaAUuiMIov7Nlvh+yObAC
+z/yMTJw0fupg0MtHBYMXYh9hsTxcQCaQi5TMxQcF3DLVZ2tOVLNQdTMKX2E
BG5mDoMz0tHv0AEM8FNPwhBQ9y+ZTsExX08Dj4aNHcsXC703R5X8MfmlAP7p
HdsYnfbFwI7b4JKjX+yvE1GLIEKPYu6uGyZ2dYv6fLUC4bEF9A0Gn2mOVOLj
VpvrzmyxtaUzzkz6BNzRjAywPg22M0RkfZcx3EkL6hoPhYfDNKpfoX7U22gE
kM6RfsOasU5O++DhR7GvmnSHio6ifoEtmbSrZ5spHViR3qF3bfKStL9x5f+E
whO8I48RYfWElkN7lLvaHXfxLBdfbArv0HK9I5Kr0q5C/KW229mxH4PXI9gt
BxomoaayZnV58Nc9U+6YdwjxKzyKASA8z6P61dg6n+hMfCi7LU755QkjR6l8
bM7tdrvmPS0Ow6X3koSv5pzmrGe7yDqvJwEyq9HkbDP+uYbVrBe3SfJYL1+a
P8PXlqLjKCPiL14YFpc906MoWS/nvhZgZC2sGAicJVKhRhoL3BA7k+UD5EY+
aFR7Vsuvp/bU4eiMZcl6uExR0KscWMaqZ/OYhLDW9etM17CAPcudqeCVTsOv
ncLy7Ue8zS3zdG5xsFLoZ/sttWKUefeH7oKz6p1X/pH9hodZvXTybtkaeMBX
T206kV0peGunAHZHh/7lQsQbaGQ3Wzs0hLXXFbUh8Gec4VkVvSJeCQptvFqh
kfMzQi+7orc7g4rGREtBUtrj9gewL8wxUllZxExnBoyaMNGLmUCxEP+wiLpg
j/nidMC5tv9cXS+SShTe3TOzS2KQmJqiy8SCZ3A/+lTFqsBYAFNhUW9aPr7D
PkGuwQBgldXtZfZW+SvyFf3yGAnE1ZFfTC/wpEgzb0TD59Y12LjzmKBnfkmo
PYvTN2TSBZCHeFidJseVpM9bIwEUPMIAIZlCpaR//eymQ99etnDXU5Wbyeu3
egcb92Xsyald8jGC2NF0QCzwAsM+IsXVnS1UXqzUjqgACq7daz52w/XaUTn3
KmhA55iNZ7B1ZB9T+0+gsET1BepX3gcGYTs62t3CRWbJYuKO7ocVFhzRggCB
mtuiKg4+A6Dtusa+ofeysE22QFtmrBc6C2Do+/2UsJ31XRVVIegc8vH34gy7
YvlV+UAuYmD1yOowm2zwPnZoC9P5G/Vpkgf9onBVvS5OMUS6U29+51CojonR
Efca+4ENX1K4h6STByBG4MvPoYX4fwDgLHkR0qvVSAlLigbaniobCDaGggce
/4et6RcsYKlqeJs403bDnsuorTHvg8gHbku/DMUyQ92STRHu1LYeIXbQigQa
nXOjbMtBI1w9cum76JpW8wnuncC7cIb3vdE46yeud0e89wNovZe5muIYETby
ZgMIti20vVxD8sYMnC7jlVNIvn/3T+QCP3yys7XT0q3Vn0O9RC5SbruZmq4t
L0uLG6H9jTHtIVKniJZT3pp04p4RbCHh04jG0Z5HKTmV0d+mbGk2JloSoqyi
3UwgCimRSjntnsz3x3IFmMeWTQexoSF8cwXMk+8N5WKdq4/h5WqfkMJx4smo
wV7DCNRuPqcTs/1wViGlumkdDmX1k67JPNtsBTUI6bi5kiqaCMzDdOlejaQW
v+d4iaxp8d7O3PWJa80kR2AMcyMJ9DxLiUpYcQ/QecC+qldrcuXzeb73GjBB
eYYglf3yytzQNsFhyUqPdJwExRTrsdT2BPh6aqlw6qIHNUyBl7UzD0fSUZGX
Zk6DiTueGg30TK6Zyvq9FJWbDG8w67W1a4mT4NdCFBIicpzOcHQNA0P+w3wZ
VLJN+ExtX4Xm4q+cOdFCYLpleGk8dGnZGQ8VbSyyq+wD/USpiThTI3XXz6q0
fZnih213DLNzKLz4FoN2TybVE/HyqBqfSFq7gtyUAxERTzMTKra28O2bXLcH
gPyFNcN2rUT83yPIUNxmgKGQdJZVaHyhD2JPOWqAmyPzb1c5Qosg8xx1XmAG
yfO/IbMNktD8psj0DJm1x7Dysdj6MH1BPiEjkKM8wK67HYgChrBf7P5/AJHE
2/mHXb2ZRHwsaAM+6pHDScdPrgMswoa7gCnad61eq6VqcpKDfznI6wbRWhwY
HF6D+O+Ft4CFlQUe8Lvn+Z64rBx/hN8bOF87I1bmgU99FAkzBY/QqEAT/iMd
N8IR9oF13fckCknKbygAGawLA0l211AdNsoYYC3KhmBvxecyRxa/wvsL+VWk
bhv9uvONXgJPcSlpDvJaolxcF4oLFOfsUFznFnFxlvpQr/su0z++9Db3Ls/O
B25t6Ct4zJngMz60sxUrTMhhv+o6f5fey74tbZGSjfYoLe5s6+3/jxF4k4Ap
6KMYjEGHs5LgSjxaEfTlcbOUEgrMC3dn4na6wNTQuI51yeAoN3N0bNQJcEex
JKkmrcutDyd+IPB9cOx8sKT0VYiWNSWQ4V88pXeGB4StF8VD0tBtM+z59J1L
7/uDJo/bNKtSaQsBIAbVrI43t4jyrpwmnGmQszX7RbPZ/ZgI45Hlez3TX2cF
IG/RL2YBztlZlzs+Hggb3TKG3nfDZhcxyKW3qW7+6fhDT3M+MksiYeMao8Tj
jWb9g0vya5SO+/AoJ8hiQfeveUvEcCjxbk7qtxGhZz7v9i4idySyZVyUcYbE
jz2RVhw1lizQMHMdb1JlZLkSKWPzTCh2Rf2utm6IcsaN6A28IXdzpTB4EPyA
K68AK5NJSvpuMVJEfrz9qiFyFs8heH5yYJkU02YqVW4GrC4FmePYs4EjJAup
M/kJD6+1Vz4/eXSLFJJIT8Tdr3aZUqiAFHW42en15L9jR5whA2ur0rtNwLpk
qF6YKF8SeCekOePdnVg0YW9vUytx6zjMEMespal8MBaDhLKzdLSeJrW8O3UF
hgjqyG7Gl1TL0M9V8s9RMIsHkpIgpK1w6iNNV0n08rBXogC98A9LLV4uESkL
sk/PCDLWWjSsFl81OrDaUcyKREi19SyijGBoBt+R3WvzB6zfHOUNYmhsh8yq
PXN1XkaE4NHvhHDOcTSMWGYRQ5yjd+ggO7J7QZRHDt2OK74LzPJ1/wLN7xik
iNcAA0nfSuBmq9UmpdqrkeSyvSn/ggGmF8Cbpm7JCVdMyQwVOGWUgLhSytd9
qSkCuVAo2doRGTNRX7X8QRAPLuwBIgYdBB+6JN8tTlxSL6nf2OxoVssjY7sS
AHFiU82LD+w6XnGVjw5FH1Vz8U60Y0RvB0qVI81tFwAE+DHntGUPuoTFJDU2
AnoiikmJuU53I2/Tq6DikPyfOaiqkh7jVipS+YljBv2ci23sYJx3rXJV3/JI
ThWl8SOMcwg/ZYHPqwlD9K0Nf3u1nRfdTZBJQQjy5MvxbhFA6KxZBcofekZL
j/lM3a0bdmkgB3pDD9q29K4mWsogrHsCf8lj/VsSez6lgrYRNFLTAlfONyT+
timBqf649i7aP8BdU6mBkQifilLoYc+pTnJCfl56hpz5firotyH+9dJdqau7
jcao1nAFWkNMcEAc20qw0AUDriNlJ9F6jTp9OH0SeP1PyrBM4SoJW07MK066
sGS6er+nLgygbV7EpXP+AQcugDbfcAT0030gjqM57HMT3ngav+v3rJxaodsO
SibpGu0+VJwuxHDLTcXzOm0t9kQCw4Ydl3o8afgiB9YKqspCdzDrDLh04d+h
gSW0xOoE6xn+7ockpIVaTis2DNrisoQ32VOJ70ctYrxm5w3jXc1GVpg6t3J0
u9h9QObvLjoPsWd6KNc4eWXElc+eC/6LFAG59xY4RtI84ovOWcP1KpIIU/k8
1Ui5UawlPY4MaqHPgaXXWnveNSwPF2AemjznPHFLSershOwn0bfB1XL/BXBa
r4VNVk2PhZmKYWfi/9UMqf7r2kfjJ/T50lE+Clb/LBHR1eVEthMUEL4RBA0x
vnycnJPz5g+vmx0OGhWLlj1Qmvl3DOK1jSTf5YAHmKpy9C+hJM7gb2IQ0MCZ
FQZKo0e1bbb9LM539ECuB8v2oGgILiI5ACVlZYfrzu/pJHp1vYKQ/9ez7y08
fOvb7cLdX4rdPZulJlKbteB3+1rAIOS2l+JFe9SuUVEQbwdkclwe3ARS0obS
JNLlakAu4zWZuLPlJx01C28bmeXCY6tw+MEZS2i2CZBHziIxVNeTPE0Kbvz1
tCiB7Vu5HS0sQF0LtTZ8oeo+JADrXIck0FiLx/FRhkOwJj+cNltHA4VYzSi3
0P3wDU81l0Il8l+g2mjDLuKoXypbqBT6yKfMPH6JkDUbey2N88sv5OirxnDT
J4B/xVTKYP8bPvP5dWI3NDAZ/nRPUGdfhuIpF2R8TmHwUMZ+dVm5zIaLTf3N
5DPvVXJsEvi61/HDe080ctBTU1PU+b/bxYIyuzY3CVwhlwHuGPsConoaWfh2
m1i8oxWicSJpA9heW+ti0gpQcIIQtoabEMVQF5pJ7oWbcC5CJNgfiQQvxR1s
Zg7qFJotTnTch1SQcdTx3vWwWV6KelQowmOoCIRx55LA1r/95ovvQ/iFPsG0
W554/4MfgMT1FkVvz+TovEyb1+1k82w4Gs7nV7fxBBmG3Oz22mutR4ur9tXw
DnZcw8n/DDX+XWfK3aWVvSOYFaxFLMZ+ZMZrI2eZwU+b/BZ6KQFNKbEInnGK
tFDAtnujFCPhhi/M9vGtD0ytD0WyUMneSDhJNcQszKRRKwUxLrn6rFIXn2Zj
380x3XqEKACMtOgo+7CiJ9XwOUuNDL3RXXqLpadeun1Ew+C9ekKnuUcF0DCX
oZ1KK4edllgPZHKVZPVerbSQ2lFzPlpe2u1VGey3lZ/TpTaZlylm4IvXunCV
LBUl61hVuxZ99NHogBGmrM561gXTMK/SJ6rt3v+NWQnzFRJaMB4OVh1e46yD
qCxc/VtdviDlQhFACv7rNjGNP4ToN6HiWtl6iona8MtxIIvYsJFyF0FBQZK9
kLRlEzLaThhNpwbwnb2ZgLKdYMd8H7etuTSz3xE3MuXuQftbrbWa5tfDDh4+
eYLfEmrLDDyZ3ME/dIa2GwAeuZcABnBXt13u0nmTugpuMkj/xujlO+gw5SuO
6Em8gd/TKAoBHc5/X3OUZxLoSsqDMsEjIGtnT/M7jbOxJJMu3MnwqLhE4NSo
J5NFxm1Ld25gKCeJeLtOWrBrNgf1laia0+Am4S3IeHgcI4OvJ1Du1gFrSDZp
WvJqiVe60av9vXSDeIQLZlCJ23azJgqYzVGFGL60gU+eLsXpC8h23gpqNTSm
jOV/ozvd37zniizq6CaY57QfwqRRgO83cmSTdR3ANRYd8gu0+PszPixF/flt
0z3js56+00oepGh3DOExYMN6f3zSrocUl7qTCjX0Ly0uVwkPsY0xc6JsUQRu
DtLXQYbmGbqmcY1gwqMU18cgdS9/LPotYDD/bJe+TzVX21/fycafR5v65SEo
Olwj9JWEnrjsUTIbnBvreUCi+QfZ/qdb+6h9XGe2ZbRGJHKMBauqRrll2ibn
5z5T6aEKpsixvqoYhJFjOCSkeugVWXiG7pBIfRwC6Dish0Ps2uHtQlfykqwm
bHsW3SRMKIlEHPfPJDHifpPIZkFObhYHvC1B3Vj4XzaezkWGUpwLQ8fWL64Y
758aBa2X9MV7lKir6HO5hP56PQtOjiAjyinsYmJyNjIZ13579C51nc4GgEHL
WMacooW0/jY8ImhZS7FE0HJdQon3wUnHuqbPwquepD0gWEWyzdLhc4SxomsL
RRBzcL7uinDuZNEfrmPiBob4He8TvcD18ykyB3MLxX5khbBWvo7MN6dKLPis
R+6iBhC7XR7jRVX0MuDtKK7gyV/QGBWbl/EJNQmQFGfVAo9L6Y2c+sCOi8mL
VPC8741YkSkBOpsuAKZVsYXR54tqBOUDmBnCCgw+Pr+k6mc7jN5pobDnZHHR
eYDsaVDJTAJBxB9ATVm1f2dlSjj0mcjK8O9oimrleKNP9bHegYNSkALS8Lap
5W4GKnwzXMxHZrs1+vqSLZ2UVMLGQ5iusOEPzmUBv3oiUslh6Kod7WtwYwA4
K41KTGe2LkGLHG9etUwMg84OMRJ4Sju0GbQLqoeHtCerbDeVxp+7KOZVJSFX
oyw+cC9eIXkbbB736vYsyECzSORoTd2aBD7LjwL34UXco+qOSU2GdYopj0Jw
KJJlw1aV3EIskbUv2OKD7g9qRMlGiyJ62OGrsJ1BfxUwBQpIX4FjQLPc1p7H
8A/6J+Vxo1xhzNhc+JkmHC/WoYrFO6Dh/t2tCxyI59CWFk1Xh/vWkMHD8ao6
5ME5DsANIT9BOGAPrv4xm/DOWDOHqXomJ1JIH8/DP2Acnw/iJ98Z8p1unIKn
bifJIggXSCdT/5SAQw+POAkci7GTzMXg/lBb/BIS89jJinGkTN1j4OpkE+DX
4XeIwmnlBp8WjlUHUVpxc8zMsMQDHD24+nL4Zak2QFa0z2J8Xu6wHN1eCMUF
n//brxnjvIDISa7dhjKCrFACtXzqt3PYlXay5r9FkyViNK1YkQOUHw78NxS2
Nc0ju1YeHP36lxH9oeVIarsKTVjXkNjssvbuzmG46WM72ZKaP7iNKQtT37LL
6W3Aj8IKcCREWN44HhccKOv2ezThvHHJuflKQrhUruPkj4FzQGyKFZDRceya
8DHmWJIQ7/S6JUtKNroedufEll3MLQ21WtswXbpwNTivCX9bUvMIzqpg2NIx
5TQWGPeIOyqsFXN2H+sdzb7RnvCL7ZiyMVFbi1HaDKt0vziTOMjevwudEVUP
UqLSeU3dPVny65mya2Un6ZnxwKjLmVlCE+rF8McHCJ8gzyeiC6Mld+Xvz6gq
jt23fAN8SKs8ScPwyhsou1qoT01infq8L9QGPdcOsgRakdfo3E/As5D4GcPD
0jDlY1HsFamE7ldZ8ZFOaiM5m7ZzJwymRGOYu9l5RtwzkM1pSKBgXGVL5ceJ
un5kcxoVr5/dkN6O9vscLP5cCD7GTN7iRphsaL1hp3R03M8lsyWg01z26gu+
sdAxBW7tRaBLElTUqcHLSd/6JrN3JAZOj41c4Q7iXfmcIMfw8fN5XnGoAJWk
N3p2B8rV8geKL0ihf11tXH9xDoYjd8b3h9gdeDqEVDSza1LeUur1oWn8yvP9
wzVWLjg8sgy7pQ0xYRHnKK1kdrAHzgKNTPXOE+5GPIT0hsuusarD4Jdxl7e/
ma0qEAuOeUCKAwUlD91Vu9u81kspBSHCKO2WCYgN2GxGEBPirovT8nzTUv9F
RfywlrTKgN4wqK8o7j+W/QtH/kszOPXukD7Mu/ABtZCybgnGZGxcM8q0wkEm
0yD2aqfvkr50Lt7uF8qY3ywYUhxYp7esf279ol6C5CMbScmGvBdt11/FOHVv
DRgz8oGDbGM3ju+kfnZPko+CUIk6wXe5eJNKXBd5eKUW6Qhjg7VFE52PjAwG
GJpeOIhWrETyhuwK/xG8xwvKHSMoJOQCbCQRy79rQBWgmMN5PFC2K5thgWiW
5vlnW+u1K102YDz7g3Z8SfeeudofFGgdKooehSgj5I/VEdcmvxbAb34ol3zI
eBTds++6/GLZQDEgk5/CRQJlOMejolDz8aHxeUfOJSVQV3BU9yGnY+ld2I9w
h0WKN3/0ZxaaWJqfqrqzbwLxGJx9zVyt79kofk9IvM99a0FDJa291TwD4IIg
XvVeCGFHmktOgkdqH+EyljpX2FwaWf1dnFMdfCltQ455UZzFxg+QD9DT4jbL
IVSvl4E7R4lYR32XAn7ypdVrkpkNiThE67qi8l4AYB0Nx94aVei6+xHsKs8L
7p/FjWRpfIAeVKrrCxEtHblk9Wd5hvsWfKXGWu8jKaucvZVdVyVNk/lE5m5t
ufrCHqiZKZSt17TWL3smPpc9+sLALJk5Fn30i3rW2XrWuWWJ4ybZoG9b8Zdn
/YGC/T62ncuYXrMk7R20HR8BvJBnlUV2ex9uXoqs+aXWgA8wNL4AkKfa8buk
yXl2UseV6lEKRbXRjquksYdiCJlnSLufX0H8h3I8hQahFn6u0uzebn7zsAyZ
cmsrZVv/gP7ahm45bmeQHtXKYi1fPwKWlCF00hpNAxN4N+VtQ9GyKJhjjYZf
PIRHMV9BfS7vQjL7FUPACl04sAWQ8gYqVF4C/dUtXH5pVhNTas8H87oqkZgr
QdA8OX0gYqUKw0t9AJAoTGX6v8kq6VT1Ws68sknNp7fUPlgU5DuhgEnIewoK
7Y2wtKFWw667OiBQoy5nLjK3+YiGWiFg3OPcvEaI+9sU+kVY5DoBHWaIUq+o
HLteMvyylXpi8HZ+8ia1EJ0HVJUGFqaeQqUV2/RsT5TI8MIqV6inGankZm6b
gjnY9YRvgqAHJsCNGJJEZzy0HnFVBJvCyBXQUzOSctxAvCk8tv62Kax0vZOv
MXR7dQmWkbWxUAJxD3SyN4ynSBrS5eJ4SCsCaRcgBGhv1TJDczWbuosUXSuH
pBP+bMW3Mx2L23P3/imIfg+DiAoOllQKqKWoFhzS4NAt6OI7b8bMfzIZ1hz2
kCl/GNVyH6ZY4X+IFQVcWwatAe47+bTm2U0Z+T0ZGkgN/UZiCRGsk9k6n8R3
xnPghobV+fR9ffSbVsYv5dj+qo5naMgLgTMUsam3y/IPoj/QPD44mOlalpmD
F1mwtrqLxUVbzDvISuRraebsucGdEX3yjFheXiOaBHIRfz18V/zIkNN61OSR
FYzqhiEdHelBVxJwxKno48Fajfz4NVSHGzApUvUQmx4cuXKKNWlwqyB09Y7R
wZTt02MCUC7MHrDzefDnuQZi1T/LojVp74xEFdxn9WPWS+/ziKneHJkwD7Le
2EVnzScBIz1oRAuMEBOfNk5dLIpB9REFoezikq+oYGoEWS9r3eUYk7glXU3T
ntmi7W2khSYC1RfiIUZmSmyoWFOiQRg6vdcRKL9lZF/q8ljrE0oNeAuNHIgZ
gAoU8i39k8wGX/fD0cmE1IUzO7T13VRFD+3aIiEmyyzfDoePEf5Ib4ORxtt4
8UGnaQrMy+KPk6pxjhNVPyHU7xYR/UFJ+UfYz4X54kKVlMgY35ZPw0/ahEOm
x/P/gZ4Jdgx/xE6INoYMX9yCvzLUrwIbKqMTbnfdXo1Y8hYtVJEeMGQi7lPl
I+8XqhD4RwpvjCY4yOotGe8f3WTvqKe4/Bsg+2DO9gQgq8uM6dwcV0HE/6A0
YjAZty3K0M7tNFQlf4pH/G5hWI9DSHYhLwLHeSXKvJleu6Ju9e3SJq4o+3C+
6vxcNLNAKsofKPHeqtcSc66Amw3ostCcAxE9w2HaZOVnLHhdue060IsDJuH+
EKMoRpMvUs6z/85v4qU2q9/dSjeTHrx6IeiTZcAeHCb1xG67siJY4xUTPkzj
G447PRjK02gHmeQeFoijj+Fd2JgL6XSlkaStenAquOSWLpYnEBnYLS1CLydi
eTCvMHM7bcUMbmJWL7ldca3ASbpVBhi+RdKdkR4YKch+28NGNPDg9xwLmWZM
jPJxl6UYGoy7whJLc/flfD/rzAS9HlQ24IclNE64/Mxr0PFtfASGfFTLOfMa
nzwCQWOYsjqkY+V/w42tBLyZ7yeRtvXULQQ4+wiILLo2Vgp2lgzSqt/K6jzH
y4O97sROuonr+QZ/ajF2Noci936/MRqIQ4I6xT5m49FTGWZ7LUV0hca6aTmo
o8qFspa0X5J68VgVmUDlOcOxieCjHFsK/ocrGTCQM64eo1kNqauudBZmPtBP
UcDOhjBG5RhTP06Wp/4SYReI4tGR7Hb1UaOTvl5rrkN6dtQ7r71bhBg7QKsG
uq1Bf9lroyZYw68vO/g+mS0d6hnCbmGNgZSMCwd7DqdVwbt+024Agd9tQZhO
/YmBSPd7SB27Iz2AK44AAVgI44K0uoLoJQLh7iJ7ADgsBBmjLxPKMzGIowHJ
gNPRfSor9e8cWLcqmHfGRs7MdkdSce8avX4uUOFKBvp1IT69tCb/vMJtudcF
rS5lhn0ErmCJpx9zYDKTt/HFRDhgQL2AspoHZicwBhvjHl3v0SrDOq9+qlcj
jTsWegQCvAShGvYTqX5DrG/wiiHis0HudGkDHE6fCWFS8+8xwtFTukFtSYhI
EELXCJocxGIsBz6LhMYYGWCFAFAU4/UyvfcN0rkQN9eDT/2QpN5eAlaxVbj9
ST+VKaN0MGHnD0vG7GgzUlVLZV464H/XSrp2bPczQqtVYLuIMJqWXL54R/kQ
V2JbcoKT8bavzznnZEqfzPCulhH5AmUP1ko7gIROB/yGPWRBVSZ4PIgKqYaW
tf9O3C/Cj+p6lO3CvJ5Rpl/0P2Q1VjnHtr4QENwnsYbjeSJzO410/Es4/YKA
5zZfU2omZ6ZyCIGxd5MKfo4vUDfJ009rZ8IKMRv1aIBBTz1m+Us2Mx7Xhu4Y
G9QKAN2MW9mv2yeWXxyApXsTwlNR9UTIC7ftqXzqxRRkROW9mWQAJiBZecMl
vq7f4k7HLj9IML7ov75zBnLPygjRYd/ddP5ncCxb59COPec92EkS483ZL+rq
5FX6OnHIk98WsnphKgQstZ/ueYIcn2nDfiAXKH2OCHHcJRPVf5d4dwoR96hH
M1/RpjbA5RoLOtdxkAb+/aXoqpV2ypmX9z4x6eQ+nc1W58XM3794Grw66AGT
P4MbIspdnI3QG5cV1/7BFhFHxZTK+sZydtNGTfyeYe8pfSnZiC/sS1cfrgBM
BWdkpXAdDuphnmjS1QwJrrIiDu6F9ZGrhpuVBMvnGudRz+hEaWMO3Yaau7MO
WDG3MhYZdRLvGGwiC57YjjfFkHr/dyvsrBPs0fSF3w59awl+tDMsv37zuY4Z
TTWiCcREQ7xDdvWdjg8B6TJa3BJ1pUxkYvDqgDK80Z4sc9tnJPBgAQ8FkDcR
Tt4P6ZtyxXJ0DJY5SrEIT/es5NDsfxGF/KSkgHan80dcgzE28r8rwoseALoe
eaKFCDe8OTxeslduYanxBl7Ht7PQ5geIUMZKDWHTQNCbK7yVUp6YTz42N0Jx
77O7Q3UGqnyGIvf7Bgukfp4v0wD58WJx03BrM8RAt2QwfYeUfNp6jKC3phPQ
aRQ2s3nUly4DnWsp4z8rLvioZLmVCrnk7qeni8twOd1XuyZT81TdN0NA4Vfh
cRKpXyd8y9sW9Ktq7KwWyAYe15myvBHO/CN19P628H7jAJZWeSUue3x2p/WV
DWe9c2yN8zYbUGdcsB/qiTo2ldoDaKD60MLi4E8VzmCSg46P5PISJdi/cina
KmIAfysjqstcDu0u5pm5eqxUDC5VFrU+j0KrnaSgLdLygPTn2emp0tBC2Dig
li33PQCqukNNzNpj4ERFtaF4foCXDOyHkuWunVx3HhVLy4Z6AZCOTMuI+FXq
s9W9KPuk1Wugcwi6hGg7xcTNuvxQ18hnAHO3nBztecWBTE+4WSJU1okOeiSx
ReJg8ILRGyf8nCs+kZAFya2IKMKxYiey9uoTOKI1pkMHKpSqKQmWiNOPViDB
1+bzO+0PTSUcHtvs4FMfP2BNPbYmz5iXVyMRTYp7lNJxk3CbhcJ0eWUZYEPW
wn00iZqdKQgs2AzWufOnMcxuUQZkNkUFqz9ly1knH8rtEGzCUaUYB0gSAptP
87RQWxgCu8O2I4DTrAp644DJevbzuIWR6NZXrHpc/X6dvfM9u6bI4CB0P6/j
UpwmiNVth1WFJOauzWNy1C0lmSgpwtwj+RGxYNI9IBh3BqLgbPfS1pNFbsFX
hjuHeuooU1pMGurEf2ApBqhPMC43Xrt+dJvg/STnICeHt8IuKVNsVCw0hv9j
RTmdfqCCH52Rikdd74U4WCeSCK/JvmnaQvusSFEgVuc1/q3BPxB7XfsSGy4J
wdlNsls7CoMN6nwAY+4UcKs5gcalC4F8fV/eOcRDQhOQkaGgf1ZsknuRoIHZ
TqevdAUdnZcfCLMjykoGzZXaSl7r64FjPLkG9y3WVHvKivpo4+mr3C5xHNtu
ntooAQBMdiFg1X15xELsLs+gHGfoixFUGNABe7Z14HRgpe9jp9TON0+6zYIg
/ryd7MtgW6C2ALh4aeBTPfT3S49u4r7X0jGC/BbjI/rXbgN+J+6idwPwffm0
i0LaWQcoZ0myQ0UKQ6LyOonok9dTXyWN+vHbsEgmrjV38sAFKqfrf3SkkHcZ
bTe3GkPtPcB3Vmg3rU4L5KungDg/gczeVYCA3RSficX/cbdKaVDNtc9Ku9Vx
uDSMkTYgMAHHad+KtQe2kjHXHrNfdvc/6iXAaNPPEMMLorBzK72H4L4YTBkB
ZU8TJrajJCL9J0yKMPqnL+l+am2sr8eKjwLyDOhwLY4Y6WY4/nnim1kA/hMN
ifLH8jLfeJxEzeyNmyiTIAZFqdlUuQiG+thbmEup/v9Ln+jhtxqkq6NQ8aYo
JJllshb51IFNtErcGnrDLFUXRQYdrosXkB1JmJn8QkhqWuRX2iNMOM1yW7F8
xO2OmNLvdGByZRokkEhHCFbqlUhqRdIX6GErEQfWG3cjvL1KWEgW51PPTE4w
EjuXB4SPdh8InIhMcpXfI1xemHEklkO0xSNAcm9UV1nSmOVErU+RJZBFRNKC
MRvfHjdjonQCc02YZrz/An6zGQf8nI0iJYxbHhMXqueDfmVZBHYD0DXZQzWM
zniyBUgHi/yQ+CcbswvPLmeKt634QaX/Mhgg/kwObK3FiUEJKopIJkAaXvX5
vEH28xNt2i3bLdNMk6jXVi3wP2pzXOl4EyV1Uaz5YxIcPxmgajXa1YrsRZPw
5rJ67sO7vvBkm8X5fVeluyUWJqQk3r0jQXYzVSnJ/veaWptqcgLvDeJFfRow
dAv2kJsXpCFZrwdiI5MND6q5bodpFBrmMWlSFJHzKKrflLu21NGCYEjCbSjM
PuxPhiwqxZjIGfL7OjPWARqQvTEdxTjOYbwfBr7zj8yFC3w4GII7PeNjF4UN
oqmbB8dq8MNJ2wbwBfF1Dj0HLj9+II0m3+Pf+3c7SDT5xYPWjXyOLCqxSpKB
jvTY9u4vvkFTLbSTwAs9VvY/X7/PQIzvH93sSRHhy/q9BYdPQpY52fXdUYui
8lYkE5BWU+ZfPosi7NSVBe2kFymfViLwuk7Q8JgUSsXtUlVeujIZbsZbLXUg
qmfDtjO74RF55pqcn4wM97Tih7D24II9CZ7yqubmRteu5W3UxN5Az47B5ixz
L6J02hjkXL5L5XiRuVtMtw6BP7NWqLLcvOkuNP2O3EH8gSP3SrSflt0hGIaj
jSZMIqC6LOKGs31B8f1hJ3LTb8BK7tGy//tJxzkrUr47gLF9dqhmXHUdZkaR
UooZS6seNL5Ly2qdosWVth+jwvIWyVqtvNYSDRUmpMTfuL7oZkuSTTeRo1dN
E06jIuWnKTKw83+5QjianUYI0/IkEBKwrTA4Js6YFe5chAKUaUMZnQhVMmLo
4YhxBL6eNA86bVW9IpXpp3jdwB97H4ygHPaNHnkCThXIdrBi4Zyb845/uXh4
vgQDs8/H1rLLBSMLN+FE6aadjP/PpAYgPLA8RzOFN2BncjuyYM2cAMBEIIia
v7lhpzL+FIA7Ns7DOvUUMCEYiPrMbw1PgyAPRwr80ekl2REdFuvsO+R3imdj
gzKx933fc+ZU3L26sXtWAX39N+jjwUnV/fQPq8iCjYwDEnxLTyafLrAtaUhS
ZIxQ3ZNJ0aB2VVT6EN6aFBSz4YY/HPDy65K5ytoAu6BQBrwEX06UCKVmNpw2
7mBPXfM5tufTiMfekjJFYEXpF8v2YugKCr5smtAcylo6lNYzjjlAQJcgQKSH
C7UMWSNneLqdiqUy4xBbArpgppa0Gt8AdTjYz7Ox/EqYm/ygKqFy5EgKFmMm
1+JYamm2yAmh74k0Fx3HOsG+CCbNYFWgDKRyh720K1Vmb/7hVMC6J3MxwPuS
trh9SbmS0A+RzlptkTcjURGJ0EPOcoDQrPK353E2tzFcjTbMd2isCggwnCKm
RFgsYR1aSsFr2tisqqZfsDF7cBUKPx2RAF1tfz6MaaDuzkwH06phXXn1iVcg
pbKV/L5IEkfekDGDTtiRoAwp20q8Kq8tQpcJKuDX0uiuyMN3yKRE9+pCElC/
2Kl+EbSWaUQhXIhmQx6nmOoKYi2lESsl0kEBxlXBl7zZ7aEUwjvxTzE4O6Fi
EOkX6yfoJQvkUHBMDHEams63kAOZoiayd2hkaWEfDs9OXuqstIRgqP885aEu
Sk6EQKtFCupegnifMspPuPi5J4OAstjSXbSdBeJVhvurJgFsxNjAvv1Oy1JM
iAbXCibJtQ7frQK8vzjziJdsD5jFniyH8DIvwqykfDAt7qtqHYqouPr8e3FU
Bvxe/em5iP/SCk+zLM8NgKLqg6cK5eCc3ilbSXE1WIa8l+ntsODS1Cxp6vO+
4CLvQ2ekYEWtaKE4OzUMcPnZSgjB1+xM1o/Kbc8SRtkWGAk4INJuOs9bzrgk
6l8ogrdGtw4ruJ5IKwhDD7Ha8PPU5umAWONilYag+b5F94/trYTs8MtTKH4c
S9x7l5wTFeAB0nyR3sqy7PWkZY5kfWzVJu6Z4rJShvVFACXoFDFjwrTdJqkQ
xb3v9TXYAzWe/XPTWmlzrEBSKR4lp9Ho1ZyQ3lkVcbXmrxWZibI1YWoiY8Kb
fJA2Rp+tAky8KHZDUqHx44VIZjTBPbHewMw5RO4W8Mw+lmkr4eINpctm6RRh
TZd+HHrZlwfl5TWKBY4vUAOqBy237i+SS2kMeMj7NqSNm6JOqg6o3AZTxS/r
66iH3hoDgvawrrJLd4Lrw+1CYQiH5BUjzwo9GQv7riuiJ/1FCYJbcdLhj29+
3AS8VilHYI51YLZmpIYbyhq/EGUj+6Tfg0KX3YVrDuUXvGLLpJX+8q8rwBWy
23W8c5WGHHx8xamsqHCpHhI7J5u7I0WpTopihN6mwbwCViWSW6l1f6+Td2Uy
65InAJ/GWuaR1IoF8iYxBE2WFbcbkOtCQRuuw4HC8KiLtVzFMTGN0kjVjqvR
ArkM51ZHwyZ+WHf37RV/MPJeI86Z39M7iAyniTNNxGVSyHh1AfHaNsmIQUqS
Mgs4QYrOELj/DVTPGdUPORMZ7zUh0jPCY4NpQ8ZN7qBouaFvNZa5t3QFERrk
uuFn16vhFpzVO+ebeRQvvCq4i+5gv6aNSkhOipQCz1zlx6gDUK1vnK0n6oGw
ImDmhZEROW8vCOL8Qdo5o8wE9S2zkJj8LX3H5aVTfa7D65j+LG850ETqbR0+
iSYlyTFjljt2W1qkltRKHK8pHlFD2meaq0L8QjNudVmeA0TTDxv9XhtISwxL
yrrjZ67f75fdUsTnuyBeG5pwTSqQX141mylZJN+Vhwk9FAMsi4iByKFsnxbe
QR5V/PZ+75GGk+CCwC82WSUTEvVMZzupvT9C1n7kT/cS7j4zOBCH8wccNhgU
ej5pvqZHt1blOe29eCYjJssF4ARWVTZl2KY3NL1OuJScq6c38d8EuW1ffbtl
QXggD+8Vppe9PwAH5o91S59ejRzB3uAtA8/BPF6WoSgVBvipsvofb7S6Q4q8
E3Dln94ZHYYnCMq9ZgAAVIehFcNUw4JqK2KCgXX/ootj97JFxZ/P+70/r7AG
C3Zt0Wa2tGtkyZaZ6xwtklTkgT09pfvC96hCIEBkwXXQ2ylLWjDGkXUX8Ip9
TuT4b/1KCzob4IDh3LhCuPrDUqCxtX3rOoHwB0Xzw1MgcaeohKPymRgxcVtK
VOMqQAKfJZC6Pbn79rceKfve4nb6QKc2QW7vA9qNDCL7nm6ohG3RFYRlhzMQ
snxLUkhmVE4hoNBPCdhQcTWsY9rez7jjzgrexG3IgCs53dYlDW/Eh88OJrD4
YWPLUpLosHciiYB8ql4ukWbX001J+drlnwPURMh4INLk9x9o9ROfPTeJEWN/
9dliw3wiVBA8a4qAUIWQQTl80NntBVrtTSPA26fpyr63p9EMRpKCmlODKQji
xYSLlcoZ0E9NayFvWm/dU9d6xgAK3MiOy/IGTJty6SnzeZzi72y18DyLRJ7N
9zmOtyRyjrLDPaHGm02oyg8wPcnToQg/MoVej/WeckqPAbbZx0U+mR1wHgf8
pM/nWnP2xds7fyqwQSTHH2VgCUCDuBJRHEccHGSz740iBaiX/HzEEx37v4JA
Dyet73PnFUXbapXFUB3f6gsFmpbZbJkby+9rLPXli79MmtFgYocu3tuvl2l6
bt1/Mue7/i4HHfCciWPn3okc1Y9iImmlEeJRztGM8GslCAAvgnqplbCs9OPr
zSUTLwn424csqjlkH3Lt1wgZqPcRgWjcPrRZmQ5KzqaKVYdLPt/DCi9LHcKw
1XhvHMOV4Sz3rn3Bg1IE8Wq7pIyaRjtgXVnbfH3C0fCmhvQKkfOWewXLEi39
ynSPc6pGR7rZ/HncvTMhfVYNrVsOU+Y6gvjQ57mMdHTe2v5pIbjYdliNF9+0
HmeWLZGbLXultqX70/L1pXscICaR/NQ9rECg+CRehKGW1DXgmyvN4n27kd+f
WAZAOFTWGVk3TpI7gFlcXzc833Rn34ci+Zq2JIGaGtFt+ii2N0vL0mgunZ+n
zKxJ6ueCS0SD1J4jHeZ99h78F2PSwLUAW5iIHBqpOOa5wgxyeUMoIVF5VnC6
1QEOj7OthWVhKLWivVXq0rfdjodzfYnaDRHFiomemTYUrkuyWwZIinlK9u3m
FpsBB6eFPkglI04KA98SC9d9VbIHNbPot6HMBhdidwzD83aBYrqGyWrn1vnV
W7a/57Y08p4iPiB2vuhNeUeD6dySsSsPDDcWtNUojooHEC4vI0sMUIWAV6bO
LW/pg6XtLH9VQO9DqXhyW2l+RqHgxclEkuKZfczCL5HVR4sVA9TzlTHZ0isO
2xElAKpr1QVYb2JfpLEN8VigoBHWv3KLY+Gr4lKenX1GXKa1PGTqoBFfTGzV
CZWieFufT+Fe7gWUUpN152gDCrlpeXnchBHJ+ACno39Lkmlk2vvy9cLmaUEm
rSFXM76dTfIGoTHMYL41qBK0+DaeX1ijvhqs7KPgW1Vjd/yn5idyBAQ2/gCs
ElZsPvb2ZfARFZwahyrLzuqrW7MroMjpzdUmVDExH4NBcvUP62wDqRgI6wqq
9GN8u75vS8bpC8TRpp+7OREny9A0d25891dHSDwl/eL5fk9rnybjZTzAYUeD
6kP1lqymik1tNJ/gETabvY5jAHq6ksBxQCDiz+HT9549O2ZWTMxWEi2onLBv
fC97Sg1QW1GQb2sLo/aAMSWGpa/Z4Y8xd3dzA42XSKoPMZDIBAOdqScXBQxp
yx+5INKXvB/37HfZSaxeaOXyNmnZnW+QByMdN6Ve/0eR4DpS06XegUmAHeOZ
8O1zBeWzv59v6sx2RDKwLOZE3Uyxc8StttRVHShOfl2g9cdXH/3qy02YDDpv
3XqpllNiDvE2I0wNLH/t2AVSMfHzZPzR5medM37ICvKJNve0VvNFVVc13xd+
IBXXH5ZY6AreiqWTBnD7CZccCHpBvlaTHX6Q4QI59uvynk6CXDkylg2jEbaX
bW2AlyomTcf6OrnH4FT7umdwFwcqLbjQTxlKphjSgX0mAuCjAki4wbBV27OA
xtiMUh8RWqbN5bRj+VoPGSbMrU7cR79twONx+cz24VzgpxFl6vKi7bhHcSzP
Tqnciv+5hE+1eit3+usYm8up1CRV7MwV4bLGd+NVSksJGJzO2zQ0B1/fvpno
yf4IsaP6SrYpHz/i2KrclduuNLv0ltVkRQJud50mqvngHqnt8CcQiAYfSvrd
lf3C95pLZeBp78QTtcrSHXvC4JctWexr5n0fBy2cyCo5hiJfebpbcPrHMUBK
sFFxWfxOfCn1NFZXTO9N/xN1KLMjTQ9otIfSwWuLGuNOY8AgiTKo9lenZNzI
qD1pY/l266F1vshM1HN7xbHzCQ4in3EgANXEHy7DZyagFwbpmnMHUJX9XsRO
ydRS3fCLVrcEZGyrXRSSqj5s0pjc53s07b4APmaRjrWNDfGMVn8LYrSQiUL3
f8gWSQhkXCHHbdXdqGGKzcV+Mljrsepzqteoa4UWRHONo5iF4pGWCiV/xlt0
5P367VRYF1lMajwrBk+Ynm3xY/YeZxc+cpjcBKtV3fJ6TTU1CDCpkZlPrSAk
lfrUMQACDsXIfWFk1s9Ppgx1T1FskYGgjanPrSioORnLuvSo96Tcr2Y8XRfi
sEjgzVGaBD64ImqWa8apCey+R/LC4ETU+Uzvmm7RJ/1AkY9890R/LyGh91aV
tXrhySZ+iCslMvl9R89BD/jmzSFj97bByjcv8uUqfJlRpeY4phZnNO1rMWNv
MiJsT6bXJGorADCjA4fiqltYOexeZmT06axfqqS+LgLVOyYHusK3RHO4ZF4o
eiFcvquzOf0v2ZDCDKWZhM1APGomUYY3/YRgZ4sbh4kiQC2hguyIAaStCE8E
2G3qkw3+DQ6KnSfo2u/cU/0ndVb1tIrGWoKTpllT0QwtNey0DpyVPdBCJcN9
PRKx3nFf45ufOgYme68zq1tRxqqvUf/s9ngPGUrnmFY3Te2S9kBMT7k3lkwm
Bi20ntlLYpBsZ+atOhdcwyrB00XsOr+fqUitxiEvyYZqu75HecjU/FgssKCw
QVJ4oKOn8ylPvjuWtBUwH6o1O094qOTgds667FdOy0WQ8SYVByvFuL5k3tV0
xrRr6RwIVB2Kr5Qq9dYyOF8bHUsubtD+E9WVrGHLbv6U82QGufZaNLiEoCGD
2fd6NQTGh2JYBT5VNvk00w3kC1SyOowxg0eJFX0W4B6iyc4DrYoFUDyZy3YF
hzHTnUd7z5Nq2ms2/dCyPpUeViH16fqSfUWA5h4CyP1WdpaFaZVF/qo+p8LF
1MI/4naA7co89T0giNejjI8aP7HlvZu/qzclkAiBuvOawFXHzYDgh2aVPZLd
JOfcJ38aJMUi+zW34G1IBdaQ6U2p+V7IlPRBDsHUk4XNhdRBJE857EQailkG
cDKqrNJVltFV9cy93A+2e3/M7aqtqof6olyo9wapDw/Buk66mpwdawmBPTM2
4nXTQsccib042t23i+kn0P+GaS3XhL4wFP7NHvSWQv7l+X6R9mY6MubiYTj2
DnoE/+Zvb1AvI6DRCAgzK/oeWRXHNpEOnOIe1Cbn0tX4HFmZd7lGWvrl1SfS
mfbSkXf9Xzkd+bxUft15olljiCOsxXqNDLkpp9ybqS9aILzBuX8YEszxPGwd
YNoYFw2z3aOsveTgiWcGN5Z+NYi4ozgzXX3UjgyKqurNCvk/BqoPHopC9qtR
gk2svYosuxAIRRebhe3fjMiwngsTQdb+aiLiwEMVGKqMXWn8SsbDuPBzbjmv
sJ6UrDKu1fnP0S/A6BpM0H9rfIEkMXbtDSgyq+OZpuIX7AUdqz7a/ECWrD1Y
PenzsTBaQ31wfxijBph6K0iG3sH4GDBpMpm37Debu2BEm0L0RS729THHjxj2
FE7jU+VY3YL7VqNLJvslsa/sNM4GcGYfdpaF3RJ5hXzq9sZw5qG3s0Ub9Yy8
LCGIFHi5175CBs9TSLjgHW89sDR6n/tcm6Aznl+UvLm49kbFniEi02Wlw/3y
8ARiW4hVC8bjLMt1COkUhHQYiFK3ha0E8hd+iie0ZrmMH0mZBeeft2CROi49
vfGRd25XoWmnErS091W1PUzWLn9XQhfDMTWY+4xYaTsh9i3sDTw8LEBDUPN5
SFNthQKFItaJBuMNOkWm3bbY3ju+qwe26vhGCBn7V2lsSZmuY6+OuK9g70iK
FhfQdLn3YGZDy5MsZEVupoOJ6zRaIAmDkRFSpZGNekEo9JUouXJ7oWksPkQv
E3CvtqTV0rpD4UwQwft/WIg5fqOVyKYeLlVmYA+HhuTMf7h6tgH8yvzq0ze2
J8k7xe+dxXvHnxaeJOCPA0LKfOnavLSb1k+XLhpWcWQsVQS6U++CAhVJIWED
AWGOeEixXXV3wVMQYwjMx2I2u8AoGqirrgkjN35MVh5XXkbPOfP3Tm1WKMb0
ANYlBYPOkgQmmSwuDUB39MDOs5lZy/nUmricxljOxxV4na2ibZAk3RblXTHZ
JJs7i8klo680FzK202qIHz7iCJI+C7VKs1i/wG1eWDZw4Jg6FZ/RsEt05lHX
SP9nl8azCF6hZGmCy8dJgMS8Q576UZ5e0uj5uRkNd1WUBI/9RYCRNkkpup8U
UHf/lI/ujxmU8Xn8mBKaD9E4y+c0f0vEA2liztLrEtWQaWzqfO+It0FoFNQ8
F8+mWYyWiKJDrulGhdogbtvHQxVWYDoch65o4dzteuqGTzfKpd7Zl25yJW9x
bv0sydapi5UxkJI4qtE9wnmM71AtOj0ZLYLCDS8og/o43TIysNvwvzgjfNmU
+Ns4Lhwro3xQEylX/woI4PvoA7cP/xRYPqkgT9mgPD7UvjsKv3szBt9SryMb
+v/7pZOJnD7JGHB8MuQuRayAkj18qNSwM4O+sCCWI6Fh/bGI+jW6ddAQrxJF
yiPv6k2nseEcRMWPATPAe6NwyeRn4awfk+IJJ2uaXdM+UdEqkXFhbASQwgFE
sKiwg4Ts4Gi52KhssbCF8FR4uHr0DvOCh+v2acUcXtY44wKAebBO0gZJPFb4
RinRdl9hU0CO04RV6AjXmPfS393M0ackYBBkkjC7dsLY4Uh1eRlc2W9BWd83
qBMrFpFNwQy6T/mtQxaLnmisIMcyd6AotN7HcpK25sasLSf4QPFCGuZq53jM
udfNaANe8wzXiu0vgalF6bh+BPn7dZDXA0a/e3XUUvXBr6BFHR5TJaoqPTuw
bqlNJBdwwXwG7Zu/rtgGDqgFsRmi4+yTaSChElm+d0wP4Cb19bFNT9B4+t7L
lHiXu92yRqTWu8bsjRls+iqwonWyhAWp+mU3f0Lt/0xxR4YTPLIXef45lrLX
ZlrJjbDQBzT1+Ez5CkG+N/ZANqEYhYiQMBz4xt7Zs/Hl4A143tIQqAttwoCo
Di4CAGbniN0hWirfUeSOHV75lcpu4yp7ZpyzyoaGd6TdbO/WS56Tik9c3L//
LLAZZ+xOtfs2YNz20aWJ+Cz+IkkCfUlSRg03UhFdmayUwvT5lAlP9UShNR90
zA4rdVX/tV82BmFNhSS2PoNohpgTXP8vuAdQBT0fY4O8bIn0Th1HhsVzyqGE
M6wb/jIrXrVnNK4oaUrrPNwCULNWwY3kv60zBypMzf2i3o0n8FsNhBGnBI8E
nW7PmdGDE6SolK6eZAySosu2kJvxpVzGYvOrN3/hze3aa1Wl7e+37iQNGYyN
9vnxL4S/5sT3MSMARY2a8E950qnCvoviUthdjm+ofDOigOWDlaarmpzP5qi0
3lsphS8A2hSv+aSHpV7vXdjiScRfpMw+3u34AmVSodHwGsW6KGYYrpArA3W+
zayfgfdEOCzA+LJ6Ezky+PmaJzuoR0pKVvhobKfGyuNmnf7pjKwY77sfqh/4
wPbQBSVOAGcRqa1XjpzPyvwO4mBLwyotCP5y77s/uX58ACvYKyresebuqFuH
g+dm8GLDXdc4nXKB6PVYOcihYRIZfMlty+HFriS3WmRcs6SaB8AUfdZ5s+z2
xGegajcRxs0r7ElUi+wHGajMQEX6v8h6z8dGbUgXK89HySzspNxra1RS8SKz
3LEITSlCJP4yzx9myzsib0oXVrfptf4RABYPeiOHqgU5tgI/kkf6f+VC1fz/
zEYlRNVx1g7W35r7xJ5YuGZPBFITyOB5WGXCYnDvZ7+Zz9LP4gy1B4MHjasX
IXiubZ0VrHLqT/91DZrDODHWCw4EP3z2ka/y24/l1XKUesR+LhUYw+7QHxMS
GDT0nRa1GlApj6eHbYUchRVbJYjy641zeqd36ZTK96zrRClkrQ6UNfdHHLhi
Ik5p5Z7AAmOwdjC2iCxXIN4Jp0AhZX1vSJDAaxTZf2+5TFuyEWyisoWfYdzG
DLiRFqg8h8+WWyEHi/1pA7B1CurCDtda9GQjctuQu5zpWVnnFipSLaB87A1z
YoSWMVDLtPbuYe0Yh40yLv9ASPe5DcCBQ3caB/9AZu1VJDBjwDVqDxB4TeTc
W+dIREj/r8mNBMN2jONeWfdCSm7e9PlTzKPNMTTw0bZxfDI2HaudRMh847Jc
2DHvqNmF8206qWW73XpRP86TPP96T+TSTNyVKnSnzNyNb/9rnmxH8h5fxf0f
Gs1Qnvl0FoVG9MlPb1ci4DaCkmOMqz73JW94XAOsDCupXCxyv28YsTzmg2KS
AjUp0+zCwKipACnO/J/MBZ2ThDExtFRWFaFcRi8B0A0KN2RxVMKe8uqmoA6t
RhwCWgz+vbMajvBwU/d+MlBlTLmFCMSAaIHRj1/PGP89oG5ZkQLKHE0i9Uh+
O/16VpLatf4lm5oYl1GtVe1LMRGJ25/jMAKE1yCtR0f1xsyUfJXakfV5m6gL
4OqJP6KnrL42hYL5Nqmj9+SFz7dGrirmBNiEiY971ooa8wJb6xLiJmnd+mwv
Ev+F3FXDFK2UhI3ulH6XfEVGWtslEqo9da2FvcIv28VVuwZLuOB0f05FDxRV
v0UlW2ToJjEQ/DZ1Zq3rBA9JSwdGpiFhqif9HbX/CZaXVEuwlLwXpDVgVg9o
+v/27depkYSo5H66zQrjv1IqWMthZqQPVnxKSLzmRrw+aTWqt+o7kMPqF5I9
9C2kxpDBa7NrYCLA+4twuzbe7Im3B7SzOyXKRfN/Z+NVOFofDab6sEPusMx3
CuYeaLE7KdutiG8RNUTkXpTKhEOvgirMgBxGPKCN3mMQCnWe6V0YQUfae4kY
NYX2OGDv8/o6SLQg6mfxJcjvm0sy2blAWof394UTioeb0qTEDWmwbie4jy7d
1EfPabiRrTAvE8pik7eROhqRJWuorJrQVSCTubc8/c0Dq0r3kMpZl6TKBfWC
ooJUYgxXFBENRp1p+blh4LY+UaXGKCk6FYEu9wCl0IJTuZFAhZCltJLPdsZz
WSW/uJIrSFVMrWjUukNk+dbDOXp3XxpgI3WPLmTvX8GoJ4JEoOb3QUFAaNy/
gsHEAevAL+k1NkJ5gkPZIZSfctYK74itY/p7rCKt2R9VJ7XDyuO7C2b+u7h6
7yyDrhGVsmKuaXg2lD8OEf/8jj3iGWLjF70w1LDUJky69t21kwIUaFPR8mnu
BBN9U/UPgcqxlEk+Sfnv4F2KI2JlrYRknRNdkDYJgTM+gEPUCOTWFc9ciXi0
uCRx/Kp8sPYCo34nLBnORqRLLSJ5PfYf7wnK1O7pwWX0Sao3y3Q4mcY5YjaL
LiGKqcH0qCCy85MU8Hd8AQQk5HwCQAkOM1K+JSKPkL2UoW9rbVZpskSVhcMq
siNyyQXZ8jdirP+vPJeK5idnZbPzxNVHdV2hFnK993SGz+YSjafpZqWT0gdJ
FMjlgZHAZ3F5vljh0YGk/Z3cbksmAI7tWv1c9G4X4P/KJgMUQEvnkron0qxA
m906+FrHgyqYbqua8kgMoYK7KRoc1BeqWROHfYYAUj8WfmJdESEU8MIQIW61
PwVpOkFrZi9rdzI1NVIuZ1rtK7ly/ImWo+wfF/4ds7ajrsoT7B6ZFEwilyNF
ha8HuJxEa2VZZXme01UhTpBoY57SI1Nw5ZJw9+UJyV/ww1er7ka6yJSOBd0l
Juy6DVexsfgKXH480oUIE3zlAKjwnkcwyCzgWxuuloFs3jFn1IABqSqnxDhr
UXHB0CWKZaww/vJw2m9JgVmcW6mI0tEHb6KInFQh8xtR/PGaF+sdCtDcYA6p
1k4/Gp8TyJZzroQ5Wutdh84EpaTNXlT9xb1w88gEiWOMJ05yAJTUHYS+lT3W
hBao+RkHjBs/qXxs52mTBRwIfxIVsWLFbUt9BRtloI7QXHByZUemXXYuX9hM
CFul+XAnfC0QRvdCUZJ5hQ7MDCQ1LuM2C4KmsBpbGWHg3HY4o+EqngS0UqmB
JBT8JjeanM0DtWMkRDtl94dy9US6b0yYmTtWj+IhTmQx/7JaZIZiYwtF5qrf
4oreJX0eEmPS3nrFqLN53w2qdfXQM10FSJ/vUF81HAyDrxt88QKWRteTofLF
F3uB+mQD36LiPfWwOO6w1pZldF19p52BGgFqXL5w61u7ui4ahsVLyUGIadiq
xplGvq6DTGrHbIwYasElvUKHBwiZ6WKzYJIpG6UHy+H4uadYAjuWfuPQg1Jg
Yydq8++NPEwDYC04gFXFGr/dHazcPxTNkF2rmZIKJJxdYDGbMR6zQw0oPQKr
mmh4tan9/TzSO82M2HgP71AhrmifPkEJ4me8JESQsnl407Uyjpwj8XU1q5nK
V9GOn627tM8kYKd/j4sVs7oFpP+ti+IhQzHCJBQgj5IkfXDj9SZOu+Mwqg1d
wF6t8clqgu5vEQ5a5QGeFA9spwOL0YCWMRzEXK3CHEQPhIs3Wb7KgruYYrWV
i5qkbQ1lIDw7FMGXw/+sUDwuRT7WOzMO5kBbSLiXDPW1N2iDOineZ/brZsK9
fngCSPViCcFvgT76j7ew1BCp8NLwzpnNZDKBCztGNP31k1P1ypK/tbG8lpfI
zEbiksMrQHHKlMHuqWjzhDif2FDCrkVvVfKw/qp6x3cDMCKWjilSuIMTtzAF
mdM2NYI3x8uqkHFR8Hitet5LKBC4shNrStNx8eHlS8hTNJW/CSV+QqXZ8cz8
zwQlGpWBUEaIB85Tdgs0LObQ74PtrXlI6xo8iTBcTTwgUwbJbIkYX8ZVtTfy
ZLNeUv6LNIS0BL1rR2dvdvz1bXPxyZj2O0nFOzTIovKa99M9FtkfVpyd1A9V
cwGSPZ3JVM7XAwWnWccl2BOKpGctvkjuOveXO1Fh0L2+76eM8cnb1EtyMVc9
UUTHTwdiTWS4I/rpxqIUuyk1BWtREnW0QimmRPLaGZEG4sqkCx1ohJZTi2B5
KiGaeA207/T0SgDG/HYznnjuqWo7f2pbc8e/K0tzZJt5zEqJpEAGEnz0a+zQ
+tIOsrJLalre6B9RTPJYq8Wspt7Q6r/suOkvzPcFu3VbYz04+J90LBSRikZG
a7fOzs6qyupliDQEM65kyWpLmgcdzMu0ApmxLhb80hCDFxHbmI5chaAyjTOI
Jv1xs28GM3ldOxsnP52ydBzb7/s3Y/hojYcGd2hYdpSh2eGCVsBBQLjXvh6B
aN4kz5B0PVenvLUdR1UaHvfwj9zCLLUz2OW3SiirBFZ91DDfPsDcq+a0ajKX
Ya5ygMIXsG75gvYviw0iPdPwpnGMqNF+QSutFll9FD1ykDdiaTAfZNOGjyAJ
09izDtdhDV7FBKEfzi+B0hezEtYKROuGu5jY3PEd1qDTqbtmfF+r5/ZozIUe
EBG9to383oxY9oBItvZodyKunz8QjB8HEbh6OYbX8bhDCYjkXNwj6mec4mYN
uKd+JCqSfdKYFgg6ph4LUL3vsGhEAjSh/V8TZK5zV2//wSKU3kowtRfuPwx3
iqDmV7HgeWasyvNiLvJ36FcJ0l1yjKpJrTmMIVSunDiJw04yyOqMAcyKx+6r
Rdvc8pAoRMc8QyOtA1OBSszA+H9ljdnyCkeQ/LWpxd6rFhbdbFb+Q96MyU7/
BAxEUofk/GDLbj5/QM4x7li5aINL3fGIoqKt4TBZKEH+gnrAofDapj/wNbwl
K8J9aYzQpAlz8nkJ5ncCIG+kK8osdGC4lo7F1k1qJBdYlTVt6Ci5ySQS7n0A
0MRyFmGdfu2atyN0mpeDjFuvO8SWjNNn/ubXLjkIqKpDtPf4CXNVPgeqLf9E
2LVcc12ct6lRxLXiamzVwsd2ESH3LBtvmokrKV1xNXQBoGTEMRVUz7TgWAh6
yys57KabATFKubVUPlUEh49OFirbvEucWId7X1dCOv7gvI/mOXAX6wDDMbdK
rbIj6tzlXQQLCLWJ7den7sdRGUdG1GKrcwJ8ngqOO2CTUa1HFngWYw6sx3u5
dteJIBwJKYtdGl5eVQ2nWRGY16d8jcZTuzDvMpcOw7tXpoZRyh6YYiBwgQN/
J63hlw7gFP7s8RUqmyyLyehNfBaQBg5LLMKBvKe+C9DK+0Yr+j9hL4OFMu0m
qdlw0+fNj8UATZpw1oNhFRwCqh6CoQbGjBtlgkXgfRX8cPnoFXzeFYjdFrxu
ut5d+vAJFjrVuEmoQOSF4F2yQN7tAZEGcFSuO3Q0v0+eO6Hryy2Ech8sM7jI
InGyPuyp+sEWURaiB/CRpE3946kzPPUt8xR9vTTx5vsFIHE/CZaAtvriL/Qt
rS3u5M4WN5rhR6zsWnM8/dXv9z5D8JzmYIq2yX+x9scEMJePraCxmA4ZgCG5
CmzTSOGMwm34SXR+qZEEoJoFaJ9Q/V8gIlTLzNqX9vfwf1+1a9N8YiDxgGYm
MD4hDgaYXGY+8NlIx49KMzvpNoJ3xJoozYP0qY2aj6sK5OXEwyo5IK0Ifb29
M5SSZUqMrm+L+TRXri70ky8kEKOT7IziyInQ2hAR+jjUIJwFTnDm5pBz0KsB
ZW3E5FZbLu5CH4LuXcUonEJ2k47Gjo2yM5jvTnWJOTxJFx5OSekYUeisIBZ/
3jZNT0QXy0h3esgy4OzppJPniMpCRsOp0i3HWpckaUxgPW75k3pFVbBAuVJ2
Wiagop4O4u2tMRUA77kcPlSMaGzyzTpr+ApjqyTLJGAN7DQ8IYNhYWxQB6E3
J5dFwjzfVKoEBpva4kbCBlrB4lpj+aoGna+NsLFNGEyz+6iODr7IDsBAeCEO
hMly7qro/1BZGEEenaytXgcgER9QcrVQaTiSLPGGKQ98iYqGc/omLAXp4SvD
ehEIIhnPO0ygaG7bbg/eOdybr2zJKYtY5dxuYnggoQgQmUiA9Qs72HeHol51
HxZ5eAjoLmlEthSVqP5+J1XXS84YKJc/9zv/MFwe2OAoaXWi+CcWYwuh4QFQ
VDMuoOXIG7w4I/qLcQozlsKjnIFSZ1G6b3apJlV7LkODPhVeVhZXkLy3p/j4
CXxtwnDPVYOalq0VcQiToVHvObnb9SD1y2hi6+yMkrPIuRi/Gnp+wC4Gc50L
VpygZ1VooGazvRVT9Xpw9GqD7/0YMNEFK3446NRDSTYE7wUaugTber+HwQ+m
2eFAxEqna1sJOG0Q/5EVTPEy2w5n/HEXIFaQMxyI7SO7Ma0m/gZycR3dbYl5
gztB77fTg1OhEb6wSTXT8gFKexULP5wUMKRd4T8tFchrJ2bswy9tvOx+TRDo
hGmYjb9DFZyyYAqYidjaeBOHPM7edSoWG0H9QkQdijPMHEbR5KWaCVtyVGAZ
e3DUPCv3UXzuBkjqvkxYowt4RyaV4EXsq9FYTWBVsUzixuA6o4FyN1479IUI
XEEXzT1d3yAYTPCXVmd71b/JAq9VWXD7fOLJwbhGTsn5R1tyq/glo466KMax
DthNbRbKx/BaD/IybMdUUMqGssD0BpKMCpw8znwEwefxwGibrsxQupEmL2F/
7xHnbyIS5Ec1FTlOmoL/3+48cllHMd1zVtUxBsqa+Gv47tgqCS0ByS3DoQdw
r/Cq2sDmP9hlrgBB9Ahkw59HgAXLtbAz5/6QfFqIENyLyUgFG/rUHIMfdWcz
0tAQcap1kx9a3koKwM+yRJzcu7neI00xoAGUVBe/A9Ob/mF+SPKARpdMfG5V
GkcntY5330GlUTJyQdzuMlBkSJK0Z0hoHZNYNkkYgeQKDKZm+LMJ+l8wfk22
WASSs2BO2o9FnlLEZ446oiT0cGPqG3U2xhBElhmBj+0gruVs4TA3V/WPK2sD
1j7oMZSy5RJck5hnMzwsPbyFvMwXZfW61evem9Bg/poBDEp8Z5nFAxEzomfM
KuJJoZN4qLr0EoFILwmGwvLhqge4gIqMzFiJI/DcTvsBK4/nDhze80wddBnG
Fv1p0htjdmmH6pvOKld9Pcvd0uZjQm3EjI3aYsYbcQisFwlGPglNo4TmJclJ
waODGXN4D020wSs45cEpRkQpYDCYMuWmv38EfAzW8Dl8zCad/VX66A52yS8R
KwGWJz4WFZhD/Qss4mEDR1E6l2s/R7FvTEfckOyn5KuAzEoGMegKXekbf7nh
JYaEkWHCI/Q8OzQNRGtefaN43oACUM5ezzM5tnRKWGLe0cj99xCX6tprqfWk
K1KUcYCSkEp8J00NbmHoW6nMnvyu4lA07FNCM0sOkII//X5tabtSJ+rqH4n3
XIgzJi9cSxqobUOJiwjs28bxTmPq1HSChU/RtcT6ea/KALdkt1Aaq06dRPRK
Advj20HGFJa6bI9nB9xT8ez7f0pNCpixlXBl1HQO9zs3TrL8iOcssiwlyMnU
f2pyjYhN5mDriihQ02HzCldDmK38EV9Sik0gvEu2/HDjDw/hsMkK4UMHUS5C
JqdV072ALrvF/B0KUSPXfgEEedZDf9whzKs6l/d+tVlB5WKWi+/xbgJtosAm
8sEPwY+R7khot7rssh9xGEvUY9Yo3PV3q17ETfUQJl32E5Lg7BxFNbAEf1Bh
xaob4p9sL9yajTnNYibu+JD5f8LEwom5OgFJUN8ooCVp9YhyN9y94ZP5RLMv
in5IhIbIa4lpBXKTe/1mVNDAsZMK+jMheuAyNy3oo0kfi346zhu5Onv/xTMy
26Qy60R2HLgEouH/TDZrbXlK3eySESviXe+cQJ6+5hNyRW5DRrKGvbu/Q/uC
AvLkd8WpRsBPjIFnMteHIw4iNtusk4b9Rdb6mn+4+Jn7MfoVwMM0J3NYAbN/
0mOOuoElONPE+WsnftUgoFrGzZMGpfuP9MYOKhAzCle3tex116cT88zOTChg
nr0dstT7IOg74mY9FTZHdQsTUnbm7x6VJZ8bhu40lZx18ozy4ejF8mrpMl2C
pBQHV6oX0PS4BPDu9OV9/nUVPbOHSCPzn+25sB37fjeG8IRsZaUAyBxlZZ2T
8hQmfXtfZcnw+hgrF+NuXnBLd7H78Gf6EwqVZmKYCr3jzWnQf0eN+F9tUc3W
pzn7Vt6dslw2BNjgGOYGF4vGVMEzXZLEm5DueW7a3AWzbD6Dom8SCjw4hj4I
8PuosP0zyatMzygrKMQvOWeLtMBPR2v2a+QcaqFujS2p1Iya5J9W2bcqNZ4n
835SKzbqRAaxIr6VxVblT1AjJHsEKK0IAXUEW2dMSKABpNxUy0FKltqjHzm8
HGpH5hFwbo4ehW1MW6HypGNZ91TYWkfQdcDphCrSd2+Ac7U3g/HbkkpAzwyb
IdnQTLoRaA+yQfyZCbxy5Jf4CHl1mATTU41kee+XP6bIvBIHNRrzV5rXS2N8
8E+XsOf8JbpKnCJNDNYM+eQSdZD55KQhJViO/P99DmvxWUGj58XrMXxcjwvw
hlp2tP0Q7EwKyU/qUgIUxhVHVrWUSG3T0krwdSW2Fq6AdorrAiCidldvbxvU
bQ8s3QV55sSyiC09se16O6O8GN1BqhyDizrT+413tNh4hZlXFj3VNpp5abFi
q1hyJp+f9INkQYgxEc2dAwuKzkTP3zJsv0URRqU0CNvsFDxsMhhoo4opnpOB
XNgoRRATs0wuorlpuBDcOUb0eDRss5h+V71rLEfbnVUC43PBniF6e3nW4ZEH
wAdQA847zVrS4hio5TifzaW2JpnpmGB8AH6EMnEalNhJSD/9Pt1DTr7pVEpv
iiQCAxfp/ZlEnpnQFLWoR4C4Rw5tiEri7SicWmqI+G4I1voRhE5MPWrhvsR9
lmVJzUOGVqyxd5vjr6eSsM0ZnRUecPaZy2dU3QcN1+vTs3YNJVqiOysNOGUo
+saPQBncN/+iCBOHz9yvKbcWgfqMCKRSmfMkevfI7Cf7CE8RAFer5hslIcgx
eJ5DaYej0Sv4HhhYbltlnSNh/6iLdjUIJOG+ch1Dep4Jlfy0W5412arw8Lpk
zm1aY38MQTghqyni9FIBrYF0arG8av1H5B/3C1QvSnf5LmQQaNUdDcz6Haew
D9WqYR/05Cz0SWIgLZOqvR2ga3PIhQKcXl+J33yCJoZI1IRY9YckBGOsX/JC
2jUDkXsYt0PhBx5tXU3atZhp4XavEkzjkQdjQDtj2hm3r8/xRCEiQiEFF8zF
iiggGaZf+B32YjzW7G5gim33QiVSWsqatMQ1CKLvp9LPgms4D96nYnmxaeMm
QdELRZ+vlnTbOognpX/kXWhoa7hl1v7lQFCFqLkh7WCc3FrXiiPy1NCttQ1L
QxrFPsu8CEqIkdIQnrsDTJRBZZ3uZbwGAgB0/l4OQCK842z07akV5giTGXoZ
T69MrN9br8l4zG80GJ2Ocb9NMopQDcef8444Kj8Mcq3k7Io9JSH/TpD6gCtp
H4sLEMJC+dQ+nmYlyDcMZk79kHLN+IgCkCaUOgj+PEEKvlNN5cV3bopqUQfd
PJsUd7+oU8iwTUEEHyg8kV2tLRFYmaK9M1Ibs/DCR/KO9p/sgE80LeuDOHc/
Z7nIXPhvfKEETNLSDt84diOWXkAqjX95EAIiCPNDV9PxpeFf2G4Mw+o84Ebe
uF+Mly/VUAfP8L4LRRJRKCCm1+XEECAee1MBO/dbtJIWqt5iHfTpo3v3kPKK
pMeq1MZPmRzqkH82RBeIyQPcngAUbN27NVqoKrFWBIMyEHnTZIVaD+H5hAkP
dZJ0QvggvRl297xb3qU1aly/z7FMQ+Emu1pRDDTujITWm99xRxDcUWga9JT1
NwXLwrbc/lTFO/35bLqVOixeyIu3V6a+5Vf9x7VRQBEaz77stMYoeolomoPR
44PkSOwmdmysSdOTFhpcXESYaXPkHCDx2A7WevOntyKgYP4sIdu1T1ChvohA
FSHQjP0qMs3uf/CKclLBdg/pDZulJWl5pF4riGmtAYs5nHP2t0Ws077hwmDH
7xai8IdgKYESppVV/oSz1aBCKbmwpJ8H3C7wX0jK9AyOk/f8y5K7fEU5nCdV
Pc8Q9DMnXlkeQBfUFzYVWss5xrypuXk8iZVWkuuMphNXJKChTgQ402wa8fRx
L1YPKElk9+tWSTBo76Yfwl6zfDr2SlylYlo+V/xiiHM01TUGTPnyK2b8FQIE
7cQAJFuzP6KFSr2j+JIBV/PN+Ao5ISdppbscW495M27jtVkOUOBdmYoHuAsj
03AP2dyHyrdu7ApYHXLYchqIf9LpRrwpwclAmIScmw0XC2OogIEl3LcaA633
WS+5zZqYiU9xTt79eBMta5F1TamgtWHK3y2lw0AcDpEBwRYXqGL4m4+qdb2/
jiq6G1KhCSbSpL1EMbao+st8UBpT05iTS8Xrv6dSSAWiyosadbhOemnha0Jk
3/vYwqivXR7XLXOOqZzd/dQKrgGlkA3JtxS3x5lkNDNquXthe/sAo06jdONt
jyxlkcr4WeBUx2Rkf3t7sIAEfEa8F8J6CAHod5wjeebH7/y6ycMa6wm0qAAU
5w8EGuvNFXmAbhXHWmXrVCiJO4OGnReCmtE/Mwa7P3m9sXzQngjYdXofrWNw
TqYTQisGDIRpQxoXvlRUrCAoe6OJ4C0v5bj6G+E05HzbYS7H8kTDMyAdZi8p
GJ1WdaQy/3faiyZMAUlJ1s+GiICp8k7nbdGF1mH0skCrRtrE50iTfnrmvnWg
yJv25wwLaHcr3b9O/6edK/Nzrqvb3UBisu9foSJ5yxXJWTHdDM+Gi6ijmlI1
F3MfMGBkiwxP5cmbQza4RzJONuoyomx2ciFv9NHlPV8iJgLy7c+6+xa6ncwy
fWBGR+nr2X4UWSakJC8ma3SdzfMRyGYygQBwdOzHn2HdtuA69NKH8Dmup5DU
JCfnRKCP9HydfpUiD6XUW8s9d++v9BorNJMyQc8y+PVQhfYcVou23sfvtosE
2ztk+Eskt/B4O9MRbMsuru3cllHxvmBGPmJcLy4m9q9pCvHGED76KnrGaHBQ
+LGXyWYPzcq36jvkYRBQc5aqMCYDoGmArim3kVNdYJnbj0jPjuxV7j70NtHP
1yRNn+ChnMZJEFU4hTn4CjiYu8iV6Y48LBcjDJrl2sspc4xpImFBbOJpbyTG
Njhs8VVambHap4Wh0FjS6mWLgTkZZVnL3pX9K+Z8V51LvmLGXnk8HF85hPE6
vy7RR6MWlNr+jCjKs8AXulHKoHfymyzegflkd59pYg7p8ZXKxN4OLJqzhk03
4nb0WWmPgWCT7qEKDUUC+uQZTqV/LYoy4xoar6EFKayK0/F2cZcWOdafGvSn
oMo2Wq9IPKkmqubF8qOIYTcqMKA9wIALNJ2gnKiSefsjSyNRlGNkJUvF7J6k
+6A7eHQJJc6PdBZVWCfDGYUjsBkfk5ZhGvWR7G0vclVD4YOYE9BjJtrJLd1v
v3dbs5p1eGvK6a9re17FSjAHK+3egPSUuhrMiFZOAQt+csCIz9Gx6BzG4l5a
fTaqJw4gzCG4o9rg24mirlUP8qTW11UguDFiHyi/KkbGJ7cU3L0e8yYbKbdu
N6w/SJh4IFdHiKHJSLp6Gl8uudmlELK0GGvxiMZk7+VIELzgTCSCOdfVxG0w
nSTuTnBnAcJ5dtZnjyAbjx3T6KAhf1G05NoKrldhENEqpni14eZuVE7LHBOY
nl3UKGpm/yvzuwRDjjtjnqwEQVZo1nyEcwyiofTt0X80Fdz2WKwilV724mba
luPtwy7nW598s+M+Fq/Dd7TI5EErRfaFaOizL91aPOnwgR7YeJVlpqj+xzjJ
Mh0AcWXq3cwzRiT0i/F4s9/7wbQo9E33OyGZIKEStllVqBzh1tV0KjarbQSE
q2xFKcQBEtAMz0p4zTWOlyZLYuOmSjPYxHDSW1k2+Caps+4R9ujjEluRF1GE
pcldCugLOeYgj0A8TwEI+UGQpIxMKhr9P8iATstgS3DpY+GHNliFCIqeo/4U
5DCVYxZGSCxWFJafrU3Zc2S3muhxd/0drwIooOCHVEmfeDVMgxeFFCUoxPou
5L85JNjmPe27UZ3AaL04v4n/oP+JQ6BqjcIFjt73XPqjh8Jfz2hYnLc5ft1q
Vi1a5VhTCcveEFY+RuQfAaQgMpE6oMxIX9DAa+IMf240QLxZsJWKoXGfQ6w3
tDQc3Ys2FaZW67yyb8j8+9rTuGkQdzc8r7QVHk9WR9t4w0zjUGSiSdt25ooS
ujZXlYFRhQQ41ShFKzrpAZLnuQGDrXe6h+lj+WMM6a2pKGRpmW0X0RDc0Axw
lzOSWcurF7HcjASfhn6jP9l5WqGXMyOWf441ee66OYoiKA8JcR2PtJ0xbCVG
oJ3Euivnc64c9dMS9fFrE4UrfolYvAVeZW1UlGYu1wFSLIcD1wFiWrnox4JM
LLB+PD87YEU7yxHh+d08e3s/H4JeZ9k6MTeKADhPJ/Y8+5LC334R2OZtjfXW
h5J6mbw0r2KHgnMyCT6F1TDxVYNKeXGij1Vqo7sqMXnKU9pFUamNO0SrPkFk
WGTUtNIuYu9kqQAv62+ajAeB5bWRcuAWwrOvVIXR1cLoWKc8UglUWeVKxvaH
Z4rJUYjNre/yeuVXk50vgCO1rqNaXxzoobAJhSvwEHWux8wFey2fPZ1LNFmn
pOtWbaZwFcLmTQIyG3HHIVe2lcntJTgivYNjJgWVUHuNvmQRYiwCDOV5ZnbM
gcX5sezliJ4DFOFGX+0iHsq6e+b0MOG6tk5RSYN+IAC5G1q5SABG2uMs3yjK
VRHzJWq43438ngszF6WBi0Qr62zwq4FZKqaUh9G/5d5L68MDD9VFbLGFPMyH
Gyv10mhzPBzMervrLH1+BRSiLW37xNjClphKdgYC5Y61JZySQ9x9nOFB6DHx
wr53CMHFkRvYoZyt+Rmx+oCMnQeod1fkRsBKznAScYu/rm7KI0r/x0ZqdFDG
YVXq3FcBiSdWcOcM1fgRHJ9GnlTLUyMoBxbBaLEEME2JWDeQYD6yL1Bf7O+a
6ZeF28Jy4ibDgBHP9FRrfoH40DjgoYu/VS5oe6P6ina46Uo+ms+l4cZLa0GP
iD6kBf0tHL7Ya/0MP1VJeW4AHPJ0bLC9dZlMchBoPk6RAtp65xU7Po0OKvCK
heHxklCfni5z5LBfzfexWFbPV6dWGM02HQC/fgiyebIQKOEmDU9glbPLfrSS
kXzyX2Zz5yrEu5yrjWSApXU+6/zPYcjxwVEueOmQSfcMlBP0VzUgjtJDyQHH
9diYutwJ18oXrVOHqCNGk7ti+cTaj31QgL95wW5W/HdsHjfR0L9PoioxMcy/
dZBVGteF0bi9RVAu5qy8VBbxtA7WbZ+UaxYHMPqn1JYNWJrQnbJmKMIiUuR1
TxQaV3CdbzQBHPMSAAT6/isV1bw8OYsIwnrNY7aoozadf+W/esVSybqY3WQP
3v5seVwGI3yv9M1RjziXWnWgFO/2QbCXQD6uYYf/127Bjz26GR1eT77fYO4U
stXcCX6ooHXWscg5UwdmxAe4uWsHdV3p2I0MSK116uzvXHpwahg8dM1B5BOg
JIqeEAEhGbZDoKk1hHI3nGCPZ4aBd5hWOTuqfJngd7ck7cCXKYq+26tVxIQk
vewAqxK7fV6eaK+P6UHgXhuBRYmQPNHWLOsxOhxWzCVgFUUFQby4yRXZjljj
bRAClHDlCY8d7sRAAs0qB2blbBAc5yGETCJwvPiW1iGEKxqSei+E0xU16UUW
1w+NQgTGPKOohovPKg+/BCjpA6lu+xf1k4Iuy9Isjcc346vD4GTYYUkJ1JW0
xdnVe2jTMN2v3QTix2Un5Ag+zJb6bcA2LK7crtiCR659/ELbYJri5/5I/B/M
cALiaStJimLslImWmssNi+xOj96KJt+nsSRJALx0fkQZefQz7OqandmyQqXo
XcYmpLvyvYjYT6jsXMpqLJpiHrQgSILYNQ1doG1xBnhFkxIbWmFgqb6Y7TbR
7pOXaIZ6Jv9HODdi/jSbQqQZuoD9gDru2Tu5oEnDC0D0GYgDroHbMK2nWk5Z
l2LqaFPdP5fpXS2HLFz9XuTgmLJ5vaBMw0vEVK4WuI8uouHwVwC6+8XPnfPF
9LWlu6sBdHXArOzZWV56n4zUyqVK2Ntj1EnTIqfVzZ10UdY96QhuXHn+QAig
PhGaNBpmCXF8npU1HZ3CspUZ8BLV6WteoQax4Bh8FpjXAFG3knLvACw10KVi
Xl+kKWYKJDRBp3eSA5QGcJmEVkJj7bzuRUhd1JF8FsnWzGaOIosx0Ky3rUjD
oH7zFWVBgOl2aora8sEuBfkzYiHCfR0g3IwwKlho1zZ1/4t82QTzD8RkUa/E
McY7BG9A0+4bTgutI88EgdVHPhDRj3i9uiCWbFdoc9kZte4sMq3dDsOwiPr7
wE516ex1LFvCXLRkGlsIxc9CqX1C4CdipqoDkYcRTIgNKZn/DWHKGeeTwiaH
ATBLr8b8jrT5AojvlfRw2OyFr4bButz3h3h0meyDwBLMKOZdcEyuZEErq/Z5
VNZunsBnpj2MmHLFb8d6cT+B7sh20gu9+IzEglsV5+HNR5ciIDrSQof+eQPi
FqyUVcDn9r0QiAWIBIQ0zxlnmkgbP56Ji8KOCHJBA4UMXpkaQuRFM/L9xQL8
FQZqF5gnjDdwplo1c23F3M+JJT6VDNn+kZZcTXJdpsm+5yqx6eEdwAmE4TCV
v1TlpGhnfk1cICopk99jf4L/YwbUH8qu/+dJzuNq9MsfHrC5B6zChi+e24+h
0Ti06OWkm4P2Ekbke2wHh7W3cMmxTotGsZYkdWgOobv/3DdLK/0AkEc5r7hd
Ust3DCwFmsvNIn4oGrOF4aT9cBgkfqX7KmaEs03OleNckqyopzGBDicF1WQj
36hDh7q0BQulmow0RbS4z69QQsUiRzpXZVpPFZLXdh4IC14+MYZEtWLV7N2E
OJwZA7oLHMbKrJxBzIgfVh+rBOsv8gMeUy3T9a7XcnZUrRr68du6k2x/YsHJ
ShSjTy/lZejtubFcrEdmEegreX7uf+J770LgEL2VSrwmcTgJjc/2Gp/yaPGE
W3JmSP7q3HuC8xCWeKgQt3AbwKoyefu7cBTJYsjH2nNM75RL3Uto/jPK1N+P
9Zr9iP1qaoyNTaSEJzACHxJVo+EHiD1kk12CJTgkaNssFxSlWbMY9xsVV8bQ
CjUiv7853ac8tTuH1E8ixD3jc2PZOzUhjzD8p7oOI+EF5fCuHotVnHrHFCSv
+fDvbeGsUogInTtXVWpVrgzq3M6B3ZS683o5x9le2ioNX8dxsI8q1dQDsaDr
Wyy0/2ugwlYwvBz/qCoBm9zpzlN7gpQcSIgWTJ4cWYnT2Vl0shzI3mHaIfpl
GCL5jsS58id3cveNQRj3Vy12aavL0wOsOXWeow5HYwA/7WQ7o28XR7c9VDM7
gcFGbQaZcD4Hr92U0Q2WrOsoUOaIxErEBzVNkEaygqcUUtJPx5Ea1xpWsnR0
QS0GfG9QNiETNmZshvIFQxBmDRlDzbRFKtvvS9uTkK9d37UBUaOw7eh38/w2
uC9XIbGprzcQV/XYRcLNqIoY0J348b2dBsmYNoibQp5QqW+bAYuMd64RGnwt
e3PqnxJS3UD6z82rri2B9e/INuQXpCcwWVjzTthdrOwHsqKamvkXiyJ1/K2i
rCpjDkg0M9EexbUCGW8JYNmYBHXHNodzL0EjAri7c+0y46euQTrC6KxeNt2t
vSqDGbgsK2eaonjXKV+fiiFRFuEmGqS3QpyFZQlzR3IcsPhnuaWJi2v7DP7Y
h7L+ynNukJJj67/Vu98WHhS6WD86HJaCKLOT1Q7t7TpXYMY4RFnrviXnJ8pt
Tx5QyZvGyPAG0aj5ioJvbmQAmJMP/Hj9sg7QDWRtBmPX8WEx9lrMZ2wKZf9X
TWKzIIXJypO65S2TenbwZBpAymbDr0WWynrXQvJ0zjyDwJ7StGNQ8NVbIJn/
wVoHXrHHcBcKTUPJ75NR8jOzs/AF28TmSFDclr+kPWsudxd/NZH+5GlYnQTL
NBV0vrXWvuWNsOMnl48LXFg0805U5Tuj0hrnaD9M7c5WH0a2L8lxJx/XUydc
f/r2cnb5v3JuOuwWEwFMX3QW0nEve/1oSus+/lyLU8T9E4+1H36E94qTLsiO
y+sh0PEfQ63hICSfJDxx0M9g6QquzrBW0fKM/X7jWnL5b40Acjbm3nQKlYMH
HHWJjtrUthZo8lKFKRrq7/NiZikBlgcrpPk5uijjh9flpqrbVrmOISK5NszS
lvRXXB4KWxNZ5HSRn5dV9ofmOXOKmYRbzIHgQhuj/p3HDy9Hy4U/X7lqNTf4
STUshOwMoE8H2/ODbCsXsFsPA3SzwcpeJqqNwfkbLXVyJFYx/PAoBaJM3O5E
EM7vtpMivbWy5bDSN7qUj07MKmYdbfCPI7BhfodmaphYBU3/4eRh1FCk0ZQU
bFzQpnQtlDlJ0Vq5Ef4wwtdPDVGhCL+JJO5EHOzdsCk6zSLBuc8v8V7FV+YK
MFbG+KIKzYomiwhQC6sr8YHgepk4YHAPhNhmPfjTvW1+MAokZ6mlD2WoRswL
2WPS9vwoFdXDl35GDzCOXle9ZIesjBNf32+8scK4CxftVzf238chWG0imhw5
02to9mlGTvXltCoGE/bsD27e5fvIFNNg5EvJNoTouBGHD7Ln7E6+dedPhHcx
FL/HrkX7LOz+jN+6uyXGYOUd8E0/Q4A85g4WOjgmnprPAzo+COwH2IPbUG6J
tuL3OCGLNNxg5D5PMYrImuJKNB1qrW98NKeDSXql7Xovkry5ZVSGxbDN75gB
zh3NroSFShsI5BSH17BvRNKH72Ibj8McTwpLDLaVhGpmN8IWCYocou6yGpeP
QZ0QPAnVK2ehEIrLH31VBmr298GfwpjviQpjTW0+qNaLfg5BXklq2Q6N/TjT
TnsfSsfqcqaNfmX2vv3NJWBd1fcsFq7Wta8C72fAljBUZ8q/QG+d7v5sBkpV
Yh+11CwGQZzz6FlWuP8Rat5nDteUw/AH/F91T3SnxnzGKd7TiRcongYZecc8
BWiaWH6qz9v42gXw3VaGOfSPfihHYvD7tDdXcZ6YVdsHC3ikF98gnQsZhUu/
ZC4J3a3HrYeyh1R0UFSNPCjg4CB74oMeSwGTxsVwQmyd7Pxc8fFa4yH74lFJ
DdQaO/FpuBPZfIEhNCcaDdjh8/ie2yhB6N2AK8h4hLYas/wUznqPGxpY0oT3
YTK24D4NpvuYnc6BxwUHFVlJZHGowLUmRGW0JSVVkr7i4O3I/qetnkSE1BKm
s2UBN0aioW5Lhto2siz2piEIb2F0fg+Pka/+W42b39w7N0q+1EQndzQ0NV/T
2K3V6mvnTp2xuREOWkou5St83cItFoiXyyZ313XZ7GrDOukxUSHVyzzQmUS+
7r292dAmRVZJIwBXZRcdRUP+7rA6ewwC32uGRtjEhL7/TFlGPUavpLJUbttM
1GEG0QUkbthKXyp3cFw6RrukLdK0pc/JtYV+PQzj0aaG6AzzoOWbKI18IjT2
PlTn82rKeDxMW0AH/cpqrDAcckfpjR0ivNr3V2pu524wlydmR9Qk3DTxpmpt
quSr2nKDa5OxPHmpnkqo3NmJrFHVBu6fW95DnW/lG4CBBGqY3+sPg2+fJX73
mgMi+Wg0McJ5714fmp7fegs6Td3si+j9Q4lUWlDVNUAH1lSxWFcT1jWJggFm
NsEWvwHEmwhQXM7s9aNgXycn1e7VUDgxpPyKk5KAgWKT9zz9dwqvJvwg4dFt
C6RbmdFr65U2Z8jSUBtw07KVloKg4hpzAzT6EB5pMEWu3hdwVqiapwMiDaf0
bCsitPhpribBGUWL+Csapg+fUb8Mo/Zi75QvxC74kC3xl8qzs4GojnhEpegT
nE4aOfm8iC2q+jxZ1tGbjyw523VIuquZfsAu55gfhLgyAygvvxKD6fyezjp+
GmSDr+D7K5i4a/GDJ0/S30d7Za4NmSAInWGVCbZB28RyYaQGWbcBP/joYqMf
CIB/rPte600l4dKacqh8ulwKtiN5Cy0OrBw/Vfbvjj7JpXXL/6ZOK8SXlzpO
fBg7YmqQgqBMvoxZes/v+SF+4yx5lxsF8BqpOpKkfNXjE2MpjiNrZZe8HL7u
C5KYDbvAh8L0hAy7Kj3E9hbOR6JOLlBmIZC0HAAkAcwvg7R42zeHuMR8cPkt
MNQyWivPZZ4sD/kXPr+M/gRmJk52Glt72II1jrlLw6ctGi4agstIxhgJa/II
xZp4C+WRrnKAOXcohhvfBijBiOvqYfveuwtGim4lHAs9YWUxIYOI13lMxgQK
FkQmat5bOML7OgWt9hgjvhsxi3cYaxB7+IbOuwXBmPHfsen9kIpEpfohpbnQ
J9aGsJOnynkVkf5Um/LUwW3GJ4Y6L6m8XFIsZBqkT2iqzt2AHncf2tm1p0Cy
yrIiw6CJUt1/dpnapVDxw1l2LsDaEyUdz5fuXx0/mGQ+dDIyW6uBXd1ya1gh
SWFpTj7urK3y/DxSn31eKS0Bp559UZIxthQpRO7z/ZqtF1S4pTOHY2rDJ4qF
1omtuy5uCPgNy56JpEOBF9MaqajqKdmz8UDdHEEzojiARa6dHTjQgqrL8oCb
Nnl1HnxSwAa6zxZH7YpOG9t0it2Q+/HCQbum57ePze2abY+7g463y07ZOjPB
M19rnh7F7m2/zjEHQUjUDpKo0/+67TbQAr7eefE/HNCYU0BjR/D/vKShxeFC
9xFsgPvi0A4qke6Fwm6ra9Ta1qt13N+Y91e5KbCXSf/cjeY9tZMs2rViX/Mx
22CWgT+coNlF+laPJDlSN476kM/+Y0zTFoluLFH7fxfD6hPF0LUvk+5yB1qY
G5lUphfGXXQiUE6v+EUBe5JtPgigGjOr7lm9lnxryhG+Ddhpn2KVYEC4mfKp
KhhrxAjahEOavkGIsldnEqVwGTiZ1mtdkH6S3TREgqsU2E8PGOtW1R7x42u0
5LpRot0N/eVORZBJWlZhNiWrr6F9yvZbJphonbpHsQhGw2N/b7Onar0lmWr/
PLLK6ek2wzbyVuaOohcHV6QkLcg7kp8QfWMX6Jv4yFgv5FHgOK3CIkgILWg5
meSoS46F6sbJui0aa114TBPJbloBUdRi1cmCcMuCbxJIUd/YTDUMASOkupLm
4V15GJHeeKKkg2HITin4yrQ2Jk8QVEfyCTvmyz6bbr74omfn/pNZUv655Bdm
LT933oX92ZdVxXQG0ZnZDTRKL5XiFRg4QGYDklTMEYL9B+ZzeyOe1EI48tjs
zhy2XWvHD3oMArVmw8yf3kGyrItvo8txmPmA3E+msYtV4ZmzvBGAw8wo3PbV
rwh8yqraXJD6lYqSUrjY8jbOimzbhO2HcVUX/dLSApOzCZYbNGpGQ7OJImwg
UlMncbZsTb8sppH7mTONWcU/dTefXrSwIovhVBUJgDvLgNFK5GDLwJZHVvqW
fC6sHWUk5JZnTjsK7wt+yHPdA9oaWCVMG601PRIdxmSYY4QRflOo87jy4dVM
CBTLYU1OS3zfTStNAgNO0AE4i0cnmcTELtEr1uQ4WNv22DePQvqcfdoVZj0c
E/XjNAf/ZysvW84rlfpsj6wZyx4SOikeFbU9nEAfD0cVKEiNs6ESgAFoNWg1
1EvQOBStGjV8B1iom10lMRad70rHsySDkxewEtqWEya1O7qdeAZdwf3nLagE
ee941du7+EshkW2yuVBpKbfJdhPHatwAwngIobFzVKXLzLKYPp/QEDC426VP
tuTY9MOuebIxiCsXembq/OPz8nl93OZw8ZrdBLgrRZZ6ISKdJ9l7EWmqJ+CS
SWdOJ7wR6wjuiqAxlytTK20Qwifk3moqHJM1R4o9ARXwxXuE3K9Q0VdIj0v5
f6Wotc0MDZ2Upj5Uq7nYLtc6NyKsAQUj2dxi2VpCrDPkU4/9CkTiwZI4mSX5
dltt+OIMgG6gcBAsUkUTshq8b6F0YzkU1sb3e4UnuGvVyoL31UVLUrZwKUzi
uA7qL/vxMvdiX1njuxWymBcEE4Odp0p7anP4c0BmWdYlHDlL61gDaSMcQfv5
9lZa2Zk1Vx2kmyciN9pcruyXF0f0i+hMhHM+sJSXg3ajPDlUOFG2iytWa/7R
E6zzK36HKoo4Audl5/Eob0qkq7NB+l00gAgTLDGjZ2TjPuYp5Pzsq+HAUOeM
e9c3+my8UKkRjP2lslWWYGC06lLaZzbIvxZkNKVrzBAjeymsL1aNcM+sForN
MRKmM6PDWqRJKwCfrTa4XBb47ZwIbKZtVW+P6fW9cfs8Hdqdg4lAJtrxRBba
E3MCX/2RjEf/VmcR7OdlOiXcrm3xlRcteJ61WV7n+Tnv50koSH6vnXDQVgoI
B71rjjwRCzz1IpS0lWFJnBl68H9B8Oyu9agy0TgZn1pbidLVfk4IxqQ5NjAn
AmnHDmAjFRPzpFZnERpz5GT+m12FGmLw4lVAOTiZOgtiVSb6tQjomeVVhVE3
u7tX8DyZYoevqbTx+7LuClcu3lA7317F0NlK50bQux0HMI6KarOT73I/V2rY
GC3PD2lM9xtB0beCEslzMoQbqeXz4xaadLDOBkBk19h+pNGnMQFZhK5aQqpd
xyfvUHsBqVo5aH7UrV3cMZFxEc7EXxoyvSoYsKsIV93WjHzxj+EH+3PodFlh
bbUvDiJnRsqKiVuXGCCWCluL7HrQCQbWHSHrWTkgHVBAp8I7SP/nBKE2oTLy
RqQKeyQHgHxe2Nl53hymI2e2BFSEx2exVfeAvixqQzQt0I8dqe/5J9/Wu8D4
r0eMSIYqflcYG1Kv2IZXKNKO0Rr/7lcgA3YMV5bKaqmFHuSphijZKExXh0Hk
FuWAXxXxlxEdXZhDyu8ib7iFxe4oE3WMu3zelXwWuIlvVV0Fm4mS1mctNV0K
nW+mv5qAA3ABc+Dd66B+WdEDl7Ol1DTVQAN1HbR1bm/O9wwYRo3z/3e2O3OA
NFHM3z+EQuRLxyS6R/qdniW8RBQzUVZj+04xRYEX4oAdJMJOkUTpd1eaI1Bf
jrIWsUevwfANqVLqNHEFjWWoNC8NdAaoQ23hZbY5yLnZc+jl34zpPjC4RxOY
mWR339ZVcbhUKndedRTif8d5xU+39GQjzluOLDEbvZYVHfrhN1m5STTSbpNI
U6WYNQZaLhWg2YwG8PW7H3a/D6ymldNl7Z4wuF0kxK5cjqFR/1Uk8xipA3aZ
OPAjFswUm51BOc7UppAnqyxOzEoopPtcPbWsIbF6tCggYnqsYUwA22Au5sms
+V5VFGAvp/ZUZXBRzyzD4DoXf+PJS/UN9BDsLxPoTPw/hz8ObC8DR8lg0IA4
0ceVvjli2EeZWnsvaJJRSiJy5Qbr78n1dn5KMcfI/d5CQN/WrrfZhHDYPqp/
H2OKIAVqiDJHiinG/m3UKPVivQ2PsJ7ca9lZM1oqncGPAw0Ia3JGnshKNzfj
D9u5qzj50Oyb37ScMAz5tDpa4Vy72LBFONDy28cht3tpKzddFKjBpqiWthgm
/tg3v5XjzQhveUyfkJmsgJS4M7JtoeZp1o4PND0rlMRio5FzE+jvge+uNt5A
DwzR/7Dd5caKY82cjv9voy/zd6fI/qmzCLTRxLu0GOdRR4Ougf5j5iAZBCX4
EAe1UoQIRIIDJLpSXRyA/TKX2lPACcOZMXyD70QPmo3ovMqp3pLyyDxRgsPQ
Vrp8Sglwyz8WbARkz6+rtdeLNBl/aPcU0omYGMZuYlcDMKCrfLO2L9BpAXIT
htLA8XJ25aTSVWbNtNkCSY9QWi9QLIyikYOpBPWGGvponZy43YrEmrV9bgci
OgJ6FIOx5vW9jyt6fsEnf9C0ijrtjoLsW/+65Gm+XPzGJP5uIPstyO32eGtE
ZT4msl9+FvyR7Vvzz6UgshZc8oHZg7ld0/YBv3GZzZZHXdhF+YdC6DQ47duc
CIkBK6TqTKgLzP8f+UMULbnLo3vvId6w1Ddg4BYoxTCDGq951eaHF2+BWwd2
dLe+RGbInYAmwQuTnI8PBr+3C4aPW845c+TWI6//lM4XnOZ/2GqX/BZJ6OAv
rBWm9Ad8Zw0zgVVs2uUnZUhdyZyHilFwZv3em9GabPLtayTlsAW+Ud/iIiOu
QHFIrI0LcQPRn52rd/dQQLPQlQKK0fvo8LKETVbBKv+k4a3wMabiuidfWsm8
sLrPcdOTCqGg3E+nnETqjiVDC4+trA73ebGs0Lw+1Egxul4bnjfftKxDUErn
9KaLnG/N4mf4HcmhTYum/X276Y0uWe/vKg6WGdAw/W4BU8EqR74tdJ/q/xTk
HBByUxfDlubp9pZC0tmEITZrJ33hMY5N0gW1rd4dSKt5JOa/m/4w7cWK0hF6
F8Sb2HAMbipU7juEUmazniADGROKX6Qj88FXppxpH9OPpIKLaBvDh7w5C25r
2V/3vUUsLQraOaRby0+91u3/UWewXLTg6KAckwfH17nzQLzPxCN6q0pDMyUg
T09YIZlDsERlHhtBy/AANDj8V79mduWPbuS06lpUfgJd96hM1nHZcdOMpc4L
4fYeVoEieIpiagmlrfLFJtyV6FJWsLyPpt7nsahvgQrMnnGHrHqDkIWTIP1p
L9ItjCwHpmQSNny/Y0hip4ZN8Eb8C5fxXfliBJyhJmYBHR6ko54QVGPLXUCR
zRUlRfaslmSPuirfvorq72tNqQmjGo0wybvdAnS11xgpirDxrClj18V7l56r
ji9VLKTiOh4sI/9hYlvu/B9jcwa++djoXIeTkb08QUxwlzMk0hYHIQ0t3pw+
JlWw2UXsmjGGJ8xffcQkN6/yezXSKu3bMIuZ/jkMQZHREIKneYJ0untTILWr
zAptYoi7EbaVT8xqIblLF4XJ7nnosaGdDqweOM4Enbm48w9eeqfZATUUyUK5
2nxJlzG773/wPd3SLCrCdnepRhOhkWYCR845ALQeWRt5YPagGV8EniSNRx7H
Tk9DH7r5OiYunAGPdECVoPMEJjW9/+geU4UnKHZViPsloaj6Rr3TF7ZZnFB5
sB5pM084pD8deavjnxfwb2BwOqxVJ9R+/o8GHV3JhgnXIa/JxE85fg8rHlOX
h7rpZH6Pu+S4nk/hZnLzjynC5/LtzfvY1Ygc1zUa+dvGkZdrQmlJolLNETwt
ma+9m6E2YHB4mZYn8g91Qb71Vq6rXWU+h1uocheqmvEqnZ/QI1wdAczLSjNo
S3Y1cGYGOT3RevtQVq9Kb+1LLSMRLqB6aN8wTcQjSGUnUEUotY7NtL5nlBIU
I6z14tlItCE6MNJmjZAbZLfvWsgKsZwLL7o6YgzQhEbKjH6zsE3CZ+CYPiGQ
arMUFQra0cm+MxBxaRs6iVIMNWloyrY2DCl05CgSqBlZ2yiT+3t06j8gas/G
iCzgl5SWqkjE+LSEo5iEzp7dqpaYZIsnMdEP/Xitn3kiDtZZWk5PPBlPtiUS
7+c145JJLDDbA3CQ7jHuLwc7UlkUFVgZv3c7AGa1Bfh1vh2Bln87e1FWyPoW
zBx2CF2YeySIWeNVb4lCuSbl/jq5N7yNszZ4GHCI2Uk2LGQRt+C7Uarh5KYx
vh7Zv3EpR4a7aEKFB7d4Mnb7dAqKaf8z5w/KENBXTpBJIyTXa3uibDsKx7d0
ohnt/WZqPaq0PC1aNJRdSR0iYKZ8HcaQ3fWhxaJqOh2c7oLHHyKtA0JMFpvp
/Ekn4HklhW5wV5/haryD65+nNo/GVYCl+yG0pduMVKq4usye9yIl6KUmDR/d
oGK+9oQ9gR69Kiv+zjTMrI1agllJSzr35Tvtq05h0zO7MtmbscwkGEt9H0ug
Uy80fI9rVtswzDsEqw3JREHMQczV5Az1mHfvfrh6Q7eUU5ReD3koMpY9zZxi
9CpbXFtZ6UkTLRQ2JQAde8DQhbyRbSHDfjCAeoYob7IUnvyDZxIuGTuiEaWR
vb/uK1a7A8KWeRwc3F+hBHMEICM1/bAiVnEicMsuinXAYmdozxK98tK1nJJ/
cUv0hc7+IWQiyTVutUD3zVHugSahcTbY+x1ZyXpwReTHNh2a0+hfA2WhaOlI
2V2JD4a/ukRv5Xw44AJHn+PQPhfqF3tJVtaGSo0mzds2cn65A2YS1Md2KGz+
MyC++iES2pnfbeT5PYb0V3lZGvdxUkx+hlCE9S1uKAUnenBx8NIAvph8q4Vj
oIpfqoZBkwymALtlbRpxoxRQekV6Iot7SCtcHGTrA/Pojp12OCijH37J00ft
9SrSHEDW8a270hSO6rLicDpi95Lqm9sFId8b+82W/+pFDi0xcSctPUunNkon
AOkmH9G86GCZEM+Vu1tKnRiASKFdlnQJy10uiEhoBYZ/rlBePX4Kz6AO+QzZ
qkIIpcohRcvk0V82n/Gc5zxBuKOWToiITjUrtjwDIfBX/CEBhMlqrgnAQRlP
33tph6gskW5l4UQMXtS2gu2lho5LFLmnJLSC8qwNpBQCuR/Okzb2P7P+EgtS
PKZZYAA0ZXs4XW2XPRHBSn5jE6EiMVanLRQc/mwxYDL6NIGHZUIKrtM6QgdG
YuVXK+5l50sO1lp/rYhYYqZ4ZJrfG38ZGGUd6xRuCvSlybw9lQW8AzLjEcTP
mcRzBNFiKb3sRUGhkxvQp5ksmQKPsmp8vXSxA1A4HpMZedTMt4+J2FBi4u3/
+WNmwGSWv9Wi1kv0sqOW2t6sIQZQvkM8LCN4m2jLQ6wkkBFMg0orU22kqYJc
/cgn9YDtBPO+7MWkb7zvXTuyJG8xpbbiumx4BcEXdteJKvCbnk+eA/H/pzVl
eJjKj9nb1dFWn0URTGzXY5VjBc2lL3Im0XIUAac5Rgs4OTAa80THavpBBITx
0NA8p/ZDIV5lzP1hqNzrGJdfsyDl1P42LNQR1MGmKqOOiyo50viK4UzjvJl0
REVSCAbEHSR5JkrYG+C3GM+StmwEuRBbEt2m3WWU56atvRqSnUQ9dl6qgoQp
CZSjLh87D2eixechHEYkgdtrPuAet8NwyB+ap/u3pN6X9eZOw1QA7jW9WE1d
rqPhgb0ZK5MXvLn8dIpk8jL4Kktjl5P++8bMWhcZEP04Hhk6pVqE06Il6o1A
bjqXXVcfaqDzYNOcrmryEysCBrXGWDs8yx3A2E5ZRjYExSxsB8ASobMGBowS
518KZ+N1oWy7B+WrjAhbp7EB8fT1DAvgiLRGxXVbqwfQvOlA+qqfufDpBrsY
5byMoOayJBOE2OdToXFgZ+9dcnxnSouSi6BOpWwcPZ0sb4miOeFM9LuOgajN
0C/QasrolGTLtLjJBZ9ozvPQQuMgSV+MaF/k03gtauOFd9rV3N7g95gPpZ3E
wkYtsmvYG9DiQsx9T+2m/r9C3EieCt3m1GimHyIXBUGHeCRU1rcynSkQD9rE
NfM4AOMFWiCemP4ARKfcVGRnyegyrGKG+7mYzUQqKxtYFawMB/trkF7SJJ+y
H1UPabERgAiDIn5cCRMYTi2TZYnCkpnDkbPxhxWuba+O1bK/5EBL2wtDqYLE
Tkg7tASfoA/BjeaeRf8WOYi3QJCARaEm8NWR273wi7kJCP81ec7N6Nhu2uvh
aYqrAJXqBSS/eDfZ4FwX+/f5F+i2/0fWpik0DnbRpx/2eScoPr5QYXVBFF2f
Muunhdf/5v+2u+aJ8EGn24cIng9vnkvVZJjKlBXbFJ3UW+lnSatV7zXl+/Jg
Zm6I2v9+Ee8EckHkTVdAWtvVa4LtVtHoMKyK/fg0uDoATbTIV3abISBjdCCS
zLIIJs9sWhk2vIVyVcp5m+pPeokgrlTgjtQjZQim0aUxxF11rE5qW3XQpXsC
vAqJsK/b34R2Z4o3Sb+itBpI6OHLmeZDOlKo4bthAhq6Q/qIA0aXgqXpPKEq
owchbPY5qe/OlVpV9r0TGtbmKocgD2LruQ0b5l9cUKi9sHvzlLis8Aq7NS3Y
SUeNOgbmSFFuQzCdCgImXdl+svDdfEYtMziZaXNqEWLCGZYr+U9tjZI7cvf4
C9WF9yHEgvQE8g6sYnFIhPJt5UiDjzk5POrnubRkquqjqu8QsUe5K1/Vxpfh
hll9hQyhortVL6m/Qaks/4Nw/A2pd/W/d2AbUWw/PKpJBaWV0Zkl2KhrQHqC
xumEN7csRphVRSSusl7U1ZXvJKSJktHNcfXZ1kzkYuxN9zDQm3pgEZof0xo8
ZnboGCb6wIQ8wjLBtodZME7zTjZK5y/GC0dsGbHmKH8ByFaOB18yLF9SJxg1
ne1KJWnG4yCg0ifsUr/mQ7GBKnAq5Nc2w1iU2E5q+OacQAAFL4u9P79LU1cf
hBF3l9K3pb1ePzTCQVGiPsgW61feNlHx/qQDBNBoQy/OFDGYggZz4jB9w14d
4S3zObarepIsQEwwZbHCmKfVbuEnedQeU9htbkGgmwPRRFVpruoTN0IlNCNS
iPL6PzhHFRkoCTOkwaFP0ZmjoXN6bk79tLTNkcDb27X38rTmKc+irHcdpruT
hjh5/zY+HT1rbgM696SlS2jMYVgbw75FP4797ThXkVrrWIBXj99zOoktwPb0
T5ZqpAJj+BS6NLiZIQ8SHLxyGQXlXTlxfwEoua3h7t1MGNmzr+hWeY3YqzA7
R7AH/hIRcWLwvTS+OzkNE2MppvNw4e7V+J+mquWS8+mS+NBeqYO6obH2rwp5
Kk3y+0mJox9YZ+/ll3vEwL8ok8h74Vo3b7YQhH0TqNLYP2rJuBj1nyqYo6jQ
2Odf8rzDlrZsm4bgyq+Q829/FK4LjqRANyfqdYDUA7Hfv9vE9HN0tepnTxvf
qKKGyPBPqqF+GNWh41e4cmi7+GwRTbyOuZ0rJrYI5hQtx0C57fAHe8Qvj+Gm
18swdo34Cn2/vSzUPaFRjKCuO/3cAse0o4eyskovJT8Qdjlily/CETWwEniW
i6HNUbNkOMW53VE+oGscvpjH6OLYcSfZck2o18JFMIf1UpYrGCHWifu5zIFy
tdjMCa8y1lTPNcr1mVg0Cr9we3hLzOGOIBBjCFyJf3KWaOTP+fWRJ37eZSfi
ZOQeQwtnftFgOo1fO1Ms20KZUG7FHlqzsfAx9V3g0FfUzWF0RSXvTKlnlIsf
sn9Hi7PTpaDwBYHGOg5KkI+dZWyEh2SB6RXD1Aff7xdsms3slQLuodKnTwC9
8VjCAVPzJcyjdQYso5KmQEfJAD9K7T4eZpZcnUnczs/X8Vk7jqnjUXjF0WWH
88xLMmgb43jHcuKUD/lDkwGUDfl/Ri37eEhd8bqSNkObwvLeB8oEdDFYm1Oy
nDT3b2SCckk18Cskjogz6u4WAp3qFwCwTdkRH14saEDMgtp0mMwBvaHC234e
biSI0M+yZWKm4JsasI8xKY+v3X83OYU8Jg0qqN3Y9G59/I2ZPC8hoASvgwiR
Jj9EwTZCf6GkIStGLvDrgv8qu94KMOdTvxu3VJ8k62gNbqWw2pumW9VOBkud
+4iPySU54obS5xJi1UgqHh1f29SXBbPuYQVVinNQUI9uaGoI7/I5pRheKzR3
T4BasOIJsMe3tadrUTtVxftGdHrH0R5j6lAiZ0KmTbHzh7DRIuW80VVgQKo5
O+0/M0Mv7mL+hvCLkxflmT0H/QS0IEnCyd752XDtN0rt8BwqvYCpMhPUumFS
JRcXz6zcC9KdVF8HdrcDjqJ4ZNm53QDD8tQhV0FVL3Tto6c15WxYvG4Z1M8N
Oinfj7v4YpcQM+k7pg2LDElss2wyEfJLLXD4RjIip24XHfLzZDHI2iRDbqVp
ZI55niX5lT8r+TVjgA9hJOCunEYwXg9ZnNyVIUYhPdE6VfIwKSr5tuvawQe9
5dYUY9SVFFmX9fZV2aBpsW745cp4wC+jJbJ376+i7jclnCZQCuJpaeWPxHNU
ZjKk1378fBB5BO2HxXE7Jdy1KuKed6+XlcHPjI8QE4sQxbaQGm1sxEPMpiLR
1xHKCcOFld45YAXip5vNuKB355Cm5PGgH3iKUeG3uB9FyRoDQkIwB1IZSw8i
5SfdFVZgXHzYAb3/BNC+gjr8UJawdNg632kYYuFjMOc7vJ6u1tBhe6/LQUrP
qPmouFP1e13zR5tiIHt46TThguEGm1FtgNqgTkyec2ciERGrVNxcPNppPjRX
Ns3IrkiwIL+4p+5pcm1IBXh7H2YtK/o57Q0sFJH/OnWIAeYKTC+vJ16iccmB
6o+GIuL5lz62nVN869x/OWMHQfEGdvf1PaSjttcYV6OTfB6skSAX5mCCpPl5
+riUIxofhnGcMdjFJMR8rRgcqgKnBykhKf3h+0OMvvbyUCRx0oresmtBCrDb
ZcHKktg3DOKx6+/wWH62sBONvLmnJGazn0oiflWZvRuaDCc3rtrxV8bVptjW
KPNXmoy9yuD4zCtgYhUDFe4BWTJ3ds7NWauGTw9kCTKQJcr3fA1gcovRf4/Q
VC7mTwP3DSZ+0HMyeu5ewCN+i3ml4DsI+8O38MlbLoWmd5/PBc5XivKveQkl
Ae+mB0opmiDwfipWw/4eNG6G5iqiKag7y5NXQrUsi8WpF14icl+5QcStvUUm
FBPKA3Yk8mddjK59SyejWhnw384NfLRZWdu3zwq8NIuXQh2uPA3+byfPh7oJ
UhBrtjvIEoC1u5vkFHUZpA50DvWWJVEMNFWYkT10voYTCqNQkC7DAmLEuQDF
XdSIIIt+VKNDF9uC2TAG/JgubmFpLUDHdlp239qlox+UX5tp/t1lT0OIjEZr
18zI41rTCfnXzQzQIHREZMSi8S8n+uqMdGgMEfBbVEvVl8oxVmFpfJCN4eP0
RkyTDTEFq1Z4Jal90jNprUn5MedS8xOMMFPvL3MJmVsu3RP4NGs3m+7WZLKN
V5l+G638KEYWgNmmVqN3PJdS84y99PeKpnML/JHPMSnDBgApSfHDLn59VQKJ
WFkL2xu01MSPlz2Uyjl6rKkW91c2mljGgczx5hoPutmrFyGvH7DMGzFAK5lV
iq+G61lcxATzKuraew5ymSVImN/v16x+KU80QwyLityt9Ht/2sm4heVQEn0M
OG6p+60peF/Oy5f8H3+O6FZJ9LQY0128hafhiUQNEANmsjdb+otiuUfpIutY
XSDIqbVGcatMsQgZoAiuFclA084uErZOff7cHZNaFR/zg0lkW4QsLAtD7lTb
VNzvt0bsjmpjwmTYNC+6XFbUC5+RZ4yWIDeGq8nr5qi8KEJFMwwkPVs44GLG
HNiX+U3aLMhco4/2ahjBDaCB8KJbtakPZB9oqI/RaMs4peIkNcTtSzYxT/Hh
+EZOrOYf38CDyZssyvpUdW+XPACx0VjGMQoV6tmotB2z3NX+wGDHrpCaqNPR
KhPLZ39YoM6Xe8IS37ElUNuyU008cgZ3W99WEOk+a2cEvZUrcgp9fDZqOAL4
TZa7pIhpi7nBciNnW5uj3kXz1/LzRZ0tD4GzDV8jnXzCa7A98uWJUI8i4wrK
leXRu+95/dmskzD8MRpyHC+H0fi7BLqifKPPsC/i+SRFniNLrDt9jdpvtOHP
gqcygrrS1WsvVVlwwclVdqnjYRP+p7joN/m1xkB2TiHdSvA6Edv1uDeLbfgp
mZf22pU/jHZo/tNXhAbhLS2FRg+2Im2pCVuikXA9ipPGKvIHmfUJcFAXKjkF
Ii9Hh+Fa5TT56NXyQAMI9bwzvyvd7wBHf8F7loY/6oNPK3WRnlbRqkmkeAhs
SmFNcU2YQhlNbi0hzylGnMyULqC6mZFqJ0qoQd9QddvdDsKsrt4G1v+3hnH1
4x0jWGicRFCoFdCw7D0/DjaqCEsMM7e/GpnrZIRdRjT1B7n9pC2VMNpwR1Mn
rZJcuRBaDtisrYtE+AOdEJXRr0WuKwWuEguJYoK8bMIMkayYt4VRzgOOt4wm
qIDqO59CJdgy0NqrEbSC/3DZNPtAXb3NiQbh69fHdox7VqBmDnvZ1kHVa9aP
/sgcNfrtka4Fz19+V3pfnl/zIRYwQTYglBRiTDQZfoHha/De+avCJlqciNym
Oii/dWIazcnDonuPpBbpU0JuiMPZ3lRT2iwTauX8CPfvSm2cvXF5myrkjKxc
224M3mEhkfutQYiASLqwqxD8wh7fpEwCQ5PNPwXtx0acY72GLk94mlpZvGKc
vxUCIPMJeWumnW5sR7hRtgFSeFdKT6N8DVVzXzBobUSDDJwso8voW7SdUWJp
Zq7j3c/WW88MzouuNqGnwcJ14k5F+dvdZN4XxtUgFXJNOmX37hWcukXDvUqe
w539WzRwAAsh9gma/oZC75Wk/cC+O/ahhdjkXKWTJ+yX5qSJ6yyYThi1d8Jb
fr2pHG06Wet0k+x/mm2dClaweVgIGfvUWfDNoletdc3DFD8ypwTt/SfxfB/L
qcm7McJ6fXSkWrYHTxC6u5Goox8Tf+MZKPuU58Oo8w0noPWoyYbldf4OZwVj
ThzPvKaJZ1dJAW43AcxnDEtojeVnXlhTB5ZDcGdsF+jEPC/vAl8k266j9/Xu
ZV/guypuPfODYeEA7JhJ/Gyxh1y6kvQn5umkbsOLi/lmWwLWTFM1sZfUt/9a
weudKwmbOoi6aP7YfL8F2278cC49NVC8JKJBBXRY0XbnY6Sb+kpRLQT/YURM
sMuRpaJnJoyd9C7651NKDaoaSm7lhMxjPnTTOMs+7CpUySHEnTOBwJU8kmmw
M2+eXFlgc4VpqhYczCe9dNJ4p4y72H4HaVYVUn5/BCgLL8/lHCDkwFCrZ2kg
g2FsgRd0MhlyNalAqXeE94N9BMV9O1d9lZrMNJ2fSB/BL35qz+nYBgEDNjWQ
W7qjOwW6n8/ym2sC8+cz8yQr+duU0M2WC06kl+hlwtC6E/N+DJtQdT8/fa7A
3li3bbyyhDPbNEele2Vww/WXQBsh6uj+Uy/ANm9JRpZ5SqwykwBtsy21qlUO
pBoM8J+4twv21UdiptEook51O3tF/DrAdMCEXKFZM5TFdZ9oqDo4XGm4ZRTv
Uzxz0WGdGzyG0Y62FWwHt0cYa1f7JxqczoK4JyBdk84xSrFL3A7wHQaIMATJ
tsmjWQXCjr/4YwvEAFXEU72UIQMeey/oXg/3mvUuBciHb0IG0HBtS1DZfA8s
h17fMaPjaVy0JO4WlgbL87SibppUpY6IweDM5LKWBJhCW3G4V+m+CR1Om+f0
L4yccv8j0reO69d14TTZgnZ2DYVQQ238wL/CMHS5mLt/a7HE9o4ywO9bRELf
F6u3aUEdXVkzn2I/RcBvpouvH4fV+eIVOyPSGdJ8mdvsukpKYlPWnPxAYJu8
uFgLuROAb5H/5E28V04LtyPBT5ti4IchNwhblBYHsPUg6dmMD9gAtkI4ja/G
3HQN8bIawc+H/zoLr2RMLYlC7rd7hZhWHr+dB3CkghIoQCGSFuhKUKWjFL+8
ke8hJ1kU1HN7u/Jxo13MZVLh/Lekv+3/NoZwtYMCM0CA4ARthYBBQTRTrfeQ
MtyMmVMNMQL3KU97hkAYkkbuEiQPk3BQUz3OuY/HEA9/fFdHGLSdvQ9CsiUZ
mB79qNB0hm74Q2tSrIWCNvZyRhdVdQuTxeQxCWEimEmjQhIZOjKP0fLGbys3
nJhJpFYf1yy1GySHs6oRvUyZyxp2qWt/71t1dtdy0OJKZCQ14J8EJx1Hjw44
qJAe0UB+PdSnbKcMVuVrwy7PI+k4pGl/HrhWi7wcaExI7vxqI717pRNzyymz
sv7SeTeB62qK/jeGWTqN1TnprRMG57vTbJKKHDAjqC6YinhIKlCs16/7NN+y
GFEvFKSiducSFNHW9NB+atcMGOo21qqhKu/U+eQpEu8oYD/YHn2Lr+QA0/6Y
7137Zh7Cba4CHzboTN5pJRCpl/jxOMtsPbcqgh3+r0cIQf/IZsY5YYSdcCap
y1bBq+mulqHSem3t2Sv31Ve3TNrlg12U/ST+1lPLRAqeubkCshRTWXZPgD39
aUYI5es9xh1uuOXs+UkRdxaOfWGY/hGanKJXw0x21+9t95stZIip3/bTLhoN
eqxsIR3kXztvw6bnH+i0rAjTF1DzAPcwfVbZwfRKcZ+KSyte5NN2GWTB5/oU
JXDi0SrVCCJH8Y6WHjQRL7TBMy8Xutg/JvjYk48snfVoKz53jkH+MWzYC1pQ
foZqGW+CkmUVVJJ7RECjwoUTLF87cx/W1Y8nhD1MT8MTrI8V0unJVB9J2pIV
OYXdaNDx83hI2wPP6hzD+FvFfaY4KsjNSAZxskHHUlTbz20Kebmvx/dQBhjh
xbDexUzF3fcJB3p02QlFxIluEox7q0oMYpVXFvVy6Hzv/lZFBXQcBTBPIZYt
Nkoq/GIiL7hgY4bhgxUVYna4YMxy+rJQQ0FXG+9bMoSWgBDCs4+kptGbeTqs
i88EgdNKbMSNZzNhbM94zPrpqKU1doqO5o81FqPV55bL82V8Y/Mdr6VTa6Ik
3if1YssVI+8uenWqKTaA4Q+Tbhnc3wMOA7RUoNgsFuFzQ+iyn+4cVvaFvvIm
7hM8eudb1m8sXC1twmOzWYGFWaIAGxHigsRhR3L+J4BK/qfKANyyo3EHmwiV
I3ii6NrTOV06svXzjCHUVL8CJ1JDElIgrh1/vVUfBldsM20BkFOYADduKTd1
7nr5ZQu/wSsr8CsfXTfMtznzC4PyUczU5CU0B1XjD3FaxmWNlPlLywNieS6X
HjoM+0G8BPRHoUY5e7bJFZzE8X8p+x0m+VOXYsd4srwAatf9jbgLbIhLJU2e
Ino+KvSP6WY1ElkFXQDUGNwAlNsu4f0fQbRMT+U1nB9mAXXjy5cF6VL/rPSD
hNkxhkik00vk8MKcg12WlOLpmGhhQtgAleMXoniTesSMnEItFELZjzmVVmPB
ocWfzOyfuWdlp67g2Makko3H8nQkOulrSS/YJAVc/Rd7BIcFcHqIY9XoidH+
1p2/nMlxoqaJfQGJXgjZ2XNH1GBoE1v/XgksWhdnQmEJcyH9YFU1okI9Vo5n
XWoPifkSIryxVF3n4v9y140RpP28QY6l3ZWltpfJEkIIsiNKZ1Dw84CPGZe/
EGWIcRBfNu5xNJbX73D4z3hxTSi/ecK7BAHh/DyAHqRr4YChS87S/WEPuDfV
qcJnLo2wcyl0l/KWaTk+sWpv6qnrUY1GUYGKrQ/uud5+/I9XU0ZQpw5ZkKbT
r6+8+dY0R4N71fUhF9s6orOKk8fkGJIgSBdr6zd1JkfbjrdAHbYj7kSJiN74
yW+EoaePchpiTHtgAH0bImr6JBW3DIur+I/djvMRE5MBn5254hk913jMsJR5
JaeHIYfXbYWb5wqAT7bvOwwIyY9t7bKXaDY9C6R+rGFWaDCjhV3vkzCr5K+v
aukm+/eAgjAhFL17O5qsiNvRqPxW34tXn9RYHlRG7xDVGsYxoQl+nMubpv/s
mEaJIiGWUHIuLqWtPWF1SOqT+yuZG7F1l90BwSEKhQFC3HC2lYFQcC+AxGnJ
6/SKu+Y8ICluk85KRDA5SUFIyKugcG244+FhHSeqhu9Ttd+EAOXBvRjW9srb
jNMIRCkVTBFhQmLeKvDiiLpVZSpXbp2q+PpN8gblmtixPcVcC+EEM/1tRWCd
T6of1q8B8uTTWdmV4qCp6hVrD1h9gR7pDEonho2SDaZ4xpcgUXjMK21Q+Xuz
Uokjt+hcx+CvDrVb+F8L7Y60VZFDCKT+vXGUKwQd4dafz5wWI9tzQgEN9G6a
uPcJwwJhh55SXveox+reEEP2f5dMcc6E0/S4eQWt9UWhguzob56pzdHb8ENl
KRPDJ1XMT7N7eUzDoKQOrPGks0TZmDqzjR3ARMHvrxTo3a1kDx/zw5qYivzp
iWnnFuZKTj77qFnXDTgMP5wfaTHjjlM0nconXTYLYIQRcg6UMJ4ZDgG6yn1A
NwFt7LWr7FtC5MMWRuH0zBzjsSkabzcZUPjkvY6s+zfnBhSj/5koJ1d97xgg
uL5QRz+jPgFk5ByGjK5UILB4Ih/q8M/gJyVphB7pAp9BCRSPaAK8dS/9KAIX
YjhIJuNTLYnJ41jfanEcV6LBfblGD50NdOKn5v+GINj86Zsmv7kpjUTy/d7l
Y5L0kWfCOpEcUZpXGcuF1L7+Q6vjuLkEN3KEKRqvknRxjx3BPFXUPbg/5Tmb
9jmSWaIzptYR4wLPJDF1MmelcXmoPkHxCLFo3u7rHoyxvrJR0/3ptA2R2U5x
jeFDqFAHMcoAlNvuY0g9MN6j78wuDFbVkcNjwMB5eBAM8AruK6xbrsVy2rvG
i2rFXQc1tS+48V4QjOaZgZV2c1TdXjZNXsIuPflfl/3A/MBFVqcygd2n5Qfu
85lQteNLbm8AUszTitkw50AM+RRCmPsjRGSL5bNTM0WUHxoEZUGxGS3ce/V8
9QKyX/1znzFUeEcAHTLq0nhiL1WhpnZz83aitvHZcm1RY5CPwl15SmXN+ut0
2uXq87kSkWJAjfqJwO71VpBxMjmiorh8Io8TGvugtrbHfLTeVBbD8BE1MRml
B2ERJkpIwdyisIzIJiPbJQlinNWFZtqIb44BxeUgeSlmcTfd4JiCgkwefoF2
SObJ6BI1/DLF/PmKm3mioXWs8l4W5d9/OxKNDyHkJdo2KCLlO0JDduv/HCgL
KXUmFMXV3gaLg1U656gnc7Sx72CFM1cD7ptr1nBkV1jMl38U/D7XymIHXiiL
bkSVka1L22XxZClIc9DzljtwKV7ZXlJTk3z+pR/FkRr61ep6hiwItYDtIFI3
nPOay8hukCZCTjc4zvcAQhlvmX0LdfwrzD3AWEdRZ+zuudAmxqDWxyFNODuW
Duki6wdLUjsd82isQC+3L6i2GOZu05ko2Yn5jY3pGCHIIWgD2rTI0RGevSpJ
5kg3NSCgUfHgfpDz1/gggzxn6N8sc0Kap/wQJBpR3F8IMoBTRBYMxzswRLeW
DeSM9487dcQsFt/YTMpQM2FiAzvtgzzILZL0/2s3a7kWuNpk+23M5aopXl1G
rwJxtstU4ofMZEUTo8l07t7x9JdSMRLLyUf1xfVLfazGEbGDIVPlfnlGZTuk
kvNrL6Sh21i4p/whJALaBpDE1RjJjQJ4qHUIQRRt3SZIu/4CbP7nGN9JaxUK
8F0IkK5jI6zN2gQuhiWCQogqp2mtbowRSL5fesbhkbS+lZNKdcc6gLDfWO6k
qscXAK+3/FQVgf3nwB9cRgtLQ2aoKv+VMNNVP69tPPVRMtVf0zpT3VpUEHOb
E+KwF7j30K4VqSifgPg0WJJZc88jcAwPpyHIYgP1/tuN3c2AL8GJPsF4ABy+
2gR8GAgcdj+oF0HbVATaeHzNDeLK+XvQSKswE2ptnr5xL+bMNLdiOlFE1Mos
ICBB+i8fYs9o+wuSTlkT4RKiNG2eoLO9KUTLxsji8it3QLjuLHm6EDMLyRMt
Aur9LH64jZs9n65YNEQPlPGMBoEpWA5ASPr4N49Mc6JuyXiLeu/m+wvftAl6
Ti0hg0cOyLK0lgY+aSUdeia98YLZsHUJxmsbB1euu+zTZwxk6kGoBN3ee8LC
e/ElIFn2zkhpZVfx5DlR3NAgrFNgkky8Sjj76xktx6uP4L0ywa2ZaRJIvJtx
dDwGelYL7NyM4YvQhxXDzlzGUx0GkjZ/nff8b+xaQT4uvgLtyj304ROrGmLo
jdgJW4ybFykvIAfAmnl7EPPGIdM/TKNO16BRcKcVNKByhNHKL8LD1xvxMEPp
eSp/S2SZqhoKqpYURCmkigvpRvZVACpxtC9Tzk2cYCV9gkS3EkL71gCYfIi0
ueWPNYMuZ0fzYhzhtplZKzzT/WqvIDxvca4z+wT2FCwb9nHZLKUAiwTzTTMa
6WvYZQKT1tS6yAjP3eLxfxJye1VgkAdHSAVJfaVkB0RK+vFZZE0K8awKgRjc
KCpaf5z/v/U5fghN75VwAuT/KdjRUlb1NTvB8MoRlo1HAGxhmLKr0ZHAX8JC
WuBVhevQDPlPHyVBbyvuocFhleTBdi1NCnZGgXzUIePnjI6F+QRViyGHoQv4
vSqjndbsYMT85F1Wbo5Uh3duR7dTuQbs+EtAyo35JXy6pM5PTMU+WZW1vqu9
aUe7fgAr19Cq7FJdpMpMsES1RXyIOFc6BFT+Y17B0rXt+KHvIov7DngLRByO
gcRbp+FKakZKC/I4e8iOMfBxlqqViD4NkFuiWdxKkp9x0jpQ4uuyzcB5I6sU
xkU2dEJXHbPPYYfRPaZ5q+oQSqwX+iJqfXh70c9ip4gDO3jOdtFDz/gT/DMG
Ca0CzLxZmoN+MvjXdfVth7J1HCeqtifBT1Aoaiqf6klDOpBAliIG6Qd6UapW
3EubxHLL3rdnLFiJn9yliZr8MuEjkACEhWqZTGdng7MXJbf5TodksveCqsBJ
mDIQNqmAgpHJsYenoTJWUwMJJpLDAm9QesCKE/UMEv+4LLuMI3dufmK46AO6
gCtMs/RWWjEjE+5kIvpTWWHfxkTc1C5njRbcmblDGNIOOI0LhasBN6ffXYeh
F8mC9TKuLBQ+s6vIElYIEHqnvrtuEgkkRDAhRdWgI8GQWsfCUU5aDv/xhJl0
BOqEaEJtIux12g06Y36C5NyZgC8WmLfthFLT4hb68oIjEFQ7FFBj6shT8LZz
2U3EFatwoHYWN8xZntraY533Gxn3oq7T56wfCsS9qAL5QMEYgw041o52Mul6
fXO0+jp+D+3ZaDUgehTnX4qMU0O8NTWkY2+ksffRJXhD/XfU1u8315c3m6vA
Yqj4FCnnN2Q5tONJoQPc4OwO6+Pxs+T8e0GSK8ZwBqAIomFtfx6in/xV/fA2
kQEV4Q44iJpieBurw8TWi/B660OAIgpwB5X/NpApH5PMTyB2nJop5pnl+nm6
ZpH5pdYbeFrRAtwbuWIW/prvfdDFX8mJ+N8Y/JM5pA2ZotgwVLC1Al4WNIld
x9WHeibYiWw+m8hHyyFtztfWuWPxHpQ28flxWVKulTIlPzC1pgnuQDzUTxLs
K4m2yA0JPlpoyNj0fAOhr8mDWGOxIbsPdNNuKP1a4BukJDr8kxg9lPN5jqKR
HrGYfSGtufoJ+AQ6DxxUGddks/Kqwx160tCnRkGFoWX3b2vqarYPjfQAzTZV
rytJXGKpWIdQ/+MiBZWOc2kbz7fKX0SCsgzjl0lgaHDVJc5p6QCOrLNISe8n
QKHY729MhDZ/nx0QlK5XjHcQPzcK/vaSxeNfHG/4D71f9Vdw2JaEBn80KJNI
xoxKIEIRKpUXSyTuTE+VA4I3kqDrLTzKHH1ZdlwBeNVc0wiJmOTOHqKmsQFs
5OquF3un5KdmYCeqGVdqq/J6+OMfXzcQ01FdBGaCDukOQezIVcMgJHeXvq2P
3AHq1+8kutSzga82P/6+a3YbW21NYDMwj+6vCZQx3SNoq5M29cINDkYQNCCX
E36kisO1Bqtjo7HoJMTvHuQNnZaA316x9ni5Wv2co7Jpfsvb2BqY0gXirHeV
YYVmIkRKvxDtggpcjUp3zdsR4BygCAG7cIwVIIMZWoSJHXKJBl8Hh8UaLkD+
Vhkr6aKBOtxTnUNUPE9HbgtNvqd4C3A6sI6Jeb4eo4cwYjhf5R0xGCXs/pad
uJ/glNKGPiGUwCPa1s4nZEFnY9HFNGbvvjhUS99Hq18weWQ6EFHz1zof8oqq
BAghZv/OKDPeILxZd5DTfbRNHeQn1TY2JxC30ojhWx2mjpgyZ9nhmPEs+1c7
4AZVMvcbMXCEhQmqVu9cGQjAx14pDLNfMAHw8ioG/33VRNrbt3sVUPNrpP/F
bxyvsVlTbi9tfwn9+jqajWgvEo5JtRM5h8YXqeDPRyxzojWjBIa5iuOTDqZ2
vXkgHH7r8RJf/xXRQCeMkejoToFvW9naHsuFZ4h5P4DlKO8vnb0HEAMNCoAf
OGUP+M05pz08CHgsRL2H0Etw+XjDBnMKETYRqiR6yHUUDELgy9SZaiU3+4g2
k5fceu2J84+DTHAas/I4j3ChL5Qn6tfJpmfhWCXzDfrO8pCBNbWRU+dFu4xK
p+1b6+lYCpvajBCjgYp785ZPbt+sFICpooxoR3OP3FMjWDK2Ev7iNBr0pZTw
Hg0MkqTwZmv+fgYitkSDbXCQbrnqE1967/YJxraoOIDjvazYAGyufMptjNh4
AuQB/oqctozsaSMUDSs4Re8HRJV+wESgOFTwoAK5QBk+w22CIUU+XVXTJ96b
sru8CCHbsTgSCXA39tsMO0rXUZ5ITMgwtD9/CqEEFzy1ZMjwTrr6CKVtyX7o
sXXfuPoEpVL8YfNZCfAe2bITCfOhI37ArSgXKOsUaI8mJihXKXOHmHrX4W46
90D0kua8pwcEJxipvLa60t+eytTajNPlGhPXBtfqzJvaN61GXyahNIjVhCzg
HG7807KkEBufQ1DfqvQvT9T+kNxwHit3Z3FkAZTwd9dIlbF4RYeU9obXMOmJ
tIiAxoyIum9oxvbEqBOzd03xvUbRIzdMyhs/QdlR8nExEcIgKsvSbWkcpzGj
O5k3m27wSDWGhwqiX5lxWmFR7PF7JzgNCMX9t311/tMYt1GTlReD46Ed8CSw
88tUVxKAidk93Sc9JiOKHKpp4Rl3TVhk9ivHHF4WhC4XMpVY/HfXzhrdTJd/
pybCuXUV6uk3B0SP1rs3gVC1IzKQwT5pk0ThDQ2OTu4OF5tmOjiMYJRAJVqK
dvOVqQdwJQ5cVNPGfZWVDLzvgxcstZtYwxbRAMPRiZhV8F8OhvA4uCy9IbPw
413BE+gykI472nHRkve2mDtsKev0SfbS4CgrWc7KulQtZGUcOrlqGNOtOiAs
Xg87MmNy8Hj0RygxCGinPvb9sFcLVAG3Ni83IxFQCn5yzgKg9ggG3ITL3TdU
vPy7VVdi7BuBhDDXHmqgp7Ea/nZJU5KvvkPeFDKCIzF27Dq/zT9cClUXPaLV
yfv6cxDe3whfLdmSSFh6YQYVsxes2R/m8B0ImDzC6F0IVTGxOo5iHkxQDcBK
9V+0jw6HxVXFHjWGa48ThxhirZ8AekhvaUM3cRzgR67AaIfb5tOMzolt/0vj
cr+A2HIhJIgNVNbUdecC3vIcqZIIqLL/j9bLWqXD/VDrIMe2IQXtc5PGmh//
H7AgLeYyhUO6e9W+9Po9yoc4VFuUih2sJdEYeW9Y89uW4CJFgx9vnf/YbsIE
9ZtnLe7gC5T6PIFbohnqqE2J4B8DrMnTEDhf66azW964QYNilkvOQZ7IY/jj
q0RfSz0/HjVb6WxvvGY0xlOieNv/y+/p0TM6o9MOZdwLJO1JuvPeky7MXtrl
PUdIBBscapEdAE84rCHHiaxLUP0SETGf4KEgVHYrpWa5cDy7RaTpUXVo7T9M
n0uo+nSRidw/aHLbebXtUJJmHLFdSLa2JGQbAwJEpfXz8n68HrWTPLkyWcuo
bzXMg/r2w+eguh64V6d1krWupNrFh2nOShM/P7ezLhYmQlHE9rvnn9GsAMmW
p/4ezv+mWoZeunlc9XTxszQQpT7fT7zdRrCb8KeIFyqcCkvyXqfpwXjSXyQn
Qdf58bx7jCJD/TOQgfgZH6fTmQ+tXkJiEBS/75kMqqgETdWxEC/bOto5uCLJ
3oEm420Lr+cFkbLkixNiF6Q3Xgne/9y0eNmxx2Ox1fxHmhdXCY/LK+BIho/u
Bo6hDW24TYpDlnqHDM/rUCtNsqTAcHUww4ujiglAiMaijxhWeHC9uCBW0w4v
OTlWC4OlhsY7/nWr8Al9L3UsIgYfumBUmJDSkkDZWW2aS6A2TYVbA5GrEoH4
Z6DMucoAg/5hjDhk5VWmxlllpC4DIhnKDl4FOyD6xvJHCjiGL+4hiA5teznG
Js2XMqX7zfkbHlHLEncYvZ+r5F6VztCviq/UHjET0tmGeaJ0p6U+LftQaZpr
/JHKWrqPgw3KM9X+I/V6Gy5iuTAGCIPqjDlQKeYF3RuLphYzkH82P+up8JSm
6ZRnBmzckXa4aDDctwTg4IehfHDjjXpWUnX8ydpzFbLLrWRyXNGNZU84ILlY
AI/jXyr9+1phv/djhlR8oekZEbdR+MtaV3mMpiZJLoN4C8GQw7/nuzru2xa/
eHBY4HgRF+SA9eCOcF5Hh+jfLrVGd4vXV52DjailIHrjse1qZRyFTw2/anNp
XOam94R7kmLqAaBkd3h2Syh24WEId6AtGXTMPapsl67vwqglgbscYrA6yEdX
3qyAR1lqW52faku6y25KyPlJbIB1YtgSNbBe3yQ93Kf9VXf3u1h8mUWjBunW
IfrcAyD2R3M/QHq14oQa065B8usKgFq2PgOs0SBsc8VT3dbnwv7kSP1ivJCy
43zdXj22lwri/Rj3TIMnr3SL6f9PUUIh0nuATH3J3WMLdrYOvr6HJAPaGbXy
g4kkKxuh97P/qguxwDWkw1lNAzjZNi0jjP5wefiBbHBP/dvzuZXYmago7fyj
rw3AoZv/RBeSIxwdByLisPfcnQ5ZQ6zAE5HD6UMC5vGEg19sfNt3ZXbsA3eS
cLOih3fSBHU2103DOOxHgB23q9XSzcZM3puVpJ0M4ASg9c6jxqT1xObJxws7
S2ErBmnvlKPMzieK4z/xS6D+f5cTMG75/jSGKN7B0AKJilIf6DKSn2b1JO3/
cJ6z2uQwERgiJMhCv9+tl5/jm9J9fvzfnqADc/vkTpw0idoHijT/b9GWoY3I
R3Ue1YQcq7UWA3cH30biuwh4meVo9MUdKGa8NZ50nQ3me8RoI9M71ohRPVIQ
7fJo3RSPVUrUxOiaOipnu8fYfB46cYo8QgXTaZArrMPs//B/5/qXn/74otaS
v49RSy0HtX2vezcRGmWO52DF+zOAdcbTi6GoYMaPd+NN2DP+par3EkIHjxaW
v5H4jRIGEwrWkpYPfOaZ3dXKPfsHiSVkOXKtsQp1lc6Ln7jZwX51xhqfWmvm
Aw0Utrn4D0+xZr+mtLzq/ueLzn/m+PfA6PDvNYNw5WKNgGVoxrhspmrPbDuq
gkcmpsOFdYLmV92UDiCBtd1U7nR/72rfg6UKA4McQPPpTBtpROebKGK+dzkc
xcHAg+4+MUe/zrWGHHBvYF87omXGopoLFK3lE1EdQfPXmYJitEAhFGS29Zuk
ITEX1g6AaGcRWX5kw+2AKQWNZowmF6haYk4lArM+Xr4lvhufwH3vZ1aq4GDT
pf1LH0UR98eBg2VIPKNixjFlmtSfumxhr20ucdxKC40cyFcFgi2rahV2w62Q
AUijAOKipxPcK6oRip/V9xfvPo1ROZpVaFds4P9wkXdAnQrFciyeZpoofU/+
/bxC+nzs92ik38CQAI9BwUZk6d7bZa1ZAnrCWjqgvCLjp3tm03r9YJ4ZfQqU
kGkGYpcKGVP+laHKOxrewHDAnMdegPqAblJYjSf6f9DU6NQJ8OyE1ZBcVdLN
6Wojv+HgYfq1QTgK2frfRS2w6Ux/mCqw46oORQFaCIE5GrMN1PE1mF6KSn8N
Bq6/QjxICeLKMxgDePw65PtwLuqf8c2g84M9xf5HN+Y8ePsyIMAniWyErTno
u4xqfl1bzO2R5hZMywLS5pXmLsKeACKKqqRN69HkXjoqCDFBdH5SB6eI4/rU
yffKhf3nXLdSJAWfeiC9Y4UwPh8j18rSN/IOekC61B2ljB701wa5jv+IB3kP
e0bs/FFAgx97PzB+zNb0cxxu3B+Kr+USwwcSRNtAYVeKzb8esTw6GrE6hvmf
Iy3A+DsUtayRUf94cK0WNtiAO/nYdg16KjUh6hTcovid7rAGEUb2yba6kgP5
EejnGLt+tQHqyIz9AGG4ZFLAyUdidSgC3RWmR3qZDVrn463arNQ0yc/1Wwlm
6lpFVPnVaad0JStHptt3e9JKaxAfpY3LE2CwbqOK71IqocGoN0TgiuilRHKi
yPztsk95wmv7ZKgqlQzESEb/7rmxTNwkeootfAnTb4hN3uCLThPyX3F0v0HG
9gPOMgy9LgHENDFKZKNPrL37NMwlFbHOajxTwgHXZPwc7UyJMh1xhy6HlbRu
eojQNuMjeI7gmm8+bkDECXa5qHHCHODzm05DmhboUUEplnwLJrMOhlY8PPjr
cknWO60FAUzBTU46GDGrDzNWZmyYQqbLQcGfRtcz6xI5r5KdgkX3R4SGrBgM
MepRxKJFFN2iIO7Ue/G4MYOjU1Xb3fNblQ6ZNeIxh3JMSMUE5OmsYaFv67VC
FQKCa18MoqZKuOSFFZPqvpZYEv7K7FDcv2uYQ2IvvTr2NwWHm8nH6+myB8ER
sKJhcsXgYFRpjcw1QUp70vhCb5Hmdqnkn19PUjIJKRcpZ14ef+wqXB4EPb2u
/AMnaHk1bjYqf8x9sSLOHKnvQWFMqEj1iSnaP57sMv1abnjHdKwJHdhA9zJu
P0YalAHYMBlvksdh8MnBDG/lEq/ClyHKhgdnjD07k7hx2G1nPKpUaqsoxO2y
SlePRVHDUDKTv/DXGcjoCebOyQIwdbPQAANnWSEKHleLQDiftYB2ZEyqf3IT
VROd62hMe5cozXRv6kUZis09/K/VOlnve4iUuwQi0lh2LzgkVAR72GzT8v/g
NOHCOyMfRhR66sBWEFJYuVrIG4XkhFCMYjI+hea3QAso6Pu14AA13wFUctf+
iy/essb5hBCbQAmtxmA2rbR4nlU8qCxPQBmrg8wovEm484W/mKz94sUpuenG
0cfeg5FR5eotkoA6kB7rS5B52RbFNn2XZyWqc0IOkKpLZWjcdHF3h27dS93F
DYKKjtOlYfIzgpZ7KQHmydHpXkVGttazJDcsFsEUaWqwQ/Ork3k/1ZhPPZSD
6z3KC5YeIZEA7YYxsqRfTAY1EoIN7xgbASTuB2oTLwKsyF6JOWJnl0QJgdIz
zsUfC9EA3A7gzHnDGw+qvvwnoxpAPvuvclfTiE7ArWoExAtBEC6VLVGQoSxK
Ph5tIH+QCmUJEqzIXWN3lHsberA0tkntJOCLeYd5/QmP9ex12TnI+o8imdj0
FvsVspCs7VRbAYTKeXE+qj5IqT/7ZRTF6dg+CSWZa6k5oklHwLElykj0j4yF
eB6MyJJ2hOVTcoOHr7FoXIUF9SZJQt/gVhIukeoyV2Oxnq5Ux7xORCXJ+11X
pdwC4oDkVzmlUztkrFwIlU6rV0OyTMwY0xRrpXzuvcRlPgQxh1lCDhwz4qdW
dRP97LFpYJnWHij5Cvu/VajWXW89tGp9780bFOzN+DBkAd0cN2RwhqGw+VFD
fFdLB+jQX4qf7hSVNK5R6wqDe4PVoTSHjVoesOpgauNGkalzQs6RFopn5l37
9nIJbmfBfPLIKlwQzqUbeK9xlmMl5vcoAh0O+OM6phrEsATwYIadhZ+JjnEg
v3JX7g+e/ntdTSDh/E3/oXtyM0mYKUh5RBHkzFN15ZjQqrCzgesTRQCMAn91
vOxNRdgZgJW3aeEvSNGv/WbZLI9s+zMz9Lml/4EBUp6+gov1R49jFK4NCTh7
XNVbsURpHEnW73MuAz4Mq4Kw+fdiqYrCq9oDhOZJ0uuUG7ZBGuE7DWlCwzkR
CBVebNor1zPyYCaGx8gBJ/Wp2GknC4v6t1iUQqNBWyNam6OsPko82JXAL5lY
3aydnjyMqtRIwky1Abm0Ea3VHTPSXOLTASCzoSSFczObG0lOUqX7xr2b8elf
7Icl63NMV18/XfTPm3+UUDUM4Unii6nZw2xuV7zlwbbmHjuOM2lh7zCxtCnr
BWc3Yb/i2QQBtqSg1fmqig7e/yI+542pdRAF1OI2B+DGXezoQWCDlXrQjl75
pJ61wzD1NEmnEEpCo9wGA8Y5p6dHpXVlgjg9yNk22KSC0ZLhY+enCefdFaxL
r70Mc0Pv8EOOQM0bOwrGSiOqRruuD3g0/mlXiGhVsY0KEcZ5OKSIYKmRSCsK
3VvkPldzvKL3O1u2P6HJkkoMwmeBtPfdoiohvYWm24MgQamqQ96QGqg1qg0R
5/qb9I9f+7m7mz3W8lh44Zb3ZUITne+vFsi9cPfpK3vFdEWFxcPU7P621tqE
GW6re/dlVq+yK59FvVp8IrIdiyPc46LGN4mwv42PYjbMR1UpPaAvXOdPSOu/
NsP1DRquUVG+VNHdnJjaYrfA+oQZeEIZDd2COoEO9i1E28hZMvHdfiDZ7zMA
lxeH+11+FSGqaLfqmOmTbLmJgm35qDY3IlwSLnjF1NEWZvlkc16bSaF4vCfK
cVituooM8qZivWelPhTxxH/RyTeV+j23iyGjSvemdyjp6J0BHtBN2jqcaXaA
QYKSlWwCmRwmE3r4DRhpR+x5ZVZiFkjOHOR9Epoo7C+v2pWwS/sqlf0cDGg9
bVPTVM840tbDTgQuvXzAn8JxXVDWOH4dlKTfPsqkGxrTIeGdVnqp8aOvmJZp
NzVVomXu4gyPzTscgrP1G36z7uxijHExzYuvaCE0xqZ6dsquqfAiGl8xinQ3
Dnb2lpacYpX6lMg7/o2P0rMpaaevrTd5U/TzF8KHdXCjMa2trmMgG+3zYHUZ
szsG/q9KUWEuMdsJHU+kZI4wtDvyoVVFKOTWv+UgLvbU4GDAvibDsZzmUy+l
waa0ZpbA2m8Vb29ilgUvaMh4j371FdbggKzj4d3EmCF+Jy6HzdOt3ERiTmn5
49aO2osUXEC+mdGtr2zNxzkDiPIQ1lscPrNXef5YT4uvLc7PLYTxyHmV4aek
mgqr5M7LG1yBlWFrl9e5s1OclXpL1EVJgnCQHkwFdjVH35oC6KtRYb1fbPR+
XNsXsy8DhPKguBn7G07gkvVZFSn5khoHWTtuut9EBxFLbVO6eJPS1ySj9gbT
zLn2wPhAgvCO9NY2rBqtLfAA+HXoGZXbUT0jGCnLw2rjqTCq337CK49KkEDi
rm8UxtZtXfLl6XUWle7UCA6rGGdq0h+yzxW/c4k425pmw+ibLRJWRE8qJeNj
DYzIS3OUUp5CGtX9AH4fyhoO+4MPq9qfvcYoYaqePnVCxUdo2+FT8/7bjcB+
zWy8aXCEShXYe7SgxreAigJYW7tT86JDZYtUJPPC5aEz1nOvQ+9MTV/4q0Xj
pfBuU2Qk3kDyynx4fdmSCoRFbRYbkrms1MfLk7N0G0/fEbT2WRkIb3N8bcPS
cQVLalBTIJDmINTCtI7HytqEp9e3KDIImyu+ggd8jO7VzpdfhKwHss6hc4IH
0mLDz4tTdhfm21W/qoCa4fAKwmQTPyOO0hgnwuNrqm63bkx8lRNLy1zYhbnV
b8aGR395j2+daSpncCLWCfxKJ8GWoi2+GcDEgWBKSgaJFVKYxK8sheFipSLr
/cIcVAV0ivtyk3h8r6qs0Tqc3f0c4npiHnYSX4lMCzl/XwdEDnPDLErlKyKy
feU0nqfLcXQpMv9UiHj2g0j3nC5Mspp++veV3be3MLNjZ8IZvsLVK1xeU+mG
QCWUKAN7kaFFF5om8pP4Us0hGLbXZf3AQAlB4EA3Wohnxk37lw/DHFNbxwDT
xhDCSdWydP4+AG2wQVJosOI5PRdvrfJVsbKuvCuh6xU5AlIvWOPLyOQbdSKq
TbIi23pJvctU/ix9IYuSQS57jtdb0bRw/JY5p1AJtAwokV2gFUZUPBJD25j/
Yt+9tDc6ic/wd+kAo2wz/SCtVXF/LsSCDVbP1gz6S2fFvPyV/1SVVa9pVEh4
ZLn7M8wGsBRrU5/bZ54QUCBP8XZ0NV+bNHOzNlmpPa8rp9kbfXS2fwdPzv0E
0Ri524ir7WHwoeCJIiowwVC2907RBRvVsVoDMzX35aaDqazEuF9YtM0604xg
H/a/o0qWdjWnNxBsErt7Z/IJ39c8V+DVqqYq3FvkOHZEP7SMqBSj1vYnaIcW
6FyYww8Xx+/6os/tukdEF0mqb6+XQrScLMcZt60t/QPPvGsbYJUrjLIKRjZ3
y0WGEwcmj50PG6ilYJoQNdqO7Y7rSwrjLQNEz7/5ZHtKvZLxYRR6aAYnZLTP
h8o4cALfkhsE6TNf9Y80H96XVab7PY3xLlLcvd2lSOXYO13Pgti5L4qPNyDn
6u3xgAkZbSWHnYu9NVDLA3l6I7iOreaIdF7JiQLRFPFl4eMWIkrepEreY+xk
QscbeGPMuz+1AfLkbylgXauU3pkgTK9Knckpida8KojNjbS8zK8LB5h0jEZn
hwOgi6vpBnKED9lZCvBDkPSO2ADd4FahhOe4rNDZcInBOTLcHKfwdLgJodUT
fGrAC7qkFMi9lE1+uonAaSnF/YPciR9SfTgkhhWdiNeFGX3T9/e48xGEZD9f
q8RoaWLUYGMAO6xLxYRtAJN4Y/r1Ez8L42gMl0qMLqu1MYterAN0WxV9PTVN
B/pqFSG+46q6EywGDTjEWXspfxQXyY/XIN4Dx4sw27JL3HVbogcAOQ19aVft
vTgeGEmP7dShRFkYpsWPzf/PE3Rx2+hb5jP9kW1y9tHGqMVXuO3uR5iVbnl9
xNaqVFkRhxuL48hTM+oWpdwQ4KiydV0uUTjEsURmajJpQNN/ih4qE92Q2pPL
jphWVSWH3QO/EXo5xmYOciER0bfEo51jsW5rSASQpljbJO8Kc08BfKtj6N75
ZQj8RQoqYS05GNzl4zOLtZtBbiwg9dOORBUKGHDokZ02Ao+TI2fZFQ6PKa0U
vlyAyye+aIJPpYrHv/QhkW1w+Qyr8cg4KkpOw3PB9kjJQ1aNJRHNdRI6Dxpn
qP2NVecDUx2H1y6H/KYHgUbbo1YvnQktYWXCZF26PlXtEkEXqorB7gB3Q4o4
PijBEpC382Ca2p8sKYKN7qKEFgVHzGcSKpfx6EEsipDyxWwgLlGJWotL9Utb
qhdZPL7xtG14ggVgkVJ6ScI3UHJyj917PhDJp/wno2ipGbFFFWl/fwH1zOG6
vyaG7/fzrPDKv8vkxIm/lgTn75HbM2DnbnJUambfHa96yvWPArkVN4LNNZ5U
UNAtNB4R4sCDEDZ9C5htCROGlz0Z6n0DwK70Tws2zCdYmRuzzosZVFPuvhR1
M2x6DYKzTDO36TaSaIgLcgQIM7AL/uL8BGLYnco4ZsB6ZsmdTzbB0ZeK+y0z
MqQ/gid5hqHIdXEX0MgifKui0Dqu240zSfhnXtsGqVigVm/o6pbDrZyjpce0
Gsg4bEyrQq6SDW0cgrln4qm47WVg4ZSo33he/D9JbbYTM4bCp82IbAy/ueSY
wVb3IzTqNhyBxXWSaQKa8bdWbRrDWhFE/zlZ9TrFT3B1fnvLHKQnBnyhMDPI
sLCh0ETyPwjsBuiFt3desbFON61bhNJwr5GcXtsINvgJIRlEmUsoeGj2EjBY
vo/CUJEWG5sj2I9Fyce56rAHnjDbFEAiE4dZtkBLM/kQfsdRoU+crE8p4PRB
5EeLig/rPsh83sEyVQhABc8d99k2GloIUP0USddQePynRENLtpDXh5RNBYrc
UhbWTMNxmr4X2Wb76//mo+g9jdhUQd+qEXrGYyasb3eu7cbX7tu5qpxmjXQL
RZVA+IxYXGB+Z0DgqqSrfiKbWI6mDlW89zJRMUoW/cw6mvf0asQvTg1vGMD0
B9U40xpKHQRlYhM8xKvxOJJBZ7jWKD82ohh88JnpaRTUl9+Ucxu+Df9CH01A
3n4taCFYpPApSLGtEebcCyFgCaiFIkZ8R3Yq+cb2cL1JPqUK66x6CkCWkuL3
HtPg+MgrbFA/0g3aWHE9YMop82o6h8ph66AYsERL1Aseav4qqd2cQD+LJbrj
HfEv4m4S1a/02CA8p6/YArCvQoQncY6vhBGqfAb6qPtrf5Yc/cQjDg3ua2ma
iBOgm2Bdx8WNbI7rEcc8o/vQMJYKPf3PWwd4ugNYIIaNkZHwYLBC91yYp4kd
h9w9xlcwGooDmLXt/WR15ra0bKGJsQr3Nj3jSUg/Sd5lCydmWSQf60Al5upD
fOf6T7NNtrx9xA/FMe2okpGnnTPOV0n9t/OvZ4rQGUFC58Vbcz2G5Lidh60V
JxVijgpzS8iyFDzilgCfEKz2HvCyD2ucRqmmaMT7m7pVG3V29gAG9maVWNoy
wW2oLG8nAqFqr9s1/H2RLrZpHzRhC9eLSSiMuuyFYboc/u8Ekn5kAV2W/LRD
n2qKcYWwsZuqsWqWRRTG83AsEzluNy96p+OYVjZ1EjNN5hVgTpt++IZxWfMz
iu4fVsJYEsT27xtR5bZNLTT6u0eoq/MZilJ5e54gxgsCRnePuIzJdcTKK7sB
EUInRyyivExqMtiG/s0Ao9qn6F1Y1AbPER6SOU1Tz364WfDEzrZAG12vEWBx
qml3xVfbAmr/zNO4DSVEW74tjzPeJX0fS1VieKBybckMyoyeHEsdL+KNTFU4
pbQsLc9Ob7/NaN2DbfZF9ru17k3p1yKvoOHxWjV0t6Aqzrw/4roZomlpuLh1
6+JRiSP5LCYfNAAKScHulbJTEI9i0FjcCHfZZN3+45CDXm0y92oy5vD+3kgy
vYb7nhQqLYSzWZhPWoekMFWhPaJ8D5xupftTelBK5s5wZP7GGoX+L5KuCg8u
K8HF8dlihs74XK6QDt/FmPYNbZXEezRXlI3LfiZjhN4PWj3sdMeChm44Znvx
YYKrXJ64BhSwuFwbTQ2p9ZUXkwQmKWrNpvGHoVQ8BC3Wa/X4Y5KvCfUDR1a4
osC9VnBu85tLUYLdJrhmC53eqDuQFwBW2QOgGZIz2dUid44HcP/sd4aV+MU4
qjqio2L1WMydmLgyhwaPDZRmZWUW3350kAI14e6I2lOAoioz1qWqw0duY8KF
3i6qoQH8ZJ6jr/uWzsKN/G2K+8CDegOkm8QsGGBfA8ed60Sg0T1q0eB0eO5h
Sf9hin19bobvz6I6uhHTpsY4UAkVzJqXbzFAW41xo1rSMC1886+AfKvUC31D
gDQ8y7TMfukfDeGxnk3M1p55+X+8Kkk3X6oX815FrvcbsAWdqUCON4nmuDpX
FcGE35gDKIVKFNotmzcBuxT5Bfm1EZWKQeo2iyQw2BKZ+ZZQcda9wPPTWoTJ
Ztispto+OKj3zRChtWS409IHdv6nifrpMtHCqewP6z9pwwIkSRnjVlzePWfU
VmhFprg84GFTCpxpfoYsoR910ANKo8PMesyFQUkgM7I1qjRGry9+aeUaNFGf
nk7tVG1pOBz1S2nC83grDOCBf8BFzkSPm+GVs/IsTXfEiBvAdooUuylt9+Rd
Ep9FbHkb3ZWWelKDZG8F7zWXVr5rh72UB6Balbi74HuI3ASJq7qF/wisFjey
hcZnbfeVmt2XJo6zOD/jnaEbJ/KZs3yqmZV99iR/JU/PRNnQCzrY+LIeVPwX
JlHCimHzYKzoQdZlgFDCvynMoqY974/YY5w37pYaBtgxABUiz6+gazmsRQdf
z4wWVn+iCzXbTqs6VK6mO8e75z8HtMdcSQa0zbUJzHa9eKmbkQHz5tc8CKWU
eYePPEupCdwOTsByHJwYbUjmap7htGTkBOqGrBMBMY5vrR8+RQEYACpWCENB
6GkosIfGAWKCBXyUZxSBC5Kfm8RX9KtcQKO/Pquhd+P9Gie56DvD0EsGI1Wv
fhU5XXSdTc5Ta3f1H2fmA4jrqurmVgKNqD6vUtfSgqYP77p1ZIyEwkeYg2w9
K3LQ880scifYShPayeNHRFbi9FrrZBQvmjtU9PSTn6sV+lBApDHkSQ8N0N3X
L0S/kYmELx1T55GARLQihlFI+q1enUj8C7cVd3YGZASjENm0a2jhmMbngZPb
M4yoAOW7/3rxidi6c3yhpn4n/mSIPwUZqggdpIjFFEE5Qdn27PCdJ6mFIBOn
R7Dfl3iai/kgrOBZ9yqt7oUD9r5rmfhTug0N/uLfGjBacoEMT+dCW2kYN4zx
Jzd8bg3PJvq1zzEtPe8YFLAYbVUdUdiDjz3ER9rOITqtMwwCeCFFVezkQ73L
0OclsM+yC0VDGhx1jdVM/qLf//N/MJydKjPjxOgc/zkHy91a036Hx8muF69h
3hFWWYxolWkx4Wk6H7lNhcyIOY2nsFQj0krpIjMgbhtu+aTzuAmrAhNaQw1A
vFWAsA8HLxRnqGV+XMWvjr+SW+9t+PuuHMbc2GK4p51TEABPHe2MLB69EC5P
Sef3TjtgYpjzl7oK2tVF1azDRHL6yio0o7C8ZNwI5fWlCbMG7uolcIpOZ5EQ
m99sW4MCe90xCmUjd6Lr8+JwiuuhFd8ynPGp3tJ71qJKiU4WfLdn/giSPKyY
PdpjGc37IaahjKH6G7BGaCJM7tM9clB/aT7tA04ghcM2zr0i5OqGRp+bO2ED
cKLZHdwztJczdS9SuVQqMNgr/ayUFfJL632te+618EeoEPjnAYhIZd9h+inY
yPVeJj9zX7mluBjx6QjL0nzxErLooIsP9rHYcQ1r+a5zpQPGFvAexk+JXq3/
tT7CyB6fwYPBFIDgfV+yAG6ilfX8OBOJf/8hY5ryMY2+sqzy9i/GWZLL6xRY
wKXDfJgcSCrEfzI/gzdRjEZ6vJjHlXAq+bwKNrx3iXJfhKn8kCvVuNjZ63T7
kSqlmUX3Sw2m5HfxQ+OFJkcDqPVQKKZJS/jP4T1utWHADRT4ZuyTOAO5QPy1
2IsXzeqOKW86Y4leiEHWLZYYVSQlG5FoT7dL80LCWxT3oFpbZeQiFfH5uSIo
LinFEw8MQpTE7WeWQN9/nKeTOZjRgVGv9KKzuJUKbp7AG6ZrN5WPQu7F2a85
Ru8FnWKbJ7ykXhVAddZD2y2N7fcCHpVsBB3QF7mvljKckU9eOtOxyC8zf7Zv
fy1qWZtYk4FKV01IL819jRzL2YwyHP1BVVMJaG7fn2SeDthOHPotiaSjSGlW
XvCF79Qv59ql50g8gX8qBVVXFIXTVTBMJBxhbxbjZEEzc5qow3ep4VsbYyjC
clHGrDv2Wkz9iE2bpL+RCgnkyIPRLs4wB77UDBq35qFTM+Hu5EU5+7hBQfJE
owcHB2M2uQ2bidGVZhaMi6H8d7rwqQSDqknGfM9IFoKE8Gi1BAkw93RfjkBl
T1perD4OrsXwfmee84iPqtPcs8r2nO/7/aBc1QJaoE5Ab4Li/UQJMPI54PGi
2ZUxPUWb4+2K9Z990OrhBriSHSd4GbREbaCWGkAhmtM1USdrjX9LuYxWSk/b
fCgbmw0ZHFWqvFpobrciNIFgAh17BJBGkVYkxg2s5B9USl9vPBHWs3fBe+g0
2PLb24ZPgx5FscTvGICWkWAEoPqg/JyZnXPOkrue3qgtmlrWHK/eclawzQaj
rrLp0aVzc7VESo7Uhg+7Kxg5faUhCjH3HJVF1GSjn2B1b7qWF7ocQKWMB96/
Ixp6iCsi+xyZd67YIZt1aAvKSTAqA0XTQY6WaqBNc/cfsBCMU7VBn/zfxeVW
3w8/AoqGU+noNgpSQ2HaSjRX7bKLagYBxeL/DR2MhWkXQZHT+Tah0XY/zemb
tM+E/BegII/WEtHSWAzorhO5DZbu9K5WtE2OG6BmY6jbQhnC+S3ubo25nF2v
hVZik9hG5Ie0/PZjsJFi2DwjkxCL70I8Rq4O6/QzmKZInpJgT4l/53AvcRcG
xc7hqjorSFiUoG8RGGngiUWSTOAWw+54MbxUubF33ulH0MMnzyHYQvW3v5XL
z1zD50ZD6/m/wW3h0PjGmhyS6X6xsWuYZbiszj/tdgzTQscQ4/yGlj/CVqwt
qBx1n7ESA+GztYVPa+wAshd2dqpzdvnJVvtUtXaLC2hwrrWQNt0L9EpDM9wM
0ZuNLiI+OQV92rITFiFfdO6ZdZn+GyEPxggjjULLZvCMAaK6jRFA+uEHGDsW
zWfl4trqt2KvuClHvn6pjznkNjdNXY6All7dna9a0FuMOGta5p5Nlb9cuO/l
5rUzZcXrWcXPQhqbKWrq2EDLyQuf5lQqKjYSZYPAO8AGBnz/hGGOSe5vY0bI
fPzlsLGyNx1VBVmYZYC0B1QK1B7vs9c52lQruIKAJz6o196LBZ2F/S2liKFo
9IM8AvipfcBDN30xXR7X7MvFCyNgLaMJqONmEeZuAfkTZzIqGAKyNKzWAXgT
/mbSpEXxTsqrP7luiVsdjoIHR5m5SslreuNk5rVIIpYfC6hf8u/PW05tZa/e
jtghfGqWzqO+8X7pjj3HGbzMg62DO0ctVWMsbLXbNcfC+H0pVTyDwbL3ZfOY
/Mxb34k1S8nn/mzD8MWdOy5JXCM/3FQ24YIaB1RwUmocOAlH0LsA+aUIDeF7
FRj6riaxl+RzSINtC8xbw/y7MCyzB8KLSNl9FImPsjrvJ7XTBkKyKo5m3a1o
sK0aCbD1wS4RflP1i1GWB2iGSs5qik26dozrxZZDJlKpOwZ5Q6neNnJj/U93
YRrnOOX7gn+XzFZveXxp2hUfgsYYxCNc4h25JBjd4mZvOwgraHjHWtiG5VrE
sz1xGBVRgqqBvxPhqPUYF0GhfQuyYZ4L6+BJF4INy4ceIu/6/tRQtwdB3cOz
jiHrtKzGvwg1X+AWKBsi/5clRf2FudNS7UGoYcenLBe9qkG9sUWmsW/tbOBL
ytA1cC0EtZP4D+NJFhTvFp0SrGmPmYcW4t2yHDTyAN9tnTheer30S8NQL6SE
JMl80XrzCFYdgYLT+zbmKWpQWyxG2iibEpy1+pZCOaktkYhLF6xNB1w4aCVA
FRT8UVCUmANS74nosHAuwvgPk/cX+bJK0GoKFTJgGL9H9sFvoYmiB644NVLz
HxHax9xk+wJxNtubfZV23HEolVKxqneXzwAGmCGhqA21Amb0ynaYDGUFLXsW
2PgoKUlY2eat6K+avHUhMaPYJpccipRvXPrZWLZKkB6q5tU6zAHLen8Qe63L
3B827/oZTYz6+jypZMyVmxYHGCX9OJNwb3TF3BkVGXMm0T/kUxDQXr8fkh/y
A2Kse+zkPVd3WKeRAElLbks6Sz2sQK1qYW1Vdi4hz7BgC2+4dPVGuao1DH5d
F/Uy4zBdCoAy7lPP19Su5prhZ1p5s3gSn/YIrz3w8boRLUSkRTj4bdHcLiLF
gFzpYnsMhl8jzIILJRgh94AXKC0SV1qfF27OeJvBybtyqwM1xNsnSrIi2tNE
Y4npHlHn1JvfE2K6tcmgqkadAJNXq/pkgxOEt+uk6XcZk6vn+Zw++6MrLa1p
GbGzUj3TlCNLWJW6+LLOtti4o+FNVc4G1IXHZTwISqrdEgmD6gn7cKEYWCZ7
QZ6uuy4iCO0uXaxxnZR2Khj/f68LMPzurBI/OAQi3W1AWKieVO80dlJOLpeX
cRcmKCFRvVvBp8adpjxOWMnjsIzUn1GlJszSRM+XZmVQjlVm2PoObH8q9Ab6
mH1Z3KWmnP5nmO+EuHZUv4kee0YeClq3jUhtdCn+H4vJlVkSg0+Jf4j9qimg
1bW8HxZL4B84CdFvD+XhgwsBlJW1BF+1qIU7s1TwXq8fqiPGNLS0pYhTx0Nz
wpZEdQ4q7OyhgNVADpbjRHLOcO4BOHwo3F0aWW3NilFF8dHA8RnqZCM7XHXY
2vEoFM3SGP3vu+42llCKZ6k6+KKX4SXivCet5t2IfbxpXFIbCTnxoHcrFA76
1lRVvJZ/0qxrJZpu+HuSs+HizRh0JSytIpyw+eJHf5V9eX8qKxJO0xLeoTxO
Q41Q1Wg0ktCYtPqJ60s6RwISxOl1VMNcVLp0kfDqmjjFxRqyfaOY4UIdKus6
ETVwNg==

`pragma protect end_protected
