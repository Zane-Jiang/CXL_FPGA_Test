// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
YEQyPA/n2+B58Y77CANvdF5CGINNWGj+8HvhHFeTP2ND0I1nvBL8KuyPue2u7Qr3
CSqIlYs/zpgqb/5a4Z10GwdgeSR7UAoOFCL80n4HcTfJbKD71TqxdmDLatRNRjaj
TiElxAoU4XWh0dIGb/3XjgXvH8QXRTWzQ0NmO9idD9QEh9QOYLPb2g==
//pragma protect end_key_block
//pragma protect digest_block
dfpy9IRr9t6EXRw/yRqCu0xVovI=
//pragma protect end_digest_block
//pragma protect data_block
Sb6CBNhx+PEGSXxpujNBxxPSTeEVUPsmS7o00Bwvp4dC0Nyd45BYoLS1MlUJF3Ln
upleAufD9uRWbMn1Fbeab6yuIY7fREKX/knSp6xfe5sr6rcqEuXVx4Nf6ChxFCA3
eAjp8XjNw1HF1ZN+/qdJb3/6WR3tvj1Y9eoCOYywXYgc1z3CUwFZGg6KIkkujt4a
KCN5g147d6/nl3/4pL870LRV8IVM7bwwnuTvo3dZmx3fbUx+/2GXfySDeoyB/g2A
k42tVWix21B8kOiMOo+tYmvKVi/hE6uG+CO3ItKOoYH9eal1g6RHlPF+PQk7/VfI
5lD/fZvMQB9mQPio1+obdTYAWja+u/m2fuc3Z0APfNdaDM3X+cd+5wda4l2D7eTJ
67YVTlflEuPi6/zxSm+25QQKqCzYyFD8J9fco+rZpagyIHTA5iRVEK1KwtLwLqoQ
sDPrRakPg7Bh49K3o+9JEmSCc5vfoG9BF6zqwXEDIUsibP/yGNB+h8VfFg2ygOMa
nFVC8T0qth7PiHW67zI7RX/vCUiCanTT+WGKAhuYrZJcztzDK1cjQv6ytAWPZgDr
400XgjsgN1OQyhDfNef2nyQllXKU+ldL+Te21GYayFJR+KvB84E0sGmZTEWzimYJ
wmHKdyOkSbK/rQ2z8pXWcWtYYJRJ5EFwIl6O9+kAggnEQ5z1FDkrKLThrFiJV+sd
VAYJ15IbUm+G/La5BG/FbuSEWCZrz5ao9hYIEPJxEKuVjdyGryWhhSg1FUXtqtmN
Gl9bkH6fQP7J3cqTpRAb87J6wfh2578QMtBD02ykz4zDWIWf8j7OCYLEILfFMjpN
ZYWKBuEGeuvNdUJXWF7KmDllVlQH2qKv36TQ82KeFNiaiRYDVZbIlcOC6wQPc39a
dtkHNMfa9HsslLOYdAAmepoER2ZEVb0PMo9pkUsjuPX6u7RC3c0LalEgj2w6RTi3
mTu1q9nahdqiZnjVcXSLu2lGCgaLluywPuRmAgg/6pUCM9Fh9GOoBGLLKj2ZO5Gq
Xt0xzYlEHzHrkFAU401wwdCFDpBTHCac0sn/eUoK7jzjcbvpOh60tQT4Qqzq1bcd
WI123CSVCFq8rS88M82rpRK0AJh8UJoS03UXEe8Hxcj5MTD9VjyNHw5oJhnixpI/
i3zZpEaR+yhoBVWd0EvAhPpD9dUHhvVGlNseqWryZyXrzRvjWmu7hdDmWRgkTUM+
l957H7ZoPlgve0SseFguCk/wwSooJWwHoBENmXqiOOtrTkSEcOCNTRSrO0YxMDzW
GPOY086jFlada0IVQJ0V44wmxmGSGz3qGEStXPXwmXe7aYr1+YQE/zxibW7dbAJC
TQOknybAp4r4NnmeiEOU5WcNEI2IlTuW+1223td4OyjLNqWQX6IngMbkVPibn+t9
RPaDNR91HfNLRJ9ZOgl80Vq9TJwZMMUphZKHAeG2CwuGd3JUOLHxbw9Cb+fyUlgX
Suy7zaKCmKV10FpK1+t62dxObyGA1THnA/COnBQaysrGP2gtmCXucMVjiFu/QvhD
Wi2BIr9VQH87tLuTq/wi6DoOEw3bwEpqWSDjPC0fpu4ifysY6A2Aogh2tXms7zR8
/OJLbik7mV1iUhYp90l6SDKT8GbYSNPePEM6AHnnngvhB6jK0pQvmGLpMt6CRGYJ
sSmk8GQAUT/9xFnbJIcfqoABXbI5+ZVqEvXEL1hh7bnnP6xwqYv+fST6q6VfMShX
UzzCr1EEI1C8cC5Zg8R+GjYN8tqtIj+UTawwC80rFORL5dQotVDGPV4lwmZnYgOL
vQ8Y84eS8FFbbNSsAeKC0uGhmAjvt7f3VchA9BpRxgxeVParTpMUoRh+YevFyzFV
hUWsG9/b2TNEpv7Naa3zqgcbmh5Mw810Q5ftxP381eNTlLNQCm1QuHuk1g3iL6uB
U7nJ37QAXOIfACj2h5XQQFVbtGzUmbdMzzeZMClX8d+0NJdA+AAzrt3et1UTdwbu
Mpj27c5awcKDxSBKYReAC3gq4QEUalf/Vy2t7cUAZOLb7XJ6XCArG3NyIrdUVotk
/HN3rxz2O7JXThLVWXrGa8xVgUTSSF/NEGrOG3uujLTdI+VYVt4IZUtCvq6fNUTZ
heSYP4VOXKRMNCyKS6CECJEpVW7lrQIz0sfEfn9l7MqaFYQwiLCpJOFjAUp0YPBe
IH4S9kTjEocmpxOR8N5Tgo+eVcWo9gfQBGHyJtlY+nlz5vT8zlboFZSoHPiFho2i
9ZATgBAm6rKKir7jwxKEi/Y1FKjWMqelO5H5f2n/xq37OsrSIltr4pLYQIzYXXV+
rem9icCjgcPgv1Oq+XYVq/QRevDkZRfr8ZX7orvtWCb78a+jbgBMy7DHQGw+kD+U
4TiLnH0xaMBNdee0wUx+4TlHjpqr9ih+yPZiABjciT2fgso8IHOl/RtxW3xq3R82
/59kq3RAytaFV7PV2NHv3a+h+IKzH2CfK/bDIzwqb/7/khN3DFAcauQoiC+e9TFb
I2TM4QTvaWFEr1XroTK+2GsbIvkghCoLskzh3hbW5n2WlMDFww+ea26B0UK63kCH
pqsn9aCeaAhUVf46YCMrfI9mpu4U1OypIZ1dPJfgBSFVo7HvlhbXQNF36Mi9aeCW
K0ROXYvPZ+m9yen0BHgtJo++pj84iqxBNycP+haHd4mViN6nPIRFLJbMwJYBaJLZ
phEhBl+tzpLy1UNv8dwteplbJMGj6YXlViRJQELL9G2YD4305b8ElrgRBR4kwRga
vXJa4pI9DpWqr03w6dwRLRnXjGCHmjUjKtusxCHhwlrpVEkTJVnhl6mvNxaoS1Zn
9NUXOGsvpcUBM6jzrE+ilpSBkLXsFekmxF4YYA7FbQmFV/02AGUVnFOIQxUI8SpB
aU8m5//7Cq1dc0WMb16CRXd9GIZh+I76DGnIZZyBD7moYsZaBWUjCsIwqurmO42k
PAmWNPcAe2MY4mQEpwJkfHKa5MDTY5vlaujFEr9D13D2GBr7LLKX+bxIEt4qT1hX
nLZYb55a2cqQ9Id6pR+7MsiMzAqiUSyTfbitHbVS9su9MU9ge9wK0ztVG7b6lu8I
9qi+P+M1qSTHM4Hx7r0XHbfLn0fjNIJptAxVdvw4FuGXlBKgwSO0HG5XGPAHsL2Y
0Ql5La6T3Ov0Pje8xInozKhkqnlnynR3jDcYEVCsHatFINeOR7KcmqkcqCQPbIvp
VOeeDCFTR8oFwZBrOBybJfxqeQsVX7t64rK7+quLKwfyQYyEkNTadzdF99Wv92Vi
2ZL1Xbm1Q57Qr8I2FkqPWUpodKfdGB/mg+SsJ3ZTwska0f3qPD0yVUwHUeT39+Qa
hDMNoKaSRVmv+iz6KilnDvUCwHOWjy/4azW4kqRjHUW2TtYgJramYtGdCp6tkMcV
LiUMA/Z4g80vhZyZCMrAJYC+OQWnw435TVnspH0Wd2DzM/bqYv3sTTH2UJUBGYI5
sHEGggIgcSW8fGhLhMFyvq/OYXCjb5FjYA0TKruJEjqEX8qe2NsN1T1XsuC08FpK
N+WL5XzM2l+jbQDhEYQVQLGwvfyMiFUWv2NfFPzGESv1RBbX5NcEWOMKs1YvCWeJ
2He6EaMGeP8AE24Ga9t07kCdsCTG0Ogc+UFr741FGmK05uAiq6VN3Ao5SCP6Y3QW
YP0Bqluv5f486ylzq1T9ooq4ao3AA9z1ne8qHyVBo+/797ltlKJFZFN2dyy0YPMH
JUmJM8dj3PhhU9E40+ODFtlpKPFneXhg1kQ7iPIpkZLYMpQisMow5RQXQdWq0Doq
iSw/m4+7yl7xuI6G9lmvS/GbExnf7C62PIYKStD32B33ArFpmpJRUh0N2qeqXg5P
dwmlgLHif5kqyf6ZrDL0pj/gowWVBAChE1QDHz/V4LqQa0mZfxGE1sY+6fYOkvc5
UlS90+TUfRh0VBwx5234vdnsSgFtIj3wm3xg+pdNfX2axe2LR2hJ+0iB9WnhsSsc
/Zb2gre8/+tMo6r15sO84y/rG5f6U22SFvUIXhB4yR54b6HGLJ4m9JUEsDDcaR4I
pUTy+LG+QalEF4LAHrTLURp+WPQsVVXjAOyIQNLa6ucCi9AOxd7ZdMO4BYRiy93/
fGg26Pj54t1gdN+R04jbZ22tsDOBkl1IfR9B5shHychPIHTiuiaCexpJ3LGFWwFP
tfXoAgHYWpetkj+uJBu4nube/jBJjfMbhPZFLjUXF6mFZeRvfkhvV6EimAUlV+md
kEI0lsyMZ4fT1whRM3zLAaIUTNzDxQ6uNYq0OCVEDhQrGb3uvjKmkcrVnqFzJAo2
xtXeLzOxezeTvCsKwelVrQV4t8dxfXi7317V+Es3r0IrrIjLrSMXD/VrNC5EUAu+
bfvoT8BZ4V+e20wz4QehCocbIv2osVC/4AydRZFrtWMeWKgoIjiPsXiuBrtRBIOY
0qgpcelnlK/fTX6n+52BzEEuF8qUJVrKv7kIounYWSZ/7k83sTDIRgXIUSo3bqG5
vyQvtieetc9WvToiPj6RA1OyIsWitbsQBv/jOU7yLV9kAutxlsCFFa+U/c2bVeIF
y2QVp8lQbbsSBXrGKn3HrIT/6PI8awXwphcr40f0tcv6rLDE9cH2iI43+nFJISTx
xP+ZDqoqD9PwrCivTHtQ2YNzgFNlo5jXtYYmC98M+nXo/Mml3PB5IFRKVnyJCtLN
LHP/ZRmn6gGnMrhxEj9gQBFNdXthVlDjJOt25YowrZe6WMy/J3HOnERnQGL4S5NI
Zk3RSoBROituRdkXOAQ7RKPBkxxoH7HgUypxmToFo0BX0Lv7X/z2HmUuPBMIN9zK
1g3hkU3Uiuequa5LSx8kyY8N8q9x6MsIwPfzXS7DPRJj+eiJhQAaMY0qqON/SYB0
AHpfw/1ZTIJLwx84PEKV5ey+8PKZ/WAYsOQq1EUy2RhV4RkR2xULn9MOqZQAyTrj
HMV1pMC8uIxidNlj8lXr9meDrLEWSzXRHEhnVFSalzND8RziMaoM+yVVRRja1yui
hrlsWxghrAcQ/c9YlwRjvCUnttBWDZYjTsZLq+It7RdnvQ2pcwLweUGjotp+xPk+
cXpoOtp5xHg/PiD/XHo+6F4bQXqbAdK8Rt8BMB5Z/yinBi9nOJhF5vfyZyvulF8b
b1sZYlpmiXDN/P1F7SSnhtJZ2EnlZ6oXLJcRpjYSuT7gdtgGJCwz+rh/w+Te+Gi8
tuWKHFbGEwExOhnmz57lEGhSRH7HRb5+ZguLk1uGyah/buRN+oUk7pylHA0/Kx8O
TLGlJ8ZyM4DX/+8CAQHyUB62XQc94eGaEVEQAE31WM8flYsbPvIQkaU06Pf/UzoW
F/v7xC6iEeAgF7LheC5ZEVmYl7zb6v1+Y6CmO9pyXtcECu2uCIFRA20xNg3FWtH8
iXbZL9qzTTtcFKgPB0k9ow6XYRY4ePU/cbrSEpPj8y2DtmSSuxS5rsfOTcqOfAcX
lkunekuxLHt0dmQDKCP9hlRCeYdLcvMfFrXCKOOwxWG/l9pRO+1XIdrOj8bhwAyc
PiHZeqOlm1Qt7fvdaIm49zAjUiNYAHwgXQ5klLwBqzlsjATLS2H05FJRDMF3vRi0
BqLuAzNxnJsd93JbnN+Gwtj/0caW8YzuMQXa7fVUNsrWQjXMtfX0DGVCQwV+Wbl/
ZnVdrCvVBceEEuRY6+Gjz/9i6XYBdPnGXI7hl2c2QLFFUDMy++XiBKP6tpnxj9pJ
4OTFmtRqB3TyUjAX6NiEIIp96TJf2jnOvW4KlKIBITenVeouPfAWouymEHFf0kj9
p1V0FU130yz57+/WjGzmzPHZnEfctRCHyjPeJD3IELZ5T+1Xko5oR05U+zJ6Dp4j
RhN8mwBkLFbgI4ingpO7rFpSIXWtgtC/vI+birLO5ApL+1VgWz5xjk3cI3UyMCRh
UMC/nMHFt+2sHrczo/9qwL2wJvstJqe+U8TGN/CTjs3bATy4iwku2z7uCu2xyqiP
eUTwuvuIYzqmuNUZq/y/qq5IlsfCQ4W7fbdywfWnjImCL9Rtx4Y/5Rvk07wrNgcQ
zzgltop46qd8CkxWv7bmafeu3mQyO4Ql9c2JcBnH8+oEt/1UJCok8LdExDiRY8Ox
9q1CSO909uGPhk4EWFWp+zRWsmgFrgIf2mVo4AyNLevysNhwbQD8E75K/xMdMwZ8
lvuLjv/A9KuvOmnbcuaLddCAPuiwIL7X/hP1K2uipHjE2+BPCtyGL8wFnD0+MdmP
vCA1ep/WMNrB6R3bJeC/w3Yn43ucUaXLgp20buwfbL9eBDcjVSFA1DjRXeYMyQio
fYqulDlV7c/HiS9tLz1cN7IRvXmKHFV5lKuU5LKPlCM3sbBJLn/Y4o4wXGKKugiL
zsvOeobR3WJxHTUolRD84IR6R0DxSMkkEKoIEvhiu3Xptp9ESvyf69JnAbaiSvdp
aowjQ7S0VnWwVEmmN5rZ4yB++8/bULNVL/9hA7otGPyNTwPFP/e7oWfjK5ToghZI
oS1Nph1cc4uOO78dZvDIWgFb9LP3tFiNOnNkL8i86j9S/TZawkvA1qliksJTyO/P
946SSjSbSSyk31OyHuK1QlMS/Arpp9WbDD3Z1l0swI2yCC5WNdIJYViq7er/sD8T
Gpvr8TRXrf7HLGo6URN/e1SDYOI+1sN8h/WooLo08JhBlfH0pfJgUWwokjB37h8D
nu88UCubmSySBTvcp+uIsz5Zr/dJiQqZIiq2Xq/a7C0Mi9iYtuEqCRPz6pfE6VqO
xoALAYa1VlaFKde6dArCCkoBsnmBpTlFOXn/2NvFEgIkXE6P4WL9CTpuy98YliNf
QzyzpWhB72UGeNtBs5z1KqjoP+1w0lBTr7tEMr1qgHUNWMorPqvyeTumISZcdakt
a0gfY90Ih+++GqZ3UQ6G02pA1RNYIfm8JQaOmd5tb6H2qPfLPaut6MR3KY5hV/54
6Tr/hNTHMFhARB5dwMIBDwuT3aXj95Vr4QogpntpvBkbzTN8cZFayTPiDHvIrZRf
zeHkp8d6qdFCy1vVxt9lJINkxFTZ9f/gXLFWT2e10LH09S0NuHApJ6IhlB9VsNUy
qvo6ju9Iw6HpzaC1Cjrnip36iw8zu3E5IPaeSr5eLKe0JLRzvkWpmAkjxGxog2hg
ptNwtRiMvZOTMZXPslJeI3oBebvhoBaxG4dJCCPS6A4VJeO+XfcyoylXVj5+KQG7
leJKqyyTx/QMEo+gdbl7n0p7tG6DCRdtD76hcg3YdiONHFGdNs7ZYcMXhlvngB31
XjtF+h9y9WlMfsaj+I2TDW7zNZiewJSMCbcZ49PGolwY0uGc54q9U1/GD22y2cbE
mpqCnnkg9xkRufnAnTNxvs21GdQGXj6IxDjo3ZMfG/PXmHk8Gx9ReVI7yXqLu+SV
Uqlv6IgSJJ6eeiTWlwMLoF0VN/DqAYgxQqPMmJFxfo6DkbKLWt58S3CP1hyzv67y
1dlSKopz1hbnMlvciHmkgWdJ0ee8lytTv/CJBzso44Kk03Q1LwpTrQmFmndFjNh4
0asqVL0hHhoLFN3aCb9o7rrkb9er4sX3uH0alAVxEtsq6XQOEClmqyvjegye+0MI
W8KtIqHzQilt7S+flvpCxg7YAHjwDss8yAPgxDQ5aFXwxQlRz/bAJCZmKZ32+5ty
FHqGZrPjYLTJ5JtfrJ9+WE907UlqfoV2/T4St60Xsupar04JQ2t8x38+RotFeCQe
ExYzJJI1VmKeSl0Oq9VWl2FTE/QO14xRBl8hvO2dUS+shfkRn64/99LrU66syKOx
3jZKJFGeSm1Ml4CyCawO7AECwPMBWGFtz7Yr634rVjkNCJ0cHK9WgxajocFMPR6j
5yslkqEvg0q4FeeCrBg1L3fi0+HHgvOKe897nwiwgDxg5o9hy+med9k6tTF34Kxc
sLHB5k5dNK9oDMOV05wpIhV3YAEsseTdp02OVJt/L37VR8Fe7uhLXfSRAjmHdVco
tvkqgZIjXQORHYRiJS+uZGCiKPufANl0tTbsRkaAelBMHOGd19ES6GbununGPgxH
dWDZyTLPDYLIbkAUvu6RjKaq74EA84kih2ONvyIOe6ZWqUxJMm2J7lpSsuxa7xI1
uSgsTLQozkNTln58WSsXh1CjIRgh6TDx2a5IEwhJASJxqrm1fF/o+gEMkBm89u8F
H9nlxyLsU9NTu3vPrq8MkPyw8a1T6FtuvDCSphmp4BAFa1OyO4h8FdmSzvDFL0KS
vDhcscJHiX13M35EnhxJEXUsGn2lBMDxly5rUJnNbkExncNKsud9PHReVN5RKWIC
QZ7QDk+KFPqB4z+8WAIqReSrJ5JGiMcMIqBtVU2GyTh4nb6PoeoNPzVEHV52kOru
GaDR/9784/L5XSAIQZZVMLVkn7E/9MgqAVqQXwLWfi95uhYDmo7AEtiGFccZDBqL
jqWH1gM+49HsRNPEqYarH4hvfScM2WyweBYmSQR9ionT/Bvefd4fnT0c+uL7pb//
PaOpLvYoeE91K3SqU88AKzu615gwrk2plptKh2b/HLM79O66nOte6YUuXdEDm/JS
/yePS4Fzj08zwnALUGkM4n3PoJmBTdnaGPDuruQ5ky7cKPnDHQPrEyJzDefX1eXI
2EkSsHUTCyyQCq+C1u8+zHIXIzHZt1LacDq/SSF9JCG8Ugy8uP2m9S1xSa1I1UWz
nV4UOdjXow1yaySGSB/I7pp0vrT/fcAJ9r5fII7A5aa1d09iNkV5gR+/TfbaGHBg
dLldT2vqI2Ndt7r5P8B1gEPQiMEfbnxpP8k2tFcJBai/7XTunamPwvxImvwoY63u
gGQXmkkQ8IY1r/Mo4btReTBoiTEufC47i5ereRGPPnZLPzbqBEUEtfXCi68SU5rx
CMgYtsIKLZd6Ez84Er5qpthWCTZqtg1ywMFSYfXMdFnqWrypeWsTlLeyTLyhWrX3
vUgqtwMshGkL5if4l2PhMpfAlkH9e4R9cML2vZchKh9UF5OXOupcdfzrwIX13Ybl
kQ2gFx8950kpWAxHrOE1roU70nfIPbEJ/gkYXrB1/1jh0L4m6nZxBx1+yzx2NdNS
mN1zs5RKaYypctcWr2JLMph0SX8y9tIYT7jrDd5IWultqrMtPOeau7QhljR2x5Zj
TlCO4F6X7XKuCE3FtVmr4KRutDHMw1945hwHx64Nrbk8Q1TL4FyksybauCFOlHOb
bAk2VRwueqTPXU8bqgm9eZzW9//wT44S++MWpYcefIuV9lkdK0KtLCjpj4+g/dt+
q2EQUcxkz9rColKC6S3LG0HW5m1FdEgAJHhWI4Y5t2RRM8Smuwg0qk2qZtXGhFzA
owW+Ae3RByGBhi6qLtKqSZfA95wRvhRdjjuem3udTbd6XYMhwJV7CcjIA7NMtsAI
y3MszJICmOFErJ+VMUp93D5aoNI66HyN+/+j7CRr5W9QyNo0ZTZkrryBfj1gzrYk
hthx6X3n70BG43P8YTOJhjxpsngYMoFf+fy4NKu3gSWwXUz3gp5Aq8wkDmf+jNmc
K7sOJ5Z31DgTyHACyijmff54ki/E3pE9ZCHZ0PxkDrSfXoIybYlOAsP9sKKcA614
9HTkrEzyVuG5CA+tfIzfPN/Jgg3ITPq5iKgqvWNS5IyigJl4NKVcp1sb2q5EXdFv
nzzq+oVaQ0/vmztyCuiWoVRsWHW7vhPde485CUULZf5SFpEbCrL/VFcJlQIQwBkL
e6x6IxdmhMPL3y7QOig0hXxTOZdX6VS9Ci3oQBRYEDDlJiBn9hvjw+ODdar6M4rh
7YasZ80mZsV4/0DCrmzORdqsw4UaNCvuwzu8SAyP+1MeAt8oTQ9hOmEKqOTTcf+R
742M2vHtr7+9nDl5bkUnKJ7cTZDqFVImMr5PTjG/AIZKBlgY9/KlNxkGUtBfFrAa
hGLyJTKWEHeuwDQDPnpSb36beQiGuXddzx4iXr6s8GpOswzsEclALQev3JDOqklW
pLWhYmrokMReJKpAucaLLGo2xpRWmnlsX3yoZG8wz+2sHK7TWYAKgUU9OLNr6FkX
4HYIb9UKMpdtmvTLWBqS03MiU5MvbkJiWJ5hc2ypegJyU3m1iQkZnV6gmukA76xa
kvxQ3iFR4LlsD2ogVr143Of4UKMguVp0/4GL0NHRvdzhh+tqW7ahUbdsBtv9NPTh
sQMASxR2ar7i9DPLPQ8/DqFry2TvQgVm3/xwUY2xmOZmk9UH992AzCIG8dNDICpO
22hyWwVNq/AdDL3XOoiH0RtSowOlx9biBbXTJJ1CIzzukypBIQWGQKXVug5H2x7W
01rvH3Em6FxU3sjiycPCqV6ZrYDuWo1m86Y8qwoqTOqFVI8eDKaN8vF5oO6mK7SK
pyzVxp/vTXbunzHD0PJ1fKzAwQPfGNTiZTu45ADPaWjwxNNpE0eVmjgPyPjUXjX5
F5RNgjGcROubgRiicMdFhfPj8Bf9jsVM8v/d8pldHh3VToKYC6CYzo2e2SlHPuEw
q0YnNEqg/BW7kOC25Q1Lx2MaMp0jMseNtxvAgvXoOwbMz2ssfSeWaFKND1WTJpCB
uqfFM2rsd9vbzVgLH0bsxhXm/S7Hs+5WmD5DI3LSKvokTy4r89dPoIwA7Yevn+Ah
gCw9ljjYIHkbxNRTIoAwFT1KOJ70Fc0OVWeKbxeSV0m+H8nNhCs14JA4Ht7KUGQY
jlmXkox5+iyxdIFwfeObIN9NYqHa+nu5ZEMDSVqmAodj8b9/+hnSa5fVsRsG4Rct
HZ+dhYALxhgAnBu+RYJUpdR+4JWxCnNUlvDOCWfBThCxy/lwKYP44RvoHcfqONo+
EI7JQIoaUNt/9Qizb72KncVEqS1G3Xn67Dac6A/kc3YzC/VM34H0HyCVQYuKq8sn
Wuea38sRf6AQnQ06WTgul694ZAcWvHGib8YDyCLaoLrQdCtJ9mrko6F3EaTi2YXS
uT6m3lyD3rgGaY7eLUKtr9mfedHoBXw7mROZ3ROKhLzS5nn61mMaxdtildE8P2by
HbdXxVEHupCrM6Ebf0A8NcdVhSUe2x9cu/9kMDt66qUA6Sl49N4u98Kt1HQUYUQ0
wKOY1r50GrPv6xYJ5OPsAsRL9F6r58+LfjnAZY3Nj+ASNcwZkUY6bBoPqCHMEh6z
gfPdNhQ/VxrxfHcNMstuu+OO6yzfbWJ1cvHKcEsyknL3kJtYQKvo43hq6aoNkhY7
EMEY8MOc9Kg7HZnchLLHwY0f/orYEpURkLBBjhheS5HCtH6azn7e3MmZgWupdc/T
jwV/2oBuy9eCk8oUpUUmmXwVWF/y9pho2cyV5xLoFvVE5ylAqGY53G5R2zGTLA7e
3ezWSbMASZJU0JYwb31Gkj4rQyIX+D7P8amyemZlQkqw38QWgb5KP6uC2CYGzyoF
puCXRsRPuUxumyFsHWqlwCmJXb10Vg7FsdI4VJHfS2LmvX9hVbVSzhW0z76+VJNa
n7g4PpXs05HjcoExosrKiwfbpErsRpNw15nc4lhPLy/emTER8poAY2sQ/XdY9SXR
2gxSPDtOXiVphlZfoQaMmPATYp9ms5x0vGqAihbJIx2gi1MYcMyaf83zLOXGvpye
97pvojipLDkYEXOl9dM0mlQLF2nBDRiLX/Cy/IPVUxX6RofVzqlc0RkkY9aMKrY/
G6VZP8AppvUt47ARJzJVd6AMalKcUHIRKuCj9isuTKPrKz5u5xcGvB6KdZLbWVE2
LkiTddrbElK/03gGbYIOaDisM97cuDrRCV//IyMcgNII1t0Z7ztZSwQRtQDcWSJs
WOPS+XQEcqoToumBQun5mPSxOMX4ES4+4Qk8WTk5vYlaZHwNnba9wyIKS2tAX9AR
HZZXPoWTUFKNzQBGybckdtIZP+Gs08yEipSVNAFnt4UKOb7+oKa6cSMmVIkEmqlS
2zJAmvdlqY5mq44iIzp2xNiOUqkbdi2rcW2giGthfVg4Pt86eMNgVK7dogfP5/Sb
reR3pLPe1pmH3WWSJQjtCYE2DIyQKnGbdV5N7hdNeM6WwFbnCUgGbrrtX1eivltl
uM1Y+oUIjYNs+0mvHh84rE3wJPtJYaPIzyNo6TQDCKjaEiSZ0rAc0kSt0gieYl6k
s3W5lCTowiCHJjxoa3p5++Nzl7XYopymXqraH2QBWOi/ImaFZ9ODc0/z+o8UvopL
YxIHJlZdvXXkWVjyXeg0dwD7z0NgHsUA08Zs8jRXxKLj3NUT5PIyHs5jqT52q640
3SMg7lmskh8ad0zqqOfsNwYLXVoDgMBAI8hspIDfCr3M0o4plN4D8K3JyyCYyz/d
HBBsoH1aNE5SZjWIsTlh+EhwhzyM/Ua3dkqGdbXi+I/CHIF3pBL/trFdlUNGGTRI
xyZ5f5ORyaQQx0qO3ht9qMYRLEsUad/yDJxzFVUYmM3WfIhbYuPkaaXeLstreZIq
XzBkPlw+pAQ5hJDb+4SqKvJ+uPB/vhKQ1zvZ5GOu8eAap5s9U87hRI5cnEG6Yckv
8oWUTv5O0+iCgIYoL/SkwkR1yLNmN9RipBfoo4c0/kJYWK1JXl4Qkuw1MpREpSGz
n0ZfefO9tLeMQsLDXGpOavP+8D0kVRx0B2kVclHOqGcqNd+CvarYlsHBBgexUl9E
2FOvAZ4CAPdbIx0SD7aDCYT9kih+Hn/tEKNeiKnOeEdX9+LNtWIHXF/xpm5CHlQn
IQIINzKGi2h5SbCiKXu/KrfZAlJd9YUldly6FHc0d7Cm3guQig+mm4/KRv5PisbW
0JMB6CyrJR6/zjJmBz2Vm3voMjnfpnBOAtFp6D2u3SeY3hGGLkV7Snn2sG9v3dMO
jkisagjyrxHIzW9AqDwgd3Yn9vI6knPLJ3lyKjov7YcXL5/ra0ACuHyDeEeOgKFm
Ppm7vIz3QPwSb5xqR74SfYrlOVYM18xFcEWubvI3NfZkgy4g906eWZMeeN3d8o/l
/qe9jLoivzpTXRcdAxDNkHOIKzdV98mOqEdtuVCUQqiQCd4KOOPxOgob9pA3fmC+
UkS99hjC4J8GqozXi/j221uI5xa7b5+KdpEqNm+U3MbkZxEAy1hs2zQiq/iuM+oe
ArnABt0YqspbdfcuRaFKuJNfztnn7Pb09HveuimlmswQ3E8n5iybQeL74zw47x5r
wKGABQSNK62tfegW4DxR7QUXB39XzsEBsGhuvDBuY2BxtN5VAteh+SODKqVtaIxl
vuKSns+zXSBomcWVnflh/+ipSkEAk5X/elo1BFcloE5AW9N3qrH7BIiQ/eYShRAf
CGbr6Gcfyg9RfXt9Fh97h5Pg6fDEAwVUsY+wG8qPRGGB2fAmF1E1mRuPNDso/aYU
QMuaue9MtSHJwXIBp2zqxccxY8rYZnjtnpn9/o7WG4InFLWJ59lDPld9aJnlRtBT
NqaufERH5di5OfY/gpw+3qYngYJHhWRp8HEH+kI7C8qi50Tbnf2hNeRbhCcUmDOY
C2lviDnSFhj7fLPUT5WdpJ+VoKqJ8mElLsxiTu5gRx01KzkBUFiF745TgV4KHJaV
ar5ZiafTrEmZACImvVhik1MeW9X5SXhLB3vguziky929CQGCR3aAKX5NvVFpTBUj
lP4fBMkuBHyfkevG4JCdJWQJOQj3AiTUvF/thmm/vhe1VorPhF49yLd+mJc5AGHZ
pFZm9IkoLt5egl6VbLUGlzDhg3Zl3ZpgkvhwVAsg5UxtRxa6nkWjFiJ8AKqjXTon
wPshAWI8XQwjbrl5UU2c4FfP5wboTvPqjFn4WpBDHniPrCqJsEDGzAzKMjlYJYx2
NhcDF2tjPm04FoVu9CwEYz5eC4tBYr4D2Vfb5Q/BJsSFcZ32qd0/UAaZZQ9mDRNT
ZuQwzpUWSQfK0L2VnEeSyADeIcWxZZLCZkNIIJsVTqowpU6SSfFlycdIKZ3W04qe
715l+nz9mNdqdfU0Kyn2jptdJRncg1AZjlXtDUZGPd2zlNSmhISoJxaIWj+FzPb9
xv+VGN5Kz+BeFFySMfGCEzo1OQnCk8t4XgdbbALORuompclHREc0ImBW9fMh6nTW
aTv7dxwUwQ7o6s88pCvx4TJw316U2V+mJ3RbSnSX84ny4dc3W2zlbR7GwK2pCJik
TghOi9PF6f0r4gb5KJ0LeH5dz6J0UAWPOmpkM1D/ybtyqZcEdQ335XeCFJRpsIO0

//pragma protect end_data_block
//pragma protect digest_block
u1Ep/M9iQ4odRVdA7MrVTwqkvsg=
//pragma protect end_digest_block
//pragma protect end_protected
