// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
BtuLGBxkq7fnhbHKlq2yVDmVmpfzIK8AcG94ZN5uMsfxHvy94YmOqN5M6aix+FR+
EyUD+fQQ8ixsqU4LPBzU0kyfYOkfTXtRqz4lOHswgYSWNY4CRTUM8ToJJSeWhmxq
QiAfSIwErwI5zDS8BHOF5MRaNpsTjW6lqVyN8z0Ee7E=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
a9MUgmszvF51x7gpn1cm2o71dgz53OkN6BsK/SprRSJrK1C65bqvEBxGcED0v5Sf
oCQH+UoDcQI3LcsJRSvH6s3H8ijupKFspaydL4RC/gALuxgHuAcEUGzE6GCKe3TQ
GGOkt3nyRFAQIEHb+q23t+u8LZxRhvaDLWfaD+naosO1tJRTRNDeOjPWtMzJmrjf
Ilyqv+fWabfYXaiQwERZQcD7xTPlcZQMY7ljz9/plj3lEYh6y1XO3zuOgoDdIMGF
ywv5U8Ea9H0h1xMKEXPMBa5XU7Q2Ee//n6Z/NTrlZbPn+q/BgjgUxLzhqyFzq7xI
DgSFG9+EW3vuJnm7OR+Gs+7I0k5BTKw7MLczWi6l/2soYoCyyia7gCMHULC3WXMM
Iptk3vEH2//f/3UpW9OmK7xMr8jXJI1jqIIBhIJt+ro4RcgFwzVGuqT7CwCy3DEl
WlngN58inJdlma2FxZhVFQGB9EHGh4agVeX6cISoLTBh1afaeRu7D8hHmJxbPVeF
dNGC2X+BKMzZI/ipBk5bo7j/qI+2XcJ48xtHcgA3HDsiRSy3qJytE7owbFLJPTEe
BHsm0K+CTx0zw4bf6KwVgWsA1D6KyK0GHtp8uP0kDz9hJ2rO2YExuzauAPcyZJdn
f9c+ODwy+vzNy0avzjq8bYpqrl+fno44XFALqnL+HlxantQN8Pp+Z8TZP7HgmAfy
cveqQn3kpOAUOxtSyitfRIU1T/bHa+M2Z4FQkyeotJ/8dus7M8xkaYtdo+kRl2/8
7M0kC7eOBQmGPjAZZEC68uPPZpVO4j9b9Ab/qnyvDvHJMf7jWgktXDFoTnThmibN
3mdO8/huhc3HnSK7BLM06uhR8jDJh7iH6PLnt7KjoMTsfOqE5kyAoKd2CPkTulEL
dGyKW4d48h3EoY6ELYeu/CDaUiRV6ESidWRBL/L35XVA9W8wGacusCfZI54RXSIm
M670NbeppS98sZJ6fOXdyZayHewstzP7k/VQbon1J25fEKTz1oGrELMqNebYy8oy
f9xeNGM0MW2UME794A2nO5RKjnvQ59WLe+fK3e76ydzwmxMj3zfu7tWaC2Okv0B9
qWro3tWOtHLVBOSm9H+0lX4LYQVvDIinc/vunBB4S+qiCDYG1w4w9ZGKUfGlr/xb
tAy+NJkU74yRQDREpeWaQakftuF3z+x/9fpAf2NDCeLbPtguGMHXBBpCv+JJ9xKZ
+wxiNt4UKGyMRLyLZhWenAm1Ez+qhgX1F/iFdIgxQ07EsAedaY1+dfpASS2sVumx
c+JhfErxfm6EOr/KLJGzN6hDVosoTmuaqp6xYN+1iyyw0snDm7irBxNq0EoBvVb8
uz9yBqQVitPx2rdViT2ksNzdyGgsGtiTnpOMeJAzoo2fW9yVZpahgeqZo17B7vWN
xZuIsZGTCZ4Fbu3ptjEYrRTGXgCPoxIVAbTZxxeuEynkHD0rgzl3svGR6GO1InsC
nwSksyoLB3blNJHQ5yEBcKvoJYDmFF+0dbdMOUirwOVpslKVCafxgLmN/YXTocdC
O6aqA1DhszCrDUdSPdEHElMKs3iEbdkqE5NLg3aHONVL4cQKO2h/WBWPhEJZ8641
ggbJuch+B/reUOxgz8HU/GjxQAZpn+PCyLi9jodSliB+SklbgmG+iYrgdCveZBn/
tZwLebnw2Zufj9bXrhGOGfZHWNy1d/2OCdN1tJeCei2rhSuDqrWIz2tqQD8BXRrg
lTg0d4aChTSuk/42nPApSWrp0W/r55Q0DLKt1JB6NmtqwPptk/Fp+ZwD7wlkJlsA
O0002r/+aPrde6y1rAE9Mm64nhkLf2y7+UrmeUFZ3bUduGNYDPXefPjKaMJUf+qF
l+heXugFf8l79xyDFouVFHglHWfjfG4MnjJXKRW0CF/4t/R1ExgIFlyt8rHiKoZC
miaSATn5v3BxR6MeejEwq+ipbCA7NvrrwEmqDEthD/M1ygQK4cYtjvUvIAwqiCGT
y1f7vfKUpIaZaOJlDr3f9JwUFWARWbmJ3T1gHOXi+M7in77Uf3i2aAXwTYmZIiRP
VV6fOlHHeTJnfesDElTp7Eo3rxN6CHtEePiPLaq/DcuQ+/s66uxwPsd1NMhUhZZx
BDfUDxYWczr+mpjgjaQXrdsbcxo0dEZI6WXySMlJyS5BQyVXnU6GobFV+TDFXq7F
aCPne7oY7pAtrIFuN7qlCYZcM5s3LMK0KMqaIOjtndpk5W8/wZ4f1fLKC0wQ8dGG
8YIBcqNcPZT9E5E20NXJ0htRhnKly9IiG9+RHh6vzKCNQ3gw3kXAXGCrAcvUrxTw
4c7FedY9SIKUiJL3EotrQYJWIqmwpxoaG9ZTbsSVYU3Ee6sHmmY84XLaBlJ/1ISR
ECdCXkS76yGBFt3FQmnbAHqX9TPihIT5ZDz9redYbGAEuS0frKKhblBr7aGZxQPc
jR4dSBHoEmOdCU+q4rhdrkMad/ifICDfGD1jKQ6mueqft7EnMXgmlO4qLguKJl0a
PqxL6cA/sFWeNmj7na8do3B8hMab947Uy+pSj+vW6/EvbQ05yYFXMIiszc4ToOwS
6Klvw894PK+hEbkfyJ+BuS3XCzUU5nzoGGv2U2FBVAxxpAYcfHP/K3vp8Wc644xc
HtAT/ksAW1kk7fN9xbY3VGdchX9pmygyKGIQf6FFOLLMwf74oDfzBY9Dd5pxovZx
Vsolzej8PQnB1VJ+JfoSvlegnkBa+FPgUIvbHjjsQ4VSkeHDmIW6daCErXmcD9Fr
rda8lSs3P6Pstd5Q6+sqRgQxHmnW295szlHo+Ngx2XxSvPjz8qVdwNa9qlrCpZB4
tC3U47xlQLjmyGvFZE8jHm2D7niTN2ZThceo8PJm0lgwm4LLVaUGXUx7mMH/yImm
oYd0nJqHfAXxf2Vf1+Q4EPeLPJWxdFK4A1pheAvX6VzXElOsrJq/yjuEOLcFjvvW
RO44dIzUoOwbToe01fhfIJ9qVBeQ1nvu2qBCzhs5J7xHqF2/p/eCFdlad5bXSYZi
09G2zLTmPtaZkV2g13AXkcNVGhiCmrh/mqbxxPZoxsgOz6ufr5QcTlOf7YUMpO0m
wAKHCVjb5kAiTlhlkftVdNgFz5xNWcnmFGacHkD4MK3R5sGRn4H8M15vBhs9CSWY
674UVIZvbPDyx3gvAxVmXEOVKeOBPJjyRdyOOB9HIZs+Dhc2EdMAEHFMTfeOKKp9
/K6xSevINIzw9VA4/Vvw7qcFEO1X3CrZHPOg6CnpjvgXcqczQsQzpgn7E0su8JJ0
UznUin/TfMokV2Cba1lhE+EEYr5l+Mw0S5Zwqs2/JH8RY1RZbw/TOZFAa0rgH3Di
QuIIGMWnAisxdAtvPdBnGZFK4MZMfu2y3JY+t1FYMwfvS83NttdEAmnh6kLtszbg
fMjUJFOkaql34qpubFjD9wIwZSalhA3TB8xYs3YBoKUNxQ4oH4CbjufAVWh65bm9
Xsb/ttytrzN/wHDWr0WEv6Yg7WRN/wn+HlRV/r/q09CbOeWYH+tvqMW4I/u3RVTu
kfydje8aiFAOPLD/HHfCjS5ar6nTs3P7sXfmgfKqwaoG98u4+gyWG4rfnOT1WooN
VIJhCI++96NOA6sntXD8+58JdWQ702zPZRHvoeA9u1Xviijm5h1Q0ydzTHwjNR64
1gXXJIFbd2MFXGb/38J3GGmu6QGP6asrUI+xXsYHrGM1AzWPH0758/oiSkcvn7EL
SL8hCT8/z/4wVG5pcgmdkYoQ5pFg7XDnKGCH5GUtKLVvXi39vDkTSUJLYv7deK7n
GL2zyBnGkDPUv2l1aumcKP9MhNWyGvAer0Ys/67+LixmjPw1b4/SN0+Vg+phH/M/
QeItgSZ2zFMaKCG1fhW3TwPndRwRele8NA06tfTw+Ob2NvkUxTUo4jBW/p8zOTZW
zHQ692TpYoq8fAB44I8qt5iuAvyYTQROMjptwHFYX+eGiAw5PnfhPTHdA8s/i3TW
yJfBvAbGVQQQ4/42ElIz5M4Yz4bgnWIPEImeSlkB3K2YV8h6PehQSHtyJRkoVFof
Kn8HPZIu2Ic5JpYZMbUUyooaRh7to+gj7UfZf8Sl/S4FoUPQFXFYIbDoiCqDLR6U
XjIairNaAqAuXKDz+AlX9LIGweoCPAlj9I17wFpfdoFFvfO7qaNWHcjakoJGIZqK
goqHnHdxc0p91Xg8MUlH+/WPCKjphwvTWBygjJzHgJ8wUH9wZuyGeoGh7qWlQlMz
qr4WaOkl20GU0JKlnENyUsfwPJhpcS2i9jiopWQCpkf2sDAGUdmjA+G7qGG41BVQ
Cp4M9+JtO0bSUA1/LcrgqBSTo4KK0gVrwZIY6zKNyc5ac+A2tjxsGseaM9p8J5Gk
5ghzt7wJXFlePRuXjKRa4JqhtJTZMFS6SeLCiDE/VOtKdMzH5gTIIiKN/59fKsxE
r8QLsZHH+yhx0onr5eK0UOHqYBrZSE6xKDGYZ4m3/BVt2C5IdNID3nVFbEUJbN1z
ekWfhw9h/bg580ckskxOGaG1nVYEpGA9yVzyz3/SCl0Y4q+GAW7QVFql3QLrwu7M
GBU6nb1ckQic1couB+u243/A0RhLuSRiLHBWFL0dTlcHef/Shy5QpxMESmQr46sT
6pnMA62IzWUDxkyGA9NEdV2fRY0JnRguNCV88X5UF9ImOaPpol6KE8o0iYrMMkuz
9WkKmGBMlzz0AW0MzSn2gYuy97bpi2wJ2sgTOTi4dhCFhlVTti2ee/T/ObCER2eG
1QRXjuZio8IMn7TdR4TZoylK2mSs9oQ0PhV7k8lYlUdfYOO9aj70SsfvWaW+FOvN
+6BU4PdCmdFZ/lOlbUl4cAqC82gce6ylOj4oBJNNFPNLvBBUD3k0l4r/Q6zoa3Y8
aHDeHFW3k+6PxDafB1SwpjsMNczdOXXxVb4oYhQjRbGGzyHnviLy8chHFWNzSpdr
ajPI81O/1gwJaawGrd+Dd+rpWPLcQOIimQ3LnnskLvUdQgw8+/lEpidSu6c7BYE9
Q1HjNz1mTMmygw6lAGfAZXOSG9jyrSXcvHQ++U4JQNTD16jJVNtDFjp4HfMfia9O
rDfiLBrg1b6zH/CKQPqPwvBki9wBYEA7LjCN/JuUEGBk5bVOynWCrXozljC2uXPD
+IoYtn65JEVuP20GDTCOKN96G6Y7TMg7Bv99hE64tU4XRkQoSHBG0BHZcX4WaBid
6MbPbygfgpv7eFQtoior486174ceqAy6519fI8FDjwBVViB8GBXN9uOTfT+PS1PA
+C++LY3a+pjkbRysmeyFNh/aBk4erA/RBEbGqR8RSoe2bFaiQSi0AnQPLW0BsGVS
Csr0a421rwW3EFKhBeAJOV5cO8fXwSVGhW2NOpLEvSr3W/Nx9Wb/JacDNeZB1jBj
euCxVlzJEIyqi/hWXUvECh+W9AaXRWLAGV7YAOlp6jTbpwy8eAff2tsvtwANKP80
0uZRkl23UPIV3Am8pX/FFKfqeFS+2ON7iDbttwuys/kZS/AZPhtFMsgp+o0l8ku9
reLXaYyjmentGUwjUiw/xRNXMZiku8Z5QEg9qcPMTNALLr6eqTQn+GajCHcMq3D4
hUlAjNCVAEDFHvypmhrqTi7btavOg2IpiN4LiJ3zsAS0BHIrQOSRoRiWhS88mZg0
pSppRBrjnHml5g0z/DKga/DYJ/CD9dnhyxQYxhvvlL+nAP/HPmK1shu7JjHDCk+6
fotDCMF1T9OSgTF2nApYKLJGDfX5Sycly+RlbsrzhR+GlgKS+p9JH7NZgD4QhxUe
GrR6Eqa/H/7oj9mpAiJpMW7ftIqqSZWmsO1EHh4kDgY4eEDxTXnjJhhXNuu9YKkA
Xo0GNRrfASQJwmyYdNZoSY3VZWhZLX6SHC1dMgKUUZ498Hb8jG7igK3uvm6omiGf
iYmY/PzL3oU85IN3i3bp8klRaMDfUhvnTluQ4t7ODUr/oSrECaL/tntFfnhMfVEL
toj00VTgoW3sSHzUobCYpvONwQHPWd5owrukOyy5/ZkOj98+/vaLFTAonHlFT8Bl
Cvn8+TIAdj80H/KCGERDykao8MTjNYuDd9CAhkhFYP42UpF2dAC6RowZA9GPtoio
aJwf+pfcA48WWLZWUTCKuS75BRFv1LrNMsthl4Ja2eN0E2YM+8pf9YIlPn1gZtU7
AijE+jsX0U4qqUq9ANErHO4GS4t8dBYitK/PI/g44rwsu/aweqH7F8b2EeZVb+Ih
ZDesVQQpRCp3lQsEAArMIafG7WokG83wFzwsv26FZM3Eb8Y1ijOGbMge9w56HMS3
0RfO/LgIPZSxzP+XlqUNkwP3hcydL9oNgFkM+4AmfU5BCswL38hWuYFUI6AqAsQR
IUVvfssVBeQwVCoa8qPX90MNWSdWYKlUpJ5CnoE3OVvLSgJuMJFSRHPN/aUvGnX/
QnLrLreij06fcE5uCyEr8/tV33He7Yqz7Wu/n1MeZ4HuY/7RLMWF54Mf8SqpAnh+
QWxgDVhaXXhpQU0KA7aUosYUKPoe+3mKmjwK5EdcJWAtC/plgL3WFV2y4/9DLPjp
YXA87g7vzdBgm1Cwfvh2yzNQLZ48B1zylQNzbw2Y5t44ji82/g1i1tVTBxjDJuSE
SzVWA9V0oTxoEkIzXHPX9CCPxK1vAjYmp8XlYwu7Sl/rgVaewg8avBI9lLMYcR80
N6TQIL/1F7626CgyenMqL9L2Tcpiu+75qrvEQacyS9OXWglgKu7OKjnykNRKE0Cu
To+skpRWQAgthmLiXVw1w8lSEeBpAVSBm/0Nj70PWqUPx/g8lc8tYGbF+R28Kdmx
cOzl8SMDyjrMvtb7yFkiXTqhOk8Db1a1NjvAythOG0s8ArGoxIq8QiteNebDxTnQ
zankTZyMV5N7F9CpWbUgg6Qw4DnYinlauYWd8+woRYmAXXZCEKACoZ+q1G5jTW/O
ZXk3oN+VZ0Yt2AG1fubyKp+UC1zCTXBjb6ZhjleShQFHzGd8NvAG6NyFo3F+qqVk
3B3uRbqfrIf3C/6DPI9btWAv/1YmPXVnHifUMLUFtLH2gkYvS0eMObRisWdYo6oV
ndvnYi780MLT/ZQpKm6GrkiomzEPcfzWDTk40KN0a6h/X/rUUw0JDL9o9kkOoRgT
lwwB8S+MQWac3u9w0jhnL5mwSXa4siCbqNisx0EqzO5JyZB6aQCpGgLRrhhwwomo
4z/zEq6+2DQkbW7Hljb/frF3tU7kOAJqike6Itzao17GGI4V2oQC3uxGDhrorOE+
q2RpwYO4iXpzad9cWkEMwqWrf6DKWN08dnXzLbB12iIw6UXqPPUzVi2fgP35SJGo
hw5UVVYueSD/fcvIkeWlxZGk1dts3GG+N287Bea3wTXwWO+QS0bji6x3VLsv1Vuk
6FZW7IV+BHvCAh/K2gvyYfE8ayNbsCDGlfxXU0B/U6AnAO++up5xFHO6z7byi8LB
SVMOxPFyGgkh5BbhUIN2+O6NgZDqSsBHZ5b+c8ruM+4KBZXNfKR3x5pP+C5IJb0O
GEt010gFRhjCdBjwUyzWXJDZy15y6Fwrtpg+iYazvM9vOJgLHAz6PxH/Hc+maWpc
hNIBNe76XYl569Bw9C5M0Le32dC2FGhbsFsKo6i+ne5dbn1Z6mmF5VmihJnn++QR
rg5YXvTr1onyY+GTwJIrenbn8/NxoLtuBxC5k/Mf5018ofIGPz7ZGLNNaft3RiOU
rdYoqFkO4OYEfzGLmKFdj0dqs+5nmtfJ94cXPmVjsOVhv0jLvdU/8JnM4cdvRSW/
FK1xBvlhTJQa0uQjO5JuB0QiVuarBICccVUpkp3ODAQzCS+Dnz00kI7bxN9acKmu
ZY2fBSMIkOBG9hRS9DFo7TtKA3t2lSmLOu+7cTrBTb+bBmrLu3CWe57HZfaWtxpN
S14qRWaDFAvBVb8O4Fo0yEfaVMBe5Fd/vpuunQiWuE7VYq9ZWGI/VaohYYLL1rBv
6q0rB6qW6WjPgm4cPGG1TrYx+CjMmmGhKJ2y/6jlTB92n63PmnGWz7agNDJu7KnO
6pN3/ZCOUseBPfPrIxUHBqt1w+YwnEu2PdOYQb338q8G3c5+nG9f+8YLke+Ep53Y
il5JRaO6399rN8j0IveUhATbFpJgrAeziKCBfpktXBOFCHqk+4qUegTr+VM2uGm0
5tQ3KqiZEdB5SJXX2sCVCv3MAKN50JtuSJMF23e/nObZa4/n3DC+wI/A0199EpvN
QhfitXw6N+agCJOx2p7ptiGmIIHK2tMDj+dF/dWYbG0q8gqVa7MxAbBmHPiFtG5V
QnmedyeZiDgj4r8z1A1TYpno7ZvkcM+BQ/6nHsWZvOyUiCpv8278XrKb/vNKJ41z
lYAeTDYIOkcsCFdTRmP5dIbRfQBpux4O4XI03YbEh3rFnVxh2GZEJkSjFXuxqHX9
+qmPDi6DdlPGITZ1yLqcVaIbyvnM4ev8Dahfi5wNZ5Fj81zMze6O/1p8gmWqW8Dz
xCg5DA5+kVupirwOqC0bqOc4z9qbieE21+hYhAmj7wY+G+qPjibYupbRBESJJeLB
UezJ/Vvxhsqy1t8CNaP4aiMEPtmz+oB45o0TU3LKZVvQoo74vLgku1E2B4PqnsSW
DutGBmO8QUe1ISOw3xVyA0ac/eR6nyu01JVQVTpVckbxCRfWl7wyMB45P9Nh+LrR
/nLHCDyD7FZg3x2RlyhFm6nXbuXDobrqJwnZgjw8I76hi7lHZ57C9DguAmNm+BL4
YGLV0MFY2RufVO0cOuu/Q9YLV5+8fjEnjGDXwHKTER4WXxElnd0AsSwJxTogPzbW
OgZJGUaI0AII9UMLm8ZvJs8yoAKKbxsiJRmg1CKfjUKAQtLplEnOUa/Gzyktcp1j
TjONLDZYIlIJ3YriVIh/CzUbqMoJYX1tZ+ThL6u4c/VsdvkXcdnQx2kLdHgdx2AC
kQReuiEJ75ynDufonLFPsJ3x2YyiCasm51u8bN+qYp+DkTMObd+BBTM8RMllcABR
NESA2lLSeCAaSce0xSPpwOx3oV+ck4Qj2Yq12V2p3b7M8qI6Ou0xMJZkQtNUEEu7
ETXuiasrBAS00VrlTE6dAIoLFO5zqRneZ4UY6Y3fXTZN4g45RawkKykV5GXxNe6r
TCugRXrNaJLnlRzySjdOEUiziv18kKMbZMt2zCEw3FvYFMYlQnW9V75y1V304uA+
T5wOTXRDKO0/RG1kDRdWoG1pe1naN2pay+ZTYBJfxG95Urs7Ml+CNgicvveoJhPm
er+nT4GnksccaHcS6X8PB7Askv0JUtGyNUtV/SL4WXad8gp2Sh0mj5rWuN5VNToc
9nuUIFcSemSpe5gkWGOziGzksReOt8IonNqy6U47VtH75x9KcWIzIX/GmH2N/1xp
PpE8geOmgc9y6w63aCE1FyWfKP+Q3GZ+LXz0AMq9zjlp3XGuR1IY/dLtUakZBjFS
boGi0yugU0L9dwKDGDuEZoT8JvxeBMnYlAqygG0Q5XU/BVZLKKgiT0KWZclSmsb2
rlxRzkd0s7yGh7Jx7whBDHifHn9Kx4C0VbXhC1YwM4cuMeYDCPQ7HDClXK1G+2NZ
BEZZHP28kC3FV+Tx+4tvwUfVSkOtg2vWHuavEftj790kRZwkMeLEYXM+KlzxuPit
wVUyCaTUFZ7flkaQXLcHBnrxhumv7mQM3ZGaHUe1Cmt3LFZraL3baY89GtzaPBt7
3LCYAPDNKUp7w+JKuCCIgomyH+vfmdXRKoB8uesy9IhmSKN7f5r1h4o5512QYXtx
5Fwj1xvIq9KnH+VvDb9f3LRf5daPb24ouLRnKxMbi6VPFGH/uHQ6tpjltXLx+zLk
7Pag657mgmKkNzUd3Z1ZrzRUyW5WyAs95l+8eNpMGMoj15YZS5ZCqVPTWTYAnDBv
6/zQEPHCr+P7xDDkRzuFM15kQZCEtOaTLAXkvn4cgp3nu3HM3shI5AoSE+qPra93
9Q7JYdSQ2nO3Vj4SZocFiUAPlemhUFQO25U9BqhMjL0KOKrd4DKReD7fU3SD7wkF
Np/kT1qbCV6TY4UwnsqaWr72kvz7IOLb3IA/LmumMWXx8JEKe3DxWQWiv+Rkmekp
Pp6NIDRxexnZ09G44aPu3fTrnT5+CYNdkcd3Xn5wjrXI6+xHoBXWcT2hRbtQfTu5
u/ZziAPwzryvvzzDPGC4bjazTfMYXhiMnFWpFXPGiTleeQ+Xf6Dkf2lOrmfDnZj+
gM/or19HQN+tp5i823wuZxBnCao+uVNZuRv9cZ4UbKAI4/S37CbzA57EavfQq4FO
xvIXgvUX0Bs2+PqnmCbZEF7rBb/3zP/pvJERYMt5iSPjNd8uGpHcSSeDInx/imkY
qEyljpZVKpG7yh0DhcExy8LgbF2vNPCxb905H0pcE8le5Z51J06MBnoRp2YnY1wt
8+g5d17Ugm6Aj6Z0um5NydCoIyjTjCchcDo4V7q1+fgDAoEnKNWkS18Nzwc5gDVl
UPTNTLzniHcBSmL9q+m/QcuvsRT/rxIjnMrfceA6Muy7nEd5sQZrgBr/CyKoA5/c
nZzTXXC+coChndzF27LadDLZgdJDNJo//xRQUpgJshrRqlUidamOCl2glrgzlg+x
mEexU7tT7Y+gMEg1HMmJrQZhVqqnaa9fplE1QGEwakn41xY7URpS5MvM9XdliH4D
uYe75lS/1Usp3IYexROjMY6MCo50lXiMVjS2Zbx7Dc3dnULRJd3/XfGr5ddtq+Mi
NP7JDFhpoNUu8KRP+1j75AbetX009e5MJm4aHrXVyVTl/vU1W0ebmaXMnJhl+jui
Na77OefmIqr6SLF9s1zehtWbzJz+Z4I4aNDbGYvucgyDMc8i4uCmVl0gS5X3sd5d
lcSlajjxd48YSmC3Wxvn5Pfg3dgV2KekKfbSSQ8Kd0lDgEzue0lDgMgs94gAlScS
xjdpkbZhTffkAQXvOUkoQV/vJiHlfzWzlmXJqmEUOeQz/YgOzc2bBJpYbZcVedGL
H3vlYM+B7WS/pDAG/+SYkaZWa8hV2c5GorsoEoDrZXSjzUCndw8RUx1DcLkBTMBm
tfOXt3GbO4EYhorwItKmj2AYsv8jbCLYzC2IYn+aYV/Sb2gavoeudP1Gbm/4hElH
bbWghCSyrEPWCxD5DgpW3id3msNOP1cd/9kmf+QTod29/teQarW3nxQJzHcdXm79
lMbbvyBn5VrDqlybjwHofib+Mevq0hubKNzkqpLLaze5fD6rNamfkZVo04Y3IcRr
e/VGDSdwGCbfol/VcVs7dh+pkouhAnjqZ/vI5pyXObc4p7LARQannpgG59oW8X1G
eNk8KfXyAnlpAPFLgLfJj5W0FkocSvwMW0lE8rqYCMW5jqSMbrLBbaEV4ItuUwUb

`pragma protect end_protected
