// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O3A1+UuTNSy5k+u+IxGCDM/xybvCEtNv9eS3/uIYM6dj37GXrK8d77c4+/vH
o3XeAGnrDUrVzw4cnCyjh8tdqKxe50e8Y17GtrhDENlQ6HX0G1Q5QNrUCg/2
LNZhoeJQe3WrRxM95M/35VQd8Xh2z1ErKdP79WjLY8/K/2aeQSlV5w3q60On
0evU00uU9NDK8ThK0WpGnkEMBhq8XAAnFo3ER83KGK0ygwDS/epX1GuE6njX
JXFypvq3X1AMSCSQNBjza72lEX5jb4DClun1q8+d8TlSDyHSYu3QoB+R3BZg
9QeWdDHdhYA5/BGg1FO7qzceVIeAMDjrNxIplCzEFA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U3aRhT8H43mJlhrUvpT8tUEGsKijC41AMwMLpmfJTlmxv6ZKUCT/5tZmtFSU
Q122M1dWIId57ZFInHvK/zJ7ds7aMYTtdabHLXYk7Pw3BXP1mRz+8U675EAS
d4eUee8ZjF41Fb5R45hi4hxRntEwea4T6ueLg+jVroK94RKm+jKL3TCdTf/X
MoHAAdvlTDuQ92buMUmXqy75ErhNGkkrqsv1sIUiS7HGizTZ09rHJ5sRn2YB
qoX++4oAhLa+4h9Iy1hZd3jcOYOCHLBsZLMBKjB+fVkCpkbYmCfYwyLsLFtN
wtAxTJDVhmyj1G9J+qq9WbPhvmklJ5zAiISG0p/AWg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Q7F6Q367VUpcmfoOnzqMn28T1SbQpkCpqgI5ObDw1UMzZVSkEGYjdKRhTJvn
v8bChCMtHnXVW5M5AfbMW5Bqrxg1EqT4NZ6mdcEPT5PRk6HCyrARDjncFEDa
iSZleUy7LKsYZrMwArltJTleFMNChY4ev16IDU/4DzIsaf0plLPDSc60MLza
qZnzpUppI2OEt0gQ3DZhdNGtYxv57PlZpbarIExveYgqH+jh25A5iG/Nh+Us
rw/XJqZNZNTz10Pw3zzNM5eLaVopjOZsX/tol3KgAVc9t3K9eJKxv7a1l2ct
hm1Q07pb1Njn0dqsqPBj21PCGoTdNrQzPeeZN91sAw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IxVpQNKFVPmO/L+I7fuwKpEcbcBaRdwbIJKoQ+9cPgubeONCtmhYlzMTtjxv
EReoyWcAolO/Y9jIRynVJzfik/844N6Ehb08XzUqPwc66KazbaAGZsB+4Dkf
KQOLUtFWaNgN8aE8wDz6ZRO+HJ9HUXetuj/qXAvqrbklnP6rXVw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
YU4e5ttwq3lL/AZ+E28eOptBmIxTmWHUbFSNqODj8lucLOR2ACivXJAowX2A
EInHHN5gtl9BWuz1XI60ltw4QgPaTArMF1iu8wHuXuuSfp1vsgeMgjcG3zkJ
XgDUNNRA6MKFJ04vsVyYnjpRQPCjpBSyInFJx7apxY6wvHqIUftJ9Go8wY0g
moGOOHi9+r7sSsPImqPko3nR3E7euuUhCK5aQR5GrIJ16KXzl26leuSoodxy
nt1DKdjwRamfgFgdSNVVrxVHZz0x/a7j9hDZhiolXl02pP+ikGLlkPHIwQej
/zHTZb41Vfhpir792tZl0eF2WC4YBRuKSuo/Bk3UVZeAilt5Oc403qjYoRUd
6QVU4FggNgxYSeZZ5qaDaJP/f8PwR6iUUybtTSwswP0AL/cLGA2frZiiulKD
lrYSRw6axktahn1O4cz/BT7nfUbNSM4rYkvopXMJma8ZUXNRkwJkRjtMzY/F
pbGTeT/F5A+2xYhSN045i9uTszu7+Gzs


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nXgbyhJ/yjf5fHCButykHdVB1MoUVYrHLSOCvzhza7mBLLDH/iBnsM+gssuU
WItn+FtFeLEpOz4mzLh4EVhEnmuZcsn+67rSwl5S/eOUWsGIkr4Y4TGqxeJ0
goAI5wTAJRzfcu/F6bHywISWhfdsVsRQ3mk3sj027KmFM4nQrbc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
o5KZPCypMnztmB1T6dpPVvM5eUceOKjOv8bbZmOHtuVRb2I5l4tyulBsvVXL
oeMC1WLwFJaAmDP3IvYdsdghP/v2Ny+UJS+xrtMuUUSdcd2qHTVoE1u70ove
Yn32Ev0GiIx+hW26n2CyVFZzAk2lHFkyIcF5dbX/QmsyRMZ2oDI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 166320)
`pragma protect data_block
JjHF1C8xw0zhCA4SiCTY82fAZYvHvRslCrf11kFAm1Xt9HxLN3l03KcH3udb
Z7WE00gdHf8OuhCcMLGEl11SOAD1SSE01Tx4tWVNO97DVJc1q0jeoNPeZ8QH
HSnifvIsM9Z8Bpy21Q6zRFfW8G/7IqL2qqJimm9ztvHx/wzpEFETC9b5NL3w
Kd0TaD2f+kf39G/pnd0t9xv8vEtWVRu7rEgEkX5RI4VUEsUbP6reO/8+dVvb
Yq+p31EUX8x+8bRCjonsDaLP0uGkq1D3PNeMrx95E1wZc4wGz6C79razNQWp
ngH1klFkoOyEsxVr+Xv3iBsY5ZosAkFrGakOD4Y2SwKJKpMpQQTZ+c3DfusV
p+TImz0vEkv2OgJzK81O5m2zEC41mtttg11WsXBz8GDMUCUIKmRfh44cTy+Z
S8zUAQT6J1d+n9n/fwZTp88uV6n1GOoMYj5kAwvljvSj3lPtgr3uPyLg2DZI
0IAlz+D3QsNlbi4LYfm+XMrDmqvH1earQ6VeoO/M2n3namquFNYu0adCgRSi
15uAuty9JMs82EamsyN3tHb+Bo+E829GqKbx4QrpdviFecDR0q04r+rVCWOp
+5U9OmfIqeQO9WnO6UR50C/LkHIPPD5HGerxWP++9n9JuO0eEefbvc/istaO
zGgjlK/YdITlI+xVrA1/qnCeH10dcHoQAv/EWXkUJrxM3UlNXSykPhJgXmZr
L/OzhBXWKR3P8TkJuDr8N4LCToIW9QCysQeCZcVkjod3C+4FwjJqs8qC3cuL
6GazuYPb6iOJvcd8GxLU1CPWf6Ew+vK87pLJjj9kcgfn8pJCkm+VUP9yjQZU
o7R3l4QnOvGA4E1/TnwrxXAcAq9PgQJ6nA1G5VThYZTOW37rSCZWPL3AEH8+
laX1EaoDUhHFinRoh3nkaIx6y8CW7cS4N3rxpzAdJP9vJ+TD4fgS8PyM+etd
PKj5yhIJzvG1PvPro/4UVlWIb2lNNVkty5AzEVG7i7VWo3Xpd2hhCX9nj/Tt
cZIOGKkBH8fPoo0NjvUV9nxeyQZ/6t6b7wB2keQv47b2x0eXcG9wrEEQdBc7
bug/5w/v8jktdSIrlcRR0Gh4ZkwAg8A7yDcigWNhhUX/5eYvut8WUaea4R8I
X9DXHMUm0V9ffW3juaM6EQKNEnKahA4LjVyjyQ43/xJnuwjNWmluZ8IJoBLG
QoFA1HNym6G8VVRn/hO/1ZsKL8jjsfQB+kvh8/rAHtjduKTH3ztNt/WAqpRE
jia+YQfvtBLZ1IlSYsbI9ff6psVMC6BsmSZ7LzqrjHE5XZpBJBsq+J/AWRel
dT9cNFrd194+s1OBjXyPUFuHX6W8fF5WPJ5WGnqNVpIKuc7NM+WTbpRKP6qE
dxLAfcrFDStVRDTuBNU5K0ljOTW59YeFSyxTLOOqA5je4yOBYo4Yl4LKIffU
yp4ich+XuT1P1Sz1BBreAETNZR7lh7WU+iGsSCtisAeDROiv8clEdDnteWEy
8nnQszowFf1C/7cfqBMTeuPW3ZTbB2YwqQfwXzZZBsYInXb4bFYcoRmv4GJ1
VQ/Dp8qrOhW7YeljW7xIXMDjrvmZuR4iy0mvYgCwVqZqPWD4wd9000tkWAJY
I01aw+BIFushTng2Rxf2o79qbrtFF8u6/jeHRAvO0VghqnSlrjY9u2ZNtfGW
k3+A46vj/iCqkHdZBfP+BCJkBSWzd5w71k+MTzKOHV1w/4C77CMGRa2rEVvE
WJrZYJcZgW2FOwMUo/EPRK4pEz1CfWWtzMqluwV4bPYBGbjMfyI9lCmMTytU
Cuk4Iag1UnMuyPxdApAG2vcFOyI1PQFGoWWqal2mJ0IIs+AGGvuV1darHCoA
jpkIYSMJSDxhdcNMFJmuuSKwFyuZjebuvqz4/eMrIiBo/PiPipf+W9+SlOc+
83D6nzqkkXvlYv7ag5LmHYRL9KHNzaEpiOEKss6xP5L9FhK6R5R+IQQ6nTPJ
rDcY0bosHT5hMJsuNmJA9ESujJ49xqB+pUjpjFvZVEzltIHEAI/RK66PdYSW
eHM144OLROSaMwX/exUSHd4QCsv70ug3USQWwD7uUo7BCNCZm3HCXCtbQo//
IErbspx3KoXhpG8hgkuQgKkw1b+mvqQ2uV2ajIAJYuFJxN5ML0fgBzJySAP3
lBnt9EzIzmR/wxFFe5dm4xpbY90ETWwswS2tFVQsQTGMlBIqAh4iPO1Nz5Qk
cKQ9ceNYcadVaRchHpAjKPlgb21/k6ttkMAzSg9KSUXgzwHwJm4jHVUI8jxg
oMZuOFyqSHEIwkTAVNEVl0JaWAJGiBIBKr4qThAMSx+GwbpCaNv5uXtzHWXJ
f+6LswY42wrhLtlPS1a6FcD8Prcgp/AWSDQvaSLomPT2Y5Hvz4zCbSMRrZiO
axBYMY1WXdhyG4mAUWrPqRpQlsdVH9vLM7HhPIyk4O1Hq3HMxxslGKNuwDny
rexTOhWM7ouWR2bKw2UXb7iEm0qP5sZ7PEUAwCLhsa8DLn/h9YXrqCjV9qvY
33loYkL6Zb7fZULIz/PTQ78cHP3deoSW/F9LN87SktTi799otWj/66ZfWKLf
a2iRSPV/ogVyk2TGYu+BWzHXBB1u5amnpLxsN9oDivV+E9VK5595SsKOz0eo
pa20As/WR5CAltw//fiZoyo6IfNaqWO0uNe0UEiE8KYTlXOALnLZzGfs/Tqe
+EpH3COsws3rlpSdKY3zCkZSS0tX7/chYHhnH4nTncD0Zsojq+41a1bCfTBI
z9VD6s2Y4JxUBXn+kR/LUd+Jz58/bWDtePkHfObWIfhc9nQ+xbyvBQx3bAWi
BauVUBZazC4JQWSWFlMKXH2P3mDHINc+T/MeqPl4g6vaOtPr5PZ1wLpVJmCM
VLAGqEH4vYCuO0nEAjG/wqt071URW/guU16gCuWQux7xNNr7tI+vhSShjEwG
HF9i9yDGaNniCxgN7o0Dz9iBIjaoRpiK36AQL0I5hHcMSBBJYDl6esEhnWgd
J+1+0rTo5ql98BlCuwjGD+nr0hqRSrWWGIaSmKgTIUFmOgJojVXbZXqNmgPG
uon65UlSWKNHhv99+KJ7+AKR5Z80p9gS6BSHLZr2xYWWdLDSHrqrRx92HUiT
1bNFq1kziJcSE1Nr8mO0zqH9v1yDzFuxM5ja039vuLEfjL4z7qGS9NJTipb9
7ngU+djiuBCar2xWmsqQYVmlegVKTfuEjQfsUAVyUZrGVsAXav0u4eSfwJiK
JyDsWVdL8S7kxWryRFGfQ3k4yM6JIMcZ2UFLT4pmYcV20vHCN56StDSdt0SK
B8PdQcI2vI6TPVJDZfhOZ3PMfC2gqaZR5G9spRKpP4rgJgCbeJbwVd4twa88
g32fGI1nOMqNvdM5nwiMeFf2oH3woqItfHdi0BYDF+2T9wyDF5NNNQ/RxM0s
HkYp0AHzihsPLdxxgtVTBa/fkUVDv8IakWx7sOdtdB6dy1h3XiuCjViGXfgG
93FYz1hYeg8COl5HfUliIx6pQpoHtcFplZVRlKSwQlptH234kmSEkMjWuexQ
owtpCyfbUIZMtwH7UobxgZeL9Gs5QGWCUU9E+E4J5T+plXo1N3D6Lg2rggEl
wIDG1j6/LNM4qyZ4vUrhHxRSiHAblBrHi2tlT5pifnPFySCYgpN09Kp4ZxsD
tbE9gN1LkKq4G4csJs7bje7zWmu3Fu8Zunk6vDQOMo+350bcrgKZ1gHdR7al
Q/qJzXPHIj4ROMz7oU5uVZODdXCYIwPnDpeRY+xhDVNGogu23jK3xo1i/Mmq
SBTIMCOEYDSyzkod4JSNAqRTPsCiq4XFYirn7/jAtVHFXbAPj4DTs5kbAiV/
6uQ1QLwtMuD1y1qkxAR/80vHtP/3uP/a8cjZ+4vMJ0eWrsFQsutxxEgjrHAw
287YRv3HWrOAVimCTp9H2RT/988rBFB0pF4vxx8kgeu/lTTaj4NBC9i9heJH
+Eil/cYbUF/O3HZ8HFX/d6I9PwCKWdnOGY17gkymk7GvmE1quPVrCIqywUEL
5/y0OjhdhMSIH3VGdNHWxw6HCf3o3+DZhGo90YBqiJLM01cj0EoPqA/mobC8
q7BN5Z+P4yFuGFm7OM1Swmhnv86QZKkMmU70SzrknbcWMiXsm/WUWfkieShZ
K6Q7Wlf4D35LHQcat58rulFcAzSbEHF+aro6Ayk/iXLVmOYMmwIjlx0kPS/F
q+8CLbPmn/SFSHE32MvjopzMaUjKrZFPYFiGiJixLYUGMNJC5WhjPcLN+HPw
9XDDfiSsg1YXStup8xxpHMgaegjk7xLx51Uxnk09j1zN6spjDYaHPLoQenDI
+hOFf0oenjRJ9bAZnigpDOGjMwrF8rQKNivRPtbQdeGPHF/lKRhQ5YZLIfYM
EoAYQdyHhaNdyhWd9Jmq9CqYJGI0ieau3HtVofUZJKoAV1+8qr9eHKgIyhsg
ilVB8iq301NsuCrHYU/r5uc25nvz6EcrkL4JbNbNCH+oBGDi0hch+hyWl7sV
09WdGKszTLbX6dm9Y9czPLBeTMFQbapc3A1kWpX5QSsltAbPlwaEt3kf+fjt
NqPxLd9R2m1tLb0rYvtPQOSBaCiWKAe5boYvLNx8B9eqxz3+4K9w3VqiiNV9
s6jRd4kKwPuE2M+YQW2lqHBkHz3Ae9XnrQi2CRa2QZvAbt5Xe3QAnzMGosUJ
nOsKTYW0BZWqOMe4CEiVhRkiarvAniPwSZVR5Qoe+Ez+315boktU5/VsPjev
TuTAVW48KYT64srCnOKL/9QGZad6y6eUVr/NI1KZR+sOLa057YVF7f8zDHEJ
oYiXo6ohb5XgJIgkD+mqpNXkd5vf90DZHrgxGAOXnM6qfF6Tg/bN3quEvoUz
Myp5oc6ErI+bLGJtOp9bJBovy1Mj6yLcyAXJ21QY3Amtg1PcxuBza6WqSuEz
Wn52Jm0DmuH0KW0mMm1GWk4GM6kf1SpAweHCnkzPEcTWx+JdlNFpPqH2H3HQ
levI/37aiGJ05sKiAo+e+qDxm/lbfUEGbJvBKcNSQ+i5xV1+m5DgIKPSXwnX
kM+Zxa5dpb6j8C+yyJJ/X+HIKasgwy3QuPHBFaQcTj5Dk5bB2mKVNSE/1ifn
PJWxyUsv7JG9DfZxjry46hIBOUpnyV/kqYeVfiDcrxKHS8Ebtem5dE5KofFI
Ysymwh91siMQFF6csn7+vCbJhaF+X+hxOqjn6gEA7bXk5ISCfOdtanmdjoHL
Nu2Svs5tfpft4yZBjR3ad7Mz8LfPSwbadgIxhujNXlR0lQLmhytglWJIlQLT
YQrmGshClZ0uj4xxWiOorWpNAr7WBNB+iJcoSxFT/vzdTXR3ubp/gJmDWgJK
SQUf5kBoL1VLusb9lUIoliTkYvIQ+UI+qPqjk2LHwYWloP9C23i8RN8n7/Bi
jyJv8uCECyj17utfeKHnzJMaARwpQV8+Yj8pfxRcIrpA+2Sy6Eq63A2qDpos
Q/Ip584G1OG/a6ygcBhzbT1oj+RamrAioNerO3SfFmUe5z8HyP8scXNcl0X7
IH+YHgrfQEyEaozw7suqdLKIAFw/p65prjw5/Pmw2qp2q7xffxGVyNAeOMvp
7qY/c8NYkx3wY3x+rNUQ/zu7wBOwy4Pwf34aO0wcI56UTSeIqAfgZpwGRLr3
nxiKvjhf9HjyiYM/u5/KE6vq+1Jo7WSs+y5YbAlRd/mxOo1twyJ91RhmlMhZ
B6eN4t6oaPRFGrOHb1Jm6YspT9UcwZi3hUUlJcJD52/Iqket5D76tZTILlyn
yrd9SMDGr/zzKPEQZ61EpSDjwiUlkxtcU8W07WBz/02Bf+PNLDgDV83VZV1C
IznHMRzGxSvHgZm2hj7jsiDiQmrKC6a0JLum4EVffEo8AIfRxJDDpuux6VZE
ymRE0Q2PZ5GbRejQZFSV0p/LSCyPwkay+jGiAsLeXTHvthbel20KeIoOzo0N
ekTBVFsThJdPjcCE8WoyyqJn0TXg+pNbGb0ufLRoqS3Q9Jwjlnjy0sCNNX4u
M4EkaVRRppTTS0LLfpWuwznygpoMfrZSJlwqpBhm2IbSXu5FP6qECIUTmHgT
6+He+LLDsK0t2boCk0fqQ4Vedol2P3fqCP68s6BX7QcX/XtqJX2+HuXvFR6H
Xuld2vqN/ZLOca/sG8tv9c6cHugQmh0C/R0wSt+CfJBaqdzCw6syHc+rHenZ
btKMjYKHoDnKyW134DSYxk3x24thw4rPwbxJaUhRRrYjdH9WP7bOws9sNq0S
8BRRDGu5BFqNlSGnFaqMgN0RicCQIK/Hpl61RD5733XrWqVVokqWXcF8pXKB
sgwDGXoGrOWcTimrSS53XowJd3msotNQto+/07fP+hkPW9Bf1bjcTzktGkEt
2OSH+dadFiuEiMgsKeRU0/B2R+mYzch447w1/RMFhkUa1QWhyHbtDpy7aEyk
5qJcPp4uWpbSM/OQ+SDjYcnnqFs8PIhjpCf5eNsp6dSZEC3BGV5Y15tbYxkO
txMa3+sK2ZioVfYaeT3C3iMvNdgzaU8GCZe/UOn8WH+6PWpmaAD4nnitY9mb
dIni5WSqUnibKkXVAS1tqZ9A8tLXKvCG8om3gFNG9TGH0SwyRqbRQQjr5pYV
phPCM7XQxSyxQDjzx9PUBgWcPAUvbutDcEa9/POljV4rpkEMKRCE1L3n9ecI
BFe0kJ+XrfpTYmT6Sp+PH6mKiJD5qdl8sxA56LT8zvO9Sy0hI7z5Kda5wNvX
W6pQjPPwsG/iXMS82fQ3x2+M9JyrEU3Z55Dx2e0+MjygiOqQXvf/hFtc0QZi
XvfgoyyqaOWb2Pb1CKynPhpA7Ww9s3BVgpHBMmwdwrru9rZr3Q3J03exJ7to
TvKAVtf+BAmGdKgvP7HmEK6Xc46A0uP6qFE7LXl84a/74T4v91spAsDwlNUm
ghs2XkeKsxySHzkM0YwmWZ2Hib+6hs6aUx1EjdlOMPd5qWAvQgU/33I4hjas
SDTgDSvI1ZBm2mJrCi1HQ6HMkW7gvWsT0KFscw02Wfqu4QFL0Q7p5SB9DEQ0
tpB54fJ3WfsYPVIQlphloc0sijaIEY74IxZPZZ4Yzq63YAMXV0DvMl4xkB86
03535vynIr88tflyex0lgwYZuuXxbV/jysruT7kdJvqen0VZdHKiI6lo5+jz
1Ng2DGaKLZgkc70Zc8yqpwZ2nFn3+a8spuTX8hVwOrUoSXPJiiJAdcqHjHrg
wlaXDqWVyTH2jvmRfUnVmthm3uSv0ucfWumzxq4Zd00+3kcUGs4eu0HnVp4s
r6IUxzHy9+70CvgvMgxONEmTbvzjOQZlSFY8DQw/exFXSdSajuiT9VcoUsZB
XkqpTKuF7r+q2+oHlQQsa5xsrUJwvVzubOnmFIUQy+0QjUHpVgf3uPmc4Jty
iqWqV/wSEVvJBtn40wWtY7EPSBQqKZlKZ7/bqufeWz71miHYsXALyv35TUDJ
HP56wf3iy4hRCBezDS8LOtmAhCJdy06gBN2fnDnBEQbUlJCqqOZ9bczYOVku
tN5Qg2+l/L24wqCvxmrbRLScc6KhkeKElYmzTg3iAGnOq96Uir0HLavOB0OJ
3gYykgYNQCNfytwXAy+s56a8jgdREdx0Vewzdo7LfXyOfqDrEOM3rtJTQQrJ
yqMoR6uOxzbJ9rWZvHd3WZiQ8Zlu/r6KmykMrkdrNt8vGVXuevLg+ImTeNMY
7Np7TJaDenFkxzizrXGFs7oz8YMka+PBXhuyujdU7k7pljaIs9cUeUkbMxLL
cWeGApAkM4lPXtOdWTFJ2FX2COWWxVqCAA3s7zkvzFfEB8D2+kahxGN53nYs
skaXdvDTVJa0gxh8L8gxbbLoRAvekKEZyMv8ezdnG2e38jofWPOhk4yoCTFk
OaOj5jZi3LQ/u9/yFIi/nq6pXPCy57hAAhCAthAVwntWH+KsE7gQHxOUukpO
JfbrZhbYCkGdOsTVbgni3d3UyRkrCVwP/wbrZj5xgXD3LA/90lV0UW3vZGm2
IKdjbaePUrOrCigurN+AxJSZGN1CbogBWBDcp4eSnBbWwQUHhhftpWnGUmkL
otu4Y+YBuaut14SSKkRLfHDx4lr6Dzh0tHV9o1bWaoqc8wD4XLgkCCUPgn1v
ZF8arL9UtaH0xDu6UM5IJwXWsVcxTiaFovx5fs0ckiPUfnREr8CP7AzmORrb
sdoOcfY+XQJky0F7MqVYSH7JNbDzA1qypSad+ylT5rKjvHPslUfY64FFpP/e
aQlzEnd7vT4tGhRjfKS3rtijBGpRpzQjBgbVWNhA7JgZkht3ZgCAVRvB9aQe
G9pjk5LKSnk0pumi7525IPhad/1725ZPoatt00ueLRY4ItDgtaNEbVGbq0po
0PQ7SztIPdVOK0NJrGiZBFm/Q5bhuJ7IXnUEDtfBCOsQ7SBth1JWxNGAnH20
wwrzyYZM3hjgwG2J/3e/i4G8KKeV336xgDzx+sNXRFYdEXDJSN6EkZUMTKAP
5jwykpCGOInIG7xlT0EZtbns2Ddv127+RdTT7KcO7Aj8g4+A4btffAclZhiV
s9KZ6PqUm8kZb/3GORCem9FvxaOB+J/p25mBWUk4y3pNOSFSFXQzLFI8VtiW
UPxnBsZp56HQRQQgcagy4xgv7vRHxLJR0dgfbnswWNsSsL6giZKVP0T5Nm6O
9sTy3CzdtsLNGlh4I+1B9vkmtwdYik+tIAGiXVX2gWiVz6IkjYjt5HU5gWLm
ASxGG0BwgWn8q4R4EoBEmtIa6GJez5fCHT7wzLh4AgpITu6Izp2hJPlzWVEb
dRTdfnnQ77dd0x8D/wiDjrUlmslVnPDnNA9dhVB8gyP02RPZZ0NFYo2nA8gC
cjCia6pgzppV3NkEYWAsiHm3MExofnfv3+SRfwSA/3/yplc9j9Rsf+br6uRk
ha47cqU949aOj1OqyxZZduBjLa7ilv71pYVtrUg+YhgIMjo6TBYadQzEWfAr
hQTxb4E4b/wmIxsxJy9WR3frEIORLVxswXhQ8rQqjr15MF8OMiNpa9l5xkZy
lIZucwLoaOfVm7WevlJKACNz51RDW4L9UZKKW6yEBTIJQLfOyTn08ygqxXZh
Lf8MrQ93APkuI3E6P/g+PvHbgPBlQ++7SRzB+28vbvYMZAVPEeNXg+XLQ1mr
Utr4GQYSrHRMCRm0WgaoHi0GemZREMcwCupjsApimwhv6P2erAu1uJEKOcRx
TH1z5zY6/VjoKsnePSX9cEJX64EsEo67pMBE2v7LG/a+nw1WrcinHZdNU694
wbHbTJ15+WB600McLe/cGDYaYujBbn2ONDWdseOSzPq46dgkeMPpkhcUk1FB
b5By1fl5DPP4CRHuwSYsBCM/l552Q+wYsQcMID2L9rKBggVlQ1RErgtLUWUv
k5WkcMOdbOvh5/Ccg3rlaFL/F8p0gNwdv9ysVM/iF4JegZRRP4tk8+/gKBEl
ywPUQ1h6lrfXyDVwPCnewg6a0X+YJqAhBwGTRq8xJqR3pxz86UkCnY04aPzD
iihxS8zTeMlWL2wnBPB1neiFItahIY7mkzgnTP8ywkwC9LInZJ+r3cYuX833
zGDkaKT+PyhwuRVrkPv1K/puqSzkdyJoTHPGBGOAWwzrwmSmLvewjd5sikz+
YNUorb1V56CTS+Jdud4qOCO3DcbVAJjfLegz33frnIspDPo3W5vCcCmE+ldv
XEG6kG8APkRlfz7IWJbbZDymLD+iUjfPxEjL383ocCP6EOOuJ7ex5PfMYLvu
zQ38pANBAli6zDOWX1hxSB6a/beoGq5pNoRn7wfhR3avi9drWmCrYR2k7Df2
c4kic1Wkd+CmWRJ+63cTaaaaveZEasLb1KDCNWopUvXtdof8UrzsD+SvCcXj
fjqZ9cjNrDBkibggZlqstHJ8dmWFZEF0e887ETctOPZgDZcyCVLA2zycAJOJ
QF1AZkydr5FOjPXIjrg/jV+xB+w0YNmtrYOrXP8NWqgTCqwgvhCrDtwHc05z
qBTUNbcce3DCXKzGkAqxtGQG4z9Nmk4xjsIEaMVXOmNbePBxJB0Hmx6usKN7
/Dl+6uoNSBMOQObltaA0AUEEWbSGXwR/SIZ1GjpqdZc8iC+ilf95tBmCOLmr
j0JVYU/hYuOPdDebYkrTaBm24dTkJpAy/aO7A22Q+r/mgIVH+3FhFPAxKLok
ee8Tm7q+gOaWOkWDAOcwdKilA46zdGOQ9+F1gNpfsAnKW8yYTcecHQEE7tvB
SIMgExDV2OoWDOPekmneZUzmUzvzkqwfx8BV4iCd/1lsgDX1I+x7eGIZEncz
NYYqxNj47RromK8AbvoFUc2gcGEpa5aKkAfZJF2KmzxVWV3DVfh+/laj4DCF
RfYZi7TJmtacbN8jmeMH4M3rOT9BztmfP9ITTsXbXUpCuR2eIgtuzpS6VrQ2
ZK4s3pFFp27hXLNd9Dzo748J32Q9SKY5sW7lQOXqOJGFmxCOTwHIAjJxtlQv
nBnGopwPBh1YLL6HHAkA/WrQjCfiFRebfZD8F3gcS/6t/8fk06gWqyXkvCbc
+0EIqreF18Fm8wFnarAoJPQQWBr8Ave/6CXpoK0i+MvsqAHJdRUu8E2+a1nB
PdoFhhQmqz58tJrTxB60Zq5tpC19wXoSqaag7uVGcXcgexq4qD1Wy+n2WZGg
cg57ZFNLLc0vlQLawh7Dk8h+pTL+moFdoMX+OBLhixcVgu2ojfgGjw17XMDB
Wwt1JEh7hEiiEeRryJihbVTN1aVSGfs4HOOEoR8xoQpWNRmKijokIxp2sc/2
e5BOLu5tBH8SnP/8awJTBCGWosItlaZ1PFDMBuvk7YaaH1td3iq+fSuR5y/j
uxZKvqAYN2DOMiYYnfmjqIM3haRdCW56dJd9J6W8wRw0954JPWZDWg3VGkol
diwtoubFI612p5V/6lZEotFmqoWsSDGw2ah4JFoIv2QPMruuFccpdQJPYJ5+
06YmFfJHtKeP1z9mj0fAEMnT75jWE2I8Xp3f99HFP7ef4zqFJpaseJMJCkzF
Xud1JigtWzh/o0ubmuj3U+QUSA+68Aasn29onDs9mSW22m4C0qYWZW8dWTnb
uKpPYDz8+q67AQnjYEUUGKhHLOCC5eTmotG0LB1OdniSLtXnF8MWLYKJMWCD
ejwytu0aIwirrq5S4a/PF1mNhNdSG8csBkhmKkSlImEyN44V0USzOugTmpTS
K0gJvQKWPSG/lcVIdsdvJkWKnWNyOMiXCx5HaffY1KF+jEw+fNt+BZZB5pNN
yw84OEOd1PhNhGjG+r1G63N6N2ZwtZAwF2kisKbBb4RkDSEFzIPFna+sSSvk
vBSXvYc/ie2CvLIm2bV3zNnMiBJEj/h6EdUOi4+S5e4VDWJ9RXhPM0q6AV7/
woRfxqgfG0vlX7pClm0ZnfoLwTbPz1av/QbyA2TNSlVM9PepkVnfFNkdpJ5n
pRUppeU8ojEWkHeitzUTB6VsoZcDuTlx8GrnzNHismfk70Ym69oUDLAoTvJe
r0c2s2WR5LiykhYw+RoAYrOi89nVnlw1Zp/DEzeTmhI2ze2MuHwOsyEDAmKO
hz9+0R2WlbjNvvJGKKB74r3J0o4XRWcIYtpFnXGcoJBKdBVcMqQ5wqzjHcMu
mC5ed4fL/6IzLQKLfDoqdXHgJy4ueEmvie4M2W0Ls8nucIyO9s3m7L/M6JoU
jNcf8Ym+G/7a1MiglAVyyLDYEikqhbR3fa9R11qN4VUS6tICI/c9rjtYpNcA
ht1u2W13eXUGiyDeGjViJQwJxRvCQa/BrsEbv0zjkgEtenr8JCWsyhvzPod5
lZnVSOTgBonH4kwG2zcqsNt3owQpQHw98td6UzJdNB9w7DEkkCVfRUzcMDQZ
Xi4+2oRBeh7QQkj2CM/50hfuB0tAZ4q3rilsrlgGXZPb7VfdDW8FfQmQgpo7
ZLokZVxs4LppCnNHMVI0XL6bxzPpecVQk5ej2vUsQp8gUoo6Tmd2gz+cXkI0
90bewbljKqZpcZ6TQIfY42EK4GWHA2U1JUZ0MN6VkXTvaA2T7zV4f2abzDkm
NeWzBosha9CD+ud7alw2w432oNcnJ+UAYHCbcmQOpauk8DVXPZwei/Wg3kqd
aTXaziPMFe/vsILYU8+1N+n2ebImSO4YrkMrpvMQA49j+DMejdTKkDuScz8e
/sNMXc80WfMG6lIWePzmjauWDzY80MR4KbV9RpeRoRW8RCahxLQvjhTKIHS0
heOTForolHw3va4zDEkNpYZHMXZkoRGE60Gz5UJSfdFqBFNjKvWyz1xrVgJY
9Nb3D7+YlPcYRWOIp2pEXFO+/3u+C5vbfkxF1EoCyPC/eHesdTlh2M4h14W7
WjbxeRUUcEL4tLmo34hQlGdE4DvZpAotcXcxuhc5+/B5t7QB/BBfTPNevdsr
7mKJrKsBCAQ5O1+iVH0VX8agVgzrDYeTJhfIOGn05IWoW7HORxDzSQwtIb1v
OIkw3p5AbueDIy4fugxo56OOjMK5xCTL2Ku3+gmjm+21n3M6xljHOzET/z/i
jVB6W9P+WwcJqWXENHeHAEaO5mNrw0CfULc6vKBKK7stBVxR48Qhjk5LorR1
0M98AjPlbnEtzkH+NVLWCPiya5l9YTmkzNYn7QnXBgzTfxBvRKNL4PGmZikd
MHRTZbu5xFCAksUDmItYVHrMY9FUNT/StWz3/WKBTkioO9wbSr2kdIQcp91K
kLAsXjFtdKajPeAIDqFchrnBzBmP5V4VkShvk4TjNpauforRvx80pqXHORiD
QDH2TJUF5JQB5RCyNz5YZkyM5Mphvz9+hmdc4wUp7iBjKajY+5r7VF3EPgsq
RW14rZnom9UlsrHthC+wj8lKvh50lPegMc8vmD3SdMSRFX8pcOpu0uHoXJ0K
DEeqboVQFsr6Y2f2LD/etwmxIMwcg0rnl7vBmIeqZUXaGZeIP0L+SQoW4LwC
7uwuShvPrB98e+jw6sAzhN86f7VyfVMzR0vQkW4opjPrSn6aeeAu+HOnbnej
Wq1fAEGSOG91kyCC6ay2RSW/zt+5T1XgFDmAFt215Oqi7wwRPacQi08pA34W
4ecjb224lL6RQCaeQda6mNOBXHAFpHCk3vytQOiSARa5tZcLXJWhCglsEv0G
cf3WRHknWg9rW8SRusermHgDIBVeUlULBc0evlDTnRoEIQ/mudJ4/YTyoJqd
r1roHpiz1ys2kodBN66yz7Wv/TTOXx66mKi1jrR/kakKpwjKRaccSLEUEjgc
fl91CQt69r3MNMWdfixR5xQkSSmh8wtvGqPrP64Aqz1Gf2tUisuVwvIfaAp1
ZwA715Z/x4v+lPXrtLkgHPj0jDySl7ExTsfF55iGx4MRaei3UTXDN+HzrSSK
dY3sQl/VmWnZIaZriLM96n2pIEY+VIJ9GVE1cKHHnEvpfx5E8qV74igvrFJn
w+Q/rE/TjCq7GiN5ppDy/IepbMs3NYjSCjn1tevQft+Lt+kChArCVO775RHj
x7jF102ytL5pZ7SNFfV+0TTHG8dIJC8qKx9gDX1GZ0E3+1gbHNS/ZjETenUJ
z6yb1KAd4XZGRQ6wMyLsLNMj+y2i3fS8uaiUVpaKQX+3hjHhXLU8BFHF5N1s
0J672oIKHfLWtCQ0MPrr9qENOkYryX2IPCNX2tXMUJTJrSi3/meu8tdT5CHU
KsNlVYZTIx5kqsZhXEcnDG0YGE7NDP+zvFrgkm2mDl54ovVtfF/MGfRr5W9z
gF59OeF9LX15uYQV91F2lGwdumswzSxfd/9UJL/NHhQxSyc2PZhK9X0NIenr
uuKcMqRE03lB9xcOk3zK9F0reIIFxc6DktGSBW5fMSjlgcLrkmFNSKuLOKWd
V/55PGyFemaNPi0jDaRPTJ1keZqpc1izWcr9eUii957fzTsOLBuBDMvh1sDW
JLxwZKUaXrLQonP1/+yir8FhwR63nL89ytze2HQjTw9X0/4/hR/KBio9l9PA
5F3O3u/Fu1GBdTRY66DFP1Oj+PJv94Xgsh0eV9ZpPT9z4O6S0YqXPtdxDwcF
OF/1wGwTnMObJLLKLJHyftg0guwrPGYeO/bkwzhoedox3fOgX+ejFfRlFCU2
vJor4IfqMIgcDLPMS912Sw/GgKmFSseEqm9MAalPxLXN8Bx2OF/AeAETTvoY
lAAkLLeDHH4FKgRfIZBKX67u6AR5Qbr/l+VuUKPUBQjf4IK9h/tJSglP9BOR
F8hpLkiuzL9Cn07YFHHpWNpK+dJxJsmHA+93hrgl/ww/32ry1ot7QyRJCRZ/
zy1BujMpbcStEh0g998L1kHYJHEXPUl0ENmqMkdtCA9ZDPOaT5ftp3uSRHQP
jgdLSSbGxBOLr/XNlP6V0WhMm6wNTgpk3PRpI1kIExG/MNeC8/lDZqs4+NAk
FsHNJjwvs0eOiNZFCMdwN9X8GOoS4WXoFpTjMpBRpJtAUDOoiBXj7sfrRk3a
MxmRSJU53LgImEvtAeNyi0gP5F7KBrnJxPGalvD6tnVnJDkc/G/oJyWA/jK2
AZuexsfxuLiklIMUFfBuIMNuOwmCLB8pKSj6bV/3ZKI7mb4Bxasly1r8UCOZ
dxgtIhi271FC6/f7Ul4C4IFtweEsJ68N/mF0wntYb7zJuxZdBdfgQ0euBNRH
ldiwR7mmdq/TCWEp9qZl9kiXKQb4SJ45m9PFHqxKfXC5HG1unSxKoKTZPiYf
0Nd4m0dK1nZFiiEyE+SoCRizTyE/sEDCf4tV815oNlTwgW9oAnOlqK/vjeR2
Nw0AqaKwoN+9rgP7F95jZVt7CCTVEjPgiWTnfKcY9cCCjWLODN2+AuxvDoli
3pCWkpsv/xFtBlaCzL4gHa3EJzaYCizOXMPt0qIhC0eNHkLSLIEOQ8r4l0s+
nweacPh5ygUr8j8Vphd5kRtQXqh+KIbYT2oMfgp28m4nInElAeCwQRlgDJ0t
QpTzSpfjqcf2sPyw0m3383SnA1EDQ1v4qYW/gSX+Y0aY+muzTIjd1FzPO1rP
QekDga83oTaBYY73nE2pq8KD33I7Rj+0z5XL+ZEhQo0xvwpu1Zsyl3UVcbIo
8yD4yqAtIJBCFpB7HBrcZymPuo0jEQfw1EbePlbkiWa25pHjgz+vNNkMJ7Nz
LUImRmGxwISihcT/u0cXkrMGDa4gMldASGd7jH5cIZtAvO2HJBZgUgaFPmw5
ebfcFAmaGrPVAttH5JvvyZUZtH0nbQk7R5ci4NdfC+9GXVm3Dz/TlYVMN6Tv
r1UqC6KlEbh6Vm03PoK4boTheQMEAEZ2lZjAP3EYiG0yPeBRkeB6RE9Yf72a
suZdzGsyy6XLvQehfUJQeCL3/KKGxYUHA3deQEiX2HbOr+mlogFmHwOpgVWH
Tzaf52s9ZF6wLyLDnGx9MWE2YB0ryxcllwh7CX6K8ylBWqqwXIlpLuts7z2R
Mc4sJ85rSFhJYpxm7Vf3t4rNY6q1sjSQbpXxpIcccBJiEgw98Qie66ZYEwa2
+HgxYBrnQ5DCKZFO1YD2yfsTVASuXuc4HLBhyMRJIL+oOTDP7VLXQoVnYkMx
fgH6Snz4rTaFbXAwHR4UaEh4MJTftRkBMqccT5iJ6t02gTrZ3l+eYqWgFq++
10AMIYbO+qpNTjBaH1gxi8wZ1qZGZbU9triof5Bpw7y8XDqd7W9wdMyc4ZBy
xCe8FSie6RETYBbhUSidxsR+DnjqP0ri6grDqHeKU7EH0F30vodR/+WavCrt
yi8Hy7NOhP2EwKpLVKSndpqQr31jggoxYsjxlwb1voBzvrrrEBy4fOTat5N+
I97RNgO8m1hdcpmR+ELfu/nUxxGbvUsPR4vhwPsRUiTnD3/aemLUdUn7uEpk
PBqjhZAYXX3kVwoJrwDBIcoNPoV63dRGsUh5dHjE6agZ7it6oTCEJgF0KS+b
vPQhvGpn6LfE60YpasF5cv05cIpanvrGDHY48vB9SQ0amXwZNerSE4+M+nCh
4SILDnxvE4UCwFEPeQ3DAasol1QHd2tMPkOq/Cjk5tIDbDfv7eAppEiF4fD2
8ZGs8P8Q1+vfXMEXJ1jr/1iibXLjdF4mS5RFLyufrUGAXqUGxnZCfPeyeaRk
FKynPRKA5yJX5EGIfO18kQALwOzc/nOc9KQLXOhh7DaXKIr/NjUukdmjJyPC
pPnsL6ZuKxajG0iBRmG0g8OwjLwZNuKMAdLrnYWk1EgUDJThmlqd6R+Skgzc
awifHR3SS0HqO4HiEas1DDfj3LeZhvfkJN7iwYO/37T4xj4HRwhNtWZ1aZO0
UM62JfvF31mP2Mqo52ULz4vs2U0AsoZzX85z84bUWMij6fJFZMvHYnclEvVy
9qSPgA2ShWh/BXo/3fSa4Jf1aqJvlM9q5zyUZzK/qjLiyVcW0PWBl93qt/FW
CICQcQGxSbU3BTHYA1n85wojjmkcuIGXs7P768Co3AgNOehwn4WMVPvgthTR
4x4qQzEyPssA5MQLD6T0iRQcqElFeF7t4Shx2t51yoTtwKmIzScc0pQFL1mx
2/X0oK8Xhu5pREYyqtWyvO1NV2kON0t9QosUMyglSCeUVzDR+aZu5vxT0qDy
6eIi8HRNr3kMwT1hRkQ7bk5aZcsx5bff4p1N82bnZDUMhBQyurdrswQl2tsO
HiGtb6uvdT8SEMO+HJHKSxsPob3PH1sPbyvayzeVStyZfoPSHr9ao1i0vH+w
r8gSiPvIIHgzKxcWZu4OaXRh1wo5h1Z3jCLUX3rYfLAe39zz/aMGbFlGIaP5
5Cyu6XbJh+CUu4qSic1Ohtn/4VhVuR7JIOidM495DDQP3Fw8oTQGi3c/4jBL
3M+IDiyOAhxytfZ9U8RJVSfbTf18Eh5cTBjVr+6fLgOH6CHqMujK9Rv/C5+o
6OosJzl6BHgpH5lEZ3TGBSNd8zbLekYlq/HpYW2ZFuEWICgxOp12tgh+mSOQ
SJCk/EKReQl8BnIRHxZIq82A7BxRyRJF1BtNSdD1XqgsqL8eX2vwsvRrBPT2
dTTtL9xX8QMWT9cejkf4cVjKnAV0HqgP6TWhw2JXSKWlx4o+qi307cO3BBdy
jGpROt06HpQHmSNu1QoB8piZE5pJ1NMMUxNXKe48xlPqW339aSQ7CESJbUXU
0lL28/FjPmECvaSkIgNFyqHyTGSYGHQf6KOKDNnrC2xHKGc3wIuD1AhoAG3n
WwHCCCaW5TgVdwPa8FeC5RT19/uOvakXKfdHe1SsxEwXY2Z1SdsDJzeffGRt
uj8veL4qP1z37kO1z76WD/aqxaCDZeO3mZDUJF/G5Qnta1UjRDgTJTlq5TJj
eRAFGnN8FXq+4lrLn4ZqR/C5psO63ukwBK17xTdHL6EVmWpYgi8hfP/LbjKB
sjgO0zDmCZ104kWJoPy+lw98oLkwSR814uKyVChxmbUcRF2gINiqvhZBpE9F
aZ6/XtO+SSUb17AfLTDt1pPTXFtBCxHUZ0QbPmyWX/kcL/REyaSyGPqZo5me
KTxkRbRJJXfJTyvEIQ9HSa6PbBsF5MNK6re4HoeEB4Dg0sxxAI8HhKKxLCaZ
+WtDyeKjlQSWVNuhE3IxslIhe6DNvXZatzO9E36s2/WUkVYKJjBBoke8MSGp
vmSmT1KyCnR14qKL21cv2PCmG9OgqAW78RYcw2M1t30wy/SPCTf3OkHHUvh6
JzEVfa68aMaJ/JkvxxTfSkZ/Fb0EgSKNPJBLYrRooHSqCqC/gnGZXxXmdzDi
oFy0PZ2XuypAzlR60YePM2gdE01U3mWsRGLd05NOXlfV8n46bwHn/NaktVIz
06tWiOGdhvMFupR+2wtivB8sdRW3KR4SX1LXW2Q4E0U6Fekakf3TtuNMGRHs
moAAp4YAarRcMHwu01q0y8xxK3KpEWtf3IMlLD+aWonfyRpCxpjs1CMWBm1W
TRlzD4G2mZ5ri5+mKng4WfDZ36zH7R4GuM4J+5tuEMoVkCwaLpZWwYDwn9xx
jYxbx+Pny6Ck7vZ7ZSPODIsm9aZBrQaXcaAIsejjNll3ZLR5Qq51/VnkeDXH
bWz3vx3gOtdSX7GtlyZgzyxvqVgGHpRA/AAbAi4i8F7rieHwrU4mz+GpNv36
DiQiHZdvmswfEmB5NyYiekO7gOrkoTxGBZLa/IQ+EjOjNQvPuBZelCqkhIHh
ImdwNokdW0EMUYVNA2MrBCdngOA+FYl8nnhDU8hlz1xuTzIZ6aNMW2BV/jxR
mwigNRa8THuEkCle3+EKtV+ytw1XrJ4DCn9FodOi4+B4bDc2jd28Of/vCHnJ
ksPNgARz4ReHkl78LPOObzVlpT3Tfu0T2NiK32asZKXHWKIMqySVR2rt/KI5
CIriReqm5qkZt6IhONbZUeDEk2wpXJJXqh5+atyCwSzW16OW6RND7qTewU6p
1dOEwwZgFcbmwyMpyjogwDHRhaBYEWFOTFo2UsjaM0JSsDQPut8LON0Lr6cf
ZMrtUVqOMlhimNS6JcGoLr3ny7D+bOwWmApiF3f7t84CX6RfwjFZ0NH58/Vp
PQSkt6Kl1WrEK78m8D6k1yr0fmiCy5xNP/odgnOzYjVOuVD20Tj3+fLs4AHc
SpehHinLC4Eg0CLdffVQSiJMXpkpFpVRwikQ9l/GI4LcwYKxTlbglHD816wS
z2wRoYAJNd2sMOtzF/qLek/oGllm1naanhLXqUXdj1idUwzV2DwAVB9dbPKz
W/a9lbyw7K9Au0Ovve512KLAE57jII60w2RC7vfVwf/HCGqUN+agblfN2nWT
YGw2Dxsj24qTURvgJXzslvYH+I80/gBbe4UG8BL4YRi8HsWjUiNA2t9D/kwX
uHYwWP34kRL3v1zj0hMTcfSPBCFiK3ha3EpkuTa/UupzTJjAAZzjU3pgTCp3
SxlFxREDpdNs3Ox4V4XRZ0IOGtwaDz7MkfJTo0uNgc8I8wFkNBGwJ/2pz455
2E3GZphJoSXn1avKIk8r59GOIN0dg56qeVtyP5rCCbGemQY2rZaFDqF8LqYR
+fz1wre6M58mWq4U2szYpphX531lqivkiHybAIq9pIohbO/JWIbitl6kccWp
XRZWM3HkBm3gE7EEpvEHPI34Z2AKz0gSPZONkYq3YsgjQBpZl0Q2tUI3xJXQ
PX4h8+9GUHZ9Clu+0EN4kmeQJSkAB/X7sRIRGMmED+pY9KLxaRMovApHh7bV
V3DompaMoTRVmmftYstw2/+c1chyL4Ep2dpNuFYMEFhad+Bkf0AGFQrC70M9
4o95mdoxlgY2/IJ0orWAoItyGzoNf68X2XzZHBUfBj1iAZj3hSQWeSqVTLbk
49sDX/xvwNHRSfcBBlNoabIlBZacGkIak+sYZohDI69pRRF0f8zYbGLYfgWA
T597i8NB1Pdp7LFM0qoVuIeg2UanOFgB6ieqewitt0qUopHG7uXtGWKeNc2A
MCfp1QTPl6Q1vQF1Xo+ixBPnzM/0P7jkZujPJgMCFU7cK5F/lMSuTxN2OxPU
Dh3M8acenoFcqhJ6PLE1e/rnD7nmugzM4sUSH1KH8tBTm0Aw1ypCv+Lyq87I
ziQhb0soVafh80Zfff5NoZOUaBXkWYdE6IhK1XHCpzP43wMBe8uiuDaZcM58
hWuxZfzQCuyLqJ/TuZPzDvZKnr/b6tctlG4OimV7iwV2asxcPn0QUUdqLq6W
oUxPkEFCw0HEvkk+FUrkx9A3okkfcA8S6jgcyaoB8q7ZJB61F+KjkZNcH5Bj
X1INsL9ddJGNMsFW1sS88Po1ItE9twWWJ5aJrGXZlAtINTRRXc6obC3PcKBd
zzkxlmIZ+6oZ/e1uo6ZAbuMa8ht6fjT7POjUvLnYvg0VfVM/pF06+1jt/G14
pdU1Ti422YHwe9k0156VqDx9et3QH+DeaNFDlXEG6GVxuFipNDP1Pf5Kss9n
cI60e380tpB7/h35MSOwHW4brUkjGiCJso4P/T8krdzQ3zwLi0a8kGHaEIF3
dgCKNjzG7tEtY36CJuhkRY8nB1ZXf66iJnkdqMMVScP1hEYDs2m1QUHXxT4e
R66xWTdcllf41XFzka8hh0+21Ek2zlPnmNJ+ajr54TiAj38Fe7r6+L+vs2Wm
UjBWhFrtParhNS4GB2g48vNkwOENu4MhBhhwwtnbYuZSet//Qsa36l8PV3Fx
jwpG2DamvbbleOLScLhj+gRiz84eJmqVqigJ+cdEFrLAnB1FBD4KlIXPgXDn
PissZBIO5RCD/ABUoiE711UpzkP1cCe/h93+NYQBH7OtG9dRyj4bHRKqAiev
Op1I/+3qPQE6/ANe/3R7iQ3xgMD2aMPrtbFrO3yVggAiZhgYJDGfrDjlp+kH
BSOa9lcwkMly/TUvYYvRA6wp35yq1OxK+kHYABJEccoHL1SWaKs7OIYZJ7JI
ZhuRTI4v2q0KiPGUyOsb1grrzh7F8zL2vOYvpAmTdFWdqVJPO83GkW6oZSDO
EalBqOdWpfkN17a0hDGwQn7qzFg1kyFlxgDxDLjpnDLuJ8MDLkzsFGxpCHmo
+9VZECGcut6mn5/TD7sxYwR8qb2gsOa32Gtoz3/uT10unYboG26Nn3/F0p/y
KVQC3zWI+6yC73r1f8vqWUtBiAwF80ez5QCTJBBDxSMQ1A+dzPUoefUsg7hW
JwNX+U3oIv0zEpOhqNmp8jS9r8xbjiysSyOFwKcSbr0dAHrDRDb3wu07xzib
Mnw2kAK6qFxm7bSNMDpNxIJMeKMvgk4YkkyhvYYOiCf0HPoxjZGuoIZ+H4gH
ZhPTwAUmiJKmmeVBdXsNQIbfdOv/r7sZXpTnair7t8w65lyC+effg1LI0jXT
4fBTQAXb9snxwUCn2dSOQHmHbsz9YQ7f13ezZOjpXdCieySC2NLAsBCkEEJq
yLbuDBEj20IJI6C3j5+00TTGcQEW4sZIsV379osb/VLBUkMT95DEiFsZmuRE
Wc3fEu7tnm0NttJ6HkQrrGzOo65Oa070kmVwGJPp3iWX3cV9Y0xR7LUuTSRb
a47sLrHwBLRMdnztWf81X2qmeHPLZpRObltt8nx4WbWWxTkYhwu65qv2mHbq
atwMnHFhHrLDoAILBfRlrMYgLbP0quRJ/5fpa0FKCEogGVCvBD59sg4y1pJF
LkznbghzWuijHaKwYlLC64knZ4DnVhrdcXkpUTemQu0cRQp8OcsFrQm3zzb7
+J2yzyfFuk0p7E/id2huzbT4NHQvpom7QXpxVkTpmcz2+RAUE98l2GLOPazD
ZEuzGg5jKblcaEZUTK/4I6YzrmoLbNYBCGuhtqjmJ5htycoryZVdQX26xJrI
WvfM4oY6GfKWtKXR/ur64g0hFaqR+gt9GwZCxreZmilreBN39fwBFmS9woxu
ureEm/2RhlVYQFUaGBf53viOiPrP0Vr+ZGoqB5ZaquwVgsc4oqHVxgZ48FsN
wpB1C2e0j1+Egkz+Wef+8xvRaFYFHjh5jVdcyDO4qpssa7FOyNnhJ+ONNCuC
s1qxTEj2r+O1X+d3C00q6arpxrra1wNIZhjKxQRb0QRVRMUEzzUnuHseXiBk
OC51EZdIijLttetQXHw4/fkvNF5S7pyRX4s8ZaZCSmFWrDn+LDwjuF0gBK+l
Rss70zVS6vjqo6TFFYW8nNYkC3Jrt9oOVjCtoAUlXuHLz+IWbK35DlNn9MQA
2WMWqvR137aO6+tE2rvGTi2nBGI/WJUpGpCwJJwGAoQSLLlPyXNwDCh4u1Xg
HL5wpQvAt5eff0/XFFjXiWEs+CqY8wKzVzjMqfrC6lYsf+g+wOr8Nk20CGrm
NKKy18pIW6Dm8rN0a4sk8uVGFkFVlvyyyWdHmLrPmIOXuZ4cOcVRUguNLttr
HpZFkMEO+MPudghhGLlUHnaFsgADD/DlPY145PWyaFRKi0FT598Ha/hgPq/8
qcB5olxP3fC0nnIE6oKCNw4ZDBSTdqgNilOhSc7gkWd982Okg97zF4dsfXwc
VhSXoypYI86RIBEfBAYj/aBwO8xnRj45P7gAZv9Cf0++3khljv8DMKf3Il4g
3dT9sopyftlaKcA27pjhpoAER9GG35KkEoKhR9bct9QW2P0MQurx9cuWWxF5
7+f8f3WEmzQT7QpHem8PRijcYPf5aLFWvgUoueOO1kqxGf/pRftWoyR5MEe5
djc5WYSSbqHMsqyouQen7lcMCfZskgv89+s38Lyh3TfEKgXQgD0m/dIRKwO0
X5l2Y9qvtteqB+f5Q7KAJGSRAjxQ2AaDP8QElSYfLtqUs78f91nCbhkCVHqS
IIVXh4vicnJ1NCRLMK0poKTKNcp5W9XTYzimOeE/9age+LRvro/ucF+BxbdB
PVJjDyMtEmx7PYOsGrUqITDp3lKXCg9jCXQYB1BxaeCCWtUvy3lQHNTLeRZD
1t9EhgiBhdsY/d6qkqlRiQ9e2ktmPZSnecmIsgbffzu3NqgUxV5kfEjtCxHv
NZFZ0dJAUyY1kkNn9Nke52MskdRdZ0roUe6GMvPB4FRY9uRIPz5tlT1ycqtw
LfcBab0kQDJT1g8qEA4Uqr0k/co0/+dfJofzfw6cgxNBN8oJ9LikhtYwkHlc
CB1qBymgi0YAefI19mGyd/rEyfLdX4yLU6ayOXnPAPxEaA9bARnwUErTRpWu
36ulWtbwAhFq7kkYVyl4y5fjIVz2YWtsXMNwoSuwVgrnMMbkpPyygTN7P5rh
PNLR4l39+PAzqDRiThSeTxBg2aSGVvj5VhqTKhpDNfIk/+shqwn4tpxbtnLk
cS72mWke8bmyezSq3j/MoSd8fTikx3vVCSonGC735EfvmNOsXTimajn1ieT0
iScdLLPrMU8oL42LGlSHbiQrm+CgzPAdIlTP8lXs8YEsE/2VH8tWkHv+jIGV
iBTZNyjZEbK0XLkRBFk/SQqBy20RSu0Quj366aEsc8JEXTRr2nNWGfL141e3
1MQ0N7w32ePsUn0qFJFTPxovXATL7VJgfKu7gHA+V8A9Qx1fV6mS2Yhw3t8O
05cco5ldEV909MnmK+qc1XaAmoUpUmkJJXv9OT+Wujc1c95Y6OBkwISN4oDE
g1G54XZGt/KNsxot2TfyHcqecdKO3/UrIhlwVjKkqz3DTlSOwdunpOqyDjkM
vSnkyo9KS/5j6XNfDYdxM1vtn+YtHb5Q+pRjIge+0RTbrQbGJcZXlrlgfXEi
QYq3MsFVEWOMWeXRyPFyt1NaYMr2bQ+N4OfKnDM95y3MfnOA2ZGCmf/Fybc7
tnbylaC1wOIXh4Mjiha7vVUk/dKAbMVgCgIoDtuuZqO8YadxFxXNHzrO3c22
Nzgi4P6R4TITq/H8r40RLhicQ1Z8xS+tjSthnoWKkpPWoxNlZGvIEnmojQlH
RgqfOFZYZKHA1Rd+sEdndI2MHjNiKw3CV13TSfulfuiqBo8eARcca4Oou+vq
xqCnTsHOqxspXIO94ZsespbGLvaZjkPh8q/9JNDvQ5ptUNqafSVkeI0l9cI0
rqxXNoOKP+zAamEbVZJ/zaJcyjbNgE7kB0MJb22lgRWCXDXrHX+3RoGD6WhK
RHIjurRbfNXL8EiF81/5SH80mvZzfNX4dyWUifXKW7oNstnkffNjsqlE7crh
Wm99Njsre2/RgSR+eigQlJ5m3bxYNivfBi8/lu4TqK9R0YuQXfxXlAYRMUqD
9DNc+D1rk71AtuzON/u9CKKTCThbGK5xWO4A4YU6jOBRbu1xgok72J7LuyoG
Eh3P9g2/DfsVwPB7+44NK4Biie5I9aOOFDqr5bl/5uRTkhFS5G6O1FBXX38X
2aYcoe4BRPrXlhQ6+VUFKueybSqCuqMf707r1DS7c3rzcEpCxX1048qJgKlW
XS0qDC5BPCblB9X9Pd2oTb1AAgu0S0pHyq2IGYqQBl6YapQ1/7WG+lb0Ttso
z+iyEDwLe7fOU1BPRApkKDbq+EivKDhmY8DiNNoB5u11UVwDkMumWeiZb7lV
rFYuk3JYrr1Yvu78U+i088riczWHR/M6NpVyg/s8AGH1GwnZCPVXpBIPzXzG
EITE6y09S6O6uWLbOhkMOSgJ9jWvYT7pDAc3R5iOut/PyqWzjm/uBCPv0pAP
G+NQBaYchk3fkihRCvyQdoEiZ84vHCxLnc/bWBJ8SZiTg1uFvRsXGz/EcI+B
hXWVd2JcibaKPHRBioQFI5la9tvUoUHzxj+Q+/v6uBI/wYPrSSNQXmpp6F8s
BfsXCy2uRtCtNuQtVWgUtd/RYBaVLEBaXOM7bzo9qCQlh9bWjnX7NSYRnTR/
uUf/7z5omwwUbCIq0d6EZB6B7POACtJjbcSXk/MLvWyVnk4NJ5N1NLZ1Mry5
NbmJvxoy/PAlE+guxE7q+rZKnHFllrY/u1vXjIwvjRsJhCL9fG1eZNtYbPYK
am/0Wd4Jk7MzR5pVxAxNPtVcx7n3NDtSqiWgXsQAuBCOj5DJd+UvckBr9v8g
dtpxfvBZ9366n3IrSUvAjhC2FYPNBxV7bsLJlDzvy4JWRU1R4wKUUBqg2mKe
factyDkoQOhMr03ZTtow9rsRmLKuLIUdnBNR8yIWGMeLVHSLrFjyKerx4d7u
Z++juz8o32PJsI2jQTkCMKSOthEB8vvFpcFj9ECyspx37F2TH9Wnea8ds9Lr
H2VFEf6xrZ1UUVY8A0Td3QHM4LDhXn042nuTRzRgogFSf5W5k++VdO/hFgSh
zOhvQ9sf2axCE9q240XZwvf2yzlVPu85qYSdzrnFLwgxLEZtZp2ZF6P99Wtw
H03TXOXac40n7We159mB0yoeHY7CuRvYxg6/OA8liYELO/YiCaJoJA3f15m6
hKxQcXaySIWQssufCTDo6A+BT4aWs/YJm3JtqJ8soO7vIaqR+QYWfFoKIh9j
SDCZ2We9YEWyvANcwOamg7Kf1Ihk4JiQnHuAt/Air3pUZxSewbX2LTKpdal4
KalygyUvxq+jUPeb2gHR+laMvjw2DaaxhnU7wOE47hKOgJXqNJQ5ex9BquKu
1DkjKyRpg3FoWXpfYs+RAoHCtwXwX4gQzildLTBg1ruZuM44OBZTXIgEP+JU
UK0pD7LlBrrzRgxmrv06aXNbhZA+inVwKaSkiHCMpY7onesJE2wSEAys78JN
sMQKUJUAf8o0kjrFDjE6xY17pettvsQlBF/2M0eUCIu0ykbgmG5mEkUzYIDc
ydQWdbKqPOXPIzQqx6PSAKR780bEXXLbyCTeO+M1mQjTgKtBbvfMj9pdRA27
0TClYnobvWET6eh2E4/pvc9PsisN+w43SeHqqYY46s0XnlSKhGkjCrsUbmy9
LtXdgRc/6bjub0WhrnztwJQoxlteJE0TY+v34ATpdfrT9d+16cD68HecZrgA
1K1V8W83DBgcuA68xm+aooVc0l4eoYf+N6l1Fknj+LCXimniuBrjsEW+Xrgj
puxlXRXtaj/CRzAgjEA61Ghj+cA4wsp+YM6OFxvJtMdOb7KOazzFAK0Z8iYx
keOVT1ekBIHX4UgyVGZZEYVfblxv4xDuPKURZ57lnDa8r2dEs/FEAYDRYivo
04WzEI7fiDBf9xfnaBE3toHp1miQZdNNJCXyVjwLd6A5Iyl+yh0n39c/A0w/
MM7LJnsIJ10GoP0QSJhZ3GoM9PEKz+ASqIV0kWE/vlZdEOoMkmPbRWzVw0zR
l1SPUjKALrhAu5nu3hCgMHKtyED3/ywU4cHwH2aH/HH3XcczrE0uoHtF+E1b
5rP/CAh4dJLVwkNNUEMxAxGk3901kb193H9hw5lsf/hBxPAaixjIisomalMd
5nmKcmjSHandqfdjzC6Qz0aM2fmnyd6cuAOT8HxVN/IwxdknY1dRHsxDlntx
BmLdehca/cRxPSfF3leKdG0wGqOT1VUL7p84WBeeFeyvWkILDswjOc23GNNA
gpC2RCPyVZzSpvaC+m1e7CTdLL4F5/MAzWXovOGWZFhPp6cOm1v2nIVCfjP9
kB4QnDrxJD+wkziM+LLSjHWaQhDDsSYcJokDtCiS00lOkk0YQ/3TxOsXS/7m
zSoNIg1lFavQlhyXbR3mmlAtFcrL4dgZiOUdVwOGYU59abpUVbe8l062v6DJ
oJbcCzlBP73azaGwuS79RdOVGeu1woXvIyd90voenB93U2K+vU4p/x1T8Pi6
TfIcWAj7wXansLFTg3fL7QyeJN5g1GlwGbhtaimk786qEjiJJAZ7P1fAr+by
0iofMD9KjeinMKhHGBEgWo61YspmsHHaiz02aPoJHZOzby3V+i0DVzUM8kEf
SskkiG58vlH0X+R9vmHKrwTg4wKNuQWLrdNDR9CLdUByK58ihdh08eXPy+ex
R0mJCIZOuCIe9PYbcDDeAdVAn0zgWyOMJfjnXLESIMcovlaRx1dvVqPfVC1A
xxhKZINjBZX0PolYxOyZb2b1WE8Jia7PAEoLMAHLOgva5Li8fYJf4i70/Xuo
ASiOArh5+FThCl7abEr5HJdGg0DwCOGBkcDS5F25XMIQhG0KMddvAD6Oj65Y
6GebTGTlwzhQVZDqnUMXRXcaChfWawKQ1VtVnhbptH2pnW2SsTFRHzgTi2HV
1650zunlrI3lJL62I4JNkqATqdAOFztlUVLrd5tuirRRYU7Ccny9q+GPLDGx
GG/vuPKB3pzr6DL/XZKlM708bLJwB/brT7HzMdy99cxcYCMjlD2R9+/vIgf5
YpYv9FJYlQvPd075jQ8vS2HsBlKTDMRViikP8P3sadhOgm4gP1Y9eXEf/A1A
/0c22caxKt4p9yfSFMOlMs/Zu693cA154SizKhodWelcGmbv85BrMQlxdZiX
kKzLqwwSz99CG29LCo7MlGXbLed88mZ0runocMgvZM6XnTr95hFi2Q81i2kD
5fEeR9YdssvFo5F1ytv91tgkArWFNwc2ekwEZRSRg3TAnnMq55xqU6wNVAt9
ez/m6JwtmdsXQ2smpM5Xo5BmNabCm83zOx/5vMymwOAYsM4j0GjHg40KQfz2
W2I28DqrgsjOk/6En+SjKs4jvngdvQ3xukk0mggGMf+/M6swJaqkxEF/10ss
If1C13xITnE8PLcbICCaJCxFcpsC1LbfaAusq1WP9MD1KDCwPzphhMxM/zRf
tGPRy0723GnxZ0HB/J/67yAbNS4bBFSz0B10muQ3mvrROtWPoNN4knRptMX6
J6vxxNNLtQA02nYiBVDfxJiBIytScQDekrzhEVLcO44RyWJBdxi6JMmUq//7
VUujbnumO9hCBQJzvCtQdyPh5p+mgkGdxeYlWUcogm72U3HydlNpZWfSRNj4
ydTbyTtzfvNOhqvZEGfBW+dmsT+Lhlz/KTX3R2tMwnnvmFiRKU/YeRInD7Fw
5Am92ga/BdjoFlcFW/5ADHS75zEyc8jU8vVulw2sBIIkEqRj6I3Xi6NPcVqb
CHQUYyhVzxLMSjkSk776SNEQlMSBRpKJPXzDoVeIVR7L7YDzxeLd+GY/MIJ+
uAqneorYn1rK43daIomM+U1dY2G2lwIXLIOpVQON6ziS5yXCVgn3tmyEycbP
/YLMC+cIpXvg1sDjxj8gbiebSsevdMI5iAtSCDD6p8hR/SA5FKP4MgBoxDB8
BfVcF6C81xHSOYtQ1YZf5/UaQYY9fRcXd9THMnF6s0Q6CHOHYqvgq2KqOQgP
TS9ykCY/0xRHiufZbIBccS6mFB4fRJy09YKxL20aooxVVBPJjLQ+0SuXLa/y
yAjzEpnsX0E2mGI7iGoYazqIcln7rOsFaj4UJ3OlNo6nWyj5JnHDchrLYGEk
9tqJhfsSIxKT41l+Lr4nhXIwUAFenJClzBUDpue9oYa85JrNuQdIzaUPYXX4
C6Kmc4nHr5cKBE+R3LNYIWEvHnrTUsQFzu4nixOTG+OiNRNYr/ejUgElNH9a
9/kjst06FKjzh0j7QMiLVwi61azMBA2FoU+DgMVA6Bg0+PGiTSBhVS8qH8dc
sJOJWEf6RVMQxtnUM0yK19GNzqS29Cn7PWEAm+Hb/xR/2pfYuFXtlTNy7whm
t1izYq0umxro+M76i7Z7HS4UNVih8huFvHEokiAyFhyINgNePhQcf7tOayLf
vsGI/x5Ofqfm68Qcjlpw4hEghOZKXaBSPEl2uNFIoZx+3yogEYT6pFbRHqZ3
bDypoFZUfE1YWvDVoHbZdO0qAVjfkbpRDqgIZG8RPxZRlzOrRzzfrkaDkVoI
plOK6ONFDqvzM14NjgRl6G8IS6IbaagpjCDqeIbXNk8DDFxHQ/v6pQPJ7DB2
eKJ+lvs30hhlzVuGHk+OIIYb2zx+oVnGAuGqX1aBOH6bOrqtQgQp9kJZjXQ3
wOCKD2ZeTZ47YE0qFATLGCM6maODX9A31B1envnTBYlh2zzGjAiSxUJquU1y
7mozsBVNwIqwxRrq39ZPiKcoV9d3gCDa2FuYx8IVsqvi6wDUvJLhsQqse6Fb
Pw/jikvOUXwFvyTEOPbj6l6US0fqgvawzZ4vPMno6pzpSXq+iV8sXU0xw9WR
0Fio4xpJ5wj0YtlcKVrhfxm5G2NHNKEfof9elOPGwC5yzYNkY7RLf11TAin3
Ss4OTuGboZMwrgLlnARYUkA3HYSfriERmC9yDUCE5mr7D8u409XmcpdsLSgp
JsQjUDppHzvLzLZMHo3R64HeF3xoRGvjm5TuUi9NkaE9aEXn0pdB40jWAGu0
37MBHXBACUPBaEPjbPe9sMpEKKdKV299xrm25kflAIbqYnlWJF/cKCvz46u7
aveWYMdMbGFpLcMb3XjmY0GD5L2l54iTMJDw6lpqSq0M+iGQTocBpUJU2sHB
fzCkkaWkkVN2I5bNoLypQiR2KehL94OAz2jnGJY4bI+Ck20fn1FvMugIwHOD
KMkCF/JPyzXtwhHcwDdoKCgKznkq+nEkUrSBOm+g1qzgfNHdHK15c+oQfiR/
7UCFX/Te1zewqprJK1mN7RSN9ZBTudnLQ46p58pMfyS2KgDdFfk661myfZuT
XYDC6uHf1Auru6nsdneguaoYisMA5zppvyN05ztvXajNdbeP3pZXqwUb9Tkj
Uaute2NH/CzyziJYy/vQf2H+Yq3jM/HVHEOdiOQtF8eiyaP9KMTzklgTIYje
xzK1rQ0HYqZwhV9WcIxuJgoIJR97RpscvNp3vMhnlfkNj2WgFK3JtuIN3JSZ
NrJd5HkHarKp5A1+IRN/v7WBoMxwEumedQqRRmcCVaY5jRpYAD8nVZYiaCAz
oiSZyP9o0xmfbUkpG4DIfTVjZifpbi+HyU4tZbVshchF0LuwxFrBii9bcGHU
acpmKUsUrXY4rDb8u90NCDFj8Yy9tIXm1f3PEmucfl0FcJZEIEfRXodnm5hp
TDlcy8bX6AeZazJ5nepuN0eIll3uN3JsW/GpU67OrfjO/hZ1kpTU6eAuaaQ8
MyDnr9G8f9vAmRandFj+ySBWYA3xY0xJ91emJFvp0XSCuUDR8bvk0UreaPHE
lrxe2W/jCPywspm4znrIER3moTBz+h5r4LeNO9qSshnLKO+A3tBY/+MQZeTA
W3BSS51HrqCRGrmmNYG5g36CKxeEtfo8IrFyTvBpk0GVv55bb9CrjZ727Kpz
ITbCiDDZ3Fj7G0ks/Ntc9d4mcjQi0ac6TMO+K4nMAbyc1kRHhzyXQHxPGgLA
pCselN+TyHa7MuB7ng8a3bD9lJLPjy5vHuEU30hx1Ooy32A08h4n71ifQsls
qYEaxOOkILdaaImvghgta8G5pTf3p/PeHgyUztIERGICe9wW8EMmyTIpFgH+
NUmvNXA04qisoJXwhvglTykSp4DS1SM2H+YG2O2l2eJDfWx8bFAqpI4AfVgg
kdpfhH5VCuoAinXg0HVpykzvFe0PJpQkqhA/8thHc0VmMm6RlT2q2+YV9XSb
goOXH6yF5GRX3I3sf+5Pfms7ejC+a84th9Y8YACobMeihsNA+TlyERgOGAWd
GIamZ95C2Y5bDxNjBjuxkyIBJqxc1aY6JncaGIQPzsIqBBEJ9mUalYbC6xAn
sX8j7XCRT8+HCGdvyDXC2p378vLkwOsjoPl1wubG3TppG+FFicH3RGbLwOJ6
6XpqT2mq74MUFuLRwCs/WlF2/q/oxKo9EEsXAMlu0DQSO+83EaBSefR5eFgk
tr9jJivwAEfnKK+XyCJtOIIh3dt/SyLe8RMdZLxWok9xWwwk7JqM7LMpHLfg
8n6xGp9ERm5c2qgg2QAhgX/ThugYzwFU2okBsUB14f8fgObmsRRbmkFarmWJ
tpd6G6HQ4TR51bJM2DOH9c7FsUaCOvj4QJJuGTed6KkKBmmqTK77PRQo21yy
/ytd9SiGvmqDVR88vPng7Pa4cpSioyWggNT+9mKjInNk03KUm62m3ThZgxGn
aeM6jPY09eZTT9mt3+VK59r1P2U9FR2MG318Y+hA5Eue/cQCMNg0CniYKWEL
Q4iWgKWW3CiWYNOEfBe7799UdC9AMESOzLGfqr+VN/ZIc+86qcgSxjAOuUI5
pW4EfxPQK5s987haEEgYnBqZbyu960tmXArkwGCu4Key5Q/PEY4j3M2ZCUQ9
SheT+OCiEPbncX1Ud8wwHg4ex9ec+x8hbawDVGcR7ZfnF98NoDKlKlhRBeEJ
hJ1zW0rAf+RUFnoxnOCDaXL3vSRnK0B3M5CRfE1r1an9+QldFxxLWkHUeDvN
100/ehuu2CDgVS3q+DXYjYKuVCAdsmAvDTs0Rbo7Jf7AeAOvO0Um50W8UYKV
JFKFxbGIsx3qwV/MWr55vefU+bJxTFVE9Gof7W6yZXijJEHXYCKwnjxSu7cA
3HML5CHWP7Pw1RSIAkuy1XaL50MPEJ7iYvmNkkS5seWjf+OHVR46TtktS7ld
v4gg/OZUqfQxXv2QgZcMCpwa+WwVbwyjDEpTCf7l6xAWRBaHs5aA//u/cOZ7
0bPMTYZHEwwAjlCc9jqI5c3CHlKaGbYVR4LyEMHdlQ/UlO5Q0W5zVLZCNVo2
VoKpFR1sn9rCnV8GE15tlesPoONnovmN1Z53uz2Kk/lj7ufO5sxCTudqUfz5
l53lqT6K8/bpTdcLep+8zdiluJHQECsB/fubBLz5c6aHBjC8XWtYGmarla1Z
Sa2IK6zDygzetXH0jdNN/2pTp4wUK9KVadU2H1nC5LjQHNzuwEQq75BHAD/o
MgLNhKKXaTMvY9/J5X/6cLLOJ/sRh8ep8apDTqV7WaS2Y7w2CgNsTXyZXIch
7t2T6KcFlNDSYJ7LpJyAb0SbgICykf6gBmJtI/+PQSan78OiYGFZlYYBvm0n
QIC/CZE3fQyYANR6ylzFVsDWiQ4awv8u+SNm+8fjtbrDL3dgGpRWo9NxL1lL
lv+flGfHZgzI5rg8WhUS3uK3TXzVNyhGALyetvV1yGWr8S9m2sHVb4S0yYwC
Eq2NknTLQOMbC1VFXZfqDVhY1N8PINIG4QTx4gQr4EcvgYQqZPaUKl//rNUv
d9tKKg4vNR7smDz50TPilpmOs/KvT6GFNGAGHAHthyw/0ROMIL7bfRWmgoib
Dbnk9zCZynRF+mZdj7+bpyL38m6AiE0k5PRzuz2g+CvFL9RKUgqtCo8H4BFT
Xm5W0uzxGU9oBGw78ouQMEbl0NFt6yOZk3R1m5tbAUJ/ZIcSzaR2E0G3DJ44
vMiT7fNNgLM7c6YHLNqGxZd7+ri+N8waGhUYuEdKDCFm+MVRBrZSi/gHqKEt
Rm6918HmhAWcHuO+RKnCskQ/06SVNUbAvftfhTQss8//mPbHdyOs/JlzsDLU
HvSlKIdk+cYAfIaV2nXB2Mli4ypp3R2VruK4VN1TguCqps3c4AubDgPUnFdk
PbDMYs8dOEnk7LpD+W72lUwbZ9NyXrzbAjv616zfOTVEu6Kab7wSVoraAPLi
QfCHfqcF3Jx6SMCjKa0JatJSD+wRkhDTKtBq9TKAsAvRQ/UxaANtKUQocTk+
8gYveW6KfRfCesTB8ciyPOJM6mpzWPNdHjGtDCWDf5pCJbA1xOj3wCtY/uJD
ElmsX1vX4a6IUEXapz6fWHLmFdwRsQXDgW7GrGlAeWHSluUY0BDFbSDZRzkX
3m1SYsXtS1JJTaRb83G51q8YYPgvQqWVj7orVNfr5gQH6EgqEvWaduPpLL4J
jrxIruNhTs0cuyZw5k7w0Gqnirnb+xgxvAtPor3vB2P4Vf0tkxz99cNy1ZWB
9NhfqZ9G/EC6GnPFe/S19RXPuIejNCOJd5YwETDvZdg2zT0CtKZK7grDPcLy
ERdDwaEWP632UxxSIz6AFR5Z802iHMvZxvlFWXY+CHqIaKCGuWWQ1/LTEW1v
cnmgPaWlU6YGYn7Sp14IDmsCMl+e79vrHFkpBLcOBZbvbMSffpHGvBWtaRS1
QbnZ4LbhHqjv+kwCzJ18tLC1Ec6krIvFemtLcNqLPimbytGMc5G7LIvxzhOh
9wJbn7k0mF12OJLcV7bbYajcD07FoJ0T4JIgdoQvDuhY5cm3cnftQaKdXFnm
6q9nD4F1x57rV/SPKptMk7necrSNt50SCJEJCPgtJWDTHOUDZq3F0GlhhWXL
KOh0mtUr7YdMemt409yXB1GiTrHi50DV6QAUw5XbIqp1cvivlRsNzE2xbXmi
TRyEj0phlbpGK+H0ypa63VIvvtqEZyU6BEzojFjhDxbQ8PcxnjZDiSgD3z9X
TFLmImaRygySmQwM7vDj/mClXVIckVg6OnDwbFz/1+WLXay1u2BkCNwMUqtt
j3TUXPl+j98mOCLY2FmRPVE2BTbAmOJbDOHBgXrJta64dTTqO/O0VSTqr6JB
U9GOVluDNDrIL9gowb8mD1Up/0iPF4H6LEJUpCif1hli3WRYkPdDeXOJwau2
yAk2oOYNdDns3Pqxgv/2yrfDF1ROTE+B4GdEoPCAIoPQwVqxTcXoYvGp3DZy
W7MMRYJj3VlXPXEJ1rGl/8k55lRPR02la7nRa/cHX3x6ocJRG+X/ZHEznIHe
zQXG6cFQNx11LsQQCVuTlxkYKUsuUt+N/UP6lVPflmYH3TpyqdMR1G074HhL
wj7YFYiWURud6drAviZDgWiNTtJa0/GfJHswPRqh0pIeWeeUVZ3f0NKhuRrV
87IQmKQCcJFArWFQ/OCanzl+jTyWeibyMonQGefuIPi3OV9oO67lrnsv9lIM
aonqvNwGOSHVDDuGnoTXHsPLiyIFMoZJeLqPWgGib8AbUY+9SG5aSl395Uw5
FlajETTB0VImWLDayPinO/n72s57SbDh3UsJe+bsAOu3GE1liUNxbWghbqpu
qNYEo8gcdfyaCgvrrwCqs8TstG2U2wQ5MhLmkrl+Eq0cHfZ3ThDzC01lk0NI
5gZm4YvzUBugT16z+/rN4Dxygn+mt3dOJMwa7kdH3+dk62imXUV9r1GGzU6Y
q1/68ZjyGtmRwQN8P5yYLgJAHIZOzkSVB04UIitmEMVr8Hayr5q+rxgv9pQN
kh35LGFA3SYZ3zTv4vhWRy1WHBt0uYd3vGnTc2NLCNC1/0IRl9aZd+GlxNi9
9uf53n1VBIBZO8g1K39juEsAiLoHu3or96SAtAcNVbkOuUIYZ7rYzkXCQVJG
/dWXX1O/BPXug6Irk0PjENMWyTN6hiX3F6AkXHsmrg0dpoJGVcZvG8dWmwal
8XqaVEt3HUdru8Vl89jKhy848DY8e0m+Wy9oAaniJymh57uaMFjSdZNg97Wu
MDj+UHVBx74xEonoNlr3fugmKYqa8yWhd0WDBSxGuF8ACp4Dth+E1T0gAGTG
F47hAChGMpZ58cdeqRg0jQ+GUJAsUmNmn6JDdq1sl2KDVBM/TyyrfUYv/NyE
Z5vgAQmFisil9RBx7etVKisPS1j8IQ5UhqCeqyszZar9UTorWItxCQX9f2n+
hGmiCnbm8X+4Gosxtb44X0kinh0uk2s8MnL4e53BVGik0/GRwwhesBiORZnK
TdO8YHzohwkqHUycHOmp68i33TBLRMuY7jh8CkZ1JzBYoqrIMpUGeME6YOSu
Z5NJlN+FASU/XaPDsaEYABsaf38mGl27LGMb6pu965onu8OqX8ZA3BqVQypE
S9o7kMsahxq5TwJRjDuyXLp8TJsQf/SCaloHLdUNn7fygeIEuuc1u/8QhWg3
uS8wNqNBDIbUjTDObNniBzz4MXizQjWjgBpG3y1DUh89F1UnHXdyKAURD6R9
phlwOj9Tc8tKZ2krAEdcv72i5nUuMcqC3kTIXzMKpOCkDNFlTC2VYlh4e+6U
ZGafAumFPIyDZbg6/e+3tmRGNDAD9MBQxGR9QQxkwc9Ejmlbt2lx7cKJe5ZI
F2MwqOLzDcLY4cXOQiKje2SDRYn04PlINc4PIST7y56ULFUvmISNTqgSHqjO
Y47mH492XKxUy3j73kmRcfYOEx9TdQ0HPQIzZgBq3CzY9iLWHBc0UVn/awR1
OFs8OL8nvloE3Q+2ObdpDmqr7glMs6CAKXScQ6uBvTbm1fz9X4UY/zk3mo+r
dFWCcARwbNKuZrWC5BWP5RubF65GyOkW4Dfl8Bat1UKEJWsYuZ3hXwSwC1yi
zUuW501HXT2vqb6sarIaenZuji4vu5a2AP5hwVxiy8gEyh3fTYhI4mGJ59GM
Hb/obN4CnuA8LntBg2tHmYazaZ2bJ/nVDwFRz+5GOoN0qA7zXtd7SL3TALo3
ZayVjQll1om+ym3WX/uPZbROcKAO5a+RPvGwp5HGdcbcxLaEHOdqvG4tnqCC
MOTWNyPuiXmgyN6wcpY2Tz7IrVr7uQRd6bE5k5V3vjtRbi3X3/6corkxza1m
iATVqbnkArpOXwJFBkzHEWxfmAnoLVysxwuyq2MDLwA7lIMs/lXA0SeUyPMK
Ls233siJcr/6wqc7IVpA27/kBkuDgx6w7ZPKnyETGltJlIqLYDxV2yJL8g5l
Ak8ycpsNBCUoqugf9H0f9AyToVYq9wy73tqm+iItXYdVL+aDZ9F0ivkl66v6
+GU2vKV7t8fJaN20Dw9aq1aO93Z4pALhdehGgO7bhV8ghtKLs9cjLVYIGQkG
itKByJSwqLx5p/HB7r+lIn906YUHF6PJXYoFwbEYCkxaejmo2erTbTW94E3J
Ixf8i26DPs0KOWUomgRwi00ZZ5SyAS6TmO8FKcjgvtc8tx+w1qSWwmeawqUv
FqbeSe3HXoBPVnjWMX1PlcuAHSUY3VixBCXznuIGxZswzMYq0reP91/MGn/v
/cS+oEfoen+yXaMowDdDt1PUU0iTaGyJ1yqdKYf0lodvOY6sHe/jrUNTwU+Y
vjfgQ6Q7JfUJO1puGfvAITgayNQZ5dGNqrRQV0TcOutFYmUVvCqzl1I+BKGz
q1MNSxCursv5/CSt3p1gf5PoSC5rSZVzcdi0A/LxxMoLERilHOQqvLNpstR0
Ja8sy0srqFuf3mLB0p6FBUn5NlN48Z1fTXgFAAJ4ibRORZEs8fODKJIdNXYt
xV7R+ogYGJDBu4KcLZ8CSS7LhN2XLPH+nX2a/FpHHkMbAwjOLDPEDBj/6SIW
xyeSZclU4SGeZC99RGDVWRu/+PZx94Yi9Kg1EKn1yTbJ8oTcp09g46bPbWDM
5ZTF6QR+YYO0dDxx+WrhsnF7VVJ2/njzO0hZft/9JHgPmxqkYrnNRkkZfFKf
zQq64TCyvrxtWIxfvJwamBpjG98c1kwg4gMmHCY/8FZvn1ikmZa4woGVKTfH
XsfKU5WU9luWkCcNyEyvGPkiWCnqQ3HJMl8/cdxQKCo8XXehXZTHXmgg3y3f
811sKkArWPGah7U6rCQ0s/NO/nx4nJ23izhpAZjj35a+BYRMJowmYiEJyjSC
CQejfNqxpMD4GJ40BNp/6qiYbhJ2WAgRKNN82DR19r3wtl4CwURNli2Ly3qq
y+UJcKBOK7qDVz5Yd4RG3T680II0qHCgoUaSGQa9Zs0/a3SvQhBY5Q9jFyLl
FbQtsr+Y+2XV0HrGnT6pE/jgAUFC+KjdSYg+qiIbr++ksi3TjWbekYSNYD6B
vAazDMjsryAE9Ao7FaNRcMb+ZG/gtjLlkX9ukWhWI4m72wSqFaSBU1rZWdqR
0zcYp5omN/xMjlANOF56H3q90t7VPGOoW5R4EfGcsR351+LXNs3AjEIq4GHf
fxJcjzET44hjoDBJ/7znGKyYwvoxqd6JKNw1+QJC1Ee8zaRFfPMFMZ7+cPf7
UD4QoRtyj539cuxXf4JzdF/iwRvGTbT1v/KQ+cPA/fiuRkoZzVWzbSr9fNxO
BFN6oU4xgaXevZ0Qby18BVju1hc8LivWAGROJCOkPoXMeNaVTGaU/0aQeg6L
PeIcYxKqXlR4vwCOUSFXsjQ0OdVeAYVjQKSlcq1l95eNOSLEJcuSnAx0JaFD
axDW1spy9fQw/nqnBZnAMoBxstVEqdVte/5FgWGDaSRlsI9OEa8cfQxkoLyO
7YKHKO0epr2reMVrI9DJFdqGUSZZ40hZEw01R4ekRiGpKqnzeZL/1tzNVLha
D4moU3ocFNckk2eFIq/q6WluSlLhN8/PA3pRvRRN1/TA4xUakF32dyoPMVZH
n9uoIh6CyG7kWgHUJ9dCW2KqERZf4esF8i2Y/gTlq+nouZWmRV6TpZJdiovT
wQwZMPzves/44k9yNslOzMp5Pz8h5+WC7IKk0O0O5+tbH642I4kSnxHNThkW
AdRCoAnIm93I0W1Wf5duscsUi4gWqF7rJipuDjrUvLGnA3BMtXyfSV+V9KhY
GojuocvyhWJecONHyvA0cvRJMp1c0TsrI27tnAeA748kUjlFnSPHwHwZuevR
27nL5jeo7SSv9+FxkQ0cUXeP3F5P6K4zfpbwHcZxAvctIjiGer6NjSjFLMdP
b4VA8+6kkClqJcuAFP9yZECrVaYXEihHcxHNNxVzx40XsReUElv1CMxmL2h2
XWSlcYJE3hZgbbGkneN2ZmZFNR3n863l+GvN8dWNR5SG7Ft0U1dPvZBIrwqd
prO7zvYN0kLkKBHROmWgxA6agUfkKId331ZTeNRfQP0M5d0TF9b0se/lxM5J
XlSk1SY+vEokpHrxMTlMDIhgzbwRg0vq0Qv8y7evvsGHJMX45G54gW4ti8G4
KAm1fjnicvnZ8tO2BWJCAv0pQJLg5tb1HVWjXL716sQzad4n3L5tLT1X0WEf
YVe4vW8BNSkMz+7TsNLvN1qzpP1AEmVZJTBl3epcGzS/7JmZru45YjJF7cI5
aN/51dpxT1nMNquPDyuMxlFtZXbwrgDUPX8MCsPOsGPhnWt3IEcYFvwxVzY4
tDh8+zW2gOue045JbPBJQmXZL0vAGpm5Uxf2mZg5k3sANIy+pCCZZweLrspf
YHFHZpr0YTDHyKuP+Aqblrs785JbA8Ig2fHBxUHtsImYKSBsscUeWddAHam4
I7bWwW8rZWA4ok2aR+7sv4SDZ/XTZMI9LmXChGAyIXQ4juBUb+OgMS4cKOnb
et36s2R4A2/Tr3kgYm2maJU/I57cpk6pgX0Bn1laZS6Y+rEKMqDwzRhRdoyt
s8UW0f2O60KGRK9iHpWZuO+5fltYLI7hYgTScjdKnXZgHzcXBNwuQRURLT5r
g/ZBWRDNDj9AY4yoZR8aZ6OD7HhdJ3/MKWoPxp5bgytY44mpc5hJ4iHGJzXh
XkaQi5bk4IKg1VNWD1yGUG9xH4d2I7iyFcBsb6qa5LtGkg3Bvp0fhrTnvgJS
66LgOScSmMgi4/DiKSs8P3VT4eFqZy8aMO9YGC1oJxFHnYxQV+/Iivp2CBQm
TOBfRJMp1WWoug4zWxKEopZEH8/lLrhdj3dVawQ5qc6iCQFeW8hkkvs7LX/I
dBxNuDJU19dknQQnef+aP0kj8RTfofm1loLUPO0EaLxkf9wHI7NEYuh2JlQA
g3Kp4UMZ1Fde7x4SoNWBfyZ7RWxENg3xBQrG+bW3rbWoZdgLxPvpcu4VOEAs
oCic/lv0vbklIp7q0FTmlMqx2IaAwX64R2/8uXYSvhNwIKLdXxbeg7tyZP45
aMVNUHcF0C6zKvjVeqhzXN6fUh4t0M+Fg4QSeosd2XrgdOWgPKEBWnYp9NUX
1R46lj9x2QwNbPJhq1g+smXOGgmgI1tj7832qSiOgcCvd8n1w+do/hKqfieU
/xJc9/+5/rJFQ1hww0di2ZOTRfvoyNPEu6e+aNZEu6LECiV9zjAYvEfBPysP
8i4CFIic01PgW0xe8bDzecr3JF+iXJb/70OFYrbNMyMQh1yWbF7AgwU+5KoC
V2RyaBpi8DTOH/Xcd8iLw7f9mSYFwP2xiUdZHtr4EtphmJxPCsbarnCg0pjs
LeJ4nm7KGSC5SJj3I/kJBPi1L1pwQ6wmYPxfvIGubOMNHzwvCCmSqD5sVMYQ
em3ZaN92u8KYadKk75Hrr4nL7hDKF7gRg8YcXyAs7aNyE6lFuTy9KEtaiGji
X+PiRJf4pRcRZQB/gpEardtNSylRh/PDkSoKp6OQSwJ4shGcMEi7xDZcIyxK
EFpLhU4gg4L8UhlbmZJnoSpYXJ8ukygC6At55NcKBc29ghPowhYWE0o+Yzkr
Uo4ovcrDbRwqGvxxEjn66DKJ6i9Zd7ekJSxWUbwZwRnyql3fIWvMr6qbVb0L
ILMe8+d02uCyaMhCujLJhtVeDxbqD2IfCqgo+EMlfjEFm/Op/YmD8a7kwJeD
qzgGN97pET3jnA0nJJA7eihlJVkt1oJUR80XImTrbg+K1Tv0xM0pq2D2vXNd
VY9ah2AB3FU/M5XyvJyqQkY0WVuzMfL/P64Oc8JzRqaVOY2QtRpqRxbjO5IK
XvJ8Ldckla/qReQioljEsUBNFELjLC86VgCaYIWGR2OuwbKTJlul1ReErr5D
VQlloxqcdP2yq69CSCFtwp/t+tKOsDSXpRvNwGVuYVAGtoNoCbrYWPJDWzIZ
BezUAH1iOBMpYEZB7Al+POwT73eqfiLd61RLKDB1pIF2i2Xf2kgBprvJC0Id
FEVPxXV7C7/PYpWdPDCwHHBuwf+y5VoIeZkyN9k4u8MSwMqzbkNLgMclOA8I
oUCGrFh13KRAne1TL/eQ641Sj1P44GGhhQPYIkQfkeZyKsHVPGp+ItJJ1rHV
7OlRnBQua9cviZICh6NMPOA+RRVJfcDTccT2V43eZviKCfv4CVeo2n0itUxF
BGUHZcyfS6dxQO6vWkKackPxrwBLt4SJqprZiL6r0VmNIU0S8GZkMT3v6/te
HxF0YdnSlwh5GmfM9fHYvtKK091aL+HeRfZ3QcF1YzpfZ9+fHVN+p5QhmDrF
yaQnXcsdlVcn6DlH4UWC+suOLVjsggpoQTTjylgTjjCX4R7e+ZVllboHlsqE
vH+TgWnNdvMPLuk3fzeWvROuBiprp13vhOCB1yjjAAL/hZ8ZhX220xpfuQAv
RH/Tggc45DEkSn3hRWt22IOpmEUAWUyQKNWzogIw5R8SEBLrba4jMWbKyrgz
Z/ybxEz64cD4R5fZI8I90rxICgxSH+yOYCQHifrVHyFadMOkbZnEwVUrTTx/
CjwFvF3+xK7rbn4PmD+Pu/D++19eerBpLFhVmg5D88puJGXhzje3KkFnZb/g
cdVwv8NBLevTp7N7pWboH3PJ03lF+dNdppyrafWWqNSV0OzoHgR4KLWAeCy1
wPjnq6p66kSLGinXFqRrUmu2vZ9jw96rrx8Oy+5BkNdqPyVFJpDsut/4+qjb
+kNwnxLljLQLFobRQByvvj1DiUCb0WjFp/Dhmuon694UfCkJXBk0hMC6ttai
4gi+ZDhKCvDjwKi39wQrC421ya1sRqlSfnJX9ge3RZcjsvEXPdfdZ3DwuD3p
YERa5gqgKM5QxRqS1ocsxmXe1VHpGRaakzYxOeRReBbBUHp3DZGJ2wqkweRQ
7GR3G8ljE1yZGUFUKG0AzRSOsnPLVz+sWRGdITl5JKz8wA3L+HxvRlqJKpz9
7KEnVD8IETMyiN54l8C6O+8xW5N5NxGu8Ba8/Fp8USjACzi6uVZHHa5BN8/F
+Zg355M8CmkrVPvA/YUiBkjuqKdYutX1V2B65WfI3YmUGuwK/FCS5lVJQ6dL
my7mY2ZMpbYEnyTi+hmxGUeS1O0NXDpvbqcJbbYkmJQ04O1g+vyg7apFFjDd
tyMRDS+m/bEvD9x7g4pMsePtW3DVExxJ2BFJe2+MkkMSZc9X00tjg1oxYtAn
WYQvP2luWKDX5rEk1+iRTE3S7DVayNFyjJAfl47lY4G9h7KGukrE0GEQE+Zb
YH/wxTM0ut5znrN8BWe9tA5lCAlrGcoEL+ok1XrAzF4luTcAT9Xdxvn+M5lg
cCP9+XzYCFTb9uQ1EeDRsTGTRG46exTZ9Th7lvWcH8f6xbg682IkTuEpvDvx
zNygsAMm+JVHPW4LbJCfpaHjCAWP7AwpCeqymJK+ji+bwev2YjXq3rLG2cH9
zEIfVdwj3GY4B04U9fPbt/ol4wIJbNLwKSBGc8TdtvY5Ur2mMroGEEUi9eJv
kU0zeRtzXt06N4ywSG2dZamqViU+2kG714UsiAGsF9l2GfiHMYC36hEUKeET
Bht3XOCLaILj6dx9HBlOOTcFxqNQpqtCVXTEZ0V0vgS45LklYxtK0+tC81NQ
E/ZIEab/RZgZnbrMj3XVr8PvyiqM7ByGIzP+YwwewkB0ZIEnIKBrMPTFAdNy
ceDGv+lJepNbNEQsnTNtvcHyZxji46FYtLP0Kojrx16YU70pumJGz+bxV6+F
cNjN2oYO+7jz8XlFHmDYy+ymEmzb+LhPxRsu4sWmfqtPeFq6y4Psa55JdWFQ
5Z3AEqKmeJS0nkQ2PXCwxl4CT6W9b0it6sYfFSrGrh2syKj9oksiODexpizt
j+Cb4N068ZXrahUKBHfsCSXHe/Bwvn7BDPY7jiWx0qFoZrpTkJ0T5bf9RTdX
yrLTbvSHQuzyrMrq0g6Dvd+9Bf12EkBzWlAYgTncQtWaZZCzqJNF4x30vG5W
zaTDRwidgJHpbKaJAMyL1ArwonnvE8OxxsRYc28CvifNV0Aw+FHtoJNjRpm3
auzcxMrgypw21fvQBIH3+2w5E0XZeyQPYUJheO9C2hU5mAfrmleShj70RpiP
vxKFOPQqastEiC5jZjaSTT/DEroiBIeNvPNQUHD/7OeI7J+Uy/T20fBiQbdg
+uQndHIijnXUyA3XTeZv+CMNMzl/PcQ/2ObGqpRWnrCq1tVchHbVgA+duE+c
d1lQsJosLNQr+bBE7zwqI88Drwd8BQOQMpqIFlht29qxfglllqHA/70yMTl0
T6gg1oWGt4U8f7ko7rES5ZcIOCi01vMx0rQecdyPwOaI+OCqqPh2G/52Rc4c
MXUK4G33HRFoWJ6h+t53SuN0fiTP8kjoLIcmkJHmuLNyXPUZrothvIf9U8a2
fKebrEV0yVWHVCsfV+95PKLrk703MKXV+3Mx2qEf1JVJV40nQpAfHSr8KhGh
+1F7t6B2ZDKwkyrQyIHGnE3eqX0o0OqPqM/Yxj024ziTHqL7pZaQqe6Qifhw
vOTT0ahaga+Hkq7J870EKPLZJgR1O/mRx3IR6Ugn4HiQ7iASMNSdHQbuNZYh
l/dxgYdktIOHmE5HQE7hZqLeCUvEOU6Z5ivIFknbqqp+izGPmY1qUup76YAl
ik36Lj6tZzkGEdMCvM+2C+2BkrYbKAk9N8ZnXh4262oyfN0lQ8H0mlWCAgc4
756z4iN/WIop486vZfBgMP359Yu6K1dSn2rBEKVM7ksf8YZkmZlCFQPtnRWq
7gpLizPA4tmG6xjlMnVUcnLR7VVKIjms1SMwhUefOsBMqELpMzhpX/xkp2XG
eHUNlRz29DldhKAtR7onHjAovkes+ffCbkvhpGJW0hgv2I6d07FuqoVeT0Xl
L5pkazE4DsabLAAoTtsx/qMUdwrVoIXPSGiWpiMGmjRvWkyv3vaK0+YXAh14
vcId4t4mtaHrZXNkL/P9fNRNyUQwZq/6IpjcNfgZApntCjleQM5MUfVPkF7p
0cT6XbOybV/AHyw3poQRfh0meekh6k58jKA3QXs1vVdM9V3mQ/bj2sciZqE3
V+yRL9+iIryaTi6hCUARPPxnzfrvPKmuGcWfpvRmnD40U9wDcK0TmUyg4+Xf
u/HV3FdT/KejOSklGeni+3AYRbnZVjiz7x+ILAOy6NIDAefZ4HNbewvZRXzX
0qiGavEtr/IlyOfVkzybp18DidH8StJW9qWJRlwCzgPi5WsEcQr/5T6BJMgT
qpNL/ATN8Mf3fa86a5w7h3AoZBS8SBj8Z4EHLWEhDiQyuB2rMhDwxEHKbUcu
DiWliwrvLI3JFof9AjyAOMdT+klLsLvCr3a9xGxaiJvlvbv76KfQo4/nez2m
9vfFbGbgbUsT/WRW0Ad5DKUdWPWaF/85mX0tUwvWX6Ps7xSLY83hbQy01V+m
+1hGU1kFNsK7v3UjrlxIMu3GCFU7Pairmj/cJmr2Xnx6YNIzAC4UA3BUTSod
YAMvJyytHCUpPOX8s5o97tZ0wI0o5GgBBidUyC2+dDaOcJu0FYf1LM6G09gJ
riodUny8r+OJgyhNgRvoAEuoxEYt19l5fRGV+NQaxd4yf8s9H6gSV67Hu4BT
AEjgvMYROCg0BjqAXkZZrBrWMY97IktYlkmZ1rTsceBhYzhDAFWK9OtYcbno
FxLwGcjiNSSnUA3f/1eD91us1Tbze1NgBXuRBgPhyEUoaDNS+FZJXeKyn6KF
/dBQlG7XryMk180LrCnTdnzsA3f+kfFvpfxS3ra8sh1hx2pgsAkJVvkQE9R7
AK5O69jFdzXdYmpIxKSJkR1jgNP+Z3mCEtgebCXgwyxUbijF8WNitowzi2Wj
mu/bgsnKEipSdIiqecjpAgEhvEqyclVO4H/PM5ACN+olml2NnN2fvzLsfM6Q
lqNHDvUKFIsfCyw7GUipVuvmADXeuUWnixlHyuA8ojfAcsjkSaOfTiLO5lvc
YU8Own8mhdnU1lyLdYsQ3yGcGasHcd4d9aQBG+U0xSG3n+bqVcmG/+aFUbP2
45x6+BYjX5wWE8Ixix3ST3H1uaNnzvNeChZL/di7j20qgIA3wmmfCSmaeByx
goOse1ppbNS+CFe+rZl0c9ELDdJAoByyWY+e94zQdI7pVCyvbYpJaIhEBn9H
lFL4L1O6YUWA4pPacSG3WnDzHjR6JokwQGK85vIsuF4N2UOnxpExQsKwYrOa
1Mp4W9XK53GPFnCkzayUNLgzBCzEUoWeQXA4h0h5knW3Eb6O9BIiI8dBIZB6
pDdMnY78LiFyA+RD+gD72UKFZgb9YcQPBsX9k93xYrXWLLgqaO7CFd/SK0sb
PNfC/DoTxsV3fwbGymr+W87UroaKYOMHsldq2St1jHkBv569wAQwivcKSBxx
cqiPHkFcrdOUKaQ+m5h13f/RkHrx5vFlbt66X6gI5nyNyws4/97aw4Z/9dDI
1ja7SuahyXQ2PmIK/y6t2Z7toB5dPpw3HHbC/8qI4sdXRvhYkATTLNcYPkbO
B6Kz2DokRGIOFGmgFWe1GXr/5xcYEoqSbNFkpxzJDwFzAdERTCujHpFN7mOj
J4YNFgJHNlLxo/7dG+wajHdhfTrGU2RXufoO4a+Al9BGj1Sq/q1j/urPMMpY
At9qGBl6O26xUI9axh0MiVUr4zgndq5MHw39UTQS7rhvCUKH00uDGiT+CWBT
uC2rCtSjGDGsZ6CFgahj5lamj25r6FeYbA420kTfuLYiwNScihH0xIO6ms8z
9WkcH2PV+AvVqquRorg0L3R6dNw1MdTjQn6UgYOD3I9KAMMWoPP5iq1QsHig
BMzRE9vr87CR4JW2/bgPLUlE4d3rnGd17c2S4HF8VEZLrjOLqMvf5nTMlp+Y
iIFZl/eqfM6j62y5wbywngOmh+ECrHbZnms7vMvNILjC415DSUf2pO11n/BO
LByRsXcA4EkPZmRMEgYA4/94b9N7rgIoJSPaarI6SAtfmwu/0cyLefAwKXqg
vmrBsFcP/rgMSmHnNn1H1EBe5Jixls5ikghmWQ1KwSeqcAzhMSbTMR90XSuH
Kk1EU2jPn1SF/DKmogxBTjPHj6u+o//V4xk1uPRWz0NkN55vZSH4L8zeDRx9
hY2Fu9gcAhyFzyGWbvz4IpGkyAS1xreRsDUsGxS0ZozfCrN4Buu7LnY6e3Qc
o3see7XDsqa8jVwvkl7wxpFW8s0/YDNztucOqAFuTvAaOS5tNIyCXkqV7WSp
JvSwdl2SApkE2S3lw41/whaNeALSp8i/NTFL7Fto1kt/pPMn29V1lsMLB29c
1BxyGUqCuWQuVO9q8m2b8E8ITUeGdcw7ZoP1DzMYGvHmIAfXO2lQ+uXE85/O
Rhh1CNlI9AWPOQvf427gWmJCf27nq79H+c7MXqlWUqhf6qryCbuOjHnrs99j
vXwfFRIhhZ6wli3DlXkkE3vxTZXvXYjB+5oFoYB4epz+7jz8P6Bvo6i17VTx
7n3DsbUVLKEq8l0YzHAjfvYQBeKzsFbd+N9EwHPB+UvWaCtUYev70t8UUnk9
mbLktbg4rnkg8dEZ0DZ62WDas0qv/gz87cFFCDySH6qxfyRpwIX7rtEsrApT
kBg5nOveSo00eHaHReYO+zrJPjsSeu5K/17xQRJsI/ncgS53kY/dtxLgeCYh
uftaxR9bi6hVl5YFEbZL2PQSL5ocXvqQWw+6o61Xw/8tVDH9jqRqfVuDrVzC
GqJogUnlK1Kl1u3r5c0amb6LiAj2VpFbyDKIAPqbMQkyLJO9DVnz4jb7meBp
1lID8xmUZQRwHrfP6TY4vj/k1MREtT5XiuvjWxIgE6XCf9U+IzeifSVJIYcE
DTkFlzthPP76Y+kX2Tt21PHJfAZZ9aEqsnt3HqieJLlBYpVOnX8Ck3YGf0ES
tzWEAtLichoHl4rygAPm5f18C62vg9p53IlAdl73ySVwETcqeYaLFMQCwWa9
z6Bay6kVOcvQR5yOItZ3lsmR62CtoLBg9vyCU+wtarnKsDfwaEfr2Qwsd6bF
N6t4xlCeWUpFfS83ZKvG8R8gsgY5JUVO1u8fqPlSN+ICMoN2zloD1nGKXL1Y
6d6KyquYEz1hEckk3W55rT8pcJdZwqHy1zLlrS8rUow7prSs6aJMPgsp44CX
GyeQY+w8IcPH7K+VFT9uwN7bvjLRfK2enVkPxS0+QNyS0sEJBe+xBWTV7BXr
KYrK+ohdhirEhOJ3wNUq3KsDlCrnkONoS3H8Zid1kPSCHvOyf9t5ZAMQ7Tpz
rrxZbakwPjM8wYeXa+itrMh4xO8KZ+W60ywY8Qf6+d6dn8/Y+70t6Fk0tepL
w24KUuyFAOKXf5dZdVdfgaVHgp516AbT04nj1wnxYYW4KX0EhhyR7sbeSBo+
9Ek9V7v+8OdMTivQc72EiMr2g5aAM+0m6DGv8e0HZxP+upE3nGhjzIv43JC2
X89ufeAAbOcvR9QO0AFMR7zD2V1cTgU8MpnxH6R4EsThcS9Mlri4aAkG+EaO
6adGbkS+zNitPNkfnQnapO37Tni5nxwvBeWnZja84ALax9UMTogcWJSHYevL
79dhFhPAI+bLWVpUeOglx4o3QklxgkG5uKUfRrS/44txQUDekFg7VBMjj9NW
dX7o1uws86ov73WHKf2IcfKkfBoLjays50D92VDa/KqlxFfy4Ha0l57awSOT
lTUcKJvf9Ndpa6Uvy8u6EHRWPtmNaj4AvLEnRHeDhbEkYvWNCK/7oBcrIWEb
NxwSjhvsfWMO7IFCeaMCSCPUFPf7Nm3pTvAVZpKA1qmqAK6xV4uYfs9NrhRe
2xBAa/harN5cnMnrKygGGk70PjVAdLB4h98KKfxVRjGcf2Grytk4vIUtvq05
bRVkYGHFcWVSwTjmuM4tJoC5r5tMVMiPlOhrXBrJ07Sp7WaOMHlWgJzzyoMh
sDTrs4Czs9ENEKy5bnEHOThTsilHmoMZ9O+u9JDG7vl51J+0onEDWZgGDiWZ
WOaKjMiioljvKarGzFmq4+NfXT+mP53twE8Fr1JO+IrVrcuz9VC6olxz7QZA
+XNB+ibmYIP2MTZHflhfjZ3Gd1H+SuGUe3osnSZgt1UduSFhgIr/jgacT/2R
VrZzBL6ecmd0vIfS3Gn+G0qmCqfIiWb4Vlgk7xZBGqHeH57lHI1NDq2877Qx
Kc1rGW94Vt0pPiZQraBhNtxWE8kmTbI3epteyKsiFYjzLm3jh29zHAmhOpVb
Vs7qEZI2v9FOihtdB530IBWh7kEvD6iaj578qPqIUD/AtJun7k39+y8jxSiq
lzoWSIvrMVheJOSsnrtwMtpVs0nNZutcyz7RQJZq6433NZ87D6zdMIMMtovw
KT8jezpNF4F0oefUDwbhQGLVemNcJnMd2ygIBlpTzvtpg2HTw+VNDVsWJk4Q
NSf9/AlVObrraHcgdGEnhJ1Kj73ouY/iYz/cCMu1XmNsQ1n8w/HG/cxpssBV
43iJD+6m7JrYTRhfAfIX2Smwb6B8mrAFvO5SCffgUkj7WU0H9N3kp0iLG0Xz
EontnwHdiQ/ZznCsv0Nr2wXlikGm4ChXbNIV7F2dHCNWmdO0tAZjIIkDwsU3
2iwlbqWDbr4ioOpHKqwXFP8YHLKY8DTCA1yxmiT3nRmhsk9X0wqbnNNqI+o6
49VCoB40a3oJJEOWtJqIk5iw1ymeyL1dseRq0fKlHhxDdT1jhJ3ZpnrEfon+
ABlSIJtVNm3B+u8mp80KnXFpA4jHUrerqpZkBzRnl3a8m1KJqG/2LyTfe19Q
1WuPGJmxLXQ7cyYTeqTW6P2OpvZLNxErGPbm4Ho8QBIB7crtLNegk+xr1tUO
FJWQbSu/ON8C6pmVVoWRRmbsQIbK38JhlXdnmmV7mwXfALac2l8oBuke8efr
F09/BInmT5Zd02LwupSAVpuk08KaG+yBDyizAc8B1IQcaWEsJ5P30TZnwuMf
FQ6IaZSA2LcLWIJ9i+oJW2abNcKI+JHV6ZLo3n0iRlh1m/wfPukC1hNU0kjV
42TNdNjaadnH446c75qA51JfMMyNLUaco5Xr5BynpFZWHlXPynU0UR4KF7k6
NgGhTWbBdqG+XAcSWlyeJU9uRNkPAJtWE0wHhuAClNIKA/HWRYoHrFxgJaLO
nY4fikfwlnc6ETd4JVBqf6Dtk6P65DgzCIXm3DMCnNXnJ0u+Vb4n1K3VNKaR
7Nno9bWcaan3rNP0hMFoEj9+dv4MmLfB8y7jQjAOlqLDaW6NWLYGvmRDmn7T
trUV6+lJbwYAn9AhomnWy1qupqOZl+sL32SWj26k0iHlPQNFNzH1BZimtZVP
h1vI/819UBl+kC6utcEWVxc7lhx+YQU9dPxqAulXLoC9jD3bUJBAWObc1x3D
phJdmaxUai9VBo6/TpXmCzvqcgedTDC6q0cPbNj1mot3UiimykgpvdVUeGsp
X57qjJm/8mDSgHpLicN5OGBS/4rXRlXNt9CIaFkZR8g/K+iVtWbiBSsyfCMg
WygOBeepYXWMJ+30y5vPDnKdAGvYOyd/JEFChxqz4qJY29Ir50aX6lav07rz
kwx/aES/mJmgJ4GOPQQXzaDy9INHa0PgcjGI5mo4SwulE3e90EohKFqdg+mZ
CynhF0jpPG5BHZfBfTVDnUPX3DsrQSHQhCErM+rE25lAb3YERsPjo84Atojk
wOY0r64RanpKF37tk2YR2MTjuJyVf52rMUaWxn6WIxht1lujo5Jr2p7IiUsr
mwNL/TKpHP4FAmZ7mIx5QrRZLZ3/ZbsyIeI1pWlP/TdTevPxkKVPnrRkiZsc
fWATjUgubLG6dFQKOzZuGq5OvKRczjUa9JJQt6A8BKyfqS6w7KF6pevI7jE5
XV2DAF+ARw+QrhAIfk9ADBpMyooH4E8HfbFVwTHZqW8Smwbjn2Mj/9gu08xp
vbEpPIb+X6jTv8OPBsYdTuBDgImAccC28LpopB68UCQQNU8o03k5qgzTckyV
UEfvE96WmefvpKKcOCLzFTYFJEyA53hiG//NYxi0ssQZARxEyw+8I8++dfYO
NXVrGXrLFpwSsM75hEpYbCNBjHyb+blPga+DCoPGuuaxqMw3PMCLEYiNeIgz
mSpE3kJILtBeR0IvW8S6dBPuRBvpcKAAeF5W2Yyi5nZJKKi3E4td37TxAAcp
31x/Zs4FNF2bhYksibOCeluzU4Byh1eVMJfO24pB737fFdI+3OfMdHH+UGs1
yLMFeDwqbLzoembczXtNsdiy2fUnIeh3C2DAWa7ixE5ErXSNhrpzIreJ4bEL
SBZrJESyw3c1TRg08IK7/zqBARd/LWI92sY/jOcD1aQ7A18ujAlTLSKPG7LO
uQxI3HZOS1z6jCqJcMmE2RrvG1AJFMDN7NCcW/VMowSEJrZ711UidmBkTxZP
oL31EpsRLRthuMDnBaCrK0/u4NHLHCFUZdRi3gNYT1ZKVJ01qnkRh1nAnLZC
X+WfwMoDIQMy7MUyrc20WbLZBhS3pjPSaIAkVCE6+8GYFnThiaL/wnn0OkmH
in8i5SsA+tlqIIdXR5sqLD68HgoaFY64SlQYDgDI2fSkwt4VcaYs+Iayesq8
u68jLRE+uqUJwytaDIES/goDmBgPRFV8jqXZy7w1sQw5OfE6NYytJSfQH+67
5xR/xbVoc3uI9ZUxa5molnbLqZ42vZfyzP2lHt0FWsqRnPYstMa3wpfPO0MY
CaGXu522wrJMT1K30B19nvEfioBQ5Wh2rNvPYdiVE9IflTs1CeUKbw/tokOB
e8WcMIKtLAvEykXcbLpkE7tZn+wbq0fh7wNWgNiS8wlmsTA25sXGllISvGR/
t0Ep05F4ApAa7s4+GqLZCJ7NotQTqrRLBUjZd0HC0L+hJSDtqADcUlEe7z21
xp79EG9mxo4xuKL/GLDwyY1XAqyoaAsSZpVlOc0+EkrjBz5IjK5oMBnaDBU3
9PGhjUtqDTuzcEUknHWj9gIRacruD4+Ih43YCIYBGvhq49aJWiZ8rmoxElfl
P1ymiRRwhcG54jVPSOX/uU232FlW3/HcdeOhu5UbPudxyHnDLESzYO2TSO6F
Ki6JYmvHz0stqByVOSWIZ8RaoBWH/+G8rRzAc/aG1MpkNY14asGttX8ENV9S
Fv0K05Jb/bLuhLS8ivSZMhwqVyimQP6bGtqIvwVvpdGVFsqR1wjtdO0+5LuN
EohRRzgtdKyCgTNlhTH4lg5eywHuHGWeMVtxpKK19AQ74Vm+oO/MpOKLhtMn
oQwE/uX267L4hptR6lakHqlb7embYihoCU5iMW0Y/TsVqLXCxZluxo1yKpys
eQDLnHCimHG0HaIKhv3Ptbjyi2jC2MB43XuY+kNxydYGm9WpbnL80hakovhr
6PBufxWjordOsRQvLawkBz2H9BqZpmy+wJbbkUqq4ekAu2OrG7YKFwckdzoT
EB49KAxk36CReChmFuX+iAl9FELjGTMz1w7fgXyaAcjVhkAeLH+uhC8HYgwB
vSJ8giVMaC2N/xo7p6OslYBzpM2QgXn74OF07rNDuAtEkuLCGgowvB2wCO9h
spTtOXC0veV4jd0j8j4ZRhMH1fkKL//w7aTbEB7VbEFpmD5Kjs5rPcQXc1zU
NU6fAR1EC7tHgn2F/SDjspGFTg5QLiLPhaY7Ohkrdrg+llNi37BNFwXBpjeK
ir8p4Gofozb6iv3W6/bjVWoWBP/lAlME3yv/onafJEMutdYn3II3lXy5lvt+
BUdF2Ty+YA5Y2sY61TOvIc4rsd2E8YCL7yNDRQh+ks2kndphk/wMJw2ky63u
noeSkTN0zDnOLhnfucik4bKBqgdtKJAxx1NJeYnIWbRHJbw6tKmOOsPuldGS
0sH9Z0D60Ped+UBHsRB/S0/R4r6GfbRlrTQttryc6Gq0Zfo+ShXC/wzffanE
+y06lLA76s6mnXQkWOvy+31jGPU7hRbua9P5Bm2Qfc9GcgIonQHBXl7CnW59
Hg3KJoIQZa28Ypg90ghyjVzgcNaSGnu7WirCMx8x4Pd3/6/991drnV/+QvDG
WfkLsmpglu2qzuhviA0vHkcExiocbLmiouLhqkq1sTWH7rdFmUMkRA1ijtGR
39PSJRdClCqXZbJwUQbpxtXyxwVlL1r1YO/8shYihGugXSCAQbDe0WBKiwEt
ayCE7YlQ1QvoGl+MroUY2a0f8z5ERyBQ+UKZ4JpSfd0/RPGyAzw8uUQzqch1
cp86aaA2IgaIrD6ZHZlwpXZC537VZ59XftF0vtOUwv7jTvAA9A7qtz0WiRcF
/pEHeIqDwii/uZLkG/GWO/omL+eQ0m6DmlB6h6Sl0pswMn23FOrqBfHrSl5T
L4JjGDm/l01fiX3yfrj6d0z9AtSLmaPTS7r4eR3CT3ibLKk+oHGzM8tUojXI
ezU+d9Diw/X1VFNfYnE/3v2KxmCLR+lUDxHDhhgtLpBbG6mnChfvR/SxCuNM
8XSO6HiPDow0kROl6OIkh7namdxgrUeOqnC+8cx09ETl0y8WV33WqVnfHwMB
9vfbVFraBjLn5viOTPeo7zl7n2sofTwDEaF1siOSCe4zSAOGzszO/LiizA+6
Ff8FnVxVbvlCbh7D9vVpg/+HFvjMyTWW7h2Ryeo3aiuzBQVnv/ZJRd+rBgvH
vmZY3BIwVcotC3IQXvyXPuM/YKCJxZRDhFE2RHPj7LWHQnY7cKEgL3GDdTNz
9Y0Z1c+9DzSUw8tQuS460iZxk2Yaz8AQo4EaQF597DfB+0krdbD9+It8o511
6vwWHxrx/Jpy5klAHkWAX0Gf8yOZantFC51qAsmxc0cTG8iOuH6mbLL1yw8T
KWE9+cx1JOy6bg4StT5N0Kh6gM+xpf0O/T7KU4VteQgD6VOBfVfbHB152lrM
bwzBngOsriBFfyju+KwLc0axjHR/gpIU7y7/qX8tSqj6s7ch5aY9PDLis0c3
JMH8IpxuMmANUlUe2dAgLpJJOxbpKq/RFw/ahIaFLKvvisYdhqW488gC0FO6
zDRY/DTAKs4y3CdFKRtBIyBG3pNrDrR+1b8CjSjVtiuEgZhiiajLGA+anO7+
8IhW/jjXXyqzHBQxrhLfQKO582UbT4snnQmCUe5ZyfteHGQ4DNmOAPqK3xGJ
aNjrB9/CSClKCsF/GRMFZLgvCG3V91Xi+V6vKXi1lV41jsmirzsW/KotamBm
PelT38/BhhaT51zK+1Th7oOtjIm8Mmeqgs9hLzxztCt07uE3qZkWukf/1Xyi
FcGYXG+QErBXGSGvhVptzWZ6gQK5+I47ruM2jUmf89n+ZgMOEuRm8QsJmznK
FyNA6Wy5WuHnMyMtc04FlG4VcdrwJL8O2y5qfwpmGw5Hdmv/wfbFsNAxJd8z
v1qH4FUXYNCXe6lONxnPvHCsVZzxeYvJL/851dQjkiIZH24Qox/07I7b7pFb
RRDss6sq4Wvn7iTpvyxWjWntxXImwzW8Tpm8yEa6VGnVi+rFmcmASQyvDcz0
tDs2xI8fOY8r/NWt5hYRRJJNWLkTm2tscWyVuUeH4wgJHIlOmEwQ8YTUeRr4
6/tejb9laLs4UAD2MvjmUK7O/3ATRaOHbuM9iNbk/5JFiEg5fFSXp7xx2+Cl
f7prn2P0PaG0MohANKwMvKjOQ+UBKFtIcuNraxMXR49K6wm71RpOqloPElwq
ntUNrBXhDAI5lOgovsQvSe4a7tQwcU8LFUuBHQOqDUck6gq2ccm071K5Vzel
azpWJclAGGzGz16iRk4Fm4vGUkN3W88P+/vx8lybhokWZKxciVydBnwRnXAD
Hgh4A1VWu2sA5EzrVTdffqEolY4eL8UcXyjJrNAHEVqKZh7prqz6Azqjb+nn
b9hv1ym9+TfQO8clCK0uhxnqx5+iMFNncqj7tdek/aGOPMMlPMy1iQhdb9Zn
SbMXtsTcxdzxlqYNK+QfHCgdAd9vQ812bpJvEJexLEX6T3lWLQYwKt1e5CTM
NGaUwsmpJgk2060v3XMeuVOSG6HAIMK/+rLx9bIxt72u1dIG7N+pS0UACsG1
ea8JOP0uGGq9ZTITbVMHgFstfrBlgiJNPJFNjelXABKcxC4Ed+pGDCEYkCec
zEbrZMwa1NsV7NTSb5LkVO1PYfIYUPXp+QKszturmpjIKjEdbfH6YvzG0Gsu
D+bBCDIQsB/QwjgBS2NUMfC7jl30RKpYGtvcBnO9mocYTKDl1v57h/9jL3Kw
IQELPONOJyl0NFLCRG8QekUR+5wqEy64B0p6q/c87mMxqgrIfd0dgSahnbmf
UPqOzc8yxZakYgoJr2jf3m4wclG17ur1zCuON9FoiCwIRnIAmHR4R3cLNXTH
Je6BTx7gg53e2GMhkAJeYLT5V7OYj8euXNFBYe6A2DmBjVbM7U4DVnfqEOjP
mQaPDx2c/Uf8ygRzoSV2xJuFj6Hb93ufp25AWCk3ORkqlD0lSVWFXEz1BjpF
2DpvVnTui1eYDx2lELVA04brn+BxcPMZvFUQ7/gz9KpCImawxKP+Kil9D02Y
Q2aEK90gTaRlUCduJjPibcoxFch1beRXbICiZ78Sgrgngi0xbhzjWFu/Dlnn
bGzra3FFe2kNA/QjditsdfJorTZG6faFxdKrftJltX/peYuiRgncpbql0Spf
HbwkxWATSK+yzvy3DKVg+1mWvM1f3NqiMpWxgoT/1UAxWsI8CVmqkAeYjLUr
Ug4fsr+8DQq4p31x8+QcM5pRM/zVwbd9dTUaN1RBUAF9CkWl8vFuCuPt9n91
tIcxgK6CAVq8qWzCIVT9Y1zlma838r8IrORVddnItyaLnSkD18EDbcG+g0jA
6C3oishouA5ewYjUcLy7G/HVnzknOUK+Nh5rSdXIxJvYL0uwmnR3dH1SHy9F
p9tXD0gL6YLxf7J+6kPhqSUNQYiDRgM14U4jqeMeQXCGMIX0ydwRB7ZMC9Oq
VUkywXJonc9xwxCmJZ+hACTxInayY4nVZSitMCudBGGVjdLfJWJ2tVfhSk7D
Duy+yc7krG5V0lObPYY9hXAMP/wmhDktZLnYlKCJSHxb1A/9PQZg5f5hBaN5
Wg4nPH/prPbjzp/bMGTFqxN/TKRZRHpePqcM9lf6CttQBDZpdOCkZnNwFxFl
eDAa8y0oIeXd4+KSivVtptqdtfX/zRSLMcgk3PajWRfvw3VGXQmp7nmnE0t4
YiPeLClat4kEdEw9VdvFgVBeVmZArWHMHDAiOnz1AwH6RLLd0+1d7OroP1+v
0iYkPp9zcQmy2p6x2hIq36sgTv+Q5cYHNO/fjvMuBcw4N9UXJQcRGz5RUUqF
T75kcFoG9Db3bGVWH8aPS8wu96MgqHTc7sfiy+Qlbq2N0HM+WfO9vZ2N8i00
kT26DbbouzXuUFjDT8kq7SwdZpA7yDxRhr+4esLiQuReEcQzRAOpOXMmp35b
YKTCh+Vt/t6CTAzEy2MT5xCyEcCorkqDakmw1xQBzfDtWpAhQ+qiQxpThdwp
Qlf6J+k34FHwrIlTNNif+1Bh1Q0tpnDI2BeQf6LaiGMFQHGuh5c3p60T/6jn
j+qDCE8hU2EF1hFrjSjVWK9ba+kAm0pwpuvBuQkpXvGrYdnE51cM28NJ1//S
yWj2iDH3lDOk9AxC9RqtBYrgOKBpBnLkX5B6RZpc2k3Qcmj8KOoZERSI7tCS
8ozyu5t7ShlpbytiMjuex3UtQxoq4noN4+QsM+8SxwLyA8MABDsqv66Hqhfm
NWysheuX3HevVe9IyW8XebNyHzoJ8xmOvWyxgDqSSnANv7Onlr22EPYn10S2
JZbWLKgLAjDRrVjf1nNAsjGCk0wp/SrE6TPvNIE+WFepSXcQfq9QMpFhWAre
nMy1buEdgNP20a2jg+Q0pwKJyLCrAqUQ71mjNPCfNQj9YTPFx7fIfjNB0M5N
vIO8+b+hjRGcJQ0uHsrLtZZdUt17NFr4tena0cUxJj5hu9eZEBp9clafqR1/
skH1OHfcFV4jHd/mVMwCJlVt62AKsR41diXkXPoGV7VIsJhEIL+CgEq7pHmg
J+vQMKSCS6zlKHVf42g4bXRauuYJrb9koySldPS2A/UkAfQD9NlNGCUloT/7
3AtfddanVczrzhZTvdbgMsbRKtPQFSU5km1AEwasin1z5hB+gugqd9QQDjGE
EvcqDyaN4/qP5kI7I9vcOBjqQN3hJHlEQT5EjIXmDcD9NIfavMjjneZWqOgd
w/sJEPa9fxPLviTItMtwvjP1GPFa3wCOhj91St1h8spU1bPW3o1ANRXLwoAE
A2dYi8NQtBxDXt0lu9hSr7kZqsRZN4n7p1nVxyvDx4iIjlFUb8jb6i3L79YI
FvWMC5i/2r0AHRG2Bwzhk9Rdyj322y80GFL3ZtNGyf4k69T+ebDZTPcLTNtG
aeg0z2A3hajzqdrWvhyjNYl/cqJYURAAc+QQGV76YDRdWx0Jj/6AR/PWsfm0
GgFaaEAZdD1hWmPYZc35hJQ2FWSBku8o3WfIrjqbro4n8XkLJsQL24Y6anJO
jNPqgyRvbIisRv8RK32EjgCfPV4NkBDJAlc4D1fe0iIhCD909NuEQgYgtvXy
1TvCV5TidDdjngkOK9R8rS4nAkdoZUCyUdemU9AIc37I9BySCxXh1L4OtEmC
Tkh6GwiY4hfBkHDkIhmF0XuZvPgkxiVItgjZQvtRMA0qYHDxcBMV9hJPK05/
wxUPG9rgwMg2W3T2m8zpHP5EtzAnIA7YV2wSGLFSJ+urWZdJpFfNX9hRIot5
KhPTvwL4ELryiJiLhoSqozxfhLa6N8rzvbA04fusBJyX+N7dHmXdhpsAo7p/
tXnhVVj19fcUd5XhK3GgS0Oj2hSrXoT92zle2eP+B4cTqGBkJu+ceeYaQd51
KHNBwR7FSpbBUWAHT8D7UBxI5VFiGdQqdHZ5OMUiBSQ3fwwLv0157cCyrv8e
r9BeEFeBMM9WaoaEeX5O0fYUrlCHEoZgvwK/BI3VhUmUb0r45caH+KBee1yE
LVrgqgXttDbmPvKKGnwTQ4apRZcx9eVLqMECScMnuA6S8GkYdNs8vHN3/Apj
gtfaHfQ9IbwPSADkTqT4RF66mCi6d1WD5nlIPOqMomx50ZZprTLK4+G0ZIYP
y6GYRP4PqRkJGtHqV5Qvfl+GyntQJD5/awq+WJnlThLq5Kvb4II4Gk1TLquw
bJiFBOwzvq/0F70BGM1+2PH3fgLXpfVZAuZJLtEkxRkLnCc+SokaYV5h5mfK
wq9Yt38IjvBLsOLTATZDxniaZKZlJFN2fP8I60iY4u7m17Ct/UyLQ6VtL6uA
uOofjZtu26NHnqziuVmlpiHUkvC5vjsVLnIORsQ3YXfopwIii5O0kwsXCVC1
/J+8hFQA31XyLKkNqH1bOYchDq4+n4IXRqhySmbMXdRolK7HIND2lj7fU7Uu
DulCn9ihMvtGkr/txkuVrlUp6EfdJ83p+xCNVNMKbD+RXC2+iNQDxMwR0i2/
GY5wrr9hzZY0ewpmFMk/HsAktzbG1oGWGHxxlRVhjtIRGL15lPVL+hPGS4V0
UwdCasWsQQjYdU0GZYR8E7nJvy/G8zv/gCwCeXoPfmrf+wlz1xJfeDa7Vbjm
nmcX6zizCCiqgFQBM7ZrAXAmLob27khRHhh9t51YmfELnp3LBfaJWHF0jKsI
X4rv353u3GRKoqRRraPZf0+698yd+ihknlfO3yjRXy8uonwgYJSc2eFsxZVr
gikqCxFNPL4Mv9112nUMFuBWJcM5WccYrK6qPKGE05txyIJa55aRKxilzBxy
N4HQcepIku7Zv6928exP4AsEDU1BLJHV4CD9OET6NniH6HrJoGKE5sYAbecP
l+2BjkIATT6BNoupaQbK0g4xzleEm6l0qLSjnAtt57nkpcmDWyjY2qMnBgIf
74vTp90z+1GDVTC1yjrtqg21o3ys6kwj3CItgqwAIZW4f94UjMWbzCin8ggv
sdXh1aS59VoiF+7piumYM5uR1DfR9wuu1Fp+VxJv5q5Z9O4UEaDxO0wTg8cd
/nDndE5OpXnF0dYxikAM+h1fQUaKvpf8TVC4CC3LfRbA0aeQsqGbefQ1MNKs
m21wbBBQhpBWZFHxGtCTo5t58zGvbKSnM/1I3AFN4dcm5Xg4Pr6m5G5iuAqJ
VziI3AvWkXAD9FQF6AwFiXDFvIPTMotWKTGBb9mmoKv520z8PixSltlq3ijE
aJmWES51/F+rwkSFvKl81oFXkQe4P/z1SyfFPf82Srzvpc84YpbNb0C2tjYU
1N3mXGzVNh6vgxsCxNfdn1mEaoKNCGLk6/OZ8PYdBEzWNLfOTZ6jloULb7JV
9qcTYZwYxfgo90kiLNpM68GH4z85adwyg4uzCepuCQQZ7yy7+Y4AWL/QiEi8
nX70lzAWfnq9j9sudeWeUrdCT/u3/wssjN543GBznxpsl1S2668NTvtU0XgP
0OpC1qR3Ybo0ins3OAFhf+18FMI6kewEy4RmmKI6Kmys+yjFx45f9CfYoZs7
+b1SmLZiCO+Uw+Tfk8r2yMKUoeUxScxWSch8f4ZHNOOaPSwa/sFvsT3vH6eC
LsZqGodgYftgKBA/7aUL3hju3WnhZNphe+/Y1hDFwbkOMgsbhCINFVbsnRPn
5IwQEnhkUSXw8Yo7E7j1NwAa0Ckd2/ufyAndxi8BM+21AZWNYItG3i4AWs5E
MU0KcLNk7BbOVFPsM/egVo0phYPglaIo3McWnOi4ZWCypLWNxkAi2+rhzWvW
lcLiVBENSCyjyvN4Jm/j9cjZptEs784DzBGKRVG4i0q5MZSr005HrPKoZrfj
nSIGnmvgxYdK5EFYiAuIllgswlpBPd+8uYUPjslEPZAXjCaRsEoNCL8XlHjh
xy1HXRfqqGz71b88u4DIZBBtnUUgNRq4r7qvBjaL6dpxclEyUQFIrV1rTMCY
t0S1kAe2lqQdXWHnZKZ23uuhtyxGNYcI/X/YV9M4v5VKoN9W6dPiZwPrNzHx
vLwth05L4yQ8JKbRvgE7lqS47Pw/oxvjzTHus5THxJ+3d3cwY4lqgIuNPuQL
mfsU45lzuix8oAlhql6wp01+SlonIks3abUnM4b8Hx2tCzugIe/RMEZEmvJ6
5+KKki28nZll8tlHYJrAFVDCByP3rSc623deBARlX2M0R2LhAQcJW2PmBf3l
tMBzFiqEYsWnI2Alnb7+gWm7K+CcvCZc5k7cXw6c4AB/jG9JE++ybuhLMzET
YQAyii7JB/89KwEJyj/NogLbiMuIydByuuJU7FG3Dobp64kLEEDCOIKE4dMa
GpZXHxIUf3aThxnvjrFynl6WC0pm9vBn7b6T0c2aozcRPSR1FjmHUdlO6KkB
ywCcBiD5nJeo7nvf7JnU6eTA7HWGirvu9U6zJ7URRplwsvg+opOKWM9DbISk
kitllzde4vd0WHooDFbTcT0jm7LbFJjQDd8HfS2jloqYjhz8CUjdb4d0mdzk
n4iXCsc8JrSWJ+k46AZYs2xlseFgxEM0R6iLCUY5T4i+QvyAtP6HqwrG/NaV
Il3KnmJ04D8zVMlHPGw99vWSkqA+bhCwr//Kbup6UOusR5/j7AMEcSTzaO+b
x6bWqjAXCeqo4GQFFxxP7MOHHCx0lk4Y4UTpv1ztJGcarPyzyWHzUdn8aIT4
EZbpOg4oOm+VB7Iv34VFoO+VhRKoXzU6/3LpvBsIp8fVkzowm9j8Iw01lKgc
bHLTrJs3da7cFf2UifgRk6dkMpElpRC+OQIfBu4k4CGKBbf9163DkQDYgF+i
sHJDQPSRCEnmPOYi95CpRKqt4b+udscggaIEquP7IBfFK6rMB95JPNva42kP
Ssh/l/B+Xd4KVIvE0JVhkGwlDdmMkzKIltKHkQ3zHNICD0jyZ+aKz3YXE8xA
8TYogO14YpdqWd9vXk1G74cPAXAziJoD21HYwXdzH0rnkQyA/r5DUvsh3NIF
A3C7gU0lHN2CnP2CmKtTKNP3kGk8LOBu3x6VB2sp3g9P/qYm1YfPjzLpDV/M
cXPn30PvjaAUyuJ18xbtFXn5p/ZREG/q62Ibw6ArSBrsUdUyCr6ShvN0LOhu
A4C/5fjLZl1ZkOkiTd1m2xz0iSYzPEB31Dsfdx9yYHLrdnjPu3Juogw+tidd
5MFhXspVVbgPrjBKbsc5DfX4Oz7elWxGc5Tz1VVIp11VGseRgG8YYsk5xW7Y
IHSR5OoHW6f0AXerhStqWk4SfGnbHLFkFl3QTfJkK1N/wPDrBdPSZPs4qc/m
a2uC64NeLYPI4fnOBWeSfYTU74H96ajp/8o8M6lMxeEoqgrshlnXwpKyWuMM
5rKfkKw4u6TXTWukgX7LOp4dmuBAt3FrL4YeObTZuFyzQW72OobNz65zhyna
eS62eyZJA+xdK+A+RNrZ+ZBKh3Dj4/WHmi8Q8Ij0Ve6A11vcSHOxbvnyv21j
NW3kSV3IWUchPMuQTug58PpIYG+b86y70RrieHfX5KlT2wX3kbcqqpwxVSuL
jw37zx1T1pTAuGgKstF2+PT2HynHGr5j/2Y+7alyDiZJCDr+3GOa8+s3uqpc
4mXbhvb50AUMfG3ribc3oF6iSZb6/KxhAyCg+v7CQCLh32rKxdi5/02MyiLZ
V3S3SSyioAUnUT5+bO16RCnfE13fZguoY+OfhfAduwiYa7dbbzrZhwuCbEmY
x9lKzye6q6gIHKHekkqlzttCsAk025e5PN5n4hPhlawlqO8zJbLwsocesW3+
OB3Y6Q1rOX5wO/jMYeLKWCV6kY+i+FtjyVkD61vPyGadfBQFhLXztKPMu7JK
AKuLN3jXoNtVqet2n+12TNAPWGTNli70h0KFJa6CcGPNxGgGuJoYZVc2HOnr
ZJHRRwG31mX5aFQkv5f57CdGCa87ic0+pgxaVuk4ZvNIpAVfirE9MwY1UBpp
tAVJOp1olbFRHFTOlLmplF50YgG+rGaallsbPaEO/F+eUo46XVQar+Pvn8bQ
rGmS5aLO0Ad00oMFHg22aG8/cTKhJ9tkrq4sLGb1vEnU/wFG9EmDBksqXbZ/
VyoyZXPMFn0ZCq1q09m9SnIFdkG+/1u3+NSe/FoemOze0Xo2GsnecuX/WA7x
J6OO8EHri0joN7jqS757A1C597j0J0KUkH+0eLl6+xWvUzILtvuWSjCp0jOz
aIICUi4iTV6aZT1nvnp2DB69pqH6HD6vixf826MaDSQbEbi5ntU1Ni0gbpkt
IKYPq6S2R86dZvt0oh97ZafSlP3UiKsZdN+guZTYoaO1rfUVaYOoSyZYQHWs
ahnIxdODuBJFPk9m1ooU7BDK4TaU0M0mElFQomDqRNuqajGYZF2mDWDk5Jab
EFDM6Jzgv7JI3Ak7It2SxbTtcw4cuF1MNgPL5mwNVyslu6xcI+9V+59JC9VU
dcbgbiYatq/dk+H1gM6xWUEgxrzn99gEolEP0glCsyihsnho7E43LFgKs6kF
A0/Z65doDEGGdq/eJAcKfurwgswAu0Oq+qrVxNrNucACrdoCEVcRX1VDuSSp
uhQ6Ybl1P91gzxGzsh7TbKo2mspP4PrsMflMJF2JiG79pNyZjPugItcnm3IN
UxH1rcDExp15vKcB1IXIIRnbZvKPA3TA+Av9GTk7Hh73QfZxCiiaJTAaCS+Q
8jXaPUqdbjUMqL/e7wwYwDmTJoaNzijI3HeW2XJQB+lGDDa2p4h3DS+dAsRh
AFNcDaPaJaFWBqHZ2pXZ9RVpaIYmIskackMAW0ojESUqUa+Ud/ScULl3eh7M
EgCMbErQ5xd5LWIz408OuNQdAwQ8fxzJNB2zIU6T1QVX0hj2KK4uYyXq/FQw
Fmb8Y3MkH77AV52pLfzPK7p+6MUlVjFt3mQjv1T6fuqfj9oXzsDq7RCUqpMj
8NSU90bbHE3K2t1kXwT/ZsZyiCdAvKVjuZCKeS4pF3ZHh/aC7TmqOWJNXxf1
qjPktkQUlD3xcp2NT5o7I9EhglLprczcdW05i/AIxJBRozfQ6MtecBFYDRaW
RdfoCibc93fvlTQcg8jOmBBIzI4Tf5uMoInDQIuBsEetOdjxnDTHBSSdN/H0
ztp1ao8rzy/ZXHk2OfYCLbF9YA3SrUgrsqJq+rydEE8p+wa/ZznOGMpLDqnb
CNClsLguTO1v9hZ7GYwB2FFbZA55zDzob1Wyvv7iWAbsPhkxCJsk6FbbJZxN
+LwBNRgg83f9jXlPEZLD7k17V4O+HjVaVByX78NA3LH+csGLpcJxdH2HvmNT
a6r4NBb87Masma06L3P45BuNLCyQMQGB0nepo1wYFBa5qk1X7y6pa7BrtXU7
3iuRtwAYJDSWN2YCiVMTqsu3rjzJkSQMA8Q+GLGbIfGZ7lY54zaFPw5Clo/B
fpDtwP6oZ7k3UNJsUXOTy9tjjbfJpEL04avOu0pKZ0yrwT0mvztyVAoBEnRk
iD1nJ82wu+Ydu1ToD7UZAG1aya1ykXa0IQR0obbfhlhh43kLTS2rGCuf+vG+
nFW07R7nEuIhBO8o4tHvxZdfrGU/2bHCI1MqcTKStTyn2eX2Y1VTZtAFF4b6
O2wdld/5isUHulwmMgJqkTEGAMQIROvkju/nyA1b6tlItryynC3dmgxZg1WU
htPRtr1aofSCzmVceX9vgPOKn6EpzZgpb2V1oqh29HT8LhlTWOJa/DRVD1KV
3FSn9cBmHvITN4BfbtcQmi0ykZXTM7LTrm8JuEISl0LxTsmOa5ak/VKHnkXd
6inBjPUq7GkCn7dzFXTK8YcQHNODiyYf+RM0zAG3RizVjac5ObH4ozfJfBmc
+8JyUkPucqejpiua2H1sLm176zA7qt783u5VKleicPCQttszAPMDxa018RzP
WsQTB4iqblWQ5P2KmASkXzYjOXoclsQS6svyb1GlYc3vmcGl3ehPbY6Hjs1D
A2XQG6XWbRr1ch594jMaRNiTU7+eXPpQR7PfPypNWNS82QLJQs2Ga6srOWNj
WAz061iI6aiYA9zQnTf2moHmuJt0Fcrnm5+fUPo0wkrYciQMbe4B5feXYyPE
7NAtQlZq8mE+4TnnnW4ui0obeL9ZNGKiMvN7MxCVG00igX7AD9/rOWeHU2kB
9yGlUz3lDIofRTVgWzuvPGd+cDkfr+4yQtP7UPURhKklvTEcXdawiiGI+L0Y
MMa8wioM0vwOaJpdVEyKUV58lEDOZj5ymYqFdBw/9hVnCTbbITcpIR9P31OY
UMVFEzDGOjOtlL2hDNyHpvFO0CzSIbKE3U9v1OHnKeoJq5QbigXoz8IOenn9
JIC4L/2ilt/IvLzLU1A7V4YGggmlGGA8LKlBETCDv+di+GKch2hXv0UNrTVi
+bZInToNK9jOiR/G8PTto+C8x4o1MiJqjAG7fmk2lMYu4er3D37lfONUUsu5
bezgi2h/cg5JFqHBpb11WYUTgW8pIPS5hK6FP4162xqF/NOm/LVVmFa1rS3G
WjZcr/lfVGVMyjaC3QcDTyWfIQwi7o+pkfk8EeMFfwxY2RGCzHk0pimq5Np4
HbJ3Ojn4M65tNmwJnM46ShSVq8bN8V8FVmQvCkw2/gkNIJv9G5fXwSSFsXY4
oK9567N/+jskm3PbAQ2adkgudLSA7cfvcRwVNJJZlABLdRJDd7LWq/XUrfo0
SPhTBedkmfrupXF273ESV0E3OlJbyxfxTGHBHeodNXLcvfQAK1V6FCQkGT+o
vJSOIAs6DnP+gfea5hH7GIx6lzKKUvIQZIs6Hhg7HZ7pFvu9OnK+EzrDnvUW
xId3CeOLyNxPegWYto2Ij2hCAymvpsB8WrBA+Ga0G5mlPhPZzImBmb8svd63
gq8cykVTmScYMwkav3ohqMGiVq0WUpMXxTZv/UPFMiIGOWkj3/LgzRvzj8/h
H0glqzmvV3D1bEuK0WnevLuOk3ekZr+w4lZIBDD8tZS57XbmLI7/K7XB7o6z
3TQwhqpIo5RFQM4ojW8+NE6JgIlzJ3jc7ioAyC6ZDCowpa9a1Wqa19a4LTh7
xwSftx5J38Ro+6TkN1NiX/gM8QWMJ9Hk3VRaypz8ZDPOPiLnV3BrZSpu6Uiz
UBsnEC3qsLpQDA/jvXUH9jd3pE6NYS/oI/tDb3yhcfkDuTlq8c0CZK9T7xCO
M81/nD5BGpbLQ6fd4vqivPB6YPO46I3Ti8iY2WxqtdgPHi8blkdp2XhDruza
YPK0WFjzv/sAX/tf0QZu60yAItpyocgQLEeRS8xZ5gOwnTa8TrbsTCFbQH24
amsPbk+7CvR6KkyFyYcxUP8TodfDxqx+LMnVx7inXezY521bVKKB6PTkzlxr
p92qbjBRLYiDhkOQGNwnx9bCCZ/FlO6aeQOzF2qIl73vWqn7INHrjgcsZOSX
w9jhicRdZAUO3Q/tvOyPIhBT/L3S8HG1TmJsmIR0eIo9WpbA7gd+AHNx0eCp
V2kFvwnEeramoWGKXsD5NE3gmW6N95v4tpytMi74VGZNYnbIPPJfsEysptj2
doACjkyo0aFxtTXXhT/QqUgMM2hGIWS1sTjrnspHpdEaQ93ivLZbOLxaP+xB
fIbaPTgOj3BLpDmmuGoTc0/qbqauAcyQtS4aZhdlLhJnM7nvsVwy7Y8cpwSI
GujqR5oqzg0/ufXhIvwyY2hrjvsmqMsJJ4R0fuH2KFWEIeLkW/a0yd96V8mF
cTN66QJu3CjSUMgatSM3C9NwvOCv1g7WgHnXfSB52LAF0BUnaFwO+YuPMxil
Ez4RF8oKwHiMTIFBu5LkuJrmkOhHs2s6emuRq8EVIrGo3yricR2EdJ32ZZVO
F5mVuokZDwT9Wiu1D61UP6jdfSnfN3/1JWVCW3HrN6be0EyouSeu3zJUhWVI
3CHondJvzLTASV6qZHclz+YsTnkbiNnMAUj9KlKMGUru/0ixHxw1bB2ESXI8
VzD8cg7qNzaWDqQT4nIVqzyM4k1/gTFdkxKQ0WzyqamBtxyqhVKDE44n5PEA
noLmG4ohR0vuVK9no5lMaNRI4mihqxEmX1CPcYvQmWYGYlmUbtRghqjlNCIO
s0w3oHnCs1SHH3by8XygbXfTLlNJdrHM6kR6UuBxf1ilMFGTzO+K7NYTETyE
edhHY2JewDQzmk6m5YXBaAltGVdb7ZZVxf4lAnvA5Mmvn3ZmF0EH8+g26I+x
Y9bgm+iroi7vg0uvAPVkWQEDJfSeTPAQD+lH7G7yfmhH4VyhiEC3pBa4MVeH
InD3PTQlUgIkLyQl4DsxmsFf/v/UN0CH3GJBvozUuq/O7lJsC4jcVY57cIpF
yM/DgmZj6KzCWeO21jixO39wURz2YZllwTu1XikfCm2freljMTz0SvqaWORo
kIP5SNYl1sWrfGv7KI/u0jxOtyIuI5hzkOEV3KstKGT6WgpwsylxFqBg3deN
gOCagcAafkg5nBc7AadQeDNi7SmhKpUypDDJGvu5HqzYOwJBiU91Bfn1FEtp
I+DENeXv1WKVqLJhIJYVZRopm4rk925EBpYbaJ06Ua8AtAITSG8a2fGSv8yk
sVl78rh83743xWBOmW3fDCwFkyv0YxzLB47Sy6l8XFW8pFJJcKcLOnLaU/hB
YUCVHSj/CJIZixyPXlZqiCO59g8+hQIsp4oFMg2cdBTF4u3AHDa1WiM/tyij
0REyGdtpQzram0PFCpAgzWoAm9pbhcZ5I05x4p4aqh4Uideg0TT8mFxrNnZj
YEh2DG3hlQ5UiWUvG4m/LaqTSRNZIUM+hZy4jnewfhogTC96r1OenNkzZomD
Glnqt7alfRPhyGIMJbEh6cIcuMtoVMWzmjM8eyjPuYZTquCdZbE7nMO4xh9s
s0Pl+JZM+4P1o5+MhILk5Puec1wA+JYHEZgjfx8F43LCoRvgFALcrE1rlsQl
7+RzUYv1prW71MnQ75I2L8HXR0kRgNsxiPv9jZdn9bFmTjVQx7lLEVYvpyOT
T1xfUNeKxzdFAPyl87sMPbicoCUMad/+SAd/ECdtiAqKzt/+BSjyNP9weIlR
xm77odUzpFQWjr9x1kxtyDTxjz0aLgojpMkpGdjJp8hCpX5Ewrcnxd630rSS
rgL3ejPY0OqdovB4idnPbf/3AXajHEaqy5Ukr6TILvj24fbUXxEOxQG+XcsB
pBvMa2q3M2zGfWLs8mu7wQO1FuqjRwnd9pmOyFGO2pTRZhAi1fJFJ9dAndI1
ObJYd6lcP9rxKu2/L7k8nkARDvkk3who8WDtzCDzVanUnyYng248d99VMfcK
0xvcdOhOLM6c0/v3ZxzsUuFax1qlUQKJ4/QlQDUj2tfdg3lMkDDtQhAfxt11
3wvYfvLu6oM6ITCiTz1cmxfFFUi8amvIEiUuJkGp63huXhuMaUtYcMjpLIAx
GJN5GU+KAOsrkfPO5cYt2yKUu+1j+GI97OdrW39Hi4tWGre/XSxRoA6msjhA
h5tJI/muDaZOtXjX8dQ5V76/163N+G6PyGTyGXQlEva4P7EUt34ZX3zqy4Py
FgVCSpOXQmEBYGQy5BDoK/HFrVbtDQKJkDyFWyM71N553rBO29iGW7F9Id2H
vauVxnRugJrQcK2u5nkzLN5ZNm3C+XmPqwSrxYTtXu/cJ3w21tL7wvJGhl3C
UmHsHX/0Zkf8WNKqxos87X33msWXqv24Psb7vNU2vpW9vgZdJWEkZBkaNQkF
QtSo2W3N7XwYuGQ/eKHXAzzDVKQl5gccIcAtIqTnTsqs6MaFkwo8zV3nMkH3
2IvF/dW2CR7ZzHh556PAH3Ib1pGcP9FY+5+5C6KK2CMHzv8CSdLtuxoaVHS/
mlFAJwPYTrYQi1eTxCjXQnwvBHm8doC6cOxaIOiU7jxVcCAWnbWQZVVMARvl
Zlm7BeTAbbd58d6QUI5x82YzbrzsKAO+mpJQxNI/MQqu5w745V3/WlrZcHYm
CguwKOWImrqTS/U37DzIZFEDCbcDul/vsdroNwa329mk254Evh7ny0nWEjaA
coxmmxt0OBUFXfBoJv9zDN4yccIfeK1Qb/61oFE2cAKjyvkXSOpPwwDGYCwN
hq3EtYlyyHCT+zrj3n0Wh/PnUsAmQCm+sG09dsQp3MmUGMTPPTKpUsAUGqVH
l/h4y2N4cTEN8l4EpDd/ul7HXx4UFaJbhCjwBHpKi+z9YQcQxOnOks/w2Ifq
Q42avC+jUy/zb3O4Brs/k8vnmKmkQvO/d2666ado65lkKaYlCkWtsFT1V4AM
ZavOeK4P4U/YvEagYZPyv8x5CbLMVlaRr2QRY4mcPXhDI5HYXU+mjZek2mtN
a43xP1Tva0/WGa7OL+l1A0Ehf62ziuEYa1uEap9XA9AU9hRt9V2aCzGkd0od
bKznn1wskTvYCoaz6GWzC/PGu7/rW1FvSpNbMF5KRCxf3JqtQmLdvZI/nKO+
2BQRxn9hDZvukNmn7gVl+Mq+Lnmo/8epTF92oERHPUZwJxClSCajM6oioP6W
hknnqk8uHrl25RmtByJtzhrYb1NcNewPPFuuuT/gGUgAU5fT8EHNk85p7+uY
8t5PLVf4fJXMs4wbtqmzEiNPZrmbT5o6BZyfL5P6SV1XCIa7Wv7r6gFYVe3Q
wOpyBskAlo6oODvZqIvNqAVxZOzpT241r/YXythAMm0UKj8TayAyVGpK0IRC
zqCU/Zjmy2Lxzav2FVfSZb9fEPIUw/eycKQn12sSB8mfgM49Y5VphtIbIl3z
PTmAAKA+jmwVlvON0fmbOdgl/rQwAfSfsYLfCJ+pbBFZQTGEw3zwuVYRq6p7
YoptGSBiZ/erEEiVhFVyHSEGiGuS4c6VAPB6hWhyq6ipK+CYLcOcSQhn/Yzo
uK2DZGL57+T+ws8qoHxjujUFaBQ0PMKHbzxShJ8tLl6PMMUZJcaBD8Bf5ACQ
FLRnooYoN0fq2ZHzVcOyUrNeUVTRFyl7oDmf548NU2E3cjJAKqdwTbm1riFT
MkLNMSLX34VY0Lm8GghcvGX4sZXSW7CluibXWz+0rH1NlbIJeNlK/rkGQiCg
bB92h0KjK+eTQ0qfKrQqZa+58sJ1XPY/xeWcI63p3vMA78hN3qr5NlIFsf6R
p+HXAvKsE8udl/Xhe0H48doVlU+77iA6xdNqJkOa6VXYLW2HWoUSqQmBPwdz
9XKIXKKeGGEAfohSDuMumXMTXPbBPZYmJDjUtirA4wGljjaYGafHuhrP91PG
/3vaycfMVsTBWjjzrcFrHen1ChJzKWqs3OsrXwgXXNdmdQ9NRMSg27I8XiTR
RQfWRE/mY187KFT14o0yz+To3uYyEODAoG/uEsGrT5H/vGj7IahWWJ8jNs/B
38N/4/5ok9ZOSFK8lceeKDB3AweMVGHfRIj8WHMDCaz4BsD4A4lWYKRc9q+/
sF4bVn3d8a0UlN6jluV/o+so0WQlUgGnZrI9NyAHhWzuTlFGh6Jq0PKIVdPc
B8+q97DzsOVdPKsn3moXbfuPMiCzXnbZrgWI6P5QCzoLWEWmxdEYBTucxiBH
6A8O3IhFRrqNs0Fjk/L+KdIpOBpLyyjBgq2PrBvhJmv25StXqbRWmjQtso2Q
9VSl+SnypKwog+zGPiPmU1vraY8R3kbppYRkLyMbgldf1OK7TXKv41s/yDsi
nG1WwpfC7EyOvy8r+LphhI/0GUOiKDZ3ewxJTgLVTEwuwXMMbVgiGbxgppgf
qS/oHzN47kE+Ee1buoZzMKl6THTdbbGwX+1in1drIRw9nOyXTmxH0+mOlt46
1bDRfdj74nzLdiezOPoi+uUk1fks8wcIFGrkP5C33wmE7UmDNqSnYxVMxNmg
YLehZLcFxYQMuqgMF2b3QK7Fg6p/+AU9Fc7n//RYz/HNfW0yKoPGOHTXQoJL
YS/tOWU7CF2qRpK4kg8Wh1NItV+IbkY7GUwTkF4xtbBgo1cY/RnXcpeRAU0k
wSDHLS0CQEJ1igj/zO/6MP4oP3prnAY25MOWP2sYH+TFt6CYVcusbqmN29H+
FNVLUTodVe/he2qZ0CtDT1eaBHOi6j7OH/xSt5ojhRv7he6HhJAxlgrOdeai
t+digmkLuf/RBU5dh1H5QIikH1zMmP7Q3Wd3jGzToFNBk5nfhR2bAI7Gww4a
/EWu0KfyS9hLN5dwX5239QkNumAX7a69Dv1xc0zn6UnOKy5dmuAKvd2HlexE
2wIXYlR5FBpAXwOn1fKMgLrREZsRsIt9W1T5hwNsTrZ90naQBpYlwczX/xt/
0Ub7R2U0jykYCYoVJtAXkyPpXxAFodt01Oag/t0Dcp2ltNa2n+0dE/etPHXI
VkOtvL3GcP2hwK4XEeZCu/pyeMEZb6JNWxT3die3MfmTwf1jmAb6vj7rqg6l
ARxmqUdab39aRDCaV+a3eM/nsboBxdX8iKflHLnVjcj9d5HajR1YZFYrdDzm
nxJR1ecR+XbVVBct21zdnsmA+KANyw3V8n5rlrs4hDVgwlZGQ9hiFN+VYyFj
OAHL4HqAzPNJn8EnGllAQHR4e/XGpUgWrZK3IK/zGn2os+MTaXXJx9dEzkB5
R7CdIE++Txtm0UDxo3nepqRJ5/hiZRTq1naIKicFImGyT7L5Ovs+3bAPlSYf
XstjeltZhdWlLlNt/r/6NdQTiB3bqSE86ZII3QDFB4HwNg5+82oIeNB1w5t9
n2DyhWRawwOmlSl5EBoZR2hREsJl0A9ezZezLZDQvpJj4PUe+0T6L3MGNgKt
jimDOqJJrf+v52CeGD08/RlxEvEjnkPU7O6vhBuAbNIr72+ouRiaiMYKwZ4G
9nrviIFhnhELlZYG2XO2pMsSpHw9a4M/0ccnQGCojrwpWpeDgSspFlcZz9iT
2J7bfIa5yogz3oCJGtf0ppa0EwxpE2+EXSILHvIVfgfmr9nmER//Eaz+HXDs
6wGf+vm+fCruBSuFYhITBgFfWyDfnrS8meti3S5zgDoNpbY82yGDtNbH8Tcx
u28v12AUYW8AiscFtpTpT9qfywHK3Ibzxt0L+FeUdR6KNFmfQa/EheSQ1//5
SRtiO8wP7vrwf4iFbLnB4n3XklCJm5G8Kccjwp1RK2qJRp8fK6r5DabM56Iy
kExpD3Ks696kimGTFEPcoyDQM5iIU29iq1AtThxEjzVEbyd5CAkfvy1wGhCR
xqyC3LM6K5XyU+DKg4zLsC4ghlR0ZWwN9KjtaIgEJW4WnC0x73HtTa9viM6u
iuYHUGBrHWjV9VYp2uBq6DcsVfQJjBYltSxng72iej78hzpS4JMhttNZX5WY
EIu0/+YQHEFtPrCdzM4ca7TsYc7l0u8n9zOExJDtMo+EaotMhHIby3iL1tVY
uqjyFCMlSO5qlix0GDbkQfBhA87i/P09jFft0b1cQfWyVvtAIz6ckZ/hQ3/v
/JkByWqFiKJqwpoRrCZNKUb2s1E//xd+yrRH2z1PlJlW7y4ChIqi+vEV5OcC
zeIH/0fhrVqZ3NHv8lOJeBHLQ1d+8mUSUWeh4Wo71P1t2gWfeUw2u02pEAOj
VyG7VZxp3EVbpj/rQw0Bphd2H7OeObFPLR0pvuHXZK447HLpfg3dYGaIdshx
pp7R6LNU/ZYmicsrqJV8m0EdYaWmjpoUwcMLjL3+i6GgTkdQ9dGyQRg3rws8
vhm/K8xONRA6Jw242dqHle/em+ZdVy3JfA50BYAEQ1F1lECs7U2pkO5di9l7
YtW/GDnNozW5tVtVOavOf0EGGa1z0sB1WwC7YifHBxs09lxolDkFip3v6WZr
eaORTd7V5aAQxJ1+FBYhf4BYhebKbRakorDTqb0JPv0GcaOTfwUGp5Cuu8wV
LEJEG8CljJl39vv0iZJYDEvSfdY6iKMXICGc91jrXp8S+ldZi+i+JiPe2czB
QKogJ12X1bFhx//5ov3EdXcPDIb2sBIcLwBZ6Jq9262Lj7BanucUtF4DF2oK
2MMuXAtttwuZL2flMoUvAZlBkYB13yVEBvpWOnHY9MD2A+4WdJEyKoVVk+cn
Edjd+alAQNVNrSXo+bv9a2TT6/imiWul6jaxO9guWqRp9SxbdQB6NFuvfOw4
z9ouYzozH2ALHnCoyscy/kwhNscFs4B3bPZ7WCRlptEc479NeJlh7Vo9yXm/
VIZo7qDXQucP710SEI/u6VzFzXPQo+gwffIuxmqb5IVABv8L1w6xL5y/fZwT
LxXjBmvPkfiG+TnC6a0FEY4tZY6W2f92T8Vur+GPuMPmnFtb/DWVPyFFmVkE
65KqNWjl8WxBwHfD/tO48AwrbxXKF8Xir6DKg47Phdm/cmdTcEkiA3J/BaAk
We5LzfDwxx2hb3QurkHaUCchOYvkNEo8p8C6T2Qi7H+UHKKn96yDtR1GOZnf
2haeNjPdOD4tmyLQwqCcG2xo+Lp+3XW1MdQJ4/0OWf4l7p/Kg/FFjlxePI4q
1lIPKy684l3NQrJjnq4WDPDHFnMXC5VaLN8r+sfLyzKtPd58eJuI+zTpfLH/
f9pHtNhome8qsYIfkF7UaIwDntcbHkwU1Xy6mdMBUdg9zmGHYJnHGyfoKdAh
/202j/37NSAz2S7oV+qe47PwWuV8C4+Y47tgk8ONbWgiJb+hY1GELm/++4r5
04BXG22y70PEzTHupLLxoMBLkH1WnHhwxO22h0ZR/2/2VIuTIssMCsZ206MX
C18CqFVea22G6kAm9VlJcLyqNIjIbSDnlFzO52Y0yNv3CitGh/+gSVaKqBQ1
cPasT38XL/J0UTyktZ4BuMxcVLwve7/EORoLE/QDKgVIfPP3ou+QQhA0w0Mf
vXUPAHtLzE09d8o0EGh8sbwobHEZHSo/uuvOP3ZmdZppXfnfmwMyYN0NScBv
RDm7HvT+xUs8AkNPCf5nIoHKItQRTeOnWGPcqHAIHnAcX7rg+MPdXutEcRTd
dhHq9hdtRjh9p3qSztOEY9wIVcHHADCwBciy25fbxHjHOG4EQzOBt0SP7NE7
93dw56KHj45RTKLHPvP4DxnZ7hoM9/JNHV8fz9xviYhyyEyLEbSXIeRCK6cX
AkAdzAYXv0gNtjiJF2nsgrqDGniXU3eceZvXPteI3QgXQcEPLyxGje3wy/Eq
8LArbrtHnkUSAjgCa0pJtFl5KlOeniQvPzkwlPzXObkNySyl6hO5mbt+ChVs
PvOM8ixMRGFMC08hfhVrWZMmRpmdbB80ftOH1+1bJDRrMi6GQqWBsY2ea9Hr
JnWAjsTolC7HGiXSojmdrdzV7EGDUY7yTVe4+yjui1aymOSIX4ip0ATvGY7P
LruCe7C8y3iSEVikt0rkBhRD/mghZDcP0fy/gN4JoQiGAFiuXahc2MMegSJU
hn1dSZl5UtGG+KC48EjZee9fgyKmVbYD3KHZU+s+B/2yIBAPgcOd7cUgQWvX
BfhlfhT9JwO7V0nzTVuhBiTijGI00nSZLJuF9P9xjpXzLWtuT8xfsuRZpeCz
6JnOrQ73BdjtLl9AdhCq83LXw4sgI3QvrJAyrh29uS5zAt6pZBgY6Sicm4vf
ProVuO7mDhUPzRkGYbHKuBlwlDD+UT0Lwuo8xXoJCXM9a9mFRqfv3zisnlh0
BVZjJe8wtqrbjhuJA6P9PWkLLm8YOzMNyHWnKhB2CUIalTOyloYP5EWI3Zbn
Z10+f4U/lWUp1YhTCfLUmGNuKP9o67T0OkfuqAzWOhEIA3zHuShg10RC0ICg
F5H25NTjUz59hJFaz8tmPw6CJP/sXnYApgnESUbuXGEGsbj+4cp4BH2VAxSF
vzrjypKTAlxtRPF2SfTFDBEn09ug0H+Hm0Rb/C5wKO531dtqXI0fYVvJVwTz
n7fA0MiUO5II1GfeOQ01efGcweyl9uNY2dBgAPSvm1vjswKT4xglhE35CkQw
x9GA5ug/H88X8HjxcndrIt1OHnCk/dmIFSH+WbYrCmTWbp4OwzulEx73Y6/L
uD6dVVSTyb8EdD3iJJm8hwaEjLIEZEMmnFfxlYdv3RDFYPkGY2okcotabfYv
BfzgXnnceKmnTYtDccapd/UorPmQJ6Aet7iF0NWKJ9fyjqvsUGbRaAKccyFp
tEMxOQAfVnCEPtsYwlx0znZFZ1cKYqREMnP1OoNUyyAtlBbnKC7wLS7ygQdE
6oIJY2mbkz42fPGSKqGhCHDXQOLS5VAyknY1AjTnQpPY3A5lixm6NEc6cWrd
Y/JFECVFkuVqPpL9yAWgs31wpDJTjt413M9jlkvFgy86BOCQWDBFCaXQFTrz
EJLgmoScYeA6wRJsF1GcWfly9Xtt6hsRVOz7y5Ahnp+HvX2StyAShs3jQ0bL
YCCfdvoeXvvLiaRn0GCC/GabKz+Gd8jign7eOcyqpIwYXVYnYpTOI3xgje+5
VgUcL4QaKkT0IcDtsUIM/wzQ6kQhh+MpvagLf5QtlcuwDSVww3fZlHwBsu2n
TU/HPloXOUkUS+ibOahXwgRNsMgrm8SkGRLKPPTThmv9VsGFOEhCPyJdWh8Y
R8Ppz6w7STdsh8VNY2Y+O+Cnu2EmJCqphItgiM9jIN9q/GYHk+1bexAGkuKJ
XOtw1p3NLT+FvYKK6gSzLVtVyBbVMV2deVhcBao073vMzNHFx6x0+KJTHb3q
Cnys/OfrjPU50wIdVQO7g41c3VjkxhP2RDHqo8gl1+ANpQ3JB+mBQyM/iB6e
V7xoQei7cM+a9NCszeOSOdmBtdenO/AYWpBTQcRmXqNxvJPwBzHWYEkYLHDT
7/B5rUExQIvXJvlUqEID7C8Ilsj37dCDKiFZtaOber0V+Fi+oCWM3VBCc30t
vHZDjiHT8azX5+q71xB5eS/aIubuifLnGaQY/7XF3njIW35elmm5CLXwCmlP
wcvJf/7+XR6Z9c7S2Kc9mmmYABOQV/mI89YVb1xTUP7XArxWQI+HqtpUyL++
2PM7U2GlSY74NqhYvSsqfe91yqt54ZDBtfpsAoBpeiDuDa3pccZlpqKxYQpN
cKyjGv0xfkxiGlzridJPixApGfZYnYhAUvMODfNYZxe/ZYIFIOo/Wni3NZvP
54eui4qZ+YpfhKS+tPZckPcmbCSdyin6GBGOw3kUvnEeFn2wnUuf2pF6Nv1h
E0wrAZmeUp0cBfk49bzvu5STpFIsvfFlx5DOJakoSy8WkiDZqIkR30vlgzYh
Kkx3ee9kReOO0qBjff1GfNLhxtPHVOJM+Ozv2qstVFtt+HH0QZXmBib5+Y2M
SIl6Zj4/jWqXLCaOaYP0bSAJ8o2b286d+YR9KesyphHBnxBaubTCwqf3nh/c
gwvHKqXfcc1V1Ok54GJL3NXiA3n341WGJhcddSj4Tz8ELOiJe1Mm/b/o8hcs
8SQS43EjNUNpkYLHhONpU5ji/kdQPqG4Q1JaEulO0jAReHP/bypM4ihstXTX
TeZWwSTzTrAGOlddGMoody+Uj+dhS/E+kZ1Jv3tpz7inY7dPFb85QXrzU0RA
w9FgWhm/2ZhrrXZTrg+QOw9RCdSYdppl+J3fBIqxI6khY2mqBglZWqCURQpb
0ogARiuqQvMrZIKDogj50Q5i9BRAGbaSfc7U5S3X6XMx9X5DHArLXgzKG3LS
pb+UmHGfcrbgflVaKwb6lbONlQ7ySktGH9vlMavQnl3cnMDGb45b9YvKKUtQ
qiDdrRhr2ZCe9Josy19ihn1Q82BOVSzP/+CzyxWCsO1O2E9FCuOJgwfem4ED
lbVQH4SuQDi5vo22J548nWNi81UVnYeFWgV65INwL54X8XxTqfUJSKvnoezB
IYEjLBq1uF/YJ1uCsYN2nHvaTXo2wJKv9W5XfCmYgKUZ0YKRhYNG+L23Bbgz
EkE6FjFA+La5p2AQsaRkZpaOeNM7IEQ1aYxueeewFjuYHjc8W+qEfVPb7xsn
leo4bWNdfYoZ2nLYE5FtSDDjBDwmZyL1xuZCEVscfM1Ln4Y3NvJ6hvTjnGAh
yWJUsSpH1WsV5H0OPT7usqUkRsQ9dH4seplfrUmOl5/COmPm30ikSmJEcw0j
R+LImnchDWRGuDzVqgk3uN3/0ohKrNpJC1tiZU14zh8gGNDuoNmy7L9423W7
9occ9bL88k4UMflhvYj0O7tKOvC9UdD4XCzOTaRtdhtu6uEGwyGUXDHiEfiM
CM6gQr+NL/ZRvotFPJNcU/SeuA1jxe3Rje+BGJOZ2jyjJMPSbTdNoEVrh/VR
P5psZMuhXwhqxjQyqP3b5+AuOZ9OSUzrJr/SuVsn+IfDFdLiGspRN5g//Wdk
wrmIlYD13WP5UFVmtlt0d2V2ZqRPFp1X004IO+LTMkHByV6lJhwSx7l2WzZU
Cka3B15s/CgMNgg+ygttFjIMn1kD9srbQcZ2Mt9ItfvYXWw+U5p/KXG1UdQ/
4w/FQiEeUFz03Uer7xwDMWl6XDj3zN9NekWR2UQGea76N+a49gEcCpYz/ZwS
Vw5CNRI2sZUaPkRRjfg7Rn44b6HspyNxTsOZxmDHJxTzj4TmP49bOmAsxJsG
pAbFSVU3Rr5GwF9rlPfATStNhMA3A7CQB/S/6oz454oDBJlv8Vi2Z4j2EaQ9
f/zibv2xCRSvrm0nMWlU/BcxGNFM11PYivW+8pQyA1Alw0TFlXPg1sdHgnsS
A8itZp35Vz/Tp1x+5LQ1Z87WkVrWJxCYA3O9VPEc4t8rDY/+D5x7ki7IbfDk
RiC53KVkbWpCTmZzj/Rd2CYZ9opuAFhT3OYGWQ4UWBe26yNNfmXMPKvwxLTN
DiXluQhuL2KSZNf/FD3p2RbmIO+QuRe5Dm8oaS2JqObDpyHXCT1rTfpWYYpY
WpGC/7zn8Dq3/MAzFHIkc/NIxEXflNiBmpj6URP2WDaDq+asx886B5dLWWHB
wuoSfsImyBMgRhJ5bTusK/8J00eXn9KqPKDXQklbIERxHWSqskVdcMPZuEPa
x+avttPMallQbNrvSmbEZEq3rH/uYOb1Xtf9qveqZ4s6TA2cGjTZwnkaBjMi
XDGwY6P9NkwaZdV1sy9FExOFO/gR8TnGSzx0TNM5G5ZUhhgrHAeDrqRb7axE
H9JFETu7uDupM/FLiQ6elITEa6GAiigkqbheFWZFnrtx+YnAmmgbYmEct+3+
jv6ds+J8T28v1swtdbOrrM0Hsd90JZsUCfilXAAspXoketxD1VvNGX2Oq9OF
CixEtVnVadQRywXoxrF46BunHtb6g1ohbiVknpWoygMxoXGzY6PDdRZonWWV
CpQHKLothu9Uu8MxeosPMFDkpcERllMK3xft1C4aR05ivmBBdtJSoglRKYj1
VJi4e36xchmQHe9lUNzD5YB6WZZ8lXMsox7J1KwZGyEzqa2FH/bPRvAdD/TR
Np1/s4K7dGAwswZjd7If8bNd5rdt2/Pps8ln865fpkZ47Qx5PjrR5vJHH+TT
eb4y631td7GFhtBFC3JWFq958zSKpbkN5Nk0SZqVeldHQDAf2N7IigB9r82u
NZWvx09iRA1wWjVWhRBEG/LCdX1dPDbEHfIwpRHQuywbEp1kvGWFNgF4wqEi
W5hzqH0XCOXQHnt9rcSbuF8dTGutp1b0HwI04s96f+qSyJNzYeYTlfrBiemB
HlNru4Q92aGCqd8S+dafOwWVJpNbh2aAdS54Iccc5eYqD1AKLMqlcO2V5RFE
M9W1KpkUGAaefU3R5a/ZHg2soegJcKhuRjOtZT5JGNmwvY/HhkTqxTN4K53b
aoElMwoc+cWyFyzfgLeRjTMn+DeTbepWjPYDGFO85uOJdQS0IYiqtFKlM4Rj
HRmlFbIhQqFfnLQTjHY9PQDx6HlhQCaXo+jwdMfJMSmis33In97aFb/96y9Z
CcxgUSAn1gWUQ51SQ4an/dNunns06SKQTnDkVMztYiRlDyMwG8Zq5Zf2fSce
d2lqZ6Epr4kRc1PbXEygWRRkyen7P7LFMxz1ECgCOc9Gqr+NNZvtk+fsZrPt
YySUQyEMtTVoV2xFqubgS8hl8Oc0OCCeIf9ud3rvi2VRAadyOqBakJvALQKp
HOBfSPLQj//QRxCDLhqSlf4PiQ//UgSCqwkIZoTkjAZ+LcObDM8+aQEUVy23
piw6NTgrhPidx0zVgtVbZiu+vwrY5TMMkiScBAoQ7qIY01/XiqiES/RT8pri
Xwz7JdlT0U7MvaMiycsKUdiJmhZigZRguLePlFsOC9b0I8A7jM/GGGgl4xSc
R+tb6SfZmlKA7Pom33FdSt6oFdYwOOo1GSKfV6SAGuYg6F8H7+qiQBLKQ+fs
fCh2lptv/gVb5ewv6ScT4wYONUfTxetJSt/T16J5FU056kuS+qLkNTiVuyTD
WZCnwWTAc6wtLfDoe8XF0tuJdjOgASQLdw/BcWj2FExsEryCWJ9u2cFH6Cph
WebAsjBKl2WYaTvyqGH50LNEqO1CjT7oRGDnv+UNdz6BIli/BMEx6pb07AtQ
wNCLpqDJgdEGtPZ8T4rDS4nDxam747Mvr3MuMi81rfdsg3fIwTopJNoeMvg2
PMw+rV1ltw7EV43fXw+vt6sIqMpth+1s1V3lSXyGYPiOAivH8jTtglikCNEo
zatp1BSg0X7voCWbqt6Nz3zXxaUz6EizvG46fP5qc80rt8N1/tpBP0Dk33AY
0tikmhMbMX8/hNmClRAUCSgnHJALsNNCl/zj8VryI7/fb7eFBlngC9LU0d4G
PdiPL9EECX0jpH+RQzd5KGrQ3b1n08fLlvh8DqdqCYEY1o5XxcqE0DCueXny
4VyU4M5SxmVOE1bcjJS5FFGUIBZZswI4hxXDNZrQwN8A3XVbx2WN55g3cGgJ
QyIf2cadK5/K/QPCjZl0jXwdbaXQR98ET5irvJAx0Q4N9rFcVYxhKDr/bTsZ
J31kgs21nNjYPXAEcKG55mXqv3xZ909r4uhQfmGJQt+E+K7s5Z6vH5j8KQa9
uCYNdlWAMBXgwPpPrdKXCl6VVdMAgPSamISn9YqSnR8Uq/uouZZBCMllxjjx
C3vB7DK4fPxwT7KM+RCv41wYYJ1hy7QXjfCMPXgBLGDapQ8vVBtCYh6dTxMC
E+fU6bNhJ2kzXx6n+izl2ItybwJzH/R3qd+66DabJea3WtHLrtN4HeTl2wT9
k1TvkTj21dURVtJJXNsbyqxMKLKUU6g0p6uBr23TDJpw+TeSD/FwoeUxb+Bt
5UtEFk7Rdrvb7f6JzqW6YJFe8T0JadB33LWm+x1smtVuuM/taQ9t3xmdi+Am
7JQ1mXq2+qcGvYXGWKm9WxrwIKMaOfF9fVe1bLuLG9PXV4LPV3najkDePcHI
yK3+iSVX32yYOqWTJbRXu7GE5+fZ40tSwTXqYk+/F+oOXLyFSuOtlTu97FfD
gTwxFfDnNSVY57qV5GNVjQk0cD6swmvzvu6eVMBtZswW3mhmtASGAGHcFTow
7BapeV6JcEjXYLU/blZBkjmElz+RBmKpZ/yqCzDig0R+mgJZ5tIMSwtYJabn
sT2X8/5gEOJ8gQikiUf0zaou3soEAaUNqszXn7lXRns77krWAmX9LrK71lFI
qRTbMXx9vZ2uMUFQQW0IO65UiL9dHjFKB/7E+YS72wVlPC9+Ia1U4zwXqH/Z
Rg1EnrDi5zRICyM4F/RMMuUwI3z5Y64F4L3bKnV+KZ1+fQhOTdKddQWtQxPT
U/A+zYpw3IduIGslVkkaUJmfJ694SjGxonDODln04g2KVNDCoWZU0cXQ4x/L
1MKl0UrlQxZj9RTK45mb3Amri3nrt76Poz4FZ94Laq7tZyPxwUYFqPWPavaR
mA6+oactX03ed6uMgD2biN2FQy2hNqm9q56xTQqJcZugZA0xARKXl3anCuTB
JymM2HAmjJwVEgfubEUasQDLd0k5I+XdA/liKchaBv3zteMLnnk6xZUcHtKD
gZ2Y/LSSWpkzL0Zc6Pe5OutOdj9v7nGcjlec/qTbMMBxyjgalLyepfotSW1z
EfmCuMltQmNz9sgjum6NVK9xpkSenEn80k7XTjR6pCEXtBPLqZCbLZDAF87y
eV5jjpS80e40ZC9ef7rolbMNcFLWE9mKpyEgO8wq9WHY6Vqtv/sX0jZMQPq/
ivXs7vv985uuTTlpBJS2Tg2XpywchRNp8yCm0A+GzXO7qTVpQ5684FQd+j/9
OOzlZPURsPdMMJ5xFbHZlezF9ROg7IUzNeHLSlON45Ki/jn1iN1vLDawDmtD
QNPZccGsi66eV1VfP+zZdDBYKOOXns3hqdUbM24p9wMfx67HZ8TrvT+UKjDT
C++jsCpZBPT4tyx5pnf67oyItWyoyZx93qMx+RqY8hk+GKWdCCGNn2e5Df5E
VIUv/3EMo3wSevJNXkkjhLgtJ6y+HRNenE4qnbvta5hukW6rv9mxt8QWYPcl
SEDRi2RXDNkcZ1TEkyTzRtSOakQ06gQ59TSLMLki5Q6E8d5HHIjEmQn3h+b1
GEoxJEjQ5LczAPtYghkscwxsSnaMBf+Wme0HDEZ4B2GD+pNFMMC/Itl5zTGN
3lefJ6uFHEsDR1wyIpEZXoZwEmbUSogGYmvV40C2xvstS/B6Jpk3F4vuhIPh
P4PXzCDN3Se257+bXLMS5uYn49X3MK0j+lUjq+ogHFYxl3fYdsCI48TeuW3E
qr++Qecq0tOQY0qGixYh0e5RZ/CMZ5fPgGxfuS8fh63xbHSwLY+Dk1tM9amG
Ur8wlRsymF5ajM3OuIS+WmyoKP5OKU2/+zS8Nm+uCwck+tYbW15HC8VnLriO
djVsxRLg2+oODdTwES57r4ezxP1NPPf6Syt+IP6IUvxRQsnAJj6BEfhElqBG
K1Avw7mJJGi2veKu8DDOew3y44s8ormXt/3amef85hrRDDpnEKVSUD0SoNOr
NgbCx4x0tPJnB+Fz/wzJ2S+rz4vQs8K2hZ89XnWIguCPFPTI3bUaXqHkLp6A
dYkpVMXq6THuLpM7c7eHKzv+0n74S45xx8R7TmhdPcH4w5trGdDtyQ+SmqPA
V4tG9HoyhlMt2I+i5OsfMB7eoKNkPzn2df2UtHsZs9Q0jRDWEXtb3uATqofR
SdpAS20C51bxr+NuwfsSaaxHQxYTn/ZfYq0S9w5ciAb0EU8BWxtdR0V4bOQW
HapHONWmt1D5Ih9PkSC7PGWmsvwdX+u7Jhha2Qs14SlTWkRfXFAb784o4DZ7
q0CuU7z8cew/MzcBRJvJ90wWJyL98wL8z8mx/FFsEb9RVLlEVVZhKKI7qBR2
tVu+ie5aSWh27rQy1LB0QI+uZT1vakpSPI5iBjeCtIVuj8IMPMsKtiKjrH3H
XnYufo8kbga1V28C5VFjWM6ZqPXuFmdr3rfZvpDNTBr0H/sunLexltblcNpP
JwwybgTHWQo+/tvcT/cWWEIjqWN9TQRKtKk+LVkcr1N/V/nXloSBzZBnbmsz
Yb/MyCW5flauEy0gGnqZ4HwHJT9nP4UBMFYtxfm5roRP4vh728ATjHs6lNHG
nk81r2YwA2VtrUeCmsJhMpZMWwxX0TIz069IO1aTEzKqUr8F8G5VHki4LDHr
CZjL0FFP9wWOE0yIcQ2yy8CfgPAyEtt8rGsR297kBQSxDgUkdvhZ6SuJv1vb
2JsTMR2/INTijRrhGmoIxOsLIJuu1/ZwK3Da/sYxMXXLd7AeCVZwQdwhyWr+
rNvAFO3FlEyKsH0NJadfYwbIqCXfpOVnlB4MioLhYMdBYtUi4ASy0Agfa8sw
Vw41gCVbFk4QT3ZPSNw46Ozv4CVV9j8fr0FZFFRPkMhyzYiD7x20zn0XzsMC
OsmHJLI4GU9qgkXMSkNxss43UBjQIWso0i0qvpdXyfNBP0VYr9n36HEUyD6e
2CEaV3HeKrCTwSWB9AUvyWda6kD03tRpLSa5dxTrY2UdXG6cdqiAVXUO7fuC
KwuQmsLHn9uWUXV97a2evPpItEFPneokUJ53wjAxTHTkX7zFZrHWCV4NT7yf
KFM/rTOZl1ur1oob4UkXXWRb3r5Aoy1PhUPuYbR/R268GKmZMGvPMRoBn+hW
fQi7V7HZztCPDrZPdbjsIP2V2YjcjNjYE05F5TsCHRcjwmY2Uaq3DFRqCUyb
fMHBVvNlJCcynYZyIxtk3hS19L0JVdrKIIet41vHTg6w6p9r8IihVRYQJ6ar
MijzrQHYo7i1A+XpoXMlS4/tVgHcr3iTjbJG+6sNYefnW3UccNaG1Z6gFirl
IZ9sN/jDs5KnNlVzF9KrbpjC0uP95yIuflPTsgaqCrp5omPUeQWwjobhgQNy
NyAmEoIP1oAHBZpahRnwnBhZo7pW6ohfYLY94hdX23pQ9uC5PYei+PiBpG2H
zMSl+fmd0GIwOHoDOJ+SOU+9GYAp1dmV8elSUOITdMfeo9dqXP+Zelx649h1
4MW1e55xIOzPMdyETrY8/7aZbLaEm+fNWOrvjx5JoyLd9uu+8SB2wvtr74oM
n7Ith7ICOrPoSsM0o74mCtuvr6VnKPkjL70cfI0PBuq/u82n/+2+Yw0OaxB1
zE+O6UX/GYpOTWs3U6+NkeI/406AQr7qpPwtz7+qOZmfweoL1TXvID9B3TKq
55qz38QytfX4lQj41jW2UNMIBaFvlZBlJfsNRh88FRim8Wv9kjFaZGj/B2OL
0aW/kjg5yqakmgOiclTqzp/SKgpOCCC17xPBStXFfkvHaCA7ytICYAdpSXen
nikyCdNCse1sfKzVlw+RQ9pwXxDOrky8sCKTY7BnyzZQM+BqVt/3X6P69l5d
aVTxF5q7imWPz2JNs0P0Gd+IbJ8u5dZ7cXIf/UzsW7Xct6wIK/hPUi04e5a5
jXGtHc8r4GaJEd8dJ54pJp1BWNTMMp85lLhtHytY4hb8NcQ1eXuOC18uzgCw
atZfnqeZIBV2qXYS+RIzycZAG0wr/tNNTauphY4FPGCRjoUKNF4/jPHo0Zqq
YlrVRaw5YMw/4GVFQU5XwwdKCP5CZONmSBljaQ1+Gwt7lS257YMOBIORszTP
UQ8VEXOPcGCD0qk5mQngX5aoXl4flOz/syHkc5goSeYeXV91US+spwxj05ad
xoQ+dOzei+GAaSBK6rejD5OhtXjYyrKWeRa+5nZHupNOt1AJbgsV/iNh0xk1
VcvRPYHgXeqjVLWRR3cV1Hwm+C/yvJn1hdrUsFuH663yXDDSDgzaWub2oJRc
hbzGt2BW/IclEJ9xByEZ2IG3bFcTTJWPfdhoDZK7Z49/42JoTniloYlGmg2p
kT4xafzsh32p2lmlrmhrlJ05qmzx87tmbhvR4OGenB24dVrycTmR3Red1kFV
SKjjxmQefpI/lGlBUi09tkJ2pDWi04X9lKk34fx+4SO1q+1hYX4n/WyNVfp+
hJtc/QF/BR65GbQ4G+7iULR6Am9U9KVWb0LiDyUKUdv0VRuRL6gEfl7HgL3n
RNCJN52/sgYK8FDPlnz7vGbVL2EKihpwZUiCn5MtM0pJ/IdlkRVT32pir0Pm
31ZcwN9C0ooBEmtqjhKmOHZQywd0qCo64v3a4tp0CmEyodQuDnwSoMIhGbRO
BSVA2vWO0slDA2JRI1O2diQtMaArwZ18nUr5fnDNUgAIG5edLsJEKWUv4lIp
WhlJJZXJLSG6TpUvQmSd05haqdUQUEfaY2ISSJmZeVeLxJc6XU57xmCS9yDj
gqzz+INQD/C7J4FBuLuH6YrJTENjaIZkI50fJQFzoUlNow8F0ZPCUmYJwhjy
JCNZfequGlmO3p8/dvobLZG1YowJ11u3CBT4eNLoM038+h+azW42H+QY0K6j
1vZSy6gZMrZWuraZEt46ZCZArypQ8pxc3gciGikb9T9EEhSJLSMoXLUJFgZ8
syOclIMkiyeZhWQTx5jGoezEqoehOVlGowNfdNqyvg3eyQ7nXfmDSvGnNBEo
1xfwrGndUGujEAX8tCR1mctNlW6ST9xj85Ao2hAf/xjep8nFtx0o/EJnyafZ
4HKorKfet3n6wYfm+nEjIYfKDCiu0linGirEHi2DzF5ZC8TtnOYSUEqKG0lo
TKTPmlZKMrNkn6GfdksCPhaYLgezvwCyW/goQZFEoayIwiZwNwnjeLdkNyZF
WIj1z3evnleb9FZ8ZwfZCgQeUExJuUlLB/84oKWShVrj6WYIyVrBq4l5PhAG
tbZ1KsL5x4Xn8rl7mEPYJaL7naRZIbTvfo2vxMqQPMP4+OQ7SFWUkMuO/2GB
zNV+XF0ORRqk9NTLwkuyIgIZkKb6wtXkml2P30Us0YNaLpxYdaAFPNPbu936
mbBP9R/wigKcvBc17wepCgj1RbiXFvH7ZzlKdTQ9rtlUNDQcbEbI3U+NU7EA
zKv5+CN3uHCeriwk4Nbb8427pTPxjHc16SwrsoZlNjTG+05npxQobnmjYB9I
3hueVfCfMEAJt3mN4oI1KADfK/0evxAi4AGcUE4NztvriPGv2d9tf9ftgOp/
DBBObEbond8vPbNwD5R2nwUDw5ZB+APlLvQB7nr3Hrqw7LqOovomdN6IgZ6h
fnHDBJvMYQIoKqKbtzcP4giGfzNY72NAXkkqjJoGDErfZRDpVNVNUq0bpPvw
nkZUiA6FlWMleQ+VWHUV1FfWXAzh8t5tQJ2DBePREt6/2Qjh3sXUhP3J6N+8
/pmxvdLMZ1hde0zth6xfQ5PK10J5+AB1UWx72mEn3lBvRXsIWo4LLHicm6u2
cEEOWZqFonzPRAXdQP8/7mXB7mSyroovjd8wv6UAcM2imqVYI83KJGbxEwUh
XE1meWEYrBRrQotwYS00LP7OAUIQ7B8tHp3vwMLUYS+dO4KVooVg/rhidDiQ
iTzKh3GTGGQ7ZhH6UA2EQangnvDSPVY7E/8b+RQN7IBN5DWJzt0j4JfAQbtJ
Sy2MGe/dDE1txCyHEifovcYh82q8QCMUro8cjYe+iKXsNiWF9RGMm05McWgI
LT6IlHDnENLsLXISvCPg1cFg6wF0yqeGYm2TKGsJ69Ugzkjr5EP8zdn/kzyq
Wc/XSanXlXfOuNPVvryz93zJZZIMAwHEWDllmqZMPe9jhyZdez3NAlz8C4bx
VhFLEpAmMbHLT98RVq7q3TIgU+APChyXUdNxQYCZMsQ5PiV8YcGJpgh1kljN
RX7XMsOCnHKnEHlyu6m+gn3xsSr+BvnGF4FZPwWizxfeM4wihgKRKzPnlnXx
ytUn1t3ORZFBtMwRi5vJL71mjv1RhWR2rnQuikldXxtttOSnz8w7raSPrlF2
yVoDa4/9P0NQ2TDSMb6A+VCBEWqf+/tAjA3hiGAHYu90z8WbUDuElAo0ZOc9
apBz8bgoqx2HADA5MsNh4yNhxEJpiKjUHDdspFtMEv1SuOFUXjBSAbMHZqLR
+QhXZAYpVCTxPti7qQahXPDz2OlPd//8RtDhdIzp8GdeZvxzcMSg2eyWCbLN
h2v1vUHSi7poNQIzICQAw8QDc+vNZe2aWeh6s8TxWTNUdXQULS+LThMD8cSm
Fw0RVjZzK9+3xb9IvfxDo8OJDNKpYB/KSHb0hlW+ZH4MjUqDd77Ym28s2qLK
BX4muBimN4rjf+3wOx49wUQNT2VeFbFJcl/kEDWYyWbXwPyAADinpRIEULDR
vusuDN2b9u/M3kVhSJP+oMFX4Da1QKbj/Omti5VwBCN0pUovm/OrAfmUx3ue
XQbAO0zISQEGd04tG7o4CK5b7UwhS1FE46LYjrbBL3PP0xWkj72bNiYcWZfa
QWG60TXu1PE9y9MhBSkdh0c89mq2CrIT507U8EYaWm49Z5nRiUOVdZLGh2PN
9fgExBj06PU7Yzn+LzBXE36UmJHAuhEfKyF04ifXc4GKNaGbSsKick4Z3f+Y
2ODcleimEuRpXlyZhXOfXJX9Zb5dqNKUUv1o69mkjxigsmRWmATPxS4VIdZg
R+FRg3uPLNJgw6mg267FaU/bEEG6h+LzRe5itbIRnkA6vv2YrUGYmJKNTwH5
bHmtlSqjXV1JzseL5KvQaPiywuNfF92XJZjj8Jm7Ju0uCZvjsFOzRZZmF52L
WkVFG3W5WMOxhMHcnrz6znA3efIn7Q4CEPeTCwqUw+hukYqDE+mLLVdDRD35
MDzdO2C+vsHG2HvrvEJOvn7nm9zco28SJjc7GuppIoZNcLWyzOQ4GzfvoE/C
JzuF8Fp31CAz+xXD83lEF/VDA2/wzSC5UjfuBdgCuEFxq5oopP3mEz4e+bWz
oVcjUDQYEcPq6sB8nteCeDJXe+GhXKLmD9MRHbZORtYIdS0xvEGxahCo4G+5
UoCA4AnVJjOXIkDP7kXy9hdFVmKcLxcndgZ1zii9o1cm2BphnP4OOXKtJYnc
o19ibLt+8MhQbDL6d+9PHuMdYOCBlvKbkys18MIAluBRQ4thpjVOOlC20thA
jp6Nea/9Ew7FF9x4Y/S3TWabGh9qy5rZigbFolIlbvMWwd5KgS+9mVtMvsSx
IorBEercGL17EjR90dLIhDgZXsLdvrdcq4HNtN5CAxqvu/viIWOK3zaYJVv2
hRf4PE3CHVf+s+kCASisT9x2HZC6XquYf6pGNMT5QcavYP/8Hfxz1X6b/IJC
ThAA7N3Z6lb0D9sQdA/yaPddbgJTjvwRtd0gC6fTsDBSDlYSeA0e8WBolm/w
tFVlZwGh900F+a1eYUb/Lrn/XcE9zhgaqoVQ7DTJvMoBl/2cWpFgSG8V/6P/
bQK0qk1Ejzq8qM6xc6wbqqzxAN2vCrfPnVa3fHlurEBSjULqukUgKhfvj48C
SAt4HXJur4+8amb2e4t0tz3TeVQUpO+QmvE+xuleyIXWcA9R4eaXLH3OKeGL
lF2jvYxpxtDLYmfnxqvALdcvJWjreLrKcdaS08I1u2W/kKg6JjQhxCmtvh3v
h9q8hFOSz8UOLStP+1uYnScY4N6QPUHsb9cVdPWK9d5ASyXOOE4Jb157r1Zt
0bhagS2Dg8OdhCCp2bs7i1cXOD/U1o/Pvgn0/HNvG/x43BbrGk131ViJhmPa
z92KzmR5Cclr/PCSzUcCnuGwTWhU8zm1h6dFKIuYE7bWCpopmm7OGycO+C3b
1OsfS3gGKBrT3vc3NSqErya3h7cLIHDPajNHQg71Hy7J9Fjt1h0bzivMmzXa
ThrKqa9eYS+JP+ti/4fE3f/mWznIK7wB9DKY+ADaJVn4XDmBAhKkSsBj/mgF
tGlxc6QWMDgyyAHTib7NG32olnafWAIGmx+gWxLNY2VunujZTkmo9jw1Tj2C
T9Uw0MUEdrr4dnT+oEmsoNkOpX8/PEGnZc9pBM9Sp/kX+hq7Dr4W73aGyAmN
AiZ8dkx3HVwtJ0bGw0sjgZXlqfumO4eobTSgk9rRGMPHCeFP8J8UaBHn/CXi
TVGowI/3g2vGk86fXuH28jspoRdjJzfj1As335ATL7kly7RFFw14Bwc63weF
hiueyJM+eVCUHezrtNJ13IFEDGBltuUlCaOhPaP1NoNVmMCmzE1rJ6gvMT4V
C5/I1olWcpeDqhA7fRZ0yhRgtC7kF+ZHUZL80hsR/d3RsodXSFd0x0tm6aQ7
IdpFEQOvMrHSWob+TMeZKtawha+Q7EuihftzfLjCYsk+sEfvBJNqMSPOb0AJ
0NtmA1d+mcYlj8cS4tUpORUXDRQRM+xA47E2KRxA3lp8l8DjGOM6qZ7EN+a8
CRRdKP768I3YfkkI/bDkJUPrHZlfyrsc0s2wHW66Y5MgLQoTUpYOmNWRGQ3U
IGF+ftGi1hVyuOwPunbfD05pC+L136JADP8PKdz8poYbgFATmN4McDAqapIg
4CmaHHeefbJZt+HQeQtDVkV2RXg7lciDrgtJZnCAw0nU4U2ssaa3Qbv1I+2Y
dqnPLYuhIeiT/Kmy36+keFUE3lrZdJyldPDX+fdN2DA9Y04XuK0uczDpleTh
DeJZnjTRvf7ndtw3qlMnvLoCfAH1dgQUzpGeLQBwJU1uwTznJnEoL6HnR8PL
cRRrtEIHdvTOavHvJ6FlTM9tv2GZmBcrI+DG//KxYqXYkGfTGUivRa7UULfd
RXq87ds6h4h6WRKde+57N1Zvq2+o+VFNUIkQrZ1sPNrHyYAE+XwJU5atPsDF
f54pFPl3qzrARJ/lxteT2lzrg9eWDNZCgOJea+3wu51akOgE3rPFofDS/tPJ
+5krSA0d+W09sSYD2dbQvsLsWk9BYuEWuM2FJcoElzIV8J1aKwAAto7Hf3Al
YLh53zjKEX13KsCOuow1vSrcaZgeOX3VNlHhxtG7zo9hJErOPKnWZZGnD9Dl
KIBaqQZePCEbEYyHkSV3DetpVAckYzYsWtFqNadka4LhnqmqOrhiAugjNjsM
HPk7Pbt8NtRa8UGPHzIkHvrAoT32jCqzd5e/brz83ZFBooGNavRPXdwCjUNa
zvSOXo7pOX7mRSgeET0UMr5nSDvgey8JEnErD0BEJI+w2FB1tB26buXsMp2j
M8ugm4oHFeUNyChES8YfANoKw6j7VzRJ8pGDNbaOeBkxIrYvkr815qkSjvTg
Mptm1QpsLBb/afugh0v7tmlYX/u5bTDp45pteB9PlTOeGfyUePfbKTEKP/ki
9w20g6pTUCZdSczQrP/GfXtJvdm3Laf6uzauMgwztPNQwS43u5HurZHDeBcs
xskVvB43k3hX2/EZfpsaXwpeXyjUW4zC/yD1tQ1o/d1NC+V2mfa+PFKMNSza
3tfGHPulCgXTAlgsPdTG2PrCBNGNWbXjbJdFiWu3opjpxqo31ce9lGFjaRQR
kSS6flG3mP/hj/+HPbojh3MuwgS1+mF61OCGSp4S9NS257O10YjATied5orZ
Dsv53JHv8OOaD/oUONwnMWFA4MkCpBBSbK/yukV+5HQJJeIgGni9PaEhb+/X
RZs2XmSeM8DtRbEkE5Jwfj1AlTV7A4ojWrUWRW4jmVwsxr1Ht/3CfA8QqH3y
jkoHjlCTJacTy4MFPIA9gLSudAo8sqTzz4Fplh/zJEdrPAdvYMWYNiB05t3t
LryYCJY3qeNFw9MUZZamr5MYX0gpdTxhdAfqadVfpXvYZgQVVJuaiTNQUjG+
AAAGdL/AjWQTwRHZ2kQeIMhm7c/vQtzPvlTJ1c/4tiIwOX6JMxVQ6CEE1Rwm
ziUx6EsFsBsTR2JZK/yxozDHwDAAPLBnWCqaZJVR1ObMJf0FkMHNzRXC3RK2
oayDjhcVPYMsyRa/awFFRKjaeiisU3VTgiNfbeOYfO6GbMeFbMSRXVMIIW6j
i9tFdhg1Xv2Qe0ggTNi4Tx4KFnp6m++PWeoJIdSeLn/v6QGDQanQ+GNPz/t2
/APqEAHgq4ApRUItIlQ3Y63L3eZbtDW8EzFwNz9i/uOpztrqhpP+5Kj/xneD
EkiMHuU1WDzAGI/gSDb8Z+WSQIwf2nASYOhgv7Q3VhwvY7tS7+H0nQExpD9t
h8J1Sin4QZyiSHs03Oy1bxPwBpgKDJ5cvee1Al+PsxNCz5CXikhydTjQ4sGm
ekh2sVydC8cjAmixfkbYgBmSFo89f3l11OavCz+oizDb8h3fuftCiSbIzCJ5
uu2eXcNZ0vHNK+C56VxI1WC1KOF28zpuHUTp+BhIbObtGR6dzBQNs6/18Gex
7lqaYXoLrUzXgzBpAnEBVP5hHUTIgdgIuNgtVl1/L2MQduoh2AGlSlC2t8A9
OTpa/CWmiepHniAgHM3p3NMopQsvJV3rKtowCxfg5jltsQBYxZP8Ba8eAMUn
jdyBVekBB/QJSjvBUxLSn4xjjcSH0ghiluhfrW2/LBTZcjH0Q1VOeXawoZnJ
+FB0R+ZqRCo5yNelbyHj5bUDdwqH9zvRc7BPAusjZetCsbGUPwT1nfu/dMKx
t/itL2ZpHbGOYuqbVkOyiiIKHpTHUwXoB+sZat3xtWQFuZ5TouoPjhNnXiCY
ajug1pmmKDxhjMIgckJcvg+5OejexxQd+Rez47eZgBLukEE2E+OKXs/zV709
Uu6LJRkjWYT/QjImIqQeO5Hut+xAr99AQA2RSJgoxrr6Ly4XfHwoDTb4Ldyr
0oeCg2GUJf1urKnM55ebNNUnrFaMm08ZCSBk6QBthiNTOfuPZJ5lB8Laa9px
aaSOy2kw0RM+mNcQ7RG5r8M2ID15Cms6iV0kKAk+HKA1dWVt3VdEPYKwrG7h
wKm2zUJyo+F5NiHCeXFFk4jWj1tvIWv06XZF96JfCnE1tRklzx2ZVswsSkxV
irpYvsFs640BgYZZQQkQN8eKWggJbi4/9pdsqr6Jir0z1HTBkgO74yV0P+2i
AUsFUiapFVgbZmz7Y/BzMlWKyWD1q0LZqcmEg+dRxWaMW3aRlUqcHTOH2FP+
2l7i6DO4Fh/4pRei3GMFu+sEo/fVTW+22qioQUaJVT+WFhvc6BD1EkPivpCQ
Ks12i4IkDuUEuzijaPHGuGe37JTPEq/qa0E+0TpXWwrKuKStWVVHw72xX6HO
ncXS9TujZzFynDDr/rSXGSlSphzLsyUITjC89/XcNFWhD9+0Og0qhT/QD6SX
SuU2Ag5A6zxrJjtZpp3JDzeO8+esrydAH4x10dIRd9n5KBaZGe6PNbTBvAuf
YW4ZIiUFH+BOJ4McJ+nbDt93qgIE1xLd42Kelt+u2eTWr+PEiJUYs9MOeI3q
wY5MYkqzdcSPQNU/yDVmisYL78zez3tC91FUiZMxbB/TRjNBSMjRQ66ACjkb
uGZnkE61FuWCUpk/uRD18xwSnaWGuVp8hoR6eSQnvDkAv3pXp9BJ5xoGpM2m
jzCLI+HwaGu/t4aPlm+fxEofa21M86+9sWC2KPpQYjDVXsDkTcEigXqfYpU6
yWRKJeJCDOxqrDLgvxP2014SBwEWKvyiWGKi0T1BuH2IDFlcRPagU0U4zkuE
aFuaFHmzM4R1cOHz/SH5+l2IZm39e5L/FuBBVnLa3Mrspof+VyjUgPfvACQP
VKjHHjotSJ1GOQlIiOa6vtaNpH6+l2E5oJQNrQ7HTz+GOF90iC8iRN5W4Wwg
d+GJJPxgqpecjms5yDjIaVc2qxfmrnHfKaFXpqhjN8CWrMkwBnPGNm3uefxJ
Z5ec+hrf2yPi1X0udl0Akyk6nntXJcc3pitb6dszbML2A9pcEMUzYu1nq0BF
xIWQ9NF0+VvedC5CuDnbH4Lhdgu8FUN5s1JNyuuV2YXf/+Dp1/CItqrOc5xg
S2bPp8hD0dOrqv4BX82fhD2ruPXoj8EluugbFsuf9insogFv4wux1OtFoLc+
K42+uwxtbzQYhg4HMCP1hFDudB7hPL9W4VXtPOxt6o4MHVQWVbP7qP2RBWVQ
DRbYlABRGgMVcDczcHoFOaTUAamGFpWyx3QGpO8bCQaSfLiGC/cOzNO6d03d
ciMMat7zJHOUwT+wMZQlilqhsriwIV1SVF9lDZnZCfzCqrUpV7/2grtS1aZ4
gUJK/FqwDkNWlw9maicTxP1urYgCZnDlOXkILLOyAaKqsD85eHDoSef9jKJH
7HmyQnTLL7NQN9dszhrc+BAu/8OQaR9NyOh4+lH84b/6tG+GTgFzSdNs1dK5
EDGzxqGa03uB1Ckf32VBuIfbJxqvBWctiOqMylOWHulYTRsrd4U6/kgofZgK
Chnlaft+bQRJ9te0zB7vAiKPHd98tlOA3ur5hMBf84u3cUAY7EgsGSijDrri
MxuPMcPAsLv0BkrVqnEfsmbu9RfhDAH77WJcmK6T8eJYwNs6hOlqS/sw7cbt
RSOg9BuILj2ps3GnZUpVoOotQ5yGihNkVP691zlSUoGqQUHSWlcteowLrBDQ
+vQdkEXYNL9uCNz1lEfo0Jav1enYs4D2E5eXc4LO7AuvQRImTUE3xsGEoaop
Wt6Y344e0BQZaobhktH0lCcdVj6sRl0IDgq89Ej5mRCRQXgdMJTnw1h/emAn
dpEaU6wuuihF3cTW8bZyW48UwY1aKAGp02LRUvJxPBr31Y4szl9YPidCInex
JdaMR5fRj7i2kcWELaIXC2lfx8qxclnNr+a2+sTPtjDvu8wJ7lmp661+WYU7
3cu4SwSicCNIU0a+88MYIeRmAXueFkMF3PEv0qRTAfr0TIRGTEpTl+snIuIp
JKfTU5E1Cc60Cug1IY/y7z1hDcK+jvrwC2Wq44DP7cGkRmQs0vyLcFBILtYw
5ihMHv7pAI6r+eTusb/vjKkPgyx/QpAhU6hCJwzDmXa59rsCZ/g2jyQMPVxW
1p9oe0WIQaJO+RJlcGy0/XeJ5IYeFIqHVcclbmOz9/A2+AWddYsZLYnvwICX
gxa6L05qoFJFqeiLkO9wxIdJtOFD8yPUPQgyWkHbuOnN0VL7d3lDmON224xr
U6EAqEFV/ywrZs14wAp82iYZ+goaWKHsauLPsSm7a2C1YjysQGuwiU/HNqj0
Gde5Ouxcs2StOrcup6Fq1WC3zKdCbAyDAMTVVY7YiWMKHsN9ERcvNlCeDxzp
Ge9PkB/oYU4zgYse0iY0DkdmS2YFz3Qzw/2wjiY5LWFwuRxQ3vEwTcg/lHSL
kdbgPEUO9kdhR3PCuIwTDJjDO3zu2CYgBqXtbijfDv8P3bQYOy2GxGH5WU3R
D46DlNxMh2RLoIy3rkxwG0t9iBOkpZ1DoDQFl9DLAjKyMJsBpjdS6KIZD+HU
AetUThev+7p6Y3yEU4xn3L/AfHp6kbcRmHcJxeSCEjyBx06FrvaISZuQAqte
CXVojvyLVvJFtJo1Iq26+8wwUpOSnl+fW0rSX4IlQGuyDk30caHjIkRS3m4C
wrYfP6QpE7RRQvGHhiyWWDTr5zaGWHYUbi0BSt2y36/Cbz3fkP0THTwR1dQQ
BEekAkBgkt8gjaNmKCNTng1AVOaSLEAaymhfEutjYjOVtOu52FszWULtLamg
irxzuSh5cnskXaWaEov1azn73kM7jnbvukPVzAimzEe+yfRNXqVQ3fmWJe1k
b9UrbrLBImr2Hdh5DEW7TfkegFg4DjM7uHMBhXSiE9VXKvjGJ68TI17ZpSvA
2nIuoHCNj4Wp++FtPgsby8fWEmCWRtyiYaNKHmi3qzqSCe/PwxAKMT3IgcUs
5FCWcXArGdX9tFJ7kphI0gVRDsvP09wBwsimI69IKT+AHyWGG302DWOY9K/W
g3/w9ZObKs+optT3auU6Alad9q57HeZJc4WwpmfdQtomqvc3nZQ/V4plDGPC
g6rP8f8BqaPBWaLMUaeGB5PUry4qGV9MC3S68SUsInjb+GxqQK+mfpdN4s3q
f6K2gTbdROULzYNooGifOx87EizlSK7jr7sgP0tcTtz59FZNWVGvFuBZgPh1
RzNGP3wgisD4rY98Zn88+q9H0v2ys3eJgvdZ/XEj0VCTM1vbY7pxPubeY9sy
HYct+RexZKvqqW1TQp/j+MGLFU4/QxxeCpHF87GoNoqUIg/Ti/Ngbb2q0v1y
KI83NwRTnEjFYcfnuxi6kX8WQ0T0OlKTh8uhInTm5cycU6fO2YFaGqKsEi/n
Ux5Ew3B1U8Rp3PrOdBy3B8muyVrp5ev5SZN3JhNc2RuFsdHSCkJmXaSatVew
P+MHGg+EJIXisdEBsZdB1mKS3earLBYOZ8VGAlBJXA8USitqalFjgrg7Fxtc
XygUOu9vLcK9V/NqFctFhkM2/EXCYNpU97v3ag1p37Gd6YHbfKdbrhz3lcYB
g0M+/MxRFE6r8D4QwgF+ELueliPx1IuE90a84ofIohr2atxqrJT33/1PFYlF
Fg1+lb/h7h6wRUZC+y9GFtqFlA5EbUOePaxSoqBs+RGJ5Yuvu/LOKDNEgQnL
JQMvEJCUGZO+QR8zEbETSIbutigDgQN4eyupHkFTLTaiep3PiX4gf6gqGJ9W
Hx06nn5I6Li2RKhSkcK1zo9eCmo67W8HiFb3EiA0DW+P9258r1ynJj1h026y
K5+f/coWghoAvZ2W1k9OkGlhgDCznAwXVz4GwiNwEmBXdCuKLUC+8NumVAe/
4/cXbUHQZWa+vISN7pWhk4Azphxule15ZFUYvp/vCAYBvm3vpVvyzgDAaYqt
BXwRiY129FtOtHwlUnhNBJPQGoTECQGqzExDA5txAkFc9Y/RFjgwiG6wmsNI
2Gs82QzgzED8f9mjPmMW+ZUU0x8KTtVrZATEI9oP8bZobJdoLmr/M3aQstkB
DVHvFviwG9UDX96q9aMvV3k2FB9fguZtM4mAQoObigSjiHo02zIxqO9w7J2c
QMY5Qn+kb3/JrgnZaB80BmyyW8LB3Jf6bda9i4hYxrYgQoJizjqhqeL2QXpw
HZEMmqj6grG2ucV8n9gSykAWmEtiSLthrurGiFRR+aXnTXr9aI+TThGKzHOK
CVkRlv55TWGeHR4WqCdJ7pDIY3mQgyYX+WlM8XkXjmHepML9UvaxDb1nPuaR
/Ky9znU4XnomGLG7VLj1wOIVeQGlmr7GI6x8vc2Tlx1hABl8d7r49q6yM7MW
fRuygS645vSHx5Q1EA13qIPQ0JC5VjASniz8dIk4LqYXLyv6avquObIjwKTU
5l3ynYfS3dnX8nrTP9T18scvYWJZTyO/3ipR8wepwCXl6eSvodt1f7Q42ZDF
JHh0iATMecqMjPDn1ccTrv/FY6sxCNvmE9ldYFT8N0mwJQUVGkERom6sLtMc
iLnLdPYuQz644QR0PT4hVyoqMxFyWwD/TKUW0eCFKh9KUcWducxWhALHVgw0
mM4aWxA3rea+cvEJ8oFTmSpxL1uKKknxovmgX7vlocLPMHmwr8vMfuth/gB7
e4ZGIBeM82Sc9kkMPxp8ZcR5W3w3Bt69GB6254c4WoJYNiFcBlOn0fCqBqUg
AbnJkxSOKXfn+XLO/4TLqNmWgBylw4yGcSpfrllEMDbZdN/mCbGBAHkHa1mr
TblmXaslC7Iwo9JldpZh4MfJEGIzDoOAfsLGJ7/htjaUqzdXuMfrYga3d1Jg
Uc4Lk5cQUbiMnEgMnn0NDjIh6d6aokxRn/Et+P/lMi0as9sAXcpVgLcPgCeM
oZfJd4FtR29oi18vEgWvkJngkJyrhDF5gg8wuP3sfBUNesuQpfWnV7+yOJ0c
frxJCOlCk/YHQwCdivUe7kLX/zhoS2BkuLq6jJltHm0YePqHKJXVs5VJmvLp
nCPvgEhHTzySw4UJzxp6fSoiI5IsQFcYcvAFAx3lexIBE4wrabXVp5IwWD0R
V/y6GqeMpEeq7k0xUwpngXHOB97yyVRZUuR6EJK+oPmM7V/6szSNg0DglWfN
EOqt6jbjCQwEnK65zLFavQvHGOTTUDjjwR0iaAxdDAHsxfkIaY7QkBMTinvr
gt31xPDKRUEQFIEoojxyGcVPFF+gRahrOeZLu2pko3C542ox7p5vpQnbXESQ
0EC9ld1x0YLzgQFuKzslj9AY+NmMfAlhLHlsxNfuVepeowWkh1v58TgQwrno
+rfbrhfaakgSi3RZyF/kmRZH5PqvrjJ9JepeEGnHtsRI2ygWTOD1AtRyysnK
e3AOiMLZ8bubGmm+g1xgl0SfA6PmEYuMy0IB/uXcp04xe8at6jbooHPk3sNS
4qo6IV7uVTNEhRPcw38wzmurDXX6Rh+qWJGwOtBWio4PB2cK+H42o1N6cRB3
DmY1+k78dsXgff+QITQm6coHTdBoX9aVo8RTaMnLqq4u1vzSkpZOQ44lDi+2
zwe7dyFsIeyiTSmPe7PjYzWDWFyZlAr8w+AzCRlVKnlNgAHhXFnwr/s0PoV3
7UNikyg3aeewFTS1L759E/iNQUsXU/lGALEdH8ek5BPOxYxGLlwmbv96FiUx
kekxzoBIoAK6gB5CC/BvznnkmP8dZrQEux5CKjCguaddbZnRigI7qr2yz3gm
G05J7G1JtRbNraUQ3kCOthANIhiOQDGsKCVYzAAW8i9zLwcZGjDQOdPwJUPO
CXYEWud8CVF9D1vfniWyl6yGXQX5G0Msu96D6j1moVkIIOpfKMLLjXGKLzNT
wIVp9zmYnN5rP086+xA9L9w+ABc9ui+bvaq9YfBcatwXhdex3Xc2Q1EbqFmR
1da8SMT7bClLMk9BJh0DtoA6olRNRsCazJdMMe53bukZ5qKOuG7UrH6c7W2W
kBfpfG/q1juWcHhu3OBRHi8EjCoHPsBjxDrwKW5CDPHfc9569ZLPLGlhMat3
y4L5j29Hshr3qYQlW+Qc7fN9tkgf/EZRviUuNbGhFD64tgegqcptBAcuFOZ1
tSfDTWyCGulNPRKL39Ffh2i7ZaowOd1YAIdHyX+uwAJpecv3D/48LJmnE28h
wY1x9RClYtfa1K6hiKCDsHpjosPJtx8PibRHUQM8/DhbBFFS7C5a5fS5u9yd
rawvI9RByOxoIn73l3Z19VcjmAIlKe51KfBUo8q6BIvKVv6uE3mgbcQEcOPx
48bBm4pa7yTzHI78BrM8/Kn9JDuxLcw+bTjWCw7w3G9wHZHuhN+JyQsBNv/b
eCklYwAiE/Enn8wS+g58Bmq4yZX6ebSYjSvewsLPs3+SH04gCrb/s22fN7Ir
6XK8jmrXrZhaG1hb6123ILRsVc6iphk7trggUMkYdB+yzod+3b4QMDa2u1rz
DODUo72Jwp0MYYC7SSqeaduSZDjSGh1AXQbfob9Z9KJUvZgGOWglO8FRQREL
ueMOAWykReLFQ5G5FM5pLmHeeDKZe9E8CaBeN9TqMunBnGwJnVv643az4QtA
fUV5tKUjJhpGJqavWJTcDFz9zgAADtxntjw+YMyqLy1r1mfMRS58OtKZHBjM
ULLwPvT3Dk84QQyQ73pAZadxlxk/FrOAMMxYUHh8xXIk6gormesChMsVelha
1DnqbKqTkRqbXgGRW51dHRcTSALpNGYcFRwWfd4aFovZKe3+QmrTdvOclhy0
/7D9AO2bnTopaC/oMMNySeH5Zh3OW4tgfzIJRXlnARNt6K7v+l9MTr4GL5Zl
GiReho3rgU8WeRG2AdC9vqHh/FfWhMmf6Pleq7yMZ2NC+lwDL0UfijyTeCAE
0Y979Z3gqW97BKbdIVzkd7tn4UIsQwWseqoFCxxZCuD+TK7bHL//n5DF6clH
DhRArDqSKvHaffkA7nWlrro5gfiumkrwuLlXMAxb+XPxcazDY8H5XdnR6f7q
prAgcN3czISW8z2vyOqigjMbfmI2e/mroKKgfRBAArLLxb6wMFlBjL9/WRKI
q2X23K41sVImWt0hQ6tj6VTWz3fJ9mI/Ev3yHlLRA/mo5NgcAw3UCyW/PiY4
8vt+mxxhIMPlQPEjsAp/zohVcASQkGvIE4mkEZqKYF/AoTf4N4zui0qd6sLW
KgqHY2eO/ov/DH2jY1yrI+B/TJbqYpQzH+3x0u94QcbkX+gFxQoRtyyEWrl9
iPnVRo5GywaNLz62mFebFWq+64LJJ7p0ONpYMUMVMFacZZN6eZoQ+BbZouPB
fEgbzlHwh185OuVR6+4JIMNaZUD5kDgITVFeg58goKsnwM1mmVN5Fg2b4trc
vXrDH2fSsNLGEcWRjjTBtvtpVwCybN9p9J3sPULa9pjVn6U0GXJGrTI6AADK
j/xsp63D/PtJ6q/EEo74EoHv2h0CgXmEc4XlKgswpp/3WNH+F8E+bPcBMuL+
yyU1Jss3ccBEGwXaLgpMooOBlyDFA+vQq31oZL115fnkyWT3guwbFZLb7Kd0
y/4/DAOCkoS6eI5wv0u18mt2zBH3SMVpSyT6pVdvK/TPb9LUBwI1pXFTIg57
jgrPZRFfMWFVAeGna7AFpSZhAKdN3HlUlItlir7A8eJgqjvGdFCW+vbVxiRX
D4j4EFvzn0glG9d814RnY9xaYYmVN40/gV1JhzDMLKMT2r2y+4j07VV9+fnl
/cpWZv0M/jGg5FK0/+ZhcsOLb0LWbTeI0P17xFv97PAwwIUm7OL/X7VvfDnI
XTrpwWJYidMUG1zlfzU0eXelog2TAMlt6dUAKIoPsuQxZc1d0yogT5DC88kD
hQ9G0qpsalp4fNxniDZJo1slyOOQWe0xy8lG8k/67T68aB6uqjZBJRLTMWkM
4gtanQZOYnu0rReK8SsJb+0QwaqkY11banoYtVAoHY0cqeJdRl4vfo6P8vuB
twLi74RvFY1GS4mU+huCplmcveg49cqLhGD5GbQ8LOIC7BS1UmHndx5LoALK
Ynj8R936g22FjlO5NSpQSLTn7e4eaYfCALhHhqpj66+4oCLKe98im7xjOBm1
8lx57T5OkMW9IA3nOcTSCFiRxmugkA9hM1fraLTr9Wrtn/nYRiaPXoIoDAdG
Yp0zPLEHULBncc5TfI57ABteGedBWiDAYWAyL7Hg+jjFpX1sN3iiOFuuxXU4
hpweTxEaMDiAjDOVNBhTnk74PjElbSUrGXxMW/BIrV4E6Xi7+LJ+DqwvbPTP
oFk4pRWE6ok+4dTqGMrAsHN4ZkwynUKed3n0vqlYY3VDbQX2x+ozhDj2J8JL
7Q6pJ4B+dGlA4pQdjbHUD4HamFoXJJEgRV2KkxL3DjIZDbDP6dXs8cNGg2o2
IzXSMlOo/dxuOAo5GcmQfc0465hqJuthNrBGUnzYVAKVB6TtnpKMJ4P1KCxK
Dot6HAqe7qKDb5ZHgzBFEAT2A8tQhjgBJa3CQczhPKQa0px9isWIF112NSrr
vmlW8Z7DRhSOt/Tb6q29rAvqIv0W9qw+1SLtvG/vA72aUf48eh1NdfdRt1zE
7gOuGuqz2zZycOHTFJ7AJk7PyyKAtQqGRUvZwrP24rBTUkF6pLTgXcKPMIRX
yc+DSZA56tjvTc+PX23K25shzd4Rkg7IrziZHmUNaMANwwTCHRd7c8YwmCnJ
724xdIzEwJDEFIb0+EE/vHb+eYjqDUd1T0GjA2RfiZeNCc/QJbVGAwGdXs7/
KrzRBMbSHxeXOqZSCRerWMAOrTlvQ+tFMyPpIH/Hz7E8S3b/q9WG/mTDgnSP
9n+dD8JbxiRNvIS3iiw9hrRaSw7H+k81Gq9OFlMCLU1YJzwHFEEgdvGsERgQ
qnfReAYmKoWF6Yt3KiN5zBvTyupVe9mna4/ISDriIAm2ofkubqsiZf7osAyA
v3HRvzCJ61d4ruWNff2+Alvga3TPVYIVS1MGj/goDJsL4I27Yx7Ei5MsHIfc
601hIubh3Y6cg8CQSTre8LiNvlKlQ71HVLwYb00cZrxjFb2h1qQ5DyRSTr0v
ueKQk4lELUHldbSoUNuMpib/HHfBeO7C/tN6NFNYjH9ohX+rjGnpi/0LyXFs
CUp88wDZ2ig5t2f2fmHHcTtSJn9IydmmcC0eL0fi66C6pZIlI3JAfuanfyB6
3NkGg/UpbrvIQlBkBPWE1+2op7lffa4G1bRD4EkmcPUsgU1jNXVbTQ4OBzpI
HkHYxhK7bUozbyiTVfQkSl5riHdlwnFngv+9kYZFMJpXVCrIoRf+FdQ0sDJE
C+ARBFWBMvmAlsY7QJwvlBwfh+0/mTTPOEwNGuMd3if2wRvK04qCt7/MmKT0
I3dm5MIEozQZ1GwOd0j7ZHXW9KLO5hJa8nRV2cwAd68h80rMw9SXry4bn/Me
rz7swpfrMTP8Vrf8WrXxDJ9E+aMI5Y0ma5FurNZp6fKPawPGwVRn/Fa9WZrC
0fM6NdrdnyCy+n3xTkmUhRYqIj3FURgoeiN0l1OdqBjed3ajIXCELWG0X3V9
LDc0SVPnHJ0XDooVq+sUXbYQnQ3rh0EooPKDRcCXnDu/HDY7xNoTOZeCofrr
b9NvsucvGjpfIrPHNS5dyuBUVRBduy2pFrZUGc1MJ+YMfmFmPH0FLjcyxjxz
zEih7YvJAxC9ovX8lWnaRZMFy+OG85hoq6s5ry8CwdMLvwGHThbiHyhk01lT
N6SPInJEWDX7S/O2ChaFNJR5Ad3c32ImH7d4+rToKjZQhMhrFaSHgfMnNBdt
0RldppwMMMABcWbGQY/xCsZhwwpGFykFrDLMS3aWmG/LkQLv7V4KQ6OApA9o
oVnKtWpr72iQqaSbrpSSvr2CY4LFwxHJYONHBKkEY8tyaENNdvVksclzk7NS
bC8MDnBoPuYLIVrRFZN97mNMKJfV1LFkYMLn8I2eYTCEjMZsELa8k7oxqpP5
Il/0IvmmHr5/Ra5w8AwjmtiqN5wmowI2UYDbAE9spWWrz6bEd/yWxa6v5hG8
NGFIXlUKbSRieWoxplW/P72oqGrroXPL/QetNvl1Y0DUW6bXzQs9maIOgYpj
ZhRb91wmkg85nmlOscD3K7VqpQDZktq5jktVtCpZ4PZBYxygKAK5P//gwTAz
kiJIH/I1prG/6gxIScoJJgbD3iM8m94tiY1yxAHJmF0UdaI5NM9CzPwnEWko
RMbsOVLsAqPZjPGc5lbLVqx/oxGxeErr071Jia7T/y1MOUNY5xrZMdo/wROG
tCPfVBAy5ajd4tGZ7GxxTMHO2kz7lD9yIJaQU+U+q8/o6IOkTO7PiL1TP1kh
Yd4c0sIvInOg7QdW3sDztF+4eWVSHkMEuHD/Ef593qyUKWitOpMipFBp5Q+8
b9w2HAGddpxOwewRtt7WBhRB2njG2ku3SnuyQwi//jWFwlSD4Q02fZLg7dTg
V3EVtXAIaICCP2iaf8WBVKfyDBtoyKvcJIT+iVCKqfvZ31tsmtagQaMapNX2
MFsQ+KRjh8Ozff9w1bfSxdbnCuFOWgcwGgJxBGJboyKO//R2wlP/d55zUhmo
H5hy2a2lL8Jyw80dkmxD+UxZrj1wlKOVeS93q1Gaz8vQdd3Zy6ZOJFqNHe5g
VPwoUuSrdjwkpzfHH31xhY/hAEZASO+oZY13Mjx/9HVd/jKEo0PmIMu16G8a
vpi4M+l8SRjQO5rjczZQ5RGz/oymPKjdmUWSrG0Ifsuns4avkiE3LbfQBoMz
weoVySZNgfjM2ur45jBTgyXMoVH3M5pfTL4xsp/sEFxhjNWYCo7fjPxoR3vl
hA6lQb3bhjT9JjRL2xMylBPV5Yjxe25wb5Kivu71/ybOFCrin/zRRximrxJp
5vtZrkhgsWUr+oIUTS2UGTkfQhN3DRxJh6WAh1NYPWr1CGKgNsH6V04Fi5wy
MTJdUF0Q5tMFn2jS/Tmc04dr49sb7My7GxS+6blCrvoINsmdyM+xeIxxVnBv
pi1gwY44THmzRVYFiKGdZ43AWSNd1ULmivO/gjeDn48PDB2fyMZ0EiEO13Rs
dfYnso2C0zgLPLkxX9Jm8+lbHRUbhGxkDXxEYteesklUqZoNFjeeq0ZLeC/W
hSFmu5vIeqDD59P8pd/jBnYrZN1jqMDEyHWpPiNodsHW8NPHBCbEd2mehsrg
rt3TxYrgOcrzJho64apue3kfSjuJEELC6ViVLibGyxfqCtO2HPsNF8RR2RRm
TFABHdzEREVirVBa8La8rkZlkYB4jmUQVM9FZw1sg3nuctKnUrLTY8dS9Xof
6H/FSTECL7UsIbfrNwQM64sosjLNPc9xPN6CkAkD1FwjJ/8eUu4fHqusqp6s
+BicIwAlaaWnbU9Vij1sznql395ylRcHr4eYdaU7nohpWbXEFoVr7/DtGeiH
iD16gxgwPQvc3ztRb60wgqwhrypxh1SSt3T7aeVbqf/4bALAhjO4wckpOV6j
1lCwImnD8TsHvLg7+LOh0enfAE1uNRVexoR9aVE9PPXCiApd2tpgEkLMRXbM
ZB8BYr7GpJXR4HhdeaygmqmW9+TjpYY4nVQ2+hQW6ftYPfj2SHafeG1qTf03
Qurj1UblbaQajz+aBlVqVTir8QMMzbXmd/9CdB8QNFPFmtLF82QYdlF1l1u1
C9lnf6Db8agPrNW3Xi6iWnAvcYSfD59oWqLSrkPQFju3vYxz02rNBrhs+WbN
nDIzzhZvs6Ef2IGdxkvmqy9J0jhxTK3Rh5WD8WSfuel/6bcRnJXFFR2tfJ5J
2j9srz+jXPQ5TBglrHD4GbBocCDlPvZAioW0EL/4nF/lJjzPyd8qnjmHBMQ6
I5GSYcR/6XhDfWzwtx676BmWhLnmJlUYj2jsvxlTBLiEuFjQOtpMoUEM3F76
CZx5oGxdDm9+6p/7WqH+ocBelXFJqPMO4Oi9vVQI/hFu59qAlONtjOrTTacE
job8XdoK3qI6e7ddnfW1d/HuL+6iVmKFNMu7aWbvQOXbj6UrKemJ2dZhYO6Q
O6tJiczSetKBC326bvgBZuYVrC6fLgtTQdX9PbPfUNl4Q2b24SwxMBthlSRR
fbTcyPOoII+stTBRwB+N9bF/M54n9QjQk0JbX2au+g2kde0UAjAANOR79WSs
LiLdpok7YUD8PZtzoKEcbvoUYbYp4MpyfjKle44hk7VybS6Zk6Vn5rQu0vZd
TvTHDOnjNjPdXQlYNugvC1aiSZBL4AP9qU+ats40QOOWpPIRhHPToszofwmU
/bZ3oxjMVaiXAWSxS/NLzPfT/ZYeKmDE7vYf+24en71tG44y0EOntzuBTiBf
y4YSwOFDQNKeAHUGEmqDNW+Ku+ZK93iQGERDE+wUA3GFsNWvTtobHLWQHDGh
SEMJofKY5IaPVFYcUHBd5WBQNCRPDbjw056BWjk4225G/KwKjQiiAbtTam4I
Wvp7j1lMl7ZzRVsJVE8cei5gdRA+sH2r+3ebx5+yvS8EyYaTzk3v/G2TUHPf
zHV88aAfWRplYDYtU1dyYz7CDVcqIZb8JlVGUOE+FRmLd+Yx6uBAzhMY1jCP
Lx7GH9aSTIRLGoMfhcnWWIdcs1KxYU5qTVsNdpwKNavWgclnL2rPhMjtgYtN
6FGyfU5QTwvsmuw2PlCR1GPLtL3jPZfBCY5tL+gykOe5bDAqTyma+ctbLuYW
Jd+D+9fgI/GnzeNfsZlfSD67gM0ovEfT1+MvrSMOIovizT197LRmhc0wHlQP
JPUPpXbOnjkWIRAvfKGgwA2XO+pLUwsEwEZgAknDCsTY2KcTuvCiHk5ui4IC
h2R0mAgGKNcpJQLBevPzFj6v4irpL/jNGooSNSPCtVAFuKHMHInmnZBw3E5E
o6NPcN+P2uVLzeYrLTw5HScg9ZYTKewlK4gBe0Z9Wf8tXcxEy/YtzfPEjkf7
j+7SwxC5GrAEFulQvu8MmSmBopLhG/bTxCuUjottSMcXwCF664Tnccm86bZR
l3tkYJd4rv6DeiM9uAfPW+stbWhUv7CYNBDDCglMNog4Tlqfo+ogSKIPlF6B
xk9CV1K1pOLM3eXG8BA9Be8OQQbl453c1SRAeNQhLmoj1VDq2i0q5F8AEYVT
zF0LpqS0yBmpEbpRdITZXPW3JrMsF18Xs9NLZeFJG4eOsM1iroviWlBS3ZV2
eByWew8eaFXtz1AInCHvuLwJY8zbwOxry1A1ISKRFPQ+MOl4KtwY35sXcsbk
w/P7woRZlKrzLzPSvREbEksBiS+2FVqbB4GEXV8hHsdXZqBNTAwKKDhr+FDh
lTkoG34bGqQqmmlSfDcqCQre9vlTdRUstt8o8M8haxhMuNvlZhmqEPyGy3VW
Ig2rbni3oI7PjaLylES7T4J82Dd4xLYfUJDM2JVEKYZTfozLX1NXqxTeuo5i
zGdqXz+bsQORq90CrisOLksnY/VSIxb2RQoSA3+BNVY23JaKnwQI1n4zrkg7
p3pDael2mL/6u8iYVUMFnENYiZDFv6bXugcs6fr6NhsRc+bXD4W+0gD7eDV5
8+DWf43X8B/k1RPdupB0h2oY8KmG8pctG2LHqzX5MkEo08tIj9CVOL2Ym++6
4aEypCWL/MIv1CCGuMW9DSRakovW9zDpUtaLGNndJY8vWHWXh3is9wCNhgZ4
WZn1P0XpBdqgkFGbX78tSa0p4mWquRwq30ryVTksiGyoSVJDEgXH3rBug9/M
K2DAljEruTFGx8UtFVTGzqmFlZoStltHjXVsRZFIEiILFpqcQKEn4evVR0tZ
ZoiTfYKySluQiEhFauXKZX0hcyStOcdDDE5Bls3uZagFRAPNuzfIBo44u/UF
+sl2F0Tquea/m7wvGYjU6wkyocTKDfmKFkAO1CiiWrLZ2PFO7vgD0Y0i+r6z
zRbi+cb+BhDtqUlu7GjMDFFFSljkENVJ4i4IFw9YES69FawxLphUDvgZJRtu
Cpd52hZqbY3zFVeOZpTqu01YDG/ZFyVmSGmiVr6mO2qa+nMesMBcw14MQkkg
3GtxVB/08OWQs8aiG7dAiLN8gPZrrPKprDJj/ucjBAPPAquCYOcF2+kK6GYs
10RXv9mxRLQFg5EceVWAKvhHAk3b/sVaRLx7CfzwSrI8NRXF7zQZ/Lb1XbRK
3KKVhOcwi5f45jV50RWeeRsbXIKtqI/VE3TH65FigQv2IM0p1LRiGfzMGFjX
dguIDYY38hFTiHJG8s+QOJoN7yidAO0qCaI1ZJNJa9aG7Ni1Ls0jVoe0EQ8V
p+WHHmf0eystgEBFONGn231fzIt3uSeFrx5Sa+VutJFc7WTN9PwzfcioaG1z
gJ/7aUUTl4XvkMx2LEVTOudkzS05XFjwL5QDgDofxITHIZwY33ystd1hAWD2
IWI9mnK3E8TTIhLrUX2TK2Ss5G3xeFDxkeJTTPmEcGoQqG4qnRH/Z0r1yQj+
Iujtno2dA3OKYxjbAKQndSg+BkcluMoPv8sGOZ5ukw3rzxRyJmEWAXntxep1
jx2S18Qe4Cr9s/OursUEQZ6wKx3t8o+efoFE3mo5qZR/8MIkWxOqWPtIYaj5
59aOJfk4P1+9hfWBj/fu3iom0IwHYhLkrVGK5DXBP42ycfyffEYEhUzpEFZt
jY7zDwFTgWnn7cF29kk3n8d00teKVTFTyDv21L9O9RohlXAeXLhfNeUzsnBe
Kl4I10ua/hsmkvGiYfDirUIgRcJvKmsZIiUITl54LUoMAyq+y3uM3TiGlK25
kP/o91qUEeNaLNBPAFM1rA88cLy28Uf3UVeDskSr8jXG+WkWS2KfqEMLm75S
CzU8WWj1Coc2VwNKNRCLNna+uXyASbcq8bqGEXXMQUr+xQlb/tV41VsF5Qsi
TDfZ01bda/RZ3+7h1aeu+zMp1gP0h11Dv6UUt1AShmyxTY6l2bi6KV8Fxi38
vVLjSaSNQRVAL32VkgR7bYRsUEhFIDsAtk7XnWnEA35MgTNKNYYBOjht1nvP
dnEJ4Sb9bmR/Rh8lqSaC1qGc6wZG3rwoaVaK/CEyWJjccpmmq/iw9cA52fTV
v7c3DsuQhrYgwIPC+l1Y9YbCHGqslg/xXsAEYP2/GR9ynZgPlzCn/mIPQIme
GX1O+s48tsPUgfhqL2nN3Uvg3dm9C0Z4iu0IWxE1lvv0tsveFYYN3s3mIWwy
4NpuXUui/Z5pyEKFSRsYH1OV2R8bGsH08T3A9vMFzq7vUCxnHEX4AVFkp+Y7
NaJ3HEg/Zi05HiLv2XCxBAQYOsgpwoodsaYarb3NpzkwE8+JR/t+AufRukVz
iDJ/xsF1CG95YR4HxPbPaNd9aAULeEq4Va4vohg3wTeEiwRuv/zZoOJr04j7
/w702pd3vGK7taEaFIJ3oQA8sdD0YQ4IZcBx5NSgVCOUQi4aPR1rR25yAhvr
lzSm7zAcyPB21MYusCebzJ6FcltEB2fGAnAN2/sw4dJRm9ZNKXDOruGYq1bD
pNKhDojrOGl2zau2E/GwADU6ybbV6i2wLx57UmiV4fEq/NY/rAdoB+dPxesU
1HtOX1WUFSHT+HnLISSC0vKZUslBIAtBrXPgDuK1+XnugfRY32a96D9kybE1
u0CIHS87mPUL1r48/YkfSpHg/49h0Y7F7N0kAbiSJnrAp/duw18oSzTO7b+T
j09vW7f8N/2jMPLqddVJ6Hg48TqUHBW1FpuzSB6PlK2+b5dRbHxRuQY1zUt/
4Eaq7iB4WUe3RilGIj8gPIKEGArS2bxNbnkMoOCfv999I3UvTkuc7lDgBwBv
28oCMvsraEkuODAxG+vij//JREUaCcFwy9zUc7RZ3MAtUNYIzetA6vaA8qAc
Hr4PjzaE/Ulz0IumRCkwQ6F8dpluuK/DYHkEDfF4upHst714tBfVHpLlnzVW
nsu0GzrXLB8wumT6U51bidGvrx0TxL50eftzKW3TY5Ps5eTqExexzooQjiRp
pOWsGmdN4qyL7WL2xVezjgUCC+Z/2Lebi1jpplWQec5W7y/SQDJEE6v2z5Lc
cSsP7aZuzGZPlpDXhmUpjlUlJOJ+4mUMkY+oqoYtUJud9FWDu8UHft0BrGdG
hMFThrvu6OnVfQKzwzHizy+F+OFzp0OQU5UsvtW4Tjmj66/LW9gz4nXt9Lc3
6Ve6cMPNu6K+gHrlqgM/eP3xC3S2NaAg2Gy5ElJjVVBYFC34MIqqj7wGVuY4
Y9NmhwCbiDGTzjIVVuVTTlVEIAssCZfzCey6Odfm/L/7F871idQTxHvle/+v
Rxh9l1R0jBH77mHHJOjIRKADrjda3oVXlX599lCLqPXbdSZpvohn9gqc/MFG
VU2pUSO6ptfeFWg2wjMrrb5x6hQgXTY1jDjVa2EYObYiueoLL2TYsaNaLVCj
b7drbvbvqv7gd9R/MjBpzE1SzSgoxPab4nJvVfG1QAY/JVbvyIUYABPdkgVy
rfb/bHUUnkq0SBx0Reo2axXF7TKhGTsIH1idCUnVGFV0nnW3gJ4IF9pPbV50
xio+4Thrh8LAnbMLYOWnj/bsWJHNzvsrOPxNWz5pmMnUhplNtHBGvvC1F7rt
yrjHBgTNtv0lkR0sQzGAqEdYL2+vjgE7HfAMllL0D5QxFpdhUPLqrAxcieGT
JiUk5pVxA5C9oZdHLyyInuQ+ItNIQhyDwLIKG43yJpm4uray9gzkL+kgW1Lz
WwSqmu3ZWkJdtpKLDObnImEAaJsxbZ9DvEJwEEdl4ycmnLJLd6zXhlQZcCyq
KkpweJIeCosxX2LvfDvRV7GQ7OR2vhhK9KH0vroX0mlC5PTjWGlsL1ZJtXFE
6Ar9qJvSQNrmo4x5mIYmHYBusYRQnPkMsSdZEXbJIcc1VNo25+YUX9ggcA41
5pMrLikBC632l5yBI0pHTtzp+sXPA33sn8cftK/lRnMunWHCmyoytOElvbH3
0/W5G49H+gR/nHK9U5K2QtYiESC9TZfkuQ4Is9zPNWMq9WPK5YNAaXLMWWNL
dMwTanrbnJiZGFyC4z2LRxmMVfeiLh9ZBhGNz1QBf3bVC9/2NRzBsPGIKtqy
XevS7HhsOw2SWvByPznKA5Wy55x45CxxZwnTqe+YdLZzhjnmX7Sjcrmgmx92
UVWnhcYhKDbyZOdSG7xN8G2DAZiYhCP7t66VvwjpI3bS8luhIijA1fDmamNg
VzNwuri9L/ByLkXDO/+1Bj+xaE5W0cJu3xoo7MOLJFT4ZfZMQ/p5iU7Tt5g5
UAzG10kc95wk64ns8q8IwLrwpIlCg/gJ+yYk5LEyndat4V/Ai/m+AL/CWUKA
fcJ3Ul3QIrJqi53XB6MmJAznq5dhk3HiYt1M+eit9vB05woex9DWC3h+tnKW
KrsC0LJJo+xe27eJUX6cYSJsFi2vJACvxOraGoeQGWofaazfXT6cezps+TZI
2jVqHG7eapDt7+9GpZvbliGrEAafp3MZdbOFnnxgQuMA6B/6iDh+uCjNiYxc
1j+RdPBP0ECWpXrOSg14dFHbpl5HCJR2koWIP6Cd3xFIKElhGM3AqaHiCcYO
+NEwQQqH6oppWgw1rJGCmhwNUixnSYEjiO8d/PWF0S2dGSQ1+BcO/x5Okcug
YrL36SQaXMdIYu/FoijATRycK37iqeqmtRKzUBHBvTYTG5Da0YthwtDMX5AY
dgcGcxYK+F8pArLDOVC8kt7BodAkpXj6VTbu9iVGjrm5ibWjd48U9HAfDoYD
DTufzLF4uuu/jSexbat7C7CweSr0UryZ7Eja3pmOVLej6L+uphYc739bVg5a
9NGKUBUiuWTvUWMHV2zQN3ERCpO2EWq77TBaHebMWP/KgIbo8B3Ro3SWnbpg
3jb1/qgVVGKr4hCxtwalEFOY2/KVh9j0KFNPuyIu7E7jUhxnreBFxyHc6R3L
Z9jESk1UOR2h3mppixHaAmfOHlx4cBgUd0CeMHxHrtXR/Fr2CWvyh0roFGr3
F39LNDiqOaM9fpmicmBVAXrNRDn4554WcPiPrHnFr4gXPBFUv0pDj8d9juH1
dpqIp4C34OxUw40Fk0Ca3+ud+3JiL9TEMmm0nRGXkI7b5rngOGgnFCrqLyf8
dTct8nMfs5nPgFxbOb8B459FI9T/18CfaF/T5EHhALTvMfjHxEJqyxCud6WH
zvpPlEDwzVGIZfxSbRjlrTIq5Ygv6Rn+73bcbPbIDtDE/MG9k9rgKKJsmpQu
0EQg2nWiQCLQMGcWt4tLGF4qInBSzOU2ZksUeG33IV/9bLvOlMQ/xB5HmJ6t
fe7789JTDfe8Or29PH0CcuOch4bpppMIE/u68U9rbdosFfK+C/5uJFnwDsXr
Xu5BXc1N3XlEBDEy0KGMEq3Ivo+BcpMQXSCOi4lj7qk2sGZVrBj4+YQ67lL/
+EcelqEZoQP98WWSgEMGH0LiOiUSFZg5E4hV1bnKLlDRwrF+PDfpdMAP/gn8
GQrDTYNqeA62eeoHE0CocgxtuB0bdEG0/seua25Sk0cw+HQfOroD26rh83TH
N0sX/WoFEbDagJZEb1m7g/vsaSVFgprL92kDZsP+gezoCJXjd38b3Kp1S1CQ
ibRypp2mS4Ne0DfFADTnh8cv+0GFByXhh/2CJeUdK2u8lM6ZM3nY8kE+BBhG
2gfADK0X4xakOSqk2QZm7LQB8jcY2uG3WnbbCOoyQgr7nbxbZ1DeBpITVN20
vlycO5Vv6WsyjWWj6ooRiZbuoVv4LjwcUZwUGxmiN8jLrBbJQY6OT1B2k1ym
PTicJy6LLIi7EQqFP8yJpe+2tzDcbQyJhASN4GHniosN2f8RcQ5ZX64Yl1Tx
QhqxGMnRlxQI1sgo7TotUbutIHwd6oipiABWk+wW0lqBBYR04OkHfEt0UIrs
T6CtkEMpBJ1qYUoziU8eaIl2SL3DOGNP/jNJS52cmTp02FgiXCBcMemmK0H2
4GXL5TrwQ5drofTkOsnH4jefcy+mzr58wLaMMte8uCOBDTwR4z02zgTe+T54
HyN+Qi/sQqiEuuMv0Qymgi2NMBLUjuX+zCXv/wFaVzEH88rtV0p/LbFwr2/q
UbqcXRWF+mi4Gap3GloMpvKgplBgRsUaP4IvzvoZN8oAiCae0NGECmzKKbv1
xRV/OHWUqlxyO171qTw/fqtQKN8PZs/LAO/rEyrmspFy1cW8HFMf8OZtep0J
adOl1VXHofuRqsBe6uMgwvJBmjJ/jbF8F0t1op8KEZDiuU9T6y6zNezGtyLp
NfYL2hr8pem33+S6f56133cKM0UmuQ9YGUmTI61XhwW2yOtXOJy6nqNR0HGQ
UyfLiwo6NaC9dPR5zrlcUiJ9O4SPWY8QJkifWxXVvExI3OJjpvG5/77fre9j
p7mpi7kQXmMlQnjsK2NRatKhkapksrOg7P+99GetnyniJgBfqyVF8QGmETrX
dBdJlRT23pF2Vcr1eE1Gxt6ikG19smc3jgkJIdEXBCxz1Q99K8gLcjiY7jt2
o6v9cymg9kKGoQ6Qo6tJCmke3FKGKFya2jrN/6QhusBSChBc4XgP3UdNvmd0
OIqhOdKe2ak045Ob/COoVOcy6v1xeo/oJhZly8oYf/LjnLgbachmUs9LJyhw
tl1Dfo8M+jR0pm8DW1cH+WckWijxcKLd2OXc0baYNc0aJoq5A5NyOzQU1Awd
g0kFXx+HhqWiBZQ9tc1I8anZk51ueFu437kAi/rM1UJYO/6diyZp2KUg4l0v
UeAmped1kbchN3smUL1mOu57cfNaSvVmt5dK/D0jHytqr7C3Ld2pYPfE9ZvW
mrJVZhUo18WSRbSgFa6HGjsQ0aU2+/LzIgyUjY69vpC+kVJGx8IQN9DSp4JM
Y+6mGPoYGvyjPPzk39BWSbmX4IjX9O42iXsLAhQ+AouxSNtNdlB5ansXdawc
ChJJT9s7KNAAdpvV8OHDpMXW/sD10wFqunkfBxR/mOgrh/UarBOh9dPMirq+
FIrEpPqZFnv3TclC57DO/CJsniTTPqIys1LY6Nc0doRHmjYfD6RkbKmhUIEG
tfcVKrQI6Yo4xn2tSPAt/ZT1preImv3GtdgEChrwy4yropMX5s+1Mn05vCZ1
xtoiEiFFOoaW+/k56PGqESc78uCTV2qk4g2iDDfMGAIrjR1llozR5YL3Dj7u
NASTcDKuq4oFhLL+7pWOTRdLgFWNkA7kE2SOO/Bub+vFKfiZs76YFuwJcS+F
8ulfBxsxj+XS0nRhEeM4AVLemYuoE+ciRg8FwYHeY+q9yuqZ8K3/RCg09Gjn
cCTPYVokJA10DnGQ2XcKpg9CrhRQT1YUG75EI8Z3DEzceBcvIVVLd1ud4S17
SB7qajSX8kP8fxb8ePcVxmVfTuimTodLYHpH3kqxcBywZnQ9muNdGK7OFDJa
nqCPB+XpaoYsJzCV6kOtTfWdYLtmZ2BOtBoPwSYs3Kj4MgN68/4lPK+49mlJ
4dU+9zNDIfvSzBD9UIccEFnVwsmB61kpQjWZ5pBfeI9yA/sZD+OQHPGzpBI2
rfq6swkX93yis7P4wYuobQzNlLBPrFO6frxPQa1Q+i0eTrrKvaAWG3jg/rjZ
kyMYtlNW/R9W2qSTMfi/FyMCgoTQnDm9mSOokGIz3b9GQavjpUVdxs7/qvzc
bXfelDth1NYq7IBjspK8vUB8wAkagVI6MIRLkNqRUgEEcd3z33/jbSV1vxuz
diaQgtrmlK+SBVuFiuBwIbfwO/+gvlt8L4mo7WWdtfyKm4eNBFF8LxTElHX/
s9y9BboalfCRaa/egWCZhR/Mcn/VPBbLvz2PCtkNCWknT3XJ+Xxg3D/vvCND
4PgATZ+niitGr4X4Ig6Nd7Js+rZWKgj4QTqSfYOeJbt0w+YsZobdfW9jjGf2
HIakXnX7e1tff6xhAxnfr7OvEjD9KBSocDv58vy3ru3QutPE1FJXPUFSFQa6
9JIJj9TY9mBIhbp6+WEsmgw/vBHlt6Ppaz5KKafub8n7Z33Gozj5mMSUp/+v
py6wwvd423T+qcm8bTmAEzAjUiE4MVm3WKRaYVJ6LRsTHZdoVOrGIAgrfYP1
FueBfb636FxzDmj0yl5xPbog6QOQVJ4AaAmAwlVNBXvmpsz9SloiLrhvvats
7YnoS5ZttDSXTiU/iMxdh/wT3whmCXD/1pd0RFnxnQxddx5V19UsXFXuhVHt
IB17dM6vFvcxMNuyLRg23GbTrtJ8HeKBz63mptSV79oSSaZogzlcmcj0Vbu1
DYryscf/r4jam/+woVvF2eGkJ8HvZSZPpQoPzPXRpb0cOOCFvXLmTS3ZxMD2
7S8KWd7qZXpKdiBVmVYM8OyovTskBk7pnJ/SP/zCkx8N05oaOYIRMA5V3iR9
Z4DtdGlLg+1QH3hXG5S6sogkyRV/Vt8w7hqsSTnjJCg3H6PHd3OtQ0XCmlxG
t7xH0nXY9VrbsJXP/OA8Jox64K06jzyxYt6czZhcl4j9p3wQm0d+Ymmutqgx
5sSqjc4v4oxYVmMjelx3P2WPZCUMtQwmZBKmPI3uj2UyG8+MwB3WLf/TXnRY
cKov1UvOYK2ltrGzyVy9MvFrM9H7npkIkjjQZa4dxDEjXz0blMU4E0z+/pP2
a45Mjf8wCimzVYEfcADz+Mr+vd+nS/5Gci1Gfjw+ZEB3d6WRIrByWctI7Bst
N1s+2r8dpn67bAmpojIXjMTSCI3SI055Zp7dFRezKvFEtm14kMr30iEre3G5
2reXHa72IaQJjGfk1U0VbJYINhMrQ1n0UMhYR3CiFdsnHG90G+R+oSwfXbyt
1oMw2iiVN5lo8XCGCWYBlpA+TDyMrkrB+AwL+bnS/AdDw9IpCotgMAjCzg6N
c9dgBcg/culpFIoTwoC08cy/BIcxC05XMdLm3x4Y4ax7v8CL4axeqsp1FPMf
hAz+o6NSvSub+pW8QFcigf6PQvqsUWfTRJqIbqmlR5cniZnn3v04hVrF5+ct
UN3Z6TfNtOCmMMBJG+pneedmXHEQuGzEa86DSBYMogoobgl/AqDYD0gKJjuX
cMj3SZpEWpZafRJ9ZvFSiXMoiuGftgb2zWgvQlt/zqDUzoSpo4ioOzQyGCmM
8fBTcR/kNzaCm4OsWBGe4yiIMas1cwshM+le13m/QknaNlvDHjlu+etra4Kq
oqTbBYTgTjd46VILSEFxqNybMlj9kINpZeCrRocO/1iianvidYi8Crnd1XD7
GQ0bO7NNkFPypluDcgIMUldAwRodMsDxgLAdc0a6p+DADQf5z/7a18atc7Ga
VNMSOfiyF8oYgSMKmHchz/qZwuUEko06klADBR5c3sbZvMaey95kbwLmHDKs
6gw5NqnRHuexseb4mEbRjI0Z8IxSncjGb+8pLA+mJ9kmeIExcHG1Y1HGBtGN
lBWH3767rtz+m5E7MahpXxR6jmr4LodNN2oOMYc3UTsD1koban1PEDCDTP/A
BoPqEYhov99yG12KJX+OL9niU3QxHjBCy7LGTLsREIgGSxHpvXyTX6EB+Ofl
QyhnrigGlGlTI4U5uEG/k5ZPb9wCO9ZuYcqvtpZB5FTnFvEX9HZjDeFznu6+
U6CUJoO79i2ydm/PFvnsHmvU0DryAixMSzSXKXp7JFV+aeMFuTNfoOj+s4ut
t7CG91zbBF+4v4fN0HnHiuwqYqqeUvsEd/sdmoqRGiLmksI7CxtqHWeN3Lx2
pYXwnTTBMX8pBKsn4g95QvHLv18agUCNwmi9h5Xk9h/RnLht2Hl6183uDJ0J
A8P/7Yw0wlsrOM+ZVDq2eeKpqbMQhLRkxpIyeAQXR1Emu1S++fkRw155lBfS
L4UeXGkqOKVqhskB8gDAREXZVP2KuthHMwnXdNslauEM1u4j8pmAUZF6lSpU
E3fKgY1a+BMkecZeSyagLOoWYZ+xVWgo+RrDNBpHq6xcvF9bI8E6mSKMeZ1t
imT5Qmwlu4FDaH6Nwxj+ENRKZo6502BC3z1ExkjFXHc4YHSY6MzzVljd+gOn
XTPqGgIREpogKOPvyjukG23zLAIkus/7LABd5hcCiaFby79lEDPFLoOUvUj+
C5e2vN3JPeYRs5nFJ2PoS9hzBW0IFCQ4ssEBYQGLrknxe86Ht52Uh1jeCwsv
kvTrRu1BBD4x4+aE6kCQKN7Q5U5SHJHhF0rKCU6LSXAZh6jOX0UZ5EYv/o+I
it2CFWESAEP0kL3Yy+L7f7G+S43TpranQx3p4+p+Cq0L45SlcYHICm0CAiHO
+7iihNEHO/rzy1gl2KSuF7yrLJnK1hKW6JaEksfUwk7f0G9ifi43Q7cOdPeN
19nFL25ztCN8H4AqnGqiEz+3Bn882/coLFdrjhzTKFlvddtWokocqJ22CQsq
81Kb6wKaHtIIp/iePjWg27NUrl5eTDFeKKkxcV2nl3ouj/gUQgPjVdhfHwJH
Y6XzDYtTMhpPHzCbr3g2VR4CgZd1wswqrMX3j/EFLHdMU0UWdLP01Iy2/a18
/+OfX5QGbx3T4HqFkzi8i9jARCb4F40hrd3uxvK3z7m/w7sn7MFAFfLdlFrU
9fcqo5ZHh04il2d7l1zVVNqsDWywJUMkmXhxH0VpHCnWXYvpwErKU/tIavvP
ag6IsemXw3gmAlL4kBkObnZpLjqBQqZ3J8x3D+ydmWb2OAoNaOtkG7lr/qVf
Eu4L06V+F2vwK/ri5dUPa49fNkVP1N6XvtKGPX0pIwqbquVFlRifmdS36Rge
qd4POfIDcENe83INoE5giWVeZHA3yAuk6juKdfsKDA+3+n2mFCuIngHh6Ie2
qSJVPn+QbzZieVd1VdojWw5Gg3VWvRK6aY1Ryuy4rGEgTPWk9lOm4qpWzexx
R7TkEiSHu4fKtkYpYIsk2jYSlwwGICvVjcg2+KwhZjExh9vGXjWlnRyGmvJR
TRuxsLAtKeOAfgoOMMLYe2tGQOH80LCRs0OOcMqangaMBUqAkGzmo1oXObHZ
Stg/CoWEztPV96VRIA2WtfNHCIuagZPmCne6+fbuboe5p7U+x5ptEy6sO29W
Dkk4mAmtJZzjq2R6joVhfcpZ691uDxf6x2+kBcXJLmjhmoevsT6nw2MnCWzs
M9mjJIt8SsgEWOV5Oa4MxnEvAOrr9dWL/jsNPufiPgb/PEmyVx8LxVTDhvAd
8LNUZDaj/o234T/YXAedpqLJEdU43Kijo9K5j2SLBBiViLx6EQ7ziwNZxxRj
u0X3+JbET0SNsqPUXjjqtbYhx5G+uQ6/2jxanEzylwe1QMmpwl2bjz+DEkLi
u8kVGAQOmn8oSJ+HZKzHeNbEvOC2mG6G9syS94OQDAehr7j0e/ag/KAS+4R0
u94uXjVxfEaDsOOm2Iuph7cO7zZzlYtCLbzQ55HA4oqoR2U0EdVq4RI52p3n
yQD+pIubfxuteFdiW6/xdWIZTVikavuvnpKhTAHWV3cCUic5qpnT56crB5f/
i0PV+IdqFm5Bb7dcDaeLDMMyfnZOBhNM4LZTTFoSuJtCU2Pgcuo867NxE3Xe
F1ZVxLxVHUtBqF37rhsND2uGitEghAuRzXxayEcr5SQ6MRq8fBiD56m6GBJp
IdsKuYLqi9K3GvFgHk7PJ2SQ+E4PNRgmwzuQ65cZztsFBHMOhkaf8Ro8Oygy
Wan1Y9iBISldaqa2AOzqzLovZJjHDzUU1FCeMgjr92HOUbxSlMzNwA/zch7j
qwfGIeBF4h9YUTtCrO0vKXRNWGhzBvR66RDSS3VpU62Nt4TQHb3qORrqM5r6
aE0o9mcx1dsDGLklol0Se4DSz9WSQ5L5t26jeAEkEoqVcZnq67ZNKLLKsNsd
5PrILPboTLK3i363HVghec9/H34wg2l/O0jzYK6M7qEZPUur/KgaNmzu0r1R
N1GJy/Ihn+Gmb38iIpR63wP7sEC60jSSmyXAvIdhRmwkA3Hy1cimGnA0bULB
goC41s2+hChpOATb7Yy/g1FrclvfHLjLRPpkDSHd2EaYkJb1iUO3ukT7ZUny
Ozt0dRfyp+4Nj9EKteKoSiMXPvXaneJVFi8o0u8gSnYBwyQsXNj7UUnAEno5
iuOt2Vply22RXS76YZYdGKZGTouZkqWvDwpnaVZ5YdrU0iANRCjb/ceAyjRr
NzTtYQp3BDMtu6OPQB0njenkg1yUpUX8OR/HbcNfLatdjKBy0yVLvuMWdqu9
a+07l+IFCmQNpeWfD2LuTudSwWcfQwWbLta8E19eYRsDrPtrDDEOBHngPHcM
agcZyihYpSy9q7v+68cWafNdLxaQ/ZY77PMkYY1Z+VbDB842Fsdh6FR9HaKC
A+nyj/SDA/sgjUdtg0S6Ew7jBmcGFmCFZ/jObzWxv/uzN7kpLFd/9IQAwdVn
K3OSMScJsiY1v2nkxK5lPbQETdZAdHrED6cse/IcsFZU5P2qOVHOyRWpQLMI
UMCzAtJUnM3WS9Ivf4D9/ZxUakgCI6Xx9vP1x4RvWorisFYXd9euvbxw/Z/2
2MeMz0SLKJdweyNe+q8pT+kyskgMGqKQvIf+A6NWaBEgwX2Ub9oYi1qYeh8p
HMyWECW29B6qPr/2s318yonGxVWPpy/aCH2k11feAIrn9r4oGgwkbc2sPvzG
4oqxYcrIkveV5IGBYF7YQsORZP9qU1eKGKIhBVT5klI/mXlDEMObZBIM302i
Df6rW0f8VVJwfy7NaH2wEKJveEG19G4M4a+KT59wMFLCdfL0fZO3ZYRQ6JZ4
n8cjMDH6DLbLJ3bo4fNAgCnjwuWveNiCkwYxcWs9Uo6Fv7HSBjdi/Q+9kk4b
oMbJY8OThmA11KBdeI28i/l9K/NXFaPmB30YrnRe/FoF8YSdLn3h/QtomsCF
HRZ5s27xJWjEJGYMB7zf6WrK1wa3WiS5WYkGcofO0nUmz48i0YQZfE9ya7Em
INLg9uKaEX1OOO6p0+xEuPCpcy9i4JDrZPPr0op91Egkn4SicVdIfgRlzuu1
ezGPxpFeKBOdcy/NdJIvJ7KkpeCZPU1gQT9OF4PWby727IRbTExlUmbaix8I
XWCMu4K3HCSjUxJz/4DqGfLmTfJ/s6OYGdD0RLc+AznYL7Jlc9OOmNQDxBT/
ql8y0wvQTAMIF6z5EzZfXhX49MzfyKrTEU4zLvFK9E2U6KJzrXekdcSCDM0q
nCCBSEpQ2peQsBIgxR9JoWBG55IMZh8Ef5kZwwKf+D+nAu9x9zOVLdcBAe3a
ZuzAywGnKA0pH5OTIe19SUnSwT0/zrzXsa6EPuOjMYA44nVf3Cy0TTxyIblS
Wv0DXS3yvP9P1MHQvXInBaFEyJeVb/ifQbmWUoF5ELEZE9UUYlr8MaeItx7r
yWZrs8AqBqzue2hMIq8CfkjT86YvgHsF7P8E+owkvMcSxi0C8QPYe/C4K+sc
otHXWiYHWh3JR56NCMGyRpeOcmL0TW5XD9Pi0ieo41EOXyq1pt+xoI8YWoBk
UENYXGaGB+QZXAHLO9wHg+Ty1yaRfivrKsVEQvaYJiusY6HrlVmfK+mIF9xu
+x/LqcwbQ8SP8eY75cwgvpwvgKGBmjPMAHMWNPoVtDpaDd1bcBHyDghLE2rg
+Y9hJkRApqXxznjiXWbJISjwOryZ6ciYOmQznqO0rOk0e/04tctbUrokvHwB
zn68N4aaTnKK4awTVNGBWqB7+2uRr9BtUinBfztEbgUawETZJRNAxGkdXdmf
VMeNIreGA4uK2WArpvjf4K0pkB5PCD9swYffR53tWzI/OPrnwyHE6XXjMlFF
dPpuPxlwJrIW+BCRzbcOduHMIFHj5pf0msdPdYOSP3dnHcCLOmnRI1cjow2u
WiTmn1Ih5/YOpjKGS/ie3p/eSOQKlOFAG6CqoWIc9XUpCGu1c4EBorW0B9KM
xogF6fNmgiaSVJVh/V7SVrnvdPpAGlB9kmi0TrcrktQu3auFhIviijFD6MWa
xdf9cBhogX3uf8119y7ITDucHRn0Sz38jC2xVQmFdlCj127jTZGDQBOVZYC5
mE2QPQKs6EpGBzNl3HKYyT/FNL1E2nZ5D9JDg9+HRTfetHSn4adrBf1xNZZI
3lzNH/+Za4BFnjLkn2ZIzjdaFyz6g95mLtLmOJmIMg1a/ElUsPBqtZ2YQiHe
E7NI/2QJuacV3B4q7VbQHKp3ZjDP9b9SWNv+XShoQiKFyrg3NTTuUZAPsSms
cmzOWnsvjODaK4lkN7xKEaUlKrcU0c92/RVRaA5O9iXoL06wPa/0sexhVyQW
Tj4UsIqU9XW0bNhjSTvFm5Fz92iH04PPmlI4TLZ0gR6ySxmj/WavuDq2lNPt
qtV4w57cfZuECq5uiL2+Z6G+8OuOD7IGVcdE74qgFRyXvkNU5nE1B2CKtnjL
V/CjsiLWBzL3PTndVGvgvWt3YxgEMZfaY9nJHVAj56vmjdLpWeOZI7Co9kLe
8lCQB9SL163XpQiWl9/nUY8UgSm/y6LSfwngywyp7gxdyJSkhhxP4WwWizl+
72Y5ABLz1SepOr3YbyZRM1uD8XsS7sWlMRM9lOBE6xRVyZemBGJRuGLP/FEX
8Fy+8RkLBou6uE9bPijrDgToXpM4NoS8Rb0Y08Of3qKy+YfR62xnyI/ottRc
N7eDIYWXuAWyHJnV/IrXIuY3qi9XfYah3xDrHCo9a1FQfKcya/NPduHDbmW4
HqiBGjOzy0eLJkO+Gsb3rWYFPldlwEJpm5YsTXqi8I1GHeFHKS1mJvUIlIdh
c9vSiAvwaD0JzT4c+qXt8CHyWbwoEmi+cQKhXvh5sUedcbjBsCJI9U7LGLPD
81lVMl4P4sqhrY+zGvmh7hYSu0sZJJXcVDSP1n3Z+lYPlYE4+MWZ8qKEdhri
diRoNvspuCpzrEWMWTRos2KH4x+OtHPTPYv9A4ZAzSz5D4r/+7XoaSVM1+ms
4X6zfXeKZUwenOTBHj4EVooDJG3rSRiEpnDPoaI1Eq7BsPwIiCkIqyalY+jw
WjxtbRYit03dUKTUnq7Fy0ZbCKaxFMhseYYrgYiNoiUofgFKVbVQTUgM1LHW
b/ILnrind1V8x9JioEH2J498IIjzJ6UxvxG672g8uT0cXSzrhFolBLn/wm8p
JwECdlZEhE2HeEmsoGDiPjtFmaB5C74axIXMIkMN77/2jOVi2xXS/+5pUWBH
exyj9H6aSnwIvES4VJOWbQDkDUjMeG9P08Sfufphxrij7la3dQc6fIvzpedA
lROriSyxCMZzoek/K96nn2Dentak7vLl0vDXC1Zmnyc7WkOWoaCpic9DiSwa
Mjkyxr5t2TKWM6HJ5ONd6C1kFPLvb/Fpmih8KVOFGdnn6SCMwrPL1Q164Vl8
slSGR7W0/8cBCnZlm5an5lsBNQKxII9FuYBLJcQLpql0KKyQqQmOO4Dfpcqq
RbEWHTo4webIcz8sm/T8uuxtY3uxskc7Suj3j50FJE9R/Y1ouVBvHFkwmsa3
5Z3eBvhu/vPxQBMfofcNxjTW9iiCcnNfwMK4yqnLOK5vsbLqxO61XwsH52pd
aHJr80QE+ugxIyK1EzFaPt7WV8qF2hSSjUAy1vBFIXONv669RtR7JK9P2Vhc
8RgKK8B6zHG4G//uIFDnnlHImNMphgEy68/tGYEEwLJcC4kM01C3K2he67O3
s+89PneTt63mMfUzzhAuHnyOjO9CKLj+46e1m6UGo2TDGeGqIpJLab9otSIC
SHOA7oax6LiPuYjTh5f0EG8X159L1boXwus/+wNDOOwvcwQvUZ4LWxR1EmwY
Zdc8WJH8NziIRDIUnkWaaF5Xmtn88/4eCJQ+5YfcnCcT7SVmbcZ3NWPnrO+d
Bx/4MihhmRa4nUsHezqDL/fQKeY46Bv5r04FrfZlUTT/ZuwSc2gjZeHCMj8m
4k9H4F6ek7keCxApImwWawwKLj348JLZoqK5I38bGzflzC+olHoYIWUTIFmX
dehzxL/GAKQn6G4I5nvY4h8oa0f2mQwW32i/eZELyYd3mdmGEMd4W8LX+Jvw
cI6MqxHs63hzvtGVgLT/dgo1OmVDaJ/eXZ23H4ybLsZQQbRpbZG3w081KvGJ
TGx1/0UEJhraBJ2yn50FeEY6vdx1aypsl5vfghJpbv/5tPiQkY83Lw6P1SGT
ibMPdIiBYNnHOW+K+gdRvSizxMCYlbn4BkNAVxI5U9WybzxWHJiuI+DfWlKd
8BT11kPUYyAyN6+Lo7K3B9yxmqqdJjxAs8cVAX0ZEllgq60xQ7GE4h5w0inv
7Z+jRu7YfkGrYGbPd1R/RqnpSVhQX6QGJXVlmgCRwCw5I4W1GiiiRqhib4Ye
VQGhSSenQtdlgZJLZZQdQhqrCEuRbxcWm4BsNa2Ry7OODChU3lT7v7+ffwE3
dnQPRuWfUxyyMmDGQmVilAQIVl140tUsEFRKyFJCkSPI4nQKTm8j3VW8L2xj
xCI8ADw6LM5+DaCmftci35Y/uv6v/4LL0eP1tXw2P9yGqAo4HAEN8JbhKWqE
7QpR9cJx7umV+SvVQsheX6U09aoQh3gaSDdLmm3ADLypgtC1mpk+G2lDsBDM
64Jugllzgx5Ron2hrnGbeM3Xqf07iPnZ0dWbFXoWv1Z8hZuTk/V8KnncgsAE
/7JTQ5PucQJviZBAnE57oJrSJRwU1zyeZ/WmVLdbtdAcf5z2gCVgvJCwnO3j
SZHogdSg5MNZ7L9Vj+8pw7Jb0NaGZ1VaPqamMzFLoSk1TuGCQ5KvCihoeiUg
iAxKDCyvjJ0X0h6E7x13MQex8Aa35qNyAOCFaMpI4GT0jzQb0YI3zyJ0FyCK
zuD22F+jvMBZmpF1xH1NNxY5kJ7CiQSfUyk/u/kb6UvsqbUOFASXkIepXHSz
6mXsQ7Fr/hFScBBEEW0tYhKgcBax1XJ0gN5/2lad93Zt0nT4PIuNuWTeCCFv
P2yanCYdgh7SIQq1w0f0Rca5sST9tSfunBvN8aahhvZOJNK9OCCJL2jqRi5t
2V6SKviZIRc32iP7VUaMgHvPZU/RVc/dDgPfz09lTfmco9jvRI75qp0LyWui
gqOBs5sAmh/JnpSAbo7xJ5lIAIOoqaAw757nRbwHsMv6K4jUXtWyN1LUBxSD
UhokLhsI6hQ2Gdss/gz05aUARNDHrO9HSCbTrZmz3JXuURVuSiCMFvf2pJlQ
unexNKQmutQsBCKD9a0+hOGGShCwED6me1biVVa8KgQd5bVM5xR3p19TtxKt
DUWgfqcAt+vrCJ4vkyXHKgqifutjnrPItkEVIF7qkMQ0Iuj+RVbJ61Q8G0dY
EdbuubUcgABJItVUFQSuplWjJ6tPJKx+LCqhkgH1zgyfr5S8wBmDHw/bg4U2
B/nuaQxX7MMh1geiYj9rUbtPjCyYaENylYSaEzYVAC9gnlUzzeXBKDopAhDC
IZWyzY6GKvprzUUGhoSEu2MRQjncxHoCK2HRMP/simR+MZaLN7zWMpKbQ8bw
oEQcVOSFqA6qJoK9x6HMh8my2/9Rho3Eu18Q4vnxA7RoiAXy/dLEsR6I7RwE
zzc9ccLKqGWnzHX+EB1k5PICAVlOwYdF+YS4n8VMekzgrIj5Qla6dF6FPJMu
MBx03zqKb0YP4hOFFCS2n1iPv77OxFe+dYxKS/PUm4IRXEWs5EQHFJh873mK
w6HkRbe7LXYZQuODVtKeKYQg0cSx/IAPbVWQSJFdCcr08+Kf0hEEUROAlvDH
gT229z3TMjXfdezCFvWVKSAp3WjgeWvno9wL7VJyw1LCMoV4z830Cja8W0I6
rtqPdLWOvktw6+vJGogObRMToD7KaIxu186esqDQENSqy7kuSMDyxcTORN4r
rkFCdZm8WFzoQUGNiuMbAxWOmd4HihYnUU0CyHjYsDoiz7u3lUiu0h17EEaN
MrFYXcWuN7NNSvr9MmFmrcU9UHMVnbu+kJ4eRZVCzghnqXCott1sne2XPM70
MvdxO0wcFszZ+KXHz0B65YrOwhL/QP6o7txcEvhi+h1tDO+rVAnZTPBD/XWv
rIJTZKtDu0IXIEqIpjHONdzbSnOC6nzQ8KfEhng/0Doq9p2Rp/e5KnCswZWp
ftOO0d4aqv+B1YPLI3RFY9OUIeIhb/HSEWc37uSzmIOeLta5WACXMq68V/8S
dPoJvBVmqlbUq8ZOT0/ccRsOJ0Mt8aaPqDYoMnq+U5wKWfAJkaGzePRX0Cdf
fkIV+fhNfLCRc8VwoK2rn/h5Q0f51Z9hkLfOvnnCUZ+n8/FAmoriWEIqbzj+
MAYsJi/xW+otP1zBbp6i3fU+uyD62diPmh0I21SvXmrTzIClr5Kpjms/g8Z7
L4uLxqiJ3idXoPkrgmWCH6BlBaNWMSfSN53rpyd8A1TX4eM1kS8n0L4OuaLP
+QW0hYRMBb/OxqdHGeGWoTfRmQfVtGbCYMvEcXcuD3l7/rStkMUypcwuq4VT
DdXm1k/YTVJ5ivfGJ2B8XkP3zjMo58W0kNXqzGLtIaXTntFkqDcWwkmyhQrB
Demd8fcRESsMrXphk+hhe8u3HhxTe7udqNtEg6Ytav46OFrz2hn5bIAURUvf
BiG9bbj6bt31RBEkW4OIv2ZqooVtTPobVNY8LCwrrOlsO4Vy4VpnlDDUcPns
eVYDliA9F2rxzEYbtVp/Fs9KnJQsmsDwkCu/5SWMkVejAOWwsYdEjOm/gvfS
qo7ztzMKJQFj9RC2HIFVxh8Ofk4pb0jzeMD7F527SQVkYwe7YYqa96/TvFPb
R8neM5oZySI/PveitgzLlM/UD01MY1D/aFRX7LGTVSbDqqsNu6L0v4zqjRV+
kRnxUca3j8K42TaMDKXma/mvqBGUqp71SEsLLe80pWoiXiAF337lPcHOHAlT
5nbjauf+Vilfd/ETVjgZHtd0jYUyI2j7aOe68X+nMJKjQEFEbZI18wBzvQau
LBboZQSMvtjuLkplSe9V2P21gkg2eVtdr7LuhAg0237g0kDx0Ha1YJswY2mq
CcP7SGRxE8TbLm6M/3Q1Sacb4AzBD/O4Vtl01eHgLKEw6/bEFbVBRr2DfM4x
0OnsDjSMlRwFoKgCA8fBLUvtmcA+bvNfAoP75YoB9W1AGi6QTtfISY+VyYCc
kJefshTEnzNFVg6FtHLsy6gl5YRebZM9crL6c6dmjVO6+LEZ+Pc67QGRZc+b
F5lFKNeFLrK41jUh6fU3ncNP58/8UvKm8CPkINH34qfvKRkAQuhRx3Wr+lU3
vYVx+PkPT+T4eV2nOkmEHR/JXWGH/EyCGysXuT/sJL7Hnzne4xOv2D9bhdpl
LbCYVElF76H1+L7wZO+zDCIYUjXhCkZAwKku+2Ob+18BqIKJ5womvuqLAFeF
XFvQiZrWQxssG9v8gUP9PLEGIZ+6wRqzambRx+5QNHrSmRFb6YC7hNebf+CA
DGwrgb4ljJnQJ6ZxxlbSPKv+PnOYSZE9z3443jo3xs+jsZj1zy6LUM0Nnzzs
ZffEt50R56NiWAtKuxF+NGe5V0XU9PIQHD0IqTwC5Nwu3ka2ISex96+WV7FM
98GwDwJ5r7UxfvcWsEzeeXSmHl3Q7xePUJNYtBn6cRsM6bWqB23Af4KALkkH
cyB4qbZi9qeTwxWSE8FUVcQ14H3WIP7hGOxcfyAJgp2uJbbllrMZlRRaQ8NI
VBHrzT0mpJEzl9Akw1egDp/S+THE/JTZQU4OGzWqkQcnvyjSKtvf3K2HUxOq
6zemFGnxnVnCR9VFxULpF2JQp38b4hYDYjzxUyWG83xO9JPl3ZR2ckIAF57K
D7UozgjePmrcZraz0PzQ0KZ2ZcvkvYfT6F1ehYH/MkwfSI4ETL1DBzK0Yttq
tugWVmVMLvsFWQggemDVKZaQn/uK86WCLq+U80tmIcfdvfMqZt/GozbuBDQm
Pm8Y1HfUhOYhsDQCS9cZI4+6295Kriqx9sz6nCZ4mDcwQZ9aFVsfO0GG+XRA
ggcJ11a4ZyxmAD8doHUKzRq9jvPNYGb5pI4M6Abe/qtcvMHQcpaPReihoBHf
1drLotrInKSVGq98FWoe166J336NpH1DgqgaPe8dOStNNbhSjZv824dOvaIS
FPsBLviePtWJiAzV7KnBipN6A+PV2LvqPpvlcb5NJtgIgc7lVLISRWVGrIzi
cQQOFZEz8WOQRBJXQJCPVztaoHFMPiFEraVd7W1t4B5HyJ0s02rbSAZlgXlC
jnLtFaKj7C2cD+ZqgzOksJjxWzSvX1BN4PTps5Vw35bFQAdS7VUQbrkqGqd4
usOOGupHoguSS8/6zg2aL/h/IKX6Khmf+6TjzeLMD3VbOnVN3do3QMpfFs4c
O9K6tIWEKQrS41w1dZi4PxeLQVzndWkjSHok/ZavpOdbVNaxVjCIcKt/oxtr
wsTmZ5NqrIAlOtPFFhY/unomZuZ+lYjxq2x2BiSdqlaP3vpApGcJVdDVS75u
baz+tSmgRvWJ8i2eI+PLfU0qsiysuwGO1wm9sMwvSAtiyKfrFgLTPNggyCo7
ytH092KMjAGngk+cbR79ssTotWW7FOaEttwOo2C45ZJh8ydrCBztJkk4Hpr9
bexaUImZL6UpvZnqpeHxEsvlRjLspJV+7Of142V6sM0rvzMjJ7+l6k1joR/v
ZqzWp3nhatbHHPg1up747gMk2qcm0rzSnEDmdRqgBYYpbPoPGSQE3fDup1Oh
grDXQKgpTuEnXx6ie2WGIAjGzxmvVnD9VmzH1/ab8uU9wG6E7+R9R503Uw5c
OWAeMXNT28aPKOAWh6fO3A08EqImV5c1pkdJ6M7hKnpywa8fanDoJrDYcsKr
BH9g/fwKGk5UzNFpoDJolmNp73ozCvhy7JjHQP4EajezXIobFNIa3PrxR4Tw
7cQpJKYE8oug7236/U2m/94YKnd1xF0yuLW5tNVvnHjXE9McMEQroL6b24cS
cAeCmFmRbmlsp2e05VWuCoTP1zbFdwIBDKA12hf0APb26a6p/0XSUZRqjHTb
vWEOGH4K/prJ9KEbCMzMLk6QdW4bPn8HQzwZTVUDxXDAfpTBUC8ZaVRm0X9R
/LGj5+R1Bf8rZ7zxWRzal+Y8K3T1SpSJstaYgSl1p9U+1JVq/tu84kANfdBc
JbawcFqyvIz95WT9Xs7LkPE7MSZ7aMPVy/lvD/ucfKXU0j3Q4zLm3elyuKfT
BUky75wbtyzI+6f9zLUX6xP1fwq1Wyw6KafoWey2NZFBTs6tBVvBp4UF23b4
0ti8AqACAEVlRCkW8YHMpSh3B0vDeiLc3Ug+QG3L4ZKnOzHuqDM5Z0OFctz+
dAjBR4V5mxuhw9TLH4tilc0HhBl/dHpjH6tiveRhamw9OR3qqwPgtWW6Ozpw
zMhqszua1MG8pmpfgRj5QBJTuoTi47qMFGO4eOKaNUyi+EVmrvav8GurXXQE
rkUiO+v7nkB1qNvX/2LtNIfms4Cf5piMqywi29KhEc1CxEkO4zGKm/d4zpNI
PapDDVG5coiV0xAvj00liCF8JeTsdg+TDTUYGW27nZILYNaLCl61RBMuB/Hd
08jB248TPbBOBbE9v6fQevgt0p8zFsBrOSsrU+sdWk1gDJO5lZ3+Jp6kRW6U
S8elJi0o/tyudpPZNh2FVwHkG0Ec+uMcZgD/krJS7ubZf0TIpyQQRvDfVWOt
2KF2n86ltclQwcMKNJa8Kw0GPzhrECjy/co8SQpTV7DNPuTBTzqqbzouG9qM
B8VmHgFQnRU0hy8l368/IqHM2Fxvme1dS9yAzHPObpFq+WZGakjw7AD7USwm
wEmk1HzenFb4TBNWXxxrSD4Vog0Ml4sBeaEbR+DCTfRGLDBwZvCJMny+zeOC
TBHwhDiUtp/D9CALCYEegb1BC3kRCBNcqa5knwKquSuPbGV5J/EcnCSVLnig
gfkevyJ9C+XnBkND4aRi/Y0VDkjsck1rUn50oMs1ZD3+qhQlqPchV6a68vUA
gcExO35LJ1a1Yh3uesQ4o5SJPFGM+FBFzuQGH+HhVwb6ukFUGQrGe5peraeC
PZWnGN6MLFPLru0LmAHPBlBJIjqJ39HIKJwOpftuuXmfht3XnlAJqZ7KbAqa
feXmN9vYDoewox5Izn8QQHMgm4/G0oeS9TyYvql6rRAhGNRoBH1s04Ex35RQ
MQYg/zVjU+Ml1yDWfs2x+VcEt+1cYd8XQbMFXSA5sCHCumG7L59BQK/59das
ccvKcI+DFEiFSKpryXCmzrxMxcOYYtoRxosNF2BuolqaODXhoxnKudGfr3xg
wHg2F6mTbRyUFiQrZuRMplXbDG/bSXfSVwg7pHDic2qhsU004l5YRj0pAL8o
MnJEtDGd40Mgq8g2/SRL9tg8t+VLGoJFb3KH0sjzgoq8a2MawVhx0i+WxPhs
8kDXfVkXqP7PFUK8oP2y9jJgVXprwWx6ECvus30jqjiyBg1jICOxqhqg5I4u
1inaCkfN1igG+ga1sO2ffAR0IRDAbqqzGAn0Sw4FN6BllvljUvDSQgUcl2PB
czdzYb/x9LEl0Lpr1nq9in08zeBEIi1WBjq7hPmfbWLFuMjidP0u9vjtsMF8
HmOi8jeox/E3iQfNFw4m4bS3ImLlvaL8SYLKCAj27nN2fLqFgZnmtO480ueO
YsTPp6ly+j1a7UaWAgEcgfRLLT+2VlWBMw08T5siik/NFYhCvOumbWECE0S6
da5bm2NebZ86TZYHDxSHvlxrE16i57X2musg7cLhSvJ5eKhf0CKtXwE5NI8Y
VC47Wir3QH+VkPPmYCSfs5eXAreEAIdtTZ2nDoQT88Ez3Om6qaXxTreGzTVL
6e+Xisx+FW5lhfugKkNlyevMe6bGSVpEubRTAKjNBBI9Z5zqeLMz8xsxTOO6
+i4pqqChY8i/636eyG4w4hm4v1ewhyao4NNBb8LyuE8j3q1YC82u6yvnaDoS
dNqxLlwVBogf8FaLpZe73PRh+nxvPJflS1b4LlEN6pHTlmyJqe88FHEV62aU
qOpyxM2+QWPBdJRsJgJ0hKBEJEPMiOmJPZAHLmjBFdwtag5WDn9DE5XgGgnh
ZMPR9+3W0WPzuQdR7LGCOoALBY3l3cfryiwC7wjSrOG2QVjpSV+/TDXPBYIn
8b1i37Ue6YMa4WC4H47MOHNrw1U/IwfYep7O3YDbhJ1WgU50dH3vPsYBdxHU
WyxfdLcLaP1adhE67YGNE4nA0PrYMc+2MUJDCYnaG8xek4ctuH3hJVmntj0w
bRLmXiKzb2YcqULdejfNwmyJ8UOEOlJy+FK4hifdIH4y2NHErsAvC2sVNf78
gdQWwKwyEDCX+VtxK/SYz+6Zv9LyAWQhvN+O2yKiqU0i2owfj2OisJ4y7gho
Lds5OzJcw2dOWwMi5s2t52dHbHjCdQglgB59tuVq2W4KtH6Yz6UDzqZ/hP5N
/tPZOdx+uL1Jdw5G5eIIeW5PFEZx8BTljCl6yerD2G8PUoOLK/7oWG/vMblT
hofxSN0MMv/lamD1GX5Ky6ND0uR/qtSvCtIPHxuBjDIMnF/RERbA6U71w4Lu
Vj0TaYy9JKN1UZAfdcVoTQAT+NAk7cnqfMdEaxxiyhiOpEtdu7PKdgGELB31
zYvJBzqXnTZsO6WZ77trinkLqUKRUE02upSSltNKQ1rpTmCBHUL2MuqNfC7k
3KVwEWweV4/0LV6kPp9tZDG7JxyplScxfLaSsAhbOsRqJwBozYL71jgQ70At
HSolxhx1jsOJtVYv68Z+du7LznkaIPYe2dqtfwPtMxfMJnSSGHGXVK0FyRkS
ecJB1Td5b8lhZk5EirjT0UV4nzy0gZ0fW54iMtiCL0J2oPhe9XuS7wRQSmrC
0/BQ8BZZZGimvVQ1Vj9w4/e4VRAhOus5X0N5mMIKzdeH+1mBk+ZNVLTDEtZ8
CurjBtDnPrhIQFCpn79j3FtMKnEVLP/MOFzLf1hWahZ1Cc4a+JRQBuk5lvz5
VCES6NeI0Jn++3tWoLAN/6TWnScYqhg5EFvJghgogWAw3usO23JlWqmqa8gG
ZufbOLELEmV7gkIxwVMPvksZXN1O2xQ1T/Dfc29rJ4dufJTE9F9t8GsoEj4t
EIHjoglCp5qKbQ0Z28639Z4FizahH4qahxgwSWRS/Wt1CwK+hhzO5yu/npzk
3cBVSfZeKN7Ds9mPqqJFTY3p1eBZp52X1l1sk7wu9dcU/r9rKc+dY3LfzZLR
Km9DGhAjbk4Jy90mnHBfhZ5U6XiGLenVXCoLnCMEg9U4WKnjm9iy7blJ4Oj2
f/Af0opFlhqV82pngScP09haQL0VsDim/9Wwddt8LYvOPxeMiI27P9vxp8bt
1dD8u8sGFl/ZnUqob9wx+mS89ZxZvzFKch58WhtYSnCpUncA9lUbRuKGEF/e
jPB+TC2t2ojXWR4qA0KNWzzztbXoVz8dATAa9/xcGybcD94uy11skCz19mK7
H7zkkzrWBuYeqHfg/n+xQlkzSsn4rdgS1BZqI/IC83qNI9wHTaV2vxS1LvV2
sedlHh/7xiuk9uafBWuY7e128IbrbfWG3tbf4Ios+p8FcaKnXcGZBhgXhaHB
1sdjmHFlgwZmlPwBojYbh9fMsFS7Md3j+nIZq+NPVwCfTm8pffp+71r2JJuj
JLgB/3Xu9NwoXUkfGfSoNKlraIZlxlT78RRfTGeqZnH2EGwzi7Rijb7h1RUA
yoUNbu+nR8Bf6TWfKUOnXWj9HRhAXZ2bLXNNQzgyIRGf55FH3TKaAKDHo6ZG
G4YkWSpte5peIN7/AaIyT8mDDt1hBq2KvOFAhrAfCSutH3pUzDCusyUa6BqW
HIwDVl0H7U3sa8Qt9nCuA/g+hAcNiUILrIM51pbgxeTaJsGg0xmcBUtXhbLW
kgmMYTUev2rb+7aC6CJV+YcG1Oep1j5Je/SEVZ/SwkA/afCpacNLesvuKz9y
afFWAJ6Px1ezsypT9L22M0b0NnSR4oYnF5Msv8iSFykgfWFCNMudqpdC7CCZ
tHp1TG5CnV+8Jh2gkri4s2R1Nfa/ooLI4F1WE+RXy4/tmO7vy3kJdiIR8BXp
eCd6Z8uKFPCOEZZ4hIKF3IotKEGB0TrH9jKxxtrdlSgHVb9CpDimjKaZ6mwf
JkprcoFBEgdpDrzfAleiv0mZCI8hQH33xFM3jzX0faV3w3p2d1gyg3jLhud/
YtIu3fkpOg4Bjf+WviZUBZ6L689+R6Yln83SpsaGJCd/g4pwXCx/dIkkGT1o
+8/zVNFoh1XmJ1xe/gb5VnR0qZ86skQnSXeJ0JPTGs6sCVm5KALhrw0ofag2
a5EZDd1W3l1Rsw5M9kGQ4TcPrBWFnnzhqMbJWz44tcPF72giU3Omz/Xlb6i3
TbCmKpLuCqXjGFQvMvxbgdeC1CPlhgA1ebcxqJ/TV3Bwkywc3SegtnylscTZ
9o+2ea2kkShLsjtAngV/v2z6R2xmqYOWRDYrQ5HgUSbWeVS5IFQ05vBsGI1v
9BmSaaqJ8cp6FAO8NlFuarEtQZ55MkEVOJt+7KiBnqRsquuqbPwBT//oLzjY
kel7IOk0x5CrQ5qmcwwd5EuvqW1ptJTgqDrD0FDtHyaaJpua75mxs3Cj7v6P
Dde6x/3fr0jDU2i810KFLTCdrBWfLWabm8wfqo6tvUZy6gzwFPkepET3OG/f
dV0D9opTBkw/TW7AiE8EdKgnB14gqRlPn5IA84fRAJXcDXTgM3gLXBIQ/c2p
bGnJRsgA5JlFsshGSn0eFuqi3j52G9M1yOuZVCl9wUv+n7uZjkgwg38uq1Ul
VBiL1HEYF1sbC11r6PENEnapPaHtraCH3k8wPOnfiQ5BUMJ7WgEIHa9uEow8
aMXT1suj9cnsHf5haklbA6aummxYF8KUc5ByJEUm/jBeG59W18jgeB8wu54k
VyZ/lBWHK4F/r4ruXQE9d4k+zyruaBTLNwm1X315m4RVHLbuSPK44D35gs5F
7QpHHoa9EXPM/x1FLKkezCR7/j7imtzrgLu3+UomyXI3DciNthH/IVoN8FPv
ehLWg7UxP7aylsT44Nt+qS7IwXkw7fMBe7QmPbKWjI+Ri4FIcgjbQKIRiTZ4
3Z+pPPU1lz5kRSTIN7yxM3hcE2zZum+zQfVcFU21LFz8nzsshsrEc2GIYKyc
xVFFwoZXsMYWFcnuiMTtAXTGn9YWA+R0ox+o/uLvKnjsi54MorAKhBMswYyP
xF9DkIDpq4yVWfxa0IFh1ZjPahwUK0fwAVdOeTA0rtpLMCGkFjuFHXa6uir5
HzCUWWt8oh/A08y7yWISyaIpruZg2LpxDThnc/IbNtXaPi+smk3KZK2OKPr8
sv9k1IAxJVbA0HBo5Wl2/fxeD2JkcCAMGsFO2+vU3LBitYEbLaD5lQQRQEyC
O1dqfiXY5iUu4iuLInQfLffkq8orY9WC5YiElr+4sJmO7aIgfgVVVp9OZGfO
hPHfv+nDODA/wXhRULCfZ38xC2UiCabFqvsrQ8h5PnngdRDf6Ck8wjoc/xHV
P9rqlYM1B+IflUzZpa8uGROhnmxKWBB6BlyE4iFPg8j3FvbtFYbbLAhUgQpP
31Edu4H2+OU0w/oiBu0iX9son6Y4ZIwSdf7fRTJ3WcRhkh/oiUErCEV4Pxsv
eFFQmLOpinKWl6X0IdSlFwyKKIfo9hX5mR3Dan9wjB+YM7+Nro4dzuE9sMh7
rViV60EH75ikqSFIjVA9Stlfjpy0CJ1AoBssidk4KJJuAhL0zi801dPAeetJ
MPQfBd5NCOIJdrLmfD6voGlMD3i4HUgQX5+qiwy93oCUQKwOUSMawG5l/sQp
PmFz4hT6FtqhbNIFPSBBgQ4bocTMblLHR1zf0rIMw1IJFvWbSTRM40D0wJQe
HDq7BCa7olYKBolUfZ/AyUW3DagP52WNHhyF4jRY6cIHJ6HZJmFt67PZ4fhD
j1SnFR35MtrmkqohzSsmy7tvfN9SyoieKxWh7r9JpsQjpbu56qCFiw7sZuaw
Jyy8lE6hpT/DmM1laK3JuIgQEnjekpqnV0rBGkZYMMDwtSO9UI8FbpgNcNR2
fm50LHJGanejfIU4EAnY1ZEC5AXMx6kMDpFWLo8DOq8p0OeOG+sUT8N/Q8nE
3VGPB8n+MXSFXQJ+2Th9iGVDqESBc5mN1UhMFyJOQNdlQhoQIgQUWUF8kl73
AbDi0MF+kJXzenWKUo3kCc/rtIsYnTABcnsVxUZulY585a5BhjX0/Pj/8fvd
A42wS6iQpGNwfauGzhtFJh68kbojEKxCupGxGlhKXrEofSzd4x3wBrbnu3nu
Bc5w7duBkXNVyaYCtzA1+yYPNCWtNRg4w2tSgJ3eBsheFajNVQQikzwmkkeX
JK3BSQAPP8t3GNXZEg2LBqy7GXDCauMFotu4Rb8QX2FaKsbnCpz1PZPZrepC
55V05nGS+2YxOwd+UBQSQAC81VJk/SrTBiw2I/+bFzFamh5W7djcjWvp998r
joiz39153tJZunC0BRcPY195lanPKG1wCJTCgrJX9u5A8vvq+OfCeUgrxvLQ
HB/B7AMA1y2Rr2oynNz2Ib/0ChfLEnXCBmrKr2BdqbwP5NDuq5pSnt3RDOfl
IzBjJt4IPdlvPEmMReIVeFlZumguEmPX4haCd+jB7EaSEH9Y8GdHjBzrBVJB
7rregs+MXsosevoKXk2Ppq7UszkKgqtltRm9AjDWibg5zqxKLDTQrDQzoUSY
H/ACQrZ49pZiHLQZ1o8JmC4NP3Na18YZ1WJHKoRfg808PFCnm/CTRbqUsV0W
PM7Ut0DclGEnMqodTeQExrEOxZWpDonkfUPIdBrotcGce+KjCgZahpzDGpsV
Ju5qmnj7rRjnHUpeU2yca6ZEuvZuS4o8yrPMYH7yQ9yqVDRfErdfo1lVYrGH
1giX61X1nC0ZVJSC5DSdLnXoshu1rsI5SxfSyebS9aFCulIwophWTFtBpqAx
IAN6i+zP+R+RXly54WLNXtFggx03MguD3q6Ylpf9qkQKl/D6k81pxgIX63by
sfAc2x749zpSA59earYe7luQH5J5BdSF06ZZn5Gyt65SABroXWLnR6ZwuTtL
XldDnG8YTf1fHLhhIYF/u8jA71FT5YyuIGVMTuSCyNwd7USAqpwiyVxG6+n4
wSOLbAzc5FiJk3UqzCfOYEs0sthN2G2RSWu/ql698J5C9YSp6ib/wGKK4G7W
HhhbHtswcrqSJ8k5H/5W0EXGcL5SnYnRwn3cV+9CjawjAInnXyQP2wPjvCcz
JuyaiswqVatL4d6bYBHPOp0MYPJzpgeVgholqwqMtQZR8CuNvviTe0ZDIgaM
T5kfxWAFks3N3tICnl8jvMeer2VnqldzXhCY54bMwCGYezuAYZVa9i9/ts71
Gd/ABtEeq2Ur2WvEMlpIxwsLWLs9PNOLFGJgljgFNN9hVSD0atWBZLYiTdSF
3Z9P7yan6XBCWi+vkHeP/vNpyvAU6KHUpNKteKpQzjYyjIHVq12aQQCmpUTb
LqdqqZSJUCPDt90mq9yN07q1FP18srWhA0PYynEDz5pHFL0na4PCmdY4xU7M
aDQYC/M8JpJT4C847ocq8QaMCw0rm3qjOJyJqFF7n1OfIZcfyg5L87v26RJq
Sxp7gTmOUUsbslEDH3B9S8LU0RIJYuDjudJFM5Lm5gAquDVrv3UKGythrxdN
wh5JPcBmKL8mWJjSWYvfy/7iVI4Cgg1qkYLwl+eaSL3OGIaEmMt1v3hegGRM
51WVudxHTkGEdjiPlB2K2TloOq/lHgHbqrEBqKoKKUZgZHc0XjEZKuqw9qR3
iBd8b9icFWsXv99zRXMqCHD8e2+M4UxoHLPkzkDgZfINty/tqa16Qdt4HowB
RwAg0PXFldGdf4cc8LfKo8dHKjOOW/TyH/XiQ16gGDho7+0t7jqUnxMFXCyL
rsCj9W/WTEBSX/YBE+SqTRvR11OH1oRNn+YFMYGtslnFIXMYk5JRhNRkwyp4
qsyzQR6J7DpdogiJHX9obZnxmQoOPJxeZ1njdmWwU5EgG/s/pDiIM05DLHhr
LbVRruofJxY93DPK5K0nwiyf2dDVY+gj55iCE4AAhI9MSj2/GYnywxvnduXm
3VjgBef7XN0+DzUfHPNH3bSUy8yuyJivMiCOpF6gdY3utDwPG9aYWMRUf5O+
hkDoeUwGo53fAeQ3sMaUlVFMrT/onbPBpSeTMFjRt///pnfiy9ZGTdhRZkgl
cCEpeBcQy+luk+SkUzYLkMAsMwcpB7Km936bUzKnNL9mVjvHZA7r47fEtdZ1
90ymo2lIpxpQACD/UVGlufFYi1/YlMVPMcgZXi8zaT+/PDhhuSFTXMsPEJfv
ZUEjBNUmtHecS9Yzh3zBqrKSEAIAO9E6mif71jPTsgaPE7C4SOhl+tXDdGhw
XoimADzJF26GOcNWAdMKBeHky6pmwgHBAX3gkCv4VCGjTe7aC2IyyfW3TTne
vyqLKf3ojC7VTcbSnlr57d/uoVBPReh6VT7tp700kECB6ryX54ZeDLqo0aMJ
dVwyvNvgBDHfSUW9s9SCMhNait5Y3EnZlqqeVkFOSMBiYWfuXjFbQQDumwUX
LweRkZa/S9lc/6mbij7QAa+opATC1F8yLHmmUHfbjrhi+So7qyHxbMfXzCrZ
N97tBswNfU3MqZijxHvvW4RV/l8H2yvueOnthuDtEoDItddNcNOCSu9XF+wl
0Ct49xkuKAcvS/DX+nTYA2j2kYsMyOtXSvq7J2rprgYKjYuxBvold4QRXi9x
1FSOG5/IpF4/wuqxPNnAnkLjDReCxsusHSkUey1Gf6IlJYlFseJQ5CvlwSox
AlgKH2nQD8haLtCiWIf2FxUkG2gXN1SClgvNZCOqb5qEEbefBAbwkzRfL2DJ
fRvgZZ+fCHSPjY+LPEiIW3StbPUEtWwVIXFiqgIV4KQO11DCJsQDhFU8gg0q
EzxU/cDjwIXDppSgAcoIvtdi9MeQmGr4cHkoO8hYj+qLSDdbnJWvl3kxNbTR
XsZxqNemlEsCrPLl8jl6p9cHLx+1vFDmrafAG3OkMbRsJiUO2woAEPqrMfgJ
ykn1RXnZGUCE6UI4q/7Hh3vYarki0facOd8xUV8lXognfP3B7CDB0yKizMEt
KYxQ4eCE+iVX78SV1ZBTG2EjqgZud36+wZ0Wjsgzvcus5a4uYttUmXgGLTYr
EeYzakpH0NGAUS337AnoDEdTNn5tRIJPtd3hIT68hoGYl/cgCpqvINBpIP30
UxViNFByHJoY2xyEPdR+3ySJXOw67AqNzLGL2Wqq8Hht0x38jgIwU/PzN3mH
r9A/MQCIf7dmePYKXbIIbbgtkgrxSO58ZPVuDEQMe0TGRZ8tqkHu9O25fYbH
Cqa18GcTzsFJMEVoEhJRwtR5ZPPn0QEOoX7NHaQyDwJvfrvVvBITcJaE0Kl4
3sGmBpUH7ZHaCmvjVdNyZ1Pn3u+y/4msBO1CU/9n5szqx8YsH5AU+BlR+nEa
rc5aKaSxZnYX8rWZS+Vj2QZCE44o202bLuoEAJ1ySQ7EMtyVABMXnIxUd4sm
r2LlXoodaqTfotTG5GAXHibdk23BD5ZQU2XawHqKXqQ2ISlt6MIhEqW01eeq
t2pM8tc6+VBztmJ0eIBrLRWeW6Jm1GVLKomTFQKC826o7V9ARCFMmg2m4LdJ
Zad9tOoQf9y71FkmSQWuviWf2uqOXy8cRMLPRkUphw5JNufZHlx1xABL+ZS0
H3hValTy8VnwbFCYF0VSKYOPjMBCknoZqV5j24zTBrot7rNcWZk1BVfQ4xUy
sPrBAzBSjVe92JgxnVjvwwdGalHJ/iZszldrS/8HhACstyNUcF2fn3iYppnc
MDL/o7IzPOOT/hexd3T4ctn1YOzuICi9yYFf3uyyco30tjyitVlH223w5+KF
7YV9q9Cs3UHPJZuDIVJgg9HvFszRCL76Q80+s1TEXnDPnZoW1wEd/8Z/l55R
iCequkZwRI/pnwXu70DfJbbhKe+FsZXeBro7ZYeTP22fQgZuH35kX2EC1Xc7
rmvlhXLMCkUtaSkrUILxvX3ox696g+1hDpurqZSoMYmwPsrctREwWV99E6sq
d9aFamCB6HWWxC9UjkQEJrrDkDVmuWQBYHZuAEracWLi+BEDGc0R1HEbwHAG
4Wb7EbfEodWvaMuZHaPIC0Pnch8ITimes86HlDLahb1jvXlfumKGE5FLkH7K
pJd8eR6BfuEfoQQqKcVMAsxr1f8dyVTSGd/I89vpSk+lZRIGJPZBmUQulvss
7eWtioZSVwKe7ACt0p/fWs2DUutnj8mVQvynvoxG0xY2TkhnIzf+4wKu63hD
NHxG9oo/G73vtuPaQlc7zf8xb9i1IfI5VPtPRCQAos16FOIjkDT/SGnVH2Dn
xD9AeyfFLvAya2IzviZWB9liPEehc/cw6l8kbSfuW+waCI/rOzaWKb5wpdWo
qbvwvaTgOw9Ff7ExH5AbGnvrze/vnEDktF2hn6MWZij7UmeqeFrzKQyIDVsO
rszYJ4zu7pUZqL91XRHyGNDBtUSil35IRc3ftlLnPVBgtURR5uR7V6AsqCc2
5CN/aAix0DV67cquEMyK5CWnT2AaFW8lVr6bWv/37pVrOlO8Iv2J7pUGGoWR
2eZd2l5k8og3riGS7aRmSX5p/2/Ge7scBhT/wSFgk/9vZXoRVtbmtmkBvbW5
u06uecIl57J70Pyf5SeBVZOAYlXmYxRNHanqFymRwMwqhy6XXoGnjQUzWj27
id/ujcpXsy5caDWGEYMzkQxsee4YP9a5GS5CSzMcKTacNgLe4BB+X9l7XfCH
E3QE9tS1soesPz8DlZioDxw4T5l01/lJ8rgx60a319Npwc9DMcoQs49flZup
dlfbPseJajTMZYnHLqi6bk7GGd+PwpE5Ir8aLdVXBnqXfg81bcDPsxz8Zyd+
HO2mJKzJflkqVBaMjvUd51IV8ZF1WSkZ5B7C7GGvE+l1EX1U3T+5pihVgFmK
1OgzvsdZ1kerHp3Le9FXd14gVaNts2rIT5gE+X4cEOBCJJ8HnQic1uLHv8sX
J+0W1g5FGMJOe83QJvJO1vYLBcJkFHc7dRK9k2QTQ2upb7rCi616YjoDh9Oj
3IB/Uyzim5BDYYu3gVH8M4SUHpLi0xg+2lL244cL6SUDNswasxd7iF/znZBy
fp5dyORduGFlq8SoxYVbF/OOVkf6EuVZZcAcg0xLwSMo95q+gYLrqv8JTBjJ
4WysfIY9WV+wgbEveLp/UA234y6DssFiHR6JGU3SJ0Psv3yeVO6g+EiIZ+sC
alGQNN6Cvs6QHc/7vOvnW1VTfS2oGVqyF64ozU3Xo/pgqIvySCkodTp2FwtV
BeXaiQzgk2PRbQpsQiFAZQB6mJJHF7xtZGUeqU19O0MpZZl0HUe+Z5Kpagsu
Hq8cgsUxeUHIaq+qFnyAXMctCTpSD6HkHQsH/lqQ4+3UQrE8wFLRA8AhwnF6
+9WZxQDYxr+eTc8Y1JEysVqpSGK1gEXO7AAjO3ZZIMmtNNkAd9XMUfJeT69M
HiGYBW8U/5wNtjEencRhC56zg6XKRXMkxPHewLEWJ2VQMVfdK6U7WQVZBzoT
2L4OUa5YwomAgG2ceBsLySJSR/rASm8Kt1x1z2nO3v9HCP7XlXEcX5DbxMEN
KCHk2VVv+JrZrD7SjXbLCAjbs8xx0ZLbMsxtkoX5ZVyKt/XH3CaLM2MARaE4
W7wvWXad2zpjHZvigARTEkWgR3iEz/aPJaxavtfMEI0JobuUp/LiXuDrtN4Z
bvcxsSkCqi08GTKKDjLH8nowP67otVR3388A3AyotmMi6BtRAetR9MqtcJSB
2DaICHVPjOKwYHuARLBz951JOUazKpX3KHaSteyNrohIMOB2Lm+OyQAmuptk
86EyJt1TsnWLKAvn3PSE78n8qXV8/WQWn1nicJJ5RrgQ9RMbV0ZWwDZ2Mwq0
JLECnreFPhtLVLptI2rw1o9HPpbRcNMNoirEPiddD8c/Njd7i/4AiW2kDv9w
BkrRpMtIjDDdtBY6+Kq4ny9juEuH31ymo7lXx/+BsGbOXQLPmX91jqtNwyQe
PPXp7gP+9CRuSv4CDtHo1hlLCJluQEMDpRfECVsIpFVpwMGgQzAGrcCvo/XT
xWe7kpKrfCHWXeYKiNGEYXSfwO9BmuwXyoEkv0DdH0KhuXzxrnYtlmtI5YMV
t8wVo7f8qvvbyb86c98PT970d3Q45tNh2cD8D8Lh3zX6wQgPxAgLE15BsY5Z
gQZDW8jGvgLdHRJMYOpbiJ1+Hv+xIGeEH1IVA1qpwckhR1t6mRyDcLduF927
11k6ejO+NDjTG55oG9U8pon6BvAaoSZzZmMv4vlHI3A+I7EjtSXtGxvb/RBB
Iyrji4lIYla7FHWpZnmjB6XhN8GJ+3nONKKrSh6DbKFi3c/BZkspuecGYQ/T
HhwnulH3ji0gvVM7opV7jgGhKKWrPcMSvtFbax4xPDhoGxoV4ZIWab/8HUbo
in2FxfzmfuNtmMpOBziMjTwQjRe617PaJT5ro7qnAkfjXQ9HdlqaHw4PNfWh
jVUOZOVC0k93RNcvZpHADOqgOwjtXpiTnjSp8ClI5BHPjAbfIe68HHdLz8P0
EvtxbjnuTvdLaRJcAI2hbKoznPqPDVG+ta9etrOpmzfxFFeRzlNIzPjDyYot
lmtUviZeIdJydm0z08Xuuq1mRruk5aYYPCOEqNzvsIVKPthRWuTpBGCZYcTL
Red6NR9DO2fHSkIIslCTkC1WQlX/NBMGBpBMPN1ZLPPNRD4j0p/uAFQcBUF0
zmFQoVW+vLC7HRNHiQZDzcRGilezK1wIwsg0QIGP4o4pgEsS3ewpwrhq/vFg
ehISijkAjzHqS/7o+8xVSAu1iTfIH/l7OZjbvSKO17YI9A4WW+h+0GIi6cN5
dw8mD41eARWNramiU6zO1ONR06JpfbtSgxh9CqQ13RwzW+YlT195WauzoZzB
dbVdR3tcMcUXLh/ivh5Oi1vKA4wM3kelloZ+3SjFGctYgHQaaH5CAImZy1J6
7FkOQCBZj3H0upWY4bPKPk66xlcnjeuEBR5e2LB8GuuwZha63VYdV0z2xKY4
prNQto3BPWhm0OL5vKiuycrYMp/JVt4I+i8OnilN1dj95j2C70RxhJCnZRIq
OWAR9lG5R5yzVq+2htxpClZsytSN+PO2QR4W02fLkQx5poBNpTqcwILAnK5m
1Z/kGU6Xh8uTAgce/a1niSXF+RMFGfW/8kzj5nONUZKtMJSBk9zGkkKucKZS
a0uEvhjuXamcuZnxq62Qc3s3hOexQde93+HKfh6FZoFv/pNvQ/SJHaZ160eY
o77sl7hQ03CkD2wFYNyBP+fJCLadjNtCeJGdLi+AmYA+oIP9WZIP1EPT/rMR
AQo5l7wj+YIquEE5G3pdZW1z5vJ/omD7AJ0gjB5RvJ7g8edxUPDpm+dP7J7f
NWXyTttKxABeAnQIsc4tLwyYESQ4e7r82GRwe7FGKfXkICDrkaThpzEl9erW
yl5Q1ZRw2JkLtRey9HeMjsTooOMRcpVQ6SesUzhtzXxeSGUlLDoNq7xvNLbj
nLICWNrtI649YkaagpTYcQ25n7MJ/XRZfWRZuGQSuVFw0uiQWMptwvgV9cv/
w61uBt9TgI4ap3aHARcVUpihuPr9US8Zwo07/hYlwxlwreTjLGIXgZJ9SvpK
zCWfv6FptH/w6hInsfO5pCYXkgp8qY5Id0Mjn7oF1oiqPndo+KUMQzvGifWF
udFt166VO81dmwRp3MQyT+tS8UqQRtFRgB1Mr8gV4tVzbh+guRExpa5RvxLO
rz1Xa+Frozj8uMZebN+HjETwbx3L9NaxooJXSQUMOH4cykAK5Lgc4nmxzxsJ
Ga+eZw/J3xExyx2Oc/3TFz9ZTBo5gB++y5tzPiST1IGqJCHtYt3DL4gu/K6H
ewXPsitSf2Mjh3fI2DuBdHbtrUoI8badsxwWdTHDY7y+Fdju5IV0Triam722
a4VIXQBJt2x9kzV8TKAzQPIsQGmis38paW7XSIRIXcbYGS4mXzI8orQ7eFj7
lB9i7L4q48v82of5Q4FNZI0Czp7lTIqsv+Ai4QjuCPzBMtAxA7tFakouArR8
Ank3YiaFpJXV6VT1bS0CAHoB3Pc+0lkBz091ARFC/J0BJ3XR8/EWjVHBSCPI
lMm3j6Thphu7VhU0pg6Wu4uVR0+3pbfC9WP5mpXMM6lJEwQli3hJKL4kRocl
eG4WLoZQG4t4H6cQw/q282k7jaH/Pf2oy9qAMoCLm0Z6rWv9YLwaSuFdn/fS
2z4+g7SLk1RP3knm7+HvMoEgRHrGsP1pEmPnwBSedbIaGDD/qnYyOZ/LcYdP
zGRjoM4Zm+bxyUZlMyYvkjn7gvLlUlpM/ehPXoJeWoWJIZbG6TeGcYlR34fT
7FvDP7NyVkzonoTAYIIzNiKR+A5+/BGes+5JASnGwEQYg/6QrO4kfGDFNyQr
/DzypaCwCRA/rWm/DKD91g2NfUVjU51FgJMqVBRITc9gd2DHBoXJMByfV/8Z
6gvByKYJd4Qy2ns3u89tvc7ds4H3dDuLAcIZQzWi6s1T1klcPRYY6j9fAHYF
hP2dENSCwhHOZ63BZs8n7VJKXjQRsbMTcxjh8Gx8+nZeN6TJaTQKKfT0zcHr
H5WpXUZRDFyZ1YezZ1MAGAzsvGRzjDeTX01W2Dbg4QzcExvfhNS2CE2c4vG/
Bv2qy9prXmiQ9ZFisbTAO6uB0jkjxP/FbQTv5guYWi3QOOs2UjLi7qEqdxCR
dsCE2wD6kbtOVcujrKquuxWguBlpx8HBCFEXSQRs1Jf5syf+6TabjBe60RAu
3bThpZ2VGZh8t4CdNe8TEKj215b4ZWacU03jkzHKwqcexBRpsYgaOsPWqKQB
vqLjF2xrvsa9onxEGRUnqvz1vqko5ROZozmKzpO7xaReFmXOvb0DuUhLdq8l
qcSdadQOaTT9lGBUnV3rzI35ZlXCyvkYKs22k4N/P/fXM5KRMPNCe4O8qPfk
FU7yhDab/f8IB8tvzytbTxgs4K1uXZo4uNEC9YKoMjjIPQ/IkabZh/EV/7Y6
FrE55AQNykQfZz4CmDuUxPQxLKt6urGN0cbMO8426+S8SQay5CFPBc2OOsjf
qDJgTO98GCo3W9HE1mY8ub+boYqLCN0+e07sGybX7YhgqYL4v5q77vk6CQ17
eHw5L+2goqfi2w7C4ymSyRtA5XzFKVLV8JTWVirm0BL3c+qquo3IXS7gA21y
XEccROg2qSS0B/wboKNSOAwlEajRdTKk1gI0hG08nGcS38UD7/+e1u+LPSz8
ubQjYqUCPyEsqr0v89DE+DmHPxlu2yRPhtmgMDHFD5HXqmgPx3mO7H/8ueT4
SXZVailjQl5qpWoaZA7CTwaPaiqplWnq70lw4pS1PJR113EK/h6mN4PaOHoD
TIYp5Iju6fHr4ZW2gRpuA/Zl3BVzaOSG1LH3gmRGW6xvAyCvgjfPZD4To4L/
SHUZVFhcA8BF1l8Nob1h6JQ1izcXhFMRMYYHW61ziC9C/heDw1HrogFQCLSU
ixTUVENUAmOO6uzc42A9jOpKCSubgH7gS+cv3/p9sptDwNs3rP0R6Cy9gTK3
NhW44XMPYYZwCKDByOp3Gz91po9DgTFMn2orn0L86P1b0Cxu7TeFDw7ReFK9
CzJRvYHQN2C3l1ndfRGKtiDKu5N7x5ZnnjwIJsT8EHBC0NWeUAWzWQxkKaq+
PfvwyeqGJncm6Swl6kc64tJ/QLU9AWmd+Vs7/NToKLecUQR0YK+doWrBHYaH
nphiPbcrtB0lzNuN2ZfVa3CfPqUlL2aGpMpm9UO7ZiBZLbSY3bQXKhZQCcEu
ArcCIORL0ydvLkFJ3Fy6UYOGNygJRQ4REVEovnjSTmm/mdtcYCxCcRjHyE3u
cDHDoJnXsMgsi/QZ+OvX5MmaAQ8JDWfbNtQ/6NHxLN5GpfRMhJhObuQKPS6n
RbHKgvpDP/RT6Q+aDxJkLBK+qOnSrS3Dm//YTaLJFSMCtJc3Z83wdXCpwrJe
1hpl5LwbU4FOg+wpllsDeysz5WBkB5WPcZIibKfrO3IkbCJbiFim5mukyLqo
lCIuVvaHlKobuFH/MpMiiwV4oEXf02J1t1gYeX+0a77opLSIc0iWk+NWulWW
5kbFbffO30vz3gpyaTcNiUxaVHzGn3wxF6wPwCZ6lrhPIiRbg0h7sEXlhEnd
vTGk4cvLQs7A1kIKrn7pDXpCJjUD2gAR8D+ZAZbP2zfEAlVzhnl++0fcjQWr
QWmd0pSEdqUcLibeLLWtI3WlNOpkk9OS5If8zx+3G40EemHdcnqKnzPt70ka
FYTTfIi/UjyfycbUad9Zbnq+A/uUp3v70vAZbS1nepeHUe2n6z8T1EnjK23D
J8wQhhHplIY80OtK02Xpvz1ayPJZyD9VQHEqsOZX7Wyr7zLdaJhK6usS/euF
otPc8DhMzvlNVRdzCcngi5lOaM2pKSmf/GPehVFt/jBIv+7KnPEwNjUnvgo3
E+gHcRLpjWbLRBpDim3qA7veUV4qPRoD1aqQYsBInGeSup1G7AJHUr8DN5SX
k//rt6FfEblJ+D/4ta49DnSwxhT6ZeY0u3OGPOavC2n+Y/GKA8W6mcF1SMu6
ofv2j/MnDEOPdz5tY+TTH6agzpsixkvLAZ9BzasZB+dlgrAr4YnbXIMjtic0
G/ic3dYGrZR1fGgMtXDjCmlQz1v5ibIrCNkKF6+mBsCoChJlc82rrRIqK0tv
6U/CTifoczF/NnkR+2x6Gl2NyBAWeHne5qrRc/f50y/cuRG/7xrWb4mROJxI
41VLAXVcAwtGLbxhGNZI6zOGIEAKBhmlwhHCcXc7o3Os/2QCxSlSXUTwq+w5
LTX+1SBQi4aSQ/MytfsY0ba4PUenPKdudVJZ59mTuEr455OfAOBh40ifrzgW
E79yJdaBO5n2KcCwrA4SlZrJKOwOnS8xvE0q9NWYIjDt18kb2zpuiSvXZyHx
a4RwYBH9dw6lOApCFcmmJjgnuK8QjlGREcgWE/vgeppPd1lNSBb7jUR0Xlh7
UFbhaW3qY+sVpW5h7KUiKFkRpGhOE+WRNnV7iltUvlU1bZd3Kfm9qxj1mq30
7WynjsUN7B7A717Re8Kw3osfeZdo0ODEMSjVPps0qzj0DjUOexs0CHhvVAFw
1inhUgAjh7pFybc4y5ELqxJGkxWHfDAJFNeMQ9rmvTpVhI3FEHqyW8f1rAWP
IM64boUXxUeYrrys3bGKZDPKdXFt0pNHeeRPexepMyywkQaWmWqHYJsf6jee
u7AV+x3bD1IXt2UItWat0gMjsEi3Oaiv9fjsjga/mtZQTIkSeZXsouVp4hPJ
QbEjmVeyKz4k/avwY/3h6sR8l5Roc29lZDPJxeSrPEMFe3YXJUuAqG4MvJR7
8oOuUmJiZfF63OqxSzReH7JoinO44YPo0+S7veIZogtAJOtEkPyajXMXi9c7
4hSGLrlQls4SiPdy+FRA84E1/d3Ddb6g/7IKibuZds3BJMneg49vAQJlYNdv
ODuDY+/sTJQ0Q6Z0sNgOYb+ZHlJEasso5fGxrnYFg6BjjdeE+lSsAA95mk+7
GOzUm+KAruZi8iDuLXR3Mw1JuvVUsYI/73/E4M3Go2HWgr/s56PCtjgdRmCU
6DA4Zqys+CABK/3MWE3g2gLYWmbzhiQeXzIPDJOOzN8OXH0HC3iSdMDFQ98Q
39vzkB3o47e9ZSSwdl3T0WWGWoPt0XuB2PJdcsZ8WtMtrZmy1YosTxDDiBeJ
lUHjLkMb8DZtMmxzW9nOeVFCft+yeub+SwY9A4u72duyftdcK6c3+GSt47GQ
ngkID/CeA9fqGBQj1aNEQg93daOGLsRYglHnLqVAZlSzfoCJxle2YpvjA7Dl
wT2CCMX4486iiC3kzuDH2+zlOJgxDF8e26vhCPEJuF2aq7LmcD4IN0Fsi7oQ
KhVR8D/I9zHdSvJIC+yv2rhdUD0kxEAyzavmpjsPtH2n2xlO8SRFMMFbEbXy
Wk/1XFgD8hZ8LPtlNncLlq2WfH4gUoTL7BZENOxsEnEL/vp3BjQkBgiEmYR5
wfMSrhKqjTxJU6ulyOiGv6fW5EeVp/ggjApuvp/3t8ZqaLIyJV/paWuoxORK
fu36q9VcnXjEEEESu0P1TI+BJhjbCofy9WUz6bQz5wG9cYFyCiwfsMQLuNgj
iVei3LDnBJfmzEI4bsWz26VTnqxL+sUFwvauAWSnJKTW5YZFCPsOKAikpFEq
+vjX1UYK5RXzHyNr9glHiOnpZX8dbgTPdg2GPUuQap8Y7QiR4JFn8JYd3T3/
v7HIhB0c1+bxk79nEy5PGJKkTqbtblMuscWe6k4SXZJTHmkiP1/GCAYQtZ9O
8+3AGYKP5Le9VaoixAam2mSJdgu0QxYE8Rk+Ihy31eymWY77c7v9mqfT2akp
riZOVrKE6U/CD8jNVuYGHwSuUZYwFF0RwdTTCxNfwkGhMtEp2Vsi6AL046c0
b6kIWrEWbm1PbAndJlal3s4TkeN+ag//nGhZ1CLh+zoYY31kmtQzz5HyLBc9
wH+WBxDvmgkXQiZQPgBzmBVBD4cU5igGntutQF92cN3LkOkxzyB+2Ih1Bm9L
jD3ciuAYIn/t1W0Wvj94t1dWG/OzKyYEwWn4qEhP4Xzol7qGdWge0B1CTGAh
Aga2QvAdXIHINO56uqz8QVWV8dSo7iG/3aS4Aqgl6AAywkUuo37KmZYsthMP
BHZPI5M4L1W5+ez/RQtgsEyE+Ko68W22JJ/giHeTiZghrdwmkLaJX9AxErMj
gL/+2IN4fUN3pK3A/c6dhrmL31zUrP/0qCIwKm0UP0lC6cKMeXPRc8f9qpol
WxFL3L7voribDNUCGztcUqE9X1rsQHH1k0o4vCfa/BfIOSKMlrljcIykdlb2
MuCR1VYezR519bHHlk/8JNZf6mliK2T9JugKOKpQOSxD0/dFo2KaZu4bR/qj
muoSMFBtv7I2cX/Q86SEsqGoDU4L4VWoooA7KeO5Ouat9ctGY4pSqZ6Om6KZ
iKrkXN8pAaBJbV2wt/yV4iU3PpSLKYhNsbxIax8qBojCV4vaaig7964EyFRY
WLvHO4VJhAHuMzmgWlOlwYOtaug6qg/39AhIlCo72KqCLsjYTGC5CXpR2nXp
x4ZxPQLACFMzuLNquIooR7zZUJq6x3rmIh4VLg6AeD2e+/LdECWfJ1aK5VMM
dEQ6uNbUxj4/dTdwpgIbBYiNUuHPvK/WtDD01jN/uue/wrAGGpv+QAgvg8lP
rq4ZO5KdgeWKZHYp3879Qh8lFu3GcRYMoqpOYS2bexjc9SRqMm/mOo1zTR+X
MzDk3O0Jl5KdXgShOaYkVOB78spbbi+No+o2JZTk4Efw1iWRTd6fTtuZS+HK
+AFnasaIH7UABHc/Vw2sa12Y8gFN82sxwGw9/Kp1XC5Vq3ogXs4Olc6y5vV/
/WT18Zuam4pbTrBx3GE3Wn/LLabJjItNADg98RMm9nRJNoFlBeMGYOIFcW75
xilLsdDigfBpdETIyo1u/uYjSYXKJZyVR69wfhgub+75Vrsomr4qsnbU5JyC
/5bu13m3NPCgQMA1ptJACjALR3DpomNth5DnVhN5uxQWbTI+TpGLkPwfzwhL
5Je2j0/7N/ujleZmNWuXy0vuQzqPyYfXtcX7J5zXR41vNi32xzwUGFjHZZVb
3VfgQbRv9Zl8bpWD/7Y3SW7FVikQ0NeLE+LiSxIT//Splu2GofG6aqb+xw/s
0nt4Fqm9C73b/xtx2OwBlaVE9y4bQuxSZQ9W2sLjVTkvesSFXgbDMZBtZAWg
Oj9hzufoRl8GJnT0Ym8CKrmVCxnlHqiMDVyRvBSa7fp/QVuqfZWaU0HoP9Wc
69EE6sQoy8IsGXwcIjO8b0Mdi5Z4Ay243Xw4QeF7Shf5+7h5CDFYJ5juLqWJ
EhtP4py2cXoVR6Q0shE6EnzAO37a36qWsubZYbhj0hcuakbcU0F2Q2esNxAq
/PWwWLKugehJ8uqJnYfKAAHvL0pYjEOhhy+HjoKXjXZFJy+p0qGRbL0yIyU8
w3GJlyE0363kV1IId0GDx8TdhPQjZZMwWwDXJZH6ZgymDbDFeqi/2K0sfUwr
HjldI+Aa8y1n385Y2FRRmlRJkkNsoaS4zb20S7mYVG9UKODMoaSdDw+43pU+
Kth5+Xgo+fqQi0sVcTxFKu46dNAOctYE4P2zyi4yJEm4uEyGzM/h6Viiz8hz
mi3QFHV+kv9jZEvcGOWV+BXFP5ICNVILjzJLQalGO3cxKquimJvvyDR4Rw8u
YUMgZJRQtUnk3rPZuA6c3WwRvWJymryWcpey59mgXnx+v+eelMgGOhVVbtOS
jWJNSPG7i9pahvsXgmPPLTwhlLr+8oTPgfV+wF7lY3CdMgCFmcr8RwSAZmVv
7NFwc7oKlVrYq4Rtm3Krx98jMN9ndYp/vFcY0Scx7QmzuhPeThAu9qHIEr6O
ZIVj+A8gl3+0iopE3V6HKG2JuKipjuVdPcydQygAzWV4zsEuHnBjTjEX8qlm
fDrpc5YVB6STOKorkIr8RELIv7+lTDUek0Eu+srZMi6gGaT4qPOZRCyeXttA
d1htNJBC29W9WFXD+CqJLIlhoKz0lfIE3CD9iAQakFVBA5La+8a1nt/3PoIC
Dpu9+/6hkdt81DZT9JS/R510b4He0+QNwlOhdZJdXtCofbL90VEC+gqWrqrG
YGzVV4QUHx3AJ4OceC57ZVNFIPojLp7mydQRRt+YoiHIREBieJ0+Vyi5I/xx
eZgFOi/EH9I9k28gsiByh4hu/WxpWzvldEBRabBWPw21/JTrkgArmQfakvHt
2ILi0lAxGJasw+fTBPc18AvPC8yqgo7NAkv8Cb63XdI7McceU7HwQKsGMzx7
7IiDKVVjdfEInI0K9t4lXFiCCeIEZNdfPuJ3D3sO2ftfxd7LyxLc6ro+zNcB
IvkAhgvvuNcwT7w4v5cgfR2Ve6EjPoeSitNkrWkQ5Zn38BJq9kwbv+5B6pbd
lo6Rtu3ndVNLKKA5ApZPfQPYgYNMFzhDbDqr1VBpNvwSmldq/R5rqJyIgyRy
mythGE9RHbElXsTeok5M7TpT4NdAUNh7Vo9+o3vdKTxXB7jOiWQ0scJsnTJ6
wc05p7kBDwAGf8u4DckPd7Re1Em6FaymPySAd9DDtS0Rr8GSBHc4W5HwDvvJ
Qilq4pzIHL1Kx9C8o+wtiQJuXW5o2aDxMjb4q+gR5iOj4oM+EsNjhLl33q3R
pzLsrVDesk1JYiY0MmXC1o2rJdJLWdAypNnCTf95EKfwqWLjPXXLOsNqhyKx
kEJ41zcJGIFWei5sK1ogGnpLql98su3K2s0XNJSYeGU9cZ0tFy08hEiTmnq4
OEEXWvHF0LINt50raIbLiIqb2ESUiZxJOcnzpx6AEaRmcFZ5uvQqZ+Kt+6zu
Ro8tm5X4+voG+pbmT2tAA0yA/qGoY9euVmRxjIcG1hAS7z0UV+BKgKAG47z+
2al4NN29v46ScyS8RqttUT9HbyqFGAEop/7zWJWWyMuOQBZp+yvSVMYSS/ZD
BExn+86/kCVu4R3CAQTYiBdjm0XZtj7iTdz0ut3LMUOU5oa/tif28mx0K2Vu
duA8gU4+0YdLkyZ8u+XyGGXT5vbgQD8nns/vKjxHFH4ftQDsVAroCt3zruhA
u3qUawPhxxNzB/rPHGmOKTN3MKB+bKVKrDZlvPeMmC6bWiB34Ub/kqLpcuDK
ZyyGyPJah3b0jEkQg+vAmiWqFJiWWjKGlGW9sWqEBOELzIw1inLA3FhCmJk4
Ckp4jETaPXuFMcCQZRtTPl9GEcDiX3qO8y9j00DrZ59OD3mS/meQv21/Bmtf
E6nZjqvbOUwwHVSNXiMIA8AxCn4eF+LMLynWI1Z+JHfHyKdBJHMeoqLQzf2i
3nOYCIpop2uYYTcC0OWLJl9keBY3VbtNO6Kyn6m2fF0FuF3O4EkRtYXp3OBC
8c5ME4qt0EOFi3yuocYePJKqEWJGHcvahfCUyGRDFOZw/Bh2sLjQzGxIPRZH
9FVpZ+wAKpOjAF1GYPX1gHwr6qBY1Zkf7urxRX9V6eJe24CKDwwJxAXGwbmT
jaWPk9RtfHUu+IaXVLTjNkd1Z+r7n+sIyQRjwC10PQ+DAz6sF+xOW6xunTgF
ez1H2yI0oIOZzheCLzvFGJiyupaUL51QdpT52J64ivs50WQ641I7rxMUlssL
dU7BuFzpw37KO5rBKSxTyTEFL6aGNWQY+EchUfKsWfCajWGTqe5fAgWydwSq
Vmb/FVNlDKQ2d1rLEzt5hC043dEFx7p23xESvDSWu/HTQpPdT4IZY6lSJRUB
BDSl58Ng8HL6i6YgyYBbcF/6qSlObWKLUgWd8a4154IGOJxtMeSAS6C5zSM3
9xB1bHJtakXUJCm1f45iEEzfCAWndsUh2EgsPQNHwOOgG8C8kVwBSf6n2KaN
R4GNOuRajh5+/LqIfafRotJPvYNmuACjaLuxaR6JmUK5jbuuO5oDGyZKucpP
/mWnQDtFpzLhmbXkkZlqbE8DBdlsxQ/vmQDx8uYJp+yCaXeC9rVvZ5VzN61Z
2CzPnvGChcIJlShQQd24ohy8GRNgSfhQBHTFSERKWeQm5s3dz+8JaJRw366/
21eeM5+7fQy8gjrVzNEJSpdiPLYbCIqW0A6/Qsu+oln40CDS2d35nONa/6Sq
7QdIeC/qVMf+ra880Hiikl4gEIHKBXE7QsIEWqZ1OSAMmg9WQ/M61WNVpNY5
PPzqA/2alcSlNdGGvLnMAl43JEHxv+xblnJFwGDuxPvxb6+CcJ17EHEPlSAa
keOJBjzYMMc7984T2bhoE10rzLrmPf2jr6cBsie6Jg0VQkq6eOjnDd9RHOFS
EI9qXlSMYnL7b3Q6WZNwhXmWVGGT7oFPA5dSpiMPbTQ9n2xH259THrxNJelZ
7GiSw9RgMIGqWuSn3Zmn0lJA7g+nQZNmQt+3xc/JCCuZfkxWmyJLdXdIAzaX
TaN7CAf7Na/k0KReOdBaoiGv+pNmlgW6D/Vvn1e7MpkGwJN3ukpNU/Zn5CnU
KhtVkS1uRCl/nDYNhbpMXiXNhaPxFrT/mL5V3CdaAYH2C5dlmQHeTY0qynFi
V9XDDirizhCXWFKfqe0MTGupEvi2UV5cQqRbIAXZIsdnHKbg20caFppBoewk
T3p0U127ibWqc1RaTXLCa79nqi0Rw/hhCItpKvjpCRSPrWQgwqpMRM3UV8S9
wPM182XZMIf+NPF3bCD0ROKpbtRjtWQ/bZIv/O+gBVcz6hunM2N8DuqdHVHZ
WJ55wFRgFde7HuOwdSRCKUZNy74KkxUHupA9oeCAjpV5vWbCobDPkqfMIntt
999yRVPj6e154hMs0jiBmZjTUcLctuml7JTqGuSVACmvc46aXHBgLH2+0QUU
2O4vcyPH6tzl6ceWbUcQ2O8F6VNJ1YPiXqZUa0/6El1zI/RbtJ1n3MDLnFsn
dSHH6jF2ihJV/TaPGfae/kfEoIB1j6Hv4gxDPTPJwrzA7LdgEMyThVxnPepW
nkvKTW/pUiyyhXPEzXMBeUocqp1jUav9CO1cq4IOrEGEzAjdMi4ozIMhaoH8
DLwOYi6ZJJOW2Jg1Bj2wirItsAMu9e0TyoKgapJ94Wh6AIDQvef3zoNoemZ7
A+c5MFa8ErhUXpMXLiEVBGHgmI2YktWog8JAqR0xctByChfkjfPf1SJBwaze
iZ7d3Jp2bKxw8xveccqyeWYi4VqjxxA6HT9ZEGFAbsUwLHvS1arYSIrxuTRN
ci5ADCkNarY2k/M59me1I1NxzNrDo/B6kUhER8oFTLtXVDhC7UlM2I4P8weY
IdxBRnTQbLvXihbZvpNNiqA8Mf2yKT4mJjOVXmkY58nFfWLvBn5Kwp2UFcQ8
3c1FDJaU1VLc/MGCy/VOBwtgiHlC/rxPV7BqSvAzUiVr7Zo3ucgEKcJodpZi
Nrmtm8TB7NM7faRK9KQNBmOEVBjvMuBQxZwL4O3uIOk3S/6KP7CI0n77ucgA
ucxmgJq4U+lClXDkSqAssr662gHj0rU75M4X11dyposPYRB2J5Q7EKu6VM7G
2ba8tUrqhyOIiREk8W/wNIGHu1pUneLxG/cL7ltNcBJ0UV8jL8c2u1mTPM46
kYQYv7kMY0aIE+AxbH609qeDocoDAn1uySQEplBXhAT8soIhKsR5L3xsS3eS
va+sEqtNFpeBKZE4R13Naxw3sVXsgoPQLs5hWlBJqVj3XvrsobpXHFUp70SH
3uOrHUAVO9ZOx70zKlkSOZvmZ/uYJfqooGys+0OYJdNv3XQ5LgJrsdlO4MNi
HO8b6mCRPlygsLKS1xkIhtuAeC2GObxV70x/ldYkEOLnT3xxD6uwC/Uy6PQS
sI/JoNLDcUwZWbeqVaUS6pZx0xl3NSA4kLb3Qtt50VnrNhCGj4I62BCgewLh
8mi2XkSAU8GhWTDx1eGjYvZyU34uVArJI7Hq/zQEYIOHkOy3sPikKZCpWJda
HG8OOtpuNaPRx/FONSZLRsFN73MXwYLqUqM5OukA0l2Ve5GotDydfNHopbcj
DSJ+tiQPPCdBp2FQ7WAaoe3H4jA4ZJ4vTF2HSRuOEifrMizqPZ24RgsMpN0R
pFQtiprcK5IuJkCN6h7u4qC0WK1OqNQZ06Xar5TFnf8KhL3nbsYmtWBEAha1
Yo7x+Po/Taosb02hUO4VMfwrH5dh7biodNB+ne2ATf4bYJWFdQLc03MEBPtU
pSBd9oCTWEisnIa3zszxyA021PAKMX1tF5Htf8Kjx9wWcQi/aiAxRDsf7HH0
GKp/YmoanjCERr8cps+887d5yrrWLfP5EnAT78pUvyGyUUZ+2o1QAzEqW528
/bK0d0+xOQEwTV1bSf7MACiGsjuJN9CEKXzzr/6MSCoCR/D+Rh2hhlyDhyPf
p+e00hVNHmqxS5bq05XZeX7ND3ak9M2TdlYBmxzoMCJCW5EUxaIfc+qQqOh8
9aPHVLMfZ7l5uGt5sVIoSh838nuoRA/LjML3ZBbjR6IQhQDxfMquobPXGClO
EDI3kHo/Uvuor4kSaLHSgQ0XwaNmls8PSW4/TK1kHbKGOd54/p2GIOfza91u
OhNQvMTZu0eKDZ8Tb9fsg6W3WYUX/hxtsjgyeygmONFndK0T7pu6hdmRM9Wn
GkvfYA3VtRdmI7wsBOFoYQt/W9sXWr0LnwbgP1SWS9CbQNYeIiwRuNPZEueL
OEVg3pCG98CHDW37BK1xUlsVRbQRBylpa87cW/yX+YzIGg2CzQ35M3SXlyGq
d03hRedpOzjkNLXg+DLiUnZ1wmxEJpBgR6Q3IelvY6ZqjgA+dIA8euyEuqDJ
tp57jDSwQBID44rw4yIVGVXsSTwylyjAuJv1ah1qBDmoP0Vnm1b3dsRvCuo5
gncee7rfDbwu4ohQOm1O8M9zdjb9HfFKk5CfByYCj8piq0gQRsFDUIlnn+dI
J+50EW316ZzPD0WVz0VKgjfHHPMiXpvYnFWEnjXT3OUh7dpcMxbjAWFndagd
J1mVOOLchEPmckFx7NZcnM6D3Ee0kIRji4uso8C2MdcCfNPAHb95CX0+9VYp
w7l12S8aMgGuklrn9KBWE1Gac3tRQ7Al/G3udBweVbeQam2/PLfGCYYolAb7
nCJ4UGuBHa48XDyNEr2yMoGxiAzYXC6dxMfrK3ULHv4S4b+KrCFYZCRlwioY
gP2oncXusPWT/DFUEk5JxBk8scG5bNliYNlvn3U8hLexFL8ie8V/bqnSGR0z
0ZPyOaFoK+17pm+jim13bR+RCd+cmM1Tt94nm573ebEqNlGHMneomEjzfwur
SGkFk4nz5WrFKkXiBi25T5YR0Xyxa561uUERiOoIVtGQn4TImzHPy/XWz6Iy
DsD/8I7ZJGOj+ICaCLd9guB5CcI24CUm51X3vKNBs2iBoEnACc/0Cg5uQULW
xxEfL03oP5keWXDRSFYS/lakxFeP1htx2ZhpQUV5nRIUL7qsN5EmXuPXdkuQ
OGqPEw5xuhNp9psyY62j1Imi09OkCt4Pwt2UqFqCL5q10YmKNvKOt/fZJvTl
jN3+3tqJy/K72YJml4wu3CiaMWDvLUaOVINZJSpk4xvPJYtGRWpoxE8r7Mpx
qlRHaNRN2rtKSsN6X2M3FO7kcXddasVDQnm3rx28iku3TPNUYO6VeNf56Is9
ZNaEzpu8kmlZCTY1pdgYHqT+CWOX1dA5M3eYvxMEWxJstSQ6LmYAIdHBfH0P
Q1gYWlhqSfZuKsG8KlS9HnC79yDxOKYXrot10CNqTxCSLOZI8hBkTIf2fCuI
Qkesjt7lwlp+QCPge7XaknWAAbq0Lt5lRMUOPAHbowcj1RWtNGEWuCKPbCnW
Ig0zflqsZ5eXRaAxf5aZbiXbPoNhO49IoGkgbCRiBx1qTQwZMRNjUy7Zbeth
cPAm2l4LqZu0236Ok/pvaReJxIyzzwntgXeBfJ7p5qLS0XYg7gvWnq1MeGI7
7GAzSXH0OCp7AnEu+nXhwR+afFB2z905+y7Y8UmtX3BqGeB6sbqLwqRW05wm
i7NiMiPr40m2l1VfbwwFiyDs9Bxe6A59/RElvhmGajIekH/Z3wA71zx7SfUQ
zEh2XmvjupuVXc1xZWLf3EbdEEFBxZLWsrtJnX3z5Ul/Ly8/aF6MCmtbOgJY
Y6KH2zYc/NStyY50NsJh4SsMgRu3eDJ0oyxndtDU09G4MF872pU5YK0bWrvC
PBTpxL2mrE1VAUcgFfwJHotYGckFFNpWlqUKm+ZIBNveDCRuEpnjHyRo/2rW
WNaAlYZEFq+qyQZg+oun3W+70ugLrxpDpqgwcOmhGXJ2iDf2VO2hF0/4d77v
ODLOaecMCjXq8N0yNIbE7NNvpEjepaEya9PWQOrJtoGoPDMEhrB/t4AnS7Qm
7iZ94a8jV1GcfxOBtINkTNOco+QX79g30uRX8RlUewlJSxTUfIB2kKVspli5
orllMpuyUxULCzxmZgubs2T2gKFQxuRNvqTH0YXjpiU8UfUJSswKbLq/Gbi2
hGUs/c4oUOA8Xhihbk/q0teSV+HkHUKD40KL+4/NhtjK5hd2FJcf74sUKK6q
cOKPQ/6SUCeBGnVJ/Jqlv9/NlYaDrnZPMNFlRocYtuBHHaKfkahD7nMPfqXY
B8Z7zERxXLWT98aVAdemKjtNcb4e9Sb5umeCdlymLDaOI5hQts1bymya0/ah
Qc+hZuIdDtlHpRtB368Hzo6la7rU20UaYXKp1eem1UD+VEuuONeLIJc7rES2
Krf8klr+Bd34IXufw6W0SGZRWJ7IXGsOpRH+sH1PpiyOqpehWWBoaBuqEPoX
a1unXWsD+eXyeiSkKQW6EZeewu4/oEG1gcgoLQmCaExZd6AMJUaHzk7f/kZD
q+Gptfop326WIYDUHZ2AqB1nPlpcQgc4tRYXD/TibsiAOeofC6PfH1KwsSjx
jX8W8nJpfEwf2B1Nx2xXof0IxBaDdAptIzqRkKI0ITd8bqh4k6Meng7A6QTQ
J+9qlSLzJ85mdGe7SFlaqjAhW2DrdPe/dt+my3jIa8HXy90UMPd8eNeksFqP
BmZGpDDlx598v/JqFBtWJetq6lnPzmUrCROm6iH7farLx+EcKEdZxRqUpTSr
LKVfDXJ55O+/n8Opv7MnCjhHV0yvUfbKa2GG8BSeJa+iGdII+QvMorqgvmDy
7fbAfdwLV0qyLi3v8uWzyNa6X/lGQ7ARuB1g79oziIHT1JiCyE9OegBcl2x1
U4vySZPwZ9Ian2j8YrvlGhR1WxH4RMewv4bIUtd8nd7uedsWRp9KPKiQD4Yh
HMJ9pESGmLkIGxsQrgeY711DIJQcCfzaLCyj75BeVC8JBeW1pjeWOGRXJjUm
hGhDRZ3b7Yo9vVxhgUQQclXFxSWBfPIDyMKCIUqekpMHpXt3bSSlUxFANsq7
J1+KF3kQdYInFtSVpyR6kdPZfmt6VUKAa95lYEZnFoVkuKQTJJachrOPpwRq
98N7eGUNAWIpgco68urCwAJ8hvY/y70Nut/bXcFWYAR7l7papK4icDTxpMT/
Qs/WoB1mg5tZt4YZP9QV/IlC4ezpUK+gDznP3hAvjOqm7yz8YmC4f8vi7o0o
ksB/pyyRBbIKSm/GoVGV1lw2DaUzGoR9zxzj3y9kyg6mRkekJ8AAT/CeGmB+
RxhObkRtSVvCpEXSWhHQ6xQtSTbH8+0m2dI8xzvVXX/SzbBlxWSCkO0TrOUx
XfRDqMtoMi+dSJBrXZbNRhEIKH8CCKMLRmFBsKfBuZHHcdEUxEnAOM95J1Yk
dEo/Dyws0c648CxS46jApy7YRnnyffhBxBe+MVelPKUp0O0nIjPleyy0p7KO
OkVxXtNqu8eJFq4EspUb5Mr9gL12hiYjYhqd5rW3PHbdB+F9RsmL+zZeK5hx
qZ5+gd/2vIt+Kr14SNh7q6KDkF95to8c/drf3TV0pmuoMbfJdi8olzX72m+J
kn+sVJ/m2vX9Grq6nc68FKXMKwnVOrz0yAFkm/wHsFuH1yB24bc/YM+QzLP6
lfUKdczQER2GHnFpDjSiaMMl44VBfXSyy0ow4dXtbOecLnXSgH2a7gay1vAI
ZfLKxuCF4oMi6BfzyYe2D1xIke9+N6aeX+cDWq+uWEuMf/zQW87sk1WGQHLK
0RcmDrtNEj97xXtOYyXmGwZM5/GE9A5Hc+5LgHMtDGbeFNX7lo/ztRZDalXW
yWqb2Rxo1wgemNIIBL9BwxyYUcrwd4p/0xokkEXo3KSTRGWUYLTJiBNUtMeH
+y+NNy1WNegWahQ3fbOShXY7Gl2dipqigqkKyBtfX+VzGRuQscml3pzp7L98
KRUKU8SZTvhG1ck8PSaPDovF6IHX0Cw3Rx/bYlYwXWgh3oPcFm1E7imtiPUP
Miae/8iacit2MaqrcKakIxXl70Rr1YfOOsmySIvrrFnDbXwb7GSTXwTvxb/x
F4QB166AwzWTjE61nGkU0hJB6FuqnQ2f9EQMKjLl+MmJb4RIvvGuCyj0/lo3
/tZVaaMsLpjRYGbWG01ti0RixHuOu4LtJlKpbFssei7ftcTpN+o+HCwzR/53
H/BPYnGlO5MUQi85NbKiUmmU4p2vmwHsv1qWxEJ/n64QRBO2HO3ETvFdhjgW
fy43svvPy1s01NWQfu9AP/v+/d8+GVgpY/uk5/QQzimx9shfcA2WZS8xt2C1
G9HKX2vifQY+ROPhaaugPBzKdTtwVdoRSl2/GqIVGjVGWl7h/WzFDK1T+66C
63DS7L2B5vNlIE0LL4f1Lm7iqn0idB8YFfNfAqgiXmb6mOc+L7dtvjMnfFay
+oNYIiVhjD/cljY/RQnmuMeruOUZLKT+uqFwKxCoYhKoQ9VVrxWTt2HeXD83
hoePb3RE8lqu6vmruNuQkNdyS3/gDwgAOnlWULQ0+EskUD7pk0pAQkF5P34y
lI6B3YclbPB92szA/fqugedfNdN77z5xDo651GlvWUpwooFFvBDb48nZuiv4
iXc+EzrrVCE1VI/DAp7KSM4zbgYgCkf6C+yUo98Wg9/kJ25g7+P21ZjOBUk/
yIiorlPRiIqYs3hz1V/Oo/6myvKeUaEpINyYhY3wVqyIJ2u4FW+vHumWVopV
AzxLRylvqfRPLkKfapXAUVbTkJkfTuxNC00OlEh11pP+K930jOHNEK3YZ89W
O9iBUCpQ0cMPswNUgCSFwobktnA9PM0Q/CPhcluA1oqrZ5zYtM2wPfVvbK33
E8tVJkJC8ctEtqmX22epmrVqKmujiN9baLRyHxPfy3JuHwM6p4KDAlijl1c+
ipuPb3DIz8IlECCvyN01zfvmcX3psxkeLnbheOFyOyfALsLgVz/en+2c1c26
PyscR0ouMjCzI26ellHJyeiEsPLZT1sDEhkd65ImFzTHB82x6ZA8x2d+JAb7
iFYEqYLZ9eqM3XWiXbmwD11/GtkFjJahJJEC3VZqY7rVkCQeZPC31TOditCM
9AYvXZfV78VbLSSo55UKnDgSNMAibNYfy7Z2aCRPUQ5+1I+/3nXSA7HikIRE
tcdUIO+cgLcg8wMRgWIqkfSxuu6Ylk/mQwGTi+sXwUNRVCpj6IvU+qiiphjX
DZ6q4YW/L8NMFB7xiPjpr6j07OMt60ItrokI21E3CcQk9fW2mjWaF1kPUJ+U
Nhf22htWFy0lYyxXU1301WmCy8O5e49gRhAqCgyfDS2p6IXSnht0kyA6zNqA
pReOFebxm4BdSbXZEwaVEI+n6YbkV2rkxdiecKbse/HsOPkicpSJQkMk611c
333C0yY/CaiZwaDo9czhwu7g1H1ZII1dT1dlQvi1Vn/RwkFQEY7fTD0u2Lmz
slB9W1cm1J7j8VL3HoYdWWnyF1QzyhdOY18siuYUXWcjl5EQXeX4d3ivPb0t
YYvmB3XY8NqKp/8Ym12nH0xDfotxhTl7dwX/vS1tuhocbbPV8/tPjn3EAsIw
U+yNqPKPQ4KWEYHTv59bE3eRfV7uRh55v0XgUJz3f9gTNoki0pCBgNnYw1Gy
+Df/gKUYzS50wqMRHK2p3atr/5ooHhxYqsKcXZSnFhDxV6iEB24/9FL67cnv
7vAVUDso1iL90q6wbIxTPvCJfIMsStqRlvEXpukLsdAlTaBdR9Z7LJE3hjsc
LfnCIAtJbvavONk4Z20horjavk9y0nhZOLbFzxzOA9Io8z/ifuSHfzapNSjP
7EKeMXCNTPVZkOeo8JO9mHVGuXRLuwoFBn2XwBoezknjU6zUmaHtKRwQ6/Pp
EXbT56uPh8Of/e13gMq2GIawzsxym+2eOGlFwy/TyduhnGuwofRpJfybC9eB
LhznLKMXEsehQomh1ttlIccR28mXoMd9ZDFg1oUyrdY3nsKHVFtf5WGTAlVo
VvMkHLKMzydu/mA/H5kblaIPJSDhH+s6+mIYS34fXYwIN0i2iV40TkfvvyY0
CHnjq4A/n1wlyvko99eV/CCYn1dPJbSh9DHMNCKsCIRr2LEcDreNOcrlDoK0
mLkCH4RraAgrCZU0yXB+9kGufZRWi8elIdUCfDdiRlst8kKHq/Ke330z9AlA
cxnlxRt2fLaI/0d8D3IscT5GCToGG7n6mFs2kssSMAPmvCEW5DBruQAIbyFY
x0hcMv0bN+pBYp+JeB3TO/b+B5XBMoPmaTFNrUcW8cyC4cLvWBZdU7C1C9Vg
c9zSjnRJb2msgbTAn7yBRXKWy69C4uUNYGb4z7VT8EU9wxcrk2QciUG4MN95
ssq/joL8oxUBeV8C4+MNyrRL/KB6WrznjR6qamsHmOnL6udh/WUmkRPzYxSc
fuJS5GgvXA8zxqn5+qSpBkgifEJoCyos7tnOD44iHbxUo4JjT31/osamOvTx
z6C5KaAnLHN2NRdJgP1NimGWM+3RH4ZLgBrHjy9IDa7dFPVrDSbawAzStjcv
x9H9mP+xQW8lIv1vgKPdnpNCB8jri/AKKZ0ooxkarBpR5sGHysAtxIR55cVj
Gm1BU7OAzmJ28WDKEFIkp8p/uv5TyG4BKLdALV1yIL1GlSfFY+5gGN/nnRUJ
aDLSRJdUffGJkwD0kcLEy/wOi4kMaSWcuts5mHcVRYh09fU2diATcIX6tTGM
Y2AGAYaHPCvTpK5vSKWlgP8qeE3oAyTBaqUlpaQoVItnL7wGsF/64F5XptyG
6YpTyxSd4NRUvo+RlLPHx4jFg0w3/DbTE0eD/0gTNynImu15ut1YD6OtYFCs
fEoZv2sDB4Tqukypk2tYvt9bamu2vdka6oFeMXgCk3tvwl0MBg5lH5e//vHW
bSEcU15A+8GtRuF7tWRdFDw83y7b0q1wZ2a3W2GS86KH/C216zTAPrF5uJHp
Irp5HL70y7KWfF87n/M6afGDmqecc8Xqo0KWoUsJc1ULzuNbLCxUPz+x6o7l
P+zFLHfQYcjT+Tuu273d5hg1XshNY+j1KTm+4FymjUc3oT+Vhx5jF5JWv8IS
KW1FKa4jvEiHyBu7Ha1GfQ0etoCWEiplkuETtNpzXpEwwaRTqfHtemFmDvbl
C7Z4ElgCrHrunW/kcuFI651UxpG1vdDa73I74dY1/jNllxgwq5mdMttdDoaO
wgj3bXWKukYCuSTkmXpLNMmNMLEu97+WJhwGXs+NgsZBXdPldikg1eAfnJR9
iorfssYlnQJNR2VCmkm7mxkGhO2pMMic6em7i36lsFDHhSlgxQSrxQwpRBZs
Tn+43/NUzOE/NjmZAxq7eLo/W6llfBQMDXutojD+S/+8UHf66ip6+e2ZrsYP
QInupXerX5zdgXLv3RrwRyTZC4HeYhh2SYv/wi96sMzHGalPaW+umGQ6tVKH
Qyj4H26rZs9XR5HAdZv3QGfUo1dZzqC5WDgFBXBlz2G8Qb7No3laQOlHryBb
4LqcN0QHtVc12TYycoAMk7vb+VXtCZgdxtIjurK6efobqpQaTxY2CRRhf4BU
tSWRk5RIVz9E+wh/b7i8MgaNBf6MpuupwXbLqAAPr66ANYtIsYBOMJFdpa/F
nd7LNlTqmuMt+MZcZV8Gmv41/5p6IVc2dOXhsScTeJ0TbCyb8aZ265b9k2Kd
5/T8N+ZP3VTBSm5DY+L36m4EWx1CZUfA/xwgnpBNuDcqLdIPe/zF+HgwSSv3
IpNj7U7CLdsW0fuallV7d49AaWvn9SnyKbXVp4Aiy/Cd29VkJiRlMN3yFjsA
kJ+pbxC8j3X6CYS/fMPXVg2TQX7jKrrbv4UA3Xm/JEFDHswC69F6WLwTniPv
ZgJi1UZ8oglsAzBdYnTrQ7KZga+NR5A/vtphJFR6oaMP2Af03FzZzvB9EKtD
wz9intw2mdFWj/7I903DFaA41KyQ+3U1XXaC9mB8SIvhSaT3j7DZLnF821sQ
THnYBeAoBMQXctGw9jjh17dt+HX0wKt7K/8p1ONTimac52Z8wvg1Tvxtc6Sf
whq6s5shJqylBxP2uZhN/3Cf8JQ1YtML9Co2v1c6LGg99TLs9vthulfw5Zh2
oGUORgC9dKf9kLZ8Jb9I9haAIC4+BSF1bdV4/emsXcOQT56QEtIpkBzGvb+5
C7fLzFRLsj4Ad80Ln/o940UtCxCKiHwbzEZde7BFMwcqUgyHQsGzG5RTR/u0
GXE67vFgp820MrZipuyRX0FcArfRSo3tvMHQ1zGjkeq/vgmd7Jvsmtx1iCIz
6sZOVU9o2Zhvrf9Kbvu/MxV1g1NXPqcTiXNDNCywt4dupZXdW17YSpugd6RE
+DlxOA25wRLZgc4XdnmHkycS/Wh0HQ852DowpYmrH58XmztZdnMsXnwkPYZ0
uyOLAsB1GmiqUHSMTtBke1vRo3na/6FvZM1cKc9R3fzyuVyE8ha5GGj66ekv
0CQJ/Se7+9eJ3TODWP3SPeSK4AKC90Q3+1fcOo/NV/BDIb2AsbWFcGYtRAPg
Qt4RkrpzOVk+O+uhq3WMqVDAfFsipCP59mdcbW7twvePqwG3OtHA8YoS8MQv
JuAkEwDYpnvQ68ggWPlPCCI/4MqreJP2KltkoW7gmKJ2KZ5lY+q7eu8Fyi9I
1QZf60CU0sxY7TMlbX6UmCJ8cfgRmhiWRopCblvWsHxCVmYCRiWLmprpC/Rz
PgxHkfkjTQa6CHRU9sTkcAAkxNQtGz5VT3XUgPOnHEzZV3hn+k3IqSSJNGkH
2VjRZfHR7A2cratW91jPB/wc/9xHI9Spb8Iqe+U0u/dX1zvhxPfoeYxacsSz
z/iCAQgVRG+irqldycvV521VJL1I56I3ADUw04Ku5Bw1gLgt+VmB8DbHvR25
sOoLayqlL4gl0xrcjLJ2AqkpP27OBBtKI1AtrdOZqv8WBEEMnciZM4vjsI8D
SG2YE/7smJj66GyUltAS+jNK4gdCUCwryfJ2+eohCJgbJeZV66lx6lCmwKsm
9LKNluPO2pi8L+OcHaaCF0FCeeKDEyO/5HD8TnZkGZoT1zaKoZSZYlqd6zMM
ohERdtUaykKoO5HQM+hX1W6su53ad+qJPmhenpjr++k/lli+JaSGmzJZWQkx
JTKvYhAhCkMJekkP3JPhaW7UlI3Y9IlUZNEbO1NneNM9o+UT6hUznL792qq9
/Qv/FsucJzeVC83S715LJqbLe2Txd8tr25tYN4ywMjh4RXTUFImyngkyToyL
yCto/F90JnanaQAcWMYmhTnKNxGDHo3cv2IQtvvStP3nvbU9GDWzuzjiZCfY
9Jlw5Cy174SxmkUs5VQHntJPJZPQOLwEawxJ9GTDTu2UDOse06VJ93zPSmq3
+70Z7us0Ue+PkaKZhJojiggraZXDnEj0nOlHLAS0FG/ZE6qT9CHLjekEBcH0
Wt2izf2S9CuCCK9kV+50/rlCckdwPttlvgc4tYLREiiB1ilmjoDv0c0ldEd6
C9Gw8DybX7sJ/bFFpFjASTE2vuHz8sYDlAjwOj2tVskM+OmmP2OWM9n6Q33X
ScZbG8hg1DtwjswJMLKXGpRvO+oNpaCpoLCEACNaKOnpxGTv+fcuuqO8LOQ9
/bPdbag0WJYkXm2dsr1zP7rWi3gSS0vSBd7+qf06lpTew1/4ZXcJMYPwpyFl
LbsA/By1vxnvUsqkjQL0YvvklHFUkOTeeJ2+7gotZ2WG1d4S2Bj9guI0s4lC
vBV0BGoG6pcXk++NJTuQxvCzagW9E/NILq+P1gUtNaF6xHIIJ6xGrN45VuTC
pEYmECl97BUFDK/UuprJdYof/kmMuvsycpQQV1QTefImcS7WdLa2ok5WRvfy
85EEo3rSYlM8Ix9ABOn+/OKanQS5XrCjH4VsP84xQGh84fWTPolrkTQNwCxu
1PnrHLIIrr6hBPuwiwbmENoeTtC6G8VXRtYNURFBg2qVsVUYKk8udQ87QR+s
9fetaVTY3UmNx62o6i3/JKiarofzlg3+aFD17r5xCuJkPAFJdDCGjHbV7M5J
12IO20pDNe2MvDOeTxKrfWZXyJ+3/VqBmdZxJyt86HR5OlcEHQXhzRajHTLe
4zGSw879VRBRS9oj53mUQNsREfz/lx13rkRckJarZdEKwAYdQR9p4cwS4WJz
2p1I+lli+m4ep5EHm8XL0qvU3hdzYcGYKh4N38Db5r5edhPAcXhvdbtS7/Os
7c3fUZ4C6kG/xvfl1E+o9jBrVSjQ28QnMztOS574DXEK0UHGb+4QQ4pE5DHK
V1yXGesSxCQ2xkugWXoEmJDhqo1Kz3yiDHaiTbNejIn2uVY9Esm16zC8icGH
lSL+fNCgYK1zAs57QYx3DyeZxeDtVZnthJpS35XnJiWLS5J1qzf6DOkFwIeY
I+GHpY1LT4ACIRrPJxpNzf56+I9xmpQcK4PBAbRhMccHZ78sxxbUk+IrwlLy
peCdsTB+AQuQHLSTrZdkKugyJthbyMnofjC4/Tt+nzDN150mr+ijHBK91061
fX2809ViM7jHsBOJ2dQDxzY5sIojqkpiG3VBZQVq4lTNnvd2fGsZ4Hdt1XIn
sbI8Jwnh4hwyB9sYxmz3ylmpxqhf0e+jK6s7SY97h2m3NUqGek2RVOtLBqyf
tEcjHOY+zGatEHHNfycUq0KBOs1izDrOxjqwH3cs2ZRW/GSQczsgqvAuNK+J
RhrXacZgZHIiFrlLCITsceKZ1Ym7QRrftVxlPSC97uiAxlxPXNJDMM9qY75Y
kcKL2wm0R16FvUkpk53plxotimIDqQSBDonry9w4G3XUsFjHQKfJ3BO8BHwt
Ya8VenSfOf9RVekg8gwHZxSAYga0Zo2oH6tNVMAeUh3iGEkOtwiQEVs8+CQl
kKqvwsX7FBcXuZwckh202h6P2CQsGI0gdFikufqckfHEOkBl1lpaiGJs8/0W
lO8REm+ZitolMw/LzUYl8rIYefvkHVJ86EoEcjsybDAy/ypHAqfgvNdWwdlJ
TTMMzdtGRdzj0SHC6Q3vAwzKWQ0oPDU8GFgkAlCCHqeCW9T3u5BrpaBWWXAN
Xy6l+wyMZ2xHCPo9DUckjUqqi5U5zaER+LwEzMHapjPStED94EuhkwbfGjFT
HH71dke1zgvOzfz7ibO8/VxQxXKhRx03tiTEWjTCMy7xU4pK80Ca9VVhDn9K
A4QL99OLPTjunqZJLBsiZC5XS/3gpHGOFQ6y54R4tZp5kCeBWLEADPHIDXun
M+92myNcK00Je7reYL++t+iRKIApW/+rOOPeV1UTokplSGlM6Oi5jY3JmpmV
69JeSYpdEnmw3FKJapbesAFiDS781i3GaQVcZfLy6LAplbFpwpzS93Y/S5Dc
CzZ7ZT+zadyy9hex5UYbUsZk9e0wmdC5K3iD2iOtNyIEQBao2f4B2RauQrcX
8Q73VjVzPYgBQr3Psc2zAvGoTGzGyBYapoH+SS/lGP5gvTtT6nZyVRELdzc0
/VNE92yyxwFME+9yXQnNfjhL7YcdUjSDkdFwzreBM+72580sJNodx+/Iw6ZT
5PUCyN3LjZ1x1jVrHrVHwrEOpVQQHCAkjlG9GMCQ4r7tTFBEhqNzaL+tEmZD
0/qxnMrcCQFtg92zkv8BDZqOKQE/MOBvipIaLpL+zH7e2NRS2X7RrsE/GQq/
uweP2ABvVIvKLtbgQz/8f/QcKWH9ozgx4KFIowpwptofEeIc/p0yOwiJguUn
7ZHo3Uit1gVhCuqMv4Jm9jNRhpcAZJjz2cECT0jXLzZLPEz14HuZeADWl+EV
wNJ0dqiaYvXbi4Ow2+kaiMTZA4Z/Znsazzj0bW/98fQtcFmHPco0n75jWtQ5
NWH8hBbyHVJL/Lrsjtyt77ufUspFmkow99xBlOOD17f2gYEFIaVLQQTjg/k0
p6C3qA6zVHCsirhYsCiMHx9ArEKVnXUgymhBa4Mv/WRAyihpOWeK+Xv8YA/6
c+5gUmfekoDLJkU16rmX55AsoLPLK/cqCPJfbylbvX/st0hh+62OEE7uxEjV
EAWy4eQject0nXuNdnsKInslyCV0BVJsmPFlUBJuv2BnYa1zhByYhX3+0RsR
aLdEHps+5LFJaCFH2ed96OyUBSn1GtAU2ppEn1RAS/wIXk+WKG3T/vvVnNCg
Pk/bxyWs7vTAX9fVTQBWrWb3xh5DOOMsHwXqhdLL+vrrz5qwi78v/9orBR1s
doxYQyPHY/NBawNPVUwD92k+KXynJfdKMfHryj06Zz5Fo7xXlM8ma9VIEd24
VwuktA1kUwo68JBBl2YQh1tZ4a48MGX5EuAAecroZmc9OcDmeZP0VAkLghjE
fUsNo6lGEh4IAOjt1Gypmx+gNqVTIXkynrqUhHJvC1bhZIAtLvzeLYgSis9t
yd+yWDXTVWJ0aJEULPoP9O0GaxmsAj9JZERXAC1Lb6o4j62+KAhAcjv6Ibbh
yhV3nF0CN6b+0/IwWfoJDd3HCBQleqBkBwQCfCWQ0gtbaVsQYp53GRTnttiB
kekM9RCo6MAmhdBuDdhI0Z6wYyjd5hDXW1umdhxgOW4g5ht2gE90bJLWODXH
+t1zS10Zkzx7+ezf6dwrWk/aqPCPeKBjio7Ta4OrUAsIJD5484+TmrYdJBpm
/+PFapJCjCEKrrw0Km19tRj5wgn7kJ50EX2t0mCO83tC34kQpcQNd0sRqAM4
zsetvgZ9XeXDjEe2zGyl3GIf1VQYB1ssmmNNVde/7dYlChefKx1xd2hoRMGz
w0RUxSjS+MpzX3cqT0tm4r98q+AoWBFAVWWgcPmyCEDgWt+ZYZ0D0uqg3d0m
VXygueoqNmFeA3+l+ERXw9aXUlJsJL1wOi/FwwEHzdp2trbbEPhvb4muX6r9
TSnot1zm9fN8XmOkgGzJlkbhEVXfRowR27ejSSACnQCiB+egIvRq4tiyNiHr
Vp5vKZgiSwnQ7Cw3Ik3cN8fQ+5xIuAhIlQ6gXT/Kd99n9ch4+MlWAQpNwFYu
GQK2mpXp6uyN7Crg7UNoaaML+E1e4+gxE4LkddavHKHvpemNUIjsWehVpe6n
jXhELS5ijW9gyNtdEz/bb9qDfSUn+Bq+YpTaOAZZymJm/2sHCvvRC1m0Ug0b
spq6zFHZko0tM7/an7sJ6m+9LNBVUBb50dg+Q4FfZwWWIZ26ExuhKWZMS/k9
l3rdvh13UVNlt3hQqK/YxZxw91FsMuyDOMAj10NFnak9RXv37iQSmnUznkgf
xpHf5IASi5nbopK+vtDkooM2Vmi0iaeXuXkisfCzvXkMpCDLoWmd4qsJF9j7
VMuTJ1oZ9pNxMxvWQgYgZWSZil9Kd21GQxCHIG4MMp4D2cv3vaQA3j5S4KxI
JeefZiG87PclQDS6aTDoIsCKiRo7RAGPM0pIfEf5+K/1QnsU31V/YAz/kBsI
HIPsv/RoFdAbxppee1DRDL8u9b7I4BmeyoGovbJwRAz/l4YJPZn3T96oJ2IT
cZR15o56qX3SaXhL5G+QXAJyHfpDanJHxahg7qb2SuzJ/fprVTfvW8D1Q1Kz
8AzriYtdOJI0vPow4uQp5f7+YU1hKZIzj9usQyH8luc8OYyQYulIsGuxjItc
GHNU8eFNTxG4zkHCGY54NVxBFZdvFuNwZv3IB270lBg0Xad16Bh4EkbYO2Fz
CQs3vCtTCgHmgN0SFP+7ls+3bvWSDHpyYh/CPoE4kVW3AjBucGk1KsznrokN
qMRggvrtakx149PEpKtdogPu52q7MV9v4gIvNJONnInHbrtk4wcjD1jSCgHy
Om+1ERsmQ6eoAEvyziJbMIGZOGOjjgRqAv6cu8eD7EQqAAZfc7Froi97sPbM
OiF7YK+8qctiplnNPtYs2oCdJXwjjt7gDwalOWvg3NsjRejzk2LfNil3T7pd
oVYSizTJ7QWlz4Mbz+SJB8RmqkLwj9XAG8ILW+4X4uUlTJkN+P0PIfyvwZph
d5uvKsupjkSKni7iOvmNYwJcjGFQ1ZNI8Iu4EXzC8TCGkLFygVMoCIBwoAWY
G/agxGRHPy35oe4B0seTPvB6IPpMHeIOBkWLWYkDcGVbz8rvnX8iTtYQArBf
ODDv9ezRqZKU4Lc7PgWwRACQdSfSbCWnH9yP40I8oyN+PPbLZpuz/2y793ZJ
dJA4dwckvPSUqvvy++Zngn4MwP1YIyAI73Fx7kggXI4znnP6xw8kHwJE+V8E
N364q99jzYxeRKDwvVColUN+JSCOHo+La12A15cwVcLEtsJV1CMU0NbVWTZV
KXA38oUz/VLYzl3Q+WHUu8FlMknRy4SC3t88gEREZEf3MxUoXBdBQpEYqDIU
DW0TNsnS2sq/cJvpP7pQi4Z58g42cYZtdctKq58I7cVyoNmRD+/r3ZxpVASV
lDObVdBpeJE4OX/+JxNSwjJBWSj6WTxU1qZZq6x2/6JhBU2Dq/C9YBc13o5m
Yi/Ra54WRr3LCrB7lxfvm6XRXk7/QS9eVzw3WuUzxKu8TIDnh7aANka2Sbm2
0RjJg+YVtWhoauQQtNV62gMJyLaJ3J11Q4NjJZMVgO9qlqJCB/ISOham+X17
5fgSyyyk2IspomX5WEMHVcPKMt9ELqrfUnKI6YxgelFuRbspH16XlwI7CUrs
kUI/pdybK3Z+zy31fCyQVTvt83AbTiOJraW791qlnE+uNJ+sLY48pjkVx7OZ
Yy6/NIl6hnqVXL34KhoTDAh3yyiDYAITx7BN9q5aT4zcDF6AmPpSDCuKaebh
a5YQesPS7Le0oOkWb2rNy1xwtCVFbT0gm1unIEnX3/CaPOcxrFVU9msINzx9
3BdgEbziEA6b7RBRqpXRgqa8iHKTF12gW4+cnbczJj11UljBRnG6o2Tr0q1c
1qm6KP7qnLpr+Bv6Tki2QkLLDpaboXniAqtlSXmlGi75uUy0vMXwZyqFkZKx
mduhY9geOqgpQW/ix29W/9mIfr9DVrixThDYwII0wLL8KC2iDYgducFZajwP
a1wRrha437BJTLrB789iBCik8g2g7B1Sf8VZVeG48hkEcf7ObXHilf1XvIJc
q7UOHUNlSEZ3nj37fNb1NIg5LBOUxwF5ejs6Q1zyEl5lIQmPRaw+g+dK2scj
J+ZClBxxfPCCA+kE2he2ytvWAbPmqVvifVGD2e6hpif/h2JAoDk52SXE+N5e
VdJiqyvtr8o0Jf6hGxQ9aGAHgbswDAgLAaE1zqY43EBTfHY8SNeeyiX4O3EV
TR9umNFbEl0JzPv6sEwHdCNAYSAsEVe9dN5ZARRCnxdZYccz+zY7VmR7SIR0
R/XIz/ToSUZOIsO/9OZl3U3Ff9Wrqw0cIQ+tiDhh96vEKaw11Q+QKG+ReGym
h7Xpkdat8zuodI5n/fdta+CXB8KY9LADP/I8KpQuNsZeUTcJDGIu/aFX0NJ4
g8QbLC3ypQ6L559Fmx9veU+gthGGMS9xMeT6G9WQmi7uGbp/Mh7Ql67nHNmI
AjdJH6HgiFQTuw7eJ2QZ3hNeNVDdOunfiwiiwOnV67PTKTn32Tkn15g3+SrX
+QqKT9BtqW9W4uOZmaSZaAO00t3Ngv3KX0lk/u4tP2duWYlkqgbh5L9XnPp/
KNv+HtbsrR8FT0wiF7WXQNGuGI8pk4YaiOnuY4AQoLrPH3gN8UeCO4KKES1m
0+gpqJeS0GbtV+gJVpJxDV+Sk0shgn0X6sVdA/hf9tBMcmu4l/EcLpquhuEI
FFUDvmYEOzJBoJeXE8rfPv+yTHggcinp3fpFg61nmN4AH+vXGrkHOaYU3QN6
Klq8timAfrhJBrwafle6YPi2y5G6p+/w4oIwg7TxAvUcKEk/a9vbSIWIYPYM
7cTMAD2nYtgzm1GnvwAzDe7y9Wl/C1Jf6/MxTQVV6pS7K6O4BjzAUTKXniiM
XpUCAzrUoDvsavsVktUKsKgLwDG+GlIXRnZYLTCCmQUz74fK2XU5ZPB3Qbsx
HuVqHt53+I1XTAa4hi5fZhLGepcHg/YeJ0yhtpTzF5zBcnPrerPw7KIMIv/u
ffoET18EuEwWlPpjFN6HQP9S1I36P9vWuhbGd+kPBEECktVm7Ou+zHZQMqlw
ke9sPE8tPkcA5ins9dwT75llRDwrMrl3Jy+Y6zjlemRy+DqxWZNGmZOaUDST
pry22Y8rUawzB5nojFPPDj0MThuUxp7CILrvE9uoJe7J2SmAfnXqyqWDjtgt
SO56UuFCNEIZhqZIbjhWsWVJOsgckah6DFQYBFbt3BL3bS+RlgbYOAp9tPtf
PpgM2v3mRJvCYYRcawm7sUvAAisnyNBwl06//NGUhd4A0Wk1ynxEwRyNC2Wo
lgsGfVxbOhlNXZLXq9bhJaZ32Kjdxk2sVhX5Ypp8oioRyllawJuETGKQam9k
j6c4r/rrh2/EEFk10Hq1lfoTLR5egDXDqaNYwbEcn0bCPjY1hLvGpzqzRnw+
3HnR/k4B8R+7NnAN8JggT4CNsdHgOf4439ZDDJNFn8JixjDsTpTGxpoC3zPn
bpTOI9J/FJrx9OQtBsCfCfS4Gf3zb3ZDsbb+XV6HLt+c2+izJ4GIKQbxXx58
Hho4D7BVB6Wb+fBfIfXhsJNt+7ffTh6sJw7Bki3o2vtr86pnRDZXamDOryLD
Vy8fx++t4RPaWBK5N5BUvs+C01YoxP9lddlHEEc64rTMdPg25uOj5mYPMIkM
xM5VG3MGEqPEjkDxbJh/aYW1RGwjHtBMQmhDZJ2wfWL2XlYKlyX1jTEzxltj
T81gqWpS5Nv5/xTm6j8TB1Chy4qQ6kQGRyuXOqNF0ecg24nNoC4HgJbh+/7r
/txz81UVKnTf3KKmuo38SqfciiWhL2jn+x22iUZ2X/iIlWKqo4ZwYXllUt+A
/tuNK7IPuZ87U9n8zcdG6/AZ1XKv0h5Tb2dkFUWVoR99UcnyLJoKy5h4Xb4I
QuqDthnaW36XqCvYfwEFA+LZNRM21tdeRRaZDHg2McchPB9ao9QkWqWt2D/i
e5syqnB/4AEpoQO9i45fpBSljeUzq1zniEEoXvVkEtAHinf1dfEtdhWBpR3D
8nOqF/2Qivq5Jrw1wMtlUMj7jVtwCjwUL3WPlf5A++22nUEwgxkxy0VS03LJ
bX1nzVD5Lfet3TqAKjyaNjYM+tqM6cqoEY2xcy+56V1nr18Wd569sW0PutkD
vv5KNpZ0spMF34gG3TvDIug3ZlOlpxYUFWQUWP8xnzFFcO4ffHk/fvm3ODyt
dVVxE2e3XuPQcCNGbeZGQmBBU8al0g7VJe/PbdaytHqmzQ+Uj81xR6gM0JiZ
33soxthCfCVGgb8hZp938eb5qQF/a8hga4QA3EhHPFkETnk++Zkwx0eKvxET
/4kW4uLALQMtoO2eYfZpxNDAIhG4X8yNdbHzhA11tfzyxmG6omf6lF62Ka/a
aR7zJ1C3K3EGr54k+NeYO9CuJDWP1KkjpSSWzhXHMNXukDBPydbHGvyAftYK
ClJKjrrnahh2HzlyD94VaFEK9cv7C+bUE+b1IE2XDd9QW2hO7yTxuism4O06
uGc+OrCEm8dDToaKCzkm/902KYX259ZF7zEk3rYeco1EwnxQzsL+8vyEIxnU
LivMf7Qw+/sA8gWnFhQP+XvShOvwr+Ur1YUBi9kUfhE4ey54uKAztSGJ6Kig
qfmxRvFD4amxbqbSGFmZ5F3SoItqx75u1k2zsbemn6OXFZkk6XNGu1PyrORG
odIJLyEQOLfSyNCm4tQXeZvbTFyT4xFg0jTDjyevw3Bttb7m9zvInefZCYl1
LntsYudNDBRI41+chDbiQobPBY5f6mbJ5GTAd+eJEVv+Bi4uTRqoENryMrnj
QZd4tys+ek1jfURJBhcMS+FikCE+HnCW3CrmOXSFm03vYYMT348vbyEIiyEj
XIVjKOinviCLvZPK3uDGaHobX3LaFth6Dg4iWhO1Nj6bXXPtn25/9invkeOP
j8MOF7ycDxkeWnzVMb11oO10koF+dNsiksN3vOK7MbdLq63K3wXmf2Pe5m0H
OSNi0WCIF9d7411+tyH7qO2o8zgJwAIChsV/7AzC+PToyaigqi9Bm5bgK1LT
0Aq56tehyKK7Fe4DAF6dxXB1nUWfWAPY9NT6tpvA1hafF35fL7RSwfUjt9Si
20TdcIjCUk8VTd0oANiT5uxganNLTy++4HTxlk52lmdAGro+p1OJ7QXCeprJ
l0NTT/xLiWUSWZ97nxDGRqi9jrCM3MgIzdHSTs402Wy8qOfAwhFN5cDCC/Hu
VlPD6Q8J0iiBva4SW3Z4cIeBJVlrJ6SK6sNUBidG5Ra+rMVcx0RoaOLeC+xQ
joeZeli+IX5GLRQHiVDTZ80R0mE7FRZL49uOwx1LpGPIj6nlPmc5v+D6NKUE
lGEGsoNhY7xbL6ye8a6eIpxw7Q0lPwhme7QFadpW7LZqtN6tdneCKcf637wt
5Gwh6AcJ+yul4+kVpEUW9ntMmdhJY63ovwJiZ9wgADCcPgw2Bx0HBTEmT/AU
9hhrZ1p94wkzPVLm4efxSB/upCoI7UsDoqQb9Uq3Z2094+yuTrt6gorW8AAj
Rh+jcdDrpCV2Dy3konDKkPqeuZ52Im/thi/cPGuRqHuhCEyVgb7PaVym/PH+
6o0dB8gNCpjO26vp7Yg5mlKCGocKsYWrQ+ppqpqucbQVjKKV1YpQ1a0N/jQR
M4Vaz8GHZy5w5ABBtXUm/E9kx4AzGveVGbH67gOzgnI23SkPFLmRMLvgCMuf
rDl6JTgnkDhx3BGyzVuBxoHTgB6zH5xz4ZfZGoApg9zU5ld9Kz8h5m7U7qsM
cQfX2oDXeet3PUCWKEYF6yGHQARQ8huP51jHJmCJLq0qKXKaglST8+eRh9G3
hlY+6z2aH04eDDBSwTk5SO1BrUzE9ppV2ID5R6D7LgdipGuVtjJeg2Wc/aVg
y8yz5qqymySyNO/4t/FiQmAFWn29PArkpimxXI7HZiCmcwgw6cgyteiIoBnK
a8NBiJ0DaNogzK0zuM8AzXsBrRgXaoVPhY3N0BmZsh0g73gA+qUH1IP4ocrz
jH6g0Jzl2JVLBC4oCxgkOueA8Ua1Q+dv0n3L4D4GegG11eDUCXyl2k8ycitQ
lGl7SA9y2Ahxp8ZFQHp+Mc2f96GOOp+7wVlIyLVmIksXeYhKuE85lVKRlt5H
1E4RKYCaD//42MrLyjDMDhdXpHoOfEGP/yVhP0yy8YVRcSdNe9rhosJwTVLA
LJehL6r29uzsAIi4GalvyYAI/zDUmwOsw/hLs4tBbiRfvifWE/EyX8nH4nuS
TQG7C64g6dnPcZ/m6YeAvnCNv3DZEy2sUpuJzd3m/ccFpeGzmvQ7BqdX/0AU
P8AFEMpZlnCkz6z2Vocg4SdRxPjLi6CmD4q6Hoetc/o5Mpo3vN2pNuCOOl8t
USdlAbaAjidM7Bylq3TztfW8aGQ/HnXGQ2uXpguw7B+5akodsMrt2btzP8iH
yrLhXjOpV/e0N7l/C69gtK0XA4iaqot7ASloucQpjoIF54h4oqBmRagnE85K
dmeUMfrrV28BlSKQGoIIi0BRJgu+SwgfStAF4YKS1OqFRXLXdgdUUIIypp54
r7HOk5khB23b3fSLQO+z3q4N7EXykqTFnDMH0h7rGwcUZyn2G+5QcE4iEhUJ
T0oZE8DBDowUKQoGBklSA4ietHAbJ3v08whNg9UXuWCSuBqHqOCN6Xpn+R3H
rpjYCNungYLfpKiwfk+aA2K/MtQFdpP7FSTgueFX7x+j5+uT5yzoJXtE4owG
Nt3AD+uqDBgN2HdnDtOa4pp7pS+SIwrZXPCSSggfRYcmMtNfQ5H3MKYtnp/s
g7VbW5ljIvn/ejd7v5ocvUhIJpSMl/KG7KTtf9Yc/2q6Tk6diAgAn8XLEjdg
Drulum1Kya34gRMkhIP6/CG6/bZRYV2Zu51cmU+gcnVLnr3Yv5LS96YICdKR
9+4WZUW6i6C8mRXNcVymjUXc5UfBMqGcjFPUCjeUpuLrafxfWI4mfL3hQzOm
Ao3o1mSw5AiWVcm2rxtDfgJHIruYzFNyKo3M+3TIHLRVAH6PUCjt7RclHq86
H0b3S1pVEOhAGglszpArpZmhL3qqETZd5sXMu0s4HfGz3j01Qu668vl9EZY/
EZ52fXH2EYIWDLJJ3kJtV/DT84Wl9YdHMb4G3bHlPBhLfeb3MNDYStJzRSHN
p9sznRXsoVaZhPMuVkwbd8GPDQ1S1IbJFzJVQN5Byfk3v7rsyVHRxfkYeHpG
OCO4fU4/RFGAUlyUS46Tgl0cB3Qcyu4b//kwF/68NTGw6jSblc9kO+TYQDtu
cbKIYWDn0FRtOGjBOYwmNieg6ydvN1lhZdoNxgrbkb7JQLqdodlzyS19RyjS
ic+QVlYWbPaoDlEFcns8fMpnhcYcj6SDCCtDQpQNY+Ujc0xMQOUn/kL2muRr
JvEbKP4e/Z8Z9C/0TdRpzrrUL3Ag+LUgBe5Mhhdcp6CrFHaBVt4JNnDEPYNg
swdLtnTuM8QKzO600XxmBecmOPAFAMD5oSNcRLx2KefviDjkuUnr2NfFskcv
02rbzdHwy9NgN5JZhfAl6+BNg9NAO6jozp4ln6mnzCxh1FSNDrOXtwNwO0FG
XBqZFBSNhNQjlpOioGx0t176kS/9itPPNQHp4XFfm+S/Aw1B67on7xvtNW6x
9dHPKjtSnJocF0hMRRr/4gPjPlJqJDj762R1zuOpxyZYwsLe9Cq5hHL3lq1P
G2PqbW8Ac5exiz8Lm5P3W0f28jXMqeOjgvMUpCPDBRuJ64e12pR9zb3IqJZ6
Kiq3k72J6F9g15g014V/WAP8ePG+xr3OIbLBGU6XSr2xL6awxxz7sUgHKkxU
KazhDVAyvJcnA/Sbg78Z+HdSh46rrUYopD+f0uCsiMw1qMGu3cKec1nFRygy
JqPVvF75lnaO9jNhtcImJZvLvzvuiTi2ulxiHSNozmdf4IFOyI8xLwyPuynT
UHcDgatY3wWpWGG9vA/qyp0HHHNyPfpF1YMbKNrbiIkn1bcnuFcAgckuWwjH
uukq4Zl/h5rTHcc27T91rl2zntkGAZ9Ib8NDAH9vu94qtmFDWfzMKjptuvSi
pkLNtqCaeixrCenKIsegASpN5RJXYnc2/fejNsr5/Z6261K9Q+z+4rQp+xM/
2f3m8liDetkIFHUq/PC4AH1617+VL5OrhxIqqFhoCrPp5uAe4rkdWgzXcadM
0kKhzDFIBUrCfj1r+sJoHD0GxK1g/Oeeas9ii24e5knHrhsdJcoFL5CiUrWk
V1jPC67oiITGknj8t+R9c5DOvvarVaPLoXtZ336RnkDacei/LQVFQE03rN1s
1vOHgKXYcqzhaLWRVEZixVmSnR2vpGorV4LKkHJU4mcTXDIhTADYOHgBUfmo
Mroprpi+WoM7FjXOXnqzC/wXB6TrIcyDGRmJRnwsBwzbomWuZj3zMg5BHahW
XBdk2Ixw8bz1wc+X4IbrKi+GrttCzqIGWDztQWkAQWoLxSIEyg65IWjbcGN5
Ubs/WffUZAn9VDPgGKuebKY0qxV4+cJGycEoiPqW+JWYRKpqHsk/PaLNrriN
VJ9ubOQVd07GSr6CwdnXIw6Qx47xekHI26WcCN7iV4zhoF8Hwg8OiFSfM1SQ
tRcDiEzA13e6m13xux6du2/Twi6jRvZewQwsGjRksPujMLHZRPo6Ie7ZK5QE
qgWmrJEmouJNAnMlmCKhDQjt08Yis2lMQ24mQh6sNMfOY0viw+mFh+MhXh7B
7S5XmSdwChkd6Kn2q0jSn/nUvkBlfhoL4Ckh995UpzS7FOTRGRtRi2n1PpvD
YpoRZDv5lDS8D8zXXanP02QlB9YGQKTOs1M9trlhUdOBdtBSPFe5DBK/nCpZ
+tNb1PXlfolLZzHrDpWiJXYS7aIwC7OGBoITuTqIjwkFdLnTXuIq4vkWiU5Z
LxSnMCvDAPbQklKfhlitaa8cqHk42VmBGCCpOh8qsCRx0oWqEvyJ472rGO11
lcCzbd4efWPZhjzk24rlN0DSbT2HoOF1SoC0U3Vpes7HivwmLLiM+0jNVuh+
Af53L1jyyT8+XHp4D29EBoGBMWJVGxeoTfinTOf5GZ2btnd8pr9XN+2OimnK
/S+66FL35vSKzzl8fH4uWR+1xYfifWBY23NaKM1q1GFZaEwVe8EL2rJWL/qj
Fl7zEsuxABYbt3zgDZUHQHNRCtINxg5lRuNyPsCJbfgoH3IG6pX04mHsseBI
/8v6MqtEe/wnlP0OV+uLid8bNdYW6V7MUtY/3VdDwU7JFzsdWj0QQXLLz2fz
l7NYDowBDw1za6KhI1rNb1RZ/42XpUnTsAqQ+UhcwCIBlK7ibZ8MxV7Xwu9t
sHnC8qvzxZomXYRrlGD/miuwl3IkMr8/r3ACoWQbndvZF9I66D7E5bm14R8D
DDrfFnlYptVgkQWwQKkxGYbVraM5cppzk1ScJjtLn8/3bNBJClgBtUE8fp9z
+DVKSTQTIwaFVC9UPgtGgo/NpcD6AFRjnSJbEu1ngZ1ft6vDpkt7fnc87FpP
PhcEidLD4b1AXGaLQ+N1wnZ6z+yNfg5weL232iNN1J5+Nvc/oQz6SNKIFC2G
uHj3i/fZqxEPJ7nzQ9CroTNhQgZi6r5rmXMfyS7lEftmxbHPrl//nGP4cXxr
dIXqZhQIwTfcvfeQdG/aEqyTjHVmbQJZd+UGdFtJ6UGuYntQHdj6EdJZDeGr
lEVK4hdfcC073PUmOjcJAy05XEjhRlj1Eb/dyRFy8LS0odZGQ5pAvQikm+kL
raxE+ou+wTykLKBPwR4mX3rSLe6fTinNsTXPtWzaHPVqE4myFfn1CyRrYBtb
ojsVRa5CJo0ZsSx5shwEIgspvqj8AC4Oe03jSmGcl3ca7HTRhKUL1CdSaEKV
tC1QP+Dlicx2TRJJWFEspp+7yTQdQt90IiCo/NSuEaGh5uD+HYOWPN2Smoej
ukbjNH6kpStciCSxd8F1Kw81nXEPlQ0Li5fD7lAseNr6paDUsYMhtn2oBK5G
m5kLuWMAG0Yao4X0+M6r3gjLtjON3APrm885odZikHLK7lAolUN/ZKA230YD
f7V6dELWj+I/BM52qYXP+S+fcaDLJu259yZy8KkHJnTMYIgdTKCp/dmn5f/C
vdt2Xulxei0PL4I0yltKJxKUwtilQi2JZN59BV1bPl4qsPzecwFL/pSQ0Ywl
AaDIaUzaP69og0n+gqSmS/u06GMOLJiun89crVrkqtU+5DqgPOzBie8HJC0S
XorvENAIkVVz7p8Y68eMXmWbOnEr/0Qvrc0AJGiFaLi1dr28thVLHiHDld6G
PJRwZDyDjmgQQ2kqpGX27uhndV4FzZoX6lgIc33wPc8ZOZJ1f+NnP7iCBsPv
i0M9OwSvn0Zpi/A6gh9NO3j321HhXw/Xf6S5OJ5G8LT+tv0zKimfvqcCbKTQ
i5VbB5oX+YhidkOWUvEy/vEKIv6NcmI92mKmlqTeI2gl6Do6KSGREEnVuDn7
dmw0A6N458pTtzPhrUcssplHpNSEdN4pdNG42n/vd4c8edkwz4BHEpbOMKFz
HdggynMTugorInRjy2932JWQmDGO4xq7Rl97v4wyX5GysdD2IgCCVyRAvVl5
ZvSxqdnvHZdUpro2s/GOpTibMiYyAsFziTVuypXtTTtKVJqtWrlkFMQ0Zdx3
cVTrnS+BD8Z/gc/rQzdrrUEFw1FogfTxQnrClTbfpug+E3A2Eguzz5YXcMkp
EE/kRli0HxwXYHewrn0b9ERCU4IQXW1kCUxtL8IJqzw458swB3aMTZmecw3Z
3HVZWg7r28vQriwqxrdKHzThhw3V4ZIts3pOOtX/m+3UAWMKo+Q/I/Hz5vWZ
7cq4JC352f6VqQ8GC4DFesvt9EIoxvyC+PJi0eATv5gJSZfYH59q+OM+3jdz
1YWoYcak+inhAPHLtPmYIRpoOYNMccjlhJpWYuyB1HjVZPZuO2E4yB8gb5xW
BNJ3TLnLkSFp4VTL8kO4N3LAI8pp/fUcb1ORZDxOjYBLdqDb+3ynLoMtk3sy
2spWSUzyGSCzvHVgtoaCi5cM7Yh9tUNkaYBrmIRD10DVXxlWKee5/1UFqq0h
X2wbv6UTNKrJxIDCKRfYspjxd/L17lJ2TNf6t5AISo8ZcB2EkWrPnJITof9b
IlLerRECVFmmOOdnt0enjzxyLhFqvab9Q3abNLsjTSO6CsxZZkeb74NpHGc0
6sIpINujNM091jkb2fqJQ6R7yeObw2XsTDVtgfPsLFk5JoV/HVKiEJxopmiB
vkax8GcJd/vtnmblSNOVNKWHz1Non99MPO6GXIT4xMS05CwPLeC/UMD65+os
+JScpd+D2Y+0ZR/YGttQX7vDTg5/WW2hwQoyhOwBxnakZUgADUG0Kr1NUq+D
dX73RmysSnTtUk9a7kKFssVPNsbKN9TwtP4QRPJCwOn0fkd/xuOPyWMn3K6P
kh5NJabnVCyxIXzDU4HO4uGDA6SuhGSbAJfByo1PUzE7+M6TvXIkOY0/O7Bm
iKSgTlKbgrW7dI5IgC9hjHsRHqJUl6c53/4VJQLIlECMz66OKJGw1vjscr6A
CmJaMrq/+ONNEGMLPpgQnmXPMuBmNg/ko5UV6+VP7Y8BjFBGudHG9kkGrJhg
FBcmW1pVaKuSBQ7Wqk+QL7IHqGiXXPaWobLSmkNiEnU9B8ARxV17ZplPFE+k
VubwVBvPK58BTlZhsprUgbcu1ccbqpRqu3km3VpZhg90eniCOeSyVtGddWTC
i51bFmxI4smHIjlZxWMJSiWRqj+E7pbccN0+vjapqjqhdMZwZvIqnNFNv8CT
tUU+jMRUEMO73B5qLEJgzNRQ8zIpx2gY0IAE9t/OGnpBJko3CZkP+11h8aJw
3YKKbrmanjAUgt/zMcWMHjxfaIslEPsOTSa8SofZtpSayRpn/aSdSW2teWo0
rbqZD4guBmBzSQodMfJ8WxoHtjw6XlSS84S9PGiN7E/AQNch651QZO7huUGj
cwYWagIsaE5xhhYRRYwWl4W4ith+ryA0EkIP7LxYkkkJeflyoKM18GEZx2JP
0GlEGt5kX34Q9Mx8pR61G/0W/9+3qx0QW78mYl9pSLaYMaHCnfH+KpRmVyWl
Q2Vlic2J+HZwd9EFsYP/KYW6dc4Su+xZV1FuWonbUG0rV9OeldbL8w8UUMaH
Fyc2+cGejufsGMLiFogttnozPImt8VN1AFKNhljhoILtUCYFmBt6G4uJ81ma
9PEgrpj7BC18+Rbua6Wsi3mNCAHM6Vu/iKe0HelOBTA+vQk46KazSq27OLwt
apvZJ0XEGjVkpD0ztMUosLUa6MKdbroEkOklNWBLr8lnSeLyqJmhIRpmM/6Q
Cak7G5ghl1vfL4cctlqouq4V5UDA1op4kvDiovjPxzVMOcp61l0PKAlX5vdF
9bNN+6rk5eJ80fDVNY3qwtsMtyNyHHz3nlJEmqcLNCzbX55Zf3GRF52N+syk
E4ZE2VSjlVIpPYYeqRlom4R5zS/jbiZDZsOWkX5ngtR57VVCMkywHpQfmwxt
RPQs6Or41wNMYgORQSaH81WOWDBR+Ogt6Fl7018Q9oeKHsXAz6tdGmMF1EIM
IofKtpuyRSd/oGXyXcdDYznh3sqBW7W2lLthBmqFJ1hPVqp+qP7aW+pkwx1v
16r3RDMg3BzneQ1RVmYMBiFPUj+i+WJ1l6fSnj1H5FZNSAZ7O8kFEK/osZpZ
bTiBjoYMm9YCll7yOXJwsPXM78kTHibQbzaZN+D/yD5cvCWJm/glc+ZNyWni
95KMMKZvfOH7ffLqJd4PU/smxy881Mr1Pst3EbaMbvIQeJhXoBuBWY5I4WmA
qJX22xSqY4mz6UQ22EStce9pAeFEPHgqKuloUXYPAR6kXKv27hdQTDtXgnjQ
Z7CFlfYk3cdX6Oak/tncvX6IEPjPvkXjPvZk4LVcI6Ra++28Jr82lnDl7n41
/mW8VnUvNOtOLuI7xa6mGSN7VrVTRViZNPa58gJ9tb2XtPgXH5Fx9T/oOsC2
hOZv9B4wYPlyo6dVASdjTUp/tdE5QvCSe29bjIC1qVxFMCD708Hv8DXQzLpf
kQDCJtco1+fifmdphX13ejyTI9XVCYH8aBn0XEMjGMoqGZ1JXlKbnDIHZwEq
Zy/PZXd8yjpY4PWtAL+KnNymP6QDgTeiYCWbm4EhsQcI2e0aG5dkxtMyOq5a
VYwFYJUCASSKSkcLA0oDYd/mYNi+dfZ67A+MYhycpM4169xmdXZ5Gx8tgF10
K+q9JsNlgG7fCpEomFLG/pk8NJBYQIKOMg4jrl7qgn+m5igDEhjqY574J8ZE
g10xy4BRX1MKjA6Y5K6NY6H49t8cqEoDMDsEhvAag6mwuUW/sROjl3dM8vi9
qg3vt8Kzo1uW26QwCarn4sr15Ybb8w8OX6zSg7XJLohbLyjHlXH0VUqqCciU
+peh0/g8Dy1zzMX3B13/FG/LDVWDTLNZ5aJ0+X9HQfwjFZdVqqFtJblOTAd4
2rmZ0I7iCvXfBu3U7cQIwS559rMChvRc2Ursu6Tc8k1EwNVgy4rOUvU3Rfur
xWuSxDTEKbSA53Qo+0fIL3Ifo4Tv+4o76ITnr11Y+GROLGA4Okpeggn9VzFj
RqtyL4XLCQo7Z7SR+bYnRj3hZNuqjYCN0atapN70QEzd0RXt153/dYUsbDu0
rD7edp2p/VwnVi6gGV9wnH3cTaocWB7yK5SteW4pL/oIkbaLMd0BioU7gEgj
MkatsSPBA5klI78xmXt+ctzSgTB33l8c/NwuqeTkq+Bpc8dohY18VdGqqV85
2reJXoY2p3aaP5fMirJoaSoX6LVdvZ2wSHaR3pyfgVcXuigB3BT2HnjWacLU
6vIfd1FAInoAPvY0P81ynDfLKqwjizXPfY/39gWsb8cMbmRCMXJYDlmn++/T
X6bgAOhlRII9GJ+e5ivnY0mt15Q596/Y2PqJcTvi4hSSrG3/MtqSgCnOpCh2
PBYfvQeEIvW941yU/H/T5EBnb0sTzpZf+2Ti/ZPiLVvSalhegVRh7+YOeK6Y
SNI7jIqagOYmQtw9O8oyKHTRmKVn+zWZ17OiRYKIyVC5cTsIe6/aQRiJw+Fb
MjjlwJLqC9ujRl2C4IaKnfmd9YfsVIglcvL3z8ZW4kmob8Xgl4TUk+QpCUh7
WWFiNmKajQLTR3vtfod33pUUYrwGk+qY0oZNN+VBDsxku/NOchSYG6EPU+6m
zNYzqn3q3FPfhKILxNIt37b9/I6uBniYfA9rRKg7m3lJwZcaSdS+Dyhvd/sx
hnobejJ0AFbirDr20NywEQtLxZjNwFa2Aaux2+XQYCtSIAUEzN/Ztgwv7JMk
wyOBFY43izulsrNPmeTuOpJJaK3fslNXHioUYIcpqSABW0VHyMHVeIvBg+Lq
dvkfUaEqJL8iDbAsBdoGAgGaVwRcC2zR/qua9dsArj3Q/OpQPsTpg5JCAefR
t5RMmLb4y6mYZc+66YIQ8sGTG0hllSISBc/Ts7UcCDatuJL44TDQRLEnWWba
fj8dVmNTOcwexk74upFj4cizsynGkcYyxB7r4fMj3Gd/aYciCsFVUPjWZxau
BoPfMKQPp5wrIZM2HdozLmzON/aQ6CXD/l209tthIqp2tWC5lvNqkwXHU4qa
tQWYs0LreBmmd2teOHXE+uhg74nqOlNRckrwv+014YRQ3HHWeJVE/P6Mjz/C
2jhytLtj1R3zfxm0WAoMow9cI95INDpfKVJ3LO9QozEm/aDJu1K/QMW0kCHV
j8XfR/J5lJ0qWBE261Sy6CV7l8IdyNrYrexLJVZed/vDVKkXd+xru0i+JDe5
++aYtHQq0UqYgDfSqgz9zeeJH+qO7NGx3FlN9EzMxjsiSade7w4Nd0i7G4v3
f/sUAbQ9fjfaYA6k6sQs0XNqGV5meyJQxrHzqRJYgbNQ5vplxe+HF7dTAOmE
EtKOjTUQR3XYrYenNvPt0epyHaMoRORGAU4B7cHxiDJ5ColX/NGcCaekYzuo
riwGZbDO2sbvNfbwvkOBTkpSjBUiC+DcReR+0D6d1v1D2rcc8Zjy2FLedmj7
kA4g+ziZaT44FTkYeeH34om74WzhIuvLVq4KC4HPeu/s7W97riqaPlHGfvED
jJGULu9h8JFNTdJs4WtirL6m3RsZMmtydb+WhYrorq7dS+V8f8GPYPb9cy9X
RbBoUQJAem6f4hS6v+Lo0csh271qfMKe80HUfiK2JV/BvXVMqb7cKD5Ql78v
D7CeQzWdXuAYuKs+d9cqP3qGRXB3r3dRetoLaXpIqd5fGALYKfSHLhLEg6tE
ukIuBL7y1AarO9NtsNqi8DnZJRlv2HMuqQnISCObpxShLxGHGINGHHWBHn+7
CmMtC39VUVPwNLDAMeUuNWU+b5VWBjYwDpT0fv6A32uKqJ2miX0uPvHlTMG1
RcO+U0EnOJs2SrC+BgUsQ5xR5W51A4aBRsJd9zA14CXnafRxIc/JOadPA7kl
UETeeYzGW3BW+NeS9odUE0MqfwtpxKqD4ysYUmG8Qx0v1X/Qu0pqV9swsoHi
cuafVrXQvFolJdDymNGPRrJkOV9TKart9lJsdBTmoOL3woEDIeLiIB0H0McL
lF0DOhBEOZ79v0QdulT7lpj0qNkcJsirJRzBFV0xbIMG9uOzfAQ6s/PLOcdU
ToFsX1O9K15dXIO2HKipTlGiteP6yjImPuG1CM/YUNxR5mOirfV8t0d5q0uh
xbNjW4+RXTIXxTd8H1erQdqjqrH2KwGqdNPrNyMPRpzt+oYbRbQbsWcDDi3E
gu1JtZUOXxAQ2jEl4ndT1Qec+pNnB2P5yVQZcXB4e/ZdDV5ukMUaM1a0w6d9
JWMo8HhWPm2mA8V25zSeMhtkJEhrC+a+Khy5kqnmNu/APEFeFKvCy8tzI5qm
tjVVkJYXamnRxQ0zrxFekLsDllz4HdSFM5+0Kx4VJ4GxjrSXTizyvMMfpy7s
WVFKZp+9vDbO0HcAeeZk70cD7lMy/p18XQPHEah0dcr1oB/1Oo3NghcUckM5
8JfuG4IdGwMPPs2Q0JB/pOKp8F5QUavSok6E/qfEW49OA8J+SJL2woNIjWqh
uhnTWIaUNN1xYUotR0D6JDHOup/GHlEnwEC+eOgKUZtPKpTCCaTuqZfs7xHI
/rAedFnyj8UZZfYI3FCFiOWpduSwcbS/oYh5BVtUKNMXPFS3sfKIk8yqKq4x
vpe3o35H7OsDWDKWcViGGDd9ZPhsXE25pm3EqM2Fn1gCqb0eh4kgJggd37qD
5+YfCwM79kLEwLIuxeWjwCP5fiD4C7TPdC2Xzu+Lp0kDjKJF7NwDCu5nnRsb
VlTZeq+blnNPPLtsepgCiODV59P2HiNstjXTIPTau+PnySRLLar0qS4kpPQG
W1yNy6J9Q8hCleT5TIjMsxlYDBFHesuCO28Ufl2/xQGObbYZ5ajHxD2eYKMm
HEsskMefwG5ely+ntaon7XWmNRceUc4kJlnM7NPTXTBjweEx6ccvtX7+bJ8c
xOIs6zPDKhNUjyi3/8q9bPearXWEnFGAKB2fUf5IffDFyi0k0bJ19o5qvfrg
oIA1P7m27SSVE//tRgVHUJwME5Q0rsdpV5tgWCUXI8IUiaT3iWrHUFPD4gAd
mVho4PQIuz6ihpFsAoETuvjb5R/MfhIIJqQ90T/0hS7Qad4+hzb7KwrGMjAk
3Mhtt9/qe0H44rap5k7z4XpdL/zpT0Wr+bdnX1zQSBHkonCl/HFTulvZY8Lb
3p29NFzJb+DRBonQP7nzx34/M1K9l5vv1gDt1Q/iSvnS+WkBLwBD7dOV23m6
pQtbhYnYG1YGMa+0BLlE/gIyVE4txC1ebWXD3FlqY0m1nfqECyrQm5i5wHhD
evp95hxtaNw912v//2e7gPGPq7/458/NXGKu8ohDjbbjYh2LZ6xxQUmRfKD/
Rh2VlD4XLx3fBYrju2cqYn8HVKbx1XqMWiGEe7PuNZ2HS0OpagbgXFED6Isk
UCaA198a6xM6MOSeABv6zbzZIcXLidCKLLb0ADnDPLHajSeaMzUzHjQ9ONTD
ka9wRO4oTfWa7/JxjJpVh4m8ZlfN4e1X5R/GHXFUmI1P5g2RDwj0l93qqHxq
6jmzdGTfVwaK5bN15bvIVKMrLaVOkhP8WxW4FymgHsTz1OGQlfHuvQBTyg9W
vWQXpC9EUwgou1zDNDCRHZmKcQ9CpOMtG3OttuQ0N6MW00TyrKX7siHHySjF
8G5wOy27UHPpP12JUXuq7bIO4X0Iz3ZBdFC1oUYfKCKPhknYwSb2j3JyqXa+
g69O0Lb1/5wrLYVA2JFUk7zhCE8BnK6VvG0MfWdLq8lc0Epe6F4IdG9Cdc0B
5rTNyUuLOg9XOlZh4gM5rEWwEQPUhyHTrhW0d5UbW4tdWsp3Y68WMQaM9wLT
PIHLIRbVRl4VLTN9qm/LYy4dc+LZmosNflT5AXPl9l9EATZfS79eYwZ/gbmO
z8otOGmhtTiBal5tQKHTwOh2FpKl5vRJCBhXYk4xG7Dgh6ke6d5iMXoSf+Ya
PAzNtjyB09R7GIN7QnIcmqWCVplM6cBJP6Uh24ejOFVk8pcQ92dmoPi+ER20
GJjloPlNcorWvKjykps/q92G8hWoC1fRjfxj3Nad/54ys9jxQQcvtgIyNL8o
MGeFtBd1SyjPS99iBbiyJezKFMsfdaVlsarnJDNq/QNV0L/IjkIvhGhSu1TX
81JGNr/IAmP6zwqG+sXZrxGUuH7ECMGFzjqcd3eC6+d2g8TUvJ5GM/Ql1sHZ
gkDizHqvktFCeGlN2w0oQnRxFLtwI4BaRU7bTwJacF0x1MvJHx2FLfv4ujla
p4UClWpQDLk8LGFUZwbrlCBgm5O1bPhcPp5bLtu+Ext6G/D8pbF0dzoyrqg3
Heso1X9bVhbC0nODBw1GS5TKPL3CDEpPAy4syPoF7sldKwqw9ohit3eoN8AZ
OoDpeewRB6dQbanGAEMKhcJZSElf/cghS/llS1N5XRINK/L3OAeCMQJPYcnz
Gl+LXU02NvvKnCxJ1OZnvRexCRc/ukLIQl6Fmi/UCbxNygv3/l1N7BubkLlc
t2AGPvSJ3TuvHWuL8mytt0gP9lBQWa3Fd2qyyBR6QyfFAcLM8l0tNkyhVKrT
lbwlTMSTxrLLomqii8Af2TyiXAldWIEK2HURA32F7/Ve4b1vqI02Tb0trq0b
YYghp8gK9p4UJL50a9PLgXXoCDtBCRlN7tDbPEN7GHMxh8c8tOgc/h/zFowi
iC8X0KGgRSWrwWu7hs91LyCVucnRagANWnHxRP+agYEDW/jdNdZGkZAN0UWu
PODCGBYZ7SfPSjP6d/ZPVqGdl3KMPdR1tx8/vUt2Dicmj14ea/Xm2PBgJ6XD
R+zYclN/lzLOnUYXWMSvkiM7+U2ea7P9+o3kevPwfuvN08DxP0ACPONO5ziJ
JBOtbH+oFgsWUSXXBajOOHfeSyauX6yrbSt5q/HR7xOQXIInGefPEJfDEu5r
UM1MdeA9HEma+JnF/ZCBWTa7TPhe6vNGlEn9IliXRbfVKmos4thplgmixZKl
/Ac+t+H4YLo5S5Xe+PSZE7jLTH84VANwLFWE+e2y1whQUwTHBeczAxNmU4GU
h5/RYvsdMR692OyUwdIsm6XTfKeuImw5v0jk33OpOAD+GfJSj99h+JeQHCmk
KC/uPCk0mQnU7oBYFs2DpUnpNum8bUeDIpm/FEiqiLPJVqbsSNiuGx2HlBPB
MmgDdAnCuapAjYsRj02ZxCE21BFge2D6FefuDt6CTQVowzB8YwUHgNljcGSB
c8YKf3NoKv45R70dniSPEuiQ1p9RLKKE9Pm5khPYhRmbJeDIeq9GSlt5tCAq
Ej4d6ptjU2smzO1tQJMC2dbUk5ElOWMY1lTsv3XCZcoUu3v5ISNW5LtTchps
ZUOoVHguPskGhjXzd8yZTTIelPw9F1f/sj3lGf+t+n3zV6X0AdRCZzk97lwP
adZcIjONDPJWTN4GxWyxADHcIvgwu2cxf7BJVyYmfLVfC1Nws5KiCQu1pPhy
rVDXH4Mzh+vCEiVVJzKdQ/EY4OKG/HcYhjBI7Jd2WDZbTQeXdcH+Tft5b9TZ
w+nutAiSC7gEJ2xPDIv/xq4mUi6MzFEChC6FGsqDjVo0uWjJLBxSuqL15Ikd
Nvl0mMhwcekQ0sS0pICr+DY6PEebZelFcO/sgy1kP/vSoi/6tPkhYdozZWAX
mjeS8OQ7ygIXZKS66HScxN0B6VO8SJVQKWtdGIWPzqNqdJTEXm564jutb0VT
RM5X5zsyBbYZx6Nk+ZILb3KcRiwugjzakmFX83UuqVH7QBebErWVu+n0NAuE
wGe1dTZksESHzoMm2laG8KFlrMg1WBBiqgGmMkvro7IDH2Jfp/n2Ey1TbX2c
jTYow4EokSmyy7+Jkzaic0NZx13FNpx6upny9XJcrINHN+lQetebq2vqBrYw
CtqWY5Hk/JJJa396JNX8QvvCKoPKCHcGKvBsZokDlPJDAYPtSLigGTpnf1v+
3iWN/uM1utF4RB59cjDqP4lBlXgYVT7ITrlTXN0yLr46UtjevPuZSNMJ5Gqd
s7/3F9+z4nr1uONtKOVHrJPnHKVgDFL3wttD/YeFlsZtwikBJID2EmNoctql
skwGLJNLlSLCX759eKxvt7oVxfT+kA61vLBW9dAJNrlyHE99vwJzVMIHWn5O
BFirjzGBR5TC9tqr9hs+DWgsuPk3Qrp+3F5du0/kZrsGTQikMmiHqrl9m4WB
bfXJB+bLevUZnEH3tOGR6Y/4vG1qNgwjjcJI2E27Chnp+67eZKGAnVxGVa13
mILgNhcP+o3ALEvaNAc0sJXaFcuXuU+47HZoSL/wOESJnItBiXlQZDuQ1MLa
PrlMsah2k/fh9BrLz0E8UBbGdcMIJJfXhEQHVIjAUls8qKOu8Na9nCZKpPYf
b+MP72HxpuRT5bwpXUl67fl/C9Z1cbEpSRhNU3Cpwi2EG/fFFrgWImBRzSKX
ir8rrHvKdW41A43E12vZdwes+lJBuMx2NtmIL7ZEx1kj8tIY3wUN11rYSGTd
XFMmFz8I7jJ8m5XYz8Rvz5JeIB/+Uat2ujMQubriiI/FU2VAgNq0DWOlTEow
9+Wrxf7xzcsxDTyJI6rkwqt+E+WiKIJc3CpqrLzGw3I7U7OFmEy+svOjKRJG
LC/+9DtRJnOIdp4b9LTOO1ibEbwiZ9ju9pq02KTUXwjhvL+4ziMMJi1UIb23
FZCwkdz22cF9n/SnvlDG65ORqbF7lgpaAeTNgyUhDDiA0UXznKUDaO3RyN06
piaG4gVAj32ecPsOjjtO3IuZSEHjh+7Bsb+SNtVFcIsSbU5oMSNMJ9S/zOCT
NKNDiE+5EieKToNL6RMbHoMxnTyjAPNTmfCB4167orJLTwjcwca0xQgqlBAr
MFXCakYDTlRBO9i5fQgf+PtrhMyVc/qA257wheGGm4cKC/L/A/LRlV16gl/J
pUZoid2CCtfx8OwQvpivwEV+vYNpB/p6Q+T/iwJiaJFMBycGqfC4+8jDJFIN
3BMvXFkXHUQ1dH62tFMVPybkkPXXCeyrNAIqTo5JKlhfYmQUZYEonj/K4Yep
abnhuMtN94TbuGtXvu5FHXp4jcMFmWoBo68gxrlYNNNdsxk/4+VK7jyZgDnQ
B3QdIqf4U17C6Fl0Bnb1LHLiuufQXOO2gOilkDhVu+7zwfxUenRlraStHCB+
JgmFCHjYrdLDWGbYQC6hEUsDJ2aI3tsE0US7N5+MbTd1DhbTOc8owxfRJlTu
RB5yTsCHKFs/qmavH/uttPIPzHWJuArjUkLMMehkVQmgQCt8yuiyyDoJVxuX
cyWKEnqMjrnKgsjR7DS0OmMBsm8pUfTsblNa7u3ZLWo9CkXm7Fx45CsgiCIJ
uhC65SCFChvc3GB4G7/BOplpRbPAtfDpNTgDN3peAgNsJmJcqcJaFv221QEt
eQ7RMV7pfjegR0AKNdv7K466PvPhCo8UOAANohxy5SyP/iK/RG/QMhHqFjYs
hPVzKX3T8IgtfMb/4y0gu16jn/uYrc27pUtCoozFelq03KPjkenotDv+Krbp
XZ3kr1TXjFGIqDdGdc0+2PKVvg4Ea+zAaoZsfCQSAZPfGpS0P742yeC+4Xli
YNu87SkW3p39jmhd7dZ4XUuxzioyLfQ0O+LbAPGohe9XcYInJPjD13mguFAb
ECFAgBII6lbpzk4OmTpAA4W2+W+SMEKxc7lSW6uXIvrbOrLxBW51E6p2Xk6Y
Il69y5M7zqm20Bpd5JsAjBO5sHrhyzMaYnp1crcxsmuogsGi52gEimz4+bAT
/3uwPBU2jyxF4tjj2Y4PL2PhSULBFWHR+OAxaDrs4tp9CgdqTy3kG6daNo01
j3S7CLfDum/j9ZIOLpTflIiZVcR2y6HblwPzO4Cq6MiY654xzETetedmVoX/
2uk28Ds1hrMMqXPEFaziJX3C9uc6z8h0/F8H6zXy+8tXtPcQPDBEPBhmNc6u
x/FYYauA21Om4exmvUMW4JHhAlw8jGhLA5jNhp/Sdhrf4CaBSAQ4at6eelXf
m4dRo3j9Kvv6C2I9QNjsLGuPyGSGUXPw3IW7v93r0JE2myIuGNe7uFaGLOHU
YPJ1bZb1aFnaFMg8tOJrVomtB1Zaj2DdODzEaxhxrNPqdLLCYdOZeZmLGAnW
+CC4UpdhEtk1ZJTuXPtKPE3jzXJTXcr4LlWw5zbbKfgYiHr/vHFC0JDgRlWI
iJfYrldnAHsKXUg/SfpwCvmhXj67FLv6Ej7kKa/zIs5v3czaERDq2RZTlClP
h+ltoILb/lXyZYSOecni3Wk6sqI7mswwarjG/2jEZkhaQsGSbEEzYa3scX4p
mYcoXF3Yhje9NUgtBrXWWHWETFCCdkNobeT5f64iuWYOwH62+yibsyV67eET
FuCb8i8q5P7NZOPUX7GTCOkeqaohcF0M9N8GpKn00T4S9bWQk2eIukDUz1Iy
keflb/qrvzujMt9UUuDQGiVlOMyJm+u5xxNONpVnPMpu0A276B7azSPC+SMj
GSuCNYEMvh8jjARxLExu4YqpT3ZL0LLjrpAzZT8emGfRnWwO4Nu0HuUEuKrL
inhBm+93PtGsfMiE3I9f+dTBzIpJ3ktIoeVs9hCJ4HOPtS4ctzYIAo4Ej0+V
GlN3D+ixELj0yby6dkvBBBRbcKz+PnS5eMpbgwK5vVjigaDW1jLloJbYtGL0
i/QaU4FaS40cnwV0psIwHw+DEDb9m91naMSbZ7jCwXRbvgngAbHjv3x+jlei
WWIb2Bl6uexCz30ZY102+JJBZ6mRmX803zsQYNKLa0yesD+4U1Lp75/L2+aA
RZLGeMH0jW9lIJWwO9DkIinICdNZdElPMoVvKrbbRK1ULsxIj3c49OUoFoHF
3hp7kT+eycW4iBlsHPJbrGqkMffENfcdZ/fmOTO+y3oX+Sm9cOf7ZknGQ4y+
4wttkrQuKTsIGFJRPih8zOw0bVp6Xa/7n+DZkY944CnG1iYzxnCIQLJmnvVj
wG2vBk1lTGKPpsXOny294s3Mh02iAvDz1i+GeKbhV67llRzYh24pVXqz7UZF
vlStAOU0z5qvUZtAaMAfZiAWuKRSS4vtbWffGQIfulObg/EaYcxU9DtrD0no
IeZMBEFdmwL1aXYZ+WhxIKiK9NWMgYmlYebl5XTYCazSsnN4SoPvc/Rwnkau
8B9yxLQJOln2k7L638gXboSomRTejqX7xQpGpzd0XppbINYQ9exIROjle8Yq
jIQ4J5+GeZVTiYnvkqlD+LW580MbhSUOSK+sk57XQsdfnUu4nh3ExREd0/5J
YbLGxp8oGFuRgyILhXqM2vUf8fvdTR6YeH6eS60OtCA1/HPLrqOso3U5j5qi
/HLQKtzJNNWieBY6OTVdro4CspySBSKyUA4WMO9jkd9tY9Akc34ZMCBoALMd
fkMyRxmp17KVb6Rg0RM5EvemOXT7GO/VekcPHfjZHLH5EHEW8UInDSp3kQHq
OJCUKdqoQSMGcTWRdxPP/ETCg2L9c/CrJk5JPvK5M2K9mx7nVjtlEVd8Qmsl
NzzprOw4jS0Rg1mUzI22bzg59LhYvlB55OCZ92cF9mxEp9t5FlBj6veNRfe/
a6DlvRMEqlK6+p9kQ24AxzgPK9r2GsTpwDilhvgRObD+rf1XsYWVMStw+Bn9
xsOdNc9YeCAveboedd8NJZcO3/0SCH/7YSrGMogXHpGl4vg5HEHp3VIpvsj3
c0THaJXCwUF5K7dwKHdlWEj4FLIqCJojKI+rsOq1fuGeyrtRBMTMfvxSIL4H
xdm8LZyL8ZbR/ynFx748c9yWXLPldOIr/mYAFg2ay0fMwOTbDUUCiWX7MWID
dj2nYCj+8qHt83yqP7OrfTCULWQjC6ztMmUpVBw0vIqFb1rzfZsoQJeZYYrr
tTT7vTdPIlJxRyjx8V8EO2M24r6Hknar7KZyt2u/Wv4iKguasX91zxHeZgF8
uMcOtpvpPUomh3McaOWNp7xfLDMIwPYZCql2UIpUzccgakQNhYQqIetsbUlQ
UwqAURCL863PgnAIe2K+EMpOHCfrMJxp4QzgQ3rO3zvG502KvAXygXNjfxFh
zwo0LqE0A3gn6gfOmHPFDrWJg6jNWOtJKdqXh8SCDeBp83RpKZ0xLTXAQczt
nodKroVxGJ6ddpVJn1EQRv9OTlx2g5uZ93xUalhnusdtHtYLduv9241NdP69
eUu+/eesy/OcwxnoCFuTfQglNh36PLlEU8p10UG1eHuIB4fkB+pE4va9IX7A
SXImCbtLfsebJneNhnwTK98miuY7ISyZhO/nG38CjbyX5iEeicFTX8fOvD7o
YPehE2fzVwRMhTH0vYY9dq4MnYnL6UNkjPIADvFwW4VirZp6BEJHQGavvXHZ
EZxcYq6xDOL7lkqJvty2sVwZuKbMHP5n5zC+japRnjG+FrosbivmnN7fJnjD
dy7+y3ebZ4ENuFXhVtSfRMfwWkiA36O3CIPKz9fJKsW9Fv/LytqPQl0+RO6N
fUNbzExuiafe0UIJEKxVOu/kGbyvsoi/Ryc1PTULauAI3uf3KG5x4rDF6R0S
TDyJ/LyyUe8g6iykDe7zh4aSxmaNqs4fMR0/usbmUXCYcDWc9Kb0pZfFk851
I61+2hkZhcDtnaDqkIB9bu5I47Cu+plE+WVoHRptUpoHYrHTaxuMfpMK3k5r
wg7mRFg3EuASsUIJpUcMM8LV7y7l5ff2J14wrjMIQIfn4DmO6BnN6cqeQ3cR
aeLgGYNdabVj/XbQZcWD5cnf5Pxy/53kge7LvKVt80tEzqF3wkKinew3pGfQ
VMHpT70/QZ0Knz1IcWQ0H8jZmFa+EYYzjtgegu8EyDtJampB0PSd0Wz5GCgs
k8ON+jKAFJSVB2H9okUt818FKTQ/J1dozeGjgGODTWsjARHH8oSRFN8qU8nr
XSA8fdXvsYLCb7cO8YmSMDFV6NOGpDTZ9x61KN0c3BML+rN4hSGbTJ1NLutd
ZkDptcvSoewja96MC9BU5k3wBLFWFlTMK24ECZ6M53dOFHjkxBpM3YFAoKKE
YaGGWFjKqVBUAI0cRy+TaFulpz+WYqqT2MLseEOPFgaKlqgkzjkUaxIR+oeS
pYphEHcDmMNXLwZmcoK59jE/GCcwHtgQZL+lwghjJdneVJpCT+WJ5PKby56i
d6F1dWMEkTJ7w0HJW6se1ShdmUoyjtB2aIWCk7YQbDVFxSkQhaAhF83pX6PP
G82VCoQr4s6dyWnOY3cxw5+Q8Z4ak6B6dWusdBFRgmrxPjY7VyO0ZsKB+Ekm
wxzbwvgE7q/C30u9aCc+byvzcisfCnM6/01svpHC2lLZIQA8gGyQjy6PbsZe
kI4qGxWHWUn4n+hm5ODdnXlTT3COqlj4+ssKnys0qR0BUchsj/xCzEMmb40w
2y6GIqLkc5ApN3cGH1Bw8cS2dGm8JFD4i+Z9L46L+vgeaMTPsdrOARtHw3SJ
j6p+N12O7SpKpuhdQoR3mBqX/wFGDwSkQJ1BVrXpWQZH+2LBkb1XbGOF3WEe
+IypGEmdLa+onY4SyrDf52qS5TqNnd1LePJEcoP3nlDk3THmx2EDzVr9akF/
klZTKluZY+GCt2yuSp7GD/5yWuECqUT13OLTavN7n4fbwCLELpV7lurATA//
VGqMjouhvWa1Dcr5vy22AIcktX0+vRfCfiMtQkGUbHoAHXvEQ1sPw2u7FvtB
3BZHL05OvM3LmmtyzBzaHx6ktbHAsERLLixw9vF7GsZukSysH6bLvNG+Yw7u
q5pytFG/X6QG9f2eq3VFDr0m96XrVEWUn8ovhgAWDCk75a01+pu2Y2sOAZFi
MSQk5L6kzNk98mtUh6EnVHGZL8pvtSUobVh+9bRR2Joe8kr9IBMy4rQtMsC4
eaai0YEdwQA6LVMn5mO5QAmXV8PxByXibCWd9VgKmf7SYj+EXdHRrr02c/WB
dFujPw2x/ABtmdsvTEs4o3jiYXFsyRP5atSXx5PSn9kryU4QXpMrYkThxzke
2dSzrKLizUnxTaXP1duZfvjJlGqrAOuh4rCjppIcGTJ+/et6ZrKEJixEtshB
y1foAX9Ll/GEAXEPsfJdTvS9x5n4Xe3vv8t41xRyuEEyiQzk5iXvzLk5vts0
gJ2FjGs3Wjkof1W5t4mIlfONeLyByLcR6E2BFrfTz2juvJgaPTDpeLMGpS5r
gBIHs1liPMcPpRqyJGFUujR+w1ymlZ0XiHMVOSB0W/4XlPuG6TwbE7t/f7qs
z4JZW3b7QG0r0W79owSkgPOOXQOXCR1QYo1Km5Kd6p9Go3IE1jnQgDNuEsmI
Ega5ZsU6Uz/YyiTCl4fFOuZ73RZjnaSuDj+2cS9ezAY3I0tB5QlvE4hl1bDx
ZcI5vcsdrJwfyBQSSqIot9Vz6BmnUyhkTY0Eqa3d333AK5ZgNKYIZ36YQygo
va01ZuGbbhiHWOjENOc8cCzaNsP2wzm8MjLl/y9smt36CFbgukM4NDrA5HFu
sZtiyuUG9Ihhhm6oVd11w/XFzcCztcW+PH5Ivym7t9LG+nBwJZU93XCW7q/M
uFabdB+r813YWR5g8XLgs+WWAf4EeDb4SJcuaEvebhOTUKE4Ol4ykPjBkCeN
K78/6OUsxaRZvA7teAE8962M/UtlAENCwEO7C5HWgeQy1vrefYp/kWqOZ+Gg
zlvS1zyRFEooH7n/cU381+X6aTGWtB4GO9pX3tzHcoLSMZuW7kRToI0YdQzB
yztEgJWtfE1KsC+OVSy0pSz5MWpfHQCU+Chr9Jb1toIfID7JCbmUC/ANgQ1t
Cs/DDH0BlSzHJ+FIthQg5UXUGrkRdszgYcYbUnOmo+S7myAHVUot8tqEQpg9
8ubXYsRW82HNGks1MavS48RQgqhYVdeUQzWWfjWLRv6Zcel+/BD0Lugyxlpl
r23L4nf76wC2HjSc662uEKL6NzKcKtADjxtPZTt0VtKr3yhSO0NF/QD8mdYJ
URRUHf42kD+curEqQDYWRqNKVJcBAGVm2sfoQ/UmtyQPVqXB1e13O/c0C/Ak
MjlMmN3j91JjVcsSCQUO9E7ATKKeVenQnMLB2FdUCfsf22Q7+vEfde3/Qstj
fiWOjIwmfgLyawOHq1QbIzfibwwLsuMMNJbNGi00QyWO1yDP5iJpnRmM6GqM
g4ojHsdi+7h+BTbgq6vRbLEvSEb1B0T9iOAKm6xpmRHQzf3S5F8VBc7gZnRY
DTmexHPQnN3U3yE9SUdezlq7t1r6MQ0d6IWTmGt4YztdSYRPkzckuR3HQRA5
O6/71nfoVwMbv6lzYwsrcpKMnmsSjwczWSAIlFt9suXMoO0IxPSYmYl3361/
BJgGCniTzC5MsGYoR0W3v2UTipmidvjk6TzBXoIauBvp7S1BhKEnIaSHd756
GDFznT1JZZUb7xHutEETYM73nlPkacppzyqfVseBsI9dJp40XzTfMff+/HNb
A+JMbQRgsAyr5QpTKcY+Y/w41O+XO7CQuXnUMbeCK/ZCEVXWTxtNrlMMBwIg
LVXJfhmykSRm0ec32iNzOfo2NDn+cy6UVWYinWc4k18OsKw8o4FQqVvpbahr
gpmSKLBwMgNG3NVhoephP95Ou3AqgSqDW4L/zg3Uz9ev3TXEiJBgiYTQvOnD
WKgXXFiKIuBeDX6FWz/BGmow9rNlBOsvEy0/hrhmYKtExfHxAzfOx3TzX1Od
66y/lIy/tJa7o4AsuJlmxxHvy6r8f25ZSmgNC3GPaIQCHZEXKWE9y2DMBNDm
vkmKzJ2X4xHo9zvMRHDYswA+M9GewOSJXZeT+XqSEkSlEAXK1Qku+wW5UjTb
9YLZQUO7AUE5CR35vCHHYxLw1xC3PzfnuKSOaOZ6FHA6fLzTrYMKLf4P0mzu
94jHXOr7bcWdbg8e3rPZ/lWcYpA7rIdZBVj7dwE9Rkv8qmWWcvGMMGKU6x9g
Mnls8qZq3J4pE2Man+AjJzKOmHMsSvXte3ZBZrgMpqUtUW1bDvmb66+xC7RT
fZhn+4vCgV+JGTfXgfTv0WJJNFozutP/F2CTVfsI1Er2DjK0n9lCwUVUTeqk
IEdt+DmI9zL62zs1kkX/J1LGXvb+5B9QnBtLDjyLEb6lEJZYmuU8G9TdfxWK
p+9W4dId0BLOvzhXyZJmLPRzSTVIU6ctE7dsBCgWyzAyynEJktFsZdyuYsVB
Swmk42MDVn3iqGoSAw3thSWXjnRzzk7Mr3aI3eTHWXVhSVza5Yl/waaCRdU1
I00c3H63O+2LsZTz34vpr99H4ot6QqMUSjrHmilpL6l4FTgH6pOgaA4qQW4k
buxr8b8IHdSHRhXR3GL7Iwhl4jvztIuEU8YOEM1dP+Rmue8eKmryzeDhpYvH
MWxLqR4D3Z/azBE4Pv2TmNenWkBR7VsIx1UYZ+ro5JrSNZLBk7yBfWIpLQVM
XvFK6qk6JNJBjl/VE52yJisQuhikGkNEIs4/N/NB+AiHFxkvuqUHs+dXh0NJ
ERvE8Bp2uFMMhV71dGgLTweADb66Crg5RoPWMoIT7CrytgHCE5w4d3MXX0MS
nWK8XUsAZlUgygPkIjEg0RRPV6TMYAuk3A6iuUonyk07nOKvxrUtrVjECEVG
GZVqHobEsqDyH7DTqk+yet4y5L2ThwK2HK3b5OJeKdTAICnB02oE4ypQsbbW
gzaGiak3hEEu/GEuzf/J95C7mDMurPofdel10CppTQqy+Bg7xR3hzsiOglYt
AyJ67V6E6vhoBSDc3dwBogPb6TN291TDSggcyS2YC6/2p4Co/4FNz/UQ3mqe
jDmGJ+fhwu/3cMYUkfusjVzItke78kt6IKzOP45Zn3QOr6iKXSfjF/HH7Uko
r+O5NGt5+xRarcvsqrkiS2fM7CeUPojYB/jzGt5o/Ahl2wW70TeWoQLT0Uy9
Eif2HIM0hsXgOmnhOBX5EoCHESflOESUZqaX+vf39S9gu0I+gA+GvIH+B98H
b1dMa2J+ZewQHGpc6GHGsz04UHhX/K+i7DAqxf4hTyRkxO/TtRWdKjskvmss
jhMMAu+Zm9FufXzAsrf9gOTEXW/W5pThj/0BkvSGFdVCNc/ys24KPux78m1e
2KUyepm9RY+asGpmaf1z7ONIk/QOZnf9BmEwMOlqczuGtmXAn3YmN5XsjXTk
pdjMznTopkO8ekbYAH00CC+7SvVWNhIZtqOM+K+QLgf9L5SFc5mM9P48Whl8
ZIaZzJWOcRYB1sWo3dpbACZvO/5LNx9usTuMa7kxv6in7a+fkrkjPbZPzVaq
Ncv/an3iseqdaNuaVxMZep9WJOngEbrwVpeNk0jMa/N/hNUHO4slxmutnH8K
1hv1mV3x22nPwd+t5lEVy5G5vfD0mSPzXNBH3JOJb5Gc9gZ5hRMEteFiqS3F
cs4GinJu5RAlglvBOOG7Tia2wO01bYojEtdPpFKWWo8IrHxtKXWlkgG6urni
mhya9MimNz9e7NyEXgnPGFIqW3vH5nbmJt6TDXwf+QMlxjg33YvZjFdWEBJD
mHQ8wydeCHSIaGj//06Y7/cgfMgDslcFHvY2uLLJ9UG9jydTrGQiJWuz9FOe
hFkYWJmvDGV07g3ENHt9VxNc/McA0wZBFWwmiKr0F2Ac4WWXgM8m6RL+YsT7
ugnD4PbLzz+mJiDwQt7W4aRtBSXXf2kmODtW3Lg8tZfsH+6zHxwByaNxTyHZ
dGSWuuEoBBHJXeYIJDm7UCXpGiFnLBtAUgDLzZa8gBn2C2jag+ehovCBa6+a
lMnQn67ulmaaFDbZgv8EvATWfuRgvfihUqNypH8cjYVZMHT6YFCDDrjJPxdw
kSGmkQ1ygS1gCxaIT7YuOnNeXTSu0m8v7Hpgzqm5lxeaBn+RZNd3zCaJrjrM
VvoRvDNh1ekRa4INvs4oV8lGKZf2v4DLguYvBsb9XjgqKwvqJJoQs0EiixXX
TLBrK3rNC2U72Hw88o2/U46eEp9iCs92A+r8vLxY4NuUnNnA0IiRxzLxLSSf
y5FJHoZfv880cWQlGC+dhTGLX0tIcE9XeDO4VPIye8SNRF+lMSEqvFwM6kuU
RrP+XokuvyXdKdR8bF3Ytpb0S2HSvvmniUpRJLZmFA2d3VEccsPY09pFepCg
f+xfNH2of7dAp6vk60fu+UpYNL2Waq1uCgFhEAH/seQjoZ7okzZNmm3O0nk0
SQ0bjnfMVqAmb9UuJ4mEpL6H86xsNspNNucf7ywRrP9Md0qBZDAO0iPgMrBV
dWYMPo4DZ5wqxogUnwmKt94ItVOQE2KdXdlJH1o6hKW02uodFrqPd1c7fFsb
aBYlftUGGLOt4/y/fT1hSzs3ev+UDbiChhEjL5bvjH1KI8vtqugsu4pdN8Lu
0YdUuVb4LFPiK2F3bErlxzOk7e8QWpFdDUMgj/juL4T2xHRkcMdo1AyL++ly
/cm6o1qTTogHTKg4LFgxuHvrfDUPJkaZHDYWUtPkLROs8pnoDAcm4O+rJLsW
QSVSb4mpPYeo47RfCPne6tKF7QsOf7zCkAKE5ftbD9RrJ3FAsQQPljKxeCQf
NRhIYhfWep9iiB/BEAX97bRyQqyAsUCu3KQynuJtdYZ5ri6WEc5/p/NtttF8
aY5BMYS4DiMFgjL57E3GZ1Pe78c/pSH/5BziQlJLxSSVwhXlkV7Gp9Mnhgvh
KDi6J7qbolwd85ZBcS/4vSpDr2CLZhdxcK+iG3Wc5DA0hOCL4PgSCWXEEbXA
VWXLhJ3evuJG899Njv7e4w7LsmpUT7OhIXhjn7xysVeLDFCcv1vA/IECgPQU
/JpXJl25mL9dOMvSwg435exO2Ixop1EMzjBOmTHT7gLjJOlEImDHWCyUfEy+
KcmrlZrD24uGUowxYC+h8XjLj66rObSw/Bg9soYoNgv2Oo2XWHAtsiFsH6h5
TjL9ITnZHKRkFXkt1WrsjrrRb9Pj81WguvFOzaZudfGB3h4AyiCgjntDul0h
58iVdM+lwxChTsHWAaLMxHfl/NgHR1dDMbfbIHROa1WtA01ZvsP59n+I9DcU
mr7lnRrOOK01e5LfoeM7B18iETdYEwpF3ClSqrFQJegqZuBWDv/ar+V1t+mK
Etl5cMISvCicL/Nu6X0S5+VL2ZVQ0njEi/ClFr7R9e7lyA+WZSxoh92N6q+S
eHJnCCdhaspvTLSczX12z6lES5+1mvhyjhGreT5NBMOplHwmEqoEwPJs+i6S
kVvKZSXsCvKDHcwhymcsgBV40qIl+bnuHFB/R5nFna6bjeCXudZgdZnGlpUZ
ayyP2TTHbIrijM4XxKvSc6PqGUrgPKwiqQuyPqf8DsiXt+qgYzbpfU+5Yy51
iYTNDSihPaYX82siZeONtYL8LqiOiDQLfHkUu+Kmnr5qRvQfjipyUme5JJzf
QvOWhKhgw2VFPYNkIvtD2yZmYrzXZv/Gqu4PUakcL48RN2Og3TNPeG+KFe9b
wHtukBLJvt3LQvOYKx6XTv07aWL+SKSNZUvVpIzVtN1Tk4/d00IiKY0cTEGN
PaWGMw3TTFi1SsQCN++6AiaZQTyDXLzA9c+abMjanuYr45uJFo2YCKh6yI85
/h14q5k4H8KFhgLp293VD9lFnNnP21T7XA9km+7W/OzsyfsI00mWWxWa+KdQ
RI2fpTq0uMlfQ7XDjk5HQdbUyUJhxzpSoibGloWZp498rSi2ml7W5gz7Udlz
A6igRlAXyMC5TMF2KEQHMqZql/d3bshx61eKl6vtwmm/d36J5LDjZCGOpr++
6sP8pFOPoJl4k+69sRmU8VMirEXUZOXPNSTiBkHK+EjOcq2Frt2MbLtw/fuX
BEYQpbcrH3IULhYYgJTJAc/2ZwhvRyValSoEEGjbdtL4K58gVcclGYL9V7r/
5zAsCLpnkTAnhVoxXf/qH8iZ5HddxqOIca36xUIjWdQmh3Ppvuq4sOQBwzsR
1T5n5SlyBszB8VMc+F9ka/iu+zm62eM5OHSMYKKXs1hARfx41QVfgA1WtqtL
qSLQJYvmz2AjPfqRZNEiNT9gqEbVl1dZueg//yytX7/m/QnoTj6pS6oonVCi
wrYxAPHBi/58Qv1TJkqvJPMJaFevPK7ruCs/sCxzquEHFTKyZpLdb+E01fWe
mGusAwEqIC2DnW2HGSA6o3NPpvxEt8wTFoLaHKtzUrCRsmvC0h+NEosOqvr7
Rz2EVcUMxXe5ZlNuedmLmwnnziRgCKNJeTxaTMhOjtmaChsnUAcBeVe6Yvls
GtYYGIpqQHy+vaGzuYLb8xOc3XsEz94RcmiGZ9V5pU+aLH0yFextMvfm2uMG
dafb6tkuB3NoNN32gIgnWOapn6UFGPtM3f3i9uPjCemwQAvphtaKl3Ne85W8
DcTPvoZZcNWutpp86tG/Bpvgq6NkirrLroQpAYvfj4mBRos3pYW3caGwzRlN
2cGc0CDz0GTOtxk8g75E73LehKPo5ksv24GgqgjkKFx8z2baoIAshiSlyXPg
REaQMNzBBEOhdtxoaFG0kUG7gKAUlXKrhS+oGGOhjabI0IRtSWZADwoyDo9Z
tx3A0S8lPXuvjyAuKOpQqnHk8pe9AWa8eCbg80LC6DdNPh9lJRfO4BspXdl6
tyXRTb0bO9bk9MhWIGKfKys9rKzb+C2f4k5PQYkAEJA1FTau0Eaf8udblI3H
pdchDASkPxU/6M4rXog8VIs1YjXCgh47Ev0yXVZlQa+KgeD/U+2lC3MOGpHu
39GTjbyLVLH0sA4uvt/IfG6ex+kRXdJxLLqexLnakb7/yi12Vn0DEM88DENV
A50VcXXV+LGDpLYgrg2vLPV6LlOHUmBQIDDjogJIdl1HZFAD3CQ/BTdA3BkW
MCYwU+rx804tE6HUuhxoBQr/ryO+QmDhg4V11VEggMIwESBGtbZyQacfZ9nj
iHoXZAhLRX4JY+5fArDZlCGZJK+N5LTBTnUz5bvg3MCOFPOqw3qb+l2z7jPX
wwEAhESG3M1NqiLcTje3toSFRrRFAIPBJPAIEVQlYqezDeT0tzB5Bkes80iN
IwHnMLmxi5T5KgYcvWqWb6w+CnOUXNI8thJmd9+BFt/l5wpe+i+T2We/xNrK
KTreCRvwPIwuiUMyas2R61gnPj0bOKoysM2ej47GRPmb4Fz/mEKkZP3xFyVw
bJw2r+B/P7+xTqo4cIlGlbb30hhrFDos89iw0xd6jXvobCfdeMGQMO3OsmFH
scOQgfuLxIn/idoIPgfciuFaCRdkhb2EL9NFIgBknBE+nUFb86wUBL+pCdCr
7dsnZPJEtyzfQXYQGltEHUgaZHX1cFJdfg4Y4XG8H+XR9sRUITMDDKQ3+/iN
hWpErWmHKM0lyHcl5QaHhJJPK6nSA4hMEBv8NpxjJOkVBqLKK12o3Br4Iqk/
NTT6/vdP3+U9guxVogXTltZjHQJ9zrsVCr+WouH/qW/guZB6SEoH4Qjx305C
6US+hDoM7ywkHJqG5XwCqpfN9aAD/4gYcYa36D/28SP958TtE3GjTiLQXb1P
F2qnaNzkjh0EL0G/eda3FPmQV5w1SmRwErtwc07/596X0+tjSWKTsKNGBx5X
xpdFL8tcpQOmJUm4kr5w0M+un53ktLjEd3PhxLVK+Cdn6NHDJQHIpFOVFBvI
8fYJO5RQ98Oizp2MwCBVfIO9frZ7o5veHDxBFNdE7x6GRDsnPFO81Quqzswq
x2S68AocWeWSsoBlfGGrlbttYCqq2YVarwHfRKSbnlwihpbWt8c0RrXLzMLa
Khb8raJeUYYPlmCmPKtm0WsYLIuZ33C7LudVndS6+GZ1IjH90Rj6YLi7reYn
jtPYxJw43gR+gUcHIZaV/BEl9F19AOy1xtQ0Mr6fgYr/WRl986jueMC5aZB+
ZaWM6CBfSHhXaS8Y2LL5AkoVspcFoBecWuoyn6NyAPaO9FTu4kpvZK17Bxey
ytnJ6EcGX9Ct1Hoess3hFpnyLDVxmp65FRVUnnMy2wvIR400MXcYZyK5RMIc
XogiCFFQsqGvwD5BqSdsvoAFglkOoombMpN131g8hsKHTe0jfP7GHpVBweZx
A70vyrUUfnlkbnObrYaB7Rgcf7vJvNu9czJiXya05M1wywhngl4OWUJ1CWrT
7vVTLEQS6Yg1Zk3lbIYcrrkSJf3OHGs881JtRNVJGvg7kLf3rSMGgxjRC+bD
WHDJ7zomYw/557fKJYbtkglQZAehW0Zpv86Tql0rjJTa/vikvAflIzWfIFfb
kLvreuuLfv+x62n66eb3QxF1nPo6gTzvMs/7yqEqyLE6XP0nT0LZb+sJgXyi
NtRUsJssCs5rbnE8W6WEIfolznslzD1ZnlDoqASCW1YaZ/AQb9nuNnhZWWj8
zKEBkSVWRhNo1UPzUc2ITGuYd4ELGmsT+Bq6UgD3K4OrnJffDFIBV0jZg/g4
aATHI5EhcW6c4YOzYt/lRqpNkAx4pt/z+K2xYGByA/tLpgxuFNzFqG7Brff3
qnw7Y4Z7HCGWfW7IABxM4r6iT6V9jdrdncM4y8lhSMg5nc2BLrgAZr31DyFQ
4RUxJZNZPCi8mpYpIcjb8wH/jyU+BUVAGub9X0qddbGApJNcwQ8k2imPX63G
VWzwXX2HMLaPtuEVjWuX5odZ1GbyItcIISAaI75dVSie7gQeHpxPcYcywMfT
I/xLFJFtknu22CG1quArtgTPCFon+Q/z/exSiz7zyauIf6DumQwTDpN/4JIY
6Rly0bpTIlDluh2BVIrvirXMIhxGOKiASn+2942R8U/MnJz2U9RC7PwRUyeT
EGkCMJV8oZBUSchkiDmt0KMOsviuq4vovVNVmvvzyW/qsmclA2p9YKhKL0WP
LeOOxjyNjO8lmmt9YuywpUpWN5kgjPgxLrbZDOvWMYrJWUxehGGxd3Bpi5uK
VGFx5RYEbktBpdvjd38+4wbr9ogi8/wcTD8vnoPWg3GXbvxz+MJvp4nl7dpj
pCwOBinoiM1Oqk+1UhYhL8jsTEScW/Frjd9A+zh0qi5RPfld2xgQ7RdMNVVN
3h0lPzLHfU+G5hpuQFcJOZEZVbjunS6/bzzLAX3yyEUvKI3/jUmXdjQQmi4M
JCRCpHAiPb+KRpny5WGS39yAg1oBWW31trN0xevnGnNOVD91f1hy7TKcabcv
e1RfrqTB2rLYcl3kbucTlTPtBvR8/QzNRom852Q640bDg7VXTZUohT3A3cfe
eDaR5c4Lf3u/WepibagP5IVx6mvMV4ZOra+SYbg0rS0CK50fsWf+J2lj6g26
zlEYWbYxJ/Zg6/1fZPvRrBXEVUsaeqAU8HBaSKHAqSoAxc+JP1su/uCy7m+x
YkuhiqpKDJTP2jEDYm2nI/+UrHR8VUh0TeUCj0NKTTAOZgT9IA2zdq0u3p+U
eSJ8/1PXf2UZECiK8qnLqCtC1auyG7E4bd7mjitc+BHpzOkLUCriYKQjLTPs
VaEgAMo5LFshJEmBWgEcQMJUxZovZK/V15LJpur/GQJADT0wgE0D+2Tepeas
XOoA02/W/4/dTaIQwHtnsAaaeHR6XiGwHW0+4GP7P8UZSR7w8WhC9yYBn6n5
7OGdFEyo+NQQzwJz9W4lPMStG+Qua88w1gn0M/JM7p/C64uJXZXyUUImJzL/
SYPLM40p28CQuDelDXAYCsbaEGJ2H7WLOBkg6rp+xB3H5d7IOTlour0K7MnS
qJO1NqzonmiOpoGyF109/WXHTXWWCWNd7B3/AqBw7pm14CUs1MQOHLBLexRh
ltFsYpkj0vJ0b9JDe4kHb4DNqJ9X7N6bPzyn6LCc72tYZDp4Bj2MXcmWocEk
8vcbMa4FALVAIh26Pr1+Sfs8EGERg0p6JxEy9J2M9B8it8FUP8l48o0Jv7VN
VAYLn6ydIMWH/Hj2HwF5LiqSnMaxcWyvI2KKlPv7WZ9ZFjA9jGyGKXErS/Yb
91C2ZX4YeND/61+6bbagtitmhxCKqAdracqKbf3FeMtcTwtdMRSJekIfdxaE
/kMrNbFQEjKsrdpgWKiSYlFAi2T5zXkc/T+QJfO2FnGmqglpg/3AAJGrp0TJ
UWdTtxkOQYrD9Xt/1wcLrA+HvCqwdiPm8todNPg82u+/flUM7AIbCynSzhXu
ctfIktYwYgPpGZo2SU6xiWi3Y7JYJQB7+VTeDo9XHRREKqUmzXNvNRZugB35
FJNEemWZydDH+WMwM4E+uEPPGdvTCZNy3+TDEAPrdurZyYSKoGr0GkkTTwMD
+MEAKlIK5kcqEOwbnmkQyd6EPawm4q8GXg65nRfcJ+LiKum1m7DWRt4nXzNW
pnUGAixwjZxlfNFd0v5HVnk3aoxfQrogTwp2xvhJO/pY24CZrxwoVB3XfyX3
QIbVXBxOVSCK36LZTayhXrO3Ghl8af+IrqqUS1ahFDM7LUxZepT3BN8qKADE
6RC8j2LmK+qTVQx55y+nYsnmyc0+QGptji6xdDItH3hYYjMiH7m/AvjPyti2
Y5U3ReyFJ350caACtPS1JOVgluSJThL+uw0Vbg27yDp9eO4q7OH3jRDQfDi+
wufAmVIZTT6HfJVrmifErNV7V7i0oEh8xKpskoxoLSg7BgQYMWfwM6jgYj2I
ziJJpTCayi1GAOhiYK7cg8oSzIAxCQTNV2p/9n5buMLanhflBCe00Se4kYlZ
BXX2zDoLLhqmevLRm1KCFHg7/a5jNEqSbQGHbwXxUoF2L0w8gdJ1xtAw5pqG
+sfMQSVivOxzQWfP8trwF8djA6ksYmi+Gn4L+SB8CUATKK++ghgcZoT07vLT
jPFoMF904W8vzPM6mtbe90yve3BhvEM07KLtJdAjIZzHLyBVKvOSXLvYFMls
6pqmnsPGqmXOyWROvx5cXm4y/vNk6MrPrO4b4v9x2LsPOzk2okDp+MWAvKq8
7KOGaD3dfWlTqAyn3+DQuThBK76i6YmMBwl9Wakjrlnq/h9aXSeo39mfAzLy
vUzASS9OxPCw8cbfOjGDdcoLn9U4ymcDt/CH6oqN18etgxGE2dMsIl8h1zky
SXNFRhCSUwUJ+CO1q0qMhAbgcunPi2R7kKJhOxwxpyO0jNCXBCbISshUpv3G
LeRG6MkIc3+CFQ2igWrV13Q1ixlxDPjblAZJfQXPqn4pL2Iltxk3v8kyVVKd
x34QpAFRSm5/o1gvMH510FyXPPZvAxK+Sm5BrNpdy27cNN+PkwCN3qjs3ROt
sCF34xUyS8cuAe41HOFnincoMel2SLeJoAldUMbJ/S2iYUNmjXzlv3Za+buO
SoW8p2eTH3PD7BgeN2dozFCHIJoOfPI6dFVDTZpnAEfTkXYYNo4c6nLqODa+
hxzcJppNrEhLqZDbfO0Qg6YSx/2r99kjd4g6yN+moz9sQYh/YSqoyjLNYz5i
9Em/Ag8/3L8zNvOyvLHqbzpdUDNWG4MsrR6Ej4quWv1fordWCdi4wGEPoHKL
MAK9CTTgoRnOEh9qgnGxh+tIYKHY+MhzSB6RN+mQocib4yso/fSfX+oTidNa
UBcltS2dRIPPnnj7exkZqBh8l1UJFcFbRKFiCnLgbbm5micTmGG3aEwwOreZ
i2nBjmXCisDhBIdfOLNA6t5kvM/wW132zPrV7yeYGy81xOBv5Z7vB6VU0nHH
71RLI6x1YDusxPSxOEoK0wUotJr+l5a49a7xM9Cm4uTVkEm/VH5ZW+wBCkod
MvkOuGX0CuVVf6M4w6YC2MeKUYwLDH74CTuJDkLyqrd7/HZDQ/l9ao6eky1k
8citLvXatNmfTlJ5hOPVhmOokv3dmYlabT01QxTkJPO2OtA4/pALjDUQXNGB
oSUKfg3/q2GSWgIXBTVWydxWz4DdvkbPqr2dUctH3I8nMv2AVA+6ZrJAhnw2
dD7tRx1CkPVatrgMR5YGXVLfUvddVZ+g2fx1VuWORtiPkKxoGEUexBlo4TVn
xwtD6cK9fOg5DbEhWqW4Ba4LoAVueSWdHenpBNiFkB/KCRctvDfb6lYuJvpU
t5HlRicWDAhjSOI6n/zjdYmTXS1lqqgPbH/KrnQXty5hy/S5N0kOHRmhkeeo
eWff00j2wyNlVRaJcZ81WfU8SPY/X0MdqbMaXo0AKBMovvzrriNVqU27+xUQ
9KCVsyYL8HnsfkLH7PNhMZvGzDMs6Vvk9KAKjkbX6GHp6cDcULUII++XBsLM
gsES6JKAmuPCZKPlKPlDDkV4kUBFvBIHd4GCDjYU6tgL4J+ZL7KCF80/Mvah
dqYF7Tsec6vDxvodwsES+ygiD2Qfy016rdLfNXV5lSjrzdmHrDtRjvkZ9EMX
yTxIuD2F1whhn+YqM7hXshnpnUC1lqBFSU6yp+FiDNmmaJbUxbarjMZtJx6R
zdmBEI0hvnCFrS1nhHb4y2TqJgPrC39CAh4yt1U87WoRYPGb3C2knAT8+rP6
e7RYnxSPTFsw1ezC95xOD/vugsxpWff2/TlTWDbcF7GGLlv16u/dcBT2zByg
T5kXYxx/PJ9KwxrkTEddamhe11FoAi8u7SL7YCpidGXu/I7+uN+FTOEitJFJ
ruqNabDvjwYu2UMPJK/SYQ9UuzDpyLof18FUiI0aMeKDt6g/U0yjopR92DZP
tgjJGkwpk205mryTm5/myJV7qU3NX6uCkxROu+DIiTwK0c2c7jItTFLmBDJ5
wzFX1uZq2XMoS3WtZxYXMjcwxfjr9u0kSfCFvIoIaFrAv+ApHLIvOIrHihmi
C23xrR0RuEJ4z4PceT6BYkaF5HT6UQeb156EJjHTybYpqGYip6z0dbXVOBLG
/jSjoRWh1coGsRfUeU+jAIJv3rVXIYiyJ+cuoRiR8mW3yLIiEajCsB9oJL2+
09unesIPTzG0COCVUpe+rl9dyfZJqOOjb6g3dTTpb8RntEmn8O+bJPcfIxwv
T+A7DB8ca+vlYe7eDY+pv7jqhH+cKJK6ZT1/CBNRYHRFbP1vrQ3fEvIGOPa8
jlyegK563mOZ9ld4MwxCQAZ09A20MX/ojH/o3HANjGQBGnhFzke1TLGBTOUq
ZMB+xsS8kty1xDQg928F4mD8Vi28f+IIwvTGGOkxsV6cgKDUxu/vGdf+6zAF
t2W4+vdf78UbhHnz9nhC3wBYGYuj1yzxAjmKsOiNQV4MYyHmKHhUmA32146O
nxqaaJg7fj8KABbCR1l3rbc+4kCDmXBqqdBxE2mRseBQS+Zgr0GRRfZE4FV1
0nPL6jM3ZLC0E1BOuAw99hZFtIf4Cr8I5HuYxSWfRohU2G7Gw09rV82F88gd
IK3Gv8ZAWVKtFKQzgIzecKOkgNi2w5hu6leg3TGgcO3xQiJuSpR5l/uLi1kM
72Ia+FKsS1uxp9/Lap6nIuD8Fu6rPWWhf3709yYMG9MuUYCJpi6MLf2JnVtE
T2/6KnyPJKWy4/wgmvIldACBG6PIRVejomXDOd4eY9BUN6Q2ADIWA54kA/sv
r4ePqX41hBMQjB0cTkdo5xx1wZ425WH+8Uu41USn1u00rFqcMd7iVn1OUhPO
U05NWNCZljuFcxIRgJoKLHJwNuWqBV7WqReayiQzDmoo9aOAU9RjBLHu0bbI
/dD92Hd80RlW7V+VCdv1RAvG+K5e+paEK1F+qTyF2Z+adFZtZmo1C4On6Yye
6ZgA96EaLftihl4BCha/H+fYSxhSefSOD2J9EOcq3oiAPNbxyZQdJP35FL6n
X26Yjp19NeV5TRP85niQc+ApVKJDGBTxXdeNj7OXeH5Ajc50HbgGbr2vTsJK
RxXcbscE+52ZfzlMxXGB2IGSMLJjSBtMdFZwVU6E/LAIK7wCwxFNb1inx049
Gg93yoNKFkPD97ooGC/XOdbGrXEfcgml4dOnPtJS4K9n5KG7McB/9Y0FZdR8
3LUndWGOcEjO1cdy5sgDq7HLu1xG9U5GtxJgIljSSw7uNyVOsSJr0hMVjNO8
xn3C5/nYGgzQ9ecHeivXj8a3lqTfT7M4LPYxNQS8kdjvjjSnCeFRsECPu63c
T4C0NK5fdEP7xXKgYcdx4Kh9cGdUpAdEH1SaQuusI0+Y3ALUAB/3JoXXGiZC
huKCXNXrHqOW+JITGVqC9Uv1sKRHGWa8v2Clo0qbquea2Arnb3VLZb7v5nRq
aoRHhyANa/o9oApGAzigZSglzSr7sSLNqBvIIjE3PWKWEs2Dm3jKvKVTS+2N
7i7rMs0aLyvmFnjJldw6Q+yONBVCySICHVENIOrLukunr2ZeN0CJ9fYU3O4w
8M2wZhTyy5ybF5+7ZtQEsw+R3yxPmmUpkeYunslRNAE4gi8saChscFKO1K8u
JtukgUWjJ+zY9xlCUSfHnJ+tWzzjeYVLix4fBvyGHLH5Sds8oh0l9UJefHXe
j2VP4wBosvaP2+lBNb0/iXuXgQRySag3E+KdyGDsV1fgb1IFdnhrAvhaHuL0
9EOZOxgVPFhGE1RG1hrClVl6FBhtDtk+dWHwllnkO8Gm/Yw02lrevRJGD73I
T+yKqAwK6QxhTYAqFVx7cwxHafRblcB8zvCHpRfjdyG55OlKCY+DkjY91Dns
NU8+uYLQmdK0YgSXzmtia1g26qbxY9K2u7TqnueAWxOEiR2uk5H+n4Wi6Sjl
TydAB6N6AYB2wt9aOgSIIgQZmv0N1SHIyAuMm/ptEbmBOFzfaVq46On/nG6+
1f4BdtoiLVYrnm5T62EzO6L5R33rU8dZN0Qy4QIc1fM2gdVrhTwsaRpcmooL
Kw/g8E4+Cge9wclqwesDkIirREIU5nk+L9VaTKR0bZBjLbmhXgt844RRTUk0
Nvu2SjlLfVZHLwe1D/qt2skVNOsQQGtcmAfmdwhlWjedd9RdBvkLxhd+0qXO
BBg7cXDHP9+xNbL9jfr3ZYHVgRH1jyNUioKNYS6/9XzcjDxJttPp8VWt+Ilq
00K1H5THs2Zc9mKYmkH7PmKrDOuzxw0p+y1/jyjZw0j1ZCUpX6QhnVEDhQra
g98xzrDlJM15am3fPYOrBm291qrLCdG8qwS0B9mHtnLEsn00upoE/igYAhlV
rHrNjKavNZ2bszzN16JxCgAQI9TBqZXUPJKUddxG1you5VUfCf76DpwkqrMT
n9yu7bgfI6LSYzjWgHCu0cQUWRgP+Fmg1avVZ9m/PTCgy995i4QdZ3L9++kJ
TcBSdxbVd+MzaC/irxw8b43Yzw3h/eWR58OdWeGgHbBpUu7nXJ1jRzyQUotD
/A3wyvO3znru+pz/wZXMacUVIPEezRaeepTJ1y24Vy6FDSjT6WpVq6Obj/6x
ntCwnzR/mKjOhw2P/ZnZpYtLZPwBmcZAR+Cz6LGU9Ipld2bKZM6ZpLHtKLIZ
eZo7ZUrhoN7Lp8CO3KdEB9HUG2Eiefhsva3djNpr5FFjFIN2+1jWiFYmFk0z
UuGCPf4MJ5jPdFjc4D0GpzresVywWm9iSr6GE66KpHMoeD6OfS3BE9ZSrw6w
/7hxfRThaCZww6enU4gHJr+yRa3LQ1NIbjJdBrowaUFSqJw6WhWpL0obfSXH
ymGTI/jc8ROdt3lbojvtdyx6CTgHXldGQqTaI5jgRto2Eoqp6IErMj2xOOsL
PLN2Oi9Rd/P4jj9IlvGgDo+bfMlbiMESkLjZBDYuCsYRra73VY980wfXuiLB
v1EyDkGdsatpZ0oIcY6hRKhfWu+VhpztHcIHD0/+sTJbmFybSSM7XV/patl+
7vAdGFZ9DeRXyLhewLLgFEbqfYXecub0zQJbsiIVyUneFq7aY8Fl0cIMJzlT
AcpvQypttirtF3j36lZbs5M609L5zk7SVpXSISz2svosjxbQQ/IT3SpWkxxl
JCKH8e34+isr4OmW7jYo0gSdNkCgE0gaAHnVjE4RM98KaiNWBRG/onoZu9SO
+TUJ/MTZkfU2fcQgXsez+Jmkm+LUAbeHNIQpCq19chTB+Ydt6fiUSLA/BR0q
KcmkyUXbWLHBkG51WinV1z9NkdN5LTUSjheirVnotYDPjYNIFDbSt/cT4ech
9iGFg+l5zlwNRlJhZdeP1KaeL3vMvzS/dVdPcsT+xdQ/J0u6wyzvS6/+oQFg
uNuT5i4ulcsq+Ie34wcLrg1f7pOFrJozbHsdmos8tat297h3ePiFyBxLxGTq
3M7jwOQ8ptPvqjuD7dKFdEBpIeUY/ZnmptT7Hc0ZC3x4rM8Nkc9pCga31tnQ
VPSD1Pe63lKLgEST2X5F0cCnFNiNF1UBuWgzIib48SVROP11TXySFo+8xmLw
m+Yws99yRvkf8iPZr3n/vQVvk7zZBqEmstg7lTc+QdenYLYBsUG0FptGvG84
58JI3lwSyfkxvZ4J/vZgXN/rQgrdTeEmlQaHW2IXh2SH1AsId0oIcOAE7YOo
CklCwjeB1p7h9t4UhSrUfDW/ST6618xRbtlJGiIEBmFKQqDUCigIBYTVQhFZ
JveT/XJ/Ubx9au9VifUmlK6C/QfP16fitqF5HX+d4wtSP3AoEXQwqVLauJVz
0xl8hjzIH1RLSTwPEXtm7jKJA70WhF5hdRLvgY0/qF3PrB/2lrCgAX92my6z
Mshj/+h89avP7xS34S7/v1SJnjbBvIFBbXEP9SMyejMm4eJ7K7Z37/w9u6C1
UplQcOJKoc2DWTu3hPqim2hLgelFWZorkWvxBCvJySf9UurbD9v56Xg2gR8o
ELRNFZu8UTqhAD9PFeNM7rSMf/eIi98IIyx7bFzQuL8OwJb0QS2HhkNugF5A
GoA6aS5R5GNNfzQ06NcS+rWpWBQa+HZmLGrXUY7TXKzggfPbJP5f/6KDiAAK
rEcND6e2s5oO8sw8wUYQ8oX5RIEvsxplAzVbIcvivsmj/B7/kpKCQccn/9Qj
YfROolh1E5PI+b3EmHjMmHe3LBvS2nxd0qe3NniCsQCjly790mmVR4Zykuur
RXtOJyuho61tXsk4L/KLBgoFKyzk9pMOHx/JF61ZbS0LWQbmn3opbZqd4bdb
B/HKvRl0JkU4jdQOyN/1HbFJFJsBEjzpjYFyP3hcOB5utKnFaU826Sfpx/Kk
IcrxfbbsFQwcxhPxEV4jpkY04dBWSndgqOQlvdjrYrf87aGQ4QN0KyragY/m
W13LsEuGTDsQ2RRzYTttZLfgP1mkxOSC8NI+WiCKLBM0GXhbfm9Rf2Gc2t+7
5L51pyh6vyXEGgDHs4Ivg2biTjeQFA2yE+wyox7ewMf1vqVZ+yDUlGo7PBUg
kE6Wg9VePv/i63bYyC0wK4W7NxISbeb/+VwmvY4z0v0OywxPIGk1d0HGG5ch
hI/Tzw4K2MMkQaSOpwwvmbKhpZQVAOXPaN5n3+w0R8PddFOMr772GPJ5qXKx
IQM/uZU6Wv+v8KBmkcwjNHPeyUuN+G2mmVa/ELwY9k8CAbNKcmEA3bsr3Jwc
loqZj9lkqk2FobzSA4+YbjavQ+2ZM0LQcM/VqkjILPeYzWs+QOfrTi5lSw0J
w35sycAFkBSGjA32w4fQO8YhFlML7i3onfJlIAz7sYlzh+NXWH2JaEPV52Ri
V0xeaTgE9eDiHg6X/XCPaYDklClTB4tBgfhleMVQpbjVxGOoxaiXfB2K9Ujm
7L1kHZoNwF4YSmudazA56Qd5w4zfGnAs6wmfHPYYVuBCZIJRRtJgwL1BhDUn
iFw6gWxd+pRpG3S5xGbv+czgcAp8QBJCGQfgJYLDfrWSTfif4M1+xawOc5Wx
r7uR1CilGBAV0WyQ/I2u+iumyUcB8nhLFKfTBJ8g4qxyU/53MbSvhrAhA49Q
ynaj3Pmy7cbYC/8g0UPiK7VGcXdefXDrvDwrXZpa6So09OzHcPI6/cK3OE6z
MXeQpmjFM+QLMjug3J4ZnfHW9szV6q5edU9X+sUB+C/26vAmpTVM02PIAEMa
Znphg/8LyIHHP3h75O6+ffI6/Drl+8SRjZoyPvXKY4lJTALexsdz+5pH3lxh
wo7m0/SmIIOuJYEhi9IGEJd2xI1otpkVYg95UFomfLxxFYU0eKV9QDZ5h9l3
eB+qAHcz98SnebNzbZuD04pdZQm6MOE9c3cE5D+nktbs3RTtyBc2sqoP8B0R
nFziBL8b9reHy5gj57xh63DQerwW/46y2Cmb8Z+Z5xybE7uuHYqMsllfLH2f
j0I/wJiHX/8wgf/Ro6x5acs/VAMocvuwt2Y0n3ZSVMm52Me4uSPsH7kFRn+V
JzTHA2RUYCR2l1pn+9CrLCIVDNCUlUiHRlQ3MiMbU6C5T9b44/8LY7m1/nEz
pU8Ny8YLhCdvUt8U66t8RnY/Xqq+m4lJNrZsj2VB0Nu/tpH9dsh9/cLlqvYc
YwiZ8iE+sBAtCSEt/A2L83vh2LlCM6BMDivRM/QB76ZJXr1qcQ2EHrnaKxm1
DkUmTF3yWnmGAdidO0Q3biWsBgELVAI2JeTd8CYlOiVBq1QWyWi6kv8rWYzp
kv66BDt3CMfC54kfx3TyL0u14/lQ37ce3GFEdCoUWqvBQFHR8tnUt14Xl9PY
gxxMOICJoJIPZ8scjhJBkLe3mFieMYpFVCd+AqwCDDWig4rLuQMmK2F6UHuI
edafN13rfVggOCRez8REk8FQahbmJVFPZj4SBeefTQwrUB2XszEyXawzQbTE
C1nNHo5daptokpGZIKFdtfRZr9C1UsosOd1GNjri/Z4gGGtuscLcMfq6x/6M
wbwWlZH98ro+r9jOPYuqGHI4mJLGFRX8pMg2uC47rG3AvSoXKDS6cYy+Qc50
i19dm3DTQtcQeItnJ6T617JJD899t6uy99QTCUvZgNLDNCzStu4/6gAGCjyf
NkGFROljo50J8LZGHMZzoYiiHok2IB0MW9cF+nqHgQ8oixboKYhvurJBAxB8
bT++XtHWZQsWKYgksTp9pkh5fC9pe80PYkx2ok50bBJlp0q5WJh6wl6/wNLo
Tkk+0tcvv+mrNld7ujLzZ7QbSO2ZvnjBIocLdOI36fCeK7zX+2PqrOE8OD3f
vnEDMOiiYlrxo4DHeYNgJJ13bpZdiA7u7FKOFNNDfwp/tle6ANd1sggjMY9M
zxik7N3PXaArMO2MHcM5d1q8VDodpZzonEY1YYFAC+OkekbcA/8v2diFZ1pl
2PdK80P5vtIXMJCEqtz0pyxzIU5mGBC/oKgPuxgiDqY+VttDwWDzlqbgBS3t
o84v+FC/P4bqLydj4tBGEKSRx7VcMtvBERKb25S+EbGkYLEjx83pKfel8SZw
PeeoFVi8ygcBQy5mSS0/OLaQWKr7KUhCPFbtNcTEyuAQqjZPbcJPuTwJW77h
piK782rsqMQdGdpu+ISTjsNU9IQSn1Hgq0nbCxWoqd8zihIn10fd9xIFMdda
SjRSlLhjcWol79h0daY6oOQD/G5aRHN9L8hSgytW3YPwrexanDsv30qJLcgQ
gWlbYQZyZTYzcna8iT1IOCTdeIDLIISfXCETN8NEBANxl+Lm6KrUDMfdXC+8
vdTMPDPovDS0glCmjrD452iAflBM06A5V8DpsMQq63ILtl6bQvKp99KmDN98
vvqK+jUHN4D/lBg5XCmXdFiIhD+1MPzoinh6cZwvAOXXxUDmL3jlQ+EyqNl2
vEgA8GkGbWONrmhW4EM/ckFNHb7QlH8i/e9VhkaO5qZ2Vd6Ej4jixuq94yW0
VMTSYhINVTkE8e10G0YVjDRkYN3kBwUsLc4nMoFNpRioLejfFoexFOoFf7Ux
XkxSa3XU3yzE3DVUdha5fO7xqs98tHIgATpECANO+ZUU5PA+W46uiTRXemz9
IYg0wjceLqwYjsUWkysIJrqKmdKGuR+83spVu8d2EBEedthYUIdlUJ0XAiHh
dKobtpvPEzEiVNYPUp8eosavlYiHTypQ5t88VZGmC0kwgbnftxriC+vfkMlJ
mMiapdQAJaDPyaBVJkTgn45LA6RQ9Gt4oyUMLu0jCqzx7RNMyKrW227+zZev
y4f9tVfJSVLogTihWAC140RB0v1x9CBRJ3qFQtrXnmzBBLqfphuS9KAYVAKy
ypsi2J0dilDlZo9IDNy8PVj7NW6QW1yUMqxsI53/8BsmnZHJBO18iaXMIAwh
ipqfOlUqkE3j7BfVSinupvRuhPzr5R6gg0W55+KPwGr6EOTRbRltg2frz1km
6DPq3ACg3ryYc0nC5MW3rVnNw2AkeKrNozdlIukUK0KXlDoZj0ifOdKV2oCG
/dj75epwdTi7yAgR5bKI29U6Ri2WFJ5rj/n5xZVxhupLty6Gs5AzztcRqtP2
hmPc3BhZtGjtYa02KaBf0SF1ghaWbgNr08VfyLW289m6AmlaYNc/0ldqmzLR
leECudCn6wGFPPB/Vh3Z6seH/YrcxXfbLVSvRTgBnmpzVPJf1SNTPa9QQRq0
F4Tjq6vuZUx/IGhtuYacoLXLlcuI1QVtwQ/3VBgoJJ8TAxAoNxBpw0THxBIY
OqMQLG9PnvNqT4+MLuGjPFYl2Iif5LV1NB20futxVAx9SD6hKSrm3tCHBBMs
XbJ66AQa5SxWxCMTWb0iw+rkj1+jwE31BOYHue+89S5TBjXK2xRD38dcs8oN
XyEFaBjLuBXDLAnAvzADTMb7R4Wu8jdAfQj04YiQG9AgENGIfm59cRF4996b
f1HyY7hnaeOwhBsM81pD8rBeoRPXypwco22c4C0gFKrSEL/WX40cVHoDmW4F
lOZjFLi2i7Ndvpmsly9UB1WuxBomJFNYYoDBV/z4AyeZdbKmoDjH1orP0SZ1
/tWjD/++nDqEzTTKXqDB5sF+gBkQnclWLPK7i1QbRnDGsWSOT6wDq1oBSmF5
i248iBWdXK7OKxV5CwJCOhz2wC92HSKsuSYWfItzu7eYEVNzOleNYpaGnaY6
IdkzHmKPZ7DR4A7dXMYFAFOrUg8mO1Yk9Hm2fJ28UFM7Bsf5Oa5DANSaNfA4
NPXdvWeLyDq3McHcDjThzy+G5UwNFg7pZhye7wmh+p/n8JD6rQZw8+oeVDfl
Csfw6MsAUyokabX1IwMiFKcVTQr6ECvXv9UYQ4UT0PPSfKx1S0gEfwPmnsuk
h9exuNwRx2dJ+JqEbZtp1DKvovn2Gc2+2AYSsPMOh47wqm5U/bJgJqd/Wh6C
RwwqF5bol0gJK/b0HIuc6gCtkCtA8d0n2nzw+1lhkcEaaGM3ZHmUQKWTqQrG
a8U2ejPqrTqG9/evwsOEshRePIMcZIA5p7AhKWFXBiSbHRa+UDz+dhfqpD8p
C8GgqrS78rUyCArqliqIJsF0/kuumJnnQbZQS5DzOghXIEI8QELY+vVF+YIq
ynaLigOFw5xCjGgihNdYDqhuRAgmzIQIeDzCNVFPRNj/IAsFI79L7emeSQ2t
jYt20QN9aZxeYRIlLAIIb1PraLOWMQOG1dDXrRHkncdPxxoXzPrEPU5kJUsD
4jBMCJkAoOoUmtRofaaMITD5E/+bTFeKMNNdrnAAMu0el2ww3232nypHxJAr
3Iau4P1cGOmr72cNeolUtF5pgnZi4G95EVC4A7396HgAxXaFm9yBytod2UMX
Jq7JuT0J8lyS6jV/N7cFWp1CwpNO35sI3lSl1iMt7lil2sJvOxlwnApsVub+
rv4lQwKTZWr/j606ymGpomQyhxLP9+DMMp55Ba1sA6L3sOHs0xU5S/1PUMXk
XEsAOYhVFeLMP8tS2Adnz/0UGpaZYiXo4DbleqEaFK/p6i2CGmvxHDDADjHV
fFhovyvnBWxWoH9dFby9Gz9dgytVHqhBz5IAGePfZUhthOkXXEVat7sM8xnn
tMGPBCO3eKLfy8EQzPaSXBXewoha/rya7f5Yc8EyXR36SyYugwH97H+zKL7r
NBwohvH3hDXLhAWNGVy7uz5z62iAxWB74Py/q+9cYKckNeIEjWKPZqJ0LKxy
0bYZaS9MkheJcSowuF5HoJJGijdppjJRMDCGxb/ci0bWJmiuG1ZtIzOaBnqL
vSsxx57kjjMHalEcfiKi1DopKblNzIJDA+7eOkFAhhy5Es33ZiQ3l/DmKbAX
fwT0zOu0ms/sbgEofEN0saAJTj3pOVzpC2ttYpRdJMZZKhyFzhAp9zH9N//j
nHMuKOKSWO6uhNC2ivG+xF4VoFj3uRWfAsm7M45oRQrdOmi+X8PGnO5blgIC
5IWYOfBMzYyMtKfqw62ndXC1TAVWy5bFFQ+C/klKMxAPJIb48FkDB90CwjXm
FfLVmYcwbeo0y5aUqoFbcOE9OiuTNLiKXWw/dMzfdnWvg3yerTq+OodVTRbJ
bF8rIby5/ToIHONMOoipd0kOajWTaBph2ql0JJn0MUbm/As/wlL0tsOrYVc2
BKohXxXu+fQ5esEamPG8LQziK4NVe4r0/YCguvJ206E8wMLCOy2VHSY8vYSy
VMa4Gr5uFUr7I7QOaEAejTILxTbwGaYMh2ZzfKV+8fYbvXT72uOAArrMSqQu
qAtKWe6m7ArrjxPLn2wxjI7UcZ07b67cXnJIA21lwMsaVQ7g2AgtS8mcmQq6
SCaXT2UaX9rvXX5O58kho9BD0jMbODUxXMwZ5r1HciNldCU9ZicNsVTAArUM
VgZKk4moM9L/qJ20GNxgHZQfmK9rwTveq/8IDkZTsTXTS3StxyOAxKyQdmaP
XjcYmMNtdLzFZbsPDjO94CLc1AcxoSBoVtS3AaHYL3VuKoEoHr7g1Xn2886Q
/tHDasLA98xFVXps2q1IJA3hEunUiokdxL5n02cSdIdnZz1MNOLGOX+PkAH6
n0wRyhYx9Dyi9hVMEkny8uQ/JmShmiHHlKzRxyN0klrKArG2HxNJSS7m8v2g
u4utfkWqWTmfzbiRMfnnhfYel2+iU+smDiWPyK2XbsYg2ysfF1J14NYlWZQ/
uBe0SKtZ49l5Uu/GyQjEe6NXFtejL27luFs5e5reX1w4ZHWHyp0+eW+s7Azp
kgBsD9Cne0twWGkrruJWJ9a1I7JAgBbypsG9nyiOQIWVcSrXT/834ueWCvm+
dvYfl4prdo9TYb08yTmhNbn2+SeAtXPzA9xErrhc0NqhNBL9L+yQ3kvHg1M7
qSKr+VXjgItb0RDQwnWnL95k/r+X+BkeLvBD84bYYouPxZ2kOLV91K3XCKU+
NpSe8VwNHdNRFEbWkgPFx80LA+pihYyYdjC6VSApDeiD0YHvm3NY8Q6ZazRz
A1ECIt7Ps2hRrNUOqLu+kkYh35rQ2xflm+LrV5kFDJWgif2KbwOcWep7wpDy
Nfq3VyzACWaD5PH/FgGYYZE5hvJttBVZMfO0J8h3fwH+sST7VfBkgAWdXDJL
dROvZdkaVFrYA9+048Pmgv3xPJjre6ULHHuWxI5rfLPUcgi3uEnFzyquURFE
tAR9Gpqzlvdro/3x7qOfAyVc9FXxzBWnWBaJZQY6+jVr/b4Vc8whQMj/tZ8+
PbB0yQK+qjiu/OF8CQW5JIaO8oLv/fYilhnhI/ToZ1+8yQT6Vbpm8h3GwkQ5
/MQlrVaE5dc3Sk0iLvFjZKbkLQ59OqmRhaMK3TxUGODZgNz8UcC1WyPqmLYP
w8lyVSztBg1NnVqIR5wEg7E95gZtn8B18cFnmGxLAJtxRB6UTHUJprwUFhDn
cMqy9SABUZUd+trGFnTPiD+LjP5CZ0+ujEZKYVqF8tWg8Nsv6KnqUU6F6c2H
GQbz5TRAV96NNB2IhwfsPFkDrlwnCRoqg1boP8AnxsxyUG7w0R9ApuA5gBIX
yFiplHnsBnVRs6kdUkr2xpfL5ZOQ9q9YbDNObmj4Up6i7IdxgTHXg54TKQxF
47RCuOZI7rgbX/PKlAxDOPS3ywcyjeSOdLBHUfoj2UM6Q9v+4ROVRe4EPJ4R
Kn86YCUSVCyaLHiKsGJGHlNUAq5r94rKriVMO5relPaCx70nd0yWBvBk3/Uu
Rad76kvY2uRWMsufgP4Cfmiwiv8dYt/bs/MFLT2oetGOIbd0JedsMxJwTpKj
hYGAKCk3GVKfrSjOCsXnUCZnU1t6kB9oQ1eKujCHTqxEmbW/esYMCNmS1seF
BCPe3LDaVcPUFPErDZA5FIrm/S5JCMyfnrvlL40O2cOiN9ctANMr2+t1l8y7
6pmF4rw3PFYJb9wJ8+7bp7CDR+Sa1nsGblDduXiUvtJYFoyVJrAG7oyjc+lX
DK0wWJTJuyM7aszzWvma5OK8WgpJasR1B7QINkKyTdqMHKmuIEQhoJYM/H62
RRImoErsk7OOEUdbs4fA0dle7KS9EVdXw6fX/olXQ+B9ScbwWW9PtgUO+u4K
Nb2IYnRJBEn+Msgy1wGS3AZ0P/uq9AIiutDYBOGv4XtRpKkD4GpKAKNDFPlB
xy7oYy9ggPMGu/EAmS1GzR24wpbd8gdUvAxnhhY7UFfqXkIcfkM9xDiYyx3D
bySEBdiE9YA4rDJnDwVyBdA0A7FjXhVzTUG7UwliYb9xHRv3HxbsrsnLpOLe
/StuUWxA0f9FyOVQrLMdPK/hxZoxjcQT47unbqt2Q3MNUJ6oarYQRpzhmsUT
xWqv3GH9USomLHIgoVNvrlBcvJ6W6Gy0h7mNlv//4vA5z80zB1f8imF+/r2U
7iZeqXNSF7Vuw6XSEv/wjZgK85vVQMulB1vqoV9DsRE0ZsYQKXA9VaKk7Rqn
1owjtjrb+7Y3LXQbXlS3jBFvuZDwong+Vr+KH92BiOBEtJZIA55c/3YKRq40
nJMlTi8uTJNVsRSfe+H70sU6b8BvQPSNiq9lPt+mltOK+k4V512KM3P3u9/p
RZldIvCoHF3DfxOGm2JJnom04J3ZRZj1j6CBAjq+yEV+bRUY46pvUqSnZGNV
gMaR218cMEK1mkG6x3L5eAYcpd46JsfqSlQgoAD4C0sGkTIM2jGDpt91aFkd
j2yPCC9qWuEoBVJwwHpGnFA3R5kUAHwMLWYZRla2ptBTSGw4KK1GRjAmchXD
UgD4nZY5w9wooYuWNbCWlrLsWKKv8ZohXydQeq3b3bivZqx33yAjKtcp/j4T
R7stSE8gqpc3tuvbixg6nUFjH9Sh2NRAq0VTlh4sF7txWkuCsxbYocm15EfN
SBOpyeZ+HddXcW8zaiT4jw4U6FwvH5ZZmrEjff8m4A8SLPjQbdVq2qnqfFcf
dGlXzxjoRhmGOOxg+nXRbNgnrA8+TeGhnX72uTrBql70uhbsTn1ZDGHTlWmX
7Eia2RU2h0UkMkoLHt2tNe+RkbWU+jJqItCKgLJ5IiJAbz42LuPZaZNvA3Qu
dKypUd1X8Yb3hyHO18852DfAKTHCELo5giFjhPF2j29FF0D5t+f9X2GEtMR9
6zosKMYzZJRu1M3tVb6ycwhE1KBCCiB46HhvCSd0omPx5ww5hoYG8hqdDCdl
w6ypZ6ZAzimC064y9xrD7KFFR2x79/SnMOrd7zvfEgiluyJr9IvEa5QP6M0e
7OCu5/ZdMjRMa/9iikMgkzNfgV//7FLpdh7BhuW+xw73zk5yG/cEU4Uj8w7f
kstQcOgY0AI0pBB6s4LFE2JlghUGnQ2lcAuRYC3tp+Y5x00e+CCMMEfyC1eb
0FSoUf77kYiZt2Ueo4dsxeini5ulTMNiQCze8VyubeBdScNVpSqMTpoDpjBA
xm+a4cSFcXGiQabY4ZZUdJLljAkoSAx+VJ0aPef6HpTMUCo6L/HWFJLRvZ5P
uJEQCbq7nK1QZkAwNgflxwHr31lG46GjZ2/Lg6JROTs2cVfscbL5CW1L2ODo
udWrA416tErVm8u+Y1aZMrDqInIJqfjcqUQqmOD8en/hN5Ak5XTZDiDFL+1X
jz98U8LYzD6lJbpb7tq5gagdtOZV/PgZcq1XORgYt+R/pfAs+Pgg/LMwpeYg
Cg8OiCEei8vMEZ7VqRVwOR+/97cTacCsXlnSoZo9bK5hHUgE6Fb65mxDBw59
VzF+y8RuYtdNiSZD3yoKAaw3m3udwhUD5F4XFDH5FAnidZTv1pHlIkXMEh67
0sb1kPjUe5wD4T/fKiGOrP7i/fiTXS2CuOGN9xzibkppaVXrvuoB0xINdaf5
o6o9JX+5VY1prwo7HO9Ujc54htBgRR10PQ0hugVOhdg8r9EITkKZg3CyhdUU
ta1p7pYtgCQS2tp2dcI93ZgENPj6SQv7LPSpZ8iohvG9Re2qIO7IXxYENpqS
Y3NQJXDdpllAAQdx4bQpyjv+3vrXB0G5clWh1A2BoNCOWtfJO9O5KnZ44i2G
tvy2YPlIfRqYoZgEhoiXz0Y8tPBM76mmHP36Qhhx9KCsV7wHbxEYRWcTesr4
kie2ptt9eRO0Eh5CesoSZyw2C33nbJjtdBXHavuCQhi6fm1g+vgREpf1vytH
a5KHX389xNYsULEBAF6Nkt7ITIc8Z4+V5aXlkDBDGE2s7ncBto6kXuX4sYbf
DjBDndEZgyVzieaTRsdaW4/nx7RPIfx5wQ1hZxvjlRduy9S7Znj8yxsNdpFa
1KxRLtS8UnlOiUW/HaeEm2g8ZonwBsuMpyIn2Nc7+zl2NaF+TNuiMmjWOc04
u2cbGlgax2K7XtjC4sqsLtVK9H5qFpUovLpkhCZIZ39SYSuKipkYQLollgnn
Lz8ysfdISwui/lsciI7y65J/gFhxLPlMpN0aHmpvmWyHCHxVs36RHNLUeKA8
siU1/cGQ0lDuzNIzi34/VEEERWHUcbgosAjFC2+g8SPoPxQkYQiw+N7TF29K
9QG/7rC6Kt7NGrFB+1lkI0Krt4mqzZ7K+QzaJcEVOcsMcDeZXGpfUf0b+HB9
2fkkevL+6FyZEst5eh95E94yLAKk+CqA6VVw+vQOgrn/nWakPC701lhB9nmg
FH6GTaAKTIkLlTGSfYjKE7LbfN5l7Q71zbfqqbzmXKRziX3lOB+7g8S68Qso
BJ/9zmUzE3y79I2bIUG+g+ExNnv5ov7HGGf715rRHn05ystH1XsSs78MHBqK
gsp7nxroG8DcIskdEt83Nk06Yu+hP+VdV13tfVJQSq8UWfXpkAGrxhxfhQ/M
/YSkwbivxJ8OiBoPmNDbIMO/GvJp+R1IWdkuMb+ku6iXMz704rkNftBtzVP7
z1MmEAMO3UbyH1qtSNPAg7iHtHoKzWREjqBEyEq+0CEwclwL86GcwWRap1ZO
uKFXOVHEoIMqUvdySCtJ/y0hzqVsLWUbNsl1s3hOV2eWjgaVM338OOPLt+Yj
4hiVf19ilOd8oqNAwAwVO+bCO9emx9wmVczk3BeDJFl8ukUkQi90C0i0VjPh
5fYAcrzXDYuwRWkjbbbfkLCw7a+ug84uZRTia9Vc+LdI1S5FpEMYu1oLt9Uh
X4am3BORqR/LPZ0iobTYvS5+Xv2G0GgkleqHYTxLz66DKIag7O/Kk6sFVEul
ipkjeW5vAR86phGfn2trYhuOsJ941vIH7Slvdbk4RFohCHf7BTturi4eTFYy
bVGqdbvcRt/B5WdxfD8LDH0CHiquF43dUWOVWTqOIH6H3qUIQGp8wcnck2ZA
ygg3JpO/8S76TwCp7A4wcF9s5zBRSopQPzSJs1yLK2WTNZzw+2UYLkFd4VcP
FH99Ncb4j4X9UL2Ug/DoC3kUqTOzcLIjqWd06jceP+voEe4YhRJIoNU5ukuq
akQxuI3FWl+E0GkVc9vW8iBmi3rPCTMJMXLMO9ZJ+V+09/GAFrAXhSW3pyhq
r9p9awrb+EQ9vr9HyCnMEPelZkhk7AQecAhy+dptCEPAoFKEzmj35nX5WOFF
a+oqz7Luz/7+7VGoCEkSFICvmaTe58ywmC4rVYYmzavtMbS6jIAjHz0hZsVX
rVNS+xcJCVeClP9oQvNY7J98lWvbTeWu3SkcYRuAd/dchwvyi9SCP98Z1GSj
L1EHaDyr1PDatokPfL9u7a7KCRoLykfV6a6pnCrWwDSWcAj+gAqQ7x51luHB
Ag8aTZKs8QKjqgrJ5ujyFg4nzkyieyU67O6kgaN7XbQ9gkSzW0omxikPtNhG
4ZLqEdHmpt1pC/pvlYXw398f3LonRP+9MHXU/viP9bIP70tus0yGmtqODWoM
x84dm2OaYzyUeCiupREmjr1ZAsqgkVzdBIBRoPbZizztPHNNhI4xifdkyWja
T5UvRAQfP6+D96EXGAvck2l89uULHlHkBaTm8pApI0N8oG/tPtCFIDjZ3ZEf
dxOgoNjL5FRLDOosrteR6lL5YaKoyi7UjDCPldRoWbv8NFMZWKNkzqQXiymE
VCv4mckQDSdyudtsuA2IjcWrSpv/GnzF/RNi8iuFoWmTiCiXod/e46SWfgTI
Lm/c45gFZS/eonr7/5AHN5xilEZ8Uc/KnHzGaRxNJIgox8YakRlvE+zAmShD
RVhR/ElL6LdqcD371HknLW8zDssnHl6QzIlyi3ITXr3V8uzlwDROcHbZ7olq
KQGq4RztnWKDm6QL2PCzWEeqIlUEwVO/UUyxAooFE/sLhATtzZpeJGJQ5zls
lJfhS28PRWKk/vSp7d82Y/ew9x8ZJIJOlLsADGwJgsmCotKH9cCvWMWRrxXR
8oieUUZHKN4/40ey3kIcdQJZc3nXtHDqtx4pFuQKa6FRmzEzlNJ7bIjaYTvt
n/+mXMu2ACi5OK5VNMITVgLbFLGY2frTJvmcPNZfXt0wby6KhA+31HlXeSFe
URI/ra5So4QMlgMd3fXmU8yjV7n234gYy09yWzih+/+uJ8H67f8NGR1lXUMy
Vs4YAPr5OFZB2n1eFgj+9PMgmOFEA7VjJMf0FTtjUrcpUqiaWP37iC3N8U3R
OPUeJNPyRH1QgLnOGp62lpZp0/w9il7Pc2iXFHLn13jGaiEOPUcEIhzXQlXO
H79280wgK+/TUbmqnUjAE36nVoAuq3yh5pxdzGUuMHpNjnUyTU731E2IuslM
MsK/+5evWFPgjToQWz8B3Ks32ywagziqbYyRL0J//QuyZuvovgT5IMNvfkwG
lHRpzbN5v+vzXtOTKrO0ks42Nhfle9USlbQ7Lsw1/+v3LhQUo+wegN20vQcB
k1lcM99fZ9wAkjiiHkmN9ciCMhLHD/twp5WgoTcnEPFszIAhDcm7U4+m5Umw
PvFqM2t4gLcssjRtjyO1J2lBcceS34g0pL7qyNfds7Q8cUWFKtRisZN4evU8
BYBDs4RAnhbVYKeHKbpYkrA9meqURmk/2IDwILr308JfsCzCzEvi+DObq+D8
GFe8bDwdWmSJwn6rdKyuokMutIalExCGV0SO+NCgLXeUZhZM/Jxe2x52mlUh
xHgAp2THH2ooxK5FKumBV6z7k5cs66jUIURYOcIccZ8snpHcdo2rsEiC9lcD
uYNJn5adm4NlHK/gtoiMKkYAMF9FiT4OtbCjO3OjUYjj3C2I8OBWH6nK19jL
4WEW7KzR05oHX/fqxtZek6FrdT2vZ/Eden9BSfd/dvQ98R7D5KXxeFffbFNr
pBxKVVLEZHJ0tI9XMcPsF9o5jggyGujXX9O2a3YBQzgBWcInMAbFtUG1j7R4
rK0JOV26BZGSwDaltD+8aHeZnGBt06Xhi7R3yQhqBkBn8NgRmfW+uSSuraGB
it/JFBGt5TtQaWIh1DI7N+19uw4dCja2hqi1GEYvIHYi12uaa0Ofhx+4Svt+
m1KnV7txhNgOu0NJ0m3vENFc0b6QCxaM+yHPythhy7RQKxFV//8QDIw36Y+J
hBWSXXufqZFh2V8g9ojpIeo8z6bEe+BxIe/VJk9e/Y6YA9pNU5h8yAjVVmoo
kbRhcKJ5o07z9sHXLPj+p5YyVgEgxZX/LuojkF9+wh7WMZrfSEZT7HW25zEr
kxS5pf32os0VqjpEJOq5HOuafcDoxloH1JzoKDBvfoiPXFynDdYIP661194j
ZXTajzObsQF6aaOZLPUXVzZFUbcpHS8vWmPBMmdbOgFVZoeluuCQpOIRsjVI
ZVIBtLdtkURO5t7kfLM/qQWL8Vo/w2W9UW0m+ujm/u49l8zziK3BW7VI2GGf
V+nxmrWo3kpD228OBvwYgg/xLsSlfKfGQ649fBBf9iBa71WLWI6RKSpRUsdE
DlUvczHF1gsiJa53UOZBJxxFBV7RCS5keOyacrotG0jD8qGlrG6J111nsnBF
mu19l/+/RDM9Ee0/xrWG/JBORTjKjVLfkRJ8/wdBshWmbNLQzUvi0mScd5GH
4aBaBCJJ2ysQUHKcz4LePDNiEYUyhtO/ktXuRmsJmJ+FvS+E5PAbx3uiRWY2
QH+su2zzVXJHutZub25xrjjP+O54Da/Qe4BVlHhDxUGm3x6rBCeH6kdzL3Yl
FTkDOV0oMnrq2Bo4Erwp//VJH4QdotkcHVi39GRPZQQpeYnGO3R3Rrd8cKPM
df+d1m5uxFBjii8EOQhezFayIiVDPrvGCmhgnNzjLDW2LtzAOaoYW/o4mk+G
W23O6TKhyEvZOsrM31w3/tm5vnxUyFks5DQXV/H3Nl0n4VougFiZcoWfD3cS
oN6rvtCTSGHdVfMunxfc1mG6T1JFvjIhKc1LJF2icys4fIQ8GA5WFZwFCcDt
0DkUWWf03PSpz+NPSB+P3UHloUNSrihfLqse4QHjLikK2xIvdxi5zEs3HqWs
jImLVzO6ZaQa3EN1i2Daql4QwTJpgakNZ9a1tnDqEbmPiIvo75vB3q3aXbVl
55guI9jZ1sBQ2WpA3iNXc7HkuaIxFZOtnpGB0mv9S7x5EJ0TQx7eziDXljym
/r9SNulZKKhVwwPYpZstWimPwaSDm2NGVldDgph/j6QA/qyDg6Gd85O35gwF
T7egvdWiRpZ4ZoDtz43aGQBVE6WHLHSK7JkGCblTk7jyjy05L3DYgho0XOye
KkXgw61mxRZ99wHtC7pGD0kkDykHSdjw1krkb8POZ2Nq+1c+YSyAAD6GF9yC
GlnWB5rpyXtTNh7V0Fbs1KSIEOOhaqbONSzX2cUlLjpNlRMkf9Mmnf61z2SX
GaFo6ZshHUmj4xaQJuDik27aNgyTxyOskt+hHdjwzHtU7MQj7c4xFtPbs429
pksjk5vAvVDyfjAhYy5p1lVx3I+Jp87pD/KVE5B0iKD806omoA7j/FQ1WFWi
d1Nw7p6WozbHRfNhl2K8PK6R6BVT8u3+V6/azZ0FaGBRpaix1Izs83RIS8Yi
cBKxD+y+feLdr5QZ9qPFk2CJFUXwJCyqeropZRsHz6vtUet9q9n0XA6U+bAX
mbQZ/BKTVkEurpyo54JU8yJMFyyfmv5BrCNO5WlnZz/DEZplcoYE+XCZ1mym
P+7Bc8Mg12UaoGws+OJ7VROw0prFtxPcxwTZAynhh16WPThgWzL186AcfuYC
R/d4KFtyvFyqLpFDS9Mr4VHtPf0SwDkVWS3TIM4lkEWu4TwJdodAXME3HE/s
dzD4UE6tuWlV3GjeIiLZxKJtq313zWd4JsGBFVJkGH3mrr42EQuZZ740YCEU
abuS9hyT2heg3JyiUs/ai/RFC4WeHj3AQSh1dB9y8wdOrcD41yQzuW53p2UH
j1ieuVmtp2UwmZoh1tm3Abgr5O820k0CvDHB8Pj9pVoVeHb4Y+weBdIUZ8wH
XRRtpDYZP0VpxNXn3CqqZuh9dmH6118VnoYXU9kRiiXYiqR1wfS+rOEm5aOP
zPQ0QnYvfAQdKx6wdbkUoiNf/2MYaWJ7MramOW8wwgGkrkJey7UNQakUYrnF
wGb9lWqYtsbhGNSh25kGyty8SOg7k4M163OB9+EzY+AfKAwHb/dLTJfCTcoy
ko78NobkWTnCbJE5qOXQp7JRfcIyuz6y3xBxyNmAr1U2stMMYgtQFqQJ98rf
OLqN2Z9lZYnVoa51cFuJ8WV3YHyelHbk2ub9uBK2geSgv4top/TgtLAsH896
WfXjIipdN5qOQDssLC8vJ7fi8Pzo+6dRDQrYxy8t7bWDiLcTZ2nuLmaNeOaw
ppmON1cuFo6NCvDmK7skn2TlLSZWAGW18VLR8Ui8u5wLD68c747+haXxvsZO
lFIj206nbI68E2/pSXN6grqglu/pvR+ZQWtD6NB23mJZcrSMLkb48bcJ1HaJ
mIY18qwDXSCf6dsXhP9FTbVtyyjh1RL/Z/h4SPCwpqhlGkF9xKQWHabMcGzx
tCYBxpyqSWYo/gRAQPKF1O2uZx81QmWYdVGp0eIuXAH6b+PF17qD4ceUThpn
WGxbtOICu//uNqw1Cqwo/axfLkhnMmUXsMiZwjKC+DliIVPc/x4IMrVHjt/J
tzy/WHJoTHMSrzZw725vkPtY+MuD5L3SKd/Ovp9vsCiSoJ19rC6HYqO85MdX
hAU2NPDj8FL+m47CppDFExkjhv/1fuq82gyfbijQJiVviugrMxHgpQNCWGft
LhkvCs5I/mUQCYi9bdryLKIAfDP1JqPSZMpVev6o5aY7yhDLaz4Mak+ZpyqY
iyuxNtoREFrFy4wvcWwPdcfymGGw2xvuBX8QOZtC4EpYj17p9/cCumSDOjrV
Khl7TNWpxEo6jjP/w7PREFaKxtLkOgkh7jCujuTXoB9YKYKSkrpOH3DGhWt+
37t2KR0tizX5KCiSTU+VtBSjTtqOI2/ESxnQzGP21sGHWcqWCS609xOF8Yhn
/luZSmwgOmRw6cpmQmLIiDG96bgnbehjqUO1kJgxUq0rJZL81ZD/zEo0qDzu
6c1u6PwT+zZNtThmuWzLGZ5fHoBuVUnKYlc1bdgHPcnWVDMmnJH0xvF4OoHv
IGXBifUd2phGs2OCPtMU1f0t3Q5ZhOSTG+EQSoCleiSYIjn23J3KqK609bCH
mlVPbTUHn7E5o5gB9HjZH83DN3iG0CAlepX8Ug2V6w6K4Yv+Adak5lmtqVLG
giQoRoKkFVUIGTqYS9jTOdzEshINmnocmAM4kHnuxvfx2fRgiwiZGzkmp/Hj
c19p9gabv7IYy8a03vwvN5uyyiwyZiVFrTnBAPo/Y+LiB73SrgansMqEexea
ZE5orpNws1aNO0tBHeKSr0Osf4LYkVKh3UlIq5uEULhmXadcZHsoysco7oFM
tP4nDayhGrQvWAUXM5KQGhjEHvE6gfjrrFhYeee3xFTgJaWhCnH4tNvl3p3D
UXTOQO5Q4DN24aCdpuz3uex5UkFNUlAK95D3EDyqNPVoHwuvPL76fKHDjDjF
AIjhCrophyFei99Qsmx0/fyvJkxe7GIZRVQ0fJGCQP1JxbNg4Q/Kx0Me2d8F
F0srKiRC7dcTS76oC8PaSOR5sc0oSkHuee2Uj08JXSX05PNwYK+X6Ph/9x/H
pfyjKMV7A9OenvxjG2/5SqLTFpcTWc9cHAagguZEaOmUuOqGf+crnOBSKdVR
UhxdBweaJiUPiL+SN5cUxxvX7qTP2Zgwtzym696a1giCU8oqMUrRMm+gV2zH
LmMTOv6KVztWETWpoEvM+Rq/4AihxR1MzUSsoqbdtmohUR1v/RiwLNVfC6hZ
lZlHNusLi4Z4qnwFYIzzcfswm5FmKL31LeS9ErP5S3wGMkx//rKZCrkSPgFM
uZYZpLCoYgoCW9uauXd7q+ZwZa8axjuWEcaGvaDDLdYU8LPd+Mm9n2TF8dDJ
1TtUBP94NNoPHMJQluki6WHfzNxzo0II7jZ2AE0flc3aYOnJGrmURk/jFHiv
6RpCJCzBASTr9in1TGVJMbJNu7jRZ+fkE5Lxq6tqc7T1YPB9I+M0VF40/s9m
5Uek6tirJyn6/O6ClzzwRuHid7XQvpYv1KGqSSr7hQnLPUpQsjKtEVYbRQAM
FQp21gIhy8zPVTyqgM8CRiMi8nn38HDU8OiYype8BihKyz/SQm6tzzFq70O/
UFIQlzFd3JIBcygv3nVu6DwR2cnei0mL14jLTXNcW8M2a4MSfKUh61aXJP8b
318aaDzx6ZVoWmP5QyeKwiTwfzhBbHRMfE+3lLJWZR3DA1bdp5MZCCmEbhec
wbFEePIygZKhT/GcNsKLOUXjqjIzkSRJqlmrGkrJo0mqz+IW9E5Y/ucHx+p9
iTyUONov8Of6pGwKdPbkENJ1FlrjEgBsojLC5Zlx0QYUPaEasgYvJzczRldY
tDIJy9fLlXBof+KMdNnXXYqOeGTmIV3+0nPQnoZAGSgJJl4MTT+ZTz3Rdd86
jNh99R/Cs1yk2FhAstAqTMRRo+ZEk6udyd3wMeBM5IO5k8g4d2WjVTOTnSbF
o24tltchibbH7kezNUZjtcxUc8YpnzDgUNI7GXFlzLLCvjrc9Uz/j3yMtQ3L
N752wvVoXrDjQq4X3a3zIngffYs+5OCsGTR8x+QO9I+2ebvd2TX2q13oJkJ9
VSYwUnZKjpH6U2JpEbl1/KtY6wgVhQnQQEI9NoBwMON7ZnoASo7TTlL0Q040
/xAZdUymB1QLDbgnnBEdeL3aN13u/YGf88G93j96sC+I+RIvEYV1TbjJlaF1
BfYZnR5Eqf0BYRw7n2VNZAcI3b+uJAefQUG7nGSvW9wJ9loA3ZCS7KqqRS/O
CSyGrOxE3eOi7d2rKWXBvfeX4SHVJkzgTmI1tGFC9vzOU1TYK5jHvD4L3gWQ
5EZdYY9+R6z1dQxNvSKAwvglO+AnL6qpoR/f5Pw0hRmvbuE9M41cNwtVyCjo
Ai+c0GgvtQ2MJMi9l5IOFrvOiZDluDIxZfzObmf4bG4jU0EpVfz5VKXspw/d
zle4LQufPxa10eoQgAzx+/9BpgitKmSqZiCT9wvVFAuDttKpI8/vDJ2JQBNA
tsx3tiQ5b/3BI3262B7PcNgURnNASxL1r3SMYKN+8mF5gVk2vB5UtuRLxRka
j086cN+bAJMODBCYpSmIgNzXjctUfl8snPohrFO3RdD43u6tY/J3tvY+cUFw
YWSfVqKggB9DdpBmAJ6Jh7mPYMVSagz2pmxJLmDYP0BP0qi14U9jd/oLnN61
38vBDkcORw7gSql1vRh4yBNxFrnRr03R5Kds2PWXwy9XVz6+r6PSHJsRioT1
AQhmZYCASr0Yf6l/JGDKCsxIAOMNoiMfZitmD1fKLQ10t2GFzkOt4cVoWVFD
Z7X9Dc9hTeltfo9zM0VcwEnK+GNha7NgvM0A+0lPRyKGOhevE8wWSjrR67cP
6UgGb4E/xlmrCMY/W9epSvjPC71SHQ+GZDb4LTjvmrLUDqkmVAdy6oRWwD5K
YpcaV/PM1O61H27VsF9n92TYTxZt0GzC7zXAbTAaBJLGgLQxJA+R8b5fEk0l
hz7t7OKMpXrn1ZsQAO8hKhC58x4DvZvG/hGwVh0lgR5dGgVLhtxkLV22WHrA
ncTbq5KP/3JLMz7oO4V1JsXJH1IaYRUp39EJ2q2pScR6ttu7tiOhfg59VQtW
kTZtaw3pxmBEA2S+Us1XPo19aRFc1153uHuROswJqvVM7reH1w8NlO9P6MMj
Xm5whkBDfTzn+HgLqE9uh/ozAsW9TicfqzF2qRnfCyw+t/fEjS/F7FCRhDRo
sfo1neUeSdV09c+a1aAPbgtP15w433RDhjo5ujNqeLXMgs+8oCBZAiHNLQgs
fTXTZwLGngelrX5iAdixPcgjSA6RzXd2rnJOTlVwhL2HliSNvtN14WPKLGNM
UdB5LWXp5g0OwyY2OEldBvWwCUkCkahGmyEeBu2SxfM9MmCOfR5c9TEX/Gmy
YFCxC7XXq5nANOtMvMQqNi7xK0dSvXAAwADhNnj+eN2qoJgRpGHR39MDHwGO
dtIs878W+MDUCL6CW6fZ8hfAru5ECU7yeFRPAiDdu7b55WbicGtMWF3sqQmc
m3oxhkFtcZOmTLuURzA9vljUeDA+ft5FcPm+YAlicwrYLwxO932ZollkcXyP
uM/ABWdEh3FDLLZL//N77KGzdy433djp3BpJtfXAcv7ru8Dk7RwBvzHKrYxv
GOPgbAez+axhDRsFqX7Cta+8BJ4DK8Pd7v/1PmK4HEpnyiH6QYFcETx6oI87
xGpE47Z3x3dGVv5ZKu4RewdXuR4H9N5jbj/stoPmymutkJhM8BO1mzQT1anF
Wt+49CSwSfRNGaCI+F9SgCv5Ye0aAngCQG38FZRXb7bK2mXMXDC8ctV6IrxO
uMpLjXlVqq4OSKgPC5T9xH9WhH94h6aD3OmJr33sMGJsdveCKslqnhkDC4X4
xG7mXxwYa8WvLSYNqyfHfcxrd0IeF5PJn1DWc9z6m+IyfRahO3AgpRGuyy0e
s5AA0VzXPTIbPoihfPuy1aNvRskrSaqLDNghma/loYkT/8VwFPEUWrAh1Et3
9ZqPaKtdrycIm+cmVVsX48FsH1BbsnfVSsYR1Dds94VmtOUimg6hJRxvUIrO
Ynq9nOb0LMdM4m2ZPGGd4AvzEMYTqeZQrM9FwBC51k+zoW3uE/zdrLymY89v
YCgjIoq+7JTw0B+GnbXhJJG19pkcuXS3TeevebqY7wwvqlcTMdYBKFGaRa8a
lX7YDVBQ/S8xYFYGNV2dp8lYaXi2dAJZCEcvEV3AmmCM7+t3GjZg1u2589qr
kw/Q0pAl3iFmpmT8e779elY4Ns1omTjN4hp62aZCLehO21ii0tnR7miiwZiV
C+Sq1o/kMQSvuKz6S9fCwbptW8tAVYKSM1Oh9Tk760iHc//v0JhwgfA2vrv3
d1nSMIjLFQdremfyZYtnI9wjuuj0Pz3/+J+EGeTlNhtNvYXe8HMNArLz+zE/
I5ZJXFmFf8CXeoVDVN6z9eMRj3kxAfpA7PtIUlFKl6sINFOvECnpubvbSvDf
ht5itC8ZlQCPUoh5IzMuJAlC0IjDEUcVw93c8jkhyukSJ7i5chlL5Qw2RDJv
uUnNc0zD3Bfy7q12Yit6ae7OR4cluEI6c8HLzGhExYYrIdy/6xx0gAXv4jwc
O+UNLj/WQvAOOxBO8SigrdNh0BnoqIJ6NhieG3qCzsvc6SaSvxlLKO3jJVqY
RlJBNU8Smi5Ne2Ni9OYGb6ePh7SRhBbXk+vTYuFInwFCl8G5MeOkG41H8aA/
dJ2knluRMHuL653kwP+ZKb1zO5scqp/iMk1A2jT7qDxqEo9Y9wqvMFMN+aXc
2/5yKqHXaqAklrsHESCTAwdxmnw+43TJ2uZFpCIPCmKjWfObYDu0nVBp4++8
ogpF+24ovBXWjQWfp9tEkY+DkPYyv2atXoUIPNPUecBvi5pCo5sTk1vRqKej
/BfDi1m0oGTpo1scdmwGRQhUdTQzMoyoLBqPpQTm6ATKbKAn48ClYl0kRfdz
Wyd96YyjJkkWDbwrqh8bjBKxEfFMuEUINW0VF1i0XHF+qdYyKj/8slABjRdy
hk7qdUqEr7O0E8HrRtjjLyR+fOykkjzW7sf921uMvVlJIJ04kGi3KGzYArmO
u1Ch+Tha0zr1RFjHA8XOklDkOpdy3wVgnkhGgAFgUHg0kHh8eZ1h5HBBLe6c
K0DRPEaI1eazpliA039ah9qfENupQ1gHlkWGTc9maIIMiREkMZPIh5sCfIbA
fAY73DNLWD6hM8NBPHXKTkfo55Bf7zuVYQ7obBZR6yzAjX3Mt198m4eof3QH
q4DIdTMVPFgyD/EuuSueMbYoKe3zinZZEogcRVwnz/cynJ4Pg9RSjb/T4S4B
m676W9GJ2ufZszfEp6DZM2v+h1o9xhvWUbFA9WTF1aAWhM/QxBhqAZt8LvGJ
6ctg6xWNJlnLJqgsfKIS4MmQEKgkFHcOMqapj0OUrF9JWzUJCqmjiSAyHz9n
vHWIiefhRw5P3wkQ9b8ls7jPd4ch2y/QWfGX4fn90HrNVCQK3t4QPVwdp0Nr
TrB/S1AOQQC3kH4mAIbUlLXo617sEErKi2AwMR4MdZyjnAXs0zVosWhSZPOU
9ub0RFMUUnn0g9VrLIKEie9q5FvQ4epV5lcdkp5d22UnVZ4zalbhfmdPvFFE
ciyvogixvhtgfXDjzo1VD3hOvFieHmrfanZKXKVaN9dw5+NRha3wOGuhEybI
Pe9s9oOfE4omAzk7jDRrUZQRWDkAA3Lm4tXRIDzgAeI/0161qZ7oVUD4oI5t
/nnwxdJlemEs/zZGRLnH2DTwm5g9AEJzOvUnLWf0hW2XtLvzuLlDuWm2UPJO
2VbqG0x4voiVJTkGSDUw2BzHr7k7oO8196zRWLfpPLAuBOz5htK14YWD+Xm2
kqYXgLKBXGu6E/UC84xrlcc7Zzd3qFXqOGOY9+8eFtIGMDriBLU74baIpTPK
5TsgR2/jSzPHlcKdoH/GelEb1xGOCGA4/nMbMRqLcYD7qBXkO9mtBtrlfvZ/
TK8KZCkCLt8jRBwDV8/W8SQtrW8pnAMwsGRI6314nbBZV4kov/bxAIB9Fedg
+8tYRyQstpcE/4/db4plZU4TJuPbOHXbS0CtsHmo1ohkQoIA72fnakinkAZb
thJlH8xdMefK9/obQ+xsME6+hWJDgg2tPSrAsty6LSCA5btSdNOlW5zJUxuA
I5+1mxspvjbOlYCKUFwl1FAzo3kfa8OgaVv84OdwevqT0Vf4G2p6Q+u4No7J
lllHWj+H6kZ13S2xg0wkEZX0jcLBUpjjyyPZPqLzPY/P9BBD9Fbmo9asOoiI
9T2ED47tzI0EUL40TMG8GhLhiL85lYYDvE5dcYWEc09Foa5aw2dGH3vLwMeP
vPRn3kP6PFERDdWWJq7feYZuhemxzc0vavnaLLjo2yy/ixYVdBoxJAtDTEA4
1VWpm1stbViYjMVI8qcxpp70XKh+9+cVZaxquXixeKWUNgiTMiGpx5YFyHYA
k1Zwo4jF+3NORR8VitAI98TKJZTEPe5lkAdYwpdASKf9KWOr0aLBpvfwbvtv
dEDaXSPO/iIev0f+SJUgaP0TQNGcLI8wCo3owNqHbJZPH4NhXvVr3OwXTPkf
cUSmLvMOsRfYBnFyJJgIlD6hd0nNNFmc5b8m2unQWgQfG2hq3PGoq0LSM7zJ
uf2n8sh09jXn6HtOjXs6MVTrqGzyS0WpEwZMQMHdoPtwqKZIccQL1CnjfVTN
jQRiF50MDEyj2Yvulo9NGMJxYBbb2QzaTSevrY07j+hv6kHwkHVX2o9bG1WQ

`pragma protect end_protected
