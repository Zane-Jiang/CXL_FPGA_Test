`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
CU4nVsGDzq9stlRciZFTp4ARZC/RSddSZyHZE0oYiRYQFrEoR1jRyl2+7SP8etVi
4S8HmKn0PAZjNRLm01OviqoRW4Fhpgi7T7bZEU8NA3MvWoz15E3zoDypuKBbJCEA
NPBoHJUifVMfSdcJ2FKYoaAGearrDpmtCLKad3SMRA0=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 20080), data_block
4fKVwxsvh1+I528qecVu9u3rNupVjWV69Kx1kI820QnIdwRF8Na3aZCZdMluD1ot
rjKLaSGlMjN7BJ5Ue/UNwx3Qsynz8fYq9No4TPp/CA80T4ccZRjRHnwrXty8zDIe
w+ReE58oxk6BnMqg9LZTtB9U962mPjF0ird6eXCevhbFn2knlLT6bU4/nqHGD2DZ
kYWMo7EyK/kUKgCQkrakzwNQqtm1dnOoBv/Aee0qjLF84R8zFzE3kfUnw0Xk5yRS
srAy28Eg/CJaTlv8NflLO7jD6kj755BfWkaMPmzP6r995/msY1Jc1SrHCSD5EzrK
vPxfQR05LqzWtSXYMMI4XVqcPzlzTM1FzgsZSM2DJ/l1DdOXTe701ysQV4h865bX
YG4dppTIX1OI7XQw4WQg2Ev08QdMa5xgUcs7PGMfUb2rl6Dhu7CguP+wkWq9fk96
TWu7zeGyCIH0CJLl7vM9RbTJP1ef8YJu7a64Gt3w5j/G8oFBgRaqozLC6LV6+LmF
WEeATxPBA7SAWopWlddYcb6VaxXGQxyJJW5anKCCf6f24V3DtSRC0OdKF6O12r8C
lb3ztGZcNxuNs9P9JCcDDTbWSlU1tj5giZmnJB2apRxtCF+7V//xvgZwOH8wTgRz
u7xP4vS0jGfaAobO3VHJnlWp7tG1HbdFwoQ3rI5EjMbLNZ3wBAM5Dj3bQOOa1pnb
ek48qGCEz8ZTfi4uufzGfZ8YjbhuCa9+n2rglL1BvpB/sgxdXIrBWxSF+NeEToHP
bUN1YIml1ji6q2QC/TChCML/WuLen0IfKdF/mJsOwpMC/6l9HfJoZn3MOjOItBWv
YqH+UC/TRt7b9atW0Vt/FfN7IUknmjhFZMkaLr843bd/e+PYo45xZGYNaAK8MK5e
kbyTVvMcFVLEuMSmKQB/imOMMnl1EiZ4CIy15HMDM4P0unzQaWZxxu56wzd1KVYE
sHrx2rSwbT2M/SMf+QT8/4ZGM93JkNhLqmuJOaEZxt6HZFYhSC6APuP2qtUb2DOr
XBUwyvK41BlKPhZ+GWkhZjU5l4Q71f/y5OHVdnsq0CHB6pNGkZf1Qb2OiFzm5zbN
O2M9ncpjHbBwhxTylZx/LnjOsaezieSiaPDPnJej1KCObwtQ85uiAPikia+R+9Oc
5bfl/dYJPItAJ9e2eXiuSUK3zQ8rbcVjVZAic1ln2l0UZSxIZyFih8J4xv2Myxm2
sfy9qjks5KzdzM36egwz2BObduK2eS5wh682D7jFgOxPK9epIintrVjuhGVdBn36
Rgs9BrDcCt80fjY8WmS5QtxAALp0C5q+xkzIWdKQiEKFfSBIreGoW3ZTpgEOEASr
UIOsObkbo4JBQ+jkf6PHgxUbaR7/s7SrWbNYUW1uUj7yCN8ri6sn2hk6CQWyAyQa
ux62ZajA41CjGbM85frcYOtP25GMUwX+8OkJXcynDgcw89duLfk/eNFgiEO7bbPW
9qVG4n3VMv1ShbiIGpE4QlhnySTwNE39WwZxuyn9ECnmq/5iZJbmbnlVbQRTQ9Py
789xyldN0oK1BJHSsBqbRuDH3E72L9tBdBeS9POK4fsCgjVMPDxwK22XC1BPJoZQ
//bIwNFHUWIiGE/wa77ljJxXIzo27JIzW9Q3yW3e0XDklJ7YAyMlvPJr2yWWR17c
ToIkPp+eC+CIWzIvSSoB6iG/+OJKg+bcuLQU2F/rQcC97l1AO/PM0WyzoaGbnMnj
2QtZ6qaRvrjQQHHHomYwvP6snzikNS3yygmUZMdv90t20hYLA/IRExQ51qeEZZZA
JJkymIjFnMlkDRiF4unHKYOam8Bh/XrbT14v+35ayiUgufncDk4B7C4FcpT8sQ6P
eDAxtnLA9/y9qbhs8iiHJioGDcbU+P/cpT6Nt6b1T9xlQVg69qZ0cG9oflzz+0P0
ZzDJ6Hg9aN8aTXbkq9xBlaukbPvJyBo7qy/3gkeI5MFi4D8IVBlVfgW+jEtUJG14
+8VGK4Ikq6DV//dJmdqQJIBQrADysD/wknkfRM8KI3gToxnUTh74zwqESFZKrGmu
5CdPJ2Wl01g/4jKnpTqeiwLfbPqkd8bKicaozoxicTu/UJ5guW0MD+0mLfySI96j
yKoeu3xXmXdDwDddRTvIZs2cmp86VJhCGIYj9kA8lsh1elVyj7M5C+gbi1R3FJ81
IlSWHxDDzqtS3ESb4J0YK8ObdJQQdo8WVgicmfqhQn4HA18wB8OmAcnOx4kr7f4C
Lgt4WdTO3vyawf8DAxjYPinCZOlxxsvMz0dyOk0di3eELLHJEoEyrmz9nW73F53B
278Eb4EK2EMrCCEBBjz9GVqJIX8+J4O5DifI4Lfeybd4ddGotqBNwNP6vEU3CmKx
RDxr6NdUfpz5/6Rvx1PSk125KayzTWDkjVoUW13AHmyVOJVpi65QiNKJgUbTiBNi
TBYlSja4a7QURPMhwETonNQKVfo1i8BTT4np3/Ls1Wwmlr4D5cTFAr/q4t3TdMkV
1Id1J2XFHsbYnGeYuFdSBIdMSGMZJvnetPnTkIrKGWLDhc6MU++6Rpi2SCbYO9yf
SgV/A1Eu8MLYU0ulAFHd2ahc9ffME0FQonDOlZIYsL2JrZZLpWRAC1A52Fw1YwaP
+Ga0vUOEXmm86iMn+PbKJIyf2azH2uOhFJe/JOgEQT6ValXx0zWtGRWw1TNMoNDf
AgqEs02lYDtDCE3gSNEl2oautfjpjPkrgsFVs+eIQKonMjxur5ej++6nnNq/OLR0
x4qI7VeQx+kIIJe8WnDyI34LMfWJp4T8EpuGSXG3jQzzGY1eG8oFtfgrMpsSDEsR
bSNyGuyym39JKwLixR5CjblcEArZORT8mFAlfQuFP0r6Y48E8hkBNzdMJR+Kirn2
ULSu1gxRVAzSYiX5Kb60LvjEr76xz/DHONg7gdun75TuPvzWqhsCrjdT3kVKgn77
IgeiNLxMq02F6FyZWkXn8W+J6KfTCsJj5zmmQd5n8/oXEoiDroLzF8Y7tiRfhN1W
64psUXJacEwn4bCcWq/giAO5ISMSL2gwl04HH76N6DJlpiqJiuNs052pzkQWbeLy
+ZX3hplHAg3PDmrw3c9XrF+G+gOGb/fiCFzkHxPYDK1x+BA/nQKN7nyiqlK6+c6W
k6ijv4dQd1vGTf4Q4HJo/l3fNBwwo3aWCsmmU/gJuebq7XjnsyGvMgLOqF1aTG3e
ppB8S2X9xHEricT8KXgfsQmeZ2pbK+TF2M1mM1TTKsU9WzJ4i77GlQrEbNVlA9xO
wm/0h72Tc+WU86UfxhaOEr+KhOyZb8EGqhwJsZ0uq6o5+6SiZhtPbKJy8zfzb4O7
r3DsyeX79VeaX4fci34A6OM5W/Yxnk/MRjcOOOYmZD21p2Zn6vUvbeGKqPuYmT5V
ihAhtZ6LufQPjhKvF4GcOZyuclSkQBkUTs2re0DigiMM5+HyShYOln5zMjTPBTXY
NiRI/e6UNr/H++/qcOdy3sFXyAAqZAyzzhCoRSaFvJF5ravlECSxDWx7HqnFx9li
4J4lEK5+Yg/y+tyCS2ByN9WqxInIhlPyS6T0ge3nO/pjNXUBZRD7BZ3DPnPHPBEE
fXnRnuXJ4WUVTSllcCtRMdzypDJ0pDzjZzzkDRnZ8shIJsRp0WN0b4eVPBya5scB
4Rd6XW+8qnMxcVK9oNYl7yewkKfJYEPOVoljNtTrx19x2f1dbUYVEw5cFihMFvmi
SWoiXbtNPV8sobumymx/ICCUh9FutRPLUFL+jYWP3U1PanrEqRqbqrOEve1cYYH+
H2GpfP3n2FQWalSJxggvJ300rfL7l63HU5wiMEAX6Mwf5PX01Lk7MRt76kt5HnNu
nANfTnK30DoDuMEkj+EquKFWRKK6kaL8G4E0Ak2y1MAMdQa1mMd8/HNo5cUeDIJo
0oEoZtsjTBBpm0kzvnYGsdKZsmgRjI/7TA3JGCX3cj2qQX6L9XFkuzIrZPrPFgpe
pb7txERFW1V0lclRlmbCrwczt7krG5bZeQXiAx7AZlihxA1A0ZI1IHP+qkP2YxZH
nb11SZdGOPF2UaJe/eW39vpE7m8+fuqPtICxuZOrE/p8p+AzBuRHR9P6m42q2zim
BqCUv6sxSQBd5Em1//nk7m16DCkRi21whDuaXLcUjZ0l1pGliLh7c5Se0ri3qGPd
G2LgC32CgSdhlhCinsxoLra8cFteisFlH0kiqW+DA20KZxldMopit2zb8t9S1y9D
Gtj/Cytn0f4YyEiMHkKV6Qj1O5kTSE8oF1C0G0V4gv0euYZDiWGAeGjMVBNGus3t
hbI309JXbaBVTzWMuKBqeJ1BsqWwgFlJqm0uDRm4BoWdSi2vl3spFaR71kWZIDnr
qUragrRdhJWFuDvpFUTAtLcyGg7h7CjxRoSn5OWoUiBKGIUhLHYaxMhIx43bcdtm
xn5BZ3gaXc0tIJv+S/DwQF6pxxtGeHfXOxwZBsXIoZEjsS0SG7CojVgga4bRrq+V
RBZMVQZsNIS82hlUOtWuhauYz7ZEnSjN6dC6G+els/KGTaiqYeMEt21xaO4jtoRl
M9t3jUAaqZabqW89cQHpKpAYDbG8pEn7tW1dVG6lIdjEOcRqVp6ahh20lxzkl21j
f+AUscNU3ZGXfhTbdmnu3N6Y9i4//o+AqTm7/okN8GZ0VNHFhmZXeJ0jazBRPdi3
3jN25zeRZen2lQ8Sx2fHowZFu2K+kfOGBxOp2O4Kl4F6Zhvy4oOj2VFfPjhsYW37
dftc6vEgUCrPfKtQLqVRmZyiN6yoQZ5n75Gh2baozulxtpGGV3tJEeVpfm89qpIz
t3bbhi6htjTiX4l5/Nyq66x8txmnTtSXfMGpu0FPVIj4vxzOZbV224AkVpJ9RUPa
/Fh+3h8+3jvHj1U25Bso9S0S7Ohee6IRczBxmdWNJBsX6+fV1Pgyua8Cmf4vz/rr
Ux664ASloXTkOvs2LmVyP1z6PExQcLFrYJ2Rt0F//vsEX6BV+NceQOdrKJiRmVbQ
RtIuZHHbMjdhp58VYAC2gnC9KMSKTRpIZk5rux3zHiE/HS5OfNDmpJ1ezqlEerb8
Y/ZNiXuefA5ZNb8wJutk/a5Z0d0JxBGoV1Gi4nBvJ/tOAo+Ljd38AORAw5YYbn9k
UQ2xF+enOp5jf+B3ipTAzWTXt8YYEzJWUSUdFDW1GosIUhQG0khvUzMCQw0Mz67F
e4A0x81y0uM9tCyS44LCEoddjO++xDKJnfxzeNX/q/iUwK3upytDp2weDwFOZlo3
n025kIqejhPtHtfGHbkpSnWe1me4sYa2wWL3QhVx5NeoyaZrdaU3QoNEgMU9gWTs
SimfFZtzMx3huQjPGED/zlW2g1zNat+KV7lSi5f4uIRFMuXwBu5HwpITxvy2YfDf
+tfYY52sUf3q2vODZpZhT7yCoIRRkARY4v40ZG8vwZIGFCZ9p0wvZv7tuFnd6aob
ieX+zn5xqqsfqQdnFpdWtHi4Pr5BjdRcmVewmgaIpNq8PmHCSqx5iOE1NaiGmkS8
TSd4+NBYiXsZBx8/aqW20DoCpQEuTmD9Mffp6Z8guKUVUujhOiTeAR8hWtMXRkA3
wmtw5NrHZfZqOoU7c1HXGBQDkt615D6MR5SRIAt38Cev8n8P1gmYxCABcFim64NN
3r6DQ/jM6ZpUhmOEF967Ix5QYukJCjco7x9HrUBNwyuHCXTv09uHvIdvZguQr++h
s4d1S4w+zhPQNQuYRuAd9ggfIS3Dz1m/SCAEW5wWvxE0fkTbiri18B/zt43znGhA
piVdkduPofS5G+IwzgXQAjgTBhebDCC/MOVvnN9OFPYqFQ2s71W3k2tL/LZlAZ2l
W8iiIPcbUtY3RUkL6txXROkcnvME/B3ReX98p+mK/7Ipn6pqdC8zMy2T4nmZ4sXT
gRwh+8NRvCiEZG+6X4sHYFh/sxTKjg6oreFKic4w3v0yR+LBltgR+9sIIn2MxCtD
xTzkbIdlDn3FiOBx1AUORja/tZRCN8FBfVDkKjHIVWnJaeSeqSMNNst2d+r9uKJ0
eCCTFH4s3oOD6PRvAwrNi1vUC0iHUH9qDXp+/xRgVHpnQtJBfWvssgzPBvnsEVeD
jR2Ml8FqINThe4Rs+G/k5jo14ZVuAfPBDrdrCgkuK6aQ7oBBAbwlpzYM7vQYJJdn
rCGwotMAFhuSmKgIF390SWUkkm5x7VNaB0zlMXmHdXgKAuQoN6+Ni4BYXX20IeFi
RhR1Hs8sqEZsA9CJ4StWnrr2L/AqOWMCr6JITNcE6b3xZ+wt91f/B9rR0FPrHjXE
ONW3yZz4keWB4NQ1xVYYaWHOQfT0qwcKEbasGKPxxu+NJnfv+WNZNitdZsUKhw6o
4Gt8KMhKRT7u0QEcL1N4u/8iVp6BZRiaOy6UabNc8J1GLhSqrbHP2IbVOioYGIIE
AIPnZsxxUKm2a9QFbjutQm9jMfFlU/Rxu9UbkqB0SZ00dORplT+JXsWLMp+ub1Ra
UJZJ1234yQ9TixSG0v2tQeBtQVM367RIdDtk5YMKdXaZZDOPXF3NmoMG7R0ULgWx
LI2RZQfCToZlj2b8HfjghL5UDQ7JPZW4RDZcxYJXT9XsUf2IEd53SbWyI2dIcLr8
tiXG1odQnLkBdSdPyZknIGwYbo4xW5697PAg0hpuHbBWEw8vlRxUJgXWWSg19ujj
g6SEUVovSuaIkoONBZRhb3dqLycekxtvlLAHliH51NZ+1Jz+ENzZP2hJmxjhz+2v
2M1VqYd2T0e8dlV9h9c7t7cLGoQIviLTOEvuqXxCufZr6MCUOXeZN7tT30POsOa2
VR+8DsbK2rKbAOfRJOLxnSUOD29QXm7Zf7n3d3vcmDRvWZwedMu8E1fesP+U8BOn
yF3xHhA/XFn9RFAzLS/PQU3Am/1L6pWPuK2Mh+4lZzbgNe4Lo7UuXYRejK6aXsxG
Xp4IiedTPu3GLuJEKp7hEGkWyLAJZJVtBwt8PX+0jx9dMlKkOgQEm1jF3rCflP2N
kFwQBNcEc8YmevHo+BFkH2n6ShVtMoJtck4hRQ+MY4W6rEfMPbj1aHipqcQTHlOs
61l05DtuY8Q0/VCNDT8VFnkRd5jwGT2rgfjh6HI3KEfIYSKF2a/Llcyf/BJdjxoB
A83UvjP3ph81+CQK67td5cHJUfbTpFLfe/QsduJ3fR4OwotoiC704e3eix+u1R2W
8FpkglfFtb08c8h22pQ/QtXIHfeLRJotC5uwqVdlOKkRN7kTjswk9LsRbgnSCwnS
nvx8I6jYi4lh2pCmZvEaL+ZEwaefMD86Ui+5AiKzvh+x9yVQjNavdziswcI49oDr
sM8/+NS/osmQl6iU3PGSQ0QbqcRb7NB76CrMHL2lA2iOki5mmyEcmBYBejtR0Tr0
jrkbY67+ydD4OGq18dzXm1TqzQ8HMdUmEr8UfiCBzSQ1XjRaLGdKc3qRlTYOHP6a
n6yiT9KAEjUNSVYkrPXUSp+sVvXsOmSoMberFz6z0qai7tBYBZMu7kUsHev6xSin
ikVliR6W8rMt3j+aTq866+gSZ6xa3syGv9g2T4NlKd5xQlq11c5kwniPL1JnfXkv
aL6KtYtXS/ND2UN8rjjqP3A5SQ3tbK3i1af4D5ooIL6YP1WskZhXcWJl3Uw3izF5
OblchIyOGoQU94UE7yfqqrrig6ZVhPdmq0fVThy7nqmvWrO6/2FLono20Kt23Lx1
v3tE8lJ6DnOWynqWTmql4Z5FmOBfMmvyhfttRyLz/5Gk7NrGMtg8+Frxn5+MMCoD
ncIFfITKjNPFRKddOIhBs9+ODL0fx3f9+AOMm+5nWrRfb80Gijy6yQTAtyo/20wJ
DnRGG0j009TYLl40BQPW0fUIlUU3FKZWN8RB0aYeADCxotROyGLmbd0h3t3SDynk
iMQiEmNuPleBwrVRKkhIldlOljc6RQb7N1x3kgLa1/DeTsV87pmLBm/6xZq2vR/v
auO3SsV9oJWselerKPvlyDR1hat1DkOwLPlA5wM/Oeqce6CKnXxlyLWYI/4n3XM4
1ROsSg/pfRWLz5AdAQFObn6sjQUPc5EKQEomz1XZUAIJICCEIaTpiGHF/JliTyN5
eQyQLNCxN1bwE2P+XSNVb0a9NHsptNZHbMApdzs/O812f9KvW1tyfULHQuAUleON
yxt6EpHqk/RoDoiTHGjHEk4gP12aQ0osuoXwWvw/QSj8ixSDYRvajhnS5+D7MdCL
WHs8bLFbTIIT3ZzIVxfciBT7R1fwBzN7sNytcaD9Qozdwz1oquruoDN+8KWv9BP5
90woy4tVvVA37hLl860tJkfoYbUZVsql+J/lun+pqdnbvEq2eUm5tBxX9+UuoAjV
sqsc9hfF7VwD0eJoi1Kc0nKrMerNannQ474w31qFZoj6srm4yrNlRueWrPTiF4Eo
dPKF6rBysydSQJXrG53PcFuGFvFUvOFYfrBN61yf13wQgmIqJcRHtDjfoG63Lur3
8LI4sJ609fqNpL0V5Nt9tUSLwJiFdSGSkdrnYF5D9BaP8S1QPd4R2cXNl+Ut47oi
UduTYYHj4MjnOod9d6a5shVxlfNGYaxKsLSo0NXXDMOl3fTvI/0pYD5tKczYBgdJ
SC2+7n3N3zpaSHpFna5MyW/MkQ5BBoCTfTUsBzkJHCtTCxOwbrhbPgo05dM0Jsd6
eRmIEwH8dFqmlVghwrYU5VLbTwYho91hWe8G66S4PFEvQnwm4C6IowK1WBVKjNzQ
SowshtvzgxxMiSgseFb3agb7EQZoG8DgTJvvlQaO3+hOfOWFv5Sw53b7m0UKoYd7
cxRR0VpR09ZpL2a7F9Z7Tfd/xppJybuybjjcEb0kEv9PrjpvnDVXjrF3nSQKwjBD
TJJMsB2femxzMaI+yjTl5+dWw7QFnR8bPiUXwKPHln27vizrMQui5q48ymodVi0z
FelDtugldXyrfuNEG8yMkgc4SlriVluhGtYWf8z6FdLuO62Xvth7gdMT50P57R2P
L9xD9a/9uSxu1Eu1/dJiUzOlgZaW/U2prbhgbTxgh8CxmYGvbR/hh8L3kB2GTG/o
T8RAlpWHhl2dOdgKesuvtxY9nikfMFtSmKGhPTBz5mFQc6tEhnozqy7PSOcnZ3rF
8QSBdVaQ+fUWdwXnnixgFSfA/J9FXncZHIH8MKkUbn9wTEzYOBo2WThDkCPcOHus
cE6oS+4BbBOH3n2y6t99Lqb1X2hNi4m4cWAAbTvNdnFqJzhBSQM3gwC3QfvxMQr/
4GM4+CtPOG54UEz1zBpEV2YEFyCHBT5lyWon6W2hJtKcQtgthXSf4ARe+0fXUieO
PDrPreF1BVfLhofAVQWaH8iRiG23aKiafsBev8L5Z6nmLjqu1YkfMvQPJa1OUMv/
8IQ2ZEG6miTfXdxLKAFeaqmEhvTGTiiYJ1FZF3EWMiMoONypngKi/MfqdGYPdmr5
EnJh1/S4HLDPyQ9LK5ZHhFbyviUil70jR1gVbzdyZ+VCOwSzR9f7FuoFJv/wBtLB
lSo5r9i8AIfn9O6nCIK8HlKjwN0QE8bfbtgOXhDK3/HjHqscQcv317I3G8t7TcyN
xUV3RB0xaF6p6zeRJ8A7YdJFMzowNI6hMEbx8cbNn++LrfN4Qm0VeM82kVUvW2Jb
dWdpRcornTQwzAM1StYBNbjXCJZa/soPCGP06pUx7ZeqZNP6yHGxkxFijK+U5TDX
6ueD771CV6GicrSFSEROwADGZ9vstLd5YZdbCueS5dQgNzuMhGuKLcnYQqrrrjab
zPJ11eC6FPB2aNhRLpvTY80p+pAFsrifPu52QwevvbMLu257/XSMZJImALSoeTHf
khDCrkwosTV+iQ75JVLF8+J0BSB8MDDL3+OF45JdOuG9h4Ydg857YDyGV7Cxpy6L
qbg7cdQzuFxqX0VG/HSUZxb31yMOO8r+5XNNqUbhfmEqGcGcya92fdhF7lvX+6SF
04efNBZeGIS0nEOf+6iySk4l+mZhpuZp6raCoL67h1L7vmylvQmvWz78ZpjqcD4K
wYU6pj4tOrsH3TGJrO7b8+wLuShe9nWGAdboDRDhBQgG5hgyAGpLwNoO1aE734OR
ooJzRQc4iJ3ObDCLm0OD3el3RRRzASa/yLVJk8U2Qj3WhlEJHgdyRifQI7ZemhY2
qZW8DyxqI8qQl+LW37L9gynFKyB6hGi5si7k41Cbn7Mj++76qVi6Xninnnzf45+6
XkLJIeYLYwFY95TvbkKlU5wHASQ9UkwyP//OSaV/ziZRiX7tIKDWq+Sd4KpO7kl9
dfyDEuIyErFe0MHtlm3U0DmcyUYbYlPTqKiuGWFyDqQkvWQWj13NmEJhBGMfsrmU
TfvGhecp8SNr8Qy3DBiUrzgPLhdreC1LbPIeMlQQYo2BVBJiwIYebr4lZg311H+D
G5TCoxy+re+QqmIv3A4rOAKRxg3xurtR2GJA4mhbKYmf1r1Fd6kcqfYQAzLu1nfZ
RUc4Db6P1WVka0aiUFm9MS1wH3Reis2k29+s9nv4GtozoN5uJucRhUwLBY12a0kO
suVKhoLw11zKe6BxGTiSx2FQavm2mH7Aod+asue1da2NovUFknc+Aczp/xyf6u+U
PYjzQQM3qe1mK110Q0vEy+95cOJiRrRXmv7W6fxiM7ziwTLEG0xWlnTwinJOfniz
ah2SBRwpx3H6YxJIENbFJDWxU9ikMAg4aQEe2KXnsyu33K0AjBJOUoWxsiyvGpP/
i0mAAbuXn3O6yrpengMFJcMrbky58tq36haBx/W4JF2LXHaWskXjmqLSd/V0cXtf
msQDUL/OuiUzGh6ZeXDBT9kANpcJxFoNbGV/mnSLugjItVda9FHKA89XoSTBSY2m
odsQen6tLtTdAP3uzPQIci2Qm3V+wu3eYKsc5iw1V0G1sj/hzP/4X2ek5WpgtmDf
bYCjhrbUZQ1EMeN/Ujb/b6+K52g9MqPffyHWMmm4DqbAfyv5o7dPx/SoL4ZLw3Po
xE8Euu1Opx9RIiEUeLKiGsxQ3EwDgg4DQbW6k4fxHCVhDqG984noT2ZtBHT0EC8o
Ew/IBzik6OlATWx6oeZ6KB0csSoc0rXIXoTar215yPHqmbqcUgc3GFmSMo66LZX0
iRlam8xyTsoX56kYHmVKliHkg7phGlh4T/ZkYIvDRGcXdce8DY53KOjHl/gb22Qq
O3lmsBWgExkxQ7nmVekedpBBhJ6+INkgx5XnY+xM1eauThQhhnna5gn2xVbjP6Sq
ZFtmnzU1aLVMzJg1olCm1inuHnTThoYAk5p7KgAeKfQvHw5boSXPonsvMSsj0h8f
yu14vWsy9EGJtsChVyq4h350e8RUOM8c3zo3soNKtBEIuj19eqkJ/3twld57DYFD
WW1u/X2qapNTYf/Z4TAQOQlR3AbOifFfkB2rWZI70TdXnjH74Cfk6jkJ3Fd1mTQm
vRJMZBBtG2rwzkV+G0Ji18MPzOPQFNvIBasl8cmek6B50V4vdxBD+jgTQzpHGfBF
W+XLGQGIiKlZ7bFG7UxzSTMH83BT4bO6icIpRA5f/tvLAAX/4EVgpDNOYnVIB5BY
hcKA6YI2AgujHorIaCTKXGufoYvcJZupaAgpzYWaGGKX8lMQyL2utViAxo7+2I8e
SWscKlcZ3mAgWB2hOMP68l3yB0pEOYxYKagT/EBBfBkVwFo5oPVdfBS1DW5fuOwy
NNKw+qdidf4JQM1S5QIUSefxKZmF6usxSo8NzVbKMxZwLKpaEdu/viLwStRj2fK3
p49vTeC/NYzTcoEWU3AQxdS5dh1hqI4h/875GP4gjPCZFE6Mo1cca6QdhH+GssRz
XJvFK7zYkMtVSzYdgtL0TH2eQkxlITrCod53nnJt+N5I9ogxULNcdME7gfu+9GCO
RlT19dS5yYsaz/bsQKkq8p3FNA/TTpSQeHgvtAdiECCm6TZn4F6iDF/Kwr/jZw2+
jjL7VsLUqeHXwq4l22okLfwrnLMud/g/1g/GStkCGH3o1iRS4vn9y6jNlRYrUuIr
wv5vlYe4s6D6dJsIm4QI/CzEo9/QWFbzljjn+HD+Hq2YL/Mik+lhBcx5oZyO12kI
GOcRe3zhyHPCldwOpRlHWTHhKUigmXMm5oz8nSx469Vcs90bzzg+mwm2IQ3vCMUn
1nnLJMS6gZVLTsPDxV7uP9TVCa7SmjoBVLrOpBV65KXHMbZ5Jb29OX4o0DCUClGn
dIiFpjxnAglsd3HAh7VuTTe0QZLPl6DL8VeTKDlBRl13FwkHrgLNc0bGIn///TVI
cZNj27+uc6VMUQKbWArQcI7bKXiUDZSqAbCOu2GWvlFwikYByejyfa/i5vwAF91G
n5MY4sXBbPf/hnbCB2gbrjCYF/DUbEBSwhQYfpb25dvGmwIqX0xWBRtzKhHKL5Ks
nKAkRan9fZbPkCHcsQBsdt5UMO5hnnJljVAZnVB5khJkowt9m+wPXfuzWijJ9Cnc
e+cAGEtrUf7zHGRlBzbrGei/AQ3lPRyUwFN3X2Q1ROOSYilkupLtuvs7hl0sSxac
bm2m/rNW5Q1HfNRySMXBcBMPtJRfQsDbTdtdyHw1QlV+q3+mzsIaH9At957MWk5l
R3hP5MdnJcELaLUctEhCt1naCyaKuE11gxpndoPY0onGBdYpkuOdkjIRd2JNMGy9
h0K0VsENMnHFWifrXYmANGqGVw06NTE0qV9XlUyLK+AffdvLCxvWB9KNnQEG/Ex3
D30yNb9DqUPPmwPmpn4R9lHU1wW6O8oPMSD0Ld7Q3E5oqM+Buf/AgD55Vtm/2Fhq
ljVi1KqWuo0kUnmzNeP+f1A4gyRSwrFBn6efUewv5+K8vj0+nNimwz70NuDR/Q7z
huxaVSlt1M+Er/sNPI+Vi7seu5IA5/vr7fbHnM2HFfNue7bW/OtvCahYb32Lto5u
qbwws50lOyORXIs2DqurGL39DeQOCpKZr7bEbPlpsUOEKSIjsAwuj/vJRagu/ARg
Y4W8ElC/55+lAPj+ZIlwPsSTYn0aOSiYN/6nlNWWq4aISeUyHr3Afd2T+gaf/DMc
8WlhzKoMyxJsft+ggkoBCzwl+xystJvulkyctJAdC9zuWzh8fbeS+hsqVyVBQJtV
OIJ4Q5pVFUUPh8t9eodJcU+fq+aZihGKh4XNvEOQrN+kMVoio3mJaa9/n9LFlOjU
1DgJGg1mUegVuY/ijnI73mkFiAk66G6YmxKMVdEfo26a4m7R+CQCnP1P17qQJia4
heslLzC3/+ZARt8JJZ9hZS7/7viWjojWupZp8qwRN1UaK7KnZmGloWNo6Vt9AWiD
LQw7uvJ6n4McIbWFchOjfqnkXzd9mWLAddqNQjRc7/2ke4EdCp8g6d/skrFsJwxw
p4cjizYHyPcQoEqac7k8t8eyH56twBynIeztqX5Sr2sgsUYFAdphD4qHLgvqiwSh
LQUCyB3UMIG4vay63fP0DaQKf7ySc9zzQOHFQIB3fS2fLhGN6KdhLq9uQYFSaKWx
udAvmyYsWSgBTYBQ1DDavyKbM8b3MrRxA0gONzmjbZY3GO25lzeFY1a/CEjgtXgz
KhdstMiQ7JR9tDTYGRojPm8wTokKPrq13Kf1ocirTXi5E1Amq4qAhHdSXED7SUk7
zs8qQZ0brfFhgKkYUi+LhySvgqsNyxE6ad3fFYJq/UUKkf+IPzeP6eabDK9UIzYI
mAoZe53Hlqej2LZgUVJpLGuGwYJHxHZpomPe6aQ/KcOd2ioB+8qeQf5e/D9VE8vN
W5VogURIJJff569wI2zNe6X7OufI1fKBNNb1sJ+ApVSnYfmRbP7vQGdoNEgyzjMO
DtkSTu8n/Tzp6B+8fnM7J8/z9NN/hnYaqTvMfAH9MtVti5rdzeNV4+PU7k/LlJrt
k9+y/iEXKUizZRv7ahcVdKdkXoaHsUdQyX2kQF20dQmgvH5Y/ShSl9FAT6Q2D7Az
WMCuOLrjYq/BD5fr5+O5latgWGJjWnVgvr3voZ0hHwIU9eBucbld2B55esqZnvJl
CFTD4ppAn9fBW0xk3egfgJHz+HjHXLeN32HuELjzRe1coeGijaHY5n6HUiUKTIp3
Voy0X5q5f/8rKdD7qRLkZkBTp9x/ytkS/NSGFPOJakji+w+TUBPtiOBuJEMXErL+
poYZD5YnXOU7+GUZW38cgTr0Tc2ZHiBa9gvQSjiTJMyK9XG+Yy7vOF6RzqGjpiW+
CoJcBNN0GCTPxRp7dw0EcLt4pxcM9d2TM2EljaN091cyyL1Zt54VyGBv4F5D4zWF
NrDKTsJ7c0QIxON/3AUbUu/czgoMNPoqvUxjCrbMoazd+5HKWFzQ4q0anNISZCz3
4ZJsSDjzVhDZjRsUiUZ6E3n0VOZTOo9Q0I8t1EgYYXXN7UqgjAmH/z/yRPCz+p4j
Xyo0iuGJ0udAUDSmdQNMoyh9bBiCSgQlm/NDi2nIE7rHY16OVtNm5zXBhff/RQRK
28tgdubjlklM0hl7h5AtQ6/akIy5ynp9TAHizy2KY5oyNf97g4ube1imRCabO9Qh
m24rsBk7PgNYGzg8r4/jErnWhqrA6Ln4JYdiZUIQK+H6GF9uC7v6vPi2vYhjQn+z
6dXW97v0sKyvXUhFuFwNNylCk9oNJP2CVuBFOpedQvMtEDatsrrLhE9DxHm71i0U
fV+1aFHeMDhqfWWhlRZyWgAL2JNxBTYPwmZSV1k2l2pgJ/SWn0dZAwEwj48/GlqL
NB0lJpvVtivkA8E2ESzAbZG6KCw/9IaIcylxwL09JnZq9RPvm/QmYP4j6JC5d0eV
/GLPjJJ/CgZSy4qP8ZhNvKl/Gff4cfPgrJgtv4rACNSpD9DgdgQ8luAE6uCS/Zq2
N5Y3Gs7JWWCAxQ0ESFxzJ9zajABwhwrPEFfXTsMqyG9rNv4zTQW0geKlodt3JZJF
PfnkIFMM00wBmIJHLsItuRTVCVZF8ImS9LAWCHNWNpd+JGm0jvqbhqmV4mGj2hkk
sBxbxf+ZgDUjt9FKiSmXg3/+242OTedkPnHokM0RFHImRzdhMAZIffSfolfQQH7S
42FpFSjDAsOlsOWYCZ6qtnrUly1ktIw4c91GlLnHZv0yO3bTFbEXqSQrUuwpZW+z
Gw8avG0lwWfp648h+QQMdqQEzWc7V+R38viU7MloLkLLxZ62aYbjWavFIAEnGFtf
SGiwoc+orolVElI/mOx3ZiJ5OhCgXPMIV18xsRnzznWvZ8PpdW/EhXgi8BQ7UDQW
+CGPG2f1wOWVBoCJpOvyftiyHP9Reork77HWX23afzZe6oje3zZHg0rnMTnIA6sM
uDBcuq281a9h7t6pbEn2gIvGe0f6w96YnVTUG9jNXYLeGxsOpRh6J8TUB3MQV0Ny
qG4mIdrBNkgdhJQLlsUFKDxTAtZ/JD1sJeKUIaIoJ+FSBWGlwuE78hpVicfSIn7e
xg8Rmvwk+Xtb0XhiB16FgO2wD3wuRYn92U/ywgY+Dx/bH5K6g+uulVwGAGXDltUB
WbkZj1ZDN98HUBFdMXUAPx1QXNUwnXiNCiP9oDBB3w3CbZIMsfvjo9dQHlvy2PA6
YEJ/1bUEcmBNwXvOO2SLXOOp5/ZN7YVNtymeAMI43zMlS/hDDTCh363p97Bdbws0
paESjc3BxGOCd3nx08IRAo84Xm0rm/bDH4esE/0w21qwQS/GPlf04XSob4FpJOgi
U4rMgsgfLjaD8MO96FAFkF540im/WqexLySs+R3IAOqdeRu0zgvUBoG9Cry86cPg
SwH8lHK5ReY7+3JItJWlvhdTmb9m0is1pAI5evWgsOhfJktPADHRQ17kWmMGGI3w
ZZU4ujfWZv6IDU0hU7+hUCCLDXe1cU6HxABqC1aMZwJIKyXYd+4U4OLcob5PzRdG
FclDGJP3MbtAWwh/XxhbR12HtYqnpE3FE+pN9pds3sP7gP+ZYTkoHVUP8QjFg5oN
jiIf15V79569vWQtebQmRob9sHCl+Ibg2fXrnpt7h12jgBZE+jyRUnY6FcgBBMIj
icPPuVTLirJh4HV/DDR3h9Aziw5oBu4CQqyPpelywq4y9RGybPPPEl/4D4jyg9Ji
jdL9+AKvJYz2BDI7EWOPC3i8q3Y26sVJuHqw8gju/dgluK2LJpu+mYiFp+kKDex2
IHPdoqGGBZgV0mVPE6LRYIqZxa7GLX9REAZ1y0H0LIhnkXT0+1muaI5XBuKhaNcW
kq6+/OQFZhKEpiNM3lN00hBumDFMl6w5nkvgJhtNwuePT2k6o0g8v3L8sH4dw8v7
DFGMyrLXnbpKy5GqAAwAFgSWEUd92k8O+CC1FYw8bUhAcBTkIEjIqxN/ZFJcdiyK
OOv4dqDYXxtpslkMGQahxPxGMO9wKoKJGPQA+j1FuaG85jxD4Jeekujo16wnhk45
Ak3cCdWYfen8PIWxZMK4NfMsY+OrDtga26oDWhKyjueLtgVWgeXX2IguJvQuYE2P
PMAkuR/Ve7/+jqcpxnScOfReoEZEaw3ZKndBfD3bd6WH7foM2u7T4h3h2zWT+qA+
ZlsNN0F56VgvufRy277ks0PpHZVyM6Mp48yL70F/M6y9pN8eJgbC8JH8MreDizcE
oca/ZOdvQnMc2IDA2eYglIY8Seub1yz4jhwFgbNNxgNfrFTiJlP/14DHXx39HDma
om3tZu7+EExdoy0+VpXgMomxV2zoJZbyPd8GqYk04TVHTQEHhGn0jRFqKaQItkh0
wP/Q0WQp9VkSGLiStFEr5aupX95possL+kP7D/b9nyruwHe1aw+ddhn3GTeXTUDq
NQh4SAtPrdtPRIRBUgoWpXi2BxFNnwJuOX3l33EtK8aj5Y3z9FN/U89RdhzaWWBR
Qlte1hRS1Zwi0kmsOGJx7D0ZoYsgGexEpveVO69f3Z/bS3wIvnRzSTLMemamrsjE
SJVRElp0QZ48aA53GolEbIvz4GYmUJck1uuBfeDxJ4K/bcs6HLNJqB602uxzYo+7
dSU9xUS5SY4w9Z3lWMtiChlRHC5cY4O8urfr4KMUkhWZuSLuvhcZvyN7fKzY0Unu
tAUnOt4GlFLhrlenfzDaE7A8RkGgSszDMUgXFlua6mnkm/pMrAGKOGnb6f/Qkkxc
wYHiQjXI8N17wlD8mYzKp/wQ26AQFRaKUy+XxftbUryyO5TWeiSgE3II20kOq7lU
rvYHzRGnNCjC+VP4Mykk486+D5+bQkxuZr1OYS4/TlKyJf64kjKjLwvpsV5vWUwd
8lAIPrf/YZUPqvKbJpyfBhkwIakUIIjt9LfDTp8erGqL6Dj/7uG/5SszxLgp64a4
RZFNy2vcw17Fkyy4zTpVJQ3VO+GwQUm5xefekevqnXPuIgU+7P6nFXywS3r+C8LO
HjGCGTxsvX8RC0+Q7mwP9VQ+yJCNQdxE+7GaPGjj0C/g/r/sDVCHiaYSeYdPxv2o
67c8R8lVzinaGkunXY19pjNGf7+uVI7YjCtgTIsSUtqbjXZX1G4lZq2rSUQmao5a
hSpXlFSbAr5c84VzWuLDWcsWfXIJ6Vdzngkd0a28qWR+aLP9UUMMZKVKk7lh++Vc
BCkLWouiDFFmYJcoDOwCwYNavEOAdn5EquW2YR7SBcE/c9vflwN2cSBSo2dC9wiB
UmEK6TrASh9G12HAcHX9X5sF8NwPVFImfNOKZQPvLpPf3GBdfnmpbHavUMOwMfZz
4ZWNQkBmuyV43/NeNLVpkeDKtREsE1rrXOPUK10jecmOv5H2RAdmcTjmVC2qouk1
zW7q2vlLV9vB0BBrCeGLu5a0fHmXJGeasiLn4Omw20ha/k3cFR5Azqly2uTbhAfa
j9+udY4dIMwTh8TRpFqDXsBQ36ZNERaO8ZHYtcmYu6OTRyTpITn37Ap9WMNRa+JJ
1IFtIa16u8E5GyhD6/vO9w1/gAbXUAPJdoGdYeVq465G26X3ZLX1wMpean1G9eYB
WXtcPxSiAyo1fXEpmlSO6QhrvKNZz4kYzCiili9+q27CQC3tky0wVg2W2Vl0vKx1
1UV7ElBwQrugDUg5KIYm0JUpNq3L/jOAsVKJLRwmKcdSb88w+vqikfrtN/4tFBRJ
ZofVLeF0L9fwcl82x1k/V2nFO1tGCgGxxck9cUWtL8wphPhtiMipWkkOf9qtV4Pj
LRPaQNLNACLwDtLGXRgKUNxzurV/VUPNNYeE89Pp1Wk0I459GW3r/Pb/p39przor
yoDlPF/xVjbhiEQWQx/lexkDltN8uSSBeE+PmcRhgJ4YIDyuR8akZKDTsGP8p+at
gkOYhRTT3y1kAPSBi/zrMh7xKObNNinyGC5UC1uBS1/x9sBm0GPjYgmce6NDMgyx
xjP6I4lRQOWnK+hEEhzFrEU0SSxwr39fHKKBDy+mZJVjBckwS/VJk0gpKYnrlpYK
5eV6zHi+bxPexIP/iaF04P7CcyhvnMIj5u08vV+ZfVEyGgtfN4zjVsN2UkTbJ8uR
pGZHyXJJugcBmohTyGbRv5Aq9H/vunvSuw9GM3ZxwL2BxV8aFPVrUj2q4R54rfXZ
SQss7RV5KJxL9ylm8aG1v+jfrVq6VdRyuIYUGicFFPuoOjLq1pAMOFXpKTekyk/w
B+HguylJmswGYsqAmqUREDCQRwEJeve67qC01S5HPemPbmJRsd+Q1MRQA/VoDDyW
9NdS/Ea3Bwda9CJB7u9gjJHSNAdhZ+W5CrAm9dwD/ZYNbcMbe3ifKbYc+euR1j6N
h7BSd+Mk+tACgk/FvkpxJdEAItel828i2RRi8ReexkBIdLWXSjrJocSthJW/t2E9
kuFfyzwsiqo3Z6cCgMPnJNaf+eDjywMGgXX7WlC8DJIvfhDcXBbHTKJTmNElobT7
AQMxTQFtI8FdLexsaz4Zy0sn35ufee2pwa4iAujZ8T4hkLfTy0W+uyhcaNvvC+Tp
yLtlmYatIOPnkuE/4TI5HEpLfxTRy3GmihUnNX3Z9gkMDDUxd/zGgarnz7YI56l2
iGsqasQtlXCUBS8b6KBZ3Cd2hkIkNPPzzw5zH/fsfefefDeZ5OEO1SA3uVRDO1a7
x7czHs9ZVvXitv+WE6kIIun++5If5Ecivvo/MENHq2sPlxQCTQqT+LGwjbJzmVzX
L0z1LURwyOzRnt+Gocu2EC8QLJnGbAU+QxWDlpxaD0wojCch70g1CdOJWWCeMLLp
NoS7t8GdThBx9zEyrBPTV47t3OQm/6Shmpv8QYXlPtxKSO/jI+q3q3Mohjvagt/T
8e1KIhB9GYsLVVLeFfJEaHrnxT0NJ5EZZP0qyLqMZByBVkQ9bOCebVN82wNnNxRd
a6+/dWfxEx7ja/Ewo9OTZMJ1wIrfRWvOJ3tgJTwVLzVUWlvK4TyWn1kBjgONN+DA
JDtSNtcU5U0JmssjHW0570zb/XKtI49nd6TeahiZ6rRRuglLBzSQJrK7jUFg6a+Q
WXLAW4UAgP4qNZTwDQDDkr8/PEEUQ/+6V7s08I6irF/NmT1mRc5G3jCyg/R0obSp
CHdMjbg0b69kXGopiJs7hniTCIW2RmTpwYH8aFg2vougdn0s5P/23z1RfE13rypN
phCOJj7TXttwoyuhDc6BPhwNRZYOyWqIkBKjcxkyW/PK5SkmnVjuCC/K6Az48B+Q
QNZrR9zVdKfhzDXHoAYX32DhG99p8tYovUAhzpW5TZQEBBpVn22ofDLWUOlEIQX9
+C9GdKUUuDhW8QWBlTDRiveN2EylOh8IZunjoDnbR4ndcU1tcG2U8nHLh77lja10
tsW8WhdZ8oIHLz7ANGtiFnSA6Flc+DTl5eDe2fgTeYXl0WU58yYeIg+Fx6TFEoLK
F0rOZRPwY0u8TFjznx5VGiTSyjkwC6BF6GoLyVpCU43ZAGN6s1SBnOMv2MBxsVMG
pEpPZ/lFdJ5XOivcpFvFDVKJ/x48twsHLmyzEo7BDJBM9AKSTQ8lTTk8yn7CDN2T
sQfuc3K5pKU6bfE6jacv2hrBaWq15ZEOritOoRvCvlO8J058OQmxMhapQRTaUzPY
1Kl1Ln1pkdcTyirtukFBMtduUolpYKxBNSaZrFDjw+fvcRLaG2p8o+txXtb7JXdY
ibevoqWlE9ePGk9zTpxH5a4GN0OZ9FNCVQFrEs97lPUzVlNtyevdswOI8N6g7kBg
faQi3IwgfPQNx8hTMPW7je9/UBMb92MSgMXH1842IuymE9No5xWSzk8UmxQKwP9E
ZWDeJLT9i6isRpMz1LXdSv/JB7x7fgs7rVuQBnYfIrbfyDoXF26uD0wDLvGDZTL1
jwC/etG6u2gG3QCq8JyvlKUG7Yzae3L3NwJP7DY4lNQRFH+MoVS8JkshIP8yCsHk
H9AReyPK9RD+kWO9pDEJiAnr/DE4o98m8f3mFWJn5Jj2BDIgOdSBApksaMbMQnwU
pl/QKXURKEPRh+0Lg6uGN5hjGvSZ8yN/eyoLlh7vyAlukeCO+8Q7VCJ+fKKSy9Gm
k68hYAiuZwrdBdkX+x5f9z0H+M8X964uIJnlZMmJrhtIQXsEJLvVcXzsGvsD4b/A
sl/SilW5NEJGBNfe0a1xjfRq4NkEU2UHvTQD03jlq/A5qyRfoM4TnWlOVytRosWz
6swW9qltNIQ+ibxKeNpNcaqDKtUMhj9kRrH/FJNF8TA/WFBAud6M9NwHw6/JvyDc
yYD9HjQaDaOYdcM/MQihpT+/p8dtT3TLEndveRQCS8UehJv2/SAKLMiynmffWXBh
hFm2cm8BRY6kQonyT4pxKeWtIQzO+dxk8LgWT7UoBzNLys2VnWoVkxgo+AKj3t/Y
PyuwrD9Oq6CtEMi78GJNNC7cV9g4MKZTzJLPJuvQiXLrx3fbbCB1yRng1Q8S+Tnz
7MPyJZ7TO43KALng/hhbFh67Wl8mZIqiM1QacnxzWc1yAbrQz3l0sJima1euXdwU
FUiwIttesE2e7s8O9szZmvbgOub15h40jHbQcSKd2Lu3V79jY8vhgLjIJhGfw01+
uaEztLVOnCZRVYsxF9eF0bfOOPSBs/s9xQD4AtJmArpPxtV7U7DVTsUXM7xFx8FI
KMgDcfbGhqfI7hXThGAzlIfqFYPS4N+R+4qLDu2vLJoqxbizBVSG0QytKuZmufMu
mHE3K3eATbF30olUrOyh+MsDpY1ufSq94TW8s/g7Prn0Qmy0S+eK9sLLl34YiLch
gZLKF7gf1yTx+ngQ5hTfxGIQDt0Jc5H+z2bCNs3m2Iy2RVZyBf7e8DCXHA/VndvF
BwntrjATGjM8JUJfM3pk1C5LZK709UqW3rQwOIqRFjhg/GcbuXkK1EOsDfYduyDV
mNHhrDwmkrdYRta4u8AA6cGmCOZtYG3DrnhO/dJr12+/P8qHPPjKHyZz7g0PwwR7
rbWCebLi/O2v0AWFm2eaJ4nzBJWF77ZW7R+82JhkZWo4atiWxEEOJdXVwCoLf5uC
6Jv8BFa1v0JaQgJNaX5bRDB3+LOrq6BtskjTQFdWA+MmawiudgnHE9pqgauT3Os8
L3IPpNGnbOXPZ7Tho8b9lQhs8sVaHBVCgjdbbisPKmQ32LKv7S1kRMr2RNpDjygM
J7gDlUNkvHQal/NARjl6UTj4RJJyTwOl5BciR9i4zTR1qo8hzuCUQgiupC3f/IZx
lBHaudYp33slCn7Pse9nySRZJKO0zTFoyshJBIXhZ8iZyGWUae+j5rCMvs5OMLKo
fGzje44qHT331fagES9DZsxmIwAO9ees9JmGDRz5MOYBO2Lrf7/OTGVB083YdK/L
w9aedq2nkVQa13zdDaPCxIJPduA9kylQ9yt1Ls+xZYHszsmXMwFEahATYrWD7XAG
CE2dnma+53iiT3raEeVchWNYf9BO4LsKUpVLHYNHMOEUdWPvX+DkOMl6Qa65i2Ak
ChHYehpfGXDxJRZom3LV1b4uYyfAEtA7LNYc0khKhGsuywn8kZGxXtE81moGi4Es
8xuDHz+iEe1O1shWwDUVhmv/icKxAHX2bs2ueiVesvXiheOWqXcOdj9/HWbre/tg
8q29+LGNwGsrCFAz+eGJtWVars/aXXiRNcy11qhuH1ERsQIF9t9DoYh73hxzvtP5
cR478RIGkfP1TWYguOg+47nb1UppYob33k5UPhxEY3YHRb0K7fJsS/KjCEWht3vn
PB/xCduYRTIn5kg3O9D3QGjh8ORocE4SqEor/31TjM4FuLTs4BniPpXWa57hqZLo
L9xNAz6gCeUHvc0VMdmmpmrR9N70axJfpSFmUAO2N0+jAcGtEAYoyHWiKB5+SUby
JnfdLBZRn9pkNaBdcspb1AxfnQRhzJoASyXO2LsNADMjA/F4BiVVdDfQdKvgKXuq
sIgfQs3oPraDTxaAV59vcFch2N4JsCIa2wXU+9ZWSQ39EM7WiN7gkWLGydNX85QV
XH66M49VRbU+kHM3voNVefbzrZHV54wzhkRkDRTj6oqCKFAWxvQpv76CNKt0VDN9
wLeDrKEiST3B1r1pRdYgwRQ2xfD6S0dJn/ijO/gQuQTWNmHJXicsxAKdyZWvv9ln
6aFRD7bReOA3/BRcfhzBGZlbjebDJq5WGY+se02U+5FqRmizr5p/YlM3CTKfLAD1
T14gCKwJCkVKsYYyDKYTcvG/FG0WAqvzx40H2oVlqodBErr2xvVJq94L64kFsaPK
S9dBeAvjPxmouk7ED0K6tf0uAC3NuiYWQQE5PIt0zyRUCB3pbzE1aPe6+14mWYQW
is+EO7InnemS1a9Uh9KW+kUGz+grmgQFHLywzeIhBCo7iJU0tIh1Tj9MvYAPHZCe
xSg3H0FPGbsKH8AGuT6OxrdpbZbga6uK8E7NeVx6vkLnhKKlRwdEOYgcfQEDlBj+
+eQjNm5qu1uBieHGGshV0PytfIa9TS6gP59CEpD/y7aC7pknvpv3VTiYydluSZYH
UiwZ2n8v4XqCQ2Kx8GVw2WdQA0P+sNyh0Q5qdztELGLQTTwKOSZQ7rSgBnhxF6TJ
88x4iXy3iIziXjK0xXaSYNJ6JSZf4AlsfGDi5owb0lrBQcM38Uax5n32VMDUVv/8
nUjgFNwZGcjOAGBQKsqTkpVyNigEHeZzBvcan4+3HYl/bj4LD9Tq0aRNA9dt8U/z
JyQz0sLTZQy+qKo9grMCLeDM5AFP9JkC1AIUv1sa0LtCq77PQq/9HxqmuYoT5+ai
XD/oTDpIsPD2g5M3dbVtoGt0QL8hoYy90rsGCCDkTSy2ps768r6dsOPppMpQSjkc
4iWXHu8aBeCxRhEJLM6gq22ufDx8K/05f2PNRadLNgZy3qWJPnnANrGIkBwVNv2V
knA8m3vueM/MGoBz3EUOMGBxIyFVjnQhgM7UrTQnlNA3mBMUvDmyJDW9rEYFvnpT
gkONxHvEPpjJX6XpKSACAi+79BIqESyZH+IpuJ7nXSo3RMNhollbpCygfYw6eVRj
F3/F5oGvF9BVUTy1xAMnyqH5XyKTRMWYvCtCb4mB2xBm7LUCOWFOu2lwhaKYhxH9
5uJUVvkVcIW2DFNz4cCrHfJjxGFt6GvHa+xB1n9ZfIp+5zZp0pVhYEb1mUfX8G5d
Qwg2wwDwOUQwyipGj2nLLRZ0B6t9nQDCqp9P4WfT3sZ7m4bA2iOsrhDae3UkYc++
8qJjQkLFFMDaOXKQScwsvLb7j99NsflqNlabgV0HmNnA4H0BE6JFEux7npyh7Naq
BO0pvBzWUfbaiFY46//WpFbayuyeXiWeqLk/aUgHXTKMKKXKip70s4oEz1i9jwBD
WYw9tA8ckIL7p+/pP09aUORlyEB6+igjjiSWyM+jgRpXBhK1GwiLADG1/qMntlTN
XBRZD1wHFgxnQZl7B8WQgK0G/I5jO7wviLy4EdYSn6z7rNiNyFISxGYahDhf+uQc
S4LmWHPuLrIpquMkVbAIpQ4mFjzkjcBd9mz+wv9PAoL2GODaFIOONPmMbnW1E5tv
BRYDQCqpYd09zrw118ZaCJhLNsMTLRdtHKVgRrE4nOm/fhRqgcrP9hiBSXgVAl3+
3h5kVuLH0dAWJDqGOTLsKPKzkKK2V/dA5JwhV1HlIvjTGzm5VpVqYyZ4PLUBZm8r
28cDGIsax0ZRClheGTuvkfbvH8xc/ScOftiEGXPBqNstekB5Fmep/n+79mE/Uk73
lGKoHZcVCLqPUIu4rU7TW3aXZSFDKM5LAYz/PGBZVPZgTGWeoSQy7ojTjFbOHMJp
yjeKu8+Sx9FN9xw80V7t+jg+cHVyuwoJ0pzWPv2PjRQu/GhWijkRq+4xO7zqW908
1x20NZ3DUtxhADdaLB+r6DgeWin3ISpvNrRRoquCMm6yUk14hgabitL84wbUuhOY
BXPRVcjqr5jGtK9VGhOaolETx6iuXvZZ+YZXi68JZs28525H0fwCzGHeX2/36scu
bh/yNYarRNEkE2RNjL80Q6l18wpdha4+JeR0K5t7DGCTcU4WCERQdEhyG+yaiKm/
hU5UnCiJLlXZlyYdPI5mfhSIK272LlyNn/H/NJs7ie8yOglU3qs4LtKogApzVTYK
aA+ktf/1LyQcXZNclYFKpPaw0AsDVuJ3QWCjo0er9ObCRXF6qvfCsPvJ1aWs/Lyq
LrbDzT+hgUiWywAM4UA+0mxCBy3MxXLn5dQQuuR3fpFizN6NQ1f7tBMAO/MmcD7o
6htRfuMxr5FvOtKvS/wX+8bGW9WGQSk7p7cTSKYjt2nvlhXnMh1b9CDw+Z5AFK82
xwqoxwa+0a5TH44Cx/W1iSsnjwJOW/X9iznuI9cUfeuI5q36fGsEz4JZcCFwt3Yl
WAuw7meQLJzhTKD/sZXeZNzlXS3zvd87mfAo3l4thozMYXz+DkpbJtdrCKmpOdEP
PQ2TDAO2NYf1yRHkQwHyQeZpGu5cbZ5ZHaz2DliWgGH/TYhNIvarxqesBwG016SO
0CljdEq05UCuekmga0XSkI9N6kCC+LhvINrzOaf/oBHz3rAxy7tiJ0YlsKVwGNxs
o499AVWI0VQ73P+dwq/R7Doz0P7czzwNMAaokeoRWLK3Nz7fGE8xF+7pZV9623Ts
FEO+lOgD3Rey9RZZSEzzxRwprQiUsRF7E+kiBH3L/SJeLkVxFI0qanSjKyKOM+CD
d4+FP5KYfH+5WUiREX8Kc7DVgDjBLmm34R0fUfi2bgbGi2QLnwWR8SohC5xjXIFl
UXhSmZ01L67eB5pW3qg6IKYMmv0ZCcPuH3cH+7U7e1UDqU1c9xfsykzIu53462rR
pX/VH4yuaUL7LZAfkTRj5kvaASxig679kR3SC7avouoMyYJc9mrfQXhjCEfSPNnr
tJ8U28nIxaF4/r1X/K9sct9HU3REEfwh00Wk89U5txL/KbQ69DKt6dBqEZMXhjtE
tMiSLpIfk2A3/R0GgnfdDjD7AF2xgYvVCt/Hm6UMDBsx4cmpePqbO/6Zj3zOJtR6
pRRGTFQcSxy616uAevt08pNvwPkoDQ9tDBseEWHNyGoEWYKyLZ9RAAokrl4soagB
W22v1bYMoslWEZoQbCRudiN80gZyQNg9AcUvopptQZ5VXarbaEXnt92iNq7O1mGD
J1npDzOrjaF36AsxOOoPwt1YHU2I2+6mItga3N/UFigEjppipDyhingAGj0QT31o
r/XAP6BN327+eySMO55VmfZUq5m9ep3YL9r3ZQdDMQA7LNjQ3kKvVFdhkUVko4+E
O2W8XHp4BesDc4fQDQxj9EHNo/WF9KactXf6yYcO39jUf9sMkZjkW0XPloSCtrE3
Qv35McVb6p8EzbnUU2pjXigeAbUH0Gptabcw4KscXJU0BTp4gYZXzSvscubtMbhO
q8A3Bbg3y1R/QJIYJmd2qPBcw5r+gnG/8fVq9UlMc4Pq8KkIC3AH04mCI0qwEQGo
aluhTUPRz2/hk5Ri5JqjH8IkqG05NFyyxh11PGqUDOp3DngS3LZD6ZXSGSV9ANJB
LzuYsEE8K+rbU2tKIXmuflBUQ0L2rX/jSH2hmfE5uDYO6KxNsu/kx3xdg88Ekbtz
9PrhPiD/5ugR6uuVhEsiZqp33LbaXwqSobh6vqRh660vCin+RdnNgLUDTHKE/aLW
nDRagayGCXwObb+JhkgYG0ZCpxpOhhoswjfzuuiW3Yf94imLSLFnvLY8oD4EdeTj
VBHJIa7qvqiu3sI7RnuOp6abjF5dB/PioZ5e7zQmKrRxzCW3mc8x9efie3O/rqGT
r5ifqn1aFFkXjnYqx1YEn2RQ0U1R2K5++E7BgW2DmfiS+Fw/NA5M7TWFhJKaEOln
QD2VjclJ9gPvH+Ik44owSHKtSIGDYKy5I31Ryq5cGDIhJSSUPsCZjUL5IDfCvOd0
3sXpUDqwKsDtNI0h7moYR8H4PqF3fiUlirEqRqhh47zFeNE4RvpQy5FIKDxtsJsk
LwcmWzpXR2XEqFiMy1xJbJyoJjbzFcG1NtOwB3cKo+tvetu6ncgoFwunj/BWxK2m
y1gtn/K+on+Z3uDJxCHOiF+LOs0xixK0+Slu4TZG4Yrr0a6BOmQqqS10z+Cdithd
CJsLzVZB4V/R1v0uVXzOu/ydSC7X8Kk7qoeBonlSfp54dBn/HJ2lnhytj3WyoHAC
foi2OmxgiYRs782RIzmr9Fg2tM5nL1zZ40zDZ16wAtP9X/GrMQMIQOwL8SjKyJZd
ujdQal+B0pArodWGVMsM3cAMFhy0CxkkKapNJlUgSYADcQu1LMrlbjfnwrZPmpz+
pEwtnb9PbRpz/8ZQZyRZSq+kVEOB18WUHtzBDyzYOq2en+6MyEEGhgKwK0pbk+El
y5A9sDZqNkehzFdlYytgSZ8UOb07PoQp7GV4kZVhQEboTlaEtVPSRmCwMLcMS1kI
TbHvqP1dQHSiWCxDe/xSksFMi2fuYM8QAnGeZG8apBpXHDkaAsKlGSO9uZ1yhVv9
qwQpdGe/40x7TTUzSaQc9A==
`pragma protect end_protected
